

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
JtfK/+1JKYw3I976gLBlwV2xqGRbyVsJ3RDvlPNJRewqWZOfwn5MuTyc+U7c7Y8NUZJKZ6RY1Q/g
uXt328ut4g==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
SKJFICLwrmXfYqYNdiUThnnX5tJzUEdqxXF+PdKpwSGA61whpH8w+itTbLnn6xyBye2kcWPZGi5e
86BY4EjHm7kmXxm6GHfc5MWAMFduB72GxoAF5LRKlUMCOdVsZag78zFjXdMU64ClBQ4zjB8EgXvA
zXBqthWa876wjTEo86w=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Ho0WiFevcJjvoEEaYGtHkcW737RD7c5clzugQBBm9an3ZkyNmpivYZbh5x9redNVt0HOAIz4unf2
BSVy7qVCwKIsJQlB2q0JzVYTIfuco8FlNbrUR7/BeLSPV7XOk/MTxR/0Dg6meFJjnWuC3OrBGp8S
Ul4C2x7zg4t68SLTuFe/LzPmogzBzDfD3+nozb8sS3jX7ZaQAm/T/7eoy3grLVkFjUg9uj1IhVTP
59FDPnvyx1zZ/V9kzMjvM4XKEW4i0DGLbDEkqT5cZNTgcxi+sBHO7OnQuIvFzoIoNFONwh8iJ8xI
jfha3bFVgIjIJWFL/KzL8e9Uwq67H4YDz6GAsg==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
tPUgwDCRFsMzMdJqCXSx12cw+CNwvndABCoiKOSYIqrjgxTgSZ1CAyY61ekJUz6cu1q3fnTmoaAx
Nh8wOKV+UbnkqjbXLltbzNbjSEawEnAI8RSn8gStXvDoHe7R6pRqYg2wbvEPk6N6UhaMjVC8JxUE
Nl+LL/ApnNDqgvTWrcs=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
EyCeFS/0OQO1er1RAmOJ0VIpIQN1auXP1dzcGUAOeSe9eyc/jA1mhBpZ1JPfDCNxALRFgLLGYZec
wCmtwGwTJ9NXiyrouRmXyaKsTpp21jNq9KLTxpWtw00JZFdcekT3NPcfNHa7nkycvsM6yWSUR/cD
frws/8FBuaG+siAqTh5qClTqkxCmbJ08Qh/l3c/D5bCXbr8wXY+SVe6EK7TiYFpV2oOMuwWw5VVW
3m3/ZK4knJ1G5Nn68ZhcGx6rqQE9ZbHMigIgQyt/y7vXemBfmAZ3xkMsYj2X3k1fFfReGPYzTOCE
6J8z+FWVfzx6XMFACHDbKayB8gE3RAvjSqIISg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 7056)
`protect data_block
PazGmhHjdES2Gmzvxkif1CT59Rt44TIsBaupHD7ii6a51oROjSHDu+HEGyL9UYQERs8jk4I/TEAG
oq7n8sJ/eS63aYmVQm/vfl5X2CGKkCsyH9hVoxo4wt6HwKRkz8GoM9zh95jqzMmMBty5tBokbYFh
v9N9HnVhJVDFTtn3wGy2Vtj3FNEIWLj0q7agbjDn/U7pGdOfTzyyr47LLxLBW5Ea+mM4IZDs+NHG
DPg8R20SzerBjToQlwaUvZPkhtHm8ccY0sy4+yr8pjp4C7nlZ6+CrkdAW9EGSvazMy3T5GZBUmbX
SmN/XcEnto86KpSN3tTMg+rhpnTmnDyinLVotkRNbN0xRmTW+hGK0c2QNaCch8bv80t843yEtL62
6aN5NA7DYq4/4qw1CbjzllliBRpcykMKxAszQ5yf643RZoelapM3zgbiXxVs3r9gqkF/RcXQV9jD
s9RclPeNHZB7JxZtuHxx7Ga9wOJ1NwZ/f+W8c0B9yRy+XEyBdmnyp/oRi5nvK+pFenatd+w4aYoY
2Y0oh7k/xmeMjA7IyHE5bSALa71zB9ceWpRw44YD32jvnoPBCjeonBLKn94cOn9Wf3ftNdve5MyH
red4uTB/6MobcoF8aSWGPT88xFt01ugH0TfSwUWN/4ZnBcYLBht4/vAElw+URNJH5vHyypTtt7Bj
olAuQB6Kn4Tp4ZtHx2YprhR1a15zDOiHzybkcwEZABI5j3/9Fg12DW31jvM0z5u1nnyszScDRsq+
11WnaJpQ6mLrYyGaJS0O4T4FPWhUwkIBleAiGQ+Pl3rHQtkIEi7ZrnyYUxpFwkGoCaHUkK3swnv/
l6kWggA/4b97bhwPdVMRNkTPTeJm+YA9e4pWIGPWAU9gWxdp7xYdgFPetClIImK03s7v6tN6P6Hr
6SmyySPF3j2oAC1zhlwXpZaxCQiiGGIJDKcRH/gafNjguixC5G5d4qO3n1INsmr1U6qwsK3R3Y5M
UvIklH+KdmyoObT30uSD+XsAUx9B8yjW77AQJnJ4I5Iw7m0rUH6hojBnETwCAxre+6iS6YyJN5rk
Gc0vTdcl6VzOsyfo+rQf5r8QfgJh31Hl+dtFQSKCw51jVKDLKYOFfhVrvBG4xlSojUiyFNgYWCfi
zgt5M1eIB8ABE1SqR8StO4YTVEstXGI1lwg+yAUY2gtOgHsTVkpjhaOY1zl8PvDwCKU9dtR6egbs
cENyU4AqkKvIpAMZ1NJ30SDDh1vEpJyOhn3ykHHkFUiYTGxpvLubMlijYCtRvuSYf93kfPGgIAS6
mJxHgT0XZzJe6tDELKlm+Thl0kD4vQu4fbYXk79VP/9j4covaYpWoCa5cmLYKevJYSZnsDYnltX5
fDqNdPYyjRgb9tWsrqVhrlvL4/Z3qY4IZBkJXXdVGa3mazxPB5/9RawV55MWHoXbLdogG0huophN
nd08P2cjYCelrIjBusXjcgYLBPRYBDz7eT3k9Uke9jQYON4Ab5MPpL0NhJho4/dNYmxztjVY5EvC
GQG64qKF8NhycGmWjAJlVM9b7fueA6V2mWCWyT6WdTID2cdPU2DOJbnHZx7ES1osV3Apm0gTVBr6
5X5TAxT553sTmhPwXObOzX/Gkp8R8ExU5HgOXQMPninLgl+8++RiBkZNY1Ygf3n8lpELpIEGxC0j
FJEN4JcXwwvR+PhRHafEmRaNpcaYPF1ntU7+Q3BGia3EbpPALk/eK0fRPEDJ7Wz49ewQ7VGWIdjj
5F7IQ9Ae9LoIBzUOU2kUMy0X+rTpoAbQvdutq4H0f/Xl0ZzT7OASPyY8g5Kb8q03jHTHwGkp/wJ6
f2ziKcWB7wbTrH67dbLWy6p/s+GYboeEpUKq9sgY67JKblYNnouwYzzT1BqZHyxxP8iGNOih2ZH4
9hfAOtYNyPGiLsG94lLRjeD36WEJQlZ2BpUUv1WGzv7ipSB6HxTMMi5ZAYYF5D/+OJBxj9JKeBuf
wZyhVZgYx65kVsEDezmU6CsH9e4dIHzq3wc2kueCH7Mnyx/a63P7iYEM5zrN0un9uEUHnCwcu87n
pZjj5qMP27XckdBU54KM23ES6H2he/sO2gOf3O7o/yIO5/Kxcw9P7qjsi8DD700jmQ47LTJ05kdj
J7DZcRbWkxpBy9T0UY8pujXLtg0zt1vp5T4Pn3eZZ116VAYuYEPUWCVn5Lju2xqjvymVMg0nUpbM
BCBsgHAG7Rv0BJG9BFn2+qbmx5RaJByCdfl5g96sAKu27KnPXkA/gkhs+Hz641qX+ygm8OnTdbLz
V+KrDQ7Slz8WVMholPcNiGm1OZWZ1vVjspQvom/Z8jfO2+bIDC/JPcCLrgfAWeppCVRikHucftQz
3qVN3/+93O3AeHL4tY3c1MPwoiVDm5dqitP3NXzfpE+It9OmiyMrFm5bzMiasNyKrBts9rcdU/IL
2Xx0afz4NbfAnR2yeSkg+gAHCvZW1FCil5fOgq8j6mjySk7SJfyPzoDCzp3yzH3k6w3CvXWiJfMS
aiVvT/+YdrRhmskqhc0hLYgQTvX34xT5dt0GR7GNB6gfZQ3Ifn7wjrt9I0UvLKFuPm0/VgJLQhoQ
sjd7C2H0TfMdfqeexCE9DGxDssXntd2BHaYVmVNQD+qiHtHil6aYwG4HgpRLXbg0N3vAMxzs3wgx
Rfcn+ahSXxkmDsQnnrVPBTZyg9pLESbG3ONN9qnFm3pjx8GFpFTcIQwYa3E83SszPcAdIXnHUEcO
ruGb+Oo9IwD2YU5+aIERITpd2XJOc5hYT1qysRNe6hONqR32aBZuFwRdntSuYhdRNFj1djBQAyPa
y9Yx/bln95VfThTNwjM+jmucAkbo4JOT056DLh0lncar8+GRxVgPaYsoxZysQZDhnzlukjAJvAeD
JqzMHCpFGI2qHzQhxex+9NHWSzeYlgnAuE0sNwYsDuPclq4zAQOKzHCsuGWas3a4eSqd/Xyalb9z
dByr9ld5ObJOOHVI0Z0CgnRcuZhsWnMPcfl6MW8oiSr3T7CVxV/AwvPnASWFYO0uMYPyXXw4V8Xb
HXM5CGqEqUpW2ptwMpliq22mRRnKM3y7EycbpMQwvisvdTb5KEvsqjs43AAmrTMls1Ce7ydFkJBX
hK5ZaUV1uHB28hcvLsJS8SN+oDXfbB7NBUn/iSSHm7Q0c7FLYy+6uF3zyYhIE6rR/gDTdJTepQDW
ZPpmgoVBldCWcLpd60HFCQImb3+Tr5XRRYMRxvoq4OdrUVt6vnApnVDCScKRSXrOzUenOilYjMLs
hmmN+8FnCpApplSUG6rLXjawUPdp6nqK/TqazFXKMrlwQhcTQ7PmGjr2+Hse3wWtsoNmKrEajSHl
xrieNZs2iuj+P3dun0CCsC9HJJAFvtsPK+QCVgMJ+62ppuBcukNR8/TnATqXqZnFbWHh1jR/3jWc
eVfwWIwE00eEMQ2OEgv7oS2K8folcJoiamD4QbJ8eDqroI8UfH3nGJUDlitFmZraVGtheIcg+W7C
/BKznX2U+/34UlzixB5a3ELCeC2ScFoSnbtBrKeVAU9gTN/deMpmAMfcgF3B56rjE70TrVroH7wp
Uv/VVkrDnlbPPIxepMW9XS7/9YSBq4W30LW4Mra877coJV4sVwe2MTSO35kLOtVeEYqIEe2VjFIo
Y/at87OOD3mtKe2id/Fpl/i4Z7gDkvgaTv6hb76whG1GHsamLeW/i2HZNFshC8vB2lIEKcFahwtF
PN4piyz/mXq3j3LZ0Q/ZpXHoddvJYdyzgZbYzgVjAL1zCGAJUrct5313uVfPsTz7ZUxhYh8NaEef
FCdriaPFjf8EVGBL3bIjUCn7B+pUGm3ieRv83ANTlp2XddcbrgrlqiDYBhm7zCbo9bCjmWnD9Y3T
lpNx0piHO1qu+x4h7jSSLDC//Gm4LHBhlmC+uU4srdlsyNFt6Mw80MyRIi66s8l76b28APdqYjUy
NOa0gv0AI7pXyvwPguf3v72TEZl97pBbZJaD22gF5e4bcguf6cUgAtHoylioUk74DlznbRIzzw/S
0sm6wa70IbRhELHu24sJjCAI4emzaOpjrQ+lO+DigoH58H/LAjvv8FsW6Cb9X++Hh50wLtoO4jqd
HSstaHh+fzB31Br3iXiQwm6091ZowN701A3VxvX5AyrKXLbOdBwr/pS1pn3dVCRzLiCGB2KxjzlM
Wu5g2K7BoqNdTsB0GmITkSbJUJof4T8HkXyoj62GKn69s6LrQSeq1w4iR/1LC1xVyK9OpRR0seTF
YZtcQ3CIflpwSb3ysugx3evsJ+BKH+YbxQaWGYCkFhrOukEehpaKebzPmFPr3GsEd9vHDAkMuTFD
YtMyeYJvZE8piLhydScJCezzlAsx1G8auASts8J96cT2yMhXfgN+8DN53QYSE1WOAs6fdc1IdaKh
Q3rXQqQr0HpLmZRkT3RTRvrnQLoweMWq+0gO8L/G7LO3CBXOB3wO1XVjNbJUYb4wnUu3fpvxULjT
WG5WctpfJes8TC555YB7QHEu4zkXr1UNeFig7gOzce6Z8Wp6+2VGb9M0ETznpNw4uQVroPzzubZH
VwLWeGLxBFNeJlOjUtlxg83sz9C1Q6hNTdHQ/a+rFI7zXqIkY56wPOJ1v2875aeApl+xyKDHxTGT
nAM3pi9bFd8dDzQROw/qs4GpHtkDIp1OGMmYBJAFYz3hl76jUdKnqT93vA17js3u0MSQ3Q6ROPau
NUjL6eJ8lLiP6Jg5oTi57ZaS+hxnyc6d56wCeN34npth1GpFZ6YO8S8+nGTD4IBzWjYNecRsqqHO
vYzM6xMzoB/IK8zlFc7W+Zq4WgxvbXmh3IsQWuKuc9bVmrCi8ks/Wt5TIBC9ioHel2xFKBs6c2DE
Mv2D7egHfawNZrFMvjJZrK+yGpIwKPRTSGj/8XdXxfgef1xgg/CFULyiMcwmrA4cmmrGffSGFo4Y
zeFtvd3vtbnHeQ9nU4Zppmt28h9GoNvc/RVMk0son452TFspM+S3rHlA/EabLC2XvA8j+KxzQjU1
8eVEHHIfjrWljcmf6KAihxNF5mSmZmHCKdIeFbsQnDPuAUD1vBiIUKuv89NFK0CADEjbGh/rVH5D
dX74QkjAm8zf1HS/GMahp8j34Dksh4HpOF8+fuXSrg1UyYMsKrouvlUT40DitIH3fFL1SbRQxO+Y
5PfCUdA0haqFX0baysZJokfQ3eDvU6q0gP5IlQr4Q4DrS82zpBL0P2nMEEViUSYHeNapfmA/REs6
+itkPdhCV+3gqf0g3uwBAnNwChzRavUezeid2IKtKK91Ui3er+xbOhtBunOF9jQFkBUfVvlEgRps
diwD2HJeQAm/Fbq+qwKqoEeHPUTfu/hELlEOCAoOkPkAJduWNkQ/DXlU0YBmxKfvAnQQWSXZCIyI
zKib1GNXIFaCJUGbWNAEUGLszIJILHZ6pic8H7WniM4P3u/xEtBdG9HkTA589Jq4LKA/LrlNQg36
FBCQGI4BI1Ib72ppMwje0F0LrfWfaRSdvtJKkjBULxcEm5q9PZS356jkTENJqu0Op5FDrMmfo81j
3E4K+w2loUAdNORTZg/s6xRYZAYe0b0yguZBhtpZcDEQIvfuShQd2dKYCgeVSXKz2bZ1eIm5vIbV
mUJVPbQ1exUfXtN30UMYlA72z3NGRDRKryKOrciIVsc5ee9eRvw2lfM/4sg1Gt8k9HL7okxCy3/i
e17fpAVrB98cylhM7tkKeVYIqGjR2XSIc9aVx/mrMM/iXtuExTdeo+GnGnNtraWkFxQ27RA3C3BU
pGjRdyenavwF+5Cpm5SqQIh75eBet1u7QHMsQstnEY7qGd9wqyjgAMTTNw1mwHQVv5vx+NunzVlF
cgCaqpq9GUg9vYCj8mGNOG6NHjlJA1D8mBs3v49xz9oxEMujLO47kU03x9JqkeOggmLJnVup8YS2
T6/dl1p0RDogIiRYZmup5cXaTUmd3p6r1M22+6fLtDmWPjmZ45A4NZkb/FL6h6EQaKOUjj1LyqPK
0LyQo9xLpOsB0LXi9YckMP/bGdSIKr0QTgN0of/tTDsRCAGrMvoxigtAAhAtfnHRpC2iWajLXVV+
rCJz4jUCIxzwTWdKfnh7DPu1KLMvVUL5x9NKKOHFy9fBYDfBqzgclkkhr/V6Hh8mVSVlMC7R3Rp9
LhnrtICkqZihLszro7Nwa3zfSV/bgIgk7xZo3QepImc59xAODREvp8cFrjSF2KqCJZrSUlPZ5B44
EZGCDFod3AOMtZMSxAWqAyL8xeQ+YAJdQd/PsEqaFAFWkKpqIZTOv7z6uBB1Yc/JRwXKhfBCBjU+
Jt/zl+DiSPYIajB/LhJV8OvqWNN1H3wjw1q+54YaDKQF3aIzq7okJuQVXyl+6p29Sds++UIjan+n
WQI8Dr2AeeeIePqmSSpItpd+E+9zieSClDhgyca2C1kyTOEwOejiUERPqGmBzZCYbZfVPosvTm3P
HdjaR/EtKVETyigVgQOOeFJREUbphzORGUApcUEEHLayi7altcktGcrKFrDvxo0uj1XhymM5Km5P
hmTBbiVQ07C6QEAv7OKz8aTumj809yvYPIgF3aJd2u42pF3yDgij8zYMNho3Gb6VtPrOMgRiluah
B3HmHMnT62LfL4/ZiMlqwl/JRXftpy90xYEllI4wZ9sZ/krtLGKodKm4VjU6NQTouCKo1p73mtOY
JefuKkPueJe+mwp0ZbIUvu+Y6iDwCtgSqn7BZW5cCRK3LRkUi9S04FupOGKGFP3i6YaZTe4QdbIa
O8o7E9etYJSqq6hGFYQlCYRHQ3s09xcX2EYX58d+eMWAXuke1VVMKcB+B2hGKL9x3ZxDJbuPD31C
o0vVy84LEIzArOv89fGCBoHszPA6DcFrOVF07WgSQbwZSxkCCfoKju9VT/U0vA4ZZlhcXbIEudXC
gf/GbFby1AyIgwMWEkMl4gj5Nk0LDyS8rRo1HuUTFp3vJ/pWOKOmSjWX1SZbbWMWdRlyPi5TAId6
h0dWejFOgJgsP8HWtW0cUoddISgNg/k/3yIx68THxSfKJ1jjDX4v0k6YcXJMFApUHShVr32D1lm9
3I9PlpUvuGJmh5sQ2CnzbYKwzOyOpwkf9yk/enIrfSiTVb/Ib0hzuVgDsddRVbrzZ2XD8dhU9Xuy
oCH1rxtXnfJZhAMWEOes1MREd1PyYzriGIm1v6mac4hyZ+ZgmXq0Im3oiLMjwlussqx109+SS1iS
IuOgkxppU23Pp6qfUH9R8cBGR4LUMiaR8pdBHoPflXsyk4FU93BGIXTgoOXVwCSwFdS669NQLAEz
1EYciHItZ9WSsBAbW9rGR7GiehRJehEyweur2EmGNsrjJUheU/UwEUWhu9x+q4aKPOcu2c5stsLO
xykMvUZz3Xd1g5NTROJV5KoEcgoX78+b6oWkQR3O2dpjVUgy2Xy+2cAnYe5VZ0Zb+qIOcHqf52b5
n3eqYkBHclR3Zx9VbzgZ3Qg+83RHeMhviyoGJoHqzhJRFwqbvLrOALRzU5KgiutYHUNp3IW9oGgX
YptUVCpglAAEz44vbuGJiraC1xXSlLWdRI94pbB36+3GsIfhZD9cklLAKlMKg4xiMl2xqNo+1Q6q
vwCl49LgGxGt4cPmQ5+7ulrKvS1zeOsYduDb78+vkF/OL6CzI1bMejViBdO3/iLgXHc4AUpa4K+C
BlS9ep5kgYsGh0LOYnL4RlwVL/++fEEgGY/ac7OM30v5DRfhISkjdNOH74nGZETf1/1BXhXPo1xD
hAMzwW2Sp4rfkValy/PYlBfghgy5B+KD6tQEvqOd3l1S7ctVWwMwsQM37ONAHp1LnW2q23Rhov/S
ii7s3QHmLTNL9FmTOOmDbso/U24P5zNMOTlnnI8mqNKy0+rYOMNgRTnLgL5J9WfWt8wbEbH8vFgz
nGauaK2qKzI9RNXuIDfZp9EixglpCCBFGTz8ju2C5aEXhFhjLNjkYhvxr3KVmwUJv/55s+o3wpw5
ujrpwmRie2ZWDYISC046/7IHgTZKn3GYeXJRr5pUSajuH/VrtOqpfI8ieMSMunlfJhSaG/Dbmtdl
tuLmR4ei7tDzZoLhWXnlVqH87e8KcJ/T/9E3BOC9zSmRjgD6PQpZXefRrFs7arNCMs/4w82F8Iur
6dVavjnJqZAj3EyJLYYrZFOxYY56sDMN+lYKloDAgxkJgj5lCkIL/bu6vQytJu/1hM+UhwmhkFW+
LezPMK6Frxz0XRKkeUv+JuEHWALPOXyW3TPfUTgpSE2zuxj4wE70dg/EeCgjDckXuH4iqqzLAi22
C6tTGfi4j85QUurFr4MeTrg6v/lF7WverMyU1dScbe0K9Rv+ktEDysY+ALTVDwRwoysrgjdJuXuI
YbqfzIJf/T7pS9ZocQoKWXvC5cc8fktDEmbw5EUonJnbyLbD9IEV9czOjjv7Nz7kF6E3wwTJvubj
qd5KUX1F9fDnN46WHD3cEC2GIXYuvO2lHgzEmLy23oK5LEWXYyYXltZXd0uRNpAuBYkzVSsc3z1N
4z/FFhUv1JPpbImhSOCqQP/7CJ94a1HTwmSxa0A2N+vmemm0J0vpf9qeTwL1kx2piqIMgbCGVtpk
gUZ3+kHtifbZGzK2656DFctUN9kRDJLQgMZFI5VfkF2Fp3ttaKjfJbiiIX+4HUYg3vo1Quer/Z4t
+CqpoFVESXCXvIRN7PeoLK8TxojY7MAnLxomTI01s2r5bf6JQk0NGMRovcx4PyBk8ofaXpvWG7+e
KpT2+ORjTr0Qu5yxjmYA21+7QG55rVZfgPodJ7Ech/BnW57VoUTLjZ/fd3RBeTx60Viy4jDVIXHU
b9V/lbyGhVZcvTyavTyG6g4iZa8uv7F9t5lynrNcK5svq0ONEIAa21e57P8pYbvN89ebirAHtHiv
qbau6n11uhkW2uLTpSN6awv/P6ztgA8H3NMLsY9EIzpyZ7yCFAVuGnlDC9ktYQa2Hjj3iO0Oa2N7
TUVT7I9dL2BBHnbaBVpQjPxNR7gn5OuG15Siw9H/TzR2PRXNVN01TQzWmWvCj3ZHljRU+q9ZumB9
vIRZfVerMQM6uVEk7cr+4i7ogLbNYVG+zqNSYbYos7tWmXMtjE1N9EOrDAB+DkJOnD+no43S2GCN
gXT6rBd4XC1q0t4yHW9lluFDgIH9VORvaUGWYUfaTsHmQvuoky16M6Ips2Q0wGmprijkDmHuoRmI
O6ArWUESz9wIB4gBhlYXyWrFLYgEA6Ho+LfyVu/CwOmVb7LBPgFSb32nB20rucVroXHzI+tVXQN5
azabHO7fNhIj/T+4lnq+99ICpb0KJr18Tn+YSJ/J9Kr6lWbCaTpl+hqhRPCS4Z9ZEljhPTkAG8xv
+HS7om8m12jh0X7ALMtf7/WE+LdptRPnib8Qlrz6bbcO5auHlqnVQyd/1j8G
`protect end_protected

