

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
RZm5UrZFV7JOtGxR4Pzih7NQYLp7LmPE59R/6o+hZN+ZT+nCA+l5YH+/j+E+cmHHWo6IUrn/ULaG
ZkaGINks7Q==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
MRNQzUt4f7a/v9KMrin25EUCYvWi/twJzLlDdceTmDN2GCvOURSU7hHpsmsqqCb1xCeaV7xbvs0c
MXpZkAPeQc5Coi1irNf+9eKbc5uIh03B/PevhS9S+La97Aj9rjHplzcZDEBFN6fiyAdKvJgOrOyz
87nOO0u5LoaEOeyC6ao=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
L17wVQWzSUChaUkUbjAqDK1dFxRQ9orAmYas8htY5fjqeIDtBkS/PldQL1EGRGrFVbxZVbStDyiq
iWMlaMSfJiAW0codwFWqGkqnH6YMctbqpTZdQPbprA8qa73Xmy9S5tgWXo6y3vZys5HBTFHxXMXj
HSJZBGLfj5+GGMkAkDYYBZrgDs/jxx605zYzRg+wKonRxjx8C7c4r2cekqFXXjEfMC6t47HLGKZO
Wp8oqSV+SdxjNfsxTeAcFxqhiABG1hbduxwcNIQO/0mgU7awDWqjimqvnE1+KO7vQU/MVpl+J+Y9
bwvxkUUMkYnqQG/HGWvvQ7Zp0u8+rRyDh2dzOg==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
yJG5RZbV6QsAW4khC+YjJnbI2jNRxPOtee58pTXfgJVvj12BYVsRuhi1xiVJgak8Vy8V0UJ43Wc3
ydXie//gOHZIACOddgGz8WdlyWauaZ9sd1K4GlV+vX4K5HkoOyunq5QSLYwU2X/ZYYkTAGg7My6m
h1UvByaO98o6pNd+n1w=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
QjcZeibYm0SAHW7YliT2StC14hkmhpmI1+m8klXbQfAK/yXQ8NfNnDZicIHqHpAbgVQzoGSkcmXa
qhjmF7JhXI4I11rujpUqz61fAf/3PeUiYimqp9l0xnePLlrRBeItzqfetftMnQ8hBAuI+sARuLin
j4+kHDvo2V/A6kndknmKA6lyd7gI8Mgzy1xgvua2Bfq25TZ30r76kaSXXo5N6hFVjtfwPGqnYepq
02yTg3lN97x/f3REjUh0T05iK9mOISMgvqQkxFwl6hBnLhp8WW0zJBjFvAguLZDf4CMBuYBnnmGQ
axcOzl5DWDcYTgPm/DTciq3eoilijus/JUHuFA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 8000)
`protect data_block
IRiwotOBADtd2IUSMvJxz918f6L9YiNOQ/YvxTpupVijmKDnQ/ZeUIqQpQnDlMPxMZSpdExhg9i5
sm9efFVOrS7u+Tz3uDUFxMICobd+2YRjrVKhUDzKG2Ge2AG2ChvDODMIh4dZ7y6Oy018ONzTJ+8d
NSP9fiGc4qJQTO8grQXll/q8SpnrmWqfESgdPQL3kkGm396CJE1pKB5QNguI29KpDYGLVe5acdY1
7zrihsRE+4AjFwoY1HOLd/UC3Gq1+qldAJRpVOP7aSYCVTiNHOoKLezGai+2vMXVtguDe4ScisAy
Dfmn1QdwPBXN4d0hT3BjSs9/eUBpKegDPnlLA3gZynsVzunia5is+92++l5CWO1rzA3GTNy5QAkA
2lWC2CAwbQ5nOstkbamDusY3of+WvmsC2g0bm89D2PWkRZLm/ZEovJCTzCxHgl87nTkg4OXfT80p
ryhZbftBMfZ7Ps6Ko22x0ziX0cBIcqpeMQbRKwNHRAyD5a6TEV77wfaBVF3rxl3scX0kalFRIhNM
6Xh7Dchw6VJviagkxNWGdDXa8teUqY6GhEpRwnT8i5iDWX2gww8tEimpkBY2BfToHVMzMNdJeloB
4xN3C7eGBz7If/DG4ijdwLfGvyy+vdaL4qvxgUlxVETtkq/5aVvPSUDSO8WqDfllJnzb/M1uHgDU
+RPCcTyZoUtYhpSbWLx21i+ejPJCfoWTgL0AnhMjKrFPPEGnF10fWjKP1DgQFw+BoHJVvi4N4yEH
rgX9NUhZXTxsAo14qptiKRc54IYLXdfxlmWBRLsUG4liLNIWlVyUNB6YRh2mA7d7XOGyyOGXUweK
JHPpSR+wCmBkg8Ab+/2kF+UzCz+0/TtHqSh2kn8XQAI2sVcQsgWRl1IG37fRo4MM9rxNSEKga3w+
yh4Jmo4u5jTfaveowcVP1QZi5b1jbFO/M0Nxq1OVoV8mZD3s1OPS5OSvmiJVUTN1SkpNC67zMic4
OT6x7fqMdlrDCVxiXaytQBsizYMXnF7qdP7+dTnDDWu3zjjyvFAGsKpcsCNgk5vyMRvBN/XzNjav
KNLjGIEHPnUckw7wp8lYaVMUMZUL3vavYDt7bvIFMyFgzNPy7pJNpgROXkRLB3XzA9YXfCHLApLI
KkqIEhJu5kwdptVdKed1qRiHpMNYr40Et6L95g/5TXvhLjF223ExQ4LVBlyBmPwA3aPH5DStDTSg
Q+iFd7phAm78tZqsstjHF6Kv1d8h2eIg+MxfDDtwgyOPCId5w/vdR0lhlBPnL2uFq798d9rKKVT8
SmphAQyuPRfoWfcoDixmHFiIsjFUIH0rXJ4/kO9u8f7Dk4tVwl3sbkVive+HKm6XLUvuXXkN3tcM
O46roZFafkcEr0fioPa61+WJO4dsMvaTf7pM+okPKGUGOo28gIRthDLmu/B1BrRYBv9X4rRvO7S+
J9KH1I+mzYjhV9E6qg0VBCuWOE61siI+FAPYmUYp/Y0uGkuPcnScqn5SbeMlDfqTc8+x2pa2ie92
P/KCkFSD5GBXbaVDI5uE22iiLOLxd1Liz1/dVX0s879cr4hn7RM2wg7sot4zZ0sKRtjmys5T9K3m
ZYGTBoFiCcgAPM0IGZy2DYaqMYw+oUhk5dmt78ZWHeo124FYNjR51mkJNcFnf/49aNHaJ9r9OK4X
cmU4WU4jrpb77Fulx+dqWBEUnuAMDTiu8MvsACDZ9fFds0r2EX1dcKGkyDfckYQ+8I3ia5AOE/vM
vl5NEA5K+vfNlVyALzT6V1FOne/dJa+WKnj9qxVS+OFvKk60Gqg145Gt8oRzZWvL3KiJiPrm7Fuq
frTM/9YNn4UGl90S7IFUdfQTsie/zOH+IFREnDVuCMgdEeBtKPWB/LXX92/6eh3cDv06sJAPafDX
oaOWBBx+LKzHVoqN+1PODGkendMV7nCcbyHXmNkoyfFLY81LaDSA/12oXAOwfNJJWqInLi8c/tyN
FpN606yjQUmyZJOiXAuLcXF/7oCMkh5r68n3BYasqLb4udZzpdJAqxKJmnMUqluFim1zBg4qyNvI
yA6TkYfLoLX/OEOK0M9Hu+bcTi2vM1uwa15WsJ1noS0CCSOq5K1OizvieGjq6kA587hLs73UwFm3
ztHG3HaXxQOueCkJl8hfrTvRv/hzZM5THgT/gFEnDNUS/boboX3EX+p0BYHae1SRaHf9chtpUAIo
jP7Gf0Oatvsy0ptxKTr45tOIetUACD5LSaX2TMxbFFQwfQaxtBawmI/zZDUFPepi88AGjZkAkywT
HQto/IOigPYeSwcPI1nHFWJau1vjUnG1kKJ4k6eLU+IDndMLk/A7kIb/h7D2DVRmgPI2im7SXv8q
xPkeXiIK+It8pCJjfYaNXkjKbvi7xaDU1nJPHLfi8gXdWNbZspPCR0y+6/nf+em1XKL9sEV6GZzZ
im44oX6lgKYMiVDj1cYFksBX46Rt35sB+9/kyoCrGHswyQXiElofW+twQie6mwvpna+qjJfsESDv
Ye8NrrEFiHgZEXZrJHREjlFztmC34FxO/g4SesHKEfUlBA4BDplSPOjKLDzLoxoUg7SYGIUD9D2z
IklmlcHOo4bG/V09Dx4iAZV7c3yOTCguYAQxK6c/SmHAbJOJs96l6Snw1aIxDny0bd1BMK0nJpW5
yKZsLosZb1mA4o5YmKxdxE878T7d0vaGZKtvo4mM1Z/bG8HzhQHbcpnhWT2oKXrho7PfFuOZ3Mpg
FIf61Mhpj3qhA19cv3zYIEA40uljyKd4ejTcszcDmoitQsVmP4psQu6L3shgObNjB426IZfglWXB
gSD2N6P+t2gWBtM06miYiLnR1SBZWN/SSGDzSywJSkugcBgMnIKFeLp52M/44rfdGCWcjeuiDnMO
RNuvK3DjudSsR97WzTBShjrS5vfmyDw6sxJUZO76bo14FXjVNd93siMdfpKXBXY/vuQOJWLYt7hl
5US0ES6TvwKycn/kZh1gdz2AXt2fUsi9/5Ag5W2ep42bpCOdodcY5iQ2KBtHEC6imJo7hbmtoxAr
kZikEvPMj4WYxnFc9zCklbRsCF3O5iKccpT1luh9GKuURjS6Pvcw/KBg2/52F4B2dHYqE/6tVwX1
DCyjKcsduuyiDlEq5nlbV524gOik05lNeryyKDr2epmpHg3Zlbpssrncdvj0JEVz2AnZefoEk+s8
qRv0bsQY/luZqKAqyMnNcE+mq8Ppn651uZhH3xR0jkYy65SetMx4H1MUsCEnhTShp9jgF294g/DM
cWf2mILDs2uld8mx+WjMcZGPvEPqmCQc9drMWlLkMMOIghbCzyTfJISDEZnq1b2wTVYWM074MikP
sB+oC42zb3n39YP4NoKJ50xP6tJPa4IOcxum3N9Cdb+oyytwvOnONzWEIiPb0quLvF1K6ehM7vVc
vHJSk8KuEfAD/O2q9hm1pDDaxDn++yA1gOmpSqhG5pLj5AwaP6ufGyDaNLTbl6WEWwz3E50XaiVU
LQM4HWRwKz9W+8hzIOZMjoo46ZmwCx4ow8W0jGBa7Xz/BrBIOjY51O2rnsyZS3XgAyO9ojEHbu30
TT2ARouDTSn7Swhp4HgkqO3j/mIWLodUBDoWeDqgkCFenUEYjAtwDBAhPxd8wanpYo+MxCpnMhyE
3raXor4i8FX2kq7OchHPYMUOH6fKfqfLZzAnivl9tjB16HNEBwN+IbsGMT0gERaROc7iCfxMYhLc
61vYsE2G9jba1elQ3A9WTOC7LgcIbK5WdSvu9EWEa4OKkRRX0UIbTyNYYbWQ0iCRA9ZPB0QPMTVA
UwEQJqK2TIe5nu4dDMHyZrbmjACDpYBkFjM16Y6ciLiNbTMNm30UFsU4uwmkl8ox6oyzwJhxYuzi
IqWK+e82og69zDb0jRTJOHeAL7FCFwh9AACRSRL2KItgQWeRemLafZ6UsAdK+43dQyQn2xpjkRN4
itqsFViG41vsacg7xRemo+/OG1OLTOmtUtd+B2eUyCI+twJDsKUJcQ7mIhb3W5VEXCMP03VAWpPO
5XfhxFmrrIi0x/vDwlUnAoeXSZLDNythSr+lNL9HORN6w8Ji+sG41e78xnNjWvtoNKR3C8ECa9Ej
gIfoejk7OW+YX15Osh9sllX7a4Mc+93R5jbxtsxWqh000TDesULj9hSssiBU1OmOGEws3SaplDvz
s3GrixZqdS1F9B6os0C/Jb7TcWCx7EsdgohTXLYawddhQJwjS0UVl5QtUiuoRAuGusLItR0YraAN
YwoVbYbR6JFLXBLN5dtwugbmNXSsjOyM0li/piLn7DwA2izhRUzEIVtGiPjlCif+sgCiUFMtfJh0
HQejdE/UfRQR91qMVy1BpqbefjsvhCG7jq0+j1f1O1Ra7JyiRGwl6v9mhIuctaMIlV/B70fszxg8
auDlq9n/aT1id1f7v5TmsLPdHOzoAnqxfKnZyUkcBtsLrUC9fsUlNcA1J6U5V4BGCZC5IHImbtok
BN0YEpRBXR0PgL/hfuSLXf7M5UWnRDObrnkfC+0Ek5ouB0sc9WntRlK31js11+9mk1NN6LXx0pvn
sMGyIhCIqHF/IxkedEKtR8jseUTGAwo9ISqL6VG8iiWJ2OURgeLdRhljvNFdc1GV/T7h3Ho0nFv+
zBVc7hysxRiJvT5M4rJSZOwXOISylHSUyf4V4+NumR//YgKKBPzEcpgAFMG32GMX9YRe7coElVSO
z40mnkKIyL65jlUenG13Ro/V2xR7+hIxOHrB+YwJFaFP2JGfO+fqd+fr4bifz0KRMaDL91MrchH4
vlBVP/qY8cuF9qGNSe4MOJr4FeIZpSytnHURVCDMVSoGMGE4gwVLY9rv9AGgYPkY5rco9GmEFXUJ
Yg3EskGV3jpwpZgHIhxgD9pWGuH5qyBdL0bKZClErVlb8wcz3+d3nWmL4YxRSfsCHN/AC/KILK2s
Zg+hnxsW/zKtT4XbHvo/S3gSvlR0zu5Bw0pQDdx35ie4ro6wYBPeUvWDjKc4RBqUES5XPpa7sJob
N5iz5GrYALtyv+hZ/9l/YMAHf8tSzo+fPX7TCCd6kepBYbpenDzjBkKGSd+c1xN8tFs7NI5C0iE1
sggzdV2tC7UdEvXvWzB7qao+6trnL2Wzj2MF0J9YRnmNAA9+ka2ZhHypEOM5Z4i8h6Ai4HZXZSIp
8WzNUVKQvy/YzjfJ4uY5+dxMAhU+PionoCsw1otFd1y40CdRfu+fsdtRb6sTW9JylKxevIllPl5p
Uo/jsUL8CTuWOUZH4jmgCshkbs1oUn9ZQOHjyPFoOT59gDWr8Ot9U2wdORHZnbX0putGUGn4hq6I
X777vzvCAqDbnAUsM9IdgJJHvVpAS06d/foggnoASa682eC7C6R6oVeuS6byo6TULF0hqS+rnGu5
oUyivdrNUhrj6lKzkhgD79yVkcOB2ecMIRFt3pR3fygQDzh8qSufnFfPunGe+hcHfbgoO6viVg5T
srAy+09I2QaDTPfHAnlb7oGuLeOdEQZ/jhyA+JqhE9G99RKjYBfQB4RRTfjpESscRHEo1l7qIuzz
W3vxlWwMJJvAapoAlLtwUYZ1kluHyR7Lq+hD3+vwpqbIf8pnvWKNYiVbGWB7wdfzx//ZZhj1Zr3I
uEhA1UarsvXkRAsls2SD6Bz3A+74+Lyox4wnehYrDKldf65SMpn6D6DNZrx26ClfviiXy0dvOZa3
B8YoLdeLF5F6THmqUXEMJUsOr6YOHbYgCFPDH3uoBgblKhfimYl62V505f/T2f6ap5dWPv5UV6qC
Hr9UxSkCfdyuMpZWR+ZuEr2KD7l2kCaFx9Xee3RX6QgiGTDqbbPzCu+8ORqFGhqUkFHYJAFZaKNf
Or2rzCIeWQcNC8vPEGvdQGgJ9NbZCwQcBPHyTtk1+9PAOzbtAkWD67XeX+gfaP8pzwYVWBqVz41f
mvwIzevw4R5Jt6oIk8QwH52Mq+tdTDLHdepIU9ie0C/4uoFUDnblv5DPH1kDiVn+gghXXW+jGKKy
HtnhNmcafxLWsKsW1dPaSQmoOx9dwCkIusOM5HiUZCfLU7HhB7g7GmQNSx21iUfaBf+1rXb1QuYR
488gotLJdu5o4xYLE7TM/hbj3vVCKyxUxGTegZpQZ8o66jBMWhSaXgr/CziSJPrxU44fNykjMkRX
Rp2d5CCoFAUoESiEg/PcYVKIfZ96wFt5ZsSq7weXREoL6OAuooJtz7n5sAgylONcgYDSy6q5CbHZ
GY+olmT48TD9r4zQvt3I4gcHv3zWwxVZKXBDlj7+v4wjRNXoGisV6jLDAS6gxv8GHTdU0sV671jW
H/tg9V7dbCLKew3bQLpQjPR0UTaXcG+gQJqUVV0PlG6zQ0ZcZIkxdnpz9VWkZb4fOey/DrA5sD+a
0d0/d6umcmWOXlctI+0AtUPBidqffkZXt8mykS+HjRk1Ee+dipPhKXAmh8V+QsWjrOPlpRV3EZ+k
qzXcLDPY5m/BEavS4TvZXVjRuvzxMBKHGOXvv0+1oYWq3GHozumXF6qwEXEvGzikIiIUenoHEC6t
sr3O1Jq5aK2PGaIkXkkpP0+x8frUagcC/asd7W5SvXzWPYWURUGCTgSQ2DU1KoMDoFbAk6t3IlHg
SR76huTIyuUT228boaRVYKKwb9qzXsgB5hTqgscy+jKIELjv7ySiGeDep0Hyuwrb1amTUtfE8GF9
mU4VRSBquqgLDF9Jm0fCW2JSxBu7W1smoC/e2bSJen3ndrNANeQA9ECxp231OAWGCKY1PONsWf4p
i0DIccH6Annt7TwkAMnBEoNgvzdDyhzCcm1ezATWCQDizbwYMTvrwR9jUzhF3XfoTa2soUGZaS9w
WP9+GuBnsOgSsxBVc3tsnZTfUO1vXCGfdhmnAX14xISifV8qXexTv9qkhr9cJIBIKdpdvgcBjnSt
B1GqJIcAv0P6i6d/f9QTMs83bHraVutio4ljzjvHlyfO3By9QuhKfV++jPmTPwiJhMmrjv7kE2NL
8ktGYx71OitHrQnH916nI6joIGCkM9WETke7MJ4R0aqkvyI1gGJGFQlgk9uvacuEQVkeEv5Jc2oY
CgUNCQCzER4kZTnmsBaUT9DIa5+EeDYBiqDpmO2tBuQlOrM8cKsxij+UJJ1cyDyCy2Awy+Mxa6ka
11xxN8P0hEzfTxJD6kniiCUm2uWdoZ+mgd7VvF/TVMm9BEy1sHOXmRUmFwgxyuJIoX4XAU0u2QYS
qqUOry7Y2Rf5fSonorITusgUvvsTqEiWdcTeeIZpCXV7l9u2B0YUDHK7qoQLoAM+S/MQqYe2/HC0
mE0XC0lrx8WLNENCpOj2S6e/zs9x+jgCSyA99VYCQS2fOrXlPtBHzsEa36O7OyKeKtRtLNf2IOs5
Voj1gU1tL+++kpxZYt0K/9W8wE2js1oLZ7edQPzgaWmbE7sVVY3JDFrwcjl1xckHOpJ2HkowXqxQ
du3GkOwRA+adKR0SJQhaXQOObZuaMzp76LCn95YkmcyeGhtkSgfjYLUJN/gghNzuL8QbNqWM4owr
6XyeNown4iAWVQ6F1pHcgis241P66tC4I0iL+bhe3fiXxv2N1EXqDvUWyo0cf4DJRqgIEFBLxk4k
xiaR+ti9bQs/sOU4euzcKV81bougJXijCj2iaisRru9XgXSJIplJ6X2bqN+vDP2ctrPz3PIdEYdX
FoecfErzmnwSt/smpubkvkiI4f6up6NEGQZipYyk0P/b/l8UAgeFKsG2dBNnfkYl3f7f4X1Gwmew
2zOGo0f0t5V43vAvrSLbVJs2UyFmbMFhKk7OcTdsnXy9s04Uxyu6F2Co96xqKcIUOVYuO2TFTl90
yoz5k0Y12wIwg8drq0tx+lDrY/GX7rs3EjpxlBP8AYqYZDXJO3miPA/SxxGXkf2b8LFalruR8QaC
pRDGNKegjUxdF7LyStNMAI9xosPs30wJQPP6rTxURj/ExvXavzbEr6IW3VU8DHUEqSXibQVjb34y
8uoaiYENiSAjsEB+MbDe62vV+LCZeiWOiEMuuwdmW/9PZe0X9KNvPJSqU1cLqL+VQkIvMtrzP+0a
fuQrISlAx+kSgtt48tOri2K3zEEDHlpjidscYnVgg+W3bE8SEs/UyvWI0DI2CB3mYhOlHjySyO6v
9c45xgos60C0qjrBqf/odmL5r//0mjEsbdlMvVCIYQTtZaOxtbUepeW6a1L3ty7pCvXLU/6im3aU
6x//FtgOuwEyqzYBd5J5Yj2gZTk8FWVpdbaDj91W9ZyvkKYCWKjMRzjAWS6kmQHE2CNt6rjmwiY9
2UVqAeZdNt1imG+f5gjYfQjvQq3EH+DdaeoeEM/fJFBGZIXkZ6arm8FOsMQu3s3fTxJAZWEHyi02
UPWCpv95UxU22hwAY5sWEzqDkdLfTFfuAcvvezCLCsrLDlkmfL8+GEZaKGG5kLyHSPXUqOu4eKSr
UzFYCtCtTnqJP6UofChGFEFxMp+8UoRVgN8I9b96Dw+1c7h3oIpo2maimstRyugeMETO4xKX99rY
MtRH3pAI9sdC/GNKvlJeOi8sq4XVUJw5bQ1SWUk0w/BzNQKIOFk7DuWzxJvmZcnNZusSnbgD1cxB
LpJwW7tbUL/DpW+pUnaS5faI80bLYoAxJSVz+jFf2MO3RgdU2TzR/4B5HZ3l3+p6uM5mF5VKsV/O
ys8NVk/XcpyuMg+THLZCdqDKQfPyXBkhXKjyKV8diqV89x8W92fjfl3XMxmCLbMFy5qujYQnYuFq
T3sPV6ouOaq1V84wvrsAwsN3OBunyRtYcsWSLPoSR0cbywfRKyOCzNMHhtd5S/XPVj/J+4eotsgj
GxbePty0Uz4Se+DVgeDI2LduIU7sNPbmY7q1fuLoCo2fSbfNrSz/ILG6wYfgcAS/QvMBc1Zi1aZf
4y7YYuOUGLD4e/Vja80OPz1cEAbUrczPKk9bnPxSrwzruxz8G7LrB3eZsHyO/BPj7nmamn+mFoLi
fMGeomYzOy7OkMRGrXbmdCmMhk0RQaU0QGyQ3MO8A/X3Na5YriLVV7G8RD4RzhTBcsNvv6IyHZcZ
sk3TpMx3O/X/ty80be6bTjBYuOnpB7ET8VhTBMAuh2vjL0m5oXzsAG80i8nHPWZaFR4y63+Owrtv
GEEXsGzKNxwklzshnJJcIKf3ICqt4cgXnljR4hYhxhZQzNBFvZpy6p6nPGlfsCOv5zP8B9bxGB9Z
pDBn3L2b0IZBvXF2tH4KwpGpLqzPqM6/df+506bTyVCYmuu54o0XdkwuVufwbmYrCyw2Wi3h+xhp
VdG+GPnKpu+B76bAR5Z3Bwg06+vo696UnJ/vSUGbSoJbienD8hvAhvoZEthTeuD5HiYico/8ss8/
kLZLksEfYIKOs/du2yxRrc5uTzU1RuqBSf5zqJZviVlvvkzmPbKZo9WESrsKVNZwp5JVPOb5ZKjW
ZZ0uy35CoZnvLahZNoy7r5p7H7YqOXlD6xfCavbb7EqvacpXFk7KnVJZlQfnmt0nqD/LAdf/5IVG
XYoVUwWePbFo7cK5WlPIlO1IUEq2IvyxlHH3i0ZIXKiDO+nBqN2alfbrFkXPnyg4h/vR/1/JfX6F
4glHfyaXAz0AqG1xNuY5220Jf+utjw2V2Uc8fagQHWC1mwqWkgHEVwguJF6zh2JepPHK5bRtCPFs
kswXnV8fk7E4VYN7hplqBnj7QZnz8yuBeiFKTA2hc3ivFcwQfz06cVXmiFl1bn5DfmuDWUFdgcyo
euxp3VZcG8YImhBm/t6w20RIp8+x0QH+LL9TbALIjFVD9FeLZKLaZjW2VL2kliR76HzzAIE9sxuw
+oVkYQktJQf1voM5q0ccmfepnKwQPwB6NBULxMLw6BU5oHYaj5J6/hJonPE1yjN6LrH3fLS9V24S
vpetgDf4sH4yrP+E/muo31UkE3lEZEZMk85V03wiRcvABZiry9Em8h0N6WCljl1OWF8IKHwaswCh
eIzFQZggdkxYsU+xLRWFMBOoPhqU9vgtw0PuJJhK08wZoSmiVjm3ajIV5FN9u+NlcgMSsHqdQ5CX
Xq+jkokHKGoc91uQUUOrkKmRNCls6zOjDcXyEgEeiLAbtTMu8Zx3BVeRpw/Zk2VvzbJ7Wfdap+Iz
YhDTzAEOjcYccuCYuoi1KY+ZXNgi8u3ckO4/10Mse//HYcTTC3kDdyAiN9mPsmHNcNuXtMSMBAb8
E+kJmvB6DDNrNpXdPZ7zyNjNN3nO9WqEBCmUHtWkjRYaJrFWXC48BlsF0ShinAA8x1/orVrMrb0s
srODhNFIJ3e1d+z95dsEnwjpvE7ZUim4hGpiLGaPN7fl0gpYgj3gKU+lWbzUj6HXv9N/YNcb05CH
XWugGAwwAoZYVVMjt2Henou2FYR/PRAUbyIDVxJvrFtwj4FY6tXBR9nzGEEePOCdVBNOkmozEpc9
JkGU1Op+EUwkGdW4WT/jpxDy0gE3eNQgwJpXkzeUM/Fb8igH2aJmHGI9uhCNf3AVQIMo5XFuIGuY
s1v5LzSDJuSDq5/naDj4+ICQ4/wINsvWQeTaoJMsfcu3KQHzbC5/kGa/6LHx7ZINa8k3wO7zefh8
uVCES209hv16xWhtvInx/Ib2AwYnytJqqReHK94JtGXJYD0gIsy9AiCsfRLcczsXNhEwcw44RoYs
qpT1+ySvmlMqX7JEiVc4yD72UuY=
`protect end_protected

