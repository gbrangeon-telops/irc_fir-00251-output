

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
DZrqnYwqMkKoBvgXgaWSB1Gvc9B94Zr8xHWYvXS3Yo2in98iiVsrSf1RUePWKa7hVSyhM66u+GP8
6zam55ovJA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
paoR3khjnzY7oR+WJ9YkW1A7ZzfFLvvVEXiP81AieLlGnfQuqZTzy9TqIBQ7d7KWJF2u8/GBJ9gB
S/XHVoSTyo6Jte9XVVsqnnFiHxvEAnWbM2e9+Vyqd/Q/lFB3TCGyLNKIFNdGxyml1xea2Gq/DUf6
P6PVaPylNEwivSbuc64=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
IuseMdZSknnKUME+O/YmMG9MKbslcWjYg4y9t234jonRTsM/8uUOZLlJPdAz0Ojsb7gi8Afg71RU
Er0Jr7fpQJ8YMMDdLQ9qwRqf4zAR9ZhntG7zWMIroK9jxtC2bvBKKArJREVpkzOWU1g2+f7dJ4FH
ubSzqp/ur3VRiEL9rSTe80jSph04B3Z7vLg49YvLUGmYKlwP09xV4/46qike4zQtuofkQ8/u3jTv
rlLcM6RtgeLWfD/CY/EWIIuhTxeQiucCqPyYilV1cA55FNKfdMv57PsY4PVV/CwLFMYY9INUTcQ5
vlvEZIaCBXiBH5TWThAkm9erewSr/bL5DW9PTw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
cyY5ZPlO3Eo0cmsRtMR6yuz2Eu2e6S2W/D+8CcC8VsHPfbx1fHUAOMrMRz8rOeXuKPOa7h1hSFcJ
XZ1TcAU5VIvCkM11jW1o53hK8qachmkkZZnfj8JtjstmyVTyWri5LmUnPYRufwJmQUQ0xqMJytkR
VTqDp0ZVnyDWp2/qKN0=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
WAcKeockg4TPNpKWNqCVvf1P8zBdM0HIqALOQnRkxsC2RA2Dy+P+XMiOG7cG04xrgm5iFejfnqcO
5lDRzw1y2vm9IxrTgVR8u92CBfbBU5si2daX0ciu3+tUaMvbyjjRBHmWEJd/+ZgwpEBd4jKx2KQp
YmRUDFYL5WDDgF6aGgbY7bniF7p7fSFQgxz06UbHJt/aNGcXnfge+DPA60LgmbiAZYAbqv+bSmqg
gA91XQkI7oyEKtZ35D6ZzgJ25i0EzUAy/u4ctGTC1xnExC071TQUx8Fakynqcki4h3cwrvs6RbsQ
1XULS0sNZpYYdAavNOXALBW23U6uD7bNRcfAog==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 33936)
`protect data_block
ihltFYeDESgZQ7H1EiPyBddpibKvXOatJKzO4s9ulPJEFznX3OX0Ew8VZCWvWV62apuLpTq05Wqw
QHXbprzY2uC0YgeT1s7cARjTe0O7SahT5P2iRkEXeixg8V8o0sdh/kt1f1aTFADgHPUd+QHTxZbg
k1NTYW6Ol7ribnVOI3EkG9NTYjcCFLowrMcqindPxkRmN4GDjERqBfsP+uBXBRTHK0xnFBBwVaDB
2W4V4QQLX+/o+Ys34tOv9Jb2HVjGGVWALJtrTf3bp0vw+N10afTrHaywBC8670fYAfrqkVF6Y3xl
oPAv1tr6VbtqIF3LI9UF/rj+ucGiRmHHMbO5hirbln44p8TBva0gS6IImCAMOc+Zsc564KYL3wwR
omM1zwm72tni0ynMmd0kQDq5Eifl0uDd8kxVHRghdWsDtaNcUX5jhO2/OHwZ8vR3Q48ySWOKsW4O
t/uapp0QKE5tMWbyHdVvDSGNdWJcyOw1eEiMlZlujgok6dfZP0K29bZ18//xMttK9PMenVd/7VU9
bwMLI+sfbdLfDJyMyOMMpbvVGNkrX7h0fb01Fonmx1/uIQT2r5IueyKoY1SfZbU7vvOWiZ1yWFkC
8akFzcxeXJoHmQ9LENf55XlQxl/daCNFfGseiNzWmhGLTNow3kg1eYm12X3X5S4PUX7lAhgkKSLU
yQiiQW7YCvkEQVfgYG4YQAwkKc8giaxonLVIzB3bK43xbCahmdoJA7wTXeYIf8PZq8lvF1pwdeLk
2rXY5R4aNcNZRdffEQTfR3UmWJxr3LycOZD8c4qTsV7W6m4LqXTrpREkk1gXfhbJnMMVNfjh2blg
ae3aleGmmpxlLXSBeQrkY8Uz1wCvH9g/OLjGLxuulsZCdcQX89UF7+Kg7rWHAuaDLjROGTZgeqjp
w7BS/xWUNUwCTUNLpJcDVuULFnImfvpnEhlIv3ZWt+EQMFjuGGULElnOuwhe1iU6czNgwXAmumui
OQFcLbrWISFIbfEzANsOnJtyU3t/+NZp2N/7A7+B0WQ352/j7S+1axQVSFkN/yqgKRQ+9YsseAGk
nbGBmw7ZKtmOvHzds/Mo38xlCIgfoTmvc85iLE/ftNZslj1qe9Q0A+2rl4RMChtX5sZE3CgvB02r
G4BAUfqFrzZsM046yJhDmFaoW9xikiCHnxcWA7rZMHaN52KPa8H8OYlAH/RfY0lEM9Bbd/mkTC+j
EHMX0cE84O2XxMF3XOzbi+DEvceLkrn+P+TIWtOjqsyNNWjnPkrd5s1csFSe/+ijcSs7BwmJleez
piK4IwXwXXoGWjQ2pGgukrIdeiSJQP8KsiRBzXZYEtywtUKHrdPSZU1zknZ3MJ0L7gFGsi+mf22Y
wy9/oz+9VV28HY/1B5nZYQLV9zvuJw4oBatyZW9QVpkG7Tae7YGKUUbP1WzATeMekkgJp9uBER9I
E13JzPP4RYUbmSQ4GQjMWIc7Mg390y5qXco53nwQYeB1G4fytA7hKRSgno8AfBf0Y2HTL0LFbCUD
KvZpxZFFaOEkK1BtIY5OcWJxH05K+HVRwHbTER8H0Esj09SjrUGS/XR/cvJ2QfBGP9JoaT1cSatc
0xZGLPVHXnBK51ILt78QBl1ankr+tW+poEwQlT/ATzV3RvB/cXOe+Mlh1OYHcOFmQhu6RDs+d0W6
0q8g0ONtndRLHHJYhx+arOueR7mIi+abWtKNP9E+RFkw5kPsLuyhf38UrdQgBKA7/VFMbYOZ7nTe
R2LttClAuQ0Seh7UuYcjKrNyPtEeoaZkBD5CxTY5FISZr5kqYObaquuZlDmQ44BjhvT4pBHMgQn4
iGgptO6EO8SsSNcBObHQ+CBPsj5kJwZiGxxXClVdf3F1L/3PAA0NNpwYAcvHV9uh2Ww8tYE07hp1
c90T6zM/ne7/4VESFqxKtjfN0GLSLf5jPMN73d2C9n8IMC9z/sEAY5hS4AIVw+nxlZX/tBVnhrMX
Fy6xWVrVRAB2b2KWWRp+OFsP0FKx+woTZNwcOwmsJdVrs94RoTK5/AUXB+objVXHqXQ/1d+2FS4B
KnNv8gtSlNRmfQe62jN0jzSUTx+3T7R1/RARhhV/1YZtw9Wkdh/MswoJsfjmUc62dsdBcnjE2Czc
c6K6wZnXQy2Z1MWsczGcx5X7Pi9qvaNN9GPrqa1IrQDxp1/iZJsf4njV/6W1vPnuOuNKR+LvBsHJ
dj/WtriseHyG3c1/fC4akTnrPpXSxG/XHBwE//HEhjqRpr+1nhs1Ke5OmP8NUn7uUul0Od32bL+l
Y18R6bHZ6VM6T6pyYqGOhbqP2yZxJtVCVA70ccBTMTqo7lLHxFXy+m1dWxnBVErKz1T/5IcpvHoC
tJBdJYm2bB/C20LrKtUFd1SZSUu/0BJ8wL0VRLkKGcHxoVS9fEC7LUoyUoD3miDnzEREZ0gEgHzZ
hNKukYZ/eIsyWRYIq86KQZviYMUrVL8yFkc6Se9Ps1NLVxj1jG71I+ov0LYPkVTL8OQqBAqDrC0r
G5WScSJLPBBA+/fIXQox7B9Syp9ITVuIr7Vj2SV2aSHwcSfTGZb/tR++eGcLpxYipMuuRwpuQ5rx
rtnZiSnxX0G4Z1ldG96V+zzCdJpB7LZAqdG+hHwYZ/BT7TUsYT0Fc65mirthnHcI2OuBKeXm9cPA
6GZFi+LIWpa3NqscNn+q2Rf5zEEKfVL0DKffhklnd2LxqJC/NBpUUWCDmQOPyT8s40j8vqTnKWUx
ffXaod+i6i1JiXYhPw5DrexUX56zGVmJSi5mYgxK4o0fJ6mJyvCnkS7iRpa7dAZnW6JD7Afzt5rq
u6Y0pJrVomC1UgAb1y46ImN0e3ZpZLG/88nzbvmgM2vJtpT8pdRmi57IEuc3/ffWXSXH/5sCYXP3
DrvRt5OrF5Kz/tgMsDCQqqcjSptmf8DdBBqedSoTkKxZR3abxN2Bw6gnVGZca09V62RV3zrRH/BG
jgBhxfenEd/PaIQtZOlzkkd46QZ6CudLQO76cLXRx2rnA9VXtXaStnjGxNtujNbtUeo2DBP0yJHb
VdluBry7xHBwfRfC1nJmK/ev3iNwJyqU9GzR4CNRNXbTyEXz/MEGxJov+AQZfYL3lfLKykTwLHqz
HBxM/ZKiTwjQTo1d5ben0DOVa2E8jjuf2H6I/tONmQ74ZCoaM7Y6EzRytE8e7cipV8HD36tb2Z8f
3ZNzfN9f90H7lJ4Dy3GOS9rjD4LK7niDeSmKZsrQAchgiP+3SsiJfratMfHh/tYGuA4W8mo/ePt/
wOOvDZzzkzDcYLqvijhMR8IulAS0K0y/edqFf3UFIUnOM008akHY5EG5shhHVLiXdcca1Cfr2/vJ
vKIaYPjdWohyWxOdXGkI2SvUvN7joJjZqrQMZu3iHAGUlbFVz8+8nzsTHbk8Qk+x4E64RVPRX2Xm
8lvL5tuwQtIFYi1hW42x9ALX7HttKNmKWa3nGhiCMnrBmW2xtxG6l1AdASjKPpnQMxSThmK7FsGe
fLa1aba+PhcOOCd9JktVv3Wgq8w+eWWgJMhnneJXLUPwb7qpoDLdrR1oSWngJGrZsQfL8kzWnhbi
oNA1XWSvghtT+JyDe8ENK6L8rCjIRQdfzw+gD9tx7715r+u49DCTK0mKNvImCA+QQdnDKD0zS3/L
d4xkpzbNPx6Y1HtHZuw1NbuZDm8Xw9FvWOowiHgT4+oV1SuE/EtqWioGMUyxD/3rA9S/Wdo0hZ3u
T1Bh5f5cGJo6nxmSdTk/kb3KrPv+2tBDaHck6HYlMojoI50fEwSCFE1oxG4NbRUx9g/XwkBKsa5s
wrwwQRBQ6X0sFzPEZyzX3si551Z9TKe+KEoiui8gMmzEk84buWzBmHVWM11QR8qCF3s2XJa454eY
9sc1yJzgiqAEHXGFXk7yyoD9PpxCCGr/PxIK7XY7Em6HHHNXuhDZGNwRjYOE0KaKUTWGoIctHgDl
8istd3kWx8M3QCfBnJ3kR8IFdEzoJuotIJp53Ok+y5YGFz0IoirvnWt0xTHwF/4Ww+o8SV2aytiA
SMFHbUzPk4YRoLDcPRSikJ05e+5nrhk2ZzLJo9TDbvb5JsVoQmMq2ZiCO/PgENJz8WzBTgFaRhHq
W5d3PHxWEJzmpZW3Fo1ee/IMkBXZGUicbuwftZfH+Sk2gsn8iMGnZqZ3BNKtax1v8No2/lj7tRIp
DWkBbnukrFcu2uO9ShXQ29uK248N43L5NKcSYqLqxF7rrV00niqNRlqA7znPIA8u0PhMb6VkYzCP
95aZmyFDB3ClQ0fmv2F9Vi2MjL9iXbAR8jQ1qD7klWZWAPdCam8jxP89KAXZvZ28fkmWeNFJ3iN4
i1EwH8D96iwy7w/cVP6KmA169gISytJN/a/I+F5l9c09ZLwc5TlkyP5TfQk9+w9WbT1nX/c0ml3Z
g4jn/PLh91rsErctpv3xaKReQDECxMHO5hyHrELkznSpZvBzqQrFLb8gloJPLR4ZMaUJiPKB/WkZ
GvUsAAy1n443lIYAgP8DdJEIOFoj5IghSTGqukDVXOFZNpdT8f689dbgDAn7upTxr33Ls+Xohy8D
nSjV4NDPFu8bklNAmAtCYnPIu9S+kVMi4HFFCyrtEupBQxIYeI4M4Cs6R+5eaalE46l7gyr9GOXD
tvVNm8Jg3ON8xnpKS+2ChjaiDimN/z1ZvQjnHdJIKwcL19uW5D1NjMI1y6Ncp0YBqMt5wqfJ6YZb
F8fXOKTz3CUXaMs2m4w8mmr8g5D3Fh6a1SpySQQ1qSehwRLUhvvm4Fv3pib53tygC6dvzhsqaCMC
9JOZ78Mk+eKr/OBcJU+aSLATp5ejTqoHnBuz1qxe5iUxXKqDDESBiifWWAyBDRbzO0ehBYq5JMBQ
4khw+xpiKvlfqmm9r7aox24crBD8gXeISElqrsbuUoKq/I1Mycr+9u8IDJwhSkKujNI+CW0OK/Jf
DA4Y8vgcr7n1S7q0RZP2dcCVBz8diq7LqRPFuJ6FfPmYj378PXLPrTOkbfo4/Id3nlCOqNTlAY6U
dn3Z49ui9z+hKqbPZgqGf0pLf3UOQoLeYNvqeKbZo5IyEw087nsfocUNXjyBUXgaN6DMkWdVbZ4I
0CMvw6pJyueDhFzV5NtToJVUXQeowtY+/4MBF3J/P+mbqQcRhJiuXH3jlUwrAGGQdAAy5A0CBS2J
t8yXwweI8Jf3xVtjW8MDy3Lp56Cg/Wk8FzFhznJ906Cptwq+smbNimP2Vug/9LH0CngEZvRL9xUx
Wy8b+GtNRguDCQcS1FLthsgKqA9lf3s6AImBKKA6ZsEzxhIXBUzUu5z92GTIFYdTdhTCz2LGVf1u
CEXLgcwbN0DWeStteoWt13KD0yEWFVoXi1Q9D4EsWYy2OLccn1+lAEtD86GxtXMGpHndVzvNF7vw
1JuZPcPu179GwdnCYni4X0dosbZOhf6fKeaKMVVLF4jSwes7WpcKoar2ERJXZ0DE2ICTdme55TKN
toCCDnXj9uITbWL1wwzq8qvHb8O+QcoUzbSgYpT+5ez9I5YJYjMrg54PsNwlrWWFIr7dNkclbGG+
KTdj4g6vwkq6WdvU/vyEhUQA7s+NxJDpDx7SgqXCWAnSYvVp4FhJ9dwznsWNzvXOX8/Fldvf+3i5
4z0d5KAzwPbi8sr3g0Gwqik8rQj4qYwd9Dm7Ezw4ug6dx3AqHxNGPkwYQ598MATdzeIwkULhTPoQ
6OROl3dx9YKL3Ox4C6TjXwTpDy9xc9C7r2NGZCitYqVdM8HiYPDTPJ+a9zFo+Rw0JMXi5ridVOqs
PZxQ/HjPln2lqV0DDqSFG0aQvn7qhvzYt1aeXr7Jy/uzr4ZQGv1uZN2chFfhewN3q87gDt4nAz5n
dNXpUsHhnWqGnTbEQlCnuop+DAuy+OjSxhct1p3aLgETXg61gSmOzP+Cp7KmR3tG1lNTGBfn91kC
rgepXpIaQcv+ks6/a86Lb1XSykNkutwb7qX3/4ffdcmvrheghN2Ik+A2i4U93vPAqno8Me7FASVr
8vrW3v+nZD7FExAJR3rJRfUeEc8RwYarX3vS4aOufNbVpkrW9VdvRMBv6Va4zrajpB24+jB0n+c2
8swKxTcgo5IyY8tcwlmldga1/cEKd+OisqwDkdOHG4+5a9MYxqHXu+LpE9NWgw9o9vNgzowI27ci
i5H8ERyC+1PrkOfghQkarO6iHihdu7gzLzaiW1o6JSKzYpRIQ31m1vZwlgJagahbSR4i60nFAQYZ
EdmdsFxjxZ9VCbyTXWM7fS1tsZ5rcgA/doUxLaBor1GzcHigJdQjOWrV93K82EMfZK1TGOQIDEWx
CeIYEEbPG9hJiEqA5wtj97961W3OlwuATjhJo0wjJfDJZ6SRrNECfGtqpAliGGOBSVUz5xJ84m98
KRxQsTlCA7kUfBYS1uNcrEm6Zmc9MdPu1L/l98zmrQbiLk8nNI91ZE5zYEtst7Wm+3g4IlBrICp5
cfyXNU/CdC9oGuSCBklVvdFX8BHmeO/f5od0kwnF6H5MsMe6lCoWhUBiVjaL3THUwprG+oE9maVG
CEcw7zgojwEWtUZV48cbXsFb2gudBVCHOaXR+JVliCnuOCW57rz+kXIff++tf5s84oio00x3Sx3j
rj6LlBWesSrukrmLL5e8KlHbhNxxD63J4rK7WjniMvSoGfzyeaiweosK3OCCw7JVw4I5QBc+tFR+
ewN+tXc7uqv6mx2bbWfVeK/rRszOfFFKDTViAM5OAd3OTqa+U8C9AZdpf5O1xKuNxPJrdezkNczo
uWFrLWS1t72k22+iuAIvQZJ0qKwaZ1dWDWmLYfEoVyztkCUBsG1bEW0qllw3br99zIt+55UDGhCb
zAvPgT38EhnN2N35O2m0f2bKln94MAXrWBCauS8QYvKGyhvcpmlrd1wxSXAnjNGaT92CHZycE4wO
IyzClzhytkus+/XJz3Dw4Yp3ChZJnvNsYotTZCfUO4a8kU88waEwlh0DHyUX6vlEWYMZgqL5G+s7
Xv6QkeFxceEPyp8xsWAuODPlWw9DkmpnHV9dHej8USv/L4VN5xchZ3DxiDHohZFgDjJqJP0wXDsO
L+wMgFgnvW23lntAJi7VbBPL3jQG5oncxSqIUCL0IGf5RLDZcZKWUZSVk/l6Vw4pwfQy6/0WUlKg
7igU1jIQHbZ6NKve8iFqL9cFY4GmSfFtBXk+Fzx75vhx4dBRc+bRhvis3s0M79oWn2Q4ZMAupoGA
x3Cs5iLGbAKVKsbUwR+kMvZvlaT/DEhxORWH6GVPftXykioQutRHAu4wkg6bZn8p+d9qYCiFjWRA
VGLpqd8JEwzuaeL2LEHNlVn6YZ8u9GAkbpUSw6fS2vcsJ4dzIDbR2mUkh7ornTVyrwGTSzwrgfzG
3KYhW/GXjPT4Bjr/h441MCKek3sOClBXjtPQoZE5nIa+EL5dVjwdrOnFoKCM8zV6D9YB7+ZNmxu6
9JdjIijaovlMrb9sdZcSZKyxvioHyGWzVEY64ELSdlNP8uoCED1KDAigp+X8aJqQJQthFeUuGlEu
RobPu4LtYw2XmQLKvrh8weIFrN/SDkc6cH25EmgVXGLqBGVBXi3232zVmyyI2cSJ3HsCAFWqLcxI
oGVveMLlKS6K7dqY++pRqU4Ioj/zsbLozJ7+2bPkNYUrr6sRzbwCZ2T2IJpZEBxpv1A28F6UMkKD
y/BzatxV5sWgQpV90o0vcTvwjRCRGQic1EFFPmRu85FSAOjCW61gfaCySbBlP1uSpK2f8WN27beb
mcXuefr6vOE390Myuv3gilUaunYgVVelie25FP+7xdplAwlZXGPETEOp0ZfYI9Ljj9xbECYKbvuR
qpTuzaxfDjE5VLpRvkpipVppyYbjCYwtIvm40JgmeGlY3gRDuSjrT2YbzREZSsnDMelm3Fh++hAK
q4uxPap3EE7ymiuMdgzCkdev8y0YwYj/CUoB/4seGp2LtiS63BaWP0GOydBXcoKwjrK2ttjwAEPe
nISVsffr1GUSjZz+H/9VE+tFcUmR9JkQsUIHFlgZ1zSQqwPzqUL8AuyFjvyPtFX5x2pgXR3/Vodr
n2vI328S8Jms9jM6qb4w2YLuTzy+fuALjKkkOUzYs+wauzk0JcyaNP8D1uTjvnJGArwrvUqWE3NC
euvjIPSTZ292mtcQVQMpLRW75X63yOcruAUG55xc8u7p/Nw2bh9pWKTkLTS/I6Tzx0Nb9lftzIMK
1nQt5uSfVBrCmRkfvZpQrG6NoW7eLd4W4TFUVm7rY7pkBGxzH/v0Rmd8r9YA2mhQjNxenqRZJ0e2
yoLPmd0l2UoIZLehKxcTuejYvqz4mSVEWj0qC4CgqKtVE5GesVqi5sA34WLxHYf8VAj+NWCGwP94
D6N7EQS9XnW32XQurnOLCGcN2h5BgTNzpOtD30Ki1e1iFM3BlmygG79yCn/xZSywI7sB7EExBAoA
GEAOQzTXHMaFTArAYlsS5hpZR0AoBo1oRDlzTcrNTeXU54ckstADENDtdamd2oBSz3hJw9y4Sped
lMk3ps6BVw6nil+8efD0s1JrbVIqZNVtQ+ZiOFgX+k2t4DivytzzDhdJhwLFHEKw7hM198TTEFCD
jtY+P6mWIruYlKPCAX4OfpzY4odyX/vlnthH5m+WrRssHL3Xngyoi33LZUxmhqtrW/xFIVYzIbCm
064hdbTfWlbsdg7q4oEZpInFz/AH26ZXssRDYTDOzvU+wSFd7jkLputhUHKGCITCBDurvyTHvRRU
TJqGib6uQQKLzVpeay/LzwtzYfQIwZ0QP3OQhrm02pENuCzjr8vgrf/yPgL4qH9IrD3yus8j9/ER
/tMcQYnTdtLXxJRvuZ0hNytn/LM4HAduEplqjjlH6oR6wYkq4Dwxjl0B54g5oj4b1qtWPVW0aLWK
twJqlHqCv49GYq79xFiMrv4+djvbWvQoR+Pif6DgqWMkK2AlP2cn/yTH+ALrnRomNIu7g3eaU7mu
F6zHFNdUHoxAfjUI6yB2SbiPOcRWHmk8cRQKRPlba1uP/smuUE70whPOTQC0vYC/MZz0aP3Amd80
S3oGyk59rZFoBqN1jMYp4uvfL3uHBlcqOPe9/l9DkocWOG9CcGR1G3icGFg19tW9aOj7D9O8t98W
hAppVAEV4j5+W77vrLEd9DZsPjMhgKt8zarUMas1BGfDKL7bTpz7HvvgxI+WSweTLCk7DYTyB9+4
buw+Mhz1GXJmPg+8n59TX8tG/51pyi6Tf5iFPX2UusCrkrCWf5rtWLP7SCGVoaDPcVpr2xu53qiK
mPa3O0A51S6p+JU0oF81O8xj3gnU5N+58o1Xdv9ZEvzN0owlW11Pl6a6kgTFGblaJwtSX9+68sbh
MwB24ymYC8jhgeF9s6HjJDVJ9G0faGZyyYpR+tdpkKDQRFHryzjC0mD/Ngxr6w8ZIT+WfXtFg64/
2vkjULaSsC9T9LVEMuOPGb0o4KZriONCvxMH4WPaO7opuXB5UKGf7NA17FWwUyL5m+wJq7J1zhu4
5oUCm8Ap1iJUVKHRG0HRetXTWTJstLrfww6W/1sRpiM1Arqb13WQqPdAsjF2FZ561oxC2TKn/phA
kTlskPbYH0r4ze91pY8tvUmFsJnpKd3cC9rSmKsRGN9vwxSiozQKtQNWDzUXqqAtZbt9aJPo6cr+
+x9DlZnN4pbMxWqyJTmJmDeWf/N51TiuhJQtVLMyTR9T27qZVQntdDXRWlF2ENcWNYB+iOPSV3hw
wpopSv3xqzpreszwhLyBTlHidgKJaKzsHaiVNvyvyJ9ZSC5MQwWG6ioSdZRmwSbu5c3jwSARYNq4
pGhG10NGpY7skQLpNe1750lWczTDPSPx4Njs6aEGPQeAgDnaCl8KVG1dwY95uB78a5M3jPAEYbAo
EplKOD4RwiX9wKfk1kDMDb9jBJhd0N7Zup2minJWwCnSB2BZ8qWVkOqowRhm0BtDSeYoQETwjhpq
TMHiTu57D5ajWrT17JHGO5HeU//I+cjYO6VyYeckVSys+rowlV507r8Os3qHGY5+WH8smwnitEyQ
BhYyYEL04vkjzrqhsNCTh0LNVhhpFv2icKYJeDF0LdoxBZaYtanjXctTzB4Ui8OEXdXFLlVBm2GD
VWIJLDNMHKchJvbjRdgdN0yuL1nzRHjL0SQH8Bzb74M4MgR5zv62tzqd3OzdXlDK356Drt7gmXwc
bq6hmmk36qfy/u0cGvo9+aZrZE75umAngf3+Q7r+iTuV9HNCySaYX7hkfji5COwnkfhL6k0K4NQr
iZk7RNJ1jKT+f/OoXx/jrb1s1Jl/hwKL2WoWhZumZXEBNjFbrgjQIqyDUI+rZgxIE18OvKGwJw1K
vrdGR/34VLbIyNcuNLymPZ8UnK00gAQ8VuqB6vqhxTyt2W/sn7RN6Bk6pmdYDdcpIbkNsqoGj3ex
NSTfr0FeZ72oun4OPDnEZeDrGLLqfIZoQ6LYHuE2FVrk6plwmccOZvrnwyrPJMLw0fA6yvRg4C7I
kW3SiiOSLGUzdNCmecRAdH+7OQaGAfi4+XD9onjKw12+2Kk1X1vCHvlqyTtZ+nYFpZ6QPnwdfbkg
KHClrMi/O9uXI8flP8PJLCZSwVCYTKQaKeRgirpAduyzYCJbDAeyJMlAFaDhCeL1R7fXQ/ClyFiy
PUjDS3fSDuqD5uFOtUMBalk9akNq6Kgfg+BNP1vGdGb/Z7wksuapy+/CC97jAe+EQrsvNESBBhTf
GeB37ce41vZZF446LTY9IrrFZLl6U5StYwd8GmH2fJxw0bvM5gzH4TOxQEQwGXpn3ydNEHm7j5ni
7cGljEERsQ/OUH3IcRa0bZBYegPeLut1pSr9QnWy7lSZJQHHULJVfxDYRCFhCTaXri3MtU1+12Qp
0mZXtLajDn4v3CJZcSw0EAaXDjcV4ZqseIVgpEZ8kI9r+oZK20Nemyi5YKKo1bM+SeGnSDCFDvbS
ATtPLhZej81la6BT6djilKhr6f8PxEoLU3vBI9UvW7nuYDoF/hR06IKDXaK+7qw7wjXLOTld+P3I
98R/vj9rouALSjFmDSC4C49mmyR0Bofmfivmz1PUVUoJN7tvGVCOyKBTjMJ9fetxfzOPM4McTi+C
6ft5boADYWqziAAp1GOwtfKAdOtiGX38kroQ9KkjPyjfhIwBDZtkG86Ei8MVJSNrlUhxe1dygzSV
PB+za/qMuSvvkXpt6oEA1R+CdPg6SdJmM6B/NacMXVW1sQfOHdNB3jV/uGZg+w7Y27uAwnrQzbGT
ptAM3NfCxvh1yB9mD59cTgRdbF7J6Tx5Te7UkwVqW45JSmzR75ohXMGeufMquAYIW2XGv5iCm5bh
ALSQjBMJa0zONEX3cyDXTnBMtWqb+LKJ4pND1DTLYs8QaMpkrDVbesgr7zBLPm88K9k0N+iubGpu
OtGBqyEytFDenm5VIEx03BwAYhU6wqWZwYpT6uEBYywu8Cb5oeerYY+DP/sLE4MfGpNpkD7wYfZ0
5ve+xM0LwcdyzpuyKQKu3dHpzI/+JgtqirT68+ExGJYhHjZRXzXld761JgHVsKptxg0kqVVtn/b4
SUp8u6PjCHw1CM2j96040+k8at46Q0weGOE+JF7ibXQW1R5P0q5QwtpwFe/4qbcH3LeT4z/tEDEP
evUi3TIVK85v1+9WQNR161gxjq/7lWxWcPr4ALT0tLEw/7MLiwVIvuD+GJ4WxMMY0164Gd5iqcmp
/YM9ZoCqcqKprmEP+Yt8xJ3vErEsqjdHbuNtGdIeLSFOGFfAeloBJN6ctnlNbLKeDFmFayhRdnVx
9qtVluRw80dnI9lUgy5TAoxKcI4vzFmJ6k3nosw6pg9R7eLCaU2LS0r86N9AGfAadTBwSRFJpfR7
fKJMP4ru0BybS5VJKM0Kn0AcE0DjfC0KoVA5RIIkP8MfdwIXzi9/Z+HbDgWjXxyQxygS56+Q61Ma
jYAIvQa2zEuimlgMOGgr5bRx1lT94MZXiK+9WvoJUXMjZpq21HsezQ1+gPDL/YuaUsIlobMYGEvQ
vH3YRCl6qnS36RTGfd46+zoNW/XFffbZhN7ilG05X2Kj3c0OwPDYP7xLswYUh3/gOoyis9YHeygp
MDebh9sjiVoPC9FvDXESGPsYhp4wiyBPDeiQ6qetlkLBlmEkaqmd0IqR+YEQbfk20aX7C7LQ3+UF
arvWQ46FK4pnz0ivQhqxkNEqRsDNMXAfUW9NXedwDLdmJmXfekn1IPE4a0KLgz02/hmP4hy/zgZj
sYwgVsFChgLmG4StkR73I0PB70aaIDIxCr/fdkqvRTUjMR/Ulpa0pYA9i7J5m80WagItb8X6Vgol
SVYwp2JCml0zJeDSL22j+/0P9gy5LgLennYz6yJkXTwaZsDaTtH70VB+ZZtFLDjt8dlds5uMMw48
mkap8eJbs0dpvIEhh4TUt1m7mGht2Lmoif8xcp0xfFM8e0TPXIe0VlkqK2iqyaJd2BcoELf5iGCJ
E52M5F6xghHMkw8p/SuMpXKMCv7SqJEbx0Fs7qZZcMqeFpbbHcsGi7ODcpnZo3B3ucB7yytuTeJa
7rfJOnGlK1nUywpyEnJPrhkdECYZ5I6BqqbgyMJRRIsI1cc1BHKegykD061qDErQlBgugCogJzoz
uVLWgtvpQ1c6zXVkUgDt38eA+xme+ZuVpdhs+afgVrQEHIAMHXn9qB4clzCI7NCPZrr5I42P3q6e
sx2f0li/ce9uxt/AksRRFDBM/gV0PN7teRIGkvPUzDZgaUs1CkNQMO++ySuGI53BJiLhNJ+v9Z6C
jbAq6ADK/U6XhNXe8wqxGjYb2Q53jIcn5+ILMf0WlBbtoh13lQAocbhZJCZgcid3AlmCeeDnxb88
Mwy1fVYcIAKAxSmQjYAxiwSTw6wxr8tNezRcAjC32sPepox3pVymnCzeLAjxbhiEHVOBEm+2Sf8w
qr5elhXguVX24XKy9M9yrxuL/C6Pl+cUF9caAAR9AcebT40iIJFhTCguv5tpd/zrZpAMQafkZyUB
mmwTA937XgKMoAGFuPwuQNP8C2Q/s9YzyOYMqxe6dTGSSuZISc//gN7bESlVHKvatkeBZXE1hPF2
lxcQ6pUtSR5TlCZFkII7YDR6s5vlzxOdS1mSxQ0VxgjkkiZ6CAsak4D+qLy+JT6bNq3ZxBm+RnrH
MWGmFZhFqs+8IV8zKzAscaWa+NK9pIktHlxz++qmKIX3d5SGvMyURJTSgzc6Qy5d9nHj+NepFh6T
cF/ofesopTaYBX1nZP6PiWe2bW8rBYYHKiCbjRRmVGUlZInqsG4iW9ginIAUDebtsE0R38SxV3mL
oOXlz+APriy5SKeY6laYnmfdUV8rr4zKZ1Hfg/tnuUMxCLiYEMcWLYQ4ScUW5QMryPfid0GYvfi/
0pCqX9umvESoDChU1qLu/VGBVomkUpjjAI4tjj5BBLdvC9K21emzPtqArtvPG0Ji2Ye3F9GsiIUA
tcJ3j07xjziwYXpBgE9ofmSZ8FdRuPW8LD1jbkbW7/idR848i7BFbkcY4carmTpbktk/KQii0VWs
awqlodGjj5co6DIvFGRK3eyPNDupVTRYBWU6W0bL1sl8Rxwc89F0r2uwzP2ZLmPaa2yfQmwe6u5r
h4n54SStpsI7OpfRx6jKj6U53lGjq2LAhPntAd94lTvFkRcwbTxJHuNbtRYX5LIHBX+jk6LxcsCO
YPPTQs0kFFAagQbonUcr4LkIlydRjva4ra3DkGAardiEIve7FBFpb9bbIs6VlT2Dpv8XxEHt+q9W
K6C1FrIUPKmr3SgfcxVRbeKjrK8QUKEih6AMaHwDLNYqBiwaQKo6SubI2qBx9yprSHP+MDNxS3W8
Cjw7I/Y6sGqhdPDthpsj+Oy90MrxseHMAT5vkUcNohiXhmwO5homDkLfg9qMdu4Lx7eVxUAMh08U
ClHpeeroXNys90gXdeNAUdy3EXWIFxTCfbtJYTMxyPgjfy5W3aCZDLJo6Eti22MgCFqpAJhpAKBs
Y5YB0Zq09Tq4OFhz4KUmzRETe+9Qg8laJAmIj+ADHxLmQFMnZodytjZC5jhcJOX4FVyK7wZlAhzG
vhVn8XvLompG5Wr5PrnBXysLzfTv9udZQ/hM3s7/Ii3fKyKkwPVEK5Dkw9ozvPvhyeQq4mY7Nray
87uExsgmx87BdjiM+qlp7vMxZuRzBNJilGZuYFbBc+GK2VGpM88Zr1Fidqw/HgHs0E8D1BEVRhvs
p5NLCrbAe5z4GR0iTwMSm9tzqYRLzSNbt/oYh6hCXrgNnWoim7/jLFV62msZJcNi6dbiRHCqBz9i
s/xF1ceSCn3znzUKHIHeI2QuuA7ea9FWjxqz8k7o69kiAvmU8ymapc5EiU6HhhXdEMeo/YwO6k1h
BdC79qGsaBODsrxby0pHA9/7IOEeUp+KHeDBwSMjwV6DFzdcQrr08gRCC0i3+gxc45Y8ks/Jb7iK
aMRua0PCbRcL44qdqfRPOfKXEfzFhWDJoSQ9mmJ8QK1v3IhDl07V0saGixYqYbAd9VMX/LF13Wo9
If7Gx6IBxceIgncDzSgyLG02N0DsbOcYBtZpByn0VnL9eO6HWIU9n43yX97XuK5qz5RG/6ssn3m4
K1YhQgL2jEndDG6gPsvC4TvQ8Io+WFCODuUH95tJeRUgXvnuSiUg5jsq2eftNucpQqGXoT2zdya/
AL3++vX6vUvdBputf1gsXoODFGmj1Gjkyc7pNJKj2N3S+sGvfJZnZD55gsJDtM6IhayVzGFSKApu
33IiDG2zrH9RPeDmz7iq91b42kosIYYsD0IYCNLIeZzplg2Xqh8pR1V0VpvpR6ncLdNn2TZ/HOPX
7ZS7I8iFcAPeSWYqNsCV0mRaApZh8bi6vOtMuiHQfqYgWI1z3vIT/9SLpWVXda+8xVSw5KPoJCVm
FyDpCxdRPd7PT+DOt+dB5mJm9itICOlnpObP1ya7N0zLMUA0Ba4jKtVVKQMgVJHmgiIxJqlBW6K8
Hgs/r1Xmfty4P4mU+8JKSxus/liwtEUolc7yqPtJ5Kz+sOiAAvNFKIpnUbbGkru3MSh0JONrp/Af
GWaiE5/e0WMmSYTFlkxn2CntwWaosaOD8HUrtu8QHaxsXJwANSbvBqpEOQI1/o5Fiko8DrFn4Qkl
aniyDOiWDiRvGlmrA3WEo//XyqbpV5CBmf9Zrdbh3QZkHS5uATXqaqoKF/FVUAFFA3WUM6Rm2uqc
1FAk0VaQC2zsSM00JQGsafhTrlv108EXKVPEdI8p5TsS5dD6tgxKMJe79X+npK4uq0S4TAdq/YyO
6Y3gnDCSTXV8geDt76I6h2gAVphhiImDPAr4CrXmZXX4IvgWDWnzY+V/UoEGDQGX0YByheISO4I1
m/cNSvMFOattRQMwDRS83HZ4SsRmSe2ihBhMRGKkFxIhh0rgzK2QAfrJgDPBMA25ymgY4cOimH8W
m0BDUpttYUdyR4epDJggcadB8jDSlM+JGJxN1QtyfgIMCzlwY+GtTiQzimWhi03A5B0gpS3nAwqE
EhitvvmTxEXSpRKaBSbgvKtzIpMBsCT4fPLN//yBXfTquE/AcIoGyuYDPwbmymb/owtB1XVtSF6o
SiX070dYQLpQ3WM3iZ8A4TbK2JLRH/UfM/GD8ZZnBOgZZNtlPMKcXWImCeiwcLAcWCRHac2V4xly
sFlEtLKhS9nSsG45GioNJZSm0O8GNKFuCH0a9IVq59q0qYE0Lo6ZoGZdOIALKyBUPEWPjMvMM+SO
372TAk+a6GGUWKL9uYXXBDu0qarHAaPjZ5kNupFQJXEhQvL2S1sSjUN9P4O32cI5zvnt8RZgwqsd
OwwKuc4T5MAj3+ZYbOVYFIAr5s411EiWu46+7IubvmLv4l6pwPtJgwxxKcbJjRZSXXZcQTe1iWAm
ScDJM1p4WWrKpegLQWPUVDaTjGfszOrhkE8xwHPfQgUNV2fAyDz5ZsO8TFSVkhstIavTjuWLVOyJ
cYN/4CoxMDpr1IgkQ21vGLYgQv5LlcVYnADvaTYXK2gKioVSIyqHZA08Tx88c0LPv8UYwXfdkhNv
4nF30U1e5v1wx3zt93XS7ZUF9kN00xfB6UFMsdAlf8X0FmKO66zYqR9Chzq3K78CfiLkuXWE4vAR
bXilYIIlRikXzUNS3LNKTUFeRPHHSOOoV2wZMoBy5nokTZ9nSIEDPydMJUv/ou7c8c3qjKRUIIaU
1W1UR1UZ44wJWLhqXS1tzZVTTwpI+R6w05wPeopnUclJQLV/Etu7O2qhwg9rh8iVOj9nlZXh8OHO
c9GiqQT4KDG+yv1D0NWnTYDnHePDOa8pieUCNhPv3V2A9YMq7mb6Kz7j7bG3y83z6gsKe6NBWCql
PqiuWoVDkYelKKrKZhFqb4wPt8OOZHOJi5allUpjaS9B7/sxBPPEB6S0LYWrEtKJo8eNNVoAaPj4
jBXH9/2z+PL6qRh/xoR4G2JKfCaWJC37c3ZZil+s3o9+PZju+Gv9A2WzOLEjgZ/KH/uZ+lx1Zm/B
2FhLKSmZIzdgdLdImezVcaK5DhmJcEQOMDOUIGy785hlIuROxB+7v9Pp/qwHB94Swk788/NWXTL9
bmcGr4hNQPQbIQb04jvBmo+9M/InUdoQUi+FA9laFTQI33JWh1NXDwEr/Z8MMAeOaTwt58ZeRpil
gEV6lfxNkfUTa1ow/812pdJE+liSAGucurSwsjByWTcsfQbH9f7Fki2Q5u3dtVyYvo/4UESI4gfn
IXWyC1cNQviqOaG51/D9uNBSX943mx8s6KeWD11Ta1tT+pGNxIAjCn+gBw+t2fLK9iTZZYDn1BNP
djG2eW3WBmsWOohN7mlP+pQX5D86fIWn77abliSeD83x6wKWnLv1OO4IWOiG0LJ3xIQgUU7Liafe
bV34FEkuCNTXfeUqdZWyh4CNKr853vMV6Vtz7IvJ4gAmcEbeAm4mzkZC2G5FM1NtV3eaBnC0n103
w16Hi14+epyjkfEQJi5I8Zf0iKfLQ4JNRqGnrBTSmWTbc4evt6Wa3nEhGn7OK/W2TsJmRs+mu8DA
rWdI/jPhZBDjGtClWUtyyiMzvTT5M5U2a3//Q95q0/Cl9/dibs4tt9k4Cdr8WgvCtiBdNMN6Xggq
5ZsExR+eTM6rNMFjmQFBD8RPqtEMyx80Ptk9XQufOhQCsO3sxs3mpk4Vjj862uKoz8obQBoB/R0F
YASO2mxAmlpSy767jiTCKZXGfw0Mb0IAWE3Bi66wj8pxHHo78OlRo6vrFPd74uVqkMp0Y/FbqNkD
/UMH6FVNyomNi2uIjPFIQHYGgQStD4MfNsA2rq9rduHBYpTWo8hsFsqsl7EoeZYDwOgRL7fEZ7ht
l27IEPaldyugKYXvKtuaCP1Bj9nTWR8hDcBackqUh12x+YEm/UlV5Y1f0DC4beDtpza0RuFnxHWL
4sAxV8Ob2yJIhLVN4GV4j8Sktal/SwnB7RPdgMw0r6uCtKBFd4b8AOuEKF2lMIHF8s9Z5qsW7Mi1
wEr1Sy1vpFtEUca/b78mjz3uUWaj+baAQG+hap2We4qxGxf0ujmcZN9wUVqZOlbg9qhuZyf6iclo
5QoWhaIrdn0SBaVB9NkVKp9GqmQRx6De+eSClcdfaCofniARm3fgcLrne0sVptMvvG5t/hmDFWES
62QPejVUqkI+ZgAwzAZN0P56Rs/9uMIjt/EwsJSVeYgqzAY/6bleANlZ9IfiTpvScCQMG6gUUcrN
0bghWWl9/mVY99hDwMNBoL6v33pP6aHbPWZaTN2pXqxYx3B2f7/idDIYY3AzGGaagQ3zFeRdFAM0
tR99IRUpFPuUQoNBNc7myDYW7ho3TcCvx8VV659zcRdUL8wuT0JacLWuwBYFN6BalxfMltyeR4wQ
H/QV8U/+CCbG5kY1aaZ2TWiFwQNPPqYadiA+7xGAelj2B97XOeP2k9RZbhWaGEetSeKXAY4T8GRZ
XUzvU11cg3vh0oIMv3MkPPYk0dLXKSU4KeIvitj2bniOZiH4VD6iYMnId1Qnl5XF4HlsfsOi2WdM
O3D1DO+ftfNKbwxkC0wlShwGqFW3MRirJxdjeJdFEzjTLoUi+ISsQ8hT+WgUX73TDinSyLYr0VaF
VvAKpyRjGvye08W9r9m9janDbYox6W4DESQ/INoAt/ZHAagtHMFcCcpX2T4/3ys7ve/6MoOFO5Xj
u4EsQ/02rFO2/orDwTK5PViE8Arz22BT0Q7uKMS8JB4R5oUYESYrJaHT3bPH77z3y7s8MWXYiASR
pfPXaV+b6qY80C9PDJ6e8/o8VatN0vCjvhZhK4VL+/zTxcR8eBKRAwiJjYT3by0Jjnrcgza167Ri
TqXRZ0oSIjd1ojq/4uZYBLc+bI93nvlK0fSovbbiHhtYSljEAvJ/Rc8s/TBp+8m9Ol5r8pfIDuFs
dgt5zcKcbmQJjXO99YO1BN6r4kEypL9dtRFNwgJGBCRHDi0WciPJ3VgqRps8N32pALlkayhapqsu
0JtnCgOXiHUHxS48T8LvFdxlDypx5/R1eOE0oVEEpiRsFNvG2IqgU0UvpMPPdbOBztbdqUSykA/c
V78r7fI6aIwD9FF0QvcnclktIqLl+Fw94OlLUX1tjGrvJKYlEdU2n2TGm01fh2zZ95igzt/hK9yn
3enjuhtSR71NnewZ6Pl1b/avPN0IWBKeZ8yWKECotAiWV+oWpwsMp0Bb6/6rXDYMHDTLqUar8e2T
2vIfN7u4WQFA+mqvgT9BVESkE/asLTcP2rxHbUFiwVrWz6528QIuQqyIpulTssAEruQky03izmZF
2LOxSpbF7tl4DK7qFj49AJ/MUdsgEtRrUqU80nsTyjRgWfocL8TfC7r+c9CbsB2kRIJTKgEw0bYp
YMzL1rFUolF4o6KCs0Gxg6GCNPQQepRBYQMXxbFWDcUFctQRuRGe2aJ9nKrWjIHvT65J/as+gcz0
FuyRg6A0pPwHow9d3saUUcfaX5udjcjUW700AZvUUjrUOCM4B3BGfun9rVCaWnT4YmVmyedS7bpk
pYf3v+z069Ry8M7O87aoLa6DE8vzVObf5lfjx/q+Zu0YMpGJCjuZjn647LpdEEC0Rh7So7eS8hVj
BvEcw269MMvCnHdIuTD06wIDP2v6fz7Yfzzam5s9g1XxZYGFfLhzmHsIS4sesgONkzfQd+jlwS+5
SV7NEj1Cf8WGImfqaiyiE+z2PCC5mqXz/YVv5d/RFKeo08fdySuXdvc9KgiqT93FBpzI7iKunquN
ARGUEmELhUV/CWlj+SsY9MuERIyFAuVgluEk0xNILYpVSqVXQhE6yT1a+t/NpFXaQ8YhhYaMB7qI
3j7dx7wOYBVm9S2++nXcSYU8Gq4MYvj+qTS4DVpDSbiNXRem4mdMR6RUkjlyFs+NAxB7Wj1igqzp
8DzB+43fhPOUlKjhY4JJt7VL7MkMl7TNff5uvkzqE1kK4Nr7M5as36IWGKPmytkRaty8txsn/VMF
wyEo+r/eBalh1CN2nXUoDTaCIjRDKJn6XrgRldHyMdUbzMcWXqLQ/oGYxPpWtsqkPn0eBaRD6I8i
CjiGWMSaphoBR8Yr71x15k28yXU8vKQ6wPm2uF3P6gxTL8HwNUGCua2MTEr4SOSZoKmz0DVx4nqg
TrPNwPpPI9QaIEOdRgOEomd23z+ZwRyNOeEIGiExHS62PWefGi+S/KHVyUtD/AM9kE6YzJ9N5cGM
AnuXWhdgMJKY95f1LEn5Fa8mtGyeYP3SucllMiYLsRLZiw+T0mPc5/56bcZCYqHY6OL4x9BAE9/o
EmiWIjATXoclTwRR6+rB/HrYSlXlRTViq73rcxVilBHKQOIXPiZY3rZbzboaVCQUSDr+SDwv0lXU
eXTonb4EDrvFQbOCHlEdTYhz0JMJvLehlxAMhqRdLrzujtqFHIps0zic87xwGsBseAWfHmNQs95M
M8UlkULj0Smw0AnzjSc8UNdb6J14ZDnJKkkU1zXy+t1Ccqbtxwn5x+OilQWdagAObGQd5oTK85AI
JSQF1B7vt+ahkbIh6xG0IuakMdWh4kZXkRkXG1fQqpbemr2M0BHG9mZf73+O0ceHvQqnj5ynH3XT
GPFHS8sP+ak++df9Z/i/4wLEgSlGZNX357zne1YUjw3kSc6teH3+CWLECfL/GknEm1+kLZdLa6W/
wQIGyV7kBicbOJ7jLCR64FyxYCtfna/zoP4V5JndKwe2aa8RXH7JU2BqSP0KaUXNaPQnGRTox3D4
jouweVmLcIpw/+msuRzDizH+EpyjsYUvaiAvC+HFSwlFyXWlQa4SFHLGgVEsEhbInr/N5SYk/uIY
894IIrVuoViO/X2ve50S42R4mFkScqCI1762KBeyQMQFzYZ2qjeL1ZUk+iwRBOhDqYi6jDT7qIem
ofyIx12QyiEh9Wxr+sF9zTE4CZ3Za53J6Jqt2ThQHzrdh289ZLa0awXReVWr7d8xnfK/xPiKoigV
6urNuXMyRGnfHpAQ069ICbRVJbGbf2AJQ1zrGf+i4kY1BBY5/mLU9ahNBARFCPZqiJwH9lj4ljrP
J1/4me83n6o9iRRSCmjU6tJdP6nKgf0AXZF59XaBj9iTEZMytJGpW78jdaDsok9f651XPGShPvz3
/xCmX8VIfwzZFDMS1M43qaHYDAeb409WzSYy2FaRJjV3HAe/Osmr8lp4PABUeTgO6uppq6PtSSK9
XazP1pE1hJDy7PLXFeG6f8duu1P108lMJRzTVPye7YmMKajDUtScHcyo/W3x9A4h7JWryhfNAg/e
xClvhKAR/hnBVii8xQBvLd0sJqfGscfBcJwF5agfHPUraO1OFRjkZ29XFEViDPSh1mzsWww2t6v9
ahSI4zBvHmradKsKXJ0cWQcrH8ql90oIVlt9/Gmb3DUIXH5RRxDiAE802NzS+soA6ULalU2roE0A
/cw0XTSMXzfGscDeWbxEMUWZCWixRJ+sXZA1TYnug/V87pme4EnLwBrsTnOCi3OXrTkcU+D0sFkh
5Mr2dC15ea//uf/gdJwqB2ko0xItVfSGSJtph3TDpvQm7dv8ngnCFPEoXV6W5YJ8yxL6Qt8lW/2g
ITp6ryP0iqlaB3kB3jP5QoETaWn1SusDNyzt+cYx0xMOpxrQeZfC613tm3KS9ZEBE4RXCRnKtdVC
sjBc+PQTxzvlPjicYeT4xTGrJNg9tmRVfjh3iguudJAsF5gIaN+rq+7N0uCEn6RiynpVTyqeyIw2
HDQs7Jfi5S8w0EU10aL28fTTsv07Hvwc2B319KdbjgfgRv0o+WAeiNCZHVMS71cVWTPO9s+K+0Mb
hW8tS5DXLUXTPetRRIRsnofIrBjy3/QLMnP566VBLMjpu2kj6/AUMX66Y7rSY0uirtANVqnn5r+q
2eKBfLhkHA1mPk3xls6BZHATZ9aNxFjktCs40hg2vYuxApXudgwnBL4i24BDFGBrMlWiEEgQWEap
ZtUR/h3+eVXdH15Osl/+EIm464ZgeilXqAXMvFrN2a5MF5nSq6OIPQsz8X4trgoUSNDYdWbmaNW9
E0siXZ8dBZDRziV7W0SxjY483QEeLzZC46m8IWJoR4IKb+SWlHlmI5tFNL8qCdSvZ/dUTgMxaGSU
xtPw/TNZzkjCO6YWOerRfYkUV/Q3jSQMsaTiSy6TSYaPYRUjFu6z2wkqn0AdV/wuvJDrXM2QMHEF
ivlZIdo7t0S4HLriKxBLp3VTyfiepkiH4iXhz8buucOKzPzgq8o2zjRH6FUld5vit9k62sV5Ex18
JUTdZQ00tvvJnnx/sRDJeitjlVJkCr6+yV3KRASSuD5C7z6vsN7PilpSEAn3tlMyAbdlvDzR+n8s
GD8Oj6zJD7ohUHlnIAiHrprPF34RkFk8v923GhQQLiJK1RBocscDn2uqToT/pVaW4LquCBOU2Chs
fxzIlw0kOoVEzIbNbhCcPQzR6P/8RW8aTTUA/oZRl3Id6gFDygNsPKs5seXna71S2T/ghmHTBIYQ
SyjB0XmwEfTqmu6ACQ1p0cP62rvanxnGVyGPP9dyDzbLC7gZQY0hiKE6v94peDNMbqTA4SWVY9Nh
Y/E/GsX5QmLWK9ivAMcHSNz0ahNK99H3eODIbjJSoFzut8hUejXy+SHuoktF1heO0U8l+NprrGIa
dXUWiCJItiPgFnRNuQi26Ymz2x3iUQ+b7nFrhc75orZhVtzGEB/lUjFnY2O+y3ptS1b0k1iR1uz8
Y0pKxfKVd/iQZ4UkwPfaci5gVqIaIgD+wEsoj8Y7YnvpOuRdDHWoRUAd7oqCNaXoUo5bm1ObdZoC
Sudhs88Mhu3QpGQLA+arJnguWarMM+kYcN9wZOnoPfbTIUah7QvKmCI4vrXCw8SSLbcJ78SabHgt
o7hUO+plcESWnES790es1oSiiN9d82JE8W8eyQlGcCjpGG+m4nJLYv8VrmwOjiUoxUUySco2uwp2
EsoqQ+4ZS5iYRtJxYJG40UErfRSG7vnxagVF8eGWiQJrw9QtBlDFVpsWE4dd8hA8HJh+Bz9Pq2vM
8/33QPD0HB3VlFqg3CB72qcdsRezJtEjZJoaoYQCUj92pOUsnLW5vFoS3qXP6PqtvuxIpg/UM8An
AByBlMCHkF4ukhvMWPyn2LGFqYgDUav831f4Yw62OWYdB9HSrAzzV6saCrQ86iApkPq/nhwQJaAO
hdLwC04/4riBe0AX3n58ffotzCUNU55vdY6Hv7T6xVaPkzWQGfOVNih4mSgvjjWa5vYCz8XFc7Ho
tcoJBJVaj+TfNVGEnZCN880yVhwTnxCgf8M9GSaP4huAFtBVEWPC7K9U4U+IVqt7reoItQuRIuZF
599L3ZRnUp8s6v10ZL+lNu6n7GV9Ey5ki8KLXwTakNMBqwu2pRQ7Seara+s5hK/UvhSXATKuWTIa
oKtNtH/zyJNXo8e+cS5v2u5YKZeeOvniVVL+2yaIF6p6iGXkYgsDdzuwGvWEKvxo8TXfN0l25Igz
T/j5XbjS+fFZpyf0G3X3dtj6pyL5OEvFdUs765WmiIIAMyf2EI4we2GYAmuU52lXU9KyAAZNoo5S
xT6uQ+VXUHWpHzFaPlqO8ZduUM89P6D2Caqk9xMXj62PpA6jtz1rwL6IfDsRGeEA4E104Gm/9gkh
pw/seZiWpMwH/uHCzEdljwBvjH3TP0m0T3xNb5cdomeMcL+s4fSSmyQbfrdqYIck7RH60UM2p2Ho
0t9CP7ctDnzwh5DtZ+R6p4X5z84dVGl+F6P/kwY9haC3fgpx0JbIZ5JDbR5pmtvvO2YSRdDCqkfn
//wxrY2F4b8SraSllRNKj4L1EeXzYthsCvb8Ndu/+ZtngnWFGudmExPjt4g2h/PKf2PKHIaGTUf3
R1IraduV4mNYohHZC9E/5WxuF/SgRiw4AMYq15loROPZMoOr19ARSac6MMh/xqy/Pc9ScG8VJo1+
lSSyz56S1wnf6UgXXmU+8QQaFIJImIWE7qAXtB8ZhXywfq1GON+ki6Fc0n5/Tcl7lPSpuvgTsyaq
BqVEQnczxZYDp8fPfXMh4J6ZsAOnlfwIOgS9PUflBpKfwfG9GbQze9Cex7Ha1SKHFN4uVUds4o0i
2OAe/16gXn5aboJ071oll4XEjgyIypKbKPa16gxQrJYMfsa8KsEu3EUZX66RAqKab92YWXnzY/bv
xtT/B/HOkG8FP09xBbvpEpuhGcqu408VKPq7sjqRT4oCK2izlckYPPwedLueSSu93GyohD6d9rZp
fArfz7moJgCNsjHWrQAjLufCFt7Wtqba1+GB/E9jmyz4/7CQumN+BS9S9qQNMVmwu5I9QGMXgGMh
gFJNK227Q9X5UYzf+Y7TOKMAHJABH8odvZS5PcZ97M/7FQuOippcqwvnCz1Z4kORwZOhvWRbvGU3
Fz8jcmDhzZzp6IfBHcfZCER8DkQchU5BMNKfGHBtn7QRguJqtSMPUa8oLG4MUmFDYh3f3AeNrHBt
m2hYKroVsMSSJOdIclPQGmCydCHtw4wK8FHuY+zY7WBuDAdoyUn+n6aGk/pyKAy8iLjuy7AJOpIf
KZtkvODWKtOLbt6m4BlzI8m03XkVXGuXcO2qac7Plfe5BGigPxXt7QE8E/hbJd7yMHWuWL9LNq2H
vBI1o5+TSLfLQ/Ep6yzO0YhYNFfkwBSbBOqx8cPIObFRME+tzP1pWHA2hJVRtWLzj0/y7rssWUKs
6YYjCjuJgYfXiT3bRHUe+9TkrZtkyt3TWKe1nZKjnRpc+86+j7ydeKqbVHHhmE7XbMk5YWjcOToX
V/T3Dt8kiyE4Ufs1aO4u48HoKD8bU2xPdvriCQW+PLvv/65XJ4asVISg9Z9o4ByUJMb76G5/LH7o
F95EgYJLD40JuFstc5iAgk3XURf3F20u/e4NulIz9Rmi117a85ca+AXNS3d16zEtLnjtwXbTZTPe
qz0bhKU+P+guaPDJnfSSL3Qa5QbmOKDtoq+sPbGJUydwX7MOGgmGpfPGizjMdE97S0zgkWT6bKDP
Cx0Ic2CBgmVTt7JXFYF2NjQFyZgFQicHs39CWR5tm+N5LTGSeT02ZO4C1TqWDpj0v+MXPD2zWusj
ThF/T5TdQoKLSSdlK4Kf9XgOt7JSEkkce1Gc0shzYLMCDW8LHAosjdIAcJ6OvdjbW6GnMi8Hb/NP
2cP2fYeEjHUkR6HoNeX6WB5GZ6wvbfe7Llee3tyigpy0ZQLyi6qADxEmi97aNalGCOy/QLysX3Bk
2ZbiuGgx/r2yH4VD1vj6mWEnuZSxl70UxpYP6d4zgmBOMEsVOvJe0nKO8N4EaPfKE+hmcJ6C3lBr
2gkAChNGJquF1VYinLug8kydPzhhkviZNou3RbA7hDEe+U/C0DJi9Lr5ggSEGZgcBbyMu4RH9nW2
BDZz7dCA66GPsgFiMpNlbnngeOwwIjAwQHocqDN9BLQ7+Lz2J8vWaI+NTQn1vInVKwXEoioLxzG/
ZzfJGlpq9rDExIjE4XLKQCALkJuZdeudzBNjE+pQ9ojXpL/OJjW3KMoJCQgVh9hURUiI8BxOAK3/
1TxO3aoLzcrv7OzOL6xNRZQm4Y8qCJDBvqOrImXmXwQweaUR5iIw+4PNBVFQXpIOG7wZZc+xTYIW
HyVYZbHYR7D7GWPzMmW9XIVHI/2B7Zpbz1j+J9aEd7AqT1AL3E8le3blQPrdebF5dV2bT0sq3DxZ
eGk3+k8JUPz0UELSq2aGfRYCUalMIB1qhKgosKi0VeWZTw31umJWkQESGKtHfg0v1lE4ww0oGPWW
jZ3lQUouu6CqAgpNl6U0RIR6y1UyLrByc1OehBkoBzKNvKcNnFh+lbk4dIk5bKYpb1JoCCsZaFCA
8V9GqoaAjZQPUx/JQeC1CVBBdB14VLxKMZWfcMKxqebNaivq98t1fz/tcAD0GUf3hJxZlsMAEIg3
ag+V+bYxX5UWhnl/vXY9a6PVCEI4MbGFY+g7sWphUsKAcHmIKk1Q+qqmGNX1qEaLU3CwHk5XBegm
vFMJLgDM7NQgYnHoWdU4IhjtEzrDi+q+Ip2XorjJpyJ6MGoLpfoHivgZHDUz0wl3Bcb34NIuDfrZ
IxztAqje/WOaeaeBtBg9jJOxmeEHy9LuhTqgCEA9nDV7K8Av3u4W+2ralFnFmHE7Z3rMy/8OIIwK
sW26AWVpczHIe32PvmMnN/65pEGpeQlJHES5yoe37cRAAMmtJf4MAbGmllHKhCXj59E2sXfARVUx
ZEP/FG1xyxjqObBSIGCMk0gYuSJAkQX1+ILltctk/Y30LK4t8so0seyu2aZ7o2rYZuuenYDtgQkb
mp+kgk3sS2WxYJpORdVwD836DbFPrr0+iyELSlcDi7pi8xMK2Q8Ax+R1X6U+eIClvgko0BOLu+Pb
OF1+umcesM4jY6zj53zZVXgCXrsQxhkFjbfcG642qUJLWEUyr5fYK1sPIMYvHpZJT/QHV7mL6m6j
B3juo5yvm5r4Ft2hkiHFeaOUZbfHLLQyBF2wo+B8nf+rS/R2wrBOlRUhyAa2c3QNtePOJlD/NrDD
YF25MPP5Yb4/hNH5vYJubmTxgqCgW7VOncofTirDWUL0jRKmkoOlZSE9wTaZ0HSiSXseQ6nv7l2x
jVGB+QJYAbxCEuvzBIu56MuZ5vDqF3wWcED+aerTMnM1vvZVm/v3IwwMQ/voxokzwQA20FcT66oE
eCLsptjM58S7zS3WKoXGhRWwD0kYpwW5QCH8SPYcScM0SkkEyfwyIsDHeM2wsc4vRXIAlDge3cTX
sCWJ+NZnAmMlCnyDYphs1/8qz0o2HQvWsMduomMln5zT2OkR+SGa4SpwnuSQdY8KYvF2nBSdJsot
10YkuV3pLbNMbk/qrArLkSoQZHOjmdteX769/MdS0Engwlr/ZMtY7FIXuYbijfEtMPla8oikwcgp
671ZP536e3we9iEsERu/2SQBc5XOQAQ1Eej6YqiUkPVX1b4tMGZaF+7I6ZEKKrBm8wW1ch6yxL7D
1wRz9bbE2q/nTsi2Xn8FtnzMu9BhAzeHymf9+IWMSLwZGlkhUgYqV+6M4G87vcDsg2rqkukh4wUd
uuajfzNqSDdWfuMkuFFWHZW+Dd+JwV6kbZvjCo+AHoPFmuKWOcuztCe6xIpqjG7dfvetQm2mMmJY
UzmbEmHKfqWlNHcn6Im3uMmUB00R6+eYGtTfA5p3kSO69TAfdDlO27wpAcCHLih+aqiEXJ6QrqqK
V/Iyajn/Ux+kqJMdTLDDTZGnb28KcM8eAnWNe+AlYqeTAD+h4/CLj/ir/AGC+mAkhGdK6IfQrg+/
PJXg6GoYENrm88NrWzckUbr/liHgVfZ+NM5HMDQqulHHOXKsMWbNymkLGbjc5G9g9c7eUjYd0alJ
cwCv6Ihi+trZRQbrfxgTYo++TF36J4+iiUiUkffPObGkRYGVwa/dSsmokySxaEAqRgvufeVcC3oA
82jAErrrWVqXG7EpM+ACv8O+zxwJisLpe5e3N9rTdiUVLlsjsqd8/JcqMGn9drbsNfjEl+a+DseA
RZCM1JUxEjfPuq3Dih8DE1YOFVBwCDUhQmhLXVKZwtecBcatYFUwsVr66EQjI6w7WjjG2sTb9wP4
NCaCiVCSl7fjlh3+x91sMiWlJy3Vj1G72U3ncLU5qTX68FsgRhmCduMuHWoqapy3Kgp+/G+M9FpM
I2ylyjoaFdnWwZ4RzTUV6v3aZXwMThbVrlw/u7VSdAgzncn2FBTSWVUEfrwq9n8tya8zT5iMtNjU
u2wshuvx24RfwTjY4D0w+qBl2p+UaB6Ot2VNHAO02kySELtrhy72ryugRJKsQ9qfQMKCdyyKT5Ib
4H2p+DYab+K3n5BwbOJKIH9xIginaR6puDiVjAAr1UObeVXJE0xeLUVv/ILuwsyuKtXZAMKTu2oB
2GcGhOW6ZSdLmkW32AgConhguaO8u6IK59eLtmSt49SLe43VT5Bsg86zdJRR7HpibNpp0NRZelvi
YUlbwLfW1TrtOfkmPax5rikeCCZjdXaI+spNsH2zCIktFjKdhTzI9M7ZsR2xCJcFPpg6UND0WLkY
VBhm+uFJ6xAnEz7Pgl1tcRL8hteaZyI/7f3fGimZe/8Gwqvg6C5Twa+2B0gXz/ly4C8ZtJOP5mKS
eTTsdCjcIazDg1v6+/uUf3ieINXj17e5dPugV1Y/JRenvKtmHwXE1DtQEk7RVg2akWaxbJyAHfOK
spaEJaHAWbgEPC2VRh7vg89U8OZ1opo3Q1xRGMy4Izo0fN0MfEvMJzvAS8apchVO3yeB1cRjnQ53
MTg6C1p98ZHpaVZOPPyCCsLsmEadDmhUAU/gv1qDUUA0pbRoWIST9oSkAV+kRl64KsAUCeBR38b5
kgbPjpL2HHgQ9OclJTyduR1O9y+vMiMG+1HPS5+5FLQec7Up6Qw8Ch+7r7ht+VNzq6/KVPXJSdxL
j+rhxLPX7vtu1TXGOi0hL1U0YU0ypUI0kEa1VYwjKxS6AmOVTf29DJNVQ5rEwycmjzBJSOWEUinr
ILCLb1Cg3K4plck52AyhSPifemWLaxd/5sx4+KwyXNmy1WoMuxKJH37XramOOwN3+vU6LD8QIR4E
kGXpFziaxh+jZn6TBBjpwXN2WbkrubYJo/LOovttly6gOAZBamcJfUe+2Vp+q6tcVpmiTtDcS9KD
Oy2BBZSd9y/bAoF3rGAwTjvxvnJ/iNoDkCNthws1jjm5ClEIElIKWTxZawBHg8WoiMEKdI0cW1KZ
81K5m7PEOMMAo+vbHMjpnr/gdnOb+hwzdIaQgB51aN4YvEUQHlZaiYIyzpMscKNk7lK4nSa22NXO
jqwmw8BnVSGPR3p2nzH6PymFUs5sricuACFhYE8q3SZkPHz0u8PiTBJCDm9zbGJiswPFChuFqqIw
6FNq1VpwT0B8quV9l95YsqsKNw4MPK4MTLgWHxPTuXOUSN7jgnqaSQ/d8HVQ+8wt9B9A1s9/elLa
Mu3g1yKb4mo/y3NudXT7gU7jpDKGpqYADLgJcj0m5uOXBQR5LSeIPKBewyb7h/gNCqfdz54hDQ6I
Uawq+XiYHWD452KIPHMmVd8qlRvbGA81OWL1/KCBSK8OUWds4Hy0pyVLlcoq064QQ1QNeEwKBWuB
GpTUAqtSVqHuRoZ5vxvWKU4V483JcLvGUJzwP+zI12/1cej4q7jLVrWfly0iVLC50yaHQP/5dzkn
EhbP5ZkSck7msHSzrXHdNiGiTCsmMgsFR4gFqB5ub/4vbfJcouLuI6KuP9cys65TxdrfLx2FNAYw
l9Cbu7tVdoVzk+FBWy4C8UDPmSryxt+cJMqjiMVASLGlDrsWFTfm7KQsqvOyFW1ZUoxdm0TiLCoM
AHpv7W1nSPqAaqRDXlINj0tEA/DBO/5nb1DSbcnRO03vi6qrx3sMtDwb7hsDSy9PASYMN04c+2Sn
rr9pMHCaOLb+PYD3V7WiYRifBh5rbOlFye5TShB0OMvEkjpbYTykQSvMmlHuyDkEZXUJcqmArCkv
+yWMftjcLvtvrhePD8cnu2b1UNT4u9T3yCwpQFI7lXXPTq/bBqd3XzgkoHpessbXDkuFOq7gSeMt
eeRancGhOTmR5yjMXH/CJcsbKchmzTzYZEJmu76+XLemj8ZrIVAag2QFxVLMGPk4mzP3KTmn9jer
QP2lndXI7xnGrEIG/I6kIwI0Llm5nKWXt0owU8nfuMlXe5ZSYoDW7/D/tOciyNkPRqDIlOvKGqMW
FCIOcNQyb71hE2+st6BUIY/2hJ4NjIlg1FWVPcQjd7VmTgsC/G0t5QxXRYhJM7TjpB198sSCryXQ
43Mq6gVR2DZCBYMlEK1gFllxiLlB3zjZqLXS1Wfws9UkGZ+uSOL9VT2oQaxIzyV7AQiexN9QwMvr
vi5EL04M6j+q5Qg3qEtC4Ce2GHLXiwSB9Z5ACmoDMpjpUzT2XL4KgtubbyPZR/B//VkyyYbUdMPy
XQ2korsGFP6MziuzqKlo5DkFDz/uc/IbiTWFpPNtJ8RHzlqVMrxo2G9VFnc0QX2GnuN5+naJptaG
c6cGLxirodUSdNcBOlMrvKXi4AeMHyX5m6sivQtzKoi8xGnKwJrEChn7Wi24BExRBiTLbKnWihNY
MEAVDvRcvHruE1iwJOy8e61ymLWBgwwLKd7yPu4FNaZ1ojFdXd19odGlkgdiaLRJJDoFKmTedaO1
k2SZb4cZE/p+SIrnCrxaTm0YGWmK7N/WdcHv9vcLVe3+7My8sb5pblvGwpHjwjgPHBbJj+qVnhVj
HH29Orddvl/hxLOzZy+WdgprHBRjnqY+2S+WPiyne8wccgY36dB46XbIwNmgzbDFBMbMpG3wRuhW
jMAc5mGl9Yc8RUChlnB5Fzhpt//8x6r7xSuZOC92SiSVv1qT8pFz5fjrkM+8TOBUuBn/G98vjs6N
S3s/s1KA7VXhkOVrTUNRxb8sku81qzJIcW/u/WkXxSQ8u24O73TfXw6O+xVDyI/02DhrH6x0O0q5
vC1U7DSe6lbAa48ht5BNBCZ3uUw1jyu6fIKBosLClVh5OdIBg5ZoEZlIHPD1jhntjYH3jWtYK+86
Fpjj87kBFniCc89rLKF36NT9dTV3NlBGF902My6HeZrJSilQzWp1xMekMrCyR35l3RloVPuzHziK
UHGxJwOLCv0giwhNQI4gPiVTLB4ZeX1DqLbX+cWlLpjRBTycxE35SXIGd/GmwoPn7UqrRT7/zrl1
hQKIEGajF96wSWZ6fzVt+MUV7ktdluTg7nZJoJqwgqLbVkd1IbP0LdG38uz3vl2xy4mb7Gy40/VB
VK1BE/RCedISDav9d21wZ/2YY43/+E4KsC6wvpl+rzcjoqBUfuHj3cyHS0mfyytN3fcP4ZEwZYQM
Itu4BnFjMXi0da3RqLdgdTWVpjJfcMB+L9MmCqPdUk8pnEjmBAx5167PKy5W1hoX++uKR4g+DJZ+
iwfVUICzOdmWEPfGAhMyVTbCnSoTQXspSj9uR411mO3VG1DiqLvjxyx12tRpMleuMxTXLtXKA9pl
7HSCyXDYdUUDszhmydoB9QMDKlFAW5JoKzW4rxs9RpBNQvbjQfOZjy9mhEfBkRa8Y2EWKOrYZpsl
p8ndgmfAhh9AsGXawWCdK/2WaugpkDbQkSxiWwoPQDaDAiJoSjcEacwq0CdbOAXUjSi/zHhK/QFp
9WwNRczoTZrWH2oWZGWBYx2M3DQRYZN1iaMyGT2fqBtlYb1yBCKatQiZjG6KL659ZFHnAe3Slp4D
SdtA/I2WIE0vPIvyoyRVFYcsZWv5MDiT+hwtNTxgqgE0M9Mw+8SUl1/YBYt2sy6FGFHqIqTeGMEx
7mdkJsuljNJwvV5731UgFvQLfm4NQLr5gdGwNKPmWxfHw1RnHoL/IzZbFHX6/AS3L41L48xbkJKE
dPkWucIkRpYmTR89MOa7lek5ULAcWwMePKUvj+oH8JVzWQHtH4oV5WWsH2cLYec/u9xSJCwb/Dbv
elMKBQyokTHK2oV8Bl3PM9jWEqI+EBoK6Nyyochy/HPD4+70bbGk4XS7UNZSTHXrQTA/p8mrdN2q
k+ckGozKeh5dHCahNOkxjEGKOmTUF53vKxWwIqDJBTARgoCYQoYbdejWxpH+OzK7LZl1nCGOJaiO
I6O8mE7JDI0g7y0/e73kPyVt/rZF3Yym84k8pifLkswRRyUfjxgbMpdrz/AR8nmfoDKsaVIZxElu
YvRYz2ola7N+lAAuU+qsslfPBfjVnKeRcqF7oyQ8MfmlKq8MxpiZ78ghPXsdKl6G6/7/YKQsP1Ty
XyFdgj+dZT2S8qoX5PshpYOVB5cYSaCDPVG2qDr4Bq4llT3P576uXvU0mDy5Zlt/IZ4b6VcZkZM6
lX9DmOTbIYH92WDEU8u1fkvlXDDr2scX5PBIZEIg3R8h25xucdLn5A5kNQgxWuayRfTfwVwR1mqm
ylOoAvCT+QhMvgPyEvhnYs0s5UcJmy016N2wtqgaF/kKYqqE4IP1KejgWF9kG/JvIIY7vHETCw5B
dSjLwl9gFhI/rN70PQNkDjMoAuhuQL8+q2YtQ/IZmXhTxEy6EBwOLdPTBZiHm1E88oopEALIfbmf
d4W7BdRup2orYPglIDYzhS3x90E9fF75l4spmR2iEjOXyXFW6UXHlSZ2KhqjFZNNjzqjwz/wtwu7
yGAYclFjMNRjKk1+ogjRk1Wtg1h/PFeMhmpHNnqGhCUhxsfouzIgulVvrU0AyUMbhPTX6pvqjdDj
gNmYM53vhUfBknWjl7dzlB9yCR5aHSf6ATY4sS4VQdC/Ck1DyUbjzRsJkRHU3tYIY9IoYtVJ1Alf
GkyJV8YLqPh1JSstq81+Ej0VOSqyt4wkbanL+Ne0779Zgp6L9ZcQ/1+jXkey9qP9P5fkEpqv9NHs
r/ewnqgoffNBkX5PFWp7M6FyitORQuVFh4HRvvdjROudOuHK0u1DXXm/gWkL88I4I2xs5dvAeO0+
wA5nbQX4Qw+kZbg6YKOC752tGiND6aUbletaVFsGDhwQmq4jdoBfMPOr8vrBi1M0kFjc+QUoCmdt
y12LI3Ptapg50GnuBkhVK5ZUoworMRKQOC+TqvUrKEh1xKXmbg/HaSs0C2eswmLUUz5fBGFNOtHo
PPj5tqTtg3MPsNRURzU6kM4qK7KTgtNqkG5IBpuR6CiO4Yy7zwZUZ4X0JAo7p7eADEtup5/rule5
0xoOeA59WeLUanjg2z3KDr9y/NZVyKGgGPldXUY06G6lXre0xIBSbaDF07N2ca05SaC+G2ufLVor
L5VRVNFhuF0ZSn9V9wYndVJRncQva/sG73I2VsBFAPv7i2aldM3X3AbIa2Bhd0f3gkf9cflakW9s
KT/b+JjFWcq30pwfr9sM0in13kcoGClWxdpoEiCHfb4oei4cMkwOasirKk+A3gc8+MLe79Uu9w5y
0Weg3StLR1RUBlsZNF6VC7nlnhgv3pRQ/tdt0pwoKzjxf26cx73CikAedt0pdWlXJQsd8efABcoy
iIRKtswZ1Oy5c/xTbjq2UkyvxaGnGXGrnO1RE9uSnSudQklW01/qVvRVvcMexWLdy+i3UgPd1Tox
6kpi/CwUyLrEVHKzHgWh6J8Heq+Ckg34QwMtvG2L0V1Veu2uruL41x6XT3cByql2mXBLaskl2bGp
uC04xk0qOM8fD3Myq1CW1ihd35GHnQwzFfgV5YORblNYrqpwFF9clLREyvWZkO8Mo9A5+jeG1mcc
kETk1oHf2xp8uFPm0FYNhK88QQKLgWjC9Z1RzB3pMFKQ3zMOQa+bvt8JX0BGYW8jlVqsrd4c0JWu
ETaZWc5KqWllCI7V+5fwAiVcmc1+D8PXrIBj4SlHZENnyvGLJryDwuqMa+ACW/e+v2Wc/EUR20GM
lCEEzVS1NkcfDDd4OEvDojuv7msKN+3AkMiQ8HOEQGgLx5TQVlLXzbVypFw2MYdQ/kc9p6iaOEjl
LFEH8ys3VNJ+2O+P8gjSv57Ee5ZU0pIRN7lDRSvtlU3kfaq4ramqCYT+IYtNQoxHtNcvakysU0YA
gKHuasS53XOrdfuoSEzPvz7cn/ZpkvaPDiFtl4jUr2R9T2LNMA6HNspUwHrWJKMv4Lv55O+X5Fvh
JF40oktqDkkQ+9lfyTiKu2j/xxU+A6sCSMNuaeM2k/T5KuikENpwqT97qkjEEfth9LWojnlifnwG
+I1b5MhG7FrGf7M/lQXALub98Y3OCdBGRhDF/TrSRCVthjqJcMSFpUnwPkIg0YebLVrx4ZSYaoEs
n6Wf5r2ynT3eoc9k/B7GIXQk3BwB/acqPtrZ4JscSKe89B/xLLFyOkYMeQ8GWa0khFJDpyJOVLXE
/Om5T0Brb5XCPyYmtA7CHY/w/UVwsFtT/gCGeCzpxKyjK6Xu9C9p41zW0MwRpyPjDAcHVAqCQknv
a7ZnWE8Zoz9JQN7tqRLUlnd3AWW2P2ZpyUC4h473WM/AlmMe65yfGvfMQRbl4drAhwKMy3Wkf0mK
X0mrjMX4ezLXeziAcT9VQgpywoMXPTcyOiZgY95yCqCs5FBRx4I9eU9ZWPovOuCXYM4fTVDom84a
VT15q6z0+ZXDQyoosuDc3fL4piwNt41PVxco5Of2/4Qy8wi10gAv0gXJPMBPauQ67pzqSA/TfNAa
Y9574r0Eo27IwtbqAaiqW5kMPyMv4rpoPx3HwlbfSjlKf/K1AfsSkNUrQ3xgMXrsRwB0dZAcHxPg
ZY0S6/Hq7/yFgdDpBmqoqVVmqtkzoNdaGFYjBNlQZjzTBiJxSYgsQHfJ0IwBlbXcuauO9OApYI6q
7+ixHy9YTVqMmetO1d86PPd3SMLfT+GUYz+LrKTl6tdriBN0uxfnw84UD/c4L64dOBX+v3KLucdQ
MqtQJry7Ip1oNMbRLiHA7ZJWQkWe38qVMBtoqA3fibdpA/1KIex+s/hKvGXOH6426ppf5p/hJatE
np1pdvx8lkc/3/Sn4bc3x+voUnyWtwk7f8Cnqj71/ttQ0/7Z49SQPZKShwRutJGu6kI2FjV+Emdz
FOjn0w71JspjhEez4pFmuGZugSau9AxOiBWDsGmOoqIeg44v5tv0/JU7/5dX1v2Pm6zQS1ZFdJ0C
PMOBgtD+sPsVGx0hLS3R1n37bU/FlbdVgOHARF1+ZrRdRdi/UJGGV8FHr2QuumPsw2ai6DzvO+fr
sDnE16Owq8NBeIA4XqF5LQ8cPu9jFIdDygd1vAS7lEbkWKt4qaMxMHPW+iMYgjqVV07x4kmfQPxf
tPsnvtQKeoqga8JI3TlR8kCxYElQ6Ld8/cb1kgTnjYoWISybJMhUfW9rSqUG24wevOjqLIHL1CAT
ME0cZwJMTrv+L2ixamC196nCxcAbkZlURrxAwuqpD+hRwNI5JV6Fp47ay4ADKSXcEXm2oiCkMCZs
MXjUnQhnkzh06xTHxGcZfbE0HSI4lXoqubL//49upnXfql94fxg37OBuB6S4FCfK+rYUY+yQVut+
oY1Y+6b2AUuuVnUzFlGhvUmxS9AjiC5Do+3/7VhWt1kfEymu0/VAkiAEXqJdOIVnaddHG61lhQr1
/rZDpMuZuqVz3OkHfAZ2dI9MqVyFnPOtaQGz0sUBq/YO9ARUtHb3PMhyPdJcVXdNX91QdDY7UhEJ
KdgyndyTY48+FEWt04+j46v5ZaeZT2sIIeIiTZEBXGCZT/apAFOuBgLMpvEIo+E8MVIm21VvWRJf
gczfNR4f/qfKwGHJTKF5xpcbY+sFkc7v03bTM1q5JClgpqjOYJ8Nt5ntc8tMGC2eO0wnTHNIjcH4
08eFwQCgFJIwmWq66G99FpkiIN3E4xGTeBM4n0aVpgKRiMg8fV6xx1NfTPTMoDuDyCEBbT6KDCg9
gSXG7B7KGggFOJ78Ebc6cB8kU9wT591K56zDgZjLOTqKkgmagS76C4Uwq1kTDDYTzk0zRdSffFCG
ICxQOv20z0kZcaRhQQ20fSQpLbpCGHjrWGQJb6LE76FrT7OwYb1vgSwskGtmDuzHa91TKru6Y457
li3UWwgmEqU5zkAzznYdYLl7AkzgMbUiWjaHiROh/csYAjiHgmiR+Nstyz+xrQvl1mf1vP86okBd
JUBQkn9d4cEezD7Y22HRGJNjtXw26prk9qJEcH5FIpzXLlIu0tyf/0AszjCImYAPjrmEHyaI7vDU
IY5P8IT3c0yciOpWCLfMGGqziFvbpm04N1vuzuSzYs0xuVtaLGLt9+UKWavygku8iruAHdd5oo1b
06YWOJ/kMSd45ch/btZNRT1lUIlBE+mCpFmi6wp+BLXYPRzLjNFAOzfwhlvYWwG4dAem7DQ3W+bZ
14fVzwx/i8cH1EjWDBYXhsidH5QdqNU47E68iyIAZ2vjYIQGg5mD7LQInM5EKHMbqobsIQXsBnXI
hH0SFu3nMVeAE5bnD7huLAktcMqiy2M42QZelp9uNpzj5SEyM/+9pHNKHwkKevYv7Kafnu2zFFl2
lJf7qZcJedxUhmk9mVeAEAdpqbqIIwOeWYiQZefHi0qkXwF6RGIkCIOOtWBAbtv9Gx5GPqUBBP4z
H3O9RtiJxciiQyrCD/YSK9hqJDImy2LId4DQn7EaETTsTQ9xBwA9eLCpRkw5VOQrpGSsPfJJFuXU
eiJZueYUuP8jevlP9Ha+AGScx6I48ZxbIgcPmEeJyNKGLaSs+proAXND2Rv/Uh0rJOC7Nie4kcXG
ymYmJH9Qv6uCe5NkyVZrdrOyLJEp7fxKMECt+aLeYjxHCyHsYBN1EfXARdkHgNc5NR/Nq7Lb/5EV
5tRW/VRkRmDGpq77r2I0lzf12wQ0oURelUxY3zbSkZOMlKNFs06pEQ3k9uPYzXNA03h+Qm5R/o/g
gd0ZG3owGaDfRr/SWOeZHwnUfc9ljsuviwRT5si6YEHJMBfflffI8hZquUbiQmfSVaziX3cV0H6F
yjh7Rg/uBRZCvobkirQlokjMKP3Mml2aCN8wEm4MOzH5nBzv2bQCfR1hHALpOsVyg/IqmR4uAY+d
GJ3nELP4ZVIyij57QKrAeoW/sWMrZj36MYC+Vk4CxtbD+7iz6U5OlEMvdla+54fAqL6WnaHthJae
V7OwMzIvZL4SYsVHLP41b9Bx4DhjaRpUkUFJ7nkqtcrHX0iJW8wE9YK2+dJQJCs8D7YCu2/Nj/DC
otS4B9Xonxq0FWhJtq8gJnBnrsWtXcCGvO3hCsaIK96Qjf9Ucv+oZAYclOiNuR3cR7UxO3gl+w3a
YhdUOry4avDwnwaLzcg9KJM/dXBNvaJlICOt8gR4ZoX6sHF0f3ne8VgfeD49YZpaIJYbt4gm5fzw
cq6w0D4IV75b5aYPql1uSt02xPf1+PE0OC/avV01dB2giqO8lnIai7ABaXWT65jyxZaLc21PnAeJ
Lp+agLu+QtViOKFM6WHBJj6+SoTqZLwGkCIwLTZ2QZIOGOafvIz+8WSUXY9AJtuOAc1P5/cMzvwk
WYUrbqv5bQ+1ugOxqg5JUuQkVZyuoy4ajfFcyKH4ivhhCY6qkXdtTVczQt8tPZ0jpIULOkvxcm0v
1c5noYFfwXia/x9od/6VxI5F21w2lHtWbGxk9OIu6+9HZCJ3u9zfOaJLZV+BWVFTDdM7XZiK3eOR
rnFNgqAwPy0NNx3m/o2+rj3kUqlRzWXSUEH8b9Lo1v/rjjWwpmDyEPZcIEV8rSnWop+fxS+89klL
ixBbrmnDcNX4IZoREjkEcZIOHxfbqq10J40wOUJjEg5SJRtbdaKf5gNatDtHNo4WcADnMYLaSYO9
491dDfn90IUmFNaIWUj5DGiHRyu4fT0wwsPTEqJ2GjygN1VXRpuLHjvcvnQl2eJR9qqIuseV6X2l
5lLUGIkVuzBYdjqQFC2Zx8+Yg8TtgEJIm9/8rG24IIzkbvQPOOwJu5R9LcAIeO7BkDvKb2dCCmjI
PkHbVouyLfwd3/8vmYt6L/G6FGE/6lVwA6uRmaQvWTnTDwRkRmkI2wQPksqVcL/h/5nBSpQhW33U
rH/4zBmgv5FrLE7/sMTUkkEV4En0p8h9FOEwmCwHRPq+tdpHio+dp3qXLXwfMjXpueOEVtQrF02q
V/oO7h082uJ5k6BmQhs7xytTiYQk9EMsytjuEnHFK5e7vgFCBKkNPgJHJfzWRc/YqMx6/3vaKWNA
JvV0Rp6C7QobiYBGsPDygnH+evyRkvwSw+h50cT8NVgpsut6bi3MY6skmQeNa+T4Ck9PIfLuV7mm
BN7PqXo3ao7sqnPdWeBCIkFRBbcy3VDU4dbrHhvBcwqwLHLy1WfJyV/rGslHMfY+SwVXalbdMYvR
6+We606IlqKc3HUh+zi8DvXxYiEGIA9Bl/4pbTw3cbv+2T57ewdm4JZsEeUjyh5vNaqy7s5MQWuN
HlmfGTeJWEH2dRMWvW+NlIHnbCCKFonAs+Xoe+w0/bYXNwz6bEiX5XBfYE9HPx6LiruhV1mY566w
dG5vXmkPAdzf8L/Z5as5RcPuvjkEbsg7Cv9CgsBf80Ai9FieaQSF/x4TI6Q5y/i2yEpsrQH/+M9L
xyw7XqNecWY7P3M0J9kPi26vUHoNj1HcEH9vXb1SZMTpWNWFEmtK69SbpyMqMbzNcZlZIrFVo7Ra
HUWBJrdCyVomSOmiqL8nlJhiAQHqOtLtHS+rskVxDD3kDppFNv0bVIOyRCkxFzKyXin1PFVz/o2k
jg+ljT7ikF8gkLDu1m/SlTfj+4j+WCBev5trSFRPAL1I0oEChi0DAfw1t8ivWqLkPZN0ommYsuCG
TdDe2ofyvqUdLyI+BF9koIeJfL5miq6Zgxms2L3m6bSqTL6Q+rXtG29xf99uavCYBCC8dfTPcTfh
BzkxPtLBN4BrmJvKSogWrN/DCxqkCbYb2IMv1tyAyxhXqFw9/At3BCtH4kSfiXH93qJSAicm3Wbu
FsBQbbHZHV8prpBwfjXbgMF5H4VOorxAOrNdw9pDviduBnjpKTIyPXMrJH9xTDPDuRagHyHyLDpA
Q6RdtHRW4AXmQdTERGBAKBbUU8O384cCZM9DjlczIfI25F8FmWDgW1nXAeNspkEmgE9T0E6bEVYs
uhNddlkZd56TbHeROidD9s76KKMDrEkLRIBTNn1MW+e2zfh1KNCfs5WL/g4y8az2551qK52zYQVN
1STyEBXTy/AotsnpwegvuTVNbrFWVLa5n3Xi4NedT17Wsa1PX8J9RE9cVxEtyc8QnEYxtV+uMLjN
RZTykIQf3c3iEuYU2/1t5o3toRUO/bu4PjkO3H40G6rjfE9AEixCn2vo7UkWNnTWhzUuONt0kO2H
MDWMkPMPotxQh/eZUWJF4ndURgFhL2B9XkSW9XDrcMXdQvxea2Ybsc7fqvb6LODH3fT59bhpRkpp
MC5eExm8I8D8HGn5doesxrsdZAVg/oVTQyj6YJa5X9wilsSEDV4HZcKWqsHFkkjDyLeRyO0ZyD2h
0oGqnF/H6b5Jcane1ZvfVBjsSP2LjR0/qQ236Cp95kQgPCZkjvinCDKrP7LOr47JERgLaV7nEF4l
3y3/8CJI24YAq+O1g3tUmcQyrl4KGS3mX7wtmFqoLYnJMMH67U4InDpW0b6Gw5qNK4xbEoKc/5Gj
qyZWmVurr2SnNuOPfpxsqPpr4XNclSv9Eqf90nCepfFqAwhIKU5FHeqDY/mv5387hZ5STZeNHp8e
TowhttRzEOMg+hzNlejSqy05ld+Eo+gGtmg6/ct/QYMBmV55KyLInbOTabtDPcO9NnA+OdfyAAne
ZslcYj6WcJ/A03ISmXl3C473j7+cpNcCwI9mcW+Elw5zoWCZJSJUiH+bpQKDyYk+xivMKE6mDokr
zBkfbhtRu4G8mA6gdxDwdlDfY0ZPjZ7/dkoeh0D9jwEG3lwDIxSLq+qnD36T6f2qOBIhWWJStTBz
oIm570JbeKd7gUV3ILADjAngv77FRtU2eFZE7lDDbE9js/CGATv5QBl7+ZRAykCKv+yusnxYFZ/o
Sw6Evr0pqEKvH7oIDRysE/NulHNegEvuPeboh5gmxUiQi1RxSJdp/Y96tX4tLaT2l3TwaBxaT1iz
NXZsb3c4ZDxffooIORQcrTLxhNrpyALYSs0aHuPPPoVHVSyVllhDradL1gZAYIPtH0oY/nFURweE
ugEzqNVZl5vmLar6i3PgyEIJZqh7SbLhcR3Sh1r35ZptNpXfv3ugfHIuCjJh8Jx4hUOCrVGVJDdU
53MvKVUZR965HsvzjyHvtKXHfW3rVOF2cl32zN+8AZHZkenR1mJV/U+lhuH82sh84559cvddQtOU
iH8BIYoKgiHamNEi9NHDL/IJcVUkHZNhwaAJjGCt3kJPMofZK1Fo6OaqZURh+i2pJgoJf222SC+F
+zSCV5CC1LW84R/YxwjgOzw0JOMkzyvUUKNm9LkZCEg2G/Pw5ZXazhCC39a8D2btvVxgfAanzU6l
1UF5FXr2EFMRT7J8CtC3bAfDbimqsTHA7B6UZEblW+3zboq/0hisuj/EgaQuYJ0/9sIC/lFxHBtE
yeOuDr9dWpY0oP3sEvpMtGNs46iyhxl5cuYpYGahj1EQz3akDq5aq21w9ojdYbbP2S7gU2x5n7Nu
QEmRhZWnv8Hb0/aS2MefTpaeV3dQB3eI3m7i/uURSsqnHRxProygvL6xdje0hLynd7Lx0WhMmkf9
/MIhSFZ0h305s+yJPVvU2M1JsgIMwTTZNM+cm8kwEfUYaB0UeEaxtUbJuWvtI44T4eYcmCXSxU0X
vbQn9TnGIiV6dkpSdNWfCjDv0ILTYFg/lTDlqVnTJ1PP8TrQOCsKP0oEpSABn9CG77CRXEAK7314
Nm3vmsMFCRLOJwnqkuRggGCN7Hrbm/Iihiwi+ssHi6X7Xy8OLM8WsrmhkiI9IPr0D34lMa/i5JeJ
bLyS8huUdgdQGe7jtehPxDFPbwPqRm/IvIJKsJh1f/fZUGYSwsHBtaMJI26s6qfG25UYD0c+MvIr
A4Ah53W/ltEEQvJFON/oxQ5Zj9bPp6F0c/Vnci/+1xDuBGcex9bq1ejL1JfeMzgVx6maza5XeOPB
inUoHBZwNBV+baphATBTjncSobv4bwIfj733G/hJZ0qDYtJ32JmEhANOd7KzvJMdPzuqb2RdOJvq
hL5dZGVdq7lduvZFMZjX68SOLnPipbc3wnROpP0aP28uFPFp8F+Yh/xqtU3PsA4WuqmZYaaxJt78
hsRFR5TzVpMzKkdk22YP0esHTjXKJYXAfqqeKJ8bMyD6TV1cgLET/x+BcF4PWVe7kj7FLuOe6mIB
ACnF/ExByTvePf++7LinN4m4kaalCwZ+lj48hbYf+YNdilw1tV1UoE5GGx6/QsCkTG2z6djXYbg2
izN1nd8yKudUv+gcaSsgGCR1bdjVZhmHUd2aOgyhVZXWvvSNNX5maX+MwWlrSxy5v1cYKBP1qlBG
kC6EGNMJm1PPyVF6jekWmD2m9UDOXhRAlnGzDbbruYo6OxUV0bLEaxI3z/ANTJk+qv6s0ybqG8Pq
B14ryP3rIGHsaBwAMfLGyY6zBsuOvJrzv9v4+0r/fWTJyIEXoso4gcNuzF03OwDjTUuCPU79dkqp
Is2tK3g//GdQ9hh8pZxwlZ8iTtzMj5LtMUuA3TLHIbbYgtq10KISAOO2k03413hzKEBeXy8nrE+1
Gyt7ghJ3oDM6clL8nfv8GnC4FcJAcmJ0soifXJAe3E/lMPIPHLIBS57ifM0kdXpCcDGjiG6mXssw
4gnhm91EmibyvzjW19fBpEX19hmxg9TjvEI0gSTg05SZNfKnBj+0oKpSY7i+xPGpZrW3yI8kzVyZ
5bYwD+6ZhzVbsnXYp1wGroRgVJCRgcwHwycaD6P5uVnulAu22dlhmF0dabDxl/lHRJt/KaGMervR
WaEVZbYI8Nun6xn71gtaBlc6gEw13gaklTlWv6+hLyFWwzXDnNdatXhXyCqDaIbl6VN41c7CndLz
PVX3MfCLSeonV0gyld1PXarPeXNy8gerHaJtGr1IySg/j5jJ1Z2jIP/k8ifsXY4e4z14SRJT7UEI
GOQZMv+I1SAn2HhN5WQz4aUF7EZsH+ZUdJ7bF2i2nHq16OGsFTbjaRHuOL2bqApvtb8m34UzuC6c
hSoXtGXDznPZ7cg2UzxQ4jCtJWkekhYH4BBcJvjBfLL1t2q38RxVLsXPKB1pF2aqPp3rANWb0pa9
iiRw872nVyLpz60uHqVQeurJUD4u7PIDoeJ9BgIoKuvDkKIj53ufYDkDIzKaAzQ6jsFBTFhNpa7l
MSSfWFrdKhAzl/2UocIzTEdBpxM/1KSw1/9t/6SUuREIY8P6O+zgKG5v9GcR/uGy2QK4iyMTSjDh
JtjP4KEv8HxjiwMOpYHvk4p8YjJezEQJP2smHxQx31kF4oasADWfOAEO26bcb0YmYf0tc3qN7Y/H
0Uy9kaX2eRllnkpoCueZFCSnqI92rFxvurbDj8M5A2HV2D42BbxMLK+hdFvfbKju1IaFumFnqxVV
DOGlC3opem0TDjemBGGOqjRcIupQNQSq6nhSyWGys2AeMqHIEOIOoalCiDagEmP5l7NBYJ1Cvn/Z
rwILFVC0X7DMC/GmWxCfsVPW/0pDxQGlHmLOFXuNQGwRNd2xAaR7jhz5e8tfg2r5UfQ/PZ5keYWl
3Hr3QgmNyuCbdIShDglMOTob3F37fr84rGZjLaTHFgRRXAeL3CcA/D0o5R4gjy+Y7iShRWpQHJcw
wvsETWJaeypTYoXY9G5D4t6l/gd9fFC/C2j9G13R0+TEa2VAhB4DvgpZvbD3DPD+vZU26dv7xn3L
9osJW0o08pfJjUCfVOt5zDswgRFUWDrVPm/Wph20Vd/7ZlGLlOv9VvPPIrSXg57+5fyICA4NnPGM
k7JkRF8bB8YRuvYycEY1kh5xsK5gvzaH6M+8P9nsqQh3uHgyDGyZmkjPB7p8KjgKZkeGrzzP84fw
0wfSUsT0XeElbocEEgdyIY2VD3eChdZVwWBeuEBqDnyeNBwGcvGUtDnzjcT/WFP4ITkGeIIFHoAb
g0niaXIBPc7dnFWWR6JeAFgKVMsrLygnMAfZTA61HWiMj2dz5d8upxVF015jJy7tATYUOkA87GNx
tAcLIbzPvVAEB8B7qoYBeAokja8joRVXDB74cHaISvzhdzasTlIxIO/eupCLv2BOIJtBTuNfq5Yl
T+uSfu/8o/rK4Tjh7d6wjUQNBLPw44emVz/Etcr8HRgf37SO0dLJkBTKfy/Tu5yQheyfjZPRznAe
QM4Eeuz8DxzWfFhr7w9e6IvuCmVrpG4rn1K3giyNp2I6ZVcPjkD/qT877Kls5+RMMgVFf7Xjthzl
fFtAe9j0JyogfSey9b8WtDgHxazfJfEHsThhldhbF4WVS1/HBic57X6ajFBO2xdqvMwMw3hLsaxW
MXEFyCgDyjfzvrall17S1fxpL8nNnDyPXUNCLMW9fsfHEuZ2Ig0dO6xZCacHOX/gbGWrqj7aN+F/
Ncq0mf7VtJmOxWyUuxOYix4RvEVbbTBiM9qVGk2Epuz5DK7bwIjFC+tcAWDJNc6TSGwj6pcuc5n/
zUvSyRLYzdeBn5XdbbDVH/duKJEHGIozsBQtcXoOonNyK7ytt7WN7gDvm9jz1j+mywDiEkd1UPJ6
EOQGdassJNQ4HL+gR5rC2tP3GvzCYfTArqx8Bz0aXb0vMjWSJSM38GSvTBh+HBiVBv2Cp33cCrR1
RKjA83r8ukZDloq+7sU1D2QhtC1lsYVsIZzQ6jabTcfjm265XswfMPY6ek2SgfVq0aBvmQdiY/Kh
M+D6E/HVTFaZWUEdFgZcJigsr/K5VcvPkoNxQsfSF+rj/xksY97n/UshToCfomU1IHWU/MTFK4fW
4pdPbQzwetQDiqX2RNd0Q+CoFhjoIPpJ5Wp4N9DZyeEEOkK5uDOtLlDLnwCAusj7IdBK/2D34YmL
vme17CPcH62vVrS3KZqbBnwdYB9FPSO9/cyqZAjYYGXGC6vMGXQieXfk1zLD/xYDyr4HnNGGB2ki
iNt0aLUtHfAL1r5R8DmyLTcgjYJWGCJRKpxVtkjXUCXq1P1/k43extoFLsKlNCu68skNJN51gIy+
2Hw8maFsbWI1HzMFOyQehmTHs6q35yfQkHf5HvhMDXvFT9BPHgg2Zx9Ewyt/J/eygi9QSMwKolx2
9dowOxOjHgxnNhCjpvJsB9mO7GWFiN881oDHMvyUwnxiZ/8NuImMKUMwERdjni9WW8ITWxGCIUX+
gyIZDHO7DrEQpMIOrUNi2kv8/Sy73M3/WOWXOyalzkme/6g6NSvl50oGXDa6cGZVNC82x8vY9tw1
6/CqOg9PsqDamFUJJQI4gfFLPoYE0T6tMU9ZCOM7b8eJNA4iTbsLpKPur68a0P3jl7vnz4cnPmQ/
G8uEwvLxec4ZLMNvxt83IgahNT7bGqsSDf5E4nslXIbMgcCganQcemUdMHxjRh9bu65M5izFui1h
8XzpyxnrsVLuO3+Tt103MfvVwaC/XoMO1vJtwKXfhKL5clGvsDSNiK8WEE5JQMm/j34yvMiL6kJQ
1X8knsfKaKCMNBOai8m2mK9/Yy9MHgVwQXOeuNE/1iGEJebySyC4/KylaqV0BfM9wHPzVIaYlqxI
YE75SHvXIQYLzAXJyemJszLvY+v4V4oF5gliknyBhTvyWGrPNRepjuNaBqKnIUPCXfae8ZbqbYjF
uCEKWpaFP6pX02t+wgoOC6J2V1O922Vagnasb+BcOleotmshj4Uv5i82ePHaxA5029F61JyBzr1G
kBkc4SVk44ZaRxFy2f6DyJ0dQO5ER/2EZfYiZZnjXrmLfZdl52Eswzvxfyk9Ru9D1sF3W0VaXMij
TV89/oXBFRIWO6IzDj/Ckf62CqjhngRUFj67ORTc9WcxtV4IT+eAI80N1SUX/Vi0PHBRMso7g4WV
CKzX0faq+tHRcmClacRtSgkZ8BM1wfuMr6UjL0F79Anc7M//itoxptotYtlXwMV3xo8anBCfkaZa
fzbZ/HrpjW/pcGjMLfdNNi+buVyxZxBoCKmhYpm6iOVpiRwQdraqSZ/WHsbcZbzQJl5rgGA8ZP9/
Svj8mxOg2FCApF3SCuRLqZxcggaYWH8bSJyGCAOltced5GsZnhJMJfXv/mrc1zr3CktsqWwvtTrb
DT2dLGg/p9R92qG/qvTABd4Ae5FLTs/d1KlyOaR1r1Y0q/ZNaPu/DGfgFCEvPAdeHWvhx4PGYnb9
MjhIGT9kzHLv21TmJn/OEgLLPgX6SILD/9j9UUdpWQtwNk+ASJ9Xkrz6zwJiN18oiBmOgFjNPGQw
ZaE2gisB0iJYnTE0k2hhW65d3hfBBJonUKeUxMLoKHzwmst7m76wxHNcps6HDypBiHQ7/E81j++I
7llYXFtEUcQ81IREEUf53OHz/JSRVva3+AFtEDrVxBaap9h182t66EQXb7tOPkEn0SLev1tvCoAR
QrneiD89E8mwRLNOp16Ybci4EW4RFhztccepnH6/HIf0Olo6dSMa8L9gEcTueveMPZ01GCwvGbS5
sNvSE8Z2I35i416AxW0R++StabRXiTuF3ujOhI73niArV+fZLa/Ytf3AxKmlZrSKqB5udryFuYX0
7XWtnlXV4LO+68NdvcEITSzPj2MsPvAGUq+sC6BnNZfqTZLsd5EM7y5dGbRafpiHszLreute34hx
inbWodsesDZPwzey0Dfjz6paplcnogk2p0xcyCShJqzMEh81pfl5I6ub8vPp5B5xYtkTh9joX16y
fYMPpTxFXomOGBI+YhyK7gIbW22zynvoxi+SU8F7B0NHlLYRU4qLfo2aMWT2cVccF27polPLne89
ZKbU8ZiJEAc6XL/BA++HbyccISyiPEK1bpd21VdLhlRiLi0+F6BPAwQloqn0VfgbniUsqUtHpp9f
4TWZ4CAa97nZo0S/Sy13OUcC6AJFhfsPDmmLJObkwby7kyOF54OK5oqLV9ey3zU2Z1wV6tYXAIld
qjfmNhKBzHzv4EuodDDnfkV7zkCHHzxcyvAW7RLdGOhdaM2jg2yyVNbSZRW/EK6ZHqrypE1Kky0f
PSNc0twYD53aB1oWtpy2ZdEn8NoBcwUoyHi6M7N33+86oFO7tzfalURoYxnXoa4tT8Y7wZ3cg/No
XqOS0c2ER6/VP8fFWVh1wiEJ3v9Tej/wqd9eievt8GajeIxL0L+6ccZ5eJ3ZHimecCGPQywDKjcm
sq71n5arIEicDByjvzXn3eopZYLwXBpHmY5Fcta0Txqis+9ECtRKVeIn7MbPQFxkLVAni+c4tlrR
mqbUsLRv+ls8/LYBYWSPpM1URGrQ
`protect end_protected

