

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
ISK+8BrzqbDVc2hIh4k9UuGvqsq6yFic71tfszsK7KRf52jFUoK33AosGVUYsGH1pmrUc2NUQcDQ
LseNrcojiQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
CxxZHetyKRTjg1ePIJzq+w/Yg+inN7g9nkhYUjpPSXav+SKIAQvdh174FZUi0SnoR2INo+rdZ3gz
yq46XymO3b/3npnRNCCU259giTvnOJxmkrtnjRyUpOg8jB2jnHg/f/BlL3OJUGGiFonBs+6rnNvW
4aiU6ycFpLQsNzqRlAw=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
HZ1Kttz7DNn3t428AVZ/hrbCqljpJfsdfcEo7T7pfqxl88ELioDFFp9rVcvvZiZMU++45qS8CpOD
SfwcEjOj8ndwnIsrDamIUHs+Qm4vUDDq8EtyiGhux+pwMtpg8rH6kCwLDCkdk848fWRbBOGctdAr
AiQz4Fie2ectzKGEhjERjquMNqkQkhNIuEu/CSTnyD7KnG+FK+llVBavN8lxjWeDvk+quMyk8Dbo
gA/SdzYI7TCZkNEFS/PvF3Z8fPBK4pBWz7TyfdHacMjMkaPd5zGsPBmQy77xwc4m/sfhM7ZX+YW6
VBTILiYtg7u194UVgu4fHE7f45jr0jTur9wbVw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
2VX2NPBJC/FYSjnVp8ueqtxuxLgenRIKbrff8tdhuTb77js7o9S4OVH2n84fEyvr3hl3lrO9ekVq
VvQQOlQBg7Zv5/tFAeI5YFisgygYrqeX9dQcI485CaCpeN9nanYXhtHWROH+ZOYckBZHUhhjC82p
LnYwoausKSjsi+rXE64=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
HdQIwrCqCFDZv9OQZsva3DMtF+8TwiePvWLQndNAXK/1V46C6C4sVLdH6SK4FvPis45PZ52T91rx
x7mjaMnTgTVkK+VoFF3Ej7xzh/2PoR+YkiToyHCbvwHQXXvv3GAu3HyqWx9b4oOndnrx5Z1mco/s
lNgEY825qOfDqrTkPvvNBXThybVoOKs2SBHAdaQhQemuYVAjS7mEC/lA7vom+55/0dhIN44Q0vMz
6utkLeK9axPmrUz/LHNLm3BFQsfvacsQoIQe/Y7g5V8ehxANfnzft/Jgo74fJAU3odGS++0PsHF5
2T1joNptoFFljB/U6DScrAB2FxigoQal7I/OSA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4112)
`protect data_block
ddPjSnh9aoQTXyUe5rRHIOnBdNr0+O3yOVd8d9mFoKQtpASCe8M7soXK0jG8nLrJMB1XKTjXF/2x
sizCX5+deGTz6bUjnR6OC0inTID6PFQ5j6mTMlT9VqlqxkpyEk8VBsldIjNB6vFiI5RJ2xU4cPhT
uc3UTcSMs/FoP1z9xBO47Gz1skAfNCkpbcxVIEtwKkM/VdPgqtQBRBpVZ/z33qcCgfVYY8M3m0Lm
n3AAmYWahJqLu0UhMd74TpgnfKpmOq5mrBds4+eyHssH3abr44YAEiyYRPGy1ZqJVUSMaFnuFgoW
P/e++AYBdH+c85o52VgCoNH9T5JMmZizTXpj3w1yiuMzeyIGReC94U7iLjtMzKTnY1MBjRmlwu5y
xS+XTqGNueft6vUEmMxpli8tvReTXB0gCEAV3O32I+r9L9jvW3VB+9E7rxSmytlkklnJV+OzjxAa
VEgOvQwn7oT8+/cpJu/j8AMLkFqrmVI6cBUjjIhLYF3wK08V+C+fo+85kaG5dRDsRvJonRWes8jL
p96/j9v62mE7GkDz19R/TFbTFpnCpri8hYQW54d3JGPvStdgkysavlZbMBHWfzpql8Xxkoxooj5r
zib4D2ol59DH8zYWqUZwfVd6YaO6DCzEjGTB3u7YqW/YmhAhRdMkO0teGjf7Ixmt99NdTkFzOkfU
HIQLY6Z5I9bkk4DKScbbGMT5Qn6W1btRNPNPlOdk0scvtMLar73DAG+aH7JNsigyxxov1RfqYXAW
LwfWVGYsmtDgeoLEoQYc2YTdpTs3/LNM/UDgq5d4JAX1824ePe58K9iRwP1bZYwNgJ/fzwNBrlyI
AG1aKOdKg3aVJ3r4pJfQeLb8AJeYWft45GubRoac6V2+ksh7UgJbZ8fLMwO8BntEwpLubBovHrRC
0dCwrEu6a8encmQYmgofOrIDPePjhZdfPoEG7Gx02xrrvsrV2T0cQEiXlHlc8ySIGeqLrE4bFqYX
fazWHKoHAO7mNWKrFVX/cBLgP3fAgHnz7G+BkOis54WZyuKNk9M8MRSbUBY8x4oyuUsESCAwMvuw
ewbtfetcTbxtzFl+bS4SkIp+7wK/ST+zRLYdEw2iP8uE93uz68BFclXtS8J5StH7/ZPp+Nf50vd0
g0xukm7gOL03byNutQ1dUjgse1ANC9C7kT4Zh5vglnldGhsolk0+ni7+Cp+NQdldeTIwlXZqtvCt
IpowGeMq/prdigabAKHxwIOzRAyhvhHCCGe2POHLETmAjF4WMvUqbw0vk1b9Sc02HJfHQUJ04zZu
q+ulr1Y7aGd3VTDnXLbSzTGtJuQmjMjftiHGAV+mEl1cMwZB4TX//APwaggUMnUeAPNZ/DpvGfvs
yoZcs/MowkO/WCPg+x93d3gBWZg3qpDHUWyz+D7OH+/isnLVlp1Xo3XZN7/oCVzuaParwuXeHyaf
sGz/6c68GCCDj0mn9DnpcklVFsYWlRe2YDkMnKZiWAWjlNmA3kDiXPfva9oLn6gAO+aQOjzEtAMh
TX28Tz1RYxDbNvdcvfhsi8B4GT1+7MjGOSkkKitSuWo0la+j8VLlhHm2ZLGdVDMRVPUuGu30rHde
fxkWuBp8rY8oB86toRsxUtV5gMoxaD76FpF9XN+Gh5m/BfakA/t2GMxJOyZg5dszZ2l68GikAswy
iCCl1ZFLufBdmSvmNRvUKAMl8jOIZbzX4D521UcIyFmVRWlZmLSxsaiOtARg5wtkOGj0Lyg3IJdC
DlTkgEIzSDtusEdIRiYv006+1NQcV5hra6mjDDtDaqE5Mo0023w8e6Sfz/SZzQbE6D2aydYUKQrG
SKrN98/CdXD+vVWsyLItrIcJWgkXnQLtN2OeOhrCDHaofsqzQx3ifCsYFuPAfRn4H6cs+ToOXNC3
YXskBQGGU+EjY36qJIlcP83YgiWZfyOCGAkLR7g16ufOw+g+oqPYR4S3xRfRw6PXOZsJMFz+j9py
zaouY7OGj9jqiB1yzpdpB+szlH5NJKePkI8VX3qDxJ9J0cgHNNMv3tt1BlAcstsb8J92eo23uTlP
s8sVNiBlX16R+8kfZ7sG8Gpk5xZJNU2KOQRnk11B+gnlY99VGFc/EXEAEiVtWl8ByEKmvKs2GFMh
pi2UlZieV+nPu0UuaMGgGcnnQeVAjIPH6gsgY5llsBtDUxoKgiY0OIaAjrFWYSSQZN4pIRCOp87m
+5hLn1cYHvHI1x5AjTfb2+Hf7qmo2JbHMWqMlOiSzYfYi+2AZUMCukXB7MsQMeb+4SZ3iQ+7Kr8b
4UOKmRvC1RVWt5ythfd9MtjJKX2We8+6IBkRRxgpQ0tO40JQEvk5lZNKgjNcQCAGywc55n7Pjo9o
3I4WD02Y0LaFq7XPAbYvBO9Hi13KSkM3sc2WI/YL6DAeWnEGYqFdaJ2ellVQQg09CBtYn0uQFdDZ
4kGv1pFTNn0SSsPmU04UFwg7VgN/WvISxAzMUtW2Mw6jgZVLt1aUqztg+AIePdwSY4t6LU4W8Fcq
e3l8treVArBRaMHIveYxm/l7Tuhi9syVYlKEK/rlh0mRWS4PFF4ONRTWDTfvDwZoI5gG/7Y4JnB/
ncbbQDHxucZm2fKdU7TuWGQG8KbZeqT1Bg9Xv8HCa0akCeue7ltibeG2fK2eJEJ7UNoqxoI4FAPd
5ds+u1lzNgyLinMaIMDJerTf81nUv7cEBipIIH/8wkUAq4x4kS+jroqE3ggCZbqzB3uXNKLEjZm7
nMjJnFbkkIxdcKXeLJx7sfXoXq2UcmemWjycSo2T3OBhmAUSoE56R0/qfT5peJzKjVQvUQ0HHMGj
UjoPBeFAO5yZr0iap5RTiUUuuwflU5aVNc24IRlICzIfY5Eae6wDXagw+5ImUIJnnVgaASzMDQ2S
HAtYjJVa9C8sqYRDaZpifCA3H6X1Z/kx68gbtq8cIXdg2RL6u234OwqahXUAhyVGgKw2wO4F6giB
95B7lLeabijtMaOxW2F07j0h/Ao05RC44c7Sk0fFk4nH/MGbdKk0StR3Km9gl+/g5repGMNdi1RY
UoCODA2+5PQJ/9D77z08Qb4CspUev9qM3usKjfqhqOZrorpG13FcqSTHHRdGLhUZ8FNO8nv4Eutw
Z8HdiFwNzgWzPFwvO9ONW1L2Fn3NnjpUzsBDZE/MoOOXYC4b+qPIcmJY1OOg97S3ph7JgaBbmnfp
hfMzTshDGtg8d6HYRqV5vVYBBXjnYnAzfba6eix920BbHlXI8/1JEluS2LQdMt/7Gc6mKg8EN7m6
1CSC0e+D8CP6QDB4PaUmC4QmPqZgED2HBpqpGRvqQOcGDc2ui8Wg0mzxEFF25tkY3QAQ2Gkfpus6
TqvS+E07GTcwRsQiXhlaxckbs1jMb2qHds5tqz1qExNSBClqgCd/nTGeZJk6gsu9VFfzBQs1EgAT
LQGfciIAaHnRRpjDO3RM0zA4xkQnkH/GOlFJ/eyjFHDmoMIi2IBekTNT2vmuhXVcCVw/aDz1wjLh
NL49BWej0iQvbwWHOBYGIhKAe36Q5ziBeGnkDQL6JoG97fbLsrxma/ssav9ARWLvvlqTeFXmutYV
eFCbxsZFdOyhrj/XTq8UnDtc4NXzeMVHpn2R+Wat1Jo6HeuWWXfNiynYQSPN9O35qh70eCFZBm3A
O3oa2eYKaVbAZ8Gx5sXhATh1A2he3VHavnoSUp6xK52ppNCaVUiCh8UTBkgZsO7ijflxQytAaBIt
bDm0lBiIQB+Ma8fqJd94QCeV7tL7HMAygOZw8P5dhq9NQYSa8iElhxGkWCcfPFzDRziYXOlpdxqJ
drjV2TXB4mU7txjddFOYENmRjFoUecRuooSG4ixpcnrAg1qbLMbH/evatMrutZqNxhLn0LuFIbDD
fbaTnYES5GGgFs6aJPl6nl4I9CpBEPWLjAOWQX9rAWczAguwTIjhYyAEQ1GEWrVKaybVKH5RROqV
SHSWw+5YJp1UySQCOzG/B5DM+DeVGyklXafjg/TQlHzfL5KkF0qkD6b4q2TLJUGlzcBJ9o1da6sc
97eySpQLg4FZbPgw3n913oNIQZg/MsU7g+9UmoZIhKxfohJ+i7zEixXfAbbSvXcO4gQmmtmMjpBD
LvKFtowk/vVAq2V2EGltfWZKsQhN29uAtooN33exYmIs50mVpwUeSQr7SsTNOMUBVCH5ah44PePw
cumDhurSnuqNYdZs8/KlVL19IXNwVfbfsD0Pj6zH2x1OwF2mtiyMFqHWtfhEtUd6WhpFcRVr9NEQ
WFQ7oEOxyIvmm9waTB+PCPfSvKv/Imtv65TCIweU+4xd0nCm6LdH2vA+rtAOgx/K8faeL/Evnb9j
ESobX8L48mBNLGGKKpGxqJbVw9QRUbY+DqbnAsInL7pkEUDcPDZsvWutpWtsqv538awLehdop8g7
o1P+MYq1dBbX/wSlztVKlCXVCgIEpTtDrY4tEGHJEhK2bpLfmSPH+K/UaqE8C+F/fjhQyi7w1Sve
FWdgJi+EJx+q9lVE3zT9ximwI7uhw62ANNmVERtqDonzj09iURjEMfW7LM2UYn46s+wRHtMWw3VF
udWUjaVORNGWRGrbl/gVbpUMza/6bmQxKzdWRWidJEHEb2U7B1BUJhrtcABAddWzYo6bqZpTO5zy
dXkBbENnyqs2SPn0VX90q3YMiZkQqRfHDSXDrApOv6yZJKqgY34y3Do7POJpa280UPCp0e/c9fnR
35Tsniq6xZ3ruvKvABbfmXkoI9AnTW131HuUIrfktQyz2pHTe9ycbuBL+fmc4rObSEYxYAtZ8JZ7
36vqiaBUM+phd+RBlhWlrqW9ZYZ1XsKUUrUuxDOjkuumMv6bz8g2qwoyJ427rJU6DpQDeLyZ+2us
muDJgUiq5kHghD/UEDKDnANuAEYCLkeixpoS1SYcyfTQ8WBkM9wxV5mc9/zJMWTeJIw4S0E1eTgd
rTZkRr/GoUbblD8MU/YmAQiC3HAA6y1X6RIH3cKKn3qVVAe4zrwWh16QV8Wa2FxRn8VKFa0+LITt
lS2StflwLK8IgtcQSj+dUy74g0+LEig1CuDMSlrYyXsZl7A3GGoD/+QpLxhTEKDAHU8tcPahpxP4
CwPnrpSoBmQmsBQkIgDtQWGIWPVzxlwntG6tN5Zbwu8VMZg4IpRbm7kSAry0Hl/XEOaYr+mmNLlS
n1LkfJy5yoc5g3g5RK239w+8nYPMqN9k9Fp1kZkzZ5GIvg5EuSuoXz6/7luj27JkX7y19KdjmltA
NnzUqcrRGmFEeq8aHfhg6a8H417lopRCIGH/PMnhBg763+7nGhMMjS8S8/vY+YQ/6JIyK3ECh9tK
dWGl0XSaQDA7/iTBnpFviNFXrTFqWNcn3FopxQcPZZBTlrYwQFaO4WW+6HoyBsjf5Yt9WPHV6j9o
IOBdVZR4X6vPorlh95tTKwdjT+QusOCYJCRsIkILIyZnB7AVUNitAgivIZffVDllHTMWF8OkEkC0
JuQsdbU4ze4=
`protect end_protected

