

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
dpj1rsbRiC2XtvMMkZeaWceey8TRzfvuZghjsYUFfvEbx0wxaUtNO2KtH3hQvHr5R05ZRpFvbxnS
y9eflHJ+fw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
RxF4+BsurVIN9R6VPOZY6IjRgF7yOLOJFH+DEaCvilnRUUfGXWquiAJNpzEAXSnsWuptbwUxy5M0
I2FA4+Rh4icthIWWJqsNOFS1K2ZEpNoHe2hVsMzmtRpnsPL9VGvgfvA4do7AYV7YhTUgoQfClGAQ
vFYxy/RbXBzM3PrDcTk=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
OvIp9LkjFoctqOSaxZyP7bYL7KElD3vYsFbzOXm+yqBzueGP4aoe0+732BJK3cSRYLmSREwKo0o0
Rv3hIBpxf0Y7nOdTTISL4pJ3qn/Q9Div9rDMzGaVxIOMLNLxqjT1ZbqCGU0LBxVzmDxHhBalP4V2
XUBBBCK3eeYn9YA+pujel3BBQ67ibuZRmgjKTwyT9B3SaGu2w8ce0O/YfSF/l+ncmV9cvUhjGdBV
Dsus1J4qhNTtraXR3S8daDpX289UCjsNh8krOgCnmBNlKeEFeTxbhmhnNPIAjDgfW1fdIgrmAH+S
tzDecIht4fghpU24F+FmCjpRFfArF8+d7uvxlA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
4ZEqShxRoOQpy+XtDUXlHHAe5v38IR2wWpAtAq2KeZ3f4UCuk5LQw2Oc5c9xFXi1a9SsCAzYO6Rg
6iBcvyh5jboOYApBCjz/4VZfMAndhqby+l7lpAzkB6TqAqvqUfdVhSRn9DQMcQZ2fMALj61IBeLk
rnvtNe9XfB9vaA3zmlE=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
CxLbTp2UMBa44c/UwixvnmtRjPsy2Xb+fkOsP/coXETbFAb6XdUuKlopddrCIslByXBY8SiCzN9B
XnnZENqObWvYgo2VDZVlPu9SL8ZNuOrh2v/bJ7ztAhTSojfY2dBi8ojKva7J9JwGsRtKubJGASjY
RHw8CGw4rdc0A5dMEVmmoAymqmzBjExIxX3UWjtVz457DADxQ6UUgPgr7ysxQXkHN2eTr8eKtbK1
R8VALM11jq0MxZUpiiq5xDX4POkxGrs4QQL6Repo1WUK5V648ZRUZDaWyRJbcIm/J5ref1gzTZWX
h3koqZ0X3HGeO0DTx9nnC43UDVfA3fgk+YpVGw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 33472)
`protect data_block
S3iRadZU0KhZgvOmbpnjvXW3e87yjJC6p/QUaRSlha1QIwwAnguJWmjkaILYb+P1ZJSDBmJ7sfRZ
T40agnrGxJWQ7ElTp9hqB5SNA8ySPghxfQc30FEWAMmBI+yeRSPEMcO6ZoHkQ9VPmQIsF6lg74Uf
EcbWmLvhq71orrR5H5A7v+Db6k3pstGt4Xp54fKISgMq/9T9bi6/qBmh3Fp2OjvwEbVKjEzUKUSw
VdSGHjPo/q+IeE1dTOPG8OQZrtJZYKutE+DS1ugQ+1A5Gh7KTmQpgQNAq+Rz8K0KPICzB0R2zO8K
tIGA0u+Df4l+1DEVSbVcE7eMl0m2QANwYMrx41qjpYFLec6hZj1xSCOaqPUmo5n62g6YOFEDeTBw
HndU2sNePY441cMLFn3CPTZ7FDwpW3JE3Mqr55MQJu4kYlYNiDMKvMRsUL0KloTNN3TN3w5g+5mL
2+dnESE7B77Go4n3eG6T1TkEHgh/qUhHlpnZD1jBpAZ5gAP25aPNtko8vErLGPP1EgP636J3um+U
wi6fM0oUt52zeN/1d6unNF87PSa/j4am+pOH6FLJfbPGBdX8Eg0tbZH4AeFDkGFfKbPyHBPkmWOG
YfBoX7TWo1XTNTDVPJRL11QmAj7/a/w5lQlMj+zoLiX+w+LjenhW21iA+d+1ikmN2S9fUAwYPeoy
cVoJTlRERFuPFp31hySPXs2mx9mP1/l8tA8dhk8CvdZ0YS7rv13ec0pJ4OIqghkHgQVfevbsB1cn
gLJtbaLeX+NPyoBJPDZ6dSTa91GtVNd7wpwbgN/1QIIJe/5lr5FsMJATMJq00JyNqTMxPrgAozxq
obv8PXGQGzdbcZYjO36HdUQbKkMGV/6Hlqoj16hRvda8+blG/xVNoaD2qIXbPOAwChyVYy51d037
HnTBjNsOY0Djv/lbuTwijOPruOyCz04OSvZ55otMxblXwDSQCn0egygVrPWKpiDNVJUp2jMWZl2M
AiEVx7Ku//ec13qGaz6Bsu6c467Md1iUQ6wwGYrvutIhcDyugPhBT3OIaf027ZvMGXhswJB/OUQ3
J65okCGDEf9qUqXSKU4XCUSy72gywAB273wUDFnT7pA3FgJ8F9O0VeM58WD3dOkhl2KLujBfjBZu
xO4IGwtYLmXfSTip5ZEpXhZshPBsJPIk117bjAScgjGpWr7VVZlAHrybqYUcDekVS1Zb3CTxEzcg
a5yWxDDhxHYu0cRwaQGX7lAi7/gb8OJlb+dIb4D1G9Kod6M1O1J3KzgMAJyBN06a6oovkhNfZI1y
ynmg2o+F4mlkjtVNPXWVlImOqKlyVD+EIjdfhFb4p/eCGUVcDyHhvSnQi8sCoFCwMTQgS/JAxdct
Wk/3A0Bo8jsKbRO3CfIGUKlLJlyv0fdO7aEA/dhZnFZTrbZUUPbiuRnbHqcM1IRrs+VuybkUg6Tk
1eS1R+PttEFfgMmdih+73jcNuX5DGZjvkyCw5niNFwJ8pbYty8syZSCfbDwBkD2CBE206tpLdx9b
i32JAFRG/iYDpTBdeEax1fN4x47uhgtWVUAT7wYXgIHiU3wPkSUv8fhUvgexhaDbut9Lxtp/cutM
Ogljy3YrHn9r0Sdkna5au9Afv+QHWCecQqp5lfaDYlKftM1f7M0vsH9UhJEpSFdVWgfbhXKNbKIC
xk3ZBl48tlJp2Lrzn8DTSgxzUb6wUQXyyF0f5f+nZ/pz2fQlxm25GPgKekpS1/nZs6peVTrAo7F3
mD64ifx63i5xW5nC+BiU8MvTiT+5XJ33L7WoG1OKFssLTt1KK0DGRn1V8TRMvv2C002ppCrBiAeZ
h1hL+xfHtTdtble2r4e038TwvRA0CP/a3uhkSi9FWEV1w0oPV9nPqLJ2wUbMuznfcODSZpNm3orv
SVPh3KiBo11yd8O3FDMEAiyrAMwwcuNPOSbdtpVB7EnzhAe0PG9R51ueQQ0EAgG35g1DB98LNkY5
8KS8WtwTaifu2ymM+U8AMpD4EHjqeUVdXvDc/iG89/sFGBN0TKtNq/fe8LKfpJPOqTynbSOwwmq+
kYAUGmEXzBz/T6vhxfT7229gsdfdv8pZTstGvDsbdoKdB8y3e5AAa4BlwH0WARCbkAqadMF5U21Q
sMjmifjSqhGX36ORW/lw5zCXFXyFp4dXg5hUWX7YjAnAC0Z/v7Z5yibaGQpgmDt+3Me9YfjjGJla
tePYcxFVHOpWZUn42vuInWCO3a3sbbi25FYUSp5et9KVAQdbxPZc0bC/hQwWHRkZVLCtQPBHD328
VlNvEkBJRHTO0NEiQiBLY6oXSa4q4YOXTqu6xqaFuxYaNU77QdELT6sRX32n5tEesqAvNxTHsDW0
tpi9/I3AzWeGf3kK2NcqRzjXL+GR6+XF85jf10ExWyKxotySHRWexv91DakJJRAWgMcNuE5ZT3Zg
+l27TYiCEBR6qQhNCq3WJDhRTfxozjUtrdkcL0fi4NzHE0szd0bC55WzMLqqU8lPt2zZGD+Y2krP
dhROHWhCQTXLQF8Wzt+0lhY9La3jv3EpuAMCqVL0c5ewMg1A6dtgeepWXOPxZLIkWurjICh3DO01
E9JxyyQG8iPkIEKwYMQJXN4ZUbQjgCQv1yuqlgQiE1cKYOgLxxTEP4ZmHbUJ02jfEDRLMRcFf4dD
dUcMvx+hmjZBFZyWseAmoB+oOztlaWmWA7IeUamp7QPvt7TA2gLNJsAWhUXsNqNmeDUIi90r1D1e
rAflBIExIsskQjER2/ZFLrTl/IbnuvgBOKBNmKzVTDDRzXxKmOE/tgpO2ZDK/v+Cp6IZn91gzph1
hAgbCrOMVgZkLXb+/YHroMXSd0dYbeb39TIjgSRnJhST1+4pcX2nU3JqaN3M2zF6E7WKq48t9osf
AI93Gc2g5dsE+jrohP6NCusgjZ/qHab4N2MQ+fRqbIbb2EMeQOQEb6Gio7MGrI/DOSmxPH0BY2Nq
WodSeRlNhavHGh7ERKFceXTUwJIdeffSm5toipwPSpXtXNmP4wC1YBEFOOQN7FP0UzsTG2caJUOA
lHB1tutjMSMa8h1k+7Dengap+Ti1AfTMXSZK1Z14yj2OzBIT3+6N2jrGKdZHTAefRMnxs7ZXpJ0z
NpmGnkXPdjcepsSdaWHbmMXaMcD18+PTTfh+XKRm2xmzwNK/RaPqd5pCPOlj4F9fpyUtmL4lT2vt
6lvzayX+0lct7fMOxqZH7ZDUeaomihZ3y8j2c+zySh3vr5BBNhK99+IBdL0PSyICOmEM9C9u743r
DRsQUywaLxUoLWgfFylpXRm0hvrg23DHA9GdhqBGgKGEIvdqST8iqfAETxMRkEHJ+xuhLqwSQI29
0aS9uhkVNpl36/bg49XvNp4jbOUf0G7jWLxbZHDKxZ8wcTIGa64atPmhQyqDbuPPPUCsXwZXJZli
M/p6QCK8yUxkbcoM63btF9j0a53drSlOO8qMvT+8Gungdawkh4w0KYHq5ba3ivkBJxxyWpfGQ8dD
T3cUe5RWCF1kA1eqrIyDzajB+SGT2XdQ5PLHnD1Blvrilpm/OQsR2uxlHa0hGJ8ZaPhq7wzx5fht
1QBjPooHqJ7nodlgSs7BosIDo4sAav5tm69Wz76toEh+2GgqwdTgHZ04iYhhI4+mVuGC4i0i+TSX
cfbYCAetEB54yvdwfeoUS0gdCKZzdjOrzccw5pVvFmFFxL0h63SlDlF6JugdZ7BUPul3I9ex9GpU
8Bezvb9I6/qm5WCyxTe8FX9MOTMKsgByFtcPxWF4ZAMBdUWj7whoy85SD1QurIyE39nM5Kq2KGDG
nCWifv13J+sWg3rhr6IQAHS0bEY0WDrS54SWnvtiSYXmvQ0gL9zVREdL6OkrbkDTJRjnYKgDOYj6
9MSxh+J42zjz70+oxzVCKsTgUife+5KAQcf3D+TPW3i8CkRL8WNp6Izfo9rlNnYIF8EDzIvC7jNZ
ToPnuGwAifauXtgrfjVR7/JGft4+V//09ubXjtw4Bw97F+ptWGtJ5ZfBGOkOFQL/ziixQP91EFjb
iI38QER6QHhCZnrVpDdxVaR3d/l/5M91qkXiMOCc6b3f5fhWuYf3zPQapzXNdteS6YfKTyhgdoxW
v27hJP/cdUEAEY378Iqv0HN32Ea31NZA1cHhhTepD6BE04drBqfrlILchp9CzZg43tamiOxIa4ze
U5bceKnPzpB+xxOGWUNn0Y5/qby/SNRpUPKikMheYxvP49QhMxs79Q17ADGnqLKnmHn2dLWtMxqO
goA/7SU3sqSS7gr5sX2mUOI2SFoCJs5YSf8JpH3xmpdTADD4pmjdKFxX+r9wClvgH42JgglNpbOV
vXOtEeA8CkVYzXwEiSG8dTDc5klnfo7JR8dWf3T5Q3ZMtEE5Tpe7sVpAyniFCTVcoh/D8iHua2qV
zU9S/J8ahEnMAHMoGxkXje4F1z4nyHBhzq/MgGn9ZP16dWgnwzy4tzhoUMIw8Vp2r/UOBG7sYIHc
MELcJ/PVGHz+N1bIFuCZeCSEHqJbWPPVH3aInwn0na1SqZDrIgTHUFpwSS3xmbNenNQX9gnKKgi4
E3Wh9DuZxQ2ltwg7b7O/FnVsrTNkSdcPCpvcfAiaqig2QuSKVEXZLKAwROlGVTIln0pivJ1ymc1B
rul9RcV0INw5KaToWlWZzO4pLINDiw6PKs+UBpZCd14jtR8447/j5F2BTFNLmXmiNDsq93X8WXkE
T3Bz/LP173asBYdM0x+8hXEZHB/ffQAlAwpbvbapgnBpdB/oBX+1AQ9vaqQuDCLrsCyjPyEFcL9q
21UHcg4BwCcpztwKZTBKzQ5Y2gcul2+4ov0aRobOKHsHsec748W3JDCA4Og7zAW+ALJRhrkVC7+i
Uu1X6HsolJyfXWQSyMrZlEK4neL7KPhA095R1RHRfN5kEufYfWU7wbF3ilqSSioD1UlJ80aT5d35
jPh7COtAJP6O1DJVFPqgc352lH6dyRGcwjyOKk9LMdMYUO015Sdy9DDFVtyq7jARQsaLAHksE1ST
RW4jT8sMWwsaZPLsCLuGHg9Dn2KCWMKYeA58P/ULEIm3N0BFBBPOBoeKgq/LftTyKwWLz/EWd8am
21qjckNCHX7uG1YgvCiCFRUNx/37VrwyP+Ho2qQzzyWAtCcH37Zr6uId6tlOLsZ2jiag0UFuw1P3
qcMNStz9boHERVWi0Lmz/SosmJd4Xer6qhrLG4dAuvg4WQvaMqU9BoZb9ixY1r1dPIMSz2/StVrb
Xeg+G3fPfcSUNAZUVNVxLa/BpcRJYfpKns2Qxix3iCjXW0mO5LyVFOOPNRin/wTQCdZWFQbPFe7N
9AKKtHEy+QzJB4BRlEP2eBPiHc8wE7KUct8rJtiJeiQ3o3kBQ1LOANbAx43PASI6MwzrNnGfXmXT
dEXDmqo5IGKKlhfqaaypfkvsEdKBNH/lWm2XffirvYRVxWiTreMVepZZ27YJ35D0sNrfNkft2xrE
XZeWa/gNIuRtothIx7tx0E/9rXH1aIJTvfdj6OWgTeqMM2+hQNPrx4tEq59FDcY+uNBIIGr//odm
8DXWtlbtAEDNaXwONDNDZaTUQBBoZYTSvLm3yQbEhfLOdMPfsuNsJbKao3Csz+nS5QaQ2S4l/ZU4
ph87ygpyukWUaez7ndD8xlzui8ERC3EFFuIYva+sm40mGVnTdiVxeLw8sAWByK2vhZ7DKjsorXnW
0dGjU88Fe/cbRj5uV4UqmhG0bzuCtTUdo5zQgcRWx8ofDD2XBj7+MKd8HXZs7hr99c8a0v6n+mSs
LL8nHiZ9/wBYOGmXmHanWaLl340XH/vcl+Kunw6/UYmgZiLMiWGHtYZbxM42T25DzDlCvExyTBal
7+a5XBTNt2C/Ww9WjBkAtDJBrPYcwJ6rLs2R4fdjIL8ib2USU/s8k4Y+SGyr2b080WqPZWd5OQkI
7qAlMVnfXuJj9OkdL54yzUnxHDNG0dMiAPDcr3+MGWRy6jMEqnuvAAUw8yUi13wjbDiHkaVNDT8G
MQ7Fv0TmjsqtVGWw62l2Ou2N3KQ4d3rxRJ7yOWQ5WOithi090FhqfAp7f/baCDA06HWVxCUM3GRg
V0Az3wOO5dvHWO0lq7G+H3su+c+eU+UdARcMOZ1+CIkR9/SFiigtuQdrHcYPbmNwcrnfYk5ZAxbA
GcRldyd8mAl511SEMiZiILrwRU86m85g/TNDbAuwIbHDkVFX0jw45o+qDE5gbkA21IkvxC0LNVeP
HyECH7d62EdWORJO7HSm5sGnikRazaxbHef/EgUTse91XvemqD3O+DLPBQ4uh3fWNVZ1elO9mwX2
jdPP0U/GvEU6RkLsJ/soUltLRQ6Q3Ne+4JyuoorHSNueJCrrmdd/nu70j9UsAgTiW1OU4xY3a/yK
wQbOnej5Hl1KeXSumWmfeEXofrlE/RiYnCPd+mmKHaneTxrFiE4bTD+pfuusY1ZPoOjus0Myq4Ep
d0IZ97DXaqgivpbfmJ6mBQLX6QSYGiDjCVnjmE263754+nKJOnSALxEJYKiFneB7RY4c2jeEsMma
pspqkbl//oTzOZV+yCcahCIz/lJo9ip1eajid9LGzzzQEHLMq5cx/PGTkQapwDI3sWw6t4iA9UYH
AqTzLf4STr66ciE+n38+YogQmvSSqnXmc00gsIML94fnoOFySRp4/vgJ8hlmY/VoLvaE5H5jmNE4
5KY7yc6gOogdL32HJfVpK+WtCh/NqggsR3dJ/z0m9AGl4Cmip+rEL+TCnduv9dXyTbIFIoKV4d4s
E0qtsb00XdW5CmEndlPkuNml4mDM5QxlKXfnxoRKgirnJCbxkIh3lbdI1s70+TZmyV2AtIaeCxW2
X1QL3fOhe1qSWUEBvPCEX2WfmvIm+DPWembCY0dooL/EfZGzpbl/v0+u51BQUoWXPuv+csn4PceU
mUUXEYnYbu0n2WlUrD1geEDByLwyEAMsYMbomMJ55AC2iy/9VYsaKK7CiGDPftQO8ITDzs8hAo/Z
ag/vtjiTr60fYqxIcISrRFRzF0s3gJbsQ0lXkJdy2aCh67f1LPILgmtr7RDr3THgvvpey3jOto/b
z4pinWWkW6ZQk859GWs5sL2nRjpd4Gp38VfCn0CfbNxELsY/sDUdfbF8qYzphGSotfUFShHXekxY
H4yDVq2IKI421UeR78t0J0LuxSAC9qmNqLHcBRVPSdUVSF+eVp3wNSRNvnK/pLU+k4YLWiviIt3d
NJ+436lIgOM0Yw/MfwZEnrJdf02AsDD4iO8fHjiuoFVeAwUerdiGwabQSPr50s7DuvQ/5BZeBwAH
KzePd/wLvmiwQdw9JSi5glxp9PhsrV14JDpu4bRzYrPkzelXDO6qyZedx+Eu5CpIODuioqev+TJE
Adbevauy12hhWaLBMa8uLD0XXaoZlIgO5vihLMBNH3XVarGFicBENvqFpX5Y4A1Ld7hL9PeYofPl
yjFe0sfYef48lURMTDlmLhtoA4xEG4oYz70Jf/jucxgMgLw/ZZfXGPHHPnys8RGD2xhDPj3aBhZD
x0/Pgk+U3k/m6cYX4n790sfvfmE3tbHfqcW7il3aG1VBSr5yR6VMq1HLY5YWZwvQHWQUiNSnL3c8
dwuqmxHNgfbwrJOlRiPspwZCsMuDuzijfgl9GAfoELLdLZYZIr5xSLakokYOSv5SHEWG6t5OIoWh
spBUWA2aRttURYNf3ZOYkWfXldzNEKDf3LXfiuNDh2eFKROrFRGJRExAcUfx+9TxRG43DK05V8YK
Gvypbo2ST5FFFxdCkfr8vDWUnC7GKdmpBltIzQ7c9jOtk+2Jfg50Xe8Ob1bOIuUo5wqg1BDUHjuE
BxDPLpZwl1rPPEDGu/smPbGHN7cTu/zHKt7w5Ik0dI+xl/fBdehyyHHiZkVuEdj6pUUYHp25S+kA
ruKFdgEwuqMNDVgkzmXUDOjQzx6IYKVq/KKV7+VTVYH1YvjPe0aXoqZaTippRlVtPmwD5PuJT5la
yyl7yRercKJ9Pb0Kmu3KHQKHEuY11QZDthqkCf94oiA3RDrRUnIcSoHc6lgj61Vy8XqKPtapcEfc
oNsmJXseMqwcvecZqxmMcTTNuEs0DX14X2lgQ854GaRlqZcrWd7cSZ2LgjmbfSmeBcgP/MV33YW4
TWUFAWoI6aTWZlQ/9H6aatQiLMhg3bDYKT5mrTBww4zVvHbkf44BTmQhcSxc1SMfyLJCFjPqkaNX
50J6khL8CCC67PDD+Lc/2QZA29ErMX1Uyys5JhyCkgpSJDD/YtTTNWW7PUD8PHvWAxgt8qG3ZSZq
qD/UTJDglO8kh36PWuAijHCUIsVAtwpdeTSrX8loGFV7BwU4JBQ7wOBhIH8b8yn6a6Yx+uwq/9ua
bkZY3gL9O0s9y8NJXGsFwhyCXk9b2n4DwnJP2ZorLzSg7eakLMJBGVEeem4BRqT4FH9oG77s2o4O
u+XM4VOmXrFNReC3BxfBVH2Xa0cqftO/wsDRyDe3lLQRgRHU44uxFxycpcmSHPGt61pcplElBr0n
fhZpHSB8oBT8Nl4aRHqcRxMu613w3VMA+MkINFgPiOJT0rVPbzUAj4ZJ9CgX2bzuGdfsH9iDr0OW
7r8+qre1n035533TPOsTxJGR6HIbHbzRvWbxzM4N9ve+MLovx0BBB1gxEbIJ/OTF07UAM8Gbl38+
snS0KTZHWFvB5jERJ8HVJWdZgEu4CrtconQIB/8hWlpcCrvPk3UAr4C9YHa3QTBvYvY/kD5Aafwj
oBc5xGU7j1kVPd1UwZPqWZpPRX9aLSnhnEr86gxCpplpOXLXUcGAn7XcPBNtNvI/G9Ap/E4ooXb3
ajKkC9J28jSyMnpGFDhuzNWKJURD8tXp1yMfxQaBnr/+0YyXLS4iFe14Lm2qDJDeNymHScz1c6b+
5jA3avGyxgBxfccJosvsUIUaIxyqpX3gKkaaVaU+RZJ3+Px7e7eCHOq9qQFtAz9GN2pO+KWGrsOd
uRI4wiY7MYvwDZd1uL7gwBeItTVQH+G2IxRg3ddZvqJFWFSBr5Pda1z7JiCyXr2+VgfnGPP8MNSX
5z6SHoZYcKoKhfR+/YR+kyvkOezHUSwuDtpQgcOJCwQpFGtEHI7qs2lbrxOqtibjhVvyZ+fSY2TQ
20DeG02upQ7PAw3QE8jha+Wg7caAU4c6oEqcG2c/3FF4RNrRLti+zGPGP2f8DDbybL3MdUmowfw/
+KCELIDSlca7zJXICyT7vqLqn1xhOzxEOuVGDnaKeoXFEDQjbn6N0rewWTVffXYLb1sSS1bpTmQ1
3r2yViEs1p7kgmJtghSYnrTCPU92R9X5+zIxwVMjuFt2qVih4WBc9oX2V5f0zgn7Q56QC3KN/nD1
BAG/TpA3LKapBILnL/ob9qUoxRhOZtfab5MOe6G+amBw/fSMRONGxZ8tqkvxo4KiiS4lbUdxO2q0
ATpOaeoE3v03EVkSl4Qs6VbZDnoNPq8kenqBiW2qxzA2ufhBwTnSVSyhdpoqdWYbvfUcJzusf7FR
YqsT8zG6QkRf1E/h7ekwXEUgZPn0FmKEk2FR4FDKy+/p0mRppSryRLaoSmC4oxMIrNXdydRnHLPL
SRFvg/q1mb6cBOL/3xg77b6Q8f+JKU/UW3x2fJuG55WKZrfmMX0lYBDM33pnakLQvEBR4FMjFeON
TmtLJ+acuGh7lIKQ6uuNYHbgV7/6H2WQBEekKwgSF6ofKpIfKZ6s4xLZOiGtS/RCvgbZYyaIQVQq
gZOJgIgTrYtW1XYSGTq6Vpp7epaUT4Ww0Lyxklvp2EnhPxc8broV1H+byOaP6z2yNri0yNsXV0V4
AxThWvEcU6j2AzLvjTDTLgMmi2uzFrl6WFB3D/JUJXGPxjybEB75Jb7ykh8AKYfSNbHUWQI68COW
OwTgA7wIGIR72QylcDUB50XoNqklgO3VCvV7KGXY2iUeHZW8PK/lRQxDextmHciueJDFD84DEe4+
p49moTphB2EPHC95fjDnuc0XMKd2QeLIZ7Y+xje62XD7JLCKJ7EwKN+HmGU0OJFbXPw7OFskQFrU
pJyfJAO4AYzdOsPYip0ryN/YOVQMiZuqy90Fg1Bv+5Ewro9ejozvLnFHIypLZBlKJjG1OtsZ0vUz
r/pQaule/z2WUVtdjjs2mUpgeyjyuPVaZFdPjrDtI1QYoraedNr0EyXW1r+2A3KnybApwUiqtnR+
zuVbjDWJ657V3YOoCV+ZNMciumu9UNcTTCx9ohGLj07vgf09xJbreHBGi87kzV25pdggky2NjVER
RK4gQmts9PTBU848bZ573YuFDQgH1Yb5kSgYGyZteoihbmgQg/TpmOOguxuToc1CkrFJi+oKZfpO
AfrVdoZdLQi6SGh9328cPsHQm/nXRl3WrXTYUI8WQTIZZk6rxTEcSwS1LmJ5+aIPERnSdoK3S2+O
X3sPCVEObGpP5Sgz17+PPo5HnQrUYf2HZRuYV8oGd6KErGpCC1xtq43zRmiZk+VoeDhJgIfXaGjg
cyPXURubSwWBZMloGi0pFE/5BdUH82PikFc/MjEYRK1ei+gCFimWI5jml7JYo8tZvcelmOeO2ZpB
jN40isbvapeAgum3v0boaTBIgKVxyVgl2mnuO6PJEGXcjJ0Cgk7jfSpLODR96+Q8mTR0euk5WgX3
Usvg2ChXvnejMPBps6dcCq/DOuazvQKY/FeCIRdL8oCv2cVbo9nsor1GbwgWJJuj6t+gu2nZrrC/
n5gRLLJV+QmWluaqtubeZ7RsTbyBgFssfvOg4A9/46Yfwv5kio0JaBxW0I9PBisOHdJ8v9/QXqJL
tkM3XQRZTpb/8+HBIoexDTVBtL5KPyLXwx6D6ZzKbaoRTBFQrHC3Bocu6B8Y44wpNS72JUE3FKgW
SeiMSwwEhyz+W8dDUAqW26ZiCM9a1RIYf9yAMJcNkOyro8+djB3evVzFyxNqQLhOTBGq6+7RRWi2
XOexRf6S09Q271WV6wJEpg60wyv/5cpUWmlIAEXdokoqoI+58Bc6P2V/NZJHyC7N+sDDieHsgMmo
7wjk9wOlaS86HXTe1P2dvUqbEZEs1kAkE6a0xgsc2db19FRPpploSXlwCUHtP43Jfy3bl2KFg9S5
QSqwtZKiu+KGDw10X++c5gojzq0u/1dq0YiOxoRctraBlUTdI8WUvNBF87Wz2BAtrSGow5DViFl1
LVnBW/lxcAAn6Hg293NEVu2K1pXva+wopjbt+Bk+blB1F1Z7VmK3VgvXgE2v2LPDaW9qZBa7NXVZ
jCg7lqj3eQAVxEQNEV7/O1Sj4Ihd1kBEPTyXouLuvuYm1F3v8iRGTktBuhe6tVrtnf2kLu/fCHUB
kk5oxuqZu7dwdY0kpU8JTLS6V5U2AKTttVbQboU80KbcpJlvMHB4hPOYsVcwgaIP2hlZufvl06pE
ik++etZRBexBkxYqIz2WoE8I7REJSIM4nOc9QGU6SIIf6jZBOX4UCv+G4pdteIxFnyaHCFh4w3JN
bZgT6g6yIzJQ+7nQfD5K/C3AAsmY+zsvZ5ioNSk+gVUnkIm20cxpYfxcuTDD0eB9UmGzoyBzVga1
Nj1VUJCmPWOPifIDinSaqAxIN5rjLzYFgS4rRwfrKGBU7+qEcaBDGEQKLhglmSyuZMdLFqYWPUK7
2FiXENqf1HY/ahH44hM4RIRhKiUb20XqKKkO6+W2eL6FRtRTNWKfM9Do/sAN9i0muc6pS61rzPvo
Cmife1xKqUfLQiEWBUI6R0pNl7T2b1T3rZuvkaEfSU6284WP96IGTM+miwkmanloWeCZzswBY2Xy
5m/aWutguXuTc9k7tkWoGVfOyj18f4jFQUcOvhxEGfov7R8YJd1P/KTJOsLvmCvr/1H4FnW6h+HD
q8ydm+wYhDq0h5Gv8H8Y2uu6rztPbwPpCUmC3wVtrTaSOhJyvgOc49PfYm0WRT3tkwX2DIn3svGT
B2R6ZmvNUq021WKjRSe5zEKEuGn2GSZLC2LENuF7cW/FXaOi4BcnorC+VFBAk7yfyHFf0mitfKpN
BVzEvilpsMr88gC92RrWon79xBH4BCjEAahaMouieK5LpX/2J4/fqSqQXJYWTaFaL+rGQp6jziVj
ZXBGqbTu85y6Jf7PeflsN1hizc93n7AJXhqdG1mZXoZn695CVYQVcbtUjHV9059Hqna6THYyTFEd
0rAmqGyVw9elfpUrA2EsuA14xwfcX4uYwzHWfq5NX3QmTuNEBPKM/MLC40bB8S137LylhyzbE7ZV
hhzjf1Avzvu7xDPxYizYxSb/MiAal41X+4LfPwhu7w6QEGtFATUkn2gjmrtFPBPLGqHVzfKeqhz4
TWSnR4T8BfOb0JEwgkBn2kSWb/tak6GxLUcofGP74J/Q4Yeb4P7tovwbLxYHUuON+TR9VRjbpmOb
PivBWxO8O/AJbYCRbERPUgbdTCMIeUtngYwj2ZQ9jo/kVn5UNm3/74819pH+zCGP9oaVQM1zIVE1
Zu7ZGYLUKmBUikHm4TM92CQMfjU92seBxil9NA2IlYf0O/cjsPqQLQwMEKWPHKhStLRJFDZAfFRs
kaTFfrF4BWJIStOnztMp07hVofd1d5a1D0MfYhwAUzzvCfbfG2hZvMVeHftBd1VB4ggmZrwzTjbP
coUAqeYZ8rHlGlorfncHvQ5Fgfc7rEYSnqVZAcBuKTSeSUXN4W5wHIQB5+vCeApIRKtvhDV7e69t
N1H1Wkr7MNHuTFw33IVVMFZderhfuiL7HZ0ODQjVEiAWVTqIztx5iVkWtC/jRgWaoeKIgLGIi4N2
VVUQ7WTx+HXgflNR0NK7UP/noHQxXyuInjp2Upa2quFpNA/TlPYB35b+77ZU7XinraJxB3FBw1aV
isMPZTZa7VuiXL35DHbGyNhSZowb585fKzmEPwzhO9Aht0HxXLsg2C7q4Drm/nZWMAygHOEqCX3q
295Am75ITJWwenS2rIUUOqlOhzUyvGuo+9RzT2NdFfRKQjiMPwklyG8nsQuzGdTuC/atBmP10tk5
7xETSg80++VHyOPTdbF8ITeDxbJ8yhO5y1HMQkZ8ISlqB1eJKBxDsDVJhLQTNlW9Ft96ayb330M5
TsqMv1RF7Dh2m4dm+7jzNXXkvudyD70Zd5x9eDWZAB4rC75RRUPB0hcldRqslP5YUtHTkbxHrfBG
2aliBsl2HUUOGYh9kBpGfSsJPWUfnAvt26KuPn/YyjC6hAA857Vocno8wC6NAYq8JJ23RUaa55xP
bFoWVXB4n8F9Wcv5tOQNAu9cVefuYwuQ4yKVT9nhJTGfgdSrBY4DveqcD7CTUMIRDwif+c8kxcto
6qsCdTm74YxpzocNGntKv080cM9Zxm0PRQQavaZY59OK9KBZiRbvG8/PMJlngcJ44p2r5YnlZkAC
80CicU52Kv9v645NdId3Gi09km6jPP0WZmTH2l9KpqZoUW3Rz3YHdN/Y4VjHQ7yUCdWbpj5XlY6A
VsPp68QDtPjNll8/HeWVBwjJiOT5+zYAmr3BFIztyoJQG1/C4Ugdu3DPDgdNpklpsHQR4/Mo8pAZ
mmkj4g6jZPuDiUSA1Vl0LYnXS6FyE3wobavM2Z/YLA00JIen6GmXUlnEBk9hCsYq5JlkfWlBuMy8
B9GIfo2Nc/k5C4rt1/4ky+fqOxWot6SDQYEH/W5FU1YDHawFllbqTB6on4SEbNs8mSsI+LV1pfS+
E6X3GdxYZLNHeNE81NsAPQyCKTzCXUwipANnVN8Uw9xf9vNNyuDj/UCMFvnQddZFHZmjY3ZF1vW4
VP24WtTcyN2yd3/kuACJ8xZJUBDTV0yh1Hpw8P1kM4FaWnBw4ZeBWHvX3Ni0i2UwnWzIMhbe2msQ
/Ird415Jw6EAiLi1qaQiekVKfcMLEjZQMS9w36yPMx6S0rNJNOLqfJv4Cb/9KQZEe34Qza1z/Q5C
G6KQcd5RvcysQflGEvvahUEv7XXReqvzLyU6h6LbX1l9vdbWZPD8eGfgCIa3cvlNnFofOpeJoZh0
uvS/REKu48qlxV1d96uhCPyEnxbmLEqOg3Xy70YYLSbqJWe/BXgzFpWKz4wC6lpIRTMHaCnBIipk
g9ezOvk3y3yapey3U8dS105nWDjHDuxIgv1vn3tR1OXA7OqifrIN1w3v+c7lM5tdQ3g9S/Rm4qxx
ev5LJ1OAxFno7QR0yM5aQOJhw5GA1R2y8eS2YoN9I+Jd00avC2u0t/BhENH0bbK4DE0H210BE0Qv
TL6KFBR/NWXDHdX9K3qfmmscxwjIMPE7/VS/CQ1i0Fj3v5vlgEcKXd40eaxcB1amNPA5A6dwjtTZ
H8scWpE5wlrhPd069jLYbrVsB7n/u+PFDTnp6iqBKP4gP3NquK8eVuJGlm5AOQhDA1UymcjkC3gZ
3Pa2Orepczre/KmWjHQZedaOKF2jdGoPqGvC386pP06bFOK199GpvUbwsQYjoWhdxkXr/A0SOpcH
Dgk35rDNsqZXj1l4DNfWIlvbhVDhefTvsKxitS4dcHNBDza7Dz/LSg33nVFMfvnc2xPB45ZXvlbd
YuBkkaiU6SBWSULboBjWOCejJ/mLonqxZ0WEXZaJn9l7Ig7DzCsW2ARa6cIjG/bOINJxlC/OHGX9
ttUt9v0AcqHgqkzdGzJA0m0T1bUQfFyjuFui7Tk6mgxWxKUi+DjS1uEVP0zKKgefu6sCWNTOyq9e
vyOJ0IXeniqeVeLKTnOP8KrRAvHto/ZEsru3YiZ1nFNW/uqy4oSmA21rR7IiukZUNG6wF8G62DuM
2cTM6KVeQupX8tYqzbJ4+cLXW88X9GyqD/QtN5s5bXtV/7dLWrudq37vPxURw8H6ctw9BZ7rXNN3
bwevhRtSyS7Q3r2SuW31/pWRGIUebcsTPCv+u6tFA2CCV+8p7htZ+88eHnkzZJo97dcXzeGVwtLj
j5KrsY7DGlfWSnTptpWIAQfAMFHDmmfgB2au1puwdXc61XimoMuiasSYyslxBU20DNPBfWHBlq0F
/6rk2NHjGJsGAGFWOERU/r55dVbHx22xhMIenm/JLl+2RnBve+KeLcwaoeXPeV3YM5VktjUbKdip
ux27UejzrlJXtoTYTWy4+haUid/e3XWsC1eSwxjXz4gcZaD2kh9sDJ16cwfqrVa+w6qnCZttzNL4
9jdU7flaV44RAUy4ffrwnJwfjT5Ja5bgcReSfikrtWFqmUX+BQcjmvTdBmzet3sp8HF9jU3eYHR1
X/FlG8yt79QIjXKWdMxhVOu3SaohO8aRDYO0KRY8idt0dPLldIlpsu9Am+yfzUmTWFoyUR260rM6
CiavViLflTrcSNFIv9QFCX/F7kDghj7zOwCWhdbMTxcQ3tvKyZkW1iIU+KlwIxLXvYCzTh9Y4iJQ
ZFilCNZxbrg0N5szJD+2p+1rahOyghVavwfuUPfQSmN1fzRYpAj1lnfaUpCYxj1Mz47AZDM0LzoS
m0gAl91GsqtJygoQdPnH5gOaXAAtbE5H1ddTq/EV+u65Kx6sIMF2X2LLx4idlRxkEm6DHnxy4KaF
2xTlM7YoP5McZOkpmDe5Hxa1FsocxzkC0fNZHiitgW0HuJF0VIvNJ8QsmNunca6BgGqU1dWAnAoj
cQpZoeP15pHaGG/F1Zk8mpkGM0vVdy+XSTgcfZ7qo3dVdsuOTHGMxGOdEotllMGdLmpDnsOlLU1w
ghNKE/AmCcyz5juhwB/rENRhVbYXp+ZULmooGYw4oVkScxRbzaKdgVwKS6EJHKSoIvyvm7dfgiNH
5iTlznrr/n3uWi8mY3A6MREcbJgRz14d3IwFk849HVRbekqPZgjVon1IjI0hiYmMzKwF6EUyermt
h79Cmz2JqovqJKWE3oeGIC8TM8iuv/uwKBysuf8I2NgiNW+0wpbfLRBtvQpbDOz3QtKeFh5HddDA
yRd0Nr6rNfFcBVkjXbppc1yRSpmB24dtP0kOrTpWKu8uGnPZDalyeXvKJcDkFlC8D5oMBJDY0aFE
8ZNZHxe3+TkbscI4X/rmbtaj5xUdbiKxHlh0xzSxCDwFfpRkZzMqxrr1pUunPPSq6rVMt2e+LzqG
s6KtNGJ/aR2cMEYIk0ELJXfNRc4qdvIXEmbq41JpwiMZc0ysICqiho7OXbsI5jlP5fci4IS7D86e
mzqa4F8oou7J4pfSRnudM9nt223JQ6spXyhCbJ7bwWByjYYYIsmQsUJigSNzR72VNdCeCoFDMaCS
LTpRhKY54w3MgvW6yRsqb37xjgdcUH+aUmNp22AZMP6GoUwgI4uBykfacYV+0axuu7pEH2Za9l2v
NUn1lH6UOfmbHJ8YBxrbSEs2GxfH+NCxS8H4I03EOO/wPRCD7KEFkn56u4TQdRDN39ZEmkQFrcUD
dnIjFI21dexobA0INowczcde5BUjFljLAvwgN9tiEP79A9V3DhHLrtZslBHCp8sAVnAA2OqAOGSh
ihp2DYO+wQXKdfCR04P6JkYJuzLEg9zAoQ2A2h+x94mEeicJd9BuvgbXZ5ukF7I78XDUg7NjUrZh
UHY5OOCxv+mkMgef+g4h4vkUxQo3K4fCmAaF181NZpCv/aJ9H/bALUDpCbl8+8QZn3nUp0xFc5w7
gcSdG20scvtXIIN/30qGYQMabluVMyJ74IFfDjx/XNTavBv9mINCkafC034Mo1jfARf15l2X0fp3
WLW2Jvz4CfkB5NevlC5a7qtTYzVnUbA1Lm7kuiZcWb60J/2MNWmcbhXUjN2mjWBSzMOJhRF/htGq
oLccKYudqltdFL35mDJxlt8Mko/3aQDv6gNvjA6Mi1KgS0CHO2fWymCSqE8DcIngHy0+38a7so3q
rZIYeqq3i+q7DmPqtr04hnetoBs8cDDVPUC7k3odOzY5Z/lteubDpiRioPxIxqfncCERDBG1fNxn
mZFDPW9r+K7xuKMN6sWnspftcUF3HXd1Ax06eYGZySnykEOb22hhsRJc9skq+PKzaq+h/OZ7zQkq
+MCDN3kFE9gU9N6mwdP9vbpT1R3vC62ak9gwiye9tRLdFvV2txyxOBy8xrdWI1IJ1SVCvuMydrC3
bKYhwZ8DnMqAfAbexAe2DlweXfJyS1Dh6I0BnErj7RzNUBzUSd1LWDGRXZzgmLALTYMJQi6d3YJz
U76bebY/6FeWvhdjIdllUKvErT4Te+WK3jIPsxTequ8WFwMyl04JZO6WpWbmW7R/Xq5umqvijLa2
LYgEKB24pVkjVm39Tqz4PvLQ1XKNR8Om7PJ4b3ZA+lGQnO5pJ1TeVZ1FDCnDte65l3VtJsPw5j4Y
cFU2eHTct8QLdxQq4aTWy9yNyUfqd7C4lNfIQCaycRYUZ90n33kxQhbrpGR4GjNo6YGyKBe9reCm
IQ7h7iQriWu4Ckg8ndDQ1rL82yQCJR2puxZkPCZMHT17+of4v/OwluHY8cZ9sdj3Oj0sb2QaGIrU
fS1/DSjnmtqBKg39m6YS1OxRxLIK/fAEKSC7LjeuzxFzca2q+uBBUQ7v4XJcBRRqwMIcLYF68D/n
brBN/FtNqeFQlZNfUKePojQpx3O4hR10FV5RJM6uSt50gRc1hAtR255VIUAAplbsULhKCVd/nMdH
YHK6LYUUzbEOi0Ad69c+MQOfpXb3phkFiNt4tGcZM7rWALz7BJk77d5PbX8ZIgDOpvgGdXZXcOUI
gOE0TFKbp5bC2UP6AagSwBBb7ZOJr586tpAjp5oqrvV9qD45h7PotwZAeEup4hRl0nRD/y4aDgyT
/Nx8beFXOZM9i/rR2u1bbu844N/yvTvnH+nUcLrmvspsXFBa5p/775jDHtS87a63X5V7/5UsNKp/
13JEG5X7aWTLGf40XMV/4WMo/K+MVAZpMY/iewNjJmN9JO8SYBbdtHXWXMzwMtZwFAgRjdaplS6P
j+tJR9YUROZUAYDd4xSehUxRmvtCZ7NQwtcQbKEqmJwT7OyJf1EjzbZygWcX2kgV2FYIfyS5YERf
R2EXL54trnxoh9B6/2POsLlildfAEBCBvMUjX26IjdgO1BtEpBrP1kEk3Kgjc6NFM4w3Vr/rjTK6
KV5adI6IsSr1dSeUqVmNME9ql+mfVUIFQLeDd1nCaDljUNdoEsYHlpUlLuYdvIcoiGNIcxalOzUS
CjgVG2HxZslcCdB9LKAa59xN26hb7u5EVNHZ6/uQCJ9pH5QpUy37EeryEmfygJCEeFFv/Dh5rlnI
riM/I8DBnPXNjsSrc5ncphHThCoTXDbQejlSjK7B7QbeXqfy0SkgQgPHUtVZSkBjRVLMC5H4rTdS
to5leXQKoZb7P/Ba7flrzlFINBDqpeOPRKxVF4OISpg9HqLwmI6Q1Q5Hf9gw/bgm9mGPUVNCB1Qf
LhYPJMrnoSXT1fauuqzibafz0SU3DsiUztebp1b7br2vi+QP75KqEV5k2astJ2gVTj8ZVsy1ngv1
Bhr9OCixEgsMPaFrtbyiFFGNhRC5OwFhzwWLqZIrqt1c9ZrKca5Dn6mLcocmvor6iyqszBKoYYbK
k0B1D1rm0mW5IhSPfknL3YXLOqJ8EE+5yNzeLFHFmCM96ivAfWo271gHBpi/01XtwB5T66TLcECw
E48pr7Uf2gQFwNt8e2Kxw8cUQHo4/4yfFHqDBqOh7X9wWOxhmC/HSwX5LYmQVF7efoYWPyIkcoAm
Kj67+XNeGMLwsD6bw/AHC3Y0Gz8qBQ8xS7+ujiyO380WwzdEj2+xcRnYD9IphePDUI3D3NgSpmr0
yCDYLSpGrIzLiHzCaItN6dAAvD6BfXgd1jxpMrJtfS2w2Orr3qQhvB8MIDhoTPRpXHpE3NWMwYqE
3aiKVJq/VDyTg0JzwFTU4FMO8l513XRDYhjM6y4OqSrwZZdDeynwxYvlFXUFhkBZGgHYwEeOZlJf
Cgygky0KDnybBXs/H7KKMbvo3Vrwfoz2kDlgttMSmlkLi1OJwerCDBd9uga6y8c6TxVAG1+uUknk
+t1cEzONEcG9/mZVpLhusIvjKInwo8/oZVbgOMOz8Y5ZkpRyME2FeamRFf8l7yZCARDcrKFpDpR+
HOqseByo0a/DBe7XNvkUofQfsMjSc4BJv+NNb6LNkXIVwYv/GBlwt1eoZxX5KU/ic7Jkcnm1AbgB
oU4+GQMYnx1jSi40gquBZ/uOnd2/D5vz8RjD5cKgM7PR9LIN9QdaGD9gSH87imZYig05O8fIiUBK
nN/Cp6oEXF1uyISNBQOwfjOkz3kL3AhieGzwEgarzaupVhy8W4pOnzlPKZ+r+uS8wpMx/iYhE1lL
joQF1rlWZiG1w3AMDv6UwGQ+59TxzPfpuXPms+Gzrm1VpCRf3xEPvcQrugwK3Xx72lSnWoJnjzOb
3aFupsen1/s+206CtclLmAzfy5dViPPmDhkw4oXGX2kZYxC+Mv4dt1qy8Kq4D7ift89QPLvC9wNk
GEs0GQnUxYYWy4ZAWeGAqnPUG6P6RpAh8mbwgJJLsXz+wu0m956saOqI6PtF47eB4Q03X5rjNjtY
GY1Wso7hqbjXPT6N6eHtkGPk7bAZs11/Puw857t0cPfwDulh4IKl7LFZj8Q73/nIuc4hGKk02XJg
I67MXKVPoe6tT5RoztPfp+YAszupUC9X7AOQVx6OnSkk+CMbOi+vW6mxmv2s1tRr0CxujO5/mlZ/
sKk7c/FlxZP6FJWX4i/uriqHqPTtHTKR3C2FMZ/wbciKpylsC2qBG7IXJGwRthjhwIQLjNGPdome
aYfbHtDY0pvYfWn05H7NFKbAXdqKxKvFiUNAmpA/Rh+DGiwcpJm3UCT+1ODnNed9Zb0c0ozFN+a1
HXiZS3OKKlkqIDcZxXesiqYn+kvvGDH+gMo4bwcn/eD6uZEyANRiRENhZnnc0228xnP4Iw5Y8AZO
3T/X9glnnsUWOjm+XcJ044ZglbTUV5oCFA7BsEJI84ABlN8S8//W7y938Z/3FGiJg3izKS7NkbJD
VBMIlBt+TVyg6q22rkXb5WBDyK3V1Fg1Bz1ViNlkGNOx4DF16nfXwyxWENfB+79SN1sssuqC2x+I
EDuiD+KBa1U5aBeuVQ+azKNr+qKLKarubLaCcmt/6uFUQgq0OaKIpw0WmN93wgvOvSZ4asF40LKw
EXV8sKRu+Zp75vPvMoN2FJBsp09GbOoR1VShzLtPh2zHp+E4MeVxPt8WnlZnXPpWMR+02zCHEeTr
srwSR4xrhwDms38/N9+o09PIQLgKo4lcaXp0tta1W0HTRUVmorpQWmla6gJSrsFIMnFqcB/faAkf
XGFwmpwvOUZgH7j0uaLXYtEh15LHXM7Rq2K6GPOyKY/HlZvTTpJupXtGWyARjX8go1p7Vh7pzfNi
pbXW+MFut/M+B9nQn3Z77q1WSl3McfLe59Vcnc0/g/vKuD9nbSoIH3q+pBsBdfwTWQ1UnWnMMt6E
W7NhhXJz4UqcM8utvPgYQrK4qXfgokdpWsL7rXQPglE3q+Yjy3m0dBJPaqThleXzjwcAtI77lEID
fol0xmAmeZUEzp0ORQW1VHxC4o5G3tB+WOcP3yk9/w3/X2z/UluI1JXur//SYMtlK2I9sTMU+x+l
dQE3RPH2nLVYPFsLQfFD+synakLkoKumTPEP8W9wLTw1PklvjvVUG1e43fiOM84mcIcQ/zYIdyo2
/w0+d9zEkKhzgt79z7PcduUvAc2kO2wQDbG4Y3QtqGojxJuvfpzQp+Vshkss0MPPoGDJ2T3ufGdF
cXhTNZ/cviVZS2RmIQ0KhudKe/FYKy19rAMwiMcUDiVO4YquI9H+sa9TVNcvfUrW0zhgSSYz8zYg
y1SMldjWUqF28GgzNIi/zpsJT0tsCFLLjgazVNCK9rUMPro5nvxaSI49YgXDPd8VaYw14q8vfxRn
nvOsXZrwYTRs4++aJYY2z1i8NGPGBzt7iPMvW2H+9B6PGVodcckz+FERSohX3iW0AxI8TfeozGiA
0B5XwXRyV1VZeT5NlQmBROrHlGPgFB8DvYLlJyTaLH4NzqVCngk+/t/SYS1l3+/pr3MPu0reTec/
txzfDo4CeYYlLNNU9HQWAzLfTaPLYGtoTiZm/Hd7msjnPymX0DxHyqYCY/sGyFWQYKbcBIEj7uRW
Kle3syu40LgGRtr499wP7UincBEa5TNfmmcn51VoDAB370DAV7Dr0QgPGXgotrju4Ud5H1hZVu8N
7wMW5ujnUR2FGRqm/Rqrk4/4GLzepvcE360Qron25V692U5rGXKZpHtc9qe4TwYZMDc6Ovslm4yf
EvzczZ+OP9jPovmoPaRyfIjQRWytTvb8a649/68IUcAt/hERMhMdgOpIej4mSLZECd3i41uCTCTn
Jk0bdRgqiyHzukVy5ZPS7u2TM3NrU/6SAcwGtANc38SWYUP1IRWsSt2IBwW0JXKiOzkEpo+so6ye
J3ViHrcTe3UWRxyd3yIn6puv1VMDZ3f/a1iAFwbS8BMsRSpB6FWAfWrMe8zIz+LMIIHWZ3ZnqFRn
v2QRpSudPWPflsqtvizcyyx/MFuB0PQTmJ/MZcQrUWKoZpl9mhtw4CpNBZjoG31SLFfyq1oi2Xhr
m3RT1IoDPAVhtMAYLzpkiLHWVLLUubWwJz3yxy/SVl0WyO0VpW2aLQKQFG4fIRbvTqOfBFk1rsSC
HoaW+evXj4hPhtqwS2UKnS1DDbVIcAq01yUl1iwYASMwC+4fHgqdJzJn3tryi1occqthwb4ETOeW
0pNLXpbKu/4MTHBqlfDwMo4A03BqS+RQnr+J5zL7Zj27qFOuMlfs4oy63ae54VQKHxHUdhr7no8J
XNzGHLrfui23Bv1Ukk69ikDB29KRZtSL3ZRARpZbBTaTSTe/I8EgxWOrI3L0eYD1zBqIsFyCqbpd
DWL0i5mcm7QF6dH6TiJP0XH9c3YdyZY0t1hb5FxB4wfx7ek01+TfpVhAbBILojZhf06zoIIPiahN
Vf5bG+cLuaTcJVKX0saqT6NGgTOaGOVsTPzKfffBYH9/Au0BnToaq9cMHKPj2kOb/mTfRqKiQ7Sr
2SZ+pBO0bJI8on0olTmuORgJUzDXAiKcRbs/LNgFsyOvQ5TAKmoDwJYkzN4hc8HiTDSEdF/hJ/0C
+UE5mBRkD+ECVrhchBAeA2HX5sFjcOv7ezyJvR7CtIpLHkqcYPVVcrOgCI8VkBkeBoCBzxzbhZmK
TCzjPzIUchcNdayFxhJz2b3sskJBxeZayrVhvSAVZvXvjY8huNw+eaMJDUq7BdcDfRGi7+133wly
YJZGQXBlPyTNj+5VyKOcUYtRasYzfZ/QXGkHGRjmsMk97HMnxlwSDC+A+7wwpo52YpbQ6pihHtGm
xJVhR3O6CfwOnC+zmccZCww68vWLpbYGllqAEO3SpnpMAQhZcUBoxpZI53uG3Oy7DuFtlajQuUGu
LmYHJ1c+a01xeZSxh0kkJcI9XMroQQegsI/vNQFQEukOMeO8J1t3WdpNTJdH5m4N9fgWNr7zWmRA
+5lgLPJ3GHYH41I7n3MeiBsrvKruIfhvTS3hbRgnW+/tP5BNArGUCpNiRDyj0bDr44gR9ep8MGA2
siziQ3jqzAwxyez6y3kv5+CnxQTxiFIkTur0RxSo2HtVeAnw4UT2ouCGidnaIDzbzXM8MxZa2/Pc
JmKadfvulA8LLjZlCPT9kCH991ej+ERd4LTuwTtRlzWqdZfnqpiNl5JmiOvqPyC1rRnMMC58eUEx
0ueWmvFUyu71QQ/WPIewVxECwx33rj0oIKAGG0pqJUpsz4ngcu1Dm5x2HBdB2ceBufxRXPhH1xNn
0VGhD3goRgyII/IG/3vSBAuHjAnWofFE5W9lUkmp01XKrndq+uaGS3rs65Ke51rtK6gGplgX/ou1
K0Gb8RtpIN8i/xvA+2cH8Bl9aKR6oP+y5WXxhrGrLa5S4zuAyqNGyOYZkTxtDIfIqE8qf7efID/H
/4n/dWO5ZGgk5Pi6Mf7BdqBSeMNrqj0F3y7dEn7b7ZhREsljF3GN1/jPhM/SJhN5b86l07SG8h1m
todRwPlIVsxXiqJ/WogZlWkoDIsjy41LjKdH4FZIGDCCPQmplUlnlPJr09uzB1UVFBR429aPEOuP
4OIgIJ354N4QWb0wEIPseRyfpUwVNvYprkcoqRuVz6yWRGzDVcIFGyb8tgT1jV30aDAJOACkhbxw
x2E444UaJbBXs7lzKkNv3sAb16jv1yemwrp0ee5bfYG7rGFpYQcKrCskGr3YpYfFFbeUF7svrCtw
iTBax6qD1JycRzmAyh5c81Tc1mh870jtzUyPH2dmrKwOF+NfW0+phES2f/Z2BQ0PppgGvHedFAa3
tv+JkEOT79dVioY9uyQME6LzUJpUq+uPI+QuRnL0n0DCVnjHJXF2sHgEbVSZjAIvQlC7cEkuyWs0
9z1XET4grnMQjmt06mqe0Wk0AjAm/PjJiCmEgdc37JYNTgxw42V/2tqriTT8xbCYMuxlbngITObB
Dmgs3lbVSyOmSPwSVSLQ0xhwMkSzlzIRD9m1MLq0jiUNzDEcWVP4JL7Hb5jMb55VSpMhiKijf6fl
MJ7uHSFW3Lm/jAkcw8MR8PPBJBfc2ZZMkPcYq9mM2SKhiXcnb3AbTGX7nhTIOkIYosFdD6fofsR6
IH2ZcScDDIyyhTYbRXjvV61RTOEe3HRvMfLEvl5kLTHOttt/MOfB5/n7emHu+dYgYpaIJx59Dm2f
nEVsT697YUxKHIgsjLDSq9Y3HaWAisE1jb0DbioN29wm0oWrH53qx4TvoGCeiqQUSHNJsebZ3zPh
DkY2QWllmNcmK4b7B1Eut9BCTHSSPpwE2CyltxB35BTKUnL+ImiEL3try7/jQ+M8UDCYKlshNorP
rPTWgPe2v0JoqY3VUzSdtxq4qBHSJO3Otf5HBXO2i1o2+AVTZEma61Hq54wTqev7ELPfOrwPI+4E
QQCZ27zj18+us2iJWbBs2xjme1TCXekY6nIKciCYWXPxcqIVrPQSxSlfRq3ww1UDySpodxIIOM+k
Gwo7sREgeAsXKereiWlrtc6GhoxSlIFIEWp7NE4m/PAMEl40tfABhpxqkfJ3lvK+cuvqGnMl6HYL
6XtbFqmfYUs8b2II3LBIx+VagxbuAf3XugUEqNOk1Fm1OS4+MCl3BZMDdbXS8LPZLGd2HFhvlMsE
P/PKnLVJIxnu88VVF8AuOQqt6sm+xSE+fbUs7HFGDLz6J8veGOgxnMPuVxjSUBlKMIgUinP7qsNp
bzWCVGOrjiOatOa8mWh6qkauJ1qwQPDRisqo6CNK2RHxrx+nVlk/xRUUZrvAjoTX9X0XVvS7z8xT
6Rq28FAL0YjPdnTqMsTanNuMN1NI7xdtpFHrsBFIFPUk5A1VyWkrKuqVlejNOUia7pMGMfD9zAC7
0WlyhMsIj2LoyRvk7gYdHBS5g7nLrx7jHhQ1fpLevjCLhp46LEhzW4PWfUV0shoYoMoJKE/66UNh
yOwigdSQGLDtanA+T7fJwQAmoFlzH6AQgnZoJj7OrAc5PdvUJY81c6WAmSL8aCT5+v5T6v8lGWby
0F6mJ4H9tezj+/ULwpoCVII+XCeCp2MCgCnRao5bWwzuMU86souH0DNnqyHHvJOAd8b+nrvPv7QQ
jAhQ0CbyU0lLU/HpcvxjuIG4vg89vYC5OJGOQM0S3mDpOynBXkUY0gKxvctTQWMfwsgl2VE5ynOp
iTD7gi0ObnSj4Fdbza+4hlZtkiHE2Nd89yam2iNwGW8j1cc+bjNKT7WAt0fT+fA8IfaEvAYwIqVC
+hlxw24CqA3lxWVXwB1pfnWk9WmS/juC57spfqSPvu5uipMTmT9wRvYvWVhL4Z5py8n/0xlDYVi4
xpfMuGGJTAngP/ZHEMmzL5RlaScv78dYj5h+W6wp1B96CQjL1nER9XBfCdcrogBO1sGNasnJXTFp
fpVx/lEYPMV5+sD0SiAlYXo50SwDlFjYAufDiyk/Cy83KJh/1C9/lihi5u1jdDt/I08wzk39TcYT
buJHah94iI30IJAXiF8KrMiacbsKjqJ9Dc0N9Uw54KxxS3lNFJKd7z8nPnt8BjdmfDwr4qMBI+7c
hWJEbbtkbWTNTEqZq3a6O+KK/bUwQreDEHpGSP8g78JT/Ofaqwljpg4HIe0ZnHjw/38mgt2y8i2r
JMEo18DF1pKBwYVIyOl5DTwcUFxO2rsUFnGA6X8X0lx7JqHyV+lJLISUaYMllVxjcnh0TaBSoFyl
1Ur4GvLJ0lySIXv9Xd9GxnHoxBFrItUhW0hKVlv4KR7KR3i6n/eMNYwPuhlV9DuQBdPVdrER1ve5
BxJCkx/U51f7RhNQuquaZzeX064KMfWx9HdrQOO70goYgEfpfLzp5e0eTFkxLRMihmCz/auvqCOV
RrR0LQAEaQ6OQ9FBE2p4FkhqWULwGXIjqNeAtkYHNy9aOjvgVa2AkOtNKLXndrBQtMbqEDP4xC2c
+Q4U6K2UHnlDn7h54i6N1wPaENVYft5UMpFZNzykMRysMDOgBy6JhlotUdGqQ6jJ8wecN0dIAHBJ
12Hl6ADSyTmV/9vGgdRj7oMRbrzEbhADlFI6dVdfwYoYnYLtEiqPm2SK/Ni9UNIiys3X1B2I+NGk
xQGZYmYCMoBUyfXUOiJ05wBy7fw6U3351ONaBk+ptfNb771nbDWJP8Y+RZ+fdMz4cWFiMe4veKun
BU8Aru0X+JFjw6zALmPfqpQoigy9zZu5nHSJ6bctkWet5AN2gDBI9J3nVFXtTH+JSKMeHu3RZo10
Kx15XfjziyquUL2OHzIkggmJFJlcsYTFEUPtzz4sXozbEzn6fQsta865DSrR9GBCs1rF+lyd3iws
Phle4YP7tWOVAKQQD1jcKFhqIBkp7242auHhpmFNLUsQEyS0nDJch4/FFFeaVOIOxTqC/Rx6XSPM
ZMGLvcWqwsZDokxIfraUsnu/owoJFIsk4EqdW8hIKAIroOUopcTUDgZqK4+G9pUrv1Dnjg0TS7po
75jp0XCdyrocSklVxTQac3PJPtyHO3uWkM75eSeNvP9D0tjelWtdJ9RsLn/AnafpFIFQJh+mSw9d
MrtL3S3t9AuKTPWoOFeuab+vEE2W4HTnZW3wr/BlfTe226dxtP9sUcI22jLcS363IS2tVtiP9gl2
zrreCpArtNICXUKiEnJvo8Os3S84rpFxt2yZQKMCA2XW8EvmGrYaZcsVzRPBOXPSQ42Zv/N57Bgq
jbwhnrPCFp9U4CRmuUus2AQSPSc+85gskN6rgBcliHxBrgS7dQOzZO7oKYpC7Ics5z5XwXpIIf30
WjTtjWca3ChtU5Ij2rknxwn2BRtpKwFEpMl59UcqggR3R1glh6uAWi4bJQZ+/R52Mw37Bof+UIeZ
5putDWVqx4Ma/Q0ycAUJzolw3XUyI/3DqI88TcW7ktfNBo+lb+3Doa3Orug/rf82i+NnOnApEme3
fXXuohEHr3TDvQvod+MGig0ujw7N/bDnuc/tcW1I4jVULAzDCFiSmP725GT3PL967+k/Rdnlssnb
V74Z4ABx35GHFks4o0fA5s4gbsIeKLiRDtJ8WSoJXmkHVNK3b4Jhp9fWzGxDr1VGHq4O9q75eL+0
A+k21VvevkGUJyN4dn2BUYPU3oy5xhrHhHRI2UKaLLBjiyj73oCrnxgm7QiGsRQbvr1KXzzs+ssW
mZpFybMGnYLAvTnoGFdoE+u2drzfWHbv6ZpIzy8oNq039kzX/dfCecty/b1LdwKcQmS+FPzKUCCL
3wyvsNR34ehFWvvpHsw4PPPP2Pz2NNVjlEQV7aEOqQB2fQvH7lXiJZF9BCdCFrsqpSkL57TbfM9Q
ULiJyNMce5kC+0d+0yjLeEhfxqz30gWVD6x8iLjeyaamv6B9YIS8gkBkFekKEI2JPX3cghztVyuJ
5pxIe3nhCZiCb+pgsBAm3jtrA7zob32WbLC8cWBdqwM5TdnEYGXhleFZLSrYPmQrF/h23+yZfJK9
ETyROHAoCbg82pnuZU43BRzi5a1RBN8nHBUqwVeW3GhHS4b20Or+tXe13a8DHk/URSSVgtjyBb6Y
kkfzmNgPVVZ8f8IDXGbz2DyQh2rzej8JYLUN/EwDbNSkKxnQvGDyqFDtPqkcL5NvlutEKqN94kNA
6I1qv5VOaN70LQim/tsS4MfobncSkz60LvvmpGN3ynLXImuUrmK5Hu9CLi2Di5WdvKK6rmm6glFU
pAlyXbknRHKSvUI5XQ1JLrFcVTyb0AXJetJ3aSAh3IeUKrLjgU1ZeiLhVwI1refs07Gz6jpDFEGG
CVmbsCJbJ1JIjmYyE/KEU2u1Ku856kl+mJjRldpKwBkngz9DmqfoT5VbhMkDGBknB5KWk6sniG2M
rJQYihbJYdPLNaqJp3wh1QGH1fgq+Jb7sCUvBQWd++edgU+YsfZ+8Z4sxo2N8butjEp/yMW65579
BREK48XzzwGQhjSOmsljqmqDsq+4fowWgngmibAKjSX3WcZ4HC0mnjJzEuiNhQlg1iiKS52gjIgH
NaOZ4YdzpzQRPwOXcsqU8CvwfYCpyqj/paoAFCq3f2245D43I5I4J4YGSFSQwemXMLh7F+k0Ki1a
VRKfsQ8S1yrigTCKryTcftJmERjKGgsVp2xZ7upBRGDRzzNy+XxQN4pPVmRhgUAPBJwU9Vcm95kd
YCFHWL2u0h7v9i4zKASr3H1eH2NijLm12yhfhOkNxDBHccVyw0FYTxvJlDi2egtwN6InRvahUMdD
X7KIt10yNm5wZQQJUoA3bdy1goS5w8nMZwMvx3kFVczbOtVNhkZgPldgQ/WcXMtlDq5N23lsnjPE
xmzd7Nc5WdHm04xKMBkm4oqpYooQ/3E72wFZe0J4W+yV92tfAASC89tDEFhv6ojlCHyhmRw1RJrA
3NZXo9B2fDiv3FQ09Gbc+6g6degXrWgFwCqJ5pxCWkqdI3zWmsg2KoC2TCjjiUk8Bkg56iLxiM04
XTNJL31vHo3g1aYNDZ03iCfm8OWn+FZDsNq99RIf3vZ1R5vfZmubZ3jS6NUQEaiJJl+a5E/6iAf/
nRiNZjfiy7P7mjIeuJxZzXoG/VYn3X5lwExiSL4bNGA3TlwnTxJzy0pkrYAVWqRWMLC7BE+2/RaI
mdOi/Ux1pHEF9lh3B7Nqi7F0PdljujvRlqlf3Mv4w7Q1aGgoYR1gU211MUalIKpkEwPUSBL1WXCU
C4bz3xo2BhtjJkVxFIhL0ZlN1lb6zBxxrBO+w6ii8NYI8Oez3ubFoPgXXWelYhJ1iLJHPH7fLZDp
vSBr6ndJbRb4DER8ilbViE8CaWrO3As4g79iaL2kZXQqQz4JByG68yQGT3wN7J9ZYeib9gAGv4lp
jnONtftJ8WAf2rvhWYqYbO3mBERZeSXpWM60GEo5dsY/MRHjhBRlUvae8DIOvwgXTNNYqqZQ/qWF
7x3SdWUqThdLq1ctucLrFPKd2P6wdhdEWeJcJeg9TxyDpkwpgFVmdOtjmg3gxwRCaw4XYwJjKewm
4QHgssuMIMqFfMeCLiSehdGWtlJQM2vPTVNLhKPCpWYt9nioa0yCaxCRhOLdBTkuFWjNM3zruef/
nHjEtxTPlJcoNdrc6TYDe6BtKSvvYuzMhMek1PNB0OHbUV1NKKOM49+1a7TLqiJSYhU+MgCW6mlP
F26Zj+BzHA9gZYx8kSv5cd9ewXlSDLfb/bPXmgs+vQ9++NZfforMHSVXDBRuZW0ZDIVpsgdCy6C2
PoM87cHjmyq31PJWHJR02xPc15bGQWto1GxkIvsCojlurXS3Jk/nDmMXHZyrBwVEQWXu6HnUyde7
/kBX1q+WZ+daGDVjwjRP9cd0+6TMv+KneEUN1+ynTK8Qlp7jZNGr08MjVVdhuZhqvxWQS7T4ZVhb
1e94s4qt6KAGoUftc3PTJV2M6gQO9oiVqgOofNBbFkbqHBEHzurqzOS1KIyF35f6EzFJwxYcPfT4
O4FMK/PMaDkDzDwhKskA5f6PuiMn4OY6Lc5Tajf23SiFjrRYvYxNxPlwIQsSRYIFI8gdkkEk2FiF
WyKXcV+sQEtC+2HNAxeXYgJUdcTUQugSY7o90n3GO0MDF15wQbNsUD1BRiIROzHnIMmjcjcjkjjE
uE5yZQtDJJaXj2xKJji0uXiTj9aOaZSOytDgpZAEruJZAomXEe55rE4aJ3zTPPa8UuLpVeF6mWQ+
fptcT4POzNVRo5+xOHqEV28GFcQRLGgi3JVm0408T4VJ34vXDTNUEHA4vemhYOYQPFGndnhuOcN8
y/o1aiWEklbpLZWomdj3262MZZMzHeDc3p/lkqHxdbuGZEd6ySWlVAki0lTYDA+Ksj5PEMxEVtFF
AI8Kithkmk1RmDDrRpwi26VPFqWvlTknzSeItsobKN1xj1HWoNxBgnvzLEiEukRE272j28Sq7C/5
3R3K+8knBtBVeXK1RmEenu8BztLziKOOfbuodh+xFOI54CF0dDgWAAuF/V6bao2iGqqW4uFSiPgZ
fZLAX95Km8sIXtl8LHIKLJBpCauFPFp/RIkPq/IFHEcWZ3pAoPUG1OWJyA1cWj1P2qX4csXLgU82
8+tDbn8lSlgBPr3UMqi1QJRbH3Y92kMa6x9/qgpsdRrQDlslW3GFtH2kq8uGFOmUM6ujXekDZIG4
Kk9QzWhjx7S0oiudVaAsQ9NxWZKdFhT0RfLIOiC3k1oEQr/Q81wLVqIM2XT5Z5Ey+K9a3MOjOSjO
fjCHS/YNN2S5OxAfh0idindOV+vJlEk6uemDplFnDWT+nrEKaGjrtaMFx/q36c+OAjur2D+DAIYg
2BJEuEQ6y0QTpSxsGt1WaJFZaVkwTxAiI6X3PVHgDzDzIOfMfXb/vqsov8w/TMTjBOzJX+gdDmtn
DkjubwdXNakqAcYBPpQzaFs072ECvRza57jL3gSBtMokKnkz/CKYkyWaX+ELa1TSIz5DZXu8sZfJ
1fbQ1P/KCkiK0mWLfZ9ltJgc6NsXj7E2GZjOMG9eqXhEGxjGozEot4QRtZ7XA2rWnrt++ngj3YVQ
WQpxHkBd9+h4p7MurPrBEK1yWFGt948asUeYEVuoOYeDrUXOJepbl+hQYAOHZCRUTSarrMZpE6XI
mhGgOUVxZdGe7hqR5NvJS6Z6tjqHKky2e60kOzNgUd5pDpEox2stYy+AgArDv5YI3gTb6SIVs16F
Af2qDcw0rsudosdLo27DDNYLUOw/TuX89fm+EuV3jWYiYRfE69DJhqkKeFaRSm0sTkbpLgRXoKM/
k5Xln6KE5uTTRarMjog06u396TpqGqWJQtDrUum8/vT2fb3UsfufPw2w6QcCLJU9q/PVes177HN/
H51dPsU/LQWX8ckEpsMInKXZMnwZZ5CtRSUHI4nX2e138DxLozFnVRLrsUTo/SuOCoMxDh7eiC0V
8L31oWYORhpzLwsWrERg8HZLeC/89J0EKC8Zd8FE6MymZrsBl3gWnCRZIj9SwjS7hMkKcCMn8nsX
Lg/n/DuVlWFDV939abXdHjm1Hs7+ZYJT/wIZ1v81QqWXXw5eQ/hE/WoeDdjEgTNPEw7S3DksjYt9
qpz7fcaYmiWFL4Vt/NFcfvdvCzCyYdBF57v7xxmFNXqXoG/fglvmjz9EL0liU5FD+5wKVrFEM2F3
F3Uh6zaiJrYkyimDYzSyQgkll/9DdXWmGh46n0KkH2giVviBcHNw9JyZ6e/GwJfiLuS1j5f1cqFA
cMB5uUpsvbyVfXoNRgMEDem+gVQjsMN+4rjeLgptJmqJf1iTYZlVweMzNAvvZ8o5+mSRmnxcPrmJ
jte01qibVL4NwVZwYuKZD4RTvzXK859R7+CNOM333/GlGeXkId3bOVbT2MnN1O9GRFgYi2gZ2b68
E9Q0cOjnU5Jfyv55oI2IEQLfRLZO3OzQIiYFVERUv2m/2pA4v7AQrNDd2IbTCpZmYOJBymZUFkf8
YpasmZrWRDdVS6r2m9d9tAqjFlpZ7bwCSkixD5iE9zrMxyA/yRpY+SyPlKBwc/Zz/yhb7ADinTQ2
GoplvYClMLnzKL9Mp55d8U1G0SpX3wcYxvT0YPQMp66Jouh9+Lj8d0RGmOF+7XZpUZdiKRz3LQ/1
OFjfAjgT5yFRA28BfdLsO2fqXmHf27R27+ZIKj9bTtZqgRR3U2AQOKeLhA02d0HkYfRxXhxF4PCu
pdfnqY5TEHyZqbRf4eMpflFZcsnoO3OPaCvhU8CdhkAxDoWZ25xof2JDBaHknKZFtwHz8ziejGLT
gFifzdplQz+MXBfwxoQe4n7P000zgBhAYFQJk5dh5ew+f3c89oKyFtWgbBNt17Xc5TKQyy0H7809
nwEJmliru3WZC5Cp1klRxr/egxt9/GxhbYq7kPYllMzMHpqd9cVtGfQbAIOP6+EWJZxHh2Ufsjug
6hJI40ShJAF+46JBSjywwvdQuH3w2h/Ck1nQcOl4qZ9RKEqakf4zg0lQBw4FZw6MRsN173H08I0h
NRp2JmUec3ycKzfsw6hnE2piAYiPGlqQrxU21+cjLHqpmHJLbjLKieOMFZ3Lod36x1K4+ef9dv+P
rA+BIo0rZhULKBk7zJnBgj+Y6r4gvUI0fmSR2iGfuTYXj5iUom1P4EL6yFFnpuFQXQcIi6C6nucK
dTObKw55qascps5RRXOBY3GzZvlxW+bYWcHne/wiHfGjudwYdgSswgmO1aFWs9Iqnm30ZLRk88dw
ea4utEO4GXrtiwRppHv1eYreaOxaoHcR7E8fooRVgaj/iJugt5t2ijg0XQgs3P5BkUMA9GtxrSlg
aojakTe6YbI1bvofZsw0SWulqTtr1hPOO9fyJA97Q3BNDLzwGanJH12vmo6ShnA1KDgewnpUggHv
x0ZS5q8A/s5Cb+FQF+jq+z+eKi0OzGTtrtKrd6cx82FvtJgTEfAFU9Lxuv50BhBrc1b01Vs/V1dP
1r4McOZTByMerXNiBMowLpKcvSJxOdjYSAmW0SwyhuSQuEhG++3lhdsnl08xao6iTovnIaaW7Ebk
ffdhOlgxGm0JmhjkK2N1KxT3rlIEAL7qs6CYOlnrmltz9ECcNmOIo1KwET+anrnyIPXKkxN3KsDy
POZBjppkVG/NzV1v1KPRBfwuzIrwpyxa0TLJDDVQe8r6kEpurEB77I///gcuiwzMXqSfHsOdcT8q
iFtfbANyKVTQrk9a2p73A8bFE5zGbmvihAWRxLroIYA+WuXeAB/jnB6AHeBnH1MNnLPkV16xWnFv
1Zh0u9NuxCQRPQeC5d10Ips7hXWpB+xVhEzLnuTcJeAFWkVPood5B4Pub5TDUw+Jlce9c/uQTLLe
YZCN4Hgli+NIbFZKtjiWnaKaDuZOa25VQOlYUNoNNp0++mv1Ptv0WegEjyATX1tTVykhwgqDNYUs
SeSxY1LMGwaihwLK1ov9UNkmcEvbT2jnoiCT5mGVOUCcfr59XmyI/JNn7qVtTZMTxupCdriygfIM
PrtOiE1AevIPQgICoYLnbbwbueWsZgyiRM94Kz2egDAorfdftSiEDYcajC3+1DJ45Xlzyi8hvlWo
/Jfkvx9f0pqVXQdzWeEIkdgUR+ZA9WhSFe/qdHcDAzSS4KvTahrMRPxdyVdw9/tOB1x76Oeo+w7+
kI2l5UfzWepyGjNAPO8HZVVcwhLRVRIiWXubhRICc0SrJSoQNQP0cw5rQd/2jhdKnbKTycfODcvO
kauDDKA/uSstW9O4b18vSjDrP7rMJpEc1dGn516SKPbnNaqvod+4iNL9Qy8KrK/DY9EAUxWPX5xN
oEQLWZ/CqMff15L8bDGCiSN7F0/xnXzgoVdAoE1DpsIoTOB0JiRKngHo13qjauvO/aWC0NoaeBCG
r7FYjfcTkA8HVwzyYbKT3RQDcrrmI2F2YGpJHDQUt/zAwW5mjH62pW5uDuL7v6hq0Gmjdz8WPG4K
khcOXWcKUIZ+mmj0g7XddClHMdbBbAr2zhR7PB5jhD7Jy5gbxHujaxjn200CwzjsTA43cO36CmR6
p7lWfTQkGui/vtotmGaSppfA9dJ8LsLYJGMwR7YYbNuFJswXW8fZJDzQv4iD0ONBRSWE6r+xmkz1
p2E4XKSQDmAa1eulIhfBy47mlKPIfqZG4aFxxinqcTCYcRP1M0BSHgxmu4SPZvtNjU1A2M69SKpZ
vw+bz6e6A9QaOMBaKC8WXfoQ2R9CnsblDrlQmb1Q1wCJLFSaJbRORGQXYO09+U1FPQP68HI/wfDW
0Cyhgt30ZJDRSgTsRjkVhqszK5YFVy0IwJriDOv2QL+nisb9Pt0cE75JsjDNYGZ4NtIHgAX0cwoK
M89pviSRSEN5JJGRARV2I4L6EWGOSrTPfzAojT283SARKfzKGWQ9gyogkQSCjEc9rfS1oG52j6kc
WLK/32KecDikOAqzvVopnrlOWaxBxy+pq4dTB/7+2CEBBTkGh+4MRp4dRWY/3pkzlgqLtLlQeZFb
cgM9k29IwetOC5d037suuS2ayacilsEDVNUy8V0P47M9nuY6X4ginogOREipAvpj6YnzxNtG+uOm
WLHXZRvWo94wdmTeZ6mAcRT1xVMvMbyjwsSe/b2gN0JmGGAM6TQxp1PPn9aqsF5a9PKG/I+vIiL/
yseMv12pFxIQW3L4a6EEf6EqnrrBoAjViTjgT3yADg+W3JiROz9sHc454qbCUX6FYJPOH+39tvY1
PjoJLw57OS9ur0g/PAaNAe+88hWnF/aNG9YwkTNMJUj2vlKgpLSzNLPA5FxjMvgS6P9F74NlxfMz
4tinX7QtOJlR3UzhdzK7ipOg78OxDc9lfDZ7XfK6qoK8FS1vaC9qlzwFFsi7o1usW3uyvmnL+UHg
4JHtBBlCAK+3RWOLLWHDCIPbKLDaOBCwdYyfIzPteEUphy6m8iW06tx6gCAUWooPFUiKKP8CZ24M
kHIlWG2Qdh6r/9vvkGswAROWPxLwj7pnbWaJnFnsFPx2gBgGRt2vktFGzLmKleBNcZFPo/4HGmZj
DgSs0WHdPDWwMHEsCxzxP9lGHAl++xIA+WxzqWwPG79d7VHRWRYbyZZv+XZj6ZInnaN/ofbbLA45
hDjPq47ppcDogcIkBp2lpXx+CwoJFkgfE2CfC55stSFjv24CR6TLKImTcGs8xjAtBK+Ho+DvAm66
VzxhLP8w8NWOsaFfNnwH8yPwD5rqFl6WEIYyXFecaAxBdJs079ZQ72oJGODzwunEqbAXq9zyQ+fH
VwXdaZSVU3dgnhiX3ZYZw+jBNrGwVIjXeT7tIj8pREDQYG6SoJLbKTvQhYFG/lMjOVVMMkRzpEGz
2TYfMs6uxrPmwlVJQYSu6/lZ3xxsno9psvNokQ9lwginjeZ54uKcxh4RJev3tUihfMjRQZl2x9Mv
W8IWLtG1muw4L3B1PysdPd+7hiOJpvMx+qvcbHFEvVkH0bJ0NDdNvEHconmLoNPeW11sNO7GRlga
tjNFZmoWYuF79EWL5eOokJentvAIQKVZp7Ly4TcjYfKC+dq2uQ/rjEOH6jEgxbHM2mXJdYjaB+V5
pioSSRliv1KqaVh3JideKIL5CxRgXwLZjdD1n1ZIk1QSrzd3jpZECQtU0uq6yBS5OtgcRw/PwgLk
G87+S8GHO4z1W6g8JS/U2mjN13IDgr2fysGB13tf5t2qlqjUjG2BoyrCoy3miOZFUas67i+CYZSr
DHbaizAKE0diSgx5ecsoHtT6J4GFPGAqCJ0GzoM678wtH2KDyDVevVFC5f9Lnby4fYqGxU9rYVdr
0SBkrlg8PtD3Czp/mP17kiAS0zdhdT7oSGBy5yILgEFfEWUwh0xy7iizuj6Go7YsfICZ8tbzViWI
gx1kN/UmPt/yqasNhJiWIiHT2LOO9oKR5YDGClyj3VGWnqf7ZS9PmILpjCk087R+tyXp7OpM5YGG
yRk6/BQD4rnBMUpzBa+9zb/7SDpyXY5ePOBunfB4Sa0/pdVuBefOsWt3GqA0G7UDz4V+qKpyywqK
bxMIGTiXRxZXOrgv8jzTqLHojhGRALPaN+w0re3VoF36PqvS6N2sHZOEV4Yz3d3D4GMr0Oi3dGj4
oVocKaXpmAvT7tXX6d2Cvo5EYiSP5D2UzHPs6p1CTyH9NXgq+NgylUq1US+2G6957k0pPCfhVh4P
AmDD8RcgLnB+u0emZP0tlFv7UXJpM2FHm7qFClTnB0qfp27+l+kictaUrjdaYciKJyen8ttLikbR
fdq1B9DpfN0Vg1PGkGtEwwoIkChLTBP3PY7wQc/Ml0rXQQK0KpKikUKf07mKYUZSEeVbbH72ekZ3
OpYNNLckEqmj+6ACHqh2RQp3kjHlCNzTMS2bod0uLTcBmMuqQd1zoJUqEjPMKm3itiSiqEuA0/01
YAqPjj2au9bbEVxvz7S9lhSgRqFoZTsC5oyi3QuN9yOfW+jMJlj+hDGICRqtKQAK6GBw7BdAB6E2
GDelJvzQec4ReeNToQmqxEy3F6NgIm7lNW6VUVKfuIjC/y5mtZElNPgi9tJl3dQ/rX/qYKmm2/qI
oQqBhtnMOoGyXvLaFw8OlFVTNS+4Ls7Ef3QVbScrtNHd1vW1OxGMnC2qd0bPCcs5bsfXR+D0nFYX
+7xOJc38TtYgle8A9Q2bsKWrAzK1SQz+yNzYtP3AicQQTVu/uu5ZoF8Bxp0csEO20F2i2JbQytem
+EUj7u+rsghVSuMMsDQwUdblTeKblMaxZLZnDHudRUbkBTzhLHVXewE4/GATwsufFH56D1ZJjTUx
sQoMHAZbLCoxfQeaWYXJCIdJAw0mVuGn+2I3Kd+7wNbokUWaO33XX01XjELQevD3B1co0hnf60ss
mGmdptUNxwVWnFhW3uTBRcEIvJk0HM9HMIJVMW3ESUFB+Rbb7VR57afnaPSVdZt1frAKGhcvMR/h
7nbdrnTwmPqqNeiFAU6/EK9zKPbi6G2XH14WunTpy04yN7L8AkdsQ7SXJixjXRcpy3m+i44rZTU7
EKLvwAAlmoy4+VI5zHxA6vANtMiD5HP5XvH8OWZnqEyfIU7KS2PFnTWR8xozYXGRSZGC5IXzVVhZ
HFcgzqFdsn2kan/buqoqycV5w9+dFw+3NUlETQBpjnDaP6PoMKqN8ZzCNciv/CAQdPFSFDYLAxkG
ZMwrmG6D9uj2CFnE277wS9GOtL3rKq+njrwCl4GQPOxvKPtX5M8DvRX93MCZsStsJmhQFJs8WYkT
mtuClMBS/DCzdnOEx4obS8kD2RqhDaaPET1C/Fe3VBIuNJ24+0fYfXtAI8HEtBBhQ8m686v5hTwt
UEHD/Ngukdm++qHmiFnwimAZNJRQmpk2v1dmx/6OsROVGr4PqPqyXHO7flTp7qDIHYsBije+WA/Q
4efalFJA/pR6OygDNdxm3hIbkKciE3wxpEcjeLSxz8focu49dZCBP5u8xsUl9nUhUoy9wFgiFEg2
7I9eoGe3/J/vcOdWuWgL/AqSWNF2Mchgf9U/qfkalXf+hZCjI7MV6vhYoUfAq/5BDqNUS1r5klIO
vVJn2xQpbaEUeiDixi8Tyk5mLe3X5cjpZSMKcdo5miqtP8dMddyI+Cnw/tkVtXZsAtLSv/pfJXn2
bzv9KFuzCcjOY9PaARjLS4vNPBiwRujvclOKhJqQiE00cBxxzWPt/elZDfTReSXXEAbAmSUS5kM8
H8reWA1IkKJInxsz/UTKzjOxL1YBqEdns68R3j+QwYdJjC9OiolXc3YxLBVr1WK4DwwQ6qF/0ENZ
6C973leeTEGkne1rN6P/SV1dot45//+8/Q1NlIOMNuHIsnlJlca0mTFqkjnNDPPDONgxEjlManLt
ju4She+wBTn7aHm0IE6YlIunvDy0IdYHr0/6q1jxOXm7G3CfnOY97n+jAP+OCwwCR0u/tg1ug7yM
wiPOsG/MOjATHS1j3JvcCqqJJGcm36jxKLZ837LS7bxtHcZ5Lf+t0pK6HGIukBCmmOkX0uuWH/0p
rvzTy4IVQ33OlkbEKk+esa83HXfdOYf1G2SO0zeTTgxqMRyPtjjLj10Hp9aIcLsSxIid4BMWtQ+/
IE8vQGp3wRdz9UnioEGF8eH7fVLrow7CbdOkH4GKLWuxAG8ezO4FCrhKaZfAFkGLGhkVY5mwMc8+
sk7KHwvkrSjKkeN7/hhVf8hjP5inJT0R7Ncwl/Fl4ZJ1GfbwzEBeDq7hROJIeFI7zhdt6KHgDilw
Dh9wZaqgZIfDtdslBjZnrr/sRGMgh81Qxn0sj/W7KltakvtDCBNQO6eXXKdLEmuDCox3BJhZOE1S
9p4oSULTWGfs8cINTcH0QHKWI6uYK0gXIy0ANGCreJXHhqFRyoaDIKD2i3Sp+BstFJX09pxpe4i3
Im5irifAtnm835wA7E4CF8hpL4kBjQMGPwGn1uwwK1/AE/o4j82Q+oh3752FErzvZSsaeH0PWPld
2xr3yImoOGG97OO0ztFM/bh6gTwdTCjQW7SadjRRhAuOookbgMNB5Gd9+K9dxQxLGdNO/K1Wk92G
k+BFKK+LaPQBhh2AcNC7+iMMTv82InSBAkQcUiFlSnIJ0ROVR7me+1ADCYMH4Rb0gX46mKmz38VB
mNSD1c+q2AeA8JNzpJ9e3kRtt3xkuKO9tJ+sKQfisy1qwVn7iAFndaiaLKjdE32gb/WuhDE4m/WS
r/Q3XS2oEKZBYCsIPePDYXPmXX1lwcNjzUYft7rqe/wSpwYpI0OXdk8eitzj+qkDk8MbrIcPjAc7
amPh9BPc7BRqHnfiC0HZFWTSyguSy3s5EgYM0tPjl8XEkLoxrMOIpTjfgrU0IDYm/T0YYiFlp4oE
fW26A3IKP8LmflBauVxifGaxhfPuE2LUHICW+hjHicTnc4Qu8yTF+E3RGZHhEhnlAJQMtXvZxG0p
gemKeAIMJG8UatomWPhBjy9SyVpgG5EEuTiucbWYNX5fldqAavqY+vlkrr2lVqaYrwnQ0P6wClcP
r74x9zgoxos5EMDvn/6rekTggf09t6QHouFKf1j7zO1Iy+gfBIpK2eS7tMQf6a0dgank8BDTiv1y
dciUowGH5tPLy75kv0Rcy/7v0fctS6Let8WFfVP5EDpKNa69axTEvgV6ZJPJCwPXEBB3kkP7AS9r
5elM6Ri2SD2Fg34Xn/AZSzl8T5Io8SBaKKkWlGVOzpzhvBnjGjbkfrKQStvWwatEPOsRkk+xwmSf
xH0ViWdk0M9860G6U+F25GNrpPOxJZmBImw3aRHgXORUg6BAn+6zEzSk2ytuOjeWR5lFw9C9TgoR
kxvxnAzOJQ4AzG3TXrh+4Zymh+p22M02c0Z/E6Lw0OH1/GxWvUHRe04jidCdYpboNjGscAy9HsOx
LXvVrPrpKlfuQC2aQHqSwDWh4dExgZ9HjfCFAR/vrr88jxRmO2EqC+q0tS6hmYdS9Pw5zyfi6jEy
gU9fgxxBIgI4lj6FpFi9a5cwx9F3U5JOF5MukWSKQxQIzDpWlXbNbySQ7jZg6Vh2NyPsFY339f+U
PJ1W1jBhgVSzeMSyKtiYcgb+2Cer9U3fYMPqWQpA+1DtGcx1dlbFzOBoeN5C30k8X0RxGXckqx6O
i5IqoxmVqvYkvrY3GbkXZkGUvdfU5dV+nWu+QfX1oWDQKe3Q+K1/UyqyrX15zTysKxKtsxTC+O/m
lq1j6B4KtWNKR4WhG6DPe/Lo0Ys3UiOFDg2R2akOIdiWSL2Thf6HPLcL9MtHLFwEiQGOeSTxNBK0
ZWgXIkZtQWl73LhbgQc7N4tgzPfsUVMtsK8FB+L8EtA6h81D+B/vir8WFowrD2mOFQf6hjgTdQLY
uxu9Gj4WQwZvYDZoj69b8aTCCYFcNy4MvJVQH2WAwbQCEX7ZnY3akkWwo2NE5/t1FZ+6mlMbrxZK
XbBrdemQqim0VcyVRE9FZlBoIuxDW9qMErfvp1h7WHwZYifgcaFDt4PyILR+pykcaOzubXOLnpXk
5WL9cmjuV21EZvz7BpZWSaL/YzV56lPd/NcrxDk+oL7MKUDssxvEBY2nyhxf+/u/JnjRHiMUZj7R
AsHwMU4gMHDa3sZ4Ndc1pi5LNeWHrOxs3lAUKZ8ZuGx5sbkLCzpDCaddWAPnVafEp0ckbqx6k6qu
B/6krDAfQZGm2nVsKDPvFiEhbFYPX43NWyidbRV0NlGtyna4I+906rWqbg5QPPbSzqxF3fUH8TAN
2w0j1jncCFNk1GlSBy/VQ9JJ2mxocbklgz0IeKRYD3cemYgXI/eio/gj9tkh5IThX43YOQT9P0DP
xThfKCb9O5BSCBH3oR9h8WHoRgFxpi1HDrE6IjsZXV7lYvjHCLHF/DJTjlrPBefOHUjJdbaCtsTS
KxOJru1lzI/jAez/Sp2gOSJqjY3q4Me64Z3FGuaQwFu5YVNuuqFi2NjQtVtIXv4wOjqYks0dykaP
kFb+DKAAkmoLsF466lwOrET4J2+7a2eyaR7e/9X3/drcZT3kng3SlxQUQJtXV/tabd0mOwarrhjj
Am6RrtWVCcnIQCCPpUFuUqJfWY7JtR353L5Hl4zWzGM1R++n0ZTOYKLwKKYfU1ePSOjm3V0eFNME
iuCuopcoep0FPEt63AfhwAXmwF7GU5RqTTIo0mMXXFK2/QGgpk36WwovzHnqPetxzpua3q5XIVdX
eyET8f17ejTLh8B5BwxuiispLrHnpheu2fWsZ/un43W5paFHsyJcllIozEtAnJosCBN32tsZAh9T
cUPR6fz//h1NRY6EVC65B5G65Z/rbZgX6r3/kagBD7PkdEG8xNjkQ4Yqp/RQI0urJUB3E3Bj4mtM
pNzxGlJGZ2MeDuZy6GIQYcj0VYN42jWg8gW4PedfdheYB6LqQLVtLg607bHK4Cp0lt9s1K/bw0mW
ghjMP81BP7lGWlCVyc47LGurX74OcxrMRXjSTqCARLovwre7PMh2+fk0T+BzcMpnwOXnyDf1F1Mk
ksOsi3wsYQrv+h253xGO8M8eTcl6nIdCANt8mG7k4Tio0SOkT7vUVCglQTdnRKDu1OiVqKawhWC9
RfDKIY1wHibl2zPfwL+iq8+csbbnFG/MqTk2xwbaRhm34edMeR8I5pVCOw3D2eLYs9sLNBT2IYNF
w5VtLn/LbeSQc0j6XLNepwR8P30fYZOcRXXPtmK8DNT4vTFm76wsr0nYYthdk2wK8Itcat/j6Ref
cuf/CGlTzGgtRHzqYAwcAgUuBaVtVmBProu4L26kv2UbRc1cj7nW8hdkUr1bnVAmV/wFmfezGYli
Cr6dMeY82rGs4XyvrWcxouU9gFZ+v+3DLXw16WBfvDCkFq2A0LqCSh8IhN1BkLLL3/NWD9u0ZYO3
R7hfHAUvKM4aFRobXNj7p+atneRnbK8ckJOJl0Xn8hw/uleKYOPwEdhNnrVF+P+KTf10eYRhNf4Z
aTov8aiV35gNmXhdFofLlLlTM0Rgf8usouuTgJZ+hvvwhjVzvYBXmXZyxVez0pvd3Gdoe/7wmTBj
vDQqa+KN83pCkDNmtcqCbr2NqiKggVeR2UrmTtIv2PgIRo8384wkBGfn+LgjUiHWLbUkEW9fFaA+
7vNtd9H83hTpK6EqVkLb0nJfxk0hfDEE4bJpT2AId+LYFXq1Lji1X806DJlAXU+ZjPH7N53xA80l
ySvjclzYjVpOIAC5YnDUmoPCb50I42iGO5S88SU1YGd5M38BDol50Ec5FqYVBqaxV8PU3ec54Lou
dLdnlQC81Wq9obELRpZOH42//cKKxtmW0LXjJwfADevawZDdxzSMRp3aqqDjLkPdQ3oL3wVdlVd/
B29CjiIw6f/C6n/D9w6gc1bFEs2H95iP90FHS7FQ9SFG/TQjxnFDga85k5o0V9S5czF6pxnVzO3D
+QquaNvN3So24c3C5j7k4Is13gFwSEFdzFuA84+OM4oWLz+fyzjA9dwW7ulJFyaH9Qtcqh5ZOSqT
C1OQsqhHIRRHvyYi1MsCb6Jy3OPmKg5SH3XFJCEFH6wimkF4C7WOXd92vkeg63VH+0JTYEPV8xMx
jtMk/SsZOoL5PQ+V/r4FcpJ6A16R0lbeemDyGR8CVq0OSNkNzoDJlQ9Y+b/D6hSB0yjYtSctmMXK
6PljHLXuz3S6Tg/3qqwCpC42osZaBx/+5thWBLZNyC8AU6KZhp/qFXOsKIuJ4eg8MTcjaeSv/m62
ZcVCQ5/5jg/Iu6vLSl0Y0aqqFXl07kSzJN36lTp09NwHeK+QZkpzTt9I4OGa5w2U4UM108NQ2MRb
O5xAbLVD5HpHXoJ8lyb3ApABjderHtMlqE3jkexPdmwHxCdY2svmhw2ahjLNqy9Wv9W47wJIGJnm
w0j9nCOpkSluNKe06zr4JIZthMoALx0CAHe83qPaJtIxzXOvxrEgZMQtjDvMk1ubPmPIz4ZBjOcG
p2JQawVvwuNctEdXKM2DNR744ArOI8JJRD8VsK3O7eNifNvJi14dUSAhCrqNug2Snrxh3OZIQevJ
jqrtkwcM8F+y5K/8StTujvrjxJJ/Xizmm5+3uCnGdkj77e4ss1ghWtenMttpCMXbEuIhy0WF5HDx
oMgBYYC91/FfVgnDSxDEj1UkkHdR9ssWCOU5x6nZnjbeCmn6gDdSG5BM/jHPbMyhJIQ/TiQBHdSC
iUc4soaKXhuM7ljQxTM6isDRZVGdbTPz5svlSsrWfkI11o8sKGAwTyz/MpPkKvL5okgcwMDUAR47
34q3XKHZJFSZ1j7sGyDbuTb7YbIBzCAISlg3x9t4F1h0KGg+AwZoZKUxeqx4qeUS8cI54xltlz6p
Bx0GICLiFLx5ajwgB6wz6SisZVfG8kPRUsupX6rGPh+iM3AGuxthCkIoKwahfKo4Xl+2gZ9lyQlS
8QWW7yTqLgGafEEYtQipLr4gFQ4J0rGDKlQPN/ki/KPCC5OGfBCS1uqRgoVLLmr2FapB3Bq3qZtT
yt6uBa8vsDJzBXnY+3r8BsRpiPZnsB7UmppRFBkGsqe9u6u7WJRw3Cy45I1ANZKE8KvaOi4AVN+X
mD6Cr+/xlQFU2AoIun4VUURI4hQN6YQ6kMoD947lt/eIS1XSzltxbU6D//Gi5uVnResCu4sPP/m2
pVlw/tbZ9n3AhWXDxpx4+3V3SDTaY8Ttwrp1QsqYY/A8vBdwnvh0VOwhaj+eeyXJrDhP1CdJSQHa
NRfruZM2BYj3Re8cs8Ss8Yvx6s1163lbb2CtXrw4ANbICczh1uR5ZIv+sDtBayMGHvtcn0siOBFe
ffucA5b+PwH8JCkDRJ3W0c3H1c6TqnSL8QJ+z7zGd+lyiOrbUIUPoCgkJ+DO66U9XYuH8KqLwsQo
HSmOM6t9dTvkXATpYsAwvntGEPYQDqCJ7bt46p0/G3OeMqHhNuZP83qCasxk7QAHBhav6liboKZv
tjghjPgtqfsVt56y4yjcgyHc7IKLx+ZnJeJMQJ7GRvI9YqOq9atC2aFSxkfHcv8LRQ8CD0eMEdjE
qFXg/0jNjcOsgh1fY12niscP9It0VSmzcXJjDBAtNnl4H5YKQDECT/SpRW+cMYhoUNu3JXDW8dIU
t7P+PE/qHwddrOJot+i5ftmuZTqyLFC0hcD6QuOHXtzMmDJ3rdVzU2fgy0VSbeOMxVk756YiX3jS
1KNtbZ0L1HwpOUjpbwNlE8SAnYAqDLM78q3aXixYBiF50nzhxyU0NLWRqa5bXzOpo3qy1ZZyBll+
kGEfyuTa3oz4qhQPW/gC8DGADl4VsrgNRw2qJzQ3m8+fNq0gB8gQbw8xNAy9sl3pLuh7cA3Bhnpp
MnZzf7ZgFOXL8VaH2NKOYTFRDliaV47GWdobnPTbbA8ujLc+qo0+/ACAkPCvRNsGVn7Xgp4FNxUz
2owUhVB3cH8ESJMlSCbvMPSJEDu8Lvy1CSVOQkDqGWG7MLgBrhIyh7B+aT8OicRemjEReaBWQWp5
LsKSBb8M5mUdz3u/yorTOGton1OQPQmx0uc25DOAYYhhOmIpuEQiXgAu4JXj7KtTRgaEk6Jb4stG
tr/ubb1sumdI+SZ6bhXDYE/gR2jGQH6mYeK0bua6ij4UjJNGXxOyMgP8RZK5l3UD4dxzWS+J1dwi
8nFohqWtXKEBZAfMy+P41e73rOWx7VuKH883xP1o+qqFccB/ZreuOEKnTZKukI8G+ppLjBmGQAAM
z9w/LbuMm3yiNO7k9SgyOCbL9bnrbQ48POb244mOoRloaWnETKntlFo/feapdn31s6CJh/oSEpL4
gD4fNMS6QSrTyRbkA8pNU3pfed39Co748gaqRuokHMOQTauVexBfaTDHxrFHMx5J3AUd/T78yoOb
hvDbBMWmI48ZjvENW6iQnLCWztFfzPf8VsyH/Wl69qoY+KlZ5aYn8CU1Dl+qRJ2Af/f1WB0thmt/
xZG+9fejXgOcBH07jhOgFW9tNlT0YLL/wX83gXlgI/XUFY+9V6LRSbBwRAqfDTAjGlIBnjf31va8
43CsUHuamgGgSVjn8O4CgWUo+q4tZ2vlFi2uNwiDjzPNbS//t+q+vysviUv/QKLCaxq+dt3Yki6O
6U39c6po/KxWGiEt8yQhwd1cksic+kNwwKTfohZO/kJBkpoIxJhTSP86tUmxbESx9Oa+3BgK5Z3f
8rtLLf6ib5ih1VRyvRsgAowWdFWkJQgv5+1rrCz0cftMxKy7R6S51RI31UZ1u4NDCYh+TkDX0dfT
iBshsXVN7kAke+pLOr18EFWKExr+a4MrzLYfgqIJ/OaG6rkeVkIStU3Alf9gia8Najd6grOQMYoP
XpZE/14MgM4sz+hROWevdfvC1J7yxXaRGK/UOj7xYR9A7t2uJ+1YqT75RXUVMMqjtzledOrUPM1A
3ud08HLdl3RIOi2Y26OhvwyzMqy1j/BksI38E3mfKPoQX+yrXGtDjo1FHrB29G4IY+dUVfHkfI9v
I7sABWhPheAIVlTJKHtkOCCCAwMBAT2dNUS75giiauJsZbHntrVQfBP3E28Sbj5J35b2S4dPRVNm
VBkbKLTpk4jCLROXAstQcdOUQQZHwAvgIbEVUgneugY6azFt09BoruK+GyyaeNMt8AEscjZ+w0DG
uNpymYONV5sE3TH6D8O0YyUMAfV7/VqHcBnWTB/KihzBTEiYkdl48VP4NESny1hh/VNFW7b50ZlG
J/TInP8HFQplHe0ndolBl6xcGjV1pSvGBUxWLn2THcAAqAHqm1qOUpV4QW8ARTqfiJr7oJUlaCqc
cjzbuq77Hltzgaw5elZeuoEe/UokclRz99h8r1lTPEcCyKBCoVoeD4q73HXod96stWND4ijGIabX
MSGBSzAVd/G4P+exa6OB2RyurJh1/gTL3aDXUXjwm0nnXe0FwL6CgZKgAaWY+J0rtqogIlSktEA0
njqBhS+dyYxUuF1BtE9Ciq8xwPTQQ/NJITEd8nV14KFNCrMnpyGD0WqMfuQP27BOpqjmLqa56cKn
2oSUQwFRXtX4VvBrWzW26YE+E0Qq/jU6jvRV+ruoGPD4hKGWZ53PNZHBROQPvwb1HM/iuo5VUtkY
CddK5uqqhdtQ5WuvgmaGN3+oIsRJ2IPZ1O2QQZd7wzwTJugwqeQNgoXbCmXi7pn78A+j7fnnZR1G
QPeRSzdl/ZA+ryNoPxJac/3Xfc4kKJAiCo3uAXzRTGcxhlaGUC9AWLsIJK09R/27cQ8enbvCMCRw
wikU+UgS6CcdC9Z4gf92N7njnVMbMMAkx31hzzTGkenRORvghwElLDTTAjiJu69srC27nxoustoE
SJuorU/gNNGDlCCFOA==
`protect end_protected

