

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
cPZ8vU4rKWICMycnP8ASghxteX0KiiSQpWJpCIK7voNSpkWhaLkY+/QNXKrCWexA6C73eW4MlVqP
U/aYYyUL6A==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
LGoeeEeMUHkj3xBumwl7JSHXwdKJWR3APWiWCdcCy3wVC6g0GScQrp7fjvXp784YBiHqjtsyG69d
mOZ3fy7Gj87kc/h2xvc4Kp6GM/IiHJc0mbPVp01AJelfAExlIEaVGoQkcAXR2aVikeaMxuRKkb9m
THdehu5n5eHx4/tJQjQ=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
aia+xx8RLMhA3IF4tHoW0Vw6LtYVDVgU/c3FBWk9RJ/SaLw9lkXng6eXJGNs7uUJXmkzrbSEXjkp
9p7xWJMhovE7nwsp+7RydSgRQ0ttqPUbPZE1eqSc4iNU9Q/KQ7cPFMFwb6o48JfKidjAmSeXX5a7
n8A9TbJ98klc/V+a8Nj+tTPfVP1QI9dRmdzaW2w+actp2BkWAgSALKaGkzvCVGa/MpfN/fdLNjxo
VsiL86HW3arw5N+Ra4HD3GVUtLt9RoCCVRrMaYywuIwp2m+MgGVDwi2f2wZCZ3t03UamXKangjoy
PBei/XvAf3p1OvrOrKNUCVdwEg17DQWfBwZyYg==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
iSq3so3iXhp8LA8lrAo4ElVWkZ4sJhg+rWrioZWefLcgVs70gDbHsh3ghf5w2wiNXalSfMYzUoxO
skfS1+28WFbvBvygndpiSNMXeXmzWGrwBeHtNO1nR5azyndKvNsun44/B61XF3kTINCJNR54A+3f
0Ezm1jX/FmstQisPDpo=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
fHCdwSqtdLKfkpdCYo92uS5kFXmPpII38bIISEYuCqZyK6/BVCrCUL1HNVeJEgqGnb0uRqkye2CI
eX2LoUaDxy6iVejnRrRRAgNtgrlZcFVc3u1KxZQXk/12l8pxvVZj8jnWgIvX3TEsZsoZ6w/D41BC
6xhd1LtUfJeg6bsnb+yBYV5+H8NnHOqkZuFtJBsUzS1+4qFALyFqcNVJhhbdB0k2hn6z9cG6wZBI
hB8OJAFj6xON517ug+qP1OJf6uK1rHsG0pxYXoT6xch+UowAmLY8V/4+ShcI8rx6DLYpPvJVhEGV
fj/RQD4+HY8CEDIrJcGjF+Rpk986lOFjZ/hvRA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 11888)
`protect data_block
uMl25uLfnUBJUXfVJY8sFk5He6Hc+iDx5YtbGl8rnXi46T6V2xOwrP2Ym1LXFvlRj2e3dNZXDW2u
NqJns2q0hb2LLhfvqMDNB0rpbnVA+LObRq7YHvJ/B2Ed/cq0c5OkUmU/Hcbx+t221GZxMyMZXiiZ
ippYNBUR7TiuSudPi0LpmAbHLtC4LqJlxVDOX+n7h2Pq3KZ1NuBdjdU1OYrfp4etn0JBS26W1qUS
EGH+fsRnsbTywXHrmzBVgQr42JPZjHxxfDvCU/ccp+4xt7ZderVykn827H9vPkUhcPU4YK3DMGpw
Fht3rG0qjdK+mkNc87683ZTguxd4THp9l0WqphudqB4IsewMFZFkeuw5+uw7lKJyio+8Srcjfd+z
kkQoP5iSBWh9PdHOXg87XQeMuI/OtyZqKN3I4NrLdjwR1w8zinKSTWEZQq0ze7zkbQ/ivk56L0Ru
aRO64DvKCzHGW9gyYLN6ZciOKbupo3MmlFxcoE3WHGhS6WeFHY0yTE7ra/c2pQLg7HVW+HZWBrdN
1Gu11XFIpAjpP1p+XcTPZjCFROPkEYqJ3b4UzUc2QT8ioGAkBWQWbc81eEXqACkozwdlWFrWPgOC
T6O/3hydzDwv1RU5igWMaRqqIN2MtJfojyhHXpS7WJ2VlKRwp5WwGZLgS6IJ+h/t2gnNJXrW1u2a
fleshLqVpG66tRjQfTbenEuGVxBjc3ffclHNdBVqK58t6rB9sFdkZMuagGnHGmwqu6X0Yl09aC2S
RNH1jjPAxsSHtmgPxWB3fUWWxFWRbyer8uBRTzKmAr+4pARxLymEd4SLPV9L4x0Ho75J0SLLQD3Z
F58J4sahth8CJ356JSjqFsGb69idQQ6bmxXFLQynnxFKlH75nDY0jqmuNGxI9rqTTyKC4NXbcdDH
LLUhE9qAWkTmME4EPRU/kfcXiHU37t8MTvAeJ2YqqR+QUCGLm8QrxHGt4zwbRKUJqCvUlih33Xfz
HFooA4tO5lJFKi5bTSnAOve3v284kYT92wHSDH+j5JJAquaDPe2pT5Q5eGD/mCIyGt7SWRt/Lhdk
0B0exLpsO7z19rmBF1v4Fs3j5FTLntmglt4rtBSu7jYahF1ZktqUGtxhgP1nKowkEhbL4tujqGfE
YfLzXENrwi9VYn2vJpIdIBY0mFOiBqMorZOaSiKm02wvidSl7K2lpYu4ImErg8EgjhzY/pQ1RwCQ
Dho+TWzh3OKhvvJpr7nWiL57wwBsfKEWXEqNPTOjsL55gRnZbww4sgX+Lb/cZaLfrn6JuzbyaJre
A/1mFs39tGTaZoMKo6K6AbNmCJdGJAF2HsNmazxl8OHtsGznRM+Nt3UuZ5tf7PbKbRCf+0Kt48Xm
SPUQ5qh9mXC+RmwMfFwJYH6CLLjwFKWB4+Ytg/F4ypGBmFOMJ0ZrKMD2PVma+QC/qXcmeFq9R5K4
gIPUmhR3m43zSBINBjCVwUsoRjm/I8KVTXa5r+3NTdrSFuozCakONEm3IGtawHXdzEJCq0sDMQoD
hP1wxYiJx4I2GExz4hzEiSe7SgoH1gGzcAWOizn/UYxLz0gBvAR9uC9efPCRUolRqlg9qkC4QJF9
sos5QRP3fVbi6dSoqVsBY61bWZADzs+xD1lgpqij7bBVawBSUng9T0UJQFEW8HVmvvGiJz+i3U5y
RS3byRV/ifYxx9PrLCqyqYhizwEGMHI0q5edEBYqKyh9ml8PZ1bDGddT9s3dWjzL0XE8Y9owk2yv
i3+t/8ChrVvAhfsbQ3vuBcgZ0UmhTkx02GIEgD+o+bbwjusWak++LQ8Md2yDygiYNXpzV56PLa0X
vQtZJcJcNIhP0cgsC0+aN2pA9R75GwSX7rkisT/IMFnLYs/Y6pbyTOjdRh0gCJgN+Uy5tyoiLa9T
+0H45qoqayVs9yfNGIzC4Nl1UMPYgzYTkwBo6bHtQokNftuc4NDe/4PPH43KR+xh/JMAFfOmj8vI
oluPBTx9lhZqoawnzQuvafhqDaiS64tdZBY/hPDpeh2ed4ErAxfj65LKeMSLIXynOSnfP473f1lt
ydgwZJ557q0nmx6quIMs9RiIwPf9DPUJNwtx4RG5aRDBXnD+UE443wTrh6h9wRQxMcrToHH6l01I
QAxiESi9BIXs0joa7YiAP9xrprKbYSqt71rLakqDJ3RfxgyNLpKhwZo3G5jveKU4zBSKXLeqxsxa
Iq01iKZd44mDSRBq+MfTsWD0HTsvST136LLX9FkdooFpZoJJrb3t4Pfe0GeLiejciBA5VI0js0kM
yVY5mnSNr9RQvyJ01tWT5gthGxqmP0ET1AJJXWRDbTSymr2w7CGNt7fcHK+1NGRkCvN66Ca642Nb
qQjOVlbDzeXfYmUTU6ZJyvjZrqC0G1wJepxwmPlmY3TqXu1k9n0sOYmO/TCoG/KrHVHWkbAEqGyH
z4lkAHdyh+63L0pMndg/eMplZ8+YhWde3SnVG8ULcobRmA0d1W0lsPaMp6afkSRT48SwJH0TA9+8
yXN8oP62WkpY8AFXhrfJwVW5Eo/svVXTdqwl/hycOVa8sNrwRxj/hdaUMQfJ8KXaoqrs7ZGg2i4S
WuYH03BL4hcO8SMZAHsf72ukLJfXvSqAeZdJSvPSN0HOPngFsphvYM7IvHido3b2HyI+rHjGioBz
vxiA4j+an6XbuTFJYMZbV1KfYjAg0efKmc6qzu4JUMPCEybPLi7pgFnQ/n8bcpmRgwJbCfCD+n/R
R/uZcFBDXzNbBm5w5Tmyk+ePYyFuC4KZzK+dDu6GAbDtMYnhkxvSgfrbOUIw9z4cnLgJNfTVn72K
yJ3FyFk7TKCjAxTf/WgXiYgnK5ioxT6z26/FEvCIM+swc/WbD619Bl0+WcanshOpRQ3O2luIY2Xn
LJSGrN3l0WkGioKCh+mbpT30qPSaogkOKk1SP8XjPj9Jw5+GZ0KLSJorM3Zl1DqIFDwXL2mAE9n6
0IgA+3fVdD3uiTFpWST5T06qtJqA7293bRuwSCSI42pbQSUtUdvCvR/FJVBxm+b6D5dbJWkQjLjL
dr2cYtVslYM6nrv7aQ0i8uZpuKT7zWxoot/4ajaNYC4Es1Apw1E0HggW6UbruGnJacYXH1jyycoI
ptcTneEMmNztuqTfxcveFzbxy+5ig6p+NkkwnR02xxf6vhSD/DVb0JzNPr+KX8pF4ZHD7bOKefJa
RLMC/dyKfP9frZyPH8JU/PEGlYLrXTz1CaDahl815+6l1nrx8seeZWx6K/nctDPuv3fNOgoMVkUe
u2c63DE74cwhmxvVxI8jGrPz8Nk/IxMLoJemXC+HTh5KOMSp9Ap+TP9nKL0PkEBdIHcbGkZY4wEY
nmXd3jdCF/1tGz2itpIn/MztJTNsIOX+UPD/Cxptx3FFmlfWuIzT0GTvqEmMcXe7K2bkhxZtYfCz
v8z3LfK1cDZNcrz5d09NG0rIXiDPLRCR7hTvXkwvGe9IwSI6lmdjrE7Yn1U3EaHczK8K8+J24q6e
L3cODVCXJzCMaasFgXpTtBUik9iHa2ohdNyWlNaZ09Z5yWkgXuChxpgP7SA13akY5cJSm8bTiExq
1ezlAyOHFaGtQt4qIT6ogMEIhc111E3ljiVpYh7qrvj/C2EfSaX9tytIcRAdb7IXLbSDxiHCV8dJ
iOmrpXZiVfmFvWtJN7DVeohTEU0FZ4/B7O9WBAbgW7wcAlUqJvZNjF36isid3nKknCV0ia/2SSVE
N6TUBuUVRfyDsyNKZrBaDhzmPK7lpmdhKsT7hBL+H3Vr6Clp7NO1p4w5mWa7I8TMwwMDLiCh1nRS
Kr+3FPrIqB6UZWjikculLcO32U9+abKJ15UmwBfvkE6a3t3ClMHPgZ7uLlH1xrNSZZA+rEJ1KbYB
tR7tCDoTDiK83RgBSVJNUTCXIxzgxxdwvzoSx0h6tAX9VCczhc8KgG4ROYRtF5go392133rA8XjS
84cuPu+zgW/OrJF2Ztcd87pEKoUSEve9der0+AD8gKie72JYvcV136CNt6u9ULulHvNoC2IZNIHK
ISgMyhY9HcfLH2rzzdtBkO++DQsnhWrn7ACLgkN5kMobHaRMMrmsIPOGkQeZzTs46xkmvU8PPiYm
RSrltfzJ9XrZ75YXYzqk3tB9A6S5PhUEUXLnT/ChVcJGzzGUzM6b/R1EinSiHQi84tWrL3HBnNvP
SfJKuIXcN8hpXs4hv/LpGj5XFFrKO3xaQXC4fJfxAsVa8DxZajuBqm1sF+rOBFaLMuGyCprnm8Kj
mqZpOWHplvDGOFWrAG85r4yrbmC6z5Ixf0ZykXcsDXt3VrOHZJ9Oxi6x6W7vfK6RuIkd+1S85Dq8
qygJVdIMSv+iHZZjuZve8EmGjvbJzCvM+qj5uyPg/4Wntaaakk1q72yeKK/DTlca9nRhyGsSPxz9
Q+vUglqK/bq7e0Xedg34zKmkNpUFKIW1IggSuZit3bTEH7Yy9GeNR2JPxV9ZYFlvefEo2W4Ro+Ky
1AEcjBMBYOxQeJo2rMLff+eoPP9vA4VGEJeQ+HsHQ/2JpcykWEEaUTrultB56CvgATsheZgcfEMp
X64LVkJhstUae02kh0TcQkCJRifJryzqA48YwU7CpYxbcqUV5MsAOQfXIKI/hWPAfbURevxW0hv5
n6gJKp30ig8gg3P5liDjAxwdaFw+vbZohAPsPUZo789oOfmc+ynKZTWlyjktIxXKKh/CKp0DZoe2
4K8GTRjIeeP+bzhSos+G1Uk/eOIQ+laETcok8dGbsnt37m1qElJ4ySPUmH8XqybsQaR98PplBju2
DG1KT53eqCLwL70fLFlsr+YFbyg0Ck2oSfAWOLZvKcfSFj5CHER3RjlHfdEEZbMhFlQIUfktNfJ8
rTe/1znzu4U0W3trfC4Zf6hgfmhMPHIIg49pxAT4WGzxrI0+RPtCEKERRt2K4zTJPOJ7YjKfVJm7
FZ0fcfC+YUD/IIQY9kuQ/unyLhRiRfcQDyQP1Y6u/U6PPKSFqg4vfI8BzyWcGlDdmgSGPcdFPfgr
hLk7JZpqmFWBuzLlu+HkFwE7Ry9f2B+dk1gSSaGzZSnU02WMitxNzb/cPe7CoRxbAOKQzgq2mD2n
hmied1J5G9igggsVbZHnhUZbAflizgV8NPpACFEk39jXij3WNyU1Hj2PaLUJlKXSg/Ln0bWFyzLn
MMOcGBiEQsK6axAgTMrUC5vCTaxO3AKpVl9KiuzZQDX4qSvYYM9hPPKz6NWvWu02p1H0rTNII+Ul
aE6zfnYK0e+xm+d26hzCVy7JEPj49OaWTq2r4r9xAkK9MSkDNeXc0UMueg2M03W95Fb9bwD6cY8o
4VF1R4QCQMc+yT3Xsl4WXQM0eD+or+HQ7TrxM319bhByCwus2pBoH16zs2aBw2nqSrVokwDd/bD7
hDnq2akptralpnvuJOMgwLbZnPAroahcbm+cd626M262qF4o/g7AzSDJ4ZZlZ9bU0pUhqabDdWKz
FWwDkHPVp1GDaq7OwMxUrQM02xZGZFwk6Hc5VRcHp26mCmGc7Opu57EmT80Gd5Bu+sG2C71ydbga
a16koFqqDSRmxEoor5vtv03PBFuBI/KQvD03/EB05i2TxMZB8tuQ2y8lOwtLl5y6PSrTk8lw/6AO
U/UsZCZaXMzOG7haRb6fpWYxx17hPn/KTr9MVJr6ZBbdSfp7ifHVzoncjkmTL8ZwGhfq/2aUSYAQ
xA4x5UA+xeyNSyHo3Us1M+sylapEHdHlQqyf8RITKCdHEg2bpa9X0aEeDZ6sB3zBHlDxez4osXkv
fD7GdiVQMirQWcugO2Bco/7FubUy1gvywrx34Rx4fszvR/QN+gxYsgdy7t+ACOD4mIozDrvqIh6Y
qVOhjThqL8/RUp7gmBADXtookUoWkFi1Ex/E464VwaJI5RVZirRlhdNOSfh6gDHRDab1q0RaacG+
/VZlYJbqPH1cQc6fBClJ/gaAaTgRQJrB8+xVFDr43c+vcPAD/fQpUGRujA3vDJ6tlrk3THQ3l8ma
Sj3FlIKc8RJhPe3eBIWvIvhwVXYK20id5OVRd+7E4dWXQZ8EuFB1oSyIJ6Zq3wtQGJ77BfgoGyHv
iVl7pDhzC9ULPLlFUqO4oqQu/nAWwU0bmNJJuJ090Ck77pOkEfGiySI70Q7j+iWCgOJVNQu/A170
lrsUobo/L9VsCfGlHur+trcV3e3/rwyI6x/45k0U4wBjgMJfVhrnaR07J19cJgdgC0O63bXaTGVV
nZIOC93xjFPl8BLb4CO/3i1bC2oYs9x2fLaYiekRMmVO+tVHS2ak+72aKDZbbXU2K9sLu4DJKR91
pWsTKS8gMejDnzUl4WwNx7/5mlJoqfLdZNeVplDNpTe/Hvi5QZtQsItiXfis30gg6280IS2PV838
Zt5caXrX70WS47y2I9LkBN08uR/F8NutI0E+GtmzhzVsfQapbhz8mZ4ookij7FcjzeryMT9kzVK5
0iilzzqPdaLi5wKrGE+LDix7481rJDbinaHojYXZSN0zelM4QlOp9EMIAGLyT7JG7qknketXaM2h
Hs27hZmCZhizzqH0a/LB8IqhWdON3QqARD7kcUS/Et9p/ExYKfCMW0Mrw2tMclZc5U3Geshi+fCa
VL+fxu4bSaG42SKrXSBsbCsFraLwn6hvYZUWXJvf3+uBCBLmDrkH5culRCe0W3CuUwoQC98mFUVY
I/1Ey3A1dDcdhg31S8oDHmoFGEd9C8gknIDiQ8kjLVXEVrMqDwF4Ca6PmHvxqoVmRGh+BU54MmSH
JSca0VXZBfBqgKwkE60/EJ49l4AxncpeNhilPffPXtdcr/DT3IRqupJSyr4yteN82LoFtWicP6b0
TBki83zlbx0bYAKGXlRmniIs1t+veAlwLHns2UW4UOk7s+J1M65RO/RL2YPotfi2zPyGsojETfXQ
z4Rw8jnTzj7Bk9YSJFRBIzEiUlxLfyCOrQEhvBxnWRaETfMpSDxAXXp8/mQSPTOC+VH9wvOZDGUd
ARIaPpOCTAt1Kp3QJ0iTMGOd1/7nGBtD6OspUSdM/orT5pYvOrwwEX0U6UBjH8p35ZMMKQPby+CX
QbPHUymIcZD8c7RqFygQlcIyukT3zpsngqlKjJW5gPNQ26BF9+8u4DJga2Dvg280rLpmsqPh2eHh
skqlHsz/n5h26DV+vC+0gdhkVVSoxZ9DOQ4esxbpyOtuaO5nsBSm1sAqr15zWxiSO55XBVUGurIQ
uddzm3xUuky0TA47mhQHUJp7hncHeeeswjl8fR0y2mVpw/foGuTPniKsohUDHtWhogu9koajpJbW
qv+t7JHwAExeJ/1crBH2N5WCv/h19zmBHAGvZoND7isSJvv5tiGFQF2HBRBHxTsI0HhCtJI9KCTp
7rcYMuszkF6lFVlhhoNhrrgzqBSs96LaD/BdrVr+lUEmaWJuICQycBRrazBY2YsP+XiQ8/3E0onS
vKpnAmyTtG0cX5v6gUM+zBvVzZ4+8WOGbS6IZFDcoxVODqD0BX8g2c4vjn6cpE7Um6cCGwomm/45
nBLJ90zyJWfmZRXsDCCFdzxcZO82WfXyet6T218tCpRIfESL95h0vjz3NKe9om4F79sHro/um4C7
8IlLeMnreGADUO7di170fM6JWtl5D/cWi4cA863C7xS9CcwgJsiAnBduTb2YirflmeszdyJ4p2xx
MCnx/7ihgtFD/X36One75xXKuEfgSxqvaf/MabECFSFd3YgDvo3tbt8s3AMmmF6rZ2Y5+RNA2UZ8
1RYoFRy9IJC2VPsRYzbJtB/8exgUDy/quNQXL3FhS82T4rluu3WUZ0I7nPBlWGl/K9hQ2TnaFQaW
xOxJ1qxUY20dl+5NdZq3MtL6FV724lejciXp1z7lHzfJGJ2pW4QOr67n9nmT4GCD1Vg0sbe6OWy2
fmtfgiSCE6P4Lktw896hL63+SwKGLZC7x2HStP1hHR/FojuhU2ZOZ9Rbiv0aPKkJpffyPKOouv64
ECLvcg5uaSKdMHwmw50XGCpHwa7yqXPRXPIipnGD/+fRi+587Uvb2k70IMPifGAAmdhn1HSIq5vR
FtYBtx04+MHaq5IwavQAy1UlO93YFegzeJVmY97JtcT/sRkntwHkObDZMdbXF4dYkw2xuX37ahc6
W/Qd8SaSWutK81cq8my2pFmUt8xvefZ7Lp5pkiYycdZv+MCOr9ainU8Pfl9Gu3LPQ+UBVe0PkeVJ
azTIJhf/lLEiW2DnvtFYi9jyaaRlgkSZi8Vpt3QPX9pn/jsM+asAx4A8jIp7YryLTXelzNBzBfQp
vV9KHhLXi6Lq1bOCOxMK/j3MGm2pJSI9FGrcQUNPe3wtP2c7kfvr5nfM0AtCcWBZnUR/okj/Wlex
WxgQ4FGy5wghnnMVzqIQODXrB3jjCuKl+69RNOSUT5Lf8FY7QiMdh4lSvwG4kAZ58EKRaGd+OAgc
2q/ReGKbYK+Z86TLK2jqx2yWAs6l7uzKccNLQtyQYgCiLrJj7woZXdbfJc5LVH7jL99FdQppkBFt
DUog8f8yg1KUvyZoGdtfs9575UqQWHQt/UU9bTh2MkGr6pB8D1/gZunaxcaw3QeIoZ6IqdxQ7dY0
08mtI/G3QcoSpnFaa+iVIUYlBEVCwfjpbbdJU1YVT9seWwKR7WAF8Q9SZ3ae0HOm8SMwStkhrJxQ
hQK5SYU+JBxdX0G/1EtPHAt9bASTtlXKt25Jy9MypTKk+sB0a/hToMvRyz/lDQVN0BV8NjrmL512
NPpQPd5zWF4LOWtx31iOGKiKvuBR0tTUCsH5hZHpOph9smnbOteMezA0UScJoRYKLS/ywFbqsAfV
QtzliuWk297qv4qblXArcUrl8Jc9z/A2PxCkZ7sbku7s/Q34HcYeespm2qkVtSguz73t/UpBTOOj
t6YlANsHfLwb7XjmQbm1O7TA4w1fzTFCOLBA5YLmS+hqV/uXmkdOtMGGXA8ohcvXmB9cPTSE4fyH
AobUWwagc2B9t8s2eMVgzLZXEoGwn7EtdyPek3Mqcm+6JhVQonxqytATRZa3CljSGZWdPsbtHRJy
Rp4tleX0VdbjIN3Dbc2oJ78st4F1zGkWmS3BD91e1pqVS/DM2xczhy9YoSNn4AbYnxIO3RxcSCjr
Qv3uWZfMCTgtaXp5JI2m3aQkSxNGzHQGR1s2Cxp8ICUnJ/6sGY1+CyWnPrAVg88H4OzHYYa2Z0Ah
JHIEf8ni+hAsRLSycBYI8UGrWOuOy9OoVD5IGGmJKwvVGkvTPG1G4LABFgqwjbfH0UXWv6MGdiQs
+TaiIUmXTvIIGKsusElgrKDq4PaIrfc0dCXhhthrPpwV861lvN/OmNMa7+j8+tjkJd4Z3r2IwDQz
8v7a/WrsDP8tVl7wT0xPgfk2bOk+tFjixRwz5d5wrWJRornbRfVPO3rPFjHIb7cJHD8ZUHmAqpB/
jSfk9goodxQ4uqr+9JNkPnKmAaXzgvYYKi6jgHhBVX18k3te3R1elAzL6S1CQaD43PWUM26myrGn
+7sWTzKaOwKBljgME5vSg2f8mLvH/O30JE9cLPU9zl54Ufq9Fmh07SPKPdrPe2S3IvoQlzKA803k
QbWnct0kAvwRJrbQTUfts/DHUM6U/OTCQ4q6FWWQToqroPvSCaTcUNvBq0CpEFQPCuV03h/b4Q/o
VITJnV34K4jrIdy/i0kC2zak2eNdVQ+EQsLuWAk3mz04377NR5UcNQKO5mW6AM8AYS5Nm69zq9C5
s5KU5sAg8H22XfVN29zQfzMRpwpjd0Fpxdq6ykCnm+ziDw27MLbRJZ419Dfqz5E54H0d/V0V/xNU
bdEJUEVBPtqSwwoWyTifScTdKgjmACawFUHwWwhwkgprmvUF6kHWhwvSaTHUsMou9rkJpp6mF2XT
qQj3LW/yZtQWp6JWb8SQLqP+2XLo0R7uXzAT9ygywXe0hXSQQwYTHaQu9txj+z6gpY1yKBKpUcql
fCapC3KaDr4vKdCwSPPeHNyW3OIO/dm401MN9zfNEB+RNJ6Ue6nWPV8B2ELac9patOX4Tu9Getag
BtQmE8bhPX1gzS94Be8ZN/Nql+TV6UWNpWQByjsR4LTm1hBTWI+pZNQgI13a3i1/mtZy61/oOWe0
TLvyxy8bk/nRiZztwyFjXW5OPw0mKYtD3d6Kk3OptZiVgFMEzSJOhZ/MxRiP0c9J9jiqZTYtt9Jp
Jtk+bZeXs30WtxplOW+lJJJBuvBKcwdVMtmqwKlTdGCspzMo0+MzQZkGr0+0IQSpzGGRrVnzdUsA
ZKEWPLX+ixLGQgMc1Zy5/sc0m0kKvnXO2N3wX1OmLvm5qy/2fv3YC0PYfUQMxKO4X2K1eekGEztW
/0URX7J/rqiVKvvcAInsWuaDzSPvvE4gA/Z5P9cgsUMqgooeSC54mLVMSlcmC/V1ReZg4c6fbPni
2IcHT1gIrnJ9kJBisYmb2v/Dz6Gv3GT8YlxFWqW1HLygR8NCqgMUd9gQE5KXtRrzk0zckbmmzxk+
vG178yQcHOHnkinaPxi2UX0KZK/9tFQlycHWP9IEpKl7AqlW9fKpTbUQ8EzmATe2xgc02P4JOw5m
Ja0psdLDS+2dPaFFXuma0BJf3DVhSF2vSQaTZ1mPmG+INFr5miMp+Fvz2jYHTQ4vcHh5ekzvrUqy
ioCr4XQXLP5GmGzMe/daJ1+fS2EvdbNLTzwxaYV+DDnJvPpff49CaTZmWpg7shVhKmqK9lZtLlj6
71edX6JABBVbWIupUQvBN5WTyyvup+qAht1Mg/QNDFqPb2xEgNtnyYy8RVzsHV0pLqt6ueOOzih/
EUjkuV20K8c2EFDGoMNIRAJsqLe8EzSAO5Mzp4bLntc0L9Ug3vCxcUBite+r/Ez69pGSJJPHTuGT
YkpLIJEYGZ/vTXShNLvrSTnWWYoJHrASbY5A25HGiv6SoA5ctyi9ZGBZPJLhi6MgMwPia4dxB3id
4pMRX3nHgt3oLF+IfWHWuwFlWkXMNziIUgyua4Sl3q7uMrcgXjxi9DLfXq8VCVwobv25C13qNP9R
GZysXRbM49My5CATCx6OZ5UvbWjxnqMvNmi2zLfTXg+/aa06L0wH9Q33xA3MNcXkEOIaYNm1n3e/
sofjiFwGh2hP5EMC9/hm1MgHLQXRusgpNoP9BcFio+1ZsWfiUpv3PilfHMxAKPs4IMlitTDAnG9L
6wQycXd8nr70nyuUwBbrdeLvY8BLfThnZmgR5zbWRSPUTpoPurgJF9eh/Qpbz9sT5bZLMJql6XBF
5tO/rvOCTlDALttgcXwX7Onc+LxNQ2wFp8Y3sBK9nICei/a7WPVeGwqVL/c8ZDGAl7xwSLs7iJ4S
c5CNM+Ym+Qr7GSaAzt7euTnhPcvUFYFzSKE8E05/tp78Kqo1HUm8XUHQks5N6+oS81LJ7TYPl+Dm
esepCK2+6gOYSuPZQOTvjSH96AVbhhiLR8XSIV+F4LbYzSEplJN+N//K4r2qW3fP6p5W5pEhLK/G
JJT6KQfkjromIBwiZO+NlagkEwcEkBofDxavLjAWwPW9BI3Q6aJFgTraVlrUCq8J8AgPjj9PRgXC
lN3gDKAAEuUWl26c2JR27Mo6W1RJz/nS5NBgQj5Q6eCmkZvWIL6GWsHp+8ZY0RwuaqQoRrQxKJ47
1RkdQiF9u2A1BheALsZjPgsOnwRk7YMd+TfaPtekRfaZnKt6Tq6CU7YIbIsWAbI5VQQUP7LTttfv
lmFwYGH6wlyG1YuWb/TgeOF30XdCBXXSrQjAJpYn/q/wUDYIGSVzpXooE1m4dsnekiZmxO0v7QSI
lLKax+EloQVZfpUszhLqx2UrJjM3qqM2+qp4hCYHoIyvscE0apI3zChjNfKoYgbKc/WTcv69Op+U
+qyx8rObIkxSQfptIeJg3YhfrDBMrm4r9h2pPFcqDROOaLzE2bHe6qcpqnPSf6Ojn31QWeppZOJM
PhqRp5Cedt1w8dZZKwtTYt64LXDF6n/8SGWd1B0+ND/TeMHeHzrokVNzvkzrlk/EdWVwsS6qSNJ9
Sw32u7LX5KM/kWXtA9pBTh9StQS1kw+y/BTBJw8+u89rUMQ8nqEyKRAJ+gVG15NIbZfqHGHmA1oA
qUo6HB/EwgH+OhgQkXrS2Aoqz/gGsmf2rq3sTfIpQFG3Hn3SycCsK9CeGaexM3oNAL821gYFe4Ev
2Rz++HlwMdQb9LcmttyhTN4kSodrXY+wf6zZUm/3x3CdGoDEsTG/4vc4yF4ikAfeBDVX2ptO0fOx
mveW4YF2XGnbgZiiU4bmYsUXKAeCWItxOsRDIpyu1imgRWBg190n3iwA7MTRgwgmqPU9OpCzZDN1
Baaej5kDSVIPcPwGXkwD5yvT4+Hu1mSN5DDwUHPdhJscf04UCRBT01F7PiALMDViLHVzPY4JO2Bb
us8YEHW9KZON7H6Zc35Z3kplE7v/AD7/Y/8Ism2iured2fTC5UdsYVqzSBWqcXYaIXj+lZbbkodZ
b356VDi35sdhVCgN0NboQNGzgTcVK1fnP+Z5fSX9iQFH4KuYBPZDRNm1tM0vMOwMXcRL9M23ADZO
LbBvPbxevct4K8j1JvlOXjfm7BToaiUaC8hT4cFXUMqjMlpqtC98S5EPvXsqbnVsXvZ7r+pDFuNK
sIwmH+QRQIdigQpC0XpiYAuuwH4Gz8r1XVJvQphkPPKdxdmUe8i30Enw9DO0S/0Hnu8tAvO3xE/G
oa70ZqG0Ofmn1R1mqdOSaMk2IJetOf1EWDH8WXCUO8W/xwCklGrOLxg7jm0ZGCYxE8jqLV6dLCoN
xxWLuTtNTZekdU65M8Mh2zOPacQXet/pwi6bEYDpahOyyFy4/SDFywTlUtvpWen5OVj+lT4x/j0J
d8EMz470E5QSobKWkNFl1oxICAhy4ju0hauOsy640eGSsiQynvCKjRMz+yhFyBBZbBBXT0Iaf2n9
Ng5QnVY4Fe0IDrDBAJhYhJb3CoogSEgxaSBwTEEhzEDvv38tDRX+caWGgjREmvs6YSGGVrAaoMiI
ye5QiUcrY6Nc8WkpO75LEITocgcVHBoPf/qXwjweNmmtEheYsLIZ1TTXOgW38jbETptkx5U987X7
l7rIjyIxAtIeactXRtOes++mYVpY0qIi6QsPfxj/g8cGdhP73MGqpIGA2Wdi5mzbJYnCHptzFyI9
qdMuazxa4c9aqMHapOiGT+lRNktXF4NexcGy0zodc62Q8jen/rvGETpoEFhnw4elOwSWk5BEQbuD
4m/28iMd3T7gRyXCxa2g9EnrW4MULU3WIzybkadhNM9KM00cWWkYjdhgDc3VTUZ3kD25eIE8JehD
Df7gXZAJLgb39Lri04N3F+9MfElFiAvmpDLTVJxegl1PaUnxNifriTR40wkRcwgRUBAZoXN+fNUK
Q6OBQl7R4piutcp1Z5Uz7wrkmhgBFty5nDfgNZfd/X9hko8K8Q80/SJKsEaNtm++PCn/aT+tQLVT
6aWZAw8Z2FSywW6rPf6GQeVxYS92KFYX8hCTy7bE28lUv9YALKxjqjrEQruX9moIsMxdDeX54y89
Lvw8889lBMMIxyHU964+22GkP2Ap8cFlYUyaKf/2cVh6EZW4vctA18mGgmtkx+m//qMlwmLygQ2m
GPiYkWOh5QtJjwKGKk5E//7jW6q97dJ4x2tUJwAEd2/a+RetwZ/tbV9DSvAbyNjKDLHBKPaMxT/M
oA75CsyFzrM0EI8MJHKDuJzD8W1VlquWCal80/eOfwSvOJV3PqyLzylXHGA3GjYarN1SRkjRZzcF
M6SxWk7JhvKH6gwB2Wcel7Qcqwg0sCaELdb27VgguteDcsO0AhIOpg7DEFZplSLBO0gzGQEKW6KE
6FivSIPpIbXAnKbs03iwkJJu6sP7nXSMF76/xKjlHcQyCm41EVM5Qy1c4dUmWFr5s7k4bc4KaUbi
Aem7Ib2KfogmghPDK0M6Oi1eOfX7uT3a3XrfC0YYL64dPcsaPZNhi+UVaTLtqgQV7vwmBktdG7LA
H1imO4/QrJSzfII4oaZjdGDv2uFDCqx3YcHa24X3vY5Q9VkYCniHZT+GeiER3d37jupK+bhpfV6B
BZXZg6W4oq5SX1bnMSItlfAK0ENpzpj7BQ9roW6xYCUuQ0eE02U2DZiKF1ooioG6SsP0tJwxZPBE
UT9b+xp4rLMk1HipGZMC3jQL6QZ1RV8gk/GJOQdXzamuAUkhqxrSqi1bX8z1ew2+BGSFKlCJLKna
Pcpb5ZUq4Q9m9mydhCVUTpS60LPDlgh4/rcNPm8t3iJsnN86D5pV1Yz8y+9FhJCtWqYbKyc2rV9N
5k4O1/eQf6G2YbT9sZns7Q6tb0dzpuatTHxQwLGrn/daN2T1I/W00l1MI2nmzlNyKG6qWMVEmYrM
qIZJ2SiqZENwZUwzGkCh3IU3iBViMxaY/fpL5RHVeVQhfbMM9waUtnPK2EP6QrpM4jgQgaGx2sEF
RnOz8TET6mfBi+Xs1F/UHtMT70+CFzE92iu/KyOPFEkFiCqL1fI5u13bAMIeyGjUMn0IkNlgLR2U
LZzEj1YpglPztCjzCtvZr4TsuuXU29kJpQW2qg2b5PPRqihDK1NaP9VXO9L0o80jeXvNxY6s1p3F
P7dl8K71QHnzbBRBw8CwcIwtk9Yjid8NShWzucu2XYrOEOA/sXsvKJmfIsY6q4+pR+rI5yrBCRMN
J3KLyaT2gE2193myfqJIpWqn7qFwiVKxfJCjNIEudmZLo2TDPvVH3nIC5SBoNlt//dZo6DBOEADC
Z163nHUrxyJjDdAHdGujIiHZvS5lgJRpxL4iAhaT/E63e1x36Fb+ai8LiWg385z6VV540fcD9E5o
a0ZfoC9n78OYAkhTCyqhhUcslWJMJ6mCU7/6UCLfdw526vA+U8QtbY2FV1Jx4TS6KeYPpFanGZ/a
sB3yjR2USdxp7Ho0oz+X5POibyPeFevT2v3vP96+qWl+MfME8NA1CGABFTsrrcJ+rNmtxIAne6VH
3Pp1Rl3ETJ0sgatm7uMimwU3HpEn725NktfmecGWZ5lT7IEgDpzbCuVzE9qptvWbb+hGydpjB4rv
4T+rv2JyPNmgO9V7ELcc8xRlWEghNY/1+6cJEvkC4ZYP75utZWY+E+ShzcLQqj5AEP5O9BTBdOXa
CAFhEN3EKzMiuAquiWYvduiQXZEDLNYnLSVgwKpDYeNfjHhHuUeBbYxy6zdpRKj0dcD/GBhhYa9f
AdvB3XANtU3fJQSz+b7rHWfvuy23R0G7z8R27t7SEkSva6cN6+JeR7F5e+m8Aw+yBNUVErkrQrOc
pskwlTXffzQwoXK7SenVvz76IjdfvzQzP1NhkoGmUQ+5iQeeWVbNjqUuzMkRtTOzohCkAemrE0Gj
I+wsAJNeWAnKJl/7zDrZpW/MDo9IkKVXlCmB9WPkJCFDA3VSMhhLYeLLxDSXwHNJE7MXlft82dF1
XAwU/LRvmiztgzJA5DPNo00hStipPTelTFR+v4MTbpGhStiloa6e5esWMY8mMvp2Q3rw7RSMO9OJ
yuIaEXiyMmk0kau+cWaLU2+N2gVz+r6SWfudh1AH/EsBSp2IBIEvMF5CUVj0LAqYLpp7TENhdTlD
3wjEk7v3K+UVyagg/jrcMt8k2Iy8ELoPqsJERSrgtpD7dmxyQrnVtak9S6Zed6F4/E5rzgkoPq+t
78SK7tX6goENA/wGd0CgYe5PrribkuyP9QT+t9/ZvM09UQkmQqE9FJyzHi3fG1FbQiGxY5o4wx7Q
dGSUmxsf0XtGp2tTFe8kPnbV095qZzaPQxDKBAwsXizeO8AmtZYZttNE12OLuxy2zuGEMZi2nzfN
VMPyt9CwGhxpIor7uhSu2zZ9Mcc0Yal4tOjPYP6nB3Y=
`protect end_protected

