

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Ksr82/EJdyTi/ZnocplaChIHl5gVfg/QywOs6WHQUUTVobYB9S2t7HfNHkvfksORtftr4wgSGG59
dqflxrTk9g==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Qqej7lC/8l20xFx7bklclhPhbKpE2SoVMnU8o5jHyjJozBFHGWWzSqcy2OHoxuRC4svtWcuXPZER
AveySsBsquyvS3CpwUhQC4HU879mrvq1rktu6YiGUKekxqqq8XWVjGU2RErpRUag/ydvNbNrFWxX
vuxu46YvGNDVpOq465c=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
439mpd6b2KugK1Dxw8VAcq35Q01RTqPVrzIbAJdjxQbya32eEZ7i4WNiFuVZ/MAk52bZBtBQiNHc
mNfbIfQciIHmnAXJEN9w/4VODhRIcUMrMjQwAjn4teKfB1tg762rR2jvGQ50Ai1Ml+OYADsAGJtF
URFceTs0yqpLMxJ8Ov/lGmeNw5dXmLiwn/XRqtS/K35VTjZyDUeHpQAr9q51KY6k59LrSFC7lxxB
mXX0In+fzXXlrh0dFFwLWzscDXHiKjrU4bwWBuzmrkKr3uCoEG0OADwjka6wlXo/Z2cEkTpiK1Qy
MmZH9UXQxrxTgtpOMmK0pjs+MfXf5/7XzeJsOg==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
porEUqarzWQ+a43o1KcgcLOOq13cwiYUyYcVmnYhbdWCiVlWWfN80U7oRzW3NODV8vTOFdEeX0/T
HiPsKQYOSEqQjf71FVXt5Qu85a7gangJ+zMjyuk8+m1c85rFqWapoLbPUbexfLeiEmybpwcybBzj
rIVwXl1qRv1R4JNRI44=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
s6/C7NZuQyYs48nVSWrZBvdUw/cGGwVNCnxc6+Wr+hB+GSdh07xJnxht3+mpM71wbe2jyi3JRq7M
A8Qq9KlqvpjZ87ZnAxTvr8P4OZV0DRnim60u79JqHUDowRtwBKuWK+fhBBqVkg+I/GuK0CQAje2N
3H5CzXagxYQGmhNBvdIDYAmWiG6ymENT9OP+fdf/JngSq3sbaQDhuOCrSGCgAWuZWv28vEMvXd4d
VKm66HgH4TXtJpDsYN5kTW6gEWdi7cV3KJRDsY6jA9RzwyOOBsMl8Gl/UvSGBWbIshxBeydyVUyg
0jabYqp6ODPXSowz5ZkW1y4reTS+cozycJAuMQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 11008)
`protect data_block
xKn7NvrfVoUly1DIs894j29k0BUKCWTY5pGCoYYy76PcnT8BlNx8JNn724i66DlZM1ykDJ7P5oOE
QUEV4wb68hyW16hDATK9/NXFKKSKgRtE62PzV6ofpTtyfCq3dGZUDXGFg00UFFuv7ALZHSpM/ygI
cXhcXr7jPKiFeK5eiueuvJtlc2PReBYC4uamieb19YWlnk+jW5YXieIj56J+xIl0vF4m5BfT9PQq
OU76XLzv6MNQN2Zx8HnnJTw0GcOO83oekmRBNrr/OLHf5kLy7folxX9QfheXgpdhk1D5uHXxaGzr
AYZn51sicjjEzxSDdofCzMIvskfGStKYg/FXDGqKDBrJgcR3Uu097jOVnnwW23HXfDSXmJ7Kz0vd
HKRlLTVYDQ3/A4nnVTTEzPmW94Z/FK6D3vBYhG68acC/xMvvLw9TBvbrZc/6bVPbddlddmbAYu64
j37U6fHjW1DMyhfPB/0ybiNZyi77VbdZtJOSLXznec/fm6LX+GTybi+oa6Gx6ZJbQtr+lMxqNeCk
6i+XAJRnL0TNmrE83FYKJhODwjJLyHKGGStshTo5/a7bNGH6OHX/ElQxhxaHNHA49H1BbJzm19tT
Szc+KAzB4pH1vwsMcgEuG4Wo2A+tIDamKaPfz2X4kDGfHSFnR7axvvs5Ul873vhm/ev+xGVoAQxU
ZYauRuk9ITsuvaLUBf59S+qutAsaP4Ch8lCsU8wrrPGKqWkqA0OhU++i+kzdyicGDeB4MgeLaS5+
K9BEfidKY1QAUMUeT40a6GFDzQlJs8f/btE9hAElVjwU//7lKlRQ8sOT4BRRDFq1O46ArtRNvp5P
/NtvINmMbgLLNdkolF7T9gjDWaDCpPUdsWK5iPfa5ejehW0IdkG32nNDx0DLJcBNLqWPGasOGYDW
Z7i1xGOAKcAu7Vai+1IAgiP1/C4oGV7EPb+mNAWvHW4fmJHWBVmfhF1z+3mkbFdeLQzdOa+R736q
qGeP62lRnBKN7rZ6fY15t1bQlgTdi3FNbT2lNyUZkRH80tGisNpsVM8x+GM035bPwvd0bSefkLDG
hffz7TzLRltxobmY99rc94MJfzwsJ6a6ZoU944vhM5R81qB0JQJPLeNZ/4v844Qc/rQejpiQkrj0
Z9qoOXohRzKawxgfnFyBxtA92lBM3UAxekDm3AVcSUoMhRXE7QoBulDgZ3/XUdJapdi4/F0Hq2wV
JTqIIxgcezMvmKILxPVWbC0HW2NgIdhwCt2prNJ/mY4QnfaNKQsnKIRV5cZTdZuEQCb4VOHqS5Qp
IQqgbUE09vTfQkiP9w2bq6SA55QyXjo3KwRBqkZyFZs80SvfItLM1nksDM3dtuSew22wsVvQEnTx
oQtMzk1iBSGUoz8CMdH2sJ6yZRocQxGNpLp2tBZuBuz2obqk45V9KM9ztKKt1HDSGZ8Z1RnHLOKF
nNrgfXY+oA16A8LoIyE+Fjpfx1vne47CnVDx1IIUogdzm7mk3a1s9/Fb82utttKMTC3hc1tnuSDA
iPyjAxXcB6WwQMkEzH1aFw37g2wIh51o4cAhBzJDnfhqvRdG/3g2B/SRU0o/wCdvCx7raKkyHGxS
K8BIvZ9KxcTtj3LsTeo1yZYcEYKdvkr/Fxi27yIzENwMU/02jfxIXKSnlg0ZZvCHve/YhuDFceFi
NRr/GkRXSCQ14lEIYVFkPRpZePRW8q7fPRm/4VTfxt1WrDQMAJUdxSJCt9k4gWW43cEavgV5y6N3
chOeEjkWIUJ1bNq/JPYVDNklojzinOTuFKFhbubeEhQzJjWFu64eUtpMYw8yyyObyPcnsn8xMbub
rgC6eItTzp4AFGBSc41KuEaXYgjE12W/lNiFyOtLDNcSmqY0OA91VQm71UGlsO7oELp4JypZTGZU
WlJ/J8q93XLM3pTrFd0j1XZekCYlAnC+CGjYdVP9XhP/FoqBl2JTrJOOEhr4Qvrd+zXeesPo4We3
b5RwpmRykrIG+Izg5tkViZOmAyDyR02ObOcDPSRTK9DEeNG2beEvIa9d0NyKar0Izn6LuJnRQ/NN
ed1npEFOB0FsbuJ+EnAXF34qpJSxdGYQICj8ZPo3JOmOgn2JuvGL9cICc3h/J7Tnk3FEoVux51Ro
GlkCMDJVk1SGsJfgFtxyUTwHCgnVQBTAiWgimIb/1iStqCZRDKKFgaytD/PlId3oBdUxaC7dCAN1
grVK77ov9GnE0Tl8e1PQD/gcwm81mI4A2XMa7WGxx+WifDxWmkBWjvry92MjTe76jl9Sf4sKd7GX
Z57qRQHy0e0udtgNq9o2UzHtSp4HooP2UdmLw6fztuQeyrVlmdxFNElWfe/vIw9ngiB299Jia2/F
FkKBhx7d29N8AV9HtvpYJWO6LcRJ/Ns0SIcz9hlqVkuMzVAsyIk1iyaJo58FZi8YuwRjAoNd/6Bv
QujtR5zGz4m0gfjW5EetcrLXLMQe36cjTLTIW3uuAk1YJdBlFvdAZi69kaaYpDLKpd1LPgqAXzsn
SCqCS6OWNZ9RlRSme/aQnBh4hYtDTnQDK5cQDvG8aTbyFOKu0Znj8xv2NylSUq9BhrGnBnEAhBHa
eGYBRicBdfZJFllukHTKgEZWuHmlRjEy71HKhxOpVBBMeQkcksnSQkFNsDMLaC1gxe11Ha4FL7Q1
QzMiECyrkyLAF4jc0bniUZIjlghKv2FnMMfqmrn24+pkRRay0ds1zd7rLcstDHypxc1+WZPvnhaH
SfSRfcSVTWz00RAOZWC+NPZro5MRzmHi1nTX9uMCqH7FM9FbgrV8FpqWQknZJX8jU9jC10gn1ZQV
8BHrzVd4YBXkPz26bozCu4cUX0orlMiTbFTfqDSa+pB0rF/0PUY7qK1lyyel0r9uMrIO2/b9Uko1
BId9ciz+gFV2bbtk5E9AFfIB7733uqzaAp9pPXOxh0B1E0QYpWkKiHVdEJsXgei4o5YnR2nkTMrs
WBoQ3VgWO+nuSwVQbKuUcnHkfRx4vpa97aEL+/PhH11GZw11M5Af9djwAITfxxGEamo6KVa4wvP4
7oRJdDXvwLN+XkJLvO7jpjgFrNa5E3AwwQF69XwbfwHKt8z8Bm2uf3pQ21P8SfSWSsHECQ2YeNjb
l57yWSx75wNn0J1N7wDOLsllznu0o5iapEhPOd8xdOtLUXoT6hRbDV1mPejJx030IcM3P/EzG1/v
Efqgu4xo5yevSXxtcqPOHKyOI2ErdHrg4iPCqjeHYQaoN0Y7fUIoSu/JLga7t8+VWcjGd5zBtcKi
U4vPts4ItHukaMX/s7DLzhoaLcSG/ICvvq25/4Gr31lI4grauR9ubgULIYURLOVEKl9+pHdQFj+u
2tcvaxgfIVfaDyugo1YrdJxYfTHX5d6hPaHpEBOyLd2TWfVYrFK9Ak+PRCnn41jEmqk+M4FZ5fku
5aSagz6Tj76+PWR2ZZB/Bz1g1ashinkEy60NWiCAQfgrve12sAYup2xRAHVJyeJh90m4a193pz6+
1TaGPP9TD7ZsFLdOPe8kfxfFJhNWL6FWDN1i4+ZUMvUBQOiaW2Zk5ig1ZryOy+TJOdNb3RpuOMMA
q1mGxKahw3iHvKsfr3cEuhREdy+iuccLTnAfcGfsFwQFFh54dJNCRsWK19a7Ix/bvclCUQVRnsJo
USjHid9LQxQUiw5MxWw/9iXffQ7loaUFsBaLpZmgvX/la65kgeSMQJvBNX8ZpWCUNUeF5QtaUg/1
BdVFRZk4g8d4zIMQvSnFzV58jqdhdOyYnGwe2HWHBNa+XoH4w1G3+5sCp1SlxfXwzjTrWxxnt6zs
jgyOGs70DR8ZbKj6LwCZYxC3qtSH/nLiOXKkI9EbdI5rOorcbvmnbPpJ254YXKhHIjfgnmGXtInK
vqgZhj4octUdp4WqFtxYa6szBeLHR6Xs1QgTwkAjrNwZ3Icd1eS2K0Vt47j6tZuts9d7NzCMG7SJ
F0koLmpqXig46uw/7UCeuRKhoN/N6iaYEM+GvkQq1t85zNpJSxCGu/vPP8sl6xwLKaxP3eb24Avh
xjW+FhEL7zdOB9muzG8Gp2pW0RCiR0J7Mw3TlUr856GpJaHmqDK1pAKo8/jwoboU1evS7BZDP8k1
DbndPUKdPR7xT2Zfq3Bt9UMoqrPLfVrf/vEWLfJapEsJ10GmRi2+tlqSQj8lsrzPpwm0F+9ueoQj
hNgIibuclCZixHMHbKKh8W/yiJEwl4iCS7nT3MBWZFl5Q2bFYxuSncIjpYv8CoY0HhCAUnNWki7B
ZO5a3kUa+gd+C3f07e6TgeMbdVUeJTPX8lO21lh3YCdJo53zNv+wRUsjH4O2ZcE3EC0oFM6HYZgg
R+9aJHv9i+CsBzhOlIg1Pe/iZonIF5OmEzX8/Z4uYU7ATh9oaF9tA1a4lVqhtoeFu1u4euFw7QB2
Q1c9dZt0Of6sFgFbn00NPivuhTnz/PILrqzjHyqJGJdTWcq2oSv33+204sqqzjeeLUjcn8Ygwnxk
q8SQ6GH2YrLbhGVlv2uja2vDQvetrkeaGrblfB3ChOJGinKkqGlmDsePvh/zTSnUE558TJ9KHADU
q3Gp8iOwPlRnoJoY7cFr1xPDicCFq9i8a+FXpjc5n6NdSsQe99M+HjzAWXycwgUQTefBHTdnhMSt
Nc6UlAiQ60diXf7tdALjb9NJpRE9YoV+NVCkN0nJctu8CUfWtm5hyCxF696d5DQNlU+YjsWCCrkO
FfyZBgjrU4szkRyk4QCxATAKsX9+2dODgAKVL404VX4yJJy8rsYiWi8rs4Rsmnh6iqN5tzYwMYmZ
b1vHMAZrirXzB143OGuyHHPpeKhR/Yj3MCJMJ0T+nKen6UEK1j36EUVBiXp5SnauM3b4W7QOw2Ou
991q25k/9pUK3zpy4sczsGruolI1A+vlbOotdmnV/JoflzX9NSdxswKlv/3l5vX+6Zo6IqlaN1Ip
rHj+fyp6Gh1UxbGfyrPiazef8VyOzoCBmntIrcyvB019Gtw9O9Agcmois4Tp2AHmYR03Q5TlyPOu
jrdi7hrw0uYPI7my7wpGZ7VtlSDydpk4RKMYLTqybICcAIboh7IMOfuHb/nqw6el0+ZlYTzZLEim
oVGvYmn6OzAbxLWwYwQzNQ+G9/XtUBENHrlCn+/1vfF8ELtZXKarXqHM8dK82OpIlz5wmlboZmuh
HmCaaFeGikWFP4NkQ3i1PO8ih3SB9/RdoQuogm5qj+xTuLZeyevk24uAkCy/RM/9ZEqZOZFrJaJY
toc9MN8FhUA/wbW6BBIw1aNos00wc/rXTrChjSlBPhEF9XHPtINjuyU7Da89CNeZZOzI+yf4447x
I2beMkB8X2nk4l5wAvOAUJdSC37olVnOGuXxiMnrI4kwT7qS2BZ3L0ktYuQiL94M+5VZthqzl2VL
k0S7+N58m4k+zL0MCwFAXHfDGtHOH4o73hVBUNXk85rPuW4Wd7duV5aOTbVhyGJxq48EKwAVHK6/
ID7FSp4fo7L6bF/FNnfIU8mQnn8W+NFeIehVNK/AuMD1IihmGb3fuhZV6aUnkzveBT+46ARaU9UX
zbpjyIt0UZo7CwEsEmN9uSX7FBEydlMfPWGN2jxrkmuba+0hceIJJZHXUbAfx30bm4NI0pYJr4hK
/PPpQRRAsTCKDXa1iq8GDGBRH38P+k8bNtyLxqira+HfFlVjPcS8wOR4y7v+c5Q4TfXAspvi9bbh
lZGUy3ez4FHaVM42kLwLdhVXxloaLj8PM6J58vDdB9SPZNkw7/9U/1G4s+Ug93/6Ayg5Ov263Q7F
cIWIrPLMegyMO0znT++1FOxmVfsd8QKSeb4N/zb/P0MgLEpU5f1Ko6+LTr7QIJoBwqQr/re9jRQ9
nvJCGRCAOkf7BoJKgWvO4PinnpCC5qjVOtkj5AEBI7n2AhnvNuBTEp8Ms7scGErnjHwfKURMW3rT
G/joROXU867tnjlenF49lmWzoC2+Romjuodojp5MTv/unSpZCRkKCkrbGo6I4AG0PqxeQxruO3gi
4aDHxG7KeaSurl4Wp6PNWyQ+BqmhyKQm3fV/gVbkwev+nCz0nEDO/FuPoufe+h525bKq5okDQ6Mp
YZItfxW/onP9CjZTKZ3AKx8iQChsiLrLr+bsaCXfkherDA9di3NTztfJl8kRqPHsLxMtwsyfb0PP
/jbQPacClpMdKr+D9ASTLL7/uUG3Nm7745SDfGpQkWU8YkNOyCbHWFnvFgUvo4IuTGG+fUuwm0T+
ayrqgfyMTzUH+R9jOHboM483gY2MNnuxMxED8xki1q3frxgt6EZBB0TDi8+j9D2cWEO2ZflUAX1p
yK2/TOm5DSkXylXh1m9c7DNn0TeV4kgnFE5SYWJCaDcPOvPK+r/xmrF5tplYSaQX1+o55RfELo14
Vp518VgNHh9CjTd4ygRZfW3D1hNBOcbJrIkk/5mWKfRbLxDFwqUNrRk9l9ekRhtypmk5MHfgDZST
Vl9kucMACA4R/JgAolVVuRHPOquvh9YK3Go7B/i15vgReEppYuevtQqAx2UxvhebTGKbHxbvirhM
dL3IAVfnzorah6nfBSZ5zJeJangsQeay7t2Kl86/9sjIaHH417gakHr000ViLVDAQQrBeExWen61
kGEj5IJ4MU0LgwD9/zY3T/diyj8HtcQSPhgS9GLgD7HTKCjzXO0bITYoCIHDPjUWXijq78J52mhg
qrE//hYrGR5q/2PYF8wtXO2RGBInPZsmkD9szxquvARTWqstFUE3jnhqnmCRNqbYsqS+zZtEw6hl
k4L90IOEqhUnFxQp/EsvYy7JAowHS2dR40btZRUGevfE+pg97mF76uDIrSkllTFXWIApf0L3Z1e6
auT7yjXv6JDG24zrxTiE56yinb+QxeoOVRGfaunecQSc3Rue4OQLa2vjV8h3etK45GfbmML760Ti
t/lWJ93mJXk/dop73MBZVhPrAqJjkfUpolJ9H2QFO9Q2eGIIbqaJ+JOA8D615MTvM8DWFXL4LSYf
QdCuodqSy3Q/MuTLUTGltC0hae1RfockBEdqqcc50VFk+67aHjurdgzz4aYZqQh8Yn/PQceQZXu7
VzU2Jza/C3SKt2hr8lyOWRPoUvOryNZ5PjyjKj94OjOdiSDTh7wWPOW2KGTAtpUz2FNjA23NwQHq
ltLJ3yI6sT4fnPtXPRdxrofg1n9XsogaEjYThNzi+gDp1oH0rWiojK7m78JSrW6D+8AfzGohYcx+
T/7EiH/McSpnSg71lLf2zKctoN06jdC3NTq38bO2lcJaI91y0LSkXcB6i4ixyIgNR8GWe0eEiPpF
GNReBXH2Qj784oL/jAYfxxyFLuBN6jxcEuLaxxuNh/6FTniK1oB8KKM0tpjTUt1jDuyGIgvRIhWL
ViN2m7/knl7waR5P00GxU8+lMmEKNf/sRCaqwpBQu/Ug89IQvHNnBvdY1hEMVas0Xs2b5tbAsRBy
OuKAW7+pY0SFX/KoWb1rep7tNagWbC7e3TWp99zxRCYy6hUaFuyh0d/MYRPLShGWqyLq9XSJRWJI
SQQL6LlwFRCFpPaIH0hZArjran/7fxYbIi60xLMUamOoyfJymsqMC/ZkrfxBGGwiK3i9eM3IoEFd
3xRoKcmXRlN2LhgMT8UPXrhkcvMXyqdajaz/g6nNS0I7tPSb7pF7iyyEnmbrd2FAClXpreQdQP9l
5iHUbVzeLqVVKLBIg8+T/r3wloTcnoRD7CDpiFq3K9s6tS1EJjfPulQy83KJ98lM2ieLNF3GfdRu
XmiH1lhOZss2TBHHNiInRauW+mSSKT2y1aDw6Y3VZuxqFkrhWshgjj+TPk+2a0ZsCJenQUL81aVR
Y2BhrPBxjdJpNkCN1EDqAslavtaNjeTWqGHJvJU9enDyPStp8I58TKlwz0k8Yn2ernIn1WN/KUn2
y4AU+spGq5NDxRM5kN3fmSC3FfTQieemymllWAcF8BgLeCkCyAScmebtTP2Ih7b0iSCiWYfoYtw3
iJgoT1O2ijCwADECVoMiyreBHFjWA5+/BjnoQOniMSDZmYTwXSC0TB4WRmGe+Agd3mm39ksS5LGf
EvDNyBpLJdRAGHGHHvaYOWU9DHNL9jY0HMJGfj7am1tPh8AbqEOOK85cg642ps+FaLhZxaAlBos1
Qq2PRwSpGHiLYrXf+mG0GDkUyg9xrX4S1SZ5ljvPvBeFd6a2Glpfrum8bkxBoKbxXo23rLl4eNXT
HjCcxUBM9bb2y3AD5sezsZkwX+oNRFbWNzGOr7v6gI7PKtKgFT5luBeQiayLriS4kdflv6JH9YA4
daHBBEu0aTPrIytbJ0klwDU2iWz6pCEgZblmD99sezfArs6gYtC0QabiIMV7zmx0OUuJnOUvIfjz
SPxI+S//se4rOmVquzYbQ0o/z6b5kuuJp2PlYgfDL+tBdJO1n9akpK42cqfBp9350gu+wCEPw2iv
iqPW7gPhasxT+bPUwOHzRjv1Tdic0c2m3WP1j0LpzpO0P6BT6hbQVEqT0pYqsFxZr0pqwo8P/Me9
YURmExvAF420Hno/kYc5mIxlizjfXdOJWSPmTKDn/M0TnTFYPwFJif6lDT9Pob4QzH5JTqZhEPHM
L3soPJ6shQChjRR39+lNVa1es+NZyewxtLCA+cq76IgUOcQ52wVulf9AtxKaNqeKtqKRueC/wx32
wq294LCoMWIX91HxV1ZyA1j7x9hQI6odX7F5bHdXm6sV6AZpy+JLJ0sivSCDnpBwWHnZGpgR1fSn
S8f3yJbONR1cIXiuQHyifjESJ0eWdgrCV2XF0VEebSWuH0mY8Ds9QAGA0TnTr3gM1/DltRGD3MK+
8CjMBBaGKlq8WjEjNyapxkOiE8wJ/R4ZGyxjw6hloKyV/2Lw38U3dhClcJLM/yv6SOzZF79A17ul
wZepiod0rWadqMY7C/cbzgAIhQWtTlVzB3h8CguD+WYdgMjqL69GYTpsbGY+kgQT2oeJR3UaiiXQ
tpcQuU++A9q1Sv1S7b94LeJ+b+jjlB8x05JvIXREazFhVAnN5RZcY6wL+mBV/eaRUHSrPQngm8hz
FBB1/HLO99dVLaILroKAQlaHbj32QMObnmBRkQOHeWQLKRwbxI/azjyqiDOLDOeMjUQXOw2Zy+Xf
N5OcW3+J2YtmYyjfVPfO3vPMcQ15eDpD2tv+SIdXjOe0nRKh7rzVvWiWH5gkFt3Q+2KzLPu054Hg
3ZsvXM2+bp8pDyCuvMTRjcacFML/U4E/LxiFwS2KcJtHFn4QJ/25AkX1D3fBu32az2A7XfDpXX5z
oqAjkI8rxECVba+KEkfezke3jyMj1PB8oXkCcVvQjtUnKMUlcFOhBE+46nqn3m/1R81ro03dAem5
sCn/vUGwSNqX89bl+2MxYiLQ5uieuBKfxnGaSn6Zz/aL4esywZkKg4FwcI1MHZie7MZqlUsazK1N
gl3ulUtaMBxcMDjcdVw2Gn1+P+1PzUCYWnEqHebiM/8FQW+JrbbAkKMjUURUCEaS6gwywlAg/+Ae
5LhpbTiULdo38BcJlRknnPM6mMc6Tdy+TIcJPn2ufT/4IlEcORmXlaHPrhUgDgU5m5vXgBHKb9xJ
Ec6gIC/YB2RNNK3HEvAPsbKuiPeuj174Rt1i88ESQ14JVn+jfLnenD/6SZm9OjdO3riYgr3nT3LX
BPRFkECHmznFwfBTC7HWIKyI1onpCjXXXyiOueRQ6OoJdtEGrHabw6yCOKR5XLDhlja10tDJMcYP
jidxW7GnCmwFZPa8yRf+qA6RhO7pGqnHAotb3JJ7t1bdnDvmWrkADrtf6kJx6JPU7ovvCyXHAiBo
4agysyVyqFPnVvUPFimgG/Gp5uLqbBufAHqcF7k4joboKHw6i9FVpcyR5fKVb8Q/gPvAL52vcd0U
7HY9yObF7s0DIrpUymrdO3C6ADYvYcJip+kH7sXYEs/EXKCIj5WRqJ0t8mIBy5qc9IMJjKfdOgeY
CPhKIkEF5kmA38H5ghgFFZ4k3wqF9MfVsrI8hJ1/ciEN6Nj5ZOOBZ/jI5kdt1WeLg2sm5k/0/mzR
zHnMfz86DtBsfTpbw3D2Qunmr5A/u/csyBrxcePYhqHKIqdj/HJWaI8ZQNsalDmxvEUM+O7oiLb/
vkWfysWf40/K6hjB7o0L1wRn5mrGqGrsAVvVaX26B+YwKeHDIzl8bXBdE6bPo7kWK4GTBlzO2y2y
z5GdM3ntfc380q3FOmoezCMAGe7DlJ/D5H27mAIcsDQChO/6tcd/cJlGLOhK1u3LGr3QlbTq+pty
RE//xWUyx3mzzBiCljaPePDLOXN/6tCAKcRcLemKJkG8EOYb9uvXnMa35x9Ura93nhKP2jCUjmry
FlKdQFF1qMGloSchKQ4Ne73y4QGL7WP9PVXnOLvIRmIO6x5pTU9jY/c1pdejQ0qLcpXJZ7hF7sKi
+xZQM9djJYhDR3MGey+/hZLDJWfOo2z9ylKtdT0+cP7EkBEV35zLEYxSaRgE8JDeBfjixLnXNSzT
JBmpkAdCBwkOCHXeVpgTDIO2DBIBTsTkbI0BN+7x9o/NbVGchvWllA/lU9ipkl1iF9JzGH1JWclu
WbdRg5EnL0gnVFHvTtq3okfrT/J0IununL02om9+W+CkMSD51YP/NoDFpyHLgQj00svkd8ayKlc8
gaiCDsQ4HLeX0eMrBBWtv+KwjKWd/XeFxFhWOErMvj+Jm98ZgSKz9WStj6Ya4PpmD+ME+juQOeXI
irCXG76MYsSDPCt2qUhf4bOa/5CpyBSBRn/4YyHMBPm2Co1oQ5zdJN2VGs2A5brxIgcNVyt1jjSu
nX8UzbXO7SiFTexzZGnNmeltKblSSEeum1N8vwnCiBMe5FCkOh9e/wZJv6eMDeFHnjcbFCP7p3fF
azt+R+hMxwOt2f98f/LLTx+jL+cFbPJ0yQAyMaG8k0daFxMwy5jkRzgR2w1Kc8hkDAXSoRr4hifH
JHLvn9sDete6VrpGJul86ZedJtO6uuXKhEhZLcDAcfOpVG80oCCFWZUDv8y+FiMHq6gR2GGvS7CF
x1xg1bm6CoNnP+s8SkPEs7w378mn6JXKgwnDqiug31rn4jbwEdvzHl1ZFOFQ5bZin1IEmozfjm+2
We+F8EZdxAPMwyWaBO/bk+Ce2MfU3iF8cQyT20GIVKgG2SNwHJIOplJM+rx3iT7rgWMrvbEvhwcW
Cq8gDE2Qwe0t9G5g5qgXpoP4rQbZ8COkFlM5HBms9sagRLCl5n31CHX/GiBi9j436ILdz1UCUIAJ
u2jw6sJJXZNpargynjH72uN0JmYzHHbfyBSmozggdEENgMGohmMXaOMZIKl0zOB51SIKYHeWfSiD
5d1BiZjz6lvqSqMBJofdQQkzS/NHaxd+wrCe64QoTYNNBrK9yGFKgnBWx1eheZZgjNmTZzafTKYn
Hr1ssQt7X7v2GMS4Kz5JfZvxREk5lourIXpzx+PykDnqb57nbT6+zUXpRhia21fWmpYbEmShlhaS
RA1BWUtRQaxJ2NgHYqmCuRLoGdK3qmqbYmGt/sWaFkmCRra4tJaHbwcy5sEww3PYRrWCxYPexhQY
gy1cPf/fw9LTW9tmCMccUuwUVj25/gjecdgHk7Tzu2TAT9zW4s8Zd8PTQq8ODRLyOvZ1xIxiHwhY
nDfoJNtxlL6shayEjqks4bTOxt+GaGJ9FxpXRvo2Do7rLN/cR10sTPHOX4muytAupIaVcaez4GBD
2YdI4PmuXgu7hgH1k8Wi0niZDrsz55C+SYXa23v3qxJxBHPKxVkU00BnNeV8WcuBNgdtnoZmSn1o
cIBr3OPbrpcAUZ53ZeX3mEJh6hza9VITvB00NttwWjDs3mXTai1R1EL5U2DNHA78IFDicX/9tAtJ
H31Kbjko6ajVL++8gnwc5vtimzhn1LdH/whoft/eFVONzzlsxbinfJV1Si9ZqILE1t5gb2z/H6gi
AYw5g8N7s06g3q86JcTk7IDEL1DE2d5NfpfrcmePgkr9NSZe8+ezWgAV0FlBaS4xTWDLFipMEqxN
zmUCklpiYBoYU3Da/UnOYnOdWCHOfAZOZE7ZlaGhGkHe05B+jhmLIeoUVV/ADHdBkjQU0hjHpavm
5dA2xPmrfdIuaAWFe2ggowYgjMRV/LNQNgmJYps0xfjywm24owMVqKohti3llhZVqrbFf6QurYsA
8clFMv4gcZkWQXPvQUUMkeuimqe8DuTF7hG5jM7nlvm/yE1Wu0fRaeq2D8Pzk5sHYerpXoDnCN/f
JuKV/csKDGkiQp8EfFe6U+P6QFduaLQlTBzMuOmaUagb3mDpwfzJVpdJvgATVkrMiUIXhItI/PFZ
Qw8GDjIiGy/Y1s9KcMCgnHa4PYfVor1nC4wQRV0e4oNcnO8DPHHrQFJaX0a0waPsaU8e0GEDcNr2
6XHQY0DsjMaj89RwQWg3CRdG+uFyk6ndoAJlUk19f9BrbJNnQAcsoLfNMBviO6BLz3YnCCQRApRe
4XaAT4DZPF/fk2V26nsbK3DfpwkOUST2Bt3aLenuSEV+oLvA3adHPdQyYLbxCh8Ar93PB/fjcMl4
UG+YW8zsA2brU4DghiCRrTnQHmmhowtuSIhaHK/btKL0hVxCWwA3L+gGTgZVmnSj+UjmskKRxFEu
jq/d6+fgs6k0XNhkTKpFdCsA0k38lqZZet97aqwseIIKchQuncHRBdXBc/gSqRLcsF3K0EXNebpc
oC1sb6sMydYkjGy/kMpVWi1wbN9SXaAZIz+3OfOt0SQfq/pqkl37E0TzGeDcL/0pHzBrYgD/s+5n
xKd4unD2YmyI38ngkia2IqzBlGVFaQieNtZJm0fTB8yt7mziZz6UNEt6cKJnGf7A0+p2eHiMF5rv
1gwKuq6PGAVlfHx1mxojS1CuUMXtA38lPpycskleQQo6NQLjDTnRsLKr+10B2vaDTGgHK1HSJdzC
hTd0NdxwiH1IiHyTjY0Dcqro/URMPdLQjXij8BiZ/+v78oahWdxFSMOpBCOSIV9HCfvB7pWc7xki
e4auh70Yn7btZWHYo6wYy/4aEt4wbOD51cZNfd0TNhecbFtc4q3wvE+3Ki2HOy6iXMiYUvo0BpaX
qRw0Ry64wHP8ohcoXBqvcFUxaNs4bjjltRitg/jSbEeNyTMuceKifupgflbjm9qG+BEXv0YXxGUD
2lQyLtAIzLBITQuWUBDG5Zf3A7uiMOKq/7KiiA/buPPOsO0y8IKsVaSgXf5KFFR5/vUTgGB1rTwt
1joLniq8pQb7VB6D144jSNQ5xCbwloYDBgrkdBN9MFg1XnJxT8iN1ZO5XmM2CedYAusquCDMzWra
Sey/C2EIBzu4OlP2p8QvrKjzqsUFCqW5imH+WU7+wVKvXU4C/90Z97ZZixI5CbtZhXkaVmf1xNc1
d/aQPdT9RBNOcOB9nnAbhTJD4MtDGDYEO4bGMRKt+d8ulaRlCN8zg/jnQsSgf7HYFTjRp60md15i
b13bQigjenJYUoUTRUW+VT2TGbXJnafvV6TmYNMibLrBMXJ3sXoZUCji+ACDYtKi9zl0EfLby4oo
fvdp2I8UL01zH+a6zWmZhU1moSOOHZ01GXMCqHO8kQcW8u4qR7j61DWmnyEzGFXNeNojXQws1E40
nBWJkQAkeQGlYUYUupXIrBPxMCuE7gdVB9lWIAPAnjgIl3ycwOwj3k9Z709AClWoqo3+/MKsNQa9
Sf7ezhUSlFYPeB8+aonPTA6/baXLuBnq4xHQf0orPg6rkqbiEIhoRKJZDhC5973VwICUfb1f0wvV
lnk/w+wKGTcQFlabDOa/dBkeTfJF8k35NDj0jww4XzAtEW6OI7QPog42suTZ1rRD1zwDXE0BzmSd
NhR4zVmhzkbYGAj/8RVaC/DGuVlhcqKCRt2aW5XY9y488lkljct93W8ArVJ4k99cyrJ2Qn/Kv5PG
uIsVwi/qOfxEb20NSMnXE0R9wirWJ0LS5A5lsbHXAiRDP/WOiZm/4/s3GtzvI427/VOKrTnsOeLI
g6az7ZJeSOtgtU9x5zGfEB6knLoZ3s3IQCJtZwuifFDeQmy/aCBWig0puiwlrdBsF/bJjTTixEtr
cImXseUEXBSVf7cT/d5jtKxY+q5Sy5jJnv4kd5M7YhIAQFS+q9eluBj5+ocY0IfDrRGS9yLe6T7l
JjKgu+eTqK6w51sZEOrR/MNXpjcW5prN8uh/YUsTTF9gB241wnY7eRpyfK32RYZy9LITAFRG83UK
id/YL9TMl/J1pB/GhDRViGXooFRXNxh8o9FPpFEwjovEVHETu5I2BlPOmGqoH19qHwT76sNEiwef
rykZPrgF7MqLNdW467nZ43pAAWcip5yQC9kbu6vy51ZjkaOPKeqAeesPzLuDIX9d1WBg9WFpcgyo
sWABd4rdbfHDfGbgfP+MF16qfy8N22b1lNuIsKo2x61QEh1moAkkT44zOXC3EN0tsY7KlTFQyjwj
IMP4vet1TtKFXHLTlE4rM/BWPG6dXz1MJOuRBW9G4SDA7Pe4f7QaO2TLEttW+DMzIzCRS8VSAYuW
DX8wefl78ANWeM27l1YAgLSL19pHa6MnPqa5ceXB3KUcgebtvva0JocnmCaT+Pi0hEBL5l3v7c+9
7hfrW0QGSq6YElgP1KzV97+0bxne1cVgfDs0zRoqdcbUBbA4s9a0WrPVd3qa07zwlj1cQUqLGVkm
DmRGmtBJtA==
`protect end_protected

