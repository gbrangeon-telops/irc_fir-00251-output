

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
dpj1rsbRiC2XtvMMkZeaWceey8TRzfvuZghjsYUFfvEbx0wxaUtNO2KtH3hQvHr5R05ZRpFvbxnS
y9eflHJ+fw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
RxF4+BsurVIN9R6VPOZY6IjRgF7yOLOJFH+DEaCvilnRUUfGXWquiAJNpzEAXSnsWuptbwUxy5M0
I2FA4+Rh4icthIWWJqsNOFS1K2ZEpNoHe2hVsMzmtRpnsPL9VGvgfvA4do7AYV7YhTUgoQfClGAQ
vFYxy/RbXBzM3PrDcTk=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
OvIp9LkjFoctqOSaxZyP7bYL7KElD3vYsFbzOXm+yqBzueGP4aoe0+732BJK3cSRYLmSREwKo0o0
Rv3hIBpxf0Y7nOdTTISL4pJ3qn/Q9Div9rDMzGaVxIOMLNLxqjT1ZbqCGU0LBxVzmDxHhBalP4V2
XUBBBCK3eeYn9YA+pujel3BBQ67ibuZRmgjKTwyT9B3SaGu2w8ce0O/YfSF/l+ncmV9cvUhjGdBV
Dsus1J4qhNTtraXR3S8daDpX289UCjsNh8krOgCnmBNlKeEFeTxbhmhnNPIAjDgfW1fdIgrmAH+S
tzDecIht4fghpU24F+FmCjpRFfArF8+d7uvxlA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
4ZEqShxRoOQpy+XtDUXlHHAe5v38IR2wWpAtAq2KeZ3f4UCuk5LQw2Oc5c9xFXi1a9SsCAzYO6Rg
6iBcvyh5jboOYApBCjz/4VZfMAndhqby+l7lpAzkB6TqAqvqUfdVhSRn9DQMcQZ2fMALj61IBeLk
rnvtNe9XfB9vaA3zmlE=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
CxLbTp2UMBa44c/UwixvnmtRjPsy2Xb+fkOsP/coXETbFAb6XdUuKlopddrCIslByXBY8SiCzN9B
XnnZENqObWvYgo2VDZVlPu9SL8ZNuOrh2v/bJ7ztAhTSojfY2dBi8ojKva7J9JwGsRtKubJGASjY
RHw8CGw4rdc0A5dMEVmmoAymqmzBjExIxX3UWjtVz457DADxQ6UUgPgr7ysxQXkHN2eTr8eKtbK1
R8VALM11jq0MxZUpiiq5xDX4POkxGrs4QQL6Repo1WUK5V648ZRUZDaWyRJbcIm/J5ref1gzTZWX
h3koqZ0X3HGeO0DTx9nnC43UDVfA3fgk+YpVGw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 33472)
`protect data_block
1nhzbJg/7juDVTAk5QsyRQZ1dIYWpTOMmK+elnf2r8i9aRy7Jy/jMyokh4bRUiUH2jLtkrfyCSMC
oyy6KmrYiG6neN13fJrMiZQ46OMcD4OFfrcogoayf07dqMkIsTiKyxf91vKt+7+kzLy/ZjqBa9YR
nYQeMcKvge6PUzDtm49T/aX79fDsz2kz9o8Cpq3yf6H7izrUzaH2ccikrJEQqEuZpBP5A3SARoKs
J5nqo8V9jUfODqPtw1CrKAsal0IcQt1oK8VOV/PRXQK+1vXbkk+cAilSfqOhkwdqel03b5y3Y5VL
XG83zjld0XnOw5cabL+tkVEcuymaO3Cnb0MymyAWDde5r41uCFkCStb7JCIWS6qu639Qt6L+zY/M
/pINzow2xhHagsAzwKG8QRUzO0gPbuLpLlvjqBHX5a6BdRV0nPQoK5iZSSzr1hjEhPKdrb3kEkxW
HucztelNtGCAFMrVMTa4R1K3nVqBiy9LD88WtXPfARwhd4SQocJXiFRDWQIF4ldlozf43a0glaf1
vBPri9odR12SaQcxzZAJYdTlDQGcWzJ63G+WdzK3kYXQHqSvOtm3PfEGzf8PP10pRVdqUznn00Iv
7fTaeaxxPxUW3RkFOFyzYthHZK0Brw2wQmI9GfVUYP8gPr+2t5jTMg92LT4YepEC1aQLsmjqITfZ
GaQ2+6cO6mzxqSslrcYCzn+INHi32VCvYKZh7VAFDcdB/tN5thgivvP/SjPdCFTLZo3yW3G28KXb
+0VQJaLwCHLDF8f1jiDJySBmh2ABuoscEkEOtidqe1L2pKATEZ0mXXdjTTLZC+LWheq+oyRwffpC
QU1B7ekPsAWm106aAULdNTzesuwk4L5/FCmkgjc2df155Q8Kjui1ioO7kTpeGq1zHuRdzZc1/AF3
t0a5tyAU2njeSI4PQnZ5J2V2chPAOoJU7JX5wv7F+3llCCuPQ5ElX0gGjY4PhxoekCFKFBWeg2sq
lBwq5tLVZCa6ohNVXd54HzwHMqLYHORxp1vCK37bKx8jwccATrJUUKD9Ev/qKY7DI1Icqim44/VW
YVi9cZ6bmrMRgG5+luM0b46D+Zd0TQ0VfZOZ3OCtnJj/UIcYhr5lLHaCRq1oz2V5WFCYhtA+SeXG
3vCtfp2kGnlqW7PrdFGXzHcDWIs/1WurdtXO3l9Di8SArW01qU/Uf8eHps1WeESZMymPdt105DgX
vtgvW1RJ8CnvLCIG4yDcOZevpZPd5PjdGmIP6Cocb0dibdjlMr+2NuugZnwBv27Ahs8EBClHwZeY
72rqlOlAfSsN1FZObhIBLoSxNBMqvmtHHQ770ByxdGybPFkGo3cmfFSDQU0yVu1E/iS6j4BXpvQT
4v36Q0AyULTZUldqkaPPiC/+xyN5VkUm+3npIwYw4ZwFfvz+M3TByU/gXxqe7jvpu6593qIgyGyI
4VTv5W+iLpiDvEvfrzHITtY/hyCSG2ILG4H4ZOD3jl8HDNu+9XrxKieTw6K5zn6wlGGfysjVR//9
3pJr8C4QFRmtd1Da5+O2Ex6ieF+DOkRTcEVphWgZPou4/bJJIsvs7SpHWYgaxkI6vUD2mz6w+aHu
/6FxBkRE9ZWCj9067a+Y5zPMm2r53tAPM7MToRAuDtKTgZ6Q9sClHm6uOE+4rBmlAOCCVispsTiB
1yGVMFhQbQQ9rjxB8+BQ8Gtgii/CoTaQT7ErA/lZWJ6nM7EdIFWfRmvHA/yAfOxpoJevr4ETRYyJ
E9a1+oT/v9slVMKxgQalbQ1s2Wl/1PHCxK0WjmF0RhzdQXX7s9qZ0E0jzGeokgKKhfPYO5wZLrZJ
SZoEeS22cx4jAiATBOonk4gDxZq2az/8AnfzlUUSiaeHyyF9gUKRDhSA++tbsiRXOl0IgHzQOLGp
sWkG5d8nwz6vnerWBn42ranvZkk0Uia5fmIag+EP22Qdqi9wGFxdMT5Kxnkp0SehT71Z0c0dnSMD
y+Iz145uRSENtdTuO3cZwEQXmclKwd1B43oxFPbzk3zfB4khiCrSvX7b/4bKVHk02ym6vYT5C/fk
CD5g/CZPE+a8glf9UUfdfJVijJWZ4TC4swCHw72d4carU0AAzXtCnN6jxevsuxWfSesVpohGyey8
quesUV8t+yLYDqwhaeZCW0ZN9v10lOQGbYsv3xncx2P/ZCzMFmC1l+XBU2AZ+GhxUCwb9G+jFoOb
CG2tINxctH++YIox0JCJqsaaQ7RIpBBMbZDtvmAX6oRqmrK8yNDJ+On8ydh/MLPeOEW/CtEW7Jrb
LnwqSv8rALCfP23p2WC8GiZO+z0Yo9ZloTbJObpwYpAM8JQwH7ijoxAvY8DbA/UVuFCXZlDAi9LH
GeEgjzT0lqC2x7d+X7Do3CRea+zzGZ4rj+XxFORaymzPiVZ/GWdfip4W1FH8fUzx/Ibx/MjInOrS
xnl9yboesczi3l3F8ggEMqn250IDI0/8TqTzk+6FmFPkP8FOgm2+tbs3ASbYuQCVpW3/KrqYSL2W
42jmgpnbSEtHYupsL9kD66MAmENYsWKDxqtbdnviBPls0FiEzJb6jAcwkfx/xpvExYo+FfOinV2E
ZswBo8pTUgApe+cxaekQIRbWeDrkotbz2ETnYUXkGL3e8aVOKexMiqF4yI+fmdLEsVc/Nn+m/sF0
B2CHII9d+fOXkrDzWAIv9S6fexqKyp9VEnfaaq9QQ3pi5zqeOJfWK3bcF4Wg5Or+4+3r90NZLMUb
9nsgDimkYJV02qTnq5M2q+pXhsmKgFvnLdq0Qk5/fCj6HeDKfCu9h2rQmQ4kUJsJBOxgG/uFaRQq
rvj1zg9Qv/EEBcFdPUj2iGXsAUrjILiFuoSFh6RINB0pxvb8j8PNT6ublf1wdHvn4DbekTgsDQ9R
whDQ3Ov9WEvrna4GX1sjOG9UftrPJPepbcVAI3NhNsHN3uPVDQMM+fioADWB/Gy1+81o/mzUFJR5
7XSLdJYgp4iSHwIfVBfGzPSGWSsvUP431yv8yvyxY3QHqdrBdW856VBBw1Z9H/MJyiT7nJPbEssC
yxO2m85qHFEtraQ1u75gkDpEYQhdmkpiv7YGQM+7JwS0ohhiV6Oeux4dB3zPlYKRg1eaDio3Kvkf
2oNBlaN9cdLDgySzkGQR59cyX8pFMR1n6h9yc7Dpa8XDdq+TQ4BBGha23kG+tnkUzZK1CwoZWCua
STAEcC+oXbzEvrKQ9b8YjKgAuA8x3ASIphmKFJ5Wf4PDjdnMGYCMjm4cfLm6I7fHbuR3yxhKxErz
sGbeuqYBj/Z2cjY6btvC+3GY7xjoXj8BkpNsV8/iB94IlVwTNZd/KJ6VE57e+SQ2Q8vXPlwZmSi1
f48w7WNynB3SwVBbdYnT09lKtyBVsuA2JmrV01AD/QF7HQLqh2oo6U/KgXUJyuJvKMkYQORPCQhI
aBJHMn++QsaM9BnJ7SR0n4jsMxHNuZx5HbdLF5PjXmAihbtxAsPTeFUby35dHMgaL2QamaNpIUiG
xN2HExGQMQar2rkBcVbNOQL9z7VO1Vg6hm0N9UrvXu1zbk6pFgiTuwIo3VbSPjenB1nSnoGyi+nK
X9XHtqghOpKaliUkLgqx6oeluuq+A7nE6O7rRusFft5PGW2UteDMcsCTSZYnTQySebWgicSwKyET
n/pgo6E+yvPps5s3zibRoYC8kjTYIKxqubsLCjnZuZFCsgZw4WQo4KD2tTGsrSeMgTtyZTtE/7ya
uI0AFt7Bk/+yRBCwknx8x777+byulaHYV3NpUhvPdfLiiw6Blc8uZMAbXne6H2D+U8ydjies5bfi
t6bI7RN5aa0BOcwETayyJpwGgjC9XOTQvACNppzawdtTJ1V4j8QtGLF3uTE+RAl9GC9xXIN0dU31
xIzQBd3WjixU4stXQ8QrlpV5/q/OuVdkLo2KY7Te7pUWsXNOx2Ke19RD3fSBDdB6vPXmit3o2lhG
Hel1PFqCkXqt466IJz6+Y8faNjJbZ9GDvpDO+SrHD3mxIsx7a8U7kbEqhDQ8FMpLMs7VreCZ+bk/
xEAJZ6fq6S9z2gozoFRB7amCI3fsyud8vN3tZx2ZsiClagflrm/w6V9SPymDJRv8V7cV2KCYfnTk
uS2K2cUy79h37Vvo22fTBc+sd2BxZzHFWsv17XSqtoeg27T5ClZRcyQTc5zYFg7FDf7JOOjSFK7j
2yph72zvvgReeBA186ubvr2a0w+tdtn7yHXuaoJGSOowKIRVao+Rq8do8A6hq539Rnq+UR0VjSG4
tIYnnBFOenq/1bVddSZWMYFnl+uXsDuMXLnMJsgK/GZCPRiio78AoyQCu5gldSAFjYxGnxSRSx29
7QVy3KJPMwWdY/DmiYGfJVfTC/45ZDWpLGXOwVhEf8P8gXperhwWGxzmZhMk0azZy/KqPQNvJjDs
h7UvlFhVS1KO4jbswKaB++fZohORmqGihktQOiiwzt63kScV8v0gnxV9FhmycmfdwfEoAbFYhQ1m
H76TMJB4zrgNx/5gjY04Nmj48XXbUKxr0eu1qFouPdYjWA0SnUxNdF4mkjEoqHvgf7un0r3B5KPW
cEAe4XaVb4WgIPCyQ9KkZ6n4k1CsLuuy+tr5uyCHgZ7AEf7IAkPGCQ71xAli/20IaTOj+r0AmNDs
pWFIwzE3Zko0ulQ/2UNJSLR2L8djD0nsDlFrdnzYIddCCsdG8DSw9B/ZhAZolA4/376sa2KeeVE/
KRMsBordwgGWD5D9AKGvUipn6DdDSNNUsBGs2R5gLzKLFV41D43HQ9q5auQBceGcTUfWqIC7Qx0h
86Tpymtz9nZj6da2uZAkBl6PlUjSsu2PtgaB16rCsWXbjzXnZUNeKAluuiteoj7hHIW3iLWXa0+f
IBw5b7C8wP0uu0ZtXv5cASlMsidHrkCzyweKLNPt69MLLKJVouHRNA11d1LDcpsF6zrjFi4QyDrl
0uCHLfii/dPPVMP/XLSufRXxmHScOlvxi5T7f96eVDIrCjHP3rx5HDFu4KZOaiCGfE59BgBJpZk0
7vzvtkOYO07bPV3KuX0EmghYXEnPpp+lmIcZO4jlI567OYL2O/DRq3iPilCFiHihA5k6g1mMdeTp
cn4IQc1nYcOCcg9eURb4DGyMYYxnnNrYMbt3haXN9vuviudRJWQTC4M0K4ukt/3aY3ZyCkHRi0JR
JuNGcf2vbvFolTKoJ3A4LBv4rTGtYiOitENZm83aPQevUiW2u0PJS2AlBwEeVtZdkQvRMO+D9cY1
T1sA/U9MUP2qE/cPOCOxlYldlg/rYmMUe66jaATpHpYh9Th/ljH3A8Rp3aWhy4XgZAZC/o5rsckZ
0EWddDufmoglCwE0LcKHjshwqMGS0FaotWrIKupyDs+D/I6fk6yBN+OjnEyKD7SRcuNgH5lU/uIg
F6XyxWZ06D3Wc2rBpftfJDtU1pcew/HVmhx/+6jre+pNvavjfX1kTml2XKkOw0EUOlyyMbSSnIBI
IMhnhvyuuklEkGh4MjjCxAor1CuJ8/R8uUJhgTfaq56e8wCar6TrCDeuKHRDCwJfBIqgiKMAFQsn
Gja6S46u/zLuEckHaI1K1G0Jj6fHwRE9rbvbgjz7ozCW8onPRBeYx+9Jc2PsTpcMahzA9tTpdXJl
Ea3qv4nnzDdOg8fEONKc0XLC3Xd63o7PSW+O8+4I0JJfX0UPRjZOk9UEokJbsEy1Q5eeNzsfCopY
NFNz+iREypPd5VEcX+fogV5WZH/rFiLdB981Ctt2aaPL7OkMl9Z7VRpmHoJobiKmOreEwcKr7C2X
OLM7hpLQNkxZjJSCkve4YyXcxKpecsx+EyY8Lb89I0mwIjlr0kcr3F230/j1FO59iFLLoDWWwN3J
NxUQzz7JoiYNM5rrcX1zZWXeJtHQ5Q67YfswjmST+iq31wNbwq7A/9/YmoiKBQy2ABw2g5dlYryq
lag38Qmn+hZKiCeKJUgDE8quvLJavXhZqJr5e/Fl9OLI9rAqb/NH/RGnZrmUSzEzPa5/pqL6BE1y
BlBz8inL7b6jn0CF8UJ3aoSnY+BtaHJtp7opVf5+P+24NN/GM/aE5k3sEoIzdFCy2JJd8nSiwxC6
MmXadVacqBxpm2VAlwQLhtM0aeiVJp8I4O5Mxu/GWOan7TcJjvBkYpTodv+n2qCgEOFx6ZU+7N/s
MoEV23vMyLmz27Adgh0R9oFQBv0IaN2OFLfuIB4oY1DhIrD6+o5fESUKQknGtRsgr+0DQtarY8Il
33gZgqnekTFq4ZoZ+QZ2akIyCTOe9/e4RDi8FjNWMwnM7ggqHJYA8hHJqgfb6Gq8Njs2D+3BKilC
TNrb6hRV/xdJtBKJyn8vCOUBVx4VGkYgHXjOc9a/0DIpn/JhcHIxbBS1rtxbwoLbpDNPnR0oPGA6
ofU1JWa+r07Fgm3nimw8YlOD9eT5sO1+q5ySlOd+3eDsyXevLAaLIp3tx6JzDs9mD72kOyYU/KrS
qysj7RE5SWNFzYvyGGRNofvJPRKN0/xGzjILaU2XqTdkJ7Q6u65bTZm8Gxbz2h0ff2IdRx/LqKJt
JxBfI7NB/wVTpSxuHmH73ZfbIlzWf+MRYjKrITgYd9N+yQwbeGzLmuRO0RkK8mEHbwCQHg6EXjIU
C4BhiOhL9IG8Fq/oiH5DUS+RwFzNfSWGsQHBfz/TKz41GGiH7tyoECyC2P/OcD2Hu3gz6bNoGwE6
eUqm11a4yHS020JOeLbln1j3iqyGYH7hQQWvadW4ZWwJKd7Yohph91/clDcpGAMk6s6O3SJ91DwU
w6vSQQml4fvHphf82n3DNxllxnmAw7ZjLMEKiscYhS4xYa6vlAedw4YkuPzWDRPmVJMEWBtZyNnI
9X5ZDSg2awB6lBFEwU8ATrez9AIUVkPKlV9Jz7UQ5xnHRpjqO87HVZqLjCz3dtyawGy/rcTag5u6
41Ahn42x4TRedcdUvZ4Y6kjIjV/zAXlpYIiglRlOD6cxk7fXBqoJAFtLfBUoBsz7dMWyNDf0N8YX
mEytIozmIDNeab/GhicESM+mK1UIL3kjQowvKaULwsNt0odL2t/9SBpU+kkgOutoZuoSFMSxAz2i
pPJVyOrmf3jxnCxX7Cs9Scw1R81flP4WMqDeaWDJZY0tCgrNqdAaTEYinvdiNQeWD6fN9GKgEIPi
yLOmym+iSvBu8VE3SVtTmWcAE8VqlUazOCMhmD0lv4nJZrvb+6Og+NrZvH2OJ2jDjuGNN30vEsjr
RfKsUj+nF1I2uExwoNnQ/2aRRFEy6GzdTxGIp4D3di7lvI/w5foW8oaX9wE2wlj53zoHOz5JPq0o
mQ0SXHsqHcHjnaWX4QK8dSPdlbRFPETIqTR12EGZdBvUwcvhC/6rJLsmFK6/RK/VVAG8FsViM6Xg
guzsBxwWDiw4LXBCOOmadJJ0+IgkoRGZtKazqG85wD29Ru7bQbvO3+k1bHPO6ai1k8KySwp/MZmc
E7WfRrtH4iTkqpr4XKghYsWvhoQPaoRSA73afl5z5VwsIragZ2hB0DDoQYlTb+KS0RrqU40KSgae
cCIwl6mmgH+F+9QbKfA0gfJYKmm8sHil+b1kaP8/m9IJiDMLlFnheSl0vrPG9sJmOrayFduTTtUj
gSjhp4gsWEzHzreND6PZkjBnLMeG7TQDxoHbVca6CJBQ4C5avit38dvmOayjqLCCBNTFkB+fK2fM
RAg/Klx6qV+eFiVDiw1rh2sR4fzKuLNHuzmdy70MnNpJqr9SeFwzasKK6iDVC6z8GDZvD8Lm8hIz
hc4Su9vbun+HPDN6u2dfyoePW2lksm7k+fj4L6TLorYOFDAzr/hT/GkheUAZ1y2iK3cZunFCD+Ai
qa4MbD6sQ8/Z7grTpmkOIVbQsP/T7p1lrvdmtIoC+BglSnuByRqZW/zzWNJhLuROoh5yew/et5CM
69n8ADqgtXu9u1Cy4R6Qapj/s3msFSg4sXGrdSDriGSM72KYGIxPHInoWjV0Jqc8vttTcjPyKao/
Ku6fEoIu1WSKAoA2WHCDOzO59PrADT7phjaGUPO8uNR2hdlt2hnk+oYhO9PXY+QJ7rR1nZVWt9vb
pQR7NMnH84tE0CA31akUPMpPmC+Rcj4uugW2x9y/to+R4TJW8fKw7mPsc0WFFaPjyRabb69RYO7h
VIxGJx3Ky2doUhZfLbGGlXqn06UL4TEopd43p6Vg2xMuqZlnSOBJGKtuVJZ0HULS4r3mGRV/sQjL
SgSav09WXjlJFRrpjl5jW/sz9F/pgcBvuneiU+jeq6Jzh8+rlBUNs+kW/z8B8W40pxnE8wG7rvUV
2QWdm0ufw5rk+mgQObcUG4QxMMf1j1Z95Pp3+f3evWt6xKQOuy+bf+FU0oMdCL3Loznk1K0tmrXl
dorH4Boja1Dzr9XsxdVTUB0zq1elaZxFMqNgyYy5q86YqLQ4QeVZ/DGBlmUGMP+UEQlWJrShygTp
SlckkRBBGEmFv5D86mSzuFIbnfreod/sljUVvwKluVh+2E9Ij0/Kvy3QuXpCGjzwiVd/e/Jnd3xJ
JXGyDAmEA6o3LN8YbFE1ytboXOrKpUgQ5YtluMor7LROozOOMbhb8zAsD20JJGeLxmUejG40x1zd
2Z+F+eaRogzZdZVnFLkxYh20CrM1yr6Od3tlPbICX1CZfpZlYUkHawnghSbrPJjsKdzPJ2dQkN8r
m63TcnOwNUDzVFg1S674T6327XObU4r48x2Tag/OLcru6UVUqyw2Dy1uufGGGWrvXiZU7J3EWL6H
yED1ViE3w33Krd017vZeZ+nPArR7YxYUN2yVt58ArRi0+ywf/DKdSx5K0xS7/rbO0eGHKu9fURhT
85Ypnr5EKI4NUZ1hP3I+KBtdM8fotfhdWI3R/nKdqV9ysypjN2205wGckj+6YZNCyl9Ztjo9iPq/
bLIWQd2xe4cX3iOib8jNPZW34X8CFBqhsAtMY9jc/SPEqi+gkMqc6kVvxvSZGKYbhAzAv67Ua8xi
xe/EFWgNPGHD+arQQtezKxmT/MyiIyOJU1gyiBiwBHNYBXuGJ1JWZkWlgqWHzwR3V7xHPgt+bx8X
xC5lwd8dsrgs9AIDa7qfdpcCaascOpeYKqM+dW5rtTR7Eykkjdym69aZ+DQHbCLf9f+S4RFsdyqq
m7cxq4XU4j1flH07wn+F8ed9qYe4wpy6se77pWM/Vc11WTKOK2NNujYcWG/ZX2I8W032JY2zXKY5
ieGFmR+17KB9OmSkOUS2YxsuSSoSpsMcKB2IMTvqA52Cm2HFZWwCrocxJ8zsJMO6EC6sDj56j0Bf
uj11plDXTeOgpJIMyR4RkD4PMRHDKIMk0jN6c8u6PK/3pNBBpr6uEeXNJfHy5JTQ4baICTiz6Gj+
99pnmrjNN7/ajOGKOUA/tmAVScrgpiVZ7xQPOtN1mz3ih1AG3TxlVdGZiEv9Yd2Lhea0V16bUcDU
ytUr7vzrElvEknOw37s2dNdp96k1cTsWtsCeBuO/EBCFHsHlvySXSs5sAWxyCPM3LfzWCq9UeXqZ
C9Wd18NTAeAb8RiKxTe9RKRU8YQsj5zSwWcjUC0ODEQf3JXcCytmUm8Ta15Xr+EJjnpmNB57PNlP
PQ3FLMJpD0VZSvOpC7NqZps142vvwjbHdfgcgH0WDqm5e1rRF0QeF5QAJvzAiooC10nlA9JtVFnB
6RG1slyiSHNhvaa+OAVN8Xtw8ZhQ7mV8Bsq4BiZOW6rQ02OLvvgFIeg6o9U+H+KkeLqFS+NkDvC1
J6iunR/PMRCjbDKo+RNqttFZOEI0GC6lt6+N70oEi9yp8Mb7yOcSci2wFSKtiMigwE3qHA0++w15
I57ZVnSKIi3LLXkXaBOYC+iE68QlEHgeVMAPMi50eEVBSY+TT+j6WQqPwT/XAHrOnrr20ZL61e1v
uk7c8+gfTT32lXxKZCzlmMGq2aHODFGWZBlXbHlPNRW9LQpnwXsWiputxsbw85vtJoryV7HyrlGT
TICqshWvWt7grkffGuNQLPwYY7jlmNU28dk+15ErfoJgcCRfBQF1TnzVg1nAgK/XmCYETDxdZnmY
xLpGbvBZzyyEaCc01abpInS2fcLJqgJfWSNJEqCrL3zSYWxyEltB6XQeBiLumDj82O2lmj8qg0Tp
KJCJYEn2fnIdWkRK4ZRDzakU/qnc9yr5Gr7vM6CebAzo6xR62tr9nKY4L/HxYXZCVAZ3qyFtonhO
I/h/AbHJn3DJtkgoR630npVKwy+0efnhiZ9c5eeg+69A6vV42kCq5blKshcduDTi6o/eGfKDNNID
HcNkVq1O4GBAV//ZRrS0XYHeqyoOQhxdghDmWc2TBjfG/d1QhY+KyMjiyFOqFCNVuXOOZ6F9vXVc
ucEHuXALVlfyrDt8Eo5nZVxMKprb+AcqzCYewGeHJMPRWiApdCwMoCY8m0qTfoGIcx/0Pn/gfQbR
/CutMY73od4xqoBgoreeX/i2DFwtZqO0/0t9Ms76pOlYKnVcGu4oUOjP/g5o+AtDlS6Bq8BCTH9M
MkPnldMoPs/iuPXQey8apfSc7I4mfbbW53cR0kLPhX/JDmlDCCBAAy9/P2yW0ZVQhZrIs3MCOh3c
bFlDltbOKbpNQPO1QZj7cANmXQPsMqif9BRGdyK42bhcVGNWanpzJKFvfV4JvkqWzVMSnQkV3uU/
b5LNEWYTJqeFPNuSVbmh0aUg/Wn5psfWnv2wY2kAsyadbL3kmXeeqlNpCTmE9S2XPrN8Vj/LcGmU
vgogPhSvDQsYjemnM2+Hu0lFNJXlignALwuT25OR9AWp2FCPqT6owQ5ua/hrTNeQbVWJuNIXBBaF
ZhG/Auhh32ddvJ9ejO+HIXwMlgTVZ964MinoC8pP5jemQdnuBlCYVzmZaxFRoTSD4b7uj0tcrf8S
9hGqS83wOimdjqJPJsguo6/z364AeUOqi0W42a8SIpeMqTeTDkajPgOcNEP9U0kf+s76MVt1acM8
txGbw4bq9HNWA496MewJy4eEIEjPKs1L3UwPTicfWo3DBEbephqf64sBtfH6g0A83IE4pDG2SOjq
XlXpP1ET28g0uE1gm1WeaPlOEwxH3DFM1lPy2JGw5EbpLR/RD77i8mrBXW4NsVOyFeiG/7A53cib
zumP9W4IhBCSIGNjgLlC0cW/e1ZIEQr133TCxHW/qXeiUSDJBqISWTG2gpABC5RsYbI76zE+lYhF
m9hXZQlXaDO6BayQkREv3ucL0PvF7yVJqxHqHd5NYYyYN91fC6/NHGro3y4LId/cVtWH1IExU/gA
moUYsk2kVvOHQJZh+CubAyexy0s6N7UMUavnR7AvDqvjpAvDXyESps+wEut3sPOPx/fk0vKkXHHV
iycjLQ7pBRdbJ8KlMqAXvMyVSjZXqcVtQqgbHCQN5JDax2N6Mb6mPOqmKg+0aMBmlasPgKN9RetF
+pVD4+fsDUL8lZvziL+nUVfugKn99PVUu1nr3Dc6e5ZMpVLnsUr0bYK47h0caxQXDC2Hvq6c5SgA
VExJgSh+aQoHZCoqICeqCpTrey7WY2+8jhMIvAxAy/apAVN08pJ1Ovnf4fEe+YoBMovkWzn33F0e
5VfbVBPcgRpk5OlOaAqpk3UikwXmENqBe/M9RXOLG9FdW1aZp9JFAqH30THwObrmZvAIi6dIYwV5
SsDD0ZQJWgf/j+f1WLYKMeBbmQGxsl9CNqHAXMlF4bnXuVCDSMJZcYnczRmn5tsrgNWf6qLnvorv
icW9DFs6T0iEvnfud5lwSsKtf4mkS2uK8u/CHVWD/BILB7By4/S2LjqgxUOScnMXJADKmfpXidhG
7bp2kz1hP9Ie/ym4UX9sB3wXSnFUAs/4kYHiitZ76/LuJAzDamoJe40/IrBNiU0lnGHrKS3EsS0u
nmyuD532DRkl42TsUxtllUbuqoKyh9Xz0E4ZV0Qx4D1wv77uUmItTB5J5beYA+dFiU58xnDmurfv
k2GYWZvd6/Lr0oo2I2VlF0MBPm8wjkujUcNDCT2zZEIcPCO2x7obSE/Exj1r7LJ41wC0lF8nW0gP
XstNL9teC6fyLOb3DqCqHKkkCBemfCSyLgvziF4IuOqpcmiX/mKZEFNW4iKJfkoSjeZESFbPVUhT
1hkFqKpSE/MQQNSFNpM65dNZVLZlLVeTUN9ZnHaynQBS7qo4E+FS1o2Uv6V6xlv2PRM2XzuAi9pg
lgIdCROAG9Hxq1s6V5bQb5l5R/xQ+nuNHMih1azo9CcHfz2nLl4BwAXbjZB9S6uUNAiaRvW7evFM
YqbveS6fLThXUbzqq0yhyWMaVjfMkg80CtGZW3ncuAiyt5NMVdR4WjcQ2sXCURgVExmqNU12sXzp
0CJzSF+LbF3TgfUyPR/qvTpotlKDv6Fw5VDvpIyNIJiN/jjWIFYPi1o8B44S7TiOMJ3ROtdmG1JH
20RSrvRkhvDQLz8zJe1W0jXcT+M9MLiR7QHIt+zaMQezrVZmgRK8jVW5Lglr/sBkDaQ6X12xLOXs
OeLRPK1XIdWdtosqbOYH6vLXYWREKySIMYL/Aiwxdmz8WZ6TlZaVY12e/v13MKDBunxoUdMOyoS+
Rm3vcq3SEqgYamhYRpG/xOmTtm4Rqfej4UsVoFQ7WFDaBVH0lizknY3+/p6JH+axnSG2d//Fq4CO
OlgdGqW+q0aAy1RTEP3Opjaok2tfeQ8qoirboxxR3bvVsTF1/vtwY5lmuYkWbLSdSUvrxjDUN6Nd
6WvkUsEgk5ehpigd+qLtQnwpcd3XkrhiITM7uC9NBkVU0gevbXY1syVWCDUZQK+uDS98xMrzOEjh
UEmS3SohmMs7LWcJdQQJARIzsojH9t2ywT4xAMnwCUuadmD+lJJY8inW0qNKCWR1xTrtOsmJuSXI
gLKPuEJd+3giey/YSVwiepJIHGSZUM0SDTCH6OqrW2GemtwZ2RnY39b62PwnjsuBOzdqf36QMej1
M+bfZotaO3rlJu7dyF1sr4OeItrCoZgYMztfEjywVcsayciyoHLWMl4gShaz1hKx/LoEyD0fQEl3
rAhAFX3+d4zW+Pa0HyD/Xr9qz5K1GXQAWtEQeuBmNz88dd5E56XDqW1SbdiRg6jNq6tlIycigLLH
JqVSPXH1KcIzVnqalodnjsPlkeLtuJsUQ/bUCTzCOuCmpX19umLoKreBbYL6aC7LOGCsehTv7hZ/
Pq3/rdg/BCDDHIZoTdj4jTqG3Gz3lGDO72GS8NNeHzktbUcU9Oeef0o4lQVHrUmJ18IEg11svNyY
vPJmDdYkKl0Cp7s+tIi+9YeNudkH8Fj5BtHcb/TfEfx5XspNLsSQkhSZTyRCtxu0O9Lw1dH4rqsR
ilmzxkG7Q3WhmffcJ+ty3bYmYRq00StLA3eBGXof6hvoSYOkSqyjyyRwzZxAkprEGLiV7aoS2I+e
FLttmYdHW/4L5LHH/fMQDsHsrxYsLFoCryZRc1aScu3GDS/pfzYmdnRRzULcO1svIo9hNzjwMhbF
sYoCRoqaEJz6ky1XURKtChpllFKpZbo87WAWRypD7sogAD5O59e2TDWlWIVKrAKukkVQcOJx5N0O
E1AuSYfJzSSGF9GtW2mwRxOHhy3lUMVk1jUsoJ5DaephEtUU5delKVC+usB8iJh3gLyghw3z+T0a
lFRrgmp/mBiaLrWtxj3D7e++rIQ59sstp7Mv7DsrxELvyA9IjU3Zk0yKVgdRDdDmNyA33epM4Lx3
zg1sXNMEoOTmR30b/AaVGW18miVTHd0BfwINKrq6gshw/Gr9/dWJzkY2IuI39bkQ6abL1ov0dySN
Smn0SGIk2C5oRr/Ega9RP1TNWHkIsushnl2rvfI1zOc7OEHvdA3YWBx2VLP/LOMKtMLJPUrtUbRV
sHDDIK8THJi8DNnJgiT8R8F/eg2B77vTedtle+jiT2Y95Sx37fXcGF7eIeGbUyKVwqrI+dJFaujj
DLKe7osWIOUHj5IketLW/3HuJDv2DfzaxahrEI2smUVrvCVOXWnq/GiaDP07gIBeN0aSn6bPAymb
ObDkNdDjzwdd1ZubU6Fym6tNaibouCnRGHl8cayzWM3S1eDnBZnLZjd/gxyNfJ59Apt3eAPjZaUL
f8FK2+yCKeIG1RDXaz++lcm0yHKpExJmiXnxeafTnl1HWh4ATC2CYeK3paInkjhXFKd9pcCPZXdo
M7itpOb/yK47NNjVFESKcOCznjnhvfB6tp6zMqnyqW5l8+PrscRyX6toLFKXC4ferZQojeY9R/Aw
+kiaGEvc7L06S8uuqtxKXfSYrOC5jooUYMTtjL+9Mjs+YY3bfy/iW7PCIXY+1mUqcveCDWvZuvm1
Bp2VU+XwHk/HKxyKw1Qn5KIKDamUHg4ZXaveaxcDlVdxGzP6GqQnGakyEBS1k/fpuQRlTUxAYRfj
X5q3pdG7Ym3P5SoMeUvQkvOTJ3T4J9mrSdsfu5MWHJRba15ZbLa6J31FUwDWsrFRXH8iH+CJ1MXa
E5vK6B3Kn1kZiIDb7xaR1Y14+fxKJ0eADBMP4M1nadMAH1g+jmiq/pjCpzqNTR27GKxYfRLMS1LF
nD9fowz/MeGpA6T32T+2dGYQ11M60oxlCBsaqM39E1MW37rn3Q9etDVGc0pkSh7bPJexVk4KDDwT
MN7Sp34yrT4Nfe3p+TqgmY4DmBqdVuNMJcHe9jbkv/nk6tXVUmUrIODmp98E4FwDGMHG4yqm54US
y8h8+5f9IikoPScTAfu9/99KQyAgu4o4PMVT56+zSEhsuukHtWbfqEHo4UMai67nJkzJNmB/JW8b
Mx3T8DPRb0Mah3UaIN93yjgO3pKYdDhTpRGov615YO7sqPqWKLmEaU4K5EUwpwxYB8YmvJohgcnm
3PVKw4ty2YwNCXYMqDZMVnpgZ1kUkRm132RPTYs9HUbZyAo9pIHLREquI4dMq4xE3N8xu2uqjjGZ
UmGb3Z5y5lHvi/a8tgOXdqZGbfK+GR7crIHEiT8FpLbF/2hHZ6OT4yU+egBplZYiCf45+87aMUij
2YJSlyCybQZ8VgEcQrFfmIDyLJoVciZj/5i93c9msnKefMy2r4rm5BU7IjEE/kpzHrbffuLDRTZN
u2r7PdUk2XrgF3T/oMnJTcSvwb2UsHILYwV5TY80svmnEvyvj+NfgfP6pBZfjWAtpYRomvUJo8yv
bVr5+D6/UBh1UDAFlYKE4LKpGjWztvngUwelthvO70mSg9kgEcK+O1P9PVuC+GIASilJMgmd3z6R
YqI3B2g7p4wZ/5IemDIzd4xA6F2GXsdt3kDFQCk85qhTnBCCii25tcBMSq/BSpXYPKkbLI4e9+J6
lysRigeX3n3/CtV5gQY7o+Xo7wirx7zOVpgcl+vsEhhiRJl56qGoGwPd0rryeDXesUn7h92FbmTS
b7OePmY6aQArqFRCk4S9NBHqrsn+6fuO87tFvgir/X0tELsbHUCMDUnVDHGzgvwp81IO5NBzXot/
xJ7MCRhA8tCrOs8ZWaYQn6W+tsVktjuxDJiw1F4vMbaU8nvx5OebCeOC6od89N6SK27k5A9g1X43
0p8UbLf/oiuCvIvNrf4DLNHuZqMzxpudFnEYjWZJLTiCFaoC9xrgnvAAgAsJ64afN/AYnrKTSnWA
xWNq8mxV4B3ysarHAqXruCw0NWtL+9Rhzuanie87IeW3jwXHl2FgUj496N0vIIw/UNTIzaw/vYbm
q9QR3lhxf903g3tHcBDZDOAqIYVH17RZ4HDzAWGU0q2h7VKJx6N4zzm9m3YYome34DUiqdVqHChD
o6UF3/Z3TRytXayNEkMcZQ/TJcE+tufh3XF5w0i0EZkzyfbhT6wWwUvJwV4feP1I5dHXNOJq/cGM
nyUTw6cpfQSYv5IUpoUoLcJRPHGQq/M+n49iNYa+13hD8IfL7BVSEyk9hpTt2zm7qFLTClYA/Est
0ejKgUyJRUjMaX/RcR0pXV0tueuD9VWwygN9LZ3x4Yo8FIBijH0Dhs6bgSklVmDagzP1/aBcIhjP
XeDR2naR6WwQlKBCzE44pzi4BkOpr8N7MCU13tNHiWVpsF7rimpIyOLGw7XnZOHfFsIe6q4SoV5g
hg0ENA4uQuOFilr7csBGk1cKDDbNvaZs3g81ruinCeT9qJZyQRSnFmiJ8cG2zlSPLAYI++fR/fR9
V8hlXmuO9h5hE/RB0kKgJIy1hZwMsAR7CTFTfpDHeALHeb4u6HBTBo602BpxfzJIIaVXzzefCRNP
KOOCNQf/Mkere2GjKAhkpkji0G3kB9nGZorxYeJcolgWeePvAmmWcnHt2LJpEvIhBogAjw7AInBM
xVb1nBmoxcBznRSIn1z56WIbEB80Ogapw9JY3MSbNdpY6fR7AmAZ08lwuQFEz0T4cJM3TAKxP6Sp
9bYXI2sWNroJgSke3wMaSB2/rOMruKZ2f47kTX9OFgBR51TSK5OjTOzH9mExB03D3s4wj+wwlrqh
ZfWi40h+3LlwhbbiUJlT050IScils8cZnYIeuysdK6FL5JqBs5FnZ1iE8Lu7GS16TbrTAFaAHC9+
hJtlqmH3sBluXP21cgg7VdCjvbENq1+Qoto+0gZiDi00it/5vvimI6gZQTkfUE3DZ2oT5bM2ZxUB
DPj/6Zj3DNRUW78dU16gqVJ7h6hoUEKgpoBaOfo0nZy+HRH8Zht5FQbjxtzp36pcrxftP5rB0Azk
wReoyGNrPIou2aTdxN2AR4ICNbzVobfFzZMrLl9W94uxbtOy1n5nKLbMSR6e6tqFZZtE4QVje5d4
f4fL6X90fpkCLnaEPpaPrgYw9vw6wzlci38yAug+YQho5B+cdYYANE8+hGJ2yMgsxUaoj24IgM9l
Shp59pZeLC9mdz/elaqXgvsYjLeS+zhWAJsVb9XV0mwXY/gk9pS2mMGrz6wcnU6iH2LxBEs0EdeT
9CQeK0OtCP1Z8IihiekqB/jcB2HWlOM/q9g6K3PROkpX8CQwnMKC/6CipWWzLCGDqvEd15AKpxKe
T5Yxtvr+ztRonZqi1nsboQtA0wUJXPhiYATuqKVD4jR/A6zaTnxNun004tmb+Vf3qG9JXmL3SFTa
bIGgBAgGztfHJ30w0S0rDVecCFI2suxkKeIQ6QCz6ZmhNbYM31rREI33xWuCpnFdy+OCYqfVHhvk
8SBdHGwT6Sy99eZlGEeqEY/QICt8LeD6et5dBIOFugL2oy+w0D1Rn3+X9Gk9wY/WFlK3jvZRwr/r
jq08xLxr1p7rY1nzeu6z5/IPBht7HqTCMwDh8oPNAiaaxv1kKNlZV0bazbcWQgeKbQdvYVIOQ4mF
QoLRvJJn25RGC3flM+LFru8pCDQzoMfnYz3iKggO5vLnNC9zxolW2iBbpwUJ9To88d7SLX8tuI1Z
DPAWKyxiDGFL0s7QN3UY9wUYXao47gX94op3ECbc64geG361BUNOGGuC+YhR4XwU+orFWSDnIuL3
vCw/WfqNM1Ppw06mRoojiLB6YISpBHL8SK5OdX56HvBOpLTWwM4/+qBZThrOrdIW7/4DhxTyKMWg
tvOMMwBX95hefp72JOSIVfQzqI+g6IF9emZ0e0zuilv3YwDi6nFoSczW+jQ2P/hgpmTaH3U07exH
DFX31KRs5/kZxYPu8HjJ0JE2n+sbSKrl/GV4XTmVyX6MFrXzK53NV+7JvFguqG4W7n/Dzw4MuNlu
JTLkz7KpsJBGyope7era16NWjyKA0DuLU4jcBr33nL0wwKPoQaYIQc5tz4+GaCFD2xvZji5J5FVF
l/m4Rt+BaY9fSF+h8m7Qlk+5s+QprWLefXTX7Z2/MT6WAp0uZ6AuDxfTaWDeSe16q5dY/iFfy4FZ
208a20hzJuJ2lMfm8Qy9i6Kn3V0J/QBKUmQ1xLTx6ewHbpmBLF6e819mmz9dhECeMDtc4RfYIMzT
OfONm4Owl4ZmFsqp6xMLwm/LMYFSQKJqRtHt03VShd093Zrz8rsqZxh2wuaXaeH80X8I9+jfSpN0
o4tSX3w8B1lW08+qWBeMmUwCjo0ckZy3TCAmNtAvEHks2cgYtsyCgJ2+S9ywtNkq5Ue93Q3e6rdj
qQB635rq2pODVil8glxIvuqzS9j66HiAR5Zxh2ZSfdQIXdtWxwo35EJdmQC9kjqmoD8tvIZ3zGkK
phk6Vrjc99qAKez+Jx5Mukor/s5DEsDSoL2qInYe3rXmw14XmceeqjwEw+J18iMviUJuAj9tiM/5
Fx3jxlc+mEH7AZMDfHIlHs80cDqiE3ARmc0TIyFedsfDJZoisM+PU/ZoNgw+m07KCfDwJWkDmzxP
Cb34WrbtbLBymnT49af7b59HRJ/UreewfbHGdFkmbWD07/Vtf2NXRYIhKX723fpUG/f/aY4s9jH1
SN1mUi9/DvjuFM1u1QjywP/k+RFSTmKeUXpB6EIwpfvsB8jePqULUVgRH5dTwvwoyH/GFCiiMF6x
mcs8mPYp6zOJlKb+YXiJ9o7BvmikMdHPdwQuwVTH0XWu8fvaDwE+24dEJAsKc3iYMNZYZmD5QVK4
zMw3wXzREhZ9cqPz8FE2+DnHuISQoqk4WBeBu34F5s7+5KORS7PU4y+VFh5HlYR3O6zwtoJwrE4e
Kc66wWeCR6eV0x85EL1pIjMusSxdaow6aev3UutfRZcA12N2iJAXT3hCB2rTSlKrZsRMd38jWYWs
/h+loQdAwK9vrw3gkXsIxiMWgkdBihXfoHeh9dqixR2qnX5HlNr/1jXwZyBc6wbm7WfiwYHznfx3
GTzwjI2tTkJgQoM5IYrErit/7g+njX5+Fnh/CLvNtkHbFklHPJc14/pLpKkMoaomtKjrAftbkhlz
0gmLZm9NOwyIWk/7QEru++OyxpgSSy9KdQkOMXWWhizu/qtq2xoXVOVLcNeKum7vEYBp4moi/upb
3Q2g/4S/Fb30W5cfgXSmbTADELnVKh0zLxgLCig7PokclrtdxMAe0HkdG862kc+6C4Egymj0o1mJ
DKMoQYqgg2f42/mXvzz5LIR8G/oPrqwJ728Gti/yF4dc9EMSmNddVvQBMzp4UbIJY4NG4JeJp7ad
wLmRExBDI0lEnNrhciOcDpidX+nyLmGbcb3UwG3YZJndlBZqrQf3NXGFwlJsnzyPNFjj/eFZgc6H
d1VcoOWKMx99cgGQ0TMf056GIyjz2N0GZdhAWIqwVPo5/aQZVzNoH1K53IHNarMUz8w0Nk8xTwBY
BNcKGlOu9fkBTfdciErfYQ5Y/DbrwR7sVdtnJz/tUlpSKpudH3Fj/5f8qiJowNIJXWncarhCZk3V
O7ZylMDzmD+bf7zWFZb5+egCqrG62AkSJMtk5tDDOSqQWnVioyd+Epdm+H0Q7ahD75Nzl9EFy5a9
19hPFIy8IiLI/Mg4xahuScBro1iN9B5uHAf1W7JE4oJK7tMjwiuV7FxVzK35+733MNL2gxDu/noA
HeWYkFiF7ZhdoSaTtXUAbSxVKSbbrF2MY1tjCKqQEBZyu8e8vWqlj9ecm5tR0iznOgSgNcrSqAgG
grLoLBLxRcnjJOWEmjLTsV3nfGkTGNEUBFo6SScSJPPBf6zLvBLKaxhyVsatlCFsv6vX/DNoYl4X
14+d49BrxsOTELqM6jbST9hv59XpbsDsbzqmNSVbNsQpSf4/1KwsLLHJ3OC/jFVVEl1b6A7o5a9O
X+TfD+4KJ1WkSmEdeJdSF1R05oVACJ/Po3BBx+eyTd/djIcEWNGkz9svurKn5KJH7f0UyXGNJtCv
/kdvMhPVVUV9apLlo8dsPuhyQNwrIBPteSn4bGpbx1hih4EeiN/rTJb5+michkgw5+xPFe756XJQ
qVw+UfIIsnDBgXIG+r/KPwbGceAxrcAtshn/UadCTnU2jycpJDzI/NyOWzY4XnuQyAyFWoalat8g
VxZ66xyRxp+mvS6QnQUnxGVfIsY/C1wZkV3cMFsE51o7DrzCT7gODXfKIKxeLrVc3fuq/17tTMCA
PcpXXg//+/UUonS5tK0iU26GeZPRPCkOENQrZ1B7xvcunlXcJofO9udAl7CTVjSBtLeZaPljDNHK
0b5vYI6TtiNc7+z/xSzGhQjZd3c/SuPxBWgB+uPeZUPElAE2LmXXmb/JSbQrK+Z5rR5AZxVf4DrL
WS1mxx10ADP8Yn4h7LuwauZ9txKqc0TUGpngz+mKfIoF0bxWeUhVOlGWPYONahx+NKYxdx4JJUT6
9P0HPt3gdUx0oXcPNSH4UT0qbpIEDbi0K+1IjggoQPSRYJTlXjt8/XXjmkfzdGqYn9QLgQSxlOGI
gW+A7UnAiTGCprPoSwiwMEwMOnPpl8VaHAcPY+R8+UDpEONaGc5S9wu5gDcurcfQmAvXQ23EmlyF
zQE6bLYb+9qAdsvDzqtojsh4aLa9WBBtdTrOV3EB2BpWiqGhm3HKB68arMWdB1WZ79p8AD9NvRvw
LMdxF/etIwIs/fHPN8/8OyZQFI+HWSKG16PTXkFAKAORdV1W7IDG0FchwEqpUIDT4Ilxaer1cREl
3i8GxuoEDIiWrGKiJSkxC3fYXXM9dRatRdrBGlAZJI6YUMQXIluI+Uf3lLTzNSuMr6LsJyp8Vk9y
gBLvTa8tyexf0mFhc6aD9B6V6qbnroZ6XAJJW7AgAKIzLS+RoyznTSpZCEKs5bS2p2BZaXMZvAMP
SNKbtzA3SSnPrhJzbP8e3j2dHtwreXz6kJR0IS6TA2h1xzfD6B+fjVi4jo0l7/61Y7m43Q5eUFfU
H9O95xd9CjAW4W5XP3a7G86Hi5mJkLZBh+q4sUdMHWpLJyirSG6cUAQzgy4Zuz0bmlb74rO4I7a2
+CAn2XqhbTNFoSP8CT7gqhNLSyJOh+KyUXwPx3rNQMJAwLvvxDTa9CfgypoC5GDaiGmjtrterzQ1
2cdsUpUNtZtIBSlViCTcCzDSbQj53HaW9gcBlVDv+6Dxiwejw6g/nI0/yF8Kj3DYxV//4HqkHf5z
bQ0ZXH1nMEaW4GnmOjxZ8fAn89uE6nGqF8mtTs9QWbsWjxRhSpByCXoJ3DHmLKoOSdpiIucz2tDh
h931Yz9ssVEcBe8GjG4Gqbr9M8Ubvs+SJUEgTKPegNl7/v+nE4w95j3BhFiH3TsdAv4xjlRwo63b
PiEmWljD/NczULvZO8IObQZZLKXkokW38H8woiysAEoPmPzrMCoOSxLMl2XFoKvZ+5+CNktAF1N4
O1ovhEEYnh8Va6kabkN+YrTqEsMGjNeAFD7sgDRjxPywK2uYJyOxpQxsNptvYzkF0EB405PlXYVY
+mae/bzCw6Z8Xs4TtrnSSZsIsSpDuQUEUhowEI/306GuaUMyW6u1FhRY2hvvHM45N3B7MJOpD3PH
7+C5UVfmAt7Szvn/U0UucTD24DF4+zwgiAKDQ0QVnC+nANoKKn+9BW0I4SlcNpVoWGbAALYvkSVA
wR3F7m//a1YQ90ZgtLty9JnaIGOQEQc9CYxlXy5UcIlzuyUSDC6xWdxVRnA0nuzKr970y/nrqPKD
pC69FqpfhvWl2XhHtYxhNbSuHKA/qTURJZgEcE6EcI4TLW8ndoKfXL31Au7q6MPAKEMm79ilKcq9
mC8sGIHS6Wp9oote1gD3uVo/w0y80nUMLcplnfQ1Rev+KBng5Qh43DRSXolBPH+9qWyb6gv7PcLP
tHNMmm79D6UFmVvsK9+Qe17XJRPp60ywyMEbygtFnsMzTnqp1NhiPdXTqdV2wWNO6zK+5UH+GYhG
sjOMVGZmBky7flCyoiBahqbF9z2nLWXy9M6h1XuzB9wiSW06w7OKNt17LEvjGUPg+tCwwEccWpze
n8xq+hQNnpT3j7j3cPbVxts9jwBXSse1amZULLbpzQvjXezHmxz1GERkU24SOXhpfbINapPgLu3o
2RZlulK4x0ITZMzilZ8xzSfhhsiT5YqxCq6YUL67IEYFP00s+5f9/1Ezgoe7U/3iIDsssabKDIcp
PP35cgn2s2cHTxs7SRUdcX4HaMlauhBJuujC8/8MCePl9/5WQ+ZMSt7PnJtQLdWET1ozaOgRDP+C
QyMC79hrJzeOraHojvfrYMKYQUqqj66O5eLigmKa3jPqeDGxd58bxejeSmJluYlAxooiLzrIwRcb
F6OszSxxeZcXjZt5AVlonisV9iM1oV2yfVV4mCoN4tfQen7+i0e89xZbRD2133wfDSWN9N98uwt+
dWC1bYMU2aqZpip1h66HYZ8pRFPY5//zZ9Bmb4ELgkLxjHv+SZJvVh9pdFNpOaIfDTUboeg2P0Ow
pGLQzOEhhIiE7m9iQfV3ftFkglSbJskOjajVjycYHuDBHCUVI6xXPGOEIsoOV6psTAE1UuA0lGSj
DYQnenj3Z79EhfS2FBEPF4Oj5uubh+89zLT9+0rXAlLGM0KttfpGXZpeiUMTxQSF5ed9FaTN8mJ2
/ivL6+pJKM4pivtrkozYdDGR6ogMyEXmnq5YFJv8jg7PqYvW35Ues3iH0mM0pJOZRZX/jiGP39L6
yDpH3uHXdApSoxjSBECC2aDBnVzfc6hs39E2/IcuCdIObzRxNs19pweuxr2Pm+OHDJJJM48yb9eJ
15F4qMIpIFiRX/2h6/tlNNDa8HBPml5XLbWFEv6JpthpzY+M5veyJuDuHyhas78gbqbOiNMgOnIk
POSWYHQ6tKDnPhXl9JPG33ISnYynDDK+tcfOgJ+LX8XA7a6oupID7i8OmkdUsvhuzNI3j4e6nU9h
+QgKCzN+rTmSSLZ/fDjYXBydYoF6EHSkKYuKIUc2uFrRydtOJ4Cw5ZfJENM8GvBGofvkFCwl7lO0
2GwOzqyhbwWIWgE3H1aCAU/UTUDpwy3KM/me1IJG3zOvv27cLFdOx6ZbDejlUUfUy184vxm3K4Uw
QgdGnsWSfih45FGDz+sS9rBttaui1gXohL0FqgM6kS+egZMEVrovVTwnxdkAcDGAtDLHUgDu64WQ
8FegSGKGbqC8DCRswfCVJYAxoe+gBNJ7Xs55eyKLg5DXkWbOllR4sN3jHiMUWlbV5t/k55EPRlUI
rqcM/IysLsmejD5mzeggOl6FRNwlOKqaEH5LCWUc/NtLaJwLxe6q0y3crX0dEHw7mWWTcqhHs5Zn
7Ndf3MES6gXWXk8fy6ydeD9mARDsWV0kSj21S4DDy/9adGJzKQXtGG9vGIPWuPfQT5IDQpJ9rNGS
bXlDQc+G2zuyFhNMZqL4zv9RSDEyn2NorzKYAj/pDptwtpzO39eNiji2Qqt1yZHWafz0PD5zXQG/
Y4REzGYhjAdnObNvWDu2T7GHNBDRa5TTqhNxn9Q2QrO5WMbH4FpvJX+54WIpJMXd0l5sEDD36xoh
/0lYL+c41gs/mZLT2zJuE55pcsFHc5xux3KvEhDla/+z8nBwx/QCB9HOvOxugfqnEfHw1HnVfRUe
vMnGWDdmTPPH/3gTZ+nRFsFiY4mm5N6UWrOJgOZUI778Q2ISRW8VZ2+hUx1o8Rc+146wAMpB/pVy
i07cv7G8gapu0pstDy5SGWJiqic6/0wksxMbRayp+4o45An0iZWkCHesO70pkZwkmEVYUv3arnAc
7i79SE217KqRTY25EnMxghUG90ni9fZEPBJ534mld2JQ0+wGzh3HkZH45HioWXj3oWBF4QuhxKmW
L3uu6E4GjJWeQB+DfU8saES68W/KdWukU/solVDxNTeggkuM5F11OwRdXQtUyVtfS0/UCvxF+b0Z
D//KqOnrwPKNJlnK9LW3j8pmKJZoqa3uv7mPoz5rWieOp2LUsLD0v++PzKW3oZ6GnP2gH0Km9LB0
0yJrc6mGlmeeWConZkZKhGvYfg80gv6bHZq6WUpvvztVjEG6o6O6ycoo4wBw2PI8bjW3qQbZfhbJ
TRNWjDAUR2aoCruuxa8fOUXzPlKE7GHgEeMsXNXfGjzEAWdvoGCrj/1w8oNxzugxyKyHwVvX+5RN
PrN7kvfyk8+AxIkJG1RmsGWDU+6RkEaqmzEUAKJBZT49HMg57ZrgDZ+EI3li9cbGU4yzFDS1R2GQ
cUKysJrwWCgwE6L363W39nOvdZxcMvYjDQvyk939zENNtBzc5J/pgXw75xXUWBuL3VLZSGwExHdh
0A8BoJYMKEsAs/kHXT0xyzgXgynmval6E1WisOAjTSockmxlwWDOZ41cWLQmI8CORP0G/7Ej6RwB
YhEOrlMQB9rPIav0HtacJmk3PmA3YFO+u5Tt51iL6W4Gp4Y930EBfr7PvmEp6x+5+OYurCIXNaI/
zOmdK9JZ79waoNJwd+WXvNRw48ySUrC8KD7V4Wxmc0xaQQQLyjt/+gK3LtyWqfx7n+KPtmSMAd+v
YuT16Scfj63DP2awseefrvLSMqKBclCUhg1fOEdnu4XIosvBdmRjgV63X8Bz22nb88QpIUNIDiGz
NkCxQ5rav7Cg/hzTb2ZABUy7ifdhjCAppwPJg6p1rO8BZCRb/Yq/XuWSkHcu2prHr4UCHjrYfSHH
Vr2SH3xxRVr5vDEZcoX68kV0l1YBdDtKNjnS3VKLxAkQOSYiQGnhjfX22lRk7U9lXeR+mbfS7XBp
MpOXpqO4J14CiXA4cw8JL3jTiMYmJHbJ/l8Gj3LNHstzP2XWpFy5/OoHZvWoew+GWQieyUXsZUux
9JLhYR2VnqBFPx2PBGotb9Iu+YP9CsfMKpm1ft7J20UzvBL1wtCcXdq2nbQ5HLWFQ3aLHqAIsw9M
Zth0QqAWi4d/2VEogk5CeGIflaMpYWXDLdRmEqj6ehhDnPWPVrdKOz0h6t/OASvWHd8pV+Vld9Ss
BlNd4WUaHua3gGF/aVgDiblB663tXqssUPlGBJzTZMzfDvVcXHo0dW/CiSGPGpCRAuulzjaxStp0
/Oj6ByyW6ywzFqumfqGAWXEji2aVeGMBUj6QMaBl2PWgROXDW1v3hu5FaGaGkhut5lPAIqslJGlz
Qlk1s84IhLOUW+8SuEeoQ8J6MQfjCyo/ejR2a85eMkpV7G67oeM4qDduZdxJzli/F5txn7QelJ1L
bL/yVdP57Cruh6uw/4QCUmcctYauIeEObTsjtJs8fGlEOe0ZJLGEYNZ0L4vs5pWTetGsD0+Enkd+
2UlJ6avUrTk05xa9JVsW80BlW8yPmCCKLBtCsC8JNv5MDQYQzBUEfa/qPQ45XhKzBDJapchtMjC5
lGovSzt0eypQParnGha1d+Lt2xsXy5KuS8jrVEAFbxXj+ATqZx1mXV0GjlRabcuOMRGABvXbj5VA
wQ2t6c1Qnwqoqvjgg3qpWAvmohLdkoD/YqY19vQsdmz9qp0X5UbL9KerHFxxk0mUyWDaLi6ZP/c+
GbmW3B2h7Td0CaZV78yqmbLtV+qg8YNa7bW94PVOwL7IGFGE+SWpVP+I/7mcwX+lMHId2iw09OBf
MogDlbCoP2qZjftNUrlwpqVRuOx6KBtrzjmXe8MZUkcmD9216Pb+htb3ZKak3rEUHdcGlFX4YVAg
xKo2k42rUzqYi/njk7OBuv8PmeoaPDbLD1DGVeDUoSLeCdfA/OSAP7str19JFRZffZmVrJ/gnf4m
ERlqywp3QvdtfCSsb+MiX4JVK4w+NOWpPCBYYOTsvJgqcnltjiErdq6Zp3qEKygMOMVdYF6PES6E
LBUKtnK63R7EvDBVb9o2AYLYrmq4KkUDKsM9UJdl+Gwqwe3PlQe8pRF0nLi2QVSqeiQzSG8JA0wS
xQqBDpzMTe4fUdYWf1FxdWApL77u/UActncniqRGj8kvWpU13Z3f624zs/ONOzHP0iE1IOz72dWI
VVMcFqG0d7MKL3BpyOlQqDRi1vqJSLU/Y8lmBVCGT312L3XaIgvgGi4NjcEBz1a7GiIEBtudPgIb
S7MuCgvIYI25tjj2eVMFteE3uOp+wFIHnrj6uYbVsG9WeYygjN60zRI1GtLGcy/OEimAYap8UWXW
6ruQo2Eja5dlFHv6TNQoOoI6TENdI62AaL9FGUpQAKAMWPNyei6jo8jp1DbrqP61MDaMb920p/sZ
2Qubh/mXSQDyhs3IASM2E3uF/MTX71o+aQTapc3lfcmoKh5EyVqO6ps1UXYcVr7vfHp+Uf12Ew44
XC+3UDoG34QRwmAAiymSTKXd+ksBY7vWaCyCBXni0v9yh3jvTMrYoRZHw27SXceciZ9/C4B8b8cZ
yYVcCrxRzPsrKp1hAVECcHUftjnh6GLkSA1kvc96fXu8KJNQUbN+Ifz46Stkt18uY6SjKAm3zGFB
CQLMUsIKaRFoLpcFyl9cdp+GTVNoS+5R5lAWZDZwCnDNkNtuaa9LEeu5icHLY6QD15yL/XCFtX0g
D+hrysbu6uP1CcYVAc0Oymt5iuSW9+zF2UaQe5r8E8CJgNelZ3lLH5RhUBXysHevaMPXmgOPQQnh
98/JnzS0RHUJ7fjshvqpiFlVTuIsCsnkdR+4jFBYOgKRc4t4pt1mgtrpVzISEAmGfnkFbIPY66B2
xbmYv1FKMQXd407u1LgNmMEtkFc8YINFwvUR5SC4gx0NS/pi42MhxzMOa31IO8ZBqo6elpR95Edb
wkw3ej69PZs7ZEKOvnrlXkQVTRB0b8pmi7r3f+YJUGB0WB+nnYFk3zRyj/qrQs9VBbfwIt8cSGY1
hQUXF03RulUh7YwWLV9yrJO44lrUiXrXYnLF0HDfvQ3wXMAL+l5b1Cfjy1tWlZ3aaNfLsM/wxPzL
QKpeAk47R8Tia5pjcx3EjAhUy+SsSVRLOL3+Jd1jAGeQcl97CRJaTfxFEv51YvjWmWnqT7qbbxh2
Lcv+VHZgF6zZ8VkpQRO8TROURlsRacVVMftIfjk4ZAcRTlyHX+YS2sbEW4EJHkVOKn+z6DjLvxLf
lZs+lv3KGoz+z9BDvOZBqT/jIEnliF5vI22kcsmnxJOcbmHttyjLfuYMh+ps0FSA/WQYHbB6K/r7
LkHf5T5U5iiEYo1Cl/j3kA5JgiU+L30snB42UgSGX/FqYB3dN2H1QsoZ9g1U1NwtJrGGZc+yXPBV
z2rz9R21H3wOuviyImgQItLNvcJOGBXqQ7mofMPI0mfZamNx92FUh/d0bPABWXge/++DhnuWYZ8v
CzkF7+ZF9G4ncp3mNp/9YKNPUXiZoAi7/YdtSGJ7/cRGomrVebHWJfKpDgFxQjVlN1pQWpmVYxVM
E1Q2PmNp+h3+ADSqo+aVRnZH2Oe4vseUPsqvG4VTyHlFDFAUthWqRyFwsRB/KxTOp/2NtORjUMoz
jrtOg5u9SUvC9wPofdDAc4bdYHM4zDVpEOG82EORzlGFuviYR/d0YKWVr02hufh5c0wmr0OlF/ff
PG+bTnbaNvK5Xc27DWLQpOqRT7Ef7DeCiusGZLTCxkzl6vKnMJazvBi/TSw/0kQhu62Xi36bNk4L
TpzefeZHHpChErcT/Ixu+sK6OFGo+jUXUyX1qRc8LCXLdSx5KkYE8UsyUK99QhSfBD1B6ypnCSsa
k5NjAeHfseVgffyUsyrdLY6xMpYzdQVWDdqngpHkCeJpTv9gCv/JZEx3TQ/+xdRW/J1mRmNgz3h/
3ht4B6Blo/3qZ4rueRLqig+m8jOIGttaGpkrqQHYTHTBOh1JDXY8Ay9KlINr59la2T/dldBet8MX
BZW8dWNo9S1vSZSvMdoNXTpyzUsSs3i9RWVNyfJW6XPqu1sfFK8PvmvLo9P3eYc5pDlVmwS8NoAb
8R6CAjAGHTZBcVdvREiwzwYhe9H9nCTKrBU/I4ntsWWNUVj+/BFPesT2cumA99aTLwPC97sr7X4o
yeuB59XhWt6vpwEnO5soJhgRP0elJt5XStwZpxif4IL0aj84UHU7fU26pDbVt+QPk4RCmHfwXysJ
638b9mkMYqUHbzBqqg2dQMBI1IgrvdnFJ3yxzSjxkwpTQ7WKImtjEZUlH78mEVHUogRNxddGkY1D
3ZjLiZNpekQAaCU1WW4jIkS0OHIgtiOyxmPHSRbObTau5VUcUfx5i9mBmunidCndEyPgCzIsdmuG
zllXBJKJWJUfM+AJ8MaQwAGCJxbvgMZi+2ucoJSROuJ7zGqKCInDBpFrXnybc9R6aMYztfXg8WIz
6r/gG4gYfFdgcCY29w/DSMHaICtgyqpGsbagUBhUyOpouMSOmExVrmYA4Kx2SLoLSwWtBGhVolQG
Nb7tzD1PiXaKJarIVnl92GKLPAFhYKksJR+mqO3tDjp70IZtdvgP1WhTYvrerOUcKp6iw2MzuCJJ
w4DC/LjNP3eVz9nKAPUH+oxBeIZ0kqao8oqKOeKdnyu39acPy3QXe16AFfZ0jbmyKrn7KpcmUxHX
b7K8XYUnSA+iJ9iVeorP6crWmR8tByrUc7pJCeg7/mGn93DxrA7fA0m1K6UPsRMcmBWk88FH8HdX
9BBhYtLW+T1UaFaA71VFNlYy+WrD+d1ny0ZtGAmybbUpfaSMYMLvaUdzMgwq4+j1F0kF2FBO7aSu
8drdmmbbo24HLWnVc+UbHCof1H9wbZ+bNed9zDEjpUvug48sNfHKy0bC2UhlGlj2Z6YBTQB6iscL
erBokGhcEYYW/r8aZwa0WiWlIRRASkmliS3HC51K+YOo8ofnXLI+xhV2qwXMqjq+WF44sy84DF+h
9A7lPEU6TkMUlr571tQ8b8B3DikescSfqWnu5YvgueSNkGKdhFenmy5SGLQAVKi/plHYJ5bu+AJi
awV8HWr2lgqd/MEMysyIDQ0gPSPGNPzE5r6LTB01SOwxUCExSCA8113RDNYe2ESGaCyK8soUxq0r
LXycK0KKA1+X/GPFyY99DRjHpL01psZmMFpnTNlVolUsft3Hfeb/K4opO9ppOgVvE3KV/QSON1oN
rVsHgj/P/18qv9bcnHZwIciS6YnDpIaC7JNahu2ss/WKwwR2lYLNW0vMTCOTAsfhSLIaY7zxymA2
y0M1XiKzA7r4YN1+d3j2b6EVLFG9v7zNbCHox4ZrKjhw+9He/2qV24DAYbpRiuvpdr7y0xH8XaEX
X9Rn8kJsWnK4o/Ro342XA0hLsIVKVYsykGiCzVBEpqVS+YbDfotnowMWs3GubEwp2D/PAXcX4iFF
QKpU4Jm5M36JHzCjqAdTN0MarWrNQ59uIeMyNVCbRbW3nWFV5No0QJXJb5LQoIPsAPJLQs408OzW
eHlPpL+1Ufm6wEjpgBwiOrXTTCd0uU2WV9qMM8VjmLPOg1zVeop4YmhM2opjF5xRel+e+bp2PsRl
9jfRBgZliGnSx1nv0vYaNZ35zH43lf0Sz66nl5f50l4/SLCsdSFCztyyuCD+njR7POUITvuL7RRp
tlW33NVKnwaph91ty2o3aJvHDSGVQF/qFDwbbKz0RrSHY+iHe8DVC6GnN81IXFaI1q68qpFvKXta
eHJvBlQIuqJqAM1n38LESH/OgDPXh9WW/xHx8s+HmINcCEnFGXMK+zBieEG8093HnwzFKqW/il6X
si9f624IBwyzxOJ5ReD5j06Egi2HW94+hMM5ZUpTQEiZYFVkGwCVIGhiCWcn63KWwc9nEk5ipIA9
ghxPFv9RuGoe/960IiFLJLI5fRdUHxJDTIy9waiw81rXcLiOuZrVec9hO8gqx/+zqo5/5L0KTuYY
MX0S+okFAWAkBc2Qooie7v9rSxsBPUGR6cr1Vxur+IegXxTU5ubktrTMX1L46hmkgTkaeWyFs2Tr
z8WEtDQ1Y/S4lSHv7qCaB4mS7u96ZSsgA1Oe8SdlMtTwfaM2+2u2i7eq0eGFN3gKlEJKMvoETLLU
54mw3TWew7Zotq4w65e1g735+MncKa4OuYPzaHVVk7A5RrurxFM3L8bMlrrV+dhb0ql6mX7FAcX6
VraNTqXit7accRLnQeoXROTxL64Bo9vdaPYg5MkiOIWU2qnrEfcv+7c1LhgbEED1r/SHxlbiQiiv
LZqCpSDgexSL1O23xojAHPLWaV9zhuClB1BDdIkvzn1Bc7jvIubvioFxlYg/MwkMjJA8ZHM5oQ2u
5sYTY4+vDCkC4hhaEDMLoH2nG8djgHKi5OMVZvqplYqhpY/uPgdHyJw445k1VKyHCh0q3rDS1rsy
QPIHNane+oTpdorrMi1I86hWEG3DFBqpA+mHTfDX1jpwbKSP2KjrEgDnvtRiTcEDQ/Aob74+fzj9
z56tuv4CZjC+78ZOS6v4p3/vTabCejTZ/glU6wKsq/zei9njZ89u6hlsJwWucvobvldpJ2E51k9d
1T+UHGlsRFU36uHdE5d9KVVxj+6PPBZFXnGdSEKA2JS21P20Yr3Aq/3evNVy5iv8U6Gj35kI/dm5
1X2gOq5Dxja/ERaGlVUEqc8nSfRyO2Y2lVh2aV9ozf+fYkOsupb0jxnjEOYn6KTmyla9GsZXYlms
rF9WcPOE2YmoeAklKjn1HIbw1qDngJICIgNscusJevNg/zD5uOw7nFHp9itr0kgTR+zCF2YfQKnx
sRSzjcHdEogSoEEERyP6o/PJ6Eas3uPAs7785wJ/bg+6kDglGKpmyHo+f64L0mXcFJJQ84gXHzS5
xJiLKg5w5wZ7AWfUNYvErkwVnuOBz51NkNgGqCDE9nk7r0gQcKIxcSb6HSxeiborhZpiMOemgm7f
44iNMYMG12ce+AH0t4p4ifJfxgi58V0mDSQ6+A1czOkDpa7wQN1ZCKS9WIFN3EFM5wctRwUuaNgE
OHv6fQETyOHGeqTrcM1Y+rdL7y1QOWhtBbxdpBCjttcITIXFnq1i5ETyzl37GUwo89lpXdyOCzCG
GIxfZgLrE/k/JVcciPd1omcEorzvuSu1R+e4qw0Qv7nKzA7QejyVWuZywKzKHTAEi4wgEZn4NLYw
uwtrBiAlXUr7sg5wYMA+XhjjXz/1B1R0Idhc1rPHDucEQxcPgLRy6RiCJF22ioUeUWE9x4gHOfeV
BDVNFyqWOlFdiJdrazbSsPEQV/Ofsm89sCurlXVx85TuSxKV828WRnnMnFlLHDQra8tWRCfQhUIN
3PxowPL/Ym5SC1HS4/5Mta9trBremPViCWH/njhRPnpUaJNOiFIuQjK5K2eWeulLaW+M5WiybroX
1o0YnH3VwNfoZCRAvBm/MM2JifEcuKxynu6JjvKRPgTFxHXJDCG4YKsxNw/v89HIToZaArYWgudW
ZZKOR561Wgq3s/iNPRIC1waYWI2bYiBOdkMF65h/ZuEVk1l2HEF0Y61n6LnNyzzu4Qm+xVEcDXnD
obex0WKALRC7GZptKMCPx0AAiNeez7GOAH6nSFANm8yEAMGlCMMzZEvFy298qpBXhfhwVjGdr/+f
2W7SvqbIkOrmM+u9izK2P2h0n5a+HpkH7if8g4ZhiELKWGXchnK9xT63GXIlP15erPVV9+gFWQcB
+mYUOBl4q+KBMDrM8h3dIbNctDOTkyd6OM0QmtXtQNLowGfejOjuBRoCRwBtOxbvQgTIXdggSp+T
mHaw/rD0xGbhc73nvFcZQGj7Z78pm7DMKUuX9zWGlCSpOoCCHZtU0hvN4rZR+wzv6i5lX5fC5b4g
lpxz0fCcR0ewlwMdOFTglBpXbMQmeQ1oCd+lX9wkdxsT3LSqKDmz367QxGgNyIvEf1aXkE16JS7h
+iv2DqTC0O4l2dNDJI1/u8gXQMGlok5sCcufJS0xPCzqBbLXexGuVF/54RG7Ib2pqZnpmln3xfzY
pSLtuoy+hVKpEI+Ml8cHwM1ccTZzwGoV0XsURskY8IwNt0wp4xFCBAnkGbVl8u8mYfpfPYBp5BUn
gMwf+2aKj+/fEvgkp7HsTiNusZMwHDrAR3U2mWlMbeqsnulKHLPr4C9YTBLKnMTEEkwl42HTJhrs
95ez6wFDThddpORqUqBkDaG4VXEKXgDcCVpPv1jZ4ppuv7s+aS5pmzejezTaGoA8AtesiclEWPXd
Dxna+TEOjJcJFTfJ83GJdmKpMS4FGSo7oZbN3oeeyfHYPz1iUGZKD9RNbsv0FTqsendJ468KO3PH
rNzchQ3N1cVXYo4RPBZYzKY2qxGfTyD2zzCsjP/dW65C8cMfLJnN1CmY5Igiwkq015AtunC3ZAY1
MKZPb2wEp1PGnk7vXp77jniV2jhwmvTf8+zgl4vkk37h5iyyZgx/44QtnPHLVNxb0y1mNwmAYNTn
j2Wg3G4DW1QPihrgu58YOMmZlIdT+xtgURPAvKD81sLmeKKAZZ/xsVfV/DYjAXVwQ1gJnCCa46mX
1/WQSdVcsVJrQMgwWRvaLMvO/cdsvSm2902BeN5ebe98uFCaYmN+UjPbpXongXqpsbh/mmWh+qAw
XNNkVwUTwsvfrUkPMUjNRrEHqri7hi1m3V/z2U2fGRo5SvZSLxKlKMTsMI/gP5R+Vy8RssYVC3sU
JugT2RaOEHKSXPzXGwjB6s3W0hPN+2J2FphEg9YI2jhbwQqRvU+n1ENTRE5xkPT0HF1BhgSTKfg9
p2SK8DrLqjVDfqymARr+RY1D6rpdpk7UFv0KD2inxFZskzLtClZJFo0pZ0oaq6P6a+B7kiTm/aUF
6CYm1jXfglXTmKcwUw1sIWHx65xvHYXE0DVOcmo1yd4u1aqMgcScIe+XaskWaMv3tIXK0YP5Kvsl
2eYq66f7cxrthbm9PD1z6dvxCyk1Hgc3kWBP3Ipny0rrhR+pm60sYd/Ytnsl2DubNqGcHpluIiTn
0CvEHetYw/9QrGRKVUfBs64CJjHNEZZfvsmadN0Ao+wWMpKA9YAaEzxfykLnFqP0pNF6HpXjT0zq
5WrjFWXTAXTfJ7+bFgK6zM9ikz5oC5gIeSTBtY0oYRTbLzariR0LaAV3C1aJrc6guR/Q99dxEvsr
8+4hIxPhLN+8PCjzimBiu9rPar5t3UP4nFQdbV5P1ER9o9A6R2mbSCtSlKUnjhnOlPIza171smBE
rbi20mrfiSWIZjUN1+ckIl4n6/M1sQDnW66I62SMrQm6VtgoPStjLmK606KK8hfoQRiD1m3Bow03
i34yKvx+CdgfY50gCsedaoo0+c0dGZYk0cTT+jwiTPmUepvBRL81HCfufypTOOfzdtgiT0IHHVDG
YRKRSOKI9/KPeXq4+dI0/AK2Jnv1PvOj2BZ/85pIwggobLG/MRS4qniQjswQO638eaSHu2kD3r1f
bss6Ij40jlaexYlHliSyyA+7U486/393KMMGa2uHKIu8Ce+R4AkOnAAFJ6z+adtpXil1PlfiDefM
BQdx/4pC8Za8qTNbFunNePv6qTWj+hRpXmCQX3YzGTOC0egVXEL5Cz+IRtjs9fE7CxGX4GxV/5lh
dfVNb7nkw0DFu1YAhfh4TcEXXxeruHtUNs/C9LwS88ENYW/IDUf92PdkmOtIMcNwnLsegwy4KF5f
6k+YVGi9gw+DLcgEjSN7ZmhQFtpQ2bVIWDsbM8fsbaiyOB5cxqWVEHDTeBiu5ymMEQWoez3UU8Ma
O3PyTGiuUTDCeGDUIEo0gNEm5K5hP4UPiL4wcSLQSmrLc/RKeX0ucRzD1cHJT+Mk1+o4/iKIjDIT
xRom0K+D388O26frWBaeD2MKRVfV3ypLANAt5pM2PgJUDJSlQwtcO7zu1XfEfeToxkB2cOy7UZJZ
n4sO2VS4m95CFI59t6xfw3rHbOhUHuEBjQJPokpnWTnAX/fDyTXIuLTxO2i4zUK+ipoH3drVAjye
r7XwLvaRN/ZtMVgu/jXHT3wK2n/Jlh2j722k2G7SS3oCAW0B2SRHEyHzzXE/uSWneG8ttFBPdGqQ
rJGanKxMsAeRa7V2YXVEQGbqqvyfPUzk+D8UNoGGWLaVAxcZ0FQivIR1eWanOpt3GmR0ygTfndd1
ylGH7evSBOKTsck6a7k2JZhIGa1o9Nu3qYtaKySffQHGgzCoEevh2vj/3UyuEheGZ53CZ/wl1JUL
WRxH1C8ZuAZtQ4mPmAP5ve+S/9HXu4WHNPGKhzemHPoLtg4FdfU6v2Jm1nxgzBa2kDBcH29DOBcx
fEce8ctji4HO32EUK0Cn14yjejc1HoJ89tgc9Z6pLIoHawddbDve4buFFZa79IEsTwvD1O2AFBiB
ClwsOp9DZ+K6vv/B9/FVLbAB0gJmAWwHaV2BqWcNr0LbK6p42M0/OaGJFfDK3OVuGz7P2VMcpqnK
/Ennu6CvAh8KJNNvqqw3Re7/aE6DyDQKwp52QVVALCC4ffApc93yNZjGraUglas4WDD/a7Vtb/lo
b9TLeZ6h+gy6K1LJghqzs4dBvqk7v6vaGMJX1LnrxLZ9D/AS6xJOErzS1ULcy2aW5B4hQStCjNhn
9cXVJbBWpsLFApvx1dhUiHvfiFvdYzbBn8ZPUcEOQFWhrs9iS9zIPY4MaVpLzn0Yf3O8nqLwZEIJ
lF4RcOQPfIfptyvZBv+X6t/qJAQAJiYgBFSOwF52c0eKOfvs1yZU27X6WFgZR6lfU7Q/EUdUkjQv
/Lwc/jD/uQJmZ8CTZTGEORY7lFsY0KldR6XwGySDumIfk7EVeFNs4kKfYDnulkcvpOhrH11VQqQr
eODXhi7RLPghztuhwS0dBwIUnMfBvoHPfEEegGLn9wvsoJI9f0G6uIc3DQtjUJQKLafVLPOyPmy4
DVdig9fuS1wzBxUWBZsU5hcT7MCnWk6DQ8LLMuyuNnH84SliZlBRmxjP9KgIYOtw+NuIZNXOPCPj
OJ3nNa5YtUSscUvcD9WYaJRUxGw1m3zOngqzcFaVSCyxJm6ZPtVZC6IRKNChrS7K781tT+lTkdgw
k7N3U124ofGPMhlXC96qKEbKIUAOxO8oHtawV1EeXF2G2Fszm7s6f6pp65hcfessx9r7uv1em06t
7zFf8tbccizXbTwDObJ4bdz7j10SX+pt9NuZsvSMXRpXtFIf/2GIT6Ib12zEgvmGmyXS6bpzWlHx
FKlhDKDvxAf3wRK6ZxIP8MrsjAu86zUCY92bM1+PgfoNzOrmSV3EkaRaHv2cDIoKEz4XzSW8VNk0
N8azjoU0Lxj82iEtN29MnuPnw2b3B7h0trwKgNXRTmuQsbgsQ6QSQ3EZVGvRGAbR99KNEtY98e4g
cm8Up/3BqQy1sdEj4rosb7j6bx22fv5aWm2AfWmLNpcm9la2EGPNH67uv56bA6aeWT+SUcypaigr
TRQpglMAW7VhAUFyOaCVkD3P9KHwHCKgcKonwrXghwsbpkMueagOmN3auvy03i/jAfjBgPY5QzFL
CHEorfLiMp3G6E/k4JVEQqciq3H8GOcalfoOGrI/lfgkjv746kxU4mS6XMBYd8TR1mRXdULwyUc+
tM8t8XHmhhBtpEYqKjKRIHyGqZTh+SK9DsAvTjeBzoYcqt7BJ6V0uHP/3XMk0XYTuooMBd7GvIOp
yhXt6Gx5rltR1vRz81dm7JWypbamxMvw09Kupst3qfFxobtaBB8ocHCxcztqb9qqfe8LO79Pzgp4
KTyCOFce09EfWDmVRwIMj9hRLcJGwyCIYcoDpDJxaRly7S1bESzHw2n0PFcT2Fyrv524qeESo5Hr
PS1RnVBbxGSKP/oe1VrmkC6PuOSqQDruyGuWmT2vak47SC1NAiZOQnxL0zVB0RZlW0yLFfSwtyox
zAk5WsQdQgGb5s23JZbuAgHHpq7iMOHnGyll7eHKwfkJz30hyrEPDK+UAAsRz3p4lf7D+eE/UkYs
MmxoMOjEAJEFGUvCs7F7JMo/pqVNoJQFGorjF2yaZDg176Lcz4tEaHR70doa979L84lzBx1ctIh9
Won43i0oZ3orUGqLfJbrEttRQaLsszQJinYau1tZjWH/xVhjmmYUACvdyKUCi6w9Q24mqEh1dGX5
8jXpsIJKMETHkEFnaos5zdNeexetILodY2E9wL2a7fepqjnl4BkEQfoUGGRmGi/DsZ/tZ+2aBIOX
Jied4b5yWelSdNJbf29XhvnuGSkMvQSB/Eo3trHmGwcBMPLsetz3goqk5Le9JA98YxxLoGMHQRqA
fUbM13WwTJLHjNLpW5xQpKmU638rVYx5mkxOjJv5QQqQtmfmcJZ7xoIw6iShEa+qrWCfK91NIpCo
WKKzRkvCkUftmlHQcxYM/HJviuxYvxAzxdmSUHsOofChhEP4NiYxK18gTREoD6LF9Zte5eZbq0K3
mIkYPu9kv0fwUlP8KyR4YfbYb+gZ0sDtpCFm+bWdpCSaUdqFrqVEov9/QuhTY+lrtM0VVeUjbaKG
lXhaWyo1+O4GJcR010K3sfL+jb7hJNssNRyxLwFyBFeRYfEWsxUpUPk4fygh+CVch6sLxWqMm6Rr
/bPZ7xMYexgUBhsM5CGC9BIO/5WniIlB/tMQoXI7YPZIpd42CPwAltNq91i/hnT5vkRYpwsB8AG6
/I67IOFe8LVuxjRLbs3BvFFpHrACTp2Vru5lJKC05SOAgn7ksMPHo1QPLWEfbeN5/jASSES9mXuV
Uce4L857KqCLDD2Hln5bVxdA4tUcQycjaMeHnBa0eezJTTaRoyUpFudkHTnCoe4tV2aU4iLTOJ+I
kg++gu7yqWubsxZvB0xKBRUKppVUPp0eSvFxx1pcIH6lp9w74Td6GwzHK/jUEid40eQDDBqawwZ5
iriP7sPoDyUHvtv+sQPCBgwQAt/0+9u/RffNkHJ0NtK0w++CwaYwE9yiPH0h+pq6yq+olJzGeJqo
7bxvWbSoQTq6LghA/5b/nX/2B6kXhNT+hr+Q0F1BZiLVPaAp3zG+iZnCmQWv/NqVyXquszyUWb2+
dficDxDLXZBc0Z9B/+Ngwyr8YYBwoMiB2uXnlsPt/SD/riRGao6crjITEbtgTBH1yJxvbYrAFzYf
ao/kC7me9RaGaA6TSMT7WXNcsT7N7ZyGZ5FrJbNDHMIsf6whkxRCfOE/r3wvYezFvkdePCx1JBJA
5VAigVQ/iDeh07JaW01ta+zqTz5rqDHoKNdLBvFArrHL6VaaA6y/4P3n+dxJWghruYXBAWsGJXPl
GtI7AsBsdiR1A3nUJonjdJnTTJTb0qPDXzNOL7gB/2rNAEqR2D0uEf/0ScZAgvXMu0Di137MdsVs
LDE2DBW/pFOWK8Du3/e9AjBHR5VOA6QHFEnfJmBjycEK81z3w0DAmoiPiJMuReN4ETkNvW0+vP07
FQJE5Oio0hea1Io6AmkEF/EfhJHnr7PUjghIbx/knn4w8JdOpOSlcaHph5KKKvoqHmtNJ87DbOxZ
8qZGSbWdK3KOXK0pImBB5OwyFvVvqMb+M9PYc3I4g6CmahPC4tlpusChO9jgc6CRc07oWhvBXhcT
MgeEHteSVQRdrb95dAzBx80vNScMO6te1ZgXungW2+ijMo7NN+0dWwos75KIh0e78jxkXQTHOyXL
Ck3u8VAngmieQG/i7Qj0MBgJqrLT1lSgJvq1aNM7yWsn+ONDDLcCF1YqH3ZSfoonMnY+jv7upJUm
sPwdo8yAhTpox71PXsU3oquHhBnZo9QS0wEIvcA7KL5oxnTgUE1djF8O6WsQMJUtFb8B2M13NXyH
oKVoZDvmDVugMAazgSyjI1Cr3b4B9RH0PHm0rTaSnFmssSAM2WwMY1MPUoX1bXm2ZEQ6YiPMSQOJ
y3U9w3N5IkBHKWZn43H4dYUF3xdset9q/SFX1HuEK1AQwwmugC0WAXFYdIcVlEzhKYtJcji6ZNXU
vtX61Hr2gZ6v6+VgIfTfQghvEb3ulZuYBjU6Ude8EBh/v0F3nQTDEoSg+VGzd6tZlpi9xMvMJw9i
zUU5Up+7nOADKXDzK81A5KZeFLGO+zOub8JyJ73jAI4bD2m2aURxmtHKuHLdWODlCDfGSgMXF1B6
NsQedMYbMEKkvih/KE3APBaeok0hCAFxlNT+3/FXRs1NIl/w3QBvKrPvFSuZV5wTsPFCZcji06uc
7dQn1bflxdQmAi38x8Gf+6oym7LAcsj5j8Hx7RKu0Q5UBqhMgeGzi99JgNK5jKG883qpMhZGmKq/
96fmTCjuURXproRioqhP8zakJ6FFlE4kuPeKeam+GATdH4F1qevcCuSApuZ2mgEwgofYk9RlCUa0
Tqdl9P+uJFFpAXAdTN9vg+2o85s4BRL9qSqWiJSwkaaYJ5O/noe+4IYi3le1tZEcxUXX3XnTu4zG
Nqm7RJUjA0KskyqL7NDxoMZvFBUW64ul2j68JkH9NGatuYcMzcBzG/s9greLM4n1aLD8y1MB7zU9
fgiWLuEFI5PEeEBuKb5IcTiGpY0Gv36iTuReigHWJREWwrbrwsgRU0laDGEcfoJv/NnjCfEhgiqu
3o4Dltk3bE+UMmU160qsm4YJ1p+8oBIsaSPphszMXyiHHiwsiZ7pIbANLB63TPCcSeYgzgK0GbOB
aCbywnvf9T7HAfGAgqYbVeP4MX+2ACOua+r3HSC4QiPSSjqYsoU4paP1gVVi3m0D5UH/1vfxlf5f
c70iu0LgHbUe6IEZVzDKuv2DbXU2BbC+WoBD2+XpaK+qv9YgGBQUgvYP88poIfz+CzYvfOJbO5+j
Si/lN0puCLyZcIUO8k29F1ijsyhPIFgAeN8pDTVlJGqODKn4gtv3jRlqtgOUMIDjE1vsYdWRbKQy
yta7tCloXoXKV0B2/XNlSk6SEwZjRDy6f0RiX8SWiZ7wIxPAc5kizIapRLPFQTzDAnG5fcsVnGwK
x4tzkd2lvtnZ+KelUB2oCtqxrZE3vqynSKhl2KhqFynG0aLcha252yVv1ZeLiNI1dmBlT5AU5EFG
hV/keY1IbWKvFRAhz1wcQZ3hhEyd1aWljg46nIYOUn+83ppN/+K4DCkpAoXA+TV7uR5cTRvGUdRE
CJ2+7goQh+u6uROYcqJQDyicWxXqmIb5gLvOXjHu5WYLxEfIxlCdzYnIqeXSrx4OS8ggVKOdkBNs
TrVvfHKs5gQ84IUAbZImrzxR8YWzZh7LxHdjezeYs3pCLZ/T34BBuquXoymLEfTzZfGN0Sz8jbCn
AaSUkPvVIYMgr4PqASVFN4yNZcxzE93RUfs97SgYkPLTkpb365su9jzW2jg6PhYBV06ZVAf+CFDl
ZVgsRAQ2kDPzt0p8jWGbEJA2BlyNLcf6+qquLrprEJDm86pGAQthhoPfFXQmRIAJDBRQHw+HyFw1
ahuXAzR13Rli2VucQ9OGr5lQfNxNnlI2shbWWEn7FuygMsVBd2WU0Rs+mHhjCv+K6GdNOZXaDwZi
X3Wnj8+El/wnzgnkWNO4Ac8iI1sJDYEdaH9p6+QJ42vFwHqlEvRa7yuP1PeIYN1QDH3qcURh7Fqs
WO1PYBOcSl3OZTK+rNb5HTwZPtjG4FyNm+OF+B/tfY/Zp7IEy5GBVa5hqX+lXQs7i14V2bSuzr3y
OOTsqHXOlh8zLgKtANhys+L4YE8vtKtKK3LziBvnFGFBbck4wypVwDnK/KaaBqouBQkX3gCzMetZ
MuulNP27VGbDXifHN5NCzvZghEgPxZV4pqNZaL/QjvZN9heFUm8Zs9GHv3ZmLd/vJuE3OeL9SXs4
C/khYlAzZkjN91+du5KMIvUvsjfpo3KBENLT6G073O29JFRplIRjQc4tgjbVuEKsIwmZWDb3tHE8
Ls6R+WU2ALUeByFNfKOINohbAALPSovDWtHVZOd0Jt0/eIqNm6ObF0p9hgg25W+TbvpqtlNQL4g+
rBTm0/JLKbR8LwHagMfsjuAEepl6mDFodY+yEyz/rym79X7dohknpc/XHpL+8QXXhLjmpVwEKGYO
iquVmMY16PxCGb82ghTIHZXhowSQD2UsQUzj4r0nYpKeQtJcIaJQij77gshRQSgAa4aT4EvB+95S
wfNirsSXRsKZrvfkXlJzhXsxCrkStLvGCkj17hVg+6F5emmFBW1SXzI/ASdzLKdH/+V8UKN2z/MQ
MMsxWI4Fqzx4jkUMMKAVy/o5UiGrxuPBpS5vMwCGi16fKhGAgRNs+noMfuRDbpCfB+QO/NG+ZVWu
oUu3ybTacIZBS6/KvgBiSRhocgojE1+oSdA6UZxLOoOPdJi9PFBhzPT/z+zwYx0Dm9Lp9n4xfpXy
3SFetlcBz69pAj3tqGfCNYGH5t+D0qWRZ1+exrkxqkrnkN73StDKAiyhKnX0hHsWmEw5bVyIH5uR
JN4GIKpGyv82Z+7Z7/eZJeOEBXFQ92arIumliv8tfPgnXjhBGwMnbN5AEy63qczKGxOasyzIhbQr
3HyWa51Ix8VWPL/Cc9dZdZMP7Ujb9mdE7ib0daIqOWknjQffvywYXmpbQ244JpyCyhuVYsvO0AJd
TwzAb/mKQCoi8CYLv3ttZPId4GGdDhBuO9SJvvVXfTePWzmUd14jzV2YHCRuSS7BCA3pnZSrfiq7
ZGNBa+XaGLppopUzFUZ16RmkdS7whq3tgBsZn7w8oNjtelAP15LYYUoEKPQCeRKdypKZo5fxh1Qh
zusW2x36DAb5tBTRBXJ0bwwymwJP8JKBGq8qb3cplaK9oDAQQcp0FLTwa8woLYIBCRv7VlChyVy8
KvtSdiYNGkwKmYOtVz93ZBRnWCXm5IWaJX1E3XSq7K2rm+vGbDHdlHsPQyC9WwqJ8z8jaS6uevVB
EEiy0SB9E2qa9zFUhxFIty2/xJrgIlEJN/H6LaoGNrouFdZ+PGEfdxPNBxtXmyZALQbwoYlauA2a
DpYkCQ9oYis4GqjfH1a6mMyBJFEakIPHDgV4zj5IwtdbjsDtzmsdL6A0MBmlmUxAa8lXM9khpGya
xBQ2c9rgoXxLKMCWODgAfuGYdxezEPnfJtoEcA7Ipp9LwY9iW/OhVrRq9LrRjJwrBNcQxRdrlxVj
oqtVyvGm2uOzlcv4qX8j0U5N5fS4CWh6TJWorHD1pOJ6+d0PNCPG1tFoa4w6gzpS87qaE3Oxnmi1
Npbe4qvhdIOtp4qOE3Tsn+/ZFHozFM13dn1lOYdPHqaUHGGL7YDtoBIkEPHGuIm8wl8rpjwGMApG
uCHFh1OsvPh2TBu+It62390oSB+5ynf5/CXpz1jgMjVnZWqpkb18DKMNpKjc9EBQ+wG2O8Y2vJNx
Kn0DtIo8T45hsUQ02moNpnCI0l7Zqdzs3nno6BKqTX+2hAMTmZPCVu3aVbNTVcNzRF3n6629oTW+
h2A6mL050ssK9+fR99MBXSUMPFkwa/9N+rTiEDLDPzTv0J9BhULPWiwyW56q9yYte2YP4NmIg2Er
TsEyChwodSis1DpjbgggRTkbjEGcT7jnVCWCI1DU1zUkjMT/qvc1T1J6JacaPNJt6+sW0aPLsg/U
xdsJsJN0EYXXApJtwSdQ2X0vKUg7OOVpTs6XMFTcwwKAj7GJ+MDuX704ZzvU3Rvn0daGNu7tKiXw
sRfZXyZLq7g++45MWgV6/E0uop3ni7+rzOTJYQpCzdbQP4CTKm4FPLl6bsZzDlnX9Xz6ES1ADBdn
xS4pty5GTqGFpYyhJt2XhGBNgGsuwApkujoNdWIfPTATsxSrmDtVWMvbZhT+dHu1+F90IKSUjFVr
4nrAs3v9YHvll6ksV+Hq+r7Mqnzhz4jYoYIWEoAHkEDaJYDKGVDmqN/eJCMziUXqUSZ4MGM+PmEP
cWY0K8tYdt9EtowWws6m0ciYZqaV/a4pQpk+N9N0do6oUSaNej7w2LDvBcyI5OMNqptxqZ1uzRHE
VcwsP8Q8HtnTajZYzKRxZXgS9XLc89H/LNJf5GVPsZVDonrqpM0vrlssCgapQ+LLrQmqIV2BrkXS
qgQNChZiGe24KMyMkDAZs7hvIz6te7hFEw+z9SO60P8j67Rdo7YxYSNDyUeZ5FY1Z/fmU5apPcrw
Gsn6Jhn2i40XzL4p2cf+TBLXA53YOUHFL90VlGDY15S1bEZPMzOVkochyWphtdUCRYQa1/7U/XkZ
+NHcglKg8nPiGqbPVHcN93istk0TY38UzZJajloXczbbw0MtWNRs/6k7vHZI4od/5xeOHFGvKazg
mhm9ZJLgN8QZHHYEf8J595FWOeak2K9GejS40Rk7zENV9D75Lv5IS4ZWNB88C1KlXNT5f2XG4fXh
XBtmDsK4Hv9jJ2sFTZRo5KzJdeIJg5I1BCcgbMxf10cXw8k1wiDv+vB2XnM4gZaaWKeOxMGiz0EA
LJDd7a30ep4r/6B1YXrkz0c0oAz6Z3MqlyEsVnQpqYraCQ9OuNci//redtK17gwhmoNsmjCRPYtq
qmYBbUXPO89G6gq/C9+A5c/JJaqW69m4773ssZzj6rpsmt1GYg4k7x2DahnYKcevUXnfLo/8pVKo
IvsnBzG5vznhOFUzTH1ht1VN4Flc1fySA5ZVvW1Ah+u5Y2+QCZD7t+ZJF3mWg8Q9xdRNk0a5bVIh
uu5tDz7ekRBMfCUYItDSnfkYbWsx9WHQtVsMdNje1FL2I/4ElalVAcDjt08xqdbGC7GR6oIsYzS6
Rrl83kJyZK7r9YHYgOwRZC5Hj7TenHHjWwb5KCVRQ0xpnY+yRdMMJkr7i3Q8hcN/cCTialfXREOg
0x/IMXHG6fYQ1mhO7A9cunYXYzfL2u83wsXmsKXTOji0n8la38RJaOpT360YFnT1oRAUXpMayYhL
HbWGNLdcD3oVpPGqixDx7e2ozFC3eib/x5eGqCmjGVFLD7c9IS1wnCn2VKmNN4U/Tll4lDppH6Vf
Qlhu+5FMs4D8niEtwEKtIIy9ckxs+x8AiW3ikZBBmpwiznJOITejD5QYHeHzjRNCZxXnT2zHwqI9
ZtHOyQ5MhjKgLwPwEZMWiZ5djnGufWOzMH+Fk52eLWP1l3GQKWTuWFPUu44LZsjFcns5w7dVQXnN
IhVOgd4slix0XwUdJ8HPrjOGtxc10BmvbqCAwz/eqF512NUoi5oDBO65T8a/nNl3mvrKuH0iKhhh
n5XPMXYEIFlju2Xaw7/6D7MyOCILF2JpPeVLhHMsyylLutKebtYV5rnRVwStO5jtaX0aqUvX+k7M
SfBgErw+bMjJ7JfxsK/0DgA7NpbDz3jWsOkHCqwnCU3o4LikanyWI1WMghFjBPpYDv2uRasEKs+O
OGRN/UIl09wxZICw9tPnvY3tu7gh9JsWuVIt48lGroyQaUOZDJxd56cB4o+ZfHw6PxoNK47jzB/D
mWZC3pGb91FIIr+XYYm3W1mo8jCuxUDjn3hjLVzjBc5b6wH3PMrNTLXlXEJCvTbdh1sKmDMkRuU/
Wz7VKLulq1HOXjfpm8gWO9HJ4KO0UfyjqrVZlNVnZ7c/BrdSGz2TeckWES/PCC5RHmS1hSWjsQxd
7KdhpgtOGA4fxdrmI18lskXqRpCP5hxkNsw0iHdYBb0xsPYa/KS3PuWia5QIk16Jr6S5X0kNWki7
yh6NtkptgLvA1bW104jcAGJ1aglc/PlezI6Xe4ocric2ztG9dJT32148VmBLlw/vxlv3WZXtYCwm
c8+d6ARGSitKq9lYyGD6hJNubdAKsWA5pgUTtRbcmAEZ+q6wznCy/USERjouhmi+fOFtWBi7Eh/Y
i72GT840GZ+3zMe3IOwiWL9zc0wn0OZoTSNZoanWapvFIMOUga3KS+IpvciiZzIE2piWTeph4NvG
H4SgBRUktBLpL+Rm98e49LJCsrg8YFeF03ymvBkQtYtujj6QjPR9A5a3UN/UCUNJkGscNjJfG9ws
h1oTK4SmFs2x+Vsa99Mq/KR4AxUgJzcOD7Zt197rHciGF73PbIyljJ89bav48tBRPy2mIPxMB1k3
E8mcRysp5iDlHk9DucZ40hRZMd/p5kBtlH8HkLL1fbhic+1nVwmnRDH7JaQF0KLCcd9adc/nhKoR
G/7W+IPxPJGC5wa70GXoSgCpq7+e40uWG2apD0v71qgS1ssj+4TUAkuy62LQ0sVat+Fcqwz/eFn+
WpaombU3nfYlX2EFcQdo0nm9A2ceiTJXFS8sj15bzdE2RJcD0iuooRk5GshVfAxM5c6lb403TeKm
o+3pKCbbuzpAdri764gIc0VBVJLQ3HOniCM/ARB+mNaYqcZLQHIB/bfpw4Sbt/qpipcGTaE62CB8
/MMTWhdNNozVCOaqwYko5RBnOYFZwBplaFUYLQpm578QXncauNTMVt2tk/y8kT8EtAkb4VMM492D
H1NYPatd8pbibEBEgdG4xuVzkMMhlowloREHlqLZ02+kSK+StKS8VZlPfo69mStZgbxvANqX0CH6
QUWyKkMytz6LiS+k+A5EuUlEnb1sOVch8vIUY1srgvSJYAxuv5AcEviskE+SdKtpohC0C9wgkvHn
D0+krTdXvi7Z8Dh9Mf1PZX0tg1rB/W4dd+iVFDnOBJZ8vHQylsm2gptNoGHBnzJZpSViWZmuSV6Q
kHSPl/E5xdysaTR46oC5tebWRz8k5Ww28rkNq/Nt3wWHmR5H7Z5accOjqQ043huG9TMyIq6XJ8Hw
K8uObcLuoVmlXPJJ2WoN27zZAzIEcJAe5ks4gLG+5g0hARIo9WmWHUzy3kV/HvWg6d8BJt2L47H9
+Mf//YV7eUprMHmSth/XrtEqaZpuHn1w23lH0qgjQJv/qOLwawFk173C6i41jqfXrVDkBkPybLE3
bxaUybfDMa8qhqnlU0hvjmJ/Uu9IcuFPWP2QY+2zZyAAU7myM0tt4HLK8H5aeA56KSLUT1XHS7co
/lXGFaRi/aHeIlBxo6UV3xCwhss/UT2pTrxvJp5+uTyD9z1K/MrJMRFltwXouZUkxSdjzWFxKZzp
9gaxI9ZJZ3GDdjyPq6PSFdWO+KwvrxaNmzph5RM3YnVoiHLxgyHcxgcUN9C7oJuOUmLTCQgn6hxP
qhxYCrvHaMO2YPuxUMa48V5lrJrZa10sdoDO036M8aSJd9OKSdXYxDJVcHz/ACLeKxP/i/dIEdST
CvPoSfcSZnxuLtT+yg==
`protect end_protected

