

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
PFFltKdLY0A82yxFqahMaWdN+zxj5kThYAcsDyz3A2vhpKKQpGJvV8/AkpYYPyltKlIzJB6Md9uF
AN2ca05J0g==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
obdm7XtHPDQGZMrK3kNZKnRt8ypfk4aZ9VtSDpnSwNdbgwrFg4uylDkc4YjBW8BFR32vEdXmCKFe
3L1bSMhXRkPXZ88hMJlBty0IcmSYNatn3RV9VG9yYtXM73zMkJ4NIx7KoDtvOCnGQpHNAJTknAv6
BNEUXajqHzh/vB/QNBQ=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
nx2eU410BtrBCSzpvDl9pNpIplyp0nHGgzB9LvwnXgdhN5HNF/YNjnH8WXRfWZhIT380E9zFeNz1
cIYhUxogcuyFP2sgar0PDv645GG14wyLd7prd/d1E3Ur29iNukQkz59OjXTEIN/U9Gy3hPt+oLVA
TwpP0P8RgeQqCkJY93IlvPGfZ/yeDQHrxDZUMFMxHHI51HM/LG6Y5RjcVEJMkX5GTsC4gSd5fEHc
DWDREOSmqmG5Gmciy22xZEiB1SI044vcLqlJadcUhINRbAw0576LfZrf0pjCGq0s1+nEKeJm9MeA
baA5VHd6hhXLwLD9jRkKDvFp76mdZ8cpvFpcXw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
my8iGpxybuJuMik3+8MRqWVv3aAmCE4oY3Ij0YIUQTpme5jJv8e5DOlNoLmgXWhUlepBCUyZ1Ysj
JGlFKQ8MBs9R5aa1TLi8cCVfI579Nm4AO6VpackDfb6c5/BXCbiBb8XeC9Q6z0hKyH6xYDDC0Z7w
m1jdROr8ONcmGBJr57g=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
pEGUMbCVqav8XqUNf0y2o1L56804gb2pssAnfqbrEzVo5CXZ9MmyISfyPG7HY7huXkJ9tWIeWtYt
bUG1XTbOUAj3uDqhigkZ4KnTE/68izmD5rgLlGDQ1sI7w5GLUgtjCBINeZsiQZ8IbdNK2b2sCu2x
1k1tcyPPvRv3myvuFaOhmiYYyCNc8F9T3cW6mq34yHrMb8GcN1rGLFkL16mdIcoRSSN9znhYYcLe
21llq9uuuR5MD7mOGEYx4bKUQGVdPOHLC411Ms5bCd0IbhTC0qWispRkmO0D1uXT6TguY5Z6gKTw
vMvXdJYpwStmSqzikX3kYI1zljpfWHQ7HMzzTQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 66352)
`protect data_block
Q4MSBFg50tnSsfVlx0Vg4myOvf8HZYkrf1DhoyS1Fbb8WITqTFNL2T3KX742AnyiHi9XtYwY+iCv
nFcMcc9aRGpUd8fkGif739qdeNPBGmRo+NfyTD9TSdzJlJHkFHZlcLWNTtjkecYQiULL/w0PYQ5+
pZh1iIkFTJTWRuTlGpxAMoNFVfB+9VJs3jA/p7q6h3VHXXx+WfcFDRTu0iYJ8DWM/hNqvqJNcOwQ
hqnKdXW1WFR2GR66y3tw/aqf8SV1ZzBOdWwZOMlOQpJlPJ7vku3AnxT/JaYaG0Yk/C9SG49CeRYy
ofyZ3cvn4mqWXzxgAq+LR4c3/gGB+G8GRzjTKuNVo/qJ6JHxoYi+BJMSmBjxAPIQgMxUKrfiOfiA
Ww7H4ilu/BoJRRo2qVmBm6i7lbgBpARdsJABlSSBkmC78PS5NWJKXWFpa7TC8GKPeQXhm9sC0O0P
sDZJvgluv4g5L9ovEmTTyRj73K3GqYYYG/HNZ6zJ82eau1v3dJP48sv/hNaoON854ehyhi6Enbqb
zgUfKwycHOgy29xbWX4RrHZLSFWgZozuF9EHTWkFll/PUoiLhl3OMzbX5pqEJMHc68yp+Ri5Hy1H
bjYYPenEouSsskOT6KzmMxOBFL6DEj0QzYuqYimUc2SGrJUGXl0+qUaNFowataHj4ftJFZD9qDBe
hApbIeKMvFpBQei3X5PhhTgxU00G8PPs9Axm40/gzB46x1duy33OzxYeP9XtHt6c/D58NuJQTCLc
v4Uxb4zylT6eUv6x8GJ2qb1SAmxp2eatNfEMYl6a9Ix3bjQ592eh6aJmxBgfM/C3gGWuwuKc1LXW
+hZzTx1y57fbSV1Uu4cdfORTp9HuTAnPTwYPXOY10utaU69DipU4gCSBjddTfEPekm+JG2i480Io
Z+NyKskBUHcwswB7apOS0Hn/d2cycqqHRrRHUiimkGY7LH1KXVuT2hoKIEneZTNL1l6sayF5F0sz
O4sd8on72Wn8dSxRyu5rNvwFX59ljzdEyFrkzcB5UPeCIm1FWU+Br6vKxulEz+fRMpjjFb4nio13
p8rHnGGjImUlzcTJgLCQfATvGOmMm5r/iJNcd0fG/YH93499eVcar4V5P0vJ1PTnyRKQuU9sHJgy
QEbtv8pAegmeUXPKiuhXXIXqruA3QzBaOeaWY54JXjqUwW2yFniC1v+NNYUV7qfpXWtRFV6CZNRU
t0P8rHt7S9iPC3VcPXH/TXvPdSOjLMgZ8yayYpwL7dzhbxTr599xvQxKxNTNO8OlMAqKKr+vzhbB
wh8EYqzyzamQT+GBUFjBESO7MdQz4PCoeBHEG1wAy5MRFRqAQQHWP8As0/gw6D1sc104EyDoIlgH
oqU1r2+lEVj1Ja5XqLGdzLFROXGonliWFiRdemxDoUWP7cqO29rBWJ4Hk1Dh/ELgcAgutnRnKLzN
IeSHDE7dfRkQgO8PCg0liJnDXKpliawdjxrGTRj5H79stfOlOW7OqOjlr0zdcfCEezz0Dv1RKEqb
UpPOuZ7NdXTv8kpYiQwxl67K6wvMUvaqZhReOqj6GQTt6LMK37dFfOuc7PdMINC1rvxcCNrSJKnl
sQcazpKrEaIjo5lalqpL7Ithl79V7x+INlP3+7Ycc3h51QFl9qwtqyavihOA7WI89DCwbKAfDsrA
iMJbLE4EH0E0X7In5jYDRWZmAB5BGSESPwh7g3gZjSXGiyq/4ePp1KbnfkgVvGAL7DXQH+Fc2nWO
XsuIJtdEzufONRbFXjd2NdpotJg9+HflcY168xLk0YDfVqMXXoBQKheJDnw1AxrpFiV7piVJ7pKP
l3fDUrhaXuYqTeODdyy6OaV5F3m5kndwmuHGOhltlGtkCHEtzCwoPxb2NQlz3p6R2HD65lWgZ4CY
6xPVcpkTw5IqddPbtSB68To25F5cqGK11kznlLZcc4gLgxAd5rMONTrpmXieoO73QMJDLX2gAiX9
vbXOxMuYrVgtqrG6seoei2+0scbQxnkTtKqyfYOJ4449MDnHqsgNb3Xq6NW0JHck8SY8cCye3qah
j2daKyi7t0n9rgzyhVerNib/lzJadorcH8rVo15+DVV4yqWRQNFnfUcKIf6dT6SCrbp07R3qae4C
cqDNPtUbtgTuq3TkUJBjNVoDR/wbYK9HAScVNZC1xb1zCUV0qkt4xPboiGSIFWqaZD1e3S2RI7ns
nfjvuc5LsXrbAKb+HiZ8Tt6rhbKz9UYC+hW2td0FXiDOrGFmdFjSRUimfy5b5P3V7orDodFXRkhV
ERKeGpGUrennuS53B1LUN/bIBGZnAgDm/L5p6NTpBUGjJdUvhJUSGIuRKraN4Qu7shvZAhPwqufl
WmIdryjIkBBS782RerFZMXFoSEU+6HUCTjZhyhdV/BLsBdUG0zPR5GYaIXH+/j7QniuWiOJvL3F4
Q4+OAEUABpyxX2zs/F5uyRFFUvwUx1HvwEeIkHg8x71uPqh8uI7LiV1plBqpnsf+PKU9TenUK21x
uw56U3DuZ9oEM1ITxnnSPrq9kj5HACbhcYL2GvhI8h5WFWQIe0vkapipsg8lH6D/01vhebtzgOEt
Ad1l96gliRPE0ZnHcGnVn22Lr0jwC6jLqSCYUc9t0Cp2ljZTBmuCeMbWIR8NufvIopQNRCW7bjmJ
F9S5O4/DpquCM9c0JW4mppJooqDqetSqz4z1s0rN8TgHTDDrNVQG2DEwU1bQMEj9mjUJC9Tmvcqw
6zIYV/hFJkasU8GS7vq1Xfb123FHq/KMDDrm8kQSwkF+reSRI60CYY6CUIEXWLXlt9sh0cWUOSLI
Q9qdsBhNb8nznDIBQse9fLjhUSRa4V8bQyDJ3giBZbSejCoF4Y23/NMcrBnchRWezXp95mkn/w9W
JNJ2UwwGJy+gw94bKUNTCqIXOr9Pp1nazQenHj6508zUJAunHlUhirYuc+01LZjKS17vAX+LylDs
ke8+FjTk7Fq1HDI4lMKsk0SghMJhsk5Yji4mg3dwymrnFDMdNSkl2Vj35m3yopJ1+WFI1p6spu6m
eMUhcTwhVGF3GONM0MwQeub/adWXBjrJdO7GAW9VjSLHIK2wZSNxuzKvxmfQ7+G/ZVjxKVrYJb7V
q//uaP7LoW8NB4UlT1Nja2iWzBuX+SrA+g4J2yuH+nFr27P5gnlLPDVyVtppzRq1YEYTm6o1xKQK
F91GW23FK1s7Rcj97wflbApA/cTGj2RIThurmoCuBgL4p5X9A/uS6Se4iNsdGsVPLRE9vmupVVaf
9ArWxm+s/CXItuGEavZm+PsAHwgyzk6rTWUJV8auf6+tk5RUcc/9Qead4fflYOspGt/IIqONyOPo
UstjzASP2nGQ2AtSAe2+owU0qkQXPTX8l/ee1fuPWtjSjvI903VtY3oOXQLHoGUQNN9SNjXXqY3i
RmOD258KrJnJ80zwHqMbVxB3ZPaBd6Qdv/lr9896Merh4zlUz0FD1mLxURAUKdYJ5KTGcTZtUVmR
ILc8NnhUsy1o/d46GcK3z0zE0+nMjrPuAOKMJeXgdCN4LxD8z3ZaX1YYNgc/MdHVaEGe1xYLSaxo
E2DF/CL8UcOl1LBAXSFNzrn2NYOtwsCXkO9w9qN7lbyVz1EbtoGJfgqLZacZE+YOQTIOtS+ce4sM
zf2XfZLFd7A5EA+s8ZkmN+HruA1R/5OMs069N6VOcUfAkQxD/aKv5e1JjZ+uFDD7BiddNHVjZOX7
Njew0e8weH87FMItSDyf7axiZ1KyFwlLBpHKXEpp0V84u5xHCmvWY5sQSfo8XCMz4fAUoD4ZPj5z
exHrplVh4aAwvCtW2lV2B7TILO373pE/EUJLzgfQiS9OX9kqrPW6rg9MXEipytnLX14tKgRivyhy
zfzuL5FYhSIsELsDSETS/bFouO3C2LmoRqROGKGMiF5Fscu6yiOyxRa7Dl1aPTOW1GCrOKPb6yeJ
fgq2svSs3ApXZXpcwS2Q6/TRMEQN4EIrSd55Bu8BqiBY4oG7C3MlBVavECRhN7bZrFa0lHUyBEFY
wVdvjBWzb0TfTT4Oz5D6xGjyo34TZ1WOdV6NaFbshRtoanb2P+opIHAQWzz6Np5VYVgfqndpjUsl
c5aHDB2bHR6QnHxYJ1ar1T59B7c2rwto+5Y7V9ZyOdbZ/oGKXahgryW9f2G3vExIyCmnDa4Di7Mi
Hyh0yNc2w1j4OFohq54O9tY6e9rhgAo3l4Y9Spv3RLTlxRv/e4lAwLPn2PTQtea88koYjFSus/b2
yTGgVYJNrWwxjBIsCT+knQatViKI+qIAuJ53gM0lkCbA5rgatWMhESiNRGmzNWIvaUGnvdd9DFJL
UhjeG14IDxUJUAsR4kACT22gj4QCGK6COT5BpHr/P3Q/tU1x2qQUkM3dZgd3IC2tb0ALLt1syGZn
7Haig52GocD3OfEIQAxv4p7Ux4LxtdXPryJtVcLs/08CWt8olrmS30StLXZXBxgP1RlIPTqdZdU1
cELLMSgxe/44EgsfotluCZZxakoh9Z7JneQBL+LDp0m192O1gGs7CqhRKK5vtQU1gnd+Y+NIuJk1
1Enk3fbnvuJVMp4n6nCRj5o633EQh1cyr4qlUzJDq5E0cmeq7PlCci3T5OOY4NHLzmPtMvl/IiGF
rPGMDTLUabOBkkg+v0uttOfY4n+hBsYF9jdpppNE+MEsbg3vQghWRDpLw0KShpfcbprtFEbAqrvz
f3Hgf05E9kWxPnieDOQsuEKiyaN2o5Jr+bwX08bQmMH5SkmJKUZkz+prCNP1ys7Z78v0enTa9LOz
lkQstHg0YPUa7AMBOuTAX6kxV+SHNni8G8D6fmtwJyCdDSdUkz4HTwHFFrqsBgm9I32iRXkfXJdW
8grr9LSyc3Hm2C/AfbZD8t1N97NwwAel0r+HPh6tye+alWe2GwYIZe7A9MXDhck77ia7cSER1Jzw
jEPiW8W8xqO/5jCIT+nP4JJOm0PfeCQ+C71GJjnmd2Zge6KPfUE6U7R7hwgaTEoFiQrmUjGGCShc
WK5iIO2pXoJwoN6eBYpTw4jJzh402VYkU8vBQFwIahyhDtn2qyn+upR/iifIpEYfcl1QyS7IUCLR
2fYn0UIc3H9gdqHeif3khyXNhRoDETfQM9SVlPe5W9swZamj5Nfk+S6yvnfAoXWrQtd21yN0Meav
i6kCnuziIGx8Kw/tp4h7xOS5pdc0e2ZzZPSGlHW//sx2hm0gZ0vkVYssdEhIAk509v36snb2sm7B
EA+hApB6UAcHg1hcOJbK1BVB5lx8dpSpxM6bLjiaA60LBhn2s8HQmlAe8bKbwKE+rbEuMkglEZiq
t/Ohwvg19AgRTPCqupSE/Dg5U7vJ5rv0G2cZclfP51vb0Xj8iYSj+ipqT0NKdXGmK8hA2Su4UTQW
ldEaVgbM0FlpzWgxG73kZBy6XTyuOszyD/ZAWSGNWawMRcegUj3kL8d9FE5PpKcDsiEf8SO/7F8p
6+zq9nLQQgNgD2ifvDdIkr9XEW9wt1dWeqbxof/tt3wDdNpuvish7KNAwdMT4C/Xg3+uhR+1XPLF
jD42hzDoHJfPi8+T9M7ASbN07d9u74sV7+7vUL8MDih/QOwDpiehwP0JqNtQfa0qrVIibZYS4GZ0
waoKEJnIE30CM945aHRuwgO1Avx5MHNEnp4Unh7UPkdk/WaXBvwSHdZo0bPEP/yOhnDk7PZpGrMH
gc5fwJyXyVJhmBEKH/ITkuAoUCMGoc/gOVQ46yA68fgndV1UT9Hah+DEjue++7L+pQHoybyvYDUo
jKQhXFhlcMCdck1HbjR8CNPKRY0WkTKK5Hrb1wV1aaZo9EVgOjNDccBtUlL392j6ANitKZlJ167+
ccFhUuAdn0CDcJQ3pOWqkL+fp66lxgNyXsbIwzfw/fspjwGfYN5AyEISgGhjvajNqrUleB1jMfkh
49d/2sBzwkjxFFZ5oK0bQ09TdDQUm4j4ZZyOJLIgq3hPn9zs9AJsW03DX3aEqwS3UOqf7FeEWHJq
tcRr56lhc7h4fAPAEchuC7oz7BbzeL/9sZMGdYTdOPYM4B4OOgLSitaaajhxHf7GSkh56znyIuUq
p1sFprRfUP4+/u9L/jXTUb8oRPCu3OTfOXDogr9AN3aTX/JHp2+YgWSZ/6FLoNP2PmE11J7dMuzp
zM3P6QHw8StbbnzE1K/oLc+A+E0L4dVn8OAkV3u4ysCPwRHx9vMBEeBHiGEOuobNOQr8XJ8xFF2L
3nPnE6iCciTcJcVjJ0qcN2qLcXtwe1QSmEAzyWF9yRno1t9dq7agNb6FOHouDrp56h5yOTUC3L7g
TabH2oEIiYs5Df2aPc8bf7v/W5mYfVjMZsyiB/2YV9AOmljAcs9AYIdAWyOhkZTdOTvT8s3KM1sp
YUc2cBJj/AmuX87q3n6T8xyr/X++2NebRjTciz5oPDzpcwzWXvdb+SBSNV9rX9kG2GUqGL8YipAG
YyUctoI2MKt0E1dl7xPbcg6RdwuFAhlUS/bnsWDCgHR03Ai708bcavECBksy7CAlStWGEkVyU6g1
84uTBJ15Do3luQFFkozjej7TMFvbhX3q8wMdH8aQlqmBFpdr/7CDacnn9mKCK/XnxgZGCsHHoc0b
ih5epp6CBoIC/L2apRV/XicM9woXgcnXuRF+4QV47kI0N4GnWpIhbQL8l5ZoWMsE4I8A7ZayuKYH
36joZ3kIyVBXhUkr7zgDVwLpXGUgivUkVJZGP5h/IXzqNCkfQIkh6EnB3Y4QAClkR+9ykK4DFOUd
y0bUGg8IM82I8yJBkpVqrgYdIf+rnzrcwoDmF4BJAnkK0yLA1ZKi8FrQAwJuvhDK1cxGSazhfk50
kK1wZVUbk5rbNcwxXghF9LDbhUZcu3T9kE7fLQpBgmrioJIJxJ9aJxKLimoDBLRpn7YVm6/9EXuM
87AE6RRqab2BqbqaXaPbrfc0oS3ZrkYpzR+xZseFtKRBHCJPDeA1dVRgPlM9cRBGmUZ3JNZDLjqP
C0yMv45MF1k48MkJ5udC6TIDN/2yEQDbzuDlj0ukL5ada/cl7S/1se2npuC52u+1YWztcF+YpqRx
2akmslkiygAgxYmsRiK3dIiHvRDzqrjhXudpSQ95NTroOTg67if5MxntlwQoKS4JYLedM3wy0tBZ
0xuG7KLQv7U500D8lMQWvJmbhNbQZ+hNfg28fs9Fn0bUVKYr+zCWfp7mvyJglj3nu6DMXS0cGC5+
azcKWk+Qo2Eb5pXIWqgKYDeYogueNvrAdfA5hHxr6xceYZx3Ns73XjX36T4QMDbLRMCbUs7KQI84
tOcuuFx7qviHGqnHnUt2MjcX/nCnt/CF48eDRSP27E11bygZuuW2WaDcwS2/k32Px8wVEiPDnmh1
z5dzZWQXiWeic8WuyRgTi1YUcbtj7wXNUGl257PTibSApMl172gbhqzC+97lIaoaeIK3okeRl5Ek
mXNwZQFuCGqGcDH2rHtQrv7wPn6dJk+Tp3bcx2b4oYUb2e81+18GX0956cxALYUPTgiWdLE6mw7U
VRt2gZOrByNfetBB/w6ZvqN4h6vrbejKtid1sVeBhAqotEuYm+gSCJadfYFWqrvgjlGTXP3B9XdQ
KknUjLjdF1+4474zWbdBMSg5GuyDLpqshd5gU5gPHb37xEPJXJn4XTghPFYXM9q7SpUj/Zv0QWWu
SfwzztfUHBb08Ftb3Qx97Jgc/+8nvQV8IOc5uohnK6lKTGrsklpmCESGqwzFMRDLFC9E6Cbn/xGc
aEazeUP7nqQYy07jf3aaTjiO32BGGMie0l1IQZ5kVZ9VBPIivUiHpRS7Cwxlj/HoGPonikmtxQmV
fnpIMxkFVaxzWWQFJHTNZpO2+FjbEabc0UyaQUYF6nL44mEODjuvT64+J4Q4p5bGLBcWQeVLHVHL
OOxUFf8kc3stXjJASBJnj0W/9q7+ZGvuveAz5U7rLfCp62ov6zBQOF5BaKKZ/XvTJ7Rf/VfY4xaj
7tVuxnclMBv4VUwiZz/8kL6BxU3ACNkHIEzioDRqU8yaluVJaCEbskioV2JCIyASaJlps2pHlZE1
XDzIbhxyNgZGIwW6YAxSO4PH925F6E4C7VMAfuWg46nZcxbkoTRdZumrU5V/qnFQbvWnIICndMLS
5N5Ra+u80Dd+1AuitupVNr2hyxvaKihfjvIVwMCy1UMTHo1n/MYAirk0V7yVOdBhmvA7jC6byHqT
Qvrhyky+6CWob8mjt7h9bFNZozych0Q57Byf11wW8LDwJH4SQNgbgF8lbNoESYeTmsxkB5+W5Xbw
4EemslaLYCKy7OqXiiSxxnPX/lqOj+vR2d2dlubnrOiUxHGiTu+KFGjBEkSsGJx4aVx/jLylSDxq
e0JXND9dMBhjqvRL+QwZnELQyPSHTcILBYC+uS325NTtO36uDQVz9hbJPfLKXAI2UMDc4mB3soz+
M0GPBQJYVDCAeYkl7nblJuhhXTbkpJH0OExP2ngMHF2WYRi52XUdSZn/DdP6wNbCSnVxmeIAO5Lq
iwiGyTw9+RYdNH4BCQWWB2SC9/WRM4rZG29a2ttnq2eVrgBTmJLI9YNKbwcnE5sxSDmiu1GwzRR5
G96XVvLBOvJQwBvFGUek464U2kTAI76xZytx4tUgF6qLLFPrNuqInthBbaFfbyzvqATPoBy9t4PM
N6gth49p67itfXOwQbL1KJR0Izfz7sZGdK4rBQBpOa6qA58dL3t1wfuVJoLyAM4f2GpXIR0BFyYj
9sVunD4UEaFtjOmTxUYwRPenk9uDaSMGpnC3HXrb4HQsXyVRFR409kWw8C8ZSiFLzNPWZLmY0FgQ
Gat7vJ/kYfsxS8xGHWGlpaqZDtd3l5089fTZp4RChOfBDkii+NTnB6Afn1+j/IBpnEqmnvL8PB6R
tsbZjScz9YC92uw6o7M1qXY9LJuOJlhxcfqKxAIZPlx8Y2t0fiINSpTuGTafX8FQdb5KE2TRthiB
3OvzW2h0Hvu9CbEiB40qlJhzA3vgM3DUl7g7q5b0SxVwynP3KHV9Lpkf/0eF5LG9SqZ205VCx9MJ
wv+SsXBsjO8JtvMgqZQmHKsWH6Qc5yvXPf9u3zO79TvfPQ2EMV+pZVRpZLH5qCaptDXoQvQ6MsYG
ezp5hmQ5X0H+wfr+hBtozmfdsewjYdrFgcTKCKmhbDUVVDoqZe3M9X6XavtplbIvzcSXnGTfqJZx
O+BPuozdIMxzBJHNzC2fc0j2tdNZqnw5zfcw7a1I2Toq+QuWjKD3ctJh3vZNncJ+pf6DKfhXe05J
HUfBn/IOiL8zjJ3TqbpwTSL/59rao0Hfsf6cDy2TxkOnIYTD8Ucz7PaIuB5CKi1Ft1auK5MED/lu
e2++mMmzB4EoMd8J5XSulfrZiZ1LjyCSp2OYH9zMBpdeJSQiXJE3PKcjNwArxHJor0ukpuCM2urf
TTIGzPiZXzUIbLAGsflzofUJKkPkOXIl+/6avYYSwhQJ7iN3ZWzpV02F8CrdEGsq9kADabCKIaq0
NW/VJpCKfjxtDSvja8KT3mLStB2hJ/qceYYgKsxeWWKAGC3lQjq4azQIevTiW8uzZd3//LYReKmc
tGhtc/gqjQ1D4weTwIwDw4KuwXjW2zvwd0/X0LBAihUAZPVQ1XxfZsb8Yq5ultnRQWRBozDslOjC
/l41zUgS1FyVC5mVcgoU9oIglhgFLrBNu31P/HHMhZ42IGUKDbqUZBQ9UOulmDzqlW9DN87rIOgm
Tsz9Fheuqwi+IMjimvNV5dLehyw/I7+V7VFWTXGgX+3hai1hsfR/2gfI4Zt30490TBaPUtfoEJRH
UgOgPGLnA/Umfbd0DvV5ZCCy5YSZaVZMrpmF58/+ds0vzJTysn3zEdSLLtYPOohFMMfVSvC8NDHr
cX6h8iPAVkX5sp+HSHI0pb5bbL3YOVt4jYQBKCoJ88Obxg4PWHz5/KkTd2+nj2RVB8mn1j6kpiAf
NT5DyatsY9nuVmgYD6/+GwIDAYyHCiiC4ux9Yk4bQRiN8yhArGrLQNIY9e1tFCOUq03xvOqy5G2o
s9/OGd1xWPirlhwVTf8EDSEq5BmYIbyhPS4xiGTMFqZPXbLx7q8j6I7imHtXH+4bDhtCGHpECKDy
AJU2ukoZAsx9koErohPXJCyyLpkFTxtP1jzGbRyG9AyzOHb4BMEjQxNbElb5RekuRWa6LJG26tBf
Xmn5syI8b7XSqxH/VFk3GCgjoBEMjy2MvzbsgIemkjdevgbhXuq8qr58o27jzAEcbejlJp410X1R
cEeBc0iL+hVoscI7TnKuoTi7NAg9SFpAl3k9Rrny3jza1MXceDrrjKx6Vk5iHLC5z43qp2FC7Ckh
FaQ2xLzF1toBpugNSLl2sXmuxj//BjTbBfZpeg52xERhtqv28F4U1NEDSl/j10pvaYOflbbscypi
4nefrl30e2NgmIFi7VLclYG8KbAm30pVJ+BktbCNegcuEJ3Pm1LFRb4QCfaODXBTvKgeVcWiqew2
wkjrxbYzn7jPB4vZBI1CWdmiEhkh3lvZXg9XV8TK33k49dfAGVIo9IzOu0PxXOP0tgdNuPMmTiCX
eDtd2sXs3dfQrClXJDqn3FibBUp65kqpdclWhdQXqseohXWav2VyA5aPO5An4mCuBAUUunpmOBf7
dEbSJuRO4TZQBSUHTBRAgeo/nRwmKuABoCzG5nkbfA4r6oRjaFQvQblFVU4qQy5lGhUcsrF3CLwW
/oK0qlUmn/DKKPh6m8HXkbAjJq5Yldqq0zsvX17JWtFwlytdZrqjLN0FzE0ZV6l321uiCxoenTcn
vHfjO0FolqTAwsGbGsHz53nb4LckDc5e86iO1NGV+6xw50d/SFjgbE9hq14tp9RP3dUr3nCX/ZuD
i4iVs6ykq+Xdl8q412iz0AJYnZt3YWvdu0tZyvbZg52O0Zk1lO46KQC/ospRXdhkciz1VD5jfXd4
2VGW//kUV7QMUSpBFFC0AFJjENEWXf8Hpdz23kgDaC9mcAPRzLGQdz9RzJyNDuhSRjbX9vtZcBcc
mCJsIcidsx/UqiEQF6ooc00X5WE+7QKH/sw1KrGlE4VgTY54efQwYrdvoJG/aEqt68smFa9R8SZn
xR1LkzG0pSQPTgtgqr1qs5M28xcFjDs+LMsc751t84vdFH4y5HkDDA4Hj0hzaHWFefHCN9Qp8zUJ
o6Ogfp0u8pgo8o/P83XixYzwMlpA3d3Vf3t5/+XND5LkZs1IgVO9eK84f1YcBJ4Zzc7WvicfsfK+
9Ao7WqSwHEsYwSCihSuji8gTSLWSq8oLorvjhoivwgU0MskFjNMw6tJ+Fck55bYQY58ypOvqxsyj
yLgAu+rVPfhs/iLE+/BaEI09E6qWKrt/SluVYb64ok2ApIByQBKTeB2flBfY0zKxZ2p5eg+9BVle
7QPjzVaHFuJgZgBnbFI2DxTkaQh/aZFWKd+707mzlMixSf8F+sXlO5r8bMEDPzNlsi+S7WHBscFo
WNWcHYABGvzbOBI2UmxR8qMt9hIRB0Hkb3c27wotfPcCmGpjLCTub+eyAdOuzyyDujYyL2LcET2b
yAjR+kC0GLKilho7yU/DyaXinaAXVwa1sa8haCm9bjp7lUdcqXr1rLUbB7MnHwQkJycb4hKDmj0Z
s5HrKcE7+NulA2MwQWYvOfubcl2Yf69e5Zz4a4A4NdtTMKczzO9HpLpDstoGm5SrB9KaItGorCEg
Y2/fj+07pAPzdSQyE8RdMGFnfj9/FFAgBs1EqZ+om0wPfK/tlK3kRdtQHt9J+1pLZCoXVI7v4Qhz
83K+nr8fnRj1YsFJzyvsnYD0lNPVGhMMpDpUnFZ+WU8TODRxnEpOE9judxVTGNaW1BnSx6lf8M9W
oj3cHjhm18SPDR/592CAhP2hacAC01GTew4eqQESXTHiqgilcHV3uMxMFD/2t4EMD50YAxUPZqDy
R418sCTS2E5O7x0fb4fylk8aFal0YA6OiWv3eodEmUBjcK6JQAtiFXWvPq8aZj1k8fXNtGFMUQad
+hsI86QG3Ao8zh62rkddBqxnjpgYu7wmuf6cEl0U1ANNZ85sLWk5wt/P4mF1cTo/SM3g30ldkqWE
BubebvsvkVivfVpfjtxCNiPmWaUVSxmF1NI/Gj9/Cvfopptd2TsPO8VdFcM2wTlw0bCOqtu5IN3z
kGN1VwU8FIPZhDTxoOJdxi8oGKulTD3hvuJ2BsPe9ia0vi2ENkAwT+vo+BqtX0wwXtn00YlhpDu9
lCFbQ06qkfYzP+KTlVhBsWtc7FoDAwELPEW6VvrEHUJBD5hW2PDxvbgt7OTxtmKyl0zhId4Gd/el
ESkaBLtfLQZtmZgAnmaqQm0mr+dDYcmWf8Ulv+nxhLocHdznTtVJxsQcV+OaKL01ndBaeT6uLIWY
uF5UnIzhU937aRBfwzJPLA0nXmy1vQLDeRQJB5atIKO5tpoxHemE2iJHjnY627vFiay7UzQRlrW9
eUi8giF3qIMAtZyjkAPVuRetPjWZgK12m2uCGH57Lga7E5LCTTgT1/NCeuIEgtKsS7aDKJNrsAj+
obPVRzxKWPY6nboqXnkm76N9CaVM7F+/z+JU4ZHwEMn49r3uSar9rY2imq+CZ53pdf+YygF9SVO4
/8TnJBWamU16Ukl4HC0Qj/TPvop+xLBd48aQC3G4gnTjsNzBg3UtkdreACZZIlyfP66eWiOylBaU
OREiij4s9mrDBzEiIsQP3N/2bvjnAhxufrH+zS1bqq019sUSpg3kZ+7s6lnmVxK53JHRAjxD7O2q
xDQ0j9RZtauUkgoT433Vg+p9qp2XW8YDY0YoSb9Z67FzR1Ursf34YAb8ki6AqZl83x4ZAC9nHAQj
eW52OM6gel1dAut5l9DpYNP6nyfHtC0Ae0IrAaZjjgKVCZavx2FU+bS6bW/TWdB/uJLRHrV7RlFp
CDd2FpdpH1EPUD2ZfVwhN+FRnAvT6HljjbcvHLezjpvFhVSj9QLtfkVdWy67f34TyEk6e6iQJszo
fRwVEQLa+gWMFK0okeLqtwvY7HT0WUU6A2kJEjB+09/zOAwcdIvuG4OGRfKQWqnht+ShkxzA2WeL
OjaAo1QlQQeugnlTi7qQMFZnZL/o1Ss6OKQNo+L05sDrivcmoC51XEa8WvNbHrT9xOcevPDzbtve
RPqoA8Xs4kWNgesX435h8Y1a6khMqfrvbJVdlX9dPZtmRDijyScDIEq+y1Zo8fNYtamkSnJgLclD
8umqEj6CDhsFzVOje1eDHgGYN3xlPdeuwIYr8FEuCLtgnqGmzOA7n7gmrm5eLveVQRush08awvRC
hTd1fMY5KSORYK5Kl01ulgNRXhwnl+xIN65+PqI9iEayJGTfIQKfQzXaQINFUEey31NiNaX4346F
B3rcZvt50I8keoshZfLIFOWlEPGS8sIxAXBlXh6LpCwrykVJyVznSB9RjZgoF3xrehzUEWa8piV/
cDlcG0hM5CuQbGc6hewDgyw17EoU0ATPXyLxDcEXU9FirxPON3Z/4a9IwskJWyEt09ni6hDUSPaP
LJ82o2ggVqsMgauRv78+ohE4Fsp5nj7pQ+ODe3Onf1QCP5rlTxsV+yRW+qYxdKLczGMvPf4QACvz
7Vzhav/ovc8nXlsGg2DibEiTCdDFs0jqH+Dt7c1PHbmaauD+bg7YYJH/R0tZVwJsHDw7QccpxVAO
cQy2Qm8LA+f3e6qOhZTnUWOzpK4t8RdFneWEQyv7u529aP46YYAwZzwt48uvUaessgA7bHkjIvHf
MDI5v6mlIgtjVtZwwLW0Y84nFudX9CqvMocahX/2iZdoVoeWi9kJVQpsNHxZEV7pDZDUeEOSE0Hf
O3HCG5oeDWL0TqeD5rGCCuB3gzc82kgjlATN417eJB2bdOzjuvE6tqXygeNZ7QsXnqGd+TYzr98w
bLteJv6XbZP6cx7EnqpzCrPWV/fQetkM72Oobw4myAcIg2eQ36OmxUa5KNvPdHsUHwKtG/VraXk2
nDowylKv6a0gYOCztKREr4/C4T+LSWImvwtzHsmOqjU75OOYT3pKFcx+AtUrNZUm0tJht29OhYpD
MGBqJ/kibkWQtWuI+xpBvVvfTVPMbYOKWF7EiSBHRBXMLD/3elmJxtTeaL9WyJnnSIMYL1lJaNyO
iIEMdKSaRHIO23QNPRed6zMH3UMi2FgY9VOO/ofXswCoO0TwXj1HQIPEE9umK3Xx9oFM7EoznDPK
mRAoKohlL3z7YLgATCPiOO0BvBNX57YaYJWUoTdC1pmiu7Wh/SOIL17l5seeNJCq3WCHwC/JIVfZ
4k2Hv7KE6oP6LqvxNCV4dO5WJnog0tIGIV9sARsjrW5BVOhZ9TIpX/Nt+zOATqJaHbDg2Kjj0Fmy
I4Cw0KY+nxhZKyM/OMg8C04I1MzaYLIIJEXiw6NUwk9ZeChfYpR0I36/hrACe/oqRPNLgV2t3nwF
M7EY+hjmVkAlMQcKwB1TKAyYS8JxTcoClC2Ck3kyfZOuEHQMZnp1pBcAPfdJhtEMAGj4eFKhUrhs
RSP8vFOSZNGgE9qUo79lunWpinM81EwVGbhjpjhfVcSzVS5wIgErwvwYCo2ievowvMiUe8XEDCQV
IiuV6SEQDV27N96ZGaRz5zJ52WPT2vG+LsY6afjZRRF7no65Tupm7dSFf/Bp3Is63VqSDldrUArH
lnagKeLSlRRtWOFbEGsG3DDEfROLLq0bj/nljcqgHk+cOoDYoAuc5l12+Ut6YITSz2fBZm5mAItI
GjygvyU85G4jJqrvjcNyLz9/h7hn8GR52W15CCSvkhhJCmiJ2rcz0H+K2InlAXu0Pom0sOE2cfSu
kvtwC3g8xNUungZHUAO1MILddMjLEhmo2MP5oMThZqLTmq5lLOxV2HuLWwyGampTIibwiWQsTOR/
h8kM/J4YNxufyXK2rCSYbt7BObrInxGJ2I2rVXoBOFG2euv3DKrkXA1mXS/b61rFDAM/cRNjDvhD
2v8IXCc7vqJx8SM83S+BF4MmUGB/Iy4OQEHgREfTGT4MIkKhZXf3YCx8Q4RbC6mAAoVARvW+lLhJ
DfXb3rDgxUzWArtcAN02LvSdIV43Tw3898SU1dDtN6u79D85GkClGCEPXgEjvG401KQPSfGEgEUH
czN5lUPT3VJvouux09LH+zWRj/WvBvRg9O0vA0+KV8a3NtucXIuEj+kDqNJUqLP2O8QPq2XnLlgK
4MrJiSaT9ZacZxo6t+TcB7m6+F0a8UFblhj73MhgQNSzD29qYtuDxIpI7jcV4FGew/YIe3F1UEty
A1Xm4Yjf6wo2JGc6lE5oakYFp286wWZKLL4jYFRATE4PmcimRo/AcCaMpIUlmZIu/SvJlUMKpWJy
fnhXJbbadXOqKkyU4DjcFirSEb1kA5MkyOqXrtP+Xjdt0EFypejO0Ef0xPszLoPM4RZKeUsuik/m
nNXl3gyre1c4WUowFDpjT5RO+xs2ce8wwigo8cPCaDOkRrKsZcKtj51V/UqWsTMIoaBCA3CwN9Dv
+uUF/gXLxacnLK8UrlE94NuZ7h70VWVSAcnQ7IWyyKfjoRp8Gy1tyhK5BHMntb9ul2EjUW4atrmX
l5IXGrJGpd9cVhdhMboBIGEwMXmyXBifRsdDXbkaTLt1/KVqF+KdHaP1+wBDIst8sWtboa4wl+Pt
YU2KxJD/81E6gg58fehTWkv+I/ASdPbGcOzzeOHApLZpfUhprPa176ZGxzmpiPf/SDpy731z6snN
dArK4TVWStvwTc79qtU3LdZxbQVixq9JuDjl8SYgHXM1qJBFY6xaUdPjCYeVn9dbcdmtpSN7eKB6
D5d6hmxYqXSURomcHa2LH0kIFLOBxHXFqaXBff30mk3N33fuXXejZue5WbPDbAN9XxaYht4U3twU
y7o6tH2Cl/Ju72qF6YfO0peJCk+InZcvOmIHGWrsKcj2ty2mgfwU6zjFbsCLmOyHUcVw6UH8ilzK
mFZ7pekxZgGnCoAOlF2tYiXm2ceb6cPCczotJYvsJfWJnM5pxm3ghT30Lt764gL9j59B/6cvWAdT
20GOgnd7/EXKEZKPPFMvM2qJfD5a0IKeEPkzpnpBimSjs1LPZ1tLAEWkjiJIDNrcGlKywYJGO03X
isZZsoncrZq6L1i8ziM26+3VYJcFf050bS3unelxkKOyo6cuN5sTa1Ng9h87xY2Pm9Gr4czaFUku
8ukf+EbiYpBLOpySiQb6WuKbQy/bqk4PQKSA7DUjOe/teo/lodCAluTyYS3nYN0DOG6ibswpt4An
pkIi4/ta/LkXCKzZoL+qiUH//vSIvkyMfQCM3uMgX+HQ+YlFgeLhKYoqbphwBPe/2Bu7ErMqrMAe
z5U19Y/JFdMq/cUBEK4hSICq35vZ6VHuWXVqFjiWyl8VNAjzE/df4tmy2C6w0+3iedMKnXo+Dk4T
ehLVbY83ToN1oZ4MgEsNeEAFXxftcxQMza7L4Zw6o5VZ7V6hG6M817gQyYyTGN44ZX2IdEgKYKQp
qgl5jk8s2VZHuKYGqmM1/CrCupjz4JimNvHTWOw6OopVWkxP/x5M0UG0UnMVTY+N5SY+TuhWmLfM
cNR6wM0G2A1P6aOdJxWUp1zoRHVarFGeo80Bouoe0o+5AnYKmwXfuK0I4bQyqXXAZ2/9WMhj19Cw
Gb4qAylqes2rDSgxnanRHvp0lWvvR2RMw4yuZFeYsLS3thbYrSyCKun6nPbwiGXq4C8OT3O6v7Db
Z5c1gTEu4aDOb8UicDTJY2n2G8IT+PB1GFPEAMFnj3NTLMOgZUZoB4iTs3B2ZUhHDfE8MPTc8qgH
YhsoFfS2ZEDCIoqK/hyvXFhYxO7KYBKA5eDUeE8UwnjwFpYeXVir52XKhPxYvGPoZ9Zdm+PDmtx7
0+MJNka3BVWywDYU1br/KGgOc1QsZc0kVJ1s1/wPZb4zIehLgXiT5I04A4VduK6et7LaAI1itc0/
hhlAGX86XKDcn3aBEQ0CDXLKrB6d/7cJub2NjKXEW6yiNJT97/iheviOlVVERt1cw5eoEnUAqhkm
Yympw5YPnIkdeTMU38Mb6vwWMsDav1Cla0Me8gTP+kZo55eIRMExxwoD5dECrkSJCN1I53TcGA5u
2t/xs2On+oUvSyuL/18yZ2PHQVmPLydPHgvh9czJpvB1Dmvrbnsy4G3uZAu2z7/lB+HjBabwvIPS
kq2JDIGVr2zyc8g7dCl+8fId99VbIlpVPugosfgrPXuVjzFfmpJeAGIgooeyvTeZWKmpvROrcgx0
GgSVLNtCNnS6dtWqT9iJja+W2/7gh41xmo2BR/Pqh0JCpcFophh09JVhuKRuK/0y1+CMY/feerBj
2kjxh8dLPvQa3R/TJCt1XzhP6Jqqfbbesp0Y+NDgwLFRBWXkI6RLYxP5tKSxuQqQduBKyrjlUBN1
3s8L/HgYE1LkK+h6fik3nMLZBCs2N1H/fgioBZ8IKKEtml8b7imm/vvP7TR8aj/uUitYBgIOwvU2
UzJIlfT1drLKA7KkZXjvdsicUmJB6bJs8z1ru9ECpJvbsxve01gT7yHTYnK5HuTlArVszDZoBGw1
pwygBuyuZHdwdfFeIi3F0IDsa0+FpK54GMoPUltSw37Z2McWahW9F/ajBbtmC76sRrZEB/HwfeE4
nArFmbokXv8+PdgdGcc3VItEg3FGDZkmA9k52CnQl2KYyKOebWWBFwaXRYcviR2xXTiuf+jV/0oZ
eZNYyoRKRxGu3CW96jrr9IhWPDnzYLJ5zw+zgowqxI3CNxLmYwapuczsuia2FrF3WRM2VoTuGW75
55p+vBeEhPCjs4OkirRCsY/cknlvn1GPyu0PEiclZbJysVZZsEHcf3y3aZNT3qjg3AwPQGjwSGFD
xJabFEeQm0VI7efeGL0FZxJvpN41OA0qdIECwM3WftYhEUTgFVz7CTA/Srd+iq2y86mcoZs9iT1X
/b/boYxMBieDJBTUyETGxhtpsAo+3KVKP19vilv/qx1tfXGBFzgleIUJFAGQUSOHlipmxqJQukIS
ijDfi0QKN2rgTYgNxciUvUhBTOAQmmYRMRQTEJjgGhSFBRBJRnbcCeqmRk2X9fOxk096CveeZQEJ
IAPvMLlUpXuYmZiK2BIKMz0X2LOpXxezFwmkBvkyWM/QaL+hlRoJPZlcJkGqtKkL+bgYsYyZFSmr
9UAPgQJlhxTMLYM8v92/XohEKmNisgLMGQQblnimZXelQ1CObYZ1z0+qJGaNzasoa8QnnliTvn/r
PRMs2Z9IrJDRPkNWdsUvpFyZl/Izmt1TPQWlKPFqdOOdhq2Wil4gXXQEb5UFIt31xPj0XJEKLa1h
m4lpiKrFdD3fEb3R/hAbiFtjETXUoJc8BcDvGqXyONlelyVa4DNV4IhllAowlAJJpqjnZEhQfgK8
YSQEP0Z5Kq2f56QoanfTMITkgPMyTnD+0nr9g7uaWGNnrUOpcyNpBfMD3vNnziMsJVQ3tNQOyYt8
qNN19TC5W48BmfwfXACrh+aB2SAigy2PDHlLMlb92ema3RjSrINaoxUZzv0m77R5I0QnawOreiIO
PjrA2VyhYIMlNSkbNGCIyhDv6fdfraK/Yf5i5jFcZr+bLvOSDTCDYBxhaaZtwCcFTq3+YBEiEDho
sRQ97c3TrfD9ywt+MHO9mP3SUnRh9/mLTCRAGoGDXoDxKHsHNwZ+DyEWrSC1kbsAsyBa7+kaQQGU
USV9sAnqV+D4433F/md3ju4IGpm40quKTanZjILDudMee3uBOpW7uHrWeBsPhfDZRwVmu6Yw1gs1
sPbuSLLYiI0UkYArwiT4C6lYp1T+UuA4+sawf5WES2m52aQ8aMIbDWl2zh3szBTVJ3F/fz85poy6
moDDKR56nsGTwQ1uGZbbk0SXCu5Ju5KUkj2sJotVA3p6pZK7VCBs3Ckvd2PE/COmnBHEYgOyYc3Z
G/0r0bU91FVMEtrKBbLlgxmUU8s4xU2kKdF+Zn36A13P8kNAQjNlM5YrJhTrzPMTSD3ZtdElPyOV
GLE1uHMS0UEo8qDcMDABL3k7cdmgRX4unyLslWDtRXBWBUCcvuREJYwfWQA+fQNIR2CotToy5OmQ
K8+KHELl8gXyvd6tGTrxkmtXwjl2kwwpqQzgD6P5lhJQQR/qrLjxKWTnXeWyei/KAELtvuLB+NZv
WrVBOGZy4+dm6oS0gNHtRkWqJDqXc5chSq8p0jSIgenyJiLJVZpjeeOtvdGjoyeejhfZUCPAgsz9
Oufc5yFjaZ6f2Xi5VHsPMaV4nT4ubezDIWhSc7c2ojDyG4xAsjfi/JFMcvGNfizd/gl/O3S0jrpY
O7Jrt3K6Q3IOHXqRww7LQZO25Y+9jefx9ym3AlZ3OgY18LR3RMsVcGtlrPuniH9IKE2gk2vq98Jp
7Y8Sj0MuuMdM9oYrckVmWCyGkQVNcCibloCE2eai15Gj4pNyjIN1PzlOgmqNkAqr4UVn1RCQDblf
IEO+qgZwKPWXqUzDAiL4y55XsGK5L32w2HNAsSc7ZhoT2nauzknkanp6LGuEnv3f6qLVnI/6MruN
D9rMvyVHdWTggW0zsXMY6/+XgxC7QGNwp0EBAZaXp1Xxyb2Km2WzVhk3gtkw1cq+TmN+c14u6/Uf
xMOM5HN5EQgbtUDhpKb/OCsSU2XGzUxPQeT90C3VXmbCxmz3NZnGTBYOJkp73GKVRwdSbqojWNyY
nrqCqbQDhl6Xh45TTYZB7sxopXmeDwpwFtmaukrn4EYFRhu71VF+owcopwe/31Mxse26vhts2Gpg
F8pP5cHXseOQpbPFbbaussRk5BbKSgQxjUT0RQX4g6wXTiIwP0/u5qhRfhl7ZySnpYNHdW3AHZgq
c9jkWtVYMqecsDA7LVwEzkzSrI7Kgu6K59EykqRTh9Rw7YmJHqUBhbxLOYcF8wUBD6PDoj9DsGqQ
AjlP8xlcrNWAfJU2aEvsDf/hObuN/FdQwUu4SxhXBuoSikU4wsYwASfwesdOxAwNZmr3Wf5wD3rK
5e6H4GzVdhY7TvDqrY1ac5x4fppH01+TRpg3dbnxFihAtNIpTNSRDEX3niwGNNz5yNooq42ClRxx
UyT7DFyiLvgb8dqyPXk/p2K7JSYyPowMfSK20fJparAurrwZYhh/Z8XTqDX7K7ErH2f4VKWTZMLR
mqFMRdryHlm5pq4e8SfRs1k2y3UXWVYXI7QpDSmGtU2LEIKAshdVaiuDZGTx1GJkYLHRvjtuKJK2
j7Tcxh4uzD53lZ9Ow4D1cLBrqIZvN3m3tOvlUvk8gz2vcJD4qv9zh+EObciKfGiQTB1OtdwPjMt+
MNvRK5yWKLwD8HvJ26YAghTuh59+OCCTPHWyrE87pDgT1x7bcBJ58M0HUD01N/RQJr1mWp1vV5nP
6GT46qbDz2gLUtQS8I+mD9eG54Kf/JcD30RAkC5FnMPXv20HKCZ0rUc4Sy0O9U0hggwu28Q10MjT
t2+PjvG0vQVKAYZBuyQ/axwM3Hu3HzZqOj6GXaSmAcWjiOOUzfX8pAGbeqgmFscMdpSUidgHD++q
xsOhEr9PCNViJRhdeRgVU0HEjy0AfAKniru7zLTeLSmM73/Xjwgh9HyH1mkgW7ClA+rkYK5Quqdf
0oev0JV0CaZyce0bA/sDldnk/65LI1ZR6OSNbfdsxoDORuHrfuUpRXHOCI3qlDopmkAEujYnPB+P
22xtWFJ7DFR906fyaRRk4hc3inBEbx4TyOzEDxnM+jXuHfYzPF8LPiVmoXdB9R9hWciqqPLbVSix
49rzYcdwRPcePQRZeGXuA8n0qwqSsYskxa9+inNte7crWBQBuii191V40d9k54XsSxBF6BLae6fF
nRiJ1DBHRIE4pghmsc5yiw+lh+PMDFCGjBFu2x+ebKTaLH4WCWaCRbZW6G+rAuCO4UX47JJflgxW
6Mh//HFzxld8lrYtEQatqgGS4JJ8dVs+CO9Sh71CsuwwMsOvtKg+LHts33cZwoq1jngRxpOqYA5j
OsHijVvE+YJ+13C2kEvl8kMKOzwDUkbjp2cXV/UGgKyiCiJe5wO60TcJqfWzFsmbD2KD4qip0BwV
AMx7PU9NyziQE3DLUKbPhc4Mo38HIlTeW4WbovkJOTmhKgZ+6DqSFq+T1qkCihggc8kDU6KXALof
2FU+hdM7xd5JOWBadHvBV970gMcLW5srzh20kKOvHH8FpMTNqapQvGItQyrR4uYK0gujAm9f4/Zz
rqVZS/lpFAolTyNENmkopzm1hrzucubODm60jnn9TVfvvgUXlu6EmKg+qhlxXdShVDbfPMokJonY
6JANVmg9zH+MTUp8Sdl86w1LiSPG/umQDaDz2XkchuPuR6Ri93yrlJQ/rKijGIl/yOqHTd0o1+Zj
tUiwsrKLQjhMEfyL62hfYr+1vnowfwq5QgSKiIMn+V7aMRKNoxWmPXb3FDBkZW183dna/MZ06Q1r
dIG+t0xo2HXx8l+IXIWJ3Q4HjLPR6nLE2lFUlpc6QYALnoW/OX7yoaWLsshfsmD4pTyw5XIA9G+Z
ItSW7QvuaWmMVyb1u5ogA3zX/fzUVRI/K+t8eZqp2hgE7eTynT8Qg9uMM/UaQt9hRiLbYkA4xlw/
PK7gnsgki3HFl67XbvhzTO4GZuvpri7xpdaW/fx6Vgbz1UvFF6SKng/V2ukgKR3p0+XNAnc5F3dM
Wl8Q1GONExtz0aNuZugHJCYaVtDTTYC9zhM2kghGyiAb1+ULfxzd3b2TXB+GUXMq/Mo1kLuN4wOT
8I/NLph3xPDW0uTXMhohw4TI7qq2npwJ/VOWuc30y6LEEGzLONnO872oR+TgJisTlP7i4ajEzgkW
ZRblPwg8Wqe2q3J/7qW9XlphRDvPtmC7Aw4Jua+SF5gI65PHrUf5kiZ3zpJKN3VupotkLeAIrLKK
W/dzHuQ1Qfb5dZgxdYIrWAsfrvffeZBU82bM06HGAHPP8SqVAlHtFf7dcRdPy+EsM+gIj/SqrrAa
8uQE+bXq8c2aE4EOyHR9TboOOl47C7+yZaNh+ndSsVNXozPK7+E9cweF18YXDU9jAS8NZUdBOXKS
U66IjV3Nz4X0aJk8A5M/KvKa8azoMWroMtIqt1lLCRjn+w1EvxXw4i/1uPX5GFkmT2xPh2yTb9hD
5KvUeEHdRBlOCRB17DeNy2Pa1CqVpatNDdgE6ndHIKcYbiTzPz+HiUT1dWSHAiHIsvAh7plZ399X
6zClw+vQPrTxKZsmh/dkUXOKfCeNpaH7J7H9IyvRrsl1ncTQprlWZrFtVMlPVUcV25NjrHMpX5rU
KHl8BxbfAFXcZODT2Onub0Ei5LgkpLbUxn8byf55bTocW5xIV7O0n/OU+4jFSvLneY4twRxf6ZEL
TAg0fz9UuBjORFXVSzmZ4+kAp09zeh24TrUS8L/LjDZPWYDdHWu0mwTCZtUCwGIeZfEhxl4805R1
rP2PM89WLPPCv4B0hB6SyKAKiU1+sGK7jTyVQYE7upiSWBrSI3RUrEbYUI3s+pmX4N+3Vv9LvTOU
qg68Mx13FXD0niRnTTUu17tvBkISRsw7OmTQEn42/14iv8fH51FQTM+P9AZ1CdiqFCV5ecao91UD
V7uogIgeFyXfsY8Hv4G+C0j2WubcQuXn9gmLyXs3ZXp/AP5844J8gGJoZQNBNLyw5IBsLIiZ8ob9
uMxaymJsSfxp/zdDeQ6Q76l38Lo2Ifud4c3blrYteY5uon0fEEILmieKqfn8nmrFYdlLLeyiPWBW
vgiFRMY4wGOYzQMFn4zXLjy7OSkN6qiD40kBqrcqlOp5+D1CToX/o/jaPne2ojbxWXWVyBDix4LI
BXNGHg3j2OWysduEoDnwBnBH5RiX5CDIz78bRqoKXmmVxZrJh09eTPkcublbxy334dNNbpXELBPR
jiQ3UgBzbyq5C6U2c/xxMFAsrdOvxq4GvV46Wz3Q0qeH2Ignp7T0+0iCWBOZrlo3OvwzA4NxQAQ9
RCVj6SLeliybYIGQMRwa2/52DU/W9ZgTw4c0yqGGAccUJslIYgOYFerqaNs7V+MSTh4LPhqumQ/2
R8Shw3CW6kX0jMwpYz+I+LNjm9ZUhhw+bVxd7XeSYGJmAkp/rio+UpgusAsE//wAYkX9oUrnyA0S
N88LYRuRUpR387WdGKRyQIDHaAipsO9kb84b/T1wnyPf2+MQKQ/xpSVYK24fym2HJm0otECoFpsG
llaoh18z2XiDnI2tMXulvZSYWPL1sEalhVNsdR2rg2sUz855WxjXsMhb2Ir1BZGvM5gFGo3v/EWr
xaK4iOsg/oaNmVbCrHfAdIAts9Wfq/FErv1FP8ueqGaTUxON/r6YjcGSf/ZVR8tXj5aNvEp2NmXV
IGwgwnKMDpBePIwZst/+jKUjLx7Q60bfbLymoc2nNUTNgfC0UapY62bzkJRnZGeOHRx0rwppQ+od
+JjkKcXMzMWRPuanNdp4m63pd1P15eIwF6jBxjpgIG8nlQbxckoIoSCm1pUa6io6ycJt6NZyd8F+
6QcjPiQs0qP3DkClrz4WPFzNCf/HFygH2xXA5RwXejbbA5vauDJtwfeCaTGpqpQQugE+lECqjTeb
jR12S999ZpMxjrxpja6/RNheo2IUotKST4N93YxkHBffalZDSTPU730HT5DuBY1o7uhvEmdrDLoG
fJ5aoqccF9IhU1Qjs22B8KB9V4wBupqxJdHc+jE8fY6Dyf6+KeJoo56vmQSkYtEEXPED4JT++/KE
buOKKeNXG0kfIwlWQkhcox8ZJTe4YMOWq7n75j1Y1JPNyo2z5X5FjEeI4WlO0g2y4OlXXdcfOlKh
00P0PPx0b1zELrYk2WnqqcGsgrL50nsLf11LwBg4tJ56tt3MsJ056xEpmjAKZx4xpSebkb4J+yf3
GbKQHe/nhNXzNqKYTPKyaiO573Tl6gckFv4QnzFeOtCtceLOG3g70VNqFRQKrST2usXs2qePR2nK
+FAcN+3bFBUCM6id0gRggYizpkZxmT3Og3pf/0dypTt4/GK+xvBdn0s2jAPEA33CcyTpNXoe1/Vc
9+nI2Fu7rDSxd67+che2W8lYSrnuHRX7Und/gss7Cj24ZHBN/ihbcgMyU/+py6lzBK2u8ItBAQCo
bowFD++e2tlwhXQXrp0MY9UUHB7gXrRv1f2UMhNTRJL9wTkr8ftDP9Iog7lv0r3Z9Cfz0vDV6BDz
QJ0zAed4xdzLc0t/dwE3Vqjomu2B/vuDU/pHGjJ9VIzJZsj6lPXqYmzdSTZGa6Py0mlX5Q3emJAd
n8Q5jE3p8kYSlDA5i/6F6gPCmJk8eE79Kr9U/dGYuQNPXQ9dF/z6d7eBhHLl6j6otGcs2LwsdIAh
TcwzzEq07+RFqDglYqiOrkxL45gF2JoTpma8cun6MFVe8LbhdvXTrr423fRo8Dkq88PxiuZ+54hJ
lzvX02+1rjCZMRXQUaZOg8EnglYf9gmCHJl5zk5e+Tmo+xx8f1Ol8OV1zfi3jB2T/4khB2HT75p/
9xeZcV7Mx4Qjt0isqO5vR6iMu+n81qeK4ciM92z9SFGK14B43Zq9hxV/YNJXPF8c/oo4M6tBsuOm
iZ0f+AhTjzxKbKqLOcX4EaxSNPVbKsg7YWev3rCI82AlFPyqO1Z5po8OsqAxD0O+VPrTPhTngti7
Zy3opMmPO3VvbGEDQD//tF7xZYTO3RhliR+XNOF+qKWVq08O/alXj4RvGfpRyFPFebuL0He8qY2D
0pPRcdBII70U9eRIxWN1ZhudrqZQjEtySeWlP0b468RtJut6m91j1DqAaTeIg1DeJPu8nAhSLvr6
4kr6uxcYF35qjP8vbT0yMF02pUcPdDhnX+jQG2ixYTh5qltTP02/BxITU08po+482dZ/AxiHjPOD
tE5HodRVh3iu1KuECa32VQbhstmKFDUMKxV/dC+4e/LwyFi2RX8WY6c8yEQgMxzhMcYzX5rFPMTz
JTLIIRew5p8WiImzW6tsAA740RCXvku1DrBlTixQdIg11zTmKHVGHxtXAgkm/gwh/mpJID1NhhAR
HosjfrhUelnh7HsXRyy5+PXGC8kLPjeX7tM/8NVUTWOg+XFOrQpjxDRe0C4fNOfD03kvX2YoBtjO
NXuef1EaL3d12gIX6uGnJQiVXDfLUIaVHPSfu5AbbBmih/Mbb55tO9btNim4huYZmgCd0tpqMEjf
H4zeAI/ONUc87+vgmfAcnIVHdo6OF0ePedrgHKojGG1AzEzc/stu3gYZXYO8AhaR9+hv31b2Qz7e
YkbvIgLvgNycJ97/XByCH0DT1vAK/12paEBLdvykHxLUOJ3TFPzfbpgZq2srCC7Q+9cSOLumSh3w
2qrA7A/NkHJkI112EAZG7dXI912PEL7DX+FaqF+fU6FatQFUvV9S4uxCmaV5CEz45pW3A3ZHdi/K
kBVTT1ypIKbzaSW/4+SCaLskGyV+ktAYX85TCm6fpLy+EjTxlH05pDAYrOC3fRkoThXu1yNyQLsF
VZjzj7LI9SAGmPXlfFP61msV/dbyr8KvCyKP3JBGyob/Pl8MtgqvoXENXjvb0tcrS+OMn9fye/bj
O/M0IhrdRnD6GF/vM5O9k4I7LY0KQ8KCYLUeHCXmsS30j7BGZZQNsffCcbTLfXNzUo8Zr3VAIIyG
VOM8TCpmNOA0S+gevEsE0+VM6OLadDJf6Biz67S5b1AWVx6RNIeDGIX8Ga2voeMX+BAZX3mGJNSE
mKm1hCgArVkjaEO5PAhevB6bCvA7a/YGbYMfh4oW/Vn973CmWJd3pLXsKyS0YXfRTNxFSfhtlKP4
mf8R/ZH/okjzeToGlXW3fAQyHOFC7WG+UUzIYszPD/P5+ZOx3x08r3L6e88XHiOzDIMPtteYU5+q
WP/CYiPQ7i5rmELaq62/Qi1pSNVSzvJxDXdzTc6Q5hJ2rRSsIowJSMj6ny+4vdoPeerJlpjpNPSg
0Idyj9A2ajydxpbItM+hyujsv1jQV5N14BucoEQGUwBeH+UgoHxxvytdRwRX4e2if2kVczxzjYlJ
F7x1VgTUubWPSmFiP0YOulSHXqGSRv6RgS467ga9SiFhOmW49SFeVCArBOjlUO2pYiOI/PVhPdLj
sonqXYQI3sOrcaorYvYH8hVUwceNYaaUNzrsgKS2yKkNImid3nHtzN21H9dRIip8WMQyqHby9vXJ
4+wxATnSPRYOoXDOKd5M57AtACHLu4eFAz+CEoC828b0gXMVe6M5glOJ9O44/SiT0f6t3YydItHx
6ubFgYkuACuzfZ/YSgl0obWMsiviFC0gQ8aZ7oXRRxLuHAz/icS8GNL8AmK82FZ/D5cJ9/pu5hUh
GM5emUhir1+WeVsHdmqGTm9woB0fECVXVy59kmUCefebQt5ePeGG6ARc6XtAD5+8kGC1qLKZwyKs
lYWSnMO7sf6NBQFC7fmjJn9aB53CTXyDhuLYqKkimBwOZRm9MuD0IvhbW0bP+6YpHGnkAWY1nkdT
HdhUlp/UlLiImZKqhpA+RVRwutRqIdhWnysotgZF2nmxosvC0UTZeP5C/voXr6OmSsQzWDwsvP25
VRzZK6XAQW5HeEp/eiik5xojEgiHHVoxLA7oCdIEQvmFiwU0fDV78PTod/20OFINGUKXDCfQbDNQ
YiLz9vJHdAGuClz+vQBRwrW8J9CJjBji0mvDdwjbDOH5NPo1zc4xYVPGqHDY1scIO1Xr+HKsFEjR
N8kJlPHS/wYbidEPTBgqkS8kehNrHnIYNGIQ71cXmdtz7xvR0GDH+7dUB+NqF2Y4XsfeYy2PwE21
BfaWaaXfENjz2crIH/S8g/ZCiWiJW4jnRMXM7IODHaDk1QyhkdWUSDyUvjl+VR6dqSlHNyuVpxuN
PorAyDtdNhp+hjAZVyTNXSxfC9tepIuTTvSEHFJKwxsjVceb1EiUS1v4mQ5qgNvpVcAX0d9lYrL2
0K1bnAKl0loHZiDuLEJsfw7UxpqZvMjhD6l771lqvxa+j0DsL/W0iKgWW3VakRWxy5yFtXJ/WQxj
s0vNGdCeSfGUtx6sR0DCx0fSXeXAzZ5Yw/lRbKXSnTupHFCoyexntLsntTa/zjmQ8qOmfzfGUhZf
PnAp/HpqdgerkhjuCet5aWcJEtNietFkLC7jNhOpPAYXOpvUJEmxG5DCn83e2g0lhcn3pQZuD078
o25YA7veqPt7L9FyF+XRXjV59K/n+SV57oYowg8uSTWdRI76SOGzejKUUxdX6H8H9qpBYGb6u/z5
EQPrFjHLYIuXo5Ew57V1qlW+37w1oURSfQ8dqJTA0ZLWnvqhiajEwg7t4T2iyOCMIXOJfy1ld0h/
6fv4bepnipZPNku6gZn9K5ibXMo/acjaRDDiuSspGoGwVxnHYXUqldaJCws2Cu3Ul3l4qJ4E3ltL
NIRQxXNZLCx8oKw1YkRY57GdH38Cwk5h5Izx9agmAMEdQMKwUJRBQ8OJ3D9kcSGpGCUV2efLTT/l
lId6dM0pzihmZR6uCA0Q1b5SwqIUb6E4X0N13RarM5/sntXMP8kEIWEt359c30pMbgb7UYM2LqrQ
1TiolJlzwSk2OH7K0a1nuCOQ3cV/rHN9qGq+Vn/F7TG+gUAwZ4S7/6zm+2R/9iPR1SKGu4oVRMub
Zu4wSMFu2RqorW93mNEdjmfY9axT8EvjjFZ2TuJ1CvWtdkIfuDQ3Ta7qy6jhY3qedqx85JoCEWj4
UZO+qk+W6L/mO1Pzs/s/bGG5gsQMI0/TdYVolqq9tKoIWPUPY2wI9MmQwdVlCra2BZdNB7Z8pCMZ
Qq+JVD3rrFx0jCetvK338WRpmuiaEJMXOaWUI3ZEUfkVcO9Cbw53B+8MdyhVK90CckRoWGKRXM18
3prikKHPbuyykavWK4nbuvFrXlCF++QxSIqZLFUj5Baytf1wNbUDi/+Wb3tDBDxU7Zzq1x3EWaMn
//zyzRhinRPwbjxlzcsyakI3fwynfvAEP1yL7s2fnEz1rjRcDQJXf/CnRJR7TPB8c83Y+h/0vSrg
e5GLgSJu7LA9dGc0edcHI2bW2/XgdX6H0KYZJzQwcA3KALd32GCzaMyHn6e8Aebs8FevX0pjWMT9
k2TVzrGFV9EYbkHTA4lOITXAxJGHVmQgqwauOrZuMwECp3zuixn2AD9BCnfXDzjpYhKcjdk801ZW
ohQ6e/eA82WTMMh2NgMO6nbDWqygmkdC75vDePxfL0rQ0A5VJmjw83wA4w5HHLhwGZeHrqlzOFTk
1xKOLniMKcUJo2aRDXi9nRVlSdJeVSaLBwB77MFR3+Vy1f2nSw0b4JXPBuqIVcpBguI+dXkzey6A
V2CwbGe5yo128tfQMNJoCnHIyxBCCCm8DXtEy5LDFohkwgOaL681msEsyCowv23G5yN7LsB77dqb
bva+kJRKTT4I9xtLgnF9CJpG+Fd0E4xWP5E8fr25f3IQoVQPBdGDEOA+umG+tf4T0j71j3Sx1dBs
41PmXXREhV+82slB1L2DfGALfm70U64bN0+lP+unf0pfIof/9+rA19yr0CDw09w36ZyrhUfUcVtm
xWmOudmjU92egWoUJoYaGZm1AqChIgCMf/OmVzOXbW3k6eiaNkRZQ0n3KUvS5u/0BPPfAjayNkZf
4DvmSbUff0ueH3cyj8c4ydTQwv2y1YwMnHQrXLP9BVjPSZPEisL5EqbDjjv+niPYpwBw59SN2XLb
B88Hj6UVIi8zlEL+O36J62GKVlXHbggIYlZM7YUWrXq5n0pRjFztsTtd1+HNa4Ccy9yLXk9/Hvgd
tUnKeQgZ6Pc1wkMOb7M5EF+kgSMBlTOUAzf6F63bMiTRlsW/D8XAMqDOCzmFkiKIPbb4zOsUn7kB
nXLcaxERZIQlJKh+Za354zIFN5FJwchzmX5isCSt+C42I2ANC33g3cpa8kN0MpzLcsY4tyJp8ikV
OYgJ/bB8A3jt9Qb3w7RQ+W4rRzDQilEuCRbkqqYpIeMJJcC/ncvwDJNpdPdgYXlETQf7T82tJ/jd
hogZVqGneJ3xlEbVyThgQOWvZD7VqTiVVfy1B7VBbbIoA+nJ5pTpx6ZSz+Xpgi1XDcaXFAiS68Fz
olCE9YmJE88aFuT0VcfP8PaR+Fw6btO+3LJOJfr38I1D6WpiqNpivlQgEF7dfrilUj9lYu6wEP3W
Kms7yGof/cBJGZPxKfNZI1XwmRfpcel1Us9D7ONE1L3df+4kfgsSWzoRLRnO+B4dqFIDy27IX6Us
FktIaeG9B3nX0J8Ed65XymbUl6gVKu7KLh5cR/2/OLKhAK4MCYpq+icn9vzIlSbqTzigmEEq0Qiz
zbKocjJ/SXtTS3A6eY/6K2xFRkHnE/8XHUPpK5ooQ4qLvg+GiZ112t8mEoFrBwm3/DBdvGPp2rPi
V+zwqCNtYqwpWR/2rwZV7mbvqkdMDUiPVGbgbfQ/hLZrfkXCASAFWufKLQwl5RpYWnyEbXzSencD
HY9Vnr3YUfnR/M1Rxetnd3ZMw9Hk8p4yPKa6RXAIhrLHhEQM7j6pe2dLZKQqKu+pIFUdB5ZJcx8F
3Jylir9L/dJiso+O+sVQzfxd2bnRsM3GQ5ruw9AcAbGI5+M5VjfO4svbpm4ciOm46fyGVu1mGItu
fheMOsq/AAs/k/CAmpItElwZmu1jCfR+5WvKxNi+zrfyGFsTL2W/+BRHQvAkcyiUi4VFKQVVdCrW
Hoa4hXys2JEhzcL2XJMEKAYCEh5D5RdTfi8+TdXn+XCgWsFPwqQ+k4x39fxcbG7vbdkD0XVRY3iK
VcfoRrdGjJXYAp6Ly8NZBFB3g9vkCcGv4+FCgcVPv7/X9VpwVv/6LGGi5UBbx+NVmKuQ3zyFO8RK
/NTbXCcKHNbuF8oVF47RbDj/A6xMJvG3p/x5ouRUOO7/OJOzRL5qNUIfcwZ0leRGea95rOiP4aT/
PtZxI+cSEJyPCRPKarwHCyJG6ioGpSLautsPMJOKnAGMu0f1td7SPEGN2pIdHS684i/J86B144WP
H2JN3JUhfgZL0riLt4nt0DQhTChdLhJ2r3x/eHUZVRXahztI1/nqGNFg5CovGVN2Q/cFHtY/Ql7l
hhDa1/GVC3n83lwEisJrUYX3sKc/ey1BD1O1xP+LdPYuhsHre8ATeFmnCKke1LcNWpYfE796fA9g
14+036pbK1DhxBkjJ6v36IR/U5WYkHQvWjm7BimoCk8/vY3V/FA6Gi48uNyRsEOBHoUnZ3GxBo4C
ZrWyWYyeFsWTylr3/Ey1rkX4mfPsQSGC1Gv/QLRXjh5aMg85MtFHCljGCsmEkeld1/o1Wb7pXEG0
Ctmt7dOOn6+K/9yZZXUQkKw0zdL9aVo1qPvoNAmjQThDBty0UoEtYZOoynaFQNetMjU32X4btsoO
p3xYQ1MUbT9yby5sP3AtSV8dkWElNUJiEQTSCQRk+6/V2eAIF6aGacX8ChmMQZfJeerYxeUUzQkm
c0Ag00CWe/Hl4NCQqk2P8bz7aWb/lMuwkS+1CyDtzdqVTU6sSPBrtspABZ1VV4vN5mA+De5cCSO+
hwC58UJ+XnXV5KUOqY6yYjCWBdgjDWnl0yJN36/62RebYoZpGkWBdVDffZA/XnL3vxA3EF/JYQxx
3MmpKYin6yusrsTb+r7rpPTtuQHpEYIf01wkWRDhDS0igP5t8dYJr/59L44iiovdAxYTFxH2E8tn
fuGy72jKtrMQ9XP1th70E+GVtHglXCLRRp/w8PVl1PJ/YTHcxaizziwfFF0OAd/jUIfiPm+7h0aE
yIDEiwl28vSXyTXtCozfh2A9ufXraTjR/DLf8cqLnRKji435VreXjXR/kstJ0rlVxP2uBpXA+FsS
wtH6ppQx18PaU15NA32eddE+02VSzGIisPZmlVrAFXxMFXHP17O0zMCjVKVOC0aa2idGC/AtKYkm
G0pSSXPm5SBIYCNAf14ZlkVB3Y4hYozsMRGIrVBx2GqklvT5eCaLOwmHcgl2YXjSEuk94Wn5UBDb
cuGp+0bjnUyHHzbKjoCqdf3npyXyHFmiJzUWS7OzF6CLhRv8G7sM6mTafbZRetuwXjZVDB8ZVPDg
XtWnZ9ghm9fA/KgaBTyoO8xHEjlwmOH9Chpn8LCyV20V7+0u9rytkUpWRqwPX9gKo2dLGNi6FsHM
JxmQVjl2XnJJSJKBenIIRPUWiXRJbbOWFHM+k5i7aSKoxtqZGVsgIuigw9qtTkLuk8fVPCvgr1ty
p0WfW04zj7XBIrjW56xoXOIU/9IJjpVNTUNIOoal6YomWhN5scccXyWVwMdSBOCQSs2DOQMUbS6P
ZmCgZa4YiqsznukOyQOT+XKwGkIzyiPEJhFwYwkUF4uXyf60QBh8Z4D8OuxUvswOTSl+AkxCCiCA
eF6aLce6phUxIMlnWnU0VTxser8dZAOhCKDehImbQB+/ZJD4l+y9bduVsVIWdKB4dEN7sbh4Qd41
YMvgDSnWPdlIf8waBfXPNd/jSJXc6FT5S75gc9N/lLifgU3wgQ7rfoTZQt5yMr+znssHmVVJ7Zxg
4LcwwSsLY51PX9MJr6jZdrNNClHGCMSoXaEYvbQ3xMX9AChTsNHt0116bnYXTr4fJYfkLWFHoXwY
YY2JN8HGnFRY2WGMd6+t9pLlE/EUo689bKEnJL6i7HuN2P1j1f76D+hlkvCPIRTM0/bVMytaG4fC
zpmAY2tT3jVKRe1gi4GOcHbrsUoT6w5ODKpwqVaaBT85KcaCkb03R/g4yV23LTkJM2FoG5bLgoRX
hwoKL4Y1QSscqHHvCHIeAnMcI2qMXqGTt33ZC2kVOrwlwkRgBRrlb1TjhPPxBop5rLn2zBZN75uy
KqUnTj/ciXoDKq2eClqRhcsb2gUuaitFLHQpzi/ODSLRkHkte9N9PSmXKL+kfedqqX7jMBjQlPhL
n25XumVEda/bzbwO1Tr7ywIuIGmx4jGn6uCNHF4S3FUSY3ySJFCkI3W2aP1yBMc6keAx1iGNSgv5
hnGpAxQJFjB4xb/0APqZBM0wDUAMaTkb49eVIdesXEQEjp8zTJ+O8HiiKS6azT2OLLjNeKGY0wyZ
I39qvI51OwJHyJo2vbYrP5BQWVLdXPIOxrpf5bvZRZFAfdYSZxekGLLELc/ihYoryMoZOd8BjkAo
Uk5cOHJL3lvUIbb+FfYDArfP2IMTPgRcVNcAhPXGrTzi673mnv+tBZgPFi48jH+RXNGc7IDS14Tv
kRF3J6o3Q0150eZA70OjNGSqq0SSMQaagXJBYR2spV9BjwWeoFhrjQllrBRyTJ0i+64vGiTeQYt7
YrFKKYfBcbTVIOEuKEXoIEN3s6lOYjD7HlWCGTQgwsyNmxS9aTXh6rwbJy8Aqqbx6zEv+ORei3kW
254DeNlGylNuvWB/WfMde3VjfcOGD3VePHVwj15GmhZCzTUTz8MU+bi/mKwVBqfnp0iBiu7yEu5f
5jEqC/ZKPfStym534tQtaO+5dNoNNVt/FWQDl1n/nFAGmCQWAf5Mr+8qc4gonGI9l+Li00En725Z
k0d4gNjbbDizg6MyEyIc8aWekP25ehdajDhCxNXD6DwI4ro/6k90I3auOOy6bPGiFjO0zxWJRZu7
4233BE8zw2rEMZKXpDfzA6LBnUb4Wmof/ug3vg8yzG2ySrX4PfjlQzbqzA4ALY/da+RrDCVbov6r
LpNzlgZ9+fSuhqDqI0xBeD7fynB8YzzEaOulrlsOP+BCMzRYYiUcjMUeClc6JGt5FyrSrea1kz+M
y11S6jlixYB0KXGy1YUE6vikjTTUu/s8CQlPBBrT7EskDVaNa+QM2pggi4Zpr9q8HdvjQDqdIwdN
Jg86mSoqiC71EjgxILJRA8SSUEUvjaMWnWvLYlgxtjeJqIL9hCPzpWxpEp1N4WUPGoumbTQkKEa8
sLl2NQ1cZNZNb2Mo8ZVVpMX3n6VUR3LQ4vs9BGQ3Zo0wpyKuRz1n4dHl2u/BNfL+diFFzGiTkG3G
TwvYvnpk5TTssJ5Wnrx6vbcWQhOPdGt4U+SV4LhsSYMCTr6wFiArunqbzXksSp4j22D9HAaNi7Q9
wrFlEwAEQhA2k3sq8JpdEIjxvvSfxIHsgCuP+pDP6YaQ5mVF7n8rkXh5p/mIST8InWHGOr+5tbRy
Y+6put5bt96ok7lRgKrIIUQDUJSwJYOzZmvrMMQVXC0sMpk5fOd11wTkk6N1cGxMX0NJLY7YxVaZ
T4QD0bu0eA7L/mJIt4ztpsTEu/Sh1iaB214M/x4mSpaRGvaYmWB+XmIRbDjD66ozoPZfTZLyjL7k
aQ3XnQx74eAsea7wt7hYcERNhMucZ8mtLWV6F367974724xV2lJNv0vyeOk9HH95prCmIghvfvoE
CcYjVrDKoNNwpkyuOT1TPP+IjhLZeq6tXwt+jd/rowHIhRZs74WNXpg55L+F1tqgTOUpHwSZC6Ud
/YE0OwQf9RSDMxT4UpcsV02AXVPBpsmVGhz1Nb4EzkSfTdpTF3u1EkZtmQysM0QKOCb0T9tNHM3p
nnJ1W8EMYs8oUEgmuWj5UNsSs5qxyoy4V+vk1H9lH2ShSnyisDBq+k6s8jbDIcQcmB1G/3VoZD9w
+IyYpcC1LWqyQhhWaKSDxZXFjOmQ+pjw9B+vWRKAJn+ASz1xWwttEiiInNqnuiFDUkHar05lYfSm
ziZcJxYiTGITC/W6+3ZtqWBPb1wL887V4Ohaz4yiQBFaYvonAkp4EA1+CT4jTtlJkssvII29Qobr
BPqlgdPbmUvslAnCCsr4u3Q496g3dLLCLwJ80CJKrbIyTALKuTvE5dK1MAMJzk4swmeTDswMWSlK
dYKtu3tUPTxuqtYlTlM59c9rIdChlY8KrjQG13C54KNM7ayTcbNqfiJyKwFkSWIZ80WWwYjjJMSz
BDOqqXRcAIJr8AeLMbCmxbO1nV9hZu2lOUaGR0z2TGqQ/bEtA2KZiD9zAtQrcELObvyYgEtMDdyi
25XsXdJlue+P76Tue2GwIol2Xg7EB17a3qGMTWaJrWZiOWBdg10VKWZbJxpfPnI1koizGxMPJfsl
76urR1kdyiB6uqoU3f5U16IRM10nW84jVSf1EjJw6bfEl38mHTMfBhub9Yuv9yfkhw4+NI8lTxGX
SH4FP/H96nEJVR9V3kOgG2EOvuDjHgasa9AM5vfuBTD/+KX16i4yP3oJIadSXQeWWAXUy9VXAaok
k7SE/PiMaYPUCIa3E2lzfABgceT0B+xrBVidHJ+5DKaPTe18UIF5J3wlVxsoDBqpR24Q3nVI6ORD
JUeHX9Uot21xDZAvidHxR+v4RLFkKBTBn//B3RbVzDNXvbqYoNUvfRoLoeFJ0gWmkODzeYDh+zx5
EnSqIQ5HyHMBfvkO21FiKotS2ttLJdcnWo885KRRMBcY6g10xyUP/56y8yOdHpWXVzip6hJO4hJj
uG1RzhxAhsEtPDC7nt16u9TT2fP4TUMsgCifQY04trpgVJyZB3SAnVblt+Uhsz6eIwipeTQFWbFa
6c/hajwUGciKrlKQCQPAaWYvMEtm4lFNQAYfwkb0emCk+UotADQyLwP1AKK+6nOG8asPv2dgpqR+
Pj4PYoNSb56Q1dZkIpWMo7OXLhjwTDTdJoY5pfbALXiPaImFOGKFxRbHjU4+/xvveBfXDn8n/n/x
EcMDA84C7RWPD/Dc97DDccJr8bFWbmEjCUUnzBOVMfr2BfVMcS8L04nXm9NGMZx09nOXuDstt4CP
x6mNvbzI56lcTUxSqoF9yksisQvbdRtIZVZ+dr7tVcYON+/hkFNSayHJ0Dm3SDeHc216amQMr8bG
tQsxzrfZ0WoAHvg6iIctS8cmt1Yq75O0QEffFgTU7cPQneJECStSz5nY9/mBmlw2uGUp4gJVpHq4
SiJutdLusMATlLyjBm3KVrKg42yxgJWMyQaxGmJqK9zx8IOuVXgtDjR21jCU7w9BZrefcHx2yq3Z
0Jx4MgwhmH08JdOEL8xky2ktfGgHU5xEVN9tUgenfn2OJtRkYLk3TMWHBJeGibYDJetjqgvBcOAg
z6NTH4UTTVTroAr4wH1s3hyUH017Y0r75MiWLCLrlL9lB5ClJKmQrPx0/pwOsZp6KJ7dcEJWZGBQ
A6yY+W0Qm3otAEJ37pNZ57DHKZRD5h1N4vH9YlO+a2oXLHYDYRVnz1chGEe31JQzQ3llUck0nYYq
siqYJW1nUI0sBWXedIlNguSoOwUAZgTIYttc8o13atcuH0Cid6vMbu9GSXmRsgjwMEqn3RFdzFxl
a5utjs9cGVDny8qtWVoDmwUkFM/nq6YUEUj/U6/vfna/fbYswJTAfMlrkkfAgvbM7mMizkzC6h49
TPNd/BSdHQFktktIJXPjBU9v+9AyOIBAr+ZYaAB9wr632haAKXc5A0TPlpgKANkPMwoPZ647CrPi
T+dRSP2Uj399rQjjGHqkBZ1r31/wm3TRTFtvD+DA4gAmspRbNCKuFstfV8lzCkZlsx54JUWzgPrr
9SxLvsh6qAd/fL4k28Zzt6X7hYZZsyGwfGXwvpQmivFSB6DqTe+NPenGisKi1Jl2QGL4AgY3wmA9
JWRJRklam//AWtXoxZl++4TG7hWVhMomW7aGcIfIU1ny524pQdB96/7Jhp5vc/hQZYQ63BSaurnb
sxKsdozhY8hA7Cya+U5MdxgJK18BmiBjsFIuXjU5iGp4fZPmCrU//Oi/LN7umSFi4htWfIhtl8oz
8eAbvl6OSbg0qfG0c7Kxu1CqB7KzBU9FDUlCltuUe/KnY9j7zJZKASxES7vFc6xo4zpNiKniu6jj
qe2Ycr7F6E4bH3fFmQKkVx1jCmIwecUpSTXPUK16IdEB/bwRf3++oXnXQqB95wZca5WaZrnHkqjl
g3avdAudb6Vqyjfb2W+IOOyDCcRY/IDzsZgaKV7vLnKM0yUhTT6J33O5XeiqQk5d4dk11G22uvob
/ISTkVkrcztH0pAlQ2n4GFNPw7q2CuWzr/LEGmzwZKbYzHTCDCfWSB3GV8dNlfuSC/ZQVvYKiW2X
jwCNRVKlJd6TBENEHRyCCRpO5atcVau6XbFl+bjHg7M9hBw6drefx+84EaUCznQUS47n9O6vux+u
YPGjylhOXWxHDipyZpLEMNOABGBL7eYYMg3dvdsABCbPeZ09UdBLgihJeyReiAjlYzLwySdk4d/m
jRHf+cYVS0qcGptKmYRsTZyh5cRTJbkkTgRFpOliglVPKIx1I0q4x6KaGMCLjAI0MEJy9wrD5c/M
b0m+mTxcjLPo4o3DxkeBmVMJXmlUFbyUai4sF11JzOvu1ry33pCyt2qEkeuo4vdjjoJVmkPNU0zN
cqsCalP+Yq2PwfxQ+CLrj132uXlP11Gl7sG2n805vh9Rp1Ye6F91JOwCwkHQizEtUM1Ce36kR/W+
AMvCElmB1aZU7epDT2+VpQvgqom40nZMo8CWI99V30h15Y3P+3xCILYZOYGYyBsJJjoTV7Sq0DCy
w20CagejQAq6PYiqitJrPLcSXE+DoMCiSlWzIK4dn+ypaXqPnu5hyaf7ZMwsYmjHEs/rwsN/cUAe
P7QhxhDqdEAa2+gejZEV2H2tMOFbUieVVNEFVxh3pTtL+5P0GGOOsGZE4xyLdW2gcjYOue1brkbq
hGYM4wxHd9H6QPy4VO1ZkSz/yAiUcyfp4QIJjC1GYOsJf6W/D+tG4+WJtuHiH9XeKlwUaUjXizqr
3ebBqTXyUThasP9DZTHJ6vyW/oUEL2/X2Cv9XLTVqs45ZsW4nxmUDgnYDLDHM+/GKHtA0cXZm4l9
TJNSsoLsXaBLncqjklvj/2ElPdNnVt7T9CcsMjjHpZSuMCfM1qOas7gclos5aABr7KO9yNh80YRQ
Z1OZ+ybJMHSklFyEtyjgy11Wk5j8ddL2SAPmC0kbwKWYePrBwdJu8jN1ZBhpxFyqDUMOseu6YAjj
PyIupXWukdPnGkTjdWUsK9JbwB1Uoqi6G7lxIr4wIQhODLK6ooFOrRCB2ZHbrtv67rDchwXmroaB
l6yaajpgQIGhzIPy+daa+n11sjYFGdq4BJC5xSUMKieGZF51Y5SyHpeNdNyNjG4O72Jz/H4Ko1HV
+w6GwjcW/0aR+2P1XtNtg4fFqF3G5HxiFPqZoSC1OGg7ieIq8wqu9iQsf4Xz9QcHbQsg+wEIgsUb
vL/RA5YN5ECc6DyLFAW2Ipc/jQuYQkQ+3+AP0kz3pePgc9V9AFlB+fQ6I4dNdgG7WFE3AN+kXc5Z
1Ary5/pkfLTIVU/8R3iW5sQYRNwJSkBJ4faK7EuFS1lO0XOzuaEI+irqENIy8GYHhLOFzL3hqJhp
40zl9O57GyQA09o7hAG9guvm5mEk8Ybm/CJCAzy/keB0D4YdHoADQGeaBYknoCwmyzxQLEtQ+i08
VJnKhRHibzRYt1OHNzLwRB8oP3JFkO4Xk0pN2WRLlZHK8YOLMbK8lyYCEDZ9JwAgHmAzm9k47gpv
uUyPsuHx1pkXBRpt1xormSecYtIE5BgFx0lTD6jamXXF59Ki0l13Ec2I2sry2VNsV7sv/5INl8Ne
F3iutqUTWxsHF5LoiA6QaSmY2MsFax4C2vEKdcN/fKeO5MUgbzJKMCHUjKGH60jBA0Pq8YTfTmm0
ZkkPAz01PcJoQ2OJaDYslYdbXOC6AsuGdbM+3nHIy6EJo4QUv7mV0U23DlZfqEkBSLbDGwtOz2B5
GvQXM+04WA6xiTktuw5K6ugIWPnz7gmCQXoGJq205Hr9Oir0cgZSwBiAm7jtz9F0ZGqsABV0gyAo
egzAKhoVirYMualvPg4XDDjIENbnJCE7hKPABBxZEXh51DE/IqHEC9hpzh7pgmMrXL5VkgOa3gtI
QOBjzv/tJ6z3EcZo8RqRKqhk8FSunn7f0dcMNXcygdXuYyPUOg/CISBDczlOlav4VL665LCYRLsw
n1NDazOPHbVnbAV3q/qQsDr6Mh8HU7lQvJ5F3gBoBHArOprrKrbSPtoJYmWS7pfa+3FywX1VVM2b
QdeIn7tWUv1QKM6u6Bc7luBk0PT/8vdinrUdThQh8/F7KLr7keCYwryfBzF0irrqsvqIwQcd9aM1
5tWlTy+H3ajcKsYCtYG2RpwjwRgPgg/g2Da7g46qeFkYcrWS8nMDwE1XDwLjS7iGKZ0vXtrBxT0f
VD4L4iL+v8DTCrnaOgbu/+N2mqR2eMoFE6LVIX0XbC2LcXOkcCpxTG/+PjzO4vxg4/tmpGCcpYBd
Nin4d5K6VOVTi4EEPmraB+Do1LJE6lawFcejVdePHIDB7TJXizT/ffE5pWBfp5BCeaJ/8VXFrYJj
/W9BCrVLbjzhUhwRczL3K+FDIF8V3mssJK0QooSh7k90aHPfP6tIIt9DjCwrvOguZsFY8qebB0wA
eKYZDRaq5EopCvsXq5+9JVNypWFeKR4pDtBVyPP8E2nFSWbNtBlBVraaUS1ExCSs3FIHpTkxKyck
o7HRPRH1PPAK2+FdyQPTwV3Tc94m8xMhionQkJzcudJZ7Qi6ljNUSbqmKVzHxt3et7JsN4K9tXV1
1nVnhUbt27VlzQXo1EDUcz5NVo1MJBOKZ2UZfI8e/SXpOfQwpbi0qSURexTXOYOfAPnNtu5gwKHc
Gk1EiCSnsB1omaL3o4Tg584Q0wWuC1VkEV+jCgRvUxX+521SWPPc+99AZTnXViYl+KagX1rwuFLk
gaJ3sVQK61vRW5LiMzUAjcyFanibelX+ROmZ8RPRd7/mNSQVN0HtoCYfKHDsA8iGHR0CUnVNuMUH
+QQf/rt93BVxR2sJj+nZGCDWEUQ212UK80rnkIoHBfCocHev3p68s0B6eGKJqu+ggZwt5sy1hSfz
L1eI9ZE8xALnZwtWcnkXyoL5MsNWM4Eb5bpEycDW0XXyyjvcMP3xT9chwdIDh2ltFdpbE7Rax3HW
FpRGEKQhReSO3YOhWTl2yac9KAX8OI5wLTD87fg+V++7MtANQIcA+217qHaLiZE0hVXBsR4t/J9j
W/E63yN94FnA4ZT2wF8yPI3nTXKfadLds46byLngGcn2uMVQVr30SLHWP/D7dy7j1ZeouUxtkrrw
2C9Pbl9mg5ke+RgOaK1npgPcYzqJBiGucOLvv+LjVjmEWlUZQ3Ml7fO3k6PDUldsWFWL49yHIvv/
QjTok4zvRvTwUvUsTRcqySnnJaF3bAP2bYcVqHzx/+QD/uXag9pSZPy5vdBIFxadGgsiYDg7eRgB
TYTAUuooBLpIaneHO5CqjtoJAWkzc5kwAT5YV57YkncYgb6EXMfOtRb79ewxHFHL1muqX7PG1SVX
0bG0YPzb+C8dHWsXO50M6Sfxo1IDiL1XpY6FuWPWCWssEQz1+mPstOF3xaiOAYU28vyjpclri8Or
w5ipRR2kkq5psJ9KLEppCIxfkONOJif10emJetlKHD66RfjjgJhtygOI+EJM9MEEEzxmAHCDmwro
zxjeAfzUGlvvrVlcHQgb9oeQGj+1K8HC4wk/a4wsX446XZe3PJgemqCHGzfdAq77Vj8bpx01SjvE
Ze7gecuxx4TqDcVKbNGCjdlbtAsgq8JscJ3439MNlqy2p8w+fc3H4vddEJnTt0aIpV29bN8nv4C+
8VA61d+9yNRzFGzaDFUVLbHLgE2l6roD+BmYjj+tONd/fyG1Plp04VUkVvNueAPtcPhVQmOUtz1a
8rUUk5YXK08FC6kmP4b2VlFyv1dhbHZO0FplZtcwhgTJljtW7wz1H/janFbSRiqnR/nrgbcBRIIp
Zte7eNvUepSUCaKQLEfn5PtLF+lUgLoFSyINZ8O8lxnBKTjGMdrSOCWbrSx3ditU7yuQ4Tphj8tg
X3miRfC6y5z0N+0lGRTZAuG5AixAoiY/ic2Tt52zmnBBbr6tJ7CEFTWbY6a+MN/6RL3dDEq11KEV
WUWUNqkwTMWV+JWfo4u/xNV/OPfcSIpIqCLrC+Kfjk8+c/hTvm5GagIXG32y6qKF/wAue1HoORYD
5hoN/Shkf12hzCquemVz9/jO8FxhhXKKNz7IT3HMTSVXT7D7KE4Bfu46W9c1cTb3DujtUw+QzHSJ
oNfyr8WJTk3bejSrkGFjUWCLHwkR2h9MleJIhxEtO/Mc93rkQuilDafAjurRUKK4cZXsa2QjBRPG
7ylngGMRxJpjZDwIQQ7OncQwneBnyDyj3byfs6rZShmwy/FSLGzAUFsSetPlF0kkcr62RLgFlY65
thzFWc8vhnoF573ZkB2XFFkv9PZoaoDMHiayFt298Fgl6QhiH43WKgbEiRpEfdY4tSnKpGzQG7gu
PRwzAndruDaBG3Lm9I6wpS4+2fZVEjmK1Z6cRkS1iMvzl3Erv6Px27JuIFHlq7ulKuwN+QNIyJAk
pWJ9yFMV8xo7G+OtpZTkCl51D0XMeMpffsbnIwlRCVuAGuDMHeM9RlS2+aAeib7wUGtNnaiSENow
CTG8dHn7ShnRR09dgtBVCV+C+lyfTfGGbQlX7vKH+Y6xmQ4gXs0XDlzswKFhrGUSTx7AorwnoGP1
vSI5E18EBny1khXkWUHJjfdBgwXsRdRCib2yXOCt6ToWlEY696H/hEBQBu8BQ+CuA4mSWYkLRLY6
M4CLAHiMnjFpoG27zyZ0HVGzzN7i258DK/dNOTn/PX7F+MSw5wjqzY6E64Uk2hA+EDMwMHJkoheR
tpSgS6+U+1aIEjXSW7gvPTVKJWq0eae7NYa+6a4fVpivI0ditqqWrdxa7PJLC4vjZqA/omSwOh04
gZG5L/Didiyvg6pdYTtPCzQipZv6ekhJTqPczjyDlW6Of8gRcG7Su4iA796otl6UhxWfOCWsshAT
EKaIX0Hdg0OS23yrl0t3m5s2INfcld8GGCXHwiXvBYpIb6+RXvq5i+eoLUV6HAPkLMfJeKDdChLZ
XJNuWihbzNAmE4UNBpW9guQc2EFJosmvB4X+S+C1VKdi3BXxBkRaX0Epd6a5E7qJCZ9N+cDTVDBD
3vISkXrrPjvriUdc8c/eAwj6LlTk9XM3HZRTNuQtSWUQXyXltqcdGK/oeVUKSZYY66wtbjDsHhpw
Z3XoBpAwOJmTehKh8Shy0boK1BgW0kSJlRWoHMWPdG91Oo/ZZ+9B+Q7Eh/Jrsty/ksKbj5ck50A7
bilxY5XqxO5MUEvJ4HO8N4Ek9fyIO9a6jMM0xDiwWC9huHVuG2G4zQsVSiXYSXKWO+jiA30kbsf3
AfVdg/THDDBKDPgowQWKWHu4+wPAGUm5luvEqC2FMSGvkBeq+XV2KWJHIJ7Yd6IGZ7nnHzqXGS6M
yzvC6n96YbbDeHuUomg6EMOkiAmp//vo/YpEOSA/EWOvmCzGO828nv2740nQScbHruC7W0DUI7Qx
CLRpHvf7wCTXAKRbXZ6tXqA72RaFjTGmR55GRAWWBB3GDZJ7vme9oJwep7joP8CZYMMdEmuShLsB
p8+UgwjJlF+3SpTcMG5YDDwP4gDT46YOYNrlWoYAqpE4nZ8cCbsdNgkB43BIaD8Tp4nRx2SjulvA
U/AHKxSjqykeQAQAbQtmJ9JBIDaGp6iY0Eh/I73VvBsqn4w4qxzCQINaYW2Vdo8waL7oIqHkIkPG
nSBOfz/8MGvZGH0xHtJj+Bqq4/sLZUBzcEWiGBaYS7WfQFu9tuzUcteYe2Oi6/zfBSm7Dxza8eY8
QLo4iYc5tp/54jyDBC25dcvEgY4Zu+OAbble3LCCTmD0kKXD5+Q2VzJG1kAZroJotC8Q7TaB+/5Q
3kTzt/T4UwKSPTYuVFtCQUARKxXGmca9BWQKmVVakqjpK2PCu32w/i80BQ37DBYCRJKtifKNwNxD
eMqU/9sRFO2Qce/uL74VfMPQESK9LgbcOJ0uP9SrMfE+9AXURTUte96sS9L3JHaB3WkWmXg9ZkKm
Ptt5GicYqsXlbUNkmPXa8Xq3lp80WroNGT8dQ1TW0N6R3v2T6JO++FuZwF+bDi0GIMPDJMtGoMXH
13Df/T6zOHxh9FaHp/j7llYlAlDfpEJx9/bMBPzo2462KdhzkCWnB7FX/NxRXXtDv377MfRFbcs5
MK7jUPx2Y2HW+9rI5cRgaORE/RJ0u57oPtRvY7XW3mJx4MLOYElKb1Vbgnr6z0RTjVpA1+6JnpVt
vu7brr+1w+PqPvSF0DYWShdaI+5JGseGHehY8sJ437zGyz0uw48w6nat+e/vyIalkQDlZT+EECzD
D1hsdgBbK7tuAG16qN7dUACaN6mOSY0Q76XUUCjm7hBE32hw4P6Vskb5oYFLkMb9e0eWrNj1nJcS
xk0lXZPq7qJL9NYua742SZGs1HjditWALb0ozkZF6e+RR58L3vlaSpPHXbdzJ+0aLCaHfqsvE5D+
MuXmIaoU5/X46HdRtdQnOobCsx+sEsishn5tudSGYye04MeF/2m/PoNlEC8dxv/ZwSCP1qfEIX3r
FYAo+cWQEYMLWrQxDleIzLVzd9vEdwZduH0olLaJQAPj0Fw0k/yTyLN/f3+BQiiPU9iwa4GbQpbe
ynCTbKuUtZetZ5PzyD5SwcSN3rKiqAZtQpN9K8WOMvBa7PjPMbJC3lCrPIC0nWllTiD1eitFOc1O
iV9z9vmYotN/eqe5edSPY04517BjLEHa1011w0Jw0zGHqfm/A3qnSxPwoT7MdwvG+kCpoJ97R3M6
wlLki9N/rjFvUbVc0kTbKoDdyUJB2JnmsB/AYymq3W9jWXHPyVSeEEU9pLoO+HFHLoZarskdVQQ8
8aaqi9ZvPhjS5HodOzH5FXbFDjJMstTOiUQx+fj9w8xCvIeuytVLxW4u7X0UkfeJwnkYB7q/1Nwy
gfF2hUEXU1Hse2md/38RWMYGWwgIZWEczu0btJET/ItKJCoQ45cB/ALUZcP0HRbBu2sgMxDILPvO
ig7Uyxihkg12+EJSq3u1cg0aYrkjKG+71j051LWnI5NATP1YEFK7b4Nj4vogpbTP16VtHqfWjRKN
yYm3JvyYTTtvPbfwgu2pWUgS1KVI2GU44MhnQrT5nIL890k4Qw1NhaFzXSqrYyfkH0gz4qyHYmq8
bh7sfgQEdgRTQ08bnn01bNKL9YSqoZoUBq9IAgHNtnYXB9mvlzFq5RLYKHE0gmkFhCOLVZjVv7rY
v97k5lQEPbM4Yj+6zXk9UeRa+HLZrYmFOQMfomKWnCJjyCnOVozdrvrdL2rAnJShEMfmllv+K6YG
TnwZG+OALILK1uEJBV0DtVt3kGyafj0wrs4pH4OimzeagM2xlT9lj3xNMd7tQ1o0iZur+l84cjPu
yJ2LcbSr1SYzqe/Se1nqD5BbGDnwdamb374nbSf/jOXpnmW0s0iNcACBVulwFa0ibCT0mjZQ8oNk
tdqd6b2hTWh1xqTfQJN0R6ylRge3Ul4hHj7tBcGyJV/OD8Gsm9pZAXipOzmH1XiDiwt2O6x+P17T
56eDH13imZxdiukqHa44WKgWDF6ieaDd3JDJA95sDdt1d+rEuIx6xvjIfpMndL9dqshELGuF9Xbq
cP0jFe0ilwK6tUT9F1My8TvyCxicxhzbzq2rcQ1bqkTftiunXT3FlNLDVMXTPlqivS60HiVW4uj7
Aerb4D6RGfUZt+7VkONoJ0iuQuDCKQCFK3ijweC1tMzwUbBf7CE10ICjDRLNdSxZQ8RnU396uqYv
UToNtn/dKa3PXPTLy4SJV3IQIE7yziYCzg2kuHzfnxR7IBjTuyt4V5g7zIZKzSmkRtJfBvYYDaTe
+inNPjZiUQjxxhg+RcOK+XgyXPRglrE73WWSqdtAuE1YRa24cgJtBsvFfpfAdroNxovnpM4ogkpX
qdKVEM73mTmC+nn6QZBmBOKlrAzNxSpsFFeQgnqyYlYSkRR2ZnocLNQeuTD5jCwDXFGScbu95iO3
77Gme9M5rK2SErokYg9lwCnFrqwD/gehi5WNcXJXSMlXwC99NgscwGIn1dwKZ/0PfxXo77aDLUrE
sjZKzF1twANJd+YV+5N5wXKjfwrIOvZw7lnSPV3EURMKpMNa94s+/lD0hAxVkcwnyhQ8MQhrE/tI
JOOj2FD4skHDiCn+GOS2TvC9UdNURXFUvWiMBDObe/CJzhnBA/m2vl+kRLFQg6aRgQL95lDhR0eV
epd3Hq1HiH5On/nzMgQVmihdoW2XNzWiu3jfpfKZS6/oKYsAbj1T8Ly/EBXRAFReFykWQjeUOpC0
PMlZcfBJYS9IaCzy22LcaBDMdw1vP79bdpwss7qO3VYEKe8seJOZ6XddRtyd35hQ8rVF9FlOS+nE
aA8D/y5kbJBtOObox0CzsyZQlGz060cYkmHRX4kpsvTRudzR8IPVw4bg0thA6AmxKs49FQ9NXWOP
W9Z0I3kRlXMMBzJ+MXPbr/WJ1fqmXcx07EUKjB4YYzhXOKxevmd3gunm6EgPcMBwjLzxgRhIMran
LGjF5+lC9hZ5MaI3HpxGz7/ycHG0SwStEyqICO92d75qZQ0O8x6TBsLFVdV61Kx2bZTmnLXplEg8
s/EmljnDofjlfjt90RkiThL0jDkez4noPS8TX69x/K2l9lzc3Q+fyjGaQLcE9KRkhc5vlYfKGdxP
KdSUO3y4X7U16igjVXjZjJ60RCpcT54SdKVj8A/5rHa+OmcTp2jb1AWy3Rf1k+2cxVfnlkj5/Apa
IzKdfNnGBvhuxytpKSvcmaOhXD5WBW708XqGBSw2qdVRsAT4AQa/XstFEk1gr8v7PRvxtQJ28DvU
xS7IothnQiLhoIHWhMYYJ2wbeGiCJEu+Eb7PKjRM5SHeHURbqj5zWZfgNYnjKg8SSa33+rh1HjSh
eQPYIhj8HQ0MAHT/fXTv5L+EifiubYvwtlHJh/2ml0sNuJJvZsGIxR98hkpeTsPqthxwIbGKa03U
2F5D0iAcKMGCOe8ZfFG0HOL5s6YiV0/BjkwKqQnotzmQa6TLrxLXDuFPNHE9h4WBtrzwFi9QnFYD
16WEW698gBHqzxKItl010vBQWEcGuA0EKY9c13tpSBk6gVtDBntybfDauO5f9fxl8G9y4A7UnPVE
QYkgM1cVPH/v8TmVarUr1E1vVcTjH2P7O8bF8/w5SGT5V798IiXAYk+nXsTV4aI0cvXqDfA4ECuY
yfPDvKf3+yY8qfwd59qY0R6r/2C4QfDmeJNKcfDxdfSNCIjF4NYT0xJX1B3QIRtsv3bV2fyTLbGs
dv0icOyMB7o/5b5HIuZbFkF9obM7hv39hmLr/6k4MT+FTnGv5h3XtMG+2I+GkdHc9LZRX9+UX3aN
872viWPVT2GxJt6D06biwM333MNmld8piWDJOCgPxHFm67X0LVR+5yYn+pD/zgnPuRE/iRTIu83W
XB9WMdnY3eC9IP+owAsogOTYeM4tqFwFtsRmtM03GMLbC7esN1brgoj5zao1b/zD7s2CNonkFcEG
8Z6USjokuOzsix8gjH7dqnaNmwXniNj/1/wOUsfWqVlEykmX5LKe0aQEvol7z0IFicbeCBoGbus/
oeA7p82PpssIqwa6YpgBkHInY+VLeGqTt5c3ms59rjhlQm9OKct+LoI1prCXJ+IUWGANZKpQSXZa
eWMQ1/Lc43tQLKyvdzdJkX+eTo7PQRMOZNFKDPEEaKjPOE3xlvxoRzLP3wYtLA5PMvW0BB5SagVq
l9EFO6MDsSQLZMHf5Yh1Fg2C3CLJ+APbR0nzfZYgfYtcgXiIavK/Go60O5DeKuP5qsD+na2mGZLH
tkjiY9BDRfKkI5poPMv4Bd6hJUaf8mnu0zOaw0r/9K3qdhBOFsyeRNq0ruH7a+BVAg1Z3kDYhKX/
+ygDF+THRHAaJSCBuMhC0LfQTk0DfFWqum0KI+eWGRF0sL7FLRhjHI0+xjgH9NsGjW/Ccz/E0atT
HOxpEeiZuMiCW+SaKfjztpCvXnJb1tXi36WOhiGd75is5RDefE+QSUD3hMhcbh0xoFZbJZQYnKQN
SrFJ3FYx6F/LtdXPJdFdXvbJfqaXGkd1hxsLSAiOCQUIhfXWo6dDmM6njljf16hOwxTo4cGYQLYn
dUb7bICj/C0mD5jpZXXRMTZXjT3kZWQTXhR+c5Io30x0dJ6AfmvZeWcKWC6ySfcjGF8O/kzZDrHB
gSFu0xxNZ1ONPBHl7v7qIlKRdHKZi6LB/EY6PVVhgSAK7lKeOSIYkcoSj9GvejfhPupXV0rRzpjX
LbF6dVpS0cueX1iHCMyTkLoyMsmJsAfaUcgv7Lu7RDIKCammPseADo16lwpG2NyAUaO2rgEFUor9
1Vwjmg3EeG5AVHSD8Uh9+AkEjAJxdIRdU1DoS4wFAsYhlor067yNU1bfXz2QdzXBsYr1pTDDYVg1
9j206OICOT2EkHYtpIkpu45D1pqAzK+b4vaGERTFCxy7PsN9xbvoSYobUa8WU1loqKX2hsAEYkK7
rGS1mHMJxhAYRmc8gHEDw35jfWnOHdyHPPULo70Kbyjar27G1RsJVn3dOVPAEpybn7iSlohnYgAZ
8DezOoeIq/s3ynB6kCfZwW67ZmqW3b4nVg+qLswOxjHDbf6iLu12dP/vco3t/VrLq++0DMDUnJz3
0nfIk3lH+NiK8OHK/K7FfEXgb9KB3cH0H5bvbaXNGmUihK1aTiPLI9Ng6nuCwQbECtlw2jTJWqN5
+7qu7fdINinao4Oqcr9Nfdl/ki2GmHMB+gOR5q1UtCFVY2gHfABCZ/ERg+Dv1Re94R6zFl0kXQBv
FhvSMAvOtaQDXhedWX3YUU/ZJdMCeZOw/c68IZN94s5YUhMyaoxd569NUE0R2Q8IFo54dfZlKtMt
d41TqE+H1cTXZnFYjobd3vc7ExSkvpU/4EzZZcPkOMYqU4X7bCmnnV4I57GFbADU6swzsff1yZ8Z
40z3ho77Iq3/vOznJ80hBJI+hjgVrOeq7HG/twrXl4InUkjrCl06Jn9s4o2GWoppS1AdN4WKk9Hs
YbZgX/knNgA/VnWUo5k7jKkgd1z/UEhjPjn8YbnE+EPIilJmbzdLfBX3DmC0Z6fSr7JpE8uPOU3j
Ri8DXwq/DT25gSILnejZBj8MGgYEmMNXsbodPE1J8KL0Y6XJDVdCHSCNyPkQ7PkiXIDjhs1sR0IL
q6CAEkERU9qFIBpjGj1q2/AkE+nNw/F4BUHngAhv3YqQ6qt6ZSxIbhkSyOPSxOvjmuU7LYqklUMa
3tdT2WrQCKOOaFM2aqvsLrqwdh0kboxWp8TIsVseDs8BL1HzqxIwhYR380LVXWpOwJEDe4gHgWV8
HT3zzLPIKyav3/58D7Xef1+yeQknYffjkE1xcRJza++SRoIqJWAZakh2P2gL+MNQgig0ZjKgfZ+I
SYFTmuPMpjVx78OppSUEU2RHvE35swJh7MR9bXVU4NILbyyTM43Nzmy1mi1YETLTNTFkTBJt6ypw
wjSi6D7KeUTSkiysN4Qhjv34Ll4/j4WqDk26wvsNKkwnSzLXixFgeTrVZtatXNB8tkYTGJYmZrat
7/d5l/3+Kn+g1nqPoicEIItrc+qMdiR3zGudXdsdCKmLFZVl/h+Cm3MeMicRtT9zdOePax9QbMjW
Od8TC8E5XDGSBFCSvBnOT3JfdRJQPYojrc5o9rM44btHS8MNTS99aRiS2rUz6TJac0v/082eUzQG
VIBmjkZR3xCxU46Ybtcuf85ydvqwm9lWtrZSNGgOssO7sia/OJ8Qg3BjIHDTX8dkRYGJ6/Lc5Sjb
3dB0MUm8vTcbD7Sf3f++eYiRj2+bcaegdeZsq8lDPgFC6UDEQsr2mLY08S77/iaXddRcF08bKJSk
2eMgrHOIuQllgw3s/HUyh4QbvIXzS5KnYJ/sPGNA4ykm/47P9UAYwtT+BrfJBweyES/EJRGcZyIH
rXf0sFD55Z7Tv0c4Z/IfiP8dM1wKY4P7Aigjox8b7gMVAp6iWcDSxJ0oNKf0UqLxqrn2KELPxtF9
ajMjELl59WkeB2xb/tjTRwF7tH2So/0dybnuyVaaFwLc3ENqrTz8y8EJtbiE1wO1joNEi0EbEK7t
R89v9fXiKatf42DKFC9OZz7jtcDMaJabpSdMpPhifVeqEI0RjhjwWXF7qMPnKHR0RpUzjPf1XpqA
QUyVHmGBEZZ0cLQ0Tbr3I1HcLXorARePLXcdDEaIMo4Bwi0rZrGAkcbr901rYREbv8Lf0yUzTmgt
i7S1kru8vuxL+OipcagjuiVwcK1vvh94MDM5fPdtn6wNzHzQZgvDNNW2fQq5EzRV5vkwoD00IHsu
RbX760qzWIS5Po0AQADlsUFHOQi5Hdnn5K815eESlnRPmyhHOgFpD83pesBItPBOFZS/nUPkZVtr
Mkxd5c8PKznhNaCUZFPcJe5gY/VfN6h5a9ULvUS7JqTigwQcN6wAnLfpFlT0dpUdX6hmnNp9C87Y
gjIl8/ZHowdIjHX3bXDGATLLD8Tlg2G/FYJHwMGsTAgXSSnb6umNaYxfBy+DJi2IdtsAcV0ZD+Qy
wkBmEUjxu2ogySKv/ztCV3W4WjqeOuaEgI6ArKJR1KOyVFtJxLy5RsTpVXmwpBuS6g8eyQUvK51Z
epZF68W42x5RUVOhceWMHH/cSlAXsaVylEahkEiy7vnpZR93f8mKdSn4YKv974NW/3Ar+UOUc9Ra
+GVAxuoZeAx3wcl8h6bA4B/V8V34NtOEslAZk1ShhRVVQCNdm9qOpcUI6cJ/DIcGSsIWjBu6DEZ8
k2X6ykuIbcnIeroBebFJ6rZPzOeYZFaZXYBF2xvMoXrD2OJw3UM1Xzp5zuPNdcqJu9nNN8GT5Cvn
ue4HhzY7+dpddnKL8ikcHvKEnO+fskJrl2xjIWtU/u1B1CPnQsXiv4aMFa3vH3cUN/LGhs1pDfZJ
wQn1XxhvoJczK2GaxMKGAWGykaG1hrWZT+Cpo1u2VlM7QKR6e7zTu5u1prMLqymcfEEVqbh6FX8H
n9w0UC94liDWnR/uUoizktemcr8jEukJ+pG1NI9AbZNbPin9EmWDG5rz4LaFqdmZxDdA1SacC3TL
3XQJEF4IhXtowONK7L9NlD23OHJkjZTB/LxaQZbxsOTmZQTTL3iIT3YMJsybHwBofKclVz1NfbiZ
ySWDpDlZYAdhS1o6DtxQIMo3LnQdyp7Ab8eJ0aRjQO0usOf+5Nqc413Jth4k7f78GSjwh/A2pMmV
gy6WaPbHgVGhub0WL0u+lD+5smTkS1KU0dPl9pM8IsrEddEBX7iPFUSNSebBp5CGGA9ihlr34fYE
XcAbTYAcUzRaEYIAwE21GhGj3Jk3ZQtWpo43Ep7SMFSof4uBEJF9Eu+bG68uA7RxcH821U9RxaES
yRWa6TMpy+Q0ZnTswIukCtrDJP27O96b/Kknj8fRZWSQQJNfNKr18Vw1hDF1Tp1c+MySU7p0ZBga
8+LhG9aq4ty3t19YRirxwLl1KkSCk9RUFb2jhMuruW72L92xt/dece/s/NekfJbeBR0mQMek8ixL
Ew+dt+tYB2Rv9UP5jf+7lcSssFdFcir0LVX6R06ROGRmUr0CcZ+IcIJWFtIV5HH/ygzANZdd0rMZ
MLhHhegLH5YMrEHDe3fxHNZSGOCQf91z41+TK7r4Ygi4pQi4nsIki/C7rYRtCRdQrB4QNaq+aS2t
Zb6qy8XXovC3pmXik16SZOgz5/t49j6olBdlHdi2Kkz0D8KrcQKFuzauIxQK0qCdW17r1GKj8xQJ
AXqnffE5DTkm+sbN0y0ByvCK2Cs7YM7rQIdGDh1BofLnl0oLydptLq4A1q7UHcjZo6bPVIPY6iS5
rJkDHrGFBUIdYGh2eqTrmyczqaLdS4Qwzcan6b4uM36GU/sBwJgvE5jHd8+r22SNd7KpV+FybUel
8amAnOVgpV714RA5XXaQu+y5UhTi6RITUpd0qzoXCPes12bu4gARyoaWBgzBsX7I+X1aTQt0E2oO
SW8YOuYOAIq30+hpsU+QgVoVtkKq/5v+R3FbOOHC4nPuLDVYu92SrO16goZD9ymjI6wNLuhrTL0C
OEVIMWWSJr1v7QazxVKEHvbe4wRFp9wAzRLCiQrooJTzYw8C1mPaZzs5lMFbGPQmbmCZetn80VPk
DkNnqD6pPbUO7KvodB9h0OF1Sdx6yCrxO3Rnkuxdlc+iKiUgmDWm+7aC0Uv0bu5fpjToBI89xxnx
VgMoVnMX4YKTmWXN6XSusLtbw7oFX/8VoBZ2PZ/ptr6MweWwmx6HG9XvFkFtk7jj7w2T9scr1A3+
9twihFfTlBR8R5VtFiMKV/mQFfIZl6TCR2e2DK95mRZlgJ5AYtdE9dc4EUdLcH5ZPnCLg9O4rxeZ
ZBFS9vN9tdBO1qCrhnba7buWEve8Y9f/JkOPhvUSZVo2xmvoTPkcDLTdl7eQTihm751tAo0JRmqn
AZn4s/XEfJxKtVrRoAZh6tjMnV4FCHITp9VUpabqbQZZSxjts5twzHE4zl0sLP5I2kS1uRFa9K96
tJwlB7BRCkkcXDyHQKmNZfH5JEJTnhhTD7hCuujDWM18rtvO4o/5Osx08fDUu9/COn8053n+5zGO
2fwHX7sI7xBq3qvFDfF9yKiRzCXcMKJkQCsFcyOnTWIM4AbqScZoRFx0CEVqQa/KE+JhkoiqereD
CSoI6+RXsvqJgGuSRmQUKRaFN13RpuhzfdFnXpOTFyMYepZD3Yf4a2WPx/CASEv7cgLeVjmCqBLv
OgmJCgYM8Qw6wGBBPtXi2SQNkzyHhCbNsQhh9V0LmZLtJtqmxJfSXLZfbcFcdYBbCh4bVb4kBRwO
cQMAeaNm7Fkg9DfizG7nyHJZSfJC7vCm3QTtCAQZQHUG2MZG4e7ywJlTlKOwXyhc9VKcxk5K7RES
MwdpSDAcAuKbSCzot6Xcn5a8mTQ5TpBuCXJAD//Yu6KPXXpNeevEma6y044FvqolaZokHUj5mVV6
vrTcqczuz5b326QllIPC6+SE4XjuRsnGm5qObdB1BI/6hnisG+2DN57K8LtqZpJJvAjRnzMTqIHW
j1kMZM/wElToMGJ4T0J/ljSh9szVnHfU59ieXGcDSxceAK/7FfsDW6rlTCNXhCCVOLnYSiaStrgn
mfYo6Qnu5gB9w+Fxj9xO+7y7/RgajzKWYiHhFL0kOHMRnh2j9p3rWOb1VYT/JtgUY4Li0k3uNRvl
/CGvq40GN6jBivw/3JtOhZY/1hL54rGxEwIitNT6/X9Rp8gLjWgqRSPB382apxKlRqc/JWRv/B++
D7mmsP/dp8FJb6Rg7lm+oabzXtW79EBrdMu2bz+SC3f1iAOmhBsUpxqLIGJsCmp8jDSrUv9WNdA5
1ZBrXmLEaGuTec9a8NHhqG64mAYrCilHhETYgdVgUvC7CcXaXQwF/LtRDlGTPQmFe7Bd9qI+K+hE
tGxyt57M0yxTBLjmS/n62ktk6Xb+15LB/kMMsuR+49ngRO5fBQq2zEL4VOMo0tKdK16lAKuRdYS5
vmlHA0nfHq2fe6vriqWoKA2V5zcnsppuO39RYH2DZREIR/ZAUlpuk0Wy8iOjFYsmW1KkfT40Ph8a
dNBle9x9p66N2d4WeDJhSF0FqSlrZ+vBelFneiVC2LC5CwzM+VdjE359yEDSe6RviLd0EMyEgH6c
3SLQQwXDcT8eYPx3dWD33rHpZ2DHnh6S5dyYGOOk3xYo77Xd5svqTREYrizclWl8HkI0P9siV/1j
9w9xq7EzIyY3wbx3NKrUvtgsN9gwJ/OTCYurwSaNStY1hv4QaMlgZ9Cwgepd6V8IilfUJxqgUCLP
sjrsn64jv1UBMezKbjw6X+foW4Id3dzx3hPR9nIT97bPlbFCO6AdrxSTpnU/Fg1Ym1P0/sGrmPIL
5F8S9bkm5AXfLYhWI3w5tr697bkiZchc4CMP9TyYxFimkHOG+kqVBRoDm6ld6YThw6OtVG4QtTco
qgILr42qWvt8b5ceF7eS9fyt0V5K+nTab6j1YBC2UHNDUO/el7TR+MWMVRZtQhbnMDAafcJE89bn
oysXSqBJE+jITN2atlwPf2r7qVj5JxCot4bfw3xJJ/sWU3vdpByza/6X6ivZwP45HmFOODmfSSZF
wj4nvqjHsZzbioptqFPXnbJ6snoGc0In7vnxYHayqvKmAJ0Gc9ic+vXbdZagPvLBbsinAgu6JvK5
YCE0AFOoQ1t5iRZwFDppvZXYzlsdAodTtx290H5VDiC0gyTbSL4KV7TmKmw7rmrZMEdcvOVxsze0
EE0vEX2kj7mBH6TW5qfXxlHOYpn5WHqjJPYqKcBenYk+Sf6cO195FDe/cPMgep55hscBPKLmNTjC
JyPHZAu++ffq9lOgnlz+PZQUZLZoqCE7iJqTYdykq7lg4IMREPEivDvrypBP9K4QvaM80dM4w0OX
4e+/HSKcsIlOOHemGQxSePlVCUwRV2B7srbaR0c/nZP6MFKWxWMiXupCwhpFxVFSJM9wT0hzY1BO
UrE8ynm7SZ6SpNzzMxozB5jSrDNOd+0FV1E01zfoXoLL1DqGMvzBsbytFQ5GKVxBeCqdTBsCVm4z
BBDZwqMfwZ9o0xCJiELabrZLiCF5LiHWNdaK9+AUBkqLV+cuccApNw89HihZ72ajSPI+LpZyD2Yk
vmO4yS0rDZvR48r/YP8dhgHzwsq36UOTw+b6qd+aPlpWZ39SWt+r/XhgmunqGBsXAAoRb1JSTOn+
LqOMsd1EDxuS0/VTTVx4tMkK94NFPNBhQrFuc115RDJ6vUBYMBabWA4lxZ64YXlCuwS+cnwkYp3s
Zrsbxo0tXpug+HWY2Pu98gr5kY8qjz458Qy2aLBmRXNIHZq0SpNnDEzZeYYMyi4oJjl099WS4yNa
YnPkiY2hTDy4YV+Jc9AiD/EbTTg5E3s4Obj21o554enobj/dOj5HBemNux10Ex6HgggLgz7B6edm
dHPemdny4pvzHd3BCJKTK6tBgTMUoRZi7eltG2Uy6KbH3EoeqQD8UpbtPYy+PpVnL7E0TDdtL8ZI
wPXKqbq5bLiUg6b/WOs1+p6HbJpA8+hjKKVUNLLPIlIQOClaNpdIrDzgJLXFwiDXUh+wNmqw8peW
OD9lW8V84kCAs7v553xtQBRMVm1sWOt+Sd3notMQyfY6MQrES4zekWy9vu+37tEP8hXQ0dXAvhNK
ZlHAb2XyQ55TMEfBdeXxPyWC57h4cG45LWgZ10QoGxd3ecEbqd8StUJ0SmWA1kGzfrnT1H9GxfbL
MK/8q/tZqdMDuBEEfd61ywaBugNfPkhN+K8BOQ5dWjE/RXXkfFgc76dx7V3bLnFOufCg9Yw8bmmi
F4Db2O6H6DG07CTNvTy+2vHoBHImK1v7PgpDK4+ZxSpCeYPoUZAv3eZO6J2kBAl9bhcLk4a9ZX8E
u+k9/c+XyNf0QklUCvE4p1NYiTS6kLALLaHAarkc+Axui1cWys/zVEG79CB2BBcVMy+XiJVcbSIP
eLDvweW8tLfD0UUKrvOyRpdIFSQZxZBIOSEC+TgtPAgLYftbhQNfhV3i7NP7xxAdyZnF/asG/Vxu
+yfkM5To6DzXI9aI/MhvwsFQiBG7QDLkaqA9QZ/HzPQMikszyukUhIOw1ox5k/z49Mz6Gwf+Sroz
aWc+2oY4wl55xkRFuMh3OYEk+IAOnbqzzHoNtLrN5GFUALzlg7z2fpIgA/77EVmgQNmZxCyi0VvO
koUzR65az85kRT5VN4PIit9LSfKYs1UxNIxh4olcO7B2T1PMlaLgt/KFOW4DOdJEhZB50ytzFuyS
emutbfTTeyenHgU0hnuenb1T4oWP3iBwdC+uwWA2WlMrozlrwSgdiILRXaDqjsuorANI/p4f0KLj
OlnPKbzWkqidpnwlhHBnOgRw4zIMPyrlDnyZr/N0NTAjXAsW/SjRkC/wZRH22wYEtbDDS30leFK5
lKveeRV9DogeOpLwN5NZcuGZ+qG3ox5se1DIxB41pYdeuHMAm97TvZ7TqdKJxq9Ke5T2hy1g4FRR
KO9PNmweS/XRowDCW7JR+2s6dNt67LJ/2TpY13k4QsKwG7u0j0ifDljDRZpQqXxnkN6sX0SVL3Dr
LxGWXPQPSMZYnn5tUTDB5sJ+vXdySfIHdl/7cLNhXbrNBDfbATaygQ9qVHpcFB0COkaReA7v+PnQ
W0D+nABBW0LiYpnOak27OSIF6mvJ7Jq3Bh4RywfcbPtM5CMGYhPgDII4fqdxyvhIBUH9BetGtQv+
eu9JdZ7PX/et1ZQukZstSD5pXdxhrI4WnpGHn927+pCQhhdaJTI6AU16VUAHsqg1ROT5qjXJxx8q
Dii2Qqr0xsIDv1oYZpWhkplJev/VV1X/WPviGSVttebgYG5DdGQDIDsSwYjAZkzxaiGb1NyT+aeU
GLsGYxj2URZR+esnPY3u/lmarISBja+czbftNQWpUiEuXVJ+y5Aj8XZqk9uBYyH6YYCQpAd2+NNQ
lgMqER/1dgQWqMttgqPqeL5ntcz4x6ARYxrkM2HlWJHuj1oN0C2xs6DrVC6xVGIUieEkfcl3uMuM
kHP4XtHfBrvlivvmppUaPTOlkLYkrUVpUHlHlfM18m0nmXVSSkhwzvI/u7pNWSUSvXS7l/2pjYnr
FkFucbr8IMqo1BPzearq+z6p/DmK/jDWzdOGFAzJxk0OW+he69xZFda+fqKKB1u3Q4iu57pDNB7m
pK8JrVb26gWW3ctQQfkN/mZi7IXoA/67qYNyMpp3GGD1u/sM33EsmhQwfEkGQr82jY3S7MOrBOK0
J5MY/VZ6w+08bmfTyw5hyOlgYIl1hyXKBMNRBDxW+6kQyiOax78YhA0ZfKlAXP9uu5qZh4jbJpQ1
t01tbw0v2chvm7nYWgdSPe3KlJZ9tlUwk0J4wZleDgcWimX4RZ3JEdUL/d1rAIG8x/hMrl6GYtBK
hogOS0OpLJPAPnEvBwvl43qYCaGgjvGQ060Zm7MtNPbJ47P7NbzLgh4n7k1QUxN4U0JpgQBhXqAA
+lTx3R+I/yXE07oeeKV8MaFhxbuAGEkpiAoiLVZLZqN9l/T4ukOaNYWCe8GewEBgDsTNKUBkub7V
tZaR9YMsc77MCrz2gjnK15/1rH0W24z+sjWcUBjfUDMXqLH5cAdYbEv9nS0pWRogb+wwc26vBNG5
9YTTtnXsnVU//lO/cKq//dUhPaGJixlqlE8XNHti2snMJMwn1kaYQ+UN3Iosqz5T8gCY52LWmvf3
qB3stqeIApi3XA63P45NyrgOiu+273wVWWeogy8vABdnXZXAyMdClEN8WDwqTP1CvOXrBQ5CgC7o
9Gep51afSAGDhhus4Kg3Q0yXNYdyvLFpCF63w1/873DiIwM6NZjeodscxuSpMBoEIQGrOUOKaKSq
EfKhOxCSEnjbA/5rvzldvZjAp1jpgy6mCdR8HhTuWqHxVXe5mmbjQDb8CyX+sc54D/XwwKi37cOF
7LyqZcvd+zhclOuoRR1LBWfwUrfcJQJgA83A6gx+eivRKtExFtKRUJFLxWlp0MKCU/Dm4zwGZzTF
AWt4mtihHTPBDkvywTYn9DZ1zE233O2YnwX7j9GFxBYY+IzunI5gQxnOimPlBvWMnqVJ0lzSO0ev
HaiJsq9wpHj0uo45utFh2dI5Wx4jvDq6RPyCFk85j3eNg6idVcM3vGUe+RCVczVAtgCWmKH/HMib
y3RIe/uL7T+1X+chtlstdk/U2axQq3icVEIyoHqbg8FvBwp0/co0Shv7bDRsXUjpMizh5KwGAuDV
P8yZmZpnegY2Ca26xZmO5uA4rVRQ7H42bhTAkqMhjhm35zCvL0GmH+mVOqTDTaletJnK076Yl6zO
3KIFlM+QbSwY0yimD7NcEimVQ3wSkrG/6TA9cvfA51SKfBvkmuWOynSGkjGEe35mjaB/lCeWq0YZ
Z6mV/Vm5Lh+rrUTKhWzECFNsZNedxViRhiSYODQn4VA13hhC0xZj7QR4T0u1EyeJ5q8D5u1+DIP7
1EXH3hCxQkv1Hc0TqH/0pLqyLJh6RvRFMhEFxSXPzVcmeyStO+V5Pm+1NX1H/nG9PXiFiuobkc+G
coeED+LMNQnggSvhijxT5q5hu1K8WcuAB9jPz77RNHzPvVrI2M7MnVWiSmFcuZxLeYPy6otMsWtn
KIykcem85SC/NXV57MKXHKjZCqRxZCn5Yi8l6Vtmu05eRgWxkU6BSqZZpggNeMp+RaDJ09vI59oc
1Lyv21UygXROGKV3vLwtIJeyrQAVoXJTUufvp4o2VG7IZWVSVtjNRB5xVwqcX/18lC5YmhyJ8o3v
lHzQcjilotQOvFeBm3y7cngcAGZBGabVrdxgH04hDsJvPW8+I13hPyirB80d/vj8A/HJVgtBuryB
zVLhKxLohCiIhWr7aug+hx3b2FbdzuJxd7QjGvymVOiCqC+/ZBfjFOvjV098lYhw/YCjH/PJCokX
d8p0wJdo0yBdgds9LSe2oC2+X+tjBkkXijTor+ATGRhlREYiSSz28Go7NoEZP5dAmrwPqCMr+LwF
po2JeAWtXUgrQr6wxLsGkUbZf030fCFeJzS0Wv3QTNRyQV2blArR9TlyUnOwIRd8wxfdAAV0Ftw7
6cgFo7iN6w0q6pPvsuEMo1ZdWc3r4RkkKNy+zAvSdExwet/uZH+Vuhc3zbtTvzzVRyOUvEqymVat
qmOFqzVmgH3kIIKObdXhXI4PrBIdloJ6fE8YRDptjLFXzKmUA+k1Ra83K/O+JbrACEEcoMxulkiU
ibMTtAdejZ3X/9u2C3ICRCtX2I3JJTyicycSB0lhJhMMjWFGBm5q0Vm3PhP2qROhA8HmiJv9EiwY
KHGvY69g/Qpu0wn5UTzzHI84VW5ruiEfHBOkKAxXybEIqpSr3QT4z+lRCeUiv18USdqxVxT9aWd1
DU7w4rQisQLuri6X/5MnYQazzHCMA9o8Vhby3VPlnpRgf0kCJyJlCcdH0tuXZa0U+2qQkWBt45MJ
IJHWaCU3+vBvcni4n3nyo/5Ir+VDhd/LC92KDWEwSISzesvwyE2hyMNaJ5fNk1KoDa4Pr4GYvBfh
rw21OYJPib6Dg05kLk4+uPqaLeGp99PUQ13zFBFxrjDvx+VCVYuYAG6c4RyIANMvL/blmbvRz7bg
3nV/98WBeNGZ+GeO0qTIbxeQOqvCOoHSqeMkn1VarAo9lELNBeNrC6V8bZID+M9IBhNlhhpPKTF/
Ekulj/Dpyu1Rf5Bvqr1/k2NQwDNjeGnjYt09y9IZ7MMDzt2SBfCvBF/SRSWZPgL1fcOGeLU8fp5B
Jgkd1HELmXy2NDi1DAP6ZcIRJyrSsJXzxFovnZ4p74WoEhBUTN9onsF+Wlc4Of0LqYOtPB19FrIK
nnxW6gt4hotloW8N4ycO2OGq1jD7mm4TzGMDNgLh4jeDN+s95rY6khBZ6jSaab+p/rCF0ipCieQC
85eWDIdGaNvCe9xkL8H76dDcER28mQXdjnTwWm4Di+Zd6ZjFpGehZ5L3m7cfAB6JZA3h7/oVE/iw
DCUiSlRA5VHuZ5RD2roKqgHYI7oUZivk8IKcO+xuq285xgOpYYM7+PK2WBpLwTQj2OBAJvKa+S06
zmcao05Am8c50wDTNsoEXhv40zmOiQx/GU1+SQa3TeFUnJDSFdJS+y16rBEABPXTnpEyyqwAX99x
H8j3FEZUoU1HHoQNMQ3/WbQ1sHs9QMDanwmRJ/IUXkq207aiBL+yncRdOakjirPqx4MP4B+sbypW
21PVTkdYwQpg/k1dt43unDqB9j/pMXhVSZBsMiQALpI/PpvMZpQm+exZd1UZCcDysGAPKXA/MFX/
Yb38ysQVU/bouilgIMRUDpZg5K39SKNMqr/r3y4uiXV7uxiLSU6hQHaQ3m61yK94NEhq1tq6X/F+
SNFuDKn1q3INu5gYTaNwF9J3DZ20DECMW4l2SZaYUjxB9ZuWmbXPu98k6ZSOPRgxaB2FR4AF6Ouo
r+MHek03qEom0CP0o5DymTZkLAxXUE4oYQ4stsFTIwjhyZ1/I715OkySZpOrJlzqjoOR5g1jzpPz
g6tiR/mNK9Kg+xbkzIWqhPcrcVaDpve6yu3VY4TWCkNJ+7Wxd9Rm29SnxBvOc5xvvA9iY94YW623
8D0IBtPFzIE8HW32BOMK1mg81HiSWp8rpOxRpXcSKH9Vf1RNC2NL/wAGk4C4AU9FXiE+1Rgaee+b
KC0VPP8sUgDFfMLyz3gXgUFLEjWR3rtfHysgj9K+3v7aUHMREcG1tFysF9S21XmTcGuLYv1plca4
/QyyiLoBLFGdQ6xxlI/Jn0NSD+U4OWBfcG1IFjx6fotuJDzTn938GE9b9U+tzCXr76S8dXPb8kk2
WAR2RfSooEnx06OnsbVA1X/AyP1l41dBTa+8yQvEfcRef+kJtZd+qsBjT6P77k/Ztb502BnR+WoK
BVilRQzSihbES+OAl9NK9ilipKHjhGSZNohECaqbPWMb5YSiYDa5xSioYOoIllwLqIBRId5wPxHy
vXNiQYcMMu/G7DuBBBQYDGm84O87RYZ+paYRrQ54973VLs/kFLSkHq2cFyuhstvBua7NBtbxXlXp
jngOhKOw+gVSDS6cerZHUnV8ItkOPZ4SL4ef/k95BU7YX02B7k2ESh9sctbSI6K8NP2GLaUEPK/g
JEME1gkY2pNJjSauCKGhYrJr6EoxUMA9Joto+zunF+z3L/BvMpfDw/nEup0oO+rnh5iUzakB1sRb
p9DKGTNO72SLsuNGj3AfastLRbPstUDHMsLexyVcFnCBM1gBfnPoUxUSrqkM8DYmiol5eqGLJmNp
iROSt58MhrUwYCAveyNXhzRIV6W75xHeTv2fSWDU3YDN2H3FJjRT8+YZEYAiu9jTeyT3FIP7m2dH
YcrqBd6m/5YA8HPKB+NAKGVBNTEt0gfZyehA7wTrQVwVbp1XXlXfxucmDNIE864Loamlm5jOEe6n
zcf3lnTkAmBJRqDkDHmJCff5IMPS7eLjuJ7q7+d6W7X5STNhmt3+vQrJKA93Ywmgv/sF40hNNH64
zb95cl5hqZdv/1M5NZossEduHh6gMqf/KYEv451gtVl0lwz08DxgmHRB9ilenJVL6dngZnmb312T
D8H/5MzXtWPEd38bLNvWQttF+/eTbUw3qM8AqIcRU3fIday1o61dUdRjVr370FCK20ExOR3JL5SS
lVxojsBRC7Iaae2BgmNaDosnV3G9cJ5rXFlb5VpTUC/f/qZoGV/Y7XkjXnPnomEBLy4BH54vtlQm
sFcM+e4GCxK1Zbfiej5xEjcovieIjjb2V6E3TxE2t+Il36Xa9+qYP4xehURj2FGG/qXND2ElpOq8
+gZDuwZLDNbR/Rl1Faq4/u0o3/kGgZyDLjLXcjA15SeNc63AQJ6e49OuOm+mKq/UthHIPruVEzNx
cERZ1hqUJTft47DG47CF6HSjPKhI/TEMFttnVtarCylE90+jdke7TOZrm+HKyk8okpszEAZwnwAg
+ImksKej5HFPg+GZn6UYJOqGmq1hPbb1aXRhO6TjsCErtrOPQ/6RmlUZgqu06iE/5Udj08f49u+Z
Ca82f5nPEj3TRoIWbNQNmdoaCKNP8JOGgJJ4uec4Gc/EgWAPizuxyAIa6MFLXZAJm+wr8Ui1N6P1
sWXWrlst1Hdd1DkiJYc+4NN3Cf1XKMA0vKQIy1UH0sYegZK13ye4KiWHKFfVt52LNAzJ30pYm7/B
CKcr/3D7n86tn0Q7VFE+kpdM2LVCI3cufEkfAZIvnIKxmZbCsjIURwdqTcxQKnGd6u9n5F726BtZ
4Bd8w80TP1VJBtacquLbRfOQW1bZFaxG67vl2o6NHBl83hw43so0ipJpmx+pwVJM18daHJartMpu
iVgxSzT5wW6EKYyBDPm94Or7xnzn6o9pBcCXYVoKFN6XdBlclb/t2nBODxBSyGxEdQO/k9hjJ/sZ
HQ4ekwCYwZ17+/31zAA3QpNVzkU8nA9ADESrzcRMJx/6KFXfhr5ycGSNFEoGn3PQmad/il903N8b
7hZJ0vJ8anK08UV0bsvu3Dn7XeDVVpm6Hr5IgfxriTYOIquBPLldd4E3RISjKV26rw5qWxQwCYFR
M55ZATmU7KwCm0yjYMtpY24BIsbNFbqxzQShcK06p7XJS/WD5FxY2Zg0TjQHKQX4m1difMirX5sb
abglh4PyunhzFL8ZN/yGGso2U1/ctjZ6tzZSy+F2+olSErn5T9OpzK3luElPtorAEGTQy2toyCCB
qdS4KfU0zjT4o71Yw38DuJrVjfJN/gv9eADretB2ammuqioPV4FFSwl0mX2rDF7o4AhvsozP1xCf
rBR1hhhgVKjrVnvTwN+HgYqY/35QDqdlBFK5esYffW2Fzg6kTUtzrOf3cv23VD97tADMbZmO3ZRD
7hO9JUjvDrDq8BBP1tkyABBz3NjoXdjz2ZnQqlbmIvaA6lBGnL9CVe+8bECh0wJiOVM0Uj9I84Oo
ad97CynoWCyNq3Ggq1CeD+NkuuZec1eEDVAnsS7tyhO8rfS+OH56B6HufDoco2bcbNDHzV5XrBlL
gyU0j6jLv75ks/HcvvooZDuBJkFqEYRPVY0GGDo3xt3Sg9Sh1fcVPez0pi5gF8w2cl9uY48qin/6
kKTUJ03HQsM11DEdFIB6j33zdvExaYBP/hAU1UlcHoIHRzP3q75jvpCIf4sSpxJG7C78J0wEmuue
nITofc71Oo+wrsYlb+eBJjMnAJ6fwhUQvWChEuXzZddIvr/IjWyZkYOv3102rzCX0xdns9fQuF1Y
9CgATRUf0D2bDDDysR+qIIJ7pTL0DEegwgEwaquuSCAwb+sJmsBR2D5ae4dcB1+C4PED67nNc5LX
q4Ce70Wa1A7ur1bazrqHafkpKIYGay7pkTW2FVUKE/2N7NMe4uJfJuv5XYRBsJI+3Ste0DPMbopv
0+OKOKNXQmt5jiuuGRRQJH7G59LlKNNb3gY8aHvOeCqy9VLX815DkxmUlxSJM09S523HAeuqvXMQ
EbDZDtqFNppgeQesxYHFkiBH8OG6Joe+EmzoF7DMknryzfi+DW+x+SgNjc4p3TGYrA7piuGIXq6l
A9tCzvx9zQLyDs0p5v9rRZalhoe3D2Xsm1hD0bVDswD50VqDVH/DvnQb0i3PWXECl9BXbQrLgtCY
49vdSkvLzJpvNPPxsBKKe8EKa4jEND93LBtibAt30xdSfinDu+p/FEYHFodI7iG9XH/nVZZT6Fhc
YLap1j8z7ZQaVeMAVBqioaVwoNx5ED9Op9zWtaCUrS9Y9JBx8PwQhKtlUIbLg1iyoBtyk12e7KWy
Pg+0Qp2oTZqLvpq/wQZ/WYQRT7t5Pl1CY2vw4lFwfbNI1gjFWSeCD6pwNJEzEBmzxXw5NtsqBNfQ
yZhjkNfcp4zVJX3OokHAixeOYhzF8HRHEt4qXho/m8KA4dQgUdIXeENBAPrMHRfPSA36u62Gy1Fm
XuiviR7tLm410j8zebxLrTwvRgF92pWa0TeRWCw+5BjX0dppxfZqHhDofzGle6WNuFFRIa9kZHko
3WjBwydz2QN4Ne1eH8whHttRw9q9eGJ+rwceRCmJL4+AEjqsqfbzAGSqPPJsIJHZkRm3NM8qcOTL
dCapb3q3RCskry7BMg7N6ZG7E9/bMS74u0pRrShG+KRDi+Psmp5dUgkl3sctBbLKUgs+1PNjFM5R
6pxgT/FynbAcBOCFX/Gtcwg7TRhAMmDtx1AI2FvqF1BvfLqiex+PkFmZg1TxJScQfyDr23YlgOlD
uu6cNQzZrgyrESxixLI5IjiWGEG/dx2bdElXHDDm0xAtpKaiCwRtliP3olw5pGoTN1FtAl0V1g/7
9X8t/B5LjzH3jyUWsZwB70935SBIKZVLFZPo/UmEAkXBCgua38gKUgofn62NWbDbiqul489colCf
ugUAiG8+s5cJwTMLw/5x3TJ0fz9CVotPYhU0O/hJRZFASAVPYxqiAgVjFnXfHGZ07BuX2I0W4I3I
2IW//FHw/cGh70ZFDLvCHZ1JCItax5pUZHY3Df8hglvGBcbZhld75eaq1RPDjJMx1/d/AAAtD2ps
95FmrtF+mmYfmo0Pt5MCSbDS7UOBWi2gKgdtBSIbx16fhkLPgNFr+PVzRMl/Tbt6vX+3M2yU/+sb
ctQozSOhLvzTrDscBkzJv9Z6QkTeGZPT6w5j4kknbpsjkqBHisDCF1AbxhGuVAMrSTI3S9XCkwpg
jSHCNC97pfwFklXtvtn2XlfpodA8VxsVwacKa6d1koYbNJUDrdMgxHZuMl4Z31038hyYoVi50L9r
2in8daBIhMZqDyj1ioLG8heDZXYH+hGiZ2UOINNnBnUOlskHv+e2/mLIrwxAwnbF5e5ULsKFcXJ2
zffe1DwcSy3fby7S5Wwbq572lQmFKk+0RqEVCHHruWETqEGvIKyhTEkb4lFDe6BneonQmF4ELCCW
PPyWPtDSn1xcnRjbBgOMH2drp/DorAsdOAcLH210uLFG1TkDJ/Xn09ZN9pJUi7n1CkGTImCqCAy6
XJ39Kz+QkwN/bgkbHm9DjwKGMo8LFoZNeiJppifV5NPqL+1dOU26xAGrTeyEgHnQo7mXeeJrvVcQ
B9Ksi7mgpFnbI5UJnlg+NTaVcBN/WlMgxF9zL46BUcvB322xzTw5aqi74XymcbanzLB+0LroDq3w
GXvGn6htQXPkZbWbfzhRdfo9mhgar2kO/9l3rCDCYF9M+521gJH/zIsIl9SYHnkTpj8wWdVtsQ3A
9PeEuRIVJs4hcCX+s4VrwzmRchXxzSBjAQ7cDx7ldFEkpr/3LOMJYuzNECSfDQoqWwrLLF8MTOkL
7chN3Ctnezofv+a+15ejyIaNafPb922c1HgPXmcb9NSema/0xoaQJh34ogP/qeIDoux2V3PyMakn
G4kO208O6ThMwwxT+nlPllLSt7oRqQkE/tHa1czbHS/O+Z6PcpRzGjBZp0mkUROdgtTa+aUyRbCe
YMhtkbS7X5OdA/LHL+zDqm+zlNFw1ox5dJj3IHRgajYazNyDFYH7kAn3PhwtmvSB+dkQRALdE9Ix
JQH8rcgjkzHmOh2DGCqJZE/MGGRHPzZgz1+QMVvAXkQ2urpGWPDjbCJKzB5WWJ+mkXuaVQv5IKta
Y13zCxXma5j9DW6LKDEusLnV0zu593U9la4gIAKns4pQI3y9aiOCGsr9x+8JHvrNCFfnoW83EfXq
RFWrHsbSLsOkmNzIB6v1cCq4CYORsgWKLPJ6QryK3KgTki9gIA1vEjQ4us7t9eFVv/BckK7BRLL2
JP4dSvHcQjbeF0KmearC7lNnvYFc8dGdtiJFEQaQNRGRa2JuGgUqGMPDR4Qyj5+HbSj6J7i6OC6W
ZasNGVfGrbbwYW+fLYiwnM4YL5hocjlL3WT4lWNWj3jYFxgOcynEkiRCXiwZMQ3TPdk5p7kJm6kL
jJb2RCfLxr5Q6RhUbMvAEZYKLvX4ljsM5sXds3IPniXKwf0aJW5qf1B0hCVRPehErGMdoEvwDQPG
qDI1p4I08Fmspjn23zCt/6fuBKJdfA6prr9vG+zVxo5dez/rkhOzbNkEmX+QiW/Z+Raeymtm/BPt
qGcJGu8ZHUtTB6MPYbJSEz0Gy2Tm0QrHm3KwgvqrDWHxgPAlrIPqPCkEnY5TmmyFfwX1X0PLgLWO
M1sml8BmGH6+pm4nsZV8qG3jbbivUqIJCJ/cKFIS5DbDD302kNU3AaGHbAubdq/xxMALfzPi76ba
oKrrxf6/RdTje8bkFi+xNBOYJjZ5MnemUA6G9f36pLDoBb4U6RwCtzFjjmsSzz3jbUfFZAj6Bw+U
iaUY1sGb8emb5zAAh5Q7NLs/cczqSLrfIpuafe08sSio91MIAzdw/2oTsRidt6B2YnZOeMMkoZcU
efjCaBCAHkJpH576TYKlDA+DFSj14x8/q6NR4mjFb5ONC9Ju70RYXINWwIp9Ve9XtIR85/NTeIBP
joLvrUhacbbu3Q/EeiSmuxhrtkiE3J+2vscuJWT4TOgsNjZ1UAwT7wy5BAj3gIpLv3fYo43Z04SO
X9Oc5pl83h9EwI734yvlpn2rD69P1CSpzp7ko3HrPolL2Atth5yp1BmIKjWYT4VTrQdg8adeqXD8
6nsKypv9qDb0denhW0QMl0Xq2YA3Bfz6FaLa5WEYVgZbVkDNh8XjPWmMrrZr6+JMyV55926bD66t
Pmr2PhZ5xEIQ4uiZZ/Z/Y7BjH2U1MarRFg9vy8+IhN+k7JXbBY0Iz7RTKMzSc6ChzcCqdfp6D5ky
NNstMcdJuDFRFs9mz7QTMgv/TNI6Ynm3yuPaYnNo1BT19xjrqz5oUdA6r9+CVezi99nUtykduBb/
5e5pSiLQe/wnNKk9WtCUNdRntfqmY4bNXMteAyRzSRvh7ir6krOq2qowj8SOVKbSZsg7bNyQzAt0
dsxl16hMIk+RnPLJrKSSVHcBNH2adwsCsLkW7ZJIOI3QTBb361QKsKwvQTa7LB/6D9yTYtr+jYUc
IUKFgwY2pMTHyDb4GZu0FcmwueorB173Le0qHyPXy655KcudAS1Kc0EEG49pwOv4G7i5ja0MpDFE
wNRdeeQXYA6wbMRnrAb7ea+0pAVC3owVYULx6fR9T6oySAs6xdxzkch0pxypLV9Digk5fbusw6i8
g37KMTtk/+w4SKnyfBEYcnaoPKCb9yOKBqoFb0mb3GE72pXL/elwQAz+tc49lDCUZs4PQBx1hPMU
vtJ1Ep3zLuxxZrUggoTZvdEws95b0zfEYjOu4GzleiUHV+aFVuO6vMgDwGJ6P8NmkB1TeW2JbFkA
hTTS7Odloh+2bDr+/uMUu7g1/h59jPKpgts+T0Pp7vG2nyGrmfaJptvEdo5+l4LWgVqilOljBcXu
Vlbg13lVrkB3Z5io/n5floz7xvw4rJ+JFvAuqtI6ZISBs86ao7kANjAGEWq2JoS18eKb54a8d3tr
xZK+BeJfsCGLc/BjY4im6CFp08W4RlnSr6rESjYe+79r5HMhy3bo4KvnP4pFMLDv7jPk1PmiM8XT
bSW4Xh21kfeINaeM6jen4vcRE537MitpR47Qo/UVvOqlyKc9H57VBYRk4SSpBdCA9KxJme3+hxlr
RpP3EUCq1FpEXeT8gy1cyaoDq8EYINB0Fy8tLfudacJH54q55j0Bm0/nhyLaa87hCoEA3pCSWbeo
tfWIYeiWo/ota/v7UCHPG9kAe9KIZ2neyk4p1T0dkIEHpfYzqpnRz4xythOjS1g0x9NsJuAazAdm
1TYtGz8xSqrUnYipOvb55FQ43d/zv4abKlpQz7PeSnY/5CDyBf4P2ZiJBeLtekwZL7DuWTHfBaOA
SqbTEwVXTVHNWC9ItuRP4TPKsSHDJecA0OPpEwmXMLBC7KTCZijOeLDVo9X3DPkuUscwZmgC3Y9h
KWWW4UY6p2YjwPox0Wl9jpH1mFxOtdBwBKpf/UlyQ8QqA/mdPeZ/NGMjTVoLYUfH2wzJmnLBVMWc
ApkkW6sChOZ+I8ne03bus1r24+qXsMDPoulbllCYO7VvGROb1E0IeKDRqehJsxsoJjHoks2IO4Ym
nY+Ti5ZVXPsm7jOvxRt9hD0mXzcy4EN7NfSy5ZRkScUS5ufCZY0BgEEA4HVRBQTMKQZm012/Wv4K
sBdGG3TpqSLbY05Bd+LMACVC9XxQaXEBmNKpj7FWN4ZgS5nuIczNIztdjf2uTDhCi7E0Gx8dfiJd
LueKUadZZl569sRDijK9AkNm1eI0Ogof2cCy5T6ZX3tOjZgRepSMZPoEeetQVkngF11uYxkDA+ga
Ud18iC7KyOyFxlA9Yw5ym4boRbESqPRlM/A729sMhl5s8JZc3jzgg4wPq717djljutLn8YxqiIOm
UD9miNdKmh2TmUh1FSp3Y+uZBUoqVjugXrxbhS2mC5tlH5esmd4lLiq7tdh4tUw5pIXetQByYkIT
HxhRnA199i/2BuWeE45WQzoR34yca/uMwbELR841reBRstIJqSDdUfNBzByr+Ym4Uc2INS3M7F/J
Y3E/7qZH3nZc8bMAf8afQlburQmluBHqyr/IjxfMS91Nny8f2d6TPVOD7TukVKzwIzfdROrMav3M
reSHkXDNC152wceK1rXChBZGqPjDb95ku1ZAM9E2vrrYWeOeKBQH9Ay2Y5RJjZQyKkQQnAr0+fXh
xOnNxJ3+9HVZqYz5x2zqgm3hiUi5lnjPOd/mjFx++wGvE0T+3uynI4RDRuCowL0Ub1Bbv+eUngeu
vJ2hly+ukLCm/ikl240wipfnO1x5jt7JQ9myadyB3YFC95t12EAqkrGl/BuV1bL6bAXEaYd8+vlK
Xo3fqzzCmhQAXFu3/Wymyc8VUun+Mqxwti92ULPeJCyI4RZ2BGpkjoEpj6pnUZaDxHeIovKwL4Yw
F1a46hnU6VhXUgM1MWyTxNIg/uW6syv8klAdsZZhVVrS049PS81YdWXDZbjD8++DTbXcne3XeNw+
ROyTyy09pt0K7eWtnf8rpXd6lFK689TsgScYZllYvggWlsxdjnHCNLj5kR4qc7lr/Rv9mQ3Lx9eT
kK1/edFUkWCpLe7Y3R7v7mVY8FVAYaBvfMYhY31qDrkTzpQGuzvq0En39DPBTpOTvnC16oPCYmqQ
1abf10frTHPT6NlvjLr07I9kugaYO2ZqAKJPg2YbE8B0qs1QiueeAF7QYI2ixvDT1WfIh6m6ueJ8
+qQju4DPRy7OlysPwTx1JmSU365rXCMxEepU3uSyE0kKSZine9k8GkLImr49H+G0BaS4X/j6rWmw
GueVOLLPlFHPxXkHa4W9iCTN3gW6Y1Hi+ugQlGwZTe1tHypgx8D+5StMsx4GcWWjbds1Vj6Vw806
YGPbmlUmpqC4r72blohZqkl0jInr4QG71NHDkJWmasZxmN4qxbmg1XP36NMKkBCkwtOoWlwXwUVM
bnDy5DXWOSXDaDc7/658CCS194invZNs3zQnLOR2NN0Xu9L4BbD/NyJCH53IsdRFjUa3vygqUga0
8dlz4T/Omgye42DCZXYFpFNgkQfo4y8uCOZVtbv3srGAQmqBfGeV4eKcthW2vi2DOZpq+6FNtI7K
TS/U74UdPM4i4OXQuUyFeSDK8qaZkiQxX8cmK1G2nHOdD3RYmVJruXMdLcovKDcyXU9Gl2GTyWXG
Q4KAPYwSWTJdErEFP32iNGlpTPNkIThGe+JjHdmgLZMie+r6qWXpZFdxIAVud+VZDTMaRVSYseIx
HW7ABf3ecIO1aLIuBuY698I4gyn9WmqEJZxlHJzoS35qy0ISRnGhv37XuMphC7LyOEJA95TFGk2I
PtrTqJFn+eULA/tngZqyMBr6IGmUNLMMV/HCL9H37276fP+uF2mBdZLhrVBkXTn85bPHCXuY5Byq
a1P4cYYi4o/qjqbQL8Wb4ala4eo0qx7qE67/AA9Ws8H8qvj/WVt+aE3uhZS2nthN3n3piIWrV8JR
hsFTW9QmtBT93sZEbbVXD6L5k42Q1IXdPrT1RzEDPjDdKe8IxKTTozdiE9Pt/Jc42EReXV8hajHj
JoXYjNOeWbsVmhjhyAOiTIhIcocxjAs0bi2AX8cXWFWUK/+hsh65mQNQ8bG6z94W1g6AjHpokkzH
cNVwrVFLCgr8ViO3TSz8FE+VlsEw3fknfzSMJhe2QD84HqR91gCll93NtoVXVJRJvcouhX8eMbig
QchNuo/NDCdxZ54jTk2qesgZv5st0PWoyT4LF1zLIrIiqPerj9/q3iK755u/BNBy0rHNnE1440ID
2cbRgLvniKxsYQc0llobQx9QANPAHPuvH0JU4fvzxpBI9ILvGRMtVLvtjzrrliQ2drDb9Ht8N7GC
mkNcBzThjxWdadeLIrcO6JP9xByyH8SyZMrGp8Ir89etSVLZQqEOgxRqqsV97yTfD0/CoJYUjZJs
A3NOqf3uqOJIrmqu9H3jgzvxd7p8ACHj77Z3v/SYVJNXVv/cX9tU0StofT30jcYDh5ZHL+ywOyL9
3yaxUED9T7Iy4ZaEasSnYrx8mOX65EW/g9y57VMt400Iq3GwLGYKOWGOx5geDwKwuPRACuXNxQkq
rkP9jT2zoDTbwDEMy9veJPuaWKMZSDjn6mm6ttLDsc7RkbEiuJd9/M84QRlotG6fNu5y2nS5bPP2
bYifjTd/ML5IQVyMwz0g71tPXrlyArYPUznVaMDwWVE+vOQ5576LH0UQt9yFFcgkcM0IAfFIu7k9
XKkPVMYVuaRHmIHlggtN51Pa0gU1FWayGzefRRF5uuN+dwzqBEGruVYJfVkkaovgtzGxj/TBWUsU
tWNY3SuE3kzFkPWy1v1rbL4FX/UMGymKEWseJyC0aDXQV5KFhGJNa/h5Rkd8XeTIuG0Z4dQm71Ma
xnI+QoTMIHrXmXEIXCO6zV4SctfoQcdP/I4ykysgxVOl3m5BoDpkjsNWhw/soh4KrgUJBCTxtwKi
nCqULIEw2s9iYMJlmjRUaznsWp2bgsmKTmmtzYPjXQQmJEeE/7f5Gg8XKdYpMPqhBJMIVB/H5LaH
kRCJ3UmknGqcvuWSTox9G82ten9DrhDo5xUwY1J5oE6OqP8PbR8oRj3Nx+9nCO6LL13BFrAlMcb7
KANATmSBrrFtLimN1WoZUKLFWRkhhQEsV+VMMjad0TxT1w23bx4B6sFqnwxKcVGzsHa1aBeyE0Mb
LReVptUQobNLOxCPMVWjZS2S+pFUI1EJXJnGCuSzqBZyJZwQsibVnJYSHhqIoZ3XnP52F+6Hb7h9
uVpkVdXAX1oBnHqmCl5wTQ8KKqIhnzm2Q8Ib5wkY0XkMyG492+G8WQIFRIZLPYjgItgyDOjJMq+x
4lzZ7ooSN2kiYaR0pI2XsHX/c9W2UIjeq1FNcjjinb4KioWFIScD0hmvp0fL7DoPKIGT3CSI8ilO
3z7HUR/GjoSwVgSs4HTTtk01UKYdm80DMX7BjcMPlaN6PHhhe3AJZ+2NvWw+0Dm6jJoRK0rk8vHJ
4ekSU4lF6o5le69cq2L8Y1JlRGWRa7Dy6ZpXP0t87ybTCibgBe0y8/Hrb401UkTPh4wjW/jOvJyH
RCEVWBjOuurzL9FKzzgsKJFjoBPrmUDkis3suBkN9upRZfuhVPpF2FoYVveZ78XnW4YXj5M0K17V
LEz3VsxOk8HFmY99mkgpOM/2IDxvN05EV+pw8E5L5TgnQ0pb8khFGPoBiykN6J9h3dV1maF3h09N
cNQIeiTlXziXUCVpNVdrrO30NfkZ/zo2/Ko3/n0EwXKG4nMtPRHVpU8SMeAd9aRw7l6k0sV/8iDj
k06406x+am1BJB22Qi3XKKljTeomgNmPX9h67C+zQo0jCNpoD54KyJ4CzmjOqArlGsEup722qRk8
vvjrZlErPOF+pyzxqCh1Ds3tb2DSnG9CaeUMeJI7p7T6ICAaVGoIovusJqdw8PgFevMHCQXpiyi+
VDqQ6ozff3USH7lE0rXZczZSz/8i9kmqUwcjyUxI5ZcIN+b51MTFQm5eWzESINadqkNMAsxSMcWz
ddn/TQ8M6rKWTSfAiyAy7yi7M6ut2KSyXTa3qKhml7fklgUHgDa0sCyKrqY0LpFeZUXziIFAPWDo
SqKp6TPNs9qwYlIEXCk+yi/COop8+PU7/MSNja7hwEN6X4Pnv5zynrq+pOYaLNI1cHe4d+anOvth
vPs57j/NZkNi4V9eTx1a7I9DpymT14OusiQO16ASyC4gF00Sr7msJZukyBDegiI8dA8/wQafxfC/
vluCQNqoWoVr9VsEGvElMsHiQ0su/SngWA/C3bdUbFJWyQyozOLME5Kp4pZkDNcAO5/899QXQzMJ
xs96ibY+f8Pd4qO0v779YAgTxlPBEhoIBNu77lJ+QY6Gd7nJvBYYV8mA9MCXxJw/3U4LVddLXYtT
h6bM4jDVXymp8wjGTd8NXzOwEuBbdRqDW7wght5/JRfo1MAaSF3lRsvw1BdabD5xgGjY1jS0ro9H
Qj+L5/n62qszQvNXgIQUQDDLc8anljoymY99r5kajScdROyU62D/XpsSpZuByIBPJqLlltAB4Dcd
KfcX0tOMfAg3zDZBbHP82yj8c/9IrqBZzsJCaMV2CHknnIsXE5wet/eTqh1wTYPfixDy3Ud9MmTo
a1GgSCpuOs6wvs3uXJm6jGrL8GPRyp/9aEjVl6jAaN5jtgNI5YFNb1vlgN4kQk3+DzIa8qvFiOLf
+o+1TfXAWd+Fhi3wp+OBnTJT48pk4ttjTWnCQzPPUimoLynQZxnHl91kefcNEuPgDSm3Lmqa0BPb
rHkxts3ufxFKG4csYrcQEAzuukPWwH1YjRHJY0RbuFkiu3HEHN7djM2DlEpOeVHjiGiR/pPZsozh
N/b77biDUSjrwIgk7v6EaZ+teVXAmbTobZCP70e+wC4s+Ddh5pS2gHxcaUtgdvmUwxxyEqv20C1R
AwS2nXVvSWilbVqoZ+/FldAqqRJIaUviwTdc9X5bKunqLlYQ3LVCIGZewnuBFzBbKuPrA0/hnfP1
MM8QCHf2/kRdlOG265gnyxMuO06MswpBG06Zl4wXZ1s4RtcpAfPBPnTX4J9bKQzVfGgOtVWZhYbt
7zaRCoY2TTP+MXLjL0umLZrrrwm2Lg/g3LvSWmtDmdCg1DTvot4LxogoLk3nKhMWvEIs9wH/hAXh
B/4y3IJK9NT99y1hQG0nedYmzHhXW6HIuuRYns0MLYE+2b1s6htpenMWGqcvRlKRkWuh48tAMPYd
0Zvezf+0xr7yW0/dnx70948fNyP98FC3JTGzfc0PhlQ1uIRx4NUuBQBwZ72Si7r4q9vUFm6Jy6qm
aTaVIpXq5iGvZflTjZmDnaUlYknSZcXWR59xEqLFEq6mRw7ywfvz3BxtWwEkI3llWziA2tcIOppD
ePZYfD0KSLq5pU+SHINRgqRJfjIE6t+2+oVZT4TxscnA1jtFB3lBlra+rGGMyqWII0FMdVMJfjbL
pM9gD/t05BeLue08XxhpmI1+8MK+nul/dV6pYE0dqJT4Ib5joFfa7AUBN5WSjCBwfC9FdNCC9la7
/I9wIZeT88bjvdp2TaDSBGDVVLeiTols2Fwiosqz4fJUZqxYktLqTy31LXenuLpkvHZNceAvh+sD
EHkV8wsQhrfD67G1AjIzdH9oNmXJ8b2ZadlVRTJGNZB/RNwlqLQkQ2xN6kaW5k68d1DyUudlaPRT
aYJ3hTOx4ZntPc47oI0xQUrKo5WvUmfMOt/3D/nR//PajpG7ybkFIO/X6dT94BvhYLGyOp74Nb/8
U0aVzCJM0WzRwzeLPTy6Ns+s8O9PriyeaQutlQPNzjsCLrG3v0DVdNT5+q/rSa0JbVo0jgNmVtpQ
S1cEZAFVgAPwZjBgTCZdn4TVnhPoV7dIw5xlN5LIRrTTCbcab9VmkPDMbuzwktZ7Db9nKTzwz/Yn
o/1YEHclxCEP5haG5CzHxY7vu6XBC0RcCdcDUIUrMM5G232e7IVCKdMDPhjYV7tpJVvSLRMkFZ3H
QOF+0QwurNUlV7Ymr2GMpN9CCBZqahlPQ+LeDxutHHfZdP3WtbD61H7S3aeVSrIlqrwewj9mJfBh
07q3UhiQKP47IsPwZVWZEalzVRG8jOqKO3DTew5CdelArJ9fltoBw7B0o3Sbf8mtwINdiOlUr4nc
9xMQPcV2F+HJbpxYDdCyy8Kz2uJ5ewIOnprFQeljnIqQrUO4ntuCGIsHA/NKxHr7Wwn3EgtbuDJW
lmpjiftUMPnYbr0jP5a3+FOQw4VTLkGOiFmUq82iaqBQ1DKVXA7aMvwPMu5cxinrzIcHEn6cENBY
/kPWogJ0w0ztwZnkwLE6kuAMKmd3H4hLz8HOq7EwEZJ5+987+1K0cCFrFMGQhlf199cvsu0IjAXz
fMayHvC6S/DmrR8oG/mdc7rOs6sk+V0eI2uKZKpeR7ls6ZPgo2gTDB+hbOBMdcT3AEUa0hFq64u6
hBIyGFBT56MisFB+cqXcRfSd3OM3Y3SiGKXqEOmq6Y6KcRBVhCQkr4uHaefeL6oBidtxCZu2tAsh
PcW2R8JT+oSei47bnWuKfyW2kwfKYP3EN7fZNWLYNbAgDpmhIr32BxCakDcPol/Eaj61HIgQtTdi
NC7tqMWRhAMvPzB68nG5kYTzBoF5WGKSN/ha0LnwJKTJiARmJTfrHcFSp1kouO4gGwQkI8ibSe0g
FRDrY20qh2PxmPOoRrfd00UcgcUL+chPZQuoLzpUsWcJv+SqFwmmSo7eq6G+LeLfgibf/MBHk0bf
IiqeMaUFXevFkrznsU/Zn3zadj0j9BoZjzGWb2z0eez7A4DltDVFSKsS4T/Aq/V+sCo9cPCJQhHw
fvrgr+sBxYMoLVe+Y5s9IUvhWPdjxPoaOTuEJTz+7Iv95C3oxWgbtUBPWPUsQ84Y5vEO68TMbu71
PY6XkPIRyUOvB2PwdMbqUT/Lv2p2a6yu/h3TLrtC6UlruzUuWPVu/+oQjJpD4WAIMxrHzIh8yqwc
umICvs12AnhHikcRThvWLA2D6+92jLJqKqqUPFaA7yG+AU09D4mFclFGz/NdPBsyB5/NnVX1+SHN
ttrquJSykrWs+//sFVBE4T3lcXo3yhU/THrWLJgc9k4OqLAQ1vmHwm9LqnZVy20Bvn74hKkd4xHV
OHCmOLYdsH4QLlHeYqmIwimThG5Gjbm1w4rNXed9HmIzfxPOn6FL2d9F9PW/RHilop5ETLUjuNgT
EjIsACFMuX8rBxhZVeo/hTC1RwESm0KQ2Xjq5gsGDxXieEhSsUk/6+OzmV9lj48AbTUwj0PEiHqt
JiyjYP0tA823hHzVsILsjjFUTZZ0L7XEgQXoai/eOKD0+rKrILYmppnel2CcSdSnzD5q6tgEemLm
npBxNCfievbzchwUO2Wtwpl3cdrLfVl/7W/X+Twgt/ISDPmZwlt4ogZS6orlHxBvMF2vKtK0GAxT
Ay697blxUpBMuGtxFx8Cc+Jqo9aJdNX9dcynkxKjuScqGlVlFh1j9y5qXGAU1/oEP0PrAet4+VOj
aqA/BKbujLYo7IWDotEL+V8TcVt1ICPNesM2w5LIo3AVqXYZ51t3bV6uQ5zJg4tCUtGksX4Uoy8m
iJXixiXNTmbiEdhkx0CUcIIalFONvQtlOH0Viy1CXkhgK9+6eUPTGMbJsRdPzJ+UiQVIVU2xRVjJ
Fl4W5PDQIhoe1C/F8665xkELYazCQIinHev8N5K5f2MKuZAWU0FEXgggPw+TCQqYeW5w93/vqdC6
esPEJExy5tH8kb8RZGnVzenNpEY4Mn94o7dGOjqxytodXWm2c7fZ9Ot7qdBwC+L6LeXoaZGo8PQR
sD+Y8J0A/XGc/gpdMPc1oeRvG28bs7AOGptg+Sgvz/1lZNDATHbDuSt1aHx2PLdSz7CktdSqftI7
96v9++moLLOK44jhESR/AdcS9LAP1M0va+RG7xsLwv0z7vNRcJzJMjaCRaE46s+QYTOd+WwwobTf
B0VylFkf11RZS5yw924tPfKPwDfgWSgd5/Izv03bbdeE47Rrgg7xKRljjljpfO4MjH4H8yeMySkw
QdWm7wV1U54BdfsL5ATFt6rbquqMzks2t0GmS521MTid7EWyl3WpDsK9WT+iLDZS9PkvG1Tx6SJo
N0A/tsSmEVRxYOZ1zrqOeva8OJHTqYQQoguHYRc86qGmwnX4CF0tRf2rEAu/lhKZHnnHIigfYHYI
sCdFCeK+gookW8ziukiCfh7JCuBiJuPxErJqyT1FvJ17UQ+WcXIdvK9/PMReq0JpIco/kiq3Ig2t
5rlTPocnufgT2Gu+u5WloUMjFKXdYjErUxoQCkzMpahD9h03JACjbtYBnDUOow2R8obgVqmB7D5w
rR3HBw4suYmAvm0/q9h1YwTVJBgohLJCyZRza4eEof9SjVGWlCJovqFQHMBZbjsP8tVaWez9jOBE
VvNKCWxz8MX8Cu+bFeKftbMZRtGEEBBQb6tx/QKnzWJEcGx64UeFexLPwnyIdCQEt2NcBMC1k1zV
5xfX908yxBHNrzemXF2RDcZ3UuFZXrRbcmKFCaKTUm1G+zIEP5j98Gjgn/f7GATm967XjO1wYnwI
P1MjNjheTcgqZjow7Ja2Jk3CJL76DqU3brRYIE+2ndO2hqzH6watknF3WAresGnoR+tmO/5S9olT
RV1BVFYLF86HBAsSI/tM0tJVpGZiIXNaMVoj9AlITcc9KdhSNq+SHccNVLTdhQE2l1vXHoaSZZ3m
jmZor/e0LNqOOc8g/OIHtPBss0ZNrvx7l/9rzPqL3APbnUwseECudOBpDkMjk6xEQPdhoo0XfXZt
QJSwSEi8WqFCKBW6ysJ8OnK1HSfvfwgOAWc2asEOkY0aEnMmTwVIFBw4GONbMnJU1xHhJphZRQc5
geL4Gky0sULhNLhpFy7DbQOe++rFBieyibivh8RhvTmm5EUNwMAPDRiumxhvtPcuRjDiYDGsSwcm
plOGEdoApruxvD+6MEpeHwBuOy5QhoeQSAT4Rjo86JMsHeWZkleptghn6kzou17KVCPop6zQhYjo
Ii6R1SdoMnGuaRxbKrSf/xTJg5hvbmTm5F95tLVJKq5CFkCdhCyKIaJkBwxX19Ehzw6kl1zvlFx2
qvZuN8guYyVCOEDaW79FXq1zoZIyGUz1dAUBxbb+kKb9PMbnVzHXDpxpo8/GXh/jbLfYaw3cKtiz
I1iuncftJfVHErJLBhbl5Ie6pcDAymq+tmKLwFdLI72pe+5UWvS/wh3udGiSo5XM5fNeI0/N/ohp
No3e5iLEk+hf1qR85UXDPE+j9MGZykX7vty8LIPKcU/ozeb7pz2JUneoxf4U8Y5sXZlh6uX/rKhu
tX7IW2lHwpZ6nYi/2bu2/CN/FTcnwYoHytyil/U6ElP4RTfTJ7aJDEtk8spoufKe1jyAhY5eTLd8
3MdQsTb3HvIWy08+WzaRTb2uPU957OhQNEmgv+I6Io8k+RBNbDGZ5AeJIzL6Vvv1WfsVZHlzHto3
Y6Em5hvbLPaJfNrrRqAdNlMOH+T7KeixbV2Pk/uPO3z4rTLOJ+Xw6JXnfTbGNo/zLGnwOaWBOZ0T
xHCRA5EujD8HeI5VYhPkFoWqKvFJUERxxMFlTM1QZVosb/daQ2cpbz3RP4eQU3MuSk+EzhyZ7uWt
mo3rGPfYXGdj5NAMnNoFRD+bdV76zR2Hbrf5G9PmK7BiHiPHLPjI7jNLCE4HvdPbGRLyXac9voFv
shPtyEMHaZZxOYXqw9TjdFdgiEpfRW7ByJgCmg00qLet4lVOVYJdpir4UTmf7I1qRi4ZFBriikWA
RJh5weKtncLmgaKStxkMB7geY4s6XVda0MFKoGefdUU+QOAzsrG3eQUDE4utVkBfnAlm4N0EDJL1
lFvsrb8IyjDlUIaimA1vvsYCJtOyjVwAx3p5SCCS0hDTTLZKHoNUUsHQqBOPOQmXUMutTn7qMgOG
LWBE4Kv7D0D6Gh3fnkUTgzhsFMKyrHSusY50GbxvqMuP/ZtksimaOm5xNAdsg5C2CdFYzSXkIH+l
Qcsc+O8S8P07njrPlEV1NOzPKMaD8Lcg1FiVW50oqbg007L9FCMYUxqVKMOIOs+ZjsgE0AwVLx4f
qPMU4PSIEBaB8xXogGIyuX3/YBA9AscWL02O644rMF8cT0Dfk5/jf6RJw2NE8e3KyqsETUX0Gp4w
+fdi4sKsha81RLfxlv9EgaOSaBli6ucnbKOiuEe/ERo3CDvr2fD7kGiYSr5svfxMhZyru1y0Ghks
W4KUy077zgW9BN0uJ54eR4xJU79nJcu0hxMXHDvHu5OefgPdQ+49WO+pS7hK5G9l+gCP2tejQzhs
PQeWkXyKyNIvkgzuYV0GPxclxbIX7j+gqCFfdz6OTa21MLfKVU77uBUqbAQJj/G8FZvvDgH8pnmn
G+s8Y+w4o71kJf+Dw6gmLFKSxAGzapia08AHt9fKhLswhwFZkqPCgKGfEpOxpl3/RTOGb/Oqz4A4
sjHTuvJbi/q8+bm7n+yGcKvW4tcGK/lIE80ty2xrCXhGxPQqfvBZFlAjB/zvJonZ/jEkCV7J83za
JGlx4j2hFWg8ic0e1h2Y2Z0U3ZOMuZi+T7zVwELEs3O3s0nARstPtLiM0ZO5VhFZZXrSmvlXP0+1
KU8pN726M3lZH2XjgpxjtvDXPdItAJQ4vp5O9m5js0p0MgQjJI0dLHwnUI72HiJkRecX7juDeKDz
rL+AyWsMQ7ZvQvHs+bdE1Zv8Aha/ewRdjUfoNBhn9h2WM6BCwd+sWpjlrsNgdFentrx25pWDA9tB
UJF4PAZnGevpwnEqh6WBxT8WgyrVQjJH2fAepKZeLM11z+pW+J3MRNQlfSgx7i251gBAX/lz2aGb
BDN9wKTiK4e1zWTPcVHEoYr4kNFLHGftvfz8veITnTHGhZslcFwjVs3RwB9YTfhJuK4YOix3FeHN
+VXf4GTaVpZIghQBFRRsCn6uwcwfOgSec3HRH1RrVXDkGSNXX+IktCK6dgGFHTZxau1Q56vrB4bV
356mBlQCsJJdXs+6QAM0q7wt5YIyHgXhNF/H68H/Sd+XMQjrS9XxIKgEHPC7k31J3AJKYy5Ahc+O
Nf9D6DbBHkMOZocEoMKA0jgLWCJKhjcz9f/+/IlqYZN0gwF2K1k59qWK8t8Ics92SWsE3FCo34DO
2Yv8PEjxnbJQok00X/OCamqH67dx7iSVDzJJSisDQBfpnFizE1OLgfWGFdT8BDgxNvwaviBXykzF
eQRk3mZzCVc5zqpv5oaUlU3iLGUGFM5WWxMCH1v0ze2rVOBAqK5fbjLvTG1DArfruORoPYy0Mql5
2ZMGigBJ45rD7Scqfy7+BK7bLriOstV6rS3aEYx3K7unvASHSQ/rp9epW3UfbqBXtSj3zMUNh+xt
AaC1Eoq/vFKtU3y39k9L//SRt5JC04MCICDq/7YdoxJE8cfexROF8fKAQXxdKnJ2yCbYVmzX1NFE
qMO8qgyEsRKNO2aEuVm1G7rlfCtOK8mc1N55uRZBUi/rFs8jAeITKH5/nNxZT1h04h00lpvItbex
Hyqsrlwb3QMHlgouRbfcNbj37bstkMEHoAsY2Twl1GawvCNudPtZ3O755UWRkUNtdDlIPFO/V40P
980EUWcFN4d4LrIzCAweSGyU+XbxuCA9d/rYKaX7N/q2u5cGHAMLVdbKKb3GgZQMEUTqDxwdLzZ2
skrZiasQ3E/McVorCD9tvZ0h4Qo/QqjCG45juwLKuXeq6LQ12qwFt7io+oH0PZgID28zjS9QcMoK
FmSBjEvkyi4vdD8N7m2IEYbiF6rmScoW3DXlMhHr2YNAUTWDVmGAVlerN/TA8yIcapRaWlmsjqqh
NCm6K3IFruEMtxDB43g5O+vH1M/30NJ0e3bXOuYb7s6S1K69hSoAbA+3xW6mBCoeEsUI93UI0mrD
b4RcPDe/lA4YH6y//sLmNZhjFNT2UVRTvCCROHwAn1GkOfUAYt3cDyyWi+IOgdZtuZBShJvKVRQ+
v/9in4gWiNV4ye5/177z/Xc6FE0rjhbIXehed44ZKewYPAIT4bdmrWWD1r4Wxa8z6cv7QZeb8mlx
S43mCo357G3ANJ5TjH1/gPJFY9ynF7/5afBu/BU9xU7jGalp7CbQZxUBwLeaczM6r3Q/5Y2L44p0
XUHMhjsz2ukf345u0yQ/AiqOaanTFgpL/Hve5Sv8zqQcPXI/4IXu0EoU/iTykjUNTVP10y8qHPXK
vVSPMZVYoAPMKEtANq/9Vsw7H0bRBQILMbhCrVCmzsGeXPOt73Kw/1aTQdjbaBcVtobsPPmp9Tpq
bx0YR8qBcUEnPfVnr3mqZBbcouL03RDH8509EST7fTnVXf/9xl/EsgSsrwUnXkK2GEupBbTwaJ4s
a/rG0ULqYSTSv9cbGXDjsZaMic6cY4jCzS8/ge9+Z1m1GcWVp47yPkCkcbirLaIKovQUJ02b/d/K
greCtjQFsVRop3/+4AmAdY9QhRBmiPuKAUTuYhZFrn0haAa+lqIhqnq2R/qroj2hHV587eQ+4PSm
1ByENDb8qLVTw+Y6ZEKV1j5ISjdE7ygD2kFYYXd/NISq7lV9nRlSzCWgEVjrMw94GZnbCn5k//Uh
lWh0k3gtpUbawGkReSZ01mw9p3OQJlO+sZS0YYfJxaJqyESzzUIumf4E5sSHR3nKBWSZfCxtyGpr
oK3sueR07AU8Q81BEFN+NGXCL6V0CwpIhFIqR5giPL3XBrIKmvi11Ab36JAEbQz726avNk+KccCy
octDQbunERe567NDwxPNjU9acZ/1m6AsjJ8BptrPzaMAbSbkiSKriWeygq+o8WkSVyCYEA5hmR/r
UJuaGje3eQDV1B5Pt8NBzJ2OFypwlWzpgid3dzQFjEjM+5GxKVAVVgz/j51Gv7AiA7B4es5rVEJR
SJ/6YUs9UDi/qwGDnoGZbYyH1nXJDYfgnpt7C3l+FAMwbR9R/j+ONH55Iq054xK1A1vrTQPo7yuW
WX401R/Er1xJYaPUJurChewvBParRFPq58nbufut+dAlcLeqWdM2YsHpKEt0ZOzhUY+FLEIauvW/
fgQDmXieAHI0Mf+d6nZm1dPMkU7hsfv2QTv+ABTHlW6395XrZr/WhCufXf3I5zLa51s78rvipCAw
LRjpDfDoom9UG/Z8QuHpnJwz2BETqfnRrCHzf2oOXuDYvnlovTSVJnjf4iLdydeHORnArrccBI5M
BL04nW+X9Hknr40QaVor6qwJvPxek7xwZwhf5GD5yZejokE97TSELTZKSMK2S4jI9pfcbae/KyC5
Jeao/DTcYzw86v0j2952m4KLX10NlcFR25jXiFx0hp2RS45m5am7xHRaNkleIGdNo7RNe1dyEI+w
IrB3GcfQ1N4dz3Ccn/S11Dv0VOw07kyamzpKI0lAa/pPy7i2gevwX23Oy3R2AMFK7rG0V50E7aDk
iQouNbWgU7mMcoOJ8VVEWdqNVpNTpfa7j8WlI3AZDl6n2zFhns1Jf62uYEJa7L2yANWt7Wn9SzB3
zYM9cxqEu1jxy1r3fnhspDWmOMQ3QGAVzG0XL8V3TKOar5ie7u7O8PJ8RnG2LhnYpFVJwT9rdftP
/XILvngIR6Sg0rSqNp/YWpJfuWlyLIOiKTlsRr9jfmacrwiluuIob3VrBP1XsTwIQVJ0hQTVCJKr
aJiFOXdqGNDUW2Je9zX2JRETAf5nxN2b3fMFFARONt3AIAqFuxqxrrJK/rkSgzi7Xp9pBqj+DBpH
wm150RE4LGTtv0hgR9RNY3BS4R6yGghexrT6fLw1sp0V7/JeMWBLXVryX3iEUdjCQS2UNJyf510P
sHLBzZszNVrV+woFhsuvqC1SdsC2MaSxlGnZsRJSXUEt2RhThZKpKQuPWFzBJp+gXLpgvVdo6dhu
C7JQ4x4JMQ3RXE6PD5egGWtgHs2CS816b3Dqt+eCRcghgdimJrN7UkNJFlsWIoEG1c0j/seqv2sa
JsCDxrzgCeCo8abJZmazbkwivknbIFOg1RknD10BdL2Modk0Ss0JswlEjNbo3imA9egSjGgOa3xX
78mdqOQlNlJqKDP4sH8secFpsDGpGhANqx0LZB9/H6FJKa9gfLHvpMYYzX2q+Ww6wjBLAnxVT6BN
n/RMpAyd1jANHmJh4VWniLxVmdr88xd0lRIbinkPFdxvlLcOykkqx/BiDYEtqwHlPWxVloOS8i3H
U/NxiCn4V52VWE1AV/ZHqCraQeMnqpyWAvGSfvo+Ruo69kJbHkmKBrhA8SDzFuTfHCrOjzRyPVdz
U4yo+xFH0jcC/fv/kZg1sRgNAB4K9wYndEiARQQM0+EvBnc4GFUJfTqb38xY67TwkqxPT2DAM27W
oKGFkSWaQ90JmlxcB3/HRcwDOW9zxPxbV/D2ttT9Ijavi1s7V0UCtaP78ypm6FHhEIFUJwTmd6mb
4BgBj1IKBptU1RZcsGFAAvNktJ7vRIULCWYVeQykK/THkT3k8II8CXj/ohZ+Og6BFTj48xsH3LAE
Oq6+IWT1euMLSysUcdWVmYQhKj/pmAY/PMYljsnr8Q7ty+RlzBMq9Q8OzafXdfbRYP5ihvDdqNir
QManWLMO9U8iTy6twuGANX/LuXOR4M7kdMsd8q1GLfCFhGj7hVZ+N3QgTYAM6l/uB/O1Ppfc01wi
E6gfO/swg8l8aFTJ8J5Y+i2QtwtCSU8xKMHg89Zb0oTJ38ZimuVFHMpt3HOszVeDhK9HDm8yTfp0
Fyr++wmewBEgkL9x1TJmqTrWKbNVdI8QpplVZ/x9Jm581l7n0AH6LYWtiFi6GFlNB5vrUMsVOpSQ
NwU4pm0xe4yM/6jCdbE7ZJMUPO7CiCXTc4CxCD4S7GhGNa/qz0ZuJo2i1KsmPXC9Ign2sM5bz0Rm
mlSWx7Mf6sY9G+Ic+K8/2khyyxEn91xpVbruwWLBOTQRN8NyNhYTBuAf+Ya6AFzlh10dNd7CvO6R
jUR0w7i4CWuehfzsL0fOgHCeELSskvCKQ9HDlpmmo7Vgz6PW9h1fd4D81SFQhApmkFrK9nim4e+F
+sUamMHD43Gn98L7DvI/yhKuhs4C3bBrGdUaoxkD8XBQc0YGA7Fvyx64z2zR/NYQoRVHMoM5FqAp
5aV33ZM1pW7uOG9i7rs6LXh6k/C7aP1hQG9DJSMmZVvyeNWs9FnQER2kuSrOSiAgd2ILuiNRAfFz
EFIj1tOFqMCDv6e+5p8cr+strwt+MiEVzYOFlc1ahdTPQRPnv0iRXMHc8+S3orbv1qHbXRIEsHFg
R0w0BSEF+XZDR7A8Tn2c0vShxtk8zSEeCpWhFM0ZB+jQyFeFoF6cNXHeK3xxssyOhLRMLztvL+cc
so1mqLpm6TnuB84piNex4kpnLnqZpzEowDaVbRqwMjnr0VyuFKGDVULqauHmgkfGtbZr1sVmPeFs
+JxM5QcgcHEd6jtF24WIvfsOWgW/eXeKdh/3Cc5u4iSJVrCgo4MVMAGeAVmAneOEbVgBwHuoipga
6otNLTb57lKuqb0pduhKRKBg8Hj1LXLdCNiNHVtu42nqZGwaH/i4o4mtM0iJ4qLqxjnFITdSeJ/D
FTfLDTuHulwqGkmYxFo3GtESReRHHE0suCdSfna6K1XbmH71kOg8DdxofFsDXo37RhWU3ctdYa+l
IWENA+LdqnK07igjoplgXuIi+Wg6Ne/mnOmpI4JBHHb2dMEbxqiPAolGBpNJED18UoxJH1A2qNWO
sHc36YAxVmMzB8qIl3grwlsSYAkRN+uCvCzoiJYuHUkxsQKnFFXgd+0hBlA41h4uUA8FVSe0D80g
VQdijbM6qQ+iuGUuEL2n5tc2B0dyoVSOqeIywGZOg9Z2pHNlbL58v1C+V1eEUF/tbHO+1v71YtkE
W9I5ZaNBE2yOZ8MUJTrLBJsZnj/dVmc3b45YLaP0joPXDWmBS4vKrum013c4whgprNe+NZ5Sev8d
pLGWDm+pysaNCg0RcIjHK0Idd/p4uS3+t9hK9xTGexFZ/lxi5h1OdlIyRWdeEqPHGPO36k5iwJ12
lnf6jlK1zyzt/O9QG4yrNlYFZjX9lPBA0J8AlHs6I7/X0i0Qhp0O5mlkT+0sNcsccFF74PN/VeZ7
RCbzWdHTvqdDeLGzDwBb2LEvZWGBOhkQDR/Zz4Hx4QvJ3uqAYZkrOY8kJb91FD9OrYiB/eIh5AnD
oCkAuL8RVUcyUAtn9srTZP5KKwy7X2BgcFCMxFqriUKp2CgAGvjXcCqQNw5j3RsqRXbQqRnHqL+r
sV8rZwNrztR1LzXbs03XtoQAUQgIsrWLsXeCOWIY82Gs9fq9S7s8GsNPX2WE1NAVcIlAKngzeT72
lG/b1+jYNWSDtKOqlRA98dL2059/ZiUUljrOjthIdtWXCNCeW4rfhshy4co8gARY489b+EwjlC8M
50t1D8rlODqHD4v21RybhDyERJE04YkiWszUfFLauaPYRUTGuSZ9GfZmYqio+THeq+r8sJjmVcvn
ADzFbqtFHQsxDFKI9rnX9+bKUCchuGL8cr04/T2+iQVekg7MTCut9rot96woENqlVGqAwLiLEkAC
lP2eJDwVSULYaHlR83Sb17jRUfVmSXTn44WKuWpCsNFUlWom2Ja4BIWyFHpKkCE3cEdDuH3cH6Jk
XZgmVbp36jZ25e/zlbE5n3iS2d+t1pqRSPHtYdnV+aez9U2sM+pi2/VfN7yifNm/+3PIlSjYaAl3
nJ9m/DtytIbRyQooTon0J9Y5/bKHTNfmenaTvrnXoCeCQ7tVdY45WE3yb3o1aczhDG0E+DpHH5N8
Jv54N9Dk5UVEBIj4ZQlh2fIp4ucvWe+HbPbrxmYZnpxfsYQzSMSPvTOaO8upcA0bMgUVrPUT7Smp
XYER9Iu5wSg3UrG0LYSDhVPxmAYsbBu6PKYRQ5JaNwPEviaqEYwixHu8xn/akpVrB6EUK4SopaZQ
bN9kR8EZDl/TTzO9vGVBHKhSVirMJZlAsflTmZahF0nQTsbh/Vwf4gPXGvoi4sj2xu3IzS86JYHh
dZ+19P2nGq6cLrDhcmGTknDhiNRPpzxwp4H2XLL3re8Ea8cdrev7C7gazrye8RTguBzr93XMzW8T
1Gd0qyM8VUIPFcXVTBd/jcrMxMgbTu4vx0NiJHiYUjtQ0UhZDjqpsVM3gdoFnmoBG/q+qSrxiTUe
dqlp2qDBPDszW77gK3l/VAKrCy3tzDv46Vz/KygIJksl29HsCGIRUQ18II1ua/sCGkjA1v0HT8Yr
ivrOiVV1TiwAgEQC23Rmc1egG2u8q3hdVGIu0kuH8wf9nR2NTEENRkbYNQv7QzUVo+Ym7ca6JnLm
ycFDwzsup43Lu3RmtrSVNUD/VLw9yxnfsjdlnSAhJDTElPy6c/sALfqCN6C4WBX8vCeB5C0/jdqO
GzV7B8695qDzsmMnp9PUgJfTNhCtazyUtR9CPK0z70RebgXXRSjvF8t7b4f7GC04mc6OxZ6kSKPf
lNlGDl7xJaxwOctEp8a3WBzPhf+Y4XzgHJ2vwx09h0aaLb8PfQM2SjubMvhYVpx++9bJwtddripn
kV/OPvyQaZgTIhJuKh8fdzOURKu7vfjcSjUSuPxlbtoSTYVOq43o5AlPDBaJ1VotH4uHP1tEtMer
RZebAhuB3kFwhyQbPx4ReftpdT3kjhk+OughRi81jrzPAKJrLJ7fAwiEKJ0s0XU83N5qO95WZ1U2
LI7Gv3q5nbFZyPGJ0YfUDg/FEtAOcDdPKUPqBupqXIz+BTmp049IYB2zg5kBto+jJVqGMRBJHLCj
l0Xy/7IZCBQhPR9UbBH1AvP5YrfBstrstXiudDDLlH3TVNaOerDzuazpK1liVd7AcpaNnEuJWZjj
99m8ccBbPKjw/Int3SnA4mAkMlmkJcgIFFitVJj/izoMCJHOljmcOC5n6V6/gt3tCdpJB73ssyEy
4dM2OF8hGWeTOPr2odLdsX6KUdQ/y8kcssJFqZ2UkgXorr+XrFosndFUrhP2Y56LQ7K21t1Qft7e
4XBAz4nCc+/HJz/l8R9Ogye2uZpCoIAIbQ7pozO1zAAUEVJxo/KPQB8H1fNCEkR9ExxN1PJVSejT
iaQROjdrgIEoHdKCd9PuCFre/v0kKbG+2dmPH/A4DVunOtUmiwIkUmKMHD/vY5dxYG6QbnSXVPdd
Un3GakKBGmmqmRpib334F+zeFE1s/DJesMI7HdgTDwOEo670gL/39lha5FWTAhSf89vNnBHENYwR
fMxr5PreVQkOm5/qE3N2AtId38SQqftFklIsPp71FRP4a39GnYvEa5b3jKpFgXbo5NVgHjlgqmao
3IQK4nGTQ2I5PMjyUlyZ7Z02QBQ5TZ7kWTS65SoCZGCkDip3k6hp0JxVtFLVEkOQSDTwm9gXgJWK
gWuIAdPip2ScEk6FZrCDDQBblO0SAiRWwM1BsrK91euzwvxJ2e6lzdJ3dFQIujpWnrJon12ubsmP
hG9z4cbcqVH3NnjV/q1WhQCp412sMTEfA2b/Hb1KVZdLtx/wolF355kp9QuppehFVF/qQrR8Ghlr
Be4jyV4vZ2y8rI+o+KbvHJ8j5LnYYlsPfUDECKrsm7ylEkM494qi9JNSO8kb7A33bD7opXXHA8h+
gl6BG10BPjxsACXiuUFXpaWDHHggvMp5XVVli4GTsa8zXjRIFBbLrg+GuANBSiOMFPcLwasDM455
6YzFYwKL0tNGESFwtHyfIuWj8/yK+0B3ByhPuUF79HNrsrQo54QWfDPTuefih/RcUuyhqL0O49kW
GHqnExD+AVbWA3wVMC7fcKBk47BwBYiRo7O3b6Npqd3UvJcIXr3+mu+4pOXA8OXlacaJjM0fsJtK
Elkwqef0dxM8hbw9ctcNfHSx3DoeTjGrZJCnCVcbYdYDl6/p5zdMUt07bPE8pC+AExgWNBjhzkUy
FJt47UyfRPXZqR07PaniEdU/YwPw3oeAMwyl5sub4buAsiIjaYLnt+4DMvvlcPXJ/gwY66cV2F3B
QVDkUWSuFNl45BQQ8NL6yavF/C4ucE9LDGReydBAUQZTScRnopORnfAn5PjiWBdP7pDZzyfFPC3t
jyqp4waM3Xam17qI3+qldC2mZTmzUhzZRi/1BlNBDUHIsiP1bM5WwGIM+I8ipv8bWf5r2AXDls3v
g/rblGjpxVz6t5OT8W8qEW7SNcyZ3fvOnW16pTzWBEH0g9S/3XQf4t1VEf8FlE2LvBcG+acIwh9K
mh1nmb+Qs8CnX3V6qXsBYnQ88FeNTSV5MZgc8RIfkyZi12yU/o487K3jkpNH/mZKrXWJhM7ibqv7
aGU9N5d4AZ7Y3uyvsT9sYKUeUQvxRpTxJOh9qVjjE7vOoyILgnzE7ZnWfQFUWU2W+JA1kfv2ZOHk
o1fly0oQq8JAZFYCmdTzh3Otn/N62bcI7zvU2QP8ne/8ZB5CYFCGnhQhVX7OUsRpkiby2fCRWYcT
xjAFAzHxHHGUT0gDjtK1xp3cwTBdtIZXQuuiLvJkKvqifD/0fZJhC0nnewNXr4KxuUMLpTK9ptgc
gr3nzKuOqHXFSOrMSTZvkidF18/x3bG/BC2HRIt5EYlbmxQja4TlvcpBpl9UALCPHKGIz9gAND4/
V4CmXAgAw0Ldv19iAVepPDBp5zEBS2NtFJgkc+WLY2nUmejpDgOEHp0nhhWdcjhq8sxz12tgYzkc
yKSbZuPk5jfQ2M/QdN1xGrn8n6CN2aYPyIXX+MWnKqwrr0W+YqwoGv+Bj7+6OM+jj+e+7p+dfaNp
rG/QSDsQ9m9oB3jr2zVoMYuZj8yU1MG8xfciyqdWVfch+gIDezOM039Tfbi+nSsAt6NfVn+TKpgD
IAdOiKRV4GDT+whBY879tUdFUkoC5O1GzctCTv9wrE8Opue5Ks0xO9XIQlWFzfjkr5aR8/jJxM1Q
o0IyHoF3IjrVkFxcsJYriqVAT/99XEJg/c7RuYDMT+EzqKuP1tmtW5Oo3cYucIQYdN9BiWTKZwjP
0xik8VXG9jwb7hNAcEZ5KVDOKB+0nKSSrjbSOQolDfI6bS70y/hyq8oEsodMfT9GoAjyimRrzGJy
AiiK8vyhmLtzdXVHQKI+M3TbNrKaV78fLUCoElbFyoyu+/94cLA8Div5j1uC/cOucILVIk6+dmIS
BKcBU1PYzoS2peofPwsI5AOk6BNdsA214C3WW5Ru3rGkSkE+KEnNbdLfhoysXwd5R9rrLegXYmWX
d7VD4IF1iFDor+BbQxm5fO6+jtcc9kxapclxe7Ctblfn9LIlRidHa51H0Fl8Ykg47lysxZi/WBVt
hA6KVsDY5NEUoYB++v1dLJIX4qdkQRGdNg/3mk3dELz4bKF/WBFelI0UiD4657EGn+y1JhX5WcPC
eVyEjkktLbvqc3QFrSxMeUO21pND1eAhACyvT5/R9sMrzGUCe5tbLMbmjyHZpzi0L9ikXgVXXNDp
3kJTCLDBjUdKtuw5hz1bt62kYMfvtb6C20XIiGAaBGwKDDuxQEdpBp/P+OGVAjBtQWg7kjbHuhfM
KwxZtCj/AXwCJktq9BOqGemogk26iLY0ICbzw/ZeAX8tZm8LiYgeuCKgwkcYNBuWg0l5dF7M3q1u
MjTAxDZLN31s3w7jVpgdVgaMn+mpY1+WHGFNbWwCjKUcnH2RL5CVdlGId1KqK5ccsvWETkStmAH4
TWvG/7htcSPBJJ2x5WSzDiveYroWdcrHH61faWc9tn3Y3BsezV80jWyGs3EQOyhK459wo/Dp3/Jy
Aw7WwIdCHShf0NgdeIT8ZmTPKbHpXudV0Gjm87lJrbX2fjj9vTL7lFRiudI7MuOIejNev/zl25SL
OYI3GzS3SuRqLqTqkkm2sY/YOrKiftGxEgM+cP3FSXxcrx730Em8PipTpL4ztffZ3rt8zuamB+Z4
4hb/h3y+eAhBz1qDmpRGvUbZiEXQUqzDS9TIbNiSbYMShJptdhRf6xZ9h3T8rOY251IwN/Vde3Hb
rr0bDVWo77nDqU83wmf34pLO60vBkA5+kgVTyYksgxli2EBVvIgbv5aug+toqiicB1Y82ikcBmlc
mC7TBjTeqis18/MriwmnNDl4Eg5yMu0D1TAcTxK/ICdc8n6+Yn7DQiyeXYN5VRGXGbSnvg3FqVlA
kKO3sjiL4vZYAdwUZvzvoIq1YpxerS9/V3a2f6sZ2MP8z5kK6dAVLPHnipJTjAZGKAg3EhTX6fl8
pj1Z0ZzbETHMMJp3g+c52DoWfZy906lk/Q04bklrpMjG/k9AkWqsZHjBG+Siqz8ctOeSR1oSx0GD
1vyj24S8XdDRuxtWr7IL0DcUpteWof2pvo5Hw2Q36yfPufcW7hASBJu2U+RRG1KbCyn+J5/2CWnt
2RJHubMFABDzoQJATeEFgy7UaA4bZL4fyrNXZpcltJuRWOJLtbhv5MWcy77WWaOjaddaX/JmnkQB
hK/0AJAVV5evLtgWifTn3BqP+GYNqJKIP+0YZsZUydCa8wenciUT1UsP1iWkvPdh896o+mjiztlV
xFHEvJa4q69Tgf3atvNch/xKRhvO5nnbvJ1u/J1hcSxjeqrS8bYuhTgTFI5jsITvXJMCwmIQJV3l
m2dveWEfyLg3mRkR1xjE91UPjlTq5aBCNUZhoQzvIlkYq0rYoriAzt5hk6rjDG21V8oCRhZLvKmU
FADxbMO92axKtID8gGPkWZ3sr3AnOea+f9fu7GaxgEH6dyGzO01KxX5r5dEwu3Qv6wPzn0UCjoNJ
9nbS3NYsr3l2y7Rz/705v185yr/09cADEqOhY0GnefqammRaxQViffs+PhyFtiSULTxc1MFtpV1j
UjSN3mzQeXEEOzm256/2vnc93PqZ/cBitxW2svLvyO5EAVQW4U5LeXcLyQhL7KSQkWAiqd1N/lsp
MuQSVlw+cu6OErna9we3vDbclwZciGZoxRqvh6KEdwotW7T4BSqdwWSA6NVI6b8QEfQFrTLKmB1h
zuP7Hh3174YCDZa06U73BUaZPdcqjKQkRP+ifVu7QirO7yvbB/r/oCXntUHZN0F7DL2BZ26ORE3I
QIG9VEz4bTljSZ5uVTGSwb6fyta72iVC2Bw3nqql2ouNQA6hwnKHarVvGNNVmJzBCmJ9tpXYQNkl
WCsjpupT5uAwBGuLkoMCQwBaZJMhJ5g/DQ40uirxmOnLwolWyeIgGudbxlScGMmM4mj4h4PuwVhX
iUAkEHEGZ2N/VKX1GrulS9UrVZs1Cn7CvcFo+rg/BfBTtMRmrhu2P+Z75wipj2TMzKcqDORRc/19
Ud21wshjv1CbTiivz2pPO2elRlRiGKeuRMO7nFOH9PYsOMSHIPAV3yp7oSbnEUhx5lyXLmQ9fECd
OknStyKEjK08ompFdzEd8mcoT7pkEJHooo2BUuPxnk4YZQfXkbqy1GQR1sp9bOrbiHL7yPzsQAau
bB0AvTDy3/9Bwo28GbxlJSAAk82DXdj+E2fI/I40StNNmHwFZoNf4+17hUL4u8hQIFkiAZUrjH33
7UVstssyX9GHg2BQ1Oh0YnImFr7NTbFlavdtBixcpg+Vqh3Htr/vQ65w0epKNMBQFPTvdo9SJdyA
hoB5a//a4D1gE9ZYDKTpj4Bv1lXsKuzQ7r8RmOQ1+6qqJNxUc9SDH7HdXX/NPaXVY3asdjgTlnxO
Ppt8dOlopeWDJoLjj+sCdBGnY2FIcfxIJYkPDsn85tdYottA5p9LxGEK8HB56O0sXFdI3w/E7yJ3
S/kqN/Ggw5eiTTv54F68Zs5zyQrYs+/kN19tcq7J1hyFzZuINX69lt0T9zF9jgCStQwe6hBp5fTV
XcQ8nXXib1IQrHfEFBf9DPWVzi7b71l6uXl8Yk2ivq/lz5DAMLn8boSerKWXPc+kI9AD69NUnMpS
m+TWis/bwvQcY9fJ4HeqLKsjdW4sy4iLT0eTimBtCTethmp9688zblr1Sp9zhoeUzqEKMT3IwrHG
TobABu1xRwzs4oY+UI8CzNT+m0OJkb5pGp+HrB7RUM3p6cMKlK7uP6yyTUf0CJRI/aB83Zo2ydUW
2tozG7gnnKGa6z5uOEzg2pfJ22i7fvU2AShMqdlyOAXODieShucKxUkwdFO23zSnFEIP4xy0lZKy
qO9lqy1jVSrKbAQA2f8M52+fScRvpSO8ZHHN1o2Btp3MhCB1Jm2pK5tznUzuFrIk7keP2ng6Ku7F
VoBBHA==
`protect end_protected

