

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
ISK+8BrzqbDVc2hIh4k9UuGvqsq6yFic71tfszsK7KRf52jFUoK33AosGVUYsGH1pmrUc2NUQcDQ
LseNrcojiQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
CxxZHetyKRTjg1ePIJzq+w/Yg+inN7g9nkhYUjpPSXav+SKIAQvdh174FZUi0SnoR2INo+rdZ3gz
yq46XymO3b/3npnRNCCU259giTvnOJxmkrtnjRyUpOg8jB2jnHg/f/BlL3OJUGGiFonBs+6rnNvW
4aiU6ycFpLQsNzqRlAw=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
HZ1Kttz7DNn3t428AVZ/hrbCqljpJfsdfcEo7T7pfqxl88ELioDFFp9rVcvvZiZMU++45qS8CpOD
SfwcEjOj8ndwnIsrDamIUHs+Qm4vUDDq8EtyiGhux+pwMtpg8rH6kCwLDCkdk848fWRbBOGctdAr
AiQz4Fie2ectzKGEhjERjquMNqkQkhNIuEu/CSTnyD7KnG+FK+llVBavN8lxjWeDvk+quMyk8Dbo
gA/SdzYI7TCZkNEFS/PvF3Z8fPBK4pBWz7TyfdHacMjMkaPd5zGsPBmQy77xwc4m/sfhM7ZX+YW6
VBTILiYtg7u194UVgu4fHE7f45jr0jTur9wbVw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
2VX2NPBJC/FYSjnVp8ueqtxuxLgenRIKbrff8tdhuTb77js7o9S4OVH2n84fEyvr3hl3lrO9ekVq
VvQQOlQBg7Zv5/tFAeI5YFisgygYrqeX9dQcI485CaCpeN9nanYXhtHWROH+ZOYckBZHUhhjC82p
LnYwoausKSjsi+rXE64=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
HdQIwrCqCFDZv9OQZsva3DMtF+8TwiePvWLQndNAXK/1V46C6C4sVLdH6SK4FvPis45PZ52T91rx
x7mjaMnTgTVkK+VoFF3Ej7xzh/2PoR+YkiToyHCbvwHQXXvv3GAu3HyqWx9b4oOndnrx5Z1mco/s
lNgEY825qOfDqrTkPvvNBXThybVoOKs2SBHAdaQhQemuYVAjS7mEC/lA7vom+55/0dhIN44Q0vMz
6utkLeK9axPmrUz/LHNLm3BFQsfvacsQoIQe/Y7g5V8ehxANfnzft/Jgo74fJAU3odGS++0PsHF5
2T1joNptoFFljB/U6DScrAB2FxigoQal7I/OSA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4112)
`protect data_block
Qy5P9bbwCPiyercJ9ubuSx7pssqjld5jPEdp6gkQ+TVhE9uD7/Ba9VjlTJyK4jgWHnAYQM2iblCM
wNEqXWPr0WAK8J2aTanKZDRbvfiKH5zeDuC6G13wseZi7ZfRc1A5rIMKkVCf+R7FXykWq08RngWY
o7vgFLRxyhiRjXOH7HkpQrH6HgEFmh4pHO6+XkW/bk3nUZ5x+UD/MwMDSTJK/Y7qA6zgFU1lgXYK
/CZlANrczpItdK6qWvNY3rnX/rYMsdJOmnvRq8Va0IsTlHfq6XkT9t6rduGO5JjihAO0r6l8NUsv
gWQ30CKqa1T3yla86UaGtWq4QLzsgBPOj8OboD4BcClHr9XhlH/u1npNseSETOr/1FTrOmOn690V
B22BFey9vhIyySeJNK3sjkMNbnPKq7mx4b/5ZPrrKS6TogyNoKZUQ+Sc+jPRUduhY0tE0mHdGT/t
p+qmGXEPqYwdBXPpDn2PtDxW0Rn/FLYCmvtRzuE/0lG2pg/H4X+U0CIBfgZewnPApL//w8LI+5rf
vuz8lBusqDy3i2RLrBhao+J7NPB78NbE/C3NzsXaEBoPLXVyABLP9Vk2A1LVveWuPERvYJp5fyMk
Y1nGieo2geU+8nC8I7qXctqF6YI/5uREpeMLxBGBIqEH1zO0qv4gRlRgAwQXgiCMvB3prcMU6o8F
BOy2Bl2bTUQZpR//z0cNEdZWhQKuNl/a0cjlS26S+s/xvwodTdpAn9umIzCWm64Oi9N0pGHKfqC/
ID83iJT5g63Y/5O8IQq0e07GUfsBbP93MonCCD4Eb5j9XbXQfx4ElqoOIBD/OY2HqFY/K4tLCY7/
1PR+0SOj36IdGccyMBFDhZyetZFy97LK11XN9N6PqAg0eieKd43PddgMzL52sTzRInWYT9/dFZk7
I0gz1UDdifZVzlFrYRXWoyauwm35ZimjOHhD16JMAAi4ry8/Q6K5ctxdsJCY5OdhnVUf3JPyqGHx
Una07EP47SBE3nw/s3N3KCoB6S9opP/2390XsAsrDDryqw3QzEX1kEsijEKWki5Og1zbwZMdMvwx
cgeTjINKV0MEv5BOEMHu+9TMB4fySCM9W66I5y62DMb0XFf7s/zxZTXvdkZJb1a8CAGN93YE+FnS
3AfV+rmrkerhoGT2PbKo5fa7V3Vvlbyidr+6D0oECoh7YJ/2HQxAbjgRyzXWpbsD5oUAEKpaZj8e
77QlrSEYyj0d1Rkk1wzqzczNjptwOb5DV3jjEH0/EYJSkyPE9pDEvr30Gyyur3uZesi9HX6+k0zn
yV1ylNITkjfdUpICfaKAXFILWZc/naJa3BIN8V05u5EwNPr+mGQfLX8lh5KJQQiuDRGbviyWyGwo
zx+Z4uHj2khRTOowxb6mLZApkhbp+NMWJN45aK9d+6H3cCqgcNUrx5d/Ni0PwG86FdA2X5IvHAVA
tXSZMLEOzvrIUIllfySO01bIBLh/I0Z7qCQDJ/759rp6Jw3VYs9b7sJ9ii9/jMMFgALIBIPu0wFk
DO/v0kIGM7deT+zwR4kCk3N/4VEY/4TMdrdDI1MhhS4HFcO1U8OmvUygDv4YEyTElszmtQoqE4jS
q3fg1IbA8tp7EMJw0oC3HPgC/gW5xy5m4GnmxwqfyVwWQB5Tt+2H0ZDkqDypnF9AsdF5sII2O/fx
2MS0R2y/3qxgJjSaY/w4pPBRa46nz2qCuiDaSWmV7MFPSi6UiNtu/hKQ5xhOfc8X0s+YkXIkcECF
/oxSCvgsJdqaRKYkOOj7JRG3nFhAuGJMAnZ6g1DZWhUFlLhZxpapW6G54/Zm7K5n9ch4mJhWTwKz
ZE/nf/rtm+GDyPrjz7jxPxOAEZSQINyec81X9aQWM7CZ4up1c7epGKJi4xfh0fKtZkkA6IL8Ahj3
RNLZz4YHRuwfmqKgyDj/da5X2JxhioDgvk17fAEdhw+2s+IagtDRU1INSmCJ2PLzJ2QVfLW2Ykp/
SdeN+YO8UrsX1udIKyA2371fvl+BvW/vYifoxhhxmV2PFYZw96AJNofT9426fi5Wi2N7iAga6gfw
ETgfoti0WWhMOP/vcxXduOTypEPgEOeRyTiqaKJ+er2M0BcWjvNchILoA/KNovE6oC9DsN4sbGPU
buZ85YVUeAl9W+7B4Uszi7mcmfGjO+Qhnspmwypb7zTkJdwj8e0nbVyJmbBNwCvKZFn0I5xSyzwR
Z6MJ14xSHgzP7hF0wGiNUt8gWAYYw9/LCXa0oD3lJfcllQsDwEg0qiGPol5E6WLrxxdpOr9EsDJN
yoxHp07FhHLSsYd45l8ErwFAzxkQDxw2jb4pwrrUNFPhazWcjJs30bwjOaaKXghBbFEWpgZ4y/iW
1dqI48wwcHL3G2Jl0GXMZFoKT+slzfIOBG7Bvu79L3qF42BM2QniC42krd9+paWD1+bCpxpvTpmC
tM61O6nG919zBdL+kl9vYL2I6gKgfmhm2JUxX+bndko3u87rQWtyPBp4DeqdWaw4bkMhXK7lP8Xv
mfJvu1ULxHG5Ofoa5keLXfS4nQrqFqymNAtuisPUDDV75LvYTkEOfzNUsCOs5v3YRYx0J9peZgfa
DxyHiEmoF+iJZPGxThLHgB38uoZVrrZqNuQ7mUZOWFVH8jahpgyogU2Mnov/1Cu3usvZtuDe3tuK
kl/khdW3T1H545lCmvJc0cr9GsGyymZxRXQUqHWWzAkDGhLdwJd8q5T3DUaWxm3sr/jzXNymksII
C73kHRDOr5rlqaoY2/KRHkxvTLBotXjyS6P0AYSdCFkHiQVODNnqQ+Jchb7jgO4v9XRUFUEvbecF
gYyjZ75R1W58UviujHzsQUR9MBmYeWQ04dxd1fo1LnTriFVRT+5tATTKTFd55TFdHR+y4HR8qeb9
5Q7FFOlEudceIFCxHBHQPmp/BVumMfn+KI54zA3LkLcEvFjt/IpkVNrPWt1XvA+m5lxPAzVzz/f9
JUtXE38/WcHazZMNEfyE2+CWKpYXkSUGgYT/zqxStxAGnvvcoDBeN/DXGD8S+1tZYQj8t/MUtvml
dXa3/2ct6o3tUQ6QcB6+uqdTmwnUHxDHbGSN01FBKfiH9nec5w/xq6L21/uQ2G0E5++8AvoO4jec
Bhj6OKfIk5COaRdEzRZ1Rh3Jyb6X25Q4AIw9s1tf1oilS8x6kUNlZNO2ktkbyzrlTur+qhUD+yX1
QrIu8cVB0mvdRZgDy6DKyrSWTGNUSaZiYNVw8B1kmVJDJgJzivo0sFmiQJSzxB7klT0ebDdW6XFt
Vh4gTxFyXIRoqwtRH6QRt/zUUAXKZD4CxWX5wP8mc+w/CPspiGnqhI7FNRS+Xj33Cm9NgaylmwKG
CBUQW9FNv7m3W957dUYV1TR6BWUuXJpAZvr5gXFEyyJVjd7goQQ/iCcef8pPiRtzp8HP1zcndpK2
Bntkfh998xvi/gc7cmvKEDMeVHhvnWmB9Vp1GMe2xPM+LAtuO8FfikYfC+rHJuz8LHZNiHYeeX8a
y0uujc2c1AKq3d/YwBYZtxAvkG5hXmjQBJKVnUAIyT78SBROpsxNXNfdjysDS7nn34l2MF3hsSF8
p/L0mH/lHdy73z8tegrDHEjCaumNhfu6NCYyLTdZsyMM5rC+8zGsrxEJ39qquJkyGhs8vGsBlcFx
10jQL9qG1OXNEFQxN0RnbYVZarZq6hO18vNGY/w7XFqdhjLXBKvszc/gzXirf5kKeVwm0bZ2HiwQ
rAkLbVDJZal9dgtLL3zoS/VkgP7nHXIuTA0YK/sBOQlSvdEsDTSZjI4K0c5seQnY7FomRDuBjsup
/dPI4be4G+fm8ysFBE6FdOmAq1++RvoUhnHL1Th1GXoYfhP9nw5UV9PFOYMjAUd8Jrops50GMVlp
itgwbxkuKsbdUAvoKYAVQJGtOsxnFG7CCcIq8HH4D4byIBuB6km2wx8RwF/9VJXdt2FA5BCzDhQx
yEYT+RBdbMEM6XomPK5EkfFXw/4QLRkcMb/7ZUA87YNSp6JfdxkhKxaGsqPhowRGH7bUOmVFsU0I
5oee/UagQYkF81CjsXDN2fo00w692T3XLs6WGSmJL5f5FJmbW8mbUvWFy+Fc2teO2MYdhFcg26e1
GPN7VScQPeEJU127P8fYOc8aZEEdr30R13saS34aCFXhZoGpD6JH9wW6AbYnPZumMvXxAGt3Vjpj
vqPNnlu2ayffkI4XaEhJJPIc5wgEn5n/o6X8aiRAfScScl+awYEjU2q7aihktZgmiOKcmFERgfcT
CattjzCWQqmL5OPx7HS6YxHSGO6OjUTg21ips62KIiN8Li9ZrzzwN5pliM2a1+sw0PKOv60rHrri
6MYO0u3s65dWq8FZGI+0KvWCQAVkYI5bYEQ/elUtoRtb2zCuw+2X2Jjvab7QM7EAUXLWcg9ZMeNY
I5tUpSlB5AfWW+y4XvcOo8nptGbEPf7y46IPLkr2b3Wo0gkqBJuZ05lVFg06LuxXUS6cCJpfXcgx
1K1HOngj3DX8LBqmgYl316mHThXJBTV3DBJKlLiyDx3g2aq49F9pgkBwwdi/RAV6kjLGv982QJ+a
n0y7iZI6pcKItDBsVIN/zXgKh0edjaznIOG+QQaVJxJUKBoQvJBURa99qinZQSMEYlGUzY+zhu2F
4Uhv39f+BH5cbi7sx/sk8dCOjnsn9w4uS8tcGXvr30IYnlGJOjgpKphS0SNG7ipgWhsLDe8sgkhl
HI30Vv1g0Yxsom70Z69UKB8O+4CR95VHfhbzdUllpIKvth0VQmfhdFZiPTATsl3wUZ2KrhnMDWyV
mnA/JpWdrngSSupeKc6Nm7hUdYDy/UynuBRs9czdM2ffn/BxKNGxchHVsjWnEXBuqYaMULpoSVOM
ggg2AxSF5at2/gB6Q4i8v8EIUV2IjpJ5t5Qy2MoRBFOnYdhO28zmjpBWpgAXMm4z6O1+fu3WsdRo
MTDVzjg9SLEIcN4lE2pCSG/+x+ooQ6HVMl8qG+tWks6qi/UZCSOeXPFYnlJi+6uUIE3PJYHOAsbP
lTiUlz0n7mDOm3lY3BdRsxArxGW1H75VARw9qcW5RUyrqKSTKJHdt7pWLEZ0Su99ZXnwcr96idlX
5JW8KB5MvJ4qwpaK05E5hVG3SaZDuoGuUJMIp3zOeiQXXQcEi04wAozRoFFr7yoyts5f4Gict+LV
sGqMLdWHCB2Bt1Ej74GG3GV8FFOkJkZ7iHzZ/dywEe5/HgL6MOAvYY5SDMCuX7Qj2ULU8ChjvNGs
dKBXGcTzGUeSxEbTc+ftmWO/dhtIMv/FtBFG2YKzLCqXP/WiuXvPHD4rBh4haffbIIa6bT7mwAQu
k4h89fc3JqbuJr3UPqI+stJgfIAEM/42h5jRpSYCwLE25ZxNZ+hncZ35qnwu74zdEFliufPliYBC
r3GEaHEqvFjrNus9ZsHClBOUw4+Zf0c/MqbFo9yVny9JeXPLwVkx9KKZUFlEMQ9YvMu9c4l7wQfO
RIp2BWxD9fY=
`protect end_protected

