

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
dKfOe1Fgzj6faSFeL/IK/IGbXRIzt9OQ8DZnq2KAQwbAq1xs/txiDbhMB5jT5GTGOpfv1lX7K9mJ
mDVaIsrDmA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
cmnaZ+nYMcuVxuKDdMnuchBB9inZOxPR3/E/irYVdWCPhl0UM4JuWPFoKMQnAcsoQ3vgnwO/qltn
0x8JvlvddPokOTwabXK7+R741NBmTaawP5Y3zobRhI33jusePpwNTanCHaHjalZxzALXRseOguzG
AwGiKgpBkrzwT+frUqs=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
sUxQSwzYYe52m4+VJThnA3rSxL81p7y01A34NmBjYzEeDRUnhBCVE2EYcZxUZHf3SzWeAqe17qZn
+OUEYPsHFdXLy5QnKWkfeT6eelEedeGrqLjWta/XE+CwvggarDRC3yCpKHD1RObvSaidPkoLOQaz
Mr6i41kRIdL7xQbC4uLsdgEZKWh/fWAVQ0EsVnkKqE8EuxaCZ+UTjEptEyr1FyibFlRQuCcRV1zc
KGcqqHxwzSvE0/TqNDvaxlN4HZAny51ra9dxL1achi8jzJgZlO8wt9Agqbh7GQueaCXon2S1zoWz
ehgKeTmxlL7ytzeVDSpaRq2XKBPlYb/82fe70w==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
nlRZm6Q4mAeDfFS8oXcdcSIf6QMcM0qJWL/GpoNfKsPw7GwRrG7w5Fv9DZ3ev8dGDXi3ZhhDXcQa
Irin1hT7IkRZSupkXr6uysVtJeCdG/feYDkdTZzOR87EjbK5yer40aqraNg1lVIuObcgZ8AniYE5
0hMf7gQTkG+H4+tX0yk=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
HiHN8/USAozrVtx8xCHzL7SU/8fs0dpiHUe+Pxq1X1HHq6PWwlbojxR2di+cVlcr3m6I0F2zjyVW
WLu1kh2il765GldD+RCzgw8JhGbJOXcaDKXvV9p6bqICOBy5WCTf6gQ/vOVRu1kKDvf68tu0aJcM
5GW26Rwq/4L2jSNVHzuzVdgC87Mdq7eVgLL1qlhKwYslU6Eg0eOYTUfGfgCo2Z6Lcfi0atBesKpT
DSbchvClt7fyjz3I+qeNhclJOyfOLBdaqFIyBSFk+zxyw4U3h7toqFVwQu8Fc+NwLgyBezl0ZUBN
S4Kep7fupBYYGAqkU2vi+UvgcgkZQxj4+5jXGg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 14000)
`protect data_block
j7Yu4TYAGnNQRO2EeEZ2l1451fZxwQ5tgtDwYpEBkY1VDMVvmq5hi1EgO1OquAmvdwenYjkGX17/
0R1M9kdYnR+xN/PM4zhK5PSUNGXGWcCKx/SqdmtR5Dfw2dzt72LHp1r6IzC21ozQRARAeIUUSfy/
l2LrjNtJciesZZABoHGcS6KFrDVd45C8hLme2+KWFqcJg7L0HQF7U+ETznywkALVanKFXCP6IBbe
JMv97PQI6NZ8VZaNgeSnuWufumtLZ5Jk/3iDkyEwSpxidbj+8Czd+wzeavGIf5S53T9aIJrEpGz7
Uwqsr3/Qe440v0ztfw6rjvisDWzCPlA8xsS2VeiRA7Inkc4WLKZeRqQ6t0SGQrHwYX+pkWXflcvh
nO2Q+tZDWPUZmQ2Pn1a2s1cDNyIV3wXfSNJ8/QpZHxi8oVaVasZZbpTdfprSd4hRvi1tVeUzTLJi
wLcL/wdxmrall9XwQVU+ZjehC/1sNyPtxvfNrEbInREg+Ve2ZiTHU8d37JLIRNMXy+Q4HUT5vwJK
sEQlRLTIMx3ffmOc4GMupM6FPYd52pk0TwjIdyBl1hSeA2w8LbXmx0Q7P749558QUnCZCv8FxWm4
4BIg8WFVAaj5rT98QWCyOh2FKnJHidfua/rtTIV3XWW+hhtaDxTCnuWIW0aPdggvaw4Byby3mErV
WGgvMQiu4Tv58LnCOslwzLxBM5X6x4ipn6pyeGaoq4fIKY8guKUpMbwn51CO48NqltSkBNLoaGO2
TuJHq8bMhqYRUhg4d7mmV5zDSKdWgartZ4Dd6v+JKdbX/7zolGwpOJCLpoyzjotNZgYECsqLaCFR
HUqLmWPHbdAMA8EFCVhWAY6fEZfbSHChc/HIZOFJXKNCiYq0u+F8PKLCgKhiafTQs5hWOt1Zrj9/
HIUBKirb+3LFi962n9tzRBGaqeoQu6gSpAsKkKri3fhSJ1lf6geoRg/NCvbMzZ3x3ltzwjzOHUvj
2zkQH1Qg3HNeqqpE4s30LUWqNNk+XqmfQ7JnHzkXfYVhwEwAcwt4GDXbnXpv4RA9epxVeZsp8pwB
z3/T1bo5gMTRfS76DsznrjRLPpzQGaCQNNN0rila660u57uimGhHbaGrOBayNABcDpK7qlu/GLXb
8TYmzvQK8/dy+mHC0By2mn9ApG28Dsxihojoq2NeQ/D6yzoZB8yXeXAqPX/T0bkYLLR8NmfgDOFJ
0TrdutOr8ofE/Zd9wo9MUxuAmKecSdkzSMk23nWtnVQbVC1YRhlmktrWmB268sbphAyd2AULm6AE
E1Ob4+PggPGkTGUkC2q7yv4UIZ+3XUIQX3ngDs9TWEcngg+ZC9Fzk9SDx6gcW9t4rgVchKFRj5Ud
VsQHN6nI4HAPCjgWyz0EcVhDt7tlTlkuu77NRLFQeDuC8JV9AmlMaGl08uK5WDPGbc1l7TyWqND+
PyCqLqjjKy/cfHuKvUc6VAU6m3S+ClbKMclEDH3Zywm2g3Yj/Xk9GHWEaT02paMTOGQ4rIHMgK17
P+6f2S9ji3PF7hDarFp54OpJANTShXLxpvG4vD8bluGKex8S1L//ejgCugLXqDbGfl8A5zpdnYgu
pFr896Ni1VnInQjuSYXDE2RW0Cgpd3oVAWYPSh9b+QlMgWh7bV0QtPt3qnohzeVSSr4SFwsr5ASG
wRNQd32EREDucaN6WZa/IIMZlWBFh+TWIeNKhBufWXnlnOBLp9EQDxt7S8+8s/JUbdxFZZCcbbUm
FX6CKIYa68eOoFnJvilzzkq04jliLzHOzv2Chlrw9WCYHLK55PiSVcuobfiImWc90a/Av7cN1xsO
KkOixvVHDYCbCiRwn4awSPPnpbTLeFhx7lNJYMml9y0fy/HSYixy4XauVra0+KthdpnATX3PvMzA
kzVzoI1qBEeYLXZy01knhGPDinP6/AzjgSN6DvjylEvJWMRSTJC2jnNVABQLXOishdTByvMIvbiE
iu0AXisDX13N+2HrxhsbQk6bsjH/OFivzxNknSibxE5DCaQlFHyS3G4+JYuBMPhfKtLTD0JeK1lj
udkpVJjH6jkk39rLqn3cOs/lMAfAs3kxsUOD51akt4zk+W36KZULbABD8xPwFt4G2VFMh6Oovffx
0sq7ecO5cRQHA51rui7e5DhNhh2z68038zzZqj3ScQcw8cP2w4dlo912HWc7rc8zgWyEQwf07+Jo
vztaoYaqJ0si7+f3KbjJynWcmJWNqoMS+WY4UuaQt/KsOeebmoCbfaKSqcDFvfmymr1l7cBiWuTN
26kjRP5D9m94eErO7i5ZiZ416iwQfu/Wcaxu6/lN2Sg7cHHYs/ARzMLqZHFZK2ix3QmeK15alnv4
HxnwnMlRagT24hPRfWVf11Fwv9s+9Z8dLMCdHxUKwvOJhzGKzHpu2xjj8YA20zApXSa2jd/Pqj7/
m0zYwF+Dh52ToCiVPcmbVMQmt4Z6M5zX9g6M74wR8iLjTgarGr8M2gSvkpYjYm27hbDs82j2eTNd
o0okCuoeKO3M10ewcmNJsgEM/GNHeyIpXzoQwfiLsIp+BFtnrezRfKeRnUq/y9xbCjrKHuq+svSw
EU0pFrLn6SQkIaLG/6m7lbg3Xnrept8Sdwtk/GHYFKazYx+uJ7ekx7JMSCVmz7JXEY/Qf+hv8bHv
2lcN2y1PFoj7P3eCcxic6s6wYDKsm+gaqa3G1gIOcsBLjUgkz/oBK/N4+v4C6V/xdVXLNDVgb/bI
tLoMd9t/EyfWzCE6oYC8fjdjihViC9pT5zwG6iWLr7iJVxF96lsCkltiNWB46/2uKr3b8YiL49LC
45yP4Uky0QvS1XalPMAHHSvYHI5AcghufjoGNTMsuwVQ2cPg21og25hTTwJwO/UHEuRM3x+64B3n
WPtLAouTene6xDgo58AocX6wJkUlWTL93jqryO2+PzTQ8BL0SYFNvo+ipHz4Gn1ztcQlNldTW4BA
HSt3Kv7DbL40ZIJtNdrcH6VWB7REFlFsm7HBSEBZPyFEJjVtIktJcHIQ3Kf2gscOfKSwuFotai+T
FK2r43lS54HjUezjhjxTtnXL2hUhp/bD7uarRG+XReIyKnjvCZd+pkOThBeGO8Kys6V8P+J7UUGC
982CYXCdilXAQaqKxMYY8eDgm789Y6mqodUZMb49E74XTIUyrYlS+Xgj0m6D5+/16ml2KeLUaxRb
As3X53DltaQBTDtfUiSDPhdMy96yto6nol6F7LNTQws89YBVyKSyV5y0WW4/db2gP89GBxk36K89
On6zdQENFBZhGfOxOzENzP0/j4jjqadVYd29Ghb8L3oE15tRsiWZFyc8ZmfYI+Gr+N92fe/ASnhv
4ajWPuilRDZupC1Hp+nk1gx4UE1B53HJkvplwNcw2eY3mkF/Pq0ZkNqtZYfbVLcmbc751OS64wCX
1/VjIxUM6IBAvH2M6Mm5WM/z3awfVit2JLaGPoxlXkMd1uqckh8sOzqszpjIwLzL3TwkLdlnj3GC
vT8M39vhCXveUd9nyPo3Yt4DUvdnHA8n2ZIrnNGenP3vS+TDcRuAbxH5lTnQSRozmUh9jL7o5A00
S8neuUU/GLAj7PDG4b4odrrgebEJ42NArzQGbbWqe6Dyz/VyQDuyQvq3o7FDHRx+MlHu2aYh1bgW
jkocR+GYyJKUVZU1Tb3se1MyNSozDL5kgma8OThOpNhEl5fKPKEWvbDIX+kDDWUhwMdCX0RRs+in
hY+aHjM5ywruxcdmiTItaOZOjEExSJZBUhcoY054aJJsr32OYoQtxB9QDQwvV3z0Deh5f+/4wSwx
SgZuIGrM91p4O5bzEdmeBg/YFm+YI9lVvQqCF14IzHAl6cQSxUmUfBkw5jXmy7jIdGCJ1fmqmJmy
gVrF0yXFmyxR0fq2exuE1MUMtPiM+xRQBQY8nEBo+WNcW0KBY1HdW4pj6rmauLkearzZf1KIQehq
IINg1t0kB57dA2nRFSHiapKl33oBse8x6Qx/D4bwe3Nz/JNLsJvgcJ2Isd20HhQYQEY/2oI9oFmV
ki2EVTZRQCEU1VylfxdSJ6UuBZoNbDTdW5ntpAigwaDuCILj+KqYGSt7Y4ktslRyLSNbj3eMWz1k
ZZD3nvwR9ilI9A0XBKteszmntiWtXi5jiIs+MsCRCRlaT4+CscP6aQjkl4xxMMV9OESHTpIjQiN+
N719XElqhCbJ4L8vEbAQlIpUvsPPjTJtutPB4Rm+WvgVauH+sywkPlZlNUEpRyO6LhSlSd65Tplf
/hmU6hbjcuw8D+1QZ7XubFjgjHzRlCplq/9rsEsrDMsezswgzGXXVzsiy/pM7mbKexx9tIGXGp7c
TrVFpUODwKf8VYAj1ehsmEOg8Hj8beLz2s+EtoD8oxFyiESGkTUCSLUfI+PsQqzyh3X68qpk96Y/
k2x5tetYIvhMGwTFiXeAfYhSrLP30cbV8o/KrxqwrwpdcrUatNEFx0wdkoM6U5jAFmJEhRi417hX
fdZOsLYzaXg+CEHYGN55X0EsR241CjzAWKl3AT8W0Tn1wbNcRCMiO4/49zSyyLKWwHZ7AbT1SXz+
jQWGNBvwXNJ0vTLw8HresV5bsfcrbukPnryyy92WMSpDpaPtRTbAiLvY/F6jrJTRk++5YPgkwSjj
UpsRoaEVjyJS6kh0z21VeT7gWGwniLNhRIQvX2Cy0PtidAIV/rumgBZI9ffv90wVmhNsl1l8ghm8
uzAO7wsubInAbVnewRaTnO+fDWD2NrD5g5gci465EveSk+WwsD9cX7gYFMnGwUko6F0e8owojsmc
BdE8F6BJ4sZ+u8nA0SJlkzmYlpEx/EpaO2BZu8su/cM0lk7a7b72/inykflTn1zm/7jVcf0/YX8F
T7kUcOWfD68ZX3DJxWHd/+2hADahMG/Bvkj3F4srun1mgxG2FBWfkSeWwodfdtm6GkNPejDIyYVl
oN5BX0hP4PNGzQlF1yApfPh0EhqjQAfQ+MRoKjERRjUH2PORlRedRtSkjLYMzXuLQYxitd5YM3dl
2X3A5iz5jSyAlX8YP3AWCJbWfoUi9MWNq2PvWvBSMIibUjltqC4RUk+YiepJoJeOjaQ9aMSZlZuE
qerRdAbNUUZrFGl88bxdrt7SrTjdk/6F7QEEDODXuR4X+hE7lEQFEl7ubWogqs+zea/EKSAI7xsb
Y0HurZmfr/NJ3FFJu/xat55u3RNGnnohpfDFESwVQ5u1gGV3KREGfJcVqKVX/SyoMGbc9vn4clTQ
1UypKdVezBgpFf+E4MEZ4TRNt6XdnP6M6cku9G5R4htIUYw7yrj/Kt/rijyowbpkceGdexnIk9NQ
mz1NUZIzadyFhpmJ60gM8LvElY4jViTltYYVRiNyJlLFLHHHFP2Ntfzz6LkuoZz7B+jb6hB4CSpm
LbYE/6Mi+gEYbYnSvXzi3dPXnxzOh8E7qVFTTNvYFhMQGe+eOiz1v7aEWJCSKEtMmL0IVSwq8f3W
+/XPfwUawLwLfNee0JFCjqYmiHlrLECbAQ23GG8fsjki2pFZZeRZcqhxIRNdo0EWBSMSLbGArmWD
z9WVSqdAmX+KBPUFcvy/xNdS923/abYG3S9jmu+E4UFho3MgAZCDfDvPulV5+TJP5UxH7kSkSPg2
qb6P+/z0r+elIr2oAZoDiFWseLBgtz79uwi/uTgCAj/x7OCvuTS7bGTMrTsRd9rpmP3osHXJf0E/
zzHcUjHgwAz86JfsE2Vy7WW3/27DfN7jiks0FYcBxaNfUdQVd6WAg+3RRRBCHTtU7yTAY2oMAd6z
WH9pXQYPoKYJnE3f43fpzvQ9UJxeKhgx95Lzby1+kKMIkWjmmCKLt2vz5gJ+jbGwMr+CAS3t+5Z+
84UhtxKLCYKXh1AC0TGUWbxTTCdHIOTbpwR+T9YCZBxN5gf4yrGmLmoC+u9md3ZjArEfi3IKUdHS
2qi/C8sY9HHq6a/Y+qKLkFfz67ZyhNbQbJkv+Ztwi0GO2l3CZkVJQvz+We8+ImEgYO/7tTun8QkD
H1PSbzgEWKKbZPBDi2MZO7ED6TU9wZgSBAZ0q9NtiuAVVUM4EJQf+Ivf6P3RSb649p428PTD+emi
1xJksi5hW+3DwDJA9IPQGTLXBk9MaOg3J4sS8C6YvsifPsSNSkUvNNebUJgRwC3g7jFa1OGu9Fxr
jm3gvPX/uhWaMflrBjc8Y037K0KqPm0rhX6CgSm7VgfFNeuB94HCojTXt9QtoASfcm5+XlaFYeWP
ciObEd+PjYQBSkR4vldmDdyK92dV3y3nSUs68UZnqtU+7kVltOO/uBsyskguud2y2MUWqiVNV4bN
lcoPSkkiAxucE8SoOzqR0nKnGxwKx0248POwB5loSC8FmpD4T6KMi1c9M1PyBUvNrE+iEw8gahiP
8FkC/RCauILUSdiHtDrToHyUmxAB8RTp/5x4fvqZI7cRe9biu1nsVmNW6NhJqkJYE9XmcEIBeScS
i3YKVx2y6iFbQNzlTbWSGsRK4K5OV003pBl0YLmBGB+whzaFWQ8LO/uwgVItep9QXBNtqJv18ny6
FN9XVqeBS0lTrhEmNbL3AFqK7fYT7FU54YUh6YVbuLCbLebIxvCF/JOOP5k8vj0pfXZgX4peVg7o
rAuBjXQAiD8+o4uvG9FACrceHk9zPGDaYZtbbcUv6Z764t7MhtBq+acQp5cpB0EVHwEfLnMlmjW3
DCmJML9EwrAI55wREKRZEYJZ5LcIU9pXttNDEoM7I8xmaV6BoR2YFW4LmdFlQ6Mz4d3LSRigjJKI
HGNVoLy7olqPunxMCQJIB0roDN9aMNljuBcXpryQ2B7HcHljgDZKw6bhEhJIdrs8X1UHwLuizU4w
WKTEQEjlNP0fwLpS8ttwIZFJm8YOo1Ju4RvgybjH7oA+CO+PbcKFEup74ibOemDTs3YTqE9sdDiC
OQ5HNKROkQHeLmzq7uT/LqCL8xFlS3L/TmyZ6VNEg5+eMCK4XYpkB2Z2t0E05+XNHHjzviAXxsIo
gc7zkeeikZBOvtQ3lYknFIeGY8VhOW73l4LbehwapTQk7+a3VnLQASEnEUcF53YELnvTicKuQB01
tYSznXFIsgWDlsvdCFXSVc7Q4cqWfruKViGJevpM67zmzI+uH3mDWb0RTi/a82MrEGbeT0mtckG/
v3D+eCqubbrCVP5l8VAzM2V4Uu9d0X47nJL20o6EVEGY10IvxderY6woa5I/4Vcc1SFSkZmnFIGm
xOM/5MhIiaG56Zbi5sF4+e8M03sxmycnbe5RYspzzqXNCWCYlJpOgqqm9Bc0O5Oy2Ub6xZFiAGC8
jX85UopXSRtnZURdludDnuENENbjhh6BYFRNBDc9oz5IrTyHn1qOJBIy8ZgWjhwoKOyr+sWa6yKO
82v5j94rOclnxIroB/USNbyzLqY2eKd3M9YsdYc2bxb3qu7135obIpOdJ3tKr5Zdk60secp0Ovdq
b2COyn5qaQsynq7Ld1wa2lk085P3DRieiYojS1Q8GTmvVtUbycfW9gSU66yHrtgvBcdoA9ESNP6u
k0XgdLPYauVXIHN5YWp7kjO1j+CRw75j5HGybwqMdoUWhbyBRVrExwERmCEPobBWht9wcFuI14rt
F0TpIrZC6RyNtVkMyLp9gP7j0DWhadn0m4TGUPPur7OZ5JOstqyGAtzXf+Rjzef+f96nW0NgSjrP
7EGMjt6L4mqu6B0XCJhjE0P3CDMHiYu78OhsdX+jxDasXj5MBjwGNp8jC7FxATl+ZyuesLNjvmtJ
lvCsY4eUnNg260mfaWUAx/+Zie3eofaYCs74QIJ1iRGOG1jjpaaydfbDWUGH1YmL/A8ToRgN1JXs
AJNpckg+QXs3QinW09dbBqX7XuwmNLwx6XPFsr+EwJ+g3Fqa5sTtkmz8Mt0+BDjpLUBIBoBQ+SP6
vzaMskza6n/7dlHZ0wzJ9TT/qDaaVUZ2SNt/Zhb54k60OIMORJ4jwQm0UJoxq4F3vz5O1u4b2EQZ
5Lm+rPwwaYDH/G8lx93IoDtnC/na7RSHS7bq0EZ6y9OXVP401K2xWXlmE38f5Fh00bXziAf2Frxi
f+pLajnxwMFjM40l3ZbxpxmQAmosd69AU+x86Pp0TyNjO5t2CspEvjv6i9DQ3BtI4H9U6GlFC3gG
9JJ7KgxQc8zsFJ3z/nnzxaXmGljzbL7BLkJXrPH1YoW998bY/ID8ZY9qA6tkE/hwkCZ558pu/UWL
j8s2yBCOrBaIySGDCY6wGxgDBJlDiu2B8fJmpfSBGcDTnFvmqOMKd9S/HJzvOqAjLW6Q6ifXpgvZ
k7EO3GFi2LS1UNctFURJXPno+wQToiSQFQa7ZCsbrJWYD6OBrCYiaksRc1Vb7lnopAO3Jl+kSbFO
D7BNrn4m1cGqsl4SZ2WQnR5Oubz1P4ZIxKdKSfAXn7dbNr/rIWU07ZDfskZgPe14/PYJhVMlgU2n
CQQzNSrlI0YremAoE/m5zQNmfAT6FCxI+SNnJX8RK9NqlHgAS9t2nvMJQv8/rKiPVwxDHfcKwOs0
K7YTQSmYUSzLylVNjoT1+pYOmypM4i1PWHZluNHd2Ar2kPBtawaVhHSNVLOVPes/l3TLAriYDa0e
QXRCuM5Ht7UBvyNeyi0ZZlHWY041jCWRaa4GFbY4Y0Fc4/+aul22blla6sPb1XjYzuG6XMA0NApb
lM6gH0AGInMmukNx58GeC9dvlYCUdiHn+BiQ5c2ebItuYvpf2KiOGgVxw8b6mVlFfQtL1R2/M4TZ
WD+sMlA7pzGsxGFxHvix2hIATBXxToFKX8bMYCHbPCUKiTDIryqb0ouAYCEy0NYhoWeG0KY6xXTM
MdHPcoJ66z9wy3mzcI8tP1RZ7UplkAk88tKDIcm0EbKaGA06QK0aWgHtA/R2ZFaHlFpRugz9idoy
ap5+ohjAla7AYFnO8aqe099L4zKbBqbf89m5hp5QmlR6o646qtKpdnzRuJ7XSegMYS8OxCdMsgDl
JZDC8gMg6yugsqsr65bECJOq0awpV3jLZ3B5aMnDcqj+tre+1jsgrRz0uF+4Qbmz/dou2pUwlqIc
5uE+AHCx4008zDFfNM+L6g3YGCs8bW3qXLJpmNAjrS8PVGEN3GQTkj5FJktBOS/5kprNgmuGudFX
I93VTdV5Kyvc1NT4EF2tX0WKT8FTGlMNTNDEV8GpRMUlVl8gr0e35vulDF11K4Zs8vhWOYUv8Ncw
5tacmFk0ArkSUFijIAznKgRJMCrXSbwd0ggeV7vrjiWqjhQa2vq3QvpbXmN898dH2u/AqUMgKpGT
KG5GvIhv+KXN+reROR8rBuCinkLvqJPaqUKN2ZXM6icJNcERL/HuPOZKaDaOc83dkKF0D1fzRloh
/BAeLNnhCrIaxHddNXhslcQxho9kJVd8kPA+UXgibLIQkbpmRnavhWKaMMOY6ZVGvgdA31RsknMA
hjGVlq4BgNsDGAlS3pm+oiO7Ru9Bsr/qKc/KFef/+KmzVU4Vs/wCQZxicv7cwuXE1+5LQr6nyQFF
dwX/3I5LbxLF7zUnbu0F5geEdnsCJA446I+/pKCUflNVVIv9qbDdv9rHviy6HNvYC0tb3BcCK47U
0cGTPkWS3QhYKMUDMEGxZz6emIvW+NFq56gpErtxX1vV4loTOlIrs76tGw/fZQ4neyCwb1qp6BnZ
T20aI5tSYTIgOfhjQ7k60PUQXLEd09MXC7YbNAq0yR78Dl/EsL9nPARIN4kncE1RjyZseigmE2ck
UnTn8NFgZYyyW02wBgm4fHZ2yYH4xMry6ryyRHxtgVpzMcvKKOuOZeOPBX143FTByVQndrw8ouxn
mUIU2oDCtg/fqS+KuSIuq7wrBVeYyoNoD0G0T61BD5oWb0IjdNcEMM+okWgSFL5IznxWmJoP1SM1
zEQUAB0dBWDjXLZKYAxnOnBxnhoR+akN1vKhvLF1QXYQNjMXwHfmpQaAzQ6UbJd+RuMU79hCzr4k
e/rHz3yanBmgLiAw/IIUpdZwGe/7AA0ZIhG8UtY/5JZkkIKJrOyoBOTu088WYzYdLXB5N0lUsr/5
3w3i4m5hA3vAFAVLcEXNMzFUmnP7Ph4m7mZOOrB5myCgVyJADe1+TJjPFWG1Od4aqCwUF5YYvXE2
6TqeukkNz6EqM5tMf13yK34//HmqyuJWbkt54GxBJn3VF8wo14hEememqjae/rz6A14x41WmhIgR
9IUbIIWIXM1xle/CC/iTggK3DOUGDnk0gDIjBYn3JIRvQ1jIoVBZNYa7uiQIHAyNbUt+8QTHoAvG
1LySXtx/I3O6mYXIPejvmOzNqp4G7Pb1b2pRfSe9UQc7YtqrMrh24yydxUqfRNhVqyPeNcAfYAgZ
2JLcE7+tMTLnoRdvl6vNZ6nQEwBfsaO0tshRNZhJOA6ggo+1PFOx4uX9VMMssA3gZIzb3+QV+0QS
h9A+QbwBTTzCwx+w0zYddnRitMco9W+wtKvm288kG3IyfSDHbD5qv53UYszwNMdz2Camc1esgx7Z
Con4ciQC7O6L+L3VYy1EKL2kATplMlWhDB5Cm1tb0ZvwNZkaubxCW82Fqinj51aWyns2syPEyE9q
FH1WFWcHML8KZCujB8tL1le3lcOuEMVsCHMJNXK/nBjOefCIXEnVqjr8YEiU/La852SjBvt6DE/X
BiQwf78TYYt1xsmd4XSGeErFf6XSIbDZk532HAjKjC2v/OCNsAJdsmMEG7IgAOxW6X1Ztg5KFXig
TMkpcObcNRft9I28e8ELpJfhKD/y8iK+Y+/4D8i6rfVQIytK1cjoZ1naAt716C1kq1gAePSK3WOj
2KEE3m444YdQmqvPDI0oipMZGowdtCXCS4r77sVBIO5B6i7vnAQvIbeEOIAgmhMbzTjHB+0AuIx8
IL2Ehx7qHcbgHSTHQ5vask9m3YOdwKs7LsmosafvPFjAHItRutYWx88FDqB1NJQJr/wsiH6IDpqo
NwGWo9PJksZNRizHjvvG8mR6SOFk5r4eqww4U1EN5TvCITQkmaiZRh/+JJ2b8M8s+JTN0jBwvW0b
RdBgq2EJfCNFcZ0CYojbPVCKBAgaTD8vcIgEOhpO689qrK7la6SHAvwDhf/j+39V2jkdT7YamYQ7
bgb8O5ylg/JUaINubY3jlHTcNjf+o6KSIfKjhQ9bFv2rvHyWdYn9qg2yAbuXKu0VBxJAEq/CYbXB
tB5mNiucmF4bZiSUhoaMc8KHPaA/NW7l4VK/POWnT+HpeZ3PSK54/EhEeFXEkJi9/UOQlLfuNN2L
8dCOYF50IRZ92Yj8wninxPm4yVbTGUPUt65wiKzqdv1kCmpGO99f5+gp61ttj3DJAFW/wZR61CrE
d8KCVnr7wQeCK26ic0DfawZg1gzL6wYXLBpbN7TroKobScaIJIWwydGLms/kXZsrdisx7A1cclT/
5t4f7YVG+NxtQ+6RpGdjBahcNb235Fg/KIdzEvPtPMStbO5d8kzr0wpJiXSBL/gU5vKjXIRYpVOy
SONCzGd/QgSoeJqwAGG4R7TD1xgXILHS5l45CMygY42yXPg0qqetbTNcLVPpg5vqP+/afJ1/tr7R
scZ47VofqwXTaUI7gt6glVaYzSqdfoiXkBiJzjxeqglb0sAKRfqmfIeuCTv9ufmRCtPyPpHWUZaB
gODA9wFjANywGW94djzWh+kz4/VzPdCs4DTHNaiuDit52Dxtu5XgxwboOlra6dDhBzsqGUNU6T6z
JyRTdJfzLS5KkrDXUai3dHPrFs787ldYBOax2smux3lu+m7OtSicOAdiGoVhYbkvbZG56DtQHa6z
ZRaFhlWADS+0NzUSkjB9OhQUOwpqOmkJ8wS6Yld4yF5jzwwjf1XaZHHxCvJzaldXaYW+fbW5bW4S
L0wGX/6ms0/yfmdYYuvWJw3sU0dDDYs/Uim5Ktjqj8RvUS6E+4zhZgdXNFt+Ywut/r6lXYvrJxor
IyK87rWquwvxd2BhcoWxSk9zFGrGS2YycSaktGURLw8hhjuYvbEF2pqASEZq7EHNc6SplN9KcvhL
QSrWTm9qeF0qRsbwfJEmzTCDWWPzf+uALImI31Csa3xNUZgPZHDEJViNyVMiRACPRj1+OCefBeXX
/AcSjHPQWZa/y2Kr63G8SkXDrSkMzlyrCsLSEvuhB7q2hlUhxCHQ9zT2DsnEVXgvJ7b9/Q+TI1Z1
WcdS2p+H4vH79uwVxnisJ3HE4Anp9FZBgsSvsuYEuHqO7+CFVxfS6w5Hl6aIVBHgt8zLUg9HzWYf
SbYqaZxHwe8OISk78bTEeqWzhvePs6hKYUWguMgVkGQi4QlJwtUC7bucJDPpn9WiykZ1bm01ykQt
UwmDWoNLRMu4TviV9gxysF3w0y/PK2k+Y7MCpfXy4LRDwZeH61dbY85tGNI4556jx5kg70LVm8EA
u6cU/nezMLpT1u5KTyJRGETCyTY7DY5+5PUaquHLfCDVWHllfAcJck0h2/R7U1NQ3Es9YJWLtxqY
yesKjtSN5paX+7MfThPmT6JGVYICRpRoya3y4LFV7szbaUKltO30RR5yXWJaxQQEpuBe5/yzLjEk
r38Dgf4uPhKFps+AN2FTdMTD+VARsW+6FG5nvEPj2l4G0bna+aRDlOxaUlVBvTxGrwVdCGZPLxDF
2Lt3Lw+1eDbezaqXktNsHHb9vum51ZCJ5wB0YkqLhEZ7Wyg7ppPjhD2PIXOyActRTfQFd09ryku9
DGcJkhIR2iZgmz6OZNmDBlnnAFGvfFSEfDySYfyt6mb4IvRllMmpdwbFIDFrdPlrdydPL9GZZduR
EHwaYRNCBBBwttXd0Wu/3gyJbpRnYdkZkU931xUqpvqK0JYujA5yoZ7coooZpE4AabHPPIjJCg8H
oRXnmCq6Kcl7UCFok4P1MKNAxyp4eaVavnQomkYpYGPz8gmwwam5oq6fmuDd6HR8ObUGT4KecmJH
DJjQ3FQKk9bHNM6fsi4ugozq1L7PREg+DdVyZxOqaVeTTVIAy71ODEI1HhoGKEkGcZlleVmk4kG7
10duDRECe1NOgctgc2WacYbyav1GRMYyVmssPYFWIKCjjP5nS4qDRp5I4r0nzgd7tj40yJmkS6ae
vH0SCbsitl24/uAHaDAM90JSj516yl6aGJ/+TtwyZJzNloJqsB2qbyfe2qTHvYPbsKLVyYEGISiC
osN0uH8VLCBcNvu81mUc/xoQrjdgPTML4wWdH2/emMUE4z4WbZ50g8HvLLiY3PGozGundn1AuMAr
4MijQJjE81M/pl9gb0x5btyh/xAkNQBRobq7grVEj1zgWlo5wGtiSbQwhKKWHDgmewnKSzXGxZXf
eO8xkPKVNg7f0ymSdGg9r0h/ckCEOjP7i8xv0NK2YA+8i/CFvjn4uK90mMZX82lEAWqExLXePaHI
Rzk8xYIWmTiinkEVCz4/D32yYEHtujsXhdSjrkZGb1wKHdA23lXd8muIfoUKYTy75b3RLkRmg0Ik
QBz/AdFSj8zq7RoJ3zrVP5fuW5O6zBLi1752VR6bZTbPAkwyrk4Rbnax+eSLF7uhKxKdtY1BxiPl
lUxc3vgi3fBJOKvVyRCVr1EhIJ7RPj4S+ppongMl6evXjkIRDOtkfjf3i/2L/fvsNzivMn8v+xTT
/vLLXEdc+yRZqXn6vvdAtpwNhBMrjca4sOp67q1/K8wRgjDaV2OWVHwhXRlxN5Z13tsnyEODZx4q
aDzRQ45MB41uughs2y6B0m0xFSKi8+KK1EPQ9UStiTdbZlKjOtVuM3mFeoNy5foCmqimbMcrFMIH
/CAaxAWAaJz5oZcb/wYMdgSnS9aVbLmCEzN17XFmcl1HA5J6LN8ccj9zcCegucXUFWlw82ihsb0H
j6nIvXvZNgN8cTb4itbRAe6g7YpIa4YzdyALJ3yVk6FP8sU9HU8YhwyGKiyjLTtHUDVt9LegxXNW
bSmaYuPJJQFOBncJoRt5Kbh8yVu+UP+XhVUEBLHMrtkaKIBt8mYWIrg5KCg4wblbFOukuX5Oq9EW
+QWk8wqbth5B24ApLqHCj5nmgjQ6m7RZMcgG8CnWmpODLou29ICIb8albrvXbcS0LOsNlJxepnw5
lx7HMyUEYkqVVy/ICYB5kjPotHebrpq8PHYMdXEb21Y6FyoSrdwkq4fLcNN3+lfprbrtie2Lncaz
gamKftSYswHAOOiBkRpLYmOjlfsoS1IRWud3im0zmAMziRD09bindMByczlhRCzqv8wDuFKjLj0w
pLBP9YkMD6n8BN8H8bxQjb0MEWyhfNQCpmf/dB1RR4R8NHlucWGoPPK7eceC0TaDtGGp0xri7MIA
vfyx1pAgQUE4jYLN7MsoC5IDvu8qS/SV+JjuLHviqfELqCTVECkKMk+B6Kgf/HIF1oHCRf+0e/M5
l7b/fGo2tls5GQe0vnaszV29KTRoeLOwAh8GDH7F/wLt0Qj7i4+9RcJNoPnyPJMMwfzEn9o7tA08
7ej4fYJBQ3Ki3gWhWifivC8YNJYbsJCcoqMalutQZ3klG1qUefKpkNOVIlSz5OBPTBkMhoq38dGV
kV6VwXhpQI8CSQwf5xkofvfR+fSatxcwXMWaVqn9jGWRpZct4gjU+chvivpHGW2nNQ/lEnJlHPAS
HNy6CWbW9v8fDbdpsCZpcICLs2CsO8aTKGBNoAjjZ3Gt7OOtj6sQeZNnVj80AcakERzcNcnZajYW
BUHXCKlrIsVhX9f+HQnjXR7BOxwhHw9E+iwZYDanWy5Qxjs4ut+H3IAn8eZB4dJZdp03//6t0Rmm
VBwBIItH0qHoVCjk8+55HrwCY56YBfMB8CwG9DdCCVZN1kK4s6q7hHYYsgPG9oRRIs0+pqwwCMHs
iW+JNINhdiClZPH2Ko+O9maeVfG5OVrC9oI8kCYqHmVliBOuSx6yYlkEd4cagis0VOH+YOdX5dIA
i+F5HA7J7BoFiyLu/cEea3T03OyWaOea/b/MUS8GH5aQfg3+j+wQL+uTVK05eb2n31qmSfHq2elj
D9jT571MuJD1uppKS1LljSO78voUhvOjKwEszU82tjOo0w1yqgWs2bRbFnRki+QwqydoVBNrpr39
AhOMsa/EK/1CvGd30TqdUM/CtDoGpIQa0hkIyGa2Vnft0n0jxSip41Qm32BxuU8yXg+p8Wfato6G
T3tcb6Qlczbeg+9VHcy/32XFIz6dHVF+74cVSERW2bWQLKsiRpfmXFhy11OqRO3hjcJ8nu4Ude0K
Nm+6upwp4mm3P0k/feA2skJwh99Nh+dxs7lVGPeMEmIKnfZrAjuRIhGot16vbHAaQPRfE9VWTbMx
YeTtiqTaeTrKnvqRSilUR7AOq5J/zwGV6KfcUKnCFLSYgw90WNUPvUF81wnrm5pZKaaF8fh9lUbk
LJwWied55z4zfe97+uoU73WSFSQZdIk9LqP740IbqziWF7oODoOGsBrrEA8wXNfxlCB1Synfr7lD
GWxyh+L8/l5y2pl7L7CpMG6EHvH9mdItuzsY/VoBGtG+DgB8aUNnM+DLCKjK2pK6uYKHhRm8exI0
Iec2ZPXZEpoL3lFSFr/tO+y6tNo5fQ8bjGba+Zj4qnPOeP9I1hWsf/ifLnONQfH9zyB3zIv4RKfc
9Hk++8FsfGtdjuvQ6iR87NUxJw+5wxM5d5xmcNCx2QE5AWIrcWSQH24TmGRhjmlzBubf0A0WmwKZ
fqF3HbSCw3jkpBS/8fanqpAsPMFMNSSG65jPQjEJuI0gRKIDlIxF5Cj3HAUb/I1vi2vAt7hYFnWf
ftwrHYgggwcjk4NHhzjQ+RPs8Y+6rStWUFhFYx8HAEw9sOXcdEvjdsvCqSvMgUxWvvDvAlDR8HJ9
Nu3BKj6Jzzg9sQJboV9r+PqP8Jao19uJDDVTwWl7NcBYpbasMC4R6jeeeOa9PJAMZKWYxOAbDiyy
6vqE4p/ZL6ZytxDc4eCu7T98qo7wlR/PqP5SYJ8cFXvBIvX+txF/DZQqE8jjlzL+aA71E3oBdj+t
8LG7Z09DHjlBKWkFp+QDfou2x3wb8sM0eg5INhj0uCP2uc6sWQ2/Umbg0IbQxeVdArFBFBjyj9DF
P38v5PU/yxd1+R1FrXp3ZhYd3VhKFSZVjSi3mGi8LadgnL4uNlb2oOdmWGLtj6zjE8WOtc8S7f9U
fYruumRSyusIpqupnzuUGlLWhKEEnL3/gv4Oyx/gqQcICl4fAw1Qrzbdg/RQgAxuDQlzSIcO7O37
51dAObVbHpRTMGDffuzT633kc5QIRp8qMQjUcUjKKBIGv3rGrSdZbKT+/zmuTetPsOhvZLFqEhUx
ihGnqmqYr5V8+RrpGSmgrtd+ttntLqTyi/6BGZfrFHlMiQ40vX1gp/Nl0lnY+7enaEMB8BqYpyeD
RO6TKd+Ul3xNPzV05E6yTwDgtgTzuatfO+WjbQGfxnpwJvk+OJD+hriCUDl6a44RYuiwPhJix5+q
V/wpGG/hVcVYqa1mShbEUI5YXA36RoeFx/GH6mjn/SSnlXzye8CiMB2dBDCHU+vNS7X5XMQc//fY
yYxyKplbqwRj8CyDvpHeJw4cH0+8oTYWq5fMu2wTZY/bnz8C3Fv1gy/rxIJTNj6Jk/JXEASEgT1G
QIxGfMSLrv4d1aU/ZR95s8+PSJTc7Bmzmx8+lRIAyU1qgsqNDlrafR2QjXv/UckF9qU8vx5l3INW
QVe/Kf30Uv2W8iBg+VHCGKvZs9yLxbp/JarblqfjFpZGVGHYZp4hPx9qqVpEaEan9s0TiR2Kvdgw
CUnQNnEQindT1fFYaGZjeFdxanFbvLkLOlPqpslgJ74/UDdFi1GIJKXI2xbITIjwVJizTaGdKUhw
XBVQysL1HsAZt5VmVfWxWCC6CswNe4aZBfQt8iScAw0330tFNQN7LFNXucfwoM2+xi8Se2W007Tm
7Zf9nXT11eYwd4SqBIqOmCdakp9AiwwuEsVF0CLJ2hizaw+TE8yJYVcaTCGKCGtmguqUutpeGQ/H
CqkWCA23tjEDN+d6cq4d8BctkyYZR6TBiY4h/kuhiL3HYZjvmOHmHxIm3T3ViUl/CkwKqtjUFJjR
HL04vau/DoVvI/sLAnuMFU+9dkmI1pQPpeNBaVTmgt2lNkaFHi7QYBwg68CYcBhZeSg1mZPMNTso
bykuvDbrfVDaVN2GwC595bYx91yOlZWkkT6gGC92ppb0JEpaznxO/ql1cjfgF3tKJSYLuCsXn7L+
RM7t5Inz+MRvPPy3+aBH4tGETs/Ed/J/jMxWUHHa+vCIhV3B2+7xpkdXb67dyxMhfyQewcxRYYP2
tP+TzXHzWyvIQaTLunQr/1cZtKgDZlIhjVj0R/bCoIY3tmGc8OMPq/SnmdKko00xUptWwQoGmXk/
65eaRqP7FjYLgrplLnWnUMnjga8RADhmLSCwYJIU8NAu9Bb5VT8pBnZOVpQExMfspha2dV6HccTg
q0X9l0yNDhnwnyMRxuUKJ8cU/6TAJlcUzo3OA/CfCSambMmxtYVMf5MAXHE8uPWSWaxYNvfOxrqt
36n6Oqe3r2BRpBEbpK1mynIBkOeXy930BB8q79MDnEoBDMEHUMsdzHmYdKe5/POXkNxX0Ob2tPYF
PFFjtFOSTnUJaf2isN/rNrtBpHexo7JGjm1vDm/Wnytv83GGYO8N/ek8L+W4eT3ZyFHdK20H3Bum
D4leQd7/Nnj+jKvJcqOJ3ulVbyrup+BR9VHdIjQCbpzy0D80IgfmUqEGZRnlHl/jo/2uCd+YKtk1
yqmBc4nUvdpAvJrYprSUhKm4wMcnULQJ0D6WVY9vsWK2AaZ9QmaK8fPUsA0cLPMknU8qPJjzHjaY
QFWrThgpA9LyLP+4ifPpGuTfeQ3Syu1dnyLvI3UVV1CUWoPGutwMd/K8haQ5fr7GnJwtUiVlz1pJ
xKCg8MfZwdPTHPtQdhyY+cRy7GgBVOwjf7Iw27+TFbSwFbs/pmiZH8i6tgdj6ik88mPz6EyITU6d
/jwZB0mYo95cnpxxGd3UwtlAe3mhIPly8ztSLIlOMJsSJIwoHbkGKs5jbTXNggRKrFp5f5OqNx63
mmhor4zzZR87DtfiZlrIAojglxCdfdMWRFh3FCNWYbjDqU7xo6/r0TQ06jwUx1RFqfD7XggJOjiY
lA1h90nRzfsLVz79eEqBaatKcvftCifhB7M/nud876qIXoFuTf4DXn8NQzxH5NjoYloa2uARJ7U+
JP6vF6MG3DiPWrC1vjmdotPux1gVtwGL6mj+nikqfWKwtri3kIUanIeMfe1im6Nk3IIPuW6TVgMa
unb9NI0vheHqr2nI2QU27VYLG34DW/lzVlRLIFFeTApRzIfXbSUSYxxCMmdYwPJPl5jOwkE5K6o5
zrDqhnGIKasRRn2Vi+gl+fTA8Uz+PHd9iqkJdEq17daPiqGkZAG2LQC/mQeST8jcVP/FmgcRbYuY
0NsKb09/gTqcVKhtMX7Jd1SwSpZfNqjv+LJyPog47Dn/kcyAuS8f3lrd7bDqeptddv+54vvK3/Vz
eFZJWNcmpNxDBuMBiCRZCgLIM8keYiP3hK6Cz2UAG2tX7kfI2ahsR3c2jUXC/C3SFRRH+khLMmu5
vsz5rSHxS1HVk/A5/GFz+mcShDNGfI7xEkUvOcOvZU9ziGpJa4ye7h0196N0iXrYLSJDjB1Btj94
pHM0XYFHTETYTvxrUWMjKpcByT+JqjpC4vohst45fotEeMU=
`protect end_protected

