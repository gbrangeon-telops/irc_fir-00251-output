

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
XHCjR0nUvMBgM1clzO9mSr8YEx9qhDtoXdaphp+J1JlsC9lSFtsV1/eTy/jaNsyBimTHmHB4CLra
VqfCr1I3uA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ebEJK3bmI2t+WsBGbhWIt2XB+F+QW56z7Xo7/vGiNjxPbaq48cjkY2KIIwhppzuYFDUdRDxp9Iva
RlWujqNPGUrxJ1F5Pa0zN6dEMkhKPrWWxZpAFto5e5cB6DM88tJus2O1hLy9PRfKWKn8u2fBqIhs
zvXwIEX3Rz7kU3GI+Wg=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
oZLpbXnbPC0EfiuqzOyPqmT4FdlvB20VtdO3P1fZux3uAWynrmGeEUk81RKG8dIjeHdSPnugG+6c
jKeGIJZZbH6MRScqnz2QBuupQkeYWE+dCLOq6/P5LV7F5481QZZ3bx28u0vHGlRYhLiMW8KnJ8Xs
JLZ2IP5YULE4cFTCCV3WAM+IdulnwSP3p8oyM0uQffeAJkOTKR9dl0lslKFBplzuTZ7EnXSmYYXA
x4iYEfwbmUZvdla6dJXCCjtKnKqL5vI4L1nHOaep2f0bW/K78py/TJVV+vsvE7+Fi81aNwDFBE3d
V+IzN5VNKD8wM+OpLL9AD+xsAbJ5JCLz2sqFWg==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
YaruXmtmo/2yQOaZLp6UQc/TTak5F2uchK3/c4SsORqNnQQMwFmjpORZM2++MrgqzkHH5KHH+0SE
PP+ha/JFKIuufLvaAIVDYgMKSDFaxIIvD/8aIAhw7TgTE10+TXTruuPFiw9U65VaBnD/nSEGkP+6
2M+aqBTG/2UNkEELi0I=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
SWJkuOmi8gVneMbAS0rfK4gI+24fr/0jQv+b5sUWbuvKyCco423EdTDwW7ROH+M/MaGP2QTzNz1B
sh1p0mypy290KKaGmvaZfJU7NOmSNGAsA7Eq3zQGPHDW45/4GXnri5xLLNnybO7r0Ndv34V/fxH0
f64f4NRroCys3EmRDJeCh0D+WDA98E/EHP+OtfmYOGeO+CDzxS2m3FIcGKs7pkeR5dgt+S6srqxz
96yb5/UwV2cpnC9ULYZHZVQa9WYc/XM+Dk71YUYpaEFd7osc9zT0azChQq+XAkJsqukhufRg3dQK
YVPZotO8blEly5GYlPFGnRW13eEh9DRYsb0pSQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 13296)
`protect data_block
I2m0LaAAa7yQCqHr1iMG5E1Hgue63hftPYOIlZ+cxfZfXP+LwuaK2/X9LLv3efA9GlKo7dDxwLHs
/Bwc9G3xcIZMbnWX4BcsjjhzDx9hRzTbuufu6vdhqN01vxZNTkF51DwbGHnghxRCfQEfsW/NUMty
t4Qy1mwOsrx3eYGvFfjpw0w0oispxFtZ5gBRcgl/6Qalywqzl+ySgMoVqiGDxI9aA03xSZwVL/gz
nQciLZ4cssN/w5719kyLlED/F3hVx4txN9Rk8LI7+Xm4tEb6MQhjWH/B/1yOb1jLXMeoA0DPzzSZ
NnLdglp/74Zu73TwSwVM9fDuZeBjQPlW/1YM/zxmIGkav9+jZK3fcYJGH1/K508tc5ukRR3fRjIl
T4HaTE4BxNIDRjFnNBc5iNaeoX8fKrgFfKq/Po0hluLclDaxmTiifc2wop0p/G61Hx9Rv3jUZua0
lp++hvNrWcqlYf1ctIiPSH5H1/EoRdins+rMAn2OPbQ42dw2Ui4z3lTZfRQu/dj7NpN/RgxYL72W
gldCjqkFrJyeBjq/9VIOkyoJ987dUjSqM3khXSwuU5LdH0sY7L2JkpYojN1rrteT9+N0XEFPlUzN
xQWOcfS1A17jZa0Rur5qfq5bMiPv8W/vMxwn1T8yILH5iEntlDV7LqYu47SBk1jbRhc6dm2VYBMI
BtA2evWks5Od0KY0+a6Kw+enxR4BZ8webzVe9itpJcuAcNz624eSbAHLXxcwqo+/nfgg1rEXUrEA
KJQZAkuLOzfK6l9ZgHwqSL1ofjzsPJQpoUAW7LmMkt4/vFmqMdPEbgLblpvKsQxeE0K+DGES58S1
4ALqaRaqjPBwT45rRJqqt8d/lWli+526e/lY+dg3EP3owX9OiF3Ubg8G7AtH6YUhJRoCn1v3E1Hr
n9Xp8aibqUEHWbQ1FMfjr70uL1TLEiqJiqL+1meToVHRmsukrwg5ot/9a1LZEK2Fn5getHddQEYL
G4VA69Yu51/PnhoAfjUMxFRBjLGsBX6QpZZdZp9z0593+x2EeBns9TXIktAWguo3Ld7tUnJgciIQ
bmiYl3AXjd9Sa6t6OjTEwSlWqKjYVJCVTDhyDaM97CK/1NU8qXwwKu/fcL6lN5RwIDcLvVoMEXoD
VjC5uJ3Zt1AWoiXcgYx1YrEALbQeFKJDGm1FMPSW2EGEkSGEbVmZUFQiuu7La2mfkorfSAHFSoE9
LnC/Y0chk58RWh1H+tulBfsKgpyrK9UQigzKgKC4AT99/LNKsfLmAeDWBSGvYuq6S2FEUFMUTeaf
3qjejvcxERLz5hYUZ3l28BlLXum23KVpnEzcp3i+B0FISWQphybF99e7Y678xTTWHavZCTt0E3L7
DmpDgtkaUaip83Ug85v/2zlH4VMoiUPNLZMSDScPfaEdrNGZi1i5UwS8nzG/mIoaUsOGPoPzqJ/X
ra4op+82uEXo79lnXBlZ1yCRz4T8YCkOCR2pQE9bV5hoPaTM0kmz9YavXUXHIn1fNpJ0PAGxQVhZ
9TlIZO0sSqPen/bM+dyF+2cYsIAb6ml/SYoEHmIrs8P/tTLbalHlAJGEhNHTavHYcMs9ZNc83uEZ
M42zyDYCHZ4yR9GyYP9w7wNmxoHazhwNPUN8jUR/MzJQ9oqC7uMqXzRc3R8QCNcMcqfVGlxIbUTP
JMXhRe4N8MuaqU9aAUSl0iNZbDNDDuP9kYrRxarWoGOTNPpdCyNQXBiFKoiN046L3E+Ddez6SSf5
w+Y/wQiASHFGKelYCOMJxSR6dH1ri9W0Yg8oUFTU2J6Y9IFpyYvnZ4fKjMGYjnO0ybfYE1VPyQpg
bSS/JqvC5d0jB3UHnbjj24In8Vk5CKCLNZtdFm1gocxcmSBaubxqs//wmYAxzdaz13E2BieEc99s
eJNyokrLs72TX+uwGzj51s7ahioym9yEruIcC5ty2v+q39QENBc/2EkVV3l0msngfVi+HwIbf7B9
A9LXWn2O2ZrbAXbCw4gBpz59LPC673Gqq0aQseLInF8Tf4Qx6ilLEwj/o9ycqE6UDfsCOvr0CUxY
x896oRnuSiXGdOBxBN8ACcFF1l6FOyOPDerjRVG8JruoUVTjMVmSnM/5BB0+vM9NX1CcmPM5aFMp
lyc3QA8NMWp75TzCqIZENa7Bp/PnJTm2YSrO/bahoLPd1I/u1d1FOPr9Uvy815glb/5g1yeb12IE
G0PhlcFv9pJoDc8rCBbXbWrj6mAmsAjxNAVX2jo1dNVdjHgxuALRtxvkGuRH6WJILyxx7ZlC/eTe
PxbQRTR0acQoWvJbnAGSP8g9zF205R682relmoCiF5SWCbfb2HNsQZ51XBG1UVcUfqKd2sHC1wVH
mmTyJ9d583gmHlEuv0fhQtjKOYKoaLZ/aqjkN8bFS7RjVSoPGfBFoMNezCOA9/1nc3EvudUT6ROv
9tm3+eb7KVnVPJXiHjJBil/egGt3dwy/SDikGMljvtiQM9mxaI8/ttqG6PgLSTOQMhhTt4qd9H47
igrbC7S4Bvk4wuc/65JH8+hwTKeRnVrt7h733XQ033U2nAdjvAjTquFZphVZrCK2pmg4g5qejfs8
jXNOdaie10t/IxzeBcvZDbKYrXL41cdlMJ119JXaZeAJG9+bHpcWXEBlZVfEfl3payNL7rmVydFH
9UyIfqnNj3Y5zxjNEz5ZV1XcWpn75NUP8IRZxNqVC2I3F0aZkmSZ9fjMUPq4ek1MtmrAx+kfMoBb
fbg6AWFlSh/2lJoiTMyqOZgS5UcFA1tT1yK5EZIAZ7jpVHJpyJZf7Jo5sK/XqYw27C78/ww7jtqu
/5qg7fOy44q1ZuBYwYuhJScb2Wh5ibtZw5FFQgis7ayQk/Psw0aKkZB+VbJCgyfxeAJp9GADZdGP
Vzr3l7zL2lX92j/bLgyIdUXq2q6MjY30g1Q/M46TYsOaUGF7oReuQ0K9cOdSZo8HGuZNniSr8iIL
VfKGYgkY0PrhpOfvzxqn3pYmYUAf+dT3UJb1pz42Pn1rv7bv4Xmn6WsyAyvge5y0B1tvtooUrSAu
Wv77BHGXhWxhjWDIz/Sw+y0TZIPzrd9m5Qd2C7qS1c/owFlyrmzu7tRcG68XphQ3U4CrynFHGpQO
P+oMVaGwScD0L/KOBKCvZvn+XgGo0rGxF4YKwXNUibD1QiB0Xspwfvpyix7YZ7Pwx31LJ/lUn0O1
BvY61um4AVcZCgUZhPX6GpqY4EZlcKCmbLK2TSj5iQEr+F+ULXdsDpxtSh9Nb96TzcRdVyGr3Zog
anXbJ4D0ljHTeI99JyKQDX43Q+JX+/axg/eItZm95Dhx//lsHNHZp29kSa9gTfrkzoztoozWrTyC
9YhROz9Y45U7jghoZ8BSA0r8vwko4VMeNSI+bYO2/i6LY/rqyqEmMGUZafc+4leZcsPhzSzala/z
k+3b4zLn/JTq5N4RgbUY+a0TsnTRyYQghRzls68zDtqg+gv5uL15HjRNk9ay3vnWn2npg+GDFnd8
1aNurWBeRetEJ7Iwu8UIR7fwTdPrTy9zzrDJ0oga4qa9SaEQJbj4uzo23zWNZu+8dF6oKGGG+e3b
QC1k2GvZFHe9qMIGBYOfWyV/n/ySsOz5n+yiNUU5Ad9qwY/uxqpJREsrIu1hAX2D9FRiJ7NGLrpJ
gz9kstt4llBm6jbfsRkLt5YmX3hu2Ia3TcS1yg1D1MARIWzRFjRjXkz/8nYJssw1HATeyYT8frAM
5iseAlvqZP2FbMmdSmFz/u9IMK07Vdcy/JPqIUJA2sWmFfTwdWQuiinYvRvHcAD2/JJrQ1dhGj1D
advUZI50F69tBGxwomQuLvVtAs1UeLGcAoPIhNLMHe96JAfJwzOyvcZ03B97motN3Bg0qtFsMXBG
jMJ4kvt0/k1P3t5G1VwzsjXrLXOD917q51aOp4PrLeEGks3RwjP2Rfkv02ndsV0mFZ3l4cwAVDUd
2rPWTWWn2m1b86xpkj4u/q+MkIBGCQy9wXAuMJ8mZ+2INpyMuziIT3AoJULj7TE53/L7ottmNpl2
fLq5kYISpbH3rzi0YN9Ys3yW1oFEfRKc2XnulNIUjMDq0HyOJqv+jDpWGWUnTdF7kPNE+bTGIOZ4
9GwAO3V46idaLozeqwnm3JrKE8YcLLlAhTqDMu46Tp6TrTHodMJFBbIb0lFN3djQg7sqoyKG3aG1
2Wj+Z/rcH3KqCfeSZ7AhM7OR2EfRYOoAGYrCkGzCGiKDUL/fdDu2ZTPMtJY9JZVpwTuKPO4xAvel
nZsNnM7Qe8lxennOn+pyUA3SiVZJ2wCm671ZicRd+npGCmXiOsCtw+0owUGSiYujW1J8q1EDoy/j
OFVHenIFzg1wKEtzyIbCzmFBggymCiLr8c8sAFNHPCSMqIGw8Cqag3MLqxa5lNKfHG5KWbUKVGIf
RBTF4RpDz0CurmEPYsJuAmeJn07Zt7mglnu9eFHCxI8G3S8FnbwjZQXeU3PvdOGu1dE8T0jhMGPu
1a8zvNVbAMdJQ1tg4/0EGt9iBXy584twETGZsnARaFdgvniM3l3dxKRvvluul5O/D0HKELAXWS4P
pha9biKcdco+RnMsMKZZLxWoXuRVnMQrG8g2TB+80jbeJm99rFipIt6po4JYLOJ/7cVUr0LHv8nL
4m/6/B3IjsHSRpfSykgqbHB56clPbdT28QIHdaetqVN6eMAqmEUZmRILDCzM8+AtCOueRu+ZIu3z
W/sN+Y2Ujh5ukE16V1FttchxQGAZqwKz4VKYPOfXV0LmNMBQm4Fy5XW75URAD4WgkT5KQ1lpetco
c49jT/xXUmzuIUSRylicH2n3IbsJZc4xwQ2w3+QnePIDN8qurbxubck/TaLUIIOmIbsUuIq24mWn
m9E9yDpYc9szMUeK077xwT5qyuAhBck6ktinGi13zYXhH99Fel7ItpeV+3m44m2skm1ENBHFRnae
I84TORHbM76s9sX/ckcxotaKMh9T5I6yejbMNhgvLwyYmzsDnOLk/X8S9xSrwW8qqxoEEtJTMdXP
KdzGJvW0/A3ZY8o9jtJiLaf4+t1h2iDd25Auf6e4DvaG+mcQ21hXIaF8qQ6SZ7+i+qP+oAxJo142
nnZxeeNePNeJMafhU2mm0xa1xuYQLQACM4v73osW3Gx9O2o7iM5qrOQhHaaOihKqx0mTcAmNGGX2
xYaKV/bfnUqg4O5yVdFNlAADbZhtm4fdZvGcpPBYmHoA6Fy4Joz7a4peww+Ja7n3a8GgFnNGv+sM
FUVFKKEOn+/pYHCwG9yMvDvGlGKf/4SSbR+AcqaB0aujNUyrlI58dR4ITsaDMUIBPNHqxpniY5UT
6k47eY+PsCicnZmNbaHhpc7QWqqlzJvop3EcutHE5WrIaxFDH1rSb+4bUi+DfsuDb2dWoVCi4f0e
4dV5KtQYF5W8CJMinniw1TclEOHSy35eZR27R3sza1kpTreBUT07UYNhU/23lcV22GxRjSDQ1BsG
MWzJQOaOZ1g1RfFDuexNEXT/IB7ImErW1YYBpKhAMHqQbHEEZDA9fMA7qRBaMAh1DiuFlSS1+l9S
ONjXbTxG9GbkH1J/B2b6XCU2bbDleNqm+hEmBp+h/PxrGnW+PORQu7xdh8bFV55aYx5yLU+WdRyK
/8WP5Xah9SGh8Zgq4Si25PohNX+I33EDF4uqtwHA2WwU3oxosSRsSk1xG0KeDaqHNWhApFGZEa3D
qpUuLDe0xbtwk5jr+DXYAk0cE9KHsB0+sarJW8WFEcAx5oAOb+HIWhrxK2RcYSXaUCn5vDIfBz7R
ifSM2AA88X6OritOzECah0tyi3cYDPVMIt191U/logPx0adVg1b3xh7G7v5whigg/bjwiq0X5DUF
1mYt+tVr58CQ/tiQcJm5rIoiUlSbgLeVGh717Kj3cv2EvsuDTDZ3EVSA/gq8V62mhDbdlfif9HYz
Gy5EnjCM8j3I2uiOyfCMpgU94rYrQv+tUV8u+R3OmZQ9FO4u1HuYlUJ/ig8LGTJt8FzJOSoJspQ3
eb2BA7kxQd6AI5ucP9Oq/3lYNfGGXorAb+zGcvs0NDG3Q6jcjGYinxomcgFQpi9bYduZQs7erDFy
TeO+rqK6AdFmorGBCc1oYVnAyacG+8GPg4OKSAtYpXie/B/JTFlXz/QsEgvZiFYejTFNO/shhwiY
6KWu4Yg0dXWDnUSVXLiRncUNK96p7Jt79jRUxEEZ/CzF/MVHqhTM0Uf7aocDrBSPuuzIYbgnGeda
ivxt9M6Dj3zwHPkNKI9Ch0ergpv8Z5KeEFZtPK6WjpGCjdQpWs4moynNY+h4REie6xUGmLcpR8H6
YaEbwWYgl7XgFl4ehzVtFV+9iSL1jezqKCxCpNQ7fzKX8uY/lDV/oWzyfIbuvSOf1yAsXNbDCKQC
+SgpcQW8foI7dOaM/MjvJHauEOorKqa0drXX0eCiYDrEUVW0Gzy4dFVZ63E5p8iq48OxtxpA8Wgb
H9BAaZBhMOoT7Pvod644E6yOlHBTrNOA9YpiGPAMLIKqrihMjgDmAx/U3L2H3wc0CAJtW1xmbG4i
eYknVVTNBvLJxR63cVhvF2s0fJlVcLVxnthDVr0TNar6oOu7n4g76ZUzR3c9eHU5FgdEXQujyoJS
Sy8oaDLNixAz7R6AEItYmn+nEH0S30Ohn8tt9nGYnV1dsIP3vwlTZeHkg0m5rcfEu9CehmG8CkX+
7WEWx3tG/U3gPPgAMaludabaYXSlYRWwUkzi5CaZhEjzn3MUO86fm6hTeMYStqzDTCjs3gvbHdBM
W3hTFzYK4zeQW5YryhcC+6M4zWKwFdi8bKZFAtiNrHH6cbw2Gaz/l1X51OSn1uYEKJLpruh5ANlR
RHPGH2byC8/rWmkCfHypmzLS+7K8EG9lNfaYPFyfjiNlx29pZ2uv7ldhQAuGhHcS9Fc9CxJYhPYv
BvlWUtLOZhVRNUy0NnnqOMQGvj7sm019D5VDI2crXYEvmjZsgu4wqILM9GEeP4kiKWwRg+M8Lemf
TIDCqE1wXX+FwT+4+cHzOCFFhBJzqheW9dtwvojZLPHdbMXTFfDOw2FGCLDcLBDCrg8FAY6cF22n
+3tamEoL0j5f8V26o1Ftuxtocn5K/7wjYOKhrADlb6R2dkX6OlL7qRbrDDVBABVxSz5S3MgZuTfJ
ad8qkNjKoOEkaOFa+zGVho/S0QVrgL5vYfwPDF61NBWkHdAedeKrUkmL1RjMMn2ajZHsxhKGMHZJ
xDXh7zJP2TUO3IrIek58HetLm+ck0ViMuAubhuanov47jD8mzfD9aA2k8cuurSc5dlzLL5gdCAld
2nHgaGCqeP62oDZYDsgFFFlPNfgcwS6iAFVOej3rm+G5vLdJLJfmbPjoS4Jz5Sij7cSSG54E7jXG
nxDDJy3mu8W1uY5agixkwr/nRYhuAlTWbH+pr0AJBvngH8F+ef8Fhf4kFzArjPfNVtGKak2oLCO8
CPTLpz9uNxJDnjNWD7VEdqH4bcN3oVJYhTvOOT8k6yGxKLEWpLbIqJtI4MNF3ZqQWuhUQ4nInJ8D
f0qqAyzXZyZn7A1Vm5tbL1m8XpPiI8rxz8ETZSph6ODWYs2CiTh/OOMontLj7LiKhBMLVl4NN2oA
utLk/D9phBT7C5WmSXKImzTEC7z2P3ZJfceDFxc7O7boV5OhkEl0ayxnvrKHR8yH8Glu0P0mlHaa
lEop80+gMDdHEPSWgnB1RFoeA83ulcCHBeMK/ot+12pUgHHxsd7tSjvJU6lcMiX61SreuINq2aSK
pfhlt1BEIcnvIcqWvy1/c6FyB374RcasTinEGmaUEiL2f2Z7rqH1krKQjeSioSDoKUomUcpqDbth
CKrXJLnvzo2aCkzno+LQ89/d+Tey1uzEzt1Wqs8cHHEphCZNNsDYtgvuEZqxYaYYUh56UoxY7xz8
QMEQsHFUOLr7ifLQ8H1XJCF57XmpizMbJjavhvAIW13L9YktkLSAS/fhoGI5t3bK1i1Aavt1GQJx
yhMAGD3MSD4hOngn6DkcLMlzoaNhIGiInvfGQ/+v6AjUgu0MrZleqlm76d1kA710ftaidPyuhFiD
pe2nqket9HVbM2/L5/u+hrCTUvfZBnjzgXjXP6U3YZdcsyWZnrT0jI8xUTaeYHO02r0I2iqBp5It
fRfRLVQy9Axn/u064ogxle5jwgh9pX5qoTZDyfnSO/T5ex9m9Unp5VMvDiHJu3fQl0AgqWeu+m6U
MK7u4OrPTBFH/yrxfJuNukcGQdQM2YL/Sj/3E0Py4SaToIRXYU62BZOPEQ5vBxV6sMvVNC8ufwd5
sOKzgHyroDYPO+kRc8fZopaHyNmQ2XvekfIQ8NR1ZAa15P1JY9zNefOHbt3jiL5FuoTVwbFS6nRe
yMFZOA9QOg9tX9fm2G+wHp5nuX1L3d6fIeKUZ16RY+15Flf/ENKggFTseKGmyaCluvVBHefSYlkn
SPGk3pc1nOe2BTZ60ix4po1x75ksP6QC8/MY+xAJO4fqtAuTIMr43iptbdTsjM63rUc4V8qppgss
q6ib4+hGKUkXuWtms+9Cs4Xnf+Kec9RGi2+z3q7oFAezoazwFEtDyKpY6crBwN2nFwVPqpk2GLbp
UOMS/7ZozsZA4VMBGaaXENCTI0hPSyA+4o4btEiMipX2JWRdjLMfm6nkPZBlu+EvCGNvdF3t4d4l
Yx/nsD6KISrjmoe9vERZ6ssOXQiW2xVY1HnKDanOLsz8MB4ZvL2Jf9xYz6I9oswpOZ/fiMxLySoQ
ub66LR4LjRsgQOyICmjUdjenNs6e+wHrk4bv4q32X1srUs8qa1Gu2r5V0hi/n3x++EOlSpUkofNG
oWF9unYPDLvtAGeTrjUU0BY0ze7oh6DA7w19l+Ylv1is5J90VrdUhLePDzt8JXL7EkshFa3xRiWw
bbonI/+fyEYjbIIb4Hi7kYDnv1fzzeFGpYYGW93IsViAZmi7I4Be579PSW+D6/xWS3z3taC/bZUa
/SldVojHDrxPJcv3DZETKp7CsbRrZgGCzWed+ns7ZNy1XlQEu4ecxibLK2l+Yr8BkqgAo6kOX1qe
ow/r4BcsGQHnqc7CY6rS/c3xRqW9FJecp4f1XAK5ypsVH7/buL+ploO2lo3h37ehTjHblY6o7N6E
ckHTmqdedyopi4MgzDSx1ruvTGDwEE7wpH/6wKI0/N7No5tCp7JcK1IH7qu8oL2pJCqsXuhhu691
WN0CQ8W72pYingaBKMEwej/r3DXuxc6ndM4eCa6k44I9F/pH6n5dwqaJJpnXZEzuLr/lolz+s6dN
LfDHZE9O9GobfxkguBjMrCZYMrnaxWMXUY6ikpZ4gHhw/Q3gkBsrC8su3R3x+7bMwIUDa4jZ7g+/
hrLW1Mr/pujY8PgwNtl8hJKyOCTH/m/O+mewsgPV5qUDJBwKgA6LOrJmYsgbODaeEjphV5i89US4
BYZqCZekjBvxEktfkQ4Hrmjaa4CJHuDYfUIZC7qWRTdgCZ44zYFtYC5eERMTBcNkB35OqDAO4Nbn
+fFl7+IMZ3yqRBkxvkMCjbNllULeDTS4jhPZDRtQFD8CDZvLVUGdnc9RohaL4QPpQe3HIXtatxFs
+1VmQ/8qT7imaeaUMGjX5tk0RUR50dLsE01T1Yc8Cr7bZq9SPIhG11qFY8iONAP9nKKkrpBtuTy5
4QV/3U3CI2Q7nfy625xJ6J9OA9wPCegRe6metIS++soSdmap87xWyrVNv7eBdsRbUGm7sMsnzmXY
m+9V7yZjtZXoYtxW0gxAyjkGT83vYoW6DZFiUsCCq/JBEASoHtvmXhP/MhOD05nNJYNI2D7JsYPG
GmMbsXA0jSdqUCRreIqLyxaIwXwgD4e9TkU5yo81q7PHVbcWN0ldZkWVcw9c8W3PTNIBzYGibJzr
nuXNh/ZWAZJAIB+V2ky1MRaD1W4ZuLwm92545r5LIhidFE30wjOMrVqTtbq/ZM4Cnaon4zX9haz0
TJnOUM9pesVW0oPn9bk/VsuOl822Q+thA7+PoDK3ZgcJDlAiDl08vj0cg0dCUOXtZEmh41b0ZJW+
QH+ZlXx+ktdQ314AaczouWwTlcdEjOaXQ3W+MP5KnLpbWDo2r/5yMxCRByPCLzDlscJKjV818uRj
GlY/5HV9pnXb4uZWJrcFvUbh+ccfFCU5xgP+6LO2V5qJNjPokgjD+RE+adECdXnvu4H7jwKOKlbd
mxMpQM4krInvnvCb4NbowL3QVS6eceLJkLt8x62wBz/zXgDqHyiSfenNXnB1WhhN+X4797U5wAXq
6XEEDcHwjjGgGGD50wSD3pdLHvgabogRKemSvCdMowueT1ewCpuq7su1h5F+NiBlLKzCP+RxqVud
9VadzWH8lgAYSX2c5g/pWX/sr82zbrPh7w9X74kytfJcUxTA5z2+lw//FR0Ro8TEiXBgbGd35Rax
eAK9Sv04Q9xuLfGwHhHpxEyM+TCYeZSwSytQ2EDfycKEabSbG+ySRuoIzf/OCPpgGhMo9yvDu6xJ
fJTWbb7n7DKQ0BNdM0FIHyMgMSNBvPYPpcI1WLzS+8q8O76BeUSl6f8Tw8DstpW43rvpWSOvmxO3
ivXlp1mswCSWPayiSh5jZ/qW0cyW75i2L1pw1TntYdV3IJhyimKxtFx+lBmG+4uSpHZvPv9xzEYZ
JQWxL1p6zLs33VDdhuTTvNg6t0DUUx30neQ5chfRk0pM7eq3Mnt0cCrj1ssft6qmr1gXBK96ribU
pm89nymovwAF1ZNicUjExwtDf57B4EjkBvWOojfGnMASdofNqaE5bTSXiOqoBinzGEVas8wDIhqF
c+BDP+j01Q4v+2BKpWeC3Miqy96k8vUr/1IQvaTVctP+Kj6f27hF3GNa057nbQVW9hQ42Br0oPEc
sX/HyTNgGgTKa5766bO/vKsle/B+JYoiOZKy9iOHUoQQVohqWYzs2GHuqt4xcBEhGUhjt8vkBDZt
oJCC+REAa8YGBlVP0M+GzWCseHrDT0Vt+sH3kYQCrAeyZSF80+r/9yDEXNpF2tf/XP85c5FEdSiC
G5OGovw3Xyr18rJELEWsOTXhZ/KtvIJzSuoJDgjQfyQFEHTT5n4ZriAm2497I5aW58Pc06JI/cjG
ux0xvEoK62QANTJ3M054yj8NVyCuty3NwWLw3kHB26ATlNfCedYRnNyjKENSmJHh+p0nU0SLuS9P
KZsNwv3l6LAltXiJz5k2MOMbOZtAW1JowsLVHaL7u6OLXJfTjf+y/KwjT0UQeZpgqiroM1RIfaVn
y4kejYkefx4FOJXaqYilhLx4dl1330y6ecUHqKeyHldBWN+WDhvJGIpEA/4X0Kzw0zA8Wo7tnY5H
DpQkB/nwsT6IglAGXkh0hIDTipCB/RpSacYeekwGTdN/UTxAMMSnGCy0jJaudJ/5KgP9x0LKJEi6
8abQQbjV87CJBGDifyGsImbrEbDxQC9es296e2AI/5stzOE0Fk38zQKjJbk7/D+fv3sUlSxKEm3w
f4ElBkxg0IIHod74q+NBsFRHlppsoq869NsZ9sZSnD97ldBR0zkns/hCQiFJ+K4ogD7y8e7cKiMI
hU2/t321sHOhS9GTYcNCk71agVFJ3673VbHZ4ei7ixTAXi8FQbV4uZNBoGilKIES2APw/Crq1DNQ
4Av1lMQedWECJDRsXfBW9SSRaCfOb98AHLTd5Fms535KWjvWaYeiyYLkxsWDpj2k6YkphYL/x8u1
hqhNGefiNNJ+yV4eE9+9j3xrMrbpSgjkwYTfuBKOI8eLpu8QP/Wdv5CkC/ywCTGDXoEEDH/oLSYq
zysmG6X5oW5U8hzJCx649N8HpdBoQNWLE1cQ9CZFlYAJEhh7+Vot3aPHWM7D7r80bafuBWJMj+CC
Qia+3crc8zd4E09He4y/2cg009mkrkvZqIsS/YtV9QctwvJBSwgozGRwEY5H1qNVZNOpL3ncQ51q
Uo+kl6kfOqXfrAiCkPFOl2qA89Lyagkd40estmfEF5+cepcH9jGfJVBXtqJ13aRcA4LvYrD2VG8n
qJIRVJgfZPpcgjqa/u7m6h+RX61bDKn+t8eiZFn+lcYmHfX7dICNT0ufuQ7lBrZoutd1v7vXzru0
2rosbn2nyXgxg/kC52YDKAc0BIRqOSCabmMz0Q+iqbvPas68A3Y84KYXItXkkSjGx4jEma0HZFPA
0ZtlpSNSfp748581ifR1wwMciwashC17DzXxTIX86UXwdYtfxpu2DN9PvEONd1Gr3CbJY1Y7K8po
0h0JUC4tAWr9LfT1NSH/WwMJuNrK83RUIkqUgHVKyv9g7jHhbvcNKaN4wvaeyxgFQ/+PEkgMTyMp
hvwEwQqCLBFh9ZD82zDv1T+WPm4fYtcUIVX63iI5jnH7dVMlHoZouKmtjU3cNg5dDdMLO4SH7pfl
DE/aITslEjpBXE4/u0GkBIXIb6I+piFMCO73VfT/J7o0gbnvXJSlt0GMOPQLHy192Z549Zp9oNnO
b7S86CcOuE7LNOJB6ZbxDrcEbfO0XdWmNX9VsfbgbX+b7ZCZUROi9lqK36yF0gEic93g1YiJyY9Y
seyQ9WuJbxOZ5T9fpW5edVtBRmViUWrxAcP+Ycu5BiRtUF9z+KENY8iEiGPq/IoRCB8FQt4RkCwb
OlyRLh2M6JQOgvwkJ8D3a6GpiAwbeNGz5niXPgEU6pmiL8+i05BXLj13St9COK75eQ/awdy5JdKe
a5lWEL9SEMNSGVMznjE8rusHxr5za6SVKzJbDBc38/jWxaiZH5q03VXz4Fb4q0cx/MKRFcS9/XhQ
ZL3AxW/BrQBB53zTbXtnAOjkIvIXyrzN+pnhxVJryW94bdlmXVWlIkNwDYpXOIfqEx+IVpJhB+6w
7FpDMK7dGQZjQUwmBN0wuTRrY/8l3NluTOuQPk/Ll4ndfLrJHRlU4JxoCF8T+/ODV+vfDu0f/sZi
kOuRuKyid0Y90Ke9OgtkA+vlikr9klOaUlEMQulxaKCGGiSZAiffQOuwkEnTuJxVT94euI3f+qqj
VwFkhR2HmzpltNd1RdiGuovKhzJb2sKcwSfQo9hm8czhE9Kpnb+hItchR7T4z7T7N5/yyiuEbtoD
yJ+5+ZRWZzBSsPzUMiDky22GFW91gql981tozaJCVlWj7p4zB9SNGuo3xpzepztl0johX2ExYUm7
/G4lbhD6O76gh45JNRdrYNR9LxR6RtF9W+F0/rDPTBIBDKCa2l1vB9FXHFpT7Ezm3C0G4G1lN4yC
arSvNJXBiqdsAsQP7MywWKLwaf2BIoOFta0AQaDrmfUyZQ4j9kdGQUy6X+GSvetqPhGnl+yXeSIo
sfKVmG5xeuf5PQMoI57NZfgceRmPwWY51IHQmCx6VbK9oa7V94XatNSP+VomXo/D3n8neRByZGBJ
jx2bkj86WFnNmQ7hr5aTGI5xKpM5SgMyzk9jHyKeSxIWvxJapcEzmXbV7h4skXzZ9ZglL4g1l9yq
7CNr3KYnqIDuEJmI9pOIbxWLBQ/X6cRM/nIgDFvFn+HThRyyUD5wqWIolI7DYgUFVgQnhTEezLIQ
I3gT9ElD2ZLBwE1a8ZtZGJpHiL+a93PfqaitrPEuhA5lmZhYJzeN/mTk1EG1rXrYLLdzKsHGlMUx
IHZyV5vqFavthEocasme9GzDVEKSWUl1aEEacdu5UnGznlNdsVqWgJ4+PGzTmrMHj0r9IMCGxBkD
4O3mGztkar9lj7HtDq+h4IBp2XEvyxEYpcdRFSMGh6xn64lvIs9yFdTnGlu+wk6zI//nwlXyBy6j
w/roBzECylTfYYo41Zd1f5GqR2SDYtjR8VdfAwvsOgpUbLfjncaAPOTrKZiweVG9mwHbme7Dpxos
/n+KormaqU4AMj5tKs8ANkrCwmsM5VUCgSMc2UpgESF7C/zrgKyxaNH5srbFSdu4kbO5nryPv+7z
5T5TGMK4Pt//BU4zHyZFiXETx00Ovf328CsHi/CCwX0YP6drbS/IW9OUxIx/McvpDjxIiU3yc2wv
jXNr6R0BoRhrm/4HxVTNv9V4DtfPGjvekGXqFYydLA0ma5cMT9RMKRwThzQWwkcaA8pfuN9jxsT3
nTfvuCOG496SUJF9RKLAyvDJe4JKpb1taiB3GsLsmudTtrjuNLwsEzH3TxxzshWYTY9cA+Wz/G1U
oe7SNbpzX7pBq3kFtw/CZGnaUO7XkNnheJzNyuhvYzTol1xNXgn3zGJFrxiNAlK2pViMoeOFc1KD
VJHbpiGqnPMX1KtnCN2oTvhGV1e5YaD0/04qg4OMFI3LdRh8zmp7k6j0npTCa2h2VKAxGAPDPlrx
fHiLjTPyi36iYmphcWWyL/J6Bn4IzCFjOF3y5Dpzj6pMR+dMWDxKbOFtgoLQQAlxKoLJzqFkXvr5
Y+wyqWZ/o+UlFDlo9JhFtBpwbAC9EDylEDJ2ZtTS+NPhNMxUR9OLIe+wt57EK2LoVGbCMMQ6w7xe
c9ttDpD/x2AFbGlFGBtbOq9LxhgUBBKdKx29KkejKcJGsUZLBBppILv18pl4NIwqCJ7zdjCcRFRm
oWZrGiv33HnbwcOCDGUztuv/ZycBYlBM+RNhqjHEBqyXvpbR6TFmPrPY7coXulDAuWxXUZAnb46D
w+7kawj6+rtdBIelOmvwXY57N+9JuNC+sxVkhcdtqB2BWojiEr+eK8/7FVMKYEdb3+RO4jRYfxdZ
78nYAiVtgAfMgTlSYWszMi4rWlFWbyRuHHYFeWSgNTfhxlpkIBqqKGElX5FHpR+SKgYTxLkFY5hw
dhoc/BJc4q+FUj4pd4TVZo1SRRgLHXa1q4j14YHKhzoCINeobfkAe5O1hwmxlL3kHXSr+6MM5h0K
Tk1cv5FVmwOT8+VktNdidbrawTdL7lLbOVxl8zk95GHSfkE7QZbsJwJc0KMl7OYei30HIfwBu3te
8TQjL8prgZbRBhR1NrQt9Dr9iVZVXtge/S5O8nrixtM4pt+NE0HxJr3R4dVjrhK/0DniN/Oiu+wI
PwIHGuWLcYCIHaAWJw8poRWVGHZqAq6HomKrhZGOfhMMojWvl9bOACZw6ZXEUoPoLM1JF0tUlZWm
QVyG1vRjko3M58J9U+cXcZuBR9yzAc/4J9UAYcM1hufcCHvQqpwjn2DK865Pbs12Q78l9fw2PQty
BkP6YPIC8NGqPHTOslxayPBpe/XMVh4rFyTxPoE2C/uaFFFG/OTlO1IsRonZcv/04dRX/QdJD8Gr
+ZIFv4knXp0gMmtLMEjlLGVHi7j832XL7uR/XB/PN4R2ne+/maacN2f78ttkYaGmNUcLPtPdEGvA
fvIMWvH8RRtG6GRJ1ifYp64nI33xRefh0wAxhY6qzxq7n0haLmgivTrAJJfFS7Xm5fIQmrUcSeTU
bH6pewP8iJ/+knCey9HWYU+jm0LcfeLTzqxEhfl4YKC0/DYmqCdjIcSbE0r4SndBMWMyfvgKqrEW
NtQRCUpXOfSmuUUoio8D/KLgvVgmFKqIf2i3nqyCMWK3AEbY/c0kxgemmpog3aH/wrKtjfAimCVr
NmMRzNUdbqqfn3GjxPUOdQiwobRL/42+M7DfL47v3oLfsf9ak4194n8GICbPFR7xE6R0zj7G34pL
5MQtjC0EkiviImQMu30o54oFBw9s8IKrETPEUqsmF8XQtL6LjPy4HxTAI0bkeIXjamPNmdbSpFsq
x8ju1DoDUaVSFqH3wQBSbNKEeBU0jEfgzMTmtszsEoJujts/KtNNnMXp0RYl4Uxrz1MF5H7r+tlQ
2xIoReqsOEzPhjWRiQa7wzO6/p78dNDPiUlgw63ew55XywG+tWT8Ji5b+V3qqq2pNm7T2GjxKNqB
STfWMGtWInwmlgRpTO5N1+hjWd8WXzh3/TUlaPb1vGnM76qL8XfbtDkO2vK9mYEnKylVZXATzKF9
cygkFS3ozKjLhHPtS/HEwGz9IPVBrIf08Thl9xPXgqRcbA7vkvioPAM/0W0wNhaUVdre/amS0LOO
16LDu2BLFc3Wvim7AHBhtsndyGBTY9fY8IN0NGQHwPLFKvgHPFQreomHG/iLONUcFfKm7zw8dmLr
pd4HdgdikhZoqNQyXkToGcETv+q08DhrsO5EhHAuBEZcanGCpXggHA6+BidJLw5LE0ioDyjtmajr
h8Rwh1x5az9Yi7p9sL0m4bFr8JklUYTizI/8Yfo6kRzgwT/kUUGCuzSspIEwg4cCUtGjnxvzN0fP
b1ZiF3tTOneB26dO8jslEVSI8/iHfviOTJLz3o8dKnC6HXUvbLaXCsic8gOpQEnbVonXjvDixbI7
FyoSvxUl0uqCUN+qTZR6s0T1ywiQccdgROIzFk+50a1ZFur7ogtJpSNvh3+5L5iOG4kf4V/Jk5BI
gliQFZsOOL9hpHosPql//yySj/YzF4749ywz2s4TR70pFrWXjIRqP/b3M9/pAjcfmKqF/AyFKB8k
oxXu5yJXaawRxCnH0G3Am3y8DIAEHsIj1zwrhf3bb4d9W5tk4n75RgRqobk8RCwo7PR7BdkTfNnn
RbOfvVmTp37hF7w9ZWi5nI+0mrHzMpqomteXtrfBmPGLF4ccOhXa0vVsoBHj0M2PmWBnL0f4GCP+
oziewfOFCLJxCtyQsL5shuyjOa4bIfeQk8s6Yvop+yJzQg8E3GK8x+Not39cYIiLrZJyDJvreJBG
6Y/YxtPPoxkZJECMQIZO3Hr0DcrBO1AWmtpJO56+tjUGX+2dgWTT83y+IlDYX6WPOYEy9UeDmMQb
JpHv8JWNP19el1hwBuO0zOpamKAptSiUxoy2+wmIFhR2fJVghwpW/GZpYE1Go+AETJE/T81wPeXm
EthxG9YmkH8dgVz4IolHjCts0FUh5vHMQ4UomkLOSkC32FZszu33jsuTgkyLGlxsJpUQ5xQN1Gui
GmOfCL8GvyjbhICvV0Y/XJ2yOKI3gYyO0Wz39QITb77x/1qFcpB/pMwAoC+WQC+XuR6tl7Mozqjx
IFefN0JlQkFl7Vm1GZCUdCdHRDnJXckt55kNJfgRu+8thdlCjeiYOQsvzmYDOeInNiF593a7lbEz
2Z5t1Fu4dVu+kgFi+IZpC4Z6UXAB0lUVt6KxYGFr9lpxm+dXi1dwOr/vMpPFZ8ilTg2uD5OU8rmm
Tjd16En4k22MnLe4aKeJmbkgvi8jMSSND3HZGx2CC794PMv67uHIjZp9rNU/5yLvWP4aM+6QxLCt
kurP1UxFoyG9lHqH8G/AFd/Na3pKNVcSFXqXYvjCgSezkCvbnx9VUsUNe6kRCtbUKXU0XyhUTQyk
XhLWq8W/UqOrUhMf2tpwVoa+2dTI3jW7t5M3yFpgE7ACqa7mea58BHeQs8HR+CxobSznXIWLwpI8
asa42HhtbPU6IyxpGW7xUOLlyOYZqsbiETXGd14d3Vm94zwy26gdvPNc5JVUF/n5+YQztoDkBn3d
55cEnSh/LSENQC7LvKo/dHQ7Ko6ktq4nUzZeo7Pq1jr+gw91LeLgjKtUNSHly2Rjv5Wa1JbsWE62
gyrBLRBEYNejbs0f91kKzTGkYkc7/W5EqAjwKsIXfrzIEl4hwUybmvNbFNmnauuqbfpA2kLfKNuR
L8btO+6N7PL1a+5oROkW9O6z1uy0DQN4TYeOYrpPVfVoECmgsQ+aOjiNRLxuudxrOCtE/zypalB1
7FsScawik5ZhlWSpttt9BrIN5uNq55Gs+77kIgY6lyJW+3C0MZt9bYuhmJV6AsHun263P+EsXWTJ
95622v9w1NOzKu9ILFpv
`protect end_protected

