

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
hajT1eUvtcpbI2tr2ZpQ+yt3wRoxz10Ck0HI/Kzj20i705g6DeZcP+FvEeRZMeE3iSuhECQss2IC
TSZjW2KB+w==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
i/I1IeDYXVmyWoncZmW1nYLxm0OqNFHolb3NRcBcmjKOMCITsjC1Wrr+uKyOyNEAzg8LAt8SApGl
0BkTt3hGlwT5vH5JpMyxisp39DIoQ/2rHyhelRgIJSLTMOjHU/hpeFRg/8m17ioym3ZBfIcVRSy/
8YqL+H+Sd5EIN7orPrU=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ZwMv3uHNJwRn2Ww5TFfON6zTPNrPAlVNsMdpIyHdq6Uz+3GTAES373CyUHUP+cjDCtRwMjqRzGuk
B23rvW/CpivFPlGt/mLvn2R/n+PRdHgtaqKJEYqkidXp8VZscndj5Jsns7Mg2gtWutKvoptc7/8f
8ZVlv3hAdKdz/jYv3JFkYYsQYs/9EMmUObpsbPxhccaLaqAcMcp2DPumqvxQeqn7235qfdKNrMcr
c6uFXng8fnfR9emT//lppNqdkpAUWD93PhLZYTwVVXcjV4e16eyGLhyZTZ2QS7WZbPAkj35kG18o
nJcfgFC/GO+Ysd8/MvmMgbWhQocjtlk9D4Q++g==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
F+8QLMkCmxgohq3I7y+DAO2INd7sZ10O4AWi5yw/qOjlH+MDCzvNaVws6hhgvB6On1+CWzlrQ+vz
8M+w5LD4ga5aEaF2/H5jzH7q3vP0dvfZN4yRMhZ4TVDJv5PjxyVU6bHIlNhOrXl3MF1oGoVIjZ6h
IEpVBqdC2ShJgsN6O40=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Nc2OtpFQZFg8m9MEwwFrTSX7PqIQjLT0ImG8RPKmLuLlbhKyDcq1HH6KjYM6DTZXkQahd7sF4tka
CU4JtMixX4Y8KRzlmswh0FCLw/Aoh3nJlGD/KZ3QsZu5KBZUxKy0A3ntWjfTg1NNZ+tsdv0ZU17t
6SODHMUk49BioUo7eB0yCXF8PR27Zd7koQvLbFKTXZjGgj0ayut3GjrNM8A+4/o3G/elRT5WscCO
qhmVtlygfHoMk7BWSkupTlNlfF4owb4C7/AqdxneLzHPlGWymyNm6olzMM4lJP0A39+MtJZjtTaU
VxxrhX4xVaQG4Msik48gN+qH3ORiExl++4Wttw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 25536)
`protect data_block
COzlGUVjnl2p4Zg1rcG46ZmsrAFo/YKnV42MGKSqI61cJcUKLXTmi3s+zwlO6N+9kH+hWiUD/yHs
w7jmwEva51ZmtrSNsCeoUuegv7o9/816wRbO1nADYYTd4fzp9Wl6U2OL0g/2LgEpR8Rl432ZpoK9
XrO3MXzNKRikay5pgCvKWLLP7qTGNWvufD3v675NrbRa6YC6KvYs6gC0LnlJxJ6huFShGANLEDAX
MCVsdH6UVi2pq1glpJGhfOVt+SErkOW9EAhhDPN5CCgt0irdRtds1hgnIU7Y+tnl9COsMJY/x2CT
Pku3i/HIv9RyLfLZ8L/PEM9hVLLUwCO0wfNSwCyl90lCv05sBt9nBdOAjvmAM7TnnitN+D4oeb8u
8hznsL/7YZ9KbCkobwPGkIM6b5tpdb+2mfxMFcB1dWUt0NQ2dipo0iulJ111H/9l0YAP9SlxMbd5
iN5hWEcZPVMigYsAob/7OEJJnLglD2LkQwf/g96esReHFL/1c8h0JElhboLSYBQBAUp4P3hnrb/w
AejZCUbq9A5kpeblrkjr28bukWfZbqcicxc9BA5tNQ6uSUIgCj85YLnjulmnH133HNnGFo6e3lX/
rbxY8Htk8PqyHUdst1S3L9SnWpdZHiRNSdYAttTxGkViXeuIVIcRR3DAvxvXYgDSJIRbw3woyRGh
NQJQAbeNb/Qc8v1u6JBxUJEpdBFwVv9gd+0bTUyJKxV4oLibM1QRL9IVhwIYOuxu4x5TKdx1N7em
ottQ/58ul8fUBPzqs9ItdNDbKzCsc7AVewTXTS/UzoF/kwtZCXmPSoccBmVI5wqEQaFHf/E55lWw
o7mBRTVfbAhv1HzuRlB2JSOKI+PwjvHYWTxaP4Q0Gl9qwXPRoblB6e9RMluYU6OUqta7evHq8M5O
2pG4EGCq9Ybyg09XiwYCYGGha0EibT+QEP9Ix8bL0RoSoayW+e+Fv652SozuK3PSAnsf/0e1IHIp
NFpqoH+M3M8GAsy/znN40IpgLMcRj4OcahYGGVL6O2kyQeor58K6bWKXWYbqqfK015byLePczKdb
KcKyOakP3SiBSwI6MRrwd/DuIehwrsFeeQ5TjPlyGm6ZeI4SBBHmXCcyGQXlmLM7CWurAuH+VvbS
CAy/UbfiBf46eMGo79Rxcjb4Bw2v1FocIjLCJCsKZr/Du7p0JiTzSR+fgYAtWB4hm6h8h9+g1uO4
zLDzyBT/yBtSch6n1QpIK/2nA8nMH4MsRBXWAAXmR9cmk8UBGsiYw0w8RdRqc4bJdo39OXHnWFtp
qKBeBWqY1k10AIp8Xr/1YC24SNADKVDPRuOw3GxLjd4hA7xoj1ah8ot2iI2QTcZwibUp2Gp7fvhf
84B2dSM/qxmBIc0J/cNhRTxVVlQUb8ROpCb299v+vGnkXCyAMbLhWgRy7MIvltTn2t7qhFga1Lzl
nyQISbDi9v1SeAruSJGFTJEsHcYYUMaB2cgySsJNlgUfoENsKLzziA2p2UowLrrPjhQ6Kt27uF1C
mo6OIZj7uYg/zWHkPltLmfIahdlMfWUHmSlCYTBUeEGyNIbWh517XEXGOn5wmumQc62GtnDH97U3
vvgtkhfo7CaZQ+GFTBh4/wQpAZ8y38tG7ZY0Gj62XratDPvvz2lR5FIDgTEilV+gHIH13OXphYlW
8OzhaBCI7AFM2hDdZsb2hmDoJSSBLMlHWAgLRiOw66mON6ZVFkLbWkBuI50L3ufnaz6RUNHAO2oT
TL/6l72+7XEHO98k3kgK9tcKj4hnxMTHXVQjMH83FvFTpLg0cVU31RgvNcrEbakbzQnmiQ9Q81JU
x/Cj4leZ9frLUaKKTwLXepp9yvCNsbuitkua1Jq7/HBt+uPSjmHaTeV1aDhCPzIAWMWbDYyVnVQx
Xj0xjKSWeKIyZtUrU47W62lpYGQ23kPkK8fp/ohCeT0sdjfNt1CFtKOAX3mPEO4w/FddQxUhkCD6
6bS453oLXmc0x1udWOYhfUSjyyoZQ3ik85Da2p8Au+Ptq8UqUU6LFm4mY5ZtlMC/lkbSK5rqjgW2
WrfT2MJWnMrcxk3Mp6YCAR+BuIioIOuGc0rt8FyuTkwez2WUdOXBm7ZnMi7zRopf/x8WFXQgf2XZ
pyqUL0yaJQQhejLLR1hiwP/xgirJ33r5RKL25xRCPgGw5lSLFnwxGdLp2dvqDZwD/zOqxuo8qGrJ
B//OHpQHt2o2B/3POd21zxcGQQfBkFMRLb2AyFruELliV4c/njufWgCwdmslV2yAu2ukIgGRgtpg
h3ViMROOLmjsSQpDpcouEibpDfsIkPADC6Xm8HTngPJ3s9m2jK32CB7vwfCJDnjwwDpJslptSEF/
QzVE+wuuU3EFHOwXvtr3SktIVh183pt7XVZsI46DRVZgRff1htz0JPcwjdkzyOorpOHtPRRokfwB
24p1JbwhnMa1nSLXG/OLIG3oM1xx+Z/vqUQOJAOcxH4MW2ZFTqreVpdVbjEmYbxKRuojDOdTBHpR
C9mqgERODBv8AlI5C+9QhfS5fuibCwgzpb+1oeJQeY3a5lcupkaVymzKEfDGpyeot7UEdwUtOVQi
PKAggZJe7OM3DMlVaALfZJridtZ6PrVQcwbicPRtgN0ZxuU6vg6NBDaSf1OWi++qew0kOBveCKoH
RGH6nPZfL/8o7YlqRp5cYmXIOAvrlSnDdHECLFdotKwgaSZjQrN4hYuiXLKhlkL4yVqC1OoxG8uZ
GLE+78jqXEyIiLU4j20pd+Ojnm/8End4wTqqN8Aqky4M7+9rFLwBt8m5Zmg9CeXo/Qg65VTlovTh
eN7/fIzjjkVO2KinQT+L83DLPlRCemPpA74n+amYJGiULpVbIu8a47I8sXaYeZHXOyAu8G214JmA
oPFP88/7zRRIFtRTzLGoGs2VJgb735CwV9VHD0VSlyMAy/YfGz7tLZVrcTtNR0mCPc5tl/fcu4A/
ZJoNQ374CV9hPyhfBUeUPDEFkEmVlotMTtrUwASg4qVE9R+vW9CkP53GvadSoe4vYupy/RyjX4v/
8UhRksrITnpjQaDLu08jNi+3BtVBUJhIRIqCJ+2/yRaA3q67JLvUGFIZPaWpZiDN2LyN48JRHImK
uR9Yw/KOM1I0E23RBaZBaBEAwM4NRTXfT4a5vdXsgbfDR6oBWZr2vU5AQiM5Pu5rK8zWMYC6uRd9
He1hPNee0P/g9ZZNVUMiFFXxefXDNgVh1Ph0sPToIFqNKPVD/a0pQnHtJWOgzdQCOGhLjBkC0R1F
EUtbO4FUUikrW9qTQjgupidIilfCY7ZM5OxpC8dFHy+HU6reKcS2X+lzCegNz4YEYiGRXHLPv90M
JXjv1tPbBx/eSO8HQQVcHL6nAxaaDnyOk4auDCc9bV47YaBAxCKCk5hbLcuZSjtjZG9sx0FAJJua
yY/U15X4zuSIgc677hGaiEMak9eEdLt2pl5/yQTSxyJqWk0e56MUFNOqz4Ptomgla4Kmp4T9Hd6R
dhYSRANK/cWnw2jIdteIZtAEScXOD+DXfybb40kIj3kzF61ERdjxDHEzKPiyvX4Ao0tkTRvgoi+L
DvPLnTdpsNe9WhBFhybCIzUUCeb/JyJquX0c08c0efVnzd8JPJqC1fHWqRbWMlp2yo3f+H0tkc7e
u76BvjwXu8VMmsnRyr8Km5w3hiFuy5tUL5idk2tgOa1Iki7ZF2paPwLAIwBH6bRbqUUhNqbF9U2+
XqAI/i3pLIEFv7Y1ho+bVXVNn4tN2YCYrHLPQgQS+LvXzPRhvJu6Iuz3T8jZVVx4sdjGoLMk7cUD
UFyFASsU0sQz+ZWgLQ50cfDM7re7vlsgBl418ikmqsn/DoKiJIkey42qwC3IP4gay6KF48oBpemv
rdAb3uULTVbI2ErFy7J6X6rcMmKJvBAszK+Wzts5LBPp/YOCJTJyUActddhonbi0WmdG3yu7IvFD
9ZV9+hWyGOb19p3cb/DIyWDgPhMMS8nj+yNDF7wtUHDjnQCCRcHXm1uEPdfUMiwbXkpmiVHmMc5S
CaTXBTIzi1s4APp4IojJcacjyf0Gqzp75R57m7jylrtFsEn1n+k2Zk9VkwKpnfgJmeOy6BMFfjMo
9QgXBClxuDD8CUzGkcHgtrQtcwcnm5KncwbRyFlAJhoFmCO5ioIvOzMesu6hw9Oxsu2hlTeEK0jj
KTG7yqXbbbwPsjPwJlVTz12cs5Xn0NkCPs06REDmdc+1UVhQJ3u0J3aQRHGWD4+zWnu3ms+tXPen
B9G7hok4vQryWURyjS8RJXxqhc6kVpqjm/Rm97qyR/J71coAzMIsA/qcOwLEmFaY1zr2i7B0K/U+
xsnnIVNiNB9RIdLTD0xbYsQg936XJF7JBzlzPD/9MDpT90BKbyjjX0fds5I4AQlT+3atgGP8O5db
vRe+vWP2ivvoOo1PQ4ARt4QOvwJIXfY3teAf8hWI4q89kurQon8UlXBU+Y0RS4W6zka2iHpB7xZ6
a4/Hvoz/DOjqYgWfQa9foCB8vtNRO8so3F0qtSKSdklV33kdHZpovDo+tKS1j98h4YqAtnJO9okc
VxabLW2OYIGsv5LZ3+GcuOAZduEI8e0yTKAbQQpHEf23VQvAVif+PUMwr8uOH6jDrUo4D4gqoCDs
zUMKBUIVdCptkXP0QE4Q9A6aGxKsMJyZpl+3AT7LsctmXAuuHYvFi2dZ+CV1Mf0t9YRaQ0JAOrN2
wJEUpwbE+lEBiAuFeEXYkzENvnadYhUxHE3+M5XWo0hd8zEGXiry2URn5r2tSOCeVWqWhCHDJCbV
biA2U6FF8B3XUfMLtNp5EAJlFrTiOx6gpllEO0Fhuys58uoo1bPr2pJNFYxMAwY8JjN+AmXCkrP7
xZxOofb6wwtp8AM+agD9jE2Sc9Kosf/4XlORegFC5tb/wQy9oZsS20YkLTnSkBIO+x1fQNOnTuir
3HzOOy2sN+SQ5mxDu9EsuMJgadBtMtpK45nai7EO/Mkn9y0gor6OAxdxHjwOAQ4qU74d5rdxLXYo
xfMIOZ4QcrXA9i2hBXONWPi2MmU+pr001K7lXNinEdu0Ps2zHIwcmAdpAKj8K2F5TMBA1bGuQe3n
nVH08tOlQ5qlODB/wt7CGlu6WrsUgF0RVz9d+mATIr5bddwnOGPVxTpBbMdFK5MOwZIqnq0UhV/2
pMm0doeKYeqF4IH4q2XHJsN1dRT2F+9RlsJCn8zXzEPj6ML1vuNjvXMxoM4aOxYFMNu+UwuObXc5
/WWbSY8uzLERSBwS5aTNxQxQWWpcbYIJOMRs7aOxuUxa6CdP2/g+ekDvkv44VC5g2R+YQtwuQidL
UEXAtryTlfQEnqAyY0TmQ0Vq9yZ9kMGFkmSzDdq8js6iCJimN+2XmDzI6ccqTtCtnaEIlnk3w1qO
YJwcLI6XyPf3WgslRrHLjKNVL0otMuYAGEnRB1e9u8yLf6NFi1IiKeoyWK0QtUidofVc72DBx4H8
g57gGfqIqSdTAi/EjLYAcjbhhXBbNaw/FahP8BKZxFv4RCZl0n1ebtivf15hS2pqWCZ53/6/7EgN
B/yzvxD2cN4HXMBbPww8H/zcXW8QLpwPNT0jeMQ1jLnI4QM6STISM5EP/P6W18Brqq1wcgMFQ4W2
fzKEccjEYld9B5Xfw5OznTQvUUMtlgZWsY7xqe980RkRjVXW9wIml+GZP7Sg6jBOXPQZv32bYCOd
9d+BFnblMFQK33Hg+OwriKyrn918uVhDdGu6J7GWHjY7PkSLHyVjh18ZNvSQx60d7Tmqb3TDWMnY
rD3HCofn5ynEXiRjxab9Q30dRvPQOaXrm3Bk8cYIV/oeJoIqWiph2vXCf5HT9ZdaSG/1ghEWywYD
EmJR6Yf4U3RzsqALWYR1uyVHWZFuQ52h+Ddcj5626Yj9qWUdlCQS1cvjW9opcyy3KFW6/UkKqsVY
KQE1UpwpF4PZPfLLSflaFdGT5/2ikCiC2qHkn+FZYGN6S3MDq90YOAJg6MC8siZDTeCnjB+lC6ST
HTKuhM0ziRlp389H3ZpMMV617pUt35FFrI4hkK4euu7Xu4MqPd6r6YAreuCsgqQ2t3Z5KoaszV5w
v70yP/RtZhA/UJI30GvC0RKuKBOFQObodZ2XtXOX12UuF22JhxSsTr88wuD4+3B8bL1COqDA7B44
utEESj+PkPNs4cUiai6xDvEo0LlCYIUrnM3Scwm542cQIjBJ8wMFNQSi+F+FwY0mZ/2IM4anT5Tl
NIKiIUE+PK81BIa34LhMuDvPbTTns6Cdd+seM2S/MQU5aV1JzGZF+GOIfFOs0QRlI3RnSPinTpLr
EXVs6tYMMFTJEDWY1WDKtmpQJYTOOyFp0nsV21aZihR8wnfWph99jeLXNVLPaGcwYHEtdej50YzC
3IkkCFmdEpuW/7JGjabBSK9QNKIqmROXqcv5sLSZgMZ2kBNKlgZvyxzq8we0MWy7a4aZa6oc74rh
E++y0+oFyxWHT4zK+KZuVmFBiE/RcQR6cSTkTrJCeLBjEdT5Ro+SxoaKsRX2n/zPOI2sUnmgJfvh
uO0RLL7CRx2Bo7qzMhoHhid6GMewaafrmgEZuTwCx+X4oZnLgtWFX9Vg3HvROG8/72caFMQgjzX7
tl0p0zwwMjAnjHcSywHSqZUiJbbS3/j0GulSOgiIVEppOE6N37TLynOiyD6da4Ugwcs2CwcdD3kk
7fMiyuLpbTTWzLvCg2kamBrA3da0m/fRKk9gPPD9pgDNOAZs51Nfm0z/7yIF5+Rwx+m++Gbcgsdt
PdL2A2L0NFij+D/dcP7LEru+l94aWOxgTG9sLk/J4DBnGmorBHH5pvpAPzd7PE/sFjfbsRuE30hO
QtYaUm9n6aKTc8v3qk1w6hljWC4weIf8qWYOfTyxvBiW4jpcKEpabxEzdqQWZDhTcvcZ2N7236Ik
0xuIE9vrt0fJ56hzoBTN+Fjr006TUUeraP/H59PkI2JGVsF7UHVweQ5QDP25TVm+VPPuV3My4KH1
JF/owZl+XrrMCQq4duGGQ+nQz6IF1puNDPHrGBPfXuxKDXOK5C0VeSaETDAY9a1pg6JCCDR1idBU
l7L2xiOS4lyUjx9IqOpTYV7k2lY0kcmKWQV1YfPNvImZ2jzxsebOV6jw21t+Zl9PEinPTbaAidMG
WuFyXNR0MaHyI22YgOCWYaaVFB6/6TVEQqAqJkoeIbrwpd76K8bVaDPfnNAlxLVMHw2Zdp/dsaTS
8IpTXuJUHRYzRC9MUa6m8hMAAQ8gOd9nOWFUctTAPl6HvsOzNag7rRhz64pjYoyi25S2BrDBif/x
hhpy4rReAKOoUIuwyOPvPdV0f9xMz6QbQYsAD0X6PdI+0q53St+SqS4IJ3MtLDcIaMKC8GZyKJc8
EpQl/9sPSQ9QioSz7KpcM6l8RL3yVyY2gpZ/Ks8CJvD1j9f91I/m6FkGF7jIbmRciud1RN+6AA5E
JLdTaCbUzyb7GEqokzhrgIYOZRww5liHhzUzse2ZWlQb09rbPNtWC0GzVJiL687sN40fsQQAek3V
t2qPP5pSqEyPCtVy41KaHCMuR/I2hTugBhhVav06MgvzaMDaO/8gkvMjujHSkAzdMbgy+expAcWD
/431rpLySmj17ov1bRtvswVK1FZZABKxLGH75JvAit8Sn531DsjQwdv0HVJCqrZnZwX5QAg4YBPu
H62b6O0lEg8kLPmtkG5ZB0Ca44UrcMkrV2mDCGHBhWWh6b5nKCS6uH0xCZXsckqlu7ziXcoMR0V6
lBwdkDtGkuTCp++TfpCQkYqCnYqS/a0nT5p/RfWUF0/evR+4JJAvSqpqc86Q7k8QTrWDXZlIsvC1
Md5nSI4KtWfc11L+hzLVhHRhoqSogJy9pjbg8axNyMwcWZzJhZ+8wqoiFdr8LO4eDoBasEcyyYAA
C6r8VesiL/iq100oFK4qiSsWPx4MzTeqCiya1HcimTW/cIaalsVcSdNFLjLsWWcDudhzRmoxIMpR
S022sTR2rqch10fBoeBL03vQSVSW01BYJVLduj4bibXykktuZ0rCWP36PcPApaUvW84Exj8p6lHu
0h/TMD1D7r2Q5f9rq6bKD2W/3/n4NhGWZsmTdwP6fr7MWohN2sN6BiKxQvhY7OdzbG20d8N/fKAG
VLnfvXPVbHZxFUHTvNTczNxKerpCd8zAYe4tO401iKeUzLKoYXuHj1G/hvSwCwaBRKT/GVCoNDeY
0oq0aS7auLl8T0Ogwo1oxBmnqOl8BM+KOjhRxr7euHDrortNz8uhVliW3IowaE06gEgmKoYP0ts2
vOxx9IxP3hr7Gy8yYn5JpEffZb3vgBuKHzwt9q+eZtncN6mPZeDi30rLKn4/k9g8a7zPxH4Kdhd/
NluZD59l7LxtT/rVqGe+hAnpBZjJDoMHlNG8kxSybmkGKwwZCCkuP/DMkJ/zDt97tQRRx+RR1bn8
hGjJAGRD9zUrESN4tYjEnKmUV6rPjiXUuDUGAhrcOFbxmJQV7dMTIdfJravqJ+Lcsz78Vl+NcPDn
BKElZvMRMaAM+O+XAqWTX6ddQocGUAW7A7KU8zY93aKtAzcwwVehxTtcquiK7ZNcbr17k50vUa3m
yUxUYnfiOx3l6qX2S40qu68uXfX+ZHzdaUqF4th7ck3dwkDyHP3BweF7jWHuSIUB1M2fKz8F1yco
0D2cUPOkTXKCRiSbQiAV+/Zc/7l1chDo5f+7jMjkv4IQ+C6fdSLBFKdKdta3037H6PxNO90yZF0m
7yLXQSkpcNgixF57pKz60LXTrXOh5ygtFMBQx54Njfj9seRLdDG3mdTvDIzGaSqTQjNtibGg1Nkh
CBHXLAve55SFqN4PzKjW4DPSIcZNoIks4gfM+fw01++EEjGfU3Jc9a7FOJr2C0BNaxfgYiZgn/LJ
CnyK59Wpvb+i+cQUWP46qcLQCRCe4RuwJXY0npBn4Us9qFjkji4f9blVY/NzcUXzvbP/aEdlOWLr
1Fe02jaX9zvcXQQAZgDxP/vokSwu7BqHQ2eLzO+y3Fwm9lMUcriCf9v6rh3GrVdnTvALKPxMWlk2
BJtsfpr/RqjNhn+ek+Fg/qsGYJ6pAjsif6rXQzRELMB4FCfqrtpwjZcQIwWrIp07CDfNvneCf5eA
4rJQSMeQjW8W45SPNYP95CrRnCLmN6e0RgRpVRYYs5UZmVJZDorFf31VmNMIq6rGeg8LjFx1USBG
HYTuBdjiD6zLYpHKr4/0UGs8sU1p9J+bX4Tjio/s4XTkuS6TzNcrfupZ/BU9eweHo78i37zsmBIL
T3eEtn4Sz6u3Xqyof+qKiq6mkn0tG8QTTROwSU62CcPjUTv52GaXvWwPi+c/2dCQpXWfJKDFEpTb
kpYOvYTfThxTfkzR0c7ttD5SmJ7rI5xO4sDHVoMVCnJcbPXT+OVqtWy0Spk4YTBzVgWML+nmdfak
ei8q+VTf/eWsgK4sDus0P7u7rcXtLtX+QneOx/ZiQb7bb9O7fqBiLohOtjohMV7lxoAdhXNf6W7v
Mt+VaxO6mQySCDZOKfl82thEm5DdmoyZYKe9U2WNiwzDIFTJfO7uhIOYl+lLjvZiD0f4JL2XrKn1
rDBGmDeR04KbG78xAHEJv60H6mApYnhPbVBlEnGQaLgTx8mZ+QcrtWrmqYoEgafUJ3LA6rhKlLDF
stDYs3nrTpqFWW1xdBX9zDmx/loYo72xncNql0E9paXoVI4+76pCyCbo6Jk8U3cvXMPDs+0/iChQ
gsyogbqYap/sR18u/BW/zincVwa+mGFainVxbgNhwvevuC5P5zubr4Sl0lsDR8A+S6rHAhYEqL1s
D7AV1rvP0Ys4dsYfu1EB/zwk4Id7vXUuBGm+dYrN+MX4EKf1BYT37ahbnduqvpqrVPZ4FKCEwNQA
THRR0duEoeVUJ03t0BEx6gobtkOcS0GbGrLR1UPvKroOsr3kCrmajkxJJGaj730ohzzt/e2r1JSO
RDeXm/gOGQ4kjVi3fdIZCa7ibmpODxcRTA3yGqf7IOMB12/RO0hA5uBxVUSdYkqwtoTBZIoqJeXr
b/0vXo5o1yoB357aWY0olt2pA/vlQOJCoIu+rkZmGtZkO6RyNMIWH4OU3uNK/b/+T6ChMNsNhSAP
pBZbKe8Ms1Qb0Xhu8GmH+AW7IR5x8fhZF81bi0okAucI0lP6mI1yvpIDPTa3xAezMS6k/I/ABLBQ
kv1MX4n4psZirkTvuW5+AVz4rydxCYoV+R3Jbo8Ttw3wyoBVj6SNeWQ0QuFrNKtGZpybWeC0mmpt
uRQAIpFRz0FOmUNEwaFV/IsvvoAzS58+4He/mn7IG9B58S/wnqfAHSf7zESJWfjv1pZasISmJRNH
8/K7EmoJUK+5yP5BLx3mmGBlxDiY+QCk39+Xoo0WIX63xwmyB15vVlsvzdgJhv9LqxdCPGDaB1tx
eVbEX0Cua7+na1TIgz3FLUd7Sgh/Z/YaumCWUPL9SVKLZRC9ZoeWDFLJQjfxFCd7W+GN7E5zYkSQ
iRhRBn5hIufYhM9LSOEo/p0j2N6GQhhAgwRddNf8EYw8cn2dNTIlkMCAsIu/jbrcsWzhIaEAR9qr
htf2kLmifrKlbDlfmFY7y9ksghSPB2TM9SVXgvnSQuHEy42MWVjz9ZgYtSXooVq/zDwDWfPdIZL7
0TJJBmSOM3T0diWC3pheK/CEENrQVjohaBEh4pK9YyD1Btz720ckd92dftDPsIlkVd8OVgBykbIA
GLldOZu77s666lICPNBBwmEKobtdrrGdAoIzwJCWvD2NBDrG6vdSNIUSwrnePY1oTGDQzMDchqT8
t/8i3Qllco0wWnhv5/GGgw2nNgrpUqRPOevQ1N7nNniPmeOg9xOCLRuyS8yB9BNZpj+TuAoiV9Lm
W/H2LboxaR/EflfYck/9mYzpBI1NrN97+4/gxIUxpkzibS3PVlwu9wuhFNbk9oXLQf+G9huP/G57
m605ncR2BJwWCfSIjIUWoHOocZq97OmWurISaNl/VOLWT+OrYUgIKGzr5bs0eb/SU6WouJ0yh8t1
TToTnKH6O3RLVjJov/J40lVip6d152PVNJD71/afWDM1fVYcMeaId3aCTI3RTXwpzDK6JsAL6eAw
obETEC+PQ0OU87abJ13BVcsQSjQ5EDF6Nwoib9p8mnptPAFRzKuBVsRULvZMl9GCIoG0eDAM4pUT
bqmEfijh6z0sxgSM9QvDcK7TmV2JSLs8HOShQR/yoqnDYe1+Hm+hOXjzexctJL7vCbSTWop+2yUm
D82Md1HyRlDTrdnbubNbjmmICZ7Hh9IsiCZS3FfICLXye3dPvSSloWlhXR1P4mI5pbX2HiNZ/KJ7
EY2QJUSWsx1JpuizToGRGVgJsj0B51I+iSugM9o74oi4ofUC1e4H/geuTF+457hEJz+SzHmZFAhx
wV2OokfTTfSbhaihQNQpLhFCerh9/fZdoDUu9F46fh1zCN1o0wIyIDuIhJZZRh46aglyL63dHNO9
VocJoTB6rvigglrdspF2cSPWYywDeez4lpqmmbCsZlIq1p0mfMlwlKe6sdx0fq8qzdNK17nWWGUF
W9jCooLQeHx6qyYQa6Zgud9hlmx7nVHslf0usBg6IjC7U3K2RM6NAhh11O99k2Rf0VCt6SYmJPTX
BgE4lmpC8OML0NliFhLvF1rzUz6utIE5mE+2Wbrrs0julnF3IyhcIHRGSs7/OzgNgSFRrclEjts6
wr476wKlOjgm1AK5WV4fbOWMqJSk2MA/Y1BiYR+VqBoPzxsR7VAMxwfFP6dgKs5jiii289u7EO3M
KEmaZnLmvif1gtz20Cyq05qCVSvlbxsBtxvm2yfjfGNnEtn2NRtMYEfPLhMj6I5v9GPQMZ8lqld9
cf90YUlkM/PXtEXXglsTUEBMdjHfiDA3sz/XZNP90bt96V6EncKBmejoTm6VT1bqfnZ8VR1uVWtb
iTRaw4xsHvWx1L4v42HfJ8N7ExP0qNU00z19jf7nSuwkGfVHsgRdzmZN7ILwX4jcEniECZFhr/qi
5aj6bxpZrU3/tTLW94m32+J4M1X0P2KLdTyLpgKrti4hWMupoqo9LTTJRG7N81svKdJrdTwAjY3G
UNuwcjVBgFdBhluTXSyxeq1yE0LVU1IQDMfLjlYzQ5vnFIgJtfyPAo7QbUFa5uFxaBWdLxrRTKLo
JgCXmK/wVPH6nLdxh0vN6Lbkb+IKgVQR/MLAIICfTZ3Eiy6d6PT15k8EPYsc7VopEf6Oe8zqZvlf
Dywasi4J+UPTG9OS4VBufCMow5wh6jnIre8m+80CnPt40rL3SNaTe2Z4lCnJhmWgO1C6YB+g+nx9
Wh3fiYdULikY4vkir7TWwKWaDTdStPvo/mIMUVzWUiKZaERg9OjoPd/3dtFgaBJGY9ax6mT6G9Ud
jdZ1cmr8jULhWJlBWvdGgW75m8ne1nUJC4V1qvpnuqU82G4YkPl1+VKZvChmwSJ16vSoeYgq2hk3
TybkwBAqWqZj4aPLsdd1PN0DyaU9U3DupuX+P1YYyLW6hCq/44E0/Rkek04RVxR6qB3x0f32A5sO
YqozaSV2v4JEwor5z78bIKOKEU6MuoYJDYAbCKbpwwIoTYtDZFMJMu1rsnwzjVAv5Fk+cydkKRXg
vHmWujF6V08q+/8l6zVjBdYevb4891LTokPqFBr2hDh5ObkoKTf5ivIjwjk0/cDHVfnJjv9JdDX0
iK5CZuWAvulPsIiFZaPZFx0MZeEkZz/1GtFcTccIwDHgF2/U1SC0ULEYKOc3IqkuN9bgKGCjvf1X
wlpPr8JjRnY+pCE9U5wgtc/hUXL7agNLBzjainROgxK6XL4n8SR12OVOnKS6AEWRB2/vScPqmAuf
weZRuf5NV6h8xAcCMsEpy3s7EbjOXDZMk/0sOkfIq5noZdXQrjU4DxqX3fvU/N/momoCmceCKA4J
DOTb0Ql5pknbFv9KUJFcYbpmB3xNc+M6PjlQI8wpJfX2d3LVTQTjz0Ssf+oBH+VFi+GkjcZkaiSM
Fz5K8A+jp1ylpGFFuyWG4JMhPTkZX2FWe2RQbrOqmZhmhNcYrNm7VVz3ZzRR+BdYYsgoFjWg6Gwm
LxjXG8aHV7GKYFzTN7i1lqrb6jEvnvaN/V7OhofT0/PSRunxBFZfZ2W2T8iV24ULGOeaxow0Nmpd
j9akvoEzMwGhLyw8OA3yyJutn4kvDZwC0pH0Xmpcbm1wh798wwJTYQwQbqbERSJ378MiqhAXbowv
skNIzaHHEdo/y3rx4SvyedRuYs0sFttwCr4dnAy+3YUnLCtgPBxGrdGRVwvRAnxQGCI1EXptdCHK
ACYB1Qcb1LYSNYvsdOhkisagXXLGOZFZpswGILUcTjaF2st14MMu8i664TUET9rbrpdkcZxQ3MKC
33deN9kq5gD1XohCZEdOGry+y1LuYl4Env2Z/V702xTjBj8GTkZDt8gTXsuIfUnQO4FJn6tENK9w
3bZN4s8ALlh/xPmlTvc9AptugHEzFWH33YuW2UOOaenEiiWl2cY/y/vZTp+IA9oSKJ65Rx7bXBVh
p+VmyE7EhpP28aGtt8YBQQ5B0vfdbAsRbPEUvVPucjwYdEm6cOSSXAb0L8mTUjAVbEh69klMFUYA
jx0jxi+DwgBMiffI8c+adsepg2xQ1Ah95rQmmGGP8gU/ppxw4hGRkG8Ck8G2OjsHdLCD1bhQU8cD
wwyRnjSS20UojMSz8fwvFhSl9jsU2XadSmVIJMAaoTcDgMuKdavz3p5NHqLTn+nhV4ueRytqmPxq
wE5IvCaWl6ExFe7GmILV7l5C5lvPVJc+UwTrPCL19oO/DQlCcJTsStntwbX+lDjmmTnweJ+8790e
QuVq334GVMyNk7ksVbooZ88ZZwwP9eKp48fOCCqspEOJO0qmbGWrA78/QaR55fRqlKCUso4YP+AK
7TQJLV8LJB2B8RO2/w6ZAM3GZpvQLiBC42WQRe22hSSg1vtYF+CsJHiPjhYkupyeHR68uHV+0gyq
KUO8NiazWSlobNV00MaDcbolnpjtFtdtvQvk3nMShnzWzoTyP1BuH14IdoJZalrWnD+8uHxkL31P
NlsEwmePVag+3JlWeZKp7eMcASSFKsCmf/fjMK8b1ClLsqV0Ik0daN9ItemDryfAo8sg4soIcTh6
7vbS9a1nHOzCAZ4f3XUn6UO4eChbIMi0a36PNtQqoB73BckzvXxcfU3xwnKypd6TtIFUw1knJ8LK
n3EfuSeluRYWhQFltfN4eEg6NXibONnEU02NvTZMeqAE7DKFgeyWHGrBguwLhNrnORQ7HiAs6VHt
7nfupukB/okbeyp8yVDrppvk3emKpcgHDOTPo+nto0F4tuBGvdTAGsZqOHQiahEKSGXnj5ul27+Q
z18DI4nmMLClURgm5uyrAjsZy/exhz2owaMcU3hrW8VOfVxHlla9YfewXSuoqc92OWE1HR7LZFwG
X4fdNo6NlRn4kMw9rvfMLKZTu4/59W1SOtlXowNXp3n9VdT5T++YHBRpfNMAIxLFibeBMdcsYUD7
bqPjLPnAy8MLPi1lV6r9BtdXKtJbuNk1wNvCBza5/A9oGtetVcNq2/6l9Xg5hcegZhXnJ+Ao7qn4
oOp555Uzk2NdAE5wxESg40hlEzQIBVjEtuumJ0wxE2Y5EX6UUuqZrhsJpMWZ24oiBtXU0RkC/w4P
P4EdYXogXA5MYr25cVJsUPHkyGuZlYDY2oiQMM3XhPYtDqJinSQYGg9ivSzCmFwk6gWxkaHE24an
ScLW1+xabzZQqaln8PWlba3H52dlQ/8RFxYmYQjwfzCuxh9aL29jn3Y1a3uCz2ftC4GK1E2cWBia
m+ybd5P70WT9+B0HFLTJOLUh/8qmudvXfLgmI2A3QFnd4UZ8Wmk+Tpkvmh92wwnhWwPw9L/yu0PZ
OkccJF1U5kzdR9QJGoE5RibVyC0XZSjgGBkAEffyyzhDMeNs2Y6rYSiOs79tpigm4sRcXocH96tn
4LZq+Kg3IkPK5hRZ6AC4dre19Q4YW9++vcgB9okpCyVXyPhjz+/2qNM23tO+c/CWZrrz9KUl3Z/L
QSl5YZTkf8tGjGnKpirwalQFKt8lUq1gbQcmijREFdRU9N1k1ca8XtzFrB5+DCy9VReduaY810aJ
C/gqZCwWS+ZX0nzzrP+HvnvIlwylbzBvmaSc1czv1nE6hqI/g61gBbBD4kePLKoNAMRtjfsQQsRi
ngmwuwbpg1yuFmVHcbCZwz+CR2AE4dISN8hM2I/CZ4KC9Gyj7gAqy8jHnbIrSnlm+NyFM2DJWVl1
wicYUHDezlYGGzJJC5B8MAmf15actRwBx040kQA96VjXs35eQ0kk7Z3bRZziR41DcPaLX+vsbcOe
Gx1Bki866Qh/+JTYDHp7myBSjM3e191F6p1/U+wp6RLO2QXOQyKaQfiR+d1d/7zM5h0lh1gw63Ge
1B3SeYfccXqB8F06rQonbceTqr9DeiRwZaw9B75SAG+ck1Y1C9w3cMPu2TVcJWfKu9OWYyIsEU1a
7aM2oGsjzFpLeMidlfYlgdWcYUFrv8Vs4w0In1f46qJq83NNIrh4vIeIyw97OCn1nkYjtbVTlZbQ
WRKkjKpum3NJYsG03zEmTAObLWPfS3MBjWMUtKzsx6s9HlJ5JZ14vQI1LDqTb2ba8Tsw2QeNjCUf
g+GFNd/103S0gL2GyssV1ZVtwHRcu49giUsBrokgE08rnkvtGbkToAnceUSXp1XvP718WsxigtRO
vOb+AGG30lhRcY7l3tWM5o+vEVLAJTpGBrcnCShOMYjC8YLASQ+fk7ZwB7ESzzs1uYqSmWPSWLol
aQACYMhNyHaR0tNcC9iJqYErnRxjejujOD0oebeQbsaEXq70BX4etn8YsYWOkGRdKC2d4C5CkbRu
hikXUMZfT2YJ89g8hR7VmXrz0sigEqXg1t9mpAtoijWpDG+E0i3BEea2QmbUuiJxDvSfh1HCR/e0
rO7mOkoIi+eQQTGS3dCwAuLiSv1Laor0WK7oF0Cz/AMDnCHDLyHiNEw63414p0oTElcbuTuVkPdb
U3FGUGhaR/KlyZFoEwUdv5xrbCURweOhMEN/GEknptv0Ihght313orz+A2/elZ+UVP5DTPgtgJ5y
wV/gvsaw1fyv38s0a63puiM6HT/42rcuUUxTJUtukxBgdQ0ZtQM0LNRfFk5Z5FQxtv2lBTPWytGk
7LmUmIS/ZKY6vrq0tR+tlvAh4Z6F8zVgn8nGR10NKPtTIE/03LWTr+sVZ8lqHUiCYnEeL7eyEwIu
dYLfKXMDy/h+E52ZF0bfPG59dryvfODUbuE3x2nynzvbxiuD9YQcRB1rQCA4/Zc9yuBSF71PWW6G
rIa7HO6l+mWti5etLCPCoLKp+jf7iSviakAWkfu2aDKmVLY0jfy2PTjUHVtNDUEBWUCmfEd/wHy7
FOApAa9lvaLgQbazqN3VcaN3V6hVID5RDE9C1f2NFjz2PdlbXMNiG/XnDLPDEcNzszufIKmQncwU
4SCC88uJnVJ5IeWKSwpfR++ziZb2JQl8fkSBWjhLJx11QyCyuEsgax7KWcK7vYMXyBCEynXT5FyD
GmL/4dWtbUyGXQA8Vwk9xBdkOOaQsCqCra8itQJ+757IokRHG5rBUI5h8/66u0ykSEvoT9UcPKSk
Suj7NT7Gh+E+6uCxmWBi7tuKg71rus09mOJQg+ezLJosLRkC6sN0cvbTcnIVOV+GguGE2aWKjBNW
9yffMufUMkurj9OoXoBo9lBwZiq992CAuQe4BKWUWru01jItSmB7OIHbkhxoL17OMxm/oUgM2s4V
8ug8gCsNn+IBonMApiijKU5tUcBBrdsjPvRV0+HX3td28fVPj7KjOcD+05821GFFvYBKPRyAZ/Q1
4A2CnzS0PuWGo094ysFnCgXg03ip69vYxkvoRzSdQnPYqtJ52PJnEJlhPoCHuMLc7YXXMoTJNTVF
0y39iU0yIvjyegQ0gUjXVn5ord89WkbIpFD8wb7FmZJ6719OOLYqkaj2cLPOfekaPfX7ni2Hb2h5
xdxACHjqYomNzEBbfA2NMTiHMmpDpkp8mP3msHDeqVrj2LeqQ085wJc4GxHAb+V74EIVCZ5nzC8G
wWs5TcbE2tA0jvgI5bKJRxTr+Pzc6uSAGVvOZGBLuE1KVlOd1Xo0HFfbxV00xCRaV83eLjsV0r2O
05/X1/+CcOJLmnXAPXyJOQNFE0l/4FeJ0+JNVxEkisN8p7fiHHFcOGfW+/yIjBcgpDrh0hxJvwME
P4PbHRy0ZV1UJANToRvOvulNifY8wS/PD0bM4Ot0RJmHBJh9jmwh6IA1sX672X6V44K6Le3pFjxK
KNkpTHUwnB4/UqhwMCMnX2Rts8uVPHuq5LKuW4ePOGHqQrXEvU8V5aG5u52ck8Ux6mYIcXgEA1ZG
9+uA5W9YeESInamdZKot94DEqJ6SZl8pgMLPhd24fm0jdzO/q8iwXE7bcDEDr5yvus+N3gNWWFe1
JP27J/SDS1y2YpjV4KcI85IXqwbgeUM2kEwpLuH6zllOtsr0DSNaL5nOXSVpIfU4ONlxq4Jf/50x
8pamcx4NmqLB27464uAyCPXXtllzimm8fn7DaE3wrbwWraRi/Lc72CkJcuSHgTenMzhfIV7EzeYF
paD7EA3X6OGvbTrdg0qcQRgsb8gXD5nsjJjjr3WmK2DRnSG4tl85ta0JSKjWyLT2dDJ4+ZGRiPGx
L8zJH3RNxiOZmrcjgSj/4Efr2iItmbehYU/fuipyoLjv3lOeZyWBwI1hNsWMqskCoQc4nSM+kkC5
74WV1Fzy7FGI2sSWL7w/oUkxcfD9oZ2DN1e7tp1tQCVIKeoQA6hQ0LITTd/AWoj19MfG5fNj/Bkp
gatFEAT/MDFCzuonujbAROHL+9D/pFzbYOz7/GIeXEKjYenmmwfIcbZyXyMgjz9XfhWC/Gp+uhSC
GzZT/4nA7QqhG+HX34AxE3tDD0pb2U1NZdgCr4Qp2i1LoHL6yy9H1gYgRink81GzGqZi9X3MLyxI
XGX6P7fqFVNokjtiYLYUxz2lwAMmKhoc0QAaCm9H+PKktavn8xozASQHfTrFBwK0KzVyReIvzS1O
T1rJ2OLnhC64jOMGV2HGMJIWxeqZ+RRTjUEVafxZJs8KcJFCi1MINhLRwYtv3IwtrtHCuOE2ny3v
pw/5tfDGzDyd3UF9WabiFHlPQOcBLfGKwtloydF0pIL717h5H4waAzWRSZX/aJTXXcOxH8WXPcx/
K/ZTUsVdv2OiEnDgI5aFNlBSDuItFUZSwuCLTplVT4rpTUS09YBFxpTMrqMMDXm3i39HiQRshApr
zK6ZP7TjUExuxZnihPAqvQ93lMP9+4IpaGxNJeI0IaKj3iJMkItnQMV1TQZN5M5+wWPzx4weJUMd
GIQHUqyg47X3CKLwsL3usXly8W+VQnG+1UPUYaAHuTHaXDCzTOBXvgVvOHDgVFWN9uyxZvSrdTUZ
RM+I/fw+5D1n0tiW3K3GKkWiCu/NEif+GcR2Rrb7w4B49rFgSeFU7C2BmtgAJf4fiVKLf3AiIaxy
SOrBg1ts6vFT+6239Hyyjq7wdlrUuPqVXM0hG7PksdTZ3XnHquQ/qiMl3QXU1uKIGMrzxC+54YmG
uWOnQ9aDryO0iuuRak7gNVUwqOpBTd68i20beF+MoJVUBqCHKtXrDt02GhqgOEPuEl3tnlhe/qoV
iUJp89VR7TbLF4US3ZQLpun7F/oi7Xk8wnTkrMSP/VyYwf8Tta3B5OGhH5qYjptm767AyzSYh6b4
xcZeWzs2B/W/Z+acPjQkO/oPZJoinKaNT1mLwAS2fbc1H2+hpKYr5O5gXSALnLRlJaNDsOJpdxlo
k3VQxJOf8CIGf/uzj0qYiF7RQ8wteGW3BWOQd5K/azgyQ/bdBLv832YrDyYxfH4JkVWevzhT3TS3
MJAX59FxTRyAgu2U80phx0BREyEg8Iw7fewpf2VX4KbzP7Iuk1+4Nuo4K/eVvoRT8zkBfwkmwGpm
fJwDYOlg9UGtkKKAJYzLwz0aEbrOrsWB7+wc7JeY8srA2P66WfBebcgmIGX9zoA7nKuyJnQfSIMj
J4eK5uYPftJezRlTTM0reUYXys29kiyJ9Sk4W9Zl5IOHKqNG32IztGWfVumP3Yr2t3rsmmBqiHCn
LuHVTBm3COSYhIHMy3tBwpuEkd78F/zN2JDwh0tlypUvPgxHQxoUT6iZcP1yZhNbmUfj8ObkuXR3
MjMEY/qAIrwT1pH+Pjf/GJA983CGKshFdYKEaR9buTqoJe1cpAdwQmmxXm9h7ITMg2avOqZwsh/H
I4nL4MSzdnaU9ZXzJiOBq0knC9a0QWD4pSs4zWuLh9/mWD8WYmxFlQRBiinzb1ke9Vel0nZL52Vx
d1FQmL/8W6tSU4cXmKezWwodL8J027XJp0zst/9gduO+mNxoHeDxOE/7ASPQ0Mf6PXOJ1v4PovoA
lzzTqtgAft9PvMsmBoo5Jl/lJu4f42gXLUSrtWsAWqS0Ba2rk8KCwfld6FZgorxHwsHvYqvCSIq4
GEa4bwRN1a1nSYMQaWhecM7Bj3XLgUeSZyiYXIrgeCjYRFUUu7pmLW7xujZwN33qWI3JV0lH3a96
vxNTs0/gWeqYicGrFxmVs0MVhpRR566NQpbWX6cC1n+BVwPSgbdpLyRF+jsfl4svxgFZB1gVGt20
1t85UDMjXq0rr+m5VOYcj/kMiUPvfkaxGkJWzuchZLP83cHiXlP7Pn/ZoUW4eIn1RIyDvvYAt9JQ
8ff/9TmvGbS4GhWSc7jNM1CaSOWePaBknee4nOFQQpcDqcWaRRPnjS2XWvBQ15qK1uTlTkByL/pB
k9JgNPvEOyPDCKFsPP7l/zhQsEXbMqrbDDYa91D8ruUckeyb1PUllNWFvxEMQFvcUuWNFRjrJAwx
bP5Z6bF+UR4+Zy+BONAQ3H0kSETnukpgCzCt7DAtuQYOLHHX79l60uygbvMdR/NcFxd082v9rx07
eYR1jCTL7F8+oUP9+Jq1+G8vQVXdpCZ68+EojWPUAxL1n77MpaReucLZ3cS36eGDz0hgQ7I/fGmR
YfWTLZj4XBNmREFjL42YMTc+/1n9F3jQxn0wllfCK82BTBPvnbIvhCuiMSrUoZ2Py22w9pyUPKUF
vzoqKV4CKTAqJr5hfLPHBWZ9DWmUG3zhwPG/aP6CDdGsXjr+7sfn0PEqtEUmECnCrAeITe6EH5z2
01LGxjE29FPbe4iJyMQymaahZnOEEblL+O6fqPz7duzlbYuYANjgnK5HYGlTR0WZLQ7QtTMPYZg+
/opD910P3ZuXn/S5Hqp1HNrwFD2eBxfrV/vScTeNhEqh2zmkiDIa+X5BGUqP3bfPScshGU5zk715
jsB3bdCIx8jacC73PdYGbmaR+IQrkA8JO5UKqwPaKMoqCWyWbAIB+58EhcZB3Llusggp0V+ZnjsI
O2M5S52HiiRSgYIMLeG4/iv7LmXuWFizycGhnV5aE2jTIly0ROgl4jAZ0RdjKBu+Ar3VHHk9vDcy
4IG/fnllulc6HoHKK3U0ohfecUQlWm25kNHDu+CUJ0LvDcqg3FWPP2ZHaV7ZoO/xxEEHF7NAux9W
e1i3AYbFDyjH7zFw1xPGy+HqCdjbSzucsr84HJEBBi6mQI8vBq04hPYNnQowmOfYhfBt5eppUbaC
WrK24wqRJUliUc24v/k3/BGSwxsyoe3NIObVlB6FS+mtZnPXoXiR5JLSQatP4KffPyL8K5Ok5247
kgPi6KpUClBcrh2gB1EJmeNlboCOTbt/KfzTqAYAh54tD8MS8hLWEGBOqaGA2ecANw3NyXGdGqYS
vOkV4XNhSurDkAG/Oi1VhwGvWCVMq8ROGw279vm5DDjp617AqS1dFDi8Yh3N++fC1lC9N+lrF7jw
UkcXuqnIj0OD4yfbszoSbUu44H+eyIDE4GW6eMAscrntesLpzz10dRKBEz6j1Z6gqwuACEeDJT2X
WWbZhfw8HtTm0J9V4l0jGq54SOgDYiJ/PMyEMEWAQStUbgspvovHx5yskR14wbmPTnvsZ0eIIZfF
xM2mV/GJMXC7bUhnf7y8i+yIekodaQYgg2YulrGKBofE+HAWOq6Ho1bP7DpK3PRvfHBGqh5WCiBS
YdXYpKue0zcIWtzY8ssSp2ipx9nD7wyHLnpfDEXvclIATsv1If3GAbnXLDRIOwURSExY5GAZbmI9
XHpb/TxFPhNhawa3CcsYrOfCf7KnwSzzCTD2GjPQS4Z13xZrutMYq/1JXHVN7SJbs3tRCwZ6IKHO
dwsBqiZaNSsMs3sop2S5W9Xuw/4yl/NrzufBQasL60VSwGGBhNdUJrUVlohxbHCvl+cLIUpLjXoT
b6DyGyZI3iEBYMSKRkDfpcdDmH6YgeulEk5AutLzyZaHbPQ3Y+38TpfLHAo1TdQ2GEgX4ev1Af9v
PFHe8QkdAPDwL+YzyzQhmgjdA8o/Ao7//sP1NCiNv1HQ4wFbzldvVt4NkuBRbIAdpFeGTj5FQgvh
Am3/jKEX5mLfBlMf/KT/rP6h0HGNlw+outo5nr/HxhGGuKrkzfN5l/a0+qQN+0unQocTu3kkQZPu
v80lZMVAlH2Nue82qv9qTGs0dmsGbFb9FYJnoOeLGFEHi1fu2V9musd2r3osseAmURYNQZnWOm08
PXObe1qPPkxuZhDEGrPpemvTF9O5zANVQMYELDsyP7NdyNtLZrN4sfz/A3GeleTL10vPZJa1QWMn
aD4PXHG0xiuycs1pOo4C+Y3yT1cS/mZGKmGav89ODuXn+UwYTjC+JTbN3YC1GGHb1N8CsEhzeUMY
pP07TlFuRPBE/y5pLdirpRSd8I9X0SBDYZmxroSoq9rxr8kK1JXakY4PmPxnSWkzH3ETYJQmTo17
C2uaza93puHKt3dA19MSvVYCYas60Mr18hwAXqZxBr/eyR/tRhB/FLkdmNZQYzn7veZsqVHQo85f
RvB+GacgJQqoRLjO19crtLEU0LVPamO/yxbgbCcEXchue1p4EMOKntDv3qPGtwJqgowF6tpuAXaS
2vdue3WH84U00U2IfazGuYIT+NFhMk8cZqZbn1Ktgh0xTc6GmkLg92HIVVw0odCGtmfYRyOtbMj9
O3YQSHuXxbxs5JpdY7l2dfiFVVu4qiCEPE+RG/LgHQoWtBcw4NVSUDH5WpjrhrRCAEDFJ3YuXgjg
zLLIun8/Xh0pujkTIKOVp4wZgQnom0ucko4PGIBNXVAIMkhCkFRdv49QxjXRqOQqTGhFsImpKvV4
JWNtlwlvF34Eh+fXnPYEgVs57LibMIpwuGSSpTr51DuZDAY8H2aJlqGCwwKWRJaBCWIT/ythkJ6O
Gr9N8StEB9jl/y7z3V77HRajA8zTWkmjxnXD/sNj+nzSyVlStOn669WhzKyspYlAF4S+GWRHjv71
l/DESKmimYBn21YTF/8BY/LzXnu431H2FBDbTA8r+mPVGZGV8RB3SAJOpmlFszCr/MJe7tqfezRy
+VYGN4o8082LywQyFezZHtk7pzyS4CJrUrTDKU+hCw2JwC7zh25V45watq1XuqAcu3zxpqZWyoYN
hbvjAF5Bxdo0M617yEiikL3ukjrDdFk6i+jiYsxW8eS6Q/EP1aubTbs0FQvP3bwhBRUbmSTriLmP
cUvygXRPdhh/QaVHiuvSAazxzyy6tBR5kwhoOS7Pf7AaxhYNXIHaKssReCzyypb6H1Yh5Lts2uB5
hUOq5Hkd0rzE72EVs5lROWChvMaiiqTMYCBMQZYaKqRQeArSpbDhzBhMHA8htn/0ynBY7pIgEYL+
qihSl2BX8woX2BzscX8fGoKwGcFtUsH+HdNsAc6ca1PDF+cOQ7lik3RlpEiNjJsfFOnyIfVy3wXQ
EWma4OxxKSVNxpdPpjHX2ykQB3YOuYssgiDp7oax5w5xXpGlQcppMNBcc6yRSaKlfxNurD3bcv5Z
bhnBCHoGKqMd59kgVJVl+sswq2aYy69iV6xkP4ZwAKOb0Z75bfG+C3BnCyVMQY5+WNWxJydOqvb8
hSAQRKA9faa0u+PlWMkrG2NrwT4ALaqRHovJYZGzAqo6ksXuG1AymaiLXIGkTAo75N5a7HHxCwCF
KLi3RQzdBlgyu7wXfdfCnpwU05ry22gHR4v/jR4RkFEE6u6cls4nFUqw7z1xuLEMaaoywYnxpqDc
zKD7Sno/L1kOnCJnL2a4JPtFacsS8SkeG9BcZRYAYhB1Bnwb93ssiXxd85WStsrhx4YHD/+bSQHq
g/FPAK09cgidAwfd10vpSWI9lGpXZ0Dn2cTjpfRVa2TFWZcmrnOUXHBoScD6MsMbMZuKVNR3mc7o
H9yiyXx5pr3GLvQ/I5PXI0RW9Vgz+Ql4bEefqTYHj+AOz35zBaatEVjKdiQ/3o7QfoXU0M7wGesz
axyVyeRUwF2gI0bfd49V8iW8/TcrDMv8n9BtDi4aojeJAR4h5gWO081ZopmrBKVU7lNDYWbJfIHM
2vTxXzFwsdRKkkQOsUIKalNLiOQ/yKIfqk/W1FZDJoDkL873fn6oS9wuXd6xGlCPQPCp7vEKuQFS
BoVzYJD6GEApZa1E4VJWw+rvdx4DUbHWXcNmU+djgxrhzqmVybsnnEQMFRQgyOWr65xe3BVa3w31
wEnvTCbj2+9bPjKXn1ALyWSkjY7FWO2WgwybO7sIe1bJsnK8azQE17rp4IQ5bNzvM9xV51JdDjek
8nS9X8QXf30d1xrLEDSIrwQoHMXyBqgKyFbKuKBaFNX4J6dFGrNGviOlYeG4JKZjaLGSjy/TUhHm
wfCODts6kUe0fCVlb+iPsApe6CGtKm8uhr0yG0jBTeU9AK3wtf77us98AWS97R0myi5FE095POIw
4+d+3M5XeRrIh5UrNOnyImYU4Uz+ll2B/txNbKpXZ0MygJz/hGqT18Q7Jxa83STEIRtW4Yef1L4L
cPh0EstgoN4HqIIS4b6Cy+00OiTkjc60WX9mOuANwxrQrnR+CABNqHkaEjREntYi8TBj2N7WIoxj
zyq2Gn1WOwOhZpNacUVsLzm/jiWCMGgzZK/RN7BMsErBKWx2Hd5R0t2/9IyNb+hsoBLRssWgLwz1
PGVm8cv/trWXPIfIqgz6m8qn5cbRlJFqjrqfkSug7evJvn1fg/V+3vn/JA3aiqFh7Xhp1nysI1fg
JrKsbnhBdIZraJHkrK/mqIof5YRFnRxICZsbUlA9auwGR69vUTP/is+vFjkSuyObcxt5ELAizDvZ
2SJoncVuGCVvTJ0r6fgAZy4AD3m/9mw14IPokzEGK0m93larIWQXbcVbTa1AePnDLgxa63S3sKba
fW/1AT9SuaE6vQBoSn0HX3IAl9/GxLuR7cj8WMwReUNBa121jhlz7pWemsJx/UQtyvwLPgIxc+Bg
+Tlmf6DusoEw/DNvogT8r8vjY7cGg02l3njQiI6yuJWIcwB3tfG23PuB4XCngIKuzFezwn7l4kfV
ZBucpOAptpc4Ll80QCrQ7UHs2zOl82SYPwLT/MILNP7oyeRWp/+uw8ekmSwhuyWqugfBbKh75ZgQ
v9WwFNJl5z9Gw2J8XWFKXxQ6061MlTtKZXID8GZtvko+ytiK0Vo5qU3BqhQ5fSF9Goi2adYGn66r
I5LBrD3tLYN4lcP7bUYzmf7B4PiUlQFgMUMBEqDJmDfZD09u0kRJIURgO0PTNp0hjhaaBYKwkVum
ZYKk+ULs2LwJVwPzQM1NFkSK5lGGvmLKwH+vtqHHAq4x0JNwr8/aqYyMoEh3SdPaRfABmjXRHs7z
+pSPSndDPdbhodzJXrLE2JReNCapTUy9n8sjtJdQH653w5llMacyx6c3cu5Rx2wQsAWtWCU66YeH
cdf4h3uDQ7jbqC4hcKSulGuvmFYJeUGr7rQWm8LN9TDrgoPtLesywn3HrhfAEgeWxDAPkob9DDuW
KRQ5cblz7ncltw8cWvJvXfMax3813LwtNB5ms7frhvbvJ/WqhSltYJk60CfKzhJcqzTBxiZZuVP8
QluxhmvS6T2pESblfdHznHDlw+7bbDCll/VbhqmcOHOLiDN4dq6HJ0zmtOQIfzvjpNpjv3cikk6V
K25Wkj9PpFKKkHy8ZRhaEsF6FdrNsR6cm6pntrS4LVXF/r7QkwSrB6ZTctpk75v64YNLwXTXpNbj
nOme+mWBXb57Ik3k+y9M17zzAHLpXSMwfjOmlywK8J6hw15vWuRYbj3dpVcGaoRsPz+QcYPGpam6
DfIKgfzM39lCHE0St9OAJGa+nipF1fdSP/n09sE7kA7XRwfgkqX7TVNKTwr8Kl12f7Que4JxYxdq
LipKzmGOEXcToEFBK8svLr1MFEIz8x73KrPYMQeCS0/w1VmozgMF1D979UYD+M6BC9ITd39B4hTY
KfZZMbcC4LA4eKRuqpouwhr3A7CyuVndukbCq7q/ZYLV7gszVbCLwwK8MQRBFeQ+2QV5XUYGc9Q6
kUg4wAwtrOi/PyS4TfWd9qh49KccxkBG+0OolUbaQoadW5TZtOgJhuK0XygtSevqGWMeyw7H1tIX
osQK0OpdFKw+Xah0OSdxUZgtfHXh1s1k58mUVDRr7elXKL/UHpG1tvCWmisLdC3NOJjAUu7Dqz7q
9UmhG0IC2B9NWUQysxpSCo6t1Np3FPrp8+PhjeN6JLJB0wOlvTCs0YN7qBiSNCW42EQExpzUDf2i
qyUL7P3QnyAl7YJ4WwlI5c31lU9t4//2j+ktwUSaelBRYHKiYRBFofVsR/iFsBM5fNlUUNc4XsXS
UM/xL+snHKrBSdffXQWcck2FN4vpIT5fRKZ0VrEsuQo7laiBC6Uoa9n1G+LNPmX6uWPHzFGqkFQY
jUlYkPdXR/a3mgaP6/fZyYSZePQyTDi9M+DOGADe3a19TqKrXJ+cgqJXsZujFcVqBMQHZUXvM18h
zfpoRbxY99LLdV9K8PJ2VnpuY/N5pHB8r99k1lWk2506bJdytW/usZLJKsufj0NyXwyTxG1tUTYz
AbPJQ/p6vUxVHpaJbvX0fVsEs0sIc7Hxtv533QeXjRAZ0wFOl4h7avJoGqoirKylyUwwRflGaUol
JFYKqEscCKlHrV+Rw+tQat2WPqKP+CwjVeaIOyI4r6xmtIoW/V9DkPpsNQSXddRIIzE/saLKQA3a
f6Bk/oDuP9iBNplOHNwAXnJXLFbR1cyHrhFjNYMJ9BZHF83tMxJYASSHTqi5qmmNjzKHYxJyOyDq
k71juGvhX4NHOKsVchiJRTFj8GTGaQmX5+Mu2L82D812u9fZ4KeygLAtoK9+f2hHsdqE7ln5UfO8
KG/mTDYbtElYHywxmg3kUS5eogE4XHDFJdZZmkqJPO4/pXwfnkGUKyYSHYh4Nsjt8l75CcJn0lNe
cekAWX3kf916/XwTlYFuAZ8eH3S11yARlgPcig8OGLHXIb+jBQtDDEIvUJaWeDJuFi/vwahcLXkY
hpHcQiEuuneZIVB7gCFRTjnSorDehDTSECWsA3Ua/IO5E6w4J/i/csMBRAU2CKcGYp/yllNP6Ol3
fhyNe17Hq8H30b9g3I27kkYm7th6IembExHpua2pwsHUUSOuUr/TxnmVYnAByQioFUF5vgyhaNbE
ZlOSGg/yTl5PAOBC1DoVGs/npCdNVraB1cJmV3Abeo4KqeKaMcvp+vEDsA43K0HVIQvs75qbgEzU
MC8X41WK5Pc8vb3ejnrVkgGs3N1C4Sv9kN7Rq0y2/dW9NBWW6NzwZ2fyLsaVOLmYWN3s2drGCv1u
kzzBlUVSieXMA1qphUw+tftf74Qf4ullHIYpCjSziJsuarXZXBt1G1qC91ZgRe2LZQPwXrKtDwhB
uoIDlADCRGRIDJ3B8s/nxAxCQH4NP2ApBG3aCMUhO+DQS4Zs4mY4Yv301FVS4RSRswPSHcUUc1EG
ZmW+UBdk4R7xVcZe8X6i7OpJJVg4YDP96tlDmDlwy5ynj50/SXd8BYu+Kt3QQFFr9DUQ/LveC6MZ
fszjeDFX5PpMZ9prPL1RJoiAf7KpE2q8kdK9cnw40NIuskneLpAZ6Jgw32I4s6+sDxa++t1saXB4
tB8W5sTmynV89hdjF6fcEuhMsOis5VTdOpWMVVfwSTOxSuUM4BwdIE7P8NxrSIEHLsuP8BPydK4x
Unp6hoMdBUkXlA7RZ5lf+v/uXDfAZO2rjX9Y8ZPCy8JMXK08vHa5RIUIA9/lzEF7qzd7J52YWCV7
VF7u8QUV6V+N3qzda8SGX48r87hw5YOwTSWYgomLTK1fYwTXnmtLY0tS0q+sIUOsHfp6tdNLBuyo
MMnnkfuORck58dT9oDUtRTULX6vekh5rZIEKlPEBhZE+Kg/PFo0Y2lvtRUp4mBtuF1wSgxSMeLiy
tOR5IUjDqAZCLgcwukNctJUdU6mcnTCy3rX7WT+AfvF08hLhWB2HDK1+KCnCrt/VY8c2EyOUq8+z
YcOQeyUTG4UFdMoRJ5R+hPV75bKqUGKwd3KPNVjq5VxjH5uRtuKGwZFpsbWKcUHUAO2UkOtcpjI2
vfxqghwHwzC076OYdD0wZ6ml7rlOGw2zA5Eo3EGzUkN5VWf/Us/9eVPyLR5QD/uepOFYANptK9Ju
NsjOiR6Y68bsBMexFVsCxU0acLm9SUvg4CVlhQH62W1oQaCc+qm+2q9Hjw7YTdZ5IsDaJi1DRYet
0VDAiOLXZss7eyIxaecmkzvbYAt/ngNcp94qIgOuTMce6421dMEv2esVj/chaCT2IBFpwZqhEeFA
AYgU+0W1CSxfaymEUHMYGfXE9rNhbuSbMzZmkSYax/qvnWfLjXpMIhFtgAG70pPgWjaktMrAaFCx
1XOU4gjjf8pYi6t5TauYR8Ad4cHLnIiMDa0JeMncgrxlLiNctxPeA3TgIgOK2drlD7D2/xv/nr7Q
DmFHwLaKDzH40wjpkQJzQYRGfxmB8zOjT9DGhWWOxFrI8F8m+00oksx96TneNgjNUUXpmfzOIlV/
hcx+VamGGdlqVB4/jXLww7zIgXWTD1JcuPh2YWoCbEhZKLaLNTOFsAyZTHzjND8BieBoJh35R3zr
K0NPFzhsVD2XS8lCGYcdXIRWx/AyxTmENuZiFtXmPTMtCuhR/w/DJPgBqAmzg1sOrXyYxJFWnOFj
C27ZPI2rWHQMUBqjL7VVOhdv3O1Y2jqYgLbKfqreKLhEgyPZcLkZDpqA7QV4WORlcLVmwbNo20Lv
wceOk3+G7CH80cH6d53c58gddB37quRoqXdl/cUyO5FFcC3s38W3VmV4fZr4F326UtVhn/yn/9BW
csYDZUn18lb8DYgKo5gJ2Bs1VgNlneq/kb43pJqTXYVk7Di1pofETkCQ2PsjMjsfCTIl4EKnxvDU
xPjhwyhvPrioP+7dLlC6ZqlMl+wA/AJZMPp6ow36okeauXuB+D8rBTCa4GqfNkfw7+MNa3FpnIih
t4utsnGKb1fsIvWP8b6Wz+Ut71GWvga5LIdhOmbGr18B587FcVUI72OgedznjbjmzDiJ8eykeSW2
+rdqxg3XWX20xoRKzTBje+nmcrBqMPLV7pJy947espD00TfKrQZhowDIzHvN9cnwQSmFzFLPz0ig
lYauq5IicPqTHenyi35je1IQAUXGk1yTrW0F96aaHhZi/0+SwgdkluvFmWvdV0IJe//ak33tWpgu
1Vko5ldHyJJefqftzMsG6ymhfsSHkHND7tKC3Gs+BESHWZU8I5i9wRM6cRyiq9E7LArY+Im7chl7
yZIpgI2xStw2uc85Nzv2XdMZHylyFT7okitfwNJDm10u2+y209+K2SQcJC0TbAzQkONBzStaeLGU
nD41gnw2cv3WZJrTKX9xkzGjbXKcRFsdcPabbA5zQY8VYUujPhLAa+McPkGRsc5fD3nhIufgElEF
NuGFjExGymcTGdr/WwGt9qm+5ayM4CXMTfoYLrfTFZlcpt/We0wlwvvVv3QK6TubXHnNJvz2AHiI
xafJEgLadRvrlw+ML7cyo4CRDGkRY17BYr4I6PeuRPaB3XCb+xcAHI4b0RZ3AbjHPY1PlyzLid5p
3bqTo04lcpXggxd2ni/QGiYxpKPFwN/17iqNDklZ9yObwxTALJmly7Ki0SFmasBWJIc6kPbaJrnB
UjBbEH8XQmI/n3ad8yveLGeAfEzY5CPO7liUORTusMUE5Qmyy6yGU+HPJE31eWJJmcUVianM4AMO
anTs26GfFcCEQg1jUxcC/e0KE0DssmQHAzXJ+10x15OBIrQHGSTG//YnuLw93T4UIJF4371dxAmZ
8rg7W4QmccGTx5Yy6OTNM7iVrbdbu8v9FADQDea8LLfrmzZe2CpXPhAOl74VPXuq9OC0ekpWyxOp
nNzaRTXyCt5ZM52n6OHbUfqSFc3+RA6iZz07iQUhxyb+PCj8gCd+HShMT5kYup7FP+IrXd8AagY3
QFLIv8h5ROoOFo/ORtLWR8Ocb84lIsE/a/hsQn2UYETsijDMghKQ18HcQPBLeGqtoTNUmebBhwbt
7vJ6BSSjJt/RR1hxSOXOQeX87Ngr7NFqtswhJfGjRA0jD+WlBkAY7qnvfNigwHwc3ltLMbuKA+9k
YdR9/TctoWhi6vlw0INBU+3jZPQo7mFgUyGBOxHp9fYqQJM7q65ziPlWIUL1ulPuokkXEM6ThZ2N
Zt4o9ta7cXo3qH8KSI5GqM3OUEYrVLqLaAMVU6AoOWXUFsYV07VmAosgiWU5qXLtYohdh5oid7Gd
5LFd37vD+sghKqeAH1KFXl3d52Z53+9AZFtH07Kyv9ShKLSHUDh5lTmUZf9wjBR/Wr5lb3r9aywq
ke8BPtInMchPV48l4xs5duwLHmNEzQ93obABrNx8RJUMiJUmzfcgjxW7hHDoU3DGCsky/g/kqu/X
in41v/XLO6B+lcVSul3zWPftSCJj0x2+R4pgH1irk5tbVFoh231qp2cEzPVN9YC9cD4BhZ12H/pT
XlabKCF71JID2l93pXsehz9ml+NSF1KolU4Pnz5Qj7ARoGznS9kFZ7t2z4bpbaJkbLWE06e3vKFy
Sh9D2M10KYmaKJXRHg4syFrOjAFe+SoGRt8fexXSlgwuc052bCa2ybd5DuiRlDySDZyXR/ieQfcZ
XoJI9P/9r9zQr2ftv3xBPBIQ4jmztmwx+QDYqYLjjTIykE/8/WzSHr8krbKi7ZypYETx0IX0J42/
WWkE09p5yo2erK8ry1+wSbBaGb4yezxtj7o9UWruaLWHVOHTxLQKm7SEyA8nmaAxDN7cczFaqDKR
v6JRZSp3RjQ6sXpgkxfdx6Wa1SmH5JYb8pAmqVSMVo7SLQ4Lv6gkxPyQblshhfA7l696Z6dU17OV
BLlhGbA+tMSuN6s8DFyF4VqPp55wQFGLi7q7glkdHzHrhvWKABPH+F/TSS90b8UWxraDb5cAH2jc
0Mj3JWOlhzfn60E2e/XDnD9kI2VqGUFNTgBuF580WiQ8FDLdiXQk51Dz0vTUHpQ8JgcKLPfqa2qF
etkeo1HSHtLCXLKKJ2yUjNI4clqy2vGLATALIfkdAnpmIH7Hsq7HG+oLBsXlwuDp/mbujOg1b1+t
B4FqOqAsPZ6xdaRvM7x8pDE1AzcAdc+glj85vuBBcQfyGr0OJdaTQZBoYkYlo/9LjFSIm2S++eUL
gVWNfWq8I4ZYYmv6tiIsTKMItlZ6BOTvByTSZfL7GrQ+8lI90QzJ7lWi2Bo9hlr59cbacE7m1Kqo
39M5kiICAfD4B8ArQKQI3Mih28zy+ooP+OWDPxtWUDuWJJedVyQ9cqK6YWrk/u5Zs2e4twq697ck
tkIqTCON/hA8KhI5FOLUkiuGMbdo+zK+ttUqsyIy3WBcJvqbhYjRRbUigY9kgLaD52YS7wJCukvD
2iNvbDx1UjL1VxBPLBZt/MQJ2/5qOAUB2yFLe1HQV4D4LLMgOJMN77DMq4zSwpgJYbVP7fwgAqIm
/iIFQgcTEp9xXWZxtO+rjXgw5wDVmxm8Fea+5xZIY0pI9C+RJD58UVUfsvASiwblURUXYLAtfGC+
tk/bC2JE9L1oSY+sZfTFy3mUvfsitg5NqgAj0XELlUXh6uKzJpuLHhZFkoTu20o6by1Q3m5KD7II
6J/3CSmCUNcx1wbYj0S1B1uAuUjOC+zMFccQc/4A2JWx4ORjoksJD1zBvp7ZDT3eO8kuRQXdQV9J
XRsQZ5HDPRxD+ES0rFvkyhsnu8jOVorANFmcc4NEwsqTQGHnIPmSTUC0QSOX8Njp90sOkP2hhJJH
iG8ertjh9UKq91EQ7OJsnjiB13Nq4zpUC5QeufixvCTdDHDxZ5aHqa3CEnTu83+3hQIatcOsc1JR
mONJQkpU5bsjz3iSi+sRlSjNFcAJXtxi9Cg7JB/G54UF4OGjDCIP6cHoBRjDwdOHavpTbG47H+Gg
A+QKo9T0U6s1dBVzPv1dH76vpkGZ30fW1r4oHSqfe50oPLeLYEynYGf9aPR2/p/CRRH23uajcBx5
g84HBnxoBPAkUpX9qgP01bCh/Gf5HPcaADZkX2Ex2vXdSJ7pnMMTblpXPQ4nn9sVV4h2ISiC9/6N
39WKFne1AlkVBhqDRYDR2hFcfvfXsGVAiVIpliTXsH+PQYi00Y87DNfmQOazJd6/mak1v+UD9+l5
NwHJ+9+xARw5XtyrikCCUdX8bdVraaBXvUW9Uv/n/HaD1GPa/2JuzBu9MVeGb/6/jh3KLcBuUX/U
S4+BEj259CP2SB8xMhzQb4u+SXYVCb4TjPDoZz6bJdx72qyNUNQy8EYGO+PeWMTuYJY9EgHqrGFN
WrrBfUzDKuDwpJeczVehQ4xbJ1jfalrxaayvhzjapzCFAb5ZIQEH9lTdkJxCXolGYbHyNLTZOeAt
0cHnL6J8BLwyEVa0K1gBL5vGXMUMf6C2bkccmItWOiJmWKANtNYMJUmbjybl3T3EyvaxjNUFn6BP
hu3RMVrlMpWxz06KAVk45v3QiWOm1YWVeTcgj2tHo2Qa2sGIYDg+NhXFU2NoPgUPnNQn7r76T8oq
OY0h+jMPZu82SiLXXlIpoZWQh15BQcjbNHuc7UdgVEeQgkrPbQBEidquAP2poVac+L2GXGoEziST
op+C57BmG5RL2Gt+wUGmxd2kx/kFyDneJqqdP/1psq2JcX7kgKeuUmGAN+4qdDrAacNBW5pztnyb
VWeYysXjAxeVIOR4Om2yzkZ/JmY5Al66PHdhiZsSsEWHua4vb4yKimuFA5udG2hyjJAYDWW3pnPd
L4GK4rcZWJEwKNcDbhskHi+AouL0rK+xhX1wEoMVcxmbxMexVP/8ZPeaVApTeXZigpB09E3kTbEL
Sopdt8do36L7CGS+fhpgNS6YvU/mlvbyUdfHOyWVFjo6vhSo/6YkiubzqoGmRevPq70wd/8wSB6a
8apb3FJzDXT6Cpqpq4LmNUSzoQ7/H/z06L+FveFOjpMYBvqiU+g0Tn6/bXNdnyD5oEUfgot8vkMp
qtvEXeSajHNhXtLxcJYm9w5ftltaZ6Tb9PMe/Dyhd95P4ZMyV2PUrl68IbekSFaImkB/vK3DdTZo
5Ye5vGsfFUJxIwb9tcWTfbSxaFe12bJppgXDjThtIOORiE8i2MdsP0WmPSuKihTV5rR25+woK+EP
YKeH0dFDSXW4NtAl3d1IjkFHR2dr2Gp0yVj3sQQ7oii4mAwBYm0llrHGLiSsTq1BSdIAVb28QZfx
l4bDnUPFy2wQDdgcJDOLyHUNayn6kxh+biaLBqOgIVs7j4sTL041zIgtB1jBhPBNfIJBsOAYh1Ay
VyCIgfUcx55UgwMtV/YkYJYxLH5DtXhqWheZWUFvzbjyhC03noaYTARLJ9NrvA1rkNnmtpB+xpFa
hLQ26LUTwF5sRQ2D6tTg6hzzSZMpTWJbzZEdYLbcyIwWOHJgqPssTALvTvHWDFtPCe72u0eBR/gC
fb+PNjaqW4VmruAFej/U1Dln8jArADq2PnFWDMhqUfb2WVJbyrYPkoGIWpbLHmlI5Gm79kKQeCyg
GKSu0eSPTJh79lYuo+jlc7L3nFkR4ozro5CJvSU+ChOHujiIGMeSdGFFzqVhLtiLc1AjURamfDKs
dA3scKeOGH8vaxjaAZ6foDgSS1peHBpcB2A2MrxN+iDHW/bRUYGQED3sMHpVy+/4W3vS7HDfcTDB
A1SOK2LtuTqHRU5CvuqBOxcvy3j8REmNV/S1jjw74xtBf64/Om50UHPFaff6HRPuWYJFgDPteByx
yGjsZ7hwehtROjUSHJ7jzRodWOqOi8bp3Y3g1+7sKi3BkADDJPbr401Iw2wYEwo9eqfbodiIalg+
RDj5alVF0hOA4N/Vs8ot60pdYsP48MxUO+OOK4Z+BvTUNiT9sVJm+O4hQT9I0e2Fpu9/32IpK/YU
zEm6KcEHCmij4u5rdHU4XSFriaagimx+IqkxpvKS2bGvSbDskX1u0oaCLDvpdtbeldLzQgkP0u/P
AncDMrWEHStHD7fbFtdLWaEtLstoCASZY0DMnvE1dvqWyqElmEWVNiAg7ATzPTWCgpOxKCjQsE6K
4nJ/fxzEzF3QqAry6d/G4G3oopNgdOTxWvrPDoYaviDF91LiDwEHiNFS0Pcp7xzP5v9AAKRh9PMi
O/fhCOyCgkThWnUKoY0YgZmRdcHJgtpe7v1Cs40YJfz6+CwFXufjvy3N4QfMUHml5ketX5EmKCdT
/PO43EX0faI0VdyWT/45o1QJVrv945AKFagu9mVSmX237xN3g62rPRCYFPi7BbOcjZZKfELrb1QV
s5CG22ZZzB+PGA/LQojnjyIL6bzbl2uFfmQPaFhUIGLx7JsZHvB2tnb207d8FY93JYD+x8CF6UFj
6X4IQDrSwgbe0ifWXQoRfiyI8O9GOLfjzf4q2dJ6N4jRZF6Kk5fXrnQBpbOp0rMaH7/m7uXfmguZ
n3EaaydpsSAwUzazOyxY3PL4ShgJia1gcwK4+8Sh1pkOEBxV2yDAltkz3L75eRSAccIixlzFEFk3
elr+XDd+/2PBQILCGxXK/OPz94pL3XOjHhCriJ3/J7F61fPnw0mljWpF5dWu0qEO8o+GW4WXjOmA
`protect end_protected

