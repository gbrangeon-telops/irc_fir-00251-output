

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
e5xVIDBGzQkhDoQ5sfeAF2q83P6A1Z/qsmlSYQJY5xTravGd4CV8IrniJyUa6zNomwm8ijfsSBDZ
3Cv5fk91Hw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
JTncam9YaU88Ye5zsiMSZerKzQZ8ndV/jFOlVBJ2+1NMrth4ym5MZgOOJUn+hqDs7WawEc66qp7n
dAXASYJYn+qFnCtyUAhIyvGYbamoaDWo5Ex6WN67wq/uxVFQHJyQE9mBWmFUuyQbfWAxdn0X8Ddd
XBKhuVWHjadjfvTndGU=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
WysH5jibOCiuNoaEF/J6UEux/f9qwkqszrQvmOG1LAQguVnzJ7+cmZtEvDLaeM5SMkI/c6AvWtXW
QAEuUSUqI7fc7s94OSdoy/EO2eWxzu/2PZr3+Vm/RDQkA2VgY92Mk7iTSAe4nvupzjwLJJp7MPFn
W0Qp6hutV366SMmocbalqT6lFUEm3BdJRb/waOPaQXsiK/eXFOfDC+OkXBIeDSI4U6bTS5BbTI6J
pFf7UmKKQ3+TO+1O/Q+2hW5WOgJzIUFjgYlL/k7HV9GLoiTkFeWQv9D4PmITDLLqEoJBQEH042D6
w9tSjJ90YaeXyJsQBc944KHiROaj7JIGL9ptSg==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
HfnNrIheX+bmcZCjcmnXLaiCn2W6T6H6Dp6dScskVGNGAylFhqrXsMMXHrPiUKf5LFkT6rGH4xNt
DnPlwzwiCAkQpMo27mNuJmSmEL1NZn19+z1IhIkgUjJMK+DU6V8j1HJvLoBzdBKXeOfEsIha7CfH
SYvgpUYxukUrvYeSdDM=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
FcdqosqcEEFjwfToDdg81IlS3kR13BUL9UoyGE7K0tYyJxwBRWvuEZwjlqyLvEdW74UEcoL322wG
MsjKrbrYQdHQMnu0VAIvQRAp+YUu8ZY/Amts9d4uoKQ4ceZKPNKKjhA2gLCTZlClOnHdKjhfnFhg
C4vFlIgGFFvgy7hYPvMYgUjBeujuUeMJVrfDQoBe2vY01NCaYs8PD38+MZrB1yBWXtoIH1Kudp5s
6rfzNC3iiU875HSyCH3s6Fgf+5qupOBLk1FOGYXDOgVB80WiCFsXlSgDSubN5g0HTJQJ5d2+rdH3
3+ADIpk9sqzMVdE2qp7yCA7kfUMNWwWOq2rtCw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 15872)
`protect data_block
6DfID8Y4XTmaaonW01o/A1JJE893+DRvospUdsjHTAqkXL4WdrS7o57Q6CLOMOcuTsdWznqght3J
j1SqhbzweeCi9cTOPZ5N9o8hJbF/Fj2wCAM92f54voHhg6NGSlvNdAnYhdNLZkBk3jblGm/HKI7i
2wS5hpZjik6OuokmF6I2BW5fZCArSldwbC+gFatDAmqiobWoHSExTs4Xf/rPGs059Qip17CK5WAN
Hw2cPaEBfDRpV/cAnW9hncZko6skS6pWBe5GnKapP6kLhXr+jNvKPw7uE81tmA2OyNGfTcOphG7H
1OPXk7ocFHf8nEfTMDfhpLTmmec2028qvSGO785xJmF7blEFzUt7dltX1o+kNjgGgk9BXbgVGLi5
akG9k3EYNTgdr1JN3reY3gtn1y0A/eooLyZLXBijSyY3u1GysMEpvrQbUDdibp5DRKaFT8hJsmD4
mUlDh6usGrEugSoSy6f4ybkKFNM+V092gC3iUSA4OMMlI9V5xfr0OjGrHENY4tPSnKe14/mqyWXE
+/3UCSV4F/WCbtpdwt9k2JivCWFjhIcwv5H+Wq0VjufCrJU4V3SQ/rU7IrSJ/quM4id2b+bddFq/
CAxoF2jtc8XSBiWk2KvW6XJKbzynWhnW8Xefcy1lKqxrZTMG7hFAosikw8E4y8ohYN8/XGhEFPr/
UWjGpAHs7G0YkVF+NSGHpUk5q/hS6vfvqkRGo3N8nPdiPtj1pE9IKgJv/w/z72YJ8j33RzzRQvgh
GMRKqpwag2v7vMQwySy9Wr6ereKJU20zVg3tcw+9mBnk5pquwi6ZAUlV1pb0mJDPbutX/nn23Eix
TovusYzIkfEeB+2pIIVWl6LnmdwK7NCETYbaDEu+Ek8+L2iJdw1TLlQAHhqJCui12mCPbFwAFRa3
3+50IbhZPV9YX+TcTOlJfJRX/kYKuSHBZ3dM/6HSM9EelSix3r9Ut57a0selOrGVR/hy9DXbQC/w
3v2uTJ+UVr32oAUqS/O8YZJDrC6jmPXg1pXYl1jLOGVui1VpOTMhQKzXuOmBMaNeEy/NA/dT4Ru+
VR/WiZTdpzS8j9VZ0L8Zo2WA0WzRJK1OpSWPTeMpRa6mx0li+Z1GU/oSmR1ArbzZfoZzMtc/ZvHm
KPxGqfrfYU+NLTCaGwbk/bOy/qqohaJTbDeqhTnW1J2bFO+7jOevegYo1A4F7bYHiajbf6c6fIoU
0F9PlDnwBQ7rWtBa2coUpetUwRfpcrcJdy4bOujalBf8PZeo5vnq5ENmshdDODr34U3776xszgp0
qEx6jF29iMra1OaL4+wIzR+7UfR2s2ct/Dld8JXRQcX40YU03tPUYC3bJhmfDYDvFvp7AWZBa5hc
nUt3rkzSWkNzuGLg0mdo1kj7K43BYnSas/PsO/u7KCu5KgiZEYGQD7aqeDn3Hl3vhnNsqR3LdbrH
Wu1Z7K0evk6ssf9o7hB+LnIpUGaTmPZxxEBW1lbZ88DohH/yqp36F77gWn3BUnFpw8Uy1L/Oc2u2
NTlUs3/KQ85iN/fgMKEztyN923/bj83bJFmnwZk0bWiGU8kmDAAfiR4/l+IUPIRNgLHES1vlqawN
dYdLJySl2rblmTYa70YURHOvF15UV9fcg0XS1tk/itkTgb9TKkJXELXysMhf6mQP59ammyzkrnFm
8HNZH8jeFS1K2OI1A6pOu7X3o0Sio+qS4PGHdKxxrfyhcBjBMJ2tqb+YprxhGZKQJfVE7FUMIuv8
QURb4Kr531Fur8fyAEoSpE2zAhUc1eVonfDhAw5xmcWTtxLn1/MLBv6rHKzdSUZxgXG5wuZtciSO
yZMjN68l1Ar5LkaTP9Mob6yUOwHCduQOxjMpx/dcRqE3WFZ/jWZzmO3SgsJiW1NW3Gg50DcDeG3K
w0uH+F+1UQSfi5f+QNoNkeEaFjFpwVZhJDP8UiW0zIWnRqEGKpcc2LwU0cnWdirLfFATVtEec+zG
6hIJvbZe74Nu9HtWBhvdZIFO6/Hex+HtxyIfjHJHOYFqlDKv1f1CZPN7tyosy9DwquTpgKHdZr0K
Ftu4oIUS/okFGfO5PKP3UYuz2XLKC3ibkIGQJA8TQEUFfdVLVQGLl+A5cmag7CY7UBVyuzxioEXS
IyTZpu2pQT8cwVIp981WPwbvmn751zzlhrNYGPTmgCTXmgHBdUdnqvysP8l0G66klvuAY29H95vx
HaVv4JMM2/KNOICsYeZPJSeEc0btBJbXP+YXqAq16b1H51R2pdLst79wtr8TmPxRmjk/POMMGSCk
lgiiie4EaUy9REI3IC8Q80a/+Ket8pYbfCj6MFl2nUHBOgDfKwa5hhEclNuah0vypgi/MIinALBE
Yb+djE7hfrl1EKbdVyuT8oTkcbTne60BvTwb1qSXxQQWSQUVzOCLIG8gZdLOqTRlZUzrP210iRFW
QOmfI0b8Zvx03w4GoORL8vCLuZkynQKxFmxlTlwQeeFFaqLPeLm6qR5gK9DuHXa1z1Z0S5rs2bj7
Z5IzHTKBin97P7HVhDR18o78pOGIYSKSO2r/odFRv9DzEeuNWuitH1HYSQnWqlMMP3kk7n0CVW6d
M0/CcW7BgrttwX32nPuz4EjbMxPr+0Gqf3lUSzPmCKMDS8qMa4bC3ysmox6a+ajJwKaw+4tlpJpk
npwFasWTJjkdlNY6u+mQwxjT3Wpm0V48wnUP+Ut+YE9d33klH5C/XQcox9KBwjgPtrhMc8Gfyyj7
DpuGKmP8PA2irxk3q01EFz3dhKNcGMwB5J6lh84fUJ5s0b0FAhK4blrSJ8plvwVQZqzY7mbgIYH3
i1/cahBUTfMNNVE0nyMbEui69xSISflFPNOXA1OsnNNvq5ixmEl67S+gADiZkDZ5ttRberU77O1R
anMV6dPJY6ZyALoe7cmqXLB9RRX+dheQHComSk/zh/fU0pLc242MiTbBoQuwZd5Zj1p77pXRq826
OY5HJKROeVuC0GG6k3mcY0tBkAvgellYKE6Q4l27PKTd/lsI3AGpQNq/ST8qbshrnad4yUttsD4J
ASj6Q1DVE8H2g+0BBmo4SxN0CVeM0Aqy4guUaFNSpFDx15z2qHF+FO82dtt+goi69ixt9kkxWiS3
zlFF+yGHq4W+yGNfuQsDHgbO6ccW3u4uND3gUpV/EPbFIqvJTOGe6tiqwCMuiSHrlAK6PVXzyY25
SYYiWQlEtMuFjxWDWE9BAfBFvHtA7BtwqAwvqgihU1yd+X9uJhnzm3Y1R9p6jPgkbYO5ya5vibgF
jYn2YKRumCJXx/7q/422jiwBeBGA1UdiChlIvNLJXqu5qpe5HoaXxtJSHYan2Jr0YMQBGX6ZSXax
m6hyWRiP0VS27MkamalWtpE5B+t9f7dUplfPTlmGnQHigux/uAjqMNzwSgnm5GG0s0klEiS4qNe5
ChXUd/KkuWA66E8Rs0mTn9SVDNvwEq+NsNvNpgi1lOAZut96vlA78EprbQMuTm3Xekw7OKCaIlHV
quF1wdTOClIhzk/WExoac/hO/bkhTtjGhpxn3XcS2c34YqpM52718BT4Foc1Ef7PlNFe7/UA3leQ
IMHiU7B7tIXz/Pn9Tkhr4xApWSvjThAl08L8t48hckvxVZgIv2v5VjtlYBwfRT919Me014dURJil
dINl+66jwVzHkMRz70J9KtKenb1U1cSevgTYpVxBxnL4oR45JPLjNnpo+9xFtobQQVMXGWJS34Id
0KNPPP2YbU4rzGhBC9leOEDccgBMoHnGXiQegy+i7I/2U9LFNz90MbNuy1vnNgjOuSgTeIFfXH0v
WxCYLCft+UlP/rJ4KnkyujTlf3AaB+nAsbDXSsfRCvNPEKrvAcZQDXRjQ57ocRDHZJ67k1DOu+2r
dwsVfGvCWBbPZ3/hrTMuvAEQOZ21Bqpvr1tsBthNx8Lvew0jy7woh6JN8z/8gSGN8ykCkETr1Dwg
R3+dg5NZqVHwLJwzVPsgYjEe3U8vs2qOFvdBvJ9NvOxDsJ39rss5l3YwaTq8LHnorDGZ7h6MQJSK
J6NZMmzScSBVYzmqS+zhEO8AJWHpZP7l+EQZKUXgwZxkwXXpU8H6cpLv5u61b5FaCKvZmzf8kEYY
9lqcHSdMpL/K9ft6K/Fq2NT5fudEjbRLjtTVpSp1plz2pazaR6ZaTzgx2kwoVG0n8U9U4amV1my7
30U4RagnW0yTiXnV1Qvm6j2OWr+d7BWGSz5EtdyNXhTJAsK3Yj9Qazyl+ti+0bBiiqrUQREX9E0k
dfhXJkKwgIVY6eq+IJBe+1EzkFuVzFZe+bFtJnGvO7fPI6UODFbJ0nqea8PpXKSZDpgTX5Sk7F4+
sfWbP0urMYLgI0YBC6pj1lNske8esz/ODBmtiruQtwBB7mwyge6gBYJ0/95ZWDD/vg+kf8ZoVOHK
2qNmTIh8WZU/m9jJCyOHHZErKoQoolYX5/zrhW0GK3hCRHRZfkDyE6jme7hreL07/Dwj+63ND2Uw
jsnB8zDu2jPURleTAJ6/IHcoK9a4DdqZ01+oDfUQ6noDJJghyBynqmE6G6j0g49e/tckRWD7fRL+
j5ddkXeFgNOsfXxKdoXuKK0Qtp/D8vnaHCAfm5OcvNJmZvKWRWmXBLgIB63wY3zIYqj0dgfsveAp
3EHVx6AMeOdqwsoX529HsipbJiIKkbdkEyFO9zKMYk1km5JQKmhoS+PNwdNkjI2vHWVLWIOBiCWJ
X6GPfB2uTvVZA4emBtrUKe5PhG3Gz1rT0TnoXXhq/ohkEPmb3KW6vlI+WOBhUUtyW1xOwkuMfQgc
xXvupXELQyTQe4psqfLGTNwZ6Zc3erH39kxPhhmnQFGrIuVJlDa+1c8bOUXXfxaOdDlVCiv6RCbo
KJKTDKGfbJNEYlHq0l5gcN9svyfM2YH+pLbZfp6kE2UMRldr/n1N/hyVhVJTZkfeTgzxwZFN+x2M
iqnntSM3rc91XLdXhJcJWJ9KHKdR9o4hWwCnmhAIvxd3Rub8GW++2a3SdvqtEMZzmbUnjdou7Jv7
mfLYB4H6vwjBnkFNcS3ip8RpF1hLC8IDnAb9iukOrjvx7JjXWW+CcxfJ933M26jKec3D1o7XD9Tf
/Xs0LQ3GRl67IUWs+vKd7pJxc3A6vZqK58T0C2cBCz01ePkw4bUdgiH4V95c0KknU+kybCFiyNRL
aoIw8Z84PNoCodi/uQUMF5wusKmVPAlgxGyw6yhmepuy5c8bJvDlqYITvHMLKaSty7C2O8ElhI2e
qyTdlBx1hYoJ/uBtbin9/gkRCH07AvqROYUzfrtvkwU49EAqbfIIlNLtjd3cdYA4Eag7IChkPwRj
tpzDAVxwAOnTCx2rmaGwJ5sgiJd1+ibDHnTFKTMrMZtDoRahF7bSArRpYLWfNqq5fvqDMNN5dh84
WmYmKfoETzb55GhWx8P+qvCiRBkt2Zm6jv3jFzrLchkdWHNhmHoYGAD7pM/iRD945FEFnKvy7oI9
4lgjdnKRx7PKl9K2m2bWbU0wLJw+7Dmut8T5qJYo5NJH2vQlZfgxmlfjeNrbfAcAO6PaouQQc66t
24z9oxNbJXCzNbunjlXMsmW5JoJIucKTH/LoLWS1RF3kQpDZMSqhi1LcswTonT49imy4xaZ4MHtk
kbh6RDrdSM1VTY317wfEog9/ViS43/+cqcCKGhEkgvbWcAOq+8ATvfQIemIwer13vHIyqJmLhwLc
Fx+P92Mq6jpJ8LRcG33sCP4voYfbPKb5y/28bH+ryGfM6WFtKMMuKnvEAuWdvCTZDJeUUk2HjIA7
7gmttVVBbx63Z/tTQz8A7zUVZF0q9ppmGRxaU/T3HxtKELbP9rco57V9XXlkyKJ57aRWS1h/mNIu
y3I4yPOA4YYBWC6z+i4XGAZnh4a8HmCMDc7sutJiFjZJ6HZDnEegVOn/xH0zYh3slgJLI12FMHO7
rHl7PQVdKfgxWj7BK66Bf0NfkEpAjcNHhp3P2xtUIlRiEyReuj0eQhhfrAiWZZePMUKH+33FJYjB
zXoPlXxZ8eBVKq5W30kNFPclxqAgHpP/MFastJwan+BtXg7K8UFqHa85gMr/Kp5ecMc2sr2UW85k
Uf83ZLk63XKHqo87z/7dzES+Z5BjZ+NZb6YleZ8Hx1xsRc3cRYeviBfMjNcIlsAjV0IjQflYnvJR
JbZ43vbK1tTEiuGU+Wpc04kgarnytTqsbprdcPdW/AlIRqFD1BTY6ksqso6Y6fk1vLsqd1z+7GoM
1AS7mK1lhEnxkXMmDkw09bYGEj4IFcmU1941zYeEzbDOfsp1msXq/NRRPmH8lFUI8NcsiOdGU9H0
sBlA6cBH7WInbTGxN+nB5xicB5PPy6nuwZOo8we3ivGXXZvUo59LRMtfI4dziKoA/kixzw+2h9EL
lUjz3v0KHNkQgtcAbdqiVUfpoMNktOeYWQUlzIzdFWfzbphuw6i0up+Q6hUQg/dFdYaYNxIe+EK9
+QkDWPsVqwszirEtlx8KY0VFhQ2PrKePPXVLGFFml4I7imsRCy24jRH4wnN2oqTMq1MvMz0jfAKO
2UA6lcS6oV6ubufQFXsPRm85kb2e2rlUijRmMHqs79HxLaDrBKe2IK6qNfF1eo3/6OKZUIv6WQQq
F2cG9jSTmEynvZMYbYOLaIcZj6C7Yaw1dVoSCnRaOPIS4FLoqDDIBE0dzPf7w2xUJYAm9tNgSCk3
hIb5+DY590Csj5+KMxwcrn1jsJBKHXaLzaMd25CmeVAo7SU3r9Bx2EH7KdtRXu2+LVE3FZm+8utS
x6pvr0D4ibpSUdB1aH63vpbd7F2O0oecd94m2sZBKt607FAVGuDiqz6IoWBKDfupYHH58TPa83Jc
XNeRCGA3Zld1vApWEpY97afH5neJs6TeUQOA0B2tO/Sk+mHBzP3M3Gsxq8dHJl3lozg9EOhqB5D6
wykmytxDAnJSF+/ZTXM6UT24vs4MJTNy2/GDqoFoBPIoUUOu0mnHiu/cbyjZSA8pjwhN/OPPPf2E
SuMWSrkyRZgOtk9ojWlfdDef7bAg7rQ2/hAHEFmqnEc+YmL8d0IzOc+amzovnR0PNfw7qtcpavF+
H7UibgifeDq2mNMjskNIvc+UIjJuqgJyjFJIsecF1dEuUw9bk1nKHhAQU9vjF485K7zThpMjSyHM
Mkb8QXPuFSxgUaNZa6QHML4LiTqzgTzEuiHeaEgKMwzTSw8/C06mKgw80j/ONFZm53B1f3eSOl1o
tTc5xqKKCe7WAxIL6VJxDGDqXjBfRYyuKyem7VKUehnwwknPuB6MTrWcNC7KGPIe6/DWtr5sKVRG
/XdVElb2OnVi8B4lcy9qLlQJcL+NNGsnmHmUdLruPmK5cck+UhUlpmuMVaUv89XtQDah0tmzoAxl
Di0o5Tgxc2LT5Cmjhp4GWDd2y4Q0t/T1vI8DwjSzap5p0KdSMT3TxzjEFSBao39LKWDhnOjam4cQ
riuMnX5LKT7GcUUEvSkM9f664f+byCEKme+bd0VF0GOCTdSvyaMpxPijQUD9TiFs5jzcYW7tJd3+
vw/Fr8XG9YA9fnCPPvtV/vd2kkW2AHHTcKCT4EDojFLABoClfxulT9Pp0g2JfCB6fk/C64mC5TbZ
nxpgYxuzzWqs4OL0thhluTWOeyNBwlDbC1k20Lcj+TqXpGDaf8QIswD0W6UKuG7278fT6WLy1Eph
6BsUH6eBthPDNCcz1ZOCXzdu59b5HLQHVclwzzjAz/pkI2xgPy7envjbwwNSUhYuVPz2UB8U57nV
CI2k+fO/A2xsWT6IW5+0TvQHcKoHUiTpTbf6iPe484kdM3wW2jEjADktNITYWpGRgPjKpLNw8vnr
FE/XVjVpbjNBsxibKFJoGgBS9ltwQslmDJ+x5FjiOQsrQIv7oiGWEK1t0WmfAlFUd6/Y+fBkLSG9
IqWDCYocHzrf9TFBKGu8KpheAgRR6jfCS0I8VACcFn/C8GssTMjzF5NU3GqG7p1/3K8+LUdq5E1u
0C/MUydP0ckrQnbIYqfqvtkQlp0ObYLZMtsg50hZHpcv7O80JU2xlekivZAA7fO9HdhaZB8jqUkj
EZxY01lF70Ch3LK6d3DKv/zb8PSJaS/aJeMmcoCk0Ci4cDMRIWfMC6nHW2Uy8uqLjfg9eBNxlkUI
uK40aBcOXLFMKOZtdrTYZH+HsBWXh93/ArJvBTTeVyshSJwpRK+W1TEPsonNEYyzxjhfG7bscVJP
t6tdLdHjEW/OwbkUB+WFmsQk9BfLYUVuq5UjQeJm+2k5XBLTl24ZyX1NgQN5GS2wYWVIiaLqyOjJ
xy/OaMNMQt2XHy9fotvFkeU4wAQS2H0nj8vTaNL9kiDC4UtPKihLv3DJ7+IxDtZoc8p/0QZmYkKh
92+7T7YaLrvunMK/B0WjUI8WZCXFbmdtGhepffdWYOfK9GUuyaQSS/2VxBp+xMBAEQiiN5l4Oyxn
NZPSCQKcxEI01ETBkYedeGoPp8FUl3FIkjIR6FguXXxZ9EkZLxsLxQN3v+WnwTd8URSjnktS84bH
49hIDN+X22epW59OJqkgPjb3N7ZdxN7o8QcvJVO4Mwk2OXEDq1kJEm3pMvRexsCOTB9bPYgyEiQq
+q6KrbUMEAYf7L/Dh7XcvEJGs3m4QHuR+lrToBSpVt1DwRi57bZ0MdRUhwH4et8h7eMBIc2zzGU/
BXbzNI45/mqslebT2Ds+7ORfUvYgqI9ZOYr1sPqsIU+ap48O1q/4fnjUhqafNKayOJ7ytaiXGZJt
WIcgFDpv8hE+wOF5mCFWQO/NN4fzfsviWMSdPmk7fMGx4PM5nu+1rNIG/A2w44Ks47txUZPZ6Z0L
UvEAB47HbsqGAM7sOcAnMydylKZlReMMylRANvz5zh3PginhuX4L/2uZ8Ni2NzVaJwwCpz+yrBVD
fd5GlE532+iAlt80kJdiNxsFg98AtxDrnStHqGj4+whSkX0U4yqsVfkZfa/MNbF0sNUPb4Vc3l8H
nleYRcpdA7+WT6C4Kv2J9gYDQqQjupce5HGijhXmk3L4ByZ62fJ4AznWZDUjZDBt/myXq7GM5aen
ta1h2FTf0MkTcMlAiDElEXDWW9vf7m8uuIakt0vbbs95sSA+zl6JEY7URbp0FjO+XOEFWFgqRaqf
+YLoysMt8Drmz/UHPH4IYkTlipiKlIOPzmbUs2/sBbgqsAfYwM6UEh6AYvzYk2ehlyxsFAyyaJ0E
3+v71O7uqTgV8dC/qZdaiSXKqxjaGQewBNHeRPouqa/xCQmKCQl3RLv/t3ugsRXF+HK/Q05/cK0V
k9y+yE9CMhtk5HUmK+nj6kiz7YjxiYrDJmJxREIZ/WbXZXR57r2loMiRZtk7Uiqr4BMRbWIDWs85
4vTeA/JFlDZZ1l3+ZOvZ7G6/UpeF6Wuy3UPyGj0NgPDXPdYWwn4GHUtIvkmFOy6fiIZIv3toVoGJ
cs0M2gqCOGSQkwAW45YXRvM0epbZzw8aOJ8AwLrTz7VHbFD5DSSCWko5RC/AjDAr4V2/wUVAYZZi
lkuUIR8f2aU8j9ymI6zioWoqIcxMqK6Nt/3gjkiXwMlUCDOduWqyML6RFL0yGFR+UZ1S/o8Kyn6p
HOwQ5draSBnqd2S6/krQuxpewwAnITAxuF3jPGojoPyENoHie2dZ68+9zUFTCyX8W28vAqhKQL6F
EyhaxagcAv2tHn6DMhNax9UfgNpTtfdrIlXduJvfUaDEPj4T+Ye/1E/7w203hGIaZh1VeG9FXExH
icwXLg/TiGasqNX2CGxIc016Dq27r8+kk/TSbTorg46ANhLtSySTwppwhx2NT5WbczEoSdySTyVB
/qZVaxlu73G5GaZxNDWNkGnvPv0zBd9QsKaWB6UOtZIpzdQIscyA9lIcfxA/GVwyGl0JpikP/jYK
tODnr1MBCC8M6Sbp4wEksFlmHo1Isu/75tUDJAjYnmjlAToAgBb4u1guc6W/36DB7HloChiiuSJf
bQNIx/3OREml/cvWloq8m1CgR8gmhLP4v/CxmCoyKUtog8US1wievvU4AL0yVc7XHg3o0TyjENsG
mMxqJUg58iIfS79ww1+eGhWVHcDkayL+pc/XWEAviWgJrCn0tmv+jYJofjgzFJGTmm9amj4dRQoF
Nt/QO3XnV2MN8/OBOtrP/IITayKj+heLkzG6YsKuaf5I97JAuXK4dYL8AI+ggSi09SQKqWgVNxiF
DQetDsaPDxExKZBuDvTy2Sva4op4dj1x78gYGKwCFb0KODjW4ei7fNlosUYNg0eqsEbadMrZm8Mc
p2HntvP70BR1R7DL03FBXX4vdEMz75PjlXHV1G1LGnALgBUW7CBOMeI0zF5XXf7YL8eFEbTnWKPo
gRn6pT67Pwwxt4H0+owFs9TtsbGx0/7RwOA4i6Sq4GWtfGIJHkTmlhdjfKY9L/HxcoWDckEeaBgg
mjOO54zwwvBXcyaLESMUzg3njG+kzp3N2U1cQrtlzmaHajp10ofvRA5F+zyMXw2culzC7ro04cxj
BE3p4c5aswuDI1SMmQBr8OCCYaxT2Upk7e058c+hnfmq7qr0HkUXn7mU5OSYaqdDdKwSaexkRLUz
PLCUnxvwgNrNUaxqer3AR9+mOzXOsHunhVVBJyP11h9LIMgAarm56tGlXRzZNCjEzUphyc+LHRkj
r/aIayI99uY42pkEWdAICYtG4M7u6izHWg9AztE+fAtpC4yfzam3mH4ZA5na7tZlipwq0rfY66sH
4RsPW1te5K4mR1mXC8xvz1A7XTGHmSpILBKuTCu2uc4TqT2jIlLaLYo2jjCfxG2c8tmdZCeGKpPO
aRlPdcY5zp3wXHYhU6r9Q0JUW9URxpZli874pFkbCk7Uwxj9OTmwtteSiVsPpyrmUfmQ6edWePhe
85ZTse+EsVtgKvvF4BAn09M83UapwncxPCAVOCnqgtoqjpidp4sMgKhsKrOUzd09oipd8agbPI3q
UvV4DshYM/x5LSZbEPqX8qqhAaSZWK0UEtjkd1BV8W0Yls8H1TSkJKn/x1abcZieLD23kHSI8IVE
qp32KhXYbA3MobBksLcJ1DcweSiaKSpc7kajaJ+qLrEdyUtiew+egjFuYXw7wAyAIlluW0X7hySG
zmemQVdwspwJ7ykc5vYp8/TuIEADRg1tHinWIjil0KOVfKBl616V3ZR31Ae6aTJdqu+j/l88FbtK
z4KL8nMu0JqMNK77shmjJCuLmYPWHQAquVWVtDhEQsjxwzNkQy6s83y4idBthc2V7BW2CKEisjgI
8nwdnboijnpcKhZ/cv6Sb4Fn6e/WwxzKS5GbAVhAH2Uf/LTN2CUIlbgo2jeNMlzvlYJ7tYhagY1e
MU5Gve0uBfr2fcn2sZ0HFmbcwvyQw1ZnEz6JiNn8wWObfz5Qtg9Q/v+DrT3x9rr4U2sNNPNeBZ9U
u0b80g0JLGgcEVi1xWjVIhefFovlI1luZPgRWjD8YHE3vXyj/pB15ngzjW1w3g2rptuU/1CasEbh
/1Dp+2vxgswkcllCBBl9KSQHriqPPgDBtrHQ459NkHn/suFmeup/tav9YRcNhDgm2KS3e8K7khCK
K4ga1a8qgDYCyDIr42jNSx7wWMh76PQYAFdZ9f7exI2pDXzCeE5gN3DTugXHeuHXxFsKfF+VX33z
LVESbwQF0XbMAFuGrgUFkcRogfZk/mFHyQARTT/tzpnZ0041yNYbfeqq8/caRF5IXfSLQoJknuVE
FqhvRLmCXZVQ/Z2qm7uo5BQuYNeA2EQ2h+UG+jWFjXprwI22Qnaz89MBDygviCnYyiMC+nIFyUE7
QwLNshGd+BKa4zh9sZV89uIivRYxV2EEZXC8jJopfABjpIQfZck+YqSSd+de1zAqGmAJtyARPLKW
TBJkkdSFSFiiCYnvZnBtX47fJVqz1SGkywixe1cLL1Ik4vMRnKxaT6DFK6Bc5ZhSSpJS/t/2TEsQ
NUNqkQPOfw6sfOC3xEzbPgdJv3DMoo2FdIz2foQb2DlVanlWiGxzZ9cHJoA5M0HGv8K0lngQXN6U
4dCZBjF0/AbLovyD43mJjCnICdYGIKGhns2SRpoQdkcoDtlWcwUYKeUGaMPgwQ3USjRwM43RqatB
ZJGUUfSZKPFQEMKchLIonjOR8nMPSvk+ShbrHSQPq4lHTXWcTPCWirtOTA2H+iBJAEN2epS4RQaa
tqi4vX4Vkx0725dZgFzFav0l/bevRGi/Cd1dFaoCmHqu5QdlZ5L3zuVCQKRxgSLqIvoidkjYYoIt
50HxRC8c7qbRxGiAEpwT8cnVDpj/yJ+BDqmjTC2qt3mLIZTY8Hum1UsrDY5GIiBNx7CFHV8cnaGe
r14sOCfIZNd68WEJQ5B5PNtgUHvx3BJsk1ZtrJF0p2aYtQQ1cQJCmpKYgifh6DHZCL+3FFupXXIz
E0fHgKo4mtElQRtAgefgmjNbFC3PxSu7qDf5bJRaVKlYDq4MRDbkQyrdxaVmgxjFURlOLjQ8OjUj
FphwEF4Nrqgu8VVeUfqe4jXsud0U/MxjW2CPC3K2l2OufUCrjh2f593HRvN8cT9ZMOLZ5IOOeBkp
j7gN5S+WbWMD1UkMxGnTTS82ZjEBhR1UUssEYQU7AD47iGR4qGbjbQhXaaVjx19zKmSOLlSog0g6
Wfo37FDl0iE5Vv0XXweavlyZXkbA6JFz+zph4KEQUZfbUx71xEAV/1B6slvn7rlidzWDkxM33Zw0
NAwCcqojh4xNrAY8PCZQCZPUHDkKWoEtNAxeiTEQBipGzkBUIdhOeuXQXXFaMIG2KRob1OxXBZ2M
JGyW9VUnPsDRgwHjj9p9X8zc1SF5lNvJzrtfXK0lbxRJaOYg+knlxJR0r0Yj69sMXvU46SbaD8JZ
jMDEf7KRkFzKkmsoPlpEOYw6ciFKx0cARztvgwjgOi7wJKBfMoosuMDVxdePhwavzxqErm6PjUPe
1JtEK8Umhv/ZdJoUjjkGz4tPhkOcZCA0KRrnYo7D6PokyiGc32T9FLg3zxvJ1Q6FT7H/2Vb6zdBO
LGu574hO6nNAjBR4vUatV5CEb4z51XTvisbFYYBaVm9g9D0FTT5AHmWufiaf/SVMAyHlfayoGi9f
RMqv+aMA+/MRbkkE9ybXeaJ6sbqeDCY78FBF71QZFFxz+HwXBA4/LRdoNPBn0c2XrHaiTffLM2PD
/WGSRdPATDjRglDB1CUszcV+tBjhCjwLe9NNwM/jdqKm8/a5UJOXzBJU2OhwRFRe73FHzDuY7BI7
/eyIssEHyT5RimnPQj/82CFoMpnrUQ5l49TFdxlJIGUye95odtW6JGyrlQpQN3buKCi184fuvtiF
2YB0T//XsK2jzZUZWFN+jxO0FSS5HqLg11rMCUYB7lk/rC5VPG8JK9ieC96dNZRFoHyv/8Nkew8A
oR4l721fAoAhLA4GL8/yT5YL/nXPm/aEkP5QIe3T6gcmiJZrP/KILKnsDVF00GOzTtppeqfcJFcW
hkUHjzK/NV4ae7OMKzS0cTC1mNezr8iMwPDrAbe2oZ3DqfTHYMrwV+QurRReUHAH+tICWmQwf/Vw
tUZLqUXJ1IYmAaGQpGPnk2bIXKlzTHG/eLR2oBbFpwTj7UR6Gpm9h7UgsM96I6DZ7SOGWeIKiHOz
XJU4g7Cj0SLPFcQj+5Q3VJletlfEa4PWbXOf4lMY/+hewkV2Nkso1ua4McIEYx2ZhgQo2ZM2WBMy
7+RHwxgX+C1WrnyqAAjGfVpe9OlQ18qIHinQRTavl4zUCsYqYPh7ioyOwa37iKqJxUTkoxDo9b3v
c6zjGRPw1YTUaux8jinQmkoIYnVBRy1S2TPipxjektgcmqzCG5MNEvIgVb7aiDchRBY5Cbko3weq
wStiI9OprjXESCPqIjPXGrIXmt/9LPYw6dGz22be4ZnVilb2hXl8qWHBznIypMd/+LGTlZ1+mqQQ
k3Uw8noybAIr0NWraCFMDUtyRgaEvGpF54wkNCiMclhZBfsBOp/Ydh7nwWDWQuftlWyUjV0zWgXz
AuSgcTE7t7J5JnKQUKxG/RlCBr8HT0yQJ4c4mmSF30nYFFvDxi+47/LI/FvzhsDA4r1cLQgJyUGF
QSjanl1v1/Dys8/NnZoI+34PZLYjvxeoQW0xJ/DDWGOd/d5NZaI/5k2RnvbdtoEWOoGtYQQy44DW
egbbUe/HAyUIZbBiPUHe1bm6cXuNFFwQXkzKRsEnG7lLM9aHnA7lIB6veHJwF4Q140o+Ywr34FLI
rnaUzIrZuGgouw0hLO970twONA81HAlr9fu+RAD82TbVP+IozNrQLxSDJzZVKDgo/L2yBL/ERiVF
7vfmKYw2CT7G7dD0AgjDsuNc2oG2UOQSw1Oj9KrKlGIHhNmQQLQ4LtT/u+Pbe8266zoByjBCQAZt
xVTk7fTnrwvlpH0JhlIKsoh6KyLkuxxaMfHvc05dK8Fs5+5Y53rwqiOhkk2bxSDSGiBJ1VwgKTlV
Gjm6Hx5qyLhO1TUd/yYJRyEbOW3qRB1cj9OrTqqKJvg3RvEOsAOsUUsEzocg2+/nxPfEzQ5Nfoaf
JxF93kYRCL6RmKrkhhjbrZJK2jd5ISuQUUmCv5YKEUW+2Pw2yIq4tTSvWAycLA9Vt4UV335Z9LAP
F6cUFx/HQ2aD1RaVh1SHvQShzb2PblTlta4Jt5GmQ1NzOT7cHK9rw8zw2x4W6KFR5YIh2NTgrJkW
habeUacgLeTbk+YeO7BE2G2iKjhz51IqKXcjokd2rUFebUk1svVEFK6trKQQfc3evbM3Dl+fFMsW
+xSI9NuTQdaUxkQJSytzUFGvl9KAfzBNupdl+7kv+5H8D3AZGJqr8nqWMBUubi/P9dpXMvYvMVHQ
+uv61PPh3KFiW+fyoAjKF3Xz4itpl5dNe1mMWsaXeIylM+URvGIbmIeVAvEqdZI4Bdiuxcmc1/9Z
Ruv+TyGUF0AHObHJXRw70mQF5kbpvSeU8eD+GPWzsn8pTIPRoY+TNqMBOdNRziiQJcEKKUuA/N47
aPONbdRURfJ2JgXhkkCBeBHtpxdZd8cL608tHqv2/Cj86wCgsCk1RqCXUM4QHzwe/b5lAryjtOxJ
VqatCEWwUKbiWx9VlQSyUQ32VcgH6Utuvh6PPPqcFpE84/CVc05Fm5Osvc5eOiRwSU0d/JUfARBc
hg97prgEuq9kx6U9/yZBhVPeDqJLMJqG4+RO0otxZmuRwTm9rcEV60p4JgEXT6kX684mJvNMekdt
wcFDVwpCt91dbqahewgHC2rliCiM4cEgX1rZQWadyICakBI7D410LDtmmtLPP3qXD2hHAilUI3vN
J5S/lMPaDGx0jsCKa8HLdf/peezvOoLsNOajiuT4tsq8WPyIQs/bsvXds7eR/+cMqs70aMh/hYc7
yrN4zuV93oXusSCypkZOCHqi4Tl5tD+mHl7IkCFf+518G41beQJG3o8lAHh/bruuYAziO+4+Ojgw
3bFLxQTMqDWRUzlm6L5OF/4BFhXIFwRIL8UUmdfNxfNA17aY5fTxModJG/nfFGERJzr/brS6IKbD
gqWOz0+fZr/rnIkoV4KT9EX7Q03LVeUF3vAsK4yvjT+AyW7v8WYye5zPne5nqkOmOcDzGhs+SqmR
rvlUq8q7ea+7lL7MTJGozCUThVS5J4DaDF+K55UyebGhXU62r2FogJzMpvDe158bGVvuTqBNUC9B
hYumg+jW1bKbX4Bx+jap5mAAK2vyy29BlkSUi19bx+/DQKRXAYMnSixsm76oUClqD55+kLd4/xOr
pH5OsxeAkTe3dNJm3TAcszVPiorT/+1BWkfnPURZDbQlc0jKwCBQcKNTQEU4cHzHX29z8FL5xP+W
ZOGLw3DOvO6hhSeD7FTm9jXxrDqbQ7UrLFJUO2zenqdszvWbkpYJdOE9IBx9MXlNe7FtB/FLwCji
1sTM6EtkHK63rh+6syQSGglFXlr7AmqaDFGwW8ntvZVDUjaFx5V10SpwlKxliLVR7XzY5NgNA7q6
HCaa1eG9ob4Gcbs5LNlcxNeT3+5fuencbTEDPN1fbHHCylXuV0ZlXrYqH2rc8fpYU/hhpdhkRaxJ
rVtkc0511LOC6EfiMH33p+HWUOcRYPrB0DEFEmrdGYPdIBVOjvwx1FWndrt4S8E9+uPseUOxiDK6
JTtH3rV9ErBEjvYf/ezCbhxBn36l12nax3YlB4oZ4NDsb3WVAvOhjDlZ6zmrK7kx7vT7xVLGuFMu
/TeLnLMQJO0KCDSvwNAsr+ypWDrHvP9kEtBgHLHhgiTye2roR7yJc5pINf5FIpQKO9y/FQyBTP6X
viK6K2C6nlVkZBCFGBIyuWQfT7YPUi6nyZQQKcCvsokHDMemF7XmzbUqi605Z08qJjW/XaxVKOiZ
ImzG+doyQiWojc4Dwc3TEM2m5lkHxB9rRSOiq/BuwdW69omYczY5lSJzQNt+PPugdDutFIQJgwyI
udSZ8LXr6URvzL6JANJKzowFZdth+S3WderXH92I03Co/lJdD6HipKDWFrUMOZ+eVl3Od0/6KrRd
uRIj6HRvM9V6vjY+i+xeFQXUH7sGisx0ciZCB+1KqJykZJk+bigvhPw9UfGcd3B38/iyRJeAC81I
xrFR/TWDorxHcisWH0c3egXHJb3YJBGLnnb9shp/3qlUfndp2Txx6tMXPKBgQxHi1Tmlv4tDZS6/
G2BMrBLH9+89McJdz/t3az0fb+EtxpKuMy5xFDpTMoG4KoBQCgznSVCRX63WuKFFvs4JyfgddwuA
zYgfeoJ82S+/iMuAc9RAm7NhHpT0LeEAnBtM12DyPWIZFfg54kO9uovKDc/NGhULhZJbpCa795h4
JUNCi7GdHb77njA2NAXarOnrwSZjQzt5LGE+Qe9bDkGKFn8a7fiCzc4Ka9WxugLcyiZvBjZaeLeH
AFaOnS0FzAwLpnyslHbbOloTswy+VkME2WlBj3ylDosaNwuYgh4ikgCRHSzBL/Qwszb9XoQULLW9
52BWNsytko5+rH3R26Qt+RYHF/VUE3pP1DMZ/+wm0+Eha2mE2Jg9AezBu/xbQSLfNBmkxQ0JY2NO
Ygkop2+jepyDsyzYXBPe8CjgcsbqQ9ErBu2cIEAq2Xcva7q+KErtgWI0DudPe7/HRwXbPDQFWOEd
pI+/qKVcoWclzIVOtF3NWKLzXkDGmh4SKQHOL18uXdnG3AGFdg67x0NYiTvMgH4S2bFFRnTFVupI
4QU2L/Py4wMY3+McSdGBeZTkxFQ2VlBw/uGWjjvcTfTa1h1A31qxcyyf7lKh/rcKsLQM6iBFQsW3
2LJ+Dk+qa7zCx6cGWiynTyj2+Rty7fXHaxBeeAa7s957lGxG2zrOPeMw6ZfMLDWZgLKzjz4pT74X
BDziaUh2dBRW4HZsJtXSEiQvSegxhfziWtYlQ408BdBApeGpz+PWUJ43UXdUMLRcBBFLSKiUKqGw
ackWwOgJuDjFoUDKTwb1tYpr7ftJdZ+1KPklPg4Oqkx3BFuejqYyXm5gUQjnL0RqRwnhB2/7GqoM
Qha5Ey50Xtg8YHx9u55o5TjlP49uzY4eLdMal5uMmOWzZIVK2cAQLqFhY6bdLTHTTO6b5sKQPjjk
bhHUEI9L9HOWBk/PQ9TLNH+q97xpZE8FIzShR6sTqL5neCBVPL+LayxgldJZCOmHG+moMSr1jpxE
EvGhBGHheCbl4kwXVzIZAFK0CiSLkv3DU94uD055kSpdQ5t8cMqTFKWwVBGoTVTmrdnUDXXnbwqQ
uzvISqwlYrnSGjhombC36qm5Tvb52T6cTMZhn3VrgwYnuvClsfrp9Mda66EruX/cuCEbgatu6oUw
CRTZLtJy02l2hlFKFx3jSBNLAUzkhjPj/U12xRL+/xznEGBNnejPyPH1jOrxmvgBp3mkLkmq9M22
3v/bsHkaKaXKmXm0hzWF+3m4X0czCLHveT/xpAzu08wL3wd7L9aEbXQrYMRLJNMgEdL3s6JQlpBo
3XnUW9x8t90Xoikdn+dGS+8H0B79b26IZqUW9on32sHKvdBCf7mgmCQOx94fxZYFp1B+FzF0mEv2
+IwmW6Y5gvcaHRsg4g2WBc5zbf+w8ZhDELMYNH367IXWi2Wpfq1a3z/W//wtQl6H9YHxhVX6Wrll
+29qDaa0rTjwEL62ztGsFAQdLoBPEGUOu4G5eko7QUPKTSgQUR0yuOIhjRld3UbLFA31dJFemD4/
S73Ge2F6JPT47Rm39817aIPmTO7hYmaeRazBeg6AqALFDnihchHxuDvHnv32oi90cn7a3bJIGwcW
0mjc7UF1pjLkRjS9IYDgjf9nLhvGR2/XPGoE4u20P7nsv8XEMxylD/hVuSyspTIUdQaC50HHoEq5
DWkMwgb+gvaYHiqDywsgiwh3rVzOx0MA2sErQgo4ulcjQnbU11WT9CT4u0Z6SW3EHQuSHnDCMwmO
pfK6hIwvq6Kr6+E5zzfZcwcB337XEp22Va8l+3bI+mexflOSqODkPNuwooGNX0LiUsJY7G/Rg7/J
iUav3fTviyysZV+Qor5+/dANc/rE8MkmrxxRlts3pdYA4oIGjomeyROt+l6RGATPZA2zDrsgjrWB
dmRBeGHTMt7dcMkl+VKpgNR+YSIn+IvRr7W9MR4EV/Pm0bMzipNq7WNVBub0XeVF+yAypc4SGa/I
sA2oBbMi3sf2zuP5gicRuVUyxN0rttY+QX2yRCbLmUVSI6L7TEaaPcdHlCU7aUe7P0SVrlQHvy12
xNqgGp4avFYXLtnA5KhlhlKjA9ZQfyHi7FDgv0I8SXCBhxcBp9KtlWR/MI3/c7a7ydQkQzKk2wbU
0DidNCQmROEkB2pmXIQBsEqeXnDfRV6lxzGfRfkIxStVEgUf9k//BlmRCTcx7xB82/GkRaAwd1I0
GCdgjbQuSToMG3XSP/RbL/idJiXOQYbvKYfwIZeBvIbi3GVHNBMoLAQZLIn4ZwfTeA+wT4U63Jvr
piF4ytfZpafQXspmLPys37R8jYYYMbxiI4wxVG6cz1FY2RPSeSOeXcL4vQYKp88BVi6u+zRM8/X7
NM002Ei3ZY61jg7Kvk4sNM7Zg5UrLdzyA8ahAL7Ig0nknQ4xPEMpUSpI/YjUiqHEaWYOra4nqjAE
8213GKmx1VEi0JPjYHyAdeO2cBYosSXfR3Gih3oVKpD7L0jKzr4JB0it51k4zHkXuh3Ur3ZaDJeW
rZfkdunZIB8UyVmLomj/o2Ms1a3yAyFvyuhWa3NX60y5TwRH0I+tWy6xUQ6ScTTlwr3LU9m05IsQ
h6DJS3Aa4LnEtzndtwwnzDl1kmjw5rXedwRaQ4/ioS5NsS8o/eKHl9feuLcDtvW04Sd22XAdByqa
nvsPyLkisBNWzkzt3+IKr+LXRGrlJuFsbZYVfbP4YChhNlOktoQVWe1quRGNnapj1ZoLFUegEpyX
3BNa0H380Q0ml/W1EMrbAB1lagODNRWBysgTG9KEha8q5rJf8dIPIuhaU2o133uZz/yywfYxAVwn
Q0mdDeAzgmtSZEBpNmtN46kY/bjL7+VSrp3FK+SzZTCYdcUritW2vMs1C9DRaofLL4V2wdEfMUOP
rxr40OFr8K3C2ORvsdoWOFiccw4V8FpZKEWswc7ObckMMfXFgTLtDYVpUz/XYAeppYlAFjkCCCIE
CIC5ol0bW/o+Ldx1NJjYC8x0dEaFc5HVs+fQu6yB+aAfY3RJHuOW9tHSNpSX4VGVrvYjl9GY21CC
mjdnsD0yzlRG1mWka3anUu4WoP0XJeaBDlERWTbNZXQsQ2QsOboYjonsb3A82s27DLxba/3soEOa
mP4bHDbkNqVj43GeFlk4IrqDqyXUHgwXVFoXhuGe0EYCZx6Ao4Vpi0aSJjBVZohP4ifLFiXONr4x
mna9sEp0OpxsX+eop51LmoEevvULqDUBnNEcfr8N57trJ3B7kuhiwITI1Cr4sgWccOQeguR0F01N
jYutdUzETH+Se+5OoGaGc+2hICTbbjpm4ieLVJZpISSFK/3jJTdwyEd3Etxa9kBQjWdYgx/TSoUK
jQ6jDQoxOYUwqlTZLc0I/kPAOkmx+gfMlXd1Dln5CqhBV+P4knSFXawFJ3Q+Xl29epLOcLvsFMuI
2BLbgVTp/IkDA7lPnKUwS6X6Y+1RZQsIvvty/cjFTrKPvSIb0WSeexg5N+rWHLH/LEgMVzfWK9EY
JfBSk1bbYefmlbRewAyTrJG8BzHBaFS8EP7ffTdztxbhhXZSTsEmPOUs7y1kRMh7fjqeQGmzWrpq
7DIpmwF6jKLLGS6W+8+GJuzjsXBlFCRmJAhdqqUkpf9nqRKJEEKDBTEjBf/dBs/nx5hdTi1d+FFI
zIQsQB5xWJlS69SG0ye5MohxaErnlzjdqLWY6WGS8KXaqppZXkQ9FghF66rb2J0rDwQlJzq0HY5T
70gJsNGfA55UNGB2C9/X+cLOoMOide3cVh4pykMyWEFxCe5y3GsWn8e4/lMY3tRGlyTu2OWCsICS
4z0X4NIa0IWytH3lMgLju5fvA/DRqqxgURsY8L+Wfay6+45P3c3mXXKDPfnhpD8BrKeMu7XpWkhi
6ChFYo+4Bwxd4u7GvrtTH/edb9qBrcQafWxcqPyKTFDbPvKr4SZRaLDa5T07oubwweMEzlUddHGV
q1f6cKqUzvkdi4e9MiaKMWG4xZYC6PJoCqdHGBSQnI32uMKH6wttawpPul/nV/YkOdpS6oFzNVlC
UxfCl9kecMLaVREVRQpgTZK1o8k5CY+yGYVdbKhuwiiOS4SWjRmKskF9KrDn+RY0qZ6coniHY5/6
OwheWvc1+9vmPCxab0qyu7AnV6ep3XgI8OxLVVa0QoECEffpDez9qlQnvj3IUuOeI7n0pIBeZ0Qn
fUxxooD7nB5G09TLjFpNhNRhxl8ULqQsCIHpEv7gXHb89dIySvoB3CjYKcPIW37AzMiXuRaEZf6F
B3OUHYY1rdwgW1BEQwlzId7hm7kqLcLcYe47ANVSDuV/a2SsdpS8dp03So611bVNIOjDFikPfFdg
+Q7/BXMbZfPmqd4jVaYTucZ1vTtxlto+uqd+BTsCGimp8AXlpSDHPSDNJXaiaYQKHMHet3gjqfQu
8GNn2xzem9FNEy0u8x4LHTdkKA+O1uBHdQx1EoJCH+jjT178D2jToMuxh5lC077MA6N3DfxzV2dQ
iQ+Ap8LYTkldEyWHtXvFh1FLTm8DHjaa7Dk=
`protect end_protected

