

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
e5HXux03McEJscFg80ZeuZznrIJptNO1SFQrz1pWkRP7P3QoqpS2mJZRj5k487CXMg1LSvaDqmT2
OL7PFCCTiQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
hgCd2yd1Ey3kW4Xi8EYui71ziVJlfu+yPA/iSZYYtw01d1xCQQbb29qdxk14t+CL2ulbT/AG/Tph
KVRTNfPiGK79TWiKACghNYtvZsEbOSiWp2tzfhZzsTJKt6Q/Tnk5KS0q9lShCg5S46ZxNmKbnoII
YTwtWH6VQAWKrWw0gQI=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
tPm67AAwZoJgqE6aGdH3UBgFSYY0hEjWFTT4t/9DwITm8ODgcytWQbTKxugKHOWkwgxnsfouuhwt
QO5L1ilTy6LqSek7CTlbPwPy4k6tJZltW8YhAKZe6X8IJvIcPyG5jVx+6vlxM+WibCk/roITcPkm
9mxr1ZYPG61/YergLsZha0lMNqW4wq3ID24jQg1utjPuifsU4f5hPPbAaCmkiuYhwkMNuj6VHmIU
m/hi3cIAvUetwb+LazrLlZHRjTpygeOmt1PlMgoOOBXow6h7AJvjUUWQmikWL+0eXLxGX1SKnX5+
Op5qf6RZYmh6jR7nN97PHzmxB7CCeLZXWlS7Bw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
as6iakL3FcmLsNV7kgkV+92olQIBIL1+cbziWnl5Jjo3DH55nMZNZI73AcIS3DfwFYnxJCqB2SLa
SuhR2kAcUXkLjAVN6C44hN7PokTEYbZ0O/DrWDwmWxnool0q47JMJkAhu6l9w278iR2KPAv+EoYt
+JQKH1y1F/+RNrZ1eYU=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
BFKuZqEfqjecGcxpRGmpCDvmWO5m86XHlx1Avi4sYpYvtXIvQdg65YGdV1jpIV3rjwKZHTLGWY/h
WohbbV2nhc+5Ruu6dAeqtH04PeCXz8zphv8vhckLjpwnJT0GWHiaXAcncvq/6wuXR25ASAvhi3Ai
lvDf+vNs8eunn+yE9uSpqndZXDEQrdOREqbbPaHrHScG2A0wHmKCr+QTb2IHKcEfLgWtjt/VCXIv
5krerkdmS143EXlDVZB7mfDSlR6bwswWViVYnH2kDpeepoBCAgyzi+PoFfcxhkn8DGVtdsW89QDd
rLaMLCCjYMVnBfrYxBWw0Bz0mfZcivLyxd+wbg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 18544)
`protect data_block
MdChJ03BwLEMVY6/i23GaFpH+Vq5prhGnGCGAm+Rly01rJV9Fh4Z/RRfmjhZfcI6t5vpc8dMWX8o
JC/aZRXQrRan7QbSBfgc+l+m8Nc2efogJw3NoZ+oNUpr4AkED8G+b7GXB3XrHYonb6WquKJS6h6z
oTfLnNB60EUH9FaCrdQqyjpgjHlkoIr1q/oWAM+btwPxY3bCu5o/mpn2wvgrb4jhbBlDzWhxC/Ln
Ic83ES8FnzJwSbKXubN5KM5ceiDlUT2WCC5td4FToTcP7HUdb7CJ/AX51hkDRGcU4rE9k0IRmipL
UqVov2l5Ip/XGDEKoIEnnLM+oKQwUofp836nhe/S98Yk8ucEkmhVPjm4klQFotoofV30OQzB/9+N
TG0rPT7W8C1SD4ZhRMaLSfmnkRKbcfwXwYDgSN/+QvDhqo4WG5jyj6djK1hf7zUBksvXiO7hhbTb
AECav2yGAuAHOkBndja8tEWppxLC6WCrs7cPctEiTPKm3t+Hvobv5rBDv2nWSbc62ZKJ4fRF0Jfp
2Pv3IrjhN1wxYO6tP+614799tQ7pA3ZbWyjh21TFqOome1LI59lc99EomxV932h1tm9boQmtfwYi
cAOUH1dQqF2BOrepm8HAcu4GbWPoLxFnB6R4d1g8/u/IvPetMnQTygfTsmikg+y4r4RL/4Ohkthj
SPelEYS+MwYfzQojwB4yN4kMVpC8LCP4MDjuowr/1c97/vOjJJ264til0k80vOwcUYoZWhqgIjZJ
w7+j6y/XiSLB1QI+k3XazjYbBGhy1Xcgtiz/dNYOUMxlu7m9WDKOn8wO4BqiB19DjJZ1jdb2647b
CcyLBghxBCOZidR98Bua+JiNarKXEudO05dQqDp9Uxk3Cepu90w/uvw0O//XzkdELf5TeWBTkL6N
/ucUCi+y+oxcvto9UhQY9ih8NViHCdsnmnjUeV9u5hAedPc+HJWhiDqKb/Xq3YrcRqCvTu2BT3l/
1SQ3RpzejyR3NjBHxzNR+NNwph4JSP4IKm1hL6asOO27TRKy7UvzrXlJcmgOYp94RHGihEg8dQVE
3ljVTlZ/UJckmABXwqOZM9SdYmLwItJO+R6wagnSQLNvpgjlPic1aOPp1GpQ/HnQK/ANGsMgjg0C
1mSpjy8WOMER6M0b6ayh2li9zZ4BsMDUL08Io82cBgrLEikxP6zFeQ7QTaztI3u74qtj3FMG8NI1
3W1RV34i3Kn/xkS8YcNJknLPpFvAhe9mu7YkPg8L5miCc3MCZx6JqVKJQ4+6bIsPs6IMgVaEQHK4
6R53gcLnlFjBR15W7VqMvDDq/SWbSuPu435synn1t5xq34fGCeJ4kJ0zQRm/q00OHWqMFJYRQ6+O
Bw3QQkM1u/xENcRdh2iqaoWlQ6mMya73nCLRPw3pbz0GFERJrsvuvQNT0H1E7hHMvgYd+dh0qAQq
L0klE3fN/qAD3a9hbxy/Vo5K9LKCTu4JUYbR46+8/rdF2sk72ZXH3z9b6ds3fpEyKhtDKzhvlpPE
1kT/TOxb1TMMERvFdyCGY2RS5/gsHWVeiarMOuERBRZqkj5MR5F8cg+q26vECzZE+hbQhBr7Z7Mk
gfFEPsbHblLo+AR++q7/fmScyjjn9fQZ8/mzzmrNG93L6fpqHk1FQFJYla9CtRnqbmOJp03RmrTt
Pv6CI/2UV7tzPSS3kvQbUBb9tvSWzZSyWJ840ClkdzkBNlLVKtJfS5hHf/u3dAZoccxAK20ZG+m9
UMKJqliWLpCqhTvDmsnep/wdTzuK47xI6BrJ8S67jAGq82g2vk6f3IeZaslXDPW/NMDekY1imepP
i/vvPYwAxOATd5wrPRL56jm3r8HFM9TsTDwPd3CgPHx7zeh5YjaXNofz7r4KPJ3NHcyYodZxap/M
6iAHoxYnOtm51EJb6k0JFZOpYDp8I7BUb3KtJUglcwDiMqhX/Gw1ApHmb09nK1C/35yQit0/7NNO
tpDjgmyjnVBBukkjmZ9bykzq2t/q/6/wf0P5rxfoVa/8gJve1xhOMZ/mvhi1CmFL8gUCu3Uf3j94
jcayeZyuXpWg6/qnUpC8Xqh3pFZWN4EbElAR5V7TrEs+ziSPXh7YdghJfElNL9+1f+GSJCO8enrp
d7UBx9WvNqd2oDtllp97bhB6F7z7q6okUK0zizVneIoHN++FST2yv4Uivssb/JNqXxdNos09TNmr
O1Lp9LZc+9RpfckH1wtKvA23iGtvunPkSKK00gEauKOIqB9mlt6UbepTBhw3/X4BAvTgrG3nVxVK
L4xXfDY8DmrXYvw1Xwe4mVz5glXdewaLg5v5L+ym59oAmDHKF9sgxA7zHjbGCcNdzZ7s+gAnQ/G8
8N9FoPFulENAbxF94e7knvrOne9MTrNwdtP2TbKEQv69rNMMVpCX28KYCFRKFMaAAAT5/zqKZRqf
glCM6uUIr96FIbI2uA5nn4AlklxmfZdXs5DUoq797wGDYmPUxSdnsH9qz1Xogswv3FSwMq/v1cHr
aKGj8x1kYKv6igU/hQ3wHWguwTubZ2a5+DqZM72YioXF8wmE69TFZIdd6D/RfZ2a/sapWR7TFpgd
T17I9kgPUOR5IR2PM8fGWKfugiqnVKiYCYzUfrof5oXK+v1IdJo1o4CICc1F8Qqk60Wa0mgEqztG
RknmvC30KVGKX7SHJkuGIVho6S4OhOiDiYTyOvUWMBpW8aRdKv4zZxkeMNYqlq2HDL/MJiFVBdS4
dkckeYkPvoWsVcElNeE5gyutoCvLEBx36glIccTzv4c9CI5qaKT+5pAskOYXNh9WqnFUxCQkIFqR
6IMBei6EbNGcEmr/SeVwRKd1KFMJlrwYh4+fEECmiqBzemC3BRY21gAXMariES7ajeYMrfNVfnQJ
x3Yq7j/VxPszHFGaMbTG9CPi11U/kZQ8yBfKcXqpByu1KZ7KripSsQTyuPXm1LJ8FDUcM1eBKTLs
OQxZoMhlkFjmqv2K3o4ttWUOHyYUm8aIgXdSHW6PjTK8UUcXmtis50tRnQAbUDjV8ijsr6FqSMgm
6ew58wrNhPOZI7t68ktYNg3HMP94ae6vgvswT993OKqCvg709/wiSQ3pkcAF/z5LnzCC2A4C92dU
jj/TjltOEAPY1sXHgGc67IEkU0UTxi3e08hn2WuitA/odTVH2Z9+/vTCJ8widWRpUHOR5td6nQUn
kUwEpSuLpY8lfjJEf5JP6yNTNlolKnolZuRcR1LbATed8iF5AIXuP2eIG73yJ5ON2CdDjsuwhVrU
FhSN4nzeQIqF6IYR4Rhv5m82oAxr1L/PX9L93UY8vhodgPneZQoeqAPMc9kPWMip7Do+nMONGf8n
T5OqxxSwWUkuM+YgqV/pjTHtDWA4BWX+5QABmCTP548zxCs9uBE/sSHsseYlO3Yd11rQBWavAayE
CMEf/Q/pXQ06RrPN4PrqTJfNnjaO6v/O6GadhLwcJ5ImMugGjRAnLPrICz+CBiXhtxg7teIl3Wpr
n7HVnh/xucKyBqy4vdGNoAeMsy9/3eisi+05WolMI5NGz+3oIw8eIsDRPxGp8gckhaoGaNvsJwCT
ut3XuvkZlQk5VRyeoZb9ChLNJze9873fJ7NiHN8NpT31a9FFaXk+BT0nncZaSAcWx2MF//M7kQXa
+yoXWxoHdpm5yMoHViRx8c7a2ugQOD/j1s4ePQRboaDJr8IdrzMBXBY9/5AW+J5P9/R73DhuvAA2
u14wILDq/mtijbANDjD26wis55Goo1y3p6l1AJQOKg2EUScKX0PL1eyQKtfK+t7XDK/MvlOHooBK
HAgPTSbd4ieOI4fpWS1hFM23MTcvwJml8+iHYTor00O4/4wLHQ3ieBc9g/iNDKVXuH2v+JEJjDvH
hV4R0KPQIihzn+rj8Xg46WGZjafQCmG0kdKPtxi+lZnhI7s7XhDqisqHVxLlKs0uM1JsP2g/SZ83
YsQirbipvCA0JcR1cL4Axvk95r70QeUBXqm59zmeVYiatZLMIorj0gIDU7//zWBDA5RZUzo3vG/O
GB7+qhZsrvNxfIgcNTWYNTSCEsw9+efs6WAdrd6qWZQwsgtWd6iphi1cuACKkd2ecEK03fTV/7ha
7YTTKQ3PKq/thTfDjnqjuw6SRIS+X8DB8G+pNvEDWd306ofpDR/hEPO7Zx8YHexnf+gnLh6SZDgb
47iKRNGb12vrZRdsMU1gftv2+nEyhxcyA8/Z/CPjxjYlVQTiOETy4qV7GWCJQjBO7eXuvoqbGpC+
fskBZNuTpX9cypLMinvuTaXej8nJmucSh1vi5r0EZt/n2jRTboM34rCEaFpT0583KOYnBOHwYaf2
7Wgcb3p0ZESKgCTxJnFrB4mBRd7DbBg5kSPKVNRZLkZdNF8zwaiKsK6TEn2XBdnoZQ6m9mWecEEu
vou7QLJMwdWa/w1rlNBNGHCT4UglgKMnpjfXz6z5f/+6X3IQLEJEq42QgZscjjv4LXIaFf2gXl4y
17/D7jzPQd8kZSoWhLolQlBQs12zGRazoV9O1UABF0X7FKw3cnXNzGRtVqRZMaiAQFzpH0jyV/Ze
/TZJ9j+g+2rFjLMpx6JFGEALMpJNalqsJkYf8MxEab/CFrC/Vr+MbSFNCdAqLHTcPVDetwGIf05E
JKxkE42OBC8DC0MEVztyDiO1QBtRUBSEHkq3XfruqrqqO19xTjso1K1XnLc0SYQiDPypgOhMEiVB
L+abLQs89qNw5hQigMLSMG3vw3FOSCqdAa+OfZc/uL5JNu8Fp4+sNEUnBoq9msFdH+gFrRDE2c18
lbTN5Q475VQcOUqHV+TeP+lB3uEALRNZdPvdj+jZ7yz2XhTqYrOPW9N8acugRTVZ1CFEzUa5hZrd
zbOQYOWNBkMoXw9IGvSAAJ/XTuyE4orgdNcXUvauaiFsueAI3Kgbl53kZOscVLpYID58K46e5UO7
xJEtd/SSSNLwCoPluRZuN4fb1Io9lFE0OtOYgXrkz1FV/AK3XeFGLLw8/fVLCZ829tZk3IBSDSAG
TFEwyKkY5fwr4wSS4mGFS9DGIAnRwgry9SAfoj44HEY1wFl4ePREtKTrzZ3cUHK5vmTgyKMHOTOH
7CQddlCWZkhBl6+mROOvPSN6W7+HbgqM3NhDOJYw/Y/37mJ6n1ZMhzvrpcJ3cOD5q8R+Xycq7Cku
jKipgH61y1GhMuuzmz0j2kxElleayRI5vHhq7uTI7B+6jvlzmQhRirqnoTV2rmWoXxaO/VJEHCjn
YVNdGXFaXlcfFcrJodpi/1rigLj4WljW5bYRcr/x8YLuLqL8//AHAUQMKCoMOSbf1ZE+zA+E0RRl
LXJ71bGVyiHVlMfTaNgvTPfr+4N5sjpT8YSe3pT7PReirAmbEq/3lPXfJaIakDXZGVPlrIJU9Wfy
qaLysdneS0m4kmtzF0WZbpEv+pG2lq39b8K7CJq63DgQFz5qJaH2k/W1HdS6xRy0YHttjQIn6GAg
BgjzmeQGUBSzmWXwSNCXzfB5OIlJsShdKwux4O7mw7saNjup35QkOEQc+MPJqV9OhgVpO7YF0aTV
dco9wi4IJzTb9Oh0jUg58PuM3GSwJ85o67MlYJvA/K2bvE7wV6rQKyY0asRBhNpbA1KKQSyqbw81
3UVHeN9HGhP9xC6BgWJTIGiGCu7WJx7VMrUPald0E/gy1ALhFs7P7PIKDjAeFQgkg15eb/KEfaKp
/BWTmZpQDRVnQiGEVt+Jg7KcKkzm/q73aC7kKxeHd2GcE0WORnTWcUbPOFEaeSjGc/Af5Vb6Edi7
rNj6V0n5zCQaKqJPgF73/PmsGs7qR6sHF8BLL9JBAxnfqxfW1rTMnB6NAPp6ipNoaU64xjv+4ojh
SO9HJYxnc7EJCd+ONlJ+vX37bN+0jKXZcgfCZu3XpJ/b8NwYQwsh3o4eTlih2gal4xNUDuO2INTE
QYbjHZD9Hog9DwW3Ou3ic+dJSZuFuHiZM4WJezh+IfD6SIBo6Jq1Gkr1JiJXwQxiCxGgZNru6kEu
C0lZWLw6I6Y6kPpxlnvJqOCenY5H6IFddFMY3zAEB3CepDezxQfBQWTHxN0RuFb54AF3F9LasFyP
o+6ZFkE6zo8UNzGLhQN5o8Yl7bFzWnY/F5Xwtpl+GB05dfWbA4gZjQHaV+3iuoKml9IeuEJojXMt
MH4djQtRsLfGyFDET8JtkeaiOmow8RYTRBoEKzGl1XiBMzRls0QTcCcJI0Mbf9O4sFA/EG7Rnp+C
BnlvAVtB4ezT1gL5UHM/20cSz8YA3e1uKbwBG+8isjBjgMljTOYgnvhPMxXZNuJ42qnMeLZFFV2/
JK3Kky7Chvkvh4xgM/RwHMU6f+B7+AexpgXChy5xJwCIKFnXtxAz3+7gnME5bZzVvWxxZkw+a39o
iUwZfgjIKDmtL5jpVoTYMxifAI5gQ2lc0mKeHXyFO9hDHCMAbsSnRx00Iwv61ug8fBC+rxOQfXFY
iMsTic03Ewp8aMZ+4jHl8rkeWATMEjtVdNyDsuw89S3VhA05V6BHFcQ7uGwz2Cw/DLaTRukaMkP6
MlPpuYYMBDelEGJ6TtBE7akaaOIMJVu1DD4j6sYU7T3RhMm4g7HIejIap6FIbpJj1AHaWgqQzD62
w2MzuG2YptRyOxN058S7VJk7iFmO0TIHZ6nhGRznN8UZpQKjtokNQCFhWHxtPjeGSalVMbwaTiLn
H9u/pHs0bK0eDFJX6R2Y5dxNi12PpY7RZvr+hgOUCu0bBXDsMV3ry4++GRqRbFACt0k2MxV7JQ9a
7Rme+qKcORIyleSU6kPfQwqHXzxINy4nJrpZiXYmRMFwHdhjk/LbDpw9i53mG8hUNlSA5c9gL9of
7xIByH5lk3Q9h2X6OxVbefyifY1JTsyqivWWiCNr11ftvTrXqFw8AIymqnLwso6/szvUQ84mEJ2H
OxALthnLNnH7rqA57qafoSFFlQWcQu9tPbpYc+bJfFhtBTElmpoNfaADb/Xtw4lqCHzQZC1HDvdM
Nbnm/im0Fyo1X+P/MWLd9gJ6aWP0yn338HuAgJPBigJsHnKgbPhV3a9SeXSE0tc6iDMmJxr1Iezo
dUd5Plmfdw4CyzC6gQ57PXhF+WQgN2p77f13F04/2xjhInmV0lSD83v31rDasilYq3+E/fyyhXwQ
mH8ENUB6jw/rhvPO+zHXawdvgsYR81nU1EYBR5OvwK3/7jhXdBkEclSV5NvKool1fBZWau0iR5sR
zEoZdSR1FTF0GEnGQY4rXDj+Dv54NJlVdWW8AUY7sW+HjCm/OgfeaF5BUQHK0vbPBf0LJdNm1ZN7
BKrZPxs7brs9EF6+k55wZdNHeXVGwuSObyWoib4mgKIIDMXZQpp3W3OrbkOse+J9k4sPJH/D6oE/
WIXECF/TApfUcDES2nbq4jcqDz+KYzeSQ5/45nupGZcyzfkwOjHJnTF2ITWF9PTOXnNwXTI+C9vz
dy76UfKD1tDQQqvw7CttJbBaBXS3eSw0G3DGohIFCNFGGfO8jQ4Edqs7KYvv9ODOG5kwskE/VmhZ
cjAdYTrLLHba49ot1GM5KisebFOpX3Vo7Q1a2QdSomlu/NHCltVw6Ud8EbEu71gzRuCQdfKyyww3
x/2SbBkWC7Zwa1c9cedwFcLf+ReJ0mDpXIlIlrKs/3q6CBRNZUrfokM7B6TOm5LxSE2IUgJ7MTS3
fyYSXIPrww9MC5l5WxRNKti8Igxb41Gonc4EG5iKf5GNLAHHCkntoc4M9aBeXk9JqQ16oYabqITf
EmhIm/erRg++q8endAEIEeb0HOxFRCXqiDMrMZUgmYdhKFscy2vfWIJkAi7xwCeVPXwGmkbxhR3T
IBwVuzMyfE2x40S7cyrNzS/vugi5q8QDK737IpMNjBQl67dqrIADBU7EWK+jhQ4q67qfGIRZXZM9
S6krw5MbQudYW8aNTY6mmVhQ6tvNZDBjXePftvKAdorkn8FZRXG1OUMcSTdn7Nvw0mQVvybenktE
P5ToAE0e1/jNL/4UHxeGzPfyH/Viw44jzidWdkbUZRB9p2JN0XoKcxUCo/c9zihWqjXVvXd94tbU
0PPV0cLzXbtIM+9icLzgu1uJ5gA/7jtM1QFB1DC+IzNYhqbzZwdMulihE8GNAsz1jqGvkBg6Pbhb
RtBG8+MstFHd2ZBjwOeWKUy9eyxhYrKSl9ExvznOG3/LVwN+nwaeDpFvEuBuucfTobcDglMtWbgp
cdT3euXWyvWbPlON5eCH2yLw6KS3lxH08Ym5UJouOd3JqScIQK2auheKE1Wrcotof7Kyd/X40lU0
nDx1XEYekjKL9T5SGkuLzlLG0WaRcqAuMVu7WLakiuntuGKPl8/EQEkOF9Tx+ym9TUUb+dIrCRML
xhBdcWR+Gx4lkwGWvumzS7IvwOFpnpMjmtXEV1e1eCqGez2+L13yKW2rkokFigT0sFjIqg2AL0o/
khJB7vCfDMOwtfDiwXNqOMxzh2eFAwMLbeUUZ8hj1Su9fsOCjCtI+oVbERS/61TE2HKurzAbg2CG
2QI+Yy73MUpxrvum1561BurD6rmxyyW25tZekvUe8p9745QKuhO3tuYYDBeIoc4Cad7SqP1KEdYr
qJZe9iksCAOkjp5XUn0D3TZxavy2XRPApPMCMuH0JtCXxpU+S3XILFx1mT/KDdFin94nbb0ZgzKa
TJyS2S0+gvW9m0DvvalZFySdAdn3kEVyl48vVBS1RnQwdFQ5JRpwLwUfYKowZY0UD9yzPOqN6Ahd
JiCoQdQ0GVZnWu0r/YJ7aN7pNlg72R/fObWRkFbBHJVgCJAhqsjOhpITxO8tHo5KRXFA/PONEdFd
WMwj9H4QlPu4VC64HOAyhX4V2lBu+Fj6OXVUGdM2wELHrqwizziYFEZB/pihZk2hIa/myLKTaoFP
RWmwcVAlewWkzc6NlKtSiSZ3Rr3Ch3LOKKhMO+BPyWCU+pK+nsP0/g8qpk4CkyRxHpt3+A88AazL
WXgRXnoTtuE7ic31rYY5QkRUShief7Yns5cStY9Geyxgiy4Ar7IvJuiIbB/SEKOkZlKQuuGM6EsC
dCPnW+GqqP1rtcWjLzE6ki2wfooB8g8SebKHu9E54W9ZX3RndHQv/krXoyeNgKcJmDvH1iqliENB
hTQY8yhfbj2AK8rzqQqflxBBCsGriQJGeg52gyNU1QeLTo4Nuw/4XOkjQjPnV9UxQAuD5Bqbtuje
YsV/B3PAhOC48oFFGdp6zIzyinCsfgmxUAzKVMt68GgJ4DbR5bRfhv2HA8gdBQDc89bqFLpJrQG9
sM/OC15rnAZwjhMdt7dM1YfZQ4v+aSKIUyL1gheEfi3gZnDawpLEU6U7XNl+J0RWjjxJ4RX9CO18
dR2h3HKEsCj4ZfUvELqV3/yXD8HwXpcLV1dymWBrhqx96uPmaSnbKp3fNs4JGHqFPEekOJ/FE1Xv
8aXlxH3IpEnmJFVvlORzcqcBddPaHxzCKqYu1tA85UvqpXXeqyFL2tRp3dPh2JalbHIwkvZytAjx
ivhctSq2rHIYMLpYR42EBL5PxOn2NCbUnmBev1/BiFaKEyWXk7Na2UHnqB85v2Aphuas/OSji+kX
OmFroSsMgLgbu9OL/lGnOtWQAVkTCVEVT1F7F27oNXiUC4bHnnGUcMdYTvI+pPmor7bhzjAZ38Ob
daVpqpslrLfi/zaECsbz+m19mSbyd8MDT+PRDmC5k1xfTgqiAXqoopzMjpex++bq9GCvAb+Cxhxw
cy2q1+MmAzy3yc4ONLchMAqL+bxZma2I5m1tJtX25mqVPexIZmOLzbbPTRWZQSRdqEZSIf9OJ4um
4mpik0pJR8DTdyhz6G8nwmSdR+AVpLJ/wJEtCP2bWfMdl6S1D4nrJ4H476tDbsYsZrkj0Z26DpJb
2NkxMl2ZaP+udLQnpnNtPtZF6XNYtI//htT1uJHlCyIMRXFHlyzit0kqdX3NuuzNjJNDBHHZ3gqJ
1/mPyWmtd3rHWBWoHw5ydn9byWuEX/hrox/1Z6Yp52dU4CnpW/1q6vh0ZW41CeUjogIJFhPS46K6
HIov0JXQHMq4aKj9ISGWRWAHz66/7ongOJYJNT21FJ6h7pPpSmGmrYLtJ20VZ2Ss1ZeK7Q5XsB+p
JsLKeil5l3/lNgRbLRB2Uo1T/muAf9RKCnbAQJhOvxOD9pPLLz6e5iiAOC44Yb5OmEQC2yrEKkIB
S0xT0T862MuwDAMTAVlpTQmcGTyhV3wUYLJTkPBwZosSBotoapM5qMyAGNm/cga1ya5EG4pq0/bR
FRg922GaBInf8XcJEyx7/nT8kVTEuWQHOX4SGbh3FP25Om9JCQHzUOOWubd+LkcOScjo2LIWzAU5
fYi77xLfyoxj/+e1rQ8aL0yiQTYrXtDjlUP4/XohyD1vLipzfDwz21Uwlo6bUEkO2PIOdCYH619Q
MgUGOmUZyctt0bkwoVkQdunpHvn7RxQltdoDJK2bRXEUPoOcFfC1EWJjY043Gp+3K6hJ6DGQdgka
R/KohChTd/DksEtJIXkJmBhQaxLAgsG6rohuelahbVRqDI1fUIxavnjMwXY3HIEnsK8+NGiDnh3f
0THllTaxSyWw+9WOBnAIugnpiRGQNTxgPbixBrS1MTVkKvsdRDpb/a4PibhFZBt269rvI1+OGZgU
SpDPqZUIsbRbw4krt9oz4OQbIgBDajTqQIp0i7iy7kqOwTM1WTUvvy3HbhlkN2R/F3l70BsWrGZh
iZF5+Uv+s+ncSZ6MTzKqlI0s8rqHRonlcIttvd7RxvHpY+4JbvOkC4Le2U1LzMoge0nRyWXypt6l
vlQpBElTA9p8rnXgU5MvWt7AsApknwF8kY2NMyVGcYtimYYxLJW9yi7Z/VR03yPrYSLSg4m1pvZA
GjkniE3QZVpHNDcQGo4ElPbnO8kK0z4LSIhRlkrqig0dZ2JbE2wjtjYD1Uxfk8/0d8Ww/HE3U1ym
XogbB11tK6QtiSS63zlUtrw04EX526bOn/wX22jhoR8LkRmXcnbPZ/wRm9/sxYgwGH9/EjIV6Gpp
V1/6PUB7OnJIZvq658isfpaWPLVk7zNK6fRyoqfO07kkd8jitWxPSuSGA2HHe235rrYaQMvwzsD+
/4ghgkWNWPCVlxEW5JDK16JhizzaMOgP1bqBLrc3Ty4k4I694NFFwjdyyvvyB59lfftmYZxXytUp
W/M3BSnR9WzmHSPHaBnBRUnuwDtKvmqde1mdGq14A4o9SL9k7AvK3lXh62+mpI/rHc//t/jrsm6B
SC7XuBEYYEDVMJcp5sPLRC+OcyCDMj/wxg/WDqKfz2p8oLlYhTEP3ZJflAQOU0+CNyebxyJHWAIh
7OCffqAJYBYQWyvF0NkAnoaw9KEZaFIlrgc/oz2BNr3ytnKVrJVJbCFnAedHs0ffRVaOnV+Z8Ru9
ohnuH+cjdsFSWEfRfiIVKFYwgm5CpGKOi5YVPyKkvNc6OjRnPMTwiBx+xUmaRSX6ZsQy3wA6Zw0S
XepEyY01FNC0EOJtWdseRKv1kdf8k1Q5j3CcU/P6svkUz3V7G/7CqHCz4UHUmQoNonILP7U2TW/y
DQkTIVMPqdp5b44k0GI7L9MOEEsa1go0xXcP8Xm8YjQH4ycvgQ8l9KyDQRLoIBIpaGjlIPJtE2sL
Egd1DVizWrj25biEQt0q1QGlNHYsjMsBNNMs5TUHKdmBZYIa0dJVFA/08w2SU0jnF8SoyRJrbhlx
Df8TNnaVBEPkYt+1rle57hf8HoIMwu8N60ipyI+g5dBwgmwiFrAKt0BlOrrX7oBamQlbSJu2K7fz
fOo/es1YMOkzJo77ta3IGCTq9MFpFhpjdsfGSsw+clb4VZVX8FXLFjKilP2XEXbN+0I4E3zPFya9
vftPKwCHlHO839NyKYm1PPaZfQTt6KO/qzhWKkkNs7tD4yaPh6J8w0rqIGcYuRCJU30cVOuKXDvf
RAeynngaslhaLpo8KqVW0abLiu72c+3GIGhTECZ96KIBClK7raYjLA6sotL9XH4zGuryEgpkjYXB
KEopHUtR7CpIE1EO8PFCBhGzNhojt2zcuxqmgXP3whDPkCF7Jje9VwzgCGgk4fZ33ObuKMOL9LUG
/q+aCzTGC4Xz5pGwf0DG1718ZNQiCUocAzFLE2HvHCJUPKQ3dB5VGkBCKO9GGx+eyGsxp04pEO3d
nUQ8r056U0ypJquqvob79FILcUSJ3ErEp5k4wZqwzyZjFUFa1uW5mxsVufIl8bOGHSX7RlcmRk25
hDkI6enYzVO+Lo/amwswRT+U/jAG6DKx9oPV7XAZLjPq0QCk7Q6Rcg1gB00jBtTrJAy5M4BU9Fdj
oo1XNZwWxegwi2A0fJ+pFqV9KufHINzUCWYeXTHfB3bozubVpAj9ai5zlnFY13FcD2cTJoitH9Cs
t2YhWmz6HhlzDPsg+/KuHegay6Kmd1eAV2SLh3udblf9ysZFGkyZpFc+hyMNsEoYbsqTf9gcuAyi
gteed+cOZKitfqE27K8qZ2QTuh/sJrLCeq2fJGHp25VZWe6jNnqRNjGJIZibevuo7EhPXyOLpWXS
gtoXIt4RK8soD6JS8HNxkuDAZOK5YRdtSgKChUpSpRVklxp1zUr6ZuXpgX7vbOTgol+klSk3E+Ts
6t6cVXjYj7aPAeCzSQxj8uhrfcZu4xXAb2VtGcAL1FZly6vvzBVl9Zy4xs5cKAhugBClv2aucicF
AaoFXWpF9tvuKmYu5KSPnJXpirnJlwAkx7NSAL/q5gBxv8+SzpSobGKhF+k3nVXgrc+aVNsM9Fcn
+9EBA5vFwEDhxjJ/RaHXf3Hf4+CdiVuym+kvKkw+bEo1VXiqERiCePB3bNewpGsG+EFh9dgFlfqO
S/zcsnAJp3GO3SbMAU8sRtNBI9+/yNkWWszFDJo6r9+LGmPhmR7RtJUUiYaCsymK7RBGqfvBGE5B
fzQ9R5T8nwS9HREOLtfOYmCkYl2hJ8dLBJUZ8G+RohkD7Vg04Tmh4T31OAJPfp7lmacPR0vvmNJE
3mU5oveCdWn7cclIsCTxXsgkHa6+kOGlvdW59mRRFjVJhuwyuwp0ryYX8N38qGYV10Y5/cXMMce/
qNCIYFYN4t7RM9r/GHKQhAKHdA2mbdCA5MqdAY9YPQroLrZdNaHN8TpYfRVAVrM/y/XKyfyHXst2
ckaAUZ+GWRwEBPO1CF8YIN4kPbXijcs0qeJZx3OcsTjX4/gv1VurOdbZYdgj23Dk9eO9Wa7xXRWb
6pdPhAEIzSdVyYpC3TCRpHYEUH0AWb//apO1ossqYdeMuyi6OKzBA+MicLdi6EaW88M3Yx0ckR6t
eY9jWfF3nhS5P4Vm6Y1v5BHNJOzA6+hybrw0rBPJhsExrcU9X+WXdONnN/yRDMAf57zwu9yA8KhT
5Tnv5hwlumWaazWuU/Nk1VmmwOeCE7kfjFn3S5QWE4CcyJgzv4qzkL5jsfdTfNKLYbw3e39EjXLC
oAN66cggP2XH8IDZkDoAllPkWVt7ycH1zSvTJhH5eZG8CQixDLZtfbOTSpHMqpR94AhLTRD25nMm
fJjhuux2Pob/cnEwtuNm8/OR+SFto1noWPFVwzkOlBqGYsP1MtClZgOwWMC6Wd4Qdnam3Q/k2OPR
S1SCP+tROzUmUcX1f9UgAazQRJBP3BcMJI0v8aVCt94samY35yEe+ESzvTy/nthM+3exXYTK/iXO
vA6p5MLGYdCJ+JGdpNYISrPbS8gcgMDz6F2vM66OCUmP1tvKe9VUok+wHJ6C7ZWemaQOAVr6GeKr
Gy52XuqA0YzHo3WMh1LqNcemiIBS9exnqxtjKgJHfiILoeaHuW5HjMkIK89+JthWGShpjwuR5KWj
afu6MGIXUFOob+OyAS3wTwX6bOHY1cBpxDazux5kMjs0Njt8+3ld96yAn/a6agPA8p3lDmj7jGkE
d4lwkg+lp4D9ceqkZ79QtIFT4o6dypxawODMWaJ6ECg4fls2Ny4VYWWg0c2eO4gJFvbHbYpNHmTg
ty+lBvkgMyUibHPHn24NvJBOxwreUBpzOCGSqdpRboXMIrBzz65/rwIqHn5A08LKlkjkgg5oB8w9
pVLV/sysrGlpR46+zjEeh/d5fbqHjhdBqzRHwFcnxaQt3oGjOOXVz1ZkajmPAWdknhoKyWrkEN5m
F7lXpXKO3zRNedfJsWigIpfVIhXD6B2F1o55wAKVGnmtxULr9al5q2cNa4625It7/ADATpkm/iu8
6tK+QZmgOJ8qwT+o3CaHGel3j6f4Ah/eC6IVhMmWbvqGQQgwDV7dkZ5lJpf8mb13XHrVg7YmUuSb
caP/vgH9k3RZANw78br/fIH6FIhjQLRmsZDQkMoDkY9/h4C3pIQw2TzHA2ajsDLloGh9h2fri+kI
G45nIpUIuJwIuR3mjThvhrkPeEzLSNjUY811Kk4FUmvxgj/aEjqhyPHDbdbQjxecNlnOsMrFwuKz
ZD7Kpi9fS2Gr9RRbIPpK/IktQoHqmZqjBIQvTd69Hlk5ua2JA6TetvRR5ASCWGBL3Ckn3mrPpUib
G1fiqyC2Ku0ieqwCHpv2IPy7dRPw7ykDO61YcgQ2olYzGTk3RTGvUNwi3zpH30d0fD2V5ielu86o
086ABAdKTgxPIMTdMxtgeoWdclM/ipIhDrOvX28I6mECmSnP182qNrz8GNqdz/WsPSiaWy/0hHN4
gztFYwLL1ex0rLDhFuP61jlxto0MSwUvEbtVIlh+CBP32yio1uQv/AuUhmMqFA8DxlHD4Z2vM7MS
yoQIoGdK6PyxXtwGqxNwPPDjaU+AmzoJquton1fYVXocvicz6su64Vc9S8C38dDd4usXtFyQ7dX1
lSCIpQankZJ2CagzA38043vopZTtt08Vz8JmopxTJjLTHoRfrdS2UuCyJuPH71EP88gLuQENimka
fCF7CVmANI6YIDBrVQS3GEobIzsrj/CJ4qk+IBxgtWgGtvGzM3oS8XupzIlotxFZ0M9KWYL7CvOA
31wgi35O0RDMvADc6e9agaLvssYjT3XKa3ISwegSNICF2ndJ2TE4vRXenfnfMvPF/hMLoNOFVV61
UmVGgRhkKGH491E9j4TRbXWqezkO4x9346tAPgGBF85OhEK6PFCgKxaeoHQQq73Z6NrBRNgH8Zud
AHXzNkZ1Bkg3ZZ27gspo057pYWZhPX0bZ+3YzeZc24uCNql1v95oC48lHlJX9vkE/9SeEXDw51cd
iGUSN56MIObO/JXbUbo4XSBrL0F+lVkiv0fp8eqXoOXTjFi6Wj88znlfgsRR1MRnfmv4RhPx3AcX
PLAJ1Rh+iR/A7ppj6ieBXaL5I8oCphI6pfYlShH1umfxbq1+dqAnXHlugI+RrRqXvEksv/rfNOQT
HqUISg36AZAhGEOPyKcs0+6HtrhFLiAHNwEIYuDKOx7yPNzb10/oElJWMPbo4NgI1ALKC5pc54o4
ldqPiKPU1j3O+dnzJQIeoE24+usp0GMrf9hT0TClCy4/Tk0zRzWD7HW5Nn+OVHJcWKggI1e+Iym6
T7vEasR/hJqQ9+Yutia3Iq6Wp1tGiDkrR+dvRJAljLyLkI+VOnIPvz1M4rfv/m1Xf49wlAUxpn9/
W6l67Z8YIQOtc5jnbY61joiywSeZlxQKPgdz0aR+0LPfgvrTJuC9jZhjtdEuAb3iuq0Dodm/8mTX
rPWwFq1uNvm3tLa7QiNAaQqkV49yE7DaRWYP80qqeqRCqKTLYjZzDb0m+qALTUYZ4XPLuImz3cYr
eHpCz1uc7L7ob515v9XO8TmnEDe7taCRub3a3MgC8G5MiZFdLx9Ts67oAgoyELqBglvjHYtTfUlC
4u4wmjJRIQ66/aAZJ3sNZPGMYRDaOmGuE8jJ6GHzOMY0BvsFWfGqFf9NiFKuvHck69+/EX2hxt7X
YupIzLmCsAi7B/Rvh4leB0tKCQiTE2ywkZnjpuFdoUIDcxX9AI30lf8JO2aI9nexb3EaIJa/ClBo
QgJoWFW/BcGVSHVVJelR+7gnHcswGrxXX6c0XYpQspRyOQ0jvVaGYc5XmW+7TotPlj/5XKGQVPSv
6ikoGIam/YPt2GOFO33vZE56vrmBTPnehkpiz30EjhXv7CQx6KvDAy0kDyI/YLqPYuA5fTMo20ko
Gi4XVT9LsQBTRFShAe+rrfYcJkc/FmO+Qac1f7MGZgxAPdMk8oQr/aUIAcNnuZZHW8DPcWhZS/8M
m1qNrtIvFEW2QdNefnsp5/o4EIFiX0y/zViiQ0vcf7ehv+UCcCZHGU+a5GXvejorhoQ1FCHkHKE+
ALbZI26g1FghcHTyckzyjF0dcKLXgVzJ3niUXeiE89ZzJa4a7QbvxmHDNPnwAy/kMEE0gsAwK1IX
3M1Pz0s9Fv+zGhVwXWxyl2+4aQKaJ2EpEwG13DWsvTn98K22Rvunoefie9tMCJn3ymonFKsbDpUE
rQgrEsmcNK1Hycii3Q03mQOcBYO29NkP1oAaWCmJ8klWac9dNDFxWLfNT/6bTMHrPRxL4Xtgs0Xb
Arofp+rPaVF7w5ECDnteCwp1gXuLqHYgWcxoXC7g4vEm4eIWeSvzaav+lLBM9ziQ3y9HYgUHprzA
t6j3zPw6qu84jdaTLoGijzT6T8ELuWITLqCXDzMI++hvG6zeiXIqPExV44COYHyVy/NjKpR4TkPn
CwzvDGnKZ4diuaPGOyJ5/XuKMGkh7JQ37DDOdYA+xmFASkhe2TEBwcCHxg/CepvrmtBV7vBCc6h0
a/nbGoB1bCS5Ednk91r8vi2laSR8mKTcBBKLJcIa2T04jxB2UyMgjqAhdAeMwaoQ1N6jfqPv6n8b
sTjLQYXry8Mk6JUiv0ttEMS0KFZl+HvPHQ6wMfeO22fSPbLYgmLW4GIvshUc/9Om+1Gt4KVoUgLC
7djcbRUwn9H8lz1vRo/0Ldd1naTSiHiu1S98NE5ub9IIEgdBtlSziH58gol41OM+RD2gYoT0RZ9v
rRKm8NWIQBKf5UDtaxxAxTlSQrveqJ+xLmMRKVGCn69WJr/QjeuQeJd7FTKRi1hzxKfHYyW1L8Z1
50kSnXQNpJh6HpBaJDkpYnLP3HdJ2CQBxGp8xqTcpxNnTpcMSFSubkT343SeHqENcky6g4QN0xlJ
67STn3NlehtFlqdygIuxJP/fbaha/662JnfybCCrpDPMZZA96Op13WlLikUEeq7IAZpqKcZxh39C
EC2aHDOIxm/yFJvn4F6E5ej8w1j++D4C4qCg036jmM2/jwapPA9EdgpcWOZ+2lQYJmrVNE+JfOjW
AAbBQ6Nko3yzb8EnJGNEMYnV6HebZYoXwboO2GiRdX2HTlyv1VRL216IRepO+SeLajr0q7YBTLgU
Njk2LI0dU2Sa6kWB+g520vgl39hECMsj34tbZrJcd87qk7q8Ppnd9dQZOlQLkG97STyrmy/VLj0T
J2K2S6Ajhb4ErZd89xS9MqkaV1LFdA/KMI2Yv1WPLdfvyFM6fN6STsXQ3n6FLpZL5M6E53n0TA0F
jkRw5saYKoE8udjbSeeabwcZG8pili7AHZyeUvdgZzdra9PWieCTugf2JGQsyZIsTR+pS70nHog7
FBzJQFUkQFrEuGXHTCJOv7WtnFF/7Kjymx76t+hF8oZDKgl/7QUbM/4dAV/4/wlxB9GxQbClgIk2
CoJWu3OJvP5SsUIcSgPUL8MOipZNdQFe+Hzxl2sP0FK/pvcgSmIdoIF1xWw35I59kg0V7LjKQ7dv
IYrIA7NhNJ+/xKwIBMO3QGZZI1zz0WIvOb81mKA7BOAYFQLew0oiSXW9c7dJvCInIHyMYqc/xVKa
XPkAPIFiQ61hUNrlqR1HFmbx/MGRtYbmrWTNn87+I/v/LtUWQUa5Qm1QxowUnzGUodg1IyEMpG8u
3orAcMeEwPHDsTLx/ji+LM7REHn42R3JWR2U6D1ITOGkq97xwL93Hz0rtbdNZJ3nQUmTbm0gnrBb
7wiMqb7OD3dicG7WZMlOmLTzQ0j3wXhDU1rBZvRNer7UJDQ04FWKZE8wso80ZmEnDhOWZ/HndKk0
oPhRddk6ouT0B8CwVMZ+ivoHFq4jxnjj0hnbW8op8px77hEjHwl5c5cwDws5OuMt4oCTVed8zrzu
6gZ09ZwV8l0z4VuKtXPtKna1Unnb2j/imb349TNKn21N2oymSpwm94R9ctHoC9qujFFBa97HdFsi
IG/l/4okdXiLqBRwFExPUvLIhm9PnsJRPRG8BQUxCavPocPSfXH6S3wPjoHtl8Jwk8BAwJjv3Qar
11DtpZG2Kr8SAmMGjSzG4vxgYBsVYVCQJKbh7rIGXcbN5olhE6vj6W8D3weGjTb1yAOOo0CZYCqA
0wI3GWFELmuloqc+67eF+tSmxX9jistrKJueyT2r+oK1jvmj0C3a2GURxv9/9Tqzgjen8F4lNF9n
nzNYCS8ZaVGCgpdbk8MtMesyiJaidmQUK5nQ9HgtxuwShDuKNGzQhePuGVRdYo/X9MaMnl/PfVYC
9dE0xLuYBCl6wsg8Fi5gOHSEvytwvNoorQJ2XlMMgZv0nBdt6bEnMV+U4pNQV5vPZvTAHbp4W0wa
FXUrl3thTw1sc1F7rejWe46AGfDUnU8IgI0QF1FO5U/UF6AFZ/tldTsB4ov7hNPgNjxzDxslbgzG
uduhidBAH81RiXiN3C8RVNQSUeqkt6f1oVZxa7MDxOcUrSdZia/vEa3xYDLILdS4azMzCNgHuGgL
7AK+5N9YqMJf3UYMzeA6VyyXJzyQXH7xPm2Y6hWlfjg1W7N2rP6Zn334g9YahUi4J+sM2NYMWvXl
GThHkqJcVxfUjWN7GWlav7lX230nQfbLKRtAzkPdI4FaSeJJ1MNPxNC6DmpaFW7sNHlnythm7Xrh
7xYWxmMhTpljuPx7qJM0smi7w0IOXcEF8NTUqTr8Xt9O8rWclZ1LmlUFo9U1Mh03gDtLIGiG4gsH
+1xpJuVDea5+UQx8irUA0/ZHo35umISNSGS9Jbstcqr/WULKyBh7RtbFhvPYaHuWk4WyCAiRh8HP
Z3/79cRBo2LoQhO0TcLsrRcjoULUGkEtQZK2OsitW214HEpOxGzsk9ZSSWWnW0iKS6SO0CTybBr1
kVmKf/svrebsKbIA5rurgEWQMWVkUJPBgYywDeJYJ56eoyOFQQdmVK+hLS+GV+81ULK56ppd+TSY
EqVK/jmKy4DP/gT6WReRHxuG4SYQWc95T1V9ZkAOM99SUwBMOKG00ftMVJVLd8woxwmbk2CKaXdt
TYf7mh+/KRJCfEtuUtYstsXwrkknGYfJPcNsDv2tfOeVVK2wB0U4cCNmPgvbGNrD63CjvyOtjkGI
eq2400noSBg8H749OOClF40bPt3m8iaMpGuyrximMVLlpaod8JtNA6n0yVeh8fgUrlJv/6Wc6ILe
/s46b4Xt8kmcFD+V2vH5khPMXLD9Vh/ISuINzvnggdWlqYL4Dhm1esGtr8kW4xC0i/EqTPp6pBJ+
b0y/CbBGZNCcAyqxV5EeePSU1b7+LKbyd4AsyiyQrPwisUnuLkyM3FJCA3uPbKPgNORrfaV+xW5H
OYqsBEakn8cDmCwmYW98WbfjWTzX+W90/SpIlqNcr0CjjW9P0K4dFMTwyFMABV8RdXU/TO9nfyRO
pix9cawFG6TfVHIAtK9raJUAEwD3EATTAaJKUjFv7Ky0liJpPtpiWM9iB89LEuTcElkUi+WHY3je
xgN4d6fbChX2QyJk3GhXzg5iJ7Ngxg/RtEevBMZpTKmLcyQhyD43jkxKgGxdJCxh7zCu2/HWnMZe
HckXKQp1pT/44RYFSxE7TlM5OiOr2mFWDD/qp2rVii/BtRWePwdgW4sKyElmXEzsS8kGiINQSxQb
iv1Onxbc3262raQwVekQoDcn/wfGcckP2QcL6CAPnrAt8dFq8j//G4Z8bFrboM2q9uYrqr0y+jrC
VsaEIFnzSnedwEJ6KR78u20CqAVIe6um1/7aowCge4sKtEU79sVGFzfYyiFGcK2X/66RyjfPSR4p
8U7zUh8rmoYh5FzPaXj+rydV8flFvEZCF1mawpk2RS25e2iUbrfTAplS4T6sir4ht4o7JbFZm9Ao
noO1QTeoHZRbgA25nB4VtMJllxZPAnJDu/4Mwn8wZUcT/dC5itm/t9mXhBNsdihdnCyDU6ybMyFG
tkh/CcoKeM5lHNZQALKFAX9xzgx9eKfO+2EGTOGXx6ztlBD7r5pmt2VbphdNoqgZ6HtNg+WVdFPY
nO9zliJe7dUOhGQk0oUilJELclH6QYuDRYdeNPVo5AXcL/K8/+Z7x/9/sZSLOIaoHZoE7sPCbL+5
HlvU1WdynyYLBB6Q+mll/+1Uc0CxNaBDqqElWKqnd1tYQcZWD2QrUbAOITl7SEJ7Lv2kDVpm7UYP
kvILQtrOyVYR1fB+wRZ47yUftXAXY3e8P4+L/v5ubyvbKly3x+ryW/mHv81dAzTcj7lShrNW0IyC
h91CoV7lG7iUX7qaq3PZxIgnk+5GYCguDI3KLmcF4XFbgxIGq/HcjHZGZQODlhn0dZV3mp1k7nN3
wsdUr0SxqFG0ni7wfPClD2wNbRS7kJzk5EW4JgjZlXQ08gxKcxUA1ew/kyfQ/Nor98tZUyW3Gl0/
05D/qMob1VadWikvJpMzQRmd8iwbFggCoD2HEg37BVH76PwVdzSwFSRQ2Quz2/deivZMj2LMAklL
m7QOpSJDJaiNdw+QE25DPno45zoXPAlxDFVjRdzbtRXVy5WWY3qZtGVW4QGjueM23PmBWVycCqqm
3WyhZETxtRHSXiQCIlj6pcMjTUSlibfoxNYssyYJeEg40ajUcpkc5GuOUDAYqNBAzuHYwGQsLRZG
gYTgLDro0wpvK3KYeVLv9iSH73Fk4WP1VcV92kuDsge5gDjSUjKBhmMFiF+2uGQe8lQqUf1KpefT
SnY8WdcPzooF7YGQ16FFSTXdlez34wR9faj2BTMsDIpc5hA5jmSns3t7SEzgFCLByeKykS7Wod+h
6X3cV93hmgHiXwEzY0dQGcaGK3T2MLpXsvc1HzkeYka+pRhENwvXM9dwR+oG4TvLT7G8zemMrutm
KOrZltdICb148yBzp4jEQOAITfrR1zw0VaALJ2uCZmyQ8EFRYlqVn+trL9mvzh3Gr3i1UodHda7m
YyNiC6D2J0apzYF5/p7Efj1AEW00ijwI9fi9o1RNyVzcC36TV3QoriWRx3ptTfIh2spZ7tfxRUwk
sMhs4MD27sN21PNFlAw8opuFcBv2EmifxdO8W0jyOfPjFDJxlyqHzFcbpZuBQdPz5d7kvDscrjMF
/gtnxUdm5efIuU41xuhUAesZSDaZDHx2aSTMsLiSLCEoTfZNfoluHhzioJ1f4hB1889NPzaMmeA0
6ACOAoAYTqfiddI/5Y1M99j64t+rnj2uyiuDgbSYTwEjXK0dWwwSWDSPcK/xy3laPwT67BybonHS
GHngJZvAiYHxgUR3iKwLn0/NKin9Grtg7Nsgy9GUEVehgkKKE87JmyqrV+7HtQQUaxtLJwZrYb9Z
uLeoq0sEoBiSX3NpbpBvzRTeJassZzmf53oy95DPeyARtqgxA3YFvQSzCG819HCXBEDWoy6SXfYA
fXu7ZYLdNRMCyF81SbDgfUwpb6AIG9Mw3MEG85BzHVW0KAZSANU9F9Phsf0PF3t6CZKb0Ph4hsNo
ddfqVHmNfFrsQzd5+oM314Q7HbxmNLCO2Sqf7mZ2FyRoQ0gpnDFz2QetQhNdH9ySL36T+YZ1/Ht5
72GJ81Tu5V3G2r2NIv7JEeNcAdwwBRh17rHCdtFSeeDvqvIrZzHJklgY31ljFDAXIalaJ2g1kyv+
OOtOpr0N5/RO1cOpti12EMszLC+3Q9BOgKZKs6MZ3WQqWcOutzvLM4SJ5PwcR4+ZWb1dlSgtY3v9
aIYzmgMTqFzWnJPcSv0Y78ssKQIHP0u3uMFiBnpeZqTJIGW8eRYArb8xfxwR1huwy6fYIL8k+okV
gPvZv9M98K9VGa918Kmwios8EIIEZ4DVwmuG4Wsae8w+N+lWMy0+UO3hIAUny+kthYJBqyDjQPq9
EqrVtnMvnDHCZsTd1q+2A6ruWccNPcQY/l13kjJRIR2zzx/auyGKRWN1ZHH70rc29H3f5+3XF3ii
gSqu7IzAc47N1TeCbY5JELoGHPpo0GcZMlPzcmfBzc/JHZSIQ3oMKjY56shZc3vs8GTDrtMrVkKk
XZDKtwS66E4fHXVKi0seMPuQD23SzWdLSc377jIo7pB8dXwuf20ogoYAy6zZBYLUEfn05gBIYI9Q
7prMk6NFQNc/Ht9HarYalxe9DIBepjDOGJ7uz+fCUucJUff7/qhRl+hG6VA8an1xBf4p+d0cEAAk
88w25Zjcm1e7o7vTDB1pXHD3jJrgDU3ysu3A9vJGzEzlZ3SwBDBqrypgVNLnfj+Qn0Wutm95A0ex
1TBdFDKyMW8AtQJwRAnUVLdm7PxdYPAtHK3VWxJcZmcE7u6ly0hoNh7wuUDYHLY64GCi6HGYDsIo
xypFxuZVuGWoLkeWzthAHjkK8AigS6xycJRcjJfwiN1W7hlDJ7A2ky/YQE1uKesgopgtFLqPZCSM
y3NWZQ9+Ch8uk5EP3gDKts4cLkZmi9G0wB6OKSVtcvPPMchkXKw0+HXrRgvFB3RBaUJqEc70MRzV
lpnAC5f5DSYamQ0BLwCC6BqvAl7RpxzUfOc9GrbMNK1oZ7ezP+2YHuCWeuTjsODzehEyT2rW9aAj
g6bmwG7fzs7h0LItC0HAb6g/SjICEzMDHjpd40efrpWrLwbOeOrScem2bVkEvzTAZNNaUmPUTAPh
MPOLN/mB9AeoAckq/G3NtMsoXBG12ipDEklrSZEAtyfDVFfVP8rJq2SFXucVopQ83z8C8Wwy+IgF
o6xUFT5N/qDrweFkRhOOx46g/GVtdfAaUzIBa1Kn7Dr38BHpdsl+JiM/pwzmfBe1bkp6oVxwrWnS
FeObQEPasXvC8egGWw4Fiz+J+wefb7/MtwIQay1mzCr/64GpE8Evx17wWc3jjem71LEq9NMPcWQo
SnM8Ifux1jcZ8o8+gth6vdaGVMzXQFK3z5X+oOC7JYXQ7DzxUZwkaHlWdjYKj0OvXEy8UO8dZg+Z
DYS8kc34QVq1vXRWdb9COpvcyMpEQW7JwBRZuSWALG2bguqD3ldwRrhftyLfZGDNkSGy6ABbRZ8h
OPZV2GC3B7qRfSjjyT69Xpajeqhtucs4lNq2cxFwtsk69S9Zs32GBc2ljKNAzZI56ePzDmNQjQDH
Fejsous85+6AJdwLnkf7DGGvIitpp5XYNIxmYUL9lzRqckjRi6IqGqUdujVEDTDQH9oaMKrBP6Ax
dp9hvpD0sohxZTLN4TV9rLUladvuQQJHOEZtbKG96sgKEUuCYe0k2Jb7rqRWnf1yddIwRQUI+not
4UBe8cWFwXbBHn/Z4WzesTZ7T8D+/g+NUkCVdJSC6wsA3fNh7KJOuvuOwGjR/nTUUH+7pibr27Xm
4Q4nwAF0JojXu4qTr/EiECKoKDHB/p+KG7ljfUC5PmAIL9wed62YJltf8YGL0DDoqIDvyVD1TkQ9
Lc/80w1GB8ioFkLmSAMcaTgoTg4ZVQMJfmG+m7ZQenaoTv1uVXRZ2M8Kpe9C2bWpsQu2kYp4bs3B
Ez53SXQTWbVyjDPQhGk152GRifLEYHIJbr836rWFCaQwHR+LfNNfDM+6UzRS3MlpLwEcWVhX12uR
jKwXHDq9nS3THjPcA5I1IkVEL3S25GgwrPC5FHIzF7j4K1tVh9UTFU1268Or9wcR4W916sxP/XAn
pNgCPnIl579dM6I5oofjYOYXLMfA7sFskTfnITxxG/s83NaO/zAL0O7Uz0vk1vXEaMk8D2BzQowJ
uItdJKlxkh7QzhhOcvg1Vz5OHza/sOAI6UqfQ2y4iisDrgmDvf0R7JiWAgdQfkpc6h9Ndvac3SeC
fEkZczc20SRjYDlqshH1cr5tZlFMiF32LAsH+Qmmh93KYvvFjbCTTiBZ4FIWrXKDXItmiKknGW1+
0YBh1osfkm5Bp9CARtZp/52WNw/z10Ig93WogMchX9Be8yK14cF8y6gcti8+52GNwRhHtl/3Ktpq
JEab/8ApWBvFB2fDNTZBrj5YB50tBwmFJrwXp+J0PzWHmUO54IWiYzbFviimtRQDf5uGLVkt5XcA
ptW9B2DuRwOYja3K5fHZTsdlRiWpAUB/tGffFLqPqyEelttd81giKdVYOqW2cWDRKijVopJ0IyF1
PcatgEqIqQCXRwjfjN/eTkoa0J5TjowT3ngA6UFWOmdLxRtQ9Yc6v+Xnqjx5Q32xxzodYkWdaakg
DPd9w/sUIZIrAjGxw4Y9y8g2DcCN3h3r1qW2zm7lq+trzPh5SZZ9P7JIdJBX7fkASa+ujf1ZtAzQ
fEhQat29aS8U2hFgKVr/AjSHaAeeF37OYnMNbxpFL9rT1ADDlKjezWlU6WNXwYe+r00F46ry1SNq
yHfkstff8LBsQPUXSwWgONOZ7QWaqwbwlFLSPIWxPmEmezzm25Rx68zVguivkAmZ1cEUYPIiK4Ox
VcU67qbwehAKQiAuhI9Rq6YLvEg/00+94rOQHY5bY/OsXoeTt/aLT77/6exVUoeBme9zHWktEys3
jT1fcaD8MeKtNXcXXsGUyiFG7O8I4ouDYM0mlfktWZ2HWTCoSyQneDrC49w5orhQl5/YFH77bkVE
xF0lYTY/mvPhDZP1DWCf1aIzeg==
`protect end_protected

