

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
HpfjZK6WG7sYhkvMgAngy3z+9zzwD77820wau9oTTb6dakSkVNELcmI1vCDbEcS/48D2LFxL/qT8
BNFOIZ2d3w==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
VPnG2AZhAX4ivH+F+USmM4TuIe2lYrNUq3Xx5puxPaV5guza4OeVGJP6pYRxsBYzj3S4OGH7b6n8
K0l2LCX8eil1TGx7VbJh+Wd7uUD2r86y3rluWkRdWUlHXjFOxoCZGO3zP09eR4IRsG+JxbSDSiqj
FoMAGfR2zks5CEu7dtk=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
u1IQ6dlJ53C6R12Hzl/XoBaoEA3n6gOO0fxU9jZJvCev68EW7XPnj0pNHAKpShucryAUuc2FQgbE
BwIwQ+0yjh3dOW/yrG6sHXOI8NvAIzuE1LMkRT00JCNCjyt9JL0PrhVhWC3cY50b1mAkSZBVfMWL
G4c5aMtB6wF50NpvOm20Ptquu8OAMlN0E+mHAN8qvWTR+CwIDUV/kvH/83yRaRonCOBULUP7XzwI
uAjFnciSf/F9eC2blbPxLHlWXLQDQaZnUw7NGNc2Ufyh7lsh0GoZzefU/JIhthv3ktn09r568XNe
kk/w7iRo/w4FLMicA3dbzrMyZkiVt8z4I74KAw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
x5ctSMYno/7jD9HwXtHguBvqXjqGDToxuRubQZySJLeTm3iuHlQTdlRRlvw3jNvFx8WWN4nEmWap
sLwuJFUESklgDZc8wPsu9plvibxKvIUprit+FQWsTY564IYlM9a003tG4rrtM7zZ9yfolbWe2MY7
qJFpoVf6XAxMMDrPtP0=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
JhbANRgOr9SOBKZDRGJGrZPWNKSEG3awknWUR+2QiYueCqJ0p8+Oq42E9W+XtOMQqS7h6dt4lJzf
s2rJvfuxWWYMk0rVRoGeqNzUfiVHbjHTaPdjhGKzIm4Kgu/QJ5ooRwBflBurdW1+74PtPtKpfjcs
79ijwPcRU18IbRTlWf2wzAlLDLkDUewye6if9pFfqGP8EVIxQIb2A7LmwWnM+VpfHc6KRQhcdZbj
LsxdBzKwdjN9Cdt40472gpQEnBtaoqRMW+4LW5rSmhm7vTXSum0cU3Afl+AWq9hUcVWPcrWeYdm+
aNrNDk+A5wRHt64iDTF82GsVuvkYpCi38y+ffQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 12144)
`protect data_block
kLHGNvVM3MIjzCRNBzElxH3fW9Lb6DzhgK+wKvq2tFGXXNKDssCXGe5/7cES1rN19CTwtUjh6Xzf
DYG7LKstmCnbjbYv1LAh0OVBthQK6Plf3Wovaa+PyB02jdJoA3oyiOg07tIHJjCWsuuYG0TMwLGD
CbMiTPLN+pAF/IKOw4s9XiW+gD0hrIlxdJ7rjMB61/+bLLF55qWEN4ciMl33++YBvq5QLtGUzgFh
N1GlK259fnYG9yx0ZBKHxm+29fKLX4kmA5VvVkWTMmP3wAgEQArml2sGJQxE3evpkM8MOpUcXrQl
SSe+VVwY0UditvKrO2BbjziVoBDBmcdzqcVD8WwLmTDTPFKPK1MO4UiKfACLFZ2sSLI84X/p2Pev
YqB+vToYDUL8vpadBPfjyYYmRD4LJsQM/Q4alcYKyFmLLfvkTTPhrStKLM71j9+pSsPWhux5shbR
DmUKWGY3/EOIar7s7g7kKn2jq9DM7HwRLoQHXvM96hjN3cECgfh7R24t/YO6ZZ4clRO8dreiNmmK
siHVTFSMeQ2vuYbRF5YK4yHacQ0WujwdShIi6f2lGhAkJnaOVxj5ZdgtTK3rGO5biGXVxBE/oSGE
zbnftnku7m1RixEvzdXAoUoIhOsxhF1Mgn73jY26Upk/DJcKJbgWMNVF5rmtZsCYoGxooJUUj4Qg
+SLhtNVEOQhabn1ZrKbxQwMwNVVC7TNslqFpmWJIjfcY5ImkeBxOZErq2o6OO//1qbR/pAS/Tqzp
ICa363MRCjIC6Ylvpt6K9pg0sss7tSZQVwKgMMBZxsNzrJRnGLsGzzYh2crnMwoU7o5hxC3CvPqd
0nLvwPRNonQKnZxn7xYRGg6C90AXDeA7vT+eaYK0MnXl0TCznHlwN+m9YZ27p8902u8GCZXlpiWl
opPkcoByYeZjMU/g5nElkQAd451rfNmpodiaYOatFopElYXtENnruM8FZSnmDcWiTxKJVlUVHbbg
Fdmrb6w3HKN3DPg28OcxJ36CENfAc/KQ1HO5Sh9cw33/bHsd1uKiqs2aaFbR4eoh3owxrp3ESQiQ
hiVxf2hjpPJQb3FIVaXEC3T+P+xje7mEHBEjGKr3ssQHPxZt3D2AqI5A9tBHTd9fXnstQxukAfg0
cwzzosSMF1JEBQRKRy7CFFaxlCY2px8Y+i5iwrcXC5FvkCrvggWWaYbGpIdKHD12Yo713SdsK1YR
jNy4VHyvD+UgHMFdSFMs+4PWVMv4clJUctDAMmMxey2dlLiKstbfcbtQi+5WknFj1to9JNHLsjAz
5VddORSKZGWSpJz5Y4t1MZCYSMHuIeTXLB3L46dfF/SpveEDkajrJqKfiL4khCW8sHH1pZS0SNKN
F2c1nZJP00RCklPIklsH6BDINZHxhZJ3UP8bpVMvc3c26B8gzYVcw0wvMctcBnQLYOr6mY/rM2Jg
077hmc/eLABwAKAyo26+QEf5YekTKKz+MCkKqAjLDZVmcJnZcVjQF1lVsM6a+61nmGenApvxmm/7
pHfQIPS4467wkPr5yGwX8m92Kn6sS2qlQAD0L6iJ+ZMyUfzD8NEnros/OPNEPXq63HasFhHQOIRL
l1rKWY+BhL7pzbRM+4b+hMdsPNz1EKd/eoNa8vswb77f85kPrwKPS2ck63xwvxEF1LXlVdgioek1
FC7llSA6IxmjuaUpG7hnUsgo/adZnl2xfOpJdMxvrdI+dVDDFIgVVb4tr5PaclA8x4pndGBdaOAI
bkXu1mpZbdFu22xoA0nYYKPeZjHhzgPWozBODyO6PDgaseYbKCr5/6ZLnZYOt11cAqR3ZSyW8/d5
hwdpFAyVtQuakqpMMMZ8hCKbuxbiBxy3EZJxS+FCE8DNFPK8d0tLpkZMpXS8VBFadITf1y/LyKXl
p5LFFfcNc+G4oAnYPB7Fj+75bdq8NjOs5eQly0JhDqMpBI8++dHHjS/OjxRQ6mqwizdTztd+GioP
GzsRqw+6FE39JczBadkurR8NUkF2qJVOQFgkNiU4XkzA2FAK/sf9fao/NYyWtZjwETzWcB71mVoO
TdCl+mLy8dasIFhrpKsGL/2nAByANTm6ZTAaLeUGH4rhzDmivAc8/npSJuCoHmaaWtnCUkCOKBT2
nudwDrqMipKr4LzTYmXTdFErNeD98oCxAI8XALBTcQfMIzaMKxsSuKSqYIclSMdi8xORMCoKmmH3
bnfu/iyide6Z3OxjcX+OGrfnTYloC7aYuwclG7lMe+9ZB/r+p1Hto0/4wkOpLwgEe4z8Sh+37Kcs
d1pC4rR3ELCGu0d4RwGn7W6jTV9N2LI8Qps5+oU8n3aIXGDgzq5WbfVBmIbBDdrgrt5vWSgv/8t4
+FzC/K+IFi/Eu6X8GaSVvs60d4tmvBExcIKDGzAV6WzHBFRDOzhpGtGcBnQPQUmW8zyGDXcz72jg
HMNIdBNa9rT09PXzQfJ0tmDG0F1jH92ZAFEOTxmY2F4eMMzHVbCm6klLgH6Z04H33tKAdQ4naeu3
RkkLTPFqIZ2SZgOOSesKwmiDcSLrDcDRJYMt7iV4Nkk5XTcPdQhDm1i1+H13be4Qbs/xLHDreaZ1
lwb0yZgf+XElBjsm4hYcwRWp+NA6HSiUE68xrbaSmF25Kki5hC7o1LjGNeGG1RFyJfVjXChSWbxl
lF9GmIJUg+9NNdBOiPfpMjBVQXBESIfRu5Ut53RaC57F1n86tB8znWJYLqGQSvEet9Q1UMIFMjku
gaGxxgNArF2m9HwE9oWrC599ExGSHx/8PDrBRWGg0p5juhJleQLWbN9z0ndjuleep+zdxLuHy3ID
XVnBMSxbU0VzR824G38QlywoJBjN0lqo+4scByW81IqAZbelLGVy45FplAdGRoPLsmRGP0xKCJTV
09UK7E7XGv4yGrXnum7Hm6IuROWiB+ZJwrXHN6DXlRmVSI2kmGlRBcPfRHvmA7yBfP2bG6wja0qD
28PSAYGJBzIXtl3o7VtV7dspz0PGIczMHf6KdopbtW+ikKyVetJoz4ZKXaBrSzeO4m8FCsXRdMBU
NTWkcF1q0UnwRJis/AryCpGfPRB38K2gAfTXJtm+Br+PEVTfi+hJjPXif7UpSUGpsYA4qNFRNpdN
tC6a9rwpkyYH0Z0wWbWUUS8Y1pIpA/62ndfEvYAPNclQA1ZvvDCGu+XGc4cQ61PWbI/BBsPfL1uC
2ugh4f0IhYIlxSWcBOfsWudDPxg0hkEEGAAUcl/JsTgxzORl2AuQccCDJ7rZ4DxsHk3hD9C08l4F
vCSHQibQXi1FQ+2JYDUFp8QTLODPYQ/LPWOjys/P4caIq8tPBTRJb3rCRepJz0bix6j5vMk0gmVO
nEiJ9X+hlD/1tQRTjadxgOD/Z4BmXZwnrY6Jk4Tk5ARG2DDxoJjLoaritcUJb2TSOzvYJa3V2MDd
1kSjLX2Zg0PFNhjHXwemdM8n0yRAvKXx8PS3f1224Rh9PwKj4R42TjmhnB3vuPHzpfG9jVo0sae+
YUHIz6mSYdTl7WiG7KhwknZY5JzQESTeuO0MuF1MD0Y3OcEfGM7EPsFboy1WKG/4nh0UniE0oXBU
08qVqDRiKlhFiuBHFvqRrvSdcwo+8GPlMup3+CT7yoboTTYbRp9F/PJqtcSv3GCuaqz0esEjdp0U
VQt4gc40WIW+YXyzUcMbewICwyADIMN1k8p6hrpwNqHyn0CRQQA0t56kftFmlqfGl5hUOqtMq3iF
tX9fTP3Q00zHtVmh6Jt1SwednBEWsWoPKczwUAd8dgtrna3jWIL3zOPXzQVz9uVWBtQwO2frvx0+
soLZOvbJYwmLIyo0IaOXc0zADsNMxH9eaviYHNn4BGU6ESVTQtK24KOIgt8fgJmHkBhmf1na4Tqv
ih7E4GPuFOm1DJr7ZRxcaYttXHzJTa6DCIvMTmkulNgtr3b3Og5yyHgdCuxxRQeaqr16QPm+J3vS
MsC+uGtXbQhTTmZ0ld7JgzuLwGma3h1vWp4bs+3Ff+ndGCFqWi6kDoisEGpkdOHsV5T3pMfRPy2w
cAsjw8Zyn5E8LP8HD0AWpPLzmeICeAVUGuCojfbsHtYiZazawaVHtcB8VfID5XR846lzy/lHpF9l
Bc2P9BQ/R1eecTCXYWhnOZHvCaJ7T9cUPTjFhRIDaL+I1LpblufJ9NL7Ly/kWP8icRfaKaadiF6k
IbdBzis19AVQh0XJpHPBsIamc5oYDxQ+s+CkNA0Yy7NlllK9/BnJCOmLVqG3WstwUvJbEvjc7q9I
FRrg90JZC3UrJYpGcFkfuyOzf4BpGuL09XOTFKNs/z5eXMUNIAqouIHcPZrzp7rXVrdvdT0ELSH5
ZwLDAiCPu25gEkuYU9qSF/NRmz3/Nom4BvL6LDWPY54ROH6nDpn+zmpfbUV87wVr82ALptx2BRIY
9RaoppZT9KlRFvfmSn/dxxgp8pRE233sHesLSwDCm+EY4+TCUy4WFo7uyyO8GWW0ikxGqqmnh/iT
Jf3Fq5FnfRzw419cUmgFzrDBr1rbBvwPxrJWhId7aj1RR0w0jyNFkHt/HS1UX0J07ggT0u7u4uvT
JqEOb8nx5/mftOxjyqdFqjTg0rYydr1KX3b060367ENdwM8YZrSsNq2ZuQfQbI8yF904JFz6I0Gd
fYx7WiNCOsURuhQ643xDmP7XvfZpTQgGCLW4C0DVonxUrlU6EAYIWY4a0NaKWZhq8VCCeO8OcgKb
XT57P5dqaWGHeaZGdE82zX342eWmlTiO92IZZiRw+4hx+uzq8iYFz6THAfSEYpoGusX4uPtmWwL/
1hsNKhqIoppXgDoghG7IUFAAdWhvZJanxXm8ZAoIuGQfvQ2DVbWUt4WHtaVvnkZJS+qEXyz6daQX
LqsIs1982dJAyYBBoOqfrwljbuR0gtAvTC6haxQcLKmNndwB2qdO3hEvYGXrCt0M3O4GDFH57ZzG
yXdBzrVnFyVB9UcMbaUx7/OMRh0s1nUN3xqI3F7id4fS8O8PANm+woowlDSet8KOrm256TwT7izf
OfDYMnDWAjeeQG74TQYHrQvX/YPAqd7Kw0aMJezQgBWrK5mXCqCpfr7ZRvFsX1FENuiYMPxYf+zB
wscosZvfX1Eym9UosuSEic6sxmIw0XIOXUz7yRnR+VX+kN9xRUyQHmyVezzRzoIcP97R6PLSm3Js
04kFC9roPVTyk194LkvE0vzZuvMtdo8rnT92mJAD7QEbV10JCDeNiRkXXKKGDZozuowWw+MC6cBy
FkP5Vcl+yv4DfexE1Mf6ZxID8rJx7zk/o9kAers6Z+BeFiuuXDUFdB9HfnLp8E5/QPt4o6gA5TbM
bS9J9yYYghLBsGEP7+3Bz8WK/0XeIIpu5Resi1NLP8CfnpZCA1+qBwJzZccQzJQJaet2OFR2/yNs
ZMv80NgnezgslcUA6fBVVkW5Re5cOAcQbAdMLQ4BK9vFOFMI723d64Z2oJ1J+eAABL1DwtmkLZPG
2Jn2+VEppHTsBabyH+TmqQ4/CP7GqrL3NWUmX2fbC8p6Zdn/g0isWs8oM0oYES1hlP1pNVOSWu6c
1o1DwOaeItjhU5Rfn6M2xcsDOIl2FhwGAtwCV2ZzjDDD1peKUtsQAY5Dfdpj56yKKVCeWBI5rPCB
2iDd3SziT0XKGYSu19TD6tlWGVnT4ykcHSNmqzCRPuiM1XIaiEcI206xhjVh7I/1dmjm9L8yNnTc
ilY5IvGmGtd+Vewn1i12jDVyIus+qgeQh8/QKIgv5Mgt8hDEbVu1ep4e3ocWK079HWAbwdflGfIV
JXZfQDgO4q+Q7E6RkuLW3vhDBmw6ZlcrJZZo2w3habflxjNTm+3RbHt/2LTVoa1DAqDjTmhJcWIl
U87iGazUlP9CrHM8i8l2K+2cxcUE0JtP8oLVj6dhLbQDpfs97fzKzXMQT05lfuDWv15UntiqaaFm
iKELUPWWok7jUw4KYrnYdzagHmOf0E1tvbVpZTs8+CcqZsaPtA69dqhCEWmPs3Mkx8S8helADCZ+
LSCwiIZ18aqppIfbrArfAgY9oWpzgZz58W3ota8+/fsEIbBzBXPW5Iq/zAc80t91RqZByO9VOa+o
oMOS41ndpGCGgz7c9ulmkEE/shYUeKl87qpYoRYbMiu2msEKM5fQ6NnBrq9T3Wei1uBNLAI49Y6l
B1WvCcgk+zQMVAJi2fbGIJ3Xs8yjKTPJcq9EzCz+zHETNWjgwGJRWhydA59q01J4VNJyvI9tktmq
UShxcrNbxv7RGUWVdMs4BX9rFE/4Ld9UllNCU8IJ2TPJEISoW1WHJTeswmonC0MhYyJe57hrjkoa
qEursEe29oRW5C0D2nd8YrRhVcUCyd7N8dAuKhl2+s5zaBFZE+MYfPMvxD0RmhJu1qLfpLtGPzac
paNYXk6Rin8ST6rR73qM6q3+e5jj08ESEaITMO/wVSVkf34p5INUeXu0EHM/Q0GoVvHTOsMgktaS
RHsvzC50dzjBY01Lp1suFF+OKQUqtd3/UjkEVPcNfPO1netY1Yy72ZlauuqncPhx0zRJDwCVSIOC
che3wfOngaj0XzjQafGHoOiT5yzJj1U0IlwzdkIEFU6nRyRnb2DL83FzPwEMNdI8vfCkoTHHh9do
rnhXVKOi7FKO5TbW6596k9C2hbdnt3NunYmThdlykrtbEY66V4NjmY/fZrgImdAA/7VH4lidLam7
6ofR7qTLFvpk2vkOHs+XUbG+oNwYnbaaxkJ5Ipyb+a1/fGPMPla2PYlhRK+IKcOB0pBiJqDWAOdw
gU0BryHudZORM0HZdBUw0hkpXzqEbSY0wqKS9r5VqDmdlJtYcXxEz3oYdywvxIulKRKk8Z9J4mSs
O8LdGbhldq4wNF66MEWT0B231mL1GF7L1xyRGrKIrXD4FgEm9E6dz/iA+6sz26mCRlNFfq3xQmWb
A4AddPCDzsWxq+gM7cNsh2cOkmWVBdVPAKzKXjgS32Qwv1uIhmmP75xSbHpw085zLrSsCifzW/b3
RPLG3LNAWuWph9zSI5WlxAz2X6sg8Ks8xeMOpYyB+QtnG8YZPIaQ194LiX9dOLO6m34xMhs8QHj8
UweH2rsbMOhwGgYSHLeabvMlkWNqhaWnI2O9y6eq985Cn/y1TOHHm886DR5YO53mQD1l3WM9mc/B
dLkZ077eeYTcdgcRj3syKnZi3ziAMNkg2e7fEdFVjYj+4t6VuWvlP/RTL0eyulrQymUm4x3lgBvp
60vOchDLymkXQrQ5DASzJ1CQe7ocaowXHkE/+ViQAd41lX7Lu0z5R2I3FbQXutoTtPC2WLC1FFRY
TXHi6lbonghIy4EHgpW/n2VuBGxGvWU60ucRr+SkJcMeAos5DbZ1O6w+//+W6/0MLCbLvksucbZ+
f8DrDAxui9+F/WiEitJEHYyF/KN+2mDLwYgW67uXtz8bVHUJqr+X9o50Li1mqimQrcyzUe/xFSAy
U+TPMb5KGuf+yEMqh9Qcti5+jS4iocoUtqtHz0U6IRmgNRA1C+UaaFOYHsZSGKMIMm50rijq1D48
hlum3ADsyV6uxQkmZiNRxmVFVEvA+7TOWFjLsRtDtSsI3KMeeHb/I9rSXwlEJzMQm8Ay38kxXXZX
lW484wXQU4a84lMEfjOT7cCvNhUPwFuY6LtljnSUaKB+4aE7Q88qiMBHXA4wVZnUpK7ZMFBX+nQv
vLq8i9vSM/wt2XXIbc1id+mauC1/ScmHKn9mWRgrLZyIWVU4Cl7wgb2b0FZRASYeROOfkCEtYBxZ
1RTzxIAJGowDPkNDbsT/c2IqzgtPKREfxrckCFWzR88BHQs6CQvbr8B71UBvBuYd/dEL0StfccSz
2+irJnvcCzd0XYFTMX4QJ8n5azHZE+o4hcnDnr7Sm3IPP4eiI/Un6bCMwFLzM60B1EiCuzj3aZYW
XDVrDLoTrWlbRdp5HoukEph3zO/HbHtchv/Ly4D36FPM9OJFAuc1PEz5OJAVSAg8GdEEK1ptvZ8b
fUlQAct2tzvFhNKjiPiTRs8Y3HRipHXMZrYQ16r8haJHrBoTIIJs0iZLoNFTV9KZI30irBUd1oPb
m2aKf/UQGFX74xwnhL+l8zwCb1A8JDHOFjzDnnduZ8yseoQtJBhzPv8uVxR9XDBUjiQTaXvwiQI/
T8dzlHdMlNMc06m7ZyBEw/ZdQem06cv3uM2lFIl9cn4Qmar/mpMuBDVLiUvZCarfW3qNyffvQoTA
ZBTh0ySy7iKY+zgDkfS0gQ0cJoULqtl9iixY7eBD/PNyPbOUPuT/pZpqLdd7BC9hxosVKi70FaKw
QZLMeAawyTSRe/i9d64Y4Zt2EJLWLWZ4SeSGCCfKADYwnMtXnUNt01EuOuJglLr1WgL5L1+7mp2d
CfVFD18rhxIOYWHZanQ3Y11sU5IbaIALnrq/P2fZKR5O6aEaPxBnnDDashQXM8kdo9KqMqi2N22R
npUOaA4HPHkJr+sEy/C8mv1wBgKEObwtbf198l8mphbId1L7Guts05DJaAJ4IG3dxZ6csgyKDQy+
lvKgEeleHgckTLFZMAboDiyKFyTRPGLwAQcOxzIu9YwxXSy97YVOgJDNdREgjIA90//mIaZsQjkq
3/oj2n0Hn4djP8ZCTpy5qJJShFzzPn69KAcUV/qyq2Q1L0jLydWyL1imWPajsXXpoXhesZW0n2FX
7/cytGxmnltsVkGv21jqDMtgbXaTWARnflAI9Ix/kzTKgICnfNx00KTlZrtLWE3/FQq2wd9lH+Bt
dRbkAfE0uCSsTMBiUjp5s9N7ma8V3P6VruqcWRxo0S/wwK5z/pyBo7GCfOdt39/5BZwMwHGKY7ZY
6n0/fefMc3Vawk7/gOWRGG32l6SrJFRKW3I5NR4xk0mQs6nTE8Xeewo+Qm5OEqmb9x9WFmihSAew
hltDR0ibTOX4in4xF2NC204v88SgmGTaPxu8JOsuWEIIcJX3P1gcSzewjJJv0RmjEi9IT2r6V8eo
KCObDUh0Mce0oYfYOxUB5HgSASQP8yd+jOIyWjqehwQo22mFIyItrRu48ONH7U82TwOrPA6axiH2
FxuwAH9a1TI60miKZDuuhpaw1i9VK0DYeO0ERZKseG5dHRvkyca/+UwLpHXzUX3qmkTUNil4a0WB
0dgKzxAFPGBibHgsTHh9XDJI01+zNvFCOtqYN0XMATf+ERYcQ0ei+8QC1E0QzdlDjW9zUpbAEnAo
4o8fs/wHh6elLy3xpPQDrcCnRYdrvfIb3PhKXinZ4EB08DV07T1kt44oxGadtUmcRqNYAxxsXISR
WAdGJUI8BguDnvGZkMRymYbc5nPcGikpxHE6i5e1nPts1h6pkTzmKDkxCO7paal4Au0O/HmfTTN0
8in17KSfG+7sjieYv+/fLSuldquL4c1hijADBUXD09xQ9ebwFcrlpYDLTCSKOTKtq19gy4fqq+mi
WtuEA8LJhnEuRTjlQBweFsRg8A2QguiiLf711WOHO3WDv/XE5ncpG4Ki8oNIII12yLa5n0RfT+yQ
VLkuwl62EGJHPCjHMMq8K9ztebx7ejmbx0lnem+KDGmwdMMZnR57aADTAbM6NYW/mOn4Vjz3Ee6d
MNT+6/JLILw3fWlL14PlgeVMJrg1ngDW3zAH9ppl/gSrIIZ4X4R0odYXIxnMATHAYnocT6r4YoWz
yJsQv06tAPtQJ0cwvkkHf9UheUN530ZWhzuSHmYQ/a/GBvI68cMkXQnNv55hk1DDuaIvyo+Bf9Qg
2s/8+W0tcCtTcpRezaftFHKgd+GCPtU0A5rRzG9hrfAR8tLnFo32nM7bTmP0CZy0tA0za8djhhTh
5jQdnvw68Hm596wOLq9f9pAALFSvpukQCXEDozJqkaFb99Y3ge0qtrlo0H0adrBiUFttDH3wkXmP
mqyrCLACL1m1qjAXYysn0b0DbLV82c2oD9pZCGWxi1wQ+nLOmQ9VEIQx0TemAHRV/qqaVyOwzul7
6VSxKFB74v6/ACIzNnCpUeSKLZp7YjxwaPOA+oW2NATGTDDFnd+5xVersHXKeOi6yEPVEE1X8rVc
NLncQ7yALmlrXf3TDuF4yTZ4g3FT4wiQJ9GgtyPAv5Wery+IzTpwczkScJmziVXuFf0bKpGC9J5c
Eld+e9x3tQWAU1YmJ/375Y7q+v7fCmvZSTo3TnA3e5kN/yyZIsmRnghbcenNCkXgi3phHGnguHNz
xVQvWXa+2o7++LYwX9gsOk87oaYkSqYdibi16dLyh6t7kovSNpKt0lp7Pj3Na8SIBJEhSp4QCJuo
MsMc4OY5HT0xLu/fg5J0rO2m524cTzjYsJOj+eyXdO2tqn0Xag/QI1R6cIWw6pdBeoo8lrh//iSW
3ALmgMvbdr7WjWCvsNnPsf/f4zWZQYdDqnkqz+LK7wHb4KSa7zrIIH/Ba6fCDkCcPeYkupsPIZA3
ffXbxVNXvrLrQiQ4CgzsANfDJbhotwaMyju6gpVexIct8wp+bye6dwsUb9dfOmfu3Gslkg1fWBGQ
IFNl6MYyaCZ+RkV84ewgJ2cQvHxTIZxYratkKv7HvMjHzwX7MdsdhQ77tLnZLV84diq+mLaujaAA
bwyYawOj/s3PhYvou7FvUJbEitexbkfEn/Dnx/R+N3gRvalecaZL+7EoZin4ZnNDBrskBQtefV9r
4R/G1tiGI+htBcr4iqYY7VvdyId6YAqNtmee8vVmWEghq8McfgCz2f8luEziICSa9Eklc5H7Hb0Q
8khCJ1FuWNTFCQTOlyTmMHNgvOI/+XBHLwW1ko7za9/caIrpwDICmuag7EzE8CRljpEAJP2YU6NY
fEzU5JIhII7twWBtdHXJX7fJMhYNjKNgOTKS1UNTHcO4+AFxeM7zc4QrNVUgHtg9Ort7Wo/vwO4C
+D5o8a9c+fUa+kj7hANz9tAjI6IRLHJMTSBIz3debZ9WxNSQY3XVIm4QoakbkqEBHjudSkKF0x5R
TIBMBDKShBdlMBu20KJaLc98x042lGgwsr76MD7Q+Fp+i+k/nLmMQM9PhzV99JsV6U9lc/19erG8
JeEArnXhjeydmPPpAUSDgQvBVvSU4nAbn7Zhw5LNEqCRqFjWgV1VIQfIcjjO4ZuJ32Efz3zSWqet
8zb1ozV+yc6/HQyxS00cukV3TIZcW/t8/QjvMsvwJBWqzOIVCjx9DcPx8x6csTEaJYBwYii+n/fr
SwCiFqwKrGFoOMvi9CWezCdxnI7aBSdCHRIqtLZDXmyXsB4W/DHQUMz+CYKiFj2FUvUxR7CXcE5y
kj36V5Kvfna/0t/fUW0KeTkC+2ZyF/qXigGhMqE8H/sib9+Mha8sUi0cCIztLbGpEnDDHkh4W9Jy
VfswAWEXLgcgsQWcN23keCczMA5W/GIPArbLs2ryuO80ecI2GUvkwyP9mSGvj/foxDCy566+PSz3
Lvb6UKXv706BlMm1SZAkOlvjgIjqHWae5JmSDCHtrivDnwaBP6rVB3vt5VT8xsr+9a+39ufeXwMJ
iDoYUF5Wbs8/6qUA5KQpoZrHTWVjs6QQ8M8CQVj1aBKQecOO0pfFoHSmvF2eLLOHyzJB5nXxaz9o
jYwu8q4t3Tjzeg1RLL9r3zc0QM0RyloQg0FCo/3EGxwSwhEwNoZDDcnDusltjU8P/mrqFUSXqtTU
snIgIfQxVpMnKE2BWjghugaCW50ay80QIm1p95rLwN0vaLpRg0dHToD1UOcY8D0g//I+uSma+p/5
wG+ShKULdm7FEPAATdrtGhuEYtnsae3bNIQx5zXR1lxgjcBFb2WD8HQ76t1nXSwVhyQJqWwyKp60
S2P5vYlOKKUdrpD3fHwySvS4+PrmUKfd1yqWh3Mgb/kCo6RyeOf8F6nKienXedrH6QX/tTcwAb9D
7iHUDo9u9kt0ua/1JpzLwsK1+jDmgk2dSH5youJtBu/8h5MJFwWZMHkoDmoRdDOtYNAuJC5aMCDS
lAQu9+jF9myKbDHJwCnOuiTL0yIieRJwckOoTYlgfUW6tbO8ZxnAEnLC4BAgHIul3Q5s0HaM2DxD
lLSL2D+gOvcE8/sWg/edOYZ+0wmkZ6hh2kaDv6V/JqfLk1WQhLZqIk5c5mvEpofHO4+WF0PIa2VG
Ea3f2X+TewF2dZd29wCyTDvesbDKWSDqH4ZavSKyGVlrfUqc4RSMrNm9UjGZ0ZhI0zI7GU6A5UUA
Uxu4Va734jV2X4e3Yo7N1r00nBD8ChNMkv6NBwwz/x4qDbuUBOIhjQ+mbkTplX+6DjzBKL5aPOtL
IfZyun/iWB2OMlS7m7nyosWrRi2Q/K+MgzGJkHx08vug0UGj1CucSCps72C/Hit1aM/Ti+Oc0Q3K
e19i5Y48u9IXlUIIMk3H96EH9/kLf6evYdryseR2RtwtOA6gUgKqOofUETyLA0g5KyyM2qWwPQFz
6qUrgsReOYO/x8GMc+w+pgV2M1e2Eb2Sdu0QpLiVrFHJ63tOZFXP4Zi2CO4dSUv8q27iq8XKgTCn
eWMET4HTMzxoygkvhn1sTEzqrrUrPE6x++cgrWWG0ctRpE6gjjqOdAEk+g4nX3oKGkL1xtPGKTiy
eTBlXhU0a3CYXAJlR/KkQI1ITIOIQ1UaShySpXh6R5mX9S3JsAKdwiYp4VOqoI9QoUxg16NkRAgq
l5EP0JRRm9XvZzzY2MI4xWpSMGP2ESTaAWHSvCwqfgogh38Z4wQ+Crv85sZ5UBwMQqE+ph2FLWfH
p5M1Uf6U9G683en74ymG6vxrQ6w2EReIEcUcw2GGGB7F+VeAza0+J0L3jQLwGQDwaQPM3evHJAfC
91OPWMuE4Zzy2M+RYWcR17t3hYq9KJvUvZnnI0MZLF9jyFD0b0Lg+q/8CmAJDkajaipLOEtgvP9k
fynI/BmlPhWu1j/vHxSEEL6iw2t+JoqyNA9/TEY+b26bfyymjOlbqFchIuiZzZnwuD3vEvYFOr6x
mu0+XKc84nq6kqiLb799k9er+H95DM7PH+4+Y1Sb/xoP7rQQnAsr2x/ZKSDilOLNKFhhXWoxmljJ
HDHnTCH0+F3KWJ7mnqBDMORum1PLw1BOxmcD3cxvk0pWAi/UhiuXl7maSYV1VH03wV2STDfiLG9Y
gAPxIgqDfgZ6mgqhqEwLDdvjneF7XLTrDorkI1B4I7OO61aQYU67L+eGMX5bHTPTUDj2yPCi59uE
mMTzrG5W39Qn91+lK9h891K0vX4xTAggNgy6h1uxOOD1luq4zhNyyZ2bFY9LJKHhRAJZdHsXFZvn
+mRqWvyD+I8538WuBcXw+/bChmHOCcDmvw4bGAXKljVjt+9e9S9AaMKOjZihJ+2WgAbKJoiwK5wM
P0M3n09FrtkCTcEfRD+G2baAi9HkAwEPDNOCpyno5a1MmOPh/dpB6SACbDBvl10Upd3/kPE27+7M
hQxWEX2U40MABTRrkTe1bQ8iXRegVKpeNWrpP/2w7fvs/0bPn9c5GvosCwiqzOiXte/8Pkuje4ds
Jd04mXY8RyIQyRNctEtN8Ch4LvFCjLovJ6CjhPf2QViLcpv1MVGIKpKokGtzyc3S12m3Ummlj6A9
UrHxOmkoNUuS7BN+C4FkXG7a00TWHRmgtaosOO7Yk7hdvybMqDpGMKQTPqwePaTCNwxB15lIynvz
9u29xfiukJ3L3Fn8XVVkqoMBzY2UZGF+67lcmFZbe8h93fA9daAiDYKXkR+L3qr7jSayydmMzyC6
7O+jkBjMHD4va23ahtdPy4w73eaH6R4QQfMpa0WtrSnbSUPVjH7GcGWkv6Vv7UUOzydqkS2Ma/7Y
7TUP0iz4/Z+aalhPOdrKUJzId40IuCHjS/9b/9bFktcMjdV4Q4c9FTGdYoJhIuMGKZ/6+nZ8PmPV
bKLN6+Yq6igg+8PKphxxWu36HzEy9+zBwhEwlwlsWgSSPPWlWrNZIWrH6zsOpMBj/HgCDHuQLjtB
Y6+2caPdrOP07WUEn/b/qLMc1nyqDmI+BfBRlYZyGqEQYjh1awkz6NdJtHPmA17GgXPypQ1Uc+p0
mrN19atfbh1nTdmvUtYmW4RbHXO1T3ZI1mRHPyusQDv1RbXjDCWwpRRFFpguUyXW2Oq2+6jg0lQO
GE5FA6Rmr8ZFMff4a//0Xokyh8SU9yTwtEwRZvazvJQTSbe+68sP3Qwuok4sbWb9s0iEOSDM+f9/
PI4HPT23mCXy2qlgccQUn39MMlbeGrqt4uLNpm51sky1FGC1y+R+3nuTT4Aw9xGMkiDqoPj+ge+W
UBlPiNh6rXwGfNNDVaVVKKVp8hRVUuYiuiT0E74IgwBqjB8lKzxP/dUjCVJSQBEAy0DH5w1KDPuW
SW0+14VrlwNsfMLhYq8yMoCeSc8r97zRBo50IRG7XxL2xVPOxBlLBJtqPD006BSsP9l6ah8GRX27
4l7l/rdDNyQZw20n1ly+nuB0DWMIF0dCuzMK96YkprYYLmw6TJbKCfYUdI0qXCAbaZ/3pu7Qym7W
o6MMPLlwvt7kGb0Uiwky/NnVcJok/XWpMWazhKpERvdv9CYewGwJPpb6CksCHtJSG523iP8CkILX
UIxOebROSjOS4WTYZi/D/Mfx4ts9lUb3GmiRHbvWzw4Lz/QFpSqOMJ/8xrvy6PHUPWX2T4eMx2jC
B1bgrNB2I+eulJkp7PpvXGnEVctkJxi9xDcoUvlsfklgoZHNcOjheYykagVTeWcNykGk/vDOewfj
VbU4H41+EpWfkCXfyd6weVwojVT13XxN/MW09QCkDbfNteAkMiiKmbevUAad0ji2XLt6qPPd4LrI
D+fulZ6lvXyBb6s4euK1gt1RavKIQRq3vDQJ1QsAfhLwN+jiBTH49E3v8eALcgCCD4qjfSmTnZCE
jzwooKK3s8OH8XVYBiRQjXCDyT6hCLiTGZaz4uvDxX33HC08hsDRfqwzvLgTOK7xGdHDNbfNI0kK
VEQjcFxIGAS3SPEbzf8pY8By9VqgSApdG5M3a1y57SCh93vKC+L9GGGNPzdd2R4hV/C4Z/w4n+gY
9/tWapR0mkq01BpiznvAcrHKTDB2fbZRfpp9edQg/gq0p2lOXgqrDJsCXOcjqf9MrEm+J2dcEnia
Uesr4NSPIEtk6IFAlg++EpxHUgPKJz6GH6h5NtkdSNdFw1gqzf8HOFpGC5iO/DckBbw84ssuq07n
48ctzovCipzmFfU4u63QCkU2JVuEBjGT2lzg2ZI7TI2Lu1GM1GW5QKorZF2rJ6XAX7utn3rD1MkW
ArUnFl97QHc//uHUNLg2fB2TRYXT+9ld+pmBgJXZ9jBuO0XoKX/8y3BaPYjXElPhGYi1w+clUfrS
kjEfkKj16v1xfHvhOKoQAcghVUD/DwdF7VMxLxJYVSQgiUJb1eS6QoaOVh1kDBcYnikd8F5JO/nY
rpLVVAvalfEVNszo82JR1iVcMaZ900peYC/DwyJtEtn1HlOwBvCMs1beFUzb0duOFeptnHPr5voY
pNAWWjL8jXqaU5W7p6hD3/p4cLskJ1R8+mF9Dv5sm9wbbDkHe7OeLW0yHcHU340Cy9r15q1Uwgw4
rsWb5Ubc9eG6DfV2feyz9W8BOtYJUOR16pNS/zzJ1bjln+B8NWAtXn8LNg6PkflX8gbIMfQmH+RR
8+v8EabXyGb+6h7H299VUCE17hbasUdMAyw+tywjZLI9GwKoFgJ4yZJIkGFK73nHTQmVdPRpPFBO
UzBEypBdgFuCnsHAenpS5GKnbOUXlp9SNqZe1oKQFhhen4WvjFLf2hiSkBSVQ/WTtqjXG9eIBbLI
vNdxeHF6dSio5mKh8bBCcJPNeno1oSjg9qlCkOZWOzEIJMFFh8ZOqZyBD/6buPi9o4cRc0bPpPe/
Jbyv2ppHX0tHffDHTUeQkYFru6rhrsH/7OkWYpmlLE4YWDrhE6D0wzybMFLkBN8w/cuiZLOzJbIA
MqgxgQvNOMNIeomFIbQkd1KtTU10EBAvh8L6RLd3GFZ1KwWbnRnYEsr0yPBqESpVsd/NOf1eieVk
UhlwtZxgnBIF5u59ZZL1f6dQPtws8pkjQQo5//xRK9vDiSqSbf3aDidDhz9tKuwbRqXUXWMzTfDG
uw32R9czq/xtS6of+Mq26En+rbRz4XVXGhh0P3A0QmBVqh09Eq+wqD40D+QnmUhp5RvKSQBUwu/L
axqKASKn1UZTJvvVoCxVI+CaxfV7mNjsK23ti5xIONXLizTRX57Nf22GCBBL761JVuXGbPBDhdRk
mrts
`protect end_protected

