

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
b5iEwcuh/jbBlgyw+948d3lvWBbFsOTNVYtA4pJb/+7lAHor6DKhd4akfRWg+MPGWaTgwtrV3Hjr
bBdLdBNTBw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
VtyA/tLK0cCJJRwkcmojHVnJYFSH/hY10K0O1xHrVFcESK6dXqpZL9jghTqU0K8Rgfgyj2mbpSmS
d3OjaMJOT/0rjwEIwUBTQhpYCQbUdyb5e+tsu6Jle32rY2EO1nN6daySTSkOW0tup2zZBsIOCr3t
+ejm/NK+miEBBu1xCLg=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Sf+0xczGTqZZx6dcqp2GTylMp6ojNl/Es91rC3p2Qk7Z8FK5U8FSMHtByvmeihj5pitp5aOxAIcO
cjVP1mZpqkA9QTc6UkTBmHGnHSpwqkUrzOtsT2ws44zFj3ryr3hssigeWwtnVK13YgLrM+5chsUj
26gA0jBZIt1YnLsbFPdAg3CFuuIkHWQ39NEQDeG2BTbW5KtUVyDTnpctdLn+1GQ9lYJeC7lVtfwI
4B4xEL5dhZYik7uaLaobO+7jlipeHv29o8EQsg6BnOj1c1kxrXtTLsKozU5mRUSyPYYAw5cgAAvI
P9ELz58Fq2bFhjjPjC0ULrxEE7cl3R3lE+lEcg==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Qzj1t+dWRPGHMv8nVaAMZRu2BQPWmF3UL/i0LvBgsHGjHy3fNoKTLAs04wnbPCVtn8n3ytCSqZ9j
YDEGkJeQd/ctkBALil+9bfKGzVPGZiyWs36ilhf0nuaehXbM+Zt3Nfkh/wd1LKqVrJhOB/A/iGYL
jRkozXf4ccRU53dhQZE=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
eo3jj49OyneaHUaTvAS2/lR4/3L9GHwLzRAoxweYog0SBxlqFd2rrO0OlKoc3GfXgogda87o4tmz
l/UHxih0uJyK1snlhQ6A1EHKpMBpfD++gCN+S5IJFV1QgpWejKXt+0a0zp/A429l2cS7KMD2pUZc
B0C4VRE2SAMGJhfx1GIRczPJREH6ZIkDU1qmMs04rSp0PaGn6eV7+euaxeQcoqowg8QlRFnxfvHh
5JrqhxNCP2z579eEXYXH3AWOzWM/EnKEFUTbEaxMGP4W7RzgRCZvuM41apmXDWTVjEj3gQq6xKn9
0OWO8TXN0ID1dcJmFJe2x6yA91duGkuqWQQaEA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 43760)
`protect data_block
4ACaOJDuC57T9QStEEELQYSbMDMrFuMGkeqKnKLf90nGPfMqXa92PfGXFZ1pxrArXfLYWCDbEcz6
9AjYH8isylctD7s/CVqLUb5FsEyvd9jnHFinQSRS2s1N01iEZA4KDo9+ORHT3ZJkAFeoOPtufzXk
JPKAWkLcLmECf8FrXvYl2rb3OFBoaivm21UX/GzNZeY/hSexJjmMF64RdgH1LgUvBQ3RdyHiVwpk
tBSJ4l1l/uPHQwSGhVxvrAcjuICwC+R+7yLJvQnVfsoTyeIcTziHbVJZcTw/2lV1NQ1WrWWuDcXd
TWaykUINYtTAqOZALbq+i01jiZlSkE1zkpGLuHWMNd0Cy8uiIBljbwfKSPD0BYCfkPx0JI/W+fK0
yCfCXbeJk2vvehq7C1LW6T9dd8VO7kO4u2uNxInZHTPTMF627d7u0ORb9NmxR93vPG+7HMAwy1R/
ucN6KLZA+JaSxdbtTMvK98pZ4Acka2lKRoLln5ZjWttpICyYCplBA91nih4JYdjpPUC/Ec534TwH
Bu2bDo5GBPUInkYqsthveVzOuswLYBdiV9YLHhS1WHOU8/9APglb6lDIHRjt7QMxIS9oVH9kSIDZ
VmfON+nnfwuD+kJW+xigYNHT+r6/AyF5/u8VdtZod6bKNSJctttMDoK1xH3zglvM2vjWUurBP5Fj
qO9WvkgKhTnz7NqFUd08lt/mDgSu36hgE4Yu6fTima+PKIQSrjX9lo4I2mYip4aGpjHE6btxeKP+
sCE8Y3U+/eTxa13+fWE/nTZq72/jcc2D2SezPJfSO5zjJ8zN1/C383uS5zKxgTp/fzzGv2saTojx
vyxSG2oo4mlecTH+Y3nQulcU8p+svgwlREJSU6385F3J9A9CSWQuqN/nOf4r6/OIvM5tCm38fo2W
hGa1mPSthgQrHbjb6pcegPEB5AY5fljQBGv6YrwQORFaiFMEGgFR+b3g7mOpoz030fpWGtXaTfrF
cvcVY1eIryXJW8/epbQiHfmfMK/2eixUdzDXlYN0KFvdwdYlREjran7Ms1bvGsXmAPU/V/t7yBwm
q2pOCr+Xxkb6+NcaGPE8NsvpwprOfj4Ff4XfXLLXGPwDZHYzmtE1R/tTBsKzSxJOpJD+bfA9vkGV
MXszSkDFxdTukO1UNhc4oFdTQCxQsmVjncYusFW4nZHpRLf8TEYUtwH+IY9WQmHMR+STkM4m5CLT
GiFIkxgEYTxxrYbhJIJH7T7NqCbh8aLewY6mUBvjejL+d0mD+sccXpQwsqi5vHD+8RCemhhWqbrD
km6O9/kQp55+4KPtnT3BB3P2G1vf31FnwNc5WJOKFy+6PoyzhR5cTjKPoGoOccAWhUp2DaaXEEL3
/1cwuxRcNIDhWpz9EAlwmmnN9vBsD/np9ztDTCanQGTbNdgBKZCzN9xF42wYK1396MtmKTRUqrJz
sGip2MW9UsiVWyNHkHKHxweaImuG9wxDcJ830eGaTtzBIkYq+eQ6PAtPj3mNxrHk78bHDIA4Zxts
O65mImtoVGMOLX0a3b34ZMZBEi0NwJ9//mYqQRKlzRaXNJyWfVMsVuD5Rd1Fy96dIw1OuFCIcjOl
x+agfFbOBdZsC3gvYVveCqa5vQ3fTwSL9OvkhqQvcmbuFicTlPiSYuExoZJkgXM7aak/ydecT8AT
Sy2qPbjy3lfHhPdnO8VKCkdS6GpmpX4ZqeMkCxqMmzZwYlvdK6TY3Lut0cC2UG1dPCSBaiXp/26+
Okzcxrd7ar7T7ixCM2fIngCAkC+RSljSgaBw4T7Et/ssTrEpshwMCRqUC7y64iWJfIoyMVlhzWTM
4UnG8e446/TEP9a3TrjseNaQ82/tGBQDXXZqw8eN+pB0lGBV2HTNciEvSuUOFdjP1jRfMsWbMeuQ
T3lKPPesIwqV28RNiu1t2Y018JPIQQstyx1G0UEXXNXdUiERhwQTFOHOikEk/L0KymSXngEJV8qt
1QN8qDZgS+jD5YvjokuBuiILNK92ZSqPL35t4a1jdCLW8wxrGGDDUC2HMkdtK7xj+bIeJ6FbFxxs
bImG+XC1kh9xiSQQX/HQYQjYW6H8Hht3+Ml2uRm2YIy/jpqSR1bLkn92tNrKHg9g5HOO2+EGTRLV
7rVqRadOfIur3nsZH2sFMcs8IkzH/ORLa6sA3F3zrF1W7xRVs/y+sXog1vyC0igLwP4mN5vh1cdX
wAt5mVn6g4KH87fiMecSNlFduvtEJe1XrFJBvJF81W5K7e0apR+pQQ6qA4WLQa1YixYi5w1ko+Wh
ipj3kWVqOG7L0hF5+fVqtrlUBRCec77pEzZzeOZwQCLBLy/e8LIr3PViIoZqM1D4v0d0sJe7Nale
A4Ynj9nmmcgp0ui0nnAo5BfajFEWg/2/+eFJZglq7LVP3upZRGOzOwJSAdf4Xht0YbmopSwSktEC
jwJ5Mr8zkYyK55imMSpQGZ8J4AEWOgxFpsW1r1bDVmupG8A7kDtwebOrKfDN/BQ7yXbhplreSCD0
wo3mJNtA9pVOaeX8pGkOnk74SbJAK9a2lxjinLdV3WY0v933zqo9+JE/YUAwISACzHjuRBnvXnYV
EzzHyk/uAuxN5wMz2ip2ewd/U+novjhsugckswld/YiJv2VsSmu8/wcJcEL1YtAhtjb+j0stTSgO
HRxb5109ee5qR5Tv5POQrO3WVCZlVdb2yDC7CBJ3SgJpg6Szr//MobkCxQXpV2buz9DmfjpyXqdB
/HgIlUUHlPDJxm3hr5u/QDXPF1+iaIfp6YM1fSzG3w3WMYm+iGhFoVN6DoTfnLadgk0xUPNmTfUA
jLxKZVlEgDAkLwoyhxH1SH1ETMZh7WkNU4q1hdntuhtffM/d6pTDArlPEjvZSKX4qzl2XMrRYcWQ
ebD0ZODXv5IEBHLXb+iOvS+cEMv9T9OzHP32w3CBiZw3jNBnJhEbFEIENjG/WaFLTz1qFnlQzUhT
Mry4T3U0DOm1VuKUTK56U0/FMRfS0d0qC2q1nJj/k3pE/xBz8L514KTd5OxdL0j5wQFFClGBhzWS
pe/RMsjG7z2eaW/P5GrWKw4xmGWeQIkU0flCF7kHzA9zA/NwkCpRMPNu6rNz1cuRXSz2b4dzjegN
yOW27J8aMOMqdSYM4/aAQiyd9gjP0E1Z3j2VfhljfwaMT2FrcPiiVHwouwCOUqrlOdFO08Dg+KjL
2RyYvQJrT5h5lULKfm9jyaINglZn0F2QdGMa2i/yE5qcxZ/7PSpJNctGIiDpijNQGwV4NomL2hy5
MN+n4q4kVoRY+kg0vbphrmg19Xwxmmj242dzSxMBlSnv3cWdJYOxdH7P0XBoZCr9DobRPK2YneEC
1BcaGVui7jWHPrGZqP/FOOqyFyUMzxzGndTKcWCGY8yQEDS/WUcyy58gWe/9pwMM4YySBeHCpYz/
GntJGV2S1hVpy9+G0wfNDLSjXSMIQZirgLS3OBYwD3t+cAWM0z4BZ44T+F+uyUqyP22659bAewkZ
k7XJWeS3IFK/9R5xRdhZvVPrDKLxrKu1ivNzHevvdKrvspiFzY45xyBis7kj4typyqEJqVrGBrgF
74XVIjZfok2WNcTRjc6cuxF8z9/5+3JteDYgifTW9d0iB2cGPb6QlL3Z24APXoI7bPUH4o6oJbfi
K7LLKu/gYKfZizwq0KGXk+vtOJPLaAf7cxJn+2bnwCbPgFrPfjQu9uJN5tg0RFH2mxKJIilmSoRB
aju60bZgzXCwxZF+dPAut+m9N901s353QU3uRu0LSbb5+mGwyBwnr5XBykf1+oNrCnEcwUgcvz6d
Nyg3IkWlSyNd7zDScPB89gt1wkz6Qo8c9Hh7XGEAcpXd3ZZ2sT3a0MxUCExX9VYpKl5I1NxXQ1FA
WEnr4vA4X+Kt2MMEgr3eQPaNxy45Ir6mxq7tTVOIPCtr0IZXCO5t1bV1bsb8FB6hOfXi/WZheJie
KuxGW0eZgMJo+VD4st1az7IVjTl7FMWdzFDtADKl/SAHjOUCHSq89nnF9bGnRSOI1xztnEXVvkFA
Gne5XfUXMTHyTznZABvVM5PQQtBlX7TZkH8FBboVPydYqZMXCrIYAAxpqlNcTFzNSs4PtU7FtkWr
yeRS8TRpkhRJTA8vGesOwdTk1SvqyizcfLjhxDpL+mc8t5hygv2p4iEuJYhEvpndeEWSzAUUPvMV
nl1hHp7nnDDrO/N4c9vkNcepc32SC0EU0Bu23J6ilHr6T900AUUR7lpX31RkUrflgjiayPfqE6Hx
Bl6QR+qhA2LzgO+lK+VDXOz7xUscQ5wjVmOXH/4OHGTv/YyarPBx8N7qn/JR24CDKo+13TcBXZ3v
+BBqijCRs8AIA+LC84lSw2ambQS4A6Q7xVX6h41s80dqUHiBJqqJCNd+qjTuZg6M81VXHaJUXG0L
s5u7h1E6XqfyRIVaesW02RpL6gICPTpoD1mIcyE+TeubM5V143Na8X6OwFKKQv8FOnD5P7actKP0
2+LNrwWSXD1ZtR9QDvRFhmv3VmygkIgXKoC47YMigKFlroJ7P7PVMPD7u+6kb6DY/3nSZeEWRBua
SFAgGf3ElsCu9Cr69Hca2B9K/JZG8lHwQNYuORZWzi223A5qaK0nYqiYUoK8NmQwpbih/MtsMykc
UOQnlNj/rZF/juHUx32GQT+UTup36jtwvtDnBJPmVv2LR6VTmADP108qLf3U1GwxDTxWCjFrMCn8
JbaU+BLjbpmiz7xx2ACTk3kpZYBD0t/VgvYiTGUf3Xssv+rkga8qGBUpLwn2u0iXpUiGWiUZljJb
1mxMhLTxL7hdAN08DeTC3jmdwyaWRD2K3drIYHKyy3SkVo/0O2lMYQIGioYVE7Va68ajyP2IGgGU
8qNtMed5C437/kbbfGXegKxGHcIt/fWrc7oX3Ipn+o8K0g8EFcUx0Sm3eqlVnWgT3FUCPVJyvTAC
eBR7YxQSn+adxy6fi3ERC6k/Z2zj41jpLb/PDvHOc8GvgT6Xy+hupyNnV3YV3Z+wj6yw9SZjrAv/
FngIYYAr6+H3OtDj2AKR2KxEByxUpt6p/TyEEvuufymtP1uR15SsqkufkwLqu4h1iMVdnh8u8IH7
lwoBTuF9ZiJ4b+nL/ajBc7WIax4AvLCzu/9RShY8TTp/rp9iznGd9EIr2qvx/hjc8HuqeEfHwb5n
qD1iU5caEJ74tEUYyyE3nBKymNMjhI+3nV9a/zDtc+A2+2dQaZjtSsrpEABBvPM1+JPJ9qRlRMJw
t8YV8d0OONfZJ4Ri0Q1cySKxF7j+kvBPTYLj4XrDmIeDw+2B/taB3GFnTarxqyElNkpzszysva0L
KM5wMKur89YAOwNhmNbHY+GrrgLKp1eJ1e1yrdgJvBrpkIAUwkmxlvXSFXAGTGNjtFE6Qppze0OM
Q4T5n1OHWcnRWnqKtZxRZF3Fn+aTrwbhwQrmMFzjUb3uoWDUsTMuWft31+Np4tLds7mqCwN+Om6J
juKwjDUgakWAAkaV9t9V/qXDyCDn5WJ2g+Mridi6deOgWFjRqW+l92DJE4qdSuh+ZScoqAc1En+y
SjwCgVrrPFf9HZdgYpS6Bn6b0ipDJMqRUkwUD4wCi3ouNdTr0gk3mcZl2cpHBlteUfsIvqZ/snU0
egkeQz1DRWC7197OGi56LAY1ezfwUsVxnLPBdbpOZ/gQj3swKePnhEJxCYCNVIF2EHw1OP8gHnle
asgxo1SXH3+wlPLarOAxZt6ZIxm6HdEYgu+4bcc8VhfozSB64u6a+sFv9E4hV0ExmKLIl19vQFHU
dl1vnoEZyrJKNcxyDU/o48UKuOg5LMu52/+CmSetqWD/l+fXpkfo3se+p5qFJwHqcJlkNLdzSGMn
pf/v40xoW3GqqrsR7M1EzNByBKmA6XpJeJn64pgilcFJA659dnMzJwncm9BvvZG85boj68H8HXp8
s9SWsFhE6brtYyt4Zd/I+2t4UJOXrYb2b6DgYnt5NWymAbPjio2S2pNOmP9227QeHIZJPVtKWUoB
+FafKrJIhieSzdK1jSv40e0X+Du24J2UeDJoZfri5ImA1xeCdQ0qxGHRomNl5mFlbxfE8kyPd6qg
iSReIm+unmaSwKoX5EVr68TpLG5ds2x1rNp5e8gO9d+4Nb543HLMzsCzFrxHjIVKgF6KL/hJ4WN1
7959CSefg/WjpqBlTurf/QjGKj055W1gl0u4fX+N9LBp7I20pIQMBnjApxkUoMdDTpPA70dF/sW1
kWXqnWIvSliv29yh/MuuNOhzOWshdGKM2b3ADf9ZaGZdmUQlsH6RxKrqPJNZbJdoA+1K5CdgdcWs
MAP7u99fraPPpJ9mlSUmIU3F8vdVIBoM7IsStgcbKdGqfuy9DnfnxtKGZCdhkZLxYtBEcax5jibt
4yATxrByT71CQY8Q8JkoPn1oqmju4d58zCa3sTZatwZvcN0UleNZSFVakx7LpZGq6qBOvGIBBDt8
XF5u2x9qKwXPxJfdldalDcRTtP/3qe34sgVLUD9HonAn5NP2xfmK4dJ/tSGyONpB5sm9X07N1CEG
uCpudxf78wRwPyr2xznxqrzLLvZVtIYvOVF5HBnPrCZjo5+FzHlxTB+Asv4ZvV4uVFPRn0dLoi3A
pJmD9SXsm8pwr9okG3h3dx3Ke/OuviYyyH9fldAf6RaSR7NCAdXDM7dTGdOvC+XY2RhzQyEGnrSN
WTkyCWyE7lgX4jnFwVyHPvDVyf0yGLSa2RFfMR6Kk8+nsnK73+0v2tQ4i5ty7UPPsv3E+QgWpfZC
67NM/hmdGkslU/hOaYt+xKzyrKbPvisGJKbPxIS2Gw5OrtWOZwhoWXHkliKOEEDOG2rqPIzHvEg7
g+8f+yMuybn128uKYHymNwvsfIk46YsIYuGBzyVLp47OdliUe+fGeSaOW8o8MLKZJyqD29L4Rw0m
Z3fZazZUzw8irXA0kLiiFbXc1JpcyIl7GsE2xQtjhKKLiuQZvEnijJ5spbrwNOJAQbF1Li6fvNg9
u249nYaRwjr4wy6TXrquLMdIOD++CjDW840m5+CBoJky8vXuBat/PHYVX91KqwjNuWQDYi9l94Md
FXHLT/MBrirweEpv6FTKa61LkYq4GCieolX7lm1p90fdyO8/Qv7J4DFERTexCfq//5t/K71fn1bX
pcYTsEPWOS4dF6ZZBA2zM+wEPLOQBbXkUZIufjKPy4ATdvGEMFXxoxMhSEkkFPDvpkygnw3XLuCY
5jBZC6ZvW0LccOf0pwgIzck5FJrvIjKG9VF5CEB/htfbk4k8w98gfUHymQUbXrO7bN8htlODyFZ6
Y1vyTxTDtMaY85h2H1iu5huNmKNLgRGfLAdCSufatH8IiRbJakFbdPz6D32EVA0jP1RR2dpyZUns
4flBT6A5rrEjNOosmsBXwMgD/BLe2MThyqSVmzBllqwhRyGP9Hgvo+z3jYnJ9/ltWEeCZRN5nbsu
Q3GWuiRdcxEto7dW0KR6BckaSQpeUc+yrd6XGIX+IAw7tM8ryjmtilrbvUSsh2MkQ0qs6/XFJ5KU
yZAgPk/TRfdL5Xs5eOAPjuNCvudup9vncYnhI81N2wZocJgbmTAuprF8WHTnH6BjZBDoOuViLVLk
z1byfMyTbG7SEGvhK5c7wIJkrIfDisq/UQARuv+pE40vDLJiK8z5Z+6hiHEogTQzC4M2QWHoQxTv
/4C+d9zSc/2X0Sm+BpC3n3QtMUlN5yNlSxSYRCDgvuSVlxrAoXqxkERwrqWQyX42Upt7Mk36Qnpi
s5Vy6ZPrVUDZlyJilPuw/itzvbT6P0PFQANezB7REWp593HTPzhOXWqXZ0jzZh0SeqGgS6eH4TQ0
GrSYJkE8LbrKs/MvVhkv6MrZqLTasGAZnq2abzcokYcP+ZiZ0e8SDXpCgdJn2a16VjBjjPb2llzi
+LegAya+kufk7yLUhHN4yYvdcdRhpygtxlJvM+ljvE4/Olgq42ODKWSBI9LEEECbp2LKj075efAu
3+WPtAjjoU6uPqhhjQvE2LfXGquKJANLdjQVKSddWRkGDfunE2rofjoq+NI+x3RaHidpN2IXfLVs
lmsUmnfxoaNYkZVo8te4DT5ZzbO42XDzKrwLlO+iwbrovRcXJAR5Zty8XS0hHGqL+Ix5LWMl7ZfE
cG49u4mU2An9OkQOjr+fqTVs6mHCdoDirYaopEHTNkpkR/Xz2o2bYoIDfYNdHtInMIvgjO6/HZ6M
fsIBnPXFD+7Zq8tmowKVUV/5T+4TqzPnVP0Iuil3+QicvEd34E27WntI6YqehUb5LO81gZONr6cT
IAy/bo4lTTmZxBITPJdFre7VdE1vIF8/wccJrotiIcVBw1xM8ZiTkaxiKbV5FCIhS0GEcPr+PWTP
Dk0+ZT+6stLcZFw0qmyl3sciNBBzpp/sjeza9zt9PXHvBOuLfAsmzRNH+iLsp8R4sOF9uTkYpzMj
bgL8x6d14kOK8SLf/EJbnxa2kSOz474kmN0j+CFkTIAaQ5HC2+BVPUgJP4ddm39ks1unaOuTUEWt
nwxGSFGGlqjYpwtgfGz2MidQTcCYYEkcchCLohRU4InvCjHCUfKqqHUwj/C/A4yr6VpriZVcIW2U
F6le8RM4m2H48oV38zljnQXwwRb3hha9t4gAuFPrdyCw+VgKUfuZlRNKSzxJwAhvYm0hi0FUkQnS
SX+kkJaDl5W36mSiiBGKSABl9JfudYM37n5UjmftpQ9W2DqLts6L3iOghRczBpD3J+tAfN4Gcc77
Jj3H33tfntBkHvNbGLCeIhtrR5kSzgPvFeo3CzQU/a4x2V/yjiFYpomhzW12OuPbP1xBYvn5nbJv
NxmQsGZ83lQ1rCF/ooaAnn0OsKUGzeD6lXl8escT3GFX0t66pwWctH7e/pnvGqtIPAxvxob5rcEh
d50y56Z6vePuBJ8YOVLaUdpWoiWVQUCwc78uO/2nbzCd/RKVFNb5+8XrJ2yvr/vApDlaEmlcaHW7
tkJeTF9NkdJtqfboaLWHhfnkEi4E0k6j0qDSv7yfkCkJrGsYOXtYU73Zl9wgwTNaNKvkWZSpjqqS
Y+ajNVttqdZ/VMfSX6GHKbVqOfGNLstOgkNzXAqTB+q4j7nG0h6183Yp9ggCbwP60om7Xe2cbKcK
T5aSwvLJfYWuwGxwsKlx7mOSZwDdiFZIvKVx6ugBeMpOdgJHMHWPUkiknCqojYmsbOsNpjLA8trj
OJ/DnZKkxafT3bkZVkhQfL8xQFpulWsbcqBNHC+W6iB5IiYuXeDEBxq3ROFQbnreDL2qa8rxA6CB
VuwDZj4UxpSSJ5Hp+6oMWndCv5cXPESIkANu7crPW0Yqzr5vQ7Kp0j4JXXkQ8n5TRJdy618uppdq
E6OpaJR4Yvy6P8Y9nFwyNzXTVj6SLRXeXgC91HJy+Z2yKdh5c3VdAxCJnq+hIX7q+S0irNJh+DOd
SXa56jACDtNQzJMwe88uPF6dH0LT1fqPhxZX4EJjYoYGdeEr6Qa9xd66QXvRkLS8yLIu+yzq3FXx
k2QiNkvy8GTGdPnGzxgmOhxZ/zelvyGaoEHKuP9xwhQCVyNFSPS8nqMxPNcR0pRNEYxWJMb27fli
R1x1T0nQMJnNsBBd4+dtU5GxN+sBRWjaCB7XxiaTxfeKHTxloJY1vFIzwliXjr0KktXHs/3XE6oh
zXpZhFSJ4e/Dij4Qqm4hH7CTGMHGMGXIpY2UlV8JIr7w8J7uwrOGYRPyfu6NIdbJHXyPH3ckMo9Z
kFlvuNA2wmxdDoI/88/9wYE+QUWnUwkN9co7+Tcsat5HDd4dAwjfeA9fHhy5lZ3aXDM8Wv2DB03a
71kV2KkyCrQMSbFV2PaJablFVq1CwTXrdqnR1Y/0oeUCXFw26/YZn8tiA61VWRDnoWNHV9Mi4pPG
EDv4cwKhrG4U9HFJojk0mK5UiMSJoybNljXGIp+gbM09+O9dkJAvQ84wSa9/YpICAWSPHZlUB1+m
zb+Q9YXCnCmOHICxrLR+KAvRF57A9g8BrDMbJbHM3Qpxc5UtNVs7A36/ugNo41yn24oH9KX7WJg4
1PcBgcz29hfbTfUFz+QeoBalbSIz43roaPgKzJvjGEXsXOYv7g0ljFOfnXtl9T7DeyBt6CRF6rfF
pUba8S0E7GhjhKbddJSPsVWSHF6mr6/CPB7LjWuVPvYAGtFu9xPt8WHEV+8w3uk4DbBVDqeb7dap
xmtg27tfMA7n8L/X0NHtROafzQi9/0ZdKLV4y7fnEngL5g4549KjeItMCxwbv2cMlpS3bV3gHctw
F5UufhtwJM1YkovHpbNWAohw3Ikn63Hbb7teezAfxQnwCgD1KWTbH/PMDEX8vWUuh5kPJyEpkmEt
uus2EuW/aPf/84CKMcwuCEPQUSWYFVvo6ZCc3Xf+lKBwYfErPKP3eC573Ig+Iz/c5URw6p+Km4wF
4UZwap2h9Ooq9UIxrR0FRLVaqpYvHJ/GXoBQxv9fk//wyopwrlykf8W77pcax2UFXZP6HMYQbmJZ
l4goV450EGWtzx4j4oy/VMr6JOfkdfaF3VoAQM6lY7S1UWJ0rOI2FR9bnTlQCveUf9T+UOaeKiel
nr3d6g5t6O7sLhM+h2HsXbP/OC74sF0C1ByRRDKPJV/oXcqnDCGgZggscoeXM6dEgcD9h/vtnyPf
9XWZTjnb3vFc2I5eQrc9w+4KTyPQX19hVz104UP9Aiha/hJrCbaP3r7alWJ53cEdX+bVKmOTqQOR
eKKCCgcDU/kT9AKgoVfgcbS9QVft3oJ61t9NpZ1THOAZ1MKSNM8m7WV22gOYEAqlrrfcQrS4VfUA
308IDfP8KlX3u1Y6S1/O2C+uyAxStC5QNZh3CwLpkdY737ZgKukcNDn9d641w+23WMGiDi3EIJaC
HubnsXYiy9rwyWhketYEMHdaRfO5zv1S51hK2BAprMnP8CiK+K639Fus4NBrrbrvsDJhkjP/lckY
W/KJb5jwNAov62QcjRYmkdh5h+5EWFLcIgT1ertwko8bIx7MhTzchYl7lV7+MCMbxdsmv98pGowy
XjlnHYy2vKk/GMDRx8d1QIRqoY5TAMWe41R16nF7Oc8Uzja0PhSOuuR8PJFnjRSNnns9hyy4o65w
9cDhcpp3Toi+0A7E7a+WBrCzeIKpptDo7F7/FkIKaarryrShLiwlJz+ou0frPplDQokbdizIfHw4
3QRP35+N1ycjBA2HfOe+uwbOEPD9GB7UJKPXuo6ni7lCC9PMbXspgD/JbP8aqHdvuSGYm4vjpujN
aFrftecuu3cVOg3pF/Li3hBys9xb6hFcvJgUZ+AkWv2tSfrJqM6oiyjScFMXBOsLGdE2C0ZIqfsV
Zg9j8x7ey/AiwDrzZVZ5Ih/gz01vKHcWpsNynnkjQf+8Mo2toWidpY+ic2Uoy1Bnqw4NqQju0Z5Q
U8A2mH6T8cq5Vf5FO5MFg3jVoQyRxQI+b4izmu3MxWIL+jksFI2TkDCMRGPP6E4/d5CINhosaKrZ
1As1MyIgXZQwPW/OviPvEw/S9V8Zh2Vn98WK+YFREo86iDxkwFqnvsfqbK2Y4rNSifADtwLxqDz/
bEMKdqg6fXsY7FVW7MvNdlmmHsRx7aFfJJy1dpuU6rVPaXKsaT2PdNROGzIqIrxOibXeTJDlnC+T
8/A7mueeywwRqG7mPA3EJsgDhJJcDKnr4iE9c5ZKXHTQDdpgpAdajC1ygfVVRDQiv0WjB80gRXPE
YbviiyMNCnHFCFaCFQxMXpv5fUIidqxMKOPNp1wuS1CgkgoXDf7zBg8r0wv0UaUsbLK24a1J7gjH
EMIXM1vjwIvnKLfAiX9pfNdmcOuSes4joBQM++yVio702+00LLpepa7sfYUKS48chD13b6HtRPpJ
BYPuQVnY9tBcz5mtl1+TGIPTnpju/GkS65NIGVIg7Om5dWm270uGXL6fjghtmeFPeQeNaE101siB
bQdmgvhZ1pYBeb9w2QK8ehthfYNCpCRorf0KwBBoCQN/5cCE1LZPegVCxIUnUbwdyGzz8ZFDRHQF
Ogrc6dJPD0QXVV9vGp7UQbBguuSBcRgzxhM1yAaPfqhVOPkAgIaFtx81XtMkXtQfI4ccnRRjh7im
RVh1zTyUQP5jZZq0W3Q21iGKOoNF2V53m94F/5X0LEgyRm9lwJKmFW9MnLRyeKvGd1lS83ziNJ5b
hR8qEC/Rm5uH94cZlBK8FVZjUBKP49f7QnTUth59vSZg9jUKIVt76oi9EbAANGXXZy1SV+4b9zv4
Mg1NaCLBl1vCmW74tFtp2Zu+whrY+IFQuArEKAljXpJed8+mlk4xJ5DeFMEYYMMioxiWcCE6acev
nXM+EcHoJCUf/hCm4zFuctdsM7S9/iNwsQVLxc9P9Xy5rfpFZmC40S98KKlvjoPLrEVtN5istiz/
X1N6/JA8/+Mq+MEWKokruAmxrsCuy2UP9QDRuxDeeMQ+upzIl/YSitsSQLkri42JnYz0JBxF5LxB
//XYuUkr+muUDN9XgXTk8MpxLrXVC/F3NzQl+ixRT6MHXndIRmmyBcpYgZUEo/rLMgRRUaqZNmy5
+j72LopjE8/fGKAeniilHgaDQM0s6G0BNGGeBGUJcuDsxoOrJrykJx1V24fRjttSYu5ECIa8P2ID
m9oNuF9cFHcfQ6Stzf1AJsYyt1zX6W9zALNCQgKPQJ9kccCqVVSya3Doudt8jb3lM9wXnQTgGjYk
7MKl5/1bivrPeIKQym5fgN4kGPTrKV3yCNymwelbfHEemmn0EWicmpumt9Kw7cmU0Ybgv6AjnHIf
ZN4lGvcyqgU78/28UEhNxGTd2u9IRYcFDC5EjH60z5uQQs3KMnoiJyUvIJI3cxp2BvmrVCFVX70v
tVlU+MzEpq3tiiwyi3AVaFgyKF7MeegGP8wsgJ2DraVl80D0XoI4W7qqVhUuLkw6KWYoKt/RxDbz
UpDvKrNq+CU6VtKbtZNQbaPm0OjHiUjmg7VQkLNdRTX5ZwmGxU2Qm0/2BIHuXvzmRsHUcA3YUW+0
byWakeTMdq2WfrgtWdr5eeR1rAAFtFd61qMNB+yqTn1urzPjmpQfGGMMbz8ohnLLEDxhWechDUQn
A6WdD7PQUUMTgDiJXqS1Ezac1G8+g6s7FOvQe092vtE1U51qb2JCrjzs2NuWe5AXH2WUq2IGxGBE
HdqbcfcPOKxUW3mQQVWMDRQhA9EKaQPlnWCNZ0sVZcErPFDMg6dl2ljPTp2tgmqUP1kq6aWgxDsL
cdnc2qUAdIrf37/IO9O+UTy/hfLPB7meCZH8F90rH1BpjcxybABijLw398N4YkYXW97fW8EHXKzt
9J7cjGw8fDrThnqznOau9qSqMV35NTuV89nUKgooRMP554uM78TcaxEr0R9JLcd0A4a8HgGQSWDC
HhccTDf62evflZsA3A/lJJcDWCPvPtxuMW2084iQv/nMfabZcTUwtS9IY4sPtEximkD5JAF0ggEA
qZJJmRE/ib77/WITAZ0MoVx487K/YIrd2eipMUHtnvYBiXpufL/78aFSUeyTLyKmx8Qo96CQ4HvJ
MxqaEw9uTuQ0JEcetd3/cTDSY0uMHzRxLZbEhliU8bumWhDrUbhGy8cNkDfVdcwdctYTpWSK4xxD
e88hzseRsQuC9o2DmfI5TO1YwIORyUqG6sB8l+z7y1U5eJh3/2FZD0JQA3ue67xKlvNZUehIPEAO
/smjehsu39R4eOUv0Z8wC+6NoBtBHZF+IJ36tTUTRm+Kms2Iwt1JxvUatQA8HAYZpPZ0sQ8hL8jM
ILNQCa5jP6o1+tWE9IhEykvgkg86WylR96+I0qU5zAhI3P301KnTAPoT8CRuqMV4tk8B3Q6pLqD4
NTOyH/moQTb4uQ8a0wXsOQ7W6Wu6SclTNH/0qoywVuJqn45TYmzQTzyMs8tyBo9fqvud/O/+S0vA
OUoWqZVyNwbQpbpA/4AIBziU1T9wMgbRI9XEv5oFr8861+vQuT2f/eqbm/QhOiG3IJG4+ptfTcTa
D9ESCQuTDQoJNzVFhG56+8/cs5fs1Gej04wQmOMy/8ybMnfnuTu1C46VbsLtwLVEQNiM5p7Of0nS
Y0gLQlzOT+2hMrkhWwkbWtfhhcFcTQWi1aqLrIZtw8cipyPfB5D5u21PY7jlIk0ORh0ltToToneX
9qw6SuNcKorJuNr02ssedyqqxvyrscFZ3NJb2COrBf3Um2uwxxiGACJePv/MXwLVf0J4X20yaadu
1d3GB7mcITv5x3o8yf8n0xywR3Vdx2sHWw9lSU/OiSXQCoGFZ2y2Pc6rdi3maxyEwxE9K5hX22IP
JCmk7mLQf66QPYFqFOQy5ea+VFtybOjJA4r0Xwm1ws6hYcg/FouSd/mPLPTmblG4+YzVRvqHceLk
gYeE75uBHYWJsBiGlYmpFdMUoI/wbLsbEyGrLLo0K79U1RjM5QkjnK0sAatMKIkFUUlcDeRamtSO
LugqPar+dffRmkFjI/SfP25f5gIh8uXbuUc/uVxNhuALIBtWRxu2hCU2FVCAk28tFgX7PAyl0xsg
tlGD46ZubIP8uDEPe4eglkpTKhzzf7kJ2kT56hyVo9VlRXwC1BWLxoKN80uVUpG51BWB2PN3CeOJ
7dy3wVxBnqbtGcn/R7jXZfSQZvyE+HyYIN0z1ZCSzLYkv6mhEgKj1k5GMgnO4Rf8jSd8AJWRlnuH
JUQNAgYdfcdxWvhAymD9mezKxHmscifELWxBkCO9s6EyIqDRfTiqNkGtnk30t2JV5cm6/VkcxwPD
WLPec8mNnNTSLl9QrFhzVMj+jk+ZUynKw4vQjJJ/vKlO72PBNiJ32rwgwVoZOm3b+n2wyTBw05mr
wWMZ8+hOYLp/eBxgCZ4mo0zVngjFMOEgzRRkxqJLYlDE6/0bh4AYYZTam64CVfJ80e58v6/daw6d
YxT492mWnXOEajfm74Rue4BpH+h2/lZM5AXnAtF80BaWiMC4SYjm6pa7+bEMWrJQye9PYpOS5nBi
CZxgZLEAoT+DbaNs+TFlIZDp4hnRu9n2eOBZYOwtVE6EdaKFqiqf5xXRtLRnnkS4KaqCql2JcGCl
UffH25aBBMzMYmQZkD3roSQ0jMSbz2H4iuTtkvmCsABbaLi0x5DBCLyP8doWA1CzmIM2MmFUcazB
9ppcLerAZlB5vyPE3OgCJiu5O1raHq8f9T3CiI1xmV8Wa6fcilCfTkhl6mJJmnn8I0fWLd3CQB/n
7gg1i5P7jxMrnMmHGZuIxC973Rvg5knmJEmiiez8rLqzODh9jBlNtn5HanhLAsZQ3ljlLzkZ6r0G
+2I/x28xc/HdFZxdcvvPcZVx6yavcBWMHaGJzUDgxKpkkCfaYlj0kaWgvoeMvPt0ZH6Fy8z8HzTO
I+NrhD/q5STMVpclzTd1KUPDX/QhZ4unIUWv009KjCA1pX4PrZs90PimBhsPOKPOuond39u9p5pK
KJubuy6PNL4YkkO0TEzhJOg0h9AvQziignfTL+5kE2s5Zo1oJpe9KOZFv4L/8GrOzAj3rI0ms4Ji
yaBSSPdzZDH0P0Kn3Qc0g0llmC0YVHrAeuew0ENuWHv2sm974cCdpY1icS5pCKDvs0aYtdwU6WtW
iyZ0RgbKD2UaPSylgRD4HEk5YJPuuDeaCJC1hzIlhKjDlODf7VoQzfbhrSqOS/1dL04rZJX63mc8
bGIx4J+utbfyhxkYhUSkBAc8Kk9exZYJdLz4RlKvPllFB+I98t1mlJbwL0SuuBcQ0WDDyALbYHOo
GjqCqbEOsEuzCWw7x3eQ0g40mLNGcjXdVrC50sQhFCwvba4D+cPQLjt6MYQFQxPH82ic4ALpr2Sk
UmBM/qa+Q63svQlZMLlR47UxRI/xzzm3hgPebRVgN3NSTUW03EB/0eOkCCZL+T8WzMb3WytRuOMQ
Wv2mQPPrWuPufXfGDC1Im7xdrmK0ddxJSYmbBfS1CkA0TFjrdORJQ807c7yK9QfRQF9Xt5IdNpFr
lTYzMs8EFWt1lwN5R3yODw3DVIW+rg6HeNE0kcwqmDcwRiS3jCL1Zxi0h5jK4QjnPQjgwHiK5xSr
0oZLXFxlAhgRYytKkUPeJF56aQOItT1Gexc79iORf+P7pvygy3C+A8wMkU5Ktojv26O/cWZRhMQz
Vi7uciorYg5t9zo7bEZ4AGlLJiN4M5miKY8OiQS+UhS+FNXkekRlRJKePbfYFVCpjR0KhiekxY5i
nuSrFTMWp+Osmeijf+qNLuYPj3yR0kw/AgbKfsbAJP7nfbdG9mlwi+hwZeV8b7OJzS3v2Xyv9KjV
R7D9sxrho+A+TQaYjGp2lEFirgUtEjLwNk8tHEswHfvqYdHF9GsHi+NF9Zgb+4I09XbXJ+0TSiKo
1sZoAXSzSgDdFqvlvjgN1zsh0P2SWvzDqH9dot2pBOACB+dODCZYNcAhVjSEud4wVh+ET3E7+cpM
cLq94rJ6BAHjRssNpKQp9n3KSfGOK3IaMy5iIrB2gr5bGPP0/wi3wvx3Dwd+/KX6/NyzIYbSzxCa
Eut/ZNC3Yh1m7AIJzp9gAq1cZeE+SawYAr/BlspGSRi5FD1/wT+D7qfWgaiSLOn1mb7xir6r3sAX
UO5YO6WP//yxycywwu220gq1ooahchFD7qZxLZMG5msNjldCXlflWhr0g/aezZgAkbdieJNq+TAk
mxVcxpLodTT7sOF7h7Sn65upcVk1jVpXILPfdlwuiMkHMuhrplqGJQinLxIoTMGJ/bDb4kBifv5o
SbdVvg9qvLKhdc9yPBfJ7lL2zHkWaE2cEmiO4Aw+PoavDKQ24bethVVqtMeKXpB6djmErL1v376P
a/urYdvneIpLaTucUkBz8IqXX5L2TS7NtnDWIIbPswmaAAWE1IFE4UGAynWqNr9dLFenNbYyYCbF
QRKT/7VRKGLKoiZPyZ1KSo95my+rVsnOhRLgURHHFwpaB8EkZ1Xa7GeUUWO+sCzmKhEU9zUDr4xq
awS+wIxDT8uE4u4SfUwD/wu5Cv7BmlA73dVAw/CHxL/RarP1FyjwODai+tftUJU0dWFsgsmPDp5C
q0cr8enRhMfjL9LId9xtmSdCN86GgrXlPhlLla++WuMMKiueM3KS8RJyqu3yiba0S/Z7IgI4sTtR
N+ePaQbm5JVy5oAQY1OesV4wUPwDOT+UqoUL1gAKD5dT54L/BQEKotHLaeFs8MjfC3wDobWoC8o9
1hJETMS71B7IxAJKT2RRJQyO7cOjAXlSduKZrOn3an/OFpfE1+CpU30lvVBC7aomH1HQiKLzsuo2
aRObIXvqb38wYRzHeq4J50RKuFA3EltRJ9kn8VDlgMSPMMeuClu6dP2iMl1nnK1NmSBsN13rJDBq
8BnmSvoHWZfvKwf24V6xKWtA9vekUlA7ZGXXPhgBBTk+aBsz0c1q1Fx3UhBfd6DTFfjMS5B9KAqI
BbN4mD2drkq2yhulEGR5Jqo4r6GtvY3PkPJw7du7mwfN7OBDYyQCPqvTvmVZIi8012hHtfpItFiy
3wVAlOWDdJGUvVWTN89eLvBsAXE2KEboExZgRHPkO1vViYzzQRxR9NBGEvRb0mKGS65j7szTIrC5
TNHJ1gthCBjuiBr2zDkUK9SsevItZA8+0REEQ1MVKv/v+PSkGLwuXLSune8Uu65mQ+uCoJ4hShGr
FXRb64eDYX2Z7QuZWiQEdQE7daSZJP67dekwCmsDc7PGMqWoZKvko4JKXTpiHLGJtPFZP9u0WLxf
CsuHzjzv3KDaAbhYosojNWtf+qFyUAk3gXXyHp2OXaWzDzbFlxnoTerL4LVCPTCmTYThvhp44bmH
OIrc1app+ijIZ/4RZQd+0sywXrVNPoKqRt5wy2IlovTVTfkfbVcGBg853i/RFXJWqqETuRIN+x7r
KlFZKDSj2L5jobuRo1K8FMhwPYk1A7dJjXsgyvdhPmn7Y+s7nwPY1T8Lyk7JrhGkoJIWJUbGrSR/
KxXmt+bE2KqrQiPJ2Kxr/KUCRV2fDt8rgIYVxEOhLeKgyBAQY1SectkCrS7GKsP2PT9WT9QS0uyf
zapF216vY4NYV1FTznbnrtrVs6Wd+MeqFAtfveFIXvRJ6YQxvAj3YA9fah3dqBbQHq0jZZp1hbXW
qb1Hec+p+0mCZXrESfa7VJ3mgKl7yhDo8vnA9aVVx72bqT/WiOUpCXbG9X2NnFluA5kw+hwEWg5v
JPJLXTrbCtrDhXPc6dJWTZ+MAdauDOZ70viRsk3QRIR3MC5WZeJzxlhKGeOZRngfFfrW1AIR6hQH
JvZ5lgZN155rYyzoCHgrgnxr/EC22agpO6wBRN9TMLNetY4JexW1R2HzeFoKgPZLMxlTNwn8RLwQ
lvYPbpGHVYYJ7+jQjnSYVj/Kqx7FudHJjXetS11Mw7C7RSa69JcsWF/g7ipvy8DbgXc7Rf/fIEbs
99/E4NthIhUwnWLeoPyYDgT1f28yNYH7Jfz4xXgfnwTisZ0MAsUfKqKVU9LN18qWc7K1tLzFpcWZ
Ci9HWSzD79OnnP0jIoy4N7cR0nUU7wyg4U8NdE1/LhRxhi6ACOs7zPyXqCDfcaXaFkfl/2snY7HC
OAirZfxBC3VJ04gdX8p4RyJBhCLDXASDjqqos5nsOP3faKlEiVNoBN2EtjxbkH7rU7DV1MiHogrs
c3YqNsHe1kC5mGPB/Byx4Gg7SP+qdf07/iVGbCwYKHPTF5IZkn2Ce92YJRt+cj+4SXtT4fsgq5uP
UFBWZKGShNdFTy01M+WdEvUinrjqZc6/hKDqkX790NOqjH/RH4GO2+9HWorYizvJcLu8ebzKpBhT
R/zgQfk48f3gX1Tl3uEkohlVJdTDvxzBObpYJUP0PMqQWEHOVxnKhpSwXhMRAZ1ckyvzazcGAL+F
H5k/BgkFaz8A+4V8kalOi98wY0aA0wURVkR86CIqUzZm317xc2iBcNH/TT2Q8JNsONy5DShNhesb
pen44L6NisAod1eNqmQlSZGgjecRF2pcMGC/lhpVcATDyit1J8yUWrhri8dG3CVyKQik1xlKxWVL
6RWCaoUkfKhL9ZMMGbiJL6wJBwCli9kOAHjPulB8SIiYEmUM/0HLay7/hgCt9zE+ZfC9r9LIB95K
yRjNG7JNhSw48aRN3+CjCjG/GjT7rS6xcWMxS+Ow4u0eIYKcLSvFiaXwyBJ2Vrseb20/+FLhQvNr
jDGX3jZIGoz60KBEdCNaeDjMpygmVHGUZ2bYXB5NVaw1JE38EohbAD9cxFyyLGEuSN2ovp26Yg/t
u4ahUtCm0qQC0EBFh2NlNLfXaG7ZOin5hZGANYctjlso8R/SPzNMJyeOTLNYdxSZYyRW+8BM0RB0
Lz3bYUWEx7emHQ4AeGEtAoU3Kxi+rSo+8/RF8ps0z3wc/wWNzfkXNHfBiPRWdZ+7pEkpL5YB1mb6
ApHOdGM4+rgzt8Pmx0Aj3ELbS6B6MjTP2Vrqt23MikYZv4Q/+g17Xe4rZiGWU9yo8A5TagS61iwa
1KDgThNUvIb1p4aPzzgOomtCiBV04LljVP8ZkDD//zCFX1kF5mH/g8u8r0AfGJlZMbhvlNsiDk5K
p4ofgxmZ/pk4i+4qPESOO3w8kWH4toCBgHUY7uvhHIa7RFTWp7MHappQS6YG8GJu1dopAHJAGJMP
zFEVZE4Qi5KcqK5ByRUcR/XtKfgVtqaWiN5E//LbEoxlT5E00P8j6bnuzSstFuy9qKNYR++yFnQF
IGKJOHOZfgskGO0UGHxq8ofcEZKzEJtM+Xxy/eL4hh9mCM45Ro5lc7Kc7cTikwJt1zA0TUdiBb2I
uhz6KQLGHWdPHfOCwSZLCKok8sus/Wjg1Np4lPHCWhr9aQVNLMCwAU+74zJhQJE12f0JtNvlvDfx
cpx3CCeYIr0M3SsH481sln21UWJVYSTdMJhbTIBD/0/KcUeIMelWLPbJegJByeYBNcbr/llR8qXB
euJ1192rWhpIZFqo/qPVMywoTsLb0+1r8qZ4AsN8tkHwyx7aR4VYMjBjpPJWTkjSjZmQnXQOOCU2
ZWujsGqv9XNGNi7/WPmxG0vBTi/uAyzSea6o7a415uaPV4FqstY97XokcjI5LBJ17ti0pEHCjaR/
bPyvJl/eM77DaFYOGuDNAU58PwokRBtdSX8H92GQXtAmR0YYcGebzXRFN/jAPJA5c70NSnQJ/qBg
trmuL9k8hbpZjlSLVQSkAh4kBc74hUE3SyNdMHbouslSFpXtojt8Bh5QwSgCRb1a4F4/lPfOss5b
n1jDRosG+Sg8oLy4WSL2i+Vpnh60g0kt1I4i1yrx5QLqe1xZXBH0Xq97FRIPjWe10/ABCJiqOJV0
r0PeGx5E3FSFb4q3UsTCtwK2eAdeRjOLyaNH/psCguFJuRwHjdy0ojDvigXiuk6EhWgCF1vZ7sI7
R01/cB0sLOm68DL2fvRqmJlqw1/v1SiplqkFJ6Hnh7vUBxSXfrvesUabXjGYtCWukpSnjqX2Esaf
G7sTFxC7Z4gweeEeEPE0JN2Gr0hj/9AnDpZhjwSDBME6GxyJCoELMeLcBDgI1Evhjcgx/XEz9ANN
DL4jj/XPCzzJX6vL9XEAVyYlt/fPRcqpGXeNDWSQCSvREgL3fTgGFqWuaCwl5Yx8Kp8bodiwb42a
y7UZeKWx/PhgKa+H5JVlZnJMW1a+SzRpTD6UQu7n1G5NgtMjdEjZKISmogpsS6Gc7iItmGI0vurV
NbI1vxl1Pk8GRs+NYbw5O16T8JL8mnzobcnqwVxCS42+Yo8NlzLoCDnGfGP+kbrEajaRbCFYMwYV
ku8YwWcQRFqD/QHgS5dZFnkUzKO8DTH4ycLpR4Ljb0KsomB+HaTM2g/eL2U/iki8Cd3yeC/yB45C
uFK3c471w4FEyiUkpb75S55I9BCLHdqaK8je89XLmsuTpaMBb9mcdb1MBw9wlJ87zqNcPicaSn7h
1mqIaWvxmf6/v+6fGvM0ivGDS/5Q9Vj5FLUgxwLkPKy8uplidSQ6RuaHzdQIbuTw95LPw5cJbDRj
BkJc5XgSmLJqjhC/ppkj4cXQ31Z3NC4an45/QNDc7T5nAc2etCQ2EtM45zBFFWlVcnvbia4BE1yZ
0f8HV1UwfMQ0sGwKFZ5+q6WL1W1d1vRW6RJ2lk921xtQz5WEldd+a36proa2637ga7EQjpCTL3hp
knfRC6MzKdI7qTs4JFjkYjQA+PjGUYxXBKXz4NK2HR+thsPbxHdU8E2YkgzwsLtbayyJgEaKkYlk
b2lgGlVfc0+APK7l6kL/iQj+wn+z/wUbQzdrY7lkXGGdwvChaPPnBOQuEzGj2qW4Q4kHvjFS2nkA
nqjAzId2ANqA5u00ZchZcvTIxt0sf7fDOis8ZyUvWQHncPV+zOSjsOrIdv7L9Vch9av1elgRjW6z
HuvwPyDunwlmiVFgVIYre2iRvFI+F/1osj008PygVDmUh0k73QjgNCml+G5q3hvc5Lf5AaldSQoR
AQKmzUzE9NFM9ocvm6twN7mEY0JSkgFga+n4Vrt8i+PzX5Xd+6f9jbJlA31890pwjjzEC1ix+wZE
c3TunXYsvvw/QRwFz5FFt2oNs1py3RzEuj792mf484Y+25dQjvxi2rp4TfB0cQBzCGIhSFJk9s+8
NC3dHmADTNHFOpve1pPpoB4VA+DgKmCzT7RTDcyS56uEG+uRs0jLvzMSHMFQB7aCmGRUoUKD40uc
tzAv9zmoRGYFkuIukgKxBzTvpsj7t5tpJuR2O2AlaEIKNQHL9rGQSH/ApCo7xzpXbFJvNkJkiNSz
yY8J59Ge0HPoP8W6LzqSz+/+XLjVX6iwiTTeO7SdEG+ccQDL09wIN67pZB8MHqI29B8TMpVl0ABX
JLarHHV4bZDMT+QQsGZwQn5e30Rwy7ekbWuSKpDvYt8cF4ziZHHF4vvXmgmOMIuO+4pQWzFMxuXy
R4L2Dh1Ri/nW+g7mDEd/IY+jkVXIw6CWAD4ZmqVUgPcdSUki3qKTetNZVq65wc6bEGHANIFI4qI5
pIMQeN2eDjsIKpHu7iutU0mbWrJ/bH1cFMka/W6oWcPC8pmuJLFLa612imsON5QqzZTGdtibXSD1
lSmt2t320EgHMc9y5B+WpFPY+e9h1mcLS1J1QEEJCaYDUrl0eCCSR3jj9HkD2innkMBNvLBNF6rt
6kioveapDjaBJM9RyIocQsPJaonsWiUs+eHoUfh6P4AdaEozdU8gUxICeK5GAAc8O80uTR+nngKY
+sgMmSzqLXvVIUkj7zEHAlw9yw8KVTwDs4amY1K8VRrVQR7vF9Vp+7Nra/hAivgB9cIQyEsiXgfr
qaEjKjwipQWYFLL6dGVijQINFgvFSKJnGXJ/cXJrdQY/O4OwDM1yWrB6qTbfdFI7ave4KK6pXfRH
X69wFJzUj2BWyS2a/asOUPZcKmAby8Mrt3bOMNWYwEHRIaonvQvaFnQPC2QiSoZGPgvxZ5HL+kSx
eAEtjHOY7sg7TwF5ifHx6/8AqswW/x6Vxkdpv2iSFynDj4zXhALti0HbeB3XhlkUxHwctpBopY1d
L2SSh6yhnXxDv9qW5vsni3NTt+UXkzXoFkgmSMD5Uk5m9COm9IpP9fOHSS+7RKtYUfgOC8RStjmm
xJFK2p/YpGnmtbWGYN9Ite/5ZicWofZF62IlfpHbIYMYQAqURVvb6V2OErHbdImi+Kc1kLb+A/B5
Rq5Q8i6VDKT5p94bAZUguk4nDCEj2RsTpM/RFONFnaDEmB4dUR7AWNSA3+2PZ4mHGrqFuwqSG60B
pnwNjReK0ZPFYePHGLZAJw54uVg4bORwBLG+L6dzkx8JpDjpoih1O2Fyeorz32WO+eau0eOEifyH
B29CLwnNZNAGFBQDqM2qL70axDwUQ5w4+/BGxjUyRBh5R4C9hTvMtP2e3EzGNMV6ncbDHSoYXC8J
t0fLFNBeg0LZ4Z6bXhT0+HOfoB9AIGmCWCdFSIf4efi1LlgtwQ2RLa4ilCd9QWKJ4jUvTg25/R+x
TB6GLoY3WEObCaER99eKpXr66/umy2eGaSqSt4OWnZ9mSL9PTS7dxkxi0vcAJuM6LEIf6MDfmzbT
AQ4XlMrb4c80yIKzmUckYGtSE/G2zc9EQczX1/18zRovRG4hiZ+jlrq+J5jaNWNRxm1p6RcNi1Z0
Kj2vF9hlCfLiuDg9ozXGVVQnX94kM6HTSB5797HTGaQ00F3bMI5oj0XjzXURmJRJZ6TNUeeCuzqn
F2or7p6Ts23bmOtSEhrdDaY4GPvV5MBoZ8VK04eNP22hjbE1BLduABwmXMQfLsXp5PfYSnVcjvbc
gHlYpcW2NJ/ivetVXeIbl8DbKt9dLO9KpMsgKYkAezbU4kGB8sTrguTJ4BtWko8Wt9ldFFQvFXTp
GwN7a9pFbgkvtQNDZmrNru2/KAHIi1IT5P/M55glYIFHaOV6ZRfGHvw3DGHFAtxZ2iKkeASS2Euw
EemKUwNGLgt82RLZfQL/VYdKtME46uU59B8iYDMzWYO384kM4ftl6+2WeCmavx6luizDrFJkcD6f
ELckZXy5qCMEhkSIBLn9yCSQGQ+vjrHCpPG6ZhBj6HpUC43Po5I8ZM+S+3wL5ssdsTyXolWPHf6/
4HWruVY1hHiZ/IV5m/KDkGQHargyeiG8loJNxfKTO2UitBuqHDu8zSx3wZQkCwp8gTKvUxoSOOgY
DhV/AD55fIIjtJo8BHT0E1uUrdGZDmAW+tuo7pEUS+5YnbhaQS8iVGqcrcdDDTMFPNECUHA0Rj7N
wd4QFh7bodMtGH2EgbaEcRCeabvAJaOGluSn+UIxUquhsr0O2tvklsY/zqSbPbvtYyHnRY+Qt2xJ
lhTH3OGPswb2K/850YbtC2DNMe/xhawW3ngv7KQhwOWnOGkw+x+cyGSOM6jtZ1KmPrnqcBMqImnT
IPKmlRU3fpgKvRJOqeT69Yuc/obGftUz+4VNYG3x+lR+JaDiDZ1oAWyGaQ2YcRA8vQFBp1ougTnE
BtOT6S/kgtt0FC+yjTEeC/h+ZBCetwIR59oA+laEX9hFRLC8HQ0Fc+Jwqip3UdZ8GHz90VPyGM94
viKD3negbGUctZJ8WHnYm93tlgDiQEGV91C51/GFLmUFKCksmek4AAnPXpOwbEdWDe4owA2B1FfL
dsAKdMTD8m3HYyrj/MeGZkbvSfMuRs9pVxp6zp1Uvu1zbmHT0eQrswnBr9cfuYA5d/ZLPEzXpWr3
Ri2t0sFSEUkCory2a9nARpXhOm+Sojxs/2telfeKPmEmTtcEp79bH0dBafOP8dh0kweQwhqKCtpr
3MUx8UUUhLYFj5I66hcrDsX5ocAwL+Y7xOXprXD6ck9HiYUwgqMwKZDj4hpoF8nXIbGhIM0MdS2E
P22AW86AlbVJ25+KkwvTTr7pi6qx0xk6RxWf3w01rCjrbTPWdNsviS8evhcwgHXfe0zgURBStcm8
ZfUX2Rw0S2HQHPb7OsfR74A+XuAzQKwwggRoWchFKSVQc9Ii2YuTxXgrTwSK1SX1ngTX/G7YA3sK
pFq935T+kaXIFTqptwNSHwsvjPG9+ahvA4b/KLMI/m7Ci705Pr54Vff7KL2n9AvaGtreR5OKfpfD
uCQpc3OaI+39L8JEbbI81WIPv7GO33biOASFfhwC3qsWKNU0hAo3y5ztWWjDSGOk5GPYaPEplcT7
de6Z9NOczM0GjDNiQkIkEwMXGu5EN+30W3uUGfM3+s0G5J45tsod0k47SMEtmDlreC5hgPnGQYfX
PpiuNkHntGFEbC35I6xJpj3dEmPLMB31IZsGHvgAlQi4yqsi49abeg9Z5hizvCOVDdSIBkj0iXz3
URyDEI1vvjE9IBk+p4wQhyIS4XhO6jC++0tPdmWCJA/u9HD9lMsvXMLbxVzuuXulm6rSsRYDIgEJ
KsPQkIc80AawuGHg72vowWsRU5GPQC5DNWjZCHMukEbM6mwA2DZBID+hM98Vgv34rcC9C9XenIV4
XrUWPuJDOIgumhRa1QwS1C8ftes+gBeth92Cz2dm/3f3Pug6IWg0dlKqqnsxP0CcEOJ/PNfyaHiB
Ja6P9Am5zyuU9KXQLSdXK7wmNBmut68o1/DSaOXSPaMbPSvt0PKKfmv/ykLrYqJK8mOH8mv92698
+uqEkydYwuFQgwCeHZxUeK6BfX8M9H6qS4WKBMxmDv7MEHD9E5nko9gXMYabQtONliHRiRIiYHl/
6puPJumhZVVHD7o6eOoBTWdWlKmnrLZxTqQsGxRUr1a36oAFmh3YeDDggwy3c0uQ8HxiCwljd4aQ
nNegNcTaPfPq3cehwqSS7PRIURJsY5zCaFN7b+Oq+eTbgQTZNnrx33k8DwD9P3vBvudbbb0Ucron
7Mx55vJkwmIhCX5MaFPnudSg6BZ5c+9hXrxpSZTfjKApya4l//5TR1kIE9cZA876QADPiH4Ne98x
Zjle1zQg56Xjpn/zAPNyUb1BBQtVMdeMbp6P6b7cPGWh3ww130eJJNtc9x5SpsEoysdHb+/hA5J4
JljdsdMGSWAcp1cMFhrQBAi6qGhQGsubWbFNwieWevy2DGBmZSrj8raeILkIczJi9VVcCvkZPuvG
m1Du7ubzZfaRZHWyI60DPeqCMfTTJ+GPs3K/9ROZx+cqPr5VuIvGrCEWtMbr5xVnAe2p/AwZwiTA
aURPemw984GLbrq6TN8eEvY5AnGX5DLrE77ari6evKVbwGb6Sz80OjtbJ+hxwCfBxdFA0yHaT/Nx
427GS2Jw/ZgAlJVhh63cCPBUPJvj93rb8wUz4pDRi41pRi2gfLPQS/FOQqJDikGN8SzDmYhOaqaa
GtjYtJZ4CHBCB8xQjmfT3QPQu804MZuTPXGUokKUxdvXhZiD7MwVYXrumLnajD+uKuCGIDba/hka
TROa9Ai+ubI+sfJ3glRJkA+hCMg0RS0rIp+MuF+d+lVQp/k3/C2nSR7j/HsVfR4fr98zv0KgXmZX
ztBz30YV4xxWQxQuqdKvLKKdofNU+wU5gEaEA3ODaUfDexfPAHjFc5568DgDH+1fkAzIZqTaXby/
F8RhXjzVGUjGrffL+Cs6MjlmUZF5wHAfwNIAh5M7SS2tT122YWYILCH7PVqKQugZMnVBV0UkjrNd
0vFErw3k9hZkUTwaYMUqz/2smH5dao1fDBOXIeGUrscmt5ryOC8wNt9qH8/g6LL2DATcPC5Kd5wH
FNe2bw9wWisRdOpHH5DJ83M7/sn7t80eRCpCo1yd3QBZ3vLymbsvxQAd+8DmsmTtWlYa0mDVg/6i
FXqGz2xk0hf7UoH7ERkppdXQ6ANl9rjUiTKDR/vo8rbSjdy0GxX3nuOqWH8lx+bu8HQHXTaNCnws
H4eym0myvJ13Qpkt4OQv7YARz+fX5uzJJr0vEwpgaRjKZp7rd3aJ4LYfXcntVe9sYbA3rsc5lbWV
eXRDpd75ggQSrenDozCtV6tD4N5x4EL3vaa8cb6GWkuAyct3bVaBhkpwVyDRBowIVeNXiOIOv40a
sVyRhRx4f/0AjO/8yhYxlSndek4tfkRUvwOAgLaMX3jBNuQOSsH/Q2PejKaCdxN4Cm0C8FmryOQ7
d6ug6lYpxS8WCYshxuI1Ujyi0Sm9ETYIDuHEf2zcnFHyFlJ+yY4UcrGT/EkcEGpzfOxcNXb9rl2I
XU5zsNaGUSYaX9ambBm+u/P5QOhgxpZ7zvwsmukEmUYwNDoG0QOBl3XDEclPJe319dBB6JisR6Sg
VwKiS7u+DUVBga1YOqzvQP79F9PqSK1MjesCWxp2WOKW6+uk/B+GgioPVGRldwTWI4CQr7ErtZaz
ZAw3qV7QPVlrVXaV3yptUNwRcNoJSLgmZl16ld5d9ijgCIzdEd5h6MOBTvuI21d1v7GvImAG4Gtn
1vzG0Sg1KXEIQ0xIpPPWnomDsaJPF6xwibp7somEuseHUjgL9dHF50BUdTbZ2Ov4XAIobDiG7u5E
BH6efr/vC1zP6AzZbMOdXIkli/HQRxoI9dLa7Oy+P2EfssVVoK5yjZwfEMwpVXcUBYJPUdlttWRh
rWOg7sKjB2wu7t6ndZPm0IM6krxo0lvdcKVN08T2iF/XqLZxQU/XuWn8zZiEKNQjB/Z7VtPVmuOJ
LnVEGc+DD7EwP+eMURpJ+75LeA3TIjMkzDSU3bW9lgOOcUeTW+3hcy5MCPVmpjFoT/nnAi+4t1YQ
9wZL/ZkVT2l25fw++439JwF4XCagMaisqMEFMBa1uH4rsvJbPIQS4mbyaTE1W3CWtZRL3fGUc6pL
tmaQzNNhk8l5GUXFrsK1gh3Merly77llHIRhq/YRKl1DRMSp1hT2rbgbdFo2Zxy4Hm0KZF+RvUfQ
dN7lsEroXq5cPatKJIkcEYEDaWOiJLctAsMxWcnJlpiStjh3uiE7cbkazI36FJBzQX/s08pjlyw7
CUwJggPdcHmQSKFii2UBTMJCyw1T1engAMvBf9XFcvPZzPaaKq6D3hDAMNCvFE3unaQ/GieL+tcn
eImHy5CB89JsHXqGGRMBp0wfivBC6BCbIOGMaWeh1wWozvxp1MGYYP5unZ3rG1LKfKrMU4XIxGp7
3+Rue1PoDTV1PvZZYsYAKtiMnkz7mqASEz9/iKaYbwhBq5IvSLptFPAqxB+Ru4tZaMGtiowKmxsA
u1ZuvPmG5ssezM0h/B0g8f9g6hktx0IhEUpqhHvBIknfVd9lauK0xwnhDmJfvdfrB4ASCTeS8w/O
+pqVKwAbfI9YvhTFSiX7ByqbZ6RJIt2OLqQSMZP/uzFFH1eNK386SC1MsKsSP3jthRRu5f5Mi+lo
HGme1luA7EYgN4zJmv/Vpg6RvK1EVAaVmT/+FTw11VD8YWdzmyOqxIFdgiAdX+we3+CCLnnMczCV
4pKLY8dN6ntdXVz3daWrqEd+au/49G15MGcZ3SR30l13aRnr4DuT3bvr3Da77Corhzqyyjl+hb8D
tWBCzbmP+9hj5LTBK8zA4r4tdP0um03lCrCrPSShoMKFV/ySyKHu/Z/Vi6icl1p7tgJ4m8D1eE42
f0oH6Kfglu9VINBzuhXcB77F32sf5vlKl4e2gnoLZO6qNbdscBWmzpf5GaBwpFDM00Ju10p/FQaI
bm3JppAbgZmUX/2Zqrl5FJ4Hc+aTCKZFrRlg/dCKLma8mrRoXOohfIsr/Z0mwfMypSGLLiiyYaa9
/a/M6kaa3Z59X6DD/pGgZXfUqs3uIeA11/H7g+jL/zEhAP++Ru3vvHKO6qpuT1KHUDkOzBVHSLyn
4V4ApqbESOJsg+Zd2f9MNIkajazQWTVQ8exPp7uOUBrDXNC7JCNPm2YT5FzSfCv7yMucUmGSFcze
AXPp7KFgCYdm242UFNpkZjO6AspPc2EVcBHJ7fYs9o7CxUaX05o+q9a/W/fnf/QO1RaaHjMGlvY2
GCUT1SRskJ1qLH02Dk0NH9qaICCSrxix8cF27cA+ste8YNBG4jQv+HwocJsdjNuZZxlRFQ2+BmeI
vtetQvlfi06yoIC7LjWy1BXUJkxqS5iZsQKDTyDPNtQ/MT+HNu2v4G3MdLw1uzE9HpNanHAjRSQI
MLtrKlc0mHZLDYyD10KUpddGAPMyljKxI7pw9XZcDeXxvTEz3zs6GLOESW5peRHRDW5I6aP66jlf
74J7pIzjA2M6byVgP9q7Thjdgmgyw/PIs9LfC6J7AUT7l38WtqVtK4sthJ1mLUD3APLhP0r2RZ+f
RU+w0vkimmVow6wGyg8zJKt6czT5fEYOS5G50h7/9nHy9ooOeXRMHjjCHdmBTXQD9FSPZPoJyl6s
TOBMj54tzdYX0frFaf5psGWtihEyX1QCbb+owXf93W9qS/prxIprjn7hifUpCx4VZOKwtACVJhF5
E7yJsbBYzTRky2YEmmEI0ecv3tpqdxafPsh01W2+P3PAUnF+ukmFxF+JB+SG3sO/kb4RJxKHgEZw
RGIq4cwqpWJxEcexh+nezQHpWAl1LEfRNpjF1nAPVtL4w00nv+s7pjY0Y+ah2XwK+s6Qz101IYxl
y/RK4MsFm0H9rshoGuecZ0NJQ/bFrtlHd4bEx+nIE9iWwwAA8qfNeRyWlYXZ8ARIVJCclQclB6JX
42wTbHcez1euqoCXjLDG0y/zfRm4HGvXtZ705zQf45ENPQ5ay7Oh9myWl1qUe55PQ55I/+akZig2
bRQCQVVAHn7lzFBmGa6O7ETWsDPhAZ0UJLzGZe5nJHnUNbe+wGcTE3ry+8qAodG6hdGuRTv8L6Ri
/Cj02ag4KUT5KfUZTvhDmOoqm11J/iNtE+SxccX6Qrt1pn8EI7ULm20TtdUCM0ay0KIjVeNn4Zjq
BOqkt2pNvunujrETBvFVP7HfpVZxakHE8QgBjfVpVhEKRnwQ3IYMOt3OQN80MPNbSIFB9LuER24u
Qyq9XuLVza5zFqVDXAw2prmo0LF3y9YVePZSuV6on8BV7GyWyx74ckHrG/6fi/iR/gR/mA8zFaOO
Wy98hj63bf51SvPArANsMyISWtDu8dqQXFjJIVJ4RpNkb/m3TpiXQCvF8MIoFE6lTT5yBczmtMBw
kg3GFy4gR5eNmXPThyfT2l0peEUYUPbWGdpLXWyQWHidbyZNiETfLS91bLNEWXplHQLm8ACJs6Xl
d/aNxfc/TXW0jjnxtprPBl3FoCTa2Ty7SsNwqOphwXGSzg7QQtevw3DgY4b4dOHrywI9xhset4YX
SoehiC4HNSQ74gBGz4erFQSHofPX53iYr6TNPxIULx4N5gSi1YSOnn7MbbLuT5l48Q0DqOkpwePl
HoPlRGNO2G3QwYUetejQ8zjiJkbQMJ37o5r9QMw6y4hd/K1N1PBPBsiPFta8LGHfDsLnEQsij6Ps
/pYynHHkDq9WRtYXv+5mzqVRF+M/aRodNSl3RVpJQ8RzZqogXwANzZDiZ7kQcIz+IxH8qL6UBKrR
BvVCq+pxBNFjBrwiQDmIUPAOKzr14lHIpvWTvTiB5My2ktxqQ6r/dFuEdh8EEgmGXFeMeMCpbOl9
nDKvoMwzGRxi1JGfUB0zMHfzyvmaAiP1PoQwNaHti03ur27UDESh0wp3U3gFZGMx/qdKIib+9tEL
1+xQQRTddlKErPwtCm2iiZTH2HhSGB3nwrY+SgQvZ3bWPKqcHuESfSnOtEFct02KgGPGfE1d3zoq
4rNC7aDEObVoBUoFzUb6txA+2BDCLVCipUHETdckGaUa1qT50baoEE5nGKi5OFQ1/dllhxaT7Cr4
VqycCYKlGW1Hjx+eXnD18oXMAlKSQAnAbaPV7TMpQONsAgVmSxM/PctvsM+sIXTw3bcR7p4cVSH2
58I/djeIW6s0Bwa8kGWDmfMtl++OANGgoMR/B+gHAZgipcQ/d5le+hfqzT3nb+xCz0zYGpkvJJyW
vdTBzUnQIwPyDR/cvHyVOB9EVlwRq90dZ59LJK7lzYwCczjHX8L/5y7GKrPJx0l8qqVNG+9JM8aU
xYTcHgC1i92keyJTm86AE8FUaqr9E92OnXPKMAo4i8b25kSSVclj/CfErR+swhaYQGf/meRcSxX8
NsZbnmzbG7QlJzZNrEA48YqzLTUkhXeOogZE7gk2ol1yQtLYnsT/TkoSNWU43Oodqbt5m/zJ6f/M
DSvMAPlZKgISA/I8nHsxxEaJbDApzZA9lYDSZGGb3s3cXzDtoBeIsIMQx4iyOtjXNVlOuAUS1vcR
0CGBlYbyyefW+vTNRq/ckN1fUHq5XumnflVaYjGWbjo8dtGANOPpm0pwN3wq4gdXTnV53C1KiSp5
OW5Y4+4jAaJTEJuVi33AW2ZyVh6ldQjlhxz3I/71dYTMcAUMp9YjMForLwljvD9aWRivcqbojAmV
GLQPPQQ36KdEUmE/gLqTN4VRvn1xj/63GeLC+Y1mt37rj7Vq9pHSv8xLK18pQm4e0EB1VoiVHBlo
DGj50BfhM9Vj2fMPjoknz5E28vnaOvfDigRmopLPeAm5SEBdiigvaJHDy+lllFl/21qpjueVbxa0
rII3JXcwSWiM0+c8pngkUqAZaIycA/IgFayBAwfnErmTXtaZA/Zd8vn/4Sw4maYd9I+SL3AANmQc
9CoaznwxaP9wvKaAr+AU58CHgxXfOUan90Pm+cMDTCH3q8QDrq24zvZsaOlFPuRAnAy9CzPZ+sBf
Wm6ftrZUrTzuh+Vcwrc+HrYLAK3Lek12HqugBL9/O+XaNWFPO11CliQUeYCuSNDQputH+mjwQ6w8
MZaDf+Yf8QrUo+WW8VmnkgkToEcpyvZIggFjHh10kEIxII9YV1juwMId4I7Lcty3BVvuY4/ip9E3
Q0E9T/BmQxKW5E32U/cJINitvNq54oJRXNx9LXSTlkEEYuJlbsGhfdOLk5AlzqIFCYnwYb1UJdso
w7xbx4eS4hN11+bQfpxJb/pMW1+a8/Z8Yq8sNQz+CDQAavo3aKfTpS7HR8AawmFKSeH05DHyQfy6
Xdqni9XDSJJ58QlrhnpaLk21Ux8XPlMX3p8UEqMhXeucnSzxH5uPgdhNADyztJucuQi4lSqF3tk2
e/k8CmMp9HPUZ36oMQN9P72nEQVQVJo0nTCCF6bTGWK2kJbYFkWStupo4gTUm+hnLxhhtarVlCO6
PFkaYKX+oerafW05cWua7Bt/IDX+GuO5tuoZcQqJioJNFLOHcPaKbvwokd19ojDj8/5WFilNRYAQ
6xy6qSNbcPa1xeYT/lQ4Zfugo6F8VD7vYe1pps71CiI1P3nL1bbska+3l9wvQM//S9ZdBJzTYdek
zErcbM+1uO4JrUD18adgIv+Sr8MD6hSEL5FxkRqdDAmaaoi3yvFaVby6SLVhT/Bcaw3cb/Ja7otW
rM8hdxULVl16nw0r8fpnchhvokaagUQa/F38S4Q5DCWGNqG4ZWugf89Ed+MEQe+0CFtvRFWIkGOY
0WJN/dnuVEcB9CtNwxjByovx641oFrhnnxAoYLVmMcSj/DubhPE8yH5MVggJy2H+2H1ZwSo4jV8D
D4GR+/y3nkY80zRzNBeCA0ar7/22GTCFAzjKgzgND0EC/6f9U4av3Ok7yzkh+kAEmXJ8zrPYqXb/
iAnzZMnSfsLwl2JA7CJ8x1VWKDNFLXZPtdc1JtcgtU4WI8q5r0UEkB05SkUaVx37bVcrmXJrXdNW
K7/aOBRNqvYdNSm1sYjVFKLSK8IFAbPlGu7C4mfWCQpDyYNv4yAKEr++QnWos8k8AJRhCtdlqNwb
7qV6WJjQekGpFB4xZCa4tJbf2F5ut0/V/ZB+5npUih8TSoeYu16R80uTp685BRBGCvR0i6IjDa/P
UQ5EwFJIFJcnTC5evvxKvPVSmuTvjtClkv3zv82Euubq3C3gjEb2ZqwGjUzMHk8YzyXBzTA51oGz
xk93HpvNIysIwq9UzSnljUa2WpW09pNR7eCjLZ86nz1hNeDY/AW+z6yBdeZSer8xWErOxMvQMUXk
0xXsRTAW/pKzbfsAK/V8fs8xHdEreSUzbRNWmJXQXGmR2wfqwJz3XAl8TCslLi7vgWeUjFiL7ySD
meAq3SKvUOcq4mrpAKUBRnDrlw0/azdMGAKVZdjEAMZ35+nwJLonx+fnf8Vn3CM+IrUQSd6m+l+U
aKc3ptIcPTq09ie5D++eRZypokCLYhFD3fMCHWghGZ5qJJDQmhuLHZXC2flTqIeyL/mN9pjfxORG
tcZRqv8lY/TCFuGrz2GlVmS9rKjyx/04IB5clc5XAJ8BZ6/OkqccI2OIpGrnpPSGFOvDYmzzwnOt
owvmG5RC/mMQfs2//p3Y1JKGe0KnoHlX9Q5SszbgTd8q8ns37EjdHiHiU0YwpRg2wYtZ1UyY7bOO
5MWV0VEP1nW3iFpWth9ZsOloqJ7ssHrD1gNNsUDDGjFQYapYhoqtjl8MyulWjTSgNKEftjtBINdq
EFBjyuIDx8KGmHSCJStEQVrPR+pWqs+tkFoQzr+qFeU9qgrr4mbryL0LgzPV7VhVpf72XGE1HVWv
DH4ioMmTAgkW2dPKYQgFjf8tFjj2i4JqpiydnluYuwhG6PaoIvcRi0lvKkqxFbkz2d3/UoJCfVu1
5yLFIE6Tmf50Nv93BnFuNciWTeuTL7OiqHAYbSMvS03tx1itQz1oC1pr7a949R4PAfHtMrNnkZDG
tgu5Kru5304OUcrWfNYRp2BJMteokvnvesV0pw6YU4zC3Giqq0vgrwPo3gX8bryICaVE6acaGPju
tF2Jn9jbMBEIbqcr0Ac7iqJEQqHQN/VGvw4pP5FYRhu3AjSwEC8NivuiBiCAPDuDMQeNe0OMq6gC
8Nf0GRvSE/5N5ggmeiC5DqIwkrxq45RBTRD4kC1HZLko4jIOiETLRutX/BXsOHXB5n+gQv+8KxYg
x3MumZkXOyhHrZMLRlrzGD60zXgPuCeOPr1FcJKMe8H4f3LOCven/BBnx9vrDVwr32PNlAZFNAne
G3HAUX2WQBz9k21PoNvd+zGVeY6mxQNiLhuKTITQ5nOXoxppZf3W8V6LfzElPw9PuOHw1jSGrL14
7gsTG4cEG1tL67AgTq3Ko+gOFntY5I3OkXS3b+aNrZKxY1HMnQmIKDPPqEmWnOgw7KhS2c3pi3O1
xd9DYov+wV983MJbMAA11gDQLae4PRZqkDIR4FSz+UbirksUjJ7ojRdyqblLz6MPC+cr/8uzE8zK
q9OdfoIkNuRWPky+KUaPItnKGX3varUOu4edFxevbar5gQGv5ozOjI7WIZ4A3zUcgLdgtP6Ihcpk
T0y+PQngPPNPRSr8/oZqnh1/sXLE2zq9WZi+pfxkNQFeSfDS9t5RIYLKHo7KQOeQncHBWUa+vQiv
SlM02PIocVCetpfBN7QtnEzmZG8m0QwJourtYZaAkRgYT5NCwPgY3m/KsfjU8hn59ujqE7NsZs7t
+9nEIZ8ciK80vUPjnynzRN+W8Rym9AS2fEpSXREtMeWJwbY61Dro0VZMj9aUQAxWsGqdgUjugX2q
ekF4u5jzKJYvzK0gqS1iX+adyxuQC2GO81nzy3nH031TggW2+lCJqeh56rfPJJqaoQffYWjOnPZB
V5bEb0uBFHc10zJ/dKTblQt45mwWBKnrI5cZhfOo/p5Z68DzxRIHFqzuRYuiFrmh/OTGo8T8Bp9O
eB9laNl0AuAmimiVRL/X9ss+xdBjC3808262/EIo+1kiSvG41SXTMeAXgxloNMbxtWiDfWG9PWSr
MkwNhbgshYnzLxP5nxZ6vNm7MeQv5UWIss9iCLNW4o5+MvKFeBbbljDq6orA54zVD87zvXMZcAUg
t1EExT+VcDbpJnz+1PmFTemqy105alS6CHBHwtboLRDIQpoqVEjbHfoZ32VCg6/6to1wbJibZraL
+yh2c12p9JVzVDmfVx+RWZzOQr8b85yKzr5iK2TlDlrV7kRIShV+fdmZRxGxBTzD+i/Y7vXJXNnZ
y1/UOGOFFB7/MtRuc5bD1Vir7kk65736hkJ6Axw5NWMN3+P0EK7weKolWdCOQRsgRECIlcVg531+
T0oLRXxHqM8WeeKuFmQ7m2aEqxeA+TVRYFIst+IhoEmwWpWO/D47fQYwoRU1TBjaVoK45B+nNNTh
A1zEDB4/MTsltzu73vaiw7O0EwzVpgzH5hK7zcOZm9wuKHawi0QVUS8N40YvZCohFsJDplFPUTDk
3FAlw8bGiqoLRGzsRwuUYzqF8+Qr8LhlXC/gf5nf28bA59x2RiHcwDQGAQw3YRuiqXvhxHU+aCY6
1X2dx4e0kD51g+XSAstBbpinxfBKzw4VDwBaQmKCExacb7mIJiOWifoQ6ZqV2Qyzh0/lRVuy8sdO
54/TEIPw7bQjUGeGRzAiJLHKR+bwcNpvJIva0FydHDuflwa6G4DUK4nBJBixDlO+SOrYY+MqUp0s
AAvztO9v5sMGFnY9XXejNUNtUNRuq5vS6X7UkCjjwfVHCSR945g60mBHIq43qzRl86iFFHYjEP0J
iJE5S2pregt2J+U1WMT+sCuLbHPtBd1ApVwYbBxkdsG4BFKz0A7NopbS6Z7465gzvI4HbjHMjWif
NqVb/tmm4YB71U7cxfZfKq4W9hCC56zm3T0s++KjPaQbGXwlg6C52rcItpeHIe38vTXejOM3BRAz
MefHU9jUAJnjhREJk2NnYfwQhnq7/h2kEreuYMysHKml9GleO9SMjTKj+xJnXO1NhzejzGZM5YFz
q0iTImF/D0/8GXkNFZyiVCcp+6vvgMy8pQ78ndTQhnt0x/1HuSfnJksbQjZZQVnsKucSoGDYwagE
qdq4WEGVdbJm0pIeEmVJWKwiGJ523LzcX5fh2iPoGPPB+sqOjWtn1ruszoyPIUKE+24cAFuc9m+B
fVyqAHSg78P1I8+RzOG09Qk7duIafZeNkCBnzXWOLu5uyYHNDaQL8fIrhztpD7BEx6XGmRW5efO0
lcQ8gjoTki9K4r0+J4/8bI4IKln+2Ie7q5wtXVmO89ajRQSzEGtVMxwfR1HKxUFhLAOmwqMEB2py
4PrrWbV7fCJqKKevRK3Qrjvgvg0Jn0rfPdSV//IIU4yN6r+IZqnkdRSOUUrvuyJH+pXpusvL1teO
3YlspsO4Q8EPh5BFn1ZP0hQYnMh6RuCYg3zJMx3dl9a9rVxEw/rTk1hvdYRBJPnLjmTu89J8CPaW
V3muYgl1CYS4dS33jz7rICFBCkJAl0eDyTrABCVCwArLNSRjflX/GxKanMWIG7P+1gI9RNNF5g/5
nha8yOr8h9+bYSoRMV0jvGFHjkAJE7zzsvUN6HPWUHvMtXmngCkll2BHKdIGJnNZHnd5zty3N6+V
4YK7a3I8eZZ79xM4CmrwJcrKa98F2PHFt/hieXT6zzHqFh0WyKLA/AGT5osCVuzO8bD4PdAdOTEX
YpPgcrDJQJosv0kQTO77od46zhO8FTtsmMbccu7BOXsssVrkrJABacuZxIQk/XOMix1zFKF+8crZ
VGa2Sau/xW9nuORA1Rm7m4VHEMRbU705tRxZtzdoa7LJVHbOmtkI7Vp29sIxL/bmC3znrLTp0eBL
LJupr5fBFPqdKBZ5lyxLiczfpOe8ADk0agPIJRqYRbUgYCpKEurASMheqYQ7Hq75JoHMQtuWw7qS
WwK7j88qW6ly9uyTzibRDOYb6FZXpl/Zf9fUCNWlhjjMCh+yUL9UNgH4o9+0/EayPDL84lfBNHLq
6kiHZgYRvhBnB7l8wElO2qdaPtePq2CdxzNvnQ3RJZx5X1NCJvyOXbeLbJ0XZVfIF5HTCRKQ2mPD
qKydLY6JjLn2e4uepHLdJf51lmwkj3mkToDtzrX5MNRkmluz/eQBzjhbxUpWNEK79+JBRh5hzGjN
hcsYqMQBSQocD19HR+1bpAL7lEX+odA5BegpXQnqK8IOfav+aIitxcpXNW0wy9fhqGqS8QAYjzaX
GTMbYwdZa3F4uYFlaHU5yDRvvXFq/XNa1FHK2o3vQxFmMH4Ua5Fn0BPAxSJRY2QTT9Eo6azqkxtI
8SRiOl8H5ys6CXeAN+M3iWRrQoSNVns5UW3D47IrXCtvuFea86zQ3Y6KJpfVk+sB8xHIxikU5rUc
g/snvheaVjkrLuDFxAfk3rbRYBansPRrgX1KcbnLLG4Ijgy4dj28PdZ5oFp8Y4td2I0Rn4z51fqo
CF81wGmUf7PYI6ZT9nPSn7heoqNz0csNgLuaUhhSPKy8BRgfZ3L4ONmL2uzGNq8iUBc2OOooc/68
VIPETC52QqtA/mpJ1bfl9lGHSnCWTW1t3nOidN0XVJ3MpWPpDrwTiSwrwYMkl0xnECWcDkemxvD5
uoqzVKROR9gyjqipfsvNHCDt5B8+duhJP2jaczgJladsUElurZx8xIQ0fLKuS9OalG9Uz36SfvRp
i8idzeX06khaECrVZ4ZQ7GG5aTyCfA9+xw3+OjdxrIZwoN2yv3079TTIVDMUDaarUYRaC1Ey/iJO
H8hVZBeFsmEkhKtiv/I8h1Dy9OvCXBr4exrNMomb0k9knEP3kf+ECLUCQhJxY90fLRWZBqhap/VH
GRkXYrjlc8c3DLynrfff9CNW2yycWb/1sFfxR57ts00tgYRfOvsfSoLuFbqGs1VNzRkng7k7eVfI
E9Kc93u1+Ln3XwQoHy7BursglayfH9yTkm6EAEfsdZXoWxaVjxV06uVIuP+X7En40ei1+y0bYiLq
/4HmoLJlrB+vCuwIt7Z/PGQLQuH33xPAjlyBssFDYd9Ck0Y16YjFLmv3LAihZHzhaCRYjltq52iA
9e+HzK2cRRyYakhjQkKCxxQAbTSJV++jSkoPnzQXeEDkNKkDCUiS7FJYN0HU2n+qw2aMUFoYWeRZ
ICay7KiRJe/p5z8nZ1M6IrgED1YkmJ/3A7O5dG7R6hKBQTXs6MbsCq6hJ4dnY/xlVXAZu+gITM0l
ADR/0FJW3FFcowB6GyTFTSyl/XQcB/MH305RiJUBZzVkTTNVfO6PxqJXZtxiAK4AgogkQBzfL43A
squc4qW+U79by6CEpPM2B2YVqa0mExHH8or4FC/4jNn7Up+O3Vk13m82ZYqRP3eIozkbxcKjH14c
57uY7UKFlbfmSBB9M1b51TDdIPU8hShKmTrUbGPlDi8dV9n0L3odSY8eKOt/j4jSIWIf5CwFyZn4
m7OE2pYDbRSWvmxnXSTV+J9UIu7I9J//L/uEZECcvitV9t5hfgqiJdLZanax1MQ2KKVvZJEE0U1w
DEjfUvWmQx2nmLTyIvblGbaeDIS6M9148i8ZoAqtzZ2tJHG/tKrLSHxE1rZCplSc7cNffqXRlJUO
IdlAlEiaZgml0YNQC/lPc6Yb2hLVwiP5dltscfAOQByrjCz2DD844QSSH19xLn48gX49YbTISLh6
itXcDX0WzpGYVsFhbNkHlk4kQ77VZo6nlZBMY2Bt+bS0a7Y30dpG2Z8fN9dpWD//O2ZvEuDxkA+Y
kUu607zSmEYC6dGLxmkcHfJcKh1HqOakspXzDz/xTs1W4fYAz8pP0DtTWxu00jEy3iRioibRTmKf
4b/49P1tRQVPdG7Hapxzzk57CmOD4JkZ1Wx/XWAZgK+cKL2PFaAOA5nk+C+JPaNccEIJt+OoxywB
+XaKdwOnotioEUrSrLdTT1fRlrdL/+p1KKWhojoW79hdatq/W3Kh3LNOuhRVwamWRknCE3VO2vFy
gEOIIh20C9nLgbmp1h1fXe05fnn+Jnfk/XjJpY2ebASoC9L584K32WJik2hxpHe+PQzzDbHeS2g3
PpxRRy7erba/Lysd48drYD7jFdypKeP3IjHxZtVgYDeeBfWmDclzVedo55NggigIjROpOcGupe7J
SSUCOaMPKvfWlMTfZdJjkdlpjrz1K3I0cISKNn4TFUvAb6zkfCjum85g4lMXAXT8iFpLsKG/vWkd
jGgmk7IkHx3UgDKYy2s5BFgVkF91bQ+UOCcPAxT7PAuadm77ufYxYBdasTsebB1RVKLtgMqxGQD9
pdiDZCAnZjpzHEpggqdXzFzK1yLm3F6hjGUjpewYXwQJFJKOZrnT2upD9f8fsKxHXYC/ckH8dl1C
wn2rkRMDrA9vJ0kK9JGQTKtBZYtj2I72cReMcxSpMB3gGALEvPoyZt5lh2n4xdUGGDVerls6t56s
7zShKronS+y5MeUIuvgvIg41wJcLG771T5irgTA9cDp8CpXST//LCahmbgWOXCBl5YNzAcEXZQK9
F+WQW8g7I0IQTvqnXfp00Sn0Zwl0ypMt86cDgnGdxbhwBANELrz2xHJmAkkROeDQeIEF9M8yUh84
1WjunIlOwYAEff4bab2XDWL+X9IyKBPk8Bzu8ZfuUclVvsDQ9N7eyH7QK41OYmdBxJu/VVP6rWCA
wW1Su0yWKIJIDmcfh/ZeXl32H2BjlhJlwbHIxlHQxLLElcfAMK+fBYu4zByYSVCqNQ/qyKH5UlLR
RQnHrYtxgLFfLbyb+nPJmD9R/0qe7I9G6LSNiqHzK2BDLBA3MGDa+RF9UNoHrhxhhVIIpY/z7lNS
k5z1YFozM8ImPYSoVemlgWp61/Gt+TJyVlsIZtni97kQaOhqZ5QEXlPhr6iQsu8YRzbMdxul6Olh
HwHYGRT2HLtoEvXJfX3WcIR8MFJq8FKDOCFpk9aCJgJfvNTlbcrXc50/XeS/NVWKymNfqa0dfBIO
B9NCPT1AzJHGfmAYyWMF31UttQ6yW2Tk1P2NBfE4464NTKOfSYV0cC576JhvbE9XU9ww8bA+tg6h
XZLspxHs2huwbV9dmkifnEQjVnJto6gZ+Kp81Fv+SKMxCm3KfngWaQju0wcFLkn5sS8182+7JMDO
vHi54Kapcznkh/fRWJCQMto23sMU9VhPPIcvc8iudjbMFgQzoDiq8geOd++5rgAqX7/wHYB1uy2k
pMjfXlrY1G1OyLhScsALMNVsOkah+ciDdBhUcd/6vwMrk+hdr1+L8IlWSyMmYZNhuFuX+2AYrD9O
fStYk+x+/lzpGfq9ZTCudgfqjuuLLmMLz2jVvAGJ5Dv6h7y7tS1QawxUOhcpt+od72Obu04xG3ya
DxPcQC6UgNrj7wOV3OlWKM69w6f5RI3bM8KJYPScF80wwp5dMVQhZFyCKrTZmKMJiUNDT6n/5lnG
qL45jb+OKqU0QNuF0kGvbJz+H7DRQFK2vlYwcxs8roBYydYswmvjSsyjKH9uVnOCfJiLmaGYSO7c
l9DtqrTLtQ9Qk7o3kTDYB4e6e18KkvXnuz0cstP0dk42TOlVNeYgNmXcWMPfva9jAq+ERv+SjidF
GF0K2ChrxflCmQt2q1g3E41OfN/iHXXslFeLfDWMyMmvq22aEpPW9jR0k9/fuXozpnsJ8rB9/kAr
kNoZTnclAgzk2PsE5voggA2GgKt07Pz1naBOEhmTUNyjhxUCqmt+XXS30UHLBwAoerhSXEUmNPkm
YzZooE1BUIoNRAlMweQtLAxmFHTfP9DosatyzcxnhAj08MxL6k/wTqHZ1qoHepY2a/UfKH5tMIAz
rg6I8Kqum3CquC7p7wUTaUC0Vqjd6Tkx6HnglDxLI9Te/DaEjWj6iaITtVQ+ryH7ya/US38vwME0
ccC0qlO9SB5+R+2JdsZKIAnEMEZmEwsTCDkSpOl/ANQ58izUzARnxXUdqq9/PMuyvATGXKMMndyg
4FeqAvE2SmIZHpO078hAcdYBoOBR8dRpIIJE2g2evDITyje1lrkcoJeTc6sAuTQ/uj7k0yZjq6BM
nUMbvE8uKcmalmFGtaUMYNHg4HjtrjBsvhOfXet9ei6jAsEVKYTGjei5Scd7zfH3KnDeeV+fERo/
HRZRV9aXWlvAA2vcRtDvVB6t6Q3zEbEIqeQ6VwtadH7FgB/s1VAjbuK5fhxm1ctzc6a3n1LXBWSw
GM64GrO7zpkeVs5w7FXeeT5OIGrkgYg+t4nmr6gjWi/wXD17etFpXAZD4gIuOoMoaOSaLfgWRlto
qFzRM6fSsiCXI/94r/7gzutc+3j2oceQqFavTExKAFsaLqlEVaTPY9QNY/9N30lNtlJuK7w6xvn6
eBGh/s5HNHuCx3Woxex2Cdqcu28ss0cGAdNKXS4xRDjEaQK/lB3wEwhGQRTVYnJRt1KRClWuVjHf
7XHmt09Nn1PK355QikHNdMt3JtfL6Og6Sh9tJErg0nC/QX9DwCX29LfxqgW2DDEcHgaSfM/bAqlu
e46NXlC0xVJXRZ0GIK6ch4ztv6pQlN/KKGhl0uM9PiN5f2qqTHdJiTQPtEXc0AQCPkbUrhi3gv2f
s0dFBuxGUpJvEJaKNXhvGAXm/eqhsKHEqW1llxTW+W6xNPvH6pLIyyad983U608fJ5QhiF5SwpMe
VF0TrpPg0gnUIuw3wjvvGvBXQzqy+d9UT4Em4XhT0S0SwnvA8XYbyC6rJ1R0Uh5kZBjKPP/KF5XC
Hy9HLqmjioMTBBU2sRJhIXRdtsdyMrmI+iTL4LVvuPGe1jR7qfo/H6wwHIgK+pJMo70eiAUZAhl+
7/7zjVNf8QEKSYJJStqXBTimjr6a/6eZH7PI3NNsf2a2JUvIdPFO9xluWZgk7YP8gXMp3dZ9WoT7
jOwL5hzAwBmqfZ52zlHHOq1jikxeQ1epJhTwVIw6hn/9LYv2laB8boTxohg+wYktrgCkSZ/9pVl5
JDIyUHF5BPgxFXUyrXfhffUJr/MyVKJfvFjXapOOqNqHXQ/3+McwFQvXLIpW2k8q5YbKpL/UYEP8
vSc7G1ezEDYk8UwbDitwAUW4aWi4SLUcvOTPXjkkm2PO0FqFJ8kGQWuXbgE9uRRm7NOlk86QLKt9
ePmFL6u/P5OXioBR8CxVTrHbDWVR+CExI6tdMxi51RqD0t297IE33zmpF1l78TamuWJeXP6h8dX2
A+kRYdo0x2USv1+j6MKTHyKYote9CnbQZYeGo/wbpBCoQXGg/sfGQwLOZrV9kE4kTkQxcX6iOWTl
4OB+dS2uVFH1lp6RiXuel++YRdm6fUUvw9QdezwLLFBkHC4C/ej2ZLW/8ogz0bkp98ojDGMPCgWS
IHXVbzMx3OtuJTKr2tfN1EbQZh7iygn/2FaBEBeiFnjPjSDO5s0gTsg8WH/SVqHZiaT/3Ic5/s4j
lg6paDt687u/G/S2B0QiVef6rMATJ+NvfD/cJUxn/NauCLycm84wpBX3Esd1E06lEO4+goHct3GL
fs9yVvPmg0NTMWU+1U7WCIdvnJGyo0epR1n48rbq6FRyOE+M93RyeApNKJIjlRcq7X+J+mui0aZS
PU96xXPFzTzsocqTiSbL4+PXordxYgxfnNcYJ01Y6JHY47VRQjohkm0YrL8erJnvFIwMeA/elzG3
ATSeuVEEcJBQFE4bizZ2zl7WrAxaIg30YBibHoaFYGPCa8zU20bGe9lsR2Wc2KIcuTZ0vrnQC/Xb
UBh4AK8FIDr381KW6ICNU29TgCzcP3kcF54OoIYghZwyuvwL4VXvXJ/ANYar1B6ofcpEovjF4UAQ
k46k04tMeBTHG7/x+QvZhsnMIpy/Fl44y4H5saaSzO92+gtSaxeNizpmSAaRhsU8yMHY8ttWahHl
JWmjWgHS+FEmr6AyYkZUBGywZJfdzV7fSeJnlDJG3noV2QTXcgAO7RqUFxShULEA1aPB4WDCrpRr
Vkm8mYZ/lrGiGeTkvogbbRaoJ4QHfiNSuVjbVlps8OcAy31VFQz9R709TpSTcQsXJfFC7iVpIF2N
f0Cx99Xm3UKwqfrdoVGNc/rvWOeb7iEPjur0vr4uh5dPTEykudZz8OzrzK8CYKSB4WDDoP3fRkfi
oAF/n1/b4wSR6aU5TGitFm9pktJFUJoI9275YOX0efsmzwrigb5P4SSqrLiN+47E1ZQOW24w6zdF
WykavbAveKNV03CHDAWt5bbHBzi5l5h1QkG/whdc1mYofAmezm/2YypRPPw0bGv7Xf8sdc/WtSM7
HGkyylvnk9u8pgzuJw7N3O9x33QOxNAQiQbOsPFggHv1plSxfTKNWHKDVGYiUEf49RLciAce1K7E
Ac3kBdbw2h4SlW/Gg5tN7Co0SZ+8gr2ZtKjZ7dlNcXZiMlHtHKYVpTwWjUT7ikSCqCS6F+Yf+Gxi
gouqmRpu2aaW4eqDba5PSYS4+sDy+jJmpion6Tq0mb5yhXUj6/tTEM6YgGTQI4PkdTiaIKa+yzgQ
gNSq9bhsO4vrzUjAHgofLTMnPsMrVaDBz9IzbiQy2tShUJOzbb9l8pLekk/u8dKSa4pae55+ZEnX
po9pnWxIaF1q3oj9UyJLj1K9KcaVSFQgNPC8QrrsaKitQ8K0gHNRjYryHLIZbF5WoGcNieE7YEfp
OX9rhaDG8zhTU5QTE0KWAHGlYHmwWMDLva7me0vN3RIavE4z91DzAP+JIqUgKZcvKMpfC4kPVFJt
doQzU2lseoPLRT24X55reB036xJVKm/r3AJmM3EzTlHzYWy7TKnYL6SghE1IuARYm7o9OKsctmvJ
P+YNwOibseoiAUx3r1SSb9cNCZoD4TKEy4pBGPgyHSCuF4KhJsCjJjI42IYEGiS8khDY0s6+RDOT
Ot224NU/y+Meol4ILpdIrazr6B/0LvhZ6RVyZLB9OtdkkqldKDCB2QxxT41HTkmt49ZdMHwGehR8
Tz0Fmk7VsT8pEzxbhJjJeae76Z3xVqluC5Obz74xV1/n5dAvkqqCBliO1xR5+96v8gOLrejUWeUb
vFBGO4lPGAfcLKDypM+W1uVtJF2w29BZ2GIXr19qdLQ6kxr4ahgrpM9loKGbHu7cJskqqoMX20sm
wmvBbKW1+xKtrP2zVUsVykKzaBmhESGttZYSJyvwBNBc+O+yFqzwkHj+2pz810KzLUFDizMYeP9c
cXBwlPVwqAMamNH8dJu47gHKqvZUAZfmDAsdUeLiebAtiO4oHuoJghTu81ZqiFN1nC+bTZLSBQBG
4sMZnRemDIQt7xR8EuHeeosCD/6UiLzQ4KD3eJf4B0pjoUX0i8fBQe+halI/LNyUq2gpUsHDJ8ad
d8v0p/WxwSmLiAHrWaehF5i2wHB9WPA4DXk/7E0/0bmUexALpfLYqp2nd3rYLtB0vAG9KONe4wt1
urQFUAwUiSulXHnwWHNv6CFOh/UL5g2YubdFtOF9I/XLsKaNbhC0w79I4GtCyP9aK2s8SBv7hqq3
I6xusCEM1GU7HusXmlLKGBrqQIcIMZjG8yPCmQa4V2NVrXSpQL24BkPAbGyIuSThRhg46tYY2L8N
rp1VicSP4P8hI9rUIx2H+wwh2SjGjpOUPGBXuJp65XvKBwdQIlil3sI7hBL0pvMWFzXt5hP7/HQi
o6MsFKcFqYBFKhu2xDF/bBuidE7jtggY547JsBqbgz0SWkTSFpaeFmeKfVTOCqzfxWVo5ud1U0dG
jRih90kDZAazhMSOhkx4TPexOyNcO+cWPYJpVqkUmsS5g5Ks9hWqgs38r5zHDbjizGwXeup1Zzbo
Zhob8eyMTzKJJ4XWs5reFZ3FXpWCtuO3m3kpOGEo/58GHY8pXnn84MudmJQiFjYB8ZatV3yklVWI
SVQpUPLQv7vIUIvcFJeBxqnEP6qP4LcgZEaqvLD1vdivXQJfrUYaYUjlPrXNXuoMPXFiV8V8kNut
NYyOAfzOc6Q/o/1djXxFFSs2O8ZFGuMyuGgTggJWYAIWdIeI2xE0ZJO+tM317tfzGRiPdGvGQAcz
ZzDWbxNMTQK9uBsGB22IGgjfFG5vTmjYha48yw/DFyOCVfkht/sZXSop1pk5A/wqqsxgJfPE0r3M
W3VbjR41CDqjJzPkZVLEai97sbgYOzWPRt8jFdmLMoi7G1ONDyyCrSAi6bib5Si7yJYvnE0huqAp
e7tryDPK0EHm2LFcxhSdWpuJ82sq23Nu7KMwSuDzMoSW+S31802nW/F7IcLJz2L1g6CxL7PTJm35
BAmw/wQDEaORZdHoEBtRcChYuDJkJd2nVeT3oqW8xKFKoba5Hvzohc34QkpumDdOU/uu4HZ71j0s
mwn8QvFYueoK6gkIrzLOUjLsRkpsbNMFw0ATI/pBydLgTH2j3Twd9xwWYBOY5sQ+kK04kahdkIDk
QKyH+3jXZFLRnlGVP3jBP2M50KnOFxQyrZJ7ITG25nBsKQyRRnUzi2FsUJbJk4ZZH/ZMRH8nRRTU
KtVosLfjzJBKhc48sD4njNUiPVNM2R42qWoTsXlD5CH7bRL23IJHVTsjBEsIEr+7y/qozk93bPct
cORzLpKpYw0mA9/SdOsMXSiUyRWI4nxV9T25F3qSpJC3iwpe3CpwOsTjYmASS+VeuHUkqAms5t2z
SQ24yyBSaxv3nmIfNA+0HjtTHJ1dRJdefY+CEGCPvCjOChcXB63Qm0sTpE2lpUn6Xpj4RbDjuUdD
k5UFLhyHkrKf5aI8IIdNrpxUEYh9s/gDymDZ5JjavERAezApuksmjVi73pphFQjyq2wUV1EkFkGj
pqzb7cd2zR43TeBjeGHH6yh8pBksetKP0RI6estg/MnNHFLybTWbutDNw6wLae9a+JdtLlREuSZ1
ZiskWBUFbprBJB/TQyv3pU3oEv9aufBV2LH6kFnaiWBMn2KTKWk/NDNNih+jAfJIkRzibgqIiSOK
lqYmxpNAy/Q7xCOeVqzykZls12SwYTdOZOiF/QbotV/zG+qiGs9gL1oECm8Qs9Ad9V39MQyBlKlO
Spc1zAZTU9/dLD4ZM8lFg+9DmErHtAVsxeAId7QqPmB3nIqKbvPPuznUju7FSMzB6/25btH7MH7L
LKfM8ijhYOIq5MsRvGmSrwPp8UBi0fIcYe7hnVJJhnGqjP7cem5zv5DEQ2HSeN24e2TGkJbnBhZx
VDBJorWiUsciqAHCg6DoH8GTQkS1jo7fnpCqz4oMWR4Dh5EOXWnzKwmzVgsCmTaucY24Ltourc4/
/CPGhbP6ARbPaDGLQPYApo8GfQOxiwrsKpWMQsCZIYuOLulXshJ65RcHDBbRUFqJsdDNGzaYIppl
/cZq3NCntbG7WxpE5FhQnDOf6U8AtKtLsQgyxRKg4bVKczII2rBAvG66UMWDuq0VBODrm1Pjdknx
enIBXDMqmjAequ3Ebbcj8IM/LUxYfBglWD7QNpra6uguo0TTd85qjq+hDRIFRV4isUnar5fBH7zq
p47YL2nK0cCEwCD3o4WP5sYiy1L5/D3OmCnP6XDkcpTanIoDwRbt9Fi5IJ+BJuDMgkgkammu24xJ
OSopejVNUa6lNwEPvrrMRcrGknerxo6u6o2x0F2wC3wks1Ztt8nioAvfS9PUmuN8Ts0VuM7nN+pY
KIBSqH1zsSgeZ+/aR7LMqLDRfFj9HNq80v97jkwASghns6bpIVXq07nNMInObJ4DmT+5qCKBv4Cc
/vnrdwWBZmcVaq+Y6U4hF3Uq2ivqbpvstgrvDuFjCQLkwTZVmMdYxoHwkOP5jG209a9RZIDsTJPP
yd88BX84Yp+GP+eciBgC4fO+lgLX5syu45lQ3QAu9czORyVB/KX0iGIUQ/xecSZWhBkFrDD2WS1c
kqpznbGTdqzJMRT6UxIhtnOPd3sPBvkQphlue/vEHVnXUQxZM6xcrqta/GV/TtK+U9Noe8Ka2Pit
cI410FySGp4nUC+bLIbD3QO+sH8L++D8EhmjkQb0s6Pv1aWlofgy8pLbX/M6Gi7KAQn7K7ehWdBC
4xE97ZGYeZGn2zQ4Ox2RB99pRX30eawCZ03Q7qFLmcL9yN6UxXP/JJ1Bmi3sDOoLnwVsXNsq8W4s
ogZ7YjpKVfSpB6gAarc8qFZ/o07QXyxAjvNylNoxcMcdjk8/hPEP+ry6PE9/MW0Q7Qe8iPtvlHCQ
EBHitS7E1gk2TGDewVo8VTekv8xqU5hd6KIkTA4xO+G9t4gE64O6SzFq7/E35IMvBqlSerMXkE2g
2N0Vu0EOkR57Nekc5IR5FuFwKW1ASA3LkplUjeDX4r9ugLqwJfr7TeKS8BaANl/ITYsUqz/xwR1m
qssdPaDVZzpLDHTN7vqPUDGDDCWHV/U9IP+IVpqUgF4x1SdDregVlDMR+CVUavbs2NSIvaD9IpNI
9wp9opHsF9iH484upIwyImFNfW99mnZhFseHA0s9hRxxiDmuFExJ6rSQxfmLUbn+blkHE1LivE1E
34MqbpzZJWo6eZsVCuSxIKqpqhULRPCbBTzemMZeprlq2RMNn3sCqmOTfsxLMebjUNkAXDSjDgJk
Byod66LcCSxAoRWDk8/SAOT4HZkb0f4FiO+jhtcWuWfbNS/6z0xcC6+7pxam92i82b28ydXxhJR2
fwhiWq/EcJiZIrAaDmXEjWVQKo7+tLklYI/BPdpB294MAgrOECREQ1Q+4hoGu9AIzK6XtlS13eHl
duX3BeWxmXAO9yguwQsPSBqCKUX30e/+FeoTWlNXzCXM5FItmGaX2KLcZYh2QFOboHIj85LL4ckA
K0ackVOpVIE4w8GmvjMSIS4O9ZU0Er8+iLrxoEvI5mpHxeE7XvlyvJWoaHecr7eiHR8cHac4+nZ9
YIusJI8y72w7hjsz51fkvCcRc+pMAhr7TOpLLg4uILDvk8iHSOZmbvmsuvtgBi1T//cm0J5rug6h
bSQ3jo0yjuniYv73Oys4ibgBtNdbrWSGTpefjvH5D7+ASiM7oJxb/UzLSQUw8G4IPI2dNQHhj5W5
C2JbnAMWGysQFolMQtg3oXi2lOwS40BzFtrKWNivjEZPECWhR+cFEczR6tSTYGUxKdF+Q2hu9nQK
3AxB3/qwBlkN0b3DLTWmKggW5BySO2c6+iDXECXDClFjOuQ7h0h5Jw4BSxomR4/PvPDkeJnbj1MX
549vwqcarUXRYDdnby84Tf79DrxX2PXicbL4BG5DaGCdh4cRHuA1rCx5ke2drzbx8MIQypApPU11
ihQ/O6Mus1xhRSqRLFlj4MFTeYk8XBgITOJAm0WwkjegIwXR+KVcW1Lm3igl+Ze7QZr8rL7s75g/
kWN7WmQlAccfrGlplvDak4ji9NvIEDx/nGbec7sl/kqIuuK+80j7xkfVqYPwndo4aHF6LbdKHfV2
S9ZPs8/IrnJs0nHymaBmFrvMmlv3qc0doAF02n+aOQHSV+VcrFtjuwcC1Dz1rc4TdnIC8sf6Ie/l
K0v8V82fOell5Kt//bjsma0SfM5ObPUrR29Sj1jCc4inOYwwS88O0GTwqnfmCN1r+iNbkaoBFlXO
eTQJ+Z+WUzHXKFK6So3pnyHOdRQMDGepDXtHzoy9BBusW226juDAOmwtYLOifnxoTyp3OvvmJe/d
3sHSSBO/WDlAYwJehhQjUCQvaekWfShoQtQNjYgau1RTbELMsGmEMNhGhi2TbhgR+05fi5P/SHlU
ROPGmO4D67RGyaH7/hYHSaQTzUHmQOFDq+uZvHs3Dj73UyQnPSGNNRisVHDXNmFjoe89vUq4k551
E67dIrzbNyrW1gWFioVpZMEzmOpiXq0G/2gF7/EfWeeVKMCX95/o0T/gLqgUISrmVqG5Ch9GsdeA
1fCENtt6w8XTncpFW49QT/z+YoYGhEyv9Y0RQFlbFlrRtXP04FKLghYXMxQs67vORvX3aroumW/j
gUcni20r5uXT5Mv1jHcpi5myMS/cFwX2vafY5ommhPkWjQLAvMULdvu257xrugVQ2UrtHtpraPYn
1KxfR36FZwvwpew4ygGPpmRAa0pzfMo3g/pYZBW7hJ410TZ6SdhWDGECKYv18qiNkm2BMfvCJ4hT
I3nF0ihYhL7a1JKaoYGeYbaWiZO2AmwEaL7/bPE7DuQfRCdTmtOcgOZDlZfnwanCwjAQULvVxrL9
0MH21x3ia+dZFTukBoMr5KkS7GvwrdyQG6tf+SG3iaWpiOssbIcyxjcENN1WjpIZMKSP8Xla98W5
a5G2LJf2fImP2IVOt8OywWNdX89TU8c0+9P0aDk3yCCh9DrADneSCZLTCUNaKQTDKikLQBxU5UK/
601cyAafip8C5Do+CkLZNCehEtLIoF+Hfiwp203XHVtQQLvgU6VqxL3ukw7VYmPsiOK/E7ZjdM36
Fqpoy/U+ScfjoRypx0iiz0BM/9iYwQBABiRJKOd2G3IIm0rHGvi22jGoyzKDrVQzUml2+0Mz523W
2PBSr+mjt+UcuHOyO1kuZ8zOcrm4IKK8FxA/3X0aikExpCFe/BpTGjgjY95/S62YwoB3eKQ+RpCr
gpwajSgeiTzbOuhnB88wB7XC2D3jh0+w9ZjhDx7Q4CMUXTckSNUeljNhVtt9opC9EVFh75dt154e
v2fvLWU5cfqa3H+Sch5CeLoONGfcx30ZxMIGTj6qPXvsy0e4gcw8oZ4s/qVM0RoVEvMxI7S/KnJE
WIDd21cVUxkhkjJBTYX9/t05E9ADJ7Ap+PsXYGsUmq8skiuRShz8GhDHKu3aYCj0LrQo65nngDkD
ozLI2t2WKaNToOgB3oZH3xsTIKHrhmBOSlridMeilhfzxzSoWgFiF3GFgpXIQOzdnJwvPhyI+Ai3
AFx+o6pULgepjj30O9RvDYw0HaPkiFsj3lgJH9XDxcuhazjB7+2yUXcWHwoka0EGCqAtZ3sq0EIW
qrI7uJ3x8/BRZFgAhf3NJPU9R0PlsBbOJ5GxF3RyNhX6DhFSbHmOueUs8XNjgwNCrH5HchHItq1I
aT/nmRXiBPpqxoFy0LgJ0e1ROIVLzzFydxeRDVBdxqzqgWcosHxPSJBLds4wRzIo7paT3xM+2pJd
dAhIFZs2LL3OmKzoaZsFXvwESfWA/2EvsNy0qHsRfVPkVjXxUKZwdqTB5IfIxTL3WUu9bCxlToVh
YZkQOOyhguR+OlDjd9eXqHcuza8LxHYeAIfuHvw4KXMlyXA/D8lGPZzfjIIBFFt/4eSSUR6h3E87
SSsKNcP6W60kYS6Vu96RmPbQ/32+2fXLrXsheHeAYLe0Rwx+1Gi02w5/lT1KEENmbaG0R0fcLzxR
vHY342wb16pdrtAHzI6THnXbzLgRxzznXZ5PgZyvk5pijcCvmHj7etWrVs+K7c4BqcWT5a3bV6ao
kfyKrGg5E6exNhbXURQmgReaDqiOKn6kueyWoNgvkhaT1XdN65Cif9TGhfW4Vjo9MdZEnGZwhIGB
lUFTkct2vMq+VjFqBekCPmhvpnDebCSgA+Uh6vZUNuHEPsMLt2VxVTI5BzzgqQCM7oddqT1sP2ol
0t/0lMOcTnTu9UO09/FfQSpzpZRMXDqPGPH567GKBMFBEW476TP7y6QQnvKwAlSWfklj4oMPtDca
0GQyCKDk0dTDDZpOCteQldgz6aNuNYupfh9v4lLWuSYSHAJzTn/7tmoqx3P9kHtTVq00DW5c97Im
mrz0xuCkMoPNSMHLdoeU0gwvbR+NDN1GBCU+ftuCYdDx3ZredQjwQqujJZThbqlXelxR3UeYx3na
6qKrH3tu1vgcyCcA8F+pXCQMBhkOECXZDODkHgwLSdZaLyo/u5je2ATGpxaFmpwkbeO9vRe0y00e
SrKdFCO7RGnnutDCCKckYrNTk7+Z/x+sIDrAE3Pv8Yd/uEo3zFmpp4qCvKKj10k4fV+9ibJSwrbo
rCBMwl6Ns4hW4zzodv7zycc8oxO2gRRJb+EImun6UBjc/xWEmbm1EA5CwdJtP3Zm8v06WUsBWG4o
9CrHDhfPYBvZeCoBE/DhpeSxPu+mN36PfqDCH/UeCBK1b/FYWqqZRK3hu+XcLnxWF1ZLuNnyN0wL
Y3i+E1gMMGMMkAWMfsfulGpbN2+UnsDo9qAMYkmQSOMnBsdmqfQybK0gVYenZC3OoFb6UIl3+vAE
ktdCgYlQpsY2+914sjXnDVLWGGBOUjPcSx+uzQU2gzR/XGk0S6uCMsbOyM0cRxQjkk8C18aW+6MK
JUBvwWxfq+pud4a+e0ZmDjtwb7wDgqAN1c68M0p0EtAQH9OVPnK9EKFR/8m5QViDVv0HthcBa7y7
lp/kTgZ/ekR4Yi64C9km5zVzvlONBtoh/0uxzijhIT34nFJyepJqzJliN7ds9ZCUoIxzzBM8Qhp0
wnQIZ0GS4+pvxZppSyD95wLQlABcxmufx9xYn+HeJ1X5fDP9D9KtwOitRt2b+gIbyt9OET2zpkro
UYjePmCShMqRBjkcFxwnjiEODqa2O9wB4i17AWKO6GoGiILq3LBK4/IeSuU1KLPYU2rYMvxoaS3k
hshuVwkRnL8XzXKf88la72XDvnV1ioc1y1df67CKrL7nq0Sxe4ZS70eUBAnG2RJV2xl73LHgQ/wf
sdfjlKM8fHgp/TIA8QMZ8UikXthpNEEQllc4CuRIWR1OYvJqof9uRJt/ey/cA/bRiGK8twTd0QvU
lIn00Gl55GfnixTWBFPdPFi8bZoLC2EHGTRF05XerkJJkVBTL1VxTkYY1RwUFWZtm4nuBFlIdTLY
FMzDrIw92/OuexcaKKt7f7rabeIJm4Y/NLYfDqjmYN1XbWfvQARdIygcudnqwzt5YmTmgWWXeU8q
hKAzqIeph07ifHqO0dWWO545hgoe8mLJjqE9C6dgu3PyuNJ2cpJiwoX/bBF6dQDG30ypThk13J2z
6YtTw2cW5OASTDJ2DLZwRntHjwJnzkqQwl1IHsLYedMVexMGwvkL1S3jjM6hu9TEQzpx0/A5DrTB
z5656GFPPGB5chsgOFOVR0JWXd2xjllliuP4MUzGd2LYmLDDAr/1EGspwFnInpjlEtwIGpZBQHmI
/mXt/71VFoHKo1wTHDmpG/j1z41e/D61k7gd4vJOr874F/na5pi344krRBo+eEGU0oKTovOeccGL
TIZfdDatMWifzVl1J/zjCidLNmcbPt4+2JpotE4THTQQjWxBoEM5BuM9TzVsN5DCxZ/ZJggkn64t
2QBBoGCdb98D4hvE/gBO6yyv7VbVj9qT48TCafUpe2g9SUnZm7DSEPDNCX5lkjMb51IsKiZbeBXz
S9K8vtvJS8rW7WR3SLidVba91xtJVgZebYRZEhvki/A1/ube38XkjD6CXXxEIDyU1P4jwPxN/KHA
O9Kd6Tc40c0JoVzKLYhT+wWUzAhQybp5l6fpiejxTZeMGVH7SQZjayj2SXeeQkhpwkHW907//z8F
tyKfHbCcjg5t26g5WoStgJrEqUFrvGbD/f6Bqyvcl6HX8E1zDztZDXciQF4f9cHCNWfHepcDm9Zv
5x/WuYKiUAEdzDEP63vKfAf2ZyRC96uVMOPy12AN70ZKKWVLppNR3ZJwAHb+31fSAJyaYRqswqG6
Cjv3w/Iz4tG26YtRo+iIM/g+W+ZwGYSwzTLqQyur6GF+yvmEbwCT+P+tpWRmu3yiG0PrH/ec6ndC
FoH+zSwWEFYkEm89RAQQFS/h001jb4CfYZD5Co7R1dvUbYhMQsFoovoeMp/xK9yEMx97WQy1fq/L
wnHNhcUghQ7by1pj+fKARyBoMCM9DGK/zCbYhLnyK26RHuG7w2mj9Os/hfSlUzgBQ/0ktRv9icnf
mIee4jUzxDhgDzLcmSLo9LCbtXUGKHCW6vBkHLdqqUHJQO2KYZCUjyJUHlmgWUnysRpynnnOljv9
YDcbg+XBQVUV0qP3E16Kj0F8xXAdURDr7qApSglgxoTmQADCT4S8aKK7d34LZPNMJopuFuTpGaRp
YKaFRQDcYGF91x0yahG+V8Z3ZGH9NKeg541zYfLF/8NgGgt3VKaBwuAiMT2OHHqL6iwNl4hcyRLt
ViWpgPjmN0nQz8/i6f9FSe4HGkCG9fBjjZMe8sIkxTdYteiaAkgL9lORxtRqia7RyzM3XZqJCq0j
Hpj76ruGR0NTZYWqSh6Ca/bACff9qS7LI0j/5TV0Ztq5DqJ2NAFr32nIT4Ca4sjC1jj+Q5KMP5TD
yM1n4hQsvYk+ETvOkFCS6q344aVeK7LvT0vcyVsKgmA+KNrZOy3Un/DV2teSLZEv+sdJQ97RyPnk
GxtzG/EdBMzqFB7pGaPhPMjaPc/OnxSXk0e9sparjvu8T7/L6PtXcVqWAN8RKE5Vqaq+5tFQMUJB
rkrSv7ctGuECq1wk7SsQ87MW4bc0rHoWmAN0aJbNBqIGsUBYoyaBmxsuZ3fSmwUIosvWNcmBQkB7
BZT9noPIPfKnfbUdfY4q5qZV1mXYywMZ6+WW6RQW6TiVuX2WpWF9EvRANcktpOhRbPi2paXKEar8
f24p0VrZ6YgsWpBjkHV8Gwo4vVHyKYCnU81J1aHzQ+Fx7aN52Mq04y3rpRWqUYbAnd55THdRDwza
c2rPM7GMIy29iFYIPRM9OjF7a3LFi2yfIKlEg+u1IIawXJJX3YDhmpMc5dF8qGjDuR4RUH9EZ5y9
mgtasCf273/OO0vC37KzgarTc+M7nkyRcNhqrxjJ/e7lYyKAsJDbzlgQa5fP5umNoLJyJ2W5spC4
szqpcPHPiP9kkPKF/TO4dKGGi9DQ1lAAZBXv1xdSUdg6w+C13a9fN70R7n6mT6J9J4Uuys9agtQQ
0oxWHZJYlPKkk1Wz9s5VtKp1sU3iJ2Ro8Kx9pjnleqZ8uzWsE+riljVspHvm6G+15Sja7/smC8Ol
k/jqd8s4fhDUDU8w8odPVmKXNkCtNHYxPmuAvMjsOCcxqDkM7W4tJcTP0iYWUlh6hropIojYeTab
hZQJ9tC11cNGGAGp6aWz6jBhspRPniNSHIEYHbjhw/l2R9LDhIQBIzPNCUUR54016Xdmb7bwYgoj
cGVTR7XJe+snJ0kFtxekN4aXcO0PuSFNiq3suQbYaXXzb17+wqbZUeisy3kr6i39cEBYqa5Liitu
vN42td77ujTqFi7DN6j8tezoXNT3SQvI7u3Mfe8H/SCtTrAxjsfNnNyXHOU/EMqGj0OXYVxCQmPK
PQEXoZ7vh7nLHvXU+HQNsX3Ey0ON+JOSSeF3yFMOUHzhtTu0Jbpgd4vM3rFw1sWkJ/PzIl0tYE3Y
FOKbXjBl3dE8jjl4ldUiknZaOLdIi45J6GAQW9WYQdQSTcl2ZeelcntfMenmDWhhOM9I9s/fIq7w
w9ter0owfI3xrMX1IE3q9G9L83EUuACacFJKAWwi1WIl+zUe2hXbzWFR5qcf+/P8fbXxE+kpSjtq
mj+EmqE45PDrnN/5vKfbJxC2i7kTU4gNUCdJiw/jHLG6oaEqpGHw6wh4QNT936gBovNhEUTT53Jk
I+fx8xOQzRFVgkX/8T8n5vn+3F1G0dh/9GkZEfDb0Yorw+Fla0iP/FWWHzoruCfBgCdmKHUenvHh
DvfZsN4tz1hdNmYK+vMXHLKndroZOyiOOZIxUMHoUSP6anYOKllk86T9XiIw+j/rZFXiyKG4rb/n
ASAFUsnXn0d8jx27rv/S/q3mZeItmF0WIdMwOCgF/Oo0TRjefdeLY2w5MhbjqDamtz+2W4AorOJT
Uawiq+9x2bNSTqu3eD6n+aam2kVEfTCdM34w9tuCNpxZsbZpRg9WbpejK7oThC3g1Oo/786oJa/w
/2LzL6q+o+mnKhPypobI6xAaGuxvUa187Evknmzots6naDH85MexAfv0GX/Iluk5jA5fEUx0cV6Z
DRnbNisywiF/03PXuxYVCeGH5EVd5CM2ZCTOs9cbZIWO52OvAv+lj3WKelvHa/ej8tCTSgEEz0o6
zOQDSq1UaAVJwNGI7Lv3WSY6CgzXku1FkHSobn49lhSfJbEUw4MObUkcoCf7JOHvGFtPYHYrYm7A
QVd16e0eTXt3Ih/EgZhCkDW26XIrH8iN1UQNBMs4gjdpZT0rQPm7xe+FziAF6xsud/cSWVLsj34j
di/bbeOcgYPhUwpdSE/a5qFrQcQHfF9jZghGT4vwsVMjF7TflCyXM4kh2BKn0ScdIA3qc4B7vomP
YhcyDZZvAuF7NgoH1UMhZyW1fDTbigFilFqs0teiPOlI2hTCKs/0wlrkFWM5y3g4LQsAqHEwYZTn
M2KOO2C8LNbr1od3wqXejQPSe9JyHWLu/aAe2r6b+Bd2M54sKHajGf6Us4E4huLXN28HG9366MBe
1VQBGrQxR1cHN/p+Hdne6Kv1Fa9g+L/yPfnkG94QoxVODVwfZGyJ6OdKuybvRPUSqum5CvYHxW5y
PCLSs78jHTv0stGP9yTzJsqOACww6vzxtKtCmQ/CYLs1JDcAPl8mIlz5eFMBbYEgzArivoaEYMzY
nFfL7WJb/YCI2QPE3RjTdeKZytt4e8YpDkCvFy49TCAkc+WJGObSkko5ee+oh/CRqXvJnOSeogdu
nhtpwb9gv7dAyYXYuMOwFDSrzqaR/5NXS3QAT+GvASCcNgRlnybKogHI/BL3KjP03smKD606gFuv
+TjxVQuJB4PCaLnwGXMlFJ2QagM7iuOTZHv7vqdFfQu3WU4qB/HM1GnFN3uLiT2gTyiF3nnSS/Et
/7X5Xhyqi8weMJ3ITkU+0S+bqAk/c0c26CARvZw65L+kwC50ruRANKwZUuDkPq7TxHNlyaqNZvpB
QTd3xVdG9c0SsJ1ETPTgMyxn8z2MZqWcWE+fJcUeL+5vhjiJQeFj9N47KmpfB8NRmec8HUrNdsss
z3smQ4/P+04EmCq0xYfVLkD7Emy0MhaVWYdzgFnIskoamsgo1MaNfVQVpbAh6Jlk3+WJniQncWpz
PLTZh9BIbPtOIy1HNTjZpsckQsi5adGQN1aBOH1U5C0sWHGIAw36A8HnqiteFVnRqZLUsboAOL1y
bBomB35XbXCv7lpiNr6gHxtu9O3cObHEOxhiO568QmN3x7RGKBCmdnPL9Vw17MOEUMhcWIjzfibM
l9Yz57kZmKCFLN9DDMvajzoabaNyoAOOC1lgl2hZADN9tMaVmjKXNOwiFmythcC2CYigf/W4pA3A
KAST4HVUdAm3jhDyuIcyt3HM3/UUF9sdtqG/lA0ESxgmNauQxkjacm9xreeREbul4tCBJVmDCNwT
Ztv3JqDY+OKV6EOJP1Jk877+b1BVimb04xkAJ/GE5Vycz/drMVerjB7qT1IRfrikOZ1H09dLlDC/
GoT5Olj3gpsVWRYS6L4YfsjzxytmcoyXk4tJCGGNoiZoRVQHdrWLnx6rmdWbVF6yqTOP5JUpXofk
iMf+LcsTPobEJdf9y7NOZ3ctHAAK9qYTksEmXFbiggPnC+av3DzGPwzs4b4gU23MGRBgx8sY5VEw
Jwji/H/lBa6j5NAq1mj9IZNB+FC7zen3OD2giuBCqUTr3TK9rwp8DbOhtEfdw6VQFN8LUrrSOfqS
nRbR7EmSkbsk1xEiLvOK8tPCMFy+w6wP4yVnbj0MZUsMHm1+B7tHlbNRX0uC5bV+fpL9Hb/ScrON
SwZNes7vFlE00qEhaIdbKI8bIq7Vvq/BB0sXnkkZAc3XZ/nQUBThV5Chrsp0CN/Cbn19Jxu8Zi2l
8yne/kI7/0foiu0zHeA4G8lbLignoD/NxgAmfQcX8Agh8Dr+z7uDvZQHNMHmn23QPFxMow99BMPn
mVQvi2lQlnWYqZPc2TMW+0zhDFlOPPUWtyG2OLfEzsaH4NkuPSbubEQv3/kY2vJKwG8PLo2VaeQo
w99A/4Ypo8wBndrhkQrBCtycl/WGPS+HjimNu8tw4I+DaRrTHwE2Ak8pnYTUH5b7ZZYX3KbkF+B8
unayCe8iS3GutOHxGoGHNL3Hk5GKTQCQP3gpDH0FI8wTb18W9j5yb+mxE2iRouq27CcTHYTMKfeg
ad/I1/UQl1MxnYMr+pmVKbHjcoU+Lt5SDk8zzbf/8jQYc7DAv0MfTMud2ryljgf4lCMamVrL+qR3
VA7W3li/jlx7eyIXFG+gxsyDzJFLwMsu7yCauQHgZlzy0m68HdY5rffNDnQSf4bpC1PWyVp0LZuy
Hm6udbxAah/kq7tG/E3YL+A7n9G5nQ0cKVF3oQT0FFJYsFa931RaofTwwGSGcxxItsL8WC9+ki1T
0M7QPK72rK+x7QRg9dwy3Ky6vTeUg+AQxYasvm6BxtKCZ+nhb0Q++m2bNPui5erc7KMZphwhS6+L
jk2x0tL/5LK32QHMCHt6UkG7PR1QlYVJMcj1nx0y0+z0cORaNznFLLx48QrubuW89IUdX9fREqVQ
37maE8QMgNx9mod/g2g9eiprpdP5sHwqA1R2YN0PYn8afU86Drc/l9bMLG8r75Do6Rf0+ZLlZoZw
KlLlbhpbYDn2sJcMXU9TXR3M3LL7CGB6dIzwa9RPedCKe9Ey+ZJrIscAPyO4ZIyAZJc99uzA5+dI
ciF3y7mtqbOnK5pTcGZKOMtvbIerEFGJzVyoxeV30g4CXx/p8TdkaZE9EJbsaqlQ/BnjOvesmkXo
HjZupcwiI3QGwOncuCgaJTvfAxoBiqKx8AmTSbu3MHm305BNJwRY9dH+z46lkWpCIS+OJ8y2VT1I
kYAvLOrWj7hXG0OzbbdlJ6JP3NorXomeA9vmNUJtJojsRTM+rm5UCDRx5pZPq6erpePuppLOW7dZ
fmh3Tgi7I7mIHxSl9e0znycZKq3+NPvDSPJ3XHM3OLjN98c7MBoMJLX/xp+JRxC/iDdKy5j+ot4K
+5JBu2u1EQp5NvUgNjY3Lg3+rKgvCtapv/isCXOzlKshaneaTChVhK+jy/SDAYszKO8pwUeOkFVZ
Rk7Yq3Rj4oH6Yl6pV6C6KV/EqJU0qzL3QL2gGdmN6PJKZpEGNvoHVgUb5HSnvSW6P1NgZEk9LJyq
Am99M2TCtxY5i8AKdnJopw38j+TdON2rLq4lVIZOBc72poYwRRfS1LCEAvPDUzByM+cosd5w3ZLA
Hkgx6n/7IeoTNJQBXFUbBWLE9DhD8L8m9LivbF0WskrLhHey8GoiPsHOKCkugZfLyV+BuMj+aUG7
5UB/vZJkxj0L1WS/O72zW/IP0Sbu/3xLs6+ACaSButscPskoST7Q+UHhv1QAm/UvDKPrcGZufYzi
7H4ituLGKEkcTlYTRWisrAsZQ1gIs/sdS9nE0vzTDsFXfvoLWhCBA3O6n6YuNcOWWltDv3+nxJLs
SLs3jBMRfvAJE3fDBUcmgjX9/B4XRcobbFshgmWfg+DsqeHb47Gy3uWzlmGBq+uyiA1sjv/ZFENx
vxJcPZsjWjO0QacozNdsvpdH2ZGesRUldejm6tbJbowPoeoB1G75YGooBbKNJi/X5htv0ZiXkpsM
sYJ0C0A1rAStuxMzIC/AMQXZR3FGqf48L0Bm+4C02wEaL7NsHcowAth1ab6jB+2s9MmMCugzUonz
9cN810wpEpF+n7eOTy23PV2TUVSbB7HnaG3HIAjaI/H9FLvnt5omothbnUVRt2zvf+YKU2FJ2YIi
v+BqlMvmkZnjcfc9gBsPTw9Jqhm7fJozJ90GV0AOyQ51ZXDt2dOnLb/MY8EZdJEzQHKOWjTsx7jD
ysEgtkgP08zkWUizIkNr6ksQmCsXxXKZKWYooZMUcb9qBtCh5X2uNVqH8b9/S37pdgrA4xp3cC+m
UheX2HszInNe3l3gcUsl4oFeI8WLf7H2nSCDvvcVKhF9wbjVy+zLSuhPpz/x8RD7D10XeP9SXhaO
ohiUZ2DGuwwrve2FtYavX3Y91sN/FtQODmrnTjwAJT6VbW7DUFjoO6pyTqCbbGhyInl3s1NUNaKg
5ofuapgwZXKJAef/6xMXYOi+BKlCeEtNlc44Z71LwjSeq8JQMBdlvYlQBb5GzYX7ONXa4AcSknEn
N7ubg24oXUPR6OLCnuVzfeMFvIZAiiqoB3NlizsgPaDhW0VJKV5f4ccUHVtFD4CWwOzRDlgF2A49
99MSrBcUh3wW8IUch5GEvhdV2iBlZi0CSh59Qhjnyxa1g2muIlSmB0+cjzckKRaH3156MPU9isZN
ORsZ4AO7FVXEvhe5pXGUC+Vx9WNCFpDd5X7uLLFJTSxOaCM4kf8I3r6zS3wJVZkxJh/6fK2EPjfO
CDI5e7CdD1bYAifQD7no8oCekIgvsRVcOhKMaPIysf90fGn9caXy9iA6/nREQpqKaYFdd0XZ1h7H
J3PQmxQp76+J7TQiTHp1G7ZTrBfpEUJWS00zHCedaXZrrOehhMLt2Ro=
`protect end_protected

