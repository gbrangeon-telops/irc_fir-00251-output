

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
CWO2bSovBvQ2ByFi3vbGk64Kz9+OlU+ol4ZycfRhtc5mzW4spj2ZUNH57Z6TD/HWbssYOjRT+UqT
ip6xHZc7sA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
nB5KuhofnITTIpXOtfG8vxQ8BtQATMQkEP+DmIE09Znrcw3yJd8Ym9iSaEwPi49QFbQ4UCNnUF1p
Ci6v7CITkdmn7C29rKsxyl5fQwQ4Yg2Y9J8sH3IMncLyMWd/eC2FXu2c+nIyMZ2PxTUPVrUjVKNp
s7scT7Me3sAj5vk8vEk=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
MNNArzGZfZxohM+fQiY689sNLR2SVnrB6IH+/5sMb7hSfawQFJxphTI8Kro2JGGDqNxumEJLUYrG
7mZGSE03rCaVpdhD6Rm70zB4CVRXmxwbIpEK83cCm08nMbZ8k4fK0avkhJQjAW3CnUztsuq7IA0K
kdwznIXZSyXH6lPiqjIN2Skr4/LMpA0PrKFOFlQVuPkT5ZvNvxenTGhCq9p/EpzKYQA/Q64z1Pcv
8PTscPeWEIpmqBcuycpxO0kwVqiQNRqP/TotOuVFkjYLePFpvLupJo2vDdC4y5SiD3RT9wZvaSz2
Bb8UYdK03OxRsiXtjWytUX0MRrf53QlD+4mRvw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
JO39BJFIHsw8fi/kSg8TBE7CDuzx+VxY3tt2e34SSpwe1+CidGWrS2YpQSFw2o2o0JVA8lhp2pEl
VW+YDwewZ52gevHf/k4qIWqrG228k15Q2kpUAiHbcd1YG0RCacsRIqlWdSiw7wc/2b5Il9la2dZd
yyMNm5GMzs0PBGaInn8=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
DxfcLsCbVgOrlbX9FvTGJxwVAV0OB3tR+6ByNYT/Wivn1M9TCrq2dM/5FWlDqpdxHIYJfhQjjzlJ
F9cbuhfluBOxtIUuGdHg2uX5LqlRjgmnPZ6fbuzAGkBvSUoSqWJpXOKWx36bmV4iGY/0e23H2hgI
ZyfwOhBcKKufNk+Nq7xnSV7GWSBSiZWYhL47CEdCY+E8EYmyeXyXT8RcA9zqsfKsEZqdz1rU0vql
DdxwHxaE1OVS6MuW2h6qgK3l9I9LyDohZgyoP4VpBk/e9sTSLxcSmGiXwe6zlvuSw8MrBIn34Ezs
uAteiO0K8WEa+5P+7J56z0wy1dst9IfRzCpYUA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 45648)
`protect data_block
POH0GBQjipPiqZTDbO2lTFu+dxGh4oQI1FiBNCznkIubPDFn8v2YwwgLFKpN3aMtNbRyXJhmDAN7
fIKMCDI6/irQMGKXmOsQtcv/aNE4mgXJOM5GQQaLN/cfeLF7+6WNEhv9R2a1CYVJ5jfoYz9kit+L
PkQ/2nV9gil5E4yDPoLSmuOqEgWMAIS65p0ytkv22tQSvVGmoZ1ynKK+3mFJOI2nDwUW6EZaWFhL
4joAU3YeEc/JHUAh82/a/kSGjUXMb6e1xyJ03NXT7IUmjHRN4YDxZObDSAMOWXemD4aEKqNjdck6
ujDIWowe2TNjMpooMf5Sfqe3AjSzlsCZKI/6+adg9qKivbRj6EgJjbs5oigS6405+koX+bGyRHNj
ip1QJM2cIGQ9C8MqJdI1HajlzrJxn2Fkhuun3SNsbrNEx3dXOM5W4FtEYwgCsDbE8xXmuA5D6J2t
vh5XOKqK7zIjNatBszTgMpScnie/lj+EqRNGqmgEQqeaszXLT9V1b4LvP+wVAn1HKYYwndl2Puxa
hLsCKX8KyOKfX4xFF6Hf7hUbR9HbbdBtCD9RnRijh4UsIBfdU294NWgHxMONLiVp23QwpEuftbY+
9rTNgQTB139huIktd7B4KHGPQ52ZNzAOJ0WZHEWzkEQ7UkY4J5snoeNX8Ds6+jtNddjUrNbi+fp/
RHEbUSASuMWZfL1NO0Ixf35TB//Ivb6TgVZhh35IfSaTlTEDk27TSicacLbR5450YVsPqEfd4Vun
MAtrR08s+NY2UiFniN4NxtUM92Mbfhygpxqio1+CN9kdOMFVMPsUNXmrVDv2zHWe9oya6yL24bT3
oWRYCoCN4BBU0vVk9L5NFycTk4S8tqrPpPk8gfkCcktL+DAmgRtFOfVQIyNjpB3fwLH73BjRrQ+Z
ZLSagX+QWigR+0bG3wgBgUzlfNt16H01EMtLOTQwIl6NLY+gr6xdoUYNmJbWirANjesRIWjBKGKm
GRtZ3j2pOWEumcFMCoZd4W6k78hmTTAFfbQq2menW0Sn4TyyjfaT/ulfeV6An5K8nJEgOphprPIe
GxiMk8o3YHqGdheel7iLRI8NPHrVOsbIiD820XYuNFejy3VOd0loJRxhnd17PGZNgdFCkuyysVfO
ajXnx0llJvrrBih9wT/GTrSvLgyWjOShUGjsH5mpRmBW7QS4dMf5wYJn3YDWUzgldFlIc/SbQ7Ri
Q/oKNEUJX0TWRwpe1zTidRDRazx6LNn/L+3v70M4Bnzy8E1O/+rotXAgMCXwjVjaFGzSnnetWVox
OxDzpDK94nxHniWt09iK8CzOdQBhCNEOei8c1vg7+VDNGMrrJn9nNUJajAqDJ9Fq7UxOaoRNyfe4
vafJfT+mugH/AUsVON6Uex4Jsf2D4LZ7EpaVW4M83bilS/49t5iV68wAxvB/5tY3wybUwxGYgHVX
JXCRp0Uwx9mEkGUtfagKUUgse3mTJjrjxt00llDzgaW3s6Jp1EDArJrfcc6li2d6Vszfc6mPOEyt
NyfbaTkxYtaIi3rOlgWcsBvvFbErL5YSt9zuI09a1mc/k811ENMXUAl5aJJA6GiaBh16qOl2F3mT
U/aFI/9/rMMgxdzol9fmBmsruksXmQK22yso0SON5OBDlDj4N6kM8f+Mx6RB4bg89ldgV7r3JNxz
9SWyFWIOp0w8c5/8a5qEUeKyboJ8jX3aqwguIMrKv43kXBm2Pb8L9+pOX/XOENRFjeu/Tmr+gxB2
HiMTIXLUZnhyxvOd4Mz10WED08+TCXO7K3HCkpz3mBbkm46KheKOeFlMYDzVoAXC2JtxRkKKefRt
ij7Mb8HWZBAuXNkZV5gwcbEa1LVM7qJEvejNV1C+CRbY1aquh2vnfMNjY2/e2TDdMXOr2j2MCvzJ
akgvD/JZDEksH29CGq+94MCjgQSlhIY7PM0vVhx14YdrNokE7IPPzUWzi5V0lNmmRhMK1kfdU9IF
6GZoSeND2NOuA2aAmLGNMFHTqBB1oTo/xCdBEz46LmX/AfpvPUx69M7lVvTzAJMDJxIJKmmXu5EB
ye4V7UHmtC188T6gsG8Rl8LQJd/q/f9Q7O/QOy4G6JqGJhj/dcyKBpC58ZmO8ouKCB2pe9v74aqQ
uYTN6eoUXEFa2L+zGSsFztHyEiPKuvP5LgIg8E0W38o6Kx0efVHXmxnlSEh81PNxaraBbDbYC0AK
Qo1yflfhpSyrP2YodHu6II6Eh0NQxdH2OiDI2Tz1jDvoGxOUVgW8kbkObmroyHTR4sDQqwWuJ9jM
DjekNIVUoUW+Tmffi3bZuMSn0VY+UNnZS+nrkFnJT1fBCk19lGVScUA2k6kADxm/myFqMaYTR13Z
sTCXpL515m6odHmX5hJzmNuIjYCHVDpjQXDawQ6j/k+7x7zruKqE+RfYXSGJi6/twqPztK72FYmU
L2SYkvNy5MhqPCLRwLmKtNW07Mc8sWvC72ZbnKkVAgXPD4DQbXqTmRgNyEN77D0OonaDgQyc7nWf
aJgkzuZbiLorj+GAna4u93e63YYWNgaF0zuUbW+cm0M6CRSyZv/lGoQ+TTvH4qXYYlVnQ1USdboK
qC5FktZ+GgqLOBxebeycYVxjVKAXQLXtJ0O+YHcIFXGQFzmdlQPAqBzn1yRi2GKHVHxfTzZsb65Z
O00/CX6+MY77dw6wkxy2W4oPh8KBhJ21kjSkfMsd2GdNAtm3kNhxkzH9imNYF3mOz1MfjF14e00s
Vr0e3K5mdEaBjIo/ePIhWITxEH56+JI4FfMCfnMVA/m2Wkx3OJmUPMtk7tV6lxmhtM6F5iEWPQFn
8gN7sRX2NoWQYE9jYtAhNJOjsxcPhVbQp/8NmlgKt4RBwQxADP9sqdTXQlu9CMUfkH4OgmOQff3E
CMpte6klTBqioCpXcC3MNJedibJtoJIfd4k85Msb17rLkCZb9nlz5Wfg75z7BJhMnnlr5XxIMMlm
u415gHJfcmaW5kplfIwG4tLH53tg3K3ddaJiDcJRqyHXqx2NQFboaLA7tgib79pHy67/FXiNdhH7
jAil+2QkuKo+vLCfboPOXNxB2PkK5vd8lzwO3nUWnk7rrfgPpRNLwEjQRXikDD8zwiruzkC9ryCf
9ClD1DNsBtPyEk3i6jAnHkDUmDkA2j7MfGpZfGtLNykBZ8ZX6Ye0vFWX5JQs2cy8Ujpohq67EG/v
++Om8qTK3qQhaWw8zrm5jc4hbKAwBgJ3OIZpKeHbcAHeRfxbPyjSAfs5htQzHOjwuzVrhq6untf/
2brI/H3cZY5v+3NCwmW7aMD3QFPpyDkX5D4TkKDt3wpPovUhzI5z+pKZPadbOKLzOYiFpHFl9JJk
ORW+BeTI2IxOUVcY3Sr7VbdCpLDeC20M4nr3J+3mnS9VJgIWsdyco1mq22stGfQSKKIDlLgf0cqt
hx4rqqSGKSKgDMDmjei3Q8Po8BRp+UAaZJWipFVPAWJUabG5353fRmRy6WyT/0vtfGwUr7+nHWaB
oxVoDbTiEf3X6EcU5Qk9Y+T9kKtlKzAgnBC8i8LELkaz/Mi31ZgK3ZCWU5MBnsZhF5vBLYJvwVIq
EWfcKzvSvrLxetEmWoAjMyx2dBrfx/fikyVf3DOgt19nvmOslJ4B8vO/4N61flZSQOAgC6polsJQ
duQCIccM8Hm1t8QdaUa4Co34YLL6gOSqkgf0mYTSAzZKsBwhiOIGcNS7rGADGUd6XIDdJ51FUAUO
+TIaugKwb63zgF8oKXIIJuXAV/SGmZ8zlTSntcXdGhcOn1s7ggYfziLwGyYtGFMxfvRtzpDf9tgk
UGN2Ty6kv7OVQL6YRmhN1eNwpW5f191dvM+8UzVuR31vBZNYrYO++EH5HYLHy3qLir27IoKXN6Cq
6Rx4XzUZo4BKDdZUw2axlCqE1HouYfAJJfHuS8AHonFT7PeS2TLiFBL/8sD/Pdxjj7tLdbwInVcW
KHCub5xUEVlSePuUKXI8R63ManB2mzKKFJ3yxboLkvDtv0+zjOMrgjWhcOLssChr0eUGu+1F/8fn
x5ZIQognakenumrP8s6+D/SD5eg7Z462fLUzCeZ1cIvEB9Xb/lswx4rlC0H0lC4sf+64MOZyv92R
lqTJM1dM3M1VUqqBOcQTFIBwH1lUiqdl8ELRroj4tn6xbRUIsjBGxzf/yKYw9JMoa2sucr33TxKQ
gg0JhZMPL+uwswUwsfMGDJOFxNL6YJl0ySph3qY+nCMpfnMJ7YmhDdeK5gTkUD8NgS33nNq5Ulks
Km8S+gBCJ+hsHD/jGwimz6EkCCDOdBoBrogdH28o7VY26Gcp/vAI26wYqhTQnK3SxF4uX4pDX+8G
K5bs8FKs+H8vCwukJi1vD06odoSMEAOgACo8DuVXGaigZu0Xwrwr5xC/Q6exMPtJW/3hnrYhjo84
s+eBZX1defbFuD+XrhrbAhO8TX1UyUD4faE6M5c7EGEuWcsKDi20lzKLJwxcEycl2E+oqb/CEylN
phmLujxcjnoO/mSyYKgodtCHXvPa/5zwgZJCrmOK3n8NH+FgbKM2qd9NFZwvpS8MAnofJCt2AWkO
yRvHf/ABFr9qb4NjH2YzpAZsCTrx4LDEMZqC6+Xc/v1AYoewQ4e0jcz1IHVY9VuNCG9D7B2V2veH
lhBLxDTDuAqeE3W1ttR/ikGBUmn1GP8cFE4olUxdhwIVHdCdPMsBEOdcQSAbqzNEQ5/RwIP+b20I
oZ/mdkcJC4QXcwX9o5izbzE2xstaNNsyp/i76AGKVY74f3DHmTVtdrye5Txg0Pb7+Zd9X4ICEXrw
NxzuNBYt+439JEkKvP3CyjD21P41GR8lKyimeVyoF0L2OL3Ttv3K7TOc6TOuHQrvGxqvHx3JbLB6
4d2cy7/EaYhRbUBf2/uk+GxFneRJ0YiEMhW9MHvvbOORpRS9p0hFcuQazrf0WwARL3YTEOqBMDMl
1MQR5+3QYCFFMz/lD4WHhMEMVG70GexQwxuK+BN7mQXujZth7Daz+8UXJGLjIfcp2c7XzR3XpaPf
LNxhuY8ASqMXXtdDdlA27I+6sjcFJOXJxAN3/tomEjL7jHUCWPMsuvQ1n6Ij4uIw64O2Ijd47LTS
FAnOAq7YbO/wn6hVcy6Hn3+FTYGlZ6ZK45xw73tVwzptRGyl6R+W0v5IvB/oJ5WfDIuzQ2wIa2Ar
dq2z23nXIKeQ/iNDEU7SjzDq2OVMiQ1p+M7MY7yWN96xGJR2ekVA2SiPm/CihzF3BnMT9tpI8xAT
Rb4uv7Kw1pwtefNHskNtZnyacnQprWSrj162AE53MuZ2fAfSXkvkzR0NlU1LvlrbnYV+Ka5B9nqN
gijtaHku57Nv90cOmJ+u9dHB1cdz78wHBGWgXf7cgDddJJHG1odvdfdz92kuo+qESYLNWWQJCZud
l2ah2W/MfnnSK50Yo6WHy9fuzkkRxyH2G1BbGbpRzTrugLddzI3SfGtqF6TOokT7FuR5uUb0Txvf
oeUzsQQb6AIKGNGTNOcil5o0zvr4cP4gGycj0wVm3otzSztTMumE+lCYuCV4E3OrZadDXkS1idkg
VK4Ks0SxaJc+hCgqStztV8I5O3zC4FNZXlXlu9Nc3ztcEun/KFjSLpknXwEg1pzC8VsLAinNIhZC
siM1KpsLyFjunR09eHu8C+sECmc1/2fy1jIar9B+JKJMH7RsrTtYezbHbBswG6Dya7g58YR2CX8v
aBZT3AoTaDulNlKawxsekM937fXa9/bEgL2JdG6v98QJ+KB+hMZeCDmMosxyyTEVvbtDyGn7Jtyj
v4QGe4USBtSv7sZRltfx0sw20ufRTzTO3Ek8prHzBMqBnnlu6DVtqg9EPto3MpVcwvJNgpzPlfQ4
BmYrdA9KC3kXI3H5dT4E3BWRH10HG/ugD8KRnAS15+nhJi6ehe8s+U4VmZSfXLH9nOzmC1Ecjman
1C8NZbOQkXK6eWSodKYifbPHF5sl/aeyJ17IUMWyf4kxh2cq3csZeOS7x0QlwZlM7Ak9zjSZBi5b
QHgsH+9uN7puI2RQpeI+Ha5yEKRnxmW2OTurGqQOuUU3tF4JmQ2nntP3oUoXDDmEZqa+xuvri6We
wI4EsqaQHaDSzT+IVgnOHFVCDWRPCxldiv2ZiaeIjU03m+ci2lyhuOsZO0PSS/Bau+9mWTqVFQ2R
OANdXxyWI7tnD2m6laSqagwMdp48YaE3Pkmwseri/UiN+dprc8ziTqvxAsu9SJvuVVB6iKoLgrdm
6NQJWBD9reNyXBfraxN9qcEd43o4PbUHJ/cvjcelkIt73mCNc+/jfFrvMHoMqijz3nZg+PzXJlN2
caNwgdbb3nAkz4J+6Cfso3V+z39j3wtwkaOH+SyfroSNHPpAzxNtUvlYipgpaktDGhDieqFSWwKm
cbzBr+qMr3jPjDse3lZm8wzz1tlgiaSkr9Og1I1qkFyEK3DFfFKCIIRBru7D5xJzRZL1gPrfHNnf
/zPgCPi8F716wUsaNTs+HnAmRlB8rw1m41e0vS3c+prxuHs4YlmDIa2aYf+iUTzn9ZScLjuD2Nsr
KkFF+VJDTQxlF1WV6qWEqvw6mafe8ZafpUrmQqmqaibD/AWOAA2ji/mcyOCt+YUy6URJ+vP7nrXe
yZ2drRgPHpAHB/n8KaMC4KD/6XotoVpGa80jkm1SpYr3PNKMeMetX12ujha/Fz/zV15+YTY6+z72
WF2J4cpaM5E2LymS9mF2BUirbn4LRIybIhdKrAhBNUVSRyQ6R4t4lgLCppNS6+Eo4MBXAIr6R/ph
fC1z3SAceR3sJgrug5Iwa0JQPDeZTEFIfjePBIKxIkPkxQ03iVgKKPniC9Tb+QT1amd2I9dlTNGH
gF/2e6aVBselh5Gjq0CoAKjZbYHw8UIp5gUCGzUNvvpPbN5aQLKlHb3YRfqvpcx9OzfjDtFdmflf
Lkq8LFfcfTgF7sUE0pwpLtBeMNaup5qv4dfSZ7vj8Jg8jo2QdmPj5mS9IlJAOXYd6kPkdQ2iE9Li
ibtleJcX/1ab74oa8o4X+Z2DBwB7VMgym6/xY3ckhZ9q9Ekx6aOSGphEpxU/TrrhlvS/yrwoqkIA
fHHCoMocsXJUSk0fTxhIWY92x+B1VCySnHj1GafSRI7OrIxly3bPuI6Da3HJc6boWNOBLl0XV6+R
9NRVQNKaydQQdcyjW9pmxTRN6+svqx4izSUkWtRcdX+5QMQtsD5uJC+aiaRHa5kyWFY89StL52Sr
W99tp+mOZ7yVXIl1HAujQvqtI12vrdcqzfe98DsqW5Bdv6arXihnpRAT9SkpPxGA1gAo4wQ76ZLR
QKxVBFqDfBFbSpQxZRlSS/0ADEKku44otH+Xzd9dyTzj4ANSaXIIRiaCv4L/JC8wtLwxj76WSUsK
15xJYWxq49p9l76vNSGWZlkaYZgQQQAxLz5DGC9SElfe5AboFLLV5gPOIAHIyPw0hPCClGxY7yJg
rNSJJYRYPi51Tp3jC0TDwxZrmi/LI2bTCMqTeHdgO7o0N95YKl0rdvUM+lMgrUBSa2Nd2JENyARU
lhggNkF3pNyPHV+hPabOa5o6i5wyZ8wFh9IRhiHzjZ4+AJUwhhIhy2CYpYdEn1Vn7aT+m4NiTQwb
DLbj/O2dsIn41N89EHxR4Sj+hj7k4ar4xFFSOUSA852O0lq3IhhgfJE5LFbCnB4aKeCAtjcdm1W+
VEPb5S36dOtfGL9e6+yxd/oUXG4U0QFRtB5euXEI3MPrFw/70isRygJRdQMJGmYfBHqG1udONJ8C
vpD0o5bhJU/0gW8KhAJiXufxl4E8dv1wK6kXI2rCjxGe/+pBiaojDZaUq7hv9ljLMzDOlpFy3FbZ
1IZBiVX2mvM3VCXH2R9G8mHhbEAwYUH6XQ+5yhIbVep77XdviU1eudVFGxefvo+gQkNhJ70MGsYu
5r5TTE3KMwGiMgufPOVfwBjWSQmv+JZPfujxzuAygNIlhDHiPryRqH3AMFhhm7LL00abPKsIInTe
vOu9F2yEXjSFymPafLepWZBHrlBxjIzs+XyTIABuUP8gIlLpaG6oVLo8wLBfudQtrW4dFfR6hAyz
8tPzee/tIQULX8CrhvSgYBVvaSbu+Cb6Hw974Qmoly5dZmKTtwwhptZiY1f2OjqrHD2rhlMCjhDt
FzjtU0qWY8+M3GnKeR0m1qJAfyN5B6XyL4Win5+jXo+7REGQAaCmC0BAs98WHvCvWPOug9gSxkFg
1BDhapy5bUXrjHb1ihlDaDK9vqd/E0xMMz5/jhoUkHlMRvI1k9qCI9nnQ8C+fm9ud5Eko3I5So1P
COT3OAjbzPJGM0P+pk4vdGV2eRmopzZjMrCs0g/vKrHyFIUsFIUAqXrbVZRj5i47XJUny/HmgQpK
OShEfnQvVtza/nf4AgQSek+LL4/ItEV0uMMWsPKdw8EhKcfm8zoDnfYDZG2mDvERPAJWSytfhKVo
dRmzVJXuSaQNXO1EAQ8l4H3DhKriZEXCv+Mndkvw02vua1UPEv634nCTYpfygLMGnd/eMOUg+78U
nFJSk9Ggd8oCjGNtIV98uh8sEDvdKnIF93XmZ+kLa529kqJ/1Nr7KqdoVFEXHNF6RXx4uZIlNEPF
hf0AiHDjdVZ8pYM9ZrcuzYV/0HFaTvn/WrNjQqatnyjb3wUa+iW/rNoTwkF2UzfjMtrI6B14/eAS
3tJV3eMQcCKTQ9ddDvgELXiEzjyR0RGCd9BqQvT9A0Shb5FlGNMmtuvuePAguXVgV6Ufps53AbJ4
5/0FIkzgRJvabjvRyLpomsLJXJFuxXum8X29xTgxK9MpKIPOjbTqvoY9ovtHqrCY8vbqMk8LSDdn
+Ts6KlsLDwPHUhQVDS3fr6RtEQNnYBmPJ8zpgQqdW2p5lsfUgh+r0hpyyxO2Xd44hfFjfGfoMScW
uNcMIZWKekqaJZhv/Ghg7/om1d9bfdgrnalrA15skNWnFebUMqXAQyTsKR2nLdpIXeM8x3H3VD2s
8DWB07fOiH+h7SAO1KyiN5KFm3JOoUYUVwg3+OW7aycvs5gyV6+xZvBRMmHirjLmHVcTksVNofek
aysAVilFfn3claXdfYZG1e2g+yPCjwGcRROChc6BWB+BKEOE6f4+xNsZnCtp278QSgYsPs4XRtD3
5pKOyRd7uJwEEeSM7knvXmJpzZIuyJhgQGGx8xHBXcFeudL0lvWu33pvc56zKKx4as+RJGWRW9Rh
vGs8xXq32hoUNFVk7/yv+OBLGQol4U58uKFqdELl2ewHVsabhENLdmMFNw1ONilfpEmEMoJqAz+y
/85MHfua3QcFL21zzXt+L45utvoLnU4wgUwIash22dK1GhhxC+YAzQEytksCZPFu1OHVeXRCfdSo
oaReBNtFPBjXo5IKKHi5rvpjQjIVf5J8v2Y+B1TyrtIn1yi9uye+pSfcrH84gwPm78IOcGruYfQZ
UeEy0WUuoBAbRLqD204gS9rZn5dUclIKo7JHDYOXOo8EaXIj0kbnr0Jmr529iQI7OQiGFv2iTNkV
H6mEG9ydOgnCHK8N/Q/b4zmooYqKi7j0hz6JHGpa9QIpV6uKEVsJxGFBcedy2MQRXhYfl1H7/rUm
huKWgwR0Wn/HP7xlM1OK0cUdOIuKb5dEM6mU6btQbYVmv/I8RO2zsxZVy99Pv3V6nCUN5+fEw7gH
4xZgPxviuRL4i+1f33YacJbz5bOc80Bdfjlo1hdMkZfUnTHNkY3OZlmgPQNunX32k2gTlx7SbGDR
NDLTWqquJiS7lYWL1Uw2dyRLv3Y4y7emYux3AlCKeRVx86YQJWkyHZOQTzYoLOPaoqmATPv7YSOf
/mKlWa1yOaZ58Kt9zao8ejfPaVY/UteYBIhr/nsJGbln9kWn3WKYMh71DmobS1qxy6N/Kykf/Mi4
qZoH/NKm0q0Mbf2/MI7u2wUZnBoKHbVatUXHzcmuJN3h50Szq+B0rqYprrWEFOYr+sb5gTPcB5RL
N9E8IicFe8rI9F+PaEpr70ZszOcaDk38ws9sDj9vhYfzMXdzeBsANzfniQsm7ZeJZuG6WJWbaboN
5XyXxXb/nLVWOp3PvDt6YaWVKCz7M24NaU62qTjBO9+GLNzIdltkvjPqzLGXi+fF1ByxuaIt3yJt
NOm7YrkOdDKbZ4wgcBDkC6b27Fr0w1CSokFsYoRBBkQlhgXWkQ5V4T3+56d5RMqwdJwRVWHTkEyR
wRaYRrmx0N8NsFZEDzJnn25n1VnPDuCp0hpwd5YXSe4C5ZnQ1XO9U+m1+byYzOXp0ATRn3tIdpzy
3NiDDpY/vFUdJ6Ja5j539FM5exbL5rkIBCVuX8ZMViEcfWJOc12+C9LsGmh7iorio3QuaiXZ/gUM
J5U83VNxJKVBAA69sdwGuxK9ZUi7RIjvExDjseWjCfC4Mxdw6Fg/jbuaii7ZK+QufUaxIOLRTES2
pWB7S4a5SIfkAnywa5+ATRBW+AIi15BZaKFa7Ab7KFeEIlt3Y6XowSG5frgkrhMDTAxhts0G2rwy
AONs93PxmNZnnSSDnbjRXeQrcdnYBcY3OnxmnueyKBbbXK5K+Fc2CnsOaSnSWXLJX1cVWZRi+DOz
ekwUt/jipxS98DS/JXOvvOo2+JYE85YDCLUyErckTU1DUXlPDMXkpkQbrBvNRRY8lM0cZbbBp+ob
hJRoV95sOAfKUFH0m6/x8VrNZV0GnNtGEqTauRqX8lT8UiHwFh8TOb3EX4JBvo8T2WxMQjjSEPts
1g53RmOWrSgNvBSd71N941SLzlQl3kERUipUchYvwriraRugFuQTNviV/MoFPPbm0DO3G7SD+4Ei
DactjwFfbFO/28ApKl6iCIekE2TMFClSVbQyMewqxXVFpV9vx4OW5bcpxc1vX/ZvUQ0vOHuzT+Go
V76p6/4lUzD9XYtkD6LZpfwXeJ5KmeI98bsP37PLdD4HVPiLkihUeAye9buZ52OUPrGKfhUTnCRR
oY7vJ+8ojCoIHVxgXCwhhUyeJgQ6OE1kPfSsUQPY0vD9C3MTqxzPO/Mu5qatSSElwf7hQIhIDS/1
a1wXQVFdzfOswMw3CRRRk+x86NKtAgeyP1OC/JQi2BYTI4zptK4Z86vWqkuZNCY0wvNx/Z/FLuAC
SMtoBzB/tYQg0XN70DBXi6rA/Tq1312runNf4M2RHygg6vYePw6LgMpn8iTTQDZzaSS3Nr2Bxlg2
LBTlt5YLJ39ID7pgUp2kKFYP4JODOwyxl2uvM8ZchtYdvSpxSGY1yEytfA0EuPoomlCoDJv1+zI2
ptHrldptA+I16XscBjfb+1OVDSO1FRvrPfN1Iy8zFK7C876cRsq84qqs1JMSqNtp9flUsMn4+Xsg
NOXsGFEXQPbcQT2Pre0WAnlYRGMDDaENifc3d9WtK29I2ECtARuTWyk4iYSYsHsvC4A7p74bgd8Q
6q82WH5101ZFfNjpMoJNby+xqO2SVYKM/Fb0iS2mw7AuFJUSbayH9JmZGGqr8Lf/IedzxHxGt8k/
B2h3w66Po9ztWEUN+dLufFdUX0LhYHWJFdAgR4E7oSF+mU1eP6zW+I/d7+SAH2tnGaD6xTU6s+VB
JvavM7u4dfYBGbRw1hYn4gOtQtp/arIpRt4gL3w8cwXCfFYwDpQjTF4D6dzfC/hqhlCcL57leoMy
+gs11dudx/s66Sxxzj/j7UAhTQtUtxJXTEToMlZd6HUXYmiAPTs7WjO9LlZfsTG/ox1oUEdOGow5
YK4ScKKaPtlpJFUe1KT9W5q9KGyyT4kJtdUxim98Abd1DcxS1I5IUGNedgIXZmpOe1qFOINfBM9r
Gpr4qQEhgU+3XrH3TB2qFpfbPjznDlyJpvilGr9yMxwH0gC9lCI9A1kdf/H7NtQ4Gmy2i12ZQ346
rShiHa4/jnUBXuLBwllP7L0qGLsJAxGhC6DzCM6vu6l2qRNy4k5C5pYlRKnbSNHIBDxn9oMJq2xI
xEAIVJ8mYUNSygBE55IIiqaudRmt/w13/oayl50mfOQJLTijeyCHyNMU0RsUU/OuLE3n1kEbzZpQ
R3pDN4ryaypi7QjeBU1j/zAkcX9Bq9Z8OV6EYZQLTlThqpa1jXo42tpD8vjrJ2Us+OeTIR6CjSI2
oXH198d+FV6CTyVqMoulOXHcTXuKuRpV0A0JEiqgTr92jszhC89JvgGwmqgPO09LfXVB62TKXAbn
UOzNcUynwB5x7D/cDf20ir/6DubHhDYwfG+J/LmEpJJsWOA7OwEf47GzK/4ISfdcm0oaLJrgA83m
Y/Oq90hffUIv67M38ULGWw748fXhMD1jY1EtBE9Hg3OabmX+7ZWZXiltP3W/oALHe6V9iXHP1ZPs
I7mPycuw6BzBlpzbecTuiPwTGFGyYFm3CVwy1UPZF+tuSkg6XuvXzhsBmmBsCiCeYNx3FQ/YvUzM
wod2SWfaj/r5MVK4jBd/6JEDR40PBTE7oBePmaoX/NN4H5HXQmJJb1PLTWQ/hheDdrKBUpgDhNRv
lL/TZQibAfz6WwqDSkjOFWx0WSyhaqwAS890zqbM+9crm0H6dGvQCP76mtecYlrLtfdNZy9Fd2pT
n0bk/32jjhqIQEcZbbha2w/MHFMMLlWvQcUSn/cxblWcsJTVo0+UQEaJ582qpLBhzp8MoGwS2Qe6
TpE/lwTFG6dDwHtwVFk+1AksRQfTR5Qx0ONkHoc6ExrIQaYJt2RIGjBDvCdIbMGPxB5WTg9HMZbH
c+2hAO4EV+45ndUeYI9fzSk+ig/WbEW0d+6PsQgqLj/T5zu24uD0t1S3nfXABOEcD4sd3svaqQF6
oTOEWztzLBiN1l6o72G4Xr6w/ZNmzMhkaYZYrv0+BIFGpZpXBY1MKtvzMxJnpadK1S+GNeDqW0E/
PrhuFb8gFFt75JLY7sJ4RW1hvsyNi+SPWs2B4vnGe3Ol6bYglXZPEZg8uBMQUC3wa0T5fecrd66T
QfUmhuV3wHMoTfbGINouQp1DNtcjAOtsLoV+sisGfnBkcs7oBY5EfIVOpF0f1HFSAyfy5WW+3pEj
YVE8dYzFza8YyQepdP/fqvZVSfFr3XQPVnmnnysqxLVPMOqSs1jSZ8i27ySfgQSRRVyeW6juhW56
tpUkRZXs69Ob/c8+8/BZl7aCjGajcYkCrVPmOYiQvx/tgN1cDCFlxopX1ACwnLrTBLkZBSUfnCPm
zYvkEiNSMDW7h8KIyUVhMsT00Yocden7E143Q0YWeWZQwqia/qOlFSdTvC2SJvQQM6qCmxBFcZ1U
j8W5TWXn03veKdtIeU3F9pWpgOo3SutEgjVzBtxhRXA/aFxEqPvdcZVqb5Oz7zSTKMTsgVv8/ysX
o2pw0ILyAVdDzB3S16gmlGqaqe61SMCMxGvicBQTvGXPt39/jBEgkcYAc2acUcq4n9RIqOgV/E+r
0us8J+r0iiz/udzczD86iBfjaHAKIwwmC41CniTzKdZGbycVGyhZyxXIwLctOy+aIaq67bufWQdC
mvwGpvJVm9DmO4cw29t0+empmXqfgiJZvfFBHdbFYbEU/O1azBsnHX+G4dB+7/QzpRHu6G6+xiTI
AZEJgYg3Y5eAJbHTYOws44HAN/cm4nm0TMjvJ4AnS2PjNAEldHvPZjMI+kUABEf1x8Cs6yahpS7W
Xo2eRI2+2Z9up9imqBubYuenz7Da4HzLT59yRd8ECZjjq8L137MnPh/nkBRgwf8T+P6/VLuhi5TV
lDUElWFhGUoW6YXI749dTzzl9Xsrl3Xl76emA7whKe6zVO9twXLaTAqN2uzvJTHsdmCtSo1Cv2ze
pfbI4hM4XrlHXUElrFD/qBnulTitMe24kr4iy9LC+rkHCjC91Ao3aiK5pTnpvw08oSQJugzZqvTd
hrkpYhzrpzFmtilbEvLYUiEwPfN5WHMEdr5qyn0KAAdE3p3JILK5gxgSLbiKJuctLXPtc11v8HNR
2h52c/Zwp/zyzaSDf4TmMKNwtR5JXbZY6Fa9MFOvYXL0xlP+6xWw4Z19YN0WitHsfW3rPTbAepco
y5Q/d0/rVD2o7GsapVatsRCSNqE0+KKOr85odK7Uv4b/cRJKSlfrQmnlhXx7J/UfwKf38fVC44rF
hgk2aP2n91dhloEU4hgZ8yQMrhmRawIE/pskevg2zpgKZMPbjsBPAiXdNQnmp+8Qeu9dzgnhLYpP
ufDTf9fMjlDOtrQt/1Xe8tpS4VBMvdV9FEr810wwaaMZjo0sxbttTiOkjIxhlfHM1HE6LPIdGHEF
ONA0hWnj58y+NoFTvWf/TE8gn6KhOqHHme/3Ntb4C34WUL2qKpaKFeJ4qIlyGiqRQfri0zhH8PVa
IjbCbTMTyX725USutnyOV5kczgLI0Is1fEC+NGj9pa5Qvuu1cf3sZWtIesKZHJt5opn9Uj0ZRpga
vT1yG470UlXlgA4XVWEQRNnAih1Zfz3Td9i0U6giw73BBTlqhYD1Vq+JfkhCeA5ttrWy9YCK6usn
FqdaJxO/U2ltJM2NytdDbFHKr0uufywUl2RC9yl+9gXWQ59BDAJxGlbZ8hVKZeQzm9kX1qT8qr6G
pYh5s7VD/CFKJED2cdShAX56npuPh/pFlwJEs7kvl3QKtp+Qe8A2HKvK7gRTiGU86VlMsLZX79+3
OZJSpBnKeehlAk9jGOaROmVL7c0+LL8q1b7/HGGaXTO8hU7uAgIspGYj46n9Zcu8HmJ+KCWybBZr
RH/dgfbJBHwSMMe7iA+WsdaWljtAVGXuGlvL++pgwr+5Ku07qgNkyqgD5RePeN4AT6yUw82MqUzJ
coNIzhsUZi3crhVbQdOiNR76ZREWWiAOWAPsOKbVQjG0tHToWpe0fxIJyBp33tOuO0UNHtikis3F
93AdEGPY4VL17KPYFpVp5OvNqxjEjdZvYEQGIvp4qyQdrICt+ToqYB9o3/M3vPFve4+nmdRn6KsC
ySGfyzkrufd3jn975WUBBK1SrPf8QNjt903L1jszuhVVbUTilkzL90KAHSs8yvRaEbQ2iuGzN6AO
o0KlecGAPNPrfhddsGWSU6QRUEYO0SoyhemafrB3IAU4IfkBIVaqwpJQsIPkqWc+GayBeQM9EOpI
+CYtyZeplAnZ3taiu9ZJGwvEfK906uW8xIgbNWqo0PFsf6KiRg4Pn4zLjJnMmcRaAkF2NSWB3cCP
8o1Gw9kRIkwJrnARL9F18LJhCHF0VdJSCX7g7zWP9sB555SHlLCGizAs5rtyS25JEDO+6Ng725fJ
5djOz1RLxVeY9rdY71A3fy9elkwJRxmD4U0Lm+zvLmzpYQtuQmKLcAqU09yCcZsn1TzhYwl96F8y
9cRndcanOrOIF9KF3zgQDhC4QzkWDX7o1WU1V8R/6HPWwr/zQVQUfTKFXI4WFC+3ZLSDV/v++QX1
DoYC9wV152N6AhSs0FAxGAePMByQFySXUeijV8DxLC370fMpaqqlQ5IfU1IKik9OvTLU45hPB9Rz
0TPwhQdceG99zH2vw7Opiu8YoxqBQdO6N75e7pwuBFs+ZVqryudD6m/8tds4meANIM3MigJz9Bc5
oFITChwcOOlGZ8/+dtttejbSMKUwvLGSC7xhQahGglnWbk8Mo2oaDGYk2C+JNCVvg8jgbPj8ZSs0
n+jYeT48HrZ7soxhTQvBMKus6ehea5AGN064FYTsgxAOrFWOiV513ynU0Ly/rt5b+92HjyYyUWa0
RI3yDAJaYidLsTZUHyVUAZ710ssEMEwtYDEyBAMKVmpHhuH4FJQZaMyolYr2qUt09Bv8U3MRrNDF
r3ivvGLTQUFos5rl6U5tIuTLKTBWSHHKnBVOLIrZZDa/kCkLNKdTO0p4pQUj0Q+MoJA8RWqQDFfK
vvrCdSHeG1//g9EGWF5s1wQArCkw3DXqasLFoW9uL0eEPSvoJt36v5j4b2JiXIIlZxAdvCInG/fp
IRdbg/SDs3T7QJZOSRBv5SPzynoxKf7zilMdwVsQaXyyDoUDOVMflhS4yuJDM9O2Q4C5YNNID+UL
dSq5qn/6zrXQ9HvDRCMBBF26AddQTyEidyT6rRBGdvBCgIOHtKMks0h88NYT0ZJJv16+/PBgF5EA
TFJ70dq9Kx3NFDtOpr5m5d26sWFqUqQnO4EBCqXcQIHp163abPaat+oCtdv+/ZWzQfDJaz7VjBl/
UW1V9QFt+1KproN/xrU3ihhtcW6gAqnlwS8EHNFBJBrI5tekkHqr8Ktkos2Icf7VpIw8LAFNEDug
B90eRMvMAajIhj4MhdKQ41x/wJ+EMDvKzTTQGBagITFEqluivD4lhiXoCFNlsaHQdrEk+CDvEim2
dkB59sXQfhhanownWpLQXTmXyOqlMlsJD+yYncuIUGuBWFCV2NMrKY1PZ55p6LMlhgH0JhOEpadB
CXNlibJGbUDL7BGQW25cFavjUHNBjxcn+e/wcin4nGskevcB+nNt+LuK7vYlJuHbtbDUGUY2Mpan
FahGX8Jq9rVV1eLaRFuS07m98MSy/+e4npNr3QwVna0WquLJ5BIfbR3FxMI2FnxJJ2OdlBpHdxSU
Y5MO8moXC0eJ9cAohfuZ+pPElMmEc0marBAprAxonRyTZq3UYR3pOFiAbdEwUMLM4og/Tlwup+qR
ze79h3nkjDOl+fyXfkfhKN+ZCfyfV6dZvfC5YFFD6dBWp6WeCQ+c9K8MARJkblscjUpwtymeJKn5
67pX1w2j5Yp3e3iw/8cHnmkvqEM0C5ZfTAI2VNyGXW9HlXjZ6GzYUCr+ZUfH/CfSFjeVhNGn7VGT
DQ89oP2av29RxCANjsAGwPEBKvcC3QkwRUo9yeDGbRsxmT/O4g/npN2KFVNh94ntjm11ohNHQuNa
NIhmlnrev8wLO0yUpmTiDum1OAdxcxyy8tEXH4U8pUwmcqAj3kGbpuXQXRG0hyu13bgAzp0QQAd6
wjnfuSM74WLH/dy7NP2rJhMiulYr498Iip46zHkCWf1SHMr2y3REatudA6TWBNg4ip5Q+93hBaXk
lYaQ0wLWPmAmuCoqzW0pBDsqYOK8T/i/qFN3Gtb1edz/XKlTtwpH8D2upqJyAkzjrXjwm7ekpyGb
iSzwGmINM6h8bFX7pVojXT11xE1aUV/6wGJWiyT+kXJS4zJ7w6bMYdgSXe62y677/ZmWqLWDmHpI
pFK0FyGF1dH2LFp4in2wG9gVoe/NFBnbpukcusdRqGqRj/CIy40HclrVgAX96CxVfxDLAYZOrQah
TB6sJCujwT3+aXMEv2adlqP99vETiUd+d2rkTQ/2sDjnvaA9dUKt39didwBx8pMtoBKdF+6wGWlW
pfEI3MS/QQzhw2C3xMbeXFVKqViYTP5/gOuRIUKvIusdyVjhh8lxvr0oaZ9yMTqbMDNSIZlt2Ww0
gcBGWC0db60DWVp0u8qVerwUwMTCvDfBy8rrGx0Dw/MU8H4IQcG/scLuCS2maDMlmy3uBFwEg2uL
YhHL2PDXYbSKrKPirZ3v9BABHVsnyMH8iPHeJjlq4Fx6MxGcpE9GfDUsweUd6jwPqU2AJvJziX7b
jqKMRlSHuqDLqms/YDZlQlP4ftVNFOetHDwlikAMLCKY22/cyo3z+lzvMNxApazXsw//oMv5RhVl
igJ9d+NQaSr5Q/eBPg+4HPltiYVwxYXGTEN6kQrZn/+uBngLkRp0N5WlDfeVw9SSXcu4jfx6cfBr
KWa1FRjkUp946OC0FRwxtuEAY37v7nhxMjEt+aidSTapMcgwfd2W6w9c6ETiIOHtJy1sBCBFSKvV
i4MASf2aFuDJLy542MPQVWbLjr1am9zIGcKqrM8wJgtl+Yoa5X3EHPkguSF1JeVflvLRGy6iuPXB
hO9jSubRejAukrTZ9GiaQ5AxUTHktrQjKkgt2hsOHg13pGqfX8Jnt7Xwqo40rYOblUsZHohu7FbP
rclMaIJhXoyNKljNcQdQjOMoo+FDYPDKo17OiUflRzzqIniNlllOF/UoOxP2nZhTIcMqvCaR6D+E
jYxgyUQGQ+fHXQKemfw95laY/RbPpFiGK5XUbhUUH8VigOpT76kGOuAzgdJ4Ec7eodVyye9w1H6k
p4W3YQv8BaeJ9Kl0ZcEITvLTaL1bwEE1yTCrCEpYQONCh5G0L6WRF+jAYj4eM9tvkgdehbAdHG76
+x+BdMB5umqOJtxd/xDvh4qQd200DfUuQQdvwHV9PzKPohWS+pNJ+XlphWvnvkw7hbt6DIOCZ+Hk
TXm7Dal/pj0MdfkIX2SqO75OOqAPK0pspH9smgOsovh0IJ6XPDjWP8aLAsMTrATTS8NGpKK05Jyw
3APSF5ecFMhcQirblUmYCe+Ul87zbcqIRjxWIwxb/OoWySxdygtJZhRaGtWH216mIESP07lZSbOX
yNTuNr7gNHoJiBkT/djjiuyc2ct5RSgpkabaDGhDCw71HKDjYuxx2Obj57liA1QOyu2PvlnG7Nq+
kd42/ngI5ryVGRLIa6GFN7wfFzXeFihFpqgsrxRb3D2y465312CEZEQ1Kf4qkzPbR8fo5+2PSBHT
xWz6iaLX4kSddCRi4nFu7kSDJ1MmHroCtc85fDckv7VL8YhmrMr2UXSAi+QP38eisnOaRqmRAU3l
QBJWG9s8WH5OZMzLoxIoBco+4yTvi78mJxFTpw7MkM6LTDW5ARN1ben6sag3m0z05XiRXKQyCWkn
OZjVMEMFxTjCD4Zo7z/mpEnWBV1aC9JRsIBoZuqofBfO24HKUDZhI/o8kaD2XmOvHzL3+b2exOoP
dMtIafMRa4UZWOenUu+tI3yq0h77YXk+reZtO1DqaNN1D9DyZ/b2sMC3UWiF2gErfbBN6WtV2WAE
NyBlyr6f7Dq/xp40mRv/GggtQwlVrdSLeS9E4BIUzjRpVD2sJq3MW8kprPkogIeSjjkRLShHq8am
jegu7hoL43LHW/4XNcodWl+ejKk1019pb3NwKcnvZ10Id8RdwOqG+hojvlvHG+kLxJBVgJ2DDJ4i
cX33c3LX/8v1zopkds0clra4iU9PGs/t0LgV+gFmXbdAKCWnBUdwue+xx7jbDA3ZpRc63dpzmjo6
9i2XqsuC9c0xXtS6TKNB/oAH/y0vFP4dvWMkYRRYSt5IKQ+Ar7JPbAKWZDsp6mGx4jqPc0PB8UGb
JiKBOP+N9jq8crapYHYF/mHXWZzXaJXrNZmAGSlo/7LHNonEpg7A+SNlx2blTwbnhFavztC0kr64
eqtuRXfVAMwjUI+HGaHVVOq06hbjnQK4o69Qyh9qsEk8GatjRDBP8DBAjoetLnE0SLNch9mO5EWy
Hs9XiZITL7WF6X0W+Of26hBd4zMuuSRFibZL6volxf3NJjtVTDduF8m7s56CYdtAu8m0Swy5Jyml
N9zvLWCBsHYay6tOMyT/h2XN9CsijXCvAO0OneLzGuNLpi0GgOMSID4Jg0MEaEc6M2KW30UGNA7P
KnalfRuWO3Zbw9+zE6DpX7OZwfh7KnS6/BrogZ9VG2/nIRINHzDVwzFhcwcf9XsemtNUvISz4gzT
fDpC4S0eDrQHNVmINkhZvOZ1O89R3anrF3NJDMg9fCVAwlf+GPJ7rkayNHlW4q2Q/FgnwHsLqrg/
xuXVGKb0gGf9zmbImUAlO0CoTtSj1VNUcyew4cpgGHRoWr4zdKUtOaRjnVy7dgQ6a/tZ1cHwu8he
Al7afP3UFSUREURj6FMX0irUNrxR8AW/e2Mn+ORwsMmsrypTCSycbrqnLekS4Oz0YZUr/nHQwL2b
wltQxh46vO6ejZuIYtpcsJHIA7K4UmezNUf0c7IX5H/D+p8AuqSSrDDLM0DSpaRXVWWYHlHYIdkB
V6Lz5fcw6xNnb3lSWnfcc49pp38+BWw9PJ2N7/YTHVDrtFElvcgPkcqPAA4DthgTdbK6Jc6guFAM
TRiyLXCR86Xol2/CapeIVbCexK7H+2UR/L17LMSWCpjEyPY5rUHNCKRQdeokkehkLR7VMZF1yotu
rqZiJX5YZhnq1WkH1rn1ghPSxaEPqdhRLjRoyiZNLdxeTJbRMf2Phakyjr9l3d76rdGfDYx2gEL+
fFgfw93mWUaxx2YPlBs+6GspNMC4aWYtR4OZijaaWUwzgsnRgQF7bg1MDH16vo0qsXlv0Jm+9kck
LxuZlMIrfjIuXSW1lAZGUs98jhv7+qrTXG9AVlwAcqMVChsSAwtk1iDsDMQxCEAahJgo3wuk7UjT
3N/lEEk9md6JXi5We/61zR86MgawTJ61ImLfVHtDeUtWoizvFc6J3vl9zPiZT4H+AH9tXnmqjNPD
SoxfEhad8OJRXFzHAXzzB1ffTzagSGwksBpwiEp4/kU+ugqyzrflUJhwu/eqBVS/0s8KOLqYbCQs
6jE/krPXDpKWvx2xI1YZrkEj4fk97KzQCdLfJaa1Z+8KunxF+8dQCZpOsex9dwVQ0VRwxq0SEf2n
yRWlKcQMGS90NvnXbUD7E6Y9z2tWQec91m0lDCuTyU5vLM/vZkyeXzCB/6LWElMkgKbWzZPa4EZB
2c/VHaJABRUKaffD/ziiSieQYVoubbDpZTDfu+87OODyfeec5dNCbfFZy2S45bvDPiXou+bAksfO
0JGe1SubZzpHJLqhJ+GDJcWSSR7Hq+UOOQXJZMDjImS1tSEbhPeCmpKmRQiPad+N1cedm3YDc4cp
vuZZWVCPu6OzOoxpY2Vdro9+3sE6R6ZPkgizaerEMgHHOMiUqFik6oZ62eRHI+xs8NvFqxZKHDjg
a5fW+jeq3X4jzszUUkeiWt/AZV9Wm2Arsg2hhKA94MxjSME+9H3C0dBYb2zMKqNyAfOx6a41MzkA
L3XvIGaWVq8Fjj20XroN+a4t3scJVEZvkW85qFIqzloJRxFMJjWJwweMCFljOxesF0g0EetTKwpq
2w7TKqRCB6jd0co6ZHY2ac2vDn97AZX7qOSiQsnXygaf9nKeS0rYgEXupKF6vu+mdODmClRALYn7
6Sbs9prGNswLv1rxgvh7sVV1VpIL1zyTmdFekKCshqTHQ5jCOzSkm9vLBL2tIwmNZ5psHvAn0xe/
zTP0u6uD87szUDOE7juOsYS+Cx8fWi7X/MwROMe0p2a+6DHIV/4N2IrLH6xRP4HD+WEHazGxXEgJ
vDlKLW303IJSFqvmxdkm8FhFo/fR15r4U38ZPmmyaeZZ3OqqkmPTOE4w+4tHwaTotSK8o64pa9X7
Z+cL3yE0xJKVke3zL59+hXfE5a26tjr3JtfPCjEOmndBgG5LMvkt6S4FAEYe1o1A84UZmAPgCEBH
GYFQFJKakkCeZQkr7pV9yCvuEnAQ1CT07mY+LTyyEkq6TMp40GTpREftF7TF2um/lbenFHdA4Rh+
OZKzlsj8haM+oGUEMJxiTttq8C8JWf/3h3bbIJFeQPE0umrwpE0szoA6/xCGEZLT/ifOpmvdJ3I2
oZ2WL/AkAsk7NIEoPKV6tXirvqx1i2t0iRLLQe6vCcfAOE8dfqssbqdqbwpOYK0eeVcyjklyGlED
Kou+a+DVwquFYofpf6YcfVDk9lpCRrqkArWv0u96E6DEeOBsIvFZklieMpVHBXQrjlRXG+kVPcD4
GBG9n9bE8yiILxnXb1QvLPNord1f6rJgFzbeyZg+77hoG1dl5Jb9CFzVO3Q22cc/fivBkHnxqhab
LMuL/FNTHWMDaGIf+ECYWvzce/jPWSGIxbCQiH1ye6GCiX/cP44UlUISgFuP/bNu46vSfDX+nrNH
ieebtE/sIzWG9SFcw5xAZoQ8ZtLYD8w7uCDyT3a2tN/N/Y1pS5NXyliGcJUW9PrdosFAacFmSKRR
VB8QLlItBHsRFGk+mfcAmKeXP9YCy74yRBm8qbXDRDFzpcqZtVAFouVGPXmCAnADR7znGgHwDdky
UMI8x00vI65r23nRe2ZigaehDfKMyt0rBSmN90jFDwr5dvzAbW4ytvQ1TAEUWeajp0tQBhbfG476
RlqQ27SJkGOnQdr7tgdb8jnbofzKp7WxijanmU99A1K2PkNmjTfJ2BsEiJykU8wsRGyu6ED9AC0t
jlyFbA0qFnVb0YrEYE+OuF1AqfZpaM2I1/Qw0S3E1fv9KnJo8q4+2mtKAL6Ie8DqCYTYty/mznHo
CyxiV3d7C66nApci5O/KAUqyipqLbVNQJG6eGh8sEorHCCIRbsY999AxKYDyiZhTeU3/w7/q49gG
PCJH3KDtB+odb6pxN9aMwcvsZStfQB+wdX8ctKzU5654mJG3Fed2bJ/+vn34/5MPBHPGP9iMTmj9
2HxdIzkbvN0VJ6S3AX2UjXoUNgClNstJoZFzQaKszNHAd9jgGUHvHZXHMYD0HIpeUfm5nlNoDG4E
Mg4ZVsLc7mbkoPF+e4KiqxQfUbTvyGo8AMVANGz475BAjSPHyN4CNsh4JKG3pH9A1mH22A9cZxkw
kyyo3wEbwYwgWeZH5lnHONzJES/3VxIVVVWsxOT20BUm71pHnuI2mj5c0+KOA9hbrHmROh2IS4cy
sNaYNK0l5QXl4aE/yVdCNjIr0iahgZqOGsJRMDTp7ZKGh+ZuYMCj8TTMfGhfJI58swVX69cSkTpv
a5xwAv4snOjV3OcBviOevs5RSrFsTs2Jdouk+c4P2TKuxvOKD23fRBfCBgEO9zIkMpHeg72qzV9n
oRMnYvOyZjPzcjG0dsLW2oTH53ZnHj27iqkarh0WBOnMiuEKAuujfQslHdd5NDRm2BxKWZWazjZk
XZWtK+bSzv+FFkw/6HEvsPnrd7Z2lUjchVxA/9v4kvCB9LeexdfLD/1Ez10SFne1zmrFGjOXKq1Y
KPsZ4lqfHL1O5Lbs+AHj1holaYvgoWlWmHxjKDawJ0gU95j75J6VKhdq2jLR0URJW8OBRhxpC4Ys
P7pdq1OaXLMge2RN7KlQlReA7jBuGtbDA4ArHSOkCTDBqZ1Ag4aXOw1/HzJ+X1syhhzVxIz88AjC
xvkmwwoyZsjQn4CkkanAhyDf/cpbOyyG08+dcqQ1Z3m1zFy3ictDZhrM56ZpkaD7M1CROtB3XM2s
n6kclrAbirGrQ3Ke1wGxE1Rl+bhk1e5nh0dG+0Fp3XVKH1PCtPIh/xTqhQt1dhPLB18FT3Pc27vj
RDEa1qeLqQiwv4pdMj1O10tAomWNIj6KADCfPcme0oDzm5EGDE7u8JlN6tHPOLviWktsIY/cq+Xw
ovYu+ilz/bhrxw7Lbvb3h8+M9gXrN0qt0VNlr+msWCBzM9yasGXZUq+wYL3zarjd/hMDEawr7fWl
1C8QC0APJDj+YkkVC6NhlingLDj8FwYK3CwgJC5Zdzp7OzdMxsN93yyKmtZfbNd/AkMBJJS00FTX
r4VUbY1lgYsneFQv/5hy1gHcuhyO2zQWrZCCSGV80hjnrRJNPrxWe/rtEJGErAps3RdDnv+ErvU4
TUVk9qOGRs3q+/WL4T8iVBLyYu9ZjYF9LLMaKhwoY4Fhk+gF5R6xBUcvtoh5l0Nc5xz0dyho+TEx
yLuZmGQKEFkkaQyL+S1LTsADfuft7bWm3T3ifqLuq7GZya3yQ0qB9I06JOttVHCRteREQVRoE8rC
9mg9HqEXXdvaal6IiX5k9PxInITp9Rj8q/sqkFZJKgrCs3yqFDexlokdvVZw6CAhZJ8678k1nujM
geciNrFRx7c4sb+mRa0wLCWhmAOnR/sXfNNy48hGJGfmfAMHb2ESFHcsMr8Mz9/1KyIc/yPJiCo8
lASFqI20iEUxMzftra2QddvO7xRiMsCu6sFYxnQoQVe9JjPveD3ATrq031JDBBpDUNLQm+DvE2Px
2w0niFaJnTDSWAnuGM6cr9UTDrsNCHGBfwW22XbjGidn13d6N4lnBcQk8CqxhWPD46Dq6TVn/KJA
XiwOpH0dTn81z0MRDcsaRYitYCRWsjILA6rJSyRzoyiuQl14bJS6Qt8ZpEAQ/EZ0jMjj6hKXrx8v
8jxDqdx2/a4J7uqhQTrKNqzG8xSJBtk8allEXVWqQgBqDn4OUyZMU1RwwutZT+XPin9zpmLKmttN
80RTHNvg/YylzApsALRUTY2nR63SP1i5aAGrAbH3OQKXG9NUlOCOTMgTHc5nvBUGNT5tgKDl/R9M
FIWOCa8utS2+EUPZmm4452J3aZ1hfRcV+4TxUMXiATve2PBkrhTM0DhbP3wmGRJxXiDNgBDt1aAt
V2xq4MB/Uin6I3RpEP9u3hTkfj8OqxU6Y3cUWMQSggx/2O2es3NL/UBg4Qf76tv81fazKtE3/uWZ
t2xOoxm+6Yc1npDLMkH0WEocsZ4jKEl6JGpPG/8dv69d4U9ssXlaemvlf/xYfuYHzeCOGttKIpBy
ZFh7KRqRA+jTJw+eko2Z462/uHUW+Zch1P6P44yCuw8zhBMJbGu1LZKBWBg4PVeZygrVJ4dKsxtK
giXX4rpS6c8i8duj5T8+YWy6Yz5o8NBukRDPvxjv1wVoP3oDz3iGWN1let1Joo20aDaROuf3otp8
ZXWWMRrYwHm7+fvacLQYRtFk9jmnTXbGS8MpOH9i/u/wb7pSZqgLH7miXpY7ECOyuM6q3QS2wEQn
wGUnMpJ7unDU5NE9fg0iE+Uf+aianCiguN0TdIOQNyP7qbJ6jz8UmXSLWSjYUgSTuZnfT89ohKBJ
tWIJVklLjvcY47eMy7N5PtTRvN8mVzUPLw111Q4a25HfeNbkPADXN8Gg2y4W26ecOmROxlcBCRhF
kklgkK9yUCs2VdbcV91m92+sqwn6CFpQcyoJEL+4jF53aMQDvpN/vx/kzi8MJ6b6r0Se9pwB6qdR
satUy9+R1Ft9xLyP9CHr7IshCyVTCHMIo8T+IuPEv8wgUFmRSnsaYiNhfH68eJOwQe/ciqO4mAeT
AJllsdbpPjzYF9gALCq+BdzZcTMnlJlbBSGMD3RB8Z8hvxhpLSn87zjIRI9dZyjAR2oYHxM07WLB
UGuqatEUo7CroBt6CMvEOlp8paueBDL3CsN/5PFW0Uh7KfAQN6JCSifLTOtdVuwvm5r1jD2UbxC0
hu0iJEfwVJvHqYi+SnWjSSa1EP/wS6uzJbKpLLM+NBGlLTe92jZE4Hy5B2gEZLrMSPr5uEz/FJ/0
njXC5t8hDz41WU4w4hQfQJ4eJJSbnYvFU7CwFXgy1fLs0BJF2tlE6dwd4b6AIc3YMTY7EdIIW0fl
O1QDX7i2IAXbsP50ml48EeD+xHCRgL6Qydr8syPUTMuMcBl9R/eXiyZrteFYgnxPr5TMRl3kV6Ba
8n4xBaC2w0BRZ0V8pbYi60SP7htRIej4U5z0klWjJsirsD3ZxZrDRQqX3hsMLzqOSsCqI89QOewy
RONIqLDcBgvfGtH9PvpHXLj9j/ElBUk3wWJ2KtF/1xIyf36O+3Pky7w/1BidQOulWe2lzQJD7rec
Bt+rG/fDn3HjtUoiUIgeOgh9zcw+MvZRyY6GJgIy+rNNGKTXSFpqfyiz1J/gDvS6UGObdFxuoUbw
iy8+BCE1je69/0lhTaGyP5+vy5PG1MYS7/vZTJGBNm4PQf1mZOIPvBegJOBkrqFGGef/I6B5kWCI
GQ+wjBReUd/Ff4zB1Pe7itYsG/+jpYaUIPOhu3u/d+JKcENagLq7O538oR1M/bRbMpqHRSHbfPnE
kyAgur7nteT3lCgNEh4fGyOUIyGIVWov/diVSFK7DyEjW1KnvmLYg4EbSmFMFohVuHZXhr2Qwl2a
5xI10PJEdAnoV82VoE4EhIIQlvoCjHphamsXcPH/+g6RukONpNje5v0BtmTgBYH3jMLcnpqHSFjA
84zClblLCHneofN6jGSsLUjOKvdZF9c5unT19jLpf4coEtK0qMg4pS+GLYIyyqs4bJuUC5TXrmzc
fbxwrA5GKQn80Df44X5YezCFXKpLg3mQpOc7kmi1+o09RhKx+ZcFHO0UoluC/dbbVQencqkQzHGD
wU+vs18kxp4IV5KV0MDmYaege3mW0WfSpLYx28CmIDb/aDyBEJKBRJzOYvw8Es6lvTvAPLxUKZDy
FLm9hKgddogoTqqyjG0yXr5yT9wle0Cl5sBlqor0RqSS4N9gUqw6nR4B/U2Qvljxg9hjsNClLWSy
3nA/ujmu6cctFhBbYSgvtwDrkR62nMquCE6iID+wga/LKGaZyp7Bzni1X+nLl0RbA3QAbQfH2Hse
Ubnv9GjemRupsqQbVYdDX0BI5ijtcU09areKkZd5pioN/CCB8XSo05SZXWQxs3YKX4I7ddi68qON
3vY0jpoLyzPb+nBRipE4yYPfHOtTdX37uhy+c5xOCgaR1hBZB+r0wHeyu2LA4jjxt2fBDS75lc88
tloH8ypV831xQRAj0+YqS+cXLfUkVuL5mTZoQl8QoEZZ06Fw0I2SWuUdh/y0ZFyTwkw+MehldY8z
09yeHSMV1FovBiZLmn9g+8pmMIrie7Xn0Rl5rzl38yFAq6PTQw/XTtAIwh7bNRdzJJJCp3vO0Z2J
LvqS4z5YW5/H+BWWA8Snv8rGfqZKt9pM90gaLHVPm8bs8raUAnZnG8GSE7UuPiAHPkgxR0dfCnQV
chNJ9jSUFhQ9MgunVfsvi0NmGfAcNnKeh+c9CeT8hSCTeb85wvQRIigJcIxfKGcNegxNW0DJnHHY
SBzhYfYPF/p42GJTSkmzyMQhtsub1C6qXlBRPlyzSEJ1+EUmiDr+5EumGSVVS/s8nMK5AF1lkteU
dZ7F6+GLLN3lYJJG+8UBNUY+RyZiYzEv03GoLzymAe2cBD21KRMchN36ofozE1k3unplZvFECcvp
02dwqZDXigNEbwsG9j5IA2Y1z2wasYnHiChRGHEqtxUwrfthVY8254hNNJRvMZq8kdWcq3Qgqpre
zWFjR0p7zE+Y/lVIFkh5uUrPY8rs34ubRSyMjIRfmN5WXp7jXNSu1vtOCeOW7KAhHoPt3/wXj7zT
SldKBcAvvjcyD+lyNGLAwYH+pjMfdHmxi0pyNjhZd30hGC1Eh4naTEqNFk8IGIzCj6SuunNlYqTb
hy6AzKPM+VBPJ7rABBwM72/3L0A2M+s6Gy1tiLkIGPH4mM5DMp6Ny+PigF2qa9ij6uW1h7DTzMKr
BFhnx7uobhQ+Ht8hIBut6snWCYHVje9eDCgVpimgzySCHQOJNnTBFH8kShtnavSD8gEYVnT5CCBb
oWravjE1tZg8eep51a3Sw70PaBlMWc1bw92kW5xZAF1U8zqcXTmlAocEYw0NH2So595Mo7iwfngf
WbA4jQzBgM1niGXEhh0h2swq4iwMezFOHq10MqZLzriuqoLZMpMyhAtOVqF9JvkQ0dFOyoZJ/f3t
ABzutOfaIGfqFoK4/2jksiBF2KMoqPWaafxkQy/DsRBIhaDqtZzzmPX+1i6Sb5lVtEblhGpVea/u
Wu9xWOB/5rQINLhnBdzgz7IAacJEbIIqDfL0OztVeUHydV1Eo1Znr3jWdVt3bskicTgne1xxPcTD
yAfKfPSAgBnsz0VBVjOzFX7DiJJJs3hd7Eso18emu8Tv6yio6MeHIsxAyx68MgwjC8y/u4nBsDPi
qMAhOiu+RYCj6+9b5OcSBjVhV2DyJjI/ANbt69rFutqljnDzcmdY9hiTsmPjMU/HkLwX3MO/SCec
hs5RvYRJxyMuJu1Jt9SERbInFLyjVwVUKcXycjE6kBUDEg1lz9BXFxZIxJ+dnNIbaWhtPyO+RtCR
14W5YHUSmfGA56P+pnn2vhQbseKxZj39uKEjbU4EvudY56bm+07mvnk2j07R1p1oxhPlx/rGqA1g
l1V3S9xl3CfUlHNfSmnOcE0+gjV+Tt/sCR9+iBEcUSGS7GQwbzSgB2dYjRcnKNJDyy6SuyrMjUcd
r/OUf16dgJWlNvj6MPUuRVTBTh5jbF/c+PEEgxfm3q9hIUtl4kRO4WDSIJdXKSM37kSBeQxPpQKg
Xc9SM3nf061t5V97IM5dukSUbAPXPdVdoSHjrXbhMlPsfMDo+OicHgx7zKHBtTryUQ8xGI72JhR7
jkgCtIxOhDprSlsNa3BuLafjU/4UUrz8YD0RqWUVhT5M+rVGNDptYgNOGIT9r1slk6c9EZLIWsCJ
UzGgRO6rLTTDlnxtRaHKVN0+EeQCcmsvzWVDKVOYtIyL3q9d3ST61xojcc7pP1AHoffRH/oDnDz6
4XxgEB0+PA6Cf93j3H4NfkW9TuUliP1iCO1vEi5Vp2CYmZq3MjAJOoF57NBNHXxi9eCvB8mR0rwf
vgD03banXCw0mbmC/v1VupSrlj/1jWwbHeHHFa6nPuqdmEptRoHJW5bpfjV8Mnwr1J9D37L4jA0E
FWQ+2g6Jn4lOX3NQWp8+BWHWNQG7p5ukONzC9kMaAnT7wVCp6xXSoevZxE0U+1Q2MKDGS1mcSbCD
6Qy9GcddQGXxEpxPJ2RIN+Cz2zpZEsQ0l0te6o3+Krgm6/eiICluq+KWI5Yv7Z4UxzQ1rr/o6YPO
n1onqeSXwHtnlT58lva7rIFJPuiZ1SfmPIM3uzoeb2cq4YgzYc+gW3BEwJ3m5XdzQ749PHOpOW5q
mUoOvGSthoNHE2N2f3VqOHRdv7d0f7qOM6bmzn1F5kJsoXXWj/E/HQF9HCbaPMB3tEt+Eiu27EpS
Zk/gRJCyy5uTZCuq8pS26ttCv5yTcGvyniWGmaLufJKot+yDpW1GrSNRODpLXbchMGWGCftXsTlX
ffPEEkw7iZkV87PKNQNCrFECjuDpX+DqX4kCn7Pt5941f56CrhpzEn5/Wyq3dIuvOzQOuO+1YYC/
20wxvsVwLgnIVWxSAB37fxaxt5fi3OIZqlB1tKEh3afTN42JQHjxhY1PKg4Twg+PEGoVZeUrsaVR
I0xrWJe473aw+zw0ffelroL3QlOO16xrg9sEXQX4xtEs39IPRec8HnJ/bC+D6k5NX1yM0BITWIln
MLWpxv06Vb9hIiKcKTELbJa5xJyRdkMfHzNrDnIUlSnaE0NW5JbKNicj9cVZnYXkHODMkvS4kl6Y
lyTbGV+IphahVxC4J+maK1SoPrlxG+o/oIpLZz7+yPguRRhVwDTqG9p/nXx6fKGJB4tEeMScJm+G
URAK0DisgnLN3zS1YGsTZ9a4UrcZZmtAv5jkGzYUCeDWutq5aGeczsGKjLsaomSJCU97wUKGJOe7
HS6iTnQZAe/UaItH1mrfKfGSFIkSaiqexWXjZnABT2CUzMxJ38C3cOWClPd+DUKwcrdDTLaEkXDL
qYy2no02nZXCvTAGUhfIk4zPdAvys78yWTFa520o1hRxIhWq98kqU8IWB1wf9P0SRWNKaC2hB48K
V2++lx+h1SsmBkrf1sKq+gSwI+FHjwqnCu2OqpJpg/XQV58J6RuayNwz0EwXcRUX8br/PiIsdZ/u
h1EIXHFCoec6pJwSez0kQ0FvdIFSvCz89lxGfxBlz8MIAZVomuYGdWonf21H5CdFb9pC+9de/zV2
c0p6gzmggdOOS3WI1N7vEdagiNY/CSIYON1w7/kDQiZ6/bFvKh5hpzOdSgagUyXtvo76r34OHn4q
QFEZItBeh6he6XRVN7HgqCHv17xz+UKlsk9LOIis+qUauNFtY+TSTHj7vuIYCO1ysDH2D8Vei3+U
Xy2hvVx8VbSJxnxaPYidrmnv1/TCp0eU5US29Q37j+xVrQ2CbS6DA8b6MoSruz404/6MgOztHcSk
3hSMW0PwrV/zCPrU88l0ZlwPu/ShtJObk0ImWjtQWbj8SPCPOtUzDV1alIpReVnGMJHoNYmFAQep
AGiixxnT63+Pg5Pu33ImeWy2BbVXTPiHposqJMCNv2FZ4DIVE38E4Kp54k1acvStPTSVirY4pLz3
p/pALh56ye60voGnqcTtKMi22OCKpMrL4K25LbJ4KACtJOjv2A5uknpHeV82jMP8RRQL+Y31wscn
yNE2qwW48YI90S9qqUq6ZWiXgb660a9/8czl/5Jxg9/ILZtwkHiV4/8Ss/jLxPLyefsxVIZy2ukg
zj75SgxkVyguNU9Ca0UdiU/xkIP3e41OK/pQ8Gqs2t6u5Ru6vTNMTVzg3M2ONjUZbgo2uGNOsVtu
csEtzwcfkx2b/fLApgeBA4d3oPZKEgRVD8j7B8SpmJbC2J8wmZVgGV9G7GSXDFBGjGAjBkZ0vyD0
t74XCDe5EM1BBL6PyK7srhR4wMH0scuVKzeXTY0H5oGrf2GlMDFaYXIiLW16drTB2sVsVgmp1+VW
PTG1N7ErfFPIiPj8IemQZ7KkHdFMxnP5xzYXd0rEQKWs+Q30a2vq9JV0NnVouZPleGeSt5jPrB5g
DdYOw3HbRNusZms+eay43ov7sIhfQPTcffXgxPeJY2H+KEb1XrUbNebRqpUZA7ZZ/wgO+S+zBhE8
zhF/AJ4Tz/ze14cyEfC83m4096nIMMmLmjENg1hYF85ojfeNr3Eb8bv7MxLiCr1S2Rz3cigi86Vz
Fp2OvSmtKsXiQcmN7mMzwMjHLWjeP882ruImcPJU7qRqwxpP5QgjD3hOe052Da+CpWK9prT2l+PA
lVON0ryOj3Qy/BwqvXbt2UQ35tjv79Fp2N9ZyPeHektE/1j1C7xk8ISkBdUMJhtPqS9s8dK4k2mR
wMMi/Rxz9RRTYjKDm4RITRxs5IDSS6+JM7vljfnhns9dPGfH7xYSU2OD6xY1xACspUiDs0zaPzjn
Kt6e52p9jGEnbCicxPZLxX/1qflCP/boSLW2WWzCvYtpW4FQuHttfQctzx+/jodzoLiWBbEyHqs+
V0MtFY/UKEhhx5M47SDq4fADvGukd9aibip+tfPjHAJGRwreSAVxsEojeubXySIYgb2gzgpsujOe
32ytH6iBUHV4vuFgpy2yOD9Kqut5jWpErd+ubU3g+DCN03/cPBapftW1c4p2aE49mjZt/W68misi
6M+Ju6ZW6pp0VbzjCjixCI/f5mAqwjoV4cxNELe3yFPgqi/sY+yOxgIVWRt42w3U1BInAFy5MhWi
xGlRhoK0W5SUH0s7Y+2Q42vBBXubx6ziYaPV8J7kH/cFWHWJodO3EFeL4KoC4j9EXbxtT/OOTg5A
NtF1e2zB4U32FZ0ObyJN2CHeqPZKyjZpSlxzWfj2tf3P9H5vyXaMzElg8yu7tNaxjGHjUwHnG0y8
dcOn92yCI9XXGNXWFkyryCeLU9Z3KveClsqbDDkVT0YkWgDj+29fwOasa6d4aJRZ19jKRhu+uxgb
LGtwKauvhBi17DTs4uduA2DBcoDajAnDspNjyyYKdHk5OfIcMQMlukJbNmIzH4dNXbHVPnQtyQe4
mw1Sjjg1SyIUb3AseBmuUa5/YGNsD7kv0sJThl3wHIrbgufNm31++YI5cVwDiFvrBEBOZW5lFIBo
dOYR/WbrVYwjkcivxdbFPt33QqiRQsvkMkP10PzqtC8hjzu3Ic6YXEbE/5IgS8pl0xDGGWLFSRYI
H/JxCPr2FP8oQBsMxrW1MiFGSPZxazXNPTxJvbHft5FdhT/rIu2avZmehIVaez06PSgoXR4Ect+u
I+oGUOfHkoYZX7d2Jw/5I5XDt6SRcq7GD0WSf07nxto41TtFG4OYYfS7nK7qqnYGM79zlgwyuby8
DS72ugC5w4BuAfVlwZru0aZZGQ1TTqq+StlvNV7oqb5eZQTrAvXgxqhG9tz6w6TGEG/IoiRPMuSl
H1OgwswkQzS3+iGPs+/McXB1EmZujEylmAK3nndgOWR06rySXNMSteUBfHoYg4Di9Fm1NBtpLNOp
YXCgYLqGLMDxbtCIqptF37WOVgI5huWO2ebPmfZ22vFskww6PAjeZIq+HGIdxk6tDiGCJDfHGLkU
dS/j6Ea8hypbMam5gzw2KgZ54wztOJnFsPYMPm7qzLfyQdNpUv3WwmVgX5b9/IUDyAoWLoAe+qHB
vGT2x3M2/b+efmhME/4F38hXqVJqT33JUi6z5lZoYegEYGY0/5hZav1nu581+2ImdpedzmPVT/xA
HDQ3M3xxcOwxXqXN3TLMuPIP9lkfk0kZtrRH+w5nNbbssyLkGskNGpyh+GvS3QBY2l316kZtAhD/
ueJso/3fk0TlXhN09GjqlOWgSqjSuY3N15mTraUbUp1tz2pjcLh0P7Kpspp7ZcHWo7woDwL0kzus
bvBNv687vvumGHxkPpcJREDSUBDCRbQ4g5D00pygFhSJOiaQPjKax9M+AI9aHA/wSUcX3FN93U1l
3PA5W+Lr4zI4hSe9G7SPC+fshODSUIRjvAwIA3b54GGFNyF9pP4XfB5KiAgIwpGubsvqFCYkKu3P
HacO5l/8JixHtmrW1REwgc8fXQ/90XMgKuHNsadvxAzgDaoDt8Cqtuwv/fdrlzBXs2gR5a4IkNU2
prkZqkqbuWYT19HpJk/FaIMxNhI/CIfv3B3oSFe3DWFTGmf4HeNdKgaBFrWUxOqdnDjsC9RfppRy
GZLk3e27w+XIUUx9CTJaXFhuxSI69DU4ePwliFbf6ojq2+NakxLj0SACMr26JQvdjQUaFmGyvMKI
0Pa1ckdR4GVqjkYDuVoiF0zqEQF6FXBf4dUSscceaJRQfR9IDiH/52+LotTYlYRbdlSP+eYnVcmB
IM9YDhTo8d1+JPMhptSbZ5MD+tswhkSeGrie4NdREKGsHKPsTelerFHn33iaMlhlyFSn323IkCDR
J2rLCvHG0uXsIgkX7CT5R8bzkQdkJ2MQ1exuSHPgB8lm3tZeQrPIBTLuM8fqEsO7ZB+yRsd1Sntb
bpmUW7nGhQZSR/uUkB5J+FrC37y2lIVjRULRbVjRBZObNqKlVoCN+s3KxGMEf/31CDGF7iefwd7Z
DwHDTuIprTZOZjVwpb7Jfwp9V/IxES4iPJLHcGmWFDMsrrE3L60p2ple5rNdg/euUt4Zmhq/z2zB
xi78uhju2AhBudfVkBEk81AgBbJb/C2OofEBu5N91+M+o0B4zL7VAvJGroXXYJoThHk5CN+kOGND
7R3qhiiMr8nfkVTaAglJ6/iCKLXT+KT2gXnRCuF+tbn0xODO5VUwGoVnXefAeqZ+3DTQiQA+CLMI
+Hyw320EQZiA+RKnCX5f0cSrs3I9zFxzUi62oF7Xa+61KQtfY+eiX85ekGtPONdjXTvPZjrGjCtK
O2Nx78dvSt7fp9eYfhI/7wUfJVy6ql32VY3nyhPCHjbfN8+sR5BeQNeRfVhfNBbgm+V7wXhNo13Q
+6jCkDRsTZ0neHGa7fI/KTrXE/l4ZchZGZNnoBIxeY7V9oIu5/bKYPbE0sPcCoLi+zAWVB1NOZPR
iC0iX7ZJhvqukw41kNNWmhBgReDSF1iU638MYJmsIyQDdhZsjxxhj9luSJBMQ0q9GFpiQLeQt/+e
GtPPYt2oI9swS8WXVYJtjw7RMzFt4W7RxB4CqOZojZEE0R8ZJ481ceAJ9lQBvmqcdiKFhbp//dBD
NF4GcUkHIXH5vf8GfEn3td20ISm8xaW+dLyrqSI0KJNRl8vSPtZWRckdquWQ3UZp9/o2/SYcYSuZ
ZDN0eZ67mCBGLtXwtVj/NsThz78EMGzio1kNmTIvXW6HcerUEoNX6ScqDdog/5xu4+FaibrF/45S
fR5iIuK+9373Oaf3uNmztnUyWbUiGIMSYejGv5DEkbMopayRvvcFiYqnMNOkRVdm8H8tI+E9Xc/3
Si3GcKZB2Qjvm2WiDagKCS9mk5E1WLetKOMRqTOR4RWIh/ECTQ+YIV4lg9AOYI7aEcCWvyoEDV9j
AZyyIxS55ZRTBJjOXiBmlM5q00Ysx+ionbXcb++krMPYNXHKpWXFM8+yHpbr7DCbaj9GsdJ0GVqr
B1JGzlAMSGhkyXaNjzueDGXu88qDobnSqFYsVP+WnaMfZrMwdzoIf5LjaI8UKCUsgwIF6yavo39C
K/vz8ujv/IYWcVChbKnW+OIoV4St8K1c2ybOVkve1ahkDH9FKr0s9TsdhIXVwjMOL5eAGxvnp4/i
OvXgZ9OWRC1SlEgWB5I9gTaDVuNDuv78qiJD9R7YIs6BzUWTXCAt10ebZteLRDQ+HKFokv6+ppyG
5Uv7IbjbxfWOVDqMuddzRdckqcF9J0ucCjskvHpjY6SksjSTkC38sxkBBRkL6fu9mlOPfK6HfmJC
vKtssGPuMR0yok4t3wwQzXiOqfi+FZBHgBKVrT9uOzh/QDLORpbBG7EpM8p2sTfbTYJWYJStU9x1
6D3VFGoKWB/2cPPqVcx4n/gczlKlvOtT0FOSVJChBy1N8m1y89b51JeSgQq9F/NaY3k+LFg7qHDl
ynhVQlv0CTBDgRbcWBE1C54KiSlcbjJrNz6q3pHuRMppaJc/SgVftIPZ1QCPVVCRI9j+FPrKh+1s
JuaaImjP+xiuiNqw/K4GJuHnCtOLYdB04SAMA4DGBuhIcflOgrEsSj0gqwiw3WXkNEeLlOtM5G/I
nTIxrDPI3V4kLlQ1PcKbWbZ+7F/O21zNfuTd8bJ4Lt7K9sGvQbc6mjJHmogm4AcXLXjq9al8sbS7
F4d2esJxnau7uqG+7CmjQYEIhbyN6bvgoF8C4OGmiZFkNzp84EoKIGxDrmphzTZwTqdfRbKnRVxi
xQVutaKcsBHYmL82ligqlSsqhK9LuCUEkqgR/qu+zPYOO3AwksjohcG7Z2ABeSkPaudvMMQegf0m
e5WnyCGgb5b9Hvosp9m4gtM52E0JRYY0jM7afpXo92eU/UH8rDc2iFV7B6fMXu53lnAtjucPoj4c
O+lgI9Yo1YQG0jkDUlZcciFeyn/iAhGI9bxdv+cbka8RiAFci0X92vefzItfRglozDuzXeognc+P
W0Nwl2qFFPvR966AdHkqw6ObWaKMg/nIF2SNzwjdr9R/pAtCWH97+djD+9oxWYwQr7EXCxj2qXb7
T1KI+HIhrTBvq32E6wRYt4+NRze7xwrdRjZn5eJ4v+Ym+1pw2BBELRXXkpNRVvIbrfkOMDvasHhF
lMAVxVPpnDWueE2wsm7rRdCOwoUl9M6Y3xtZWLrBLiQoRS03nlLeBrQY0Yku1Cev8pxYgsVbfWXR
TfPhqG4l812eIbfJCEZEF8z3ncElnDDMig3TvAg6IEJq1t7wFORa6fFcXuGqr+xAQJucgLinRwJX
QldepqUQd28N8TJrnsIX2htyWGTmTgIlu3WMusHes7CFc9kZyrIZUIpd/PrcZywR0oNqS112wGs+
kksYs7B2yLXGtSCwsexkf+madA96R9qOPgPGJ8wg2g1KLYttvkHytc4L3mpGLZn+zKAITVYjTMbU
5nD6lqEiS1ih8HSBYSi8g/l8wV+/98egQWj+S8SE/TozgC7fi6j3fcQcdFJ3vjl5vSySk5q8bFqk
7Te4a9Zm5vkrxMwcG/egVjynGOEc63jTfWte62/QZE+ghwa11GRz/acHGBACRvYaEzZlYg4lWF7X
5sbR/gMxkB2sAiXLYxULpxFhpI3/Xr3//zEt675UYFJHWMH0Ly4QG3nPJ2ur/peGf6ozVG3jnQ6E
jZoIRm/NEWPG2wiGRHxcCs9lIFYgLQFMZ0rEV20JvIEj6hiTVo0j3Ezo/R5bj8bRlVzWxf7mwPEN
7Ss1KztlLbaR94oneD/FPqr4KwOPgVadfHegGhWeiVwlYq/hOELPTXwm+iP3Or7hEeGYQOgYAOsc
dj3tByJMUmNoCxzNi7EA9nYmx13r6LpIFaZU7Sg/uRJTQdR2LDk8PIRmEwPjUmt+Is0T/1wT+eXB
RxGAwK0dLD3+k0pap2mFz1o8787PS0J63oCwv37BVOy/w6o//jLGwuJItDdRtGiyLOAMeoLh5IpZ
1Z4PYE5slFiM9TapDNYicMba5hBQXMqC/H9at3fCOXP+gPrjC1RLgmZel+Z8YKe4jy4L99SzPnqC
EXkH9Cpx5x3bnsN7C6rZhIF8SKGxs+H/CDrO87/NOwlU6BvGW9IdMv8zMjwTCtPY8vYAWb2rC/Yj
AMQ8xXt3mbx0heqGdpXDao4bFJBanRCj6HEaNnDuUTaAztd/64tMU600/nyFZw8/OWTq+EW+5dYV
XL9sw1PN1vYXw/FykFZNsgiBOPMaryapoMwzsDcJtiS/vR2i7rIlJEREza9XkU3FIAyVzpffv97I
DuNEYJf1aCW9M4s1b1+wAVenBQqjKcQIKOM3iQknlu91w0KCnNYv/Jh+hn9fpFFbK37hIu4+GaT9
F4FiKcvMT9lLKeKh2I6S7eWZlJ+mYc4CltYTfwSjxQWnapXhd0wY0Y095qVcJUSqLOS0GOMxBG5O
6blQhQUBSDpOyK8Yc/5WtDqI9KSag9966wtesdLpCMAZg0DJr6UA/626M6+ubdn3+OLCPx5QzSvJ
jCnu7EYqE8rxttdHwMXNfWk/EBmL0pCrIYuFeaerS/GnJVQOeWeRKZtRVF/wrkIo1M4zHrhs8Izr
3El8H14p7RgIjf7heT6ZRxNwjGvjDqgvUTfkY9RrnuSsotTO2SyITuNnVaO6ToqLHS6uiucBsw4x
BE1z5D8rBXwrBudrfVbIAR4m+jRf4iyDCroAyryuAwaK2u+1m3ayWygvRNYjN2Rt/aeh1vwwHM8D
nsUI9rimZMXJxQcl1xNRgOLYOdaAqTqMFpoD2cLS59S3ESwrLGMjzy/fVFsJjXdfOkZXhIfor8Dy
ykSVTEZT/5OAcu9rYGmXja+H4JvnOHd02uFiwTi2/6VAe8UvkU7JKIKFeJnmsRXsDThpmqu4IFc2
NDmi18Uo3jnPukPFnLfwgvG+qkGqY/0bEwChhyyXYKCeSdFF5UKgtQd1jBSlc98LSKSJ+8fn3doI
1hIKhmuHFoVchcglrhWuqH0ETzCi2050j7SA+0vaqOcswhHCiaUgmOLTMZ5M+wcxA6D+i866U0Ut
KN1V6wIiW95hGnsxqxpA9cgekcyqu+PwvZXUVKIL50YqsvvxXFr1gXzzdi4xscIiYoD7PobBu6vs
z8vOQPA6tts3YUyeI6R97Z+F4p/L4LfOqta+AVlag62HO067MBWdbmbaHhSVRNLRWgbhlF0yKOhN
2Qt3n15Jf3NrAl5VQWEymGjR70rJAL5Tf9CXLQAEt1E58+wggROvr71ZOyzwYU7At0H3RDtWoDeD
Miz87SU49r2blSlIGsTIoA3OJh0CyTfnqLOktnmPeMJvI2DhlNsUwtJJoTQjoXiC5lbWakGDFZS/
HQaZOocZaqbnfYpdEWYEduHQGY58RoetndAKSx0p90YWaGCikxeDr0MsjpAsbIkfKR6Y4+1hw8kv
IZjfLxercPCYTjUbsrbbmthuxGoAyTuQ6V/hLntlxDmYfwrgseOMVpHrZMrqVbRS+X3SumyzZECS
9YBResDX8qlQswWvd6x/KhODyBQWf2vD37ICVzMQfxujLkja/jLq9WQdIyUS9NR5lOY61mVly149
Rn2hH6sCvip9rE8vZ40jrm+0h+aWXKzjOu+a4sRJHUom6XyGqY15jCyjigcbEXmhFavvhJbLtGnf
TA36EbtkJ07iwgzdWdoprjaN/H/HIXwso9S2QdVDur1uKc4BcK5UNE63epkmfnnw8FJuVcdwfgai
IgPvH7/qU1woVcwjWxon9QYQsfk5vOEtQC7udZPwfY6v9TlOQ/lXudN7SkDRx+VkZW2htwOy8mcF
PS9BXWsBETfDNzftkkNXCpNfzv0DCrzjfhhdJOJlHuqivP1Fo6Ju8Z6j7miZf0uVv9Jj6ukGcEtX
ZFafxMPUsqVk8k9o0Dnw1DtRTf0jTNIeJoUA6eFPC4+m39CyIAn41MqKZ2rIeU0yf2auJDKHmK25
OXoQu2WbpVXm3kFQg4ztLIuNdUiBTaTko3UojdKgfXLGejBbnnotb64cGmM3CrDeaEbDP/vVgHQ4
Y8VO2RjhtWkSk6qZHfZd1oDCChIyUNKuVgNB6/5eY24YTI0Twoud8sL9LuamZXuQPXk4yEV+VacM
Mq+8m7oC3r++rq6yLONrHCPLSu/pbcPfZuiVxdxqT6vnuhm38mR+aXN4FWf9xHY21n39rWDOo7Ql
LyVlLeMvpzilPMa6dBR4PKSqHiReedePMVLvgANOkYC9rn/q5pKF/x17DTDugwU+zKYkZxACsrb8
cjYeB0gxnu8UeUr4f2UK2VXzCkYL8dJzUXsxwK5CiD10A9zt4z0faULYU7aTO5p1F+IQSscTJFVC
JNk/EQMm/bXY4XoSuix9od20XdH0TmFLZ95vZTKYUeg0Nju6ZAts7h11UOzZH8HW5peBl4FlmVts
66foaXCHTx/se9Fm9PvbeWDH1MsUSZGRMPxFOGqvCbqWPvpC2MogVyN2C+U/TbQ3txyV5Ii+Krkg
4VJ7UCQVArm5mBItu1mIo+YXw8uuXCoKOEi4qd3qYTe9f8dNsXAKtla5CIcN9E6A7C1lwXv7y5v/
pD1vDUXwTRAMUb1GQx0v8ReKOOFNhEJruM2DS3d0prgiYgC5yKJULW7zMy5Qq0GBizgBZ/VX2eOO
Su3/+1r+g80tofGrcfIYHI4qGl5fsA4G7Rx6DmSRNmjmcmBPwm2/C1qsH1ySWJ13rMLuYmIayD4M
itUoELfgMFE3e42+SkzuA2hs8yVfZmidIUguAtBqHmk4oLEO7JJBXzs03H+lsEF6pNi8K+ORfwby
ZZz//tmpMTO8oSbvTMvL9AS+xEwA/eJoyvY7sNA/JddbqI5OfBxFa6yBhm6APvINCfYvbPkpmiA2
n/gGl8HJxOGN1HU4VpO4WWAKTBNofgv/7ne7cw9JMO70V6iq6OZHKrxLuYBPpZQKoPccA+EjCxUs
590pRszspNAOSx5TZZQxEqEpUYFy5fbfez8WLJJTYXRVyascgasWjJpFXZa3Cjtbi7j/SNpYhXgU
CFkqP3eRzPnFdkkkHBDCkqdfi3DTRJtPSO1EP35OJiuH00hBmFGvLWNQufpc7i21pQwW5tVFLGGO
SCVDNloWUOMZVaCI2olBtfClwLB48iAls5VA2hf699TLeP+pVLihsZkLSMxKsTeVpGr9M6JCHX6k
NTIxqYnAnxtlhsxXNyAbXrTyltN3DBIITFxU5ub+n85kCMoSZjYfKeqFzwaLU8Ewgq81FM/EeGwJ
B1HJmu//rsK8DKNvljDoRoLtVz4TAdISC5Wmw4G0t+LZpVlowbQQSxrRFdPNBlDmCNPxg33Vtggz
XbP/KjxKCmlSs56Egruskg4toreXhRvtvKIeK9/qvgi/WXRRwdWy9eUpzrH5G7iphBRC4lGDzDfw
Q4peDeZtyDOx4EAZngmDgg3M4O8W8OxGXoay4x5u9NtMLR6IHUWWymn9uiQ+OorBXNO3lEVPppLh
dLdODqF04eTpDfv+Vv4calVVk0B/lkEwuOOdivcSd6uNLxuRfY72XxhmPj4JNvxG71pCs5XhVv3n
Jrx1lwianBjOhyDrsIZek7Mz61sgK26RX9XCDYyzfDGpX2PBDGXDrOdPIS+4SUhFw6EkvdwdD9oE
Ne8PeSD8ISzLYj8NhgVvsF88W9U6jqTYZYE3SinXc5o/g+Puvb3WRXY9FE2m6VTR7GjSO/1iqPE8
pgkWzbh39AgxDq97ZwyAeSoBZr+RNed+cCaKYN909W+Uw59Q3pHkCGTNLYTteWEsp1YeMB5G7GFe
shM8RrLBzwRTiQkLgBQ5XtiT1fCaOuDsDXcbz6czEf7olsXaOD3zrmABOarZsRXZLHzgsihpJbvk
EiOP0lZbugs+N/t+sWB4/23LjUyQgRkonJxyHbi2u5voDPGxSYVZQuBf0jkQikT3/F/62IX/ZfDF
3XLqeqJ4oQHUGrdy0zWVHsJWGOQp57hTlRJeFZU+GO3uFglJ2GGCIoM1br75Mpg4D9OghpWueGUI
HJC7Jqy1QJitbv0Jijo8Fi+kVKKWFR5xGoSnFnYnc5uXBTCu02kH1w7cq4wNXKAPAWKkyy59bU6h
jkty7wHYzQDCGd3xNiBSwqgEAA0IgFAOVniSpuYoWDA7cE6AzOCNSlRaguHmfvgmYI6T1N6xanQO
XiCqlyWD6lphEpM3z6fOxvk3sfU42JfwjVDUjxuxQK2ExpID00OBdBKWvprq1288D7p66VRJFWph
BGvrmzsGzJ5uzDg5spDmJ6beMC833XaghMgsT81nexJGORwiwl7Sdq3nBgC49pSeQ76zzdkAXPG+
7KLCAJckMPBhhtXMtmV+CoI5VzKsxEpTZUgxLtv7st2xYfeTcnkAlWtvY0bHvc9hDJvtmbTkQKLY
mEFsiKCMjorveWb2tGY1JyMsvdXUokikwkS4/+TgNnMV3opdNlNK3yUmVVuo4fdzvtVTMwP2MQvr
x+uSz7io2u2qGgG49z/Nmxar7xhaDSxceSjFv0PQs1jl5NBcNGjf0G1dzQ5C0v+vobJWFTYG85i5
/Lnxw/JGxsROHIqeEvsFdlwGgbWnX/t8wbcj5MdQiEJht0XzFHe/2Vu3fVdASfPOVaHBwbxzufll
ml+pSg8yHw/3x1RZW7YSFG9ZmFCe7y2lnfcProDttpBOkjjNehAWl0Zv+i/Pp25q8kv9HhvJ9Qrn
8NgJXO15EtAVVleywD1vlJ1wiYSR2vX673Zd87AlDG0Uh3+amcVXVgD0T8hTMf/CPLCkI5t1VvFn
qxv8ynN21hOitQQi9aGSyhK6Ygoh7jVdOmnl4GShQ68zn78fLkTCrY+pdYmZS9MjI5oW+t8JSrqv
eC/0kFfTaBkfWoq6MKs0iIbGYiLtLhfTt1o3/SoWgD9ae8EypWFlfF//n2dGOa+p+00Ofa1g3wf8
TuAOwwhXtDXcptTzo+zeJ7K4ShX0M/S5WshrpC6WXGP9+1ha6tPt6PukeTLxDKn2FHaR9ezZHzU4
iYLjZyH/DKl6zygyskBWtrReJyJo26QoakzdX2iZG1UGIcgg1DeMQ3VBrIg8adH7E/Y1QZVDVOnA
57RidGs1Hoh7YTs/u8f2Asf48ZaNCvZCcBmZ/tULJ1igwc5ET/ctSnn7SvHaqf2Az2XPbPLsohvj
vKJOPx74ryRk7ZZ5lQAS8FnpafM59IXE+RppmV2Ox/Vesoe57bdfY7AeFlHWUvF0pFEk8KzILvSu
SnSoCtNoaVpgzV/UwFDlOh9nE6xvRrWY6dcChpdV5WNHJssFh6df7f6EbTHn/HIpakHicVFkn1ne
1h8SJOwgMbK8/cjNNf0SRwLt1O03JvEB0MtBGJTHpPPBpyGP75h3nPHOB78Exooe2EooY2uPbuZj
tJhJtlFNUUw8mkSS5EaXtisIt9VSY0YqlJ2xG7XGkZc8P3RoiZ3lSbuwKbGbZRNG29ofVPyqysnl
2aAqrRUpzPQFA8/c5JlnYy1Fh6BBB7uf5K1tvGFBV2Co86qhTqQj88Grb6+AaxOFf4+hCmKYwXib
9Yhy0//KZoE9gqFSIuPrwQlJryo8WkqqEs9RCWx1OuyT2sHDvAWUqQotcTpIA72XDqUcCio7MnF/
DKkUBVg1Zy0pWSvles3t7yGuVfOH60ggPi+OaQTbg1fU+d/WpruKZIXohwgilIi3R1Qe9mQX39Qg
jkEQZvCvLsuc4ei60hz760gTLGSzoehSqjQHBOAt+8LEI4F/84NiPWe16nVs2vKFf3tj15DS5LHi
0g30NW/WNqowo9T3UdE75XjgrfClzrxX4V5nIZ5WOT6x37ozVEtFrhtCnPitygEyktOyOJo7nGHK
bag3qDC1wpPnMIamxqral3Dv4FJfgqFtHwDYuuXCCR2MxWqYyAnsbnk3+hjE42NHAFIzqCtPXhoQ
jA0W2J5iAQ/v52c7nIxpSD2G0tOFmeRXd4m9W5fUzDMQ/uO+o9FoVTCQEMY5MmxZmXv6CVjW9D+e
jJUb+Yjj/jjvhSPlOv8w/tQwNjErNKV6xO705wfLSCX4v0X1ucsPOaw4gIFSfSWqYE+IOqJ8hghM
bdqwmWxI2xlreCrIkMJIHSvrxoOJVSY8Bx2kbhOZXZ43dPf1vOfGK46732qUPy5h5A1DZypVXZe/
6gyHh7ZOcPUw3BGXVV6jVGfSFDDsSx28Zti1p28gJvQOhpehWDNT5HrTbhM4PjEKi8PDK5UGo8tz
avlL8dVTuXgvrqO1FEwt0lFcqajmQWLDe3IZVjik4CwgIox+wMbNtN+f/cE0R44VQboO03ePgyGR
mX/mvC7k0fB8O/HNw7OvAcZTeFUAEI3+G/uyTQ386woHcUJ4o0eL6gRkk3WHhhXzVXwKR9DLhn3S
Gvia5RSqWkkIlskB5k8BvMEOX0UthbqbzGJsK2MTXuro5LjNrn8b8GSiAsgNMeOUp9SOqPR6VvAe
xU1ycYiZmaglbCfVptpRVHBYLRP6RWAhIUEFPNIazpu5xxLH6MbTRy68ArtqM7y/aPgKqtphatTf
x3r4jl/43eADdh0AHqdwnzlZZm2UxZh57nJxJGMS/QhFdLrGKGRc+AxZAHGFxgjkMJjufuAGVuHu
h5ES3CkwJ6ps4Hez+O1wb4lonBx0LG4nF5Pr1bIMj6IWZZbmG0emZYQetvKg8T4/oPqSMRHR5iPH
w1Zrl75Y1zx0RHLrG6IJs7svOUbxJpJw7v7f7vgc/4TAUxsX9Qo5rz11lEoMq0KifhozdONoz9kj
XSHA3ztz3IBjZsabXn+bh++0xZc5Lh01vKArjxYlScjVm+f/MLizJ6T1aLtDznvpZXKFSBpi6nkw
cecRcf38JjhvjroHjkwlUYcjdmEs3omUOvu6UIWkSb2jgFcpPfMhN3XCmmHVucMGD6XDcxETeDzn
CUTuKcmd6tsTVgvFhQufWpWFeVVzn9siJ+578Sy1wK1K7u1puOa3k1jzTHOqiK98z+QAmI1rsHjU
+37DoZQd03Gcu1g0CGzjYlQqIwGwj5TOWAbdoHhl3MEM6+rZl9+ot1dctv67O8NuRlD39V0m/6vk
dXyVSX9SWznv2OotzwfYi4Y+KZ/FV7QNq7ttbG+DraAbHVvI0cdTq2fQTXEHwCu9+mvojxRn9oM5
ngnWgpjwsMu0pXbEgVu3+UlZG7szKBpaX2J7hyqx7yEsPPcPrVfXtsC5irJJzkfZTMvoqVeRNsKa
YMEoKz/+rcEfnRmmxp3ThKjWd5aUdk3oUs8GuVyYL5yu+DP2VCXXu4IGwA3YZJsqnEeL9UgFDS6F
zPIX21xauO6cOxmYU7apuT10G2LHEBLv8q/6gxc5RrOYT7VJNPcgg5/XiUpGSt6IYTItZLCsaIv2
BUnpbwidKjcq1qp3Jyc1JSoMGVwr1Ef0dETGR3n0EKVhxtqfuwssFAOX6TKJTXelqzHNzt5mZoWr
xbxVJGA8Wu8Tlh0UIfJNflIe//M2irQaV1O/i4Su+bpwkTL5dXPOfxxlVCMs+ZHTJnB6JjwCn4FW
VbtkProSIuM4cDwdmc0FcYj9LoxYdQCzMAfNQ2OQxHuUSrWRk+qYFJfAyDSH8IkYkl0SwMWSUVfk
x6I73HQHnwHSHOTyixyQvmYbLTkUJY9TSBQ3S/JjfifDbsmKsuWnN9G/mYafQZnCgRHJ9/qqlE2g
5hivW1Jf13OpWjZvXoEhtYBrHsiH2nXr04ZofGMN9yFSUhr0SlaPfHYk+ZXCNJCAcTHJfcKJ4Id8
fgntRFTTuOLwPTtvFZT3IYF3S4FNvbwgyjesaBeHfUM9RaPngk0TPM9YB8PjA7iiEzzEymf/aDxq
ljcyCWM9GEVMz2aoQ0yykOF/QOMLztdN7xM11X69GNl7/eHw6kkFV7qdlwPMpeVr5JEojQujmah0
faHQpZqrsriE69jAsfpwpsyFAAx5R9PvChC03vPLQ0Tv8FA6+3WEHjknr4kIq1LbdT1YaYtspeKj
qoH2ybnrnKy1D078o65BSvTlur3vsbB5L5/VfQVc2NmJjir9LKFvax6tQM5waWeiM1ZYuoJSrFUd
Z9dhDYwFjSziwe82Z7NHcHAMoXEjHnVqLD3O+KcvIVr2pY6TZfsO7eDz4v6o/xBCoM2eLL9WSa8M
IFNfTgrdkFSrs2O9nl8V4em/cI/5962ngMxQu7la3mRv7M7EYakoze3QgQuyqKZhmHaHXCFV4auc
qUnxZChXrwxiFE5iWA5IPR6bpVoYAG4BgNFDL5pqYrENqpiE2PAS/EqQ1b1IxwP/Y/gVFl1Ju7jW
wDeG+I3qwSEhDRtUl3GcLbQkDLa/z/kSVgBYlKpLa1GJevlXDKyz8RYWyPC6nTt+ZqKTyh5ZdbvQ
QxfAtMP8jqD9vrf3fLoIbpoP7Pd9HK9vXmlRQPpygsR0KM+KLtPL76MK7H80oohXxcsOsUFUgLlC
IW00GTU8XXiBH4hxMzrnHqXHhQ1NPHsZDn4IV1Hic8ARIog6NrEABu254Y9cPYruTHsFHfM+LhRo
3EAARNuJibbthF3mS/HT8kVb7/6ugzR8XtH8ytruTB+IAoqpR5accJTHnXJjWw0eBukW1hQkHdJv
KrfsUihAXQwCBRzKuIQYYWc3HixD4953zaoL6b4+/PwZw6UFn/9jImsK1e4E/JpAZs2039gVvonT
iQPVjH2m08sdn4rvbP4kFKpXGtr6irmtYpHHdNm0bqLCOy5EaaC55G/BOBsrAsKBDvcgwEf3Jyt5
za3L42dlBpCRr6ill+N7mY4cmoAGsAmDhlAeQqfDYECfH6V3ZKhbcp9UFQy2RAx3/JHc8yjEr9ts
1RDzF8Wpw1jEAr0h4HbjnEyzd6UkIfDP0wH/+CNoxqzwZnrzfkmCFV5zTbwxld+GS3kSDWEZE3zN
g2YdJmvaAT8PDXpK6JpeVSjQcPkciFBS+8na4it8yIk0JK/ha8MCigaRJu3GeYCMp0D69OZArrHW
4tQk6Oh+QE6VTEUBB1/7wPJRlOc+stEeif89bxHbCoYOhhbhDSrgEArRpGhxTN/nhNlTqXFbmn9T
wsXF/FpXBzirU/1Is9pJdHz4iCI+5YoW+IfAHgBKu1haVhc/f2zx8OO2aTPYgFQgxaL2abpqnv8g
/HspS458tD7TafanqtUOJskuUjH01d7hDzoA6Ya6Vo7LoC8OfuFmYDF3CgeQ0u8iA5tNMYHnvRkx
xgfJVJjsRlD/mAgo9kGmjaI5giKjsm/zajjuhxXRSQCzmjHjPlrlWjn/Ks5Y+TfYnRNb3WbgETe0
FpliEHgSGtoOD8zFlNhkVBHxwOIC2LMP+k18TdmXhtBQcOXiswpuE7ZVPGRRmhcuyXsPSF+o6njQ
unM7Zzf0hHt3tBEWegi6XffWpbnBCm6OHimswEL7Pb7HCfmiZ7F8A9bMsC0OLTQYX2qNBq2fafRR
GBIFfIdDKRjsYQ7wCchzfMh8cPgfK9Z8mV2Ilqz7Y8ibCPO+NhU6TGmRMpCnHN8rgj1E/UUs521a
bxkbq5fknLP75+Hf5JEBroRqIwpaNDwQG6HEYSigVH5nCDV4OXUWvw/HJuePuw5DGFY7VNdRGvil
esTxlwyxW/TGF32APyjRTwFBCgTMX2pMCGpQjpP88LgmKEAgM5PE8IQPMWeK0QoqFvpWZ/mNs7ya
1Ki9uyBrNXfh+YyEf77id5/nJfJX4k6a+ScBK51fvQPZeXe7jjnk/E2F+S9yseCS+68N2wk8b2SS
pwVyDWAed4iuy7riArPTD4gEJdrN7At2IgXBRHxTq+0t4lQLLu6T/7Vy0Cs1mRSGqARAey82BME1
CLFAzLFP3Ighg8sMxbvBP87nLvpILO8kB5LTaMJNuYOGeMc2dI4/mvtff4p/ksPZuDl1jlMKa1lR
VnUHil6VkNhgsyvpnj+YMmmghOadT2noxh2AfoXwR89qr+m14M2D2y1ZmEoY0PzcLdmMB6Br+A7n
pyonoNA2Pvwy+kuHVJpWmhu7LNJLmTbPxBJcBdiYUAmk9qDarho0lWIrLG4VX2XRrzloit5/AvUF
+F0PlCPGIzgujVN6lAhK15lHO7JDcptpsDnZ+k28j7il8EKF+9HuKXk/8lG8AGr6ozh9Y0kfH1Gi
foLs4OApcvK+rGE/BAEaCMyaD3xBBMRmV8Ta2t28ELYBZ9CyGTftvkF268QQC47igbI9nQWbXR3A
SX6kbRMhvh4OmopGiQRNevB1+ZUYi5Q2Yx7SSjccOVhf8hF6VsRjqsKvMc5ycj8ljDQSx3nQlVGT
X7dIUCAhOm8SL/hl4jHZUyfo8neBO20CjvDZFal2G5IlVrhuHq8RmwtIPLb+aeskR9MoGhKzH+G3
DuXU9IRmCSQXAz+TVZWDTnuRLB3A+OlX74ch79/wxuVSMkJN5k7tAs0pyXdL4H09hZNcaipZeH7K
+/DsM12cQlCHt9czXh0mTKO6/wL0wTSNXVm+NLuIWgNY3ZJYfy5LqppJ1cKMhDt9ow2cYZJLxt/E
v33IW+Imb0Vz4YhcvbbsnVf51vq8OJlv81zfGgVeQgeJtEw2fetNFqMWQMpRQt3FBpD6s4OaBCXS
aaBD/b2GWfL4oX4qyP+LnfwEE66TKZ1YchzJjayQIkY1f4TqeElCVS+5l0lzAlNYGzcyK2Iu0rjh
16dXieERbQKbagLnJsxDNeZkYbCwXAFtbD1NJVqsn/qu0FU0uDE9m5dHF80PRQdSAqBMRfUCP39H
BgfCPb6pBQMyz4QOUxB8ad7WYYpFlp1ipAgbRlNYoF7Jh8M9/yaHF+zvNR1todeG+HjUYn/0h4zz
gQcN/Wo2n5ukTlqrogwEBU0kRO09DCf2O/soDpaGWwCcXrAUIr57EVaNa+0S9eZzXSUxfnX3aANT
AUEejAGCmTDVzR2TADn8fsWjJgqhokihjAGqIpax4i3PWIYRSr70BqOmLoNHs/uIdeJd8VOWQHgK
aiiSPUyc6iAml1lEukoXUHCfvYA8GcUyUYwShIIAQrUlMQ6HBnPb2C+cRx69JAnmHVViXBbgu3Dv
ov8aSZSQSR7aY+833OLoMvdbJnt8f1VQBOgpaSdI6WNNTTZPS3z4jlRNEFA0x8/1sKLXBN2ZMHhZ
STrchcCtcdeM5MQK+an8NxeIVyxf8yph2E9Y+y8qNF2S47uiy1hj+D64m4ru5Uz/bQn7QMqaDGyV
jvLbVjc38ZsOSDAqejY5BDAgTCnOBkozsZ5QE7fcXGYmbkXrkKNp12tJjo87gGe8h0hFNt8Isn12
7D9ihJ20EqPCnOcZ3VZwEfkJ4BLOh6yjIGCAKrqir2BWJc5QciqiSVngvOH9ma2ZVJnK4W1YBjG6
HPvM4Hz46TQUOrfhsgMBsiRmFlzqdRpcO8w+RzzWXinsChx6rGHZgheeaZTTBhqdYZ/p1XKkeMo/
5bLTEjmjfukM3YQE2bVSPOOTh5qHYbKz6JRETWZYRTC7AOTbL8XfP5t+ql+j7IFbd/kowoGXIwwx
eZZy4mjEhw5OhFhJKRadeyyd8jZunb+CGanmKVEXYURPWgVx58EbaP+oknD562r4BprHPw31Mf3F
+xz2TNE6aJjjhbpyzixJsmyHR//6B1xCposMVlgIRp+1B0VtVT6WNRhnOm8LM3iUerI5n0DOoAyx
6utShH7V7MsIFW6SGrb2JQv4LtkAsemof9I11dVxMsvXJHotDDh1V+XBb4LWJVSZhR6RUDe7ZCNU
8mGcr+tawp1PZ29Pmo4GeW4cOPT82t/ToxFsb6hV8ZbGTGlxHB4God4Gz3yBgNslnA96j494PtxY
VCKeo0+0FSx5SG5TKRRUuP47zkAobju1bzkmXNlMrASxI5ENkTbYqDEKw3ObJsO8e3/mEHMN135J
AwLQ9ML6acB/pGwOrvC7YPwt9Z9sfndDO9fV5e28HysLdSyDy1zVDdwKmCmW0s1uprfdcikwFq2p
OwxCAD4XKCMyZT9rGxKyjJmQWfZPQONbcnaZL8iFCRO3R0W2SmMuHzHq3sLecyVBlfNicFcitTHS
Re7Al5o95l5ugSlUDizM2qEkQx+1cYDisP1yOhBMAq2HJlSvTA4czTCRaafBIWgLdPULIs/wDzFB
UV3EG4rvNWWJncD9Ka3meIc/DHXBDPKS9RIU8EaJKuZqFMdctLXSfcAprG7cdNWgviTvX1GhkKvN
L6fVTDOnLgRUWiWWAKfho5fCKoP+goHonurg4LRfTbQ2bDg+iBxpymMV5wHgC0UBiC//KINdtFpH
h5QsGW5MYm3jSOek7zi3YR8noNYgLE/QkkhwgxHX4g8PBbhCFUklX8xCqm96ji+IyhSZ9W/kDSMR
59HJhn9MNQKZ8u9D14NudqbhYMyqK6yMMLj0JUPh7RWv5evWY6AUEe+AACFUhkEGp6xW6fPQJzl/
JhxW1gycXb6eYwaNJxiIaia/D9dWeVI2gmzzEfIW2ioVAdmM7NanmSaPJBmQodkDY/iIjUEa6ke1
9KFDRDxCyXqGDMsfgOk6tB0lmzSDQQYPLGAFrf0f+BmiHerYe5lSyhxMC1LSZMbOzjijD7om9ByZ
4IJIZnCdmu2L1xvflq584QyI3qm2yXh8/FGA1QowG5VuUBHz297u/ge6I2sA2iwFF5nlpKkHKwyh
jNGNKyDYI4B5GPzfH69mn4oKm4xp65i/mGnKNCdDFOHATGGEFcq1tYmD4eIohj3ms2KXcBDKpzxZ
MGMR8OY3Gp9QLq9W7HtJF5FNUc7DUNQOWbgccS5D/HOknZGMFphL2I4PKnvfDbTXVb4TiluxVNTm
ilb+mt7hVQLqcLp+tAt0vDPROVlgNs4ZBiUBvlWwmxcJjv5lqP877h+VDEoBZlrKNNlCoSaVdj3U
n+skCsJj1Kh6h45p13+06prWmayBEeMmV4ecfkMHbQ324QCWvTiiMhQ3QpjggXtc5KbaD1QN/a7B
s/RMJ3y1U22/G47sEkvhz0WFw19JE2UgPh1Ue3JjtVym30LSufeTu7uFFO2ZQ9cvIFJTV+qt5Lpg
EkBemK6w+zMLaG87ghUkKTQwnpYig0JkL1Rxil1SEAFfev7xuRd7gyl8/wdM0+a2pubCWpgvrk+4
5NJ3OhNw8NkuOXvbfwHH5Rj/wf24ITY1L4XfxrMjGolKlGRw0obSuZMeDBmgYC9ysab91G2upps2
tZtDCFyEkOh/huGd4PSN9+SQuIwjHoweDvpRsEqsLsF/ozHVyiHTgeCcxWwMqumySE8ds26/dRZ0
SFo4SYO3bV7XW4707TO5aRUfREWPU3fYrew4iNcjCqJv0YdKxYVYgdqiVwmu0BF96+r+naGSc3H/
LxY9mvlwYhy90/f373FZ1ybFo6W9cwAwDTy3dZivIIDpgJCC++fN9BYyEjVHBl1GAtsOJqfiapAQ
znLsTT5a+7hNNsASIBDsjy4X+9z2QwPeCh+tCndBf3d1pDshfDtP1/A3GVayl2PfoXoyLS8EPtPj
QRet8O7CvfzZ6oMB0soOVeQhdBvB1dbtE7hgMAa1RTbHTAO4lLhSLmvIbkRKkF2Lc+6pTnQivzBH
0nBGZ3t7r/b5nn41azxGvePBud/bgEKdU6Rolg2xHnd7l0Q736Mb8zXB2wHTcR2P1l+WDNSSrwCB
x+4q/d367ZMdRSjqNhS5sL9HwI1H2Uly0q6/QSYWJKLGQgMsgenWN3GWkjIwQkDeTt6V6INVkDyj
zxUPD3M9ai8Fqhg9qjhy2Y4fI2H/AHQkRQuMEaeA47SotMAo5oDB8JwQN0NuUyJ8i4F2qL0FIFrG
qbTmtMnbgfFwqm4Bo07xbFGw4ohkqTAnZ0DNKdF7Ehl+YFAerdIx5OYKHS2lJeZqN7KjF7C7Z15L
7PeIBhvmYl+JLOTqvRHGP6vcvSITeQSZlBeRE06wnvuRVeKQdiqBU6MxW9yY8zMa8/zpCxSl0PFo
hrJAPxkWJgBtUf0yqEgcuaZfg8787cOpiPqFTDPE4hRp92YkXWyb/o+jyrOsURcmJzIJZPay+JUL
BVoVbog2v5myIbWmDLXQfnN51Mfzwn00tMMm/htrUEB9zj/Jv3R/wUgzlFxo9NPtACz+al70lL0M
rNvGGoV3v+kcTmmekGkZGTE56WSUUJe2pDPJHBiAyzz9qN50CA6EXvn9eOHcCZvNf9NVO6bvzMXa
EZbPGZwtGIWW7In2r1LsEDOe+Gyg5RuMvTtrUV6Yj1bZ8e7riPevkFgTjGLi7tEkihSRs1SG21T1
HRT8/XabmaaBnxUxWWYYhDQzM/0Md6q3z9IzovZXRVp0sZFGWTpXq5D9VXo0PvbhZSlh5PMLoDtT
q5Yxj2ZKYxgSjBmy/6PsTz63CsFZs/+dedEpD7OL86eZ8nBAI/iLfc9LGdaXCm0nPBlsWRjYSqmk
Nvot5kURfOzOr9cvm2eoa2IxOU0JK3gU4Zax8VRSyxHpfTseI3v0xWWLTgA4hhsVV/VHOzTNsI/r
xTMwrweCZf9Wm24Bcknc0ZMbFWFWj3wpfrNGsXXs7V28Z1g1cmDWoTdMmSN7LnetSMgF5VvCZ0Fm
LqZUD9HkK4qhj46ygmZ13Vpn8Y0gZaZxjMchKSFjt8CSBuA+OGf0i82zlFagcF133Vj/jlxnFSeE
18IJO1u7l7/Z3rCWputbAg1YHIxiZRXtLV18QdMwpM+mf4N1p4Yw/d4lceXrntrqsFPy3I9biMMb
Haoy5xfPsv5ld45gLj+FjKcCm6yMWm1bG+Bg6Jf7NzNrl28WFXG32n+RRVAvBdzRwDP8WR5KsivS
jKncknMv7a81NesMWcvYubX5pblFqblINuNkH36+mu8E1KfgFti+niRL+hUfQgrqg3WCPf31fGZ2
Ox3isyJqshQAYDm52hc3214MMam9AcWIBCUCepQcNPCBaIhmUE9RR2oCV4gMZ13RVl3rSazJLbXv
U4F9D2mh9znrJBOR7WRdnVGk7nFhkRtCPNqUSYM8K2LHaFd99dMFf4qb7zXY4HBL2IdrPXJH36QA
96Fwo/ZX4p0g8eSnAjm0dTiJmzKc7EFDHtSysXeZ7m8kgApkc8+sUPEXByCyxzyom2JfAD5ApRCD
NCZFrMjUC0ZYlc6jGR7PgmsUFhh09YgYNvwts6d5mg82/3D8k0pJ+/hnE4uwObz3qLXIlGLpRicX
tmijoi+GfliiufbwwMTu1zbBi0pVmk5LSuePLKsnvb0nG6RK3yJ7v+nGjp94gSAT9Z37HZwRo/Hi
TiS2PBHsLICkkepBj+ZHmp13A3ap5Ns3G2zffySskQKE32OGpMQQkl68mhtOw1k4hoxZL/MxBDXo
ldfpKKQrXrDRt8mBTgBgYwt4F8LJXRulpA1ihquPvNj8rbf++0eNMEfSIwr3hHN7Jj/0HCX/MoKk
8W1SBe8bYAQLos0Uu0InTCZeLASHJFyJwQifY/v8Lx5vo1NHZr1zLipmPdFpSGHzMH9cQ5kJAhMC
Sq3z0lqNCl9A9tLOvLbpFAnbUPgmyQWDQZpraeONcldZS4rdNBhRTPBWU/+ZIHMa1naCt13/smKN
XGT+zwNZ2ysNnHxaTFyHizh58afjEtOTaVsyP9JloaD3O0fI1AiFykF77hx5DCdJj0bB3CYS54lR
3ilBu0ZHaWcJATYIHb4gn+5dy41yO7TevXIeOhu+bFmsSr4Xx2Ck8sVhKPnxEKbcS3ynXzqXija1
iFc9Br+zyIJ9buNdcBpBM0Qkrx/12+rFqXhKcuHQZQs84iQewA/2cVjkDwymK14Hmm47RmI/dXFa
hG5+urj6vFJ6M24qqgWw/eJkeyI2Qreg5u7cIsRNa4jzAj8QqRNEUiR7W69bMxF10UELH/t9PLUF
JetxTNCMiIVVaEKyKhpf+H2/YvmJGm6D9m2+CJ2uQU92vP2AK11opj4ua02yUK+kpWdl3UOJdKND
t3tRMWgb83InUk3AChjwZjjTHZQT0jjFQdp8EQt0fGYKByZ2/R+Z0wEPoh4Ht92iPXKUuzJGRB6a
K2EHuYtNta3di3mM+WbubTuFabloY94nnkADrj/776k1Xg3k4T39Qdj4zxKERHr3KW3tsUzbFQ2H
Wad2XgyOSg1DywCDW9NnAlzdyxPgWJKmSr57oaSBt6pv7EtfsEn6JKsoFwJNWAzw8tqaPzrjEcwa
4HjGNdZYfptl4rTxi9myBkrRz1rb/8XBl2t5TUj7QRnQgm1QPRz77lS9Ht7a6x6zQX5IQGTXBqM6
GPJjVGFpHgvdFBzfLJODzgkinEteBD6xLEMPvPUC2SWYCnNGmMCAX9Yixw4KS1OI0bQ12JzlG4EE
nJtBGP5EI+v4R+Lx9HHylAvfBdlyQPuxfgZnLd324Tl6My94SYy1Rk+p+IgBsXoS+8PGaAFtnXtp
gn65Rt/6AjMluNHDniNu4WuPnO8MtEIWQTHyw6x3igcr9SG26jjJFfgNBQdeTnQoLeXJH6yey/Ds
toQJV1UI+Z6Kij/tn1jJycPU5WftxlnzeKEmKLO83IdsJN4ymAotdpLfPjQFJ447kUvOtLDRNa18
u3D0lkyHiVlXVFaUfUlAu2oTdxItf20O3mNKbNZV08IzTJWxZlW2/aBreSh0OTPDQwmh6wewxgEb
BNqInicY+M4juXX+LYQ+EDfEf3jeUg+qHphiX8UlMjsYu0ZGXTAPvPTa6eoFbsbve3c3CHvUzxa6
nwUq8mg6m8Dg7wLgI+29lARvLW5APBfTXyUPR8ZXBfb8cx1N+OUcUviqX5eGSHuh3tt6+fOR+27o
dEONnxGUiEj1GyBQSibtaEEYlHClazERMg83zHPAqO+dZd/FipNtNuAPnNRfG9aKH7ZaOkEzhT4Z
o3bxWZQYmSsA74Qg5iewiFFgQsWa+rzld3Pfx6MmXdKjWCY3RHLdfykVQjplINXAQG581DEFA9cC
dZCnHS/nzJAAvyXiqSWbQ74B+rV8XaNtsYddzy9fL+bi6k0oABGmDyupNtzGiCNd43G5YZE3I5oL
PepjXrjAe62eJwoJmS+UigvtqzUJeLuHvkA79DaBapOrFBXhEHs2saYRJk/eB9cuFzrTVqHc5KUF
CneuZbT9Sk6f4Tzc23Q8j7jy3yvi8YUw4onICP/Do65SeQfBhvT5CjaDQH2lgpb6HMMr0u/TdvQP
8y3gJR558XtxQpdvyGMlM/7T1UPRtTKVC1Ti6K6mZVUWNd7MRrUmQP5F2dLsfH15ggYsgpvVeUKP
heRzBRzJFXRdJCrhK66rPZFCDgvdDM9BPLtEMtR6k9d79hkUrv2L9C1abQA6ku6iNWvORCfqs73Q
irqkNFybdO892FlMg6usJYJmy9P1Oih4lWp9BZB8VYoA7Y6JFeRZutwE22kl6cY00Rfsn642Wbnj
8N8oXPllfxBId/6mWcNjP7oefhhJfGn03cu+Q/a/HnyvUwNbnRvecjVl0M/pnHDLKP+z4OugEfDY
4YrCYAI5JYGEl4yb/O0ebxbbqKgyOcswjqpo+aHUuoisfGSKwLEu7K3Cc9pj25O5jyJPib3OLqXI
cifOKZMOcnKuNKSJ2e3bHT8P9KIRdvkbzxAkhgp6c14oFF+FvOzGDUAlKQYgjmGru5aYKdDwQS+d
WhYC+OuPckkPvlGMkHnQSekDVPoo5pXL+v4uS1vwKNtmzDQxiqCDiyWOD+K5A+xlhXQBgtifcDkC
q+uNjJdwBDxT/Uw8kOAuC3x8JP+YU8cjNTMO6BPI9Mi6cYEXHBff+9ZJpwcNSWJTYY+RhHqR9xCG
CdPHOI1cGu6olew5CQJEShNEYZs8qhUD/5cNLFiGPm3LYpIiVYvpQRl3Y0ddGyrolV2Nsl58qJZv
3tekZaVe2c8lSrzQV3B2zHCgiSl9cAuW3HG7TAobPxOEfd/OaoRGm0GseYNohF6aTkAVeHlohQsL
QmCF9KhaEAcgyK2VyxDavELCGHImP05BDum6+HKIbgNRdu0xNhJEPUrgBGdrthVQvWlTc74jkRRK
q7ta2cdA2RPNGtOmhWRyGym4hGBFtJoMLhYEIj+INHHwxC0JXxscSITfmfUUH60nqzGpFKV9z4oE
Uh68KBfwcfMT/jF07eSKrRIcb8JXAbK0xvuCDXfUbk58b9x/DnHQd1e9kp48aThs6bBPRi0wBnUU
73IgOzWRvJcZHG4X9pU9Ci2GUEluEWKu1jzVc7IpdymdmUjUDIac5n3d6EYwogLtDFJi/PCEYtrL
TyRMJs9IkCKndF7i95nru5I0iW0sYPYM17eMCo2RGIs8cdkn80uJAfVYVr8822u/PG+OwubEpC6G
sM5bAZFnYEiMaj6ktgnPNQaerM+A/xK1M7VN07ply0T66/Rvf3ntQSm6XPbP3tDYUS7gKXH9FVbp
HIDXdFYMCOA3Gmz22KpHf3iRrwN2KDFyR0jFipDa1ludI+Lj8AvSHxTvyZa9RdvwHCspr5V5WH1z
9+QVLAAtqp6t3BJFbfFAdaMsX3c8BE5Y6UXBxbGCocVE7proCkcc/L0w/5UeLowvrhceKPl23IYR
jjOJP2RyXRy/6VUbWZFAhL88znNwCDg9qy7gTDbssGdaaNwNgmKIqaazS5iD0dIDa4EeVCYjKXhO
bFirlPES3LUVNjQ1X2Kw/YRKJhxs8QMTKPYWeUWkc/R8bWojK0mb85nrzShLwN2gAjzUBVsPwQnr
USRfm2xMfKmenamtlBsreXorjKmu5RsEIuBcjOYd5QTnRsEHsZNpAPU3oZpsZQ8c8fxXa7jHRCQ0
7wZhuS9iE+ojyDT9lTGSsOCo1IWLkT52HpXmt9gwLW2G5XHvoga06yuXW1C58xnuT3DMV6oESHk4
capJ0yWfizLrbzIQsesdlNYmoB+CKIW5Y/n/HcGOcZU4WvzzUowwaUEBymz72Fv1oTgdPG5RgS0E
FKUNATxmMdaibdMRtpF6W/KbfDqVxR0gmxxFHI0Edd3BSOMk/Fp51SD3SOh5upHqCM4XrfKPNcd1
Tvl6jpbYcmX+Z/6HkKfUSWSrr6l7v2RxtW62T+U2SpgtvpVjpqwxsSMrOz5I+UGXsxpTk/F1M+x5
XwR2ffZhUwxUFimwEQX5W86wB/n1pVdwxqgwgFj7vF5/axlUReUm/ejyagCkFtZVmfZfi9bDaPSw
GDZA47uUnaV7/bDcHjc3+8U0Ejd5OhRh9iSKk6fWRTNBP/disREkD5zqzH5jmS0wJsyT0X8xvqI6
jKjW1W+7Fg5BNtFL0aI9a2rnIx7BQbwCoZKK1mpzEOK501uQPu76Zg+x4PipRgswVgV8L9RbleMg
8py6yybk2Slj5T1OaLB+7teNWX3w/dYcYHzFnx/SPaGW8eE1cIyzneSMx/Ug3k3OhkihQ9KAwZfP
I4OILhV66PAz0bgKXub34SdAvXlH0Rv/f+BljbRVhMgunznKJNyf6FoAdTJXUrHqzIK2kn4AYsxv
Z1kJSGtAsSUDwZ27/jV2oMCuhkUjA5pvrMT39TbbAl3S0vNCiXTza747YYxGxj7gmVCtCaoqcODk
xh/E+cFuXf8sfhfWrQiqXanHQzAJAfI+qLIE0E/+BVe2dP+LOk/g2Yrtq+WjXwqO3Y9ZNanhWCgd
MPaAg5wgpyieW/5wVEg7T0rGYZYjJddCxLTbY1jaQwCnsdIH7ZRmN6xc3NXKOeehBht8aE36U03W
JIOF6f7xjmcCaMt2xjjKMXSVO+RAw2r6kbUznsfWXk0MbcVPfv4cYNjRhUP0B/AFGS8jJ81pQEF9
uh2picDbFG+7jwCn/oPQcLaR7Dyaioe6+uGCgBsdtOf7QTy4t+AZ6coUA2MKWaH4erPiEuAjb489
AFuRjSV8B3SIxbRo3ZBwDdoFZMGo8Ua5tTvyxnpQdvcJ9Q1SF2oRUBQXN3DyPSw/O9/f9q3WHrnd
rLWDpVGeEIWmJOGQZLZy0MX9B0sLtqz9F2NN0CETTt54ZoG23w+kfqKcz5JdvyOHS+rogrtWN95t
l4CY5JyYg16DOYMLqNSI87oo+h3QRj6/wEVNMAU86UBz/+da7lARtsYTPZKmBqdnOLhyHAkftkPi
A3CoyPdkCssE3XoL6vg/tKRBIajTvjlj5KQIkhL4CGWpt5Q4m/2MJg+rhVHWhnt0pDKkeDQtlOKp
k1Yh5bsetLt4U9c18gDnbBGsMRo7raD9A12Zk68Skqxi3rFH1jZ7Gce3pvSlLwuoAMtu778FSiHl
0p3xbVO4mtDnxHlwc1HVEolkqge0ASwjcQL5SIRpOgAfp5s7DLeF7eJAGbDC2PVHth3kR4GQb4kc
h2xuNCe/Ko2S1SsIZU5EzgVswwIux5NYvSkimRdrJtFE533ekbP0QBKRA6M8ly7GnwPLplGXCjta
cqJI3tbAhb+BrSWwI1lvWUlRXq9tjY3nM8LGlspboEA3D6IMV/bRqyqTh0AC6gjCA+UQLKAWTRtC
T2eVfL4x6br3lz2TuEGlwUQL6hi/PL0YCKyqdejeOxmiNaZgYN46evoWX3tMjSW4r28HPMjmmyEU
30fJtUHuNIii8O1rPwL4aveUI7V52jHf0prOINNhOqIG25Uxh+yj7UM/7zfc6aJPUr6NzBhpDlfG
eJ66wb5qLb1yvpq7ld7EXCcv01iiNY5X1ItdasblZCUdP0mEkCtrqbrTSsDFbZQWqTSQttkZfLC8
borJIiCH6OFgfg1HG0pJSUR7oZfWV+rv1DHDIdY570FxunFR89ukRmRJW2KOS9J/ZyJmt+nyFP2k
DgHoZQPcm+a/885z9KB9lr9LfH69LE0DKRxu1cpNaQigjvMPXjQxJSpJmQh2aR+2vanojNaRM/ST
NIvedMSgvMMxVW8dCp1iKAnlT1v51AW4X/MwAP1n9n4FLBg5A9yduzPwy0KPs0kiNzoeuncmlKB+
gk/0mYphglZfRUpJo4MQtfT1PX8D6XUiF+W7TZvNMp7XRmQ0PoFjbvlQ3IGuLHa82voVV+jCGlI5
HBcdUYU/ypuPg2X0IuBXXmEGuSr1NffvOvv9AO5XsKY09llmrkcscLxzEWegkVE85MdauJOeCVzy
hr/Z72J44N4KJITta8YaDV/krf5j6PaZNkpAO+xittWh8QVKpcoU5zscSRsVmDbxlz5zwT+P+gZX
07oyZnVQjZ24+srbbIqU1xCmkKFrPvRxHDV3LHEnxGp8ad/NveUuopNWIwsOMhDwjmrWNx75dWpm
59tsvSsgb7ds1CX21py1V0CAPRMNlR8J9J3ZwfhY5/AZSw9OuXkXyCcbC950AQsYfUsz6H6ok++s
hmu+Vj/IiEpMlMpu/U3daR5/dGalC1dQr3BJnWe8xgxGGRhk0sguriyqCkWRk9mBgVTJEoDwZnDm
gPNO12bj1J/SQt+RHd49LJvH4UlL2+VToUUyBGz8uiYFaWW0E+Z8j1GPJ6plvYu5kNyD7nNAluJn
Z0KwoVo+ROrP1hX+2bQJ0sPzJCjlcYrkYz1oDLQoa1WiSLX7NvifEu99Rf/PjpayDyEWasaXnnUl
GHgXot5GRR7Qr9lKI+eVWZUdMk83NGhyjiQgM4CjFRMDXWOJ7eFbqb2fm2HulM4mCl76BWTyRnKP
nVdSsy2XtW37pCO4T0iV+Q2W45RAobM6VYrK8PPKufp8k8PwEFmaYElcdnxwqjnc/u6QsbuVsKm5
11vuznSBxV/hQqTPKUpKgKE5M9nai2bAp0D3+PlImk70VgsyI6xRxiHe1k+XcZDgYz7R12yEY7UK
EO68tLsMSAb2YBrna58ysX4ABPaBEwVANmq9+N2sBQ4KD4+oeTPxQrTBgtl3oZfGJlTpyI1aQe2c
dfwwgl5RLSXsMfq93FSWOqm66YlmqR/FbQKtlWnz6YEmsuoJobStd08s/niSDe3ubNmWGI2iasOf
tLPN5pdyfRKM6zN7el/wXKZ0DSsbjPXJVZsY2jEt2lzjzOMz/TqPe5WgYnC9jCpwCkfXslvp8NEk
LKnJMsVQWWkQxbHhECYRuhifLeEmsK7rclX5jddE6IRfIj2yFzs+gMufmaJREoEACFDxoYzwQ9bi
zlHLc5LW4trjWkBWrqU0Klc0CeRZJj2/PxS12DLcZz3BYOoHJgKXtxhUosjD6KF7AnQOTmQbRKz2
Z1s/BEjS3ZvmhiydVn1jYrlEbHXu6B1GNtZn1vqrkN0OhGvG/2Q1DaQu783Hz/DmdNamq4NNuxWT
kMMLdSlpZd6R2UyI37r/9LmUHBOh0A6FtoCuc5kZ3s1xouqy5zpbaPilAtePeIz8s0PP/Xuj0ZEO
lrRmhNo6Hyz2HOWVjruyAgF259V5CTcIjls1HlUmJZr2BfBn4NPoSu+jO+rjb+67gabhSaleUu2f
SWdxZ0YWnFPY8WAZddxVCAvOaajOCJtmhZLCRCIbdPkhdeY/6gqeWPgwCR/tLja35SHA5iUJ5L44
d8lMuyfspLUXB5svmjJZi5Seeb7YuFEu4Krg1gCpHQfOa/+3RZEJBfn228xwZKDavPuFA76Hsa3M
TDTLqf6EHNX8e4Enr6LbkxXc4FFBIRzoHU44eRHMxsi/ASmkqmkhsjU1HmJqJmeZv44WLBQf1GsX
H7aI7rTuNxqXZFibhJ17oZUHwhOU9wNN8tBf3CRi66TGMs0vaDVs3XxhcCJgUEnvh9dK4BLaVVAK
S0Jxqo8p5m0tNyqUPotpsYfRGc05rNZX6JtOROAiqwEL3Xo6Kwxe0dpm0ZZbXDWIok+tiPBmSw6o
Hjd59ewjdNJca5eMytjwNiUwJcmL4qRpqXx1IubssXaccw5X67EZ8pQ7xmO4+SWTaIkMF3qIeTKt
7abk7sJkVWJB7+tysVVj8LzRpih03rRWbd1G/hk5WeKiAeggjamGB7fUAWUufxYTGpxCb6UarYAM
mWEEzUlgSwbgrIgdyUohshmOKofq0Aa+Swl+etnoBo+1OTZW3hI+S/lXqKYhUhdZXiZPGrwzIc3H
7A/6vJPSASeZYx6a+q6DeNCqbmjDxqSrvFWFZ8523hbZbnpwnOOoB+DTpnIb6G1VDaF5So9DxoJZ
E2EZdVPHiZ/QJVfqlEXv0mY776s7egbIYh4CJ00Sz+0SEZxx+/ZuT3EKWt/xWUSbJPsAmW9tuyvc
6xQvwZ/6E2nzE7WlP3oT6OHxazI0dOzU9Je5rtJDrAyMBrxhnk0KLBCaH1nKxLJxX6ayaEEgBaxt
qlVIE4hJIXHe6PuTeXfAGq/UKns1P/nxPV7AQAdJTq15cRoPta3Uhr05l+mwHajxxYokPrkt5rA4
L1e7dXNZl0jMxwWhihDV3TyKnyV9r95K9xDHUyFsNPNUxfE5WF+0eqhhU+O2ZolkzHVg+on0NAoH
n8vF/J8GPchDiEo6OGO17gEo1Hr/5dmNlXyc2r4ai8fuPRt03yflqgyDFV4UNVJvXJ+yGa8Qim0z
Qy+YavDCwgtnrnxMzhj0arCsNCRW85ztL/030wij6KtrDJghjt2KPWat1k9mzk2DvDxaNnGEPEXv
852ds3FCx80hDivGsMKuqyAl2ow0CKmcwCj34O06H2sPV3vOJDpanSVEGLMlQoTgWoZrqr3D1zgi
hN5L3SwVDmZN0NUvLx4g5w8C+X0d75r9VzjKNsocoIu0qU8JdHoKjN26bQ0dek2foChjY/GO8n26
BBGsEOrJCSgFxtmc78HFc6UN7NfVEbfHGmYGMjSxWoPNaJkre+l5PMQI8C+g0P/LcqdTEd32wk5S
Hvasl6kFCbA/6TILFNYgJzpbz+pRMscF9BEigDRvloYruJY3BNhyRfj0u2m8GYQGyFdO3lZ8XI5Q
gDXiCmA0wt4YEtKl+tNsGLOcuE5Z2B7ncRBPjnLG9iVQvVIQw1XYoHrL47qeTlEN7whH6sdK/OG1
WqI5rEhopYOOk5DZVASZEhTaaL/okuOSpXb/jFZExYzIcG1/Ph7CvF33u9ZYGQoWVpE5ijc1JrjI
0/VjOIbbTqT3QBhf4HqogaM8UemPPKGyqrzV81LemOVBW1igvxmmn99gPn1NqjcYsmrpkWzjr/VL
QWLkdm7WLRXY4jmqexhgMCxXfuH27b1rNIC7IjR7sAcLjWU/sl7SJDnl/NZ50weGNqhlLYkfo1PR
hJqf53Rzvy+MgLDQ5I/ZCt9fm6HffhmwMx2exhNem59UxXJQ5IdWOIYX7u4erx1OLUdFZIEN4zxX
IiFvmHfKpjfOFwi7hutTKWjiuUd8bER9hIt3hYr8pc9uzAd4m/QGJtUJvFsIOTeIGYL9Tcfl8OS8
0qI9vpkkK5NSyI8vcLgwu/WBxP9y8HN1DmREnt8CkjgRthZKCVbn2xOVPaXtKR3h56PFfQkBv3Lw
vdYT3Zaq5bAK7VURBfZYxgmx5TYjphskQv4VnilyRq5kcn64Mrh0m4nZvUoHWWwhL5NbgEFxZx5E
Rd3fH/PZHqVtC3/hnm1RaAxtIGLrJiZ9UlNZCK0NRef+NPUzYj/v8rhowNoUW+XIlV5AJDJBga4O
NC8KLz8he5xR1nv62snLj1zadJxTnO0Z8FMhlu64yLgBIPduOlnWEbNBBkPFaL3QHpWosgO9NlDN
8FLwsih2yG0Tm21Ns7JiOhL9RR0/GaWMr9LR3QPxTjXmS19sUj8jN4+NbTRKCGesOPm5XLLmImvJ
f5rq2BiyIpHbR4NfWHFtpUHq7SDtOH6SOnDrRr1y/3S3Y7QKMtA1HpefRtsvSXRvMUlw2l0DYdRt
3iVhAf9p0UD3ThhkLSQueNloS8WNmWsUCbVNEioeFxTdPzd7w6gwTd26CCGcoy+a7P5vERSxNhCk
kotcOGjvnK5ANxwdFgcV2H3ViOmDb03OTOD9tDVyVkp4yF3EIENG/WWDtxdds2fVymp/5WfcMsbH
eMYEn80febjPGWnZoA6FkmHJNGnpTQP/zUVVdBcAHZwaErRQMYMa2w1kQfCfc17EN1XUL44eWlCo
xhuX4Jsn/YPfO7IcgKvygD8EuRkKZoEgwBYvd3KiBK+Xju2HGjREHmKYAlmSC94k8bMFWUeq+Kpf
kN/lEecW1XiGqiHpCvDz52FbH6rjxkivcorVfzMuHw0/28aQ+ALWpKk0NtL9rleNBeMM7zZSi+hU
BY2B6UQM+vAbuIKQnX7VE81ozjSbie8IFQfB7+i3i8R1oxovN7iYhLQo/qHpdOIMmz0sxKbtybzF
WFpu8u+hhAhDJejMcRV38j374maSXN3a/Wg+pSg8KUcRh+2AS3OsHZgxwkgowUi7eyvw4CZOoe3e
PSxEAmUmjiXyyJ/FiAlG0bXoRc6sBp5E0kg8kBU37e8CHLB/l4weZdcfDImFIdnZ
`protect end_protected

