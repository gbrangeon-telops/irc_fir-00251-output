

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Ksr82/EJdyTi/ZnocplaChIHl5gVfg/QywOs6WHQUUTVobYB9S2t7HfNHkvfksORtftr4wgSGG59
dqflxrTk9g==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Qqej7lC/8l20xFx7bklclhPhbKpE2SoVMnU8o5jHyjJozBFHGWWzSqcy2OHoxuRC4svtWcuXPZER
AveySsBsquyvS3CpwUhQC4HU879mrvq1rktu6YiGUKekxqqq8XWVjGU2RErpRUag/ydvNbNrFWxX
vuxu46YvGNDVpOq465c=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
439mpd6b2KugK1Dxw8VAcq35Q01RTqPVrzIbAJdjxQbya32eEZ7i4WNiFuVZ/MAk52bZBtBQiNHc
mNfbIfQciIHmnAXJEN9w/4VODhRIcUMrMjQwAjn4teKfB1tg762rR2jvGQ50Ai1Ml+OYADsAGJtF
URFceTs0yqpLMxJ8Ov/lGmeNw5dXmLiwn/XRqtS/K35VTjZyDUeHpQAr9q51KY6k59LrSFC7lxxB
mXX0In+fzXXlrh0dFFwLWzscDXHiKjrU4bwWBuzmrkKr3uCoEG0OADwjka6wlXo/Z2cEkTpiK1Qy
MmZH9UXQxrxTgtpOMmK0pjs+MfXf5/7XzeJsOg==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
porEUqarzWQ+a43o1KcgcLOOq13cwiYUyYcVmnYhbdWCiVlWWfN80U7oRzW3NODV8vTOFdEeX0/T
HiPsKQYOSEqQjf71FVXt5Qu85a7gangJ+zMjyuk8+m1c85rFqWapoLbPUbexfLeiEmybpwcybBzj
rIVwXl1qRv1R4JNRI44=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
s6/C7NZuQyYs48nVSWrZBvdUw/cGGwVNCnxc6+Wr+hB+GSdh07xJnxht3+mpM71wbe2jyi3JRq7M
A8Qq9KlqvpjZ87ZnAxTvr8P4OZV0DRnim60u79JqHUDowRtwBKuWK+fhBBqVkg+I/GuK0CQAje2N
3H5CzXagxYQGmhNBvdIDYAmWiG6ymENT9OP+fdf/JngSq3sbaQDhuOCrSGCgAWuZWv28vEMvXd4d
VKm66HgH4TXtJpDsYN5kTW6gEWdi7cV3KJRDsY6jA9RzwyOOBsMl8Gl/UvSGBWbIshxBeydyVUyg
0jabYqp6ODPXSowz5ZkW1y4reTS+cozycJAuMQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 11008)
`protect data_block
eAnfH6LvbCwHtxD/e+bM6r5f8xJEAFZ7wlE7ZqokKzeP6TuNFfdO0z4eiVZDhzjF9j32HVV3As0X
rL8hX/SSIrCJuT9pgHgj0QYpIyrkURPB9g8mGq/1razGjCvpvwl+ODRd4fOL1IaaPTp2Ae0XQLNj
BnCCE+aEbSTEvOOq/R/Z2gdgt2XWBhcEbyOI4L22L+AJcnCLvOjoneFGPD0Nlz67LWLGeUFIeG52
6A8a3eX1t1wzFHEtK8Him/eENz11kyHje6PtH+s0cICyrz1PRZQ8PorL6tKIVFMR0FBeRtRrqY61
TtTLO3Amu/TmisJHsva17dxzehVcWugaF+r7lN1h0Fnv0sYA2g6K5Vwxfo5jK8KjCxAoLvuBMu94
JahxSYQ6WjjL8dihn0O9FwyvwvRDQm3+8J7KMOuRXr3kh/+cA/9Tev9kLfSPOLqbYhRSIuA+NiXZ
FH8ORQmMk2tEX+yv3XHxMa46cTAmKffd/KaucNrdkV2LyXHFLKXKwOsGgq/RSai/gesCLpBXtHBa
uwJM6iHTRsAPfW2gJ61gtphK+TusItBIWzwmb4qM1edEJ5bdIW/YjcN4WaYKFXfn45nseI7JnedL
F871+2wCGkBFcw1iKxslgZeYxQVhn6jigRg+4t/xoceOw3+Ku5zZj5YyW3A6A+Sb8dbUl6rUflVT
l6uHNSoHxCqzNjTvpDO9E7coZO9a7YTha5raqYd52UaId+0wS8QcoMkydkkxPzc6ssgJJu/v+U3H
wvwH+YndQbsvDysAcYnwOZuK/muDnWMQyGNVgCckFiMse983ZXpRAUv0jE2RNGgQ4+DdZ9N6pce+
q56O329Bizb627M8FY0J8AiFEMxh4a56jxOgUqv4kiC0Xxatauq+SfmFj/e7vrWztJZTUvVcfzHE
M1Q2r8ujvGAI922YfIfW7uRFYw1v1/3GpeTtXGBHGwyk41l3lEbEccGCUz/QOSdGebbmfDd4o9wq
XMo3jUsBX1YU9cMEP0BwDabiHWYL7FcnCkYB2hMB8h8Hc0bEwXx+KjrXddmU1cHpOThGrjjLLaSU
2NAL5WNcIg//jmPg+IpTvutNiVs/L6pawBL4Y51Wtq2lZe0OKinTTBaSIFUJm/3uwg2P1Qzln9CU
SfWcA3wLj0ub/XeI7A5O9tshO/9qcBLH4CrlEf87UPmnZWG/PnEV84jv0dkdtdqIFdNlYHbAczqD
etaOp2XEIHdR3AuHxvAWwuzohDWiylZKWLg8/sfWGrrty4bfa4uCvz9Q0wrGMoDkT54ED27fP1Np
Icw//8o8Z7/sZdyeot+1GmigxMj9MZmMAfBFH/sxIClc8RXw0QxGPNPkdAWE7sDYo8gkG5Zpyarw
eh1aDkmUtuoi6JSM9YboOdgIcI3fEIMo8VwxkKVLi/Y2EzG2oyZDLiI8Feoz6OZ8kP6/NfZ4XZ8v
99CParJPE1EI64IaUiFLhKVN4Hzp5JxD0on+dS5HOnolPr4Rr09Xv/nZ2yVDadWnaHT8WRVWmCja
8ElModTruWGhivec3GeD3aZKMQoLSJ0aEE5xCa4pHz/V47HPuhkl6dJZQvKAW92T8e+ifJ6c9MlR
l5dmClA6R/X++/tDBTCNKiLcDJwHy4JKH6S6/tiUNfgG64vC0fBylh7VNPQQwU+FM7EK3U6/AI1f
8lbkmH2/oNb2e9TvkLHNYmMwzJ6oPmlcOKoRRHHAMz+DIAdNF0IontDX8rLu+LoiQWOn/uf5WrxC
VEqHpoqpFxy7FBWMCHBGCVjKvw0CXJ6jup0uxgdY4mAylEFEEBSmKPUGm8kO5aAPwS6EO1tnHDQr
NTA3A6RiRRMrRdB1ZABU2/ouXgbJdcEeBoTaYOvKZhErbE1/jCIoD4ZzpgCcrQGOs59UgS1YmJxC
KLkIT1rF9qPDSq9G0HVSvHfwBWggGUe60Bhx6gX1XDP5CiTs4kTRDfR+T+8ajossc/gSvHeG99uu
cRrI1X1BW00QI2stk/iLaALxiLUshQ60esxIPx/KtFzwQ8vaN3t/kva69FEqinjPjjcBDaWx49Ej
QGXM4lgLjMkHdwVhQLLe0y/I5SwXiV9APTrV8gNs0FMns9xjD1xZ027n/4ZY93FEGR65Z1PX5AQk
OcJ142XVsM56bxzE+eDreCzGwvaTB8B7J+m9GhXLvI3XjpQxaII4gCDP8qRhNV01A1I7y3iuhH4A
GN1I0plQ9q6XBQGe8c4is8aArQyURGXwl+EQi1GOFAWkfMFQVpF5zzn4CggjkVB/3DjK6exSCxwD
OscogGuM0BoVQ2P7gENC4XEfDDlEEQMD91DVW6SeKYLnqn4pT3Xgys4KLHuH7udqtmevQ+3Lxeqs
2fpQ0vEKidbHJuUvZb0lxlmf/sSGBLePpN0qH/xU1dqTP0/gLCqWrkDBrgDB/dKaMwC00UoQfuo1
Hz6QaaGgrfwzWcqVIfoDYgokGGKo9022xYGYIEZdx43A8/tg7kBHqfiA8hk+SrT2GdofzsqWJLlX
f18vDAR0PjlpPAP0tHoLK8qZ18y4IDG3K7iVHd3RefLHcen5WhSzEQrWaSpW3vZ6FqBrMb5UEmr2
FqIdgAoBknabJ6gUma++4XkZxM3mgyfMc5IGfv/DA/o5AQIjcfi74V7mi1Wt1HODJWWOScBcZWl1
WfzKlHl8Z2xqIy59/IFEO9W9Kpjf45LcmzmBlmAHoj3VRUSgdRjtqI5Pr3GPSNDsko7l80FUh7Dy
fDN1Ktw54U69g8Y1h5ghD7LIHfh+FmDlvTdiZBmARwrUaOMmJABQyj+DZEZiK5ugA3qVM6XbiH41
jeWqlZAv6g8U7q/heqVdT5N/GTCboC4kDjGIvVgcAAZtUayMm9gkvXXWGLgo7fc2V7c937g1Y6at
fAtDCZ26Rdc1WEIujSMc/xN5TGfNwE9vtSUywwk9KBrt9UPQWFrm5Cjiw8M/H5Z2tdvCpnmypC0Q
vCjFC60J7nDKJoCCoJMU73t9xqv4MXhsFP2BxcKEZA4qiW7nEISq1uStWKMrNDpJP42bXM9JtJ/I
/zEFjj6eAlkcDv1ZyIwNctcTE8QWUhoGONhc+Y2VR3AKJBVUGpCcX2ljVpDS6i2SV6o1dAtJqFlO
z8cV71a5CMi06ezYfYFxdHkufoII4+Vq+kJtwy+rI/hv2S2uqN09pu8A0J5P6cHXLaRcHdFsE5qL
aUWNQ2hBAOovdjHuskjweiGjWmlhYADBk+Uf6RBAELVpbqqRPAjDCTwB5UTlBmYVDXPPjOXkN+NQ
BhyWR+PWb4Tk/Hd5i+LUpdCCwY3DHrGXeHYo5JRzRLeeghX3arkp9Dp75TDTIsyhqnYW5FtgINqA
/sOxQ87JRZFAxJJNSzU/4DQLdsBOqkZhKEzyt/V2nE83R5ERjEc2WeWVWu5xTb/ppD83ckwP3ajw
pOaeE5Ydz5ysUyRXVTS392ZXuQ27lGmKbjYn6OLyRrFC7K/u3oCZGNlt1lvlUcv7W3kRBN3isylL
yNblYrELaR4yhcdRukB9DzwRweIUMEfQs5ptWwBvMhp8vY7IiyhYNPUeWovThBxacvYiIJ3oSMpb
awkdwT+1pnANL1W1SRMBnXxfaSXD1RloFNOwdhq9nlz2ZBIGHqkVJWlXsTx745uoVtGW9xu294jJ
20IJ4WKjX19igVzg0OFbmP5FLmBAhTrQdjyVH9+s+Bh5deXGA7uf42CCcmAbesksOh3KZFDbk91M
jNJM8S1JLLiruat/0DJFl26dol2705Ok+h7EfrjehgaWoeMEoC7Sne+fc7s1hnnVmS6O1JtFC2mY
5lvV+VsZK7UMT2Ju5EkugN/amoVujDtFEgZpaloOzCOSTgNN61O4vLwokv/KsVEeRCy2beEp1dK+
re3EEKeb0vJTHsdL4IKT1un5AApa6r0IFR6S8qBSQo7wtE3yTm91DOCJIJNF5VadgSIbXrvBbH0P
nD+sFPkp75UkD1UHw6hu1rKCBxkhsVu9yKtvlWTv2TCvN0KkFg9Tj2ws6QkC+ooMb035mJBnbt3u
FeeMrNbNs5rqmhwCKJiynr7fmojWW7GTszkuXO12TGjF06krRUrBShzX/ymrzCU7oJJqXjK/7/vb
DcS9e/yCrx+5sWLSg6nhLCHMNxXjiTCrsHeZCgyvChuQ2vQssKDuwS67K9F/4HpykJX1DVM7bzZp
Rh1f5W7NItpe7Li3C4VOYineTle4IcrVQQCkM2gKgWhbqN4o+0+oFcVcvxeb2AlqrGcfvLdcDuVf
+NXYWHjsOmXaCNPqMHGS3tu809/Y5ubepnthLAKhIDX50q6RouSJojhfl108VuLr+YZs/RlGLJBH
Iv6JIweMg4mK26sttRYRBTWzwAgKgPZ3GoI+odpOrldEH91b6OuFn8InL3HBA+scYVNJzvk2EbbI
caTDVj1JSiN9spcshNygIPxTHxpn2MdUPZsAtBVRoLxfWFGWHpy/cOxWcZxt3GAXAC9vIutGiqG/
4JJvFWC+l/xv2+QXUEmtChlJi98+ta5wxp6i0nQk45A5js4THmoJfgMIu9fN+VnVcd/obC7sxpGv
hcQj2qvGHIDvpEt3ouVqod9fK4TD6NqE0m0GszaCwhZLbBJeNcbtcUgPAsMCC1hI8cIN7AwJQX/h
ZypmaEtEdMaV8m3DP1oMy3tY8tDLFVROuPuYe591Zmn7pPILMQUIM6LzBJ3WqxAcR+4A7pmM545Z
JdPP8Y2kKLeBaeNbfgxtnW4xJUvS7JpUsOd2n2k3IJ7zSBAgf3bWaLkXLHWTUwUIQTB4nDUC9kWC
Jzpf9+z0piUhS7B/oR2xSgpgSl3ClhDllEMq7zKRJ5p+QgEFo624dn0565qKAjsRHJFmUZvpr14x
3GLUND6XOE1ZFEJb65b6AkjNjRrJtm8Jb7zR0G/Aoc8J9xoxHMFnIXV7YViHYhe5yHk3/lKxmdUt
6vFlWhEXtBPN+8Fu0KnNtsqkwy9oRKoX/3hi8D7dTLrggCLQK1by/gI881VXFNH7ApZjJYSYVthq
VIZowfegFd9oMdHwz81svf31RMQ935QWlk4cgih+P0wqYGg4vT6YcbMwylE5U6wXkG/2uCNPR9AT
hUwW8QVt4PiJjZ3v9iXd7Ia1R16YlwqzQYjVfupvJOvufalTNJuikIAZ0qPYAcZrg4Beb2IYzCMB
oLN20zd2hM50p+bkm5T9cIsLcIKsY2Rf24aHv5cO87m0OVZjXKIG58cVBFBCd+5Uv3wc/V8/avHe
C6FXvH+13IFVOJKxSTZ5T6a/VsDsKzrb9EuZ2WOkFwmxIxdTzxmfEzQeuJSyr1m8v72mjkt0R8H/
9gsZF3tlXw3XiuQWPpPfh1E8mqLe9NFGByXoYBqCuVtU4ATumP9HPD8DZQ3Wjjfh7BJlDeSrDXeP
0BhYB0nqQTry1+fovcfOGoo075iOJQwrLOqF54xrZbXwWad9DjLG7cM2bQ+0EZAUINxN3cpFHwos
Wg/pzZXvsRyHtA3QKTdr9EhMY4VeJVg/xV11RkIjAOSamsN+l6Each437SHruHyb7aIx2dDxvPkL
CHXtyZkpKMwc/Xy3cwGKVDOtHr+IKNic815HAYjkAi4WakkVQdmbLe9m2uKRbt4rO1mhKs+kZV3z
5Oe6InpokVRFcdEDcMRYq2f7rlZtsIlP/7nwbB+PnwpOlGJzHoXL/q/Gtt88VP+EipsNa/VA49dE
3OHpIbWEyhnaMnTd3Mls4oNF51svUbOaAuvkno8mychMA/XZl78jBe7WRCVh34tLmbqVdzsNkACt
fad/RVTRPVhDQlUAO2EpUulhr+xEXvE2/cyUvfNPaTSMU0YpopZmXwmv+KcrjO2KdJKX8jRkwl5d
2iDtNyeqG1HSnmFLEsChxhoGPpxzlGbC5A12pExpaQYJ9zTKS9tusSobYlgsy5JWj0qJ23BHjVdP
dEgzejFWfmMEq8Vs+FAdE70vhMjx4HndfdjGQeZz8dpr/eTAOegX3F5j+PkhvUB3cEr5mwLywE/E
/8hEHE6AIaJBDB4DPBhMoR36rVMVZB4aiiOjxTC1gLTlrCRMcjv1tI0G0b3gltQnChoVbe/fS2X5
1fcBm760K2XLknJDyQY5Co+VT/3DivNFNf/XCmOfS0O/5Tq0n7cUmVU0VNpv/TaqW83nj8pNzGqF
niGF1j3Jd4M4TcmHJZhNK74UXqYpawZMCHOdlZXH+yjrzRm8ZegIgeJCqGcIQRXCnB2TaUqnvu0g
sQIFjkB0VcuuPGr/vYusrw2kn8f57+TQZupr9KNFkMK7Nk4a4YFe5TiwoRV3+6v4MDFwQJS7o+c0
3YmoE8C0cUd6ALyMqxrolXfT35YbKuEjt7yJzZbZWJixCR5t/9UxHV2lTCpJaghKYLQ6qDfx7Qhm
jWJDjAQZ5QNFiLikq16lXYS7q1mbCmAcAWGiI/pV/xVPdDJu5/PLrk3ptyalvFJBdn8O/9ZonH31
78R3YOTaE91C6MTZT7qdbDjJXPjKIudO0diyMz7Q4v6oeKT+pOA98h+C1iLzbbHcTijKgyu409eP
BIUMhCeg3H/uI3qM2QeY7sX1C8OwJfpzncxgCzMk5ceoz8PBy/mx67mt4hBtJJATjmQL9Ld4F9tH
CQntK3AUPLYpcC0xh4lTlRGryzt3Y6GAvXQg258VzumA00WMSpkr73ywn+xsIURxLSxCRHnb457c
PXKRVAwKLi90M4SiRw8bTAPx5cMMcxnZ0if8gl9HAUYtatfodvItuCx3+x54rtWuNNh/eo1Jqqbo
xFIjZtIJUE6/bfQ9CA3cPljzQEn8Nzp1yz1ALRKGF2ijfugposqOCvKYcglPNeJk+BBBBbKLLR38
QYOTu7ZzY4iWvPxJ9UCNW2OCVii/hZAaSZHkVFIYVqFFLfRSIu3v0hHfrSrPjT5igv5r/pqBl2B+
4TJtaEZKZ6R5PQEQOyY5I45d6+mIKvcot9TVsBGod33kQr3wCEHXx7wZzvqEuKLbdQvRjX8nXJxv
5cziZDgzZMnceNnOqC+37h67GoMEApQ7tS9F2uKtAV+gSW8WFyxoyXUbfHrdabKXOtgOGokiQZTk
USor4KpDPJoJbkSMLLTlGSH8rv5qArARIFxT3mC1VXLVRenEljvoRuBq1W3Auma/hrrozmQNQFRR
GmCtzDML/kRt85h/+6F9wr3fgG/qslemvNenFPPAnh1wsXdAPWp/Iv/DPkJs/BGLlD5M/zW8TUBc
zxR7LtaAEnB7kAbtZ45VcBIF82IcWNfZiIxqTiXQ3Z0kp5zxcpblRaSOHaCSxjEKETrol9/iYyFG
whq155EiOKfWEtF1zLDBsdxyDgIFD9ME3eJwRtdUvq8VfB/uiJnY4ee0tgavTbXvoy26BDVGfCpL
lD6VD4EgPBfqem1PDnG6exOtR523Tij2gqxPJK2NJtGCFmRU0ybMEkUC4+sGdRXftTqRMuTvUMpW
yspsvtmmIW7J0uaoqEaRXZ4ATT0/gYr1up4GBaeEplKwiR5T/vBFKLmpVaHWmI9FnHs0TS+2jKxp
psdqgoVKADguOrMcOfhcc341IPukep1DaUleSqXPwcr8CXpPQEeimQmWapwcuDgcretnWWA/RmPr
eY7ru1aVC35LOmqB3pM6tQPTePZVMlDluci0KsWTiGebxe0LaOD3PEefiCDXPz/M974OpYox06h+
/v3US+J1GCe4F/ShQZwQHofzZ0jfjqsa9lrekKy7B7wHmm8RrVO3okDQZckp17k5V33D8IS4MF8q
WNvsUlxOX3tmjn42Z1uVNIZzKTuCc9vjVeNuuYtMMZs676arM21h+vZpB0q0Z3Q4W+ELgpvuzEbT
KQUj6fJ3MxhMBrtyvbUo792ABJm6jKLJUHC/caO9DLpTOYylduv8oJgVuQ0JpQjYXE90CJbxtEGJ
La5TzfbveRrJCPb/pOKx7rnM/1Bm4UVbhxSdMXSObvwpe6q1XBrRVtDLxa3zrbY0QI3Ay4nVMt+w
IfIBa0MZ7Twuof7oif1z5puNKGHtAYFPkedhX+jMaZyl8To6kd84CIa30QLmsa7/K6K2qJwMagEy
/Y48sGsuU0ghjEXaUZLqMTf6qjHEeffaPJGQyFCT5TLyQxl2ZxI46k2e0RStF6YBwXXhRSvT0CP7
2NGbwWVvHwGqL1EizQ3g4l7NVNkm1FJL/saRcO2T+aeYwzg4hRbgzr8W/JjFETo662lZX2DWPtAC
6iI5AVhk1N9X83lkUkbwc6NC3VMbT3BvQrkSc6DWqHQsBqmbemVGzUSJYXdwf/MahthStGMJR89n
FXlfFb7Nveo/tOb7ItzoXQOggaN3nq16nIe1Dq7seVOoLpjwepm3VUYqzj2NLIjRf3xhKtOA/6Qg
G+APNs+txnf7RbRXb1qf7XNR+V7s73VkThQhp82kFo6MqXBbXd876dQhKPbPGgUfuCemmMQA7Sqz
Sfy1ROeCq84IBqWtIVJXSjFtJ+86F+QgYx7Kyf103O/lXaz148SaiCU6OdxJn81noh4SkvcsmGET
+SE0pMDhrSmEHOD7qsUMrOB/z6w9+amxD5HpEG7fc3FkyAPsNNVq7CyrqltXCNXl4vusqKdTs4SU
EQgYkutZsyDybB46dsFWT8MtY8wV99ldE02c3hkFr55sSOhE/kazMJb9HBhFaq2aZv7qmBazvx13
/8gtPQ8HrmXjvP7G7dsVaH4mLac9NwuwKjVL86RbC0S9kCFEwfVEeroaPEFSZ3CEELojzNcNINAG
3yKx+tK5MfHGfxU6foJDWADknKcLgSXLz5Rdeno/lasVtnikBNBOlMvLLkLgHPoBMmBwH8ZW2oMT
Bl479hP2VaTzH9L3OpNaZkcmldmvlca3S183yF3neFVIbofPc2YSbhFlh70pibLRn05ah8kOg2Gl
h1sVGnO5Rh7vl/Tawmk2kcbobMDYoYQwZJUa0VC0eaDpSzTle+BrprjxGGbyfthkRWjghC6PKsoK
/IkoltMm+Fvh3Ui1ztDG2aoeAFokp5t4njCXv0v/fkaJbc568Yc3xc5q9FMCBBlMy2ZjKdnZo/p6
F1g6Rzj8pAA3VfYIjwgmwRhP1x14Ae2eamS8j82Q6J6t/3UNWe285UE83kE+/eyW+eJi3bXX0Ixa
v25StTTokegAsQKfD8+Ru2QmpTXXBi0jg5V+Y5Gp50OJKo3GdF7TEVP4iD1ahUn0m1sDCsScBQDs
QjbCvsbbROEu8yMtY+OgfAfXd+lv8iofroK+c8FaI+2CRs/MYQQNz4rMKMxddgIoo5f891TLMgiV
i8PXMvPNJ5sJcHif+wsuO01yE1Go4IjSoKPzD8R9KB5QUNH+lB4vtfNtVuwKq8Xa+0tnE8ERszeg
JJF4srYVWjzmBTxTWxpyOV3ysQrF+2feXZQu1YHYyU8BUI/soIvP9HWet04RxR3ioykqwcXeFXjh
ktOgqLjeV1cPlOgKiV/VZ4XcZJ66iU6KCcXCTE7mOJ/A5OBid+fzDiSVck1/kKVXLU/3GlHUFVVd
05I7pBR9L1LFiGMo7bjdkwEZjuJq7+OrZGCeCfvziVrEoIbNTkaDjL7xTNKyv9bFWiup3C5ed03x
KX2D+/uFpRFK55fForniO/78QWViFevLFBAb24pfzLifElNti9VXkq3ILuOgdR1dmuJ8dDIdR5nc
6Zw3QHalHjhOfKicyRqpdisgHyArQj+2vcPwtFZ9Nlfrhh+3XIvZF6fMeUSPE0/Eb00oT2J9NXGf
visfyj/FOCDeF3Dx9JxoKOOA3TB7UZwTZrwXxyQlNoxY2xY7qz7S1gSgSAWCCH3tZ75nGTpdxkIZ
oKCKiNsVnOZcbj4S4u5J5GZn8/tU4xc0o1zofbk04e3GgmsxM6p0v7bxC0unJ7zpB6LVBpUYCemJ
sKRJQ1y1HywnNwLvwimR/n8vdQphwPqexErdJS12N1WwRpmmspYuWU9I3I0U0cvakxZiGX2qLqQc
rNyTcIXbma/ckAuYNAibORqeH1Zez2HruDzyU73I6TaL61LAzgbDkpCyck9uEhgusBbHBXj4NuRj
MH1sDTpi0a4ujSNCk/nGXn112cnJ8YkR73Mlb1l0+eGnSRM5XuWyq8jXM9SwhMEs8zzQSf01LEE0
U35TpMpG2Txf4guqCG6dDQt+AFRKKqhf9jujN8Ea/DqVpqgCFYNsUDuAKy6XdRWm5ohOlTG3WF6C
ZO260yFUkBoY9qU1M8eDeUEy2RcGrXjm5efbGadVV8QDhFgotesn59OjEDhwLM2yIDsPS7ANRY4+
LxVgy2vLue+GnYOm0jMXFkndscLdUn7BJzsPLDCgYpNW7KLmX6FHmHhNZcnWdQcNJ8He9cCX8nI6
5nTYEm7SZVlcgeZqup7sp1OjBXBj3/F6W8Sy7t6yyOydl9ZgVbId0LcT5gmPrUFabXvib9rSesw2
ZRhV/4y1UM/cwIgvnsi7lRxo119Ch9K7QW+dSosacqTZtT9Um72p3WpuGbo+wDwJ7eBRQn3LVfYQ
PkEFy6oOQoshFYDiHDavBClHXjmSMc3apPS3tPd+qjJdHm8lf+/gM0IBgIQSCzoUSqpFRzyV2+9q
l11Z2tocKwJ6OBdk7on8v8TBpu085NBQ/two7QRHGuaYDPI/VUKYEUiaUnZx2CUODFFWGf5Q6yOz
Wucza50ytt5g4IzHGQlHDOVceaXdq0HiVLHjuqKqBXoVfqW3wILJRtSsT6oYJmqrjczSMr3LYLit
PqluEWuudZym7Bp5dytCh5+qYm/6X9IHKn33czu+/Mz6smN/75GqKO1rMEXfrROqQCfCYT9jBrSZ
YyjEmFwqCp9vJS2HeIQqCVN6dMzOr2c8OXcn6iHdRDmvB3x5PbosEP7ZC+IR/ZiQ+SgaEwwhelb3
Zc0vX4HGXzu/KzBl5i/gJRS5bVsd7pZSVOTXla5db3F0fMg/z3vUtaZlbULLffyOcx4/6MlG3P4m
WlqUdZ0+nRkpHFNOjqzq51R7tyb9QClvnrhOCOju5j7a5KFFmqfnsrMMPlGyWOLyZhKdU13BAFxB
tXVvfMJcJSftL05TWZSnPf4doZ7sR/YTQMxuIz0x8U7hwJf1644tQXFEjGrwrHeWTRAhtsSMg9Ff
Uxb+uSCQvdluQ4MWvArGieQXLHaEYvACNB9wxaBh2GJ8rSK7Uvt6pn3+LGLZ6dtxDEOoFh/uPUmC
S70WqxcS/63mK8wqsH6PjuAKHaXB1XO87ajVaPuYAIDNF+GYqD0izJU4uIC6NQ2xbg+EFWqt/zVc
ybXmcfge0q1UzXUYjdNCpBzZI251OFOm/EFVQllqnosEutvOlubWFP7lwQhnKftTTvQ1pfYDKLRk
eMe4hAZf0yhsnoa18OnPD7Q2ZEzKQ9w/dQ9caL8wsfXBw0qnOW0D2aG+SO5iDEs3qwty2eKSGeI2
RfT00HUsxg6hufiSYwRZ+XqA9AcaTlJ+2pnx+oXvjPDa8VlZ0w7NECvY3+AVOwjSQ5l5c8us9Zll
06y1Oxa67L1MBKuveFtuvkfJly4jHhd1w8QuigF0Gvrv6CgnMXeEYqBk8bG654VcFznkRrPLnx0I
PZsjt7oLiRGfqCGZKLjvmEoHMOYHqKrtLhDNOxTAetfm9LyVHcQxMZH2spuChqd32ZgCGk6wc7MZ
zGU0tD0SLROgX522Mf/JKEYXqVOYs1jQAg7rsfEO4y+AWwCKRE/p0SNl14JqArYKuHP4ugcT6WEo
Jt++bxdCKVtf1ZXmMBiZL/BbPZy5VEQr4NrL54Y2Vooum64xVnT7IJhcb2SJwMoKeqVKALNULObp
RaiPlVVgmMgOPi6iQBLtSPA6zMB+/uu43gUipfJcipSRts0TurkGIL8sSsl97xaKDHqFiMWKEX3I
45ro+R5KCMeyWoWdZ8s9d5R4xeczqKOi5FUKD5XYvVfp5mz4fc+A23FTEs+w0HnQk5KVuLkdCH4p
h1Cj0U2SxCae0MeJSYKeS8TVdVModMi1DPt86NMBanHcaKZUeHblqIkJv236OPFoRyvlCbpBRjr3
+qiB5gYUrx3OJMKZD816XMTKrZvjZuqBMe79aaGimWgjcFXpIYI4BciQboyD9bwM+57Ve3EnA6SI
NCm/idwwV5MPwKmD5+WJtUUtPEZixySMwyKhMm3/Z3DRKZL9nzJcVSbvrr8oGF7JOp1Ic4LEJ5pY
pRDhes/sphGINWXl7/LLlKNRbVhD9p+vZ6y0uox+bTATSl+LlAALZGEpM2XIk4rC53KUIpe96FaT
kzol0vDvONH/bSbPkdr5B08B9gRUeJ16tNYIF5WaC4zBamEjJ8NgJd2BDFf7W6b92Hjnyhk6qkVg
Qmux7qFhoMJYdIHemqASCpWufQ3AxTb+0XMKKhpskZH1PNWJBFlb4oGzBvOZKjFcmXYvojFSIteF
OEcwK27itrj8tydNfI/pMlVGxDVlP2I+hw4Ao649F/SR/kt3vrAUTY/wo757G0XtuFu8KIusYAFi
ON1qy14QOYwOpaVKvCB1l1YyDDDuH+8R23nMfqFvIhY54k3V63wkygwofh2khbKGgB4mGNtf/KDb
PUGSBUqE4wqD/OngEVAII5rtLzV5ipLPSvTQOurO1nzTo9XPiQuCJTv+rgYYlHoYvVaCg+z0VJUW
3Duq1HygBkCUl+dw3WMfBbtAT5AB5MeF0Cd5EUTP+Fu0HJTI6ZTOQvqaDxQT5z6BbKctC5U29ram
yqpoMtWU1U3c4dNOj2hbMpDugL5UuL/edmlLPaAtPGzEzJC4EaAa/0J62opV//joR7GD1dsGvzSG
SbuyZLg3z7GdvWjg+zFKIKhahQX4xZMC5bbnzP8VH+7ttB5vi/zy1HQwiUsAdmfnxDNIBAF8x/NL
ED45nuitfk7kyBeevVUwcRkw+sddLjPWLv7v1qFyfKSRKGGGK+tRHVHVUiFeqBnuFZdbw0cfGlFM
LkU6GyNBK3UxiESvQe9I4Ggrfj8lPDGFbiO8b8pTSyGaKJGKVD4iaccz45/07pvZC37WnE5cqtiR
m6BUOc2T3suyCUpVqvk25cFMB7SpiIFFGRiJ02hZVAK0jm9j41oaJtKUeVRlND9UgcTEhOHeLOFw
dZYz9bGHSzwq0N6Ifcu8M2HWQp1TGsiit/cm8ZTnU6Md0NaYdLfFzmeoN/RMKLcoTeEJQngoFTSn
oUlZvvYQXKztcT88dT3MNoTfu+bri0Y1UrXBaKpbrfgolmSi8XrR423Pci6cTxLPBTVLl9p+6Htl
hrWW6q/wNQqi4VEgBElNzG9TgG1iDYyMTrYr3nyYgd7FFrarZLsNyB80JSjU41qlQj0jq8KRIvHv
tUf9eDBArRR2a3pQFu9EDH66zJ88LCouLj82ieKSkPfdig8aUBt3HG14fqYoiLgXC13vvuIBvGJF
fRZz0NVrNAJMM0qUKKb+QtSPrx+90OA7ZUrns7QGTde+E9GfBucY2+kjPmMOnsY2iHUSAakssnq5
MMtv+46pJA1IwOSq2p12aaQUvimDiKCy7TEqw8wZ7FEQ0NMe6bP1A2sqS480AQumFGttiCgej64U
6/0XzTM2tRztnuTg5LUDouG697jxu1y9cg0BkFvD/+EOLX2jHd/alEY8LuL/jsXZ2ynSchudTBVx
KSpMCmb4I2Hn7ZTUQe4HtZagtavLzDbDJLgNVHXBCtP6+KuEXsVcrRvGcQnCg2y4cuwsVoeJExI9
f8MyXioUxvEZEStsgHEPMLD0WAYajiuXR90OONfHi+1RzT3mp9rpz/dFNY07JnbizBtFZJpPwthp
6iydmCI/bHUBo5CKV7vxJYMKakLQzLEALe9QuFMZcxLSuld+gBxpIm8iFWliJDND5whqK1lGL6MT
7Y6KIBko4o80mKh4dsVMjIsVZiQggPtSmYJIQHpH/CoObnaAjCVETyuWX4k6m/hWA75PONh7QdpX
cHEzZ9tFdkooL1c8CcCOWmfhZ4+u+jCC5i4LIKVFzT9Vf9ElvigE2qCVZjIQFIoAeelDN+telLDq
OhAaxczL0Qcr2AMBKUwuqfEn1b1SGO6tiRGxmPfSX+C9lfX26M3yyrNQpKXhSlgWSifezHwfpqq9
Zy5WLTOd/buv1CEM+ADz167O1ZzHRc/CsFDxfQYret4ZuqOm9Ic86w7+1uTwIKPp3lTun+aOjcrT
yz9tCfIjfOi+v8M2arfTggOYZ/kKK+c+K9ZguV5ro8rWp5qDSSuuopbuiAm2ZpLaaBa2Hw4dBLE4
xCzv+DazzvGtRtnXyp6UcpHKyDWKNA+mMfbJp9Kp1uYqFgrg6Up7oQs4I/tLg3F6QlV3PM7IIl/w
Ouu8oWGhEbuyKx+qsPjor8d/UKNNJdjUWu0D99HPF1zvwSIPl2Rk9vvXHxqHN+dQkEXGMAA+WQf4
d3cIsiGDZsmlBpuDFnjSFmOCGXLmNeh3DrNKhnUI725drG4FsMEwc8uIaafME99g/0XM1E5Ob2jJ
eLJpO55peq7gSvjt2wkUkFF2TuvR3fRnPqNqSDmnNnWGNJyKMTtCIiTyiJbL7yl/9/98lU33nOYW
6TKZ1dh/gm+DPCCNtQna+R9zdo9HH48c9Nyp0dmDSgFb1KTE2aLZ0P1+vtzHcQPN8wdwkzTKV4sV
KQZ7M0nlFIblPoWn4YLklp2tpkNto/GwEe2Gz3R+2H1NfFgSWvGeEzcO4CGpEAyzYpX++zW4goch
2LqSjLVM2A==
`protect end_protected

