

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
DZrqnYwqMkKoBvgXgaWSB1Gvc9B94Zr8xHWYvXS3Yo2in98iiVsrSf1RUePWKa7hVSyhM66u+GP8
6zam55ovJA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
paoR3khjnzY7oR+WJ9YkW1A7ZzfFLvvVEXiP81AieLlGnfQuqZTzy9TqIBQ7d7KWJF2u8/GBJ9gB
S/XHVoSTyo6Jte9XVVsqnnFiHxvEAnWbM2e9+Vyqd/Q/lFB3TCGyLNKIFNdGxyml1xea2Gq/DUf6
P6PVaPylNEwivSbuc64=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
IuseMdZSknnKUME+O/YmMG9MKbslcWjYg4y9t234jonRTsM/8uUOZLlJPdAz0Ojsb7gi8Afg71RU
Er0Jr7fpQJ8YMMDdLQ9qwRqf4zAR9ZhntG7zWMIroK9jxtC2bvBKKArJREVpkzOWU1g2+f7dJ4FH
ubSzqp/ur3VRiEL9rSTe80jSph04B3Z7vLg49YvLUGmYKlwP09xV4/46qike4zQtuofkQ8/u3jTv
rlLcM6RtgeLWfD/CY/EWIIuhTxeQiucCqPyYilV1cA55FNKfdMv57PsY4PVV/CwLFMYY9INUTcQ5
vlvEZIaCBXiBH5TWThAkm9erewSr/bL5DW9PTw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
cyY5ZPlO3Eo0cmsRtMR6yuz2Eu2e6S2W/D+8CcC8VsHPfbx1fHUAOMrMRz8rOeXuKPOa7h1hSFcJ
XZ1TcAU5VIvCkM11jW1o53hK8qachmkkZZnfj8JtjstmyVTyWri5LmUnPYRufwJmQUQ0xqMJytkR
VTqDp0ZVnyDWp2/qKN0=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
WAcKeockg4TPNpKWNqCVvf1P8zBdM0HIqALOQnRkxsC2RA2Dy+P+XMiOG7cG04xrgm5iFejfnqcO
5lDRzw1y2vm9IxrTgVR8u92CBfbBU5si2daX0ciu3+tUaMvbyjjRBHmWEJd/+ZgwpEBd4jKx2KQp
YmRUDFYL5WDDgF6aGgbY7bniF7p7fSFQgxz06UbHJt/aNGcXnfge+DPA60LgmbiAZYAbqv+bSmqg
gA91XQkI7oyEKtZ35D6ZzgJ25i0EzUAy/u4ctGTC1xnExC071TQUx8Fakynqcki4h3cwrvs6RbsQ
1XULS0sNZpYYdAavNOXALBW23U6uD7bNRcfAog==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 33936)
`protect data_block
rVfLZQ3CJ5vyoRiq8r34MVxvTGDq9x3weOWbmfE7I5R57OyLprp0LAow7kBsD5jagyk0HIXzQ17b
szQyW9SDCbdUditoVP4GPAFl9NjzqfFevh7pQQzeoEWTRi6BLzVdYlmp8PLOzDC8oZkLogJShc7V
fDEX98R09q3eyhCXX4DAEFxmSAP1CzsWb/4+vgrl0wZExHmni84eul3orrqsuLROvFvH7H9TU4k7
nADvUDjqBXCzBowP6oQRG6hWEZ9dJysW43PBNo8fIugfVmP+NpI9Ck7EHRovgkHx1lQSdtpW4wmm
XFXHQwTUsALAN9gSAGSi4vck8BVcXv6dDqwOrlzRCpXFTYroX58kw4mkNllsJ0dI6DcuWuxgjuQn
drb7VtYToLqGL7Lc+RuSTv/qX3B2HIP4fbgC/L2kNTa61RSgS0XdcZ3VOMGoc3B3K8qkWDUXUOeP
25iU+SqFfhXOd6B1qvYxM+sSJw7VryA2S1TxOL77UEJ2kW2HxBtV2OSp7GKJkO1rcU6EMR4WHhJF
ju5UB7LP9BoC4Pj4iUPHApd/NUoDe0S45MM1WoipxLaoMBdKF0NScaVpuSMmY5ak2PZJZ1L7jhxb
EbUBfD5k9pYliWB0yfQoA61Kg2eI3NhrDNKKFi0FOMCSQpIwclp5ze3b+bDLpzakRQu+FdNYfGu2
7B8IhtWrY7OLrgcW4Yv1ipbVW/fmLS6QEwAGhvmmVwQMPuu2nmiwcrlcrUDrVDE4JX5vA1QmwRI2
tt/AAXfsY6ndI1UnqCve0vhgxUhFRNEvCegzcwxUvZLrpyfa/iCPeFhIxOf/u6qX9MHZiekGmoJt
K5qqzFQDNJUvbgW7jBkQM39N7WweuvIxZVtei6RE9zZdzT9rE1sy4h5RunOLAb+UVGCebet1OC1o
lV5ueBL2PL/ReDRKLN6wiYrNcOdVFj3Ww+BUeWAmP8jRRQ/osUB62E2zVnCFXeNiz2XiqZrZ7FOI
LflSddTb80YYTyfvGVi7KKV0pqXU0XReL4Q2qa7hO7CH6YAy3eeXshanP9LYPKnyFP2AZjNNROy8
wv/IIBe8L3AFL3HwRE7DkUOr+VkjhvSLG+ESPKT6sGTjBtGgXp1H8xIVeYIYBQyVfO6XVf0ewG5m
gaVfq6oc1C7vK96Aq+xsDstxPbh4CTYTktdPPacSJoLC88NrpPccLsfxdxkxSKuONZgyQrl8ecH5
nJliP0PCIAnmt1r31kQzuhkCRj5kOlF2wtUksETZ9THZReL8FJanvjAsJz6Qdh+5RGLi+xwXsYKy
EHq1I5YlNyX0NFls6elOCBrLVPyxO2lZwtWvVamLhl+8Ac+LFU18D61zhMywxUkp1XL/IFkfZeh6
U83a4pFNrSLirTbVdbW4l/ZKbwyNm5oXpGNvajzRpnv6u+HDUj6TMacW6dAmppIcI5b7tI+r1Fij
mIC1krjiRUFCWmQj5tVTFiinuOqCWTdbR7WvwK+jFP6L934ITNt1iiI29tYHO9MEvGcqQYSNJ0/B
+0jCmu3zlWdOumBqRUU71POeQZZFwGLaBczuvKCOE+x0Jl7fe7YdLpb9p5p3YjXyL5gW3CU5ZT++
9z0LETfGM46PWNcjJVXhc2RNDWf++0pcbJNd8RKqxuAfHkXXJHleHI8oil4AgiBIoAfxBlOA0WXf
I+IfI7S9s2rtguDb6QXTL4oY0aBPYCjzlGqZyHB8QV0xRmzqSWRmbmvUAEGidzDjG1nS5r5f5zEl
RAbos2sWT+03Jc4gvOtlDGrtBGn0V7SU8oVhGXwGe52PLZnGC5yb3AVBUoK4JxlYNBhJs/WyyZ/s
qxXKK1SWhhehaRMWRtNJ2qs6nk5HuWciawwivSPuWsqo46FKDfRpYo9F99febJz4tR4U/1kb5yba
/seMW+EaPmbS9Dxg9Mj+teRYgik0fsZZ4ysldweoctpHxlMv7PqVn/b5eFVyQlqFC5qHCxGBpB+N
8h32W+V8Vbt393jCKLeIL+TzaP8EvccFLwicnGrlQ77bBwLZdRCRukcmzL010zms2d9S74OoL1eF
/IR7oxcs2UR8UQ2i9d7PXQWS2V/jMbN6NJdd403HfG59AVyqtU9iib1KmdN/lHVzAJMyn68MJy+U
JDAx4+gzw9NaLynDdqaUEI1hEWTe70FS32TdUa+eFIdJgj3/Tqvz7TE7oTxK1E+sDLD/DhugfjIu
VzWPmM9YN1/5ozNvgICjgT5kW72DhJgMbON1K0g4Vd0hPwxyXu4mu6OK3H8sIccTDsPFcyjS5Unj
+9W0aqLCkTTNebgRN26K1UP7Rc804O+zCLI3y8wN4tVLfh0JdXc1GJmvXEnnje8lY62EnlIbJ6bA
jtKBnZJ9WIFc7wzEVhqMbQcRSYetfHB/CymPrR1M+AC0f5LhWC8Whqll8HUVSymom90w8RzS6f3E
+h7eB2Y3vOu+HMEkEsr+E6hWMn6Eho+hGVBUBmtAHVmald2vhLGyJwYxFNRNkGiDDU/s2Hj0vxVr
FbGZZLaY6d73E/aWoHkHh09yDl2RLVHIbMSggPM596K4eftIkCWmDVjGwRXeG/QLoGo1pWJC7Zrr
Sna+gautS810HztIeaslJLoH7Yxj59j7Iv64ityoH/YE71fbWf5y3Q2dNE4rJUKshPBlVdJEO03Q
LxFtiIJixTUSaVGrBUwQDixCQSixItgEVkhBKflWSf0Ca4GJXL+2jX9dRVslio05ne2Uf9WZsihN
6756ECA6NbAjtT5Z4V3oAmp8D61avSZFqGp0LGm0XG3YAeCRPodJh1VPvlqX5ZWBDjmd/cXgfI5u
NjaMQNDK6wjiFmEVwYGzSNTEIlWV+TDJO8jaC+7GRu80ZZMAXdHTj7+w5SJnjyG3NF18Vzs0BawS
Zq+shRioJisO/SU/9B6ikcLqG+RqzGgAbgeDwdO76CdEGv5Mj3BIwrhTGNL4w+58qmcg+zDXHlJo
GKBdqTAfr//8SYDJTNIWt7scxBSJ8isrkN0EtVDLs4vgjy00/Ilow/4NoEmyTeP4ygU8aae1KuYL
2GyAQGOB+euBF43FnAxcYAZ1aRc+V6SSd4A5PjPedXqF4CXugq7PJxBPTPPLNYCYjk++kzEWVz8C
yDy0gUKrqbAnd6EiMoZC1XgzEIm3ZVT/9XpMcPXHhoeUEkf6B5ss5CMb8YFSpoJRrALbQez4EN9u
h5WBBPFUGv5FcC8GZSKqwLIrNRKInat86et4QhA+tr3RLiEWHywZfY0MgBX7n+AhR38zKoT447PR
6MRzp+b7htL29gbVD+ie624GjkPeBScR6Pur4igYAYJ4sag3d/TaAEkF7AdfMQ+FpxNH86BWswt0
amV7u/BdBedAmjZJrHrhlnHoVnkQ/HRJuIMcZLd/j0+Codu1+7RVHJxzYtuE14oX3j+QWVrHLJ8p
okNkTMsUN3BBGMQ5vhX1qg+hZqN15HFob0MJM5Ps+FTxMbNlNrMdgeA23wFah7xlwiR07vLQjmDF
ziA4dfYcZE2vW2VfRZmIYSQWilhi7RLPZ2SCfKeo6c1kOTFA3xLIbJ289v0cLSljLb2QX3VSqnSk
fowZ8ZhUtsbpCtLJRvSz85ietxtu/TKyPL5JcGG9mKNUpCOX+RdYz+5bvpL0GXvgz2YUcXFO9Fsb
WS24ixsLmU9Gzz+QMCWpMR5zGkwJZEtbhjfmiDEt5oryqg4HnKdijVVFuQkZzE8guKs62QJpmNpt
ZPWFruHbG1/pvNO9/cvW6HovImhgLjXP8gM0yaDmZkxe7E/h4iFzh+OVfD+H+BFtKuA4/h24hMWT
/8StPcVGCjF0CYvsWiUUQCdIw1iV9klfRmJ9MRGtgyH+6yDFYGKy3DG6B4tZed3A3Hqu1XHDd615
GKSS51atAReXZMWA+A7U9gkByFr2VYB9UIJVQlvalX/p8aPqJLErdhQLrWcAenj6EsTZsARUR3vw
8LcmvtQ0L1YhgyyN8TEUBowi0yZSP3kh0R4GO8Z5N7EueGnQb0YRzVvh3y79wr+wL470rQXEeIAa
oaBdCaTNqhcv6mofn4c1CRORJzW4gPmHix+5KsAdY0eWFRmUOBkDXmsODZYeUr3Qo+BOhiRORnF4
ekcSkboz6iK/Lk6L57yzFyphJ4FHnK7ptdpcNHBLMucn1B4yFe3aN1Qqg24xi+VKxSzI9GCZOR1n
/hq9jMaIibFCGBBaVHClImOrY4X+ZNKH6cZd6csaPAR7cVxBF3ahHuEr2Be3oDVuqEzSWuQ06Q8a
ZL3xPnl0Jgb3T88poPTH6BBldSODMPOXyQhPhOg3IbBUyb0bGwAFK+Ex4uDNoZOC6vvtsm/8STEU
6aYhP1MnRzwEMnZqXb8a4Sf9CarKeeTNX1n5lQWyCHON7WxH7NH2Ma3ru+Q+q0N51v49pLrn6sD4
+o4aVnL2EByb4tVPHpqXQK9ypOoe0Dk3W28GqeeVNwMa2GVnXMIsK7eJArvYTCGcy+SPQuyCrmkH
ycKjFBcWs3UQnNb8kOODtphzdewbGHXEXPt4EW/DwClq3ZxyS86g1rQifIGLqwNq3WoMtdE95YSs
CjPZqj+jJ6L0q4Na7ibbZ+oR+i5JENDoTrnZ3YjpEjIf+xhgXehTFZ85wIO4C0o3mJek9Ymp/4yy
CdbvtReyDSfiUjAM+nlJcVMHTZ6WvAwP+j4d3/9EWLv9NfzS0zTfHDHGlbIbZbls8LXWroRPDxGN
DFTx6m7jDqF+o7gAVB7Pn3JpiwkxHuN5W8Dpxe4vq8e5mWi0aeeC7ApJMydwwyrBoPtQEfcWxmvZ
LsQYS6pIQZPfplYP+RTsh04iDUdBN/q8rgEKGE9beIcBuW23Veuvek9vDbNG9JB4NtKE6byyxpBz
Ans0EWM3rPbkJKehF2LaTbdxS0Zbt1VfY2xmqhSW67e2VRf0EVTUW4nXBRDR4EHhkJQp/Xx7Loel
3eTOMzwSDgsG1ASSxY/8lUSwy7I+T++FzNqc6YXcuZIN9KZyyBSDsp5zidE5m4zzfi2dNBOl5E/5
94XsjWve719BOtfmxvf8IPtmH6uj5L7Z1tckAkdca8XtE9/rCxqLglW+D9n0TMTjjhCXmFzVPHS0
x3+skdlS2ISCtFrhZuE6Ppwke9r5fnf9Ibv/lLV5xD8vCIwhsKroKNDplXxyCIdk6kpNRpGMbddx
++NxyI8nfJGK8T3EFXye4I7QWWlNsmxUrxXqOTqLSMA1KnpTxWQoguJJRDh8PCfAqUJXj/osTuPp
11tD/boe9jcHNLhHPnVXh045Vqp2tYnUFziV6KGgpKBPonpAEkP4CIDlfSQulNd36ce67Xpj5iQo
BqxJzZtkPz5akPVmHu+2aDvLWGdyYGauTX2ywte9FJnzEAGeCMNtAsErxR1ZCosE/8trQjklfenX
r7NF+HZerntuAFScsUvh+lPfU/PeajQ9K/q3Q3eXD1zgoAL7fIfK+FW1jB3ffQoF0MKJ4XYMCzuw
b4vZY/8pNjxTqeQBL/VCGGHVygoU6GWSHVQ29W0dcJh4X8wksE6E3BGHElY8VX8a/5f30PmvF0r6
dTTZWxQ7TxOiTrY/j3S+Op02hZA7E+bYTVTzeVZX52VW7Hbc5Y6nBthRELwbJtnuQGJU0HKtMW+d
Nngfzp7Zu4uRCWrldw+RoJL1qZUOIENmVUt/ptuszngbVf0kXH/VK+kbreh66OFNIQdFPLjJ55j3
dKpSMss6Yv08jkP+7l4vuOG8QP/D5P1AlXpeMpUBib5iOoUhP7sWGLp7m6P5X9ItvFWOqQoDmzUn
TlDG//l1ESi5u8yhxm+Kslmi0KXo1etsTsKH76eViYepvRnL/rTozj1Cgb6/m/Rd/PCwdCSsmhUS
/oFgLU6m0HU0bs3/56U2X9v4GfvJPRn7ZyHO3IneV/m8eCisrcgngKJiBMm4nYkF12SMhM9guT6S
ZQUvjQOkNEMiZ2VbjevBslFeSoD4Hbq+o1cbeDYMKv2n6pM8Sxi2+gvM44SIRfLIKkKBk/j9xOA+
Gl3jIQ/3c90llDP6vXDoZlXTrcMaoN4jjVkMQDV2gtThfdFXqaojP19zJfI+7CVFW5lKZLWIreE1
PvtpEmIfQFmUOisNl1RjQex7fvFwxcSvAbO21jn+CtWjM3bhlZvLwwvTRgUT9z8RtjZCQtL/RovN
VABL+XQkO4HiSq69ILWXrnCmbrcb5+t1SetJGzQ+FrXlf2BJM0+hnBOCZE7/khTWZp24BJ08WCe1
7NHA0tjzVma4UwLZP0hNvoSvyIbq44N0WM+uDFzoPSrAH3ceasBYxpsumZN48DSaRGMs9Zhi2tGr
7XlTeXS2LnlKqTbWTEfF8vIwSnolt9emYcbxNW5HpcmUiBvsk9pDn/s8PkWxpiXkIAi1Xe1cGrPS
dpx5sBRf+HqeCRwEl1bdgmhOKZh8TFG9kaYp+pTe5BnxFxMBj1Gt9/YEejdMzxaHohBMM8u0nmrR
snDWYY/I/KHE12bmmWv//MKt/Gz0sPMiAdaoVRf1ojZrPvmqRDylC2XqltJFhivCeIh25jssy9ks
h1NjE+RzhYGoEoUUtthF077qj+IK+gFoqs4Pbl0dhM690H2kg0kmWoLNKcaRtZCOHX+jxcmDaSRO
iAJLLlvedIRj94ZzOlSBT6pYWPmJ4V1BK/JU/a1Iv+GUwOkVLkNZfr8lmZnHZve+L11cH+P44l2M
E3iuVbjYiQEFyzU2rvSBQnAdHZvoYfb8W0vT/E6BkZdOAAgeWwrt8aZ10RDTDE1KLbmwEI2Ox+De
bMBuQ5oWR4Bt5qRoEmRhIAbTZ281LCSY7CDWJ9/i+oItDkC2AAWxlJOA2vpCQsZ3fxpY1wkx5xYh
NKa82tnz5N1K2biAuIx6QIPu3ACykk3SfdmqULg4hS8Vhfxg/DJ39ecCkcU5WQSAc2X8PSNURh/z
ZOB1DPTulYLNtSJ8SjA/XuuCMYDjJvgJ0KJ+BpJc95ROzAhYZdg/e5jlHTyYiRw6eIVkUbcQ/v70
sW1we70CK/roOgAfMrSLoK7+81mCdj5JRi895JwJ9HvUjIWZyo6OMbKf30yHflbcIgK2150HH/0f
kGbIEFYSbxZ+/5DbwnhqgJ8+wTn1JI/CkQYbty4dpPSQwkPO3w3agbPkPgSpoNIyLDbWNVMMWnss
f6kExlzCPZHbL6q0Fo5267HxgG6CE8bmTJkEVaBSLdAP7lPvdyjyNI7L+6qfn80h5MUeoOa3U0KM
/DhXdqpqAo0TIgRdcLFEWndeoYlQHsd2g7ywVDQcZA/lC6cDnKDHOxakFJ14A04nHEqlBQfBWyqN
TDuAolkt/RvRt+DmRE8jX//emIfg0uikOKqO3EQaNlO2ctnjDAH5Rx6CwSmgszB3xWo4/EbGD+4o
pJLehhqzwb+iytkjeAp6uWdpXlI0NRnc4ZwkUbboB++DZhWnv9OHK+QJpNC+tMCllfB6pyW31fD6
wxfVp8L72a3yaisx51OrV+finTE09Faw0i2dyGiICiJIfFSbbtJiz5xR7/tT6hNCLZgWH/MCB+yA
94AktfmJxCBIiZ+K3p1UTeAOM6J7SzCODnjFtZIkEWXAfOpBopyW6rpa2rD7wfi8q1Q3oEC/BeRK
1WO4o09XblzeZukicC9CaDmuJFJYN/Wt/3/9Tu3VpXpUprGSn4qAVjPuwlTVflAItELBLDbYOvYV
lllV33/V+ybvSNKIuwMy49vPjUuESEKtEsp8U+WWzooCw8evcHi1J0LveUlYV1Y3v9+Sg1+++itG
m0J+8pry/rNAwUdtb8fuzPAY7gHpOBXye+hwmFyCdtIeLYaxCDcBy2oeabO+gEmdAZV5pnpZODsn
xitN7E5RFKSkPBzHI/kCp0bcfRaedoRmnwTdUhgITDVTl4KC4AhAhdw2ilW2KK9uZe7c0fjgM5NM
EqKbtPj9ta62qLmArFHGN9FWf8U4RizrHAv9zVI2TsHwkRC3lYmlaEwOgqvxHoSKd74eAZWfykXd
X1pITv3nx8Mr1aD6ZAkqbW5/CMc3a+p/0nodBT7eVzVLNYQ9f2pv3OiAQ/MIwXa+S4HYCXNTjf3q
kbn/FRk7IWKXq/YOPg1SPVfP4o0tXpd4DeY4myDLp21Dzm7yCUTXSUIEmU2XHsxTB85bFZHsN8ho
LBpESlB3riJ5twhQIDzFkLSqYRLQKMuVc/s/gYfEzNJxPjxMdLkVDiY2h0Cl42joA9B2yidRs/04
1HIZmH3Y8U65j7MC6EFnEB4b6XQ5TQmlj9U/5DQNIKbSlW8hkR3nUQJFzhzWnkWC8gXhZOX06+uK
fbXFN4zCkU0SRJN616448Jkkg0tHN+dV3Y0jWOWO8kjW/v9OH3HgeG3WVZxm1qxZLW1Re7zC1YGv
H+GrA2F7kr4zLV6rUdCjAlXQkrvu3MVEf5fjVIqIyxVz9eTLaxYfdrrqEc8VBZJvF5X5FB5aSSC8
a8E+1DXGu+KftDmuX5vudXxDmFYvIkgtXoShwKKjVb9xYOjC+rZv4qP6zZrqrrLj/8Rda0KcGQLD
dlIeijUkGGjo17V9vZ5vnE0XQ8euYMTNIB2KO9QKqYWlzaVaGofEBc15Ns/ri0Wk3yfzpDCYqwWD
xLOMsCJba7ssVPrVaKqk5cF+9cycnGbJWmMkCZxjIyLWKLEzCIwHYUJbYkobUsOQA7oNvEhYDPXq
HcHuvDep86FZvjNezGL/rKpiI9d9+rV2w7CENpgue12lyAW7xGWZE6syrEnnThHVZla246dxZlfF
e3bj5Qzg1Jd9p6AqpeDYiQcdpCX5CfHkxyvL9TGJhtWSF0pqBj3WLuAI7CzorMKRmFunG/N68UHW
n5azjzP/doXduWYyKjNZyRqdQSfgqsYwrhGY3+vQeJmybNZ8KuhlbbiEQ7thA4g5I847MbuyTEey
cWlic5hs0xqusZjRf1i0KytdCnnudUhdaX/3IT8qTD0RrsrGyhjNQ0m0+1Cf4zxJC9ih72tMfdbc
ctYwGPnx+GjGe5iLdubiUR+ic4hzWhJMougLHnmNWPCRapTScNc3ZSmqDBuxsIDF9jR2a0L9ayef
Yk7CWNqW1IWmPNUKLZlDmUHiPp45jX2lhsOx8eb+P1W7M0VBdf9e1giaIBUhqmHVGHR4JkwkzGGX
9EFsaqHrHixp1xjQrNszjcZwY0RE2RG2W0zQ2bWSP2/E579cBRrM8UqF6KdtzHkqpnndOwLIf3Yj
rlqnUcmB2YKVM3HVE9tUpLosSx7imD+ea+tJT4q1bMdJXjsg0VlSMZPZnSx/agUc4stH8OKpwDgD
KSkxjol8/daeUVz+A8xnVwM7/oMRHBLy2L2XT9MqBaszgYQXEmeNlMOyVc86/Xf8+LAMLX6A/aiK
4fr7MGPBCkltG4gHFcr1eQxFGiyyRCv/gaiNssvZATXTWHtmQPJuHEaXNIN29anu+D0q3q1WeVyV
a+mvAIiKe7edUxFSkvsKLcdqeP30YoQFYU6NSUrLbR/3hAdqWVi00XDMBSYJ5oLjHIt8fDFkNXLi
7A8BRdl912sEUOSd0bCesf4jcnZeacNt+pnNc1ccc+ZBtgyPqKuLeoSo1PdprFUgYiE7eq5yAJpq
JBS8HgBPt14jTyN7hLzAMCjx6o3t4EW49h03nPyl1Mbh1rCpPsjYyh6aSPuTiFgigbjAuvly4O+y
qlI03HK0O0FeSJo63H/0N/6adasG3zRLs+52W75qY7SvA6pbCYRTkBlIK659WsGnlRQACwzDC4RZ
ty4Vukhd5enha22P+G12GNZep4jEx+sD61j/E4q2Nah4pxfd7b0lL0gOKhB6vVxtPz76Mq1iNqnR
Od2/eV6AZGGmPApUOFsAfFCpCY9x0fAeR3LHYYoTLXrFdoZniHCG7IgU18osxAL0U0GIUEWDeLG3
Agvl4ssdOAbO2ThZmgmwK81AaddxbuvlfSlSDlTxdC28TjU8+sAim+34N8QOuduMm1+6hpOdlpyN
TqxSKMwivgOfUonNctrlguvy/wkDHcSGnS7eZpiGl/T9NIKeNLeqST9k3ZnPSpw/1JXd0jbYOTrk
HDyw9foQwoDrlQH1fjozL0rY4jze3g1/Q3uHpRp9NJ/i/5mReROdZSf+WP6t6nfhsTGIsNIK0Dbf
ObQyXS8jFmvd4gFBGTJXMioOYG4KyomNuazhUuYYJLqbSOE0XSeeNuwtVrY1X0hraQ0Uhle4KL1H
JvLh2MIE+j8wqnexMyJXYmBQ/gsH81+ARWyWTsDVltp+BoPgQMLRSULP2A1C3LMfS8qc+2S/crVe
Uo6jnTXveAtjcnSjjciYDCSsa2lmndrlBsH0dpj1inmDZ7y8IKPkYIQpDxP/wAK+8sbowKGfWcVu
sC7PSTh4BbKXoRpGmJhj3KcnE0untXws7ULy7hkylsl9a3KHJPOgwh1JT0uC3wWWeZteaEeUU4xN
DgCp2H13aKKs7AXv0fMa/E2T2OLcx7Pq8xTod0zR1+isWFm76UQOYlzCElSBUp/QCxzuDCidrcYT
whhcrD2NtApLaQ6DKVR0RerufZLHRu2XAdUnuU5d6P/96vP+smjbWfO8G+EnP2DbV4S7aGrYGsFx
+ZcY28Dgl0Sou08xwV67Fkh+V7ONJcxhKPgvN0u4sQcDOctootZPWmpK8idVPDssmxFLMr6IWISL
ArgjBiHX7GyIkmm2u6JFIGUoTURKSUaww8RDJplNzZweEGltrwTaRj5BUBWqwFy8LhtaLGj8ztMx
W32UpkEqS4xw21lXfuoWRAloAUw5zy7Kc1w1hsl+bPbSB/jzv4c3m6YWNBwleOTneCboHlwdgstQ
dC/w73j9Qdp663rEdvM04+bquM4iQQzQxtcCgQloX2sh5NOQBZPgY9b3Tm+ZMCn79svPgBGVJY+S
bxD7IUGecczMMpAjntxQGc2mFqa0uHuMgzVpVtSjVeVpTqJcCdtkohpuw1qWnUqyrr2X99is12+o
fTI7lP4M+BQ0CxSdxlFnIlNdKTFf5A4pzumw+Q2wqucGziznjIrHtz4b4WPNO7Yj01lXu9SO1KMk
p42VJfWjxcaeAkP297i0+F5NRO9E4iLWQWAzIeF/fWu/ZrtVHAwgske+prv0HhqG9CPJFsSqGa4s
NdhWy7zRPwOFvP9CH8KG9/HZ+YU1ks63HdDCSIXG8ow/erMe/xc/7NCvxRZXfJK9t2SsCX1fEIZS
p6BSvw35SVEgmf+sLobDvOVjNn0HLr2EnwTIjeuSkf8CzWobfrX+5NSmoZB5wXpVlU+3vgr26WfY
/bCD8uAKGHD4ELwoHJeJbCoLr/CgMdefX8Bu4cl/TCUBIydrupMUhqAdz9sZ9en2k4sT9jq+AVHv
YvuC0jiwP7qa81+VAZM6ELG02WXQPzVDD2iAzpoAgkS8uHA2j+9TjQrZoOq/j7wGEjZR1OIOI5vY
lM3gV7rmgAighjLiPR6yeEmDX+uVhiHO/FZSZQa9Qt9vO4aH0jJAEwj7cIKCl2JdP1ivjdNeHGNJ
CQlcsqWK1j5smRTslclBv01rtwiSTqSvKcjwJTQhX7OlUrz4I+c0NYo3iA3GJcsvvDv8tapSUxAp
lS7IAfek1XlAemZBk2OJwW27JPEdFZmRCZbxEUghLfhnDKPhRLmcuMDcjC+7262yPytyKS2dYVKs
FYPgPWjgvxL0CXvVaZBeBlX5YjogFOfGzLo9X7u+ll8rzGxvf3+pAS/u6W3Vu8jjE9FBNU6h3tAd
41S8klOlP/uslSrOrBC7O3oFoacoumM4mwpL1DUHzkky+I1SNCpWbGp3btKJJP7Gmij0kuJxAlST
turHcvzu/9NGo1U/Dj54obof9XpPLu2gzxp6N7/PYfehpwCBRiHavtdLH5Vmj7FHZcQ2qiQagx9v
Yjumqk6XfSPFYDDtQEOzUhP/ClVpPGg9it/nko1qaU6yQ9qXJ7YnSLAEgyD81In2l7vM3yQzHw0V
vzT7SKHw7kDS0yIVcZwAU8FKy8FIfo+motPeowoLeqtjF2qrzX5b+sisPJqXGD0eL0dfRMxbsxXN
lSZY842oG+UdQ1YQpMXwAsn5mNFMebIEIPB27T/pYEJ7GifPecKDqu6Vjt2UW5nhn/x+JHBGItzB
QLbp1wAW3IIZtW74RHW54fP1yEUXR0Y/XdtLeVW4vFdTPCUq8MSEHugzJNhlWjirWKlbVXzWSPJL
gOoo6gZPJ2sK47sVOc6yUjxtfKevG8/XFb3XRVy/Xyh9jJOuqcbdv7XgiGweRaaGE81JVrrJv+RO
wSpUDI1I5yt0AWteX7tpGJYudhM5pFFZsmFJay43mKFcRiYGeZjlol9BWk13+Y79mWg1vETVqrNk
R8MVBb7LaO3k5pA+6nMGHxa6eDEBQay8xw0e8CmYd1e7aMIPMxJKQPBgSzY5WuniiHL2PPj2biMf
Ol+/6Qct0BWnau6ubCBUnIL9c9voyVTszDXUooG2wOYc1+lwy9uvsu07r8nwo1gjn9SQp2Un+qzK
pzfWd1sEEdO68SM+5y7F/avvFb0JAiJ9bm4UlX2+G//HWPmZas05Cj5e90ROjnaDgRvD9uwBDom4
wvOfzQR2uQA0doJeqlVZtmJ/gfHp9vFYIvxLiQSvqCTxNMPOJtTwjJEv0+Vl6C0wun2Y9/zXGuto
MaiBLK/OoNEuFXv1SkgH/RtBzNsimgLrdTTyrSf5VGgB2wwr6YPqUkCskfBDMoGCI4rYWl01cmEc
Hg3+0TxMAwxZLyli1ARcgqSe1tYmcz4kL89UzYGK5ArbGtTdsRGv0JFdvaukruLAROI8nN1Kpwkn
/iimLVKC+jYmO7DuwrftuZ6o2Ga+KLqORgr3V89qohLo3ngCmn9kDfVsiLuyRm7TFgJMZRsE4FUl
iQqJQEJJ/wxoDjaVVeu44kpMmYHLzASUAeXYlELdpys16nAhFrlP6Wo5Aa0s7CxVH6fxGX7zW5lW
LX1TFZ7zmaCaIbqZHPqfnrzI/JOEDgjYrQwlFyX8w4Ni7Iowv6Kjejwkv2RunVRubtgbE+eO07Gy
GFZe/oOoNZ7Ik2BbolNSSK9dmmTOnEIdtk4n2YNEluKoLfYH+imkFx7sGh8BXmqyzEoni9+1ygHx
CM5MOY0exPKIB05pSJb6FoG1DlurShZgoNvKL7qmHs/wFEjNyEhF01m9IHf6JZvuaiMilqVmX64n
xA4HcTMTWoacMyJHw6uKPLg7s9aTo5ltBCFjcEDhfgp4Sm67TXlAjmZT6QGCV0tL82bBkdjyQ4Rc
L3zLfFT+O0FCFPJnvsrl2XHa7RvfuywjfPWUjIcEYpa0nc1xsbTQd1/qkH9Dw0egO9qZuu/ZxRhv
N71nTygg1g5zCdmS0WYefDGtr/lMmN6eFaYeE/lKtolHcBN64an7UqppiVZdDCOMp5tFkOJfLSPC
oTpJWeH68LZ7M/EsKpP9Im9dBRjCaJVoclO72DdoHjjfCGXTlegn7x5V45jra4Cj8sikIBzH+6rI
vvfJl2Y6kI3h2w51TFzLLy5Jdhw/geT21elEFhpfjMaXz8CVPnnmzdguKTI4/o8oVppLRxrhPBxC
mBV1YXCL50GIhlnlkTGtKCpY+mlZArul3qcsWrcgk+iWUy4QYgRZc+a0feqHC898rnwU8+06Ei8l
s6XIAHygm7fj9BeEa76gYRtxfRJ+55RUg/VXkDg940u5acwPgPxZewGozQvxM279NEtP0s2dHWe0
g6MrSd3j86gUErTjGf81mpsM5XC+gjrWpr0vDwTjyVyLzsA43+yHuMUBoyUf0r35Z7Kl8zZoqiRP
ZhcKSGcw+7JFXDja6/8Lv2AlVLgNLU3lv6+AEVv/2T/UDNSRsTvhexnjvVfncT37cXvjr8Hr/hdx
X/7yCkWtyVPoQiFJCFzwteiuB6j65dx810zeKYr2egAMkgjIG0c6dSP6UVYCncvMn9dhlXFjONC9
BlM71runzS1WtTlMU5GFzrdvhNHudcISC5OC9lmdJNVWsEwOYQgxdWMKpqN5pVL5ueFFpT26i/OD
Rb9hPwPth0ISO05Uve2wOauA+8oou4ys8gR7Z2htwn4w/NYpacSM+yU0pxbvj6DDmtEkTPKeoS0M
1vWeQPhyuvt9wc5ykLKTL666Vzkzk9G0E0G0Ejkh2i+QOGcCoCuRaqPBa7sPbLCUlUavAiDHZSl+
mmY5fmXiSZc4w80QooWtdsvIwdu0LhWA7WTiot8bKjibagtc2ngYb6Nt4ho/alvoN3GnNVDSAxoM
O3CGcByEbEg5YQKEDO5Hk0zIWdhFoMbX8BhwWkT3sDxwhe3j2No4IjRKc1UNBG3xNlYGqIc3dxlo
SEPZBscT3VbZblC+vEGA2JDH5b6Fh+dPY6ndnnInqyz8Zt4I2EH8pYdZb6npYrPrsAZcicfkyNeF
fbtcy6OdY7+Lq9QBQeOCTyxOgXsnxpySNTSOi5+kEsPLYMeAunxe4m1Rte25z+/AyCJns3MfGSZH
GFgAZnoatYk9+2qSJr6dIE/kozqz+wxuXogywmBtVKjQOPqSueusZfBFvczk94AyYOJbNs9S4cGB
rd45Uifu7e7bKj4sjm8Qr9UQEtpJKUGsly70VeK8V9XepZZkfSv9IjaVruouBfUj5xptOXyiRT5s
gAr9VLK1yRurYGBneSuCf9rcdTcnC51N+xQohay6hg0OVQPkBLoTfajyr7btlB32ZpFv0jPj13xx
h65PUYBBJk74GMAJXotY068upyQq38qf4YFR2NVI8iqlI8RmOlQ4wNazvRTlFxP+odahOiIsJKS3
HYV3LLrdUndevCXQgWP05AEutMiF57oTVTKaZB2w1FYsJ36UJmPU9AlX9xBTJARPTLrFPNOefXg7
H+vuVeeNbPvRwSdQfTSsJUFKch0BXYeK0yVZ/EEZ12PxHs8u4+uh7MNcMPLXVgQh5sCNQu3p5kO/
MrLMl1oxBa0w9rBJgguI3OFBAapsvqgezfGhe+zuwVwadIHXiJLzuJBDp0ZRXQ5RfPKywXwp3BTk
3zutl7Px3Td/8ISNC7QAuiZ+VLxghtd25iKTJzEzqmkGVy+Ud7sy5gkoGLruMSdrs7Tfoee1yZZX
I13xgVUP2PsP012Z/XoYMrz+p0AiQTb6tF1UrFBCv20SHjCsFwQtVysY1a1lP7aK6SyhQHUk/kon
FzlB8Y3TMdAmIZ15CtOl4F1AB5ItkmbOrtiP5yh9a3HQV9jSvr7uaqLhu+Dn3HlluGrrpgXCMv3E
Lr4dATY2VZvfTcMzBtqBDtn6Q3011StjD+UZOonOqw/MVPvyKNzemZi8qg59JqWaH4gk9tHD08cl
+y6AjEq/xDjAX1DGwlMRTnbrZSz3UfdE74J6AK5QJykj/8qZH8UwPl6r9qmZbkvktKIrcNsInnzG
dpyVIIP6zhkWxRKZ5rrQWrfHzp4d4hY+5/+SQID8kKCWNnPtBH2WSkvOLTNrO4pbXaDdISTkSKV9
vpKAB9sf77H/k3/EDR++aaR38zqmnEY4F3B8DI8snDZ1B81ZSdQlo0m5zwYfASkFtMM7UH8AVNmQ
rwdkWcVg8rOALD1O9sR/jWrBgnfJ8q5o8qXk34XGPVGsSeBQIj4huPuBUrZkqyhtaO8hAEAsUGEX
HuvCEkLaGsak6bikoN5jIp7gvbLuP6581jkaZIr7vCaf5qikBvo5V1ul3Dnholq6cH3jbEfyFlvz
berZVsBSGjw7pm1Mq9PmjID7ze++xAQD0geJDw1YOvlAPYOxY+5qempBUCkunjiwYpsfwSeX2CCO
O8x2KXODmKbRq+RK4FTb1CH5iWvTp6YbYxv0J14qvyz/kJ7EFcU6HctcseHFOLmh0LbZfXYTBcbt
kMZkoR1ejdzr+dhnjiOrmiXdB+QapS+VJuSB7XlB6/1aE1bfu2ubDt/x8WKDyRta9UJ4Tsi7wFsV
9oDdAMRoCAfT84uGAGAu+NCTfCviF6R8T3F1Afrym20dH2hUKz8d+54hoZxcHNo2yBc/PGBLtIwB
Z5y9omsi5mEBldX5uGWAOZnWkuOJ7lmoXZ7TTCltY6nGqdX9O6ySRJtrx5ewxywawWiQZmmJZiAV
o+IIIG23mAAyY9E0S18Lmzaar7TzQWQ1aGwsZlXVTm9/5EV2XWKYZttjJyx0AztbUpYR4Vwb3glW
ifjsMG2dT5Y6efMJaoNvbuLtIqwrwVKuwLKUMUXGv5tU+GUgWESOaC37MCHhMDoty7QiyezQLmLQ
MtLsvezzMQd4ervuQ+tGnUIuzLrnbLooVAwyCQFPM2z4x43QK+0knjCSgHEwmLGchmQVqO9okmoW
eTpDjaXIEpHzsyPtULdUjL40zo0ogQPT4k9ViMJ9bz/9VRgeLuKUVaIPf03rV7CjwOm8R9sWKQRn
Kx6qrjNj1wh3aeQo3YZunmpuHi9e+wKhfPPAtoR8Ej7/GJSdvnVmpXkOj4od26CE0I+oLmSbmhZq
9wYLedKzPyFILEetb0Eryn/KOK1HE+ak64tHPnfCMnIcbmaouBMP2Va+MiT41zDwukoTMZjoriw4
rPOy4iPVyK6eY5AZALQ7M2bHPsFQp/lE5gj5yHwzhOEPhCScJGYkVlGbIgNcO+nmM6c5p9w7UGuH
U2XWsMEkjUkHUPAATfVU2AlvZ3Hm12H+KvleD47LMgu6DK8foAGVyEBxBG+9zROcf6DtKJm1ZpHG
s4PYhMLuOv/rz2fQiLN5mWBM2cehEh/BNs3aABC80zS5roWpgYkLx+rl+svGL7YK+zLzxPy96acC
+lZjJNqDyQk+83ohgAeOk/Zgr3t+zb5FfPisaBRygZH0vS+flpF67W7BD5fVmZNIN5Mswi90XvMi
vHZllM0GITWA1Bse58LNPgMFMGjVxxAUb4Gv2PhbK+mlY7G9ZXWrcL9sLCrrX0OiJmc2bLZqbUBd
lLXKMpitMoaCkqlvde8JroOHS40GJKzRNm/mqB3W9vko4j+YEANI35Cx0Spd4Nb1A0MS2lLdS3DL
JjXDTN3cYEREwjaaTm7BT3S7iRwtOQLQcLO6vYsLHUkaPMwKVSilq4pdHPRGAF2SL3/sAcAtvSg8
U7c28MjvTDXDJoNuJ1LVl2EyMU5jsnFRYnLBWir72TPNc4VGtFwjbM2PnMnjSAY+XAzYz0VoQS5q
jqrK6NuJr7zWCwaDCf0wQLFJrOj4HI2sh+AvdCqPxg/bD4Nc9jytxF7LmXIDMTZd7sFVs8DhA5tt
37wNeT4t8khud5aT5opR5KFUPuTlnju1+SBxT1hCLmSV1zgrPlUfjLcHu+eKuGfS6DcmhrtbJM8e
RKueGSoAN633rZvt4OgiZ1XZ8fdQI8q3uY/bDIaGTx0rpr4ahquWx9x3usJnGs0i1OYmlB4r09YZ
FyK6K2AREhVHFGJY+LSd/ALhJSXCapAP75L5bzu6MVXjFjQjIFgJdXvLTk7zuF3gk21XFnQSXCr3
rBzYKdMd7qmJXxt+LN+F25HWvS+slmxHZaWmCTAttSduI2bTPwb3PqGHR5jo8WjuR9Ye6SGhjPLJ
AQ/JIA83f0GgN5pYG4M7p4iCjGYXS8cYPmnfJ7GgrxFT5n6AQ+yXSlJRUajBp98YOMt7FhRPPnOY
K8kmJtUmJDV5Kuj37Ny2L2lIM8qJKT0azGHeivPKm/BWIafonuTkwX5ksifRpxOgBjG9iWAnjyBG
F1mUU35mYqgIIL4N3zvMIbSYuDPimiEGOKy2XMJRB2yeJXkLiDIT5qdwv7wbQ42nPggWUBb5GjaA
00iQs33NVuVqd+j0LuFMl15VRii3adNGj3Tu25Co6dr266nf7eny7Zx8SSeuuy1lk9Ai4cMZtmrO
zBtJpVb0BaQj7PiGQIcKh8RSbmqEWo5GiHu0i34wPcFZkz/n449YU1ZlI9vil2i1Kse4UrB+HjYW
w5EVKFnnfiwUzTCRRl0ephmaBWl9nxT6eprCscVtE8jXIq8yjD4h3ZoCIaadDTcKWQ5dE8GTHNYD
oF/kgzAqOkw+AOJoCI7fSV7JNebhcaoZrGRQFXHkvb/WgGmPhPOCF4aIw+nwb3wCz/9Ux4FaMyr9
HyC/aSC96j0FJdg71BogAp2zeJS4/65wZZOet9g0Y2q8Q8UGj9LFjy+yuPY0k7gAzmLiEunGV8VU
zwxKoTBs/BRtckeeuj3Fg7KIGU8v6pKYGfD1njiptX9ngWSpMG7C5D1WsVQcj0odl50ZkrOY6+RW
Sa4ckNDe2YwWxM/s3N/WOLxuB5H7tk1AwPdS+LZ3nctyZjxKNeKddNlQXQ77n0WriGgDam6HaNGc
ogk0ThvZLAyj01BKxRxBuQg+HV1O1DmwzhKsARgYJ9aDvdLN3bswe5tod7NacYe1pPt4I0KStzoy
rrC9Efb3xi3PHQ1uU5Fcu81gmOc23pF94/iA6X4nLuhYrqMUeg8BawSut7jjPhIFl+4ul5w4V2ii
P8qD+75uz3Am0le0isbT2F1Eg47V6hkuzWQ3g7hQPjl5p9ZPpFLePAFgXp5g+Jg1r8pioGtOTjbf
JVXlfofpvcKziHvJ5NPUs2nux0lODGyJyZWIxgbjmr2qISFfbLeouFgt7KhS0eFsucrtdaSfaknm
6yhYjigGx4frrP3fHLudBG542YgVEFs7CWfGPy5nr6Gfn4sCaON4nBBDBw7Etu7RpSsf0yDj0Z61
LoR3B2XEHdT3LYz+lMCpRdWi+9TxRbn/zpISwNLPiCrx09biSbCKHVDgY9a8Zx6SEdg7hjmtwtJF
kfKiazKPAAT6kwb9KoN18DmBLOSuBOih2hIqx68xhzg1EB9pstMlqHE9jTJY5mAZ7CekZj2sog9Q
A/hk9BOR0wx6vgC24bSkGg+CCOA13gViREdUZ9VEFUpZ4N0+WKuYGPlq4Zk5G3BCNpbUtJ1B9I4k
qBEBoqyrWpvEQIHy9OclBurUv0g3eNNJ8TZsYVZS6LmztdAmryeaIQ6RM9TCTX6mTQSV2vo3RnYs
1wkiU3vxtH3Q/U18cyqL5nLNOjmAzR73MKXB7TmdL20/yEkHY9XzxlWtxG8Bqqyr7UCPKEM/2SO8
EpVYvjRhtohBbKMKqayh2uv9v/C+22YyhqdLhAs4zyRHLQTN0juLSIFdL27vHFUVPAPc9vQlLyx7
RPLJsdqX5qB9qzw/RoDeYqMYaN/7mE/XLZhaQL6l/bkVKBGN1+9g7XbjS04KicWhMleYzo2ePnpm
wwQj+MCXwXaR7UE59DzELlPnfcDdMjvp677PY33Xr90FnE5IAXFLymRuwr77k/OF39OBvsqtMcdc
VryUq1UmW+7fqLaVf9M4/F0Ju+FT5C0B08bNkE1WxxqchQy9R2y+8JOzc5WJQtd5icWNEBtV8A5q
vKlLnigWe+lBRNGDb69hQdOzDhWw8W1sJ5KhBAdEfbKB0eMeq0aZ7TC3lhR50wAVhEi/bD7WDnVq
GAoTBenqdtkLtlneox8Cl02UM672nFjJv4lrnmGc4LowvnHQVUFHL3veegX0JvPtlw6YLmiVOxBw
Y4IcnZOzY3YqI+8vf8hOdsjkYWIum2iev8+G8/vsyYGyLkaiHCZAivtp/JCNxy7SYW5XVwgO4HuP
DLShQHuZx9IApFdw+DI/HQiDBYV+UMVXax1tIw+jkxKsIrWHFa8ToigwKoVaHE4kTtrIxx9kepWo
7qAkoER4xfWhONCRda/WXEeI3+bCMdep9Zw7EHtay6ighzsmImf2a2rr/luf2RAP602bZbzdjZkC
/LP1F6+pbeFpiw+BabgR/R5ozp+60yMDHqhxiMjWXcrVMRAZHpXApbyDHfxEHXgWapi9OUvmfYnl
f/3G+YguMgYaQ4r4BRxBZnNIicxXyHVf+MwA0OVPpcJcH+b/F9wKWMyAlv82RWKeEdiG+tPcPWKh
uVv3TJc6USSlZDSlK574dAgNfUqvshok9qr91kN0lhj511CueNF3qATdOnfzApF5Uh3nP3U5V5eH
L4EdQmgAC1VFAhwaz+Esv/Aqga6sYAgcZX3pIb1H2hM+sf7sXxRquRePP0Hs2GL/371y4jL3AaMH
BZAfyISzOd30ffQd49RXP/CZiUfyFq2a/DXLwqsFwgSrenrCyvlTmUTJjgd+/KiI2nKmpz1qbkQE
F5fX7bceVGj/SmTzK2w/8hKmrBURvfMCKD2+sOdNb9JDmfANiIb4K8Q2LQuM27zXMjSAFhlVabM/
JXzqAmp5Ej7p7HDy7bnpbJ5BVxHwEijRT4LGgC74n+ixFJ74AuVtI5RMbzor7KV6DOwIovCWnBGK
kgYgmnyQA5P0m5vlyXRFztO2gWXZIuzCrKS6XTrxYOfiijXFocXaMgatZYh/a7Dby6XQ0br4sirO
NtwhE5wJffeARgfm3xpaOR8AjUiabfeYBdDWLHW5SXAoJWLJxrtNDRgWlg3oPJyXUp5y6rZ+Bf0T
ovrYVQ5VDwqMLUU77Qi2HlY4i0yHHzIGBC++0tIxfy4NDnEoXIy9BgmWrrOXrukG5owRCDwijBJW
mjdtCeZTOF34UuBVLE5e+y5ifK0SsygZ3Cojir5pWa7OlrFN/4hJAkn9h/3PuNcNzFTQvDBm0MpM
WVW4ZQvM2Fiay7JVKi8voMaAdIX6H66/YI7nEvbU46ex5TZ2MMYtVWjpAq1psKbmrOb0xOjFyrp0
HVYubRGrfUbDhouAbeuNLcmvIwUXyxbLjIilvRSZ1ZoIIz9toUe+Nql2Do+ILRe3e9LBZtFMnusY
XradLoes1R4qLfLrL/VOde/uw32hGfQMf9xUyCGeG/th00lSLo2iH6U7XdmDAEMZp5zL9k74PoAi
JyBXBMjGkRuy5sPyPmo4JRc+tP7clsK6tmcI9fBlULKCau/hdANzfG35+X7b3xV7F98afHSQAVxu
DLy2eDmiZxc3iq3UxiA83WdOl8zERoMz6WYA0yjljyA59IBGduUuB3WYctlptJZjfT5ryoVlEQhg
P/peCCnsF/7+4Gn46hEAvvpSz59e7onH7g1dZQztUUvq3L7KkJ6cOjzZnp/5fO1yzBlgAPR9a20s
gSXGldJnT6kb+zNqpwSTgWpGQCdnAoKj51efcE6vlxFvE470AjYIv4SOycsW9Gx4CaI+pkIUz3GH
gpynB2zXoz5mKVxrge70/DkFD+C+bh9T9+qZgn5pg6VftLJU2pK2gCKzvp6sGDcpA7Aws4g90zyY
1KhcuKcTIso9u9zHigah5D6iIGOyH3Wsr8rUZN+ufYh91+3e9EWvgueN8Yd5RpnlWIDi+4pdh0mB
4ZHAMGNu0lZr0zQF8wedjKdQk+0LsH1v3txhCcYhvgmzQ+/S4cXj0hN2CicfZKUfBzyPN8pbAZME
jdDrFWQCrYNi5eMpqAXRzPxm7BpVqyD5lZKuuBBfIuAKjnGuJrfStY0t40ul/ozj8uhzaq3IK+q0
QXCHtkMs7HmTAC4l+Sp0Nnek8f4VFfIbfQ5XIzljtCuvlRZN9ertwQ1Z9FEFXAvvNqor9jdBmS7u
toHvPFGXSkYeSSMgxZG6UC9BvHYXFSggGVg1FgofQ17btI/MaaiWyLw6XmHwIKgT5T73jvBB9vs7
q1lE7kkM1M4riD0lSExku4L53iLqP142jf2Gc2vli9sCIZZvIn/ukzbxkiRBxKqWXKctTu7Gb8GS
Bx1aL/OdRnFvWqduSfi6K8Njfs1MSMUgSfDbMHQ4qH5Ng53+53Wsj9E4LxMYnspLn3qHk45vqM8o
aQRN8W9mXZA3UYjXhVfBDNpdYh96hxrvhd41Te+T8LqR7/WlEukypHfhYRL6zQVTdrstiw0NZgKe
h6hNkiA3P91nvcTDitSvJAfiCCxwqynUaq4a2RiWtnshNskz3wBt8EoIQ0KOAIir5P728iYcwBqK
ae9d/ORA+62lhIGL0EeRxhOqJ3MTdyxDjrUUuy9YOc2KiWlo17MY/Juf8zfmIk54q2v2GHHJRY7Q
OTFfjCCMx0+8RLWmWU5JfafhbjSanT3ZqD5Ququqjm4ZhekDfXEEqH2u9SFrL0ROT2oeTuPBXuiP
uYF3bzJHIkqyhDH7Dpy2z0U62BGa3Wyq1lT2oqSX+vJzCt4eINtNMcD47zxYyfryY6J72lYU03t7
4oTzSJ0pLbSKCDlZ2U5K/QM0rw1lTODq9/02w4MIZkeoprWpI4vvSurb1J7lIx6i9Cq09kS8EzOp
6gCZlVbbgtOnU6QuvPxmou7x082DHLvDnau/R2IKC012XaV6MJjgULygw0La521lUYrH13NBeY9N
KP94gMosURZ5JqZ0YNIclBHNX1NrU8g/b5fshse6XM2HWAtCAfYwBXhWe+w4R9W2Qw+dgwxS755W
lowY0RlSn9dH0TVuOV8mbvJx8pWfAGZWc1PHassGZjXgMNb6H9D+hpXxddVGy2zxA78T+qBVpilq
vTsRq8Qw9h6qNC7o4Jl0qaY9OQ2wispe74CnkhHdnUqENk9l/ISjbpXmHD8HF8YuDrnuMG/A6j4y
DIi9AxkiMQwTPq11f1SbiBtKJdeBvvw3DZ4JTRr+G5CJEmkBreed0Q5QtxXn7Zp5kQiupkpw9dqg
H2llXvPPHKf/s/a0GgOSttg75JkmO/wDgVzBN7w2B+iF6wI6F96x+NjFttY4seDsK9+EfFcjEUNE
kN6FKacoe3IC47ts/U3O7XWgVEMyenJ7ni7iJpi2RIpjB0/Xjr5hX8L4lZmaxQk2GEVKjiTR1308
ULtdAyxPn8zSL+ILtznl4nuLTK9iC5ZfWVPfH6pLAiN08gAORAFa2TbiHUWCky8z8YGRQ6WAM5ST
STc6I6LPIyAWaUbzEkKqwAdXcVsYigJWY13wz53PIvopkbvWmhowAFRV8ErLpHdMrKxg0jjmCRMc
M9X89QqC3uBCO2XieEvt51VGioLklYxpDwSw/g0tVhowJ4QcmXHhlFLBOuvzbGxvUN1ELm9Nyfxc
JFEk/OU4jYIaxWA+IptmjWXP4ikksQ6X/uYdmg8SaKUwqls46lPOVyg1L2shdQaTKZm5aibLLxsr
hLnDhYuPCU1cDwQxgyKmnFIzbkXK2cvZl1IxFtOIIcXEsN4JsfkeXD9P3m+LY/3t7o2JAxBuAvoA
Q3wyoP5soJM8rg7IG0vEXJI3PY26neWpRucrmv61i6Ok1R8tvGZ7gLjKujguGx2FZPjEEbLUTwhl
+RGHcwWWG1/gyYseoxdK173n8r8NvSCUACor16rVXmG1mM/+nvdHo57i/3ir6i9tehJIrrp0cYlY
9fug2U4R5CguQSiPxzT26yoQ44UwrQaOdRGEumFLham83Xh3S50emxKtmhggxezSWJXAEeXrouhb
kTbJu/Wbn/pqC7VZMoKYZRseejraDvOlxQiWDiMy07Wyh/1JNWAMrLc8sth6Bytrn1alITnnf4R8
QeVMiAaVVp0AObeIQS6mNKUv98QoilGw0m1KHCoqy33yN9fy/1sOKSIOC6TQVGs1yO1HrGrXX//m
stpctQKvzOiTinaMkJ8cq1GddjGKncbe/PbvXm6DUt9E7wkJhuGxHeodUa1rog1gLbuHJ01LFprj
QREpfDbqo4uhfv8mc0wGS2Usm7bjQKZJUKGrPm78RP/KprXjG87TmT3PfeLHUTGSmu4KVjwH//9U
7MYxnEdZNJlQnzTM5KmxKWXrl1xejzn35P2nIcnCX1Y+NQwzY3zXUiVauEfbqsuyZGyGFn9kr7nW
KBck58XaEiR499+wPy44Op26dV8r2meEpjVyb+DrvpqL8nJv4yWj9EyVC4+E1fM+R+b1yr3iha9d
pXKc917J/bS6hIvlnueQUR6OSl0uEE+1Nt5LqXYACfO+m46ywPBLwAFhYutkUx4OrTgR6KAzLYzF
5Z4fmvMzSyRtsKl5nq6SlYKIPhAEXXWUdYn3p678AgpUPPw5ohLMFBUiRdK+zeRmFX0tldFgAdOe
aUsz3vHtrfb+m5HHNVvLGxz7TH3j/u1FfNdVpQNgqMWyIBo6msuwhcCFXoapuXPw94pCqFC+8TOF
hYDwLbOIrFkW9yqFEpdtfM3esbNZoSXHzNxvOJQAreRSXmRl31X66E5DUEUBDr5qlcFQT1uLlotW
f7AYbUePzVr87vzc439Rkk3ZvIndlbfGXdXtzeSLHshDm7DOGqTzgithQ70aDAhvX7939Ty2dXwi
nFMF6vXyJfbPEjWDQwNSNZ4931SPKxi5nsVRKJIDt+8gsSfMzb+h9xYuyKYjeWFcDeYqtOiQZh+2
k/4HTuP+2pj/K5OHwC6z+pjTvZwKG691Xjs1ttkWA9g5fdzHJg+CoJpra9svKdH7OV6/1NJ0lg+A
ludR80dz0ZI11BxpBsOWuRlRHhDuB7UYIpkinPdV/n/3IcbcB39clFPRS0iJFSftpDZOy7Xj2kNp
7lPf+BRAHsx64tq8MYWo7Xh+XE66u9szUYv9VciTDIw4wPnkFn1YKlssxxGgM28QGRlmGPHw79gX
YZF00WiIMECF4bk2shRu/jyCAJsdPEJJE559yEpYawDyMQ34tl+2obTtCEDbKJa2NfXq21Ke+wIn
w4/S23KzNOSComUghJOX9YIfPmXZrTuifTcOsK5y73O9dJPowpgNdMSZOTmBNbq74b1WTcNoBEI7
JgCA7Gpg9FHaB42ULeAXPDmF0IT0j0oFkIwZ9SAlSI1AQniXqvGyIZf6q8iCVR9O1inFKPukATNy
LX8MCWTYHorRR3Auz5ccortQld7Rq3ERbHQTshuzgLjeB9HXzg9v4ueJQWF2GLMYMIsZl5tBL5kD
FM1dAMC6um7dtwqHQl3/0wjdymB7RKViHae+H0CIfwmM4D0jRuWKqnsgnF2FBF6JcA77TU233voQ
gXm7hfxK0/LvPGw8HoyRCvkai+d+YUrIZebfNfsxElfgrs/co73YKq/ksiOeKeaUENHWx4uDVRLb
y2eNbH+YLmSAtJiaJlunu3yuCAtEheuSZc6BPW53YeGM1L79e49z46DwvqIhFWD7bcrMKTEGGtsu
43T2dHSGbicFATNsgSDLqgaF3pFdIl3CDu+u4Mz8o/y54K0PeV2VmOXko5b6Elej+LUgucPTSlFi
5nk40tR9MGkZM07zHAB82wqluedxe3U0qTv2h0A2iWiJ4L2rzxM4yW+Kyhr5ZOcONr6tEOGj7KbP
MRtEWvBx4Mo2PAMnK4YjzLGqHNN5XdFQqSeHelFUsxfrm3tLkW8uIK54y6TvDuwgseI0L9ses4mr
GbmVLaNDISE9nj/3wh9HW2o9BQzdei9SXJSYWnQIT3kp89eA6dzfzAyXqzPzorWz5DCu/dU87sD9
6AKYP7eMiRiq6K7NxkOY1M/Sm6UlM0wCyj1uKErSjvE9cSsfEKvsrry7xyclz75sM/LPV6N6otJN
3sB+pt3I7yL86WD/7h10lTzLHbfa6cvGkPHDjXodm9ZhCHGvy9dhQkPNBdmAWAdXtr5JOhYfjN6W
IrYE/qyTOkWgyEAZ9mpvXAYHRPyL3CTYqEDG6jMdubmQxbvlJWi+a/rsRodGB+OIh334bC+1J2l5
2OYqi2N2PJTacGKHjfmwSYkQ5U2kx2llINIhCBotfUx5duNWxsXdStqxpy9rG6BXWhbaMfI6/FFX
A3oQqocxex0o8PzSUsq2KUz3hKG0b3i7tfdkd5KDvdD6FsxxK3v0a8Oq9t+KmtIH3swUNfs7u/k7
zUisoYA1F6T6ucG3oyAidqxhPeeYtkz5kZH0WVqrVLQYQnC+pOaAZRFIG6DK5z7/2Z/+gE8hS1ew
eEqMWIDhxX4Pe5dKNFFBf0Z2GR7nJCFLYRONnLwbrhnjjfG+VYdaQLG7qBQbue7hqCmTOdZ30rdF
boq7IvxlXx11kOuBpvP67ZOGTDTTE11X1iqcbg0UM7mu0ZC4PmfqD1UUA0c+Ao/m1HhhavbqoB2n
5qSw7uuTZ3aDXJbhi5I7rbsQsQiG7HLMgtLfwoIHWj2igJjQwePCseFcNLZvrBGyd/2as5U5R9lO
b5fM+4EOLU4bROpiQ3bUQavK19HHiVQ9sXeR0La/3UMnGCf6ar1V+HY5Ink8R+8JfkQ6+vTEDLJd
lRYlcAgUgeB1c9EaRD/udonvr4wS77Da2lQuPAa9ADnWNx2PRbvfW1aPLR0tOcuZAA5eO4gpzLvi
E25RW74vTBh1TELhHXibbBX0kyFvQ5wu47T2tPaY5hDMo3oZO0PU51FzMDdh5ry/lyYmc9YBD0FX
wZFunsmTL+Ed5KarWs3ByFQVxdF8gpunrG7F7EaCYpQ22XHhOBANpxeKOpPsnQqzu+QODWx+gyUS
/lR2ydQLQoMhPYt7NjUF4I+CEcDTjpBv1xVS9TOYr1sAWNY1ziWgJ4FJ7ut+xJGib2zO6TwYgR5N
D/iPtYoIO53uK2638uKi/CT3jDFvcOvQUET1JRlhu+iu87EuDLscR9T2jCVvBh+Dbhff4mMJawlV
ui10wiHNUhx/+ztL0WOcV9IW3GLhRz0oR5/nmZw5tfBlUa5OVlKYOCzLAToQrNks9HwwlobX5Xks
4IBQdHDr5GEwMYqSXQn9fjDBSfE/N5qu+LwOqkL8CuhP9gveaiFvz1mt+YfslNgIWzeyoM6T7G2X
Z+YgmrhK2LMsQpxDIL9vBhBFvUlFtOzM2J/1zFNeD3Lc1UjgaULmeXIIhhx+8MsDEH2OpqOGpbwJ
gDOneRyBJb2vDWK95tt5MpmBKbu4gI1RHeyR8HVrh0CAocU1plS7kKaJagsWU3M3n1sJ9NxADpvp
kp+7IfNdAPJtagozn6Vfic9jmj9RxqoItb/fZP54IVoNVw+RW0RInzIolnQgXveklnIhQMsUUv1j
WlOz+eNKhHb+qmjNpEfjp2mwc+KtebCQJigWlcQtkeTRWAk3Skya5gpNzaEv/2vwfLoy3B5/ge4w
eLPuUtkCZsBoSdwJRbXpxue33mn0V8xRCYMhQEmh3nc9+CxkCl+i5sH9EUX05zU2JGTFh2NuF8zd
Fxau7Fct8ai0hiqn7O7wv/rsY4Pjuv9o2JXadDFUqVxJhDGM91+hmT6fbsg/7h4Bu7/Tq4ei67ZD
jEIg0g3FHiSOb17u5QHl7R/k82qaBZq/+yTPLuKopSx4gesM4liB8MS/rkZOhP981BRx/hARtlQ5
/6FQh02in6H80z3cRTuawEN87cDQM8/NXaMuu/P9beA70nbYXHYNGmb0R35y4Y5I99qg9Pjw2NhR
Ao+u3N3xYTuVRb1+g+SxK5I2HDAs3/xbIb6QdVcECaAiaOOdga0fOgFERsHPm3SY72ilIUIsLRnA
DjojVtaljM+Aj+m7Ka9PlcOvVFXUN07DA4RLS4EFD524M+nkuTH73saDSnpH4mxc4wxe6iRjXcrc
HwVQzvohOa8kF+oeDO+MRkug6RNS2VNldavfIKxIrnfeAnh90eIwN7J3j3+mLfAFNiO2jSnrkVsw
Qe2iKYJJMMQhz36KqId/FBpq4lBTwtC3Bb1kXPDWTlJ1/6BSbwM+vBSDd7WwaVH96JANRCpygTG7
lAElCd0+kZtNboR5C+FF6HAcPQBK/lJF2JRICW/YpLP96TTF2CZJe0M+LmcSWXbSBHS6qF5Eb70g
gIJ1wUVQqmgedkRz93fdXDp8iv6f0FAWdX8KMBzHlEECwz+mlGdWQDNF2QnJ2FKzvrFSVScDJd1O
yG1hG0QmdCwamOFtTb+Viw1grB3aKTVUVJgNfAH2RcDdYcMWfNO/cNz9JHp6pK0cEheXvgKGzfz6
S29aEXsAU813k5tqrI/PeJk+vu+cRXM7ey9KfFXIKY81T+hk8THMUEiwwXhjWNADaHMRVbpIfFN0
jQtbyjB/wz9ZmpBRiLWKt4pGRyMGJxCu9GStcJbNNaf+PvjVc/3hkq0eSQdFX8QQioQEE/I3grvO
NH5QNg3MdxXPLFOGVTu/6wpnfH7XySzaD2xLC57NpfizYiU0GsL8xkrJW0uLw938+905RoYljZQb
tLlwxRSWMkpn+6AXnGNwY0mRP97PKe2vD7YSjjEhExuyTPNuG4Ekef0vYNACJSgFX4eEQC0hmic2
DAOXQkV5I8rjAn7JNrhzVvuSa9snGiFGWPesak7EOEs8sAf0VmQt04tq0zuHZik1ULth++n5o8MM
wtOUuEAmWgGhFSRKH5WiCX0X/GG4GrKlW4+F0RJ8TJooUa3hfaUmpUKymJNtrRboZEVuBURqdtsB
qTloh1wQhSp82im4ziKk4vDFuYAc4h5dmBjIXXP6PdBaLtRquIjikgD8kGwWKDODg/82j38tZLLq
aLdQO0skaZu47NJFw2rqONp5pshff6ytOO83H6RR41rofnnk+jjo0oOHR/fX+Qg5JsRSSUEpWd8P
Um3HR4kgkOSV5gLuvyemC7m2sCFswGvGUIRHJ7SiBB9CsqmQ/jzuwcMJ8LO/dWGyPgxyXRVjN3Kc
oZl3rNo0/Nc/b4VfcmI80dEritqFjbljtRL56KjpeIh+VlUz9EY3h7+cfhOoqol080WVsssPoVGP
1FJGDbKoxcJTYtqmsR6LoX8zQR4unnkufBmFq3iBH/Zkg34lV/4EkNAf4vSzyvKAffYEyoP2eMQD
Rhfsyx4ZjjXvWAF0h1mCs5XzF3nNwOJDq+UHzRWTXrWO74B0PyDwFtUpcy42UrXme6owlq/9i+Ym
RUpuY5e0u5hQGpe3TvBm8+VIoWcLDT6SVKsl5TjOZizI2PUKKGio8jIUo/JM0CIJ1Zf7xx3v3pUD
kMbgfWfVMfHN/B09S+wI2sMCwT1RZQixWvroLJp8OXa5cINyKbdfgoWdYRA6DlotfO1a/GqidRKT
7v2J5k8XDiokZKSAtbArqNvkswfHxxI7Wasx8qW87cJJjAx7pxukq0Mp3sDW2TJMicehH3Qs6lqe
jT2JzyjJO9y9oaKcy8FCFEwkFq6JJ+80fhaKaxgDhMQsUELPtYSeuEEOLHdUqPPQgYp+9tDdoJRe
Yisq1pyZlk4IjU3vEdENtc7M/j4SceuWsrRXaLlo973evU4jJCxyoewB+4p6wM7OPaP85IUbtfQJ
KSjRff/oznZmNXDzIOkx4NHGwMAWYq49XMqELi3GHBJ86Ya4h3BoEY5wlAxkeYW57a8xbscb1Mf0
1m1i2N7l5U0zfLVCr1e3iCwMZjxnvsVmsQwLo3lHi8M7zRLCdMFEPDbeaJaG3q6cHzAhY5thblgO
OzBqbpbYV91ShJy2Oudo+R/ighay2ciHBTcwv6j5ixZr816KMqUD7SlSh+ynBacnSMTWLwmPkIIr
piWKESp+Lin8npykwVdH4LyUCcRF2wDhJeKl9pOW69CqZXvD0SU8w/GKTXw+k6UzQ8U/l5r9H7U0
ydPtxeXbbAkkebHFr/wWXUqTcIkTdVX4IYim+XY91j1o3LFNKzj120frGjjl+5SDNGgoPcv/X2eD
SHMQPQMx8gr++pjB0felVClzkWHRpGlp1cQ8lqyCbLSP6NGzHXRfk/Oo3u7ElBCLIfuw5YqiGBBY
0fLR44VX6Blh/IEKLn1JxaMlN7AnKjcyLz39xmRDrpekTxWvb2eINoDlDVTGizMhLXkMLQJY/fi3
ufFLNW9FR0PWMfPCUPqk+cqIiAmjLoaxBMGp/W+3/VYw2LTSMsw7Qy9jlquLELo3KJJAVyEYiiwO
QpeUZ5YupBSJGs3nuQCvo7bqBNhEK0f3xuTI8iKEsFIb0cclI4x6pZ73Wt+BhMriatbCYgwb6gT/
85rMXiwuxQQGDClYB3ipqoENZbhS/isrj3o9ikU+6VpKBm8pexoEp3ZIbrJtM9pp1uVYBykmy4HG
LAaHOgSxtVCk5wrxM5ZzLohC2jwwt/Ps2f+1K/W4oryBj4HYmYoNVYTJcTrzoXxCIWe4GJx3wQTt
/qRFrOVdutw+zIBvfz6F+PGPPfHfubhmYKJNWufrbOX6TYVT5cMCBWwPTXGE4cQiAI+NCSObj1Yl
/BLHpuN0b2wPK4FcE00k+9zsQJuI4+fi1kOM3VFlgD3v/8UK38e78aI8P2Ae7pZN9lueQkXceeuq
ff/teIm3HZdRZ6D6+ZxYUrjjK06GsB0U1wjiJOEWICZnRB3GW6az8IuIJgi9RZMysl5MUTsaY1S2
u2rtMBztYJfdBNu8esnMikYdsFyDyYfVmhvrSyTkFV/MTXUIpe1yrlZ9bUsnz3U4bczZlBJGYWlu
b51/NJjSYaXiEhv9qjifUCyjTrsgWTlxlm6hYx8uT1GXnGtFLMFr4aYoGmuTh9AhAAuk4KSrqy8e
iH9tmr5br3G3czZTrafSaAul7sveVBrG1P1Xcd/ZgB1K4+jixZWBrzhu55azCkQjQFyChaHAeNkJ
/zgBeSGYmXy/wCnJxs/u2w5lmTlamiDy8jamxbLGRm67IVxYESUMoO1CWIRuEG6tyuXV5eTiZP2w
qAnv1kyNid5t3isqvlws5Kl1kIt+HdoS51mPHCgqIf+3fS8ViwD787RRAFo0ZINCwmpOCvrufIFh
9zHYueiSs/a5+CyN/8B2p9J/Jl67++RY/11ZdUzvgqPQOJqfrXaqfWpRej0rywWwqtDGIkg25ibJ
vrj+0gTZXNaff5hSeTORNM/58Wxn4fEm5WMJWgtYI3bpQHPGampgGr3z++Y0EQP4L9Wt60fJ8Y2E
Dz0Y0rMamG8klbNC53AXlWmbhG8l5WZi2uL/2JdS81GbWdIFnU4CYh9BuC6/8EF8y6QI1LDz6hXa
2b7HsH5aBOhCPsdbpg0RjEWduUErHWrLVRdQhW8SYhxhXasKd/+g0Lgh8jshKvTu45uMx/PiXf7U
224blkieba7p/XQWY0mdgEwYcCZtrC7AB89erYbtyhrfX/0N09TVNYqrFwmsuenzk9JCc6dD9W4P
UdRcK0/59bskBHGDJegycKrs4PN5tyAscflgPL5hRKGMNMCFlk+kSTuaRluo7i0qQ8N/nLljNbdB
bJnz64dkl/BpomyQGxKySCtLDzrg53tHEvcTZ5g0T+3FrIwtJVDd1oIHK94Otp7TtQafE6rBJ6zO
J8Hfn+F1YcyCzE9wU81pGidW7ByRW96vj8nk+JVPR9HSRHQfVKgKw+5aFr5o3BvWvhEmwE0mqL24
rcsM8fqWKY/M4kgrHlplSObOaNer+38BMraj/74e/3Rf1xAMFSuclb3cv7BrKPrIe/JZj7SXimAs
fT56IT7NdzyHs+uYidQ2cPpkimAxn8iGS9M89i6GWRZKefO0dhJkrpomWTdhwX7WVHcT2DCDURz0
nMdII1Fs8J9htxFBagOqjKooV3vvkEQwWzgp6tuuiATakMM/nKazs5/on00NqfQY+4ezRB7hiZDj
bftlzaKFNri2to5KuZQ+Cr0TrlWnL0dmP91t7aAth1dalWvUH4ZTegg+feX2jCLIcolGwPHpJD1r
dv17bkEHSnV2lXOpuog/VNv2j31S5Stg113lYEn5+HXRbTy9ZO7vDP3ziYPX+9h76ynbdZzz/3Wq
DQ8Ec8+VMVeaaCk4wW+v+MIFHhhhlLXTPjU2BbrF3xxdiw7QDuM8Oc+JNzIrnuC8h/V2NFlw2Zjk
ZhFKDRwev71jso5UHiSjT8rrvvxRN3fVH+9LdYAN/OKjjGxOu/qJtO6jHtNfTMK9g08l6ZKqZVkt
z2DGr6Takz3YL4+8TDVTFrSvOf/jkLePGNWlcKvmQtNRwYLPFZxzPipgp0LYqk3QBAOG3aYywKhF
HyO/6FNNuz5fDWtS5+cz70bcppvZCZC8I6usrWDv36x1hS79NlQ0PpO9TB38ge+ZJKbgR/8lHeUQ
da101B4g31OpNYIlkp6fWkzfKWKqt+5IOF3R9DXasjqyDaXzDkZqD7TZ9NcQZ8WgHz/7GahDb50O
Fp2XlrSCWsqqGzqoLXGldGplpMFKlOwtBO50rk3XYz/uc+g+V0bkgnZABmZ4YdwsLeQv3/yiZtya
w4AsYk8Eacci3Y2hTauFZs3rcLniV8jGD8K0LKJxg0M7MRifJVi1pz6TTn0wK9f+36PkPYqsQ8q0
0HCs3Cq9yN4Inme6sE1fOdtT+RQbr05nn6UxGSLeQ8gD/w+41F2OHLPTRxj4tlwXueBAp/Spnqkg
trXSHAuMEGmxBkIQJvu4ZUiRqw58kwn3BNboZDcNgOD4My+dtIvSo3hieDL30kGNUWIsuG4dJWKa
DikW0vix+BE4W7GuOYAkKocEr2cile1Q9tqZaZYDUt9pdf0ZkvPRPmASxWADOks+ekiAPJwKM20X
R/p4LBruJrRZRZMfUkOxgOQNQo8Wtm9SsSA3I2i6VgwT27pjMSMKZcTDhMRXd8e+uw+/zwB1dy+v
vaxjPWVErUcAOrAhqTTxD4lWECvCEbuMhBrWdLfBFNqJ+7IYi0kEfamavV25fLxJWU1u6eMc+8ik
bQ5whHShLIHiZdW0eUORnmEFWfK1m3o155IEbcX1Gy4fIKY6kl/9ajOEwBv8dDeg2LZ09CAO7236
8NSx8RuFNdHPvBy8PfbxrPTPl/eY9vAhAkMlYL190kyW5o1KpXpWJKQ1+b6T2+EFrWEV6OqLBCqH
HGoh3tmVRxjVccikI5e9OchVGBvK8AXbXUWldWqkSlL/nBI3pC5pUKy8spA5OjV1oxdZOLecc504
f5x9NjYoUztd3ka3QX6fZOJ4xDp/OCd5Gv9fVdq238yKlLeCTPI59zqadMbByT6IJAkhwDSyCU5O
Sg+bgJ8/wp7NZsioqAFX4LPdR5IH5jJIrl3a7fQQvYLSExK5dP9xdBptmpY58gz5uJdtB1u4FLji
jI0kxvwPTdfaEfAx+OtE/8z3o6VCa/8h01p+HDaBNKYyq6sbOCWH/JL3bdWllTuxJ0zq/X3qqKsi
xv4EHXgK03UXozjX75nCisJC666pu0XuEPZVRmbWA1tjOQY/kW0OWjOfLYHCPUvOr2xPrUQAeZVM
wdc3vvvHI8s0lg3YHxDbGECbaDg7k5ojFG8YpYNJEsBya+L7FEIPwwjb1k0FQKoo8xye4n9ELE+i
+W3CSFoFElBiA02vnUFP8jHpny4EEVmP4hgxkAHmWpugfvSL0HuSga91VAVwi3/uU2V/QbtCRlxN
nxEqFs+i5VnYG/YNyeNLjSYwcXOeiFhTY6l8eYwejvzqa0xqH71cgjikJCKXtaOjHw3YUg25ZP6X
IsGIzIM1av5/fRd3Brv9j5FwRjxck9uw9PH1aXgkDAuQy8Z8I968XqPPRHYTLLYcdzQiuaVpUe6V
0W/O9G96YwtaPqSGfWD0UY6NhkzxrHY17F8b9yZ1uw4vz6jErWJkMcOztiWzcnK/oSlodeCzxSWx
Gkvz4J8iKFLVOdEqfng1p5c+ISTrOpCIUEBq0hxfyqdNT02q05+toDgjZowzOAHaASenpUyTbm0N
7nT31pMU1UqGwkgSlex0BUL1PUViWsdImEQDsaTcGGgkhKm54V5ET1PFQRHc66WSik48jtbozrNj
6A9UNmQT4DLwB9x/4h07l/ZCc4hDpCyDRTLdxw4rmEnPFkdtdnRvdJ3V+hPRA4DSHMdA8EBVNDPf
uM87MTpn6HCcoy8FoXuQNqeO9qmJAIVrQXC0TTxZrl9XWPC6cV4gqRmSqP3Iae9sMJeDBiR/rupD
yQYSc7Ghs/KAmHV7ozAkOaolSC95nzERCRzpkNLup954qlS3jvuHTlbc0d/6+XqSNzmLO951U30s
CYXCRJ1ZdFzpIs1kXb0dmJ4Rzb8KoFk9GXnYYPOWBqeQzDvabdh5vOOP3Y1LFPm9UEPZNW6AR/to
oMGzGmOoEAG0Dhh0xD8X2exHkm4ozR5qxooGgZgwtCHIcDv2Xeoe0klGvY/lsfV7rL8vVK5Bpk2j
zOFCVyTRVzBGZA4u4sA1m2jKN4V9mrMBq3DXuVlpg1NIrXOxmEG+qKk4DaDEPRhfqnqTuQDGA3Tz
iN1LS55wjCv8F6KlYdcvQfQEipApjlpoARvk+aZHSCOmp3yuVylovHcE5Dgx0SjGlNvoVMXyKTcM
i5kCpa4An+X7ZLSENVz9AGpVi/0Edt+Oz2pVsFpjO/TALCp7EO3UohNo+FI/oExB1ruKJsw5OKBm
bB2RuL3ZM05mb6fqVEalqQV0WaSqygqzaZxJlUIwHav3b4IX3pr+UVKrXe+a05of8ybwN/BTa8Lp
5xK7nD4EtfhzbapiS0YXbFV1VLQx/lM+F8XEbBxrUuI3XWKG7H/EzFj0sofdV/5+qVA9yIKbSxVR
FacFqIppOnmaGUAMSsfa4vAwS8IIdOucy1hTGwEWPJgttePRFJIx3QMScavFQoQM+njvxlQziXAy
FglTxsmtuqk7qGtcPY5++iKLU1YFvW7ozgdQXkhg13HVdNUqCWNJuU55GvqSUg6SxbA6vk+Z89S8
a19tOlaHcekJDpX5DfWAjkL9yPvWxlzgbVq1HgcgjCvmc5NKeD3yQGGD1NxHzs8Fa83HfLlB5JcL
0bfkyzQw0c5Py0o9KHZ9rkzG0CEYxu7wz+WGxHF9jNW3xdpe2mhHc1tzdVIFdPQxNx5Nl/H/Jlss
U88X6x4ZXDNPXQKQCsOoZfaRaYSxxPAjwm7cel2MFp0zBl/ScBjhMz5Kp3mNSQ2rjh7+h2/Mz7qq
Enj0uyBF6p+dJh48ERky+Wt67v+gdz5QThCPJ+l6kQl/3mAhV7UQ61wzPLbwM+wv2LsDyOxjnnjL
snCszy6TV3UXZ5uUuijNl15UPZ0YZuBR7Ikb0plncPRMS+BSl0IX42nBSO5tpU64WqRb4104rbox
UG1lqXlM1fG6HdocWVIv/fLTYbfl5FKKgRCs37LanmE7T7lPJKuwRL4WedtCppnnwvgIA04h+GwF
7+te9jPVkldqPQuxASZ02TleEttz0Vw4Rc1qOkyLlUpoK0RcNYYpxuJuUbqSF9uyc5Tu+6SPOoVu
ePmmeecjk+QmT41iJyw13oadI5smnVoEWE9lnqfLdCkTRRDgiXk+WxOnzKNMQYOgX2eTj076PO4Y
TyJfiO89VistH2CfQZQt/yXeQoT/o2elBICNIG7233CSCCPcm1czj9JyCT49ZBAazemkVv9I5O1X
U3nNMCwDuWUjRzbneuw0VFgIJ98XqeEFj3/5Ko6Ef7RsgKAW/ibqqKXj/Zru/LT0tV0QgYhXo6Jg
w1n+KAz4ucr3ofJqoo5eOV2CqVvJdMxTg3D4iLP64YZo6jgrrzuIKk62gH90wLjd1tUXkqozT19H
gz/6CGinqKwYpL77Ib6GAB1WgAzFnibXy2x7no6rjP6e+4vXq8vGkjAcO+jUft0tVH5WAzOf8N1Y
WkxFA0hzMsb4HXlClISxXuDBRc1EWbpRP6/hKxo6JKobJdh8/J2RzGaAwbooRS6yPqlDtr9Pvhft
asgbDoPk24TGXFWHFGjUKBg+gnIYsdTLNm6YCh/dgaWF+OiIhwAcOolbpLgcNRgdflAfrNLLEKFJ
geCOlfnx0sXekUor2g5UqFFvtwgdHJ5r6xXm3CEd6dnqOR4MSu+02+wF7Sd3N/XjItEOtRMLFwZn
E3c9ntBoNfRfvDMm28wOXCagvCmcq49F5NBMe9igWeZxRdzMO7j0B4a4XtKF84mNBAbzdhQ6A7BT
5K9tY5cWBMOBlQ66K7TuHk/6GhRC82/YBxG8QkfrtVE3NDSX5H8YAW1iwScwgFe/gFqLDCYURC3K
AtGc9gGGsRiwW438WeEugsGEUHPAQCBb0KgF9R0Sd9O06MrcLTCkNqrRGL7lR9fQGFa9uCDvys9F
u04QDmoDV0eNUosob4ridcGs0FSa0AAFHFCx4AwDDn6nmximUmqvcd1etAb5NDPyFOfbHBjUdyYZ
Bo5oa2WSoA6V3ch1n0HoNLTks5HgpQUAHNZKZCr0svPqfbxxwV/hPtt/c/IBw1C5DGIIhI3yxi5B
8/NXDcNyet2i2WvIbFJcxrHGAIMfCBnNt5Hz5DmYKmnkCynm2Nk5oDrh74DQUS6Emh5b7wvuPJ6n
TshiW4IeQ7CR2p/63nx0zfQhN7U8IGKEV2NPgEBZVUI99J/uz2vnbVepabkgRBhMeUnltlsRDsEA
RaHz0n6sDhqmg9KYywD+Rt1tu4souPGTWkQdM1h+o8HoLd7og8pr5APzKlbKxzE9XIfx5FOh+b0u
JTYUImhFLGEQ55z1cY9yYos4+PADhSEihdRAi12mtyFrU5WSmn9qr1NExw51epMZ45cKVLVUZyhZ
8l3WnWNIvcIeLDheMMmF0BQF1wAl6onedwksvPaRdLpDHb7CjsqCuv6sfNPt03y67I/83o18nszo
yP/6y78dpoDFH6AL5ihJuyuk/5Du1A6TMbfsLxX0bdM3wrI5eH3jiM9hX42avoB7l4KlikY8xDXb
P2bW3Qq4jpZf0tKWl+TUok6Drsrv8ZTyo2s0m5bw0Z7rcvHKdiIrS7t/Ve3G4ovZQJ0Zdm9aDdBk
xKPZImRWyQqHLMJgA5YwuGNIXcdyyuqDhfgo9urDS4g6EejCtncr9rysCxae50uyFntGu+9VKb5W
lGnNeooAVEkb1/+bN24/zRVJURmLXFwxiIVR7LKutqnDVxVqraiiNiJh/c21qrHHo6+7cYgFOInD
qjwH1Vk8IvRkdJrfYDpYTqtAT9VYKzhw+JJhw480BRhuGWucNoYOcBAV4KHHXOh4ji/51fWm3OHj
3MnztHy7krDD1RhJ4wBZRTE/MKIL9cAbvRk1XHaP18rARXO80jLn5Pw5JP9PzKbnzyFaes8fOwiy
Tst5/ejvtsGBMXvUH6/fYFGF3L6STli3zHYldxUCNxVS4VLmk1nrTaVJIU/S8j1uk8luDRefgKzg
PJ4GFO1Nv1fW32/MCb779bTgOVmf5pHspwxUFC93u8OQywZEwk8llGeGrrKpDHZnYQD9dTWXVtBz
XIO1BQP7fPG2ovd67mDMs5H6dCXtrwMl34udSE4ZNC/p9bmSRsC7tRk2FBTRFfo1xZ2FYD9Ev/Fm
FOm4H/+zrythLrG8XWIgOHsh1Jso1/08S4+KpixDIdAS0SfvhcSJn8xWcxBmAoGXCUF+WzrIw/Tw
cF6pJP7XDL+EpFSNiqBs9nnpjToq2R0tSmZvn6I+4FQ+k3gQiE5X5CZsRR7HBEmK2Qrqa3S0QXw+
Dzcvx330jj/1V2SU6bwUvWc1SACNUi0+87CboGKXbv0Vdk0IyAT7aWMjdT0NmwLuN1ScmPJNl6qX
rkMEVjvBVw7pEaH2MrWFBN3VJcKkwMJbrSsbv553fgwgMJLpJ6czzRkjDmjPUHvIceCtxd5I/16l
vNiK15oCQf1Bb0W6fbruipCj+v01lQ55SVPc4U2TVAS4GGBEb5DAKy/uqLDlT5cSj2wITT050QBJ
zi9kmy3YAs7EHa3zJMSUcMqRwlXSB3lRVRX49aK9qTWTd1wSSHVoRB5044CK/o6RgI3XZEgsBQQY
6ugmkIQvleRYbpdFVpSulgPWsLtUfZmwh1hu7hlGfOJcVCPVjOQE3ovNem4m50GQyHPIMOTgUH2G
/qFMZz+QB0Oo7HJ+lHTqi0mU++ek/QfO0ZxmZ86lzToki3srfb+tun4rdyL1SXEkftjzCfWd+mkK
4kbnsaJ4uu/n3y1eLMntCa1Axnw9Z5WNhL0Yigvkj3D/RaWe4aEjGnwG8d+6XCtStWO/PkdXdCvH
1KEfy1z7Tr3SpLDSu9aCrh2gBAbzwH9Gcw5cKXYKctYoU0VAwPMZRGpyVa0tCdkJqRnJgPNLE1xw
QQ8DvRZAN2N7dR6oWfD7EZ3+t27athanJbntOQB0YiytVwOusko1KL62+RcQooFtLg3D7G2EqkFT
/0aBXTqvsJq5diI288JXZvvM0bscCZ3d1+p8aLwyZIDA6G2FjC9RdOIZ2gmlJ0Il12DHQt5be0MY
84lzB6FiVbdmB8Tz/e+dcYRG8Xbg5CWNLJpHSym2OjJF3GRbkU6YB5oqP8jpGLl82MAnfUVDolJz
3RW49Gcx+w6rUYO6JD5xoJOGAJ5OrRSaeg5KDIMGQMOzo+ptKCKJ30HAsN0iiBYTIAk4MNit2RZZ
QurXmocA90Wf6KTlTPrFBTILdQVTA3AsOXC6QxwDfjYd4O4GHMtUkZtCKHwBqZ6q+sy3crQtKugS
Fg1NLsRHcS9IoXT2weFIoPKN/3WAqXCezVoheTP6WOdSPI67Mw7MT+Q9xQjkaz5RJDo6ET8SLBxZ
igHXvpjEkomrxVobIWz1DC/Tq3+qWH5J1k1EMxGh1IXjT86B8qqTHFzROpQLhds3D05M0bvXiuGO
bmmC5XCgWU80n/9KuSW3kvrPAE5CnAIeD2BCOKzcA32IS88brD+LRk2dDb7J192W+fJNmqnxkPzx
E5c2Y1SYy/Ge0rrHvs84IxGbCS5+mFbSobfm6s+UE8KMwBbmFtUOnkJZEREAipiv8racscvOjure
kNimmPx/C7rKQNvVg2J6y9AJpRbSoz1lS+r7oNlYCM6k97qvFiDQO5rG8iNeTOGbGxZaJ4D242oV
Hb+vz+CuyYsDHdm7nvGuKGX4XRGApGOHZ1+UyGPw7NWQxemcwwZms5O78I6zQq6bYSgCFoVjSd3U
ijy7ZRVEACby6lsVaNvdNxwItHlyJKVq5bD2zle5oYUJ0y+sJ3Qm8k4l4xW/shEhaCff9yO+aAKO
YJkfoQfQRfRTUOA2hoMfPrPUlS7IIeE8GrQO9Zh+Q5sPox09zP8OQmt0M6VMsAkrzW1ZOTd5GZgN
4zSfwOSRosP2rIWU9QDsVkvWphckQPRtC0sWlYlKPUpt1TcYiEt1q2v2cikHoD47K97fFujKuckM
lGUM5MwmoVR/+pJn3xlZpcsdmR0TIA4DuO/qpDeWhSl818OJSV4N6rI4/mlgig4B3zbK3FlWuLNS
oe97dNrb3VN4uFZcrjoZicmCyjcme5/1rJtWWmi4FaUvU83oXzBcGA9ydxg5wPWtnB1thX+pTyvM
9qYjTx45bVbNbWQhghfy1ZxjIsvzryQ994rZrh/uhtfcwnz07Iw8yn5Vwyv6E30adpGfTRyDjSjM
K/bRN2X6J8ZAZZg9ApglOseVTxXUB3lEeviZ1oK8Sh+Em/hn5jw533/Y+zMzyd6wE7BTU+Zpo9In
rNPnYEWTkvmarrI8fUN9nwqNFzRuZZum6JpJIJIV1ph5Xpp7V6q2DH3yaI8BO0o1yyZIXhjTb4zh
Zz/1dHWELFHTZS3j8Xmd/dCS43Zv7xicQVu8+d35wwcebQlXZjIV/ZDHM6J8o40PvzfiP1sg+wqw
vzHMJ8uZNgH5zrw9v9icNfXs31ewNg+8F8AKb48HSgatV/2NWBnQisb7dChi8Ny5GiPQvTDvgc3Q
gqbPSoUILl28zARr9jKX7xRqcrOtco+OiIYtPocVhuNCsnZeaUL2QdK0RI5179bBIAr9XDQOqHh9
VW4m+BRDllP4UlXotWVis9GqRDCwHNyvAUB8d8aH1ls63OwMNUBM1t2ffJMXfJD3N49Z47ucJ0I4
InP9MmbJCsbA3zHzxM4K+vNaQcTKdz+NHyftRdflnhfZ2Tme10AtgQmTdGhqk32xdoC1LuNUJHZK
fNyBbxj2NhFgzLvn98W6+4rzkjSz+xO3vMD/Z+zKyCZYBJEiDs1UPa4Rhf7tnqf2jlEOJ1GbP7XF
riz6v6uBv7jJiru/7FhFqcedkIjEfJjN+i8MUoMNmhG7SfagMNnLrogNWybADPXVGdiKUOz5Czx0
flgNUep+RXuNFYRg/3UJFujNk7J4cJ2BzobIN8bnendHvJBdTS+ojNnADPNYyo+D6a7rQ0WV1iS3
o+yR5Mjq1MwsWJWd5QlbSdnDw0j4xmOWNQPTNSpTUkaKzGxqCM4eUebACJy68Ec2Eofge/ifteaw
jNk0DkQ+IIbJvcgUwnrG2v8HKsONIT4tXcKY9clWpGZio8WIUKTo4nPCeSCAqKc93YrYm7H6YzRX
5KyAUoNhqHTBFeRhK0D/l6H+mWp0E/azabpOjPHNgDeOE6TdVorx+HE54CwFdS/v3gwZ9ZZUFEX+
07wwU0aZwGb/QwvDZqdEcNZMgEZKiYyuzFYdVdsrWh94sJoaHcVZcVuhGJYaHHb9UM3FbNSSC90B
JW9y+WGbxVtXL7yvTSfV4lVjJH8bh3zcQ+RI4IJ8asDMkBHkLMoIGFIeOtazi21Xq8iB7QbsscPP
nx6j7aMQ+p/Qxi42rFMfIKH8GOOCw8g+9S0y+57ZiYdJ/qO34MMfA1zlD8Jp3dFGuarGcw9eZHMj
0dnkwRrVyZy38qPhny+7095Pp1QfoRTn1hVgOj/9DjkQT8/hNRCfxckA4l7D9NWNvyucLJ/URrD5
Rb9OpEhpd1LDJBFdAJ633d+rNQDVzjxC9619ztf0+8XddcGn0VIuY4iLmtcEJpPkdFozw0GQWayL
7lDzGL455KJmyunu0T3O3fstYDIPgOHlsG3KY74dPOpEnLiAW4BYRTjOErNZ12xCSTDHNiUIQyW4
A+5zRPafGd3COkZsDJ7PSNQd2P8kcP8lOxCpu+j4GbHWKdMLYRztaeIVAAdy2FUT622CthVo6fB1
g4hpBAlv/lXhGCqmrC4j5wAsh+XCQyhIBCHuMw12gphmCtC5fnc1tqnI4kjizg183ra5giLlFNub
pbg8vG8KancWoePzciEf9lL2LJZVQrQ4kY/jnj6mn7l79tIGC+x6PS5qGX4pWpC2/O/3iGS/dKgu
XOq3hprsqgf+LK+/O+w3iGn367lBIpPHmTHtX1c0ztebQ9DivAclSiuAszIOznIL8pj7E2NXufDW
//mkuZocvEP7sTp1+dSrMiyePbcrIn8v7k8JZAgwSQ+VVMnUTr6xZzq5ASBOF4DzGaiOyW+pNINp
LVdcpOJHVnX3LryZDa3iYUxpCk55R8h0So0+WLwm0VIbRqPKfFjzkDAD+K1HLZQZlC8UbOvxRX9+
0o97XER+0Uq8kFVdc3LYVnioNIpbjP38rBq+Xh65mMySQuukplzb86KjI4fPS6R/Ax7vVcN1Jcs3
hEL26YtwKTolLi5eMUuUA+63viw5THUiTRtCLTFZcISbCx+HRIwz3rxegA+T1D6voRbmBDdcvfcv
FQQzY7akC+5xxbmOd5mKLfayasCGiKOHYq/ZZOJWh+mIj4PZ4KO9FBo1bROd3x2EjXprzx370xVx
c4kYED3Cpy/nsxzp+GnAwt7NxqUrXCuKPj9uJn24i4L6i42tfPA4IZRi90FAudsVVaV9uM0hz7vZ
2J0mFqVdPGVXLIGoqj2ekVkKr/Jw4GLGiUGb3izBovKYy1j6CJ4pTj0VdTTF1/r9om/b2b6iPUdK
zZsuDKlwJ0fh1s5Z5JkQZj/lzbRUOpjJNzigDp2bZFN97vyYXsn6NaSkZM/St4+oNB33naZxj1d6
uXUjVqFgM/u1cCFLrRtgqW9lYBBoBKf/Dmec7Tm8OvxDk+pbtj00dDvgX4qHgeR0zqtMLjFSqS1Y
NBZTH2uLJ+2//HNT4xjRjQ7symMA6QfbO2GB0kkZP+jSgviyPTYmb4+Rn/FVS0+XwawZsPMhc8aW
d5G3DjYcjk6twbTR6r3lD4mXK1AdK1eusVWeKmGCluyeoiAkh4waZgGowe7PDGvPXWMQYhZMddqg
mDE9h910utmIn+oxTe/AHS2O5uT2XYyFyILy5ilLUzd4UIsiNo7aPJryTIG29vH6n2wWmUGV1/go
2dNu412a6s1B6P7MYqhu0peH87pex0NYT+Ea/VHQbBmHoCjeQDG6Bj0OreD7HQJmXVEC0Ql8OOBl
QUcp7pHHzPQrh6Xgg8al4+nTA0aLN6felL3SQTnehahiXCeYoXpZSePHLMemYD9RvRCAzYvUyGRS
yyLS3aRrycHNUI2pMnndnIPJ60x8SwX9nA6QP3kXlaZdRQNMh3rVEb7uX8p3+yXLh9KC0vRfZzQq
Mo2AyZZwzn1AOZX5C/HKCPN7OROpuXYA7NfSchAu2yckJmKugNZVh9STS8bDrUJWQg/AA6f8cWpY
TQMFh3rbRTuAkpivdh0CJv1JGKYHfJwaM0oJwkQM0V59Ur7jtOTTDio2k93nZxmqzek4xzfLvY0b
HOwglj724g+c06ZyFnMvX98WF6ejNzYeDFzI/WU1PfcLhjzUKocb8CA3/m4zpp4yIoCvSq5VNe1Z
dPvWdDBy4qK48RYdUpClKSq/xrBJwDRquN4/+dfy56Un1TYCgMOprjEuywWkGo3FxLI6/3NEFEyL
JDm1CY2bYyn+LsWhHloaJkCySZKlT18hGO3pttxm49zqJ0p4F6es99CUuMDeQDCdkFmJfB1c3RuZ
fEVZKiR2fWga2K41rf7eEnaQomJLEZk+sqkMfZVBRxLOHcGgWjBWmGBhmesLqGeyBUep5qrZR9qV
pUZcDwv4h8PDo+gWf6jOc2vtK+fWZtDdGJUEpRZMcWLEPntboObY3UcQzMtOmWIRviMO3rTIKUn0
7+pOtBFF/9lwkrQWXbjwu7e2Ni0gTwyE3ag+MeZ9o4z3dQ4tzgmrJPRrI1kSvxSV68LOCQdAB55L
P305CUsz49XmntKIxTnaAqV7YmilrWYC/5JeD1WWzvH9nwr9dyOyBIxtznn6vQGbggAVOzE/bPCY
CJZSHyg/3xkhjeq3SLNe603QOow2jg2yexDXv2GPI4LGcem7Ye8rcwduqPqaHXg0NhEZ6HGABowd
k4tfT7piv4w2tEMJhigJioMuLZv2UyMvgkOAdotOoMCAj6wkLgAny/XmJMXijo/Ufa1oIfmsbzSo
82XGkwtuVbMloQkKKdEncYR7j+uL4AWGs5h2DT2utkjSjCP9rY5KyEk1x7w9BxUejwW5QFhff+bP
jZaeuqpiE/tWSXF70dn5riBqV8HzQzq+8TQxOTBiXqtprQibsLLeOM0ewkZdpVQVAAKlz/sHAicG
61FzjDY/BMU/HFZMrOGcX/7A4jr1aoD0yI7pmMt5BNB4+wpnWN4l9pPQxG+C4eU7RmYyBBTc6ZUl
8bUWgRnJ1KHPJNbD4CzZT7m08EvSoYfUZ7gjkehzAkelsN1bnIRsoOhSv4U8WmJINpYCTikZ5hs4
wrgXqsL938LFc38jtGNgfZAlOMApcA0drB/Kdern87Wwz0eqoXKtPsf0zR0PvWBfURK7TJca9BWH
I1IKAUxYqphIvO6ks++/DxPZmUlkkZOi8JD6y8zfrTHiJq2B+0kvDKFAd5MFksK5aOWTMkg8vIKE
KkYHJydOBNdpSa6qPLTqESOcLagTyiWmluHtsKapZm/im6iXYdAmN1qyU9doG7EDwGOrvM/aCGc0
VDYxrZkZG8wg9MBEy1JfFIE9bCU/E1UxG2mb81negCQR3HT5ZtF+6cA3pF3diM80ujMNyCs0pe4Z
kh85Xh5iKkBhHxYIxw92xhQ4gT8Mo30Rt8zqUx4IL2IV5rHjN5vTZN9zjuiMXjt+V8Xhhfae4Rfp
73F0/h4d7YG5ZBf7hk30nr9QP9ON3cUwULpeYx/Baiu8exkKm3vrHyBQ/DQMbWrV+TohPLTKv6Zy
fu+GXb3m1QkOE718mmAuMMKIezP+Al//W07z1zFZpSbhnY5o2N61adCRPDDmi/g7kubpU316om7S
BaZTz9vRxzBMGh/HXdJrGd1Wu3cq3OHin5PSqtEFNnfsYMfurD5ulOT+NszoiRN/4CH2QJzTJdET
87TBBfJzx8G2MOmkm2DaC0ipgMkgRKZSqrqxJ0OCiITsU0JVLrkW6JNFOaj7gGaD5/SvgKqqF2y1
kWzAjNIjyIQZQKr3HbbG7VruHWAWpenq0vfevHVRvfhLXlw+hN9HMtezLXYeK5KNxb/tT6sInybs
cjtkR04aFbhFeTgkoYvymV+Zzdct6kyqMzgw4yFlN3fpSk2hgthEtr1SkI3MXx0OQPR/YbXaEg2j
3NEQFRVsNUgVFc7EV/R7DsWayRoau4xrGDCkBEM0AKoPbGRmCiluThw5Knl4u7Q2Z8nyl+LZVoz0
Cfy+RLJwtBx+uEfDiUmSlKx/s1wGunGR0kozPjaPgdAYVGsziDouuN1O+fksHJpm5F18eel9KHSS
i3G2vICJteeZOkDct/2jCLjB724UEzkn0jXsUd9UhBo5OM7YfY1STWv7LQmLRbLkJUBB0MYPwroW
R1Wcp2zs6wA8Z1Q+a1Y1Xn5BHe42CTqkWniBKwKW574VHu2ZSFpEgwwGZN9BUYura+QjFX0I8ZSJ
cwYxccnHIzkx89CcmPvQgNF6QqdryK21T+fkA3l+yEki3DwH/Eyd/1344snGn9DxZyMv2FPr4h7+
w3DQuvcLfzVCQh4dtFKXw+jCqN804mtFvvwLkxw/t1SLiKE98U1sR+fLyLWWXOQbpZvMKpQT7KpU
AhjIwoHOALE0s7LXSCXjcrZzQ1ASkEGL1Xi4ZbkfJ4IPAIgc0biq66LKrZ2DV0CwpojkPhwwgHq8
XD/+JPk7wnMzYDW7sR4S4iNLQ8OLiUi/tgyK/4hm6r0QJUofBRw/GYs+LEexTuVg7qdAPbXTix/J
pnrVvd6jct7RwzDt+G23CStvWEX5QbQxa2nNEqum0Lc+RDAiBmBmyTy8QYDtheRJlHE2iPaIWt0o
5jzCyKJwQKXYwIOctJB9wWJBja5d/uwT2WCX9mmkSvVD9WJAs7vjhVKT5F1YDVDfskqpKEPffPNW
kYIFLRfxD6S3Ri+AprZzPgXFYPr1YUcMwCoh/+yqv8+3I4OMXvyHfptCABxuHuwvHnvIyusZjUkZ
+r8llVys00ORkHb6UOOqLH/y41SgklmNnygR72JMx3EgVzjWOT4ezdA+tcoyXZubD2T/Y3Sjb5NV
fKaGlU+etzBobwiA481lcLCUnE1Ob6UjRvBAA6o4wCkKSfeF67JaZEYMoZpbxwTakQe4tk4qQjGk
ts5tane49vHDJUxd+34M4zpS8lttoXqNqEDKLqkZALQ/0JXiqoXhjM57i5ntticMVCrl+DokixBn
nBcVFEm/KLEbPHcOvXpH/o797/cMOTCYR32DVSUDhNZIQPygFtIuWZp9WNXDpCm+L/otRAumHGes
hVZ3MkAP2/hcb/V0Wr2ZEPf+Ok2jRx1ovRfumufnl/m5zXOI/C9kYrBUGjSRENRpgjC97RJpTGS0
ObRh2cDJEVGDb0NsTFg4SZX6yUOWl9Mucd938/Unlkaq3GtmjZjpKW9NkHI9R/tmyAR36a/Y4FVY
eYpwBc045L/13eZ2lYxvVPjSIW5ZP6NzPokbX1E0ZEDECw5qK0GF4D+2P5zxKsLANOSWR4KMEVZ8
Ud1vS7aeN55k0t0zEw22X8jdF4XWlZYduPw45PKWK9Jiyl9SXsauffEtGXRzZtnQhruB4n7QE1sT
7QCkCZ+CNpvquggc2medSVhL9NVj
`protect end_protected

