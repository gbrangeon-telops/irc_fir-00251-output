

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Jjl8vAn2UJruW+pwbvMAIo6yT6bQgTl9+ZqbT+VaAP/dcMa9HxI5w52bG1uOMJkKjbI3shaTb5QH
+WA4TEmwBA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
jY7USlQiP9PR+LALAEYZsrKak9VnF4tfhT9SQb5jLUPXs+eC5ZbIVQkPjdV+4wzhB7b7ai6shnHa
gEu6kUZZsMTRIotEQn7SVZESTAIMCGAU4lDLU7RT30ySc+gN3y2heOoScYVxVF3kYNcbErB9g4iU
iZLVkq3ZU0fP1VLA30w=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
W97r968B0QPwlTs1emSg8mtee0qHNpQ+/n5wfXS0R66Akqy90VsNXhnqLJjbnGJNqaGSMTKCRNVS
ox1Z0rkuemlJn0dMgZtmRgHM/NeyMTSbsBwVvTSeFdA56k6PzciIIQ1S8150Bxbexnd+b7l/UMK+
JO8+KzzHPEIPqou3srZGn9dog9HSSfTUIqvBgloCeGmDxxwlsFwQ2VsrffuE8mB5Kk9lHG/A3rMw
tbJURgYaS/b69KLL9Kc/urEgbRWHU1HQCQDL4hSKE79WXE68MZJ00kcWMfNfAOR1zytQecSerjXJ
iVVvnEzEtzUejpnuhHCRhS+b62dMTzf5a1Q4Dw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
l6IXa1kcvqxcIuqXI9bELoLDvGs5XxFfhbXxOKBitloxuDBS5IYgW7AXksTedGB5rM+6jbAr+PVa
4ykVDtx+9n1RZQ3HKQZNsRywuW0+Fcm/MhmC5isxnEClP56JmzAEyD9l7nmy9JJJI11qQTy86iSs
hkUJMmO3Ph4Kz8ptLn0=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
gEbAM0PoYz0kTXyuDtZRhRtQJeO0ezbVNuHzWd2Q6Djxe3WZnx453sNsfBBqykQPTu/zHrWi/wfe
VIPTt4c20XjDHHTidMXhf5YGMYpytIjNmzV4g6PhJehJgJTQj+T/bAmaDaXLcqMDTjUNont0w58X
XTjVYtxQgjqcVftNf5PS5GCVpRxSTsKbT4CfmHhBwwsNC5rLtE2tRCpmB6tKw/7xf8VLLD8a23zt
cVvVNX0bw3bWCGFmWZjC/1fhYI19WFrjQO9Y/0zq8T/b6JCoxXV2HE4Z2dJ8uXvV5GV8EStC7VCB
DhBS/R4IfNLPojIIJPxvrbzkKlmuEkhgwflRRQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 57936)
`protect data_block
pYEBbBK5dQEHQVgDWrl5OiT07/XY25Tas7skSPjLnhHLd+i4z+fB+/vlL+WbnL2LIgkl7eX5hQ8g
9Zl3tDpiAZPFjV2TVSSlkWzMoOxfDWVk6dNAajsogEcnSeCZ+Q6y+ubKvbDw4LaUqpzuQe3ZOAX+
dInK+F9BTTxeCGXm0+ykcvcFCGRa9Ylkjb5DMs1DSKPifRHpN5D8kGnA+QF7zw/2K2PJviT1l1g8
waK9g1Yfw2lISUrEDKMdkTAMeIafdxSelweMr7jJqL7x+bQOR6Rwm4hEtsmiFHfVDySHHSN8aIc/
BWkpew+l72srcNftUtxfEqNhredbdZS7SG9SNnLjLjdcgGMC1sVc8eLR39oB8QvBLjsAzLTTR55D
5PADa7E6oxnIQEPaG8YaZhY9KORSDz+4UjSrRfl1PQEITyGq+qw0jKgHvdj+UxsK47dWfqdGy7qj
x7D7v9TtcJxCdofoRfrBlF/2euTSQMcsvRKhJapGBuuVD3L3sWKflS27+iVL+aqFibau9YdJkmfo
hu46BWX7tD71bILymJ8k71/71ro5qAMajagBT6O6bmTJlDylqlkYAp7gaSxqb86iWLXJfRRNP3cl
mGc4FBQz4JFh7XbKDb2RfiPzTLEsi4bBPZAUuVSCpIig0xg1+aHNflSCdbYouHIBBacMsH/XvYzz
MM38Z8nJPnhHA+uINGF4YIWdqTKh6141GTUMcb2aPDXZ8khq5fQupDFvFRn1D0/bgmvBsJjazoKu
hrvfwlN1Lb9OemwmYKiDaD9HJWQ+264jErURH4iaD5Lg/EQ2e6Ry6pldFZtdAltJd7ARrVvvkF4I
6M5/gYLjI0ZQLPLZVlPtdvIafV3KcpH2RKrWmDu94KqGZCqs/lWuZ3/OuB3ePTOs4XFenX12is7N
2ecobWcosUgQtDmFkMAPbXwcKmEx/M9t4HPvVr9oqP4IDh5tM8x/nQ1l4NFDH0IJx1x4t/791G9W
Q0Myk1/KUJBb9guOXmp1qT1o3G4W9l0FrVC4ZgArPK5m+rotRw8CmUn7LP4m0vDk0QKXPBacCRHQ
03lHoI+gynRb5Zfqo3qbQF/rpWCcmNAt/yjFtydsU/KugXvL8R+ZiAfgE7T+LzPKfBRffFku5ZGm
vGwebLtjhWlszTxcA65XG80J0tTzpimnu3VNKivVVku+hchlMLIKqyy2nMEaxgaaHNJQHrCTHfGH
uE170NI6uKev+Nr5s8sbeEZMW32NvNO1Ay+F3jaYrW59gTmXoor3qqFCqELwOETkwj2JcztUmEIu
JkMhsWjy7hajQwCLe69Vut9ELXDTWpRRnzNy5n/k0M7dRSFaAHsk9nceKfJzJg/N2gnWFabtyje6
i9rW6ZL5sna1sk3GpdHPyh8LEoYV5nfl7QmgaVEoUv7L5SHxGBe4Vo0Tl5Wl5Xc6ZvrkB0T2B1iW
YZmrtIMCzVOp4/+ohrYbch2QLPg2m402s7DxqciHanm6Pfs4OBng2L/hhNvPhwkKcDMITD5Fzk06
khUVziqhDlKA/9sLmv1JDD5iGj6uLQuS0UoIeSshcDTetmQAFgByAfe2jmnIe7jJEUfCIvLYKdDs
XyHXRFUtOOzDjT+GvDiY5FnHFksYNoye+mwFHCc628otRt/I68bp4PYVmzRqL6sRaHRRzm+ZpUvR
qUoiSWEhpf01y0VRGI1IoWBdx24gsVhCGgFNkf6IoPaPAvPigDi1ahVLqOcDAQDf2u272LWV7jHS
bC9zBG7wmBoz44rxin/5r95XG6XbAOYKVUg4E2bbbfku8I8eNgNGGgKxNV2351nOLv6eUGlAcSj4
DbulHboysuQ0K/jsUJwutO+jsEKau5KR4b0ZvQCr3ue9WN8PKdl/wzSlduwSyxyFFhtISxfvJSJF
6Sxs1YRZ6PDnlhN1E3/rSZDJ4dwd65RxZQKgos6kTz/o7uiWwRvDPn3tS+P9DY3Ts/kxt8L31vMH
lLYHk9Ez7DYolHyTqMT51o2woi2ipAugkbHnibQhIdJe17zHc9wbX38P5vLvQwR87M0JKC6M1T/o
LZScyi5g1cQJo/ZJZ1awiAREy9XlcveUhWR0O2q+Waon4JVNywuhvgfs1YC4FMVizj/tIW9rwNxM
Gmg9QepYSmML/E2W7H6/2sBfURJuoHsk780r5hhS/Tp3OnjHu4WIrUHFJsYR0xraP6JLnbQR69AO
8vH6gYkjxNA4/QINbkEC4pBHS/P6It8GvIMO4WAawIu/rrTqQBdi2KsrTdiz1ExUoupN1758OiSx
79F3u17mrFp1B+4kKCXLDIQS3geHdrsb+Z9aimXbacHgeJtxXp9crcG0+UHyE0nx+nSlzV1VrlnB
9WCldn4jbxoqWjZ6J6igVv8XgnOuBJH4+wKjKJXrrNMQRsQ1v4UxcSN3WjvwTBIK/Asig4QRu4ZT
HhOcDfVdYE+uToLeMklulhVKPQCZqoim+AW/NtsgpxUorVq23/LB7uUpL0SPoIBIS3w3a+6RRwg5
+NMwQHDiLq7f5GqSPikpmWbZ4NuLo2haJDuw2jjgxoBtt0EtndQsBm+y/2oqkg8WcBN/rsg2xuR9
hl5jRpx2DnnUDyI0erIZ2BHZNDDSq5wwiMSQ+0tEkM6kttveyKRUHclOUZm1MxJVvk2Bg6UNMwRI
jtGORa05R+0HgKoU3XgdF6vcKzPJnMTfc46XMknfksUs2tzABtDOitrZB+n0LUi6ehLoit+asX3v
cSimd0GJelEM4KyPQ/Y2LUu8HVpvhq3yuTDsOIOqC6rA/p5uf4wbItOO1rMtM3RbT1skYWJlHHhc
0rSLFQX6Q3TQgS57gFdMxcyYmopdQarevgutd/p8OMA/FUCZXUW24Xsg/uH8khN/iAUaoWl2+LAB
Bk2bnGkih+HTrJ4GbVeyJVOqxTC+45q2tayR6KHovXYiY9dBvSbEsx163ainTB9wlg9VlRPL8Iym
eZd1UVIjZczeFjMWPHk7gb0j48FAOWbjsxs+ZSsf/M8O5ExWbu0RpBwA2KQpXhrc69dKHSjBq1dL
Qvb9m1dSgxM9skuc4rE14HmdbmHvrI8Cpfv+2dDDAaOxv3ii+Z991LyL4/UmcSvVvxUXp4eKZ8jk
nQLJR7vOsZyTA/Fi/zNECIHmz2sssq+Tr1XCx/yWQ/6l9d2QIfHRz8lNcma7LG4hIgqmRX7opV8g
a1G+02PYQc3TvQEPvQGjjP0ah9BhE4KQ38vSqQ6T0Tw1a8mcwrYs/HkyHQ8zJktFXJ0mo9rwy8IY
vnWnxkM97ybp0wLmGcxzcdSPObBSkgekafKRfM3GgPGU0FadvUw+fJebxG/H8hl+c/koGv28LLnk
uBfbNV+fKC61SEENpm0MiOF3PeDjWBJipmzLVbOUxO6zsuoPbo2rW/8ZKenGAZtTNrOxLpgpmmeZ
G6Xotqe/ABJD6/hxAl4mya9Wcus6ur29f/q5UJv3kmyecJjkFvh9om5mLWP3Yf2AJmjg7MSU7e9U
uowImQ1FRNFbUIuZmf+O9OzLYidtfbypbNLca9Eqikkaq6WABdUGXijSKpJnMXSWkJasSBeg1+QU
NWitSbiJfmY/YowCmFiIVNiqJAK4zMGiakonM9aJrrcHpuD0ts6RhcwrPCLkgufJZbXEeef8C4aW
hkFY+xcBSNRD19BL2luFkklSQUtjpqn0xOg2CCZcBN243P0zOjAutP4GdoeWeO3BNEgYIoTHXJqg
jLzAfIIOpmRE/PdEZ8oB5TL8lqd42CMjirfvVGnCh22uvnMnUMoK+uvgP0pMF5FL44rPux1PN2VU
gYwbIC9uLrZgXL1i0781x+uUxOvUa1iXQzlQQxEUdUw8TMPfL8t0fsUc/5wox39bJhs8JfhBc9X6
ergM1BIG6/Yj0lkjM9GKaL6VGw9ucsN6h501t6HanM2muTeGhaSWElBEE5aruMz9J/LzuBcYACUJ
+XpcONg066trIQKGesr6330lCL390GlxTpd1TqZdu6qsjzs78HEIDzIU92Z8EqeLdEAK9af1pzIK
+/xBYLFZoCcSesuS7bCkbwVwYs1Q9XdJlLv5CRpPlRIPNYTGJ+MYZuECQj0/zxoLrQg7QZL3e4ZE
F2I02PcsxAHrHtrXkKzO4+6BcmV98IHrYaICLSE50K+1y1XIqbRB9CRNj63hhSfprN9P8L6KhczI
tFIFBRS5HImNKQFmSqElGB3ZEkKD9SyfOS9Mm2BwcT2Yk36GTK09uAUS+DOEeIVFgs+xw+JsgA1b
ZxPPg9KjoQNkqUTUYrbypLSh8WtwDBKuCbPSzQFKVMd+i5K0IxYhwMAMpcKl+40l/jE8lj9gfKbz
Hui2TdTfP26cLnY2xsFoP2qEe6hrzlJQ7r1URcVqIy0ZdKRxieDkdJRrD6Av4ydjcMxyJRrHtdBx
ZclrXypMlUka21xYxPAcZKCEPJRBYLuYJwb0WwCOfaBkWxpR93DUjGN/YTLsbgHh3Z6glUzALEGk
1f1KDueODBxde4+ZAyMWcq6Tf4l4ooLQfrRFNWFlSByrBZJBHHoO9EThRO3GHoDQMqSySor9COdt
WLSZG8D8vEJcigd6W4cD1ZYqTdHg4/Qr543EOeCMJrsOK4S37bQk8E+RP0r/uL5StA89M1LeHift
DY99gDtAk1VPXDSahYugo4+SKjRYExgkDe6YpUPUECKsqXhrqaAqsq6Pr4ymSTHayb+8ogJiU2Hg
5oDxJxzF+JJ9i5SWAsUCgdHbWShOO45PXuH+67lve1IZ5u45z/Y0fpw0oRh+Oq63Mf5KqzSw80NN
8W7BNQV7xHoyE/yxGe6PTIglngaYZWNtFGAKF3QcpStg2vYQbu69UUvOnmIGwhUyID4Ypdd5lqfz
80cMePxaZ/7ELIu/Z+2/G+wsFo09bFbbPUV4kKT7lk+crpwYnepnwJmF9RXxZ7XvqZtwxP4VdWFs
uiplJsyo3jdU73YIlA/RLcib3g+papPHuuVd1Un7S6N56+1lMpy4Rba6ygsBNFi0qQqKs2N41hlX
P7fUAuCel4ANFtgYS1aaNU43gcYBBKkb0CVJDtQUogcMmV/1a1pzXVgbKsdZ5raDmU8OfAEF+p2I
9Q+CIm9KSTM0ZVuZSbTfQr2OB5sp6RaR6ej9/ff2VANTsGYuiPZcocd7CBpBBl/NarVgLC/vS8Oy
5cV8F058oMfk1mWH4x5NyFojNYNeUiSBU6DeXNjdvf8Syzxmd2jsUB6gB7MVzPeR6fQdHkBnCT6d
E0UwrLaviRWAU8OKdSqZLKr279EBZM5RlErTIAYUu2tKeLLVZn/M2F9ViHsFoY1KhVzIXOgHJAUh
oXBRJpSqLQsmZdDknKAPaiTn3Ux3kmZ5OXk8WLl4KB97FAA4dN72u7oH3989FDYFQHVnbRohcJCG
28jMdQic/7RqBKTNiAWaGM6DID1zGnDLMKgCMbcgSmavb+f3WQ7ax3rLUKcfrrR1rf3MLwTi+N0u
oltU1ACYJw0LYaQet29vADtrPiCbHzuytM3kxiBhMsLRHSewZH/Mb835Gn2b0QrkxLP3YfyAI+SC
n8B+ql6zTHTUNSItTvecEZRyO2O+f+j1scADLlQ6yzKdJtqkdYnp2Von0YpED25xVe5IwoukBKy8
AoFHA8JSWMJrC1fs42FWlrpbml2kHgaz+HY0Ee7+3BCy0c9h/kOstwNRqQjMa/rwz3uRfjpyYzlt
e+K1s8iEpIodRT+woxUc7kM7FpGNBLdRb7IbRQ9/EIH6b9dn8+3qz0zRzej2dm9uvScy0eLlgjLV
MLmLgoB4zl/kXAjEsuNRDyFsKQZLjZFeSxRfxY2yJUrG3FHzcVEJaT/wzFb3tCF9AilBEV1kZs8I
lhQN//e1WclscgoS2ZZLq9NXRYgCxe8tTTBiDPzq7OqUUWB2MrTgWFWUajQkYoXiwQnsPAR4oXr2
sx85ZnMNScSMDln8sCB91FgLdCquSNxFx2PcxH8C3xE2x7Va/RpB0cwA4oP6cvUjwkKyoa+gDuWA
fuvjksVoFGQpj1VljHMMemR3Ys5z2foRJ7aXNa22Zo+TjSHyYJiIJ09HWjWLDh1wPUqj6+pGEQzh
E1tjor2sJfKTHXNmapCg45X3OxtvllNzuXlkp+AiC3HjZVVGf47K/eUOT2yeBUXmipS8DHq02JpG
K5rX1nIk6IazGA2USSEn8NVDmnhKmtBEVYZhMpq2VyCUAL1SFPmMpB0H1Pv/Ee1n8sGmFuE5E7Lr
yl2kbTwn4lt570ff+Nc26/DhSp+Cd5yaog27W6NpmxPx6GlSdPHfV5OSK3K3ZL2MEG39lUvs6oPh
Wo/SSNBiN6cs2U6NiTGX2f073P+tUI2qV/wZRzOD8i0m80esngVWVXgB6gH7IHrWgca94BroEzCl
k4ECa2OyqqtBNUOyVebhRrCL8dFvhwPkfGZjMAYAP2mp+Lfxy//8W4atZ3uf10ZkDXq+OiBn5ri5
RaXszWcfzAt9MAFKipKlUW8cAASFRDkSTYSuf5QIkvW7mkN6AzdzbmE8kB6NePuWOVMD3z4nu8YV
oRmdurmOb1D674412KIT3Yb+MsM+tn1hDy47uIMDpg1ziz5yO5R6j3QLXKo6LdHhLEMocLnGWLVa
V2rjSyLTZ00Gc+DXx+J0yTRS+yIykqwFEgAf1Fkaum+ozM21T9vTBB1sgkiOVrj8eyKAHDMrVT7h
YthCgLFckRbGuMbK82oo6faSwjO3FV+4KYQdJ3I/Z1AyK0df6stDU87uNrvwoEKAkNRD+QHYAjoT
aS0v7DkCAVooReY7FB7vqZbG1IyqWTdpYk1cCFJlAy/IrtjajmfqaKemCCA3Hfa1qAJyTUiGpUdz
N2hNtc+GRmiWILafvLQ4VJAKHbsz9c8sa1c4i93pEw9aCuHDPydsvCNXziGunUgJZNo+PbmjUF+K
ce7gzFPoo05PWXzb1Vl1OURR0zWa8dHeSk8dk3WBeQozNfy62OHTbgkGf/sjSm1wWzr8kwhXr0Vi
rIRgkzhE0uDGshcPtyV4QKo5bLrI+rsuWMlCU1UDsCNoXFfZ3gz8geyadBGqABJVHd5lWvOGO5ya
im3erRBuYJthq3u2wKD1iNo5RSEPOpIllovrp59yuPuLGtmSgr0yJlu+Q+XGN5iiN4X5AA13dBki
rVl0ll8+CgqzdioYEG6+xiX/fGFCB5g9y2RiV+RawpF/6c49PBkXOoLZhci1RyHUoFlimeVs5/Tl
7vwfh6Ck9WpIBOpvMnKgOEaFUMjlNClr1i9egmP5S9L5X2JSpdnF9g0lAutABfMNLSQM3DD1P6kV
gVt+xKQPs9mt7mC7FMpMlMIX8aOylulWQxBcX7/z+QR15qlN2mfZr9SVixlcsvHLDghAYVXO1l3o
tQa/vwU2LcSu9PPrVusegQV25ZRK/rSEUqlVjuc0gHbnPlaB3lJ+drs/+w9L7uhTttYEkOCXwLho
8f6lDcwg6x9N2iH8YDHHERGCWJmLsXCx0mSZnj4DFZv27Gwvl5VLfYcxp6d4H6vlbj0q4BPh1khf
U7ReDKQgDKwEg06ivYFBK1oitHF6+lrzOvzxlA5Z8w6A/Sc7pSFvA1sqGPszWRPEOqctWdSECY9e
J3xEzliTA75C+AHZG6I3HpGFe0pxUOailEgtlwqtu0ZO3nHc5MX+fzMhsKz1udnKy8z7HHS9ulzk
Hiu2Q0hMpRCsehVtq4b+PpIfxAkdgOlMB9A4ddubJOKT8qAVKXPbFjki35vsGtTC4L5Nvfv3hRwk
AZhKRbHpEC+EmvMY00Quij3m+eyl8aQDS8FJsP7qSamxRD3ayJ5ktgmtml2QGcH/4CMQVknMLolW
RpbO+zjtr1PdJL7GZKa7MMuPxnQDyKzN5PcR6YuUW6ImfVHVDKE3DnsvymB/zV4wzbaGmzqtDAFc
PZFnJ/m0yTY8NFXkJ1oCov+TdbVtjLrdMVUbvhNYaSSwWxAL+sqdTLptTvWUxq5V4tXmfVIIvUkv
rr97kdxSZz6jw8QccDI/3SSF7URaeL6niMJyEj76WhzCrOPh4603GaUh3bKrNuJ7TQ+nw3ovkT6N
zve7r6fRujZnFOFIQA71VlJBRB/uarIsV4UcqZEjxtl3tdd1LZJYSdiNKYUiHGhaQDb9TAcL0WXa
Np/NHHbD+vZ9vJN+3VTTn5XVgQ3x2Uzlg2JUh1VYHgfdh6qgj7TkuHAoborySht61KvdCfyJROXC
cvEAgLifsfQfNhKUhRWqZVUh2Gqa5tdzdI6lnGaEgeVJrQ4jkyckCj+bRGClCVk4ucphq95/NdcZ
lJLxGTagUNqWCTzQWx8BzG/DEgkl7LmUU3t7rBhuHewVo+Z+G8cnY60L0j+pWfG6ox+b0MjD26Rh
jF8G7ck3xgTdKABDLWmmYU0G9M0vDuxJKuCO/mUeyHLwKvvePNDvqw/kdcQEugUS86zHkxiMhnY5
WwqVWIAaa33ytC0E4B26sSMXaD3jbLRzQrS/lI4tfifiuMeU834fJIC6kjQbxMBinLoOu6SKQ2qH
SOoRauXY57vFoLahkBE3EkYNlHQOOdcCer8i6FbQ+d45cbt6rIX2lEDMOIa1NFvO9X8pxz57vAdW
R3U8GPeVO4Tx4D6q9Q7MSsMwM6RRBdadIKgmp0RIAzl0/fijKuxjteBtTCkU3NIhyNpfCt6qDbHn
VElbyYFE+C60kc3tymUELAFQCo25A9ZxgJeKEZf6R0thKWWFAVIhPYngQIxrRTu0lkDlNHSsvFtB
LDk1iwNKKxQN6KxUZD4Zn3XVRv2R0SzRNQ1qfs4RQO1VBy7t5CS1jVfMdu+RPEkvGqrHqiyWV5kF
5oYAvS2JaVNlFGn7FsqorJ69VWny4BBBUP1HZoWzPRCBtOx3AgyKgk0J6roSinEpAPCES9btr6/o
MaMYtMz5PAEd09qoCfNdMVdifMJoVkwrJtqTpP2VM4E2oczhal285Cp2J/Z/f9dKOixYoPgYeQxx
AEOcdpy1WVpO5vvhuCTtd8jr3dFQxF/b8i/75HPnUV8X6jhg/wYDX710N7/ghukmK09/mtBBAJ3P
v9WTlDqVma6eTS1YEqeNV8KBFuxJMazik5Wj85jdMcEbcmETbjPnOioJddcjT8+5wXtnunI6CUqj
kWXF96TKt4GDJlYN3hefUpduR1Jqlhqr78TkD/I0wUE7iP0YCLKAklXHw/LPlFU60wvkmqbDBI/r
jVJrgIdlTZNIQq4JQ1pCKXPGEwmyoMbMAXmJv/5HyfKXr68/iOfUdxmqWPgrnuy5zuvQ1ziBaNHw
bza9fX9K7pso81aYp4Xo2bD+5h0KfEny4fXpHT4rjuT6npMvXZe770EZVGOREzALnoteQIUyXEoL
uGfRh6KguekeAvRAsol9fd+Y09LtchcvRx2deVT6EkRRWDUD6wOsx/0Wia+Aqx2KMXyfNigvZNZt
CrpGnJD7D1HqK0VksbzeznMavp2kdKwQA+crn8LRmAy9GLTYHAxPAdq/tj1i/ijSMVU+UHJ55YBd
9/f3pBdilc7j5ilsKTWCsvMYV5y1WJ+Qg79Ye8SXohDIdV/ayqv5EKLk9drJvYGCUuoND9TrVSYH
ysVYrx94tXiMJVDEgyrpOTJuo4vnHdyypCr9KxZcccrH8yIDk/Ycg0CSmnbyUiUjoKp3eS+sdAEa
0XsoJ2XQF+VAbkt5wu/CwFGxr2/jALygsHHu0/ycFjd6AgfgG+aT4o6AMRsRZ92EHfVZ6wGOBwBk
m/rTHWVB3Cnd097TS48UTUNrW2g4tTonHQs8AxgnXWQPa8EqTDr5G4DODmb1uXODbTgjCF8A5bJ0
0q3Y0uZuffu7q++PJvKgO/5LAnqlwszUrxbjfYE26W0sa1//09l8NW1LEvDsYWh2h7T5ho6jS3e9
geANIJd/QpDYkH83m7+pPoDinpRith9k8NoyZCEqy9nxgZKX61Q4ton9Z7b6g53iUnjTEr/NgohK
J32dxVpoCm0Y3228AeSv9yCt2m2GGHJ9uVdCsgexmxufkgu7ykSktTzQJbj1SE2kEIBm1HHGmU+0
NC+6fC76iDoMQe1pdzzwMOboej78xmGS1NI3Y9r7n6sm5LkQkUAlBJJmVKxbFae+P5KqTbbYTMUy
ph/6c1Y13CGizhz5DXU2Besg+zjZLK+JoZLykvkIEZc5/kaQb8ZEp3zCiayExtXcN58ExWhTID/F
Ke2Ezf/2l3eXNlqYtUAUMxTS0nLgh88w+vpirju0WbtDTm/NUC5dxOyws6tcBur6knktoYny3CVV
7xooXnBh5MBhjgzbBQS3LGi1wAwiLITjK6b0gmdvJJ/TWXTknj8InG/4HsYl+LQiJ/zgBlDKpiJ0
UlFaJrFj3xDxkE9GpBAFLNkrWxnr9P5M6WH6OPAmmJWzhFj0xjuu8HRcE+9MObiVa0YUTF1jqwej
f29EVXwJJzKrPvewNRvYCqq3OaZgJhA6ykJnA5uoPnD3IoDfUgBhN7lovZTaPJNdhnNiKrx7ATwa
MtNGqPMa75IRPjJRW2jLX2lzn7/xnQ9MvSjnm6Cii6oiZ9dIGZ2TDDmXftVMVIRRy794s3NBnoUU
sg3axqlhiENdUO2l0llvdrO9Q3qXt5dHH3AxRNQR67TPT2ZPN7BMHWvVGT7eSenaLrxiP0f7l5T/
aggeZzURZE0d31VV9bLAGaNqvmc60+nwjYh8dp+21fhaTiY3aM/thTRQs4rbTgpaEyWS6BDDhxbO
YMF6hgsUc0qpTq8K3On04LrMqhXC0ybTz4znUf6aUbDm5tvCaLvdbNhBLsaIx6Gkq0Uhm1XE6y9U
8ovBDFCsc9RYRLDB7oEvnv3Pe8iL+v850rpaVDcc/fRUuhYLPEK3Hy/9W4gRTdL2NNfpJRZtF7pM
L4iknuMumy8XxtQOAaIfbY1wjUuilstwlODVV1YAujUJhMHp9UqciaohC/LZ/1dq7ZpZF2Jd5W+G
aD7VJOsTHB+34sXZtVc69xwYeFOzUCAQtOvxEW/5qKefwX/NlGHUl/NshgnhF15sVgT3l7P1K/OT
0GDdrIhlIldqJuCgPD49HphQsE8eXqSPjxP+MvMjWC9UVRINugtlmPDRrU0yfj6fI9zDZBABxW+X
R3tDJn/tMwR9qJP1pPwzlJA10OImjRANAVTcfeogAQEpyXNyJbBuQocBcJgmm4i6X8ojjEVkJtMn
XHQ3AdyHSQKMqYru3HAJ67mzYovXJ+pqNmL2sQmLD8nr2ZyNCJ5c7FqeboeCJvqLGkRtBAIFEBrk
LseJNf1xN/k+qsOon5pgRGhchEgNdUPhAw6doJ69HOl0ZjZ653Bqp9IyakNHHxrVT7S/qlh/Y843
puavVQ48Kh2MVGy/aphEpyL5lEBCcjrh6ql5yDZqAgKh/e6hoFzXQiWOgv8mi8bKY91ET32tqNgd
oWl8AHqW56Zw9aAd2hCbKzDI0IhJrJsQRn9aMMiE4Q7YsQiKyG4KHY45V3agz/CmSxQWcE7c4l9P
E9Jx24WaRvEuUDgerMd+6sQ4A8zemEnwzKXuIul5jof0j+QNhZ4DOCv7NDBwRMEYfBfbVGSqptgQ
vUFMjbZm3gWBXikPq0S8tm29veJvldFo9ozdd/OBvEmnwbZGcsEZLVCiy7vMybPknxGef1r9Ju2G
jXsZ98GcYtZDyf/BNBYGz5+Xpmwei39tZB2Wjrdb2P2F86tF3l9KgOlPVFgeviT6tdwGQGIjra+0
bg7LKGNOUwzVf/e8E1GJBNEq4iG5GkBhPMmWWIPY5QvYOBQ1iisGW4p0LlFT41avI30EWZN6U27U
ucxnUQM5qD85JU5DZex7nAMTeE+OGAx/5WztvXDJ8lYdY2FaUyVBQ9mNW4/5C9iB1lv7tyE4ohOQ
YuLrzVfplx0ZfGX9LdCQBy9MNRVYelGceRe9BLkVEfOPo4wVSQxvp39Kr7kj6ZG2t7l7hofWO1+E
vYGn0gltB6bToF+AvZvont+D75Sfyjfyeh1Q3VX1dHxRYAKCClEpNlMByxoPohqdnIbVps9vA0V3
NcTb3tm5OjwHUTvr8UnJaVvfcWaLs82cDjE02zUo92SH27vE2r8yLFmJoUwCSgFLRSsStauxWTWs
mXzr94TFggVfOV4ivUnRsZen+tOAaWGt3Ijss5Z2CcSN3eUw5BJbwlxVnk48DDrhDLujBkFkq14X
Y2Lv81lqrByNZj9IYYI77cAq7xW9rI25AxRaxhXyxNHFB/tefEXaJHOA+do9VKywIxepZFvGo80k
A02nL/rpCh74i4IvF4vboLns6+l99hncGbWjY/wfoadaIyMWEBuVO528v8xvru2AZbNZNZh8S3pg
92RwpUu088KEEZGe95Hip2ysUJeQuQk01sNaFBPiA56NWOXnTXQk5y9eQ1mZY5hLYT+YmQwf2zY4
TuTR6kk1jeiHfVe3l8e0hypnOo8eL4jTFFzFytzX7iJePXTb83QdYsfk7uyviGO3ryQyGld+sf5L
ByM6Ezr57QaO9GclQRd5Z4MGetbJ2fajPAQo/1FsKfYkZJMxvyhVAHLimDe+UXPIELdF0yV/k3yO
aBbLvtkGx2dLrbWd7st2iWySVBTXNAO/tdqda6bycO/fK1Ml55oVlsWbygRwZsOl88IVcg66AzLd
+0AYFlNz82dYL1wogElRUhSUJ4XiWm/5ye1qebgYe/99rxcAm75VaMeCT+VEWXoWxQZi1jXdvw2x
QajlLOfK/qQB+T4RsIcdOkSXFNqnwmD9skwnTJVTebbfPCmD49d+1byo2HvCu3zM6i/6zux2IzrY
sO2Z6oLqRmpbCnhhyv188NyRDlPZlSTDtOfRuPVOheZKF40JyQLhCuvzeKSz0Y3Np95HMzwynEUi
zy1VLWi0kCwFcMLQ8dC1GvyEjR0vZ1ZaV0+S629XJ+jNI2MamYPmM10fcZ8bfkSqUsKlvrvbwEiE
0eLJmCnDbQKLGfasf2qjFH22kraru42tlikN8KCumkygAnyIEN65D/ViT2CoHdC3UNFQauECzH43
3TKj0/F8QQvEzxOaYyPAgvB/lg07ygVMPTO8A+vuF00/Yjez3qFnmSmJU1WBN+1KsLwUsjpk2MN2
5cK3VOYOBd/FSJ69PKMN5sJi/KTSoLoqtK7kLPTWfeDgMBPZNEhQXwJACWGlL3ctdrZKguO8ILdJ
2Te2omswF7wfzX+OxBs2lGrTyc6KYP3AZvMfaoyBve/WLnU8/6w7I5+7P4SlANQYWIxWsNAUpzED
W9lR3axG3c0Fopk0JHGUSwL7bCHF35fE0hPIwdfN7NptJcJww7Rc4Q6ItbHQ1XdgNnQHeXoDieUm
wvFUSDuhPs303zDKJXHt2sHVkTJNH6mV+VRa3Muv/tX+UtxiHETsn96niQjxirnYnNe3x/woFISM
mwIDrvZxU/bTIF/T2HMcCYN7wZgYxcSsdAKxUAYfa/radwm/qVPJTNbJbFSuMtR/F7eeFdtpSYau
9buLnnssnmx9gKFzfrOp6uB2TcHUXrzR73raifqqjAaS0uM9qmZV92hrfZNAzIUeX+Vs/46vgI+B
QW8eSJxx/BHdnVtWYBrKC56cOgkcxDDaufvVQT7oyvraN9jppOfp9m58/PTixqSv2SekuliUN9Do
p9WWHquaIhIR5+223hCzva0zKdFmrhqBbqermsQ/E0F0nyFFilByjow3cN3p2OM4psXWtATDf3Yw
LUerpBCLeTJFJtCg1XwoPQrxEoF7LPpS6ShteKa/MIxTyNBa1QAzwov2VjmA/GCVSNHpHH2ru+hC
uHkBt8FPp21C54YZ3qYX8GepGyGc2Ni3d1/+tlJVM612T9AfrQpDWBkrg4nc2WsiBPvUbAkdqy5Q
6BXE9lZLw+aQUutbw8NXMTOlR7LXLdIsNYhMUukYLhWMHchmv04tpkRBWYKDcKvcCLaRHnNoKwEg
KAreopaA7OxezaOzQqSmjZySp6h+rFZZ7crWWfioRDVKiYdKa8EJJ/NUoTva6AvSr4LplCx4P49a
NP/vSJvCA7+clylXVKfoW6cdsOuq+7VDIWrPEhUITxb3f5gVI/oBYdpj00nZ3qymHvQ9kAzQDL0Y
7BhvO1B1jkRQGs5UkGNKFZgoWjq/ynOwaWhWkoIwwgI7KV5O9P/0eOttCHqweM1NLUMR9rRJLj1o
sYE9BgVrgT1MN3Z8V/VN6RjzfZ5nV4EjcZ5V3H5bfF39ajBLdT/Pu2TjcDOHqhb/WbBMLkn/Oye4
sVmPC9eDcBftANz9j+M82kyz4yGzUeeqIvprcB2XmhhW4BpVozVT7QFrchd2R8L+MZ4sUwFh+LiU
VUfzn4/cxpzf++QKhWLq41uVtGsWnnPOHH+rKbs5zf07VB4XUTUJYKnR4wt/dNhULNHj9NTzEQj7
QsruLxcOWFNRjlVD8DLsB1uNIIwzEIQSx5aKxOz01Gk51p3Xfv5p7WbvUUbV6PkqFD5F9roCC294
+9pJgvz86J1QZnYNE+Q7at2e2KYMtK4iFvmIlT016ceqllHqCS4IlA7qT0+2/iFNZ+dB3AsLl5wE
3BiuLk7G3FfaOZhbSxLzwvKKar9ZK2gg0cIIGz33PMwJeLYyNNPznyElMiTv72zCXwT0jkIIv9Fe
tF0ahJmdNHIGYxlse+TNUXT3qZT+Aqn75PP3AIF0Qsja52C1+lAh5hbheX2FbRM3iaDMmw4DPZfW
w5YfWGNG0nNnQD6j3Ds/bukdPQ5CRwge4D2JP/+fCWQmI3G2Qcr94t/ABlkO/+G/n3zJPCy7qTaN
03wYKacvDRoI4etOWopsYpiDcB51m23oNe5Fo4Mf//PksMW52fDlh11HN91e0ntPfsH6HNnAvRj+
3oj+Ju+RF02MVkN4XKrAYAyNJnfUebOY0LVz7XHc+D1DHJS85caAQg1mFW/t64VMeaY81+azUpyz
LhkT15cUh6I7A9n03E6CfQn3Uido2oeL5Hb+xKgU+x3lgO88N21V+O2qE7wdnu9hFtqh4eTV7u72
8R4/D9Av083YAqxkJyzYCZhqCZB8B0RqbP2usoxXAGCxm5epb/mguOQKzxtBrNJXeUhrFCqMYihc
Di0aCLQeGGEMvbE+4fqUNqa7HI7WrqTES2D2MFMLrStVz4NBg7BSVZbjyHvIYiNUJ1m7+3IGcWLo
zdxrX+qi7Z7JLG1/MFILtRr5cU4q31fqvSy6lqJTwI/Hsmz/TUZMHcc1kiMmPNXG5MQXRTQt5jut
nxcAuuuAy+1yVr5l9QjF963UNMu/KkQ+T7MC52yVjUJN4KuW1IxSOHBdBbpMrMip5Q8FJZhM2BWx
WWLn434FEmUZyFJUJ4d7OvxVkd8xBr896j32uFzYrewanQKigqiBG3YU/dGxajpa3HR9CliWFdrB
Ui3cChqqqLpAHEikCku1vhFxW08jUapIbp7ndiVm9HB+YYd3l2tZCqzEnis09saYrmYDMPi1TImF
hBuMKjXWjR00r5303s8cbqvGTV0+HHa8rpKNUffB7tUaEQo8giRG4cRPeWhbmWubwsNnwhhGjgQQ
6zT6bVCVbS04gr0nq5TXnuYGDjvKyqXHCUloOhvrU7WgBqh8QSLfOaGbCIj9RSSeNw/eqZOhM+Pk
cIB/gcqlUecxanytWhqAufVWb8tuevesyTbWR1YzHhmdUDnvcg4wlJe/WYD1cf9fOE8FwdhhrJHE
sct1v8umqpUgLoWIFUIBXm/hf83a7MR8Du3A6SzJpNaCt2tqbb3wJj8W6MrSSXbijGjztqsUJd5y
H+9EY1IouHCNAOoRDjMhYxVwLDPMIObo62ObJ4oiyrHiO20LtBdfbIlLeu8hBx+0uAAQfMCd+sgC
Sb15k4XxLlLzqN5tskn3ltUwWhKRXAlcXlqFuypicYU0Ts0RpeXLqTGD22H5xQ7SQxiGCKMxQGyL
tgHUokDbYjvwdJhJEZmR2A9df0zDeSO/NHL5me7d1nsKEq2dCeNZFQQZmjs/ogyZtXWBrheWfr7a
fOiKK7KVOzLzHle/2LL3pCjqUYjAfTOhFilqA5ATpeoulFiPGJI1nSr5Nx5R4SUGnlpuFmZZnnUs
7NURCtY6YQTYxDbLahVJm7XnHHIRxvYCQPWupwlenzKTV7iLdZli2FPjNg6dhBZJBifSnjzui5Bg
s1Ny5tAjr4OVsHsJaBmAOnsUvBGq0/5LPQq9K2n/npKBIzzMkP6LdStpJd9xZiOmoBjnZJGfRS49
1jj1wV105WZzeE8QBFGC9WQM/21xIOUxImxxtkWwe4zWPVnK1qniOabjnxY5SlF2VNL/6Ln+hcJF
c+tdTr29hxqqzV8NLuxrXpJFpl3VaVT5rI8doKwYhEZSBvFAhaFFAc6/3og8+jtO5/bXWJMcNxN8
XzWE6/qqcj8JcIPdy1HeT00oxU2/2hwuTCxunsTPNY6lj8Xdb9B/NLn2vFdDxmlpyB2MR4nXmUF0
rZntEpq0DQqH6iYdPck/B4i1uwhu45ezVBS1x8X8hiqslkFq75BNNPObdwzUejLyIwB5xD0xrWLr
s86BMWcs/AMF3E0Dp4xpbWa3n34d+wHlLDFOijHPa40ovdvsQUSCD/osxZ5Vw7xRdJbFABn28M7p
D6l8w6SnGjU6an83TQmGu5PBIPuEOXk7DXVf2TWaLKvTQ2r3I53rSJLnTCSPKlk2X0LA8PD96XOI
74jB4Ksfis0digaW2RNzF9OO+5G/EWbFxZCAeFSZm3kOuixT9fq6tCncyWQIiqZ5cu8UJtW8u/p1
AXQlITuo7Naa5ElVqHa0ZVforOLwT9OfU7YJAViFbkb7dOX5gt5uIoVhyyY/sjj8rHsEpcHQ+LTv
iAlvaLURer23+k3DcYe82V60/9TYtA4PMPEgjquP+3vXi3csLNSRnOMluPZc6IM8U2eIrG4eAIdW
C8ixX5/2P0C+lL4QWh8ne/EWtHWxVGfZ58iXK1PZN2lQYvyqqWQzPBfuSMsqxkcNgxMApfIeNlCx
p0ps8SIC/Peb9elc0GTaByujp+vL5f6TyOVAxx7ITKu947Ox/PVafF5ixSLyz7CeVqtasED1gECM
dbGHqFxFX+Fi43RxBaFvmn+TQYjXK4qJO1CDpJwNyyKOqB1PSg9SXAITdcm8/cbFKoAqXZ8rPPgd
kaKHVs6WSakChRtuL2lWKQO+EZnfyT0SnwYdVkoTbPlBVI9Ij0KVLoxMPVOV019LpLyG/V0GCwC2
txoA4HPzpIGzqiz1ooc0UdDx09noPNRkGb1X/saNNY8KMUl0F+gVI/jOyzvkzmclQHCRyse2f0fq
a1ucm9gcuNr0n9oxlRKZsxrASBM6tsDQLFYOXnNqCOV3AqepfS7wVM9o46hS5MfgG2oY78fmZUsf
2aL1qIrQr6d5pxeLCFT8JgEI3fFQ/JhDEBhhV6Wszt8YsOwfv4yXP/tQ8pPsgdpeC/emIcJmrwX0
vXURboLxGfPKFkrrU/opdNKgAE6Y4BUIH0VMc8p2ZE/0owWQycnDU8YTMUxjMskoPv/orQ0rB3b2
qzVMmTA0l/QPUIuWG3IlmPrybuNM1mxbxRo9oVusYtgj+biTldTJT6X1bM+AQhtaZH3R2NEPDpV3
fhgS4d2bipxhNS5+MGj/KfEYvrYBm/qIMK183SD33KAtpRTJx5cb6QJLV0KevRnPlZ7LSPKPx7R9
J7LxJ2cqw4iw9UXiIoJSCNhxy7GdaK+baH8VGFjeEtOlYYP26QFtDBcwptq6anl+tHzeqWEz5IFr
7yH58Cy4Sl9TsN8Xj3isWFb6XwTCHVQCtMm7p1vyoOhp3yfFQda2s6tEqVDU0RJBIF1h2LOEuxr5
724AEZ8c63+83QPunQeAZoXRwi8rqDQGbTNW/jXI1fzRXigatBVT5V9tQwQOeIGbsK7iFSs5oq84
lsjj2IswJndOJA9JyKaIAcrO1d+rqh4cBjMCGffl0TMyPIncPmoA85FYXNvoq+vDqxpa8BUzZdyk
OpR0nA1abD32Kvarhp9POoSstB/h7CwM4Wrzhdyz2PL93+tnwp6u/3oDkLGkyhCWwUeHSY1fO89k
nHd1+w1gD4obA/Qqq0RBB+6GnuZN4GMmQFPJDMrptlo64D+/sOp3R1GupATVrRh4ZE5J+le8fBHs
7S6/W/A21nOHvnVGXswoW7QfL+2V8+2j7DaLMdBgNMexdOkOhMM1QnohKoTG5qQkW9Hs7FmgiKM/
rffzmCfHFzvJLAiK+8sCGscgTwJ6RSM2a+m5nT/OhlT/pfxwA4hD9IKOa5QWxwm0mSmgKfrOA/1F
6Tq/wiBl1iuAa2ibYWzaeCMhecb0vk2z15UotLcmVUexGs0zfMtJOdGyOH4r70RJ/TTjA8IrRANU
znpJeVHuLFd99dLgn4uxRXLCPZ4PDb4qnaGCiFZa+8LoOMc5x2QXIOxiivdXmFaGru7Tqt2cET9E
9auB5m13reCzAIBCyhjsprgWvUBgEhRcciFdg/Z01E5yUHZBpzpVcFu8zOTxeAa3LmhqkAwd3IDT
0hFEF8Oz1cn4pDL9YtQEQmKTAm3G+vjxLiw1Bc9oN1nSYv2UKRoL/ANy/oe79vjkTF1GzBG1gQS1
FMUkXVHs5bsJzhZpYkxntzG59Ielg38MV2qfgzfrS3NJKW5fbU2hTrSY/TEBJ1gJcTxdDPNdHIva
wnFhmjulumNCpoVHx/W79GsUztE1qyhWNbpSHlwj3wK7R7GFnm9+3vv0Qf+yH7wuHCbmB5GS9FNb
cGQtjKrkK5F+sw6v8KQW1FMxY2/pIIvJ/M95VwuNM8dn7JcGC8Uopk4pfyyaF9AXxion/Qh5W6m0
dF14UEtwYKuTmY7Icl+5ivuZJt4n+rZAXgKZf66vqgfifz2qqT/fCqEZjF/68fQg5ihnhTvk/EQa
QKM0862cOasGSTaPE7Gx88gtCoAwI3GbpAgjPDFIsYz6PB7mwYIqYI1TSVz5eWOVog8TBtAF7lto
0bUOfr1Zj4Q4Or6kyVIHPet2ZN3/cdCJr63K44KtWXmaMD/LTfu0JS6L+qrE3D4OLDIy6VfFuA36
275dQybxMgtB9O7mnMRaEVlm+to+WLR5Leh0DD2UCq1WJARKOZCYeS+8NiMVQBa/Gmk7Kiizjox6
QHnsjibx7RHboga/Q6D84/+9fm7lKxRXHLYlr2Cb7ev73K1i66PSAGZWBLg2uDlDSXckGnOOrFxF
YWJlZFbewESeFM9f0895sFBP9Jt/ym+O7qwzIbMXMCiHr8Mjix5828VIdlegYMovqvyq0ZaSND4B
iN6QZxVJmvYy5Gu9RzkYXKWT1JRqsanYNIxocLzbosirGgUCiep+h4hnTsCBxQBslcgjmVC2Nl3t
3sH798ZMxw6wc3kqE5lIgjr/LcsyDhM1QGJls6YxuiUHuQD0NZx2S3rMGP+AhpjNstv3wHw/d2KY
5+3zLcbDfjO97y/74StTl5C3QrV3qiZlDogZ9DYfVXs2sIUSJmDGQZbz3bYFWtxko/JniuG6bDJ2
JUnhrytLxFJgd5kxZ6Xmre9UFpjZ8DgiM9CoXKrVqEBgP+4BkVw1jmbjr+dq2vzKwRVXKqE45SGf
sJ1sB9rQjtj9lTCDTyfFGWKB4SbC1iZPPCLaKM+VE4ezrCyHvCtZatcNxAOms56uZNJ+wv+Qsewh
HL59Dhqk/KlklMlRSWNcyEIop56CRSPXY8duVOCtOmKlreAvgAnbu22ZkWzMSHMVi7PyFDXoSnXl
MhwmbTWYKH/+A5y3dkXwdMek51BCx8nkfEC/IH9jkfgAnKDT4WRfDEgC4WHMHS96PzwuNpW8OX0U
BGVdJWcQaV3FJbrstnWSPr3W/txu9eMeNONlajDAlN6IfvZzBqg3E1q2OIDKX6aAiNS+7LVSaBiN
xYrtmM5l3eGeyttyuPcUX9pVpFwlkC3hsWAninWdtuRpInrmRSGZksRj+N291A+lapSoDe0rOVeQ
FWxdyOTXXkqfEYpAsi2uZ/8mPGFXy/57VAANpOHytopVloO9A3QPTPSvL7jJRPiNSNuYI+Xq95hJ
3NvNPvY5X8askSL1o4kDTj79KY5rGsyY5JizD97tmxwB8IVVy6YMsjYEMY/Wz6LVFG7/puyAaD7w
+Bt+Kzr1M86fVOGe4VdtB/0E+52Bi8vWy4ML8x4x15f+DvFfNPcsIDMYHcFt8vth7X8vl1LDkqIr
7iquh5qI+VKUkEOSGPTghngM6wmDRHTRxulGhPfGD3jl5k/FiDV/97y1+VuEt8Whd4t8cs7S63OV
4Dl10NXiJVmKutkQXVuCzR34msL5yBG9ucVHejjXV6z5LZbqSvVYK3krVNDwIk5U7E+hhfMr3D3c
sKaVW5x0OycN+YSojkh43KkjvRdMTwedO2xLzJXLulp1jzJGwPI2ec6+E69Vcdd/nglfZzcvSmiS
81E6LVRm3nOMDSwH9PuyE1XYNqcR9hoqOGM+Q3i+INVZykUMAMChFcNC89rzR/VrVj0uBZ/l4uJD
dX5sRuJh0NiLx8EApIu7qkqlL9ZFADIsgj7vmNSthaPei3Z+2qrAUMhY1FUvD8zNYk3g82WgOq1Q
nj6MSyLenmC02WTM/A7OIMfwsp8DgAX2ELy6VV7tjUiMgTRuOTNbCqKC8Adfqstc4TASytC6PGOE
C6aE/ReuL6D/OSfEIOy4OElWZuW7p2eLlDF2ftDhZ+8XRAjFxH70Z31rVpKw+zzvYd8dCLg+NREg
FOXYWhfL6iQjVudL6sLJ6o/hmkcr467lPG1VetpJcL1z3Xrm5MJqsBceg8G+paLa/mAY3wd5EYPh
1oSfC8jWkeCYMPhhD9nHttjmzTtD+BfSXbZdWY80XY+UFd4KzACALE0QRTKVCI4teVFN6ZjzlYH6
P0GKqPcil3UQ+u2wJYKauThescm035zGC81iR6zTTEkUM4ke6GH0x00aZEFn+ZN4KzIihVZQWzRs
vHC4wnxmqBqiI++KXL171FYr/XYxlWX4FzOWw3B2c3mxwlgkECVxEZ6SFz5MrJ/TUoaIoJIrujQC
WxG970rAR9EK64L6FzXRV0DhBNMSQIiVxFqLwLjF2HMkBiwBts9XWAKlOX9Ych6GoKPzEI2aYVgq
3fVBGEExzVn2qQqaUeTgKui3kLjULc7tdAJA2mVFvLxgwxm9DuYT72KjZ7SIDPjsYEsvBV8S77KS
LnyoyPxke8NNHDaGUbEPF4xilKaZCsPhsT4+GdSX86IPaAWqC/oc5mNNL4YtftZb+CbIgPupbxme
rJPqh5fsGcdqakLPXTciUYfGcp723j2pkUnFQqkiGp31b8kt5m9nvbbuf9EvUeDr8ubyU0Zdsy6h
sYPh5JfyMrUebA8TgkAHDOokwPYDNTyNQCq7svTKopnzjKx7bPwXvSGvctJis4sskctLmSgEZc1R
Lzo+mWfKJo+LIPRFqAH3fznlJwojT+sRWl3nJtqqHyUQ/zJJh7Ohve7UdKp0TDBeuzCsKZj7sc2O
0NjIjyFE3GPsnGwcMfxzXGhvqiK+t6XzoKl/fDw1bzZq7nOBu4ePZ3b0ZrCxztldMybKIoq3nxXj
UwPXU9HmeeV1R7xzsB6hSDAmLhPVVH82i2vkyu8CaiSwhRkAm6neXO34lW8p9K76wVr6jSwo76Hj
TKrHyKhyb0iZI9CW3XE28TVfyn5zsweF44ACw9pmjBJj8OD1BqrlaSwwb3UEak1ATjX5ohhMWUZC
kauIsqNoOo0VBw6wmeQKoGRKbs4Tu+NZtVKAOlmVug0bw6uMmIJZ72Ha7sC2Fdt5obDPBwRR9Ajo
NzWZV/ObSXxq3f40kSYZqeV9CNUDqyAfM5gCsSvSsvE6IYmrPnCJrJZ/pVgURkMo0plHzq34W4i2
txKlplKfUNqFNX9l9ZQgyMvzzPVK53qv38yMAsR7GHS5V7QYfeDAgw6ATcPYtmOOI/aDqjJI7uVs
xFHsqtORHr1Bqryckb3zr3z5IEbEBqBHf889PPiyefMLYn0uF/eVQTOPR8Scj1gPtuSZEsUblvXP
lB/DMpHVLv0wFQX3pOCXvKBjJlUVlTMZXQCobHRgLuJ5QCt6GMwQTYYWK1fiK5lvUSqp9dRfZYVz
dzbuXNdAZqrbp0Bdtk6D42V0fcgxJOW6DLyaN+SN1vFh/t8/KctpVm0NtX1qwt7Ls0mwrYXaqjdX
gbA3uqjWKKtwQ8qKDeJ83xOfh3dOOYd6Xm0GWhSukzgefKB/QF4VvzAcCgIlqYzqFrUvNwuvjHjp
VKWT3M8c+Mjb6t4S0WP+o4wRarW9Ta0f4sQ5peJ5byvqKaTxhdUt7kky19Iw50C1He48Pwzh3Wsn
vysM8YN/PJX3UR7dXQmpi0KebvIVkzZqNo0bEmB3atRiP5Mde7cyh9LHsTRZ+GYkaNLN07cYjOtH
laDrvBgBcFyAj+fk7XN+xKzvHgCsz3SAR1tso+2iAKM/LnMs9hRFMPsVBlsNq8zHPavLWUEcIoaG
zXpewOLg0AJ9zJ3RGJSvdkvME1Nk+dop3Ef32On6fTUDwCdfuqBm9uSQVxQy3aBCGG8wfkljK+Ol
eI7A0YYgQt/k1rRpqAcBS62XD11omyLfAel83Qp7qJC4LfAMQBQxcd5g9wp+AlLZQRmPbEdFgKdh
K7Y603jEFU+YhNibVDhjuU6Xyf+bqHAMTyMOjHKQzmV7Mn72UO2i0X47hDWfFv1bQOIDV8qblRB3
cvOt4uRB721/Vr3W685LXIHhoMQVL05lJ+MBJoiJmv7Fq+Lrgr3VeD6OShk39KtLzmNL3th4wve5
F11qpw/T62ZIWPW6zemq8iSm3VBDCLgFjwcNw49qz1X4Dz1mPgiC9uv5uY6fb5bL5cLwGCmfe0bg
wef77vD4Xtkx3RIr7DAay7gFt8jnUAHEK1N9xQbKq3hXiyfbD1i6TJ4rLK1mD0F3N6rxE9Y1fxzB
H8q97nGCVnJdOHnQUUJ/AxtnWLLuZDpRaZxhA/9HYIgnKjIy2ibx633jEi8efNJuHXFz/Cw/MnDq
Kozroz8J10aZIQ0MF4cDlWo/Mi18Ra+aqCEDyV2BE5qFMryaV1T9Bppps9fvCCX2B3xb0WE6k3Fd
8md0ODq+O42vXlFOkBLn9hU8eyuRuj6DeiECB9k00dNxmz/2QgG26IEXi0z2kxR7DgN/0p9aEIIv
Q0wGTyohBG6meaF6nUUJK/+Ragqivq+epZ84MIE7YIJp0YzXxGyNo1iDW/Ab7HAvVXZnXAvjx1lx
fzii25EWAm2+MAU9rH4aEIGDtuAlEIFZofHyJ92qCSqS3rEqDf7Pvc4Bjsz1BeI+FA0wDINk8HU4
afqNX5F1gMZGrBO6t/o5nNzlNOU7Z7Un9KfMogZs66BhUpKNE9TXmwt9r7qmcvAT0MYWgLRSYIS4
vq9gayQKJOritrYrgPPf+wl3Su2A+EtSwxzzo4TyEZH7YQl4dyoM6irgaXpQ22b11W/J9Xq6zisj
lJalYg1fnUij9ypTxPQ9uxso24aUnuHqU20jvgjo12OMKvJwg66EZH8lwxcDYLZgkARAcVt0PtXm
0+SwH8HrN8bdZOk/ZLzr1s/tuhGm2vcz1CQRK/tNB0vP7RU/2wIAQhfbaz5F+vEON941KKlMHMKk
Vn0BJA0h5XlS2bDjQM8XdNGh4QUCsKv3hEav8hxRobV2d1otgKhNaeiyuwfenj2Ns3yKs0IiAtRf
bBpU1BUSIVuV6POf27Kiqvz5Jz8txdAyGwbZLZqr9u7CXnH3/XlCrvNULzbMYCSRyjbHHjiG6xEi
rXaZSdCX7MpTVQYbey0jLBuD4u3lAd3wXHZ7s5UGSkqabm/xAW7n6e1vcODSIk7Go8+RTJ84OLt2
JP1zbeW33D+9619WS6iOTEoUHewuZ1e/oOTUQi0rw3WdNNfccrYINXpefSkEbMZxeiQub52xVsmQ
9CWnjQxm8p9lcEHjJwFXHoX/GRcFMeU9wAwzyq2vSTU3rVJLIumuRdOMsWiLa6S4QvbrsPsPkVmN
+4l0GzICr3nGpMUxtyAm12CAQfAvNN9SM5/Lo3BtRJz5XfpitAoUxU06gjuXgRuDI/68gMwzMsya
TDdjgkKlJaRHptAHJPDjyNeQ6nPbAt10G5Drt99Pm60ffhbatLPp1bgecVLSM6l/gK+E8vz1tS3+
zpM9FetRIBNHO/IQQCLkjJ+9SLZGeZ+WhK0FXgHFPB1zqU0hAHjz2st8V/JkLXHizIY/Gh9mn3pF
3Yblw/Uxh058Pvszs/O0PcBRUzJxcUycV1CKv79k52S7Khugv1TwcJEvo9uAxciYahVGDW7CWJC/
xBYRfsszq8r886Zg8tPSgF5P5aM2exmVnHEsNrpft5DYoG4OnCyktK2y5LLOu/VuID8QUIdxZFmO
J630XgXQwaQIMZUOgXhI7kkfOhmGmj8xgHnB3VxWVRev94nFu/bBaP7HKxnfWxyc0RnRGVpsBbk+
2PXf3i995ue6MMEeIOnZr587FRJi3Dztxnd/ImzeoYWzlG9f5/zgXZHD6Bv27A+kP4qwhL/sf4TA
39tS8zkzbWA1vhXIEB3GjxcgKHdNbiOECWHe4b6Yr271DJermMWDKnXMXI0HMjIYiYUY5NNPxOyV
rKikZ5q5R4sDmwyM4btFbQ+EqH4loG9Ljk/8GKR1L2msgl5f8rVF9zPL6sIyqD+UKpAD10OfCHTE
TWK32jtZTcT1MynJBI3TRDtFDudLALmYYvGuPIb2kPuCebuWea0ijjAxdeLWUrdHMI87bpfjSj+l
47IKpDzwCNQLDZqBEGNrQPU3kykV1S7IsZWeObs6xisJUd0hXEJpHQkkMaVPJs0jEtWAkMwkpJm6
qfnwmAlF8XkDtz3CWAoMFYTjfDUPk22t7QLe5SGvi2dqPnQdt8vGcu91hH+uEF5tGHwPKrx5iHPH
+6yD0oWzprX+jm7V3cyvOuAmaR+vHr5fxOoR7u5v79qgkGgY3mMyziWk6TYbLpFiYUyHIGwTQ8WO
q9BAXqg81V8ylti8Kaxoq7FcZ+7L1tUOU/4TrVtFw3HT47M0RNeEYxgWJ5mUXXzKFPRiwBpXyw5C
gnNSZzfOpCc6CmShWTUEpThEq/YHuNprP4RrPI0QnYBMUocoiiPJxE0CUXizs4mdI3dAha4TtYKf
RqSo7A+y27szIIFU0NWY+3TqvJUejyTLRfk4PeQBCDUO1Ce9Pq4V0I8O+raNBt2BXPrjqWGmeGbe
niWjtDjDN+y+TfMRVLJbvYe9NXiqQKJg6e62peaH7UmiBkAC26n3peO5trqb6W8esKaS+8zlnZ6t
sKSAMudxavd+iJHglf9nuIZvuqPW1zNqKAOPSSJ55QcIjPH3PI4BDEfuVayPPrBluuyDOzE5GGfS
1d7cTQjHK3peH73ZmfWaI1YlcFedzHIkMBs5QXX2vkIoyTojSdqn1Ge7AvKm3LBlMDt3qVFYGQup
qepfchB+3z7PrW54HAzH7sX9aqcCy+Su35fH9V3ObkoiZL2gDAxc7P8pfeCOAVszMsau5DDa/4Lh
i2llJAmeXvtMISa8jLdVdoq/CmRaIsJsglCuc1HzgdHM1a2kZhxDG4erYxM2VbofJD00s+yB3InF
fsn4ouWSxzoOJNKpaOgjta5RXILB+nQUXPn1JlZebztRwwKP7zJDqKU/kY3BViQtdLGnnSlj78Kq
C8ogb8Cex4GcwqiTPZ2OS9u2qSjT/LhHiHbg0A1/4xVOSpBsBxAb3sd+YRsgjxLjLu++fa6Dc665
LGew8J8PtZuLSnoJhV5QrM4WVczuFRc4pAW+dL5IHLG21BnsMthzuicm5FRL9pKsmXfHnHHkf2Fr
XKL91Hl85o7HzrMNc0dk2c3nkrWGOUhwdW7tfCb7wFhvoNW2YOjJJuizU8bCmjyH0Rmq81Wpa6Qx
AuhfmjHmNvD/xXFFiRq1CQ8D7ytS5yIrA80Cgj0XRJOJtd8oRo8Z1A+IvK34wc+uGJhADyYyPxVW
5KY8hkqRVVda9lsLZtwx1p5/QNMtfQaEXKTEP8krrRP1Dc8UvAmUdf2nGB+fI7067Hy5xKV9h4vx
qg3vIer5xuwkoFobnzaM5bteVo5Eh7cxhzLOhjGo+qhYOSLre9vhBdx25wo4xnJ8C3V/XrOye3pb
r6k1AnxkN+m88f27Vh3nIgbiD3dMud9dzPfTUbWh/7w5EKlFd9eLATLK+vWXkdslvSHt8PSnjaEV
GV0dNOv5nG36BOMjutY1joCFK0mfrpssc9wOe5qXqvwajVXEv+Z0VPTSfW6vr+5T05DIg2nUCcu9
w8UvskG3SfNDalSAi7ZYer6Q0LkTTHfCYzMv/uLr5rFJH4Gw+fU6r/V0GBD+x5iwYi1ot9E4g5Sp
OEh88OVaRurZDaRXeaksd+/yI1Pbaq143UPL4W5T+bdlD+JYWUMe4o2IzncfUaQ39TkjE01TE5gp
bNJ0EoyXahI0TLvAs93A/SgRoSOZWpocc0MCbz5mxXaqMRbO3ChnDWkQKZU4SUxloCjqAMcYFM2M
gO7jERxnTY5n3bOlIy43nuU1KBnhp/SWvnrN3ICLz5xrYEWByxzQzxINxqKId8+ZdILR/OHdetF3
wWxYlzeLfn/OEhmwQburGwUpXSAUKYAyqtdDq9Ue26lkXIgak92EuyPrlY1tAZP49EqXaqzXNoDu
pQNJOfr/JsRunObFPcrAII/fhROSoMx8zg7gQalWQr/31HiFphVjL4qBs2nAnftv7sytrcnCz59p
Aif+lJdUxtWvnTgb33cT+pYaV/1YWH+qBfv9bIxo29ZS4yt6r0jE2GYbd2Y8WuIRm9tDRcgRfZkG
a9eLginucAImb4ejsfibcp6wP6kVmw8Qb5Y8t0lsz0Am8JZe5xsPSqzi7zNN6oye0GcV/9daM94s
eGzEemuE+v9PSP8GaRuQRXky6wHk5uLvQ0vhu7Dks4hgORI9LyKQRvaMHYIVGohDyuKrVr6SMqif
2TwtIQ1MhuFSg8F8YO34HW1o06AgVOknrJdyGAJLYnkGMBpENoDHUTc5UCwAxg+I26pvKwtn/a20
oDrUcsgJKow8XpYfYwsviIyPRM5JMKtmMSxjsN1ce5Xe07ruxjsy/5d52Xwrg8lrrj4SZzI5GxKE
w5/EkuiTe/NSsQMqx+9pNNmtXm42oEET1pZvVh/pUMMbsosLf9ZesdFQ85HAy7HPPEaXdRV32K9P
/JNtxOtAteIO4dotTxW2bgZr/IIJm97ke/Uli+kXd9N4v3/KZABUGsv5CewY5nJg0OTb0erQCubY
d33mkvy698zPG0VFU6fDlT8qlg6PwsRAQKLUvC3de8oTgzzbDbwkR/tUoyZD9AfyGtHad4MjQAo4
qBZgSH/WGdhNzt+jFAVDkbIx0zMPQA2h37vJ2hq9ZB1XI86zOLOz8bNi0N8YmRlZF/7l8tl4Grgb
mXVz4OX1yKOkE5yOneFxvcbdJpugZHdUtyZeseeb/N218fUp+XiHOyXkPNzkn9sMxtgsrXLOHZYP
RlfWI/noVaUFtpz4bdb22F2GP/D63/MMaY0BZmLCJsevmrFuY394Cc6XRoX+kj51fiaLFVM6H8Yx
02mo6sp6CyKmWyrOGdnsGRcTdGFHcrkYcANil0/f2nz3A5fyH3EjzqDsWGOE5pS9W7gC0QN6J0Su
w5mYRLJEI0jNaxrOdlGMgmqdKCMhsvHDoROSLDIUNUlAGn8+ay+3cp+KZSftmnvxjyXEDNV3J12z
F5Fr4QnkHBQ2zE070ieThlqRrvTkOZpbxArZ1SALwYhZBCWW8F35pRL1bggkukWGlg4uRQPh6tjY
RVOgFaeJkRghej9Buysoo8DMglb2eAgzRfe7VffJDMiBgF/mAu8qmiqSSxgmi0Q4s+llGhTqXbJ5
wgQgr5i8OUtI/PkSbKW9a8Weh5erv1FFnAI+X4ViFasZ7K+HU13NJPiOh6FipDftpg90DGwzE8Ux
6TY696ClXEEVWt3Y1zkLJtSk+fIlG4D1GOaOv534bwjBwPgUGyOyBZ4EEo1o39zNG3epanHxKTeG
8kmBEATs7KOotUcypaK9AVNXCl86BKOSqrch2GoNcA8LF/1sGXoYmJV/s+tDjAHI2St6UMGdgF2A
5YbL1JnNGPvH9K0Z6hVv82sxGOTZxAdA8nIicYZ3uKJMdrnMauuDWn+RghrGE0+pTBBMyQcLKhkB
ceTDVZBcTiQwIvqFb4ol6R2tqeoTPqX50SHo4tfNj9C2pujRiWOf1zSBm3JHKxLdMKO63B4GFJKy
OFZzmXGOlVcgZeTVQcLIYcnbE4cCRaHqxgHugvLFejbVlbvbYoMIr8G9rX+W6wa5dAyTNbiUJA8h
0DqqXlDp+8xg2vb/crvw+f02Ps4Am//Uh/5N0SDDtWIDzTTzxbumwHowH+RnSElIMjvF0CFbWABF
cgw0LUQH8eysJ435p/77E9fFvJL/6uFZhwRFU4aW77l13aPRI923Ly/mCzxsoQUSxd/NoRxi+98J
rRtMN8ncyqAubp5Didf0DrkTxKYkbrF5rDv4B9kU03ikvg+r/00MH05qpMhW0JCEP0DVXnVpD7MV
9PCzXgLDqC93AsTWPcZw6j2unedMm5zZupU2sfrSDefM1D//XuPM+46shUrctkO/pLOV+HN3ddCE
q4FsG8DjSZL7WzRLaiSHZE43X+qpsrxrslViTsC79NGAsxng5lN2C7+TiMhradA4xDlVnYYJX3GQ
xaQI+nDK814JXaZGmvPY6UoiC0I9lSM/hDMCAYCVkfVLcv1iYR4+zzkYxqkuaPrCeabQVbnmDZob
miQGT+gjGOwiuTpTlw7SbKnBOzC3AXaxF7cZJMwo58wBmouGu3QhgPbNzDOeXN99iB0w4UzTUYbS
VYOjlxX/hwntTyG1am4wqI9+CYJHBfUey4x0sy30D/gUvKlN5SgQCiMY78/V+h8u7DJv9DW2DCXc
x7RiE4snBB6goMmRX70/S9mx/h99GFRloYDAzoAeeIxAVOUMClU3B+M9cPPGdAQSc1W8Nj+On/+7
+WKnIEO53XpKXlLMAAFAwt9ZXw+hmTCZBEOVJhcjb9KYHYIP1ISxUAvL4ATWcH3s30Ea5haciljv
Scptp5Ox+JRkXPJwM2KpsqTGdpfNq3tYRRVM+H016S3fC4bx6rjeWKVHaUyqLt9wN3At1p4zoPI8
sW9MVe1dyTq0EkoFscUwe1DfQscwWubIeEf4L4Lm9CmXyjjwx1cr3R9kNK+O/KNWE4B6HLq7XKer
PV0XLN9nW3IZUjcbFldgNJtmPfvw84i9JWIV/H4pa7fppXymOVI6lB/AsAKZ8owwd+Kqob6XfIA4
skXL2nzPhH9/mhibiYB7ko58lXs1o2q+bcABr5whUzHTqWcu2ZsOkLxH6nzgCAfLwffYN6atx9/T
j8LTk70Qxzc7tv0KzPhTuDLIt+zY+K2b8Rtqq+zhnDOFYsJdUjZxrIwZA2OuiV9AKsNW42HjLtho
8i736+KD8fReNL2BN3zQNKFEZ8gW5RcMHJCEUte6A4fFLhkrmOawkNm0a2soUtVTYO2zwIWY5QLJ
vpZd6KKqi73vxWy/4D3Z5ZfZ0Imia9KuPDqlEaU/hswX3kQ4nUvx48FpYTyrtX53iw7gUIkofKSe
2cfSQZMHuYXOg4qLhsqoc3A2QRpOmhYD4buztTtyTQYIBwCMuVzowH5qId7hYUUnxgCzaRPBSgCo
B3jRRBTf+zdqaRxY9Imh0arOxYen93ygO216pCCF3K11+quVh/unoMBoDqXO5wmU9/tD97qTXR+D
2g02ucHIg7cthIqOKkEbdrBajQF5gpdYIu8JqpSF01/21QxiJY5TI02lIvU9LfwwReB39867Zzmc
UrdWqdQha/CFOSdJLqKe+0HFD/NrGkorzTzddNQ+UQzuAvDZNSPyUK3PjrT54AsI7I6uaJt6eruc
jpvpRkCJrx7vdhx8Jb99Fq8b4Pu50UuIaZT+7MQGNxxSW9pvZdjzvXiBKo0yUBsz2JE+id34H7m8
BvsIVKmfzWH2DLKEeibaFQvfCWna+stFX5FrHZYaIaiymiFgDQzVNPzIghwhmGE6HsGt4PI7AJC0
SiMOXFyBpr/Ms6r0JIZCWeQ7xGZH/0+AajKy+F48cBvgAIirRnXGotLQvj2adiYqMuLbnknTLlv1
Nn20DmoTD8TVqX6qhZlX0j0r2FJ0NR3rcxQYywMDAnoFy8P30A0AJKNsYl536UPaWHQ/zItth7+A
nZ8xLKeWtLAzYsR2ShbN2fKQ1veoHTp2Y1Kt7YAHTECcIF2Isf7AJwKcpfxA4qdEIfA2PDJxI1Dn
ZSlOMBmxrFSPMRyXexDkxuFj1qPUAypyREiubhLYQ+BWWnKuZwvIXme+aE9UqZK99fDmtna7+P/3
x5gE/w8fGChuvWjieBPVsOMaMlZPs2oDHsB9R4tDPCfOt90N8hPeLuTGFoRNiKaqjVy4tIlCXYxu
N4t73+S/tzcLMSqHmlVyUHj9LSwTp6+iti2LfBcLKbn8BxmxvH0IwFyFzH8dXGN2ctCSCO2lW3x9
OMcPBHWMM9EPxcbvZbdmudZvB3nQrDIsia8wdk4T19OlcmAAwrTgrhadzFYKTifA4XWzwY3H1h1R
3kK3tsdyKflWQ0OJ+IVAzES5j37WigdWSo6jV8mRzLEAJ6tywb5BHaRgqNPp6hWRzsg92BUTKLOj
LfHITpdEAOczwW/bInP+P6HRbVLMwZNi/ZXfaGTc2Z1ClCcMOOnVyHs6r4BQUKtr9cZ/bgLlfsXt
VX3rZgwb2Gvk95z6e3/ryB9veVIMxSxvn+L+5T/V25HiT7+MA4mLB3XoI42UyX7B7U7Dx9UranwV
uD5bkawJixqMZoycZiXiXOvpEDYH04NRei+TsdLj5jzLXffY6MerwkcMxj6w9USkABjMu3ljthYs
GYHrM4iDJbQwW9ykzfgqbVsiTFs4oQ677afVV0ps8Cc6c05qm/okPXyPQL2jjnCp2g0tyEt2mMNr
IGEL0pem9dOiMj9tPkSzbB/XH5j+0tuvPGnfI5mwYmXSf+ICOzu+OQWox+0u9xse3FvfxwM4mtev
3HPFdJfEITem2qnHv4sTDMLmD9SsI89FjaSQxkjQUNcHT5XvYwLqzxrnvlSNfpbYjO3dw9c3XDs6
WzVf0QTD0mcomO6jfJbcOT8iGS/khSCK16jCOzv5q7VQtPThO1xhDtZu0Pm0Jnf+T8Lkxl7KdH1a
DgWR+iAtrIY2ZfO1GLOBz9iTDp2pTowqB8S8N3wpSktcqHjfFoZ2vrLrauKer9ieo2n/kKy8fg+k
wGcowk8TpLKwh0ddOELElqVH0BJ7CtD+Y/n4h6+YQ2lNBtn3f3063Uc3ORabCLCnQ/zJAEY5MCF1
2tYA2MiwjiO/7CjI37LyGxV+sQAL+35uJi3KOoMCSNdRNclMQUTtCGwMCKh0vq2bGXWvm+NsILoT
8zUlHS78nHbhEhsWfQN6Qnlwg9piFZ1p5cdKy0q6+HlhRAXXlXtlXye0EPzUcgWcPI3VUpons/PP
+hmS4HxG5sEDFgWsMikZ9B7SUgY00bllFTXAnQpy/z6kzXu5PqD3Tw8YSIXOKX8v2AKPgYpwPCi0
apbA7LUFPIUfUR8OwyImA30KMfGySea8w7CpuGMH0MT3COK8LuaNsTau9FcGsfQb6lc9SxKVIk/H
EFfGLFcs/yRqmEwZHm8t0eC8WUBf5C1YzO8g0xcOxuBCozR0hUUJLZuy2Xcg/Y2/V9LMkFv7hXBV
7Vs9k8+gOB5O+tLaoe5nSmziKkJehffEb6PiHVbKLHechVXiOmmdiKXC1DYvdPwuLqXn1Vrymnmy
Oxx7OebQKsJxALIc8MFzOuH4Q2pgVhEQ2MhXuE48ktvjOkrf+riLvo/DdwaxCPFXkt+6Tys7pYgJ
aeZhzOXkRaer/965v/3+OHo2Kis2e1xJTiMvUODIHc4nPWdmh2IQrD3wgufCx3DIhFX3DIBqYJD5
Jtff3wx9cN8pBB4uGH13a1yGv7UtBqbCy9+bDid4XWBw6KU2/J5sdR32rh/XdygDOmq0Nq2RvNLD
3cFidNIbfhTlCy6qoeGxSoLiUNOgKj4atPpJ/iA7TXisfjYukGEgZc/esiFxCHazm32b/kkmXIVg
a39jkXvdhvDV8j1K6eV7uhxr5lmEIcuuHSTBMzUJCCZTJYBVAUvgqGiCYMtzwrTr0TxuieifuxyX
1M9yax0xzr+QBjIHMqT+diPAWwMKl1To0tVE2mtZTynoBtHDUISLccTC/ZGkvSCUH9B7HaP2DDcV
j8RawHO2vjfXCmaKQRmwxgC1SbhXsPZsZU4bUmWcjQUDOTxZbqj2amdLMSc/DkwJFslT/HdfjZzB
F6j2L04XHLqMjHRYQCwtJcXuoB6QoO5F+lryrS4+/Nmq+eppmHpyBRwYrrEITDBvXn2KhjbK7zV+
nxxGqka+qV4a2/srhLlcKx9XKErTI8n8f9kdnYzXBErRn8bgMYNpJ0n5YGoZraS9DZlmoqVc+FA2
1FLa7ycSKTjSI78HjfzVVP8F44xuBWCIpYxkvBxGj06+x6p+o8IgCR6Io9h9fEgThBrQsA1VVsGG
Nw9cg8RHh/KxcMLdd3X9To3yGClYTt+1FvrIEoREytblKxigfcYp8XkNY9x4KGc+RmrMnrkupCrF
IZSlR2XH8yXGKpQtfaeJKSArH7Cz6XpRSnGW6mV9zv2+HFO1EOrUAmPoXkDwNV+V1salTZtqac4b
1GnnWdMlYsXx0cN4Sj+pBzQOJCDcxZXSvZqmdzjGcFmy+W00SYZcfHTbvND2rO1GnIM56f5OaRz8
PDeOsEJmGYGcol5ErvON9UAvu1HsgWgZHFefaVMjUs5T/WyCBDzbj3K8GODSdWahAjhP0Dbt58gC
lreV3rcIO0Dn14BSAIXyVFTUq2fCgq0ZJpnyccyLFjbQbQwzPlgTBIf51WKaupU/lv0PStZyDBS5
OZ+MowVOJ2AYs43hEolD8SKPWOnBiSI/Ie2GNnWp9t/XUHJE8LrbyoKvzufid72j+im9H8QcQhDW
XP8L0u7wkXW5DTBDz+2v35PzuoTv0lwvSoUhTx9f8flb3WcckwFBxxYP2QQHzc4oFvfqUU2zgpS+
iQW92xRkQMfYj/LmJLK20YopOTnfxT8H6LbnzntdO2O1yqL2Bf1DWJoxeDdtyE/L9c4UhDJmkBTb
D4A6/4W8RQWc1827cHlo3EDokM2cxsdVT1Cu73GOzAsr3wIvMfIRbX7m004BifK9jhBVJdtqgN9L
uv4kZ+QeXqvKJxp45zssp1r3YDTKt3oKgV9jOI+0xgC/VdDbUmGi80I5qIsnhvj6T8j4DqImjco0
ZSMSyrvk7GfntQbyWS8tbyttUC8GLlJObulGlVYTWG6GhB9gNK8wGXV3epFI66HhtpglApfyJKgh
LSV2ske2xI8hOA+to/PTmOvRu36WPVgHVzG79NM7xLE3EcPdjed2tE7yTM2P1PcsH5r4n8ZETfMq
dqmvuXpmVbIZUwU+131StRneaSJVcRLkeIeDhcvSAOebfn0obF2DbG4skf2k1oRRX29UZ25zgXqV
0zjHSp7l/Np/0cCwQTPvHWcLj++xto1WCBCP+TG7Rw/uLoSrushm3VhhHFi+etaJFWzLubIHGCKa
JRr5lN5k2aQitN4n8JLYctJ6LERQlfYBphExeeCVQMnv+oH2UGo0p71Ku8jDyGobqfmBS0lzWkCZ
AjmYSxAV4f8rxIf9mh64nb5lgVQRwSJreCgHWJq1v9GYKlv/tQw/cTHS/WB22noQkKFhUH82ZvGd
wSkcHARk7y7XgyeFc1QsiLme8jrsLqN+LxgJd7K4ZO1k3DnuHy2tbAMqlKNGHaj+gsxwyjudNLNu
c7K+l8xhiPw9hWpVE83YhH2J71x9lxEBcoWK99SUI3v/jnKYYmgWcp+iJ8YS2daIGb0Z2ZZLWF7J
cWVCfJ4s0djRM1emTsslWUKmBF3oRr4QP5/pbDPfoj+JllTg8GG7CGE/imU6sKmo9QmL3yRn/ykc
VV9u1txWLG1GCehP36HbkOYX1Rl55iGRtwjl4J4eSjdyWNG985SvyS7W+hKgPZmEkQNWXmEPSD0b
vUVozCP3QHkbPJMzJA4kWGL5uk/a7frOupvR2W+qRjKLdFi5uJ5TMgGjPsMhBiGJIqBZkVpZKZOi
YcOIvw6asz7nG6JpFLPtLLp0KwTEQQEuCMF1W7d8MKjzEezY4FXv9nwLbiyjdNaXx33n85Pk4IPB
LNziIDuwkio2PCMAt8O0vYGsyls+Ors/4hKdIeynDq7/x/MdwlWlBZ9Gj0Suddutd9oC4CDPbesa
OQY5yC3MZrthBihuoYOfClEVURTgLj50cQ8BumcCWQdp89SpHVvEwp/qPMq5zEwpM+fNqblLQpio
ZOgEB7NLfv9ahG3/Eik5WdNw+aeETcUWjEGFmb+6NjNnld2QAbqbuNOT0oLFKoRta7hmlPgyGHzd
Cvy2ZbFN8FZ7QQCIdNVR8N9GoDyYIBeNM9nVGIPrVGccRlf05ZvNBnoIc8opirCGaPx3WVUI0ZR1
6u/Qf1xGuFkj/HELMMuQlyO9XajCH+TvQJlSfEUN/slVsr+rklwmHdrQQgC+kUUAnIRtpam/1qL6
eYBl5ItcPzaR5jmRju63TW+UUALp33yS/P5l+XNeiRCcZlk3kE9S87n/SPVtaWZMpJzXAPAcFDES
GYYvokwS1SyXMrehaJbkVpMOUd3LQaxaE2Iw8KJ6UGvxSAsbS5rJKuhHpwWU6LEri98oqbNf19DJ
Utr/+vuaeI+dizH2sWRAeW6G87nFYm4klDuwLWVlQ6g+V0nSl6mCC7/IMsFbjQ8UvF5yzWMszk8+
rWuho2sWIYp9Hj0l2Kp2t9pHN6/Ra4HMF/S8fM+o2uMnabByRcXuSCj5pzC8lkE5nOhYO9Hx0FkB
lJ+Tiqys7O/YOm/SNI8uuiZlZnd3AhwqL3/PddpStfLvorrgrEkaJtNBGz2Zn2yCl8tvkd75I6SK
8gtr18jtQSSZAfHV6tFMDgogPNuYBOqsCbdFyI2wninYv+OdYT8rur7UhRZpgbUfhPpQpWVR04FS
5W1q3jH4SJ3X2KcIA7XnB9+RB6lhQEhoXdD+ucrzIcJc5fPOOnDHiuHF2wLnPeZnsUZ04oVY4j7K
oqRYQ7mRfJPqVTAKaL6sdFemJxeX/K3931szntMffKTghJ4hfSFSeRN57UIZeEbRyyDDP6XgFJEg
DsLuzoWFxxmRUTbnU91NkSUxZotnAYKpOp+qFhvuXO7RDAqU3P5rkC2Zp0hMQqWnDkzl7SM4Orlj
02RcVD7JToSlZuQ+uhroI5m/9dh0K+WH9N8+0WW6h1xvfMo/7Oi6Burbtc3B1+uznK/KWoDLJIzd
wBycl9hMWEBUGiBSdGMiwRgTYav60LUQuh1xV97wiumFOG3BqehvlOwCtUzutMXqkPaSyan188FD
mFcxRT1stvYYek+mIFMF4CcbPTe42/BOpVwdMzHV6/43BwcPERvNNMNxIKgWfNVDWaDM1YBdDvHQ
a/FtD0tmeYePQGr1yHzceAD+lF2+/ByrW1yRU5W2sSQyakhOn9GjNc/ajosn/B/7LPKodLmrmf9b
MfWzaQ8rF5FPn3W9dq/UsCjW0sJAnzklavlOI5d4QAkF0DOF6me5Xjh6OPKFl4s9kmKhaZ17kp9h
baq7oW2rObwgPH2ZAKLdISPSJVQQnPbtHx4634xe0WKakuIQ+WusdgV1gV/9Om54jp0g5wk2fc9J
6X8U5T+XEZb/i1dnF52hSqNHBlmfhF7mTQzXNRPcZgQhCL23F/LYPI1FAvXolJO1cRDHM89ejO66
/KM66Bj6Mq4fLOqF5GGMVsGrhYpSZWBuTzjlV3ofLDANnvixgeopBKLp+4+ZUgOJtz4abLE1vYkl
QWfU2kN+wJoJh4BV4OHGYWSmmCbE7ClR78mMoAN16xjJ2drww3MYtN6kSGOo4XydDxR0aarH1XpH
vEO+Gsh0s/t5ud6nclUzTCqwNlbHan5urAofulOwGMvoxPXu+4LFK3GFXxZXd8cC1IQNrxq5QrR1
LxD78xQWMc7lRstlw6SzrXZyi0RT+m0wk1uZgfIEgEzQzzpkesH8tOAqV4nhQPScjokglwJg4mo7
/VL3oabgPBtdTXTuACvcHwFeyk2ra9cP2CXCSaWDv3AHUZ9yWfqSjxv/bqNCNA/ynSQavM/y2vrl
+bLVyfDhoVC7gkb/UlwsyzzzsIeickQgq6d888aVkaSymM++5Lr3lxDjwGhO+WLiVo76FMuVf3Hw
+hZTHti+kTZlNpYugDjalShCcKRda1eAP2sjLAp8X3u6Gk4miqwe50MMENQ11hEwciXpSF2GVbYj
YaMLKpUp8JQwA6PXoWt0uaoOMaxWbXgCUpu6nSen1JEKVGGw48sFXJtiRmn8mg2b+fuoAD0y746Q
hN0KpqYIGiZXoTJ8V6s9RszRz3AD6BUQ0VZmcGPyJAI7FORVEWiRtS4g0MwCWGYoHs5dCXPicmMT
hnMDE+7jxC2U1OVO/yOusPLvVhJuEX6ePEn6rtTjmw7qRG2i/anHdiJmW13cilfMgeHh5pXYhxS/
2IStrIioPTuEXeIL82YbPy/ViAijJ/PjAIpT7mA2ANF1V+jP2rbjFf0uk47mCxN0fYGhv76GM7Vy
Jdp1Lx6BD6OMD6BnebZM/6XapZ/6PW00TjZkZQ54tQ6JYcxDXqTnqSkxxypOW/JTP0yztYxlwrSi
97Vsr2UIbAA1ZmnredyCB9dbOQ0UGhvI0N8O0jGpKZhpPjUsDfLlCvORRYHwnTSzLxnP57FYIXVE
Jeg9zcvsLADv0PWCoZf0m6Evck6MDiS4qasT01RKf6Ud2hQRCacI2FAqVpDgJnmc+Tn3IptYnJTg
BB3CX3QTecTvdcjZO6opfbTAOqmlhlNtPjYVpY5b7vSh3ZFF7/Nqql7rZIcAHs15wNJLiYufHH2h
rCtoJ8ncWDapJMyoJHcxuEfVe6/Hp0zAF5ihzj1hjxx3cc1pRGGlp2BSVl0Go7VUV/nsE9zKaSOi
YRFnbLGNtiBRhL9jVRqbgyipXdVUuP4+znq/q2hsIVEMKooN0Dxl5MkU/fvpWjJdzTls0d//bmyD
q30tohLHP5Sb0DlwJWM5pfJGm4JeIo+d4Re/7btD2KtGxn+uVJBjK0fsgiWfjBfuEBtkxg0Nmkyw
9togcJ1ugHvt+0Czgi802XiALDafGHv4BdW21Z8EgRb3WwLkTXx+QYR8hoCC1Xjp8P4Qvm9hsDU3
Ds9TB3Q/7yx5CEzYW5qtjFAr5CfSY5L+g4QVMdJJLvaTfzNpbAOB5cxxtWA48CRjMG9gPFCryQgc
6dTNGeiSyTOD26wIJjzj6oUgSBcQzOoknPex+BhGVLSMFpCgtAyzO17yjR4vUEHQ2RhWJpjBdyGm
Tj3QJX3qznVUsEdVRlgv+w0Sd/5FqaNoBu2Rhjc9xC6sxwcfk+IXkDyOftTvfmlsEk4eO7UMloAr
emt7yQTavkLD/bG+W4b8DkQwgAan1m1ARHlBY+7EUY3Sn7vzPcoS0CP4heobeAlA9sAkL6Gacgzn
0hEnxZxFgov3IpDCHR5sB660QP84pPGs9Ns+SCJkly0i1gDhZZLXu4D8OaVDKZBxK9MEjQ1Oea7I
IqLnK+VZDMBUhL3zXC1wzqdZa5lSBnYq0PY4vsFndfVGVKDguGOiIySIh00OQAP2XfkK/xK+Qq+B
4xIBs9o0a1g1G9yoeeli/hP65ip/9YlrLi8YbqgT7SYWfgIx2tu2eA7yAZjnJgKfilAlxrIEVaAV
XNhDOZzfoU6PolkVCwkyiKB8IS32yNL/krNqTxfyi533quqJOcdMuDgtlqwzphpwdamoXBlDxZYT
zJ7OaoXUm2wp3f1rgHe7w8aKiZS1fDYB5VAwk56+NMgEdNe2cd/oPL1hah5+Cpwrzoyu1wIkp3Xa
rbGeFe4jvzKLlU/cbXlGwroOHRABvDpv83X3df6u7Kh3VsF/nuEDZBpbJVDtcO74XYN71K25XQxm
uhYM+XVahZoLkWg+L5H9w+ptCI7etf5qWn3JSQqUQK+Ss6xRbz/kpvZ7RaFB83BXU62qZ5zU+wKd
A4pLQMGVlUordd4zHjNVM5d6zzIVNUVf1PLJodfiGksqwlYh6OIKyiWcSn7R/j8SU9z/Ii6Yxd1P
MD0se3xLzi1bJEFT7zepX6sclwhCDamp0ZEEabnEAfPbRstw31g1DpRpUVo85I/VDmPPOEJkjdpz
6hLtvksuraLqFGzjb2YbKgxXcPJSJn4Bk2/6vvCMEIhC/hkW5F+y0DFIksLz9JKF1ZwwdMZU/nqa
b7Jax7SpK+jP518RAFyNVkseYprATKpVUWQUxpFSaQbyNRQXiTe0bnGm1IcRLyUwv7qHoUmLFcuf
QDGguVJFIYGbtmW/DiCBydL4VFZDJgD9RjCeft4xwcHn1CD5AxW5f06/4MoITgKg5Od6FlfxO1u0
lZnC9L9QfKcXgsg+5A6smkP/tybwv9G7JhDrNjBu/k0Yy2UBj090HpmD7CaM3PNLrUcOU6hvJykS
/3dzQWzHCTc9BSW0l8Ax9BHNXPP7v+PAlmG1WuNRnbkTrs152ST31upYME18KFRm/O8Me36MibdP
HmnOB3m2OvI5ieU8ocDSgXT6DDXQlt+7CsIR8LortFufOkBf7r7hQllMbRyz+fK067mtj/0MWym4
g6zCXsPNlBjFEqEAauhxduvEGX+A6GmWaxDn18T7H55BvWEewTQfz40/dxFiqH16/3vQZCwIdXRp
e3uMYfhWT3BntSHGoHIiYnh5/YFIA4TGp7XpctLTrJmnRLx2r37lwNFWZx0wHMSZINhXtrRArlZT
l7diBghwJTtJwx/2BAuf9mr+EGOONbKeG/WmPHrx+drSWxR8v9gcGpXh3Dv+qWa1Npg8sUSQqaXl
qDrZgdVTuPkIX+LA4k/AJrMjG3/shk1ascMkDZwRZd0aS/j6ckFuZ/Qr4bvTg0eXVaddaIZKZAUH
d8MA6w6mmaZey6+hSOwNo+2OMLzrKLyMXDFLQexXaY7HdGnwVsvmuLgRXCzs5bBORXODwADgku0U
CFHSk+tq1HprDGQBJVvqrG8NHJwWKOoW35aSCuFD9DeC67gDMVZt9H68t9KJ8xP/ZviQc1e7tb9v
viZHFCLL4mWgXG7tJKwfQfgoQ7sk0jk8bHE/gIdRHG7PzGoyVD3U9Y9h3bsF0C5fjj5j2Bx0fMa9
jZaK6N9ZUOO85+zgPOf7Dx9n6EVH/I5z/wl4L/MbdEmAq7rzs1HO3KR/MRbgSb9ZFbW2i7HRg8Qf
v7g8Xagpu32yy3YwxzwChRrsHDkDWw9BbYAJfuqSdaWg1KCyH9M6HNMjrI8vWdSdZa/e2fOG9SfG
nXLmmpxCgh2MMK17YD4/CG9h0O1kg444+KJ3w/9/FqToSI/LHIK6i5VhcipTN/Ko/3iFH8w9pcPf
3CKO69a8o3M+YXmDRnrltFwyBkggDxYSDtoWbQPkj8oMs+Mbx3thu0que/cx+IcRP7RpO/gSvZpF
hk2okciZeEVZvjZYjnFvNbny7cEFyH10y8oe3DAhWdqRqwcBG1Tg0Na9PdJlGv4Kt+7c6RHwT+Ln
8A0vEUzGXNgvpCKChenM83PRtQPtg8XwGp4eK+k8+g4SC+flFfB7HpycaW/dHXJkP0zhDelLmODd
Zy9OW7QA44pViQSqWk+qB0ibrVdkcE67eQh/t5POMkLYTxZwm+Q6XRwKHvKLeBJMvJAmIuWFfps2
QnSyJUdpoZu4f1GlTLOftKFpnRzQD9GTD6s6DqACNpGfSfFI1gSXYcl062qjdySMej2CNL1u8DND
p7pRNVYEkh4FOCi4zMZ+ONiaO+qdG1JuGhxp7ys36CVx3NKB2JbnciqPK52gorGRmqpy8vio3e8p
PjCwZYbbHpAQXQ3BL467VOA7VyduOUw9Tsn0zQuvJwMsHch5ghPUXUQFFJckumguiIPYx5NmoblR
jE94antcX/PHpHEg0nNFjdBFRC7UoWMzA2kTLrKY3Cy2GLOKoQ6TTz/QGMh9Cba4VjWaJxmcafFS
dsQkSvqJ1u/4lAuifM+KhoujqQuRycpkbx9Csr6GY3hv1lQhO+v1iNILXGBIKCAjzaGm8ULEcm7/
9DNAxSok8VFlOF9mt0XAm+Dx0JOndB2tOOp8YwPSRJwtyFYEbP9LeMItUWBLIy8PWydFD19I+24V
oYyPMP/PfCVkT545YWMGVCtrHGPuJMEPYuPfT1900a9Ih7/u4m4UBNm0WBsI8Ly6vbzIgg8/zbjA
/2BabOjEKZngXH3f9PX/kHyqO6ysQsuHbsS28Kjb/nB9mFHxCKZaO7618tNrfTxR5JCHocBhA/Ps
V1zA3GIzfRdYrl+pANYVNZMx77/ChqdlUdvIze9SxJZXeNijrWC22wJwptUyynlVEbcYpHnXegxU
hfrZrr2nKU6IB7EpDwT5qiiAIJJVSb3whsOs1xUjsAYpwxVSVYmrqEPWGWevzDx3hRVW/5HkNj66
Dv4HzPFjqCgPreNMnJAYGF0inegNDPyLVGixSC4QK5VFFqC3DUE5egMsbIBUom2NdpAh3DdwhPZb
ColgZz1ha+7WcZNPUu3Zcxy3KT2Uadr1703YIxVjyXey1IEKtDsjDL989+F8GzPPx0LliBVX5vbJ
8Jfol+WnpUE/eogTNJeI5MJm2V+nE2wmNm3fOy6agNjYdv2KfjHlvbNeT/Kf6NCijORLLlEKYXB6
WkBFQ7Xb5Wag07nP+xI9cZ3IyppvGf9epZ3RyH8WtcPJz6YIPcxRtEb2qpVXhAppqEtXSQsCVnO2
O9qSZpTAR7/8rco8hfk1r/i+AwJtAWcxat6AJs9+imj6NE/UN1PBf0kaLwNFkvN743bpaXxm2Rw5
shlGN9L9tOuYqF8SvY4sYSeZM4SnHMx72oqexwyn/46+xoBdIEJlvFDMUgq8/jkdRu6W05QqGUhG
0ziM2DriYqRsX+NQoK8Vu6fUEpPDL9GXTRbc4JkZcAv1kVZdLToTF92CxkDkN2ih9EQ2aG0A2UVb
LG3PtVibLF43n0U+0XNlPjD3H7mWPTalRQgdCD7Q9d+rsyxVh8tMqYK/ewH1/b9WPKSvWRL1xIM2
1KMe8wgJUx5ZqMwZzONmrqWrqCdaC+xPZYQ4oDDw9GB4d3J5JtH1yx8N1MPbacESvZE2f85JwkPM
wNA7TEYonp3B1hJPSZQu0icWgHXS+OnVhwDRm8HoqWZjHbtojp6Wn73bOS7HEY1jCpTxx7rppyFX
PRecukVgb/W4S+EdWzDyGk5RJTuv+2RBpDwh6A7VdoomHyI8YMYaQTIckKA+6d9YMJf2hKPZP3fG
Ogj16mY79Y+yeg8HgoLbVGdXfsIYgwnUL4FzcH04BtJxwtzBVTyVcPpUGIFT/obmksQwkVdbyrE9
tumbP9WMTfF/xbBvr1A1WJ/Mu82g/UUC5V4+VUSyGrBU3gWM+Z6q6hHmNwJ0ZMagjUUv4XGDwdVT
3BbBbe5y/K0sItv6org3rsGoy9rmNA6Hn4z1A1NrNbHhQ9dF6v3fxcJd62WFLVp+jJWejAWoD9vM
DBW+vZpv+7cyLkNiF/B6RxVWUUgy9qyLiKazBlKUaF5gjlaS0hYJ2Gdj2wL7Uaw7ZqIpO5PUOqIr
zKd7ziV2UJWYcQUq+iN2GppNS6y7Zaekdlje3quG6emRAPnBS8AXE2Aei+Le3CGhFJyP+E7/BZzc
gadeuWWwhmBNjhDXrQzV4uMo70IiV3YnLuTL791treRpC7ouvJ4ae/R+zlWJlJrftzKrBR/K/LQs
6U4+IvfVJWlo/tGkLNvI7CxXs7+aFa1fE53TNKkmc6HPhpYlmgwrFahEckLQfexhOVqTubzw5k4y
FPRcglx2Jct2YAY8PcLIhywu8zLDMEZBOtIwlqqJ7PHxirGvOqd/gZVLFnOgdcTRiSnlXRyEfigu
kKnPue64+3YVxWUKswvwzad4miBD+bYf9AlsgjinZTDJSEnMkuOtLPdfnqtv9dMOHbz0guqYbcMF
i9lCp3cXxsbgLI14NLZZSQ+bGa9KfXLiaSkryoFsW7Ik6Z9II57U8KzXiwX1StxEpFN0eeWCqwE1
FD9VzaLQNX5W+4KU3Z8lMF2tpVWysiqB6Gb/Em28XkRBeAamGNrDC7lacIS70fXvlGGi8c99zNky
J8vbbb+eVRoYBSf2I2mUZZJUWzP8J9vboWUMO4CbiP6m2vmVqaHw9Ka8O0/0zUbMDhU+6EGIQzhg
V+bm67tcSzQ3v1QxZ87TwM1OLSX5ZuPKb0is0cOmpizRvd0KDgg6s3466MG681GifolFUBf34A9K
fORh1JabYE2+xlAAZPn85n4AmdvpFL4nh8p60pP6ya8dUQ3a8gctrbInWzWqHWhYHzOOOk5AWeGC
2+TEwiAJm7qMaV9t5JuTiRXU39NtHzbIkd/6yaCFkyvdjC1t+4pOKu4jML9GEpzpJ7+iFmL5plBg
AozfSU5zZy5XMGyKX1pbAv5ohKZePMLTFuqUAqO/HCSEvM/jKF21sdWBxsZoDlfeVBubrA2SpBoR
DgNu16JDpSvKXknV9zOfDAuLH9A8iDAhW+DAcD8G7L1dvpSoUb3j5RYZagca8zYuKctwmyTw0amK
KgPjUtB7RN6mNajnXzb1BLhIcOsfXW3XmXzZ/QuP9Fdbrwi7WTAbNJU0gmd8phzeeVmMDicDsFb/
bsT09g8i2X4SJ1XRYhrslxMPfVT++q03Og2wcgHLNS9/Ed3624aLW5ZpHfkZjUpGdbQJAiG1w4kq
yQbS4I75+CbfIsyNo2WnIjADJ0Rtfhm6RF2UMX7aPYXhaV6hJ4Pvz+sRjsq5mS6bGMKXCHA5kJRV
bGE0KFiLk6bjnwgE95BJ77uqWQiZAJmJSjQMTWCSm766NqkqmQMZ29EtX4Sx5N49rJSVgKs4pGAy
7/SEvGDTLltPng0rsIYtOUGDZl/9A6vxL8hi8SlFIdv9ddWuPqc+M4bfDSAWFIJMJfxdPq3888P9
N1NuDWUY9dKle7iNwXaZj9N4H9F5gVXbcMPcHZlyJg+tk8BbXTH+9gL3hrXqVt3g+3sZjOgaRsw1
QCZULduyjdY0RHnR/cZ8tehON+UtkIOGC7MEZ7oGtm1MNc9GMoWYNNvMq9SpdrByAigMvChvh/xy
7D+6JblAUAhfYuKtA8+o0UdPAw/75Z8U2kjgkngAnYt0X5rRvz/hTLRXd1OzJLItZRp8IG0qlSB+
ZYYjrmAzVJMtn5wtahmc0ZsN/rz4RQaMBpekNeNUhVlwGdja5E5ahQL8xGA2EFOUeViMYsbfkWDe
TkYk7SiemNfGCiTIcw6NguQfVDBtRzcy9n4+bQOJNA/KEXkqA1XxHxiHLUSX7nZNpGSZg6zAqUfj
sdZXxHAa8roeyglm3fn2DrMisSdhAaEAko4ZFLJLx4HcKi2C0H6afpqagNgoT8R82hPxFcfPq71c
vKtpujC19dKeWNvhCMi+ofD2OvmVUYISgMoVBug4rbyxfIVhkW2BMdNX49n7YBkGIxNpM1ivQ0DW
YftPDhsb5uPdXscgU7h/olhaEDtczDLnflqDGYd65A38KoQZq8ZkruITnHOMQBf0n373ENxvfXDy
xFfvWKsoLGiOHTUUiZW40kYSO6bH+WU0tNdunPzxcKzsoywJW8kSZasBSCwwvccaw+hgzH908SMC
qv/0B1tBO5Bqm2wqm3RxIjQOaeVDwydsbg5ZSUwxEoQbHbns3jRpOmS6b7Q2wQKqMFevkrNRruXg
rYbzqt7t0dUA4itNuRFARyrhhpmNsHu8CqkXTMjxVkgAy84vMW8/QlwfU6AyJ8PXJ/hZ4Jbq2MBk
Ke1UezqB4mQlmMBJMF3s3vAheGdhRyC/GGrwrC4C5OD7yUtIovZMNu0N4xdtWdivrqFIZGyJD0mg
OJUl8b2I3FHZpFAe/4mTFgfMEV6o6EZ1cRfy/mS/d9RhNCx2lbufvV9ZffuXt0vTQL5TquhAAs31
zkfsLV5sj8zTbyj6x8nR5zdpcw8Q9kSPsparMKd0OzXII9Y8pnLubkwvpCl9MWgX9GzCGlz1LN7T
qx4GKvYR81r1On87wxk/UqaFXO2ECljRU927wIBSefDvKrh/uIT5GsJFY+TPwta9+1m6V11BsWzp
x0BdQdejs2wtz3MfRjkwQEksjYxcp9d2fAUU+qHnLCut/RaWXvmm+y1VM5l4goXAXFOD10QrO8oQ
1RNULaXVqohAzAUGLPmtIK5QKaOHulHNbh2o2zkMYPbwDqO90SrpT+yrp1qbt8mgLsNHkQvj/YTy
wKMmTrnf2Io7U4C3rH81k7APhPAuI4zUWuajQXulrxXR6mIviS39VP4cdiK2/Z7bBYP1oKND3w59
BCvlbINGLvnxwOwFUVrlSOiCLb0aekZy0XWEAQcZ9Zky6d3XqzDtGnNvOVJgq4SzXfwvdp4C5o85
kXwY1gCesM0hN7iImMC7RX3uYgFl/9HrY9wp8AZtyKyuCGfzZXTJkr1F65vy1H21ZYc0AI8ekoZd
VpW01nruFmTLRiLVUNIHb6yoUUOv/tXF44jS1oC4jXbqml5+ztCYjL2Q/LgqP0CLa72gZ7tV/ln5
jS1GaRPPPs3EAuT5HFxxcjCBMrPfNhY1zOTlW3eE/ll+QBoJzBrrreAXZ1JJbf1waUBNdu6V2/yK
eoRvyq3EGglrK3efQjiUn9FTQfXWk7qUpSEz4ezXl7/x6IvRiXGKhcsZU9EWxQ3+P+whtC3K/h5K
n/Z6QaivvvGt7KVPkehIYf7aTZ8DJHp4o++rUq9tcDwvBdpd9AbqZ39+D1KhvbAyV7Mnouba3L9Q
XuhQGodcPmGLvY1QK3/qzTlBlcyMkJaSWZ58GGeapv4ZuLgmlk5yM9D9DHpF/6hvRXpVozC+8KYb
oS0/rc2aPpphNZPJAKl3EOq8b/H9c6GJX8EO/1wKesouzQminXhdJzNVDJdfulXqt8XCreLZQx7x
rjD4qXqf/oLWctSomJCWkFgXpXnNiGfFccKYYV98ddnJTlv9dWrVlMB+ZiO6qzckpkUgP9SPuHjr
2qx0uOtd5jXQJFcUSBwGnnyZV+tf0X07g+hH6PEOL4tzomNTNtw878pbn4Tv9WDrmfgLytIFMvv2
GoebRMGbTng58FrgDcz1JE4n+mkN0165qPASf8/CxGaDFOKKX3vM+nUGUNucGGDcZ3yaxjOyGH9A
QkeHzFWQYcAam5qXHXNkY396gmzTBcPTwDFJSELGZWS5Hna9mlkGoS/YSKfR4XSNMLA2YhKyyUJe
GmXZ4v1rELr8dHJA8Hb9uIBgzP5ZlWmgIFvjOJb5nHXBKmRooWmUoVkDcZtuVC58gngq3WO5dE4N
Dp6uxs4rrxk4qU9VmFophQkJatVMDPFYxb8lzPruKd9rX2BxxjcrhVdKJk4a8PJZgdRfvsq5vGFv
sLm5d/cdn95QHUktd2qi3utLWkZPVGV07wwKUddX6zYRY+7z2Xrxz8sHt+90UtiygtDBZ3MV29JB
1Kiq2/Il+J/DZRQzIVpzBPONehNv3pURQyo9UbT8fwC90uG13Z8CPmPw8m/BkyZ1qFqsovB6hZbk
HhjC7oHatI9XLoPm1Z5VfszM8a2AEQJml2p92zQuD21detiI6S+xmGNBzkMxMfjMtCbSqLLaYeNd
2bqmmdAJnUmNxAlBDl+QFsKsRze57tgWjUT1URUbq00K5MYz+qoWnRfg9Y2XCXJzr5LIbaAXYW8r
A69jN/q2BIKm/QJOtYlUgfiKdzGaEv3BGVPMyeY6OyZtyvzPjpXDp1KYUXDfsamHEMOR1RnHzZ+x
R+f6vsATylvO9RddP9bdEi365yS0bl/+y8HDqm+C3ldvNFxFHfGJUel/JX+1Z9nXoU+q6mFsdPHf
5uu2m9mxSR8SBz6+d0sBDEC4Qj3gfED1uQbNwNGPYwvq9y19ILGwBUswLLfWR9Hi1RAYcZa+iHzx
W276nL3JHHI30tKN1qOTic5fbMmdAJDeiygjBw9ZEwg7BMjLcCkZW1LBO8tLvk6CeekbhZIBD1ig
+IvjfVmbiJqhXSVEQfQRzGz0pnAw9tq1oHof/DWnYg3sV33PE1oCPLt7DQvo/T+SzKizrebPt3Tq
EUkd7Z9CrU+39pQUZXNG4Q8iO548+3B4spJTK0iT1zrLofWnJrqqkFWmpOpQDFMrKP53uKjdlH1Q
hFg7IjMb5Hh5trFeCkS/EsH/n0FVV/rcV4JG8BBiKWzGEIC+SdwvSPLly/UszPkv7Z5C92GF2Oh1
l6H0WmVVTgPqrkl9vdeiYWdwXAI3/AVWwj2IrYmUqZYK+Rs2Oj3ncrjGdffjJ6EVfXyI288ZG5Hm
wB7WwvbIMs2IYtXz4jD3zTKx5aMa3MeNsG2mRLeEZUk+LzchuvZpmfO6lnch9be/pzfUN3MPHk7x
aRRLKn4OLke7cxD74eLYTOZGpe5FKVsqlMXvTnCckTM/oKVD19kv3y5JAZm16kpRYKOzh6Hh7YWI
C/1JdnACMk06DY8DRjxmzYN7SzScxk1LK3MbcaiSzvmAeOb7fGuDGC0nPONs9uFALKqyOy/KHMAA
U4xOobL4gGr6C6ZPa46SVya/rjpE+RQqkzXbsV1IYFqV3GRFmYx3+J9vlFckN2D5PO9TL7ECeSH5
VvQFwifE5r5M43Vf+bhH6hIJd70RoOi0IR9KEGBdNqLqcrQZqPcCdsAah6lQ0jpDLuuYm2O+p2xj
ciXpdTfZN6tIS/DWajfq/wIXlXhAYz9bg8OHOYInK12SEQZzxs4GlUo6NM0aRPS/0BKeMyO0jeL+
pd5JFZ9bhaSUuzfWdUSfFJCUC3oHQvhvRednF2tlboIATgK1wmIiqR9NNUzhkLUYu4bMKmZIfYIu
WxcUBvM4rcVhP9VnEwJSBBZ1YhHOjNfeqySy0UD/RuUDfTn4NQCe+9JgBgQlSLjSLHybHSjJcjZq
z3YgAkQbPEvX4hbK2IbvVFjEt4kSq7FUaneQ+P7mR0kHIlMQRs5DWDb5F0tMoCdsXrTY+PrDNBof
KNlAgCKY65t1zFteEIqrUobXlnRORzPCYjGTlHgz0fwzzrUHso6PPdiGfDubFskfqvylWuyPpJ4b
A30Gikspr6pXht9rf9wYtm6gF60zxkEUSPcChq6QylKbzL4vO0eDwwWXrCuGcTLg3nm1YQKhjrYB
Ol4dC+Fkk12nIPPJB9mhV2s4JtsMEnAWf1OYQAJYAwUAUFmBv2WbUKMY3Cvlo3OyDkD9Ltmo1xqU
RKp548YOfKA1PHNlZUSKxBZlLCg4UWPzaxjcwtSairqLcZ4SiMW0D8V+x3fUzefpcVNTw5swVN3A
BDLwdQEvpjhu8yZPo6BoG9AAmUE/I+f6u1iVYeB4gLWAh9v+t740vCjAyeYtb8reJkU/TRV3oUsL
FAl25/kYHoFK2++YYk+g5BRljVdSA9ioS1axM4G0zr/uMclf+SXpQfozFUUu41irv+be4DRT9/aT
fIpJYn/cNVovDOmkIOpBAYWvvrjo9VuExmSLzuri4WJWR9bsQCzeqAaf9FOPojN0b8ClzbZzQx+l
H0BeD/oLOtItqnfO9z9mFANKY9gLr+UhnpjKBw+dj4xx8ut3yz6tDl8lOV5ybO7wcyI6SLhGweBq
cPRVH23fql2eXkBy+WYtaHf+OgCFLMQqSHSAT0O/P/z7arhrzdxHSUJjkcV2mi4m1GiGleu9N3yW
je/XyUTkAdB+UR0IMJjtBzlDm3652e5n+ZnoL7xGWPFAmH85gskao2EpVT+mspHLcatnqFT/yV30
/Qc8qS2Mh09d/juDCCsIeqC27SiuJtj+YFr0cRlgfua6r1RSNtGvJlGl8QJEIxCIZUJRKenZzgXH
ykqCLHq0qvOr4XW/pE8KrWqlx7y6+9ALdy+jBztsJWZeJTKfVzTosJJYL7nBATPP2/MI51lk4qFn
79podDbZq0EZdJTC9l6tuDp8NGT59KuoLJNrpy0dgDFlasWgOpux6MTUkwWt7effSTRkjdsNntDB
d3ISTMkVA4kOYM/ddTvfYByXD1C9GKluW8QDh9WGNnM/FQ+BN/xmEL27YsVNBCqiU9WzSugd+Gaj
0KvDugX2lWChI/KP+mp7yvXVllz9hfYqHSQsNfJYQ1Ar17Guef26c4egf5eS3L5PzCKnriFVbjFP
Mbg2Jp/ROtMxknobFaaAi407ceAbQ6XIi8l8gIZdDDmxbRDvqaPIEQuitwNmgz7MH+pTLRasoK/3
BNlDnMNR8vf36pT1vscJFVCUqlEPjV6xzDx33M1RCVvCuEQR84CPbxAvjLCOEW+oimHWmA1s/o1u
fYHYEZWKo+Z/C6knzcyPKLZRVUD+uBoF6dBAnIYjDLDqLwr9DfvLKWLRWpE4veTOGvihah78Wenw
McewqIB55XQ2XI2MEAoeLJMg8JsyJhaqMf2k5yn+GgWY2YLC9N/PoD7VgMqTq3Y/480YnFDeyXdU
PVJichTUo7bkhMhTBilVrfe1jiWW8oA+f8kmE647PrT76dB8r9+G8DiuZ6yw7YKZRTjzV4kYMNf5
Gk3W7viBqasM+hiaT3br1p4O3EMCnd1tMFTFUblX44zK9zBYl5InmUOOcwh5O1y4fuxVB22X+Ioq
anysg+pf9sJHNuXJmb0hNhcoBdCf+PiJqSk0WhEiO3ioq0M5iYVNaTF0vS00+2E+Rt2vACJE/6hH
s32i4a5i9aqNTcH9M68xrE6cPJzDJRZWl4Y1Tcm7ohF10Db9D+UX3UcO4X+RJ6DZjx6TrJvcP7Ev
czGY9nkA9JH64PqrtGoCG3MM3aDw6CzC6LUYkMwMOEuDoZTVRkvPR4NbqhsgG30RplXBv2vePdxt
IINFPrmoZaoS95yhw9kJ4jdqhqv5FLhgU8ma9OmxHiv6YxgngxV9a6WFWpPK0V6syRQNzNzvFKdP
ZvtsXCPsUg9xWVgVwP+s/FOMZNsrf3z2P30ALhH5v9/PrkGuWVjU1FfotFeqGq3HfLUEtH1RiLgz
lCI3jc3PaWiA3WTNQMp5yOU3ZyS45/xOTGRvshkXKWQF6nlnG2OktVvr2eSK+ADciog/5vspqP/X
7h7Sjdivjk2WNYzj+llI9/xHMYyFCRBLER2K+lMcPVFHsgV/6xSV3gz8zN62GF6IHMQgOmC/kOcD
PSGYzdHckOKIztUTNxe6Rfd8/E9Xnap+URJk4Of61b5oJVPDetFf0hn5SLPGtJicDBxpIXMusW91
EDTJZRRUw12sK00UnBtTohi9E56nVYJcW7cOYz80KnoQwGB/IyJRZqjPNMvaZUNHvpfPVlAMT1Cu
gLsZgkoA1Jk84i5JoqSAx/mbwaJrdxg9Is+xvxwk3mwuubz6wn/AEkehzNlnR2+/0yPiu/IxdIMe
ePAi9B6/dknk0TjN1xzFclCeOgLhRQTC8sipH83Ln/I/ivxklv6ni00tqfURITbssOCaS2BFZIHu
BY0DfL0tkbDu1FbOVcxmLqnzgkx0hyHGUomCQIX+AUXYY3bDRRUQ1RCXr5ra3fmBzxhtVwKIXSDI
VBfjhIULkSsZZb8LfidTr4ahzDefgqKutngfy55jKekDoidTJp8J/5pWBv0EMwM3nRgaymVgP24v
jpthSfIgWIQosUkM5yOIYGxFwsz8g/hmZkafsv8cmM96VSsr/z2sF6QTjBUIpEdUzX+AdkQ5oOaY
3eXPRhCxWrzsrCWt+nuWa4vrKQRmFOU1WsDCUXF8G3z7lCs1/ILlZfjwzPDse+EXIQpIJ5qNssZi
LHx+eyprs1vWS2/ta5EAuSX38YlXpnXOArec32+0eQJey0m1Z/zQxENvKStV7xR2nQXLJEWV38ma
hQLTCuPBraR3nZfoBc3wOP0kdPaI7IMzoplsWVqH11mOCzFcp+TvkFv5FoAAOADzlpX/gWbQpIHZ
ITaUchCDb1v8odJ/M9/4x8Cwd/hArWQnmf9qIRLpS7GOuC92rXVZJ0VWANaQImxxSvwFuzDUkOBA
A4aeu4H5SeNp8TJbfv/0M3HOXhKpXnedHNoXAJ2dCj4JydfRBsGRrwFzc2vz54IUygPK7P9n0Tzp
miPbGP2x1jSbdwixQiTu/QrdVT4CGUrkya5in+TKhy+Idct7HMCVSXYtXtlO41qMPaK3MRCP4Jve
zIBBy1SmYoN91Vv8Y9RlZhAq9TaxAp1IPoS35/JT3+k1b8ijznq6Iu+axI5/95cM17gqNdIl65aD
NREvh11RIX7XMy1eEIH3xNLdpZ5tlbSybXC1ZcSLX5gVizodnrOboIccQ+t4oUz7xHfu7lwhksdW
o68C69fgeX0mwPMr/KdzYCimAUKM35F0g+IZJt0Ek/pQO5nsNamLmsmO7m8skVExer4nmcgD7xm3
MyX2T7G17qMwyoL/PfhVk3pWZedv6AkR5F/Ur070esxudr+RPF3gs77w/0x3ZLkfjDutTZMsauqR
t5naPrzYSoeZ3U9NDIk/OQFgoe0ZpqZ4PBssIaqkXV6ZgqYtQXwOnTVF6SUUOL6QVn+fu3b3Qnbl
TL9ItQ7yVRttpYst/yvV0qSx8BLyXR/oqN+ocao6JBDTjwggcYT1Q8t+waCyzxpe9bG+pKcmuEX+
XPGK0oi0l8Q7S0sZ57EZc8X5A+eVJOAr1Q9JJ7vA17gFvOU0nzRkxCkgN7Y0gTQ6Xl6Es+oSc3hb
jEho8ez5/YGbvhcMTQ8s/Dt47f9neeLyjE1XlPbONiHwJ5eJfhPjfBwZXFF/Rwb2RUNzGXLq1iOT
69WNQNrbKcU+oaBDYq9LYPOVhYhqYsk4cQzsvQDICfL9Am/mxizqhQ4XLzZ+ViGYb8zyz3YO1eRm
4tKcpLW6MTjQNpy4k3h5iCi8HSuRUjaZbrrTzCprCu+6Rhj69+l43piIhUeZwf1/4bhRmbXZxKwJ
AG3Kcvhnn6tUWf4bRrC+JPlVQejwl3DLLqJW78WCzqPU2kLKzKNoPpsQxxPHREg4jdPsnlIl93s7
gzxmwpU6N6pwrjX3aSrfFgdXwbuvlOw9wax8lEjsXqRsLSbfRLxespw6H2vN4c2eRYghEPI0+2aG
K4v2u1saZkPRxJzeBNf2YEJTNGM5OSdW8fZLP04HHSYwjKH8GxfSxQxIQaotAFBlyqzuK1ZIVfMs
XkKqxDoGFLg8Kj3G9LOv6btBh7xUXZ9PfOgg4TnPKv6Jojl2Q7B78u5vulJYvpwS5fmNhKijwJ0C
wiVNbSnCns1aGpOQTl2Fx5Swp4pAHe8Y/Y5JuQa53fn1ESx9J4qZKc1Acvc+2l9yHkmY+I4wamsU
u2fxGvI1msfvKWeFEPNEYinAOQm2a/VLxvvsKv9iqSec8094/FcGLZYwsNjks7nzcBCpJX2ePHJ3
xIM1h13BXIjaJIHQTeu+dM8lHs91168ITXowBP58fEu+3FK5et7O6b71hMW5HsnSPVQBo9InI3Dg
rov31o/Lnnwfr4NLxlWkDu69jD8q87kFVfOHRowMEwI5/0aIB4ZE2MkMWr0Vs7mcWoJOLKrRaJjb
YlbVBlQEH1ax2/eV3XVOjUN8k7fkJlPELluyWkKqDQ/5qQDi/3e0NeEOiPdPfNYkj5yNRRQ4gqbz
QxeHMcLoRDUJuznCLUGWTEdESyxoiZAXeFzzP4fj7BwtgiUa1G41X9G45v+TMCpb9GFA6qJQPsSV
kosQ5cdypntLtC4dPvfVbBkqiMsaTpJszqJI0Gey9gSfRof1zoBJHGI5n2IIxL6GOHYwa1VSP6Uw
6ARZrO8uEEJHTiHTH0QSO6jjvjx257yGGQ27WtQrCOehKbHEdoMwqApDgfPP9MVTS7cL4IeXXLzE
8VlC4zYz+xQzBt+/SdQhqIdv8kg2/8am3WTdyHMY0QajS7qN+1lRvDREaPAxQ0fZXrMwJqyTP/Ri
RVRk5TTLKzkrxs/rlyu2qDF/DRM/mwFTRqTrC5WtarA/UaMXGw5vxNU42ptwW3h1zkpNpKdRJHeN
ncWXtQ9rUoaTh5eYBxo8bbLxo/Xsz3UBCQmMvFmVrgeVKMEfKk2Pwf5E7SWr81m4DHknImz01xlc
ju03ZP5Jq/hKpj3jo+dhbYGS46h1Lvv6sHeFKU1FilUON47INuo5ftp8wPmejzlMKiqiowaAqKWz
8kB6KcS57ru6wFZKwGG9oErtXKV6UofFTikv9P7+nAHynKIorqxhaxQGJGpA3OCFdXhl5lxgyEon
3OYZcVrUdKgu2N4H7z2JHDtfR+lZM8Q6Zdh4vjEF1dlRDW3M4UdUZXX7WzrvfGIS9ulcpM/DRvAu
TcNL4sTW7Rcj2rUlzcFBlorahbCYCUD6oR3JfOkGG074BF1pcBOqk/h69Lp4p6sHaO/kF6AUmLni
rj05+fxXgY3war4wrs8o1ocpaWiGjtBvAwm2vO4Pyg2loMjODYDlD2yVgfHLvQ7r8ZWcW4fbKGGJ
QO/BrSxtzxlFuobB+aiHJ9kVQquiDHEJwxzWemFpgUNqGzR72xjCm0iYmJXm+iUmcnONzFdy74rz
vOkWFZ4YZw9uw/7EcA1SvLW38QT3IQ2ItH1ZMqbVINJHAqSvVmJ1uPKo4B0jsZBD32KfTyZFrQ3F
kkqqxtmiyo0S1kM9wFwGlafkUiFk3DoVA8359CKZl0Vyxxp2tFMfT5uEGn27XN3gND5I10UAomSg
3mwcG5sjWQuciS4x6fhBKC2OFr4TyEENDhrC7cJqkOIf30aqKMaOqfddJl7soebk6k8Ex+ZDmz1a
iOVETETrg3MOR3LZLqULvzM7QMqy4VChLUB12x8h/PbXmcmFqG0227bjTnDGo/ZcDra6tG0f/D7U
VjOJDIpn8MBgRC07PB/BwOuPc14T7oZVAiaDrf1r+ZaIynVJVYAoHgKjTqnPy0QHmdyYo5gPHRT0
+caUhOUVbViaEAhK0B99f+4pVSeLjdl8IMD6560ATodP8YCRSnLZtNl9xD2C/s62YaPoieRjSeuA
SN9phMzUDFk/TKeuAYrUGlFFgZzWkZxL5eGyFtV2iJwBkNHUypZu3g20QUiiwBdBgGNht9L7unEF
OMg6M4fDFxC2iJnINsn4kbnGwxjlB8xlnU13FoR2ACoehCaMcUgg38Rt1cltponNux9h1eWa+Iur
5qSKnkfT20u7ZredqhYgOSkNQZc/xOBHThFMh3nimdtMsqJ0MOhp+W4hnu4/JUIjX9MZ8clSHxDU
SppAL2yNvVJvKVLUXpy7IkODPYryKckzfG3b7zYoubH7MzFOBld28aNiEf5a8GfOcasPfS2cL64p
BvHXmt60LNYZl7KdMwg+mgogAlrT3IG7yNdWZ/RpCBM0rHrsJh0LhYlD+vM3OiXXGTH5p5oVIu45
fbEdjNJ+BpWTX92c2wpqrPO5M/NNSeELH+qBOIq9FkiAXHOWTYT9HpqcX8nFIiWBe8SrkEfLBgff
kLlphswfltBSiDnwBfLenEueF2EAGUimhrXLpnO5DFtmettQ2nAUMGrGCXMDiUOJM6wHA27gj69p
o4XiL4ze3/Vul988dXY1XGoDfavM/fugSx7rLg9DVkeYLCkx0By7mwULXr4U7BB08UohG6ur6ka3
X2It3O+L4UHI8ouo8xP2GO8ydA59uDQ728g7FhCCKTky4upO9VbIz7U4itZMTQSLk9VNVdxxuQrQ
9c+gu2jzHLHiSe/EXVsYfhCzwmY8IU2vykmqjWieZGqkv7mOphL/u2wQH/gRf8uBgADtBv5hk0C0
LPeIW8qbrBGrTCo4N+VK+ojEXRi8AJvIWmHxVyKrO3Xar5JP1D87FIndzwlcoD5Izk3vK9oQoOn7
lvMSvoFdaOpOywv174Gub35heAwuVyUGHmYtqqDE4jVz3JmxYnV+ku7Iyu3eXcIF5Vsq3xPQSjF1
vB+TYcwfxMih/47vmV/c+SnM73tSwcpz/i29ucxP0tf/i0zpbB6INoxhneYOPgAyjuLs0fGwtVk6
/wW1m8WqZhJU3hXHZyv01l3JVWbAXr0I/WFsejhLHZYU5sTzmyjWi/OBJJqkkS4zxvi/zLIqY7oJ
JLFCYtHPtN/TfUNEX97C91/OO1e5cEu+fiW4mcabkKKsx+oySZZazKiwXi6zT0NZBGa+a6jkIJb2
dNoSUiDS/0kuX73OwsAeIU0CxbUSE0PTVrVQ8mzRN+5Y19zajNiFtDWogVabMy2PqnY7s7w40i0w
bzQQqOQ/YOaJggZ3Rrwzm6umPzbx9EkUKU7oz/oeIYmDHfvIUK21SjTePkLvvg6dtPatehI5RlZk
0UqHNntJdVX8faNBM7Itlnv7joLmnPOK5m4SAr69wGzO4sEQewjW6l7hoZ/Fpn1sp6L/jgulXLvK
DcicMRyVJ78RYLboViIxezhHWvBzkgjGPj7jIKquz6uq4IKJ/Jv/6Ut9k6/4eUMXMEz12Du/wEKg
t353TgWKS37bZfnJBzNYKeNu162fRc5iH2jvUOc+Y/J1KACCV1rhCkSdVlluNQsWb1BcEc4VTYyA
RsMGE8oFY+oZGAylEqNXCOtZ/Y8TZxN2wmuHArshW/LcDlXZAh8yZHkI3mHehgZ3wBBxizH4mNak
AhjJ+Qtr3B5+ySG1Wb2NQAMvxs4aLB59o6wNc9j0QiCCv/aLZwt0DexDfIFSrD6eW9d1i/invQhH
NXUWRUk7Mph6jnCThcODdZQwbleEBdYcnjp303bG7w0sZ0mwhLEVcw93h4Uw0LD0FOxB1LQJuRmR
lWYiYxyWv52p95pa0Xh1WdhnajI0+/00fjWXFeAL/UatTvsCqN6vKMgBKwt50Fdbac0ZPIUCTyfd
Fk3egVU5PrRZ71PLeI05fTUc3NteoOgA4YW2lkeAeL1mqNPJL2/7Tf5bnYvhG1brhdKYgl8Ss0HR
Y9CWMXRBsESnzoutH4MhMrAoNXQowPUyy/9mQGkZoEJR8jMMXhYLvt87k3/HPhwPXazI3zjC7/HG
nPwfoq2QJsgwcojeFWh1pWDwssJ2PQayuk/Kdy1MmteBp8vF+/dcwXPv7i/GaoRXC1gIV6/LSOfq
xjcwWxmsBegTh4zu2TboGQsqyljJlYxKJ2tt12w/+0ArfkhqHyXIQhwGfAfI92Q690aH77cNh4WI
GvkpiH0pOm5h0aLus7OuGMlzZMqg70fzjXJC/IwLc365PQtUlPnT6SMAvBEowkwpXeQZN66O5DBS
g0OYx8FCoBhK5+9ahKXsvGob+9q0YyxDmkFc8QRu8+LJuK9gVuBGchiUAvFqY1GN/zas0HO4azdb
ispioB6j2MEefIpmvNXLJRDgCjHy1xQAlJKV2/7xNx0fYIsL7RAa0SElxQjX0xAcRhEZj92b0Nxv
f5nJo9Vqa6YHnusjerQyc5Cn+es5OgPlIT6lvHn2uIf8PZDOUhG2qwDN1JiJOf1ZRPq257A8XY8X
MB2h6nA4WjBogxQUXxpMhk5CheTMVgogB2ojE3sIYlXfOGWp6zcs/9MK2sB3X6O7vYYVcjDVipkT
bu22DEn0INss5nbxpMQHm0CPHkzXL2vTEC6NYvn4UBdvxPPEMlWEOIwVGn0C4QIUsqGp3UFGkMMZ
0vWCJhV3g4KMiO3vy2aFRsTM6f++2UwkuNxBTPk4pMWzRUZ09+1SJykuFmR7+TJhdqrvN8zlsG1u
KN0cq3sMr1fBwUrRpNyWNGThIWJp06wUGAaLGHE5QuuXjA+qs7MUi9L6DAZ5W+U4AGUjTMFs/iPZ
cfoqveRFJ2FMgIQX2b2oJNUCKp4MneGo+8GlU1CIMPa5VJTbKPaHkuPfSlQtTNLEAJlw5wQRhL26
vcOV6s0QUVSmBkm1Iemf1aVFJBblAPUK3z9/KVgr1DKwH5658bgClppNClXvJZuOlNgq8AEioJzD
iSSdDPi0HwTzfbkkIgUU42CCdNb1HDfkJ+mS4FikWsn/j8y4yQ5yurUG7W4ADInQoHzq0NaDWRFd
e5YzGl96O1/WHSB1f7ASmNWflTfrKqRZmEDw2VhKngee1uo6fMIjszT34/uUxFUXxkFORzvF4pAD
jCiy2hWsGvqLHMw0AEW12UCQ1x11Hyiz2IXES5vS5UStUiPcjMCm2LUNiff8dRmzZw4RF4wjcSxw
iizBj8bf4b1JY0OyaOQ66rkEZyUHGeMfQ4VMncG3D0TmB+rTDEuUBf1lkbZ86H1q6IlciGTpNwA0
0zpB4OIOreMzdJvhuosOUBobx0ntHRcQFwBYQJIeafnNf0E1kC0lSqkbRGuYpd3TQ5gddTLmqvuF
XGJX9LU/NDTQcpfApItkPdECyPUUrmUDkMJTHylLQ/nFyuR9n8trqmy4ScjIwIwRTKVZVYJ9NfTt
vGANIhinZ9lNvLTv8ylu/TNpgD8GWU+Tuu0jX/+m6J7+eHXE6hE43Z6TxLDVmOyNpGFfQNr/u2cR
OnrQ/cz6eB/EBefe2thLPCVSCN9702pRdkBvZWSdFPN69auRfPU5tmIEWKxIabFEfoZIg5lXoJbO
gDQ1is6cF5f4ePScP2JtnaqQeXVGP5V0k641AsjVpm16A4bxdqEEHDpBQXUC/KpI7LOAY9mbVgJC
/Q8iiBynRR1nLFCvSMfkF4jELi9IHMnePwClsxjVh5AvyUCuz9Q0aYykvXLtDgQfPz7zFXheem2p
xe71nO/LIwmcf3b1KozJJUNdBDHQ2p9GBTk4gh94BYWh4uDwQ7R5pDQ67R7KS6mAd6DfE9P7oGCm
JEMBCMAx7uv7Pz7tmlFl0MhBtKtj8hrNHSpo/QkBjF4VzXhHBejlXIsOjGWow6tkvyV1jB6v//4/
dNwL1CEtvzyt8qLbCHig/U5MEegf2HZK5fzRzbFQSYfxSDa4xFITGgdL5N0PKd+Qr6vsgBsboHcf
AVP0JrYrCVMmj+MCBQxhq4K8uZh3zs1fqFwoPJVGl71vUVZ6qaIPtYLpPgAKHzQ45MB3FTAIXCqa
yF8tCd6WsfNwKIF7Yw5sxC7qPVbJqWOvinQVyxri3ppldbCw8p9y2cI85SZLViaeBmdbYSUjJAU5
xTmGR6KeIsPEaRozIA231R7BCn7BWeF5kHuIr2W3EipBHucciY2PSwl1SHeg44yLHZ1WakS7QLES
sXV/m+QjWwMiF6MUyGgj7MtDMbdbXlUZ6Hc57jVJOO02cAM46S/dNmNXzU6oir3nKJ7+1fCb2HXj
PcitlyC+k7XmTpHYAgwcAH2oRhMsVtzcmXVkUKA1qHJHUeGKyLofCytSvlD/SrYm6+lhFpQIUhd4
lydgzsfXzzPMIe9nXsGEB4vShG7cRAOTjgNR0ybdyspAumMcC9bGgxhysMumPq++PjTIzc7evXSH
9w+8SyywzL/MsX4KP1/YmF7t/lhv+NGiblDlgv9XuMKBmx4JagJWr0W6kH655iux0xbdCucYuo6m
fxYleLJjk6oblRt80k7Bbjfe4q+CfZ7Wj3xjDwkDOqkq38Z34JRG7pi9YVz51lcPNc2BHYpu3xEl
NTZGngW7gxpcgrw88OkutUDKyoxPzw1hufpWUvfuXzhStq6RRI+/RCH8Wv/JceBLhoj4klQgCjoT
eKkynkA0qPG5mhW4S8WRsh8FuSmK//uveilhaPwIFu2oXeP4ezCFj3T3oF87GwXu6Ze7LcylvWl1
3lNx2uEgy9Solrh2vW3ayH1fsPDZjTdcYkszYBP/wSIBF9oKKXK5tQ+vWebnyfrSd/SdO7+iBhpx
vzr02Y4p84Iegp1Vgnc2ZjJf6iM8kV6L5n+Q8osT+r8s6Qkv6eVXqlLn0jIRYfw3SlhT+6FyNDAZ
lFv0KAZ4+owp0lzST21MsT6PAeDPEgGQSsxsJlo3U99oiT5/AhLP6XohDK8JbuSC5SMF6L+CewmZ
rdJudA1LUuhhzxoqaFagqhBbbkMKI7WY+1bz3/hp0aJqbASkxMd2HfRO+MeWWF+kH6b0iTw+Jj5U
glMUyTluRzY9xEq+ZwQ5+cOgNkM8a0DGxT1PiBs6Wy3+XR1p038EhYEvAhTgoacGBix11hHMgDV/
nue7RSZt3KHVxrkRvO4L6pQ6dx26gduIyk/orMK7YXmQRvN6gCMOWso29GSGUkUipzC/x9rYTFo5
MJuPhxlyE+66BodHBuxe4330L70MvbxOhQuOCtGGXR5Mkg7qUvUZ+A/6ztRQtBOPX0KHNyM0S8Kj
zwoxK2kccCw/DyLTKK6NfWKPdz7dIw9qpnqfdUqKpcc87ytnc+2oT5ZMbhaIL83N7wdiUu8k1MTF
ys3ZW5gH4lBt91GIOrb4K5/9HkPklMpGUrEZuHdYPrBIwVUpEnWtNs8Kbocw3pj4KLU5W86LTAgg
c6jd6CblgE1nY04L73VD683Q1HymudtXtdhBSsFalEAD427X5i48pxavWBlfpx5dneHVUPcmKMnM
tLb/OoYQJkCcxDYyGQhku2c/WmKv7brESQrkVVeWfEFn7/n9RQUt/rdUpP59lea1kaEBQWgS1QqR
qnG4aSFADE4TmxwklNTCaShdBM7l8l6LmkEXXeEdiE3TEQjeicZ8Yno9HXmeKPOUPM09gCmHXNnj
Lw1pj2iWdMLZt/GPyRxLJTiaRuWsFCa8NGm4zOQ5Dws8me+9FDqK+/XOYfheQiU1I5r0jNUhMlZ1
v7WkrFMlKmN4t3NjV/tOfwvoeEOgHhMUK+aOiYJUHK9VCyu1oClx/cV+42hpAbbtdJlakZ9k1w8e
2H5w3bcst1MFWouJ3hykhubZXuwr7h9O8PXmymBODcCR4cVbkaIwpGZNYrxoMS13Bn/SITbW7ymG
8lttCSnZg6DiceLqUfS2c8YvQa+jgQCCIFQotCZShAvEJDgDsj5zsLFK7sUIfWPaxyRdEvi+Qh0x
hXe4gWZpdPEBr+SvP0hc80TvmZO8T5lqp1WnFy8NR2xpLzFD3dPlz36THXLKMRX9ITwg3DJ2l9tc
QU4mEvaCF9h0XLCsLuX1rBEq2tkWai4rd8SjjCP5xQK/rzpolHDz2nly+IWtCh35uzBVh0IT1Lq6
3lXU5pAHMFG7EIqm7BjG/wKZ+vUBxmPIBAbwAtzjv9gu8cga8vAvOv47G4flbneM5ZCwB/yQeOEt
d7NU1lXim6cKL8OWhnm9nl0RCiN0vEfdkGbrjdSDszg16Mjzh3x5DC7FUpSWOJUHF+iSKHiOnvTz
dMb0d40JqY1bcHHPVSnR0LuOY3Cxrd2oWlWw1KfEcgwQmc3y/5DCom1Vp9L57mCQ2bBKvxTXxZQk
fl+AdBaOLEBkDNTEz5bbgfEph0XXzylehvEztTY2NsZsBJyEXE9d+ZErE81T/I4RL7FVaDdX6LTU
FUyrFusAZYASFndiDHQr6VhTCJ0zdKLJAqzNscMxeCKRgvB4UF5z9UZzMaOjRXSMDcc0w6EqebAw
SqPK/uTUgyolsG7H/cSmGC8frsjswYwDYdK+7g5EvvfyaLykS3uZpXucWLRFuV/FPWNN1wrbU4K7
kLmcucAysbq7NT8QwOHSg3ySMRPcprNaYxpKCWTGkMVjAJmHiqPaDno5gzYAzthI1p+5agfq7DDg
gEGO5REu6yS2ezUHBIsCpJ7Rv3ZbMMYO5o5qEjWde+YQxvFb5QKeR2BDkOWHfdUjHbNlBq0m6k7Z
nZ6fS7Wbo/MAALOwPIRwMxy/FlQczO82ZE2gMxK94JIwHEy7CWBJS0ojCRxPd/Z551GyE0vFCQ3u
VA4AH5vOIiUTOSK6KOFFEoXA039BT0Xlhe8NrF4qsBIWz98iq1XYAZJ2L688E3Oy+V4HfwBSiHF6
mkvWW8pRJ7HygtpDOrssds0gp9aqwJ2AtnrN29OJZmv3kcTN0h1U83ucYcD59eE71+hRuxfS0xbE
xGfpOXJlvlM7z6MvDwsd7c4ubQOqMwca2EEtpqgt1Qs5Zeu/rEHg40KXa4Qa2pFkmdeMQM9JDw0B
djfKeJGwOA7Ely48noH5NJ4McYj5UvCStzCJOOIif4AUWN0HUnE+1lMiTeYBF3Vb9/m+QkhYajVu
3RAaHpQbIVmbzXN0JKFuR+eciD7QgKPTVAcstYXAHwW/v1e9QSB6/MilHfxyf+y9I0q86YSGaAbo
x995UiV+szZx1rUEwRTgEcyuaDlyE0URFXrPTusnAi5dH+dDTyRoPgtu9eYIMMgMQl0U5MeULEJv
3WOLczEnA3ad3xeF3AhSUufLmvrF6pUgNPyinGwiqy5cC5mGcBE4pPJzwR5SVb+sbC3/F42/iAV0
EXox3jEhly7xRiPEwjX8sxzYl9P599EMzOWq9onxJAjBuftgNRTAHhXi1Ky1v+4vk15NNqQv6xaz
JpkWkJbV8AIXL+++XvbBMuVcziCrAvVB39CJv4UmvoWxhcSmv1YUCy54TkDYxE3hcJy4K4TJ7Tul
FKjZXBApNCbIWCRinuJuR0y4fmWmuj3qH/++M6kn57YRfukRfTAHLXUNR0111hof8qJGFVHxvtNi
41ni2gvBKAvFyH8H7Uo0eFQJIY9ccuIqM0gAGSh6qTR4qwgWsH2cJSsBPHkebVvujPCD5xqZ5RDJ
1ExlOjCt2zq2pfsopXxFLi9aqurF69GzLOz73Eyh5DWkqWNTiG4+3KSHHVEvAFj/npCgclWLV782
ULc0CVNAPFxevz6uxYb8DN70ApETYgLFZop3FGl+/foWOwJuObRhJDZYuynqei0w9ql3t+fW5Y1V
qiNoIT7etYIS3RB8XbUQjC6q/H1KfJMRAjsjCjHjTfzoTn6cwV49yQt/zNmhnUXn1SIPYffTZtI2
10deXX4rQoDxxFG3AmgLad7gpLCt6sWlsli3zR+I47kZqJa15jEZS0tWhiQkPeeNlvlu00lk5qGC
iFe1jSA409ylsY5+lJSo6l+YC1yq00mc4c9FHNvQm9ctNiSjT5d5QvxOz51YNpvIeChfa/TJw8Nf
b0jS+fpUy2GFaP6OCunFr8bEWgPLAT7ReipkOP6rVdPSBcNWD1Y/3VtY6jDLixmILhHEAOn7tS9g
0dp8HFqot9KEgi/kTYd9US2geMLjHF2m0hxy+NJoNCc/Z0Z0vvnyGvQ4V2ekhD/Sl+5I+mlr14sb
rtjx0omvOSS7sD4F3+nVOOrksA3HtFtN/bGwhOpP1XbNeJakEe1LP3RCb/4QynW3+eDXijDwVUDV
aslzMd5utPXwV4RzL1qgmd4yvOtxvb3iAiGOFDhqBQm1ngXc8lNFb8+K3Mo8Ez9trl4mDwWMAJ9J
IW5+9HBW2YYt8wstPx6WTbfbAhIcxMkWmBCDLaG04P41vUsMHSgxdRFn30IEsznAUfx4+4bjQXHE
ygdpfnn6vPtSrOsthjrF5bNWr48aBxyhDbM8aSxH2gqNhNu3M29duQUqPfx9M31n2FA9gp2ryjmV
tBR5LH32Cc25a/flwty2pW7ZFNspvdAb6T9xFcCk+RE0JVmC1UZ+7cjhAGCi90y57eWF3nWq2nCq
DXaadKKYBKkx2gVEmwvmYzexBx5EaB5d2WfUXoReC/YzJtMNWmkckPjZ/opRraEbtwXRVy3194QG
IV3/vM9yizW3BLsYmXG1kSA2PfSkPvfZI7PKilfmCo0C21ykgzAcqchYBDPrOERnqEgLtipYmqgc
iGpOznyArTPvnjj9vVw0PmZVe86FuxVGgTGrhqKrQdUuh7UGXO+Gzl7lXSBPsZdFCrhJqUsZasF+
PE2C7QFLO5msNz6MC1/zlFhPkgVxx0fWmCjlZo4hfCZffUze+f1O/GNCHMMkq9MKycy4qWJUcVGS
l+keLUpxnfQUg1k28ZoSevVIacgVG05KBnkCWVvNCvkA7JboEvyJIER9ENuOPF0c7wZNpqMTvcqB
j1a22LDcB3ia/LrM3zkU4nERIjZWzrRUo+aRaV+aK7a6usg8evto8uMH0gr3iNTa6Ypo5pVx5g/l
EOvZmxqVEynwZ2875HHpQ4YKhuIbmU1J7rJ9iFB449LxaDJjv9FqzcK9BxxYDn2NQB4qL+TdSozx
0WlzHzbU0uey3fR/l2/3+hKaa0cmBqrHVWnhG0TKmNzkVhmzbJrn/sHeyTW8LomTIR9xSv5NFldz
yvpLFW/OaOE3Bxe4MdDcuVa6NYKM+zx1MH89Wmjyt24rMfs+elSZp4DCnF7X5k/PruwXaYwtWu1w
oWn3HN8E0RYMeNUHu1jAWCoHvSPOYkV0IEafBU5xpxsNFLofcWnEa4TXkzuyW/El/AvFtw5AGg3t
Cr7aiIBYi5fDVjKeM4VuRATPdD0Cm3XybJ1JzXFOnxk2uwvLVD2VcDRBU/k/2cV/oSy1nXYtLOWY
FfzY1QDmHibpfz6lkTDK3Pmt1t77m/9NtLir7/pEdsxF8OB6KjEc96IfvOIQgCDEjhNfz9zlL1Qd
Cu4ZL6cKJ+PqlkB50C5/v2e2TxyMbQpB7IOhLv3kSfVZ/0+/8a0L6TsCxuo7JXeUdhM5yUV1Udo3
+E4gf5S+mh9U26PRoq4UFnTwn4E60vYRKux+3msIhuIhW0M6ddOPamuUTcQMEebOIYwbLFQK0q8x
OhmvE94UqMlvfJ+3tOHkDUDwSeR9bTfsFhn8tJVFNc9bFNFi/dA8tqYqOGxQrHLgoyVWWSiuTelT
RNwxz2CP2tUyQ37zFsi/1rswTfBlG7Mp0M8cDKENCZ8R842Z1ikCPUxiaqWnwTNwTEIsavugoWHk
EZ+WSJE0oiRJxadfs+pfLnIz477chKDPu2ceUsHKE0sDimfg1EZUG99/t09qcNqKHKOnS6SgBI5K
8/QjiL/bEHxMkk91+jIs/AKCkGz5adY/GmwBfV30oYDQA9UGQufiKxyW4IJZA003SOPivdDi/bB4
ILmHtZeEoAC9tz1RCxsjM/xyFZr8d5HyxrzCZusxeSMidFwGyADXbqycjjFERx/JMqtnAN93Znw0
6PCQL+QetA4yEqBfd/OEJ64TDBpOoo2ifeqjLEbtcZaChjdWGTtV5nLxXXbvA0p0ODAk+LBfOrW/
T5E/21csG384OduHeJrNYlYl+ovZnXrXwKhu3LNkPGdTNuSJ404m+CYPNludRaTa7xB80JrrCghM
UrioRtHcrs4lfiEblOaR2AAgLtujlS2vCR7D4+NdhNO5z9Y5AJf0L3+PWGqog8HAyxFYRA9wWV1G
q/O7nbGicAdD1jr+lb4hPmg3kufMFWxD16Jwt9I7I5YrSPt4lKk7fHQxKfA7IbBRx0NFl7BQvLQa
3JI+LYrAiJ1djQCje/ILYk4qGxgPS0vW896PH+3h+MP9N+ZfGp2mW15EWJPEuN/YidS3qtpfmzrU
1Oe+E0CrjGWiAWsnd9qSlwm0fAXlGwLb12HRaOtlFfeiHLzemFKIaNF2r/ByRTekDAGf8EFCF6Ps
vD0GmaRrjl/+7dkWivguhrgi8zBHEXYH7cPtQiph8cuQnznp6K5h9P+AvobreMnOPidjY8s7ri/R
bcATRkJUGVb/gBR18VVf20HYlj551fa0ZhicKfy9wFlBxvMfZpQmzU5vAkMlV0w5TNgANHsIzu4k
JgJ8kKrnEOKOyIRoODb0aZVnc8N8OwXQx1BX5M4gR0n6wHACBZNhn3XZ1dJw/T+DVEuDTeINK/4O
gcZmJSSzDE0ElK3+2sT6Kz55wJ0tF1+ONWTPJEP8Ajo6EjhM6RovX0cf4Umu4Rqr65YsgFh0gVTh
mnKzZoNyljPdMGNy5Mu7bViiuN+tbz3AmWf5WLRSSR28tAZAsLNV0g9b9UFJy2nMKqmQ78CU57Uy
rNH6vcmYV2O6htuqfEnsCQYi3UwqmtRHGtUW9x7jeiYap9uiczMleFbTMtjr1TBUnN00zWohRvU3
czb99ZG6YRo5885fkb9qUB+xVRswk5rx0+8LJDKun5cnf88AtAYzCYFEp7pTcVUjdy5TB7Ti9n+S
XQVYIDwUSy66ETbfKAluVWYIYBBHH5+zmzHm0gWPlKU3sSEG9CkxKcoJDoa/oU1lytVigFP4ZLH6
dT0X1UwuOf9qqgI7P9CF8CONVuZhEL8FjieVEXbLgjh8SqvmRY2UjO6QG7i1ANthXc61RYTfhh4m
t5jAxU9N/TlsSL9NO6tBwcfSTO5dG2YNKGOppVmtULmUdMh/oeylG0mwzo51P43QigA2f0QXW+bc
xG8i4IngTN8tUv2xYaoMZuwU0VwnkEjPDgPVJvsxFrm3zyRcv7QjQDvJ1vJmtachY4F+8C2nee6Q
oAm4H/PNeUVb3KeFZ9HZ/tXDK5/VUrUKOuDiAZhuRTVM7ciE81RjyoEsbQyRCIjW4mK7UIvCFDDG
w1uddz1bmnmf4Zld1kS2MEZKRAiRsNyWF/JIojNOs1qUc0mZSXhK0Gtf70fyi5xpg0l6amsLgH2J
wgMAQ0nfwnsNsP29gQfASG571D/HJcUOPF5nO0Qt8yIqFJuZMJF3l4aPJvCoXgnzgTur1llcOcs0
WXE+V5BIgvsg2iPKUCeWpp/zTmb/1qMEUyhEMH3LQuSU6tpNafrfWHAgEmLWTlpc7PEsUL0LhKQo
0c6ilxJ/wQr6KK7Qmi5Dp1hAQ7nraHDEuf3RqbwjS83OsMMfVsaMjewl3PpIliD1srzWYKJX/vov
tShusiheX9EvpM1DcjlqIZbXlfETF3PEwsZInHpmjLhGkitPuerz+T64dbD3vCIlgDtsRd647h10
uW331ozZzZzdcZAX/tddDe840OnUaiz95nwkW82MqCDED6pbDCe6GD4NqIMRDvLNLzFGOMILHj2z
tBMMJTxdYnT7y8VSMXGXpC15AfjPrV0jDq0O41oTjJyNulyfbVErlmCOYOGjq6vutVWfeoLFYP9u
e9a5QxBYERfdjHd7atAGrOZk37hhBm+sdD4JpyUHcHCq5sIpIUPjSgfSMPwWy9Rsc/kOFAiyfGSj
OCFBv4cQLLK71Z0sN2ke0wsi5FE3pzbZpH8FoAqpCJpfLrSm7IxiNP9cfrtjMBecngZf6LRVhptg
Iv3MjySegG3ViTO4a5uRuZ97n68VfLeAYQkagTj7w2E+r86P9ysOR+VGAdSDZIBH+KYRjV/vvJi0
O+3wwx5gkYqv0nDapyDbvvB8Hjn6t23VGcGwl78Varc2kCS4rHWvqChVXyWRxPWiv6jwbr/6OoTb
ImwtCNUljP6DUV3mWiAAebjHaH74gITthKqXPVS5jwRazLJx+oXH5d4gYzpvsGe+7b6Ve0bFtY/m
+XulO1wX959/kiK/iUrs9V0JSr2NcjtKUsBkPbStjIm0cAUp3ZkP6ioNUA5fX5TOnFDb5sHhTQuZ
3teZ//4meOztRqcRzbdt3hu2c/po41pzc4zXRNqRqxWKcaB3aWNdMtd4w0Ylow523KqVv345c5gl
CXwHXnKZ2lP29at0uyoK81hqr9L62ux12sCgyHRsF7X/CMb/GwycS95wM3kfgCQQhyC19CuShwmE
iSKbn0/ZUXhxQP7h/6lfFAb/MDc8aemKJV/ANpLaW7XanUK7+bk4EgwPJqS8GiWrcg78tyf3G8S9
EDb2sREQ5+hcSeDc3vEY0iPt1MV34D94D9aKpSumGez2xgUmMRkyQII97584rSIyz8wcoY+mAQqE
uYTaq8j/zYZGpTQip3iZHvXTTOTCZvUB+m17pI3j3/WdGG9Rlvt0h5eTK/05rOTZujD726z68TUL
GQyGBdRhDCM1c8AxotwNcCygt+qcL+oPpLK4ShP3KY0nRJEXJDv9zXlyeg8Du0M0uDUH2/8ppwUE
XL15PRXv2ah7KS2FztNHT7IBx7BYR2OVqr/+uB41DlLDOgaRwrwtOxKgWG9sXR0se+cPwp9GVPCN
0x2J0C3ifaA31BP5s5OjqxpKGQ0kaVnma4p2F5UZFKkHoNPXj4tyVXM3F4oksIihq3eJOGYYi464
JrjO45qiBAgrZy5GExK7TZxU9hlOyl89oJRWgQuCRj3xj9tDkkUtsMC1nmZgrfEOyfMCIhPsR1I9
1Zb/t1+gYh1nWnbUYJpuydhiz/YLV3YU+Q4ALoLi5fbZqSYEKzCuhEz+uWCOBrzliKT380FAEgLP
oKE3PuU4N97Gd9kkSQbuMPfgytAH9Yj79S9vxCyX8AZDtbEFdIciWg8qG9txiu0SceIteTrvu7vw
8bKyq5Wv7P+9krHDgzs2gWDlJ3ItLvDbgJdUF/+56jfR/FKwrA1UkE01D+9C/L8uvHRP8EQ/kIOc
ZMo+VJfGeTs98iTacx94xSnc+4A0yxhF1uIySnfpcD7L8Fa15PZ0WuQeKMLn3f4VWdlFMb0a7UCf
4tEq2aAhG9tMnoMusNQjDchwDfEUdJvluqklmpBcaam+6PaqYEssgdw6mnO8HtILLLAKOqneqUl4
MZQNatrBjTPryOsolyiTVH2Z3IoTAGmhYPPpPiiELXCF0Uk9gZ4vQ3SpDyp8Q4rWCRB5yDhmgrtE
VrTMilzw8XlaeUgkMiR7ke3dbn1kkYHbc6XJHuroLFddXBkG2hjmZDMd2MqInEqMhce9mT68eknA
w09Yhlfr2HfoPtTE6WCBgeK9FM0p+qfe367JZei80b0nlpIRzq2K7k5HU27k7Oe5s/g1Ex+v7K6M
9hOY7WiK++ZUpjyGtyAnJs5t9CPqle06nLLlRwttQfqQsQtBz8fhf5TE3JEpmnvqvHKyIsMHWeLe
oWEYCa/enpQRySK0Qa8bvDMovU+0LPNB1VimB31Vq6hnSra15sEpd4AAQggb7eagMC20hEWHo3Gn
ErveqYku8nEFkqMc2UjBt7U/FfF0MhqNrrvFLSiTr1HpS0AiAyCpKAhhycBzvBDSF45+MCdOzXol
Zl0NjbCGz0mQYLCxChsv3htOkSjos0dCjTdAetpONlWHcM1clSxjRWhmMzXSQv/JP82WOH5AS1Oi
4W8kUdh2Vxzo0w5zPzJ9PfpTiyZFmnhDriYKZC7yf05EE6kmZBW1MJzuayz6Yu/Q3QrTxdV5VbWw
TuZ/zpplEwfih6VBQ/YN8cFndjeox2pwDuSeawA4UkegJ8bXVQgaAp+Ojg86TqC5Io3MGZ5dfN5U
jgX79Vt0dMYXt+OH/9TJFlzR37ArdwKkNo8UBqMBRRjmfu5VkmhFF8l4UtEgMKzlpOUpFVTFXks8
1edTDRB9FWfEdAz+daH0F3uPzTDcMTAANFP33APe55EianGw9VGfDy1WOLpnbc7VhCBCgZXGlwjE
iaRfsyr6QNWNGgqKYWOTAq1pXbwOTBpWpN/qlYyNGXO4AtsWi0bcqMTB6nJ94EWdzElMHFaTlC8A
d2QWnAUZHeJSI5EmRdIN2lLzpK5yk2ngq2Yy1awvfkm1PhWHdg4Zn02glZd0i61oWW2WIFKAhZFP
R2E9xPur740JzvNwX0RmejEywyVF9Mh5OSCWRAmd9Ljtnu+4dXHlYaRiqA+tKBY8PcoZAhU2IgqY
j+YJF5MYuZQd+x69VmcW8J2JrFjNIy+t4xFmSitL/fRGs6pomc8CPiqXKkv/4zrc2aav/vCarJJh
gtTjhzSzMxquY6Fz4vSf27ZMTY3XeNdWmpYBlcp3hgQi4PW3vQDArv81WIyS5QUx2LCc8FSlueE1
3fNSXYd3GSqUjeEwaWlHoJeD8FCsur8IKlfYoKgX0/JD5wDgBPM/5VXS0vZvVpg9Ge69/6sQuJiY
tNkLgFUCdJYzF9VGhu0A0jstS0iBvtlkKyiOB4L5YIdDirTaIRpOLVgWJcvcTTSf11FMWW4RUXAA
AInDDMKV1Q7UumehztC4i3Y72Mh0aIFD3SLebCLgDZZe/w1PrvZDKktN4cSRGOVCu4gRZCkbFLI5
Xhhf448Wy9IXFlq9W8AQsVp50wb/UZ+UNgbXvmZEzzkdqFPWo/5vimFM8yhnVdlH5+cyo68dePWN
gMkv9SBgqqo0daNccLCzZ0cDukeBAZRjSt7kV4Mk/NgTCexosjx62ayQYuKXJdAdxn8s4UKDxZqo
YePoKidsI5mkfg1ScNJU7eiwii5cByPZNPKLIrvWgZ44hHdz7Fzv/O7jw743bhJktDUHIP5nL0/r
OBB23fGnDknULDYwac+1kVFtIhC0boKFxkDTqwa7qx6nEqnfQksFlqQZbbrLLY0MePAjizQnCGrC
XGpuAzDPju6gUIwin3Srxq8zigrzJGaUA7r0O479ySO/07Hb9ohe77u8zSl4LPzPOpgrJh90XEq2
kN1jqLnGmWHTvLkX8QCWKN0cnb82/IK0okaFkvlFh1wjDJ3k5a4LBIxCov9P+qr3qYNAN4Ad9cuA
f4jTq7eH5WX9og+sfqqiJUUqh9JT1HRAhwdGqJ4cUb00tci58Bnai5wBS0N75LMBruHjtcLgZbjq
JIL3u82iONn2qXxORFZMgdHvYOVLA8owcDm8TOt58vkavJ6yOPb0r5D3iLWU30WMv1F4WlKad9xo
TxigT/kI+JiqDuVMHnSHWnv8A3X48YhwUynih86W/Ex0xchWKWWMhS/incArYA7sVF/7eebTl5jZ
vkK/tgopNmga/VTWP05oVJZmfeUybeCJ2CssvRByRxrorsLNOVB4+DJhB2qLAcXX43JIT8Q9UqPg
iyB+FL+PyUqiY2mjcv+owcyzBImDdwEmtpvQAFqpzDy6U87vEj+kYe6OaU7hSFsNpmREAjwaV2DN
PKHBV3uL0bR+NC4ck7y+Z5DeV+8hzbgAA+5111wLxWF4VK6r4CBarnAH16Z7+LHkfyHaRrjUIP/G
/g/thPje1pzaCcdH9ZiTZ/IRiyYWhArsFVUF3unl+Ne6aL9fJMkEHq2JatXtn2vqFy7zOPC2b/r1
IzUoP+Q0AWunjskF6vkL5nB30DYSsn1NzQ9lXLFexzSxtVLLc+Np8uQfeLBBswUdQK1lFddIRart
NhoRs85iYIm78RH7lHWS+CHw0SI/+A4FiWr66PShkWlYS0JbDUCrZ65XLigSQYzlqiSvC9g+SnFt
MWsZDGpfYDB1ANI76/P/cKa4PxfFcyZ8YofmHHU25taZGul43IW9ZZx/+Da/nu48WfAcBNecW/Yf
AGXMzbZODRHpq6GvcMmU4z0kyyroxtXSmvNllSdgPLofp6DTn1K1Ah1m3ORkeLnAyBzXP50B8U1B
PuLJNjqflwZ+VQ1oMfj0R3DSmWuq3J5c/uyMUp7FsJJpd328Is1bpM4YeRhFzqzDxsr3njqZtcGR
T0Zk4uRhX973x0/YX77NfCHWuEglrKsqus/WMJmoPzGLJ0LdfqlekSWMlqiw7ruN4Gcy2T/Grucu
1i0dC3dJ6uTxLtVR3zKl/lTivh9MtpT3ldHL2wTCVIIsfHDnx+JQSe09nnObvFxnzBtXTb8zJEIu
soVPQaGx6yuRejd0DnVpSw6HK26TMiXU/1KRGlQDT5/+R3dPb75BJi9XSvAcCWRWdJwb3fUByzGd
oAU5nukWSv81r5aiVsLg79S6//mHwT4jHUUyUoiXdYW25IgkfSZaX4RG3Cz6xyajlgBSbgHgk9J1
bxr2xT5c9k4r6VqyOiYC+wugQrYo9DNwYQpMKLgJrV1hiNu6hC7zE3AT5YRGXPSnUafmqqzVkyG/
s4/rV5M/zjAKZAMKynzpd/2S82fs7cfnXe980bQhkR4tT4qoAJisfn658D4PrFL4AbXz9TTNnKLR
n5v2x7NZsmgPjjCOZYeQmtjaASpSUHfRrAZbvYKVSOMTAiHBjrf1jZVCAl1r6PxIbP6aGbGll20m
z59jkbDjEP99ZB2Rk3H/ypSNZnASUOfeaFQppXSiLMfAFJ7x7VCtRjESJ3vnvjBrDVTnjefeQK9L
DeH58EIaYD2lrgxdu/IbVceeMSTbEaF2AWjH8P5G/R+MwkOSAMyDnSfFwnL5teEYggGi3t/qGg98
69b7yGXg6Cv0fDekvkhgJaBfVHcBrViP5R0Xh05bEcNqFqMfdWz7NUJvILUfPdyRHuIVD/Kzq7oV
d6hxrWpkxRx7znyC24E6ddYTwqwn89S91wz6H/uBfCQKwUKeK6H+XQQBtmP7giMGiIoezaHkgPBP
QxKrC/nCAyNssXaUvu5bKsyZTSA7Yh6ZRpyw9EuW+wMu032gzzUtr7rXr5cL+Z0k2NdS++XS8uah
fXrxQ8UosU8Nxn+LOIkCbdKlXdukHw0shz3PAPPlFvh5hMMajV1xmiVFkauKsvE4cpddplki8sz8
Y2o/B+f+8D8sqUKOf+eeKdY/ESW3wLNAdbKygW149/9GrDV1EjlC2i02rbZaZed2k5CO+hYDCDzV
40f3eoatesqoeeb7FxKek9xXs3PCsW991asruG3iXgG/otGF6O3bxyc8+acsaVregbNSLHmaKQzc
pLEdH/aYiGhzKuykTD3U273AnvPxXS+aJBeG/ieKjYI02rG8Lcmis/dX05kq/NJjaYqAr2dRL9H/
kizfa7WYYv3pWK91+EjZM6+Wa6i63e8J1nAi1Ijw0kCFIOsPuHmoOvAagUT9m+mArAg4wTvfrp8s
Se0CSL4yCNoSsiHKtUfzpJPaFb4apjIn4VB09vLGWvvQe0PYtkqhgoRdry5FIR2Si2w7lLkXCFK7
2lNkLQql6jzpWecI6TuK1BHrOvDz2jOXx93zHdv/IcE858hzcdFex3ZWjRWeQjY/pavfEilpHSk9
QzejPii5FL/3W1wvz8UZ8MScfmgpYMOEc7iTI2i8114fylLYVkaHfzeBBuMpvfR7WNjAY+flak6a
hQzAe+EqbAjHJhbCmk57OELYAAEedEnbTOulWYjgi8WBk+tmDiW9V5TXE7lEkhwb9vGWpK6VCruk
xII9SHyVydsjFiv1RnFbwCltIAfOvnxE7o/AOx4wJgNDRqx/CVfX0Ff0kfrBD0vqKg4ZP1nLmTXh
BEVpip9lMLKcSQZ4bkcyBTUhAj8qDb61p3u2AWZCYUjnf1VwG0JtGbkexhn1Lc52AU5FI8hXEKxf
Ka8qUo5QkgLTvj/IGWVJGvm00TbwIpkX8wygg9dzE17R5YejDUkdS+OHA1THTgF2+5gJ6cMQ9Uz4
xxtFwGYPMI4/t/EET3XnOJnodaTYmVFF9bpDOyhdNj4tjeR3ZIi19qsldtvkfpnG1pM7NAgT8PE0
Lsv7DpxLTsyY9MUPLOteUDRGU0CwmpuQQ1F8R4MvzHTpdyHFuAXYQRAHq7/tGnBjfFCs57Ph6cKC
PPuRQZ1Sngv9GFNjYj9T+wgWUFI6jNwDjqTCQq3UQAj+vgChpjNEvX+HhmcNkzTd0VLb3ZN0MPpj
w0NbUCiYCyw0TbzXgVYmaAhglC3FTX989x7pZcRoYlxB+RDW8Y0zqqmW5r6GYYqPEJSbka+ns4Z0
pix511DaxwQxt6F5skbpXaiC+AD4uC2LJaBPhpEekP8Jy6LcT7u0kHgNmv9ufUFeV0PGYa/diMeQ
cFvztmTwoSC2nlBHYFzMU9c1irsEM6YlzNooKW9/Y8zAkDW4pms1NldDyEmuNGwzL9sIPjnBiq/x
kSXHZUV99Yqr+eCoOtlxss9spNaS8bXJINUiUVBH9V0cvDfibrdAXXsyz21y5EhTFMoIIyee625C
0VoadLVLMoEPAQebQV4rA7a4r20gKj7BWxnPnv0CtS3lTlPbaSDRRBQiAGTZhu+29C4moksqIMwb
M6+WD60DqUpTgRX3DuN7L7R7RcmKZ1KYvxOxfG0TQNYChkKb5ODtUxm9x94Pbnpt/94xrKJeppOJ
igD8LhtjxbcYq+ITlLCdyBSTeq2swVQb3VgCU4CJ+RkC7M1ZVMZO+WOVAhNpfYoJpvAPbfHqV2wG
grzfMhLAKWLpFNo+KiYirGh7pzLDgwKuazvCVkuiOAWWT/s5vFnKQmfGl8lPBz4r8DzlQQCRZ/ee
Y65X4XKzHyBtt0rZn0a9LFr64HWPwb7f3Vtz6fHTqs0JB7T2SpWRyms7P8EfnUh+w3wh3RLPV0gg
SfXw4RvjGscchROCoHGBMiUEq+wAvYim5HJG3vpZfpVVR9uLPtAXSQn38OuHXK1Xlw1pCgYS42aD
BUJfhrLHEl8bnZNJANrhofneQs39fh6DP5OoFZwOjW4BeKZ0oqFYmcILim1I2TKSSdbPxKfdUrjL
xVyWGeon8wDI9X8l0IeAdsMD2WXP+TCLwhRBG10b2ukogJosikUN+V/4ILF9RE8vvOXwOxNV8Fb7
MZBIRr79IVt6/MC6mGUV6LjhSH35ypUQIYr2Ov9De/OJTfcq/IhHNfSBHXY7XU6zBfgTLwoZ8OfG
0lQnS1gwPlji8sCJ7oL0Xrl5pav5YYPfhlDcu8UDDoKvtGEz5MmG+CF2/UfkESOUal5hjI5ROHG1
DpqXYp7+VXh2reYyNAotWIskAfmJwzQZDnbxECUVORxa9SWHrGkvAs7eRfm8WteQlRdwYNjyINKA
+BXqZZ4zFpr1cam1+F0ahvyXF3WBlSmx/KxZkwxdA/75kCu2ulZfLE8VukMEbdo8Yf3vZd63MEF7
V6w9cccltzX8x6zIYHMZUvqWNJOL4FeUbAv4ZduXx0zlCvQ/qj4J/rdI40lOx0FdSueLyfx0FEtS
w2fGyhhYnP3dajFOOpu6XxK/fphaxeg4fsa57dy7asfQbXCZHPTSOl/ALxbYAW9ehJu2700tGrgy
/GNl+zEgE871RKuhC23JmJuC1yah8Pp+Prz8/GGw51U9Up9Bnb+qD16F+fPWmgyEIGaem0MqI2yH
E0omXA1iA0t1R+dDeDaKV4tc3RYuSX0F8k/hUKiAfDuoQ9Tp0jlJhElIMwhgbEfZO0JhZ6LQLLpf
yShRfHU1jjG3FdWda2L9XkHYHy3wtNhmUNNTvwNgDUPieybBsckm0n5WoFVXmiVDeB7DixNMwM7k
r+ksacKY+/r1yvhHsEcWPLVsEQrfMBeNyFaktl+AxvvYBDCtKzVLytUY2MhXpkhxbAJ8JJ1cVcoy
S8FEt/5rjumuAb+GTfH4fsnImeRCttzNdB82vp6zZwtxNTOVJFEvVWap0lMdvTPtRP63LpGhhPV0
DMi9Jf8hfSOP1rFix6p5KBuuG00kvq5b8NJWYLN/MfjbHD2euov6wTnt1/QI0vbBDWGSmKUg3IHG
d4pazLkdCpXyng6BbWzNbGvmMPdlHdG7vu+E0bFZIWmQrsnX/sOGm6FgfY3YDXN8EP45GOTvGu99
SjRcwVmQjEysXMU+kyTQAZJneV1YNi4AxBgQmQyYAcyLLu6UH4VVfrg79QJT4d/vO5P6gnU3tI6v
RN3mdZv6ad4xa2RHEiWtOMcs4Z9OqMCmKSUnLiIde8ZPZJ4C6pwmHUEAY7mz3DVCMdrIN57UcRee
3fLUI1MCfwaBmIMRUjrubJY0jBCcBBgx0YyVuRBxBDL93/N5Sy7c4xGX0gonomSy/buce1I0A8t1
/D6qRNf07pWUPlRsxuINIRRwwxVP40gLCqAlq2EvK50ri2i5thSU5F89sLUxJyuCFQu1kWH8/f4v
5BFUAVi2GjIzXl6a482fV/b70ZqVCiSwpDNL0lixub61OP28/dU03a0fS+CGv38RczVjjRu81e4F
F3w1lX8NlqZWF3iTwSDN6yi6wLhmHkSvABvHevNiCCinIC3zX0yW5QJcz9HHe8NeMeq/l+0YU1we
Uutc6pjpmp2+Y2goE76lBgH7cS+xWHQFSEM5i8WckKVrygKNNzr4Hn/Ok4e6hw/fZts9GaGYsovK
YMcPIQiS6bZXTm6fN0AwX3u8qLxG1TVF+kCo3ohVlhXN/UyLkY7V1szKiggdfSZzSuetJY8b1VI6
7nn6W785hHftoYtV34O6CSyoqQZsLvIfBdt4mUt6uSXZSZw2rCI91qGQdg/slx6xmhdkqn18j/AF
yGBNmsBDT6op3Gd8NGpFHUEuUEmkO4O5tcEjRFL6lldxvwm0enQvmZXiYHhePEoUrvIiiC/IM15h
0gjIoQQIXe4t1kvXHXnP14bgi555RS1My5a6BmReqb5xBWMwvi8B4NeiwZ8qIKT1pbZMFt0hyfAt
umrAmdoCb/EXoigdUZuBXVVFmxtlmTUOCaaNLJxllN7HVfqvYJJDuEve/qhP7flasNNsvweGde5v
RW+np+aKjCYmw99xoMH1C/dnktG/2fRCfR74K2Nkb3m4bhB0MuN6eRDzptVlLx0W8d8kJF1bkY/w
ejiKODuXRtwv8X+/kUNUEnh1FYc9HbY0c6T+7bahS46xTVURv8EL0g0REBSr2bju7842TaFa2VI9
pRzbdQjwn2iJwuJwWZSHY2lMrX1/yOH+RMAaYrrIzbiGuUffraMxuAW1zNDZUa/F4V/qTgkblN3T
1HAlt3USPnAX+35hnjkXJMHnyNewnpVJs5zx63eSmvlJaeBd8irRrm1mpZNGl1mDoXbuwU9vzwed
A8WNpIbv61Duh8JpzvUSnY98vM1iOfyhunAAKDlo+ctPIOoJHaQc2TGf4k1CtW4leKu6tt2tcAAE
wfsmruw8PjNfOUxY/8Sx9TC+JXrXJ3Q23kFjxI0uEI/HDjlDek3z+w49R3IdawbkRRYX9Imf4AlU
+8qzc3FjpLoN9nw7GWnczf3Kq0AA4KEGnO+XQMc+JzwC04umUFnYSis1iMBTOSA3wRunICqxz2pB
RHX5hl0I1S5XZPzu+bhiG6kmoHnjLEZoZfBYpGqGNJqwpNYeXrnr2u6y+yRqzxIYIfu8U/1f+LeH
SyXI5H94r+gWYnECDEIR96i9RNC001RZBPrXmMma0oDzmxeF6GYDZ6mDix2NUmO3M+TRmRBXeAkX
+ZWd7RR4DdRUjsYXgyoLV2ZskRVdIk8G4ub0skrGQ8QRYgLMAf7E1ZQicYnOs+qS/8/4n1/slRmw
CwnpaVLy4TnlUFKiWnH4XnqowCx/vQXXzcaucRX+XkRBbjQjW04FiFj6Hb439rEiqFJPb+/R3nNT
zq+nkOtjj2akVNuVigTJe4RlBdg7B6qc6Sql/dgAalEiaTsBf9DVXJH7L+PbgUKAguVqc6BAB0er
k2WA62PeSUFHaGdvRpup+Hva7Y1blVZYS97ycYKjdGvPbs+R2bBxRra7IMPoQ5a9TjY40tR3+cS1
cPjvgPofzk4ZSzpcBgscXF9mzzq3UKZdXCeOFbiwJsfkjt2/wlHTJPFMbHeSxPSuNxh6/gZfjrLI
IXKL19hTM7Cln6YLzwVjr+kG0Ez2Z+ct2r0HCjsdfAn1sAOhDhYV8+RNEMkxuHxiMgzeUHboLt+Y
Oh9jnW3EqXudiWI5i87kZ4bZstbt7W8dH5n0QeKr0I6hZ9owwtLatlq6oEJDHgKt6clYa5bk2E/q
8NwtKFkT8gXKZ33OBjvPZx2iWFZrTgIvt2o/wJ48we9WfJA2wnA0vUHW0OwVAUFBsUgQiJxR1WTG
jNYLJeoCZaAoLf61/v7ye0S7lVRQiX2jxzbnJVD3AO4LgQekqNBLQ++WPQPypWwnx6S2EKkrccsm
OW5A5mVm0FuVg4cc1c4vHQXwPqqJfQ9lt0GZMlcOBs3t3p9+jfLZ8NJe+FyOU3Po4p6dIi+VgHdB
cPWqs2qX4Xa6ZyyuKgrXH2etXAe4VmSnxrQb/wVE+kulIXxA3YOQ2fqBJ4x/cIuqZZfWhtnAK2bq
OOI7Vk+N/WycUlOfoJibw3c8Ou/4IXJAWBHuUnXbFvXyTodXO902uDz5Lv5nBCwi9C4AvxqndZ+o
ULsxsP59s4ws2Z+19+II6uBHa0Wt5lMAeeZDqi4oGfTkG4LpEngUvoZEP+z8oKFw/HDsP6SCaxe4
9gxWhnscQ+60qebAM+zrUExNA9AbT0jBKI5sSYakR1I545gu2CD5tpRFdWk0pmtpr3f07MSYPokP
90nkzqaquPARkPQ3V02dVcNVeyxJMBwUTLQ/Tg1CzyfMczfOIsw53s2RVN+N07LNBcSgPhtuJ7nT
g+30c4JlFP9AOM9Hhlferym2henUliT1h+53AZUTfAPtOfkcLZfk4YR2aNAjG5NDGLRJxZJYuKkP
8fafXXhqWAodY8KDnclVQRk4B3IRrghgwakOoueguUF0sp6GHTNLTdcAIjgSrxT74f6Zl9g0Ej4z
Aybe1pfjiGaWljiCZqsU2gpTiqhdquEsJavVSmZeGQBZ3Og+PCpF8cl3/0j92iqMekwxEM9E+7h1
Btl2fp6hmlm3jXeUCg9h4QrIJYq1Dga1pnxftaZuf5HJizysemTP8+4YZ0CJ3kX1Bwsi7fT+X4Sn
f+nTxi0k9mKfMFiED+VVaeWcYm9xfqEKIjVRfGMNjqtDienEcOiC275q6yxCRJixiwWbIB/0g4yG
W5oy1ixepjeOdaCNPLfkDQEU4mdRqAKbsaNmJ0G6FFBC0OSm3v+cK0aj5EUI7iLF+vSNct3K7nOY
BrOaHLg55jpc0mJcxDTpjYgfAWvER5ib89sgG2auBhLa7AuuD3nyigWe8qzlU8TWezp/vlb4/piV
VQ5vqlr10gL5ZILCkXgx4a3jv04p3kvrw5tW03qa1up2w/LIS4G4Wrv54hmlRuw56mwSxfVBf1g/
52TA6aHrBLnx1GaQZkx1g8oM63DzM1mFwMNxFgoAb7+Acjf6oJzjA79HrUbS7ANTGh4yRTNwXtnX
3+69E9t/KeOW5hYNbfvwhzCPGlg41ZRDKcjx7EpQCUyYroPPJ79Wd2SO0naF8oClSAV+IN1GPjj6
GJuKMFHrlNLKKYx0YHzip8FHGjm1YRFSpVsIvYfLZWPD3LM0RV3LBNjAbNsPu2pdvxOyfLtMs3wH
Yamko3u5XtaWtMyf1pRBqKEalKs97REEle5QwUVB9Wns0pL40vPZY2Rr2HlNNZkBWP2ar6vMCM5f
FO4oa1v+933gQ/1nPA6eco0FaUhY1c1RSSSUs454HnvZHed50486BeYNEiyT3IntdPs6YVYyqwDD
OPXXUY/wWLda5VeTKJ3DtX+yXFG3FLYh+Xh1ntayO4AwEKqAUSfsW6R1/HokfWjGJBP7t/z8LJ6d
t7Lb/HEYkhSfl67bmxBmCfftfOtNtz+af1iDKcmv1z3zqgNzj1UbxxF+U92UEsQnd6AeNEHQ2EPO
MHBEjdsorU4t0ufgVUlsSxSJYL72yfrajM+Iam9E4N4TBtOVPN8q9GO4affsrUwvq8+U4l3k3Z2V
+RdOrY/aDDrTVXJ8WWD2hoe9ZTCIJ6mhlkGkCW5RjsSER4YSNcDJAu9BHN4PA8eS72IqbWU4Yq3D
0I3DQUt0TDkAW3/6Ly7vgvE9a7evbFC0C/iQvciCYtupUvnt5/NC13Df9AOM+/4Tw1SoKLqK8xBr
Lx0eBz68YkioMjJWmzASh9adBbjnj1A4OgzuNHtzvn98Tt7KEIPtS7FA4W5QX2kUrfKLE4aFbiyT
WxqVJJYgzsFsGBsnjIQcf21E+qHQgbdf
`protect end_protected

