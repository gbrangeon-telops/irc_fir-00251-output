

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
gQ4CxdvWgnieRLRQ2AMwpJaA+X4QUP23A7mcpTzLH1nina2JWDwyro/SbR0koY81VxQ8tVNBYSg8
3s+EjSEjvg==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
gPnHmBrjBHDleV2Jfu7AAgNyinLiMa4GswbueiHBD8y67DvELbF4ryETXsYzyyRC60JDgiQTY9xS
mNBL0n+tguqX8nripcl2WvUcK2rEIU4vEmrY5Xa0k52V9uCE29ruqODz0JXngqZvaosAn7R3hB73
7cI2IgLWPL6sayUHq1M=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
bim7wErRMWV5FSeSCuJLdGVUUYEH+U9HzwEGlgElmMU1LE1rxBL3MWBw6E1Qg5kGmxPZcrNQKg7b
PLZUD5Dv3VyvXW/HR3jI7P5DnwdmPcuCjrrkZwCh4jjzor7rIj0AM8ubprUHwkpicj6rKGNYRGRi
+lmT6hjwlretXlYwE1YClKFDSDei0UBfS9a5tRfCcNpmoCaImXf0uTOJ8unbujREQZSIp1snYBqM
Q6qvNMpDqcLoVSU7OrgHQdnonXWYqY/ILDCjdL1o02B+xcnkuGf+oGCDs8KSCPuzYvirbLqI8N91
feufkvRKEcc9+CQ7U9kVuEQ2Z+MB8XwJtiWwVA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
HhRynIQ+TRImN/1ISEgCruTQGOfZ7yQ0AeSPRr1UgeSXeBV4/j+sqUVwy6KpjxjyOB8/Up1pUaXk
C62p4kvtT61bX2llnNuuYjikfaIxGUWJ2S1a+GpileS7Ui7iwtZy8qreshTy7qb9L+4SycH2S0Vs
ofqZzZCA27OgdUdAA0M=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
RhnO7aE6HcfX9+ngWNOvpaRDGHOLotkXich9kwwYcDEBAwcff538vS/s9YC3iM7OnnDBzfIjK9PG
hZTnV6Wbh+heW3iD6MhhmPxC3a+3h3Xr7G6V/gV+8tP3qbjwLdyiI3Y3Tl9GXzeddtSNdvaD6764
1AS1CtRtG1cyGvfnXyGxmyDzJ91rqIOqSJbBOVjL0a+NolFyEU0BYVthKlZ39r7JI1kVtcM5XAND
LnFrRp5p6iEzVZDFdricPTs3V2FwNDnZSvZ0QADHlENUl1ofRaFRtXOEIahTDRwJJzBMRTba/K/s
3AtKBuzpWzTyvSqo+1PWwgrrClt60fAvHko0Yg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 12608)
`protect data_block
SiaVsfB90jjOO2rzCmxrlDXZbq20M4EFGZNbA4Y9sqWf8p8iVE3rm4hCzHAmMv1pKGvSfw45IxTY
XZdg8/u3TMrkcNeRaNx44uPTbQpTmd6lmFFpS5VYXir7bxrVAl4g1w2SH/uV2yA/+ZzPMcFkLqVJ
MFORnQH1D9gpX5rR1AbxWMu1n1mlkypIsqjYtpzOrQIgpk4V/DhWWm0hOBVLUkPnvCIrF1ZEOLbO
riMVdYElPrd4YMngi+Yfuo5g9BPZZ8acUrfA1KJgoKeiiVMXJXzuF6psleuKvZjloeIjxPrQsE0e
cIdMyMalZNLnKaXAgo0ZnUYRpt5Nddk5Z0E5Ga9+yAvXYR4A/+CFUNGK2NklfYiliqCl7QeceCjy
Ku24j4M6whjDTjRbhqRXTDhrIrA0mIAFrZJoUg7Vq6IEJWP3IhLivzGblcT8KbE4jE/dKaztCcpx
th3Rdp1UVpnpIpBn5KJ0KNqijzBGz4834+fqoWv5Tk2unxRIzWX16AH3zQ3+iDwUbZkkCVci0DE3
bZvZTf8FV1cMTBK0szFraIEdtKDdKr6mMRRUddX3HZTx8eHFCZwa1Pdg3ToYnmnJvfCZrpB+vMa4
vBCN/DHhWW1blN71JI7X4maqYjikqx/0n7G/X/NEsmA4dUlbBAAghpacgqlhXJkSvnzK3u0+dFEX
mwdU3ILSEwu7KaJcBT850J/IO9W7PdbBn6QGgwZZZVVWi09tvPX3FsNKUN4Q1tfzQu1GR7B91XA2
RT1PSLLYsxO/talWycVWP7L3SSZ4js2BANHpV+cRgG4nCIGfeCeaB8ItSJaSnjIbNriCryUk+OEf
uyfdC2GeBe9FoRpEaqjytOoOBqtv0T9VA+/XXlLmJsNWQjweGiNm62kMkWHtZnNV2WCF+anN+KNW
74QNUrU2L4AxdOtnaHvyulu1r8TTr/y90rHgHjc/nCDHR3ZLRXSkGLvi4ze/iera5OFO9wOoqb/u
LbHuHBHt+ZlACP//uVv3PfK+uCpNN4ykULnYMFzJ65RbdueSDm80vv4z2ZHGQwT2E4dWxprh7gf5
Rx4YKtiSQx6sI1MFJZJxDP1BIivLoNsg9NBPvBQmkzOWeJnf1YwSK3QbzpxYSDzlp9bDrYpuzqe2
+xby/SpFcDdQ0rblNhW5jkYbKs+i3XWFEUeXWp5POpds43Yn99ATVPyN3wueT+zEsFHH2LMEkUyb
eR2zLISkBpUO8systrxqZem1OueqsYG6e6rpHFJkVI2S7owUWfNz3qrmjBZtfP9EKj3da6K07Rkj
gFx0WsyPByyAK8MloqZTRkm30S23DLp4QNxQBYuY13YH6v+bWUuGUUql/XtFloWvgNz/2a8VRxQH
q2c8RApjAMHrE6sCw6SPGmzLaWuRMAJVVYi1GpXunnx4O9iJs4e+Rnq7Ji2DraggAJRaet1WdtW4
O1KsvN3tbhq0K4y6VaZZpC3wkNCL/tYpDne0ty4F/Qhk8zFBkKs4Dd1CokFTZ7omaSgRfe7q7BLC
ASlT4YOE6S6XiY7+kq9ka+mK8JA97Otlsd434I0wvL9RVoFJc9CoojQpCNPY/YYvREAhy0CBCmq3
A+GeNSHjagnGhD0l0crX8/v1milMxzVL9vWWk7XpkwNvKwno0oYj7xZHmSRaRYUcwHxzxM/7YIMp
f0MIfHpCfM95bUMqvsi8AtMjS2xk1prw+nmU0KZHm6M36QjpZ6rm7Bu7nootwpop5WL4gHA/BuOf
+nFFd6QXQnWRyF57LaWuand1MUZvWBVSMxMI5+LJSZyKidEwaG9W0ezhDD/X513lmjDASCZwXcaY
eAa6cYWcpIDf/zYU5TdxGp+q94q1yaYPGwelVh5MRDNpIS9XZ/HcPj/9jwtDfsYnfXyLLInZ/GFQ
2tcEbyIUM2yQJ6UFm2lBH8c8gOH2hE42YfTI+VW0oNd6tLNNZHlx+0hFJm8nlGgBEJzy2il1BLIQ
iN1MdXJXS01xmKuayjFebeHdLUD9PWBEGd01eKoGkY/08YRAXz9m6wd6sBqfCLtKcyiPT/54jbEi
FW0LDjwNK8OvyCyjYNXqPTR+3CN8Lv6JUqcafkY+BYV4rOFB1LgBp+8+EWgVken6pqf4OnwhMROY
LK0+OAKipe6SCSDzB3TtBWSE+x1Fki6e+ZO+/TIiBObsZe3n5bFj4oMeqtNoDaYBkrE3UTq2hrnJ
MUTvsHBZh9/UXUHADJIoqVUTXk0c9lwkaFBO7Sa/x9tLfjnoX2nhgAjLFwyGqXhM3rgfjWzkjXN8
aA/H/swIjoRaBYmdZP4Q764pNiVrd7TyLrisFO5mvVXRKvFCGamL7x1X1sOC4xHZ4QRbZVuC6Dg+
OTGhvhLyN8H8zTSevOnVI54ovHaiP9THf5xXo5/yz3d8Gb1IPhX2nIfBP9mYIp+0b+SdifYWKl2l
j2X2KIaH96S9u4LTXZGSS+Q6lVkl4gMhFXDvSwjA/+U/Zj3D4DoHgsmAZImoUFKSPCLbzM4K6Taj
yq9up3FTE6OLdoowxVMT6IqB891oqmruwwWNdSh5c8zLU26PqrYgcech5OrciwjrJ78HPWR/Qf7m
ZbAHlGk+F0iCReaiEwsS9EqvtTGwI43H0G3oXjIhMyiJboG4b2/jmdYw2uomY48hT8Y8yo9F+WmV
f29/EgS3UoUVX9B64JDLRKOFFF/zfpB8w6cSShFPKriIFelVqwKr/ivngCYPQlzJ0kVJAJ7t+d1J
BBl1I628tpvx169g4Bx04bT+5MYZIncDoIVLsFnY4r1fx5eCQlPh+3iEc8pxwKTfDJ4qHvqVrFQA
KgTUDegkFIZhflHOgcZjxrQHuuQckIhOYyQCHBHhN7JyRg8z2QFPkCUlUV3tjuyt+YrGCxXbaf6Q
0EMsA3X++QRR08lt8JwxE9xPdArniWkwqmuRiJHqy28pBXtgjKtYkWGpJXYSMp/tHnPu1n63B+5D
RhNoYPD8Tf2m0b4RPxaLiPBdny68yFgPJGTPsalhU9h3XMJIJTqn4WDr6dxPQKhWw1kFuk5woqU1
/aCH3na4fq5e8tRaqT1XbWDFFUjv05N/si03eUkN0gzj+1C4rp3X0ZCqvpwSse6ouENJD3kICAeG
3NoYAwR0/EPNXQRlmXsXhdpke+727PrZMsx5cDdUcujP+0sXjmIkF7zITvpaXuS+CBdgO/k2TLCj
TjDCOIGifcrUTuL5hIPlxSM5rklp+93F4yYeY7/BN5bLIzVABLZ/JRj+vxDX9Pf8TPA0wheueIQB
BcLs+WSo9PJIUvnh5WD01EtTakIkIJMrh9onGgGRCKXre5lJeRUt9fERILIq8dJpvwLuf327a+m0
hk0cLgHK3jxoRVAlyYaO/qTxfDQmaTApV74j0VMtZ2BYE10G0UC8Cf/14XxatALHtcHWDHW5rBrk
8z+keMGUAfebGtD9I0dajrS7LGSsEk/Vie0Y1HfPQNDxee+GDZ0pan62tt2ayV0Bt2vU2g6gB/py
9H2cQEGouQgZJXFPkOTgXJzjFOSPbqpuUEmr9eq1WK1x6UtX42KfU2ffMwrNqjtPhdz+2xAkv/+U
cysz6IX5T51C9jfQDeU6H1xsrYZcWBiDsNn59EHFkAVr5FG8e0nlGUd6silyaz5J4KupMbMrzCyb
zx3+VoB94vaoW2RIyYFwI2fSeYTob2zxv/jyRn+GQ7M0WRZjJm6rFjBUtKt3+QMHb7hSiLuvnqFg
7R/MZ7aT/jlvV6sBaV+LtqvDMm8hbAz7BIlUWXtp02k3VwVNlyabl3DxjKzOA/ITcn0Q4Zw1Z74z
ijFuAXVfTuyqxgbgmtNkAeRbU0TeQCSc01LNt5rnNdYAw2Gkhb4ScOIrgzXG/mlnINtbMXg13KXx
YSDczHjRMQ/zDPuCxENFh7Tg18e3yloJIYL/gChwi5QT/KvEmX26rvTKvY2kJ2whRUuP5Q9mTbR7
bcv76sKH74oNzuAfKirox/XPM6KvQDrO8OI65TpYfFrquzoqaYZhVayvab5qhMoTbQgwE0MlIT39
ConbUw6Hq4+wImUysdGEiCqc5gquB9t7Iivrv6HvvK8uVwU2dCScWXRND00gW/DBfwSIhiNz2t0h
Xuf+sH90VlurmgRAgs79DDd8+F/5diRa9NsaRIabM/ECxkSzQ8cmf7AxE45V3AW4pmTDvE8aKZpx
5qk/H4w66HbNSv0qcBLk+fD+JLMh7pukNYuPb3bo/vQ6/k1KMuE03iCSVidazM6Z4Gy9zfnHzhPN
geKklE0Y06of9NyJsjpzx7tmsv8HYLdsSbuUPM6EWu5xGC3b6mtQcY3loVWs8zC0s/LiRltrDPzZ
HTimjlGc2S/9OplQR4jUQxTteYybHrdB4ZUaYnYM4+FCXLjxXhF/Pia1aAbyAQEBAmlxT9khiHkE
8E8am8GaPomGn/TTp7uC0W4mZrcS2FDmRzwlajIj4JrlsbwpBfhfGXWRCAjiAdR08uuOExmgVIuZ
yyETeDnEv97WxV78px4VRdHftQ5evg6j0sS24MA1qgSeHqNksgPi2k55dy8bxjjEJnwqv8W+cEk7
Wt70xPTkI833W5cTwSktxK1pwVEGLjGhDr6bbkwPVDGqAKN5nfjVnuCW+iya9ZxjNIMEU7o8HSho
Dqhh2/V2OwFlIOkANg4e5040DT3wjJ3uGkmzJttBYnPg5o1TAxwUZ/Kb/zGUgdv74UJN+ZCtc1Gd
maL/4ZpBC+VdURcxLk02XSEyyyADhMhug41aVUb5x4sZO8n5LDwiuJaUYMhyMGd7Vb+0zi0s9RZf
iXUoLhxEsknmVRfP3EbLEn9ROOy0X70/t2znT2IzKnr/ewCVfRciFaTpjGdT6uw7guPCBrB4ITBO
JKFpEOjqdIlIM1kmh9oD77FGwmW+tMXM7oS/2TBP4DExusSTzHyAnPEEIohmunZsRh6LRt4TWeZF
hGNkvP7tLLZg19IdFCkkC9CPr4a0IJ8oyHG/xijHDNo1FomPjg+O1RWHCRXSDRlN4ZotRisSwmQO
QY54nwyQKL0x0cyJrHXzZGBOLeI83pFf8dgIgCxBGYeabXXKmejNiR0teQwBhidGYWPvCWH0rq9G
E5FiX310uyZi5/CK8ZIXJyzdfNfERGQG8Bk2W+y1xoW0jrVs/9VQ1zfF9C32H6g3ZVfEh5GWp3Cv
A30A7Bb8U7I+VMd4iBLqE/SEPMECJb80A3A2GusGLdF4pO+maXImNSEBi8Osw1fNOqY2zkh961vU
dNEAIdHcFMSNDm1qs5DpSpvqRlKaBuEEC58Sit+CFqr659HsPm/l/uy5UgsIMPyugVI3qDvg3A2Y
Sc47djyWDArMe7vWl5zWbl20aUwx7bJ3SDRyC5aErnDy/WsIFweuiyPhoeteQg6qABYrMcJDc2xB
bTVulOnMqVv99Xz/trrEsU+/4zDfmUo09TCjEyKj8M1uv5yIGgeWdr3iCWv0Jfm4/cK4T8b894kq
8qHx4HXD9M5Ixnnd3qJtHsPUyDvx/nkbKYcPpq131DGUIBV+zKCk4dkMOfjAJ4WQX5JqP+PoYFi/
GoFJSjldWDgKv6vwQbBgyW9g60vO2R7/U38q6pzux1tnV+31aY7Njmw+/7FYbv35Em/QZYUpjd1I
ksdTnE0EyZxkrGC9laeCGNwLv22ultbagbVxyW3Io8CwopvZx7LXZgQiBvDrJeq7D1dNm5lpt9Na
kDxYcipSiwx9OJ8DALkifeUgLdsjND6H1rv5Dz8Qd991+n7yWisgPSFJIXEiVacfkHUcpM3kIt6t
pFhRD5q7a2GiU91QN9zc5vsSSASwCViTp3Ap9dGrQZKtqj903S3huIbvnqhmFAdJTFzqEYfNez1Q
280cOGJxkSp7eifWYX1imHK3DZrac+29XpFLsSOFhKMDw55iL+/JDdfJZmdbvzdLpVvUcH2e/ayJ
6dDpU4QmYpH3Y/LEoulCJxbnnkTUyUc5k9RdC4pSSc1pPtywno9+H7zOs6RD8RMt5tOZVpBAMQ0I
zDxAtq27XCr4EykY8xhd0NsEWLqAQN4Zc9CHVLUQIkJ80UEORjDaz7kWCMQ8vxKQwF9zNduVWfhR
Qim/c8usubB/RlutzE04oWst4eFRPKXyJgkTddvTb/iauQueF23VsgPaP9dgw1HvU54XAVnUbK2t
xwiqEINpYxqsQoQnsap92jtw+av1jEi115bLcXAxtQdCfmP6qDEkSopf3Vx1YRHn8ewejuwphjPg
FROgrUD0XLtljWAd5O5f4OqTAdNFFXHT4t/wz7+E19+8gK2GpHFTOa//SMzvSG5KLf/rBDCoFTMY
vMdrKC0hrCKBsvmC/uNK7mFI9yihpzz85yFgVQErO+5B/Mui0S2OUDYVHk+zVvk3gpAY/cgypluv
grgvo+GbuIUDRsW4ux+eQbXhIwXSoF5vJSAe4KICo/SYbOs5zHz0kGguRVRPJMj0ily0ofkB04FO
nK8XzgJTn97XRcINEYKGOv8kUMgw9k2sxIpt9R2zxrNpT8XZT8bNCfji9k1C8g9R4CR+SGD8Stxq
h7ltChFJkiTFc2qsyYep7ZFJR7wKwAFBgFFSya/sV/Me2OI82mobjkNiRRqp6fbBJKqc8w0HiMc3
ISKtzesu+fVki46f8mQSCaf55e5p5izm3Rp1p1zBVBUGehnafSFLV00nE10vtI6B8+IVhsRCBSMI
kZlFOGSLIEN+Agtzspjy+DRdpD64nkgC0ht1hDvU1c3ES5Fc9sY1FRmMis0FWIwDlK5e7DJ5tW4S
KZPcH7tkpyn/BsJwi0uQmzGMKwi0FSDpLHnMzghCLcIzMaSehFcAQ6HgmHaouB1e46/IP8X0dWcA
IJ7MhxfSPlxshKZkjoNC7xVmL+ofOrUMvHWNtV3PM1AP/8CFc46wKF6RtUbVG2M5kxMADfKRF+wa
7RlBZ6lbV19lidg7s75WRoj+gT4FdLwD6H3FS+kB1FetkswyhZYWsH4oXiAAYBY5KIRzEDzMJbWL
+ghPKxz+6oQzCDEG+Ez6spHGOT43f6rrQQfuVe2Hy/QpFmmE1fAvfHCFPE4NAijbhp/VnxoRRfVQ
jtQ2pHQlmq638ROPaF40DI2mT6PkmW0WSB/eQxfQtnnpPpHuuqZgwZco7du26kHvHMKmc5UmXg4l
48B0Pzq3DkZlnTqHbMWuTBEGY4l+6VOWL8s8a0ACZSNqMCqhaIhc9yKUdkBFbuf/9ulx17Pq9Tyv
pUxbgQc9C/76EwkWsF5evMQjZo0Y0xTxVL8CS9jtoucaxHRz5FRDhji3x4UwqoBgOo0190Hd3OFo
DC/m46bVpXvGIMhl/aSE575IJuBPOhTrcci5zjaDHdfaQAP1a8WIVN/u07vagh8oRLyiT/OK5HWM
/ym2CuaQJFytMRjIJDdv+sW/2KqHcniwOrXBn74ocjlXzikSYKGUwJG45QQ1pw59OpmxQ5+/BzLr
NAz3HWIWm5+Rb0fGLbnkdbuIUGAHx5Mz+KL+z5tYtzkfhAImLXHSWDjarL6doTTFSA3acVKCYVTN
Dpvx2Qbe7pRGevcZ7CIwl4FPNb+bspCdTy3HGd+epzKeQciU+d0nCKDTZLhXMgN0SUNVBc+89nb+
Ro6plGAscOkclKjKhsKD6MI1pTzQUB49I4GNPZPR0HiP+KQhAfE692JvGgsUtiWNDvKLESNo3FXX
PeSRMDAXcu1xCvzs5KOfaNMgtjBeTfMiQis6ABeV1VmcQihut4duOlUN/xD6f3ZuJL5ouqxvmazX
93oU6HnDRmGbLn6+Y/1iRZoRfX5EsC73S7zdaz2LF1fyfELuDj5flGjSjUIz27VwT88CFAQyjK0e
t9TAUHYTLQsyDcwO3MsNLul3wn28ktd49Y4tc2z3Mca4rTQm4xJtqPfpWgO891crcuVhlZc+oApI
VZsIZtSlzEydg1TEKH0ESpBAKSJd0SO2aO7yFDNYyj2YL8C3ZfwLLlylgTkWpyfcqxPLYPq1O5qH
PtBqHncQkCCOAw8l4mFoB8JWoMCB/HivvX/k5h6j+OVAAVUziPeJ2VQFRIMhDHRM4ZiXexIQATgb
YXBoiblDBjqBSG+klNUexk0GVrhu3fQEbwVozu7ORHcOChnLNGvlVIFvuDqNZ1w3iMZR6CAVoAqv
0VkRwbN46xU9j/kjpbFOD1KqI2xi06uIt7AGfttxOo/kneC/tielqp/f3YNm3wy0SNNNZHSp+odp
fs9/QwavhvILF7coJcL5zH2yqGdPyJ2eBVH90jQ2Asyxah4JI2/ljoW3YF+hhN6kjCKh7PyOJl+H
PT2ht6aRt7u8Mp/eubPaQhSyBPdy7ZOpCbHKjcwaLNjnwJg4p3AZis/qJiuc31Kw1ddAjoJxRSgH
rPPTxjH78aM8by8+UlBEJSQiDYfZW9F6S2WqlBaZ7Ttd3eeBXmLvg/M3jzzlaZYSvRyTUXVsHKe4
sXdDfNzKVnvrpGbqtVsQtmHl8xgI4X/VumxHdY5rz2PZqBawmrrP7qtBsJHt2Ss//ySqqoc/upW9
CBnfTmsUXpbfiLYysIdlErY5b7Ft5jeSNweDshP5OCcBDl+Ckp9zJMZFPOub1Ri6IMZKk/ZIA1o7
dKd1gkfdmJHruwzPnFw+BgOo8TSIJFws4JI3qfVpCPTE4j+dew8xmlYFNE64W9obR6ws+kHndCxg
VNnBuxnYKSC1PBpyBdq3bzqXK55/qgGCjb4f1BEK+VIDUtnrMGiu8+2y8r/08J+glh1/y1lSLvNd
J35C5YC6u7sLvM+0P9nxeXqJgbn2xepsMO1ioijhRY+DhVIZ0RV2PnsZci1RLTHBY0L3i7IoWXkX
+8Hf/ty8P/Yn02N9FbSXJRk3ho485zTIreOyL1yVztNICZYdbl31qStCLNetTH9IQWl5mcbORtrB
g3h3UYVeCRoV7emoKfkmpGbjuPpUDmIU96uw6+eiZurIficOfiM40k+d1BeBactQ7ZixGSX3H3wd
n7FdgS9buzRRT7YMBl1dcvyPnWmys3lH6pGbK9FZyrFw3G5NVbK+gGXBkwPr5l3L3iC07NpuWrGS
s5hxWyYeVnPnBE+2HGKoAuxPv/Gl4+Ygf3qQyYgEKGAMoOBSwS9LpEbwbJOakhFBgVwIu1agGq1t
8KUpaM88dI17y99SoaZJwwz9rpSjUlELzTrwuxsWAnQY0uRA5296XfmnanP71ljJz86pJRURVaDW
WUKUpUEBM+xM8uwpEnkx4TygF4keXmsfw0FTkZSfJqyLoFgDgpYo9aYmeiAyUaCTLj/h/lvFzS/g
79I6N0DRlAK5/fsSi+2AL3puFIU4oQOmZ8udaLf8IjVapgHDhr3vMQ1HUEA3BTgW96+KxH6M/LIX
oupSCB4HRVJnBbusJ0cejlCYHCtnrp6qbjpPxkElJ3dsAw28ZiHhIRgicA6ijiuzVA3ArDYk6yQu
ER4e9QJdKFX9k7pfQaYs8WOPvo0/lg1m9c69AFb1GHpSgHy+r8nSTZAo+1LiId/kb2JfrAWR72V+
54vrOOxfXO1SCspZ8o29B9rulQesjl43rs9RBxh2u1Mx+r9suXv2JQ8kxza1Epy1IoRNffFKT88h
MvPwfK8PZSKpPRPa+cowvaaW1uWaZICOq9Hf9f/G2lhla97fRYYvWTTMu7aJhBht9TTtV5EeI4ZE
TtGy6c5qhIU/xCs9st+0H+38/lmPZRav7/snTVneWoLpb0o1FZXHxlIurVFEHQLDyHPrCJrWwEuW
ARCN0w1G8KKBMYMXHOevyeOamUB1PPnRDyypBvOZSTSa2h22OfGe24SOasXhe0W86R9kj/pcxSEz
44/ru3jfM4a8VETZzlHEwdCZgYuybiSwa4lsHHDM+YMRarFFlMbhU3Z1GYKYY4WIB3mFJpNeZ9iu
Jah5ZCIvfRKDNcn5hOA7/i8p9Csp36OxJCBOw0t5DvHXzE9OpWdAEft3sENfMsgPb21EPmHLiKcv
GAHr+gDErHS1vyML4ydlwiqFEfRnEvt6In6ZkIpuMjLdcE8jkQazytqkqGr9kl5kBho1wddpzsw0
r/CRoAnH2I4zrqOoUd76LeM79LqOMNN+IDX9AHyCREb7y+M9noruroTUxk9uNnADMtUdCWIY6kYy
RR+cILHUG7jtvzupyj8C9kEZtBjN9KRqOnTjDeyPWRdkfqKJgktN6P7tPz9O0oOR5gjru2F1AvNu
nJgUBUmhKrhnnQomF7TerVl/SDPiqIaOiwwH8r08i0Qf0F3+asLEEBWtTQCVu4c0zQL8LEuUAhTA
jjUyK13TbMp3x3RFaXSYxqZYUY+RrluVVqrdpHDIeCUZm5IZ2tjrycBX68rmotc4x+GUE/CktE2d
gOykVIMMHy12iHO9tfXLajpFKS9YPfN2Vb8ZUdXSc4jbJ9vYezRqYz4vCa9GOxIa7uPljnogHYfX
U3jwnKhFrijOvejsoD0ykGCWZuBtxRFpyFR5KAHzxGUHM/WXBuU6Jw4e9jce0ECVx3n15KtD/hVE
qK3PYHYsjXKbsHpqJBKGU3B67KNSGlsYMeId0bfx+XKkt+kMxIOZiKVbk1V4FTX6xIzlRis/ZMLc
RKJJ1gIJVqWdIf+JjaS2KmiQzhmQ5hMCFBcljoaBVhLDKs3k6z7JXfNbsAM6s6zFrcmzxdEFbqYD
R9M2BQELzHi1HXgVoE1gSCMkYmyy5bYmU7awgmKeFgCrWQ9c5gYWtOO/B5R/6fa0KC37+eFgonwV
pSSbnSPqeGDCi8hH6Mie4+oN6WrdvnYDXUdSSCs1b/MJvbTAFgvCWyAlPu18lJD6EMIGimubFUi3
ml9vai8qrqXdxSQ61ac7veK1U3h93UwDeRPulJAbACZ3OzG9f3Mktgcli+Z0FmfVd/u3J+LGFHDc
hiFJalbaFWC+r+KGqp5M+trdKtnp+07Y+RocxRgzMpvUGoThT943c7lrTdUMVEWGVS2IDRC+2JP+
HoTx865ayL07tjQLLdyV69StXXdMi6wfa1X476vXoooU3K1xE//IhhOEdJQGbVy39acGokhdPuBr
MpP+0n/bov78aVGTiOVmL9KzR5wufT33JyDicM5mXbuDCEGsxQ8sduTMxeDm6LbwethyLNLkmBTq
v5hncrrnJO8Qpwdz9gMoUtoDwFtf81bni3fp9XBQJOJRzof5xZFGU2dRw56nuGheL3uleXVBe+lN
/JB6cYD6U2D2mPHPkZByGgh/Yq46rMyBvlfq4RapbDnU1RnaeqeUqYU6Bc24TiD6x984Uf+g4XIn
RgSJ8UIUpqBxkwQZD5hsQO7/6DwD77YVcwS24qzidXXxRTBy1lfe+jUhfDpOhD3OoqMHNsilw6TA
zXLcMQK0CD30g4ALL/TnIfUxXA1TAb4qRscUDVpCVIOlMR5XT2A9w6StYmHhIrwuRxM1oCpOZIAE
F2qh98gWRDD58RZKZCvkzh1fuAgYFJoFrWwKCy+nL10GN/ocAN8fXQ4TstBZPCANmS8WFllWq+oc
93IwJ4aLA+eVO+LlMv20LA7bxLAR5Q8piPSmsR7kZoLshzimMg33DMP9NmSiMV6226W/IhCFteJ2
mpMcX3wnkIpSAgOSLwC5XodX0Nz+985LrDVR+mm9ywHS1hH/MDHcqSO9taKdDDYCOyW1mw6MFLWo
9Im0hoUruYcWRq2mBzg+dC1627LkIBxy2oy2uCF+yCKDoHUNbbpI0aWpVnz4pXa7Z/2qAmLOQnCS
kiNN51KXJ2ELh5Goy1ZRaydXF89uq2NVgrDm9GHGGrKgz2pl6w3tPaKIccRZ5iHcy8cOWnvHqZZT
uAv5ZLfcZ0oujnG6PAdtuLC/24hN+4SlmkrdwWpnVoA1BYhPzX+J/ApsD8JRzFeF/JpAPrLpqRWU
GV9e9H5tsjoV4VDkBgVMuuH3cC5wCPjsTPUidywWYXkCS/Mdk64WvTu7FyA4//BmufLfZJNPCNPm
RvoX+KpQizA634pqVOoozHV2OoL8/WbyJux6APGQEcow/qnZ8IylMpxRv85xryn4/kg8ptiR7pD0
FX0lnWvrZWerdLdK1MJHCVr0nQ+AAh97aqa1cKsLA0xa8RU6d4MzFshP9uuNu2q8HojMkrvLIq7+
4v/yvoV4Imq1ga9dyBV3qKqPZJ9Pkzbdt7xI5gDUiM+FaFfONLoKU++EDE+O4AZ8ivI8p7aVUYsn
l0RXdupcfB62chTxMFEP2NgqlHL4tDLTSqv13iq69vyqyB3U8pkpcubFF2oDdGX7Tbw28WwEHeu+
DwT9dxOeia3+hpp4Z3Mkm3BFwDqd9Zje+dqyfCDkwfJCMgGsi4OkNp8UalXp0CtSZf7s9X6D7qri
P+QD+vyVZ3D9m4USkpfkkNR1DJkbwNqLYD+pQgFkdc+PPhvJyzioG4Mw+jffoZRtnU2wP/FLJc7g
rYmi1YvVvyDWJpMFh5tPHqTG7SMTLTG9scC0M9EUZMxjRYWFSrt6rWhIm7UZPWqjPuZOqhGbjzAv
tDryHQd9h+fvTYgQOhluY5zYrweDcXarGY+skvi4rWQ//t5Ydwawim3t7+KRyt0HrdER+68KpOJX
G+JT+OK0aPrmmlpach63oV2K29HziGhBO3W0mpfebFFM9yU8YA9wZkxHt4RbYowLz4V8SlkjmDzR
cPDZCeQt8DIhdYwoSyfTY7Fyvz4Fn2VG82AhQNnkQreihu2vD40uIgI0u0yc4M0qdQ/uMMDmwfEN
Ty3udossHKTK3uBuAQpsXXvGKpjOe4VD3Z186NsoinRziSKW5IG9vCK8A2H3ebNZWQzyeEEbtX/I
+Dp4XMhPSs7guV1IF/F463Gdr3ojmLoqbgdaaMp+No8hm7Lmycgwu0Beqr3Mb715LPWEDp/R4pFi
xakHOuAwFSwtvVAEa/+sJt4ahnkUXstWuWaE1XDq7lJKZLEEtK5QABZvQEX7kggh1+2NYgre/zKf
O12ni2OFmFyNLEos2OcqlQTxka4+Hsmvs6sgOgP8pee792usWe3Zz5Z5+15wbaMajgLZHlVb6wu9
yxOW1+c5T+RZ1tvYManf572nDUh+sMXLmjkIkCEf58mYJ/4902iPDddH6R4cPvifzgKH3Uy1zLq0
WbeffgpdEJlFB+cUCMvIr080qnrlwVCRuRusiE/h9zJ+WvRYgpDs2nqNQtTzaxJQTa3LnusvYSqm
43tvy0YiTwCPaaxdehhBiTAysCaY98nEBlnQOJinzJQhlDmNnH+ytdEv7k23VL0733t9mslk6DfR
BdTM55QpWNX7GJM5ZxNfVxtnh3AseBRiY4vvMXplhFWi5BSx4Ziuc/HC7h2ei36kz0/9yp9yD8ok
nzXpZGmcUiOQ+W3S1g86pZn9nyuKW0K49D4TLqcjxsN6zwWcD5ihusDmVcGiGyBBhFr7txuEWkwC
5v4/xMXsW85vGudzLLU0XR/c5zEMhlZEUB/a6VFGvXAp389aKVbG4JpURvqrv0oGOhZxY0LOpLvN
gJAWqXKDV6mQwrHqRdSwqJy9YIzUoZfvJrw9eKr2iedpv/Wg5rq2GB4NQKOcrEsVwmJ6lYMQr06Y
3lqCFuNwyCOwQLv0+AoCY75Y0fdN4g1T7c2moVbr4ac8qU/fgpSNmAVnSHLNMUOyfglMcrzEkD90
Yz0HpZYBNRnFicrfm+/MicAizFdOml9JLjjJtNwqNvQDCWgOwkHl68ydXMcgCqekUtvOcuRXMvdT
305j28ZWBH6/idPcaJHJwM2xHCKSVwXVaFQTAO7W01H11ANTbFCTqiIvrnmGCMhFqe2/V7EzUTeS
wX00EMyf8mRlfxQBQhkTWCGSm2T9k552R/cBUQb1CjfrWOqjwSXsS/TIzWKz1+N4CryGgh8BcEw3
WC6eoZS7SookhxtYncDwAV4Qw0mptE7tuZk6tKDERGBYeF0ONBoaZK3oFEprY97s1gjHqRt/l77D
MgQWysvxpEjoLYUrSnv5+Af7FzieF5iA2Dtnl6yM+e9tiDXS6fQZA+y1ipCs4F181XKlRvYF0ZWh
kESgTf3rIiXlwIuAszYF8Ovxmf4eiw4Pyzqisvl3vgNM26/t7w2yTo2BJ5krwhT4h7Kp6Mq5AxsF
RYhbS08Dkq/cXav/Nay9i6DWYBXCBLunVjhpDiiYFRmXvvm7O+cg4Z3Rg5xk45Q8jAq6H6xE0uXI
Fu+GGaYNyF4VoGfq1aWbMf0K8lcXP/VnWV3acOf2qxKgJhxHL4uvl6T5XOZZimoNSGSmwGNIRrM3
XPh5eX0thf53wdZZyY/9g50mZUfsWOF4RFyKcyBfgsPcO/KyYzrXLakFRqd1JEP/fG+MJouAM8w7
RVl74Pc8NIT5TOLQqV8CWWotOSdseGjtx30i7jdsQQqDEfBrlh8zZDeTRApwgeMvYArXPfS3vbT1
PG47oAvERDbWzHZVNAAeYU3ycTLHaIW4ASObK4e9kPxpsT+xwd6jO0hGpzXvu1VCxSs3OldwGnEi
NcTmWuRXXYJtrsGc3INtamu3y6F8NGgtS/g9BmcXVmOLVTcZynMMLHs6x8mOMtIBxsKDIs6PYE+B
hMezne6pPy2uqSf1X2DYuLRBJ1Qo8nzuRfCyVBcABhk21w1pQdTR5IQdA+PPQmfNDmRtRjyItXbM
evIf1idOQpTjJwVOtmbZn4FZE8wyIXBl7GxsAfeRh+yEg12rvhv/6ugFQFWDwkO08UsDvNehhHom
iaLbj6plaKZFRJkMnkpbpEI4VsSqftdNsgN3MnniMybTiwiU7eCfGgGXdJWpX12eBr/R6VA/Bxxc
4TX66t8Anfg3l2UyuVWM94DJcMhYz6y2Q/onPNFaZ1rK7S1RrZ9kdb/tq2G1CvnEL4ejDX5aV1on
qaDgR2ysiEU/qM5xOAYXrHN6xiNcixYiVnTGa31D5NNdG2FtEUhtof+OWhlDyo7wfjXHx9rB4jtH
O5JgJD4fDYHh/XyMun4akknmjTzdfzkzosY70EL9gqZL7Od69FqQt6ttMVAxGRca8cXdDSvYGOlS
eM4tyffBvQZC8IvzUrYt7SMWwJ8aKbliTOPo1I4V6V+OxYxKxv/1wxk2O/H/LYJEz+M+A36piNeQ
iyZXgJQCBglOdmKO6FpY1xxhiThmhdsXHSTtFf+SF9nLji09Irm8wsfPGi5VTakqzgEf3u229cAy
BSt7DzbDxrQdAMCJwZzxZJZGrFDdOHuc2Es1ToK9f2od4KULQmj6CKkAKW/psEVpa7wcwrAL3Z70
+eYV42kh6xkMUN85xWDxJtlzk/ClbSRr+WvePsV4qi9DExjTEBLrGxK05za1VcSAhBpMmDO0eooS
34TJSM/0TJB1QR1ygI6EgBRzE4r1WUh83DHttt5X1sY6TjzjkbYzONO+dM/VaMy3oXIZqLCo5o00
nj1SUHP7X4JqHliIQEIfp1zhvGSNvFGpUi4H/aBUH0d3BFxtqZ7p5KJJgO9eegvhzi8GCsldmXfU
Y7eo9HsiyEoYMoGcO0RVCfwPQGqobKGyQES9ry7WXXkr7zRSP5/LVPT4Ae7e2fM+eHRHyN8GIv0A
ktexp6ZERO0eLDJDPwDbNmS+9DoDs7Hi555omSJtFCzkmihXKL0QJgTpXUVXUm1rL9Mhd+EQ+xLT
Xgqi1SHV7H2SLa7eXygatKufhTgAqITxrFJAJRKesXRfdXQcTyL081eZdChBbVdUZx+gOBvx9zjp
pZkGU7d1SPF2djfrhNiLMuRAP7y8HwofSlKXu5Ym7VBww5NBg+D2jBYP/AbogyzFnx30FAlaeupX
UZyeiA6h/Vd+GPuuMy8nASPa9qonvWMnXztwaCOg5bxOsA+uNRblRdFr5pkAYhYe96x1w+QoDB8H
aKk09o0pQ19bi18tvpKp8/rfO5jFbtdSpcQCm8fNxYBz03gysqt9H8Yfg6cpPODkhNiE81S1uQby
A4YllJm9LIjtocwUYpSwKt0CVNVNPKX9Ob+v9/xx6Ckyut12vw4X4LbqwtNZe9GXUu7Jra6ugIfn
KNLSdx9mza9KqHmSEH2309TYxLqHzaOEVkrIuvxTW0HRldvjcqXHRgJP7ePzJa/JCg6YfDEvY6MA
Ze87McA/CR/emO4SB+BwTw5yFVParhLjpSBODv/iOvTpkyKWWPPAJyl4DvirDIeUFxMykr6mx8cg
l2KslzGaolpRM6axKNZfvjJ8obYBanG4Oh7nW7HwlEwPsg+sFLjbzi3pov5dXBpjl1gNstYm9YfM
g8C/BVe21pqm/K/MoaiOxivVhsxK+Hy2ovTdewr9TEoqOKIaWisyNugF1FCcWn6uPTkaJldX+pFg
TLldcqsFjqDbwq8GLo9ij9cZfVGwIv66qWYf3jiLPLQVVQJIZM7OnC8RHRc8Hly6mEvie6YetMM0
oVGESik3VchYP8IRfMUSaHYxk3+AihyF38VyUnR7tgSAcdJ4Jrsp35LFsSh+PiBDukaE+RGxuw4I
n/xXu8GjWUUE65pXe4NxUiT5d05Imwuh48UBWDDx5+E86NP6ySmc5zTD/KlFxwqvEfH7hzehPLID
GNBwCZszNEP1lxcHzYexhcmdpnGEJ5zyQRm6x7UlR1uMfZK79+tFerh7djWRz0OeU7hy3Dln08Tq
ChB12x1xlcVVAhDdgbBQ3EpyqmOJAIKB7X+qW68pa2pHPAJT0O5sD/NI6nTlnCSH63elAYnScRYe
2XwDpFJ1ixfBR1KOPjGAgp/VQnjyGjj29FMLGKLf2aNYeYN0RTLUnQ1+65CasIUM/VoTvyVruu+f
FP+Vi5smO29Yd+korVGhKlfl7OjGE5LsRUxoA50WWLUPsiVmZz3maUB0nlDy3Z3jvhP02u0doDVI
EBQQ06GqmXOsW38=
`protect end_protected

