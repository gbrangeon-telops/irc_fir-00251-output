

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Hz4PNZqDQYlRQ+ken68CUlKtwl5bD3KVcGYwK7pLDyYBwi6Th9L/PQr7ts5tJoXAIQRYcIzRxOvE
bOvIjO60PA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
GP7r+Hw/Nq0CwA10fCvNkrkcgK45iHUPRmPqoCkPDKd3ozfduaGFS4NbQcQDFEPry0eRmQ2gSn3i
AGkmBiS/ZMkSitJxD/EIgYbO/fqPeNo/xyESKAW2O+T1ZwGwXyv6qMAp2gFqycRAbj6T5U/FUq52
EYpn3NB0sMc8yOEFyQo=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
le8HFUmlytAxiraEF0H5rT3qqsng3b8xZZHcvlli3mx0SdV7s39NBBuklCsi2z+U5UKSzgnk8WIo
w7XOgbkBH4I5bMmtC280eEWQOIcj1GSezKn8Kq725OUTUl7WIOM9hdaAEgsyYV4aegR9ufM3pfv5
jM49vFUeG7XEd7xqdKUxYcrZmsZ8CqQuOZKMv7+xnku0k9eaKv42hAQ7cL1uIXuIFvzDlZHyC8MD
e2+jTkJtzyJMk7U2Hncf7jaM/O2gSIFGoRR2sNNwVB0ATLYzGBnoP+wY1MWKJdSoIbDQ5r0792eb
YO5yRbe6PhUe2+UdG6sNzgiR0viGJQ6R/9i02A==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
tSJEOPsqlnARL2Dz0wpm4XWyg0nGSs+Wnp+fpstkJG7juRdPH6snLi4H3YFLGcOIteaUd6+0+nV0
HNDEDrgudSIwom4ffSyyotXElk+U/5goIr091+0B19LyBlVHPMfovruJJsH5yPOjkIUbE3z//OG/
9D90RTj2hDW4+5DRikw=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Y2U+pnaPqDjEYN9Ag4nM7UfxJ44UWPvMFi6W/IpytPtcFc+Gta7bvyNellM8zINHBtaT4/XvwpGs
zz9LduYm/i37u/eaLh4notjKL1KlEzSl/RQQCOAWEkJvBF59EPqbeUalx4NMTEi6gApYczcwU5ry
jjndsvqks3Obkc3R6uXlQHIzKbPFQM2kj8SV74srGUscAjTY98txOVHFhIk/okWPW2x7ScPBZlnH
/p6enNTFgNVy7YICPLQQ9SjExe9hKly0/QrbtcXPdI2+m7HVD28iWrn6JNqPDPmkYTv4lqGhGruw
jT2AigpLW8vV0cP+HITHbLQV7l7eN+9WNmGRNA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 126368)
`protect data_block
3Bbj6HkZmUN3IiHRMyjAHVtrS9GG7V7cToH/5dm407tuKH0FcKuf/1qmC830Yjq29WKhiQn8xJVO
ege8l05NV5HE9l1iGPqRfT7GuJVyyrbU2qde6ZVI4zQcFO9P97bJEXJ9H9rXmPOitiVpMs9vx6RU
Q3GYunlmlE30n3jwVy8HMts9nlBjb/9BlocmnwoDSCeynEz0mGQ30OHZGo2xy/YrFtACYOTrXfcl
zHlCel0GKEAETZqJL7khwLN9Yb9CmwQTiODOGF+Keaw53P89oNh21tuago/PkHhp5NdrrWhO6LcV
geWQpWTPMYk+j5v03srSS43iYoawEUYfuqZcsQl0lr2/iMXkh5FUdk+5SEKwS+49F0qYyHTpExWf
3PVew88Rft7H0PpFrKYyijpVOqMzarHvaUmkUItA5JlOLTdR89QjkH9cEcsI/JgcTBge7O3jAbyW
z2o0IM4O0oIThNAlTp3g4k/UQ0pRpPNMhzOzWor++DEJg9nexGhu24L3Sw7spQWwrHIZPLOft3Gd
qrAmpJ86St1/TTQSX0j31PqzIGkWyx+UH2QOUzfyuUVqng6HoNXbYJuUF2YkUbuv/sQo0by98iPB
J6zDiz6bmj8/ZIzVIj2wOz13qFYH2rpt2iVT/oDEFDfmkEnBN34QmkWWYKkDf+zbxH8C2hTxo8zi
2lQgvsP+yAdixozIYcKepeKtTRVpYzlMHNllfuyV+sSVJOHFisDx45+UOmZnZl7NTEkSc14OYH58
hjyt9UL2KF/lQk5bIyUWhJB8relV9JmpLhDPqIiOxKsX9BjcDxjNEuJ9e214cQJH6PVjOKzH7oW/
GXWxKQ0OrkIUCrqFi5ypMyixMc24uMKuv4HW6LIjBbQj95vafRu5E1WnNJ2Wdeoh80YwubTsWBjd
HsmxF2P8NzFXsKtendhusB9/+xOzhHVYZw2aAfuqyMQQsajmnUqOUXcTVj96f/roUG0UsIdJYSNW
WobIkECNIJ0e6WFdBC1H8mm38+NB5ukRj3jUNdG3yRyM289T3+Hq2Q1kvnN2hD6MtHS/HQ85wQt9
gLoI/s0iCXuUel7KKT0JUhGTKzQbjDKlR03iVjfn6CW+pLEbly9xQktN0yi/I3V6dQ2fVE2oB4Bg
JwlKHGFM7KhoKE45iINbVTBEXGfuXkqB7P+tGatZtoqZbLCUkjG6n3gHyKF6p6PzpqQvSx99P3pc
vtC3YlYeCszwpz6h8f6sh97STwnJGMrm547FdBiMaxZfJ6xOUh8Q79W0Ee7Qrr+Jh/1/Gn2OuQpM
jBlrig+X4gnSKCRGnJFB80NhuhA78SdyM399HkRBqkbU6R6t/CakWX7n3U4zlFv7Bt3KI4mi+PWh
X/FtdRCd5uwvz7XaqrLzIYI3W96Wt3laXjaHcjq5V9Eb3/I/MhDpN7NsGMDn1N1o7SBEBcoxxWBi
kuFDrAVF3/VzbHesocarbB7IWDabWzXXXtc5jxmTqIhkNbYi/0oXsV/uqYwtDtMlPcOIYepRZjPZ
Sxn5c5Js37B1R5Y7qnvI1N8zeT8iXqc4BS2RQjcn5gSNgweorJJMvf8pPvf/YOwUHLg3Mu4NZUGx
qxObdlZsWoHnlZjqNljL5fS2rzlIVCsLzQlZmIxc6Yuk4nRczFfOpRpaj1CPmIqXSNugqJSgLkX5
/8lLK1zKDW6SaHtQHhhL91SsWNDjHkzSWggwKCZE+HoRJ3QWR5FS6Y7bn774ceKoTF3A473UK+0G
tfvzScOasbJJMW6rnL5uZKxzpfKy7yqvvwlgK0g/i6gpZfP+DmH4eVuni7serT69rF9jV6IGI5bB
c2jWwL06nqO42goTWBPXUcg+fpTbY5SF2aaAU56FUutJ57MT51zH6dv3QzLwEvQ/FN5l/0WB3m8I
sk+sfngJRt3sssX6fWTMlWGI/Q4FQWOnTduGWmMglkuAt+EXfkLSpckmmP90quNGUqy7dUrpu1is
+Z1Y5a5NHWMJ6XRaF9H9mVdjvJFl0X3u7XDCtv0SiusPGoDINk7F+n65RYZUCCiPIKiyk7CXfQdQ
kSCimXKtpGwxMJlkPt3n5LdrXfIZJh2ZknRB8cpS1SsobdK6TysqtzTo3NUuDTjXBUpOnzlQrdjA
03sIruzWjoMp/zlynlg1dhs/VsX04K0JZRRcEBLBEhausYa+TUFYivR4U7+c3mBApGpgUVbElggS
udPsHVuz99waX0HX6v4yqXn0vYJdeCXdikRmjbzmnIUmQlYsvQkD+Lq9ZV4hc4DHbN/hhfMRh0HN
+E31mZKRUSMLnbkPR5IrLJLK/qQ+Hy2zaxMMQemQJHaRhlNMIOLMSDSUCid9ksl7/VRfsHcp/OOq
CnEOzMcD2dlk9BLZBGVyJTLRG24Equh5Iyc/sBJwZc1ZeDL2nghGWm5f27QxOnwqL/qUv0gEnejN
ikW9x8GjN7fXU0dnl6j3S5HuhoQsKUgFcLaWb5m7RT4wGDfx6EoxZasThZbtCHHOmc+MgcCr7PS9
wkQoI/hflvsUUeZlYF7X1885ee19RJNfwaQ6dyY5zXcV5L7Xe9mDXOgHPvo3r9DFAxwTyZjvfB/r
ltc748uNiHnrO9IwCoHPMKXpmU/8lJseTkbnj37dYWL8cOSbbefhEeqhNNmMqQ+r3vxtcqAzxLdy
3/ePZ4uEX+H+R0WQraWQbBSxi9H+mzyjEyyCWg+4JDYyU5lBZtHQ6x+MAqtcxpkNdvhHLaLjWl8G
/5dye0eMP10vZdI16n2cvPK9gvYhrPjuO+wcqV9/KfgCb9xNqVHnVLEiRJNKEPMED/kmzs+Zmwky
m+D9zLZ/jn7KpwL9hD/Unkz2pJuZunPqDpUInFJI+uHRSegGj9RH41sTJ1O87HDfq46WnRnSR/by
L2K4c1aTrC5FVBJzbLUsb9phovqW3MaXgK7VGmos08Kj21PA4WIa4qs3XcOEXRhWjVlN4jw1U2wj
w1ifAk6rhtGE7IzGrP0DQPUd3eKUH6Pewil2DH7YrbXcL/HRLDmZprhVpkZUA55Bu8rdGu7pZtLQ
pjUoo1PfKNMd5pP8vX2BS+IJln1jBS7V59uoWplQDoGw/tezteJa/IE8wEyRRY78/OH72krnUCOD
bP2N11H2+Edlvme3KHG5LdyVHmcSVpal0t89EivxqO//v2TdEN+E3g5jyki8DGOP63Y0PbZtMvrP
eWikUlUVEzUkLH4MtBZUcYr6bIMc5QqH7jq2KBBY05y/vZt/qXK4ICgzbnK1zQH1rlP0a73PdhQM
1U8aNZS181TCmnyAf7hGsDHKzd+5ufbPT2CCds+913KYBWtFHEBXJy1D29FI9DLXHzAJ/nUX+3T2
OyLqIeaudvVs4p1PpaYWsVGNzyNd/h6/Ze1/qttRvPQls+CszAg3WzWVrmsGGdWDqgsWLGwxx1ss
nLycNHiB3gvCGmGtmTZCK3XunvqAWwt3NNwnnoIZWUMPP5WggA/8xsjzDDdAnfIZLCgd15nefU9o
3EjJKkRo/TyBla9vl7bc7CbKmzqNuNngPEKs0X0aV5qJC3wnQVb7Iznk8czOztLDpmUJFeoq34kl
KrzTW7Dz0//H2eey09+H26l5gMgIj7Ld8BvrSDIt1c8qy7ojbnxvjghGGSd4SjR6JkS1rGMm57Wi
Sy/mu1tqxGaGxvsaLz1ZE6GtjnT9xG9drFGSVbxUoKQ7XgHfw7J5yIneneipN1+lo/wwTF3YKCBA
LU1aqr2o2PXLQNIs1J7/ZdHqZzletH8eFwiCsAkLsk1n7TEwq0M0RY4SUXVqzNVdouyPsyosdqv+
ucy8pZZ5agPq9+1uB7BmHWtD4tKMR6FS7/vVqqJh1ruHrYrMRWHNFLnyJvdNV54zqOi4MaOwr2xY
7AtJCa6WZUuJDaRgAj5PnTLgh7AlhSXJjoUGuWIF7f9dcGof75bRGhFFoPFvwHq7/YFiSF1HokAn
3VZCcpFqr2J76MsygNtLV5xDT5Ez3rKbKv1mccZ/+F/WGN7vLpVco5LtvpEa4QkBkf4qpvODU3YU
zPK8feOIL1Wyfu2kwjqfc9VNDTWQEVxQm9Uo4WJ4N4lyA12ttCKeujQium8p2hEVTltHRczbCdHQ
KLZpN9YNpTbxYM25TrrxCnw5zQHdj4o0suR6mKwa0judS3iiLsx/4k2m+Z4ldxX+/U2dC5ikcZmf
/0dS5N5gDumcEwWTBqLxNkd3ZTNFeF1nGGwyuaSa41WBWWHBzvXKo3HXycNM71sj/ujQeEZyNMfX
ujLBmkkZD/bikQ5iODo3THF9esT8iRkTFeS+2JII5FAgocVRUk92/tMXc+zIng/+0LsS62zinkTb
zXYksO8UybsM7W4e2ZHDovmQASVdtUDKfRhgISqxa1VYjIwp/iRd1Guh88BmU3z6PEHACsJo71s9
p02/74wAji5aCx3bT793CxLDkSY+7jVm02XNjeAn8OMGiXKJE2qWOdKgECuItS/sKBuA3HPPAyLK
G3k00w9E+LpUG89WO2TNEimgYqbNfsu3cjWp0rvfs72M6o0QewZ3/oToyChfV6iHLD24tLyExJ00
xJ/iNQ4KHOkQhT3Ao2xGmMFYnoidnixw6hncOCcWYOavIbsydTCDw06UyYiCW928DB8IBM+SiZ8C
ebbuPkOB8KsOrjRkgY5JVsbJwY1gZKNw9dMzc6jf0PbmrHeIiN7qvsRmHpGHYpPYlB+7heY8rWuK
hxw2YORPnig/gHqK6b+f6SlMfYlRUo0q+8SFZXkrywTFjRPUEXpKLsAO65HpsiP/eQ6w6pHxugB2
ujwIGRGByQV/vUKDnL1RKHsb7/nIb/pkTCX7nbOfFxxFSUkzbFmBa5JRqsZrXmdp/aA4HqMFcDdf
lOKK5mK6Dmh5OYFFXC1WjOiQB2mlLWz3hStRW5V+xxUSV701gd8CxS39he9/82IQDIzmvFutfGzZ
60XRD5zIhgz0F4j0kdGJrAQqY06K6VIdJ+L/eemisTn3Qji34MguaRV4H8tXSHl3YzNrq5Us3ekH
sE2rINLis4Lx951iJQ4XHap8Jg0eB9kHAOd6lR5I4Sx6ZajOpBO6IF55kkKnZafOEHY1fOW24KOg
MT+Vh/H8CbPoeN2xNLGJ12LCn1TAVSz4TgnCMcnpWQmkNhmDm8I4p1+FJ0oBkMhDObEFzHRq6BOG
DNpQI+WujIL/ZxxjLy+bNrfSZw42UO5egdTDTguPwYDzbHILnoJzLiIIMQnR3vgboh5XMtDU1z4+
EE/IXRg7S1G8zpYIg/3v1qmQcE//0aaxWBcmpm6TCotIHDSXbElkLecdJmLaRcq9F1dcPq1BN1g6
5Cx6J70VoU4ibCQLo/xQzMbDC1ZSox/JYzBSryt8rWd38YH6oLQzQ9ZWdApUZS07WB86s76hHac9
9zb9h9NB4f3NNtztcg124396J7xtpO1KyP+cFa4dnkZNmDgrrONJJGKFXmnUO4SRAiv5QdMsK2Dg
EFS/J/Xb6aiPaCwOa7vlIKHyqWpIfpufIVOf5PVZX+c5IZW8wESDWrNtvFdMypcWifrrJzCftRRS
ZV/FNt/xDkzfnOFgpzVqMI/v93kfi8LnZ19lG1EPiIDvOY6mBZcPwxKUGnb6owZUjBTPFv4kzUcP
k+Y4gWcWh4NQ1ORIDw2aZ9PmnIV4FPseeq/xTGLrJUWyn+XmoRMXB3pzHlqh+mxGr/28UUm2nYCV
EjbdP3Rvi9MPgbyrZXudUYf9MOiPpjVq9xrZGOgjNYS4Dq9t+OSBGKkcuHVeUzkSpJlQmPq/7uaP
SZxx7hsCr7IEp3Mq4HgD+yWLzcM50xodV1Qb8fKUS8TvC3ZxghJQ+TwfSU/+W1IRuLAQdiGhfpU2
Ovl3pFCEgwKgOiQACiq8X5e+FKjEq0w9wgyndwSoI2lPVPlShVAlv5KN4CrExkMTSE0q9zxUQ1AJ
jihk679O0kp3dE0oHwXcNdWnOG0+vlbwjqws245bSPNbq5K69c/tlvses+7D27h4AMois1Ekokfl
GgBpKPpXhaSWdrM20A/0G29olBr5MXBYpt/El+hr91SUam+9K3rHwZcGYRMveJMPqkgnEfNVywOM
xuvtR772zH8CpSE7Ps8zfJ8e3sNn3E5HIqdVvyZlDEL1+Ox8c5pWHcZON8+j/dcpjj9G+5fO1g87
cMygqW0gFXctQYbdgC6kvp37WviGkUtQk/Fr0EAd1fNfEgnnA1YG2xRZZUK45ERUeRw8zQ+7lD9A
wk3b6IaNjEhyi20pIwvuFL8wf8s8k6zJk4Sg2dz8EMFvxOTVv4RM4uxxf9JclWXSnY/mZcAfL/Rl
vzTyZ1nJsrUV6Ixsv8E83GspYZm13492wHPmcpfos4AVBI8bpxwY/kbYKgxzy1pfheQn/yZsN1Jm
TjzB6h9P4qGbdt3DouABtQF3vdpLU7mu1VsTJ6ORWRksZF0h7dzPCAuUu908TuJwKLGs0Zh96yWi
KQ9Cat4oNtq6ICDEVIFPzm8FR1zcQchLliD4jFI1PnPryjuJInVsJM+ramxgs7M6LjLyUQm/tbIe
2jXl6nn6Fpb0H/svaIvvOtXupY0rBBKIOO73kHRh6nlmcIAgjuBhbe8vrYUuZquU8bCSm2wWCvOX
3+sqodGmSnzwi4DakyvaTvnzXTQ0mmkFh6mDazLzzk+o8DfFWnP2HtqP8UGBgTUZsGz5bEaK/Cs3
4n69myS7VCrHKmTbTEugYvOKqAYzD5CcZwt9wi3F+r41n2LjuK4o3xFLMgLkkQKlCBfuaiw8pKSj
7sSX4NPlNt6YINct75gbvPIWaASTQc5wu117kNWZBbFQMDjne633kKNK1S0z5kvRc8f6TZBx/FQK
y8r79rGnJYpnYf01aH1aSZgst0Mcfu3VtoPVSab5prwHGv5MN1W+7ngSLit3GDQGCSTpaYojDfVD
5G41tG5WIed6SSPm3PWDhkngLmzr1uchFE1mcUfrVHRFwZ0N17CimEcliLizL76QpfKxrX+7uOgz
n8tK1MlMf8ijAZKxeGiSr6X6dRUcxEb50s8RaVF6ChiokXvHUGIkl2gcCrngalUEY2mSzAHlJpoM
W8VhUFh85epvXTlz3RkAls7lO5FN6kT4F/pYRCxOSzyq3WDk618QG+sIh9yPBqK9Saj5aEZWKJlf
T+NsNMmN9xHTGwPxaCCooY+XZyPLmk+SvBOSclazpadAtYeebJXoWnFIHe9V4fZx1nxlWVQqhWuj
+k9qm4c2Fa0kgdeXNPZKaS+U3DiX6G4s3v5SXvyjT5DZLWpDatvP+uW+MstC3IlB9j+0IbBZO2o+
p7AxtITCrIbbk8lpOcN7EM7/kpmL6/qbiNRwqhPcbaDO71QAB84VN8niG1xQmgzR9TK5+K0nCO4D
/alEbxjcHIR1+Uk76S85vnfqHRvBU9j5WaEXThvEokCrFAr9tUA4/xYusX7HQxb632UFD87GL9XM
QoMN9xD32gpMMHjUYVxehk6kXs71vTKXkxTxNKbv6AgRdT2PANGmiIFuMt0SI+1eyEJ/Y79eoSrj
8KeWseD2h96JuvW99wNO3t0bWQvGz/TP70SOsWzeTgeaUhltWvtX9GB9zpwjvDVt3JtlYgm74lAV
0msXSOxrpJLOaCPMkhET02hn7dje4Q9WcnaZ2KwoDGXanw9h48IwQNuN2uFHoKmywTlkkBq4HMBx
yyLlislmUGvIo8OJdWkJWustKAFbCDRcup/qdvG991MKCxNFNkrP4s5rwkH+WXReLOaloBZEZ0gM
aEG9L9xzQ7hhLXmH39SzOwmGIPGa8t0gtNF8rPz0UFpuEf4t8pPwep1YB3tdu6ylgK871esbcg5R
xpRX2O+J0JNcWf3jFQAGNJboGr2UWIS1dIAYrUTI5yNeQOMQfat1dEAAY3v2ctp6s57to+7Mg8To
f/DmJeKzQaaFocyrFspdGX5TLIHCOn3oJor4YsGu/z5DkmFdZmDPhQxJBTYec314DzvGRpZskOY4
ClBmo3iTowcKvZz0iPeDPOY4RWuDFP15MJ3kNrb+c3d7z2eelYEkkUTT88f3mi3IMBJ1ZqzK1V7G
cmFpe4+KQ7Pbrb4un/oZkvUyeyQa3oplSVmVCZzuwHUftwFFMp1EDtdnEC5yNMCAl437O5F7bHRv
vv5K/meMEXG/PN4x6uztiOVogqxfZUBk30KerCeOLGOUe26EP1JiWg77e6bYIGvj1pF7dfVXKh8f
eaOW4EILeWugmY58LCWaR7LWClDMU6U3pNrs93dmlMHDNoQRcJDdd/84EJP6qs23/1OPz8Pkp0wu
hY4ZG4CLxgvgS6q8kfKjIG4zi9bt+MlgZWKYrFBHQ605sl4l5XkdI8G2sUwKFsr9Cr9iqcUp+4a/
ZCRMGZHQRfREYalomfZMs4oU8AMGyuuzelEWPEJZKPLtHdwhzsGYPrLgPCKzdZZo7uEY9B3a5Bbv
2ezu8F+PXZ4LZW5zwSPbrbfGkPLU3oJBYEjPu/GInnYZ8yEaMufINbshtMum7o60fK2xeHbfm++5
MeHJg3gFHZbH0d5NtOLyP6O7rYwxwg+KDDtoKt61fOWO1SUFfEtMHH5En/2yfyR36vFNAl+6ja9m
JzyoS42hzbpXXFOOojP4MFM01ZH4bkiJk3D1pBW8lFq6kHsGOpeLwgpUlLANrNKiPa2ZLyspZoNI
mCRVbl6KHxq/Rbj0PbzWanIJ6i8gw2djfck44g0AsP5oji0khb8q2/YCK5Cz6oviDyekJXBqUbpV
GJ0LheSRl/n3Iq3kAODqR+mDjazPwBP47py/2u+vlXIB8YhDGLWQgkvgesoAzT5VYR7DObUEYSD5
Ko5tYnQshPabKBduWZxMziwor2i4QUUWsjlXxfZ1zamJlsYLKF2bbeZsxTH+Vb9OhEtaU3kr0tpN
v/6zY5t7BWthIZ+ECVjQbQWZHAQGjy7bPh08SSMYiPV4D9fpOKwRi0r/U39+OEA6OfE+57XbZmAp
bRathHnt+ppJtslYO0WfwD0NmvM87wjbewmvV4tE5C2ilfDVMquNw0aIzfO0LH6vY8iAl4tZLwXJ
lD9Rds0+wkzLV170Me4TpKwNh4nr9iUUiJ3w06YX6EhrHS66YVoQkz24PLwPz30Cng99qDWfkvd+
zP5Gv/NG/IG6zNzUYUdPAQb56Va4qW37MhcGs2ABG8yfqDZafeXHkVnniK4k7B5vL9283tNYEm62
QLtTcdjmrnnGAPJ5+cAygA66jyCVXM6HJMvnx6W28HhCipbBq4tRuwp23nkh/c+Rbu4qm18/J84H
ddNhC4ZNdm4H33KPg+WrsgQqLVGRWqWg9TBzqu0gSMDD9CRLrFOBEbYU84pmnReDdbp9IRFXBK+1
eIwk2z6xtM8Vv6Ff9p/tcPKEEW3k1kbaPFzQJQTmySgmnd9ReZ45NKXzlpezGXhr1SIs1dPEqg/d
rOwLVwCtnDUivHmZoDijpCCIVfk+1n35eyigVTXwDgNgJ9pUMQhFZO9/02NpCgy57nCQF6xmLOHy
nocwDamiFIqIjrWchLDpMKy3AQM8C2GupxF2lIv71d3DuHVNL8sc+hNmer/Phvnylze0LIHOdKKV
6p6xl/2cuUviOc0g541FP1QVCWWUk/zXKKYTYCePytw9yrGDv5exZhGKkYt9IBGksTlMv8pWZYU0
C5b2V/4SzGiEqIHV3PCnKXrWj65axp7tiiRbZK/wgkGIsBH2BuCUg6XfNCoB7WuuHriYA/wMywrM
1AMiA/bUM5elqr0RIU5jiL/NFnbniqCsKdOocsG/d6X4pXPgkOAjSZpVQYS8nJRrTZT3nMd226iV
6Pl7hoLQjluwTv1KZW0yRCTjvGLg8mORHj/sI2KDa0HqrOvIttrrbH5Q6EpR4dt6qSJsgOirD4I0
8pnpw39MGlIyz+bFDMMC5Wn9Mm8GRwlKexmE0nZsmZz+kictLrNWbI0FwCN3pmFjP9NJv1ukVGt4
HOenqfm2TYsa61RXRCRbX0ukmBpbfllygSaz5zFLvlElJhs5CFowg6OzNUbAJ8DWASE5T6rjuSOC
PzY7Ih1Khct6edERTLiX9gi6cUq7pk/xrhteAb21CQ85MRL/eOhhDJ02tdyJFUCZ02VUZkd/EIPu
uPLf11vjh91jDZ/llmca2fi18o3senHGsJJixIJprtax7BoHDoJ0ppHsxO9PxKno+TmbLt0X5XUv
ny0S6DIC8LW+BMKTm5JDiQh+koKdwMVVUnN9SMsHF4HQRLFPBFX1LbwlzI03p/12LZ0cqkwEBQXB
mGLrxn8BjPdkqsUq7kh2nR4VkyREvbxNluFrmZBqDGPnrvx6OXIpwdUTaKXCAuHeWOZtQT0yJumj
qNuB4OQXXWji1nbdfOV39KEVwBKeH+R6JdiIfM8Dn2QtAIFawnR9f89VPWXpRpkxoKNYOCd+IrpZ
OaH8FaFBhQZT104VzrB797445JZNtXF61M0mxCKgy8/rAKLhKhE6luysBSeuMY0YW2yxnnlSmIYT
ri2USoyxqq7jWm+cmdCEIngRzfJd8XwrnhowgLjT982rB8GBsDeAJnTsi5+6Q3HBgHuI0jxAH9M8
U438cnNnjcl/zpp/VAkcgkIK+aZtVhY4NXRPt2YBfRs9iYck8KESjgeh1aM418f7t2jvbvJp6MAm
99XWdKR/zyyeSj4OtAM9iNBj9co4YJHAJGwc/+0iAm1SE3zzYWNe4Jv1Ha8jpezTq8hpzQ4b2dVH
RTUk3DQaHsPfWzJkq218tx1tr80rSqYjzOWPpR263th2jw4K3UF4jPnVIdTqboXDtT2xiXviRiai
QUdmLRs/OXPsNQjkRngfHA1wJDsGpUyghc88a4l0X9kbpshppoehkGrQ33cKE0dEtru1dYlrk/Uk
KrKz/tHCOd2Qop/iWExfGi5HQQPPmlrSb4COwJmvxEB7n0NELW41GuF5aJRquWiyVxUpnzhDwfTQ
KMJNqyXAVX7X9HH/UhKZH3Qht8dSW/gwpfeMsO4s6xgJ4vP76DjhKtJhRG8GVnTvt2sScbiLmMcz
DJQ+ZIdty/6YHEHhr8zRtHAjkMw5n3nXaIXf0dWtAFJjudH0C5PANNbUPsCwvCOZ5SltM9Ok16jB
f2koyhb/oU0OsxfaBkFApjMMB+1EZxxN3qbRtn6Gz4VP3Cs/z3Vq9e0GYBi21GHdZ8I4rNjFDJYD
HZsnQJ5x4EXii2Hv+ZOSs4Ai1P+r6esow0UMI3YxrLGlwksCtNK16cZS1dGTVN7On/QeFvAgRW0S
TCN0P8eX/duYUS6J/JwshtPasvzgPUlHA7g1eu5WKtbJQ+OttDt2ayb5DUKxT+FDzZJmftwPJ8S8
tZnJfPjI40cQm0nxcbbKE4IdAanB9690XlLWOJ52WaVvXfk9j5wMc3V8ePbuiAEjddqgTUIbhTTs
ZapmeFyA1sj5YP7c4xe2kj2ykCOWH6wR9eRBnxub5RJ1Jr8FyMvd1n4+fFRQs7qLjlmzrhpOi/vY
el2rV6rYc77cRiSEY/rkkGOC8qoK7jgPrkeXolO4P0l/zXvc+3v7y3Fmxm+ihs8/N7cKtjwh9NI+
z2m9BjWuiL34TAdgx8QMZWLNMGN7fkpTd3oUbHJ7N7fmQ4/J8iwNSafZJf/J+w0yhTUVLbm1g/th
f+IoKzFMu00xNtRTvZ/JIiVguCIi9jo8+HSd+e3mtO3hNaNU6foXpuWIf/kooingmHj9bEJV56tf
PbXrb4iuWG6msyk7h0wL7v0+5kO0KiUTKruAebsCq1W/t2q1DWy1nkBVrJoUUMqb6j6P4rFA7V3u
TLYXVv/P/QW7uuEdzvXhHvmq9WwURSrWRBvF9M/V4Flx9TUwXFLwJMmiTq6IFinhhhvSQUnaT4B9
OLCiublnFqeG973JGByBYgqaGbXraW3HO9GgemRkw89B1UClT/WU29EqTAAKMHwxomY2jPNcqIUz
AN31cMQ3mXM6nK3UsKmpWedPxraEnaAfo87dnI/Wq9OgRMMcHfiCx2K3N1BP6hLn8LXrriXc7MJh
tOfCBhiljHbEGxge4hFdqc3NZV0tiZeGFuAft6F4HWvsWoZBmlvW7L2pCqXWRi+QYm9cWkcYwK49
8l8DOQjUvTEmJYcdjbTbmhcswU0nE8aIIkNgZqD0SuaJFsaoMTqsiHsgg1hSf6upZ+aZB2QqxHll
cZj7Q4HFcoWrY8ttfssaKSwe5nfky0jMpLFyZG6oG+e9Vf7GF8qHLBOcrUBpOiUCDXx7Bm+2IlDP
j7Zu+blAryzm6hZmsMx+31FcFcoTTyrvY8jHRvpvNVQbrctUPmP3a7/F9sxLT9DbT6J6dCCPN5uu
k+NtVdGkOnnJ03r1q5zd+GA66llta90ZGf/HmGA1ZOM8XRyrYgvZ9hjqtBCLpw6vgIb2nK8gx7xn
rMkr5Sl9nPa/Xitn36h/n2AgyV66cZfZt6d9W2kyKLTR7f6VOsznebtiFiY9AdH6oQfjmWqkPNO/
3znFGALBJKl4S88KksHkbK5H2wJoyqIOkkRPgUURUUz4FrPVhAxi8Yi+55TbloB/PnL3bUqe8oNm
Xmf3DR4QOPatr+VUp1JqkKjKjDiEfNH2j2sDI04aKZrck1kaeVUYs/P5rJ7u5JXiEMBZVRfnu/Pd
yL9YRIsNEf8qPYgGkBOMcV67FAroN7UKoL6Ni2r33N8Noq3d48w6uYGo3rsLolLEqQLDygYhPIMB
0gKPddcOPl/qk8NZ+dlSaarkJplZ90Yz9E+u6XkJV8cUf5Q3fhUsc1n8tn90vZQIAuvrWwhkw2Xb
kdH/QGkny39OAl1GhzOjga/VtSxlVYUHseMiOVw/V1IQy4sbXuu3Bp/VnIV6TNMnI4rt/5UFjjBI
4R2ZFUNlcPYGIxTuXKl35igaC2jPXPhIkLgQkIZpEj3YDPyP19wgVDfK4OEN003bfAinW8YqqTAV
Tczi/AGo+8k0rg8H+IcU0+1Ej06XA3R7M5ODGlfx5+DY3hrZioPu7yl3scwqgXXV8jMsVm5o+aZv
yIAPf42VZ3hUOvkWMRWIYPJNhP7nE0zlsv66Hx356HQdgWJ/u5TjWDrucQoU9DEn0HhnMm2wm+mH
t6SFOkeSWqM7RbaJp83zZl5yFC5ckSYoOJ5TvqRUpyH+ae40H5kDb3wVvYq4M/hrgHghMBWs94YA
08ahIcCdJFR36jx5eC4C6WBlIGHrNFmbZIBhbZkfVeoU+QZ7wzPQr7IkR9y3ZO5NoJWZBaHe/l4Z
ogpaQqe7966B770YhpdwnP9Cio8d0kvOx9T+jEj6qXimzyvBAzi9bXDJWd9aK6JjGyBqJfKvSe9u
u8rInbjyPdllvUQ7lB7C2PWnUs244q7kQvC0B2GPGCgZnic4sucBEUDJhtc8dA7X4pVj2a35AMdq
ZupRm6tkwe7xjcKwvdc0LbA701o6J1GLy7DsOcrNTz3wwa6iK2NOgwXoZSPuYFo6GYlHn0HxAI5Z
0XGvGAPkrZvJPR06eHFYNV1ur15WEw8YHubWQ/Mqz4Vdm5YIpvBORUWBcFAf+TdW/b3O5TlPp4Hf
EK0bdQb/PQ4CnKFWAunSbE/7ude0ocP7gfxzoDGJwQ0L5ohhxc52ByirbpZ2ipkoQG+/C2s05Q/Y
aGKT/mxCk6WM6KSNUryfPEztpzzWKE6kzP6ydCzjDdlCtK+zGGNTo7aNzgW5TzJHDXimNRFJZVwg
RTbFHYzZ05Z2z4Ogz5bK3yeHJLqfLe5vscswOngz7jMsunYVUQbfdkbU/RlLYQN9WTyB7gy/FvpL
yZW6iZOvcvQWCgt0ARtRC7pFQ7oES3brIu4VFryJ6ZK4xIg920taiG9EPimjvG93wkM5dbbEXZPa
YpIgbzjz/HpsnJ7yYjn+36BTjgu4DsHCVS60vwAQmRuYyLeuLYZcrQvHnCVtQ1Ih6CYnWvWqNDCs
/4abbq+Dj00kLI/pqDVfojov+cHN69w+ZDkyRjxJSEpheBNv5TX8HmyfB1i4Gk0br6jrRavRzjm3
hTdq6D2QLaujOSYcT8yObVGm794ze9D3HIzmM578ju8qOZe9vVcDgbDWVdAeom6HAlH2GsEywv12
XwiLA94/0Cp2zQqzueXmD9g96LZWOjqZkf00mR3FMbh7P6pXH+M5+jlaPvCvj/ni9nwbHqw6omRl
fKpCtZMwrw3KRN47bTw69N+oXneb6rkpNyw3dFwGT0wMzDzzcgXyen/kyD6Dyuhxrsj+sd9GG4+R
iOaB1ZomEWHhffZE+Iwstz6+Bp2wUkByOq95a6lDxFVC3mcjP/hQ54MlO6Y1HmHcLG7bWRlFo3zQ
cYV5R35lhkZ6KrC1b7s2kxLTmMttBpFbBqt86PfdHG37VkWYDhBQgim6WeKmpANvoH23/7YkeXbN
KpYdTQfuC97cBv62U/LYp+E2QXKW4qTT6Zas+geXc/WMyBrOKon/AmIQ1Ewx8Ef2gX5tBpYbSpEX
oxhnNQxDelhsYcz8GbKUfxWjbE0cu386+vUfrxPpz48KcjmyYF0doEegrcY0mPj9sVEidQHmFplM
d+kGNdB+6LJ5RMCSdLQBbYfc+Ipbzs5/nTGeITqnwIzsZg8WUuCb45xstSxb0+VQd5XXREdo8myI
zhQ6XU0QHezY27QhS8U4OZlTllTMXSZRZQjEQR2oD6Wj8JvabLewirnjj5tCdH5WZMI/3P1UHbVI
ILwHUiQaWwtkjjs1RB5rRJSMEBuDdjh8y79NgX3EzylCKfC7sC0d+c3wBVWZglj2gww5KoGaurVz
2fgpwTQZWeF0o2PnhihG7yaRzmTs8KJoK1ExaAlmYnM9QOC09wOhs4FJQBGNTRrCKv3KSAFo/iq9
TjV8pC/F/Y85XOj/6ZjaLzxblLQuLFZGEoTf9m2Zfd4mAj41Vq9W6Fc+0lJTg9bcq3rQJlxfiIfs
cJnDhBFFtMbtbulYwH+oA3eq1j2dWwNOXv3KMxdmR+bhkQAf7NoW8FBte2FexDdsB5CTXJm3Wn9h
WMITMZLFt38dZKwaD6TlqioZww9C7F8mGU00/ZA4RXgVTt2OT7FwD2FHS7TLUjmtUOC/OpsB/GQK
65uQAZFZE8Zz/P4O+NM3VjrLJ9f378ijac++Qogapa5YEISfeYzDzN3ZjNhiHkThZE7J0NBg+vsr
YsCIK/Eb04yiDME7BAaFyNaCWVkDjtoit6qhKuzFa0u7B57GMeV6w7m3vDhg2Cs1c41UddoTjcV5
XkqcQ+SVHkn8xQcn5K4hTBD4fl0SHspqow7CmafCvRepi1MF+jad/5ooSPbn4uokUgN8AwVr6Yc1
tvDH2RasPWuCc5ZKagsAQjCz2A15VOuz+PLamSfkwCWYa2PQhVi9hTFp4d2f8VKwQFOoaUes974J
ZMSdcIqn5KJ/Q+VTsMD1biNN13K/75+AY0NfTNkW7uezLtsa5wdDHK7ixuUDA6DI4h2ct4jITlV+
NK96ip3ZIrlJ7A1+w0FC69RDvSeKMn/ofXGV0SKX0d3HKFjYUnyoS6iREUNvGRef90Q0X4zjYiOr
C7y+15WGoe0s7UvwZ/XDDLixlwJU667lvKAfEFo4VPaQJWt6qeXmJJJWHQQ6DrB6SIqSPNzO/qFu
bU3sRqi4R4eINwAeaYm7iKLkQBhNqYRhRUW+dyqIhVY/zK9JvYctdOcydac7yeGKaOXgmTz6LQ/y
u7XcZqrx9jCE9K6nDGWFm72pnBcibYZ1eMtlrTaYzlXjlrJbdpDSF3VR5ypet/KXMlqHDQ2sHMZo
QmTey8UlmltIkO81pb5OcLjUB+xumlmr+aOlLudER3EBFr3LNHcr4h+ws8DUsAoWoRHMPO7DXjuy
0BOIThuExXTCSdCzWsQ3Cpq7TP8fqxdYq6ehF/6E8WgQimdwzIhNDKMgSpTeAEfK9E5rmqKv8P37
lq8NJS5wJYucLmoyRQSfZMsE7m5XkFmrZHvdNkjowwHzQEC5+b0gGMd7h9v//0hS1xhvG2WOtT88
X2bergIRejhCvQ1Y4zfyQkRBaTSC0XgTr0qOUSbb0lmot7a8/I0zVGR78EXk8CGj8n6xUmt0hZgw
FaoRqoqY7Tfor2y7BVwGP64lFlaZtpNszX8jkx/ebnq5xLJJ/dj6E+5jt37cpPVYNL2WQGfkk1Ob
XfXEEafd2Tu4ZdP86yaw/3HHWXD4HhDK29TuW5a5D855sjsm9zDSK1JXFujwYEpD5LqTZnO1wUNK
L9BXeYSGXe8J1rFm36/FXSCQGNclBZB67/2acWB5mGdLDCTlwfUva7fL2zNGzbO29ZvaCGvs57rz
PfBtqcVUHBbdQQLZ096GMxH31ONFG6THG7dA9vK3I0kC4IOInQ+1K6AdLXBt4ZscAJ2uLPPN0HDP
MN7Et+Dms77O31RNiDYgkFVQWZs7uxiKsnRbpcXmK8vdZpPlskXyZ304xofAVFUEZt0LNykwXoxC
JmCaCqeIHgcPgfGeFBQc8M8ikvmjGdyW6Y3cocN/ohGYG5HGrE8wdeI3SuOfD2+n9l1PALHSH35n
cf/sy7CTb8/Szlp4j/9IlkxOcfMj+hbLnDCsbBJN7tL9b7PMmSeKE6GXbp2mnX97QVDzccTy49wY
HotyFKx8sv6pbZREHAgQe2nGi7L6gMW2hjF9AonvfgOXBLhbu6HCZf4clNWN6zVlkUoZji+mCe3s
4uJ28MWAD13EizxQmkAcOaBlGarvi6aMlBUtmTHQjxqUjSJdvxff+M7qKc8NpcsBT5juoiMIDEqU
AxIAEe4s13yrzEBGVnF/EiT+kiy00iaM2ql1fV44Y/CF7Zs4owyB36X42gQIqt0El1Ez1SI1VYKP
Z+QIaDyJL7lRSXQZ8+RIxZpmmknxt7XUCjEBWVf+33Y8fxMDXw1PCkfMsZfs2nJRVJpqbcC07Iso
Z8LaCyjVgu/a+Go6mq64WwVXLnibasv7O+aRdGDyiY6UDJgKHLQZTEZV0xUlnFgxpPggqoT9NI1R
wGPIh+0neIrC+BLcQ78McIVUqFZkFg5ysUVOOfk0qUEOcsGuSQ6nBVqTKxeWUEYXZQSYypn24V9Z
vQZO3nXQGDNKhi+HDSE3KGIWLx390vYYgs8khnd92u7NFPJ8Kwn1inDGR8InmI03MTxT5zX0xHpj
VlCtJ9jma7/DpovLj0wz5LKsBsrdRijSq1MsjxTXj3qZR6Rp28WJg7ft7U8liOGSBmclCJrKa6xg
sICrbA7SNdjOqNFLzWiPvWfNxA4Y00SBVUG4F8jsEJfciDvR7dSq3qeqQ6t5gPUNU8c0aEg2taF8
E5qyEU7Uvcmefmif8IICyZ3v26Q9dpkMxv4R7QhiBhRCbw9yF85eTNcF02gsOolErt3IJ898WDzV
wzzkoT76QC1qW16rgxCNnjGhUgpgyMeODPlrzNIDc1DtDP8GRCyyM3sF4U7eDbE1Xx0OBzOqjy/j
BmKQ+Am8HNBcjRwplUH3+mhFRLeROhe6eYTcEt+dnoZVdgi6jAfAaOJnoxNOCdzQe0JqCrMHUnIg
hdQW1JUoDEvQLxKzUNtYmbRuetB9vaJnvkC2iIapAi2NZQsbZE/96fTUtlGXSiFTPsLpGEIGzxo9
YfRI32p9opkGonRS3TAWM9lw7LLYr/q8pmXO0u11EWF0431HtGYV7spL2IKl9VQ3Tfe6QVHgPkkX
cViA/S4Gn4dHpGhjUKh9UcRiUATYyiykwBovVj4KyA6iPgsD6mpv3SiZ29NyO1yh8XcCO1s98zNI
V9y4NxbwFcFHFZC7+Xx6NOcuYrhC+olQ94xq4q3WZaeUTQZj+09w0yUdmL7FjVVFSbqw449Y3Sw/
2TgANn5x4ihJ/LDbTWqdK9x79aRT23+3XnvGF0jE6zHn/gR7HkaXgbaB7L9l1YGvy6rZxnez7Io3
7EDxeoEGPhGB3P7py9Qr5PF/XsUflssPB4ahxvYQhLy2FGsKb7Z7fOuJzV3Ddzvp1iTQPHuglnN4
nH1hKZjFrBeapyIMlIinoT4h/t1KgVpjHU001qSkub7Z0s7Thh/I+DxhQKJRZreqg3hso3y9PO07
ztxGX8c63u9AETkNghw2KkPBVZxdiIvHVHxzQV8BoBGTJb+PIfdFAZPFFfiy6FOBIG/mgcv5V1V/
1gzxrjcXFxUZUVpjda4Va13SSMOTXwx4VRa4DdtO2uotKL2wWOK8V27QCbfNsRraQM9PtA4lWvXZ
CJWxsJhcxrP64cTGeZXPcD59Erp0wcSn/EWFT7DP4GNZnVVu/RsG7dh+8XLQJieWqZn92lT9Q/8+
vRh3WftKP2hgoGsg/J2XO3n+SG5NXdT4IcGhhpO4FOd7k31OTQXDmt84ZyHI1nPK3eETJvU+COv6
R1Mk4eHCBBSY3XRebHYQQTfoUdAokksavEe8p084t9BXeNvfzYi7KbQ5UKqalMGPxPPPcvwOtd5f
thc810NNiM14f0PLUrDQ4QxtIvPIUr4NDr/+ErhW1hqd0tGAmsUOzA8VgIxTswQjdCEmus4OrziL
eIGhdUOkap3xkxqD3hizb+vz7+ZzBoVR5ioDvdteE4UnnjKa1yn7qhKeEQn9xMWq4wiKVzU2GhQb
ie87pmGtrOg0AVKvsBZshUgL0OrspCj68je7EpMXFbJbWNieP0aDe9ddMxFxAhEW8It9XqX5z4Sw
JRixR9EolpWDmdFnnSljK7OWnDTiEKVGEvRdBeGLttslRDBWugc33nn6bq4R0PBLXUcokvQ0gfLo
adn6+W2X/3o2xMfFqukJx+QaLjAtRSSxFlBoPrGnOt7IV/BQWtvM+HndnKJnNW4kESZtHaQkJ1Xc
2KqHuq27f9CtAw4SsugMIridukozHlVnSnuHs0OBRjLsIAlH3nV45cOy6fkaVqX3azym6pZNMNvT
Q25wjdch0r9NCIFP5ZuhlrR8QmNiKWtkNO/+29IMu26yhNqoTwfI9UQ87r3fzM/MiZW07mtc4RtU
J9D4e1Q+JxW8bjSb3WRmFFLtWKHiLtewZrTvRcu87TGI1GCovRjOBPsQMTyJTL7P2hNmLp/kZ7Be
NmXjEhFM20cWXHTZDNbhqVth98RJ+6eJjabSuT18EzlOWtj7czOSjZ01VGmBtEyvOwjU4xU6VVPG
QEqsFSGmOMoUUm59OArl5eusmkL/I5nROszd0xRCPzKuGgcGzVVoWnTXVZJ7H5S+zyuLwrPw1e3Q
dkytggSck30tFE32zdRJ14GsqbbP4Ym6IA1N+eupCvAwNcR0h45rwG/hk5X/CcnlupleA9rNTGqr
By5dX21NK+bya1EzlZKQd4yZzsAIwBmkcj4eytqVbZr+tNFPyS4gXupyvGp63uHnt4rkffWOOC8F
QNcqXAW1DGcDgdoUklT13I+SwlfdaTMkpx1XiOzQ/PUHHR61hm1120A5tQROYeQXrBYqe9vRLrUz
BSKOwWimlOn4ToDyCTWBlLkfvP0cGis7k/WH3vmug9gg44EwxfSjvRddw9OEGSyMr4NnxxALyYrT
sewglI45MjvOHazuugUcjGQDUKfYN1Kfnbtz5K1t5muGuXESyWabrfjsnYJF9NDKhbKAZ4moyZdD
iqFDJVdTH/Wk5YYCTtMYtaGh1aoDTUCht3jLWy3HKcPQQuNd3DFCYAHo4Lyg+hiVSAHQWvPU8Cnr
+dg5cMG9eY1PNG1RYwBN0I3V+3h7/eKhaxo0NyNeGqlB/lrE6jE6tvw54B+F0TjV4WOnl0B3NhCv
BayWJEMABD//igJjnTnM5nKRenvrujKpDkn1wFIwIZVdPFw09icn0s79nYNrGUBL7nm471jqZh/F
rcmDyCrBj6e/Xmrtc8+KUSpOw6qrZDRInd24kOdDMv8qADBdzp5U5Wf7xrkWl3VpmpjbdOxJQ5eZ
i10dsO8IKubLnehDnA5dvjYtMnsSu2IY3J/fV2k6xe5q254OpkQC4yFoYQ667IGY6+4Y7RmLFt56
gslw++IeBmbZ71k822rI73W2WYBhtIc4UIG0j2cLys9fwMTBcmPeck6gWFJMmus4VnF58rfxlqov
eXtKkOVZTP9+GHyb+3uXBhiNYNCAIBOgvDQ5qewnM6yx/3GAf4PHgsqFDubBmjzLLfMuwY6/+ipf
sMx6jfjMC6zjM14AeTf8s3TiHu+mZtmyYwTzZfWwATRvZrEn71tu1R/woiD6BdMjulCxertFI8dn
j3mq7nqwrF5bCLJml18u4qU5m6ygeBF2ZN2R+pa/KT70wI1MszjKX/WZ4LjPP1xp+00HHAvbMlK5
JFDLu5ETQoRVVQL5125io/1mUaoqA2/WNVmZa8D1oJLJerPc08OfoUiEu0/gETtPaoeuu/drhvo5
ovEzL3LYe6UWjRi7NHoRzq36pM8TgCAwE5fHegLCay+KYdGocWnmdugYN0O2oKmxCGC+JnvoFQpL
p/Mun6jV0caCPVCZlbY6mFPgXCLoOG88kwGX5j9yyivT1Y+b2lkoTJ1ay3zsdg/FsWIOBwSU33Vc
94XC/MKfpNo0aJ4YHM+UDvXENR2bQk4XHs0iTzV7kDr2EFP19Ke5+h3baCS9lu+3727L2ugJFCw7
4hqDgcgw83TARoyCC/PcvMVF7Wxat3va9bmIy+lDXi03+tLC8vCDlGy3t3R/oF3X09/64DH/Wu9p
CLbDAxVIUIY+LY01HYvRKUkKYtvZ7rpBE3qWm5o82JBnu9uozHZ0afMpS06z1V/HSEAYcSqikLsx
1xe9cIdvbsQAXZD23n0w2JpYFtpiYYs6eRXZsnK/GSFQm2+Pt+1s4W/kPkqwOz2Fk3UWEJ0++Czg
/yekekwA6c8dJIarw/GBSh9IbTm0J36LLb77X6u2a0m8bTsLLjf7wYRvyP93v/yab73oBbpWThDJ
H7Gxc49YGZtPLBOZT0s9HZReD9UUTGhWJUlEVPt1C7SfQjgXIygp4/MCx220hc7HuG8WKc+hpfhF
ojqazf8EdwkZKejTt387tCVEMUrICZKXfh7vOFHub3WsUR2rDhphehwzTULGjBVsA+AsA/Tl8Iwe
7Z/Jca0aU4wh5JDiC5+qchYyP3OgvS6dwf/WRxchtXMpIUuloTE0kSNRGSwwAGCw2JI4tSFm3fm9
wP7i4fQcL3ShdKbGnQ14tR0shir4KR2i8vv6JLo/oT6OQKVYrifk56+fzK65Sxf6uCU5zqJzTmwk
wLdDKdOtrWGpG9YzTYLBHNcwcvKUrv6mcaRfA7JgPzNL7kabn4kduKusoX293WhzwmcMmIvKtTJ8
8TP5eHRwv5sVO8ug0VuwvTPjH0Ja2H1/ElGRwpg4CSLA4GUO7JlhRxZQiTXg/rEBs4EyUH+vTNqj
IMirrjklFRaMERx2r7NzicAoLoTe6aZsGSOiz4f1XrN46QCl1kb7gCbqJLiksmmX05VGWPu+Ji3/
b9u2BbzpUcEEZnR7AEV+8ry0BmAlWMYeFmMkPiKTuLgMmUzrlvz2uWjFNOM6DsRIzrzH1XUO96C2
2avJ+FztT8+h9+9YJanaDHhTd4n6Fmr5yGG3H+kwaFU79gTNXl+bs8bilcWjmTY8heeujZM78FpW
SJ4vpv0NSopOPicTLlkYlmpwQ1/w9iBGbtjBVPyXU4jmcfv3GZvHi0NhLrAKO6qlUf3mWw8SNZDx
i5bmihFkhFSMNRVV4P2m/TCW6GktCHHKDR1276NRaFhb5Yy+WzWAsoCFc9z0eF+P8RdtzEwS2GOq
j1Tq3DtcQjxqP1JgMZu9YZLtMOOR9yZNxrk3QnEjkmhfA+502TZIzB9cIeqwJDf9eYo/LwmfIbJh
9Jtunw0pV18rUAPFpoea+fwdF40BHfFMS3qyiMWaLOWrUr9k/aBbYxNJ/lwrB+M/zbBxO00aMqIn
45imDXa0y76QN9UWyrwYoIOdtSDEf+rUJRcI/v3dR6MJQpIQct7DDoMc0NfByXXJ0qT4IJpq3m8A
ZDZH/VOdRh7a2yrLnd6MDVgUtxr0CgaqEudieMhaUx3N9zu1bGoK8UXzQzcF9uk+wQzvo4aKzu+P
p0TB9p1gMuoZbh3Mg4URbwx8H7sogcJ2beIialjzmO5TNwk2feksOIgZT6QvLewJ39trnhDEUJjG
Iim+Oeat5ojzpjGuFiOpSlUTxZ/9uk7tgZoqIL3msw1IkGLQiX8FaHOjKDEOzGxE7BmvEG9GijpV
p1NgBJjjLDomo4IeoPTO8NZdoJQU+WPYFQtVRWEPRJf43tCIO16Wk/adyOZ6IyERadRFroNjVpke
6kg5UYQdMYlddIW/N1cc7m2b5iPVzmB/bq5gHe8YpmRsMdwLGXY4jjAjAZ75d1owJG9fIyrk3htR
l4UZxfT0SoQypk03/5HiZVM0gF59Z3zLwZSWCXHe4S57Jtv4+peHQ2kziQQ8Gqt0fPHFMWE2lqYB
UxU0CnymcFClsOpKSHd9nkOqQWzot9RC8toaffK9HAebZ7F3Mem5yXAD/2vLW3rjbbJZqz0E7ei2
Y/wm95N4GrpdyMEPuyIyidrrIcnu8HTrv8i1V7UixcKVJg3RlvdA3WyvwynGLJfyw22Akm9ZxH79
4RRx0dB/r6bIJDKmwL7Hw8CHN7J1m6RP0DOrBV6uZphsUUkHkVbPJzlQaBxJjYXKNcAPZo9Qfji+
X1gv8ptC1Y5hLeSb4vvZKL9KCbG1eFO1kWGhIOg3MxFbb7zuUXi7sF99YXOs72goOUsb0SocvZ6V
IqLlU2QMoWH+r+NlFLUkOhPYvWQ1R6K/AJ7cCftbh4N110nLbTofHdMRMZzCPYT6u1PDbmvnmA0f
ZcFUNbGpUoBEMI2R2BBSyRO2TlRJR3kVb9TDPwbUllrDfxWfGDAf5YjOfFQD/jp4J52DroZJABvm
R4o/Eq3Ng7lLA99oJymF6Dswb5Ahy47duZe3Qr+AUe6gLVdOWWgdGrGAQN9/HOJqiBEgZVgI8y7i
RCfGjtn++Oa0W+VGkFaEXwfwcijYVzytoMCeM9VblZ6dCYEwPMv5Fp6IPUoM0INo1j/rVLUhO/Hv
S8xSpi8Q9BsK5Xf+Er4BU07lqjcG6Pg9vq3WuDk2Ilgbv9+HynpmeMcg8csak9izPvc8Bz+R3lGz
eD9MzvIsMO0EjF0hJEYlE6WFczWs2aveOATI9Fc/It0Im0QIZwWpbr6SH+MBTUQEh4kbWAGdfzBo
qZ1mDe989kVVsjTwsadB9Wl/20ZVmujGqscwfLg6RbMs/TbXuGRh0DpQosZIE6YCfIwkP2Dx6vQb
/fjEjTUpUzlrt0S2XHC5c1yyxHNuy0VP2s4PFL3GYo4bhhYngxr2YqnBqZsyESz0/cjbVScQlwrc
q76A1de7ONzwF0Ytn8QnfbBfpepZvbXnFafiGGENlrVrg+pX0WMLrXX1tt/fx4wZ7VZcCOic1sU5
1p9z9kaBK2Q6Q0M/lYelJIvFrovR7oltwVqDGaLnK0UZZro5BZ5zeDOOzeqKgElqmEPcwrZQuK/a
uKFScH1rCCSAd7lcS1qwwcyXzwnAJu1Z91ff+JgVsIP5Oc3Xs/BdYIDoGLz5HPo+gNQyBbRrqydQ
JscOdgqUpYjPGpJYsd9TQDQhwyYMMhCykgdgA8+FU4lBMnXrdfikSEW9gi5tLPHOmCmjXhubnDq/
OBhrGlkW1Ef3Z3+Jf+paXlTV1TBR7gz6ffrL6rgq0jqWwqa/fV+RuyDplWwsMNNQeWtF48W9xY9D
z8LGY99oZQZejTZkkpQP/V3kHU+upRjb5y/9JsOLwVYl8lE+STHsKuxBIvB5o9LLFTkvbgsVRp+d
aZD8OKxBA+25fPEt7ZCE0mij/9VPDoXy0BKjjJldk2f6n2GzEXxXCYRCRs+jEH2vY1Bl7+qEJu2b
S87hIqG3F6FYPBqDK6hpNf3Eurz9jhhZCYUDrpj+Vca4ez6ARX3sc9DZgw5KO4mlbKrzjMTknKvM
h/+VcD+JFkz/GPF1rCsDcIcykZCNn8ro8Hqo9kDQvX21RBtnU7UHxHu+U4VB1GdQBzKPcVW/aqv3
6JHkIJ3aCkEiKhNC8jt4doUGqqc3GzjR1yok6x/KXunlonGZ2tVthETqzF6FXMOyuccLQCGeGDtu
eEtNcMdNvIn1YMzxgShRRShvUBRxXqBnM+kME1ZjwZN2nqOsK57WwKFYNSceLeHrvvRjj2+m/kC1
UatJFiaTSRwBuhL8FRIsPeD2Hae9wBa6rkArYHvn+dyQGCtvRQo+akD1bhbpav2gQNCS/5wIDGdp
G3GUfi4sLv/fbOwsyWtJVsckpO86Vz9W22xBR4TPQoMI2v7EIY6rrJf7orMaDDFMtPpusrIwEX1D
PhEj3NL8FE8kuN0X5pcsbSEDmR79K2I3hOCaS5rgUqImcGZDiFOkpJO1+6wgHcAS2LkXL89svJjW
njJ7lJUN/+Q7b5sIMyH9BsjD8k9NaUNcTLT9FK8WqKAZNK1w2e8uQwKzGJW07+Cun2fojzbpgIGd
r2ZPsRg3+tUPnpJUV3bfibT5JGvJ16FT5fxMpwEBSaGO026vtphmi45J8KrTQ7ZO3bR17ptiLZN1
jI1d7upwbYhSCH40eBMU4mBJFxDPYGhLIW8Qh2CEfFcxbYXOC6FQIOadNWpEAl4PQ0u5VBcr3mYV
9cRNZ1uQMg3v0irm79MAmDF5/F5O/TK69nqnmF7Z55F1qVNKlCO5LCR9YypD+AnP26t7pNetUSA6
glPJ5n4SCFyI/gjEZxNt8cpl6Esfszds5FJC8CJKzDgmh4nIwuZq4e+faFSx8B62CwJ9q9tvLF5W
YHPJ65d36pMahJTY8BsCT6h3W/tIDug/gOS1Chk+tg35FtVua8GXaPDr4iO90N/GMVxMFq5Igunp
qopoAs2EyXNUqn8lv8deGBkePgYLRRUtU+GWQF9L/rXpy/Hc560MUxx5QxZY9WZNfB5uarUZQEuy
jNZHk2HxB6cGJC2mnLLNr4kVxCBb8QxoZVPFhfOy7Q/ZhSX3HzrbYsVUqPDSK7QGmna5yuK1ZLQC
ORCBjhJPmL4NLs9tnlcgCbidHe/9Q9q24JOrcYQwskniDubs57tQgC9HPfHkvJqd6VSPoelxGuzA
I9AvQ7LMneeP/7kZdaTJ9fZ4nxSwrvSsULtUj1XksXAbngR5qdOvauXQqLhksC1v/0iOp+dkwM1w
OjE1O4KVuu8yXQVr8aTKk29hAm37Qoo4QeR4T4d2xIVgNamXPQGlg4HEuDbcUr5zR6gPvYH5ODC1
6ZE7XRxO5jtaPiy8ilUaVWGqrqgOsHaUI1CYcXAEkx/WowZ5Oudgf4xw1YHLUhYr9hAYSF7HWMIk
1o6MMKGm+cbI7VMDJVKWxK1fi5aOCC7aaRPq63FPBHSjaU7U0o5IFEYRQo0WbEk2jelvgLezD4xF
4Nj4A4uUSqU5I6W5vXVz0NeLRO1DeChacDDpIpR8+vnK42sOesxywvVI+FWGWXK+nQ8rnAkwEqja
YFaVRRHMjU/k9N9nkUCk+SeCDf0CYJUUm9NAPyC/JrkDnxfqLiE/wyT5abPItlw+3LZQET0gxkeC
YcYwlRJkqH+A4eWS9FNhlt7werasPk1eFKDrLqKLneQWVfnT1GbHPtEriMpoYsKoTYsmD+qPgXcK
iHZJfUt8mMlHGTzCaBlAnmjNjAMViVPM42wIX2D0xh1p+pYzzm4eLk3hIeaipZ4RgV8XT5RvWu2O
QMmcnWJvRevCkFRa68X7SqKBGAOw5QHUC7AmIXT1P0FazJ/CI7VUiHuqyasVKpl21690mRd7BS9k
pEfFxDAD12mB+Sslvyx47U/8/Qr2+etP7wvkBqC987PMI4qr2FuKjn4Qa5Nbl4PAOoic/NQW5AIT
Bzl8wl3tmBDpf3uvZVrw65C0rIGYlglSKS30FUlh6ZpvyinwCcfWxJFAE9JqGxobBL2FmUYn5izS
VgbBA4+2c0HkBk147w2Z1y16rEGoAFrXjtB4uYh5lM58r5lA3UfSWN/diCCHo9RHnN4FhrSYfBeQ
373QpzClS4/8df6nO7f4OM6+FXfCLSj5bX6Xx0MyS2MVphMIh4DqDtSs0fxlhI2GYVdqg+MXNyWE
9lYDBAQdPY5pKGqmXR98Yqn2xh4ZaxD6rmym0293CJhwvaA7fMxmHbVjt5LG8JRk1xwmhfetY20p
6ADWLMFwI7K82K8e/T31z7PaxSKY7S+98VvmYUdAGM9lF8JaMkei7rZGNMOjWSestYsYwoeKYsll
vsRvrsSF9xqWx3wKQ4i6kkAxOD8GdtnRsozSnGw/5j4YZAq7uQXrZcRUL6sUbZigCBAAhzNgRvId
M5+Ynsi+dS3uy+hvwbdVyx5eIz7TM4r8T1Z3LpgdEzNIoWbiFvaLKaqLbOfhP4qOffRKLk+uxlxi
g5X2nmZp5qJwBe/xioTzgeuAGwvZqqdXw614iYrRdb3wjUgVBbJTR2UnbltpicRB6g7rPNWiPEzE
9SLRTek3o4ln6YZsODWcWLmDI6JLVdQkRhKK2b24GJXzwaANlWMuZI+zzyxaiVZeCHtl1ySMR7vv
CA8x0XJCtPAZ3j7ufMM7dpM0NjP4e1AdDhoGV5a/zPnU7GcT6AW7J1Cw3UO78GWtqIo/upWt7Y43
rfWbGjZfyaF2gLgOQBtMJW3o0joIaduCXwuE8ALLGw/x6h/2dRrQqpRjhmgKUwbh0gBNdBjtf5gc
ma1+1BAPnKVAYIkj9GdYbMw1W/KL4YPROMTv6ntsdH0r7exUlXLDPIbqYGRzJPqFI+F72KoW0z0k
qJkclvJ2gMOZj1/uQMAyYme4tyzaS3IBZ7oglxK1zoQRqGrgdhDKFJ6+ElXfGfNCBSBj1qT7ySbT
aBX9woQPxfHBDq8Fdg9hzNH94gCm92eImXWL61hzn/3vA3b2OvWtMShaKWzm80YszTNSqkMJ70t7
TJIQyrLvo0SHKqOm4TLFySI7zS3uBcSLEHg3SWR5ewGz/sN+3Ke0T/N1a9ERxu8LpCQM2FBMEl/1
+dNeMt5ej0ZtvLDOOr1yu0ahIR71SQU5vjrrdPYqJwusAwf1bcNCVYjClOex7SwXGdNn2+lB1osE
GwCDCrxA5ksnIbh/DIy91TI7krtb+olML9a5V655kqpddSr9nxRKhNUlSYCn1If8Utd6qhoikdeL
uvmfchePpI0fXcLE3YHhGIJMUtWGZZVPNbSrOp0c5w89ex71llN8ApV+6DLGtqoAbcDydPhVBX8e
Owi7UpJQJHT7fVFkTn7GJnBNK+CLtdAJiYMH4pZQ8x/3QM8u6UXrSFkSZrc+KlisiXIqeYaCpOUp
6uYiObg+xLPAprGavkTnSCYL1t7eGEzNpEASMw3YQGyY6YmAc9o/qJqVyRwQYuT39GMXdZOcp1u6
BOku5JWWbwTrp4gSlH57X8g8sA5ccFpthkaa97nZWbUIaMcbc6MpL4XlMRkcu5V9UJMYupuUIZg8
0XN4Z6HpkEKxHUkZDJaOs0kUdN1VtGDvd019e/K56uwmhBavCr9b8eEfp7rlf+NE637DFD7UkKlN
5b1tMJDX3Qz5hUGeSKNNKF4w1uSNSLQ+L7B0EraN0TxXCD7e0LLyiF9S3qnmcV40nBqNNrofs/J6
mKjNpy7NyV065yXDfPiwF3bJql+gFyC5sx2tWyODMciu7NHxT1sb6UFongP94NDsOte/A4RmZCNG
IbDsC+rd99ozZ1/0OrTPzi1oCUbrrvo6piCEtg5JLWLLVqLVy193Tp6b6GPzpOWooiCmwjDjesRP
+De/T9kkmDy1hNPdFNaaW1rLex4vgvqbMpOCULfn2m9TT9X93b43LuWXG/ApcU3CroKMykxEvWkE
QTjUs31K5jF322dG51nfghOsRrkl+/6ZeAEcWVutQALNsZmGJDU19tAUG0MbsPHRNzb1FEao94KK
/GAaBzxG8/GqyF5gPLe5hbT7RmtaJQU8fDcXKGLrkkawuuYpsTibweSyVsik9yWuV+ug9jcM1IDh
pcE+CQuTNgR2ERBKeIMxm6ZczWMdutrkJLpeDXhrNqIyx2l+WKgNAOXuZcfMgjY/tR/URP8tgfpA
DdJhkoU3T6qVyvwlBVqNfA8qNcg43BxQlpYB5M/ke9JVNqzPtXIYO1k4A1wkdT6u51UvOW1WJgOu
9zIGasH+cO7fMfm1ZpugxJZhCZZVRxMz2zPjx4+5P0+Z7WuTqA4/+bxV9S/CZMecbVjWrbE3Idt2
DhiHFCCEda14h/eU2+9PoJ9K9YqjV25imRA1IOrHU0JogaZnMm4/iN8UcmqdPmT8LGK1E32W9wTR
961onfQw825f+zOT6PiClM4l7gFeUY4LmJOCTg4NEBqK7eeoaVVmCKuBcwZRZ9KILxrlGxy/PJuC
bmAZsVurKx9BKpHiRqvgsQWuQTYwFrzb36U6SkQ8PoRaHs8/nrv83TzEHb3M9PhF9m/9Ww7k32zH
xEbhtID4QHbmmwEfs+ayXmkVv6BESX8VZH/E1os0ZVH64Wx79ja1ByEWzfxY5TU7yOOmHcXeCd6o
uN5WL6OW/xCK9J+7mprnUrvaLPLrt61ZTNzYIqB6Ot42IEA9pMsjvZEHwt9/SeWVxzyVh4If17Pj
V8HqEGVVRaiJ/PzGBY9LwkYk3rqNzOLmf3D6rLVRXJQTfxG2IJtTi28rJk0oc+8jrUn/Pl47g6Bz
J+jQ879eTqAo8mcC2nq/3XS/0KvIc4WVxuol/R2bxzwK/76n8QRs7OU1WsoiCAAHw9ZMKJgfAkna
7cpIYKJpA22Eeg5IJ22hUqQ3rGwqhY0X2prjkMpVUZPKb5Ewk7FKdb+VZ66ZOQmVbL8c9JBAfaEn
k5CmZz/o4txPhfsX4vWvzlo2/XZE/Isp0EwydMw54T/nJ/vMCBJza4+L7A4VtyzBZGfDiVyKT5Tn
ei5H43RVo6ZVNzb/qTGJWwADo2PG9k8lUmHW5gZW2T4FdwpBw3Uzv/sg2Gf8t4aiuhYuhw1xrSBH
VenuShPjIp/f9SAYjp3+DxicHrBHURN3lPLgmR2+HkoBTdqpIbvvmAbzYaLPIx7NY2ec2lF0LLly
hX3oXMsLMApv9VHMlk/ixZU1dcK6H7dkpM2Wscz+utjq1ORWNyEPEMd0cwVtpfGwKdSab7jBYHXc
81K/0n+g/Md8pFnsIwRah+EFX0AKYyDexd7Y8jJPlVcD9188XftF3lbOUNFZQ6IFvC/Ji/DFLDtI
RqQq3aUOGQ2zQhKCN5prF+xwQnwZVe6gAtt71N1qm3eWstqFrhndXCPJ6hJ+dJtOiEUxZZw8j37o
liVIG4dzOgrAQRFFKqmeVgcefxfLJkWir4M05BHj//9ce7zXYo35o7OoUoE3MTqQXKxMaiGPQOFA
zS3zGXqQ9PQabhv+CXabSnnrZVgwGC7hHOIfrVglTSD+WthUhB4P0/F6FjC9e/xKSKnfuCnBPWBa
LoNm+PZJUfhST5GpuqSx3bky+gfF4kSgHgP59IwkNwkld2ONwscJ5lYivZ5eWN+o6sE+yc+2MtbK
684xu+5UZn0ObMiv6x2WoFmvfNG+MyvSbcetukw1fhks8bFhOWAuPE9dYaVcRxyFtaDCmO7wK/TN
vkcmyT/r8q56wbHJHrepl9rVFJC40gj84fc5gVBTutN6tW8vtnrEo5uzsb/MMJmQfiF03X4CKj37
QbGRg4JNTMR5U6w85eAUxdWVROaer3KDtzMCJNSqTBNe2NXIWm4v94pZrVsfbIVH++xnORPBCBb0
8Baoh9YVJl00t2kZ3GhBhJXz4UZqVtD3ERtUv5ZWXA8nWDcWMyZeiQoR1nRKoUOViKIL20ODZIDI
xZoQKcneQgNsqLOEQdHhl7YsPI5n7ujq1kngvJe5pquO8RYBgxEcg0d5J7x2NlGPL29TQdhZdFvD
bqvtuzqHdMBdf31F/heHtST2hCQ4kPKvXex3tvngi0qzf4jNFTjqm1L+wGTQfo1YlsOC4I0lDGWg
DM+TGgiT16Q25PhPdDBCR4eA9Yisx3egIA1QNiIzM1p448JgfE/Lu3PDuMCcbxSkgTOJwV3dUPLl
YLczQ30GnSpFR1ngdAxxIYykxkRWSL4PkynZZ0p8IfTilBzUogOYD3Uw8BnSAjibgbt73Hx3ruAS
DPEe6sA8IQn6DX9YACG6Go89zDMSZohOd6ga87N+q6LPQ1FDwJujzXXeP81QSXD3vwrfo46LryK3
snLLv70bR3ev6QC4Hr9nHJ47+h7m/ccsSDX1PJ1PWaNMvsP0i8hZ78nE9gns3/8i6L19Dd8qV5UB
JvMx8Q6ioK5p3C+HMjiW9CiZTe8zO8o9JVXctJq8aGbThlSGHd8IxWRT/U8eleaSXj3jbRn3Vbtp
ndN8RZSSKwGLCjVW3BusZCazCxm3TpbTvhUZeUecLNC/tl+e4RS4Z1iGPhph3Z9PWV25mlJ1N1h+
9HPhWG7zjRtydW8YeS6dW86dwEZecZ3ulzVOQbhRONX9cY7Ce7Uyx8lNQqdJKmyQV2toi+ZUf7tG
tvb1aCFZ2ARmvb8HdKietypx28+e/1TFFqZQxzUN7HwQhy+UYheyATMcguhSUXbf9zEJp7aEa9Vw
YtkiMTxg1USskMsvkT/DGOGjpdRdYpTesDetY1k3cjOvgjkuh37MU7zEO5a/215Q0QenITS6Qxqt
WCIOpZM2g+stQi+apkeTWRNWEt3BuO2z/vhLotJ6lXKqi6ovd6UAMcEKQxnvBDfUsG5wX1CeFXB6
zgVEPFSa2f1iiLYnHKZe8jVJz61/8bWUn0Fw/Jir+x14LD+IJ7xXYTU+vwhPR9a9X2WEJ0gSP6g/
bL+mdBj3fiWHqRfApeB/Q7XcTamVDSSH0dtHkOf3onKe5+PnP6i7zn9nvVRL9b4FRffnSZvIiPyB
VTjxJXAtlvoNN1uEOei5VEZPAlF1uzXNWcmZvOOFFI9Tk5E5c9X5G1XplD3bqN/RA7ATOkFJ7JSr
Rrh8c4cweF5170EpB4r9ywv69QRo9nfUXz2G43oS4Vicl45pGWKVeE/Pyy4xLAVvQ3aIHmd/YGgv
X+Kwz86rXYK4TNBgefR/iSvExvxbfpdN3NvKBq04Va9zkPEN7qBxOQV8tM8XSpo4ZkwoDmY3B7/u
IUNVAng6zFPKF69eVPq4KKhC0wcvn+sa9pzl81pX9x6dPf9AGcvma+bE22cXS6RelLEadr+aXHt1
WFFn4t9xY6X3rH00F3rC4DWFPy+IB/nje3dksSKO+alkQPVas5w55Y0BOfd2hGzXAeQu3lx/ELVb
HipwDEx8QV/0ZJ4rI+P9BEpBREZ0gPcIH6A5JUytrAfIqonOJHAa8Njw9mnvl7uSUO8RUoAcExFQ
pio7zh0SKd4WZNeHcPBNve/kTlgNo2OWnxHSJdHj/XpEInfxGZOI2pb3vgWXSfBPPVlhNeGkQY+j
WF/5SJXPLfu45DHNfVdrYMsIwLYJt92pFu6hcFLKXh+snh3RYSi0mcoPqmNBXJ47fUwKgXkjbVp5
pPm5kEHUnFnLKvpBEUAesYV4PngZNqYlMBRLED/j1jUMKBiST5RYqPHGhuYRKSCjNYf4QLqLbO2A
BfiXxNp39GcNmaj/yyzZbK4Lnq147+Vcori+K4hKoDrrUiCNu5Yew4V/nGSWBjdMrKEvOKxuFOcl
3MgzAVmnolxR4V9E4DOwbUCTtLhiokZSHzI7TQ0jSvtOLTBj8XmHBOek6oZWu28+/+8vhdwSBs3t
vOvuFlIrvBx4pY7/vujdvEySjX6QTYud0IUV89F8IgF/64PxyM3sz5gwG7qybI7LWs9tGqQ0z1cN
zsAzu/RslFUjl8TS8w0IIAC2TUYyU2O5ZuFkqtSSbHnK5ycqLyLXTV2f9g9zYOjj/uNP2NgSO8oc
dZQD6xvWyWQ8+PHUN76OAv/0d0v0waSdSuCyqErIB9Ah0OIPa+E3KP4NfacD3yc1jX3IYCvgXwig
Hb7vMUHJUQoS83bzaqvhbE2wHTqlY+XOf3FDSUIuHwtTZsab7aAM8ISpRQA+kAmX5iTYnzxas7RG
FhX042kKG0zVTzrkUUzSuhf6mwLHQIHvXXX3ZXRpwbBM3sfnB3yCqsHNUmJVDfvw/Abu89Pj2y+h
bveYtF4sOre8CnRB/Ew1PGuwvacFnoJNBLOJmWq7L4uh/VwD4k0MfsMeScxjvgWXYtSlC1gZDnJl
L3aWynaLe7nWbDN4yX+ng/D2Gqn/fxxdC7TOIYVWW/l1IGzVbPZDsZN6zRZgg+r3bpv/Bsqtq3dq
EOHCoaBAxV6/9d2+zSeb2RXHKbEd7nGiQlHTipoKfDE2j479EzGkCUSt4lbzfXLlojEtrYdaC3Ix
8S2uY1NFgNcIbtYpNvuaeu9kpYG3Ht6vzRecGM/HsagmVWP5jkOu/kKL1S2o1pVOEHvS8nbe2NuC
x0iuJ5yNLa8sY1NvTtI+CZrmHol30yLoR94reouXCT1kvlvJH+/aGayVLrACrwue24RVc7aS6nNv
fs4tuxdeShF78f7Pe0v7OD/KgMZwPk109USCUtbanDlzWhs8Lfc52kz/I1AkG8p94pdp8x8l4/uB
sEfesoV31kA+xREukAwxRJMqyy0sAy7t0aji6Hn2kH5+D594zarOSURLKkkkTN/6lPyA2DM5C/An
9lrBDQBVO83Dpdcwmkwrd8FjRMnkkiMQDAB4joM0dhaSn6AVsmUAyPyGH4TdbBqcACFbQxh2lzLz
AwwS53w8u94XNk8XLR5Ar3hxRuOdeD46QTrjdKbA4Vg1ICngL/DQF4zfta/j6XP88XDBPJSgp13n
exX5p8XPDYx2QNRL+6M94pf7r1Zgbewn1eodNzKMyeDLXcCbtP4XnkdLNPxYyhqPiL7oXxOMOdeF
1TY/GiH47dJRcb4JHJd5uUdWjeRC1yqTIFfMKarQ2wEg9znreG29F68cmBrpVR/ZWBehFRvfALBJ
ULUspo9zGSdfykeC/gDzd+dtH4j2xUHC+U8Kofe48HvGyekxuMVhZlw4Xg6ork4ARasTGwWDSfro
I8WPguTuYzXWnS94NahC5vtrHULGAcEWZ/fBSJ7PQnSMkxX2OmMrMl0D57htnvxB2hOz3tfGkihY
T9INftTcUP6Ho9OcmwjScca0TFc7uIvpgYb7CxKhbd7CBk1juBraJVXGkmAlyWDvdGuUki80WIY2
w6UPp1Vf+n4BzgtdTYnf8dRKWa9bkkXYaPgO3BeUG3lhNes1shBQS9vdsymZ3nufqCsmRmQ3XSnV
g9l9aZW/3Z0H0O211WtepNEi4rKM+Odz/pV5heoJY5HsiialEylj5HTI9XbCbmngG8ZIW/i3peUe
+Mo6v3P18YCy+Rb5ep5GVHZ0o+nLycaykIRBh2AyFyTsEXOjhBES7xmLXrQHUi4irXh9TqGWn97y
LYX6b9un44Ui9knBOAwgY67pC+/vHyHSIlF4cewUZgTCd+QkiEwHxZeOk9Y25GH+742UqpRyUowh
haMfJw1Q+dL9agANHyzVN/3wK7uBtcC8saurZbGnQqPAcIGfRaSRSyOPuZLsNbF2DHzGPrqOiGG0
djoHe6tijqLXXGSAXUFMWtAL5qgI+rUtIBpir+AX3UFKI/qsaOsyjqKawDpn2OU+ByLF1qeSYdc6
NbfIwLNfU+ANctux6u/viyErDqFyigqFKJxHZFgIk0DkCzaFrMttjbYi/etdyk9koTV8Us5OOhxr
6bibuGRhNjtGGGdIDfN7n5L0mTQSLRcrANPrm/+poynjZL+U+5ccQAtdlnqelLK3qtmWntmW4vjj
07iO5gCCrFN2TVk/UHt/JmhVKXh03oA3jILIdRei2rwHlF9wXTuixxQ+L3AGQQIC8oD5oDlz+e1P
7qBNuEPM4sjrZ75a+dEsG6Ci3cltOA+numXkNlj8Inxwy0jOCaYSURcgc5y3dbg2CgLea+EPbHao
25Fkp3XyqfJs3FcciSEqnx16/yqqmYKp7kmcz+gJs5qigoFowMX167GEJHpfi1fVTFxfGuMF/1EX
Yp5I5Dw4NuoFAdE8BUHdaugtglRiD7eWTI0fk8Xe7B/7o6suuAnZTUhEpLacA9cYWBYtvSkaJvsB
6PmHRZyfuB92FMvRadkLWZGJJL8WdkqEiTZEmWuh8boyX0gH8b6g0eh4nbeBthoKak56ReAkiYHd
Nr4m8jt0t75CalwyDze4Vfce/kHiHBpyiRaCjyLDQXgBnrSzvHEjWHAQfKCg2JiOsTMDEA+B4vdq
V/dCH9jx7LhDy0h3vHTxQclt0OoIwT4t0+GPYR2lJ6TYNcrtu/Rm20Kv5nw9C6N4fROJ/HkTYOAM
WOjTuxPfyCv91+ihcciCXejytdQxSNPH35UvSzbbbDss+Fux22rMnPBZhVB1DpWwA51XYMF30QWQ
PS0ODsGsuwp4ONZatBhFcOPA5tqPY+eHalgXjSV0yus34JDZefPN+yK0cYNiy/iYcyj3XyHzRhzm
qzj52b1UXGc4Q4AJRCi8TK6JqwRZmzNpi+YRKZGiamSOHXlc3Hd7V+pXf7fC07T2cDsX5y90iIm6
O1BEGpuTkzMoZnCivCqIIYOCcnvIEGxunztunqZ8qNjc9pKXWB+rRQr1gstnRm5W/tk+pCvPOT8I
PewxuHKJ7xc5/A43JJXURUFlEvvF2ZFn68yP943IEv2j+mhIQfTHbl7xgYhzJ1TEcZEGeE+tfaH0
LDLEJj6w4QuaNjc0djSqrZQKiSciSTmYwovENxKi9PjwB6S4SpwjD4qRsE0kZW9DeHcQ0xHjFqci
56Ey9EzSgFVTMtiDXX55hJKPlAko9KSFeZE74lSA9r8jXHlIK1rUbHHbnxTc/Hnl0LGGSPZ/7w5m
1KEzYv4p0vfNNna6k1vwwY7CrLvU5RNxyrOBQSc21V14GWwzvT4p40ZCAU836MOdgWG8m83Jj7YT
kU6cRIhVYSnnZ3gGkzJeK4ZCIgp7sW7MZvuR+NXcQC8SqYXj8szjLBtLLd+mlas5AECkjAYHRd6r
sqclWC1TlDgp273hTVt/pcDwbqnTGLA4rxFvEf6pRut+w2uJO6WQ5xgaIoVWTr1w9cmoaScfunFC
KAM0CIVDv6iQ39py7gBz/XUF955Y7IDtF4GmR4eyfi5wmfFnqi508zEHQ9P/L86zU1973O4homTY
pPx0CHsPqSBPGBAv+9FvY+0MrzHPoLmgEJPrRAJVSthKWWwGufA2/7vvNfrY94tSSj9wsBx+euAU
PxtBnVFZMoJ13dfDKFVVk9y2VYkYDQdFDWzh/MM0j9zFhZfvpUc9XroXGWImHHh5fZEyOZGwYVCf
gyT675YtHompzvukeznsfDMGOCUsPDKzlzSMe5CALkRRUE7EnVzcEOKT06RxW8k64RQ6s1kv1eiy
8fO9Nub9LASi1kYLtbe3s0QiTlHsHvnNmdAW5TyS4LNEXyiAYSZ5sdybyrVVJPRm0gHAeCX7OUuj
OBTC28xA15UziOpoQFesphwmHlUIbODcCWOJVvwfP6ve9CQwYJvrc/BGLsQB5N0n1FQZUfYKZ5he
4T5uC0S7BPLNVeNgStKHIz6BItef95rxYMrGEvdDucFxHmxWH4+zKi8qJPClwQiVimKkDTl7Fcy6
l5+HmVc0v5PTISmEqvwAmDlp1v5rJc0Uc7p+ECwIJ2+knf3zDAYEzVSJIm+RW9dl5Bqqd78CLm13
Q8od+5yQtUvuluVG8+Mf2G0h9B3RWOxqSn8zQhD+Qz68gUxqSoKn0cxvyq6tQv7q+FLHugWkBAJz
L9Wu+Io4TYR96rXhYA6ej35L4R8obVX1eA3K38KUwBtO3BOrIPvoOTWpt3uV6kad8CqdU5MrEY+q
OoIi2SczxtcErohBetsL+WavscvSsWKUMoXrlFQq9i42gh2a9/eNexgMSNOfE1vZuxK6LSP38blD
ytvBfLzz5hzMnUbzQ/9wkOv0e45LNAxQfgFBjvYfiQ5YK8S2MXFBUV4p7RQFVmN/IO/y9miUpZzX
sR/LkUvM9IBkbt5qD1oJCZxh9MgLLDBw5yIYplKXs0lfouNR4XaowNI0LLlMv7RMvwMbPxkYjRln
EXIe65YaBxFe2WBpKOQ0xQ+Sp6Hoez3OSe/Teh6sLB47uHa/KFjeFJn+m+fCsMZcAYKQXQQsAXsY
tT0pyQNbt+T41FLNtqlFBzHLGZl2MeYW0J/uoNUzm+S/MYtxGD6MQE5BCSPtrtdSknoxItRTL1k3
vooCLbsQMr1F2sQ/QkNAW4f0qjNrrPUejO1WPQKWEDdV9J+c0dA6EvlzWQoq9gFe9b4ZWDJDEnOy
DdHQwOd9hAOQseRR1C7p2abHqboLPaboSK/w4qb7pTXzQ2+n4lKRjPjf/bM7XnM2RqocHPw+nBVZ
3+y8oJNMyNA/tav/tcGi2xrlbHjRsdi0DZntDfMeOwl2veZWLFYVVjFUjBbcqa+73H2VHSw6ok9f
cGL3ne6DeXRqtoBj8Q4zahdzd6RbQRT+GnI1o/Akv/tutAlZjK9uzHExFzmkQMVGeHW8yGxqQsui
OuMknigI+cnEeWCFtklGwDL5abG7YIv7DIAYNW+RfuF9xFQMrL5Teu9ZspAquNNcgRw3wd+7woD9
tDs9j/tdWLEaQYlhE1N8i3GABDMZpJyMGWU1+f1aY3dwwCuqK7Z4GdNVyaW3foPdCWcFgna2GzYK
hx7ThxuzcXPRcRDzMtmbCEh12OFQGkZaxUFxdeofTogkAvhACAsFDjotaM4QyoL1RXjYaa+nwCgX
EBQAmDZ2rB7Ylssg6g3rNgIssuODgTwNkifAFP98AE+DbHn7D3uSXVLAB6F4bi9XW/U3qhI+vJpQ
+ikY7LLK8y+dhsqSJpPy8ugRE3+3X480US+Ckj0gtE6C2QbQmSCNQK0w8rjHrdmGiVnnXJvCyUC0
XgpPgSWffKRN0M90ZrJjcACbm+ANOaSLbjkUAbWmHu5dJQgDX34AhE/amthFMinoaFx8i091hlqg
H3/28qJzMQRCZ3p8qk4SaxWehBeP3i7sSB9WEw1tP1ntxGQL3/1qrbv3V1bVhB2t7QtoUI5QKTr0
EloVrG9aBECMiUbYGcrRTTdqL6W9obzEnOob4U6vO8CbipWI5SAIfqTLR8s09ojxl2REJKOCLd3F
nP+XKuQrZwJ5L2Q9TcjfN8FTGeXJpHoFw+pLol6f04WE6MlqlKLDJJ5dNrwCl1t4ur6LWkV1+ri9
ACmdqyn6Aki5z9uZjXpfV8BXm6jsM+7CVip9YrMEXCD/Fjc/y054yOjyCs2HV8DIPryWtr5agYpa
7bv4lbKG+cdkqPMZH4HXSwwJZ2cYzoM8InMFwcqkeujJl5pm2hpTdYgtwHr1Yo6hF9tUsrG5mmNW
yMxtZpFDIrDaSjE3wfVnVxA6HZhZCvoPbpKxxjwFjzmQdp83IjAeArakWEvVKHly8vYZjRpNoBjT
V9vRT59i0uo6AUzdPrFqzmg8JakJvJLtiBEOfqzud+jTs2i9d7F2ia6O2FqdFQiBvly4G5sCnvGI
uK8fN92oH0zXtKAfwNS4unkrCGf7GNbcJSaYGk3+7CnRYf8l+wpOAWRZOoeGvwYpvUnzltY/Ldus
de/DEm3SNunYv1RrxuZqMbezDcZN6gDYz/w9QIyQdZjsGeZ7SaXBlSur1QRWhlf2R1iZXsdAZs38
Pvi2MHqcdJqBafriut22rd+qxWpCG1M7IzyBwY3WUhKEF0SGdvhM6gPMSONfL0waLSXVBNXqpu7E
ILwLi5gae4m7cTyZuJzfRiGsUwhms/6XC25Is3CYBSF06F8OPj2HTe9VAc2fJo8EZIC6NNbB2YNR
oOkwzTjM49LZ1GhJ1jsBzXyrliWt9XvbVCVt9iD7v1L2ZVWZHip7NIeyGRLpLEqoSKGlOd6UkFwq
XsKPjQ8SmP6lndKQRjO9SoP2UhBoPNDaRJ1AAKE/M2HW8Vq0AO16KwN3yYoV8IShRmC/MDiWXgBU
aJPTL84TebaMHNtaAQvagRA3x1DUXuOQoPogZ5FjGUa0/4AsWOCgv3OROQjtBMS85tX58riJZ38Z
gHr0V08HUTTabNZprVqU2c7fcXImcP0iKck7gL8clOJUcKvQayx9wtkTMpxF8g3jvIZnnsMUM8sb
cXvqk12hmynOJ6Nuf/2XLlk3Hd4Oz3InecCOdugxKUGg5ha6we4DJdM2Wemcb8pEw5knIJRzo85J
I6hfM2wqtR6jkR1qhgRwspbPl1cziyPS/+pZcskd9SXSuhwUSb9/b66hdlgnj5EDza/89KHole/h
nV2OCgatTaU/wjeh1MY52bnYpTHD4JgxTqVD32+XnnaHV+KwC+lRVxElvRo2+/j7PnoUPxPSLplO
EGU5fecBcPYiM7ED6lqzk0yQi7fQE8IlynkESer27TEI97/pHdR3yPW1N8RrPvFNZ9s8AAiyV/MV
eLbEtQGSYFjcYwLxjeszfGBdp7CWuaspAP3AQW7ZXAaItv9BPSY3DkvlKXymDMWPPUL0iATN17fE
/7sPsxT4X7tKBAq8QjcJlrh1l60zCBAnJ8z/QkmyWbLdirh/LaBLypT1sbNLquDNWLg9L6mM8z/j
Efuv1sldDf8USmjgQxCb0FtfYEnDGCHxlsdjne/AM43v8FZqR9ByGjnmQusFdpv2/Qi1hiz890ks
/5pcUMtsmwf0ghZMJjCr7DMOTMMkFGLID0Hbhoui0YQJ9moxfoce21OvxOv5GBtvxL/wRJguHZp7
2JAzwokJs2MsUHLwVCfQKg3a0tRC1a3OtPczvrzB4gFrH332c3DsctlceE5b+JHB/sjfig0VA8uF
nY8+cArM9HD7Q/akxofa5o4bMykXzinyAEnh2Oe3Ys2Gqs5fBEKzYvZFK0vL+/g2DBBPmh61aUUa
1PiO5dfmtyKiUQQdUHHYmJs0+jBFX3gTARNbaJY0pcYoHeF2Aai48uiIwRoIR5sPrkadTbQJMG4Z
eVqqHiLQ+0qwcxq0KcI33EthzowcqmrKfwXUAu0qYXVErb+qslKbud7+qxtkkBWFrpnFtHno2yV/
wthpXwDfpxrZAqm1vJPgS+i2vEAAMvPDskEmEskqw/3ho+oOMmn6G+PiUarLUpbstm+To92VbQFc
XBxjSj8gnbPxLdcd6Pb4RL/sCBiDpY2joKOhmb28dnAUpOBkAKUWl6h1W4IHPQgRwZ+FXT+2q2de
NaVPvCREbbuhknreBS+m2HlAFJwCrSXybwwCjUf2k+uCl4aJEO96pBW/Tji2h28nBEz119Cy+/QP
LptApGZ+eEMPcpZ3TsTntSOjdvcL+QHMYD/heEQ6bosAXLG9PJkjuKazzYo3/uL2u0mYW8jZ4leK
+jMbdtTBAcjq4yHZBJtVOCR1oblzOABXg85zATmLf3cixFi4ZL2z34YotnMVoo0kEdBh5AeyBFqD
y7vpelA32iefU8knKwo1bkAdn7dcpheg6LwdSlXfg4nQuwXZkcaGg45fNZ+ppxeFLEqhwFoJYD4c
ijyLLUuW8sD2PX7o45YTWZf5QSrHDDz8e3FUPtA1VhpfZfDwAgUB8Qzmt6iWRhxZM4iRhw0SETvU
kOaD77Wi1MhGQYPdpKXGPCN9/ceg/TQ/rGRRo3HLf4IHGFfE8mfFJNUG7MOrZhPS4TAGEm4wb2CA
46OAGFun/iffHZtTmJ4oxkZlBxU736xtKWtB2SZn21VIVW8ii+2qY2Rcx5P5rsnuvohLanXb6Cnz
eUO0ffMMTSP0SNzMphbiWrrUnK5hs1JzXYMGIgWTokCjisrg8h9e+nbzMvXlyRYXCLK81eaD3tum
/1EXJvgMu2x57YfPS7LiDgfiTuNFKUB0mCVAUMeNNuVZcOAUlUvnL1+0SQ6Xn8RoLQvkSDU8TKbk
5VjNTeajTGCa0xlWBZM5UQ05VwfKBfCsI7JX3f9eadtIlk9/iSZc4N/Xd8hHEKsnmdbUD90d7sxU
siTehXNwwSpr0ugnDQzaeV+k50Nlj//FjWuPg1UE5mtFFJlPOv0tSUWpoJAwSNqlr98ZbAM3dNRx
/Dlgz5EoVdwA9tVsqg4KfsdGVH9DxCZI5RoBxfdlnmFj/1Tv9Np4EGWrXaEe1F3xJi0S8eJGiiBG
n8aZE2vCSaMi9p83F6T3oNvKVjrbAsZzSK952W5yHIPZ3PX7cgiGF6wipGxVx9kOk8j8p+WFKDjj
+Xh2y6wCDnrxKmg6NshLA+YjlCqjuzVvwEUzq2wNJN2U9BvnAJPaxgl/Epib6P6mrqlSuOX2qXHe
jpuq02O0uy99rC6SIQFbKwIKR4BrNG7hY3FLJcpSpSFml72pRDaqOaR+Kr3QKcfnhk/X1EaT2Zf3
gLrUNN6dbjQQ+EbnN2rnzr5cYeby/zxCp/rbHwhFffBHAA8olN/WPUBcfVZa+CwoI18Up1CVvyIv
3Yg86Hmd2UE2UcEEofxPByjrFMOa1slDpbmMp0uU/1/Hm+FsPeR0X4P3y5JRB8kC0Yuyrzqv+aVZ
w1ashCsbgQEV2+znRX81i1LvzPZGwgnJ3cM2CGGoP4XZUurBWQoICxiuk7CAICVp9zHYYXAui/0C
dCB8SEpQ5MXaMwf+rz/PR696bt5i8D8yZ0e+f1bEb8P1UsGBuHdkWf4wEJDbNZHjGGqSPJtguVqX
fCZqMTzj19jYL++H94hggeeT5XUTBH1VxL0ECPDmcHDZi8gDNWzLTUPJ1w6C+9rlHl6TubH2EPZb
ER2dGrZ0wzMNDPHhpBxUaREiZ276vQlJnHfQpEWi66xPB8x/I0EtLNiDAkUQO0t5HMLiQmVg8tH9
OrhPw9OcDbkPntdmoUKsVFG+O44HQNn7gHvELpWbPpQw3E07Z3kn4Fb2Iw4MTkq+yb3hlG3W7Ou5
EmIMdkTi7gOZOToiWzu6emAyDINdz9soPj1Z19XSezEgl6C+fWBOYrfIEkSStJHv5vkXvzGt6obF
YXwDY21YhGxDLI+zt2V88HtIGfLKYri/jHIKb9wBn3Q071oDrKrHQw+vZhN9ZGyf+eLWTatYo59Q
W8jg+YVsYXdoI4tRPX7poFYNjBJxrYWBewsUftLl93wBy7Pg4qpiHwno2PtL4v63vbg5zDv8pRRw
Md2hZKDvWRu3+QuH0+hZnyZIptNbhfUqCRV/OcNia9PFTfcPiljTcRHdIUcc4cmkOkq25I3zBvao
WPwxpX4BYMVoeNvNYCaUBDfglN8gVlxmBWUFd1o+DQmfz2Q0gNayG55mNj0YSa9b/9wUG3YHfosF
1xl+MCNdr5bCiViIuYVN5U3B+pNO8IqOiD87dSdqHz9N+ksgNGaIjseFJFSttatCYVkBBVqp6TMf
sh1JfTIvekkw9iYeFZyPG4DGSjVZPuq7R28zj+coasRHJYZZ22kaG7MvNJ3bRdwCyTmRt1TKfDte
zSSBdyPrj3dXsEVb8Xn/4TJZcOd6JxXB5CTjeRCnizcnznn98zxMy2CCBMY/IH91y7o2O4qfKfwi
Gc7Uxg2iPaB4tR6UNaJ5HMH7ejatlSHbZ1/GeUtBSFlSTAC2e48EU6Zhf9XNk0n1Qk0BquLY1FUR
isINbaydLtH8nwVqb+aRBCA5dTjmqRhq7+EhQt2toOyQ2FkVmlXpxa09kPzXy7TnH16kP93S0B7+
3qHN99xIObpgnn0BBze6rXsFi4RHHLprBJrABlY4LekL1Xwl2IN1eZ8olsNq5zO6HaXRtxamT0o5
oIXVKo0NFHX7jEnq0e97lzULsn34ECx2Z+rywkWqjOOx0nWiTJOL3JwcIm0opHwFePJIVEjXvQhy
uVZ9FMjCjrNB276QR3MJwXCdWWPVvj7AtfJPI/XxhSgyvG8VDUP0K31h161KP2pjiMHo+iErQ5pm
pwo9/AwQdTFy2JHPnDCiCgzK2p8hxoOw6ghTJS1OTfKWo+NjkVpBrRey/kvvQ6VxOLY1ilm7mwpm
7L0vmOljR62fD5B8TaISGt4ee31L0XZYhqGHtQNcPo0dXbut8sItJtvloLDtFC+lLl8Zc6Drsxgc
g9wANhDywV/PcoVA0PCTpcs/Zvo87A0iihbZaN0v+3aVn/Lk7I2NQPXBr/Xy0pNITgiHF7gLVIo+
DoTf1NOT7vDspGkcDB+9UxCShj9RoFzu/i4BblQ/XtlbeBC2DGsvbym6xS1dyzLVGjYMxqn6gGE0
D6JIkHPtd0vFmlX3mn1clY5UL5k71urQ7zJQhknYXDeEZt8LrYsHEYo10+BR0y3RIDNlKxGH3IXE
uIKorwhwKESC7GApBcKFsUPAc5aFEWaJ+uKPssS16GtHAgKyH2DkUvOCzyJ8NV+vg551yRVlMdNI
AzLv8kLYUP1RBDvN6DwH17DjsAxNgL6r9RP+7sjCy6yT7p4V3gPEu47Y1i2KVKz9wAAQkGaAhgor
a+LoNbBUgNGzBwR7nZ0+Dcp8RmXoe9eb/WD1mKkd2UdKYXfF3v0MGAW3jO/r/fAzn9ZXoZVtd579
E+UHdjQJjVoskG/oIYe4M1RiqUWBkT5asDShd40zEu/ZdZ1gwOkMu/ZbHKnvozSng/P7ROn89jp+
FPMNn1kePuVruptwoy4HIXTS3Rf1NY6EQFUhG3aS7bNjwuuajkb1EnkxVi4dcJr9oZPzxiTJDo4M
IGXCxpuUScmZzPTdgvJqXQklSJr79ugLNYupSqnc+cKKf1MMCJeLiFy7YTirxa8znZbsXbAaO1JL
VQhSQMctwrJ7sOtaoOLuyC9UDtvS8fyeCyISY64Fm+F7/crZkRd3AviN2Ld+/7bYJU4BvL42p9Pn
rlTFRzjjgq/PGfVmlMIxBigAYfe1queDxO2p/6SwWibfeRjsDMXY1H/HS4AbiZaqc+LaTHxuE4Lq
2h4eWNdv00cspUEGQKDv2jxCmvE2NQRoT5T9QecuvVXLYQBkCyS8OHJvLfV1L50wjdxXdrUXaM6K
uG4RMgOF/LshjYu7uoja/EYg386Om7x+Zgu5TF+NGHqnBniT116YcFfmE3lKoOCx3E5wNvUUWcAb
b4nhkBibb4QiASri0lsJw6258YTrTwLfsNpWNcy3skSoEuAVm44CEujJbEDePQkICMtk1WarZ+7A
8Fh6D8G4OdlGL1Ydi8dVAJ7LtOGHPSlsKCueZyLLo93zf63pykY/+nDd5wAKA7vMnH/5gw0SxhXC
gXuxCrg5c4l99IPYcX7Vewf6ILpooEw25xqKVBN08iw5aXAL8SFq+T9C3MklnPdctnptkzMiL3eT
7HxkjlVy+UAh3Vuf5k9G2GFOsrrpk8TzprWgJ+PCDTkWxejbAQ3YqKW60uquZBIX0TaMMGgYgto6
MvLEAUxHfwG3oEVbG36hpLQTgmtEreCUdttzRcn4Sl4N6ig3qtzD+TX4SMx999ts5ujOpH2HAZwG
l9HLb1CjtleQKsvhSaw2vvKyt12siJbz0jfAlVZ+AQyhcHo9aSJnAe/Lkx+xPH3L0gdEo//G9F+a
v+Eo0r5eDfqf0zocB6cqMjoS5eCFIWuNptq6pp02UtfRsvvnh851x2oRdBqPwPR4MxRdPILohXMJ
8ydGmQSTKIiKWAZkOB6/HOBFNBclnbQ+ep+TDZMygUlB8JxeyVzagibaILLXPOu0N3zFE4Cb23Tm
R5D7/cc0PK7S/hcs9IjcSTTpsSgDk3yfnUVqzFYdKa/m/eXKORxyZQq1Y2gcKOXGGQf5pKN/Ztek
97Pk+aNcBeY/e4TQgpFQ7ERl9zqKLUzFwSpwCzqMrGItFVPBMD5rQNKx/5xjhkf2hnz9vZBQbmkn
fsdsyeIe+ZmF3hF9Kafv9LvkZ7/S6Bq4j/yxQcNsr56WJRX2FA56dqKk4kTFOO/RF4qP+dFbiJ0/
foL21hYrfVkaNUpDGp/PHYOlC/wRP44Fb9qsuSoWYZCqQG/1dcOWF3cEKDgpu4QuFX7EDJd5MJWM
xaK2ydz7SKoX28+l2KCSFZzy0AUwJnRUL8422QMUN3aQntLAn5csegBY1NyIUpnbn3fVMncNmm8y
ase3mLWgfUDKU7wdoyg5WDnpLM/Xo6X1OYqAQeK/9oPTyAIBzKx3bsumi8z7bbKyakpK9+7zpZ3L
ahGmGUiIe07AKndfYGOcQKvnm18HKuAsFDg5c19xdNyg5GdCxrNGqOwGSgCZjzLxy2Jd1f2belbF
3pvxLvSJpetmwOKXujz/TCPflNOiEuDzWu5s4LnC2/wuEu5QD+Oij0DtnMJ9VTujdSLNfP3/Dn8Q
yU9ma58fdlLxspZlAuorNhWxfwQ+qLzBInnXFWZgK6drfS/94LEiVWv7jlURV/PcKZJJ/Ht1faA9
y6LoLn1KqNK6qJ1TLQybqPjW/N8pwHkTl2414KD7UIaL5WVKNBbs78s/7GmHlt32VS5+jkL74Blq
NnLNrjy7PrN7PqT1PtxK+jYwO4FnPM6VrZyvQLGbTHOhjU0mpiB9bvJ7cxAMuzXtRShXFyyfPdVy
om+Io5oTJjjdpsKau4YR73pQ4pMES4hNDExU4N42nh+ENXc8+Ps/T1eQvXqURPVaXQgashdjyoNa
PnZ4oq4ufarow1Uc4Re00M9v+mNHGBs+vPsMiR450De70TZVFRQSkWi1XJ1+n/sj2Hsrzp8CUbvt
i0Ea4y2ZIWEtKcoFQKepsvbjjrFTFdravmH9wXwUd2fcbbp3DiIsFaUXWTwFygXgshYMYvyCZwgc
VizogHj5CT1WBK109jY5jEVCQJTikavp0KRCBeUBoDZ9OWtVsc9E0cn0cbvfi7RlEg/SqO7yb734
l5WuhqYBCIjmcJIE7lcBAvm07ZanpZKdWzFtDrCU6jwKNl9URYPRhpSX/Rlq/tqSvyYNyxuA0yy3
dqDLBVJXXHK9Y3vfPDlMreiYLjL4Cajys7D2zyVQ/5hN7DSESImiZ/XWjcC77UgXz88sIOsAUz8i
cFgGNnKubAOySvXe0RIu7BrwH3un3uMtx4H5xRonbKVCnt/7ZFzqe++zntkDrFdu3H2M90NMZMAc
4DkxOZd2SzWt5aRGg++2s+FC57FOJzsQcHDZGNu4Mz4ROqalSRwOdbaVmrqJkV6fF7cIE5wuAoY+
od/xPZbdRNLTuBKnjO47e11F3rnh8XK4KekQHMB+wtEIfTqBC5ASOk1XPw+d6LUdV/bBkud2K72/
QTHJOj/22+ff7g7vDE73spiDs+hf5BcyMZDzmy0ouVmcNRTwTEqmiJW+41ee93cRLkydMkF0wlHE
anFXjYUEJbncwu1U21gDsHLxUMnKz2AAG8Z2+tFx5ab2gW9SEN83W4CC5TeQIlBTOhjHR/I9w/nu
rfEdNdduxeBVVNs7zaWBG9AV5SFt3uZoLrRkl+PECSw3MpWjVCdA4aXpFbeT2B+lfd0Vgck41QdH
irsEy+qLKaFKSjkdDrlZ/NP6PnOvoJuVTbq7csa/jQVcGl+dAke1+ZhCLq0BNjpcKL9H96oc0kVv
DLx6R4wfsAFdRJMQsD1RXdJhYftdQeFFINSENy5FCgHeuid8V0pVMvIkiXsXRMma9bCrVE71GQ8z
OuFdRoAKYGIYKC1ueCEoacOcwKbxESVWlGVEcfp5VtOIaYsCOE+YE19wyGN2vNIi/gO8/eHLhW+6
0D37sTKCZ1wSw2Y7ChFz7eBiJZYjbtcMYJzt4QzS23QFuXdl+LRUNAUzLSGvxYdLrdQDW+GelREe
n/snSF8Lvnu/pLEOYBIf1I2vLCX/zZC6+ib3v6+FMrEVqrJTj6jj+MU4N+dG1TUTd5xeTjbWMRHh
GaTPqyU5qOKEe+MPedrbuIbKN3fD6B9tpMAVCuxtojIz2StHagu2Lqs0/HLTt2zqZpJZ6Qq81pN8
ILnsJUR86PZpIOP5O/fg2zRPV7drvzKa3Hps0gW2VTzy5sKPnvCdIPtMlKaaVHdm0DmbjLU9Isyu
+BKmBcaNqYl7jpLhtjv6xnUQ1Pj59dbUxvITxv2jSS4w9oxfb7ifj6jdChmTu4pIitzChvxYXhUM
I34Rjkg7Q0NhJMTFEB7YO6K4hn8of7f0VcbnrMi2NU7kGFyzdegdhvtpBtyUHWKgaRL0eeW2eT+1
m9A22snAq+USZG37uRqgQOX9Q/phHpFDpEOHp+jM/sOQaozK49tykPBxe2IvM0TZ2o+fq/btEtJD
F+OG77IYRJuxTU0uzfQ1Te4Hno2cCYybaXUUFNpZRuCOncWsLG9AHPpcMmVhN9HLb6Pu7TOjnD53
EQ7jZ8vxA4cGgznwvOKALIO4yxCq9Du0tU1KP5oVuAfk8rbmk1Ftl5c26Ec7aSBRE5owRuCZ9EeE
waQQRijziy+SLyjU1REw/8gKLry7+BtKwnuPXysULpF0hhOh2hp6whzW8OyUobxvDH2/RJ03WbMN
jndHr9GQfTbjTNXlgpxO/iB6gYpRfxZOZz+eQapDQ18BEZwsdsTGn3Hb02p7fIqKiYGczT0aQGst
46GV7swku6nuPupnPT+Yqffs3DV1TWBEM2OECp8N5ZAhRDkTtFPiksjiXmKwA1G94nUGmMR88AHC
XBSz7xpyoQrW4Hk+S1JieTu8BYMvkjmXSVMjz5tiawdWA+MtxJbwlCH5n4lMOMH4oscvdt8GM5Xz
Haj3rxtc04tp3V6+qvqyBU71Ze+ooNBEd7DCJBUqPQJ00np1HId7+KAI2sYjSTnv/uCEfZFbmOjY
WbvmYO8T/lXyAW424kpIT4dhuk16+iUHpMmbzlDL+FC+U0ATYc6hF2viEdtfzZz8HIPOyUhIpq+b
7vBK8rNNcL/SyBngHPslphv4ud+GFaf210dvUUXafyN4SmTE4SOp64KZgvT/z/Wu8ZZMe+r9mc6Y
1pPrgArejfgBtmc6dI3KB7vvwflu9bc3hC1HjoPcPfaYNPZAEUp9Ej9pdUsFD4u6MlXy0ZIruyFz
rGCs2RlrBXsAN6cGvJNyt0mhbKZnKmMfFG1E+JmmniKfe7V0RgUISCHqAFVjrkB1CV9yqssX9sQf
3I+oaqU45xATQSwyaFlAJOgRCo0eLQlZvLFzAioFr70pH4qjNxjyTWAjjUfPjVez2uG5+Qx92zcC
NpqmALbjK4vH/v34C0pvpxTwkjVUsDBtUsuL28EsTfDou6CgZ/GeUFftUtS0+uh7ezA0LE4lNa2A
hwyASQyUBjGl/abBnffxOvcxdHJtp/XLpBu/fxzqWpOFgjJKGfmoBQwnWDAKA8bKXuCn0kbrKqEp
qQpgIKNEgO12ptHpciEWfCxqm08F2dFJwc6ih/aTHJ38ZBRMYamZ5+OG8vw2wuVMa60Lzo+YmEo9
Fw14g22qhzWEAwVBgo1K/DTLDnWDlETOveg+iQnOGyRu7gGysf2bnXupM/R3E/qwI3P5IaNynDnE
46h5yNzzZfeuE2VH2DNTaHZ2n8G5s416hacKG9JCPRnPMEV8d6KM87Wf5VcpiYQ/79l2AepLrbAF
/6Z0aj6p1SezLinnH9+Bf+NztGoVTks37FZSxyCqM5hTKWh4EJeESqSm/QgZaA7rQSw6ydX4eoU6
4j+ZZmqACy5PJcPuc5Aq6UN0+E3aFazGJSukFA2Aghhx4j5tGFOZOt+3vkTJ7IkrGHDlJMm86IJq
5d+HKDvKIb1xvsMupDMhJQs+gVbCxhLkKrakUG4AIdXW1oKqgy9XHeewyRgkyDGAiSHJ3YupskWm
GuSN5IT9InCeMHa2GDxqX9DWBvfTRBul9++w5cgxNiRj97FrmP1ZbU+hLU4nOh5h3JIJ61TCityh
bnLkmfuJSWk9OB6uLbsKKx89+mO/RF7OOyRiLHAmopZEuJ5lerIzMmpYFb/CvUklltD6VNpqwnxI
QgGuhIyioiDQkWYrgyd+UDRIx/RaV6MoE0GhRshIczNMLAiJPruxTPsn4cDoCpfKoHb4cllAXP8o
3yruNktOH//bZzly6TRDGCmOgOwYnCwNvSIF4CaXXsSkimGfjsOER/DyiIX9dX0EhB7CSLjnhrsO
ZAU+V5QyqC+tl0wjpDP+eAAobrLmYn0s5eScuFtN18t3Pz4zaTipcsLdNUB+7mN5rGwvk3W8CS7r
EI00VRcFxMqkfgT59XtgMEh1rW+ZGmVB9SE9IuC+Q10cB//459/Y5iZPvgTT9KMb/20khpChfPFT
mB6S9LWNYZGaC/Y8ampdjRekBOEh6gFS473lWOpIz5D3pxPEApGJd6yU4esYub+LtY1qXLdDFSK8
EYjJRHnKmQg3PBH+gmaMRItGCAoPDVE8V0id11ouaBEpVBgCknchPaKZizVeTGFtRyYERygKRfKd
9G6Wdsy4wpIICVQyqvQQ0nmWONyWO5Fj+IB9BcA7wAIJOnLNr4AM3h/NoocKyHROwIXhexYRNvtA
eoCC01EhGUzirspyGjjXNuwUYvtAObR8SQHw+ww5jNdH84cxpUh75T4fsxgPg/mg6dmdb/OBGS3b
A2sbbw8LZVkgyP7SWwVKtXpClsDLIP5jI0kro4ffbWtk3oUTepvDkaNTHR7KStJfBWLW5xAu7DGS
GlY3mqwBE/sJ7WmbJuZr8wu5hS5mZFNNbwHBOK443r/ew2ZJ9t/Z16Q1t3NWlTa2GhAqb/kzeh2P
++V3D5MDyHVqlXb5fao/Nsr+un70M2wNtOgErJX/ApbzHdrAhdNI2MzbQqoAtwkW6dm/bwcAyAiQ
HpTz02MR17zCBrlLfm11FWWumaQjRS4hEhEs8Y5ipWBE6XoYv/oEpr5VhSasAI3sPUAm3EVAxDCR
7V1142yC69GQMEemCtDup7bBgqFLPv8szGUSRV4WVz8Li32TdT9EAJL3bJE+raBJLWGNDNeSLR1q
Zxc1eciCyDZmqJ92QBojDnt7XB+219z9n+7si0SUdhUNWNMP78sW1P67qYN5v+yaNSaxTuw6F4YF
u6uMv5Zl6beAn7EM8iPl4WiqLbXFQCwIYfwEetB+d0bGHttEvhnx596a4AvkkxtaCD0qqcPs/xV7
msP3EdIfOW7FKx9U5zt+1L3/cwKF2zLsjd5bAblTJSnYjj7vPOfr/P1o2cq2D85T3dCU45gANwGR
F7O7Ge4UicbywCXGrTIswM6ldmhVJuHMi6wsZbR7PZarbNnbXHr2oWCeMRLLM1y2njlSfAmO4tiP
lnWkiN8Z/JXqliesG3Ab+jtwLXPl6Hj78igks4kCSWEYKOSLCAOTl3S5KrIPgEVACyjJu4i46yzx
ESYFU2XIpBxqezpHICnlke3arrCGf0Z1XhwwAlSPleecxajyFljiY49PphaWbMlh56xg9xnGF41E
Z/TLpr4ZcPdVSBvUiu3I8pPq42DWhw7371DXU7aUtp59n17X9HGDn0nClWpFduSYRObwqzI5wihz
4xzpzvG+wSYzN2RnNLThSURnlKR9q3uvNGFQjevkr0nV4RjFA91ZDv9eqbdz6HFt8kKW2d1W72iq
32/S2qEs0qOYQOWdRfXWo2kEinCyIILFX2I/liiAT1cqRq0MPoq9VJf84psMRBG/EwMQH8aUiNc+
cpIlnMPNBjMUGdUMhTwVLRjzCQUdq94KboKnMbEERpgCUPtOUsRnHrSY6XpWPFNIOzE7NDPkcFtS
zk6HEGKbivFJ6pwzGrc7lvdImS20VzVHHceeJDxkJd7x5VWxXuurun2V8po4GIZUHDL7sxNZCLQE
3nqREvF2xh+Vtn3BQiid8Q7I91BlHHMsyZFXmqwFXbSlSu3Gdq7wZKxDJ+ywAQ0bc9ANMwi4T/hj
rLg2+kJcHS00XbSCQZf2evY9ZnwKaYXQ0xPhEY29vHo9Tm5AMcf56y+OX3q0+ua4QWWcXFHs77hy
2vEl6yAKaaRZCbLbiHg8215/zg1hnmpVYfMOSy4K6Vh87GeNBMDE/RvVZD+LqfBIHLNd+LZVchuf
mp0RkmJSB1fadtmv5Bw+j29bmtLk/j70W/r5RtCPs0XY/scg8v/+v6BCjXkB24d1CC1MnVrVOvbo
87osvyycQgJ+lGqI2NIMyis63mmLjgVi7+1QeRySKQ5wZgb7iREPjaGjN3Huaf3zWzX8sLuZek9Q
cg4SLM5OHPhKub+CgQATATh56rmLWLAu/1aknbMS5/YsJCjAIwaP7ZEF05Dm2JsoDfLgIDC+vhqh
HfEIZ4Jyd2nQMyNst1172GN49RQRBbX1b4Jmqg32tu/ON8yofiogzAtnEoIaBp8Rv5uy/uT98u/5
p/7vdZb/yTustRB3x3sfN8KtLbaqXJwo4PMgdVpe9ZmFtwal1Dadea+AqT8reDi9S+bNCmIopj9G
/c+e3XmPaSPUUIKXW3uHmMvCWwyzM9BG5Ec62qhwIhCHzbQXLIpFXjz9FMvKljuHtp4O9ie1d/pK
PrdghYr8eFadJ68B0VrsOx6Q5EQ7DzJP4zXAu0xY6QwQU0Snx7fIEeadD0AM+i9wWAE/hyTJuGFy
OP5MiDJ3fS3lcUmEDQZ/kHMZnVAxcIFUZTAAI5XphROnyLD0EDstqPfHicKIMAdz9bmc+rTAsLO/
h5DFiRI3YUEGqotkYjRzHocHkzfF5z6X0rDk5HFCfzV3PnHm2kB3ZPT2bjnYMO7G9VkS3INOUohV
G88gfe1m1MMU8pM9wWfhV4y4CsqBhO78iBILTQrawJTpYnQTb9NxCRsAVixJJuuv7BE3DAs+QqeA
bNM2G/tbyTT7FTJd2ZKW62UUSfmLMARSUlbaFttPwYojV4BF+XJpyO/OEvRAe9BjdPF3zgjnmKNt
p6PptUqSwLDkMCmLgLWK1HXYqvzGSJ+VwL6yy9ohuR5vqj83enGCQJyWDwm3JxNc0Wo7Ckso1/W1
2qOPuplwg+Br5Y90OApMV5KUmdbeeKKc4GcWW47ldT+ziQjEQgbwbBXSWyo6mi0vUNP1JSffifnM
Ex0F5dicUEjgBUVVVsLifig3X6+NSgVYFgMLwxvExNmPLAJEV4lThcM2TU91uMKA97Jb56MMM/u+
xd0HdNh56gEsoGzLWOhdAhdE/6nLjdEf/3eSUZkIY/HpoKJGlI4IhfGiVJCmIRcKoafkV0gB9TW0
ksXOrl1Z984mL7jDj/ul17R1uL8U77OMVkHZnAGdZCrairF4/J4yDDysXu27Cti9xpGkDnK6WI0w
ISE16XkvN0Ddu2q+yA6dvqypM5tuywQGwOMbXokIkWYkpK70CWI/zBigCfTWWj6Z1f08gnBS4xlO
/MbELxWM4Cw1vXCG8TSjEemxvNBO+yONFuEf4e1QUG34VzTID6Nupe7GjGbsUnqvBf+pUE1Zdoo2
rEuMXTQFcvhdvXn5ugBxn4f3MZ3q1NQgSOmhHzb6eLHVXzmB+NcDd3DC4ekkJfk5zRbC0k24eRzU
l6t4zqCKfkuS555ZtsATYy1LQgVz3eEoaBmpFP7Z4BQyxUAHlBYLXf6s7dO9sP40Nr3XKdUebTQ+
yE/bNgLliHZ7BcZAf/PpzteZ4cPQdYTRIWaP0iH3WxaSPOP8TYI7BDs24VSSEGG4Z4KPJT6zqePE
31W7joSFxeBwWjDToR5NiV7Db0WL0JOc0MbESK2yl0ou1Yz8H0NudWQcytw7uV4lywXK34T5+hHn
jK4jqnIvtZdHmJhnhOJn1j3GMAn4L8ya4rT9D8UljDThQyxCHCex0UWFA/Zo1GUyDXmGLl1OIUWJ
xmKSFs1v2Q9mwfbSrR7JYw+mY9OeLVhjeJpC0I588S/HN87F0NI4s7GodTe3Skc98KahaekXnskp
g7YzB3vnnSHX0bdRxYO0oI2OsVYuZYWz3YAaF1EpvFzQVFVqQqzDKmYr8kITrC4tzr/GM4CDRPue
e7ZR0RFL0WJl8+247ioJ2uDQmdxl9H3haD92k3JIWUvqDQ+4LvG3Q5IxSGyDFGkU5SVKkcEIs9Fx
v+G6pZCIUf+Fzh78Z1ex6Yk1XtNIUD3lkgQCJ4Az5OKGsgof+d43VtBtgG6x6xt2e43XTtBodP44
n4v82e5TUpnVXu2SG9Kggm5Gomp5UjQgB7HDvTgX692/YRPXYP8q8/UEHjVygEgNeDgQ9zidKGCr
sTGZaHvsOYpoidWWHBf7F92QfehTacHg+vhx2RfgsPU/m2QNZEFRo2RaFi7MUG3iZqyYsSwW3Mgf
Wb9P1dW/S3Z+W/nFgk5X//KojmUehvT6mHX7JAjwhzr/GHspuUqbeDQCctbX/ugCzALtB+wYxMGm
JN21LlewhzbJnYnSiIan9M95JTQ2OE74W3xcW6wqQ8C91tJeww/Uoo4JjbSlWpEzg0cemOwZUdB5
GjWdVmtKCblxgglufoIpnrQwqp71HIm+2dEqrTWBFDXBBmRT5lOh1au12g8RdbILPPeXVlpx5oWl
qQKXp9NpQhbXHP6BGkHvEVAPxvMRBgQfzHHqNSRUafii31Na6bf2Ytxgvn55mzPSF93P7ca3wSUr
yXRkCvrxB/tWxn4PfV3Am0DQ/2Kh9hSa30V/KbX4F0sxE6i7p9CWY6gMQ5CuQyg/nk6s5nBpRIOK
gNclXhCFqWspzKvc2hveQf6t5F0aCXNOZsGW9a6yORL4ejLH5M1AFoqJSfOB+Q186wyKJ54UvOyD
LJJTKzozxD6xm6+bUveJ59Grjb/vy0R2jH4KdtSTseNDRVrMFBvWj6+juaNHv0jSJRs3MR9w4lah
KzE8qO6sxEGyqYkVBM6hAkGg7chj+iX8uUgCXruUw9UbSmATBf/RxmBznSR9cTa2Czx5XumkLPto
kkoc/c9xosIGU2pKYBA9hCq3ssI3AYGQvBi87n4HS4QdW7fWJwWNFQBIY2SxJJdAy5fqRUb+J901
sJ093eh89QuEirZMgABUQELM80TBh1Vl3LKqP0/3fvzMF0f76bPs98ZPvJvnK9znLxIR4my0mAon
z8OERif25YImThm88dmEQ/xIKq0iKERbFrtUGScyQKx9NrDI3hFIuzyVcsuFlQ858vd2hHmNS6f0
Q2fp6PIkz2LnKGPfnDdMte4hyv6q6htuzWraNWE2ZSBxqur9Qsf3d4eJbTCuHXm/vRs3DoLSMhIG
77VrQPFprVJQdw/5d1JURwx5SXF165JBVr+DJv4iUhaonV3pLcezKZVcMuqWZjZDWHyhsmdei64n
XIrE6G0w/e1EUcFna+nrzsz8MOeDeRcHsqIxJYcJ65k4wOZhFkD2+yRQLkvI/oJw3y05Wl6cWkyG
ssP2ONh+g+gOetxVetQE3fEN/+4Wb3xfqbO3+bhpTJGGf/sTkQ6wWyNfUkN+mxS8sl7Z0flL+nBp
zKBZznDCCy53A4iJIhMUjrPZAHGFSXUvCYqfIJaeUyQcilTs5Br4jG5xSDnjSyHuZzIhcJN+XSQn
UxRTrOkXci9h4MwEgkMEQeDtGcn6taRg1Nr7KGHdMgpjI9k8Ke5deudl9M59wBCTXyrjlDCTGkSt
rVAdJsKY49hrxY4nv81vNs3elG5rkmfTovXw+Kgmkl3k+hWjrApXI1hEQxHDem/+iy7UKKXOSSi/
Y4XFzKpgy4z2oTF0V73vjGdGH/JT8KrE26PpvUvHEk1AnM81Ca66zTDRyFef5eOn8FvzBgY0XKZO
XKVO8AwArbqndz1ca+TI1l8uk8hHQwH4su6BFp+ufEq0K51I2rzaENsJDU6SaaS6n8rx7xzQHpgZ
2ckV/bsfInwe54VqRuZ/0xUOdztK11hvZdGDf0eTmyWWRPVabvBMis7ofh2RRP+mSUK7m2OqPSim
cAgVm1F2rkWtKa+ilVGgcxYjTc/09yQ1+vkq/7BgXBqagUCA81BDUmu/tzk5m8BAKj62QXXidp/t
DjrHjPazqo2SvK1fSKg5fERv4Bmv1o7BnQ69UYjh36sI3MXNHUW5axwELXmkBNgoFXzr9kW6WYcr
4dBJ5AyMUZ6V9FSYW7Wncpwtct9Bd6kV/Q3aVu/6BJILBfHHb7/HDmjcfDLpUwmeEk2UmLgU0rlk
b1Kcelmv6BpQfvh0IzPG0WGrZ5LrSJSQi4g+3M+BSYhwimID0rMLE7aKLurS2N/r6ztlmQ3A1K8x
lUM3vJe82lsXFTVfNaxYrq062RvaxoXMjYXrcug1dxhZFoMDAWC0PxG9AizId6sGUc/ewAVHpdB/
tyhnL58hig+EwhGthBlPrEK9Oggd69RCz15n5Mf2PObYrZ8rW0mVOza52Y4KUzkZelotS0AEIaCi
P7sy6YnGEwHTiMNxJfHEe7z+caH9UJDRKe6eZxl/rtHtDybZvSncqv+Qpy4mlyOhx/G43lhyB/zV
yZqUUlncUemqI8IVJMCEQiRt3EEeBSB5fTN9UWmqRXbY70ALBensNXHTtwzpZngt/HsR7uiu3HRK
FXCuE9D8TsCZuMLaNsiKF50xgiYP3tW6iy/p5djpiCoGyt3poxj705RL8LgMUIUSx7HiYBY54R/D
appknJqJJFk2Md3FVAokRg+hgSZEH3BcuLF37f186+OkkozW88Fni8dW8aBY+RPDV6xh78Bp1u3A
hXiYwXyNrFOq8+0/MzfZiaAvymj9pw/O712kbrMwzppWbxwz/XS29leGHRlRf81BVu3UJ5fY3PH3
jlHSZzpOrG68i9Bd6b/uHQ5haXIO6SCN0ONVZAur/VTzjViiSHq7UM1TsSqgwJybNRszMzs4uHol
X1dmnjF7YfkSVhVJZ1+PuJI5p7f4nuSJPUWE3rLBBK6COp9IjD1SoK0mSAeK2i+M3goKw9o+vbJ1
Vh0aHoaNtwjY+rAi25qRRYijoOM8q9zzER10rBzvMfZlNQ4zbZT/u3FwuaumedsQHMBrMOOOITKb
+SbpoFdnFPeVav2NTX8nKUhpkU0+8D/9XXVB18vGmu3gej3HY8Ra8uhgKXJsNFv7ap8SQ2b+Ezux
dRvpoqBtSxPp1Y9fCHOCD5mB4ZIgfbs2Zn0Z0oi27o0LzDcLUKDED/8dte8fImbSTILqM33jWo5O
HjpdhYTMZhsAZCQ6q8xDjmcwi25GMFvlKoOaJzWIb2PgJT3Lw+H/0U1OgcbMQ+PCt4IFW5BWmkmk
0MUWCiMf897crVP4ZLLwJae/QfIQKnL8ox6NYeIBVu/LHKGD1SlKME9RtdUOgFDaTAADvotjHWQd
X7VScaajBiK6AVLMgqgAI6rO0ODe0CoBnC3gJLrcD++I7ollf+1guWXLr/FyEmbnuJlmYUibeNJD
Wbgq9ulfSjxIAY22rJSi2heN7bVnx31KyM0NfbHnnUgb72E0I/FkDr06JI8XwIcqLVIjJFLhqXWy
Oc+fMxhQ1MuG0eo+uuG1xcygXk8CdXZc1ku5zBWNc0XH5NLNnOpiWU2YkMJm+GcKIEU6H+gErWA2
Nw9d/TYDiKU5Knvjs3l8BtetzLzxsbfTKTtJgzUSHOuJ/8i3TUGC0OiJH/8Ytt4z4oaHVe062q0m
ENTTCWKDxocxNIfI9AczZrn60hpQ6zi8C9HMFMZ8+LLpxxLRNuVSfpTflRObgrZQy3z1WU5KaXE/
HaQmjoXcWXJuYoAy/3RZ9KZ6xAjmrYfKoXZkRZeTk7RXtZ41zijrqOXjyGJ1NtUMuqzS0BOkRNYs
CWpuei1GGE70CqVAaHJMM1lNfKeMZR7ptGowK6ploW19gqcMfU0de75kenh6SNThCirebY6RJlTf
d1xPsCXmAKvwoK8wjpjHA4TftQ7p8agiViUKhjLJXZjYdQxlnGswDc6c7cTBIpRqaSak1R2PQQmI
vzn+XG3SubS+ZPzbY1/Eh0omFiANK5d+8iNgQgM6qiUIVz/fyTwdvgaQms7rmgstTi1n9hRSOYiG
f3HnIrkAklHAAMgGzDsnZeCrdIk2KD2r9RhqAvUNOdHlBJTwUpsKHYR3u86qFCFdK84zFHsf6oAq
S5kYdUvAvnPPvxZpgtwbUy0sfkq8OVQmwHUegSd8t8i443Jd8lK702SeDHPwz6ZC+LYJtvxOcj7F
QCNpkjmkRLKHw7KK3QpI1BNYbg/tlJTyLyb8lNiVBy4fTsn0fUSsGCUCHc57dwwk99dynm7ICTe+
mAuiIQM6jjw+3QUO/uc3+I+VjsPP9b+XjaVUjRJXNog2NBof21tHYTNoAPBcNrcnIkk6KzfOkIDp
8/JJS3ZnQxLhqY4nRyKiLin93Q6QXd5bOraspRvtY9PqgEJmYRkN9MrLIq6xGrdwlYs5EWK0IEPZ
eHHc80b6owkIjoMvemSVC7OaeLJdLu7PX0FTNoZsm7OoZOdTRK8iNcm1FS6R82vee2cqaK/jP5O1
sSF5i/JM70Zsf2L4OGtXMA0MiStlN5yQgQMBKaLCJjauHKZxNpX4ENZKG2n+I6nx84uTN21APxt8
ca6tO9IdKxWzFitBJ0COi5kzkM2gj34d1Pz+5CmvxoSA6LS2gfs0PyKfiaXBoAASJR2Z+TK4HKvd
oZ0rXxGlLIndkU+BYNZzCFFOQd0+l4uhCzk2ZF4RC/fWjUwSW/eJ9Esb3s6sCd+3L/Ngijsl53WK
eZx0UVzkYQHTsvlPZm1WB3LTCj4JvcnNIhY6A30v2yXBIVG5JWDDBHfNMf7lUGVewAvazuh2bj1s
OETzdy57cFdoQBuAl39MA2apu2TATp1XC/ptSsuEEZqzAORdF6HKQ5HwqCObV5/q6iNHqt0BfX2J
YaKlnoK2RJLVhxFs/c2ePgXBNOQpJb3Gm8NfcqjAhYR250nPGJzTouSObK3hsZe0hD+vXonaHQSl
wHd5QJFwGzfd8s0IgVMNot9nP6zuQ22WKDFI/j40b2NDSQZnQfLqHuLEPX06/ifN2FdCoyy6lTMm
2YHF3L29sVzKzX5cTLL5KmuDvF2cucxnnlZekPRlBoQalV+hFzIqZwDIrlhnsGyXQhpTid38Vn5D
6Yt3n8TJ1F7GiN/aD9D6aophUO8b2M6qED57TUaamSpot+wds2iLMd7orOcZgKYeZIJA8WC4Gmgw
XzDhFO+eWHF4fpCN27VzKMNIDMjnTY6dBTArdz4Hyt+Ap5ZLiKkwX+/u++EG6p/WJRrupDshDrhf
ZUZGBU3660IDX8yszAn3NFXc2MyRNyCKJFrnzc/nfKWXPpZDP6oAvJWzSuvt0ssZK+PoG/63qOzZ
fI/jFUXhx9ArH4uS8Tkdq7aHIL7CEhc+uisFB95QZCGumJWP5VNztFCvN21KXb1CFihAIxwWAhIL
61fQ8pmMLuYbx9RMbiX8aZJYk+ASsnorq2rfC9/TBO1ktyNAad06DNVnPcIsJhVJHBwSeve60/ey
ilHtpn/1al9NIgJPJUwZIemSjzXdMxDdapD0EOMhiPtJ/rgn2+lk7T7ZiCdzDJv+r8hjllL6YXe6
eApuRmc9QLACQEPN9QrpL9gshdubs6JZSU5ecmK1rR+TXhE7kTXA0OOsMhBHJ+00kmFkby4Ngnag
Yyq1z90oxZJqhGU/2YM2/4lPeIkvyPGGdLOv5lGYc/xQY68V22BOmrrYtALJUEPlejhStsMPSSXs
PNEnsAY5+edR7ZbKxvn5/9gs7XMB3yQlllqiLyNknudz74Pk4Z/OgY+eE6MPy1GJ73aIYwzZi0aL
K8Vh+eYGPN2SZO9Cz30oexdZzIrPfClgXWwiVVXFwipxunKdDkvu6kqn5Z+Qsb0GlAZF79QSpFVC
hHU3r3pZEpPrZ96wpg+G4TbbEHaxKrvwbcI+dZpN0y3m3y/G5zoMqVRJLsWy5WMCsg77TeFfCYb7
fLM88dt8JEzZ55Y9xfmW/q0HMeW1PWZH7UDEDPfuGd+D0lBVLm6Nuxxf+nzFdnA6L4KcBUCUChs7
5VLnxzpTyTSdQpd0nYmv4C5ZpfMLDMGO8vLFPrVnEdo/GQG3pMmF1VgeSgZaqUfvwYFm9em+Gfsw
LKSI+MOe9KI8kLHzdSpVN2h9ZQ00Pjjst6T513+DJjYVa2IAI0oZY1lSVgblwjnMWHKeKVdUfdCB
L5r2Q42vy6fsMMA3TZ9wFy1F3SV8P7pJ0wWFT8EHRgU4QSAvxggkkeKUB1P0digPbGCqttM3/MaS
W6fSw3AlMZ6XnXKtAEcfWrKtwOf2f9kCV67X3SCj8i2O4n96C2l9MG7SHgkjhXPX5y6kEDfpiDm0
sV37kWxzX2hRQclQCsSrdMpP34Wi2nFuvl9sx2odNHJD5VOhVz/FXhxc9btOIu9LzPLNS8cGnhZ0
UEO5oyhnLF2z+Zg3nkLmiEw05O68daym1i5OklW+YuFSG9O6wJGkhLloLl27TYpCXjKqlOh/y9Xp
2yMJONOyROzB4Y0d+5RjRI0+veP3dOqau1GnsMHAQR2uVXWOzrdqtrnkHbtvZMCnb5ZfwDwI1bbJ
gCT4iAxds9qFFci9OU2ZZDNPwxObjixxoltLiYGqAVFzHah+lC1nrbJdYg9GGaeNny9YuYvVu7le
bLmz6689Qdn8bmvTcLyAp5F/5GtxeiUWVDDy2WUBuApYPz0mwtPMov0qX38i2JJg8rnKuHQXutf4
aDD3nNZ8IT7Y/UgsspgZyjiO0XFT553LX67pckNmNvCNMlWh5rED/Ty+6P/Ken0zCivmlCLvs8oa
AR0NjQ098OB2aNi/4qJepYwQUSQ7+5oXwBenArXqGTF1uCTVK99+Ej2eDLdtXheTKF6Bj5IdSjOU
6b8RjyjzxNNs7BYcQm5rXAlliltpouwYSo0XkJWD+PqjfheNbH4f3qwdu0TLcZ9+tRADd3aqp9sB
jADflf5acMyIESt6ycN6NrHkbnT78KVKghdA1AAVxlYQRMhzxZDyRt/AnbkwY5SXo/RoFOrnK4T5
VMB6oTBX8L+AKET5X9Gmdihb+NPAPtCzp8XbxEU0GNZpXNAw/VlYGO3QI/lBQQD5+fMtrCS8b9vP
Rijc4FKAs4Hgfa2Hfef4FIGzZPTCC94H9HtSkdnmYQKLxYDNXOE1J444PMsA9rYrTngSM1KsYGL2
s//rHMJzVm5xrLRlnEmsiIJAUB0CqczMopTE+nbmW56sIU1EUjY45W88HaKXThIAS8Tse/wUA6Uh
yzlAmEOZJ97oStQQKNjkyYZb7ljyVNHMoIbomD0ESKxxBONhyGGqy+/mby70YaYXs42Z3HCL1im2
+SafTP35lrXKBXlF6h96llma8Y8lZAfCd7su/AJ/5aYMaAQpuCBVfoKWSUvSajmSSWgAKgKGn+8J
YZoVB+cscpitr6fgsF+zl/FRWqCz5JDmaD8jEl2+7pe1LojATZ1KY9Zaxd15m5Ymwmk5Lk5CjRgu
2PCKItlA1vyy+A5TydDxpHQOqE+fGWqvBzTYJMSZL6vAsEaf+XP1JZnOPi5JVhkz6QWl8uNEFo1P
IYkkSt6ZshanFAEkDkLuBMdmXfeGavQ8iewgZaOaRnRgauJypppzjL+vFa5kOLHXJ18SFIMKTmuj
DABaQSsfDhWCBYVtKyeHSp15mf3UxNYR7sUb+BcwXD4MFzRDk4U4f/8rdY/V6q7LFwawIrRkFIsj
0EInG3NRwqRykJuBGeMvI5Q0NAmTNH7Er39Gwj99dbE5jjGlXSWn0tV4etaomBb0ITqzCYEuGxI5
MVM/RBnhBOKlVx7rOKiBiETAErFViQ6hZoNe1XXrwXspRDb3QFJhLJj/aBTQiuIe4La3DweiQ52Y
8ZcRVy56+S/DpJcxL2YJOJclSBBHZeG7Y+CaZ2CmLcJ7DLrmYSRSZVXbZagIeixGla07ppwSodyg
G0uVyJoppJh1QrpFWldf7GQMGP5yRO2d+wkCX9rfS5nRXpANCATC8H0eLB7lDPTAIbaft8y2ts/r
ko5ToIyYyX5NqNri6wTsDtaheyMxGbRmXDfKh0nvVRIElmLiHvvKtQrksZUvwoa4uwv/caDokIFR
nLPeAKXlK/RgfPLhx0Rb+btKjyHuLX5x1XM5XfAB8ScHDfDqCClBj/3MLIl2IiqiWZoj5FjpZD7N
rGiUFuzcIavbpsWlxgqwaQOO+6PJWM13Y801CwtwvS4ewDbWnkD7MFqQyg2H2XiQF3cHX4HmZyTX
6ioEXZP09DfkRpxFUfZ8jMnS3CCzxAHgkuC1lXVQunnl9nET3s14eOov//qXOor86zvKA7ZJ8Eur
Ujoi0nvTFNAzL7xi54H7nQR0NuS04iYVFcIM3Zpam6w876FYl99rVexDDEoYLCWz6NG4sDKvoTFW
2Ff5S2c4lFgx7Bvd1RRXw2kVyZ0+1rksaW/4vrUf5ve9UJrHXa3nCzeume5fPTNUkB31DICqWdS7
rRcm4PA6HuvVJ/Bn20pOUnF8bb5DlhXPr1fS/3x8QWNSjVzrB1gvX0oZUKTLz5AXKH62xyBSbSVj
3SmRbve4cHZzHEamVfLZF4tKXSttNvA0YAyL6bliwKW/5csZMqTeIVjHlZdsEmCdbwkWI3b9Mz6F
eH23BrEp7qpcV25Cmvl0TXGPn5KhPPXmIVYCGFMiPvDxWur7naRSrriXpKSOje9GV26COHO5j425
6sVLfWz/Jr6qzUUZeGPsYqfnha1/lvRZ+UcIKzZsDmn3/l1v+g6QMTKxW/L6zTtTeHGNzfR0GH9M
ILEQG/ID4YuFxVKdXFL7aBk2NvQU7ZYLHrgZmoUC1yDTYlXFQ6AVFgsWJa+UEzP1ehqJQv2FjnsE
tYc0aXcRNYBgeC098MxN2KUnnsyeEhMPed347Q5GT3zDtDsv/laWSVNxyi4qTWPQSnKJuyNCacpr
uCL86ICmMzXUfO7rSq9daFruJ59waUKFQluC/sTipJ24brzH+WgFbQ3Nuk7PVdVBqTng9TuKNlun
meUEP5Ld2Vamf38Rev0Ta+HTjinVmgZUMtdcgHkuFQ4wTjPMC4oJE42upQfX7uXPceK/6+WeVxZ5
fBAehsX2l95Cbpy5IcAhpc8DKbCGbxNDPVwlwfb8RGn4sKZ0+b274aZ4pqoW3ejGdr+KbzONoNXF
4ihL1lHb3GBMl9hz813Zan6/ZUQhx7qTHf09qm/vyyEFLtb8vYpNhqLtpiNYpnUetixJ/eJapWAZ
rYPImHTXbfGYDNDBd3VrCsoaOGw8KNiQZvChXnJf3fpQbfPFMhZMSgVIWOe6dIw6BEzp9Uv1JS9F
HBV/bwpgebNtQlpNKHc7o3NPbnZBJLi71BUjmSTTABK6YcqgNcI+dJuYL6v+Myphy1gM3vD9al0c
3nzJ/ldC7ScT+RobKe4hwh3JyNoD/FQg7HHN9HIipaFyLuSp0/QKBLMuSZJHYPCYfcrAaQ7h5a9R
t77y/d9w3b24NzZfsf0Fhb39FDzqCynjJVMkjiJYB8VPgFZGgw5TuDlr4+eNpr0Gb81RFwP/KoUt
BU56v/erdFP2QY/46FNb9ABFq3OP8xfcXYBTzKl3X3cO1rKcxn8CoCBDSGAUFM3vbvvQAzN218xv
ihp67GKSH/lwOF8MBeffecBfXAT/FamoSrvoMw12ra7xaKAbywvKnZBEFKZq0Lgu64s1jBITKwki
+t810Xi9GClnsbsxfZLIXKl+b3S/HGnb34F7UHhxOJ1VYT+XSYnTZ5Ox00/NmmJzgm3/mzz3Hl7q
DXhcQbUtAGBswow6hrOYZc2+VdviKUemuXsCr5JCm7dJXaoIc2+Tt0rJra6n3Qy/HI5z6Lk+je5G
DL9OuZr+k6xgukIguaJTmC+vbOBj76d0j/6IMs2GgcU+A/uWu3hjwctTsujXDzKGiCBT8n+M7rxp
t553kUoP/c5QyZuRbIh3QOdDykakaqv3FNe19ctbpSXVQJHWqpxk5UP5j2rYwnjf1ORjZ3B6g9Mu
koKM4AZ+HTb08pijtCH2nvCL+27u6wkWPxvT20xZPQc6XpceyentZZ6PjW/XWbUbP6UHYZb+pV4X
AYpk4GydaZEcn1l0yd42mdWXRn4Y8UQqjb065Pl30QLQR8DniLaMB41ESCfknrqq1YwIgtB5l42t
t3lEAoszeDWsz9XL4MTEU+OXlpBe37j0PUpCFn6BDPFAnZfVP9Mv+x8uKV0aN5rl9gPANnPsL+8o
5ofKK3JRpzuycTdP7z8ASkkiXepuo2idBAY31wBsga42jp+oaKVJlkFgmmQTZXiyAUBslyLvKhdG
zYFgTX2ygXXDXsCs53FIPoIgGX529jA5sqkGRNO6rLaqJ5QTs4LH1W0UGIdKlNpdaM5rqfrmsMDT
daeM6ycihuu26u4krKLQLcFVcfT7MzmIleCcdi0kKQUdpnQRwePZYEPaK6BqxRn8BPAVkqrBeT2y
qKvMhycXn6SnsvrTIBhPgqP7flz4RJG6x1zItfixM2NbWbYg3McCWJKX+PS2sHq8Ol2C4+LWYVWO
fPEVjZQNwYURD4Qqy1AjUyZI9MKIwR1ObdPAXoETIRC9WOK38LSfBjAh4Cv6P4RlvIvltpEKZSqX
FmmnQ/nPsoQQWybpoJozEJcse0n3WOSgdE+NJSnJbzNfZLk5VetyiE256kmtZDe0XTWBK1+1rNQI
KNf64EWvQH3uxaeneC0VGP1Q3LZkydLBIkUyFjtX1g4l2wVncatN4WMeC1Xp9ryO/lWAxwkM71j1
X7Ine8TZ9sXZ507WApQIOQ3fJkJZcr5YhynbiOzkyUds6qY0HJ0ogZ3EGL4/vBi7kD3gTEXkOK1D
j4ZmPAGm1Uze7uzqWsWZ7GN02WJNRRYfOWaxFfKn8vGCBxxf+NtxJdmRdhNzabDTQ+lmUizoQFCb
NgXEZ7Ceev2JRs2RHSHf6IEWxopLVXFZVmIVt8GpkGSfotOHmSQfRvpY1VLSIW9H+DbfLxMLHWmB
Qi0jjy5mrOsR8Z6oX8Qw1x76t1I0oZK76Lklqs1aTqHTPrwcgmvkxq5zch1Huz7YaTRCupE6HPuV
XmoWi5/eDIEV9TTAfxByUsuX7Ip+K9hVJ3Eb5bRKzFK8E4kBeTKCNDtAmvY2vmtenHwTisBckv/T
WdehTJXP/sLJTwv+xnZBF6+0OMliJY6ej6WJ+SMy1gcqgtIFQBXA6revT13+6rJq3uzgxkr/xAFA
oIoI+tAoYvSakFqknR3w1qcQ28fPidoSvVyfOs5Y0GpuBujMKu6wQSQUeupA9gWxrqixW+cDRGii
XQ7VpmQunXPjd5zaWSOqTmJeMTMW+ZmDe6oMgTAjSPYc/hF0K42MBuqEgHNAI6fjX7boTuvXlQNb
yT841MZ6gEXTg1pvIKN27erwvDigN43lel7q8gacy0geehZdSjQK3TYt3JaxQensM6XHo1HkXeHY
XQr5T27jXS35nHD/IR+iWSNgid04+3XpAI6WPk4of1YnBskKU2Pu4vUKtf1ncoLZk9DxXIML3tvK
axmFpvtYFH5gUkhHNjTLn/XHGqdnRI1eZ95WX27dqsAeDd8nVio7T/1tVcXX3WI2BLce1CjbSv6O
niqzWf+XCZ0NyZMeNXibiiKXiSJwoesWT1FHEVIilTdGVpkhOsfuqOprC8fWCY2GSuXjP8gHWWkC
CuMHcMVIQCnD/2k+knefRfP1nMKiNAvbkV0NHMVqb9NRLK6G8e51MZ5d7SwOZuKSopRbnR5D/FWU
X/pixeQpDQGwLP6nFYgq/9BvWVK7BmNPFk1jpTEqSf7KY8Z1zTTUShpDTZaVx/ikRZ8G6i0Z4DXK
YBxD8EnJrQpDczuMRW4TzdNIBMTtLo6M9bYxZg6VM3nN7tZiAFHjU5OxCrhDBAJGb05BOC3VRbsM
obYpHFIFDcKliFrrGgTXZzljUQI2ymjLD7dMWx0iw/6pBUiLsvAAFZXm+4Y3059AYJEUTOimJSeU
0uKxeljlA2N8YKVi1P+VwvdcS0F3tM4cOBaHBAVnu0diccpF4c+an1ILR962R+IIqbwckknm/QsK
TLG09lZljE/APXpf0hz1ShncFUOgouk/trN4xxpvGxXI/y0urDQXHdAQc/2AO3tAHfOZIuE31JuZ
Z70L3qMgfDlVQJVW1WNPTCi1pQC+4bzCdOZJldTntAwIi5M9pv+h8bJAv2xqQTwgsy+1vrhsjQYs
oV0+kvngd5RYRayk6uZJYAB1mRvgzivoFab2CBTTCkAkw/NhUT3XTnB6iuIif0M0GrloSo7YGKfC
4rfFEihMXkfyMNb7OomrWlZrcr/gO/0D1a8MAXKEJ5gKhK93E8b7e1VIVvxKPaqx6fP7HLP9cyaY
DKCjeIaJGNU0AqJcwVDZvljwex1tulWUDc6yDexB++6vuHOmjeLKGSrrmHmWrWFM7wwWYWAqsHu3
u6fg6PTccmOHIY1bLmOs4dJcHmCN3gdrOY3XE1f/4jtz4a06Ju42/H/qjyfYQpAyQfOWFq0L7tLW
NyqNXnviuc8gT6v443EmAMmzu3eVnA6Pv1LsS076E9HPmcDwsl/BqAbMCStNAdD13k9UOxgj/PgC
I3/Iv8IhaCITGI5AlNz4vUQ+evDr2P/VPXlEi46j5TWyLq3yaN2MnkeB4Ta9loxRtln/bz1F1zUB
UpAKDM0D0SDVVTVy9SjOo1whZaHwYpaKJwec/mhinc+zgtP46keW001/elvFJc8VipBYqWaWtUD1
XlHNfpHcvsPzg6tU3Ss8zV6J4fvEsk032OoqZCvquZSFBE6Lh7Gzu5N0I1EVJ7wRKbBSBtg+lPIn
GyoYNBbMxSHGXNXj81S4cTLa/cI31OsSesbCpZvdLdJEOXhXnXcoJ5XzUKc4yS6BDo2S8QAV6nOb
BwwAAUTh2mdDYrnPaSU5e1o93Ee4/gNZP88/FBsLe+7OlIxVWxm4zCFy548TgKOXNNtIEidksxmz
sy9Xr62quQ6cUZ5wBLmrj311W5AzCxnxS8JAKCslzd5qymUw3d/AJyRBqx8E1LZ42MaBakkazdkJ
bMvkq0n1lVXW6qRjOvN02WhWSxScS5rg/blrOHw3WGyS3OO+TIRWGPYwV76RWG7FpcnTOKbEPQOA
I33Fl6AucJaI290vaid9sH2S0KZRvxrRjmc644Ql9gbSWoLLJOz+2ezR9iG/1zY3Nh0TnZUSl+fV
YDC/fYKZYxOrrrgwf1wRO9SDFmqaus9+9EmunhTNyehcv9rTwHzjOAM9z//EgOMfymfp40hp48Ak
XIV/yCy+XHQhaivG85QIPVCeuOougZcd8vzbngqBcqapBAmwEsMvytIb3w8kLIEJvRsB7Ulkg/99
J3gl5rieQUpadFDe6/FwHceXfI8C5cHKF+/tenDnjFPiUuCfR8++XHuNIYvDgh/cJzsmfUsYtkTx
w+GG82Odpi5GEM/HJ9J6KkYY+HGSpFEJ957l46hU7wQhk8t3D0GYB7AYOqWJ5soUvUaAW0W9QfFj
MQSxWS8+3/jaXJ47XG4TEafiS1bLTBggV/DLalED521Q2Y3tClM4Dax2BuwJpJb0HO1f788pjoEy
fay+25zqi6NtlfDRyQKl6HSXKGappqtBpSMaZwmwkHFXTi0mS9clRqKrMwGElaCoD/u3aGKpwc7a
d3bJmj09Rwb2Kv0xqpR2iH0FcYXKMia4+FPTOFIIkcfgPjeS3FMYgI7tN9qSMDT1bCxWcH5usrta
z05iPRY9xy0llqWseVXlWrI/HTdeiIkjYZjgbAsA315vbMScp0anjPnd2+Ix+lzytWicL4sjZs8h
HHIYmeVRbfG0HMDhQ5miKgo7BIMwdpXL7oTy7vP0exh64ownk4v7Gz+wMZ29JQ4QZk1bYlizM3K6
dbIzRD449NluEEX2T4+1y+jS7feJTyl6jsJ4mvn6Z9zYV5qtxlLkSjFcZ/Sxnx7PzWf5EtuJG/QQ
FDCDB15qIhnBJXA0P8bM7pfyuZgppmFFh/xnz6UguSUhbKtxrJ1N/7JGIb+tkrCpQR8adJfnSQbH
eKR39dJ0o2g/jrxRtZYFtbG2Q+rCPUHV5551T6cWCHWy6ANB5eUvKT9N09DtCEUat/+ZXm+DzZJ6
s+oAgWX0+pBO28Xlu6AVRkCQFNZoTHuc54apwqWBg8wJZhfucQm0WMrpVrBsbHhFULTtsE9oZcwN
+tgSsPOME5fGJ4AiWWEc9Yyc0IbqI+/vUkmmCrVrSJ5N13LdYmp68HGLfPxdX5gWI/Zyx9P//G9o
CL6BM07QeJq9jV8TWD5EzJ2pMoTV/ZonuWOadtrjDO/NuF43or3T2zbtxLksk6Y8a80QnqpJsaNM
+98KQRo1qfY8W4j2O86ud4J2sNd+EMh+7HiNV9WWV4QkjerEnQe/2O/b9nryqszrWsZVEs+M2hMa
hEcKrwVAyq6NeDcr4tWtRYpXOoF+vI5QcLUgdBEpCNegGxjiWfeemgZiI1YDPq41qCK8aM0xvti+
grQAORknCfQWQ8q6D9HnbaU5yr0iM2ay85S5pBxVc54ater6wATHZQ77iIi3M2eifiFTGndAGzMx
5sateDYl5iH9c9uVC3sBpTKp3lcu43Vo/m/LHCZfcFACux3+KbnBXmJfxSxWzxDrhiMPtt8nFJD9
rlkPhc7hXUSCWk80nF/5iHoa3eO7NZRSHPLLcDsDw0qNLERLr/fb1par9RVmwoKn9Gr7rMa+g/ZM
WKbADaTGJ8FCcsNeTIB87cRa+2t28oEdob6uEEHDjoXhdTAW4PIzM3XO2Ww+PEla8UzjevKK27ay
EmgoDDFvJs7qqT9/y6GcKb5SNYvr1ZvomsU81g4Wa+NcnBaluMJSEs/YKaJPj0qSLbNG8ENjlEXC
LJuzu5nz61aQ8gZge76eWfjfLMqKp5se2Kc26MBO5uptNY57FwYHhNVC+sW1tJ/vazmmkrWfesah
WeMddxnl1dTE5oUzMBsq1Wn5Q8FlC/Qs4vfDEriQ8upTxxDlHDUHp88cociWb/bmqwDmxUg8IRkC
+Kum/6NrTpuId0T99s7Wll4mPLcVD3WcXC6etXbxMDVxujTqaSvdOKDAx4sN8Xd2YnA41xstzEhQ
qSJps4nmsJi/ZJ7svNpVXU7lSFj9qIf2NZ36J4ce5uijIJelQhVRXVXlxRPJuQP6iWIYZ3/pW2CV
E1xBElGNSlWyIpT+jEEu0hRfVhJGH6d8CWZK7m/lp1x77CYokDu1H4JLiLWi9QoOljZ8as2NrhCG
N5mA3J/F2PGITGMyiQjdfPXgQMq2I2/3mh9pDIQgiyTdoN9wym520Y8JZEOLs2g4W7umCAI79fFs
0C3TJELwvwTQDfcOGscF2Mmvw65YzhnIuqHu1fs5jRthNPPth5RUhYp5tl4CPnRhXsiRhzNMzX2W
3bMtjU6wMfPswLd5L//qnEdHbi8NYpWGEYU2/A3Coe84CHDimJJkHBnbRZfpCBVEriUGtWOMwEMh
9P7Br/kqRchZIP1qE4QPz0g8UkgccwDD6j9fnqw5bMirGCeRVDzkj9znA4AoY5b6xls2AS7V5uC8
I2Qc6gPlRkx529pOMHyAxlnCh7Eh0jTEQCQDp8GHt9XJ+nkabdKpmBzqKsTIzvs87cEMXTjLXDJd
fEs4KS6NOeNwr2SHeGP3hjGWzXDokJPiWDodegDAvoyycXcmKEMlPIpQA1zrEWcCIW3UO6qCCSX9
x2Y+ZAoefd8J+tWEmVWr3Hr29nxfI8Frd557cghbVccAsXaveYOAgv4D+rA8uyU+S5LtqpC1rRp9
Qgd8fVj0zmyKaUNbTrLQrHe1VaCr9D0qdycavtd65sxXlhiE2v88HUoCtcdkDwHcAKqv3Pybs067
/u54ESX0uhy+zvMldU61OBtgtkFULjHqTPq/2kwJ+s/Vj4Wm07XAZV4TOfd8nOYLiae6uVgt7w6Y
dwqJ6wJfMCo8ECTRQZPKMfpTkR54JendXrMcGxgGXKBSGnQTBCDCWsRlrngNH2jhs16fjtzx7PYI
0CJOq6beuJYPKrDm1hYXZq8s3vJ2FG4CbARBzKzCl7nBC+d4mHqMlSslYb9ZWNavTxKXii24EifG
vTaSJLu9xTy+8MMhVJYY15lgYaQ+5CglLEoAzDy/vqef0h4MPHvdp9MV60DLBxZNMy/E9jPmXhLo
Q+QTQBOgr8ffEc8VTZyMDSBoDQmL6OkMdQns4tUTX3nPH/bEpWLp5elNm8qhJH/xjwJ62zAO6Yvc
qR9OewGXfZpfT37iM+R3NwyC5ps+Ar2WpPFAX6Zrgyj3CHYRQTrEwnhYVVmTSK8hIno3MvkjySoN
j5sKJrj0ZNTvoSdzKsYUDGmgUgMstDnHcLSUXDYTvDkUhWM/Y7wtEEJmNgZZaCbb2zfixFUpXQUH
0wN7m+wEExnts42iiirJ8Z56EIT6Lxc9Np1bqjbS/EVamxjGGh3vRR7FDHvZaE1+93db5AxzkqQG
L8qRDrU5jTdn7AL6aro819F4p9ZbzbKo+qr6Ht3jVaXt6CRE8CvE//WpHzX+C8QQp5lIG9jdqvLJ
0RVAqPwApP0unKdqGlRd0us9XiJzb/JE0P9OmRsQ4IS128s4VRNB+Op51NctPR5rbZA+XM1nqhP2
SJ4tVZLrAGSmADzZsqDKC0XED8oO1kf86NL+cCsMi4o6jPsZuqvSD3XPMj/ZZ1+tUZaMsxAyH30u
HfQiH3M2MFE1CfCizmsP+w2bBDLuGyZ91AuBROw+y3vQEf2SFQv5YaNfLeTsXh6vI5cJTZ1Tvd7m
CVYeVdG5vjryMVLNyF+Q+XLxhSw8XIksiUAg/cEeY7geMEjYvxxv6R1wF+reiyvwrbe0DeF3lU7v
KuSHezPFUuSeXDpAywqtPRkWDFjI6h2iT2sCFEJjVYshwOEp4ZStQALW6Ls6/Be9fG1xJAUNR3S3
DSaiFGFl0hfEobiEZvL4fQgbPxccOIbOc1nQukj/mWJ3p3LdjLeBC0SYkjxmE78us7m4OC077S8j
mKePHgSpNI7xjn3yeuvbbNOac5nW9NvahgGkXqaGoontvitb/49ZuVBD5Bpa9+R6XKQvEx7ra+rz
r2Qqv+6lXKq8ZwbeKKzgRExWB8usEHc/C9jNgh/ZXAHNoKx7jFs+jXR/1RLZKFQSXHZ5iQbJ8ltX
Io9cZkHd9o9FOXPQZZxiSUWhj9WgUnp0wIlG41A9xuZ/yYqIgmwznu4Z0HNHpRK6IzlJpiZc+7oF
gRYmiVMfhCRMqCTifbAxT5lJpWtJjNy7+GSS6+jD7s26vbb2an6yCDaxn//TQZOyvcelu7iYI/sj
Fhjhjn27hyOilVO+/ggHsv/NGSMP1FADni3fTN21cTBlIL/mCS338WLQyI0y2g9TASC1vrUxoPxn
yl67zKlIPs12jJn4lHFNfU03ffJDipoiBjtNUt7IYShlabZ3wSq4OMyBxpygsFKI5+t7Dbq6o0+y
r8jzZhrKrKZAPGgFvWxygZL91adij44nLCnjvSCaNpd8y3WE3LcD23eXCwPGnCUNpm/whOyDdxlx
NWZ/525hRJEJ/3LvFtDSCWeYMLz+5W0VdSeAy9F3uOZ/MVtklsrzIid8O/8WrphUFZ3KUz/eX5cd
fsS57oRCGf0K1RdjSJva1w0IV5XYvL3DbITpgwpYqI1OPXbu0u9MDe0Otr49xXO9R2visau5BWLB
/LOojNQD2vim5I711lfOxoFBP+SyCIoGk7MRlkcHaXSIzkqjcb2lDxAXFN0XJqE7LopPRB5lq+eG
TNYeoeAo39fo7W3wUilqCSWZYIfseQ7VYGXEjzrFVhijfYu/rdV+q/bSoTjPam/jYNhi6/q6YL97
1xaYDwVT7fvtfw5j08qF4LrbX+EJrId3bHxKL/P7zJA5dG/mM6jxPVriJ7G7hcF1cFHRWM0cQOlv
gJgpnZ5DzfQVxCAsgM4yNdS3gjT1APsYuy5ccLRBXff7aI0UP4bGO1pEiz2YcLFs57n3R+gkF4z6
JAzEHXvg7qmzYpg6BgSpAZfbk7jHOCdq25hGLiDl0YhFfTOo7frGvG0E1ZFpReEDhUN1OY5ThWka
TB0XwEFYUVISIuwp9vwdrU2Phy1FEMFfRVbsuXxXFOVS4eN2lPvulEkw4yuoXAQg+hVjzGJgbW4z
UPzv/sUOQya5OZeuBi3kbkscdd9cy57U7A0VzSS9fac6DOHoZfaejpJUBp6DLu9LeGUxy8bmYBh0
ksp1qNp9FmjnrhWqoEYh6rYB2ggw52kJV2icYgGmMv/onXjEGxsDmxO6AqiLGIL6vGNaxz3rUQo4
g+7TMTcB/NNa6qMxw8YPa2ctFPII8pewFbTU/QD/dAEg1UbHPdMANTAFxobS2ehaAnZqGbJkOo81
V0CHX+pJBDvsXRhXSrDhOrW2cJc8MTEWoTh6RIG6+l3JldNXu1BqVRerMErLGrwp7BTtncn1GOsN
qkry5Ms4CuiO/4asj8d9VOiEi4thdcWVpinVQCVbbb6mcOuBNRHGe4VlVxSYgD6HmhSCGeGIsM9W
IMHehLE7gA/s9b6rCnt4LkrFcGlIPOa2aSKhS4yNJm4EaMK1ovILc1zWLPWSEOIIGgc0IW7xMa7v
CaQSrvTI73Faqqng/+uECaOkdRNLMFNcz9IiirlXJ/sxudpZ1fhnXR03F2KsoYEqkYSuCD0aY2Xm
9/0LYU5aqzPbiiyA1nykbKP69EqnlfN56Mk9XZ6Sg2KaalGngEqQEFVbMTzU8Q069bRr0iFySlD7
LfvL6RoCDr0RO9uULLZPgSLmUWe6Ci7OS2Cyi/Hs/4B2eLh/aS3IVIK3iP1Rydz/EQfqwJYX6H6B
3gFYxOkrbSQDQGIHE9CnpPiup281dVidfoWAYuFtLcxYg7Hqek1JqoHjBlbtSVultbrAGdaoDIWc
RragOctjxqo5w6ZpFVKEDbnNZ2VzWaYDLnIbdHzY37rgd0Dwyg8FTV+Z6D7Aupil/4MSy3jUW6GR
iETTsKG+rMxBZRIE/n1EF+BM0pWVVdUj6P98+8dfuHCXtPqg66VRjSj6JlrGkHGbpe8m4Wz9L+CE
9sC3dhoayJLtx30IKK5kr9eVsQWeTJzPQ7n/K/ZI+76yqb1N4/N+lWBVyNBW3mK+ac2UmhyslCh7
O6zwPqr4QuRQ6Q0LnylABSHkI+vjskPa8bkY6bZTWGm2yUEpCFiMV2nvq2/BKpO2Xa5VpS8RP41+
pFXEamnFHB6PRn9S7MyEDYP5CkacGLBe1XKp2vFkWuegkTyreXrncKuOkNM/PGANnyqWSWPxmX0o
Mo0v+nBQLT4bWVVx/QG+diYDYx9C86Dr6Islglp5Oj/gldTTqXZNuMirQ8h1OiwnK3aQz5jAad9Q
AQm7NZ8lUS62JbeSQkpQDAJPIsdsVkQoe5BKGXi/CODEjDKXea8UwDh4k/Mne+oxoD0GudQQe+Ah
ZieXychDUTZkM2jWt0eUBxeZSouv4uEJbtVR9ZsP/oS6YGawMZeboZ8euTQhctl0FrDvbAyygMeT
V9TJE5cVoawAr7XLmexdOcn8R5cxy+wM0u4f6Fm7I2dyOgDMNcVy2qxq51NxcLRMrXCx8M/B98d2
Vtze+cgLoXk18LmARU1dwR+nlz8fm0qY50cNTBv1ztaDRYtUtpyCbVg9sZZV1Cn7rGqvpWvOCcyQ
Qu8RpttOiedlCgriUlODNxMXxmUUTG1SmZRvcFXUyEUopLDdFUCN6kupZRt95ENfVHBS5DZaIxIa
3lAgtb6SL7ejkfIdS/P1zwk6Mlu8K/tFZg9MFjIQJDmLw9k0g+rq4SrBNq410G2U97Lm3lXFvSgf
QJyBdNiS8wQyO5+boxI/JNQd1GQyB+bHh+HpNvXsW8F2XfkrOF/iydTFnx4LVZ2GU1pIAGsdxza/
+qgiCjVY8c1+wU14MWSzUCM0K3eGnDVcu6StYP07g+4zYvkI5829YIooEAGjanmRk6ttGlxxiSX3
O/opl6WMfhocGDyfR2b7MvZd1lpGIMIv3+F9Ne/5zy79sdI2o50EJenjzPKK3IKgI1BhWEKQLLra
U2JcsOJlrzsQBP9OMG8iZyRWmC8BMsfbXT2crSyqkfRAylllWWKfbXOowKyaC3RAD8Pi8wA66cS9
cnAEBXIhzIfDJMkgh13E9U9lsOhxyK42i3fuGK3vPcuxyumG6T0tQwWzUEFC4NR87/My1NJNnux9
F0v6EE+KmcYtlrI+4n7EY1U6lGtcDM/5mrcunfKxFKSm74nqCKoWYYWA245O3LJLsfYG+Ju0MEdf
iYI7aZfZWKc/vlJ0Ap30Erz1iYYOz+jfjGxapVuqgBPqCE95zb1tmiC12OHcC4z6u13bX6uVa3kz
7/wHcKLKN+7EjaduxX+60UoW/ZAfP384u/TLSxfGQgN4gpdKfroqUGrlHqkkC+YjRSao7yAAqWrj
xJsLUqwdaygBQjtVQ8KJBIMFNGb2ii355pKfZJcbn2Emvc7tcAtL0PAiZsw1YnZYLIa0dqhclvyA
d+9LZXi6pl9UBVJrVAj1EdfKZ9jd6aGX1WVocx4/1L67iqfxY7w66yCrNAvCY9xSPIJH86/nYORJ
IWMwvkps9RM72MSw01K+zTUlM6MakIroWd6VQY3rPPmjNjeIV4OJ4L2y9M2PP4uSjDS6U+XXsK0o
PsjNLYBMA4ajT3A+7hp3iN4TvwHk4y374IEwrHTuUMIIvN0Y27PQE69tvRl/E+5dZ+tlwDVMKN/B
CyydxLQuJUB7WxKIbkGB2EPy9wd2PVJMkbwzsX/5e63nP9vcx8x0OaE/1P7Wo1wW651QxmWaPYtv
uXmltquulN3/+aUnTljR39Xh2gRdBJBIGpL9rm1vSkbl5Z1m2Ywi8QhiTB+7ZsEfNkwFNrbdujPO
4jEQny2pzwesnxSq/oTUqZnbAvFl4TirrdQxZSnQh5sFDJI8N+e/T3qzFYgXgs6B4XMhSHFxyMKz
peLsPWDkWYAZIt4/tnUJ3wkecpF1elF0V9an3wVoLCUqrEtkBp1Yj9xLMyl/4duMgWZcVpo+m11a
cD5CrYKUBmaHApgdBQUwe/N1GEf32hnfjYtcac3KQWFw2NCGJ46TKSChBdfefGX4qAGkjzloOpYZ
8LvzcDxOREXJWMNAXPcqXtatnG3z4FxqTXMuSFBcI4KeTdHn/42EvgHCmS06ypr3pIYrj4Ykt27b
kFVGqA3rLURwGrwAh/fPBLQ6ujAJHV8ypwjjwim5tPe8tTcy4z0it8g051hG7qTK5cmjui0nKaFu
u9ZNtX5TdqqRjn/yHe61qVCWCfgmuG3XNBqdWi6CFuZHbEh9htgBjFityJ4/uX7J+mSluVpFggvR
+otL0nOY1cAFQq1pOVW1j56BlaM3BIx59cfLcOce2air+GXESiZanqkGl+VV+jcTK70Z3icYQ2WZ
Vj6EH3knsAFPM8pBddQxxUd8Ch+zKxXqqtJFrLtcIraAQZuFUdCWajrt2GNMgDA1NZQKt8zX6mzM
n8jtjttOBLV61GDkPVg4DCXXNYfwtrLvOvuk9aAiqqIVwVPi/uahgSeeE/j7Q6HtuVQ8fgl5cnkE
pqhSM0nh17k2MP7psJ4dc6dNlfi9Hnr92xZvMb0FuaRu+zPjqkBY/ZnW3XY4LmoH1TCbCkwxnzTU
7RybkvUrz49U4lleSrtwlo5bmkU2PhPaMyljlPTHcysQpD5IiHQgk6a61CjlK+sSEdwkmXaPqCM3
3BTlh0eibAgw+EUVlpG5w+fxsIkZM2QO/pK3EnW2y1zIcT/luLPxRQq8zJgrs06AieUYVsgoTkPD
6DSGQ7nBp5tMFK2U8SnQaOlp6S/8HiOLY7vzQ/fiSmCc+ISwrMuWXwVm+QPNgHicMkEb2667fOD8
lVWijCjoEBw6lPSK6T/svTI/mgCSDrXqjGHilrjynJft8X5VGFQK7XT200XrnRbg7hM4/aUv0/ng
mIB+93Ii4xKGbxvUfposUfephWJgqVUR9JCxRtxRTK0PL4sU7MV2MuzvpAvl0JmLt+xPCHd2iM0s
DdrbWW8L3/wmCrdjrB9VwcjKYyUkALC16POT2QOrVH8V5HPQBZZOp7PC7lovyNhYoxnlgDaeBkI2
gIeB+LdfqJpKO5OxajqTbnrrTQ0Ck24cj+BvMrhIsSehe2bX5dRvEqzO+wjRFh1bKqBHD3esSnJr
p2SDRkduQpzmfeLw5zesyNyckauzJfqrPvIcDrYCR3deXlTU2lOwuPXWUoN3CqSwYdV0GKThi1Co
VlUsWOLd8mUuOElfRQoXk+uszsaPvo6pdyhg6iVX7BfjcThlXgsTWzPuAH/Cnfx+Oa5tJDfe4xe7
NuYuszJ332Rg3/oLjVhoFVALlO9gqLQ2BEC8gD6G4MDdgynp5h9pZoURq2z9dI5b6sl0F+HHgu2o
ydNbOg4lJQHJFdxS3vEjhKs+CtC6cziD+1iv+ezgX1SBU6ltdOXwJTycRI+lq1sJOE+cJI39dB20
YjUXzi0Sbfz4YXyFw+lNsdcLXOSqm1AuqMHj+bWsw8pxQLYwQiqZ9Ot9XeRh38OqhYvYvQ1iKx0j
D3kNdOY+eHTeUc8EeNwjTt7iTMosSe/TZXIQj5zhyl8teSVYSOLouc0ITKWZYoRXsQoejT2d2NyD
ZdDCpRCIQ3cedK6XGvl4lq2RYuBbsu10XlXiwp6Ni4OqNmAhdoDQNWO8TwTpHLbbru2k1hvl1J6a
uTeTcOfVfLqAdYeSkGFTKZJRPk9NFsyzbxwUw0HD3Z82wpYmfaUJ01Blwb1ffc0YDbm8Kalr+fm4
DUO7ES8f/TcDA3Hh8Lc/F03M8SIEtUUaz0GNvuJq8cCyN35ta7Hl95Bjh5gr4aUR0+8/sqfEdifq
V81pmjISG8uJQHrdGykWKcYN68i9wKvgsx8kCzCt0a00AU3a0AyRhJZ+/GN1KQE5+/1mt9BIWR+v
mfgzJTOpuSjS+bYRREweppjvakUS1Z2MFLG947Gpk0Anz6X7kYPr2ilnlpoGD0WXS416YC5goL72
MIgxFLsAqGPbD+FhpUbgUjW2V2N5NzDJa+buL6bithRXdU+811zQPlyy2+H3Jq3Rx9dsCqOGL5N6
TTtO66TgB63ggStF8wSRqIgUMPpBRxefOktoFisKgUyfNoIS5ytoQGz9GXehH3wBQVZXsmkIZ+wn
K8SLtE/wBgGVRTqVKv5OZc/asDwK65eoiOeKVsYCYpYktj/pSGUFnYvbh0pRgXuIMDC+Fx35kV5b
W0R9cvWAbJVHGkmzyzd8KWRKaOAJUcDB8e7+P1ot9OD6gGeR5y6yHdAbpvsR70n5TVowhpMLANSR
o+xYfGwRvQNQK+5/twLsGVkWH7CoQ9Nz+J2TcX7jdtsz2wY121OY91Uai/iJ91l9zeRfmJ5HWrDN
Bxg2Z3rt80wYvsMF3/cr5M7QPSZ17NkLIdzlHkXuEoOsz8rwDbaR459esJsyOPg2hn8DanVIyroE
iu7wbJ6yIxtjEWAsayjVv+8mZy/r07LMW4WTDgQHhpIv6ZIObHFLi5IO+1OviFKvj+OWUbHXAQIR
B1j+f8ehtBLMqE+bpNdJXtmoqy3osHujxJ/8xt0ec5hiiCFcxbIIu/0Xsb+Gt3YulCV+ptCpzO9r
8DqIxILwDkFUM6KtiFXpUDgyNEpFmSmqLuZY0rHhXvC90wadLXYcF0I6C+ONE6bz2BleUiU82CqB
fydrPqKqJdeeokXijq5pyJ30laZS3toXSTZA9KPtiRbQbggp0j9MpuvtbzCB/p+nNC0uys1VSGCS
tg+sZGM6HW5M73PNI4o4p8Yf3+Gepg734ounlTXpTgY6IQ3cj7cRcE82QelJcvyHAMqPyMG90Mtq
NG1/xvmbfyy34Tjefiu+XFVPHwGd5wsQ42QOJtmaolz4AfLaw/RNtlwfOr4Djlyj2Mjefy9c1AS+
BPAl1JJg6nh/hN4925JlxWqJotuvMYpLjqH3yo8+OSJX0Ad3f0YMcVJ5FTscz7zJBHHYRetCLoIf
eK3diA9/fYYazyl7/dlzxCbW9DvFH5r8/x01i/b0mymNs0poEXdyjupl00OqYMLPAxpa7FDykAM+
ewCN4MsAZU97tSz+Zl6d2ec7DnaF0O1FHZpm818g1OyW1PakfVLfmB27FlZYmrQ7rd9OA1C5ldM8
BZFP3nZ1/PVcVW7+x3X4Lhv14Ov4bP1vgM8Lajop8zrUe5nazp9scQgXlv9RyqY7eHGQo01+2Swn
1mBmplX39ZYVPJng5DDqrubXMMn2hNVmP5le6gDScpeSegizH1l5kpWiWhGU5Jm2TUJ+8FlNqcTM
hwBdwjfYfk+1fcsvG/FSwrWBW14cLPLrDtqq2SnG10v6IfWKl7i99njWVxRgDtuIK4XlzeGk6JN4
UPlJnmcxe3rTD5HpOcDB8y18iAqScL5CKSYX4CRxPgyy12QYBSESOsEA4rsoEflL7ABuUhXfzTSo
n0FeM6lFoMb9vH3rHS1FUSqCCNpjCMos0IYhTMb6dG5g6F3HEG8FburAKnEURXPubpHvNS6+dhuu
ctgHMQw/NigpV49/s8LguhBWAmzhqf7CbyQ67LUjUsjUau2iZKgHVC/ZCDzAApTe1sit299mSJPd
dIzQPFWIoQmBkSYbCgDOXjv0eSGvBWLnFjCLarD/NNxZ6xulrfT3XxrYx7d3XXxrfXUEZg6vX+Sc
4luyDS7Up47SAvNSGRbQxDs1S4uce6O5EQATHece8UjcWP7rni7rPHvY9IEdub0UtNphtmPxu2c+
vMYkM3VXjFvMJlYhkbFYxczNEObENOHYuo+p7tYRKMUSc1SW8mmG2etaprlf5Nslz+3+nc7/SDIY
xOLVXnqnApPwefZz3SovJcAIzbYe4EBUzodxqPozLxCt3Je/gFvDty4WIn2IyhOWRuvmw/W3mEYh
29ixQyU6B+owDno+LtM/KKXwUD49Khcrm2J2U1w6Ptovc7dmQxBf9A/H6nchJXrGMmm4FpxSMf1L
FIL/cwToVRvKkJGhsB0d8EmnfZjTur92X5SJiXjEiLICMQ2gdCs+pNafSTKxPXNURtr9GC8enc+b
C1Gx6/YfLN/MuLJgo9NvYRT9knmpEyayz/lS2FEaYwqIFPii/TTxqHUog4pm9zKiMfg2sLl4gE8r
iNe5c40HwdEQtjepxPaTD2QEIUKQHRNK3eeAYmOUq9d1sme1up9MyLFtr0uj76bTvAieOF647bZR
DLfoM4fVLT85lizy9ZLw5BR46bleU9CiYpDMmwDjoIVNiEOEHCuEW92zvTJEZbFBssH0M+5dJ1j7
YxmBqnfSNDUrg4gWkMDU85qpddPeXbqZQ3y9MNdiVrZ0hTERmvSfkoxlBN3vMIzTX2jn403ncmfo
7P2tooBlnwddzwA2H4kEPkXR6AOl4yNAbznr/6ZF3VIZ2AkZ4dyDPcPDRa6rOH/2/rP5jwAnAQLk
5El+a4vvK8bIjCXYWSoFv0DlN03acPUFG5hh/HYyFM6/NmgV2TDA/bHN+w3fYYMTyWNf7JXu3EY7
IxJJXSIqWd9f9tMS91fNYPKZ6LnYqr4Tnbcnqr9FuuzGPuESbvUdaBw3TcHfahrw2wXxFUSvuJvl
783SV08xEw/a3Eik9FmtaZ65xFlh6cPRwTt92uhRQ4HaPyn532i8QzLVkpHzttKSJQWS/f4zsLTI
4HmhoAXQwfGJYTNXkXeZS0dtXdhkxg7QUp/Qq68Es+5bX9sFkgQOtuYkkkeFdYwC96X/hpVB+1rn
+h1Y/2k7JqCtu6PApnGVONjZ+olJ70Eygm8M17jXsk6Hp7BVnw7gJQsmruQmLjzP8eNvhuPr5B6a
HjwJIDpToElihtC9G1HVqhvTvuporgBJK4qHjsxueXdgQMtUq3de9zDSZqaO+oXw3lXM186G9seQ
56dSfknLVT37K9rTH/hQR2/046ooMtQN0En0n+vpfPwhIOmYrDImipWW5KRSXKmWFQvgzxxwJ1c2
We96cVYq0QbFHPVIJ4qtL3EZ18ne9K93xPamV37b7v1E0WQNsGnB3HLlUB9pk4CsHfIxfgdGPdta
bDhwbui+Q2OoOc6jFpmORjQ0yaw021sMZyfIhb/2iEWajdLXJTA7lMPtoIsX7efJAHqQr5DYmllh
XNcO0t1lSuadXYIuBLovIu2Sf8tO1uE996k7KI65zEq/2Nv/vSojtyymqXnN0pG1YCtZltdWB8gb
FSPHtDq/pBVVXhkMhHmIoKp7r5HM/mVwvKgUAGfyrO1TUvet2qt6in0C9/sGaPa56hCcsGWZUCFs
BLe0mabXMxG4lPOISKVizqMEVWzgxJSbPiKz03mjBDsCFf00iDlDqKDHOKu42j+0I/PWy9F00dET
LO3FfXsqcTAA0dgAC4LOPzOjEieOUDTfIouwzk1jjzEmnpvD6rhZNChIxK3pazF2w8JUh/Y2cPSg
0BhHhsh3iNTXw/wkRbZ/MxV+T9ZOxQpeNFLChqVLdAwKIWq1xCWmFIC9vfyQL1co47JwkFzB2LFx
JoYxmDdAiRR8LF2hHbPELuYBmPkyQd0HbbYEIpQb82EaDzd8UWumiRZhF6acg3FD3A1fKGKe8j31
uAP4umqcvnCYD42lT+GD7m3SwbYUkdQWJ0r6OoxmdcZzC6uXad1Dygwl+pbSi40flIy42vDXZPLg
4LDwaHSzSbJddv0QfSsVobCclIdpod/ouzcQyKFQmnXGQnVudaVY+wsmCIEg1F2tuleu8ixbrdB7
GmYipacfx6062zWKwFQDfxufzPU+dxt3QeO2fOcZCZ8HmiVGelrsizXr/tUf7ASHXeie0Q7v4ncC
x6xzacgHp7rKA0qbM9Zb9aLD60359eNRkog/8vR174RugYlM0URji1iLHZVOLcSWrZsZwO8XUdS5
1EVm/HtT6FW6LRnPajYpGYzNNptbidq1BBRp+qjK9MCl1TiEzPDeDALzn4116g2PiExES8LcdIJi
aZKlU/ieZmXeOnSPSM0hIDDQ+uwCmv8/UCl4mTIQe/qISOtMp5nae+/sOILwKvczeaVpn3KKOBZZ
oldapsjKtZbdIn39VWaLG1V4Rwi1ia//jvdFKIwR/89+QtU/mB24+EJfflnhp1ktF1UFWcsrix6k
XYsHgb4clQ0ElxpleiRDo7hcaFdOiWCgqWTbV5xtQYkLRyMsL+7Qlo0lYX5M7+6i6Uw3MMiRO/O2
Mq5vujQ+YEWmcbSTd829HOMD7N0ufj0UwPvQm6mNPkC0GszJRLDEvmJekHqNtQT2E9/M+LlLCe+M
u7Sk3xXPVFK5a1/xYctkknPU1hyYGphnBaJYXGLg6XH3XusrKfIzpOUCHst3j+4WDNbMip82ACCB
FOHEwG6deUrifnAIUeIOr0MIBzdeYYYAq6YMWSuQyBugTaVcXyfW1YaHDZc7pqdK4yLG8A1UTjk2
5TAA+AzHk4MqtVYDeNns63ttZ6YPEFdzUZbsHfKNgVEhcUBhjw6gjt3IrlD0dbiYnutniy4WKoLb
dXwZ+ebgtpCkd3cnrCYFe4oXz/1+3sb0O5x6Q6zD6HZowdn4Mvp4/w4Okk6eGqVPtMmEkV4fvDT5
wgAiUJmTlpn1K0v1lw3C6lF8N2Y1PAcmFnvDPrSN5eNQZqSGpDJBqxqL1WN4N6Qzue0q35kKVkAV
xwewWnvURVaiaPlSvSfYlZ21u1VVxxUHLZA5/Sdk3fDCNEyeJOKfgtzlR589xeJct600Hoazy9GM
1oCNLnQFswDuDx3mCu4PAtoPsk5HE/3uGEXZ0lLppjWy9kD0MPDsyvxMbzPoMvx/wflBXrcrACJY
16S2XKJFVUz+I4ThKBH5xETXU0qa4rJnNP33npBpEKwHLYD6tBbz3FmUPWzJpvmLk7dWyp0kPnjO
LP/Zf+gtyfi3StSuHkDL4Ioij41tPW1CHkgiyJaRwY9chKPmLESZiIcgaAwQLz9CWnwI/4l67aph
OrodkWpFpYJIXWtvRuAKv853EkMaNrqVCUJOFYgmaf3EgWzPwcdHHcbeB4eu8es7LHEZRDN0QQUp
4Q5oDc5F8ZV8PlWAwN1s3V/alTMfHpKAeaJf+fqH/IzxdWu7uHb79gOdNfCq8rLGJVHQ/VgqKnT+
p80vlPQ5b3XczkrnYgZcPbx1O2IrIlXMBSDHsBEs2/Hvn3CrUWyCloTY7BFju0Y1hrhOwsPB9CW2
m2/zIrI/eaPbxmkY5KD59X4TiOR/YUppcmsGKPbp2cVccw2iB3Fq8V3aUDd8B7IQwc1H1eAV94y2
t5qDee4zrtMFb/rYeQ3Msxwi63WBm32YecMuYjwkEYpkYdUs8q8qJGb/e4nX+vZnjlky/gZnpm8M
GoOlv9vn12Txzfr/ux10F08JOaci7cxRz+6iqREHoHBitP3ol8nRSNudK4NGt31qgIg/ndPlGmqC
h2C9M/hTpAblK7ypzsCH3qAdPK8sTcKDoBL6Ju5g6Nmj6zyU7uDNgiSYZ+haToiCRM4taaEaWnEd
wYx+gc5FMma1xtzOjTeCaxLRg4MQbtrwCvRUgJ41ImFuq6Km0tzMuxMLy5uXdf/qtT/UoXGD+/Qy
wK0by3uqFkzzoKN/1hLQC3g2OmUZ8Ch1WQJdqVIsNyDX+6IVn8VkdNHxjEY27Jo2SnBHenRUlGWN
LRgHVLLAS4Bk5XdfWkFCYo/mHK1JIAW1/TdtIkYZ2WHAUlFv81EyOLvhFSp/rs3lqYy346A7of0t
J+9eK/DqHcE4ZQDQ4KaKAlDbO9HDicibOfK+bodH65HPrHER10mjg8T157VFQNAKlFxPIzn02MhC
G+QbASSM2ymkzc8pm56Xux5r+dplMV9gUi9KL5Hghx6g/VH+zPQHZ5+EoIlO/sxQwN+fV5fcCECl
oE3xG9Rowjt6+i+3G69AVanGM5mKQ68Cd7U6VSFY5ZurLqOgA7pp6n4pXZwDeGVSP+FBdtlfw1Ae
0IqewFjwDlEdAWkf5u0pCIC0rB+fhNWWfc2PvOXBRNQgQkWSPiYvQ+eMJZmbiC98OtiZ/GTvFtOT
YHkguO3xO2nTvbtb2IVGGVyNnCskJ/+WSddjuhYeSiT+yTdNDBl0I47yrkHvGECDVumlcPmU9i2/
opD7/IOs/f1/TSnhi0uq9H+75UypKEMO4e3VdOyQ0Ahdn8YcLObkng8CEZ4u6kphJfUiKHFuK9WO
k5b5ahjwwO88488iR80gq7K9NBPCiuqkLogWT4Cujs8sMgn7mXNo2n2w4dybxBa1b2zgBNbEaDDH
JUZnlzvtK9TqZlgOCxMGli1aK/288zced5OYnokJQsSES5r9/WaLizmAEJ2rSjra5SGTsuY94/l9
i5OTQ+Sd51rE5RV4tQou1HmdapuDPh0uKtN4Rggde/y7NtIinN/dtwkNcUxBLIPEwk/6geCI4esG
lQKX+RXXtUu/9LNTaNebZF9fmUy/LJsTuY6jhbqcyvB1ICkVfDICTc2vShzqpzl+FCusXpEIAgMF
ocaFgyG21DCc8mQMxapz9wQkplgZbK+IxfAaG/YRe72CNwv/Wz1QKHq84lbj+1Zps3t7JL7tRmO9
2vvTVLbUKOU06hMxnvHDosjfdglQpKQNJXp0uU5Gap23qBV95Vx1T7VLGBqkiwH6DqWIshF7RztB
PLjEuFfuscTaz9ug+AYqp7SJ9ANawx/O8AX6xHq9PP5xHmZqbGR9OjX4j7v1joxGSsnrYzX/sUJD
iFGAzTift+V+TYNy1Bt4APSyE3JlqqqeLxLclYwK4VM7wOB+uyKmmy+Q0Y8cH3aKkmCOFSO1/Hi5
2aPixlLd2Vj2DMjeKqABKT+fwpgLvfDqZA/8QAkiL//StC0MwT888ecLsIBBSZD8r40RUmeqyJ9Y
ld82iSeif2x+AwYvBjq3Xl2Z88ZxFW3+TAovuzRuvhPqYs3RIbr12qVAci+nvcZMyuc7THpGnKeP
VxDdvckBYabzZa9sC/LqX9m9OJcWLb7OShuQ9u7Oiji96Nemr2AWwbFrYJ9ER/bk1ZCVhAs9E8DT
wPkxXOVvrG+1o1mWR/GB72RXH5SYsBKQPhMZyvhXSWwTHsOPR0WKMRp5VpWVO6+ehtTFPfBQIM5Y
DpSklylGqT2Vq3z+M9rhxEVwSGu9PzmNt8pUq6xIUBYb/IYutnEwW/n4hlRw0l/pdpyMmZWeLE38
lUqEiCfPoaxllzDCPfPZ+9EzOMcOSh0m3Ry+i5en39wZYSI0p8z4s5EzUWG1cISgxYqRFHiFcX7n
TvaND7INgagc++rHVWqPiQQvlZhy2Mmi2nT4buFC5sCaHLiGLenoiz1Z/KEHy1FHzqvR8QVT5Pj7
LtP0RUYKe+5Q4Ac5krTg17zWNkRXZwWBa+3O880LnjlDlzSKvJvzAHp4Arvlz2fnCwDQInFnNz5N
7Fdr2dBwNngEWRQ6HCl6LwL4Q0/jy+nuESwQwmiKL+e32FZeOrhyq46dnvbTg8FoNjvMKJdqU1xh
6abSeWRXRKsuRhoOHKe7vbP2sWynuYFolwQNCeGsq/azjvs8D6GdnJHythqp3D1U2ShnbN3zAs/f
vO8ueFxzl+D/vmdLOI2WkWuWpu+bleiLALhvZxQz+klZJzOzqUUGyAdCHHDkuUtMCMIkbcLQtRt8
/XnNHq4CE4uGAUpFJR3AtgwfSSbL2LRwiDVIuOPWTFWEXMPdFhYPk4fUrSFhbAZVIdZSg+1AXD5u
+pDVBST5rOBDnomsRpmkLC7IO1iPMb8fmjuOv57qa6JNnjtrSGm2SRQD50KwNeBBdp8J7e/y169i
2Qpvj81jnBNKPus/Qb1N2/JdYQjQ9X4y1FyjSqHinNTodh8Eo5I/UJydsCnShZja7L7T55rCXg52
14eHTpfVomzad4e1dJ1W82peB1Qk8Xg4Al6QrJNfasDK3ouoZHSL1JEqHGW4diw8c+zyndIQpMH4
meEBY9uDShJH+yyQ042Qmfy3HLmCTaRjRm0ze4uJthEiFGtdFlGdsMcBgxbY4OvjOm3MZYFCbC35
+NPSazK12W1xGXqzB+1lWJ9oCeudGdwAj38R8Bj0eHFKxGOL/hY+nXHoiHzxqAp/lC4WYefER3Y5
PEb2nMUaCNTN5RpeZMC9AXcHlHKFPOhTxqnUKWstdE9rUHLPWY1soxJYrMcWlTeaAo1ADAG5jkH6
/FG4MwVwnd8yejzbn9xmArWiaX40e65AIE8QfA/s7z04eQl3L1ETHoXiWQXV7bEl7BQuh/96fbNy
/XnqN9KWrl2DrI68JTEJGMYTFDQQhTbrs9GMmDX4+QSvRni+GCMEvK3xk0/4oEGU5YZVtCRDK/rX
92V2v4ZaVGzQu5Jg9+qhT3mR0pgooOJE++zFJ6CR2KNXsj9Zi+bdWpHJ3yO0mPwS4LdTBEpb+EQa
QlveFssv67vUaZbpRjB3+AzqT4b8ImqS+0aYq2egemaxMRsodbovzPcvb9W40Atuk9uqsov/OZlM
nS3JH+68UcLbahI7HrM4y48u0Yu/r+o3VaxL7OJptcV7RYwMravmAaMyJ3GgLBhZp6RG3yo5cWAH
jKCQ4tsA6NIpgG3ervXILAzSJBFHf+JzlYwQLVTAYo5vHt6Ge1JwrgPObn+/FId0XJjum9YdWmZ9
hTjVvTshuOYGb+INLi9WgiDumktwKtSlTEQvp8s/slhM1ZXLzrdnpsckkmYCIQ2+ZKmZTYQKM5ce
oCHvBlc2fcoPUPvPOrr03JiZfeMD2sig2GZ14/hHbMI+F84cozUaPo5fwgDfnl4pyRH9hjBY2lP7
Hosioalxb0o7ANaohxs0f3xS2IMbT0O4elue3h+mDNQI3HvHikausTM7i979deJHET2rutW41eup
nnbpbVvd7SxZWLcrUDtpJqnma2/BYsPOIfWMh4TOm9GQOU/arJOlmb5BDSeUskr/OykXfQ24vWXZ
okDUgK/LTxjyn3qQVEYGXfrOA2D85hgR2BxDSdG+Cfi6LclcDdaEBgCytAi/hDO3GVTJV2UzhoKN
kaqEYr++6S8fCAsEZS4UIKJ8aqY6XNtYPSba4gXJ/C5/1R+bdnaEzb/1SdO7UCrVd3rNFb6a/RH6
CY1IluigNFw8+a9nz63jEQ31GfpteNCSyDpDu8tSWwm2zcYmlX60bolOH1jLmD/v0ovW+WtdV9qh
U1C9+S8CbdoaWFHRW9gzt9BgS+HqPWooscQ+mjyWMfeapzZEVAGgjCj+fnpDffuFKCJoHIYgNWOK
RN91zdKNSKMYgUqjVy7fpIO2a2er5qYR9/GFFQjfUdZV49+V9TPwwbUtWz+hrrThnHGwN6YQ+/6f
ZGCKyZSeNXtS5ORU5tftYZ1/fmoOGgh6YnfYnNtQLnW78eFk0s2XWACKuFUZhq2kLTgVsrve4naX
WYcA8CxwV8hFD9mDxbuGUQ5ZpMgf7mUUzYol+Dm00ukaZWlf0pAcDsNlCreryMb/iS+HKHFFefz9
VuNY3Sm+qES4XJ/pj+6Hgozt84+BZ72yC9C0nCbapWVFnashyOms+gxLBR/I7HBqBCaNn4XsGgvR
cr+cRdzohil51+X1TXj842ODqT/h9satGhXLP5PoMYX2KfGsnrHGtrcCgWR8u0Ze6LYAo8CrNA/J
8roWYMQOGUp/4P65Hx5PlN2/Gj8hzsK71KLj22WOElyGy1XWrjYJ9Xzfu8LkVUMfJWfjN93TbmBq
ry8BNafgMSEC5kOiYdBy2IuTmpWNe5s1yl3/f7ZW1tn7+9rLrRpobqmezdAS4YsbmPPhoPf26pie
opOfdmfq2NewPjO6L2ojk7tTs19D8vBD2YK/8xAbIaJ7I4FU3u2fVQu9S95ywlo9yKlsN5IRfv3j
NdoGDKUDHwsMq7iLr7p/ucgkVM4Q8fBzvPzeBC2duAgiG1OKExZitNeEqK4SHcWDaQYqGe3lOZjG
taNXecTkK7HG0ozZxswzA1qEOaohCoQ8v+Oeo8lhiOP7a32L1USil4hnpvaYRUHGCpb/HyNSOSLi
vD1K6tyX8qqaKYywcRzr0VNerq85mUtbWS+OxSGXN5vWmRyYgQiIcFH/rTwtZQzbvPIXjCfhET18
U6KoBjnxWJGQCaAw4kjNeTEIPe5+o2gelAiBHekAAsmse8U3LHG69FtvBQekQ++UfXq7V2mn7jKm
r4OfMYLNzX3XsHJr9w2LN1kDjo9B83S8WjXeO+LjAkvkiDLHZVnuTLcnTenzpKwfOgDjVVbGCz9g
yziJuKH9aLeVoRfseqLhJFopP2o4GwV5I9ZLRUNj9zgkcj/ggXhZtqeXe1mvEQLq9U7hBg+HYFsl
jS+9niRKyoKFJdXbs7Xn+6lZyY1YT3yuA5g9tPpy+RfJCQ2Psp6OSLfoV/t/YIOrFCxsXVH8k/Pj
V3H913SKYI82X6xabiyGgDOrZXHgDbNxwzHIId75WpuuvEi/K5mmr5ukDhAr6DQkdGzVs/T6ki8R
GG58vn4zXdbLLbphdenPj0HUzUfq+/Y3w+2PNKng4aI6VAGUik00LVQNL+W8qw1XyCtuuTTaYJWM
kqVOXe3q5y0qppK1Uxc/uCw274wWfPN+7iP7GBJoOWK0MPLhrxdSAtZuv6Wo6tn6W2d1gGbFyWcN
PSDgd2yXWGxbncVeKGrhKSO0sAJmVDvhEhCGEUy8R5sBiD5IGLqXOjLUwPPpqi+z884sr3LOQfN9
V5BxQ8saEa2c4p3BH2KmhvlCAVhT3RGGpVzTOqRrnK72o8UE5ONmZUakPCmzhBbMqAt9yUTC6av8
0EpOJj//e8eBzvHPA69YHf4hF6/oP8k+bqd9nOy4vnWABkFSMSnKtXXbsjPM1aK/k+f+c6mBOVKL
XZ4XbM5het2Z3KRYHcaTKTLmNlohQ8JPDAFgC6wCWE2pBPctMuWAaruzP7PFTReAJ9/T5CcjCk/r
C7+WQquPUTPEJ7msa2VO0tbvFmjSTeBze1Y8JpXOJhITWU5l/7lv+6e5kS7YpC1hsbmNDmLD9oV2
dT8KSyJBe8C3EuYDVXiROQiOWEdmhHNjMDVH9xCpmDZELGSod/ro7N7Fh8Sui7zpxifa8LB5cpn+
rrQ/ohjsNsU1p0JJ9cdimF7tcBpDpfNA9ffI1P/gyJuQBvh9/NMCWJXu3LZdI3fv8/PLbXRLkxUh
C8rv5lOZgNpe61C13sctOeWgLHBX3gl1MahHUEgeFaVi5MsV0DWqfUwVd58L+ui4CbjL6D4UzrKY
GzjBmw3+rI+iqqDXvCLkQxE4AzeR4siUAAphseVwInRDp726JbpP8sYkoFqJdQxqnAHi/S45L5zD
b8xPJc5/+5q1yky378kvqhVGzDiogkkshlMBWBKmw7ELAGnwhsLMDM1uul08z756IxxE29zzX4Mv
DEInUG0sTUKVYOwGO1evjYXvZvHCR3qGcGVwH75rY27+W32yfQMo7XiXTIPyVno/qGWyUOFmdbr7
rovPpdnhiGp+Gn5DYC7OxX93tu+hg+CBXUuJMl3Y/OPLiMqKGbfMaUOv+jqnd/04IaZ9d2hNJTr2
p6LLP/GML0XJNg8zaCwDw8MP6XEXjL7D6hG5754guSWvO0wANrpzrIEaLE4XhXh72Xq7K03Yr5s3
HDoq+FzPUdwvLdELYUe8Pc1CH8wEcDCZA7Jk6FS3bKJ/pLgzxLrAFqB4ApAggoOYmgDKgzXErunQ
6j/mEwDvJRJJnH+fYMEL8lMOnQYLo7q1JVoYLdWHXwKZ4dNFkBgFf+WMbRIukOsUZAksdn/RW6da
SCCIVFJofMoUlVoqeKGisCYYyzvvdCUvgdFCah7rc2gTAGm3cZ3NbeGWDiwl2m9H8rNteWbXWKRf
8zm2UQIxErCeUgKZuZBtNFYBl7McXGuruF1fx7Yzk+CqM1NM5cYjdycPBFu8+JZFE4gB8decLGsQ
e4phZrG6g9qzWGepmYyJkTU0l8zR7O+u/NZIGKYwF5wX8HmTXhMMArokDiKNu3WxGxeOXKB9TQcJ
mvC9dBNU4HJA003DA2ex+p/oqFgZiWysbq4q8Ww2pn7Sq9njC9OM0f9H+9lqJZ+xzeqOWQ98md2q
W95xB3K1VoTThwfJ6j2+B2q68ZiKyPoTztZpnWFzjRp64mJccS13Zh3k+BqqivmCx9WmcbboUUZK
cB8p+Ng1rPy1W4pAEJkAJdE/L/L82V4EDMZJVg94frazt/6pPdkDql+C0uBz8sUZgcCqK8pWux9D
OYHZ9K4DyhpcgQnZUA9MQSS2tvWuB09pnzMiI/jlnfpI9O11nCkZGYkpXJzzX0yoqbvOSLIqdf2/
erjh6ow/4rSiIbG7sDR2nSrbPlHsEjau9tKJwMJyCpltl9C2YHbU0eaDnSyJpUC1IOzEU4zLOWrW
iogxlDCxLThY7G5e2wYAmXcnYdaoxfXFLUTzCpfScKe1sB1CwbGVTxTQd2ZXijCVzmdEewGFvZCj
xg8GZotnSW453xD3e1WGUZ4DnpTuqepBr6eiFCICVvN27wNpKVNp3AQ+VkppWPva1zlstn/BylAF
kT2MNk2A0PWAaQsGHM2il7CRU6T/c5scqiyE3lIzrFiS8/J+Dr7qQ/+9IPAxw2Md2gpLC8kebOSN
R0r2WgHfhtmwDnBUd1jgSJl52R3Y/DesEGZbOfv4bdj/18GAUMKdtYFTa8QlYvYOoRj7ttxv+Aaw
QOKMBRK5PMp6pgamtbWqWQy+Z04LRYS5w9TyjONrLvd4rK1j0vceswTmIApLNTLoUDdjksl0bxgh
uec5bM/BlvpGhmLwsEB5loLJ3tyNwrmGX0zZCt5DW2G9MB1kPqNMnELhKAw0eIeDOMmaiuw25tXz
s2dKIZ1eMaDSu8CDU8Ov4uNV19mDKVh2uiU3rrzKrbMnUvXi/sJ58wlb6AZ83rJhx3BTBcBYTtnX
mU3cpRmt4YPzXsSROdVuSGII2fmaMaivLpcv6QOrq9uKSvXr998AfjOc5vFOWE7ydvibBRznUxEe
6PsIdKc82McHV4XN2QUfH9uy2t+UKdeQypjZanjZy6sGz0AeevWFS7QxXSoLGaqUxQHftF+sfR+a
1XHK7dEgTEF5Bn/otA0OFq968fFvF+Zs2/GkBwThMZdExqVmai5yutULjxXK9HzK7u0Vt7onspW5
+/FT0YC2yT3ABxNHskUusqGHHuIFSy3qzciY5qkegCyiCAks11T8KoEBxxB+2qJ/Mac/1UU7yXXR
JaIm/FBijIWyvdW0g78rHZ0wVUVu5Jg415xecyt6B7aj6m0vP4LeLN/1ABxD3aTrXliXoXwn7Ojp
bKoNmh62jIyfz9mc8XzUoXCvZe1LpZp4GE8yo1/6hkEUrDpItakE0CLOKC/y/L2cvrnRWo995bIE
jgmz6AZllw07Rpl20y20wpTGC/SMQIf4Pjvz+Npd0QoGR+w1UE3UjmmaulhVSYgTvrsMkAgnawM8
B8/YqewJqwlnMZ/QeiYDUorQ0bHpVoY9JLtmRdmTt9LqELPBfUJ2G+GxJvmeILmZfMhSG4KE88b3
dyRkaiTGcHOYQAc10ucZeDHuTlL8OgW9uWzsZ6J24lKT4WUDJR8iZ4LD5rlh+B2iJYAZm4cjzd7P
8SvED4lh1kj8AWuUm3H0ycWFSeuN9tEoaxwhpzQgaClkwJY8dFydeEc+mZkUwdNKgzxQW6YCSt44
KPuRKqg5l/3TnrfmMKAJxYbLEPi6BAciFD3Jok6gDR01nYuNpUMQE2F1zGwgxcUbTXkatUOU+p3+
lWNFf4ka8AAAhoqhU5yEAe0WKMgcjthGPrAnITSOH9Tl+GTiOiotsaYV+C492f01FFJx4dD/mOqU
1pnhY4mYiN02sKSyARBJboF2FiqG2YBxgSrG9c1p+97JLCcuFN2LwnZ5F6rlCXp3Bl/YgNyHHvjw
IxMhWe6qWaGK90lLSU1zPYyd0sjxAq0zv0hFwQ9fwY5iqer4hXtqCYgFkdkFqJ/W+7ctfHKPyjOl
2lDsq51FKdTOsdjOdjwFjub8matZkAPngaOhGZN7ehMQm4J0M94biuxTyYy9LezDUNX8ARN4s2xM
0vFAyRpx/UGPKlj2piUl59Y54oGwr8oB0Y/lPFy3ONOKwDJZrZD3oxLs8lKt5VujjJMqqjCuzapd
x+v7RkRWDnrmQa8m9IYestDfU2m/q4Vq6fWnGv8J08aTzL2vJmI+y2SjcdH+NsiQcg1ZmCp/j5jl
HdbJ5fmSfaO+xd3pSWwBEitJP3b0dzSMvmRdKT/col2hj+vMxHOSG9cqDJvHEYE3uMuv7Hvnq/b/
YiQczhbSGLV5zcxiS1uNo3C1JqVpkv3s5t3Q7tyHF+7+XjhbU5BhfVA3AJ3slONqIgyYq0AWGUEB
zeF4dIjONLG8LpAGKtKg0U1LlThzqWLnAf6q4Qn9TDUfCEKpEb772hP+WmpQrpJne7q726JI5OcQ
+oG34BvWeG5QhmZos8TBOINhuv4Fh0u9L3ww/h0C7RzvwfwCHFmuuEwCWz5tXb2vZgwOGD0wSANO
BVS/yjfi1lUpUo3bPIuhWIeth4B0txdA/hHCuSDsqIIw8oFYO0PAdLVFVTSPTLcx7y0OrP+RS1bw
Q+iqxRNpvGyssfy73/qx6jkyyCyZ4jN7eWPOv9sffP2W+yTgohqkzmypNwgwuxW0v9+WwFLy7fnh
ZimWWXauia6X+h45U/5th9AWU6QWEc/fttRoLADZTLy60ddlG1KK9/I/RudHt5CLetJfuIqfUPJo
W3Yz1NB6Ch/7FW3te33Aa5qQzi0MM+IPNlkUAU+rO5M3kcGKtoAt0BF6VKpWOlpjFCCYnb9nxYI+
hmUOyNyNW0jvnhByWmtn7O9mUo8CyWblRk+Kv+kmZlrSdhLIwzTcdPEYdbiiOXBensDVHR7riajf
CLAHuhPupKuFGkCQv/1oli99JG5lRlDrb5rMmd6j+lWLhpdFJFiku7U1B3adQP1Zm/OZ0VMwp3L7
O3E/j79IOdDyOWT20NKb4KsCaoVZ6KrGwEjVGBnTPnLSLCS2w76BJYbURq4Pf/Jb8xj19WNWfhnB
Nb2DgNVxECuztqhkkqCM+t7YVlkbqaJRGZBmTsNt2Ei+jwzd+PDdbsADdu+Zmvxeepj+CBQj08XJ
I5QamhA6YJz2sDDAbVJjRXReIc6ntC3MVOeGOQwR/nb79Mco/Maps2nXo+BvbGY5wsP9ChdfSOIE
1iwgpzRL+9QrWOi8kZapGSIale5i7oiyvtHNoI95qbRotFRp352lru1GNvMYEKITTjVhkxNUky80
wBjDP+gPZM4ylKwXjLEUua0AgdUlmA8UonpmxMwySdQHYXLUIi9Eyc24lWr+lkdr3s4zE960QK6u
im/IDiwBD/1jlfdelK6MUUfi9K+oyRNQdb7I9X9iPEYYncqXKyqhE9qSFoBvX4oX+QY346TihzYp
yunSQzSfFoT5AEcD02MznJscjtmefeGZXyy+UCET+zSaVnMkXTFW8XwBk+IjNaVJ4aL0AnOIWNCE
9bjzC1JfsjqmTAuWpPj3do54nxa0LBOqOIw4hLprizFDAmPLPwZsQxNc2r695c6RQuOfvn9o2RO2
hZw3seGM+dAH8THMiHhnIQF7ITVpHVRDmcGKvthVg/pPjNOZFdL8W/+xBaEHj3xceIq/B8EXVTZK
VSPBXTpZqosAVJgWir0pyOegI2vP5KJmwST3ZYTqmvmpmGdZF+pVtrhowHRMDNsVRjUCBOPW0uVm
KUnOtsK9b37Y7Q6mB4MzZYobXiyffmKkriV/HQV0EMM+se2NXDqWqLh3yU2uvdgiTb+CLL8spB6I
DT4mfA7pR8bLVSbBhgVp7gJs2N9DAOEAI/+TnWFt7qteVjgp3ph20Vojj+NFIYO6g9E2COE8TMMU
cWqhDuzKgI37CwFW2ga8a9MYMxxD3mf8M+q5gZJixTbPNTl/4egP2bVvNYHe+yQTzmcjxbDmT6FC
nQoxcIkTKFQZZ+VFILrIwMXpMfxZ7b7mXC4QUB0WHbMkG1lprbX13eMZl0CaqRMb0PK+jJVP2XB/
wK9SaRqn3iZemHBRBZMmvhKl0skgp8vPysUDiFLg7pbZOH41CJUiuZkwCj3hIlMlurzjkN11562X
2A43DeSQS5nHBQlL8yWiqaG/iGYUXQifOzk7/XJHMutP/q6DTS7avVt1M+SF8/VeUGNkuNeNHX6/
1kmlkL7ulbjIVq8n80T+bg5kV0GD+UNwEKE4Avao5hgheSC4UZEovQ4QjgDJFwEotmo5pV721l7P
98A5MMLSFogCfOEIfO/s0dDqwR9WvR072FcyiqB46TkTOzKtTb0rQEpYnsRMMv64tx7lKK6n+ZmM
zefVzLHCO1qiv5V8YDaUGKWE2u+ks1yuOd0GZgf8oU+EYOkSnPHjrboJjb2Sof1F+yTbhs+AcjQ9
dQ3pZJTw3GJWxlKQV/Ch03ZvCJ0YVxp9YRZL3TGzQM7/jMv39WQFCc01ZzAx19Xl5Nms4+vbtZBR
YQiLOVi3Ta5I8CGVMOfMGLKWRhJNLRqm5sg3tQYJmLcnTlmACpx8KHkibq4uQrj3ogdtvyoCZvdG
z514noHSNpQ3z0JXPOLpUKRyUr8Uf/XLIJV4rQ7AXHeMpH9+c1yoldVcbxRZK2zTxtcW7cM/lkxs
pZ4PS7igaVEU/RfRhY8egCoVAODMCHXpGbMoiFtiYUdtUvs5Bp8FnwiCavsmMD5RTp6myD4KXOoE
GWx5R09aLSXMl8iVbnlxFY7wLGvuiCPfSKVrg+6QmEUR72EymyCxMwSG+j/b/FFc6Cgs07aeS1YB
XmmPbtBoN61v7ezlxshTMU1G7HR0cxp/TQuChmnE+z+GDx8vEBmx5x8+6qVPhEVP8JZEfMS/TCVi
MvL5j0MhNQSG5Ycd9fx8ODhFi4ctB5JZEfiE6itA1FAMSIac9egkPRglgHQAHqlyUMzL4DBNzVFZ
IGmMBjk3hB8OdE/am3KLC3glc+CRSN73rPujuexOt0uCqWyNd8MrX20SCzuZc0C1ZSHrAgf23ZtC
O5uFwwxGEDQG+oFKKLopwtHt8/ihQkchrUwlOscARvGA3d4Pfx1sdIAqwgtM/DLQ/O3Vo41RUI6o
iXg8gXaClxhdwcCmSv4MH8DDvqCOAW7YPaw7VlNpwstMqn3IL5HsI3QXtMD5JkTLQMwUj4eho4ji
OjYsCpg8lsyy6vmNnqsxx1jRnb99BbmOle7OLCqvmlpjD46UtpyUHfRVT/AhXXS91MU14o/xki8e
b82gY/tK/+KlTM1U1fwxhbuLetQpX6eEg8j+k4mOGDyV9w1kECYC4Sb+teLNpXc1USM3Jm+qyX/L
jc8hnvdeDDfNgZQva78kHMq+C0HsVVZmNKiIMjKUDKdcT3/alwVYPXLSUWrx0KlMica81cdo466k
8iJ4dLWVF+glwM+z8iDd5A+y4qNhHnreOJtO4Z/s1rCcP81Hu26p0idrcZhE93I/Vuo0/rbdW+KB
laQOxMpOt1TfwSKLSAtXyrIslsSqJ40TjISlGRDiArp4BhSDdZIiu7/rsB4ZFDbfRHMhzq0GtLYn
o7TnTHE3uSaUjxvlNIyfjQF0+dgTRY6d9nkRBPVujfinhK1jB9wKxhMYhV+G/oJ0xWA1sJyKEbJc
u5RNXofIwXqP97Nop12yljEf2HCSHUXFmZL//LZ10xNojqPzrX6KFimV0w4ZmTkh8eDoYUgJ1qlK
eJslaTFPmIVkigi8FqM41BD7XJPIFDaKv3vlDig5pS2igYIWCK5qZ1LY2IJzHFqXjSUF3B2lWwTY
x0hqoLupZXSzhS5NNZdCF+OtLt/8QOXa2wo3mz7551k9w57L4ccjgLF0ewOdXmmH6H0HvMV/RBwh
kcu6vtyWk0NcR5Wr8UxZl06BEKNyIhkvl8WwTGByWqLh6fiGYzS0lqrMQUhh7s0r6kAsqswlwGfd
9A1HSXfjC4n4EwexO+pKqbgk4axfyRSJsr3jX0XwSFCOgcvn/VvbElFyv+XYNm2xDsM1xBt/6tRW
+g0g3P43v2JewZ7LhoSuyDUcjzkW8/aOQochX9ppFw2arcnS7JH6NyzRX4sxyeBsxRix8kTHyNOW
sZFzq0YEeiD9HV4O43EzefV/fgzLlAlhmphs4yuZ9vGd0D+xr4WFL2ZDPNBFg2RRDbKhQjNEipN0
nCUgbTU6aoz48z1MT53PtrOHo47iCza+Ja5fNDxqkT8D87WMbwf0IlMZKUyZ0uaVy3NjGw6aOl8W
R1OGRgu2YgxWng5oxbB6eppfrIu2Ti+buYvdWeB5AZUhsa7fyFTqFwD37R+QTlm628vFybsNLGC3
qZhm70AMqnkoDWSCc5Y5+rhhW+dcckQwwQ8WazkMEQuvQvDXw7MVR3oAIpnclWuvFzeaouxiDhjd
VhCsGw2j/R7ZcAcTHOVGzuBAEqhIUaZ78X81zYTr7BnxixzDf7znhRcje1HqO4xbFi9fCnUudDqb
tOZSG4fuopi+nkMwNMutnn/N5/TovzpkBioIPeKVVtoE2dS3z1QKXB+TLTMZ7qKcE9/QFdgMPZXt
bgIRtaSNGlZV2FOq/+Sj7a7ZIgPWA8TnKI26seHYw0aktlz++TB6FvflBQHw7SpmlqG9VrA9BUc8
NiHbSf5Pp0xPBS0jY0lB5R5+jIe0k8zjRoKoJsilRcS3TsRP6otAlJ+OAzMOaxVgiqgFiS6QK4eu
Fp1+Mq/s3GV+kUZRz2WcDRLnml0e9qRxX0vbM1rXJuL39gZWUBYwdYv4bKUfFkox+9qYfqn8/e0D
m+xTKx1IlP5O157DKTEK+NLmyPbX15QKwW2i17LyFEHzOtg71i6BwSU4jTJWq623zA0AhZF/Pon2
vvvCz5wYGRVrZ+K3D/aGlktH+bDY6Un9h9LCpiXzRSPiErbXH8pNj9+ipvkWmjV7eFG30ZpjvNhf
Swbo63SwwiDOdhsS3jJEYhYjVaMjmEr41gSyvFI7MmB+leKWXEc8xQEcaCT24GCbZrUu6pyvnmIp
N+0IUaj6KxFovOsWcCXD8HIwVEt8TfE2T8XDFFcISe0UJsPc3cgiHAMKsrNRNjeReuHVu6c3QjQT
5WuChJbVg2UWbdOhgdtRJV77uZ6MExh9iSzb+5lwcCYNVLpMmGN6kXSyeKs2Qdudh9GaxqhI+EaW
V6qsLdWDw6QxbJLI2n2mfjU+lJJnY4kfR3SKryZAAsZwap6/C4bWomrA0xK7iVzhEet/DPro0Kzm
edWd52b4qsu1uYaWxPtKrmLdWw3deWRMNSJ5NHLoIhGHfG6ZeM2+d6gYyXkwe3QWYKslqR+rlHrO
ZVmLt9YBsZk7IBXxMCJ3rIu9JJz3gVD79IOVJ6AGwjKcWBHnUgOTstNioEa9QI2D2Hkq8NIxOGUV
l43laCD/TLtKhTAaFbukVOroK3Fibvhlp5W2voh59geVN+0xz9LFDLjvI1kceqetyIxVH4YKjmHF
30hkF96SvVgNNcEdXMooPZtfzWl9M/SJgK3rGKxNstBuVH/t5MBX5lLWmfonOKJjSIW+Ck/j6SRQ
qaDayp9r8zHw4nG6chl2sHVs8ONIvKR18z1ykTrHRMY0TgeprDDu5/IHccV0w6wNz1FIxubl3not
koFaLX7xw6SyscX4W5ihivI7OSd3I2Vu0It04wGHJrrWFQS+P2ZXyyRlb2IxBezpgVFc3x9af5Uc
Hpcjdm/QVf/XoNzZpRrqZy7m/SIpCtoElREDV5eddEXLtafSLvCGRmvsjg/HBSX9TPRCeU2MqDpz
DjFqFbeHBby9bDlXkpxkx8t4CaA/YvHkwNKhxvANyIAZu3l9O8kDoj78Jm2EV8xOXOp0k3G4ro1L
8NZImMWN6U8pp3fhgzHBnDXt/+LbGheUwGoA32ymis1CnNwYZhMFHjcdafhExD/22vieZlKTtGze
OL5LPPcs9RxP1joMs3CaiCznzwrp526LvVzigvO8rCbWs/FXu4JXG1OZjBmFC8kjRU3qKQVVlebX
GADI1v+80ACOfF1P5V6NSqmu6CTZ63+NEVgBzdkuTcL35JqEzPDNGInVVsvDECSJJUCcr09Y3LhJ
uESCbPlSgxIWvlp6NJpBrWGT1KBSRQPP9JFE9F6ENHsljxkZCXB577EFZHjAjqBxzedzDst9nFuU
9l9lxQ15ozrb/1I01316/Q4tx9kqxNOQIt4/dMng/8VSTxgi7waP4Gc1MFdL/kc2s6lPVkKMhgC+
NvQpN6Oa5UqkAjiT9B/dvsaeNb2PiyqtjddYycL//Uyu55u0hLXrvzkumA/Vxk5EDDhwy+cmz/qp
CFL8/IAAevznpqze1qABteODV5C6MsLyZCkOrN5ywlcXofDEfuFYTEf6XHVCzkag+qsxSFJezXFE
yEfY3GF/JLrixcilcTjkq1y3q9mHeTNY2hfznePkbj07Yf14Bw7FS3a8ykM3t4RxvgNSYbit3ZDp
4hhp06cZNDNxLnYLPMICfbo2SVuXCbrkhcCZdGoR/Exm34o+QYeqauvOAh188X/plxREM4p7ombg
eR+P5YX9q4LgcAK3a+2OHwlkN9vhXb/qUoitp9aAojUqA7jZLmgYBqHvd3qRz/iyO2aBVb7Z9eZL
mpzpRvCayuJPhzTIHIcqnund5l1SC2jmlyf4fiUbeneaLiIGF2qz5enHH/KPN5oBnIppmdCe3waQ
YpJA1T2O71OHV9hyFH76JehVWHGIDt1o95kmm+vgcBfHJCFlTPp3NOFL7mbC17mZy8/ouvNoE4gl
xjssUTloQVHD0+PsW+htw3P2X2+hdPFk5XBOQag9ox8UD06CmgP+mWQ2n/+2sSW2Nc48Q+vmONwm
EQtUjlwpCa8xdzg09GBWrjsLdtcvBVn/pKcyv5qLWm7R2MLF6RdJeOX5XEJ9l8V+7k7qaOuqCyy2
6R6n+l+/D7aDhPX2PuRCkY81xaE0xAuIK/ZRXQmfUhOGy+Djjc+j8MUUf+jyb19bzHoqXFaY2QxE
nEhXRLVuDGu+aw7y6fpaVJorBwPHjxtK1scTXOS9XtmEqKj2CueRN3qVhC414EeVQ9j28njP3TLU
X4TKQcacBrRiM/kfolGcxNuDOiUpgNs+6dUOZdrESORboK7UBkQEvNkOYKijkAyLb8B4D6sGLNni
NYoOZ9CmbjL1ZLlJqp1ZDGfW4ozTPj10ygcB1mmthtccvs7gYwfqicE30KNt8A+LT0bgR6RO8Drd
GKHQqj2mQYZGDJJuYl9TG2/zV93RL09zUWAYR44n+Bho4t8Sow0z2smfIQ6U+y5hJj/Kgjs0Z9Fp
xXnDlr1BYoTkdGsGh3JDGqput7yJf+CWF/RTJVbRrc81FwSMzEzhEm4zRIHGv0Vd3FFdX6M7x68F
akhe2j0pCeI1oi/MSEUHmvoSHRpKRP3ATuxBMwb52xsGzTTL5PU0xe3ohgFoK5Z6K7UuHI6/sXsd
td+N/K5orJeNGRUElk4EOyLzFMgMv1EWOZ1KEosaYv1vAi2RnRKnWG0TR+Bxg1ZZCXxASA+PaDub
5rMBh6iTvoStkVoCFHyXWv3Ct5FjDnrCqK6JRYEKN1eMMF+Tf7Khy5pCQVAA6/AuHkHN8uDmWEMr
iyRZIarJ0LC1HXsHzPl5d0nURA76E9VNDPqNrr2K252+9Ataf312/odEBZseIxPaeQzheiiCLbg4
IaI8gU9TfVXywUYF7UQDxsmPsI6JscC9IT5+qPw/soAYo01d2Ahjxw9m+uuevw2vJjji9d+Id2jj
arhIl/e1MTNBjxD0QU6JxvLn4r/pqhJvNpwWw5SYN9KgpcfBnx3Ibq6Mw8JzONBeu2j7xssUWXiZ
PUrGnZ5ZZZr6MP6DIV2UD/wUjvLlzEzkVH3Au8mURb0vcsKkAH9e9jN90av844xKo7HdDV4HcoVj
PDqAKzdaIjH7hN9Zr5P5zsIda3PrnhAj1925cGwiBHxr+7l3HhrzuXdpmg2TqBMfeaij5EsviQTq
5mXy/PhED38a5GMLak9anPnpCXvRnL7AK5pkpf/0q8qWO82cSxmkNIeI1hvY/hi8Ug3SS590obfH
UrqiV1ve5l9dxfA8Y8DZ9uXqJKyjRRdAUyI0sFr0nCQkFY2sfO45+x1iWLgb8/D2IRowVQZPUsLF
uuKR6gYMIWCYI8UKvbHpM6MycAUjYWWUzoi0LtKzGay+9e5IGnIdJzZuKt69RTjkMpgi9QFNHERa
6nNBPzmpPe0QemxdhFj8nFAMNapIi2jJ9SH9l15EVEqJaWxsEDDgGXCqhqM3Jekt6/0/omNhe88F
SV2yqkURonGOflIc+5w2hCRI/0lc+2V2YJWfmvf8lNPPY4Ce9o43KcoliUru02sUy9vB7jjHayAp
XnMRKXS6w52zjPZrb8WzVCUFhUpnwf4izGfbOrj9TCjzBKzW9es0nmZyDOhH98esfEMvrSGxLTbp
M2SB1qjb+0qQZySmvU0cEcDFw0ihq3QGgFS/HQ1BWkyLz2NUtP2jZwXKfW6XZl4QsRzOKA5dz46s
Xbmm05TFHTBrfzxuDFO++a4Exa89jyCktx/WoLsywncI2V49SJYbztTVZYK/WT0xDSkqLITn7onO
fMd0PGgWrixGptjB/NZ/hICfWrdx+mBiTQXijFIUIbzOyXfcyGCnaOqmGE22pwLoUpFq4Qm1Y00l
qsBQykqCmwvXoxh0moEnbDL6j3uHhuS5mOhu76iwUCED72YQvf7zPWHAs06YJzMsoxWMFhjq/YlS
as8XwfVuRRvc9qEjmKD9d/Zjx+Kgk0HWAZggYCxTDZilQmRpZeN2xPOObVtvV3yNSZ3a8h28jyie
xsB5TqQqqS+etn9B1bXep9doFNFBR4rT4PGgDlEZxZ6gSst7osr8aU1DdQdKREy8kO0zdLmxk8Ur
Ey3ZzZMCylfFWdK1Bd8Ib/G/gkHnsnCynQ1VU1DtuAwfpf2R94GKhB/6BbuY4tDhnqjIm+TQOS70
tGpp1KQDg+OzYE9lyOhzFP8Mq5x3PufXuTSuOIZkLUYjo6XvkyNnoXCZPr5n8959UG6AEDlj747P
7BaSHoYXtlouMytx/YJdRmhlBzOhVXCaKDY550Ckw3ta7lW0MYRvy116mDjWsgzR1wBpiMohsoCI
KhgiKT0Sv4n9xYRSr/vLuT2WIlOuh51EuRIwAIkUG3dOwzFsscxFQwh8ERBYxzBxaC0iBKKqSg0+
2hEdRAssgOl/0ygzBEYzddC18/EOGIrnrHKx0cx4W0kPR3p1G8vZK8dcGtuXD7CzYwu13smT1LK1
BoiDO8DOBcJ0ixHzd1vwxtaaWMcbO5n8vI7v2ZUFSNbpIV0jyE/j580WceQW1HCU+XEXOkPNmG9N
i4kEV85kZDUNnhpi77khmL69TZS3LXkaHn7V+SrtRcfPpR/VXH00115jLHsrKrF+7oiBJQhvL2jj
n/6TJjwaDJNsacDL/v79AgTrWNT4t4kfGb88hLOq9DG8TpsIjNT6Kz93QH9jYTqUcrzPH+C8HDmF
s3194N3IV04SE0o4VlbnTQr853fnhQNivH0u5HoEbiigFDKD5xC6WkExt6sDJ648X9hKeNx0hpt8
LeeH1eXyTmU5kfvflMzqcx2sHSg8puJeg7ArZoKDcDqfe0RB9/RCAxsAu07iOkrBI8uxMd115u5J
tqqlInk9ooCUwoAT4xXoYC8AVd2dog0jkqEJUJ68InFnKUgRfXku1/ersGFV50vhKI1OADJrTfMt
K97CAba8pSzXnlSEOWkC++SIxhEUWU3l5HJJdyWD1na4qymuAx6F376A8Tru1uIAK256ko9sA9qW
U1wz5ewo7Z2PXUPeL2OZf5mvkfLezB08m4s85UaBJZfavUEgmgv3o3tJ9mfCCaDiHsJ9SpoA5ruE
TW6jXpXbGoLx1akJ6TFMIFaYhtnYQTGO/Ors3Hs2SinUd+lrBoyR/WeE81mHbMwC71/DO2ce5hCM
9eIYC8z7yECHyq0q3WQTMqOm2tAb8D39uhtCBiRHMvlGs6o6y129LHvC008hLUPyeeQNL4PWsaXs
A8kWpeVU6Hh27znBqInPeXF7Lcqo0vdD9tJ5+A6q7fUs6zjMOHfKPZQW72nCrIgEwPB+pB0LDtPo
2R+7qWyunFx/z/XlVQ1cWBqt+nDVkS1zwLMgkGc7YtO/lTOaU7itGd9fm1d/HUyjaZ44QHgkvdtr
6jcQakeiVIreEmYS8bzNjOsMb9ybASc6OiXCMNdIFlMEA+umYMxrIKK5HEFBIvbuM6aeBPv+jjFs
kzuBPRPbipNM1pzXup+a4XBnn/8n3+yipAM7rmICVUDNm6TFKKyonj598b6bMMQoABl1TTkUAsJC
DYfyH7/N1mbrSwHrgVKadvtDYLds1hgwWj5kwCkmzkv8PO5aY1Fyk87Ut0YfnOvfR+MoiaSkSIIC
rDUFH/wjQT3VE7y3qfp6ZGNeqLXfELs76RDN6PxkAJaAHtKt+wNolOB7hRsUAzT7KWyNyqQgda7c
6jBjEF61PVmEh6lKlar4+Mc6yI6ARj61W/cc/MghZoCACzHIl5SQ/cgCg9LWyctKD+9AC8/PB31m
MmU8rrV6doAqIUMFI5dwkYgwE+KXhVqPMWcfdqRBWYdJTfrN7ZH/vgEyk9BExfLjtqBSH8L+Ia5y
SKBNN8s+UY6wU32I94xmincCyRn4MxjCyK8a//Trwh5wib/s4lS7+X7ct078Zt/5qrQEI09Q1sD+
7LA+8hX2lYV/z2uMtAcVJTYtWo9hKTdnJ6cbPGypw4vrOUGRz9gpekCYGnqz+vKk5cv6NPlzYYnj
w50p7CjkD6LY/E2e3TpEU5pvyaQnP3h81lNd070IeTp1CjyuCdgN+3fdo/pjc5QoG5FaJFC9inNS
7U8xvLNvuqL1Gs9YGjNC7MkbU21PMpT1dXCBxWlCiyPaDsTuYo9jcTfX193SR+tllYZbvvdI5SZR
LcUnxzb30olfT/rJWsYabIDRU2U+Z0mSVkyojT31bzCHIpHLE4eL9ECJ0gaH85M/7qKI5EMOx7Be
wRATlWHD5EiC4Gn0Qx70xeSU+qeHTFeoqvLS5+hHhCP7wFl/z26p7l88eBYQc6FZ5JfJ2DA9t2VI
fUhwQ9Q+4XYLT7AA2jQn2rYOAm5nXWwqV5YrlRPBjj1Iy5v/DcWV7QMBW/ueP3l0FZ3TjqMaud6J
jFSq+ztf+UcKZmNeWNIF9OBunwu7lqW+2pimwSkCirU2NLT8ppDSL60J8r7Bu1UtA6590maQyyd1
93pv1hI2SquSQLkDn6TyMlnOX+uNqJNC18reCtXcNHODlgWaw2RAT9M5igjopn2OT4BdaxtAi52d
TXomLNEWyhdAH3wcMEfre1/6e+cRQkF0S92J5YTdrYj4McHAxgUXCF8A6eWnEHlXDW1woMCaXZyL
wdOTPIOU+wdFH2drH+Jga3mstoMFJJ2O4IBiR0xHYmPjH7bXMDkEKyPAreyMKfccvjnflS2Ia9ua
JPyl/559W/twUbeVoZGhbd//yn1QZ5ECHQRD8qf2UAAOhTmCJTWoeHefgLudd7xEJZpPsGXc76qq
hPF61VXea8CRVhOokRzPB7E7fDIDa0vEJnUXXfY5BaoFL3CUG36PmE7itix6M4rHSiFycgnRLwB8
Abj9zyharAiTAvyRGgQdxgN/vrnNTxxGr7zCZG6buy5zm/SS13oQDRtnekMMTgQUlYmLTeXz0EwX
o1RZGzfPmE6RSz5GwvqxuQrLYLq2FLG0ziJRyjCxCy0F4fm22RqFPPkoGan/TZ1Oj9b9jL+nuYsf
URVPDFWBi1jNCMKKXqDJJj4/TlJ7XEwx6cspVSxMcUvRx2TBglgvmSEZlWkpYi7DC+jSi7eW3Smv
Sugn44/XyfQa0I+NM1yZecEzvQqJq1iCmqr9U8CAjhruWAL0Zbi4lzb6k5E/XBuA/16tEW9vmgnM
P8yrMcDzIXnhqKF1+fmyhgVITbvkuSpzrNtR15zOf/CJ6aris2PTYYOXXW191eZOTjF8jDuVgEfG
piC5XTISqYcmS5cm/fidePuVbd4mcN4bpmP/3i+LBpcRybgVBvZ7HhlvSK6jZEoMUbr5R5XBHamv
BmI5Cu+OQHAu8DlbL8uQbi+R5IDo3UfrnXfZKrMe/MQXF7pmveEnLd4W7RVD8LAdrikaIEuidWIL
v/d8nHtWbVz2fD9jvibFjk25aQKieHLY5C/jiR7WbuAFmcdtbd0UgNWlrr9j1HDXhs023IpdRED4
MshZ0u8R9ImH9wdYjdP17fLWvh6rR4dAENvIJwxzmb7eXej7D5ChW2Qd5gEJ6VkZlQiSS9IvjnI1
ZMpzEusvZFVnyNu9kgbnU391ujYDU2aq5sizwHjfmbTI2dsoYIHyq0hWnCUwW9CFawf0Ujlyexpm
QixQlJKp7qF3rHOp55wJZNfUkRlxzuaRwmzEAnGgtrXCvT5mFs1boyUJBd2tLBc7bJE5jKT4DMSd
l7U9Z3vsLSkhHNGIFIrvbVAxoixkHX9kd4OanXZO3acr7NSq0Hci3NEONkYFOkucwfB9CJJ1qjXp
5zuZzLdH887EU/8u6CdrPfz5Uv7mQbOe3DZsBvdbvTM7Un7tValsHCvOsh/hguADnKYv8jQAq6h5
y+B0aVh5Gxe05TrH7i5ROHZwoI+ZKqTb9kSOX+E29oI9XBPfwVCSKR76G8y5vO5rNpLeT/rr05yV
O88R0BXQ+z7NYzbr1sL4NrEJgio0fIbgTlg43o2p3WLBBPl5khx4EiaetVHYc7zIvGdzeuCEYg8P
YkOmh0X6htmHalxvNmkCDiqPOTQgLRC/DjOT8Tl6bNqEcobqHvKgA145gCIIvoPM/iiployLMwv9
XqA53cX5IsgkzKdq+hq+r63MDbVPLRnGGZqD9Tszk5jDBPRXR07/HSRv92FkN8chsXMfzoVZRN4m
A4X8fggf/hTREKlPEMd99i5nk/JKDNLbkkfT8VPFTKCJMvAvgnmDHdCkHvuI5tuDKkNZuAUeiXVE
R0VbFS/4Bd15dYbPcV2kNuvOQujr3NKL7HBVJdGND5pMA2kDJADDCjq8Qbb1TxzVGp/09PhqRTVK
6ajREIB/+TtJlpIpqmEYYCFOKx6L7nHV7ogkdkqyy/k6IATkU5qBJbUUNlYUglD6tLXj7yuD80E0
RQfDw5boM8Eg/0vO6ZJyY+hv7bTOGV9G6OCrFWhZGhDexZPidLL+TeEKPJRU7qKWrs9hpl2nETkq
tdltWX5hUlMBHij6e6KDaM4WhFJk96dYPYDeLo0xLgL6xcUynrgzsXDsPl9um4x/gSe/RhywpyLr
jVyr4IWiJ+ETKrAsm1LMOZ/2l3dnAEVDK6kQNybMfj1PqPXjDHcWcIyiCw/zynwbYUBV5vMMaQq4
t/2WwHAuRsx/5SHXO2dH+6pDdSFIsod6lYpw9rvS/0gFcGXHR96EX74UmTSGJAUCzZg2Lk54WrfD
QGO9z5KMgNmmHQo47EO7iFH0L4ZHTt2+chq0K6/Ae1Mbv10QDCoJ1Q5XdMKgXfcVBGLa09QZCSYt
Ftnb9OKm+Qtp3F+I+l3ad3CzGt58/8LxUXwtUTEPUU2iKQs78To5dgjcvStkJcPfGcIyVBoEFlHh
S+SvUcJQKTG1lThkOsbMPRAaSFIHmhZ9ac1LE4N4GZs/7y6a1+x3HtNULA+jrKrdYUsAlqumw0QV
5uW13AYv/bDwYJu+p6EoVGHwgK3SdLRBfG/dmHk8K6QWf6l+jQI5KI5TJvc/pSJdskS4cdHfrMkX
IEO9N7/33Wvok0LLzBnmDgMTT7+mik2IzvDOoAnJ5fZGC88SrJGBzGYtiVy00wZAaGejpV4K6aJm
Sr8XkZI9ZY62N+qnKDBjcqhvJOmQbOdGOVhfRUB9PCOoXeZpU+WF8ZeIt1dAyn2nQrWNYK6y2lCG
mWD/2OW60KTedRF/8Srz+6LzjlRuwCqWS3PVxMTKNXdlJkFPWg+esEMhCz5MzTzfKCuGOnQ15mst
libfa05uV60x6DCobRC532rDBJiRWrcNuVKcj+IcFj7psULqoMU6mnDKUf6Gthf5RAKa3u7MutWR
ILElzjm95MPKRvlD1Bh36uDEBrweKaCFG2W9+OgASDlA2/TeNnkBckIpDffqvsvKHVyU9uWbzzIR
rn5Um825ZXaZzR5g9xacQL/nur6qPFPg4jSKf63g2/Bo9R+zJ2yZFcLcqF7Sd7bmcmMgwmVxeQg1
FRvvehkmTn0u55tjE4jS/kYJoRDFbgpH3PYCENsdf04KF4Q7Blek75B6YY5Uv2HXZdXK9J23Ir0J
Bdp93UGzuv8cY/xbRXuU+KjCulxkj1QjGYBECnXkANMCzztQJSTnhKpSSYJvOvdzzXtDJT01HeuR
Tt0iQrINt7izlWdSWpC0UKrezXiuSqDrapYCQd9kxFqrDckOq4TxscBoIwZveLE0Pu1TikaPhgfN
0xLQNNa9o9Dwzacou3QnDYVRzMwbXFJXKexaquj8w3Yykfi1rgI7+FvBzPRrj0XR6EgLFyJEmyLe
RZgv+ggd6ZOcDRCxx9y5w4N6lmoMkNfYMfDrj/Cx3ReX+GppYgIX1e1twAvaQ47D0IuYeKKStN4G
6lkG7CXMZgyKGV2g3OZya2vrl2BJqHv2OGkE6WlbtBL9axALS4g+FLvxLX84h3RDkyACdQGCclhg
5reS0/5g+EXQq2E4IZ8CwKDneVetOa1oeu8LzeXQkbpz5KPXhIr3ggKN6itJ+wopr2n5U5S2K1ez
WTzqeyEr3djDWLfSOFlNCxjzsTlouJwD/R9F1v97OMMBGPpoYJEAyXUDMqR/eb+OLBPRHXRDt/Mr
6PWAmvxgk7qxmMS/OoDkELWDZ7M/supMdgqJjjHoa5P6KxgSp/hGBadZQtcVgLq4SKAzkNlQ5iwJ
CpKBhVCw+6eRXUXQN33xja1YtFQRREVXfXqd8QUhh7vPq/mekjhczspeg556v9H/b70oWgI9hq9O
zAo0BbUzwORktETZnp9o2MK3/X8sbQP6XKUfzQx8yOgFeLWDplZ8EKfwuF+OR4WS7a5PbDSirDHZ
1YrxrIkFWLSiVc1DC8Y8x3FoC7yZvdcL2SdPyTMJlYcMOiEZ1ZLnRKEdNpHMtBDUEwTJ8dq2R+jX
Dd1ivQTTsCCjtscx8CK+VWw6lPVgWOVyvjYjYgJE0cGq1mpx/pvvODVfXV8OMKy6GNoXg2IsNlIB
azEosow/y/RoeOHpOZ/UDp5YXfclBdL/ysZ7n9RUp8WlJAwxRvx51bNTsITA80UwxIv4QmrCqc5U
8YSdFLhFcZ3m0AyoD0Ff+xQnOv42GG4VJX0mx4nwg0OCMqzqOtyjiO1bRB0WvhkCogvImsv2Ylxr
i4i/s0QKiK+t5X8UPOaveqrGUXNSjgiR2idFzcW6kuN7Pv1l3WKKZE2uRtBNy8vnYX2hF1COCt+e
UbLrQyu021ce6scIx0Rb3r8w/PA1N6Skn52+yW8DK3+o94akkm5qTOt1eYgkrlTxUU5wmwlC3ZGb
nT0kPRIva82cua58bh8IGLBY2UDS8OuF9u6s6eUVOK2UPJJKjpczgSS0eFsHxsMWjKi1Sf9IGONR
8umMMDyPFV4xpvRtaX7EOmcD+ugOVRo8bDzp+JZZ5VldSP9TYHLz4YiB4gcZ3Ztcldu9IJyRv/sV
mH713O+r3juQeCVLwHPYTOwcLjY7JGUGGMwm7urf+MLeLLFA5iyo2nA8rAy5+dbuxhoRjxAPoJQh
K4Fp6RL0zodTARx7JpDO8DzTJMjY9IgRAxvrspPkTGGHxuNFsFEZ4PuzfHygi7rebimCqp9NsFMg
xuZsD5sw6QQLZljijvbZ99p/zH4asPQP6g1q9ifLjnZDCtuWqUQIgIDOIpAG8Ko9zCWMhBMPMH4D
i9x2XZqywPaCEtDLuAQu+z89vqkDRhYZfmCUuypJ36vCMo0CZnA34mxnJ+EycH+0uHRzenorjTMo
o4fhrbjEXFcW8O02+K1WPlztfy9orCz9OcgzDceT/RGAimFuyXWrSFMQ43ZL6GSQPn4ve5wZKK04
QgHxvrNHo4FYDTyAQqKaIPtQ2tBYYgwjkAHzk5mE1al463bEeFwRHTAyNGkSxxCANy1pgZsYT96n
E5RD8++YXdzM1gHf5UbTlwCgXlO/kPYuDydVirnYes+YRb2WGik8Byy+Iu9AofxDQsPZlXB7V7X/
2gUsPCS2BDXnUfa996IMYGob/j3/MtKiRwS1oouoAXaR89NxnEblyslyVmisPP9cWB8zGt8/Ufu4
CaVbETdo1l+JoNwLQncZeTpyE2IW8eC5E2Gf2NNSBpz+sPcDPABA0RMaXYGnDIKQSdo0YUKX7r5s
J2vYZsr6v9Lik133iUum6hZEYu2erZ0bj7OA4nLqrcMIuwtTouCdaKH14x6jE1t5xJTQIlTPqTrl
lXVCSl76NMFeScXeOvBYtqVh+r1LmQEBYPknfMgxJyH6dj1wKTX9AYfTtPEVgFX2jtXA8U6cQ/6t
xcvSRze1PsZNExGKil4YaFgeg/Jd0prfmHR2guOQaQHJjp0av6YncA5ww0z+kBdqSQH7dAFpp+Yt
3B7hnFVCARqrXg6NNqSUxPkU7NWEaJElL/NHWydzCgWBGHwLxQvO9CFL818Fnk6r92e0pEAIuOEX
9geGK3qdh4VzpKKGuENqBSRf7qiUciwkePeDKeSKNZI+kv5GRzFULEDBCTWIPmZK/ND6GtDCKarQ
yoHJMPQV+r3+Aqq0wXieb327X+XlGl8hfMalHF69sybQypxWU9VCWAyZH8k8NLfcobYmnNCuQKCK
6ILVOWFYTseu5DGavZUBxpJSAq5NPwgYTP/yrgLhhihMZyrRdLU0N2EUQYW+kK8U1eD7IvAMY+Dm
9Kw9CwR6RS8pcj2XGy2mgG9ylWdiXxYtS2uxSXbKzjICa4bwz/2QDFHr+rM7YDZt+X01WdNBTsBh
3SkPnPFr7uKzWwar9L8Tcr2JKbA9pgrXE+Fbvc4dQk/FWVyEjF/KSkC/ipGvb9uN5N/sRJQK65+x
irf23QTUQ3ukEdamD3UBGEmHhDYj9xRiFiaNB/rHJPa84kFo6IOk4sG6+q1jjcYYCSR6+lkS3hsT
5sBPWe4FSBe57jWRjWHCodV7DrVNQPjoEc8fYPkGxtCqDV7CutuFa2HYVlmObBBh2ZZzW42CypRX
zsfKA+Zw7qsZLbjw0AfR9LhUgRaU6i1QXOcwFJ0fDny9s+wqLYC6pzNpEtGtVDe0AC6kHB14xTRo
8TC8KxnZLo8nyPRNWISAQbptQLiIxFMqU23ub8CYVgBwfhz5PpM6rr5QS+N35q7mMMyEPDZSDvfE
4940FHJHiYyLslex9OPTB53fdMciumugGc10DGBen0yHRk+YpKjvuUTnWxBCbY7Ce1V1iWKRPjTY
XxoeUksc+fI5+3S4dEFaoO8sGmgzDmrUXKjo0epUVQiYh75nQdIxA0W+byEjmnNH5Q/m+E0zvyda
1MKRAtPqTyO7VhgJAqaKjgc32pOcx9LstDiyQmMLTcMtP6KbeDh7cCbleWZ4uOAgoApfBc/1h7PR
JS5LS0yJUbYwHgEEaSeC1FRC2066xiucWjKZH4SljTFxUMbgF+HH8ejaEuc6ihfW6Yrr0ZKJFsii
lg+3HVFUqr0tkOMRuq4ycOiJp4+m2/iBnQbnG/HovFl3qFVnO3ygHfUENMxIHx6BEgj9wsvc19lc
jR9rCqEFmn/z03BVqGI7Q0Cnv2MmTjq2jBb0XCJJS21IabNocoaEHK/fgI65of3QS2/ghpHxHnrk
+A4eUj3aC0gwLfVzu8C9e3EgSQbb5IjH64ahUeVJheedARfuOgtDQBj++pwVVLhSOjlx2I5DKQS8
vfegp+Db2AoOkeWq56aboNyRX5s3vKwLQWfCwbgXVNXe5ZYOzSX0CTYadfpBbt4sJIFb1IITDNWu
yHUuPoFAT64vrnDYqpimosLdSOK5ohRDqgPqhxbmm9d/kkYnYYbktVljKBPrLuQFfVjtui23/faB
U1mzh9BI4eBqpln+66W5SfhQLns7QWsiD/B1Zw1C5cXYcWxIMqDtrOLWfuH6+J0OtPFicUeudbWq
NZcoQnXggYqrNy0eXioIga6+56q931Rm+BMkyQqcVg+mzot2Eq68XzR7SqtphyUpHKdjfGMUmCm9
3Iyb93gfVY8QeLn+XcrZsu9+piXupQcxf4Q1m7mKEOeNTo9mcK90k/KgxdKxCu7jdVJpvVNwCZVn
J46jNvpisUQkqubQ7qFuISzN9cNHF2XFLRa5Rk5/g8M7uSvGJcZ4DhWudNgz77JmA+C7i8Ftc1Fb
zSuPL5MEkz0bCFVrU2iiPz6qRrihMhlLdUTb9Nk3uOiPvRtafTlZpXykhlB3TdDCB70+faV6bTtV
uosdkOSd45BokVlzL2DJRfbdviJeXUnyweFlOTMcG1SJo9YLUoMKkVN2BxH7yAmfTH2HCSxb+3Hf
pqZuFLHGqBkTyxU/6c9uofNgPiLwDGu4vmoWuv+E+TDGCBPtoawmdRWUz7aG72ofA61+nahlhg0B
kxOc1XbsGmCdQZt0itdXU4e2sxih7FE3UCUMVeatQe0jzRfc1fvu0MoNjvSUq+hR6R3p2knznKsB
vhBwAX/7TWe+Nr8vKd9mU/9zOiPLcW1DQ9QqiHoeSJHoIsOrzm9qfy+Cr38zJKExyNtEadumd6WV
uLxjIRIpHywOxm2URJRpTTovXDhQtlGH702cjuav+SK/ovriW4YY/NdStqe8Yr7I2vhfHV7G7O+F
qR/VHGezGNOFzAwVsNXQRnMhbOOMwjeCs3R3PTd+2n+g1uQqSAhCI11riCUeA6RpesmGJ38/3f4H
XRic3QWwhVLKcgPeghF3XFtxmDuudpv4xsnYs2haA7tEpgnot1hH55O3Vq4kWV6jW7XSHTR5CumP
DNlcubu7hk5OKd3EM7R529qGyt+6+jUWo3VWHCW/07d02WwTKqhu4pOlIdOgH8m6Vzdg1XwJx7OO
mx9jXJ/qWIdNzcjTwUfAueKAlq8bwMGw73NZLLuVTysPemF0YTClC0+dathOLwPZXGBDfg3znYE+
j51JaQi8zbfeqRq7s8mzPmWLea4ZbLvF734hyiZi3Dj6AXJVrMwvhR1aRrVaOD3bOHUa/wchr8LH
kgefIF9HmwS64Nc2V0eMho8NYYD3MZuFj0snJFuQrUZKyiEi7344xi4WvUfPZQsToKCEqGOIY2v4
TGc0BtMtoyNYKNktuYDiFk1O621vnBbJvOZ62N4aMPHZKpGgu+kXDD+B6PU0iPo5lt/Q53+juPWV
F0MrlF9zDtR3HENENt4HUsywySHo4mEjdqSsD1DeDg7Xa6ksmdY7lN539zFF6Zig1ktxNxPPo0zO
N0DrJCb2hy/yp5xyU7OzWkNx25IDBayc6y3iyb6YiWga0oKptEhQqrF5ULkvm6f1SNTSk2AhDAeO
OOA9Hd8RrONlchXFg3Baj2yOW+LAPMQBr2jAfSikeDxa0RPk5wyTlM9Enr7MO3Ry1l8Hp+On2SQV
/xE2F+iWxJk+itofobO7W42M6fHM8ENCN392Apj7eDIKRKHNP71xc1KOYKdZrIYpiH+MebUn77lk
+qYwy73gDkkT5zK6yRdXViggzGm1yY47yyqqVEGWPd/eiLHjf2IgDx3RckXLOkiU/a8hg5ZkY560
PRCcQD0pVt2PEdeW73Ow25owPhJHKM2ip8TdyOvvNPVSEAfSIAHCY6Oj8+pCr+k3aDPLtp54lqRH
Qn7MEGr6Wd8yokKzLR+PnBt0RqDqvyW/fxKxg6x1qlaI+a4H8/HHUUZjG6MSTYlUbfV0lDEDGaHe
Dm6uU0/y4aolExwA8u8tbiu6DwgtGGsw5IhMFKfNp3Kx0XPzNXoHKQOI06EJyRzuMGSnCHMSReL+
2/Ed+Ocvi/PmXgqiuvke7agI5S6/wXe9Qn5n8aQ/ihfh9r15gNeDhYCOMeN9DtJsKihgSiBh7RhF
cIrFpTeJ58vzK0gDtpaKjUHFfJo/a7kcISbFLtqAjZS6AOEHPz7HT9OkrBsHBWNJydPi0MT+0m+l
rmJUQY50pONbdMgVn3rUokCyROfJqFM5FKyN8+nfRyHN4XxUiST8fiIVCGaRNwCLGSG3T1a6tSQe
GchXbqRuXnZOaJQnlVJm30at3LdXjR7rgNh56WItqhrEYjGi6rminJqiuTpDBIWw6w/cd6CNMXFs
39T8aWW3t1Pb8+voNqRJ+kbKzxlJsabr1EBdpYIdsloRNWnE1ZLlZysGTTCAzx2WdOs/68pwTptR
39JbBC8RDKZCsBlz1xy8Er+2vW7NQBniBJrRokdpj847JO0YVjKLfs9azN3gHBdCRnZqf5AE1jie
Maw5YkM9o4TXH2RRrDjVmPPxp0zkKQm3/Hp9gFY+HMhoM9vgtvkMbwYk7UvVsR2FH/uOLnbjsEgW
jbcuFV8ieAFhwauR5Wz6LN4yFtxpmzjIwlAAbvX1vwjZxI6YH6jU61otr+jqEsYBhA4ZtSLyPUDe
ZTca34WHLAoiaa48CEUWovxpGgBo3134QQQ2CgAdB6QP/ManFW72XmQDZE+90zEpukN1E6+LmN+g
xTQqjqRPxGjZmSC1Ie0VxfwG09JSST0Y99NaqNf2R2NII0K+7fBUZcgoKauAteT/UzLMNyM77QqM
Am0PDMw+Kr1CrhIBhfyaSBfNRTZRunvpfynr263uPQ1bfr7BN3MHGYBapv4ZX00EG0cwbr38Qar0
D33ax3m79rTAYQ9s+zqqCgH7EpkMazXFjQvX0/bDND2YjEmlBljqMh91IoeXXMiOHNVyhXtjXd8+
CLt1YqUl6eV5B938tb3AhGOKNwD5O1Jqs3m1VdRRkjDW9txR8X74m2elK42Hvyn5G/oZxay5cL5q
givKf+KEKjizzQY9oyz//BwPXpSTsynreZS9ztyYC2fCTpu5w6PdfjreK+gAxna7sZcVfCl4SIkk
b6dvNAHm7znRnVJ/AeKbpNlbYFdjt1mCmsBkkLsyQPbPlCmWeuu8vEqF9vKajtXqYei4zpz9YJKA
dqHkBV/YOY8n2VrUO/8PtAo5ZCH3l5D8kEBG641onGObLC+8pa4sfMeeXyLr+Z3PlpqYw1Tv356b
VpsU1igZFleSBVftBNkNTSukLMXHKhP6ywG3zyiWYUN9/0uaFava5FNCqZsu94fNOBnEzNJ/PysE
q7Uzk5vDGEPfw+OFneSHr1aSBV3G4MrwwkPmSDTbe93Skv2mIE0Ijs2ddYQGzujzztq5kkwpJUkH
NN6u4+4ZGIFjcooICMS39Ng0bBPvFy/pqtZaKy6+4oDuy+v9ClQOo9cmAsuz+TA8PAKETDklN4GO
RnKfL1h7aSyC54WZ1DUO1M6BkOPPceSJHIbo4a7mvG1L8F2gYkfyfmYerRrMWOeSBD6SYZYE3G8S
IdapltY6hhY5bNXHCoS12wWr+K+OxdRgOzkHVCOSA6+gmZqorbRKzNbHAqafLZdRACc/ooIIeMRv
NKTsNliw9vOfkhe0xRZt1JBjtxb7HDdw94z/eGSwNe7UYY+OUEhabSAnHXVMGZstkmFM1FBvk3Vp
O8WUFngzDwmTS75mvq9sTUxOIIe3FVJPeY3P0ejYT5QHOfJhltP4SblbIikK89LKcl9xqzJbrFMC
3WHS+jxgLXZpF994oXj3EKK03819IB6t7bln1gOTPii2IuNMGHg1JcLtgYlMk1Vb+mb9jMX/F5eS
g1zYJHhreFhOcTJ8saI36VchyJ3gmU8euVDq8mUGsmOSjOagjeqUaXTbEITo8+1Nb/e9sWsntMYi
cGavPbMdAz4qNefELaLst7Y+GI6mjtD79r4LIazmCkVFDevVIRpweq78PbK7nY9F16OFrsLSqqaJ
RIfnZzIZ9VlTZCI/uYEVVYDQz5n+eqUx5Iv1KCMTM7p+SCMTnsV5IInYHAhlNJaabAncHGl6m9L1
Bxz+AKXxD4FLsbcLBFcrTcGkyFUxrU3f9K531Gmk0tu636QPRw83MF/WLpxIdi5NxxNpUrqXTb62
TurxHaX8w37ejaxGfElK6eFktySqSsFtYKJrco/FdEwI4rydaL1kU5CAvGqNlE9UJKC0i+3cJ0TB
zZV+r7gFWiNhvilwaOhEdAfqD/wctKhds/00+aqKtlnsR5IaG7ZxWqHZDF/LJiyfkkP5i+3ot6u8
4U1AB+0yKgO0r4rA7NEl28QNqRLFEUB1lBtvwlU0MeFypg8fqYHLJti0PsaFdCgRPm0Z8r6XjQ2/
DrLU90V2jR1XHB5ZhXQzPbDSUSdbVP0sVdjZSXhnIilM6UJ4JTNdPiHUIhxgV4Ck41Ixd++Ypz/8
/czFi0mg1nBg1n8zcfL7+HiNRIx/26kX1GFiyLKf2RifVjSn7VvtEFz/34W3d4Ny1GR9o/0TiST1
L0mG1wI7sIGw3rSfnVNRvad0E+i8v7JZw3uSjdtVnpXPIm7tte/aZwS3dS6byJIc/XoWOgtKWq/e
4+mILpvNauL7DHD5Fsr4vpPVsRoP21VqdPEuxsni07nqakVx6esDhD6zOH+FqfA86mtv0c3CLI5G
J13hQ7m/I97YPS3vx8W1OEUY9/5mekCALgslOyq5YPw6Gf9MCagBIP7uRzq10z9bZHPiGXao/blB
MwM5HtxrQ0gcme4CQM3Go49U9xK37ld9WsesP06JOZmgbPSiL7VLyIGpxJdj4iQG1L9geD3Gfdpa
eEmrDIylEDd+b7KlY1pTd92Zsf2FaqKz55xeS4zNMYfIDLe9T7BW7wdVf0cMeB41oJfkk75igiAM
zu1hRcdDSCmCcNkm6Q14naMQJ+F8pjTZSs2VwQzJURBKOrsXKC8nE+iaQ6xCp9SHH+0j8HESTlEw
/LSfIgvufYVeYPELtsvI7crXikHKhpU9yAxeCv4D2BqrhwtPrJ+g4hPScjLNziZzTFH64AncWMZ/
PWRPxbWFg55dGXec4fOmhUEZSvBP3SoSHISYXqLyuvqTPzx2jSaHFZeMlU7x5HIAqrVZbifZn8KI
8Yf8FzXAydBpZTVwqxb0+ytVmqL1ptyiGdvblHCL0aOOmSrHs9CpNzHQhpsPpuct6vMvJW5derLJ
ZPpKrO9wp594TqVBRSmSrP56hZFBObOrjjQJcv3LYz9nsXSXSL6SIGtW6PcdeJzlt/nCjdHFNdwS
MwiclAnt8iDNNrI/tswKXMG2xm0xLabB858wGKdDYA80olE5fmArid7UJLK+iWtj+RMA/PzNRGVz
HEjdjl4nmYfJ+oyzGYH5WaDXznNDDoY07UqDpqfdkUlL37bx3opY3ahJS8W+4lMPiXAlpiRK1lg3
wkVtl7b+5kD9syMP8eJhGGW6HMKl8IxWgw2qskSYbyhoIKpWBfGQmjxJYIlGAPuegO+5/8PHjWoO
iU/o3LHHgBtS+OC6P9I7FBeO+VqRgZqBR7U0gEELPiyUiGREzHpBBUD0ddDTIKy+OrK2S0A5gzl+
WKNDqR5o3YeBoOsZW4SiTxxjHveZ282K/Disr5cOP3rqNeFw9lHkCBsdgELMYSmVPJ/XrDj9hOYz
b6ZMpNsGslTsf4c+ZB6AOXriJG9Mni95xhMw1KZ0fXg9XQoNDs0y5CSS1iOdiSBp/Wf370Us4ZHR
bxMxZlwRYvexkMy/B+bda+/uXOOdkRLdkSNHjB6025nqW9TZy9MuWupfVVVAjzOSYRsOba+ztqjQ
SdRa9dsBwXq4hvh0dftedYu5pex2vIVWFdwcAC4BjrnEThcKwsiPFCsjkmCXzEzo+kMuVcSQvm9o
iVNihJc62VRm3mPl6ernoy9RCQAmFkb28PXXYRVDJTJ2wISQR4h3C0ENDyJaqyaG8vjrysQQ/SF7
dEvPqrr+H9rzkk5lgRX3XssFkTeIzfdGG566Cwub0K/HR7VgAa6sEecj2j1dLK1gVRfQAhPyAj+V
/mn9EHIY5wqjkrmExLu6eRBzxfu5M/F78D7FzVOSXqbJpjMvm28LeWrYXlnDD9i5rv/zlqO7HzRh
94HsyCxiLHRLs3iaWsHmJotEGV5PVFTFSncmYx3qdPZyZuoqAW/nhCLC4bQXLNSGr3Is0r5ngixb
nX+70HcfiWSgOttQ3uxrdHfqRGugjA6ef80r8bazVXsUI+A9dfgDS6XMq0qvap+v7NanD/m/6PKz
mpDM31kNxSkS3npr0VuLhWTDJoqf9C4V5TLnpWYwTKMbsXnMMOSEq5N+GfJYxv/DcaayAT9Xx2tc
PaFVEumZmB3YLNlASerks2eHdbFknjDxFSN1xFXRBR21ZBvzJ5qzIrpEummZ9Q/r4ZXdw1OozjgN
NjRgeB+bhRpCfuxq2Z51/D5r0VgG0XBoT3m9lKicnJhYJ0PdvSJxRG0Rj8Oue+U6WJTTwfxVfCfx
WxwvakSRYR0gpTfJf2tNv262BcjWU2V6wsIdfeaEc7ZK0+2aNro9Vq0JJv74sk/wJCP9qexuA9Ki
iQvKqnNpvLNHNl0uxGgZt3T28bsmVWvtal5c3cXanH9kX5ZmlsztDK6641Qz+Hw8eJiob05ydbCi
nYYFBjjm9YAyzLlePkNE6Luo9E/Ehp+IldKX1WmN+nt4oEbsToGhnfoVFdraFKfz/K/q4Caf6Kq2
gzjwfc73Xw946bgvXat2YHCKMKidXrcwnQbTBOgE3fNFiTBy2V0lyw4McOF/pOL6DYYimguv7O2u
2mQ+pUrnzElDtbMp6HgkejeOuGEHKpoH1rimvJiyPVodY35UF3CpA6rnJe6IE46xddlTXlzPJpq4
KV2Gub93YJPSeQT5a9LuiboM1bPUKiTg0f/pnXbWESAv70GKJBBmLWtyCRmsPuFGZbzckES2S3/u
1QrnxvvDHSIuCmZBjjgMrUhTQOYQ/SeTpvbLZ0JMG7ewnOx3v5T7NiAOnd3NvHa4WPQIqR/Qv4l3
h9waxBAaPqLCGfnfxhnPNHAECUetPJTn9X55FwhoMbhKBikWcFPHthp3/hJ1kx9XoZE5Q4xsqZyF
uLN8SCeC8KicDUYIgBkRD85bKjJ+M6cqCZ2wpgCZC5zb3yDpae6SWAIwtMo6wBrrSajRzn/+M2bk
7/ddhNV0fisMkijPnV22hm7sOxuxPMdhdzZAgBa+tAWDJDJqWgDUFs14m5LfLR+3ePLppjJ53HJI
+SBYulKKfsHDgPOqHnKsLy4LMBSuBMa1lBsKqQVa1CyQJ3I/ysvOdOmQwNW1al2CyQVdXzsNjYwL
5AudeqGOGuaYrThnuhWn9B56hZcsGUGO5Htw1x3Cy9uBYkmIRljWC8XyH1BYwFSCsK6IR/tMt6eL
BteeFV3tTRRDDZHbjt+idGvfSFLJyMA/KMndmrZHgCqxdCmSosgsU2C8fSQTGR+NSQfBU26l9M3V
10LMjgZyG5Kc8gV87LibnfUvfynsiwx6o1Rxn5WxRMa6ZqoCSfFwFHMNQqvDFNxQOBdLh2gdvYut
q6yuqGxG97PR4zV/KxjVs5frY6q7Leq7HfsrZZF/dfe+3WkqMlivQnhrXeQY1S59g+FssKzo7fPE
yQYayD0kqATUIjCQ6mYWwLlxco7CVVBOGU3sklR+plqxFL6Ce/Ewm+6B9QkOlG84/7ttM/ezTqMl
rtTSq8lIqM7n2zhf3zaICVzGRnZSI1Vf8bjjHF+xFWX/u529vaAz+2tWEKHqi/g55JmnoyroYP/h
tpzVMtw6I4WxgA7pKToPVM3bEOQdatyxTcUh4NADhJwHe6iW8BZpKnFwPYSEkulKxgysWyLrfygn
juL/LGGDY6DpCrVGKO3iViBryNGm7mGRTxim38ex/crqGz6EAlDmMYcebnsg9BFZVvrsGTLwVsRO
TfBGvm+ed6O+5pNqvRsY6AFURq+/GwlnTfd5+CtotWt6SBO7rNc+c46ocWrvBeEW0XMNxoIe2DBo
e2b6j4a1yxXUWV2TioEcr0xUqMjf6q9+VlYsP7tlXUeuwWz6nKO1cQAxLPiPfkiSENYvvpbXRbyd
R3sLmzYoAAmd5zh9371RoeUJDnPDpOn91qXkg8fk1TD9g4bSi6hGKnn6eaXr6fJqgu7c71O1j29a
eogZ4BfbYHH1tdFpr4K9i6pEU2FZUazEwQV+oWhs6qH/gGk2xD0y4OsvP57s2VGfKDyLtA3uYGVZ
0k0z4u7UXnZ4RBGHEcF3TGyde2n+jVqr6Pwk3gr5vgXrBSnsPSarCQl5j/dDudocT32K+q2/ZPPj
Zdx7pJD1d9ODMR61UYoPWEzoLq2YiRoMWWMEcv4p+zI7w2FKmnVXUac1LGstObjsAI0MZNCESVeC
QKHUy6i/bKe4zVLLuFatsPobPXvCzMj3kY7pa21F9115pOVe87eSrvj6qsltHYwKnKCBDVDmI3lV
soMKBa15ygMdq+ZpIJ1ApXCLVNXRlTxs42QB0dJla6tGceAJVK7t/UFH/4gi8wFqdwiGr00QCDKz
onLA7MDcf9UQktv+cT16DOQ+udKCTOLuRxfw7GJR2rfmzDhY9iFCFWaim0JELjGDCU1eNV0/7iXj
0jyIZ+tEXdDYSz4UYMaj2xwZmb/xpdx/Kt24mDdfWe+zwcUfEuwzOPZpN842t5S0YiS5WBogngEG
ETfk/0tv2P57SIp1iB8aDzyDT1ZVkXjPA4OzXH0+8Aoy1AMxiTTFAioYEJQVE1h7PBmtY5b1SLlP
DOxjXa02A0xkA+CfmW8ksVpVL6DYy12T88U4xaaqUeo+KQHldcBjBQs+l84LbmF3RvgbasQpZyQo
KiAwX2Fry93PxDPMAejnlMiid8YkPGbJeW6ZfRJC4J4/8uvFOhXwRegI4CIwmyGRmBoarpjiGuEn
loeR5lQwSurfSxyb51SW5syqVtLQbs4Y8EOt09Dv9I9lP6KluOFzzfzixtm19d2jet6mmi9UveH6
yUdT7WeQUM7wOqNCqcuj2K5UkEyX6q5mCWiNXiouY+aSvsA0gh0jGwNJgCjbdfY+11H2TC+78oI8
yFtrauoHjPCdolhBtFAUGW1RoDiXoIIUxutoJoW6t/oetJeFBpG0NVq0xCAzWNqRgUK1BOD0GIwx
arc6Du8NmQuvnBXTDDztUevK7Hb5sW/jfPq8VwQNJsexgeZRjNMBwNIm4+0dK41WTYb/0b+vG/PG
E9ZjEjIAybutmTiRBAV22sZdEUvctuoMsdZ64am1V1PeYMskiPz9+hwvJlpqAAVVy88GO7ECMsoi
aSrzWac+h3VpJ6UCTCCochYgkGdHQgR5vAJ3vXag0/a+USMvQKGaKGB6t/gWuRCwp10KHqxXRki7
qS3jj3lPVOVLRyrgtpO3WcXTm7kAo1UbAyjxFZ9bGInFEzLUBh8NpoiGOtoimx4xoFnADmQHGrVP
RjLyk2/UJIdzLSkDW1lKIfkvJwj4ZqMku3g9lbJJPLzK6MXe/0mvuT82G84PmAu6TP2z+07PShmU
t8Gfhxb3aeX7VHpLKA5X+CyPZFsketL9M/xbkx8oQnQZTGePeFeEgvl+Zhq4aQXsTUAqmZfTI6dQ
QUkYF00Fqy0HMMLBqiiPkLXW0z6hd5cmFXbFeIfbyTb0kyE35pf8cdRonYkeMVjCFtrj1C7V1bVm
mJCwSui+0gFI3Ie9Sykko0kwbknKk1F7+Z0t1cjVkWZw9zYFbvCtvusmES9xARNvDjdNCCV73/y+
TNDY31Kl0GA+ZlEG15zXgiisXyPU8RNxl+UmC52F8WhKSUGLO7B9+sV+O7MFAO2uJQbF/rZkht+H
FgyuqEdciDsi3wX5FWWKtrUNgr/0pw/HvVnf25WvRqopPq5F6es4RdjOTAXpc/xmiUKKKwAna1A+
1Cc9+bjAMTwchm2jNUrHaj8o7PXbuHOiwLixsuWJrQ3G3sEcrdYzGa8hCT/HiVlkYn3229pkq8Lx
s/QMqPSzSIwqIINP6oj9VlRvriVdm8lJGgReYnqLEZet2lgv3d5cELth9f33l4S3jU9wFXdwKSEF
42gG2UGW2rtdVpBztgvFToA87PUUe28sWnpGSxhPj2WCo3Ssh5Vh7/Ddta+RoidGmWQRXoke/fdZ
mBSlGG3EbQZqtbdv5XjYPPdUplBtU1MQ9miFvwQta5w6OlqNiK/lohdde9bdi+2YloiTLlhxJTaw
29nZUsxyVChI6aSzkbRVG7BMe29XsyBFzqjIOhkiFVkPTosAh0bT7lkiUZdav17X8cwLAhgjcgJz
B0uyFXJQ5amwAszDvfCbQhfpmCiwN2tFrV2/BPed1vh3nqr1QxRREUJDJDtBMQQc76X32GJ/ESkC
EbyHZ8cbRWcn8zhNyOJpoa+2BsZ+5AnY9kn8OKkUAOen9bnF2xlB3Kcs/HlS60dx+o6xopvnOtvu
sL8mCIyySSZdFvc73+odo1hKaD5syd/U8iLcI/Dv0pwcPVAV/cNV/jcQ8S1oBqWpGsU0B9mjy74H
dbVppq8hpZcTCMFXC9jb52kz94zihHME6xskkoH/csnFc1vyMyRWUKTqr7gHJ83/9TVWVsM2U8pa
Q8OFXRiZvvJbynFT4VCSKFkocBlV/l23IG6vw/8CRpDFhePw5HLtdgPhCm7ngQ/w25Yy/cJUVATg
21bGiAi5NtExiJdybMYLrV/8JBHMclnZM/aXNWwlv/cjaSfg1ZkD4i9xRneDVRaOWgRFnc3WYKxH
XkceXAn2gGyMc+pdXRa7ll/veksmEjf9co5IrPb3/sGmJt7a53jvOO5jg0z+glWlu+rBp6sQUF4X
MVfAKZNNHSXIa780SuxVeTKxmAKb907bvo8K1zjl0hAifuDQMECeuzEslWUGFKUXDbEMgweJIDPx
fPXwS2D3SZv7TQjzzmikX/uJ026JBrjzIoBnJrhaSyoGcfRTfAs9sH9MZKvS7Ry1FmYnvOUp/X2d
TDrYQEf8yjmCPp/6wCfTv/MrVRcVFCsRCgVVuD6xIF8Y76n6jJjQ5toYTgLL9xKUg8yalagxl/c/
/Sbu8v4LIOto+clra/8FFqSVjG/Dl4SAFlqx8A0bUcWub/Xg7ob1rOWWeGnHhBoJrKu/I1QqGvH+
j2vUhiWm1XGr0l5TuP2OfQ8lKQ5mOqmuXRbwunBsawZCtqOnNOrsNDkVmEc4lSE90RNW7u5pfMii
98/Xw297g9XVbKiQb3/9TyhqLD/fYORwMHKYf1mf6cRut6P+M8AupqHxuEC+zDyKUQi6/W/AcyvD
wVFZ/+pIV8q8mHtPmgytvVZNMPSEI6V2LoZrCLipDwZWVzomgCN72crH5CUf4+DAITqSPICTLxA6
tlpSa601pxwquOH+l2lEtaVMnnEpIjXVOkFtrchP+3qbLvOg6tNx7OLiHYjHTS8/fzc8KvfHCvSN
7W4RMaxRybziVf5KRlpyPsVUJYc/h2b2mpfU9cmb8vGQG8zpSkbHa0Kvk9oDBr9SIaTpJBrogY6x
hsk94MFCP0SytvrBZaEfuXguL9NVEDEMWIqMOfIiXvuA9zw3J/rCTnJavdL+Z5ElcUViOr2XZ2Cw
4BQD+nayHg3sEEEc5cWSvIKgdiqqLerHqP1iRbpK1OxoIVAqaFRZTol4EEEe9Yurphu2DyAUYS1K
9yNglM0FGrupPgTSimX4tBcp1QVFWAcix0AFtygej/KBZYIXg2NkoCWoXHRncjVGRqmtmonizvbZ
QUjcjCbnWxh+bbp9OAekatEssztFePjzyCP0NocSoEnYyE4fvLtvvRL+WiHO7Rt98XwiiGQtF82k
qyWfYB5Gi52ObCG+sywtKidGXfJm8s95SZKk40asgUXaLvEndC+e+mtF0/eMSKzeKqipujxLboNq
aQkClz8wtRqzk1ZeVwbZ0vmDXq77CCGQs+JkEFTPuuNIbZQFF8JNBeoeXgXY27OEnEx3miDRIS96
wroKZlV2v3z51HopVEY2sow357wvDirrLE3Mv5Cb71RfM8auCTujKj/kmusTwzFrjaMwzLWvLrqh
vcahTpGR3J7cL2YyDSAUkNW5juNBWSYV33wtZejqFywp6szgC3kUDSrUlV0u0L6afbvoA7WuFShD
3V/2vkz/0aUEuywbA4vJiLewxl0/9hLQJu9E2VxM5etweg28PBpo9NRMXA1lXhXayK3hhZP2Zu7g
IRVTTN2vMw03gQ2oa//b3oJocXQHZ+eiMni/8esKVAJi148YOyZFVKUgqBqdssehBpleJ5JLy6cZ
kHme3ZHTP3BaHWv9o+rZpofppUQQ7a9bH8DHajkBMjIBLJ51zhybIRGIldzxAWqQ0TeQyAeBCrNO
XLQ2vDGhu9IWwTO+GLXisK/EWgw/UTG9AKpaIhkaX+rsh/42m4DAUeDY1G6Zq4xuGVgZMjqwEF1m
weBmlkiwLIeWtYWOXqpd5CIBRUQo+EjAsVdm1IdokUHL3Hm+QPTYdw2ursxOFW3CZ7Di+mV7zOqd
QXUxSD2goRL7YAiStX6wCycBKd/4fa0ExM1Xf1M4HF+nKEFvBiyYJrVnKoXgLnABUmpK5qwlo8yt
NwQUlkeIluTXjnA+ck1E7scARXDgOQ+9vZKxhEuuEoqG1DXLNufDfZrunj/5FZXp9x7kXK+0JJdx
bUF776eCYZQTuJOnJk3mDUNNEUAe2vsEnboxlkOQ0gkwLhdEPe2XUNYf5GPbr3rirH531ZpMa1mo
MQCU+NRXHFBuzqTGNNWji5jzNx/XDQpK7Y+zNH7R0m27AX4o1bcTOq4rBn1mOWPaKbckiJ0xalNw
iLd68udtfURciXgoiBZ4vHEk/OJEggZ4S/4JY0owFTfzMsCagnRQRQvml3LpFWkagX9x10FyuLSY
Qret7u68t5PbYyHp4tL5iQlZXQbIu0YHTTEC0803V7E+j9LrUdXl046MCcNXWRM1JHSLliToniKH
Exh0Rwiuq5D7pQ6YBka/sUrxk4PxXGhWdEyG81XCKg0dITQN8q0wB2/8XVCL5QYjcLi1OUBkm55H
ndGCK/bEv9TO+ztKbB6xAJNQ2B+icQ3bpHQf5UjH92frNJIVENbz6I1Q97J2TV3gCdgm3NyULJ4X
zdmUlAe9qS4DM1PmK5eH+kuKwwrM2mdemyXT7Ac9o2YlfbjET5BLdSdv/M4p7jAvSdnWwQ9BYPa1
e0Zi7OU35gkQeDuabO8XEooDHw61maO6OyM97PupdrxoI5H+Vo661oB15f1RQUXNm7GjDmvhxpoU
dyEnMe7ZVZnJmRD1KPWi1YzsuzXLVEOxKc0WpOulO/Pk13PT1cRfQYTKWiQkQ0W2RicLL+9vpMxw
UQtP/FQt08tdwJlqw60tjJ5FXlUjI5D3aVES496zaolNssJ4l19CK5UvY6m8cqeLXjb5y/06BMQD
w6ajMiqx2+obFyJR8v7EwkZNyXNxr7XrVwzyHBnL/+nQnTDDHtlvggXBRe5UKq0xuKEQfN4X9qxz
0RqF1DwFqqb+FruL9yHXOWv3n8sdg2SohS40wSzHHElZfmI4TJZGrUXkDSBIFZjuwkEwvmAr66gK
symTVOzrIS8qneN0M8ojd5zwPNFwDPVwWd//24q+hDi7EPjt09lm5IqcmRkYtIGhC3JTn6Yla4Ty
03B5lx7vLf2GLU3zG0kOMCpgZKMElYtntFlSIWIK67EdmFUFH7ym1HxGeLuYjbCWcmCsSnC65+zn
I5eq9eAAAs/YlC4l1+r91KKh2mSDDuVdDUqg21WsD6vSMoeMXMxT8+mhYdu9AQrNpvfG3u0bZ9jw
kph1phlykLHruZtp2i0E6jTi3rLWSb8aC7ennOiPo6w0llDmEooJiX71fqvNh4FxOw7gQEwHTskR
AIvg2KO3uscTHFqN3YKWvc8HdRn7UQyIZWo6y39Y416bAoEu+HS5Zm4hhjpVe6xO8gkzp213O9Dk
4wyB1rhv9+Ht2NUMkZzSgMsKRYuhCXOod0mym7ahowgCKDqrzOu4xiPx+bFo4sfDIf8WuqGOlZBO
rJ/mBgL1r6rMlSfMBEwMVxJw2hrFmw43w9F+8Q8VSfifJkbwMFcqMx7VLKcEGCrdl8pnG+oKujoU
PbD5C1tMY3TUgA/KcoABXOjCTxn/2W3X9aa7p4SWMw5GfYeRlLjqm2ZwCpGJ4cagFN+V57M5XIXK
jp4Lk47sfrioJjyNtTHxEh0hNVYdt+ECotKSZqTDypHol/BsdtJ/JB4/ary7Al8JKYQrs47Kqnpk
cO5EpS1zSSPNF39V9L2PU7KOe/ios58JJZcRViN1EcsBDeY4fY7o9xGMs66TtDJHlpIYjqSG1MHC
18eCOlNCAIk8zElw9jPfWVskqbkUixDj/qtaSFmAmhXDGOrx9asd21+OIV1kyZhg3Xy5E5r9uc4M
yWPqVTlJbXCsJ/f6c1GRAEeGkfoWWPKzHvYLYcGFh66OPbVA62c2UmMjROZi2gQkJ+FOhD3yVmCi
uxdTyJuOQ9Kii4hrmZZ5JQEeAL6KybWqseKfpFd7uXmR7s+5WoDrbVdJFAcqYz6qy0PGL70FfbJA
z3IXT9sbJswQOw+z45VB/Q/T0QVgwWkGyrHoqM3MjlGdodekhuOXO0fc7f8fcFUHOM+jMi1TyWqv
ghiX0x6Z8e84VP5IMTV0e0N4rfJ/l1uGuiU35cuV3vk58p8DPKCApSJiFgKS1CWGE5h7+EbQdje3
/17NgZYndEU3NfuJk38XrI2w130Z3XgCM+uDZqWSLszHfFqF776EUNKa5LhuHx9NBaEtrxFc9lA0
tbCN8omCNHW+FbgSteh6n+KNn/9AVR1qWS7EcjKNdWP59q4OfG81iP+kCZIyvjNDudBEGuq7zCtz
BTZCVm/ftYhM4VX4UvcIa8ch5yrg3C5alkA25bzHSRzGGdVoo8QPK+wPRlZTX4GpaFFjfoN/YDSl
cBd70l6H1eIVT5o9FmSCPqZx95J49/EOOfH2nXWcRK3NTFnJAk5TX1Ks+kuiGi/Fh7S0nOxqBsmI
8Xzez7Q670HWtdRQ7xAChA+eevJCC/ATEnbQpqJt6DRmCEK1R8G2LmO6uPatWbIP6d2iA/3/NqtC
N/QxkoFjWHWLmgVOmej7w+sxkCU5Yq+92HrY7LY4hMBAzYPU3FnayFJLawItScsvaazhUR2ruYPg
R+SjQP6xS14aqKTxTZFbQuC0zkeTJX0ytSszNPCT3d2oWgwXNtkeSz0nEO4Ppc/aF4VCUt1yqCst
PWo8GNjp3gMbRwFpMqTi8/sb+Ba9ZwDO4jRXpNG1wEGkeGj4JZ6JSrHT3XsUXARYSlFw7Ym528rA
MOI4aqBFJd5pL685DOvU7A7GeNlC72G6c+zLKSFK6N7n+xVbB8kdJVLGzHguoZh27aBa9XoHD8MP
WSvJ+LpE9UcnjrmZ/AfJky85MP4wy0sYFLeduvco72WUuij2B967t8nKXpJ7RhyN3HB4wiu52b/Y
/mc4Pqj8PTPB6oF7zqQtXUrZh3TMlkKN1Sggh99kKaFXc2d8I3VuyTZ6PCS3dVEr2xVnDmf8B3et
X2XDuYPPrc34VMIZUdBf0cKrQrvKidvLEX4d45BiWXDcgqOAdhyOq6+3i4s7/bu/4C/yEVvJIC6l
wQV9EAZihkmrSe6xP4sbiFBls7qFFBR0T1rDCQcK9A+sxyYxWHC45ZnJmnaj7MfMa5/Eq/4JoSQ2
nP/X/lY1sDbioGj/n3UINZ79qmhDwgdd1NmrI1legq8CaEcMK9gmdr1+m4ZfvQqU5T06O8tSTnvL
n110OxjblUXQwIGOqtgxR6HFJ5FFew+v52X+8mK/8LyRJAjQfioEj7M1wFBfQpWhzVR83t04t1m9
0uhqe9/tc4ws18Qhvi+WwOHbwtNxSiQSvEtyPOOvMuqYTn6jV72fa+MfJeX0IcfytjEwyjrQB+Az
UbgktjwuQvWPjRjF8Py9XIQTzPAXaDN+DWUTU+we3l/eju2f9l/phnUbNTql6Oj87osmdF1g/pb7
S5oWLBmI/uyYSn2ZV83hh20vJOo0KGVHNcIjAKBfYmRdPTdoHW7vu+/mHtRIKdROiOAQCNmFdN/i
WIxULZ1BX9VG7/iDwrEjVR/VJqQzbjXlJ+X+EAfNpsUv3wnixhqVRYIw+gewhv6irZalUusSPDfQ
QwUlQ9AD38VsptaFWxZid4I+seuTCC42pHHYVNdxuvJWGDKrsRnIELK4XwnIq+ufe38kxiXnlqIY
6R4mkewkAUnkTNzbOsJXYjkPJDNnIa82Eo1BoPctUrhlmr2qHTFLwRN078uw5dJ+XprH2Su5IYih
yCLLEBjmrk0Uyuw8QNHp9ScYwPukWnmpfPFspJNgIGQCpsdmHsI+R5OC8+w6qSoflFkIrU7vtQJ9
kRrGZS5PVbpdh5McT3Tq+Ex2iMWlsNvalBkSpSbHmgT9M4BhK6vBQyZL0nSlEIQm3Bnw3UieevoY
QDSdIgU0qvwNMvZ9Tm5sA4JcRPn7queEqLNWaph5vwZ6TmT+v/f7Qz5ajI5lyvyK8E9fHAa4iEVu
IOijg4jMpV8GUlQOvIypKGkxXRW8nf0MZPiyBqBNjMIYalOp5yhgAQSfPJ2bX7XgXZLtoNnUBrcT
A5iGJR5BXS0cMi6Nh0ymo+JtYt5+tgM2dkQZ4Sqfw0Nfh+y+iY+fuU6q2HQeq1PHoM2xg7x0Em+G
+/SBDjca9uUsBUShaeG7mp2RzBBpzO5pgEhXQoujs7V7SFvJb/FbNtlT3+BBy4PGzu1N0bdiD0Bk
51Ca7JK3UVbJIPsrcGmWP+QyQeG5bTMOY7gan3NycK2QSF2NZkwvvOMCZvpCSHGWYCXr+3DR6qEI
hQ2uQDKHOztYr8SP0na02C1/JNKCcJOSlgRsUAtu+qG0qNK90+6oNLNe7cfG7ESJfQ9eyr+VW1Q+
MuZ++xN2zVXnS+LAVsiwXtEsqnCsYIYHCV4G7lRzOuaz+YEUL5vgrXpyXJVEfliGtq0mod57VwhZ
mXqBc7dlJQ7qkQ1ITiFhZy/fTdPC3QoFoKfgUvDfuNCo7zcV5jmcukmkMROdnOwViisg/0u00Lnl
zJqbeUBC9SW8OlviCMWeLhLGasO5AxTXnjhbtn+EXE61iMF67JOCoEeYO2M/9m/VF9Ttihd7smD+
aaxe7m+zsp1kRt41UFsQ/LZPCZK5jYdyQEILtc17x6pa56ROjm+G6lyjGq7GMr5dgBL4f9XcTx6p
DngtvaklMphUhRT25WGMj26Us4BUGVVZbj1zIG38WbZA4w7bd0JNYAGCkKDMOBFoUcJJqHJA/bUU
nytMMPYoudTGXxFgo4+I3DNXUk8OPFYpYFgsiVNv8KYup+vx2E5Ix1LS1fhajI6laFCy0fIoIANv
UeoL47hYsJ1poRRxND2r90UKK4Bxs6+hZXlMb2avn1j9ciHvGpJu8orXWPGzhdhcSBJCxsnBoo20
6mikuggAO1ODebeowcfAjDGRyhr1uL5Jt+0HUiVPtWmFtxsmcLxc0rjV+lzay0aLamp6t9yGrJ/a
gqMYVKCM11r1zBX4fOrTWYsotpP+lHM4bAeLpelMj4MMtM+XQI9ztF5Rp0ndTyg8YSaGfuTNAqRj
r+ZvPIdCNmqSCWzC8p3p1QkW6vDWMMskeLkZ3bsxJcVm7P8N8jSIiNSJk4aRyxEszhL3b92N0Gv/
RPZEdL7Bi9MKQO9WSpEi2zWtVN+L1WERQs1Dn6g3v1AmYgjx5DwIsAX41iqRpwSY1fEfaB5N/SnK
42GbdNCH9x6BcWVBfwM/pFJJYHs/3CSU5rCgxgEK7kd8RdV1Au2Li09mGQoLhGHKB8ZgAGw9IEjp
uoibZ5JU06R6hhqgqGiEW/GJefIG5AEsZarg9HorF+RM5x3tnnHWCkcQLIkgcFfaczsQ44T81yCZ
Nlp85jEcuLODBkOzZoxWhMwDUfDz7I8D47EmdkzBol5/KbbBAGAopfE7/DNEfZhy//buCfPEtmAK
1X0pJ4Vmmh3e1CuLIK9kcCLMPy7QbXDbY1UX9cNovwslMHD6EjP/s5iqq5BTGxc+7pv9L0XBRNx5
tCKS8HxEdJWcRI5MK6YFGXZ9eJZ1mMLIC2J3QEAyDMkXAAGhI3Me0wlO41JAr5HD12CUfZl601Kf
QrRHaAA2GeZ6LgsCalmp/67PRFfRBhnvFa0RWkLytYDEMXWtTl9McWafUbMDdk/bt6sYgTHAh9d1
YD2UqAVlDwL9uZ4iwU+y8D4m3w3qJFqumhB/mT71qT3WQ/WUiDPOX6116w+WYKeTYr5q8iCHOAaS
7dvRnhLOvfj7J3G4ng1GLSLzoTQGnmJATXVfgEoAE+3fGMIMBpUTgMMuYqMGYiJ1BbYz0rhdHv3l
qVm72q4UVFYQ1V5gJae1mz1hwxXhFvXJMd6zzAT3cFIMO4PlW/s6cHvXudBEs/QdUefsY2m69KSV
5nYIuRZBergsM6YJH+vkM//OgwRAKfFwmFxN4jElxuc3K8CSsKOPqeIyCRSB+CKk4ACnoKAhpa/B
UPi0c1mHNb4v3mjnaB3NTC2rnu8bt1/grbPskZKDVruMI7OwP1iQ5adwIoAKQ3DhSyqmJsdHkq29
KHLu1tYNiQM1Ftoiur9YgCeJX7qI/Tmxczt8WQ3cBsyE/13nwp5rBCiwgUABqJsD991Dx2R2fRqW
6wlUbxhw3OaaYi/C/rBTNR+Gb4nV9L6b+fW71JvsI9JJltemnUupsQOq77F3pUTFLBJY8e+8Z6Tk
oqONreKM2Y3eJEGTeibhQgSqNMO0DZYDyg7kCI2E4q8FLftFSI5elfj/zMuG/61WLqIuKr98cL/l
/PFA+tOqZbyVjkN94MnHWs1da1xNxyjmUgfcSamgm5ouT0s42zeTMKUyzxzaZeix69kYWTebTsM5
gQjgsG9a2NmaPsmBsnrgWiVFZkf4cUohvXrBVuiQTTr/Ro5GTLgOA1zS43yjYsfD5K0xt1NGNn21
6308KfpCRNhjSkieUHhllMwp8E5L5gPWGD2rN9IiZ36YPpj2BFaBc30wQ5eHX7cUttt+mkuFzevm
fZG5Nl5pD2ZvIaC0m6rWi8pH4zkAq53IcSbATsVOf0AlfxwzFzEhoAw0005Ph+8fczVN0hz2LMaP
RoDPHZx4erLTaoj0qhmnMHXfmpqBG/pDDI7TGOFZAmx6VrX76H249JfdMU5dVjg2VCN1eeik2CKO
WiEE63HhkS3/I1QrbcbDEluz7YESP5QNu4fpsKVt14Tm8cRUHMCnkdjZKodmMBQhCWNleMiwB5k5
8G+ZDJIUDiY01hbMLeBNEFBa3LLUS983Tm2/P7menkkbDAaOJG8qQdTr6mtqzNFngZXuZOIBdNxY
5nXouBO8YESDHA183WuN9XPDO0GQFuaaCAehrrgOrhIWo2MU7xpFlxzm0wThQzX2cSZyWiKQ2gug
/Jw90wnt9b1zn4g72qRLRVbFjAAG9yfyn84aqHpbMGvPSQGnizc3MJopJ7bMv8pc3zBzQ53dj5FO
4aA6YDlPRpdgGXhECF7zpY1a9kbl8ARirjU0Vg386YPTRL9AHJcXvFIWsgn8UqsiAogmazIwzECb
RhNqwDlwztNUGnaLFd7FbwWEAiUf4kZlRBVSM1cl/cjg0PsIHFb/a87NG2tq017h04dxuS1mIq0L
c2FRM2KKr4YE15bGP55qSsuhqqX3Wdj3VH0lo71NeJFDzUqrBYdorEodwaBv/wSawpN7rDFaVrH1
TTeK9bCBSwAvHjJke9zcL3kcCII/FfEQIpTZCc5KAKamsa34TGdBTrXAwPNJMhxEDPI2oCK5Z5Pa
LrCgKMGpmHa02Q8NcKaEW8KZ1bsr8cCKRZnF5OB/lrgJdt8mgaatdCfLBksxBeLM3R4gSf4j0OVe
XpseNsKT7XypG9l91qqMvhrL4/0twBiSPs4DkyRxTbvJPR6AW/alzqXOO1AE4ckbJg05L7SkTw5c
at6BJ/5cx0sBbTlc8AJ5aJM3RfW+beA/Iu0wOQLnRLAXfbYtf+rifgoEO2f7yJCUOmOVECq3G0kW
4dIoKN9mRbWj/aRGn3bEaynDunALY3dJjOdkKYaroZ/sCHAMeIFhylOk0mB4pRitz6zG+wSuV/RJ
WikGLYva/DVGOm3sWAN+x/JYRHF0bEIUXefqFccjQuEktJ2TIfoR3Z5IaWieLe9SECAvLIb2+ilU
FlXuluUtTIqIrfZhxyzcOEWGYJCG1olhvfF+k9esSbH74wAYAsJO8udRf2x56kFXdbI9HUzMdaj+
hHsmG3Ui4P++wuwLYBad0SbTI/L/u8aETAk1qWev6yjcPE4deZc52odXVIDX1b3TMYDGQjLArwRt
Op52Um5a/pBwuImRsg8RTwALis7JLwawvgdKTbMSzhzAX/WHKmS5OueNQ2a3pFOnW93SNV43Yd2n
utDOPqJKQUSxz9VrN+fqOla8A9sRl48KacVTqkK3m91tmZDu27vMAPflGcAUuNgKc9A1eJd+t8bh
gwxZKNOaTbJm+ho4ikfM9qyHvQKdxH38kiJrg6Ipui+ScPIUdwhgnDdNdvVPuHmNbNxE0vzlTKIU
XEUkQwYNiKc6KBPRE8s49O2SXhcYgXy022cA/cKrUKxK3XIA1+J44a1KCTta42e5jTXTW1dVfToA
Wt6jtSQe66Bzrl9JTbuXzgfb4PZ5puZwJpi12GK13MZeqvRK1Vm5Fm5qqEyTqTaQrQGyz0Nvfcbe
PS5KLHPgqqTIK9W9ZHjsD4OWFfYU/VkHPZrENdlTZRYRWVeTtlXUuvZypjNypNAOCh7CFAxttSEq
e9bTMFNGYJFHktuW0DG2XMy6FjLE7WzYxzgoranHOMl0EdoOtJLJIkWkA7f0NBaZBNWMsu60XoyB
n5xyV0rbbBksC7fJtKF5U/kvQrzCgnL12Fi2mzS/66OTGtyupi61jEcXLp9Sj+7Fr2Yfl+yiLpbC
LHcQfodYOFKsUeYDwp3InuA39ySPdtJxbDTE1o5X5Df/A5A+fH7ohHhxEOAC7xeMRBZ0HlDWoQp6
UpEzcFx7ddOBrfo2V+YZWnBDwDrP7YTYGNpUkoua/XvcpmtPJfgTMMb7giNr7oZoHo/yQEFl/Isv
HbqUAMg8+IV0z+j0UzrOGHinASuuusqKW7lfLHSBIkS4SEiv0KLFpgRBIFw1AIKtRmiS9ccQWPWj
09IqIwpG9CB+szIAz1ouvQ2L1lRTLu1QCaH6wqAD2VScaEAIlLmnwh4VX4gVC8VXR4ai4SFKMmAI
jzEo8MOtyejW3aiSqYU84xByWesmafnSDBCtvRq/YsxvuX1bMgdL+KzATg+kH8mQgibnLhIRz9vY
aZQugmD/zjos7PLJ6vLXAWfph7zxxYoqZpBsD5zRF9xbd9o5n99hjnzDTr4RzbUbqszjr7P7px3Y
inFo0R582TlW7UzVGpqqdopIkiVLdnNDCbA57WO9yrc2cV/lW5VO9zwij/nI9+uAPdKqf+W7EJS2
M6djWT4xxNo2qgk79s2mzaJf5nCWSXKcHXtV8wI1c2sbmtUt329IfIKrnRRzWRjbwqNsp4zjPRzG
5w5JQheEIebgzAGASQ/yLCpqSKC2BVkiik1h/cGoMf71yDGm3apRU2iDrQZB+MdSxWUxlzgF/jEi
pdSqqzMUg01PrFVfRFO3T7Uz7TKSNDtM1d5FdY0Q/S/JRI+MntT0VbH0afw1JnNr+nWFT8hbyJN1
CaZz5iF9LETm8cqkJ5DEz5/1t3f2GBYvvKxL5JvdpnI3ad5+WEGFmxT6ZeVjUapMFwDOnpmEsxU+
r557KNCtv9MRGAnPCHS4w2k4dJSe2qxmcqDTADkKOmbwXnLRqeZtJwAFOS/fXVR9lHZt7NRTftei
I78PabAtc7ITbGoXN94VNAN8PWa+YTqHoXqenUJrTkCrH/y94HcLhZO90zuThGe7sEphOazq/G08
SRAL9YCkIKbaEEZDMSXqj5mhEdZzCOR/R+0aRXAYnK4YfrYgHuiXM1znRI3YcPx9jaaQzWuhkTKE
JMDJiPaa79qakQAFHILR2TQgxKpDN5OPvUNpSBuFQImBkFmUg6z4YHHpkL/E8Le9qyb5sToYXcN7
e9whJqLZbWTeA+R9LW6yw2CvYNNFE4Vf6sWwbpX+RDRpG8bKJO5fyVVbB0UtXDWZDxJoQUcH8Cw+
Vq7JsU3VJtLMGD6ehDYgqCsg3qwU3V/B4gTBWwlLdhXsIg4nXlgzJj/Rs0l2sVwVtRwO5WZ92FWT
yB+eViIHy8lq2OJH/+So3O/zDcz8hwRb+uhmK+jcbNsR73DYmFwGs9yKdd/7HfzCnt6wZ+2RmwYA
WFrK0wYnEoJjfE0/3+kEfLvOtqAX1CpGir8Px1n6xSbGzYT2YP8Z1fwEXpDQpt9eFnTiIGV4spcn
U+aXvh9iXQOu1XIV6Nw48YtM5cNcpxnsTxe3c+TkdvBa/zZiCzLW5h5ARn2U8puz/A8PcQVu1fMu
WVsJEMbBnoM6zuiuzSOgbU0Qs8s4c3G+73K/merNxtNP384dwyHuGpdSqhjuleZGB/nQI3OQM+Hp
L33nqWr2Lcm+GA1oIE94Ai3GDVue1bQxOJk6MJ9o7/ndQz6ea/AuqgEBDyEAodXg0XfILZwUhlTv
9evkN+MPfjCa1I/wl1g05haaAF0jDk15TjyUWpyrKJ57+dIBkvVSfwgkE8rA+/cmU6vYCcA4CeCi
IA8gWGBCRWjzloP5H2e/xe9Q/oPzpzvT6QSi6XK/4AeZrwEw07MnsHQjt1azQKLaTzQeonL94+4c
xVBtxkeEF63sbh+PH91tvhs1ZRAN5BUrJYVdv+PUXT36FUQSgoBoVnNSrFnxwQ4LcyLMjap/LPeO
82WJ3lNKl4lF7Wm/snb95vwczROPNLuCMy6TQX1dRHcZTrd5v6Z9fKm+2rclPPQMe2AaFRNH+gZY
Zk2+Enos7akRuz5hWL7cnMG/ged4q5bJqp5MiCx0XC6N8Ue9yv6FeWw/QQ/p9neT2iQbV8uNmHlK
0B4REge9hbHi1re2kNmIpEHQu2nWTijaJv0MTQeR94N5c49KjJl/6KZUZFNilS+5+L0eRWcgnZpX
IyUPB91vCN9ayy6a6QT8Kq0yMvFa7JiOk8b8HEl5PzgLUONdy3DN+KdqJyQYJpQL28uGWlVUNkOj
LnuCqQODyRCOIlavp9zBayGFrZZm06G5/N/e+gC2LCS4M5uKCkd8D3H+JtahnDXh5CVJNs3l9L0q
xvet5K9RR7d1xx0F62CI2w1yql1NgiCfZUxt4D7ZdwUdp8B4s4V6yldQhglicALztuTxw/BxD2iS
+6pueiBSnNE2BN1Iy2+KOlVBcOb9RncqtjoP4H/yXCSP7qyJIwSgIJQ3rQgzfgLnh7N88XO+5th0
+xP4pkwRxBuCCbfOq9hKdmT/aCbAalM3nWKQ1TzpA9NRE4R9vqfhg+fvZWvmJXNO4K/ICs/aCEjV
2z629ohArJEagB2xtDG09A6lzD2y/umZiy0sQdpCAyYj5Km29k2Ren19g2WMty0qh9jUSwdMJEiP
a1p3HgRyrAoHe4KfuBC6Fiue1+3EKnmpB5lT5WWJ8f17FK5nixEao+LvEiOajDL3CMkIQM26oJY7
zx8zLVpljWmIOdYPJ/kSzDQC96uArsjbFOpIIWnAdK9hO51SMbhEg9hJeiPBgsRx8YOxRMhZdY8l
GEKQBYud19nonef5Asc2ZhD3njFyezivG7033pdHG6g7mnK6joKtZy9LQf/ByX398FE1quwQR310
KJ+5r8owh6IQo2lSmijoQqLXntEPst1Goox31vSW0QKMh2B75bozYekdOav3LP7NfyWJ+JDB7iFD
UCyIsvtlV2pd/41+jWxC40fvs2vxr2vNjpGisu7E9MkS3VOQ+ctugRqRY7t1Aoeck623OEzBB6np
/Ebf2pqY93tVqYs3BIuNzRlQkw+naId51vMLCsmKyVq9jp9INRpIJugMKaxYz5TqxcR+f2ktNSy3
ceEZoPeXcQrBlju6IhKwWwqsG1QT7B9P0p2fjZQx4wBixXVeCISgIWrxeVytIZnpmcP0j4IQKYBW
uWvFJpKyrcQ2c91jUlAREBgmW74i/H6jTEItFGU1LgqC1MqWyg9h0oWfzJbRniXPLqk5RMXbD4+j
fcHlGx2thp/9zhJectaK8ojAyWnfG2HKXFl5jsp29VxGCo8eGVV4VGLWsqFYfzEbaqmrBGSz4Aey
0YN8eh94kie4GvIxIT3IqeWaEIXdAhvj8Zj2BTccMSRFrEnWoac90g3B3ZnV3crHvD22XJPjOuUo
SeaBAIoTubCauhhhzyHR+6C9tAn37z35pCDTU6AXK6OTrXLLjxybRFGjU/p8uDNT3zj+L3YoVOue
j04OoUKEHHo9fGEQrtxiJ8AItJIuxONy9SfaaxUmZniU+XF6tZsh8qTBgVbXkLnhxaUflpcIqSrM
OFB+vEOrmB32xROoKiZVUOASai3bIxo9zmO59M3FthCk0M46/nONw84+aeWE8fxBhmBaaW9KPr6a
16cQRFENEDRQG//YgNvLdg5dPu6nwvhgjYBteYZPGAQ+3AwxyNv7UDPqCoVXYJ7Rzw5tEwBHAlqm
6zynAVshE/wZUCdqC2qmIn24f3rT3DmBPcNvY8x+6Ht4qm6xEge4d7T7HV5j+0MDbRUFoIB4AydU
+5G0hFpPBydnbLRQ+1VpZ4EpdUdP0YKAkDTGrU1f1HSyVxuDEk0LbDF5xvlmUpbXLfUSChc7QaJv
oleyR8V73G+sXqqwuJYQ98w9gS+OPnm+Hl2NG1lHPq9EtN3Rud43E/2OXQVdYT5rA3L7B3QjM554
8luPJqiezFpYprzGOAmyKTHq4ps1bvwcwyhIvrSSxFpy0epiVEWDP/W1uTl4zUPly0kMTNgQjk1p
ieIBUZ+cSC/wPiSooJ3n1nWTuG78IDiFHT22RnmQqJ6c4bb6q1sDxBXT9kAreLM3kw4Lqvtj9tD4
skp7ASk1Tdv1aNlDVLLNJ5JGCw4twcjtHV581GSGicjnzYlEqmoFHP6azrRKZs/+1MIBLWJ2xeYs
hg6VBiyENBWdGf/hX/POdLozmzfInlw141/B0Yt64grphlvp0HInlwke03Ox5f+UsPadg9ekULzh
5qOcYt6i/A/iqS1tcUuamaAeYjT0gG1Sn1YI+pnQPtYKfceUrGr5td8cWtrP0Ur8oMe9t+vn+5T2
pAx1fD9xFs+SV4RePk7FrrHOt3Gv6tw3+JKI4mt8sg2b+w8U5u5EL58Ap2Sx4m9cbgGDe4Kmxw16
kzmpfAO9DvQMc+QZfwK8L917xLmO4kjkv/pBRfsxhekQwGVGNx4gTDRb/xXaIMvwcm7IPV1ztHkz
mT2ofs2kGAmACXyLrr37fMvVXm/IsmHpPWc4nzOebwQL+hNGC8fgeUmachfKEdsQ8b4N9uy6bdDF
mhelrz8cecD+NzbBcAwSjrp9cOKh/kqEoHRl/LFOtcCsIgBBwZ3VNFMffrYxhxXv/MEIYf97T1AH
gZF0GLmLERdWcjTgzcQGrq4GKA6j2FA6f330r32tjDmKL69p6xDE6YMu3Ksaq32s2AQuRDpk6Qqy
qLE9edH+kxEeRkocv0DfCht21SMSnuM3NgroZ0pqxXE3mP0E2GQQcKXJXQtPjKp3UVPNfLMu3m4x
5iwKL6qKpY6QK4zwZYKbcBNVTLBElldCYruUEFe0W0+5JtGBNq9BAddz+7YWcz/aAOoKmy/cBxk0
iW4tVLO3txFJUGSoVdym5EALfnHA2UuX7UddhV5WelT8hNwKdy7mG2RPVbw9bWfZvFh44N9Oof0s
m4PdNCOnTgwH2H34uK8jrk3YMwzrYRQcIp8/3ADFhXG3gFpepFmmYKyp+Aar/snukXIFNUp9fOjQ
EpydIfQhg1U3lD4IYwHCXXHhhFXFyGuj2WR6jCssPttT1zx9tGzHEVO9IT0uMHgZT+WyjKodzQW6
Nbwk/gWZUC6v6En5DU1bOulT6E2VZaJSpeVgDDurhayABeVXO1wYvoOis/3Pp2AN94wixhbJDjpV
GXFMisP5VzBqHGnmqKCwKMBMwtCx5/6ItK87vIIuw0sCgee6zs4wZgZt0n+16Z1wwUM+ufxupzw/
VOutD/AfKz9pQtY9PD9m1kqINw7IYUJKxNp/MdL+faNeM36+uimQRF2O5Llgr6dPujK50b3Pp46U
Oe86MJozswLVgxOlk1SE8ep/5xeyhPjTZcBRPKVmoxCbQ0Qqcy6p8PNAY8+MvG5YsOEgS916L0By
fwVmf1Sw59q8DjDYvpr5XqMY9815I3D9gxzZUq2YPCT75pdA36hrfLa0XQ5TAVcvHvgvK+KkAsqs
iHBYZELnsR4z7z6kaJcE5U75vg9M0IYnR2mdpyrje6zMoG4Kt3CwCwyrno10fSEz/lrhxeeIXKqC
9kTXrjZ0Bhhyf61X3bR9Pxw8sr4uWjIrzMqchIqqUSQEJKH8lUqRRw4sQYZpaSoRGHEcSNKDAxfh
6X1ihg7ucL8G90y7lQzQWCTIDzpMbwQ95Kz7j3DWgxJUpiWKmaltrdvdwukAj2+4XcSGmZNz1/D5
6tfc28Nm1HgRLvcVwYJB7+o5tcwG7o1QGSKf9qZoo722R5dmXwgYnLLbxwyZI9cr3AA8BorMExFt
vHxVBCcHR2nzbT3LlN5pBWW2x8nImYxaXwXfhdTM81ntEWCOZVGcyqmLqXZeapCN9nPDekVxWDSe
WFtbuH9coZyL5JZDhQLhaItC4c4mAr5PwGo7V5kw/tvjRube6QyQa7AyS082GqLm4inu+MXGvJF3
FTGGIWSGms8rfTVPNBU/qLuspMhT2awhU4TMji4oaqb3db6iqf9ZbpPEp9QpnNC5NT4GcvOAh9Q8
dSFw5SnlCT15LlmftuKzs/Xxh0aOXpVaKbT+wEu4ZpMOiDvbLmao71t1lPYqHF/FSID3wXsIQH/5
5/tdL/RwMZY739WN0uqzUKmYRyOTzJRQEAxgn5wydfa2COvDo89ZNk8uuNsesftef6TcqwxKLdTU
HUpPFttDFc8Kr8kGZSMlcw8HZELl8CXGU/evTNlqm51avhtoydPYz9A0avrGfvcEgoGdpCZZieUJ
8dP8msW5iOOiMRSIeT6Q/FE9s09DbW4+DLuCTVzVLF1/lHOtHYqeZGlnKHl5fmWP4T0RRuZghZD9
fx+/Q2CyxkuN1Yh78Iacx1t1AXt8snqrqw2MUEz1bVWGvFr5d3x08pHNxO8Z2znCz5u2jO1V81QH
cZhCUQKZQKSd5jU1onKyDBgVS95pRJu6J8Dl1u2xBHdXoevf+H5wduDIicGWdswfG9tc1KhObr/B
KODM5V7395J0iqNGyq3Anrl937vrVlL8E19I7zF+Tfphi+TpXky+SRmRO5xpjv1LHr/tbr5WdCYZ
c/fJYcwGOfI/PGPzAfTK3iVUpDHZuUOsU0lAgiSyeNSJdcO8jFNX1gpUrqoTWbobHHmHtKb2rSLU
khZNUjGasdVNl+jplxXwoO5i6dV/n8QlMqKkN4JSGvowNZXrlRTaFrXK8pxuPsq844UUwKKS6qpH
+vjO0kl/LH20YzZjd/RRtI+cSp7o9JKForNIytbTu3c/Mgxr+dPrkZ+Ei2prc/u9q6PlHHt0M1Hv
oKumSzEtP9M7kklc0UIW0vcGcjJul0KUBKWbY6XaNDNJvSjysa/wSn3r3mfOtEvaK0Wr8Szq/R7M
TqLP+FtY26+ak5Xp9FHxAKG7mRqxGNCqMm+sP0g3ryRcLhardOBLgo449keG2rd9VroRXcH2s06q
budLyKFvt/X3L6Jh3TNeLRg4st46iHEX0WYwry3jt3hsV/1LwLTSS/CwLnPgacDPqnJPehDXuVxr
fGtsUrBN+KfNRanhzLEDsb6dGLIQ+cslBlfj5omattz7OiD72zhDKXWyyh1ZdKfUE5uYCWCquDxX
dbbt+z9StWdshXYSSPCfKtjHjbSJ3tCuiemLuoIu31pcnixYGeml8wFfPuhUXskbYHPO/Pa1l9S5
vIXhjOu9joEbkp7m+uNWh2m9TvH25BvZ7L/2Z5BJ52AzDgOAL3ztYz98B/h+YYGgvC9d9Os0VUGx
sYtT5Sdxbu90Fy0TumNsd/zvIKL37/49O9loxwGzzuL9W2HFE5F7Jmlz+lwUfJ9kMVaokdx7Jl4F
CQoo+jBMs6eCWSw/gfb/NOH1jnuc7JvNVM75t3NMONuKNfJvbu+sFARB8l1ZFV7SdXCczEzNyy7a
tfhqET2QhwIJd7IZQwLVkM3+sp3Q+0m5wlHS5+m6hBiRz1ogeoi6n2VQlEXEk2z7VKnsvpBDg0XJ
g8Gwha4COVZgJmBHB/AvqO+AS4PXa+0daLKrV7f/7b714fUaAL0v80gKMWiuYV3nLPjZkPWfyPBw
3LFOciLmGHOrJou5sqSu/lJHG+rcaK9k7OlBPrBDsFYeEg1JQPLGcYF2qm/XyzV1gQ/jGrij1TQF
ey1pc+6EayorfNdWsXGtbLixgBHK08TjBItE0uAnGxgJGIKyJI3fjyJ0w56SjQtVM9w5mJL2phum
Q5bAM6409E5ZjgATnuH8v3ehIR4ObRSoYqPnOQ0jwzstGiLa4501MC/+6skFYQu3hnZY+JclTttg
bEffAJFK1Nzl+hKOS8W4TDLMoDhCiubdmnDKS2yGL3N0SA5LVxJYw0Hj8uYDXABB/Sw1ioAjvGlS
/0oI+eWFPyPYQ8BDJeTRzKvHAqdkFgmccUSv54jyTgZULxjW41Go+sG5hFiK6s5nOncB6cX7sxS0
Ncmn49qEmdUAJhixJagyaiLq1jF23DZO8WJVc6LfaQjGU2mtmqHMWGFoDU1tVoTYQHd2cJyZdZfW
7dzztlrHZbUsV/6VqzFgfAx3feIB4CR+clMgL5mP6f9EiOJ/6QsmjDxQ45fO9eNoJet3f/JuwW84
/uOi3yzYaME/qm+gEfZxgdtD3DQwqChjbc03YWXw46lGPfInesa2JEzCB/nKaKtaXlBASZahubN2
wNGCzztL5HIN3xZxM/nt2mc5XW6R4IFNvjJJTls7BVmccPgx2nL9h9DBLCR3cJe8a4MX924hovdy
uMUaHTatlQi6EnWeCLi1/3DeBi41CnyI22O0whimwOQVIxa8cF90byiIA8O9G8cqoj8Erv6piHsD
7PW3OSJaEnTA3z/UQWzR0ETY5LLtILEigIlEyoGetUN0RZW+cBVsplXN97/GDv2cLVX9TK4NRV/q
sBVwuo+/q5ke6Z7vF7SbfrCyQd5KTh/FvInGZr83hz2ZRATv/dJ4YVvb7SuV8RxCHf0440cMZN3O
MteFXovmHTOfUE83UGXZ93u0/vrgUuA44+X0XHrrzQWp5NCp3FN8q0r7tbE0R9ARWkDQfZNzsuLh
6K8QlQaQA1Oz57qLgDwj3moJFslKkAqDjKrHrVP/coJHHcZoRsj8+eVvwcQh1n6gJA/bCJkRy/93
xLWuJP8seZOKL8hv4VFsSXvkoKet7NSqAC37eVjYSjeykK6jVey6wo3zFmerqGssBz0Kcgg8U4Pj
cteNJ69h7iycGSUQI0DAqLHrBQnExx13+V6mCPXPjHUY0adCuipIVU/oGFD10dehg2dy0sjYxAN3
ftdRagr7Vl4FuCpBnTvHVFsxgrgzpu1Mev1KfpCPEMJI8Jr8AE8V0qEaksuTB8wuhsgOZLNIIZND
+xcqupf9LPxGs44d1/6XMeBJCNrFpLtzvEeKKWyqm/QVLYaGuIIakbqAjxnd4PGSmjYizBiYEpY5
JR2yPG4VO7z4fz8mfteBsWW9NlxBoDwDN2BGQbLtXgOygs0mXg37zup9hgAIx4vtBwq6l143rwHF
jYLGS0VNPxUUPerd6WRlY+pkP4UfD/yx2Vp/DjnxDuvQwrkBNUJiBeuQXNUwUaeoO0bnhDovxqXN
K9Ci2lkqJ6df3zaG2YVRIlP77ld0uyYmgJMQQDezsJDE6AIVLWv/yGh85xr5jbqWQlwi0L+kzFyo
GoQ7KMrWMpk7DyQdtBqk3+X4KWfiXGv6BimEbUmzPmaUFy8Vwa4BV/zsAfTX27BrVJtM8wPqsEta
fBduUmC8RhOrumzKhAa9OBLn3kAQJemMGsTZ/VjZoMbq3X6U4V+eekEFFiz++yMcQh+vk9PLXqzk
4kMcXHfSpXTUKoLruYkN9+iLWFjPkaryMG0tpHy2Gv5LaCqhUtohwHtu5AWv/XR5C9VfjmP2hryC
fv47tuzeo/PLf9wSQCdVoUnkwIvPHcxCPEe3snzXu9SrJtYpC2TsLhBN/et4pCcCOTdGEGU6icph
TLzD6Wdrrh6v3FulWeLNSKj4cTgOnGBsZAqOoxL+CcR3ZmOKmGjTjnABOgPsnXpTK+TKXOlX80hh
EZD8SV+GQJA5AwMEmLLnbz0rIYllp5IE5j0b5QDCeDtzIFUoilFkkrqCSK7hHmXtqSXdEYbRtBPL
tlx2WOevQCmGB29UqiI3+BnIPKDxB4D5d9YCd0sBNegc+wTrBEAYt5H14srk09bgZpKfK0XfiNvQ
HAaaWATDsEwxvNWZxOV11GH4MbbQqQF6J73pwJP1JFz5mpnjMaqr3u+RKcgw43IcrQ6TjLi4DZEJ
7iEZlHbN4LO3IUPmXj7/5eyG3jXGjqtVU94HLdbxun2Ux3T2q9aOIbxky5C1gMdwIKM1zsn+lgor
sNmge4372MsQjEEMYdkuqaVhGDwAT3ShLsVInExtb8eN5sZi1YMN1V3s8wiBkGf54FWVSIAkdckJ
ya1Bm+vAWKk4dqyANxso8PQmaM+vthrKQwBocTZEzY7ASGNg3p46W17ERiby1L49DYgmUF5J5XEP
uyoEhrRVp8GMzzWfcnA+kVbd1MScHXhYfJfwd9LMMieIBMu4YRrE4ADe/VGmws2533vDD39Ao4uB
ntCAbEm7eGgzUXuAjyXXDyLgUlqIgqrMG3NylPIIt0yjX7SCMyODdarUmOpx4oKKdb3jog34NNLO
TZanyRz3H75vAg9TEuNBRgwDHfFfphrWnH/pfx2cBdUmquhyyQ97a7vKgS28TtAckqGYKpqwU1a6
y/uirscRC6bLzNePXDJ8CR87q/Vp4RtD9E9ycIQmiNrsBWAq+KlZ4i+N83hP5nBo284ICg4ezzDH
OK/2j81ZG9Xp8OGtuVsnYX0aKuDh4DInVqWtX5FQj+PJXTdSREH4GnYb8jYyTLykJl6q+dxhA6Mm
rA0HCnIXXH8TKqlFOOmFAo7C+T4HnvHrba7m+JbFu/N6axaFlgfJJCA9rTIFZQu5t4O3GeR3gI6C
5+trupzcwM9RLmAhAcNbvfGyzl+P9icDQQaADMhNum/CQTFK0DLcVTHk0pVRALRljwd8QSzt8AQZ
ay7m1Bbb8/q6D0/4q/LvgyrBC7RTEOwS4RIXkwJKrblg/jMwdwxVcVVegN9Wc/8xeRKh8vQNByFe
S8EVtZwQRVHwdY+a1jcQ8NBrHuVWVvedyJDqmvdGyEzK1NuSUV1exXHYboDHKkZFzzza0lKRDvmx
3eEaoO0KTqwRm2o9bZLpKfZ+n8sRoQDjSnQQ48SrAMxMpMdTsrFyxKFLpKX2RrmUNCSTrETKi2KT
aFVLAyd7OEw8DguePgrGyUSL5Vr5oxkk9thxpmSSo9q4TsuT2dQWLyal/nXwRbHSp8etEx2gtPzy
RPFurz9exOqKy8UzGxCuwB4bwtwRUSB9/FVTBwRLdbUF21ykfshuWy/gtd+OeQnmX8Aasl4Me/va
tb2Z9vTduPut2fv6PDcyuqPc5WGwZuFTlQpgLrXLi3D5k8SaCottrtAmsbtfpBArgKgFUOZo6zHx
AGJ+IifS8uJFNrUEOxeOUxd+/GoJ4ee4ZZSU+xkXqP9vTmA56/arSnSakk3idDhaw+A2FIfC6etg
DBRyfbbXCerkbn3wKjI3Tv8ufJt+X1gRO9L39ZRoCp/JqYoMiBxgk0qgJ+Be07S3rCe9n3EWeUJx
OxuYO+cpoL2pbDqgQDFLG9qcXHxUsxc4fhfTF/TWN7SKItVDSLWwb4K57Mo29NRT3wE9coYNG9rc
U4kg0kqR3Z6QF1q8fDxhQ6tCouDmyXJytubqrdePzxaCx2XZ7h+/QdO4Q9CmAd1yNPTOsezOZG8j
yLa/lS82/hvft6k7lCTnayQJYfF/VQAD5GOy/26npKVHURbkap6H4tXMjweXHv+eCBBk0GgzbEiK
Os3QoXiz3gTl3L5QZRX+RqkKkYpw8yJS9bIzgi2K8Mbp9Dg4e8uAuu9DLejzoB8ZwJiKhADteDVC
pDIoRzJdWpBL9sU5v960L4Kw1japfm7oMXTnmHiE7r3uJGY9Zm2dAIP3frMQU/q5OWMWRK7UcUzc
zHLYsEzoTaEtFr5Lq2i9ZCvvAk3GyHi9qahAG9eLW+YC/N5I5TG1Ac73Nzr8/Tp3eS47/wHT87oI
vzcEqEDt7XAtolQ0N7TPPjOr/dXVMWlWg1yeTzgSJ3y7CQ3eT09FUlOmsaKjZj4m1RP1exrAEU3w
Epar0RAsfKOxIWDWn+4PV0xzI0vh5miKqDxV+3nGdDWzEK2XZzgREP+1ujAnorhUZBTg7T1fqeJc
QAmYbaTtZeLte0Kt5E7lZCNrQqJ2Fc+U7h7/BSVfq0sP5T139F9WE7Ph9ZI2bCCH6ZBWfyf0TIpr
K/Bk3Q6xqxLe3Zqp1dgFrKDlTfEJVS6aAL+l87lobEGtCA1x/qgReRwKLO4AwHWBsnECVfnNnNl1
RGbvzGMVeaIcDMceqAUt8TssfpsbhPEt/xHMrIZMeblc7xnZxkXOu/FQ4BFENW8FrJQCbzz/R5Z/
rUyPQaT0QkWxOZ2Rty6yk+6X5i1UM8gZ2fsYvxKapbe4EwILHWEt0w7kP1/MPo6EppL9BQIusLCZ
pSdhfhc+8Nvherf6zBDpTto5Eg9iTVnZAp1W16gEyIs/7HxdPlSRnSOD8vKu+Q8mbfQg8AQAsS9u
yhZXBU/o2iARCa005Ge3nGvVoC6l7WLJZYhhyiWfSaopPu28O7SFMW1Qx56HWUP6aqbMxo/OrxIG
2WRRhDIFlEoUp1T+67I6qoXxo7cZFcFHsBWw2gie0/xR/Rx1bjZSHyt1EAG4/mFzO5YTYyi0CLze
Gxo01S1vr5SMB6ASfi4pqzzaxScaGGnjamGqBs8M5O/izjIJ75yPJT77+7I2NLKXdNv5cohRvfTh
JDU6w56p54XimGy0FKjKuxeCsEU/iUFL5FioTOn8V/4rgX2hMMmdK3q/VmaU3wy3tBEQFaIQyKrf
SToKyfTiVvUtOsdiSfBByUYQqErgkjjuyIdjdiYMe0J8WxnwDij9yqojmuRX8NrydAyQBXXPuDmM
muh+cm0/s6NPuFW89abIMdBo8etIHZZ74YVnAlJDumdFbLvL0MsHfrb3nng9pqGlGP2OSlgn13Tc
lT/Emkp59VZPmeo+BZLA70w1pT0pH2tSb62h7fXA/TK6bL/eQe1H+UsCwSmk9uR6yA87vXfmdmRW
tsRg+v4Eujn0eQEgG19BpUlndmItUKUGh7MxnJe/E1WZPUxqxVZmovT7DrFuGXVO0+e50Gwc7yfJ
ody8kpeUKYTDXIAy3rrPcaCSi7Vt6KQz6aVeQpsP+emwahZT5g4bLhEnNhTNL3M4LM6FwiZ9fPnW
Gq1pLVWy53eBC84EudFBZqRLu6VrvnLLq2bWQdwTNCAFdK+QIfch5nH/e2wR9BhhEMAxOASbMkJz
aImV7WEokTp18QLBA+1Cp0lis9Bzdm79VOsHgv5OM6tJCv5kVQERx6+pH9xnyFaImKwRjATaBOYN
IW4taJ/+P4PntUdR4PaAGwF8RxyU/InxagDMRSkiutbckGZ8/l3ZTY5M9zyo34J4POmI9pgCGF9S
WMjnQtAZ/ZZ7JG8n9hEVyXulUFOIJHaanc2e8TnYR+rTEz+nDFds/6SLO+v/8QUw+VITfwFAbb7z
v0OEiY0Bs+PluoQ4wMqMPBfMDAQXv3E5G3wkVBeW1af14ZOiiYWRrRlKIwHXG2UebxpdEqj6Vsyj
axbHaodJNSqya2uvuU0cSn8xtYEqzO8XyNC8gBrycP7wDc+xb8ANYNZYus0n9IGeVQjgvTGQHSJa
5057j9zb/tr+CUv6u3pRWa9dsF8NSAPlQerxJpZeGpwwdArZqCaVNAljyUPkbAoPfCHLT5Wk83Yq
n3AGf++jjYBiSDie+XWw0RWhKsm7oeSfReh4dTHpZczxxf3VHYzXmPGXe6q7sLXqNyLU8FbwIt36
qoB3CaucENpM65dKrsrbNDz3voBMSZzPa+0CWEoWOdVZny+a2grFBNUM95LsnhD2DclJnaMNrVNj
WaNhLLhI/bpvwfW5+DVrgfSI+gJqehdB0dw/xbgusqeH50Y3Qw7q6O8j2B0mi+ko+Th8xj5dpcbz
EQYFwQu29wZo74pbTrLrDx3x/S2G69HTbJToMifBAGYIfJKSQ3FW5h79MtvhBq/6EpVHGSkCIcYO
kb8/JNABcMlZS/k350XUifjUHaIpxAWfle86N2G49oZjebv49pbX9JtU1TwDGiT/0r13gzhHnxnR
w27ZGSUZzNL6/qPgCiSIYgXioc/ihIJw+ZXHt9Z7tBJE0oSp0M6kWTfG56f+vfVM2VwyAu7NDmzu
rfqyR/mkaXOfxW6P2r/dErgzY8VDuEIgTJ4eutx4PXdKXMHXyidffnWHb0yJbiQDyZ8q3Lk3CCOW
svNnlqJVn8xSKN4d8jzrwIOCDVpp+v4FrVjvI8mmZK5844Phbmm041FhIcinzUvpc997BMN9MKt7
i48OENmMDAaurNUbz4PAoImDjsov1c47pkpYK9qrwlM9kdrJNM1OpX3tHSDbDBJigaAlVgWFaz1C
WgLKthYwbVBYxXyfw/M9T8LlS6/es7jULTVCV8eCtgGuqQccyLJVVeuh7IDDH4abC4ZAY7tq7ZGe
T4A/Ov0CV48hcBDGeQ8Q6ZbWLrBDk28Kev9S4sk9IZBjtVV2O0YPaJTKZiSgYcA6PhWQb2pPtOD6
OerN4fAVODS6ddbXikd13WrDxt6cFhYdOs0dF6JffFyvIU9ZoZJ8Yaote9xiob8xWWUAFg0h0P0S
Xw+SPxcsbKSqiGSMQ47LoGXbKLMFuTS4KaFv5J/fOzsvn5W0hatQ01dZ4eqRuhb4LXgYH4MTlE+c
elwqxxtl4rkpcLPYBpkfdnKrKMTzCUpbqBluW3MsSYank6GjI5en2orEnce9SGz38DaCY0SohWVT
q+tdZ6CPwROLRyQQqFAU8piKLQTiDWyUrtMS67+ohGNe0UQSaIRTvJUaHFXyUCrtM8cdsJiSba7w
rXYp5E5dp9of/SHux5oH4bzoC37SjPFQuXT7Opbhkzujuzf6+yHM/MCOlxn+WCf8qVhfwVsjSw+A
CklHoTQLwMLApMopLddnWlVPzcdLdCUqShbD4uxLsR52Tz8PWTILx+TKU3NdsIYUVVg1n4wIw9/a
sDiF0nfPmawSAJ65T0hzMAkvUtct7cht1gFlsDMh+gUSr8fKBe594r9n8uK+qHRhfpCgWFF7fdbF
CDgRxov2NvIDuWF/mFAfsssQC1LqdbVqTps6kqKAH60fJqxOCaUj0p+xfyKV3Y3j6KBO/i8Whm3d
+9ZgXeJ2XJvRfqvZRsGdjPEIkrbMI+ZgYc1/hJo7vaasa155DoKBCnG7XihiotwGd5XGZTb0qcPn
BguN4IybBSumlhdptUy1rpbwu/boXDbfx3frUSOB6ggXdBLUpXSdMLOT1XigEQEEVunzyu1FdGvq
ckk7/Dng1SU+rI2Pw0Lf1HwXINsCZLHIb8Ot9qJAwUJ5wWLuK53dnuh7ze1c/N0CrYQFq/TnCmeq
DUvtyOhXetdh1DEK2xdivjmmjPcQRtxvLhhNHBIba/m7RTTPaugP5EHMHBgDH2B+lk0sGvdMBtYB
iQvhfmmYyzaXd2OTP3L/MW/0iqwXUqjhU1eD61zOl0QzcDuWj8kJnWSK/oAc5uHjZ2BMv6lvff06
v+o7jORFoKOUbShLhlziTSqTj0x2MxhCd12FBMq0uJPMehK3/8l5ZCeRAqKLm9XwRnDlwQQcKq5u
S0sbrudP5P4tX5LacLkFlrUKU0peNZiAfIN06ZLYCfbtFaFTDDCh1Cpuaff7+xXTloE0+nATofAw
Gpvlr2UKjnmAdAtQlcN36DpECHDdoL4rXmFwA4i2Lwl6egGN0kkLw9mFXCQBS6iXhuRWTScCBjw1
i23un/Qs5K/PrG8GiN6s6/8HFmLmN1T0c5x98gmnRhpdCVGYYNZd/JHPNWY2Nd3CbNz1Trc4aKjF
PXFoNKdfj3ceX+nufhbpedbC78guAYPRsjtLTOicE/qF2ovxY26V0bUNQqHru3O8cpj8ksGo06Ee
UKFZ2y5X21igAwFcisDjS86qRYk0QhFeMg5o3c1VQgFU3VaKT3LY6B0NWX7lrn7yz52UTmTwjdwa
C8Eg6Vf8fj1nJ/BVTtZODS/8+vXQiFWaLPONU8bNLfjB8KjmdK3OAmSn85nU93W0vrQU/LdFVzKv
C20aC5YWpOePN6fcNslLOqAPWDEZ+3iQjnCyRJabKtNF8FGenR6vCE0W16B0vXR+RP9Gt9F+Qc1y
wklk3h8rgpi7LyuLUXw+pvVMdxrHmSRBzRgXQQ6r3O9hDKTpAggu9C/7g/xL6SJXDoHaOoM+ZVay
YwFwkWSWLJokt++F5lPet7do9ErcGHWIBBxlEgSNvaoeS9Y8SWo5OowJzLTCpJR+Beg76UeiNON/
uCZDNH0jFwMgKAmvTs3rsL0b6kdmobysDhsBOyZGtJbOshLC7Dn7izFvoTNhGX1KNaBnTACOX5Cj
/iv3d9vAaxp9TFOprLjqrjqRYDWKnQhSvFb+c2hBrkz1QBx/uB7hm+bxErJy4ZCQbtXgPehajUbo
dCLx9cjNKo8zzyo8u+KLd9Xbt2s15oEK+zLaXQHgC8m4W8ao3c8y02RLdn/d1a/IzSPShMnX5suq
KMdrZgzPjZMhl2LvfyVlJiBZP8drusLHWRAOvlTyiTCNXjv9Fdidlum2Q+FxugoNYO206mCBOpjE
5gz7v3UkBlzBOZcmAKeSF0MvH2nk2A1YA2z/WKBvZjirUXDO67hq6sWQudfmtteNTFH03FQo5Gw7
42UhmDSRuEMlJrd0LoLdzax1GsFCsfHCR8WYoAWGW0G6CAozxnij6+zHDwaC61OEtSQJlt7OFZBu
c+pVw4L2SaAJrQKLvrF3fZc7sLxsepFlKYAIunn1oJbnLWqwEObFTxCL7LbqW40PhgpfQ/QYRlsR
683WNcT36coa1aA+nvzIoqcCkGzHbjC0GjWm4sv7NxlFPFPSOis4iPBjxPp13x+4i3bqUYUNQybV
AR90ZvQwgkKJ/h1nNyORtQfxm8/J/rNZnRrI5CM8LCT86aFQ5NrOahfLYRIC5xKdRdl4gCBH/p/D
2mfo2kG4Uzry8JVgq6aMzCHIW/mQspLPjDqHQByL2VIRV/CoMlXyUpd+V2yWHBb/qrmDqvI+gCEa
QS85N+ZbAHG0FAVwJXA1LFqmhqVP7SEqPXuUjmbdxpBauL2lPNOO501JVZShsHmQVBVT5Ad6tcF5
BSH8Ma525znhwlEP6U1fY4cZdjAeOZCCy8mvwvs852wTfSbjaktBPGEhZR2EC27GZMps/BnFHdYp
oHh4LicLPHoaHdzkI1Vm7snMfKzTt3KgKMEe2FxrkR4Ye0oZt17g59G6jjxntBDqWM3hdB/5lsFd
exll9DszmUTqpm3wrJ0E6fHAn1cF7VO0lpAe6oM0HPyB/w714LmKJ66SOHUrc6VjAOKCBG6nWXKi
gPe23XURcTKmAX+dwuhZAcyn6CrtrvwA5mAVXlRvuFPkBSaUv/rSTruWY8isdXjtiAaHgsFDqga7
7RUiuuppN+GTaNJ8kX7BdZWlIQKo/rDCD6Iez0tv4vaU9pS0S9MXXZhZBEXlvpRE/pybSKt5AxOq
vZkdWeNQ7G48tEbWd/3vk349jLhXlUZIl9lw3n8v7Bz8iT4kfTI1l4eACRJ4YKWxG304aoUYwM38
DmHk4maLrOr7FtXG/ZkfiJTgQtlBC6xdO/RV0R7R2hiDM9jJQgRqUHcqnx4o+oti0lfvhUE7B0+G
NikCo10YRDbMqHMsEqgthFdBSd7E+MtU8ZXzF1FKICVpZit0EBO8DqUYRnHO0FbQBNa8NNgDwTGh
lNe6mtsI+3TC11EqATF2+o+HhK81JcweLpOKPZgK7Pn+cBq+1laZ0xi4SFTC0cinXlqZpk4JJq29
5bYO98Y299HAw7CsLl+kBRk4QpLXK617abE2j/5xA+I56ozxr3AMiGKeA72MGxrEj2cJbmm5U4AV
J4JqrL5V6qkvZ532/joADQL3lbyOhDXkWiOmUYbcxJDfPxmx0tvSSTbzJfN43gN/lFHLIQ3TiuBs
9OVK/sSnPWC/2zkxnHGmAIhZ9cENMJOnUSr/R1xy0Gbm5tlyia4OK12T7nXKn3apdfGOyI7eXHSy
RqJiiaMY0rA7pAxWndwBNI7UUEgW1AlOUd6+qvYCFasbt458tbciNSUnUYjDvMiHRqUteJXjzlnn
ra2x9yVmeeUOMfc9o1z4xTrcmxVXrB4tRMpXhB1odHt8AP+OCahW76qF21QuD2ulVEEWWtGUV+7p
b87wk5IN5Kxzn65DVNZyN5SWFb740z3Egm8LCxg/mC/romaCyqWiYgYTjwxQlOSBRL1DrYtAvyOe
u2lWBerqGB7P6r9smQdWHJTUZ906atIOH8LTuSv03lIxEzaQ6YlQxaPTPlwMPf4sSOjp4KXJo2TU
Y/DG5c3fCWWUbBzIE/F16TQhLBFqZkwnseoKTi07ObfYtMV3cjAtXkM9nXw5wSKHGWZL5vDVwMf6
D6/K0jLDU/BggofqQ0JPkgofLY+PTxg9weiJozwVing5mUraD09iu6IVJQGCuO7jECySJZn2AwHK
rTu/VY8nJYQs5XeOryLeQv130REhukAocR8orw5NOQLUjZ4xIXQnoqAA2UYB6fxb3h/dK+ItJ8Vo
bOvIlHKj7+ye8f75mbRJV3nfHJgQAECA5EMdXgAjLiZ4JcBWbQosSj1GqMUFpj5Kh/+HT1enaVsi
cMku7+SXVE13jJTF1vJJpJVcszT0tpKx+VRGO/lpMn4eF7oi+cszUCo66CHnvKIZ0VrIc3eBxDqd
TPi9FKVGSzIYCwK/68MGydb7yvUPFLyBU+Qs9g5KQUytggVhxwYPe3nSoZBGC+Ge7g6QkTQkzCLS
qMQxECvBcLxehx4iEuKoGRNh8vuqEE2ha82R4LV8cXfVmPm8ggPS2yDpkUhURROdz5Qhab9OpXix
geBaEQMC/j5YpYylvnAl9dblWg5+/hK3ZiD2KmksLTz3oUSZpqHs8f167uBBEbuYrncZ+Yr2Rhgp
310m2iMxREF6xZMxrxQUT8Th4hbQqvHHF/iOrgvR0cly37LnPXmaQQrFGWcW3fll1K1CgQ8BA5Ub
FxUTdR1U5sWCpNjCcKRc+1oxW2gPFk6wvrWtHBZbcAPR23x4KEgrktxLppQBtEFORzZrT7mqfOnT
VcbfXkwNcD7LK3rtM3gVSSQJPpI9SjDIsmEgksbODrmoHDy7ouDRhGAWw+DTDDsxrG6+TUP261rd
N/n2GoW2bGtZ2UC7Ec1RcB9/8Qx5+O0FpxmGdsdK6+l3/YmBbLhWNL1yh4Lejzsg6P2xNItOLosw
rdRyAPMU2VQBX8mR61KLu4wFbNOGUWhe42RArEZqipKdKnh2WgJfvsjofMAHvLS7MoAR3Tf4T/Gn
iDFEUiN/3OVPzKw1N0heHGgRYoyPHq0zdBnLVm8yqWGwdmSGzT4vUKdBh6JBYmScVGDzDTGmSHZ5
i0DlPgMsFZ5zrfLu+zV9Ghw8mXf3GPX20Snbxch5CiSfzIIGTYJhXjwhKDOEAFV/jyOFm5d5p6lB
Iftf7aO/Znjqhi0SOuDGGsHGUU5niANJeRJBBGHZ737WREHyWNaXS4FA/hzp9FH8U7S8uoVWKIpb
D4xVxOzXiNtvXI+S59UB/HI7wDHcJnASBbfhEPY4Gz6WrTJDBb3/lbBoGLgB+237eKV6TTccdDer
pFkNO/A1LzsM9/RzqmrUymFAXdEwsYWNEx8Y6K/SGhFrQkovRMleHyqd6SF2Q+1XTa06WKAPFJC9
gpkMSfW5CY++EYnsXurxyBgYHqOP/S3Tiugge9CesibcjP3ESoxvW47FwNenH7XIlbbzagc5Gb/s
uIl6ZZDC0Q63kxz2RFH92TWv99H6tYBVVsDmJ/AXWp7ERn2rffP1gEMldrXssOGiMfMYLgBLc6EQ
17AivtEFDk0ML1WcTR6DwSRguaCZjs67eOaedM9hrMaLAJe5Sh83OkgiYhOnG7HVfA41PHrjU7/M
u4NIDqCzjcFsPey3iFmElbr8j4KhD1wK8ln9qUMm1p5nvb+2FdEKcJgNzQ8F2zaYytvenQehBGkW
KebFRoiOLlBYvj/a9KT+Y7G7InObwyWiWmOkpTnsmhPPJodHwVANOQLLTmI0rFIeBUKYPvLZoxQE
qb3FIhBEyQoILDdSlfYfbZQB+pGSwActJKUg4cNxxc1mxVbTfDNmqdcj3T2GxPge0RN+DO2Z2Cfx
sXUY9/GoVjOffaO5Q0dbDUqHBnItIoJFnBcQBbV659wbPwZjycCLUhdxu+dMBrNeC0aeVWAPXOOy
oyctdtLE5LvR/Pp/2GWByT0e9b+CGNyr/1vt9XdB1mOizKap65fwWW1tzsOYLbbAz1ZLV5RweK5x
NbeZ8ga7jAIoSjADziYiZEskL8gdPw+R+eFVr3/t7UAO8ordz/Sb6eCpqAzfyFrupNqdSOkmTXAc
D1iCKy7g0/ZX50QK/7xMM1RG9kHvXQZmBVZ9RPqlC+aU45ZqcmLcGsAN3J7g0/B4tDBIZlcRQ68E
QVGfqkjjJPGD/0yzE+ldeGQO1LvkKzvIV+wTwceLWRse7PYW+nC2R4XdBcc29GWO+Iv2Vlxt5ZeR
HvS2YFC0a/w89uTeQnj2L7wqokehc+F4IOHHxhEF6FiDPXbLlPepuG+36p77O2y4/WQ+1CWMmOms
EBFi8l5aZPpkI4E8QYJEa65wxPqmpUJM6FbY7hF+lo0WS4V7U+VfrpuU8RWRRYXQaKwLGHRU8WJY
L8XRSaVEEk9IR3xHpEcnwKcqqSCL2OpCOTcl95ADdnWUgVhU/JheIe2DDEZSqZWMUNWk3heJVLu2
acaTh2a4GcYRon5so2lf3RyxspQP4u+BvGOWhgD2W1UljQiLdKhnQUNlx0l7OmSLnAXzVDpQm6ev
Aq5UXmWl5kUI+WsDFvgHWLOUFgU/aRSXbspkF7p5jovqcWW09D23u24f85H7GNJj0bRe69SF8KVx
l+SPov1QasNqLQdh/MYpynEW4Cude3rJ9cKelPVboN2vopjl9FfxXQWu7cDSgrSdHgxdOX1KBbfO
dWW0CGmLDM90iGNaV06uRFDGHULiI+io932BFVhjAVEWdmEIa/G1UWEkfqL0XqH0TUwki0c7LaSz
tw9NgaLT7yOY2ykAVAecLFfHmN83pjcbMjpBgawnGtdvpnLIcY8R7gD03DA8PuotKooXhbYKXKqz
y77ZY8KVCQtTEQnE+KiNlu4zSHL4cBCjuPPf95ni05mtUFAySMMDhjvbYDRG407HuLkEn1iPe+oQ
45pg5hkwpN/eQEcSyyMGk5daPSC0aMeuC+WBiORzQakqSJulfRA0n8jVJeg3mt28SRqRGD68w8Hx
z/2o8UUNu/Sg2O0cTkq432fXhEh6tkKcwmgttbTP0B0X/fA7zqYufpfpWQMEHjpDDt2o99vu53KE
M2OT3InQWmFb99dfjQ7L9B0p9i5sMN8yaWtmN47pWiFB1rZeFAhA/EyXjT6Wp3Vl0pUlxvxANJQG
wpv1jjfQniMWfoeGwMKRc+WH0w35Iktmek9rGBj+msYHOfwb5fgkXtFwJGVr/52BwG7dIYdvtGN2
dPxEVbvVqIYx/+KpiWKT5j7tQMPvWDZeXOvc0ExEavC+K7uy7bCRYejn4d82WLbhr/ezD4kLwalt
AQsT04dp8Wq3+IBn6yALySJXuN8bMTfEJy1EfhFJRJFCa10UHkCitOPqDvuwRQYKfb0FVNIgCfNu
+2x/5FNWFbiUi49HHotuI9wF9qAsla36jR6/YrKVuK32GE19rrmX2ubyOxEQ/A/BPUEzGWjpNA1Q
3xBpSh71OP+z3E9WJqaxzfYUdOiI24dEwxUGvi32bh3bAl9P37ZrJiDDBWNrSBUaQqVbyYpgbKXD
omwdBfiQm7OdbUBkOxOy1vSyLfH6FpO7IOEsrLznV477ONq6d+ADuDbI8af035zP6fXC2BUozRYd
VlUaVf1c9eUTUpBn031edWMJao9qU9TliOWy2CCkXCFKokKZ7jowdlm/e+Vq4+c6w1xDhKFnDpdy
pPGRqaMPSp1iljE+fBAZDr+1iNI5oJDsC4Y4ENbggLYmONdeDKjXpFNWSYP34L7VJh7KPahG9q/X
qkWJL2t8cgt737ylO02pamt27+HirUMeV1eCw9eStXu8tpXluq2p8yrj/C8knxrufwi03A/L7Pcg
836zXDLt3oBS5OW6QESZVYiVx2SWaD6c+N1e091E9XFD8nG6YIesejcIhaXzj3Dcyeq1LWb4b92z
n9NxGyhzo4G792LB1I1RScD55tYqDOa8bAx5k9eYZ6oQgs4AXO1e9lugfH8Vs4BgwuGERC345Y5/
1sQ0CI0FI3cRCYY3hUjzndu6fJ3s9CyY0869R9MZMuB6kfZ1cbdFbRmfoK98sZn6TYeCP7/WqH7f
6ivOnkokPlZxWYHuPukD52c6LmTqFO6T5r4WSkkHE1P8dLtnYQftcGHA8sgUCdBgD/lzXYjtcLNg
jT+NH4DCTl6PMl91Sktfwo1YxSYUzM5I30xYTroPtjpA734HNazoXlh5DE5ytlHJaMEsHlLDB0Ks
qYfhe/NXI2f3+gA79zJ+tKO7/WnjbtqFE/gUeI0zscqlPm2PYTj1B0/NR+YjafbYJilZIhm5kJB8
2HaiZiEPy8iqQkVIN/84aC7yu6o+Npw1Clf5GQWC56VBOKBTK5TehvVVXSsxJ/VwbLRUBWIk8ANL
4Jj3OtiLv3kGdQoAScUPb4q+dH2aHtHAWZvT6H0Uo9CO61+pq45Y5A9VVZhkdGaY7+I+i//IRHwQ
ou+bi5s1gPNfshexpvPuyq4JtSiB4tUb+t+WH0EeUcRf3rldtU3OGof660nhjexs5xs+dVLVVmvc
D7QIBgHPaLiPQiemux5el57MT+2WwKy8SUPFJ5oRJwxVUiRam3X3V+tmQXUh3npYitNYcyUo86JY
u5hlpI3PAJsBg80i8UOllvMG8lD8cay+oGKEM3HaQZBqWycad2PqtvFjpUm706I2M4+Tlciw6VIT
v2VHHxtVDnhYgtaTKedaVY1mTSSPaNIeqjCSbkiEBdNFzs6Jz1+u7nVp+lc20mCOkhipRJ7q6h5L
0MhgZCckitsmw+TZ/pvmwzrNXe1MXwDyt1mUvljwDPf59/XmkGsmO+A7n0/E6YQmqZWKwMHPHweh
dj2Rrt9guZ/HkMLsJi5JHZrbeSzojerah6zpiZJp625N2hfxZQA83eFM5mEh+Ur6N+AYnHNjPW6e
iYyeTrocqv369pdBksbwZP6pC1t/mzUD7DhHZx4L7clU8SSJzTRoZgJ9++Wrtp1YY2fDLgo/I/zY
gdyaqjNtaTevm3/z3gbINk5LSz5txnZbnjWv2pvq85jlVouC2e7H8siAKdKPFQ2LbbViUl5MSy8s
Lr21KKMvLT0R+qBL+P9SfHn4CCjEeB47kTi1zmixoZ2rharApmKTkOKHeMErIE2TWLfCsToz9o+v
BMi25xZ/wMwRSgKQoC/4imTbDf3YmqMmHxk+AP5hvZsP/5QznQJ2uOjvdtPSDvASfAs1VIYpN1aB
GlKp+F99OB+U7Axzy5YLeV9oB3Wl6NBbipDbEnvbnEaFZsgg1sD3PY7s8ohtMt1bt5kVWYDDL3xa
yOy1UTDdpRYqK8ag4IzWyfawSjwqFWEEnhS0pJ+5FDzhkWUBJCnC2fEPyaLyJJMnFdnKAlKeh5gB
HIpoffKNYyBsn3PKwsk04DNKDwP++ATNyv2KhaGML4wIXNXrQDUEgCezA1s5EjkG44mecy3qJb7f
Dw09o9ko4nIpM70uRyQeOa6Bt4SFvg6wyfDGo5GDbbhS7ori9z7LKaGSLR8xhtJGJSpQLlDjiwxH
yUNDaarjWQSAdCUf7wwTVKmsVL0Ux3yDvjx/amHeaUBB5OqDV2aLlO3DNECOKIgiHGaTSjRkyyVe
XL3c1BdKBtIHUM0OiR28rX44LC3KU271m0S+uQ6NjReQIIAef+CPmJpWmgE1856WclQ05DyYyffq
le5bE3cyhCzn56jRFPny7OI26sUsxBfME4rzGvrVbh6uPCNF3sxbJssv1lh9KpHTEjPRs9ZD8cZQ
ldhMNYtYZSExkB3wES72XNwJ5esjcBMA9kX5mNZr+1963Bjhz/AbnZbkaOdOzTNnwHS15d+UG6ut
4XfQHDr+dCKv0W1UHQZSohdEOncbJLprMIWsTS2IQlvymZY8e/hHXu9QUKAx4ohuzux7Fc9l7tEy
Ku//ZSORtbgqTbndwXxzHHlTS17g/hapJoZDTCczem0v8AF7g5x6yYmPZFz/KRTraZMYt5uDnbZF
QMt7XjPH5GqYIRrp1mtQSYysz/oMCmqoorqCyWmtZFsOHqVjOMWXdd8bGb+MILilnJIn3/rNfFxW
bWpoM0PkyPwBY4F+3UzDbWqOYIQv06rr13dCioNQOX6n5n7EZQ8HjgkcrNFc4M1atEHeEu6JXN91
8OKjTOeHBAnDcE620uBFICjRvkBEJomqX/33b9B7dGqKos9JE0E2cEhtIo7o54/NmvOFOoMShQcF
7WbkQgvw4rO9t+3OagJbtnnuG3pfxY9tQ0EDtGnhxfRK7Mfh3A+sMBHSYRPN6K6vhXXJqxiRxwfn
FgI0Yb892Z8MSsx7kHKuRzu64Mdr9zHGxkpDMXKypsaUzLT+uWxtm8RMMUODjcIsucJIhT+hpnoK
bchmBeJgQc9U4m+XpdSdqgwq94i81QQy20b48JyZ0O1uMy42KtBYRu/mPLi0QjgK+LdiOmtHL0qL
M+fD984+3pUSaPAduMhrcjnWxdFSbGqbWI4mrPrRGLSByJV/ppq7c1+sljyd5XIyQLQUWXLNAXZW
FxdPWKUs8ghzpiyyU+SjPTccAypF0A6T/lmvKHzAuQjbWZIB4wehdMlVcygHW/Xcp/J4SBqoAoGY
g9ACYuXNwMX4tkCGdUNxB+/REVj5poAC2dv5ezptZ6ic7fQ0YI7X3/gWghRhby0/lke8PQMqILbs
iygz7p463qMrzFYw4P/4qsWEvjZnpcxIHQciyJhVfJ/hJ4fH7oEdGAnF1xsggYAxCm+tqj9LPmxa
QCWJfl2xHWZD0ooQv53P1tAB0v+dykgw9kqcBTYjFGh9Ukk1whCVfPwLvA6ewveW41FrOQFVIgdv
8cGPPIpuUdbZ8373KwWLK8yBKz6zMpvFCsvqdBqrjbPLBpv00woWdhztsX+u9cthXpdTba3wwX9D
A0X26mJFhkIW7qlyVgf+haDi68cdzWWZvHLE3m17/m9LSKy5mNyVp5UfNsiQ4HAmBkq9QNDr0RFu
Ep44lA9ODn5U2SrRXtYshTvaFCAytko1wZ3WgbTwrbPvIXB4Z827nWPpcs2uomGe/+sQqQi1mDQ2
nF2dILWvYBkcaf+HFaSW7jM/cuySsLSW41we4/2BK5u7ZABGt5lvroh5jfwby8Hk7W2TpHRaYMbM
z4qRGHgkbebqMPzEHgZg85PyTHKpdv/sRysJd4V2OgovTY5bsIq0z2AFKK2+ho02XtmJhFFLFq7V
KG5zanwQc3SSq49ihGUF1zFiqK7EohW+ccgCNA5WZOhLenWPo3qgSQ5B6q74Hmrkm8jXz7AxRKOM
XvSSjvYOWhric7DbHsaAJh5zT0OfYWS8LALNVjTxrtWrAUFOA04U3aBHRUBS1wzr2cYF5HyJP682
BElKefmKOC+GJeE2QhPHM5QdTuvRYgMkGFzsZ846IZJZs3NNgLRjmOhLeTVJo1QVSgmDbfUGiBlj
TN0N8GSIvCttUAyQ5GjG+8iaOfxdlFtRkRpLDV7gW3f0U4OZh77IXGpcVCGqdjR8sR21bZZizeL5
MNPYF9BWU8me2vDsrFyNMoRlb0AL9THTWjQvX7ZH3fzxyKVwtv5gOQlHljoRnBFFWy+sMmU4+y4w
udkbAnyIlRTJCDr0vJWfcsxqc7qz9/kuPJeuInboEn+IoUHRObdvwi0jzhDo4r4bgBQFyS2BNeDW
58H/QyYpLBlgJSTBykon8Vfo1dIyGNZl59WbmDe1V5+zAz3N7fcxjJl+Xv2man7yie8lsiEpuB6U
7NNaHwq/wbAz+qWb0Tq8dOAbe61yHQN9SunSX3mungzd3eBLVeUMd1Nsk5Eyq9R2e4SHkN3v9ARu
RNEcsNP7zT0cJXl+vL9XE5kuwzG9+F0XdU8RcJk47eEaruEr1XTRaH+NpmXv+8yjUdk0hJEsQIYe
GOi5weFR6hUt8XQH32ffBkfE4nQ7Bk2l4h7GPZr0bXiLdpeIFC17FkTN6xYp/p51GQVz9aFY73Eo
tTsBJrqPfqJ4CPuqamf4WlJ/yOcJLFM2d7VTLqhX9VeztkkKQD9tzW+zBy9qDeipXqX8YG9IUUgQ
kpnYN7SHrTe5ubF+bwZLIGwn+pwhuG/Ix4S9ZPDdYWi8N2k1WNMbnlYIkdMtd6jyLIJ9PUwt+F1Z
a1mhtWYATlKPLoNYdJozty5GlOe1vJyex+HFkE6LVxOAzgd1Nwcvje01nvijUevDk8W8HKy7+SCu
zX8cGNnkCL01kGhBMHoEdbFY07FmDLIs7fGZgIbxf2w504qbrnpboNj9ibDHyVXZwzR7ENQdbF3D
rq5zEXq8iAFncyKw0XgT84ROLiQg5zlVX2uqc/+DpO+JrKU0BVE52QVrCyEyPqWSnzGSaWSwlip+
evV6VpZFVOfetWpIM7p+Dc7fJp5gjpikXzx3iiJZ/P1PRzKsEYk06Z3bH9lDKiXx4icnv95IRtmj
Aorqv0znmQ2vJ5GcVwJwXQ7BYOd2ET603FclqmkW0uRtegypn7JLV+3CKq9aBNUZUm5UQrwL8smz
HouxXbrSy7sX8/3JYdoPsJW5Jg0Tbr7t5UjTzStrybjRiAikBzxVH/hbLfH5Z57okoWsNEK9mewc
Zizw8E1fl8SUn7vn9MeDhLefOT4siJ+ul+W5ybM5E817yItiJH7bHYmNdYBNpKNA7xw45X3ISJnR
Pyk6CM2fxnX+dK0tQJNZ8lUmJ/n5TuaVdPMeUAJPqi9a5vKgoUuFewYmP7s+/nbuFS21dIhWStj5
OzoVpiMOjz5loauyqY4Imnam3n1R7Rx7JecyeB1mavKLInpC2+eiy82v1D4LaDRx/fXb0Ht8I3cn
IVGNR8EbdM2heDqRHHm76hJvo+DJu77ulxRpFRBcrRPAjdEMhguByHPLxBfwULmxIrx0dz+ngBdR
FHTB0Z8jOjGlxzq6i+kvaYRmJr/rf3/Vn60AMPAhZs8eu3eXLJBmO2w0BbZwZZ8ZEMjr2K5bheFs
mJGDpCyEXVmEb7JCbEK2Xgtf2tpawrJHZm7N8acpy4ly1+mqoqiJNH3SpC5idLLJWIk2Q2YuAJPB
H1QABfpbd5pUxTL3bA1O+LA0nOBfyWvxGHKVzT6lKzq/dqe5Hj0KSI74XwMshSKg0orhrEE+Yk4z
NqETetCZM7UahiWVGZKhKTe2GT1mIYELIxK0oWgSg6P+zerLGBQD/Spp3D0eASwP64iniktgRL6E
cnlCtT+y9aVMGmUc6ZxyOSO9qR6XwCPftlvGICE/aKu9W9ah1a44aKwGn0nJbumno3x84hnTYDnW
pOv7MbyYTwuTwLl8jEsrKSSNefmqt1hoynAkhShuQdSHowI4JEWDfIs5+dICajKqs6085DDqK0EC
U7MTgViFL8jEDsZG6iF7G5Duu9uMRxjxoZYRhcrH0nQKEQ/sa2lR/h/nD/qlZw+igs8Lr2fE6CDv
PTv9VQpnNoZBFMyTBf+aN8rAf+pwmjiCg5lOYQ5XVD02vn8854VBu7kY04j8hxyJHSYumlW1ofgd
PQ3fr9jhLyYJ3iZoxtyP2iTJdNj6ioyTusk/8iz4jzQ1DBrgvcWT/0ckGRs70AsHG3ItQNi2yXR7
NjX/rWnYB7aaZXSTlVUYrJCp3GSL6n0tu3xX29a1ivPpLjYvD8LuF38PkYE5qlUjBiMySAqmLQ8I
FKUZukMKAFFm4gKAmts8y5Dv/Ls/uChSUOMJ9PrSxgj2SFTWoP5lq85ic8cJA77sW3MqURoBqlT5
94EByvvjtnXg+/dzM1xQaE5+kXwHeLFhi/V30tAmLqCN7jd6T1dOwFdq3eUKQHsuZOgxzrvEEEgV
cDDstCcCGE9EezymD/rFETcOzprDs2jygjeuGof+kmjtA3sYOpMm2RN82XalOea7+u5senP+ei63
65NrF6XUx6CXRODgRTDNnMTlEbPlkstng/9NA0OStepIKDbjoL0vsGAwPJuwGMYabum3+xwScUI8
SSTBOoiyM07xe8nFtGsVv3ePB5LBDpUZMpZzOtLdkBAT9qOLxzyyhRZ1+I0lbvXdA6S03D2S5lhw
4gaMTf8sFIiUq68mrU/ofAOCkpGCvVcEuN3Z01N3IkhV0iVVrITqP5d5G53BdbxS9dyhyZBJgGIy
+biYiTymjHrNhJhIR92ZI9Bt+tjCGUULwpxPvbrow8/qB1bkB2BMpGGjEzqjQZKMYBdDi8Kj0kHx
Jgyb8TXpWsRuCkrRIXDo07oBIu3O8+Bqz3JQXkU5v7IvGpo3H7CQXSUeXES8PuWkUuLZZbR7zcan
qcP53kZDt5D1doQJF6vMsEXndb7LOpNR/Fp5zljH+Top6NbCSgtetWN6AbWXgxCDqVqOV52qxbJz
EkzJaWelySJZlGZHj4jzjdAp6tkdx6fKwNbYThViUkInwmyezJxWVi6snUxPOcT8uA7gtlowZJR6
yphaOCNYcMy0ayZjcl3xcZSW4bDonvnZkNOg2OSfP28q6NJ0/T+uINLg3kssIdBkXRZeglZuZxvI
N/rqBGaZj1K2Z07fYz/yltNg9hSFzy17QAkD0zTquBjN/7Wi4EI1JfKe8/ervadKXwa6kMpLdnZO
rWMZumIxP4DRtA5fZIrLFLvCis+isVGfkx9CNSqLOhiBzblrIHPdjcEAu3wAgApXUPexeeVIane0
BZP3nNZ0t4S8X20zzbNRkGBJ/rgxp5XBWe7X3TiSp4dhLOqcC1+QB+dAr+0slsg82DpNmGqSQYt/
491wxK9HxmAMM1J+bms+fwz+D8Ws0cwuKCplnMTNT9iViYKvB2HPqywPyMPl9R0qGDF8sqdHrbyv
O1nXVyPrH85XVIoSOX1h3YPVbPT+FQIOpLW6SjpQ7W4o/zT9mytDx24dXC05ux+knekz+8GAJXH7
YQ7NMFHIZWV+8gAsqNKOijy8X5H+TCksJc6Qx7ipzRf6paJ/6bM0419BraPJBQM/gf+CiY/1/D/U
c5UPtnBIeeTPnT+KuHnh/DxSvkrEQCL6Y81YDK/YEKhjQMWOAoZgyLjlTTCUNvGh50qVf7cJdSRD
aO4DTSCrcADbRTrzY4TwYHHa80+VPVS+DHSAkDUwW2kTcILdyB7i8w6ZBTU/leBzS99SuiAeMBGv
5Of2aLKFfG24G1BaOaMEc2mUoqw6Gp1hpeBkyEhypaBJtGGX3xXvVDaTUswfVbs4gQmiI5kWfF5x
LbI7gXv0BPVkEuc36/9YFdMNGdLRH4EXepQXufzQgfGrJXTv0PC0csIN53wiAVE8NaKclXX7doGF
ESQxqlBCsBMq5EduAWcbvlXd44Sgzt5UZwjE3Mp/8OgjD9n6z6Ba0zLsaN1Tdq8caCSgN+8FuXMr
B9ey9IcYJvRETsejytGn+5V82aWk6MZ/NLhmrUKRgvxqGEuT990qSeQdm+Hg2rox6fqxhfIThDuM
HtGO7tjpLZ0lNUAhOJ4s1TBaTl9ig59aGx0YjUOz0M4vyhEuwlUlAlg6SG7WZRFPEmaaic5yiR+F
JxH+w+BefT1XVvmyqb+OL6hDnZfB/XBH7EBRTQa/+RRjcpqkJNni4SHUIppUGPT15yO+2rnJc++c
oYQea592zYVhIuInwsYUU0ieiHBlGQz1Jwi7mEze+MePHvN139gneJl/D3K7eVWXQyvOu+lO+Wea
j7aunWnHIUX8ECNcbnqHVR1QZUDnOhnqMbj5A5avpXEzljT3qGx6QQEfJo7jkuUCL/6Ef57ipmC1
AlvUUuBhS1IQXUTBBMqt+B9B9JRCojGRtRmJYUQ56y17sFgcXJvDYHuCvntgZF6cFVF94tIFZr4N
Om8LusMbJcLL9ia319A8JFCOM8dX92BO3M2+gGcYtxV5agz2hKj5Hcs972IpBJbptNxdkp7a7jME
pXuKn0wETgYftNW7fwz5KLXiW1UvNxJ46kWT5UJJWkX2aErhs5RFOUsbEGrvekoTVfOMM15OZmU3
cxbu84+IBWaBdAhl8crG1lhl8NUze4g8AP9/YESjIBOYEQPAPRphXcla6bvwTHKTE06FryQftFF0
6qQymAzf/MYPRC7Wa/cTdmgZw/QnrAGOYNSMGg2iSh4omp/8fcBDkKu7haJOlKcIbsprD07QG90i
4YkdBPWs2xYduSHxGaxFCfSCPXAEYe/IpoChLuPqkjV4xEZCnd1wDVg6yAbBTZKN/MVivJEvMj8q
Rsea83jZfyY3AJro1sRThXVOK8A6ncF7LZp3v0Wyjnfhc3dp+eLd6/bs7mmfwzlOi3bxQq7f9F5A
msUuFdkaheywt/qBaeB80aBcirqKCItoDXXL6Pq+tR/H/CakWSWaC++Yg9GiPm+f+xd4+Zt/Qmj7
GfHgHfydKGIznAfxJBFOktXAWJm4RRPXL2R3zms3atCEuC2cBQXuwAsx7dY3jn9e+22KXOFI3oNy
IfJf8BdvYb+awz9NUHeIzezHDj0903VwEemLh4rbdQVf2S2P2LPWKEm9bYxB0IiIg3eTtkPl2JaB
7R9klTXnuDIlXZBPcHXq2s54deTkB+pxuK3atbQko5q+Dpx+xQXrQ4WGUS35hUTqyDABX9m9v2pM
Dap77B9Khv3ezWEi1yCiFSCHhX2nTiaj0U2mtg2DOixlTBBduFBKDgxoGGx+TaveiH4WwHMTm/mF
fuMnaVSr+LU1FNBwmkBJ7liJ4zT2HokSgWtPi4WTkJ36Lss7IFxh4DSpKFu9chLFVKDMpB1MHT5K
qTEaojMZDJZdv8CMbfAuCUbNAQ9UmexbvHkEIv10ef3mq+4Brxk47IKQxj8oG6o6+s1U5iZzSXZx
8mhYsRsHsm6e9IAxUMYFNYEenLdij9tlExvAsRmKpEsTlAaNZLv/8CPUkCZPLewDE2tEoVHDicZf
MWYXex6czvXUO/WgLeCtOOq+NRIh7v3sHcMWPH4kkmkImxFL5hGdHiLf97Vywm8FgGLbYFOfUFwc
jW+I5Khh9ghg5tjy6cS8dOO2ubmQCUnIuB8/NM8j/JxLE85O8tdOM5/x4XiIltgbHbCFI0ujztOt
tVjs6pCdNk8WIN51Xi5rcZvL92muyk3NRFNVDd5iPHCsSEovNYdJxcawPzE3QEt4yGo36cYC1qiW
FxD4HLHWMRe2m8UFlPlfx+w5uO/6t/+YEeFQ03FC89IzrhEeJUmLPulGIH0mpMSXJ0tkiIPhnV4o
rFXH4HMKA3HJ8fri5NlQXdkJpcDh13JueTx5dte9s+pp+dfz1arVp6Q+wpfvqFjScnXXeRkcuEjQ
UDuSZD/bUYMIpPbhd88A8dAclJjtoA2LxRT+M7iEU7N4vqz+0y01bI8ED+oEgSP4xrr0AKKQH70i
wOL6YxBgWR4vjZ2LA3a+I7NhJl+UjuCtG8knjGDbgudRWGtjOz0zcBza5TAXpSzkQ/PlV84HhILj
DdOAIdNGuUq1ZV5XnhkOk/swOmgNYZKVXAm2YFxXIOEriefBly6I6GldiK7jRD/g/BiPYTgmcDKv
j5KtSpJkIzI6RVrGCd4h25xriVkRJgf3Ye1wi7beo3nON1V3no9KUY+2qjKeqT39Xgj0Mn9AQO5C
EEiAY0n8kc0B5q5gxaXKNdH/JMe8A4Ow1XmbQ751OpWjBNJmdOP++Yxxyn2oozCIAsrgMDI+kZmU
gmd1Qb37URvQXwnnQWSABoAjCIaq34HWrDjFrzgTaME3PTyG1e4A1zTDla2kBRsOc1XgLhAU5LPZ
q/V5N7rL8KWM3G9XP1bWWC/CRK0rclBSHJnCLz1iCwjFes3R8gaIAQWZ392jJ4udOk2mvs8LE0Qv
j3/5DaQVZONbJSgk8lpwd4lUSuiOQf6hlQJuClKo4a0K8pzl5isI75vCOpgdc2M7q1IDpU/KFKzN
E9hVKerIPD6AOjbKnJTIhjev2iTDfXY6cVLxBkzWcOkmPTk3fDupVk9Cf/iQCSeEMvCvksIKSKQC
iDYn377oAjPcxMkr4qiIUl5HltfoO1UaF2BluuGwDLt31La98cDVfo87W9i3xG6I9r9qlTm7UBVT
qBXBd4f+afm/ukH22RoxdwxILzsArjqja4c5KIJ0M9sgEXb729h7NYyegx73/wOaAHZkdBl1WwRL
YkQyQ3xGzdOdArMHrX63F3gLBEwTarRmabGuhdc8HXmln2gh+WOUuwQbRt3pAc/DcnuWAsR263zW
KZjX5bJ++nkEFgyhcMplPJd/GK0Utaa6liaqIIp1KwDklL88CseZ7TLw9Ufzbpk7shc1hGyddOIj
1lnSY/mJLfK5xoFHp15pPnV0YHUuGRHyLuQXrvoPCCcByooEzra1aFbWuqzIBzwvTufbtE5R/pR/
+BQB4AK51AfWlSnH6VzTS6BIFcjPDrvu0AxqR3ORrym5dOijhTyDFkEAY3TE4BDsc/3EtLgMEmNs
8oV1Z8WEYTSGIlA8yw0MjmBu4VCqhnLXE+r0GRyyAO4v/8XXR7OWGOSUlLAL+pc3kM8hg2P3vsOE
7N1u5cntop9Hvey3nubKgJnAuZbY8Q8V2sjDIQnD52AohEtOS2GdXyQWsc42sGr1WLXonc19Tda9
Y9yqB+gnhg8UCsUpN3LYC3cSvzeIDm9tr7ewhxKy/ryrYthY89UgEYQHfLfHQO8P60ogejgd9xjA
7xknYFBbeT5YNRb2GwF8PrFV8jrbsyXZvApaanWArtvcy4LB7rdbvJa5AWcGacfXbVcjhL2Pl+W0
ZQDVvo9bjJTKn8uuSjh6S+RH3ZVed/abNbdlisCvw0gOCPY2b390e4UZCoHNJdt0fvMjd5vITsR0
c3SNaqXAIUzo4qmi+dXObxsm5GJoLCdSL7jKX/CC/VFgS1a0OLIsX7zUd01r+3fWZ98Z1tzCEKs1
fLf1kr8AVW+86as2RKPF1zmawdpCFt2QCE2iHRDmwPpgSr9TFIwAtuNhlf3zH0C9XLdmEztGDGzN
bSmTe/LfAsDW6IKS2vGzaupVl2cTHvuerbDMcnwvnirjzPOR3fRkJNxElX3z9r8zp5PqVczprYSE
qCbpeQBSwZ6YhdreLqQmvZKgayFw+EoOUqR+ecHGbuLj+n4ihICxc0a+fxByoPa3kbK6eBw7Vm7e
5JNjDlDdm5bKmL+8pcJoGhB1aPJd3wdh3eu+x1NopOhqDYnd4ClsXwe8afWelahipnbVTlfvtsh+
rcjyiI9INg8zBMy6xB6YR5QESWeBXfssVQ4n9ejJLUPyE3GaYHaCx9UZHiMWjUvZamOzGY9+5XUT
wk8M/Yqh7IjbpVHfIPZjxqz5ic2rs2oc4+WqXJyVcHAV+VGhiI434wr486ZuJ5kG/YUJBXfl9jii
QOmLIotOl7qBN7Ndgz4/nEYCMRYbtpXcrm/3t/oV1Fb8WBYwvG87NOhkgAwhYiggq298OqkBlkK9
f6AskQRZFLjJdJK1pjqHLdL9vEitRLN4Yl5Zl0JebNM/PaeJE6GA+Z3XkEmXfrsfL8YEocawqKIF
1jioDbNMoJPUTwPJvJYrpjeFgu0y3OQhxYHX7ZweEaRbzDbXA6USI3RtcgAzJ3wKEhgmX44brm2x
l7Iqiaw2BIkmzOcCEMur07kuy/5lVg4jOvirE6BDznJKjeAbpo2YWwET41bBgoUI41wKAmvRGsrU
6/KW41dPONFhIMplxE6riKjfA/LG6xWCOdGBt5lilCMnuudIAZdSh+YEDdBENKuzQ/ueKDCOKFyJ
0x/zUcJf1sWxZranrkQdf5a6OFhsn1Y4TrPj3zWAHRjj8Gg7B3ZQzWC9viw5TkLn3g819fvNf1s4
JDSANQ63X93aOrR6DeRHLnwvqG1JDofNq1PfI6i6L/yD7/XfjLEASWEv/gfenI8gg99mgCXK7XoV
ACRnn2vgGjiIC4S1muvb5i4643ZtueK4ZE7Mqkw+XL4lWIOYrNbG833uwMqAxizJE7hDcReAlXVm
AwX7FSeaHbGYnkgQiwthi74ZDCFfXbopryF1pZKCQILL55p6eGqHaJT0muYM5V6UMVRHeGRjcvNO
tt/yKAb6z9WIi9Bq1OvBgs8eDXPeL2RWPw3HQOx1YuIE2SduwD0J3c36+hPUEdV/H3R9bz0quFR0
xVCF2MvCjywYdO0eotlDsHdrEeFF0VlLmXvcFAXyACm4CatKlTUfOgH8NiuG0apLOBm4PttuHvSy
MXfiaPTE2URRVHAaI5XnV33L2fRvbrluIaLC0tYfqgefmwerDPEuc5KT487LPLkPHAE/hq7ZgaW1
5ZjjXo7SyCUZ7DwKDUCy2ps9FGXFxWtAAauwZFyig1jFlBJdMIWgFnoh+f+VMlk5ow+RRfBuH7Nt
rgOFsJmHTKK7/ulIwDoaq2n84yKmaJ3shBgLnMSY+sBTeQZT/r5UoZRyPPmYKU2TVzTgZ2IUhHAh
O+qZm1OjNsDufS2IcQVFtIVMdIXMxtcusq/H4vfUzCY+3jiI+MKfaH+FhrczA2ZulH8ndK+h3t5u
2AxhOmCvp0HRonJu1lAp73+AGmvqD0SD3h30tC8qYBN1VBMXqDgUvIQOHuqYeRIL9X+5TTXI0np2
fQwcYct2NCpXof94GrXcXBaV92g4ah3u9pDJJldEc7pcByg7RzNi5AeMVNgokF3D4IXXbWSPSPzB
rCIGGa1Q24EcxJKDJzmMdt7wf7zmBt0H2HLEAen4dpWYQTvOl2tO+Nt4cjp4Ex7B1X1bWlZwV9wr
7oQA2uM1egs/XuqUvD3k4GGeQ8vcpJoqEJsBzRgNlg7F4tUtgRd2rOCvdnuHZnw9KpOcom6WNy6y
iSz+OA0m+InGqNbJMPjPQzpbFPr/8fENvfltAftiIN/8G6s2SFMl2pzPvq3dLSZCFnQ5DsiXY3/S
k+i+DZDrJaLeh+yBTSmnwKd8Km1/5i3+zpBWGPrcWV3jOMIrSb3b7hPIZoPSBeF2N/kRik5oCGXp
JKjBfsEhF7mcI9pltZvRkAywPg2nQTSDg6Fd9yie7K5UipHSGS4pkNe4iZNmgwmiAOtLrbu/cJKo
4qnoordZc3QriSxZedBeT4auWwS0L1XeuJM8p9GX6KUH5r+iqlyqkRsT841q2j+gtibzx/VEyN9y
L5GyibpkjqkHIPPsy1Tg8g6U0pEuGdZi/1/mX6RGZXJImSDkt/vIT12TvTfJveIdk5HnIxnaoH/C
bDgROGF7lHDyZM60/1oJ0lvg8+PK0sK+ytHbwERDiLKHWYjfHW3kgmJ/8ovcpbUJh47K9ZHaozca
sR+coGsd+GrduJnaDdagRBgXsltxPlLJll5X4dcBawH+7sTFwd0mcpUnd++4cN/fFRA/MIknyvdK
3i1iVBesdyfAh/iaygbeMDH1pLEN57oilPoIjUkq0VyLZiQUQRKyzhD4KhGp3q3xW35hXS2dngde
pDPnWAydd0tJnUayIqCWaoGuOwBWptnjKfEs2SiHCpT5It95h15SBGDM7iRd/fk/+ge3j6pO+I8W
hVRaVKeHwjvE4wlEdcalLw/ncJzMMu1z4WjIHeuqomHoGURaf7LGmcWP2eDQ3rKU85J1yfPV6S9h
5LlMZrxys/b4h+fDT2No80kM7OX9CXWtouXqv/N2UUNvKhi9/xda1YBjEmYWMFCaPF6h52R6MJ6d
ZdVgoU0SnH6IbD61amsj95fmNtWnMsBatmYScLSqI4diaUDLOr9Jeg+ubaQUOSDi9+mZE+FlRF6p
3bZ6YBPIadKbElhsCaj9xuIUTaPkObLHg8hJkGdYsxxjTVc55p9NkWwLJuKyZs0KigtrcIGBd4nP
sxX5bT7A0iBjoU9SU4IWe2jQAX+YF2h9Brb7DHnsB8UAJR0rnifYp81HxQNwiUb4rLxRdgWuOGz/
6gpHxLII1Wx2WTGxgayKe2Jr7SulCJudqB7ctiolk/NvTF8ZWbIami8f2hunVmBpEzfYGDTM4mED
RM7UBLFCPGUU4Tbt/LixiG3Bhim90OW0IsGrBe6SgVWU+FJUYxg3GYw/w/7j4RHHUp/rilZ1jVO5
2rtqq7lygpqPY9XvO7AByDF1GcQaCXK/TLgKageRBoNOn/amxxbNqF/lfi6FJ2Mkcra+Sst+NMdc
tTTTEmXdfQghsihc9OYI39UzUMVEZ4+ji34uylGIB/gwUdyT4GvgMPMxnKamR8sBtEnfn7Bniu/L
onZ3qcr1iVJvQVYGmfZYACW5B04v283Z4hoYns9Eq+Or7Gr4H06YaOpZqTr4STwBoTz4/fRwx4l9
Sb44kcFKSywtGo645oX6FxVJfclEaFw1kJgBdlkER5JDMEfRXOvkiAgOHKUtqaf7OobLJhgWhCbL
5rkkitNDpkXZH13zxi31zaA3jSRoAmHzRut5Krrndpmk8GYN2wXmHT5yaLD//PYOpzPH3mvUJSYY
596J4sZyU/KHJXVLis1G1FlKtkrhpRv9kv5M+Z3U4kYZsq/PGKMzuTsNQzcSqJjBBOjt3r4tZiev
FDwWVrsu6OA5lhZVNcstMpruGwr1xR/Gz7puHz4Y+m6Ph9LajhUsjB43f4qJBvgiOky0GozsUsUm
edsiyywCkYFJwCopPf+rzjK+iQPfZgInU8nyDJVf+oEiqR3fNds0qVhBenQmyH3vOxCl85yZUhIT
zVRdbPhTtjdysvFLUyETUNq5nVQNeWvFbotkXzEAK5j9ArBxAmB80hkYm6wfsE86ZE75L9J8OK5a
Df0wKNzPjmndZPXDUQi3CNQQtL4firu9chdG4cU6Zfm9ItWm4gz9V2YvbCi8xnrN9mIbn0sMYcgn
YWsEUTFhfXQQyAThRjfE2ig4CFu/XDqRLrYXhiQyKbSS1PkWPquXRjDWwrqzNMy81ly6TFfhUx8b
lPrOGV3ypChXCjO8mJyUJWzjs/GfmES75nG1jYLgKwDux767AFjIPnr2YVinsJgMEl0nSsCXKySD
V2U4YtEOyGRoQuzXtsaKnt2AFaOWRTR0g33TOJz6MNFRA1k5Jdi3gQXNL3KBOE/k5GXaCj1D1kS1
j1IbRmcbZdV1X2FZ6XatQpSmy8IVBqy6kNlG3tz+3raLtYJDQAx9067nSva+y23TrTuOxJ/sn6i6
uLeWu1pM3a4vb7yGzycVKkdFCFATmlNcmfQ9SwO7gvROakU61tEwBrZOIWNDSOt237IrATAxmPp7
xqsNyh78S17GH52br+6tEf6UIj+jfk0AQAsPHZ00oTLd1PLo7zuG5dt9JTSlahn+dTn2M7AMqfqk
D8pdv4/Ftib8/L/nXSvYOxvf8dY//rG4b7Y5b4lcvQAeLgndFmjM+V5hJkVZhklMl4HdlQvdeTB8
72OxsEwXhJBDNZQ1ZqwiDXHiJL3U+ZXzlEkKrg+j7//ufiUfGUpH/+4h4JY/naaUc8twU2IDTuuT
fy94oYv62XBwXPsnQ4z1dHyrVqGHTo6WVwk6U0QG+tGcGoSiCkeQQxdvm5e4JDr8ksWNIW2jtCum
Q75ZSIWee82NFiGRv5pa3KX6+PN3mJK6TTeSWnlqGH2TjHRT0diS4mWSyGyNSK79dt1LK9L2ZeSb
/B9Q3jMKgpwNCjXVIRiwfepUPSCu5t7VORfhrIxfdLGkxEsQuE7z+JBGpYuz6WUg6nnK27Q1PRp6
wOFkWcXXvOayp1aS3+z6zZBgF/Bk0B3MxAB14E8gj1X6LC6XzuwqwnHy+c1HCVW2JxOAwbrAOL9K
tTrgyjrVatyhNm2zkoC7FwkqCkjtxYXigPUi20vD1+nY8xrtS+r6CswWR019eBrudcIToSkHwD4J
4JitcIO4jHOya2p4/Br7iyq5B5MaZD8td610hkXwWxa98/2vOnIbau30yrc2dxvPl8qFijwWHhEj
EHKGYbEOVjFXh2uJUpM4I1YXY2rnGO+mPAQ1zw3gxi1lzyVl4KUY6NFkfru653QTQDEJ7ABHO0bJ
XuDTfSksbGOG8JOxlQnrY1Za/HZq/+MIBz5NrTtV4+vGWse0PxkOknEfOq1JXPY70hWPFNYWfwAE
PsFCuJXHiNZXITYNMkkgZkSeg/eHt9KmoOc2KkSOjPIXv6s0NpgSFzO0cIgixVqyjlE/+LqUMMTp
Qrn/dDTHeCzwtXiqETvjdv6KNoLV1kMBp7xGGC/0dwPVAx2wADPU7zJp4ef/sEuS8gkgc6PDLO+D
kWWaZj67uPitb857GLVS1wm+jixziFjqzaPZoGpS0+j8En9kAQKp8EO16PDzXNd6NV8/PdJouxJ3
0hmry58NoNWPXHrLy2gfORaZzFbyNJzMTVshcUutiUf/a6WgTGYJMiFVhL0qo8bG3OJPRC20z87N
fFirmQjhHjUWiRGBrMblVRAjHSfBe46EAIahphKoVv3aTI07LofLqv72YaVbo3MHAB5VopJmSGMT
4oykI09nrM11ZAlpYxnJ7TfHnyHjPodKBbudlwXzVfhyKnDC3MlNEYxBDC7kSGN/Nk45/5oD10vw
OTVpGDtPyAh1FeKoun2pzU9sXpbUw4SrP9sfHYv2MwKOKREbesJ6ROCyi1Nrc9dWnDmjcA3yaNIr
E0kKXs8n7NU08xxpbJAZPpc+lvr4M5ZNlBcMg1qNhLQx59d8Ph0u+ZR3CI4MkAWFYP8kWKV4oiv/
eUl/8GR5U9I47ae1vGG1Qfm84rmzqHAzgflL5W8A++GmZ90p6BPg44hFSZNg8a/V39PFAOpaLeEa
9YyEto1jl8cOE8QofLRUUdmQ8GiPglP2PDIez/ed10mFMGhWV+adFN9PdPxopqGxkzFK8TvjV25L
kLxHG0ply5Ui91drHgP9Cl/J2tuK9VetmcTpXgidfY4NtFQcm3xlO1rzV3GilaPz53x7Inc9EcQ2
FwrkdVyPWo/xGxvyeB6z0Xakn+rwRkIzvdaeW3lgKEFsB1nE9OG+StdLM/CLCcJbxPUVpLoNjZA0
MV7ICrmT0+kNoABpleA2JsRVRc4FsguT2UNznyYcxJ2NCN3cl2TSYr5Lli4S9pojR7vi2KIxqrDd
hNXGBVtyb8iFOkx1JYz4C6mW2EmC2UJGt7pMnH6jW2DjehA08qHx16vLJ0rKja5tspHK/XNhx9N6
32hW75dU6Zz88Hq3GldOjharmGMu+xAVFy8NjkGR2xopU4gBvW49UXeREkmLfWhfh2zndE+JDzOH
pRDUEIJqFUb/WBnA6Qm1GeN81ZwVAMAPhVAcsAtA8c3hjI3NtBxVdiE3n52kUSLXH+mNQ3Q02lnV
mSE3KMhBL2jpOvz1sLlmG7xO2qUS33SWMax17si4+hPB5V34MoL2qR3J+EqrgG+shjcSdLaLBhTn
JQSYWx246FGcwBvRbtv1z2WTIkRaOQBYfQuN46WCo+9ouo6Mm0Z/1lcNEdQ16ZhHFHL7InS6w3/y
XPCCy0RvNW53/Yvkr4TV1SIjkAdrNNw5aoY1KDJaqfC7FBeEQH6YiDCxL2TnzmVxnjvOY/7lvy8R
CGyh6BXEQL5ADSsAFa1ivv34JPCMMBPc+jftBYBvEAAD6F/v45CLbIKF31ENEOqdZ2d/mO9MD7y/
XFe1x2TkjnBnJKgH5xwIqTJ2hayipusoOgSwBqzLAQyIoeOgQ7GoVEEvzF0RuaqfjjtlveZJh0/A
V2F7lyk3RR3O0VGrR+AZkKYIS9EbAT/W3M+UC3noQJ/Txs3J8DAVlysSaangWUWVv9gM1HMMu+Dz
3qH2fsbpYdaziM6kC0kE1+osPzFn78pJHM/WzrAQrsB8OeZKdYHxSTwP0MVD36Ew9mRHP7Z6uV39
FjgFN9JFsEhj9e6uj9gxNFUvlMRMAMxkEs+w7cBF1fAFI4VWv0HU1yLzm0zCAE7xLcJEz6xX1PGE
QZRvu8BjejMOsgPO7olQzD480ZJaAA0V2/U8m6M3nxBZ1SoIYn5v9VwFGWj4zQnYAL5o7wBpyOgx
mareJqLbB/iOem4HmKbzjf2zg9up1fVe4JF//Au+McM81l1foJOTpoOCVo3n+Q/t15VSOtul/FSf
QtGOxJwbbBcwo8T0gS01oeBAXJGRYWYMB1OIjLXUBZEMEjddbzjLFAmj5o3oYSAFK0kb3M8tURjn
49Z3T0GL205nir0B5gCXb+ZQdgfru5H9wtKuRGDp0CFUgzeZi3/LAZmWJndawEZ3ljzMnQJJBL7l
ljbWInHucn8PDQEjIN+rhpIS53BRSsiCUjq4lnQhE03w4N+pMUsXw7S/mRaMqHokygih3Qp8KoLx
A/eghiavpMcl7AiZ2sw3bV5WkteiFgH1ioBNQLWxjf83xpGVo3LW5Kru5SY/9ApGJ4udUqBP9c+7
ZleVqTuNVnghY30VTa5MywEBrjh0YDz4NgC+3cmtprTViE7mtHOf2fRwUmhlPL3kHrVoPFbe6nDE
KmCinAjUkyOqyE2GmXPjUJ/9Yqx8679PM+qDGCcr8X2cNc3/GhunQwJQgCGG+4v2accrF/uiKNjF
93BliGD29+n9r3Jf4qXl3j6Y87TvDaBzQTOMYiGe8lSPeFBQSfV7KLKcHXKi+ice6PFXo6IsQZTT
EoT6t8vv631Iu6c0fzPpz9w04EmcocXEh19C5Xluef9EvkWJgpu7ZK/P2pEBxfrg6maxjsfA92Q+
6GR4KbW2p0/3c8ajuqU3cqtsQZPD9ZRwa1bXJ6+xCKMamaWzkWVJ49SfQD2C405+pBrfbrZNZLOx
mig8gNsoBI49Q7l5HTrlY5eZJLSMUlwR9DeD2PtAU7q/nAarJdmckiwHHsGC3GW/JToBdChnQnTi
Jc/ja9D3UU6rss26i9414caZwOI7rF8HZOxyJ4E0Xquf+LBM4JnMhKdUcMQvbr2kn4pSZx4R+HSA
AlFs4jHvptFwtqrOdBGWR6FeLhYyb0nnrczMeDLiVFGcnjODXjZUv4MO6NO+dqZbOJLku6zkDEK3
mP0X7WtaEGvIuiBmbuE8jURARBRV7lwmPLyW7JXQNqdWFL6d+CNOX7Gp5VBekXiCmzTpvENm82qS
mKckXVfj+Ewnst+FGqGulg0hODZM0PhY3BEKXhc8MNJ8kFHepYcer51+sQHkvwDWh0tIhaXoBRq/
iCi4Lqq2MAmaPNFnAs6Ju9Ry3enti3NcJTpKKDVU4OY6LnVYyKHLuNcSVkAy6IUerxFjc6iKSrZ5
X5ADMTtvy16ueuwIgiAFai0QRy7PMB4qt9q2onnxbjgmFT7uiLUEIKlhXKhfQsx3F9AQpCzWFzMi
ia3XUYHAu/tdTXAQ3aAjmlQKuqVUC5SJPF8UOZ3dldb3GdgmW119HoLaFuvWc9x264AqlddFmXkh
2pNY2RT+NzORJuSxK+BDLOpETfDtCDcOhTY863Y2GgwqMVLIpx5BppsoqeKQITvOuVbLzD8RSVYL
lToreC28+bGDE2NNDWh+N08RKjLFlFhSucyfS5nJxWoE29jVOtbUv+gF6xWI+IyN+nJ2BPObdMYd
fRbs5b5+DmLeE/DN6VRjmVCIuOIQMcWlGZ+R6ZtxHUYM+mJMYZYd8aKRWT/t9XkMRjZJEV90aspJ
LtX3MzvSm88fXag1OFImH6/zNRZqW4xwzq/BeQBMNCRGYmoimvNs0OH3EV0ANGgEhOM5OpVPwn8=
`protect end_protected

