

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
BwHHaRYHij9TGTVh7NqyF6fPKvSJbz6zXpDQ9T0CSRjM0Tr3I2/EoB+qBgzPRFij4R1VpNLIhF/W
jnZk7ILw5g==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
EoffIvgX5Yh3KSkMHr6Fb+Y16CSwhqKyrZiel9vaFNUa3EtfX9ml680qKyH6k7Lt+GT7JeOZ8tsv
GeWg3Is5mnBMAsR5XkmKmU1Mf0hiU70CtdaVxbMu+l0K5NkyBzps5GWZFbpBi81xyWc3mZBrsdOP
SKFV3jiPDhzIXFusLNI=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
pC+fmAQpqkr0vqse1A8SFfJnAErWB2cTBoy5W2fu+Qfel2Cgg+f01SLqdiCqUwM3sdVOYKq280lw
0KlccFWeISj6EGy+UhrlckR4KPE0XJ2GFpTDwr6dIxS9OpYPDM1MXlxttLYJRqT3qA2yEzsidST6
0i31grVO6qNsjmpW2d7uByo9M65VEOheITjyvjEpcaFShH/Xo714T1rUj9u+HOahJ+Y/IZt5BXf5
ifgOOsFSC4Urhn+vw7WBdTykWaXAuPqSgZ+BAzkf1tn2a5qwxdC/nJyffVluJZjwqKsS2qOqxdcW
lV8I6VmHkVrsFF7Im+SIdtLtq6ajfsK+Fu41Qg==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
sjA1wOpImDpYBBRjnwY37zkJTSoQvS3OSqKSHwre5fBAKnkrgUJxozoTE8i2Z5d9g73A+Dh1Khan
8gYd3xbR7Bt78jJM+PFuUbVx7c2wSRcHOAp2KIXVLTpuc4ycdBn19YJhb2UIFhm80kkNGNgavUsF
mOqFyOQQiDU6WY7JVI8=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Yt106ecWVBUI4xOZZkRHweGkZD2nlI1jRN4H6Fzc3EkfIh+DLe1c/sY05LO26DhXbTC0r7f3V5kn
SKvkly14VHuR+p2mt2PXxY2kZUcL6SEF75Sdud7O3qeyYyxwzbLXhAk8rv8ESHYXdpJzGlAIPVhc
CV3MBlzutogOhAPHHcbRbukDx/ONHomfzueq+JuKHmbmSP3Sji52yPtcq4iLW/WcLghIBdR8EZ6j
UoWFDA94p9C7hEbP1WkZCFdBxukr8LSVfTsZyILoNCYLGaM4SAN+KSvY/r6FcDftOrSTK0VkVrNX
POMgLw4WpJ2xpIx+qCPH347wGbfYnUgOpgfHdQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 39232)
`protect data_block
IF6pmlZ9ieqPNyfXXpMMd9K2zx8SmVUH4Om31Y0WmeAjnijdvyoRu2qMbG9J3jfuCm5/62ehngUW
RHYu/Fuj84lcL0iDbq84wpouAxfPRwje9dxdgVv4HvcVe5jVPHiumExj6vgUahGrnXTqyE9Qo0B3
AXGRULQh7hwg2PdaSambTYSeG6r5s4oYsA4J7EkCtQ/TfrfzJCy5sb70nlXnMOtnvVI5457gTGx+
8AhPUncQQrYHz9lmaG5pxx4XLRLb0vOFEDQeSm3yn509bJmlGtuW8yK43ZLidJ/3mW4gTJzBXhic
ppL1tShUZOHMr7s5t77B14wsQ9QKc0sHEiuFN7V27G332k8dlC7gcHAnGLND+R2k99NnRgOwW1kU
5psVnf2EyxL+Eyxzwm6XVClRkNX0164UmH5R07+pjoZ9UcZP+2XxzB3Sh80oeAiMk87FJBRUllIG
cyAjmMPOlT53ZwvOZOuBfWBreDdCo/G5iwE+ZQlBhtAj4I9ZcLcHumirU0I/S8cIspiTxku0V6Uu
YVAzKkBSt37u+Q70CwWyBetJ4a42kRTJuME6AcFtFR8GbSAvg5AoHlrKfBWgt3SKGeAZTLAIdG47
7rdbf2Lk8tsEKlRg6MTl5X2mEi5S96HycQ9v5foBW0yMDp8pP3Snbx3vekDnJewuWS83u5pgbVKv
oNzEzfO17K9P8BfJ84zD/hkeG1SjHdubcMm+B8EdwKWEKo4qHy0ByX7/z2ElAwql09v/OZXEqm2M
r/S/yPzYP3LTjor9Na/pPzsLkuWXA2wJGDvCRjQT7DdcGJx1QZoIbotde+fvBFib6mct5TuVS7iT
TUKt8TvX98ZSh5ELwsTBrF2iE+1wAoRJbJMC3JTRh3YlkWyU49OYMqs+KgPMIZ4AXSP0L7gW7yaE
WEW2tX0eTTXUzopPF5Vft2pDpCAYQ26UDerBlibb7H4ELR0oZjAdHYaBQ8bxsi+wX4XnX0ILNO9i
JyjAnp9uPd53uYUvOe6zIVu20ZA4Y6DlEpVzYgUsFOBFlpZ2obuQIdSHRl4lvSWo47X6eyLtIAdi
knQCnoUiERiDPMCXGEChpgVtca7WoN22CNTZignQ14Y6I/zZE04nbt3z9JSqmp6V+vqRgmQl4zTK
3X6rQ+cjPmtyUqMIcsvTyFq1WqN97BVwxKnjNPfrc93QsdtqGI1mgXQZGseGmNxUPYhEicUtiMAk
VeF4yjWDjHESCntuJDX0l37DiQK0acuz3LiBdjR5lCC9sTlt82u5ZapnEnIGkH/3FvfZbZeav9EK
QNzHxyho1cgWAhO3aBmV+6I7HeO44hxVmQZ4CTc3wtrdtXYIrN2gmUCzY4w18hjblR75AuX0q+lQ
fS1muqCNPbKYmEEVosVmq4uQ98KiUN87KbSqv93dL29TmurjafaJCUbxmmWCyAk7UNNnjdVvsamt
IvSAjlgK3MYiofxjPS9tLWtC0u/1gOEuRyk5GLYAvkVNmYzjjlzJsqs8/I3KLIATEKE5eoKgqcnM
PPf02tN2l2z9AGCWQuCMkgVWhcCfzH3+noZYQbm0B2Z+ZL1eJoquSAfIZ+41ucNgloe4UB85xlTB
QTYmSkEwzJgA7+Yr9qcyZGeYkJLkfUqZWB2ZQPgNabiFeJS+FupOaI2dbmMclkwMQF2L+kLo3B/D
PFg84S50beE1xb35qeb8/v408vlze1Haz8RNVGNZTeXPOttPZRGKJsa8XK0+6enf8GZPsji8UVJM
N7RM/ZLxXtm9XvU7maZYKiePjCvRx5HMwNe7nzhb6ezTGju7+hggyFhc1nJiQxYp6ibY7zaCdP16
wSnIgS24v3NfG2b9bTTu67FTJjoUZAgda7zvRmmag7CcNc5/JL4v9W+iINaYJoA1d4En0OgrV+pM
+3u12oaHr2yhFsXlKLy72/yqhCP5xOvgAdfPiTR++mH4Un4MgrdWuPY7WsIiBGnEf15m2ypQWsJN
CSXr1nKaTwCVpWgDGKQ4K54Q6Z3ywZwNlGXO+Z/dsxkSnsCXNQOUSLykYz2ujqBNIk3qATvcbCk8
oMJarcvTae3vOG3+aDNryrWBZeAHro8fzoVTJvbjnm8L/7hzWosXNZD/kBDWNPrKGBFzh79yHoEk
86E3TBjasXJI8+Gu6wsQ9QlbbguyTm3ZH5J6VZkhVUVSGTwHV9vYELVcG2Dynv+wpHOfrELhs90f
jP5SE4QhMGztrunLqg46WogTklDHbu04YbyAa/e4qOJAOnrRuaDeAMql+/U2/GQO/XuXYrwndIEU
RRnvEAv2WqXX/e1sC0+3WM0PKHS5RUyYJpEgobhlCEtM33jB5Pung8ncWeJX9g+AP414bgByeBf4
yOtd8Sb/OvTFNlgYuHdEWMeCrIAj+q/kPPlR0nW0GgZcET1dcWNusJaDjPe8J/XwjwcJxWCJnVGp
Yt62kLduvvjn5vQlhd3hLkusumTgFEaK0p0GJLUtDUFyJ6yE4w9htVW+q0D3vE7hQN27W4lZAPWU
kA5gFHYja+cdwdjYhgZtKf8WskHiUxmVF0sluj3YGm8ZaOAvyQ1rQZp/Cq9DXAbIFOGYnqZlHQFP
1dJ69COT5EBkjtt96FjGIR1x5EjSrqumo0JzANo6rHnPnGtIGUUNrmVBJoshfg/ZEw3nY791gz6e
xRVc56Df7jsOvqjq/lAga2wmQ+SzNBBuWiWtr4qmylyIKV3RqikIv3ZohK4S3H3ix6d4x2nppFL+
cNBIfrY6qnxDx6QKPVsz6PorKDNyHl/0a7kUL37GVvgyAQYFX2GaSOoitkSRPk5ZS3s7J6gsZJjn
Q+rgNvUqPBx4K1qxqYJ8Okrf4jMt2TeAAW0bHF/sL0OBAtc9n59IcwfL+myxp3pDVXLuqgf1qI5E
ri7u220sHuYy0ynOEi12/bgShG25gGnFH9nQe/iLQzexRM8OF3RF2Zzq8Neu5vlQqPNjnkRgESpU
781x5NHvchDKBT2wsbMmgGvf6oZUWpGNW6uu9A61nYfEgxYKMSZnPB8wMb0nrHeT6nnz37uFZpgr
0qjOzZJiYE3K32JR6d+9PYUn9g3+isaK2VGSjMI+OwpohUrGjQ6gBEQ/EoovRtI4pnUMQGs8Mo+m
qk9gK8nok12pO+12YZnNESkl6cY/+ItQ4I0J7A7us2uCpZtVVieKc/WQV68YGld7btS2zdVkuBRC
qr+aF+7MUnmXZoX6lsT2d7ZCV+7lIr7CZ1KThtyMGWLtwxMQK1XAZq6WksDB5BIfElUIJWjjerzG
wUoJWpzqu4I1JMK3KHLga2pVtOLCkkWE00r3VZjRuDAvLaxiDlEMwiZxKDJBAr+gm2a/nWNJBU1n
D2Nx4hzliLAN0CMTI5hm0QZ5l7pCVJbCie+3gUDfkMq9I7a27hNl7/4EMr10l6nMRD4Ky21AeXfv
cf6VOBwoAx024orgnSnTbj8qI1JArOdFZRPFLvrheh3gd1S++OeQfKwnlHlSx+EfjTvkfUW4ykzj
WsoMKnVRnnXALCSLy9tpYSj9CESvFovQFze2GM2fa6Z+pFl/h0OZXBsAt6Ousbyx7vttk+SoTiMu
rC8Pr/6gvkZCkrwh4QSqC5LRJX5jD7bBEM7r1UQ3EfuJnnxS6YkojtH2QeJQdlg8cHWGlaA/BwZy
NnnSO4T8d49hnQxyiZmLzD+y2TU3aXix1Al3T1xAFcx2eyrzwVtce2iBXWjMLNyrf4fhbqln0ZQz
5HGLoJQYcYQ6Ivx4uoeF0xG1BX+55Far4dSl9kSH3t72XwQJHjxLZrp1JuPVFKHIrfpUC5kpRvLn
cOOk0xWg6aSRihoc4H/q586aMJoTOU7PdFdghKP3drcVIewmKGZBJJFrh8yohnvQFZ7NjEcZIwss
oEQzyiOKyjdPk4av3LwkQ1Jyqn9CGWQXrcrHVwt6582o16nbdU16nQcJvkArgV3HKxnKei3SVYqK
YdNu5I7XoaWAayBsBkXbjCfuIoee1/eptC8aq9m04JSObCn71oFUWuZp5OsbehI3w0Quqb5jeQFo
QAvZdo79bvztY/x6ViukoM6E6EnZkJ8Oaip1Eh/XfrpgVkccfu5eXlM+WmcHHMs27aQjnS6n9ZTK
8rWl0NID1XroNFkQw5zMVbkFIy6vDk2Ci3gWKpjMasuQunBiMLrngdCAnIJP6QRk1N8yykjZWTf4
xRCVAOuTJSOxfsm6GO/P7MiYO3bvp6mfttPekj3q/R2VR1gHuYsHvuUOeTUYzgYbS/yBQNz6pkN8
Lawa0VZgcYmZRcKJ8SsUlx64rM4UgvmyU221ure0eYickTuPh/mTrdnM/+JRHtUw0BOhWJw69pjM
saSJrZR4z1YSFpigU9WZliPTwbvzIWtw69Gg07Kc0GJbSLzUeHdDzjJra7A8Q6sBFWYILOaN9cnU
EoFieO1mLk09rNVn8PKVhtiknF592Y+7OvMqva3EDTcavvfWOLE2jrzslRKAQsyspx8tbbveUwdH
D1FdPcnX7gwYptwySM9/ipFJ28Zwfio9RoYcpk/WeZ7hFm7OkTomududHK4woEHyL8QONuJ/EtkG
7IRha8PrU5ufhcq18BQX4FBHl/H8p+0XlokZ6jl7uv5W2FwqEvtL9DFPUwDCnNyqojo4SF7bPgCm
kUvq1/kPZav6+Bt5+sbJWCcu6XOJD4wH2snpKXJaBvy49frnto4HoBs8f2jyhIfzxA2rxdVNfkiK
Zckhk+1i9VRG2qC0THYS8LRSgo+bM4qZJu/jzADDAnNMMYyk0Q7Of+l/aO7PM5W/Eik+S/zSa8Zy
c1RSFltrK1d6s8sLzqeEvEb0fc829+3je3umgHc1IBFeN0j1k9sKp43xGaMP+Ni5zxuRCtU4bndI
g94W+gtKFIMoBnGH8pFisWrfUjps0JlcVDtqjAlbnZ5w2dlSIv+r+5+6nNGevZu5wL7qmjv5f+0t
BbsMH1xGG4kOlT5M2YzLpAE4Ct3L7o0zPKOTQQ+I+9eQ5NBzzbtSQbHPgJivuwlYxcl+7y6sGf0u
UqfGh+qD8e9dNOCi+sOsbVl3JnPywcl1SGAVKXla3XVTvFdnGKz29s/lDMlJwP4eCXUkUOkMKNIQ
cxph0hKy5Z/3Fs6Yt/GbFNoXzmlbCFDePYFv8u6MLf3mIRNoWUM1kNoSoWVyCafq0EBMNeZi5OsI
JqJuBqb4xw992eZUSI3T+BJKFMGueV3HDu+hxrtEOa5Hg9AizBiTEqIDMyWhDhYNhQG8iNEvjcBt
A5APYUXpTYyZeco3mKjDjXdKqDEXdTc9YfOJaAqj4X5SX5NZsk1FES1hULGPZFEKoTiy/0ATwk3h
KIC2dSHgH+XTeSegA0ssn+jTYU1SIvIr6Z1qiIBtSUqZUNohDK4o2ZpXovBNHkrkwigW2UZam8KO
To1zAV7SvGd6JL5Vmzw4nVTQMkprzBUvUwIZnITaKtAgJ6RztO8h9K/EzWP2o7z9l97bBtoscqs3
gdTQheI32nrHDmKqq13giuJC6IRfmFyk1MmjqFnlcp/2DlIoIm3A0Nv0/FonG/x0nLfd59Xfoltj
dVVRh7Wjv8MevXaFPb0UG74Xd5wo8ICZpjR+VMfGcfwT1gAZcBVyADEH6LtFkzXodkir0AzfPZxS
5pCQBMMtgYjQvu3DVVyTn1WeC+7sArkHx3wHXCijHrglVym/OXj04vPe7AnRGTmnJ4tF8GEdf0Lw
hnWsm5PRu5ilIHDYzp6X/T8pRy5G2QUMF/xTE8V7x4uql9kpdIGAfwDiTZXE5r16Fs/LBgMtkcQ/
Z0yXoelx2RFMsvZqLr3GFqOJyHhLktmqKobTf3rwoMEFukXwCEBmAWjinOTAWFak88jG6RZBf4K9
gjShqiMb94rsgw2v2bPGUv7DFexEqezVkiVI1Dpz7yOMtYgyDF93JYxRTXWUtaAX27HPtA6U2S0Z
am32Q4PhgJe3K2sznmNXlrxyWbXG3n1Ula07tG94Oks9hWbbYCMS9Upo07WhqLKOkIu5fOXthN2M
FH25eTREkMBFZPtvAoyDq0mvuoSKFVItvmxr1b5i8mrOJ9JX85Z9YAbm5pP3j4O+0kXrD+ilmElN
XFeTf4oXHV9Sa7KzrIoUysAJQ5N/O5A1U7SLXbCnTjA4lfe45XBXiyEbXePIlXJTOOPWvcuF8Icy
xim0vYrtdBmeR+4rjdzZod5Mi+FWywTjlrVfiwzvilagh0Mpocds1qPjHQ3KSQkcWIeqjThqFRti
04ePmtiZug5PBpnY8F5i/wENC1sRHLfL2ph7xLD4U0x8qdjR/VskdhIG3ANLINue//JiXaeaRMJb
1lYODrFEvDg7f7fCQsWk+uNv+HsKOap+/o/LTcVlkSK+pRJvDb6pfSG5D+vOGpPhwDpCzzj1nP1R
IZgEeya40t8EC2PzEHnoyOnmBBj4KeXrALSiRW+bEEouv8c/mQ4qHukB5981ynsPrUeNfS4EyMOI
W6vSEtIOas33P7oFk9Mp4t8kWH6TtnLr78XlX7P1hFxa6YLoyTrbndCDjkC+KdDDNgFNfyQYsXcq
IDnSwehWtwp072XE9QCqYon/PG0fA6cAP6WE0VQjeGyRLjQSsZRn50gWw31HljqVaE+C7shw75fM
nTjcjidpeVTPL7lL7sr/zq8mEsjcCiG7JYgSi5xer+3jaV8sAKLggXeUZ4QzYrzOuW2CxNeuv00v
WRgIOGSz3WHuqau8dXYpNezOBx2BAeUUfrYGkkapLLx0+QdxRaD7gPYZcGRG92/uKR1gJR/Jj9O3
Wf5UUpDQdUbIQAU/mvBt5GWohSxQJo0jM1UscYiZaF8WFmTusB6wv91pW0Sm8gAzQ+PkN3FTnp90
mQkuOreAHk+B41vMJ2ZBsyo2rJJpyCTgo23Fb8kCRr0JQA233y7JeVW5YfephLGHj6i8VZFiVgrd
RVIvRucASJaocWE45rloJsjkqhuHXMbvqscDmhhCK+qorMV5MAxlnG+fT+RaLD2jrQcffyoz6KtP
zBTDK3QucceHT1IRQXb6ppCA3BM5O1FJDdeHDEUmWZG21asLF7XrvK3YzTn861Vv0WQcYPoSbewW
wKoMAHQQ3gnyu6CGfPx87aMYHIhMlwUjTfxAAcE0KbQyqG1TdmDu5g9vpynSof/4BdmKBAOWolhl
yzR2SLxPfQ7eQjtobH+pVEraGu8ourG+HH3mXdOQGQX/Q+qVpAjKGVNqZnbyjGipAZ92vBCFBdja
zZ+LxkJUFWnwOWS0yGyhT/0ylMSuuRdi4tRSlymWRhcdnvLmN8NZs9bMK3vvurMkPOrNrvZkahmb
TG96lQVrwjz/81lSKqturPMv2HaXY1s7SefSH/6s7vxnK/ezL7kT2rIokvgesnTRdw6JhJYSEIN2
B6x791N1jxyWfo7EPfovNHoEE90r1fcnQnQ8J3/GOtuKvc+xPoI9Ac1rrtKT4m12Oak7DEQ7DB7n
UyKBCpOrlfVbx6hX3Quz7W/S0py+OJt0UHaoAB4MkL1vWnRG1Z38vm0UNKRUcAIKOStXdKnP+25W
16+CHpdKhhPWOc/JUtaFSfzsuKAuJkfCWcL2ECMTBT6ndfA+kuUbwQdjmVo5s170EOuqAPgU25jK
GHPD7YU25hE8jdhcAqWBgGJvLBXA3gKltMGrz3kwsMZwXXT2IZY5zbJhhDn586IoZR66lkVtDJEf
HCVJFu1b3qug3KuT+DMvM99kugkzj/DRvdRNEESbrS5aKKwfvUnrswJ5Rv+IXtVQkmCwJ4DLzYva
Mjkgtyyq4EAAZBdghFrHaFBfHSnlU5Z1MskWuNovJA/HboqflN1Nqorp84SIAhigGpTJYU5z2H+i
2SPMt8yGfFmZmQn5WZrM8HMt6I5So7sK9G4TtqMsKkFwSsLPb8dNYxSX3eITh7sSyd6FriGjmRc8
pczPgvqu3mnzF0x/mxgVHHt8RET+4AVRSxnAp+a2ppSt6E5nAIUwe+0m1AF0YONbJba5Zsm84WuX
VXu7q9k4zrxJ5/kkDYmfn01cV6TyJ/C7xVNfbrdrkWaUTAG7ToJp0CSGKCkj85knqf5gXuy4PeS2
htNMN99IBS3TnuCpOSmvVPD4kw8COe3T6Uluz7ypWlcWQgMb4cArvak785jOLK87YOS3KXF37Njj
S8z6YbSvo9hGGY8JCxjGSfDjCKbRZ0BxsuCuBQISN/p3lFv4Shtjy1ZqAwDkACabZZ2XCNKJEs5H
OPFhff3lBhU1IrEy6Fw4VocdXg/04lM48D5WV2vK/rJIoq6sawNpTQEPtxBBPEuZ+f6VzHDl+WxW
+u+yOvLHXoBLllALH8unIcggwb+Iu6Db7+dMONF9iLDYs/Yme42lX5/IFe6d3dzikQsEfZxve9q/
flusxsiGf+92ir00c0wEZ3LNqCl9IMPC3GrXKg+t7Umq9bVgelfWtJtE5kNdMXlMGnbXkodqU+jm
nEBhNwykrVVe2dw1Weict+wu07nyXGXp1S/6uf9mkVXp9aXuLzCAN1/x/AcjhKlXg2hI0wgLb0JR
CcQkP8H0Uk8Y1GMI8ZI4s+J3cg+GRcpLi1lsvrXbPRJPIaD5EWVPcGRQedUl9cKBxYaBY3m2HITW
QLu2JcwQBBxUq3N1g3q22t+NjCsQJq9xXeFIbH2idvOve1zW3EgGX6FlSdFiXPDVMmEIR3aqV+vr
wEtqwkxWp4YeHDkySHt9hjs36Lh8qGLncy3uAMdO6HaTuaR1mHlz2y7t5U+FDjADsBX+hQimoxF5
bgsPa/H9E31nwOYrjuX82aif3/NfdnDJTTWKoeB/zaLHHyQ2JouHD0tivnTLCBSuGgQHjaJwzOne
uaShfQ2ie7GtirAdmdm9xqoEDmeuQ9sR9C6XBOVzLiM6HISs+319h/QDFbsaGqzJi98YO2ilAE5p
4W+a/WZeLI7ztm2Z9ieFKtnRrbee7jDDyt8vE7BD/VIx0KYyrfVp3InGOvupjOlleGeHrQthFod/
DW+xFygraS7Uktmx5FrbQtTvfwd5WpYzzl+89MkEVgphnoElad4JdYypE3TpyKZqU31tOkPxeqWS
GQZiic+dwAdINSwP06hzZs9ECmqu1W/uk/0hywqMV5voMdTOciRp8x4EDCSlZkr09fPJHHdwePck
TmK48extwslfN+BmFHp6ecCBkHaRG8WE9MeA8JRoMmHyH6z+v1EL62YNWZkrtFMVKT2bX+0LvvpC
VWZIcaO1UrutUlqy25Kcr7SDJ3qg1ZL98Ahg2QCe3/ZzsjmxNd4/1Ul/on8gIxOM1B58oZSJ5Eq9
TYkMFtQj+qoRR7tix4XErwmBFAu4PfOODTod2N5FbsLxWhsAfZ3kKymaVsrwAQ0uO74JhLjPdHAd
+9iqoaC5lZ1UsFZ7q9YA5f4FbQvbbLh42qDPsH9M8ymfg+YOXoWGQGoVNswO7OcGs1fEBr0xPr6+
s9pZlEZgqB+A56O3sE4Ic8ROOi76LO64h9hzoyylBExFu213R4lTmHGsh5tqv5mCxOk+V7/nB/jt
2QKppsBu5lKZg6/FtA2gxf1GjEnzWeMjzhGTHBl63QVOTDKBelESVFNyhcJ/ESlmhcanisdxfrwF
j6mvDz065mx9D9kHhE6BfszBopDTjduDRSGgLVl7xvyFRXabBkfXF3C3r9B/eDF8mvVRDO2pdRGr
F6Q952BCpjrSsBsKkG3hq4SlaFQXiJD4DqTVU2rxEsXNGVa3wb7FSVTbxhdGzarIDhVzY5Ib18fj
LZCXr8Rb75u/0z4uJ+HN4iQEF7I2oO4em0z2xJFmbBNwE1pK/d439otsgAOy6vnV/jIrf8PyjXkx
Fbgft8CpqXWI/UaFhtn+FivpwQlcASX/MEgA3iKTeXTpM/TF4ueggzexk32pTSHfyL2ChKnRA4wT
FxZEEG3tlHgjkacnuGaujmcvosnZc6sM/YdDWmuClsJO/pMeCYZH22Dp7Agim2ot310McHzsqiMB
2s9H5P9DYNd+hNS8aWxuulHz+PBG63H5Q62NyhGWmpLhpLu7BqdV0WP+b1M194B8O2NSLwKSUfZH
GsM7X4w/xVTeAPsK/0LnpD11Pd0TaUpvFomRAFGIWw6kQnmVY5XCrlYBARpbqGjgg269m34KW0t8
fJgseLF3BX+kNufmcV6i1BvNyOB90X9mYctTyQWD5OZdbiczsHW6D8CCaGSqNNQHwPtuKugMMDwm
2fTRlGC032SS2Xpv8jO8remmLVjWSMOaNDAyAMbGF5FoQmNYn6H8EBJbv/PSoi3yip1oWYSMwKu1
EtbVV1PZU3GfwyJnqIyJkmRvM4DA7KO3wOIPJA1YN4TbCEhdMGsA+84W1365Er7hCJaxmplDstKY
4AeF3iy4W/4080yjHXMgNx0q/Xi4s0g+3y0oH5KWVHSZ0xhsKhEuQicxXJ/5+ptEz3CDTGOIFmtn
KL/ZXMvOpNGhTMbYUST4zdMzUss/PowUZLpxBS1rsvm+h9viqI5d/GrBdsNpQaQ4oG2TSQctgFnU
u55QOnBm8Y73uM/tfLUmmpQfBFKyIQpR6zYYZ0rmtGXlN7XxuvUSdQsmUofYzlU8mQ8PNHIf+Oct
n5k9p8sunu+KcPAFh57IXs7upcWJDqvMr/w8PW67Eh3KiSTcvlxZhn4bdl4KK28pm7Kc1RMkSg9z
au4ybwptoEp4caQMUT7IgPYVRIYsVpu/H3D4OITkbVDYHFmPM1eRqINfJJ89v5v7gn60eQx5AQDd
HUzrbfPbxrFd6WabLb0CzFUQkWspyPtk2z/w1iGqp811YjEY93XsafsZ7CkLlzWTTmefTd08T/j4
q/LDFoLiL9jgA5TYIwWqqFJjFjxlAEdffvBmEmX8GXwynUEE56lJmtIOyHO4erO6TWNWHO9qe0Ec
gcso7u4M0lR1o1I50w8jGYFachxOftfKC8/uabBHZZeGylrFzEMIQ+eUB3Oq5vIXzNxXqIPrph+/
sadn/vkFgxrD+pfKxh/t+ygTvIf/r5YoJRf+lzyMQ7MhUbwt/QbhiLsl4NrOF73nPtvp1BlanrsH
yunoXvPzssWPTtkP5p+UptmUayOCaSda/zwFLGg86Zb9rbo1Rl5SZHXrJuBkFkpsrjWSk/qwHeo3
khesUZ/MRMpdr1Xr1/bvfYZi/cF+DsgksvYWsEX4pXXQyFfrz3eGFhaJN7rgpKvsOrJ758bc0Hmp
WKX5o0mO1ieI7XxWXcS//fOT/6VRPF7Z/rpGDlrVDGe96RJSvqc0DsiBcE8J6w1TVUTq32HqPNal
6jBLiHxEnkkGWgWW0mIn1FcfAI1Ac+Esy4uIqMtgqCuHSauO5XnMBrxL6m7F+jPtBmxZZ0BNX5gR
PmZTxF9JLFYn4LijzKTTeJ+8qbQ6COXP0zEsA00s1tMtrTCibx2MFlj1bR2rVFX0cK3M8m1j8Qlz
UeljVBjkxBX3t+7e00ypWe30ZRmM3XRy+fifXD1+SNyL/D70W99oo2dWN5Ui2VhTkhw3gMu5xWi9
Qt2hxsXg0SGRSupTNmQrzFcfc5xUPaddkXYAc0jXqInseQT3Xz8cH6drhu/LDXjsTV3RwwPoYlgz
ED3r4HB30ZGZbeIRQUgKXiMKklFRfTsslbBLNmIrmEJtcn2RXGJ8gielfNIzuTAv8ocj9rJRaPzq
z0PzDCbWtQmXdOZT1wyymAvmr2MO7FQd0kIiq1AiNMlWGAY/prK905Bi1Ai1o3kjwKpVy4y1fDR1
pYOSdR/W8FxC8AHBjuE6J9hDPe5OQCKVggGuZgOk6LE4sPqtTxT+pCCLY6QV5Bn6lBD4KGyfghub
jh+sgmf1JWuIi8RtJIRp4jDEFfeQuqiabSfZKKtXN8dEeh0HQ8FTZPNkpa22VwDzbN06EnQFABy8
cBjecL6a1OV4i8uRQot1ilCgwnsjx2n5+CDl9MSoLAnKjRql1bAhQD5aGQvU1g3VTAbEHcMe431n
R+Ttob8UNc9L+bkxM/VegIPOs9q5QwwRwmaxmpo+qZqaZtmZRBFZUmOd/80D3NWW4aJtbkXGDtZ+
7HM4G9jsGDcma5Qe0iv1ez399OgFWUcBNw56uqn9lbpY+d9ruIQsXxHfeR5d0FumV0LE14u3+7cE
z04pyRTmaaM+HbRHl9ZNL5gb3InjTjjvVWjGRk3V24+rs6RwKyaOgoyZwv1ZCoArrDC4FL9YBfJC
pFPupU8WRDNmmAC7y3Mhjml6PANymBg1xKhvCBig0NIwr1awgYcO74mr1nVZHh4+t0IzbqP5ZLyS
/FNgTVw6H6qN6cwBIpp8Yp96tI1QyX2a9T6U6gxSfHkx83SXE92Rmsh/lGe4uAzsDlZih/d6HvP3
seqWn38J+xBlbz4DQVT/mtD5GRbPQ9IdMNOQ51deMPlpdW5Jl9OfFOYcPNoLZD1peh27JkKqAkWG
a/OV9G0+RbWHA3dKa9gGa89YYdxvaiR9WBl+UZSlIFB5JWFdE4ja+OzjNeyosOnUTnjLp/7RqugR
YEfB3R8jMO3rKteOBD0+tRMhkGbqVW93RfRDXpUsbrMHv2FBVZOTQ7iA29rJQPR7M3wE++bLn3Cy
ba4bP86l8Nb3XYuRKHpmvmJHlf5n1R+fUackRtcdUj4aLKg5GAJ+lyLqD5t917v39U0NzVd03pPc
hoLdPo50Fm4vR5L7/om6FCQtQUAsFKdfUVzmU71sWaxsvB5ihbb+htozMvG+P8Gu0QjbHvGFQBes
9PWEth6fXbpvMSlIp3S5Oa1ASBQW9cG5vM4Qix7QtMu+fEKiDchT4sowJ1r2eSvzCNvPNuZxPQL0
Kjiy3ZI8IwA/QNDvY65tHddlvb14S2ZJHSz2ppwUBl5CZNGxi/OA7CLj9EndJEariO6WDergsCgD
eK8xCFTXwMRRX9EtfLi8m1tlmRqu91+n+eYpWcffrYO1ZzKZTxEjT1xuZ2s4p1AlJcP1aT5Bsoda
eGEiGon9M6zt1dFTIMKiVSNvfcLRgbMjwZ4YJE5lI6NruZ592gyYsmJpSYAjp0fJTAnoiPfwUAFO
+COEIbtrdUMBr7GxsBgJKBZYc9H9z6bmpQzuYxMeNCmPz8HVXAoqfTGYySp7GMAzloZY3QmIv6rJ
UUJD9ller/34OwSLn2ZxK01o+gSLN5I3btgcs9LoL2GRbgO/eFyyvbvV3KI7+cXTrfbIP6fBD5dB
zQa6yOS1Y0dtumSGv9nyk23z2FX97fOpiBQNTvjhluTGfAkcYUzm9eBowPvjA06tt9x4qH4l2Ars
nbF520WDHxMg0e9TOIfKWZ3W+v2tAYF58f5jKih1LPIBXVipsZPs5UWUT4aU220A5r9rnDv1z1pm
AwIYTSNW8NHx7W/zOwZgaIkoPEOcSqospO8Sghk90A7nlKFy68hh4vK6eVva2hJDFM66nbLKNJG5
wyMJkda4vOnoUSLQtNoMoZyO1W3xWQUehdceDaZa/7mutCMGLyZHJAhepMS1Z2SaZn8xLA+FE1MM
NxEVXoN7X77Eld6UEQUlCKbx8TPmE0JUgaJSlkM9DEzKETZFyAsvLFgom3cc9l6mzU5foUkJMqnU
eWZ9AjTYGb6O0fEF6JX1v9Q5Z/hLa76Nus4drsZLT+ko86RezgSLcjWnN0gLiSmKnv32IH+gaOzP
WYlcHaI5/oBTwOdgF8BzO6QqFxeNPsZu/0/1OOxvhfhwm3WlOsPOKdiJHQ0LmU4gOGzVvpcpfRp4
zMnJe1UeFohJIYN39tse+B0n9ca8Mp8zs1ek8i24u9UsdLczrRTFDESDhxfdKlcS7djUnhV5ejZJ
DqL+PF6fMe1k9sywqptALY9Zn8arZzgPSK/+g09J2sfdI6PEjqocAMjirYy8uKPgV45WMvCRtbC8
e+A6RkrRk8+Ljs+QW9FHUTU1ftTdWuK7y0uEKFIeXL8rixTXAt5LmaDVUkIjJ/qHQODpAdrAkSZQ
KKULvlwe4KqTUwrHLeWAEhcEm6h8bgnBxDMixI9hq5atI0V9nBfkOKWHrPV6ybv9gGbdBs48iuRJ
07HY+V1BlNqxh7oEoi0JX+LYNbqiI6WCMyJImw1EcnPqo/FtKpwhALKsBTxDxfnnTan2rpGUTvE7
fa/g1Wj7CEeyZmy1lYlsh4iCTB5NRminiebsHb2nEYtod0ESDZHlC2rPSatcmrPTn9fEFQ1X7a6v
2nwikH04P6R3o7HUS+W2MFEGgrENbvPUJ84thf5rsqorMEMyclyZ3AKRcvUhe2e531Eqlqy4zuuH
Uplzz7sf8ROF5J5IQ9DKMFxUokea0ZeDqvaKnOQ9pylQl9kOwzQSUzacAlgDOjsXolA2tiiN6Ij/
sBItkEGmI5rHpoWDKQpi84GStzBaWmPpUD547u0WKI8DbKB1ABwMqSEvBKtsj04JutfTapeblkyl
UTXNsrvOVplbdupEe562vyGaJb9aypbNWL79X+9x1zb9UWqHNd6YdV8CNTSEtYHsOg95mbOzIG/l
d/c2d1Wo3nPnGXmx67bmjORHnBQOEM8FOdIoPFNCFfSiDJz2Pd+/bDI3p15mNAVmdqJiZZrRsTzX
qBELufDnAUHsVCZszqDX7raMu61VQV9GcVC6qWWoEa1WuMmGl3yFGRWVNgJJTtUTLgcrO0cmP9uA
Ilit72sr8FVwCPxWiuDJzBr9gNdLgaaVtKChqv16Yx3Q1p17xt1olQdlYbSyA9HyXejzNa/rESJo
9g4AFCqf76pOlsEUpnF9lONv10UlA3BxlsEzod5f8jBNRuGuCOqdSMt+dkYvrIiCKMT0aDMDkd1i
PcMVKD73Ru0AZOfviDw67Xdk9RpkydMffbAobf0PUVv1W8Ngp7er4qAEnOv3STPSjatdlE/odlaq
4o6be8Y56yrBJ2J+vEwc3iJ1ggGLXHqUA7DSJ3/VthsqKblMEQxjSasFlSiwsTN5m1iKLKCzZyy3
s4bcOYJGRzdjVyic4wnAdBfjkGJBq0Nq8y1NsOLSQ/Ql6bBTZLgeEu0FpfmjkqBi1ZpXRGIoumIp
EPDAMVYlbrBkOOzfK6ckCVW2fAVvokT+sU/DoW824tn3iOZaertbzHCp16ROGkLZWPoNJ992PdpK
y/MgmrKT5S5zT48q+TVs7A0A6laqbfkJc6Y4lAGDOLO2+UF3HB4Q+qtjNmjJupwYy+9WUSFcZwr9
flgpfTXxG5AqYJp4fGLvwWpum0tz/4pLqxk13EFNm0Vhyf+ss8jy4WZ6B62xpjOOFH/FuQd88fkz
aOmIwc5QpKDHOxqUaQ+20L6Qgp+tBXGoWz0YGjJBPIjktOOYjT47CNjY82Gwis+9DRzy4b5q3md3
d0tfXEE1pIZW5UKFskXvhkkDinsuHFpOecFJel+pH9hVrAQ/wbMZgwAhExugEipxXls+AEZmzkom
ftd/swzGyJuuH3rRZpP+v5LA1QRsHpYm4vRyDu5RA08A9BYYvRoPSIUdijGXGH9Gf/vGbNTprtso
oejHCg8Tqol1wwVGM8gDqBt33TCV4/1C52LIK8hYraBUST8JzM5PGI+gmRtfhe4L19CrXgmQ9aFi
Q20Fe8eKvjLoqnbclLo218WZx0FXGTzqAkQ1LzkGHEZr+MvacEWZNMc0k38XcpN9d5GIIjsJwvZq
M/pNnQRzoISIEgl5rqXw2DBG3R4Im50Z5UChZzwAere1OzVM4zVVmh8Z1+kpyKfvT6yKBOG11/2T
wHiKdQ9RlZ5fZmt0vbcm1Nqxxkp6m4ih+TTqW1abK00/Y26XkFMxkARKu6tBUJDuNzxkc0yRiEd2
RzCQbSlOC8J7QPjgAC/k/bNus0XwoduaIOKu0+t5RwgwAeyHLG9RO4slBlX84FOEO689J7ONA+tZ
rksCZmOfvqR3w4al31ypetQnZQltaXfti+5ruPAiaWBu9TTV+5R+twNOCCqzWv7PvLzgwfmS1dOP
Zj9huBJBFAUJXOoCJBZmf5iznOH9UBjTbDsAKs70eOlHqAylAhpWJdxWe7UMBlEugy1++jc7+cI5
TNlut3MiqooCuG0mYdc5iYywbmGfEhMin+jnAkQ+aHxNkzzX/HGuA6jrAckml7FidxuloCa7w3pZ
73aQLun6qwpA8Se9L7R93mKQ5iMmmqLHw0DYOFTh2BqbJv+//karuUx5MtLd4cK+cWIPXXDzLd3g
KI0cxoKfCwN0fE99Mivf8YkMa83eHfJ8yHByOW3lt2cJQye0kCA2P9TVzhaT9XfoXt8UaH5+YUMP
ybz30jVTP+Hf65AupbRb5i3dhw38bDtlTYehViQH0tlVsetJAKL6jTF1ZjbQn/7/aHIMLhbqoTbf
eEVLPdGTytAvE0jeBGq/CxaEdbEQZA5YEL9h7/tmCffgrfQ2fIKGiHvdGplPTBModKDJOPvDcXL9
Ehr5J80pYiTNpq5PQDkyjI0Swk3tdPqq1Mbx8D6uHMAcrxbl/RXgAUqf6QOr7OiC77jyBVjr7DVq
z5Vgo/uZguIcFP3F6/9K+iT3BgwWypaTmAx3w+KL/cCME+mpwhjnPUAZj5rGwx77PDFCuhiNlSbj
k9c6X5Lztl7Y5utpShFqOgZC3GpCverYrNgjHfygTC/qVmbuK7Bl4ExkKqEU5UC2JcqTA3SF57i7
vt2YdP8BLgtULtKq9qgjiGupR+VlU68Dj5iGlAUpC+RtsfXOF3SYOAbW1v4tpaTtUY0ToTKXHRHA
jLhjub69R3bEfKOpfN2XO1q2k9FNo9XPUFNxnSG3VxhJuNacQb4dRK2cti+A+GKI0Lahef+86q+X
/SSiNCzT7QTFcDHr998t8nqIyWlVkXvmAJksrmCvD/ethWwIsccZPOvZCGVBQDLnnQgguQoGkklH
do8MUmnijdEkbjHCjnA+XWgkOiN2Y/U8QcsiHz6QJJibyO7yqKXh+QzLPl2OEvCImx0jCHSiQ9Q0
LN5SkXz61RG8rmKeDQ2p8QPR4ddHRg/JnY5beS0R+U/Nc9Ey0CFU5/KPbhfl3d2Twd7JSqxDdM6f
ClZsGb3bnVkQxc4niPJvEy0D1jYaOibUpKnGMcAWJm12a9IriBJgAdXWCmP/sEnBFNPyPZn87bFK
CcDYeYraVN0q7s7GCI/p14YdDNT3zl0Y57hsmCt347W5vNrrCHFpupnfPkPQx8nJdq2B6JS1+arN
Z1OeGxCspX6yVdqKVekYPGlnFVIpYHsnRXbD/IPmJ19V+kRPDiBsrqf07ZzdALRavTIXPWzzdIAV
LMZGeobM6fPLK+Vsx+3KH6tcmM4XmhoUnGXwI1L1kk7gKXjrGSQQ/dcuY4VWR3m8oflv3FuY9/rA
uzFeyFSDhA0CP1SraJhPwLfepthFgGpc04hcNvP5Uo8+OtMOc0n93Z0Gty8H0omaWdcBs+23gUGq
8FjeyT1mNDbixphbb5Wc75rONaQkQ32pRmW2R1GQ/jQggfCRshbyabPBVe1GzOF6ng/t9Vgqukx0
a/gQ3TEDdk/Z0UWmDpuwAIzZ0o50k6Hj8GVwVm46rpbIRZ1FLQqm82OAffYdh1IHWfMI3gBUKVb8
4P7X484G0zKcPlZSlahDgyVhwLYVfFUP2L4YifsSVZ9RUNwW4/KFHzqXOkx7lO9N9zmcuWuQ27uX
6JG5P66/KUUb5cvaDT+UMZcR2AibLCDEHGU06O4iuza5S4O53AUZ6JW46DKz6NkwXeNEUhUQWLV3
w8dtaL+m4e0/dRszNhR0GCQAhnqx8JxkbysWSZFcpctCN/Y/l2RRgM/m5E4AY2kteNE8v0EU6S/V
HHpcW5m/KuznOkSoioO9WxwGQkRc/2lDksKct9pX1QnIw6vUXx0u9aW1U9xzB7STm5p9+fLnWCKw
PJM+Xnbzh7ARMnoDacJKc5uE+F9N75GawaYnEITMmleqU/VZRr4VqV7vrXb/Umfrdu7fGtUZVA8q
WNosMR+NKGkD+Ul3IqdgI/LdaihuScQczcWUFx6Hzr20Zhf9vvgyHrscl3L1Ff7Yy5ox9krokXCl
D7OKPQbulfmiebQq6wMi/OrlVcmjFwRX2WzPgFDG5FDIVpOCJ5xQKttIyIYSg/phM5qTlEKPVUO/
j4bk/iA/r1AbcpwdaLI5GJfMTrSSE5g0/U67RTdo7Q3XRjBNXfCHo1lXUz++xi0cYK03E+1HSWcO
TAnO/1SDq6oO4HgG+YbYNOnCNyKKmJfdmH6fYY3xo+a3XrF9sab1RVOrafEx/sqcxkjqKJ7NYPNF
TTmcX17dhRphaw/mI+k59DpJVPQjeWMtQ27IvVoVfiiVpnjm+LEFBnJOHR14/bQwjch2MOQ/u8en
N6/BQ6LJ73/R1XN6xIKOLapAbPQmeJiBDLYij+dQoUCX2g2fym5HMxr6rHBTq1dAvPkVa7M72fWJ
H7q8uKGq5zvMKa6OLdSRYNNKNQslFbuvSSNQwECvzfe5e8ITTGM4H+9J62CgMCxl9vR32UVDj0Ak
xGXQXzsaz/Mgskw21XWWYDFTeLsThicLjdQKSvjqLxKVf6RqazraStsHY2x8doFuDC+71QNNLkQs
ea2njmJVs9e0JIGkalTjUTQOQTXxuopnfYg+aizpz4M3dcyqicC4b0tw4fJyApKpIerhUBEKGQXd
JuPj3/fPCZSIUr5ELDEXoSOp9sWtTsOciad90/Oi3mMPomNnJi6plaYdku+yfIi/QftFHLcllg+9
h6lv8E/IpuOSAXNScI1AQyw92jUtQqw92jOqoY+FHtLVzrADSKY1NvdF6gQVCwmMdMyaFxP33+6m
bH3uyIQdYtMSRDyEOUxLNiLMEypDqXEC+bTkmWRP5XpkL7ZuwYLD7hCMkV8BIoGvFrSqu4z5Xp2E
hxz2X0+IGmNzkZg1VpLgEMbC4JtYE9mDcgscPOCPgNiPNfOeZzD/PRpQw2w6Mjn33wluztS4hsfM
+YLYJ57QRPWbAY6Czrt4Q68otLHSVa/zjtAGgYGEu8XU1ILxlFw07WOQb7Y4jiv15pHn/czuy2lG
S/18APdG8msdD00xYHWte1K5YHIMvWMuwbia3KPmDw9CTk3XylrpZX4Sz6BFOgtqJ98xvrHwEv/A
EJhJ6mXwtX0eyfovZy2mlrYXd5YNIjI18e1TBz9AL9AIi9eyH30fdJ16ABpPCpW5JMB+MKifxX/e
l7Qxt7JlzfUBSyXwZIs/06o5z+agN7nGtyhtz30hnjzXWRTR39uBpl7V7QkwjigGgu92WUGRc+FL
HDfSzQauSSBzr6NUdLxqIuU3nIs70MVLmQY2xahXgynHhiHIRkOqKmjIqy3doymYb2g7Z7Dan0PT
sklXDBKk1Xba+4RVw0CZYUhvyGOhOcOf9AKVIxc9pwgo7XlqkafCNDxvHSgjnyoQPUgGedGySNNN
C0M+QrEoV1f7QXApjHDPz8hGrdG6gV/4OFRyeaW/K9LfDRewglKD7v2KkEndVozmgAP8jc44Mrqm
40UoBmBibJi3qWWp5Dh3nSGV8l85KofvBYj/Qh2QhL2EJelPBIcDVp+ZURJjPnLWigQLrEZtCA+8
k9VTIoaGpr+sYkgGlrFfTXXTWFyBOl9bWQotwxrsrh2cPkv58dfwqSEYk/sSOheZ/mbUDmMH0FuE
wykxlphVYMPff58MVbabqRJNZX6WK8R1rToksb1/udrLXlSQG83TkIkDEHT2OYGKXS9s+Rqwfmbo
KilvWT2FTSrfk3zkzpPHHrdtpOcoKMT97Z763oSoTGia26CwyB3A5U/WLPezuKhlvFzyNB6Jk8fm
7aYIryHvVARO90mf7X65AO5HkrrnRPp9m/l/IlkW2OFhPfKn/QzcLp7/BHHA8PzkxEs8YFxAvly4
Jp4LvhppdaOgtk3mJ68HIXxb/ePL9xETgcqvy1s5f0U2Y8j8ohNc+SxUw0VaiiT/hOqWCgMhuBlx
TOXCB+IgMyxqAKZqBvwAb6f2rO9okunWVgncsCgmr2eW7psm4esucG7cl7Jcok0vx8JAW9mNRuiU
lTPaVuSX5o94OUNRlN8t2YD1Ome7ajyu8tsVy3mWeofl4/zs9IHJwDgDmb6Yi60JRT6M9AlDZNT3
kkp4lD5DeEOd+P3J0j5dLzRXsVY4Py5K+cci11m8GjWaPOY7pGXCBwvu1dQn30hTwinsLSl5HEWa
B4Uq5EGdHfC+64VVR+YnNjVAWWunTnH4BGeKiMwrMjGSUAcyKr7fgWZehei1ngeTIhYaIxWDnYuA
U2NR+wt/WfOD6FJ7bAq5kYAtWgvSVGCSEcU6GuLsrNGZUGishFEXtGvV16aIXZ7B/O33SKwKCrJc
s9qaylBxybaC/GPf5Jnn2Mg22AU/RfAuRIs6Bq86jVNQToFtJaVRi9jiaNt9zE3yYnljCqiDnELT
GoO4nJfavb/1Q/ROZGkXqFxt17N+wiS41ye9Ht3dcZoVxJy5hd7ogKNOSSXHaloFpNJvAzD70etM
tOl8ehnYNhHfSzZyJP0basZ7/FbySki0tpgVvoNQcm9cRfbFfjaSRDHULZCSluasM6cjILJCPQun
lieWJ4ged8QkjOiHPc9rw6s+xGc9qwtFZDmyZkLfUmbq544A63BoyviSAbUuKPeDP8/3fFH6Z/xu
2/7UG8zsvyeqvP5UVyenpo1heJXUUrJ3B3AC1Ktvya/TCNvc6hsAgIg8jSTq/efpROhWa8aIhGGu
bY9XJ+c0I7pkU7rd5TtfmbBLn+bHQqNIr62eqckzc3jfKzNOUNWzplucej7FUD2PM2P47Qbx3nkJ
XwCBWN7+L9zGp61wNF5bQTxa/v+PM9pW/4cmHo/CYEvOUFpGlgmdVppkm/gXUApv6CbJuT+MXe0e
L7H9KwoVgbd5oar1MOnacveOd1NnM5AWS/sf6s11SdrJgLLPYdBq7zDGjY8KvuIvGvXUiJs5TLLx
Tgp5zX+feoeraD1nU+dsmm5zOQ9BC2Mc76EtMd4SJWdT2m9CJSsc/LOcEc977thZH25lr+aS9Qoo
EcHeyHVRYPCX4pSJRly/iUOMVqzlCJ23qbP+gUcLbKkls7DhnLn0hYT7m+hY8jvXfat7RY78fpYq
6u62JG0B7jdQNQ/7Y6WuG0Tz3TW7wCObpHA+TJyj2lz8CAyHJzPyUO8IvWxJSPp2MhhyQExMeAZM
QY0+2FtCUDBG3ca1QRA7VbRtyhRpb2cOixik2hcVM7MqvUIalMBmHWft0/RB85r4s2j5+4ZgSVVH
BWXzAtmWV2FLLRFW6rbjbO5vuJnAcGKCY/30bi5kJaIxA0Av7C8QK51XJ1jczvxH0foz942XKEwY
JjbwCZg6KLLksPY3R88WtVrzNhV4T4CFpS+Hq8/dDP/rDGM0IIlitbD9tTmbXzFGu/gorsvQwRW0
npHiYPnNTZrrq8aTmzxHRih09YiFDhJtWS6JmLREJxQ0nRRUVnTQOHP1daTbNzRTK5iu5URTsvSh
+k94NmATSoxf/9avmQvXy3BCne6KylKXiO6lZahfiOZDaPu4aDUVfZXmudw0f7TaXMlmr9jvrsDu
buYwZZuyJvi2NHiXHuuB6a4y01KT0IIXYDqb7Dgoyo2+9hwYV3i87A/eQJXWnZVSfjEOcUVSyzax
f13zG/q/MvutrmZvuDJEkgDu2sNEPAY+G299dkqdBOmie75nlyJTZTo1+C29UUFnQ2778kBLD5+Y
zPyqOanZd2glatg0csPAg3RTqLh+pMWCwV3q48yj3qjKqok9hWS3iGXmjs9thQeUBW3dCWctcs7S
XLp/O3DKpF0F7mXKdtjN0Y9QaP9T5OylPJe9+9i0jwyUc9u4AV7nuuxET4bEbjW9sBStdTrkL7D1
rUr0vRBhyx1lfwGarc4HA/XsYN32fkkXXtXIiNzXlWnS7qaQPX8HY2VYRr0rL+0RtK6h80L6X4u/
fPvlKvn1aErL/nWb4Ac4iEQvQkFGHjbUN560KUYHD4HkG37MdE0ePtMWgKZCk/QLOBlh4Fmwbz6h
zsIzoDU0VwoQ3XlAiGCzH3YVbOHb1BrZd102AujAd9u9A45eQNlFX9DCSljIToXwIv/DzI7noKHg
8QC7CMdeN6rMHz/DCSKlpNbwKLBArSkWHYC6189knbgoqO0QqiVafzb2rqfVljT59EhycI8HSREB
9aC9wXdz875EAI8i4mSZQVAUDnHWueAKuWmM4ZXp0qAC6DCiYOYkZVhU0HPEEIrt35SWFBc5rcQo
UORuzm9lJEw0m9k8ZuYR7tDj7mhmEQzJ1CQLT6NPK9w++HctmzOZ5n+DnxeMA1Dcqv5Ao57bHbbl
MGR+uEZzMvfQX+NHyFy1/Xzm/QbINw0rFGPCX05SHF29TTM4r3GzgLYIGccIUe3zcZkTf0fTzyjx
BRVi67PRNCFwYKvEIWzqqO09/yKVeBWr4oWXaMdHwbyUtkPV/HH3anxAIJNMaX8uLGVLmrYm7sT7
68l3VZ6aWAE9N+ShSv9Jn9HSKHGna9WIuQ+2jBiEmvU83F9Y/GctwFXG0mVon6/7RxAwKQkyJEom
KYCTbyQAC9XjFgEO5YY+2Djvjx136OssKoJLwoUtzRzlkFi/d1A6p1MwGzUcJ8q5KF7nehsY5OpD
YmpFDWJWAaPeb0xgv4iYHCXYG6t9syzyrG36ed+xZj1G2lgiNuivNibFM0bzB0jVsyPf+18GC1lZ
arAX4y7mG0iNq6j8YX+6Tt2+mHo7ubavIK9ETUQrFBr5G3WgUkxgQDnVpdDgI6v4GhROcd5WNMl8
5dp0Mzv1IgAw1UwR7eVOIjHmDBybeBfTgtvQIxDTulG4xQtSAuU106t9HH/HHDceqDCtm14rjM4o
jhkpizGK2XiLT80TWuLNLD6ZOwATNtpYcFbuoYm/2Nl8Yq4DEelj1VSlUOJDL0HjGqXZ6DvRYdLn
d4+YpY42pyaKrPaxlE8S2sF6wyAWLAAD7taG46tvsXCYZnyAxtG+N7Tr1uN/fotnTwqkFEzh91G6
wHsUlC7mx27FA1O98Yq2NJs33WRulQr16XfyD+UUIcvJphc81BrwPTEvJbeQR/4khYZroT6l7eQW
CIb1KROS2V3E0n3ho/0XPt+XHn9nuH6/R71J0YDBtn/A7+dGzV1rwPsiM9g/v9lDC5U/WEeLJMen
E18QYA8XtbhAXwHJgHUmviEaknyJDSjSoWAhjEV5Req7lVB0Is4xT7tmjAM2JEoe/MQ7phMFOmBt
Wwk9wY01OSH1MdtkTZGuQVv3P6gFjrnkhdJTotjyWCBxiMp4Mb4DWXI9ztR99VF7yncfdx6Lv7dY
lZpEbb+yNgpyQlHF8VmLPIEAyHjGnnVoI2GLvERzvDrgN2hdqT5B1J2djBMt+nWUVWr0VDVAaGxD
Zf8jBH3zMJ/D4lS7o4SuaNJVG9d2STQngukHhE8C1WHrGkCQbjh4vYNKbQF8K1AB1Qk0CowpNRyP
PZwmUAGnNO01LRR7hwwCHmzEzZmBJcpK79Vw/CqB0q4qrJdc8iFmc4qaxEaexwRuSPKjbTNJhyTw
B9UYveidrNPfRZHarWvDMfUt/l1y9hLQulnh4mPZCle+btPay9etty6vfI0Qg/Bxt52B43c532Gc
g/uAiVGvnvnjJggRUhM7D2iA1heI6q9We5Tyy8rSPtnQ+YA6HXVIKaP9oY9yaqhZVGT17DbHd9N/
28o9XG4O2jrTsQuW4+HReA/GgBLZUr4ak+LVL+mJ5QH3apJ0jyNZJiS5L+xdahpOKk3ZXcpf71A/
lZPrlmuMUO2VxxfxmlYy8qbH+gPUX2Odb3RMyxGhksC0kWPJIOZITYHU9ZBTleI2w+zFybV+EuVS
A9lSCz1kQH3vQvsMKncUFOZrYx0o341piSgecQovRteX4TFhmHTEXo4izRDMrx6MrSXLHfoGXK5x
r6SaoQZXsJhuMv7QOgR4YpWvkqi605aAKv8v59LB3iPOP+ddE4r98gF51h+azBoFED6vJdQ+cCpc
cDvJVepSovcx704o0YXwGWt9JAE2o/tV5w8uh5Ci+N9w1UWL38YKs5eLyn4s5iBKJMUBt9G8P3jW
x1jzRHYsleoKB6496CRE0V3YETfhh3pZqz0wllDUtEQ20TEtp9Y/MYYVXh1Z4kZMHZ9okS6L3od4
F4Y/G5rn+7QgdTNHW78eHPaUgS6UBBfm4tLgi2xhOK0mWbXO+TAKJQ7K9/pqcltbr5kjNy8TVdh6
EbAErVRdLmmwZneHoGetQaTtuBdtPm8HQVKHxp7OsnvqZF417v8X4D/fhCk7yw7AhRL79zl/NtEb
Qji9W/xt75FeS8koOCrL66M31nEppaYADRxmc2VXI5to38uW2AmGQrhCMFMT8nIbZCnpnbpeSkWA
wfAko9eh5aKx4xKCKhKHP1TubU0ymNjQBZE0CY/30/wCzVcLdkmoAUbOKKYd6tkgqI546RAzF2h3
cDEoGXSNzIX6YpO95JMjP4+ReRRd8SpEr++4fftAY+13Bz2BO760xwFWfGH92Ad4L0O11ZNMhHWz
NtXRs/ksmiWhxgpUyEHK6RlujHTg0sHg463QK9ymfNkZvd3TzO3hKfTOBdAXmifSWL2q7lMxzjT4
iUNm9rjHybVKJBdQqqw6AI346mpUeJNuvMmWZ7OvsDRZQNrZOT4xQ+wOGUGnETvnmIoK3AdJcUYO
ZxIQvRkDz+31zsT7kmnaWiG4LVy1xwudYQJwY/t8Tk5J7VMraCpPqIWusxq3hNiUZPGW/t4zzaei
p1/YOY77Td6mSLD2pqVhsXk+IqFIq1RyxfCm1kZOFVqaU5kuM72b3ewsOOV4XY9NrwK6yNonHsZ8
v/WJSGOa1VJwqrlQ3MaDg9arVzskyWiSjU+CN/ottIMFSM/TiV4dZRUF/CXpIKCpyJC2QfE8X/oJ
nUTw7bkJ0fJgNy657gv6Hy4WvuP/hixVdM5O87y4RgPLf77IrUx2PaIbzshaKKo4BT9AEYLBqSGX
7G6yoc+n/td9s9M3hNctvuvjswOQ4oxNrks1ea4gu5iR4UtVkmQiI/Ywn4Z8LQ1qmxuNoPGEWQoH
fpnArdHo7VGr4JeDGK0T+yS8BbY5GM9MnreXErG6sMVIaBG5ujgKDu7gP0ZrDhRyu+g8tqjxDBa5
gT64VO/TI3HqWzAhQ2itpK6WY4vsCENKm/eJThSwkOeddRuWgVpD9JzjCu0tCW9zbCt2GSFk0mTg
dIYI9xRCpQ3JVUMfwwJASdQkKt/lNPVwj2rOBure/XDwPRpExW7MKqG/A/WqmuhI32SveJlioZ4n
ONl3QI8EXG1m66G8rW+6XsBwTGMcmmkwJOi/Ma1GzchMmikqx9P/cnCTgDi8fqJ5MAzjYeCSbQ6X
SZFyILNqzJ2xh+pp/tv7Zn0v5iyW0vr4PjJbMXzmeEG1AFv67FRu5FmvJ8pyxCJFeJBSENlycorm
G9bxzotYfUl6aOINuwnmif0uZh4RHxZeCqHMViraLb99u6Xoff+XG386cVQghkKY9UMfnrP/GNMB
7COGXJF2+e0c5U+tnk9ofcvvke6MgSTpjhWD7dnQUaUuCuP6Zw+t+y87XAPpAVBWy7KAo+0LpYGz
oF8TnlXCFBxaSHDViQUwmlcN8ctx9qucArZ8Tiq9lXQHyu0OIMEENrQcQ/2oTQWK8PMLaosg3/Y6
Ipb1IxUZmZHt23KegYsymWJYQNsfGyl8CxcfFXieX/xZ1KN9HoJT/Yt7kpWHIxfBPHHZiYZz6twO
QT+cxIqXKKNujxrSwDP/SqRoY5oW1DQMujE+VSm4wFxmhNtWCtTvZ3RMfEbc7Jf35hGNCBrNsrsm
xyPGugWOpC9z/TNc2G/mF9G8wcLYQP/WMF1qMY193EpXvjYblLevjTeLpWUp9CnHofwlK4J+xiZr
JRvCjGRdPZAmL9Zpu2nHCh1UlXpjUFf+P5K55B1v2OMHz+nW51jo/lxHmqUn1MrxE4DrBXc+xfth
Nixd5q+qkQX6yPlppMehdOPftkzHgSS83ZJzs1ftjIpMi9mj8dKy2JlgzRwq4GDFcGJ8aWUsg1p6
f/pvbTNLIN+0ES+r3DZ2cOJyuctpOpZbv/iRbnDJBNGMGZyCW5SPKoH7b+F+fgG4sZbyvVYka5ti
1tlQZqsNu8jtSOTnCayovlLG/nGKJqn2e+VT8WYp/I6uBzh4lPSXgJwZMfWxCtMc6wh72PsSjhQe
lz4K7Oy4Curwdj+h4XgjJqFJMKuVpBceJRLOXD7WIzEJPsJmfnX3eqhNKJ4tSDSRNVw2UCUYukHi
k8kZU/huMIUg6VQkgy54WTQboS2UtBt/lIq1aB/ZaK2e/WKszD/Bi519UkFijrKkxPtAR2w20G7f
M3nw3vHQbpVfC80WpBsCE6PUT053oyGJz7zFENk7PAeSZoVSvVDe4ty6FQw6qQwsYljidMo14Ahj
sBUIL1fj11YLFYqhOLHuK17zmxq7KK2GadN7YPFQ0W5Er9xlHZ2cv1Xf9fmfR/Xi1dYVc01S/wgA
l6oHDcffQRjoM/5hGUJy4MmFNgvlBGA2sQ7ZtpM7JuPcYQj5ZUPMRSjPnFb4CN9O22ERK3rikeeJ
t0TxOZld4vVjPqp3Ak8OT3ULeH3vwN9mGx7VDkPjpXNTAwdWIh/IyjHYV8It45LJm6E/yWI8CVxj
HZaHXvwFNJbYo/A077DRHRd45gyZ6VSW8RS+iXV5kbE1PPMKW0hwoAaiKcc80PdmkvgDIMPg5m6M
hTT/M0E0kD+X6QsF2Owv1PsPNOpCDhQ89jaTku3QfdZmxbG8b+XKgp0hnbMpW2gtoI1WRZFi2fEn
TPuR9G23OstgpG28vrLWkqjpwx6NKsPUTmxH83nt68lHhxCJB2QYXOKqnwAl/J7UXi8869dM4yD3
BK8KtxaoA9/A9VnQinQjj5o5ut1i7uDqsfqHPVYgxcUW6NVVrkZy0EcJgLoWWlYDSFVAxZ9+CEJN
l3PX5B6QDL7W0tc2d0V/MwP1Gq1JHzLoZ50CnNwlViyr5HEBjxGw9E4cBv2cw1D4hBhJ9E6BAn2I
dqadpzDlxVRvviXU24mvgUNSo1YYuSdLaxogh/Z/yRaMssP9B7MnMqqX1EuPeLdmdbotJ6w7OQwy
+J4k2tXZxWYBL4YZVaA1LLGrBwjm4jG+iE9PXHbg/q7O1SZ9MGnKRm2MM+UGr0/i2MrKRvst1Wj+
YR31F17A/ygNoOpjyV8r2XdBqlrANpQYEETNeQqprUgyRPSEp16fFTtkiHLlewHHDlR7hXtuUKNN
b4eS1JJTDd4mKb65ednbhN5m9llS34IckUrSr9sgidElfnNIYgGRbI/1p1rx/VALbwKvzZMsBcC0
ErUIVcewbqHTc4Fe8aaqxD9ZaejjLQ3ADLeXSmSS33fW5v+oIkHB4nhOzgU9Kxec4hvuRIRs67q5
1JtP5urUlkfYEeagQiD9N9yhjOP9ECwSVpWwQERXUsmDjjYRLjmcUTlc03J068GvIBZZfvewsMOb
eXoVZR/D8pyRsaGMVzycbzbLfJTssvpNgmB3CTqOxQsCHD8moXSXGmDYXrMFUP0AjmufVvu6Zm0j
ZmsOn64p2PsF6ChX4abNQ23t+T/Pvv94W4UDxgLUtUoeCajWwRpcQSbHFZlMFJ8jYzdDGt2GNPSh
bjJFx5FfmThhdUYQ/143hqdjug5bhEME7THbxWNcyiBypoaO2phgn9b/gHuWX8GLsGb6+UYmxkiH
OVXgii7vMNlMW31HXOnN4uF3GQ6e7SQozCvErssfnDUXORO9tivhgCthWjgjJtwEqklegq4m/emD
BcDcs2h8NZrOk1iOtU/O55FvfPNJq5PrLxK5yQHkovbZSBwXAx7v+X+d8afGAOkXPhooh4rB3fg3
5Ksqotgg1kugvd0ptjoqzgwqq0C9s5bJo1vKyE/7alVjZPm/eYWX+6yCShcxj2WObJhtb7c/G/cP
VPl0S6Lyr0CfR9p8dX8u0PfP8OyDTHbli2r7PJiV4x6ppmqbcjw3hnaAe0LHxsbhFLfYgfY2SRZf
7mbbYFt0QSI1WKQYLIToYuw77Zn8U7hGsH8zolzkSY7ducFALC3/gFvpV31If2MPKaNOEvGTwvuD
VZbrBO5sNnN9IewsUn7CsJhyKjznYznUWV5uX4iDuv1bfK+cLTTzPYFCcYaCyqF8vxDDShX+CuBn
qsLaxhdrLTtRBXQHfl+Nx1/x4a/zwthC8ma0dBGyznhirkCPizOaCWAYUXxqZzg+0wWjfxKdEP+g
NKU8EvhY68qqUNQYch/8pgrTdQFT1m9K9aecB5/+VTFQvwYMLtA7Oq7TDVI7sZEt97qSDIYeOnmT
GTsjfjcqnGfX2eQdc1KLb0YbPcBH5PYhR576D5jAIIuw0lPRSfq2BjxTQcU0lLrEm0wYXkS/gGbH
n6KAzZVA3Qrp2GBtyHVUk/jaGUb1dGxtg7MNLZ9i8s0ye4DVgU5yYbvxeW+TtVfZEiO6tN/wySjP
pBzCDAkJ22/aKgAPEIUU4ul4Ot9VLNtynTWqt/mrVcMJ+HYi2ASv7OeayJV99fou+xiLRbZSS2w8
EWsNu2PiwY03S9le/lprix9ljJxV8cvvYtnvaDhqg4pp6UEfw9TUjD10UjBRuWuqcsa4CWvHTjiv
nOa8MVVJNKAPAg+KMCeTZyKVOkgzvYbPwG1nFD9sN83NuVgl/Nr+ouYjUBJqjvSBrgKSTcIp8pc4
8oLIxe8By/YOlq/aB9ZwsrolzTNXRrSs0ZJQdWs3qStlXSFYuihBVBr65XrRz/dqaFPDJyofFY1/
DLEbJj4DEz75Dxy45w/Kj0PzNypStSjaWRZkMAehz3gotHaiZ8AFdN0U/QtHMJCZpmPwlb2jOgOd
5QZOw+7CPhp+bmaxHXFLTTeFBiRAejIzwIUhDr9IcQs6vGg7MBn3wlOpkLw/hlDsm5zu0aKyEw+t
JVZMmHnTcv7sC51f3qbMRO+mKxFzqVfw4th61/V0c7NpLG1j4LxhK0Nm9WgiMkh/iXcOhFnK2SwX
S8JJ8CH445vvJ9lWvi9h2EHPn/GPA2FZOZj8IiCtlQz6v+vHXntI9/YPC1NTWh5BCrBiRplfPaVV
h1BB5QiZakbAkrPtXbJ8d2+cUnEnE1rSrCjvDY44MvoAOt3MvdMWGTRbdKYY+iHcXjwNxIrMejns
UUJhbVHtWTV6ShRizVgy+eCLjb2XOWWsl57zZ/drH4RN9rE4viNFzYfa+soUQWe6wYbJFprbpWT9
AISGYvqeil4LAxvT2E9ue+21EhqCKYBMtjLmRKrfv6TTf61KYNheJehrpzhyqmQU16RqSTYS7LbC
7YxESsgXUrACubCT9+6sVmIQD1OuaYfOSruJfFkCg4c5a1kuwDNjTO3z4eDBrtnwZHjwgT/XG0tL
pIkyUn1vYFW6szGLMTpPlOc4Csww3x753yfPFFnwaIxkB8oqFhWPaI9hVtnMrSZNW5FzFNV2F6jm
hxPipndrFINTb8FZCDEnsxHEHj1hk3oykvePrfUJ6D8c6Fpe3xKI18w/HOKQBa20amJEFgQw9k5D
F96WjT2KupaJDNVrH8JdAfKEXAwO2FSe65jQaiKau+xeC8PBQX0FFTtiLOA4xRUPPfuoiU+bbZXf
RSieam1j3svR0zRLb9JY0H5kCkw7xFuSRKGLcoIno6gW81NhbMKWSTuosqb+7YsVkDeb9vQLnNh1
lJ3JDteH852OKChlhIUCvDp/Azh0D0IoScwtPLO/q9Jl5rX7tSSf0vaoILld+tFudEUjpAKb1XsX
rzEVCJZSCdp+huVAITjbBoDrjhHGoO4MnqrXxpP47jwvszdJoHtuEoOB7B+f6EZtJHRqMg40oAYu
qfwGXkSYwSQt6tU3TLcGq/y1aEkqivbyKzjJRnOE9gVvIzo/8l2JATZF9iEphylVeNj+jAx9xGLw
87rfkfbBIJFEEjvfz3VMluaIP7zzyeRaCm++/Wl26PEqPulmnwLePUvIA8c/xpVeS9VUl9PQgucn
Tm6OKgPnrHzHFHpcFrEBYVlJp8SXd/IoLSjGBaLt3AY93dazWVNSjgWX6twPdbc80OY+lX0VUdaa
zvGPkLC+3w4R1qbq4mBh+c6BlhFVeXNWEzulqzRCIsOW7yCWlAUQo1KV/MxydAQQwieuNhqex67b
43Zb6nZX1y1RHvN12GovlVac5Y+XwW738v4oI5jbbj1gPqasatBm2gx8KTYcnYMI1aRtf+XrkUfR
pGivT8nfpvswqWl9HAO+ErF07H8r60bUaugLCJapTsDbq+F5MQgTDAiS+iGB2QTMrJbo+r3RqDeV
rAJ8s67148CuYhHqvvtA3WivSvfxJfhQKZ4hzw7pTsEz11r2H18m0QpUU+2tniTFSdJu7QWvN10c
bHGB+0KtoUFXnr6W4gAwaIdm5chcoY2/VLivJSjlcn5iF6s2SfbrQBR7BOzvtzyc8YsfonMfwSgc
6FIu4wXk3MbycOfOPYPnX1CH0WD12fthnmukbhCLGYV8KGlsZ0uJ45T5f+rMHLPjfVdbJv4HGhS3
H2Iuto0absA/NJIgl/IbBJaDgRYyh10cywYfZSo/eY6WCs1ot0nTh5w2Ev4ZVVo/H83QkQVrHlM2
pJXgUd3AHabZY7iFrtpRieBTwK5ZvemPoFoims5TKfiWJWUA3GDBTXofeBrxHmBOwImXhHN/CSTA
ZSfcBJ21R1IOHaINVBdBb+RByuWQf+VvVvCwLLdos0sarxF6Q3L+NUOaY/FXjPqsIC9iOYLW0ijo
S0kbmL6Ybvz4vwX8C0FjhFnbBj0rqjJfMcsDqgbCJsPC+BopzlNh6B77JxolbVMNhhuCO4ZG60Zv
Har3Bcn6C4ZZQ5MJBy0GOlOYsEWrIMtAkClqwqW5ZcUet375P82El8Il+Im/98Hwb0CwqFp9oQ92
hQw9jz9SyiPoBpITRwDAs5U39A30paJvaz5iQWsFCHx79dxkcXo0W1TPT/5xHsA5y50YwkyIohdp
0fMT+MraIUk2ehzHFJDwkZ/0Ahfyc+npulrFmIxBCvF6aNVOJWhGLBtg48X4SNIns77LzaN74JMG
b4nRAvt8pqTiVzip6ppWJXc3kn5oCFI8DTGvIrXE7goaLHWHMxZWJkNSCMEzl/vmDAAZ1IsPCdKx
DZA3t9R3uRkBmFaUdE3dcR0GbNHDuGXivsRwQ47dxZJqEK8XXX8vdkVwLsBohoFdx7iReu22aU8R
rI+wN4Aud5AryjcyrfTWm/hcBJoI3kZ29IdginKSacNNSYArAiM9S29cMr0TF1JL9keo6ZMjp3je
2SH1iv+TmXet1Fkdl4f/pcxgZDuIUs1OTHIORDO+zp+R0MZ0nzFBXnnwdB8XHabPpaxmZECYEY3k
lAIkr3XyZQXmMd8Pp0pz/J5dKuI7O8v2Xa5dTmtP49Aptd9XeoxA5qWV3AO/Amt36yj8CQ4jJmwB
1UesVWHDPkphbrCzets8ZD230KJ4Li76fXO+QxnAE6zr1MQVqoELpgADJW23Du2VbR56V24Lo7ak
NowoR+ctcW5O8paP7ESn7VQqb0Fhk2B4OnokVFssoVVesRIqlaTMrCg/7hEsuLr7qqhJlmPgxcB9
4yEQiDWphCP5hWydH6itVkGHrJ0s5hlTYivjY3CxXC4P0p+3PHk5NX0moNbnYhxjwp+pmuV8iU2F
wvijfqdQPd515iNh79Pd5cy5h1Li1LQY9RzHeBseFYq5a+0JOnG8YPwXStQJUX+nIUTvqGyUyoc9
RSo530EdWRGHTI4A/Lf1kcQ7n+MUUI6sbcTKcMAk3FWVBI7mUPX2a8G9IGZD6gcPL3f73mp16td3
EvDh1rAyBFQy130ofixn5Ni7P9yYVPxxx++ZsIsWUeY65KEFB4bmDJwrnEtZvf3x8CCwT4siaOdu
TJUbzHN6p6phW3eFqj8GWXInNRJgAJT6KkjOjemNUS3bOlM4FTUr2FZC4/QWJvt9GBEmP2Kenzpg
0eT+moN8p3s1xovXsKW7jZDUDPCzjp+41FiriLlV8Aah6oaQuMwaVNog2c66nHEdpP46U+inr5Ky
9ToXjcpopJTc65fS7FUZt9wJBu+jT0VhXMm0OE7gBJ53MJ5ZEDGMj+Jo6Vy9TMCqxrzWJiZKVpr+
j/J605Ejab8cUQPbDNv9xN97yjUvrbUcbgQYogIivvVPDw5OO87wN28BXgXgNRhSJLurkOZtXs5t
eTitrGeJmMhPvrLGIn/SqpGsPJBKdI3QtZz0pD3O7XmTWhLJRR/dOdls1tkGw0ZnUsJLK1YiBxOj
38ez5xHrshmEed9s39H8+PSFfdNn8/VhcJvrz4cWFbcQr9jhWn7TDQC9aWhkP8NPYwzM9PWKyWKf
XyFwFPSCmvwL+0VWWMvs9HsZB2JV8o+eVdVlAD7k3WZ9q/0TQHjigDLcZrlgLhCmXUlcjn7pAjT/
5WPB4kPNOiAHwKP8+pgPyl+RwCWPdTD5x6j87cIDud8Cn3/sUNM3ioH9Eoa35jqbWTu0NIqGxHKt
BYSKYCi2vFnZL1pblnQuqShDvww+Md4ybhkcDcLzOcdzDDzfsb0wPkjc5eNtilHBQ77uv7QHImV/
Td4Nu5UeOhubNa3zdiHajAyqO+7+F4m+pjVu6F9eopjkvhI6Y9rXJPC4UVA6FKZBGfb0OQK0foMH
WZXZyxFk/TQbevxgvash1sfeO4sCdLzzP4iKlA6mKa6SCCa9Y/n4QmdnNEoeVVcWqbxFHA/juMBr
sL7zzwcXtSv1Z8Gn1WoHOaqmA7rRRA1F+/o258MUz+nen48kzez48KATy+MgEww0tJqbk6SKg1Lc
of8H8w32K4UW/xnbmHr2aXCxMlkvwpfeZUXMNazSXhKc/FMF+DJTVqakgU+XRqiByAqpLotZatGn
RDKGtk6EjL/2xuCVUjl0aKY03MZLFGk/4FqVJGUoEVWJf5KCL3pMiDAF8p+SfsdJysDKUkP0w8/+
H9N3YDqmDcj9s0RZeta2Gx1+35OORQju9Muxguvg2Vef+XqzTcKpt8vuBT/ihL51us2uJat3cGax
vAmNL8RoZpmped225ADumdaNYDZFAWCFTOp3u9NvSow3xvCMtYmKX/1maScVoiLbL2jWGiW0C0Cc
P0+4F5TXW/O1WaF8bLhMajGJ0oZOX25l6XYgwyT4IRCg1CdXarhxOp+wpp/n+6IagqlLw4crFH/B
DzAnXAA6gDU7B550B9OBcoduj7vQTsB3Nx3ODRfcHVNFGO9lWR5q6tjrL5sDM0OK4QjdS7/LXsc1
FEl+5+muV1C0sxUXrlpC4jxtGuzdLO4mNMBTcLl3KL2WEHHCfKNwKVt3cunRgbwP5VczIaGFIKzL
H/UHid9RBT9fmX2dJIWcAvplexCOS82r8FjUhky0NgnwJgSmg4CpmMY2ivOtGm+4l59etePxUpTb
1E6s27P+/B0ibkG3LKCoN8th4KPm5eGYvYy2zPVucNizOFwc1rIvS/81BRt2G0vCeLNbQ0zAVbLk
rtW1M/gX9AsWGZpAwm2U5njUP1VE4tHsSSs8xeFYQYjk3nOYf9enJZE3RiPnGmYyJl5aEjcEA2j6
rGAUcFYrgL7K5qzfue+Seu1RfOW/b4VETApP2+W9dsrTXzEmrUH8NeyHB7lUE5r/ghf8UB5o45g3
903qgD5v1HtjMVaeV8aQwij5HaEXWkg2JbwzXT5J8h6ObAjLywxmIpGCFEzik1DPL+R4hbADyR4t
EDS/C6QG26WzEwnDpA+JrQK1yH7wt0b3auwNMVHBtoIxvW68MnCEtYiKiHAPxekSelTpbJQN/zCt
djk9cstdV6osOAQkjQ4501Bdva0lVGvoLv8u1SLFqLBokCTcZSGKhk/Kl2rQAV6XKTpjCxGNQAUA
5uGT3/SMVbAVTDO5OTkbAVOZaymqboiU/oEpzX2tlIEYCtMSBkmMaPX30zCPKOm4IINdOunXW5KG
wfHnW67XbJDHgcoJKsmNUcEHrZOxQ+l0+MvRKOJTa+klHwZ+y4BPw81zpKlYDJbm0P4d0u7w/lDI
fwkGk4A6J69roCyGTEGanff0MsjEzju8gQl8kc8Q1haYwZa1eKJhO2V14E6TW4zjtcg4AiqJHMZ2
cyVJ/BZLgrTYrgzM7Mqy7pnSQjsCLvOK1HE35Ul08y7+c0IneyFbjlj7BBk/CP07CUV13mA0cIgs
cUwk3lKxvUTAAyPNmiJ2jzs3wbxrF5eL8GndtVVzTF5nnOmMfWvZM/gQ1Bt2ECOeoJmI7zjlnD+Y
qrEK1U3eGZ+poRZKbpkswNZgjd5hLjaTUILZPUtWcICnTwSZbH8BdLFyzNtUnOpkuloxOYQHEOOP
wNPiG89K1BcN2IlVC8sq/No7anOklhmZ8MW8/nQKYleBf2vCgTZu7Thk4qXFwOm3z3UVoWi3DFMH
9RgSah+iqEcrRAPPPjUYZVtyGH97uGRIDZBwBmWjrU+4vP6eTZqeAd4i/CH8MFt6SxHfTXHIwhUp
+fCTTWUuDl/kLrmOnocK7+obERqMQnEPguZHQQtU/jMk4Lt7ZMEHHXUuviaqnQn3U4EVcAKPzCq+
AeFYL5be/mJNMb8eJQv3UgTHRRfduz2kqLcrDndw+uxlqPWAA0TWCw0oArC6cgoAoysW7ikBMXX+
gCS40x2Bj/wXIXSXFiTLJcUt7PR2wH/VhT2LWUymBrbKCLpzUQlEdFIEr0Ci/oYNQvUb8Ne5HdbJ
GMrNjd+ze1XyJXKa7le56cgtaj2JPI5IK+uoo5+WzY1ndRwnNvMdpEpWfSxwhml5nNjKeIo8fg4r
PokaM03PY/D3t4E2bQzLHMKjfHx+dh6Q+cofxgB1qWZi5KjoYCRQaFg9TL1iLcgKv+CIJdAUVnQA
gPsWm92VoATTLSDpPggQ6/1H8aP3ijNn003k2DWV8Ybcc4YfxvcZ8vRBtJAU9lpRfBHa+NfCELRf
4KWW2VwwObBXhA1KSqx8/kcjeTWRrq1eR6WK+CdOxLQyOSBc4Zz6KDfxcEFL1vFZcxp0x/ZosT6j
Fr1nMBRuVdA5013a8WAjJOE0bOZzWaHLxaGtq9thOElnATWp/f0OpON2B0HdtRwM5YcjNJcOhTbu
qp8QNbdr7BQ3W0csBLwEPQYlwFaLUXNaHUHMYvoI8bcHjzILHB20bpdPFMPQ0MN6uazxVUO179xJ
Se0SnH2YpcdgMEoRB4hcTGjFsCUbDOQWbqRHAV0GFBPpryS0uWhBWrh0gneJr++Bstc1fT4JkZfg
4g9hJoXhtfDwV5FKpvo0UfvWa9pHb4EM/KAX9kny3zxqS2Hh9WPhZHUm6E6wNx3TbvSGPyygoDnX
ZLONVK86MRSICGqseEQa4VgbrfUKayHrKF8YZ0qW5PlQfksmQHF6Bp+DH3gX4UbCzSUDfbIPc+S/
C3FZ7osjYYCW5ZlKJ1rKgh9eRb/vBdolDRAhqxkSgP0UN9F/PIUMXvcd+Pdo7falARsEDHozQwNb
3N/1x6pWf+29P6tBTHBJGcss0D6HNCJedcqvvJcVt0alSfKbaDJVwF9x86zgSdtMO2dHw0/vFmlo
U/xejJgq9+KYKRP1lUillpSsQCHbY96Kqokjwbx7gnh16PpomMxEoWiH4PxheJvQCY6wgAqzWUPf
OWH4hb0lMHlUE6UnIie/PCn0x4RQIDBUwh896mVEB57F1niqQQsF4l3n0pK4dBhimAHj92p5lSnV
GG73O64WY8mRqF673MBdJqStfFFeAA/FxmWFxQ2HX53ytXtMEhmAO9A6nDzvVNuLM6C5ku4yGo3Z
xFw35TP++cOWyYrmKJ8Y0eSJc9riVVrXNikccAGD9ZFgNymnc3SRWBZXkUmnwC6MnntpV+D7jzZD
F7Rc+pTz8oB5udFXHex44eZ9mmCN9O7v4uDcVZf9+mwoLVnZ3oazLKf4EH/1S8486zcS7F/ms1vJ
+9HoFHA4szwJciQRV4EuWII093gCwN0yWxu0yjpzENJLrs5X4lY0gV9ejQsjJYVuEZO/WF11BwVI
vlHHeFjB3elxYJj3UNlplPVuLRps9eikmz6QnMjOOJT9o6AlRtcS30XE4V9q8AOhAAPxngeAKZ5F
zpkb2T1xOIEiUcuOACyy8+pMxJpy1K/RwQy0RsEg1ypM2hi6x0QJ7WNIv6sE/iwlv3rRjFDFK2Ki
B95bzTI2V/7LTLAfa9yaSdntHZvd8Fw42hYq6VgtKLGtOpuvXfijrD9x3jKaW+o7X8YZieLoRIGM
EEsc5q4OSzDSwuuLvZBsL2tDW1y62LjS/JgUQeMj8yXhDkFAcons0uF8zbL1C9l9mpEzlRYfDVVY
4U25NTKIH+IcC68rCZNTk6Eu/iEDk6OmY8Enf0dzJCkbEeQU6L2PwQ/GuPijMeCenjKL2jC8Ad3R
HJFds/o9z7Z2b2Xm3QInfq5PJCkh7e0Vv/wAj9D75BX4OeFia5ZOI9z05SK8pWpShy1BhUBHLFSz
ETVIvWGtrLBJArCdfSmEpfib8K9gxut4eapYn9PNC3PZGrNVFVR2T1KxwMkThaaaf8t7XoiRXOj/
AUnZ8wKr3Fwzb2G1FaQNdwTid22ph6Fm6aO+yNs+7vGLATMjCRJyPcIEEPlvoXBna4vU+7V9qf/F
UPmHhpyiqPTwWAixuqBkCOtmtAtiavZm3oMVysFlSLajHEopSEqQDL+TP1SKmMZGdc/qts/6CaIu
vC8TsrU5TFb+FKZJm4i+ERuS+WPK0raREuJJwKVPbTMERrXhnPtidGkkwhvLC1GWuDl1qpITN7no
X2SOdYinxrErTVOcRlQmBzqYK7EMCWhW0N9Gd13gC+SXDYwZ3T9E3oIZNv/72Kl7rKixtNkTXotp
TxWekottH13cm6CDUDCOga6xoLLAvqKyDdtpAv/jrTIx8BIW+nOqeHF1Ekkk4+WepHpalhUbrPGN
7sjBbsCzTkO8UZ38J9zNDrTEcmxZ1mhfWbTu2+iMp5HT861elHjZDlqAz9ApOVaAgB4hiC3fQGHb
je/pVrqR4wSD+JJaGU8H4w/VbuMN2xduFQGp+nM0WKnYk4gE5wgsrxqalOdXAXHOh6QSqWV6fuGD
UvJ1tUkR/RMKlQXGsttzQgucIztQac8rhcOLhXveXBX0wWPxbdvoCAtYkHy/L2R0dg5IPNsdFPy2
uBeWiKO9GE09SumA/zBn2+yRqaLrV/dcHiZbcJbSayliSQESA8Oxgu0sgKxvtRf7qgxhtYb1md7G
/bfskIaCOlMIwKDmszMA0qC2UUaUTFPkbtfyK0Ietf9ntKrq6yf/mnup+XmbcADPVdPpMVMW8COe
dMHEkD8CwZVuc0ioBvfD471hyDD5CwnRaGbtCgc/H2alVkbaVVPa6K01D7acvmafcHGNfLdJ76z6
JpqSbLZ0yGLHXqTKaXRsqSbsV2kp4+8JWYFwd6NG9IKwbfO3Ee1BBjsjFRef0ZhZXWELCM4B6MEm
sJXaHmra1uW5dczxB29Zex/Uf5Bi+5WlMvlUphNye/aOFXy65BjeZy3gFSIfbquUjStbGvrQORT8
vWpgqwcG9BXmXlH0dUq9kVxj1dHJRSwzqnqT83lQUboGm86Q0+kj8zcuvtk/dB1CDMoPs5AjP5oZ
b52o1p5f20XUr/70ClF6/pBzOYqmZhEBWbtu+5KE/TUDPF4pxjrOKa8B+AxWLJDmdKNZoE/1uPGc
oZANrvutTUqLlR0KMiC2PSxI+M3mAleCH0XZGMZRRjI3urEBP3IPANUZ6e8SVJH1Pajbz0rOQ16b
3EX5kuOhkJSsfuXeE17w6KLVECKxWgpsZRs7QCRPUfIZPKFtECZ2KlMFd/nOliTH1x9xPvCVzFhB
tfI3+zeEG0U20dW4rZ4daQk9fEtMXRvvGz9kU5yvVxbIGWYl2aqvv3Wgjv4vpok0dVL0i6jbOkV7
pIVVRpSKa7qfN9r2K36nSaLRYKRJkBCCM3WeLqCcqrlgynMmAMHB3p3xsmj9mZ5GY/4BEtrm7p5O
ngPCu4lV4X6MFQuqLtOjq5bt8PqJq5q3xbslfPT03S2eVphW5VGXUy+jAFzTnLnu67FJqx9kouMJ
N3EwdhD3SAmc+m/7BT7fmAdYN05GDHAg8WbFstU/JuhUInSg4dgNxvv77wfJb2WRNU9phXh+q8OF
E6ETAwhOaJ1FBJ1SSS/xDOswBlyOgLKZglKdiZdQ8njRl0/h2WHncrV6//UXnQqAyTkLT21vEMhh
Yg6Jcvyscx1vwSOiuQT2u0ziaeT5syZaJW2QtYJ99PSSU2DI9AjlpEshIaqsixQU62GAs/SS6Byl
iI+RJpNOwqxcHZaoMSzd9bWzKvG21sn0c7k5FDRmuiks4MJoqiyinjADPV2OyIfi+zjZuNxw65hj
5k65ea6IltLnfUCtqVgnWyoKxGhsnH3k5LqiBIL34VCFOXqT9ZG/2Ol9pVwiEDcTbO+IrvfmoHJQ
AgppFT85zoGbRknn/GjIwu6y7+zwmcHmTGowzeOwkDc5csZODFHfRts6JgIEvCVyXaL1f6l0LtOL
Q4layeJVzeErqFRgkvjKNu8SQO4A7CfMiDBy9pdKZavzfo9DVJvk6FoyMwc5DDtjH5v/oH964Q1s
hP6aG4vC8QSZJgX7heGbE9J7EeWGgrrwVrsKjuNx3nd6Tdvtd52mxQ5iRHxGFfO2dv+b/WS8g8Fu
1jccH8iRaxTC/owSk0/cxRo/3XkjpzI2oAchykaqfCYpIsN6hckTDl++IhMNCXjStR6qKzFH9Mbu
PDh8tB7uAT3uGrkDiS7gi8uY+ArpVm96+ZHigGEn85TwIbfsoCG0pU5V3CNZJyAmovxidYab/hTV
3DH6pp2RCgkh1AMPfBnQlDjH6KwTPZa1c4isMeMBq/sgw1y11jWfcMSEUoNCLCxrUoCfW2cy0kcN
OfSEVi1fUT1mAlYT8Dod9SHe9/K2egNytUQ3sLohuj4jzw/vI7LmM0GpTU/LdK59Bk6KUkpUZreg
J4jv++PfHcX5YV8zO6j09ncupbLMdJb9EURPBunaSSYy2v2rrZTsidDo2Dn0F8C1vTbwhLEwLhx2
9Z3K3jIEd/GXLy6EKOjS0f2y6KxLUKjHJjiDG6f20PbTOjMCKMv8/MSw4VDcxBmQ0casUwewLoAB
jtOHwoaQdwcj3K8sqx/SuSx4ylGyRLrNU+MxU2etev+sfh9EuCyxt1wzBnY7Qf9XuN21VDZEcw3T
zz7VYNCt4WCzISG5R/l/tCPKma0GAdUXtqkBu1Iuy83tdZeZLlO++WWuO5x1NvXXkKI9s6cZAtGD
4bILWU7d33f4mRDBnOC+uPFnRhMbZL7GxTOfnef0BPjNAKS5GLdMTulx8U6he1pfspmuU4cYi8NL
RcbVE0qwTgAjtnDxKjt2TL7UV65S0vMlEp59OA8MrbW8NyXmzEIyzZdDb8EeKRkLDV5VH69HrgIZ
6jQvL91ei3rxSUNJwEWRRKo3Gawpng7W+vBisQg95jg7JpY3N/LvdUHw8X0XLyOAfXqI8XTkC7z4
5GdX2ucVJzrEOuw+kIJLhUymTX3UHjUJbnhV1jlIyjLcoV8dPcKf3W1RV1VhX66zCYg0iHiWafWG
uy4/axbNfuY4CY3iwgJe1tjRbS/hyr4WfmTE9MvD6OsaY5Tx1F/RlRYtaiH8SoXd6i6P5HTHXTML
iSUJb27/jOFqZ8ZTN3WUI2j2WGBfvXncsJ3dnT7PHFKlxlqVsRNNQ20cAPpQpEEoOkuHZqR3bFu9
sNPXslbfSBh09lGvmeRlxa99rlvntycCLX10G0U6LwoWZ/oHnPMxc3+hVyKhWFboSSDA2xoSN8c7
JRelnOn/o5kJiY94Pa8syoQ5fu3b876HnPpFAJXGxfurn7gJoDnFLx8hgwD/oara5MY+cDSuOxnM
1AlmASUYffd6HdCL2rBLy2kyM1GYlBTexsTmfB2asuzu/Lwoi1zm+ZLeFNsCczmrbVN8UNK3osYW
P75e+o9lpdYfHGFx9mYmjQ5vgYocYkiW4sbq0dGxmel+Dq+lVJUbjGV3wqfdcJW1vDrbmCR2eAS9
LWAFsEETuO+toslGKOJsPdRYw4cS7EgzGAg6ZRToVvsSezO1INU7o5kCD/xR58R8xluesfo2YncQ
B+RnYol31CbiGRopAslfMKgNSX2DHhxHu5EtKS8SATeHEnRWkaTLeHZorLrLBn32wphDz4PqPEWM
tXUE92tmDq/eifFcWdVx+01HtL6a+3lju1B6kvAeWxoROJ1Ytl8700Za1Bb7vSeZiVXHAr9cwg3I
0d7PL/M1x1b4XFEFPKsPsVf6/SA6qPrEoZu1Qq9bYZGnMQYb4DIf1kP/p1a4zpjlNst2UI23GBzX
14VnxwCaHS7YerOoobIIjWdFv+oRCvPG/4+oK2s5lTNShGWObnH71Q7zIf6fRfjRMAgGstog88Jz
ypmNh1X94ita6vfXd2qfoqSMN2OC6KswIoW+04dkpHQ2VSwDn/O6q470aKXAdq5MtBR1LuJnc9xf
FWPjGORbCCTprMDxUrluNuO4ndPTItE0FYkI7GOlUn3+NlEUzUXlxbBMG97fQi4o7NePiZ+vCvT0
AjgFHOwp1qwIE89kkWOJavJvoMBlm6XU1Ffyl2tEvgqul1fw4itCRan2b3zeNF1EomshFtxQi2tL
1bsny1Q5rSYTkorPTPIuBVsxEMSkVEuys8bpHdC4rgdRU4oGnfOo6UY91PFINpAcxJoL2eCdSVyU
jAKvqvKc1qCr76qcGlsDTWZ2F9kSAafM3ELexCW+NFtJidjEIGeBvxNy6vR1qpOYYK/fF9bm0e+x
1zG3em6hXSqs4CvfHRQEWonrdJ1hlVn60fZurgMUTCmfV8OsF+rL1/4VCuycxPK5OBNm7ItglrYe
0eryiaFQRVC2sj9H59CHH9Uzgr3GSM3+IQvfoR7RsGKVIa3Hu0n1HXGVss9OFBP16CFcykdSbgPD
CuL9qeyZvJ7R0/C4KEBsaXG7woxkJ1PT2E2Af1RjZe7zHbQv0UD1oRYMDxMhFjCqslaaP18UJfiw
tnhqnh2mo6ZBV4WGIAPzVnpaqkoku7r4iN+dLVnPPrsY3dGlKQvvOCbq9gVCa06Cy9ptOc2q1LcH
CP13LNLwINcoCEtqtkaF8U1nscBbUiDWIBegrPP4CCpeDXSRK5A/3Y0NrGpaarFVnm3pch6Gr3Sj
hPyRjwHue1nYU8cAcTZcbIkhaR4GkdWyqCfPijo11HaURWBweLdOalGZnPafeIU2P/+zxIlYKdJQ
d3l1l/u9RrhBUVmSyxex0Ny6Sv5SpuTcRhKWpbC9Q2qjC/S3RDrfYbdgm2sKEhn0njDQlm5D+q1Y
w7GClApKqtNDDoMV3a6bgNgJHBMAhsc6iWM/BemKv9utTsnz8/pvMLXnYM7vYmdBIUU+HF/hVs3L
cA305adTtDmRjj9T4tW0xk4Szej8X0s4ZlB+7d1IQMmEoYj9q6JfNwDB6OSfU3lvCG9s57CuIKVQ
hb7PI51z5wbUcxsMgBOO5oDdRfrrtwQpZywMg0sxiXRXvw6YfP4Kw9ZIsD/qmx5QqhXjNfVUCEp3
w6pKVp1wnmZO7xbDk5n4M1f63hlwrghmmyyd+LBsuHeiLSqtCqzLzWhga1DaofdDUzxlD1VB5mR2
e+VZdvJvkzwhy7CR0DjevbdkvD0vnRcFOLCyweMSMCKlowheyEKrIx8C54GuFzCody07hIBuhACA
Ss2o6R/ThK6LSej+iFhoe4ieQz1FPMgZDIEoZmJXC2em4ekan7cXSQffgO9DjG0sXpr7BFcI/tme
RdKE7HKUDTVWFVMkoLWqJh/GJUwhacGKjM3MAm9xL3/zi5Fy+7LsYGyVizv8haq5tL/brycGTL9B
jEka9VGdatfpQklLMs/hff8jimq+SeaUOSLU6v9MIxt+JCwtkEwOCf6fWUchARvOnr/EgSI9N2To
K5IN2OTH/UK8GttE+6vBLnYoxdlwBom2OnBGLi/q5IIx1F2HdNloQvuOd6VgTUCQwRvAYNjYOiBF
guEtGtQZF3k42br34OpCmQEch+fec0s5lQoIDhajq3KA3B7NBaJjLPvYiT9S8/Ei+0NLPDZ7p0MI
yfA5f9meC2xopxfiRpyQ4K1rrSTxxyGivw43uOE+x0WjTkus5n0vsdha0TopWA5cjCBkiSMy35I6
k7z8BPjjHyVRqLZTvQ8WfYcyqO494qNlPF/a5y7rS7QkfEJq9fE+i604ZaV9D1KODEV5QZ6zbwlA
FzybJOTAvcwzXYQLtyKuH8KJ8iYT4c3ipNnNJtoDE5r6IFzAyMnxwSYprWir04Oxp6w5+j78Pfb0
0nwZUqLkkRx/SMVn92ijxoo5ZdmG30ZZvU1dHyxD0/OgPjU9diMi71agTi15AjPprAcLRVmBCmaI
Nw2KA7Ab7h3AANNIg9vmrgqg8bOEbthj1r7s5gvB4wmYXtIgSHxtRzBMYPpSVdK+ckWYV0iHtlxl
dMcXNwHSs8YPdKINXeZZ5bBpBqq7kBGuSVMBnKThXkqkDr3QjHJMT4U4xqSeOh/nq5At7789goOl
MiNUOhCceR0xLsWlzWxzFKGyzakGFYQj7kPgodWeTKavodpoOLiRtcDfsQWaK0v3noizPxFGUK3g
bF3VZbVDSjPZxCfoAk/ZDWGM+XYfDByNF1qaRj1sshe1QoYRs/HIo70hPMkcDkqNLkYHeyDQpzrg
ewcncWkNxGVsE76N3F7s6xPHzRdSsxACre3oOZQaKuRJjRLH1B3Fh7eKtP9jTEPo0S10CqX3+LRN
nLykGpaU+bfNA4gucs8n5dxU+WSfoZyE5xpSihQil3F8hHkLJCauGAYkIvPB1/vkB5r6G242lEPL
iN7VUiLnmawg3zHPCugitsL6OM7tAbRjlgr0gFzerfkwQl8gtIkhN5QQgELoKj6Eqv7fLbC4DkWk
f/wStcFZ8sY52GZ34S0wQU3GegOtrICaC7Nq+ZsYaeMf/ujcXWGW/QN24BPxE8YoSIT4EDhTGM0F
pBQu1QVJipXfh9Tc6wEkkr8bMnVNsDW0DOhoI76GDAXvw3GASeRqDO/FYb2E5iuTyg6f5q9KHVrZ
klnTEoLesHKWCzkfyR9UaDNYSaHwXenx+BDG8ukEnUnfOJhJlo9097ZpvRwcT4oO9zfYebs9p8Lt
MXhCzsIsCrsMZ9Jy5tVXqYqPpLkiUC1SRq/vwiQy4aCsrhkMs/qK9VYjHVIVAsPMj0laAXtiLZv4
PItsXGq7RBXJtAAzVGL30XDNDQy8t+pNdJWOYsVPCiHGOffW1ux2neZG0l3/tV8IZ8Q8wXLwBmdq
DINO0mjWFsuD0/x030mn8AhYsriaLNN6f0bhNJI8WjbC+VJj2K/YLGj+MYm0d7WNUiazexEVQrhi
jeG5iC4b62jmKGdm/JqzNdDQzR8rfgTHtYFVGOzLPhTcPUOMbwj9Dv5yMrrfqUYDpKv8s9b4rTVL
cHlYYGCLKjMYzgjtECO2mMQ9CdVWoBIjdbSNLasiXzD0Q2F+ECErCQuny6KPTjLjsa9OeQvKDNzq
d7O2uUsBTGQOlCMoxvtCgXeelNu/hWc2imq2PQJwQcP14zyXOESQEDM/AOfZgCoVDE0UubHX31Ud
byJtN3zB0yfXjrkG72dUoHdtNuv3R0P4kpf8OvH5PaTx4G4LqRn43Ex+BqyEYLxn1EIp5W91tqf7
ZG+aevleCo0YKiUFS0kKJ09cqxBmN2r6FpjILipu5v5JrdyP7/oSqEMYkkkJSjT4Krg/jkLDTY+l
JhLPGHEONYvHt8IlFN0QFeYUdOg+zjH0Rs7mD4thyT5YBNNpn17QtrHs7x8EX1Obl8J7Ionsbshu
qbHRhHUBM+ZvkL0zMTV8z3RzVEa2B6udOvVpcagZzK+tPy6eqv/qkaFnBdB8bXD2Xw+/yOqP0C0I
9P8JIzwTyd3O3somREvivr0u5mBzZ9iS7fKOfk9JwpUA9+E6j5Ov/w3mLvDYDRcWAaGTKOHzdzWh
oD+jDiWEPK7IVzyCylg1TnJYUQzbm2lFJ60hzKWd+3KAKf/9E9wVo5YTj4nzw+oTUCc3NhDRyn1s
/zNQiBm88tI9Jjl1CZ1g6m3Qao8Pxnwelk8dKPSjrGtv5KfscwEAnDxThEbzj5S/RqCi1KuyeOmf
0uhIxQxqpzm42rg30ych2Bccfbx2xEw8KlqmuKCnI6975A1OjSrfDKGPcSd60Vm8yl/AakRljxqz
EBahcHGkiW7joFPFMtreGGD4qBG4+28m1D8Z7kNbCKnAnJC2otfhHqSrGm9bc+wk/udC43IL2qnt
Rb1Knd/bTveALLeGTsXkP7BYHXtNrh/b7iXWBvu0Rg7ML5l3RIoHnGL/6lXgXHF+sDcWjD++RZQL
i28SrUvm9J3769+uK3jNRa4yFVgrHEAaOc5myOdnYkqTPCWSKYDzULXZD18GyJbPz8xQaMoa3N4p
PbL70/PueNQMY7N4CTXI3+r+PVOlbdVGfcpuwovsclJpa83+6eOqxoLOpYzv1BU6/QMBSaWEpTpB
uKQes0cX2t90f/ufEUenYmGGVMLRBAKzZn8t3u4DYHG4fRVeT9/xlsCJRSuXFPr+hNDG+83hRfyE
4lD+bgVN3Cl7r4zh9hxlIjiUmkRgE1w2zo8d3yG5SabsNKNrU9QxPgs1suvbZiLDXB4EWJI56+ye
3jIMVFsnxKb/gJMIsPlPGzHNctZGF6NUVG5K7Jo6K4o+1YFUoNhYqjz+0YeeXX2eeS1tNy61tm+H
3d8WiYdME1ReqpeVsT5fpu4AQ6DvmCi3iJrnthASl8CeABJLQ4HTiYkCl4B7YG6qhLdQ2buMrJm5
N324AqnO56lUwUzBUKG6LH29ZK/ZZ8xLnaJ6ehyn453xyYLOlQKtFrjVHyfrNqlYTAdQz6PaxxwD
D++X2tUX0q0dAAtbV6tY4/gOQMkProcrwEAhmVNU4hykHyAmgBVHRxWlxJYvzHZqL9Je6wvgfZi7
d9wcBsjW3KzHLHV/aQWs7bqgIBQPzMiLcK0TBy0cmB/eyI2QBRENOXy9eVWKZ0ogH3AKUB3HnNMh
gpdQ849VjUbVNthXjyD2AcmPExzjCMXSITfiOHslVGyRoZc3vbhr9SDnFmrGOyPAEbOIT1fOotj2
JAbzoR+Kr1OgYNVpjhGtYvxLPPkeZ4RzKMNTGx6R+GvrS+2zC2iVcxXUQ9kzFq4eBH8yaT07Kv41
0s6Vl4Dnep2Rt7xtOhCRQ4IpSXQD0ttl3thc6wkzBXyKaGf+kfaGCDfdg8sLbFkUpBhT0nYZRsmN
EaEmZZUDB+JgCCwahSo5HNXadZEjKxD28ZM54FFnnwETzMxBoIXxO+0EikkWep36udEqZuLHS0vI
MEFqIqPZf1/5AeRT9Yk+DdyH61K/N+McMsqWj+wz2APUR3uGN9vACwZKk57vVNv2D+aIuJQg6yWm
SoMMFW0/7uHFUGuEc6fY5attTyd0zZwSr8NrkJdc4Ke7t35MWrxfVhap+bXqsMPhyC19Hl87Koq5
5UjQZBnMk5MLv1g5BYbhgk+r8ccG6NfAc9xSTy2sAv9LxLDcLDm70qPl7QHXr1Q+Oizn2wqKQ58f
T970yzE5nVVHnxX7HV5ldsu0x8RmFtRnoH/GD1c7CwRm+Wu7RF8AaNsrQg3bdxN7C08J6K6oSHAW
vVd8Vhj2suOrQyXAut5KPs1zxRjPWveaIa7mH86w4GQIfJCCzHoC1hbuvTqvr4nDOVE4Cp6sSaAQ
em3sXfK9fnOOizGUX4HuFyPv9VTxqBCordtOXywMK8X1FOlf5K1cPxJU3VJdRqvCKov6z8qyHjC+
6k6MgTcBac3bGrtCDrNVUY1qtrF9A5Fl/Qvf3v/T3rL7ml9vEwU6i+Y6tTUd0l9sg7HPl8TI03hs
y6f4oNSWRDl0DxkeNRV1MCxw9uCyJi6f/luuWyc30ULgcM4ULomHx/BXR1kR5YbGJfmGdHXSJOPV
x9vsy8a44y53YvHSPQfuqggDD52UojqGmKpCOPFV+KQWZV2S1bi3AWlWNuC9Zj56WTunhDqp+HYJ
lbWDwxk+Sg+PYs1rj7DFn8v6UlmOYUSWx/txs5wTqDBZQkoh5Xh73/TXjhiy83SsLwTkBWtc1j+h
NS569Xhy48QSyZ/L+FIaZBabEv4bDu611Pxu08RZZfjPbjN4SL5K8yk0Yo9j63aumELOEFYrHBDP
mARx0As0Z5puuQ8MGC9nbQ6sqmBoTKO5H1TJut92lltRdEqSpYxU0cWOx8BPExljcKRfqhsM2pMD
sr+raTrNuuLrd3z1K46SxMKsZiky7H2su80RgQCF1R8PjJJVZSvkf7KfREI6O3SV50XSVe2mshAo
t0We9SI3PsUHLwAD8EtsYSpNFYoOOlV8uMx0nQbaLren5JfkHsjf8ik1W88Jh8Zu/izOsLVdo4cv
AY7CT2YNz1Nynf8lVldiI6iafkL/IdoWXEM+v3uLTFddE4dhivv038Stun0V1uzys1QhcSFl3Jww
W+o8SWS4Tv7zz3NUHgp+rGEL0haWTbjkIqLitlE4y0yb7QAxS6tr/DEoeKRGVgQ24C8Dt84vaUeK
qiy96sZTj1E9cXuj9YRElhDf0m2vn4Q47oPGi5K8PwQt5LUCsip7y5ti2WKomimd24SKKkwIi4Mg
Ld8SgSrG1SOODVV6Cndj4kH30YJgydvrf/DzCASx5Tm+CNqqdPDc1cHGry42fEdZoQmZv2cjdhFs
4xWcpwp2onX6Vrh905PzkkmxYpcV1qE97XVaN5KVhEptWbRQZAu3Zz11SAczf8SNsmUhNMiIWOPY
RtU/Kv6OIu798zCcckhMqW+/5zPTiDTqqA3pAWyb1sJwawbNsZudUuERnMXlSBep1A589743Sh4u
yFUhfjx7XlmAYx7DenkDkuUSQsQ5HNxK1v+SFrb/bXZdIVvpkfapIgBko5rLn50MvWEoKEVtkMZx
vHLvaHE64ucl2Hr5slDAzwSSmYGxkwlJRBgsP52kuxm/2ge4kXmhQq9XtIDiUVxT616DDttv3/rx
Cj2wPlkvINT9hNJTcABace38Q5+SWONEyRWzvyU3I38ZD3kUGvshzWoXOXSSYZAx6j0CM+Ve5iLQ
LvxDkJK8UsQOC8zFpBTpPWiDlhImvlXq1YY/4sVcw5IBSsHN3YzO6zVNjpM02tiRxyKgyz9+qtKu
zZo7OEopxkqSJnkoA99Nb7GLp94grK8PRrPUWc6gLr9rIXUtXBpKVD5pr61TH6GXERMFAtUOP20x
Igcz3Drz4XyKxoQKNKG341b348StvcdjqcyJF7WmukZpM1+gV6UPi0TywgBnHoxEVvcq+QVbdNST
B5SdlGxStYjG1fLlvRkSkNo2UsECZ2pgiAZ51eiVFZoHMvcuEDmallSaZ7IM879tzuRJIp3RPOvx
NvWydjfkEbjTBJe9ZXDj9a6K2gUxAV70xo4mpuHT7hdmEWJE6wBPXV/uhcwO230pglCi8KK660fA
V+bIGNE6kICsHlNfTslj0A/ZBTTthgOSAtGQWzD6vAAYhc4YLwgouFdZnNSH7CSdrJymOWP+LgjD
eA6yg+KGIGk/TkuAjwN/2Rjha/d9gq9bFnoD1eaZeED/DaJbaNzLZgg7mY9gqGjLDvswGP/KHdpq
hykeDUYZL3mHfbOGMblFlCUpn0KAqDSf71ZfXss9ZgEXjsKB7RDBFD8dlqkZ9wK+Wt/qwOMjj0d9
UMGP7s0tRUqsVKOX3tjq4MUKIIiityn71giYyaEqqsX3z7jJvc0QBhbZv16xCjhk9rzupk8YYvI7
lxM66XvZIwybS2g2H/QW8lbgzG6FmWCk6cGKluEqynJJFHR/hN/flE2qn7u7td0vgFw69hBgNHf8
cL/6WjryXAhtpNL1ddpvG6qshl/fcL3/UEBvZ7WhyzBtrb5jsgXjq2JgCV8Jyzd/baAJ3MgMhZIh
0C+D9ncuMWHChr/wKqBaxuct94AIosDuIoPTEF2dsox24DVdYHIXHWcCqJI5MJHlZjKHfagx+uwz
nSKeFBnxjJI+3Puj11A8cdHWEI1HHPkjxRMmN4M/GIUZU/JhE+ErI/5Z5Wz8sL7+Be9Re5m4LjS8
lbBw8KPl/OlsbyawazRoTyqJtUZPqDkmV5buDdofn+xAFOx9MEVDNUDwZVwtD6Obwoz1fiMeiRxt
pA3VlIjVdpNg4AFxdXpTye3qMwKIL+57YcucuSCFPPJ9QI4klH0/HlHyW/zppp0x1K1l2YK8N9rb
lCmJkWqeqg7383lv/3dYwMKsXzA9cnM55xgb6gEHS81l9POMnI/emXP+A68+QDN4afaxS6MOVWo1
1ibaWicCsQ8juRkgi6j09Jg9/sPTPeB7nJejxbyABGZVDdC/i2dqZAD+V5OGl8KhewhTm1uUbXFq
ZvKyiz+Q9uauISXn8Tzl5ZQurKKNzFMkxJ/WWg9jOMSBiWIoWmaVfkdOJEYYCX5U+x64IIwOvGFK
BLErQhfXwG5WtAIma8obYwJ7nFdGf5oysLEn8kjBAsektYDTzkGasOqSGxERA5iyjKy6vNedy/hC
cGafSKaY4Li4/0wV5zwdyL+zmHLLCjlRvP19RpOcFv3Q91Gnf8X3ApSiWgUa9+SkXQm0PKTyRjnQ
XElLpTpdfslS7ZCFFMQ4LOHfmXu0yJEwyVij3EZdQ2QwYKPHfeBxBhbFJdTNeqXhbSZtvM/vW937
ufnImgXVzEJr4BMvBwoCuYDrA3HGe/U0AyWLuQJeELLbLg4oS9k/G01Wksrfco5z8erCrvCzHpGA
kF+QAMBAvDIhl1EGJlJaFWYlnjRU+ZU1JCp6Z+X01iHJD8Si/yXAnLy6oWPTYT/mgCPFTky9tXU8
rnWWIKdqB9gakT4W/zE/BPcqbvrtQcBtHIh4TQK3I7k+ShPyZJ7V6c5FebQfK4ig2wRh4TDFP9b1
RHikBtRL3YY8k6kLoOYC+BErrQyz+encX+6WxFlzFVJxnq6cyHzw45ht0UK5Ul8MmVMhHZjvPRUd
wgASR/W8wf8lax2b04p667n4s6/ccFWVolffYRB8PWQXMCsFXAuoSKSXJujALQjYhqlsvwrqH5br
6xUvhAyYFSFw6O4jbyJqGi59o9YDJiy28MJyBTz6WOtd6rvegieYAHCJZpjP5sH2qKGrx8fhsWh4
gIkV22410tMczjsoUDbrsw15u4JPk0fdTrI4sGAghC5FwqNpfqGZ4nJuETC2bn4tYVk6UXpVAdye
q117+4dB0E9agfV4Dl1F5+q4DymsDHtvv9q4lapGnS0jcw7Ya+qQNeii4/9+crxdprMjjKZ1Ht7K
Z4DD2sBt5FjacWIm1Yr67T2uke/MqGwPLRWjyx6dO5StLOq1SV0N765g/qYwk1GqYUqiaFavPK0X
HVqDqAl9Vhprxw2bM+CifBm8TIYpHKNGGr99w0wGUzc3WUMrCERyvyGMNg8uHwKNMbpfYGVoc0vy
QE/rH5edritB/GdOAFNn5d4ya014Ne7osnZ//T4AEsMQTfFFdaqKqP/V0zvUXLCOcdVQ0q00roUZ
P2CXd92Ax8ANboXUadN40TiK3GSLcGaRF/SWVqfpk1ezNK9QTJAXb0ZtYsmmZbVSxz/5auERxt+7
CmcgGL8QJpMjGfliSWwwgeSif2ZZ0X7/Sor12NTRAcGvyEqpwHsLYhlJMpd4lxTC86DGN6Tf/xfm
2gocv1gLexoyn9LA03a0IUSuOpRD8FpzXz+vfuW8MNTIGqAhM3xvtQab55VM9wAUEe63j15ZnzJY
SLjLOnnQmV1YcXi3nAwfiO1Y/8MGw654NudZuIKAf+dGIW4cOYP3zRDxdt4G6rTVJZDWpn4qlQaI
cighOeucgbiHjiLNJFHrw3ThdMYv53sX2mSs/BB213C/9fUm3kFwDk+XB7domWd+WJxgZILs+sja
a4YpWlN9bF3tk/VTw9n0h+C3F0Up8MEw5NU0iWjVaFA5bTqRl1XE4cwdL0UgY8UsIxZ86A1CAGCI
oGLfK8uuuKVtHiIyACsEp/kwKHo8QeRyYJ1kELJUfqz/tY/q/1UpU6sqhabkETsRduxY3bwpcXQb
QhaXyLSYL4cTX+khsMUobaSEqFoUB9v6UU2ZjS9LQFhRkAp/dIy0+Ev4OzI9cNbBtkU9z/8qLNHZ
T6MLh7C8qcZezNotiJbBk9UD0c+tcmSoq3Z5aTbkckxt1b9b9U5QZWCugMV/cx+AF0dX3EWTfFjB
fO93YRo84979G7hnx+vK1Rvv+EdoWljQnYozQHSevTsgQ1n9vbBJkFbZcF5SJA4mxoQAv3kDY/sT
0MN+/Qy72nUkHpGA+7FnaJzqieFu73Qyo/NEZW6xuTNcpMdZErxlqQTQy+jqb9gEVLL6592Afdpn
hy++OMQFf824onMExRUiUNMrhw0J04Gfq1UUCr7QWYUWliWjfv4tlzy1i0SKzPBh4wQlufaue2rw
l8wmiXJcz31o/0qmS0nbGyROsUJhTpIUWkqsFbOnFTh9zZHJCw7DxEeTemaqNtjSvxZ7Yvsl465U
MtnwjWsLz2Fa/JJrYAaTHhU98xM1K0+sRRF4Um16DVjOQ6mNy0N4ntVCEij1SS7TbvHGDTfpEOgQ
pYnjMQOxSbaTPJvHesZMP4MnebEZRNE1cAOpMA0XEWGPWBOAj0Zuw0OC8stgN7iGvYsAn6xJ5jun
qHyEdAZnzPnikWptPPIx3qQblr5b2Wlp98qyWRrBzetSjJJdaDHRTCHSs25pLIrcmnkT+ii8Ppgl
mrPXBTV/Du0t2Mf9W9tRrqhgEYi4wbir9KNJARRqEqtMnv5CO+Ki8wAWuRMaXSMSAkRKxM2FWumK
6A5reYzk5krsVH0BXBzrfSZQJCvxhMi7GA9rzgK+95UMNyhWJG2lTwIMg3pBmSCU1kumxjt+d8Y5
URv6oB7/D3YgRI7sTmwxBubXBqmha7UuNVHJC5tfeOostXsQpsCbcCzQVjDjkoKkfj/K6cjyT12u
/f90SrTxMemYDGFF8ryw6ulMClAGruAKN0hYs07QRGE1UQQUGVFeZWOg0oanU2SZyJ9f0KrHdWJ5
sjRCU57m/PpfiOr0vMP+KSsso1jYiBjXLkbu5at+IRjDEn6TqFtVYw5c7ZbIl1bbEzcKdAazynuv
jBTEcBHx71u5MOg39/9wbHF7YSPsVHmosQcirjV17hJ5nWQGVt/qNtgynoMp3gKL5D7s8LuM51Fw
yxpHrUPEEIzdH/ezrP1n+Ij3RVpzi9IZiNTm9ygsU9Lvg4qM+wH0rN70tUfs7S1sUebqQFfPC764
UO32nanYEXnXMYfsnuKpxJEgpweH6cXcjEeVuGyNyyv90YhR9rbagE1J57AmaawzZb+e9+JGA/U3
UcPzm0tB1cbbcE9nG4/dnX6sAYjbBrZp0huG1CKi9PxAaHc1WYgzzmP29amwBNjHjwoy47euCB1U
MIlU8VtoMxXhWukioTiQDp7ZzInjRRqO7ddKiDMnjuv6AJVdA0gz/hzPvQ8RF5nbdPjiEfvAnATK
06hPEbd6KowU+5GGdlqRrn/4ParPYP55ybA0zC2ZjrjPDmxpy7WJ1yhsuNrp7be9AcQRFPKW5hiy
rJX4Sj+tRlZ3mIQITOH2xm+5OF/S+o0UzzqL3/apxMLOZ/0OBOPGg3i6yXNoGWvONjT5tOt0Dkfv
XhlxtZ+a8D5W+NdCyLDhPgYodwFuPjNG8EjwrGek6W7oz4Ask1IffqOjuYvXaBUbm7APxvrnMvx0
CskCLDrglq7MmuTHBCtDydHaBVwykCAStjhanc6/tPAJ5sIE08efUGgw+hEXTr/mw4q7DjeMBZfO
BoITdq3XfseJmZrZ6qpF65sGpUehYdZyx5LD9NMbEnIuvm4XpPNbMkVQwlgpoErykAxNV47NXKBH
qowmA4M7pZwBo5K2QUDo1E2ye7oSpXvf9otZKx8zFpnweI1gZP6nbnZMUeI8ihqcpbVLQI+OHcFT
zY6vVmZvoFlyBKNmMfUU6o2opmdfFhFj85kRJekwLDVY35DjIkFK81EodJWx/dyk8YsFCQgPYJLJ
SXqDjHP1+JgOaQuH87oZqqYBYRzStApnHVOSgI//CePoEdqA+F/HjPdhnHQn3mZoxNO9hMoP6i5/
VL+QE9r66+oyKr4mfI9MrgpkE7qZPGmKFk39MXI5v/fGppqYo7jksNZXcmlXOaanOIZZUMTMMxe8
10IOo3kDaZh3Nrd+Kpg4yZLCeneuu8bIYlYlIjIMfFNi+OPqVbAVmnMwb+912lwQssla2ulE+8nO
ej93yajIuf+f1ouIVCH+0WHz0i3RaMB3WWTIz/n0buYRCcTUYomWT2lKh7ghmpTwyBTJJKXDKlmu
w8OlMWVAi9rjXxzfyH0VaUzpAFk9lyrIUmN2dq/uQ5kGS1nJeqg0nk783LtsTy56X63u1PjfFyhj
l1PRMznsMbm9G4XymMil4Q==
`protect end_protected

