

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
AEDf93kkZknTAYDLPy4q67UmP9O18ta3jK/RtCkxR3ZqpY2KlRt7rza1H96MUf+qsK6643W9A0n0
TP4few4v7A==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
erRjv8zI0elbdGyufePGLqKRctW7EMRy4ag4V3lsqysjcz2IbkoY32VNXZB9TkYq6LxuID3xgPR/
/dbN8HKNlVJr4fTV1LqzlQYnx177n3iaEwIdtrjwP76G8DtyrbDzV/JISwzd650MMmyKJtHnC2yw
alWuAIIBdbSW+HbA0I4=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
gdHY5LRWuJLwhBPcRYPMx1NPD/GuGCtHF8ywmbYLyoAM0rjTxb8zBoSHfJbS/2vKpgG8RCdZOknj
FMJ+fOkJbpOMFaFsosZ9XfIryZEhroI0pt0zugw4Ha2XsmQGqxGDd3IyGRBNvDMKRw2cnjSZz2Oy
H3SrajtWuLhpP/vuSzlhtnqryvgbp0USaL81fja6LLlPm2jXTcuqgEPsJwwUUhxjUSQyRtABTEvs
3Vjc63pIVZUYkpkoaKpA4243dOoRhazlhTF1c2Dp3uyCrdGZU4fWhJHW7m3Cq9Aw1murzYGrPLS4
eQrf4MTXbiMtIPpNK49OUBbEpUuLfnDwfATFaA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
fCQs5S/zt//IgxsFc+FuMl79LHVh3Px9B+S0yADLC6MfIDCRddIdSKbTMZ5DlFrngWDJwpd1JzqP
cRXcul8iGoVMrVmrEStKWXi/mhtK5UkWTAd7hoyj5zcI+N7wWWxU1eBAeKZQ7uML2SLN8mYzQYLY
98ufqGLyMQeFAWp64iY=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
rLzkYB2xv7C/3jKaA9rJ0Hz1NLTW5YORm+QksBhLo7WkyUXUd0Olk6yTtcSIC82lRfBo8f3njqY3
dhmWfikGbTNV7gixnGfPYVUvZg+xsJ7adfqwnApC/cK5eBJGeWXZ3Z5gEbLOhuRw/04o37fRIoCo
Rt8ZH/C+LE5As0rIpYw6uzjL55RYR91wP1R/rUwMQTNJ8XwXPkAbkuyw7FWG3uW7vEvZ/CGu+T1f
VDCUznG/Mry2818W/OOR+t5yQ5fYiXNh34gzkO30FRWgtIR7ZfOn/fgLqv2Iaq5XPzTdULGOHjv5
Pl+0fdEaYyo+sJ1yt8Il53T+ZdgLTjEgv9cjPg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 30320)
`protect data_block
RE++apNNH3vCx3AEMdlGD/s6c/cf/1JBN7w+qh0nuRVodPFNto11CB19WTH8jcFFViQisCy74Tbs
q6p23uzId0LCld8a6nDvRkNzVQgBy6Urg9Hzrql/LJZY+L3JsIHKXKcMVYk05mM6ZtTZklxlIwlf
eCo05ukOpfSnxOScNMV6tkJrsfwRP/XZM6zlqkouQgiY6qgBkqR6W7XbJg7XKWBdBQEK/7NDz7+L
MQ1b69cvuCITc3J/vF8mvhXny8tdnyLEhw5dbAtSAnXhk+F3+1bU1AhFRdJYB4s/4SU+snv+7ujg
9XkDT4haYvwJXD/dL6mC+qvct2w71N11txutE9j604o2SBDm1C7nc3UUD2olA458rf9cYswKGkbf
svR2ufCV9Kikf+PynW/WAJ+qJXtyZ6AvHTt/RMBy8VWIGQm1bfoOB4bnyP4i74m0ld7iFDgNF7lJ
yPYgchUuZsJPeQ54eIX9onLsoI0Fj9kCaYJL8jIQuxadz216rVHi8n6aBVJPFgs/ieFk+QVShpna
degP4Tu2aYJIMKb2FHiduZjCC00ft9vEa8i+acLoeg2ZUABPczaGyyYJp01n/brg5vkLcp3fmkWy
Cyf4Fj1vlFYysfpgP4/coeyCSczs4KzyRzJrhOmqpIOCMsAcv61UMuPLfQxCqS1NM6Xsps2qjjxb
NJI1BgrCMVvPON/zE4TsfjEJ2rEkbux/q7g136MAkv/3acTpvLA01scZdYFGPNTGflndGoV46JUY
iyFDO6YsI1y249K40NtRM+FYXMtDll1RhNCv8df4XyG6ZtGMyIKprfQd/wxRs2MQCtzxMLvBr34T
lrJrmOn6XbvMAQNOi9PXjrvsc+91X5yWBhaV59oW4+faHV1uMVZJfp5EdMomR6nM+LjY0rQilXM/
UfetxxLpj2LPK7P43F8HApIvmXO3H/bzSxsUSLA/vS4gk+wqthJgU7nltljkqutNMojAyjFkAQg/
5GrYho0bOpQTD8RGf25LXhlumiuu2OACF7YFjB7AtHdgIqb7thN5nT6Rr2CnQ9gtRkJ7POMv8kXS
bB8ImxTJ1PGAY658/IAys6AhSAoL3ZgVv5IWjSih8kU8I93ZntZc8APk4KZaibOKN0e1VO9V0HEt
8TEBvwiamN04HIpuyhDlx2lELpOds5ed5gQJTLxKRZlSpwbmJfWPYNlCKRlL/GXncvpnXgBcpD1I
JrYLH17RNI61l2PjxuaMNr9iqQ9/r51dqXggUfq/Tm4I7iJG18lXXpaM3L4hT2ulU13qUcB+rtxF
2PShjFeedUYAJmlEPNs6LthoECLLnETf71JCD8GRB7t8MmAlmy6g75dYiWvZwfMIQTFDWKVyjYYd
kqzDTbk6CjOOwzpsfQu0iKa0KVEp+BQAsNtSe6/bZWCv0TqNo73CFNF/W1JUdUW4onYUBEgegvCh
MuJrkMO2Wix2DV+r3IAibUUldwsrLbR+S4TdLdtN/59GSSxA49Lyh3d865e2HvcWE1U1RkwLv066
5W3/8NCJ9iRP5hmBZXTNAKWdbz35jFOdm3X49SJmHn1wYjnNOk0uLoXhaYHnpkfQbIwLkKQK899D
mcYfBsl0PiJzevCQyMSSIiOATR8tvmg/u5KhFkh/01QESUQv2WQDNyAKeYnIkY49AMHWnNfZxSWd
fED4pgsUPo20T7XmNsd3ds8O8iPXl/mRinfls0xu7ZYtAmqRWSgRBEEduy+Pd11EHgr++rj1r32n
K/+dboAK7I27CJrWms0QxuqaRhxMdREj/zuSdS3EmjETcorYfpYRPQVj5D9+mkK0al0A5brHEYnm
/AXG1RR6MYsuyGfNGytVq1CiEtCcqB1xypPRCdhjmNaQlQb45l5xYsepsBT/e5Rr/K3dF/KcUgfr
47VL0MJ/MlLDcUCSuisAd9UFB0IQoVeJ9v/1w1V9FnjSFZaG97ZZqx5vRCTmXGb3l1ffiPrOyuPW
1q+QWyAuhbIcHVfR5nzcbGsDynyenkvBOcsTk5gidLb/+VOvuhkQ6KsRpfU82OVF7vkQ6G3guxIj
JY/qzXB7hG3UyZ0y0Lr73ryn8nJVEZcRBgAt3rmNTo13JBsjNUvrOmG3HmjTILJfFRC+ZR1Q/kOy
zt3rw40LtxPOTPAF8DNZclpYNZDuObGjSduU/39hMGajBafW6sbqVp9JYmuvmsFCbjAvoSmEWquX
cneFdmpmgS/kVqrrDNMtxLc0Am7CetumnuGCZjL0KeOGNA9NkyvYPx4iyp0YzZxF07y+DE9mOehl
VXbWTK7oPJ7lnm/Eo3F8PjYRVxD5Smqv/GoTXfwZ5yBNdOJFe9cvQvdxaonVEjt5Cc4Z3+CggLlL
th06TCDvMcmRpPcfZDzOoWt2Rj5VW8lEDiYacRuhTVhGSvDcCHfi/0V9wKCVvMmDWVrvwb3Vf8gv
dDYqGmwsA2jrwqeXAh3pnBTXanp2w3kHOXLQ8A+ni6ZqnO1CCSArEzQLBphj0FSQ6IY1mU6BF+RS
I0aFohz2tzXqRywQWThMOsDa/fRVxCn4XJdInFjG4srgyGx2z4e98fb/A4r7T7kcdvLcmRp/apGh
7lk+/+pKnUoqVW13KFCwuzLEVweZwnXkWXoO/vPHsD7otmDgW+6278XvJRB3NxFfd+uIBdp/j5AP
h0t+mGsfc7kjde7OcaoAGosYpsNgynK6FWPM5JOmRcXgespIW/vJJ9CJOXqQycFIoMdRZlETUSU4
JKziIOY4AA3pIOsHxHgj3riKMNvzg0gNdlgoKb7QVoe8hDkz3a+G7SZsBRKh6Y3E1tvcKkyyBQiv
G1JivO53pL+mcrki2vFufxlvY5nhrM35HybxCwOnRnTH6QLN8vvHGaz2qAUvTQs056GG3qofaqRY
yQdLd8HxIM4dCC7uszkf2EmshHw3+kt7deaLm4WHVsEDGLPhaH2CZNKlq8oA1MdON+eqTdFbHNv3
WVC4EXwXFfINSgJWt55CG2fjsqYpyu0/7+TmzQH8/kKupbzDaupg3uWvwaFoAnfsqo8vU5hLNiEO
Zksfjzm9Y0g0sGR03pTw74S947RAe5w+WBpnB1Q4FQJTp8yjCJxNfU/Y15yu7ts1r2Ov9P92nREN
82UDkpFA0P7NvYGdu/AMFV7R+N/RghWU3FF6bILR/Y2hD+c05XHmmCXtkM2/dERBdr7aCXcqDS1I
noFosECnlSL6eWPT9qbBS7k/6w47gLRhAaDtuJP/yJSKycGR0WEWdcIWciXj8w46e8xgaZOtmdC5
/wXxkbSqUsWXfiN9Hh0uYP6O0YtRvutxeogilxPiUtJlyKLCIxYv2KksgdB8K6oPbJR8+HgDjVVu
UyXHWAq7jk3XlxSHX3+WSR0/mrawks0jOGingvYEZEMLqFy42FnxlJD4DpU9RgkVV7gH6Jjs0/Pw
OGgsOsoNz+AT7KvzfpqVCMvmFGJ1eb9ODIKKskyV4RAXNX0eQ+KXiIHAo2cliT4wikBJVaIRTz5F
ZooUcuGBPwT7pW2ZfQ2zJYsNK52inRKHCsxKixrQgDkEuU/yCzoND7vQnBxc0ngnVTi72cyGgCjN
uB4Qa10IGz80kCGtxicnfiwlnV/TdO3dFJTu5G3L7s4jCS1HLBpGXIRTwaOcsu0IEOXUULNbZXFJ
UkkMjRYqPiDE0rYw89AM1Gpg1cczIn+bfn0V5TFDhfqRKJcdUIPJ+ymxBnqx1Q/jgjiU0z2w6RS4
lmyNS5QFGiYZ+uH/wBke300vHKH+kDIZwII2e+8MpCSutcpkNohsyU0LO8lc7NdXb6ytKc7VZJqM
o4ilTxUOIez4NQM5QEcTHZp/V5bKNt97A7hXMZw0jyj3GiixmTEa9U/00vwSjfGrF1mAS6gpouJR
fhmm1O9mM5rqn8UT5Q1BIrEacGMH7ifFKf9zNsdDND1z2PoSBvc2ZP3YekTGqZ+AYWMEbckigvlI
aSVStBhHjIAsptEgfacdhqBDLo3LNRfp8Yjw7vCpNwkvpUwwD/Sk2utNVyXc0IL67A42qVDNmK+X
tNAv+i7mfGfBJatolfyiR+Kyih30kZOJWH5aXrcn5PwW9x673B/CbYHED/BLGUWvRAVfKFrSYPZw
5ATW0wmmIXZExbBMRjEV4gMBPn5Eu7Cnec8FRcbPHyq4/qwmUlvnEUmqjtx4ZnFoWf3YSdasvUr0
HN0oFHaD2LhP64z82rcTpaFSW8ZWjQFyX0cyEN2jYVWlmI05av/qo6u7rXefsC41Cs9RxdnHqalg
FLRCwNUETrnYeAXsrMmHh0Fc7gk1aYtUx/TOkGZMQrXhipgApyu9e27PYf+EniOZOKtP8NEJ7mAF
hAVphmKirKJ3IB5Lg4MKdlQuvffMySxLHgiGT69eFtCaYhrtuZ10Bkz1Rl5mX+0PYkME39Si0FMu
7DXKi8jIXruMwYGAuGMAsRwv2UpTPcxIrWguRSzQvkiXv8C+7VzfbwKIa8SDj5Ekr9gvMLF8G9Rm
mAXrAC2GLN/Z0nysGWr6sgiv1cPguNWLes8Ft/VESreXDcnnBHJWA0g2wRFvtd2cGvVFH4MbwUsD
CU2i8CmTf9V+QKs1f/Dam+p4SV3XwQ7kPx6mM2BdncgQnZ8KF8m3H6+nDUbQEjZmKk6vGcsAneXT
ethlE4wCtnlGqW7GtC6dUK0EO2ei8ZvXrzdzJswsfL0M3eq1c2tIXxQlW4YBRNPxYqD9n7hbBQRN
LD10SGd7PNrpxXsNMU58mRDWELepaBqhpI6A5WBiEgGb2VXHUDwvDvSXHooxnI+bP2HZNhu9CQLS
xxeEPnvWr5xLS+k+qoG9RlXHO5geVlpHuKJPfIrBrY9sc4bC3f/XnS0oyQU/gjYBL3XhU01OmVeu
2qNtjXrwWAeGspzh6j6ZuR90DkI26vs3DiTpTPJMuJWYxOFV8ggOL2SIgs0RViBq6K7vFt7lt1AO
i4zfw1K2rQSpcaNVKHLfUArSeAswxtrjL5uZoUdLNBaeUrfHcMACB6cAIWmlwhMDtIj8qTYtgY3B
CCABobi03AK/fT63RH1ZzhryK0hl7daS2BN8Nuylhn9pMYMjMfKgH6xxD4EvigX8mVQLjeuIZr4N
L6YM1VBwEui+Dw2SvOPAqajZjmy4lpLCSNdJTrJd7s4A9XB0S+V0esKT3JzdyO0gR5PYr4kgpxIm
fmLG1+nJPAmExlw62AytQ+UHHMmMjLG+BXFctZKPOHXBdLsiW6+zENAl+raE+th9iH1kfb9/Mo8W
GCvUJfORjn3oauPUySVPDHv3GXAt83m9PpvSSw4XvtUz6JMvO/zc+mogGGExtrd1fJz3Au+3qr8H
S9AbBsYyLg8XLR58/Ettw0ZPOpEbW0W/dE+bmAtqCUIeKvbXP/wFlWZNh7K2SjdDm5ii7Gnvs+NO
gRAa55tsDscWR0yDpW3Eft50QaEmuzwdUVwWcLqpzbhm9CMWuqipWwQsyH8gGAxqHsMkNzqfNSx0
bAkUeFWLkRCPmMjBYTRsQ9xgF/wGJ61CVeNy3w9zCEvk9SNPEl+P2tRr7XV/cj3QgoLCknb364cS
sEMN8X13h+hA2br+sE9Oz461AUwUBj0VppNRx1V4rlUAxRLeS2TupI1j44AUtLCBdwBRmbrUnP40
zLyOvBJxMYr4VjO0mWdxcfercsGLAoxIXi7E+8KwZDwQ0j+omk5ca5NUrljRN7dJgOtB8AwX7Cab
gheyeze2vplLeSSLEdiyQE3/T3MCYHkyWn7HPrZXC0++ACRBOaQodmqC65KwuxULP/JeyQ18ozA5
I9uSEY5kWj7jZCXmxu9qixJmlFRgTeFXxxjXp1ZYUQsXVis4PtZ/i2R59a7ur9oFHftE4U914dO3
AP3gxOIquvQxrSJrqCABhLp26iO9Y2IHahJtDvkWAMY3CKDZlbLXApWwYguTGjyveK+cN2uGlM8l
FN8Bf+F7XU/rbcKSQiTHl8njoEHK0hyeC9Q5A7raTdSz+CoFvMPyRMMlqku5nPO1jJv1TKwtbpcG
WkDRHAfS06RM098Sfr3RTtyr6OIGUY1FOGH0ccKWx3ymYb6R5kATujU8G/U3hYAgf5PWrasTMzZQ
G6lX1GVzpc7P2S9tBtTY4XHS/ztul2hgJcsVZv8N0b3y0U049eS82maKE2NgX+aGqAZgoDbm2wep
vdXD8XYEl6Aegd8CIYKtLfz8U+/PqM7844uWGc87ceWkds8rPVtmhZsA5Kn9rUI3K4q/VfzE8O+K
6LTHjta8LCb1bL+k9qZeo4DZaSZttA0TRVaPAvSHFfz+o94wUvuYemtRaar+lOQcWUOs8PN1Djsg
tNHWr9pEJa5TG7/pPsCGeePyxpOSR6tTWqxVBVpQmjIJfAOpsOmwXny46U7TNr9jfzBpMfAMEs5p
X0pW06lC0oAockNnmeZ+KZcWHA742JlKJ+TcELbwas2x/2DXKcmwT4NEfoFTCi0yvyd8FuqKNzr9
PuUoUQUqhreYpk2Cngkl7zyCGvP51bNcgoeuA8+c446QsEC9QjA0ZavEFhec/9t/dILhVIuYWR1p
bUMwSamKKmUMEc/mTi+ORCIsUewtbrwnR0ijtkRqSOZVdf68oQ6/3BSpQB5ARAvTiWo0FqztoLGg
8jo6MEJLoInidRSk3/COPAHmyu+2hhDRzFEgnSHzgqNNzfTx+GO89f8oWm9p+DirppU2X6pslmgr
48m/qiogZprCo3VjhhzjDL9NyNDOgv+XTvcMou4cO7AEWIOrhjG4U2wpYq6xqfkyUEPSnyozo+Cm
BlE2oKYRZRQ6NARKLdgfyalwEm/3wc/W0zKcrlp6mtCLXLa7je1YuacE5u+vaq8AVJwEp9uW+8cF
22YArq7350NuStGQfjnwFd2RMg6k/3jLqCQiIWyJOJdJ7iYYbYtoNe/7+dwmfjw96Fai1UsKFnuH
1iRPF2O2PnHr4Lc+Ew3WezkCigRIq4XBYUvzVh+jR5WQ+kWWJ8oKzw5mLkr6veiSHjMq48V8mZg9
XSS4Q9/MFun746y8BrqdhIvIruMNvQaUyf5tsVxrHcw2BZGXAPWi8FIOgpA7AToj+VSrgvaFJsMG
8NvsC9WwuNLkFbdR/fYdvKaolIwLGjp9ZJ+GoD63QhoWIPd0oAzpgCq/zvbOtMEtjjXq1quWHBuq
H1H1Pt7M4P7v/ar2l/4b8b41ZznjpxvexkYU9boM3hp5dhQrf2cnl6SYEE1V3qiExorpFK7WEM2u
YHmU2+5Y86tY41m4NqSCTRVh0BB8f1rMdaVeelUMYFb86aSlG8X8GN8L3LWvZmTKcoXdn47dkA3A
DK+2YaYeH9wLeJ7xyvzspdrdhapGxWRc4NNFaWV77aNzP/aoXyossmOEiXK5F+t9EchON5SRJ5iN
y1RonaiS3RzaHPmDE28NrWXHQhNAuXtr1rii0llaXKdoZtlEtckyA1hFdUvz7vJA6e2RAXTaRQ8O
T7oVMhcfz25UE8qfnMCy0fEPvTIPBSL9zW+iNX6MV2sdOrPpirw7TWk9vQ0KoSeDZk6iQP8oOqfj
FeDqomBFjWRJ5r9crhnT9cZQrKFTl7ScKVnHWItSbqaWd3HWAi+fZPnBcHoN+088mU4Iighwz7Vw
5FuA1cQHUWLf7N0ExpHVDBcQfAQSSVY7Wi/73M4FK4f5a+XPSGo1Iat2vJB2jfSQKuKEqTwfNlfR
LSG5/RjTVIu9+GiL24tf6vcqO9xGWhAk5Mw5bCeXoLN02KYmERZVifCNo38d2A+lP8iwWlLR+WSj
RToHHhtKQfpKDkqoNcQxHeKn/iXkp5UI2U3igWwGSYL8ZiP5kM1T9QMKskrTB9gIm4PQ+SZrBQcb
kEXrJPjzRDnQhPoeYNjjbf+XARR89CQlN2R6wYS3EZG+gUGkcw+P3LhHamEyGcglwNdsZIpvh2O9
iOHzJrPPno+aRS0rJMAk7RyUDUunBr3iJpFiSKRMbwwKIA8V9OmWWR/ZEH0cDOv1yE4UfK5fTjo7
oFQxQnJXLrbMDKjD6+izPVn4bTA7ZhePw4P0uupNXvzI0DacqlKpRLbXtH907nbTGnXmMfeYpQeB
6DkOZ9PJNgqdGitLuxogx7K/xdU1eAwa7VqnPBUguqZ2kCoynRo+j2/NCk2Lu1BOv1rBYd0YzVsm
JxI2eBaQuOiXJI+Xu13DrKk+IqDzQfJg0c5kmOVqqJyzEaaa++zTyCy6+ZT4p0m9i0P8NSHphX4O
nDnLUAH21vnjWFw3fTdv5RQCSiFO6QDHhbRCcRn6XtLEJS57KPV2m1IXBlmRPNlfDLGmIdva8cpG
0L1KCAgbKpShUcr4zRHwY7GhQD8SL/mVOH1yYFNQTwQ3mrX5j/vDQdGQB2bVJjPoCVy+U78SdnkZ
haCEW8virPITXPE+OCXHRObwxRulEsWV9s+jJ2Lt2ZzFUyphkEBztaMjwK8s3OvVkFjcO8jmhfka
/LClFxDz+8TOyKezVzwgwZQ3wVk/huecgae6cDnMhH0Re6XcUn+5wIkbzxPKxokwmmkF8Kw5jJSw
baYx8wTEVH3dVxp2a4cCtrWbp6A4EYRJMAD88yuQnupmP/trntyo+3wZCVCPZyHBWmJNzQsYd5jI
Xad1746UMQp6ipcHNYNxVXtTqTBmnj32wMduPipyp4c8oUzk9UzXoDUbj97t1Fha9BWe0VxWYbCg
/51uU2i2fGP+b/8cl6BK6ZTxr/ktUfbkBZMa+K9VPlYShPWPdoJ7pMnEfUFHkICDnQFdqnRkjAxY
FAzi3VPdonufU8ZiCDbzFnVXS7gukHLZXet+hGDhIPxffD797sjFaAvCaTDtEcsVxrh89tDbpMv8
17AqaxmjeFtuYqMlnUCeCNwHHZy7c33UrHMSkE17TWRpF3cRkoM5hZZ7RQ1Dss7gxJ0Cr8mt558T
Ao4fcWBl5S/H2hAVBXJ5nPIFtgIJdfPvDf653tU2D0eOhRTqU82etU4M8Vh+500jKLv+lKfgcbEs
t9cyuhr4tnMQpMnQEgdw1UZ2NT1K1gOCxCa1BQZTF/U2qsB3VPPm+OXkDsOhjyfsc3QzvlK+R/ud
lhhMf/2eaOs9UelKhqS3VZHA9U6Gy6frA2rskSJrPIXzmgffQrbkyEmMlOG3cwAMp3nM4amawscv
XUfJ6IKTZIlBckhL3yCeIi2gCeUzLHAQmqh6HqhpBh64pGCvoYl+G2FaXNF8xAOQoudGSOli1Jjx
kztgeZNVv0J1tly3xxcOaD2+4lAi68drcWA1Lu+eYI5VHzWpovjmcagF+QIsYqdKabVIWkrNmNbN
R/NoGIQ8wdAJXMM8o2KSqjT+pqBWRVTRSPgbzBG1XzHA3nMKi2ezR1uBa+w7Nm+G7bwQwpPhDqlJ
aSX3nudontCxCE94tqs7IuML+KfQYkUc9ockdX5L4EDnC+jHt05tffF/RO1RV3+Llc0XtXHmuT6y
iWv0+u/vBSJKhuCTvOv/YTijuOl1widfvCTjszBXcqs4sen5vpXfHxWwYbWOMFS8buqHfmTekeeJ
RaDA2DIUwG4HQFp+onZO32UhtePKst86rI8wIu2MqST7VVdKisVkmpvy5gZ8nDUQKmO4DrmWio/U
cPfcu9gyvzxAkLeii4/kDSJsvtiGHMvbnGIf0PQEtnIE9gAWGgz9mF2tAmT7PXREj7TmDISdeNZK
onwE/tPmmUQRCvAyy+AIJ9oXYFmR22LVug22gJkfd5Nf/6/MbR5W91bhTORrmK7gn4D8f7eFowUL
EE9QU4Z9Ulf7oK4r1Rj7q1ZqxwGzN8tg9CTdcvQjbsiWxttQpCz9wXXQhKtYkFCetW38eedZLUH/
YyC1CEHx7Cyb09rHOuER+48ZMOk0wIr+oZ8p3bN2yR4V6egCGy6OG3LOTU98MlFXNN76UuUJ/A2q
b3Ek7ou0rYVqPQ1Tkz5cUQ3vfWMGTqTY2+3CK4qPcFGeL7JsYccBEm7JapmMMa80TDZ6Z+ONfcj5
FIZzHeiy3T2OKpVCHW7l7hpp1jgP4lwtb9dA6Is915AKC1RAC01Xtix1oMARyHjjLdBKnJSLXehI
Grm5q5BjgYuQsNlqboUqrBJ4jj3ayvzVw4DEzHOKtvxgjVjuGKGcpCa6zBU4Fey1ojRIEBGbyMgc
p4BYQ3VQ2auUr7pNNoXEm3u2ZtaczBtzmsI7OgHrCH4z3kWnf6iw6QQ/In3Fq8MjUSqU38Ha97Uc
WJijy3dQqo7cdE8DLVsvvnBx64D8psz7GwinWyiQMCaw0x8FrNWQuDv0zRPT7ssXurhQJttkfP6S
gChz6lBnNlUl1gIsUbenfF1mu5ZYHDR39IGYSsIPv/xvcNDCEvuAX8jTN/NiroUlqWsslvyGoy0z
6uTjgc56ddA4g5tIzCdd1q8YhdET+7id3qR/tt7zLajQ4G+CDLAEUGQnBs9TJE0COUG0bzPQRo+h
JQtcjIl7tbVAxlUlvR+hSOBSfGeLYMFQYYnrvzpdpZYoYuAnJZpa4y9ceGp074oPlkAq5gztf30R
aAT6dQ7/K3hwgQY3HFAoRygUqayKwsa3AZTM8uCurrO0U2+iDXPtmM1i+WLfXqRIAtOIXbpKuu0Q
L55tUo8WntspY8mWY42PoWR4LMC4+ubl2+0uv5K3mbWQuGYwGImo6tIu+0xkqPiqlv09mD2gMuaX
qtJRpQSeBGknlf8Z9G6FAY6kSMulB4jFE1odGkLNoOtMo2sroNqXILG3JRL9mdVa9JEwd+S+U/l6
BFxAVAszyK/n/D2wh3v6zc+KtQvHr+ks6pG9XE19EXS5HF17G+iXPq2dplyC5UFr49d3PxRZahsk
MUU506ZhKpctaCOy5nC1WUrrorQLtkzFDWciN1gKGps6mR9Z/fsvyZ7aSDEg/Vq8Fu9JKksmh+GZ
kdgyaf6cy21blJ5yOPQJCP3p92h3T4Bg4fHUL8ziauSzYKMdU6VuiKRIllqeAZyfoK2mXT+NVYXJ
pDbLfljWOi2mj2+2FE0sKh84JYeJuXgXATs6fgwQPoiuzLclJdtWRQBQpTVDrIvvnhUK3f666XcK
xkMkfXgdVapaQwbUc2BQaQ26omFJdEnmJexhGNFoJc2HtA8znxgDxHU1JqFrtBZCv6hzT5U7V/rF
qi7nEF3mLhufSKjUtWAuWRva5Lf8rCz7eNsZCZLWrVNe5NtjSvKaHFnlLgssKYZ/Gw6vqC0Pi4CU
91Hdj6MbZNM3bWe5Dxa8jyKr5Rut2qFrw+6sl7vEnB0Grh3ai4Hh9k5Yl5rKhJvEGBgw7FLba4O9
nF9oSWaMrJTiD6SH7/4M6F0609pNtC3ztyiGCdoRTDIqvHKhEp1EUkIaTsmmyniiubzdqLF8/a0N
gyCD6pT9Ywn/aGkglZYAdzXVHi50tIywYV76H6AZkWLoE0RPeYJvGQwM9akREq5nnbkekC2bfYUm
GFLGzRd1eNu7Sjdr5erSS3nrRxyJLqHEPGiryAaAoMhmAf5B0AG1VI7LzQgH4oglCwF8lWnafVN8
Lztib8XToC56qzwRnAB3Z7Q1H4K4FVO45fO/hPy9QY+Wg1T8In5wFJHCIfKliQ4s1I4OaFj1mB7b
rbY5O1mjDTYV9m4MQ1OjyuvVPpEBPDbj+Q45qXo8OY8Zw2nUkRFIgZWd9IpT0jlhWda3vPPdYYST
aPxMCnlY1e4ftwZd04vxZNqWpHkgzrgxA5QVca+S23OytcPjNEVb7p7NxRNBsUOuGaN4A46te97i
7XpnqJ5DRnXubF2O2WqzffUUml2iqwKUe39lsE5T8zMh1JdqbkPM0DqokB76m0qC20HkW4xpJs33
aE0SBPA1j4HyxF7WCz0Fqlg5HgEMnyh+MuAiFvHE8bjz9EDl3AaKXC0SxY5NBecGjqtIjPk/Wvtz
bGXl68ikkSUSrgYidURBesChwCtjDiHX+gPSDC1mVAPB62KKCE6HskI2moQ3E4x8owJzP2tRcPa1
fMCeuGn4wXPM1PNe9uKrNsTW44KK3Gc2SGQ1Et+7QUsRCB8SPENQqtEsuFrTyYE5h6+UieC7BFK4
AkaE8mO0uTkst/f4fzzt8yhWPaH9rtn7Tp4zrLbav8VcgI2bqpCkpuRiQhwiYDUeQ3CvqVKfFene
RqaXo3UJ24D6/Mm5eUAHUyN/WKsiez7a3hotbXFxmy7cNO+e/MYG2VaHIRZHUQBG0gmZ+Xi/LAaT
bEg7nTvUnizsXU0T9GAUsqiTLiRPElixyUwzJqycbDntCpZvvXE7pO39Dv0uDZ4Pv+naVzCHzyUx
zyp1Fi20S4wsWZAvN2ybTSwAlZ9mtQcHmB/eIKwnCyGK5uVyZ93Szg37CvWG4ocKbKA3tlrCzBWK
1siYEmoz2+GoP89AsYINgsJ1Sk4pzvT7p62hnQzaialiafXQ71Skhh6SbpApYkiljRvEvuSBEBpO
206llFASnvGlXISR5CvCgnLMLohv6eELaD4A/YW4HxahuN2FLpKJ1buwogxpDfEapPB5yjWsuSfy
eZfmmXi2D6920tcAx5Y+jjRO78K+JsZajV21gDt/ryynTKM8i84sUr8eOZY1DUKWLft/LMowRIc8
/6awzMox4hzP6vXI19Opv+6nCUCbQ54ug5/EJZZq6SqiOIspgd7tYr6iEzwgFiQ9vrdmPkR7Ebok
lxDEaiwHa4r2TFlHqwWu1u9Fzr5U7rtUx/IQT1S5vj51FPcVnSIux8zoEGf6nWg7eheDVg0UEQ3W
v+4q59V3xqdAOsgu2pOp6VouZl1R4JtPnchpaq7CWn33qMZxM2V9bIkIfw6QhQblRMJa1q/hcvOk
j2oAuHbiVdjOMrCSgikT7i1nLBTj0T+y0XRkEPDkWAQkJ/rf+ca0/rsjbz16zwEn/j+gFj1s6GGp
9LTWW/stkEM+UF1z1+Of9FZduPQ1K4NyCACyPRTTOCYTZR9YH46yHqWMTmo/cLhlsq397QS/izgO
QZlUtUuYQzWztD40plTSawneJQUDbql9IyLcvd4ErS0JSRd5yimqGc9N96uDijuYEa7zI+bOnqF2
mI70vxDKgvyvzGaYF77HB2EptWesnyEwZAk2dpACsDlVK+bnbcZPsb2b9/8/9TfENIaYTdPbajr6
MTUJrHaJnyuowYpAHC1e42nAi3ltUkkYMsFfBap3FGDG8duf3Bs3bgYPVPSyzW2Qeh30RMVe7AbM
5wjErwGPXUcmHgVAf6RRNcHuHcRoNOnsnezxD+pYuK2GOIct6WpE2fA/VNBYGzXmz5mdHrCunLKC
8hFMAOmlvWpkcvW4rxlv96ydkB0k1K95p9k43qC2WWDlxg/Cc8cIpU5/wqSp9LjkjxyWShKIKJBK
X1EuG8Y3qYl3MzVx7FR4IoPUZfrY+aFtaSRkMmq2BjWlTBO7GnnkCcFhlzxjI85e3dy6YtlPSKRc
lnp+l0byuGv2ydZikHyUfNKB896pPuHSOGfrT3+GnpA9xN9srhWKtPkC9px+QmuMoLC7uA8lb6MA
SKUkT9XPgPmvZS+oLZB7nUZbYchS3eFilnjcQ2+BKQIbaWFc8tXEGcdKbmGePBysAlxCQD7XtjKi
psmovP5ceag1qzMM0jXIMekmEhFi9fUGpcvevTTvD+0PgpbKl0bE4CHqP5UZw6HIGXICSUeu2MH1
PW47mxBejqOJRwWeyCee44mVb84OoeV6iG59+Aue9zJrez08hF1CsHzZcXSb2d6olqlYPyb7rdIG
ZnES8RP87TX2pZlZWaxoRDWR5Tkyqq4HlSAbmjgrI6hz81qGMTAWkL4nxJjO4vDFTVfl2F0+W0a5
M4CG2P2QxJ3drICYdAKIAKrjw4K7cdz0BFCX8D6HZsoK4XxY1Vf1VlUAcwYZdhrTJzz1BTBN8tcH
sAbCBs5qwJfpOtuQPL29t+6kIIYHlostAOLach6SPfaNC67GaP/HxgGLRh/pjUV9vLQZO0Qq1Pse
slcS0XQN5nWj7K8w8s/LZWimxMbS8Hjs/FyoSo+oydDD2k5R6WhoHVJTAnk97VCq4RgPvgyGz1+j
Oo7UcqKXnyiVMGUKKTrdDUD7cW4I6g6Bq9qI5Tz7pHvpYaqcFqNb4/hKpYre19ovytKiyY6qMm//
GOBNU9dQmhHe3qb4JgZR1IRMLgQrtkUWrDWtpSDB7dRSKkKDP+YLC4qZBhgAhMAJLEXK3zt1JDDB
9JUdUAHW4AYFbKe5LzQQgw0xOlaEphLWNO1jOup/YxydVQQaeSfB1o9N5oaAhgbg4Yg2WeoH1GPZ
bXCrOOKok3Hn3Ec+89mxszFPesEcNlDqhuqhr8SxZdlZuebVyga5CXgBvbId5TygkMV/cADTzdyb
fRaTJHBCBXFnzG92DegHiRa2GOyoI0pCft4ZjHsVsSxrvhF2RugrtyaTeMgGqHVHPd940y2yJ9MA
X4lO54SvdmRUzDaB4iszPazOKQSwcuctGIcOik8v2QLy919UAgiazsceWXc+if9pgiGNqIotJfzG
8QGUyWIO0M+lBj09cW8az0W3didKiluBEY3XqdS8pnFiWvLbDzDCi1ReViT+El1ZGfgw+xwX7WIb
Nr9sN1+9fKblG3aIfqeRwc5fdI2JMUw+NdrxQRy7Lb7vuMZa7oMMYZeZUiF7wpjns20l9MJsXdVV
AkJYHXMxJBj4mL2/PJxBK40XlvEGHrb0AmE5R04OTVV0BLEYnaVksutir29yVdTQWkvB7fe6X3Pu
UK7EhdCDj485W98GJEjprikUFTdwABVkNnqBQ+LuGvdSzdiUFkS3E9hpTwJvjJRoHM1dHqF6Offp
TlvbvJwkehWpMilzqJvAejnqZzlJGwwCtxe5fNXTIg35EZnzyl5rlwkYieLouWULX9nHRC3UWnTV
snxiJeZL/OY5Em/XVdaXGPetlBxRKD9qXHhOey/wFq5hcTXOK5feHygncZvMfOsTi+qK6ctl0Ej/
BlQj3vSFQsbRWKHIFFOUe6kvXI/kVP1EB7rlvo5h3dNEa+GBHbOkxFUOxtdTlfcLGP8cxI2HMY5H
33J/N87MXr5dOFYNdp26BV3i+qeP31ORjQ55BgVFa9ZEqJg5MXwNe18UOX/JKCtGyGbggl9kyZHy
7vhOsSilFj7x6W4NbAA+bAdbvHfva9Ridv9BF01b/9vRy3DKktHr+AVRA67gbfY/Zpy7hfWLJZBi
wqIlwz4OdXx4iq/G4dMc9++lqkjrBSO8WXIz/MToqY6+YK4Ri5Pvcaw8Ks9bzokugq/BcVtZrSvf
iNf9LEsqdda6mmVChGJiJ77DKpEuwxq/KhVZaJaigZ2k66LNZqYLb9DLKtfWm7V7icS7GK4au6lP
O3L35VKzhiB0pbZMVeQEP+FYi0AFPh97BquQR66fIyLGcUlyoYT87YH5zLEJXq+E+AmRzFA7QOlL
57ZoW0V8XxXlDATtODT9Z/4/CsCrvsg83NxzKdXVU6IyJwJQMrVUC0XM0w3G+QDhQ8wBSdEUhYCx
SlYj0GiWimrHgGZA4oN+oewqgMPKYtcbbrRbNltzbZTJHf+hAMLTxeJK+nnErvOdWj6iYofc+V9z
6F5KwsjIpO9YRMpwk+UJnWGN9y+5F23EHpVahGc2WOl5qkst1yWn0L323zx3LCGogeEG0iPsWoRK
zynrl9TzSo03+sdqsZ47c1QZIhJVTafAh7iqOi8S23dwAHWyvmcqErkA6doX4/uJyBVMFhA28SmE
Z4NSHgM/+ydaD/H4tmcdH8Fc2dHooedPbrDYQt36QD7pnahIDTAwRm/FBwoddhCAAR5qmOlxKxt+
3zNcb3kE5K2jFY/Jo/UY2CxvdJZ5NRx7HmgbNy3vN7KG//mKfRspelsJRpS+4+TAY/xQ/42m49/a
Peaa6J8cDqZhsGb2GD1ma0HbX34azqfrV4s7CELxrSQRyuM0y6EV2H00deGu/jMEke1wrYCxuEpb
zGY7xjzjIOdjwQtLLLITIBRU36iUEfPu8E78ncQ4Ec68zX8uaMkLLzA4LS72qPiP+2vGy7CYogjg
Fu3QGa0jBf+YtGcSck0VgrQ85FVg/jceGaZwPzImgMVCPgWXJLZ7lC4W+hzLvQA2PXi8pD0Z1DZz
QmbLqxC1d1tQXCF9OVMWIhwMmoAsGLlHNYLiZdLc4ip4VBVs6E/FFjJ9XtoY6hxy8tUW9/IpmgFp
iCJZW1n0xcP+banye1RXtFVQ3+VLeXR+90IxViVFmJjN/XcnaAwQZuKxzRd+ZEvkM/mzQGIP60RF
K2Y/un+V9ESzWO+DGsEFU5f1raBb11uYW46dA7xSLB63XFmPhk3VgtYCl4aodvFI+kbdimfNVf0E
TWVi5wVMWc3/u6ZTku+5ZlMYal4nRuSj04xRPz6cjrRHb1iZSv+pcxVGq+yaB9A2OYwb1kaf+2SM
Fp0Uv8h0oWxGfGnzBLNwLHd2mMYgZXG8j3S+Ls9k5H6Fibd8pvEmKlShtgoFJc9Bw10Ur3kw2NOc
SsoMamlDeYX1fteOuhTLuJTvVMBMfTwLx/CzNQnWGkJoeVRwZlKt3a+L8tkd8rkn3wwPbG0mFA2y
4RFxDjs0/HvzVqzy0VdVIunSPtnpl3b0cqWqCVQ7Rt8us+hDv8DyohlYAYUQ2GBO4Dsb+y0Tr4Fv
bIZDG6hvmLzjfDB+SXxIHVbnQ79xuE1ax+JavgBTdrYakm/mN7vMRi6OnZYFqrA6FnGMBdb1bmzY
cklnKe1sBRwDRjizdfvOaj3gdHQI6SDf7l2lCLV3P7EoZJixIBzoY5j5IQXPtcht5VJSCB1sYqh2
i6tHEn8suSTUadPAjziohnOghU682xaPtS/UBudLZOpoF20UFiatM4r/up3DKDUiCU/SqvL5bmDu
jrvFT9fNFX+wfed2y+ldD9GGlsAJ8aBb4WjVpo000Y/WMyxhgRsU28lyYIp0akA+Mz1lkGmnZ+Hb
aHSt2MgODqpCJ/ii+8aYvg9EK+j5Af9rkpD89S8AUNpWRRXhhS7lBnVZDrIbpoAdugLrgiDE28S/
sQtO8yUeObbPu9hFUp08wQOyu41LLTvf9VY4oM6Ul9a8xRhiehnNyyhNOID64BYwmcHIzjwNkuWf
MEATj2iYoumYFcfhz8cS+aoInQjCAPCeO7psp10WnCj5rjU1aCOHk93NHCj7AuWM5I9kapAdfYIU
FBsKGsY+W0N1rVdhvm/npU+vD98LN9nZOB2K29zVAS7dd2Zxsg7CwHtVkf1Bx4Ym7EByV7Lav5Tz
kPAZAEr1idzE1QvRoL+7hNs1BsImAMl/UcE437GTSGxjChDDSdRCrtIDt/mXm9dgw4VVKJm2eTQb
Qaly5x/7sYxc0HwOuqzbJ7uUabgtQnbJpwSfDJZ/dr+ItEYIw3QHt4afro7Wd6jRv1gVikGr5nuj
uaO/9cE2OJ6oISXvjpLvmTDGS1h6MH0SpJfFUwBKVBGe57WRDz7nfpKjb7BjP36M2iJuevVHxbA6
cRTsZuz42IKdyUsIoEbnQe6UKgkg5L5fVwGuu484VC+L3lWrfPEHgpK13/j7DIGQEGYF5JipKymb
8skX+RCi5Woy2WS7EnI/uJHfhjyykJL2NZo1EcedShIRjyxK4+9CnHtRwqUf4s6auzWELHQ2WgqZ
EpEdWK2682rBBEGJLSUsEjYTNZ18QUjdIrU7STlsjCRbLqO1tv3RaBTxIBpRuXhJM8lePMOeNEJF
fqGVtGbFqIvBUSof4ElDj/j2aBBgZDdu4OWOcZuGFI/l/zdKxdqKTrsf6oEdvA1UFBWdEyv7glow
r0o1yPmVRN/jlJLBRf8LSZ1mV82OzJW9StsYGfE85XBqnr1aqxaH/xwJ0yukfCpEwIGFYIH6Czcd
YadRrP81R0HnDo0UKOTU2YLHCybz1rxraWZIN4qNHmTGoAN1gFWIbMVGvApYRGOX51wBZYHrVA/j
lKgVvln9nwvdwTaHCNYQEEXT+Afi1OOfzkWSuBPXX0A+lzXg5BUVUXiIasl/dMVjdP/Mnxzd5VBr
Zm40ua0wA1bD60D1Ae3ISWSYULOr/CAi+IqWRRcIhxRVknXdBFe/evzbbZhigWKlKFwAzrp+blin
gB0Xrmg1288kTOG0/EwAOCPgKCzsdXs5DmLcbfDwf+rRfQyJ9RGoGD6qhGQm3FUszLJkgQVNM45p
shSad8omb888ejqHWBzScnCSPBmkeYnsDIfIMOH0HYlJ733nZ8w+Niucz6bBe+Ki1WY2rMJ/6JEv
dT/jMyckNSOfzR/VbUlXkDbqef620YrkN3fLrrwg6sh3081n+QCZu9MB/jZWc/6hMr/ggcUgGLgO
FBrMuKT0yU9++6lxCjY7Fzp6yp2njeh3ZlUDKpOBeyHPw4VoeyXZNAUmf0CWCSoUZJm7xE8iJD1Y
XUgmToMygxx/TxBYK9xGKJDs+99TQXwyX6I6kUkTp6bz79t/5auyHG30Rw/HmJ5TfD41TfLh/Szd
g1YSJt3SFl+74Csc2TYQlgcCnfZxplAcppD3Dvx9tOkzt78BtTupeyVzDV/q8oTXb1tH0eLDzIv3
5oTp08lfLfU07YEINSjz5UBTJe/bTyTvpbIs9A8599l511022/qbHuxhkdjr2jRI4+KtpvtZ/4y7
+2FsDuuCKTP1xhg19PrfO/5Rs/MbB4O6vMyAPb3LIelxFskC3XwUBPGaBcsCvYbN4riqrYK2P6YO
hL8713+KityvkXXhaEJIXVlTZCyVaRAeUETNMernc0+MFKZLwkWYPsQ1SkxzvcQzJ+IB+QsfWZXZ
X7eEu4x6uy5Xgkus8QZ7BRwqZGAyvuJcLjz9TVH6mu3kYs1wkQSWTCScRmsr9w3x5hmW0hjsWjj2
22vAFFvKkwvW2Sk7FuWEiGRsWg5Bm7+9KvKtFJM+nB17NzjYtIzXgt2aBnv+9O9IOtUuNGZwH6tb
CsoGNn+o7OPXsG48QTu8B3nwlS/2w7IN55OBX+F4dS+zEECU82zEaErtaIY4Wlf98CfLQX0130Fn
aHU+yT54JnwpDFFsZOdGrORM6Y+R2JKZrExnSGkCsIrndwVZkN/7GS7PmAty7cgic91ouuAXUX8i
bZIABSKBFSRG8VKuEixQNHlKOuDJc3t54N8rlVUGCPxoYgrbOPz40vZ2o5tu5g2sR0tfKT3L8Czp
dZLMFwMv4VOdlJO85mxi3n+FppDTZKR2mndLesK6BIrQjeed22YRI3YMCQqiqFtP5dXyb/Wf7gEJ
vYiOuZw5tRK8ps5oDzpQInbiJANbxk9ROqn5FPSyI0uyYUKwPpxoj+eW3sqC3mDVgZ1SHncBw7xD
6/am4Qn+lHtycWq46LZKV2EQKmRp64XHmZv3VOP8wuF2lWRr+L8aNIJWkEQN14+oOE97b97v0eWI
P6c9hBeyMLO2HaJYxfIsV+m83a9G5d5aytt5tSJpyvZsDbMWas1cezM52pgwoNGKUO4CQ95qkc89
hWa9DQ0mhDTsMIsAkFHtw8pqO34DzBtHTDFk0ZYOct9iT04pCl2wvZULwoCF7y/4ibBz2HQ1gf/2
qBlpw2dsXuxXvrwnI+zSKH5IajU+ESInnNAi+HcFYwrWGjl3PCxSUmOEq4iahHKJC9Y3ODKikpi+
TUVCG252Cf+dQiKudWHOTxbhyLnWgUcJWIXM/TQWzFwFYDqf7Lc59L4gUfXDbwDA9rBdo1azX2b7
T6awthHmKy9kltrvSwRJoOsAQg6LDLK7D1T+QCKFjDCJQU5nl5TS0FuEl8RAJV3X1gfOnSc3IIpv
60liUNh9gam+deGchPQl5iasx+Rf5ZYpG2YEpVma05H+VHyR8h++hjyfVyMe/M8fy3z2oXi3eLG7
C7KQzMpleqyK6JCK28dnBrRhPCfR3IBtrHluiV+4ilW6TTuhsxlqmUflZcPT+zAmi250pOKH6UM0
2df1u/xnAZTfDW3eOYWI9L5k6ExSD/Zw3UV8ZGLAhByzCoHtEwzgALRm4b3rqQ+WXagb61Yn3g9X
Vo0TeRtpUblpvfNfpEboALowHII5n9ExziwT3b4iQi13Z1WC2o+fBzgQCB7kYhmelqDgHWVwrfio
5w1dKKvPo9XfesglzigUB9JmuvI9WhncDu8sosyEWhaT17gp6gztgznowLNEZN4Rxd0avYi6SkaW
dihQI3hhMSVnIH7guV1urgp1VtdIUpLVD4fN/7XW1N+Sy06jFoHzv3yl/n1Mmy8AGh3l8TF5DViv
fiEM2h7Ffek26+ri6LJeHThm92uvQ7i3XM6cTiA32R9iZC3L19AsAremhlU4663Oo6KS/Onzn5li
Z5MPHNCvYdmAxsWjTV9Os0qiTHaEUcpbEgQcXcDqkkZKd9p6Frj6bqiFCfRHyfickgKDGtw5sKYh
7lrk+tLn9im94cYQW+k5wKHOfz3Noky8r0TTCJMKjEXDw0Mg4F6jRIqZKYtze6fbogFbBNawyYDN
ckar2wSLfyLBflcy48FS+KmDpQfJiuCfanPeOCn9xxPDBHWPocgoszZrJ4TobCfKoROx4mvLx9BE
jTSJsozquWPpt/5sjRaIlVr6SfprsWepKk2+A/El/oQ15O8kgnWecU9JmAwQjGHoOCM5wqGG7sdn
jst3Q8qust67aBK1rHOEfyc5H8gSwr3paavWOs1s7VidyNR3tzF4HPFKcNoFXRvGdJi3HANsN7Je
vZ9ythtN1yY+vyXJFyFEGuB3DhRmlmAHYSP57EEy1AWhGgnjsGbmjrqxmrdNQIrAeeao+nkTpg/E
t8CGRvYZVzxfFCb1jBod275XJ8bKsu1fwoBzRLFZeFxeOoKYJlzWlb0UnoJHBazbOLpkk3shdZFg
Hw2p5/5KiAA0KPRUGQ4muxbrHdpAVkRmgEeUJeCzIjRAtdVIT1Qz9AHhSxgxKARNXAaxtgoGprSc
LD2Q/hJ3+/w0cuR2GTYbDIHNp4Z/uaqJr54FFkfT16Cn/BSUUv1udSFVKdeOQv84meLAfxAH6pq4
9rwNmZJNpaBm7Mm5lXruGIT1fxz7qPttx3/SgPrkc6yMvnRXtJMvTWN3aJQPiDYlG4tT2BfOFTX7
wt1rIqkmRs+biVqFYJ29vqKgL3DtWyWkbLX4u3/QNz1f53CXc6USHEqIFJxgYg/GV1djCI26m9Oq
xlrr/r6qlw2rBTF6oqxr99aLxElbguwYrKYg8wnskwDIAwCH5j2z6SC2TNXmV86OOvoChVlIC/CH
d8mvkce3gxbBQu9HYss+TYCIDsHjO1pE2HJOdO2CX0xhj64FVTmG/CNJpd8YEXd06UiPRJXgb4ZM
IMPrJ1nRJU1CFqs0XAF18s8f57U4bEY8zUUN61WhduBDPDgW+1RD0J8ZrLj8zXRjKnT9jHSi4/bl
1IUvWb4bGEAQHm2MHREfPYVrdKo6PKJ3aVwK6NG02Iw6e1no1luU0k5d8IM9K8StCm3eKyi37ykC
7AToepemPDCo2dEZ92pBkxS1cbrrwpL1OiRj7VDBdZ//XuukAHqXMfhmKVhpPm5LyDy+nhBRS382
VaubvLyB6CuYLJno0wtlzLILr3ebclIUE2vvNIIU3SaRxvjyq1p/cLPYIUDP2pdaA6SgCtuCF1MR
d7r4mXmjiPe7GV+eVLepsLdiseOFSyvvzI9fWQxqoO+cCNi6JT+N4K2gGAXGK+e+4MtOBNCU8dQD
SEnBhr4pwam3hOevn0aQimmihRpjs5GmvPfkl9xkZoxNXzHxhCw0O16dkL24Fw/1tQIO8thShP/S
CIHE9i8EBQapYxwoSCTW0VD5sXpykUJK16VlOrMVlEPwkOuPkIF0EcHTILDIHYhdNPhDxL5GfHy1
kjPMf4T3V0rACt4yjE+63A3ylksBCCG2j8v1ta/sV/HxoWTgoBt0d1KFi7HYFnzhRryng2ckVexY
i+0rwPEdtwVq6S5k1NQF+tOLuHWcKQrTYLN2tP+WViPsy6B8cYHkKt9TBTYfEl0+ZDch5kzDqsxy
Rz48dfvZMU6+mBFOA1zmklsMt6vXBLB7rBVCR6l/vCkUSzcKwC1fKNO0MG5Xy70qn/1P82QNkr3V
Cy2LtMpNBGkM55bFyFOpa1N9ZpeHwDNbyLguT5cakHC/jWAe3Pv4JuZDxK5V4FQ6uEQTYRN5mfwb
Wz/F1USi0SHghtXnnR4BNwkoHIKesf4AMpl/GRNhL//zIDBallf2E/u5xMTl76lL+3VZqn2GKM6A
l7omxCt296rv3xMQbNE/hjG8UXjxeQDKyXM1qOvAaCWdThkW22xNfkBBfPMTXvCZSNoELwCumoxE
Yk1f0U4NvCiYQtWtn2S8fOkWnkYIKlRwdiRMUjF9vsqV0hyE4BRSwlNfRzeNfwMga57Ss2qnoS3f
gci/JggNqS/raV4+ZRISO3D45ztX6BbKzuSTEu5Wcf4gFGTJhdCOWQzp4GJcgo3yfe/0mDrV6Jtn
oZULnqNG9S9KtCl1Kpesa2GmKk/hKn3/WXhNCCPCaJH9RPhygZpgwV5sYg8+0vcqJjBml+OlTfg1
xsemDZZY8wteUZYP+Q2NrHvkmMUtgNGFeM12Q9bkQuGj14J+cS4BWCBFLMYzmBh2QHmua8WDZGAi
LFFNTsfa04hzUYQXH4rsZDWq+9ABBKREm4O9Rk26Tm4RKfOC4GVwwp1H+0RAWYKJXzxNyMIkMhXl
ZtlaV8EFQKDQoejKj71vku36/7BV6qZPTKBUEA0bvSZwZAJfUa3gf9gBa/sk9i5oY53LkMeuCKG7
pF0p4JJhFYNc7nZWr+54JHOqEQwmgxOVcztoVmbhjYABjkB8eIyDOsRBvU1G6Pbh66iJdSz/rYQj
M3P39HTwZOIX1CXQdDL4mD0Jelus86E9JZvla7e1/OyHcqbaVjq0r8vvK6DpmmX/1EZrn8A+d+D3
3Ajcpu19rtvYYkLnDExS4D4OQVZUZqSEzFDt4KHMoC9fV0p+7UKu7v4bSNh580XBIb9D72rwIb5e
+aJ5LKYIcLm6/94zcGylEWNSpVUgSYWUMyCjJzEYcW9Iuczsm2vQt6KvMUtd4ond8EGGPpG0XK0N
h9qZm2xRpK+bhXEByIXxkEIw2Ot9ZzkLrV+ljTyOqL9taChxmsz0/xGANFFYuTsmi8fdldFNVf8k
6zduGwe/ojvmrrP9Yvg+Okyva7e2zor2IRFuM7eWYuK1MsnmIn1z3x1PYoIdmCTbldORAwLcuG6E
ATK9FWrsVDbMJPcUcRAl4c4MiL5YISlR/AtHMiTDNgD/jt8Xc/Lgu0ouVa2tnujHjy7x1RKmyWi+
xiSc7A48jLTedo6Tl6X7hFogCsEopAwwJGDRn+l7hyLumeqwGD7Z4eIfivF7m8yYCIKPLLfYw7nc
z0D+rZDPmRkSas+JsbQ+R0fNpVjsVi34TJ1AWoGlbkuaYiox0ozQVmRoxlxYpdK1pTQ8JdMsweDX
RTfbSPkdgSM5gRf5uy62qUnd0iLvjhnKFykp4IxqFO+KQPiSn2H9aDpt73eAFx/vR6ECkqN3NYiO
bl6hg0M8kmatFjpgE6kLbbG1i9g9VDGnbDHGg2vp01NqfyEpjdlBeVLOwE9bKnGCTlXaPmFYeUJZ
yeUXHGyX/hjsGjEeE0BQCkqmdSLd73c+Lm7O0fL5K8YikXgMpnCU4ZSMtIGeejJf0yD776jY1E3/
ozilKrCW1OSwucJ9OMVA2KcPnMMA61L+6jeQ6SJ15bI5AM66UuPfKygBIFH28x0HwE+1/tUCvQ6H
x/Y4rcyQ1J9UMy84o+0EaTzdNoyi/5UzVCtWarDPE6eqN8gxsLaNcRNPFFWBDfUIlLCFmK6OLhQI
IOpBI/gvdnWbj2/rKYLouhZk/qC4bQIuDblKnzId/rCX2gVOV2ulerpQM5EWa6lYVzPvGDmoC+8c
9HWc7TcCci44AHfQSHDti4H8xdbwZlo8rqHpKHqtQp9PGJQE7N3vW3uekGMEhSjYCi6Qmn4MO3+O
sw5QpUH4d7vJ5k5sdLT/meN4Iq8eCwTrqyA4NDaloJRrob27Alcqb3h47b6yLGYH/Phi9qMNJuoH
+fRJ1N9/gK2FhQ424xhjwwER6p+HOFtDWWse0negwmnym3JDabeDZMl9ZvV0Y0OcqFIHX9Y29vKn
JUK7kAv063JWAcWbVWNLCpSKD2OemVxuKy5LjbWnB4b4D7WqtPaEK8E2zIs9LY3QeQ9nHg2uslS4
NX4im3tNn+l5xEITK0ddY5DZ+eJQoAvSqELQUC8UW0+IwYoX7f8k3GfGZ6hCC98lCqunYJGtjf+m
RV/fAF2Wa6qHdsDVRSyrwV8Cu7hqtMTSaCnX4hq1Caohh+ocVYYMvtB9GGPSEZJzqgyW7so7zAK7
2AA2FmU1jXxuS54K42u5U8peVUZIMQLdZ2/1NtzXRLF7SOTb3Ipj5hXDHYA7eLmP/Bg02WayWnJL
8AumCCc+zgTq8pO8NDTvrzQy77YSQ7ReTJKzv0ERP3eLTNEIJahRYQ3fMBRybd9OiGKHW9+ZTtW2
d5PtONS3MwXg7sMetQUF/2mKb/WFigDEQNKj/6OAeZoo1r/oqzg0q0/JrMtGVEZFm9XcQPLAS6p/
RMtVf4iAmoAq4Xt0cR1n7x+3t2eByeZfU9NhMgEuKsrf+K+5pZa1oh44VFhLji0na0D58VDc5+Qv
HdVs9XJy/ub42niAMz+wJ+Z0FKmZqUw9E9uQLnm95+l3S6BM/JMqrRCLzU02M8SeBjSC3T3aYt7d
rGSSdakkontzItwoebLy09YA/2lKrnHxSu4ZjY401nGS1i9asyytQ61PXGuqOqQugJXtjiplZLeq
6T2zXr/WmyCNQreUfh5pIfaSSV2Q739ECC5AHfaTYJcdehrrUCEleOigX3h8e4eNg/J0qUaR6lha
pizaOQG58QfV6Mho8kIp9N0J7yZYp0JaJzwq3m7P4VSathGximSyZKlzBJVFTrQGO8ZKUiaqk776
L2k6K7iZfkNfZmlY1FSu3fZ/QJwQiK5Pl0WnmbRgfudjJZO2AQyAEYjLrJ/2e2nAMLs9RGrP4OJx
8OVCJy//LXr4PM2ARm1h3F3Tjj/uW9fNqvrMPFG5M+S3zGB0hoXWuM1BoYxYaShgALYMHNMnYrvR
MdSU8EmN1bi4z/AgpLDIN1PhNq4aS9yNIMkh7WBNZQXR6zA6P0qkLNKy38/nHqjnqV4n3Vs0/gpT
qsWhwDXcog7eHLltfFm170SWpOhnOGlAs4jM9EZkNf+9pqmoIXplISQEydnTYLiP1UzydPNCVm+R
0CCC9sAnkWJUqA+6HHmOqDith+CY5oJSXWR7jW2Yn1D2CqUgqli6NqHMD4vBky8I1ujg5pCAPd3E
doKFfph+TtX+Ij70ZTUVjCiRdKyIcuFLMVZxNNGHGk7JaFMKROt4ZhEcm3p5vIOvzeHhT+Py0kwr
nwxLb+haxKq7TkwsvCq7T0ZfMrPv9f+F3gT0Tp/0gDVwHE+b6WuSL6FoKFwxZp/zeGGYlZ+jvZ+y
2n5dTFmrqY6CDyYvykdt1MbtLF+8kT1Y/wuBDf8AGQ1VHUesM0V6lZGHBw4TtPLPbl67N/rmvHrw
K5TpN/Rtmr4OsTwpJoKSc0/P/2KhDLgOUjE3Aj1drM5vhbVoakNndcq8MhT+IpglV34b+UTEX7s1
v9SKv1npZp8HrziUSrEvZhbK0D7e+acXK6NxtDYvWJBAzN2E/S/rwgpHY5hxv6Ekt2/3OA6pq1m4
BJmCbh5i5pvCceEo5iKVjGJtScTT1s+KPp1OLRuvtmA1C3xdLDBX1Fhkns/VuY6zcL9YLBiX3KMB
4rw5aDZDw5CfWqpp3ThXJycCBil41KbDmy8lqBFw4VND83EPH7HYe4dG5XORaKNRd5pBKcBX/oPX
+IAVmTYCjmVz4LvZ7rsFw3WDOiNwjKqJkjBmhQLUQw6V59xI72npn5K72cBLVrJBFIV8Pr4t3v9X
lqSK0+hZ44AcUhyzblxIC4iAaXKlf2NImmjbhHIw1iezvn64p/6oTr1K3XJZL+DGyNDN9QNXypzr
SshkdGA9FyRlhufsWudyB0ro7A+YZBuWw/PUHG0zcXs0SRn+btrLYRlk6TOFYsBwZf2VTwsEjBqf
9MStjcZ00DaXTHVLqNTMoAzvaXLZm0Ftwr8MlHXlfmVot0cs8MpU9hh1JiiYqcLcG1ck6Wym25iD
kQJPzIyLlbATf5/r+xyfIYrRUh2ZwICiW1pkFsqVMcAF21Ylq33GMPfUS4r1yMlUDtEy15Wvd7o4
hZNoGsRCVPCnliFTFWWyGNJeXs0n92eYDVtf0+VypOr7E3R0Tt7PkpthpmV9NOcTrMMY0Pq6aGik
rMLElO2qLJnt/GUn3npXf0Rcg/rrv+ZOsLmDWLpSKPtWj+btklCCTVbbkmNtbueLl0G0eNIEGw+Q
rrBYZYuynK0xnEX53Ye03jh92LE8MtYR2f0v0NOvrBubXjVnEv0AvPe74kJgS4/87GPMBtz9y9Qw
62T2avgDcwVfQ4N9z00RQeZ3Vr5tos0BZCeApE9gOoGIycEsG1G0jIoaYhSUBoYKA9n4SwNMAhbe
X4zuZDD2mXld/9y5uy4+k/d5dX/GUZcTXyoDPJk1GooajPf2istgG8UN+3JCiIbRrkoOwzOBne/V
s6JlWy5d9pJO/jowUW4hClhtO+K95st0Cxa7Vr2Buw5k2ruEYIP7YmqyKHvmLLNSHGJstoxKzVan
iZ+hgpJjMXDReeNeTQBU9hWO6cC60ZX3AJxfow7GGa86MEIniKFr3lg5rf+FEIbXp87AqIjYyWwo
6CYZxRO1LU9QVk6bb6cOtcLUJm9tUXk1YgKzwlcCWNVgSSql0EZEhUivu28YptUduw31kBfDZvXd
Xzb6NYZngzzV4Q+Al/nXJYNYVwk5wLo8PnahVKrY1hJ0+yl3EEmAau0lY7RIqLD/A5OnIqfLh/eu
sHG/uSr5mKvwgS/59mVKFSY2eobkgTInqxHkr8cWVwg6CqdtOMH6YjQrMomsqMB+4onBUbKZ0X6v
mSnqsPF6sEGgKbF1eP1y5B1yVv2ePk6lKfmjnXfsvCZoJXNji0NlZ57p+yBd7xmCtqsdTC890+J2
BoBNYpwPr2RKQ0IAPmy18EKsFl458941wJ8b0ghw9WYxfljJRqpeSrxSuwvjPdIw4jCrPqgsb1R5
3xay29TA40uUmLye5L7VWFwYbyLcqzx8/E+5HaEX86uj5/vvqQYAcNW2TZ1p6RYgy8QOoNkZu+65
eMeqzkibciZdcK72ZqFKDGwGhpAEtRivN13LlgwkMQDr5iN+RNPrfOSlMrBJu1hEf4kIY+aIPnOh
EwP97Bkumwd6PLVGrWXCuC9jLSqy2b/skWyfEqXAdzISyfZwSjtlAL+C8eV+TYBqqDPCOk3nQMwj
iKbh+7I/a1XtJzYJ/KL3Nc44fLxyyfBFUSqrDBBIp0r7ZoRoHnmwtZ53Ba0KdlO1HeLtHZxRhx+z
RAeMCG1229qlg/xOqTZ3xTap6P5MAjWt/YWrl1aY7SL8HpEC9TtJd69qU1S8FvM05Q1fyCz/HIeA
7tDL7mmAjkwg3/S4p8wtru9Bur7Qa8MosAmRjSTNEz0wdG/KciUZCSO1NhFfhzEFO08A02JoONFR
2DLr7WENBe7wZjKLul2ZcbMSdwL/VP2IuZISHlt9WYtwUUHXV2Z6VKDBUIR5cXgrIVEvxesoDKGn
7mHtLN5Krgrfv0Sggp8tMxKltNkj92zwT8yf2Ggn9nWZDHxpAvt726Gssn6m3Ld+m5Z/jfTDTj/C
K/ZWFPoghL6kW+ZoFDJnTQLEM8LWqO4Xy1I6mIMXVWqFnNeBhCxZdRdWS3srYeYN3qdMg2fC/0/k
9dxXEeDoxSPrb/c6lKbyyGzJs+4BC1U8tP/c1l0TGaasEvBvHr77RDOORjLhH4LZR8adAp0Pt7jW
Yd0zU0omxlMrsBsd8fAafPFNe9rOP2aZE98tCps/0gV497NEVkdOPyEoBf44aGNCrYEHOoNP35Sq
ry6qpvE5HmstcD/CkftvlooOCejWOZkHgyCbm6MHD3IgAR2VHF7mTPyftTwb09AHxP60cRF4oW7h
jQX5FJe5qc4rtLSwRKqLsOUNF4PdhWP6mmHxFZoymKF7Z/wc0Tzj0vYjKa2IX+uTf4y5eUrim2GC
B7c5jVFXc0GARuPgiTHIS6BrqKSPzdTgw64dfv0F/RuzbH+6kk3kANfeaba0RiFRuD6ls+8oaSrW
cNYO+Wj+Pz2noi048aDzb5QtDc8xiSFS4GEEoVXhcMZcE1LwrfLQZXKo5fdlX1xR3kqAEciW1Oj1
2OGgNfBLBIOqqlhk99juEFqLEAcKscAXMAEDDi+bi8lWh9BONvX7tAfpLDN06zFqW5cdRD2umkdw
5S09vwvEbbV0QAwfaj2pzk/UblFh9nYt9sYdFiiLoaHk/Wf33omCx1qIMV7sTlnonMXvbMqiljMo
hi+KSMgvDOeg+4yAKM2FnjGRSbX5NVCTyVLWXEHWs6gB1PzzPdie7P6eVf9gVbrUS7XJ2/2c/rvu
dLK7FQT7EXAA7hMyBUipOIJbZD9ZdwNpCCdfx5x397t/zcUR83tuiwTCSInIxXkE/olNikWhkVTz
E0wGd/MsYF/U/8/YrFvddYr9IPzIsp7xQ4qolX1xYSKYGE/9nZhUgUpRtDT7faz59Rey181EfDSX
iWod5e8K6l8aUcDLeU+BfjS3kPI2eqmJ/WNt62Cu+zc0mJSDyzikV9vRmIk3Zg7HA5+yz81d4nnA
Qfir7xzY4CKhaUko+rK+GH2ecLtR+dexlmQlzxQhb1Fas8kD3oHEQqtsdyJk0kTzK+y+LS230yP8
OzPrxc851seOaA16ZSbXu5MoZv6aIiIRatVroX8jYh9ztQ0lW/Qnq+OEoKbULkkRv1XqBaQu/eCI
heV1+Jhg0qKYcT8UTutVtPkybORm1EdlM/jB2adfK42LejfjymLqc3oXaQoMqNGjxFw9j9lfZYCk
0IjAnhAhjAz6TcbwzPxbafqxzpkRvoWaBZidBYU0/Tf9K3r2Q9X2sRsqZCAe2Ea6McJLVzwkzNuD
2U3+311qpTxcOBAJ9YP7OQKcDa7Ne8KcsG5DTlcPPYeWof3RNcKDpmATN7Gek1rM7izdwBH1V3eA
sXp1CyZNwsCIclHIVrHLMgEHQYlOoNBNKvKqqblLXQziksuz6FMM4AYeFU8jC2DMmkSlhq8ZcVhz
7nA+CjfHOkJE7n61BV6lF3coUq+qnhLKcmxdWN3SHc5gpCD8Qz7Epjk8jEI0+UTgC9LaG1Nputi3
UZK7PL2CmEJQH2dDizsaUrI9sMfJgEbXuFJ5DMgEYmu6rqtHyXzN/WAxTS5iEVNRP3L9kd6manCX
08WnNXtCWFGxi6CqYsyL/ziDYsCHLgzEDllxL4fFeQUUR1vgxEETy18bLeQOx88Qc2YI54biK1gR
h0f9k2oIkFNeBgXMI2FaUInyFkX/mGw0BAmf4zZPQgmT7ZlQXZL9WK/7lbxTUANR0tjNVkyyDhRF
3mdEhoA2Unudcv5zhnGl74IaxNOaWJBBepORAgKU3u0nK3B6WvoCDpBHF50K7w3QaxxzFDhouhfJ
2hYab+v1+nFyLdzSQcyTIc8u0sDQaHAXqEn8TAuopKpkDScHQmfgUhgGq5EHJgySf6BGJOqVBJpi
K/xcG3DD1dkZv4mHhCMRiTOqM+T9TnDPSpSmzBHcSFCaeAk5vvc0MbiECmqVZkIybsZdVcnki0Ck
gImYimy5lPVNXxYMV7/YxkqlMAHtNrkmTmCWfUUsQiLdmhCXByimWX0wtlxWY0zeYhfQTPWWX9vj
gFf7uKL0JfR271TGMFbkDkOKBfF7YaZtUu+rnu5djcpTWBHmTVrpdnWbYSmkUbVJ5OPYKY5a4Mrx
P3IGLQVwiHAFjjf7cc2dVMi3N+DKllV6+vOknR5E4rWHoUNijMmT4yCaopY4gDbty5vp59xx/k+c
EyNJfU4mSsDnlUklNGMb8YwiKnYDXmJsbFtsME6+NkHba20UCTsPD0xle23fcOGn8SwKpJzV0lzb
TtWM2JaumbNAthXQpVI7QHPNQCC8QzraZXSEuwetEG1qwK6JBdnGpbzvmDwd3UOXalxDUJCD6Qho
cPJUCgiKP3EiV57GNfL1urrhR3aGeFIfL7PteKvthI8J273BlIx4VIjvphXo/unWaDecmaT3500/
oJOH2PUr5R9Qb+Oc0V3lx/GNdBuGD064y76z7MF+uLTyVyc/GfX9y+xAtnpfmTuJImEWRuo8k5VD
3eHMMgHtjm6oOq3jHBtxwQp6L5mf+Xcc8r/Sp5xcX7ChxQ3qZQh9l4Z7JCgn9nTfq4+3nAZXqMe9
JyfP9BV6cklKw9HLZ22yLmtx+8XSIxzjn7tXykskVL8eIvjczpRabqUGJsHgEC/aXwq3+tTmCQD+
qpJYWGujEkL2eiLqrdzX1ABV8j7yh3wgWZ50hgYWGjzrAOFlrz34/r0FKN9uyV0USrpyFp5WNWF5
WFL7AGfhYqGALyPOgREW6+J3+jTiQvBxYRAuz0fPiZ/1SsvBqtanpB0AiCJ+JTaCwtWp7wDee93R
oGFtaN1rSv+a2LEzll5ADFyOfWmo/yoVj5Si+hRwfOp8S5IzJXD2RcHR974U9Z9f7HAGHaVzpS2k
rTcx4rH3TBc8do3zfW/4IYeokJa2tcwHQwVGf9Gg2AerMuqvKgraTNV9obFQMKBH/P9F8u4joOfh
Y6AGHvEyCvGKcSbfHXYlupJnWfyFttdSX1d6tphINJYFegpZT3J26LpkBbqkgsopmWi4TAdGjTaO
c9M9uVysQdX2RLWSWC0tLkp1CMf0bNsaoAO8Q0JOJKhotj9mcMUcYPCsIwRS/8gYzak+DFa0mfaS
BBfL7k8us0bwnjNXN4aBmpvK0/nwjQTm6TD/LNmKCyaY9dPWo6Q0CJIJ0wEPAAY0L9o0kZvH0W1v
Eibs9BeqoMP/CeT019ZiuLq+A6SE9BGcu7uo9xtxxNsIn9ILSTOVcZ9JrggXEpvwOgR3ol60UZcW
kG0I/xvKCqyCdCVv2lR06p/JCEvUBgjBB2TTMVI2XDFbu8pX5Dy35FFa1V9yp0H1WFBbcGS7YI9Z
F5W9DSNSXnAyNNFDFjIJu+NUyUwHiagyV3F/KPAT1ZLZiF7CZ9AZ7bGvwe0lzHrGMQy0T3EGBSOO
JIaUQhmmg5g07/uTiHrf1FRh6F3UzvVFaCnJly/8jiDbWF03MVbz5EMSwjTUo1hBsHjvso1lsWfR
rG3VVzISSygukG7S7aBQ2CdviI2dENrVpxnj4W1EJ5wbhFsd/8GLJ4HJj9i0rMb1jw4P/XbSGx2o
7hDvUd5XNkPEK99rVczx6hX7/Ep88Bx7khZsmP6HuZ2g/eEjgqw4nLzJEWaloIoqiwrcm9MzHEIE
9bxVuQpcCji84BTvEGlXFNaFxqXHYpiXGFIa63Ghu7JKzTflmRShVQ7ohnLP3WAzWk6lU/SF/u6L
snV1UQaItei0XosfFqru+UNUicHgJEN/fXFK9wtPsSW1YUd4hOnVEU/s9sRztcs3t2vWryBk1tH3
JKajfuZJ10j5MAK6a+5nRkNh+mEhKB+UznTPzui52D1ITl1Zi9CaV6nnG+ZP7puAkKKIHH4PWXFC
UHmelEzmUSTTeM0BWCzwgySLsYjQrfPcvkWkZIwlLce+QcaMDe5n2YSFc1f5/ii9khD2F1MraHfD
CHy3/iEadq8ACie15R2molBeoO16NccGXNhgtBJXYS9Az7viJxyLwXZEofancm0iB7kMcSwjOa/h
iKStRpRUyUegwEggiNGzoc/OoLjvGAo8eDzTJmFR9Ou8lXE4HFStUcUP07FfmpZNAEWHEeRiX4xH
njw6Vec8WVlS6ZDzrSFifY10a9BtKbmhlTqc69wwYpCbAnEs7HrFblLUufrJ5QZUHJgO9YDHnwKV
aSEbYsPVvZhoxRWo4CVHLIkQRSWlVq34Uldoxi6UoQyTuwvzIRktnpa08rqk4T2h4CSIG+SI74jp
zI8xuP0ZOC/Hpc+bU2VsTVld6Fx0aiMt9gvmS7HAGsSnPycLQ7g/7jMEnzYDgqd7pRK+Q63c5DuU
nxmw/OubDvcPnwhlksZO4pmmXYjT2tZScO27ovczrXku3fMZek2Pn5yr8iSoYFfe/E7MNOEja5C3
QlKWX1YuyFnXYtzQmv9d9lUlmRfNjTfVxbXVi1JqM2aERQezudsy+qtQrTYtcpK5TaV8Lo8DHQ3A
rrqLrA2ekLSrrsch1rckHAXdkVFDoKsseFgpKvOANlWisiYiG9k1uKPwuJf6naSwF/qdDAE7lxOy
9PlDuFBlpGzJhqP0wuTTVhGH+UreWGlQqzKX8dBwLLgAxpViFFBYFVg4mrvHkxt2QjTQdTF4vnYx
3RusZB7vxngPuPD7vdoFCcD/RTrnb6QdDiMgSmlSdcw1XC/7X08pvtNSs6epZxH6BSGlqUGQeGHC
lizId15xrUqKlmYDZGb2S0B3kkeBk4pFmGM2gaQzD2tbgu+aI/8bwfa8oVJOiTP9FIpt889n4mFU
M5Hr1wnkoTzP4lKTaI1HUdthxCz9iWypx0QpgpmkbhU7aubB7+DANspVn7GDEYa9RmMK5ZNTfrWv
qLQJIZ14GBwuVKVJNgM7c3TEJZ3CLLoqiVZvfkwfidAsxoSM7kCDYHBr+RpWEumbdQe59HhjOVqG
6tcXwWkPsb2Mk7RPc6y4wzdfYY9Nw5tv1gQRAaxPbhrRVKNZtp8k3CHnJ1KFE0gLiW5ydGsXOEfn
qX4HwGX+QmscCMq5t79fcyWB9mNenlo3Vd08XniTcQG/jlL9EabIoW7zoaMZGiTesBlMTbgGgU71
zn2wL9twYB7YS1xDig1v3ma5rqrR3ruPp3riTMaZLwYtYMW/kdCbYZ9jpSSPjZ5lyD1WN7iPRZjQ
xOS8+aegO7zYjIAbyntxpsK0Iw6U9LtYW/so19chl6n2IKfVCL14pxOCQszkOalMOnp9MQJgdTpw
2di3RuyM8X14A5rl1HemqOHZWKFlcHkL8WWDOxtnt91V3T+rrfUAHk6UZWYnjPyZ1q5pPilRxyAs
BhLaxrSacz7klMJf340H9mwJ/4LQURWUdqshOfgm2M3+vbe8SoPv0LwPqFQ/Q7NaM8lnUr2bam70
Yl9poYuMKOKvcbWQuH4wcHBBaSwOBkrlpyQVr3Q3f7scWssbI6rSbthslplbfPScDSWkO5pux1Oi
7675c7Zgw4QMIgQvnlQjlCCqoehOebmEOh6x2Ejk41RS17yYFUkgMGiJzAhqMrq5XWHK/sy3V5qu
/mjX9xOgZxi8e2EMVfhO2q2F0Nn0en7N6muybfyrYdGDhK04/eJ0r0c8DmNoZAFy/FljyrApD3fs
v+42dAlP7Ya1RfDpDTuC//Kx8mpm6eYyIpLYMDQ0l2vleSd6iNouNMCn+l/4zSUnn4+ANuK4p4Ke
Jsd9zWrwa2TMq5pFcPcXEtkO2geKI/yEURDVPGiSqxGlClcUz1cKDink6H5wN4VvMiD34OTLCQES
mjviW90nqkhu10lWlcdeswm1gcpPJmISyimEzagQeJywa4srg1VhN60l3WgzaFTb2QTaf8hp4JUC
bJnt7MlJFGH/JYivG0HCmC3qwpXq9Ho15CgPg1EX/fEWhT9hclirqzC3F1Nc5nDwAZQhV9Uf6O9n
PC/Oh9IXj18NTzWRw4Y9WDhZ/Ntf2tUvucar8c8ZOnUIpLhIDhU1iuE2ijm5AcJ0Xtt1njA+nB+k
tFLYskdeUbbQt4APBrYWWNIkxuCcmfI1cMwoW6gXmgymud+lCQs9OUwkgsAJkcQTHzaZEYmLcLSx
fvarGmUucwmq584IiIQfZg/2d5yYkHqmOTeMPtm1ZAw7uxRbeQuQjkntyKpRxNbjdFkBxRi+iNMP
YmeOXV4jXdY9rgq3jNyj502o2u+9s01LZCKDOZUxcpHy2xUafLgx47yLA752ddCDu88lbshh1U9y
NotIFs43JacLOkSZyqAdT8j382lsCK4pirrEwbNmVW30FB+oYSwi+wlMOPVultglBTm3rcatSSzl
hfRhK2TJXCC14y+gSDhpH3kbGx/aR3B9sGXXJzg2XHL+5mxFN9NNzJMmUQVGPuA5CvKunFWMgN1G
7g+SbVKcjenZ0xhtdWV2D6MypKf58Q0YEdALti5rdOQhlYHfLIKr3PKKF9f7hM5txtezzm8lqLe0
M0hPZqh+sutbnBq/PlK1wEwEataX/xS1htTpIJksTz1Zt4lWchP/pdoRuc/Gzf06YU1DSw5RgNAZ
8m554nuuYSMwH2S7S5292duxQJVg9iuRcufGaZ8SZuRdYU5a8/4I5xt1oUDiUrur1W2h7hCWtn8r
ayY2bjuS8KTgiAN+ZqIRDgLR0UYEpZ62gUysVNeL8OwU3r0oDto+A1bxGPD7+Q2CJpFWh4BFD2vv
jsliv1i1TH/OB8fAEmChX5UxFckeqxgQI1cB5Ohlcl0InyV0A2ii/O0GGIpDYirvpTUpWHH7174T
FVlCmZ1uiPSc2Yj/ExuwoQ2kVFXD1Acu+x8VMCfNey1zkESP04ui+TZ3zlsV96O69s/O/kcyjUvX
It0LbX9xSZqn1ItN/YVt3f5XKd+iXwNX0lHWg1GJDF6MsvZ7DNZtsd6ma22+X219FP/VqXtuwMNF
p+lUG5kAhwUcm8Q+vgMOWfuDCGb0T3Sm1eOD8Twa00YbsfKYpKOc4YNempnUYbRpL9x07e5AhIIw
F0m/T1XPplZzp0bDUeZEIwfIjwYhz5R8rHpbAsOw1EyeJ0aIqNu1MDyP7rpotK1JAyaTa6O2SzxK
ghEnyWas5BCVhDgKROXR+Td1HdfRajGk3+OvEmtZW82G1EgrcOFgSCyzNoTydKC4M//CwnP7ZNZN
h3Xq6qatzwLW+4KzIQ6ziDnvql9Ns/Tj/4lvfR5gN4yibTng/XyfDiV7u/ZEWvWz1kaj0lda1fIf
VogUWIOr+C6qwrE5ErTgYedlt2v0ZqH6CFjfsGWND1gHxEkDCuYpO9qgnnD6hTHeQtz90t9KFCMV
AcAubhR/nZaxOb3r+ikYe0EF6t6AR6y8YyHr8iHiKOTeh0pBi3RqLSb3C14JsRYHCdygXxyERQO2
LZ29Tj79wuMasVN3GPIV0RUMQ3ygyODDvwIbeenGQGpitIyYHukZT8u6NP53+Tl8JYFJ8a4fGaOH
EjHUpt4kpNZjaWFKfoUR0MUsMINW9sQ1AqWYe424py8OQ2fszbr1+/Hsdq82oojbGo0ZAr49+HBo
3zz0FqUHpSKJtHCFphIn0PfojFD/RJVaoqWz0p12AdQ9VD7xoc8YEk0Pnw/i9AqTjJghT4keiaNY
pvkBpaND3qMcmJtIoXkq3/K0hehBW7WGm90nf3vunv103fDrkj9xfW20zxr5c/M66mIcpFZuyYT1
18OiXSF6zsGP0L851cDnCBZIkyFgAKifau+yU2j8vwTd/mkO4jKwLodz/z2lH4cZEHblVBXXVNSY
uBYI4q/UbK5ereaU+bnjymK5LH8kMUV9+Q3B1S+oiKZJ0mleLmKMhcx6dvBEsQc9Yt9R8z6Kr8Ti
I+u2m9J6EBeN82i2fjEXFMfpJTWZQKYpww0OO46+x7lmjz5mgL0q/E84084FmwnH/ODnyz4ev4IJ
zbfeF2sXuJ/zMaA+ibqsqyiaicGJUQpSlTetkNSNijQ1+N9BxcaLQMrlAiUvlRQX3zpAN/5+iUys
bSvc3qQ2Z9deyQwR7WmAg0IpnjPmwXV+4GN4yJNsl9hubiRAmDDlVpxC6n//bqctYPgCEVUrLSnp
yLBFiLq8fFXets5crro70PZ2+ZYPgQSBTpU8ZGc+lfW2DiKdXR9+6k1iAO8+/F7+XOugxhSKBnEG
0Umfb8ZZorML55hTnf3QXdoSEQ4FVN/7v23LC4tWMViId7xFD8wRy6hL3pk/I5dWWU7PcIVz74IE
x5CjJNT+w8xrMrImrH8GvSvjkO0WvHFB5qmb3HFyBwwk8EDYsxJkEKGjjxuHCTux1+rPZMAnNGFL
17oajMYAQoIifhdL+hHRSYSFAQtgBar1oRwNIRDhsOwiD2S/IwY5CbIuKz1AinKVghWhMyFK/YN9
NWYbSzdZ8gdRp8vFNABTEShNT2H331hD1I/eDgF4AxMXewcNe2vb944stT17TgpSH4hL2xTgo4YV
bEIdczktEaIhCdZXNsLsbRQC5GqWancuMAimkB3Pd1l+Np3uygjKlPCPbO+eRuRo9MOZWTUXktgU
hKFXZRUOdVnYzGLS83pnbqYyFvmHFQLHOFoxV9MOWKlsxXiuzD/ajH1mHzvNlUKqGWIP46fccA0R
VTaV8aTzbrR2cPQkUdYasYD1vSq5AEGkdVg8iPZ2sFK423WSvdyyvCnKyGV7UVKdhdV4McYKiE+m
rrm9eS8iOWfnnTBPZLNA7e7oh1iiMvU108zYHFL5x8hnQPV9pBfOgTsietMl/LAdPrue1fw9ZOR8
b/zv2AtCSpH+7pLJZqBkVtyO2A4WbsyrsPnfw6Dy324yEB6vvGJheplVTi7cnvvUkS/vKgERBgTV
nMnQt5DEwMPdI+MF8Wrq5yTsrjPP0vLUsMpgdZo7rfVl4khN0UlaeYH/+L0VuKBNyV3Exhf1gFRJ
Q5fXFM3u0UQJSoHYTNRx4MRW5adifuV1b2IJJ0WjEBN/DZ6m3/tPGl9H6ix7FYOpHK434IauSLci
/DoMmXjwu1x16yE+vUcXlMCyzz3VhwULSwEHVAUIvF+GjZSCccd7/wo2GFShTcXTTf900Hh5PKGU
yl8EjhpWWsAgAMfh50j8kK/9CJr1jo1jaXEvoHqi4ne6mIzumkR0apkBSxhVsA43CLrcoG0xoe31
R+s1tCkt8qX5TKNphWx/IkqqkQDEp2wMxlKdpRilinKaNxpLKHAJeTq8uRyR3mZhJY1YQgpCk2MK
7Zu4/0lKXCo4b9ArjZR0II1EM071X2OZlMPjvGdYRs7riJnDmRfPQPAHGbsxQb6ym6XVUpTWx77e
cIulqNrJh/ZJ1bfYtUBEyf+VQAfuIBznlGlpF42mKEd/Pa9m955n2qdDT9jA+/G9Swrkt7ul1mZ1
Umt00j8CaU9+i5di48P4ZYZ23ipfD5YND0LSlGGvrgPRPx5zpjGSlGf3t8RyZ0XSN4zibaaZTyQx
Uro/r5d7hEWXqp7Mq4HYyVMhtTJj9afnq95Ypz4T3/lauhGAk/refhjYRATUuIflGTO4gYfgotgE
BAVYg4s4gh6CsGPtOYCcxJ99z4RMw7ouk1CsOPciwWhsTaY8fsSM1lWeXZIrtva2c66kteKmzlfA
7jQS3z35bsLd5Tizcygqb8jKhyZnt20HV52PSt5/Hb8XguuZt1FJ20nQI8ETxZsovLkVvDojoIrs
QSZHMdlIQz9tnZpzge0dzvGTbK+3q+yOVKHvXx1qIMOQlfp3f2hG9PbV6Cz0pWLjiNqTxyF+SZh/
vAAcjl8KpqX3yk7n+8+vTL+aN2meJEwjbTT29eu0H+ShMb8JAsZf3o+3YwNxx77KyuhuSejWfuUG
TJcSBYis20xWyrBus+5m98A5DctbUC1XZSlt17p1xN8jV5Iwm6ww3HqteLNMTnPTu9ReFv6kltzA
+W/GFJ2QkUg8EwFu0I90vITDCJ0ESNy129bJ6a4Wztf+CUKyjpKW4fJA4SNz6ODRIZAFlE+0FUoa
Nhirtj8UUDK6JHqo8zNUzpftlXBPWwCtMORaQCIWdQH9y/KU70xtYhxaXoTbjf8uGzXLje3VZHJi
XdHMnTjGXhgKox8ULkjpYMGLbS4QFX5EGmch/qnT8TSK6QPV+vweicKupA5xo0y8y0L/6oELe+E9
v+G6sBQP0WqN6fjGPkj45EE+pzTNy1ywmHd9e5aBA6mh5ZOvoe1uyoDHYDOzRPIFqF0SDHDORw8t
lSHmOph77lwStdDE7PJED+a2MLn1QLnJ8oP/8bcdxJXznsKyBXpeagmT+K4fcB2Mn6WpAQzctfiU
uY288YGNmkbHNvQxOYfuDg1zZXoYL1aSDzjDegh4Y/jQHPLd42TPUOvqo6niYIJUpmWSwcokyTZL
niE0/PvBQ8nIef+Th3RoVYTLu2wdFTmkcBtMcAKPOoK8vXP0aMdYs8/mXgPusfvg7NrvhjyZ/p8P
Kv4Q4+WwtOtRoJGkTqGYI2bx8TDMr3aeNv+DlDoyfoiAnvikfp4IKagO00axo9nRQQTEIjseZo4T
tjy5zRAjjBs6jVusmQu2rnm6QqOHygdYw/OGAeAUZ/O+Sq5CjcbyqQQDkl0Ow99BoybJPqrbOEeO
v2dmlzBPqUxh/JHus12Lg64yq1DMwIrthFDkuVb3ft6lKTyvcDMGVcyJvWwhPuWFKQid0kKqcVAp
vVDqHTibiRqwDcn5Q7xZAQ2IGvBvDi3M3qRrpPSIniqmzie1D/JZZyHo/NnkRSUYpku+b92M+pRh
eggrs2ydjqVuDapNyp9OH2iHhRFbro0bz6aUsfuVxrQ2dNasrJzzJCcO1vwhPuwLkYeDjH0E2Eo5
hMVeoPpTeWUqiX2W2EryXBOM20F5LAcuzNx1LAQI9iBkdIZRKZctf46Jfw7HT/UrWeVD7k/s3ZP0
VY/mlH+TzJAae9viqJUjnrBQlCPqE4DsNvUsgomI+F/XrI9rTaQEexoWeIgFnWxsysnf6/A9GcvF
QX4TovL0lWApRxog0hsN2tK+WMFSkWpiFgfddIC9pEeBwMT8unOMaxEKDhd1LjdOhDBQSLACQ9Rm
Cgs6BI2iKgCMZI5dOskUXVjDwOXJi+7ESkjfYh8lP194evwlHkbdOjUULb3HuOaRLUSn467A7GsZ
WRnvxJ+KoUHFVva1UVkf9UU1xFdHt6emgOCKJBGOopSTq18oWw6Z+jl6O0uqtQReLVc2C6FlEECv
2Ixvg/EVri02fn/6NRWtxHCdY1xs1cC1tdrVO2ABStJlR1BZcjJ3yHFVlpOz2Nmm0jkBZHfR33WY
VI357r14ubvcMvuTCY1Vq91AlvgEhd/97/qKNhwDg1hliGNYap9Gv1oebEtmZztbmZ2m+B9eN9jA
s8X03AFdY+Fg4NYbKPXQRH4KIXTd1GfPK8q1HmtAfwIsazIlPfelv+aGqNWeZXJoj1DhZKKODPAr
dKpW0I7TjG6c4HtgSt9+VNhuJbueoFKVAmicJw+utDA7WDd6Fy1N046q88uAVO1u7nerFEgB7wuO
qflSpJtLPfncKCa5Azpy7VBVJBh0lsA96KnMgrXFw/I7poJKf5t4EDzqOUSbzbgIaatE++id0UcD
IDFxBIriozBTTonXL8SPnwx/EqmPegNcbB3s8u1nUCPRsiaxXFR3OzBIHNEVf5yQm0nLFGtE0CLB
PUfbB3eAlckQtqoWCQgD5Q83fZATMFAGNtc6JHHD/ysTolOD9neb4WNpLzRsMKazMIlK5HcwT/n2
Gc+jQ+j8UGpQ8ctZFkMlj64nKvpY0j488uEz//X+Xv/jxHR0AV1sCvtDicV0ImUcgYLRZk7JmTrE
o3sqbXs9YqbwRlCuHrOD6w2PbW/S8gLdDFGe1vIZUyPD46OEsgvTr3LwR6wXxL6M/uXkOMdW9hHZ
BrVZjIvRT6QFVSsj3nwjlS1sb8NNQSn4S/LvphpXHF0wreH0fWdiheXOQ6LCe/8tNhpLQO7HqsGd
zkBmInAVmxlHdCkMU4U6xrYCnnWf1y0GYIQVlWXIEvU3x4JjmbY+VW3ShkkOR58dVr95vhR88VTI
2xB2S230altgSzbsMX0j2H6HeTQi3a3Rt3d9IF9Tnlwhi4Xp23kde8Um/tFjO57hSUTDf5jHLTue
NdPZk/rWbKsiR2ovfHgptO1z0BgyPfjsqK7rkeBtAuwqVrXbK2WfgEUA1hVR/cEc5SehknfaXZop
9C4Qr3LMeEHdXBeTYdNjveiWPBmZwiDITJUT0dPgOWGJeC4vg0dyv++gv5ZX6Ea/m0x4sMU7y/tf
MJUXy7xtMzOFXcVHwQBNoQ6t+68QQ8ZiLWRTJoxgY1b7gnvnvCmQXuU14xZaZl5RgHcx//IHZg++
qGCbA3PbSHOhp2VOAYorIIvsScg9qlWt3Ru5vA8eJT2g6poBzfpp5DD3q55ZkdDU/O26/uhvEpAe
4HWyB3IGfUJKcZWjrQevgj31bGNjxqzmNB9go4306hGnwhC3Ef9jMkkWD362QIHCV9Ga6vqvJwKY
U1QkhtqJ2qdH5OHJHlCIYBcPCSRFb21chAPg/0RIGPkfWH588dh4IjzqC/ot++HVhy5e/sTd2aHo
M3y3ZaAnGwyYWFFZ+E3YCxDWiezknU0secug5ZUNHQFlh4Gb77uo41spnCPhVTyUfNkQVA1TOKMU
3xX/TobLD1g8aIIucEOp3xlLE6jnA9O+U74NXs8HSkw5iyCXqReucMWcM5VkTLvAvplLukOdGs4X
5jS404ScslmfY1i7idpJ663rYx2aaN9fLun48Ia3LtH4am2aGH7xpsu4QvHX2L9gnZ4wVes=
`protect end_protected

