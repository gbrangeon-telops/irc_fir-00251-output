

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
p7Rd+JJS6BPhm3C8uEMSjtB2IOpOZImN8ABL10O7dB2/wknTrPPVnggIUugEe0Un6rsHScVa0yw8
WbsjeU4skQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
bancDuzOXzE/C1Vj5QpW3wyih2C6ymZ1vv70urQ985WeT2kXc7KQyN00fbod+1ycgrcEzdZs+OxF
/cQLUqqV1PAWyHyEqXlxABFUHjs/nxBl/f/B9V0jlBhAzKCCHBVtW+DFv8KpHE75Z2lg+r4JTjg7
zQiXYHxUisemJqUJdhA=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
rZMEEzwWFXOuo5snJgtfZx9Urf7eZRBCxLhuSc3DgaT16zNB/FC6Qo2PLk9pQbhTwkt+6VFrAqaq
rIuJ+6NqrQaj6tzRnuILLQxRIcZaZnlaNGPM0QELT1/pgSpbDRVs/w+jfcFf6hDgLWdb7+lF2lZt
EzdkUS2z3RzGxMw0dEl0kPzX4BrObwXWpUb1u4DD6JMZb6O50zBS5jLIs04xzSPqxA3PuLRWpuc8
zAMmWK1PCPqsF6JmUA+ToDlUTA4DP+Qb/r/OItKXADHbpGUiJXq85NgUc8TOMYazRmcSDk09joNa
rvnt13K7ONnKnXu7DU1cLEZpB6zC/Q33/JmxrA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
fSUvPGwGSOzh5U1OjbBgxWaXchd+ErSm3+d+gvsNPzEzvrhBDlsbz7cjXesFumQgP32hemPRlsUr
lFspe8TkimNAMoMtRIt9Rpr9MJxdvSAJ2AckK92TaQKYGICYWnAAwRZdM4hFhKQynq8onwVPOItS
8G6qhIBnq17qx8rO48o=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
MVMseSXR8Gidb6hUpBeQo+a3Ho0qfbo2cQ4XmaaPwOf5p+bpngyRNVgFStTGlS9V1Gq9sxZR8m59
KVYbqvyTG1F7VywlVWjcCzm53JiHqc7770pyh1TFlHFmlBkxaKOZI17/BbAJVPtrgC1AFUgqJIKl
KWFzGNfBnaqYhwSBpkZVKTp2N/RCKh6/dORV7jPLmH1kXSt5iI647oKA/xzmV2IPvCjRau9wfIMP
3BcMw9SliL4YOeA2gPuyEVJdJ+sinBGqyYpGCshGE4syCgACrJDHcCC8bST8+Ee2RwROkSw85PvD
RmNqdRJR8yBkuN8MggDeHwsPe2oFAGN33DaQEA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 56304)
`protect data_block
C8ENXIVzBgfZ2FUj+Svuw2jG3g/WFFmP3es5fOGiSjydw0n5fNQh9gPpxIQiweSnBKISAD3K0kzW
kxSrk4h3asghFIJvc9lb1VOqG+lzHmeqGnamyOqBS5re3Y/ImEEgJYkhot7/l41U+aEhvLbNFIm+
/fa8d2xKFxCwQI8ONPqWHdBt1x3nvbbLIThigUawY4A90QS5MhJDTE7tXV8bnO45L0bRGLuo/6dv
TN1V6hakD6wqMzjeCrCRpfbmtlcEMRn7U8KqpUzBATBM3pQmKWER7Cb7yeWuBvclt84GlMG/V+eE
FzEPoOORzAAMkLUOanX/tEJk948oE0ENuZlMlKg4DQ8EM6v5eAuuBgxzZ0xyScu6baml8NhE46ve
N9lsvVDm5SL75sjc4THmysZDVuZDUFDApVIJ/wZbVz0CnusWSBCrohLiwhshGKO4ai7HIWNpPNqT
FgNrn2IrEmKO+5DDX+E+8HQBIbMCglrg6wNVi5o0qlUviPy3Dw+swQY6buB/559hNTUSICoN9Pva
I+gzVeJZxGYajOpkUESj8gOrXO5L5rrtPCv10Y5hK7i0dPKWyl2Nn+zMNgcenr9CJQMgQkjzcmfq
jJX6vYr0VvuLUCMlpIZMUUb3PIz0TxnbpSrkcPemmqXEexf31lsMm8QdfBAd4DYg0lPLQ6kCJ9UH
RfEwZQIvOLtcR/Qgs8CfvjUDg0zfx03x3L0xv++Ds7v/cJrIAm0F2jN0Lj6PWDPu2iZ7+t2I50xI
vxlrtWbsx5C7QE0WjUxDLsccX0JHcGFpd3Z8LHkgUO/WEetWZJmDf/tLmqWucHi+5D/kr3UiiUvN
FHfhHV95H5UVlW9sCdlFh5Vr2AXLtbqWxG5CqUYmBAZr187ioDMZWGsnHHZ9D/jOR5I8Doxr6mCi
oh7UcTMXd6QM6W1TWAI8USC4tFKkFthrITLnXPmeay6biJWjILC4eiU0U7h0/HKtplTZEFTXtCTW
ipbXedP7XhedH9i5BWXcLTvbl4V04s4/MCilr7M+GwMF+K0I2b4KVUzmjL0IxaAvOXNxwitBfnUh
+2ovhIZHj+vxMN8Ik9+Y9dfOV7yR+PcRmVWm7JU1oRxzAkQAjq/1f0BqKbwYc+5jUMtM2a/5louD
AZY0dho4eE44KbYehwHNCv1lGCiii4Ut/7yWKNLlAKRiPz0/c+BI5r4niyDoN5oQGkBQvZv68AvO
adauLn9hGdhdlKPCEWImQBQd4n+oXS1Y6Etiq55YT8AwMqUb2ZgORwLcgPzLB1jPYANj6WMg0ICd
lpyQ4Db32H0U7zaKzioA6ugNSsFdmzKZMc3KZZjBHBW5/It206uNbRPtZy1zgpP+wJkQd339dTR7
u6gQelhSrsEeYkn14rkcqTX34r+e6dCIr/EACHkyceteHCLrPVDtCwLrsm7jOCrLpSktjFsTD4h7
OyieM95HWERXztFQla3AewJJjYHoEy11SSwv8CDuJve6khDMxBlAmLWLNH+f41YhBIcQHATn1ufH
oIC587wVxPCF/iE1x1uyAZ9ZFDH+nVZjw/Xg5H45wb/19vGB6OviUNV4YPjUC8R8qeH8ajygDltp
gQO2hw9GXauGjLr/2dTlPk0nh+TrH0DFzrtb13N2TBRAPYAvecxnTTnrPLyaK6Cfb9ghyDooSjGS
K1pXfHCaUY3AKh69jxx563VjyewpxtOkeKQGbCi+/sBoLpVfLDMFRdkoPlgCi8b60no7RTccO2QR
qMrSGWyIpEJ2Z/L8LkYbuBvv38XzrevTbYpBiKVGUD8ihgfrHte0gZxvHVnqZbNkQ2lH+oLvl4RA
jBrXkMDIuh0a/ljP/hUiuaN9w0lSTd4plapm0DTzBOZ8BZ4twGyVmT/DUYUW0NrhygRUps9zLZ1n
A2Tx73ycn1hr/7+MGcV4A7bMEEfe5phVxIuSwhvx4gSMLio+TMfhOC/5uUkO3Iiq5c7Np2pdl4Al
Ium1s8s0EF44Ah4ogIalsSxShB7EFEtq0RHlkCKX9/Toc8HfdWWyFBTuLkLQPThPVIplh7c2RehT
lbm//Oeb533SiLZ3uIYYmhkCGIDPxsoO5vFzyS1vjLloGFbzXGKkffydmvXNM3w034sk0/mIZjT5
vQ8+eQgfKcX9U9KAFIiimA7iNRALhRIrSu2cP1+Q+8UymajaLMWfSKMwaMrb4jVyPuCQX1PYB7ZO
RzdmNasdRR21BoBbTSdpecaLfmdBiqUqnz6KVa7wNo6ScVnImrmRwcIXqKLQRTpxXbqbfTCu1eum
XMlsQwkVgzzO9juzETsvWgqsatM/qxIealk4OqzpRW75L96CNH+SoSQy00DPVbJJaemafC39Ba/g
+E1slUQPrBzNm6dsQYxvRRZNfUN3GGrwLx4BBdXTqdYVdFvdvbAUW1lPHIz6z3fQkhOzDthYGTC3
SMccf7Gh+xhGVWPhb9jyTm7lgwfKurDzejksoviHDyPP/3ZVu+xgHCNoukHhVgCVlCauhMAMxHH4
8UiOteCXd3SNiuvfRfxGhkWbbcrTp5jhe9HvkgX5hnHYcYJyOmWTnk328Th8BcSEjx/gya4MFpih
86JRov2SxzkDEalQcWfZpsOBKs+QjLiQ0RvJKmx/oIqrcbMGDbQw28S/hwrfDwDh4+t7erh94k5d
RHupLvgkYOVImrbS0Hr3zzrlc4EPZfxT/ZLRvwJJ2bPeADqV70Q3ALEha69q1WrrADyiFFbVqBQv
ZadRA8GN9t6sEJj/KRzeK8xbwpxvjEXjeeyVffQDqOpS+dEqpo26o7DZID1fH6ciWbx1gXi/mDCo
Y90L8GKp1mbl4PGJY5t16TGfe15Uff71Yils+zmvPkkYEzuwc5BPLg5oYLXjYFyv6VIezNKKqyht
9ACGka3r//cR46t788H2PDz8SKaRBW5MfOMYjobtExcjyMWJ9NwSl2l4h2ygyv30SoLJAcbqGnuB
w6sBZ05uz9mMDkbFH/tsstmEhl4gmqiPOLJxk2DlIFPODs37BMmKnlY78tXamVSlRugrXQIeYXjt
jeoQNxBHWbSYjy5MsyyjCsROo2WoWKhlYVft1MBBHfhhTGJFyyyAk6jtTsA9zSo8ozGWAqF2TQOb
C7mu8V3d6HUuvqjsQ9FFU89UkRW4kIDMfXxrV95Jo/v7xSfRc5OTA927Jjo3ZSNPCFJ1sI6w2uRd
o51gjMhg/oKNSYoq6vgbnEnLqE+Zo3Gks5ZwW4NZOJ8owJzQ5Q6jjzZ4wj136yxNzUG0f25plD25
yz0neVQYR+Kk9Yk0Z9/rqm3KtKzwERHv09aTlTKGvqpiCWn8QhnVXGMei9iXBCyAO4fpgiaGMK4T
Ph7azNnG0EeRn3TYw470BUZCPKcEvKXgbL6NrOTLT9ik9LIVw4Z4ZWUoDAHksj2JX3fwtlcYgcgT
aJhvyBGXgRSXlpou18YZI+JXZJybRGU3GBapwRirRAaZezKmLNFn8PjphqKxiOUvqz2jmaE/HSGg
AoiwB9+nbASoRjCsh7F3RhBdhwAmH7Pnaym10VATgIXJbpQxHIK/HjKb5jxHj827qZPd8eeVRO/n
1cQjvzTYiemDCQ1odj40GqEQqJ/j1EG9sLycMQ/7PL6BCSROpxeArjFRyvA3X4/ZPAR/TcNCg0Q1
uWX9dFQm5ffKgAdyKNNR87+BGbg1v57XhU7Y5MKKA3cXBvEZL63AUVmHJLr026KSVHhC+qNNK4+Y
uCEWTqFE5fxvbhewqcZf6CQZDXbsnJIj2Xcfgy8badBAlt8sPCpBtS9C2+zyfbayf9jZaRcja+MM
XwzdMQpQOqEmw5/Y7XKYG1fLzksQzs7tbYpx6kX26tyydwvWwgz4kVN/17yYeV2VRGhUGmpMaW3s
i9TYGfyHPUuS77RjfJ7SvSJWhqntO9DMp0ugpklD/QE0GVkkyh0Mcm7ikcjRweT/iUZTeV3yNdDq
o26XIsIdg9/Aep8xaeDC+s/eAvFV2E7bH/t0jGYs64y47tN6w4iU3A/NAItXe1BvJ/xVZaWd10q7
BBtlL+RcPWE7U9Y1Bbw86Lc+YBwCEGTMKLYEIrdPrV3ZPqWru0q5B3NGs4m/Ae0BTsl3RTvlnwUE
Zjktggq5se9xRZ01jg0pwBonLxVyaY17k3vwRvj2TLDAO5YW9wD1sXAGZUy/UE731LQQAoS5hat6
pFXrfzxaFIc3HuwB1V4Peps6vvRpTBGO/NtBu6TXLRNNjSURaEvustrn6ZoOFwUb4nRMlDMpU4UQ
fb7YXbJlx6Mm70hGt6gwkeTBLoBjsYBJur5H+G8WZMU2+rgbHtfVnY0/vZmPK2cp6IRyhHXz2atZ
o4OW2wg8pZulkNQMb8x6OtJl1HifhfvGpSpl5z3HZmV55HvXQGUnEZ9ojjWTrx+wblob06srB6Wc
mCNN2AcTSoA7lk8k95oQJhWmvjRVkA4YFLyAB9rWxvy9H9OF5B2MocHUn7Zv+8wXFxqzDK40O1Vt
eeVACnw97uJ1IIMu/YY/vOzX8BScveNMNJ53Co0oVLDBWS3iKZjcuKsX/kRQxDgaMrnsopvYkXUb
FF8oj+rJLttu8+9DNhhVhis8n7m6eBtfhbgBZIFTl9sO4KtCaFJEczZFLfVgpYK8qvmghPOmeoA4
mWTu/StjXwkUcveMvDSpqATbKWLndDziButb8HrblNeIaXwNWHsN/VBdaHHIL9hx0Nzoft9l36a5
tElQYoEyd03+PCwRoKF8WZ8tZmRxTKb3/5YcCgEqpTYGwFS0qplCZMwDVqxfAF+AbtbJOtIg6/5H
FZce/nk1NC/Xn0teXx4PKnB2mCudZ5j2A1L1e02lhZfY3ZcEZTxENaAxrK/dbbYDTcGCydjudbGQ
H3MJAUuxSkjjdMDUDDN5eRi26NAkQCYm1YxTc6Be0ST0IsLTuGp4opdaxpmRqIP5a1L1/JmSbVQt
cJG4MnofVQAPTmjPPtz8HFibxDFO6gwKt3p39nXmao98dPUyCAopahQtNjQqvpTTGGQOTv90e5Ha
KLzizABrYzZGHlKnxXyGixwbm3twp+TauRbu9USLERv95mFid5hjMtL4bjxYJTKX7sbeFLZO5L/r
pRXvzCAdLXp2IvzEXL2Ju/OQFFkWl5Ax6jA4CZdflwHUkg8IABKWNVGHBpG/g9sMyJPj7nz4UOYm
4ODAL1hbdwUVJnCd/6FStA5iiRYyx4ufx7ZVzjTEx92Idy5UA7WnlC4cGwFF5hYDPjtjmfDnIwdW
oW83Z0ovYtsdem2jeG4YuZ/FuSFJtNpQvDUv98Lex8r0AGAI4pqYPCDzHFZconcY3QC7dSebd9lj
ge+BNo/E0PzvL8rkyElCuBiorKcBr3SFnW6C+wXDVspxcm/kTyYkwUzwW4Qq+3GTZmlSsxJ7yEid
PbVJxS18ZSPf+oIThVbqYXNAdIA15qglWiIAYV+/BOYjoAe198zfzzSI+jHhTVcrOmf4+Hb4YWOE
tXY7cbytzzbIa8XxhWT20Ycq5N9AUAj0INfgDekbV5F5UusIi7N8zicx8lTKw5rGJ5jrag5afXCk
Bt2oKRVFlrAbp9RzgPVHZkXwagKFETz1ONpRGrcgivxIPdje3jtI7MLI/s6q4wZYk6akc1KzN/P/
Q0/kNjnrSjqWMbadtqX9s1XSCQuIwUkTo88g2fvLqqpzU8D2peQMMwveMK1lFnXnJxz2m+M45VtW
EN0bFW1DohvHS1ypfupTrKsi/NLxdQMHe+7dL7OcpPv8tCtqF6abY3/j7Ww7XjUGgj6gi0OY+Gvh
LtkZMM6KsH4AxeskEYR7RyeiilomYYBtkyvDtHUMzfyjBrDdxB+WvIf2YrwfVxUx9wkEk7g/7PCG
ciX7LKWrUcsasP+v7wW/g8L+l0onOvMf387XTD2PeqLdmS1LuufTMS3RUtc6R6sAQ7ZdJTX7JrNx
TsddSb9V1nWmritu4+ukDCSi7hNqNJA6Vc5osKv/LGEI2fGaxyTfg7yzzXpH9UiwlMjzSBUcNrcW
wcmEaWCNM4vrmlPDm6bc698cl7D8Ih5hElFKLQFUFtsgW0vNY5TuODSHGG1Xvc6sei/2ouRUkZN4
GrWPPovgW4IIHUzk3qIvHD/eSAKsQWxHS7FcYOZBvdDrbENkXO7+WTYlOfTyuuprZw57U+9i/eXc
MCm+XrXzM1MILb3TAHY+AK4JM5U1kCScv5tRaqNf+f4KQK/qBi3D9PK4PJasY1VdG7hp5syneBno
LgwawV+s/OB5B6MwxE0dtbYpjron1CpkA6PrlJWdFe0dhjYXrKbdqF6NAgA39+VzWf7vdUV2555w
YSMBwpLo+W926UJ3uTYS/aaZ/r8YymYvbqCABy/2ecvoj3O4xHcyAZqeKIgVOWRWlFP8hb7M/1EL
cxsbtegBlPyKQCM2TZLPN+NTElVxDR3hTF7+FJ7IdpAPCRw/+37MLV/VkbDNu+G74U1yJ0jSkO9l
ER0Fpyz0wok58udFQps37HzqXXA06UEUM7ufHZuVBSt43PLyigLvryU/+7VPn/pQu3xQ7o35unCj
W3P6+6W6Jf2uRiDjfLleB3cu10yrZPmrirN/a3m4PGFKYklitP6tZaOZCMKdx0Inqhygx32PduRk
OER2Wd2c3NWDuef9E//6QkgwhoBUGSDCITMeMGGIfN4ZZryVV0mUEoTMx7kc4AT8lDn8UtkPBOOo
jRZnqf8IyrEXvs+ooOk5FgAoBCEYzrUu+14IGYYgcAgeTGdqZUhQW2Ch30R7NcaywLbgm1o2YMys
aRWZnfrGKC5htpRhGI8Ps6erli9YyjZmmYzexki0TSxAqy3adoEWHYlugpM2Zlnwr2wfz0rRphOF
+tbHpC+lP+RQoElUNrRsOnSr92+YGdBD4vU0VWbP3ljp+/nVXFcTqpBL4bQyMK0IUfoMrgNVF8RP
wTIb0VqVgvB+smn1q3ES7TlZLZeRI9X//BOW3YR1DP2rXC3zGAVjXDhI0E4vm6M5sbrksAWDtX3C
6FLBpK6rO3xQNN4b9W+LcyBY+lC4nrbmZDYaZQxAq05nHC8eSuI16ynp68Ff/O8ZPTC3r+RErRqq
utP/+jWecjwv5Tuuw/ediGWH+oA3FEhKZHrvOah2OeKC1dronAREnasakQfuE6AtQEYqXvnI7H/K
PHAPNAYronafm88AFadTl52kKe3n+n/qJ+aobb1MmTzpC819ZvkWYQ3Yow05HPGfCVWHpd/cTa4G
cxSp8GRWm6klmJeJrn8f8F1YacXT6tPsTXKZ9pNKjSwv1OsaJIZ368aJQ/+/ITFGNXShhfc+9D8a
mjsLge8dCnafekkKLj67EqCULC9xFZ5S4TczJRfzCxyttFty6UZHPcpDNV6hGC9MlgaGLmjGAaZl
y9MTrYijGpZkMF3IpLfaURjzh3P8qy5khwXy1Qt3/gsYgM/SU9mT6wyGSDtF23q2By8ChRlRYSs8
dTyUnWurNY9aoQHRiVeecHNYK/Ivm0FaGkGWOmB7kq7rbklNocDmff3+auSI9Xk+Z+keGq8oCpZw
PlYWNINXRmo4dr7juz/USAdzOXlbGKk2tbW9Wa2+HC/Oz5zOOZYjjTU9ZdS/Cka8IMrBVq1i8XkZ
icMrVG6rbpDNsrJaqdhs3PA2K3wf7rcb2mw0jg4XtttHF8oRzzj9JvscNmE00m71RcBo/F7fZejK
8+Ck+2ITJk+OZ2uJH2DuHAIfTtdCISjPH7yLuXpIzbBodZcpG49O4TcpYAh075qjtfSDq16LV/UL
Prdw5Xzc3bgS08gDeqCELyyeXCSWawGA5L32aBZdv8H78za+9r4rzEzNaHBcWOtNjR8XBKWjvhap
xx//XOIb4nbjqx3hnvTkoVFcm9ZyRU/Joofi41urA1YKSS+AaIpkZcG2JE9ymqsIVHKOAQDTp+su
Y4SyxOPBJNjNztVSF6WH75i0nccph7j+vy26KeMOypakPfduycB6nkBFLN8O07tvrvsm78qSBuQ4
ENf5d3rYK12iEKL7WF+lKaxFxVyBaPQwjNCkuHSWZ3WPNQVZItKnsV8Vs4cUdvXu6+QphAKIDsdI
7RhUHgw7NkgMZJGc2MQBCRO8d4tBaUmDUM3iIYV169iLy6Hiy1I3CxxPfPPiuVuaN7XHybU3loWS
doE/Hq43Kn6DCDNjA50++Jp3peRKOVH2QkkQwXzHIR5rteQtJerueavoXtn1f6mK54DGhuXMyUhZ
T4sxa/7jDuXZNoP/ufGK1d/3Y9f2TEX8VjB/5VgLrf875JneByHpTCW/5dTh0YI5anfub67J0Yuu
k3pFNPMW/yKdEEee0TsCS+/mNf/2Hxsh9jlXQLYr1dyVeV9pTK6Hygm0gMi/alEgwMb7Ien2GQe7
0516rcEiunlTHDY4Ei9KzuUrO+LL8PzYEDdmxbwiH19hNMsPeDxfdwYDEKdRug4vE0QQzT7WFlCy
6gi/yccYuylYaYR+r48VpzLvzrMdjIzAervBSNiuHiKbkxHhq1LqW0c6cbNYMOxGohrH1uKURcJr
GkTa9hp9VoZY3YmJ5nCdoLJaMHtek5MmKcXAcrjeelQ0+ZtHskwC+bCjNb7A370YUiFvQ4eZcXnk
sMPlIPjZ5Mr3hfFFCA3yBQMZuM3Kc9z1DVuqQDzk+gT1beeGcymVWhwbesUD08L4vmi0zKrenPAt
/bKkD5oAoZuczFiTdSsN+I3LzWGd1MzZZ/k5VnbwYWlG7Uxifa/GMisbMLV2Zn7sZ5JW8f1cjepZ
t7eBDQ8RISn8Ksvxh56pYivkNTh18IdmiNgJHv0xhYkMA/mSi+AjtTp28DlvL0i00ZrIR467sANo
7oU3ONtXRr4lIfqFtfID8I7cEaY3PZJwTanyFiI5KV9c8GsZnVQomtAeRXGCsSURo/JR3vIMHqRt
PWbkW1Hok28rF6PWFbOGd36nVitF9GZwmsPBsdXUwSV0wl2W8hQpFWQP4Q6VAton+tPHMLy5KEkS
LTUK9zskF/fp8WH0Lh6f5GiHTaEsZ+XkHDSta2xZCirC/HObqJV5vDIGDUR1BSWzAbEw0XpLjIkI
y5pzNKIjySLX7NYbyJVri64DTgUKOiQMHaH1Wj7VKbBrFydJS9IfVR3qssueDcYK7yaTP4ZZKphw
Fb1z0tj89Pe9BUVVlBmyQhyjKTVvFh3owp5/VWMR79MP6utClGI3M0y8uRkpgaGSG8//Rc2m01up
GJLv057D3VljJDMwufLn7yH6Peg9wr3qSKyfiGnFI9KKTBrkF3W+5CFZzUzW+D7uoPTeKGDZd6Fj
P+qHobIMjraTqSOqYZIGIqnRFM8DxM9kBZ0BqIpGXG1ZMYjcQuM31TO/0PgLkvYQhlMzIBWMmvuP
fQz3OxgZ/OwIbMuwZlfHid91XMVDZ6uW9+eZSde4zQ5OJhiE3YZOzGcrbVb87QSCAZozuz3r364p
i+SxlmfuhQF9AfzCJQWjPVxMwvDIrieG/x09EfsfZ3q5RCO/PtKUY0itTRCoA5Mo7b1SIqnKUfOc
KjO9z5iZ2+zvuI9xFGJ4RrISYwx0Topuo6Qq9EnOyeD/izQuhKJf+JlGXwatwDZBSEFBDFJnxepj
49Z9JyJ41CGl1QP1bSFmScAXJJ/XRZXA08sEiiXvWq8YF+BLkLvJlRekLq3ss7X+Bj9ziR/9MXWX
VU+BxX226QnyOmblIMDtyHR5OL+cnzK4YED4w/XKSdd8IVqUHvCCG3djdoYSaxhlTKIwdm1GK5jG
ofoGnUWKdu2aMgD73HApsDgQC6G+TIUdsV+FPCLzf2YsZQWEY07Tb+aAn/lvjQUB0hk298wrT2jY
Pbc2BkYwRfFlSesGcv7cbWJzuFpDu4T3MekhAmjdgWnW2PNFkHtxO0YbTDZCRuglDhUs0zq3Bdme
Us4em2UrwaaKccI/OyVdQ34Hq0eJWFyI/3MeOEC7pNPY3496wZ9D9B0Jj2/3VGKsV1uxCq86KtGl
p/zVaMrAU/vqzLGkWiGCSWjZLw32Sdj28aumGZQpeoVGz92DVhpVhOKZK4fmmImgnwMZ4gXoY/0o
yyhvEGkEqfM+KII4zKBMIiinfZJ23zZHLOEgkbA3oZTxELX3IDM2SMne9yRJYW6Qf9xpBXsD2fF2
xzT1vK7fDCnr5XjnwdviMjhsqYP/8i3OHYKctFH8A0auCGyLSqFgvpt94lmzwXfAQHqBUKESIwNf
O2z5pRJf3oBoxE/h3KgBCx2kfk4JbEG4Rxv4qznyukDMRv98Nl5Ru3rL7TGRzrViT24kC5wL/nBQ
CGSDD/Klea1PQw3ScjD33CWEHbY6Ph+v4XQynV+IWxLmbDZpdhhfdCdaSrsiiG2Q6leSO/8t+7SN
mBAC8ZYtM+2Fgge+4eZhHAH+qpr7+y0L7aACX+68mYmQyWx0+dFUa3A1SZ6Lm23K+NZptBcu55rK
pZeLd2HeNfYuTEchIt8yfcdin5mon5TC92gY0XrmAEzLvG775ztH2raAQxxpcKT+B3ZKEUfa00YG
zyeM8umK0OOoXDqzPV7tLgpSODVQWTzM2N40RdEo6eArVP5YoH0TXRMdpfcnQuK+UqsPxkn6jHwr
HEm+1Gcd1aqEN12kNGzG2d2HwtC6NvXZfq9FkFjao16zWstOTLoyoz9wkoG3KeV6yKbiq01qliuo
B9/dbuRMvm3iSF208r0120x/fwoEEb2g365eagCnkhuCxvjbjPP9Wn4s8cvmA67KGCgWFaEKKvz9
rkTHHiyH7kwW1tbZrYhX1MYdUV38BUWaHMy1STW0h0bIQm3+kp+VTQ4PO/Vzg/gOQov97iBjumQT
sfl/etfIw8P8YUrTlIUCRfrGbhekE8zCPn/KFhAyZV+isT02ZMyVnNUSx+5JMS2Ogct+FldcFkRP
CU4WGcpViEj+et/AQ+kUKhwMjRo0HImopjHnT0TWpT4CK6QLu6tOf4gHmyNcsVUZ8gfN+s+Xfm+d
Q634FZRvcCa8NchzKHRdEi4arSXBgjUEv7ShqW/lBUW5/q/2xBBHVmAYFiqptwHEyoRb+ZuRjnuF
8dZJJZxD4RoPsJD/zohH6pMIJ+yMhBa8R3Y/vZsM6qUpKwC1dPVVqlZmPaIXlvg0oMoKdJVmS9AS
B6MjCun7ISmomT3u0M+chCi7nwNHkiTkJ/ysoYDycmIOPTVzt10j8hepgnlRVhyBVbBWCsvfxtvU
dU6d/KvF3/EZJ8FOuYvQcKRWDuX0amPSUOymNx17DKW/6FIc430Zvh8KiHIZ7wC5N3cr/U8MAlPr
AkjerL0bfM2ii61ovCc2kgMcLW2uZRow117cnIB77wm/SWHSiRznLiNsGgC+shzy9eNNHeV0t77G
F4sZtuJT5swUSUIJeuZJUhtPBnRZ3Mwfl4hQ/SAzOapUtB7H817KmUJ5rtE3e6Lz/aiHrMRWEsZT
2hrNIHVgrMeTNPuxyCXQDIwifT0QwDRzbGonKJPWinxUBim7PVqaQYO/KsBABYRKGm3g61osH/aj
gKHVcGsGw3HQhYEP2LbbjLJWi0BD0vWV/gC4jtScnev/MTB7dwkvp1Jmrnwi8zyEA162vUlByIry
mC4xWeYqVb+//pXzKz/cePHtongkhWO87duhBeh/0SGM8GRoeI/CjDI4qN6BRh1cOh+DcXQn2khE
2DbxGaZkPgkxO0AbAuAC71Zx0slAyKaZQaulJ352QtGNYcCI6Zv2zcmxvRud7NxJCycn+FJlBy11
zz4o1oa6bgT3cWiRbBErMjlx2njPMLum9NNh/ZeRmXg1MhF/sWFV57KdCbbJjNwpuzw3HMaujYzT
Lrz78dZ74OUFXwgaDd6nwz6WUIbOy2GEz3OOqYnKOTG+Rxz28WsLsypxjfN7A4mvXhCw0JaD+UcA
UJ8vKvQq7BG6PKOR+InQ1ESHXjq3oEGk+cD/CccP+Zdz5mdo2YXTvBaGMQTsg/AC++gRXIwjIrAw
NugocAva6tCpTTryieDCAOX3s80r3zscxeoiZ/fXLJzwhJnDpTSi76MKtfMED003AxDXI0o/1LOD
uuP4zA1hbLydmHt5sEHE+ljd6/spO5HKZQzjnzkdO5uVAW7h8kpvhhd/p1NZHRDm187f0miMpPad
/J7rvCjWJvqWRj1fw9BxMhgEnafvqdsdY2nM7LKrkcHLRjCLgkWW0Z7OM9RYO6CBvPTekcO3sHM1
g2uiC3ZRQgBAfYYlyjxxEdivpsDzxJilYDdHCZCVVQdZ+yJxbfGLDExsnv2yl0EpRw+7yBKeXBpO
hKQsTOeNmh/PJEMXrdVBxpbTdxwJN+5chDtoCcZCle6pOKLi3xcfdEOoqeC0OYIL7MU7LR7fkXXL
txmKWY2ZH8Tr0aYweqsfIF4myajpKG0z21e+WGKqF6ER+jcFCYNUiuyfEz+jqlStN7Ra4xjT03Nu
OxFwKcmcQXa18EpSngw5mC4mYxdGspkOAAYxjJRlF/JfcBfaPA9bMWWWY0D3iX/R0IYNKeP3hfxs
iGshma/boJY58E7yG9/+md+1CKxJCWAyb4pogndBizuoUnb2zhhasSqLWM8vOXjTJgBo2zjPm0fh
LBIZRUCa2bafMaKpZ8CHsQG2UneAxCXsmvDyTlgBz6198Zy8KqTgLjp/RbaBer625UJ2qmoAhY6V
lINwofyjrn/h7tHmWi0Xez6wkRaXV2LIUiUsp3k3oy+ElhDKOVS7F+ZWo66eo4xaBiyOGyRxrZu/
1GV4ynDR3BT7nHroWDvw8zLhoWJi/s+4UDozP/iJWEcqh0gmO/8SssszkjvazuGi3oun6L4289lm
WFJd99X+yolpKevkdt+X9MzQEw2PhsLMvQ2YQIUqCi3eZkGdus57OYbhsFJTAd/ArxbXOMbKYAG2
UUPyMG5p7FThAnXuzPYOV4gRGgG/KoptHBuCa4mE0eg4Mk4hvnOdypigeZJgD8fFX6aohcKlTXwo
68eBxUqjcj8izzIU9o5nmOt5D6lufKPZvho4p0sd9hrC3ifI1ja4xWZYFtd0gIcXo6sadr5+r3NA
wnqQ3ntaeZ0fn3gKQJtuBhD5FVHd8bQwjF0Tj6PTTBqIQRVVyEYCo4EEvxzZvuM7ggFHtCUodQ83
KvVJnOfdZHlqE/a3+5giVb7n66eTtGpuPu0Xy+V3UUBgeC2XNIfZV+gCIJL3eB3VzFNHwcxkw91s
M22krdvsMvBp1iRJ2Qnv6D5gaH/X2rej36FlkVNPrGSFUzklfcxA3BeL5ReWi+Ex1mqcTpVEq1tc
bwWjyDx6/c36jJG5G2uEA3oXfVW5HQDt11n9iqxnfrSYhsx9gKTxSKYshdAVTtWftHpuV3XiiSEC
40CuArNtPqT6i2FV5pwB1567cAIHdz9oLEIDIsCpUvUJUh8RP/uqWv4g9U1DJECS2vOboxI/ToTZ
Va5tsE9zGsM8OPiAPc+XukoEzHmsktvKaFtLeHjS/23QiIBh8EyKGSnVT787AQ9Cb5VS2LM7n02V
MAfB6DEGg8TldBAJUbyb978WR+2Ntl8UPirAlqDvnJ+4gpN2aZWPchsER4qFOG/WeBJRiPg5WPuO
AVq2WsZb41QPDEig6e1QYdiYai+KOS2JVtpSo14rcLySLbeO4mEQEuqG/gkTFfxohxszVnPIGgEL
lgUu00qIdsUMMAGkyrmsH0Di9fceOTsB6+0C8tCnkC29wv6CMj94L34GQl8u+Ng+kaP5Ffy8use7
aFx1NZBF9Jr5oODkyzwAK+8we3ooyfwigUF00k+TFocQGKVCsZKTA4Ng1KPBvVkF7DCth8aJ9GB4
Ey3dMo83pM479FHzrIXOgHSv3jM6tI6wMXFMf/k8ps3pwRyhxq0oviQAMXJjmCW0xDvxvBqChj9V
VtBYmD0oPW1ggwe6qWdaoOPUF5EFgOEYsZw6okJ0b/TCvcs5vS44D3IZJPfWp/CiMn7qnrPMEXNe
1SgtKEuLoPwJn0MBnwfPvjc2qL/tVDeAPn6hi2F0V1w+qt3RrYWRe4fzPiNq67SiWr3XWAjPcYSU
sTOqctLu9nLif+YqvNw5caqHu5g61WVmYBuecPhsXfsSUY4CKd6eObOzxWs2mu8tpzY6Tgt1mBzF
UkpuvbVelqhSLI005O85JnZM0oP0RKRquMb2rDaXhS3nQghPgbDopNdhjtxHdyIkHuojC4GGOlhJ
ken1EASv3XZTzG2pg89hNJjJXO/vgE+WigVrxRhCzhMBkRDsT8lL4GvDcj6ICP41KUFB/fL2vPwX
LcBse8Z4BOYhzV/EIDgsHojm6rfYXuKUkmaiHJ4OLNQ7TsrK9C0Co4HW68MJuTUyNGlkTWZ5Swql
nnswxmA0XhqkZEneHOmQONn+uUY4MiLoMwjj2hsP+Co666eaR/ZK6K/toJwlMTJQv3VrYrjmt5To
ovAwiyFFvG8ne04EW67uNnvvCUrvQQTSx40LK1evuNFDuh9shZzjnyL2ZfVX56HfK2iwM9ZV4uZH
9RgtSJgC92Ctj+wFMxd458UDVztdNk5p2c/yvZwGtYfQs2hNNmX7SZZ64nRT8r4KO+Z8DWzs5nYX
h8RKnDrMMJUSDb2yYUx5HtBP5UpTr7eOP3qBz2qV2k/AExpIjtJuQKwH/vn7VZmQ6gK+ELi8O/Yz
Abdz1oU/xv/Wjv13Il+eTnLoR7sxCvo/kLqXJMnlECwzMsZaX3sqfL7Cw7+nfVVYDbf8FciClKb7
ysH4d/w86DPrzWi8l0swjECR8M8G/L1K9L7ttzRPnt90GdM9hJiyjHrLAA+ZJSUXt6D6Mpm3sZYo
14HAtU5mP7+7SOCuM5PXr+eIlAp1kluYCaxSzVLc8QaMKLSM6eKoezeRNkwsGbQOFTiiwEbFn9+U
I52Wcaz3SaCgC7zHnIJcqwdZg+v5xNKf7D7L+O1cB0mH2/XdNUOv767gLnQ23BKGLgTcKWkWARFn
IbTu3X5u/87ndwCAX8uat4Jh28s84sOY8Hb9tbY5zcN+mjKwvI/NfP2DH/ttDkiBNXZwcs9/5n2M
t4s5xr6U9YkhwHmdf0ESlk0w07pCV+4JogD3R9pCqR+Jvw71jtYL6b36n9kYr+CUQo+liK25pND9
lKNN3c/SDoysCoCEaqcnD6D9azSqVJ7ZccWTXvg/5SHafI3X+4SYm/Rc7l5KvkOGHoOs7+RD+ntG
dk8HwqxYv90YcRURCsg/HYKBa5/+qgbsBOuqbKT0F7WKQSTdq6FEXuvX9Vo6N9nESlYpalTsmn2a
I/OOlDshmWCjRtNuMWBUKIHR9GxMb+PnUmGBi5qrOTm/H3si19A4gXGma8QDhzOV9QQS8qEuuP0H
X9hKKXyRNAEYif88qdPG/rzYB+i51+5w/RXWCqVyXDvqZIyKRcta3xRVmw2V7I82q8/9nxamDUkn
H9695/5sJh8WDnXJln4MbuE7gWTts3VYZ9wk/SyvbnZRRj2+LRYKaFq7iyf0GDgjipLhOUK/bmkJ
V0rqnf9zs8UeTbttoFSawTFuu9Yb5WrnbjRS6aqLEuN4hx5+jA8X+buT/2aapKLRFx44+ZC8NiDI
pxQh/QeRfZZx4J/ImdhcT/z0rG7Reg40p47GyqmdPzu061S3b5lHT+vCXrQAUc0Xyk70zFBzobPh
+IMhcOcNS/Ysu5DRkUCyY2NGXYMFSjgCaXPIcT2Jr5KSqi/Jz1PuxkeO2VOMBklQ6KhJjGjMZ4k/
23w9qcVBAR1078Kh4PsMKRXlwbUq8wQg4Ikwo3WENpgQcB3PBgMdRsDFGx7VULvH/6ikhb4mlir6
KQLLAfbqImNL2fou4EqBkwFqHbBH80wnGPvnR7Wmk+2Ph7xl7eJregf+68I4XTXb0yPLOLFX1q9x
mi1+2hnL6AYE5iZvJPb9dGwnXZDiIj1eMqC4r2+hoa5iTVYwx/uzkD9UoqpL0vKQWYtryUFykEGI
4471L0VTLkBOMIgySTjT75zQ/Nwl17PlG/cvV667BUZsZI+TI7NH2KFvShVyX09Or4ER83sEoiNh
9jhOtk4F0u3lTcR4Ho1fL6bxkhFZx0yaYJzUP4MAdtmFj8fiLX9EeGUpctxHk4XYDMXAZdob9gmV
MgUO3dRlGUkYGfk4RyMDOJvyRI998WLdSFrRuxXgjkGzp8Phy/xDpbERY1dH5/OR+55XlcgGRu3S
p9L6zgFazVDn0PUX3mfNnKv4AC4Yb1rOluHheAJT6QCXMJszkDZpADSaCNmKp9MiHzOxj+h8fcat
uMHgFU6qN3DJp7t8qPWNYfajxd333ksV85tYGINffw+Dnky2lOczqaL+uKo0ORHLSIL1YUZ54swt
fRMKxluv3o93lEkRskXzRlY8ryYYmVP2D0k4dnHacHmlFzLbmyW6sYv/RegagGGLwj9yX6m7Ydpg
XuHEV6WTRNx7LHJFni3dqIAK1hhHSG23cA9ZIfEowqwusCqlyYaTwVrlasHsNtckdIAk5aB67F87
K010KmC9nO40ixGWegfox2A1ChQZ3Cf4uFquvqa4603TRynnHsRADMrmeQi7fWwHyPcCmmB2VQbi
Kv+LhAjqgCZmNxz3PE/H/DH2rcWSjCPE5f1SJesTPLW5dTVQbW+PjAD4Hxp3Ne+j3WqcB3HC6H/r
n9oYSkuGuyjjRm6u5xBilP1KYMsdwWZC5YNZnvMqfHZnwNEYcH/XG83QlNtTCgiTT4pDaRzvCLrD
otgSMA/+oAQfK/QP4bhjfSgKHX6qrYKk042TLS37xRaAj9xQ1GY+fGVTTrrAPEMhfE/1v2/ugwxQ
pTsqqW5wNJL68pJ6QxsURsXohPXaVjw+nbpNUnXXS6PgBH4FRxfJI8M77VvRQ9qlOwqU9i3jxDcA
lSTBEwa+Eg2WqECdsbalQY6XxxqYx3YYhC5j4hEZ2HpoVS6NxZ0q1+le/oDEktifdKWRiAL35SiE
NWf9zQDtK9gRSzizlbk4bjYHizP7mx1OOynxi68MaJMOwatp/yLf1yhRSpnM0UbC2OdFcugVhG4h
t/Xiuk1kpnS3wJ8yrliLlWZLQC7HuYEP+aeEyUET52ks55DCMtceP4V1ovORecLjWBCCGQNVkdmG
dqiBWga4XoKbD2MiPsXkbRaYY/yjhoFkToM1rphT/hDoSnLnrKM0xQ9B761oYQBhfyal1NZj5Von
F9wYD5Y4aH/a3Msy9t4ITevWzP3lXRi+9J9wtV3h6XbDL5m6iXF9ht5+uYV+qQRPgHR9QnNytB1C
6bbfbs6GvShDnK1/YTrCUAibs7Yq72Lt8QLbnzUJhwKCAOLXCGpm6Xz4M1SZIM5H1iziKfmPUD/L
gxjJIUqKD3KcaFdt6sDrj22YAazOHN07WhcGjMFXN+RzXZvjWM2qjnSkK1hUPCaFiq8ibGIfmSvH
83G7PVL5ZX9/1IpA7z8fTD4GXQFpgp39QxKlsbi+z5dhlYPGxQVfoZkh3qsRD0jLqhsAGX8WvEyY
nbTYI/FuVd/1gR2w+wkeMeZv6es/iMb7RJjA+8OgZrCb/+CNT8izi6uxhbVsuCKjHxPQBY3UH0pA
qQ8+SN2A2Sv34tLKrBb6Q537LNLe6lgJjHorfRc+eaPFaaGS+W5r99d/INPXRE2ZjD81ELhxoUac
hbBoid+qRDaL4OtbZhWK7olTd2bCIEYx/xPdSslMxG2DtQiUvJonTa7ixqLRQd2E5dTZ14+QxRMY
crUMHIJFg73jwLKFytwklWXgGuaXw10mBSwWs+7C8PezF4KGwT8EBSJyVx7orEfyM/wYLqqWx9bk
HTTEkoHsnp4VVn4+YjDAZmb+OyJcsMDb3pbiFddtx0lfEu189UI3mZXfvThfSHcLKGD0dErzY46B
2ZPUgErXtuyOPm29d6UQJMIoDqTo7DMYkyLNgZtwjy+xJWOJm7ZzJQZqQOlOaTIZt/aAdOZSzqqg
myxBEYTL1q7uB0LQM5EwZuGQNMvJ/LjU+emY87Iw+RKI2azl4OhOexj7HflgLkMaxeajbhrGjVYl
JGqGlqEaJvi8+MyV+ps73RQ6+mnZJDcindPB58zrLdVEuQdYPKc3d3xmdhR0YbsM2wEwQaQsSlYE
OctvRuJbTt2yl8xg/PrN187aV2lX7vtYlw9kT201ldW6kJfYuP8lZjtBckVcdpGdmzPsIxa3YSdZ
tF4xD6BFqftZ6NUNatSkjOYc31UOaZJ68H5udDGt2yuZ430pK+52iBgXARXILuSybx+a1+GUWTjn
qXed02A6zLGGCv4uEspGif2cQ74oFS4W8SYzELh79SThmqnG4ahkMYDHheYb6npygP9iW/hfmrBH
9Qry281jUJZo7BUYwjgExRtpEbjJxpMrr3khu4Z1wRB8XbYZClFzoqcbVhHtMOSLjjzxXlnHvynV
pEM9JeuaDdQQRDS0gjwUxqWSBh3Z9PzEjWuQFk+wIIeNuPR6GDBOYfb+Bh1lzsWBbEH0p9nlc9ZK
tP/d2KC9bTUxt0ali2Eiz+rnncOBB1Tsseg2w+ZmYFS+ESV22Z81R6X+YcfFsjeLnR1sm95I5w6P
FaBXBOrNoeQlUVzym/lhUAjb8F3Ye6toB2AQJwWy7EjJkggO90ideeh1ThFcEp9RQLenHEn6o8+f
tHRWKTqI4Rpu25mIe81K3T7rvDyDRzzEjJ0t+OV8sYDyExLM7WTt/+obsAWjK6lYja6UpgM2BTcj
wR2p7T6dicFBck+MvIZi6xZW1Waa/truA/mfqJ4iOqdsqKioLN2Iz3rMF5rOu9BiZMAR9kWYzGHX
u/QrdNZ8kUYUTtR14fiAJYogbi4VfIsdSPfgwJjZV1ARSKiqbA7Pp2n0teMXyObZHQYQLpYKwlrN
j97letEz0tcSJ+5PCXZn/cqlJxmqYrVQR9ZRRhpgtg15xGwg4cckonPzTr0x9pu4ADf4nAjjvE5H
ws58P842Oy40+qNahfc0wbXAswFSVEje1J+d9RuqdOmOVDfw1aLIuOBlIbxlx4j1Qrm/ckbG6bhJ
x68XW0eM7H/Fa4DN4vdRYCuSM8e1sfayc18fGCArxELp8ITx5VGDDUJ67cQ1i2o3GKi5q2TbH3v+
xsjKcXCTOS3eh/bSFauhk7KpdeioAtFyMxychsjjT7eD1xY/57uISeLKI5MfpwZQpb9Q2bJyNGgb
ulJRx6rdPLBnkqvjwK0KfTdEfdrm5hrXkw5NMnmWACoh9A7//xdmfFXSF5fyNcruw7KNYSQQYAy1
cEL6+rKaCht6X5D+xf6yPxtOlUG5c+PP349M5Gd4r/HTyP6YJawvwp74AmIGG509WjX9QVGZCE/w
MqoIPpqFJpt8QH6IcwZGEJ6gj2il+7h2CnTVcCMOvrTYl5n7sCG+5MRpmlZOncThTbYEZKTPllVp
VhkeP7qfg39nGEvYpTwWzrkF2vZ/wI6LISyALvLrfcwLLKD2bIrAOeppQMG1Fve5wngE7lIxvM3k
8dS6plQFnF+5aQg5d/nAa54bDR+ndeaGWmahwSAAmyZOFyJnoJe5P8PP4rA8nxsWGFEMNmRt1t6S
VuCr8KRK313EVkaZKOMRYuYkaQESTJz7ysj8KiQXc2sGH/RfGQGWS2fO1/PG6piZgXMzL4NqVR/k
FKzv4lfghgCOAdSpkkb35M7ojlysqRJmFcghJka1pLsvUTIegCs8Ezn+zsqHDueiDrXl9u6Ch5KM
O/7+gADVzMiSWVCGWaq3yqSYywyvNeqNxdEBsBV+m1jZqg8M+8O8ssj17KKeyVunN1tXHcuCx762
gZGAHhnY2RKR/Xhrv3BAq2x1tjaUDu6eMV5OwXWQMv2ZyiXPMmqOTxcPXRap2cz/HvQczsZ6QZOu
asj4qYKB4tvELL/yknA9E5T5GFZYKMu3HNOIAGyNjOZylz4bhzhDep8wrpmr75KiRkHi6GzuexOo
kUpDhSWgNu2ylJTcY9dEPGHCbAJU6vX6q1+JTvdoYa4QBpuOY1kX8MWicV/iTJzS/vb2FW20V4X3
hu3pmEMloSQHLMzELDNQvt+85102X5gMshQOMxGgD0o4hCNm/V5kIWop7JlJEM114U/MYlpzlAMn
PAM1I3sLf2rGNXJGp1OP6c9DEqAMKK7Mmy+d5+nE+1VB3xqCGHdofjEWWm5hNUmeGoblVXEgiIqt
s4KFwvXgbMQfv8eNDgC5tFLD+4LlCqm3kaGrjneJhQfjtyBx8WZOe47QJiS3OgiQEXLgjyWvi3wl
ivUqQGIRwIKPsx/xgyifY3sTNnHrX3tnsrSHP/SGndzqpMQqia/Jafpl9OV7hCzcwHI0tsNLlYQo
hqgb3mRdSahXj+Brr5S5JDPTtTh5pAZ3cLSLvXW2xd7fAaSYf7k8zEIFifXhAOqFcVeb1FSWf1bG
nLaLC8kfgttXcxR5vW7KCFZKLB3C1mgzEwbb7TGJxHMu98gAlg6pouNPABfIS/9oF6T7eUUzzVK9
qFRlJDNg4gkGETXPznMmN/c4o/6Tdr2NE2ZvgbITzWII2RTgxflyWl/OXZIJpm8NeHki3PVVBuRD
YuuZDAR3WyRPZCrNAAaN0+Jh6UA8YaskpYszbmV6/i/SrFxqqRdtpi8l9acIu3MIbrYjLdQuEkDx
V66hf6M0O+CL+yWf+hi4jSxPLfCPkcQw+Ha5HUeW+SEG5f9caueu7/e1bN06iAoIuHUmXIT2jDPB
gxicc+c1B8h6+ZnM1XhwxCmIzRVY/KM8oSZP8isM8V+rowWL53RPLLHO3tBdkZDODF87VUUQGnZe
Ig98ZMpCCC4mqd7KcOexZ5nfRqwiVX6WsUf+wBRW2heNXl+GbRPdww70Flhf9ZwjSeA6EQHdaY+O
0w0j37SOKfimvLieHYMOTqtxaz/aB8xcwuJUVd59+7u6HTcKZB9T9C+yI2k5aTBa+Pv6WP1qwTBR
d0dBVn624PodVYXXGvfGq6NLSK58lJPKq1R/EHPD0n+PDXs/aTiLfs0OvHlaGFTqel2QdVoNMqUy
sAcSsA7HK7/yLzlLXzc+RtEFL8EPxJvGVl+uA/1TQK+5JWM47tUfq6vJ3kq1wm5ijIcPRhPaSO1H
1g7ib68n4rVTPTz3u/Ct8zUWbU3G6XekKpZFUaMsTEUVIV4O/Ak8XGmLTGy4X7jrFL2FO2OFUqpG
FP8iJp17+xWKTSW4KZHnL/lMXUrteh2SYSOS7gU+3cHRIYg9R3E3/8kBJ3KDoXJZU9mm46kh46Xt
/6818UAKMrkdDwH+OXcSs3FuAgnX9/Z9LgHIE1/YMMF7ytNgJxiKRZV/7b10MgyQCOesKzBrH/90
1UQ00hSzkB3roAaCxTfYyLi+15V8h/hBNMJxYpCF0P5iyE3GBq83jG+4Ra0PxMV8uFy2p2LmOXsI
VFZDCpV9aHpMPnADHmTskI8+o46lY1JDp4h+sWweC2/BTtOqQSsGyIsktDQA34UJpFNwOCkFUfOg
lXWig5QYUbaGvAkh/tUYxbvyQlamDZIBMc7m+UDiCE6iBD8/iFq/Pya1g+m43OGBwWRMntawQz0F
wRQrQhx+h05q5jDM5oDcoaatueL7ZqvKNR9fNCyeRm8XlNE3hNdZj2ajTGPPv3yLw43+Y9izZojS
vpLk/ywmvJ9dSkNRRVaKoCKtgLGYPwBuSadhVEjGRUCGgU4ElAK0d1Jh4UrKE7BR3cOgiiO+/tPN
G49eCJ38Bsxww/Cdb77+WrLls5dmBVbujJj3TR3//ZuqvD/VNEFYp0wKNLXb6j3Ar4b35PSE/ose
z/ZZFw6mU6LdN+qQ+qxHadoMrPTM5aaADYP8EU5a22ej6WTO9niJpYGtLSXRvzqfLBNBzIKNHdAA
jcbBJd6gNNzrqAZTABoHIB3RJ06v7N7O4ZDdITPsWgAzo0IdtqhdNKhAuQZxWTTIbIWEEZmvOq1w
wYjUnllCdgr8aiYXyCOwpJ10gnEZkjy2va5TX6o5kSslfa/9UZ+41naxT7ylUzv2pq8hNvi7jQq0
Uex3roOAYU8C4Qe94g0CVxzHSnA7vwUrFOCQsLP4slqz57RBbix4Q3MntZJgiGvr0GNwqrCwx9zH
A9qQGBV22swV2+yay4+V11J+6rTZUUvRtR7ikCQz3P6nZeW4Jz1cpDWQqwx1lWjJ7MVFO4+O/vBk
R8IGiPpQVy/vIEnHYNgZ6tYgfm94IeSp7jULD4i0Rb7fjNumQVL6I8LKQb9E2Vthucxi5lWMek4x
rR2l9UKMYAOFl+M6wOFQueXzI+hjnpFlTGfvxIeMdMANFzk7VvUQfL79O/vIs89AClX6N5kKIVQH
sHSWeb3NvLOirZU2YTLvmMu5o7LDa+2xYtAk8V1oudcZeb2xkbEu1zqfzjp/+Ne/wh1CKJBbc7ii
w+EvJEndWohgQbMNfEdXRjPz07Vsk44JIPF6m9Z4svJ9Np5dJODsodSD2ti5KqttyszKaDrkigo9
qvf5RltDbw+/hvIe03IO6aprqRBCPs1DEIVzTSYOOou+ZDUNQxbtUhVAR6SLB/nwwAbG9+BLvve9
xMQVURIEUgviN6lTb3uowErPFotUBNU1nfmBrtp0jMRyZMqg+S5oXFpeMOMxMfn03G9J13Z5oFbz
h8D8/tx1/n1bDjJArFxnzfJzCWzIUxLF85GnwRUnrqNFQGvI+pCsu5MVBbhaTg2Wf+jmF4nlvNUB
eEIp3FyfaWudQZj/Cr1R41GBI0H488fbCT4TeEWSF0HcJpTYAlT6weM+HK7+nDQ0bG0tXoOxqUaP
hfdRpOH7pwH1Iwon4vmM61I98ZIfPaTXCmHXyc7W27xWm1rth4GxevOC1SjSaArpMh7EY8rcmwQU
rp7Bse9pNQN/pmFxlnOKBy6lx6j/b410UBtJCs2fVRu9YVc/9JJPEO62DZvAmF/E39v4AnJ4+Wai
nA5AOlt/7OH9VwEF6OQklkMRVZNyVGX9tJflwdQ2ho05g4iKNhYS6ImAbUEtDkiR/syUgh2kRIMd
+6NpTAZljHHXYCqyxP2PfxyMfPIApcMEKhBpBypw9T8EtgZ8Ah94Oij4tPyXBktgTJE37CgkPFIv
obe+fU3NO4jApYdyEswwv4hQtI+pbCLcUiEjFVe/X0GxjEarpkXnW2xRmAeGkTY05Ay96EFMYkxS
nXDZaFHHBHigelcrbJNnHgYq2kl4Z+GYKv0DNGyGk5gmQNFfYAlLQLHgrmDPK6KOgFpNjXItXPaI
6mqBvwiyvzT2JwVVsoJBMRssG/QzFAz8hZyTd9ycI3/5/CMJjy8SR61bylefbOb+o2ZfPxqJaaa/
k9Tw1r4EpOZbyyV48szdZ9ofXCl1Yqw44aISljEZCynJmeVbK4E55cG9H+zGpz3m0G7TR+Aw8Nhq
cldNqOAUW/zO55jkJ+JuhoSCIb3QGqLOKoiXcK5WqUCscQPtUIfC3AlVXEbjcuQ0zkr3hvyfDnqA
mZBT0MvHIZDGaXm4y2h/Qe45WtQeBTwcqcoZPgpvQr0mwQkm1+gw9On6p60A/NcVyaIIr5rwDTjL
ORHRRt85CKs5ProKAeCV1VIbteNHk+VwMr6kqG4egTMv3TaZ4Ammu9oiCaxb0n/dLgC/V4IQlvIj
WvW2aIUEPsvIIugQmtcyFT4/+/Du5raq+/xjlGyOrK1683XGSZx7dBOScJNkCLSqT1s2b6E4UMKi
jpwzVJXBgmXrlvAKECeNG5oW6yw8t4qSt9DeEXOzYr/S9jTc14YGWa1dM2FVZKKAudY50nnQlMNo
FYDcS5c1fmW4+LPoYjy4QfRyqRQ8aiWCP9TH9OghnothPv535a3HtLb302tlr02u/hPgiznoJLJX
UVw8ur7Y1O3DXzajcCiXBDKV75UjqtklfC8RRCT0uK6n1+uuaXt7q4hxzKWo5yS90vAPFXz+bvkH
H3imBykUVpmilyFCLYQJnSRnbW5Nk66kNODQ1AQVhBq09opW6DClVPu7oZkynBjGo9wiOqNsjY3o
PoxEIdaKQBSlwAZlcn7ZeNYUOHuguotv7iHpjquSUueOcr2FVR8SYYPkm0U4/8urI5QC5pnGQJN5
nNypoqBjQYUr9/CpThmGC4k06QdVQWIQJh2aJs7hF/fECf7ntkwsTZHbk9eqMQ8G+e9rSVFV9STH
oTv9IGcvKvSa5vDSRAOPGcSB+K8Uu8Hr6pDgYhPKf/MOGop+NdeBJs2P1Cgs8idz4O4hNyGxNU4e
d3HQvD3C2YQSwKmbGb92DbAARHMvp8B10q41Ydq6n1S4O0oZ050lbIAqcBa+BWVVhMYrlVat+NOs
MUzhU5DWjzcbLFQ/bF6OgE1+wGfH12dM/uVk8814UJY2KEE9iToKx9OliMlJt1mewbHAylcBICtd
t0NPBCVTsnjGIjIgzw5Ivz3VLYcBW6wP1pmwvRgRrx96NVhQiuQxQGpOVgZEMWlx+RkOv+IjuLOc
gi1RrnGrkunnlVpzoRtIkqT8PEbCyLCjMD1SQkuU2W9PLY2bGysyWrpcL3QcJD5Nqdz3ZVvX/GaI
MEn5GHumOwnncg1ynr6KNSf9+nRk1x7W0dtEEJsji0n0/aJrPkfp+bI+wZ9uOo3hBWmfIjYyFAab
P2dRvzWCjc5kwjQWCu8l0bvIasGcvgA9HrDDQe22U8SWa2bdpKKcMhkGwGDRVyoJzN5vGT7qNv5t
Bz+xDSVgen1LUabrk230IYI34LZvtCjjnIYeHrjGLqwjXx4Q7LwRrBWk+4a5dL6su8PHaHwRNp/c
LJLECSBmgxAtiicpzMw8d+cxj57CmeUgCCP3qWXomGkjjX0vrdyulSNsS61S1oPo2CoTyz0BjAFt
M4LdNbsA5MZIkp4FjUW5r3S7gdhTRTNu5zzURJLNt3gsOWSh9GgR7q8ex2nk0pGEoLBXcKhZiIg0
f3eUUr81w1k7wYHlz6UAvJrYwa1CTaKfewGLNhki5e8SIPrKDMTsh0TFd8TZsBcAVKJsBceLbraF
TKyuYdhwYj0ENn5dy+X8CJxQnxqOMP001jpqQhZPjJhqc4AWVm2684OnIYO9trF+P4v1QzXgYDuX
Z+Bl9//ukUCBJtXxgDgHzQ2yKeU2xu4tuHXFJ9SHCZvu9HMYFCuQThCMFbwdEv1lJ4myOAeoz+nr
Np/+bmvFUDzA85gps9XlDcfLiOwtpKtkGSK4Jd323FIwxxxHupL5iVFzP/edrklMjR21C3wcal8K
UO43FUCm6N/5tfC1bPwlZvFgzsVuZX+ZJ6Wmn3usYRLs2Btfv0aeAzf3OYywv62VRjOtEF0oGGFN
hHnRzEpSzSDMOykC3X+KC8+sBW5xhiUATHAxP6wZWkPAa49KJwzM33u9Cf+W6q/xsYpOcWk8jah1
tQldZNIkMkyOBqmJIj2WiBqYh4+DxSxfQ49UKdPWwaCc3FulKgU0VUyVMcoKMzvvP0ICr5lB/ZpJ
MsQbRQ7FLTyEoEAjUMltFXW+lbp2njZg6nFquM6N2iDgE2SmSoJm3Zry+Kq5VgjrNIIt7007EOIR
pIJ/FLQap1b505qDCjrgaVLTXdJBEr7gxFDEutVxybfW5IUlWJw/wPHef/6j8YQCXkAv7USVZeL9
QyT/icNdyR4MioiWh+uF0pKQg5E7TpJw2HEn5D5ARh/L+gJsfyOrY06Y5GNcdjbe6iXZncgSVaj7
gYyxkPCoClxW4lSKbXZNlCn1tRcgXASpiBnL+Y2emW4l5rZmu9ESj8gMzbTZ8V9zRZGyIy27K2Ol
5eCqdCHu4aaCcXVP1NbTw8vf1lBProIc63oDarRXWfMrg9l6cr8XdtoBVquuKWEYKlTMxqBLjsxS
ww6q7iNIFCJU7gYSqdu7rdiLi/1Hf3Ls1BTnNg//s3VeQqUpFG+B5HKkwISB0br5MQ0BqBLCs/Ee
YChW+wN187zQqBgX+icsnYiTQid6cfJLScNCoDuY9aUlOcIdIfJUrUqiE1ZkXEToERhvWuts4mCg
pZxPTwnuB2L0FnoI1AMRJoDis3/l/l18Y+hSSjQNlHMZ3vKKbf6vRfr1JebSqJ34zkpdhahvDfKb
xGI8Jofe2kZNM6mbUt34b0Pc45aM3UGueQBx7eFNIlO8qa0WC6/7QiBdo+27wV0N2J4cDfcP+l6o
XGlzibbtw0cAaGM9yZ/P0qo8qA/klf/VzY3WwxLh2jv0u8A6+CtE/HSWwWks/V8Uw0uUVMG1BfLp
E4ipFVK+aMhKGK5k7kOVW59JL+cHqJ2tuhOg1AGVOrI6iQfuJgxTEMaMqR/gHP2myTxF0pwkM6dP
cOejRwVXGveFRC7fjkx/aiThC65dExA6EX+8eIzV7mKBl1CpRhJtkRTjOE95vrA/DIZ2uGIxhBYP
PjV1ht4GDh2q60eOyN8GiSAO1eQhWZQrzfv3/QDbis6foQ5FuNW0CenLEW1LdTaY5NeiIWpPSpAP
SaE42h8XylLSTsD1Dg2phv0pBJRRmK4LFC8+DrYptAy8H++11N6vt8HIWvNS+VLBL7Z09/DIaxIg
+Rs4avFW0lyRxHDaiBIJSe+zpR4ZZMF8wC7NVVbW90MrZlTY82eqTA1TBAAOsdeIISGUEv+FrewQ
8ELPRarGYfC7PajZfuq2HqrEhM9OQ0Max8DafjFCWnUcrdi713v0XuIYLNtAT/BPQaty4/fimlLm
0JOR5pQqEr4ugNES+PEU4rclxK0AE4wqiQPYvDXGoa6sn+1E0w76Q8guXGxBJ5OOtftZu9rrcqEk
d1tQVJko73poWkDvW12TMHiHTM5fb8bKx/UHGQFn/A0TGpAFED5O5QDlCXGeHUafs+twWN99Duzh
ME6Y8CZ9vrWbvdEfPCnOVJgFr1qRjHahrtGfEqxVhunRU9GQ7XzSo7ozRo/5uUsQWLqrOBKV9Mdz
SU+jYXo6UyHlPnStYMRER5GqsbW85IX2dE2j3sX8SBsr3/Smsv0R8EcrFoq6qIJGpby52tIV/EdL
Am88Azwfte9pg7Qfs7CzxgYDUdv8oVB+MwgxH1jWa9dpzaAp9SeZ0DTdsNTYmHp+vJcC6OrTfs5S
ITDE8/DEEOM3uXQwSYEj7VOBvCiUfZ0IuVSNVwdDVBmS0RyRWP/4q65lvKS2vyGKYHmkVQbm/2VC
emd35rhl9RMlgnnKvk79VY5VHyiU5bmJ4WGTlDuJsb73Fl+Df8D+6J305zqYWOIMLIbRAXN19W87
ei55nUp9yYaUEgmk0ckazqjaV7YSUfr99ZaeNZeVSCvREU8p7D0cfJuv37dCg9IlVhycpL9aMs/n
RB8MZjRA/OY08p5pvzvwk3pFEFxnPhjL/FIcKFAIfxN9+Mu05REraKD4cs4FbWltCjVZIeUFTFGk
E1vTTYYOQxnNapuiWtcDe08HpSKtEW8SGfXNGQYiBlBTvL/pV33Y26yk3h22EVtgTkOXYFD9BS+A
4xt9La4I2niSA/cIfvrJvj2UGWTcrSxEMAAAG9MAE1Q7priWr40wxIl7yJCO4lM91OmGMB8AOefI
KyP6KI0My2CcnJURVxi5eKjVUUZuRZoTK9tOQ1u3ZruGuB3xyDRs2PdZD6USF0sD1P70McOB+w+4
8wOVxqye2Dr9kgOvBSGCSJB6ZbMDd/m1mhcsR6sjOK6fhBrjeusQJW7/IZ7DdqKKAEFyXLhSBhjE
aBjgetLzLGdyRwTdDAjtC83nw/BKwKcu88uzsURL9lBQ2VfUzQ/hy97yGR6UQPd0Z/w+CkIFyNo5
48SREknkryZJiRXb/6zlpSDS2K8Vz/yIk0k36pTl2fJj04BvUz9SsKTQOYV/3rfoOpm4aVCYJkV3
dzBvull3j4ZznGWNj65wLrbVHByXGVlWwnRgpYvwieMu8f9JtuphhfxKvTvkRn0c/FncsG30G8uw
dI5N8QiuY8vt2c2prxCGySatjAW4phh9eRLVcOTR9zxT1POKcyUgM5LJjKuQJZgy8oE+mC6mN2rX
obMoEA9arxwVnSP2mQaNuVP6o3LI4XSB45444PTtF9+y/9PwX03xplJa7eyto/D35yubQsKB2lgn
xkSMlYyiG1KVqFz5ZR+ooUpavXoh103KPOY++pkv9Ap4nQJOrsVY32svhYhL5BnstjjpeGTPwVI1
WqFPfq5onPDlodyxJ+WT3hsp/+I+zelhm2NAN9AZNYoziNgnUiecslagdccalI9OuPyg3JjhcsGY
CbyWqlKDvMxEfiS9nihJsC6nn4wCTTy0pTK4mFERH6zkn17zCPMacIk604Vxv+BzLxuz/HcOoZpW
UmcuUfI35lpw6clCW8fCsf4zB7uRbxjMP/eAteSrjlvGgzZyYBCpjxI5t6aszJQrs9Orq/Nn4sOe
NgtIE5pyusI8fQHACDhXh2shGKmsAyIhXEMQUVEXLRXRWtK19+jSPJa9ZAJYmbZhbsNNeOCa6HVP
DZPcPFfmyOTzIyUGJmv8+m93H9NTT0WTS4J9wKvQ1XBZXu2V15jeju7qiqaPp5TkvIswN8LbOZXc
ACNEvRutGQeRzsZiFaJu9TDA1j06lAKZSA0FVMJiesbQkfYY1iwreFBBQbWWvLjP1EbqcyyMzPXa
qH2grvxt196+Oze4GAVZMqDE5xv64Fvu2YYHSgUaAi/DB89dD7g4w6kaEESw8r8uuGI8zhaPv444
E7iTZlsd3ipCoc6sH+xLq2dskS4AnezQUD/HCTyNwXcXY16iltv0vtRx5dIUCX+gNEf1rJHVDQwS
kefwBqnpTugJ0lRJBGi2W2BqueCgmknM8LeO21mrC7oYMZzVrvinRm2cRA5nYuLq9sa7mQd1+30p
HsnzYJYkziNnbXpmeZEYhvHGZzVOyTs/v5F2RQ0ow0yQAQzwAlyriUSS50dfvxVTM8wLBsEP5OBX
HwjJ9T+kLWH1b0a4KHKRyc07IXoJH/KFgKXSFlTB8+9mK1QHimeqQvTsXKdVjrCLbNrkZDxvgAUt
0HNGqbmg3zdBvTbBsFgmBA6O+Ud2f46RgaWyhmzf5dTusRQV8LjFXGz6lBHal8jLVZIPnC7gFi1Z
3YYN5D6xcwEHVlYBHJberNcXrsT27hXFmW5SdzkkWg8oMmrid08MjgIZIWdnKEPnc600oRv2J2EN
t6qo0V57/+gxIBxBYO2smpQUcEUW0QILpeC71yWxZ619Fcjj/cdFiRrj//EmiTOeC8u23t6KO/J+
mjKdJUAQ/29LFYjkKsVYOj1oPY+3lfJy3XR65C06MaCn33dAIAh3K+PHD4RSCGuw96smwf6IEKan
9oAd0QFZOCBKmz1p/0dv9qxeHyWv5aHi/yik/22pXAQ73FFpjUGetqxT3Qqr4WuWC+DeUZ9LhHJ4
QKm6al96MSs5LCUShy8gzxef4zNqumsLXHOd814TGDJcwBppSqjtpQUWJcUicrCIU5XIeXgL31J3
gUG01As8u3/sgXRoa7y1oE4YMds9/PKNRmNgkhred25HhQEJBalrbstb0h65koMmv6ObFhnTeb0D
QsMR7FPBM1741IYxXrfFVcnTtKq7QTz1aDvmOmuz7zp9vY+9u+uWbeueyDiqie6OaoHxePMGrVJl
5owRR16ulQBffnYWOHXFylIE6HODwW5lk0ypUdUTX4DfljNWcdCvF0drXdzsBWYhvtdx07iuHujX
JXL3BV2PYDpp6Tchh2i/BDmjbylJsxUqfShE8EKZ1686dNWX2RyPRw5+USkQrl21HzBoeuH0wwnC
AdcC8ZXbsiA/C60R1uQu8O1JLfvS82XcptXUgaAtdJrDVfXFaN7+kwl411PA+N0cdq45PpM5jsLJ
U56mT6EMDZAqs7xn8DykrvyoJbZw91f0yOD+9ULyS5NdKIJ14q29f5+FDuRzwH8G3v7Uwba0+IGe
SbRxNVhiNKS7ouz5ogRhVbBFr0Qyox10YoLsTwWwOyXEFDnkRrRDvOkPXUXdf5HB6U1cXyxGRtIx
gQ3KzlvbV3XFmNjB/nYoqv0BrTc9AcX27WMz9xCQXNroutDk4mGSELKRQohWx4tTLZABNAKPkFhi
4HT0+oRW7UTTmH9tQhEkNekQp251Vn0aos6HVBxgEZx5ePLpBkpRYiXPEqFh0Ni2PyGtmuVb2WY0
QOBRsI/jW+yeiP5RuQgGG4QifNYrO/jNKCTbWFHrBIkSs7nTGy778P0SbSErMFQOkNPWngabO1yh
LmOINVphTTzHSvd50kCStIBlCaFDY4E0azBtf3cNrUQcXhl47NQIews6CZEizBDryfhwKCPk/glv
NBmtE1sxxAS0bh+Q5NZTS7L/fjd5NsXfsxGvc09AfiysSIdgKg+QGiwZ2fzU8LZK78IV5ZKBh4QR
TcGDCfj9MTsMQUWw8pv/YD/r9XyeKv7pljakAedk1ae4C0EiK08rkrppDKPNUy7W/HoqEOXcu5YJ
DbtX4VFBx+U759mfpR76aAsopUlbBFfGpbtiKRFyjpzoab0NXclD00qkE4Ia0O/3FonNI/vcHYKp
xAT+X6Uv+6KQp7LQ0CzP+naW0ynvjxKRgs/9W/WDnH5GHxyR7hjdaH+seZHVZYS6cE9RTV1OiF+3
krL01UxVBaoj05zYpL6KKq1wDeQzZ5TR9zM2Lyx++P78K0+YEjzWnN6LlJjn77qN+J/qcELTU1RU
dRxX2f1qUR8SaRbEFJl1QPcTFH3CM4w57GImmiVSC4X3NfA1JuqmapTv5VefQa3xz2ACPr+bjeKS
Ksg31ezMBj4uLy1/AOwWMPFQbzFrzog5QtNaDkHxrVux8j0PUB26E0tQ2K+xFIlpnqSuZ+ayPDQa
I2+8mOWUM84jYzwj3Gn9tDOqq0eNfsIIXYHAWOrQQBUgv2zzmI+gCQC4cyGUrbP4kVd9kwKLypsU
FmOaeA5TmQaSZ2bg2ZokoUbodGeAT9htjDtDm/ktigDeJefzZb0zLkcWPboSs/cEZNovok/aq8zi
umqdZ5Bs38iJ59rEq4FjvrMAwGQSRrGMliJX/bpp4g7jKC3fjnmA3BDc4QJ2LbsBEVFwhw9n8Shb
tMIJLD5G3hS1PS3qBJQwIC1oAq0GqT/DBSZW/677FgeLxonS+Y3mDY+BNTZIaLWnve1rr9SBZnL7
vtDROZYZSvogQ4MIfNdo5E5Z2h/sQyGTuBvGEXlTZdKaX/MYDbukNYF8TP2E3jjpjqw6KiRNarIX
xwXpsERROe3icou8XYcfxnRbXCYh8YOlFOaSNU3wROCmGf6pvNV2LIBQb80QlaS41teYltsYBNft
RaIVy1954Jctris3jWiG7q5f6IW/ZyGhZ514g1OiJ6jYSWvfImKXjTLlfs1f88SqYHPwpKG1i7Hm
hohihIwrypvymRFKnyn63V0NoCc+3fkFv6lZhhUSUGW6axq2PsbJV72EiVOkih5xcopXk5pV2Z5l
vgo5CqIWrflF8PhIwIdKbBnXwPLnxZc3gYvwih+ysLaSPsicfQc9JVv3D4bvHe4gWpIFB2NfMLma
j1yd3ZGOFm/iQPJcD/ThaNCBz5Iqf8Lf/bQhK5O+g8kVo5aaCuy8dBrMIWv+qBPQUQQY/vXUXFo1
iQ5XuKsW0v5NM/pdtyr+68pWxixF5WeF1wvpRY7SWpeP0JbwrR2RNFDk6I0S/9BxdrVxM+kvglzP
BRjx3cNpsW+aZw1i3+q68G9tN4DKo1ETqWyde40C2fIEq/tvTo9JbuUrHtGSMMfY2KUVu08qcGt9
PbanE1/LaeiaDGNkY95KfveLAQvn86954JT2Skf6xDZ1PwNiw+R7hGDTvEn/VABqYg/iJ9yn9yTF
tgE2l7hzuz1RTFb8+/9Dk9NdkWM4Vz7i8lvf28/v1U6BvIQtIZEEaOrkMI39YPLpNWl7/LrU7sBx
g2OT7W1jSWl3OnFNViZ4kXwvRmHO19EqhZ+bq0WMANlMFVeRPeYcA8ROIpEIwmaatnXYNkkejWio
Sm5wMQIsQcBAVayEsc6QVT0SoV8dHe86kTSTHaXFMniQjtqvmRZmgaeo18NyyIZu+Z0DCuuwG+Oz
+9pZCI7aOAx8K2c8j9qfIfzgnd3enNdUEMQ2OJgx8ZnzOJaVtP96wokrBBeG9LsRjh5Tan9xXcBo
YZmAzuYXKDSaDO3X9tG/JpbGTkTjNVq3lTPEMy3xFIYDuL3hhXptWZo/cloZPkWb7Q8tquHEljoU
YEMC8dh2ryppvcI9qcs1TveChJY/usZTEEenXCrZ1XINFmz1iKS8Ta2jApg2V6TreL0pJodu7oHR
z/mFI0yzrwbXAFnJ0IMl04yHHfDlzcGaWl67adwUS1UVBQb2I+4H2oTIHTtujc4XPC8MgGEZ2Lhm
AfUtMLKGU3ze1rY9iirYmTdyDVOBmhYfOpeXsUKvyvKwwzKCeApRIuyImqXOxbUEGSMTyXun5m3P
MvLu0bntZ5fsFDEo0yM58QUv8RCybBNaGjU7YaVYTy4AXKku5b1i2e13/B7LMT3dSP8hfgoDx/Ra
su9nHoFyM2hXAZ2lZRv18FFpOSArBb/rN4sd8OxfATX81GUzMI3QNeRMRqRt5ru39ADSE7tkI/Kt
ni5tSvTB/qElfnaN9TBTDvORh7Fyoh6DGpoFzbFHMw3P0RnKSSLnGAm4fhF5CTCb7ts/8/o17KOw
+DgXUdD6ZqpomsDG0/37paNiZCZA4/dym+ygIcZ4PXa0juTARGDuYThX9yRVfjCh1e9USnoX38Ak
sPtwRVj8lFtksvo1oKBslXBf/SPUMzkMIWLMFDuUbkynooOkbT/7PVPqSdw1FHfkLpWmaM5/JfQ4
Prmi6VyQhu0SweTWCKSuj7a71yOCNiJtzoeLeUQks52iprn1b38g9aKf09Fry58QaPEosbquk3LA
DJzT82AWeTOPEskBL9xjsgL1XBjcqtZmNV0tHy5gzvGLja6X0+DFOiGBFCoZTUtIyg02s0thZ24E
p64I5VTbhwDg09/QinlFfLAk8N8HFshcpWwMwmWGbbb02QeqAItA86+gpQfHIq95B2zaiGm7Jlw/
9c/H82nUVgubbz93MGnT140rHeJVp4JQLXn0KwMNVFbBBA6E9NLpxBmBhDguRtZRTqzEAT0bJj3N
wvee5S00qbnQl98oQ2x8Jq5nS9SIV4Bsis2vDwNhvan4cYJlZQQlkDCh8zNndIblxV/H5friUYXm
noiH0Y54kLNAVqLF3fLENqRLR46buV8VdxJuo1vHxNXlYtBVQ9TTRJcKBU5U8EdlQeGgIZPvb015
ar4IHM18+KwK7k0Z5nh7gxUrtj+nRxZEkbcJuTwZCXn3H3e07d/4tRmv/83WXiM8z63v7FO6oFJy
DGi+8UfH8T5f6zpZ4LYVi78VmcE16t3diNrWcgWPeQgYPf9h1EFRAX59EFrjvHUZji/akjFrYrxd
z67VEgMOvBCrNxKssddp/WccpGAfiCPMilf35x4D1JN9pd5DEEwAHBI4WUgLDtZE+2PkGf8irsU8
o5rzsRvU0FHA6X4wEiDtDNbaxh1ZLVpu/3fVaioxGYa+Fr8ZPQN/CqnW7x9slzYofBleSAjECEtO
w/MzYKc/UGtLa2KA6eVTikBmphjKb4i39PEvFxpbd6FzmfJ/zNyauSq7t0zCn1On+4q4VaFAwoT/
OfGhwrsFaVU9IeIQ72PjqoByWh2o8kbSItFoTMH1l8GGSEQtr4BTJw/x6Xxbpuq5GGb/CdMDWW00
EUyXyvfls1A7L+9LMFd9oVkyzBz2b9QqnzPIB/qg2ZRIuAqn8FPWWm9RIXyxo8tje1oQImyufkRU
GO4g78PhCMN+JRQTOHo2NjDMNYfdMhMKigcTnHZp54Y051OnyiLdeFZmjmnua3UA4yHdi8AgAlIK
iHduxPLbq03sIOczYhMKrfBmoiGnftpKK8byR1CILSNorIZnvxFi7brwcELI7Xj9/2fJ7/iFiysD
hVc8nOsdFRpLJPrEwLl7/kyMVJa90/vCfLLoztnBNgJ0VdsUrQzxB18fWeja8qKzgp/rjpx+5++b
pLicrvUBpgw/QNp3SZKXoxIBSM/W/SKXj9uprh4+75nn3TlmnIs5kLs74gIe/HC5gIvmE22RYRVc
7CBqIaEPu/uvfwJ1TAmVale1HdQ0RQgPA4Q8Ez4N8ZtSeRS3Q18/kzbgg/jzqJlWrJkEpbnEhIag
57WQzI31GdEbop6CGXGodQOLoUMuuwMmY9rtfVyZRZYYoJhBp0WPdiPEY3fQn617oiZkyu56qOFd
FT3ma5L5pAEVhao1GBi7r26zlci2d9fLZElfYtBHH4FICD445zRcYTbMA9r89BqogtsfJtAbCCqt
cTkm6dpRFQ4m5l3bKohOXy9RGbquJYmtMLLXKup+z/plfcvUwcA6hELVLujIQYUvvAS87SIYpdoI
XyMnK/bU5zuEyn+IRwGGmjyXl/95OBPk2UqkpEstvB/WrQyVSNi1+oL5DBQDbMwcYCW0MSrfz7X2
BhxsBSaFqiCl4F2W5SLRupvPmD4rjSjHyyNQBvQdp0zaxnfcQ3FBzjb9xp/8+ud7G0khz21JHPNX
Qs1r1UeASLONx1JVu8L+0w8KU92ipVsZEHelf3QLsyJDBBw/ri8/c0hzh5Gv5VIl8w4irYpVJ7AO
aetgQHSrjWA4KqlanBDWo+MfJyR5t84oOKJB5kPck//Rq4Vq/kLqRbfLOK7KAXB5Om/vEE4cZy6V
d/CryK+EGWYG9fYDWsOdcy+YJzLwWzw1bSHVBewh+F53Byij5O8WcnwwBkLxssVJF1Yn1B2iL8bM
a4XVCpFiYKqGlbVNLPyFCatd/F5Ba+ueHW4tL6L9eU79W1gN6MVlag0oz9barplS0st+Smf1fSAO
5gsvIip1jDF6UP+uvhCAIKJJiWhtNfzBkQVUGfcuZiQ/R3sQY60ZM2ID+C7g73M7lLM0RHBX3Oht
38QhILtC71kv8MD5MFWVVnLesHDh1ODk493piNNukFsY2NgUxI9mnpEiF6+hyrHBu6vDdqtadIu2
6n0dFEHOg2tTYPVxbgr4D39vj0Xv3vca6ajT5IcCw/ES1vG6VOZb6YjBLgEyZov/eNL90YGnjGp+
yVaF7UG0new3kKJZ4JNzTdJ0+ggkAToXEKLuikkGNaA9PkBtPLqqsAjCxvvLAyPLwWvw9N88Q1Kz
o1kY0NQIvFqgwO78U74uATw+pkLcqqG9UE0HgrBRmhBJ0+OANS+9YmBEOKdF6/IkjwfFHEfHk3Q/
ZWvgnlIvyU0QXGO/KSJywGSyDLAHkARf19ENERs9OkHkPzQJ1J5ewrfd7BpRHrhiH1Z3FPZF1byp
vLMcquIASAEx3HzB4MDrFTVChYTsBL/X5AvgGdrH0s3qfqdupgVd6NrWrqe6fFXmCLSeqD4oLbv3
ndb+oEgk1xqMbUpvlD3N7lwWuSJc2Lt3Nyu29ummysUx3W/Awbujub5VXTOwFmT7lpcFgOobz4+X
3jrFxdZJMhG4+821xPg8y3lNl4ENMkG8+DAejjRCixSNsOVTb52q1VSDHOy24Vm4i0TLXAk3Z8ht
n5WTUooX+wsP9/uUfns4wNhPfHf74Cgzo2NcFVbqFpFDYFqgPjN+/1PJIJPVADQn446lMvAlC707
LDQMYNfb7ExeITJ/MVKfzPVziFhR6L9qOK55c8XcNP8AVkqHLDH4BzgKQgvPCaHB8C3ZfexyXfIo
YCf1YTDaQTw8o469a54OP+fdDZsAAyUcg2j06pCaOh1XNcmFwe6tfGYmZRPuaRjtjFh5zerv2JNW
TB++S46YpMbEnezGFIALJhWZEqPrWjtM17306H0N/JDpAhRfvr7A7UOkNbZEGskME5gNtQuWwK+N
0OIZ/1JZU1+teBsL33S7nZQeoq4l2z6D+fnv2nHuFv8aj8nJU+SDGtu6VAqQts7IlkEtdIqLdrIk
LIoAd88KHFJY+EmNjX5xrKPXRogeN54GrlGxDHEbHs4/FdrvUSZ+CTNZTZjUlBrCmtdbv+e+2neX
kEksl5ep71Nake3uooe6W94rBWr869fnDJMXN0r7pgukpkTlWlRzm4eROppJvaPwLNSt+fcF76nM
RiJQtvO0kIhdi51CuSa7pOMi+ODaUyFSvYyXTA6zRS3kNn8GzUw5Slvr87ESwFqotVuk10mRu3LH
05W5WD9eAxMMMiMOTvPPqR0Fw47fCEU+qsKdSYB47/ktCwPcwzBDzF1f7Y+7WCjP4uhvesBitRw+
V8UPP4WngvdZGSDGml6n82VBbpunOnUZOJtX3jlYrIeLP5mwk9Q0h6UN6zxvZkOlmYxj0xc6XOkU
xEBI4oW8SWIUF22+gwhjT/FKanotxCLbLOekhgBBxY3M/AKpDvhQoLK8Tj/mRdsLMrO8LdeHKKOU
fRlQGqxGlNHdvjuN44jxchjHhQ6eRJJBBM8zO/GXaM0LaPexrpLaX3PCdhNbR3j2f7CpneU5AiIW
Eq82rpUKjZ17OwYgKcG8mTzttUlq/THDnDeVcY3Nvg0ape8kOp8nuLvHYt0XNZvCrfo1Glt5Fawd
LPKr7wx+3dAhGI1rR8CJ4qU50beM5CntrQYzFi42/o7mp9D4gQNlFxtrxjpSLzYjIH+0FrkN1p9a
Y1FY3Xd/DxqIpT1EnWa0tc+NSzuWdFvbl9FElqTysStuNOYFGllGUC8l/G4H21WHFIz9x5YqqOv1
eFgJS8i1oBNH4SubI6fdeKj5K2CEMZ2UC+wgQD2O2kv3hlKx9L5YJxDWyH9MGw3j2Fl+XnyJn0kV
g8Opa5mx4qVZz254SnFfJF2K7jWdcy020SO2nZX2SF9DSY2IztgNhBZsRLIvrVT+QIqUtWpmCezS
Oid6m8pOZb7lFmWK5hEk95tG50ixJ80iqJLl0T2FCDtKTnHFyOyTWDYJb5YovucFPGz/+MrjUWfM
+zHoa9ZjfI9YecW3mTbb4DDlwoVQK0h6OxGrzyEKX9cHndqdj+6EFE5RKK5rGGV98J7tjK2H46Ft
cuSG106+R8vVwTposS6KFnKpLHsrwI9wzls1eHsCaCo2BN9fZZzAudioLsSSj4H8H5ozyoyhHR3L
LdMHa8kQ99Jhwq/5I5cbwo9Q44WgBhiAA7YGznek5BJvwM07q0yYRHH6210jsGNsaFOVgxWX7ZK/
rrt5Z9qV7GgoFCnMQyQ8rfNbfFRqWavQu3S8ACppozrMP8Y40NR8O6luBntXQjGz/DTdfdLOPtLw
yWYtGsBNfis3FVcQSK+hp8AB/z5xWbcbE6ri++g2eL4O/e372H8JD4jQnrOvGlaQwrbKVvOw5Hu7
9a+0x9EKjLNx+0DQEi9iGfV6bFUxzOybbzNxIv8WDU9QFTu845YhoOsMkWFk+tN05YMfb1b+yY5R
nU8dlDUGPOjMgSlF4ynfOVwfBX9pnkbaDJP7X1Uujqoek1OfgVBRYWJtKfl3GDLSV0EdYnvh7Wok
e/Rw1MYpEUA+awG6Rhp+omgvmDtBO+Syl7AF/hX5mX2ZebIqju9/txtqxvLMxKj99Cv6q/XvpQr7
mt6KEnE3M1drR1m2wE15y9sPt4owGT7AaM2tH0fbGKMc41fKWeRTXuXnqjJY+BKdSUCR6prrvZmH
WWudHaCA/G9bI3X596QVv7LkDQACqgW3JBL6Ua/qhu8ix6iLJBTMUl2UDQEA560z+BHRmtDswC+t
QoZ9F4D5zIv6zbb/LCoTi3kntPHoOrEmWkef75kZt5dNV6YXRj9d6aDBzgf/IV2q0lbuHoG9Q8yd
0NfwyhS58v/vxmQsAvC/poiakF3+wD6D5J49fuP8yEct7efsjlNXYTKvS9yqlHVJKWKkxVVxxO/W
lzMsljZWeusygP9dM4VnNtOUJ65U9+0q8imgglzgDZzr/jGZps4JfXgNdDNIGJG+8alg1Ohz1K5P
4HnN29OqaHXz1Iocs7jI/F7B9zSuOt+wfwAEZbLnsEb6mef24Gs4U14U3HgI4iSgtRusOKiTcbb+
AWp6IfwsJ362AxwJtNWhQGPpBxFvoENqGOfbmfwNY2kBZYNDt4CUXoI/PAa0UzgniSZfgSEh8E17
JbIvckY3OS8WH3yDihO204EEXgoa3XUdgek3VcM7BQ7b+qt8qAw2hvvZGFhdg5DCd3H3QavNpkNR
l89m5xCrG8LXhy1a2Ow2ss/SoP6Oj2IGuisvkEj4hQl/2ySDZwBUbDWam3PjobP7IIGMCLA+Wx87
tdRiIk4WpVxVzzAFnt54ggpnQsQc9gxK7GXl88RAe8CQ34y0AXH/0JVjLmmsrQ9HB+V6AJuN3Apc
AThISXLuV3wMwvIBjIEFEguVPnyhBcmcPDkf5Ci9rtJTON1jMxZSkWszARgJeu8NX6Onq8hBoTmT
tJH/dkm+emnfriunQIqGri/VSwrlXErYcdXsOgPNP8NyCntS1D5JwBwFGbYpJQTJma83UkGp6Vx0
eac0rCspBMqHMxLNE/5ovZ4uApWx+Dem8JHnYUMUbmEquzIRaavM/iTQlh8WKrZI0EqHH7f2zf8A
N47+MwC13Ku8Zq6l5coniR9bcrrqgC6CWlZDLUIjc1cWdx7JI4YDCl9az1Bf5OLLT7ULaoddRp57
8vHZQc/yNxAyKBvLV+lWZV8FVGKdBewGPU2dsX7/eHU6D1sDhMIWtTn1X2f9od+ACfq8ycNNuo0a
5uGTZ/X3t0/qrfe7UoYzcq4WgAhYhZjyUzKUEhVgookKKq1Nr7hk+gE/1SOlJVRwKs6u9WqJrA1e
Gd71g3+Tq6Ths3JsDPhR9WMhhIi+yVBQJa56+OYfpjH4n58ManYGas3GWofZpupSijgpqtVytp4n
zhy3C5DwdkJa6MuvF6oOAJgltQCdPYNybYE6HF+Tj213zyGBGk+ft/H+xp5iuhNVLvW1rN3Xhi3C
RFI8BSMwZo4crKD98jPYMe6ta6XxwL8k49H8WVrNyADaMT87mDIiL+kTFo9fU7X7wB91RVQXs+wA
lul/K7tV+80A3w0rBuiWGSpVwZlIjrhZLA5emUUezV1Q07NvHf3s7m5kn6ZUGb3b3sd6HTVtoxkP
COnWey5AluAd4MdI/W+qNR1GyhT2QYLn95X+WD1FnLzdagEyGnX4riuO9//TGrdVOzH6jR4zHmol
0pQMjTeDcO4eBKMYA4u+SZ4QzRWgOzNE63P99C01lVyx8jpUN6WN+SsnY6bxTZLrHvN2kHfY3qr+
xWyeVv/n6pbLFJdIiApRHJzICI/s26CeroNgVTle6sgRNEu6EyLKH+52E99tFcudW6DfZXRZY2Fa
kkF/m2SojHNuE/l9mKUfyay3clA38IDdsfsaj4dKcceHdyUyxmJBOYfEDqXcDg9tcvmBHBkMl8mN
XCwfEMHCPGxtZIfysdg1xmj1JVb+/M/VSm5+kg4WtJkIrwvWowdj2tcEwCppkRXIj70hrn+odyzo
tD4p8fYcXp8Jn7JeMouBGQ4rw5TGf1PHOEy1DhvMc1BMPmOhhuI4QEF4dDXSm9Vf+oxzvZfgnC8j
dyX9+lruPLqNqd30yPXxXX7raC8JT6MZ9WOhHtHCin2IQ9Mhb3C3aBoJw6d9i8MSKpFjVxHVSbye
PALzo5QTWqq7DBfP8BoXLo2RqDxeiNWKMPM41vYwFC4eDy7I6tQ23Hw4vKOTVTuTvr0ktHPN6OLm
3lL2dDYMdhQ4nLwMwmKHexShhdzVdEDJMPFes59Q17FMhqACQCu2Iju02kMIqvITACQMX8KuUOWW
Bw/DkkyF7rROS66ooR7kxZgCV/VjZ2UCuxF/JzCK/Ym8XGYxDB4kJWVryGGpj903yAhp8OwobHOP
WojCkOVME+wfUt+yvbSVGJ2NlFLrs/qe/zTy+qhgsJ+Z/bWj1c78wYqtGmSYkK9cVbRLF5oWdix+
F1Mli4+PFhFaTcibL1aHdKr5adzptKkienV/B83jhLUZiuns/RqZpGgJ2UPKe+K1xcqkmJnWESF3
dcXDL8tDsA1y7rcFVztxtHVYGwRvtdGuH5W9wDfj6x/PoH8zbEZT0RlmqFK8pyGv4NlfG8kxEa/i
I9alVMe2ljBSKpuAKRlZaFODmjFUWqCPFBNXiLJrGw9CjpHA25wafT30LgNTqu96QFsjDK4FWQYT
y2SklMmuNQRPfaylzJCF+K7sx4jDB4HL7lTAxI/iv3LTLABACXznVUaVKhGd83gKlbhNLu55PJfq
zxy/L2jQYVpyO3sSBBbRkfJ5hk55FH6owcIaEmH+RRC3x8MI3SKEfZtKG0mZ3WPULNVnnqZF8Al7
LA81byp3fFpzCl0oWd8Ki7qTwoHz/xUsKzRX7CUhajWXqIUsb0lgGoOBeoqGUSdIhPXcuddrs7Pa
fEcY5l5YM+kbGzB80LaiEEMude8aUn8hYK8AyjTGXTkE0Rnn+VI5NyVreZES9wtJZvcyvI+iJLc7
R5bGniF2/m9Mxsb54JMqeploF7WO/JQ7VzePY3pDxbmGK/c/tkRQD45RVvQdXQlzng/1rJ/Sls6p
np16sTLxMTqgOBGT9MxhNyLfjNvdj/sI35ejNvTQPa3p49DPE3GJmII9vi49RD+n6pOcvo+k+teo
SOUFafspqKs7oi23ydCmMRulwlye7ciaF2q9gBEaVyPEl+t5alJx2oemE+UFRmXPmGAENe5tLUZs
lLa+8se0mTueywvlTgamCeIuzzB5aH6g9QbsZoAvTDP/DnzCNbTw2+ptYXnQS3aIfrbW/Ef5DBTL
aqOuj+34BP0T3VO+TDhBMfCFlXhZ5fzKc6jrTsx61dS3UYK5/3xD2FGn9wQYsu7rUTgiPVIm0VWy
tRNniOhP/D/c2Zdm35MzB6ZQQJz52FQktHEqi/hztN9RyPf2PTXAm68Hsg3JrUObS0CZgZbgBtxf
qxqB+tNv9yI6c2PskGPQiJpgD7SrPPxLB4fUMaSxqk1GFcQYVayznAaZdW1432SyFJTi55ri8xTU
UIqQFbvfTRranD3tHSe3LxvbIjK8NNmG+cBJ7Yl2BAccWcqmRaj/9fE7YDCnJliDrCRwqptzAMMS
dOPjzvJxyLj4+g6pshD1lIAehji5yXCoNGFNpFKsM0+NRdHcArr0o/Bgg0XePQxZFQEAuZCvGH0e
V3w7Ed5vknXCO9bJYNY/TzFLBLZNM8dAKzNtCqsuVaLPMqe+PTxB9hJXtNzOWxM4JqOMOkQCMLin
380RfR+mQLpFVTq2+BzH6hS105pIIbdIjQcvDFJq3dM/j2sCE7u0CACAyQ4vbhmPinAQWIJyhnkB
MILDFWaXKwKJSFy17q5BOGlB+xXG29ZuwHPDC8nyfBcE5orQSNfpQX1pkbnztw+XHYJ7eMuG1owc
2OkWPr23jqGpXMKT0E5tF1XqF4mAo31Gt/Lg8SoEu0bEqP+eZsD5IQMXXyoPnpujafm9XmGv8CGS
bTWdN9nfW6TWD8xzeM+owRhkn3FY+HQWj7Dixgc9e/n6FJESPhzvMvZpzEUTbWCcNTpao+cGi/eU
BJ4viLwKOJLwL+WNVAVwSTfSbnNJpxHzfAs0fMlexyj1xtPFIS8vWqu57tknMqBcSS3sbfe9Y3tR
YcBwm3VsL+cgNNP6G5kPUCa1HcXijY3VAi/XlwZZljbI4kvW6jYmLRLjOO1co95hxdrQY5iYBREW
BCRd7mAaL3H5Bm/TM+rbatrIzID5mvNA250dfWHejMctAggURo6ADycrQk87fZ6xh0if5oHBhe4s
+FS8P430CSzTeNgYx9DMYwKPAB3CeyBX6SjhWICgRGn3j1CdoSTbRpaxtGeOL6u1zCeX3f48tc0i
L/t7LYAs3SKDsyAcR6XCXIMVqXWvTISFVJZhks7G7VNq5HaDL84WS5pwOjwrOqt9FgFpwk1OdNQu
SQaICpGMKwNmpqpgwHRClCTa9i+8vPCpNCm7yyiAZuKbrvVKseaFzIWIrp9AESV351ZyuVGh6/Ex
63Lp75DIfcswcH67XxYeZe3LsRZNgoI1DQ/FuzE0xjiscYZLBg9VuxUfxmx2UcfXx9Tf0132u69q
QAXcpeFM8VbiUBXcePKH09ChQBODWe6sqQtJLJWNujowGaoS1UsB3lA57GRjnaNATYdf67kU/2jp
pXMv0RLrEnNx5FmU/VMqWFRkhX2W3iM5R74Bdu7amfjv1XwevaMquM2eHjkMrr00kGQPpJOctaHi
Wlk+iYwd//LybRXpoW642AOFASWIPSxHimUiUy9bF7ITbrM8UHlLHXzA9RKzoeDkXPv8F+OmOe3H
ZSpzGDY7QnfHFtRmrH8qQ4gPeHViHHAjazhQWrGizVQ4drVAux/S3z7WDL+eSNLRd9vdk4Ctym/u
5zJrJVpUw1Uh4+/QWgVRpYqdjaMMWqLkp89bCVqGgsLNFpJ5qo08RFA6s0IwpEZYnXSqxOHQvsc4
mWRmsPIaCT2C2MlwSx8bNSmnPDO0wabJhESxPH4EW8tEj7TFSAwg5+ktoj9adgwZH5aHOd9618Dh
nJKMNzvR7XCH88XTqZEIJ7PsBO86xRFY/jseheG7zRcdI4hWXaVSxiuimx4znbUlduFm123KkUNy
BOGT7hIxSus21xOdhRA/f6Trl+i1sEPlC51PvPETdrcyEQhEC4DDcmcSPzOjo1GVu8RxN7u2YRDv
BneMDedlLhXPqfedJJjYJg4wa6PNRSKDufFVDRDhgv08gsS44WvfpW+K/vhfMHOsOH/dGLpx4CmK
5TiBWvx4jiByc022Ih5uBYFLJC3/5F+U+bEJY3wAsPXtNINAjI59yz3OqfMr1jz1CfS/ireie3uZ
LDosNaQfoXVMdlRbTImcfFBJKoPv3v2Rt+0vZJnEFWt3r+ohWJL7Wc8CV3+qdoUBgSsy/jIlRqY/
nFe8x24hRVr9zbmilEiv20BkoLDYogm+lnbOMtlnWmbxs3EqWHg03uKUXw5TGKA2FdJXUT32boNP
aNcY2KHnERNPpY/typ07o6HsFZYSAsUAc40IC9HR1lrnIgoS6VrmdXEM3IJGjEjwS/Fp35xrKr98
iV/yT3QLR4c1VDdTyRLo7G2uliPLGnqTezlgsTQx2uK1TXDsUpWgCvQfLW6fLMJR9HjKoKvOGabQ
nUo12ci3oCiTi8Orm4VgoydRi2WvC0GE8R0+c0TnG/QU7VN3hXHCoGYom6bs0KWVha0oAl++KY+1
VUkbhDrnmgcGxtoDDS6zOUbZ/g8g0xPLD1i1bTppdrmcSvbXSk6D6icfPFphzxRTodEmH0Zu09qD
EGfnYSIWmcijN7fM5wJG0xSEZfVhERmhB3TTQCnLikHdSUJ8j9YxDgwshtnhKgu4WPBQGIY8KHUS
n/8xcbVeLubSE+CKkg9q8ySzgVgxt8Z1GMszN903lSqGRMw12p2E+o04GfDEhbyz9BHhmPdQFsXP
qxZsNhb4waKviI6DITj/VCzzNO+ZD4o8NSd7a2gsjckHGJWpKRYtk8d5MzXT6Ahhb6TFs03FSO6N
oYIpYOI9YY9anNFL4AbzPRZLf7fHHxLFTuwLsnhHniEr1bjcK1Vlb7K2qezjSPf5851qNzbQ/ZtK
ogop6gXWJNbeejbkLfLKfVVeX8lM3eTugNRqNEDSwMihIktFQ0OagGkFlPl9Ztys8d5rzlEg0UWe
GcPPK9KnfxMugTu4/mtvvwMSYXt5wgSywDx3JZZgKsiQRzSMcauSj0YJotkyqUxYTSijUFACbW9K
KwUKX39uXeWUC2tJVkAwbUhxbv7p80A1/37C21p/Pg+evSnJTcvyGpUvInolEAg4V2fKuKtTSxJu
quM6hsZJUESEPVsqyL1qyiPZ+1y+fu4WK3d3N/Sj0QylSu/zyzSQ9IAGZJjH+jrZ7T/2hnuXaZ4S
/blxLapKvRcrGWXflDQTscrZ70rJ+/bBAp6AzU1vyRBhlyYjF1jWzPkjwRuSzzb9RHt4GRmEmtSH
YgCAcibJ09ssXDps4Uh+5rpa8Qh4p3nlQG5g86fmR7mUACoXJ33ErqvX6w35nWydgEh6Ld6ZPvRT
vIm0Z0TuQGlbxxhAPNufMQQmitsvYtcGcTukhZKjDB+Fo+WwDG4WK6JTffA65dEE33XurWlCp/i7
bV2ux/jW2qLBnZM8wnnmfs4TSfB4DRl/I1mO0PEpUdtZ94Qq4ypA3z8tuePZzPFYh1d3GvsttJ3X
EdSoYZCdidQuLbsjhQ1s4rfRAIdu2UrThXDkdU6LaNpHJhBceiAyeRCK3SbiNY2Qb87yYilLOCy9
KcQzvF7Fye3HZHMh/MoNGNy6C8WnN8AFWmN/F++aoLVkqw1Vhoo3x/OSaQ27Ns7a/uHnlvUP/ONy
3TPcQAPNMy4UoCVlg1Sz1nat1ECg145d0diHG32tvLBEBJPM65An6acU9GscuNMkxCKgwc174mJF
iAaXb65PHNduLw1HhfACRh01PH9DhbeuuzcVupRWANl6eMRyYgJkLnWk8R2Q46wBxiX6tLTWnWgu
2elZNY9lnhraWZqfG9yWtRcFECSz8eVnW9Xot7Pp9yocn3/6+i40e/YMOOGePN41Rh3UXh/QPakK
YTyjLwiD7/QqrxKkc0VqhX5r5IKNxkAyHNl61hXUZmAGFfR1qEkCaiigwpo8MXn2GGycdZmRekwz
4VRhR4YxWkfgGKmA1Kp2MWqWOPca/t+nxaKNSGGGBXUGoK2MC5er8tvSXwbPEk/Bfaf/lof4n8HW
eeEsqKueB8cHyxC5Rq2j/JC3BMtWaiaLkgrGu7Vlsj9ZIjRGIEiRk6EvziT8HU6gz6EZdBBD28hN
cPOXSKAuopk/yVsxivFL0sSkU10GQScW7TAtPbJnpmVAoWjeE4VsjD7IVPbtXnP7YSTpIHBx6MSL
xClLGyxys5HRT/+ytYupanxJYaUn8FLEpRDk7yOkAejhWTLzBWPQW2demR4/ftAHWJPFJRqDU9vF
8Mp10fbNAD2WV1VkCs11rsDEWpQvLIBBugQWP/u7cljR6LpgmxysLni5CP3aldQk50jZ8/dgSgrG
gQSl99fO/AhxBi/LufE+ffUeQjvbPlcivF6xvgBhan8mzYvCEwQFztaRScl3GgnhQo8QNGgWaNW1
V9pN59dfqe006cNAloQVYfNNlRTL3Kfq4S5Ki4A70VzZ02JZ+sKR7zt5ELhbRWfb0lDo6fjxTirv
a9LVU0cQFqrHDYAOoki3m4JjXtsoVDJPPlcfhV/RmxviY7AtfwVXHDR3k9dNhLuE2v/jp24KE4+f
UgTkmSFd/V2u+QVqdNxoRI7diUSihz/cJujHddJsmnlDoEfmGVnpX9LyrJK9ee2cScYIp0/RRNxl
IxzvFmdMGDjKaxV5oGQG7Y3VpI9+OOgEKuWLaCTP5bn0g4D4P6TiA67QWQpUxCICGQdHGoOVEv7w
BY86v1DEOUO3PKzvgHTYV3G/jUuy/MDLScI9WfFHLVqrBTTEWo1JjjnaB9p7dTRoSc6um9CM5F4l
JeDsqAoWUBK1uUQ6ELKQmmACo4a2lO8VP8jlaWQGMhaLt3KjaPSYEUIjdBc9nIqm40pGDkqpSLkM
LGvNuraTvMqyBQzewirvFTbIWanWsxTgTUiDV5UdalYCZUMDExibwxA3HDugcH8698Xm3Az7Zna5
oOBWj0Uymlwq6Wq5H59fH6/FM+5m6s7N+RD9h9TCTWsuHdCg4AMYWUpUzF1J0eEa2EdQn/eWd/ji
FWuSIgsvI1brb9ho6ItWuyqs84ZDzgvupr6chMn1Ajwb2N1bST15TbxUo+GTzPV8GM9gcPEfrrJ3
41jdz5ruTCXWMyGy+CwsMfAUrNw6qT8pTtH+Quy2gYzD5bRS8XLyNrpeOmCX4bvuY4jNXnPL8h0y
lheU3d6KaBpqXYjWI6O0AY36fN69jKk3Azv10FNDK9e2QEe3hCEAmTMeHobniWKNCF4Wl0QX3dpT
DpzlAofGhkcVlSdWSBB77S1eSvQknXPR/afK4A/aOdqWfbqKvnnvIInklWOBGb33HpbPcHM33e4X
NBBeZs3VlUtxhIxZOezaskwggeFkOf0rwIQ3SfZlSZbrZvVrUMkDidzD/G9H81U3T4fYKCcOV3+S
Jx+dYzwB+QaUO1jh3oho7kQiNrMF/HKqo+ErQHszBKqp6ovzMeFopH4rXt66Ui6MtCVbo1wkI5yI
TI5e+yqZETHUFBZh/Zcl3PeAGV65hCmnU084NQNGDGrhFqwgw+CUuWmNEZzq7rUYW26CQkrM4+94
6meJ3aWW+5iqgKNPHqrc1P+O7cT2olXj0j2FDtcuQ0B+qbp7Q1PNfri5lewBgUf8hAogiH7TEnJ8
fi1I4DthUbkGetZUNZ2c1jYcBZpjRF13mjTVw9JV4l1XY9Nsr49d1+9jLRx9IKwjVsOEEsDllmMw
7w2wVV6odBAiuE66C8GGLciiOp2g0OGuphUlAzMlnORjSJl8kUQ+mS0AydtOwp7ssxilXrbuTzIM
Wxm5S/b1l/xt2IpY02aiiXShjroAvMY72LREuZoqP1O/aiEc+bxXy3vhsHs2ktgvYAr0pW3PSAm8
2+KGnC2+5SYw0gFaFcT3HTLEYLFBh2/a6QLII8LNaCJLXmDFRheOIw1/DXS50bB5dVGtU7Ahz5Hf
L9ya8jfce3M6S1kbUc+U3N5+AGtNM5ObTO0nj3MjMxKMjBqay7fjMYseXZVh3AyfRVvCffwepK/g
YhyMtIpWy5+S/FZSV5f9M0aLU4q7GQuL1cehtwWDilIgxoeJGSRyvNGpVQS491J+pMfGFbrM5yS/
CM3Cr4KsuksM6hg4RPnXOmbzwEAABDTNmpPmL91sGvOWEoxnb5dXhLW54FCzAieq+9WO8WB0I+Xn
o3WghnwAlJdqqq0MTb+e+f5w+L+8z2zKoLzB6K89dxWL6ZoIZxkIYDBQEByQqcN+CCWLmYxoKz5X
zHUpsw4OETt0xJdK+g9ezPz85qjD1WDMh333piKinvgqqQWmBk/D+JSD0rWQhXauNVBLXvZUDYhh
UXpma+j0ic0yg+KJ0Dk4Dxre9POC3b45y/4zXOC8WcowpDVSks7xNFF6fBHahcJK5enXrwqXp00R
ldL5Ym8a2WBTP//C0LBa9E1jBLSDjcuH5E4CS38MWvbKLC5awekpEbyowwmlRATr3mPSgcq4nnBK
x7GnyLx1ly1x72tQn+DW0AL3caPT+ZUzUZ7ZOyjH3eB5d4ejwdnQxy8sVfWW/zmuRuOVdC9+uVeZ
kMAOT/0iesMKhDq88HZvJsASM3dQbfb8L5nZwsffnTkCVKedmZzuqpftHHFAD8xaSVMmnRvqoOfP
Pi0XR6N8fFr2KPp4UTUtAMZhmj7357aUhLel1dcqqvd4AsD4VVxx3fJEZc882N7zT8BMbqjGoaR3
VukeYSoT27sCF15ZzVEyywVVr/DgkGqBRmpVYIQm9XEH6Rua1ngSsA+PJT37vf7bhwWhNvnfHVr1
weueax+4eDwG8BIJXxZ2u68XpEXpTLAkvpS75xLz3MVDFqAB6r/2ZOSv3N92IhI00LbQxMgeTEQl
3+bAZqE8/P37A5U+x4NahPu2hlLC5qef7h3JNzvsVDapbbNmgg8/8nVLcFmE2kObM7m1e3jUu7Kw
Iw7LYIhdOCE2Bb9wRT1OJ86kDfYyehc4Ochc04cK8PAj/SszZpiHMni9Y1fjtGp5glkw/5yEJIQx
tnGyUOnZzvFzRunZCqqZRjRJyOAD40R2w0CeF/ngLR4Kw87+owNz23YzxjEt1XMLT6baGVOskCIt
+r3wps94n46I5VFq6d8pUwqw60U7w4V/dXo8RkyW4+h/tQIUdIC38VC6CteF9WOR8qWRWIBDsFkm
LZkFM6RKphwonPmSk1S3FzgYYzuLg7qifLPmboRO5c5oC9NDWcPPpPagwP8WY+QlBN7qSnH/Dgu0
CgfWGljXrNP3yLq8+wp6ZLIk+i8ubBIgTiRBEOrvcKmz7r9h1ZnrX3YE0noTniuhB2DPPjJT9nGE
M0sr53XS3imva0jPNFHn6ked/FBCEFqvC+tGnizZKp6btn1S2ciYmFk0oeKDLMx40UG15vg/QLG1
AqMDQjeCMy7TNYoPeybkgYbAaH2P9DpKnN2F9cFWJn970HwKT+3WpIISVrrXGFUGcRWpN5LtEP96
RZGI3lcefCl+M95Rm+Tybuc+XC1naXrYqx87FaesWYTO2R3dI+tuYwwE0OUiQj8O3SFSI9RqIM69
i6oqDtU1ErcexZfDf2aogmOBxjQqJy2SCpuBHqEDkrTPRX8PIY759Xu24JCUGoAPs6uP+tC2WVWJ
kbdF3tNTMZ22HImi3QQL+zk+Pqo3NRrXpD4zpsj9LhLxU6rVROqU8HUsOxZvlYc27NOLUJXHJRHr
o412orytPhtbXc1gMOZiqabAWfvkj07es01IsX8lzGUyEUM6ZcWaBPaTpGMsAOs4D9zThYzBKiul
Jub1ThFwRk+idvbYvRs31ASvQH3BMez6FvdxkErAy28lI5MCJRVarbBsnP1tc8l3AbOKyDK0Pb+U
E/O/tdKkNBkfkfYs4/b02Z2lNgafWUqo8Q3PhoqqPQDzx3L7n7Th3FLW3AkwgPhU04SruIKzQbZI
RCYEp26PRLRisuiYVRrkamdc9x7FtWcyzf/dBAsXzjwQci50iuqYs6m44w4xFdDB1lkuJPMHw0nE
lDM4oV4L+wGonfwNHv1I+DnHRCd6H0ss8FpilG+ObYvIE7YbCzdHWFeTIeTEaFhokhr0EpLG2hbO
NxKz4CEF3MMaO0VH7EOTUvspyvmDQzolhyRU3drBvQMcWJajsMsKvtd7vPJ0AH9+GPLvVA90zwh2
lTim1h6VtG/zF+xkuVwRyx0s9hRH+oDB2CaQNtAQKZRAdWOz4mD7c+5d/SnWCHnv8uN9R5CScRCV
UF1SGpIaCspADL7g2auniRdLeyLKg/E7L6abM2JpbSZTgbhHVmSHDQmsFoHJo1pwAVHG36qAO8Ga
51tHktr9IiHty34+Ogp/8DMYFpiqYiQiEH5VXpL9R8YaXFtG6i5xcHY5Wxyiz0+IOGA76bg8HpNz
qLMCTdBi0YqsCPDtRCr4NktEntEb+9/iEqP2ZCPpj5stvpDrxzBLRnc1NQZNHJkm/MsayYDSdreV
Rgnrfq7/CPUqeKRHCeLuvbr2ypQgQTb2K/8TbbpJ86pgVKI9p4CyPOHFqk00JegZHM65rsEkLdx0
P+sKdIKNT5rbUNtXiQQwksDFIjW0eLzHaAOvb42cxRpcEGFZvj5R1ToC0/7MmvSOPo9QLrChi77g
rkF0exkZdvJseD9Cfb5Pjd+0Aqkvmm0+7MOg10hcDpXdvb2GK2OjqrHyz/gPJX1SrYhvYxqK8tty
BDymEDUy/vNLLE4S5NapmUjLkhHz8VWgt7SDLnAW1AYDg8CsXA85+GyCJlyw/1ruDsLn3EtWBZaK
qom5vVjKA8hBzzNyIOE7a4eaFfriMMaQXaOWlRIO0bHjDqgFQ6bDIo4PUL9aI00CKH/KTyYekuTc
KXHw8TNt5xn/RGtT7ZcmxSki4/C2YYvERn6iESYQV1TnTTr/Nxmv14tioDCSMY6kQVkdPJkbeQMK
enTylugqvc9+B5Y8uBeafM/ZxkaPr7OM/yNvyc8f6Kd8inlQvxkm8JGQz/v2nn4ibJ9tqYI3XJC6
c0ZLKjMUBg4V8D81+OsSPKrb1/IrG4LOHJTi9uM9rePZ2U3V4B818pM8RJ7BCBIOgk3YYqBYDAbJ
pyZBe6axKy9Rz7Wh7AAqn9vscL+Z77lZv4memPULRI30JOjpjKUaeYxmE/azCESeGQsQiDxYHtqs
P1CI43eXaLtFlSSXdHOYVApfa0Fbr/6R5YOPThO5Y5+HL33dnOBNpVzpuyrfADU7ou3xo+wAy0tP
sVaMjVJYPVxpPsI9VaxzlNcbejWQKU/+8v9PjMYJZYs4p0Q9bw7CFjMWKalg2Z3MwvOB+9oWwIqZ
P5TPDvJsPsa3EHAw16XNc91BW2T5GJf1pAPaLlhO2lYFNt6S2J9jgdzTFDwt3i11SClkBffOAqJK
4K0lmoVu2QUC+ildll3/OgjcG/ZIL1Kruc/sM0Dtx2izV4Tq/z4Q9G4+zUcJK4xMGkd1oxId3Y6l
Gcl+Ru/6VMWioXHjDkkibDfmLDAEPUOjwqMtIsf6Q0h0JoaDGXEq4qYX7Y6DqacMceNtueNAuaRj
UqkXH1mIXET9COoAJLh7KVst6KR2TABE9aGV8awFrFIVJksYWO57K5GXqCZSht5t7ygECMxdDdeF
RjYVHVB9hRgC+t9BpdTcun4Dzj/UGjGpCLsxIUdGP5Z6YWEUSH6TnswRS0h9YUMejpXMsoqmng9S
as3L4Yc5wotm7oQfYMyZKcuzgMI+sswPORKy/w/Oorq4s2iLt5ER1wQX4qKmXDPTz8SO7B9mjmW/
4cKXzsWQsGIfo1ILhaKqk6vPl+v/ue+yONPWhXlgClWcvw8zqz6r7WbMiQ2Nrc4SJ1BlAZPPv49d
vzArI4RsrTcClu5pxJRUslmYxTBU8H1CyzwLIHKAaW7k1BeJFTCsHNLiRTdogjHHqrHuLQdpX0ZT
d1L6tgR4YeqOHgovwKB8mcqzdFLmNxBu0Q0qYyduW8XTFndeswpEIDAeN9nI46B6AkX6H1mpLTPo
AKrQygTuzxYGffIg8Bl6spq4+/k0GcZLwlyQb5UKsRzPvcvvcIu6t0uypbA0bmxsMQzWyi/xiY/H
4coWdNH11B+1HKfuUb85YqMdBWIq9eeSj67Oc/GrRXg+T3czJZ/zkDGoUf4RqAl1hLgEzDQzjtan
WDfcsvIB8PDfgjaGb1at/BVu7+UZ3zyJLspXkw86I8PMognB7byZFw2deCh9iaRx7BAR742GlmH4
vmDpx/IGjffoziQ1qSMYBV7ITQPoshoKXFPLN+rDRjf3yZSceiyQUZz7iATv51b65UD8XVZoRR1b
r84qdzo2raOXgxRKbqa2VFuLjXyF3UPNU0kIVKMRaScYAsa2pKTVQ54gXWhuITOvdf8yA0c8gT8L
1bKC5iT68bvourFFshgcbu0pznCi0DBNA0XWkapazteZfK9raq98dRTjGXA8tFEH1cretr4lNxh5
k2GYt7QPn80+52+V6y7tERzoFtL536Wx4obemXIFKY4pfnJwZGxCaLuWHnF7EkXuGZ6+ZYkEFym0
MtXC1n+lQFOoky5uRinWVZYDNJScNGCa8SXzoq1TAvrdegv6Thtjlcu3GC7VXyTP9+RhEKYb/qDX
EjgnUqVJ1tR2Tu8vEXzQ4HqSrX4pfhi906W4B/7vS6FvJ7o5m5T53mhZsn9qq0+D7q5b9WjWKZE/
/AxdZn/+7yP3k8Rarl0sJa8WtSJjKCH43VdizSnmfLOriiseQhhwj74GnF2YyWrCPoXqADINtVBg
Jrymie511J8Ksn4eeunaA9a/2KOKcU6+GSVa5+FsFuoaeSxttM+vBiiUm5URKUpRJzbBCSEm1ynZ
UYGXPMgl9LbRr8sUYzR3+IL6ABMdT/ZAOkuqjQyjtAsB40tCvJtSEdEvFVPBnowf9kfjnlQDHxqb
VsAy7vdh8RLLzjB/QcavPznFxIyWUcjGiIQeqRCJIE/pJpL1TbE5HxYG2vsrUOLYdNEW7sxnghuG
kTen4mkDeCAB79bA6KlTuHsXZAuwNiSgFBbtAviIa0LO/NfQXmKi9iHFw0YZ73cJ6Kfnq5bUZzee
1nqCDL79T7R+C2uW/PCLb33z1RiGz1cBARldrr0rnE/FymMg9YdMBHLYjw9B+liY/0uxiC6czotH
IrTK0mE3IaXPKSnLPlXMOFsgBORpKkAKCOLV0c/ZIteIOzaAdfUO0Xi+rJO9gLzqosmO/u3Bu+dc
ffB5D1Crdn47dNb7f1vT4KwW7E1iSfhaWJCODfqU5jCr9EWrdn2eJDIvUSIyvS4kVg2wRzUvITbl
8nHi8NmCeB4qmjzaDc1jB+rLX+saJ0c74xaricTj4NSwjE80rceRMi499xeC3yMKwLVrkIlrXhbS
NMNrHL83FAVD9rAAlafieTN0uknKWRL6E6AFKyKOZEJO1uCbprurH1k0P2LtqS9/uo/9A6t7Vw7x
+mp6ElUjJxefAmKH8zz5QpGqt2eKzgG5GUh6nGyNteeTzO1vQSm0pDxDjErIwOMoU8BT0GP5h7Du
ZzvBDEcQyvw71j8VYzZLH6GwihGHSqulKd3mkM1nC7ayKdfb8Xv2FwrbX5NHr01PShjjLDyQ+BR7
jyhaPj3QvVq4d4mvnCS0ADmDlbco/9hogQM7KXf2lIJ/64G9NihUEiqXAlja231BTqaKrcKlccqe
+F0h5xcFhpF99ETildjG+kjH15Ene7HYRlUIlP4kbT2jzpRHLqiXOTBNirEWShe1Pew2G+O7Pg4p
FTmIcqoxSOl/VpmgSQCQU5je99d3fMcaYQ1ikaRHOjDj2pV9LqRVt/Bo7KYO3Eqag/6xJtrhZRDt
JHMg2l0vXQn2WsBmLZZt/PQpokP2WXkmhmZhEIS1aI+LlCMTvz2aDb+zVUabbgcWCs1A7TlOxyUx
2hNhxa6Wef722JYoFSFnGfgoQVd7A4KhAMPpA0Jb0RQgNlNkjUz6Ylr+GJZcLgJntncrNqu5puhP
ITq+Aa0VsqG9dKo6l9OX0luvIhhsYxKz1czRW5J5hx0n7ka2YvsZnZhOs0IsMJ0nOQvNpU2hm6Tm
DkB99gkFM2yLNT75X2qQ0ONwmt6jo+h14bfTvJGWzWRIWN/ZtkILCsiRU/p6QzLm9F2PKSoD5klt
8FCqNLksBFYv7Eb5tjYhv1kQaXwpyscZvS7jO5c5NJ4lLPppzGOXyUMZm9Q/Ivagx/kbLD5Gk7q7
CU36D5v1Zt3ckESbJf3xcDdYZlAcBn8do6HgsascOZbOH+bcqcj3JB/vAh/XfisAeRgQ4HDL3zbv
SDoYVAO3+C5BXrlyWxbZ0+/FIJ4N7BIJ18mo5Z9l2V+hgJqptHyXn3QR8xy6ByPVVDgKImCrDoeO
2Nx0+OKMFlHSIIl6w+QNuL8IbniA7bpgXk3Jss5DADuYfuzOOeGPqJljjQvH+o6pHVmxQoqK9K0k
D38+9/Al2DHcsbo6GUY0tjsuTjwt0tQys16yfnMyIKsbbJM3Qkrbl5LWzFJCa0zegsuZtPMgz9ep
q68OWgbYQFc8Ffi0CAH1cwUR417Iu8uM4C3sAtyz/Yu61Nc6/6j3X2XclEYHvM5JEU/qrIL2+4ZU
pOxJD/37DxqxinAxYTp10wvyIyl+6kNJ+DR/qn7HQrmlYS+Ty/E4PIXXalznsSARpcWB33CHXkRT
3A64GnoS5ZL5tGHCj5wPb+VhbYil5FGojrZGvT86LAls7FtHTXyNNglUnmrI7sqpRPBz6jPHrcXU
yoMaRFejID7bgzemD+g4QQCbzyxWQ7vxO0qX+vAHwWtybOsknWikA+jTGuXfMG6OD7aJVerlCVNI
HnslL0l+yGCU+zOnwXQdfg9BPXLRxAyc5eMryowfPXK0AnrF3UgfPCt71k0nb+WCDQGNKeQ2I7w6
4mjIdZcgamF2NHR7NxJ4VsxMaDiM7NgWXrVt3+w6MH/ILc2i+VGEzfBzdjarTBp82sKVrHgVvs5v
yVshadVjjzzLXkuHt+gvkAmmQh4/kr1li9OnkgTcm4jw5Mp0gYbmYO2EjJ1q93ESdpYx5TpT30j9
nAb3GFc/Eek7CDVgHXC/bOuuY4DBwUo5aBvvsQ9AnbJ8AAC2OZVw8WrSwfJUIDNJD2YH8fa9/tsT
FAq+8WHFeoQAwuLWY54LM256Ni7SmUKqMFb6gJ/cbkNthamkv6SCYWmhICoshpf5Ghqu6rxrBfuA
zfgC+/aIjOEwuikH2f1ke4QWWXY3lbjM9DRALmF/N/IVqF1HBStzPWbms5Vji/sLLdY+fOGyc6bH
Rnckb+iTF5vOsoI52xKfJYPdyY5Wz7f6EJskpe42usPPah+uBn46F6+ZlRUhcsJ4XtDYUdoNlo+7
7N4aLRd0j9lAeBTVckxcyhHbUm4dgKQg3LbLKMoytZifsSwDVaRsiDJBvTLpV7Eak/wjXTPaPJm8
ox8oC5tWbDRrTcpjbg6eduC0rp9D0qioXXH/LGlXlWk5VZX0IMEMGdqyspRm35kfFdUylrjsDy6k
4mUTxjFRxHqTgOx7tB+itMtlgsB+JqiyOe/tKAzO1IZZGsIJY6Yuc5Jy33ea0qXay9yXUUKyadA+
yb0EQpwp2te5nHT9/g/6g1ViN0JTnbzcxL1A9LKeAiUGNzlFj1TWUhX4FSs6xOGHXSTA6nOEVYBX
MhsPYUxCvvTUDCBD0W6iVsydKZNNsZBuSd2OcRVcyXh2g/Zr+RmrGO5FBAFHaikMhgn+/9oaguaz
i6w4qChNxY2mW7OiLMDU85L/xW3LA43ZPSu0PTjXfJ+rrWjPuN7YPrEF9Hbzu2Nt1dqIVgUd/VHB
2Qr/pbWDsju6ksz05KmF9bRh/d49VuqeOKhrTiwktyD43ZpmQuP6hFiuM/npIaERsRVcoSiX1kGj
UCzHmsPqzUN5+63Q+BbTG6j92o1a8Z3a/cRkrB95eEeasw72rFNrgAnhbSIfZy9Hgk47vyIwNDb3
ivpohqFEQ/pfEvVIFs8CgS5+BfpMStvQg1M2kY7K9NGcF8xiax+7W4+TTGek20Fg///4vKSWuAJx
ue1fQJLmoROGIm+NiLyKGKelGTeXVESp9xL8IwMTFlmziAEnGBbPdfbiWIuwW8rsVYw6WRLGLmoX
evDVBUO5LHOLG/yk6SSPzCCHvfcrKnN4RD+W2iCQdHMriC+mQcRBMCfQmaMDHU/zFNY+NUOJT831
A3lREUTtvBrXn8KxdzgVEAGG4OCJAVwJyJGubtAhNDHYvKY/wexdMSgMPkEChBGrc+GuWrp0O7+8
p7+BvU5lFBT/K2K++hnBtTYDc8kiVTa8CRpq5wrlzcfLTD4bVroB65sAR6rsCvT9bJS1CE03jZaE
doG7UfCQXkji0mTOeoFsBxVfUqgO2AbIDRmMLI2vEAMKcfcYeQVEfT2mW6hbIWGIbW6fxuluTNoX
hVi6ZiRgg/56kYIjSpsAgfTUXPhd9LWJ+hUqJdxW5ZRHcksuA0OrzkOuBlE3S1djLTAkCE7Lp6g5
/gMaPW7YmsFu6uOLVGMGHVnqfkLs85BkQfVZON7Huo37+lMteVEP6eaECHNfVK8PClScgG7rFMlX
az+hj2b+B/hDD9OYtvTPo55cgXIXM4mgBhwzRW3Ew1HyGl3LioRBhKH9IU6y3CJk8QYUevlci/ah
S1vd5L10qW2gm5mBUKAtSTChUtOi2epcA2bP52I0FqXea/GQom5oO4ZqQeJL40irAB4D3Fa32KF6
ITFt3B4m1ake1ZvzVBkxxjdjnpYJitqYFUBBm5fX+b6l6m5LcX04qTBVfhQTc4ip6+UUKZ2M4WAU
tV2XGLK4XgYAd0E8mKZtvFJtSlpIY7ikUMbU+DFvgE5z51hVX7ytURmienZG0spiF68B9SH5sGx1
UovO+MSpfeZZg1tHecouGY4zgKCClnQ0bbAfrWpGknSYdo7dXULDeayvXcOE4Oh1shbXhfveyf/u
JvSMGmY6PknW8HPyCw/WWud+uvIRgmTXpsA7OjBbLrttUPySB9CElq9iSFcv8vhzg22Wx0PrmMG+
nu3o9/4/5KXs6C/nGu6e493Aeh8vdJ3bRqNgPy6vPEvuRAiueQnAYXHQkgSjslqPha+SK1DFZl2t
Qa70ccqJt5KJIqlr+mVP6cr84TR0Z/29n5DTZoBBA8tgqVbgZcDRPcsCM7dVv9bQW7bW36qMqTbt
tw8BJP3tvI9dpgzw2xUgyNEwUDPFNFTpQgoV2hlXkLxM+Y/A3XwzFJg9/45Dn/TAqzPak9O7bp2Y
SZFGoqcUf3guPcFDWR4O4BhKrT9ma3i8R75/CQUGedHiVvfpipqd4img62FfNGCwyqMUEbAqnWST
pwph94bsF86Ky2/wEchtWvtdr16NoDeR6FPfIOz19mpxVyC9NlxjzRMKY10ZNOsMJGClyb+y7K+T
zhHqrgRrniTmvQLNl5fP12gPEt3I7KdHV1ThdUlBUOYimeD6HF4ZIgRiArOQXESPoEDLeg3rNcTO
6I9K2L2XArZoRcJlIctabaQ1kaQgvyGPIEEEiYHOi6SgzCKhupPJoiKuxBXHUFbvHK70j1kHe4og
DC86ZN6zZUSruvuLjQpakcRJ9BqKpZrgKySSI9yaUp51r/Inz9NJqiSL5ifwtpWwDgAQCduqClxM
8/71LzM8ePV7Q1SXLuTkcYE62YkBuWSouPK9+dAmDXaVwms+Zysd8PdPzduJBn2Bom8r0GSNhOB1
gUjsH1eFMOmiW/WJwgfwQPoIN79ZyMnyj423TlTQY3DoUW6yGvqFHCjtLwHu9PEzwpGU51QdTUsR
kJXNfLWUcg62Sm76znnYTaBooO3nI7hJ9OKbLEpZKo3U2+4wJXO/ywFz/FHbVcs9+/SZU3bbxRHS
VVwKDT6na9GTYOjGSgcON1wkGFLlsas0SnFIQ7rw0I6Pnrra2Jtu5AQ5n5zC5fuMFsFXXMGugtIf
F5UBX9QQZZN7oTKV608WQDpAx7fgX1TA5QMoY2U3vmUBGNohsZiWMs1CIV5TspFwzielnBT/J0Tt
YgPcY9rMhUqLvF6tFvrozoCnDziwHkaBeWvZtSZfV1qQVH6tewC4ZXJlk1V6bv/4v8oYdDdnPNOy
o/sqpG0HlVVxyMU/hCf0AGIb/VvCs6+t/J3rkuzKRsijS6Zbg3Fdrm8gRZ2R9CnsKU3BjVvwLhpo
N1ecY96Ysn5DOoUViPB4nUXNfYR6bBsn4HdfQ12HrSXA0+q/C7/3aie9m+4+w9YfUyCQqbWxAOut
v0att7sdF0WZMpO8T2qeIPyAaYJdFRcbkjw1usw0A0mOlp0qAhYBJyUprEtGWE8+J3MouH2lG6mA
MniYB7bq+CQEilLhWJIxetViemp8HmwvnCIDCbGnBq6tq7Z996erLWZOYrFJvb+pHjGkDpmdHIXQ
7T40x91+nXxOGEPBqWPX/hz9WeR7BCcN1pDx0z17elEFIQMffo/fa1LlhTDhFq4iM0UCP0JCXUHv
FEemxtV5XOVzGQQkUMLlnVWgJm9pgE8tUobRLFqFSiodr/utjpOtr8OEWY+ZRZ7Gzkrmdvrz14UW
Lp+9YhNQ29+jHYF3FkvT5hT8cHhy+pb9phTWZgo6M9JflTFHyjt/GqMLPMfCdAyJBUp9xnQsIx4J
I7rwL4pjcsxEwVLeVUzSqBcQw3aXotk7TEgPrM/milNQoB9gfbn5xYnSNvR/JAdGZ029h/OysZe5
Tb6Rx8AZYA4DL0RozfLnisoTMdmpMxYIa8uFc8jMWgB2KV1y6tOBNTtIEjQw44X39302ZgBjXA/O
aOESetGPC8nozFwdPiv1SZiS2HgrX/ofaS6Wd99zrch/nLBvpIAcjtO6v9W1ymgZ1RrxdAihhaGg
N4bJApf5zIfGyUHFtd8mFlxXfmsuFidMghdf5/pfEacnxBUB/rIIlf+q3/t3r0eC/oYHCf2bniKC
9+QdPPQMAd2poK7DLcBATqQgB+5r5JU/kwivHPNoO3rMvv8upSiEyv1WMVKmEnkm+6cso6jHr18z
+2c+mhic0lzZcaVyxO0rWI90tpTPNmloBJh/3aJlW1hdI7sBboIut+vqthvYzAo/0FbZtnoMBMps
mvKEBCm/IYW4rIkiBMMFD+1T0CDnLFi3o+/MNVFsmtIUHnUv7gPhjHWynsTYLvBD5y900DCxk3rc
+Ja3ZL+U3wThQLeBipiWrDLGURgffGWCTFztwpqKUG8eDazPIB7OGjSi0R/J46ok6ij2oX/3iJnq
RC0l9MCgIY511l7oCQmFBlj33+gr5i3TTC52AMhVnm4LnHYfSIDCwJ51zkf/KnOwPAAyYZRRej0L
OtS0iI5fMaGY8h7HGgYNDkocsBOVm9y79dPtDS+vX03D5ECkNeCUWye8zlutshJe2WiZaImRIlh8
QeLwF2ImvNzmJy2KZX5kHtrYITRVmO35W+XFSoVxomEgCGO9ki569UGPVsuz5rx01hkI/6w3yfoJ
yXSnAm+vcm5T86qnnOO4hrGBVqtYlmWKxMr/NWT6DdA3sI9Z0HJH5fQ+AOvho48ZS74rmgxZXf4T
oCUD8uk/RMSgx9NK34+fdeKo+8J/5InBB9zShrvsFhGaz5uZrRD7pvMPEHaGkn7Lm2Cf/QmBDZ8d
7wGqIr5lXovXn907Yuhhc8IzLZK82gkL/1BZT+tOqpJOEBgG2ROESr8fttjw4Xr3ltURMezkFSKk
8D4/PW7QDBnoLWRt9BBAZZ5L8bZ3S/l0ri8Np7p+gYjz9+cXVRvCobI+AJMnvp0TfEtx4K+gR4t5
Yh4We5eUEvfeSzK1QpoAKvTeALQSSi69e24CYUH59SfBzfcPDtI+/zobkDBi32aV/UAoRg1J0wG8
mRwGQjmRDSfOdIQGMATt8J3B4G/BkHqf1QaqD8Fp15wOZ89B3WtoEuQ+y0lpKgiijYMzZfDrBC8N
8XFQyv373esc3m6I2VkbkblaF69vcHskp8L7vJ985D168bhqZODsE6EbsskwuZfoondA9ba/qOIK
Ua7mY2EOsonE9/F28LqssaSxWMTuZym1tb97GwRh00jNMv0k2AVwLq2aANXILjiy08ifS2eMh6el
FWuSQ5JmPfSzvir5PFudGZNdRM3LS8gcmXtDsGNLGYRiQT6t8/wIej/pANodWfw0JkBMHN4+VXuP
kf3XkPLzy+0yvmwYfNWFSaeB5xGLI56XhBvn3VmnC7fF9mQ8FMbq6aeawOvDKn72UnBqSLixpLlQ
edgw1bNBYGiLjNC2bfsGHKHubj/iszHt/wi1PnP6dCa9oHQHsCJVSbEUhsLDgoSP3ucXQjgUkwhb
qiebPeBbC2hx9nq0DvLGX1rcWH+QZUoRKFmUJRxtY7P8ld3dDdq+lLeeTU7e8gJF6bBOyVVH+M35
0C4tHalZhjmyGHwOVAjxrXEVRDMnYQsInT16aXZCz34NF3ihhwMv+NW8HOudwjxyWlXyo/rHIFLd
5qNw4eZ5qMK7FHiTlClyfcssbkADimg8ydDd6ljD1ceOS/djB16z9mYCuVsifA3CjnaMANoBa27S
k5qSgvjHhhgYazR0oTgSD3brGDAeCrox3aRnW64OfPZIyfCGunyWFgMwWV2VR7l6J41AcxiYelxK
jnItlSerHo+7fQuSDw7u+A6d80OKngJS1Q913f8/HUDTDErh0cLtzbK+fAAEbPqQ5TUfvV3RhA8v
zL5MN9SakzZnj86zlOKaYZDuxxD7//0Kkl1tQM4dbYHEQR2hUcudpMPNgs60welpZes6+ZbeiOaj
TPrwA5ZY0ThS7AieG0MUdp6n0Dm4C2BKbCTGGdVb3sZ8jfvXL7N7/i9suRYKgHoBApld3Rxc7xu4
9akF1wqfb/zI06Z053JV8Khys89UYcKcmVSePwjwCiblFUuZz9b2p/U6OvX+Y7v6B+cp8L8V6Y+6
ZFK5Dbvtw+9Rs5RKuS+t0KlD7E+4SMkFpvzQYop+w+Q2rmoXbDBcYt5VQgvYkrehfIM3JSKqGilR
PuI8pJbiYFmPR4PNzuL0SNASrrxKGuCAeidwOCWmy6nHX36O+CzdsoH3eMUhErV8ZDCjPoIiNAKU
UYzcUrHwimgPxX2BLHBQkNdbQfc1hbDCZ+17kqKacMWFQcQtF1mnUUDR3qSm6OB5HccXplyu12o1
nwM+disKB/WxWNE5lGklBxKKwwJCiW1NYWfO6IDOQisAQK/qRznFOrs8wR/IXT6Ow3b0LdxUxM15
ozDdVRTiv+jqKMDe9p3jc4X7DFjGN+1cyuWHLelxgDMI/7DK1t95HJSwfZ6fiAjYu2LRgTfzbk+I
/7iJ8B8emV9Td4JkxA8nIT0CLdlhN+k5dhNuUAE2SRkpbmHHt/wF0h7pbVrA4p9XeXLvgBNApqhQ
h5ROMv9xg6KtHJPgjpBWg+wOKY8lo2mMqWARntz0d5RaESPHYErlWVWpEDiOy9wXVd0so3nL1gfn
7ixN2QIIly79b+nAkWHRU55HLV1uQkw5sUwWd4u5SM9ughYlqm9RrQDxEWAoC3RDFb49elILcklq
oBg5J/m4zIFkhm8702YgERdMAJw6vpqiM18LDH1Tk7GyMkf6ZktKzIvZZharwAu/agGBU7hg+FOG
kkB8Rz51cOlgml+uSDNUJ5xLdUOTZvFHpLCPJybir5HSgGjb2uE4Ax+uld/hs7M69aN9P8RXrhmk
ziYmIddQEpl/XvlDh8yapymGXA+DzNAemq0RDGq5LX8BrC/gftXbYKdRWMdU1CQAnr5MH4K12Yo4
0vnmDqIYRfzFeFcjPDOdgVTlSHDJWayJbDa1R5AvCJk7LGZLb8+YH20iVVFa6S+3Z7BkmBwy0oys
Z7+0yTC2xic+HHxw2eratdDKXxk2N6byxt+dlxEsBHXMaA6a9t9crCo+A5JTD32KGf35mcDwVd19
MViDyXeZXWojASKfEc18yjJxQBNlXZtmx2tt6jTWZ0RG4V0PSFDZqwMfJDyVV04jaQ6C3kDsv6Vu
jx7dbKWYUj08HakHZ2HC/QiNxciVRgo2UWpLd6YSjqGxLgr5g23TJ14qAP0C8sr0QWyYycOz6LoS
/cnFZzUqC7/DWPgMCzsiRhbmpYirQKGHLjU5NkTzAp56InLr7TtWJtnKpM6NxldLjXn5hPDflTsZ
DGoSKhiZMbk5inyAbkijZesRAwaNOGGAxBy1C0l4o6Js+mn06nPpWQL+M6b1HDtlolhbulDHUNLD
W2APvPhv0XyYgMJL0E7Pn2IGC2NLyRX5Vh5tvH8AZXL3ad6iwImFFAuJDFvEW4zjknkMROPfe9Lh
XXTdQxwfU88tWkVSImwRQil8zdXXXa+E49Y44kdGSaoKMN1baAfzjIw1BtoA/805M9sjRXP0XotR
3Ix/Dt0XIfcs5QqlkkCIVE/9yI2ztx1aAPyttrf8ogmAsxuU3ox8IawEk7LSCvwMJAldotY2/6/w
75cXBn53Siph8a4HFPf2//Vrg+TtA91VxsCvQCdQOja3kjzyqFvs1/rXeVREwhFxu4lsiJffPdnf
3wVorF+d0PHTrcKgQkf7pc085dt2eU1lKsPvzoRp58dPNZkQ7c3T1JmUvXBpAU3yoReGrDzWNIh7
JZ18pWyrYTFIM4l4ulo6p4OZkX7WZe68iP97r+5EoH4yzy1zFYUtowb8yYt73tlzKfEqsxvxGz/3
n/QhSlSnAK8iRnFfXxE+HtP7qr5QXznFEPOJqfY2U9wkondFqAUneWUszBaT58HTDdohCTWXWYgi
lqH9wqA7Y3mcO5KSx0JklM8emfzVIYSryUhOR0b3v8CifcKJY/ah3F6PTnx96PZ7LLuhWSMtqR4R
/CmXgij9K6gHuaejO9atvMt1oORqhXLUFoLJ5wDC2unmSicZyGWj9hZjA1473/3CTml0C+ZZUxl+
h+TLUkpyAI5TctcyCDpNpwwXMCHAHdIMBcMjT9LhKwiryuKjHTyQU0ALu+KCh3fqk+Avc/2k+mwT
gQJqH7s/Rt4nPYNY2EWQMmDuT+x2MbynTILqwF5wdgR4PbaR+ZFjDCeVaiuyqPuOWdFqjxBDzhmy
CJ+IEzG6/KU1tjpt77u/6JPOuNpEwnXDWj4lX//VThLlY/JWjCDuy8WTkKa7B2gBDkFYcSZm2U/f
hllD5qj8QfLha7fY0mQowWaIbjUxoJN+W7mk4otYHql+466ibz9soiuvP6cqBqvFa2WM23wU8N4R
C1Xe5WoEhRnN+sc3prfx3G8Qc93rQz4rn6AA3zNVqF91YHb4qk3UlQG3X+O5llBM6q1DGt0d56b9
ZXoLZ/pA3TV6EwpF+xR3AqCMMHlQ/5+Zbk9QFlK4cgTC+4iua/g51HlTRkF+oRoZHCVFAqYpubQk
oYOA7L+U+i7uIB/BgW+1lUzCBFEo0jVU1sILcLe8PtKcqFAYeXKSITDQz4peRtGY12mOA5X2jQTq
oodb+5Cmoe+yd/udpct6yGYN2EPYCSUbKb7Yz1+FeeXGBzeneGBI0uQRcdhPYcfr0sQyQITjPjjw
t9wFjW2PVIYl4bGQyx7xXkwekorRlsEv5XIt6Z05M+LUzHDPhP7vQ+q7MzYbDRzXbgDgJfxDELLi
VXPv90pidZJEueZnkeQAkL0rCgaxukRhQNGEOpytaa4tJv9opERx23yFE0wEuyu2TAs0KPjIamSK
WFlXO+BZqesW8vrFWkZNY7lj8GuGOYhYibTu2azC+vb2RTKdxVQzVNm4hfK5aThHWrc2CudCvjAJ
8A414Lv0eFrhTZ+9BhKSJEBhyx4pGT8GwjWW+Ow4if5yV6+eMRd9VhRglGr1qepUDjGdsRl1Ylav
HxgDrzr2cXPECuoiXkXazUvjjkpXjVBXqJl8QEOZt7O/v82VpyccNDy3PUzD9dYHPcw1Tu9BGseO
IHTEMoXGj8qBO+RlVbfPJt8ZTuDuTNxaUbBYnFi+gbTShJr2pe1zzQA3rG7qdnDSxilmon5y9bDq
6JSR3yfO/ZC+8fY7W/HTl5YN+n/yoobbhipEllw0+MKOT07w4w6+FU6UkPnfy83Hbn2lkElAgNrj
6I07z1wsntXCvZxZRELuM1tvB/Md+VUHUzsF1Ln96n68gdYl1+DRXPGPrx3ebk/9aUUTHqypzMES
iKpsSolx0jz+09u6NMC+QDTUbhSAVql+rgUD+AmuWKHK2fp7bW/oV1V8bt6Kw/W3jE9Fdzy2qozJ
dRrjXmWH3Y18T0TqBuG3xPPARrDRkPyG2jQHEX4oI/G0Af8yTOfkwo1Md5fNTyk1h2zpbcEUguQ8
/jnXTwiBWp63z89zRtpiMB2Y0WWyNuOn9B7qnVJ3gKMtjFr25QNBTmPeIaF08IqKPBF6ebGM0Y64
JdafSi4EXZEPfSpe/c0sjLrbH1tQ+iQC3tW6uLBOGH1Yb1+LuRLUewMeymbtrxkEXQQoP6j+I/8h
YSOkI8FFLM38qFU2imWaG2nZO4Jwj13Toml0dwhIHTKLffm3kc8j2bVx2anaUS33+MUpl12CIgYk
1sp/HzYggH+71to1q/UQlHhb1ehK3KVekSdme1MTZp2sSblWQapMJOEfBLVsUHB8tLgfwmCZtfDW
q+hsDzOOBOiVgwae9GDLjtDM3D4PBiErn3ZQoiTsNcyU4YB/vol02EETrEJJ5TCXkKUkc8Mp78+I
FCUlmwqIN/MyWZWdk84GbSgH9moYBUQPNaFllyUzPjxLb7u3B78aB8MsWWSYTwi7sQsZ8kjlnsl2
wPnNW8s7CNl9siyTi9zD+E+ZfAXkB6lz3xcCDkxe2S0+YZNSnSJlFIz3oGHnCNMVjAkammAuBvZW
PGc2tBq/tqH4TL8HOdpfg9fvnd6UFr2X/MkSigzOUTBMLQ6pGbYK7LOQr8M1T3ie06qne8GOrkbO
DRp+dhra7eFjD1JMwuXLyyjjQRp81c+C2mFcPZXO/Fc5jvUv5oH8fwq5Tb8xjVnoCIICZvHcswr/
yNao6gchVYAauFf5ggrkU9AzJJiBzzgSUy+uC069G844KjUYhD24AaQcgPzktfzdOd8o1Q/HWCgJ
k1750dM/ko3lJhOsveqkHvgZ2a9ebk67zWPUyjbaw2yJUp3be8iRE/ysBlzk/9+wLEKXbleCkQoq
X3dPf8cpR9aQ7ZnE8QK8dadqnCpgenbMcxtFa9/wFylE1I5nEQ9plKfRWROQ7KDysX1u3bBLMuPy
07DdwH+5gAVDBxHQbTTHGDeVeu4EYhVFfzLvfwhll0Z9n97z7kvS7lqjNLy6oF8P6P/NV5x8qgGj
wpEYiBVUmo59zTbOancEcx+gan+rqEID+Ie0ub6UnMdJLK/VwI4THtKZyTMj34EIiUbPfq0cKX4Q
ccM2HGVwa8jkYf2jGoVXraTjubQPeAsjXfr1epKx1uHxp7+iM3MTUha1VCzevieUTPgZlCsqywZy
7q9x4Fiw9z0GkhptAAKh6T1lmRLXnWKxFj8eKOOgVWktiXG7Z1yoKB2yxhNHBMrcl9+6zzdbfGFJ
iBzm/Vx8qBRuf1N5OgaqWl1LIHfi/zmPUFLdAvNBZ99X+TBreVeo4GdM90pmWUg3Q5XIPRr5kK7B
Os3IQDy1JojanYsPAs5YI+V/RXIlwYaPCO0kmoR7atBVjJ7lLtBRVyRA5Z6Yqbr2XAYohwJVHKNC
0sC8784fSgt76n8bw6eOOJ9fBWY2c5W5jaFVecIcGs5NgIdj17faGVYl7KryUcLyxcBylnkbZkK+
mmeA2KjJoAztafEIqyw/ba2fVPL2JUPB/q4snGrH4CsgGvqIS1BttyjCtXNy/9uDXmQNPQKVCUXn
PAoerEk47OdpDPmAzGzpWClOEtT/f4tE/VQRzmHbkte1OMXvn7+35jJyAdyw++1n12wdiA4syOsS
AlLL+1itR4lKOr9mNOD8ohNrEHmbx5BB9K52vxApuHBkuJQZQ5zXSkQP4QDcV95AwQ2Y9g83Clnk
lqqCAefwXLhnvamP4S73B3HWOuxSCYy+nDYF+OUpncVcbWOHkodSl2LB4GgOjj5D/sEJlGguuEi4
VPFgHYINZadZ5PGWCS4MYLIAgrS9xgy9xU11SA5BLTMzoSCoRlHD7he+SX9kwl1XNKmlwdy2kHbf
hIugUfLuN7o5XrXCx8NoAv53uuD0P8hcuRsgVX69ji+1nUsYJDFft3QTESYYyLM9MwFai9XLX8id
K3zgSRCXXWEEf2bwO4I6MpP/H0dg5a+XuvwwqinEWT5wJsWKeIEduL/nD9b8TAq6fxkJx73Ypd8O
xBUk9/3UTIStrRou4hEVIDuRXJde9uAHoUpeOn4ugoWcCdK03MFmd89BkABztNGHL21Cpvv20yhu
jOtu7smhGC17kkOcQGc/PwS6qn1N2E0NtNYwgjueqY3h1U+RmVfqNWGIRmGzBgLdWYVxtZeBUQn9
HQSlWEJUdDJyt3twSt8xfo/Rzbsqex8+PP7Eh1jyAnBAZi02sIsa+o2gylQ2C+h+NuIaLEtGlapr
+hRKiGVrDOvunpbx+Rp9qfTvVj2fKVJ3Sgc9+LQbOVVDsDSZdsZQmP9WCRH2v41AKsSNqq/ASkEP
asEQ8qOhwj07EnXOdzlcLyNYD8RsiT2ThvsVXl3RFVYINdJZU6hDW7iPfNv1gOGp+b48YrPA99Gp
AvGuPP7+xUHBIRYpo1nBQ8IYRACmDZ6e/QjSqy7DG54LR260hD01YmLR0xR8Urj/iujOhIW/V3ia
FF/k+hZHzCnPp5iUEnR9k/t32tCu1PKun2gkjIu+9K9MQ0VZsT/NBPeXyFPTNMPG4PuP6CfO8oqu
stdeMOMDycjIC5rlMJWpt2LJ618ffa5or9AUCY3cC+eIAkjvw5lHAPcuQsYzbvMEsGS5lVWS2xu1
TKVS8O4xWnxwcrRUg1KRFVSVpAIUyHFbL6bN4xRDMTthI/+FiFuzeNWULnub486D/xzEvhmYBQdr
qLyVvBlnn+qB8gPBEDOy1geLAmqaSRQ/vkT/bDRiKCvjYzvJpvpB3fbKuMBQv2Fa+jubxoHvyHWN
D+Rl/BjuaCvN/PV7fsVxzeam02bx550L/HRX5rTKDop21t1EZ0+V9PCjHZs9zhBIkBVvYH53deKw
aBNRBtEjUBjscI7+5WtemrSbZXMLFpFHL7QqbvjpE1wqlaK7MnUvkno9lQUGgOeJN50G49bm099Q
YuB9ZRNJthqLP6HKs4mzeIV5IeNULFGmbBXIKrxJWLVJC8zQMuUtrIt2vDYCsaBoNfl4Y1Zcuyi2
LQq4rfxTrt2jbKLR+AMKmeRBpJdLE8fxMJbRyVM2lKlHCT3ztilELesHjldQ49qhP2xRUkyE+qiY
XPuPCS/0gq00I5rPh07eDhEheSAap0fB7VH9un3lsASZBPEintBEE1hGhviXtB9KrueP7La8HDGz
E4+NK5UTR2D8KmTL1qvDlKebDx7IO+MPk+Az2Nesh/AvCFXE3AuKcpfnSm4IYOhDlG4byKfLhcGu
ky6ZaummrGbKSvP8cFB553bMhu7oeJlshxxz2l7CTrPLQ3uSW/J8f9TnwpVJGmdFr4B/XUTSXAwm
Izw224oOQ0R6GiMZQvjPpxCe4HhIwTWCiJ3EA1pV6sMssJmOOUREi3b7UU/fQHk2+PmoJQlw6YkT
ejksrICL/j23nwn0aFHgG09v4bIUK2n7DRuPU1ZBgJQ3MQzAoXDI+sBviRr4uVJQ0PPPyZ0XuLAj
X37EdxJnmV2DQdKy/y81aKwKFQpMrmJIVE4Ye6Z66pD99iu5YA5RBYJamStxzYm7YjrFUiR4SSGz
h3hcjnjZqhZqP5PCFzudqdeYbrqNWTaD+6tZvAbhyxvwhmayNG4Uuebhq+3u4byqOBVnnYXB1hHg
VhKkt1QjaNzJo0lcNsHgfKphfhHgTZgyn4LfMsiIyoyoXC4GQkolU4ZmwjCXBhsnr0wyB8x0AprC
OLjwMFnuE6eyl9UGHijoljFCvpQXd3D0HbLLv8PxZ7+59vpmvy2M9v+1/tBQOP4cpV37Pk4axKy8
6INqyonKyH2xJPWxFLnx+W/hx0athhMJvhzVNNWL2+uHUkcPcDnyKdRNMfpCUarOvyowTvLKeUoE
/8Zhd0mbl7OxeEvnFtHizqllKGAVhfNg1l/d5rnh+X7W9Jf/nOvpmPSPc3uvAoIMU0VN5xQgutSv
mziYKCRCVZR58lR8F54iHuntwDFQiOFbyOXGGqFDwrQ+1u/8D8UhAH5Tuee8atD27rlGjmE6TByV
mfup39vDqgWRNYSCxxfwDy4yicCqIJjNmDzE3oLVDpMqW3AUx+JjVj/7putVFhr2yWwix4Po8bAO
aoCaQly1O25xtr+RhY6iFdiGo5WuApnmhgZUDmA4KKOjyMbbVgCC4AlfFLfRrZs/qUQF1ze+TSoR
HD9CDfne9XdbyS53HW8XUknt44j2cWU272IziYjcdqMVNRlgJd3AonR2bTaTRgJneSjTFHtGwDex
Qu2wnmlHRjAYAXbnC+RtGxVS+G2SsEFlRpcZH/PWp6Iv9EAdtaNavv1DvbMZplmdM9+G1kkReLQr
xe7vfavYWoWuR2ufaYivfzZbLYOzBXLIBy2rQgYWsGiDnxUG+aigtnQ0fJZVhWWDgPFm42gp4A4O
lYTrDIixMm0sIyOrPWuRx/AtiCzjoouG8YnrzTG+k8rc34118mm5u30q530I3ZPN2WNHPo9ocpu6
5aqYVLSDmCJF2XgfpJWBz0h//tzL4nO7A9MROimg2pcyOv+mMgp3pICz7N5IujwtAMfLhSYqPHE0
Uh/HeQS38+g/iiWlx00NCUrk0Bhv3Fe7sHEpxr8iDCDdHvGSSrcK19gD0sJQFbpKhb5rAGuYPp11
TzFDDqtWkoVDMGhP6Rg0C8n0gHWyU2Li0lSHHuB/99SqYu3c0o4pgidkgMA8daSeKKicBwluP8Ca
FjtZ0DP/BcUx9/xsemNDYAanJremMn2wZtF+ZTH0FNfwOZlemZtC9oP0nBlydTB/ASHc29tqetCI
pmVUv+m4czg6GUAnouLXsOhDpakDR0kma0+rUfpMWHWgvAxgh9BVg0w6EyoUBdPYo7LzdhwMr/Bu
2zHtjdA2qk1z8WVGnTjcQhaDocOs/t2T1Xsitz2wZnRMs2oKvcRKsT2PEr6xnA9+HLtdAWLinicM
iiOYj6WrWNzUBi088LBVLhQddwToQRHf/bg1ZH+gF5URYUCgmHPScL/MVxfa/xde1otWsQgkuDcW
fFV+4fkIBoZZB0efLDSphx3KmtAbB3U2yFoox0GAIICxGpQxKgx2+Sirr3yXKS3I54vtsFfcxLNz
D/bNBrerun1SrLrNKQ0cU4ySeyhM0WxfLtAtV69CYdqjjZaGVD/cs/hvDv4raHa+hC2RfpC+pKr4
gxRxX/CD6LshLQrTdTKDgJBTl7iMuZbYByKXVimXLenRuRROZuae/TbOhosIJ2XzU9HBetan2qTy
fPez1wUeKQxInnSi5c5tj5t4n6UZVI7qjVuKGbPvtoPS9cbKn39/LsS63NuUY2qcAqzisiVCjoeN
R/m9g4Dxu3aGai7Yq44kWiX2LSbxgPYI08TW3xSE6SrnrnewE6R3EBS3BO0KarKic/h/nm1TzNQn
UTCarZ0pWtyO8qFvdpBeLhQwTB5BcepnrYaVJAGDwY7LFNYWvHgn3g5tBYwYB81iiD2iFQiQ72Sq
XJ7GrmUPSnHusdPNVawP0D9HhYdYTtzFypO3YXjRGM2qpAURsVMJeTXBMI+yw3B0OUS/YKegZZZH
K3dcmr6kKDbPgykRxM5DD+MpxZhLjKFeEGx1EFJSWJY7Yce7UWybTaiUZMErrzde/5o0wys9H7Q/
ewyTTwTDgci5q9d5apK7dhdlDQO/ovgQSQ0nmaQUK9mS2M0nKphQ8RFmPjb3Umow3cGKEgRU45qU
TwJ34vHWqPZPVJM78IDAPbLPwelb1f3UhtdujYdLGs9D2ozNrm+NUpAeiOlUzBKbfFOt+TXuKmK7
ZyGAF+UiOLobupoH58bPyhi0TfYb1FbL7sR5x+YKpAgYwA71iLiNs3WkTePrkkD3F/ShFlnHnqsJ
sKYgfnVlURS32JCMzbYXxKG+Q/JKt4bF0ZknSlnfQKW8hSkZth+shN9VqoHE5rUa1dDniMoDRM0/
cVc0cnyRL4QuxZ62RYbjMdtn4sR+YZ9KhjhasCJ2V9X9YbuYrBVR2OB8uHYKbZb9aUH2a4Vm7EtG
VYMYBFTBB+JZvDfota8Mt8XAasqUtTmFqLVAkBtfxm3zmyHAgvGu5T5l/eaOXn7AkFPZWvdZdkx/
yQ4GSViUEhewMTrClgfbApGvo3MgYETHnOa9k7liVSJo+t2QLZcOwIQ9sjbrrquaYX5RV+Eznfmj
EZOe+TGTZAofeFDRJIJJUemX4zk8nXfUYKICI5GcOSugZnjFZKG+KWxOxGmhT5dZZnZlc9+0f2eI
cNJ/5yCGHLTVCjgE/ZpIdWKQ/KQpmaI+4huIioHxrTWiz9t8tKQIbBj6RzYa1RFRVRs0flJwFscU
0EYlVN0cUI5hLbmxyC55vrvXhDe2tuBBiCa5WIEgtQg+0Fyen0sQzW4V6WSN7AcN7Uj+tUtqak3J
OOpdHAYWM6KHHGQ79XieTq7J9XPQynJlD20DpDkVdjIiVM5Z2DTuzULJmvj/ujXOpjzGLAfs6iJU
iuKNyXKiPXhCXG9YRHrAMmzUTCPhiQQBVAi4a4ivLjqLd9SkBUaBI9bKocvCkfONU/XQDOKW9f2v
9/aNS9nxjD6MhlfSc9wpnw8YjCnXpMM9TeKHv81SMiFfiZMHnS/M6WrkmjyEU/UkKG4NJKntPMaw
OPVfpqo/A3T/QnjYaIhJNgQvXp1xkx/FYgKaq8YURvkpN4RKVhD9rEQMWmaNpuTcyelYsn1JHJA8
gUkEqN8DrsPdq2kom2WRqvMn/mdoiwvapHjBjISBUnQ9gzN5dMDmQAUiY1ByoTvOIX2iuSogHq87
aQkzDSNvES398XPB+dutEDhdpP6XsXIV/PiNolO6akErYp20Y8JQG6eY7QLiX33rm6wdR+JJ4uKI
v4QdPa5P6W02R26niEh9ynija85s4vl/YYW6UR2k7UoDBvcuIxa45zmRPo0b/ejMkLBUdMD7mlaB
hNhEiL787su1aQ/O3AlI4vkXhAIgy2bY5+eq3fpeNN8GAy4SaPtO8xco1keKMtQFc2x1e+pLC6jh
2DOK86HqBDnQMegDemd77Q9Ujy0c91SORAllEj54KuDDgVin5a+XJC8ec3NT9SxNkk6DEArizD2y
KieyPRKu+48IJcv4S4redbFW3O7GmOmwzVAwiWMZUUr2Dl9wfbLSQJrv1J/+OjM9AglVOpc1EaKh
MJmtkJWwHLNSP7rPZz/D2oqiE0vGTlciSuW29/OU2mjNpeVSch0uf5rJ+gWQa/PJRP37ElwvL2cl
6mmIeVWaGTDw3O5SDMmsSzuzysfZr22+b7rXJ0saBk4wHgKKS52egXZ5B+4PeSBCO1GwDGJeqaRu
VSyFfSAH/75KplNhGtNBA4mGqipRg89PY8P3GeFLi7qkW6XZnd4mLf8vbw2B+8DWflKP7tQ0W2Nt
RwdsrnPZu+jDwFceOJ69Utu8acr7JRGL7uphJFrdnnGWbE6mhjUX4QhKJo+SiTqpcaBFBGH91aZ5
jpbRF/K+KOypYMVdgic7fnuy9NWq7ihzQljdjzouGQK6R0C/CpvSuXXxCKXXHzj7S1K4rwaTgUJo
p7TsgQctZQe/6OgEQGjiS6FN7XvysapO06FdW94EraTWE3dxRTaO6KnN55+u1yR4xu4S2ypLXIz+
Ccu6EIOw4s7fYkhpPaJV5yHQ3K7TCmHDoZUytNwSU5CTDFeEoSVR6Io3NPjDjZPwqzcaPA/RU8FT
cDfcGUjie1nbfc0Ie700OKyzsHSWivd8d5V088NPQnOQMGHcGIuYEzaj1lUR/lbv503n8Ap50qby
Qs9B3+MdoF5M5gK9gAN1IYiGQU6Nj3IRN/Bfg0dVmCHNsl2W7rnXGqpktr2pm0N4nwRChNC8vkqC
b2VWGXfn+WVMEtmWWgJQwWIixDElIhIA/tfSeRsIx1yfIkTJRwT+2FLaDToa+4buwkqDnw6sY2RU
07Mm4OFrpNHBo+2fqhbTiHUL5A82CxUfmkJ3QK7B5buw5RcX0P8oaizWbzIyXo8hiO122XvHqHqw
sg1wOuDoZtJKjMZfgswOrIShgjhV8LCar9GkhgY9E2UR2xZRi7cPCuZ9/5Tw2XfmZbjew6VwZPob
2qzRid+UaSq1MyGFdZObyLYa0wH+pnHpUIPSNwryvF2aKQlCDELw9FsUIWL2exq4wHD3P6gokcpF
et1DpW+tk5Wl7Sb7Ml+oFZYmp2B//VsBj2/x+SJr/4qFmfq+1fRDsjKPIeMyy9Az1PNq8hClii5k
c+MapvOMtqnIfgCcmoQldk2u/aR2Jvi9qQukFq2znLd/oQDdG894a+CgJXAuHbClrf3m9Qdy13Bh
MH63ZPxa7Oa3n0uIZ+Qfh9qObw5IPLP2nDrzYcV0auekJiiR4kH+6R0TKN7ceXipUhyHL1Lsqhut
FtE9J10nCFmjgZbxUwzmlL3PaxVQ0ksQyKscA7t1OVDkwtT8qkKZN/VBM6goCve7/fdTLgQQwtUK
O2U/XB34oe+RezuqtdtVMVGX0dGwwWIxWcqcwlj2chZArHCVFeIl3kbOjpaR1qt+nB5LhjBGlkId
R7PPj57l9QD2BDAiKTVUp6BIwpCFc2qlsjLL6iLU5LO861jl4XQGwz6cC6JCV6vFpkobJLZnSjqw
gZ8hWws0/u9Fo4QsWhxn4Ki3E8xV1PQkHlVsWoXzvMrn90lhZRjt3LJFWywi+2xPwA2jvHOctRKh
/8EwOUTBbCiBqHWR5OE/AXCp16WS3pBzWM4Z/hla3Vh7u8euny8dtFR9N4ydPu+P1Q5xc0Tpe1nh
8kxb806F7/mJJ7P/PZcYvmsklZrDkWplPUMifePJUF7xO/c542SmNpgdsZHNBMPW3g9drORBRtzI
PQZ73SknXLvEqlpoi/lzaWYxnqistdjNDz9YfPBjm+c2+xUzegR4+X4U4qxe3AciRdcI294+wemO
V1t7pThgZliLDKj0DXI50tSgoVhj1pr/r3Qs7COWTq5wWzToYsqeZcV3DTQP4PJ4rFWbVlhCLbWK
m5v6iTHUB7FKCAvI1GeMIfOjBtZZJ6eYe0xhAZfkl/Bb8XREGmbGSe/OVDxnqhC+vmktBQsMhrJA
3bFjNZvcK52wxAO/k1iAVLaOvI9LIanhzq3igZ3RKxyKa6Zg/Hls/Hguh8H9Ju6w1FDcGYgL4qpN
AHxMkVh2qMvyaq/YRG4p1ooi5COcEuyefhEUKVJ9gYZkuylHEXap5zhYI5Xz7ltrLv0qMK8jSlm9
SL5NgLwhQe+kOxd75dTuXJ3PuzuH5f8LgisXIcdjRMu8eM+KWiP/dAq4ckrR6kDs24FHYUq/ZdWI
MdvEHxFZ6b0TgKxYqp0pMVBybD7xPlAqaphDvGh5f5tz49vRVUhXTtyIN0fnWV6PVDTHYoXKFTMg
qxrrb6I7wJAq8dLiT1V+zM0IVoKyov8PNPBMbe9ewMux7+7PDZER7K/HVnBbw8zTLnXeSfxCzHJS
0TyVLLrw+u/W2OlDBFCryPI3yivSNJmTc+y5/egTAri6HE+DgW8F+XetgZP7k1pZ9JZs/qQFFOHF
qmUiRiGuG+kP/ixdH9Kd7CIR5NVwMF0eBoTFRqbXJJ4htaiMt2RfMBH9rFuI3npor3zfQIqUQsr0
ADshGXVWIQgWoMB1YHZQ0i4xxafIQsEpdZ3faDCPLmxWSNfAoZ9pk6EBcBuGEMeZ1oPn34D+0LwG
cneR30AiVPak2B1UbzvBkCwrF4dvvske6ipf3iLljzvQoyOLguivrfsEOUJ4E21FeJcq7g6XuraS
fZdWIpeFFJNB/2hN1LvzY/AtcYazKuSYYUu7wXIwGGHPKN/FGiuZnB6sKxTBXG0GPDo6V7/ivaiT
F3CnBy43+CCyB4V2lo4T/3acEwnaQQVYS/Y7YP90W5oPHLRwnIcG94x+VCnGI91WBhXV0Wvbi2gU
y2VO9vuZIy0KzY9p9GBmYMARrTLyzKizAMsDLORZYgSplP7ehmDRv4NTbXZhZhsaRljavXSEvDEz
amYc+J2aUBmK9qObPHLL8r7yE6sklWPaiSM94iVt7juImt6/3RMA1iuyfkXG4ZMJcMoQ2pAwyXxJ
atxVWzgAGRuVkccKne9i2qvJfADLU/6PXFKlaiyliMlD8yf/dGf5VkcJj+0wv60Q9w5iTHSA8gZH
9N62KQeShURXEVlIxX88z5KmHp5MGhQJkOBIbL7a1ajr99vCwoeFmoWpPmQJLEG+jK46PsxYF+QD
NYEAuAaezXkWBu27R6y8YMtG4TEyEtSrdoBuOLv0KnCHv9xoqlEppsw2xKujD518A+qEDKdeEoPG
YVcf/wojMoG0oA+3RDHAlfzeGzF5nuxw8aRX6ff/uJfjRNBJTlvCvu4nTgDyThUYWyFGNNYrvJ8X
ZCj8ZNeL1HO+5ZSmPzEYunKbkSRjDj3u9kzJXBRCN1rt0o291KXjftZRycy5uUx1R8i6o/7K2esy
1S6uOEbZqDJT4b1OrGzYUubNsZM+iXNg2rE0gJrdZ+6hxJyilVqJ6Q/0EpjCsvLQcSVPd+eKQnQs
aDds7cLBZ675v2oiKrTmf0eR4O+QW/CVP9F24YvsQ6uPBSxpz/eFYZW/TgA2TSAJQ3ziTol3Eqyf
AprVc9TfjRENuZBScQaglj3FZxLplGbHzFn83ZjTkRmDEgZE6lKWaT7NH5laYREzV8VaYxbVK/cr
9OPe9hNF4VWnPqbALXbsS5ckCMJjwMQW2mdUIueFoJ0wohqEiGNCGdBeHArgAM2Q+cJs+kwopGVu
1ayNUvJIiSWV3oVp4i+xEjw0fp3G3ieOzh2h2cxiiUIfGpqeBttg8MnkoI42PlRX8MYdh+LxlXBZ
8JE+yC2OKcJbmPzQ0IVGb4yrfUqPEJR2vIhDBZvlLzxrMBmPzTTB2bpN5rhwITt3gSKvZ23K+5Aj
GD4CwwLZ/COphba7B7euVksWUEPW6V27siqX3xqpNuMp4Dr7cR9+GLmw6idX9M8e6S0O11X/C9wH
NgrFLGT/a1Y6+y3F1G1A7sDlqqi6qJMcrvjvLCZdIQfFxHRmSBPbTeTQCY3XTeYLNwCUXdABFnz3
fDI0uw+cQHUD9aKLL1R1L5ThrPpuOHZ3mbdyW4AqxiFDBWLGLyz4S7A1GT5apNgYvdR5Qyh+MRTD
FT0EanZJcFPmgnXy+cWhl2vjY+Kr0OYZ2G1dzptGyGBxEaNs/LiX5kUUBxWDnIot+QRyZ2//Ur8M
2YdLfDjO7LSb/oRJwikkfZrtDc73YOQKG+F3L0oOJbuy7HOtQV+LEzuWoHo3vU2bT/5PMKgvf8C/
GQjMhzYLDJaAoNnw6HQc/9K8BFwz2i8mDnWkH5UrQh93Lp3RAMkTnFlJHqMfXXVoxec1FerkHuY0
EbF4gz/Tt+Sms7Gk+quZtbK23YoM6tRPVBYUKw/D89hzV5fYjEZ56x533+TcLtyqUtmwKmZeDAO+
AnhP9hwFmJdi0M0o19UIFgYt1e+BkElighC0cLnD7aFBWCGqfEScR/DwJcy3Xk3zJeUecHagI1PX
iKZ5+zTGmoTWLf8pgVspaL14dGX24ONC+GDRzNc4+XOtRdNOIgQpxXhf9k/rcZFrBmsvyLxEMI9O
b0lgwy0iewUHCMI+wF4KxSVlizkE5z/HLrgNHNW/YQQL7unc86GkZjLQ7DUtJqeK8BlttMy4icIK
6lbG7OyLcVVOJ6e2K5e4Q4JTCFwPd0L1kEUTmnVOoSVqLBALc8olryenqB4+DfOmPqe3lOxOrPtD
Q7VOcMKJoCLTcdHtOSHaTbbN8zFhSFl3SwG6iTm7RH/Z9wZUei79LawWB76qtCKQIjfiNSeN7+C8
d1Q1FA6WIXwWC9fBUmxXjoRzdQlH8ZGUaq29Ps11VtJ8xDTB8Nj3HgnZ6Zt9WeoYzZTn4e6X0cSq
VFNGIclP2EPq+DGlQbD+Qph8jULjfTbxmKWEUAZhyuRqSxhUR5bJGUw5X8hh6rhMTWPk6BqtIZz/
gqHTkXo307orvBkY42BQMnvrOwYrmf98u+WTMNJydLE3rt41P6Vq2++ptTnOJ4JajbZCkCtSQSyd
2mWb5L1ik0JD9fs+aUDghrBY1TDnodH900ci/j+JeiJ6yjt3zMNb1bqNk4BOvL4tUJYyM2YMb9Ii
ABBh5u2R4fmhVW3pfxSNhkWAVNwNylxm6arkaN8dWEI0cURLLBRSjvCg6eGg8dSlVTZTkJ+GZawE
bgx/I1hKRQJ+Veb3fB6pqHGpWiEHObZGjK79xjid/E+VpTQhdbniy9uYjVHDRNjhciGQj+Fqc/oP
dn4YQsIcdS4A9+GU6v9Gy9W2mRo9ZUfijbBl57F/vaAxrTAU1f/B0/vwoga/MwkoyqqlXK1SYFHW
nK8Ofe6/+vtjn7BHzlFloAe2ciU0TKj7R3nKIGCPHq1xCr/1hkRzyQ3ToXMMZloFeHOJSy787wN7
YNqLiE+O4YDiB1wQPNFjWjzZierUI/YyIQ+MB9PGxQdun9Z+cCSuOdYj1WeFi1colV8yKQUGLFko
ORhtlmpQFEXUcNEijM0zn+GXCr4PPWn3f6MaJqIQ61e/QS2NS/TqIcPfwrH1
`protect end_protected

