

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
XoDvqNcsUAMVrCepxGZ+692mBkX+rCE8HMYzKPm5R78cJ+RMc0dkNWWZsdClXOY6y1T5UuLnfOdJ
4pIk+MIfbA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
GQd6VykDj7htiYnOl+4WVHQM4hKgz1J8Md5aI6kr8/Lamm+PnYCv/9ATHhzH1x3ZwU/+Hk75nShM
Z/fTah2o7SNlXBmxO/TZV+Cu1NdyZPM9aMjSfxhjbc4DdKhbt2eR/JXlXgPN+qqN+l8aDRz6dW1r
rhTiAjUos5V3YtoS0kE=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
1H8fvXKZG1QF+UJtGmRK0CnD8bm/+01l6RcgU14qYFFE8GVuJpGQyW5h972p3ANLjy1WRtjYQ4xM
/dkbNa4PXjLXaYaHj221vfSd3lB0MAvfi3uUVJSvclNp9cIhjsynHt6eX7sY3mGpxNDMKipfks7Y
7QsvE6SpbzMkIaxn/W/Og06vrJaRobnXPbk5O8bulSLgRIfqtOFawh2LDbI1+cySFds9EMjhPXGY
R3cSwZrw9voRIz0AJIAvvOBrLoxc5eVp/j0gskNHjRbPo5Gkm/B0oz1Ia6kiZiwtS5XXf5fYsvSq
8ip/JtlfeTs2FRpXweWaPr5rFOg0LxkGg0mLCA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
A7F7hPxr1ObCyOsY3iC3Phcz4OOcedLcCp9ggSn92l+/8vc/8WokvA1XgYsChaRHJl3lXf2X6jfk
OU2I7E3QgZVgyd5+syjWVqouw27C41FFBeCuGD1GtzyBYnFEqdtK4Wi9fPab76EJM+QSrUTFTxOM
vNsxaERzJOCdVgQoGH4=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
DAf8RFZxkL4Com/8UijiDJflLxIdfhDldD1zcH1XeixMo5g8/n+Yg5p6ecx6wthzScLrbvkfxjSo
INrqjZhuOy8JD1hgSySspkuAnlB/pYzsB41QYrTQXDdhODLQLAYA4QNlYnc0Hld5QRA0QsNa7b9I
jitn7EoP2gA5KtAm5w8Y3SJ5GziR/wWC7+Oq7vo7hHrOsipiX4kUa9vhXNaEzGvrcPOJN0YgaqRR
HJt/OxiJdqU+tEWkUefOFMVnQWevf91iZ/Fb0oG88z41wfeJt8eTwCR6ZrUTPInU5uj9Frdns/GT
RmMrsalABVuwLraRXdip/IKnMD1dw9K3eH9MHA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 94464)
`protect data_block
XfzzjwOhx417QodPj92W/R3+LEioFNFKHUN9laYmZJRps6Z5k3cdo86oQlHIoLbxpzznIvcpUQmK
llYhrW2fQBVSktBchtThYNh51/k96CGWjMlrBxF9NOsE5jNbLqtR54PTplfT6+E4Gv2oYZhIsKDm
tU6rmzic4the90bg9FE9Tqdz38ED9g9u74lg0TxSb16rR4cuYpKgRKQoms+DB6RdlZcaOHSXBSgf
a7TbCCm0mE7aUzWsDhl3/AKDodyABenCtDeg2wp9kX5n1osetR8PR9mdgbmN7ZSsO62Jg9wOtpw0
iv+RzNbeQqHJW3SYsOBfgPG8qqLQxpciKZAar4DdEda5hitADmLQyJXNwNCQCsZiaZEeJDovj3OB
Mve1orR3ngBvDjrNJSOoGsp3tDiXRqdwJXuIhITKSc515b8djlgXdvDhAWpDmxcWrX9xcVuOI2Hn
reC1z/aowSNHrvP+tiJU+0JzkmZgn4FjCFmyRdgQ2TyG3hAwdFWfWdWhYZVazmgt9aHW0AFoUmhi
6fEs8TsKlPazbJLhttO8mxpiYR4oihxzWEuBRCRdilL8UfeZCQvJTxFiDWePOIl86orksYD0kKrT
RhS18q1xWgPCcpOi8Nk1KPIqVr7wUH6D5vCKKZ5wgc4YapPeND6BPZxLj/u+RluUZTyq8IzUr7mp
j3O6kE6Lks99nxoCSXZiW1a/s8Erv1pMtq82ZdMR8lmmxphjURixmhSK93LrnCglWQC5XTcZavsn
AdhzZsI2ubTrzGOATJ/fCgrQlDUxUrpsnYgp+90GN2pd3RccQ46mm5WSAqM+J3ek8Xpjlwt7gZBV
WUW9F/HsAmXDMm7Rj46P8X1ARWVk+LdFYtx/QZqn38dWZ3lRblGcyOFU7f+U+oBa26ZT4PNoTNqu
NTtjaNQji7Ilx5bhwkaJ23zNWwZrU7d5arlJ9J1LBF/AYz8Z2/vj8g8gx53OvBoOiRYEnxU4/Afu
TcAwpPU0GV45E2Cln2l3wLO8LsMCfziDvtH1BWw0rbpiWSfbU8pFP/eQ9+/rzuateihMBm4blNqd
9lmLvfd9LF9pE5ig0AX5xl3RPhsF6OV0eFEj35fqIGfyeZOte2TA7jVENiU/wpglWbpuYvJIVn1v
rfSyuIUhIzkqFXavsuvorGbtCDv+dGIgoqkC3cium9qbGBuisi30wm7IG4G4hM2WfDGB0OPbjT/W
Kbcr/QOdr6dWjyOF1bp/nVTBXOo/fYlaQy/kwsle5y6TnOE8I4aQsZ4RYAHUHYCl+53e/lQC3nqI
6kLCzfI/MmQ3zX7nJH6RY/ZNeHEQyykDuo4oJi/SRRYmsoLTiuxOtJZ3XxuR2KRpCvZ6EQThWXlx
F99ayloTiGDpnW37lUIETCODsBpxq8sNCo7vzFMWl1BUtarVT6A41eUPC83sYAFA6bXoCQ4MoZer
ie5dDRJOOaq93GP930KXGmul5m55bzE7NK/uzf8SU6L9L/xkXZQvUNpAt2jas51HCwVrXYSXgoPv
v5wg5uQUz9rzPAvQbb1ApPiIw00dzlMB8HqKEwYlCD7tSdhJ+qe2kMjXQOtGodibgJvpKC7w2Nxe
37Bl9W/kya2Pw4BYgdcYc2cmcU3+WTTQYc5yKM6oI8CLdOnIFbMaOtrBAVaViYUt0YkDo6cN19ud
s6D/7ppGTVUpeUnuaFhl9a8k7NbDU0Z54UYZLiPw716DchFdSLfDhDNscass6BPUCBA7zkB8q6bY
REll4RQdbfmVUCWiku5Dd7oewtk66c6lKOqkpsq9vc5egVK79M9TA8wMeYK7TQPZzLlECoVS2T4f
LKJjxQTu9WOgERPbPmgI2NTqR6DlMJFLAVk31D87a7mODsXjrg0Zboh6ugyfNvYn/UUKA52onIcu
mmryDfc9RNiCodRl5qQSY/UM2FvY9O/JsJZv1m5D6D7azk4QgbEwOGg7FXS2QAYXYmakHHEgCAaW
R+Xralyj2yGmNhqdTPDjLRUuw/YrabRsjjjy5kibz2GmCtKdbCpBVXJYg5oitcehaKYC2JoT9+Qe
HuFbBR5bPobsodeixc/HWkqIFVUYhRx80CL8sIPvB7ocnbNSojUw7Nl4vwwt8q1UiTKXaWPHU5ai
Aj833duVo9imUrMcrH3MOIlSnib4Zi9WMuXFWpsm8/RFYViOGbsUEJb+Yjo9BsfAbsbdHqelD7B5
ymgk2X16pEegbVicQaQlJ7TfVr+JX0z0XHpkJyLPu2uOtOOKLOSPSZP+llhp/a1iULxKbZTYanSG
jkUxpxgxWBtOzEWUHZj0EUoD4cp5fbnSbFnBDy3s4nmKqShUrjuSvyOZzn8JLA4uObhd2b5UDWMl
hxDgJvhEO2cpmxgRD1SkkeQtMVZQUIx7Ed2vaoB4HJOhAI4k3mhDh9sTNonF/ZlCUt+uQ+kn4+Rp
w67Zf8hzUt8tHzkLtWE28Al3dWjaHfi1NwPgkf2p2GecwBps90puhJyJbEFNsdFL68KMtuYBKacC
l+ZYZznrNwzLtJFxcYdNZ7uSpzEo8/RowzhyLeDG8shARZR20hmQah5f5T0I+7a8nLckW7U4qIiG
XiQPmIXaOTmXIFC8zdOPIOcILNlBqCVKQC0VzHChY23850Wa36/NJBKxIQ7S5wIoTK8pD404SzBw
tM/rEzmEdwM4VTOMOGR0zqzNQFkNnyWj1RBgzSzoWPsg/mByLA8MgATmzI8oqv+ETGL73bwiRiTC
ltx+7u4V+sAjyC7QAj16FGi9xU5PYBLfEQ45JtAufK9apKQfQfX6OFKqSj06E3D57wPT3HwipSOl
5AVWuPQ/h9JnUXmRBDziTeTHgjL3TKHIdMV1H8gMlOf97mUPs02+ntIQwuAPZMc7py+XPmJP0rL9
srlcDS8FQrplWnrDHT2u+YDnMuUk9G3WjYb2wCHZBqqg92GDTv2ZZnMiHAp0nfbGvyct1vOrg5N8
8wGzAdyU5ElTux0mmJU2cJKeFyCT91EX/Ineq6+mq5DYV0/9v+nd6ztKAFaRLg7+yPNFplZRl3cY
CLgVC04LvwU/grj6nMDeuSlnJ1HkKfq0wf6OwLZ0EiaskTXWonT/Uztjqs+smM4cfi9a94QhUs+o
NrGB5zm0zhlQaBGjfuREUEK7mf8A7al6ddRP91lUTHq5OUBK6Y5g/qGgpJuJjD3exCdSzNzpQ4HU
d9Jge2IfuQ4jGA/w0J7h0l0KSZ3gg4LQ+UDNeoHDgBGZvcyYIKMREeLl0/s7eC6zPaxKGaNpzQu2
DrxcyYdJ03eJ8O6/RoPiwYrF+d+Z65WuVcgHhOLto7Z8TdI7NLnuV7LDCerUyQd3T4pgDW/MHfk/
75xyk1epvcCYW3hGtBSWc9NV5sx7dbVxqVmqwgG0NeftdUs5wCDZdrityjQKFuLdbpx62yhzUPRn
ZDefcoaOHMFYHlbWyRUm5EJTY7SJSQv/oNSahRV9oYhaRvoJX5NlxxAkrvO3eUecbZuBBf0l9pot
zw8CRF+6k3Yp/SNKbiK5bRlsUIdZRYVKtMRP5PFku+ZkRYZcFaenaz4HYcKtIRMyq2Wad8HQHlqQ
4TUPzJ1ozI64S2RnJ8oupQgg9iGohUuay1j7QoktZ17yw4R47b9Aj38Ecak0RQeDWFDwHtaZ3qrt
qS989MdJMODiqRzMV9ZmxaoBXj7xlL7BofT9mdV8D1/ynPNHaDvhsAtil2YHvzZQV5vgW3P0r46f
MK72lH+PInhB14nzg0BkisdA9PTqMDACZgj/3P4ShT2OB4wAjewRhkI5O6x61AUGOQNyHzJMKKjE
SAcLZaoDimnebNx9UOxEe7keBMXgpqR4P3WXFhOsGmw4jxuCvymO1Ma9ILcqBFcgt/4LjZEHxCAa
6M8wmCqBK0u6ed36LF7pFmz+nLISUFQbVmPbhdJkaaG0zpRqdf4tV3vXOGT6b8Uud2D5WdAgmG1w
l57g3ycgX2jUAZscLux/KyThro4194ATuTi+a4U8fmnFKPYB2atef+4m+hGTpzptIvWm6VBP+2AG
IHlwOb83sJis3utVjTw59Y9u37SByzA2xerhilux7SaZGpver7O9QsQvqCOFeAA5erGgW09+GGvt
O8ZBQ4nx4bNqT+9aA+++vIQGkbzKGRNsSpHII9x2IGSctkg/NYePu/jv9n/JN3KUnOqmaktAPyqz
AznnihnmwBYEkR0SKd0lZnUDnbMTjuRYmat94/H8nCUayy9+HQUfmI/bd9fgBYuFIo4hCl+P9RVk
rAAdANve2OvS/hwoU5Ns7GTGjrjpYMqm7JYCYUlOmfww7j2Imq2bsN+Q4Hid2msnw9nJfZDkLAYP
Qi9wvJRPS2ypiBbKTL744YBJg2ypNxwqZT5GjjYpQysZ0O4e/QwJwGIltZk+KTlQVWN403KdyC+D
nEvKnFu/wv7Qa1PQiA/tnVr8D9ewdU1oO8ZQxSdCfQGUer0d5v/nYw82ZdUb380Rz+mj035tpv42
YkvcEyicZjW+ccWVH0y2f6b/yAshAR6WbKXZvUVOTt35FOSYnNyfANTSNXrA0XFw1SViRcTbMz4b
NOFmM+zJEJBX8L1vPuobTsXtxrVfU9/bf+Ht8gxN94fdH2lqP4qTAHrB7g/mMam70OIpQAjuDpM2
/qe42BgmxaaTw2D5y1gC3DtLIMX8qIPql30TA6RlXvWyUBw+LXvL+ndVn2/GtLRenxZJBEJWQz8M
nFjizJ4EJiwB1CXOhx95QyL9mlLF1qr/rhHX3geKxEw28mSPvtvA3py8ffITCO+p0yPqgGe/j4nf
Z539S9QX/zqfx/8IFAgVNcjtl3+1EGnjKvdFmCW6mkobu8GluxcC33f4kVvrFqk0szfHaz3X+FlF
I1qviDUrHNEo5Sg/DL3y8cz64whSBHfigrJdkBNoEVqJIS89zfgWQOa65iotFzKHz5HXoRztuolB
5MAT9Exn9p+NcyPQRSCaKgUHWX+BSUr/mlldIjbBfky+167+nsOECbpyqAt25d0L5wxjWE6glPdq
JuGxTkmx8N6wBA3bVswsnZv7jgap0ccDtgQv16JYJeuOs7mfbg81vyImrscLZXG1pZ/i2KfWLugZ
WCx/+Yiv2qTHj2CC3ScCIQNVXRfG3aH+1aWhxb0nZ1m1nq0OqORy7frRioIeZVnIMG4MP990tRlR
vHES1T7ev5PMDvY5gdIWDuNvTg57qbpYRc4HWXtE4vwIs++FDWVtC8H6HgK+gI1XiXPJYt0ZrwuU
xd5+8fF3+qMAK5sG806E0QUEDp9fqpafGCJbfN4qNjcZaCmfrr82lnmxOFtzIzkl6BSc6UvR1bKL
3TUSW21SGcOjxtoRGf8Aeu+qEoXX/A3gqInv7oC6XfCHi3tCOaD3Rb0PL7xkpDW0E+C6GOxL3Bkb
Uq/HtMMdj93l5UNZEDRaIABJFTlsoYxqmBx3R8EEpV5V/Ln8IK96FE/n7HSZhqygJKjrdbF8lFdm
vN3myv7wZERhScVz7qFkjh9RyFjrYXYnJ4odeMJfzq8X3K5OSKkUUX9LrMLtw/752xIH86IhAunE
TgvEXUiQsxXpy8zn/cmSaiW7WUrTW8LCmBdTaNh2wDJxKfMYidOYxVeGAyWhWyIA1Rv0J41PAvCW
GJOgfzh/rdClQx6ZkK+HdYtAAwpk9vtI8ZnN3Bia4poDPom/rCrkO1wqXaJJ35tG3GxjMYUFEBXx
0PmGzdveOO8U9WJIsFARwdoDvF4bDk1awik9NpWayoCgn1xKOW0J5P9ZbcwL/YhiomkPTW5OoCjH
swYN5MpVVx2/+SqVcwLehJB4gQEE6LEEF/P9QVkNYLURIEyHzYSBjS2CPxWD4X+ZFa1yDmyNnYkZ
t8ywOh4TxhjrtjgnbHVtgAkjvRAKXe1oWCSRKUGAxL5j6A0x40fFjgLHTrSs/mYAH1jwGnvfpeXL
fJUtAvSPqeKfgtdGpvcegrD7sNyjYszAa4jfJx2vnFPI3ILIO0eE7d3wPTlOylfVfmh6xWnebALR
KEP/hX1fCs/fa/Y0JYE6k5AhplFlhfVaASW7ng1RAhhkRXxoveTVKLkTVa6s+/zRE5uUew02wS1A
wKtI8Q/wlbFZSYX2f0jXoPcO9IYu4818I91uCuK0610wH5NbMoKuf9PPnljCQL1T0zVCrbvZySo1
bqMe4kFNqWG/M+cBzvA/aHhmcWbJGWwaLLjVqg2s8A3xk9MJ5H9BOJr6u8A87rFvO316+vvbBz7A
b0Eb2/NOS/E3cEM/MlrC0PqrGwzx6dQ2XCdkKQGCQik/OzPEfNLTh0hcLFQuaEZ6o4mz2QhnNZrr
KnK4skbKY8xiRrea15t/72yVfBo0+ow+hiftVizkIN1WF71sFdFU8r+6/VOwUdrY9yfWU3jWJpaB
vk51hfWERoEDaXPTXYkHz/6pOvSvlcMNm8w+7iwK56SJMkjyyBQImygjDr+VfwaeFjSlsyBNp61i
gAAA90Eynm6McdjJq3tzfnyLuvkDa1I8Sa8MJiqd9y8QUIjxapfsMluS7eGd1cBtM1pnPOaQTyTP
BsMOSZhImoO9mvZ2NSx89RjS4FAd2HKppRvTsC4GfglPE1tK15usxPdwqIMFaej19FigpKTBvrdL
YPhbAbX2IkpnwmhSpW/JY5ab5MzS80iwO8kUzV52FHAzSqcs1iAtzcXy1MIWakMKj8cBmMhkdZ5v
40/InFSpCKYo8RRJ75w8jkbAT4CBtApc9Wi2Ue/0Wh+/zhz4jATZDq420yRnN2848cJttaa/sytZ
75cZpHc0jeGdBJGR31VsMryo9Eybuoywfl2vvXiQTgkWK59jjrQuin2JmBYHdb+P/KZlC3YbUmUi
dhmxhc44W08kcM9wMinqc/d42Rol8lJN7DM3Q2licFeCBVMWNybcGX655R/3bvfeGaEZkGnTYupx
zLy8qEedIxuN844LlsMCyrAHEPHJe+d8ZNufRVNoSzR8WjrN8wV0wSwqx3AEesz7gDOTnOERuRIY
0d8rmF6Reycwj5IujyeHhebOIBpYjJW9b7LRnvIzJBHF1lFMlozJ2Iu1rZKw2gOEh6s5TkcRCihg
WuTtggz4BNtPTcSp4WKpIiUGZ6+valxgGpxD8AmKZ8TQjlXjbREIAjFxDDpJAt0HqF7V9oFZFt9n
uTHbiNjQld45gGGjzdidv4c32WGDtx3FX1jvAMfMOPcYEujXh9ei0UBNSSs8eEZ1EIa2NR0B8xZF
k8QmDg+dIqbIruLvTdHcJLmQgQlme/4OcNyVcTYOtgIxflSch7djGilI1rwdq3dq3EcmVcLCjQrs
5D3+Pw4IECL2VDvGRpI4Yxfqr7EOrd4mqX8A1S2AExzr3gXLzw3tFUMOSefSI/AEn1VNM1PiFPRg
7Mg81oQh3V8vTFwFvF5ucIGTw7fboDbgSuiWM2ykjTFTTzFMXqjMcfJoiWLprZ5ghK4la+r/wSnL
pepkennvLHypdQNJsPPFAGuXUoV66wk/88ychdzBVOP0RS0icgZ98MYCP8rLys4SbMP/sfEvyx9X
Mnbmuw8/A7AWtyhSj8uEcm2oTWbE3E/sRAt+p78GOe46maTd4Z3ZktVQjI0b/RSeSzi81yVLCFC3
SEXegwVi0mXdBPGsYmpTn/Hm+MXWhgubBjZlPrg/a0hAxxmBRyVxNuiVF9SZwFl0IUP+MqiRNYg5
6G1n2zyc/cQ/V00HYtWab874RwAB31gCbinEecbfw3LjRNRQL5YnG9/QUn5mxrV0bugUvKiW9/WI
/uf7hOsndBkbRbkdLcRkeowN7U+k9zGzlLhhh8TX1/9ePRnkMJao7ue9uZc7KPGNluAheMC+AMOF
oJ7VFApHobLRUycdxzOiB41wwYbmKZS081G6aR9WJHszJekD1T1/Fszgi4pSZKDLsWNJnaozJzi+
7RIXVl05Z5HqtTExe7HVKhe1gUjTzcssXkl5YdEmHHXTGIe/j6iDYVjFAvEiwL9V9BsZi0MoK2Sb
Bguo4WqPobamyGRRuiQ//NiGoyWErXmT2I67cv4CZ32Jy+ZH9b3VtUiVqCOKdGqd2fTN3EDdrYYY
kFeWyDMUccZ1sUuBzyvLmt4y6ZmjvgQI3wrhmL8PDCWyqSLgoJfxlm3ySsh077ItNL5hodiWxx0n
LxkBZU1/TXhomTxmznMsW3aRMk40zj1/lWtGh4IXyN40Wz/5LNbz07it2dIn2Q22B7m2hGk7I7qT
4fwNHyehfePHxPKhat/e0vbPQv1Q6YotOZzTkrImP3Idegnwbhlxgq/3z3fYkHWQYAnkHf5mJwqR
VHkGfQpEUtVN0x4Px5MmGfElFovAITbjw4NPd4VfTJSsRgGHOe1lxT81Jzy8sDwkyT92B+va4/Dl
Mtgl2UbZnLi5m4iVRrV0n1Y4iEYRO8Qm0O8aDj39NdTekJvCFBLAryEdjB4pxYnj46T54JziyXcO
dKlpkyh+mzyWXxiqvs4WsEO5QwfyW3ZEVo8v+krPxM5titGImAM0s1LEjqHhAwnok2ofgANq7vHI
3peZr8QZGc0wbze2P7/bcZESZTagtLt32BsXqrVWgh6YYG4ca/jBbI6xjY1db0eBcXfL53LNozvD
aB+xqVkfftLqc0hVH82shnl8dAAP4cE6OkMGnq7wPx2pai/hfD7Z8G7WbQyoyNLHkWrtmqCdN4Zm
oAjSLw8z8KtdUjeas2vlAiElWlz6suZJQTu7PgnL11oKpG3BCnXvVNkS6a8E+fFxE6TNtxDnGg5e
hHYSAhA81n5k1kBE+AASJLHlCOR0hs6TdXQ8U3AzjZPo5y9MYftucpWxTVeM5nBAs+qo1wK8A/D5
Keitfervl/0Ln37myw2k/ucK45fdVr0ZMav2+C8yHQuvpIresw6OeTPfKSbH0wBpESdfhGqyHO4f
TKBTGrJjiEatbcMkJPcP8OGpT4yVy2OCpFdVchxXYwuct/n9d1xJrVT+HXZrj2wCuPCpOrVUJuy3
T4BPuu00dI5ebr9RgavfYude3+y6TKTytEyWQ4AOwpzUfCFlXjGXwK6vAI7lpHT0OHAFX6hIi0fN
uU3sHD7f7sSBBxvKk6ayW2upfKzLqCoLgmCGvLbt2swalb3XlA2fzJZcsbA0v/AY2dIaup/avly1
8ayS6n2uNFk4PI+kUmTdM6+wGIDJLjX1sfsFYuDQZCMh4Qs6xnPC/ANbMb31yG+mZwfjgQ2ZBlAJ
Rcaxv1BHgNBgSniL2xctSm5Tnjw2bPKHYrGcpnsiZTEmB2SKhQQiBH3P8+oWelLBms/lW28EhtBh
L+Dr6h8XoSLfPOKe0NJ2lYdQQPYQqYHT1cHjd8pMTdxVfBiAJ+eCrXB5h/RqmoPaEMwdHhEYhWDc
//ypU6ueU5BtL/B7mlX9n4J1V1rqkzPDZ0nRwYXzvcWK1kjsSmG79aDzK7FGabng54C9Th1iurWm
BbupkkRQEyXD0J2nfMD8aqDbRRTOG3KyP8r0YiD8xqcgBKOd3sOAxWcmF/SrabC24Qpgtx8Um1EG
Bvfwz9YHX7HP8s48UJvDvBUy126MqTgA/BSnjNC2CuPq+JsfT01+eW2wtf/AKqHrjeZRBmq+GWD8
U6tIGq8k2ObRW6khAoUHIsfk0trbGIKy/RqQFjn5npmNwEsU5Sk8i4wuphqF3eFFzuE9D/u7tKnE
aWLOrlkc/xtD85ash/O0/f6/assccj/TicOpMCbLcTVJ6YymijTIxG66MVC2k/icRXrjcalOPrP3
ck39SANsBd9VX481I9ngERyEoUTJEENAU2psYKyktQd//c7a75fQgFwT2Ci0L6SNQNd8M/9EDumu
zx3ojkPQ0sb9OwAMSvcxkYJ+19NHBw839mkLZc/TDdyZSkSbTscVdLO6JkDyRk7B0GaUzEBGAkZY
91YQKH2aTKctIc1kQY3TRQDDSPjdTQ87ebWaw/2WB8UuowUX16c0QrCGJ2Oq3QqseRmfy69oNdRT
4zvDUdt/sQvcUfDaWLogdMaU7uUxAxoO6tUA11MNHV028Mq02HDZqskezHRjGsgXrwF2++Izb+51
d/DvZINuphup+2J0Gysxf9Vei+x+iMo+JJwpoJPpNWYZa7oiqOSdvb7t8npLOjBBgVqNY8ZKrac5
1E33SPf7QVluE9oJ4dr2V/Wums1BlMZMlD60DXZc+XiXJH8ibg73d3j6kLiYNMTExB/iNFRE+RzI
v93Lz4oAfRsZt2I1tNN0ORUDnS7mpzFHO/eFmY2Wzmk5jUkZX+Zzg2t2NKwFLWnCcn9e0JUld2L7
obsnGwWOm3gfnMD9MmL3xPVg/FMwdC59zBcv4q1NwtS4zAhphK/njj/vZw0B9GC9/Vs0VB9PzVTf
1QkPJwYjBsFdYCR8pI1RmgWDV27PcL9KcoXY1Np4VxksLvLAkNcQIuH+0kYcJWC0zA42vaBQvZm+
o0nnhH9OBpY+3h0049YaVYAPWwkZd8jBDFSuSAZVwLmd747psShVdcdhZnzRd2iGjti0eL8IULay
yskyYqeYv1J5/75dI+7wYr0L5+AlV3yIqlUjjuKf6zvVOwxHkGOb1IlAPzNfcecHrH/Z0tKBgIyH
hpMTqOzuqjtJBmXcX2ZzQXW52qlz7VrMFCpCxP7UxnYAuBmGcW0S92AixlKuGORM4mLU5us8/W8O
x0hVayj1/8XNTEYphKcRbDq6D71iZgJFpJq1cAFJ9jKbZyz3UZoaKWpG0CRhIU18zv0EZvvZkjQk
LwFjwxOXcSTWqwELkKy/bvHQnC7q9Mbv7WvtV8kI06+9dBGc5gAfoF/pP/2CNDsxZPC0rKkrEPgF
FOmdYBVfnGpeRxKX15cTjOIb9fZn2spJZkQbo79AtI7bunib0vS9bn4bjCgdt0f5jQiTshZHFlET
PMjUxZyILVru1rdcq4RuYBl9pcqIBj+VSXjIctENafSUcBCSlZXiuBbMBRn0QV/R1rOlE1oUmf+w
sLXlHdjAQW/Nt2YVSy9eCeV1zrQT9xOhAQhrMkPL//Hl35+KzQaXXxn0CZ3OSLKopVxzXXVCb+jH
qES/VCnmabDqLL7PtsStYsecOeF3ZylotEIF5l3F8LgnBiHZ1XPPwlRyCb2mCpdxYTIXgI1TBNS8
fi+wzdCDvWelcYi5EluiahKuFZ1xxgEuLDLZskkHm0AQyWVArRROzTzOKHdqMuZ+OpXcwS5tiXk1
Aj+Y63jOhY+YgBKWgFAeg2t/LdW7aIflxkHVz2e9pBlnzVrBkL7W3qoc4njKvWDOvmFswgWSP65b
fYIz9cvfkczM2nQXAkN8rCC6wDJjEQ8jYkSuq1KXSkfDip5Cnae0zhdZhL17pMjvaA30bvlmQuqU
L96mGcBIiwF4i0w2By2u0/ssDey+8i+yT9DfZuW0Rqo/Bi9HNh8AlXhIAJKW8VVU2vLYBwYEkUXe
FldgSOZA6IIexkk2LIK3zuUBLyk7DR1oAVcwNp1lpNDdEbQAWJaIssT4RzPZ8pv/iZN/RVQBJwZW
HqRLmobWXbZ6y+EDk/5+EPZEjsk6k2KiNSCgrXKNEGx0h4ukUIXPkvChBf+iLbKJMeyPzry7XFdB
1SVV6iEp+j/XMWXMXvsU0Ag9rugMfPGQQpDUU638a2v9IF6ZvOhVyGOYNR87rxbi10LF9KMvIvIT
hktKtiL9jbcIlxKEL3Q4pcERzoxFQRElmk+4psAJFRciCwAVMnJ8g3V2O9saBbSEtaGF/IKCarMF
HFOjlJqlsIzqEStPG4Q5xT46tvYvnrrSB8FaoN+t7w9kqAnx5JfF7zawQNyGFD0Y9PwSuZqgXhqS
n8Ut1bo7idrh4CTe7cyYmL6VELou72zZXx6pIuo5JkBtG/A1oVpwkuHAInBfAB2jpEnzQ6Y/eT+5
2YofIBVB+EhTa4PVAcNEvP5SdWJkfQNkLcZGn85npTAYODka+ZAe21i+SxXKh+b/x/Fswsacc8Gf
FbkJP4MHLJVykoexXdmILN2lxL1JBvb7kwvZTnRXeibfoWo8j1540ZlBa9VDAD6ZPCaHeSp99/v8
lv9qO7NS0bwtO9ziyKiR+3hpQPtbMYmqWO6wggZgJsGhijrmE4xDD/7JzivGnmw/7W+nEfW3B2oD
xIKXq835QDnAPo3reoEqTpBPpqI7SLt2LCXoNKpNVUJINrc0vnvWeL0qYdRPEY+QX0iSur7Fbnog
zrPUsGU6N0SZflLIYJ9eCIE3SAre556v4CYlR+n6A2TFswcX9JRI+CaeVYg2sOB9NKDxg63swC1T
9Rzjg0g4O5vzV9+yXK93f06n0etlprEe4c8hUk5cnQ4q9tXQOBWYi/KIJMbjuFE0k9bJDrfVv8yr
TYDksJLnj8Hm56+j48W8OPVpYTW8b/c3JdG1zebV2nsRW/P8jhhe+M7wT9EpVuofzWVS9PiukFaM
veexYHkfAe1s93wsQaIC0sTrHfw/PIzZhXgcSpcEC3mlbtofPGpkSi+RM8yzHHv5cnNUwZQK18uR
FbLxkzdjxvMiBrV5yCN5z2c54BQij4K38y66NZemtBf9INyYlpq4p56r/7+9GJ+I3dSSqpknAT3a
a0a32wNAnzAZnJKQhuMgZbyTeDa+uQNMMdENUVlKCaHey5GDonQqdp/McwD59YUiglcLOHwcKbUV
k5p9kwgMciaJEWMoz7XUND2kx9hvC3qcfPplxpKeTFGng75yX5pF/9qbOZpaBqwFKu6kLpkmImr1
X6xUfhqMRqxnbyuQ6cS7r0G7Uw4nOfs6N9fGPsrivBLRdDD3QHZPxBouedqXjwlJGFV1QZkp00HL
blhycHbNGiqfSe8gIGgcjptZgSTaqjFTpMzI59DotbD0Uxd4d9C/VYkYK/NEgipynn0C0xGTqGpK
E/q+AAsts3z4kzX8yrPBgVNEnKt6b4P4TiNk0JRgKA16aVRXWWlBPFkQglCO2BMVuOURTMQFfCsx
/6/5vbcMfRmfXTSDfwEXj/YTyKVwuK4Cq3Xo5eTX9xd/mL06qGMuib8oaJJcQCqCfAsy4IDn1beW
mmdOrZ5X9LCPZb9pyuAgjDk3SHH/cheGWnB1DBIG9pXLYCoA0rjG2zFoa7N9bVMXeUQV5KrTkcxk
GHxVXdI3Ox++QduhcKNF2+dxBuUCZGQeApUmvNxSLmyVE+zx0I0/nEazpYVPmOj7okFrhEfQv8Gq
mt04MCRu1t/06w7zRyN1QeKAFHFLw9Sdv+cHxyi/GSbo6jyY3hDU+cZQc2IlB+y1ebi020+NcfOB
jjeM32EKDDeGVDDuguqsvLZbB599MEDZVQERyx4qR5Qt6oAWqLaI/xtFNRCGDcFsjBLiSJzDrxV9
3JS2cQTHnXmWz08nwz9XjzNrjNnNs8Bqd1Gv+oN2RDXEwY3a1xLWCOW4khAcNCs1i4m7iGipJybQ
BcBzdp8MPQ4A71CAZH79RnJjffVxQlTXaGaEdn7fxYcBt3gLnuJgA4I5f4venhT1kPMN7wyuuBYx
PO2OSS4AyJv+9k39Hq5soGVswDj8JsXRzh+u6HVInsSIU50hFciWSYlHQzG/O2dbGHwlIwNwCv5O
brXbAg/FY9nHxC1EhBDQqGzYLZ8ZEHIyFZx7ExVvcFStdP7/t55HsKpCPp/PGzvWpooNUcw0KC46
t2MgTa2dK8BmNUe0joFAEVTePxqEm4h/84ykkS+21uYHCrf5/A0/SvwA41qGQvGq+YNB3TC5JOLS
11sZVld9DRnOnaN9NBjfuOPnuv1wMCkeUx6Xh+gatyL0PWxM6oCi/m0KS287WDR+oyJ6nqKe0PIw
hiDDO12yt2fhprz0xbmLvliMVNe+0eWSlfjAUQcssfPm7G8HYdI+xcVo8yRmuDioN4LWA9z7o7v1
ouN4QBj5h9o43ysnficEnauSeug1LA9d0LUTEwLdLmS+QRLEN/ZpdRoV5rw+1UWXpi+5juwL56Mn
oQ/i4eFthqaBZO53m5GP99FgJmN74Ao2YGIBh7dbl2cvRb/pOp3xPkArhuIRL40fP+ynGLHl4QXE
3HvZZzNiv3WjTbT2KNeRaV7yrcPxoESDu9hJ8kdbNKFQrTz+CgRyLn2uDLgkx7NCGF2SFzWJh2aB
9ycPV/CtN8RuBM5XStFztNxgYmEMcoCDyJVUB22Wbo2zomVxwjj6TyyhUhrQkzlNx15qn0TUvz3a
xTh3pYeOxl41BUBlfWPOYkHNmAqaE/HAK7FMZebqVO45Iy2KxkJv1puj9Vk6b0jfwMl7ETInKisx
pJTnc8nIvtx7rnfYU2Z0xs+BYi9IjJafjI8dYndG8huC6lVy9EowaRJZgIosJykVtIH6kpzV0Qn5
tNVDtuuVQ4eE1VDxXLuYyh8zDTh2+KsbdVp/VJhB3KQ61+uiCC2E3aLaPziRVtM5HfyOcKfi8c0r
2TQib+HclHCHNN/7WndLEE3zLxlu3T+wM4PuwM4cHhFSHFmp9/eyiuQ/YziCZEU+mSnkhoYqsucp
nPGndJ70484rb/1iFZn5CgUgfC/sNCo3Kae/4fsGmCdxg5+p1vS8RYdAC+s9KZMecscS4SdUCrtv
Pur6Yu1u3HhJiqNB6Rh0AygHpzr1/+/fe2HZf19wLv9tgnGrVJ2YKuaGyyP8DkEYAu/Jex9QoSLX
sLaKOacGfQqxXCPe07nMfycI358W9y3LxcQh0vFWQ2Labuxkq7S/MkJbH4Oj1aEgs0lR7ZkMB2vw
m0jMDl5JZPU/p4NbqtZLoGdiSwrJQ8uqWsUpVNS4CckzuqQMSk4E5zd98FymsAzhJr8eIi9JkNEX
2fJwToWWavJzNoqB8UDd7tTHVsqAMmcW3qL4XN+QGe1EP9bjGGwEmHE2LRjEv7syihc9KK7J12mh
ymPB4JmZgSsS1oGi6F0xWUOF2p/pe10WVwcK9SAn/njMBsZ5IvXtgHIAYOJNzWuZWgFBcUNl9Ajw
wYLt1AARho0HsULtYbA8K2YHAXIIe3S4Xuwvg0hbcax5mfX5yU+TgZvS7VAzz9eRuEMx6HT30g8V
JAD18PMfU09kLeD4Ems07cr98u17m2A51vPvTfPPG1qGnFoyfKul/ZpGuRurCSovQTr9Rcwlu77+
iMbe1RLITVt2CqfEuM4wkTu+ETarTrhxKvsdKy9L9CCQQV22N/MQyzxtdJKYLLJiqE0zNkomEpT/
Jh9cQvDJ6jYiTQg/toagoor9vWxkVx0ejlXRbmbTacJ01q2V4VFx1kRP+6i8/40X5qMrFZ9Bevot
oPziaK8fDcV/n7knXb/QyFA4vcLkd/pc4773a2iMKR8+0/rxaGgCK6BNXVA1VYF9lb+MsoNeysLq
oi5yUNxrpbK44syz/xGDaPeiyA/Ay8rtGE/gEc5t72AOGtlSDhF5IzWU61ngEMWG9FbtHMylypri
fuVAn7VgG4eNQ1azqPd0xO/7n6tp6CSinSiwjGMCDd/69s9gzbM94KWPYl6+I0ecnIPCkp5HN7CH
yYJKZ8iNEn877Y0VPPFbeLyynL5agO2e+U5A6Ysw99OYeGGnpz5mdCqtZEhSakeBOmucwC6wPl2K
JFdO6InNlR0AfYhhdskVwjYjnZbmyXA8mSLvCpRv5yxu8tjlpJNJW9cyutpVCsbDjHt0foMPnD+3
cjH6QYC0puDTvQ9xhLxjgriubsiDswoGtee/WQNQsQV507jU0umPWOVtC2P/LNrRLuSgItE4oeBS
Wi4+xzsjWVr97rsZBUfPAL8CCvwYq21VQY160qf+b9L5ZlNBepkML2jycNQKqhTJD9jUOerZCEBW
0t/EQOt3BqwUw/pdXwCPQqqjBOBvjfgRJJoPX1kLaGk+sPXBrdHHizPNegZ/RrjX3L8ff8HXYAP4
ap7h70oZeUNINbfCyNDG06jBj61gJkaK2mDZj7FRTegT1dttgr8M75c2mkhVj1aRChXgRx/uZo/y
DIwE5uw+CakHfWe8AX5f8eM4THbrfJ+DCMY2VVHRoVbwmXqiB3+CCf6a0vu/C1xJQCyINvpIJHGp
Nrw1Vq56Q4nXnsvrXCWxRawapM8CWXFFjKpksH7t6P83J8AwIr3iRzJ/CGL4ZWmIDYKs6eycM4No
XsdCzxuTWM1QwcFA/DkI6nn8oVSPRDa3SpZKYk3RrInhys2DBfgI4Hc4urnU4OLcd2c1FJ9C8oho
irymP03m5cZRB4/HT33ieV00hnTfZvVdfD4xfLgsCUddQl0MV4VA5ensC5q/9HSLucZH4/splHdo
2PX/+zJAw0no9TxzIpEP5+F2XXn3aEUMODfVHgcgPkJj8ZzNW3uV1xMhl80qdy1Le9BMV4E1lKXq
HU+9rSlR25y47JlHZIndY6lbKddYFVoFt09RhL3JQKgOMfe9er3jvKNWb5wgvz5p4ejEoJspn21C
3U5d81kL15Gr9bJ1DGZ8i0uFBkot2GelTUPpE32AQr0JdtKHO9WtCh8rrktlrKwjXQSGB3LQmnSZ
O5wk2nQxVSkpUBPOaVF1r8NwoThxB+GIr5VCLlFOp0Upxh+zxaKmpI9WsRt2QCH7fPw835eTcVTY
GJ/vXbnT8XnqbpVOSaz994durqhqbxFrnGRoWi8+dKQFVxhyBNTyQAYnQ6ynyncwu1xoCVYnmbm6
Gr4e7vpbY5i7hq2e5kdysxvZ5taQJCZt8/A8domm7ZJrWfuYwv0ViaLamIfygouvkkAz+AcLveWU
mONeOzIkIyM/qQEGt71jfM8MzSn/pnp2M/v9/RpEpths5u64Mf65kIG0haAZfusr5ZbY8PB5d7I0
y9PJsMQ9Q3Wms4kzWbW0EgqkQNSSztXLR8jsrG+GjQUARWjO0vrwinojMY9XpWadcykQT5FOph2M
wUNIGHzHb7B5fNZ0f9l/gFzrYiHqQ3bXGFv3h3ZHQjMSN8u3I7kBSQAYPx18YqD2o83TWxAhvWU9
Cjk5lUVlhOgrkum1F8dH/dRIzWjDajiewg0ufT7WKd36LoxXZrMr0xGErNC7M6S6ypqziGp3GKDz
sER8bKUxyexR6P1tylpM7vnEEvp5HtrHSgdi6H/G3Zpcoy09gQFTWzcw5tqS5Jg+KH9DxZYbi3X5
YXQwTwu6/QURuHWJx5A26QCS0yWuE3ZOoS5Rsp+naZaSS2xWBDRXqKYO2dzORgHp76v6x+wGpJCU
gB6Y1IRblzllQIgdzrQ6qY1imBfzDh17mpLKO2OyauDcnserULHCA5WjyKApK7vGf/9MpMRLnMML
JLmCmH00dIBCD/nv+hcARcru1h0Byf4bXo7hwAB43tI62HqODTET8zO78RBpRxvnmnvs2pMIjMPz
Rpds42d7ltz0PnpTHkfBJG4LO+GwomjwWW+bm2VB/sOtUSW9/AoFpZj1NIl03B8Ic/2sxNiHZfVH
CP0w4OtMdcd18hjIuhyI8B/xS23mb88BQQF8dpi7IxN1G0juIwzfsIvMrXR9Xltf32D74s3intSc
cmr0p6TkkQR8UxR+P/HzjMcnrc6lTl6kHvePXBwrNGJ5D07mvNpvVKTAGR6etZEh5myO6I8ht+o0
IVx4jJzm9pDWNx/wcE9OkgiyEfHp5tGt5eSBYo5qb4N5BeSp+MTgkhFemMGp34vPtPE+wtwl3NqB
Fq1go8Lj5enQr4dud3SDr/WyVYkfHtUTCneZHPEcaeAUJA1vLsmlZojIJ9rarPty1anwvWe2CV+G
QFe4j8/LkYEgOpOvdRp887YJBJ6ibHOMfl6VbJZodEmfsx/arVylEgh21Hl/NIYFhJkJn+ZV7C6L
9p8iTv5pJOPndmQqId9iVZKf7yH2x1IMDk6PKAxx1BIoZRP2F3qo03MiE6R73mhmNK93BzusllkQ
oRICVPADiR1/UQTVDUiE63r30fB6icjX3k+Qg8lqcpoy0fqJlNWNNCbLruzN+ChVitTxIMubQC5o
hcanZv/ykzLEz/hLZCc4viOUEegww6fV3BRU5AJURNSIAKtUeGIWSGrl37hoKoAveTRGzD6wK3dR
fezEdh7+wkMEwZOtxa/zMBx03ch2VVYw2xL/RfhVvK+ZNCj1eTJdOyb8KbpStAfh8MiiN+VFlgpG
6Zqsyhmmvw+sRTqBLUA4IZW4qFNeSz8GiDcUQg/hlJ2MxwXbzs3P32J1fdFBE6U357kj7iiiNk4/
UkOoaNVDQZ7uGzHtUP3x9kL/BRuLC0gPbgQH7KmF5jetlxqIVWpQ8dabl8zdcI8n3/gXhTVdpPKM
9zkb6/8/KV74Dsnn1wDPe93njg+iK5LjP7CyhKV8YaH4UM8xiPIgYXixxOEqZJKEziW3jEkuvKN4
05CRUGXm/HJneb5pCmSmM6tb2xiHvw4i9WTOex+EmUvbYYIYoRvCbkL1gPRiE8gtXhvcnlfHDv5L
qvaJENHXiFm2bnnKxiEwCGOHb6QPOqGedQKRGeJnlrMCQ/gBti6BIiuA0buGJg1FxoAWy+xlvuf0
wkd+qmJBS4XYMm8gXl59U4lOEw/w5c4hw+HLwSIchXisrYi7btQPU/2uTmu2xcMgAEnsm4bCS/mF
z4FRUzT20btgo3IicrVe+ofCYj3DZzywxT+ZfI2R217aq3tg+qYPktVwuRXv6I2W6bkTDktcuXhn
qMbVbI5wq4RuAxA4Uzeo2SzdIpU1Rjxhij5XmFV3aw8/ycVMGDzH/DyiOri7wQNj3PKujG3+Q/nE
FPaKixj5QrXuIuY4E5RV2mOWu9Xh2mZXU+MPKdc8iISyESW5xCASpgJmqo83K7CaDsehjCKltdhk
ItBYgu19Qj78TGYMHSN4iBUqDBp0XfgMwzSrCS8/hGMDbPJd2t1HDU7CipvPIll3XW9h2y+hSmyd
+16kZU8MhNhGq5HB2PdxrnDZ7sJIWE7iwZ50A7Orw0Uj3M1CO4POxaXVJ3fQALhDERne/6uvEKfR
vjOOhqRgszXoXn5sfRsiUFrIisRoSZRKIVEOC9E56MiK0wPJHsC/G9c0YOsSYh4u8slVjKKgTqnR
XL+sWKV4Ir9XBWgBMKpnK1dn7x+YdWOSmOkTbcS/dulwnrQFRj+w4aBjmzGpUoSQfJUpX6fYKivV
TS2rNWSyBsts5aOLYoCX7gv9zg550JA5E35uAUuxR80Z+IJWKVP5IW7SIZTpJkN78P8fJWlimIiu
dBtWV7hP/6IAoH0X+imDf7RCQIyrCvGASZIZafhZbBhex83FBifmET9fpKG+1XI4fqeQzRhBCGK9
gmVuLN5MALVPSXs+rR8oI8l+0pUi5xwNx2ywfAcqVu/UU3vsbeVe3JX9LcmDaYWmh5GVUTMvNENL
3UJ3yzb9LodOmGiV77wAHGWY07Z03c4P24JroeuFUymwCsO5nbcbvyO9Ke0zNjaKitUNOFVu2V+p
w4eLxlyEXZ3WrCnD1+lI9sncBIMMpR96nw15jjVRzL3ozQa99XRKDqrVSQwbptwqMK8aWERyKaic
ISOl5eXlnp+SUQT8hVkWYT3iDm0+OhbA0rrXpdk3Inwv5JaYApnUodBQGHjwpU2NPPn91PXKwuaR
LI1MYOE8A3rOTROG3UcYq53srgowm8pTpf32Y6eb0j9w3K5/NBRwtAGKQ+S2r4fJKtzIist6hmHB
xeAERTeeMiP6mgnqQU4xrzRj5ylwT9JHzkvRNkChwQ9q8Z0OOhzp8Cf9NcpdjBtpBdAHnO0we+sB
cfUiDnfxC3to2VG/+qURCbrdT3IAjD2SsButVG4GuU1mjdVLjGbtT9wu7mE8yBoyZxge1k1++MvF
s32Ksi2gifwo1Bt+Tmo0hOuMOmbk30jNN7p07s+fdctG38tl1OVIKgzbrs6o6A1Cb3DlsxqXgvn4
dYoBGGxcFm21NfjDPsSseTTH3iP3zVijkzhC2U7lbHCpNjydwN+tX8/r0bFNbX3aLPgQ9DK8NQY8
XEXKWK1As6K0TGm1AHYcRosIzRGELtxhdxTF/vSHByg13S/iuqDLiNEu+LomaMrSHSMULz7rPllO
Qb9RCji8QnW4QPUgNAyXTt4rKfq4CVD9Pn9OB8Oew4ECzhkxqhvzO8PUz1OQZza0mdIgjxF3ma20
JQ0l6sTArhbHR9Ufjp+0Eg4Ne4c2PRv7p6eGMqIai40PhvHgnjk5QZiiZU2/kQ59lP3bf1gAkg1P
YMoZPZoueMrMh66T7Z0bpGKLzjg/yvasSQXzhPw3j8o6j0SHbyPNOfdk2Xo/Y3mOLuzBNEeOWzYh
cpvJxDeR7eqkiHF+QumSPWKOhXlFPPqqEHrdmEGBtMmJih3ddHuPAXnIPDudjv1NEbGhJJfYt16s
kRsjigqrj/ldxmOKRBk7IeP+H5bCjFwREMDzBE8cl9/QgODy9YLf7tmE3mESdjd7sRjdpZcEtMqa
3ncFfp/XJctJLwP9EmZjanvW79TShjseGRm/P77KOsCEkFjI+cEFNzkAPB8pLGXwQAmyqrAQrIRE
cni0539/4kVfCQxRC/IXgpFqD+M+mvehHQkYPjw3K0tNhwN6R1mb3wLtu3hcuJ0Lp20tp86aykwC
KEJLcu72WQcnJqFCouqW8B/aowpfplsLzGMqf63h/LfCEtnDyDCLs6vGmEx+7K4W4nbmmkVKayLJ
7ajkf8fCw//pQlgrfULOTdIkPi8G5O2bFJmff714YglqIrpPS/yyW5ToxsSXDnTF4Uo5/ofZu6m9
gdKFM0YpH3kiOGQc7YjET/xzKbQNkdI10z2wrGKtlSh6WbWmGr0a0pH06VbeiTOAtn6VoWE/+lLe
BMjjyHVj9mCzaj5WmEzhj6MLblzJ+oTK0vswhsFBlSIDzvIueMXHWOf83qjkt50oRdKVWiqAhYyF
2WNlJr74BhPwq7qHup23fiRhufZF3JK/lSJDAP3EhpJXyYwXjjmb43+Q7mUYtryConxzgfGvKLNs
YgXa6q4YilsUO0oEUxI9Q09Lze+8F4ZWN1l/rK9zYd7o5XHEjmlqh8OcnxogkWTXbx650vVUnVMW
MM/D87bdDkT3/Lvfhc2bZdGRZ/Djbd/T7umUl0OBaaw9GLo4fMMPCzkgFyZbZ57DL+lk3rWQhMMi
WlP9C84Faluu38EaMrzWsIim5fQ6SEggvx74GuBQp8TfCAKC6Ffb7X+L6CgPUAGGpKORU4Tn3G4T
sU34DCLx0YOWw2qe4j/YvK1+vWv3zDcc8nnLmOC9zQVkRyNmV91fwoi4aO9nCt512zgsPMyHzfbT
XD0Mq4XUQ1Q1yIEnqVqix6ON7W2UZemYgKXhxXcYaOrPavdfX9n4svtA9lm/SyumjFXvkF1BMDQd
5MB+BZvE2yUzJbRNKnfaN6kNxECtJEx712cl8vBF7ttXz3OJRkZBz99Uj/3B8fQYvp6JA9fGZvIp
go9+ByAYYoCoWXizUSJT5m+NCHBhjQ51RRgqitUPMZ6/Y2F051WuHZO0eN11QqVfh0q7YulBdlRm
NiiRVtPI5ZaTYXxIwWzEoj+BCIsFbmHmLxnBhHrJTIXFu7vlqaBB1KZY3GEJM0fBWev+085q9ds2
rK+zyoj1s1Z5QQyfZEG1Jv0VdZfvrgQXe9bng+XZEyeMcnUCS6Qu1HZtxi16S982gwF/pcX5zwLZ
8yWn355zk2UNc5z4sGV4S1pBkWkVtxFZKGhRt/768NOHRf8wMTNdi2rL4dZ8tICqYPL3jy/sBzA8
Ud8sBBlxiqWpghw3ci3RfGMX2U4R6gqcmB6Vtb4UHsiN7US0ZkZlTjNG9Q2xdUDPAcLBlYIVARzw
ohumssq6wabN2TfZDGV2L2kV9DLueKjxdUn6s3N0NrwWeoPVKc13xdvw6n7PS/qW4HHQ9ScUXoGx
R9oe50ui7SenjSGFXUE8JCLO+dc4ajAhZfWmCtMKiAA0rdIvkji1FATUqlYK+Pex8BIImF8vpyJL
5jJMTVwdaPGFFHVq1GSsGw4QUGc9+468NL+XmU6/WCaZQ+1V4hB6II8G8lurJtzo7rlHjlcuOJtq
PWICCAO3a3pMyk+2Y7NYERlBzDN/NhLED42J0LuozM7F1IvYAOWtgJGPSYnfUQEfrX5esbZSoQ88
pOprdeISYel6IeAVmiyxwVsR/SssKWkFmuAE1Z/z7PEaZ4SKCI0RZ2TXsevjHFgAu8GlyP4D1Kh9
f0ObtsfKCfjQjrZjX57vDwbEOJVSOI6sbl2T2W1UmudT8ZNymjmIvsM92Fx5Z+FTOfS4cb+C8B+D
GdcPkelaT8oBfsRRT85T1NHgF5rGjRmJLhFsw12mMryWo6S5Ot/85HMkVf8Az+6ag3WNflLhPf6p
+CweShDKwmACeaplnEN5wcVs2OMSn8Fq4Y/qEVy2T1fy/F0ppxtkaVoRtFZlCoZaAGGBQcBApB6r
MjucqKVMRiN2/dlVNSgbY3IHqZdeEBLp85N5PJ485qQSTHl9HFWxOMHxhQvVM1LvF1H+OgTWhTHj
JE1hr5zpiDfccpYbEx60eoNPtr+oafekyXOLyEFaCNnMfrb0hjPPi2HpKn05ucBuMpvnJUrAIUtx
9A2M7zL5NGqw1m3NC2In4GRdOwKrwHRLXYJ2H3N5/hb8rDde3W7dwElV69HO4KgPtlHfGuNqKJh4
GH71NDhOwDFnAxv+jkAGtjFJ/c2gSTX9rhe6H3Bw6TNOPGhj8jZcnliIISOtlQZdtIPbThAyP1Sy
WM/lDv5cFB3dMaxp8pR+w8vhrzvQ+2zHOcLhi0HyhwGJC75X09t082VB2GZtx0r9OorRSjT8SkT2
NqQlT+mQ3NAG9MtUy4urnKQUx/fAFoVW25MQwFIXJB35QimMYZ1NuuiazObCZbYX8DAut2qKEhTF
b5bhDcgOcb41NSwF5nkOIeqZEVZIceVBb7pz6Fzj/Pze6L+mrW/KKuFsDN507Z1Pz/PIW6o9H2C8
43VylBWnjxWNPn+Riw8+px3IbFYiqlJozGfsBLT+g60duzBbP8kULUz8im0GuNPLc2rgP3PkI2ER
W2tT0h4FFnN9Z3m8CKZAIm5Jz7Sn2lEorceZBPBNrqKNQBd9fYoiyJSnpxOjxA1j3Q9BDk+c1hYn
Rf/tR6KYP3WcYx6LYYxo7+cb7+O++QnN+mQFjr3Fe9LY3C3R98q3a4rkXt8N1Q5AFuKHul6PT0c2
T+71OyxOAmrnBjyHMvGwhvTbpb2NYFTa1FVqAbkkrPSnra6eDVoDDO9M7pYg5KyF+od77shd/6A7
hIpgnVwILp0fAFixJi63JCRGV+MxTPI2yqNNqksX6RAqaTh1ZyNbASNgNleu26Juiakjv7iLz2QP
rj8GnKLS54/vU8FKno4GXw2pMAe7xeXEUbJPedFtDjunzitHdZKY/XAsO1dSGpvb/rV+qQDJ3IRS
yuw0K68/zdjhaltvmFu5lXPfZ9svDzO6UGk2YhtB/GR4IY8VQ6+hHVnQDyvomURo+/ZJaD6CGx2n
xoxS7gpYUsrZqu68/KcLNXi8fPsdfTDlJuEpXx0MZNHmvglBeFF2E3rGFGzB1JkJulneR2MCLN2s
ssFFpUa54SGyleaNnby6JRDmgnrqu7utRZWhW4T9Oq3Xdbqp7CqPaVZ9PmGoY5WOsIk8OW2ZvmmT
czLL6ShDT8AnxctLrL7zVS//k49A1YHmhiRbalj/z980SynAJcOwUX9Cc0i8FKZ+VGvuu4FBNNz9
bDqyXDlzjhzuyTF2B7Q4iByKKxsvII9HUnI8lVw1enVCVf7wrItmVnW7M4bwsNM3CS0Buz41bUTN
ubIsmMHTqGSsRO4cpbH05+653IRjvrfOOf5EDEMYBWWCuDYbJZBj4zfYOVlgzqBC4StmadHJ88rN
10yPe/OGjylxEPcccjRW+3xCafbNSjar8UAqRSSS5fwJ6LhZb4b0m0UysY8puVhH+ibvsXZusmMK
18Ert/KdFD8qpYYdQPmUUWQs6YOpAmWOvQv8l0xmy3MxMiem7hrZozZntMqD6ZL9Vz/z8o1qB+xI
bNp9ij2eOD+HxEnCD0p1yZ3SfLwYvJZsCbAnvmdpQGQlU/l/PVYt8vyC6lcVhfS+E7FvweCETDSo
BeBJFEMMHRsNyewf8g/JEO7JnDUlqTvFFhdxtoRpwzcU+8dXrgJIxsF7ICvklPoTYtHqrlshzSf4
kutZAj1iqmHiRUTjS4SMmRL9nIZoTKat/RM8wIu2KXYNnVKW3aOaheZDihTfc/TJYGxKwuxX/9le
6y6X8yJu5XcH3wGnFZOY2hug0X6A9c+UP3nGjr9nwedg+/9iDIDJrAtHaFRMbmTx+i3ZknIPLdhH
av5x04jm2ezZIjGopvxaichOnG3HqwdZeSoq2TwuXMFmhozIgo8AQR2Zh4nZ111GC5tcYUl5H5JN
DKWoocRYBisdACNA6Gax+xRvD8cEF1BnTNLQRoQxApH3VY9D3vESNO4zjsonrnUT9KtVADE9Pdgu
QbFd6oKsuUez58jMBjzmXzuTTHM8TkyvBtBCUog7JjjC/HU6PZvNmLPq+XiWpg6iFDsJEvDydrgj
u8Fae40sAQY4wIWeNxpkbill4OT80sUqNTbKr7i+Zg0NKLwhOBjTWoZ+gOr5qr+eO5UeuQsoBIRV
Ni2tKBE4+9tOyhGdANl4U4fU7gZGzXzY0ZRrGUTlQg6260kLAFA7TFno3mcBX4ASUgwRmFcTukXx
xj5WDZWW+3CVtTeOGNKWLWOg1ks9Ap3G7T9ayy+d2Md4ap1dVPYR63/5/NUu62WgdrDSYnszZMDw
/tWQ5UYP+3HWhB4rRis/HJ8F/1B+/Q0xAY9c2rjJs0gRqHT4ur2DCzVQw96ZHddnQWrKe/OlKIEZ
DZaJhZf5C1/chVOphdGUFn1AYUXeZwG3Skh1BIqq/eO8cTBm0jlJTrL2biA7zGvlXMKcg33e5hCW
9pFQdjdPCV8isURQWywj/gvOainmVMCxSO6z3yjB6tlkQkPQl1JQjiDIuEvpngfySnRp9dq1CtkL
MeRb2TJLiZEVYSgmkUwxlgSWzQtiniH8YZp93wOD6gSCiLmLxzoJ9YQU/x0gpru0jN81GQlM+aWq
L+5mO8t3Fxeh3ucwPJ5daCIN6uwIlQduOFk0/lN79yzj8hjh5Lq8onfhoeUpkinbGOpm/sT2TVU3
zqwfz3UtvttyfuO1wuGGWhKzVOJIfXeLUwQFNeEvfgOrkPTpu2+8kfSCcCTRSFSMGusWfortajRn
9/rJSZcWEJKgSQx6nE6Czq5kwWyCkNQ7edu9WK3VCEb3Wzr6gcdSeaWLBH0WNOsj6W9hsqcSKrea
o/ayNOqo3mpGOsSFtIlhec9FeofGyTtLC+irj0nAXp6+upaLLD1HzzV7PrUajlFYF1Wc6a3EE0xw
k3b7Z0crQ+vEmLBTsn6BByCJRHEv+00vrToRrLV6piPZK1d7M3YY+3YJvZwh7iQEyrQp17cB46LG
eOiC2xBAdB+nd684VyyOFxtTediodywkRmp5RHw4BpDi0khdNnxsqnX5hgjw52hUDLqKL/VMeJOh
Lzlss5skR6/OteTnGZshT/v0ZHANOE7OnSG6xCLloimHesVcQKbe+YJ9S4TOm+AcP2U48r04vB4k
6nZsC6Hk8phU58nw+OBypQAIrw9iimg3IC5+u2bt3f0oati+hbiCKL7CPL5dF9qVsFrIwbT0Bo4d
Xxmg0sMQH8raM6r3tPgO9sG622rJlHPUMa3xMFnX3j67jZH07y+uFN/ve0lJDS6BHWiPXTbIwQw7
oGtjerIXm3pekqbeBCLGNscQdwKegEz8KjJ5JtyXlpwbCLe9Od9XIHtJde5OKh8zOy19fQ0eOVKd
zsFG1udSSR+h2ypG2Q15hbd0NWoKbIK/UOJKxjLvBeSr849Dr88ZL6u3QU3QQ8541X4/Srn/BRFz
e2KSuk6jA4hysAng+9mU8IOGMpHJ/oAXGpUE47Mo3JajhqXiKl8Tl7C3cU364rqXZTuOgEPGHLAJ
mQVxC2Y6tB84HcAMY9UYzYMZ6ZVOYOeo/23BSlPyiSbj5iJFVPhmTmC1OIIpyzUZV6QBou37v3nA
nhIAa+BwqylQABR3oMmZpqeMaX66Y2oa4lw/ZpePLbvUqNUZ/h6yQcI5xLuyxlEIZEy1veLVfTZm
9sHQ9vbiEPqsaI8QnvYeEtmE5RijR84Of30ignv/plzaXGQyRVL2psIUQ0j2/tDISut//w1X06IE
koRv7GkOm8irJwXFh5kuGop6AzFvtOlQJZvbSLDVFzJskdr/ku5eGbQ2umH8aBQLYrWZfsyyUJpl
c4+acR/KwzwG6mc1gkz8kXQ0AbkoLfTTBdF8UQ7zP04FeefPocjH3+vCamkg4HsdJ9TSsPqZtLlt
f+NmPTXBo710VzxVmD4OO8ez6Sab5MTYtdWI47cZQYMc35ejy42ywB/59Jm00LgG4zvpeyVEI22A
igAemZOzsRbMWoF3sf5tAGA9alTyXk2/SmZHY+VcZgw7kjGLGahPMLRnUCClLCoZkg2ms9NHDQHn
dAl0+QXBh9Z1jaAPdMkuIP5r3qDHKdeVcylkGNamlzKml3OO0WBNTWrwEtYVqrWt8Iviiz6vnGkf
gL6B1HzYBYekkcIBSs4dV7XU7HFtbH51588q4J0+EAJ/C/c3o1WsJpm07FrVxzd5aDYH+r/Uojtm
NL63GTDIuHfiyrKA2cxDXMMOUhFTzfFH3UAHBQo8y9S22CJ6013sku7kKGkANiXvSm157mZpe95y
nkn+5fGNy5DVpqsX9fnvNgKNq704dDYPFq8U0iElHYb+HZSDVKQhJ4xCiysRoYI14PQBCqwDD3UL
KM9eXKTnP3lYfON31m8lsvHcvzkS0MX2MmDOZZfuFFsBsvvARioF/fEAfuak6H/kvU7ZycY2Di3r
4m2tmiBToRW2ztErFphanUEGonffBXRz/vtqqGui4m+gADoP+xQ3zPrDM2HtvEWN5Twa72wzLf/O
0Zi34l0gvO1ClDKR3GTgZZn8VnB5913WSYe1vvctpMHJ/xfdYpiF4JxzLNVZ4zFIdaFBXyp+GOi7
PYjaNin+KTvpCblmc8qjjNOVs02JSKj9YTBRul6yy+s1AK7AbP2Qzih4tFcUS+LNM2j4KBzI0mK1
EYRGtKgQ/CGl7zm+sSKzIB3O3vJ6KILjMzE1iZwEoeK+cbBmLmTphxquSlLdqY3zOM/twnn2j6FD
HN7Pa07qdpGqGlmUfcpm72ZuvXqCIUUo2no1c24fsi39bUt9QQLkGKj4mpX2zi5ZRB7LeVUYEtsE
8ExlGcddYLJLeSeTJT85k1DYkn5RuR2zcMMI+4hZ1BEHXZUI5vwj9OBCIYYKw6yYkSWqfomc8fU+
6DSN4G/c8+oRgi1F4GWqSVONQAULlWKUa4UZE2A9ukcUnrACEKbCnCzSCuv9H78eyu+FbxyZrDUu
YN0de5E3qe8nBlLHPhl1Tlv0XJO5WGK23GxoBC/LqpQDv1m2bxJHKz76IfitaHUFug/6j6F2FD5p
YFEFZNLQjKW4jjwah6CcMmqBRfdUMfWgDtUzbkO46SPNt8CLxWabYYuWGYyZCIhwZqVxnmqYcVE2
rJTP9iRAa3XAqP1NrIdUoXN9nWiZ7VaoMhtCtX+9pezZCJRZv/KIBQ1rYphS0LV3ENmDnFRMpfb4
DmeC5gi8QhcSeP+Jja7kLIrLsxJSz00KFY6rRf6QmX3WI2MlD3KG0yEmWU6qH5rOuQDx4Gd5azJP
X/tdhyppO/oPx9qyD666nzkDSQ+25MXP7z2Co4DIevfjwdLusVlI71brTpsU75w4GccO0TOx+wBT
59MH6KVVp4A6joxbj4T5/7+0PWwFs2s8O0GK3Q7YX3XfJNg48Dz3hhBLCiyPM4cAMuRV2jg99lX4
Mi9797FhGGbJZl3XykKf+4KfGJi/O7EkDbtABE6uENL2BlyiDNzQqQ1X7/ehUB3dlMqqT9LNsE6j
5KeJpKR5bUp0R8sKpDUT73ptTjRwRkMEJf8kjTmSg4l9/4UgblIq7CyG0KqWS9r226451QYVUC7N
KeOsza1IYARz4/il8i2lEv6WqdIYoVO3e7YiKG9q535mY/khQhvGa5mRzXs8vMFSsz8fd6KAJwhf
llxCthhisoU26hvrx4+jA17Y+sbw8mRSjoEd04ZOqFHCbHkfCs0XnRKxFWYTOerpnw8zueTkJGob
de+wOkJt/zLGPFEouPbX8gZA0wJGAczdvJ++j4+OtXAGEmQFvkKKKap/VNaxiFGI3lGtBAgUCVYq
AUi6jjoWuffz0WeT4R6Ug0ZBNWBUZaDmBiINXQmoQJbL1CrVPJyy2qA86o2wKpv9m39DdurS5GY5
2g4rFDgycPN/5HKVR7OANMphiAnmUkKJCdjqScWiU6bp+pKLCF+F3VxypDODP1MkMYs1lOougo9E
mPMrxMorVNihBYthX4kWC+wcKlnOuhEfuwU405X6p2rCNICgz8gc41kMGo2D/m5/G1kRpTZFXNuJ
fXL29Fy01esnkJxspWXjwdaSWRg9Gn2yqXxH1ntNVh14H8siM4iYbaJHTd3FlqAH68YwwDWGCxSV
Y2BncCIhNSNmK8HeJ3LkfUSIbUJjLHoFG/WrpXWhzb07q53BhDjZKZgUedCQ7d5uiOtVBPQQNE81
fxLQF+VIPhGipkWFifeY4VmZFeMn72/2irpMyeyRbNTH3+h38tPdHUgQLlNVHES84vPF9XIzqeHW
eZRQ4U2wN+o4D3tcihwsBM4Noxbv81wwCmyAZUp4YUlPUF9inbhMzQLfq/pbviZIAgvCPiKzlr/e
IucGzEVUrA2rdA/+FTzGwI7sWAUHy79EgiMGnRP4KwFGTGqnGVO2HTkps9l8/B1iH5OyXQkIsZV9
M1rvFBxUhkKFqtM7BfH3NYk7UDxZjEoWpq98wJ5d7abAjTv3fLD//Rhq9wKKGYbxs3PpozOpnpmi
OMQF4vMwwHM3x5NixTJcu4jbM1Um9gVQxAcuuu30HrYqJ2AkCxIehTG1AawaXaRCwZv9Ue7pd0RY
L2JUF0yyZLl/FsclzHvRxI/eV+3aBxpN4HGOQOl/RmBEjWllHkc7YIrxQ6gleWOsW8epD/pk7wUz
QIHD2aE8fe8Sg0wycPnkExXgxp4pBijQiv9rM1MvRRTAS1H3CrIc8MX0q0DWTRUwTdwxeFzRdVBq
ppEysjwOgWOGJ+J325Q3/mIzRNi/5M3tsyMvpizo3kDCQNvsqT+yu8DN15PzOWEnCGIdHXCEhBZZ
AAt1D83qAmOdYoOQ6V8XbObV7SWd2PtTek+BhR3FlGI8rj4kYATu9nANk+zZTFlgpFN+C4ZfQXuZ
1KydRfuKR5xaj0b13lU8/6BWzztcOD/4QyY0Zv2YITs1uIMK7X0yM4EruzPAVNy4D+rR1SxIk6rz
iueeHVytNwmZqQ/3M47p8RMklMTm6mjKV2GPw4xi5CPICC5mApJT3U2E2gLskqJNJUHxeudLJQkm
3fA8YoueDGJLU+5ejIrnqq/NhJKpwtCTnU3kku+pfmKHLG/x9NoHq5o6+4XtyOstDJH4Q4anbxEH
6lq+Coihm/AiPn4NmBb3qiXExdQYQHA1EDGOCBT27rQ4H2nYQtVdiI5hOGi2zdgaTDVtBZKM9pzB
8p8dv1rR+yiKk7OWmAeSRHx5VVZlRk+tEUw+1tizz/l6vYXlmAq0jUgrHNx+HsXC3ScGRPvVBbHE
Vu8ziAGl8lzs5XhbwkEbcN1QYp6QQ7OTy7xieftHyOd3Yn9prJL48P2TqGqg4tOAtHLI+cp9AGi0
PnbXVlxD0/ZkPaIhmKUAcbrDspA+sXCrf9bRPLyiCMRfZnRoxSLYdNkqkzk1sS1QG3OcxowdYKqr
664tbCb77LzcW2DHAQ9LReEhm7aO7AfjxabZ8FCHa9itwTLQG3FV4xmgF5kq7CEt75OGHLL6Q8Fc
1raQJBy3t/bod3JKT+9SVRTwxF5J5VDaTZZG4ckG5Fdyo0DNXUM5yeBOHticWl9dz7m5V0/bzdZ/
crc7UNk+OezWClPTLWc0+3gK+injoa7IuJplEEhFLRnmcnE+YQNdCl7mDiMFLVjXJwZ0lQr8EeNl
nmJ/J3Hh2ZzDAvuwipSagoOZCmjU5afALgIQoXUT3H6vFBTDk4YdtjqJ4SOCB2vSIlLPxJmRwpcF
WFmWbA9qSYg2WQigoc7gGJdIo6kpAxfpfPJSuVF6yOS1zb8azZbfPVlZO0ou33N4e1gvTGuTdcxu
+tsYNAfXeffr5DPRY3XVTnb0+AB0p7+6X115NDKO01JRU7FFfpZfBqT4XuI8A+opCMyGaDXZBrEd
wWalI7BG7/Hq7i1p8gy1MImeQNYCAqzCXlWdwBVb6xAujgyOCreAYR8j22KYKFoXqIyy8FACvP49
iXEUbEAoouxgPSoRY8EkLWBytf25kxs8tGW8PpIIiU+Xdc1kDLulcjJLdjQ1I4Gn7+g1razkuJIQ
Pn3go0lK57uLRiG0HJcCrrELysxLAY9tahfshMCHDLwceauYrDluB6i+qw/e4RYaJAuB3bOL0Tw1
LDbLMZhyuqGeNdeQ5CzY3G9+ZNgUyOz8dW9AYNZLN6PEnfhFR4mqWxx1RZnX3vbECh+KhdvMIiiH
lROkLv+b+vdcIBaFbr8w2nUYg+FNk60Xm9klAYl34UC98hVM0JUYls68Uaqr5i/Oxx4pgkfADmX5
5hq+DJDCzcRsVkep3JbC1hd1cDIjNVc/XW0NuOM1Ehp/mEZTvNxa4tJkcHugeDhlyAMg4r0O2BbZ
/HsU1wcVdjvUENXSkGCEx1SKlikGnxlyfvKPE3AwpC4sRI6TqS2kEyxzk46cIX+q6P6HGACW0llT
LMoWH2kLS1wp+pFIdwnDP3IVk6gR22oEauISFOtBnrbB7KUq2Lq5mO56LzQsxJuTpF4uK+x7T1YC
ff/tXdDc3gBtsYTeTC7MOwlMOiZNztgn5CWyvuQRuQlYAksh5SxJFOZDG8+GzOQHhKMcedxggD77
AC4yTBskUsdwT+WDhvL0GpPiqGZQPmBjrnjMO6+0uT7vSO9UMi62J1fy/HunkHmpEKsbnu3HY4Pd
ToHunuAJ29wryVHs8whFwJLbSdSBmgQerPjY5v6TtrIEZK8JbjNHDa3ijkZg6j0Z6E9LVAIiSMis
l6c1RVRYTF+Ep4oHgs7ln1Vw0PLlkpMPWRdkJ/N0kHdNNYEaUuRfCNRsVpaN/e7aphSJiCKyBZiW
Nsw2yBY2VYSLNnxq2HgInrgNsDg9WvG02dnh4B3ofd4Qb/xouGUBxegr0Hl7fYcTmGRshJLVwU9f
9qRnLzv2R+qeQX626JF48fXgggpUFT3fgexkWDr1YxZRlXoMq9sgrOMxvJkZUPamVj2tkwvCW9qP
cjWX81eoXBTsruY0BEnc3lSriIhInD8sZmV1hwND/nkDdKfXGvMYTelpYNMqsgOUEKmvn5kisuHG
p/aMPE24tkIJjb3AFaLkY5w6FpY4/h5RMkkjdcq2bQhI16E3wp4/W7N0VRh+ouosUU4QAK7hXmgm
L2wwYlEGHehrjwbm+Q3MS2Sqf0hXf4+5lvQJW9rs+C945i3DwsFY2XPjC5QPEFBMMO05u5SCCE/I
aaKf7AliDegf5SsFavCsT7Wcej29TNehfim5P9OzG8DoUeoi5mIt7D3BO6pX22uWjFphOWr+LrCx
FxGMqAHKMquZRIMXm7O4SBmVJl4b/6DguGo/2hj4Sr1awXvjRS1MSRdYo5HT4A+hd2kzYD8pfk55
c16WEv5uRDTHztTS28q7Ljp4E6FELcuhlezegqUaMyMsqCsjrijDkZavv2r84t+GoJzOuF1jxnXl
wuL/wyg5QQDyx2GLpaUGcqPeI2AaATtf7d7RVJGZaYhJaBq6+q7fK5H4cFp/6LapoTBN/pm2VxZI
Qi/r2Q2Mkqf7GodKE215ncE1VwS7mtUxcTZEcvTCEA0tSehq5VnPFAo/4XUACNVysHcmlCVs0bQW
wJZKSRZdVWAjsJAZCKYX/pRmvjYpgsXT5PPUgBPagMgbmL00KFx7fS3GehyA2xioXnpvY9/pZUND
g9O0AFsW7XbTPGPhwATiekEF3zijdVkdRUiVzuSbUyzNO9/8GDv6kEUKDdivRTtfjlNcNLvWytbp
1gsIzJnag469jJr8VcOerE3xICcG0Ciapj846a76VsVarL+M9Wr2/FnYZOYe6TqSeC2k+ii/UuIJ
M9zhifLtmA2Sgcxzh9CRplXb0Mfi6EwkBDstjFa7fZzEdciw7wZlLsZGAsi/18lno2VnfIDHgxbC
laoCLCngXjTnrf/iEEhqeza1N7rBkgJD8AnbaEkgiY7/Z7c5fNCEy8aY4m0I2C41VTvZdV3D8TaQ
l7f+l+6E6kmvzCmNPWKtaEfMpEPK/1YYHEYM5qvGhkr+kjoQaVwjY47MQ7z1n/kb3LMb8omj+r+7
ivH0dB9kxvC5vltoB8kCkgMYZcCSdVPXAairogD/WHlcrNQH+6QWU5+WCUYGsC4yU543b8W/DsE2
81FXnXhXcq+h/AJGBYwr1HmiIwsbgZgDax+UDYoOK7QlODCLaBhVOSA+ym3PZcx16F7lHf5N34ii
RZV90D1B+vqvBb/pG5rJF0WBaTK87i6K9dEJBoLSi5iD3CLKM6JMY+/0HOv3NSf4qVGxsJXjHndE
o+O72DCszsj38Mp0oHgCtafG9LJQEddBFWx58LyGmXunLq3Ik+fEBHfFtmRc9vJQdwh8ij5cxxoR
5zO54tIq+/+qTOJBWW9R31z0amcq1Nbi+Snvr9E13Gls/rd33FeGb5T25Rvw/SXHGdBTh0gMXgje
Q5SvhnYDmY39YZKY0Hia6dXlxacpBrE1yvc6810laclKZaFrEGdOlbD58p2QTJwdxtLzeMNhdZj5
gi9TPJ77hearUgkuliQXg9dcXdA+T2yE77x9EFvgtutrRZMnBzH4i3P9uLyj2Ibbp9Q0HjGc6dJZ
4AVGRel0Yjd90CuJ+Ks1WW0IqzdgTBnMHnedzwtprisq23/CPloYvplEezeJLU31A5vqTPpRtvEf
58GUvRQftbwPvXlAuHq3tRMuTSD2CNKeK4mJljxwTAeT58kb3YcjSoqRldu7sbUnFryrxvCPo2Lw
mm1CYpnUJRNAjdiwHW3fU0yea1V8GM8qupefRsiDBJsVkMbXlJjcMi/j2TeStrlKXBdXy5be8IFm
IPjYcAHHghhlKFzpVnIdyZnT3vaK2R/5Nj/jMxuWMUvWHQv7/GGfgZslOOfwGapoHlEthWrVdAMU
u9V3031C12pGVetf3YasveF4iMyblR5IOTF6rUj/IpLfK/xzbhVLjTLV/JpI07AGUez4SSMJDLNT
ryrmuiKJFP8aidLvjK1h93zjmsJBs9cCjI7p0CZBLzW6EWFfxkjXQU0yQHFTzUhBtu7prPFThQQB
anVKLRXYIOJarOxaNG0MXcSYzG2fW2PcgyFwHgXChKxoAs3m4ZLYxz3fVP9o80owux3ifWmILF0G
F+2OERMdkjDckvMCjAPzMcYoBlvbmF/WmmyqzK7CGHauIYhfbVLzA6rzbZ6t6zRj+QKhkiiw/itu
KkLYaGfbuyFamzd6G/owjaOJmj9zA22qFp0zzfdv908QJ2CZTCXOVGAjwcbxqGH2OUbU1w1ANqPQ
mrGkYplJczO1ailHfEjHS+SqjiEk0/3uXUr6JXN9Dzsdlv+aCEWSkKvVj1rtQ4UOkpUeqLmA139k
LrkxEhAQsHpV9fGf4SDxqI87Zl2riDGQIz3ow5N1lLTIo6QhhNVMm9snqzlqNWsBemUwCFNG91DR
Gj2peQLsrGFquaBhZSyogJfRZOw/r1AReA5KES4tI4ITlprvY6o9ugDMXJAxhLX7GK5W+DJF9bX8
4x6r8aBmnkwBm0dBE4VFVHiQDpxbLU8K5OsTDniABTy4LsKJCrb93G+FKYHErBp5kU9iFZx7EReZ
HdkuaZlHmDlFQoejPE78amwmFUbLEBXfjeVVRy3ljOajTm7PjfMR7N46zzml/e7Gem2BJIxbQadO
AbBi84k4hX683zkCgUzAlpfofsv9SgM2UHPWrIwkKWfISIafNiiybPLdh7y2jWYVxVp1fIfAtQlv
xGCznOvL6lC31qF0A1m/BFR7LO2mSrqe5kPlMEYhqPn+2jmH/vgA2y2NhPkDRt11XO31OraTE01G
lQ31kyNY9tqhHZdxi92NnX+6Y47W+O3+37eiV5WxcfNfGTXAtmQykwenPA+GZ4tEgpwegC535Zc5
Y9IelgWg7YLo2vsl6bUxhwF16opju/preiV7XYeKnI8BdnNwuci1Pu5WpRbjeRYlCG4DQ+8tFnYf
+qeaXjcaHWGDOjZKu4R7F/sZ0NVSJyT6sZbq0ULkzZiqAXG70WW3BeuQkHUsHJnVIlYrPen6YHuq
d/OGZTNZhdCTij/I+WanuJt+AnwrS21XrjQUYtixjJgWA7r8l0DeIsTQdFGQqds0mtt3T8Fak5g0
CCm0/2z8o6DyN06orqUQPQRddAdLc69HXdLQfcdTeajJtoO1E31xtoomuvmiscIuVFmv9I1uu+6Q
2p4qI8orXra9wEwSxhKQODgc7SW5tx5jZAlFsWYzHDzut94PyXvIK3Ojg8K9pWF+DWFnKKsVQUY0
LkwFTVqwS/zoHof/k3saV396zlyQkpK7Lm2Icvuq+owKn8FibsQDVKr0Mob/biMr9vairdhuor5T
C+sN0KIMDQ/hL5aeO1S2L89xMpYGhjBjvMz1pf6vwNM9IK1VafXJkMXtEdYo9aJslNWLn5FNwFgp
Ukn9KKLChOVZE1m+hAxO54brF0ZA1yHzSrgaJP7VhwWd+xBhPI31pz+qRmWVlCsWGD1NVKUzfCy5
FIpqMv0oWGGwbEB6ccj3/ei58P2MuuTTVzQ2uCmp+8iLd+O/DQKcXQaWGMWQ/UvAyBk9L17rgyYJ
OYdbxfkw/lYZuziBcFYjOM4nzUuvlfQ6bWa36hsgXPIykByZthlE4Gm0WmPp0bq6xx8SqIBsqZbc
4HGaq79XUq7oQxwF+FGNZPYKH+jEJFVzmePSRCBrxO9VwbmTsXWZDkjJfelstV1aemOdGjbjTMym
sgVUtOSoUhFghoRh1hfVhYLEodQGbgGUuhD3HST4lXDv00nI1V+ttJ1ji+haZgjPDFv2HvYg4YCT
pnExzl0K7nENdw5E5WKYTX0WMiaCiZY6vf6LtmPhcg9PSb4IjWhOGmnNob0R8KIlrCJF9sWrscI+
Lsdcgf7BwYg9rIAIedgS7eAEH5ndbUmS6aFbSuK1VU8l2L1F8A4qAzMC8EdBgOtV2uPMX3pVp5O9
Y0IzFy/oApSaoBYyulzLhIVQf7Mm43D9HkZGAO50SUsRiokZsNsaTXVISm2th1n4XILb7xg91KT3
uDtK6z+8druNFjMev4Sb7D7YkY+PQBlIvds8RrrUSJsDOfe8PuAU3TGtzUTQY+wy0bIoSQ6LeWrF
/aMSim1uqf43dwEqE6gDE6+ZPkH9p2pdejZbEj8cMOzvEwCYrrersV8fTQBNKx4dFtae2PORbcpO
BnVyfjoduq8DjfsGlIrOQ4pU0GyfuxIbirdP5CNq8euA9HNKJI0aIu0iOawMuQNgyzjy0z7peshf
wPQKjDkU0fk0NGEC+pjCqnsyZmnYao6/46i0zoxpbFX5kY4fxYwHvRqrJQqzJHO1zhf5xGcTVX2a
LC9tsHOZ2+KErteWXpjTMOdyck3JSOxis+cd3mnpRtHxrNouFkHqDpj/i7XZjiP4m/wrCS4evdtg
qnAagZ49vyL2+PTAxhztwr98Cg6NopkwgwVfSeE6Lbz3eI0V89sLFTub2Xjrqobx2sgXfI1wg1by
GiecBMmVMHfdu0P0E6fpw142dLCfHG7yKZs5k83frFLhspCHrPy6xy8y6OD8Yyfq/WqHuKyAlARk
w0zXk7zLITNdCFUeUCFBUhPv4WlGwHLjlHrbrEbgL7LFfYop9abE+WUfGM2DP485rVae6mJsXfsF
8oIn0MTC20B82m7PgSRAhjnUCNmoSJu3V71bHQteAgPaiLtwYYhGxUyuHQL0YdO306Y8xsMh0f5F
XaxZTnr6m1yACZxGTJIkx7X5b1x2gsnsfnnu0rmNvjiAWtwaw3ridy8lpSOydmu61b4GxVnB04lG
dSM/cBOZejbDfHxu4o1EFG5BaGCzxVgml1xZq0ssJOZfYNfhNTfbBzhe1a5gG63yl4PdzZ+Kt3UM
4syxFuRJ5mYulW1KFuEX8Me0Cq/i+/ViswlcTvAPdaff/0J70KgePTpT9IMzJvX1Y1ujXtAiYy/l
Qfx161/JQWiDPEgI6om/zpkkPPZCwfkHlAKs7sqCgHPaVuUfcDr3YytAPuWT88c1YCIQguyYd6H2
DOofsEcsI7KFJmpODLPgU13warVYnYoeMKPo6S3lwIj2L26pQopMuVyjm2QnkADxiUkr1RT1wUHq
AyvCc1NbAIp49HkHzGvKUsxsR+nG305sQWn6W4epIT6/G16h67MZVtu1A8QJ5zZNKvtgCibnPd1A
Tdihn1+JiPWW1hQC5er2Euan/daSzAc1Jy4eOPgeETn1iiDEzATs1uP0I9EHmNjkg2tgaHbjj4uo
SaIErGSXMOKGEnhQhEFsVsIWnn4349mVDsUIxoaNHHIp/0Kl8YHBfP0PCEpqdU5hXW26FhaOwfKG
U9i+CoVEhl6PjuKVyF5NwuCl+TpoCcWOqhZM/jgA+2qAQDqiDHt/JOijZFkdzaY0fW3dAD4K9sc2
hs9QWdwV7Vsht3GtgPXQJxXBuv1eFhraWS2nJazpU3lh2hfXe6FbFbc52hrW9twimM6GhlCYnivP
QZq4ZiYUFZBT6PKO8in+I4M/6Uj1Q35BP4uCw4HsklHSp38JIlih42cKH3IRFGqc/LYBCtiLdc+Q
wfTqW+QEp2CtcCUPd2VSvAYP0corwgTNoKf+ouch8UZz07YY1Dh+zdh/mbS4AHQQeuj2jNzmErDb
KXrZSNDIe02BmD3mgQZnX4LqmSGWghQsVhxhkSISRxt6ARH95KwdiR/VkVib/56HbAZIjbSQn18v
+6GoyqKfUGbcfM1nEllfSrOsq1dc9d9sYu1jenftSfCEfTBm+301/qXNj6G8vGi2MRiydTskIqp4
xhYAyt9XNL/q0lemhNxNKt/C7yy1F9lTni+9HYCmH2dJbS6UggMXZ6T7zi4hJDV3fk6jifhb+pKb
Q05LfcV2wUiwP2RXjdFeSPD3FQGjc6T7POx/CqJ77kICdchfXi6ZbfVcekZEmTwTceGON7a5IPy5
8Ono19bzm7FRNqqmS+jGJFvlR0a6bmjEHnUcXCYyyso5KKROSlXKT6FJau85D4Bzu2CQTNbxJGf9
K+WXPXbLRZPfFCGHSpxU/SXBMjSFT0Tx/mNGGZwz3/+/O1koZDD5il60TzdilGwRRRvrXkabVWd1
9ZPBq64u3rm+dA2iZo19zdV0dSbKV9rhCTF8MX/lUlwRkCJ9QWyAeRtu53aOwFW1/aCoOc/y5Yxe
E9tj9Gwd2AAtsyWpuihBFNdrRjmMB2i4wJHII83iJGG1KagSMr3a8cKh0nS6pr+NqgHIrhEIyq7t
Bj87p8N+xeBg5QZT7tKygY5nyf4YhR8cRNYfGmteG7Z2EisUCkdz2ZUnzwq75VaHujkZYJ1Eg626
QJYbZ3cXzOiC4PbV01VzD+sR4eASXl98AnI1vrsb1uC4rf3JSlkgzYZjCu2hqRX0sefUNByHvkLG
4R35NbCI1VtmAHiDx8BLTqCZD16VVfc6XLJ9NXK597Zt0iLP/d5vBxUlZKLEb50PI6KsYVrUte2B
kAjrIMJrIMjDCFRtn3BuyTRq0G30S6w57sVtm3wTXMK34lzNlUJRWdGnNT4zfg7QbQ42+2dkkSQQ
s4mS+hVkswHZ4donW08u1xLeZioXgPKl6xsw9ox1kVJ6ixUbCDgWgxgheeGnkxObAg6TZT17iKXZ
QyYj8eap7HZlTuHsd4tw8ba9CmfnZ4KVepRHl3mBFvrhHDE/T02aMXHVpT0BSE7hN1GL7mUUt/pX
1u4SOk88pWqZ080yaVwRflDvyXXt3izanu7ZB4E/VlNUDuz1uMHzLWzhktcXo/pvuJMu8WBagucb
vwTrkXSBKYrnYdC9R7MPAFex2pKcfkSQtCSC6IcbwBw8k7TPpgaMZgROI1SRPxK5ClrQg+B4yARw
pgO4zbb6iXN8vn2kRKMko9V2LR82FXnChMT+GZEhNEtyobJyFP5Ecd2Z35gu6s4b/tFk1QfobYSC
30EEy7MzEWf9m2hBVu9AdtOZyuBkHv+Ko+PxaPDQmWI0Rqqsf2w5J8peZqVtehGiYGVSdAwILOMP
7jXSUm9KcmLq7dJY7pVzy9Q03wd+vcfxX7omh7x+sLeWGEXHxrPuP7OGKPk4/fXr4toD4LTHsOfQ
JAOVxUuqVGrreW+LboD+IzDCGKVy0kHMX3TALQvQDucffXtZBRc6HCopqCaO/GpGTg7+psmN7DrP
BA+W1A3aYR8nWqtXFedzOuXM5aM9PTfQ95tq3XADR7OcAaC1j1hRZIMlh8aQD/KdlJRYruWfSner
IrhXZfYeIIILirPAFZDFDNZsZEgb5ZlUNTG5VvXLyp7ZtOqFsQi3CoQX742rnqXzMPW+4WajTg+H
o5tpKil2e5O6Z03mTxBcGvW/DDbQu9w3cn4jOGDpF49z0yIT1KMO1bwGQr+oDPVFahooulnVoVi2
dTE0oG9F7GdLPiJCSJP/zSEo6zO8YkxvC4giKc6ZvxYTmsdchYT3TaYfJe3JktifpoEg1WA94fOO
/oydU4DOqUS4HOgwAAQpEf4VpORkzgPXdlB47HprTgi3yWQHUXZOO9xC7HsKl4UECGF1mQw7oIFu
/yv7BcCDvE1ES5opL9wK0GREWd95hYVnfB27BrA5s9slW5zqKfGgIV+AUuKqQpDA3BB81T8JzemG
EtzgRp8325BA9bQeSFLF3ux6tDcKRPMM+W6aq+pB2YNZlCXtwypbMylicrsGiU3RAHGqIaUB+vJi
bMC8/urq5o//9vbhUI9PXZA8UjMuvGC5pjYSI+SAVEMBYXn23j8ZUhiSvSzdQVxz28/ueBg30LUy
kv5eI2GeYpc6SfdXLa0t/N81wwQ+XstBGetxUdXZyL6c0PtLe0FofbWk1JLt72gjL7Nz5rLtZvPc
eXorPwY46irKlEyzPpHczV9andjMUu9jYLTaEBaRN3n00MX3qOBlUsrDIE7LFMTj+fa7zlJVbhmu
TpwlugIewqL2gpOud7YCWmDpdVYOo6l58XfjYqZcipZafKVCoBrojz/hRUH/8/qSI408y5z9ba68
NIUj5IF9zyq9Lo/2BoL8PAv+kbWwBJLBftCF5RjSC9tDr1dxJvZFTHkTqeZxpisN2UmZ9XH9SqhT
cQtEIdY92z9W7f119Snpgum9MCak0SSH/9Mb/7fjW8Qq/s8ECRwB/VuEOGCNJh0WzoFypOKglCd5
PJ1CjN2QWwuGk76+129NScRYvnryXBmRdTwUasZFzzFe0zs7dUyMIJKG11+RL3OLxANsna6Hn1SU
ou84pGQhQKhq4RK95z/wNkSDux8t5w+naw4LB/6EGYd1FdyD9x6nS3OAAl4pOokaD/BgPtleIQY8
+hEiJpZCBREeLrq0Qn/sSluk68y5jbgB2PjqwgA3kyFb0uciKumx6/DFL9F1rD03VUWlqBnolFlK
8Opgk/MQTN/UeiNsSnzlvJUevo2iT4bXqSp42pgpkG0dV0Bebfn66vx8mGgQ7jBd3MjpAKlmYysk
m/V09Z9CPjdAVZcbDPeszNRDVMUQnWpT0gjUCVAu9lZ6/4FFICGRpXOATkIR5CE0SoX4/tQRHTq+
QoLeWIMZntSYL2062IgPY2RFx2qoR4JUV4RCj5FungpAo2ozToz6g0YsfnUC/KmKYnFHVzkqDL0m
M+gTSxY8v38zKCeGjvmY0smxtuF0sKi/yY6HKh0rrKXpmkcDFRPqo6JhazbLu12lhXJ5LTbLSOy2
zEvbUgjjN8k6/FYqI0Xv/TtoWU2ebxDRUkaylC79XbD0dUGNFglh3NQ689vHtislIpwBAKYPGkBd
FoOTEzdO2Gnywd1IhmCeSUBNUgP/htW0b1jRtbw8FXtwKeq/MxU27UR3fP7rOzwBlwCIpJOlc56l
Nuv1BxOXNbTy4UciIrqltyeG6G3owvVOyLEuaAATmYvAcgDeyDD29h+kzRDW1jsY8JvN+WMKOdVm
iCu3y2IDUhvv0GG8Mx0bNatfQH67sinodTbbdxGF9ndKgTZaIKn/ItxbPQ9mWF5jAXUM5qmUavhG
UvN28W6O2soScsTCDARgQcx5a9GTzrrPW/+OC4hcc2WWFx+K9hs1MJ/T7Xfe19QeYS0hbRELbplf
iN2kjZYi5rVrH5WcTqfmvhEhbSokLgw6kpAHe/Oq5HkLtyYH+tw8h4a1+DwtFzYuafrLehhDgrRm
nUx40OlhAY27f76GlCxzw4dE0fiFJccN1xH1vqIBxHPfbUdyGbbPhMvR3VYNOHls0v3cRRPbfuzv
j5SEXxFbPrnlJ6cKW4/DhuRApgjuEcW9gFFQ8iFmgE/s0Yd+6azGWhDQdpAPsvK3DJpabsBTnBkD
3i1dhD707LhFdMVZ8QMkIt6hA70GgoXzrr1LDafxycYKSmAvX6ChPNpF38/RyYCeFYbhYhJQHUCK
Fu+Umc2UWpJ7240HuuS/LLWZCM0WWazTw7qpVuc4+tpRY1vqqkLJdiYS4OFIusvTBgEgwPivLC2I
u+50ImR+e5gDpAVyZy0u/DPAYfOt8CdVYaOfAVF9gkImpWu2Y9DIfTJWEPzq1vX46LQXHwLMQafg
dGo7Io8h+Ok0XfheDpa9+B4LBxD9I457XtZGbf7Zk5HsGCJl0tDPuvUAoG0WmUfzsVFUIYEyEhhs
0XdJ4ISg+GxQIFIQEr3H5nsbM00feffuIy4UTVifEyfrBvWmKQzr6mOxIlKwCtG9epkm0t7fl8gb
UnnlSFgalTh2igy38lf+x+wRjQMo6airLcAicYykS6/lb0yOxvc2eyP2yCab3nfNqcmL2bVTKbe3
nCQ9labjsyn7cBUi7ijRLnyvPBvaeiS0JRzJivFqzwnzmhrKoF1KKZRM6pgOw3tqnBrNnwHyir+D
GIY945APWOYBJtJRzkNNop2kI+h1yI+e9oGBbTFX4rUf0PEvlEqDRdRwjkEtJHncJHSYa0fcBiDL
ZEuMkrbO+x+QAqPpJv4z77T7Nlppjbsl02Q6WFwtsXlBVMpbjuYZpH9Q9CegK6x7Vh0dUsV4Yfri
MRRab75re3aBY9sV4KhpcEZlMMru8Pv14G28QOHh3GbUtKftolurZRAtRtMk3Jasg22fnjnv/wDj
30UM+eWOeUsJZps/LrCVjFYqb5yjBww1QuQykZtoUo0pBZWCAsR5UBQFc2KDNFSSCa8CyNwDmiOy
WvXrJ86oGLW1ZLIVR5NYqWC52xRv83coEdNKvidsqEBRuC03zpplE+/wpDrRqjtGanQydg0te6FC
mEOqH672zRwAfii94yjaqyUv3FGdyPTqgcz6dVM8tfV3ChjOFIFCMDuxhJWyowtTSxDNaEVFEO4K
St72sAmHY+TqqLq2a3af3/Tl+217VGBv5BthBjcj79AVQXfJUvEa6QDi3mjIbWj11u4SXQ/+mSf0
IY/m68G5B8BC0Q0rBrMCtdfR0m9J77cghnztKOSwI+bO0kUasWJzKQVEVPxuP0DWEBHVhqOwMO1h
XF4EfgDpFNTt47ib7zqIy29Bw8PYCPs5I5u7IY9Jxwu+1R5T3E/CrDSotZZ6x5PBs+JSnD++PkRk
SUShw+apl0Xug3zrhrLhxc44rf2cyho6yKnn9uFD8ydIaGUszSqd2HBdzJ36/XrQJTB9RuQYV6ME
rTaJ/2hUmg7SCYthRQYMraIDq0KNUiso2H1IPTq1Y95FKe4Q05yF40IpQIK9hAafpe4VCQr7ZzCu
hBhQPzbWtEBqjWCqt0PeRY2aeuhstrcZNZqxZurnfsxfHcnuHeBrvpnm8KqFX+NQ6Pi0/Z4fpxmQ
3mZsqu4mqITNkdGrIHKyzL8hRfScUxR2gwGgIUxTdVN1hGl+wxoMh6qXCpKH5NGi77FBpl5xhXqE
VjnHKmKK8P77Wcz3Xiis4sp70FcRgjfpfw7goj60nVTKowsmLRrlLEHT/qIjgGjIWvP0PkNChKly
t65j3kJYs/Bjksq3GBMJoZ20DY25wpNrYViGfer+gBPTLd1UbpQRV1wJgBL3t3fMYhSxloxCPUM+
5ZD2Sjds6IVf9qPrOHF1SOAxfHIegnIo9wlgVNWpP3ZudFTg+KFjrgHfKTtTY3peTvBHJCYFmdZX
+8623xi0FvZyHSubRvASDk216DjsviKCHd94k7OGlaY2+qOtoSmrbplzagNTtFmvgF1PlM7QEDwj
30/5LwhB/Q2EwpL8WDXUUOqFPjV8t++8z5kq5B6W94H/MFpkSWU+dI/zmqF8yDcmkRf5/FJhaRB1
tp7AXAFA9FWj73I044ZXeAhsfWc9eGVaEbp1FZTUoJk9hi6MkqVds4cXG4639wyhUtHuumZOH6MS
qb6YA0o9yRc7jO9o4/FMIpThbS0WHGxP2KxonNL9UNuyfsrnUcHjtKn21WxmBQDovPUDskwNxXi3
7A3ntv9DUcxpU5TUMdtA/Fz0OumF/umSzidKpcmq5YNCUpoxff/fUuMfY+/NpWk7U4C/ZV5cpeAp
ykwR4qDm6AbHaeWB6TWDxCZshDsbaC7N9gyCZA8R1PyUquPQ5x/PnkkRrcKCnccfuiAwsKYT8u31
iDoPcDpkn1k1OHNxZPgJR4O7DTiXKt0gtTI1veAHlIWkg4NdGmp7vKV6Hf7abisIZUmfuwQcAFDp
mgGd44TpVLpz/xH+YFsePv5tRycFhQZPifD3U74UzjEk9y6u4+T01e4ZJeLcB2zWW7PO3W+5doBZ
PE9ZoJroWZKncZhmQ68g6rx1tI8Y1ZZFi4rasJaioTb5V1Oe7Ub966QauC2NSwhqF1xwpGZAUbzi
mSMgKKILAfVvONx1vBVv5Ltrz1dOwi+GJCHb2HZ/JIeKoY+gsTdlgwIDQfugEOhBxlaE/23LRSLI
4u/9xyfzdrhm50O8gr2wRZou1rpetfrtSgs70XVzBCGD5cnZMNN12wf/GYeGxn5knBlwl/2ZWloh
fGtk3+/2czTR+KOujjKev40ctMrBcxddUbGY8h/Kp5ZE1LtsGLEHbXJAe8AR5yz9I5qkKa3H7V3s
MxORzUYPDSif0B+OkG66I3i3E9uegFrS5KLgXn4z2MOD3I0TfTptRhDW6nFUyuNbREspib201nlC
C2BAgSmxDXfPTLg+pzEHUIPvxLIAx0FMdAUpqaFdhWjd/2ktTXKGt5O5NRxlG9Tc2eOWvoX2l5yT
tnVhIXbewMLIO245N8c2J6AhCfoGRKfswb5f2mijqtL+sKm4rQMMCCuazXsO9lweMHv0P81BBKtK
/z8Yny5AdF0VttIhhNLxROq9qL7jXRgxNZOJ9Kaoc/A++0w3JNW8nj1hMahshiK6ETcWh8Dk8cIS
CF8tXKdzW97MyS9qa22/4fusrasiOrPC1ivn4n1LxPk8CInJYzARfoG+iBUpjW99+dEe4Xjr5LpR
rJdBCdrtx94rEH3hziN28/o2ZOUxH5CkMgyMVFYBvLz1SvTnWQd0JI2Zx65ikwY4ldRqi9SI2U8N
euD/PJBggCHriHqfEhiC8nC5W608zw3L7+Wyppwvf8vH+A++rWcnrRuf2cnxdS3Z9KysuONrZGeL
+wHNbAMpzn66nqPKtnoJo0rM5ky7lW0TMa0vtVJHLPR4kuk9b0dhGm7bEHH47+qJ/MrLB4rKpjfu
KNMm9JEb7w/9RcGWGJ3RZ4n12jXjZSNekEfFQ9qbIdIcXZabMnXZtSathJNS4j9AxVsKFeHD+hLb
wrtsIiWZ5qWd7WwyqaY8hIFewa/Q2Ab/t4pxKNDWAikvI+e/T5ztrk+fXbTAx0UlcfR6pLM8HWfw
DcZzUhgvFJVJTu+GL9IMWGWcmIw63P+2nXfu7WodURrheHOt6dxhjiXxtZYyHsuO3g/JV7tcS7xb
LiKsWe6WOYFInwUAwRzRsarnKtL/dkIAwI5kcPDQeF6fBKW3qnkDky62wDoeSyhqsaFrcbRWgbH/
2NfdwqoDy9OzfRt8sqYTqL+P1h7om3huwrnpvIGqLfVVRTyMoOidl3KvoSDv8hXsVtimTVxNwrxm
K0llIjOhDyE5D/PHxUkgpezm4LI4X5osuh9uqnE/2OIbt4n/f3MDax3yZFvj70vY2xZdI5eHEOPj
hajv5ae+lR9YiYtolRco5wlVi2wYxNtgSOlNqAeGh7Ng58HaZW8AuvI7W972nMbpfFZKDLdLUldr
ZR23pJ+2TP3wQ95kyF1exJQ6Q4Geue6Zz/ewzwJqj5qHObjfzUjR6gkmW1Jdzjbv1M7u3Dzvb2vi
qo1i2mHy9SChVl+VidIye0ceVaCB7QeFkNU1VwgphK80dBxFtlgjRbi0a9VHZ5V/ojYOmZvGgFuM
22dDoUnYh1BdJ6WnLIAAIclObXeJIEJMqezxJlTywmnWapu2dN6i9f0U+MYTV8FwVwhDWnihoLJ4
RxRtdTNhweNyY8MuWh3hmjePFApSyhi9bOMOD6b1/iWUKuZ4Uz4su8Vo7ZubjCez6Y/dzR9qujjU
wyMf9v1Tm8ksINnqjbGJgg9LIMGEjhNoUjhSjE5cX0N+aX5++VMTHnyQgmJnOK6b+/CoaHHnj214
BwDnOocWshFB2BBl7G+Rn5UGQcl9TBu0Fm64AMO01LUJwxFr1/vIpYOzBXEw47V/QVJo0cetQpQc
kADiDzmeQrct108I4I0v+cSKx0GPN0sVZd8SN9HXwFEQvlqNoKe1uVorlUlm1nEJL97KiZq6n5fe
rZSDh0xEDjrAVgg1+SrQc88Mq/zh4wSKw9y3GcjR1z5GkGwOtAP+/I4FdoBnGqsWO7B820WeWLGk
FFDK6XVTnOhlo6+VtkVZ/rud7AkK6VCFNm4YQoReDaPB49QoMOGzxYO0zSonGBDCsSszIyZ85I1/
rZ2nY+m4lsCLdzKJf+JJR1unLrq0nLxWdMUodo3djBrlxXYl5IkVeqJfBFyi7MjfL0Gn7JbDdMex
Q4EsVTIjC7CzmpD8FoLM+wadX6mcJrItSxNGaUpLw+bI5tD+ISZ20FYCKSZC0dGNLe+Pmi2Sl4Dg
h6886s/CywxPeYdWRJoTU/UCmwE4G+2NsEfgaziGniK0Qcgogsvhlp5IiDO7PqJ85aHgShjizP/j
8zvl6dDo2hx2wxUkaqFU07DEcTCE0kwsMBWegQ+id3SUWRQV063CX9H6iisH8h4+9OnMbBj1Vrmk
Lknk0RNnB8cLJivzOjdEtRqlDuzSN1/j00zzBXN2eZ7p8tf3cKyZyUCgL7+rGfmL0HhZk+T8XWYT
oY1GWRs3lMUWzHFIG8nwrkQ1j6NQOF8I260E4UUX9YtHGsQYL2a1860t6W5+L9I6NmRV2mhhbkeK
843E4ftUp51CMyfZuwULOsQwtYyk0CHXnsQDcvkWK7EPNwLa/eGjK0a9ULViIPtRLMTPncXN/nXM
V2maaiR7FS81Vi1v3Vzj8WDKELJxrRPUMsWh4R1nPgv82gpNarYBW/5iZFF/jH3V1kELeKrVr7zg
bf3mq167jrDUVgmlNJqH7TsGjriEIObIWlJvlWzu4eJpbVn+OYm6B9GshjzQhNs71HSnK9TyHbUC
SPQqxVozs2Zx4NqOIppPIX7HovsGW1BdrsNSQHzfF+5oj3fD+p6o87wi2cT5KeBHFPyBL7kPOFD7
Hu1F6TZVkCKeoRoC0RnjMguSGvJmB4/x+jaU2crH9NedS79VvaBVIZFjXTXmYqXhR/hrb1cSnqgm
8Ts5c7li2jZEQ8vlWip0KKGDIOacKoSO5WpYEqpXhjFOvE/xs9XmMZ1hGQy+CBP2Zm/Y1NwMNmwe
MznPSYoB4wW3H2q+uPv1ycMpHBctsgZtLX6vfzxuvzcCxo3jvTH0xNOgmpjCKHXC1UOm5Y+yXypf
7mlISYBW14whEFZOqcrDTHVioaGrKOPX7bZshIbdyi0BQH79e4qVd8UFdb77e7cQhHO5yvRjI3zH
LVkl8EFBhqmyQwGSoLxr8SawXWzm0BMhBsAQode0NgaTtcIGQ44lGSdqhLC6kh1lQ7aMEYBvCi7z
8T0nCobFY+fvX7pHslIvvTuOAAcvVulP3CY67RVgrgiY6WpR/OjA+RrB8txNbroossDfr6PksJ1U
fqIYPHbqAsjvD9xNQW5uz8Tj7QlWz3UOka9xj2Q3MZnUCT/9bzwtGEUGY0dntgq/nhfN9mFeH7yV
PuNpJxy4xa2fQngJMsmTKUz4NZFsEgcocSIgS2oq45AznlR8g2/dh12APzpBdoptl/etZGe1DJOV
uAcrlTF1BraRCU/sZgh9u1UGVetfx37tIbLG2L6prnZpbwVSIAodyl2oLHWp0j35435FaVciWORP
LYVdwPRh8QQp3gLWsaE5t2IY9nuwx3Oeqwzv9jIf49TBIaL5AgywClzmBHKiGebCwsgX9Hf/c01Y
eqnh1SmtLpliJCvbwy74lRNpiix+sZ4kY0YNTk8V4FBnLjJ2mM1OX1BgBxE8U0wo4g4GHSKR/14m
0Xc6XmpQZpVJK294ducxuGr/IjD9906acnN7/cU2q8yVUcQj3ySK98d7FtpfS13z5zEz1aPo8/6Z
1TDmwgnMCGEXax1uAg4F0nRrAGgQq5kthERtrVYsjtujcG6qzquHE4f08PBQs5M35ZlotaAxR8p3
NqCdv/Mwgc3PfFqwPQ83JlSkrnR+9oIENhbISUF/NL4FwqDqkvmTvqjHoyRBCb4Gjl8Uib3JY0na
z+AjNN9scrzrKDKoshr/jBhiVoqppNiUTI8I9rPlhYn/qwjegoJDeIurmjrDt2DiuDY9Bnsd3SGk
jMWZKE6QNI39328AygaVUzy1wS9rtwQSxF3PtpyEJZ1oPPHZR/Ox75aCkEipQMitrsVqks+oaVio
5K4mv9FUImfy6vIu8rb9NUAOKpq+8kNzvjCPygV9E/qydWX5JUWdF4ub0VCp/WMAwOYmjouFs/ac
Bo5GFhhTF5Qes5U8nGnSmA+SZS9axekkh0z7//gngZV6uZsRQrT6Rov8wL8kE7OwgxggoYgeKGU3
Lj0RX8Gl3fn2nKgUZIbzIMGesGnomJvieHD7NeuzCfN2Uzd9R60doktub/GbaS1lmDT8vymLX1ZE
Tx0I9R/tjemV0h+VYoyPg6IYR1HDt/yw7ET7pGmBiqWzx6Z6sawuUzLdyXIT1eU2+h5uf/yk9MRi
3Kiv4/k2xA/q3ybTGDtDGrY0KGop2RhjN0TzeK+J6CvOlDjxc3JrKgzksC3FAiyRD6O/Jf3hZKG6
4FESDaNKRUclACv3VyJ+iMs5fBem6vr2wKBkb3orDveunFEw7iC0OdhGtyucV+tCcrWV+pL8LEdO
rFbxlGsZhbDnmuHjVKg/9GaBiZ4fjrE1w/xgeGWt3MPdcmQb6maPj3XrUR+F2UXgAmRwk6f4fdQB
CBN5XURcKL/EORbdik0XBZgiIP3uw1pdjl/SgEi3bKvYYSUCWHAafwRQESINSmRBXAUtcJ9WrWdd
weuiop6MF+9CoJesOX4dfHgs2cfJv5e5c6zctyG9knYKcNRNQEMZDY5qNTDTNC+ChBJcxcQC42L7
A53U6bDkJ5R7RMf8t6c933JA0r6gLXtBVjrVtm2GIeUAFQOl/JMf4omVbQnQKsv0fFJ1x6w+U2Wu
Xfx6lFoBGW7+7VzovXr40XbV9GvvTCOKNjI4WvWPiWSdNWkUmUvT7cpJw/RK7tRNZynRCO+Avd9K
1p0qrxbG7gEGfRVlIRC+A8O2fTNHUoUpZZghBtscDCLFUIkEpmY3kIgrFD3YS/zH4LPhtnQ0w4DC
MIKriphA7POfQ17KwHUyJx61EDTL5VKvbv9tT8swpD4Dc52Ue0G4wAfw6Sfyd7hW7k+grpBgEAHu
W9c7Hi3hxJmuLgU8oq3j8iRW9qN7T5BvOrcvcRZk2ncobHGJps4mkfmA/VWHeHSVH5xXZkS49iWD
BI8nycTAUU454J5ujuH1Jg3hzyLCwyl0wa5QT4Zw5Dbsk+a84zxJd9CVLtp64OVNIKfMZs6sDoJw
cesH0PTu9Mo5AT0BwW7GuRXszySx2Tk+OfKZ7EusEkVuVfFS546ED0hpVWPB/dz73oh3RgAyTA7h
vxx9JSQXp0sQGidN7fqzCCtIU9DP88uMN+nXiCPaBrDrKNyKzpnKG6gyeXOnllP6xxS2Ukft0/PV
A9a6+GslLT6VRCeo5yMRFj9vmie9mmPeRfUWKlerZAySySC66xthX3bCe3xdwrQHOC9uzrzXyVBp
kN8uUHIfF42cPbwU/Kxv22d2/pK6JI2DyIXwTh6GloufEL9SVk1uI2jFcW52bryR//aC8wth7A8U
LwntzFhJDagA4EwOmep9DFuZT+M7/W6hrFCbKvppliJpjJCVJRPYtd8B2Y86laGjJyAAJuZ8pr++
fI9sCI/gQtKjMet6feukfQShPaCWcNN4q8XIuBDLqlba9v5lZl4fLYCp7RW0vlc2werkbUWg+FRt
bEzgLu+C5ry1vRJCFnPzfD+CN0XEBp+oRUzKEtDL54+PN03ST1Gm3cymA+F9cdlxENvdW3u11tvp
oKMMN8rR0lUSy7fZrCEm8an8OezF4HGUAdbL7MKOIqLSigMtE1908s/CMRCyYm65RR+Nt+0Z6qmh
f2o6UOgWc7y/MafCpo4QhMWTcQjttl/88Mv67BFjhksICVcd9ozH3N7ToXT8RIHyLJRJyYYTai2Q
Wss3vkfJBNnZMJt9t7YLpAaIcgj+JjSwCjpw0Gty02L5KGBZ4NKDw0URZB/Ob99NCeUOPxMewpWB
5oyllQR3iDfeaYkyrFH+1oBwVTbG8TlzynJoAgViRQUf4oOiweB2rWfO1+F/IRxSa2d6D//+KuEp
PlhrPK/l7DpvIe3l0Ez/AH6fSxKv+zFK9U5fURUEnGBvqDk8pH3wdSJ8VKYrUmy5EYlyYGpa4OqM
4lgJQmpPlbdz4DuWXY3gKICwZQkD8GXnmqDAAED/ESUDHLAmLN+psj6IG3STJAgRG1c2FgdH9nYX
V6keWD78cdlDaG+LitvJONfm1u4Usc//rEXOFV3PO75FhHZlBCyDRRZrpKPGUUmZMcO6Eu+5uqX2
FDgO7rCYZ53Ye9P8mHIdC5YUqYvKjEqpFOqjbIBFQk+nffaETSu3US9mgNjriTDc2EWuE93mgBu0
GVivRzF6i4bgtE+q9aQTYHZxPXWm68BwA1zlWqW12roaPFpIJ0qL/9qVFNnMWVvpIUkjWcOomyml
PyWY+JomFw84HpRuzABklQa257q2H3glWnuh3TH5ub9mQKmSyMDfARXLyTHpYBUdj/tAcS/+xKYK
TtZRIXjTsk3XhMfdU1gOAnSDKNqxw+xf2hBKs+x7+GXGLCKTRQhUL73d+H1E0jrNqas2S+1xKD8a
w0k3jDn+MuO9Fg1q9PF1SaY5pUGXYH2wYgqW66WS8XsHACn6Hh/61iw8E5USSq+vdfAo1yCAy0We
bm2/p1f4RM1c+l/g/eCziy2VYb+Jva/pLMvMG6cR4mmXfyncYf85rfbJUKqFcZa4768Qy5xL6Bhy
rfpmfm313VJykWqBj1L4pL/S9obi0VbdDH8ds9hPUq4kM0XGNJnWOgat8/0BYgxjWDlV133ErBZ0
3YfxSpqfVIKL/k93qykiG0QT4KgqLpp6PhG3p3jU/bzgp1X+gDS8Vr1zYcf+/Ux8Lcfsdz2GfnuW
kHNJOkNFy/5woZ7Kc6kzZ+2Aaowd0G+HgvEEKZUtyKNhjWbTwMsaVJdumwE/xGRMcZE37rbsEi7z
514N16OQ23jYMB+r+nq32R4RkWj0nMUTrLRM+rHFeFMnnNT2T7ix1+qE6wbWuC4RMzHjVtflnI+7
LVl4S7i1fTEVu/LCMMczybJbo3B+FvXJ5PzFwFY4hdht+/+pPuFXc4yBVzPKH2cd/YeKxGBBYTmp
GMxGDjnUhENeSZGO1Jg4rBj+XsoShzdnbYsU90PspipianiVDZoN9FVdSFz7OAa5MxUQMetmWnzU
9TCgJunG0103U/RGvcvj9FaNgQAH0BR2AUoTbCZVNXWOWPJdhk8FyHmM0KajfIrXBhh+SYv1iP/v
8s0tiGPuz0jsp2kELkMqEmdPvvwgAh+T/a6FBlhQMEDYyCuJA6BY6uqqKViSeluxkpwks1aL5G1K
0hEaRGsuI57Wwb79rYLIRYskRVZCgeCMCf2Mf/9tai5N9QcO7qqAQ4pkx+RL3zdb2xOrEcZ6rnOw
uxn4bjJjbp9fvyWXUdLMskfsmtdjegR+k/BFb6ACfWFBi6ojWpWjWU4IKHbpkh0w9wtikrkYYyQF
Ly1EzvAQW9eTBN50JbJInZ+fGwEk+sV6wERs8O7iV+9pgEH6M2WO76fx8mxY5EWtyzhlGswnIRL3
exGtth+LbSJ8yu/NL9DzNirWVKUF7UvwnaamUqTTyNtRXi8dV/zzZVDbC4E/tHLYWp5/Z3dNGB2C
Y8usL+hleck4C7C+YTueJiBlUNFfIA34pxtaAwn+vtSfXzf2EJ7Tw5MZRzyKwI7qWFMOoz7jOfv2
d85KgtsBD9RSnVwfTT5B3qKdd4JD+QTImSab/ezI4RRhXTdQbbVQW4m3cO9TRNo8wMxgT3cPI2oR
+FRdyiyzF+MeluEOd6oJCKQA1ynduBThd2gxoSTPqjSJwsaN+mBF6dc80ny4OelkVP4JKW9r9RIU
iAt1eFjvK3nnfPIDr3GgR9sHAGo3GYnVW9EEM4oEenThpXsJfzErNoi0ANbDC0xsB71ApHy51TET
YaPSI3T5VO5jeNoWYd+To0NTgKsWsCIfhNppjdluqw2YdZz8pdk+OLKioeY1rf5j3KbVFXOY0NPN
hdyDDAMMpQ8QpTn5LWLqvAAflfaj84FPCzWM7/VSwxM5ST3SDgkQBtW6ZDqQhR2a5bY6E9ghnYZW
S+L+aXIw+2nZYXDkBsjjJhN4d1fcPOPIOO1kYTrEfVP9Drpd7WXNQRebwLgfgp/9ZDwqdb2svJHP
vGTdl8Za1eIMWn00F0dNYf8it0WloN7/Z13sudKjNxAQPIoszA1MCVB1yVQOUJv7+s6rW8AXi/0R
HiwG1tNgJQrcltXqDp9LH8yb5nzBoQJj/7wnAfI6vzwWzCGlQgh4ZS5FSH0VH1AX4+EiKOdhiPxC
WuZhgE8ketRQP8AngJ4ymOdTVKIjtScNJrdQlSDt3265rFBz1r6tt43MW7gQj8GDLoLaYBA9g7FF
MfJkiog4rb0ro7AiPrw1+HIXcu0hFXVpJZtz6hcWa5y5wVsWSAg6FV+xRTBCJTXiuRfKSh0FEAv4
IP+gw4+ucwaxFoMIacZDlzC4rM9ElSSV+wEBkBxpEkDxKZhUx640MjJVz0ysjC5Ac3mB+NFG4EgT
4dUvOJTAruld+svlNGRUfKu1s9D9p9oaK+BqVWvAfRAfkzB3TChpbWTgQ8sKoYCVbKJkBxYZv9rF
inARZXM1MhliT1kPX6x/IWacc27+/gRcEWXKyze/OdXAC1xkNYGSPIEA6wXgPvi3sPlrNyoBqZBJ
Rqp9myRPv7kGiTLdI0xRR7I0RFpu/cV4FtnMw35qeF8u8vLukHuGpvVtafv+FhhZqdeNMWyXvKvG
cPDNl0UF/Zo/dVkPR5isDuvvna0buDp8eJsd9iWGC+cWz8EJcknzZjkR2UZCdzsRMWLIfUCS/+II
XMAbYr12sqg/YNYkPTNvjaBrVcWbsnCDqWG7m1AUwWJgnyfTaTGBVZgB8DV6zfjr6GqS4swmVNWY
9qSAn4dt0xpGEV2OFoy/n5HC5oGj231Ax8qRk9Qqds2zPhzKLdWT/sZpwgLQuCwBjWKFeRJ0QyAE
cHdH5dgSZBs3P/6Y4nAOPsHl8Y6h5RQz3zE5QZhywB59tl05o+gec/pIoZN4EGA5thhw5o4/owad
GrjT0UGz0skcFA6FKh5ppJZ85L2Sul5BpW7Zk4ClSbUgcEdQ/sNM2L8ieo/rPttpRa9rG3g4ssrK
PA2XqxNR90mjaQMgpeItYUzKpqxXk1mTK+S4sebIoffSY+afsK0rI0CAwAMlq0LZUD6GFdAjigE3
5JTZzgfV4pOxePnoQo++grscr6X673cM0figk9Z9CgpBTxWf1J0mkSJ41Y8squCFxI3gxXKQzaoB
OveWQf0bt9ltgyAB4Mzj1+1R+C0M/SsmTRCQ9WC0ICp17cUZcIHLd4rnnycdGE1DO4fIy3cxYsPg
YrkdzFBuhNdRPu3/NGsHnHEAodJnoFBjNOlQqITvwGcNNh4Qel4D6tfVfTDEqOEHbwCeMlPtVZEV
bjAMfwNYGnaWZ+qSJM6a2f88LJ8feg7wiUMAGG+s2cq96Iz0tiMSWsWhrhsWzUfz+YLaLWjPQtEa
Nw41NNy2cn+BQGTqmTmaANjSMSrxY2kflPYLpMq4BzzyWPmE5zPahX4MC7a/+jZKmURrM9nzieAq
KXaFILaEiGG1EEZ4NGdXbtgwhXwsaCnGm9LbGuE8G4Ao1NCnwupxKteHLxlK1clXJnKjX0QfeGUx
pG3/Moy0VpbgF0JEw3TX2CcXq27qUjRCRSzH68KBCWCnIXdJWVKdhdlEUY7uZM8KFPjvDim6qXHW
Dw0eo38a/dFvJI0ZjFzfGYFkWae6sxp+h0cebvCcJmbeXQjePowSp8QpY0Q5764gSY/y9ULKHSvv
bceRUVxzl+HSrC+f90C/JghJL0gRs8IuZBqEZ+DsrHaY/fq7mcXLtjmIiBeCxos6463eFT/fN3ws
vq0ouQcPVyVa6rLdgeR9+EGKrTv8fGDtXyis2NW0nMVTNy1LtJBzEBvXjv8cerF1qzyheL6upL7k
dKRc4L5/yZ9Vo4jQQFG0XjyqRQGTLsi/bRRzVLmAOIsmcXAzO6SCvup+xybS5DpC1/1eVS4EUgJB
0rqkq3lBQ4f7q0Hruk5DMqM1xpJ77ferTK5Ll+Npo/6JmTAtH3n9tKHyTvkFKA5fhhUpcbTkfq49
VvagIY9wrPoSFcyPJCbjSHB8Es0YZ7GGPMXW0dpdCrOZVyZes1y9yMXECv6gR3UiUbmraNfqlczG
L4uIrS5DH1wxxIhvOkgU0uQwNdjHmLd3BRIwBITCUhT67Xvnk2jhYr/rAR5fpGPgz09n3Y2PkWoQ
EE9BE1GuZCF7DB/7L3xrRJiNGPISLRQ5PIqe2nibYR50yZb14heuSEwZtpiiXeUdvf3dIcHy1Eka
AGRCeSj7aYI7m+S8Ef3Kl5hoc8rBVygxWPGtprpEivZGjBUsRsSpL+vecpj/E1U9r5OXono8Uu6S
cTvOdZ/6pVqxXmdj1qeUwfQcamQn/vwJEmhANOlPldrsJotLC86ofoR0pVpT5x2nP1bqGmru9GJh
J65Vj63LuxynQGWKRcsbE9hkOJ3xI41JGX4kR2GOYMTpMGd9UDxf96GxFzaRAN5kyDsmbZg1Wb4n
68nVA3cMgrRecxUuOLHW7cQmSHw4SyktsDwNqoKWF1lF/FOKtZHQftMSzfOAcmdaTkAQAUohzMHu
vkmovLbyQ2TExxHPsCWDZ+wl2M66xeCaq+UxxncSB+3f0nvzr7vfkUzYr7DMfqBX2UAcg46y6A1D
OeLLOwu1BBw1mtunUxhyhkL9pb0Di0YZYhQpHJo8ZZzei6ydJIcp62UG6Va07gwEcAjWCtZj0F42
FcoLX+YXqFR2vv2wv0UrnPmwmp9P0nFpXThljn+1+gD1eKPcxxU7HAHy4MLKAldV8CJz4aPNvOnr
CjkwjbHS2SChfxAcAU1WX+7l0nhKb9lxF4hlialyHe98fnRRPrJIHKkvyavI2F6LQOgI6ria50d7
7kcY2Xbq0AWLxZnWDHgxWWHlalTsLWPiWJYFqUmlsVXZeicYCxq+fWH83KaXNFObqAg/VK5LJvTR
9xr6ImE0J4sKGrXeNBkZhOo4i5FrHNyLUC9UM308sA4PiaMlOBUkssdQrG+1KPglNXBKKl5cKvkc
S4sITiSgOOajKFmJR6fgmy7B/gojKtZZgWK1U12nSOdmF84ohnwRXqDPV2zYdng+OC1NVnNG26wy
GGCAGe5PBVIC+8BtrQgb5+VqMLafIE2aw162m5db2HVgg259A97Z8GTNck0SDVfZqZY2nvIAQHPL
jkBemT3h5N9WCNNslAN1A7qB6XLl+dvb+jXp0DRXFBDVN6EXPUN5JmZx/07rnvtg9nJ7EUQJW5Hv
JBskX5ABxOepp4Zf99P/bbKsDSAaSCEUpdKJnHIdqkWOW5hz4yt0uHsB6pI+rqRtjqT2JClWPjze
nvF6l2/h943CYmbuRCjRleRRnrqgmpXVLB8Wp8FNDGs6SlKjgA5Q/WTjzqaCkCggMHqzjEavPNQt
Cq+/SHizVJhj0ZdD87qOR8YsvsxX9Y6JSR8C7wG37xK/FFBoyhcqkbn0iAcVnN9/B8Dm6L3APvnk
Fy64NSJM4fQjjH5x2ZoTHdpyzWPqfD78vzl/ISz41QlfW9iGKJeQtOHzdPAWBsMZB+W+NaoMOBgh
d+DGi4+XgXiC73GPiZ8+VnxjQ9c1YE6hitdgUynhVAtArs61TghiXAwQjAW596Lf4pZKDzUtB5j2
JlpGla3oODNWQu45C6drwsFNkCBeC2E8tb1JnJ1p4TrmSS3EbX64pM00Q3A45V9OsB1tMWsX3Cdm
wQXw1oXBMBVuG3orKr1L8xo8p2dR2sicNRcs7+rCFQK1pTw7G/htdCUhnFIffJe/+ctzNYHbSOj7
92SNxoIxgs+VVGc1Zyl9s2fySZF4RSiLlae63ZpcXH9NFtOLjgujgT0N52yFbGM2aUzEQv7/t1QW
k/PZn729/HjyOL3cN7cFE5BsamNGJRWsreZcb/SrLq32CUECnJMTOYUZFFnhPny9ByMk6Sp60NGS
IVlII/3RO8C0roNfCqXlZpNlmokl5J34YU28f0wnNNBAj4Rhx9OcEmZ8/hUrDtfGghp3ukt1cOkQ
V4++UA66h7bpna1/VHMa+JmWMqdpr+DcV/ViaFLmZSqYjcfk0QmvlMVQQNuxHd+VkaG1/BSDq641
N8kW4rxYQSy+tJBbgyeFxRTQpqVMghMEd2exP0A9v+ix+o85oQi0EuQY2KqxWt7ijyx8BJUd7FRc
FBkKHWZxI0brtPhlAMZcBd9VUr9SS6Z3pYQzJxDubMpMuU7XHScRKDjaRzXOdlCQh1xb8f81Pzsq
rCLs86e+7wXAL0Q+pA0yWcPNP4LXQcpmbC+XKGtD7TXdimJodC2Q45x8KrvUW1w4QE+3eNHoHOde
4NaCL36Yyed9Ef4905jYvcbf9DIhwDntUgIPRj0L55Nl1nkaTMNU4HlctEZsrEoBdVA6VYIqyc3a
0Uu+zwVnMRZgyUyhWWQGarmfFzZZpAwPqUs2NQhi/59Nv2zB4/9mUGgflzGDuwkdn351lb2Pm/eS
MLP3VAQbY3lCNr9b4tPAcxUW7NQFEIaJrLlH7XK16tbsbtfCux6RbphTWllkQnVSDUMHhUySE6Vy
fVehPIlpKNLxVHRPoQWDHjq7XpJT0vgHEizc4h7rxxCbtw9enMOfkSH/GahgXHjxYkl4q5Ees0Vs
blTSYjRRjOp6Xm34sdmxCxqWMh+8RQqqL1QAW/Khxry8yD9w1iXKSZXo8b15oSEbKPoQDJIfF7QE
3RHHtl68hpfd0QWxNQpD/Q4FVvqPzy83i7jvDxiXlkheU7DpO0MGs56XoCYVLplOtO8DxoWm7vn0
f5r1nzZ+gtcv0KSGkwMllqrZZNFJibTlBS30UaNZOl0LL9ZM3uo+/0nesFRwHL244/+MORICZdWa
MVE6MZIY5wtFkT7MQ7nYzWQLmeSBIQRMCHujdUUwt7b1HlOVG/72cF9lmM7MV0EzZ1ie5Jp+Os2O
kjnK+67bUZoVBgRbJMgRHcf5NMPrPE9ws/Mm4dq9XeX4dej+mZB7u5+m3Tx6cAhqa+ot30MGPFMc
AcgvEdcnc41Roxe/wcU4AfrUqYXpzGgB/Ik2RfNceRMY/eY1Da9e6PjWxcjA2lss9GM8dj9hQFZU
XVwJh6RqAenvVDcS5pATIXsaci4SPMT2bHYyQ6kRd4h3U4gGoPPVhgTCRiiexNSZ3D8rlgZvaT/q
77ky6NRpAS/lkF5q9eUu9lCghfQKPumneAy8OWF1fNzYGmdtk71IysutwTr62qpVGZGTV1d9ujiQ
javHLAwu5HK9w/R61ORgQ5a5TBnDRdvKzrSgNNNHavOjL6mCPLzFrjqVrSyTb4lNhXsUFFn/tLuY
rMFR7dT8en938eyP1wdT37ma22Et9yiwiGYK5x2oPE4QfeRGIZqLdKzioO5KAvvfFkNIStu9s0JI
4GZQQhi4A7q7k71CgYCZkZgvTqpDWhxzg6zh+qx7WuUr47XxeXF9kdHTGJmI3IgdlWGe+0SO3G+T
p+BDErAQK4l5RMzu7yldLUzUD8PI2VoMWfRqs86H5ZrCrath55EH2kDZipVaXN66NH/IjH02ibIa
AaKcysLXjyZyoySrz8geWWrzTBd98YPT1FYFaqFfirTMZ79AdehkYhdO4J0Qeqx5pwGcE8q6tn/5
qNdP0mTe3V/cZG/uDUJfh6dNuxbXxZVtXlvRyhced/uiGBDY0mPXyNtFNEJuLfRrYjG6C4aZvaS3
MzfZKYaml1F2GDncTfU6+/4HA1lCdzCVAgaFBfI51bsnz0ZuRrd/yX4QgAbNahYOsI4M5WVvK022
cALFR542FQ2VXgpHI6YmqeZ4Y6WyWVTGZ5LyOHajOr/1/uEIWb0b9rCUuLIAC/vdjgcgxMRoXNHJ
vrhLYvFJM1eeLtPk9qnRRh8dNqZffJh3gjJzDe2zBBCf3GE1U50ngfaWPIEC8bCekadh/WAlNAo+
XG+P+UHLDDIlmjYepeYFBAl7EKvHTe2PENuzL4hohXTegKUfJ6VLpDF7oC4B1V935PgiujgS/38O
9LKa25qxEuMAEmgYGDeYoG9Nc4nLXLMLAZfMn8mfL417tWMyYXDF9s4dv8BSJ+onmSZs0X9qIifQ
6obVRWOQNzlZ1Rdqh8Mw/AgfDBxIWQ9/HzTLw9FVxOjfn1PKGALYhIl0HqG423VaRiLvJXmIxkDN
6OTyEwPeLjsNYLArWs1j9lD7wDIWwiKuTz9mwLczfigf+RavTrgF00ZG5f/nScTb7Xj4xnrewd3Z
p7v67lcfJMo5RouQzvO0LonvSsXBKhEF8OiTsySDnsG9PDsn2LvlBkNTDsM8+b4E/xyXX6Tm6pNv
bWRXkgbod2RttbDmOoO/YKUHk5zLwJT5ynwegng7TUbi3ShwqsJMJeV1ieKZiZN78qstjfMExaIF
kNSqYoyXivOvQ1KYE9B6E1Cge5TrlGMunIAJuTRyegk3t6RhtqHCaUfPyGonSSJEBFgNHwH9Z9E1
Fm1e/oebva+hkF6EfRcErv6+ADmOt5lizwcIqYbsOClnPNdApZzfBQKcuQlqoYHrW/p/8uKygEpt
4EmBlqQlZP35Rwxw8SAVhEoE+1ZRNw3ke4rK28SEKm5AExRRY64uzy0Hx6imYiICmpR8lXtyPIdg
dKYRiEglR7muqWHWOZCyZXxwe2IcoBCEPRXc+o7HvN8BqmNtL9BU9+4XNlHKwtbQf1e1q2yv4JfG
cd5CfhcJwFmULQL7jl+viNLAHn/4MsQYb9U4igmbR5Y1r3G6nBFmgU6X5OTgZmqdzs6vo/uuw1g4
AFUDiFx5GgoUoq55bIfTLMCtmum6e0+XBTj+aqoP49sBVZctTpfTnxp3VQ031dKoxwe2TOTuHqIE
lRzW+mbbRG3HDVHJ4aK/ZKXo1ztlCIDPAbPHtPxzhe48V/xiMNaHGsB4JK78VKfzQBGy/5j0fBQU
UyApjBkxprvWSNc80YQC0xNwu71ZY7BlcUNiryRRiLZ8dMX72TXEpg3CLGTIks4J7w5qJrmHQ7JI
0n/U9Dq6gWmj95l0JWo1DqfMRsbzW8jbB2KvmHt1i0grRxGJB1zxlkH3wo1XrPtUceoEqvTMXLJk
dzM1YVhkGTCXqqXA+R4nUzOQ2FnIYnvWSvT86JGio3J6n3QJ2Udc6s45mf1eslVtBO+tynyKa8wK
lUAZ43cASundufLDhQURW4TWDpGd2mxXMu42BIEuBWHVgN+hiG+SIkMBJXCgcsltsEmNe6ivPYvI
7JUmAcQxOSjaWyTcoJd0k8/d6WINtklvBjatXQ9bTFbTP2coQOi+zWY42vc8/w5wmml8Zoe+8+fB
roqlFlBzYwSTyxKCu8CbyawQOsvjYlnWoYqw3N1wPjssTQMzeXGeMJUz3BhIPcKc2Ly84GN2AIbr
4XGfC7X+8grC3YE+/qKFNhmb3JdmAb170Ulr4tXORrJVlqrh7EJHKVDGdUBI/e5ZJVJQ7wHjNxOu
wJ49NrJFFEFu5W+1c4y8a2SNYMEh6GSu4NEUwJZrSDOu8FX+58fFFMO7VdrYXEdhfMSaHHSKwY2s
sucfwCOwHnprr4pmsborgmu+L1QO1To3DmflqntiKh/aK4lu7PNthR+UW1qs++Cw1gNxUV7xQI6l
YxTouMpcJnESZZ53C6fH17E4ONfcqb1mw/hwk0ICLEs8dAKS5cRCVJ0Qnw6TnlXs7q9gCY8JBSaG
il4g2auezAJZ0xpjyUp7dl5Yzyv0faOSy+ONerPCG9Aik2/6Jg0Y1xQZK22/27xJMJGMhzoasW5+
Wk19rmBeT9UbvHe2JhPtC7jOZ/NNX+XUriEaX3pYdEl/RLFqCjBSGUUEMt34jKcehqWk4tqiLIDZ
9HMxjAJtBBKmrr6fXEtiC5CqJV0rgTPm2msUwPf7APLcgCQZC1yK5+LpvNk9yZIblde02JaB3HSb
NFvAYstepbksQR7nXEj5x97vqT5+tV/30zvjg6Pp3uMFpFTc7tZreD0ROEAKbhSGp+6fbi5MIS1y
4UNx05GQFzybQ5H8DYhFX71ARzZCV9fXeLBMTKra+Y32EQ6SABSUis0J5j6UrHSYj2s3x8JkVxop
5zaqAXz44R2f+ZeWuScnsd1YRIGpgHowFj2B//ChgnsEQpvEF58UPgJnOv03RumtBkE1M0QUzN2k
lQt6s8UEvvXXYEYnsgoX6ZzQViI2maVakVHIKLlX1pfzOeyVkM9x8sO3tYnSnuSI0NTEOhT7hnvO
JvSvfJXEC1XFKDdTKFZjDe2hsIIREfxXhA47imbwPPe0FYxgsttjpobnLtrlbgwm7QuJ6Wz4XNhA
vGNwunVXYmx9H+XFf93tPOloXcmSX4clnHlo15PJI5CT8GCoQF1Fok/Oj3vRais0qKn1mjig009E
XR51IxP7VV5WHwgbUVhIZTNa4XqSxtY1hxEafjU4pssnuOQ68ciE1Uf1kaeJTpHs3uBDPHPEnwpY
vzpx29V9UJvi+kactACtTlJ5SmrFdwtLMEO8bn/tm6I2lCpjP+ACmuKsiekbmpmgz+kAmscvCBI/
wPEOWTt05L5b1zpXMGRsHhdNZGH8aXc4m0Xe/FHEBxQxIGRNZlGqJYXeBZgrXMm/rVHUQjdF6lGu
23IIBoE1/qc8Ykkx2SRoxnXGGVXHEcFSyrKi27u8+K8BtwTSXdoOD+thstgNMJVFNzy2S26SKqbr
BMkFuHrRGvtZ+fpoWWB6O4gWFgeN8GVuzUPUZtyvoDtrqLO96kwK/vCvSbHDTGvP3/1uh3R3GJpR
pai5/hq7zndLB0NOgq9UMza8Ph0AeBYemBb80T6JXy7+1/65ZZqr4tqeOSgaBn84PB1388lJuRsz
bdx60z2WYDI68T7smLNjVbLUeLhYqDpHwlbaoPYmy5dhtVuoIgsRxXYJ7GCPRVRNdK1E9F6XWjqB
3a9fLT5oSku8Umx+fJb4kIrje451WFPlEFxhlrbOSUF/959Sn53a8tmsIrOSJWQOUY/SwYKzjalQ
u9lnqfyltNtNf8qrzfnqKu/su6V1fcyzZrS9oxdCMCbXHdH3a+NLpZUjqV2O9pDdr0EfM6v1BNdT
DQ1DZ27VWoJlFXGf8E6vBVcO2ihl0Fg6E4LkeSGhvq6ohEIxRwg7EwV9yqKNkMK/LVRlO6zo2rR4
iW8w0Y+0GKC9F8ziJpBNjpC8WoGuxaIoP0y7dMz/+CnYYeVlvi3uYQU169ho8CydIP8kNg8wfzPv
Ljgcir9IXtmlqKFcgMzR/nadXY+tGopSWruwvoLgspnPjW89U5iUbPj5HxJX/xQRFXLcm50+6c6W
tt696f+/4wV+bknZxmOye67uT8f+IvnvtyPoP+tEBaMCl1DjzyJKUpZP5s9zCmRlig3QN2TQluSq
BbL6TajKbhTd7dMCORAAH9ss2wKyZputlxElhwK+0FFpTfVOa7wX8u300xxZwgXHuUZpqH+p4fMQ
IwcHflc1lj4T5HKopb2Fiq9+4NaSIJBF7eokzd3cYerD1pw8w/NzOHB1YXqf5l/FkWyypIJS7cx5
i2qODLl7GzSGNzoOim6W3NsfN96oD95qRBB5WI/UU23M5rAgM0432G0jQW3CXu+D5ynKUo3UiAO1
Qxs3UTxxA7HYoc8a/ct4x/JoP8LCICVS029bToQFZ4SVxdAhtCg4O7vGJy0IveoYIPxBMwCtdKf6
og9sIjsGEJKmjGw0wPUpVYnSORIFbjYXV8wdHL1oGkONJTxgvsthOQN/cYsJQ0KE7GJkaTbZ+Cmn
1EpDBUrswRPOkI30emPTBo/RnT4s+48StpkI1D7aS6mKIwm+MNo9i9u77Ogkq0H0jTP1TLvaWK2W
0dgUtJmeTpR82HBU2aQhMf5J3OiBBENIHHiJjiO/eYfcd8D9gV9D6hTNY5IdDH/h328YUxcIn3z5
n4cqE+MQbARhQwDyeAIL0h6qBGQTjtSLaCjPbIo3a232uZWlzBDkjfO7w5vuqcWsG0TO+AkG1rux
DpB8oEGuej6qmDmmKxMSWTJHNTE1guFH/TcM0rBCQQoL9ryw8LqKuxrM7J84zecpnR5mQZP9lvKr
2Io+dBK7mj8A88IOWUEMI9qcWoSd2B70sNTw4X9m2brAR1ICnZJxsfcGLIoojYpgdUpwzYTR5tRf
sHBM3EAOZHjv7fDC1AfpRt/7WJcBwf7gC2VMm9iQb2x4U6bvNo/AYqfjecfipB1I6m0+pzH5Z5Ld
iAIG11WjWBZx5hGSlBTtBy/kCH8vqwXpnYGrfVZPabDtxHCQZSsbjPaeCVziHOy4sU6ETw8bxGwo
z3PjfQIWqhbRV016mcO1WD2kk6EsrB+zZ+2LqtfzOkQO3yth0CHRpV8bZQLXD7AzEbeiNRvwCcek
8yWZncBR5PGYKY5ZtfGV43yjLOtB85RyuXZDpvUUbkYZKBJkhgM+ujbODBjHIhb3uAYgn7yi3RP5
4fcpHRjcDaHOjyqA978u+grQXtN52vUPdF8Dn5D92zS81VLJeFZGbYJ65MqZ1OIeD69dmPmm4NUO
o/h+tAx8D+d/g0ow28VaSqigDYv0Yq6lrEyBe93gQzowaatxze2DLf0V4+JGoAsYKDKYXM+JJ/Kx
6+rmUlpeeTapx6PKEcx6YjziG0xRAHnx70QaN0tZqpBPOkR/J5ZMYJS+vIng8RdvngvYNIgS+ii/
CSML/RI763tjFEpR/x8JrROZ3+A4c8GW31ZS2BPBLV1BYWKXfD4DEminu6w/GjQNyLmaQVOeuqBY
ovctUNuNwfOPSVxtGWyT+gHMO7Cb5R3RUy6WLzPYEOX7qeewYfl9OZA7NGX+lLkCijnt6CX2rnpQ
4NnyMe7Gt6VGYG6WUEy4KFWBsXUYei30nrtbJkzVnjquZAvcrvXmU3zGYTl24moCEHRdKiFJMi3k
m035OSsYDHf8apeVdBra+Cjou2VwF/uW4DMaH28SyO1qGE++hkp7hWPpsDAV2c2SMfI1hSI7aW5z
F6hBegyi4EU6LqkKz1UqvW2KV8MKFYrgle3UQJx+RpcDd44f4kWcXFnqOYBUctmhWVB39hDeq2UR
lph+LlyTBPD75FG8lPlHlrmb0+JvPsm2d4PPIf17uYUxOIBzZVIDEMvo8ORfJ0fr74JujLPgJ0px
PWaqeul34DTf3BDMShv3PCvhyzarxZ5kZFAcHsTo9JPOry67Lpm39NGdQgqL4TyphIcdzanJ4CwY
OXT2XZsUN6HgQv3uNM1+vBYBMPCIm9+/B2tt2P/TAvpTmrKKrC86Xn5NcYFdyqtx1dbqTxp3CxIM
o8KDLKAB2bA9+EHIXljhtT6OYmou3oIm7WsZBBlXwCW+Yyo5WWMUpj4sqkypWx335JYHpF+8u4xz
FwZ/HvCDuMKVIJwy+YQ9bLsxeTz0dOlf7EqBDZOiq5PxVCS7qLCJm+3ab04Zm8yTVwqg+VdJtJ1K
UtJtC+7qqbbtgJ8jkedIJw1R16r2eTe7VtAybhy3vqgbV2DIf/veaOvyfMKnRn58VG7M4BETk0xw
/B5EE029GV/uqDL8lQfyLp937HXHX3sQRIk/33VqaA22/fSCjuv2NPaxezz4ZBAN8PEUpIBm08so
8crVT4Mcv9O/11apKt6TfNWZUI3EXDRNsHOlBtH/VrAQMwKUvBcd6UPO1nlM39rozZzqZp+nSuGv
sSCk0HX8nz4ocnIT7fD2QDzWP1zkDNKeXbZLhSYzglVylQnRsQMjLbcirA0aSepp2rqcMBWkXNcy
jXjtzQLb5I3vvpn1arSYdO5kUF/nPpsIgBo+JnV4JCtYFbo2XLSzeYKiSSOJsko8QPqSXHO2ZmtM
l3dIxMrFt9LzSXQxaOyriHb6Hzu3sa+JNCP0B325PLZ6CKDn4jkoi9tsGBHkPKyHg5s/m0iVD/oZ
br1o8Aoq4N6iC6oKzCyMlLRSFmd4KhgkJ4FXlz9gxy6qYUQJh+TokhvR6tk5FACesg2qjDB4qPnI
wpYQRcd39HQwBNY7QrejeoSsNtXg7HOZV97IuVxt5L2XyRH1LH9ZQowRIZMUiKgqZ7QO1vUzk1BP
+cIR82TaNS8FbKJG5fuMjINlb970bwmWAZxlpbWfgMWoMHLigQnw0wyTXco+Xn4I5G/nLyTh3Cuj
Btky3DbQbWib69nxVumlUg4KfJkO9azIS7Cpt16KVWhgrsCbUqTLzWdep6LMvmRIs/RIFpkhjl7C
UJ+uuRX8qMm/QeYMzvjMqQGpL+9m5+GEZMy9C/Gu2q5Edx1vKGDrGxs8fzK8zY2qItoyY2acERPx
kPDSQdwdXswqGKus+PF2M6Xov+C1Er3fCV+pQLFfLkqJa2yaK2cmbCPd6X1CBhO0AK2TId+WMDfT
KAwVPC7vwbEpEYMBbCmb+LPW72bCDFnI/B/A+p1QY3tQvywzg3e8EEx2rq0HLtH1imyLtGOwiqFn
TbTg7Szqh0psAexsXXFSxplwLlVhh/2NaNblg2MgitGAgfcNf9bRz3iU5n9Sb797kQDDs4S7xs/M
T0MdMtwgHnwr+5gcrCM0HEzyMW2WdraSynJoCZ379XSXj8h/mFIe0qZBFIXOFsSjzNFcL4orbeUV
kynK1ZdVUAylyzX1uyL/POIiV/dRQlC/0OVDSGIyZ4zCa/egJtF2Na/coMLGcIJTAFyGYVWhph5Q
uHbudR/3/DuayksBECod8H6YcaV9qQ6aRjgB5/OCSXuL4QKim79S2Y2PMbF5RFDbGALNc4jHGXyz
Q6MMRQYo8GMME2MqMQnh7T98X4xtzFqF9zn6j/neR5PRua2tbS4UoFdNIGo/w9AuYMAQ6gNqjOaJ
JGKY5LI8v3owUF9kAY2aCaMBrQ/4AGb+xk1B3jI469E+cJpul7AB+sR33BIjfasf83NvKW6ft3rD
do9vgHmbanknh53J8egd3jFJ+2gQS8WTabgUh8tt5tH6hBUF0WVkzMmSgeYLiZoh8j+iTt7q1+Ry
N+lTkJi3e5tQXJJd2OfCZSfJejUOADydZJP4LzCZqf3E0G97yrlmWe9cTMwcjfJihJ1JFhtN25Db
c02DN2gjc+9qStW03wjcHtNPONbthmf+JFDJYjioLDEqvg+rUdC7tqg5sVPjDmfyhk9Sdw+bjGv1
nf5TjCP/SapXs/IeCx+n4+kk19COYZIEkfdQ7+64xitRJrF3Zb2AUlr4U9bo6DC8gOq1GZ5InSO6
DJUhUMxXwxOCQPlHcbKj8y1u12CPpI6puvhyQchn4WaW+zoD/q3itOUK6Wa+kypWDdfQrescXxVF
TFJXm8XKPyWVWH6LH7m4J4S/f68EUun1pQ4U0saw2wc04dE4GI34lIUaXpAYzHyxOn+jnmYIEDjM
KCib3neHK3TDPF+6oTK7z6n5EOlhYJ4hPLtwVCO6+hl/fq+owxfbDXhkn6hJf7rk+QwgMI+GMmS8
/HsybH8aZZVqqui/6TZzSwarA5derjYxVmsic1e6qV+KkDlYIGARccaqKW+aWUGCQ6QRxn15J5ms
6HwW8VO52aUg4c+MBddQYLf0mdp23AeNY0g03llrHxz1iNhX6DeLsHVS+AN0sNysyIDe1eXuqMWq
CO3eS9v4yML4ZuEggN+EwK3pWXvRFRlOQmsRfi0S79ztGVJIGA7GVmbFsJ/HbwwWM810zTDLqB24
tdI6eFaqKICN1QtXNjX+FV94XBq2D1q4zcYLfFUZQMIHLI5DFopYdo9xqURrabDwQwz9KbyOEGSh
h8a9OyPSm3Hf2twVv2PWDM2zF99pirQUYa6nWBYq2yEinzsf7MOqKooMMp13VGiapJJjts30hovp
NFdZS83/WTvTi+yeguC+w4MQ5D4lvQisqrReOKYMSKLNV0/HzqZ98bVtJtY5PecIRjH6YJsQWwHw
eH6Sls/4RCaumn6KVUqEymPg2hFSaZhTPQHuay0YR97gBg/mdkhpG3ZU0/cin1wZFOWZpcCYbx4Y
v+DJxw3Jh/+GN0TuKLgjh32Udj1Ergc294/scbF8axiXlJoR5X3jY3lTMz58+zsWRNckxofXQ5k+
fC9VJhHoCd/Q6cUEcDEsBegjL4tCXHrUT2I8HuBt15pgZQqumaKdT+0a0QLybqNVZc6iqiJZEotJ
DmvgaHGeUaDqQ6Mk+WWfXbnV4/oRh8FtKrNeOgd98ltTsZf/mvfjCJKa2TpFIdnlkso2AkbcHcCg
ovyWn/4vsY/MzofH8YwX3l0DbBeM7NaBngtD9tbQK7aNqcvT5O2eaR7kCweHhzsPBmzjXL0mvsWK
A+Tre6QQax3RNikkfvKN7EuRyU9M6U1TLNxf/WMUN5YKZsLzzVYs21RrnUmv6sP+1qugOVWSmrwq
4XWjO1U1ftSRmOJhCMbwDrcrsa+4dxOCYOPWf77OP9QA4cUdPKOT6zD+LyrjV/YQbBdqlvihZLub
gBWbWz0x4hWooUgJkUhWhwPghRvTHx3X3/DfZM/YR3VUSVpNkUT5QggqGGxLGWnHA/LPlCkhSP+R
cduG3kGhcuRze8k0MweViQGQAdFa6Vdk9aR/nk9btqWcbUjUOG9NwSdbzYpoC3oYVTptEmCSZMbr
kvBB7uEF1551Q69VoNebg/x7fS6ZP3Zg+J8j6Qvsx6pH6lgZolLjCmbTX7U3jhbp5C0RUrUPDHCu
KaAbkGb+GSIt7DhZnq2V2eaBybXOTEMJZX9uicVpVBZfSKl04JbP4ujsS6ZSPJpbCz4IlDTsGsYy
TlC3+E6ovKjO/ZtjLFm7y2Hp0n4bSwlBk/CZXHXn5q6YWoJaqVJOgCrqLGu7IcQReLhEh4ejPZ85
/plMRUfakWnCbGulLyg9FsCqO7qfLJSzlyGvtFECLm25Yn99ATc75kKZUzzY/gHOwHCqX6krbeoY
mFBdcSm4PT82d4vX+iixSgfqVxw2gzGGqLZzVkOjUx2NowUBBbx8vvTmlQMdrbMH38/fownrf/fM
42CCKIWDivt7xlZiqNBReD4TU4FEuugmDKOAWYucNrebmLVgT8Z8gcb1IHhLeZAS7ez/vx0MxbFM
ihLrQ+b+icttCAENlSqW4Z8kfyjFY8VnO6unMNdswm6U19U7rq8/0y77yogyOWrjBF/6MAQZ+qtg
Sc/R818DrLjPswLRmRu5BdkLUo6rWJiE5s0tpuvvdSeWCpomvlnlLNcmJhRkyNEyusOTUmd0UABk
UxqHlR88H99dbFYCa5gU8R4bX5LBnGWLAPLwsiI1eA4FUYSLzo/BV5HsITo8qDfG1YP4hY4Ac5uE
ptdTjOdfy/vordiNaxgQSJ2wnt1AEApfFYeh9K5EXM2fcw/ubSeTS12BeX46X68l1sh96XR/trBk
AqvJDo+lLZo7HPP5uWt1EcOUJUIe3Zd9R6KguyJPnI3Uaxc/p78INa/SLX+zrKWq+wJNfI4PY/tT
3UwyFWPfJYkhQqRIsLlizgnJBQk0rLPlGGxtu1vENcE6JftqC2eUBftiAtlfnnCAj8lGyIl7DUzy
jB9HpFjY9jzba2aJ5hkLlBL4POTwLNLK8xJ7ilOYf3Lfb2EoaHGMQmDqOKAXTzfTH/GQJ8JvCWTQ
jwnQCYghnSwfpaewAVBh+0PTgyjf8GoulkMTNbXoyN/tVDiIInUj4gq6/xMXy+gTSZkqve6KXBnJ
kB++LS5KLvuS+3epqtfiVCs9RVBOpzYNP2a9SdhKNBqvO8ss0rNv+E/PzkzitmyoQivVcDv486if
3Ysd/XCUEe2XL9GAzusMAuzIuK8N84N6qug66iyUqI/DbkuWDyXG1b8zOM8zIcNr0w39EqNA+YP3
q7w2jaAiK/VCXw/gkwGz2eJHgyCHBJiBpOzGasRLMqwJWmPkjE2rtfr3t+1YAW25i4I5yexfNubb
JXvFQw6KrGi+DJRdjpRUpwTWnu57pX5H1cOa8sE+491eRfW8QpOTp1qd1Jbli/E/F+H8JParLInm
vcytPH2wQk3ARj+lHs4bsc+ZqPBZcJKK2i0Wp/fpc6VNnq/w4gbzmS2HlESX1j68Eisa1Q1TPmIt
+1paCEvcrwGb9fHuSjoScLzZsP0Xo38lYVjGJnd89yD/rcvu9HDl1NSzWZe7BlaZMr3wqHI/WSn/
jyOcAckKrAc1kjITSfs7ra2/3PO63adCnINV07j+SmYYpJT8CiICIb1kVV2G5O6p1VZPlOok0DJz
zPkdkRMe4cmsOmuwdzFJqgPwRT06bHtdS8z8u80EhstpEkPk3r+fG1qfH+vN50jekp50PkZhlPoI
aGw5up9ufaZGcfsefq4G3YOxPxIpALU+Xm2gTBOIS5r9TGZiORJtHU7gfPR8hZfK28AVhQZD5046
WdOn8JFQErTgto9gkGwKug+AZu4eELYmxFAjDRaJPXnxr1oIGjyLcEQIl1Ie0f/rHaYZ7g0PlJxz
TBQHdDwSyCCW9K6z0/552wgeB5A1I7cdMYFm/bYl9IL8dgd5RHS5WxnuvSxQLJHhPf7Unna8/c8u
S05oINTgSGmzWYyS8OhH5bhmAPhab2O81LraELFm+W69d5ziEJnAbsGU13sxEg/P7yEm1BcdO0Oi
0Y7Xvy6RBCOSaz9/vMW56LRt4iarto7nHyCNOY/1459dxV4Q/6SW1iqmB1Vybgjicn+NJKPgCrk9
CAyGgeHhzKSbFG9N83eHbghgOvghwxbWzDosbkdm0qquNT/3DF1AS4fZfDlmfeqNaBN8fiI/bYxr
PNWx6wRbVDU1KC2O75SVa8OdspIvMiGSrrMHimnfzxxj+MD3m/D9wV93TvE7cirg2G1nge5fMv8C
wgguOQ6VA7KGjfNHr0M5W5kbbTn0QqsK6+ZHmSC/1+w/9lzzdNdyDWtqGhvS8rQ4UKd9hGAN/+KJ
8dKAxJqVRP9o7XDEHIbcPBPCO6tvFXModlAGYGeW463EXF7JKRmnLw3PugxzG4gydtva3GusjX8o
h49je4e3JkgiS7U5mcFOKGjV96DTn5a8fybwpMinqsZ1djRslVJLT9epZvz4yXBTWWXg2RbmyCu6
Iu0fcGVBIK00MKH8B54L5bz6vhpvaGt2oU0IzVIuyVHChL0i1UXjwXdAKFv+4SI92jtRaZPZcgYZ
RUtK3RR9pqUvg1NDFCFVK5CnPKE4rjITuQAy8H58CJIxEUPr0YrvAMNk2LEbV80xubWdBma8TnQa
UEomZan+P6ePyE+PBFInG7qoCNqvBrI/m4C0S8mWlmIS/YzI5iQ1QXMt5rBVnbSJhAUB9Kk7cjGY
wLtujbzmWMImLuromj/lSc7TIxSur8s6egBzk/eeQusll5uCziJHRNw9qgrBWw5DtDDffnpeqWHV
y4YleEuYHiOG8TjD3WwV+M375/LDV4wYTMUDz1wJtw7i/hwftnFE0q70rGC6fm1RfXTr3YHwHQ1u
9CNqag0/UFbK3UUfWUnUPYF7tebIrShwUjZ2y5kq6KJXaNDospaZsums61cPARKvSrFKnhejT5MH
c1W+UqV1mhmZkACcv+NjvOB8dTF1zyyoSe8jw2abfujE+5FAg96havih9xkKNouz+YFX/1o4J+Bg
ai6+xpOgpP75LT3sL6TCfOmBcmVd5arZliq80kjpdsBp1VqkEw7aTW2uTfpkWQF1yEToA52neRSA
uFrIG4H2XfZdFZ6YgCdluWHlRzHuyUEp64KVgVJEgGVLY1dzRxaNM04xZH424Lom2nTr4HjRnKwL
BQ8Tyi8hTHV7efPOvXxk0oORMzCJY/kiIYT1i/feVetWQG0ewqOFItRrTsnZTXwnR6z8Q9PySpAF
ZC7/D6F9OjP2qYrkkHd3ymLNLuK1wnhcdlKSn5HPrxqh4VvvygcANjkpQBUVYX+pnaik5zBY3m6L
uVatcQ2eaLWEEM2/WYBSq4UE7ONXal6PKye5yaLtnkfrFIJs2A2imQs+ljhDnRn7JGk69cmmvANk
z1FmJxr73mRmlaCJVKVawltfV6pTXijqTgmBRdO+CryFA/czaKMbjfweeQKluYeLdHSAYt5aX76j
OYabuqPgm+pxP1ovVslJBIrZo5JJmuXvbfc3/X7ZqmwVGmESq7UYtIR5kFN0nyqAeHEhwBYbwruS
UuWQEzcB1I46oBDGUFAkzlLXwKEllnf07aXaFa5H8ZktDTlKpmk7sFzFGeihHSd2RpI1Q14Yr7HW
JSlcnIHA00UaQO1/sSE2fJ8WL79GlLzFABfqjCXVUujY9xVDB+TB0ZPyLIE+kXaa9cinJCfPuclX
BcB0PjHnm5P4ELOOfllEyCw7j2WBTRq+67gCpZ1ZzT8VIvcalf4SAPZ0sy1hYLpv5LcG6OQtCOwy
/1gaQ7s6ITvz0hXOxORB0TxVirjtEJwEWEE9jqmIbKhNSAiVfUp65r2XNZ2tTQjsRztUy75YzuLA
nBgoAyxTiAK1TEdOeytRjb5Rer1TXtvpEtLz/Zp+APDf0550be6mjfGkdQHKS/+pUAFdY4M0zH7w
+tlVN2fnfN1OuiZPIfQxhlAdX+W8YdpVvC9/QOHWEqO1/Zupsw45KGhbXOfOXb3dzSfk7T/pd554
pKRTGzxBBmgmGg7JZho6BEZYyV7wl20FgHB7tk/9RDkvlrKWVKIkNrrXZ/cfg92NTYx6lFRgR1IZ
rYv+sjBO4aX9/0y6z6e23twWWF++QAmr/k4qk7Hp4jbghwilmV8wB3lMnVOuJUqIjBD/d9BS+e8l
/C9EW3rn9mgRG99istKM/8sOdy1auJK4laVR7v0Y+tKsDNbDRydyD1/34kiNHmpixk1YTXSpl9+P
Ju0CNluSXYstR1TC9NPSk9RuNB+JNbL31PF1jc5kqpW0BitL569BM6nsqbDXoNBx9mM/pyg90Vq4
dnSFKnpH5YN9K3JNjmFLEKf0rlfDdGT+9TBEAbj6HgjYiOOFEKB0asHeXWGfNOhR/6Iy5ht4DCr4
DgXCupsWjjLiC2oUJ8ZqyDzqIhwRbLOtgAJ91E3yB8f34AnO6ooKxsb7mChK7iE7JOXq34AgYrbb
6PoAJaYJGrDFgqUSqDdp+5AA9oj/m1xxURLBQm7OyB91X4li8ckJELGKPft5oj1vBa4rnRtODnIc
dg39M77g9aIPYsb0z0qcF5ss4ffN2L9pD2gDx2lvZ2Dm1bW0PUzOvsqA2f0eQlNqryU8kiSWLSiq
WvP5c8Kx30klznZa9hCLxpx/JJqAB/6LkP4FSs2vp5nONoOWZ0b7EWT9dLAtQxpbHUVnt2s4Bmam
zcQTaqAyqUHkDtYd33VIIfUpNYsoNjRz0HontehF1dCovaUaKdzrlH6SximXK3pR6Vnto3ku2PtJ
4DVUzZ1E4vO6BJdlLRm1Sf2Ao/KKushcx8Q5HIkqBk+cQxBkqQDgrwM2sH3ehyMuic2/EWvJvCJl
UVtvg766blcPPbOb4sgNuSoYRrQUuiqX6nCDm/lXNZ40mB7DVR+sRXEUd27gDpTvRQrKqZx/fw9k
IGQOJMNRZsrGc0zqjqelk/qjme7ZR8I0lIjHxpUh8FHco8UyBpBH5sWnir5i/TJLC0G0QxjBJfTB
mnHdOnNOyf64I16PBRlyK57kFRFHWCgVqjDXRakUYC1sry0P2UcxKfHok7yKJ2GjIOt/qPcMsZ83
SQnh3CwnQvN8NkeHdYmmasMJhU5VJGtd1BfeSqsnvWfzRdJc+gBEQY+eqRLwF8l7+zyHdi/1fbaP
h0q7l3+oagszSsh7aWQCsZjxoi+2SiuQrNqBlq245qsitebVMLOQ37QPrsTrqN6LTSuoBW/JkJ6Y
CpGx8W8P/FJyA15gVxD6usoPpgOEIya3SBrffUvRWu660mzOedbcWWIHtjlaLrlwEA94ucZBH7DN
/zZrCTGPUE3TVr0jc+96+8Eueli58tu5YAdoySQMrKKrq9/jQSUzu8r8VNrltfoHVfdjc5ly2Z+Z
nQOwSIiOGVISJJYGzQnsjHFB+wl7+JML0XGYnhj7IiOlMDz0pQqjPtj7kKuaaljUBgb2pwLHxmIA
5uumSrWtMxIOHMb0uyFMAPqEdJjY1S7pAv3FnmVvJd+hcfZGBbOQLO4sLeRPhFRAvd1NYtsnUk6N
7m/0ONr51/lMCLXAvq7Qpk+Z66zYHl2CC5B13+dniV/TRh902RUz1eguwQ1nuYsihyP/X/YQ+Or6
iUDqU9sBL0zRpsYKU42TPX+JJtzlMYbgdShK+I21WP47JLtwsSuUm9qbjOCUlcyRHoCvCTATD/Ay
zpGf8ikOO2e0gNeNXlDZSJRuzTgJu9PSwDVWhzxDH22eh022Q1Xb/aB7Ahb7RHQ0rObqICWGeWO0
SYqbqWmXGScfVdxm6kHDYP1zrgKF78oYorNGZJ7NzTMjKm+N6BHELQ/cldHM0FS0YGNjQknoctIZ
SQdO7A0YPB2w1mDknhO+jxxUBoXnRLEkFLvsJUVNdWt5OyErMyVJW/2LkbxS62s+GN6FLie8j+C8
CU71taBgGBpfuXgc5PLw9z6xavU19e+tLPDKafsr83FdiNL2Be2+QCapJuVNNRBaCbmHQUq1eceb
YE56gv0J/HkH3iWF2iLnjEwJyg1bWDmH1eicz1PDpX4pm7j2QPIWufy7Qoc+3/6jKAzunlwnucAq
Ctysc/4qGPGSOcq+Zv+Vdu5oK0mVEltfJ5dm8/Sgfy+k4WafDNy42fOTmTRPud3a95xJCjM73+3y
k1G8mT7OnRgDuEIXhcP3gH6JajB4etwh1vPQewmzptFzJMt8iC+IXgGxU9kSFx+Lyuhxb1ZanSeu
hxmdYa0a+iBi2ZiiNvEQutCwYCmMRW42pkSL5XZ9vNG7Hbcx3dXJelL2sOJZvL0dOp3b/7VWlgn0
qHev6JYo67n4yVyzr+hkAA+SquzOpkQMFk1MkMusyohm4mlt+2O/4yHVUCbv5pcwDHatFbI+vEKs
QBRdiwjLQkz25BGVcnttjv2FZZT7QkTbReExnqI24XBixb/B1+wsHd1FgXiiZu63w2qI6EZzcmnX
+s5sPhWAj4xdg81ONfqqizR97y5/JBCc2fFhsg5Qeh/BhqD4fA7D472UIoSQwnm71bdu1EgRcYMi
M83JeXPi29lYs1kj+9aThcAGnjmIY13jQPPDNWzntAw7WPLH/qgpTheAgbxoejFArkH/GfVOX1X9
SfKnFiCvJwxYy9KBdxPxWKWz4pKFvmaYHh1p01atHMzZK5DURbH+JGgwLa8+sVBWIOqoQcIMQV3J
+ecxEf5bFufdVu7CH5XWuMVO8C38Sv6ZYNWgrv1ripQoVFv0M69kMWXVfikGim3dKwOxchLle8g1
gg5iNxgiDVV/D7vUV5sgpILsva08ydOyVuQQMevx1ZWv37q2s+rDPh1GqVJwIvr12U4hLM1pFSQP
y5mTMeqR9Q3h9hKwsPkD6FrUySDeRKeDw2PP4ZX9dhcvEat1UucH5atKZLJqkoj/O70Saa5ERuCr
TwRYVP4s+Bzx+NOW2KdJr9cqC9KqF9hEs1/PWcRZa2P7mGIyQvd679LNBiRj8LlXSbmLawYpKTqV
/x/fH0wi/m6HUv7TFVmLYHV1IsFBDnLjwYlNvZQfcJKtXAQnZZ3OlRonXWAhdC1AhI9Hh9NRhUxB
KybOS1cClzMHjERwADoD71AsQZZ562hvj7EzqsbvWpmXgThP2X2nWyEFYQNDLccK7OIPF4Qeunmr
0nikf8DEaT45jAQ8nLpoeMBiCVm7GwT3zc6doAdKiaIeD4jm4D5X3jKSqPOhgCUAHmFMh7BmkKl6
dHukSnbprj8tX9IC5ZMHaxraQLWxxiWN0moktyIQQnKHFSDefMz2BrHd9jH7tc+cl6dJIVZHLA4l
2WNsio1BnkrX/pbt4+ozPRE1YL9cvTn0Qe6RG/T5UGU7KobhRRh9t1oAuy6qLFRDhgTxrRte0rQ4
kwcs3xG5/vkloGb+WBY+Ay9D8khshPPP3TVlrRfJbzuSQBl1XJHhMuu9nK07y+W6tmKf+lHpgX9k
EWF1G6M8dACyYkNXilDwKwOyg8+wxMf//X2v5ywbU5FEUdnpG+JFdTHqOotIN7f7Cv51RGac0sED
0qAV0DSvKLSVPqaBwc9/vtL73l/9FTK64uY9kJG+U/80Wauo7CS5+4GKn4+XU+WyeiXM9wljsihG
U3qH8oe+Pj0G47/3ST76ulSp/WhsxoUeezJRrm2dmVkfzkLKQYxbY+JFSNuUIT6loE5GH94JRZoZ
Uafy0WzM4KBfXHxxFKvretKAl4hxsy9DAXEwSzm2Sl5iI17HLr/SqhAFghQxyCZm8qIVSGBnWFKl
NBkdT5Lny2IyWTYzTDscse4mjogDadL2WeYAxT6OYA9QY2rv7OSdV8mi4uMZO99kCrjb5vt1Rb7D
NA1o0PXMdr6y/sEvI0XQsLj6M3Om4HAizEokzJbIqaCyZyPyE+rkTzz/xz/g2NN1/LrE7mg6K13n
re5Z/m+6En9m0NrunSpTsFdt5uiXH5h7YOSg4M/DYtJ7p/Fty/PEk73lwqieQV/VxOFoi/06U3r7
vzcza4Doi8Zi69XyO0fDs/jjDTN+q7bTUXAfdTac+GGgA7H8lKC9/ylwuFACpkgBG8EtCUIGFVOX
yrc3Taw1gRcNwgnoBzYSNT7Opw41N/yEi3M+E8ueRihN5GQll8R9Bm6+CSvg2weWw63B+hEVin08
2jj9lRdn4frsVAQ+r1oAIsj4qhTxEwes1IqQ1RdPeiDKl9CQGyn92otOyh0nLn8Z9pYiJSpmViAo
yIQvczGkpa1pPq3HBtMVgR4b8u4y0qkih9SO+7OjV7ZuTMZTcnnMTRAAQvnNW1ff3kpXGfI76Uo9
O93OT+sjIUEaMtiCiwM42PVEYe3wEl7atQdhf478Vi7rOK5cUDcx60d4MOOQR++6nLJj2VZ69ICx
qkl2o3VYjwfjmQvKVTtOJeFShONXEvXqN2hIcJDcyKwgBFdFVDZmMZ6tq+VFiylF3BB7MrcqXE1D
aqJLgDGYRQNE+m5tnfutrbUnqnGQn8aX50LohUff9VAgTohlua5I/9SDpOVdfkjxtWwjUaZp+Rv4
qRKt7Api+EDJvc9y4VDUZU1so3tHo8OQCLvrFKNxSaPiKMV2JbweTM0pP944YaNkOlKfD3BtVTa8
x8PlTZTCbarWYzFR6DMlBxcQtWzrTFGD4j5XU8DxCOPIZq3uI5mADxgZbTXxoOuZLh5zjdpVrJwv
wBTSfeHtDyHofHYnQsAqf/GFq8vnWfB4lyU/O4AZKWxLtjMlo8BsN1na3gBGjVjpaaI1eveDQgIh
GZIrVFn24JRw3MWPg7xBaA65yNh1P2uuEEAaKTPWEUkNzgTEOsdI+7csmjNyZLHUGPtt5HWzmeRJ
WDKHNvecc800YW6vOFVe4xNSxHJYObnV8MeiGW9Su0eXoMIhBHlDnOvlFygI8S5zj1DD9G/uFYFO
17YW+McILoZA+7wi+Tt55MakWS0wE3V+lrepzzWg56l3/ILvfG5lvaDf6sBg3haGgneBpaTf1tUo
zRyURfk10XRJOPmr/8STKBkCOubnq60QAHsTsim7H3gDUXYuwpKKQ7KlVkfABpNFTCKRNL0O8MUy
G8Vsv1hQpz6vj+vsbHGliASecPlxEQ9d5jYQVJzCjmDM0J7yeau9OE2qOcYX2RAp1smpe+okPFa6
H/0h6MzNRymlwBxeztsEG+rSE4uOxYT016XL+NedVeYuXvTOPbYzI4Si1qhiLgkQAMHhTQ/8h3PI
tX6UfEmrpAkUen6UDPZF2gKUiCrEHue8Dk0oiVpYxVoVRfVDTrv1VujSeam19VALfdKdr42buWzV
NtnEa4AF9ZwQ9a3csmrA/Yd2Lfb0lSQdYWfzt7TACR4nNNHjWA9l5kQiTsQeudinSEEcs5+6lsXk
ai5cqhC9xUbfnWV6LfCEBI3+FM/YYAUSESR5T/T+vc9tDyqLmqmewAo2b67SPbK6U6k3UF2fX8X1
38Q3f4DF53JnIePT45GnnLMj570L8WwoVirLFpNWsZnaZynzTBWh6mntw2utPJulFbDF5jk6YRWs
UeRFeNuX9BQwfw2gVK1KuEgXOqzwMRKWjBsLl6LA8JaqBZa5wqwiBlju5yuusIzJLdBuwt0p+Qaq
9XraV8njfY7CHQlRl/bTI5jifPtW2WSISt+iO7jC5YJDDNJXLc8Z5xz/I17cLGO/N43o0hR+Npb1
U+LlbQ+D6mcVuIjABTcdnokunNftEbyqiX9m/Nzi9ylU8Z4eeiSWZSgbd3WiPF1HfFm2QR4CZsZQ
V1xHLzKM4erzyLmZkrAbHRpuGszvRKYzqNwQFeMeTwnlwcFmUn87onECz05wHU2cy8cOkqtfnQwW
IQfEuui6TCeI0secfPnS7WwChGSvZUs7gGe9gxU57OtF44Q55O4ZBhITSy3jdK6xgi72UGA7tCoj
5qpDltLmfqrb9JVLpIsqiG18WSQt6jwNUHLOXrxmm1MknBP/qmC3Qv6rfv7OBMIe96tfo5ZFWMRu
Pm/L3wdyjmEjH43IDFVVpwPhm5ZtSaGZE4H4YXJLpHVKZwejLGvirDUC4lmv1T0jLj0h48UiAwtA
VZp6upnHA3HOxCyFHA7d6WHL7vzqI8dEsHpfZACNvaBI0ySaDZqIzQhfsa700Vzc5YLmE94Sh5q7
Mi+b/m0pMKvNqYlF8zsjLs+bIXPJC7YlOSLfIwEGkOWtxmJSWQZvX4epQ4jx1Lsc0mWxY9vzdjvu
zNX+IWcQHc2FNVZp9xBlPGHD9hdivjS/3VB72JLIBYOHPU+kGlRF4ZjLSR5lKYxTx5jkT6oKSOhc
XyqFEJQ/ADmyEvjNSK3epdvQdunGJxbCSCa2gudRCtCz+6IKxTM+VzTuQQfc8vw/Q1gUvRW12ng4
KvDqinDyvuet3shLpq7Y4sJqKDg0MKnxnEJWKR+OCDztTUUjn/dKXT+lCbvDOc1RvERtalXT9cMJ
d/983G5/tz5HZcLsXPq0YxcZAsoEIaTL/0MpQIa0EvooClRK6BOmheVRNGxzL+S+4zcnXgFO+VmV
Xgzn0z6EqjixXmJgS01wKc485d7Vt8u45Ls7vzCVcHmzM0EiR+MAhnrkjpkq0U5r381BLIbDypTQ
pglFA/SAQ6iqkquPDo1T8gzt0dAZxczYV4kXAcuYgqIzN+dL/wvtRe1Xy1yLIiXftaoa1m14AHni
R8FWjPOq4a7CSOJxh5pAqmZ4Nxum1FZQQyPdmeUK7Ivx7iO6RsQMdoklm/6iFKgrHGnaUesQDsbb
t6t32VJ9SuX6DJgJS/dz4mcCSmtJ0J+aILcNOtSBRW8oq8+6tfm+u2z2dTo4HruSIKsPpWyVJbqN
7KCbgO85VWhb+xd7hgVOPZ9GG4pv0Y7oFlnVwXjOgk30AO62DZGgQ6/Rq7NIy28VxLe2WM6BvnRD
EczXX3R9LGGY1LoFoVjyInx7qccySel8tTeiBkTicxtUhLq+qIgORxecf+wWKGprXSNx6+6mxOej
aRiAcZdLab1Ku6LXp133aVeVk8T6nnj7e25cPzk5ndsOPr9EXWM4DmbX12XaOZDPeAhd1FUoJpbx
uNTca64ifKlAIbFoBysw9lwh88ipXjtpRh7kvp00HnxTjZItkFD8l3xKMPSFU9smzT7UKAPVZGib
7QIc4q3W3pdeeVJbv8SAtHgTcgoFcV6PbxK/0HqIAUL6oS+NF04opSU1CNQKZHIb69OSiv3++qKi
BwL17430G9xnKM8OzE1U4c6J9JK0wLB76Hcwt6lXXXRQag8Ocvv/ZISuQaOB/bSaxNLnXudMWtPJ
SqzaLGx3vLiWoDmax0Si8ydXO/kh9uQiE+12INfVOwfOjjKoEztcdMVdkjA9nQtzO6mjkD3+IwQ/
NxvdHKVu4/vRdqUmSccE6eJt+xDQ7WMY0mw/DyuGkRTHDWWhP295nFMFjg/nyoOEuH52RaYtb86b
IX8eoQb5/L8NtVuZH94TvEvaWFTr/YWaHkOzHGSix6huoE/dOvW30j2fp4on7jcW4kfksS0d/wx2
NYf4UNUY7+5R4gCCRoWFmBEzOtgdvBdrDqQkTw6nTA9HbaMprEAjJU+zHqtx7Bxex80lfWndjrYZ
LwZ8pv4x6R24F3H2PO1J/ZGe84Uhr5ySanj8N/Do+Aq3ObC2HlSXUhM9QD+/W4mmV9D4PDHATUXj
n0Mu0Ozr2hK1Q5bcKFO1xvsRWXRSeiXkergLVvM3daRAU/uMs55bRzBxKcgaX70CexRn3ZDvj1iT
uU6mOhpXso74t9d2WXQqk0zfDkKE7x7yTW4p5W34Mw0h5PfhlU275bUSJATlZ7nPKHLO862JMKq/
Q0v6Y7rkp4twDeZpl1xh8Ybe9ic8Y/TBOZIKhx4SBEmVWzIxS0VD/eft7oWuLGwc9rj8WhHQg3M2
X9G9IBn0ADrjXSxhfVNAyJc6onOlncJU32pGkZPvYAAo/AWF5y+jxQZZfP6HupXlg553hUopQbYd
J3/KBRbVoxaoHB6dVhcyIYnxvRRe8vRVswol62ZomV4pyCuuYep87WCYZipWeq91u8yYd90NL7ld
febQOcm/l9DwFxyalRi+ZCBSPvhSofcOVdFSb7tJTtRMjGzTTy5NqA4HsdFVKNgU/P7ctZUY/lwL
cdRDOmnUiE85zSyLdsMusifpIGe4P+KCZBc9r3abKPFNAFW3LJe1bXl6XFTpkHlfeAuUVQpe1Sgj
pYNrejbhQcrhUcEst60ZKifdmcnlce9X1nHw/iMzi4OQWveu4iMxuNyzO38xPFwE8kxjQQk3oEdB
Ddut71M+rOVFxV68+sjDD1ouQSIN/uCBa0JY6rkaQU9RCsxXQ3baOAB5/Jc1mN/uLX4txQ19FEw1
RvrYDSlF5q/zlGS+M2X/Ji4gB09y71EEF4/8oHHhReetyCnKBAztrVpOF7ZWhquNCEe40m42X23J
HHdFWFz1cNMbXr6hBw4S6iSgoADrcC76k/poJ5V4WnchJWFmCW9UzAcNBOz9+CDbZw5WhAMLQN/3
LEO9pFMpXQJwm+MbIngBstkbWCjLnzWh8cV8RRDT8EIEKz/Vp5csB+LavlEHmhWjyamYflFZggvX
/Hy2kmHr+GwymFBl4mEwAP/vNQl+Q8ZrmIvXnZXQwI63Xonc6Zqoj61OGXmZMqWTmRR+nyrvCEab
3BbkRGDjeXIx4pO47kalhcCsWlMr6DyQWRpHR97RDXGWlURbHDeBp/mREAlYPzhf7YMoigvZWPUM
WLpIbMoq3o1Ehv0ceMcNSOA1KaL/2bbUy1gH7lifBoK81gEXHRk/nXveRQV+zv81WUEZqrbtvu8E
0hteTt43Obn2MAc7uEH3PJTUKn2XiSO/slh0dT5KKIs2+7xn7YjMtH97oslLGrzdCX/o4r5GJHoj
O5SSDGWvxa94ONiE5KcZevFkFb6P+Rk045nOt0exYkNUARP5jV5uHnv9DpYQy3CousJVqUxcTDVv
ywMu5ZpeSmsv6ljc8bsjbW97u6xVsFy/ewhNGvbgqPH4nJh2pE3Di4BXb20W6XyaYIpR1VYtpdYG
gWLMXvQS2jy2SjdrlUEDmC1CtJaPITJ/Tn/VSQOLgKJaI2qCQTmeKnriPaywnKniSINti1JhjR6d
IE+pg2ny7xmt0IQlTzrGhynR1zjpiIRaAkD0x7ExFW0rh9jr/bY/c89OaXVXonQWzDvT/7roWnyR
rynwn2fz0yW87DMt8RnQ+EfFobyuB5okGRlyFSswQ1GYorhn6wmCHxSAVNVD+CnQVkTowz+HeKX2
vJyISZ0JYhqgTeTN8fjNLGf/x10LXvesg4Vsz2/IkZ0JY3gIH0FOcX+ncpsgkHDABECfAplUtMbg
MM1e8B+7hop8DkvbwsF+LAIBtrEEx/DXOK+TqsqIVR9GqKtbep6TvVPPAUEzyzwQ9/uN2QgvC7EP
u4aXYvhRnPzeRPB9Y77tKRRxnz9pojbPIQjCtH+mXzv10LpWz5YhqVNGInYUkdqxOhNgDjjbMhae
Px8rXBztwtKqbxiqs7Qu0grzgRBG6d66+/Blhoqz7aQi2xVmijdPl9YXRB5g15ooGIGREYLuUWrY
vKtR6HeU3MQtl2iqMeQyhUfwpPr+7IFkgYKGFgRZDOfuxUL+KmDqJh3RZqTpNA9PcE/2IIgi1ItP
TjveogSxHXPP42nbyrS+FA4aeYa0I93rGorBcpCPTsKy0zRQVehC9Qjf8WyLnDTPAqzl5H3mRMFo
kpA1H7i1j1FqoggIfXiH2d5b3FS5bY0UFShzehcKxflLGCkowMj+XNSwHSaZFQ/QYWiG+Vc3wxSM
nPJAqdRt2Bdfxmsuw9zhqcJiSehGuvJogL0CXqMMrHQLOZJKsaGn2VF4xdqZktZOGZ/NVEwVTcYl
/W72p+BR4dU3Y8GEzEUvPRF41gtqH/aFoFAAWqxS7fLzYEPDZRBNfKKzXTteh4v+BNwmdShHGQMA
10oOj0EakQ/sdpDE0X8f8flVPnDwgQnFuvp4qJC+9mdQ361tPdLGGHEpxfJqiamv2u9JlVQs2DsY
dhiMGpOuSVGQvPEuljsT0RhGzRwJ7h0BKj0n0XoqEcAT1+OOrudR6xBdxtYX01YR8NGLM3b9f88l
iidhbU2qWTaYJFkf4bIB4WuxIyp4MJyWSbiLS1ZOunIoSXC8UpsfjAzYFY7DqWRdAjSwJ3b5ZU7p
wnY3TbEzTkNXjeKmtrCoV45OCmNFZIrh4phuI2Xb6a/MIj0UXWhDvJSFthRfQuBphVUyDTUtZtpl
aczWLDeP1bvPZQdgW/THthHTax5OxbiY2CL7o6rEAxiFeNJ9mjpK9DYETp9z6GWOaCV4745Rncfy
yZtgmrfh5O8njWFUY4KQlVZMnsiJ3qoHgPziwfZAYmuVhGsjku0O5LmklKMc/t14qywSkuLc3e7X
RNjNwWcy8Ph+ZGiejemj4DJC5+eVWuE8sR6Uy+WTN00IpW+zg/Pdrc11zI/986ujsk+o/HlMfzR2
IWqy+H3VsE8psOfMmsbmMylaLjaUa3ZuBX9zFxL1G7wnQyiQ3MwCqNkNL613RwU2AZ/iHc1GYT7G
hQa2nIzr2uNHmQxcwsaH/RxLk8qM1r1KkN+E7fbWFnw3mHMrCtF86wlGDVbqwJVWrzPAdOs+B4Bz
ITD5KNWMSjEdL71IEUqdgWOCtEkSw5MGDsBsF9K9xw3YKZy5TT29uNKHZ/x8u/tjPMdCH5dzmwwh
xuN0DtUwAU6wk9p3SrIyULnzzXn6EiqOmeHKbNbOxhXLAh+sIQIpttd+TR16bmuvwjiM6WdTtcit
CiCmOczEMmOEtuYReZEHfT4gX+UVc92Mg92ONy+m6x72ze35NVKd+3mgLiiUDoPjYe5/o/gLOe+j
AQAY9sQMyNsqDESCzzmpU63JKYlzkfDRra3wMYoH+z2GTcOGlXV3PfHU0m0982i4DAdX1q/MbCbW
Q/6gctYVTT/a6LjXVQbTVQxFZDH+mPcWnwbfImF4mlKzXJvlpkjbOwfIcESYZBOg7PWtBqoMgeYX
0YwQ/D/eDm5STqRNHDnATbpSEeqcsrOyh4QA0QCt8Ttd2sCcM38C/dolHVx/jpUNr8x4i8SBUJaE
Y8vj26qu9wLLxQZYZRh1igs9aly6NEoFJxWVZiICALte3G01em6hpOTAHEfaXQ0O44/gS7LKVq43
xALWxbPlQ8wuBGhkvKUcX8JFdizOozhyALpy6DQrShH6wGfo92x1eUit3nsy9glaXMN9/w80RI2Q
QWEYVOTOOPwURlbIVv0Vt/7GNAmWrmKO3t3VjytvMgE22yOOd9h7xjq9RLtPR4XLFKj8E0i47Wg3
oFW2Ud5Jc3Jdu7P9fuj1fkRo1siULq+rvocsflQpUeHrr7u2q7Vl2eQYuO0UiLaR2kcsXsfC0Zc6
VTFIkuLie28XkLXDZLQXVLbRRLa+llb0Bou+mrJkp5P/f6RlsfkGQ6TE5LrCske6YXCgez8nRwo3
AzravPrYuaZE8dfOVHeaAaHVgN1m/VjTA4GLgh4LxvsawuAKgP2l/IYeCQ1aK1U3CCOAgz1vW+mc
jrskCFaE7n9J1GvRjLdAVqSk5QQTl/OBIR6rerrvoDeBSpilVqF8yDMMRNl8iE1jEUHDHG95MqXu
SPrv36Lkiydjri/UOIYCm+SIlQNx7h3ANgdM/NMtB/pnnyIeQiavbEpRE4aI0KLXrFQBiiItUVX+
+kxGtJ27OjKr8DnXWUOLMHWSIgYIqKbIwFQQCgrUADJU6X3tDAxP2AUmSyHPaOekrfSQz+U2psVH
nMhrfpT+OlQmCRRNlFFl/3Ap6ik0tlVhT5ZRwb1NagVb59FYq8Jk6EtpJuFxDM6hKlY3q0QGCCDc
x1HIAykHri5g4HVHKRbk/3zWPnCcFCNoezRjXbjy2krJDXWOi+XXVyHFyNVc4vqebSN96k2eBwYD
++eFp+6sXMPJqHcCQeb8GEkUzPxWUz7vEt4jNyOMiemjFw3CYTczQeO7XOp7V5Qx6T82oZIVojgO
9beLP8bFPaDaJI3G2hzjUy78SFQpS3Y37q/KLauLElSULwAO3Ixn66W9a9GCg2hvjPD/sSVgZFbc
uIOInm1L5E/0SmI2lLFurb1FuQZsnF4I08+jKvutLr2uC254vjqO/lCQqeX2STTwZHmQFBMRbFYR
c0oA2vDI4eKL2ssgLUyguxXOl6BFJI0jorcVye0oRHG6VkvAXanXecyu+CtP/lzTwtQFL81YTIKa
mrfQOBYf9HxEiQSvJGBStMMFJrNdaHqHSMoNYs4nIME2tEGJESECmElSPAVSirODAgBrxsfI5hJ2
LwlzG94jpBflovZmsnCZrILhDhsnOKD3xBhrQZvc7gDCp8zoV8WiRXJxohf7Ca2gpZ3sR2Pansf8
xB1MY38pQGUaeWj8wYyTMa3mmwTnJgTp9BFd5i4t0j/B/tStd0LO6fxzh2XCNfD5hcGXFxOMOUtO
fTxrHeSSS0lb0E7kfNB4N7AzXRgjdaC3zl+B5NA8LIzNcse7CJMYj+mXvP1FCcdbmReAtfI+p5go
Dv6uCcptI+4xkp5vaivRcEytrcR8xTZ8VXLQ+FUuFjfnTMQ92tF2CgKSx2GOuZsM+Bh48/fdNNtC
emgW6mypnWuY8MjogRyY7JD9cMhfvf2VB3GA8UOjzV/s2HiHU2k3OTxY3/daxOM0uWn6ug6xcH0F
6efxgWFl8hpXwUzTTDYif52uaoBcqJih8QZttvq4HPDamKr8knKwkEFQTq/xvjRz+FFw8H0ZXijY
L2Hra0mAq63LvyOtry31P0tOB19nr4AMPo01KyNO8B1xq/T8rRcv2oTFbNzI73nXRmzmQPMsPev0
nX1zreFaodTIq9ahgSEaVZiySbthlm4ySKNLRrkUSnhvB9dweB3PRszOWB/OplSsxyrmbdyub7nc
DIyfADGce4mKnI8F97wRym93H3n/aSyf4G3EsJ66HRFjcTU5yhU+Hu1bloG6S7ZUM45LrdYQ4gV5
ymyfJ0Z1vz+OROnCpZc/65MlCknGZz5KlJuV+abjJnbGTbTV8+0KrRSDn6SKsy4Lhbdpl7cQuuGd
uM+AbRBxZK+ReRstnkZiDSbRHFmeGOG+Dx4o5R9pVZaqafKwo0Gp0uXLX/XOjSTf6sp00helPXVM
8d+5xeCBvgyuaTIKXibiR4O2H052fo3iA1GQwzvHtpbzJkgp00xN6RIuxlzIZCy5Zg+vT2kozIo6
jsGSoNm3FNOtCc2Ns3dEhttAs3glDFqeP/xN+L3DNQqyX0ezq6bEWbz5UAoNnd1Od9UHn1gFmTVV
jnw/hDOdUmWQuy4RyFJkCEDDMqHarZOobZQCLD2UEHcTAUMQ1FUE/wGclAXccvMcsC884rPcikcJ
+LKntXSo6KGmjXWX8PsvO43c3tHPE8TtKCHFYYcVl+X7hwxb3Awde5zSQfwMK8E4fD1u6rKil4FY
Z5On77B1fL/tV23X+vxJXkL8ku7EFkOPpf6bif4N/qLm4YRtsrcKFs9QG/oXzZ/IfOkYfqdxFuGD
Oc0Zp3jdBeHQFqa0NmpSAlUdqi8hoiovNsfoCzCZ2CGnkawIt+6yx9DOHh9sYE1Za0dOCt2getUY
rl+x4gETLSeCIVjetTB2IGVoJ9D6e3HdLQweKFUhbcVFPAGekIyFOHK1Vw4xpErmjSEfdSzbyw1v
dAzEL8JsqQ+1Vs5l6lRwKXTBqgzvPBTKTsVa4rUkxQ3FnXfXROjGwlLt665Yoy190IzRrTt1B488
ZT1378QjxCUSzlvjY8MzAmqMlwT9ibHgkRfDeTbX3DqtyXxKCkCcrtaS/hwzGkbIQJqgzn+ZHR/p
usoyDzh+/c1x7nmKyDxJ7znQLHdcbhRUETsteFqbpLrhZ9hKbe2QKdhP7CpBPoSEG1wLnNGuvZ9I
lEdhnKaaSe7glt52UGsTND5i+UIiK5Wt4V7S26Fyed3vvqeJvsIZ813KZ6Wn7miUc1ywqUdTc3bX
lt4aMuPfR+qkdubt2+9MIc/Lde9z5Xq26l5VFKRlXZr4jVCUxHjt9jXZs3krAd5R3ohU2UrzTmry
XsjPC4t2dA0HRo0I5mn58/Pls/DwlZarUdHX5c/kgkpSLAHiI59RXE+vWhNfXkA9aCiW9pUx0lYa
qY7d7iVGjqWllyBXhtMKk0Mmik/ddNQsCLstwaonMkMRdSfzZj5ychMTwXDi4ANUZsulMGN2pH1R
pSYqsIL7KVExZiHUe3GIjiKH6bEws6xAjZeMqZRWLGay1AYRwCyCDCkI+AnyTG82apYiPnfGU4hE
AcYgrbCRXXMfoPWi6nygM49qAF9pIln2sjPPdScYQ3pY+YghQwep1/ChTi56uZxNpCOMpL7iw14i
y3Eiu7Mk2yJixgEMOjpZ8mkaQP1TRGSAC8YHXMbCV3QlJDySsaYAmdRmAOiqyqTZBVkyNy6ETQQl
MT1eaIVLh7ZYky+P0XLeLpnS7mimMmqOkA141FxULhT4mq8LSXuCF8iG9U+k43HyI/nlA6xz7Nr/
w3ECNBnTG9WB9Yj+D17YRSEnF2u8DIY6vOoVzYlJUMwlwxN2GCISxn76KC3lhgYkD0VTvf/Eq0WB
+/ZwlQFdfDmGMrl98spF09UVWX8Wzl/Tk66Ab0PVhyvI9WW+MSqFbzFZ0LXKnztFNezRRbsnX7hX
Gq0hIlsUOdSsMdovNliSZ1FVo9VgoSOZoKZ/Dtog4KcuhxYpJspPDv7rc/ADbrvYKA6pB/BY1eFL
aqcc4kyBz+d3ZiXkmnMsMbMPU9jCT/0eIMondqZ5c1BOvXnAaQtmdxhkTdL3VGM1rbj5vlBh6GEp
oRk6gLOIXGgenSMhPw5Sbs6xc0SFSnj59b8zUEtJKv1p6QFDRVaGwoMKh9xoVTvOxzXzia+LGxS7
QHDZRFP/7cSkHgf1DrfOqrztItkSBc4HPhvz2UcuZxIcmnjzZa72ZWzUq28bQwNTSBDuNZR+00jJ
rRDsmnA0PIHzwavCds0PJfd5xHoc46F7aYoGBec6JbJUn3D+JqOu2LB5DfqwCVTBpKZY4b36dOi2
BjRkgaNqyPWY+I5uqeQao/mcUl0k4S2aTTz3ykDnAbKBAC+YMGeG5L2ohpEj2HcrNyUVCfCjwgzR
h9sn0eddjxx77lNhtjhNrtbkAVtiyLVrfy6NSDWNucxn3gVeP+JbzMhNLSfVbv5143fJ+d8yNAP3
0TxWarOvzZAr24GKPSva9u8Ljn5xoOM5JzRCbdz1Q9jBD00QP220NCdyJyuuFMkg9oYwwCEumGxm
Jg33vGf6N2Yp/vyOR9w0mLYGrMyo05yWtgy5Zu3hl6QaZdl+NUNemiT179vPN94CYtxidTSajSjS
kfVt+RGxwQpEBfTfZX6LBr55wMHnlUwk91UmAzNJW8L2RYZj0U2vePSgj1egdSpVB65s0qb6EEM3
qiY1nU4tlyvFSPNusG5QNcg+OpvF0E6+IXnoVAgXyiiC9JIJqIrgv5X7xm+7mttnpu4Xz4eQwnZa
tfZg5LD3AuTvFb6cNNRJ1bWHbAfefPtcnfwNI5V2zqvOHRWLjWE5OUDX/GCyk2+61dIipdtmnxnx
mrNUOKgE24HjDjz/Zv8i5bB4oCU+JNMo3fyKxNoPcOeyNr57CtivApnNbEKnCWoLFOBANXNwM/U2
2GD5V277hhGsNNDAM+b2qPih3bgjvfl+xvlGirZegh91UREqu1G6S/de8gbccp9n2n6GV+fl23Yt
/QyHEEieWBo27LpfbXX/6d7meOlFP5yA1WyXtc7DKh2MwiHa/WO+PlMSACqEV8RzwgjZnv2Q2c3z
8xXYz1Hoa+hghZzOGLXpVDuHJH6Xit8Dw2VPMyhUCAvWr5kuJ0AaXnCYIIblW4I3MSp71ZDFoG1o
I8+qmXhtM80i9x2e36STIPEXDLtIGmht/MKc5zurcaIwCUogfBgG7GyzJnBRIIBK2t10n5ENV8XM
J0uPDbGFtZCqEGmMpC4N2NccLiiw2ZE+g0Cn+it3xN2qSqZsmXz7QoCKOtvKebwCPOF5rSotZGQg
2WCci+YIWFEqoKmjHe06Fy8Ygz3NGCE32HGHJkphYHuZgXGqcIR9Ipib4/wAUcds27XHHx0mUaAG
NpAEjgQBAQirbm16fkuoS8YMGLoZM3CycqtNTvR8SWSttu932FBu6OItWazCGDEQKp3tjMVa7MPp
mAzP0KwmqCzvNP6WgLT0DYsvPtEmFHpnydRhwrccTagThA6mGYs2eCAjhpgQvpEdov9Hoi1J9v/b
4VxClKrGoLWbMenDGWHR0LnqtpK9lb50SQVPaADn/EuZELPpKRbqUVD0lI8CddN+mzqBYzk/MEaL
5fEVizKEiS9xsZ3u3XS3Xn6SWBEXKfThuzrW4Rz9pO8v6zIacmk+OhbFo4jLPErApv+4Kz3ohe//
X5VI8jhmwF/ArHaLHTCUPGy3nRnnXGJJvCWa9q6dkJMQbhFRYKXAbNSsmXcfC2AtbRniEnD4gsa8
ZGTSLwGN/xdfmBnUdnKD02aLVKAoXV0jcefOoFUf9dXFz3OhU1QMS+N7qcN5LG79zroGPl7Buz/w
HBHcVBaCqF2dDDJVBY0s8uqnvO4JAMEHuEw3Os++bHLOo+6w+KPRW8iOdl/OQ8PVU7lsIrkv7SwO
U+zg54bevnRPX9FGrgdaE4twYcf12pQK/3RvtZjMVZ1deQEvDz1cwLgH16nHAQC5F8FKfVsaU+fY
b4IePzVfGzevQpIaVgjJl/ag71B4PjBXsb5sj+0ZWjGuEY0nTp5LOvnxMvq469Bm2XFCU4CiMxTJ
zkyqq08qk1i0lqUaDXNcoNyB//AkzRC1gM6AsluGL+Va7STODtYiFebPo44RioRmVtDkGiebmwnv
LyuxYX46nWwTpOq/rBsN0VxUqaaRD6IiiT85dm4E08wskNqdIDuav//uazuVt+vM6mqZJQYoAXED
zrbAqWfKB9GfkN6KPthJMyaZIKxtWHOs7PsbECsLUvB7TmPZjTgoRUa8G5o/WTBxceFNjaa/MdC+
xGhAEUZgMDeFkmRAJFD1wa/zdwi85C6XTODkKo05sw1kWh08Z4T7lD2i5MYzOeZgUnrso/3KsDW/
HmtCJJpqjrd7hRVdvGuk5Ktq7kVQLvVMmJNBcbtrFIEKKgvUP1tJvhwGAE00EFctzU6omCrukwGC
gppctPGW0QdVMKz57hv6xRU1uom8udqRAmqwVIhVHnHbbtN10TFNhx4TF0AiugeXij0O1lZReXuI
UQK3T5SSBeb48e5DBDSH/PA4wnktUZ8/VPf2iJlaS6cC7Hx3Bh7+1zE4dUeU4NAQGap4GPa10TVt
v0vhPCXec+MZbGBOid2hA7as+QYREZQy0X4EYog4og5SVzZKHxG50UAM+G1zGqNTJz6j2iMo+LX6
UQBK+YHzgdbzSN9FNYzrpiWnMb36yKbfK87NMl6WMP0VSS+jAQCpow3ET/pnRyzaLPsuY2dlHurQ
VCpQ7D+gi/Wxxq+gEK7zkBYvYeJ1DSyn7F5NzET5TMSUKVLwZN4lnqbrx1ooFRCM1Dd3BJntJ7u8
Ibzlxg5kKg68F7JIdTw5HbfFsDAP+tQ5Y3wm5Dlj1SrxMW4xNCwso8MhNe9DTmTUFYkJAZFUO/JM
ReXVvwgDKynMXaVREcNscTPldJ+gnGFmpYNDp7zVf5nZen4m7P/K4lzYUOK6Zq+Kx2oJChAaCJQu
LTMoFDH0t789zwctzcQ61GRxOGtVPOTr27iieG6QAdn91wxmsWWE4zWm1XpEwZxVLudZE8uzROgD
1tGuuRSphMDANx+GrxSnkOWsKzl8UYCmoBnfOtCOlkkEThyGTrZenU4WMEFzi2WL2ElHSuqsPUT1
gmG20T+xDQ8vEOam9Pkr/pMSMuSI7BxfnLyoZ+inrMDEPG7E0ZY78DvCuYeHelWnDT2F1YK+SL5C
nuikBR+TB/gYpk0Nh0JsJu1aOpjbfd6gwCwkaX9kYfDCzxhmo9TXsHZhTkf7keiRkCqoWJkUzCg1
9JtbTNbPvFmdtPs3NpSqAsxqew1bfOQry8zHC3lSLzeqpJvkFD+BJpl4JPqaSk/irZpRmzLZzGTV
q0kJA4cln//NbqX3Jm577s6wcKEe2jL+BORsIqqq1+wPQsYz2eYqPH0YII9sucoK3jx/54pfYzPf
yjbbX9vJ9NfTb5FjTH9F7drbOCfEfn0SSfI2Oc4gIJcG0u/wjTkEo8dLPBJ1M3Ejx7cU7VrSYisi
aIvax6d37cP0HHVetqDXOJMTx4+XhZSncarrbWGLCJolm64ww4bzhCbSUTq6RJf4qE1IhHhXMHVr
OcEB1g7CsKRa0i19EF1RdUty09Zmr+Fs1+zXbJyWlO00AaCsE2wGSDSDb9Y+/HXBnBer+FCq5wCG
DYcfDLy03TC0cmKrY0kR+RQ8cfV69Pe4k+/4vMwvhNj5xzc95ukQS93PVL2cbi5Lx175ubJuo2yF
oShaH2Q6V4IpwnCstvOXy+C3zATEysYHupTmlsNBSE7H01bCHi9EvDXHIzK8YWH/VOlWVmpy73R/
5NaRo1vAMVZzUP50qn83cdXiiuYx9HeKGgBrfUiaPn43o34mjPPGH9uIWlzfoFfgdVLM1tg5bWbF
aoKWgwXjIf/Ple/ADRxkpjSR6TyQITQYXPRIw/Zju7x7UX1cXaXcfaOBfxuqqt6b+XBLk0vNCEkh
JDQ8vb21ZuEcPH6pFSgzNs1fXtj4VmWTSwhimBcPKBjMdTpjW4CgcCQrJMYHSnkM2anjkf4lDBnw
7Xp9YTFTM4Afen6tUzfLBb/UoabnWlQcGU8PnKkPqDrDc/FyGiiPKmI04ROM+hBqWpQ8fYxmdLlb
BLFPjt//SoZxlzygLshrEfgRVMM6M81ZXr4XZ6c+5WWgdqrqDsiRiYorFCeBxsSL10f+yfjUFqRU
/RBbCqQNHCoWmvaNriC5OVJoZkWsPRPckEZWCavholFx2FQMITPUeYJunqUujl2Q9S5/Ilht1Tro
rYvgGR6G+6dVP2U+KApOb8MPKrgfIDAYWCTbIN9MOVJcmIEYrWmn5FEABhC/9LIO/K5+F6ITAW4H
ugCV/F6NeZvHfyh4aBnNiHqrDtDBZYFUdJSOvC7TqlUvRq9J2VkyR42+G/9wJXlQK6f5H8uP2vuC
yELLztYOIkRase47vqlA3LdR/A3rG0/8hep9n0pczPg3+ifgTbET4r/pi0muMuRiD53xa8HnaR4D
JnUkb8OavW7JSTsQoLG52/CrsylgblNdbK5dwUjGaiwQxOu1NesVkiakjjgEp0t4xk+3WJtBzoDO
acWWY4DQtcYsOCvvBzs/lXc9aYQ8fp6SBlRTuOuwjopls/mRWxKKWfrSLePlaj7htCUa/QIl4qN1
Nsmt/pFY4XBMg0s7jSwPl3Jj9X+GUzbaWdQNHItPDdgkp3j8feYF4OnWqOyblchP5yBULe8oJSj3
qgMLxkbUfMCu6k8ZRo6XYhAyLDbRS4RJLggSo2zIlJQ8m9Mc9KKcIuESkqacEyr2xBybu9wr3ZiG
ZESBgyvaEW2Jeg5bjrOUWGOu2NWpz1sovBAF+1qJqjdywGIJs6N54Xte4ReKZ2XISDcHKzkN3nM8
+JLOJfwAqO7HO1FDEnhh0/bArFLrnboHaGVn9jo856okymBIl+5Y9RNMCV/zZWrqH0gUiv1akT0e
uwNoglhvtGAo+BDVDq9lxSoR3XYzCOlSDxlJrdR6DV1BrArABrR4wCeyMl6HefwStbRlZoVvYLwl
yFhJeD0kr44JoGnLnrfuQiy/bL6eBa5aq+lVA26R8gGzIbEZsL/9QtUAuOxpX/CILsTmDmVZUxuE
MuN6FUzZEFcZcc7NGGolYIdOjXODDLdKgbLlT1q2r0qG5TjH0O/zeN/WQCyopeYpmoA+BQtmoraD
wmsMv4QD2FU5LcN5S9TqAuxoG1xxdNHlERyCDzEV+Qd1ItrnoFYVQAyCKLKtYICqrBOO3tvm4gTB
lUIxfyzxfYCgR11AcVRkqFQI+mslNzskFYQA0EbhPrALFj4FjHNNdCZTkqFCe9l4TP7adSlKe6ks
R2PF3PWlotiPwEfYDrrFDs5N0hLUKzyVFkSh7108N4ZgwXyvig4BCyLlTuQCxIWvauVmPb8FCv3P
nWF4Z6XulPAr/hHmJrFHkyYWOxNoSSi1egC5ZZLGpTI6Lxjl4HRGJjNwy7fqspOrZvNrYQSK5n0J
aG+jPULU7qXPb8ZlkDi/2ptJjTJBG2p98hcI0CnpNT02Bl0zU1miKPZIzmoUm2ic01PSB2vGsecE
m6cHmG16kaSJfahtRhY37rQVclwWZslTQC/RwLF4+5kopvciTFiO9tiQSaENw+PCXxj0mJquJUw+
JNP+DErRGznnEg0qyLWureN0eAy3eUsmW5r0ScpxDh8LUHuCzjU9QVgu1nomqv7C4vqejmMnyzyT
B0Y15FI+MqrMkspkCFIiHX/8pAx0ek4OMepzANUXgeKH/nMN6hsI8pMyvDMg5yTert3eqEDr/sGx
BWlwZAjgPb9FiWU8p0jAF/wCkrUwdxOkXMQc/A76YQG505ta+DLxvw8ZnZKO5g1OZCVEn1rDegZF
AueGzP71+SFtkd51MRLWQcBpY1xTlKTm8epI5vWe/C2+sPYcjeUsA4DWwFW1V4XMMN7uVeyZ8U4Y
lU/Mqvh3FueUhkTvooiwUorr3k4oIgCU8cZVh2cVgOoji/qT0qTMh9QkEbxeD0Y3NlQA3Ij2nkUZ
pTywmliGjrihW0tadz9taOgtpJ2WuxCQMcsih+BHbj481XPGRsEv12mdSyKKgR4zXcraZtFayn1Q
KyNJvJTC3RfOKUOE36xtqN+2klBPooZwUlmMLlzdb07E3qCHIjC13fG8EEXF5YMmHabkVpRfsmlR
1bpzYQmdY4+6alJZjHKRwRrE8fbfn68Mhr4GR+3ySbMvQuxbM7p051eP2eHhJ+G/wvcklEB+Qgg4
5jD/JIlhyV8acGpiftlyqc2yj9Cbrvg605Wkl1bbp7IiVDpdJhlwsRAQpXbPjgdAWihCmOzgoNIo
qi2EyfPtzdIclsJzsyJFLJpGwFjMJ+vCiWBzL5y4CPlawEX47aJJNDafqR/+ya7iJboBNjKvj0JI
IAc1cx9atj5lRxLmTP4WWx8Et8rWk49oUU0iYAfngBjXZMj8dTtertQIlOvhbk0ijnXmtmal71B9
KYxvgpnHNkOio6ra2wmFnoqh4CJRF2gcEbupOr5XpBpQh+qcFVlzKJsByEqrYWauyezmFNHE6s7p
hSxvygQyLcD3bJo8VmH3zS01BNAeRXeXg9Fy9G9ZCOSr06en8N/BJtCUXHRCrr+7bSR4mY2q6CVu
RGKHOkwgblRa0gSBCAsv76VRWH8iWZ5OTou4SqcOK+oudz5BxfTs0p4iNEEMB8VPsRPErzQFjeRS
yDODdHl3jAWENbkkDZAW65LBN4unSJOBV3WEC2CyJYrVXlC3EQvpYDGrj7FR1Jog+b7GLCw1vZU2
e2wo5ZiHFk1A5RRO5/aUQf0778y4I9FYMPg6FQrhq0SERVtpqhRclzeIJBhHtDSVjLE/g65DEKRj
YQUixwMFPbX3vbmSue2khUObmSV4mL80ZpugUbDSdtrGlJhM1JE8dKKMepMlqQnW7xtffe9Of8KE
bQCdPJVQ4tb6nYV8QcFhJAHtxp7ekbA7sE2LorFZy3FIquM3s2vGDE+hK0e2rKejFs2oFh27ugtr
4oeNEHiZlu2xzdun7lXgtkmwFX9wr67J3/DutsHBPU/CGdffvshfG7snULiJGmjkHVQeFlk4DDlX
Lah788V2/UYUsz6DKJewQbjaw3UkQEag09KKUpbZQdrclcnayg0Os73WeUzEv3qxKPpKPDIe0vr7
bsv9DWaC66VO6j7+NHx9daFuf3xMTe/hWSJYD0UxvuimnXcgUVUhdtc06m1SUPveDIFw7bLBwsS8
NG9WfX/8BU9wlGG57Aaj5OFr7n6AjWGfgWQs2QyzpNOsbuptcjSjHqiR6JOnx7v9k2DvYrBkWAPd
VUtWczAO635KixmwKcg5/17cXyGorvlh2hCxZtzhBNsOFy9O9FQ0CUwdlhcFlFhLkWadUlTiy4jl
A/PdZaakYWlFz5/+hAYNPezAV3bfFXtTcAi2YQ1+8pk8/piOyiWea7ahGFrBgpzFqrsuR+vECOfY
j/7g5Qk0OFoBXF8mjbIs8vHdaxmI4m4sdjJa+mEKx+ElY1rzvUOZIBySmqONhPtxxd65tuDrGkt5
jn2Xd7jABQ/M9tXxj27eL4xQ8f9R33zPm9SebWgeoEfDECCCZGuXZIulEkvF8F2PGQcWUinPECq5
UpVH8Y+9A0RZUDuVXHdI9WT/APa40hLtWgYtaz1i+Qc1nt+QGieJ0aM0XyTmw2YSZjQYytARSrbp
mG6mG/a+gLCtUVh3iPmuXL9JrM/PqA38e6oOWLUrT7f3AVBE6MOebyd0qBYGstgiMSKXGZIQPgB0
X49C8L0fIcQYVNifN5bmXWNndd4nx2qsM6bY6jXFfHbh5rR5Fb17oCfXbFUIB+cTMG+aJSmgRaNO
AR9IwUpboomGRKsdfg8Nio4MzWBGvqaybwZXxndA/bDYGtx8Al0+VMgIPlIlyWUuDDyWHSCzKg9F
5UJpHMrJ+jF/qxF3nQxGofUsZpgSDUHmCDKd7kUs22e1LW+Rrg7WAEMPos8UgOduQW/fJKRymMHN
P+xfHa9XCDIMjiZn6FXvl7y2tc3EQ4DXQBJx0YgJ/rXhfwAU/xV3KONLQzlb/gO4eE+FMu6XWQwa
a3/fWmmCz4oZSJPcXqduDzLyQF63oLyuOT2e9VQ16Dd20s8xOKw6v68Q+mm4ZfIUFv7XlJ8jHu6L
X9AEOxRqtkYYiZBKX3JzYRO1U9O+hkWGm80Troqvd8WDaLEw3A0vw99skbwp7VrIKS59D4eoqGeb
x1BxfnLR86PuSPXigo1fKTcqNTX6ecsPTgBh3bDtKakyzC2gm3P4dAX/y8WORJ/5/tRU5KxEuG33
y2Yi7VvGD7XJzvHoCrSvxkqS4y0HpxaSFVdsFehxFs6qXtSPM7qcLWHh7VhzxDwxr9TPh+tWM4Ha
PrKBQG8vDRe5RkU3UmpsvvB0E2M5XLTtcrNJ+o1p8RHqqzMXL/8EuQr0OHre0du8T3/VGfEQvSXo
k5yTXx/t0qtCxumiNeeVfYJZ21tWb5EgKQ0FXoGknYaiXmonA01SS85gJjeky9tujVr56pPGy1QG
wMNhywCmKSjpu8AhR8NEQtDJqfmDgkYyW6YJNGKoMVeTOXAOICK6dgrs2Ky6E0cx7SWgTBmdaJ19
TEg06uDLYRyoCOxZR3HuukkYh9+67gGHeum3L7yjqYmxZWgqGvkrgFqdfl7Ud9aylDUSX2HVXZZU
JXTgyfIzpmOGO8BjYYgB2Er/6QPTrSAOqEJjA64KlT6N1tMuh8d9zk6kxN7fVBsKmRlVHkN0yE2t
qKgcuuPnU7kUZ8QTJCUPEL9BDK6m5ZBe+cm5HuDjH/D//Ag80ISyLXKYGgdthuzm3E7e5adXNE6y
CMvjdJ9ce+1NndK3MOAcLe1D5w/8Mg2S9UTpqd9ZGhbeKawBcZL5RsQaCswyeZSuX8w6tJnhxD1d
cqGei4Hd8elCOtxVz7YZUvReP4SBxdVDO2H7BdEdM3UIpnAxLEqoBtqSmozDcr5Uz4Y34BCrgKn/
7olljtLGuJ59ZRDBU8+GxCPHTgwHiN+/nmV/iVc0YtxZikz0avSjpJK+K7k+93984FCLcvmAT7+Z
3LRQW7acfHnfl3gQVr/m3C2tXdsGl1NiEl8vJ36E8DcD41znyMliEla5YddkYLvV2UaL0VPtR5Py
8yDapuzyw4swYXAwem5BDol6DkEQ1MveZBYMcnMkCXfUj6coJFuPoUVtkV1HPUb8zrLqw3/qMfsk
FNDBSea/WuZ/c2AJf/NPelpHGoHx1jKMv5G7D87RtckCA612VcyqOBGpntx0eXL7kQPRMMfP3/44
M2Z/qwQ1QwImcuff65927QKiwv/0g2URfKyx7N4LI5J+PPmb3gsOQZR24CR7NK/rNcHiYDK8FqCQ
Z055YSkLmg+iPyxAxMgR7KfefKo7f7zKHBApg0iuHk9rgrZKDCXVTDZCvtdqQoXN8+s8Uesjp8fF
THjOcfdTa8tmzahLYART/8N3BSANLq/RetJbdBbYb4c980kjV9v+gUBiOxFd1A7GCb2uo+rC1Ql0
krAgB1XeMmXgdMuLCdHucawU/f5HtAqz+YsVnHsmuwgP9OcqQnRva7huBdRzqiOP1oLOvVgbRASg
oRC4qtAKAijwdKneerGrnxjcsLO26kH8scOyMV4L5cREa1EgSx+6PSlVElzFAmHY8WF/CfLkTQuC
Wpb7Gf8C3tV79Bq/mYOmUmow8IU9GkUFdFmVx5RArL7CAyNUpQkEWz5wzfAPCSL7ocPLLwAm4idx
X9TOpjlAXNvx3WLydxWqtaZhU05OFj7UBiVbBYAGUTkd9RQnxrOQpQoG7DWqWBelh4bb2q7MAu2r
2KgN002yT6NzHsr4c0rby9AzHJxmUaZMspIU73JURVZNbfKdhMYP2//sncP5jtgtUDDwqU2Z9hYC
dkgPskJze6Drwnn4yj+IQoE5ST/mEPFcIXQYvw0D+pDLN++4nWlfXQvO4SWzc8Rm0KNftPC6M8YI
0R6+h5ntADIxKCvAUAWafqt8HD+/m3XcMesqgTw9wpupcTcDHOyG1eFcKNOHYzN/HFGIcF0UgfiQ
ysSy/kN/W68VllYsr29j+Q5OBo/sFcNMsi/g+YeAEIxZy9p7PG8l8qJPVUjpFDQv4zZUy+4wo2Vz
vfApHKshWZoqpu8JpKonLSVXcGVwTRUzf8nMJG+kRGjc3Ew/SvVFp7Zi/JN2Q99yLqdCZezfOIzW
85JS2pEOs1K4fvL9G/ie6rAvEJ8Kx7m7cQcvdyBsfBwN2YFELfw1F9p0Oj2HnlKq3HzbeM9Jm7ZN
uQDIYkysXIgVkLoe9mwohJ1sUoU9D7BouSInR0SfG4u2m/NgJeKDfsAzlrON8FU64CcyGtJqPNO3
kXeEBSh4RiVBgLlbAPGJcQx8SxdwWtXuiR0wvfqvAQ9Z5lpmgRyLxr/H9gYtygLVioK3BIV4CqHb
7Bbe7sGnwZOKmCja1QxV2RGkjG3GyGsrSl6H2GVWB9kQHQa4tPOqfEJKQdx+OTu2JrHQcUcgfOfE
8kQ27V04bWxG1BViQEXdRxM2lAPUCU5vWtSvJ21wCq+jIooALcl8SLQGxBtHOIEpJSpEzgJjSU+8
EYG2ImycPmWKIZNGx2xDo66Z2ZGVDI4umc05e4nbuzhzur0bDgv/2CwvepYl6Qr0sFSReHLOlsxu
C+yrv/Wlx7sxxJse1ek+zHdWMib+6QX0pnIJ43DoZCmMS0dFukc66JHSAaVYSz5sf1A1l7Lo7hca
jIAjH9YJGRaQnjM3oEvTp9kjHQEmPvyTbQWPhW8YQJAx1/0GPUw0AMDK+jYanNXMsPRkJAYkTmuY
DSbgLxjpzTH6Lx68qkYBOG39doWkLWZ1cv2xp86BJjMOixqhqhpBJPYWPAQBiMU6u8d4+os/zCN0
vdQLJEHFifIPugBzDB+/fM8mr9fjSG0rErJfMx4gqHM4BRevq+nyy9Nf8lc8UEupn+bQZ7oT6TXp
6mKSETt3vcNEUp9vjFwk/Qg+TGZRBnLw6F7KJQoTp0Yf5kHKEAoardLWxNtq/PW71RqpU/mZEa39
zaHa5wF45SWnXBqXf0OELK4nDNMUpLRsl+PtUZUpKeaPZgZ/866gssydw++zyGVYy4ey2hZn2TL6
2twRmJSNLd1nKWY9p8xjT9e488WNZBxcC18vxLF58nMbgpU9mY1C2xQVqyO5q18W5cnCm+zVc7zP
7DljBPmy/uVgojQ7Ty5hdg9ueG6J5AGiTiIJlhAhjtHwue+AmstJcmXgg2TRcgzUEw80yH0uCw+i
jVPGtKaN8KImhqP+FCXKiDomNaqwXqTPnTBqH3+EOoHMWO7GkaeU8IjXY+lhIjMNmShsI25CA1bv
xz3upNMv3MdLcrFGxvcoLIzVNkkoFTKVGy2qv7D7En9h5PcATTmJ6FOnOBF4m2rahG7oV5sya+2B
JByc3e+au+s5DvS6w6IDtGlFg/UuwvZaxdBjOoJvEP8mEp/Z3k6PUx/HC9/e84MKwCuYjK2tjZHY
qFzB7qlRGtSJJ5Vf/R6BqZJXpMVytLin3B2S06chaDUSSSpdEV4ak/hf50MGsIM63WTskfUG3OXG
OxhQZfq+Oz6JpZy1ddrfS86+XBhcoZ9PvSUAobR7TgFhM3LveQa3Lgq6T+NFU49PoSr92J+4hJnV
BCxDtm4CMzz6j2Ud4eeT30/dcSCfFNvob+kl0rcdIGMMXwnX8SktlywUKQeD4P68D9Yvt1k475Wt
ycnr2yiHXBG2JRDlXgAvMa00Zv9MjZ5Kf53jLPMumfSI9Z+Er/AUmFr/XqUDlAZv0kCHW4S6vsIs
IaWbwfK2c3rbZTPjjqn4BcpY+LCQRAE2GbQRqVMzbLP9s5zHwFV50VoWiWcN8jEquajVTt5ReRI1
eIfTp7hgk3aOxc8xVSM4Nh4st5B66mk58JvFjmC6awXkeDEOcGheZ4novVFRchMV2QhhuPJNndoL
xctNWZGvN+LAmr7qd2FGGyhMsMWDRoYoyLY/ORx7NB/zlzmoA+8MgjfKbqEETFe89PqCyG4SGUBJ
/yfx//+So66Mp8KRYb99FeQh+QUTjqiRpH+rY/FcbQuuKcTTL6SJdlIrZMAN67LCj1bdB+pkKeoB
h/cuT2FPi7Y8P9avMJhJjY2DjNmaSoDQpwXd8Px+17V32MUWHjvluiRVbTRQmifAUcLFnN36xawG
lpQ++XHYsHTSCXw+0FHKi9SQjXF1v2um5XnlThOlpH7BvIkpiS9oVIcsKDYaqpF5h7MJXPjEzeIR
exIoN78OUXhvkNKWrbtf+QoKiqsPpHMxUG3meH+1q/OT1vjIzFIwQVn978yyZlJqCz0wFyBdQxRi
EQBxO0+wU7Tq08gCoaDKxciK25x1ID4y2tufZFXyUi+QipBnfQHKaXK+LtBb3jXspHTWMldlfbeR
Zi1VzMJjopGqdGiBuuZeK8WTn2UzrxvhF6ZzT8EL+EMNB7C5lpqs7NWA9YcLXpW75rD034SKYvXS
AgkoNMPoYLqHNi7MyKEbC9S+DX7lL3qaVzjjXJTug8v9J1SvFqEMD2BiUnGU0BxxoDQ4fCpL63nR
5yqNNKOYXTPp3BeuT+vdAXGib8JcZcSS3RCXJMnEG1dvsIt61DRHXU1rREnq/KdL/e7Z8zD9NYmh
D02baWTg5vXLrzrxf2b43uNaqVoOS8rlby692ga5rtQMJpTAB1VTXMp5NToMbaqyGmq+JfpXmOlh
KdCWcjvzUDTMZCJrO37GIpYXaqO5OmCx+NqbT5qq5xv7lS3KOytgJ6wJ8TfCijWqa5CCS/U7FZGn
ZprImYBcTiu62fT7/5UJx3kpRyS59XkCmjA/G3dRnPaBnXTndO6/izwCPGFXCUIHCfurhxDadbxf
CPAZNdLGSuyoybLbuw+0muDUbjLMV3SaaiT2dI8ocmGE9bhRwxdXNHO/9U9Yj7irllizvCkPAflj
oCX/lU04+n1NpLYykCOfRsd1oBfmxCNBsRydTpNb978p48X41jCRFLB7wrgz35DVZaXDtwAeG6lu
rns36c4lkJcNl7AFz29SG0Iyv+zlJlZ0zBGFWnx8exElqtF2u5zSpD00SzN8/R+SdrvoL54q56P+
JYYIWn2OQNjqqIAKy34PHDj3zomZL6t4x1c9TrJp4IVyEvV65RwJtvj59VC6jBXqGm59ssQFyosD
vF0WYk3tlJTqn6MuK5IUOXibEekShnyLYfyYpnhdDyuKxHH15OZRMUklQy36nUfYHrlk7LbJ+fA3
LVKyhpwSNwTaXLyShuHFLYeE/TC2qopFuFXfeXs6K5hgSyLoOkdA6L5FGQ400W8SbTxSlz+m1taX
CRMgcrVUIib1t5zg7/cQ2FHxai7CAvn6jC5ijs9wGIxfCVidfVh1pOaQiXkKUEu4ZkN92OWrQq/O
JLskqmSetwXYqXklbEzuLkdNYKXwi4Ruc3OEnnhMxHIwY0XIiaRb0sniIpwUs8ZVw2xH0ZJSbBSh
J8oDr/5joyymIyaTF4kvzvZ7mGs6eS1dsxmobF9clIE6xXwJsVV/LSoLrOAMXz8cADjd8tEQ8qET
b41NIt0b1DFgfz/U3rHLmMCUUGrNb7z02srV7nfEVu6As85txDDLrfzy0cwZAQeHIMQHc6vv9Xt/
Z/hNdF0dBe250YFpi/MK1dO7lkTCalZfQ/gF/18n6FXMP1ClN5hU8ibk/EB5LbWcYsOp1TOFULG3
6gAgb8EOhZBbWSYbeFrlKo6huip/OWYLj+BcKdlUE0zhANoiZxNP3O5m04CSxEXGxrFkWYBv2Uf5
B1nzGeEJNmWC5lM0BQUxuJivUisHDa5Ph8YxIknh3KNj+BBszlAV5reUIm0MYPF7+CnV316VFL+N
hno3SeMicCfV+PhA1mAF/oP7vclJdyKdQ8i0qFgaa+csAAfIyOIqJldK/63gewS24qYQjo9M+UMU
EEKWn4sV9aLmyAXv5H4ao/1jBNCAoqB7qYqkOzyb7GO4Tf14YIbn4HoA1gxTqYeb/ZIrdZmKDA59
Q9lbWi73QP6P2zs4BzSCpnF5WuidoiIujwl+r72N3g/pLbhQKd0ghQtWbXhD8fZjJ6tWyL8XAX69
h4tfIaaazy/fA7NL8Lwb2vFUDA3Yzv9emqsH6rrc3Gum6hKHP4MORgj9qS1zhaZX4QQ4fTajPo+Y
V95U3Ly+MaVpNejglKnsVINB43/exrWhfnBJX5jghMRp4YlJpSSNoxwLj8Eokze5plQhZ9WBWsk6
aFBIGm0Ru+uq9jhMrpUsIAKTcnuHmK9EdGos5ZBHoir+MC6keAulh5bJF/IYsXE3+BTrzaxddi1E
iCc3+EmLh57W1ug1qKZDnzlW3f/zM+W0t7Un2f95u3GiheAjyMwR85TmTtVaIyn/7ETkczbTcFIi
wXBYEMqMSIiAHMCO3GIB/0iqmcWdY0x/MaNBMMZuoBx0v87oN6646Zddx6Cp1jNBQG/yfM5Ba+le
d3Nc/0BXXS2+/l9TrLtRGCWmFKuQZ+lCrpFM3HtHsngk2JVaXYBqdhC9uAnqgw054v1iX3u4CJ26
VdLYHZmlZAgYFiNQrzUolob/B4mh6xTL1Qr8h7onXRhdfE7acoXtIQHjMTmyPCxosUCwZihtSvWd
KGmiKnrpGyVzvvdGccANqFEKvJTa1VnIXG3aqzU/wxjyov69LfShhgJraZSHPKg0eykK3+toIsC3
DQEmUvYrJt/puSSzxG0JJoE/sb5gnwcGmWZUYjudJkj8VS0HQnaWc3B+a2LO/xMTEpM+opG/i+uJ
VT0X1zAd7YHNKVTnG76I5NJjneXnf15ciMr1SYkftXa6Rpc25XCNXcNvU1om4iSN5WRroYCNC0Ky
Mty1ef5phC5pS4IiTR709FAwKA03km8SM4nuRd+Ma/srKISNdX/5cUKultyzwCwcFQu2bbsg/gjt
TjusmdQagfccdf4WO6ehR1Z1skOGGD7u51cNDSBlfCU2JdtwywJ8FI2ADQ0KOQKAaaS+tTUTCkYv
DChhxEr3ZClchAhL2kd4hhzepvGMEohaA9tr96U2IreNKmZnmz4R4MzCl6/0NXg7nf6OxqX9p5vv
+EcLIR64ss/yNQHoeZSGxl8fdVmNNyjbOrIJp6V5EDGO2pLc9sP++5EGkunN9mSWOl8EZtnEVf4h
jJTzga3RtPLjqfkHhmzk5r6ieKRqt+0+alEvfxbTSQEKq9Cn9aj0K1T9kdtrQNXMBr+JC6YZ4vSc
3d6vvjGEEOIWZvS3dAGWT2SKj8zGggL6YchyYSWXFpMbxFMHqSKWGhX7f7VqEOvLOs7n5KF6fmOX
G4Q20+4LTbeW5MeEpZ+tAasxIAyCR62f3WM93fi00OefsjcuR0eN5KNPKPwZQdfwI5DP+d5hDtjT
cFSegP1k9fZxexBt5cPrF/O7GVtww1SojWH4ADl2YeYeBUt7f34Tn1AhM42+Fa19wVzK0sO3X923
nfU8c4vqzk937elW4A7/B6O0uAO5MKiW8vek9ZY2wiqFqv89w2W7zE7cosKrtkO4UrJ1ZBtTiVr6
7uKE0FJqzkIJsJl7OeNEXdEBeF/Hu2kPNjPNlyqSeh7raym/izK4bX5WY0HIB44lt/kCDAZ3r1QC
wUMeB5lGmh09HTPGWvh5ncB8/xDYAOyU35/POy6umKKShDiiP4GnIaspoXNwFt1ciJEUUMXZJr6G
gOJQ4uokxY8Y0BspLiDOucfqoHVlRrv1qo35LVNwUgR5To8KlFcUKVBLkCTxl7Nc4/uJwU1rqqQ3
5fO6j8n++yCWPkDk3VJlxcvxqsWvQp53gUG5A1tTHbVB8EhCO7bE5mTUR4C2oEugTCnIam0jyOeH
HTUFVdIzD3JhiYeRB+M5qztkZbF66nx4MzCejF5UsCLtnGorrfwUBw5EZ7/l1Iy3tizhkX0KaeNH
f/qweL0yq1gbfnVdxPjeS9vbTeLmPEo7g2fhQavOAWioAPCFlzdmoTV/GldCDiLV3skNJIriw6oD
W7Bn6SJwqgVzUtCOqA9wSgF0V5q0/r05i1xO4R3BlF26bQOr/DYeFU2aVcIl9lm8MQ3QaUk1RVXS
/HD5pbzQgxLKIczqIsPT4crFlQXjcr+hJ6sG+vAvl3mtbht2PFPiINP/rtdUznuN3abuc1hixV3g
8SNhLL75MHoeDvQnh9DGI5T7Lo7zFr97TRJ7JndZPe4CVFDUsZ0VYg/VSO6MazaG7nNIfD+So5er
n9gb/xQpi38obwY7+VPjBAOx+r/nPIRzpU1AwXa16SyL8tmQR4jNMRGnxZzXsIqF447RNN4oCYX6
+Bs8mVoOj1u1cqcwgVLDKGXbY3uDXcDE2oZIN4aW5MXoMtJocpESCzfMMNt2gkzDKhAnlVa/Xraw
jO4pBaf38sr3iio2UJwlpV47En/SnKKX4b0ABRffit36f4tteOHFyQaHFl2hhrtbP8vvJNpNLnXO
/R3uK7i7iqV55T2mckpa2gD46J5YFHyKn/V8qQkwDH2la4LQsBx+I8HJPcolo0+aQzDmB6j2R9C8
yD3a/cXCaMoZLe/9MucKw87wJKuYL2qHD6eyQ4BtCJ0AQHdqkLD8bL86fhGKIgMsbJA/vz1GKr36
7ksGF0LpCS6qg9ZIqRSitWTJcryZZq1GUuFZuOjSrRAqFlYXbK/tPAY8MqLQSLkWq6THOoyq+HaX
Ns2xIthiPhOadJNUElOdAhzwLTWun5bn5BrgmeOmPeXLooCtoqF0uGybzyPacUpU0BeBiEQ+mN/l
NqCoIxx2Q20wKeaHYolp/UuKgRAosdpuYNAHqyJknSmTlycrEhkuNl4CvMeWTM5humZqTl/1ZvTv
RU4zPBt1Hljm3MjkmHsrV+Jd85WNGl87AKUg0ORMab63yOrxZT7SKeNJ0jAvWA5a5emcKQkO7QF8
3HX+LBEjqKbAzDcT4dixp46HsmxYLDTk8e5LY9X1CPdrMdVZ9RqY0rlIiZLN4u+d9bafc15l/6f4
kxKtGOjm7lyxu6B7lQUT3GmoNgG9ZUDbvyffP7us2HvSQp1aYfETKZbDhmUWuC2wayn416HYCkaz
ElHy3UTHe/nfgFAfDfHjY/Ja/f64FhjLaN2Lh9sthJ0JwQElZW1Yl4HT1YN+xEzAdxfP+B/mzZLo
R9nBKL1fKgax54SPB86o+akSqLGO/YxejLecTn1bDghEwTmT6l4Qk4OcldFMrlS6rInaAXDCm7NJ
34gQIzUTpE/IvkTEDjUyolsR4r+CKkJwE8Tkcdvjqgch6mdL+MoxNBKYeQCygLiubLfVsgXL3jhI
czv1LfQ5b/BtOFJP5eADb3ry6AWjGk7AcPQgf20rQpigtP+h+jd/xrLXuayUAbht5h7W9dnSfV9C
uBasIL5ZYjtQru6rUsmzaJ1a+U0iUsHF8MENH31oP0MY5fWl61l2vDWeorbeBA8E1dmjczyjM2Uh
xRpy8mIv0oroxJxLJP7FcQZUE15pUdieK1sn+kxnVOOAJGQs/KpVDI794edlMYT5Jz14k1ei0Kbs
tC0/IXc0PisV+lkPJpL4GIkKUSWFnDtSL2H+9wSOmekYqzjqbpIKuszcDS+bY54H0Y8FE7Z9RxK9
Oy+0/Buuwq9tRCdi6gugDSuOGk0dSoplsXwcFQxV3GdXREygcCQykCbYLJliIUn8tBDmD9uIba1G
GRfL81taYZPxRvxsJfJ0rddl62sEOKFIZOZkYOCx2C1EICwmaeRnQsQ0gbl0DfPjwpQQ8NKqqY//
LGIGjg1ZIoIM7tOUN5cwihY/o+zDZuHX1gua9dbRuv5j7KSfYzktqFTwotd7uq8imZqdK8/VNLiZ
6Kg9Laa3YwVOlZ2oRE/zzG9+lKuEMTCtiO6zt7qo+DapUdBZpHEk7HevFmM4sYbNbb1Q924yLxRk
p+vBcUahdhbRkSCOhlCMDUZrZnCbPsh376kDtGZDBHfbrppQfQ+xjxDtzBgyVHdlm6DP9AEDxy11
lSCUhvs1LO7KyHmUxlGuVxjFPlX2hvA7YBMB6fgtWLJchD/88yU8bLEjCjtHVYV1RkWo7+FFxz7d
bHSLginyFuVPYQ84tzOn/kSsgylMTpvOYCUDFV+Iaj96uiz4IxaCeKbOjRH4Muerf0T7b8uk1Q7P
viaqVsSGscrqFUNLfGL2i2IJCFHc1vdvM7G9EgVLN3r+LF7SJovzTw7L1jrAUEI3LVhA2alppcwn
LnzCvuvAeHobeeB+wdsDUDjEzPkG8PYtMeZlZZHqKT4K3LcaVFGW3SPhLaeXZ9wP5jFJzsKaLBND
0JzRo8hW5JEC+O0SgFA8Nq0H+jeB06S3GX9QDTXF3jZqbxXvcPVeucpcd8BHSZEvXU3EcLJzgDjr
GynuMLAvx+IoTAaQo66NKglhqCBmxSzx/rVv6Xs84l2MvLxTfY9tLrXfayhd5KRBILyfP/uYona8
utyfEzEP6myZRTrl8Z6tlW/pOUNieRhK9byEZf0aw39kZ+vTdtlP3F1d7scegvvGNAJwGKXj04SW
eZUGr9ieB9yrSRpooLt4Wxj0CDLgh8888lAd2Ffq740zpapDwlngZ8LxSUnbRne8kJWwwFYv8v1A
qvfDBfSFR6d+8oVC1caIyOxgDCEmCVQVCHzSvG6WtYMCeYEKKNBtfqOMq8rM8GDZZOoi4g3o54rA
VdjOKpzj3aQ1rd2FrbkbNyXOOuktf+pf/5XVA9GamOOpcLiLncemrDGulwiF+BkAepPoqmp+i/yB
jDbyZZaG4wEg3ZVgEHGOCjjNoc3KR3ulpwOAvDQmPiXGOaww1lxrNJdP/iJDCWFux8ND0mXGWyWX
J4OpvJG0xrB3Aucl98zM1Vhw7oWAD6qQnXgWJ8cpkz/kL3jtg3fOfexB4iDqFJeseEgg5u79j4PG
r3x/H0c3DQVABgLuhmefStU9e9iGZcV6L758cheooSSyPy4/GUU4dNRmFEKXReJyY4OPwb5QvSbJ
w4uKDI2nBAqb/nblPyC889aPS39S73oldGOP+b0i5p8Ni5HynH6DyQy6AmrovVehlkbZwE4dSDaQ
oWsfSufKNc+YLW9VTlA4R2lSvriaBsRRT4ij371LacU3+KJXPRgFDlLgmGHTBcTjAmdID3sM6Ne8
xHJvqEcjCh+zxe/DNWDp4zd92kEH7gbPIkxQyrjjLSKmmYcktzQiQpQ6u4FngPKBFdWRwpSfWD5S
uzSGsVRFD4OD6GPqTDNMHpvQdj9Ae1J6D8AuWZH9EnDJWnFAFmn4gk85Al7Trq6pk1tInm1VB1sy
GDqU6QnUP1WCXUusFINvHdIQDHvrj07BYqFQpwUp3GV0kZzAoIlNxulWI3h2DlxxVYnGD8jiOWm/
985psgDdQxug0/4HRJHIlL6S4drM67Rj5ulRU9YanbU8GZ0JEgDng4TTVXft2jpQ1AnNf3PNmOBv
1ahgakmGaClSBY60yoCaThJecei1agWdlDqIf7OWCjy5EyeZdQceWVBZsdkrZt9C2+kX+7Tw1b4+
enAsmgm85ML5dr3GPQ1l9qIgejuJaQLVmtMqwwUYMANC5akgVt7Wzn6stTf34A90/3+dFkVYm5xW
qqGl1llnYdvPWUxR/6/rLA1ZsFK15EjTF+/SUkdrbFzjRUCotndocBDC0e+2ygVJpAfu2VGj5jpz
+MKAK5G08YXcNRJQhOqomaYHDsu1qzGCRhfLOOOXZJt8fL1Lnn6J69bPRjIUvLu492OZrL4OVgyd
ODKC7S/2/NR54DxpZ5A1vF8rLfSKK+3SWJm6LgeMOs/NbuGNhwJkOuDQww5mFQg2+E8gv/trlquR
AaYkF63aiYQUxz2Mxlf+VApKLSnAhLQ53HTdkPnM+doAzILhZyXIyQuFumzvCurGghCwZj7ElxxW
vbo8aXrVlf81iNKQ6ROBAGRARng1VciVBJlabpsVXaMXVKiKROdQ58fnr6CvGKo0OzCvSZwCf92i
CfAH8Y9bJKVw5fu9TQmdB0OXLbw3mpRZQOWsmEQIvei/ZCwQIaI91KtxlUCe/1LjHrf68ZYBdYXX
EKv/i5s6vHL5SW8s7SeqTSLICrTfH1Y68yYD6WGORjh/uKMF3AJY/Ahw5jcBtxtwAz5UaAHgpbiQ
B9v+nCzIecP+FbSqHjNGm19jFTIFt6/0tAADFKhGnmnoATVuoy2OTbWsV5nVxZ2m4eE1nN0Wx9Yy
c46kJwv6mF54klA5HGbaToN0r/ad2k/1XTXOwhApBzUhG216TMWI7WpVEx6N/gdoooyTlZ5Y+q4M
ozm6xAE7zYwOfWtPi2keKS9H16x4punlURBtgnPtx21VDvNr0lBeSOuw8wubCylg6CaLL/qT/Ufq
aUdSbDWaVUcZ4oqqb/3sGvlXvSQlej+tyctB9G+Ca847P+uG8BYkEPjyc+z/AmhtNl+Nj8kZxLYm
Xd4tqhbHift8eLKV7vk7gU5ub3h+/ulc9SikMQdqFTZSC4FEBuYqKOLFTPoZGJrsXnrNPP5UjCO1
BOx+Rlf9OBD4qGVQcCJspvutqbgz/x2OiU+TWT83uVMzYklHX9fHP+/zvlrS4uhrH3ctErbTAGyx
ATUhkhDmEPUCRG3twLLyEdMxsGbmOIKkJhWUDWGNWX/BLu4RkLDO50k+GWAPshiRTM1cyF7aIMNY
jJVlMys4tXhM3rCLpVeqIxHdigpZSF1THqUq1GGXknW/YQitNyXotCXMmlQg0UFC/yuidVlOD4jL
ql3Ul+sTgNdRjbmzLyI2vsncuxs4ZrkKOWudiHm7oFKNvrhFYcWsZxTwh40XDQYFog8OvUmZlv6H
KuqZskUP0ouxfvTBbF3/QdPy4D2ULkhFBgrTFdQ2IIOLrm5LI7ui4Rg8ipa/RYYm3tJ9VqKcK/S3
vi2IRLbuu6c4HFGRdbYAN8Hb2/YsxU2dXlIfNviyteoUa1yN7ZKAXwh1tmsiCwPDhYK6AkK/+Ik3
XO9xDZwadY1zYQgvOGkrVOHu2PkzEkzhJWXbnn2rwpsUAa4kXKOx1h856heAH/8/IS4gti45NHUS
XSnAVHSY70rD6gCck6/vfd+XVW/3s3apvkGGK7BdhxEBdxQB+do5pZXsz5Y6AsBoFnVrd7ezGfYM
ktGBgjS0Aihy/ZYcl+PFrnN/4oshAdImiQpZegwDRLOkZ6ZhkdZRqCIAmA35EMaoqhY3Zm+j6mRa
ryY0ZyQZpN1dg/JITnBFeH84mn93xl8pIaS9I4K+cQcLHTO7/ZVPqtIyPsqsQvLelzdat32wo2Ra
fQf7gP1ojscmiEupuyRu+YC8Lh3CX0KdsYLFmTrJLmf5G675aNuROAMLP2uK8KCfStMVDf8gCNeg
Gahat/EdaRKqQGgJbV6SZ4amtGmFECw2gMeSAypv/Yz1M8vTH7TZefwk/hmBwscB0VQqaO7Gk89B
kKLgVxkp/V6jQQo95ybv16hsFLgj/BjppapjrmFh86m5PcmNndbqq071bBGEMRYYkEIUtu9ZYEwj
E8krPd4h22IU3UPxskQ9ilpnwHDLilD8ZpSQ9/KK7C6D8QJj9H8ugAmp4O3jHbZLs63SXf/aP/B4
av6C3ZY+CJDgBuHNEuN8hYtTwai3ppYBq755FJBI4mFpuPk+W8b1pw+pJWCZGjjSAz1TgOND/TQk
ZALenosYlM/WCWApYynpLr0Y+DpoMa6TGio47mQq3Tnvam9VaUg+XEVixz/Fr3aXTuB6s6b1JpH5
DUjoGXMMf1Oug+iCRXwILj0dcEPxUREG+GYTnnlB6Zmwh/gQK75tir/gv/AkXxE35Vcxl3lnXI4O
AeM+J2MU1tjXwV6xh/ZM7q6zLUMT6f3amAq2wbjBkrXwEMqEgmxZ+Bz9rV71bDP6x9GhInP//8x0
MlCt6guTvNqSzsu84CR+/pKhawA6MCJtC6RjE4XtAIpmutKHTq+UjWq+oUePN+ivcFCD3gulMmUN
OXCVDhhyve0/Qx+D2rDn1nxhQoUgIuot1mb8jIiVvHxI/JkB21sbv+T9+yNrvFSbwEqxNT0KYo/P
YThAA7REbyoV5lxxoXlsgYcBceT2w0Y50wSecuFgWb70mCymxI77EnmN70xa9m9gW5fwQR7ee1my
yixpJMMDjtwGzfqV0J00W/ejZXR7N0EYM0XacROUsnnZIiFVZdymb1ZAzQM6MIpyIqH0jTLEQbEP
Tvd4hzWPbjqJY0obC2LT/SyH8sX6RaRSYFuPnG9JiHcMs9pcUkNMVntBzliVp6hJECyMHB3RrxeQ
0C/htZ8v0DIooCKu18nZ2WxXHLGb1f4Hh1vDhJ+JLboQKFBpcXatCr9Lq3kmSX9YWtTasZra2xKn
e/YD22BjTbJ5KcoZW+n4Fw1J3phnHMypIGZk4tDc2NuJ++sLWmamWrzF5zxxZ/PlwQ4zMBG+gsVG
Hz8KvGh/+zn0o7ZtHz4XdndATNe8fq4q9b52NjFLNbj5g92hPoPNhfpHQ268MvRuCDeHW3Lb8YOt
88bT2FtghfQDclHLKfZxXJ87XJqMCeuPNahtsGCTS3SQzsdKhjN/owRn8QQUQzLeh2X5Nk5FnVX2
MHf2UQqbMitwowZbGOo5TS3VrtezGlTIXe/eaqLJhkPaPD1pqqpP8YF/wb4qb4VZ6r9sYmcQRP4p
RyVooyhWesJmYfmp+c6ESJ4dPMRVN3x+HtXmLZu6wP577RYxqZOHlU81lb5Ht2mLQu6dcHq1we52
F/T4YB/DFbATMWnEpwCCXrbLsOrZILlsjYug7CaHfuQiytnUfepdgSONOpzcgHrRIketm69v0p6o
EpUUhBELRO4Mjr7uQuTDXvYjL289r3DntT1YeenADEWf8TK7W5vCzoIG8RS4F0CHXTCSnR8qt0zn
PGfFNuUEtSbKwoeD2KCDFTwcBEpeV/XkJuOJvMZjqLTEp+PMjNtluQzuRF1znqQmjtC0b3MyrgPf
pcdaa7QDkFPpHRlS3+LhiJBYUnP1j0WooJmaxzaIIUF6M2+i4W/YWGTQtRQvwUssWKAHM+1L5tb2
OpHdHz0hAOSl3M9HQqZQKdGdFNmm6lkywc9vVpMzW+hhNUaqIbuElcEF+Rqjq0SdXMfHuAklOWnb
PV5WmC7hp91yTTbyGxp01JgwvyklB5ksvq9RLyTOlQ26ojzfUQ6qsEDdwnJek5N9CH6V+pZ6qLsX
SqUhUqL/lQdSw57cIbDWS6LZxAnqVQ3dfN5dEmkjV1CvQEvM85lcngWLMmfZg99J7oDfL0WI2OHa
KeDVNnQjBiD3dF0zPp8tFmG/JOzhJYRhpg/l9DZi24VIscKxtIdEfX1wHgoi5vh2WKwBdTFG9ubN
FBq51SKQHql74Y4Oe9NSRP3k/O1tTEQzdYvECZxdzPfMi0pesi+vRy/9ETXutGlEmXBeAe7e1rRy
2mxIoYBz+ANA3hUMW53n/UKxXQDzf5tt5XtLjYIGZHC/nXfS9G2uhDGcVthTpGJWOFLDZ4tPWxvs
G4svwiyDaqY67xgSJC2Oyoznjcm50s3pujeSfHGoOzTiNKLCIYFMZJeUlo8zu2qi4Zkufj9wSUmt
Px9REu17xXmgfryUlJSWGfNZEST/rbH/Hdj5krBx0ysuZq59U1JtJkEUocUCPDoaJrlc3I633S9n
pmmppVDLbIthAkdQ5DoBixVbaQItdu4c6ELF0PgdmOSpKw6FP313QBNyfJoY4KT/hXLbdZsENH2k
5Qr9Vk2xlhNuIBMwNQT6tvsc3Zrvxt3WXXm4kEeeuKy8oFLicj7616HzNtOQRqUZb2qN/Uq1CnnX
hV4UspkJPIAlq71NoRj+fq1Ra54NfthnoMk9IXwGGNcghZAG2o4roOBKbYAQXe2bAV1ngjzCN6il
Xj+Gqa13TC5F2qTqz6vmbMTi0A9QdNsTU5LZtM1clY3GHTyviriIfQrtThp1lnlwrsiOzUYXSiiq
WRknBhpljLgTaALwWuU5DLmoWg/Z4cI9ylD+HwE6zawheyiqLBAU+O3OC6mzniYOnXDCklYdEX23
1vXIRR5K26NHkepDK6PDwuwpELUb6pacWPSgSrhpPdkkZLJcfxqZAv97er0FVTc1R8RUChgFV6Dc
L6a2JBLA0lueTSfXLdbQC+xqAdd1roRVVmU5YgvAscQLL0KSVDbFWB4vA8RVBHnt6iOuEB1F9GB/
MaGgXpnzKeboim1BLBwMvy3WSGEa0LErCfWbOhOf/czMFYDLV2Sf3rkERxsPdhkSFlOelfNd3Kvz
obdza6GyVlq70JtAB7lrAjWN4CvwfC9v/bE2ZvHljU8QPeOyU4iP5ZFZoeKFUETK5Bx6CSWqIULP
lTn0vQWAEMR8u7Z2zz29ZNtqlg3og3RoeNoxwOIVl10xuTQzPw3JM3LVpEWzc3Q8Hu8M24Ga9PHi
P6JJne3bfC4xzcpzLY04HO1TZHxCaK9xqIkmzHHSI66pYmUIwbqtni+xuQkfaEjhVJojJVJwPEt/
gn+J2Bw+ETp7qBiSCgHjuZ7Pti82KhqFF6bSYobz5QR0wBI0MIElaJ5qgL/jHmGYmi9tn8PVHxlW
8SO6ns9bgthU6O8qJVWe3OWq++m9PleBMa5koI4FYMGkKuG4knWa0nqR1LwTXiIl3/LTEniQCNq3
rB+dfNYX/k4Sbn1yGYaJ0gzyEWH/Mab3RULOzHQb1uytFGmKqNOwpDglMWN28pp9+asa5KVncjZW
S4qaVB0AuazUpTfF8SUC2r5wm2Rn7Aqnq5klv0LZYM79tEIY1yRBwDWvr7OMVhu8wHj8WXKXpMrj
KGDj0OL4sqHgIM37H7Y0RMCFP718d4YYCZv1UvyQU0/YIj7t3YEszgkthFE9kx5gWw+4g1z2jVMS
DL1hFxpycFZo4Rhx2PlUn4BjemtNYXdShz1duOInvo/dI+yJ7hzWvfiBTHuibWQvcNHP+gdwUgpF
AyMwh2IaqoWkVQYumHV4fof8xW/Gpujhb6Xs3BEG4WBxT2zHsq37T313qgi6rLnZutr51cvlJGpb
kOt6N7IdLgl4LOoLJdLZNNxrxpNQcoP0o5xYq9RuFFLtAqDGPwVBWOXsSmTVxqaJiEpchEWC/COv
Jq4asrKMYUTPCh6O4PvFe12Ti1IGuIijkOItWvFEYdYAVCoTxUo7E589DJIBE05JLfNlHpWHtNkq
+tXAsAJlHFavk1CGsskBIpC43OxTaengOlu0sfIYkTDdSTd8p1hJtAXqqwKiWAajpoW1zvVEm7b6
GQ/sE12k1jcR7odBuGw8MiixcAIOJY2vg7vN6ezqGQyfAN7ZitqLpkt9zknclafOq5qSZSUApCDl
6upG6iX+9brn+VJiHV388gptdNLXhX00qaFQ934Y+mniGuNkBP6Pt+5nGGRvBh0eGXYi+qG8ObvG
81OruRb7bdfhnPV4HCOqPs08/xDa2nS+dFRPN90EOYkAv7uiL2f57Cfz7yJ8ZTTAnTUmI0moQwhe
fgEt7BhCLRVKQYnbUuvMEFKi5X+qjsDrkG/HfHlrhmHF40WZEiGLqtQcqQffysetKMy9gs8WmJ3X
PY4LoCZS/+uOmLy6IhNciO0bTcGDpqZPAu0lX3l7r2SocP4B13Ojn4TeG63Fl34NWYtopH1Lg+M9
a4jqKeiNtyCIzS4GHSB1755WsPOM2voehnOQJMvI8yCwH6uuKf/y2OXrnwvPi7OTc29DBCPsYQz7
ogiMvITXF37j1qrQgTH63ePZji1eZcJ//y2VLhFW+UORae0TbGm5ABi9N0CsSxCpg/dnxASy7CY7
6T1jLKpmTHdDooybdlZpE7t0wwvhXO76o3dhBdJK6/nkZD4Cmxn7SwAeRL30XtACSK9ydf0oWhI5
YonHsBSbM811ZS3SbsdfEemGTQnSJMQPrBpExebSxUssvQhj1aK0OlD+5BiD8Ouzflw9i0+nHR1g
WBYTzCPQB7ouSVBJNhThwM2NBSPZ+vZwVRS5deLBLXim35urBxgLjyrbS7q23FffbgbxR5N5MevQ
ID8WpwD0ex4WclPPeNH+T3jng1cA1ck0PvkfjrlFqRgNPAvetNrD/Veq6GwFpUB81C7J2+aApr5a
OXYK+5DFrlqpugafrcizBlwosrkhwlmqyMs1oJhIbQIG+We1/4RjlB5teeJH6CRIux6E9zF7UjXW
IfgYFTxFn6RJ6wus5EmIc2kTMqjkyYYOcpkZxNWPhBLvY5V6dOXPMbjukD3QDyTMfJ/0uCsjViPR
2QF1AZmhknEqGWGNTVrU8cV0zJgn4/H91VUiqDF1F6EPMKf2rkmHExFwc+G7YqPrQbs639RYQjC7
E4VOdxsEmB4EZ7R5e1XMCcfHp9NHwyTB3Z5opdksLHaFY1OMyz5bCaWUwPK8jpur3AqVs2eJw2a0
2bgBQzmuiY3a5R0D26SIj1LaVscuGr0oD/hnFcg6e9BfcKRWJq6XawaNLMDeerTbF7ZXQ2jfFdKW
DTLuFuffNRjDVw7ySoLMNCvMAhID6zI1Q8oJO0JRAFDTb5k4MfmllfR78NvC57SRVE/hb5HsAarX
gGSUcchd/gXtl5bfMXn6UIt+Bg9WI6B1JpkNTPf7fJQh5e0xg24cEdkCNyA81LjrcCOk1gFmG6jm
nYxQyTcNOAtc3MF7cYbHDNJDjXOdGE/AP6XygibJGs/ghneJ30tmvSu5SSWkms/uIjTNJUTqF8vF
Td8aiq/bRy68uVWjXiRW4M4/7G6/uVD7nacav9jeiOUZJlFPfKXqiNmmD2p184onHM14+IzhtCiI
JCwB/ahdwFf43XQKKBqXp7VOeAQhXA4B9qJyorSZ+iMkUV2Q10PicDJh8TC6MMVFuxj8LpV2EN37
IKlpTbyYEp0JuFjCOh+GbyLoLke5a5xjkoQBB6Ypj4f5d0RPhJ+Z1ZrwDYH20u7ahmroQ1Z2Hwl/
UYM5iYLrfoVS5RW6wE8eyNI25/N2UQgCmztTnf58GXyFLFDa+QsxvONNqDJh+KJKQI+TbVAauIkt
SPGHNTS6UM9DYKkwH7cOcF0R6BeRF1KOH3RcjkYpTe9E/l9NmPNUvi64r68okR8eWSZdeL10colT
Az/uBFxO3OOlICMc2WvPYgXwbIBdMh0w9EmPiguu/SVMuLrB1iv+aUyU2Rytd6/r/VYXNUVeTBxy
wYVlt8J4meyv6xQ0XnF7YX2zGrNpzv5wM6JLh8z5xaE55kOQhq8oTPJ8oPnMtLDmN47sZ3gEzz/p
TRRDA50QQEL2ds+DquEALgi9UG6HePv0fB2hVWgbCBqJjBdfXOLukYdYk9aAlzU4ZKW8F/zOidS3
D+YiJJEwVrZsZcK38H0fzYRNkISHb3XDgAGCwYQ12WjowrPpFCz0AOtxp0MaxC3DIBBtgFp9LLTV
Q72V6+lcrn3I0hEhM2+8seXdOY96Mz3nTFZAHKrarIzkCm1Rls34Fh3N9kKI0noj6/0UVFEhf4BY
5xS6Z9pLXvX9B5GOulvPVsf4NPVzg1ZB4hpacwtbnLWzE/fPTjQnOpvJ9n7Dll7sp63MDmQ6cZy7
0YeAOXhvDKEvaZBsEfR0ffsioK2aE1lP1phnjLxBC4BCF0M3EVgsQFCMx12jfvgx0s0T6vffKJqO
3TWwplM222uMrQP27j2Bij7dSpfCAmaruY/bJsGPliyvjGgcjNISIMtWT38Xdzy7z/LZpTFKmI0B
WfFJ1uVOECQeB5ukNiPpvbZQiYzF6BvMhRvXeK5x9i57Y9Mw/GQZB5J9m0PbWu8MVhOq9+qtfjxk
WL+m1EL59KDB9D8igk4TTsrJzbD+i/tQbKQ1qWOTMc/YHT1/XRGSB7Bl2at1srXF++FUjIaXeWjd
UmqCJD8JZ+YbDtNSrwdAtyZ73fWg4K274qhg5HzsYp9ny2KOKfx9OQhG7UM3VCygS1PKrzwtMZBN
43VHTCvK0AXsEqy/15j6Qn0whLdTl+UpuXmtOFS/Ja0ZSJ0+S2TAN2sHhuTizXIz14quxW45Zdo7
TESRQdDKdCNgn8RL3hDdKSsluZYuiQjkNrygyKBjbE/OJkndYChTbeJ0ZGWo9usHLTZfa2eAQ+bH
GxvEUgHD8W6Xxki7dG/YNL5Iw2U0L/tm7A4SOG7F1HZZo5f7FYWTB9w1cH1/A/tg6j7GQMY1pzRQ
2WsHxZVkegfMv7Xib9sAGnVylUjah9aqgT6of2q82WlnIezDN++6Vz56s6cNryfI1f7qLpLWUsP0
6sa6ydJLG265QaADhs//ohiSXcc1+33IpYctZb+goODRs8HoYKGdFrB2+WdxSlubOS14YLONWVgO
A1vMHabIDwk9cYny6qO1aZTjUSWnW8j8K0XayoyUxAalvnB393FSqV+31bc4R2QKQqEWT7iv6bNl
o4vIME0tt6TvJYB1RumtIi1i3I/fgjeqE5gRcYWccJPv6in16uN1UZrMpSCZ9lESeZZJby6V5hn2
49YiT0jxQ28q7d1u+TUq+whNaSyawNOJViH4CMpshvvsiwJq7oacmwCDzkDtBLUJfF/ObkR3A+L3
vuktU/H1HCfaqub98U3pi5XwwXAevWPFr0eWLWe09MNPZNBFNuj/fURJtJekB4BODh5ErIEByKYs
pDo1zWpqlFV02bywB4x5kAlF5GMUaZ9/VhZwAuSw3iLXCLTPR46szvkRugBTruMQv8nRgcRgp8UQ
4L324ZNh4c24YuEgRHeOHjhRAyGPUFkwFlIemulX7ZP+3YNRjZ2/xaPZMF1TB9e6QFhV+qkZAjff
hI0R11mOqFOTTcSf4cNKcjl83rO37/zPXkv1Dx+DpCU6ajS1699FOUAWc4xclUJJpVnNYqoBTvNl
4jmM6OyaVjRwl5oQ7zRqespWgY9NZPFjKc89xylmcKkOqGRwtZFtPmsjac9xoJ/XSMNlhPYk3Tz2
wn83UmLMEjrsiqlpBISU0gWJGGtNaDYPiCkazIoEhntoc1LALTja6dqjIi9/Hy2G1RvharLc0kEL
9v1R1wOYc5BaaJzNnjxA35hqOvxK0gJ2cRC1mA99x7XINuDubPlLVAw6f2NgSPEZkW1l5RtvInGI
B1MkqcjKsEaa+mQfx6eAfcIQ925UbbIiDPPtPpclmZ+2R+ezDTbh5npGF8OJGDSeAlDsML9ZsTub
mXqCU2J2k6RodJK9OGVQFpGRYCvlCi39aNBDhaTNEgclyKU5IytxBx9BCI3ksx3AHPx1HXgWpaI3
Ns0JQzyEbH2jAZhIjK0ApHKQFcZo38bN/tLWk5nC+I7jwjEgmj2CK/lD0EbQDCDuDokiJIUZAJO7
96G+EscpsHwJ8GJbQNjiVTu3QUL2Uj3Ifh45Ve+3hAFs9LFhPgQrKaUOH5i+juKO1evWZPQWWwFB
kvYTmTOR4v+QINw6eNBkX/u54Yvf+ymlyhd/RSZwTJuyzQ+llGdBfskaM8vlvDgQh3zjHIpi08Jl
ayjy9HGZOnvaxdCWiEW3dQdmgYOXXCeT00fMLz+oiNi2CaNlRES4V9JPj0F0r3+WD1/0yg5coWFg
8H+H8Qm54qPc04w3mCo1rbe+nQpDkHdF1i87PyGS267ifniEx2TpfEGSMQ6LI9EsdXZVHo2nTKIy
diGmRfYJCXmNmEuAuc59T8y3d+9chYwQTX2baDXqtP3ti9emifBY/SrmwpXnI6aBPnnmTVSSn6Ip
ZjFlohd9QtrQoMdBw7eevpdMGEnq91EqOg+WBUEDgh4Uf8dDbCDv2KRUyi/LIHaHCDap2wlwFvbk
qBqPhK6zfXhjROZ7SI4VQZBXni07302eGTDXuU8KQCSJprgOycnlWXUR6DJdhN6xDYllT+OdDRpa
u5Yw3ryMriYQUa/3V5TSSnvO3J5kwGe5xlZg9QEjuAQYnzWKe1in3mpqF0Ac0OIvAClglHeSTp2m
ILxd5UjRC24/9Db3r+z+rIsJGqRVY8+LkXUT2/um4zGUCGCpsYPIKxp+P2taHTw6Jl5SujPuWvGJ
83alsH5DBUpoHqc1539A2IlnH268erJYGM7LKu27p3lPQPP3nXmKTsFWtFGq5yQjE0wbcrLMRkKS
0ArxTKIvmBkAg1iBlfNLorRKhDCU79gSPA14RhCqDdLpHYaLpxKwVZzvz1olUsbNyojFlu6Ii6Ph
DOomB8NtL2Iq1onFvXzX/FXLJ7p6hrPP27sPG6nkzzJBWFZZc/KithozSwGXgWUY59epzu3LQSuM
dq6whjOPdv7qB8zEucOTquE7I+li3QfzPY/710K+6KCloUWa7jUXmJDn+ZEUTCJjCcC2ad7J06ZW
clr1zoXG7tg1/E24/AuTTFVrUdDczgXw1hpYHetOqw7I11WS5QNV1mhdCtCiJejvrkA43piVLPxE
Xj2CjyTQrzsCFQiSs0dzgvFE/0JPI6BjW0/TQIjN5LuEzBYKAmEpk31//VcRAt9eqrrijtNH6fzM
rUb5H+6Qc3H/FOR0WiRt+Y3INs8nkWD27JYtMFj4EJ9xgBjKZR+FyqjNA481HVgKN7kmz4+Lq65b
nsr2zcHKLtMmVrctCTcJ6dIAHfnHUvhLc9SzWt3Q7qL3iHeaYtVm3D+2L0wSRCN5kHVeHPSxLT8L
1yIXRWjwecKt1U5vjUzK6A27P9hIiraEXxCSc3XQFSVgqFNfXcfdoCJ++CtwwFXVxSm4rCr8xvEO
+6oJwcOyuH6e57fKtLccVfiH7kmcqnW7qbmk7O4Ts2pwwKm9JofetJKB9Rv2seKa44pek6mrTlu7
+6sDqWE/49UdifdBK47if+KwNcqcmas0SuBsX0vt37/sa/BjTQEqDiCPxtWkjYlotOa24xxaV94X
G1b75vGBQZO+7BYp4AVALmtXYxfUGPVU2sEIKRMD1TI/wwOpCXdR5cvsODyNdyX8lr3jdhWVKTS/
yCwhZUFdGe0gPz0aXK8CFDuLKMvT3/O2cH5vKQR8//bm5vcgKYfvgjPuo4GqoqaiY6xVI3t2jd3j
DkoOzDD9V4dXXeYJ5LZ7BDe8ojo1ScPo/1HYYRO4JddyUICZjPYfp83W4/iubFDBWHst37bjPlVe
B+kOiqthLZyviZkRISHlsSnU+YUv+8RqmlRvKwRw6AEi5PtgSRJd5H2jqis66VL479SDRdUiOzdn
24RNxcVA9uLZnDvzzxfOagcaXHozO4u1HFh5hOrQPQRU6sUnicp9m0mFmhFeZkb90fdo7khiJhU8
kcBw69zjUSemZB0nBAD6KQUuv0OWP20dhjMOblnjiuzV593Ujnr49mfFl6JDV9PPWkFFv9/lmmf+
nCw549M6wSkTdDEPyGGMylN8ZKtn5RGW+HXuCoSH6iZ6bPnwl/Vq1S3+L63H9iXDWc8Oh7uJpO7q
DbcDhsBPlvNTmiXaUI+ZPrsXIVgMRpbJi/9+EaApFu72uEMKFnUus+3LyDYo+F9TSMTbKdYHY56Z
Y0wd1HF6fdli02WWufTpyw41DLfLQ0PbUfmjZQkSImrc5UVVICjHoFCuda1qsi45/RtQ5ABgPlWK
8UqKvnlh75SGo8qZcxTecgdKJq3PyZ1L3ORvAHeExoP6Oq7I43+xt5Jj+3BR7sqTrwZAg9RXOt2s
wxe/hjxX3uSrAqzGVpmtj0zso9jpCTaNFUCXU0fSCheTfCXMNg1LEuxVH/QjYZuqQPgIZYNXgs3b
8GfmTXscH1coE6GOOSgRGsBk9sNncTbHE7wm0IAGMHoguf6EMjH+s4N7AfQeJZ1JABaOyzpkqWLl
vUXf6ttqcilK2Dts6fm7CLQWrMWus4gp6scp7pVtRa5zCL3T7W5vj9/qEodHSlEPSaRvU4IemSqF
pUfhNWeemM7Bpo4sSyg3LWxjYfLOqRRHZoHIM6mWT0iICooAFKd5iCc7/Qow1VV4NM0thawoenIW
Saz3ucqOtoYdhvsJ5x9+Hhgruqo884LNfCG4Jawp4srBcmN5fCO092XiHi1p5SFAv+cp8RyebOmE
I2M+21dPipFbOBU8J9lNA2mqnhtBCxYQRtf86jkL2/A3u5YkiOoNnxrwM0FxFBzllV7RKyuV2T+S
HKx6aPFwf94YFQwb0lAjfuNBxb8fVS4/vGidLe9sYeWgdBobqzDkJNPIpZ+5BhyyVSqCADQ4OmqZ
VLoCHbyyb0I/od4HEXyC2K6kH4EBUbdhIphhLaFDKN5a8ligv24/ygRn69T06ZUWaQRBklVCNnpw
m/c1X8O7YfwNeWtlnko1tmrsMyOXhSDhcZnNaXr5YvrQxKZIl3hwMVhMOXfWKDsO2SDUyO1ckmjK
o1qO/Jk5ME58l4w13KxGePzYswT103TeOZDLL/79cJw2lz893vxyCUPMvQRuM5BmoCJ46ZRuhWs8
AfzeqThKgmSJD7Ux1AU8tfySVxhQajA12+08KeJuhK55xvHedr2D1p602urxrDpSqpbbDt/P5wHW
U3XukmhLDSnQ2nSKFmG4tvd2TgQ5wJfE7CH1lc7VOCYWh402u58rEvbmocdnPqURvYA1U9YBqByJ
+gPMDNkFsBZq/yX7k5esY4xg1pW7y3FrOvBdFdwzBOMn2bkuySFGh3IJuTSi11V9WYdSCmLuGS8f
SbjxZ3t7Zfxh0SHx+ZcJO0iWIK6zMrE4xFxcf43ryOeADwnOqpRBPT9W6Km0KJjbZ7Y30GGQHMpl
3W0TiduQQt6JoShUFq5s/5K4cl9eWGgZ8tGf9gp5SzWWz9LaIaK8c+VsXkGDFq6CnVx3bix2e3n9
FaD8PxOU2aIKHbgRb/M2UI5IArIY8dbMZnNreao8dAmyYgPfP26CyN+CohmbQPOabBALYP+4HvIz
vCMfVvPryEqWdtnR4xmkjLo0H7TB9ZwCsX9XdBxECECMuQekR4Le2dzHBQsUhL2wvtFB3FxERDTL
RkceD0a+qHaHWx603KN2P6kaD2F7Q2E6fEXfnkFkAVaDBipfcE0oamJMQ4uVil52KBTnlQGZ4v5y
88szM7DOINpC2cIK+BzwZRtm43hGYlUpQ0Lm+0Eqn2whubSD9t/jYHEpfen4SEqkQAeHy6Lr68R0
odIbuen9vEohu1m6d6eKr7AgaAPDn/xEnL46Ju76Kr58M50GBsIRQyfFMI616ohFiJAoJl8WP7Uh
m91w8w6EKhOViBRFvrNhrYvtLh94tUOYhGKADs2DcWk4ayERWW4bk48oi86M7ZV1u7PkDx0OxeL+
I94PeATxG9t5LzJdEhXr8ZsMiY6xgVfOVsK2PD3vNFvx/I7fFDqjO0KCSNJz/UbJOOgu+axU2F7U
0LiZ7NGvoBQqN2e9Odfc6Eu5l7fC9Dk0AH18Vbku5bBloaA89m+ylx4AjEb9ns+RFmHaRTw7l5ux
virf5qfN85v6IRpyUk4VCfVW9KQa8G10gyWzSP5SJv6RplqDehzsdZX/CEg0STUJz0KSR2zms1YI
a/mqRcJ7eBr4P+jWBvGcvwDNBc+2eHSEWlatuOuFdOibR3HzrgC7SbyObYIssnChtT5Y+HSgjogD
rYDHbT3LIHzKgNiag9XDSTrQlsG1OEDAkzSdI2GOj0LarbWYgWpIMijoDpcpxO+95/UjVDKs/85W
FG3mM+0/ZLHmKq+OA5l46+An6wEsDZSpPMhQcZ5sCQrPs5DscUmcq58oETFXm2cwp7TkI1RsXWGS
Qn+8jsPtsBGW5x/jjJHu8/xkCp68P8mGs48nNvXNGU6hlFcfXNHp6COVILSq0unPMrXk63MfBaMN
JoTY4jtiUKz+GYuGECy6iXgv7XpGLyUnibfRxF8eo0RQy6qoVCupbtDnfNysL54tQZTp8LCGsD7M
9y7iXD66nzjYuoTtz3TmCecNXmsJ865OdcmtIWvsGRNZyTn+aiBVSD7yGF7qivDDvdLDitn5N6Io
ixnW9c3Ftqs/sB+yCb9Dtqe8SCpgZ0qsJWd8zkFNQe9r+evgjD88qJLZVWvXzFIZ4b4zx0ilnDk7
vLvBdDo5NN8IGe1h2NHeox/9/f7Ev+2lepayU8g7/PFLYA5nJXmI9kLUuza4cYWz770Vlu5oC8cX
YKzZLGszygAe3TFlk0bVa/Lpxww3YMX19xa85C6n0qK4yYqqO7Tz6Se/qgkW5Cu2jffsNty8Bz1j
p3riC4wyESdXBPWWs47jm4n3t84WZ4WhD6ymYg0DuWO4UuwNxWECEChSYLAU6f47V6KfpGmKwJaz
EiG2jkkFZaKl4OdmcfD6UZAG2B/gl4xelo1M/G7aYPW28P6IpOmEzunWvwjY5kXuUsS3+HfREOqq
QlW3725YuJyF/qC2EgAWw0kGNpuvLkkuho30F/nuyc91r/zJKRmyaZBjYluH2fcf2FadclLoZaqK
f2XI+bUlECp74UYvvOk2CKNvZ6TFGvWmphrXsTkOe0SYkT5HQZ5YhnnUCmDuVkyieN5BMJVtBxm/
72DHXFmZm8fQsq45ZrJScR2DWwbpqv5IxZ+Uap9ofRaegLOLOWSdTqpr3L15m5UcXt8Ue7/jJ6+7
j0idOkG7iWqI8IiSMUwwB+ce2RUNsrVfPeCfrZtwdlOm8kuidIC4g0tiXVqgxJugGw2kzinu1YQd
Y4MPeN3CzGZ1/PVeGI8Aa+DaxpfpplRjdba2Ktt9Zee+ZOi9SbP3ynOavW+7TG0gmH4JucrJtVI2
i6naa3IA8QxVszu9KdQ0qpT+whda4IDMin7zTf7WrABrYaBLlinCatT9KF94Q9qmuPPBfJv0Y90d
+gTFR7hK+P02FyHtv6PbYaHLu1kkYqTEhAkzXAhmkLlUfuJb/x4eZmHCEYZ5wogspYL3NydIEetS
3BV/xiSxmKaszvk/lS7Kmqg+NZxxEbsxKVi/qrddtplnHNNAG3Bgaw5deCMbK0AH7IuX4Qp5yJsL
Eq1dOps0s7il4bZs6Nt7VmW9UoW18vayBXxK89gX8wlJDSHPOepR7i/9dAAOBxrSKXATsJO3sGLb
4Nln6JBNrZFzWBvf99YnjdqId7MaM8VybYBwqsxQ9KyyQO0k5LDeD22EG+A7sz2Qa5BeGYc4yFO6
zrNvQUmw8UfDb5p65xQh4+qHiIt/qvLb4qgY8KqdyF+YLX/TCF8sylidAKXTwN11qoZJo4aFNvbC
skmi6PogarYThThesTIvXD9Gpgt426XHChxhS8ongdlIuQnz6bW86PNHqVNijEfSihbcyfVMtC4U
gQBQNc1ixo6om0bIJZFF3czOVa6vLg5yw9knZGWcnyrs8AO0tDU+edIq3pQyug/3J/mISZxWUVz1
3kDsVt3+mn2IylG9Z0rt0oAMEz6MioQQRewudGYoYpxK/APza5NcD1s26h7HTf20Y6T3WBbTDDc7
xrljg0hUc9Afv5Kfc8MBGdJUzX0+KiuDtJ3FHiSIzpa1J060mcHiAymj11NKtiqu7g80qV/F6PMz
968YnMBRxUS2YFPGdxe4KrIrM7yiGEd0d8Wj2Q/aUQSENdU73GU1bx/1QHN5WYl1uTrYiLisPGKP
zlF/mepLUaPzhHMozg8YaB1Fpa/rSFAiptazGptQCG7RVLubJwltVqe/36HR2iQg0XW0o9SH7C2+
dE1M4YNiU+1LK9oP4xS1wy3E0yTunjn912pGfr3DM3aSAsiMMcqWxdWRsaYsXdhWYmA90O1H6YLx
gcodTZUjCydqY5oXdhJuxw/pybh/1S1wpBUsX3h0KwNzOcnG9TKfEdV2dciJo0irjg4X1pQTlsvI
yBbIEjx/IudYExq2NGTFP/8nbSGTVB6V+qbJ8/8URmELGDkuXcVri7rXh9Dt8+bMTBC86hNLGsts
cCYFH9LGN8GtfDs6GLC63iFXyvZYRsZzVCHzlkh3nbMfvPW93CmLmO1gc5/Fm/63amsUe/BNFJqQ
5tbl/cdTVR5kgf6CfyMuRxtz/zF/cymAVSd9Nf4sJ4M8hhjo1hKdxOgm7ozCobCVYji2+KMedwtS
sSp4KEsTTZWZo13Y0bfDfygdkXLHcvleeF1FeEw0z/P2/3dGKgD9XTL7Q2oI31vqCCLRqZE2kWQb
8lTIhGBv8QGAQc6KcVKlR4TsQnTey0R5QKCGE5EuOgeG1napZMWpGAEuXL+OwRSUjmyAI/dvsJgM
3KUtKXgegvQBvRmKQWRrVmhJf1oOhipqqBfB+5AroDInTxUG9N3n75DnLXG86iCp1WIAYhYz5hdZ
l5+RNrs5KkuBvDFUYsgjY71vNJCEofSzkGkIdOPi2QgnBY5tZWCvQGY5+jqRB1XKlQku2BxoRyif
K1QG3GDMeON3kjCMbipwIrvt+hifrXDhTQsddSlLzC+yBlSgZY152/W1APhX0AuZy0IdoWoyQj4N
2mhQXuu+WEwTowM+Gh3Q+p4pArdJD35j5+od0lTqAeH6GdYJmSmZINS/mDNTCBfI6XzRhWJlLPWB
8EvyEIoex2VwLUI1Z1Ro36+8Gvcz6tKyKpOciKM/Y3rbpk+2r9Sa96xAWPvdc/WtyDmdUNjk6mvv
ugfAu4ntgBB2XFvmaSqncXWcnNQtdKMGK5BjdmlgEhOj8QLJH3N5RrieLGHAjhdphiainth4wzE3
+xSw93rw65i0M63BdCN+IsrwwZn9UJSsPNC+GzuDfSpcWxb2uFKHq4mgu4OYrAWfZfmP77bczMKT
IZSNa3LZftsyo3JNG135USTCl9kA6nU/4kSj2UgRGH9zlkz0x41NmQ7YOrgl5hY6c+rh1beGA9gm
VNXSL9LIPmON75YSfWbCHn9Rs4GD3QuQwyuQ0X+d9m0KWCROqMV2yjKjGBJJM+ov66URV76NZ70N
8PNi7vN+53nxUGpmO8IE5u9a/VVarwBF+MMxgcV2VimE8vEI6nTzbvAkIWkDzR+8tu/DiJc+z8wO
0t27H43/WEflxSS6HzWPNdY+01/yjopzQmk+vc9OsziB+mTXGA9oKRC2bFOb0f54q0WKJM1le9aA
dNPJTC4l9vfAw7Y4c9aTBHDMDQ89PLI7+X5oE5fbz5eZWg4GyPukiETinRNIB2oXnKg5sWMnQQ8l
w0lWgfZlUlDaINOPr+r/2Z4e7GsEEpnnLdAFuRUdwzJIzCei2cgCbFF///b3gbeBWdCtmdxCu0Ed
b7w036YocoUdWc2orygK3ZUDZcmLuceNTObebKrxnd9MzhiRCgEIJwzhVj060bjOcanRNW8IOZeK
62s/9vwwWCEPufR15kpFKn0aWCxa/m8zG6NMmTmjPL07D8HvG0gVd9RzXPf9LycH2XJK/ByAmvIR
LLTygGOtYbBusDE272izOe3WjQhs2MyXHaeLs47eRuujuHPKX6NCnJng11zDFOm8xXCxIkOALzD7
plIUqolYZY8ILUs1HrhZHcmF4NXhgpq7ir8s8qUgzpincYKB/SnUYCRkQhJw2+jFC1e/ZZeoV3m3
YSOvBsSm1GpmX1XIldjRr69uWqxF3jVCtwDWzNmEAYP/SNLAl4kJSZUNAnoakaqn59mQKX5/9U9D
IDbrtwJwCiCQTU/f1C/o3K4x694QrMWT5lhopu23b3CjEyAOdjpjo/q0KTma8zXzdY6nUS59BW1H
csK+920S6SwB17acK+VizQGXJxo7BytKfaGjghGicViSvVuVRB0U9wB4VcYR+6ldz/1DYtF0kK8i
2MT9Op02WUJQXsE8jjRKkPwLe7xvj3AZ508j2Y39rVN74FudTxvu1k5aXMnrg7t4N1WiC3bsy/Bm
Hh7CMf5YwH9Y47MiCyyhx75WvEg/R3TS+/ilPfL/OJIgYBc765hLAVDDPwJ6hsp30CYWfNW/PRoj
BkWcEhnV7W05DNG8s6wFP/g57RsAh/HH0LDVRMw550QDRosk+pwxSQb61asV2tkvLihTPs6nCj0T
fLamG+X/Uujc51cfl0M1ZpA909fAytaWrqugwZVb1q5BUH1tdmPKsL10ZWztzq6D+UNQVzly0cbP
STyaETi7uq2hleQnTeOE5VAHDsq1BCkYF9ATBKzcVGVTTbyqQRHPd29hqBOIpDcLxq4GsGCaw4uG
HIOAogFWAoL2f5CFdX1gYWH8I8JCVBLKM4g/zQx4wsQS7ub7mLJDhDsDzSZcVpj3NbmZpFrBeDlB
8/59+xW37piUjUkKN8CbpiSCM3IbYd8kCVi8GttU5WzxGk8IBkQK5/R0DyuVo24ws3u1N0q2aD5d
s4FzINW13nYNs+C1sc6EVzrDpiiAqO/O2RkR9c+BG4qSWkK/bWv/2hfIfVfQ0pzBLo6Lac0etI5b
C/B0oD4WtAHhL4nW2YN55HhpFH39IN9kwGh+h/XZAt5oPbS6sb6mEpmdFrbyAe79JO50T7ukz/vE
nRdYc0B4g2cFMTBzAMUW/Km8hpgrZzwOCU1YB7q9u7yD6AV5sheJAkZyKnDRsdYs8v7eYLDvig/P
BNTaucb/c9DKDMEkTfp2cK1ds0doI4T9BmROeJhaj6kcp7x6/mjVAsfBDqXo2aDPgaHqgzv9LMPA
wR6EH1BIbli2nPLlgimZifPkd82H7OA/+9YuAXgQKme5SJhbBJWraezHqJXAIK7ZR15nam4ptQv1
ABn0aWgJpd3n5A/DgM6ggSJOKnPbYhPZM3tzNNWF6lgN/NcVKTx4bVz/qFHnPdC7fbik5YyczwBj
Tven7M74P9gPallyZOfqMjfrQKnRViiLFYVsNDkqexKyHMHbbtDPT26LOuC7lyoBfZtyCcZcRTZ9
y7+G1PhM1RIaDEQ0Yv+79KNjo2RzdtdZTP6nAbUJHLQq8/IjjZLY/QG0pHJRTEjxA0BMMla852kq
GtZmda8Yjg4+RVMmhfA4JpoZhudvzNG+06HlYkn9o6bmRdqS9xYt/ZLP3kc1YaJ6khkJIbdhmFxt
q57jh1j8Hns9BEI1Wndf96TaEywPpSJM1hYJ/W3RFfy77h/AtGtsFwmerCNhEbSqwg0P25XC8f26
fjn5C/NTIxcCs35ViXo+HrbTvf9fR8GFWKHcyF3yjFELAvjFUpPlKIBB43acwjy+7dOitDYwKzNw
G9RDgFMaays6USjVCVPBBvwajHitacIJi4x3YC2sBWwzozmhMlkUA+3a8XvQXKFEXLuennhOpHfX
8/1DzUV0TmtNMmei1sAnnD1c1d8E6qUcJZkyY66MuOpcMbCKHdHof1EW6LHnz+cGA55Cx8ysn/cs
YdmR2Dc//56anguXf7w4zpC/3remIMB9LhBv7P8LMV6UgEJ7OSZGzzKmIKhy6wNVWh+8kOB9kzm5
a/mfMP9mrQwvtOLSsRuZODQbjv79oELC+IOjYaREsfkF8XjsFESW2BPda+bmscGtuhhbtsV5lSYq
ONDD7ohyWsPNtGeDzZacD5XYkGiA34qZdRGttL4nTWNBhGBYPUZ5cvR75DgbZXEZ7S0lIEGxx2Gw
RHE3SaYdSta0giEiXPSFxU+SkQccH0o4Sqkl3SwlruPViG1EWD5XKQBS6yj2Y1YX7o9NTiONpfSB
WzNT5qaid5K/iLCtfUM8yPISXkb7A1PCLgeHcA0qbK/3Hcmx3SnwYzQRags0a7z/F1Q5Wk474Qg5
VDW9FBn6wrwj0bVw+XQ6LQ2WnwEt1oLW1lHrE2/fijMr3SpozgCcnOpgxHR5g8RoKVDUbSox1/A/
Wg2EM++6ooZLSIT1dAiL7cheLfwWEocE1stdCj4AO5GsT3H9Wpvv/93+ix9r0pp+83W5/7LdBPpV
FZvwMnWpNhFaF2+al9Qiy8zVcWdioreAC5Bn0YzCkX9QVG/FicCZcfOzwCWXhX4269P93zcTsMaE
RemiXuAY7buU0Ss1DrgXTvokmuuZRTSuxSVat2Thcvu/NerJ0qmyFDDR6Uqs+O6VsXi6QAcEiPQy
xAruVa6DImJyMaT0rrd6qodki4D/cvChpmusWDMLs/OTfMNu/e7BZ+toR7gWl+PWDiZ4oGpKBq7S
kb4TVZrd2mjr+AoC+0CAxGm/4riJ+WJJbWfUY83zjW9PIDpC0WTQfWpT6DjXbqA+mbI4htOODfSR
J71G0reMIa72Jbn7pGUrWDbmPFcHREWMoWow4vWDAIi741+/dX/tN0xFXdNutQv6OtKX+2povtfn
LTPvtQOkGbdWjtrKHQ2eYAEyv8sWOzXxjKiwgbjVU1syImgs9Y1uXJ+kaJ3bSwfCr3xzTRlxyk7N
4oPpqQpxA6hsVW7PWiP2fBmQSZrf9DyFkOGlyrz+fWxTu6RcPawLYzMQEc7mYo3fYtYNFA6i3+b0
UGCfUg0lPaqyXzUp+mVGm1rzTFo6kg1eKOCYDyQ9X0ujDeZEzPQI8Osyvq1AayopgXodCelfBMDE
Ecj3dEybZlEbTJqvlqjTDK8cXxWaGksUdEatuTx7vFBW76O9Akei8ATM4najdmQwc1uGLzEplZmZ
8MVIxjqhzYoiWYKb0b/aSKUTEYS/N20GcLnCYmtHCdcBxk/7t8ODWtVood+O03wA5+j4cXCJBNtW
hvbV99tgquJu0MBNJw03HpsNyXHWLkJK99iohO4C3SdQAZ1tjNZPZh8WJuRA8hdBHsvM2qCXAOCb
6K/k/SL9MNnTtCMmyzGUBcjsNHbgF0uH7PWeVHocfbsCgu1bUbj6bKiZdF7JMd0RyKVbfRA8+0O3
YIhdTpeW4a9PEFdu2HrHYOtNaCqe4Kr7Y4XLgTLTnno2YYAV5WPKa0b+1yJic7h89I/I47RUPi32
aDg0joCLxP15QntFGDBU61lAoLpPfVarUpINU/0B1Vz83ml8PSGtkAP5uZ9Nkmw0EaWwa6SBwKFt
IS0Tx82ZN6fMVMdWiHYs9HtWcMaiq3bUrt/a9A5Yv6f4iA11RKXcu54N63ue1X57QlulWbTyBy1O
liLGhgWoj+PrdKQXVkmUI4g57WXDx4d6C0tM9jYHBTnhOu7tDpxQB4Rh7lpSamgsMdHuMk8I3Qm+
iZY4VnKwrrKkpbRWz7zcW2RkHYx8/GnO2HEEKsaTmfynVZuluW8ADpw9yVStRQvBa3dsAtNhK01k
pBCPA5u+iMd5jcsJreS6ZpfxGg+Wzjh2/CJzk23hQbuLJ7hJ0mnI+qJ1T3IXCIy+VquXJ8K8dgHi
YrHX+EbBSyd8Xtg2x+pmMwUrkdoAgELpJCUaqVc9z0/L9h3fNx9bTa8upjedRl3njfwYcAUU+8AY
K4VfFP4StPn/EnJBpiNmAaYSHMLVmbgYWnz8okglSsRqdaJWoROwktRqWCkr/ZyG4a3Tzj6UInG8
MwaRyqvJ+CTTmQ7PN7wY65+J7wj5eZZIB1hABFt9et0G4Fjb7kYRpwIaKGRqT5zq+TRjdPFrzn9I
635qbDfamVtDLb7yHUOw2yO6pR66939F7QiDmFDUELJz4FOnh4PYRKgsXv8Cwo4SD5Ji1U9atMII
J39DtDT3BBTSHX7cbqfpzg0YCkdoZOikYZo5ABD6R+WcRzmUb3ezkB3Rw4nlUfxY0c59AmMZ2hHK
uu9eBN15keaQHdq7sdnXMCwCfVMS4+5Kkl1ooYuVXNDxYAqFXMLUvOLeKJRDPhH+cZ9YZ99HxYGD
XGCyEnGZCFtPtvzb9xKBl7TrdDHw0O0tyG6lO9qPFel8dSDZLH/L4RBAFHNBUYGdKKf+xUzSZQoV
dJdS+xsfMnosrhE5p2HsPDfGmuwGFny7ytWFQNdYjT9c7HWfG1iC6IQOqXLGwNRH0mkIp4w1EthO
t7PTMCfWpwlc3ys4I2nfOTclOZgOPNv6id1iT2blc99UFnR6pnvDPqL9Z7h5ZFCn2XrGpTNl4mjO
vmbVkmZhqud9gVcNNZ/waXZ6UeVTFTOytZ1cynu/s/ugnrlMWiOv20A9W8Sw6ApuVnKeA00FXVh9
vgS2+pjDX1CjYlGnmuOkIKSTMtFqb8s32oC4lP2/S/Pu39e9htFMXF86anRN8JGpwu7INgnBD5lc
SJugCmj8QYR2LHxn/8cirPCMS+0G4G4yyy1a4o4ZnSAhzaqDPbnGR4S2HcDaB3YordMihBbYJMri
hDns5q9WEKBubhz8GUvR
`protect end_protected

