type ROM_TABLE is array (0 to 255) of integer range 0 to 65535;
-- This table was generated with mat2rom.m
constant colormap_value : ROM_TABLE := (
x"00000010", 
x"00000011", 
x"00000012", 
x"00000013", 
x"00000013", 
x"00000014", 
x"00000015", 
x"00000016", 
x"00000017", 
x"00000018", 
x"00000019", 
x"00000019", 
x"0000001A", 
x"0000001B", 
x"0000001C", 
x"0000001D", 
x"0000001E", 
x"0000001F", 
x"0000001F", 
x"00000020", 
x"00000021", 
x"00000022", 
x"00000023", 
x"00000024", 
x"00000025", 
x"00000025", 
x"00000026", 
x"00000027", 
x"00000028", 
x"00000029", 
x"0000002A", 
x"0000002B", 
x"0000002B", 
x"0000002B", 
x"0000002D", 
x"0000002E", 
x"0000002F", 
x"0000002F", 
x"00000031", 
x"00000032", 
x"00000032", 
x"00000032", 
x"00000034", 
x"00000035", 
x"00000036", 
x"00000036", 
x"00000038", 
x"00000038", 
x"00000039", 
x"00000039", 
x"0000003B", 
x"0000003C", 
x"0000003D", 
x"0000003D", 
x"0000003E", 
x"0000003F", 
x"00000040", 
x"00000040", 
x"00000042", 
x"00000043", 
x"00000044", 
x"00000044", 
x"00000045", 
x"00000046", 
x"00000047", 
x"00000048", 
x"00000048", 
x"0000004A", 
x"0000004A", 
x"0000004B", 
x"0000004C", 
x"0000004D", 
x"0000004E", 
x"0000004F", 
x"0000004F", 
x"00000050", 
x"00000051", 
x"00000052", 
x"00000053", 
x"00000054", 
x"00000055", 
x"00000056", 
x"00000056", 
x"00000057", 
x"00000058", 
x"00000059", 
x"0000005A", 
x"0000005B", 
x"0000005C", 
x"0000005C", 
x"0000005C", 
x"0000005E", 
x"0000005F", 
x"00000060", 
x"00000061", 
x"00000062", 
x"00000062", 
x"00000063", 
x"00000063", 
x"00000065", 
x"00000066", 
x"00000067", 
x"00000068", 
x"00000068", 
x"00000069", 
x"0000006A", 
x"0000006A", 
x"0000006C", 
x"0000006D", 
x"0000006E", 
x"0000006E", 
x"0000006F", 
x"00000070", 
x"00000071", 
x"00000071", 
x"00000073", 
x"00000074", 
x"00000075", 
x"00000075", 
x"00000076", 
x"00000077", 
x"00000078", 
x"00000078", 
x"0000007A", 
x"0000007B", 
x"0000007B", 
x"0000007C", 
x"0000007D", 
x"0000007E", 
x"0000007F", 
x"00000080", 
x"00000081", 
x"00000081", 
x"00000082", 
x"00000083", 
x"00000084", 
x"00000085", 
x"00000086", 
x"00000087", 
x"00000087", 
x"00000088", 
x"00000089", 
x"0000008A", 
x"0000008B", 
x"0000008C", 
x"0000008D", 
x"0000008D", 
x"0000008E", 
x"0000008E", 
x"00000090", 
x"00000091", 
x"00000092", 
x"00000093", 
x"00000093", 
x"00000094", 
x"00000095", 
x"00000096", 
x"00000097", 
x"00000098", 
x"00000099", 
x"00000099", 
x"0000009A", 
x"0000009B", 
x"0000009C", 
x"0000009C", 
x"0000009E", 
x"0000009F", 
x"0000009F", 
x"000000A0", 
x"000000A1", 
x"000000A2", 
x"000000A3", 
x"000000A4", 
x"000000A5", 
x"000000A5", 
x"000000A6", 
x"000000A7", 
x"000000A8", 
x"000000A9", 
x"000000AA", 
x"000000AA", 
x"000000AB", 
x"000000AC", 
x"000000AD", 
x"000000AE", 
x"000000AF", 
x"000000B0", 
x"000000B1", 
x"000000B1", 
x"000000B2", 
x"000000B3", 
x"000000B4", 
x"000000B5", 
x"000000B6", 
x"000000B7", 
x"000000B8", 
x"000000B8", 
x"000000B9", 
x"000000BA", 
x"000000BB", 
x"000000BC", 
x"000000BD", 
x"000000BE", 
x"000000BE", 
x"000000BF", 
x"000000C0", 
x"000000C1", 
x"000000C2", 
x"000000C3", 
x"000000C4", 
x"000000C4", 
x"000000C5", 
x"000000C5", 
x"000000C7", 
x"000000C8", 
x"000000C9", 
x"000000CA", 
x"000000CA", 
x"000000CB", 
x"000000CC", 
x"000000CD", 
x"000000CE", 
x"000000CF", 
x"000000D0", 
x"000000D0", 
x"000000D1", 
x"000000D2", 
x"000000D3", 
x"000000D3", 
x"000000D5", 
x"000000D6", 
x"000000D6", 
x"000000D7", 
x"000000D8", 
x"000000D9", 
x"000000DA", 
x"000000DB", 
x"000000DC", 
x"000000DC", 
x"000000DD", 
x"000000DE", 
x"000000DF", 
x"000000E0", 
x"000000E1", 
x"000000E1", 
x"000000E2", 
x"000000E3", 
x"000000E4", 
x"000000E5", 
x"000000E6", 
x"000000E7", 
x"000000E8", 
x"000000E8", 
x"000000E9", 
x"000000EA", 
x"000000EB");

