

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
cIiYfk3Xy6N5OP4pq3GmqGiiVNUZ6H5+UojetFJBvbKolIu21jc4BnJQVK6clVlXeOqxCwUuMeWy
2HOHrYFv+g==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
lIziGPDmnLk8lYYpZIaDaMbL8fBzq4Pr1Jhh0ulXet+pjCJLyV5jakxS1oSptZ+tHYCT5i9DwoXk
484l0YBwGxIV/F50kQ4mY5SmovR5v/32XWyGw8Sob1+z/rA/iYbfy53jpQjBFTMhONxMl2jPMKOr
8b4lWHN3CKPgzR7gpH0=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
htRzDc7r6AHMWLJSZlCSE/9tAboPhTxPArTqmJzMnfBntgIxMOX2YAPT8iZ7gZlglNlT/Bmc3ZIa
nj4bYkmP/Ed/Ze8J5Af7OuS/hLPfbdPEIMVOJrAzPKtgRUGYzZFakpIpDVbTLnXVCXGbnWwhbHOl
N+MoLyC3ep/1xGkMFlPyLgKVegokAfOd/5ePZ6yal5L+KR1ET32v4t5eGaONowzpG0O9uY8LtLQU
iVJDGAf4BzpePmtzOyeo5v68FfUFTjm1d6csF3e9pbQ9fEwJazksjJfyX2XYuUZH1eu5bhyJMU/O
c9/o5sfORhKXoxNo0FDKepouEYzneEXI8uuD0A==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
FHtFxX6m7YezwdeWAQ6jmWMHTTCQ3ATyb5990cCrfHVNkzUwGdq1shf9GRL+uR3C20sVQ7v4/+tb
aJQn0JjlSYvQTO2Q6FVyjXNHAr7wpM4t4p6I4KuMXkNXuNp6PVpERQgKViWQe974sEr/n8wacl6w
0ZeeyAlvAxPvOHeW8Sc=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
WrHRD4nLu8DRRwrUtiyMH2ZN6Vs3L2kgyFgp5P9DMlNKTdIDDQa1yTQPpciIt64OlniyoYCatBqg
Wt8N5KlawExwntwLmfujXap7EAFuw40uyJX+yki/gczIgekz/25Q1+NPVfIAzqSReCro4UUW45VQ
4oIxLBIF53PvEJm3CGD200yoSxIl9Szkkq1FCyNtIufy0im7xj9CnEg/iFEwxzn8s8Ge79lV+lhg
fO4H7eA/Qsx28fzoVv2RYnMwC/Ln7iTt2527VU0KjrPDX1WGbNCJ5ny6IM/daMbuTMvJb5fz48+S
KUNyOcNxuhu15WGxxGlN6mcj5zB0r8XxgsnOfQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 25744)
`protect data_block
id/M6fGFzXzGBIHaK7OU4GsxrPoQiEA5KNHXSgPzvYMdE5jK+Lqh2oFe/6s/7p7HrKpq279uGawq
MQncLDyuv6Jve06AqUfK0pYIvRxN0SG37fWWbBPtTBTpJyNI+ZYfQABmHRI/+isTglpi1OgVpJ8W
MRPd0ehDF7Gv8BDyM5jIV1htz+yIK5rTpbvO5AbaEdGQPOEzq3aS/44+/iM+gApm1SD2MLyLocTE
a6WU5gKlrZ60Q7AU6jRZxKU9Hh4HrFRf1//7lAgrGe109XloOS1gJP6sXPgBHITB+KZ93weCKPcD
RXh0xwkwg/QGIeRYumn3mpLa2bJWULgmOqKzh8VJah2aOr+cqBBf0VssPOZyYqLSKiwWHYar3fxO
4uCT6IQXa8iKI0RQq6DLTlk7ZLV/So+h7bXYE9aeNqlw2aCgnwNFj+qFqJxKuq8qh1JvdMNp8Esa
xJgKycfqaZHK329/OmXN8W3tgH/eEeRBZhRcgNng+mE4hvOvIpnNeoBSFmefX0VYqTUVsQjZYQ9P
mMjIKq97duuLPFuVcF+IDXkO6RnqHUorPX7nop4MN1ZSgt5iGXyt/rESNb0Yw9pmxc96SRkt+G+P
Y4y51EPudmj6kBWDVwli9Gptr0MWP7DNn49PecqWcCUVTBJP8j3TvQeZEKuF5bYR2rNbCubzdm3j
fn2ZroZwNk49CySPBPeIOnmqTxiLn7uSu7vDg+jDhsxKCOSEtdXG2tZpwhY3laHnUS32Dtn1Fo58
qFPgwYD9rExSceKlu6ylASlo8MV3IQG0SkAwhL6WV7QVNPFhCh3R9fVkBTH7zI1Wr6S0il/BtCFv
M2kPmsZ3u2llAerTXYT2MFpVgTnHTD1/amECR+LY/RRdxvGb4Av+MJA3izdJ+ZFvga5m3JlMZQ4/
CIISc9+6Z7me3r0QPYycYbTGy9GioxUN5xj0gr4UeeMYzsQIhxa+xz3v6NKlEnNLJIejvV0GHV4z
NSbXzW0VWgloX2VxKBAVcKCW0JMaD9GOvoI0pdi1Ff64oX0qJDqwaeJM0movXYWrE5rDjWTmICCg
lTkGpuL4vku1HbA7Wr80ebC8+QwjKcaGHiMPT3oEcB7adct6Ccvztxr1JKDzBK196NaqtbwwNMOd
4jn2UYXSM8okFfDCDIX3lkdl07Sh5ztPpBl1HQlhb1NRACemwjFNhJ73tpQDBYYGAa1M6BAUOKcx
R1EKLOVh2OnR8B0Ge9RGpnM2xJOSKruVPMiX8B1uWBihFmHWfPjRokYKRFimgBiMIU9O6t5Hm2O5
mHzlR9ROmsT4WushfdHJlpNyWfKAF7tzNNsilpfic57svW11lRrM5reJPRdVPBxdwtg3D3zhDXRK
ue8iWYjVietOhFmgaQbvf5NrKnU/t7ftSOtXXnuxrCwAMYn7nphMXsigs2fRrQpEkr3MhIa+GCY4
TXUmDR07zV2qVj9Wz4ls+WKc5fINKpZozc20G/FG4VkaJ2mchb5/7aOaIrJFLfD+gTFEJBCx2xkI
EVYkEanp3tivR2d0PH8FbAKsFWAJKxtSb0Dd9hPcSbwD8PKTyx+BrMwew+J2EXrCbGv2ALNIGO1w
qwT0q3CzJ1+eAOZB0e3ngY55E6WfC5LYRM6DoEeQ7IRnjFaT9yJuP4yxCcB7IywuZ9+mACbjU8jK
0XdzIJzbRWVV0RNN2u4e0k7Sr4UZxg8HTXxKotMVLR4VZave6AfMpqe49aKeMEiqnDyr2TaBxDap
/tS6ygAdRAxRYJtwbr6N4I4qfnC6C+f1puQ2pWeNwn97Y8n8Org0vI88le+v6kvavJpj7QyJPjHy
kk6CaNl+nhVCobZz1U1a7Q1FDIH1ruleWPH6dW4jvD9NXQnS78uczuijRg5mJ/WL4zxrAFFd1pZh
xllS2DSzLe73UvVpNefUSaXInP0otA1Wkq1bVKh9Ju9IM5zerh4HseudS5omildADOA8RWQrnKAi
31YlKhS7tpjdG6dun5J8r422TmRqAOgZovPt6CuRARYnfA5f1Dvj1NAO54Wkcfqsv7ICSY0kQbxV
pWT8A4iSydQl5JADZecnAApKK9ruug1HWTjjOR1IEOkpvKZ45X87KUTuRQfc4sb/R4Fnjtl8ws0Z
vYBOZ9XQsMaZKJLyvAuNOm7HlpjOslWU+mmVuwKgRFRZBGml0VOj0TnMfMmINoPeiK1/lnbodbHw
zu08n07RDczKVZ20GfMGpEmPXAH8+CDO5/9vWKWo0UE2h0XMuqNQB/DgAEIESLbISd3HE1xYhvrk
yoxpGnTNKCkIwjmAdQK5KmvJqSn1dkKtJBks0zy2TXKCdn4uOttV8Ey859uM2zlprE1FjDWKQpna
iWkuL3HHhiOSYmR4HOImZawzjIJpxqykUlb7hIG3itfgB7Evc37Oh8Tz1aaH3/dVCBDR9a9yC8lO
GrLH5uOvnFgT6mRhRC5i60xwpR4XZPsOnYCrg4G31ODmnVw05+AmokRtFHA/aTAt+v/hjmo52dUi
7CRFL1KiKQV0x9OFpU9hWGoBGtBJNYoOlzvbBewYAkTCb4RmRyDLSfkoEJqsZQNTha2PvnCRFhVT
hy+M44r2DLMwXldAkkmDTeVnSbwSkZfZ82BvuPfQqbClsiMZyPj2CVB3SnRfD+DTaJHbMJ5Wfd4c
ktVHo+lRKDG26a0q1UnoNmpoozPNGLMbzyvnZosVE+QaUX2JeHa8ZfWq9+/CpoK/d+pFcw89ATJB
4GBW8xoIzK51CE+Dv/Hfbur9FMwNy1EqnxkHqXzk7rGd5R8IG0b/6FQ7S2Hm2k97UFEVjZlT1yYR
ailuWPn/HogD+4FGt1WmnAwmDyoaFRoM/rbMefhj/NhiSSQE5LpeLiqAm9HrLTOp8Zxy9hLFpq+I
M+zVtRjwmd2x5eOqur8D5Snxyvu7VLKJVSq59hWM9XRN+K6g2crnEp3PnDpIc6pp60rACTMFG2Z2
Bz1v0+GSDfVJGfD9lsxjANep3bRch8M/kAHrihXhgj1LllnYOEXS28PeHQIdV5/eIfwYu2/GTRr+
S9Sjaedmrwt3UVcUoIzujp3zPlgZSbqJTUQezoXM/rbx1ee3E7nKuppIZNyVleL4JcxRdbVPCpga
inF8OG7r3THvN/BizeWSdrq8RLlJuX/MILhgSQDXrmMDPUXbq0vToEdXvLT5oqfsrO/UKZ1+ytyT
UprkuUb5aplQ1qJXo5RraeEd3tbV5rO+tZ8gYzIW6S/w88QXywE9kzjbS8dujFZL41LMsm7Uf8Nx
FOAFoCDUonhkI49+7jWOH4A0bTKxhZsCAQ5QUIsBnVFOFsAat9MmjhCtMKC+6kOfyHKO9uLV9eFr
xL5kHZpWFAJYu+bN/4fXJrYpRuO9Eq7FL11MuAJj8lsiHIuaW5gLNPAz/7GR0d4FQ0fHgeK2DlIU
vz641Irw3lcuy5lu8Bo7cGYfhvIu8uYNc0ZwFJDzT5LbqM7T5S2R48OcJT5c/W/bFu1mg/77k3z1
UM+dEISo/i5fm5+plEEwqbeyABeTarnzf4D56jj8B8Mtbx1jZ/au+5Aas633CXB3jvpw07QTu+aE
FSLVempc548hHVE+ZRN1gfq8za1+QsmYvx04sTkYimVBvCif9pIszahJHyDEet3WOmslP9Vxg3S1
6KnT5k5q6yGh6WNygh/UITPlBAWv4PnFbpPeFozUXXSgtE9pA4e6LORr3ajdPGYmdkMwLiUWPCLs
U6uhemynoPI1GKDJMunizb4mJneZ2pMFbK/1l9+c9ml0GftpF80tNuaAzwLfNsFnPRbeJDciYYv+
BYQMUVwaFIfiE2dnLo0OS2HseZZ2lOOe+i2ElD1IA3S3nyiHKVHdq3Mr8VmakihveUz9YyEVQ3ir
512T13/nddUuow2f0zwuVMKOAbaD8JBJQQtod4kHdWCnFiQKV2ZjemODO/jTaNV5pWZtha1D6ItS
5wyJeqkXHoR8Y68s0B1reRx7jcEQDtel4CsBu5yxN4NCrDb0SLvHhITrcANYtHKjeB7gfSzsfx0x
dXkVKpPNSVHAKbPfq4NC2jDm0frqnd+I5nqMI1/0rz8K3/vGoqv2f3yi40who6uLEg0ZLAoTAqQN
ibdG7HV6+CpixA7l7TeSfxt+O9C6SN9i0CIEEl2CpBadj27ZCiNtdYmRkw+LwTuMco29WbggPP+n
QfpEztTpVgPTO6M1pxLNKOSSs7OyEbu67a8xKY0ia2Ae/uzmRnTRcryDa8+ytsSxwiQEqLlhIV9F
RSenVH+CBIKdnQSdEqV690gwKVOUMoy7H12bKgZxwuslt7mGHRFR+0aBlSGPIwFi3dJB10oKHfGd
ee19hAu740DQ6QwtsTiyTqy7+QwxdW8AConU/ZOv06Q9GD1C4HzOydrFsbNn6QdSM90K2oeGyh6l
noEsvV1cWMXXauvsU6vV+w+8f9I4UppKuBCR8UVN1FlOK+l1E5DN/wqDJAJ1sASh37VxodlDBANd
x6pK9wn9gPWjEdrQEs5OP5vCngn4/QlHcFAmQb1gspNFVO2rgfbVL21QATbn3s5229fd/efzKxRH
aw1WrGhW+WgkEKqpaB7k4EGLXu+3nJpjBnHsxkiidlTJoHUVsM6Ki4srEvEwAzor/yXWUiKBf0ZF
2/G3LkKjmtGTY9MJrI2xWFTwr+i/ZFMvEIUBX+AAhb7q54Q2qzXw3bSnSJWAfzC7moULw5nUkoXR
rcSPLm33ThSLTcJtT3hKoEnvhaAxiPYJgb4gJK0Y0Wn8xfwd+hHLpxoCXLGLgwGA4CSvLOA0ed86
mN1ggGFJT9CkL3bwH9JsduRFsC9L/oMf2j6E/97tZKpOcw180B6VrJPO3ZvVv2/nObKi42hksSTE
T2mqxn9VBEU9SaoUSOu0wbCUb5wta+XBJsxJdAgHcRjLWCvKyudZOE3Pj2Q0BgB8S0vwP5P6zqZT
bRKTbGAoiYo99MjgJ0CE2JVbhyS9YpaEkoMUIs8JG4kYYpLRoSqJmMNpRKjnT485NpDLQG1fbvH3
W+vQOLHOb4CT/bJG2mjfI1+PVXkKxMURkicJFdwV2HsYu4IP194aRKTSoCrYQHEGT/gZ44TOGlOf
137K0su0xYaIyiwsk2+ST3uaDWWIM44xn5dTA1gi36SvQ0TyFqpL0jiDxdjQjFubHkLqmueIh8gQ
0wFGLOa7aOuXjdSolu3exWpzI/OM5ysTWTe+lz/o62OraZsvYkKbukfCoUV36bOWLzqIkqKR8YNg
m2IuImMElD2msctYEyJUYKg38cpgDCYZxUCL5+cLZK5u6Y1b09jjSiTluqG1jE5pSbrepO4o+10J
8FE2zddQGrzbUSZsTryRiHSrE5m1QnJz+WDkj8ednv6ufg71eSOFuq1/sk3U/kHGbpvsDSBW/dOI
J2HNQ5HGpQmfn2b70ig5+efLBNySeQrf2kEhiN7yg/dU5o+H7rvl1aEVdQFwfK5cJNsjrfGHvB/o
iStzwuun0YhJjNudc+amo7TkHVdtueKbuP7ULolJ7FcASXtr+mz2Gmk8zVoKTPiLz4HBRD3nhjg2
yUy87FHogHSOX0Ue3p4qZbQ8NAijGcjoyegmSJpBrZ5mxrIvI21yoLZW4f6HRNqEwADz5xHUb135
0w7zejdCh2iwWvai6LKqshmOzA85sUOMeebpMbN/4Z9SyxgUaNb22QnzXbZrzOsZFlvNmi7ue580
J5XVHfq9RIHbY3pQ1ueE5vu2kRSCMOEC4At4RY3/x8ZHme9co6FXI/mV09FNfwt76smE3VE4zA9r
ZrcaIaMZKTcuBiHGY7R1U9JDi7QmNu75uDZWl523Zw+gSdruCFELES6S2fd/lb+KBOzqKOuAvKgF
qlI6eJ8lUrGcQ0mAW9WjQWBgMxL3UgdoeJnB/kz8mJBjM6ZQyPr6JaQuzncop59gzqYAc+gbqiqN
38Cml7r3vp/rloRyAIS5lDizPtQqjAN1msK2V0qfqg1YNYRy2+jEH3fHFmZmKNJMvoWBtSD6qSm9
n6fd3kXbEWTgGMXpsAlRYZj5WA2W1Idac8irl1F5ahSGAER6q9tC1+LHpnosMSrJ+O16uyIZSFIC
LJeAFnVe15ktvMKzwVfGLs2hV6PzPALprpH3ZJLH8IuVz9DvZcLjr3TXI14Cfc/W+zVZbwt0ATeF
cV7MROSQaL6Eaa+Dr76hOIYOrop6ZkdypTjVRpUbEmS3GQI0b/CfqZomNEtkbgWwbWLLPpxOQv9W
F0gdKsQoPGnDqeS574lVMbeFyMdyP7wM2wzvUl8dhwQGItB7zQMB1t7H99UzYFDTKaROvGVJw+o4
jBgaDZyGnOw/u+J8DAwJoB7FXbjnnXXxyaPd+ysMRbxwrV2+Di4gz5YlUPjesCrBnqb/JpuzcM1H
Q6VoHB0+7RmOyawvIgmPZNs1stBrGoBGt288OMJLeUGtLf8ejBxoiEiTHvD0pSXbX6djEylHMsy+
VtqI9Xcn0urUODHYekc1QLQXiAh6r7b3tAa9pQIbHd9HiD3wQJrhPeCALnJE+Vg2Wa3geiP4+AYN
sTU3tvScsNVY0olwrbL9JPHB/Aiuey4FNOcDkGVkJmwgEBq51UZjwAEYHR8/iunXQ4OFWHgLSyQ0
AnjILlmn+2W14EaZ77kcK803NE1zad+1h5GDF5bUpuYk9B7DRXPxyCicpKR6gatU4odIaAmTNUA/
ab2GUjdmd6MsXMEXGGgYpXFQKE74pzEIZiRomHTSCb3K15gI3QAYJZfC0hHo+ThZ8kNMPAISadLy
514xKPEY48Zd3sn4wDU5IUhFb9Qbihkw4IxfAmXB9pVnJ5Fhgk9isKMsTz47J1dV5Y16XBYVRSsm
Yky6cuP0j47dqJgPVhBBZup+3KaKpf3H9KNf2vUeqPZPxfsrv6PxfUmxw2/0cIoBdPw2OYxLIYao
gN/GsUdwD+tdsUhsbnH1etv8HidlYqg/o9V5UdWZmoKhl2XrMUvnDW5uvE/EQ5rZePoceoj7akgr
2BG5r3e3Oyfo1CKiIkU1egoMjS8k+QBONFMLMOcakS9PNWzuT4JDoXji1kguGeqVL5Uq/raPFFE5
pF5sR6rSJiJxcJ1iumrTVt6M+kh0ghwji9hkcFLsttHZawlR3nlsX2ehGhF7NGzfDBZYzoz4acgN
n02r1LbmHuF2M5tvRHNm8+bdTl9H7ZWZWh4k1Zh0OXPdIbfocXxSYD+7nShku7QGmTYw5CaJeXqS
eusFPzMwozO87rJ1uxTeFg8NoeqWHHbNlJt6f9pLB9EKFa52PrwF1FGxB56ciK8WAOde9GBUJARh
/7+IrUyyEn86mfCHG1efIpn1FRS0rCJg0QxQG8jHIX2lnTfVM5cFbZvjjFyqJF3DcEq3YYTAI4mm
GnvYYBdIUyubW1vuBb5EbFFdVaSZKn2ZDJ9bTqjUfKq4ahfrv+0T4i/CXI63tb2EbYQLXeVTCU/S
Bw1Is0TjA+w0msdA8W0JR7YcOiB7ZZnj5x4+V4PfLD5L8a42adW3aPDRe5fhipbg3sScfUi0ukBL
cO5NpX2b4OGOk+RtI/HuQGGAQ5VoAFHT4kpf3qyl0pyQ1kjddz23sNcIAbntMrA0vdHaEsNdVWcC
UsymnFLqK3MrCMQXZNV3j6lmrpcjpB3yhQezxy6asGNEl29pQLn0ZL7ijgd+y60jaALvYuQYrqLM
rhWMeUX5at1OSe4/s0r+cXDvyYDqLUdUFmSxNOkJk/cEfJpdkVoSk/JbdV+4/j0z04zgGeTlS+hm
pkEyLW8f3BAnGX//1Y/g/KTyG9+ibDzAkHA75fsLpH8UkfPxdvilTmE6JOaC86AJdJM9Oc8pYQr4
FaDVNTiaXLbpfBr52CPd+fBm12Ekw82fF541MPbPRxK7PFdotReOXkG08PuIy9j1RlrDkbBPC20C
/fz3/iQZMrby3EsJ5jjbaLfho1iZLRCfOuApDJscN7pdzv0+5aPDwkHiCBAZyCFBsqKa4OZt8A3Z
ekn1ZQMwwVHDqChK6HKxNvcxY8yMW8oO1LhkrdpEuH8KYSsfc2GhGah6cu6uE3Y8PuihAPem1f8K
eNaTcK12/2TLoIj7vaw30/9W0B4iFiavhjOS0c2IPXprPBnqeKm9ftU3Sk2IrMAes0ZmqXzo/2EL
PBic6NQWHBhpse1cQVLcoydoGdbrHi9xCd+wp66lU21yUd3tzM/x9uNyGJlfpWqivDCxeRpt95vn
Z4I5a24b/2ovAT5S4D/Xwix9GbYrM+uk1NpRUEZWTxv8LxFy8rdvOvGMIOlR8JSBp17z00WS+SZ8
Bsdlroh6Ypt4I/loL/8x0RLkyhsXjQtEZ1IXBvhj1F7VDJ1DgSwZwLOtHVikHksU/2EKeANKZe3U
rlAfvoCmYzV5OXP0l4HR9n2yu8l8CafcAa3RSOUSTWBWwyvUbfn9yww4hNcoKhfvEBCVf7SvSW1I
WAI+w6Y+oT2QXmK4+GUdp7ghjqc9SrIWEmFAf6/b5BYLpQBWt8z7SKIpxrTxwVAd07CgT42+x66o
p9fsXW6W4hCKWOvC0uHQWHLunY+E1nuuxXXHoskAqw8EZHsgVY1UhYEkLb0pdhdUIZQbQFO/8444
kkrLvmSuX4MQKuN80upTujBoOGwBqajh5BYUtNaN+BzrqH5bWwTmkDeCOnR0uY2WVyy0OPHAy1y9
/mRxVr1/rjBdz07aVKxEhTxH4VH8G5D9T/ARi29sINOZSzdMvSykI6GTYtRB14kQ3dPifvyJOSif
YTxOBThV/DYQzDZlK+YcFFOYrxOmnTWHZkI7ydFvOxA9O1Q9NuWgIq+K8WGrWgwVMqiZFrZPyadM
aquDi9s/Npvy+9KIF8NvpY13EHC7Rl4EjaCEJz8csP55dytrDADChpmr2XVgcaS+zuJZ+8zaN9Vm
d+QhDZJr0eQMsOTdVSD5caOttVvzi9tHGPJrFrT10h4QglvPSbNbgZEeUZn8W+c5VlEQP1haPjAM
xlEE00mf6Lp7HOP1TY2AizIzmxTU4KLYE2MAjPDQKkX83SBZ/femb180S10e34PSfBuL4r70dZLl
tT/gXTCAV3br8UBZ5UuJHdHKvR9lMT8ubwuIZNBqvHNIWvT7lXy7MYGt9/4SszYHXICpZpJBScMV
TutyjGzYDtvP8je5DWbaVV9aO9pmjb2sIaTEqgLZMW/zf5j4G67lb4OgHMv4R+wcLIZLQULCulzK
8CcGLCRh2/H86WPPtJAyCAOdbI3LPptzNMhPDbufTtHJ53iWLihh/d9Zkr8P1mX7x/D00/Ev8v9W
8OXu3yKGxSsEOMG5wbt6rrQt8E3dZjLS51B+sik8fDV5gvOa6gMVi5VkHPSXd39bmWtlLgfQciux
25epZ2cvaM45YDgw8xSSFTuBbwpVtYaDZEWD8dB/A48fbVfJ06T3yoKBL6zrxKBtZkuUW8NCVA/h
VVQQN+VMqbLV0nX2CnA1neptA47odepwwHZ67HYEzEvlvayJkM+szNiKnitBEGYiYSBvsbzCo6hS
fAawjkcwE0IVkt7MCsc8xu1orbQhs9kPS6aCf1nAP1KAKFLYwfl3UfkwuNcNTECEzL4Cn/2UK+gL
RrJl3DzAK7r+SgwoFGw70eIWSf+pWa135jcwh4SZ7T3bV0+sobHPEkRrKBcFKmwEiJoVLP3doH6L
wQfkYcZbHv1vEsI52Ivz8D6yDB5azftAC0TRi+CFjfzFgYaLilfw/9XYo8HjE52evf89685iJFyx
MvNoK6BVbSpS7mPqj/pz4DjvWzI1rhgpNdDEb4O585Z2Kjb0axZb/T4HynfByr85kRD+6eQM8SwA
SiMnOP3rESl7rdEIzRj7RUjK6kzzDbnCdNiWbPPim/dcT6gCS6bdur7ZdGqUYZOUfrjMsz5r6Ta8
a96P7FLKTsulUdKB2ZHR8/x6KnZZ/LsM5eK+D2EwrVWS6Z89VohxbIEFJGrtz3FNv0hqcX+GJoF6
KQIfpkOU1CnRgWobtX5jm0/n35PJIu0e4wI+WFSj0TYIiGKOBteODJTzTpkZs00xC/LOWRTB8uKF
SgLRFb11ksdq2a10B9hdCiXH4Q4a22GL7SGTRdLASx+2ClYogaDSGjKnnNILQ0J/qUe3wHex8Fv7
94WBAV1wRYTIvV+kS+FuwN97XiwT64nKzcx7XP/58zHJSmMpYQQH6EBTyzGTEAa2/N0PM61Yj6RJ
peRkEITaVt1jAKPf838toV5qGttTstrBMtNeJc8wsfYDzrcOIz3yraHGc8CE0xPBElFOHMuZ8c40
JfReEGMPgaofbp5SFzNAKv2N5zXjoGr0ePYPak5xEFVlL+mvFKfEJgwxdnpB09p0azm4cp+ajZ9d
ZiyPuwTVex+TqaJ9xKI9n0acPA0/siNsEBHfg6gJieE0FtBSRyAHrAYwPUOaU8UZfF+fmTwOFHs/
lJDhc1Kv264VbYt039Hc4KtTPte/OZBkWPHGTqYa7Wph7ogxNxVEO7yWKarfhQb3eCVSbV+kTovN
RSMurwjlY1YCFySK2kr7vAQAkDI6WgEMa7Ab40nyQcmJRFoKCpEfiv7CxJ8nQ5LhbinvNi3pfqff
BwxVgQOVd5sa38w975Q2znOUc0t/Pwk/7pJ2EgsAQM3SJkjcgRRZsE5Q1SLgQ6+O0ROsVuiqNwWC
TiEZ6+Hya3hnKN6twWL/YoaqOl/ovE4rB70snkcenFOHEl2En3XXgqJjJtUUbFf8hkXtdNfP2UAz
nK2sfefyysKcFLTirEy4uXcoOuFe/0LZNUAaBwy9kxNyV6dWkKcL220eBygZOFnGpu1mOYI3Y25J
9dgkI27R0E8HSF9YHvMJcmtx/W/5wBuMlwW9bZ6ZMd496k/YhpVcaHS29E4NL/MdLo34XdTH4o+g
sH43a2NslN/Vh9DWCIZFTOJaFMzmcC6QLHTtf2JPWRSWi276lGz9ne96wy4Va02USn5vqfinXQEh
4DWVvklAlHyh7O8vV0egHWzm3WWr/50b2PuadPoCM5KZWxo3lLdqIMVfhndnyOb6XTjxY02AJDeP
nPNdDVgUvw+Ox9862mP9CJI4MCMim6E4uCJPC8LviPLoPwuNM4o2vd2GNxTnfFqiQ4s1Gn0U2a+V
EryCjUUMuNaiX7A+uamufE0Z9R+5ZjwVRKeprzsYquSPdlJCerUjYGAbnVDAiyjfKKZd0VykEDpF
J+djf5gQLfrMyznYfPmB4BoHS0honoYBHk6cXwjnMe4qGKan1kBXKP3lpIoOeTaIkrJcJZGOGnw6
/9hIGjX9STQZAw2IYJIawlVPnae0+yQomeuVQBTGXGJb8yzbupsI37btDW5m/Y7YDwy8s2quyyDo
K7VjeqFNe+oEXuFmrMJa4rTNcc4q1mLnDLDXjvurkEFrpN4JBvpF1NZoOgwhtFtYj9BtHTmRrExK
OilFOfcOh8lJ42KMED2srpfn/jHk3dAQmdCOoKmzkjUkcM8z2xxPeYzQcMRKWuQFv8rNHx7R90ks
iJM1o5QoaLlNKOXCsH2QAMYt2HeG82H8ERr4p4WQWu8YFXS7gUxT2IinHe9zJPn08829Dh38MBxk
hNxolfrLjoKjWakiyZ5fImjHEmj2qxVS3UgwkmNHy4nZ7WiPY9oxlXSce5RiBBjoCvuH3caghyRn
lU/psADH7yf+QgZEDxJiz+/zQSAg0P0edmLwLKh+3160tqJ9QaHze2b1navV2WCMoEJr4g6jzA5F
cmAp1e6jBfBQQm5bF3cSjw2vmfzEdxXUfUBmYBuMKUmgf1NAa04VZg1IQDsYLbNKyhsbnl2pvNG4
R4wMckEggQZBgmf6WyrT0fiLtcLoC5nqTB6mN/xBJ9OmGM2xJkwA3CfwGj4952ixE5q/h8Oou3xa
783bhJbhBMYPQA34NzBOL8SilpbAvHrMCykxRHJvv2k/XHVJ25jPi3ozEgMGONIpKpIcPO+0TVjj
BL7fawE42pEQRqIoJk53Lu90uo+dDLDkcdt4UvcmygbCVryDaa6BbDXcUlxLrIdEFLcRKdx85Y/3
WfCzKMGL4ncmLWiI1sAbyl1DBZXjA2mJWO3vBb7ZEC9FidrhZQ0AyIugQsDCnFJ8S0KOrUopZ1Dk
zcKYiBaAOb9YmHCWI3K3x3A9ognjsiUcDLgnsZ3uny8NFmXVNfSKw0e1n4z+1rkx5hSK9HkyvJ2r
ipeB/dHb0AoWchu35Sl3NC0AzTgY2ycjRTLucSEzXhV2XsSD8dLp28m1Huamo0x/oQNnO7TzSvUG
DydZgUAQVzell/4hpQzNxZ/rXIkVHawT4f+6CjLm1xHpPuaSW7BKgBD2k1j2rjtjCetKm7Fwkn5N
RA/BbCK8xHzrIylzhKeWHuv7sdsqRN8FMAMS2/L7B2UdTeV2mqL7H4Lq3PJwaI3SZF/6g231dfZE
a1/zDUIkOlAZozvFQToEn36+CuujwHqrjowFjFzeZhAv3ya6MxXC/61jCTUYo0bbz3qi1ufIyVlP
jEgAP4iJA+XHn2HkQLcQ/I9taPTA13q6/7tzmkLPxRuLSn9NeDe386+W6AKudlyoisn4TTCBq84X
Go8pYuU1LVANvDrGbBOfysimBzFv1qbwqxKuMdCsZsgj0v0fomiEv2OpKp6VvpV1xeHuNn80H7iY
RGwgIU1AYDp8YJ4BfbbPrsXhZtwORuikoY7by+FSzgj4WFyb7g/QdAPCjoQmFnMsw0Hhx/eSpRhi
AQnUKIvKCWo57E+Cuov3heQ1s8I2dojr3G5W+DDyhQJF3BUfySITzz8a7eMPdqt+ONrjhiMot8HS
FTEIG5v/hz/gNZ0RI2EbTTINvHtPigoZ0dNCrKYigfUKSGy4KAIM6EUsGw1kJWmU9Q20EXENxifV
Jty7VwxNWI2TUyjYnuw/DB1uE3oJW4WEwNLGvhI1IxwJHLD08qhoxSJvhumTmfY0T8Di0Vb2qNma
2cx2MVRDL/3uTCa0fdGH4kQnuFV4vmwL7t5oKE6NKiqH9Of7Q7uXEXgt5mJ8ExiEA0Kt+zMyd0BA
igMUQ7BpExbbyaQq8USRPzRltE+Hv8u03fVClKM9LTGIvnfGP9bN+M8ipZh7L21sQ7SVcy1HeFSq
acZmi4N9K9jYzta2hfQXhksWGw2kD2D9DOqY7JE4cok3m/+pPZ4/qRu7xVLX4uMYFac2kt4RYZm5
QUHb+q9TKvb3EaFiSTT3+aM1n14laBuWSgUWmz0ylNoJOPNrjW+9J/eNZl0LvxL73gvXbHvyPiu5
CvcPhhN45G4Ag2r7UkHqRqjpcxli6sgVwrc5DgjT3r5Iw5XafSVh0tNeN3WGhvnnqH6Ixt/7oSpt
W5rWyONGBSMo7If6bM+tiDh0XWYdma0bRFQT9aSikO9kjSVVriTX+CKSTx6Du4tMpASNcZqdVJ9u
ZbkcHwXqrtvN7k4zariBvUClZj24yrDsCBTu3wpQCMVVhTOq39M7gRDJ6rNRQwLZeoO4qbO6PZZm
KEUruubQ6E6MDE02ZnV4C6Rpoaae9j0OhpkBIhnEoDo8hA2O9p7Vtzfrf9S2L/V0dGD0WMWi/vQ7
AelVdvX1dOfu5uXsZsRMf+DxoV2J4q4FQecp8l+l8zZ2YOJvOZ8KXvGQJGg6BoXO8/PZn9FtT8G3
qNo2qdeuHN3Yz672km54Klsr7AE8li0AAoYYxR7HV6BlplyAWTw29ksfOWF5YUEJmBbZa1LmmWlb
TfxdqYOYE9I0VVzGmqb3nKYfOVwKiIodvkEqbL0KuVB3OFjHEqoSHwj0mP300NKhZv2lw+a4mtWs
5OPRYsjdtvxCU94uH6LkghxcTG82cAIApaaekDTLoLVXUO8D1b0CY0tojnFjmc4Z/NtQ+4P/IHD3
7einaWYAQSJlJi+Gtdtnsneus4SJWHy2FOCYh01mV9c4ifGrhNR7neHnsKBDaNuYmUJvuWku/11T
IE/To2+lGxVcPsBLeCK2djHbESonFhhTp8gwd4Byzd8OrqfjDP0tH14oe+o0XzzC2EepOCvp5rXA
zHbXJZThXkpKYPWE0eNuT9FUf2FYqPA3nD82zLQusAZqDeTAQDqNCf73WVt4s2NnvErc2AH0VgCA
L+ONTOJtaNeoQ6Z1oxFBjobSQ38/vDqE37/CgMQs8Dy+/bZIO5HKBiLqlabuEDIqDwp7l5VWGUVl
MU2eo38tAH4zda9g3u8vtBaDN5aitvPJiTwV3oGaQz6SVIp309HEtLAOOcsdzD5clDkvlB8RZZjn
UG56XQWsgYe5B032HyjY+W+HqMt0Vk75Vr7n6BgCgHztRuwCLUJwFYzXvmPHL7AtwpD3eYaoJRI/
AocUbn1C8Ml6o+r9ZqMx3RrS6Hki57UawDCguDGZOuAUYcTD9nXiCXLd35eZGtFarnMOVKaku20j
3ll6P+XtHiGQYXvsqgPiqqwsdJi9Su637hGvb8l95GHpzkYuiDTCDAU+9aAqjPaFamOBHkuvgag0
+H+LQDc8lITOpRpOuO5Tjltx1WftJQxw6ga2Fd1o6mF8ElYBB7lfmkp+I4qZg50RI9/8rs8OduDL
odaciWNZxxNo29ojxxGOnTE86niHl5OuZuS3GpzSIQrSDD/ylGfgVNGS2+KCs60dKPT+H+fxf0Vl
2eH1wkrWT4XEmEajAbXIZkgUXpM9ZvEL5qN0byuL4N8IKLQaCLOBjXgYt5++4AR140NF+17rX4nv
Mh4btLJpoy4xyMoMjxZUAfkycBV9/3N3oYU/Hanjp+EmzPtX1fkuNQpNySw5u3gykM9SR0BYliNp
AkM4av8OOT38YbrUOQBrennEV5EN14vy1xJb/Blt+eVoD/HsPIUkbfyXr/98MOQ4gyMBJTSkuSO4
7eUcPIwfw0n6qZdEZLVixblj7z/AvGqHscdF1k9+pCUjcAgvlKUgjtYRLtfcserb3jKVJa6gWkYS
WSIiixj6A4lDtTmgXbzv01gIgf5trOzC0PKx/20EOiM+115SDHJOf4ijEPE0vJU3tY/h92Hl+zuf
Ozr0c6+JiuFfyEFLpZnjsLoOzrqrtkJQDSeqlGbUXxlkoAbiLrM9fmbFdGK9gQn1Xva1puKc11Sx
kjS+b6kP88oDjArmRVD4OE2vByfa0s7lq9pLZ+BON+YMqJUITTn/0B2pkQLdiEOFH6DYqAtIZmCT
1HTvDmb63qDVCXfJ8DCyFNIzlgI1OLQLNtEDx/wecJPuhgvG3YQxKW26ozQ7XpNYiVPcmh+hHQtU
rqAKi/fh1Z0HxD9vKnYMfbwX++vbH4602yhXUF+If30TWvhT20t1DE8/n6q/AcQhNqOnK5g+ObYq
W/y0w8Uu8KupWhzOLeXeTCyEP6hcKVuR1l0E4nWy0sVIirnUnwouTxQdmD+NjjxNBKv/sdcYkWQP
rFbqvDBL/p3XwooszoB+dF2NTuSU+cQE0pXuj73c6RTcF2Z6pmVBGsp3esVmu7KTqA910Laf/bp7
2QqHAhmLQpyRYeSrOWzWfVAhQ/tJA1kwJF+NfJa9HEmbVGFLoudDZNHEpSFC781+jT0FAEh3KfAa
Dl+Tdko00B7QGVixH2nUrrxRz/NZrgV+r8uIaM5Kq0jQCIYHmNkmUXYAT5R3G2ZBUONvvjJuOCxR
StWAjhVMKVwaGokJ7cZvaPSGu5iQ3R+T8aoH/Mm9obBuQG0z8EtIJP246/YdeEqy2p9s4Kc7fSbL
OymAo/iS77tjA5j2VBQfI82MXvCxEzlszQQJgcOUpHHhNIB3IatPlVv3sfumkiMmzMjBgBsSqb0U
B3H506ojc7E3y6xo1P5eWv8uXrgJXRoLQ8clTGXLjVRHuSvjxHTLRDRTcMY8kj33Fa9XZMVIMpaI
3w0c5Rid+FAeYqrKW2Mq/X7C3sBbySsVVsaqif8JM9Hk8GOWXx4dFHI5jkgBW0mc2E0Onr/EB1rW
3IzOs/4/luMco8oaRfN6l20zmAKt1vBAPCwufLIOUr0fjN8NIRqxzyRlvZ92X0qlhr0rDHLSdR6A
2Kvc2+Jpj+N4RU3rylRj91II+W10vPqHH5O9sVZFhKbhffd/S3MF7RgnnZy5mTtlrbOBQpCLWgd1
eQnilVxsvLybW8FmV780ltiVrznO9iIVhTG271W9w6lsE3u2YuPbvwzVIYiSUg7ooKy8h5bErMBc
V0KNhuVB2ED1l4MNuKmofPXMFkHg2HR3asjUrx9pOUJfMyVVmjHGiicOFgu5ZQ5zObtji+gh1tEr
uePd8ac49pH2p7WuDiV9gJoLxJDhOkFRmT0w5+R2eq4K7fytRn/QDv5cdkId3yE+QrzXkDf7D5B5
mNSGKBjm2YhvgJ2RIMynpa0Juy+sW+1iqRwQnb3OvRQLHeXyPYocYosuoxixxl3RvmzD2Yt/Cfdg
vplXaeFn33qSx2t2xlIeLUvEeSUpzeVjB66U+NcwEIYLIlWHwTn8ggnvU1T0DAmUc72jsQBgqJIN
gYaCtDYbZO6hXtQwNCT9SvF6tt7FktaKmUvqmy//ma7wLaibU8/w42qVMy0T8SwNXYZYn8ROO2Vw
UCw/kRa8vACsTg4SzXqw61iEwjxyqxQVvJCNWBGS0DlbzfbaU5OiefM65OxJXJ62U8L3pajocPDd
auV7ajo2ynwMrh4heMuhSjGAtbRSbCB13gLudEy4b1wMZZ+kYG9gdu6dLWnER/Djl+58O6GamqB3
cHr6vZhK6YLUG9YVsjSrXSQj6W6X3p9fdsxBesPsEjDsxtCLILGojEcJhCs0BAQs8cDYjCFUBzUC
O7NdXyOzOGVLSuUT6jblGxM0C+QXKI8vJ6WSyKLsGaHANl8+QwqHhpfxIeu+7RT0srtzrI4XwPC3
mXIbjHCpJo5R9bWP9x9LiU8D33Q/QDfxAV6VpFtO7InvfA4F10vtllRNmpZOZ7B/CXTfnR0Py8kP
UoECrmtF7RMMZ/kg/3e0rnUIcWzyCrCdsGmP/d63yPCidR2bPtZtmVI1SzxNOAK+GxFamljRrD0j
LlUrV8FPVCOsTEnLkrc8To9bnQZ9ajTs6QLIawYkYAD0IWHou0FHWYiB2x6HmpSzRdq6b17tA82s
ogIJaemJGM/4k4a0Tq1mwFEkh5jzq/eQhRXCB2mXyd/CkK4P34xP5Y4kd6bvMH2T4QQWhkHMmCsW
/Umu3YwJEP5VCKCGqVWtYcosl9ab6dXT983MresO/992az5CjcV0Dwy7cIJOk5sChl8tH94XuvOP
VwvDWZQfpJuxES+uhSqDSRuCFnwuelDE2LGbIJYYTs0sfeMR4Ypo7ksdGGxCULpOjctWRrf4Ak1L
WeC+yKSsGgCstEdq0sQHW0S2LNapPUpVxmnYNMGL0hsmqG4TN7uWp95i7/HDC3g65gB6qYjJEM7B
TpxS3/UhixRmElcueZk0JvXEzWgxsR8fYvMi2dd5rVOJ50yU8yuhT+IiJTkOrmyk4NFj8+FmUDBL
k3kAbPqo750gyCMiqzVs7HKroA2JUNoZ5CuskesB3ag2ZlLXEGIL3znYytaSOu/o5U2l4N3vN4Ab
KSnUFY832gy1gLaTibTh/pIi2Ccxv4EIeqZozaBN0qYQCdl31LLffX8P2so4jVdbSA9JwxTlvRDd
I6ppwSbME8TLB4iGdUfZ1XbTCVCIpeAhaEaU+ASQdApVbPUNt2Rym9PYIp0LpN/CC82UP+nFXl4a
OGRKTL5uYSLWS2ojiVuR+UUUsk/TinepWl78q/bmlfCIz0cVbL6XWsaoEKKCy23t1wIPtt+kDY7p
+smB0BCvd7Mnvo0m2LQpuMuNN2nu6/l/WO7EBGzouVHQnElmio6lXV2DgODeDBPc7wrCEms5EgWg
8eaODgBEWvK5WEch0M3I7y+ToEFju6fFuw8bABG2ZdTbrzNQyvTnyoYPG7Omb7cm4c619X5AFBT9
Y/OJ5dF+U4DJSaVUJPmmcufVHN1beaNDZktBSM3S3kbpP+DqbMcU+3qzPD8kf9LB5cV0/LHsb8ZG
+jovttq8o8pIV7bcjT0Atea8SWU+0vGL2r59vArnkWCOgqBlLEr0xjx8wrQNPAdYjJrdVwIKzaUa
VauFsU2KaNNus9VWghMQ3gww1jhzYetvFEzjvAlKjNxpXYj8zfHTgGYoXcvrTjIBaBUM6semX7KR
FSO/KfCGKl9pUFImAlKFWP1kPsjeXt3dTxMYzfYGeBoBZgskRJQDYHxEtImWaYGjDVklYmS5Z8/2
HVoHoMYJVOznGBgxTa5e2T5K9vIEnPmpYGs1yFkZ38lgOKqCFTPy3Vuh3WWHKyP5U5ugbma6wdJw
hENnMhKCkfPI3yrGj+4Ubmy70k1Hvv2aE2eyX2MB3C0M4vBgXPIgNzC8N9lNCpWumohscRIAiMX+
m0xVPvnQZn97YTbqqkT8Y2J9ucqNHsNAks49G6A1kDA0YHWqtsTO2gXoSg68db9DU72w7d7YG/F7
lpUsV2IEKh6sDzmwt/s4j74HI6Syrl9aBWS2kWd11U3mVZJdBTTN5ufoljtVR0Rmx0rDaRVKzVw6
buPgHZIPppTuGxS8M7lZROSdNZduklyuzYem/4/Vc6Xd9j0nSJ8e2tKOopQGLLnGfAhFyb4D9L8w
CBjHoYCpT/bJKWF1ovaLrMhpjW6t5N7PdeeNWjpRPvaJFAVzjc6ueS4WGpyJmn/Db573aUZQDrLg
DGmnZVwIb33Udlh+sOl5qs5CdN2i2I9OcFErZG4+RIS0jXEbsteI+g8lXIKnFEbYLzWkrBk/u16u
0YLgZ/ZGndj/qYBDv0NTDm4f5Dyl89wGJAFsU/1Tgwi2tk6Qi5EWd6dKELkdToTqEZxigNIZSpVM
m4n1/Il2BBmQkGCMLdCtgyULNdE9IRRNz4ZY1VV877ihjvbMgds7+vXGbhraq3S74e4IzsR7RBaV
ovO430GRr8VDpivUKVh1aPmF3vW4Z98kGjFUjBvsrhLtvvIv+YUCJQkgcySTnzPTcDKYiIXea8fN
BPYzKapmtR/p6CzBkA++YKzdi2BaTU5xcwkdNQMsVL+142WeDnTS1PVfAG4Hjawxl/vNEqmWGGAN
hO1CIQ/Uy/uxJDfMZrlvrvU6vk/Co6NFcItrxV9ZCSoC6vBJJ7+9+4ZwCkLVClT9JMN0Kem6ApXT
RMM3y+A9NqPkeUhdGs7nz9XuhUHX6SIxJZVAPQzzqy7558lIq0dCmATXBiiAbCPxa2oeZu7j7EgR
9VqsE2zS3XrQhEiAiL+njIRQiMNT3SU80Pgxv1PPHh5MAzB3ueNWmBpZrJFEqQxILQ0pORk6DQlO
WihzKYF8Up3pvkLZz1cSiXFJipx5mpeg5CVX6Jxt+cG09B3a01PmjFqLmciwZieUjwjGInT/AG8Y
fvzIKpLtlGcDYdcTn9ST63OGrLXAgobsFo9mE/m0QVKvJqpxSZcFOJ1+57cgnGmKdYyK7WReQUdv
FjGvHZ6u4yqtNZk2GFlxkHxWLBvKhKVWcCCEtQA4lxCK/rgasqxtoYwKOfzSbfFNg5lOZNffFcDM
sVaMP3pUX2LHWfHJm5yr8UdQ+sxHdo9T4Ac8eL1Bv/p8XZR0oesriMF4tmxoHiDQJdLBb2a4C5fv
hl1RVRlM5+VSZjTe8AI6U8AiODUb7yLTzS+MRxHtx6SkOVWuamDPe/q6ZKtruoqv8z8R+gUDyccj
kH5qRhidpPsILm/Jl5WFA8qMzbpsf04hdCKzU3CvKau5yX4OwAa7HUwitQTsZhrE/jRaKY4hP2K1
6iEeLbsCGQPSiqsQhQs9XZxTOTIEFnouoE42LFWP30RRvSYSJP8zaAYV+ui+nDNt3nioZT7gYn0y
vUlD5m4pszhMhd3b2tdKUoBc95befc0gn6k4Cofe9UI6uxSULgywLsGHIdIgSmc/gQGaDc1hxNxB
guaMD89hJC6+J8vebxWA4E1fxbk2UiAl/24lt2WY0xwvucRvZTPwKLTfBtnMLDu6t8F72AJkaFVg
O7cTzRLcpb9pxlwSs1J7olEzEh9LbEyAFwvtWKCZhFHWi1gW0LOlJEbvL8mtxFqrsNOPugAIIbtk
FdQOVXCOjP/ZbJ0I9HCz/bUvM5Lo6kA32+4LNXyqjNancU5qA4XVnhw3MGMZT1PLqjGCEWEr4l1Y
xh4T189yYK0JoN02zcMiy7M19pb2dZPgrJ7lYHoyp1qHot5wT0T8wvXKP8mMbx7fErdeKebc88ca
ZFDHatjHMl4rqAzU/+T+beNtz1Arqub7auk6gKZlzLHrLDsq2CSRxcIT/g5fFRLusuSndSHwvIEQ
PWOsnH2DJeVmIfMBuxvDFG5jhw0gW8qRIyAE+aYl6F/YQcImz91qXCUJo0LQaoc+cp6fVrxw2R69
rcjul87StJEat/pv772uXv6uD3DhJI++AqX3REaCP71pdKOXfI+ygem+3hiNq4V+zLYbQUZ262Zf
ZXFBx3aqvkZHr53v8vAwXMGo94LKF5qsR8okQpkTjd7jwYx/qoI9/hUDogpgBLbhlMh8lfzUszOf
b9LlUZE6qdfjeZuaY9gAJ2ubz3OnnIby76M8t20zqnjDZR5tOvW5xPoSf6TAJ9SpSGQD+CImJd3z
kbvMqblOyooDbMtTOCXja2yfarG7CUg+fEEXY8vOFLrNSssbAaMsQKgGDIk6HydPZSekI6nGfp+3
Erg2y0v//FcL19N/er4TyIbP6TH0OFVvGdkPDl4ebjOuiXHy5d9fMmoc/9CjFNkwga7qYlXJShat
usdnPqwGMuOODjHrorKMrJigzaTM+OR0O3lnVuuy7YtxcIT56SzdAh+6Mv2aZ/W/lHb9SDH3/cRf
aaVjUxNNjDhwWtJQcTUD+1c/lY7eWfnWwbIXA6xUy3A49QOM9djlbQPbe/sL62xRjctas0CXjVRg
yeH6LBHtEhwn9Dq4z1gSa6IsaGNUWYt9PcXc3KDBpetGHc8vT/6S0hLpXpSXWtfaWK2MNsAhMUib
p4I3QQvukqPRs585rmlPuqlCFnEy99UUnXt4bpg5DLwJ4HacU2J8Er1lwwGJZnk76K6rpIYCHR1S
EyyazPLGayAPC6gNNNaYs60io4aT8r3jhOjQTbh4cbFVAiIp8NchFSr7snJ3H4USPeVgCtTISVIg
RXiYpYS6vQr9r3EwehZkEtNMkskpyK5/7HYw1sWx8wdDfvmfN8mcGrGwy3t/6VVQch9o+mcTdJjq
t9/nL5jKFyQihm5iPy6h/GTqivunNPmA3G4TyuDv0QfWEDh7L+wu+X9zzQ5Orb1JmJyLuGKkkS2W
Whu9iykR+tJNifSboAgQuRq6F087t8URpI13aKwLMFZWKx8S4lbxDIs2xENRI2WqlilwKAMWqJ1k
Zjn9A6gDfsWYceX0jgPwSbe8LJJDC9dwb25L+BqE+VsNmOEKYoybRwx83xIRbQFUYNREFEjnZhJv
w4hNeGXY4aFzXBccJalz7QIeDLlToHMTzk/isROoj16ID2Kl+6yTsMXPbFSuPpb7qdm0zM/rdlFy
3z1T9MWZwOlgWACIkU9Wn54seLQWllLkuEUlA8K2RYIQ7mk8LyKhXZuq0rNXkCftSewcHXvJQRRW
RRBSq5buGg93YNEIAHY+IZvtBZtSdrg/VkLqHp6TxRHt5WOV1PJxyUKQflasbOCFvWHPJzwx+kqF
l04A9fwfqbrHhH+UEsrZXSvTlgWdgZKo8VO2OQFwG8Evd9PcABSCn2IfHqWZURFaaEo2g8Ztp5xy
9rMfugLnOq+m3fVvN4chlnJPpIwXrY/JDwzLH4FPfkczgy6h8nKMscGNS6VFYJfG9eJsl2h9BMEK
/JkZaDjFF/p7n1TklIlyB72lFyJWk1S2Siw0ECFJkIVcE+mgb7nr51yI+Je9HECzYs24yzzNPz0D
ixd6IXREy1kGWGR1Lx680xqzSPxaPPN/nqdK75aYjkndlqeFeYBu6H5mU4pf2oQcE312FZJca3OG
gsK4lApcpuaFYvkOUg8RWa8YFyBL0nl1fTXE9LDpvnfOzCqTuT1Rg/GliMozfUaMtwVbLFF7+p3Z
83G9K3kosQAga6Vn/sNIYjpRKs211kfac/MtNSfv5kIXc+/gPvY7wd8CWBh/+JzwdD3BRLJsMVd2
orUEsghf+538f+E31+/zns8bSlLkNpPIRhvA0nzssKX4XWm/MSY5ryYOqQlHCzCkQxRQVQ1kJgGD
Ijajr/tNQkINhvVcsXuvt6+XSoWZc/qPEjY1df3r+dybPyw++Hgz6hO3A8KM0tmPGJNH+3aY9t2s
3TS13NWqAS4Yy4egfXhDvcKtC+8W7fWr7n6W+J4/mL4pckfrFgdzHaHlkhBbWw15Ma7jb42050gQ
Gvqwho4rVH8vbhfTcHAsgYrtKTF17RM9wIKuTCAzWFfM/4RfvrjoNEU7WwYUW6cME4Pn4mOixy5T
q8Oi5ag+zEcO17IdBCFdzo/UO68tKyJ7mfppS4ZEdTh0OwuYHnu1MEv8wiZ9E8bm8IyiS4w4wqLr
jL5Qy3Jak41jVFzo3iUYNTVLMITJgKCqPqblP4sT9oQQ0D5zOzzi66wAfJSGjgJnZrv5j1vmm34P
0QzfedDjiamjRz+7dohAPXfUnAyTHxtzeIikux2tN7Q6QDpOg6k/tRDzVBk+W3PYxEygK7j3KVBR
wvhuW6qB5khy1wz5aBXNO+sgNcGyTOOgF5D20vmLYsUrLSLQ9wVeqzU/H7mLgRyNVhWBrNcpvpPV
NikvCw3BmwkpDbxwPZ8KZq4zu+A1BmZoxK4HPpmkPoUFg672+XC8X4o0ejulSB5gBHnaKtk6Fiwh
T0zV8gkJFbbrKJ/7l4+5xuaTSpCBymRKA+vSZG6qGp/vFzaTRd93IqL+YANvd1Y3HCZLtwNZ4J9N
8RVwanhc5F2lzsvpEFSLblb7JGHd2j0eMEa6MK8PHFhLmkxIeA/MCyP8dxQS80+4Y6NBrpiUDID3
xct48PhmIw3MNewwRCn8Dq0EbeU8sro/aaSFFxVtDx+pqID0q7NucQbytPBlK9kr3s0UTgtMuL0/
AxGpJF4QhR99e3mMJSye914m55kj0HTiBqwwqNDuGZuyFLBoXBnKKhOiW4hq9Nhc/VtNo/MVT44z
nzwTXQs6LBtYrwvq8iEpHQbNlvThtSQY9ciu5TH1v+c7v1gCdSbLzT4EKfi3opGuOHviBK7FGXsl
UNDajrJTuv6xQSvoHVmI+/B9iqFOHeNJ2h4TQkj9jP/8zEYVjbrp6CNngjlzD9J9fqXh9qNT+tOm
V0kawcpfSexg4gIt82FfeF8Uvj2cPuBcOA/C+sb4CbJ7Tcmt4AaMjGPR/cHq+Y+A7tMhXZyq4XGk
uSrpHzNJFg9mm6zBJCtElqFuNA3YOWza+AL0J9f/J9UhSSHDk2a6u8/woxYK36/Ipyv/ZBvE/IAY
mJNeqYw8QUt23wa56PXPp/z1+beBju7JsStEwPVvL2pt6Hp4m74SYM6CpETar90TD79fFKZ61Lth
4/FXkH0xHv6L3tj1V4W6/GEW86gMVxtyG7/Xvf3xM6Tlo1Gd3F5yJ/hBqjh2heXqYVncnoJPLrOp
DonMkmUZk7A6eFz2fTmpOI1c6LWLB49Cn+CZRylRt44TLcYTOnsJMJTlskt8RijlRD4Oi8uofcgU
iQ4FXt32wlAYa3suzmDIEJCdmuCg6dpzd8wUwl+rmdltfGdmrmhZrKuDjeMhXl1ohEGgbn3cUsCd
H02mA18Vgk+Ke7Iq/sTbK1cr+jSbRUJTDwBYZcESNo3PHczIMKxYb2a+p6d8nVJqWR9/jk6o7lc0
xAGL2SVwqsB2qDKmIYtkk9Y2NjTF38r8JiKvHSzR8bhHaLdl65sbM8sARcGyhJl/PQHSDe3TB6m2
DvG7B3YB7v5MxBdJqZcQ5FVEeQtea/x7Gzea7USKLuyBq+1MhgTZeuNwQTO6TELhPkc01DmZIoAP
Gl5YLyd1ZW8+ms/XxT4QP9NSKeP2kyk+Cxk07uOtxkyJnMDv0xamWU2QlRRE9UDgqRQTSamF7JgI
jZvVA/CAzey2thw4X6hq11FZb1c3sTXefD/qjM5ZCEdeEF1qUSYCuHVhhUhQrRZMXKkP8Db6vtRe
Xp5Cq0Nngm5S+22pYxu/0SX1LKlVHcrc8DtIcB6g68503CGU1qhyn46VcKIj8o0XuGEVtCv8rmVc
DRE8TIHV+OuM9Isy5DyrI2BoUcLCm4Zx05H2bbc4het3obmxTSEHTzr/hP3R6XFQ3H4gajiP7XjV
Vac3KqYttI9o5BAd4zgXo+CB6OnEhzpViie0Fg1E6GuN+43c1vOyzojGj5/S2fxGdaQBUDtRZoww
TyF5y+bGrPEbhR9JjkbuV9TEal9Ck2XVmz1dxDqO6p0tftJDg4HAxmW1uiIfwGAdIdzGnwvObeA3
nYcVmWOxrdguPoqFrPFh3TFesvRY4B9jxB6nfFHGI9qdwoM5I3nK8uItJM0Tq2GXP6dENJn28VqG
ovRTQuwnRme/XeJZdCekpop741REFtVKGaaOwWkzE2KxB4wWWfihT/JEny77FbaLnYeyrBrfVbMm
4nUAsUxeDzOw/kRqdBMoyN9kev+NFBN8/t3wX2TqwOC+0AcbzB2gu0677R7a0nr+8RQNL8kioiSL
PlhtXwDgaWPJXAm1eB2V8BeiHIA6OZReXmJy3lh4yxbCPkVOgXqFUg4dQqBkKyn44GeK0mUHvwZU
60CCDqHzr1KXFeSUaeVDtnSJg/ttkki93uHzRmXFG1AsdrxrUyw/eef0s9sQu3D89M4e3UMafSWB
r5PVH4xRXBlJ+g7belpGhvMCk1yo/WZPw3Hzo/VFIdMhL3NjBQGGLbB4qBbDVdzA+ayO6BxwpbIG
GNxvnravcndchW1LXTnwzbi7ibQDDWs3Rcya8/ipUZ8VyXPDTi01XjtgKqALh3lI/wotsyzy1oRM
HaNsv2ENMDTE864Qs+6V2+0wki8Riql8lciuAlGzew5muE8rKhwx4UAw1Vibh63WzEr/vINJFwm5
nHQpEbWCS2aRapkR0uVNqZjKhwRsv0jWXgeVuZkAwfg2Sn+K/swUgqH/Muuk5VY0emGz0IXsSHiu
IAjssWyaLsRzlVLTxkNJ9U1xFFReYezOsMJfot6J3WLOgt3roK3/nuGHVo/2YYnqfgipGYTrB9Ps
JvveXWAu/tgtZCxlei/2tloWQDnN5ZieK2+KsdIpme63jaZPG2xOVrWJHjjqm3W/O3eUF623cSJ4
xJgt4tKbcVdwzBQEcp1o+Q+bNKZzQqALngiqIUf2wU+B9VOdWseMVQSRApw6mdzbTnkb2IpsEZip
80N6DkTOVQhrq7NgQm8AXgsOGXnKcl+vocoKuy2otW26pdjCxpERtYuSJC7iWGRf8zNYap+1MRm8
fXJbZ4qIsGQkDZ4yiszG/uyqWKX+NfzkGZgKpK2Qn6tCu4nRhzrzf4i6sEt4qAK3+DEVq951IYpy
7wu40aPc+8KOf1XXAYCLeg85oDtU6lZGd/fJ3dSMpsgLIfxGXur5mYlkrhFMuxXRFkNHVmYUBkU5
CbG52GyovTAQRyTKmqyYPlb2XXVwu0H5fAzI5/w4hRr5Ut7bwfai4yeRtKei0U9P7mEXzKZ21USm
AwTstLLtBrQfMqGcmyP5NUt4H/aJSufY9x1YzPNH0XqPsFA8jRX6eN93O7zzmdLu2DdsObZyuYTC
1wwcQAOaHE4ckgoOp8vWOzTVnpcHS1uorz6bNf5tzPzkhMsbwCa1rK8hj31Xq3TVco6On8NaMxR6
LVyzI4M4A+uSFYtlFLE6Nc4jqlUJb5msmkxfomxBX5C31ElNUGAOpBJra86WxYqfoEfx9jLA2iin
KJ1eDw4FimI8H+dRLtN8n2tXJ5MKSzKqG0aq6UP72KTZ7qw/OsBeyJ6YPpPtVEal624rxQsFv5jA
Wz4LcivdLF5bB0Jz718HMLKn2ehOZg6EdX5dfzP38BcX94kha7beEU9sZLyrq9CwBx/KAKmZ8+to
O3Xv9locOttXZS42Ll4KH3NZu/UsT4RJEQQmsGpqPzi33fMzmf+fs08RPs5lAOEwhPhb480z+oXb
0gqyz8Y1LmI5v7BFuNONXGd3EXgi0SMO0pBkPg9Lsf4f7J81Bh+vMmBpqTFnlmwlsXUK7Frzdl0g
m4kDY6nnmGBPwvClDLDHJfshiGcBnRoorPEk7QJDgZrVjHbgDTS+zBeG4mnr5Jt6pqu5z2NByjuS
XIlFZpX9metTEPTpQMYAoIrNVSmWv04PPw0VHBCCnPjpbnWlutM2samgCpYn9VOfvG51xI3u9mFP
rLEmMVG41vBPZ/j1XwqnIrPj1bTmxqcYqNWwBWBgvpIUALucc5/SjcKfDxF45+JA9zId1MG9nWKh
f85EKoFGHLZS35B66KHIceI/nxrRlBvn/UXL1iHrHod72yliUENYl6GQRQYNyde25UelW5NoxhmH
Mfh+Y4V65IymlHoWtXjbGmTZphEDc5Qqq6VkTvLGmGemjR1I/fUvQ9suCKi+iGStpQbXL5GP6Vw/
llR0iMf8tdicP5rPBk07uua180z5pPNVM7bFzouYsJqEgsoVnIxE3VPYPnQX2O+qI7MPNYs0PQlP
rsbwPLudKvpjMEXxwdLnG1+ihaaxQOHlKlc2QpjCTFDts16Jn86cM9YaEzzObJtOcXJOARBua3BJ
DBH97+rOwkXN+rEfOfsl/1henx61zjxeNKHd+Aup+LrTgukUw5kHxQ1xzE1wjYQK8FJO47m0Cj80
HKT7jH7DQKcuAgcxfRWBAMC6MtWTnP//NTgpGT9FNpgtPC14ZQzJjyF41+yw9args9rOjoJichQd
JFWtrFDEUhpMnJ9y53mhcdmfBsyTrtLBkfh0UfC7FA7DDh2koFE3xyYO26Yqup/SUbKf9pA9VZpz
6XYsM8gtdrhwEhrux6h/kGrWeUM+vghM2+Khozl7CURUbb21VFymhKwSqjFrnl2CBFpuwmcfBdtE
dD/tYYDM0rnyae7kMTyAs5bDau3LmY6hJjIC+VXV3mtHtS0w17ws5XFS6XZYSCpbD7O+AIr1RCYq
gJdwxJg9H5PU86cKXpxm4SPX2npGDP8EAxiFxm3616F0aHpR3mbiTkkhxDhgvSFymrPo82SJyIGq
x74PngaZMEGKoXdbRfPvofRXQJYOl67pJAWPuZG5sa6LiKDX4clF3xHux/OK5NUBwIOhHdGgIunl
Rh7hv2OvC1Erwux0395JtinSD8NiuFZ7VBfMrR3uLw/EHqIM0oBx7Bh5L/knQ8giGb+gf7uJS6i5
I1fDdWtcVquV8Pg/wnrxNigXOLk1eDScxVCMKQIQCGnAMw/njEVjPe9jDOn5fB20gR0eVv0vClkl
edu3Qn7UhMy413NpZl8pqcp0AFj1IqGnSTXiQ/lBsyajXQuLqsaYmRuh9wVeFH4bAAzB1sBhukph
kpT91fMKCb3AJpPNo+PhvKSuRGGLYYfZ3lp+UpSZR9KJG0sxHpgJJUOHKqPh4UC2He+KfZwtmTIT
FxHx5YQgekvbBxohPBSXMYbRRTz6o0j0MwwfY2F00Py9ERV7n/WXtOUxenAnljDu5pdy7kU+xruP
hzktiw2b0P3eFbgCsqvLvsueL6cNzLsGvtIMctTKh0zmJxYbBmIMyFvfrkcuavAUlGJ/ekv8gm6H
N/mF1YiDqUDkB+NxscDqggewUmouaGmm8/fRp+UZldodNw8603N1Tdn/kc/5idHW8oRs6yaytOvl
pgSp4fG9h9N1wJGGRpjshBA4RMfuzK79+89fTwH5a+kXuM5y7LaaqLFSjPvkX1ocOttPlOqHJAIU
PeUJKiJ/6dwIGvHYS+vfho37P9JfBTkE90PMT37GifkJ16/VpbHTAv1uwEatRBqckIiJklY2qGI/
yei3FFKFjuBDSv0A2YX8ZZOltICO71MIGoQc2R2SJSqGr5+PZzREa/LEm3VDSenaaohuqvwSnPwF
l7+lpXI+a9QoEcLCbE015Sw+Ttw+p6ys/WQ99bSnqZwSyQr/aY7nmHmFHpJN4fcTbxGAPb4u9+o3
ZQDZ6+drrUfBnKc/jKafhqsCYmpH7QTIn5NWykDbUNjJqzV6bjg/e7zfF9wQNkX/mValK6fsPUwA
NfULVK38OLOeqoui4v5ohT731Lvjw63T0RxUo1z86aIN5Au91Pz25FYIj/vrq2O1I7F6jNdnPOPX
vV+XDx5w5vhCtGG8JeXFSu2m899ObDxKwjNmA3Mm+YMCMPEdcsCaQilmUy+cQr+bdw51S6/IpwVD
5MwGEGw5A43K3h08vpzkdSSkpE9b333uC5lL8Lnw7/GPqPrbB7CVgOKfJSI1fIEEqCyeuLrXF7XN
ZUKb0IXLR1/Wnu7esKb2G0PGPXoWr8yQZuJi118+uHrpbWm1X4pUI8d6SJqnJvn/fy7hVqh9SN18
R1vpanYmF4n43vnHXcdEnIXKI/06DAn/8Omgdq1VhL90DU5eABwrIFQDWJR7QxuN5OSKfuKuLfAY
uRsXxI/oPwfa6QTkNHp8fhfjchI+6wGi8Gq1941szOr48qfohLYQvPmNiCQ5LV94BudfodbLYP1Q
6hs86YRayCE4gb7PbulgefnZ29mfkExu8SGQYaJoSsYJLoMbaYhCtdoiyJvFU0j/v+8JOtiEcOVO
B0Q/aSFGUUBrc7Os1yA/KMk3SsmzC4SuEKNrBZJ0YBg4F+ycA1+WqMo7/ju+a9hyQO4KwsEG2u0b
MzxI9YRXgYGjUt6ivDve8PNojaMAJjSIeQcpkiynbAK3HldKMR/Sz1zo5DQfnRlnkXEBRygsqcL4
jtfPK1JdnDlie1MjFqDbZMLgSuFkpW6iR+Z8B6gSxToiVmbxbLux8VvWJGDclTr9dwA+Oyew/f8h
AR0y58Lyg3kiBcYI/oeDFJhM2HGAbADvdmc0RLl4K9nCJqZ+g/Aa7p5ZXWk1Qm27iL3zPQwRNtcq
/PFCS8g8rrWn1R0w/4Vc7U+ueBQ8ILXshnQGigtkfbjOScQX0R/id3huBaeZhsoQVe5JO3C4Te90
2YSZezbRB3k5V5dR5784+b+OrXL5hlUBfL6SMsRtBUa3XaUFhVkgcZdT1y/zMnChTHnBNbtV7TuH
0dANdj3AXUUZY0AZBCtD0a3E0meRvzT+IuiZpNxv7gsusBXZ9K7cqLiyCzsA92HqG8tWkApYj/V8
ACp3yZ8rPzcLtHNsSZIzH4EtOZM4tIeQuq+6KKfZfDLTnRcgNkY57EylQ1+ZR13HDY3ZjJ0V9wDW
6s2c9UfJQuXqchziJR402traUf22pBiyTTrvh10dNSXxsGmSzNhgfLLBhrNHBgY0sBWTTpq3cOLe
McJUZl9tkQCkGYQK5e2Us6acaGuOEEbpjasUzeUw4S6bfV82vZel1lS5tQ0ei/G3Xj2mT5dQxexV
c5YqaYFVdo9tBHGmZ1qLKKKlzQ6fLExYdLiGiZrXzc76Fv/YQEnwteRKFxGVuSHZUlj9yOkQ8hgZ
EJ77OV8G36D38PSZe+1Bm4CagoRa0qT5myFAw/R0bGTGR75DAA6THCSBi/cOFGz4JaGRa2URH4VT
JbnX2LOZj7bmSnzV88j/VxhxrRqXLgBNN4BKBj0z7vxpa7yxGsA8Yf4I4Y575Re83n8Jy8tnj1/E
qlsjx/kPCKnMIhI93vOBBvrE2GwVXQ6xLkb7gh1Ov3RffSaOfi7dhZvc2BLtzZZQ8nQ4rf/XWeE5
MkiwSG46FaDQHHDPXY8blFDbLi1phVz3O5j4pO6wVfW/JL2+uF6YGTMOiJGkzoATVki8ydUrmRyF
rHPTxF/jelLFgffhXRPYdYh8GXnAiRYqQKbA0Fs3e28eakqxO0oR6mkqPZ84wiLfz5+VEITVLqas
2gP/FIYbI4GcJSxvg8FfP1/IH173oB0Ki3PR/zA6AmcG46riMO1A+EyobcbpJ/QZLyz/wDMY8GQR
b/nEpuEjoESOnVfcvouzASRryMsZnpJfFqVRXDbt14//feEaYfaH5VffScBFrLNUPx291q+TpsrJ
E2solyFOG8XZ3d6jAovXYYfBRwbvoG4L78vXT9BRQGBHBjEA0CqSN8iz19jF/lyJUALFbuUq+ddr
9/JVlU3rJw0kDr9/JIvtk14cUrU5fvNn8J7fMf2wy7udnINvoJLp8xKVoSZn99ozM6sahDbGi77m
7rr0lWWKZRBqKM/RGovlesnjVJQ0TdExXMuubImElbcpWgaqvgTnz31HUa9urWRIxXeac791Sbdh
KNdwK8Y/M2Je+LSO1j0zt1WXdI2RK5lT4z4J483RmS8REeeEodHUeQEh29En9oMkTYJoGQlE9UTR
MuZtYzNQNG3NB26CFkI2eFZzklathjOX4UVZEJbmJHL10aok+h/HrYbKbXlYwGqhS1L+7yUAs5F/
vD6xkcNuBERiB92uW1/dmBQb4onp2bFyQ7ERV/68lr78hvPDpijvh7hvAnseFRQEsneExTayE4EI
XYXeBEUso6XG/VUPKipcmxUpsMwEgdd3umBat/YpbGnkuEtE1AGHdrFXDQlw2GCcARGxIiD8V0sQ
qAo/BkfB5OuPPklYJLZG2u8TdAc6rc8sr5l8H47LK9aT2UolG2JoPPVI9+NuYT51qGAYP2oet6ao
/u4lDrIq7ScHPwQA+ZUYomTPnPyvu+zvMirXsQNzrdjTaHO6PBigWk5QSAcvaMywGmCdqtsoUAhh
yiWAcFTTbzEsisI97hH6nC8aLO3EIbwxlPEV02GQ9gpARppKW+BAXQ+KKi455yetQmgAmSBJeGyO
faFULAqTLr6bwTcVdluFkvmPeGUjutwlXM6lygFrK/cJK3Zoqa7KEkZwd9qfbavLHDS5eUe6XfXY
6juv1TNaaaVbP5AahL99QnG2mNw8QjGVqLgcX6NvihURo68Pf8S5JHrZdJo/KJ8pqq0vyHzkGXio
u+GDYP9uo6IdmNPS+lgE5poPcFssruupfuMgthBRRhhOR20v4ZYVnagRiTw1gFtloHl3vvC1xY+k
LFY2ItXSj81jIOFKiePO5D8XBqzM1vXBrt2WWupF4F3w8Dhoa+yWFEK+43uTJ0DAHZBUQX4d5Sso
1EiAYr9LSB5u6pnCnygMswL5KWd92Ptmw8cLbNOTCIZVcsSycRwHiQTQN4aVX4EwO1aFJ2TdPNeL
ZwdL1KSr/HAZr6dt52toy5BiB2iNcKKPuhWuyyP1gPBUeHk+/b1iSC3orIjV6S56p8MdImZTmB0C
k8tpAxyka4n8N+Eyx24+HsFmpPUqxgckSkQJ9J7BH/KfEQQphJtJvQS0ZgWjl62oL+cnPgA8bugr
EImhm3PyEPMnHTecuYa1YW6tT0XWhKwh2E7Wjjh+rCzpijWRUPDBnkqToZEhkhQDfP0JNoOHuToy
QT8D0Dpq8cqqdW8ZUW6QY9vWQ3M+Sq+1+zEA1AfkbC+C/TvxX+KUTQgrZETg4Y/SNKv7EDRZ4InS
99PoEcI0Sf14EpMPf05iCE1f2zaQX6a6Pwfmy6zW0A3VwLimCPrDgAJ9S5vQM5R9oTxKtMn3w2Wz
+itWRXqfj2nhaj5fIhDckdSoRxXWbpb6RAQptojh1NIgj6wneLoTf+yih40dzBf943Kc87gAHSy+
yRDXaO8KHiKl7h5RLMuybmY9ZV2zYFpS+RvXNn4dHSo81gQ8KUUoc3vWY10nx1F1OzzG3l4rCrlR
2RfzdrSgssHUyuiZ0Fcf/QFyWVaGaM0G6pbz4XPFamhY1ZL65ofAkNe3JoxVdQdYI6UpnF/fsazw
vlXI/7Xaa4Sv8WIv9fBvr9BmE9kYrA7yDOl9cv4MHpxOBitkTTViTeKPu3d9ZT5SvnJMwXDHUkNT
IHZvO6UMfVWnJHdPJXeREQr2puyPNwO3goKK/rvIbF+I4ZZue79/VB5p05kPSi1snko/jLsxTtTI
NtPt4e+7pGJQpb8E2zP9ChMSptP5R02i5NLdfZz+0Y0tG6MmuYJG6KMLUV/4SxUJlmW/ysx70sK5
tRygNdNJkgkTwIX6wsdt8Qv4tkzgSeGwbLwjiE6CKxZYx1yMjWxyW+R41jiSEnrK1T3tMfaVUC97
3EZ5m+7RcmW6k0iqU0EYloxf5YQCLc+Qc39eAH/MiIRIgWS3FqeYuK2N4/ENCXEVi0lYJJ3MCjOI
bqjzX7LdquywFF9loKXqmm0T1DuIGxe08UbAIsotefs/ncLZRFockt9NRO8+j6jc1wtAygUtb4Ma
kTXo0lbs1uqcN5UEZuuMLNADoM1eq7+xL3sjH/459sbqJ7wXUpetNBPWqCr2IxIwueHKAvRk0gSG
PPDU2sGwKIvNms50feneV8Lxjs8ttbZJdrCvLuqB0VcVA4Qbzl4lMZ6kmJAAg8lBdK9bNCIJuK4w
6bTYpjggI5qarByZ9Bk+Pg5vnLIZAcv5ZykiIpGbXevUfOEoVcqdtR+JQIyZxJcZqDLhd575ZGdg
naWE13rJU7RmBskVWRn4tLNYEYYMPfB1j462OU/D3W4ZRxzlLpJlS0z+CTGgErtEPfIOFaqBLwrC
iYy3+OFF8TlbRC7Jua6iofu8uIEnaXHdHM8IfQrTiny5xWM9RJo3/L6o56j7yHgWo6DuixnN3pVz
9uH98qfUsfZpQxANX1CklteTkGSX7qpiUdfnJRq6RwJOAK38aee7lHjGXAQGTQIWrQRbosbLTo++
W+YUm8EGEPGTdUAP/ENvwvI+sgtc8SmgCcNGrsOp6QmpWtzkIbru/QK97zOoX7NUSLHFtWFvVP1I
g0DvfLgCosABChWF+STZgDsHjmTNiKx1m/oUqvL+QjFBOSRnrBjOXvZ6xYbVgi7bJiE5ssoRbftg
CG8sI3u9mDDwU8EaYncg2s8QOIevaA2D6BM99ZfV4Tzat482xZ1+YXlLokjwCVsjU9OR5/2VsbaU
7EgFm5z1T7GTVj7kZK3yFdWFyi3GP3mirSSSx0KByBlguLL1jHnaw9Y1OXOC1K84OkdOYai/EMlP
M8Tk8MsSLWqZ97g7DZej0A+rzxapNKgHj+Ed+fcdFQ2nCx5iAMQ/imT1jDnDlQM7gYNIve1OyBZ1
J8mOzVKblKIt5wkMyf607m8Afw67alIan7ngqteGBOKO5gwKsOdX6FJw1UfJ5yemI5TwxOlybB4H
37fZyAWkUedyYxoZw+4AMrFc9/AErevpopdksjIoV6JO4bASvZCtb6w03DJ1RQulyHfc40URAcF5
9ENnNXwoUyMcFZs/9cRcijZjmnCn/V+sAcaA5hOQWn91Ey7eutx7C3dDqQz7zT3sxJ5g4n3ZAiCS
pamDXCKeXh2HkCB7Vjv0/6IQYn41kCJUWYh57zalwen49ED0kjdRzLWmoA5NBQcK6a5YrWQQ2Sey
BsKqz9LZ3NcKRq3J0r8XaZpm6OaoxhCCNmEh34DxoySrPEIaCAo/2Ds4kmef/j7cjen+sEkCoW0k
IeoNKC5yBCoiBNa3c+MMpUt9qD9/w3qZBik1DtcV/AChQzw3/ZAcXyzYMKg7UHvvsVK6X04m7IEJ
cJhpuLtu/uXrS8sDIp78E0issvxqW9GcTW8RNowF/lng7d3IHWnHTdqlSfPz0gPoZ5cC8fdYipK2
eRxROPOzcpCqJkGjxmn0VTXynBjGiDdzgoAQv1ZpaoP5Swa9UYZQ3jO7PJGIM1q7t76LtXT6MqWn
eVybNSAITpFX+uo0FbkSVBLaLoXwsCszA6MlljOsJGjSB/ROTy/ZUiN1Z7Sv6u1aStaTNYTj4/fh
jA5O4JGugnMi9wrrG97zllq29E5xMI7GATVqSzxVBtkkNqxNEqo2OTalBY2sNn6tN1ISb4NzyXk+
FmyeBlefruhG5hJ69cGRxltxLvzeEaNntiXtICYMCH4crlXv5ui34c1fLgISmnSintGmWpMCnSDl
V36hZN7TmUTd0Ow1JGVVfKLtbY44nQl/u6KPY24pD7sl3G9ia3Sb1CYzduXDxM05hMlGa9Jk53mK
/z7fnE7lFQUWXlN+XzJETPH25boRPT6NUAX4vPg/tTQVWklt50FxmsxVLfYVK8Hqq0Q5rULNrylh
nWUaVX6PR2Ulf6CALuIPEaDyLRxG+lZEgG+fCqZcuz1lJIdlwrVSZwZvHLvcIyS89n7/XNluu3L6
GIQ+ve0kB7+6YBOCdS9Zg0p5TKisz2xMfXhDlbiDHR5Npu0yvU7rwAT+9BBUHVVN2uOkTX3PnRXY
f8GpRNmkOVpz/pd/APd2turw2WzTt7/0Ory66F+Xk/cKwASgHzKuoNVQwHbcFEYLn8/49VcdCHQx
JVFtdoXNP5uiAw5b2WlVBbsgazVokpJrzU5dQRKUAoocaXhtLGs1gJ+IUxZ+17g7+Wgc8/jZsqeK
UO6v7rxzf1xlHXPOPu8P5xw1ua+atL6A7Fwi6sy3JfbAzIJ4IA==
`protect end_protected

