

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
PpoeUczC12+YQ6zcBW/hk7KVg+x7UTioMUTG7QSkaE8DKLm5OzMFnRnSP2RdM8C+WL55mLvLDYfA
5lOC4Ruqpw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
K3yZ7/h8XZC4VnxKqSX+X1dWQEKELq4EziAIjvSKKzex+MM5ch0NyAGabLWybM0VZcnyA2IuBQRw
LXtEZmU52Vw900CqGAC8j1ob1JJokunlfDgROKOp9VekmhrNu0zlywHl+eh6CQ/t5W76EWfCnLXS
TKcvUxKzMPqBkiVg3Y8=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
NSAGB2MTAPfuv2AfQtQrWIP89UNTneL4Bk6/B2TdOO+6mmG5j3iveazvIvg7qIHwAqHfCGACbbAp
fGS79Be+x6ilLMPgwgbPlwYl5oARsjb29GILZJJbq65kaBdWWJCFrRmIDIFHXq65c5qChGV/7EF5
BRY2p2sjUe67cd7MFOLVO0mKHurU5wiieT+wdpbGs9uEgt/pGFeQKlj4ch2XzN03R8Lg3KmqOC6w
j6pa6lYe8j+sQMdh+WMN3EmYurAN2aA01NOtdnD7EoaLrP3ByXrwCKFB06hQfAMKudCun+42nXbW
17uiY727vjm9PIB2xOmQazUdPEZbwz2Eeua7KQ==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
NPiHNhu2YI6wz7attBCDx15tEqFL81ie9/7cRUJzlr+aO842fU7+GGF/JOlqWsuQg2RB92onmIR9
gKmj6xIVPN77wRnezyej9aQsYy3bBfOSvbf7a7d2lZQT1pTZcYMfp3xveVQ5gTGk/1BN6rnnT8J4
QRALHC2oqPHhQZ427wg=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
aHttOHUQP+m+tZmSEhqIMk3Jbc86fWQ1/2LKPbbHBoOHb+XyETCjDqnDo9IWfpo+m+LC80obW4Zd
cXgM5NoQ9F1AYdG2ggcdGNXeaparpheOz+XWEe8nirOAN+Ks5VYo+yRWYwO3R0Y+0V6Yw8r7cd48
CXttfKVhu2QOlKTiKegYDKMRGhVyrdNkx/KDldRFk70rkBceBbiSjdBniOrozyhG2imBoMkKkCmI
8TwlLhPf5Ra+r8wceN6j4BjOnyQ3EtzJgw91ujnHo20MZFiaPiqLQIavDgBT1y7leXT7TIK9Z2uu
L3Oj5XHzPc1v3FMsMkjnu8xWqC9pP05Ha8xR1w==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 26736)
`protect data_block
/XvKHXGUTikRS3LwFop6sNy5tz8PCO/LED18g65gyUXlTFzEy5+5KaTMQUecqLpCyFm0cNDZUpHj
kquObW01A+40TxBG6lhL/VXmPAZS16Z8VKlzjA5AOTDvEmIJm3FAnUpdblkc9l4H4DH/SkT4J0Pg
AUrHnddqWaJpi8DSPNWBqO0MUrawkHbgwaAUyh2ko0r5P2MlvopbQ0GN7P/0e9dJhjowbzTC75nj
WBZGaRmy2cflbRIGbFD7XjXYxUQnlQF4cr3RzWdWy2DHDWf05Kl6rbFj31Aryrdk3mgBXtlGkJFN
m5zr3GDjsM/aKBahJHrS3qOGPCXovz1q8q1j49WDex7tma2XQMF1EhfV8shvVEIzFLEeQeQuTT0b
XLKMdo58xYO6K2Epa+2sr18nEYhU9q1E419tpkHM/A3Z244kAyDth5RcLy/IxEew7UKo7JSu1MSD
T7CHTfFgCh2uzWpJvqO7gNsMpG6cDE+TP0sXq/9jY1pGgnTfgqVAfsxpqG9LCBqQcEoUbrFo/yqD
f0nd+lmVoA7uMBr6X7L8eHoIRR/yqzgVvV5OzOLYecSI7TjxmZDS+7kLMtGeFMkPa6ylrIuTC9pd
PARRXxCqWtw5MPbhJncyA98I0Cv8ozgK5Kbxw/LvS8+YBc3fDkdOWvz4o5BZTziCKrJoKoz2D9ok
0lONoqx18IYmXBAa/+xJtYjSkUQH0db5ZKQivPlg8ww79bCkqU9iiyCxsnvRY6NqNGFMv9W946DQ
qNhgps929Ab7oPDKzfA8KMQwnGn68eLferD2jwo2k0a8rpVandvCLEeZQniJKtsJ6MAOdhNFGiho
j/UnA/z+yMW53oULcK4VACZRFgUwyW+GuX9kvXbeT4IyfVPLBnZtAUySOKSmyWlHA18/GJIqc6JI
SZwKGfmKaEkjwYZJd+VzBmqN2VLMPeyU+7+vMfPHuRj9R4lgjd6t3zoZqLwCJHXRS80BALT4CZJw
9HZOSVT8dx5FvIg4YpMdcOChoSSvUIRwCGUf3RaUzfTDdhVIEF89zleTFh2TMSPsEB1GrvCSP7zX
yqVn9UfQOoroaKpudNe7nwxqNuljNu0zNG/QInyajRgZTk19vMG0NubhjsdMkXUCtx17Il8wKrLg
ThaqrJ8fmyCppuHPEhUvHSw7DWTz5AHPhOMMiRwEfVyWFdHvqyzQvIyF9A35oZvCZAkRoBL/Cuim
zd30TiNdDkGGPAXZGYy6dvaWKdpXdB5MWiH+aUo3tog6xmY82rXluQpepNeV/Ma+k6tj/oLxPJPj
DTbfLdqjcQkudqNCN8dOJehIkMTSUpHRENRoh5f5K3JtZFJTyotGhHj7Wlz0rsxtGZBnuaT6h8RR
RaaFb+wNYJlGm2hgSqJhZJyoIQ797GSVxT8MJLB5TPX0yLEjer8IklL2c2IgzvEFV14AEZHOiD+f
hZHrdhiiy5ePycCaTl0ArbND5nyorwerKEJusQZQxEhUpebp4SO2Cmz4rPgfrqBcASd48tFVIT70
Kq/RTwfOVBUyk2BSVagbP7ulVwEhfwKq18wkG0InTl3dtFXnHLTUStKBl0TFxjsHaxhocWYiHjZL
0XNkEL9xSHByb4faN9FEi7QNfsRgLh3t9h8Qnuv/ljh5+Wm/XDuyjPnQcqBQWc+eGwX4CcIL1Wxo
vgCxRvhZNQfkS4wWuWmpYppAz1zMCiOoc0FIdi0D16fI0qNN0u0OsruhnXRYZwQ6J9YT/KLlSNaM
e+7r0PrYQRLvUUbnaiM89r9BaUXHlNgAU4IpEXFPLqx9XYGrLE1B7fuz8kU4drgTLLB2ViVkCzYg
NjPe0DvPFVMDaoeqpnEpuFA7Lc3JsnY0iPP5FLufLfNMBfQy9a+NAuVTPVbmG+PSH4ALWhkDo+31
T9wUjqljLKxf2p+I/USW4a4lo7l9Xk0coFMZKo7XetNZzKJ0366xEe1QHmZpjrZgWo7BLkhGv4Lb
bpvsF+FjbInFuyBSja5Uyj5F3Sq51wnF9BL06BzkDiT0Yp/BTpm+kTiPAqZ1vbnoX1K+/A9y0MkA
KZSJjc56QK4FuVLHFz3zAood4kgGOBWpy2x4Dyalq+7kLfgiZnDM9+0oDMX5RNYbMfS5edDzbeO/
e19lDlbPCvHfa8Xz6/r82Uy2Fl2FgMPVRBNnbPdt9OMXD/58Elf1x0XMWgEwaed2a987vonweQxh
ZskuKfnf486DXfgSSLlFEq9O3EvGDKhYCYf3bh4peWYtyg7QbpWFafe6cOpfwCh/nPNF+snD32xq
QNYEdDbVtRyqqhxAMScndJPdJ1ukvTct4iXMWTckwRhtbT/fjIIyDhby6QJ94eecgLE6mv+ODbpZ
Qgol4T1n8Eha8y7Alp9W4g6NgY10Ky09hepWkPRLhezxeYYjPzLM2UteYIYnOrV5V1YxqN6mH95/
tG+l8n4PM1dGxjLbXxX8Y+xdzj1m6ZK/CfJbrx2P+S/dX5Ubp1UDeNyJV6nIkme/qwdN6wepJv/o
fOv3Pyr/KJJwpDzVb82pVms1PSXrEInJkAQDOcq2nPbxlUL57dR4INi1hmRJQU+M/Ysf1DDHKGou
yjV7MWLqCQY1jF2mCR6HMQMHSyOnFGhvG92qrypqLAPMGjYdwHXSURby2mF+rY5THbMdvLeJBYHK
5ZF6AbmSxPoqHmPr2A2HbwOUEb6Rm43R+XKIR59nbP5kuo5i0vsGWG29bXGC7nrilNru6y66vL6I
PGYofRYzUPcUMbYGHU7V7MJiilIbLxfTiDl2e0I3T7J9iDfG8aI3UTohs7gRXEi+qpQ/PDCZZUdh
ZW7W9WMYZWXNxL0UxkEb09SFS5DnpHbgL81FY8Ltf5/dQE/uL0H0Ydwcnv3Fuw7fmx/U1oW+PVn/
xfCNXzOvKhTA1QtGwQyEzFJCKZ39AKmISJgFNKE8ipSVP0f4FKivp4VBc26mBIL73BoDpws8q8Gk
lty7gHN+FUqFPPqralSagTJzpoPCrCiA7LUYdF/Evb8NcqxfuF78bZEq5noLKFV8EjHH4vyJQTU3
IyhE3PbY/J/Ba0Z++F5CtDZJH6PlZb98hYmSPkHbAEblPvTIAD9e99B0bRWuJxqjYenINnj1N4fg
MmGrDCfygmAIcqNbGmm+E2oFrlRQl7XhcDtRSxmM7KyLlwF93E2jaCpqzooSyQ6nrEfOHeSrMu1h
CjmvkmhLfWmj1Sur5FsoQ8aUku3uvKoEKCo0U6FLQ5CivxLuWlNXaKb4mZpLl18oWz4aDAE0AhmW
7FcZ4DDD2V/9OETaCaKrMsnSoVGn0IXlD6/HlC9L5sgZdIla+YrF56XDA3N8yxDzJYYn2bpf1bZZ
p8I3B3VrrJobK5MUVlOzBDIADLn30WQ3Y9X31P9Jf3lCFwvVA1/0cFAdAyZsq4JWJWJS7rbH8x7w
AsCszWQaEj6ZpuMJMwk0L/z/8ZeITcwodjXZ4FQ2hzeE+t59ohDmj0zNAvW1HdB6jHltMnW1aBBr
BJfG6F032X7Z5P9mKNoXQMuCMqmeJ1IsYkIXh19KEUjO4/HoWvgFsSMJKOzEGDV9k2uee+2GXEN3
cZikARx6WCf5Q2XOM9Z85ddWd7NxoH+CmhWAtzDwaf4JT1H32dxs6y8udaqwgR2kibXG//raC9hr
7bLrciUabxks8hbOkeB0hxLxb2W2banBUundsjzJ3CMRs996/H1SJuz0nxzG3jYVsSGBufJ1KhCg
ZDtY5LfM5LkQ1GYkzqQZPRCy9aNilyI+7zB9mtXxcJYiuL6WNyFGEVrP9pOlrvDrn2cmf+dUMdGD
dBzsyWtaRXA8zZ/4O7yA4zgn7EgQT0s0RZJWdvOkO7VCBgGhbyUGh3tC32OXMtRLcf15/GAr/z+l
AbxzIed4yrVJknlWHDpZMaHZR6YBBQlPSqs3vs75x7DjhF/sYrc/na+R1qOSrVmc2vHCxIYcU58U
wo9NcSIQdubRiYKdhS1lzGeiIxFmvGv17dIvS+OcarUbbjEc5XP8XKbnPSjl1ZvZltpYodp7JWB7
0VUedg0F0s24g3xsGIUDzTGYOdvUmSt4t6cqyB1SNBuDmdp1ojqO14P+rK6Zeh9a2AgFUVx2vEPh
GYKO9z4/pokBcnM0xR1rVotvy/AolE2raRzsVb/I070gj3hPu9p8feC5k2dOuMHg6fmt3dcP3uGn
gKZTnQj1O7v/5l/fg0AR9kH9qmMqJSugifH+QxE06DBqftxCn7+QUqKLk+PU7HIM4FcF9jmJExjn
0ubPre49PVFCCH1kuiCOYNz468MNOzOq+ZUyacuEcG7nQ3HL/QHC2d4pxhaUdnfpm/z+t2llCClv
UFfVLaGUfX4C/FefaYyPEnR18V718TsgXdhNqLjkTAD2mPzD9vwb0mYlw+e4Gc9CJW0KOIAnCvw0
4feo2Rkg+Ap2l8uzYQdiLu54tl8vlSEp9R4/Xw0DCAJbDvNc5xlAPp6K/2UdDXVIm2Ai5+6NpHxz
RMLo8vounjuM8uNVLk+xgJtV9ir4CX94wx5nvN/uKgG0ZYx3Ga8ZPHqX5f24CMABlb/v5onpIZ6e
dRlMb50t478h9AXlNTbLNmRYZeglsF1Cv3MHae7OPfqfl/a2mtJStw5jRwtmo0+sMms4TZYD6DKD
Tmo3T2ymFoXAJFVaNTBIOvvByBQzYt9Ajex8qPBbsf/Dj9ymeBu91GJeFtTNLBxskbOCuxD5icK2
I6RHbVPy3Kl/WSoUh05S5IVpjPsnW3r9vSqhZuDxdV7ftkFOJdJNXiTLuO3mxEDFoksrq14CVI7R
GdRdEVsJkRMNGRTwSojwNVN46clCjI/rqVu5po6I8rO7sAqR+bMJDgDNjkZFPJtBnuFe4i5F/51q
vYQOJphSfO0jHbf+i9xm4Xf31u6S79IvX7/67ScXT1tV4lR2xkOIZB/xSnU17xG9BiZxfHeFV1RM
nSE/Erb4fotL9DcRyZW2FU46I98g+hBNUqc224axzuqQax+6ZkumJPvi8OEBlkZdlkXYAmI6lDa+
spSF5boVn6W7vGLcyQf1aBM237OYZxJFilI78TxDX2scfEYtbSkFLZ6pOK4KsHAyJplc5EI8/PuY
rHW6zd9oX4C3Ku0jQyJWTbimOP3vUnkXCG+TW3U04FhMr4DKTjJ1WfQe6eJWtqETit8O8oeu2Mz2
uko9BRYUaANirKjQf9htYOsuqrLNxFk0eDIZeGj3NDMjk82yrrcOd3t+K+lORzzkYFvyhQARJtiy
uQXyIcj2YCpaoUPufXYjWJX1nJyJ4uJnAHleHkh8gT8aWrLZYabjAJvoNwfW4c/OoeZt34j/qtlx
3rQARfuyzl3X0KQDGxqdp4mEAPjzb7RTNh75ezMu9HgCgC72/xfYPQvequN+fVOCv/LczfFULnht
fG2Cvth98mfqYWrQ/Xc8/reqrrTfz71eu+NLt3AXPXjP7gOk80163rxNpos1Jq5AuwdVJgMb6E9J
QpRXNW46VufnG6WskjJlegcWQF2kFiYS35YVqORY/YInL8nHA5KIqPoK4YdM5u4m6UZtcCDn/oIV
z/cPwBPv234TX/ydEBEH33FK1MfqtAwsXemub2w4sk4Su5mPOJz0GwUGxrY+dqpP6JPGwO3aleQZ
R/3ipiB7eAlT5JQaIDPtWeCRo8deCLzcKMMTMeaqgIb29RrLh3q7tZf/3qtaj9hlMrlSRyZTnA2s
eLVJCPrMHxFoS7Ep+Jt2CAK9SO9I+CpyznDk7Rl35sIX3cjKMW4H2J8+w+sYePwvOHqSTY6BUgIb
H7xTFmVjPpb6w7+8sR6zYDYJEHoIUTYqp5pdUz5jbCraYblQ+htLCqu8zhZCBVUHb+eByF8C8VTv
9btYckXjnbxHwBBKdTt1CHKZK5OlzGM2ivMlNm7l5hKkcHGe7cotaSpygu58U25tL7zZd6gzAjYh
ukkdfMDbJEVL3AU4P13WEPnAcwyI0VwsNuc7fkOuxfpceo1sco5plHMiX7MBGlGvDnU0OssZTZkX
+32XOWynT4AujFKfnhMSkSqvh7RZzev1VSD3adzVhPrQemDwMAvT790/oiTNy6lRNAnGmqkI8Ryg
ZVkC2UrbryPosfKFCH34kWPmNnOaH8BcQweO1SABCSTNofo+JlfDmV9cTfZ9lugWiWAFoG+pa7ro
SSMmfDWrNa37a2OWjMNlxJpfQMbMyRIWg5IgrGJP+jzHyIoaGz9Bs2Wuc4cWkqc2ahMz2o/Pr27r
xCbtOC+C6yI0CTbsndyvVl2BmMubCMyLxfH1ImThf13kDIB2mp2Iu/JS26HROM+eTH2+EA0meW7k
UFVC+vhKlQHV2fj6QpRwcYKYHRIJFxvcwyFMQdK3KeBX5Rlh1JTmQUcqM1WzvUXh/yzKrPyM/bgB
Fr1xEntm8M+eJdzvmIo26Z7kAXciISNqSwxwed2nbyJWGz/6oaHtZ7MZbwZX6T2pi6V+smkrYY7i
lv0oCTAR5h1nTPWjJ6mPczCQA6m13/6W/XJw2joXhKZnnRurCDSG9wQrGdIzcw4oWLRf7t+jr/JG
C9Ya6O32h5v1mlN/tVXGsGEakebHZ7pToDLEOyFAjJLwDJcmbySRTQA5VkXi8ZA7svvvMMKL1L21
BVJxCwoW2j3LZRMVIL2prAGCwc5yiAigvMJWI+XKClb8wX0hmTSeRssgqHHQvs1RL19mogppuo3q
zhj22CMS9vXnCQLGK57HX+YXVudVP4U7pg9dRvx2dKzwLzjYAjYYabNae+viL6+yt99vXGz39HdZ
91I+vYLl46pd47MK0XGSiH/ETjUKKpR59wdZjRCAdZme6BHvUVhCwtCoZD1a2DmQWurPbCa+iP0Q
okbX8GW00nBAwCswct/75l53UUQVHBeaSrxUPDWKE+kzs0+nszaMOWiOs3884VwrbdlwqdWJkncW
joMLIQxKm3a9Zh2qC/3AV3ra2LWQRHeUuADy7+L2ejUvXn8Pz/uvjY2kuUKECJTtv247PLpVjGrW
YHRqUdEZLuO0Tm6gB+gljajvF0tn05cm0och1UMfHHZ01uwdhhVMaSpQMQnzZ0wKXUAGkX5bSxgL
tkTPvAbkiGa3EqwWq6ZOeCwPi/UAu+zH4sZtLhLbK54e+sgDUjE9fmQurUPJscFs9ATz8cKwioYw
9ONokks8DP1oqdXy/A0QFQu8WHD4BpSKF6szmw7hOhkO0LfRb46gWWCym+o5qqyXOiSnQETReKQ9
YfGJbyslrP7Fj/y2qU3rDckukFEP0QdJvY53kws5g9KtEJisVd0r/equPCW/+OZUlviRlrhwVTcv
th48PonFfZboDIgCvLg25KZU8dmMQWHdBf/UXkG7x2yLSWekNH8q2VcdQ44tBGYsFJkgvqngQ0QG
K3IjQnUxt701gftUXMqM0TaLzYZCZH6LkS9eTrTVdmOWb4SMjO25m6T4wiGQaPT5X36su7RkerK1
/iUadUSrhK94KrNxyIQ4/nhjgDx055kLMMCBiK/ZWVwr0+c1uF0rE1ATWaO5g+bt0rDc1IEkhwfT
D3hIk7yTp5igv7Anx/iScvkUEh5J3rWzwC+dWLH1g7c50cgKayZEcTJzOj3x07UZQhTefTdOYQyR
b9ICs9R+C9RlMbHey/1Pluxl2bB2FmLz7xMHF+WTtlXpQNXFRaf8nskpDMRA27ysXB24USXSkzLW
9B1y6Lk2G5bGTEqnMue8ueRD2cwZJrRfW0Rt4lN4SiifkKTbXzl/arJsjB2ZQTv9fto7rFFYgkwx
N5n4ki8y/IaZ+rExM0NFl5iHk8dqaum1G2LJHXtzQwfgTSyWu0HAAXV8yk3ZQi4NTEm/ElXrDJNC
S+1LAx029xk/apS0UINTyC6uMEVj6G3BG3+28ZUxB6ADYy8HR30KFMKPP5zjZpTD9n/stEF5HTx2
spjYpLEuqSBb727MEcSbSvVWqGlUlK5pp+4c3yaIWcX9e1h0VjiESM7y1+O1egpW5ws0ywfkFxTx
xFUmonvZmhXiy5dtm9NbeFiIOhU0QcXxbyV3qK54PtX5Q3jKXnDJul5UmpZU4ymNKPct8TOXyjq/
yD1jpKRXM9aye53RThjuqZVLyCLUQi3EcsfPJo6ogv/ndotHX5k8kXMht+o5qG/l1EaJmgGrMVaT
bTkgd3Vf3Vh0GD7f+6Ufcdym+pJ1FdpDbK9jjmyvuAfdwQuMlxqlHphx+x4XOFdFQvPwedgiy1Qk
hpGza33quDcZ6jmdkuKwD2h6absAfXKSsRDf/SnTQks7CFUZmWMV1DcqAfj9xEbN6xi84fJTILab
xVIxc526T52Z140BpvP8SlphqLfIgAz2WD24g/tjevroj0OsHYjtZeVWvNCtw0ajtROp6UQTA7UJ
UMIAQ5fACrNU1iQEwp0qwuIMxWwOcx+NjVVzrIsz53zBWKkgWtOf8doUmeZ6/A/nBeobDhZrwdqA
c20l3CZY36pLQkihiJaqEAyb7WMJ6NZT2RtfdCfkrqV/hbRsA0/8S/VT42+jaJVDIgw3Oqq7YKPj
BGJlnQZW/GhqOem1UKApxuTjURY5XM2bMC2+olGmGrD8tpdpbmFcTz/2pCjR2+QNIgM5Y3o8vr3M
G1B/xHTWGAxbgIlcQb0MF9nUoa78/Prf9t+VooDrjAOpYm6G+Ni5h/wKH5mRSE2cnmhc59cR12ox
t0jwkgq4GAczQTKMlJL2j7bHOifJovAh4ACvR4slIwVpE3q7MX+it2/cwa86h+DRhfdl9CRuimR+
aTTr/eYmt6ZD0LYg71LoS1/l5zdH7MSf448ECM37X25OsUzq6E5e3rKQnkjYSbdWXCKYNOahNKqi
S8oq5jZyoGkWuSXJjmSRuGaLZdtOnOV9UwD9Lqpufa5IlzNZFm0StSZNrLXYJ9jTYQBSwEfjmlcy
ZIAKjktOeNB/pqXpt22HANM5mVTm0yGOa5WlcmivCa3VBKJWy5XNrQ4+VBGSuqVO61ybwVopKx9q
jYztlW4HfjH4ucgT5ORbKvwbh6MwsoQVLdqPqpXA/rX34z6VRIVr2uEIuCcM1zHLx0EEkKh8/SYI
Z1Ax0+Pu7RBz8AKEar4eVunWyuOpC/OA/CQPFNx6ym0quUp42T3nxV6k1O+Y2R9k1Q3k9gdziEfx
iCNac/SnqhKb5yiq9vJBjqVlMJMvQMmTf+AuAmqU7cH0Sh/D2DuwFF9uINXQIHndebk5leeClsuE
9S55ZskUBl0813ZCBF9LdfLqzBXnz0/u1Mt8rq+3k8Ko8LNo67PJ7nVScIyx+EEmLG30FQ/pLS7L
dV5bo4/IZ7vQMWPqWkl/xBgPLivSNYpWb8qmT2FU1XNiSvhRveGBEm7BmqXfYFjCJykWJjnjdVNh
rQw0DK+0InEVoeqf/5BP2zjiwIPR0dRlz4uf5YeDhX/uhNTOvCgwXZ0gi+Ak0pYWI2Mntcrw1HdC
uY/hYqscoCL503vs7FBLCbsqqaytk+B4uZCf2at1Q7R7D3EGRc6RmXb1jQzmcsRy2S/l8aT7PMyF
wXW8QMw/81rUaH9ATDfFo/2nmeWgolac23GbkFauer6rosUOQV50nYT/99zfzLjJFoX0IAJSeRXi
5SeAt2Ulx1nDT8gMfZgOWzOPEMcZnP0PLjUDE/txI9EniTrdIF55jupJYbZNzHzsQY5lWy96wS6W
JQv6a2KIw2sg4qOIQv8R7ycw+JRxhMHDM0RV8tkI8A/nQxYqYp6VbIPFyzKQu3Ytc3akYdPKNnQs
l4xCugnynuZpAPpqbx2AFdnQhy3EZh+nE3afuq3GmeOI3FjJDEMs3CbPtD4i6wmLxwd+DcirH6qa
JJXlCfEZaWRScIj6tnbhXYc7kAdRY2miqQHA1Y8eLPk+RvFWSfJXUr4qtSV88HOBm7XCHoJLj48A
909Xb/VUQJ9a6HlO8LxTXB01ph1MkzsvpRh/UZ6d6iIHZjj0wqPuqYGdbkSPgnju6c4/RWDhLtnO
n1BQztNpESjwBAiDfeCy5+HpZTjPQTkcJSIAehQ+PbL5ZGrfJ0GZEez2KhZ1hz5DR/0qBjzsXkbB
4HpX6a7QL/g3p3LR4KTHjPW+1wH33sP89FkIDyMcL2Vo1QZfxmvbgamfHiaenM3PUGjvEXmtlUYn
7Pi4dRW5P6erU5ir+in3aLQPxZ0xW8FBECKAkkMRdzP6iA6oDrVHpArmD80Z2Mpi5+eLjiOmy26m
27r5hOtWtkxrhkX5fgGlVIHoiyjkbnp+kRqHuVfWkq4jbcbmmVHuG+MPOIJy086VJcqlYBIJ1XfM
FfNhEVOgVojpCfJQMnjCGbsDvSOBft7DvC74IcSBmwL9Y1/3GIFBq4gijwQ3yGPXM95OeHO2l4Oo
S3z6NIETYQxmwO+7ChQx+QBVaxUcESoeOyRU3F+I8fukXOb+TayyKo0DWdGPVBfnjmbOWBVDgypS
Z7B9ptU+jB88lhgqiOq95Il+uY9Zc4P/oQqY0VnWrQ3UF7wOotCec7UdLjwsCPtQyWce/89wxK4n
fuoCK9NJG8JZ39mX776XwcbcCAJxYapcxunkXHz7ZtKXrYOpr+Giwd+oKdp4jYkMjKxgVMINiFrX
tdtEVLOJuaybvII+wmbOaTYZmY2+jpLzNZ3ttiJHcTsNJEmsc2WQXccazXR3rsISW9c4Og9iBqaO
2lUT4guG3I1W+5L3BEGeZPxOj2K4CGUYDo+ixGRJBm8G/7jTINGZXhCx5xHsH00Y2vT0VnZgGeT4
gqMx9T18BWmoq5cyiCPIkKOpdDfRoAfYn9UZeV6iE14mCIZicET5pLGBTzKiBrm0J9IZ++3HJl3m
+y7IqQzuQbhMKWuP0hykA9cYoKBCF1zQ0ewqoCe/qcdT5+PEkkVP5ZG4svsNSyUVvB4oJzZJKTme
MJRJ+VTOW9p7djj7Nd8jWxny2TzIG2SCw9gddoVQWZI/WQXVpA/QAOE5G3iLfG3C6+Cw7UxcYHBx
DBQWrLicos5YhIGhiuo1beHbMcPFmR4ZLiOIXUu/Zg6wWXJOcFAsHd0zSSVgCt0PlL23akB7VKee
dZCNInNFdC9hTp6UW9tzeAIQ1lAu/TG63zCoDSKrR5SsNct57Q39b00DyqY6peVhwvgJRt5FBrPV
PMfymH9eQg+NSVZC6YXxGfgtdA3P2r4Nq7DDVf5qpQLdGhM7hVRW/FIjV8XKzIRL2198ZJid+1HS
lbS5eBVFyVyl1ERB+Fpf22rwhXyODVTbd9rt3U1WPDJx+UhfnMSL94uN2wm1YwhW2+jljFISCEVp
pot2gkp9I0kgK/XuIBK5Gj68MHlqaxUkS8RwzzWJbqQLUo26ilIocsv7HEStlecBYXfBc96+NbfG
Ffp/su3Mw1FmuJjjghEHqpALsAAgw4ySYWMko+06NLMsKOjfMWFL0UosJy/EY9q5m4B7gL+S/n3L
GDG3hucj/sZqPGeIdDo+2AyCI9OmaQP8miGQk+cC1850P1lmDfKxS54kDWho3QgTfQ6YIhcVrL7C
kI4ykOtoO90eRYJABEA8TYBNhnWlR+ibJ/wZk7AVVk678yJnqKBaSTzm3K2jPOC3s6sPEbGswelM
HABwVO96bGpg4eA3zRr1X2DSjKUn20NWQzDq0t7q0NOCI4cgK4FZCR9cOM8iwxQgeQAwCrblKFPe
VR9mHPz0vfTQDxYf4lFoLtAMdDdD/mjTsvx0hBhxGvAwPPXoN6NXCF+5A7JKyImHzvYBVddz1YMC
q959/Uj/SW/ZqQKg9+/8XkZkwZKS8sk/OuLDy/BjtlIFwsEvpqc0HwXSJoWnmesKA/eUdFc4EK28
BX+cIopxkDs66thiJFO8If6l2gDa9+5WPlKKKnsQksz6HfZoJAtQn0zy/v9m5d1d86ow6cGWKs7Q
uDFH3I3sPnTZPRXeKkp2vpPxR4LgxbzqqE2Y7uDhGEPIRwCl+5AGSCI31zm1fLvrmDhx8M1ovqsX
tlDEUX1AZLqBqiIMAuy1JxLPp2Obo7459CrxEB2/EIZlKBrDlCaZ8W1oHOmf6PveB2TXizjm/mtW
sL6jLOnuCNJG2+PNin6V6sIens6htIB7Blc0yMe4VrfA7+d7zFmOr3R6/gQ+gKa+YUcwE5DXQxPR
moKtzSAXpGOWMG6J3/aAZbJ8gLgTOZ1FsKby/V/dCd/S2uhBr1yqcdWAZj4wDGLjjwzo6jPpYx3p
0HBJbYH0MOHsTFuVMehxRGI4nItPbz1Qwer+r1EUl7YGOZzB2W6u5psmgk9x0Rm2ZZzrMzdTmvxp
Fj4HpPQtxH5CmAkqlMTIr7u2kNjuGf/448ksPbnXhYyFvxc/QKKTx/DMJebiFsODa//MkwhghHPH
nxpemvJ4FpX1PO9gDkp40E3qNJasAwwJDJElznbC+5+XzVxyzARixF3VRtNCVf2Jfn5DHj/LiaAo
l0g/xg1o4ZAvdWo+zhdJmkboqp2Mfr0Fje7wxq770n+u3Ncv1kRtBd5psTH6dmrNTQB/PskE9xwe
z1KKyrYdhrMY9cPQnslH6l0aHtNYbAZZkbLfbhBI5eUZsNoEYIxg0WqatC53X0bWvD2uAzjPSObe
q36M8Xw0Tz/0Sky8Uum9RtXMzhj57pQx5PtjFB9/heIgR7vuK0MztHz582Tf2cI7ZnGa6NvGBfhl
pwDfiij0ggiv8xwEZbGblEgrWYhNoAwGfAA8C7d7sdU+HU6O6/OH2i7TsLSh0Cl7+iYy7HPUPSqe
Aj307bamFRwnEB8RuGyALzQYIRu0rKyEI2Y6/yhvMG/hIT1rcJamj0SCk7jwu27YHK+uv01vfpxZ
N6Mw48B2X979RYTsJ0w+3I7y7XKj6w9T480LK+ge372JQE4fVTfDLeRNYSH2m24JLJw5QjU7tLD7
9QBEZiXul5Ba2CKevqg4Swq9axlSQZDLubQDhGUfLRu4qj61V0zzfh4oZEM9+jS11GFk0R0dQfM7
K5mdqcxKGjkjETZ3iSnMPkznicH3E8N6gKRUIRyuqoALMw1KwcUeEQc70sxjU6ZIqpGRi0I2ye5Y
A7Z+eacQNSsHay2tKo/5OIiIbq3aNdb8QB2a920nevilDPczeUK+dPTIdLH1tBU1wpYzPnbsMpiJ
6SSfrag6MQGfIN4S4FR+C+pXvTe9w9/kDOwDF0z2W/JRsOMqVKea7fPZJ447PtZptDeGg4sjqsV5
puvcSjzVAsIoe3xclOJWLZXpkolRjuhVqsIzzoHTOVFPRqeeO0yLORFHsa8/yMf657/ohu+9Ikxb
b2gTooFWBYJrCUjCrYEjhuPmT2Mq2AEnpRDtGPl0YZEWx87U3hS9+b2mta/B1JCbbCyZFA8/k0yM
XL7wzUjJDIoGjjSMsSNj7/UpPiPNuqxp9KVppix1T9RwWnpv5XNpXQC5vUBcAVRcKvbutgFrIpSJ
TdT6pXxwJKdaXVCy47EwrZVb3+iuqfNqXn2zZg7Pt3LkozC8FALLg1lv3CzJM2y+O5WhJh5vqXw8
zuy+V5f2FRRa9M7uc57mTXbCzeA/xmkTc4Z8w/he/ASBkD631ZZhitUA2dos3pYYKG7X1CeB0hs9
655JCjtjLaz5gFHRzCgS/F0FHNaH4OM1HIKbiJ+viJJuFw/XKDLxxMtQvYzvVWk6MjROCtlZZIDr
P9T1cbQuRmjYAPUCuPdSW0Ym8ec+wkD8TSxskbYw4GYgA7nS2O+PZkYP1APXjKlDq+kHGNOzZE1s
qx5TkeCxWlly5BrFp6cJKY0T0DLse1JsMZojF5gRExU17+7RxwFalBPlyCuHTTrDHvYVE8PRDRou
ny99gLtg95+cG36W9bLPY0eCOy8Q4gwQNYyemznoWR4MbHPJHQXEVK6qJa7S2YPnhMRsiXsUPo5A
d1M2grI++ZGQ4COTsCn/8h/zs5lZZ/LJ+wzW+1yXfpb2wEarnZGiU5vZdrEjEbTtyVp1Gk1XXCCe
BfAYm48eRf7am4LeVq/OZMxUTpj9KsP7orM/+vrCoPBubqF9fBkkXyuUU4bpAGcVp/d6wueSxjmj
MdPc3m42KzM75umXT1dT/06/pmmkK5v7XILSujXXw2q37vF7xDxHlMNUncD+M2b3gVSN7RsC7Nzi
KvxJ23k33LLei3FX+4TtkBWRnBUQKzFdyUul45YHfspBV2mW7fISUfWT6UWIDDw9p3Vj1INyUEK/
mDiBXbmagfDcK2P058X3eS7krOKLLUELnMogdRJMpbFC0Azi8zqc2U7/F+G/uyuzAS6Jc6IGfPwh
8CsQk68yF21aFdeR1PhDfHCAEsZWDmRnURidnbtKY0OcfHvigttMKyuG9kzncyxKkm629WXBveu7
cZQV47jgnqM3zuas2J9WsBJh32KYUVpF4T6o7r98wW8jogdHGpXnZJbMRcSE5y/A6Rxk7B/l/asG
G5puXfN85RSySigkX//J13qyjzVAus63tvo7kUE8RhXfwoA+ImikdH2jnLHrq5s3HMFiGStqo/1c
CBuf6Jf4Z04pTILcX4m3Nw0fLOHwHb7g7J9nsg9rVxdqOENifaw0IKX8x329X3zMGyJ8jQg4kKFf
lV8/tPbypZLE2KEtTpfr+/2cAsh4+nopHqs+dTqsTN1Dw250IAov+IAgnU+PbVZyVwbhzOflsknc
yjAhEsQcU2mOIpnZtSWBlATPv9bsetyPWkuygLP0XhbJG8HY6BE+55+C4DKc/05UkNa8u6TvQhYd
O0OW7LiUR/zNMUp5nMhq94pVWA4c36hQ2mjiM1P12VcAyXCyMXj0OREeUZFEUseGWMS92Uo6y1TL
2wHBa3rvr/52tOFJ4lT3zIa3ylsV8S7go9ZwZyZY+jj7xMbi6rj7tTNwTqXkFBRqyp4sT3D9aovd
TmyNGI/QaS7pLsAQfYU1dsDSnfV4Uz4zFe6B8iXK33S/uPNAU1oNmD7mqucCvyO7vikufxgxFFkT
QWb30QXdCsrajbnw1RxfYYgF2vH220xxPptq7BDMthVTDUVTncrvbPaAnxIV6Vfi6KuFVH3nrCBM
t/kZqOaco0d+uqa5sBNVLR1vVIPmYp5eWy1AQ8HSAiFQR9oJmKbJbJC84iO1QuZKMgsooMYIR8Yb
LsUm/omCPFXMpPsmmBBDVxFuTkHa00ICQPE3TfQj++WqSQsOZWIfQOGLt9QjEE54C3mZ1GIaieEa
/SL5Gl3WP2ZArg5Qr1qBrzitvRIi53md/eFsMxp5kjQqeGiDJuM7YtXMZAsPP/+Wg4Jqp4Qob4fy
xDzcKiYakO0yezkFWACNoRiUBQqkHniObdyASl9BYAjZ4Lk9ZdlVPUtER1k9v1y62YdeL23ccGJO
+1WdagpVjnm9RJ6blIYFc2QDPD3p7OpoJpdk28+Kct/dSHfDjYEJ2nlJSdAJjEDwpHj2Y0pkK/IR
EHQOlermjiZg6OrLoKLoEeyara2w++ccRjKG/fSD91+gDT3gkC0slVAdgPrrAN6rkwneb5YReD5J
km2pb8UuWvaW6r6ESw6FqdWdCij60L9KtGz3LuSlQZIFlfPxf1iHmHIx6Qy/Yf9Y5VJ+zGa38GL/
Ha8p/yVgwbOsb+AQgXNDb0QMdpNA5Y9bmMT5zdYB8pljSW18bGOyH+wkkcko3n8tFEmoybvIEJTq
xbHTXgXsXKUEMsndNXqz4uadnAqHSGTESNbLUisJO6o3QILUom/ibx6kwV3AXDhMG76uKxrH2qN3
TwFT4sUmEFnOyMueghbzdxVRhrH+wYDHGKQo0tQDaag4gt9pZthmpjqC70h9XwxkUqwcrH4M03B0
vbjtdKSP51qqdYsfetOdOcs0OWkQwNNqREC0jORarKMZMzMdvKFTE0PZo2YAoFZT+eRtcdqgelHl
gzMp2jw9Pg87zu6vIhDu9yFfGlYoUzmBUGPQBdSb0Emilf2SjKW2rWUd7tSKC5uUI0azWGu8UfSH
O2b/AQiK44HSW2wQ/9h6HAT3A1H77QbaPoMeCyyz7TR2qd3fSGVsXp+KJ1xoQBaZFmyiLBfa+NEO
NMJTYNSy+rGHFxGJXIODukGVLPyRNf9cZfegL2+CPqV+8lYcHjj5uQ0yFJltqg8IiO6CyvJslcsy
e6e183XbAYZqpoundLbrdbd4c+oK+hSXtz021BSG9YvZJ5R05J1tugAVBh27rDjzhSyRqFEe9Pk4
QpNvrXLNslueEBuXm5+uboATJREuO1K3QCUUWnpH03kngQmx53KJ7FgXpF2E4CX4nGeKPtCM0nMu
BvmgHNVb0eS0zxTF3AEaXGis4GAG1VpiB7hu+LPc6oM9U6tVf4lcNvaWeKYf25lo/RWEVXX8ZjGM
rUJRIoqUCOvNP/0TG1kzOva6SRuvbzqQrEbsAon3woXESicf5lg0wfkthYx60P3itbSvylIphCJg
cDgOZCofd+4dwED7lsI4VgLRpZ/ZT2lNzSXNjtDDPbS5rvhrjwnXLHbnxlnjtMV4jh7FEoMTa5+c
8iOxtS3hk/dMkg8BDqTXhLQxWAHiznrwvNHrbWeP0p9h0pEslnDtvdISyhs9yC3GieBhn9Oq9hA3
OsyyneBDCjby8BdMwQABTtXIn5awtb0YY9xwT2ueEeBq2paCdKCZR/1bigZmA26EvCFRDVq9fgk4
JO861mp0Wbzqdb4EHm4eUYWJqVe9gaznBTnbmsyY4/l6IVjbyOXTVr4bg2fd7SXgy5feWPWblXNu
AOeguU2ZzRBVeRM4fkGr3SbX9l5fxYYrpcpY+fmqCkmwU/3C/e9RDqmyZSwzmvvR/M42KsTLhWYi
BNI9eC/C9TLgdTgURv0TXCQL7ozOkJr0xQclDiqGrjN5O5qarPuyJxlhdi/AjTLb2rZwtxhcdmS9
W2eeiRovlVFvUXCNQKNCEXCt1EVVdcXikKud/1y7TVeKL/52JGrszJY98G/h6xPtK2al/znJXMpQ
Xz1NdTaA5Fe+1WDaDDqCA7HC85CWfr8IEOhM363dEfixGIUwBgZ8lrG8KjdcxK8PA0wKWZ11H5SL
2pxy2eXiO7D2ssU1OCZ04w4rvNuga/G9q1jnU4K0sO04okBbaDSDm/XCg5X7lruDPSJhZFK+l+q4
ks1JYxzubpGgTCgnNGfTKmfhJ7WbEr/lb+jlUjjA/IizvOYHW+2v7MGaxN25/P51Fug9ktObFNgn
rk5eSzEzq/pePhrfws40xf4XjXUbivltlK57ymb9nH+PUOVqnTx8xD0zXk296JT7Io+P8TDTV2Gm
RD+mPvSMfJ49YartUvB+Rkklm85SxnZTj2cxHjrG74z68fjOAhk5f8wLPsIAn6EIDsdvjlxjFacT
8ZGXYt1gtIZx9VxkW6E/mo7KO+6QFiT9zp5LI2FBcLJkTQsNWBSORNcnb2Y270qh0tw+xzPKPegi
OGXaKzktnrlmlkU9o6Wf0x7bVxAaCUEr+JFFqSr6l5OSF5HqJRtsUNCKeIBi1MHBjFSO3iRxHpXF
Gwfpr/FFcq/d03QOnVfycd4SKzzcM3t2dL9xwjRqZNeQAEiR03RsCwg2A5rtSQW1RHdwJ67TcRhQ
CKnw8muNM8TObjIGE2FF5uXFMmh4ta08KQYCrQKnD6BohjxZexcBf+mfrh0OLMPzqYMhEe3nezsy
b8WSSeOTANQI73JcYAf+K1G2zA1ByzCHTraIz5tNruvgoCFbTs5lkcvELnrS9ReMUJj7dnZ6L7FA
NhLjOdxZ53VWcO3oguXP1F8YI/Sd1t+HBYE5tiFi3+qVmKcsrdIrkYgkn7PBOkWUsv14emBjrqv0
cj5+6XduVvM9AS0Z3HPu0vwjrMfa8x5eUbWN/J3Akwmo8AAfRDq0iHV9czmu8/D0JtUvBOAwPtMt
TbMW0FfZpz5ehsCDyBBkEsxUWvZMMMYY6wsx3hzmy/rUKxCxOmhEjB0ZGFerXFo6CFMEfXDWiNW+
GdzP5ay2DR+Td8iWD+PpgzAlZDaID0hDvnnLaiYzZ9S588LX857LNEXj5lZ5CWL/hTUYmzYNpgA/
br7wO2pHnRYTpR3z3sGg9TEqxgoU3+XP+NzRL9gvTNpOE6RcblH7HNLFaNFD381bfUj6S5Fw4m9a
D+l24cjVTv3Xafui+/I9fmCj96v6aZLC3GUEEB325ezzEtW0VzMtgHw3Ebrh8+UayINmbxukzY4H
YJDQ7Lcx0Jgjour1ReFrw/JXKtJjDa0NmDlzt8ELXcd0ZPZS0cwb2GsFQRPGSR6Uug9lZWLd1aU3
R57p2CKon30Q31MeN3TIBQfdD4DuB9f5yYDE3BNHT3TfqrYerb4XjmnFJz2RO62a63ElaxZ7P4DJ
4GLjwSTaAKad4ISXg/XIQhx3whEqDLINJ/6PhcVVtNAIt9ct1cEjHiM11aQSxEgrzc3ZhNO/yDpy
1ayzmvmeKLBLPmVKPZhwy78JfgdiGh4t88rkNj6eZDITyz+NaQXIXeCQ0avm08DUt1ARh7sajANo
4NbjOYN6oWJW27z3NdoE5ORlKTyWzlzzpi03jldAXZBhlOSbaoivVqM03i8jp/tD/unh7eJZSKzO
P2060ymAxOAC3cX2TkUly89qm5qfieV/7fS51deGz1jwlOqdDpMFETzNsPsdbur5pRUynUTZCToA
A6pP/6pIZoVe9BJkYZdP1GwJ5/bubUO5J4kBWMWzyq/6q5Srbljz7Diq47dzMZ8g1gGWF3hLlLZR
djaLawfGNmw+5S34N5sTKgQ178xdxMIvcqAIeFy4tGi8WY4aV7u6VaNtm0KVu7IXbld1Lj+2llx/
dl9P5DFR3grAgnKOmrk+MmLB7vV15fg2oTx8wMXPXRHzmZhTtfq6pSc/4aKRKj8A0ui/rrlnSsT4
4aRuLMzin6iAMf9Qu/NNoheG39ixFm55bzl1gQ7NRSps63ZisF+f8SC/pICcXDkZlz/QJw4O2RaF
OQNb1SpoqzUBiD+eh/tN0L5IArgxYoGa9HVktZeepxn7TtbIL7QFrVCxaJ6WJPqIv4KM6Yfkq/7n
73TeNR8UZ+qzScKFGbeSG9Y+SoQh9GLU7/7Pwm46fhnHlykRCfHP84ATrEHwadqgg5b/wjIWFQu5
MftTEdfi789NDVMLjujbKkfqShC9hmI9CyevTs/iv6Rc13bn3YX3ffCo2aKMWjI2gel6QRFUP8bs
mzBM8YD35lZoH+alsa9mdGYwq1kcV0KqlUfqmEyA7MuITGUZYH6wwgjF2GZzamsE9uwQKajyFnu0
lL36BXerl5o9WrhcJiyvQGSLuAQ5s3OX+W72PZ2TVnr7lbsYDPTn2LSQu7dbFyaXWWBfmapEY63j
2x7klwo/Iczf+sGeFktKc6LJ+YtfxKymGWJZHWqgR03o4svtPSaiHYAYcCDbPBuuvQpd3/64hvsw
l++UbktB4LJSVoehmA3mOG30zDrrX35LFo3wK8agfR00FNIbPKuvfBSlidfJe5A8Klqr8/EH5ya0
1uW+NPsxy02kTUAc6rhpI1NxY/gGjFSTCbq9ewYWmgkDUtpaGhndroyZpMg0FcLpDMYaEguBtG37
+BceQTotLagRyu0OFub44mahR10gnHA9WYOjZxOI2NrSIc5dfoDsrlyYtq5/UJ/PuYSEjSmmxMCu
quWxIVqV5TCovqRBmKPlpY0UqBsxr55QSDJdhCl1Hh12WhGv/p/56NBIG3SqA+oJJwoqCGobI1lY
o75x6h9C5Yke/hLFI159R5orSB7DuGLjFMq2JGEtC4gDL2z4rTnjop4hHrL7jZrdHjGZKIQ4Pj70
vuzkXALV/VlDnXUC/qKKuC8dJk6yO/2ZevU+N+qzZg1NsBU8XwiYwrrY7bT4qOi1BGwAmD9qyz4m
TQpXItb2RLdCzavHVVfV/EsZ31HcHcwIkRQxk+Lb9AkqeuSfeywJjsAPl9JQp0mtr65BhZ+8DqgW
+5Z20FivfieslJzo2GNWpSaB8m9W4KRD6lqCH8aXC5ZWFzzsJ4PdWLwAJfVdZa2+7LVZ5XbBzGKR
1EduS9JAWgiE9376aO4JCnct2yjrph4CrVvtHPbmw7RjnlstEaVK6JHwRi+JQUdFZzOyiKd8bJaW
vAgmctwtBGxcr8moGIZW+YRPM/b/mg5Ld41XtkE3J7vQF+9LDUVFC4QyWE9UryLwzf9+CmFQVixd
YcVyatuhDUSABpHruuohuViH8KtuRxaV3dvOvw4brq6ci1B4jG2c2cInM60gtQwpUKvnaxpe2FM0
NQug/Olz70iPzTHklFDABUVXvNIiCBO1C0HTPcKow8PpfG3+RcbHwu/NtAgiJ7MucmqdrO0l34da
/bTui7WeHjfwC0utddXJrcVt+xJtVLNCrUpu14QurWeypCegT7BT09Se3bXoldS3zuBgbrjOHtS/
sXb1mtVZ5wdh1ey+iszHM1+gdKTxXOTvTcT9aMrXUjURFKZw7t5KYehfdyC1E7CqdcuBRYIZZ4/h
FgO8FNSa3UJ0uU+dBCVFQRouSgOjYAMAuBCdIRlthjaq2n4c8clAyupfBH7Q8IMzETrZgjaZkGDD
JfLm3ljw88sV+/FxJyUh3Zcwfh/kREU/hDg/PoEczISrSIboMERV9D1Tj5fLTImVcMabpHGC7jNl
M8BwiF6p2eZsuq0NruSlajuPk36L6236rPvK8kU0FOYU0BoDAtEkKaZlLHEygno+CPqMbSUIopiS
JJSD3J59aQocMP1Zc5ioaC0QRjWXiXYysvPDsBxBf1xcpzTY0rtJc8D2Ft51pKs6AFcOO1OwZ6U0
G7Ltyv5+sHzklr1K4POuV/LdGGFDujAbnsGemH/BJfX5WEVlJ97HAzqgy3rkjS98LaBxIyHMg24P
9EaohtbDNUdRzypVIYbCuantVbjRkjFDAEFrF2irEHqfLoxwkDMiyxgT7Vsq7ioOuW96zdsIkMEI
HVO5h5KJuxAW12EXzaxMJoqJyGSdjHOkzmtvHvdx/VlBF/tGQq/tBsXfQYBMh7UdpvMs4WSSkUGM
51/o1O6v2Qb99j4DqkvySd3wqbwA6D1mi8xNmn0pbLPoyCq/JrZyKy+/wBvD9ZfZ6wTAREDgK/lV
9+Kv6/OM2n1r8Eiws+rcptx+m0prGmRJUAc8in2d6kNqF2fkmFchmW66sxNA7v6qXTmiOqcw9blO
Za2cRTI2C23K8hlGspv+sBBxaObViNSACDo1JshZgEIGCcf/2nbonwas7bTeur9eAvCetjswteAx
2ZcYac2aktnJEwlp2fnf6Ex7bsxQzBX9FAtlC2zmyB0NOKWoUvaFNzC99XyGLNQi/bvgStsAk+dY
5Ke3Wn683K3TlSTRKoTKKVJMsXtmL1Sr1I4rBWSeyuy6V7xAKP9IXSB20rwcdGHw4JA4Gay3Z/k9
FB7z6aZlCTPSI1i+Wu3/C+0iFyLx83nogPabj3P4LxW2JCUCX43EHl7TvRilqyY/YLBRcgxNoQv2
vceVxMCQGDQhQZTvBXX1TgLo2gz9RUy2+AjJDpy4QzmV0LQ19Rma/flN92DrCFpOO59bKPpx7B7J
Yf0TlFnp7aJ56T2xgXTI5qtCoo7y9nduVYCeSAGeDruWkIrRYI/zQHPVrq+2DM7GpoWBicGiUk9w
yXp/ZpUXDAIkfhoyYwvgER38KXnMOd3y/mUJVDTuOvMcGpwTHvzHNrqxMUE9Ct772NMoNSoD6zAq
I2abUMwypENX4oeg5E+5Kc77oFjLL6qwLJtBFSo+1hcAZVJw5Fe9TPCV8ibohh8vnlGKthKJfZ5R
/kVI6FbLITVW6Lhk65eU8lGLEXiGqQpy6491Ogjrlu/fYTyyTRg+drGR99XLiXQaEfaqlCNZ/0kM
dFGZVeNkwXxkl7GLMzX4/kZZdH4r6TC4o2Wr7NjkxzR8R5VH5aFsQfcJyn5COwxIXFKkKN+JeZj9
SHETO6lWF5S4iYxZhfHXaKTZ5KytFI1OyR4F8NKYgBuG+joTkfjdGZc23D9y4P7tLHBlfaXEsICr
wFt0S6N7OQJ72PiHRokPNPeqKKfsQsynyLcQPoFUSqwj6LHG/3OZ9o6dwVPRr8xRqERRz4MPDF7E
uCL8/YzxIOllOdwFSyXdI1bCKJeIZgqT8JbvODWwyZ+Px7dlVrpJN3ERHWJ9waVwa2/GLEBNu6kT
Fe3GVcn83Xdh3eX9+1D1s4wP0Bc0euUMHPJ9Oj+327f9axvys1fxuFagdyeakN7HJFSFFDVbpi0F
pTH+YpSGL8nnJzVOQ28Kn3bx+i8ukBpxzLU/Ke8FKninIEIE2SbL6352E1LoM2Vv9qNtSIh7I4kR
3g3FoulBNcJDOG2+wNqKK3V762bCqppvaMBcWDGuzdEEHeeIt/WcVwgdo+cpk8fmG/Yab9swEsUj
aQfzjqUcVPmhn0HSBC1rQPH49vWKZFGCWNJVouC2QJ4nHCZsqdLplDQTVGXqRDBNpGIa1dataIuK
6y3lyqUCT2OESbhB7n8uZ1nG5nHkaQ34UKF4g0YfcnC/yxaNHq9+/5NpU00apVWBTz7e9yZRlSJh
3E0DzdBA87mKfa3xwWgeyHQ2CyUIK6L1gwct+7bXFWKammbOi85udfy40LwSUa60Y+Enc8UoATGW
jx83uqfFggEjlgT16f0qJj7nUg31YS05pB2z3HGDU+Y+tnivQvzS8p5Ba2my3jpX09tA39Mwb7D/
jpQTjdWeGkbsSltdclETU4X8EZF0b4ETfnFhtDOvWLXdaYLNJlkoeILWH1JDMe1SYC+zT0Jk5D0j
buHlUBlFN8EX/i1KJtG0hLA2EAFJagNrNTy5l0EAJBf4v4nKbzx9Ssmf8mNZUSFMWRu8U61205XW
x3CdwMf4A3jj9sjXgLO5bQgWJ7OpIKQ2/s83cBy/1j6KGClavLS0WWDPLbDaztleCJCOYA8NNP3y
uC4ISoDyev/Qc6cL/++Atww6wH96YBoHr08Vpk5mL1j15tT39takcyRyxP2OwquXRHsZRlugAN2e
cWhgLnCIS3yh4I3hZjn25lNuFqAfY6DwTG+VRcGw9W413Uz2WRT98KlJVIoUKOcfjiWrzJkuJYHU
Y8uE+7Te7ErPMnzJhbeGxu09VVi5fEslctMOmJXSrRLE3kN2BEy8eyACfw5WNjjFL0oXGbjI2ubz
lCExDqTDDzI7gvS2o6f+DwlkpW9DRtOja1sQKgKFj8ciX8lWEPIVa//iFpNOPuQjR7jX0y0flrLC
gz0IaC4xmdO52k+JDulWWSa597fcGkzQgQgEjKFMLBUGBxPr2KIosU5U04s/jYwzylFymr5ZugjK
HVapZv2BEQcK6t8u4HZxEcpTpbhdGkZZqZ0+ZOcrTJBHQJFjj1VCeJBh/MtkrxPuAsEnYD2Ry1QU
U/kYAtTEZddMhgNarVxB9wlkY/iLgMeHqutsKgDUMAydMcDGXyCeXFlbsX658HDICd6FElirFLWd
3kEouyuuy0CobKkagzw8Tda2JOUTYwedgT5dvsWouFWvmFItmSRYg0VNGZG01WYsXFGhO0/xmuWc
XEwwLrCuXZrvsq43SkWuuJ9rmzcuK2ookSJKV6NJPrWNYBw0SfEH70gf/qOrNdnMEH/INlwa02qK
AZn7LMN1q+Tu+cq5PgPguzL5iKSL6Rwd0KFhO4Rz8eHz7kh/lhwAc2I5bmgPmcKG2qjAC5dkc3PS
Ir7fG6IZVhpFOGY06XQHxiqPEGq70va/JFkdl1OfJzV46jJqgbxobI+XJd49SiOuoUUcl7b7iiKX
0B/VTsxLynFOuuSw+y14FtRGhE3la5BHbIf+rHgrShlutP50Q7Y8lBXPm9e9UQwVaULxC2KjCpC3
XveqIghrELecByL+iRs2a/7wdcviBjQ+VL2UD+QpK14AREIZHURv8R1vSCd4EGtwgqvaN012hTWl
2ruNFQBAhqrMB0y/4W8qy9S9kG7dvSyaYNS4zI6BLrp5EgpxQNu4uuhASkmzNnyZeEpR4zrdCLTz
33e6buyevs0ySuEUCrOZXFIDLIJ1IVEjs0Vc49AH0VuaB/GTjsItQ/Jo9L9wqKDxV1Vudf+iShhq
N9JFecpILagEfvNOdOyzg1Tl7txeiciZwK6QBjAMZlqxV587ftadOD8H2LzF2rS3UuFPg6W2wpEY
45O+L6KII4ZD+kwEbkMt+wg/r2eEtxPzOscnNhrSRhPThw+jq6ahgksQlPuQ5TtpNZE+lcW1CFLN
px/FoTZGAOfifTPEitCU7n4c9wiT6siyk1K9Rq5GkikAWllckChhAI9/Jk7WvChzmaoKAmkTAwma
lcmAaFmotlSWmv4eMrhJS8lLq3Drj7mcONExFTpAoLwDlJ6oDhSrOwGIQbl1YqVTobAQ8sDSWLnq
e+yANFsoWXfcLVawuMEj43cbWwvPOi1ikXZSPIHduLOU9IcKrayYbNF5wwZtTXcA3o496sCI8xOD
r3Nf77I3yGSZlHZHn88QT70VSc8HObhdKziKMvgZiMlmgoExJfNwX+T7LU/WxDy1jpQerOzfgB13
e5WSQTFdeDbEvYeSMkbWxA/9lc0qwuSZpIOJ82/BZpg76zl+oGNPPH4JFokEkIsj2yl9DEigu5QN
hz/VivtLDYtSWhg/xrHhOUcO8F1gLcXyohwqLadAXcpCU+GW3XF3MuYsuSh9dSQjvIE3cKqlo5mP
I3TEPf6NvZIYL/SI05cQIEwAkG0vHXA83aLzvc0N8U9PqqE6HDX2lSWxkvuVyc60eXtslTtfZI8s
KeJAtS7In9OF9qp345XZ0YaCaQl4XCEq/LYtSjRI8r9Lacswdm/os6ERetyrlYzxJneQKfX6Af18
ib1ix375uJ+GSieF3fPv/HcKOBY7vwPO08CqGmwdrz8JqyjFxPkmZCJpy9bL3oAkRYiZ4mkr0ZCZ
GLNNUdta9JTx65JUe0TNrLTS7g2qOfLk6udWhl/BjlaeR1Y99Bm2Dvw9qF2uV0fYcL1hO0ZUXYVS
nEdt9Uw9XUB6NZ69DEf5WKDUyt03dZW8eFXLHMV2NKCXhQy6x6HghKjGOE6gj5lUg8SMZFuoZrwN
dGGxdYLkeWB9sgpGOJnBH74+ii612CPzxRwq38z0jVIKzQtF1cKtrFYQajb7LP8mLNv77u/fkKIQ
coqTd9Z1wj0Zp9H196fyMr6wJ9X2kMXY7wds53cTF4YP8SCxrvxfMtdb7DAkFGGziryUQwED/fpH
GL3PTyM2xrnFYqgAOBp4bRqPThbsaFMG5OdPThp36Tm8kBcI/PxBoWwRsUM2kk63TDND7K4Rr7h2
PSlJCCTonJ8sQeY6nQGheJNXMiku9vccLObDZRHgiQxsNWidqZO7W1NNKBzS96RTsTXNUumC/pxl
+jLcB0ZxyqPgfIk5CWutVBbrIrxVX93TzO1tx1e+fVKrJDl/scXWzKGsvObmoRFXBKZGLqaHSmo1
uowTwHFzxHVupHRxLfGLYlNoYuTnd70A0hnk7gK4QDzY/iL6IR3JY6SpWwQU9GZyGx0Wap3lQ7aG
xZzS+ACdsjOVDr8IHInkrUh5NpmkVDQvKQEoIaLCJm1QXuG6SbEAOFK5WJFxJ0Bwnkim4n94iXrb
TI58S9qa1bfvHieTV3bl3U150Imj3xLdYA76Hno+DLHTo8/e+ICAbeYK+7ZifnPwol54qcKfYbHp
o1EVvEuG4hGJXEIu7Pol/CFIiTvpeD4uHLFcrZKszCvRBzlWp8fVzIoGTB9vCOQ8bRU79JdjLsev
2gWNtMXIefP+IYbcEhliqWWAEYVH3MpK+0o7jVQIZES2Xc/yCRBywi0EJyJt13vyf4nuXnXoyEth
PCzHBKLt8gE2ph+8eSIXOoCGEMys2k84FRqy3KapxJeibvNJkZ3hLL4V6HJmzW8OAMrKUsBrYrPX
G+wxNXLekX8VXXG5koDeoMDuWwfRl6uGX2by6T+rFMw/0hMokeC+L1HoaO2sh5Wg7nOsMMSNjSI8
2ULdtsdaxPEc/52rnYL9YiJztkOZPBlwPT44kGShlMhVBbM5zwXPM5d15ePT4R7gOJpQ8daRb3ss
Usy5JKVo8m230Ly/Xa2AfWBDtLbQxaGrDkl+0nyMmarx2IxDHKVoPlGtAXgA9bPv8/K3XedybiKi
f0ZdRqkuv6b6/J17Y9pu4xbrxbpQsE4YG81vWippbAClNosTdtZ/vf3rqdlHBwDo6fvI6xTTFFYG
E6jPTKKvs9sYrM+7Cf9QuL7SxJconcGKfOHXnLf1PqDDVqnLpQ8a3QkWcaunGatJVD28vSqO/tW0
LKG8/OgNGh3wxdKdkvOunnaLIyTgbcFC1FVO3gBflwdRkfKAdRzDu6SDrWqjTVrQFRCLf3scq5x3
yNrCgx+yaI3FuWPxvIKmRm7/FgiwskBOZVdf/T/BUqFzUcIbQMvXnL0JuoWRhl2bS52o4I2Et3Gg
B3ORzUm9c0FleLNCs6LQTeVrkWfaz3GUb1fL6wxA5PDT1Lt29ZN57K7jkqD5gQaBCa1GhhTl4ql1
f8bc/SGteBcLxalBqM5RCNXXNkrHPkROQC1cpnvAISoiFXYquejEe5NBjY7CxtlRPrEg+HXix2FV
LmmqaNxg4kNf9LySqDrNOaHmuxBK+QMKs5U8mMeS6yqHurVFwC7JAl8KnGZuS4xxeNRzoFFD6ZDH
T5MTl0gd1cZznAT/UxqJU8cuRxGla4eHAsh4aTnLdLRrEAnTqRfwSQ3k6tE+FSi5e+Xe9+XNo6Tf
qLndUdZXv5TdDgYLtRtNrrAzVjkrTQhcE5h+CbO6qLj72UeVe6BymmVQpSX8n51Ld+Yd6gM5UTBv
t1JhtofsiTMp8UNfia53MNnsM454o1MtM6XjGBv0C7rDBXq4qBh2ExUXN3W77/MEOIRpRRgWRyTG
JfND/mqkydMisczi2Uk8ruGg5e7Lb9qodm20XBkZYggboqseZGockxOJTEIqHqeF7s7hyWPnmcq2
o0d5muw2an/RiufmW48rW0k3OSMwlKVJfMqEVM0jPEa2HrdISp7h9n1OWMoDHX6m9B8OLSsg5OzC
khO+QKjgLPxpDeHqeKqrRGYs8N/cL9IfE5MHLib6xx0TKcXSUJr7VVDrmfcKyJCneD4cKdrOr08l
9bp5u6xKylfr3aJAclY6P7sxFUL7Ec/O3PtfhOGweUGSJe75q0uPBhi5wrJz0ekUdyc8U8Tqf6Kj
OHpCtr9uoti+fFr4YpWEI6s1mvbjkg3ekHGbHoSA1G7V/6QGDeEsdF/ugtkuV/AVDoN+9olQgN0k
XAVhymCfxayRWOhks5xaeP9F321B65hzHj2mY7LXE8IslnliL9J4UxHbX7GnW9nHC2fhpvb7VIDo
ZfbzRHRHoO1dOoV9hl0GInH3/ceToJxCEybYVPV9QSrEbUo9H7O740o6kLecbDdIcfhrUyGlGWpr
cKn6llUS8N2K7+mQgSC3IVapd5GeVp8sk7750K8v4Y23Q3jf9zhX3QpT9op8jY6Y92hvdJ3ucWO6
qXe/xYZ5uGKJ8cVSE4hMR6SxHoor1GS9nppWw46XZYrQxmElHFCo2gyzsHI9Via+KI6NoyTCBq8z
GY3p6UEFijMODdYXX3+sxfb7g/w51X8VSPtzMqkbFsLiakk7LO10Ubyo6CNcQujqlHuNbdE0ZYI2
uQeZVOuZFZ8AYzluzgBfu9UWT98nRzGQxg397fozxDOdm889Vphxh/3OUN8RBcurDUq5rmFOM6p/
K0T/Tv6dVg5PZiBABGVaV6pAfBG3TnvWPlLEu9uhd0ybRixsPoPWWjMLiOkoOQB2vtFUkntssyKC
8z/HPAD3/Hy4gS8vyE38bBq5dP65+0CsqQQ5Oo2peM//8mZBq5Lr+RmrctIjtdK1zmBSwUn54Wxx
X3ahchTlHj05n8gJtH8KJbahLEWyDXHHQ/R6vylBGhvaV2l6F+BhkM63L1OfQ5eeXV2JKf6hsAod
2O+9R/wGf3lP361+fCiaVnrlRciTfoJfyaSPneMVRgIJQU0QiA5IHg2NX4MV6R+wKI0hqWMk9pdL
AK8zpk7GAEGKVrQVD9z5T8Mc2dVSeMT1COUY4d/g+DbgfTkDVyXnVmPwI/f5uAB8/rpJz9AMgQzy
bpW/mdPiRoLn3hKK1XPP12N57342UA9tJabryW1GSOj8kAwVI5a7go1LCF+TPBoQdoYjHxIhBvbL
kSSkm8gfMr6ceJZl9unQXYlSz9m0DabBinkiQWbnj2h7om35EfmkfmAtErIlMGp7gXGOGTls2/wI
Aq2ZOssmFP46mVHJTxD5qlF5hn9W+f+7oVFZ/oh6h+RXBC2G0DvRNYV41GnMeSTpK6aLmiQa0mjk
CL3wpMA/kpgZoE1n7P7Phhljy2Y7u6OmDhnjf0wIaef/c3kB5Y6ourXeMl7fuS6ovU2UjmiB9iAK
ic1+4Ij/h239KAZtge6VtWo2bkIrEgrkOPjI0zk9qPmtvji0jfgHdVAG9PpBY/VAEm841PSnf6YO
3QdYRj2laT269xmpn+24oxm/FcBqFrTsnuEmpahfVK7Jkj39mZlzrvaOrqFlU/FnnHppDLIdqmHc
hUGKS+BUfag1q0wKZcunSMWFAtN1n2zv6FY/cK3fDuiN2OaKq5LwZD9CmrAo8eORgI1OUAaeEJWE
MO1C1+m+P0gdSH6c6wzqKrDE5MW1enSN5oJSy4ghDkIIR4G56TRmX8+9Wsa3FSw5JqynF5StbeHn
K0X7JXmI+c9CGLticPQlMxXX8+iLnXYMDM1BeabiUbstB8IffPw3onzGTgr8GZn8Ozuy5fI7Wouw
vvIRwqODv41ZWlFZCR4wHZNXwWVOigB4H323k3YeN+UMGPDDvImbhVAW+lzj8tdV8u8NK+cn4kBG
+ekdZF9sTdr4lqNKh7/fQ3enTSqNhmsMAAPGJmbXXqUBKlt1BTwunNH/w88CKIM3k2m/2yvTsPqQ
qNZ2OghmKZf8XVUjYfDkqDKLDSSinhXhfMhOn5Zntqses4bsoPN0CR81KlilWoYVTokRsnNgQz40
w2RKbAuEW7hq8DQlco6XSFEbLOEgg9DFqWwQXQ3QIM7JzJ3lvj2+4Vm98yLjwp0JNcdSmqsXl/aG
Bz2yn1Qw3SUhdk8Lo3QZ9+KzTdpZDTlkECb+Q1+ypXQaKlxOEMTqBJ+o/7ErD8NvVDzaNvWM8/x0
X+KFsI3gTtYqneXUhKFrfgNIOIkkHoGjI8EoIZMuEIX2ZxXtpffZzGOZmXcp324g0J+t+uNxtlD1
LLKDtII5fVVX4BZmvacPnm2pGATH4yFjbmnoP41oq3leFpwWlRmsmA4hB6W/E1/ZwsGCslNu7SRB
z41XsMJSWhQODzscF7slVXO0D/lQWlycEv7lXz9dQXRGisiI+0cB8CgQLt9ThD+pxsn0Qy46p/HL
7UPn5Fdk4A7EfexqqkCFlcLimCeT0pFeBimusBCb5DKAKkeqW0nU57EmCu3cRBMKxBhP4AFmerM+
S8gK8OnJJPURwvgpOOG2/DB3rfcK7j/FRC9q7XmIgdMYVPcwOUTu6Z4xOh2m3HL6ElfKtsEbxSxW
zs7CehOSRRZpgIWI/MNQnFtqxZE8KvIqLLjCryqf1yoFdAYCFvGkeKdQHcQNZU03y/+m/e4eAHpI
yR+tZVUO5PoMQ+v9loHx7FAQ0oEoy/Engzo57hdaKMxxzD4Cdi8PTRNiFSn70aXpHYw6cRYZra47
WWVOZxv3C/Z9vzJYvMdQpG4iZZ3sRb88BPBDwFxC1EI2l5N5eMxj1Aq+sdGhrg4qF9UqY38zaz22
Cjw/pag8N8/nnZdVGql0cmpfH3yGmbISGimH7z99EQb3GOOvMaMq5vYRLa1Twk0/J4D5uKyN1ViK
Cckc4wlFKwYV0ZiqLZz7UaeIQkTLUfov9U9uKDCVZuPb9gMtDAHBOUoWmSt6kpkHDUrgpnn2tbgM
5MP+6vtIV9vcu3nJqE7+UZdkE/nqq7AOlDbbnEK6grnJ/plWcJdqDD5bWGBCkeTOfrFf3qgnz3dU
DCHCDyhtb7IuW28/JmHsFetPX58YKPDpfgnLEWfM8ejGsECFtkp/PPsdIjvJvMQCmp0YEmXqa0X6
G9UgI7OwIuLk/8MjD/ZPDMsda1jVG2XBShfT6olcYKAI4zv3VHU0NMsBbsbwQWv6y0cNaWvnSsZp
QqGgQDIu5HkT301qUXZcH7y8m2DmMSNk6hDZXQIsOsnHeIXj3+/QtQynwRa6Xuy/X0GzlhpBCllL
23LlSAyvf0H1Bt69dhLuiot/p4axTWaeH4VJUykVO9sRC4U3VY+Q2tNDF6hBiiXyJg53JAXzMXIf
XZfmYIdXdWPWR42p8948xwJa7R++6D5oGJKuh66elmN+/hswsh05k31K+hBZJkHQDGvPFzNLdFz3
KGdqH5NyUO+KWM8Tb46sdYZYH7fYZnvdL2vRjhFy9Y6jKl91/hymvS9vF/YkAS17tLnWVEHsb0RB
bAW8OWnyha/6RN7U6XpvQHNGAkuurg1b+VB8osu/OEVxO3IKkMLekz9QJ9zn+4O07llRj1U6xRWn
59cQIdiOLEm/Yg4U7FR4D3Jj/NdMTlpYCSKTc43SDEQh76YUOlOqRhxxWgNn92YGv9eAGtPzDOjy
pjqrOFXZBn76rDZwRjn2nX5A63AMOHUCWhNNTu0WpaPBlvGiTJzi0RnzhmTRy06vfvWr7poRuxNe
OS6skX6JMXO0TmqcUdRjQ74PnbvF3Cg3MzB7x9aRoKt2khiLIPWZDTrp50DuWZ0I/adlvYRZ88K8
HzLRF9BNZMn4GK6G5snZurZm1/8jBYVKU6oYOxcURtuTHCBTVm2/ObAkX6EwfvQPv9M3m0YAbW3n
RO5jFo28kt+malHsuUVNewRBj3nUvip2bmQbciF9+sadMOoD+09raxrHgbFjH6KwDXKqsbqEMkQq
/mB2xSnEYffVPP9qvHunyN/GSrAGIgFWUhbm3QyTNvj5Mpdep5cYEDyTk11ZDfj3vjgk7U4sx40C
fGnySZbexkRV2iQnA/BdLIQWYnZOO+dOxUKOMV4npqoih8gIj2SlMe7f4LIRHW+SgQvDj8GCNuJq
1GkkfCXO7g7dJbB5EgyU4lEy/pZCaIsgBak1qfeBj4gSJjyjn9vMYnzv3NV4yHkG0KoI6U9V5hhq
LwQjTH99Mc2657/hwlAg86Czu3QvHCbLHRcOUKGiJDEPoRQ4R81Ewvxv5dNQrRXGoMVnZgd3X0Cj
kwhQCeBI7AYuqEOFxnblP+z7IDV19UrpLbEyll8EzftyJ7KWGIV5ON7qFTgfQgIHAQKtJnnyBjZ5
CbV9jhfNSVW92+jsathUK4aUv2Bx5I1UHrfojeGUdo0IVSthxJYnQxNkHEUg/Eypis1WWGMdPqGg
ID3PYXwkhbikU5C9QGt9W2xXZ0+w57PzMov4lACy/b50cHQbQ7SrpE1vJ9/sRJkjIw1z/SzlYQmS
HcWuFHu9733TRHENCL7S/h5jIUAGdiXvf6HacS+Wwovd6lrHZRwKjUCrCu3dTjQ2ZrGobz+tOKyA
H385q0QDa8OyxMWhDinHpP0nAtLNw1HKTBlgu29bMLHwDt6Jc1Vg7DgYfVb/ghZjDN6s/QF1X7IL
poL3ad8usTaLtAOe5dt4eCaWVqVc0Q7UM0J9EjbtDi0FF0NK/5UDBW9zB2HJzVU6moG2VF6pWcnN
v9qrqSxDB5Dk2nu87vFhh2Z2zENR+KK2lGUC0Hw/4T78JFFdYfCJsJ3818METJ7HYLjcMLkEIH4E
WOaKX+LwgJ+jB7z6v5J+TCKZQYbktZtPUktlWeYe1Az05hxSV2GkA7rJH/8fHU1AcNnDn36q9heA
vOHisBuMAEH+a/Q5XEhSXJCwkOLEyr4Cn8/tQ9CX28G4yd0xB/WP6tZa7penUvsvSf1xWBTML3N+
C4yN3Gx0G7CpwhDNE9YUw6NwLtRy1Q7VKXI66/rNkImeQ4fUR8Xu1yNlI/1EynDFUzF3Nr3x+2wL
Cgx4wIV/Nba1+1VmfmCyrFhDVFyrKK+JguLVRfgvvqzOfZHyTMVqK1MvuXYEz3bsIg3xnvOrDJIV
Ie0n0izvXbVfFG8T/T1dwwIv02noPyGsZZ+5+BkNurkUxCGfHg5JeiiTsLVIe4bAHmlA96f/tji3
PL1M5dN9Iyr7itieB7tlAhroRD1IKRPlrVVL3Srm807hzGeHK/Z3xZRrGABNOBeutjtnbprlLb0F
DBw78fqxMQAxmdQ9XJsBc8SXx3pqpctmNhl95sLGtVImmf/4nDb2AoQ4y6OFVCp6QUmQQ5Fq8HlA
PNGFE7D+kEOWS2b24wYI8hXgD3JabYrWZ3buLw57iQZvt9WF68eNY7epnb++3pDfvYUPvmO/VAmK
olG2OjfHcANJbkN/6fdMCQufB6TlXU6CJgngM+vIMm4nZlfVZ5lK+MzAKdfnf2CplSCAx18O1Z6j
hXlfK1zDDtoK8P5e9Z3BGgqupJQcg2HR/b83knAea9w1xq0nz0Qg7jHsz7OfnlzM7x3zIOZRathB
g107OgAPOgDvuClWzUMqoV7SbfJ9GsuQo2vwjEvQZwFdxATmScMw/z+LSTPBIaVVuYmuGf4A1uEs
qNelRv6/O3wrX7vOZWkiS0+Nhfoc1rltAG4Kk61nJzxyA6rLQ1YrfBfMutV/cFvSWfnG/ibq+SJf
gLezUx7hfN6rCjfbhXm3wQSqPykG6iICkaHVEMA+IBwkAnHcuvprd0KNvOCYMZHhk0YTqO7D8vfG
xeoStl/Rh0us6MXUDNOypJfinbHK+8I1OQ41JeSEAqDgq7OfuaXICoA2G4MmeEMB12NKYFaY+T+o
xiclcjs87qFS0Hyv9ionlZf7k0JvlCqLmRRxf8CAyODnZXAXey2q5Q0tVO+2qLXyqcp1haW6oatP
6qSHXeo5Bl7WU9Vcnxxde81T6NZqFrjlPHLpPCEkR9etEfdtWZ1lZzR/B42OXnDfyCyxEdXHvki1
QisVdF8306XS7O3iJdFILh/Ir1h/pLmFKCGOLLM1x9yHm9jbF6Ue23kwqCGBctzFfW8p0S0uF3Qh
swa7p4bPfkbZHTZ478rAF4OakzmbgCnfvzU1DZNP8CPgaHcZUx8qpfy8sp4xZwXFcD0YwiDlGIDg
JcdbMsboxnPsMyzx9UXAABJNedYuptcjNawoR5k419TtqD4NzBkW4FoaWnpGi/+Wnm1ZhYQP4gSc
jd/0Uj3IchjOVisg5tZysrAcBab/B+RpN8HGy+lcCD7h1eywHqsmIUHVsssdcdEAHBN228X6goq1
Le2tBbtfHGbjyIrVEVlzutFytCnwl3uymtirPJVAMSSVotdpXzl7xqbmcdS5nj2D85OmdItpwvzu
S/+O2iGspsp4d8OuILsi8+i1fIQaHka32AdhW0ylXoEH2uz1lX5JfAV2a99VLaqBt77hRJlxvgI6
lMNI2xn6zewRG801CX/O8q3wrwQLk62Ry8gljQ3wCvDKqOqlQiwVf1IVP2Q6O/zPbjJH1TCmfEPC
njYmRMoOoIwAJxojfAUtatNdWtHz/TtqOJ5vSVhCpJgRkkbtY1/rr8IJjwAylNdKodrJLqA7GW1j
Rh4hRYOTJCqb/LQghMD03S0UGzFi2zztaTdssaUhVrONfVw/MOEw8XuEDR/u0rMLaftPQ9CMYO0Y
nhmexracDkRiaGPhRtqokuLhcNQj4bEaOCLQeS4RG+pef0aUSEBfzA4/yG0LgEuvQxbbVrwsZ5yw
WNLZduBukJORP6R1dwW9jUn6iN0kqUF06tefbfYB6lgllnvAyYF2ls7MtKg+4DDQ5/uONyKGYvzV
S3ObHLxBr02XiyR681MNwbUkVmMNBiZ+NWfBQiqhZPVCPuQtjS6HYn/tVn0/OHbU51ON9MxJGlno
QIn/KotogeRCGs1dQFiPw1zyD40fxZ1olRR2gJxmmQQyAI7NvWKknvJXkh26nSLs5KEau58kPUEX
tylOyVvUzttWn9zDioC7Csui/JoCNoFeASi7/Ogh8Z/FHO9o0WPzmtkPEurMttpuy3Cz0t4cGeFU
oieTEBn1IirMXSwuwd9PQX2aWCdi/bfTDQu1Z+KH5ASbkxuNoFknz2k6katKhnOqJ5BxoEb2fJRw
1/iaD+5VgkTFhV3sy7SW4pVrLUwxxatWMxMoO1KwbpkmWCvGzpnQRHduMGmdgyaccc/4DnqRTe9W
OHaz9dTv0NZ6KQ4Op27WB9iXIgDJ0eQTAupClJUuKXVyjE/HB0e14ctZDUBQOWw16Pjvq+bJB7PW
2FvnJ+zaIPOiwok1T7eZ8ViUGauBzwfanCKxPUaJpLJB0jmKiW9SwXaypNAuhXXxZqD9GnRQrtPq
bthcsblfQj1nlyUGslEhACwFZ0UuL7FUSE1+sLRPkEFxvEn8SmPx3BwkLvf+sXzGQD3Gb8zTbfZg
yy6MxQN7p63N8y1d9xVkg6F9wGenPiv/VfwoU1eeQo7MDWbwRMXDKbWWhfuXrnNrAdhQFxwuizro
6ERB+Hd1dWa3RW/aAk5Ubll1NXsV/VgMk1QskXQvo2sd283JOsxsvWEmzVpZnoO6dhJ8R8RCHcMa
6cUpnyfrfVHTchi531lP3P1cZjzdA8k/38XxkCqhHfeLDlBC8olEntQQIItO9zaIrjK4kM21WgIf
FxtuNZHirZiK1GWM3Ut+aA90qWfw1JbC1YlyetKny72mkZBhyJdGnoFc4nWP5Xy/Ia0fB8AcdMAA
1hAWUe2PwEpL0WtGT8y+qWoUSd2mvdV67+LOb5/J8QuVGstwiI25ePI3+VWYd9BGxasFXK3wFzeL
RRNROUavSDn3Mc75SacZpdkJNv/5FVPcrNFRdU8nSwf0GAPyUIGc2D9w3jVSaNl+gZ30uiFzF7L+
3ahnwQhaHvMRrenLkdVmyFwSPivTGtE33CZqzn6P7/s4A6ZVC63icvdFZnaaTLY/3GYvSqY1LGxf
P2TQPVAUa1dfM7B/VpXnwAUHKHadokvSO/y5rVOdilmwWO06OKo1Ewq9VDVTgUfySyzZAgBKbrgB
iBBem3y81XdVz/Z9JQ1tNb1g7JdEe5xPjhrJ+otEzFGAbNqa/UYubJC7bBCXn1thHrVnrVrjVMia
L1kSi+hJRdWS+vLmeTkMf1BzwDVt8mwktImEjsRM9NCtROfmooCgp+rKdyR3A9ZO83FjbXk4ye0M
LYo6QalzYz9bniDTyODXBAxzPRoqVl9Vvp/DFARfd3Lb/AyvxM9MJdRGvaidknLM3gl7TJ+ExXAP
9VVNZEhfhHRMsuyzwvU19b/fhporu6oLH9BZgq2QXRO18LsATkBB9+EJDUMA++jufVwbRLXfaPDi
9zBzOyiM4DNkZFaNKWhdtBUv4RvpCkZU5rnKR0xKdgDLo21Fuv/lsYVQ9//qHE8TUvcLSfleoPwr
nToMylLS13Cb2+Nk+LU6WvWiWB5mThw6mMbAVF0wnOyxljfBUtvSxdcKYptkRds1SEgG0kULU5uD
XRYmaNYs+O7ZwZ8LvKHJM/quo4pyd4rdiSUhXaSvZ2e4saVX35vbcVqXTroibwcUSxTxkyvN91lr
UJk5T0xv7faQZYUoFYbETBn7UhKHqiVkHNVXZQT3ita3mTKjyu33Bo7hMNYsgen98EPNUVYxmATr
Hqtw8P9djkgQF7pZGoTqQh1QBDtONCfG0F/wcymuFQG6Sre+0Kr/Czp+s5Zj3XJxrtPNAwNHIVMn
2BLHnbNtDvKyto3AXnnYdSgDAvsb8HiuB493sTGJIziVWpbAgbJm22M8oP8EJ3+TohDVJY9u3O7q
1g9Y
`protect end_protected

