

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
jPOKnt2dHOagW4dFov86UptHPGMdrE6d2ZgqMnfJehhzqeTiVLl89did3kf45SSrRMnQy9YGjxY6
jqpfslmzag==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
TbXlwhQ0d0UG8+CBDSNOnRgRBfh1oNNVi5QwoMGV3zJAlkTsnTywwNiy3IArHTxG6Niq+d59upyT
QOuldsHqtyc6KQBpxueCYJG7Fv1OIOGGq8mGjrkLmbJVhJEwBvPv4mlhsXKQ+/UhmQDpF2ZyKhkK
EbgpRIm7ap2EmEdPduA=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
iaTK7nKuH82rPJSrGYALVeHLyxEbb+9Rh0wJiyQuCqzY3/f+ne/dT7ytF39Hm0BXD9csWKwQp3QC
vOqzo1FyLi+w9Ik3lkb4njvMdZauHueYbVoku659dslyFGV84Aivwjcg0Y5de7FqsEonjWrVPTE4
0oo4m4QHuK8VN0pa+LmuzTIHDEzIPM6IMp8H0IstAk4VaGHg6wlCrG0u2kbbhcyaOKk2xzxiDfSu
gcUy11TT1zHFME/fHUU4VO3aHMSGacP3N+kgMah6x7bBUjBd2rfEXkVcl+/1g+qp0xW2BzItYrMY
Q1wtoE+N2GipiyxU+AmrXQ4zQNqO11zaj/N6Ig==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
QkbQ08NIPb90+bNjwXDlVNk6WbvhfydYhJZqryulAczmjZMBvdwitIPmanwzKj9BPStsPNHXyOKf
9PFA9l/uvQOwVNRTz3G2U0+6+YFy3j+qj97mRopffETTpncxm/BoroKpRNN1DrgSjygcTkfrt06N
1lOXW+551KWRUPA+fGE=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
LXGnS/C7HF/SjGcWlSWMUKmilNZr5UhJNWaaWr/ybus0u0ctzmNkXcydCyfmEQe8OngFPF/IKSaG
XMrlZODcxs6BdW6TBJGvkBlKfbvIYg7iCmAit8JvgZpuYsROJrZ/IapJ9XCUZT5PW0Y/S/PoGs0O
fXalNP4hoIYlP5OYjMaSowkFFmCMq49fHUdBBmi6thqlMFhrdpbAhfGoJVYkjStWry+O4YcFvpKw
Q8WXsOAh5J64eppUG0x86EZ8HpsK6EGAeT39tAy+jNSSIcnklat3mhXxMF+BE67OS/DRt5H346yK
YrLlKC5qbVgH7HjzWMBFYeVVtUec0iic45xLPw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 11232)
`protect data_block
AFeK8fqX2SnD2KqUMlJJ28Rki0jeS2n7Wzkuf0IAzEai8HxzQEitqT4Smw8JcpwuTyZVRELrtBN6
cHH90IZi3mP5/TftQ5DJJJbn2G050GjNvY3tohuBo9ruo2TsZu5EMZzl14XqciD3JqeZa9XZ6zCC
qtyk3IWua+GDaeVXtLaB3TTXwqFqbPlGE2OF2alA4BLDOaE6eN1mczRI4VDZHaJYiMUOCygoH5i4
6MysAmHHHvn8QB+wuGAlJRLfpKhCIK8oDdD+Peo4/uc76W3hHbRck11rVXM4p4KZUJIlHcI0gnZZ
yg874gM3sHN/bAbgs03J8w22pQE3zZy/N+0Dn+gcwcD0HqSWlmk/2qdZul1VNtnbVMt/5PC8Wq7Y
LU2kwZ8rhRudeFN63Rxg1KlLDjgj/OsXF83uYNqKYEz6yFPd01SDe943FUULs+POpsFLBqMDyPRW
QhmPnGRURytikeoOFAr+AB2buN7sW4oHXLVqFX8oyyRlL7j5wLy1n07w+NBznWSQtXyDtsYVEjmi
Bme2EVGZiybOKd9FAGHEH/JqvJ4f15ZExoqYNCJ7mTVKPTaw45zMs5cxQwFdsozBw4sKRstrd4lZ
2AObLw5Jg68Qg5ZohZgll72bQGqzF70woRe//oxncWm3fjjwjaIMKJ33kmRmOJ+JoErGLvgqLhSX
3KQKZ6/XxuMVlvG+dRCQX2oSmIaHFkCkAg/HvVLllscYUf/1gIygYbm7fpAjGYI00jfj5pfCf3E2
769VNg9wYfZjeINqijJacSyvxIpRj4FqHJr4cpw8+zY6mkhc2L1aBZ1E6f+jDTfLpUj98Oqjv1nY
1sMuma9S1RVF9b9dt8paf7JZXaNw1pYNKOo6b9N3E01lpjivshAt+9Pina2Pd4dunM7PD8XQFiF7
aeIxjNPyHKdBNI8Ny3eua/pJlbd9qQyHEYOkiRsVtEAvZiU7A/Gs5dVCWAJcmQoWGuw51CcOmJ+S
4HKzGwUspv5XZc3iWJNlwCOwTmEVxvvjRVCS+bbbrzEdt/bCIvaP2wwma4SDFnWKu/BZMv6nfxYX
vGHluhGdHn540Fa7dfVZ/Lj1O1zHeqPJqSbpVgWKXGy7jj4hyp+SD/NHiNmoZmwxDtE6UU5YFrnD
wRnDjPbrhM1fvLPkrKBYhu6j7Dtgx9exIjcgWQ1/bsuB4wgE7h/nLe1+W9ENV6WLGt8fuILvSxqg
nVO7PqdqJ63yIpXH+TlixXPTvvolDK4OrWrYHpkfyIxu0OrU+1nK+mjwLqYwjSHlOHAbKCkCqmXP
s9RYDp6KBb9rkz+SOgFDyr/GF4jVwtdVJBKeCEcUul6Zcy2R6cUNhNhcXWeKDd7KiyU3PUbKtWIE
CKDzOgNCfY04WhhR+qhXWidxDkyGEiATMVzcK4u0+OtQvlMcH9Gvsnai/ZRew0XkIkW+7zWe8N2u
9doTYzE+Bb6hPQuoAygxBfGbyuimbsWN5Z/rwUbrmmlWtQnhgWRoUi6fnQFTRXOFkeRE1bB4LOA1
AKjqynk/rssmT1cdL9alegQAg9JVcRD9DHIrLCcllu+1sPu+hie7zpUaI6QAjgjIJxasLHpr23yj
dJ1JEcozucKegKMQoD0jP61czLpIQKfJvbhrDT6mvVqjisE3odJkMMZGXz+tFgkrk/ibflUVrOIK
aFpveX/ognQiJncubl0rfEM+NmA7gF3lAoW+pbLWGABp+s+IZNvUzjCwnTsMPICNw69WOjrGFJ3Y
MTDbnd+YiERmmWJU1Dctc0JbZEmbwEFHN3vqyasG4ShbPZCXTe0JX3ipOL+nD+mNMG5lF6UqolCz
riq22S83ybgiB0M6bNbiQ3C9yUJ+Kbo4WMlA+Fkv3DKi/NUI1yOk2L4K0x05pxf6HSGiqco4z8R8
7J9eLz9HSr+Zw2juhJYIneg32/oSqYiLKXXdqTUEB58qVIG7KhLETggNoq8ibdTv5lCwODBElbRt
ZQComBgTky+4FFCUa+wzurd87TYpUbPcEoYy05zT5yerYvSnD58HJGSn3vKbe2ELWWiuYQpgjaf8
4pQ24pvnZck6CtFmVTpJ7BubFD6NunQYIb3VjH8LSuTKolbohYPaDohLmrKAJ//0uRt2yda9XpP4
zcf2U6herJM+B24KsIdLVoKeXoWg0oA4iJOqfv6wnnEVdzSPFx5Ps7vshCenauE9RjQIR2uwYfCO
2uMlSPiJEZwc+9lPtSbrZxgXWQxCCbrQMm4zYtf7rry51xnIjr17c7XnzJRI8/ig3n2Fvs7fGcnU
9k82D2NybwyIdKQ2oK0ZUV6vUpvwJk4wIe3eQlFoVd90GeVi4qDISk/ZSG/XcISi0/cUy9dmone3
1yKEmSxW9izyNQG2/DdBTlY4IjpFguYdT/ifRVi3wBsigRgPCduoR+9cEM6pRsHaFiYV17LfvV9K
Le2rdwfeHDcgWpT5Dod5N3ifTuawDr/1mGqqVBgngy9JuVIfPn/fTpxj1rpeh8ZlBBuXZsXZ3IN5
sFsxahkwIDnonEdWWsrO1lilGHQrZ2olO5r0wDyHh96q9oL61qmByjgk3wo7EHsBWGPWYZMp6h09
xyOpPCKYt5ueGYP7APkbwRLKmNB/lF3oLSzFZ1khGB1e9d3UcdHas4CaMsHoRoIJUbGqrZJOH/Dj
PrN4NLZFh+Py6lUoRQ6SWoRHi2uiA4bLHFP+PqMM2hDAC8UtoY0AdDZJe9p4J8TSf7xsqvZ6V/UF
jIaZLrfiss5xRimH5uzrucUhScNH/gK3PcTbH1zP1YOgAlt7g/ZS+bPQP9naJRndCPEGmgCLRZVB
VrE5q8slsIV07dt5DRaQzQfV90MHxkUyHBiBVGYzED4Z9Bmzj8VAa7chkEO7Cubu56d0lXKGiaOC
g2mJAZ9uoakxshfuDRVc8i65/nEMWps9ZMh3yiUYCK5clObxLarlze6SU6aSbuEJWfK7nmGESZQM
0f8vpJhkVTNcu/AzytZE7EUKDZ0XB6+ix/PBeejxeB0A3BRqDcVBJwPh7QhyvpuAmJ0eA0YCvQLu
wdU0o05EyE90BT8XbE66KN+f8zDGc49CjfhRgZP6O1LBaM0kkwqigmg0fb3zOZmH8clmOZE1Br1C
7Ag0tcehrdKu0rFbuO/NGQsLna5dTxMAgNiCWd9MHztIja0GlNF3URd1r0cIuOvr6nblgy98Y1ze
avaDUrAk9C529RALfLjoWqLcebdRnS7LEt+sQPIm/gMr4LnV+O7IhuIWJ6TPbhUI0ucyce/rdOtB
hKiEj3ZlbTuiptc1yFhNcEROWFYx0aeoMP61k0/6EvznmefkPhLd6MDiZRHZtwlfV8FPfLVofO5S
iDMt0VPS+/mlcUQV+CeP/ZbaY+uRpr1adTVpWDAtIM+EXLnxX5uJfZGlnsJ1AorKnCbALw49GvTy
04wpKQbhljMV/0FKT3rMG77RaNej4MslIPidAEacbMVN4jU+FLZ8N55y+uZy0TvbTzkc6JFKW32T
y0rRiIdGNQSyFnHlt4Oa5Vto11ln/gFN876ZoA7a6UonFgOaeJK3HQbWNAPFr0Y47KGb1EAKPLWO
eSvgjTtEpoaTGnmwWArDWd6x+SlPuJ29Xu2ujjU7q6N1KqmElRSYZIz4ZbNGB599UnytLz7WdADz
Mgu0B+I3+GloKdxG1jOdYckA0+348JvvvHBDZi5vKChFvkfoAZv+LYjTtm2DqhjpPDAtvpCOY1Xf
Ld/w0ki1zeN9Ljwa3zxdYAgiKMbMPfkt/NWfgTDs1D1dmKxsCJeynod1GyXceTzRi3NL4kkMDRLG
PWIgRpR10+J6+biqfyGM8/WRLCyzTQjeZX9Dy+Qewnmf5J7dxCQfg83ApS85vrEwwApDvkx7jX6D
NHizoJ3bGmKccQwHFm0+g2HoAx9v0iRSggyQHex54bQWUIGawuU+Lugd8exjREEf/53tvxwRWq3P
+j1AHYZX+EGkF5113JMyeWh6e5GfjI2bVTX3WDWiqEOErwOU3ZWMWyGvokj2bS5zE9X2KJviWJxT
QCMUQvdQdZEgJDaYDrwhhR1/IDDUqJW1QfrUC1J+2lMfgxJ+xONnkvKKawTtxuTf5d/8SNd171lC
QclPR0mY+j++A2/JYjnFvigJGN1RafOAcesT7i2ZXp2GVgcGPuWOetl0TbSilxjPu0z+4xL3S10w
r9b5PzCIIZaYRRaYtSonVPlLR4hT6CJoe5YLnQzHugXvZ+QzYWb6n7GcPnPM8ZBZQmj0OZz5oToa
HzJu9BvgKo/p2hbBozb4t52lSe/PRNe3BAy+wdkxwpw23qeVeI3Ng+nvclVfLvrAabXP/dh1yJoU
kf7i/OfTXK1Ov0f6UxNnj8RFI2luABIZ9f1FHZaQY0pGwxg42BsK54uclc/Kb1EMXHJfMz8s+7Jj
038rbwRAOkkM+gjnP3dtK0Pb4LE39RZnppzfovyR6fbcB18obe+CjtWOU55/6OCiV8KJSf7gE6rx
LmchWYWLLHgK6tqSYN6Mt7Vl65zW3r12L68TN02vxc3qiP39CfoTFm8w3/CrjUt8Vzv0K/LptZUF
REMgxzKMvB5x4L7P3hJaxNjS2jdRGZu5GIqnm5f8/pCl1Q3dGG+OIdMZL6OkUBe2m2vnc3oOxo60
X5O5pEr2/gGAk4dii26T4AWvVSkLA4K3N+Q4dfYffLWN+Uq+6hM6KG67FPaWxm7xnMItWboTMr+b
8TqD+gi43zwKxyEaf9rjAo8Z4Ha7F0CreSu35gPFpoSec5+BaJLhc/AakEoOdeMW/oTCMBL1tn35
RH0o83dnrkIt7GR8myrqJgxvPuw4nIRlkr5lWp4qpisGnwWFpdHcS+I/M0h0sv6hcgLri5uwm6Is
yKCoaCZlitc0GTJZRqX6UOSOi164cIPlRtDZ7KlHe7HVjhCw1MBAieIy/Kbqgkph4MiO0C5U1rjH
dtD5J22PQ4ih93xP5K1/LClRES8ym2Fhepj/MH6CnCCeXeEBH47L0sHerjoyo97KyTt7EWpTQ2TJ
6tsoEmNUo4e3NlooNMBFvsz4q5HrVDd92J66aAkzHzOB1ZUHc1fQzNlRhMEpUI+xvjoalJcW+3Pi
eIe/gw6qQt9QCKwO7xh75ZI1nBvfwW/bct5E9Z1kKmk4x44XMdBLUOp2VP6ydVwE4e93eEtv/gZ4
yeoonZ4Y0QT0T0jaDap5NuAQJSS45GzKeX/VVRaFcaoJYzE4b3CRAujtl26GvKhbS+C7mEjzUlxj
xnlkAqOCXfyk/3bQP7Q8SuXaMrrzCZ+hEDoLDN3BXr/yh1/EFU7yBTpeqLekoXCvdNYZPi6co2SR
S5z9G3cUTt2em++nhF4xcvpL95A4bhRxZIv65ocOfC8rExU9Hm2qb2b8kEj4d/IV+Iys/FmYk/W7
SZ4Zb9sUsxekOveD4Pfd98QpcDwTAQTUfLUnE27MRPiTXsqAFNkyrPjTH8BVosz00ih9A7k1aKst
k5/lL6C+ZZQ7oMSWKfVMdsvkIpauIWcIq0+xASkbbW1fQ4lWxkLXddvS5Xr43tGZAcspKwF6i+nS
/oj4UdommSy6sqqm8qWz01y4ti21/gqwthInBnQiJCei8xTg3TAlNCIvPg/2s7u2z3GCmD5tP5c5
OcNpmeE0tMssHBE4/0R9TqUOiN+8YIbfM6DVsRRF+ytY33Zuhcis8imHTKzfRgIGI0cqR6mDt5jq
nsC+QueaJdzZYvsALYNy05vNpkxWxOMCrS0CxtoincWnnJT9BDkA13QsEchuyt03aFQCU2wJSTtR
y4i4+E+0UoL8CRuVBKN9t4ZkKuU4W6DrRNoOpaxAU6hRod7uDtrxXSJSbsvdzjLiRYjawjIDLtve
zM7+4Hz9t8Y7bn035yGT+LigDyDQ5Xs0ex8AayRrBpWgxBGADjwne6p3gRq4a1L6QcwYTsQthruF
qtaPZhmete8mQ3/Ykm2nijNBoZGSYbD69EHP/j80laM8gSRF/lbZ16q4kuOTj23yT8LO8LBdroh+
JI8+w54+1lAz/aCXXjc9YM/OR1m/yh4FGvKeFJDuZVQItHQOPcaOIYuSwVTYsFuUlp9SMAN/+9T4
CB6YiBTP0hwTx48IWEKCCV/bGegv01avf2vyNRI3eN++agteVl0zpL9QAugW89j6MN751L5EBKq8
t8/bfvYoYlcDE1ElkU2mY3ml2JVK4KUaZABVe0YPwKqWeBDA0gNxEm6rwprgFscK2v6c0gohMu/X
uSdFooXBMziCYjNhm2vPksv7Ias9GKT/jouVr6+NjKAAgI8czKsccY7POOKY4ka+WPC6G1VSRrUB
XEj688H3vCWv/6c5jcDdf8Aogw45oHnLbOJOkHJFM7MCasAS2CkfyzSfftQLvdU2UdhesUFlBUI9
Uz/KWaOL+TGb8Oh91U5b2ddJeBDMjbeJ/C4Y7rGomlcFFcdk07W+YGiYTa8ac0Ynbal7kNlETKM/
FBTf9gggNRm7VgoRFPaJcObTO/6JnhxH8PH1YQXyR1r8jkTR/oIDW6wrFQjRJCjNs8d/e69sx9r6
hrRdzvpTmgS9JkKFeUDT2DgyNZZf8mrKFlM6SbUFB2nD9IDnFFrcKzIt4qo/qCIbUnsv8c+RHBRV
iXOP+Cms+FdlcZEY91ZnBmpCE3/Yy2TAuzbg4b7BF4XlKlD7SB5A8i8sxq9YKjffU8O1ylkcOgn3
1ZDY2o1rSX0KPIjO6r6IawMZGM7j5vupJso0ZT3K9BWnZCbdZ1aQNtWoyI9/m3wJm1twca40v6yD
6KykSgVAE9ucLf8zBNXxpsrwwJbLB0i1rjyvXKrfOAfz7rkBolinggqpNEqhk7Sm7lS5e1M02aVG
fnNcjwKezBced3x9w8aSdXa3VZPr2h53FcsXSjC4rObqHowl9W9UM2y6+BYtYPLlcwK9nom7ee69
I6RVXPk+L9RPnhES3k2Ep3HIsF7qwYEtUuYj4uj5wmx+/rdO0cqwJzUywcZXAydPsem/nG8bcPG6
caAQNNcnrVvMlo0KsmEsHASLue8fntmnapUdXCtX/8SAjDam/3mg4rmvf/HdVyC1+myhZhk1bjjI
6Vu+xCtCjDPaVhR2hP2q3FfDXLhnZpRMGqs+xEzo2eq5BHEM8Q3zAmeP4RxJZH5fy4/nh0dHsQIb
scFfY/uxJaHvMeu/ockkYvPTFChrFEPgmFG2Pi8aBJ8PIrXkF2Lx4RjU1T0j+RH57opZgV/Oqy2o
47HUCI7BedSrJhhTudLVmUQXKpiluNchLtCv+xcwVB6+aeZ30XNusYT97ldPZfiKBrbkei9TENKy
yew5xXtlXAVej4hurdaKq3lbvRTD+h6smN5J99SMGnpwZu1PUTN8IRnzGrY51Fu0LiahTbwXpjzO
NWkt/tIwUhkXiAe7l+wDKvX78qu/983ADQ59cHQf6Khzizx3a/KIeW9Cca6q7M6Lxn2qEj7mUjim
mxnGgCxnbL9WGdU3hSEvLpLpd0yInHLyj0CEz82/Uz6VGKsDLHpdFYjscz0KP/wZ1hJMDhKcnLY5
6scPQv6T7Za+KiH6UdkgHCdy/l6HnV0H7apc/TBZg2/evUIT0oHVsJ6U6aYQTPbtdjqEelXBLWF3
BN7QURbh3lNQ6pFgmzDB9vCHlIuaVcuVxshUJlBsG1wRqb2vSdn9ra5oSsUE4+2NWBWB7Fz+Gt6u
NZ47HKDAGj8CmkeLO9eWrXanZGFceGA07lPWdiIwsc/m3klFw/nkGW+ZT8rgVEx6NMRufxW1dNo9
X9gjnh8RHqM2qwKOqZqda90siqRXigzDeypPEwJnpD9D4gPs1CUYeM1/XHwjFHCo/PM5OYYmk+UV
KWEaH9hUoCXuJydeA4TA1fSyGugijzh6ag8opp4vS/ai1IWYQoOesFHXaaEfwYG74B1OdUAXjsP7
DJwR8xSidSw7nfMiO4dDLKc4WY7GkYePJYdAtL1WYYZdKBejaL3vUkLnNhaEPvGF99n/EAabf2Ym
BBlnrT5Ww95nzGG23I9hNri4FP2EKxwKQllknL7qpn54rL7N/1DtnLaPecnQCPnpBStNgj7GkXXj
MDi3snEDCZrUZIfRogTwboBwjAafggfR17rsWQbcfOGufnsysEwQw5dmNKgRbwuZ4h6ErT6P8PBD
Ja5y2dKbjnVzVS/XNcIVfAPV2oXBRQS6hFNG90P7m3ugOrEbReqod2mHAoJbiD9ITNQSDHWvL+pn
mM2GlQSph3hUs9U5xrEz0wGcEGlRBCS6HjH97AqoVewhI6hHAntnmqwgANYafgxQ0Wlds8odY39/
66wEp9TLE87DJKHqPqXCMJ9V9/1iwUfL/ZzSLjvRhlETQfZTkW+ZFzFrNYj74PM70Nmko3YFiqmY
V3BzqFfrL1XbESbq/PUCIUCpRpVua/5/iBPZzP+TUsPWtErBMUb3Vu/tQJwDgtWz13iU/dEJLNz7
C5iPVrQTv4s79uzkqqO8nK0XnOjVbMoxmDREeQ0oYl6NBTbsqXxeNnZnkfE5WySofSyOO8v7z21X
IuiZQ1aPgCuctoy8bHL0Aq7evwEkbYcbZtFCEutnEX2uuZBOpYPIU/NpvumchzNV1IxKxxnh/KFH
B17ZKiEqyMmy4C13HUUW4rzpSy98JE12JYZ/TH3PENiKBRl+Zc7ugkk5mAIXOG63mqXUYlVi0xUQ
WM+dMOFzCfChtmFlktgaHzzX6URwvGgA2C18s3v1H3HKmx0mWi/e188wkTA0oN4rkJT1H0lvU7V8
DPEhm+jhU8hTfzpdNwnpt8avAaQU+5JVMqNu03aJyNxeFGWIzjvcwHc8PIfeJ3Z+RWUlZTNNYWpp
xLC7Us4vO8rHeqlNKi1vW2wbOWBomjAW3VJqouyyk8Qdnqj7U9y6SvM/mYrFebwTnYwh83kdeoZD
uR/6RMdPzrt+ntJXZeKhdoTjbZFxz4kBgTZkDM9uRnjLlnI1FL5PGmldhWmIpi1YU8pXfFMnHbvi
bWCRuRr1Ly3QkrFJRbUttArQSLHfcDAHQgWmMMon0+w9rNlO+n7KX8YhE84nPLkX4FUfXDRM7rve
lWD82nzrFDA+Ew5PgPceB+2DEf4Ir3MUSO7KDojNDsRMa2BcjsauwlhN1ZMGu+VvaVHIC98ZsWdK
B4QENhCli+1zT5x0A6gj1d1tII2Y5OLMYDQ9hCY1vwEAbOdhbzsPYeiTvRsXPquKCu9txF+rFWjr
h0osbhLissEbsiVSQtUwUbPK3os/qUPlTRv4m0elhpgDkUYtI37oBqauWNcw54c/HGkvSHJiQ/8Z
12g6LzBE8JOultikGQ+rZ/vsMHecJq5t5hQ/cx0d/u9SvCAlQyZPC9HHeRHfuAHqpNjzAHxg+7rT
F7Dk8FlhRU3zRtmEjrLgv7bruEGHaWDmV4VAM380K1PzmNoMIkWCl0y1nE0FUp1eIPV8Mk4nKj8G
0lZ+4BGx6Nls0nTpmHICZRKSWQnTX2Ioly9CbjtOnoJR30Q49KG4E/mVuLZlF2mwZG5qouRHns6P
Q/OvYlGkPx9YTake0Jy0inHN1ZwQGufdxOtoZu+SN10bWPyhJ4TtjXhdwAlWolSF0sWLP7IY3VAe
ZSxdB9AdjJohMSrJaY10Sklx4YsFwo6WMO134H1ID24Go3U56HqwhwInx7XwJaEn9anj4l7u3dwR
PMJgIVme1FNquv6DfSmGi7J2RNTR0FmTqbgELllTzqSGfT2RG8St/oayrPBChmd1z9CqwYp/MhXM
bDOi65SpP8KFHmcwsVI2aScf8XwzWaHM1VpMTrkwy9rFOnAt8H9plwvwuhwMT8b+4Vuy+FSmSIgU
pY1wAnUHaScjfjyMzhNCIx1X8AWFB7dTOoenFUoOYQlA6AV23IOBulguKjaw2GN4ZKztO/3H9nfg
rbG8fpGj+5XmltZIgV4HepHoTjpL9HDr9w9jt/LQUCVOnn60kKiKhI9HrDFNKxaCZLNVddd7WJVS
STDho2rQ8oSiR/7T3/4DDozNSDPa1R9qIEDSDK25eWptC7QVYf1pbgqzwZr6FgJPhS7+J35nIsNh
i2N2hjqlmZsCZhppKY4mUd/hFDK1ybPVICnjSdANTL90xDiA6eVWtslfQgqGyYKklM7yeQr/G2vM
uSX3rhVWbI+nku9FwJgvcjmxILkqjUsCmQnW8LTtm/oLwbWesXHm0dMdISpksZ42zRuRIeQIbIhW
t4pIi4JxFcN1seyQQZz7AMpLXDO008zOWkpvhDihXGiZITawdByScsM9b9C9QAs7V/L3psPuHmCK
bRLVcRltiRxftFH4YcqpSORuq3+3OGoyTeOz0X+q8hkbRYxepKZvyz1cY8M+1mEJ6NiH0sbzqu2b
4igwrsWaHNETHv5pYMJdJN74uuU78kouClbf7e4wVbVdeBA8dTJjd9BoajXHge5XzdgIHDKy/WsK
+9HIuQl32dH1ZPMdnxIxeOfeJoxncMcLIKXaOeD50f+QE9a7+3WvMrJodK5LG52iLcFNynD+e+z3
NPECX6gmUynY0aB7gZ6RizmdRBOD1GA+WLN4/CjLZ2kVBnNB+QvNAMHMbp0oupjc90Wlkbg1fEvY
q7Glc9l0mBX+Wn0OjwrIgs/n6PCTwYfH77rPOMtQIOrXZW6EmUcXoqnT1Yksne7AR74Czc769Z4h
asILyDnZC7gDBVqgn08plotaESPGeXlSTc91hc+fdcB9JS2KGd3EzRLgEc8S+vrKAx3VrmKkbkGT
oaS3zD7VuCBJbiRXkf0CTOyHwghCwjh/nSyKtY1JzL3He2agpkJ35VU1eydlYtDzKRnD8mfGG4Mc
Jd8CcCj6Gdq+OLWiusYxvqQ06nra3MZzcacuxVhY8CBkov5uumL9XLzvGZk6tcNnsn4N3dt9HLSa
HwD8ZyW6xhA0DPyj7S+Pq8sOrCLVcm5XoDJs2i7sVl2v9YA68AeeThpsmH/P9JcAFMkA32Y+2Dvm
S+dhxL65ybmoxSJRCZhv2T3A8CqwChP1yq203vSSBYREW3JUq/dLjB+ut8FrKLlfB7NoWJwf+2B5
QkkGxdYoS66KuC2NgRU0HYhJSwP9pcmYEybPMW4VmnNoTyGmeIQkqKqybCuUsSczv2bx23SNjlp5
RUo4XC1tT5RHqXY5cv8YAdoO3SJWShZXuk78g+3XIN22wJoJkPQCYKfRgTq2PcRHmw0sC/8pBOZZ
QYAEhSLq3SeOi9gEHfLwew2FFsDBU+bTIy6983Iu5+cGT8UK3kpfAeCUVZCpc7Wq/iBQLdJtnyeO
PYRRw0KiQ01sDmp6ZQwb3+Z9bckj/bRMsKykujzd3e9POloNRA93vjDpqhr7cX7DtHsHyOC8G+19
2LVHMRUn49UD9qnvFDV43toToRyk6vYULHmgaVkuhiu6XYq93ctk/g5cgE1XsOWXt4jSMOqwdwNk
TnZS+3h5mTOPd7vmCfVeACfiokiHMrDs8yWzs2lhr0VCk8WRNb87bhIy8djuZejNe9wtfccMMzGA
QXH2EOjEpDt0F2S05d9O7qWTWctW4r7cNpYYKa3CQPRNSDK2N8bl3owh7UBtnt6KME6G1AiMVfd+
NpR0QR2N6k4S09dT5f5192GJ7CHEVFGp3s5aZpAS1Wqk3JNUTFu4RKEdGOF9yOlWhkIqNhGxaIIJ
yrbTjfFmG72tVMKOYq5SWMHeoK8xeHB7X1RUzmXX6t4Jlr1EGFyxauCSdrzXLC4OJzOBbl2lWwx/
/ZFr/sOXYv07mZt8Wx8XNDARZQ+4YtPyzSP3iocYx5IGyRE/xPlrZ7pZ2DUoExs7zt6GgUjU25Zc
NpQ4vQuApvv4aI82ayTwK+wJWEZ/3sOitc3Tf6+CXQ50KBPrKmOGZkc2R9sbHVtf9Y2tROS2oc/X
7PnYXp+PmUe6MZexSZsTrBJzDWDDkziWjFHgTG7rpj7JaydxMXIaifRoQZTjlFldnuapBDijmfUr
KiRw+Wi9U8tZC06royUOl0LLKNSS3uqe127hRF5fBwzR5bOOitsOepSnmtnFPC0NkTF5X76f/bA1
w8+gjfb019D2o3O4WeSMv0yqjP+VrwmXxdBO7CvBC/VkciihK7yPRQtDSbP7Lzi9W43J+eQ05AAs
ozSnx+MiOzUATeivN0det5i05fdw13WtFOyfxmX2oJ+CxsVwI/VrCMWXpqJoH4aqOIdWEteAZvQD
PqBW5coSWAkAuutu4Ms71UsQG6gwktAlkvVltfYhkqI7sNyQs9vQDGSLCfXfqvN4d6GCoOdkk8Tv
WgED1DdiwLVVIzToXLawgPEXs10xD5eP+EAn5SAkFweXjKCRpdwQ3fZM8rYoXuXDlicEq+sznk5U
oddSqntU5RVZGII4LJHE69SbrluRFoZ6WBZndTy4oEx4JO9+vQCE9pSdMNNbWfeYkbuRErBFHJNp
lQ8ICYFH4JsGxWFfjkm4qvURwbIPjUHVDdz5BtFYJqEEhNUQK1BeARVj34RAEKf30J07XERqqx0c
Sr0AtT/KtA0XUMCsb1z3lNNurP5dDaVixAacI7O7f0Fow2ixj4k0YBogbx5xvaQXIQimWZvcAmex
6BSo/jIilToOEHdAInytOGs4Ck3q4gdQzKrwc2HBkqQ7XTItC90rObdhSqtiPQUTLtu/nA7M2MsP
GR/9K3J5CQNbcudZpSbVYjEzCoLXdjQ5ctx70RgTsmwEHrwiUTXY4AgrfgYr+CVmgNF0oB1FFRC3
3AhZCeqVbtTRkZR5/f/IVTkDDkSGWf0Hzqa7uDNiwlNljmq1rg8gcCTZYwoqAWkK3iREF6nbOhcc
2FIO9EaPBwW6pZrGbnkF+Z3XIy8VDmkZ3jUJcA78pA4HkV13f9mem50lbPChyOrW14CSYiRQa4Ja
BssBcs5oKb9Hl7QmdQ0e8O55TyR5/Y3RYWjKGlAAeeEZdtkqK3mc6TTz3u+zzm+2fVrHwmOyiOt8
135lKLoi8k/OLDDLmuaBaLBgiPKPunl/hkQQ0b5XXHwm5afPIpQQHnOGCY3CBlARBXeJI8UYYJmh
qFTDiL6UXAhmfSOvkSX9zRxFrBuRe+Yfb7e6G7ZjbAZxAmsORMVHZ1EzfSX+koh5rzvE6Ix+mKd2
F3c2NLWORm20cl9BaPQjMlG5eW0uYMLhTfHzqMYK1vL+jfutOWC/wd0gELOp9/L0DxIFUSGY4mJi
R1uxeayySvXwRmfMiVU0GfDyPEC4mVAIH5nIGsKv7jB/jf+wwaQX65I+X27hN/rJM5P1+zhcjHtO
HxtU7GyCqaE3SFObh+ZjnlGXGtssOFm2N8NndyCVIxpF8ewxRrCeI5jn4ZSI82xnRc4vx/E7d70J
aFKPxq++7AtPW0gWG+rCgeAf8t/219RehmYLGhTMiR+P5o8cBLzoKlIrOyNCyglwbYCys0Wy0+m8
+jpBvt2QguNvhVZfTTY8A68bNI04R3e3XD97WeE1z9Ruc+MHFzSdAqgQCi3Dxtiy3Lvs2WnZ+PDj
fTX3mNWA8jTUHW6jnuy32k9svAF5nU4VVms7mBD8bwnKj2HP6qGJerjtPxsEiePJhTm0HNY7SsJL
RTEXVpHljt1me/4P+es3rFrJHsDju6n+saSHQTN5ZrfWWBOKa6uXYpKvZ4dIiuxVYJpTsQ8wGujl
8ljTuNWrzNUsXLL+b65aUFy6AyAmDag7frk7nSWPusRgsZXLDYWF5tqeRLWnlzTXdu8xw56ySGmo
hUX9VU1+hdP9FE1uPcmxiDA/rEU/bExsgPnui0+0qfWgoHZMtvXQG2CNUVzuNvQ/82blfJFcTxCk
19HUJyu7r224YQ/m43Ze9wy4J0viaVidwF66h5gpdccllOEa7G60AEGMByhES8NMbmOEEcZPt3B2
hvMW8nYSwfVaVyZj+JYzEMUWGEToCr6mSrPHAlVpOw8vr37RlAFKAw4nWqlQXgJnFrKiDlymtRsn
7BgZX0sAaoiQXxy+k3G3nAON6DxCsWTpt81axXximQuAWRv4lf+kWNkf3noG1iDQnURgQKKPyg/1
ss/T1q8dyLwX8SW9LZfF4AmWWbjMYu9e08rLOOL4TEJhsgnutgmN+KcI9Tw9ZtPSb6Ggml/V5bfl
b5GltI7wnSOGMRzuQAiI/+R2Yl7fihhjX3KcJoIkeIqCJ27utKh1Ot3nSy78j8BokGYtiD+IVdge
0JtnRAEM7oxGLsmJJknnCNNZPFTdO2I0HTvVUSMpep3o1K1o86T6CQAePjIut74/OfRa3dAc2nAo
/3ASRrXrJDclrfEKUF3y/44DB83pBqlKupsTq6INLuVpOn7xsmnC5XcFeSUW65aVXh2wOJV1lm2u
3WP2/zIG7rCUXIXDf99wz0SHa4coQOLigB9GrFXfgS+1Xa5RPftHRTTx2qZu5rdZ7LVPuU34om+s
7Rc8QQ4sIHwISGtPRyB4BxEHU21VLp0v5NRCbvc6IWvIqEC3z9zHWdmUm3e25P/bIq0mkALVgnvA
nv83s0hvX3/OSW2gBKaFDTdYItcmF5D03yY8M8InMvteHPIM7yFBvkzBKWQMcpI+CvQtKpAkFAy8
7mCS/f2yhm+sU03J+Fs54Lou6N9+H5apfUvqeqWrUuLQ+EwOF7I3o2xoeqYoNEQXO66v7ERkcJL8
ESkuWwb6+Jwd7cO0m8Vde8mGRG7+USN+x0ftBWo4ZN00qbD0pJ904iWXwcVnNNcW6GcW49KSsmQI
e6qabwNoutr1n1oWtmiUOKeEc+fp6DqCL8r/q/pa9a6yexxQKBcMWLFNzmPf9TYOo47w34+gEJld
3XcM87RasSmCdP53GAr3l3Av+xp3is3SfzPl6tto/OijbN4wdM+nDq7d82dkOS2jLSHN2TLO8C7S
3x347C5/1a8GpNil1ozewoO+IY6KtiS3O0AD2N4ffBCtxBplnyRis9vRgYP6iNn/DLntE0HGxihR
B6yvxnQp4Dq0fr17oNcn9AW/nMdMPBZ8JMLjKtcmYJ5XA0ERYrpcAeied6t/KXo0jJGKPFamZ+oq
Cw5+
`protect end_protected

