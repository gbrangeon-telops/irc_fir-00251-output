

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
QA13xX+R/ACi8km79qumYiCoL95/JTNXmw/Mv/Sollu1nSewLnwk6qQvytLuy2zqP8g5ZHUfDkXy
dYJVTyRzKA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
nii8tC6PWRY1wcl+Yj+dJQmorGaa82N6txtyUcQdtmyxn18ohe6n/SpcWdMXBCN1HiV+XVlZhDEw
KvXEmx5H6nBr5/f6eVRIc3k7vZjXpluRFM7lDsLgIpfE0fW00UnX/0rMYgmxn+5+4dG7smGpX72S
zm4Z5q7tYiBa+z76ex0=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
yppU6wpcO6vEUEaOZTTT6jS7XbaY+e5Jeh6nknICBRlkmT5DzQmd7eWK0ShMWSlNt0Fv0kuxSdt3
PRQVKoJayZoHlh1UH0U//6ySDV8PrR8ZKYbnb5G7lC3+6hAsVS0WEHoXFsxe3QTXWezPX8OXISSE
YYTVzXqeBUtBDqueK1cvQyMM7IWnXgyQ/0dRh7UmnEpiOonlQALl1eEnWSxVZ0L5cd+jDbcSlWqj
VgoBh9A+IbjGjOjE8FOaFLUMzvKXmpjNiGzhwyN1qXczrRlE54AWkRUECVVEGR4zuEA7VTQH6H/B
e1HQhNsFNtK03nDJRyhoiacaeHGOBo4yneyZRQ==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
xoEHrB3Q0Yfcf3MYYTBHkrbmS0WN00JVFDeAhGuvxPP5kv5812Q+oIM0e+z8RwGLEwQ4F0j3UPw9
LR04YDkbyd4XfjRJQED6GhUyhlVHkeZ0vYn6D/hB6y5zA45LPFz5aqbLudigfR6lDZgyof50XSaT
wkqaJ1dNbsbYXDGYiiI=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
SZoZou8zrLQYkyuoYxGz7q7TKCLXDf41gJHR/eNOYbjhVAUcJLojwHpmGq29Knnj056DtiEpAnUR
HkNwqIIUQ/PzBp2ZRgLcYUhgAGFauW9u5fA3Qe79SJmVAKU55R6eP+5h6YaMx1oo7Myp8ZHgv9LK
0atkww+rNUFhc/kS4ivaypKADJgY/Slv1X55We59ldg5OMI3+jFcKD4Ow4Gbs5tHnIUzKQ507yjR
1wg0oIoTMEm7GhN3wZnee1A7XeomsW7IrTE+3/M1cRWhdrj0rq5nqrI9yilbmzqQyqntfJK6N8Y0
QQNZFJ8oCjr3X+2kFBb+Pd3/scpZe1PtOU8TgQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 20896)
`protect data_block
zKWn/puVXY1IR+Eg5ap2wTCgRmQPr9fxj88E2V544BE6x7jbgUsAIdWp6w+BYVTwX+IvoVHu94pG
MWDZWk6czkeXcR7kFssWVv6uVpB+/xeKck3vvjCEVAJuFIxZ9qZyLlXAbFp3AeUEEv1IUypVExfE
zLPM59ZgL2QdZxnBpDlpdvc7BPBUZKFSWo7pJp6Gx4MHYzwn5NmUY7iEG08dUA9FRYKvhGJdIKvh
tVBENKdrOzbt885pVOn1aWwBPRjGZFZwAbWM4JTS/aR0PfIZmnRH1nqbsBtCqJFchyPsP/OCgcfH
m+rRjCT1xbHHJ+I2yfUeiGycQ/fRZ9e7jy0OHA9uiHFT6ebCvSsOoSUyiHKux8+7IGDbGbxWyzJ6
sMbyPDdVqJgNSAF2UlHV+hMXkcw8SinD8ojX3YihxuPVc0DRAqx7FcIeTS2PYEzW/m95QIaRZqH5
QCEfoL7wFi/5SYnMw7r6y1wFVkZelfSOEX9ciKZmR/3H+2F2Uud0B2ovSORZ5BC5RBDfDQJwmrmf
0kcVB0BnazBOAgyL1NTWHtnIMsk1xO/ucpudo4Lzi9D8ebeEyHd/VRg9EaMyoISKuOqwZk0ojrsg
Fpi62XDE7hLkRWLkK41ptn6S7efVbVzpCfx8FM92MgGLdvfeX6VgPZuEF0lVWQpnB6j8VOTEf0CU
jjLZVsUf48QlgaUOiKFk+oWFx0W79fCUBu0AnBQTnPxEGsLYGygv4R7uV/n2+9XEWuA0qSVJuSj9
+84IJX+r1mEzvrybLHWbjwoqbAIGufpSR411NROIleo5waQfbTtorqV0ByIhOnWD7JyYq57/A8V0
V6/npRMja+Dpo4Ced3nDKASBBdPiJV+pq/mFPA0ZbcH25Wln+dHR752BmaAW0UbGwrOfz212t+s1
eBlKLAsQJrSIvMbyr14QkoyCSN6hcAywniupMtKaCpN+WIOdCn20YuqXIQ8OnZ6MnvoLxHFuEmqZ
iDY/TDYr/eCkDv83fu3gSH65rSZtt915fxNugWMPxgCzezU5A9ZD8z7fHUPQNcOe9c0rZxzBna6N
WnRgDi1XJglhoyEBOImr+eRndnb9SX6BRe7B1A9XmdAMTEAXJkRmw/exa/DLT6HAvcUD6xrWHuq0
5b+qi7LJlW+R3y59rJWVNgGUFVds0O5cwIYqUP0y+lUFWhA7fqKvkEhtUhNJbDKnsz76k61yEjpB
GXdXdU/KTWW5Bo8GydlyGREzA5t2mN1l2VC6SQ4sPHYPndXgfSzBUDBSEWitgKsLwd8fidDBdN6b
Cw/bh4B1tMRA5pVQRE0Fx8l6+HKIBQPnqHDX5WoB3NVN7UuTsDUjjz7DG9Djb7DG+bYIch2gsRWQ
xT6qWSpTDEEXUTRtVH8REZWN6IjDXewBSaxfkVkcKoCxB5Ol4wfZ6cEo7npxzUf0Gv5sddU+oST0
pXwXpT5hrvNHwrHAdYx3PhPhtzg+uxP4i+l5644TAAM2SnZEd87T+LrgOXxC8KTsC396DoBBT2o9
vPasOZreuRTw5eucUmRC0kegIb2xaKKeASOLtJYVoYYTSZtGNolEGrptpWqcah/qatFzisZprc5g
74Vy4Dep+CmP7pfVcfMcrPKX1VgdPozTF9sIwItl5EeSrf6WGKMhePSciKigSrEEpQbgmBtNpPAN
ZZkhEGVtJZcvFhzhq7sVLIJ/NWSQPyajHlZ1NPxpXHmfQt38uFgfWMwiep72YeXdpJcXeH48oU7V
1zREBzSorZAIwln9fTZIzdh7O7wXePVBKPnko6iBNFoU51/yRgPi48ylu1aCoBgnlgfteCxe3KpN
XEz1yno1M1xYFLYbuT4MCb+gb+zm5+XiL2GsUJvWlYA9LL/gkb4BYSRzQ8wir4D5ZPfH48tpbwgm
Edw69ac5hMVjdKju/GO0DQ8S9gHuRE1ebXmKnGt5+ZPKnK+MnXuUL3f/SqI0G28sRU5Isg8V+zla
7j/TufX66CNK0WqYZ59NptwAvF2aFJ75T6WcqL9ZkfNxjIexN9kpA84FqDLM+1mdPTtIfSkpGXTg
wHlDa6XHFHtqSs57lR36s2cAPdAB7IDZ3VQHOxNoHOnhiVGLM3hMkrstduMbR6J8hm18XJ25b2Yp
TQWjZTtDBwHcleS9LE2tJs5FXp8JS14BzrY9HEVomMM8VRVD+h11XDpYXkTzqEFxhh94PHqVx4I6
CWmCqXpmWCILIJjqX2tExuhMoLRLge9uOIPLKvJJq/f+8jTuOcZhm0EN+f52mTTjw5MoYPoPNT6u
s/oYBcbNwdESGTcUFc7wGhMlrFOXOps4K+HsTTywDRQgbzLsWthjRfDygaWKgYpmyA8hWaVrnzlh
uoX7TLrkWVEPSClRYmUmLDkGqaVb7VRUXzGVUZpPuSGcGwjPLbzdz4EDnw24P/s5p/V6NxHKXeUx
uA0gvq8SvWEo3tM29wDScLz2ZdKCavJgJ2xshGzXj0AZpM2uJhJE34ogSnlWqK8S6t2QQ72bYg8l
4BFKfuj/ng5VjHecTB4ux6xVRBTbOvU1Mk3EiVcE+4PdAMFYac9gaj2Lj7PWJOgIhTfl0mqqflUW
aEN//3eobjUCg3SxZhey7BS8STwP+BTSFTQUbgI16NiqglWDFyyJP/QR0uXXn4i2rYenmyw0z2jo
3fMZQqtmrMzU/w21olmWK14ZDpwfV3QX8tUGxgn9jWSbN2oGKkVPQ0VfwSHJME5UHwChO++YP0G/
nIo6vxTGVdQPdoiaI2KjeOBHGG9x80U/Vp68zAk1EGJNV+SI/zenkNgemxPhB5EPh866vbB/Cey4
jRwMm17z2wpUU/iwJrFnTUsRWwusmOE8HFljQ7hE6U1tEMGRS0kbH+WKZ+GqXYUVIDEkx/sNnZ1D
okBIHLqsIYRWHs+viQiKDDwnl+bwQrlIAtG0R70UE6cweQoBvQrfS7E6TPS+xd3oW8nY9reN/Rza
s4Ik2VXUbg5WK+cYvnXZLtXdP+F01ckIoxsA1N+uQKP6wFSXsodlCYy2Ev6YrSBzrIpGyJsvei8X
r+zmwBqM/IffT7XaqCWgGaoaK38kOrv/BlegEQ/37xMpmtYBw+sfHGIGqi/CClXUsf0j3bv4aGva
OwRSYPQYht42GuGzDAVszZBeIarOywSMP95oK/NZv+c+mQZdm7AA8PV4H0Kh0l2mxuLbS6YRcqbO
fheAQxH9n7TvHAZyTE+t65q6/02fFuDaGCjWGDAAjSijCJ6m7RK4nHH17QerIxjjL75VAArYYDHw
2kBR6BvADQZ+RbHEXcAYyZuFcFCoc1+C3l/UNy9K6cKXrUzWOYUYjiHo2KY2XGi4ij6FelpheFGJ
slwcj9JciRjCbQMDeLWfNrDFetvWtiFJSOqAYGI57G2l/z0/Hhy1uZBbX1o6tN43zMpxUOYmwi2I
u3N9fhBGmG4HKU/GMkOD8bfO4zmM1B1Uw+mn/6V+IQms2Avt1hb4EB7DMTD3HAuS5/wqhgY6jo0T
8Z9sqlZvjPJojhB3eHKIv/M2MqTL2+to3xvnNN22fEFAntoh5TW/8lTCLi5mCM0RmEYea5RYXWjh
Od8ZPFuIfWRAFV0l/ipFLcddjgI0fUgzyQBTvfjc4f/2NZisi7rg1F7qjtVNWfLJBa0J0AcgkB1j
r/XEMiS4eszCF0aHvcq81Byyxlze4GfqK91TZ+8bsN2HLDGEsf/z8FEZWbBjA6w5g0OwtfMgTgmB
qIWo183b5c3AJeXB7A66I3OB6x0m7PUtwedQpc+fmDOBTvuF+1l5B9oHgd2/deAD8bzb5GJezYT8
VW0GFL9T8FcUBuDnxFDd2JcMeVM6vXzAuiCJ2CHmVPpSC0JzLom0bHglZIvYqlSjzg7lht9ZzrQf
abDAUMyZco2/Wdpnqki2S5Mobd07uSDBDwSwtAeACAo1VRi5hNCubAw1nJQRgnOQg3mYa4SESTmE
TIBCxmMlKyhpKC0jpadYANy81FekBbnZ0HYLAQgdn3Q6+ly2F+hjZy7KLLEncf7Mmgl8lvHSHln+
opNZbJ1rRPv969vxsFfALZbZ1eXxkZse9iTNzxw3jV8gE/Cg8qpY4LFTD+6I4uGNoHGcX/WsHjqh
8qkIX0oNNUguJS7dI4cF4zdiJ1ExRJoeKPBCVIIXN3jGPiGqzFTlHJFknyYYK02hxWi1rDluUQBf
auKzTleESpfWM4c8+0jIDcMv+iZ2YpmLbtihBI4GrW/3a9IKEbsvgj/FHyydQr+huXtEMj60iKc5
UKabw1KSZEM1WnLJE+7aBe4y7qx0W2ECy4IK/ggo1hnlfgM/I4AcZr8zu1I3e7N4oKAvj9tyuRLs
tkGyh3HmdJ9v+XcKj2yZ51oxK9TofCBasGacw7PLK4gJZeCqZMD7kVZHCadZSI8j4es46icru3Jh
EPiblUtPbj1nJ7SbOUDl9XBif6q688c2iiNJw4//SCGq0ZL4C8saqgpL7KlaZef+j+jhfsQnw/x4
/pAM0dO5tq3n/FsbtrmBpJa6HxYYPIjLtN4SqYhmucHgT2NhK0CCOsrVUdMS5iPGIYpCgWIym/UZ
vM9shX3dCarikY9clBI/SmbBL23ZZrcE0c/TvIa2AjHW0gcxVO+uw8OQhF+ODZOgVkDupOV2dS8N
sCPt0iwwIMh+1CYDQw5dN/bCbC8fGspb5kwlTyKcgaqHfht1soGvP29GREh9HWbreyUukTenlmay
lMcNvH17WWCtvIxcX6g41wvqiL93HEZ4gDyZATqK6IW77HOtH9Q54wQxchbKbyKg1P8r+RIVAHU7
KCqR5i1Q6stb85ps/w5Kpjg3G6+CY2IQevc/cbGQiS3776yIGXaJsBauQIIqi7IV5ZksUBQM4NHP
5NXskyIL1OvCZOc9QXuKGO+i+lGv9CTydbk+xTuVule1MVZaYNCvg4Ipxx7cU6LJDghklaqzlwfD
EVqpg36Jb/qebKPKZUpicJY7Lw7CBMnzd19kqo/59E6wZSSKnjmpLtG8uk9LCstvvOf2D83Toj9v
635hujAh2WfGupKsBTX02H4IBPn74K8qaXmpvvYPMiXBOE/5GlCxm7sN/OEwYkcvP+1iATbmq+PQ
qcZmmfLXtEOfbckpEK8p1NUDq7ek7Sgbj+1xFeou5NyYWP8PNY7LxuQ27ri2fBTH4PiAFo5r9hMz
yWwFqyNaivbzB7PvNUgPm/izJCkywNL22bjO4NbU4wyLaqrtqqroNsujJg/Dw4j6LYPro+eJIbIe
QAdK99IkeAF2CKb4o1m8T9waya/knWpUCIu3rqYv0RS4xSIwIyhsFRzicVUBSPggD4aA6iNxokmY
PVdk/CDYEWzLJgWS6bnw+ROhzj7zEErpawPwpclNjGvc74gtpTWh+jdPEHaRfU7myYqS/dDTNLE7
PCxt2HITTjpUYAC8CueMoZZ2W2WmlrqpOXdaY0zilJZGoRmLsOZQLsTekCtkB9M2X9IVdOx29mlR
Wtkb6tjEh/SG/zfjCUntD7TiF5Y2y1wxQ1kqU9C3b8TothueZi6vrX4zVtpeGyhNkvGacV5Bs0kq
DnM3vakY5JsgqOum256f222t/k5fYush5kdCeo2AtlAjFF7EVC+sdzj/GO+tpUsDxg7hqhOn++HD
qw5jS9sspbjhLihvQgDdfdQpKDhv3TAEBlElquxkHhLjWPFrLSI7cM1GPmqGLj87dWqI4ZLNECMe
GemmYcHM1/ahuPH2zCBo3NphKp1RIEYDlPiWRmDrhczlFcUz7TMpV6EgnfsYF/MGB9nqurAPWJjB
Azx536Rmz/TkNIR+ZbMKWqP/mcy6f32vQwpaQflw/2xwzjAxgd/GKRgCWEgIsm9qv0HvpbSsZs+y
mb2gVcfRCybdUqgVncHyP02XPTOliHsxw1oNyocASowHKALy47J8Ylj/ScrV76L28o9GHNZ38dVX
J8btwOTuX1s1ommWdbyzJyPSi5NtwRxleDRtKKFIX691GZrsjkcrrIu2Vy1yI6hLwscv8YZ4Cuyp
ixKmOgtxDO+btl/GlyyFuX6RWz8GK8NcTR+mOM5OtH3yMG3Vls18iPEZSDNKn6Bl9NMSsnnLuGVs
l9F6v3yY5p5kcMExMT6hS/2XHehkUtfMImWtRUKBDiXNf5ARyTBP1xJDCzCgkr4oInsDFkDDx5oc
k9XSLx/mGGJK2sSPNChz7ozzXcMxzSjnYCldfm1xVeXoAKS43/GKVQg6YnSLLMl8AWthyQCCVbAd
L/6yD4u33f53RVYdowLgya5e1m+I9S6jukRc8jeGtwFt1m/520866yl/UJR0uyjz/uANOBkUqqKu
OUrXpW4bmZFnUqSbS7roKPLI14Lo/ssEnbLfv2TTc3W9dUej4nPkkWLjM0aYw3J+ZH/kitnpaU9l
2FWUononswI7g9c5Lv5OC5Ucm5IAUijyM2e396YJvQnNjyitnbnxtYq8VSHCwVxRkOqptsOuw9HP
7qALX2iI6G3j8s/oVDZLC6cDAwzS5TvDx1CpaOwSi84O7FxQ6KXQxdeF0thmoNkuHVhMI5JygTMX
zbMoO41DzDEPMwewecBaJMPGffX7CGcVko9fZ0JaOV8u+En8qzntyCIqdlEEXx9Swi21JqE+HvIp
SZ7jJHz5Qa+txgERtPkRGvUyCgQ2OcNwD2oxtYCH1poi+FPSUSq1r0794WSkbSkt+8pNgdOwnxc6
DWZu+v58cNS9hF3PkaZOEuWSVYzp+EfCYixupw+RCkIL5fpV/hFAgjrh0lhQV9yKzi3UITQEbXTd
lqbX6Kts2jKlAP0MFU8DFJh4ZQmziNnJXmdIWzQhsx2IEIYjl2SwEG+JEwOr2Phj5SESKpWyhTIW
khTuXFBvDoJh/mwOPAnC4XxqXDns/dGqDAhnyNOFZdDt39A9Ok1X/CkFzy7IHeIAQBbjG9BntdSJ
6get7KlotIFXq7aPXfz4Dg+vyxsRHu8v4N5Ii46yK3JgymTnJfaljyBBY0+df/652TYqWeM/GQ7P
20wWYrLB6kkeAoklDYhUerPOqU3fYXKabSCLM9nWTllUoviH2V4wCkPPBGmjZnXnTncQs5UijEdY
XhzWqCn+I5D4ua8nRZ/t2ovuGI5wjJxTZSVp4S45amh2Y+llYQsNxzOjD34YAaPUFnXSgWmFjZB7
R/IxrFa3pPVpSA2cF+671RnZi/amXH7e4rODgz82nCoPqMV2sYpbFsO7KnsVKFb47Fz4M9wW9xSX
teFtSWsfqFhE2B+gd+ycRtNC16OxFZBLFucRA7z8C+i5F/6tHiqwwsGF7utZVijecQVLnTFA9UeD
Eb0g8xlcbeU3Y6hV6NJbuv6xOBlopNm/2XercSsEOj0unIgtkGuHzVtPEk7M9SXjOqHY+Ls39Sgb
qRp8P+5LzoI57t0gE6Swfx3RWVhejf/jMvmBmT2HKyF5jG7rouIkuMCK/cRDFUCwYRXywL+/3Igd
La5iZZW1Hrri+raBZMMU1PJYS7mzruSMjxAnSLYJuehbsLLVEcGuh9l2V08jfm68sz6WGyiCJUNf
htyouBYyx+MRh5f35L2rtODxwDLw/u7rRK3sL06HexyBf2YXZOqaGdATYX9zu+MYdwvlBxyDGt92
bKrdve/tMdTS4uwv2B0552Fu+rhfp7cZIQ8NgkQpw3+FGtbJOU4un9VRZmUgF+6Qm12x1TMnflIo
obVSRjUmKsAChLnpnRxrX8T29/CH7g/VYIwub1P83naHKVAZXwWwHuqVLITm3mHcYjzJlmhPGS4b
CDasvWyaop1AGdKLPZ0dbE9SA9hjUvBsC+Pwhym/RIMVJuWl3nzPiI3/UKWdHZpAREkN6iNeAplz
pHxnlbOc7ABRe+MJdzIspk0JXOUUooeU6M+2nkWPqoux36P7klVoQ0n7v2j6RY8ORsL3/uU2RWt4
PqeDyWUu2JN+d2jPvlMMNcp1Mj2qQvhX8og+T5lZjSubw9dD40bIuexJ0tVf4WJGZE8DsSej3ryb
0y9KjmT3YW8KpAHXME1RJfLsjGaemX0+fMiSBLUVpE6YJOUkfSivhsuDmJNp6+NKsZlAMKSQExyb
QOa6IQjJEpCLGHQiTg3vushBnd6Xa5aCXBzeBAZQjTJo3lufB3RIgziiYvTJ0VJWB/j1ALknLHtn
kzZugOOo4fDqvZV/4pUjExatUhTTfqGHqamjIMfRZPWMVJQ0pWyNZ8GA81nxUechiGGYxcqLbt7l
976eSLCKki47QWp12EMQ7ZmPXmx4WjKDAjH7s8bZXCDKOljLu3Yky2UB3fdp1M0lMvFFNEWJM/PN
unJ+yxONu3erMAajAtzGxeqYO3jg0bo2rRAwj7nYRIMj0H2lU5a5WhZaZegP5UCePH4amz1DEjB/
xZ881RiO5zNeQfYolIACQa5jKPcIMqjTL84EQ5e8ofnJvVV38srMFj456Kymj1Cydl137L85qwVL
Pa1eueM+0Fc7m9YsDOoyt3xgwlLUfTOGQrUUaBfdBcHcJJxEE14cDqXv3+CcuvdyVx9shfahsa+X
KCZ1YPMBb/oCUYHPxVgpHtV3lHCmMscbqswE0B7dz+DIklsLOKeu6mgkerJNQ8n3dsDkF7g5nSlA
H2S9ynGnSQNacHXzBURpIBJsiVp0L5J8Ci6rbotUO/f6+wbHk+cfs0YE5cNp4hbvxxqs4XB92Oz0
nejYrJUbvEqV5jEpCi2yvyY/E+6IeFB+G9ZZa7yL2nfGY8nFDtXvVKqCoiNkQKXMj8vHajo/jBd/
yYKhI/RGoqgIZmVYOXX6pCCD/1HegSXaqLEdFvDZwsSRKZ9OksVD0S0GeQU2aPe15FbiRL892FtB
LdrpJlCLjzjvpe1ueXedz4TWpYe3o0ElR/d0P5HICwkqUh2iyPBwNoLirm+/tKNg6uDMHC8NgP1Z
vcSwQZQbXgWljwc+RxdqwTNTQMpGYNjwQLrtLmw/m6q2kUynu+OpNvp3HhdqjbR5vK0AT1OFu+Hs
YSGMCuHymuIBgKLe++keKaAnfyLSUNDhRBaQH0ZjIqH07IrFI3uU7tFGcmEVd6JU71b75XXtOLq0
KNK85qyWCeSxcD5/k6kieeS5fWfQUsn0ngncUp33TOXgodo4BjHLmp+Z0qKBLo2hJc+nCTreBVB9
0OFgfYNzxlROAofHrcC85eVKgfDG4TVq2lTo0H7eQ+YgJQGl6MJkdumozmSukLQ3P7NVxlJPer7r
CZP31ZySkWiTuJ6I0Y/akJszbShGcmqGPipDYOxmtz+eAncGSteZHKVDpY4f3FimSB3FdDFrbVbu
YWBfA3C0nTUm0c+9l4mF8heidLv5nIZ4u16LC9cZ675ScfrXEPSr9f9l/ekJBod9tHmkCbi0FChN
o5J2BMExYwzkoC8W1wMCBM40CpGMltI5bKsurgVAWUQeXLH8gDm6PUGXrfnlBlsJSdplizk97O0+
6d5fLRh9yef0HESFrE+JoNRaFDrWoLmk3QVtYH7Ksue1mvuZsTtFwWOea/8RyR6ExV7uFL8F3fQ5
FgT1ko+UrT9hX2OuCAQTl5LdjYufN8Fn2gAvf6u9MuArpk3DU8NDR1+YzrG8HMu2mRHsTAeKRmw/
kOCRfCjfTV/z6xIOUVlh7NAu2gd+RPg3TngW6ve8KkrLUQuIEYCuTV7LCdomPd/yc0xEFbgfJfDY
YFDT2wRdGgGLsFJHC2hT5MavBAvhJL6iFm6qumwtxY1+NQ06/4LhIrf0Uvz28hXroJt3Op6mehYV
GvHPxm95vAsdY4P9PnHkK2BsKIDfeDd/Zrp81374iBZVfmIZAO3LfNgBvGhuLHSCHmLcmSWaVyBe
r7QA+1UhLpoIfcXvQhI2+REfMtsUShKwLYPSdvCWmIIRVrCSsrFNYsfQZ9ub/d8NMhFHIqnrCbpo
90baZGBxsLrMxshBXHDi7QjG1P04xTRuSPNpPZQUHBFdoAswNOf/ccD7xr405pYbt2K4Owr5tfZY
OsCLKVuENyS4V8QTtL9Mm0X04rgb5rMi1G6R6KRx7n3DxgZkPfyulL90ERiua8B6QMsG+hL/OjMV
UnQONbCdzke3rXZybhijtag3ULmC/3QrTgkNexsCj3f7eCSbXjY3wecMrf3keA1R1WHx2V+jOEtn
UG9A/eGzLBTOllXIjD1HCBHvTP1NtgXCWTZWgufDEp9BDhL8fK9eYmb8feHw83eZjgo8g2P9mRnF
kwOYlTFgD+UUBRdNIZ4oaTSKSExAv9mwb2vX7aGJv+7Ufvzkkypc/HNFOr5aTNYiCcmdBTFRCPFY
0GMtFVezQeqhGNLnk9MJYC3R8NKRNd0FO5mfQpHaQ2pOz5miUJxRexo3elvxJPmB+YtFdQ9CnkMb
ChqS0wNk9ig+v2Ah3DrQvC2JX/af2tRnQCMg72szVjwsVceGBRzzLCKz2lEkNQkL2j5uKpzQYART
Gjxt5gbYY0JeUeKpgBWIaIwg3NKIMHMzXROxceV8UNfZy0Mp5AZc2CUVIkO6rb1IBr0FEDzXoKjw
3VjsZuvyhLxeEDsc5lLHDcAu6eBgCltRN9WOCK9yhD9A1M4wYImlkMzsX1vzPYO+jDV3vPDtsMbR
BR1mD6nmcYJ9G1wehsv0KgClKUNhwf7Upo3LMwCVOn55CuYilRfMSyojEBXAjojC2GxOt2cZgCmb
rt6uGpK1uGxhcY3s4QM+lecdhV6uu8oKfLPwlG4LTXh4mIIzbOFcoHpCaOQBbl0DoEhWbQf0mybT
mGnUktbyZsjHY9fwSyC4wUrXugrh1xbmdo0DcGC/6cTw9DmRkflZjRiHkx96NP0D/Gy2xYQ30s/1
Jq+9t0vxATOqcCCmuIhlE+o3UHrJyqksFm0ijUrqceG0dk64PVKADikCQns4mXyb1Hiy/eDf8lcZ
I7vTrwkIYdeyIzWlD7SyFrIrZPfLIVpoPe2CttFTZ6fdVr5SgxnSxf/N+XckgZoRFHSQVNoTq1Q1
fEZ615FvVCRo6+54yVLjSvPKKOv1Yn32dJWiAZKawlpijea8OBwfXSOZ0XkuythcrQl/9MjOw+3s
DuK6n0zNFDOno+1oxRhGzJQ1vqRkV8OvtHK0Uns87+s7g2DSSXMveAYaAgWzvyFh5e6LVl6tklen
rNN0UrM2neCTe0tb4NlJCI2DWqHUoEuHWqRDd5P1z6pzz55k8ZrfWSTjPktReqYz4LnnA2A+3gKq
mFMjiPIQ7KrA3vXktC8EPlu10Ipv3ard++hwsj6u40wclCy7jmN0jEBbP/qXJ8JcJ8a/aNMZY8/J
H6mDWv6NtglJxhsYQQn+zlgyimEykk05ap4LiO2/PewDm26l1J+I1mpBEPgsnMWdYgtQQUo4SsJn
IkhpZGL2aRm4OgniEnVpAHCBdgyidYHZTwsleGpYF9KABlDMoij3EiV/wN1HimsBLny6QUHx7O8C
nzG7P/OqbEv/w8MDhSws6hFo3810a65+meg6P2kw821pNCM7QtpIBTJY6w6obbkbAjGeMXMUOia0
O1nYNgiO5wmf3eWT53L+4qMA8rGKhCZvfRsoC4NpqAQNfh5OupxMqOYboNEQKaf70qtnL22e2VDG
LjandMX96t6eWhy7HC6UcdTZ5b42bVT1vBWWFPcB+gk3BViHlZK0SSAPjrszhVQFj3evSIw4RsGi
7JyihxTPTFS/CkLXi+aC4fG7e/xiyH0Eu1GenDgyzsnjxkewpFQ0fyg3b+UhGtaaDbSWgODBkFRz
+w3wBUDoIlKGZxokbowcJTJTamX18qW9WHaNQIisk08ZTAHO5f5jqoxYuuZFs0gfN1e/l7lkTavo
m34kXh8jH82l0V5UxBCu5aGITlOvc2OyNmS1LN+T1DI2lLRt6sfkh9Y8c1q6d5wha1z1RBeZx2Vn
I3S2K2JDDN95b0G0NAim7LkkvZAeu2z0vTA5z155evLFZ2YVPiqh+ZDB9kQBdlxTxqgm2Cr0/T+n
OEgASvEKbxy7lKoHodITe9CgWEmMkzXpnH3CIC10fzcRYHHqM8I0iElUkPR2uQsdo8JCKF0l7pNr
n62IcysHArdCBQ42J9pqBHlEM5penF6J3bKeMgN6YRVL1WHQX1jSuvI4hbq5sqiS22iuOo2ymCGA
W/3z3OxDe1bsFOg9e3chWbWoJmpSiFdUHhuEmfaZTgOBfBZpDAMn3POlAWjV8Q01ymARTulwL0Uz
uhJvQE9eIe73Y9zvTSwP247g1CO7bpOUi/hKbeJoIr4UlPuQZQosfKgrV3y/z3GjgLlZU3zz22Z0
kp+Fhwm/5LUe1Dd0DD7aFfW/P6hLS2sWj7sPrVrvAgz30OXJX2ueqVed39xKArE3qEOpGTzHEEHs
PVDGgitAJ5hDRuiO7mPJqhWAP4+KW1NWnUXgL+uXFq6A/HLQjoMo1KYPZsT41LE2eSKIk8XVwuH8
Ev3LkXK3QEUKH8+cUHhbVuCLYapzoAHU2kArGznDONWMAYIM5xR6RAws7txRa6/aj21aI1UWUZAG
R/ZiJWTLIK8kZ3PgWRs/c1eWstpIUtVPQGgInFSPuiljmalbYKX8ou9Sxdk3TLzS0xg63Teht7Sx
K4S6Ca8qyCaqFr6JjelvKOfN8PKvATy68OcX/NcrtklmPz+6fqz4Rc+eYpPWeyxSu2H+gVqYB8xF
V2YUcKA7Ir0PlZCocE/JLKPhNkRVdHaoGqop9u+ZHQrN3DEnMCIbvo7U5nZ/lu6dkUxxVbnXX4E3
9nRP5zAe+qixV4laROuHX82gKaQjSom0+o76cah8A4YzJRdMYOUStx16jHdGXR5dHphDItKUPa3U
8YkzNBpqS7hq/nhKscan7tBGSu4Y8aWNQFkjbuHeRjRjcvkfGw5tNs9gXfN0rAMpouUCdcw3Sa4g
MaPf+xLkJSj16ztxxrrCUPm/oVeeK9/Qos8qEMBxbfZ4UhXfo6NPl/sQ+fljaMwDaxTTk0NiqBjY
3ppWUgrT38H4zzeagF/v4bz6pyo4JYK9OijEIVa+21QskXJjWK+9aXIEnf7UKjDQrSp4b232UBuT
FttM6a6P3m2uToHT7L9aHYYm8de2v2L5WlSlqpBYwtH0Nt9aQKWmOOY7dqsgUmIndLwOWPuarEmp
P7njog2LaVGqK6o1hRFhtpqfak78uIZN6hy6pnY18X8BgDL+AQiGj+6j1C3HQqZJ37mFvwqmxLJz
PX2ofxbBt5fvDuSS9kVU2mgqL+Mf0pIJEgyiduVkvi1fArp7sQypcQfd3agmNxwEbdMZY7iDhC8o
LjOFePIqzI/cvicP8P2eVU7ATZcOa02VVA428jyhLOGDEH0ylYPalLl81hIlpCmH8JpxbvTygzNv
3hU7gLMNFQ9nhH0JmKAZrH1e305jUZXNA8JBFp8mtp+GvlfH0ZeocAzFF3/1ebK2ESrRVSuflYOg
PICva/LP0cQHQRRanxFmqML/bYDisLGikRfPHdKO5OapaKP0zwz90LsJp7E3I71REAvauSwWxTWB
GENQNnoSvjee0XNTJMlVT9yNwZqAdVT2oGmWLrqdvHhHWEzrGY+HlUNPswx5dQR7WLYXPraMc5OA
zNoc/cB58KbxMxxtJOv3IzJbYv/gmn5wJNxWo+55055hm8EiuuGOiwemZmOGdyIo2qoPP5z3dXLf
EFCUG+4QRoEkJ3MjvvZexxPuskzGcv6bZnSHSr8oan33jHFjHjVu5DcWUG3P/Y/tGs3rgl0jmCFb
65yN5yKm6pNIPyvuCppaYw8qzlsfPKjp7ujxtNbOyyX67ZdPZEZ+Yhr8fN4RwB3qJvirFAxcAfZS
boBGP8dZdAhChHYTnGO7eD/JhdUMMCqnMD12XY6Id66lgfwzWf5rgumTHYaMm9pkPRknIRqznGjD
a+y30815OCW3kghqRtFmAqTL84DUvjC9TgVGVi6qLHbeYPLWqGJ6Wz1EtU/WhOGHRQjK2ZjJh7V5
F/Jt2IZdMdNjpwRViALUufYkWI+ufbJk1kN4VSSKP3yMvAonkOSOMjCEEnz/pikFtY6eSBvo3MWE
ACW/mmE17Cp4VCQcuYn9YWuzoyGLvpBvHkSDjVw3MC7AKQRt6jBq7Se8k4TwR+ALWf9Zr2t+ibXl
hsPRlMbLPvjDjQA/Q24UYFXZ5uURLkXY7k8erU5emaImND/mIha5wtN5zCTkANSHVtgwMfp5oHiL
B1Qw1Rmjbx/9dt9d2i/VlRkQxgdHxu7uMM9uOjEOEoXFn7ujpDbpVtNz7sjieNvARnv63vsXq3KT
oAKXYuv/bJYf6EUywZUdsraMRLs3GZWA7gHDD1Etakr71mnEP2oOxb0RUenxh9qDKHKSjTShnb6O
9dlzS11CqXB/KDX+ocoqJyEp+DBwogeTgNHD5T3o775aQ9sZJSTwHLB6H5G3SFaKujdU2WYaewLM
skJLrN5tRE6gHGc8WyxH7DiEA17OSEWRwciimIa8w5jodPkPkvPAp1X5qXMJa52LLIwWfUkpd4YR
uIoF0Gv600CR2+j2gq5tJf5p9xCI4bN5ka53nSw/KTF6bmIw6GqTzgstiEjesfQPelva/Z2dOkGK
vbAJiQAOQQ1Osqskk+L349Fh7M1BFM+zHRHJA73ztThHGOF10LApKiBFlcfPYrwsUrw+C8/HaJFe
yVK9FA+EPS1fieSN6+g+Z7LHVkAnY/gzW8fAr9K4wvRVOD/l0zgIZnLkOepD99KNikYVd9dUe6D8
7p1PZKtRBjyOiM4slUzHqNi5/PpVrPnPUWdDuVCjKQCpTX+W+o1b4OT74KvIqDh9i2mhPwyRB35V
2t1nmeHy2QVfj4rcSRmCbm54UfXcCOvQmdzQlpoeJ69IKpKKH7VoxrXsRN6ONxgiOZzJkWKGtQo5
EUxJ7X8JGmanQp+S8jx7c5E6YmA7CD9Sf7LeERlsCJIu1k0Qilr+2gNNcWG1+LmXUVpyaYOmoIk7
fYKQSiblDp/WuqKGTTZGAUx8TJzvbnjsy9D8pQdE2oZw8K9nAFJOEsWz7yP1cIrhUdfUOn4bVTNn
Q/UZe11UagWhdci23ImUD+JfyuhPW6WYFtZcKKO2w9/9FgLRa4vGao5zZPBqEm4WXiIyT57nDjTp
9eYdA0BDKRkJy55en9E6a1H54LV9ZE4bL6nZ3dkU30XhM4uGJGcO6dQ2DiE1gr6wBbbSijfDPU0b
FdDPPrXZo9J/HvzxBtM+4dOG+D67HTdpzgbuIvKZVlK6Il1zd9JDZ0Ic8knjF5CtzWmWERMTeGAf
V7FdHCGGSiAkVbqCa6JTOx2xPyTHakj5t+fyPNFH67gH617aQSeoBPIPd8sQZthCfrbdIqgb6+P1
aAGaFiVL076Z2KTN26HCmHNw+wAaqIqwmpLwpJ2wLxf8eb7FWao2yGoZEECCagfuxhroEM4fxkQ9
vPX2jGkI5diZfVupz9Fj+Ac0vyH9iIFAjaWD8z8afh2EG1fSVBjcTa4LRGecPhuMgiOW+ITB6P6Q
80Xw63CfDEITV4Me3UzsnRPEhS+vCtUdlzjpazKPeQTLnxmFST1wahvE+dXYe6faQ85LqAuEHK7D
cJqXaHhekc7jCP3gJdLV+YCg2Vs2mbEjby35sR8c7Ed6CjS62m7H4M3dzXQA7Q1VCcdC6zWAv2/E
k4Matfvh/QgcWnf36s1OahYGe6NIVQIJNIcrCx9QFaFwpVlaZic4vYNxap58aH14ECG4J+7gmZE1
FZHGKPVN/ub5CGu+ESVQdOPmQr4OF5iIVDONoQA3SFyRjXL7tcpcMfaQM6qCW4ILokNPt+CMGAq0
2G8XOhGCFdhWaxJES6cFc4vJspLnja1jOTp7fAGo5loQ5msLc9ylfnZ1ulTxUwnl9oR0bS5OsyDi
P/sU4kmlX442nwtsVrflgZJoIMyYBR9c8yVKLj733UYdj5/NeL2Dyt3ChUSG4Xf8gCeEufF1xFVp
9bzoIAu2+o+96eP4PPrTTiINBxEtnaPWfUqpx0+m2Pq7oJgDfTH7DeT8ViPaGhdeBXOfv88KIh/u
Upr7Tyns9TPcUNkNJetvEi2Pf0b5tZa/plQh+kLe0UAoO9Nm0PTgIakLT9k7BDtzkTm8ai92ePVA
OWmv6Ztxl0w8OOXUuc8RFm1i1GpdUw9OqS71MrLPZVlQ6txozuX7KEIHiZ9hd3c7aENs8ak+oB2M
fdKsxWAXykWOm1JznQ9Rp2z3N7eAHqg7cmeZabeETCyc/4mjCtrREhkxId/2kPadlHgaJOOW3E6j
0kAPI5h2SXHjCM1creQdT1vyK1VhDzDNSGlbMG2w+S34eSBHTW4TeL/EPITQ27B0dYdT3pA5wZ07
UjjLQYRFxwmFAX4pCsXcbpzw/0cHoGRrtDsqLSmeq4PNXFLd3slQVLQC62msnyeE9BoRuP3gq/GN
kJZujGcLHgeI/eKs1CyGSwV1XrIckhNI3R9vGXhDEhV1RtrYOeZ3JAbJzqywIzybAUtCAmwu+vqp
YSYZP7OyUPXD6AzCgAKzpcb74KOLjwG5du885844KeXrRQA1LoGmd/h/TRQn3hogtsmeal6wsnyx
0XciaGogZEdIY4SpqtUr1QAVGZixhKwSN/9KK8OypfYP2r0Z6IJMDib5Cgq04mo1tgZSas37j3b9
eCYwqg9tZf482zPTWvSqYgMt3BOlzd+TQjjwH2Y8JrgC4Tzs59iqYAUKOufDU/cmN5SS2ORriiBW
KFvO/NjDkk9H6Vew6T1Odcl0QvoYlM3UuMWRQ21us3r6Q4LA+FGolSRbVnopHaUxVZea2x8qDUg6
2IbwOd0LIgSbaS/i5HxqkuvfmgBvNmNCF1LY2yfB+vFvPoDSrNIK16Xta9Oh0F0O2+55LIP175N3
/gAW3KBgch4GvzU9g3WKAxs/R4o5Ar9YS7V83uUcdhVZb7Va5p7suPxb6kD01xeJU34evdfV8Zn7
D9A1sBpDFgmaaUUsiKxW9x8I8ny+fVGaxKzugBs3eynHvxRAtPG5rdBCWikxJn2I7CH5RF8kHuhD
xCZSE1Wlc6YgO5aMfI3f+uKQ/nwOeeU4z/b15ZiZUY9XsqZ/cfPMB6iNOoXKW/yIPAg9hp26z1Q5
rxciomMu/EtcCpr1Pb4lNQCQDNdEhO8cTtAE3W+eOQusCJdZOQKf0s9Qka3vHc1q4Ep2X8UCdSRu
d0UcrPBGx9FYlwea8w5CWSOexKzVEGaH81JWAur/RzaXF5ziPUzmmkDx5oKIwFieXcpUHiPQ7UQa
w0o6CPa3BCY9HJ8fzL8QyeIeaG063TtGu/qx5kwGR9s00tENqbo/ICEgLhhGYWqWmJ1CGlNtm5Aj
cbhDZ8kYTpzTCq1XiPXxavk9C0Dp/TJ8Y8W18u042TgdtNYu/9aofkyg8aX5ESVRNSgH+wmUm+u9
hjqxt5jWWY1y2UgkXoEtx4g9RqdyuW+rv4ioyHiAi1fdAmAvxWSBMIaV6Djzc1O6j8bzrrpHNZVZ
zabzkyh+JAee1lpNPPfG1CPiOUYc1lkUZH8NBPrDhtkkQhU7dP9//4y88vHhaaVYTGYothDAvB0k
ctOiRXsl/D095FsdJjVZJD0Bw1HfnRYyK2ykVieQqQe0zpzMwO9gHN5Wiwq0YX9GHP2DtFPQ9yJl
zdzL+xnXwD/4CyN0NJBF2YGjrTOFpWXCUZpteeYSmmh2iPL0O5/uKAO7xDxUa80hipY0jjivfywo
+ONIB8TuNSA6+PchbNwq/0Qsi4BO5q6Cq5zVixrpqLXUugxpU6555YST3cYVUNYigqa0kpKAdGbj
5EkIhNCi32lPVfpyndpgAl+vUiH8c+o4OQ3nzimIKf+fdzu6B0unvcD22S8SHzli8BwERX3HcmD3
4PTSPbl8kAcKRk4J+5+r50J3DWS6h2YXxjtFublTYdTRT3bFbtd+7zZvd5AjbRrdmcpdGL4YOzXc
7gjvl4dNmKi1Ru5ti7btzIaeVUiBvWdHeIMxy78I9A9ijKn6KNFkQuyGS7gJ6t7xWMGg6kczzC4O
MGo/zz5D8fcNd+4H/dLjK2TJRhz8X3yJGGEYl91C/N8u8KXwRdDml+7QEhVIzkvGm4qG0ud2OAA+
sUm3YBT41V62KsBfzulSoWMR8N4H8dIK7wM/SaqrHFn821bxEpTCTtFYuJvK6h9vWrGl7lDJRF8C
2ZpakjQBI+USockx0azaBtI5PVdQvj4/Awr3tIeS4UnWGnaS2Z9UJH0PRBdh65yfvSs3XCAKFlhG
RwdA/Y0US8pKbSBqcn4SmQpRMaWDbzxcg9zAx/+MuuwIfSxO85xckzxEOBT+WZKs/nbr4WvmZzBq
LPOS7nr7lAx4ksMWH6qQmd/ej+HhNLNK7nVvIDWGjR6ICXZSBsoaFWdE/jNoyF8rWzx5UglmH6xB
UH2I3vdp2iDwHemxopfEzJIaAhPBGVS+mcSUjCl5BU5w0gSftUPYkYViFvnl64PnJ2jJxnHQ597E
Yn9UNE/icIXqRKsoCkcAiYOdniFc+nhVjWoUfU5Fd2H5V5l+lfPqGytLYxcBh4Jce3KrrFTqBxvy
0EccHy6PyjJzLHK0QtQEzA9X1rrDfdWaOL+kneO8hbrb5rdErSiMtVanJylXas5AFB+lYj1kqh/q
O+qCRobJFa2DBLwSSxLznPEO6zmZ8zu+LcyLw35eKlYlHUDzMskOz2JqfvWt9Uj2eydeiZRI/pRs
zDOI87BZjeCIdJ7VGhu4ISFJgZcb0aN3WECz85a6tQYLZQjSAXm7Fwd5lVJyCKRGIwlLgepEfi3x
WZgP0wzoeLSrQpuKuHGRE88HFXwUb3GamTDCqX1byWTwfTyERTHG/KXPQQi4nkSiKsgzQ3TghBvt
Cmmez2RtCvtZP94YT1d8QDUGYACxFv+yJK0yTtZWoOlYC/ilb54uvvYi5IKRNQjcZEzWk73JI5pa
suRpUI6vf8L4gubZinVTZjjGNhBhQTUFe2awlrAknoVKp3dMWfwIo8r6jvywIsvZ451HLgA3exeg
hgXlUruTRI7FXUD5iOzGBM9Gzr4iXOo7h+niU6c4HHTCm+Ir+SM0fuXymjOK1jKshhtv33omQfUu
iaCbc9SQXA8bIppvM48mJF3zXO1LzuXahRMSR8xnXIEVnXWpl70nJcnay2WRtJOrbShusdBxIbXC
2iFHLpFn+50SWn4gqiyzaDMYfhMMLgWPhiZVJ+fHcIzEH2KImwtjBNeU+gDKeNwnC9LiyluD1gxY
bPLieP14tquv7Ae3K/ZA8VW8NbbPoreNkhwTs4inJAV6jFD59Ln+D9kl4YlQPSAFI2Zc6ZZZcTMC
eqABJTjDOEynVPAoDbeDgtmSF4CH+ddmyvVE9Ex15rFZU78lkWEFIIjGG8x9/J9T+y/Loe6Hqy8m
H6r3yL2EUJQkYbyrttBezlC9usy9zojq8vnbRxJV74TMhqLrXAcj6pPoBEoZd8hJvbxGsK/1yUAF
XStqsdAKpKLrOvsJtR0l66C20NinALSemH32+5lbMDF+/nmKD1TDXl2Yd5/ZtWu44OqkoFXId5PS
6JpjlpUuBshi8y1/XY9IraZgOc0EdEhMhG52tEpeTLhOxMVi7TyxqrGKyuOyRbvVgx+CH+fTa0Tz
/oj850DCSD5m122OrNFAE4G48EeioLXeAgtCNPS/34S1UHSFwDPw/A7pJPkJ5ouCXFDEMef3Ey0f
6Cvtjx2c1Injb94BbvqOJzYbCAX2tRq2QeML5+z6dPUSw5DVt1wbb3ky7wjL01RVYQSuYcfZHXrf
cZ4gT7CeAdgs8ANOlhdy3arKihNxRXUUsufCCEdJJpi7ImGCJSn7a2xD/q5fOsrs2T5hkduXfWYh
KGUCtzDAQDU/TD06JoaHLK8ES3cOO5+LP3Y/ADdPjUesljkWzJFXdn0D4WVuvnuEU/KbTXLgGyjF
HlfqwvCorCxUG/hZ6XqFEcjQDCFveBnzplGBkEaR5rkbK/2k77/cgIf4I2WMVDHumWbO3jlcGq1f
mDW5gb7Ybl+9p6qCFfd0wo3PD5kp551SAsQiOthsy1uXrB1EmqQZnc5kRhyzoTpVJ+zNSs1hnYfK
PNWGbWZnZNBwnxHfYSWQoFPpnQXWW731zE2HKyrSrjP42zqDe2AfNSZzej4xfKjAgUxY8VJgrqpU
ndK9E3lUJ6RdYMGZmvKVyIz8G7ZiXiBB3J3bUSmYiAOO4JdDVdg6fTNZBRaiReB+eMlohRId+jKT
Z8RwWjfw6KaBq7QXEbaQQh4+EuPuZZFrB047JeqAhdygznsndfQ/EwFTIfy7JvrCMYlcx0RPJ3sv
x5xod1LzI8ofIUb6t5DTs3tFAdsLfqpYX9Iqi026D+04KkyXq1QGOu5+3/28Bje4dH8XSuj5wCdF
mtk7U2QEWTt+d5wjGyLLDbEEviWOwRhbFIQrnRJ+9u322gIEYeN/75iCe854JlmpP5F14HRZ/tP0
Iv+u/I04kGidGqgj3p+aOZt0WJ+YArQDQg9072HvNgmaFhMBCijAdTwyFrfvMsD55RQ6irXRyl4x
ORO+ufxYV868Yt/YkSZAZiIhIERPBEvO/I4DwhL89li3DgPsBlpgGCiRUCRNmfZVPPGWxI+mQUEs
99cIKHIe+52jlxOzJ+c4JBfjhK/3g8hUeyEAUN77Iv9kG0XWzVlwYUaf9mhzTMx2SXx95vWP8/l8
PUY26hI2kQEuKiRUwuIT3KtOcqMFc6xPrVKxomUcDXQXW/Ig5klBo4UyyLP09ht6cCZARYcSEz6s
joD4X2a1w0k90l+Odnv3KE7e985XopTH6LbmTZ7RmnpfUAJUP6RBWsatGnuA9maBrSFlTtQR78I/
XmOfXBVPlMaWlCkWeoUV+BUbT0Vm2uAgqQHkexkM0HkjclvaR0r19pqliXv8y/x83Z9jNW+Nqu0a
Vq90TTxoODglsEc0wzHufVbITE0SJVZ9nTj9JEIVFBC9ilA7gqa9Z+GTr207ipXF72eFAmNcSF3l
zlr9L4dujfrL3HWpuY4pzppAZjjVVL2Z2fT/3+LnvBpppPTaTkWKia8YJMgHrB2IDii6ABylReKf
EnQhziUc7BMDrVGRsZIeqXcZtzUP2n8QvgXu1Dn7x72Q62BUpPYe1OVPBm2hkrp5Xv9cNuLnzrZB
4a9/lja2+IXKV9eVLoKpq+lBUi8nQkMGNcEAV+56kEnOz3NIn8WGP8diWAYoCIDyx59ZodDxZc1c
cLvzpWyLsf2+LjAlQii9o+jlbPSausEdpmxjAUF3BdNYPy3MDHNJOU18EGsuHa1JLFCf1FG1Varu
z1XVCy8sTjwZER8bAbA7qk4VlsAwIVULKwiZR8o2nesQJvQ7m1QrrmUlb5xAIQ+xd7J9mFglSovw
8hrVDFyxErkpSsPAY4mygmc/zdq3c74rfa2TAJS0DOjTEjXwNsWn6CrLlwq/1duNBQDOIKRMgu14
p1NMICwDbgaJ4yotlnmKGk8RiE8k7GXbLIw+67YsP5F2+iN4JRDIT8EDkqx8ZhvDjr8noTMR7xje
YHvccggN/D6HwjHHy+8AJCvdZNBiuHmYNBaZ2Hk9ReDDhVtOcRDpgQtqM92+hajctWBuGQAmThPS
h92maULqXEub0oOm90w3eEudEdCwAwhkn9yRxMeVbpuIh9w9qmr7zkScc2AZzPRZ6Zhiz1b38Sfx
/pvQSeoxKFDmT0MrLOR51CcyV1CvDZo8g4R66QyyGjPXLFnk0s/tz4g8YW1TINhs6bKEmz38HRFP
6W0dJSZRpI8POHvZQMbFrzTaOGgPGX7OaOrIqhiCtlIU3MDEquD9ux8n+pYM5tN5BT8/yfjLsFmU
0mSRmiYV2iGouyZo2NYcLwKFknd2yRfNfwSeGHgA/nuWCrQh1PEj29xANHMkm4YwOLU7wMbrWiiz
8Wv6BXTVGUigMd94dtY4ewziQtXZTxQ/tRVuVTZDaCUVxk0LvigjBsqpz5Hi5YW5ydXJw12YBvq4
Lhn2D9Iw8csZrf5/dhhO2534CsB8U5OJ5UA+6mINPnTONCdgGcuV8LX7tqJsIGj5EtW4JsqrLzCz
dq1YUoPIT/LUSJNDM/IFO3Ugwbsij3XQlLTfC9s7liOrNZX62kIc/MoFbtDQnJeosDoWhAd1KK5E
cZnQYejoxZumiFVPfTf64CehS1zUJlM5GAOzXezzd9gvqLnPZoDptqAt+60TTi83L8yCQAtlxw8I
T++yrsPTm1sU9WYTt7Izv5TXuQemyQ8dZWa2UGGJQVS3liDMLKc+u7Zv3T34NauW2K4pJLj3Vkb4
7y1sOoxMPny3AQBXTybk9I8PJLaAHe69+vDb+bLLlzY/IGncjc3cV1qVHmNmtR38mZt8AOPbVb95
CiFBC0GI5SlZwH4CTZ0Yw/GbHj3sQ5Y1/T1FiE0DNDxlnJJQ+8rUEViNR51NVXdlGZIR3rSBPiTK
6h6H89uB51NsHoalffdtDNjYC9t9Ers3iHMI2avOG9D9AgTiuZUOp8mRIC4SY0TyzAHpEnFcuCZN
J4R8fJQ5wz/tcnAwjOoHa4n+Tg8B1UFZUYLymbm3v2eld+ZaNGfl4RdYoQetRkaxMsoc9ZxWWAqb
Kwa9hrbrNd0naMPu/huJuZ60UMBATt2F9w7tjT6CWW4WIO8nBudMKRANyAY5+00CjnBc62rWrwrJ
zQqoGnC+9y6MUl/5PpFti9k0JQLzqbHa5nKuZRjQC8e9c+KaXhmsp9Ef2GZ012sb55WgfhdLZZOj
ijfKZuus8ZNX+d9Qort/Xj0TbId+6TCHhETQTH60dDpen2pi1IZmE9zSob8hOEDLrOpG5JgLtl+I
jHKbCB1+bcqjg+4G46CrYFkfxYiUBnoTVqZ3c00Xt0cOe53Di3qzjaSJGvKEqPX4Iqh53VWrruQU
oSFLHkhcEhrENvjMNGMu3vmnb0FPDTL6SBRtotuP169+ft3DDODfAqGsq8IdjuK5xEvYUmIJNM/q
xbmpwmsPl416nZK14XHfTFV/NYIUU0CiBo7W+OEV/j1c8c5AzJM60oFBuDFjpn2+aDFLdbGI4v7H
tM0OOh5TXrQl9SF7ZlKeNexudO1h860Cr8cIpL1S5wqjEi3OXoQbOKNxExa9fz3VwCWn+M91Rx+U
vVhA4kNpS0hmP4BnIZ9BPGnXX87l6DjEMqZXHkXF52JFREFLxk1RP8066r1Pl0hOlBz+ChF7XcK8
8/hKkvX+tzYQ62VW6DMD2sLCDq78BLLIU+CTggeVSHqQUPh1ty5ZVqvSTuty8S2GZeuRIXeG6X9O
pJ4urDGSEMIa7K2aaVImmuMUBLABC3limwWxW8q9budT52DQfqSwMvx9JJVLKjCTKf1PLmI3TE5B
dlz1jmAwjrlbofYtVLiIUpRNQX0+qmIDpNb9Bo1rfy4YfVkw8B6ox/iRYYLUwsJDkTA3LX64o/hh
eWQ1w+pmABWdD0BL7V3hkL2H6TZ127i1wKEPv+u5viyseu5gW/sqFOOH6UHO2vajWEf+5dIBvGR7
08QONbQSS8TcF/Fjqf5/5R56cTvAAgIIXqQxHbEo8VJ6N70cn3w7HCE5HkGnBzylYcw8gUEsfvDd
iIvFYqlh3u0nmPHwdajjhFYNCOEVu7tEUXXwgshee0Kl5eoU+bOF+bUGnGXhVQHCm/YmTDi9pbCb
OXF3v9YwgScpvoXi3P9UdMfMtI6gBgnqxy7bRR6+I4ntmgKWanE2ummbtnq7madu0+RXB822TCaC
gaqYIi+uGyjzmfSTmT3E7udonxb35A90fb+DgAzED09NpP3Lmg9wIIJ8BUQgRRdKlLWgOXGCZ7Jb
ehbMFWhkaTctRTRfZEhou/baDEpkH0jlYDmTYO4Y+hPvlER9StyMS80a8j/iHPRpLdlK1kOP7FST
/QlcXlleOSn5HatL2GHHvfOCr8NkfyFpl00585dt18feJkuH8SeqmLZ/WhrjBQpgLjZNytnz2css
mkB1Av9IituzB5L12vISwefzvmOTSCunfV5xUuxVUqYpAHXhQiGzXNaXscUOHUc0des5nCy4E/X7
+r1dVgNFWfhbrHRmCDTn7bqWbMgHt5J5a5pkrlU7xc0LIqlNfQhiTYaW3qS4n/nphZEpAlZTBA2q
Fpq5Dc1o0jhm35aMqSDLfHmpk2QpZEQ9GSgsKAwYzKlAcP4BcsEFmBkpmW+UPH00zHJ5pv8vBbGS
Rb92qRH0EGa0KlVzEPPI9dK9KkHAb1PG87FDGfhKQ9+AStm/25/feCcNK+D0pYcEayY7CTiEBqhZ
OlwaGfQ8lRF3ih24I/ozMVY+UBRrtncAQHARH2EpKgC4QzEO73D4x41gIIKE1ZPcU1SxMnGrYtx1
PVwo+6pGHeUkiz3Loij3wiewX/VHwI51DFP7y7eIIXREnau1Wo2y4MOvjkCedWIekklHiRzvNeW1
slCYZCZJoVYzYahnsCwuI40+JDf4CNwFWJ9G3mtJdeTvy4SRXz5z9gqX0cYXROusFlW40IHgtvFg
wK3XSQeUpVSBfik09iqsSrS/UEP+wITraZrwWF2jZCsi9QpgfaYgr7vVFu31hhjpU5vzHijpRMcD
GzkUnVs4frOFAtD47V2sCMRKxWigIkkZAOZ7+n0K2O7U7Y3eHq1zMqsTttR492oE+kv9Q80jkqBv
MNaDmY6TSvAW4GGdZ2+Vdu4lrkJkMOGVSXMnX9+uroIL6kDwP0cC0m0qO8Iq8jCKkTO9dgiyHYkp
O2FZj34GhZwlNAMaRVxvFoW2BEQWjgpeAernkGvItleWOCXwpVlTaxHo98N/D0kn9pEEWwfY/0K9
LPGMq5pqwFihkDxWrYzBYf+O67tW/t6SuGm7JFBuCE7uOWlBb6E4mLpM3k69ZV//q/gmqB6iF6Vy
s/OiETbXm2klDjL2qjQbwnuN7fE0/6Ly8n3RXt12N7ZM36Lw02JFD031Ku/uulvhx/DGwp2BJfie
pIwYIOZ9u4MhQ4YF1QZO5rJARKa4Uk0uPvyrYIbOkimXm8If872znShMJQuhi68Lypf0WDMMgHdq
fdOrGUGr6pkGEFmfqF8YskJbJdPvU+sROTlHkf3qW1jmu1IjfZUIjHf5vUBPpGYIvqWW9i4FhQeN
5fE1yW4DTrqdGkTJ8t+6qVv2FPnAh11d50HsnbQUzhCn7eT+eo9luXpdqgIFaIfum9qhEbU4zNgE
I6eAPXkYDVHwtUoX8q3V6G2pD3BuIJrw7fFt0fm5tkIJQajpXEBAg9QtQpvTKY1SM8DZGAuKSD3b
/ac2gi7sQbCMptxSitgL0vPryqWnNSYE3u6vU1XAxoMbbzsW93Dk4M1fEFAu6TACz1OSciphiuN8
UTa11dH8Mw33yI+cqLyCPs431EClXGUlSc0lcdfYaDV0Uy3HJSEbUWH66LVU+xUlFM+No5GsAw5C
h1PRviSIOY4vnPKC1RKwGAUrC63NMlEg0DxPV47AgCZaJqDnZk0WMY5gXlQuNZQ3OWGu032M4EWK
zQ+3hzHjlt01QzUHi+GsDsjkyh9088S7knwzyghdAgwAhjixDcUVJsyjCtSaSlGcShFyM2y8YrFu
nUWya9F6CHmwjAjOgLhVAd2N4h7syTXAuMwfm1sXETYS8G88xUzF67ay6zBTQg71gIMA4JoxYNpI
3Fd1BYtjVdYS7XjK1p2SXuweW5z5yKsnvvdCojAzBmfx60gId50pVRTgmDEC1eoq54TQ3/mTuETo
IbtweDQ4NYff1CVR63wOr2x0kklVnqXdwfjjMBQe46GRCgCUGbdesnLL2gau1y6KYbuI46j88whe
BDMsgzFMFn76RUsYhfWN4ly9vBQLeG3UVS5J5ORMix0WlHingMTno+cHcpLMvC4sY32E9hW7wmEe
ao/xUdEdZNHBnfAdZwCNfN+M9CwHbW9nJK2mpE7gdD+6Ixbhb4INm5ZW+IZY4sW4C9hn2sIG8Kur
n5Pq0VinibSTSeGVZxt5W3U3wqJ+BabXjhZnM1BC5UUcJrRBi8wDo5wwriZgzs8peIp4ZvRDdPXH
xak5J0KD7aJT/C43mGZGhur85F/Epgz0ykRQjNLDB9rrgxIXaemYFf4T8r2gC3APc69rRjcgw5SE
BmABNPC+ZOuHMF6KlTmNPUgyqmL1/1Tna2JZkacM/Uhle8RZbLonH9JR7eilEcqudbRhADKUdsH7
Z89R5D9rAfI3Zc4wHBnSo/qpPg+EgHaOQwax+t88U1UVaBRtfLwy5SqMam+IvVOEJ+VX4ZarblWE
1XTDpLnrdQf7KYJb2KkE7eYCXe1enSAHT8rcXDcm9dliBjaYUD3Ak38WGSBOYpsrQ7A75tqUueBQ
fU61RzoLVBpIa342/KYsMVC1Kr7IgwZPYuRRhVZ6ACLZjW0pQ3egOytL5gQm+Lu/SnlEIOKurrBj
iwTFzuu/qSpaLL801lFYLSdYPZWvuDQ2hMwp3EuQ8Lq50GvafgbVvjNamJ8znt+HVqcCqa6q7i+9
+sBK59S4ht+X2eUDMc2p1/WefS2KgDu6e01IBn3o0qCWQNo6CbpwnGdU9LcDVLpyOpMT4MsHmCYd
WgiJMsBPH7ETYPd17wFvgjvaP06JJAKBnGPMltRu4X0YkxhEQb0+UgiDz9+uA6BCw7+EqG2Uspbt
HwotyUbgxvsyVKsiu0wQJwvqZeN4fV1PY4Uu41JUYEo7awtA7srrBTvMEDFrA8AhZQPK8xRLAcPW
I7F/V1+5jPA+EcVLdpH+hV9FJM4rEZne+OrlWupQu1YrKLFAoFE5HbRjB6aDHDWeM6Q5HDSqkkKD
J9UkL7CLy11iqmEJrUifnxhvtM4BVXhDfAhkxihkHF3tMj3Z8dGnIcQJA/qfhyS+sybUktdZxfN1
g+iCUWJFgsF5s7YrsB4PjwI7SQ+ZoAY8R4v0h0VavRxyWF/EKt1LezwGOeIrWxu40OK5JhRF1VEJ
blgMSYSFwOQGc4PkiO8nhpXsnznXEuvj2olF2Dld2vISQUoAqhvsc/Jg0teLiSqEV/S2W7FHnkg5
yGPPML4anh8c5UFx8s6ige/zvIUBZw/rWf6qcI8cusqJam6Fp4rWJ7l9G/vDbP69weXYAqoTi2Km
dLOXeUDEG7oJKOoF26MXQzR7RrcLczcFRuW0uinhpO+rFYLVLD4VoTbc/fhBFHgP0pd6bjRvnFZx
rhUmzRY3pOmmz+SWSoDDm4XYnTkLuM3IHYBBoKmfYN1uPhg+QjltJHoOxlVzWssjIFf/jBhXRj2z
q1Y60DH6O3j4SGFETDWbSgpO0JbAXwAOsXdiyy7TrotWlx6tKERtYglxxaIUqcd2o/u1EseQMy9U
nTUt4PU48jBqtXbDHAr31MG5Nn3ksQln1BMaqIgiXDHkrWm7Hc4NyU9V/cMmx7xLGcF5A/Kn+nYa
bRuHoC15tniBfmGdjxcrLhJMzgAIBDBFu6bHN/GwKzogkKYv+iZ5URvCpr3DC5tDZIDAqJXhyhBH
aEBErvGG3rPj3ixHLzVKSbPq3DdbYwWW+gGXcQt0IjK0ndKeewFzs8E5UztoFnCpkjC5XPJ13OZN
DPVHDLd87l2492TsTlY4mjPkawvIP5813510SWeXCby00gJW6uTIrG84M7lDtow2ZzUR9wiUwQ0Z
Zw9K2AdsoiXInRTIBu/SsKaMCvjUwpSrqSIRht+pwHb951Um75DHhKQNIkvuBbr5XHhCuOfBpado
2Jjzwcy2kLeZOBa0qKMSECHcQJMqTzq7CGX5R7JiJu7P2/qkhXY3tO5iLDrJnZkFBqEtlGcwt3Z/
s9T5R8gHz+4o6uuFoeZU8QDR7hC4K4C5iUtxvrF+B0bURbHnfidc7J5+qC6WLLIBUtMLVsC9r0Ld
MesbSVWD3nmhUq+QQIimZvm//mr/8twWYMZ4VqfHerZngycC7lpRFsYJLk2d5xg5VKcTIYyfbh0e
rXzMdXmFVNP574ZFLpjk9BGcaWDuqeE9jV6iM5Shf+6PoA==
`protect end_protected

