

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
JoMCOWeb5WJCBfHoFXpAeueDDgvCDiGp3AckCc481MQYfkwqbKzf91lDJ35VGRkR+lnFDdba8hVh
ebdPAvk8sQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
bZP6jV/nU5x88OLSeX17wUzGVM/1H7fFl1OvjJVlfPM0WRyEzOpDDBDAUuNgnxFvzLOKKYEuQdGX
W9Azus4jUwU+zlgsaiCb1S5W3YMjUJKtbRQ/PvNNulBlTlfZaMHLAox9gfCqP4OK4hzymuRCwSK9
PA7SK6I+FbKAacX9y/g=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
38Ya3DupjVbpSJ4i6CmxC3OEuL9qNwdAvGt4GnhSmvDhP9C+krqPc261IqfCwYzwzxzaeMibTDWx
/h5fHzYF2I5fsXilkoEoRxiVUecJo1YSbQfTJW8OEBtN5aYD4EfWNZxg7GXemsfNXYAT3IQ9OGaZ
Z3OnlMzYiNTbG4DNtpaaHWOF6C1ZcpZaMxg6JA0ZIcSPls5SVALLcDt5FUbDAqBNYpV4JoWo+qsc
FnhESB/fKp4TYpfMu8ZebNdGwLZE/v7NBBWsur4E5vgpE96o2V2PrhB/yUkeOaYd/sqFfOVAPPYH
mOxmomWznEckwZ7yWdfaca/+EES9Dh2xe5bnww==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
D5raxCdsBjNBeucgp+JNk0QydQuZbfT0hk9FPoXi6WfKMKGXanrHw+M0M2EvNOZMUencxzfv6CtL
nCmVqYCrBCTP3KURzHM5DqNYzQyp0kj6XGMA+Q1QHtCCtnTEsuFMkRdychCBXeOcnfn0sPqhPAb+
dDkLPxvSvOkSf8WjYwI=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
KE84+0MQOal9OYCn+WiAXywM19zQ4xYNV40iodnIlowR+vSp+kbADs/ClNTsY+01AbPMnO8ZTgZN
CGRjsRjKcpFcdHcCbRqcEDPJE7OK/v9PEqPDH9NFgGw1pSJUkP9IpUNC9/uKTepjTRYkaMQQIcwb
MA905J1RyQ1JTo8+T7ZjypavwIpWqfh9+/OtTNQBqe8xPN3IUu4u+7M4P7P5w0QOtT0XGFUOVu4C
5WyMVCFrGwdZoGJ0XcMR+keGC+lH3zgKGf7XDuZwC5nPj50Jr/CWT4G590JXwyjmGrh+LuEInmJ7
dRdHoyo/UrKvxi9s4oal4X1UmgumWAW7Jj7wfA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5824)
`protect data_block
MrM8eXEOEx8dwUvU3OwFf+bjjcI1LBHFpEX+2Z4mmrmRBM5pwtW3267C47UwgFmHJl/vB1ppyqJb
RUUdb+qf14pdM29kBzxhcNFFOLFIIvkUe8FCgdn1M+Sj1W7Att+kvl9MYk+bxDoDZRSXN89TIqjC
Mkx2VLlbA1jUmlIZwtCBuSzRkrqXSTrZKUy1yqiX2iwRibAojYh8tg9I7UvfyEglMmRTZogTc5NU
EsE5cf13FOQxhJ7GKsFbELLDdqaiXmOcPCymHeQNnEfzPICSSlnwpV2++eNuV7/u6XX3CF5cTdPe
iij+YlTBj4OGvmKEF/S9Y2GKKUiFXwVc3eKU2ck3MOcDR36YTobO2806IJY+5ZZAXbXoY1g6bzSE
C+qlUvTvfhdVgWpqCQnSYI/Pl+SpB4xSYn4oRBuM2nxPuR/kwMqB1rayAX9PzsDEk4jDe5s0Mngf
47T6FF3KyUDXnTPhO45G6dJ5w9gZrVi285V7DkGd5ipglumOb2uXlveeSH7KiAW1CJggHyZD2rci
IAdjQH3JEWcAtuphTVEPFsZAz2Pf0o2HmO1OtUfU67A7etYbP6hujoxJpIokLMMe/F6zFmZfjE/M
jtv+6ig7blqtBd3pWsMBJPbJ+BUzKbvDSZvpX+n7WXhM0JBZj3AxWtylAf2GKrThrkX/96rB2hAP
rb0QlbT3kzagucoojVlf31pp+bgPLdlULeAtLRrqO2sWLEjfK32kVoNxgB3owJnpEBrI1t7cLdAO
L3FL0KSJPYgoR1uNNWk6em+fKi+EQxCQcleHVeb+yp8B7Te3D/DUn8B9qEfKb0r5dscCA5no5OdD
z2FUEUgV7bvwZvaHqqPt+incltPa5jCjeDDjRtf2LioFV8V8MLBv0jO6XlwuMXyLtyoT0LumCaot
BBW8ITo4QPT8ckjGsI+OwiMEmoapmcPQA0hzzOCKd7a5J18e8HHlbdIywjl/AVZPw5ttICvCNDx3
ADVYHMmrzt3ZqQdAjEI+Qnff8UwRSmHq/kFX35vJztnbdbK8pfQ65Ld1lAbs6XntUnUSwVbmd0aO
ptujnpZateKjJnYc7VV2ZcI/GApoPlPkVUhOM8bjmhzehNO+IJ+K/WGud31o6qZwuCfZjlsY2g/f
t/J28xTZ1L3iLniqQRLhEEScc+UTXqBpQOcuHzZAi96e9nPADHC+f9jf49Cebs/uuy7ZcabEGvg6
Yntsw2znwfNzvh48fkuawnqSprDiYzSxDbSJRigGete5ByJ1pdPqW/lqrruikQxJElrJ6cswEJjJ
XJnCww9IXOOEJt7HFTDfqzFixng/1LoR8/GkeqzZm7cynDv3wVRNKABY7qQVWyOl3zJStgmuqviK
F1PoUCtkv2eBEdtnrzOX7sbwQSnZxp2zhwX9Tkhtkm0X8qRIEzpjq0NDHWDSgmDHl8k4CbrU9BQ/
kH/inz1Z5QT+f54SdCTttSyQOjtLEFXxCEJRlTptD7mxU5E33S0K5fvz9SZc9GVK0UhPQE3iTvOF
xneJ/M7e7MYRoRiVlFcqhO0DuW9XFR7lCWz1gIw4uhhZ9T8QPVuZJUMmzqhYrQY/IoChHMqxI+QY
ld7k6/Vl4dH+qK/yHdEcMbVArYexM+bDQSTwWDNhD45FV3qXEtd/DqQNBMfoHYQ0l0/5L5vA57xg
Rbtuf4IW+AJ4qVojGWGFz9NeJnaLv1MyR6eX9BqgXmAtUPH50NAdcDdlM6Hpfba/ONBr48nYJMPZ
jARWOTGgODP8SUQE2uoeC+SBzBjdnc/NoJyOnVRlA/oRiiVzxm0tTx4pg9uMOgrjjQYzKXy+DiYn
k4FboG8YlqmEiOgGIVlzFliwbY9NWVC7rE3PYtIQcjoGPiMhzjIG098k9grYQO2l4h+FN68zaaeK
x8MHol3OIodCLawz8imcKRojEkXJZQKS3ok59vSW/lzjI2yD5gjKikSZ0IxjiEUPWDf4JmfcQ4GF
ZPdSqEthGIoCunVosNzWTIe+Hs6BKL/AwarX8JyV9au73C06Hm92P7YS1KNmMEY3GIeD3B13OqdQ
oDTsbqKDhZv1R6AmCnc5+ArwcflVVMbV4Hk8pLgEm02UXYav0in3aEiKeJEUgCfdVrdYk8oQEaL+
f7Qr0tm3gv3SasXxzV8RrEyAdVQ/s+ll5bbe3MOe/0sm2gtg2Dx08CqduyKTkbeHBF9VPzBWQRKo
+CuMH7tSS7VOXZxE4kkBFFU4sg/IrbH3+hC34o+1bscyTPtdPl5Y1r9XpwBMXhIkZYou16bPGzkZ
UskTRaegGKHxdsB4ECCs9uSgwNQS6MT03TMQ4u0E/iF4yH56Hic1vIUp/UWscNC/SoF6YjuCFEeS
h2GpBMEekSiUmNhzQzH/EX9xtjyQzOzTxcu9MW5447HgqpdCe7LFvit4J9vDdJzpUmC1CU5yMYkp
S/pQVzPFEikGUCDnWkGqDI6os+1icF1giYNWZ5uLBCgVW0/GP4KEatsVWfZYpE7dxMO2z/4frrDe
5bT0FO36rvvqaPJNwbX98l/FmnjSBa8zTLYLdwHaOxdhkDUGp2wKZ4Fb8orbM9lUxh1nSLKGoPMn
rCKzGZJHonD+fKHUp6dCVMZNuRhRMwNkbregVfQmn6m1YDnTaPFapGRfx4HNeGHmkee8/4EUGaRD
sG+go47efbzVyT/zk7aRNNmPqFfSpG53m2wwbSOS2MFKbTrJN5WFaanegmbxWEO0hYg6krrYvOdX
Ei0qCB8JC6xHbJGJ8HbUrGpSZ8jWfxje2PzWfRkvfFl5vcp0bkirH37bUJ97bzMMAxeiN0/QT0aM
xQ7VRagPQu/ZdunRW17cksVJWdJ0KzyBr1/lPnX34f39RCxzz4hJPYfyOop/RYBwGslrY/Y8O4/J
cBnGYQNWQCWqUwpyT6oLdUh9w52C8JyQ+QOFuBRrvbKa/Q3zpV9ZOGEf77quK6TllrGA+7qZUYOc
6XwgmP1aPUoO3zf0wvnRigyYsdifyOnzuTAiQVzvQsJPLA3U9wLarsguVvy5rg4v8VDtIXRb/9z1
iN0Y6L41uzHwDU14bCmpkGFD/4syvsHQYE3Yfl6FMtD7udnPKt2RJVuxleWzLRw0nzY/ho0+gGks
GPNyyRQ0IfvQk33coOdn7h2hIVoSTirKnxUVNZruRiHuiY76LgWRm0ngTgkL+0L71HFiqZPj+lHX
27yJspkks18+KMaINIZ2yX4EuUcjl8CNLxeaNQGlUg678CmZp8b062VF1fQoGzqmrjV49mWOh27n
nR8E3uWpntV5PGaJaFDJHlo2+qMd/3Wp7bhhRhBj8z0uE8znk7iIp+5srtBE0pKbCZOour/E5eCI
KSIKe5fRdKDTV67pGG29dBkyhA6I/gxX8EtvzBzZmRO8XPRSHncr/Ep3HHbsjRMd0/BjS6GVzMg7
6XhnRokanfRLnJjBCgd7w43E75Gj5WuPN1RDh5t1dppEtnEjIS5X6r2vgUrPDT8wBWlMju0F6rn9
PVJ1wQfBWYTjck+6Ue1acZtcg6tdhjtp9p/A7IgM9zaclzGGwywK2mtENE1D3dnRGtpkla8UzJ5l
SEnvVKL0CHPCO8t0SRlE++96/0G5tnhLdv/rbR+Fxz6QsH4tjbUEezNZlvbrvxOahM+MHk+QPLmi
04ER9NubUYK0+7kyvDXzksmPRKZHRxZQt/2Sr8Dxq4fQjPG9fPzRhacFqOW9XGw3MyFMM+6rKdih
KGr/HUwhkYQykEaC8e5TVfWChB7OZWKZx6CS8RsMBet6fiXuD2PPV/CTN5brbu39OgKgRL2CJ+Up
qf4qYLBvfnb51jcvQIh9f8WFNLzmRCDdokj1WNIoqkZE9YB0uvLZtS695EWf1d1PoCwAniV8BFq6
wrNErfEAik3derjNE8mwvFRkKnuM2RR11kGdF0hzLI4kZIW1H8/I1Gf/vwH6d0SFYo2gfkZGfAGN
xtMn9w/mKUj+i2QAQQ0dw7zJH1sV4bTiSKx13gM8/BxmlikDp73F9xWJ0Jq870mLQ97OP1gIX3UJ
6Sm5CeyDlV58HFBS4SbDlHMP/bu3+NrG2ie/5u8iGn0fjMEWFDYdiI0GTAOsb0TSueWEGQTEJmIM
ef268B/3Na5PUJiDsU2A9w8YiZkhbhKLn+mqe/dZe9evZz+J1iJVIdK7Lfk5FYCA0eEbxz8U1h35
/PapfhjHVYeKT7uMvP+T3+KKv+npRvidyJmxhJ8+al4Difkqv4rJs0pjvOjTpNfqWuXl8+VDN47l
GMnFr0pOv8Z2MXzJdYikaAR+qL5zDfwdCweITfnWntfWBEErSuHOIV0i2HKYKzpPSfsDduH7qb4H
OTAj4+1lp2k+Poph3jjJdN8rTpwAt4x/Sf0eZkN6yIEo0TzoYJpmWElnH88B2nly5/sjVpVZ+FB0
6YlOL3KmfUKcfc+AThlRIIEWsIKncWSgWUZs/6B+84Y7zqy+2ZacSyyoURUfsZCyVSMzwr5zTClh
yBf3qDI3UPjHPR1KZEXx0OZ6dv2h7QS36W4NiQV5PUBXAAFnaguPUJsgtyCH5f89pi/BEBFLo80z
UtMa2GP5PbLPH5W4Tldr20rgoEkuUog73pTPZOEcd2LOc0R9576R7nimJ/5Dp7STqae7qHf9bpnX
PDVt35sEHfFJ3eLzzeE7sJAldqxxRN9+jhV3giEaP2BdHwDeFLgCXNey64/Trt2fM7PPxSw6Xtzk
C9q3mFD2FL71GOg5s3SFYdAMMBpUXy9zpYeDSA6vu896LX2EqFl9wNFNxZdHQrv9X9NJ2GnTV3lh
/MBlIz1l51ERjAOrvT+22BDK8LaWg00sqHsoKAUGEABLa1u4kRdh5fI06Rafcs3X87Th82tDGeEG
k7+P9+g3rKXDM0yq6gnvbe0Rn4JbZwNHmg5+CvUgPw/inway0p5gu9v3EefabEaItLsxayMgbW8o
9unMM2TYZlbhE8Eu8dZxA3YHETvhGuqmQtkdM9/DLpLQ4FeV7a0RAr25oKcVALU+82hZn5LzRAIK
ZFOvShTQAOTtHbC6FyqJ/0Lgd2BgkATTN+Zdc6eh7DPql9HHTIju4S4KOWoy8rkpdSFu1ZUQ/KID
tCU9Jvc2Q6wF5HMjD3Gms+7Hb45UzLti51NzLMCB6PCH8LFsBeTRiTdKE2VC1TTEZIfT0hFsDnxa
X84KWbHrkzned8yYgx7FG33WHLjH03BTZd85wEOCxPXLcMk44yRkaRwpHLSe2tRAmkuE6R9Q3Wfl
I53RaqxIMfPiIX5VHBa3dknuKOHhmHtvBLZGiWoodkZgFdh7Bd46765zlnGFYWDrUHfVN8L1ARru
nfXhbr/0CDAIB88A3eeQ/7zPighUedxwFMGuhZRjv4e/lccCBfzUYMpO66W6dpO3rSx0gCBGdtip
Kr1KSM31f2u41Tw+T1KQb641AutwQMj9VornwWKY3AI5bO5u/01F9u2b2MebY1lUO35LhzKjzS0g
YvrAPaAhUUJqfZ14hB8HtzNyQ2y42Lj/sKgF0VbU3uTpCgoq56aFX3Na38j9QcLnGTXdqpEw1Aae
lwiU0RXiUPIFBD+Kh2ZqLfLfDp8/gjBo6/G7sn4GnRZYPfitI6u4Y9WqvHxlakPjWUWVPhR6XYlx
uVU8OEVU9oCaZyEay3Kv+/VDnnus0PdB6dgann3mx2Zxq9qITVnCQ4EGqXJcl8k1l98YPf2i4b6i
vwppskJt/RIIFU63X8/q8bMrn9b1Jd70P5XO3aInC/TK0kMOYKdVV5VFm3nbZGDfhJopNjXTNddm
DqO4B+NyJP5HbJvEtjzC52T+wenAFvcbEDXjlCt44XLc0yUqQwxHhpqSOgW7CLSFogPS+qNIiyV3
WUMzY3BsSNOQbuzr5EmZY4009nm7tmkGonlsQd0wYcFR11NvqMBwkM5IXseUxqmZw5Zb3o4A12tJ
7B0jI+CmBejZ2yZhayJAy3SB3rXc1dFs0lMvZpv/Fp0OV1PUApH4+AiWKbcHW1msBr8xJdEkgIPX
AnP5wzCtndNjsjI3s7gZX3kCq5KXhsOv9uIR+FgueMqmIZNVqnwH43G84ZH5/3WRAfGmEuOEhjjC
V/gn3+o7sptr9uJwGYaVunwlmuiEDqgc35wj/DEiKD6BZdZYJ6i3twIgSPzIt6Pbg/PIg5+5bapi
TVWVb3PYOhQUslCtFQlXPzFkFb3TPVdyhfk/KFqGG8YNFfCT/hGg3qMf4rNP5fKxv764KzuWmqr8
ao8MTh+Rc5hUWCX0xYFhz5YvOe1Si0+zzOUBLvAWGk0cfcyi9gOASwgQMYeBadUW+hlPmfY6Z0Dw
kbul7c9A1gBqA8dGT9/XLP9KoNyiGYw3dPOILM7MRT9FLvGgKg0osWMIelRw81oIRW3mZ8zN5W6c
EZ1Wllz35kX2D5NJiEAAVP+4T8gEw4hrWXv/Kim6F27MnHP41JbKP9ILtGudfklMTQe8Bw8IaBZ2
jgngYu7kAosMg0TSXy/AqZZpzsVTF/O13lEo0jl0P/3mnMZkTkKrXanKWQFH6APY+9mhiQSVDC2H
nz85zp1i9D9hPc8nTDVLcOxhY7Z1VNOGCEamaaQFv09WtHwOMByBupmeXbpixnDIeam4xrhRryQp
8n4dPvgkPC+l0NXmgM4Dbf2tzMxu0GmpmCllYK1+ff+3qNmfBrZPQGjVGlaQRopQ4dA+YKiM24XN
x7ddmacw5SWyG6aetTr+zKd+qipxqZt98BhV6hLxvmSV2MCuZMmu1TLrrn0FrjOawSKVWoI4TLyu
eKNrFNpCW4Lm3G7134TKlCYn2nNpSfrwxbpgEXs8s+RAvXjstEDcRCkm5Po4O2SJAn8pFPtQcht7
Op/HsOkO5EzCWrbDnTuRboJWMY6Hxo71fn+B48HG807B1q29ddq7tGn2y/cOrKijMiYeISPUoxK/
eiteirQZleCDFdH9YbtTYsku/9z1HKDjPsp3hJHV041ZH39VRCzibJBhKBCfGoSbJzDExWeITOO9
rwfdua8awaUphsMIF6ft4MlUkx1x9gndVA/2y3HtBec4euRM/+Z0reb3PbGiNbHbt61LPdOoJo5o
0GaQ4mgFfSnqTdfJTJBREgjE57Dw0OsObYWPaDwFEzTfuyqlhvolZPXif4OYEKfIolxW1R68fVa1
/K3d+/Ej5TmwbH98PylGMzhQiw3cpRuRD9GZhhSPnio+8UNxuw2RogtpntdvXgmUVY2EYxx37gZZ
taQiQYNAgU6SFs1UqQiTlJookpHDGmtYsKFcHpXw2Q6l1N5ogo0JB/Y1otJTGQUTjLocz+905obf
XTUylAnGMByNKo201qwCMZ6GKBRtO8Vpn1YhP1GbFWp46fu6Hss+Cz2xw+UYSFSQ4isyMeZiLKDm
B7xceWbo8L87dlOXBJRHDoUhYgECBkF3+phKqyvlj/X4cB+Jklylg3a+ILHD9YlpvGpVBi/hVKAG
SYntrAkXvoBkU1Xm1XJ4af6Rfd4Vt8o3en5W7mOGefADASbZasv5oritpf0BhJaYbaqvM53JhQLt
xzYxpnFRwizU9S7HZ7iLJvrb/azQNkqWv3bYQCNsACLJuX0NChTcyCyCETR82kpD+NzPqS3+WiA1
dqbHkwQv0kHr9D570uahsaErEpD/0FTmnXgN0nYFe2xP2rR50wNaaKVESWbBzfJkIULCPWoLyTk2
nfAPTjrhnlDkyfjEOpMYVvaAj6quBQUiF+RNKmnyLbB+Np0gusfnSIykv6sz4zGTu2YVM97FYSt5
KQgh4e+E5/P/tA==
`protect end_protected

