

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Ksr82/EJdyTi/ZnocplaChIHl5gVfg/QywOs6WHQUUTVobYB9S2t7HfNHkvfksORtftr4wgSGG59
dqflxrTk9g==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Qqej7lC/8l20xFx7bklclhPhbKpE2SoVMnU8o5jHyjJozBFHGWWzSqcy2OHoxuRC4svtWcuXPZER
AveySsBsquyvS3CpwUhQC4HU879mrvq1rktu6YiGUKekxqqq8XWVjGU2RErpRUag/ydvNbNrFWxX
vuxu46YvGNDVpOq465c=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
439mpd6b2KugK1Dxw8VAcq35Q01RTqPVrzIbAJdjxQbya32eEZ7i4WNiFuVZ/MAk52bZBtBQiNHc
mNfbIfQciIHmnAXJEN9w/4VODhRIcUMrMjQwAjn4teKfB1tg762rR2jvGQ50Ai1Ml+OYADsAGJtF
URFceTs0yqpLMxJ8Ov/lGmeNw5dXmLiwn/XRqtS/K35VTjZyDUeHpQAr9q51KY6k59LrSFC7lxxB
mXX0In+fzXXlrh0dFFwLWzscDXHiKjrU4bwWBuzmrkKr3uCoEG0OADwjka6wlXo/Z2cEkTpiK1Qy
MmZH9UXQxrxTgtpOMmK0pjs+MfXf5/7XzeJsOg==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
porEUqarzWQ+a43o1KcgcLOOq13cwiYUyYcVmnYhbdWCiVlWWfN80U7oRzW3NODV8vTOFdEeX0/T
HiPsKQYOSEqQjf71FVXt5Qu85a7gangJ+zMjyuk8+m1c85rFqWapoLbPUbexfLeiEmybpwcybBzj
rIVwXl1qRv1R4JNRI44=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
s6/C7NZuQyYs48nVSWrZBvdUw/cGGwVNCnxc6+Wr+hB+GSdh07xJnxht3+mpM71wbe2jyi3JRq7M
A8Qq9KlqvpjZ87ZnAxTvr8P4OZV0DRnim60u79JqHUDowRtwBKuWK+fhBBqVkg+I/GuK0CQAje2N
3H5CzXagxYQGmhNBvdIDYAmWiG6ymENT9OP+fdf/JngSq3sbaQDhuOCrSGCgAWuZWv28vEMvXd4d
VKm66HgH4TXtJpDsYN5kTW6gEWdi7cV3KJRDsY6jA9RzwyOOBsMl8Gl/UvSGBWbIshxBeydyVUyg
0jabYqp6ODPXSowz5ZkW1y4reTS+cozycJAuMQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 11008)
`protect data_block
X2Hy31MD4zQ8xzUd/k/NB0PwPB3idSFzgWygCaDOLASvsT/VUtzMEdQuvdE0zkCfvPoH4t6nSW7X
U1xsvQimrMDjnq0ojAodHUtriY3fzV7Gdk8LUKWTh4QHwt0WlYolgQsE5n2w97Xp7/HSeD3cT6Zj
oUEcRfNRmUiJEWJxTwVmYKy4K+lrBtnRAMLspFG6MZjyU8STN/tcFt/qKMdxYXqwW1IukxJA/7wa
5pw+Zw5rHbAX2wPprrvNjfz5bGJWYD/Ao+/DXlLbTM20gNYXILWa/xVHpq0kBQHd0NNI5B4vgmK3
KBWoDsVztNKKpHyH4vGAdvKQhcOYmHSr9ZEOL5dQ6HfYk7X2M2BU0gpE6jf1NeHzdlXvfns+/lmt
vG6WITQzl2MzLdr/fsKHDpHt7Hm7DJM2+3kOpoYZJqAQ7gyGdLakil9/RiglTjjv9og6LZ25akrP
PQFkPdZtVuZDYPLYtnczJRuUzJsX5aSaa49blEh49ygqXcBQ4Xzmxy/rYGEUa8sf9azO6+oNRbsu
zFjL+lY+oJCKPln4gxXux9fFD9MDlL00X2k5YedP5jagXxjCD9Rk3YWozB5d1ufcoVy2Fjkydrqd
PG3eh8p7M3LowxgBCG1e7HZPR6s2NgeN9WF+7rzkdnmrsV6wLFUPLI/iZWL4vFOvcpp/KwgThWhZ
uE+j28uYxiRGedMIojrUfcUNs2THTYDALNOBQR+jXMBWUhyiXG8oW2lNm6PaYvOySY7xgLfvLWkJ
7g3IGCcfXkxwFcpSTi+O8KRUgqg3a3Z39hMO4pWmwYD0bzDYmDNfP0hpddlAgCPtplSmzHFJT7Ft
dwMn79b/74kZHgGqy5v3KUMTnfd4klgEZODEK7He6uIA1wK5pvYdxuqMkva+YDK+OB6Go+sZ2cGv
qr9wF3nhoqgyftUWzZczLMbjwLCcmHXAlCeLxpRTw6j8SVJ0fm0QBWZnvgDI5bl45zNrzwMpeSHx
TuQ4YIn2Kbc36j2XoNA8+9ij5n//YEYV1wP1Nxhvt4iB88BLWvXslnQ3rFsTmQfs9rbroodvWfqD
d15hNl362eMJofsxTpSva6wBHzutt6pDG6gPJpjWOZJIZhwXDBEC9QtQEjWhyLB/7CnHZH/JwQ25
Ay7lNwmhnT+EnFYhUGQH8blJ+RhQ8UlNocRrwCnAVGKvqZMKIRRbiq4A5LVyprATbfcVnahq4FVr
U7ngUsz7sD6h+VEZpKxriBPMGV6Yoa0HolcLil2QOGxOKNqJNo2PJ1ezcIW++VaHQ2fk7IDra7Sf
qg9dq5VmKku/SjaWAa/+QbnQr87P7jWc/bKlpo/6OZ5Z0dqY5nE1YlQPsCW/WaHOfwPNCn0UpR65
9lKziv8wq6YIk4lt28AwGid6d29X6OrGaudhNHcVgo0oEFsxEfH3WnaHf+/8QWI0Wh/9/PtIilRY
QHl8NBPd+HqUZexVSq0GJ73pQiIu4S0cRdgccI/JAJNDItKO4WUFC4rGlhZxO/OAPuE0A8cTo73n
RLuhC61odR3CuBAD1aVcgvDTCUUPb+7fiDBmmmROZOJcZyfjSQAn66I2LdvghLcFMsI/Mb/yW4fa
4mV2dSdy18C0F7vxW02nj4jswFaKb+7/ZV0etC+YJzxArlfhDtkG19fukZAcJnO8BRhID/nwqAv2
LYT+Vs4PsHEuE9iFBn07YW18QNe6gOadr0ZxhI9ZSq8R5pDaw1bTCcOrODm/pgFE064Cp29in6Zx
WCABWviPM5fhkdHujqBihK1yr9dM7Y3CR+2FqV8fY9dHJWrXNThvQ4bkilY4T3qrd5a1yZs+CXR+
YkW3UbJ+U6dKXjbnCXV0jjcIF/6vHeebCSbBGAOmYwsXYMey7OshUQr+CC5ldr6hp2vdK7T/S+lD
oJNRgAExpGmUcwE3slOGoqbJ/XfVOhLRgwsH8J+UmtJL1oi9jMheS9oEse08QX3qfO3fI3U9EPE8
mN7KqrN4GIL+cxsfe+qp0mEt0hjXowqCq9NpyBz6I5ultzL3FpOAsSQAbTtHbIe0RfJ84PjfJRYq
9xSk57zx8Vvv/coITgMoQeL3OUH+pjKGqS6quHk+MMHSLnJUxRhPArAEVwybRRJS6EhNBwydUzPH
RqQQIbc/irK+RdAn3j0oGSzIVGW9U/6lUD62Z6XH/7hxcqsawP4AYCpqR7Y8H9wuoo8bUs+c5DHR
7QHO2sLAKK4kZGuovNXk6JYPGCsXbnZQb9oVBaaXk/pAffFikzGN1JQWnftCnTa1Du8pr2HZKn/9
qqY2VEZWSoyawOnPI4FFpMREiGiJlCEuHX3f8qv1xGTPsnHIuG6wBxEEoa5YuoAze9S2k2Sf9ryy
Iyya/x+YKBzV/r2elLim8SxXzYmbwG2jQsrRuHYeig78rhfQ0FoBo71mPe5fVp2EA+VYNEHypDSu
H1W2EdPDowByFjsii9/qlZelbmPTfrmjXWQsAwWIZ8NPuUpgsMeaDuKm4f7ttc/0Im+X1dwsuMTS
AHF7Iu26ffGdU17nvXhU7wAySbscyoRV7hYr1mfI3Se5YklA51MlwInk3wrQWoxDNRmNdkoB2IaL
a6Y9zqC5ECcZxswL/VK9R5IZKFG65Fa/IVmzT8OTAaWfefCLV3dX+SmfZkr44K6IjwsR1SHgkybg
I/QmJLbx+9bfXpvBoFzMSJEwbpF/kVKG+THjUCDPRPgqpr5c9ursuLnoOG4poGSRfsv5TjtMAl3A
cQTd14cZfZec9YhrF7awv3QycA4eCVkwbuLDT2kxKZK4uNgHSQTYuSzWsQXZO18ebhsbvmhjy1aO
j5lICHPTGbdzOqYID7N1NuESAEVw9hkRmrZcL+wAnfR5X6TUwQ9NmsH1JaxybrVhKlUb2rf/+c0S
nMcCaTmA4kE+WuORkKrDVkxADWyDRssCkkvu2C5TGxvCsnNqj5iTtqIOPDZRhKHX/f3SVUAmpBN2
o9dtPv5Me8/LkY0WDu6WVmQg70Elm0HFsTr4Lz0Ov2dVdTEJkQdkpOAaimm7SvZ4RD8asAtLAKlI
5xqSMZSp+QORvrIJPWsauTlpUrbifAcK3pT5ZwD/zwSR9jaZSyesEAxaez9lOtwaiht2YPxZ+nKX
zbNTwvjVoCPAIXf6ezWp4NG3e9Ck6t8mEokuDn2OQN9NC/bifuddgnE4ZrQG4O7yiRoGRn3zxyfQ
Vp8F0GvXA4T6gsM7aIK4UKab0bzGz4Bj0Y5HpvcNieTdOi1O/lvPrXpn9MhgvlpTyJHPpzy40m2b
4KzOZ1xjA+amsQ9P/t9nfTRJ6JQa5RvREXVIDinePEyh1kDzr73VIJMwlmwIsHDUxNbl4X3RIrkX
Wr8wtcsNPcbjH2noDVQq/pvq3GWzimSamU22mMj3HjJpPdCZ/+IHL+U61baUvEPbfiB4ZDOipnc+
4FKM21SWCXSIngLJtTIBqaknWQ1HRnuuE11ArMdkZNh+dB+IT6ES9jRrSbBmy9iHkV+Mb6sBmd3u
TISiaLovCkkp956dG7dyqnZZ9D16gtxlhBOpB91jDvCEaRVi4KMF0YOh35yfXefWuXR0zs3oZ9/L
Irn22xkvcsMZnv52yy/YEZmUqgm+okhC7nw5tZhZHbfiAa5zrbPVPYZbMp5fctjfwPgYpJSiJm2Q
CL6+MAv/npjxMuYVP2oaUByStJWRzFiOZ/A4/Z3aBBIpb9KzZBYplv4YC16xYIXZa801g5xQuU+/
yxwo5cCvDOzwlmnqLp14qN7zL7V4oOmykrm23YJfq2Ni4s79im1cZserZBvCkGeMxb8ZRImAJwo4
+3ZDZ64h85cphODF9cZgYoUlCpLOFgPKY4OyBDmmxDhMdR+6UtfZ5hy8V9Bg6MSoor3cVh4W5qSl
JcQ2FUsGnbzwkP3lpdUuJbVUZ+UqE5FxsRqORvoyGGvMGa8/jRMp7dzvzl252fSrkEjkZPIJ8im6
w2C/W4wZwEt53kMqUzbINPm5MC7vS0mCGAFFI9gOrjeKp7LZa/d4fgJbpnFp+rVOY3eQgCC5PJbg
4pmroDSctjqHrtaCwme1tgNz5GcT3y9vkMsVTogABKxMunyxaAAcQ/W/hQVnxlVy6IoD7yIOw6pu
AjX66Wfh6a+kPRqiuEgzlhEoH1ygZtxp9dEmOWEfXiR2sn8iqQFEzYtDtPmyxtAc3bZ+ND5dny3k
nVaPnVLXNdGVrpEoeYte4ZMFioPuSLo74LKU+uJxvPP0oIhwqD1LdHWF97oWttvhF/xmbmXx8JL5
5jJ2/DSpdiGHDOlS3VcltV4a1VldXXyNQAegSZeFRcPpva9wTvlK/ZBoSNdkg/2YRUrCSODIlG9b
zZNp4F5qWQI9iVld+2nyjr7TdvRhXvqKuNcpCjyi60pNdrgbmYAmxAuWoKywVxZ4NuS+aXy2K9bS
sJF7VKaiQ/f211lxKBfoxiRibRNUvhVKoJRMoARj1miTfBJKXaITxoNtjFpA9+6nt9pielcUugLa
1V2WKXUp23PeUIfglrl1YMXW+GU5TAmivZc7RdFy7Ij1uQNbZtOTT0cWedIcsVb06EJXUO9AsOmI
xFzpmxs6wrFEolo00F77vtGKsCb35GM145DYqg+ABlLtW+ndjnMXJiXtQ7Kfw+64S6/nQzpoYOby
F/JSXD1r14VL1170xlJA6jj1Vsq+T2ZeDm+pB3Yo+Z0d7rFrhcxXA5QwYVS+wtBUJuljsQ94KMxY
uou30B8d+5lUR87kY1xocwUWB5hLNN5Z/wgId0zQAEUMyNSzKWXJ21JDhgw1HMiLsxD6VDbV5ZJF
unB7za/fSdvWqoXYCkDBmpDlXIqhB1129yPugh9J7o4YD56ANjYfBt45GqumaPwQT37oaVPZa411
qe0PFRC6uF4ReKy4v5g8muZcxwktPDVUiLqYLtltTDIUZWYeQGMYo09+eNEdrauctbkween8WhPb
SP+YZ00kagMJGwq8ugZZZRe78POcKxci3UkpHDBgM+uZzKlBuJuayrMZRjMupr+S+jiFizlre3Oo
HyXhnwVRq3sNrtcGxEw9IxjK8mLhjd3AYAFZTvbe0uHOYZyat/HKgPW5mAQUW+sptrVIOfy38ySS
Pv613Ddv2CEoa4Hy7HQo7SQs6AxM/Xkgj1riiyvMMaglI+OXGqbj5OMUsYxerkVv7+cD6A50kngL
84Ig3lzoTJ9comsSmuM6vvGBSV2slP0EBKw/vA4dSbLxnbJDdcECDIgSWYPAB3WkyHlezXra+ZCF
C/+cgPF6XQQ7Mv82l7iS2NCOQZT7srTKupV0R0uS32wHamB9aomEpRKRk/SaZ+JioMvEdA0z34gj
DVXlYLUI2h8MEu+yhcuFPmQXB133M4kS/rgsnc73I+GpTs6GqdKzBVe75qpb/k/vkO5KZ99/YNwN
qj6hEDZG7XccQB/Hp0UsFVzlMiTMzFgC+hfAb03SchZaQSalVfb8QaDb7U0pa+UGlhGqulGPQj/n
DfEXrfehv4/8xpEF0ldFibbD/xDXH8z5SEpzy7aEveup20T2hSBLUrj3sUY2f9KM98hlrkrLP/Vw
uqY0uS4OoKhwRGppAPRMFOqJNGVzY6oPoJCcbRxXYwO/wKtYbOPSJwGgdPLDbvjA4YjR4bsL+KVg
Yu2yJeHpT8DCgT+w3uW3VoJ9tFnz5SzQqvdPNr/zPndpTNqBx4SLPSfM1tIbbk6htvm4Q+tkfE5e
jQAPVhAdvJIrlYAplJazlqLuMhOfNQfQKeJ4kd77HpQC3artzvKVuKSyeMYNybiPGoQtI87Io/6c
CCqSV2V1K3/jhzsKxPt/kg3hMlBst8BV0QJUPTHruGE1+ytl9PRKxjaNLG9VeauQi8U7kk5uZG43
klq/vQcS7oECXjIq2rVJoDHkl1KIsgh50NlGncATyZ3V/zhxk1kQ7tUxheAeHBYtziAXR5/sGeR7
dtFCBdxDmC5a4zSJ0niD61CP3HxmwhV7z9xrYjIzfgPY77I9uxMHcrGvdF/fRCfny+JshXxDmIYb
q1IggIKDoWri6rDAMKqvBlZ6cA8kALwWIFSTAByYpCNzsjKCxuMbcRLUvDAbUnPbF0Q8AAvUKzHO
HfwPiliyCZ8OOZX0aqRIoDMugloqHaQU5r4306qkxi/u3QgQGQDh0O16N5SIMXhQaEErSQsMJtmd
KaUFSab+W2XvBwdBwuJLOQzxoi45RYzghlJ5Rhto3AF2xqzfVo7ESeLT01u2VIaqxJcb9ms6w/QE
b8JngaoYJHdwMtQx73r3qTBTrXRg3YhqYiHuyk4bEd9J0CJ8rquNVdK8JdNiqNQBjpD1dbhplnW1
prTTVstX0V0rB1nkEMkqqhK/Ptnt9D5UXMlICuOYgtpyIUhLJis+YRGvhA4JQc4fqyeQoPCTSkVa
DvEvMZiI2f7VjTQUh5mcM2ZjNNCn5xouW1viNZQQ+kz8Lbv8UvJr9KQi48J8g/IvkQfWhq2mbf0g
G9bsRC2P+oRmDphJbSabph94hJIVm/s6QjmfenVl5WgFfAqtLhSJIC7sbqStEFtQKhUj4p0Lvbvw
AE0JWmij+5idTTqSxhM8T+Q+67A68JBtGIvoklxbRHWhCSTsUEYh0vxLBwlRQahM6kBGwOfSxI9C
QOJ5PBIN1ST+oEn6Q+Vowdgrgpw22mMlYhvEzQ6m3tmvGjYWUqYZfyw+STO6cdQrixmsANlFde/c
Xl4izpyIL5vXJhdyKNx7NbRc+uER9gZiCDMiQsSmvdIKJS02qg+eTVeMOOdyUPWhuzONK86V0Yz1
KfcqeybqKwSytt/qAVgDMK646vIiW5Dl04plQVedypR7zXON9VcZnH2AFFQybE13oKer07ZIvsz3
FCqeuYsk3N+Y4+bq/BBhLgVXFhbcnCQ3jn0+E3aKYAt5Gvw0hbBJvUWfKlJi3QP+XhhOvEKHo/nm
1Yrc8Qy9lHwa4UXtNxe1NGsXHx/3eK90lhlmZKN5ej2gWC0h2kW1pN6JEbSz7VFPJrb5GkmpickI
lxGxb9h9upFRZ2QM/u+HDJJeYoVaUwu1ChxxsxmWvMuSLvn1hUemLFeMJDT5PW/mRbYTUqbMCVzB
TH4BaYwoptNamJU1wQmgZFvYVIpcTq1ESygbNoTUkh51VogcJqXpaOYtqEvQ9qTcr7LBov3K7WyO
9wMT54Ng2v8S9k/41yUUKwKzS03yxfcz2gqxyQL3E62bKMg/zX2Fe0PPhyZCf9QbgoGIs+OxE1dQ
vICG9HoUc0u+5XskHC6+JizCnPKev8gxQNBHmkSRBkPNKJ355YzJsrezaF46txRSdRduVM66WAzp
4ww5yIyq5od9lQZ3bvxO+JazxgNcs1fLdvZQcwWLqKtlSMW5cxqH3oO4/GNhPT5XauSO5MRrsk69
dmVcKwC5aA0ItCEgqLxBpIoJjJHJ88k81s771bOShBqfWj5QTyhk7oUUywK77Ai9jDQJHQ1DH+OO
ZlyO7k9DIfjMwUj78OP8KM1Lg78ZNHPc13WMlmKARzo2YyKuElbn8YFAalF3QngFbRqFFGtTDl/+
wVzPgkJ38prAjpbkYWpyP6EXBRJ3NHTg2G+Ziva0k9fhiK+tyk7ivK8ikg37eiILA/bTYGLSYtsO
8H0CYtvYx9R0E3F0or+rnswQcMnIvU2HbXX54RvKAHgg4kr6IHcOQQ80lMoDl532zpJnT7jmUK6N
Ks0O0BNCnxcN91dyHeLjeA9t0gmorQyZ9N0cjtinJQBFiE505KbN5subO+LlGopH/VHu4YPELPqT
CNaNLnS/a9D4jd9uhu8lVhjzBpfrgKZqXHFyNMULgQPsLRN0p8OofrnajzQaEofozVcqnU66k09o
Xvw4HPaFWgYiDojPsYu9HLwMS7DOv7rLz2X4vL+HSGuXEszpvTboMLooXLI2JHqptvMaK5eETU4k
bHSmzFg5BiVuNZnX+5RlWQ4ZVYw/PcGVRVOM4I+04ltpLSJ+nGf4/I5rI4KQCWx7fn5xCkcy1DIR
0ZPhxu5ftNGBewG/pwTzQq5SISxVirj2Ty3Y6+gfnWTrL7q0RT3Wxs3h9RckgX6B5Drfcb/JJe3w
bAvIcmqjnElHUYSKVbNvsCHq3MOhA47T13+fcb2BBUYQfjm7FR0leCKqbAULTEYWX4VFXO4MEa1s
SjaD0Vl7vDxrCszl4sCIWhdEGY3l9Al6vMQuSaJQpojy23FIqmY6dw1KgquIrzB0MxkZ9SRxoxRk
RB2tv4ten9mnkpXzP77RuM/EAefbkjU7BgvlXyMUjmRqy6jyqNjnDlMET+/8ZOcGRvprEF09bQwk
6LcXgU1sRxS7ersHk4cal9jarBiniuqd002CEq4+MkbpsTZ1GmlbM33rQTmgrVk7SflJsmRhG4sa
/4cuzolBlFIMDyCV6v9ij+tEoNn/lY8N1MQL+z6Rt7FghtGpTTBNmXaGEP47Y2xfQpfyD+OZ/rXg
5RYO/Dy7f6zaVeBVMg+zrCVNwp90oBOH3/DTTjizdqOkgrdwR0tyYq+PJtUUKPv6BxNRx+lcKFE5
figMR1NWtgz8XmE5S8mqOPHKXQzmPd+/1RZYokF/kzxvNXWcYZaRIqxjFljCiz24JNeaRy75AOAn
2n6x9krj51C3IE8kDJ3um0474TrtxS0GOuHtz4txDaYaQCTn+SAt5JUbpgl02UI9KGwc3T80EZp6
uLKT2UZS+7J0A/2y2ZwY+Y+3t8qt6dJpDbR9qgNtSFjFqAXGyzLqjH9byQXJolpT1mQXhx/Btf1T
1CXrzhif6qwb9dCdUY52Q/sU25/7q41E03NCNspVuKuCcwiVDj79CCgjUA9pn3akdcfkGxVWqwAa
wp/+eVnwbNcfYlmTi1ZZjd3I06x/SABXbqzhtBTSeC6XQ3W+hKDG9M183OvwTsSX5jLcaCVhuOld
Y+Y5EaWOACcTXSmi371sd1OCrM/dpyCbciNI3aj2kgwQb5ZJ9KrzjC56u++9lvPQkrrkxZ/GwmRX
6/1S3DeH2zWJrScfz6FYkPlxPwNBPIcYlrkFtGotJzOMz3T/RXU72uOBGPexsf4fB+bQ3DkVkQCp
YSxL96pFcz5BLI4YyIFAHbx41r4B2Kg9kN139oOoFxgyd3T4c6fLI3+y5Q5bdMTuxQPK/i035CrJ
N+EgheZUOBsbwM6Fpk67SwCfBpQchTWg2deul/USVvwwTP4ptr/CdS6AaP7muCXAPWXns8NGjW/2
Dm9udpJi1f5ZOyu5odxgdSOJ2eFLMCJ9Lu706MloJyWsETRonqibAMk1SBOyXcDS8Yf1yvq/z4Jz
a0uStUnjkZ6P/97k/ez/9zlmiparPnTih1aeDRNCqDlyBLCwGHgwZzGjyF5UdUW5vff+DeEP+EMt
W0MX/5Yk2fPnddNF/s93Mah3cdYwezUR4qJScpplwAvAHk63NPnM5wKxN/2LIKFmYaq/OKMJ/8Dn
in66WBIn38es9zGpK2cPRHPTIzvYLleTTwTehqcl7Am4S7ffmQlhy4oPb1tiwF6zB//QjEW5d3X9
6p+2mb0obppqLn7J9YljG9XoMQ2jWzzmJCRsQqcM7rGL4rxDxLRlEdpxxXbEU0IRTsXHe8YzYRna
So6xpvILb2wX8PUH92gWtwfmpoSoDMdBWf5QWB99pumfDu6ReTG2JwxeQyws0NaHnNeTln6aH7Yb
aathEdg0hoaMTuAlNUrMhkGQ8lF9RjPJDOLFRaWd5ky5yhvqzIEaxfLROApqz9K9zf18PH61rX7m
LVRe7yYGkRUizdBjHFwdXxpGBxGsnFjV3ozSbL3ijJasWrq0PgH3+cgLB5dPn8cNNs35PpMKKCU3
NJBkIZX8Liad/U8uO5VYiT6AXUJ6V7MXGsfFrjadgHY9ODsdQw3YsUzjz22zzDFYbb9BuhgizqvU
LeeyeHeeODjITk8wcLYxsbaWxL+Wu/20WpratTSe6+aOM1tjK2/NJKW+HyzgYlIaLPFpHlYSP7Sb
jmgVk2NbwrRPo+g7DNrMRBdI3BpxMnRWSULk2DHTYBA5OVQ8RjBfC94RsNWVKhDqRWE6HaO7fYsp
0U41g7jp4z3zDbSw6L/HglEVkjbLu80sl1jwpieVs9ZaTI58nGVaqBTEOwz4splXTtOLK9u3sR5j
MvxNyYbUdJXHF+Vkr1YW9LNAZYUklcWxONKKs/RyobQJiuuRZQOSMz8EtTZAuuyRlO26xFab9wGq
ysSfwPiBYSKBPeravC4fql3p8Bgv0L0DOw0hsHzcHloBZoCSG0faSjUFNmhFwKdP2Vr7kWO5lCB0
aI3FsKMeElW0yvbAqqxdfGP0F/9lVmYu7H3EQW8T7OCHBWw/OfHtvDMNCTSM8sBF0fI5CNMfEY12
dkBE5ikN8VMy3HzDylSVIn6v0GBQhN8IhAtwVxE3uAMfsyPqik0IwEQm+XVV1ViOpghksBi9jotY
8Q7+KG3386OP68w3dcZwS95aKTGqRYqzvpQR5O7DqImdzGOV/3wRxrfS6L8zfZYHgle3f/icDCEh
RKsepYPYTSVNtSEh0YqptPfb/yotmy2WJlxUO1N1fbFQnWR00e/fcFI7wzscCnZ2m4PAvwW8WYu+
PrfW2fTDyDtn0ZSvgpzAh9Xy/jQwxt2oF4K5mGE/gdRDIaZs6D0BuFCidKzvf21cbJs/PBw8/GB4
Kd4F+mTaKN8LDljn1vsv5M1+OUa98gWz3utvn5yPxhtLpqlyZMuQWZBrKDzuDP7X1DPxT3AH8vcr
CtawLC8OdSORHw6sCVEqbFIymg+ofH0Sf4/otC5BTwnVDQUG4H0i0kRgpL7HC/1BqWNP43B84S6x
3oTWpaw86RNWz3c19tcFirIhBJuYIpWZ+9yOVWOrP6QmwoqROd2A7uQGcCIFHXHsKtvV3TqBSTr4
NPhi74FV9z7kk5Wsj4jFAJBs9csB7nB0IZT12leeYdGWnKh7/D1aAhCiBEC3c2n1RSc+nV8+o+2Y
QW6bs9v53V3AjbFhOSmrp6VLMcG+s05/ZpBt8KmHApTkUgY2HJV4WRHV0t6naO82a7xDA+Bl2Thr
d/Juu3GUwZw2+edu6nHK8wEzEii+WUuiE5aaeWhN/BebYR8V8a435nF5X4e81x88VIlEwbyldbaN
S9Gh3VXf3wt37oHu9YvkU6+/9X8Rk7/rEe6VDiT3xlr58gWPFBruvnumQX7CYf/n99wLRO0dAfhc
E0qfWVksRZurndwgRcZEGx9nElQbod1IHOFyoHo7ADGovLaVsHbmiD3QYY86NTSQjhwkwgLE6uob
4k6tPgxtxeuIoxSEmK24Ly5rYYeeuTe2YyZ4AmTRR0isK1p5LT5sbvzO26HxIcmFXt/TzT4aMI/P
aHHf+/LKLdguZE2PqoveDhsdRlwJe+uFHEQ7D1JD3mp6xxTXU0c2n+sh5hXyQV21tpqE37iWCCOt
Zq4VhGqCbFajF5zO4b25GdFaseXS8psON/rcPfVWAiDf8lNQffq/LuF2f7fArNUuaqYW9tDzs94d
3PiQQ/s0G3v/o17vNl2cfvueabtIityLDASweumd8pn1Y4YYs25LiHLge+RMR+lX4uIDv3cM9WPf
N5IL3VMupvkW+q3Hp0S0pF4exMIEEi199gEREWUdcyJyr0Axxw7fqX6zEt/A5TuI1qt5jnOU8iJK
lmWZCpCwTjTGppeD5MV70EeRid0pVOJeTdueIAjMDTNFJepdCwCpDeM+CXcGJXlSBadd45yKn9c1
Vw/1u0aKYo4EeHcReUhcbkdixscPBNzHZ4qIEipGxZJ0WqVvXQEqjOGiuKWfFbeKfYtiW1QCjqaL
cfNMWrAYORAUXfW82ULgsMWiUWim2QjbT7a3zND1ZllVcz/B7rVO4+TpZoC3NhJx70PgA+8gdvdd
KMd8zmLzSTg8+glcvBIiIiQYfx32PeWu3rUMkCgIr5OyAxI6cy3n5Uc1UMe7vzcOGXOlCEKBgkU/
1L70Fah+dhSiUp2f6qgAib1ryevkcIhNPySSh/DEz0IHrQ1doUjUoNadimPdtNfQktKOdNfdYhL+
oj2fpTW/QVL85a42KsvDwFeyoS6kAAzCK2QpBpA6Y2xEO+slSDWope6tnyEU7wI8rZ+N9d1MTHZ9
P+eRhefcL/oFQ36YbMjExxEAn35+Ftgnvh7FPUwLQ81zGy5+Ge5DwD4ZvD1QYhvT23LZv0tf1CtB
xTXUY67UowID6ZZzNTXsOv61jyoy3kBKE1xi9I3tQgDLK9WVXsfth0GFLt2E7A/SvIjJMxOzmqvn
cc494SsR2HWjU6xzFHpIbXVRgGBiQjRZxVeEC0gz7Mk3tWPdfTeFiMfDDdlUcBWIwJxrKrFVZlQZ
JHa044qM7VuHJSrOIkQW1TBfkhSAL7c3WXZX6chngHOlBaGGv7gP18YhFKdbhS6p2STQqZ0nEYv/
EO7gj9Pb56NYyBRp1XxW/guXrRFdXwmrHVOdagO+VMqQT4IsE4OwvOaBS+xgFoWY9kLgtpgpcYXZ
kzKU39nvX4WO8ufRPDf0YN5iSugLgmLluuc4xHq3HU7KnaVmMohKZowhPHrJ46p4cUm/ScKERyvE
FzI6dDFx/AWeBYGky7jfWoXksYbTGafum+y1esivHTZYLKV/dUAp37FPzsY28jSMHl83ttRSGPUE
11z7BZw5A7wariSazYheIGjRqQZfNCC23AJS53XSAi4EqI1pTCpmE9oHb9NDKqJhGrAFJgrG7uQX
ww6OHkdsHrwMNPWQaF8rH4lzWc5efV4/TVuMDQELF0b5mzBvugBq60CxKT/5LQg0XAyR49roOEc7
U2Ou4CstAqml1dNrGUrTKoI/i6KDSXyFvCn8KYWZX0PaU63G0iRREuTTHApaypPPsIJQRzxKxmEg
vPz3wRGfPi1P6S9z1wAzsHb4un/JurgsbEeHfObD2KrWqW0ksujwA68t798KT/U+8dLF3nYEQENG
jEzUtU9LR8kJeDSRPF4symCGrFttkdMbxRQf34sKdTH7bwdHBcMkov8LyU+8rWfuCBLBcosKY7DK
ueGSohWNxvt1ohiZ/2m5ah/DH+1kcwXBRIVVAXpKR1j8JI2EtES0GoVjReleNsziZZAM9RlaGUMx
zal8ObWgnp50zrfgOJF5YhoAZ0K+pNL5hbvZ5MW/vVHrxMXmXo71CobeEJMTlbWHy6UHul3fkRmr
VV7BzbvTg7+dbDc+ubi5eTzdyluYyhM/I3AAaBI2toyabsI3IUV/Eg3kRSzZ9N0VETmVG7Ed9cA1
jWsJWiYsTQY082LlHoH7UoLVtVz5N8NbNpq/MhSntB0Z73E2OxNGphTvGdOfoheuFQpF9iuWQ/h7
LMYHpEUJ9XnNXNOqzx47gsY5pDM6V6D/vbSrFx3uDTxSklYDIoujIyoVt2OMiBpxmLk80Ud0xlX7
29BdorOwYd3qGafafDGBV04qGAaocbz6ZqZWxPI0ks9UzgSmBfRsJRSrNs5fJv4d51mQeF4JURji
uoL6QMs3mgfv7YwyBqx7vCssoTkydqyOO6mazSjLMYCDiZY9Pjc5Fss9M2whjI55lEMxwxpEkz7p
cgo7W4dnBhjo2diPZz4zT4x5laWS40AGsqDNJ2bXnMjchHuGOneaq2mKZSLZpWpK+T+W0jy++izL
pp2THaEBTWgafqko5tGFLSDNsQYJs3HNK1Yta+qkF136Z8XYQ3Js6L3mrKqXC8p73HOxR4k29nfQ
y4x9vewPFnzBQX+TquOlBAimyFtspcmCOxlpof9rflBqTNH1iafpfWxkfJrYBPCDy+XlfdOc1A9U
4iSvZbAOg51IVgK+jASZkOSQJ5ZcvwjZt1S7b2EyHMbK2f1C/3dRw4GxLXFA8mOfFKz0Tngc39Iq
ev9br4Eql9MU+Eca+5aSlGyG9SipS8tiJ9WJCBCer2FGKyR/czZaIklJD+jtGE9nJZLhGmCGG7WF
t0BK9ku0eLqCK2hpg8OLn2IIvcJ58T95jpWE48OGpjyo6I9oz9RehI2QH72XIyflmAYzdufZbpLE
Sj3fc3Jq5kLSexszYhv7I+0M33V9DQ4eLKt3q70obJHSjyUaLUZmT0iUEBETVOzSc8ryjxRD8XaE
NT+YR+6zMBZGOdNkhFaNndG7H8SE0yOfZeF/6iMUEEnqY8G3gGbsSlhcqG9zQ+hDw7ucCx9j5DGs
vIaR0jZuq4NXgeZbz+CYhvKgPym2jUQEEHUzB8UQcAjlYaUxPJ3TdofT7W+IwTe8h4rmenNYICkj
m728VMTnPGDZqIdc7wNLytU6W5LUQGHYhzBDRVH1kbUEMq8SxHrFv4LCuEXatNnDxYMmqb/JMowD
dnZTCvdbMunIe+HGdezzcdur/dudMO8VtQNoguynSV895u0mvNFQ5DDptM0l0qrk+dBcCrn6Y7tP
EvEtrLHaHnbqSpa/jhwZzpVm6R9GkIUDOXvp1aCE7w9wrHBi5uflKLy6p5qEgadrSUvhmKPrFBWN
Kp8ruBcHu0jFNCmZqvwbIIj+lmftd/IshkZvwUWsqplWTFx4fQ18w15Y0ri0UuwEenv34xkHfRY8
w+BE2rc7tFOri2P2OZQLp4dZLasMaOG7/BWN3TOt4frS8tog1efuB82HiRvFH97c5rbaYR+AbkMV
mcNPeIJWZ12hwoL7jVJ00AnNThd910dBHqWnc4dhFE+Uleh9zPCVuWHRiJr7e7n5AMaZ9mSDz56s
c/TQQSVwpA==
`protect end_protected

