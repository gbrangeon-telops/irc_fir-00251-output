

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
jAc2elpDF3eoKND1/3jp/zR+PqlylbAiYUxqPEeJkonmmMj0p4wWQxczZkP8HQmv7tuBnI5hb1Re
XvZ7MbtjgQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
NcCSQniKJvfmu7+yh3FyGy0Ym5XaJUypJ6Y0uQPsa1akcjYi0ta/33mMsV5QsYvu+JmAYVNroROq
Kz/qydAoj148DuSUxGpr/Dh6K6KFEJQ68T8sjkHECM7M9i1ksK/n3u+J02M+jecJiy0HOyxQBNjN
TYNC60RH/oHr8eLrkFk=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
bUAhd9meaxo49J9KB0t7maJQYPBZ/miilGsGpP50LlxHKsJESMzras37N6FY41fj0BrwI2d8gwNc
EAnUne+xYMqJWaUJpkx5tkU3/Cq7YHGk19i4FrTEgtDQCfuJmvvnxIjd1KLqJ+tz2Gc83+JpCcen
LoaQjHQoa/X/vrkqv+GBi5yvXYw3CmPRVPihw2cyPAHh/aKqVK9U2rN3QsJFh6K1GPjF0J0zEoGU
HwvENWUy5CJqY+RhFtoI4cFMx4zvZ9LvGAYIaSHNcjGEuPxJtjqEiRDoZaxAPs4fPiQgVWKDuDze
FLb5NkzGHVW3Pw1VKV9puYBInovkYfTC4nb12g==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
yj/twyTkVkmohkM4L+pOFWHFJL5INTv01+xvkfId4SWEcQdYpyZZSWwRohyHdzU487emKgHzTSTy
GFDvnAvaZMJxmURlvGRprcX/FxMbqrYJ/QXjtyclneLv8hDwZCLiXegIMxugiwW4gYlZjMaOoPQJ
gs8ya5IBC3x9kMPV5rU=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
tu3CqLR7y72d6lMu0BtbwhwW0WER0YZdVAODwj27MZbWzMWHxGpAy3KeDW2xQMQiri7N5lQ02ec0
GWpokUjyJkcJKOv6cAVA0bMYymP9zM81k2IaifDaYhtB5Ah8VbDj/ArIWXDmp920Nuuu8ntuPKBS
17ifrJikBEgCPNkkESl85/+YxK58m3UimCI0iHmw3WvHkIj/sAUsakbfIOXt9rbFyqcIak6vi6kx
Gi83B53duhddmOvXqbhgzW3SRCCdyG0CtC/tlZjBXsJNv2kpjQBMBZf4BiACBpRjP60jLswfeEZE
bWRI3cRILGIwfm5V+sLTGxa0jiUVbd3TzGM7gg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 14464)
`protect data_block
P5q4BG/fVSOWvdRh7Pnb8JdXck5UOzCzmORAqPX1iTZ7Q14Fy/Gf8Anbw2mltNaVWJWMUIVeCWmf
vKe5cgpf2TAOhdxwgNYHbabNA52qxKOLorOLolM/p7gtuXIUWzpsRUQaVY25s8joE+epeiwyfsPs
ZGnutFmtkGkMZKdRwLabvetrUIgiGc7A41jrR0yKfcTbHMjecCUEO8tl8XI/7+J3ANpDfsPeX9hy
BNl6rz4pnboaiM3EdekILYhAQ7BMsnyTEc0x6zoRxhXR7qfq5ok0zpsxqnctIFsaSDaC3E6k1Vpa
rjXrqJXBMG18koyAVS3CbJ5hw4MHJUOVAqro+j2G3ry5tu+hBCiS16/kxIKQFUvVFKJ8uLfyLV1w
hFCHaFBUUkq8Cc4zfouC0Kbcb7VvCjiW4xC2TDYc6NZe4q3SelA6YRpIv0LL1eOLwA3ps5MjDnbm
Yl0qEQae24jxc/tx3k7rBR9+Exq5517tKtN3wxaNCo+mJ3VXWPWljGDs4kPQRyaMEadoBmLbC2eX
XnQGKlhQ03oqa4Qve96qC6VV5HCBYpxTsTLSorZArFNZp/7tZVZ4dT8Ed2YIK4UDqD8pWUD1MWPY
DFtgY/kY7nycgskSo5h6WTHUmZgT4ekWsCR7ft/2TKW7S3BsKaMT836jMDz8H3qkxNrrOjf9AJ+s
i2A5rgDCJh1F5cE4FT6jW31hbnESNRMbBLmbh/97/MVcs8vg7Ai7sA4+MHI/lpX5ym+4/ub5QsaO
8NQkTdFEAu8+o2rlQ5WOzzf2x8rAPrpRaVyW6ij2XVjOKQFUE/+MMJpkkKSfKkrT8uak62BUNyKY
DV0y7GUbO0AKQZL3e7mHIw+zXuwmw2l4M/PLj/Ej5aoO1Ec0kLLB74XvAHtHxb6aC91mL9KOs/eK
FcppHMJsTQCh3PWM0S3ZVYDrUAKLt7o+1szUnnPUtreYcucvHYVJTICvZMPrEmvNFAeEF9n0lxdA
PBNEQWeRBpid8JieRuVsA+a61vasX5qukCtWTAXNRBO9HNBuEFadw72v2wWBSfh/hyrNUZDrJ0Ka
0TgPbWuU/7jBiWY05X15oHPTcbhfIqxQx3o+0mkmxAdY4qCg5d2y4xSfIPIxpGl9/cIuB8mNXFvX
h9r1NCMGSRzHOWqwFg1k7EOjsE+x26Kh5SYd0U5bCpoO+evB00JxP5+fll6wnq6k1ibkh4fNz3gM
Ai5BI3W0HwNZxTIpUKRetLyvsFHVp2TJrdBvxt00uL0b+UE0/QhS/HEl2X6xja5ITKji4DqmOr4y
xGQsAxY2eRHW854KgEp2SaRXd9McqHn/np62dUFmhfvqxzqc1LXqmwxdPyK9zTdNaXzNot4slbld
FTZS4KCLW+AMJq7qOzm8MP2lSF7qhn4Md0iwzmh7pXxXp4eJDYOiZC/zIRZsXp/vPUnxtbHue50/
MzroTfCifY6guFbZ2pnVI7kd97RS9AoYJaDM0kZ+vxIr4g/dD38uTgRX5t6NvbRYyP6FSN6uKMVU
NI9um9NcyFht5CaWg9RubchpDlervtEldxDDxrSMS274yld+D36BS5Wakc7DykRnl81s/VLnjlpW
RvP8j0dNBnuMIClRy6kcXtxd2AtTRVWLahHsZO2/vplAdxl40m8Jbtc6n/zalSJHs955wMIi/gbZ
LzHTf4EwlyTYHsZLhzCEgp9aT2Z+IysU8YsC1ayWu9fqzWPqA6637t0/ii2gmHYSoCQSUzOX2y1b
eXJWMGdITX2VAVA+7w7uDZvuIX5bdUYwLNOu9/B2D7kTzI9jsfdgYk6FTZlSs78/S+ezSx4ANacv
nTCpVvd+qacLQE0nu1J3AeW4Uj35JEbQcOoXKKfRKc7Aa7UdQdnS02KX4ncjD7lvSogr3z2xFFG9
3YIYSek2wpwJ+S49G3jITRV9YIcStBMzXznbhHUj3G7GalWMsFvVzAASCtKqNFZRkGCQFcTBRXyw
tdFRDNbNUE+/B9WDmAufPCvt/JNOwIT36PzyapsEo8s/W8nHAFqUhTujo0eEY4djUBgjoE09gF7T
+B0QYVqq+xuDUIXtBGC89ThTvGyCJFwYly12o/ICn2HyLkuapbw6NmSol3z7zSiqXSskNLbOS+cD
aTERiBlwrhcPzcNiyd7dlDqolqZZe2MWlnAtkJ6Cz1DPW3kHQuHeN4+H9mqlEYM6yTTO1+nNTf0t
9aPr/qfPFaSAxXtaHacPMPNvpW/a6rNX6YBp2N0CRVAOnNiSR9H5OLP8tblsm4i2/faF0pSCSJvE
cZ0v27ANm9ubgt1QnOGVFuoMXwkN0vdpwlxT5+99W8ys1GJZV1dxrT2oyCmMz7MRd0AJ9m9kAW3/
Fd6UNTYoRDiC4OhW6qIdvOlsCH38QhdWQaGMGBFQhPWAVSx8yPTOd9OIsxxTZtdj7NL+1Xup0m8o
D97hKhRtQ+Mtzxxuwl5jverPBE1uqGN9GLIB7Y96aj7vMMYkZHN7l8GCbpNgcsbUBXuijlNo8ZMQ
Bq6iukvSDEqGaZjDZcMqqOCqLikPfDJJe1JI67rcAGgtWfm/YCN3ff3/1mafQTx5ruMo+9wR2E7d
AMERIfQ2j9LnoKjJtCMge+atM4Z1WWrOdKdOYKxILJN+LTHjxBAXLuVJFu8yectCgVZq4K+Lqyt4
gQAG4e97k/uBdoRAbWWDdmiEP8yJIksN79LqcoffGfVykClJSt0L+mU1/r4Uwjzuof1fekdL7z1m
OiQAdti0R9Xih04CPk+BKEm7xvD+ir1xT021v3Zq+RQh5AMNLB48auIN5690YK/SmFV7xoPjcg4a
GLq4WMNGZHWsjpaYHOmfs9v8wLiaLw7lnzMlx5UvWeqnoG2egzP8o71oWNEn/QFVnxIWGsBSZ7Pw
spNgI1rjlLc+y9g9jMZII2BIDVno4jgFyrMqx99mZIPE4Ot3dZ27+lfbcOWymHZNHrElwNj0MAC3
dAtlEQjaa8wlkdPrVVyEIs8CA1mNuxGEsegB97gCCWTUhSNyRr6nzc9+/5LoFU9WJUwjtACZnb8J
kwD5teAb43mg1ag/qhqa6oMl6oV3ntd/JLGIGqOs1+Dm6iu5BdxG3CaCh35p7bVwj/03JKon7CM+
Wh39GwDNU98vOj2TYg+2cSCOAmIDDcb9nes+VrXBxf2nIENQvNuA9gUEjHiCHL/7mmhfQNJu79Sa
Gs/nY7U3Tvg2wOOlZw0W7gpO8ZSCSdSd7IqWXEm5hypOsBhs7swYyzRUZjt0PvBY0qLepnC/stA3
Fcli5mZMyBjLs3GTzHPxJxQm1PxCFsse8oddMKA6bL5VPSiM+P/DCMaEh/f2Hl+VUPD9rNIckTKW
8W9G7egnuJ88LF7Immp/h0jXmlAgn5EDemWI92Zuv9ZTpEqegDmhefC2TAVpZOei2HGm04SBQyig
AX+Qi1cATDRNYOXuhnzI9UOKb2b6Ekhx4mLAPjIMyl3mxRK2ojpyXOV08JbcNBN+DXv9brgcVFIk
U7Ku5xrAgrWNdCKxan8PCIuaPgAh9p5tr8/e3ppxLBZGIMBEN4zFeaLZvEJyzTxgTw0vWqsYhiwG
p1gCgxm1FUhHt7FdpzZPGBsZQ6gAwiruXgq8qTQ8dyTA7u4LPhr/tRq8jazTStPnDS4no6DDSB2r
P65Upf15a5AthvPSnrSGnvVXwcO98n287MaB3rt5Bxj/ofB0if3ECkBl0xFeYj1smkWq74IhEuJd
KwT8Z3Xvt1g8ilgmRRbQHwx56X8uhjI5rnsw5vYrB5N45LuSppNvsl8jHwLK/SihsKuLbrMZ6cGn
gJ+SVMjiIFK4q9BonWdHaI8gDpkRL2f8OS8E6gi1jvuy5QubP2x2R0sH79IxO6iNKtjWN3ycQSBG
g4VuU20n9/e6ZZfMg2UReAslsq14xQxG0qjd5HmHNwhSa/r96H6oQbRijM4CoNE3e3fSJ9SA2lTy
nEGRK9+zv6vMnqnLRu/7T7Gj03IXiQkuTfvGThJPzlHGQvNMA+ShlFA6EpnNSj5htrvSUhzB6T57
A/oh7r7EQsZDy30CWG5p/F01yWmIQCoJ2piOK08WM58yzB/s1bit9yT5u4Rm4QSkJuEmqHuWVWd9
QtlRx03WHRE88r7zavu94zRTv0INOxf8+A04i4Sgcsf23Qm4Qc9L58TRkwBPLJyXDc/qp457vH4C
UFzWyTzlwwJUvHu7GloJEpqX4lePbD3gH2YMNCQkpKbydEgUsFhSWFimgHpAQzq/wFl23X/W92/1
fRYuXs202l/hOIsKdgyc8ksc3VZ+GgO2wG4a0BQH01UcS8Zs3eMoI0DsaDqlu+iJzO8dt/iw21VT
QEIobGl8tgJJ/2CbO3i6zbUIHEwdEgNh+UO1rom5bDMjhp0a4G1CJznwKE+UtPxK4OxEEn2KBNcg
hS2BGfgzTvF7xoAyln45hFY6c7us4P0m0oyhxxQRSbvXnMMeUzIB8jcUG5w1mspG7JwBZTlgPn13
nCvUlZ/W4ibcie4IXEdwD/u18PH9jb1dsRH76kv2+ap5OJgD+tknu2E8YaYTuS+6nwW56Rwh6uE3
P/DzkW7vsUg07aXDldBfzFrjK3kbi+ZJvpwHjqYNLq/2YbfOdcE8l/jPq/oyD8MrTyb1w9UIBQ/q
McyVJdfpyrrUn6NnHKXzt2MiHkzOcqa29ysuip+LLr8lrNVUgVqbd1Cw1QYfgKiZYFA1Qr6M4JLs
98mww0D3j3J2Y8ANpcKEhSoaKY6oe0tek1elZa6QiFkJ0GiXKAf3FsIN3mLBiriPWCzU/+vd6BNC
OgpDz95w+af5ppyE9yP4pz3wyH+MYm5cYfDGBq7CSuAV6tpM7vvWxuQiJGp8vE8HY1xQ7lgWK95w
l39czC7HZ64hGO4W4uKxnOmpyLaYUqDHSzthfv7kB6PVor2NFOR+JBmpCLgSMZU3WbOnxbcj8Fah
rg22u50Uaf+OoUB+DRDhQFNIoPZYhdVJFx818NazHFJA2FQw5naJjyWl8Kvhzxy/Sot/d8IdRz00
YwjgaIEmPDBzkgfJ931rLweW58TG78910V6JBfy3/9z5dt+jscAh8+CvQUA1AU+h5n42ahE6r0Ds
lvyZH5ri+dKUYmbA0+sXmQSh9nnOWnZXWOK21932atb8zTNrHl4zdrjdsOFVjQ3hlcAnUSFUgTbI
rGFZim0Zw8CieSaciQkx/T4tWQcrb7O4wmhJzcL6+szvj/7iYyQbsupC+WJ8PinZFl8U7FzBfaZJ
Tevg3lebZnuMc7elOS68gziS49W7yTQCYtyUArhWgBbblBlumWgIVLANcEoPXsxaX5Z/CU41oId0
Y5BellBqpnAInQHcnPsiJ2Cgqr8SJZvcGQ6e4SCna+JIjDHhrXpOG4u+CHQvQWJptPTtKxkjDIYK
s4cK+3CErPdUyWR+tWQpyEXhtSWT7Hh8jx8Y8pobvViuv0W0NXZspliYGwzAtPXlhV8VMqnZ2sa8
CFiKdlZGCO9LV4zUWpkcAXe8Acy/VN7fN4KPbAIJ//iv4cG1j5wdzTK3BT/1urGNoMRe2hKOiuL1
2Rdk14GOG6HbxmRB+qMk0ZVwlpZjyUfnrBRbxt4+zvUAdD7W1d5pYlviBuEe06tFdrrXm2aGqEBa
9xslzf51Hlaf6wuWqvz7W9aL1Zv1i2jx9Osp+rrgWb2WoNXSUURfrKigYVpzmkXwHMyCA304d28Y
rYyuhcLElG/ZfHLNmzSaNo+6wxlSAHPclNdnDj7GvLFERgDsOP+ZfN0er/34Xo7q26XWx6rTFKQT
XA4MeJXXxjY1+RztzT8as3u6PVCEzB4knHciIfn5b0eqK2NlFsT7SfBoypVR+u+aYHhLG9jQwG8G
ikYQQ7H7gAdg/UhduObdyCIBeGpzHAFhSJ6DiY4DL+ZtIDbWkNtINFGe2Ny2vc/TeIrdGvPzmzky
e1ZBqVIW428cDcvRiit/KcqVVCpWp+U8OZPps80zp/FmlnIGEf8yj4YFHMLomnKfHmBcBsy9e2Lx
XU/3ldqDSwJv0kPkoLS9TQ7SbrXZgp8daNFWQSGwroeKsffGa2hGjFawrAN9n+FMI31oof8RvK3+
apUTCJjt1sB8+M/Pu4J+oRQpq7/RdCc4yIxTUp68BK05miGfNBf8/aW1I863K2VuIGWsmffQAfRc
RXDZOGIvro8hUC5hDSNchP3fOCjZbiEaW14qp9AU77stbL3ogBb3vJGoHd9kMvoR9NYydxDnWHFZ
t7BT8nOIUXaPZ/xSYpNpv+xxEQT+0F2A8K74HEILOdDfEQXHfClqQUOUYmFHgm8kcLLttVx0G+cI
gizj+n5gUMu4jTif1cIeH0aPh3evbebZ/R7y5jEt+9PVs6b9ZCx0WsLz4daRlR18hfdXia8dWpBP
6rXm1wMHvAcSPCZmd0S3lO5b3xrh+6ntMrlvJnwF1LjVGv9MTcjtx6DEOJgw7OZmDe1YJIMm8NfJ
LvMxIBHfsEZA+GmoKTFqownoP0jsLw3M0Cb45XxT72Xp36Qk3GvuJ/6Qz7BL+g6rPvx06ZhRaMSx
UGSENZdBSC+/7vJP/0VX+Qj94z3oVAEydMhKBpKz8hNAUEDlcMWPBMwuglyP/Wfru5ogRFSmbgUB
JAgOggga/fRRy4tmLmaCbI+0ih7Pxgp8tVC92/KJwhcaWhvdVbOeFNCD3uTYpX+4xOm+/cHYGoEZ
gvbAezDQECIu8uyQ5Q0ll35z9g/gHaqgr3610LTH8qqH+P0aeLD4ynp6vVfl0zSST86MCaks8XGE
mpbh/m70kqLhIR6tW6aEiAmz5Mc6XO5lUr+VfFWGAwpY/K58u4h/kAT88GLe5xI1p0krKx4APu6T
2s2J9EVRl0AEU8f6PA7MPnwc2BxzUfcsM5qew2YbkBP2UdmjX8XySrQL/G0u5A6Epa9okehlK0Cp
npZPX7IIYVSgmCxUES0+U4LTyoghSaHwNlDw3X71cFaTkltcDcFJHiVXRQ1WkTlINAn6h8qnZAa8
w0oYvzgET6ASHREOWhRn1e0i4KAT1cU98khajxhtEuiEj8XHpOVMnCTBxUcXoR/LCD3j9WOKeZ+S
MFr4N0l7UoGMYX/Jvg+CH9gD3zXLZmwYCJl2cJBpffnUCX4j/xCC7mKV5fAuX3hLX624bBcnBK9y
GoD1jdQFyC6ag4Vm4T2i2ai1WYk7bdFOE6HyHAjvC/wqDyZsKnaYUqAjMHw2t/Em05bD1xCrlQdr
yuGxIA4/TX56b8frQnds0DDURp+RimrGPj8LSeiKJD8z0vhpmI4/lNz/QApKflJpRB/plX0UfV2Z
eSTPamjol8DXfgxc4L25Kjv2zlJlGlHtPEV3S+L+lIICeg5RfuOXFmcDa07PcavPj0Lq6SxQ5bk2
K+t39YE1e1SqGu7II6eoY2gCPkAb/MKazEPuDsXdQt4lm820cg/6y0LISnC65oEGuNm1CDAtw6YY
LkB9Ur/e5A9HUv6tm6h5WULANF6Sna/yOJKM1kUPm3txCR+6bUuN4aEKZTP8G+VbFQXtf4iskwEH
zo2y8+0YZTBnntfuh8N6HENsW7Mc01YOb4vvmqZhk/HuNDiXiyfetXhp12nXfy4lGFtEJWsaxDci
vwrKg796LXGwy98/y+J7Z3BAhUA925OHHRro8Hgxp3B9pli//fQyH6clVHqemWBTebdFoR1AU9SL
xSqJNC5xdSk6RyDcePD96D03B4/q8nEFf+oidTZk4ym9NmgeU9Hhptr5pxGbs3rKK8T0v/3OHANV
rFC/6hMxEDti5LR3hEwcm3a/Gdq1fJxyI2EIiZnB8DBTRHCA0PxSX5ECoTbh4+sHgrEhzG8yg3KY
dXw9hAgnXIwLYQ8WacZcg1r6MEgqUCtxsxUi7BVEnIM5Wjo8fmDHVwa2WGBp2+Lk8iyb4yXm9keW
ZRgztJ775LjcrEBDRvrRVAow69cMi8H3MZyykWwEszrsXHwVXwsFdfLh78t+0qa28l+JAVYKqx3C
FFMzVhE6CGSTRSewUXs8PtcABmYfsOJe/HatzrjADElFMHh3r6gjf2tfaMikiE5+pSM26gPDcPcQ
WbtIkjlZmWmnI2tV30kPdmiLVTIEBwGRIgIAPsuKJCBCuzrQnCH+wd6uEA27MznXnvy9KJVRDUPc
38oLJmitymQiwsBWrVp01ELS/BAx5zBLqjfWg/+yY7vyw7twLvwyKp4Xlu4LkBrYgfEto+d+fxPo
Mg5ET/0eNxWJ3MXT9GL7kG6s1t4QBwKPYt/tNDKFLw7cGk++pSM5Qof93s9hPgCIfZlp/icaxrbv
UTzsFuSsjOLr7p8fFvu+Ff+brmuCXk5XsuHRzy0T5DyTHMQsT8R87oCTl+xh5oigEfDzES5X7p4W
Ovsv+ovSmfmKfuj1E6ZvQeggqN3qv0HTyIK3xz08/tv9+oYo6s0/V4uAUCcwE/XpEV4mvcvcqt4A
CqZod0Yc+j6xu9+2GuFL3xStD9nK8WDvTl1EAxoSjx46PVLXkqmRqiH0B6NbE/EgOXq+UO+VoqYE
cdVw1H7aExxtiiZiPa9lEx2iVwizvcBluKXkKJEpaijgxXv8HyO2ECMAllkThP5nP/FfRRrgre3U
o+Fdw8euuI3yhsy0KYa1wLfC5QeOqv9+2vkEulqXXFGxVwuj5A7JZbamWHm7puTZgc0zpJmyniAt
B+75GU9AJK9n6pyrY8QZi8hmWUInvgyq5bxTuh3i+WbpIT4VKz4tN4qs7kDk5bHeQybX050QQX0g
nzzaJjjha0kWwmhoGz+RkzvfyZptQWQvly2Ic5aaZhFxronXh+6cU8n+6cnjlEWowUjQ8weLDOyz
0POPskZWtwfB7LgkgdmaWE1TYL0gC0U/zA5Q9pq4/qW4XEIVsat0SNQMlpAzaVHMMO4hlEpHxoUv
BezGbHvBmb5PhNYV/kj62JRSX9aiJK/vJoI05eEUuBFJzinEbj76kxRP5QnNhcR2K8wKMa08gPDF
8K/I8xUPkW4cCR3/NHiHDZuiGqOHGlJeeADaFUbkh6GIVuCJPbw65+WxUY7qp2yKBPZZWIuvJn6u
aFjbt7aw0NaxXhbOEB5+NMTkhdsQdXytFc0qvSWDQuy2z89THUQS4ZYkrHWxghRx3wP/wkwpvrej
1Ct5oauxx/SIWU7yWm4sN9r84wtcJDolIaNLtFnfLon/ua2sDp+dgeMdAUJfPyX4Fqq5bkrG0qOg
2tvTzqZeKqyA5Nq6+7cZIpjm5NYRGWjt9bNJn/74tHC9mRDWlDluQlCcDPn9E/zccu2vQBPWpjtT
ZhrQDfvf33CVB9iSrjSZCFfm7V8k/8n8ruBNg1k+TIBg8mVtG136G/czyf4RmktiuXlS1grj/xVr
LJKXmbkSMySpmZtq1JGPXUTZPFVePknysOX0Kd7mQY0QKkwHi5yYg6PzkAy/6ZSGyKmX/xDQEWBy
X8jSIGtWidwEEbRqrAb8SGy/lIerRGJ/LYG4yXY24m8+B2rdTHxbp2sf/LQ6QOJ5eA1GCqrQNu4w
Vo5Xsn9FWtuV8CRedYPM1XagnTv47UZ/pTXq0lauiugGk5tgNjzm5P+P8pn4t46HwfdqH+habEId
McaQ8reYBNQHkcKSjEHb7SC7vXaA28t9nIx4vkjwbIpyuarth2zoxXwCFL7iAgf5temjgCudmhLD
RL66REM/uWhb5kpyCDe6ZC/j9uHpubfAL2ICUFuAsDdT72QnYI3cVEx9fnxCd0SfnWMNBO38lny9
Y6P9FNHrnU+Hc3KfQNHiafmI/rcwGncxZT/M0OtvVaV/GxfhvP2o1AQJ0x7AvS4aVmDTE9KmzxVI
iCGALJ/PLgB6drfx3G8DXmadvw6ZlL32BlE/rCAF8Ge/drewAwtSx2aTEZUS+krWTGdUwImP3CmB
y4UaVPUCBP25DGY6sutgMHOy4dmZ4iReTed9VwSLpfQqi7Kmh/FDbpYOQ/EQcp8wU9qiM2e/CTzA
nKQldB3iU/Xdq/b73PRu05Q4TXGC7yXEa8dxBQ3/NfFOejcSJJRBRAytBNsm+n97iHDQ84vFqRIh
uRyg/vrE9f6un6PUykw4jI4vVAAVw2Zlhzbc4toFVy6ufxTCyzbeAQnLmSR5VekKB0xin9Xxu/nX
Q4fQ+wWFq9Fa5tTyCgYaN7KzeaJrJFHoynmwDHrjjFKfd/AVSWb1CTfy6cMGFYLzqmHOCu68xraE
v2srm/+ZCxvDf+TFjC59plO+hLdc50xC0b0EOmE8ADyWmwS5SwpgokQHao0OQQkohB3oPQW/Fmfj
jXt//BDQU6q2onffGmu9f6OB8hhPWZ5Vm8fhj7onBXzsaC07DgMwLlPP0LVIqsR6QD3MNjrvGBa+
4Mgi1aCN/DP6VO7iovmYbUTU2YIdN9PrkDk8rp+3QcSu1Iy6ttYjSC6c75bTZXh9PcNc9/IPpqLc
/HDNQCZjCevJ+Dmg4DbxqfkMVDzNBhWZNoiqwusj4cTw0l/wf5hW6NCPt/yEsfCdDM8gqwP3tICv
qYTt97uPWDpDtuZRO/CvN2APistXAhtT6jb6oWZZ4i3bUrzY1Ngkyc0E7lBMOsxsMPkTvvBQV5px
S1I/jMgvn+IJeDsiDFCBcq4pGo8EUYo0/5hytpB6OyxfbgfgtH00A/bYCAnJ/vC/OMtMchvH+C2O
IjMnDCooBqCoBMwqz3VAd+4+MZG2Wkc7oJsZF+IxOiCHjn0VksvvJ2dxftzww2UYKgUvcckOzjjf
qV8hccZ1HqCWqxvq9C6yBSYlL+0TIlGZ0ggPTcQMQ2SkRL89J7xfprr3vgUcaVc0sg8anR7M+3IH
fUEemdbHdsutpopzpBGhKPfe/a53qvkDnlc9t9Sj/bhqPzTyyzMIN6KcEb8WwDvteTS7PAHjEfB+
VbrJPh4rxZs8OLe5hEaloIioI7jkNrqlqmnWX3BvD8Kbxz1dG1B8tBODgyo8UBMl/u3DdLB205zK
2FIpk+aBNmD1XFmQPni2ssGcGn2eQ+WkluFrrhJbjIFbZY4o37u1xsvpQkz0FiZAebEIzNBCri48
stxNDI/fDbhRpZYfmms/Oh8cyq5+Ftp8yatfcmxU8mphfPH9ax0iEY7Tb5PQ9CShvi8gbMUk99eF
4bAs07EIr28lDuAGC9tPkrrBp7BRzNVDBqLrTBdjYpYquWY9A6Rbj4MYzvoron6CFu48wayH5AkJ
5xKm13B/qZRAp8IqgpFPiGZsh6kxbgwUDc+z9i1d5zFoKbdLnwZGlVL1D90FPcoUwyuF4mO28LY7
d/b8fFbbO5gYEaHXdNvusb094g2oRTtmpti/HRO1m8+etCczt2SYGRccTFADrYTbKrFwLBvD/Y0W
TxWXdZI4aIKhLcocMbBMbjooryPChRtrz8W77iWGEJdISxR3hl9DIvXLN0osSBI4YYzU4wYIi+fI
A/DTpDgNNOfL7f8os2MrcHFllYvFMTosMbvp0p1kGdR8+e6OER3C/uRpZVX/do7K/GSM1j8BZ7+p
7p0ei5c4aZsv/n93U9lDD3YUgrgkXG6CFaN5PPl5TFqlUE0ymC+GXOxCzKEpJ/vbn9Oi0EdoW94x
P9FK4Kq/1/eJOIxZBXxlw/LtO4y9v2y5ku9ZPxXJJ/u7W9gBDgc57DWDOepfzx9kXE4y/4BkRFtZ
K1z6Kqx08ueCEdFtSFUAhbkBxtmzMBswFxDQYZCFfWQ6W5w2M0SQZfZi4bxSO/yl/f6P9UhD9OvU
kxjDPchutaEKy2+JS4jJgoeIddJzylpNfry2yTgi7a6Sobc1/kRfwTCdu/3iBFR3eNUEMJn85u0f
6h7+C3VOUgv5IcXIR72dFWX3N64Tro/AiqGu2hH3VK3ksGBx/gf6CBqTReGAfeAKCrp2PsQpZ0RL
vAfw7PIHx+Zl2y51WOn3cuOI4Gv/AncadC79Aa9kr4zeVDN+3TlcAstxWCXD5ff0mdlS7zEAuvyg
gxaX9zog1ZCLaLavvmJqltVhtShC5AYOG1TKKEiOHY6n8UHtL9W68r3F0q6llLDsl4DVQQUJRCON
CkqjOz8yf62N0S/nn84s9qF+4sf5iWz74kOZadkrJIxDuB7TWEg0q2hA8k88YT914Qc1bDHOWNMg
a/bt6zWE4dtSdsOmbFLD5QIxxbLVwGHppRS1ZP40E7rXWsi9ca2cm7iHoQa4t5ltp4jQ+dIU12pV
fBk8XsADmV3dbU20CdpEKWHWmNMft2RgMXhI19Ygd5YBXLJJZlpUcADkeMTcDm4VvAtfdI9g2TTm
/lDMxOBqgM5HC+QwSdu6mWD7/Nkiqv8d8jyOU26bGN/3HqSmIPRfzfOwaSHEAKvRT/i6kEhHNY8J
R3Nq/1lwruoljQ4L7LSmoE11x+ulisDPIZ2DR3ltxixEnnrIeBLLaoWaiEobpNx6UxABw63VMZOt
U4RF5PyjfyNHbKw6mHMpFuADyMBxg7UZkQOK7TQQi7C1RM4yVGDvBhZzNs+JIW7pmYyT3WTdW2pO
PXrXM908oRRLgS1zFlqJ6BJkRr0vJUgP6IMwsiSKcG+Ovu0ptN+aNnhFw+/bLmhvzmzw0sLR/5eg
R1NpXbDdvB3bFNOGgQ36HW9f0PaNtMJojxnDpA0JfkZn/m5ZHxmEIfPtCmYviEb1JO+7eowrpUDw
115ult8DPCl5dM1bKGUUUfeBOgFLRPebYSLqyfPZ31cwcYT4kqUfWro+IHcDLNfMWiMP2A2T4sG5
HF0Hk15PArsYN9N+HWuQdR+2e8XBgZd/c6YoZQoSU1RXmJVmBZx4ej5rTwsQvLZR7oopzmfX4jbi
TZb9hDYe7uhLbZfJwWp6KdR3R6uNFFGL/s4nH7ibmWHPutyffuc3M2VdSKlY0nwJ1jYRhdExSgKJ
ds9KH2gG3GvOs8Q6NbLMHmfr6b1RVwIIbMqtwdlcuYEpK6gmOv87eT3+FvOMW8PB46OWTo/TWY5I
/zYKaV/dCE56R7hNa1+aSuMY4E+5hizscLmYDuajtxJ5pPYKAJF9WdEmeQSDjYojxs1TkyJM+Vmk
q7fW+T4SKTMyi/PvyWDCimCno+E3XeVCDrGQdzZgBKaUSozR+4v2Pu7ZYTtgwjOj16poE6+gL6oO
32Zu74Dw0md47naSLGMb0CHGFwh3ujI6Q3/inLM9o/okPdFzag7TPxhhmOhK/+WyN8M9pltiF0Wb
PsNUiwrYAReq9NJj2EaneDjNLowQHFjFKUAUMEIBirmYDCQlqZJECBW0vkKm3kxXhJMBgRGHAVDr
HD/unIlAm+kyAWvyhyxLM5MI4bExEwA4kI/CX5wDa9tUB5xvUR8Hw2zetkQMCpmvjh2IdFEFSvC+
FBYv+ENENnVnabpXlbYSW74BE5qhL+s8Aa84cKTlT0/WfPJVEF+8obj93qKKtVFfibqn3anv9qaC
SE2POQXARHy2mcFCtxJfdrxPruFAfX7R5Wa+7vKSclPNbeKdPfSnuq43ix2xt0nRHcTDeVJ5PKTY
zBqgEWTaabSwBJ7RBfPB+mSOxtJg2r9cCH1LJAtI5iv0A2RtOXyB+B3rW3UnnOaEgCBEsRxVm1ex
ev+1RFd2fME3EU9rmWfvBY+IL8/+C6Ge+7T9C3P3Rcy1NnAg0DH4vkLBps/uxOwqweq919TKyC0n
QDUhP/Q6vquvKhxahwbQLBG+5cwjPTTOPqrFtFrLkOAPKZBW3c+HuZ0VrnWcQfQuUNoBs+IAENPi
mk1Ktq09Sg79SP1UjdV6bDfillN5cDnfePT4v2436q1A1SkVKB6uC8kJeoBDISWgAbIzn1cKdvKM
58kC384hb8R7QQSHU0BlCFpH+rhPYETIxs5rRp6jbyZn6MNqfIVp+ec2afpju1wLOZ0rFVjT4Hg1
NHGAQhXgEM2r2MW7/cdooLiQOEuR4S4jV3n6isJxMnfQpfKcPBtHoLIMj0Ty12HSCe8wjb9sCRHs
xul5cYQQ5zB2IXkmnmKJyuKdZ/pIXAmQPQu+4mjNoqjedSa7oo8aAHWkE5/0PWf9/ND2U8VFP1BZ
lKQCrjwttrkEusM+nG8yeDROo5C9uP9umhaooZb1X8g2DxHzZoiwfS2on8qE7E3CYMdpyeiyMVCF
ldSvPRLKfjO/8dmsdhGeP7drbk1r1g5JaSTJVoKL6QU0YU3q/NWXwbu/DBE/I2p6blUIXyyszzMY
yY6sS2/5J1pxZqTYA6LTDIsHAf7iPgSA2uApRvU833lm78VnfdQc28X2N9kKkZ3kCAHlSNUdUXMG
axLW+s/OS7kCuDpKbkjXXb/ss0yJzxkC1DVrS5isVecXBayF6dqFWIXo8WqN0dsYQb2y/DYpO9J/
U0qS48fnr8q2bEVMj+65Mg5VCi49uWsPUPCDkq+sgVm8dLINgFbx3Pq7iPuE+TW6qRTwh33qkbBt
f+yFKcBOuzNgMXLR0rFDuqnI8JbpLfgVwTkaH6uaiQDcGfLNvLFTmnytAUUIPAYmQana6j/jJifM
yWnTOekxD2Dc5nOxNqWQqmE1v9dPkG6SE9cnqx6qyvkJaZ7xtPRjFfsM69RX+f231rz58WCHbNW6
mee9Eph0wzaoiidnN51EXEu5xJtCggqQ/RKc4Dc9MthX1AKIpcPgrKoogJxq9BA33iIUvDCpzAQI
OD2Gx3WUvxARVuIraBTMV4a70Jz8Z6tFg3WFzH03ZuLvM+A+GvFGhfX5ww4hpXOn1gDiGnlVblZ5
fF2k8z5AoGoVZzJXJsO0/6GnHsrUDEcQ7kiipBp9qqbz6p2RLK5mt6lTUmEFsmlwl3JK1mioCdZH
48JMu6Cev7LDyO/GThaFc7V/jkGBE8grAUZuEIH9FeR0rOXgRjZBH87Tp5i89zrSn2PTfZgIDriJ
WHviPI0VpCKztGo+Aq2CWCEDSTRnJwlFJeA0Lsq8Etg8oLy85loJ2ZKZv1svrrJP8RNBzJCHkVGI
Oaf048ZntJs26E+jB5+pdJpSReYNRlLLQLDoRINXU6mxEMnF8Nfdui8TcjgBAIXi3x9wEmbHV2lX
2SGTQtCILSzeOpIGDFa3jlhLam9Go6edQ8viLJ/BlRzxEWYD/EdEXhUEk0fBNriWjiHNTb5qPWF7
pHOsFmMQFaXm71T93kGK9rUaadaFqvZv8UOjzeJTUIbR6iu5NxHqhfSw+GFk+KkhRPb8i0IjcjTl
NvGblqyp5R3Goji32iuue8Dsb80UiNGGIY6IAoC9sRsTHvsJsYCmKSBmpolHGpvnpLgGMShE1orx
TmFGDfEAOX5Hv7XxnVYhVU/HXvJENuZtKTLQzzH8PpsPWWOuoTFd1Iz+Y+P6Zn4cqlyCNKgRkqym
B4CFQWWkCJ7S8fQK9q5XyO4onerxK3QtYfb3T006sQJ0AjgfIc7HxFj3dWXr2KCpszIR4r1YiaNU
yycFgTvDbuVbKCuSdf57ccwkl/k7FtxnEYxxQTx+TGw2TCjvsSctmszxjIBLdx1+UkK9OnQmcnX4
oIr8/Rf13Nc7wE2T6TfD5CE6rCpGsa+/2Cn9JMOO6tuBXv4RVRt2VJlb6nPtaX74mgcn7TFAiZNS
uo3T8FaUllNSvQRUxT3IwthcIwi2rhnjkucCPaxp/+ITCYmoyDqDhNQ4ZCtiwO2R4iid11FkqUAc
31+qqm4n35N86fO0JOLktiSDe8kGMxTEKqu+b2sDpjLm+8bRyIR62Gxws5L69sbk0gYXvC4UyR7+
Xf9VOlbs7BG/AhtThbVTKe1rVHbBQawxosClW1BToEhA9LVrcfDxW2BaN5VvH/9vcdfpM60GuTpP
4Z5aeEk9PJ4wRWtWrc0X5Zb61G8YtON/U/+k42GZLYvS3AcrOyRfKAtlEjwov6meF+yuXcP2/Rmc
eoeiV1gWq//DrWi3fQGaiM6DXRawK89hFEluAztlvFtu2V7z76BYZDkAWITc6unAOgLpvzFIr4Of
gZ5mLoQTCf6VPQWMlSM893bJYG28u2yn1/Fo+DjvK87Hx4AZoK+Bqi+MFI9psxxJ8VMHByQHd9fH
CKsr2NbiirlgG7vK+/grcPUF9q775B8kksjd8ewUbYdexls8/x74uJrJq/1pbo5HWOXmBzKKrUws
tl2zPg1/u4GlsWKPyrMI2ZnAEatyaB5nLWuU10xgqs2Deyr86MkskspED9WYKqG2aMdsp9bXNawA
AZr+fKcWgwXkxoUP/qMKZyjiCQCFQriZinDCIHcs0Awz8mTnd5glPvRi8UHj7tqbiOmw/jnnC2Sb
10H4PtxwQbzQF9BxZ3jpHZC/BBuKvSpADcxRiZDx6UgZUgqb3PQlznJHs3QJU3dHNJ5D0hR+Maov
y4iyKrN6DdCGYt/GqKbW+yBRn4AZc+fpIrXpP4nl8+cL7fdcNL+Bdz1m72Jwwjpp0DXrtgDHKsbK
GYkdawSzdFHlDdYoVnTDIuWzICNMA+qZxLfb791w4gcLjBT76tm3lCW7Xo0vIaPOZsMhXxfsX0JU
bfSU30cdQ9Fh6gxtDHRve1B6OstMJD/TQ7KehiewfXGiwCrG+p1OAUBpyEJxf8XxAECS48wxxdDR
BXcsaBDC8LJNEGazevaZ+3vCFkILnSb707O7oTRaBWQNPxGDCFuAgwJkl8dctjqGOdn1ySvOYX0Q
d6B17JZYXbbnQYDJlWbk24ANgbUaR2burHmik+RhBOA/q1tPUzlnB732Vdulj3sYLYPwQxHXL04H
f7EEaMS7EkZWaP98tlpW2LgUKM9QDMp/SCh2PQedM/hEWOYQ5tHszHtecJG9T0CESqP9DrlRd4Rb
pYEOfA0NhlMvOAxk7TNNtvuLCbD9tkIj5wyX15ij0w9LF6twGniTiczed3iJpDmDwww+cfQn/vQL
TcUez6cAdxVlkbDYY+DZRd1teSnBIbAAa2STC3UV3P0KdMx1Hqc6nkSf8SxRYnFDrl/KVYid7Vcq
t7ncYXpxZ0Q5UjDbsjAIImzmcDmvwtIafF1vs6yDHfQWx/8bhvJ9EjSo3PquKW8HhUVqYx8nVvhJ
boNxlgQmgo4tur/B9fwUGloF3Cf39lN1ydtdIg6glvzoypDRE5cecpto2X6DfFegrXsGuQzolofD
WMOTV2pPEg0vIuOfNGQlbxBPPjKvwigjXFtAHqB+OK/+jb3xJlwx/HDpZzo4GjAE3kRaRZ9ISeUU
fmWs/cdpaJ9xJeOdXBprMae7U4K7lJ/c1lt7Ddb0qsuH+WE0XT0wtQsBoRxPSN9j2pNTjTS1n4lY
exb22i+W8tN31AIssUzyOxoiNl+UKBlomaAJr6uDOqaDtLblKUFxGhonBOPLTfxRC4jaJYygBPLL
ssCjrf56ZDcaFWGq4uCW4p8psTsfmEDsELFgLBYZOB1gc0oD+HYqwwt3SzXgqiluHuCBSpMMmJpH
tgp9IbLO53NUASK2bjiKhN21QsFhScQGWBXJVXbLDF2A2zOeoz6XVfcCHHofpmyQ60fC8FG1GAv3
eDjsIyXmTeB02minIAKex2GOFhHdTPlS8o+CpMaCwhB0EtZfa43HHyR9KfvfWSzcwrZlIWzPcqp4
ixRxAQ9mEqbKbjABeUfUnd8myUwDcQHlYXEAhaZsoQ5Krhg6BiQEw3rJDmPsH3nlgwkLpMdDFxu5
vDPsoahOz0q7/GMHld1KMK3A6QbGYdZj/laCvLBjgTZB3McB03oaWcDL2q4CXgY1NvlBJLB2SH6r
M6ARUcOEdlWMtP7U9D09g307Y2iiFIgLkgd/L6HxvX2wOI0RhiyDG1ZDy0UGMqAj9/PekhE5P9nk
sfeAZ4JRSZMrIsQVPtsRTKM4vpIpCfU+dsvI7ZmfS14QL1HyrK316wMD5DDmk5MV8/DwCreabgtd
b7j1T+Iby+1C9Th7PQR8uGLD+Grz1SZkwd2QjMBGqcyK+gs6YXcxKcl1/M4bhYAeVWBKtr7vBTQh
KkC3ZVFNArd6lu/FSaoy1DAIpoJV0gfVuyGHrycT3lpU2/c50viK4ui3Q/uukwczpM1l+CiTwuss
oh6IU75BsR21nO62jZkPv8WkeMkvBPQzraxcx3peDAA0tISP7CEueVe1u1S4uGYCXNXv3s/LtiqI
0UQf+NdDOQqD+Nk1llFkjZ6R5Wzj9Htofjza/FGHOCigOweDsmdBMW9NdFToN1TdNNAo9bCPqnMI
hlCsIdaEYHLO4Zj6Uh6Gq4dZpOl5BfO5OumVNHitu9m1ClDFIzypS5QPLhDLquvElaJGvpqqlKMQ
4ZC5Kgtf3dPxYonc81fF+mtQs+8OxCJ8QbxnxfXjXl6AB7wU8lPmrzo3cHhs6vzhriDC8dN3FVyg
m1r1WkBTxl/lVRhLKXm+2LacfEo7HQOYwiAWqUcboYWudGUi6sgLvWalkiDNqYzfZxOCL4R1bIAx
iwmU4M30oksQMFj/k0CseVNCricDH3zbh6BHLfSVCVhietZNs90R64d+bfvNKbM6t5BehvofEYR8
I/wBOMGSMac/lU9QEQQ7pVU/KAlVPJRuR9KVDZo8P1OhoqoQZrmsjUptGNWxmQomSzMLXuAC+x7P
jeCfSoKS40XR89sK0om4fvONHNgOzU+X2ImnFfcCLZG6VWE8x2Ydr9jxRNoZ9QUTw/nsoB3NZl9p
mfTXG5iZsR7SR+EuNpHw4FtLoSy+1r5SXLG17oaadxSIkrPLJwkaC8rlwHPW4zjM5U15Ryk5bDsk
XgCO+awR84LSOcqmdjYerVAnUiK05n347UFw8gc2rLXzEl9Pf0VsJwfQIfwl929/GsBszsYXmw6v
HybLgA14I38sZpwMGG/uplHAKu6QgfFyz62eVHsLUiKKSNKgx3K9hdTWQhIreZ/wW9rla1KfPf++
mcl8SlT41DgA0TFbmKlwErpjsWRtLKVpKCvCdoSddLtFuG/PBLLFzOb1FgSvc4MxXiC5+fuDfa1G
oXrkw1/knYFwZ7clofg6qTe0wVy4uP/kG64CnQwAjY+sk37MpioPPWVJMl/Ki0E//6+n0Z330YR4
RZLEwsiumCDua/WuuoWjxLakqYHS5o4dxSGfjbqW8rMbHNxIEEDsPOS32SaeLtGd8LD3Ro9z3nzc
X9FsvtlXGADCLcSUPQc1fjljqXoqj77GiUMPqiK52bKgXHQyViQ7yT6wlfBY6fceuf+jCEko8Zyl
+JYWFjx3FkD4GF/9J5H7yqJ4JlPJ+iRDK04bYn5ias1Uni0t0y7Hy2TGSpSRajWK+BROBe6+4BJF
n/rz/gGNoC4cYjm4LTtrCkS7Y/EgGkRtm4Wy7WrFW2EAOwcHCtt6h1I6J8kOK0blj+fHlfTeamZ/
DIpHIQ6SEZfLNbanlCkBymUyLKRtsG0bsyjHTaslN9UVqo36Lt/lVnItkw==
`protect end_protected

