

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
eRz+leRSRPpou0Iyb6bnhB8hg9kPbBirrzFUAdKqw/be3+N8ZrhDizYaLfXqnwxlgZsSWJCzRfM7
HvMw/rTLhw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Rl74r1iJC/bnSjzA+Rx4NZe56NnmjoVRFzUux12uAkwgT++rVuZ0cWQxVSY31Gff9TGn02lNxavo
U1xWF81U2u/Zi0XY7ZHmbpbdUEdpSv9huiEIrpuLuTgWjBSUwsGYqRxHLx1vq4vioRXFlAhPk9JA
iYodwxjKI7YbbZElfVA=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
lO1ylq105LQ/xiJNZcB3fPTy1RngsQ3yQ/KJ6FM1qs+SoXmUQjQaEb6hJLPAypYN8r4VdJAzSC/U
5nFe27DWNjEKmiIleROkH20okne+9N7+PhPIZQnib521U3SV/ecBImKKPYRpHhAeqE7OE/DzQFWx
10ISqR1I6WBii4R8gkz5k4dkFHhiTU6fgkIHLUXXclJrpQ6fHHlk7MPcpQDjK7bXjIiQ81qfpVmp
P5Kh8wiY7VppUj33GlIcYsNio8GAIV3e0kBKLoX73uDqdvJ/2zBzKOZoDd0As7C4AHF8YSixL0MC
djalIDRCSOBX8Rd9h057rIe8ZIXNMu/BHoKk/g==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
aJoUzTg4Ju9hNY+ZPcuNUmGg+rCD8aivgSTst8VRB5/g9QHuzghA24ad2z08gxWDFeIOT/HFgT6H
g4nDsyLlbHK2gxUijkJ6ORkRfGOxb8UwHTzLEIRJ5zmkHtJXYM250JOsiukrgEDT40HqdtSgre6O
kXXliGFm9MU0LwRby+I=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ca/+TaSll/KHF7mIE37XMZRKDQpSdluwuJA9x/CRPHNmOrubSxRKoPtbXlxVM6ehE2hXp6yB6qBf
Fup9ZI873BFwgulDsuQHuOSUPGo4bBHwDnNbSi/4G2je8uxqj4KeP/bv0RKunNMT/FTascQdDh6n
SVSARZi75+ElUvhBfAjPHB+yugMvSxDk7TRPn1RomvNtW1CJTL51/PQt26FoAtnxmwYDcU5wo8WT
ATzZmP4jq9ClSvjXHkf/VnlLenBFunDj22Ef6vdvxByXWMZrDdZyqqIvDvktra69BBPdtD2LNyW1
FCI6v17qDRdmShLAB1bJHs4PPkDtQbDOwcgx6g==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5040)
`protect data_block
ZiFiA5yVDlnQHGTKYjf6jdQxbw7Xzr3XewlqJIPmRB1KFMHMr5WlXRhV0l6Gjdjar/PqyF501arE
uFK04oPXO7Ml/QeHzWGkE+GwCMOQl/fT/GHOAZ5lAEM4OSP7McjnDSYYyHraU6XtOeR/a/VUiwj3
skaa0kbxGQBsnBSfGMMvns+Y8Z4PPtn/A0wvAOiIlRM6KLjY1Ldkpquf7E5DGDTpkv1FlXvHKRAi
Gb+m+LEpDnW1hEsmOZ7qBhqV405akvItWWijZDneW71UZpVdV3zYDoHhBxFr5EeT/H7w/p41x1g3
CxaPuSrPF6UBfk6+XhKzRXl9Z7tTruhwimPUikXZ3jNTYrsqh/07oZjkfwCqufPo+C4Vchi/QAsn
ME8ix/aEbFZLaVB/aEVQhIjbglr9qp446mYpD6eL8z23Xn8qm5/lYMbrXHCHrnZjDU76pCXb2syr
CF5z+sHBgEulpWGtsdt+eepGhPP7KhAEO+zPjWuc99w1r80MZzMVemmmkZqg9xCa1u0T+1uYKxyk
jcOF5NMML9cgEL1fma9rfbjCMjCDf9WJirJiU3YnoH+kZerfY7N75W8bvjB6Abg799B4zEt05sfO
mdhVDHc4F72CBJT0KQcKjsdoyk1q4gINrJ3bkzWzLVl+MMYqjmY4mn3K36jtehabn+wGv+2mSRJ+
6wyZdvZqjDKPMP+2w9ptgk8CorLn7pjQLu9rKt788c25edajHNaPclcB1Z2xsSy2j+6aXKOveUiD
323Q1P5k/NNewgUFBbz4ABmuQOEQlStL/R+4pDQ92QPBfXE1f1aSaXqTeO4H4HQqrylUiRyohvTB
HFziTzpyKhcFwewGWZhfxMrUcZBWJERj256HJXEB+oubKHGbB1CmNQ7F9p1Bvd0fnqMEDx8FiXj2
I1aoOY8OXATVIqc1ZMz9z7en3xW8SJVeG0Z9Hw/9STiOZXl/CbT6S3Rqf0VIPFCiKMY4yOblW0nl
h+s+9otjqNLGSZynlSGpNAoUOjJPaZMEWXQ26VUcBCFnpvt33feB6CJaY8hEGmarfyINxMMX9g+L
ai3ARHHqKoLzlypCDuYJlRibxUBJYsqVEE++5F7WMDVxxL7UT8S/sIvIyYxDekeBzk5NIYr1mVhc
sdXqeLKoz+0TciKBmeta64z0Qlnbv41eZwBNUyoksQYpltHjdhLerJSiQwH05bzkmUxf5Zn/NQYv
fItGb7h1P/nK3v0XkHkf1UxnWjtvWBWD7o7kqAjDq0quwpiWQsciurfEBfrgF/twWmAWvGsdwfTW
FPysSson2BiYkBpRdjWvjz6oB5hbsTPhfozlqGl2s/YnJj3siN/uD7rt/fjnpPVP3WInZ8CMWLe1
I6jXeOg7ZxqGivq6Hhqv/w9J/SvhJ34DeqCcRO1AtnIZMptcspcq7Efc4ZI8xJ/eVWEg0Sr0t3+X
fmACLdlRvPzE+6odHNoZKLTzJRoZ9/nMfHfSZJQ03XsOooGmX7jhoJsaGWAMrhAZKFhTMPSb4klK
z4Pw7b+LHduLiZmIJpAzi1nRnVFTPfkfYR6I46kP0tGV9qlFkVKUqFkbzRDORa6RHG4unEd/2Wxd
fV0zLP6rDzu1K/0CreC5Q4qWHpScTnIghoKZpSD3RaSRwlrxxBVxsyyXCro5V3u6qXB7SYKL5+vm
JGwcft26J2QqXSmoGOGDb0dLWkctXb3/TjfjIJFEMkEwEQoePkycZgqfHErLC8J99+V1AUsjHoSU
eUii3MG7eDubTMR4YwunBM37pnZRYRCFHy0UJg7dY7WtS2MEagecV7bkctcJajAQV9lSQqj5QH4e
awdZLWOD+EJxkR1yV/+ilV2D89ObDi5qJ6c5CdC9FR6s0dMIRho7K2rDYiVGrZHK+BKFmH7wS7HS
QYMwsge/7qMx3UDeasR8XFZgsaBwXrfVvZzS8cobH+W0Lrs8zIdrJG80cLNJXjve0GEyKPjoE19z
FmbPptissW8sxnR2gOa/83WkyubcaVkUF6haUR9aLOUX3yTRVLd0wQDJjVtZqqX5PaXV1+/2wbML
eSNP0ZW68bfvHmuvB0X67+5YBFQ61bczQwffOpesyVgpwF18LZzFtafjk/YCV+F5A3xgaHVqBBr8
azvpTbe9KITzcTzg6KvZglREbvhTNvrfiavdxJDaf9+VckmbBLKy13vGZMxrMo06fFajM0riICYc
4j1WvNRUQDthxibwCWs/o2Mcwq3Q6b5vU0dAdMSGI0e2OjyZ0+o3A4WzzW0cyFamXcVnIdZdbZ05
emfgKhSUAb2HPcvZ6tRtKPgtApTuP8zKC7Gi/9JkWhtjEddj2gePDaSlHeactRvovzccVYOKgn8c
yhZ6m513Lo5kVQhTVkDDofIsTcep+csTNN5xKzn7llzyTV6U/w0iJCIFyyZkkL2oQoG8TFd8Qr4r
c/reqsZ8gojC4ncpRvp2AT3DGBztWiWnluF+ZjPAU8kYtcCUQAPivuLqKfCoobp2Yp8cEEiJyR7V
VBf7fUBc+1bUKoxsq51NELq7lqrejvfrs9rbMsx7k7RC/6apoZLGpwL6GIG5wxC2zjq1kpKRh801
szHStf5Juj+KtanwFpeQAsECLFlNIVh5oA8nG0/U5rFY3JsWKWVPM7X3yuETn/jIPRMatKhaixi/
9HKROaUVfpT5oIlAulZaU/6533HZ7YXQ7s5M/wEYDzFmc1w0AQX3IGjVd64inM97U8/pURATnejr
R80t81Z/nND1ObZkDsHAG7R30rds5aqFv86DaJ1VVKEuQ6PH3RZi7M7lkSws641kcbOVxFhKtAnh
8cTLhhj7NUNExsP2/gMM/pw8/3AfVXUdLZXqQwBlg0t6eoGu6wE/1TRQOz9gpTLfk1B4I1DCYOuT
nb4QSUYMG5NocxDq82Wp3q3JZIFE6JyunV3MzOCQ3tUAx5O7KqvyxfqHQ8SmZztB3MFxeUfGDSbo
DfM51AwOHcYVwDN8GxeG2KIBit5526vtmcdGvWPrSyrZNhuTEf2SabXl7Ib6kpgCIjFsxESLc+AO
C3QSOEW434lZVQwR/r+t3oJDpNvMzDBmw+zdfHqY4By7q0WqUOQcM0DLPvxPOtBMsLpo5fK35F0X
B3D6dSndsKmBRGSsxW6HiZvrjkunyYiMX7We4RYgHOLUA4Nm4ByKEZ440eEHZCPylDjNcTeVuAQW
umFeAdFhfud+Zuxpvf5cmxVKBxcgJc41PtLOSwOuSYSVOY+j1pBLVY8+PwTakwUIQyRsQ/79Tpz1
p/2peMnG1Wj08HIvr/ICaNloRWuO1Eto9M2nCycAqT0llhYMkvTAYJTMTr2wQIe4AqdKpU6JZtNq
fogQJO+0fhpmXiUWNWvquGpZ5yi22t+eC+91Xf09rKZFJI+8BpMItbhuRfAuzWy6/AHSVd+u0ot7
0HJvrC9CWWCUnkV9xlHzvHEvTw6h0Q6xlAod5fw6LkV2I76yRtBMew+8DReRfYVIKr36XT3blQN+
/N1gOMGfSAaAYCvxKvU8a3yugMAx5mCUfUZDhnnBi0eE0kKuzpsZUEVnqpIQ1zkXqowy9eddRpEv
hn31Zf+qFMeMelcEuM/DrGaMO1AeNPhNzxnqDEhK4RFVoykcMJnD/dIKRfiMc7fGE2uvURq/e9fa
D4kBkviw6KRK4BbifOfasWoFLNW8WY/VNKbkIM9u1m8OYCACYYVdI71pF0q2YIk4A5RI2lxqUTq/
+YMO4tu1QdbgjVRPhsLuCHMNdXOrfM7B43Qi0mEPnA00eGxwfdBKrBpZqk32xf1h11fchrNFi0lA
u2yRvj7FxJlRPaXv/euub3qnlaSIroG5kYgnyfFF/5v778FWZ5rOjJOGds9NzktzV0Nn+PBVgOYc
Hol+d6I/Pe9+UBwt1lwCtPE7ojiXeAADHRJI4V6HSr1kCGcB5BlyTK/8lE/3wlCt6TTCcI/9S7Wk
eYG4q2YdzZNc2Jukqfhk79/wk/ZUawl8LnyXDdKiqUyaxVQ4s/+8EI7H0UHgdapvFKLg6yGHYE48
39irBM7e02cPNeR2uDf5TrzGoEtc5kh/bvY3R/AseaNyyy4N3ZPOb6R4fJEI3Wkz3wm7f8aXMp0E
aCfyFJgIAsNhFgPOYd8K+G5rvO+NyV9sg9FJPqkMJB2rPsp1L3bmln0wIwBX6KVsz6NVrmVj6VPU
FJfO87PfLx5eeck2lhzTqiFzEZLBrhTtBYh3sHJF+/ZZJiIVtw6fkMf3qi2S/CyAubxkYIyrhwhR
9hheN1FEnQSzekH7k4Nlbj7BMzBbILQkJyRLZPwznqmsMaC4Tu3DzdrraGg6Kivktfl6t1BWF9Hy
5FgUBYIzxmqJh/Kihzlbnd6Ul1OZFkUYS7VZ+qUInJIAADxKwCaGqS4gySz6exr3G8QtYTzmMsrv
HJ3nPXJ1rUFMK9Ik1+Y84tNuoSFqK7A9hXrtXkVIEC4JGsvVo4saLOxl2HTkxUgDTJgwK7zmwk+/
O5qGsluXrBi/X6n6wXtGalhHJhVWCiPiNr0Oxs/fYwYqk4/tyq2sSjTaTF0wfUdUL8101f1xl2PU
3HMW09zJPP+kVf55pD/jkxoL2N73lUJv2b3iVesbDevfQqTdqA1LNwkLg0rRnx6qHYwK9nsDKaIj
6UdTx19E3f+/UJGVKluBT+DhqL9rxoKt5gyc1D3o59necx7+iZlj1a3ENf2c34KVo9PxbPTjCWd5
y4Oub+32YeseubhA7yiGuB0qPbughy8+OzzIpsXdvE/UQTsv0dJJS7uyU1qEIpFK5uaKzPaEl5Bm
YdjsEqDSJty75i1R3GfNcZ+1Q2qKpJ2/+/cHQRLhEMiLC8rB+f6eNoT5xnSrxbAOc1XqBn4fTu3B
eGp13zwf0filitD3pEyH6sVlz25QVf1T13Jsy2Ab6zhAItzj1jjyBQNS2CWC0na6S8gYSNk71PlU
1l1j50GnEIwgmbwEbXRDtQqf8e0k3A9UwneutRBkhqxib9waaiU9fiWHql/40Ip7AzdttQTs266s
rPA/NJL82rh5sLzU51eB7s4OCw5R3O8z99g9NimgIvnMOVBKBrhH+zmXw8v1HG983m+SaG6X1JYc
eb8fZjY7ZsSWOQS5BYdseLcueevL9tHKhxxXTh2mi1fZrD4oKZY8FTpzDWq8wlL7FMOblHDH6cnz
PSYHMIstPQiUHKPp1gK/NMmEip/ZXYorT7w9LNSDOuZZL8NKS+VXhyPFdVpQGcV8ni6/QqAPOqkn
qlp5Emuq+Rl25R6srF3VKp4bYqSenvbqZXH6n1aqAgf1zF26lbUjQS74HUma5f+VCs3ZkSwW7u83
cvG0JnZBQBUp6Ihm4j+WO/bcH77wiSlsU8OfyULktrGlNCyeQoDaPs6Ciqb9Eb7dIdyVKeszra+C
QucXmiHD42n0utbhdazbdDMvRwaxSGjvGmsc7awfi71EcZ3CDXAXFODXLjxp7mHh/3H+25thxkg7
ZbObAH3kM0eJiD6Q3dkvbH5jvgiOJABxSgtxlZUJbPCxufRTiV7V1cwrHn/dHuQ+uos4p5LOquKv
A2rq867SPZfwU9JRzUA0o6zLMobJn18XBTYEYHcBEm0sHgAsrgRR/A8T0hVVLtAdPbXO2YdbIo97
87Q/1fXXo7GU0qWG9zVIVkAqQlvBkb7gtHA7dn17z8AEv6D/KdB4h56AHxLo1+CC1+kFB85lNHy6
8I9V/dBvlht5j9zZC8SDsMpJ8fQ8U1aSAFPnlS2eDqQBz3smBsD5KGERb2CpElVTMiz4f55C1kmn
JO+YzTiBALWQiO2qMfbuCHrcRDxJUxwJN7ssnDIBiKVa8xM9+W+o8ohH4BSI0L1wv6/ZHbW84Vqm
DIIswe9LdoY1eSRM1St9RF2wo+/BSWONO+67KTxQ0Ua6Xbr6xbJi8MZolR1GzLYIE5GgllyqTp3L
9PANQToPzlsFBzUq6/2CPpfqlXsr79tL/hFsF3vMxbbWaIZzpXGoM89O9uNuPArN83f/pKJ/I8pP
/xFc/wQ4daiX+Pt4meYBaYCV9XyUspHHuKm++jl6+jZ/ZfnubvZp44fHXVObm0IFwAyLGokdBUWh
/1N2t1LAHHMrUvLodo0c3/nHWxkmPXyq9nP2bYCjJdPWZhBOMcUakCubCPGbqpktgQHb8FFrFgLm
8Af7VI/RypQ22ZrFMF2R6+UlttRoGxdcb+ySOdunrg0udX/Ihx5Sgb8bfPBytEMSVxS4gHuTKhnr
fUdZI43uzTTUnMPkYj7A1OLiLp19ma/4z1P+dzb7W5wvlPoJK85nLG8Ol2rMtoAm5+GM+M27hUyk
D0aqX/2Gei1uw6zVVW91NNvfnSRj5pvvi5LcCjT5Sh5AzlQJBV9g7HueJHT8uZxeuFvDnQl29ChE
C7+PaV/Dz0rpFJi6fR8IQhqi1JT7+5rY1bpfbYMTOz+kA6DwnRUggt/WdNmEu+TvCa6RQwd6HPHi
+IgZ6e80KHzoWA1fjmd/t4BmnAlK8HoX5dKEpu1Fa2dXsbx6w+9J9I3ZXOMJvPJJfqKqeovHylWY
IVHfJRvuLSSaYbNo6x9tqridhKPDW1bVp2EoSWWEbuxNUFos9ujsubgqjowjMnDMxQksf7I6fq6S
B+I2ki9SWvtp49rh/3rUbyR/yxat3XxTRp6rq+Ndq+3Z8oRk6j2QftE600FI79o59irGbFbFwQIn
E8W3UNnWt6URLWbsR/U7LQKCzngQ8fld
`protect end_protected

