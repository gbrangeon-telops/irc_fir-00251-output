

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
nqqBtmqfflVo0LfdOWD2OeylbTCJPLX6XaSqFQpCXkHX4TF1QAXZspyiDVaQlwRkat06cPZ5E411
bTzbr9/qZQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Q/X3qbnpTyRXgHhmurX8chlDRL2XjwnbHjo5m2aoqrTNSVAUPYEYGIGJVoJhRP1Bd27KZbGI0BFX
fZKfju5H4nz84jXPUC/rcsp76WTu945qoXwdo30XI0Qhi1w21P6EhLXccz1l4c9zfTwlHtVuYV2c
xkxHRh0F8KrrR61HDHc=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
jBFh6UBl2pQmyl/KNdwY4r9ld/Frb+RgwTVitzK9Y6Fp+6xDwrsib4d9Z9Trd2PuW5z5/ot40n86
vR7VZpJnONM8UmDjWgdiB8rXNXaI1rBfme4TQ3jj6RaF803c2cAi4cdZ4qM3X7V29W2B5HXbYsfA
+fn+v+caVjEUXZHZm4HMyIR7TNVnvmCWeeLj52d+u3MrD7UjjkqtqnRWdy0ckM9p4TE27eiu/nsz
awiAJoiVLZNTMmdaTdZ6vB/sS67SAe0JjX1nTwssfK86UYU1+n0NLZ+SLB4lkqxmhepGPNojfE8p
9hJaPKOTV3d/umJbTV97L90iPloNPMXpGK/m+A==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
cwUUX8orCEMoCaO4wbzIkA5h1G/QOLlup3/J46IxMYEEhFnVuE82RZ46tcCa958uxg+L9/l1SnQ1
1Qa6GFDzaEz3zEcSDS+t0jFMPNI7VUppaIgcalGdkOXBIX9fihrhASeWjqmTDrUSlTt7Vzyo+3TY
n3HFHRbTrCchXcVswqs=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Z1XHzIMnint6AvJuhSJyN/+kraiZwIT5ZFNyZxcRS4ee586ZcCrsBlqjvo3awgeNWb2yZNQKbtJY
UBJT2Ww9PtMdwpg4MPuZFMCTECdiBOLjqX7gX0K3iBdA+35RXRVkpnaon7ABi2dY8SU6a03iv3ph
ed9P79UVGmdGucbzSQNo8vkiW9pS6ZJElXKmEibSc0C9Vw6VmCNdLosnrss+vUEVkPDu65r8MqDO
9/2zcjIio0kfnpSLOaIDXqGefGNR89nRv/NxKymzLnDjvK13FSfKq6qNfA+cXOtnv8oRuf0tdkh7
e8F12j/LQajA5bXDfmPQ3bNX4Qv06vuQ9+MAAw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 89616)
`protect data_block
S4JddA5BznzXyxiV3gk7ru6Zfd889A3j3YC5mbbiz8tlWHa8BS2M6G52yu5M618M24yHyiMBqKiA
oXu9jIiGSZ2i09As8eacE1a0lbXxTDhcMKrB7fOZchrv9mv5z9Fap7u9BWCdTkDMhcWrdtYDbdiH
11uXLp1pYJB7MdCV9OYlXPmOvNDqaW50Cvxb0iQw3WOzzI3h4PcHcxf61u/cc8NoHd3gh+x5hZH2
s+drs/wRg3xGq7Z2kV/Ezf0Hy9Mjn+5vXDyORmHgTStqCA0QT3RxHZcFcnoipX88JB4lQsDHZPkL
lfRobi5wK5D7BwvkegHLRh8YTV3LXdSohfHdtWvE2ALICmE6c1xJMa4V8TwCfNiG74T1uZ7IrnRN
MafvRT3bSYIRFgz3fF/1z969+oxxGNLBUaxiHgKlJbvT02VNmUCDbBVJeoTbJzbRbfNdjqwdRGmc
FYvr7VoslfMhVNGvgwtTgq+BWfz0ZHEDEquC4+3HvOvDdtlbATbWEFc1HpWKMxxLrUMiro2NtCI6
VDE7FPDaOoPDbRNUnROb9Eq2JdPuZt/x9NGklyqsTyTzNklsWAiYFAQNfeLJKsesiRSuAjBA2Awx
H1Bwq8QIQp/ggmOd+uaLOJkXBw+ps3f0/9G2c4NbQrT1Y/qrrD6XQ1Mb5i6P1Y16RFRNeivjxBNf
YdNl2u6PmkzcPLhZy4r5DcTfQlXh/b24UEYb8Bf7/Ag5Yt91g4Ti4yTDl28mtWsZCPLRy9TEb5hA
+tPmhWvTvBA/sYDX06OpPOQVxwXYzyyULZAWv6KDEMe72v5Pzfc8socNzM0U058cdsfyaRsgrun5
BP8P5IhBk/bQezEJ1MjcPjheDOFrFayBOsKKtC6K/QQOwJ3rF/ovWPMAF4E89kDT0c8soBvIh/ba
8TJe+LibcT78eyeGLEL2VMpwepe1cCCHiIuQspeqfn7/kCK0eH9gHKbIkcY3A1ZxkpqxWpQXecyP
VEuy8FO+lpDJDjp/FyRidGu8hhjmRt9O5MSohJ2jOqr2Q4ZU96js7JtKi6/z4mJQPsCGL63vxtH0
2BAjnfh3rtgQ/c7/x5cJ/GigogNZ22Pg8xX+gjGh5Gju49CXU00pUejybnUSLQK5fxO46ZH7q8T8
SZ0J/GKIKwXVtRRfxDZJkkopWFjsmqCTLMCEYbKF7MdXdbkBsIGNJfvpEC3MCq+TuNJatk8TwFp5
59iQGuKKU/l1iyKEXQuGHihcv9pcGqadrDE0E+viaXYhFrFs2WLjk/rAZPWrZLvYmH7Y0hP038ED
c8X1fwJ2Wp6INOt4dfi3lRr8LVCRdVbq9x3BJzqrMY9s12nva2lF2VG91Z9zKkSe5DkVxX1AukXZ
hOUg0UyecpddAsJjmhOnTMEIZT2c2YiItbe5mWzgP2hvLOlXJB/cDlkS4ft6Og+IFIGH4ApoZl9p
o7Iz3FdKhhSULLgb4nL90Ke2cxq1xy+EJShzVrmnLslGIn90g9IMnJryjjwfHpT6B8/tdUYD9klB
ZVbH0Z22k9CKXbcEb4fGkxZLKWa4wLMb6wlKzSRxxzOwD0sBO7PKIX/wpIrY0HZ1imb2Q2o2X6SZ
PuXZ+VrbFATChCVjNmqnLiw9T8K65Y5ABkoqbX4yUdlhnBJt0garwBZUF7R+fba4m0O7B28nikkq
pysWfMPCytPSIfEm7sKI1aESxoa1NBDBDe8DWBtgO1NPJXZy7r1+ZXfTj20IRO+tk3GblytnlZNz
3L1HR/BFMniAgaGCjGTOQhMowrIz23ylGmhrbixmPIhlhiCN4vNCrIC6DnVBRuzJ+E5cTdBR9sK8
bPw1crFGu4npqNTwPp1vOU0s1YILf2URAVrRqwTbRlANG4LUIBSCJNfa9lMILjmbFtMK5nWablmW
1YCeqoi6LW/Y4EcHq9tR+D+xahPmvE2kXMV9s51vqr4KGb/uDibtMcj+Wl2r7OYkj+zx4DkpYMlA
T3Yi+0MxCm8kS1goyk0nWmAlI1ImR9tqP1nxqfnQmt2SDS6+fdMT8b4Wr5/EXod/xhYPvy95/908
lkWwiBksnOWk7JvNTmxSjXXdNM4iA5bbX4yotMhaYMvwyXuFnlnDdBcNOoKwPfPX48TyZziONfJD
K8snkH+CEWvpff1746l9McRUOXfIpvWI4ijowVh9+mtpclBkNH/q7ojuJHQdoySzaqMxWueys5R0
QCrcfOF6X7cJPM1QuZtYu0xLq9shBn20VFUB2tmp2WcGMa/hv4MQQcXi3+VUDvkRbzX+ZRgE6QeS
Z50KqSSG8OXY6ZQF2fezqjLGmrGZJYzeTxEW/XMyzXCP6SgWbdRQJx5q6Sm1JpCY4Mzb4X7bMmPQ
o5wBUiPsennYmd1JDy7YonVIS3o0AvG0HkruWanEQxxODOfljWAtwIVf1yJQdHkYxoxqx1mqqsPF
XDSRzSbLWySd/+6Lw+zs8x7DY1tONzzPZaBCmrm8p4MeJSUoeofFLPT5PBibH26RNqykcZ7aXV84
9do0x5/iu6uwqcoGD+TWvepG84hC2IX+5VEsWejUhl4UqHlwfvIE3q9ZD98oqUFL/8p39lpVgx/r
M61puFVxrOL++nDwmvewhrNVB/fFxyN06H87mFGgR+zuAyLmbhzXI/V95bGkdu4UIUmSmP8wQAFL
J8BhAC9Hv38rum7NemYu2fEn4YP7sL6CXqiPsSbwo30CscV5fJHXleT1HU4nOL4q5Ju1zu3YEAFv
R+P8ZUbgYXfwqpfIYT1Ce920aQRIZ0qOGpen0uRIWOYuxvI2IW4ZnkX6tcDYip4K66Dk7tZepa67
R9p6BL8S6SGh76TN2wKkJD4bzgMzm5xj+Li7eYBiwO8BtAYCmTP6b8Nb9IyPkApCLwpMhRwcMb6l
EU9Z003tqoQARhdVBj8cuuWrPAzmOP1QotYMf6qMePnmd55Y7NhSs0d3Ez69d9dJMPHbpJS/PL9D
Tzde17WebYvPpg0XijJnybuH4FOx6SD8oMIFNeQue9itKFLORKso5BqHal8/9+fZ21tKmu1CArwH
UwL1kHIFYpPj8W5id7qxFelmUIKmcI1sZkIssoAdeh+H/N69Rny8J45B/OJwcFfyAoFKI69ViTbq
c7tuBHXMOsFeJsrpkL57O3EoumB9X06KlqUduLz24oKfZjnJqhhbU0OcCJ6M/0TMzRHBba462ILe
y7TBZ1IiuZ94+BUjm1Gpk76p/tr2Yliu+HaLvP29O8eNWhUhNAzyJyTwAqY10ZTRXLBqjTCA4mPU
iF6YoW3UXLsvD/PJSQqh9Hv63BhNimAc1kzv6zGEES0sbag2OrGOoo+48cLKNnwkocIWJlzpYbsV
Yfxi2buyIsXy7rFLeBdrx88GOhV4h8ZCkLK1tbbBhcmW2TlqAkogql4ssu8J6WNTSXixV7B73vjL
+tK5q+ACA03Pc27Q0d8tNmznISWyX7cHv+qwrlBGsAVqAjqSQPcgI3miJY4xe0wm316EUaixVeFQ
PDnDhLCJs2phPGIudlJwr3jr4k1mTbIo1TqzuwQmLFXR+t4NmRAPcLve6NOJjFuKwENhUWaESgnh
L94iDCOE04gXbJynwEmP7LQ6R1ffKL4C5H/zJiAX8181dqZMdLaiJ9IE4GpHMViVckoxRYZ0SkoA
VuYhI/no+BK/ekAuYKv41k9V5pA+jTyRI0c0oykavKMR/R+HNTbMBBDw/87+zU8rm3UmTYzdH4pZ
IfrhXqP0QvEr0Z8HBV3p2AGawHH8YAtjSnGZhhiRiOI1hMr1BMN3B/BJVk9rRE7/WSaaNV0mXSBf
iWH3MbPnvyAimwPwl9ElMFVmOvJnEW+6qRF96ci9diKOA4K85Z2a27++PCVY374q1RvuYBxOXSIc
aQRSdMZvhMWp5V1Khtycz+G/hCHeWyQv1Vi6j++bR4VkzldGg3Ev0nZYdlPxPh2jK9IIucD4IG9C
UTOufSXNpl4fb5AkzHPhsDohKDmdsQWwTI2D2FV9BRuk5MVGpdGrujsJMEKRONs3osR4AEgAPGqR
cmgIoJ/Aw4F2ZM2WWFsopUaapg5x0KvQYSX1Uo07S7RLoq1y7JxIEohXVqcjpZR/evaR18fNH8km
Tfp8ztxlvf1+7mkvPqeDRbBKZ8hIltNPO3F3wlBRQ0AtF1ANHSsxcsQLKDiWDwgQY8h2M2cQMXux
7LiqblJqWxfkCakomovPjU9T1Lg0Bnq2+okplDdacwrFN3KyKRr2gabbLxtMj/Bn4f9k7xWgJP9t
z1MbV5DTIL0DH/U2d/NKkaCvJilGqS9uStvJ91TNDz55LaGEl69IaUVG0mARst0pIedu6t+R5ifo
e1xy+PStOGFu9Yyyq9qROPwSV7rItd9ptGvMkaMnZCz/sBlJVBiz5P2AGp9ns57CmfpkAl7PoAbZ
/9XaQhcuWACuUJVIU/Rmllpseq3dWysfrNVpVKh5J+bno5ioQn/daKSdyGUABXlwZeaZqDvV28yy
2J72kBiTszYc25c5c8bNeRiXO3VNJnowK5mN3Toz5ZBWozSxDfxJ7VNsYZ/53TxHrbQvMoRY9jxq
9ybf2r4bHCXTJkUvQeCnlemZBLPZXzTj7ENQuToU6PhqHtIevW6HyJ9fVZndTo7KuXU7Cugrb6Ft
Br3I5C7hVYd4k/zwndBsnHZc91L5QOGWxezAUyRpKR/1s0ntXiPvlL7834hgo4cZnjQVtsM6Btl/
8r57bSh7bDJbBExdIXyybDQTeAF2NTeNPtJLh+M55D5loivQsNJqcX1pONRzePEPMsxRVqDQn0HV
Qc0Lkzbv1vy3CUUjCzcIGmZI0U3RfJ0rljp9h/bJPyPrs20SKlpCaJTOhqs5YRBqgUTrh+f//hN7
X8TI0dtJdQA0VutRJ7eMwXySG/bIFWSV4PcyIbTKsOyFXqu095ZmFb9grPlR9VBbu9oxz4OUgvS6
tZDJN+T+PzsM22yLMw2uyMmne1c9FxKqMm4dlHYIVpTmsgpT9V2dkq5uuX7qgrkMTuL00uosVPUF
cE3CPM6eWcf0587asVF4+eVBxXT1sBIo6v62uD5d9tyz/cexqXco2zLRZz4G1go/eGPE9HmWPt0V
hYqbGjwet54ghO4ZzI/v0IS74yY3K3qVerh1NpAjc8vFPoS5i7byg12/4LifMM/nWouInuOCocUI
SyumfdrpR6wqaNMU7xvk8Jp2PHQJxZNZKOpPC0r3OnvSj5mKfbiFdRAfcSaiEnCLEJ6EhM1ADkv+
Bzhj2OMEF2vV10P9MrVF6L6UoIYlmhIzzE9n5cQaOfOg2sc1Y9aLN6iEF5v8sHnLer+ga8wfs3Fj
mrtUbuV5n5ZiZEgjrGcDVZzyoD14dg4tNDTDYopa4gM2B+zK6Xok6saenDgLABfXri6p/mC1fOjn
iSFkHRTPFZuZsm34gzvEYMoOo++IsfDORg7Uv/kQqCQcyvkHyX9qaRnExS+jPsdoUOj8SgHli0l7
6LWr5m9QUjYhwXoxXMs9lu5GjC4oDYuzRlvj12uqVVyj4ibppVUbSv8Ivr8vQ7MWk9rcAITiA70+
/1ysMwsnkIXCFzzJvv+49XUac0v7SjweB6ltLRDoKy5lpLFFS9vRB72hZLszanyniaJFJjZ0/PpO
5VqyOmn4PcM65OW2J0IP6VntqjOBVLFZ2P293EnB0G8lNovde9ZkBGmYK3yQVl+JCUdOdkJOzg/p
r/ZXQWT3xorqwRVguXwMLyT6P8TQT5avVgJO0sOvaPjMezf7KyXCcYbSuxWwaiWeSwGXJdyO0YiN
EnvngvOyu7toXTCwuhsmSTBEdgicbyvrtIDjEllKPhQ1aTUB+OU/qRspUfAzHwtZ7Q5AeiFw6ixw
KWbeuwdTlx1cj9rSm4Vw/VAUy24XhR3f9USoZaZTf49tbYALsmDDdVDwEKqYaJ99hUI0bFgfnibZ
HjM4BRt6AXiMWCJ8uWpIdd7QK/NkXx8SLJ5py4LCLH3if7XZgyVJSqs9GVLI7IoTi8X0b2FKzfJQ
HHXggz1WMR5wiMSlsaQARy8tHhF5qcAXVhqgDk5CR7LTbgyKJlgB6EflS0j943uiBzNK5B6t7c54
8vRNAbQ9umOpoU+Ny+VmcK2r8fKgoTDyi03ASlkwUlTskEzCc0TM5+xv3z8K8C6InIb/HwiPMBGd
kFIMeZV9cJ6DRlRE8cp9cfD8B0ke2gki/khc/O0VALvf6HFF68zqTXg3gG5vYpGBa82EVmDN9OuT
qPxNRCek8zQpEtxJrh3MKOlqSCRikgNODs2xA28Hs4R/sa/b1MwANID4CCIO503epxeFhTkPWsDJ
Rh9S52mYnQ1YEi+4tOemOaULcpkLdHYZm180jg7URM2bMjJgiV4gAXgpa4KkM0EeVV6v+0VdZYPf
H6EFuxDOChV7GrUpePIeAWRKzVEtDlIC4A8Lw2AY4I0FZE5pfkJn89+TmhpGDHMqSYCPJXg7EfTq
2zy9mtzByf2sJBXeDZMG5e5W8iRCXUEVJ6zpEWrbC0+Gcr4FaVuuL1LdVvHa1z57ToGhnOqTHz42
jR6ggyaSh93g9LmrRdBxSETx3G6Leo3Erg67BJnSFkW0/KD6jRkG8fVLLDeDLMLvpCGFtSZaW+YJ
PP88JLidyEnPGSmra/wnEycFIeeLld8ThSpIG93QZNL+t9gT9E5mA2ANOc6lF++llTSyRU7eCvhm
hJm8hpxwUH4qwIK8yFDt0AhZVRDs+cwm3CioqQYkcG/JttM/7bTGXgL7gNwGBNsGetr14FPfviIx
YhCvqoJoO2/Haqs+vr5ljlVv1vf0iurpRm8eiB+VEAZFB7w9RC2PYSuBOAkdVrENjlzxhZROazbo
lv9jtrVEwWwtNgUXiQiy5OCUOy0p6+u6xNpikk6WvZw6BjtByTIW66WriClJPox+0VGPubsdlsKO
kqkaH5HD6LyKF2q+XlTjG3qexSaSski0bjzFMxoQywUxjnvNv0gSasSQsUhQie7weDpjmewok2lk
PHycLXpEv7vAMVq3ne5h/UU0JHhLxmyErgpQTRAohmsJ47kk3cbj07xfNMa7Aa3evnxlIA1bz97G
SffJOz+cyT10GIOKhmvfTzu7e4YCMfeXdBpAM7GzKjt549DhIhvan9qJDzrq2F9KmC7GMjaTFkmH
DYKzBPP/zOAwyrSa0GapBZKVxZnODa0fiR63UJXT1M+mlBjj408uy9lju730Vj37wo9JjlYt4H68
VX8jY4fSracbnrDU8LDksyZfm6K7geRg36KZ9QXKNQwTVLRcnumXV6l95YPgsfdg/9SwnxBjsN1p
ZSK7k4FskVZXv2Tgna6K/9MzxUOQE7WIsWvI0WM8itvikOl3k1e90MPU4+usvvU8FxL+FVwmFLSn
9JI4wUym2Kom4WBb6jRW0qFVFZLWatrQzWnjt6McdVHfW4llohInpTmUU7AOQ2XosfDLEw0vVLhh
m1DnFkgppBMw382kVoNVVKDuXO7p0PmaVowkH/xHmXj4xDOvwv79N0//B4sXYq9tIR+s7efBGPDw
ozvxM4jXWcXneiPYdzaX5XI3BG3wKzUNdsK0NlVjUM/UdPMev1HlPkM9RPKzkkuXFYK/4l00YER9
AtEyeP/mE/PY0esPvK8ppK7bipsmCiKeAnIpRx2u4iM6+uySpsF1aLAH86MkQPUACqeStfdO/5fg
9jkTZvM6XKz4moFWk3MVF1EvYLke/6AV0rRddRReZY3I5YXytnlpLqqTJtlZVPEYorCtlMb7HaOF
8zQ3ktfvKI8q4TWEqKIKOVCyg/Ww99GBPnjQP9eOCm4Tk0iCxUhW6sH8mM/67w5RlgDIBHvmwQvJ
XuLT91BqCOjNb1DUReiHtVDqKcaD9KwT9ACkYJTvYGZeDlpa9GuqhYTJgOTFCDoM1xsArKVpf8Ut
yXRjkOH5TXug6FH9LN2fpcnPTC4JJOy6o23Rd3fJJ1NqBBo2z9Yhk4igP7Pq4dtM1p57RJXsNZgW
Gxel9NWgTNTuncvflEK24fHBJnsD+lMWTSQatGaKs60ckQyrMdvl/o/katITstwWDoanVBD9qxwt
OQ07QCyHDn1HiB9asAq1xrK4rDTY76HXkzr64XjXfQEbn5UYDGyfzDlYPSPVO6ljhWn0BFBA6nBs
TRLByeCs40zcx/lHEwNjRF2hntQfB9PriX9yAI9zi5TEGHsXlEeMmbcmwboecRQVx7Na/JfT249k
1sSi5C9SRiPMF2EaQW6CSW/FqEgHFnMYI5fdmMgvh7opa3YIcRYN+SJvPb4wH2azaHXmPjW/kuHM
IwRxo61AOQy80LO+BE2DXH+LFXgbe/mdoDlkuLaxQo56SJDaSo2ZyErXN6jr0zqB2W3JWtzF8IO5
JAPfkPDxIS2Ww/5WVu0nHst3Wx8/yyy+zsZDYTlBgHY33rFvUeeWgKwE/IbTNuVZy0xq+ggq/uNI
S9AW3FKiGh3zSkz+DoIUPNLpun57yoh2bdPrzX4dHWtqy2v88btOL6xyRx9FlB3CoR/m4ggPeUYB
fA08hH71Uc4ztENBD6g5T38Sh2Vg2XbVr7FEqxqRquCjnXBJzeLz5beglEKGaCLmRd/Q/HpCC7+P
TAQvn2HU60O/dqtQCRP7nheFDLQ4V75HDbXkZUHogMJdmFDGuwFiG15EADVVVI5hxPskH8zDMKb0
AtDe6N0gqKpbi04i+GJktTXOrv1txWkejS1mToJUtpLOidKl3JDJz5lvIPvEHerAXAj74+ybWDt6
GhiFFw+jGYx8ejNIsBtdeUK8rVRHbB3KGl2sTiLzfVu3Ah4ny1Xe1u7nyER4ZxZtbCF3xOEMRd0Y
78e3EqabnTctLT/CFSKoqjfvoVsEgaBBFPZMfcoCGjTByje3IoP98fSSZyxpSrCD5lcYN6z7plOC
AscxELD+vNR4lx2jkMJ8RpYWAtJULKUSoeBe8OzYcbLZuNSRmXU8kEkQ8WRunlZV94rzLYddvDW7
7Di8y2jFpSB86Nfcjvx6aNBu0oDjJ9p5cYz4oQf5m6YLdGfRXv0gCOMg4SQrM5e4CkfEaNgGKHlm
afTmiKF+lMUxwqFTIGWOlte+HeAzT5x4J+Xtdz644EVpAxOvcW2OVUXZbMzW7n4i3g40fNQsbCQh
O9Cwkt0dB7cgzrL88MTKMtzenk2nHYiNGytaXsAWL5dDISQ0GujXVlagh01WuywsC5Vxm0t+Fccg
KP9jJfRXkuuoKaBWZGjxvZ7n9qVV4N9tVxPZiWudANLfr4HXZhJtpqVnkymP/A0lMjCLyGD9t63I
YGR2CSpAs1+d4v4uIyB1kozfAd93R1W5yv0U9zBOr/7FJHFE522ryLn1q+aaWwKCo2mldbUMIoQe
xxdcROW+d4D4DDUGuPH6rsSqiRbJz/oaOZYRDtRtuprPysa3QYIfb44SLKHFbG7kuSAHHGagKoD2
1DkVS9wEX5LeYczff5/AhrrjQq0FIeKEL1EO9ys3zGOp0zKSPnRHHI5R3UlgDHA453addo5pN/zN
eDo6U54yC9m7o1aoKty34HG49WbRWF5Z+SuQQB2wx3zGXoHERYHDU13FvXVTxbW80wOa1LVTeN8r
5aQWOcwS8u9eSGFADPE9J3okdQKhlzqhZ6LJ/nmYow9zc6Byy5tpmzIWjB5BzBrU0TCAxPqyd22y
V5eRDFA9zv7vogxmgYxFZQ0YhOyjX2WtW3/zAFfxo6L/qzEVZUI99E9NtCNUViuEqhg9lfnddRN5
eAeMN4h26VKB17P3JJ1LvPyFZQpLmJBClHJm4Y/H1kaPLpswIfw8D9aSsZfJjjrED2YtZd5rdSo9
CeHipzfMWl4u7DeW5BmyQ402siTPmGP6bkntGTknohwNZw3MwSQuILf8E5IGDDEpSnIjqxD3plHB
GHy5o1xRgHb9rGx/NkTpwmdO5fEsgurb9moP9Ge/8+AFQxx+o+wVgycCnEaRn4SKfvmsU5KdIJtk
n4HIXUvUkaYd7NpAAir3oAdjOUU41z72EZm+uEv4du7O44ktux0f1wxV7fCBl/VoVEdE0f6l6Z4W
0yQ1fZ51PswAsema9kPiemFAW4rEc85M8oqJQ9hgNEPwMKNZ5KHObe13QKTpmomTMhEHWyFXyvxc
uLqJlU9kouSF0LUmyGmpB2jfoa5D74qGIRqMgHXEQA7gVGsEtbXpi5R+DBewSc1ya6z599mFR5lB
ccMH6YwjOKkG2Ft0+j0fcenqHndx5EwefhBx84HlQ59U4suRFjp1K7Up9nVwbrH5jEWN9a6Ibe26
P3IDS2BVYSUshtvMPXbTwko3Renlogc3/PQxh+NEK/Rbn4lo86CSFQzm7yj7Uz/RB4v5hIWlzrOJ
T3WZ/0Z+o+vyU9Hhtzj94gKoUEC3IwuYIBmmdauzcVZ6Egp1FIXd/ygiPoByJ7Jl9aD1ZFw+2y2V
L1Y39wvOfribGqYXimMKjyLg/gl997igElVxIktIktt6XTbGK62Zduwg0aI9H/chMAd5ZdE82JOT
GETNqzfdq35F6Uubl/M0mb44Tg1sFnCcaxE3n2f83NnZ/TVXjs9TLjGHJVIHI/ko8qeeaBTlUVBz
Vnu8EmDxbtHOFSnIHvpUeldwKLRa8L3lCKwa9HD8lI1DU1Q0+mfg/qI15gQ6ClnfrjDB2onhaZtT
oGan71M67p0HagjL3GO9Eu7EfrZHEO7RIWsTo0Rfva+sTZl4qSL4eSnHQ4bw1lzgygox3YMG6oEX
U8nGR9hAPxdxpsLMTgATo1KX+N71szZJBmka0XSXmCVc32AKSdV9OywgSQRR3EAsnIdeJ0zhE+D/
DbtrjIMnmq76yaLMfa61jjty28eXBRM0I/zxIj/HAqrE0VOjsTRM+KvcTSZ/UjikQmqz1c4sLb4R
yrhjA7nntkshVQ20RCyG8rk5mXnm51K++Fw2G4zlrkj0byes1vHI44Icz9cJOlV6CLL04Suk2WjC
uT5pr0IgFkiwV/xlsUunJpvXS3qIiaxpiPGFtDvoYpKpaI/EPF2RE5WpSV1obSEVaotdweVbISQx
ywS4Ccf9hDvEoo6nR+aWI0zDi7WTsADD5nt0CSCDv4BjP31EgOry13RyATjzWPk2IwkiDnum4VXq
jXvn6eKIrkmO3yM+FTuKkGzvnKlJGR6K/qaWk0LQcu8A7nTjEH+D0C8bartJ9mzaLI9Hcff03HyO
+5mgl0vvYIqylfPahFUfB/mc+KoxC6TYxynOM4bFsf5XV1tAtm86Slf8IdpKHD/A6VtCQjkxiUDS
T0dMY71FeBlusDILL6NtDWBJzA0liY9BzpEyiJCNvBuyIjNjdjZ78JaA13IW+qBySm0nyXc9IMXw
VOcFOIhOKsbSArBlIm/ou2ykviU6hXAyTPUiIdp5g9o/s/L4BCWpHI+D37xs7eoy9ilPcdKP81Hz
X0j3FEmH4hTlJEMrGICzXlICwrc0w/ZENA0Kf5C6LSyfrDl7ve20MYPe6RPe895A41PbnSZBiJNf
s+KpHd8fbws8AGEIFxx1E9nD+97EJcdhDCK/ibvTG6zda/9ZXfGJih4bSaKxQJ000yzsR+EYN6Ey
Pivvqwia6zx/93ZCOMZWUKBqejci/9OEtEwF+l9uZcwyYPGQSpSTjEWgIVg47HQtdvAyXNv3+mur
UBcYHab1IcLkhhh9/NYcAo7PaYcgEtoJs1EWHLVnoeOMQBGNoOA+prQDO2wWCEKZuIe0/pvb948Y
hywNtGZFUPPpnf43g3I7JvbEedW3QKw1pClcTP7k4mCE6PhSEuB6S9dvAesFYRbNBU6yKzHlhNc1
TSaBevV1JfJZVw2u4sTOsYvWbqlRnCNqvLf2rKIuahmSPPO7Odrhe4ztBYS+Xs5Bedktyu0qxaCu
HTjHpuoEINf60i6HPrViGCFu2OigKY4BAOKdt+XOlpm681zWBH0OP+OR2BmE7cqb18FrKBBolUOu
it1ZGgyJgZpGG5PURwR7Sly2HmdYIlDLx0l0c8NWJXMyg9Y4YoDRI7vqzeuX5J7/b4F0WC0ruzzY
VkHrWxn90Tc5YKdFc9jA1lHWz/vEIc3LQxpPdzlCN3q9UgdJ5FV/BJMr7bh0hxVTz53Zmyoc1CQz
XebG0P0a03c/xWZRwOS619JH/JoMBNMcZm3sf4XKboXUS8EXzVM9qvbOZPcOhjC9GQ5iTimmewx4
Ek0Y1gDxt/6X5IU9hDC/qZBlD3ffrKbvaguBIMnHdkIKLZeMfqtQCuMqlAIXYXBFtR4FtGDw9Sph
kAvmlGC0VirGcfQVjU3ZRD9McpRMX02UpTenccEx13OR4IBo1RfcvbX06y0PemBk3pPVis1d74EK
NN6hatc/W6SBib6vAV85k2sfa6JNqyi3u0LdaR0RpvTL8pP1xgs8dXMSOGITM9pCqgLXPCpJfOQo
tIB218wqztnrBwXMaNI8L8Kt54QNO4INJ4BFcOL9NRJz5DBJvgT1fPWALzjMUrzHy2CaepsvLzfB
qINmAA78uxmB3fwWt8lSn41i/dHbwdhSZPrNCay3rQUQrTu/N7bZ3Jw7iUU//khf9MQ6X4KtUKF2
iVHCPNB3L+/ktxN7NG3hWctBmUkPVbmUpP5dxZxZbZnmrm8lQlt4AXnRdIoyk5J245IFEO2uZmNI
2WHmrDc7qjng6naeuII4CicEUTsXAjUnl03t19WbrNFagnaJnQuij784qGFPJ6bku25cXF2g33y9
VCUS9z/nJIBXJ31b539DD3QkzDUTO8+hbNbkOx0iZHyLYuSL78/jjFUk5xM6K8AFEOgIV54Q77uO
QRUlLzav6RXG4J/dJvTLsEKFaDKzQCkscfQzKeq4BUcj1hhfPFf4TCnsURfFbRSWPnQK+jHlfE1U
9FAR5B8fxDolsWPOoH+Y4rvg2M/+bppb8GM9+J/JKH8jFYFK6mFLW5qzqZAXQlqV4o/QFezp/oxi
X+WxifAy8vhW2wLaoBf0g+h2r57g/KmvJF9439LekghpjdJ8Zc1nGdr8dF5Dso+eY1R7KkjBnxMj
X+DOzaJbD7KoeGztRL1Cb23ApEsShZo1NkyyMQ1EOgKN1kACvglMvEIM0ulk40otKuioLigaJEdT
imgWp5/tOPi3KktvRWUPIYjAZJ3fNXXXn3qPzJJjpBUADKeu7SnEFczBi1008fwn4/tkEkTlu/Q4
zGuZhmLldG5375bN+mZ3MmFBsPFc8Gvo7k6EdjtgsARnUHd2+lMS5Z6g6SgxvsimXX9672JJ5RSC
NTUx1UBd817WMUrtdYdrhZmelJH0pVuCG03kKOUIkixHXRiaU9Z+dG0IlIxntX6OndbqNGYUn1ns
KIHfIP+uOJLR6MUi0u3VUXs39ELla2fRPNp9f+pk4yNM29oNzFDTjgCmH3hdW5iCnbJLGZKGW3Q6
MtTk34+6bwo01Z4P2G+CVkPjDtUWUuePbRswqazT/BDG+w7QP26b3j3BnNQJ6d5t2ZJ6SyWPhJ3g
+20qUBWAbifnqrzD50X4ZXlLx/o9dw/GSZePTlsd3Y4oJLmEA5YTJ/c3raOJRf//cPSLNz+wCqWl
eJ9F/dpnabt0cSlni2DfDl6Sof8UOe7XmLfBr9FQcm8UoZ8SAqYu42RMOdw2IVlhqiS9822PDKVz
kmfo84AuuGw5vdSvmnBK3yvRswwUUqpy5R6v0t3JjHtHJJ28QxBMXczJTWQL4RHp78ieNNmoO7l9
4Q1G+gY805p+C00ZaSn61tk+hM3EXfJ4tHMy50+BsjfzfKj4H4mfgRuU75edaGquBdG+bTDYo15n
gE/ZaX5APAjDdF7RSrvbBZ867kDng0oTFSuKXFNxp4gg4NJf74PQYVNoQHXBaeL3WcoVrOOWpYhL
tCyZz6eNUVlJmz23EgxL5Ccglh13lCQEQORoTEvNGiIo30kXssAbwk1IQAnYHKr54UNidYaGd0v7
o0lCwteGNpfWlg4MD2MLWHUtBGHDQ9kgCQyRECZeo+qctCnGZQV84lI6JQr8Yl2zcwPhxe8BtSC1
frMX3qJBuxJU+GE1bthdOtQufIP2fyvOit1Kuyet6FeOANgl1Sh1TJr1E4Cos260jjrLs8oJfa4c
wApnrZKrU8tVwNt+vW1Iz6ZEdkqlyvXbn7LX2+gaQ31qcVxiVotg/WymM/UNBBxC9/hYHPWv2Wx+
NWfuCysEfZoKbhl2MHKEMgWWpCNdz8wT6Mz+kXbs1KL1MntgDwTus5GliVeM/IoJB8v8aiPjrL+5
i5rnk0tZeUbJuprFmJYcc08FwrnhzVdfIDN/Vx9lev4EkvfsTJoFRKXU5CjqKdUGftlDzcqbRB/e
h16SSuky0cLMNbnlaGRiViDtOwakjhO2xWJbYq3ARC5/OUE5h2Dc6htdE09xmQiXA0T3f+wWneaP
a0Rxbs5oi03cGmfVcyyk0XYI08zVwMQ40fa9RubzHdqE6Bcjwiv+9tV/sYY/TEM8FqiR1RvAXprg
oiD6PzABgVMsL9037R00P7RW49sCNQqhwNAmYkQ+0ucBkJpw01HyCi9CY04pz6sJHq0r62HY47tK
BxNeDIU+JP2WAPfeg2K7nTyP9SR6tdX6L7Pp6Xyvz/yUMfWUSO9oeF2mP1lYEMjVuu27ANgZQJr1
n4ytL6We3lu2MMWg7DMpRzTOlJLmM/2SBXzNQ+WWNU2YO1rxvKT8Dn+PUYb+BR9OtuKQMwSbrdsu
xvrVfwLT2QiNAuUI0vSzfh7rTWVDYay4u8kxM1XGaNw93SZ7zv85LoO8n1Morax0BFZXYpLKoPWp
6XfBABZ7/svKmD4e2J3IEeZX8ABLplH/OW/A70mQ2jhZwKYtq/LoQOxj21zp0gusVrDNtcVAkOrG
YOxpu5p22Y9+Q2QDExij+n5ZTD7q3wlmQkEdpqRPIIBeM/LjnShJBguzMjvyA0EZ9vmku0Nag0lY
DMMDa7U7yzP7oyw8zxBDEVyjIq6YzrtOnB9S0CKAYP1XANG1kOGDTYKHMjpD2/KGRKaSrFDCIv+w
kBJtkSoVqMdUTnJ2llcwX6YqpZddF26f4uS3pJDC01CgFVs+VH9Z9lBJHic2UvXRXm6zP2KrRdDr
Po97AKvjK8XNYsCVYVCkd0Z2ixvsLXd3/bF3pAz9/dOqQM4dlV8YSz0x5rRpw6+E830SHt4eWEZ8
9ba1obRbp2ThFOUM8kSCm4wTkS857aJfdIoSB0tLndiq/mpPG2AC/7t+EXcNmS3Pqv/OErGdpVMu
55Ri61FMDFRjHAzte1wf3nH2ZTpTWW4gD1PBEgeDffyOA5syT2P4GSPf2UAtD2xZpOjCSH70MQIi
U+Gu3+4XB/PEI/tYPOpdqGY8HMECqc/70lJNg5UED2BsqeHnVEs5dTP1ZYF6PnNN+p26DEvhjJxy
KZl2+7aHYjvFk1wUEy7OTp71wT2hf7/VzQbnryu/sfUeYxkRzI33FQgqZ4FGaUgt+MykUG+EnPDL
YXYwgKEX+QeS6mNb+qhdVNSm6dQ3VgrKsRGiys5nkTxAKRgPcstPxn4P8I1cK/oUiNPsnF+5SL6I
0ewEXtF54lumOaTSiTRn/NdlnPrHfkoTNH4frsQJf/nRA/qffxOtmV3XJMgfA9WOIkVP1+3D8mhO
B16iQdJHRpLHHcoAT28l5Tvf3QlpJ4BoTzOKHJgApmYXjFkgUnvbp4IEMeXykoKh71LkeYojn+pk
qvNfnT5nUUJ6PODeYncrT9znkVVVEFc9YDzpywUVsgz+klBSweUbOYMxbQeylz6ig+nohV5Gy/Ho
A6E4q2q+f2K0s2jLfN81kAtwCKgXVfiWSpKrTjej46SmBW8P/n5gGTVRmOB3Od45V79PpxoVX7G7
uO4Ocpa0znqjTwSXqNEVmwzFjcoJsc2NljqGv2D+NEZ9AwIto3yyz04DzR3Y3njji3FX2GxB71vp
SdBKH9dRMdgS4+3rB3BQRS/z3PUoUK3rZymSjaDhZ+YfFS37yv0fwnhM+YuZ2D/wr607DU8lGwet
Fa6dGtl7vdBAto2dDxgRWBnUm7VU6FfRiYIz5d+rwsGn2hAncLuON7gDrkleBjT87MKVQcI3oRWp
etqShXHPiQ2KQ6MiRF0SEqxHrVMW7XMQZuZJYFhceu7xEeXeei23/gdQMQRHc05MRvOsI8E1rt0y
4OYg0bOsVSQSJzHm5gGVCQvzpordJGb1XZG1TTAdk+KJTr8oPuQeemagi0zZgknpO+vBHxdD5bTX
3EFEN2KW1ciziFtuYFf08C9HmmzOb84SzVnXXDCRmijtqcm8BJndE5rIPgwJGjI/W3oq5S+UVq6r
dIfaWGTDFZN6PwrTW1uf1LsNvaxA9XgjYhNHciYFeZWJ2KrY2099MNYpbVY03ATeNdlSpsaEDh+E
4tCgIViJkxCH4ibquHhu3GOi6iIwiolmIlPf2S0Um3r2wMGcpihqldE/jQQoEscFGyCjariM4ZvE
kc5juGQW6ByjQimr7khvBgxruLlWW5siSeHn8nlARlZTbGFD9304ZXKxeFRyzijiiKQuKbRRN4aX
kCPvL1z2nl3CKCs3h+XNS1KIIWGkVMDbkCX9DNKCWhO7xRz/neKNRKS/PXSPA40frqIguCBFABDx
i/JEY2EVpMvT2SaD3NiwV4BDccFLnPQYGbhYFJ9r3KG8Iv2YmpF2Bss6Gg2h2v0cy5VL+KieXN7x
143CoDnVxFvV2IcruyFpPumG8I0eLau1GJgRd0igeSVITl6xtDM9K2VlKvL8wIKx7eOM+5cMElBE
yF1dgNE9iePGej7s1A1Z9DW+dHWjwDmOe+ilPDsFV8YTS1RgsURh44H5QGeoW1rOS0ioDBAMF0v7
fx067W5UinguCieqCwV0yOLK5EIl4ozkLnmJ4/CSqBVbLki9gQ6lAOxuf0jqEpyV10GUUH7i+DSE
7jkPekQ+UUUd6RIHwT8ZT89SrQexpGwU4wyeDoF9mxRFEGbJLGXn0HqSrxWTqGP7Rc0mhuH/YEdR
GMGSJiqp6J+Ah/U9vUuVAiA+q9Zo7bpEcnbsirwV5rypdPPHHRU0a91p2637NVovjkUFowP1knpp
p5qeXUbEjtOiGVY1S11vngpqHkTw58NjFeN0ByXXDCWyX3wz7FZm9HEvwZ8W4rnXKQLjQFDNkRpw
NvR+RCubfCtjNKpq9H8nWEQ6/5CKivv1i1SzKO3mzNf6piPCPipxUKJOxzvgcTo6JbEgWTzEsesb
S7wRwXdBDvr3/rWLmpa1NhNzzUDf7qU86RP4duQM9GS+KatA2xBGLFI/wZSVtLSDLWBYlUQtpWog
GTqeUlmUCz1eLNfqBwWmGCNaPcTPmxI4edQhZzRSCTPqfLGcePgLMiWHuQqUuJWB4N/x4UfVca7T
R4UoDArlctJgBHhsl5hnPJPqBRNmaYBpC7wwRPWam2vsd7dfVzMYNRuLECQsh5Ks+bi8MwigE5Gf
/Lhj9+hireTasX5Dh1y6ad8zC/bAxD+wuBre21VET5Gmcl1Kxn4cuexGat/DN5QfVeKOBOYukUch
9jo0l9RjlRJVWk4MG3SEMJs4UpCFfU54ddcdQhK0b5yZXONlDYtmfwhQORKEz3WsOdDAmoeq68KX
vXlgcuedWy1GT2BxoQn/GugaTx49dNVVLUN6+gDdO0KEPAJh7lHJQ1GLOOlG2j6gWVQWhqayvtXJ
SqRCAA4AAxO5wh3VqQP+mF2+PB0Ion3Hbb5rGz6Cy+qYfaZJH06XAfUcevhGWA6RBWtvU599K8WY
6rrriItWWfy39EYpp/yZUqKJX164P4CO+bsDWg4PeGZrzEREoR4TCfc1dC+WPmwbvja5A1xRS/r9
PriehSme+jIBwvi16whnS7y5LCTysNpyHZzDHzHRGbuzd8RyE2fZdbNibGs9q2ONObqxlQLOVcmg
7kKaiY6qRFtZZkWnDodrC8Mgv0rZbcKOFybGKxfF1mb26llaqPcYmmNg+yy1jZukNrXoSNVRDroc
d3QTy0g4MrbxMOI/30xEt++q7GSQayvXpXdld2iHTWY0MlRvr1kJGw8FFOb6v3xe/I1i9+MLWRmA
M45t285yJ0ISBImmLfDbsL72VtDjcr75BlpO8OplF5Ij5iGQKPnAVXDb+7/PHL0Nns9fKDaro9wr
yxQTqdLMpRL1Osp46DsAvjBhCzIuFPBO1J+M0ZMp+hXQrPkyxdO27v1WHlXRO1Y5Sg42svNX0VPo
S0r1dRy+izI3XR+eIleW+Hh6uOrvck6LR41BM2n/jjUP88J/uytUkGvud6DLdH/lm7YCcRX0/OZR
nTbcj6giK3BktTstVYXqqf+aJ1wmuGZ2XT/lErCNu+X8kHNEIzW+OfpqkPdCDRQ950EY8Zcq8JvY
IXEQXbA/d7c4ip/lGP7AEGWvHJQ8F+KwEjlCPqylW8HCX+NCt4AnKq5nMMv+Yj0cY2o96tFRX9hv
xWxkP5wEYLrqC0B52zGh/zwMsxhrbJmLCXeuB65hvQPiTTYrAQHm7IxIohDm+0f21yOZ2UFb8PkX
wa2J9BD3Li8aBXCUiyHaRDLZmYJEwCcBm7ORHvvNMvzkSuLVckwe+RufrZVgbqL8TVnf1V9t0nRl
bJ0P0vWSMpkYyKq2fmqND91rkAyDjLeN65N+APMzCD1Wp3GpEKiv7rRFl3sd+9EKeKjFPbgINDU5
U8jn8aDIV/I0fOHHIXkT1UPeQb5jZhwpCJkbYLF98jXeLszAahXeK10VVg46SKO3nNvA9/PdoQRD
ydzyKpTrq2RwVRfwUDHaoMusIIdCbP8VafYl/aFqlh32c30jvRB0tpGiY8ACPWXi6fuhVOmSgVUH
6QPfuSFXLhjE5d0TkKmXp2OXDLA8vxQTVS12QmXjKQrUDVcSmOryttG//iWLZUXSaBzfeK1GdWKh
E09hC7zpIxh9YzB4wAlV1CNzkaD8ZeOwQPIOTRdsAKA0yEm6o4qjKPOXaOqVVrCKGTBxLuV9dch5
DvAufWoAKYXC9N4jtGOHQ3EnxQPQG5ZefvYWJHfGjvZgPQ4kAkCA8Hw0wdWWq6hi5RA6epNl82EO
gUP5OPNkm1YyDml1b0YdFYnPGAx/mUGMLSWyfRt0/KV2/ih6Cu9oRrSzq+jd0MPBxYfj9bGp8sx+
6g+KtLzTBHBXCIR/E1WNCBwArWSuPE2BL6yBWzTjsyQLFAyCY1NjE+niyexu4UdcBRkX0KDiyubC
GG/9QKj5kjnyunZ0TGTOgDWRRTO+GOF59dGrG4QSVlGxpj/1GAdXag6/7OWYytfqHuZksUYKpeXL
m2q63FY9khIOiXwmucARHrABjuhsA7pJVMYD0jRC0jB44OP5Cb5kbIV/AKiotLDmK8CFg+iG2BU4
WEHqgRD9pxUXw64oxnSa6mQciV525vyDj3+BRxpXOb+hJYk7d6W66l9t/9ApkvQso+gZKeKo3lcC
1B0M+I7nZh7l30IRC091yPgrLiNl0OyhMM6G2TrVd9sGfxPdCtcikbrOF7/f7q2qnA4xWSStNuxj
VUhALU+0Ps6tj90tpWv3ilk5oJUHD8yx5Dla/4oTjch3oDgutjL55Ha2SCNqFdPcXil36MttrjK9
adQhH6Ob7mgXpQANQigr7hu/lGgBfG7Fr0byLAgJh2tnD+ACMIqjJT0wTYGa51axK2/pYt8GoSw5
1D4CBKhH8jiME2hOYRYzJX5jtOsTP9Fsa7RGn1QU9ywnZMNoq8pufUONzQ5EaIiu9mQ/8dSKtfln
RuYXOr5kgYe9WyjWcbm3+aSwyrtnC7Qe3RR3DX3OlOOjZMra6RiEiUg6j65IINPz228W44dDBLeL
TsItLVZcxWacVP45qB7qyYSBqxIqDekEfzqbCbOiB857OU0jZMh7f3kRNt3Z2LQ8BHofC71UQ3uo
/2dqZ2TsEblZEbzrdQJFUlJfW6UBETIeP6lyGhKVvR3cC+9Qo872QzAjQ2m11YLIyuXaQ13Y1GZT
jeUNESWKw30Fretat1rr0nn0XSC8ORYR5Jv4VUWsMdk+w25AqdgCpBzgNdlDWcd/L0d0z8j1ApNx
0dSXzcPOUNc+56siTsfJAGcPnRF1S/1m/lOnpd+buskqPUtwA92Js+yM3w/c6nG2Z2oJYmtsaNI1
kaWIJmF7/XmwdqWlj1hDjkPQpGkGl++oYfWZMLQPgbHCgK0vdHGaQgi6IjdAhoaahhVHNpG9bzah
ftZ0zsv6Hc4m6UbQeq3QC+PKcPkZv36v5BvgKhyG2vo1Lx8BmX1e8sM+KSOYFlnKTf7nPkqf2tZN
ZmfJcWZsDFF70/KXCtXRiEFUfYbJx6IGGtOzL5Ssvk8GGtG7W9GocSFTdZgCiXS5X+Ub+m9Aht+2
ClzxG2eQvo4xOwMrIDo5wpwQq6eZg+ktMrNa0eNAuBQTZOykCdGRxjA3p0EOpi6jB56gkGJNynHI
RiFSgPxVE2ZbysRM1q+TK8gouNOHduCSW7PAlEBRaEoisA3g5Dx5y3P82XX1APev5A1BBFyjaKCi
mXkFvfnB3tNWlXsqUaXywIUu7YH9kj9cRSTyP6K9kHljA+yQaoA7ojfBmDliIeHyQvp81x7Fnxvz
B02CU+80/Mt5Bw4uofm8AaW/4RNIVk501Nzy242D5Fu6ysDHHF0gbQ3r32wRUkI3CEmuyP3/4DMn
lye/AyHTPktD/U1pCQymMVeONApsQ7iAMPITtwYStfoi5OHaXbWbPV98O4jplf7RoB4fmZVbk1Ge
mEgNUALXgcd7z2rCo2/UvNWX10/qaYu8HFj0dof82f0seen3j28T8OiCDmDVNbqr3eQZOQSawr8w
tNS7o29j3acSoG8tO07XMHgCSza3fwiMyz1s91e2nGjlI3KRgYutCb4w+ONa2anlv/VETmP0KBBU
X17DAV2nKJs1rEBqRk3smynipDNFXXVxAw4HSVlR2Q862tGTjJ18IEX4pCq9iQoOHSGl35BlMZT+
KEIBVGQz5/DgU+P0GcljeVnzR4k00bF4dXwpQeu3v25vOgOcue8ytZ45puzEEZYS/zTO/e/tDlLa
EU5K22o911bjosfO0xejSL+3oG5oguj3TDPcuif8tpwD7xOZ2OePTVy/sWmwsoHnZLqywcgSfOsu
Z7A6Fx3DVp7QZm/wsZklIfcMrE2S7IxgA1lFMII4/rGUhjOOFmemDIX/hEnUvm+ajqNRWzzeDqc7
MREMSg6DEo22vrV8FBxvEkpV8j93cT6mzDiS/tNpXjS2rTHCnHf19Nt+aKJfmvn8VjRRh2ciOHKS
jUfuvfWmQnPu/6CZFmht5JP35vEdVzOrRNEB4DuR4RgK3auxSYrwtAznfYYMIadqmL2nZebV51xU
QVFNqDQ0XYUZ19AH02ut/Cf4ZEWfv02oElsPyqR8N7FrLBC63ujOfY2vCz5GWjVNfIkq5oxyzGxn
dJnK9v8ndnNjmVgQ1HYpSGAXjIz+ywT+CU24x/PgtbzF1N5NXtmlPSPY7BSWlARQ0rf7eWrb5xIK
lEraH5U+9uwxx3hXvDBbkSaUpm+BvEF5TvLVTjH9UgcKieDjuFc3pH2PCfoe5IX/RY8C9eVKpjP4
Agfm+k6jFZq3727e8rffB80AK9QmFbiEsy61S5y/dLV7B+FLdTh/QkvBFoqI77szj4RryHUGLYUD
7yrLhRbNVScx4DSMdG0BVh+B6Syu7RgDQYG6obSRjFcKh14q9Bl8j5MKH2IE3bAC5ew5BG1t1zgx
n5vqr4fhRqI2bMNyRQ23c45zd//QMZZOfqqm5AMhR6/kS4cui8O73vp5muHsi11zQRblBthhKUMV
CZZiEkWQSUU2/mhP5zGj+ZBrILcaqQ9ihvlQnWspCPGPD7hkVPmwPml4X+rwclqnVc+g26KWk/vP
SkcO8q7VZRTJhACgVFtX4j3SCC8fDBH7pyzQE+gB7XMe84H5756+syYvxFMw+YV5T1PFXVjyPdvb
J0afeHKAzL+F0GIWVOG5d36XFj1X+LHRHb/Rl0iMHrxD5VWt7SHByB26VDkTmcC3WbOj6A2H+ZU3
dBB0IWn7TZeIMsBe7idYIcrYfjS78qmB9OqSf0tBr+x3293tCN7dLuvUoE+RJvaATs5FsLCEgcgJ
8KSQflLCISjybD1ogMzHUvZm9vF9Rl3wMZdDKQxPG91h32l6aql8NTeZIh0eeWiZmFxU76dlmm3G
m5+7NU2ikDcGR/JbGje8qGhsSvWLGGNAxWqLTKLuzpWdw7rYuwR+9LxCF/Dg2iaDlggWYK1qXqjx
X0pR4lKDP60UvooRQ81ASQKgM36HxDIjZxgEJEWB+Go0v5MPCbtsc7QuR+lIFJRthbLRSFv5bBFr
yP9Ih3ty4qFfZDYcoP5xCTH1TOISPTxkyftxtmjfmpX/x1D8iSBaVx2JxvZTJFXsNXYexoS0kiD7
w4o63uaOLzD+TbD5t0ZsNkRxGTFt5N+88Am7FOyzPbDJAqXLncrxADl6YPI1pQX+ibhOYq/EsyVi
+o5v2BQgr1ZMchhtkIGL7s8ADjYB4xv7dD607IdZ+aD0sMDFRQZ44nC+jrhbivRf8cLGbKcgdJgW
kkda5XR8oawtkaJ52oYr6SvJbiBW+9worMAy1jbxxvzF2iRH1eA3YHDmd7FNqaxkRWvAp4ToDtG2
rg6S9wT0dCzvK7sHiND5jH//lhF4lzHU+zvV0pxqHPhco9kEt7AEcSRscTbjmdeRgFL5OtQy+zmC
ME6nF7hh9ZJbZE/5amH2I+d0TzFMSbXTdTsm2Uu9VJDz9ETd6zsBBpe9JwBSAijXM+7nbPts3clb
Q8BdC72tOg/PfgX1dMcfcIVaGxAtByxbtVwNKV8lBuZzUkqk1DX3KQKZ+FLR01cmRBKIQpRmRgyD
j+gd5ij1EmQaQJlnxNWC+sCSABhBgIcbnqDQiKpvvLPCMxAAEy8xeLi5osPJeTWNGbsp3E3UmwWC
GYLn8U3S+PDiOltB3dYBXBvHQg8gNoPQjcmlkFcN65v0FMV+SG0We77ijp4N2tiDErWwwObbkL8K
9XIdeeLTfWkKGRfIItDzKod33PNsaoic/Htm//ELSnwdMVWywEoYurt20iwBXR6NilhgVq6Wn8U9
EHtm/GYv6M+amfC+n96FH5biB6ViQ798k1PPMXVFSxJhqTQxtLcXkub7jnHk4QU4ElumE5ZfFnKJ
a2vs7SBah4K5a+VvLHJhIFCA1t2Ve4RaKmjLsQZr4SIJHBTvYjmd9qr4cLGERrtBtDHZLex3l1D+
yC1vuJu8G2UmFgr8mCyw5ks2W2CB/WyYE/7UBrhHiFSp5J5nsx1y+pkyett/vIypOowIErGayOzu
Otrd0NyjAXIbWueWN9Jx6CJAS4V4Qj93vpICoCJyk/O1wfFoyzr4aYpRD2RQHYF6Z3MwxbW2F5BQ
cQkiQxPRHJqr87RlhA0fq3PwbFr0RPPSncndAeYmRPDAWnQnE5UFGVrY/oArNBUONMJOJZUMCXL1
5PW3xOya8IvrHnQhRrS/9yWqCHMJ7Pk2sEY/7FxAf7xjuKjl2QFTXwf0DFA38QwDjoHdCwQqoGLw
TqfSLwNUkXiewrBkiqaRAQIT2pELQnzcM3oy3BopwNHQkOFDb9jxa6Xuty0ak25MzUR0Y1qvBagr
iYz1AaGr2JUqxFWX9NCfF17MnDPtsufTPBq09jys4gvhHqczidurAjQP+9oVT2M/22nWOevmEPbG
heQ0vdCdy/mfzjLT+Jj54RYZ917OAuYLGjXTnetdhu3txp769VF23jVUwidOOG5VYuCeei+uWWMN
gjRSyi7SIMOu2sOG5D+0jEopXDD0slDmgRPvqx/otM3/MzjKzFwMU+cKg4ty/hE7/ulR9v+QKGoW
afArXU9uZKrK/ITxUxTRrOdOUd6XE1opxWZLurxQ5mEHO7cQ3m5OFO+X7yWuQVJyXoY3FR85hZnG
XLz35iUzX4kTocR2AsFruBtnIbqwOago7WrZyCsZmolTY6SQca6tRfwwgp4qLwF7n71WYbPO4VVu
cyr00cCsXb1ktDVdOfS15Y+La/R7yJxOhWpi7h1RtNXeqQONNvZ2Xdbxd+mSyZCitTVtIchw5TJo
CSJLxpaZzLHzqYsBQmK5rAmQ+a5Rm7yEB5UGDL8mWwzlGhioUJ3EQ8QWjyPo03hyT2ZmW2NFdH54
XzAA09kyvpKQ4Nv5CYMTQEVofv5l2VjR9u2MRzVm0UjBafVSjBSHxm8zP1t1DcUYzjrdAhWkAkm1
cCNyScOgir1j8Ffw2c9grNNFR6utayz87mYaNOnHq+G/TNeaEUbbrLzbExnqwQOmGbBPVdxZ95r4
Un41yj8ye02HA3ZGqwVkBy4cjR1wcjhGKbYB5mq065e+tv0KbHRyTxAodek4zrXYnD4NnGtsFE7Y
IjWrCpA9O8Fo6kwcmLIcGDYoSV/Akat9MEiGmE/l1y58RxynOxpsDQcamszoxQCvnKtfxAJwhLfg
ZC5e99oFDFlE8yfmoIOaS7MxeRi2qUdjh6yU+oZzlV1WAIxzN1n+gcmNLofaFAmbQJb3sblx3md5
GA+KE0p3alc+VYs6B2c4ezf9hal+pF8B+3zSgs65gQWhPDMD+FhO9SvVin7PRcmDVCqlgj83FbUM
am8/vxGe9EfpVFwvyBBebb3ztPmJGZf6au/8JsVyq/VYc/YmYiE3560xbEL+D+ERq54YbILXbdm+
jdkCLUMcb5If1DAWJ/FtaLseQyMUwIC9yn+F0YBdcuevslTkwO4GhU0gAAoZalattyo3696GOPY+
AW2MDoLl6rQN02CP5BBrEiI5msjqgC5hzEaRO0YZgKMOEITk9/z8MuQtjxWD+K/C3Vrqyc7B58RD
r6XaLsnUjk460FcPUzGsznn/WUNHh4WJHasf4H33b+sawYbGc3p7TJO2aopJhP4xMgxHPsY5Z3Ez
7r7y7+MXdh7Fl7JJThilemKrWlnwJ3gvGFVKG9FXyHaAq0sO/3Ug6s/OkkdVTdMm5sAMLoF5854y
aTfR8HyN8RODP23ZwyZcWum4Z88verKWLUOBtWxzvMq7RFhDF86b2Mx/TRD1xcy3BhNxmOLts2gX
K4gMhlIZlRgucyW9HgqaaxJ34CY4KUfRPuHityQd8tW4I+V3RhJPnRzAZtBGKO+xuldoaD0Bd4kc
3+dslWcFDuplyLjLX7dSnS9ig3aKD+Hrw/44IUFnzQqql8yFRK+lth6l9GkJCwMR6Ma2uPTq2HPg
m/4sU4kth/3q15eVurWEoW27852HnRk3gy0UJ5In61f5P8TEJV64HjV+BYOreR8G73ZQHuOQnnZG
e+Uc01iFZMjpSmx5JAqVBSl1MsaDWJ87EC+qUU9/LSwMye8g/96UxKdkoXRYyje8FLXoMrGvtNuG
a+K3EYrAiTRP+1cOWR62jnjMPbLwefWkX+JSjDRodR6mQlkINUAurOowSEAaHaD95/nHfBW/asgi
H1xQfn2oVC5vOZeWBKlrz2TE5bI1O5nRIduD06VJJSxLZBBlduUkA0/ILJ/WB8krMKNq6ZMpB6Nn
cB7/hQWr4qWRPJ/HcJHOc+FqZkgvqBlfXBdyV0+CEzzILyfr8n8VfFVSITR8UOIZ9TK3qEKrKknZ
4nTcnl22TMEJjOlb2J5j/T+2yTAYQ2bmnYJCX/OG3Izcts8jL4RT3xGgFXwXrRRCJ/4Vtsz556J0
XaOF13MChEufzXHiuBAi+bYUZIEa04Ezoto58Xvdn6jfj0+MDVvjTobdJXy9oR/4G1ag3iu3uvHN
HC0xaAP0Mm2ZQtnbKYumG6vOyN9VTzzrgQbd/axSoR5TORGzPsBNtNl6TVtnhdNYr9towULzaTff
xhkR52b9FiXzPon7idV1/8bGViNYPAOBK3Sh3up9zvG65qZD6hZVaEW0vnNEkvDXRj7Eozw8LdEb
jz/oAMjTFYdV8VTOV/XfVvGPrs5sQ/FQC5CY2GD7OzVCCppEnUlpmhhjXdREHC4qKun8a2emkOGl
Bs322WY7SH+4onPNN2BCNc/sTgkObfQ+sNNLuGG7Ay/KrVnjRCzXgSQNahTUXBOYWjckptye+YhL
s7F5Kli+qeaWis7f3Uyy97jEYhZh66AFV5k9CQFHmgQgtIE0LBcNHwe6AYAIVDqy2lrMnNNWfNLo
Y19lIC7WV1qh4nWXUze/G7l2fzuT48MfHzdbYh5LGL4DRhYLuuIQHKwjcfmO196xYon7HgmTKvVD
JuCBwdCTWuRUcTTItvz3SfmSg225BeI7sXu3UrBtv3c5oP8lQilo0VJ1mLttwTZq9xUCmpUjTP2b
zxZMqytQDPZHrpdb/GlSE/u5yytICjIqIDWwOL6Rg5Y0UrQnKWqFAaiaNADJU8526b9HgcZfX6PQ
aXwv5qlKpxwzAeug/ehFEq1hihPtVkrM9RHuwVFEQY9h2VOZ58l2A398AbK+4cuiDFwaHuXp/OYk
d6wNWqVmh3E8iDO6/qP4gDc1WkIvj2ZQ8mQ+hTpUwBih1HYO81Hy8a/WA5YJMFZpbmECVIqhLFtr
sAJ0JVmpIwNaTHQ9oyxd1AMd46LBZZF0QSlsFKITl7TdWR+sAWxyarHIlww54lx4ChsA2uaELupS
Z98+32g3aIMMwPmT3VlVmAznPN2aOeTZNribzrOqQPgOtE6iqzWQOtYl7a1r+Rxno85l7pDtftkT
T6TdyXnhnZs5neGF+GzviZBiRWBiktaBBxYdmiB/vkqIJQXCzGO7lfPR0LaBUkzAJM/U1FhzKlv4
gmlLS3WCAnXCWXhVtla1KZkTVgEfSnLiL/voKwm3AP03kl64MqXCTme2ey3ozuatVyZl596fy8Sq
xePzZdeszTGFIOnSeHnLxBDdn4ygFncWbLnoSjHgJUSnvOaPAPLqj3BN1qrsxhRYC5yOWPfvj+ps
sb7/lgZeFtzam2OyJ3spHMa8M+gsS+OcejlSZJfbSLJNh97o0a9z8ryLjsA/f7sLS2r9yzO4Ge8K
d1Uv6ax/l9NDTYRblyKYsUYPSyCTptAutDjMtKA1jY7duRYS6HVT/1IYR8jTEVX7xu6un/YeXI4Q
VJct/u4BKChex55WHVN/nrliWa0X7qwQsguP6NacsHHFLR1VRj/0Fb61ibMXAf57weaDyXD0ZcWb
doxCf9neirGaHbIA1jUbGQD1Tq62U8fxuK3nAyFNQ0E7SPgDKPMWa2GlF1i3Xbx0qWNIbffnPwxv
HR4mViNSoR14aCQ4RpKzRq4e5aKslA6VTpe1e7krqjKWBZvXulyylrDj5Y07lXLhV388YvOGBsbU
Ip1Qbh3USq9yTQvQrY0J7bZ9kNQDAJ9AAHqBAxNHYnz+OJ6BloMtVvm/9WGZ6/3B8oujS6v1Q8Wb
qms1sRg7G+apDdCPe4i4lFGpozEZSxaVc1b9siXuWP3W4BRrSnS0oyUaFZM9wuU5VeyzcU7Z9D7i
5G147ypSm8qJ1C6+bYj7HJbzfkH5zfj3PKsllP+WJ0llMnNMsC6ybtyhyYXOrHap81zHvA5pCHHk
kQAXyob7/rDtMLGEEX65eWQGuDs8d1NvxnYvVs29kQ7QdY3GpLYwauI4YbapP1lJZ4X3DjyLUksr
wS8bwr95YVF1OLzVl2yUk+LNnA/+mkC8irZOjF4HYhgSkSW5ekXEjIPrRXzFbTYMLDb2JhNmJscq
fAY4zgW+bACTeQRY1GnNrRq1kT4dULSXfCfZF1sSoQYnQDWmhLOiva3VMryn3ZWV1F6IZfF6KE7Q
yqbMqpl4t5YFYY6qCNlJ/VmKdp2DZSCBfvByWIuvbvaluwT2M9Q/mnymVknUFY+qbd/vTFbkanzc
fNtmRxAPwgT+wxVQiqCmkQopJqq1v0/uVFF12vtlUVVDElftABjR6hZqNddBd4SAXRV43NKDRr8w
stS7BqQbUN4CVE/AWLagJIqXLRxQbJIaFSYEG5ybxDQ91oSXfqp5VlcduqFOHhy9nx8FAdJ4Bj8m
M2A90wJ/oYXBRLm3wzpgKR7BDKVagO0AaCeMswt5GboG46aSyrvDnoBawWVsL9avajDdn1ZjRkev
3FG+ztP1hKfMH57TJ/qbW3EEr/T3P9b5u+d3YcSaNy6CwcPMXWpVrwAeXBQfB/8NA4Wg3jAkqMUD
HlL2PIsbaG4oXuTG7XKGTN1LKM2MpHjBrt3CXbiXGkEZXyCzaq9w1gHcHsXNoWBfzsVQva7WjJCa
qwDOgHmCyK+Or0QxMtRl0Btdj3MNJFwIPCgMHRjGjvUekhyg6gS7JUxundR4EUP0h6K7j/t9qa1G
qxv5VErdtYfU/j/jLkUse36WRXpA8nKkfROMz+JA4SFGcHnwGEutJATKS5Or+vl6DFqY8tNNyuOj
ZbeOCb+zHR7BQ5FE6EpISrhSGTFr83Ld4UVJVV2J+JUuYa0fYwm2LA7UEooRcctBbiMvEwwyw01I
CkCWMOZMuhAre7qo3M/r0k7g8sym9fI/uCx6wAZI8MKzNWWDR+o70NuQ0OZrgoiStrywszsPgBuy
P0vGx5WU9R2ee2AM7D/z14/1D+bo+6b/Z6Jp0Ih/h4/emRLZmzek/4mWUDCPnsmxM8iyGr3PZsx/
5I0zj/UG+fEPLCVXtGTEZVmUtU2kjA3OpSdKkTRuWak+dLXJXHhvxeduC2iluaKwWM/py1JTN5at
pMWyxpu+8wmWQ8Zr5tgt9qq1QBpEq14QMJJNDc+U35sBvKauqT7VQ+bfOZdUzEprNmo/tHoVWkpz
YAp0e5+4RA4E4Ax1HNC0pZpnln7iYep3haUyfm7NrAe0fskJGqMpUOn1++Kgref/FmFRI6k9lBwM
zfhk9KMdzcZQ5eEUqvqzPhO0lw3V5ZmfA1UvlYc4mA99cauP4So2COi/dFA5feNC+3zH/ENX2V7B
dM0uHMjnIBkc3Ui4M5+2AbdWOagNRSwOg+OVm1IIoTCPhnTSdtsFz2xTaO/rw13B0oBHSAI7UP43
qmYLaGSRalgGEO7tt8fWuAopkhJJM51i58qHzRO3lv1ioYyOtOxqE3AhYxOmezqZ8dLlNLh1/Aex
22eFJxOsZ4vNIzq645k2EZAm++qF/wTaoEsogbHZS+NyC1A28ogwxS3iH6KFMOTajuI9V3dTPxeY
wddqs8kjvUDLnGD5gJ25VGzHrwqZfw6ztKIpIEad23WXSbIpiOqzpnmcbnRHptfovxmMlgSqMztb
OzwPYDexMjFlvLnzfbl1MbHPA2tmKBJe6V1IKuEF4092MPcNMKHpemtmm9PFN/o3pklMrEyDPMSe
QhMKG2A0LDDyEauLskcW+QEyFgZIqkiDdzeQV63FT33sLrWjulX37qi2UEDvFImQDhUO9v2gsn69
ShFqCDDr7zzdEcNrV6Hx+FcuI7h+ytLwesNwP4RaCEuAIN2o9Ej8lVtZkrbJ0Mbhcp+YAJR5v2Kp
fGGolua2wgGiLdK3ZB+Czz8d4M1ak5x/z2E4/8OFb8ykv2USTprJWTQdAH5NYcfiYUylqsiAKn/d
xtdwGXLW1k3+IrcYfriUspXdhJX/JfxIrEbBpxFOtRfsZ4f4JblQqEdbZAoraWk7wzeEFTcXxCdu
B2n91mriy3UHsvMorwt9oJO3EBLxtc9IsXytFqmJbL/tYCh7+1aR6vaetJ4hkF84jaluEWVYi4jp
RRH7HyNLfbFjWniq3qwVpCZqtPgSgal0et2OOMlJkePooDp+yIfAQk0lnEvw+JDOsFZH5qyBt1UN
DJaGOBwq0Z13aZ35mOxJadqw46KoCqxuJj244n5WPn47KSzQvwbzym0iSuuMP9aKDee4wp/vNME6
foGf3DhtZApP8J5aBVOw4BdFwahwEfku+ilhLnllyjir2oWji75iveJY/I+RqI4WgzOIiX2aPi69
tE8m5R7Oqy7ptitnuEwKPAQjqat67eEMKhznK4fiNAi9R53RkLv94x0RCmYlqILuwU+bTw7kp0I1
lo6mNse+oa4sr8YywMg9FzJqC52eKNRi5sV5V02q0ce6ItuTQiG6C6xkFA9zz33aRtn00es2Q6bj
d/paHT2KVz2ZrZO7zRVTaIfLFy3wiWuiLQvPfnlibYWlG/50E2cYGeLO+pl2bFqOr+wWTg5x2c6a
e4aheVi//vP1/I35ZWdgmukfubdohGiQU2Y7s482IWky23g+yQG5vCNHYXHoi9fYDFwz63mSCrfK
rtf/VLaT40UOkmV8iAJb+MoLNs0OoPJFG3ue9BcaqZapCV+xq+01wIWltqInYrI+tDBP9jYmeUq2
IBX2KKu545hC8CfD34wiyUjnEx6uClT8otL1tfiuzYRyzBYFExk9CALoe2s54W4yhdmUfwNyNzVv
dArwOJX56msVzk10nHworh0WIR4H5fXkCCA5R2avdOpB30CuuxElE2kpXfjtgx46hO5iZs5qhiBa
hq4EthVExwSxYpcTedJGbLEL4JEjEodozJSoH6yuR04d5v3rAYd505mSNOE+J2BUgKrr7CINa6Ig
JhGWawdIVZpks50Lukk9W4z6ARykT/2P9/tc4IZJE3Su+X5qfTxTOW6x6XLCHmnzZF0VKLXjYgLh
0NTKqB/MHPhDLyHy/V0LNwEZg5aBNf5wQlI2OYyghsPySyqN0dkPssZJq5Q8e4wo0zcuK5a4SotE
+bfDxclquXmMoX0wn/ude0pIf3ZR+IIdyJ+jxtb4Mm0IDqrUDKrxLyEX0Be5Yu7FU/T41IR3joqA
Op5/SW2KjqNDrvAdS0VVTbkv0U8tqXZmRFV39Mcpcxn1BMzOL0uvP7tWJfVW+c6wifEwXDQRRQch
iNN7igsTZ8D5f/EwGW+++8a6pglz16q6v+O2OgLkClpZimCwoqm3B+pRpmLAS+EEHee/qqg1U2h2
m6RTCJt3XTNXyRWLNbN5CdYH3QxWijplC7SS5E+JEPe1D5I24QFIxaUJHWbRggnCq+UvL9Qo2yAx
ZT9iTVHyQU4DNxdsi60vRF2ytbSKJ5cLW1XeBG7WNViOzfIq/Fena8PLDecAI6LdH1GzNVbED/31
OF1GOoFjGMOygJGzxSXyXoSwI4dE5YGVnALXafxOud+SdZKrv190bZ8Va8HgKbN2mE8dyeSq/NFF
ZcqKnSIK5q1lfBwr8ZZ8IPQTUtu3+8QSGQ7gdA4R12FrvNbaKOOB7XqvuvmfveUBUAKdOawmTHAG
BEWUUvuxx2rXydq3vIVYkGctMx6KMw8udEMOjcG6gC9ABnE85/9x4uNnB2eg025buB46OQHLTNkI
vguZk39OHCoCpYd34YMSZhItPSMpZ54xSf7ujmLWlYa6RIICWMDg8drrOIqwqLt44OoOK9RunplH
i37urMkTqBbH4mwLXviJ7UyZtApE32u9f1usL1EzVmOgtEemxQPb1ZS8n1KOTig84230THQbPZiF
Wn7KGu1+CkGZD1tHqHcgEdY4RKyExzmSZivQXfBrUSClgDouSgJM+sgl59xQSLo1+NgJ57aTKzVv
Dg1I/yBa/ap3TBr+FMqSWSFOEdLKihOS0Tj7j50rsj1wqL/HtdW5lTFhDCf6yRo/ewgIYgGs8vmo
8gCJYPM4C0lwXdQ6BjoY1EBydJgpOTGueByQS6oZQmZjGScpwNxPySQCDS2PgTPn3vhBoiqHL8Lq
qyXgAyz0UawVz6mIMJMOnJb99oIh6ntH1mJlMlVa6I2GvQ4UlOTHU8K4XT3I5nXtu66Hqg0lnOj7
Ee+Fx1h0nmuMp/iU9rP1upCpOgCHb/W31jmxGV9udwnRKyeoQlMKp9+K3lGn8ox9d1jSZ3NWa0Vg
n4NnSB4CbuQCxFpfj2ApJGHasKdCEjW+TX+EtPzTiwjYNZCPgJRCyqEIG5HGRLhDh3gPmNZuQQXu
VtzmuipSg5drO3YIXyfhX9MhtAJdMOL1GnANr/TFPfHSHSacV97pBxO8wqItSrz3a6JCla1BGGS6
zvc9W8xnKmE7INmVjbAjJM4RvgZN6F3hITnf4OnxsKirHN3flfNy1mHxl8XEWm4NhZSLBxPqyQB8
ZGPvpblu55zJ/EX1JG49in1wunN3vap7RB9J9m6LuC9zy/W0f2FGVbuoRKZqyTWozgAjrZFaLTS7
WOcjYm+R9M72Q6Q2XwLiRZJR50s48IeG/dkvKjIym4SoFfUdq+QqYWownb+PeIzpKD8OXdC0oaQy
TI7FZtG7OSRaFGvNWEdo2El0u+jni7kedJQDuYNySbHkV04maN7F6Qi1Y9Y1wXWmi8qnmwS0TgNB
Ce8z5l5FwIcF8OJ/NoUJvAsilsMpln0IExLNTBd1DfUqEBomrsp8c2ANEJUTi5RASGEWGU5L1KF9
7M9U10OSlFdvOOzJeVnED9XU6ZMJ+i8caq6gS+eqLjyPz5EkgqP/3X9FPKeIypZxNbwlKyLSwHy+
BLqA/8ZB6tjLhWdXvL2W27vY55Kx2LQptiiVwZFoslpRgUoGLtN5GmI6T7FIHkw5v7LxWrJSk0C/
qnmcG+mzu/Op1xMQFwzdWvjdznzoRSPsvTrHMmtIqKvf8a7c2GGkb3oH721zuAxTC6rdwG8BLImo
maem43kPeD+oV76RfeM/17sK3NZ9EZ5IYNvNrIfRpWFAMsIq1TQ+2eJHeggVROBXXFSW5wYdZxFA
VK2Afyse2+hlj9DnrwwTlxsglPudeA2DqG8EnZbhhtH44sWhNmAYegVaKa6h5QcL7XnSdIyw/eix
Ed8jWXqN8Dkeqy0uskrcAGgewBkUPzMIolVXbawkaSKzJGGpq7QzJBVV8QZruaJa1xGAL7RABpdo
v4WTJ2vUh5R+kW9vbk1qVW2DKdwipuIO43kUawFjr+P9jKyyZq+LTCjaLNUW96qTd8XdPukoAVF+
sHUBgcWCU2MBsEV9GvXGrMb6TAR+8bQKyQuMXHDxp5nKhp2AH2L6GrRNHhvLEVtk7TEuM6RLb23v
hmRlBj4BfDYWDqUzWIJW+ZCvBmLIab51bp/B86mxtOZwQ/wSuKJKYsUHqb5wci9b2Y4CvKQXw9Wc
SURrajHPgjpbRDAI9igkEEkuIe/+VsLHDlMOePGpe1noRUoACStViEmef56qQn9mn3bWNzqn093i
Tiko5GxFrSBPiEoeLBa+RSQ5+ydGFNuOTy0wNGli/qchj+JP6v/RrH4WulaMk5VlENjTMxoubIij
KP2zMr04orG19IHt8+QqAvbxnwONX1kWyoEySvS3fRT7PVsUrE9E5+AI0a9pcfWDRnF1vX+VH4wY
kXhDblhIaPXM2iYNCu9nEgYnYkePWsDfpff9bdkse2xL+esWX/DMHzsnV42e0HAEJ4pI+Mx9qvU7
aIWcbIwj7fl1Zr1Xz9ABeszNQGb/+76GXU5LmoeUP12a4+Br9eY4upk5/sAdOTPqllYzfSkFni4Y
mWyXrdPboU3w3IJRR+nFVvHQdNNP2g0R/8J9LX330JTpH/oNpKsxM4BzCpqbXUZX1PGIMYoYVPL4
4qqhMGnjN0FrA9z475ZWTxi88Wn6ascbmiS2tozipuqDXUUrbEkmv1V3nDlW0SeiSkO7l5ZkP3VD
R5WnYJ4tG/M3UabZk7w2inLtLjFebOFQvuXMHfy7FLNCmrPMTypfhoBoXyntADtqmhhX4SBFWpBo
fyECzNRYmR3y6DNHT77O2FWjKQJeNXBq6qDVaa/nHeCK68B3kzVvTCBQNtF02m/i1/uIpODMZVyu
8BbpGBtVLk+txBG3RmKiT839hz7um4+CIgjjEZ+u5eKoRAlwXFeQdHrhtnOy2vsqBks+Eoqg+Pc1
zJPZjB5X1WB0GsEWox0MzEvL0sRs3NyGlFvs7NJYETfW/yJPAVryA4AyjXCVEfSKRdf2LCqiESYb
fNhwnWIFC0iIxF8wk2JS1Paeryzvm4+mgEjXwJy+oIa+91Jng386NvBON+dII4Pwp2usxrnyKEUC
nU41beWMpp6uAHp7JBSdkbm6dUhsRSdrIFkPDrxI28FQaOLFS8rbIpZdNI/pFC4YlucBQke7f4qw
3EsysB14r4ZR/Bp++Cf0WprBOYB0QWN9gvpZ5hSq8kQhTGKFV2jUJjZONrE+7pUH3WB2vA8bDOX6
ZgyelR8apN7flMJ9JkXOct4AxmuJd3kB6dIalK2lvd0Tf2Gj+qaAWm7JhLEnfbICWbBuByOGN5xO
jL5s293tduTPWdfLDFOr++xGxnlx+vThA6NiM/+Hg7Js9fdtfLIpPULnXsCUFAuqLkIJs7rAwzPC
izj8dw8CUlxyGaSBYCIiAIz/6lOj9fD4k4Ibpu4PskM7WBTGpya+/ICEaGmR4nKEcXw6IZscAsh4
wZWvu5v2oZt8jmtFfMOBgP5Ngn/z0h5q0nQ+yr74g504EB49jmAqT5n2FXkS8wmdbuYrhyAnDnHF
Drxi1+5e0OnkUF/8yiW2Y6KrEbtsvVpImiVqZBy/sKRI68ZDMbumbfMqU5HFOOs2SahR2ADG/T4N
bfOruxz9QJ1kc1K1HQ/uqjkUzzQFC42ER46cqTmNTkgWFoi7neXTxQ9pDjrAPvDTZqRewsX/y+WZ
MA1CrfAEly7ZzAVYSYIKtRqR7cqEkxEJVJRFdooVsrWakDe8xSVd8YO3gT6cYoK66cidAG8JDpRR
tyBgOTt8L+06P9Y8FpaBv/5VXhL2ZAcGbTCRDB3nLI6AH2yQv7B16laocZAPYe2BAvFvFcaDXvw8
woWV0awS052/eD/QjQrrmgOFhBoFnThv2otcfD4s7yREOD9rdnCY0c/IxYTn7uNNbY8id3R3NPfc
19ixGIdRvOpupgXyUAJ+sd2Rd0AXKvtTGqV6jstL7YkFNqahbkWwYCYvI3ahbPOwkiZM6KHYasL+
4mTNU0/foXG9Wbgp8UgvzW9aDT2K/lsubE2oBYa8D1BlUwn6Ag3bwdIqZHvN0bvrZ3/DytM33cIi
sXl/N+EnsGTEQ4Bze4JXniP6RQ42Nyx+FQCtwSaw8ljSlp1Ls+X7J5zH+QQenHPLIzonwXtKwloA
Dy5PU0QyfO35X5gpMvPlJPkg5/xzJwYGp3ZD91NqmqJxEV2NSwbTgWvv+9tKVvaHIaMB0csILf+V
obq+FS8Dll5Ah8L+dINP9wuS0lQU5JE/63nkcSFHWGgkBmNLAXLT/DGwJJn7uEgisDA8Pq51E43t
jH1rItkIW1z19HVK+SXGTG0hFM0xUcVT0glKf4qB+94ND1waGrkx4AoShAmfRVDSZ1jniYfXY+zZ
1J+IfZwfXZXeoFCbZzpvQjDbn54wx2yKRkF8iPbFINqyN/47FMOal3uLzD40Qt1Yp2yj5po3SFsp
3h7w47HHxOdfXVc185Dyi8XtXtos6u9siA1xOyDXYVvz25O7i3Sxu5MS8vAZN5LlIe0mrgtFdMOA
H6DLU2EAvtDq4FcoEbRmfOOZW7nCvIxRA5mqZeb4H+VPozUF+sRMAte0DzsBQISIn6st3pu/XLBA
w3tZ/Bn5UX6iuaTt9ckzdronS276Ol5OkAmtZqZVFrd2DrxhM7R6ohQrq+nFxeWcQKUwUbQ6RDbl
Qi5rn1kBLytdN2n8iWZTFJFL8/lZevPvlkRVYHvyJH5zWtpgH6m85WnC6Ah7PFOwPCUg01Bt9z36
vHX6Nodoo6bAvrLxYjjooknMx//BjKDojA9mNp/pNneji0cfjrLc9XiLyIUB1nZEPd8G0HPJc4uN
NgwFmL7SNmjOPqpmByRkCFKjmIm+EmUkYfLzEzxWbyHGbttHzSSYhmKpzuyM/r4vofzfLoip/57P
SfOc7jGKRGpnEYMI2GCg+d8fJ7IYPC+JnSGP0MAjbEt8cupAtO9W22sr8DBHy/oQgLR5Qb5sYuBn
Y211BhSbUcfM8KUAmhySXr06M3HMVpieh3LQeozq3HA4Y45v40ZcoGjs4xT4wa1tyRZym33SB4Y+
QcJfL47guvrwqFCKQXB+tT/5cFyv7fpLm4xvmMwTOwcT0OsYqiS3/BjgycKk1sTCsJZYbWM6v9XU
fHfDRdOzvXKK+O3I1wCIyPH46M2om+TWUH60DQrZLsqguf6S5F0z7SDU0/iWbkMh27mKc7cjtzAl
SjpG8ACG2NnVGjqv8DPN6Ik6sBevumlk1UBy6x/KIVigbFmuEMErxmZtj0uiiRMSOLC3tf0bDrzT
Im1agejSQkwhC/9uwOWdX5Yt8CrpSt4Gn/yrwi2EjNSZP8c0Oc1z9R5SWa23er5KICDTf/Yt7UHM
GnHpXaJbTveE75g3973Odn5pnlAGk3fFEEJo7mHSdpZaVWWm2Fsauz2UADnwPQ/7Fy4v98Qr01Av
rjaYg1+mOC5LX2SxVOdRVo6lXzzXmXhMC+loaFmxtCAgyaVfyhvbYh51wdmD2DnLm2ZCHkrgdwUb
LjRUKz60IfIGCoBS1t/cqNyki6jj1auOMscejGNl9Ppw7W7CpLMaNrePtkWaZVH8gmhQ0hlzjcUy
WwxCZTcG3imnQqvm56mWCauGKV2UX70hJp4T52l/Fm9or5AGEeITipc5QAOpejIrccQrHSIeyZct
ak1cXAflWRjhufT8yOZjaHUCDGXL3kh02uJaB9RPR5XNcCU6mc27TdcCA0OjZuwYER2XPEWXY4OQ
qQYr+LUbsX6EwKsfz/fq6AVvJ+hv58XAv1T/IRWsl/6/0jsIBAmkBKQR7un8JaN/rn2DE2EbPv4w
x7sKsJvxf2k0mg+ech6HfjFDqn0Ja+CMbcG/pne1+hN7lSj60exR243Iqjn+jLL76Ds4m0jAhh6l
EEc+Knap+SF0GzmwoTv/RjC/Yb3p7tncNpgooDRl3twmftEadsrGGxmYxtZ58u4eH4mL0h6v8vM9
q7TmXw26VYsiGx83lk7ypEQamincoe0/e5PLw8qBcdbyVlMy84D0PXzt9KI7Z5XNclzidwMD69kB
hqKwZPzdvkg5GceZepL6Fa0ysxl37/nc49DR899WmJaPPc2rHwqdJdgfGiKZuYJS9/nbUoEd64/n
sRo1fmyhttJAo5l9T2JjB/yMGGIURs9pV4bvYplYfnZT6xYwiUNqiBbIfCjy7HZ1glYCYDTQV4Bh
C9Fdn22YeXqTk04lfcG2YUyqJaLzBT9206noTVBSMZ9/kr9uvO61xXG8NS6M4tiTRlcfEbc+dFt1
gwiI6PLuTINUbFZuAYAoSECwGq+J+z0O8RKicpf9OMdx8F/Hycz3oRgi0aHX5UsY0qsWAu0Kiuv2
NnYlhwB57qnfH42DkvIy5f8v2QIiKJcgofUMzcVbesqRrwX3EJMnpK6BYlHUCal3v9gSdaVFJjM/
3r2AEtgglTt3DLbuyJWf0gL3y8Pq57Aqj9ccHe5twNADm9lhgpyhULqD1gJWm2X0i6PsHnsg9GEg
Pf2JhwPkzGSqMYDBewWNJAgtU2MeDrVzKU+h9yt/uPJ1sB8pXzijclHH/umQ8T3SF5VRyLojKXHG
3zb61SwhTaTkVvyu4OoIi80lyEzISrHzcoph/rVScnEZRpmd21nQlU/23lE1uRJVdugUx8cnWo1r
YNLVP2vruLiaNZabWECxnNq1DDVmSqYMwY8ok2pEYTyNJmv81xa1b82HKTVf2MLn5SAPpAE8mGzz
CJSUvWA2n2AjR0PDZfIgGXBWSn80YlcFgW+WZTqytN7sqkRcD80yEAJxvBlUbiAMkIi8sqqiukfh
DnWMbX1CqKNigis0ENSn/PdPHPtJpuV5sbzianFIpN2tjXPBE6+Y9nFJE0T9zAnrtxqD75x8qx/3
QHYebopioza9z6LhOaDsPMocOWiRuYGhMZvmzgxKHOM/SmI8tY6RMUu7hYMNtRJADJjh8kq8Nz29
k+O4pX+qd6UxUhp2kxury+dp0HFwFiF1/YYIyGWPnyNKYcS4x1qN5wVE+lzwry292bEK1Mwp9CfD
XIHVaAzvaMkXMaNc+Xt2QcuW7Asjegw2kVSALIHz/lV663xhgcmv04JCQ9Z0fvAknw/WUJ5Tj1BI
GV/1PvV1X+LIIYexSRNelkbQeaZILQTu7Nh7IswmY2wT6a6g7TEy7tM/88WXxYwjuPoDMrO2shDN
FGEuiLMtIqwOxTfC15IyHc9y6aCBF+KLt7BK1ktOheJ+kJ6Dlj7FRfE0RfafHVg7GXaC//PJLKZB
xk/kFfXrpxIrKm6R/PY4yaCaw8Rlpv9whVc9Zv2lBxNtkA0X8HoT2R926oWHe295u5W8AMIRlDEi
pVbUrJFBKDRv0saUl9E3siWQ8zhV1aU0VpIW0v+9ser5Sp3dsWul+xGZJ6BPWfqHr6usfX0izhtG
Rqv/mjNnLqW+yfn8yI58u3Uxahtm5QkNn0ayock70cNnKDQYoFOS2ALoF9OX6Fi8Zy6/hSdeg2tV
GdlJ1rAXaF0Ct5wPBlcW5MVUXoUmLcYCPP+kcMFtmJrgfn56T5P9AqvleJ0Z6lFihPoXjciPLfVL
9rCLHcU/RGeD04CAvsp7yS4y4MJOM9ruSymzryscuqda8+vCPUXRRsB1qjAm4ApsHDNTLwCRwRca
4buePmZiRp9sKX/e1EttRtzmtiVopR4qITvklSHcHxAEI18VjCDHD3sU0m48djsN8TqZCEhenNpW
jcpQ1uFk0GAJKKFfq2zi4kyi2jxFVScj9Mcackuet0ktpR319RCobClCKbyPOU5LZmAo2o/bLWNS
p63LJRHgiuVrECBLwLEQmW67bd+J5yAuFKHyrG8TlyDt8Bueia6VIs6Jn639qbQA/mLvxtbbmOTk
cZkc1XjNs73IUSD3kfRtnCryiw7NqoqMLnsFymaHzRjmv/5OInJesGIjmTmIK31YjKt3VWADJQ4Z
Zb0M0AE+ioMziSm6i7AnDEQRdZhzrVBnUov172WG3mydx2a67s6DHkFqi774xFO9t6SKJl7IQPCn
BIHxZGFMWxD9ClpVzfNZW6FiiJgTsXqA7kPDVtUajWvJmYVwCXOhgQk2Ph8AweAswggXt9XqShxE
09q+qiKQV5qMEFK7PIsObx5BE61u9qr2+GKeOXCQjCx+tojwqJKYqA/zpCCWIt+RbVDD7b33SYJh
4Sn30SGXtUqIQ1OrNejnyQbzPSprfOhlJIOCifFgFG+2h/IpWF3SXOVQ3Qzytv/X/v2oNGUz6a6D
+PzkAGjmc3Qk33xhk4Ura3buZvlh2kbM+r8lrCcIR8lksTUhQpvOraiqGFAqlbBGnwKL3afODiT0
tJ99AwpWbZg8r9sjiKqAsuF327nB3b2itwBnp928Ep+yyVDvm3x8RzoKwoVkxZ8qhAHwghK1OsZb
RIPwC+k9ID5tPoTg2GdPH2Q43TvVCmNqByTHJonZFzQxlxeu/CeoGooEh6iDFqtUPDSMVnyZlXjd
pROAJx97ykuEyW3YVOmhfWnpPkwP7ZMOXpkiVGyzeVlnPipfz+iNkVIvg4bHwu0xhIWQJyqI25R8
tQsi/ClHyM7Ijf7tpsPa6X39x+drDcxQyYrTYa4ZAv7bDNb/p0aFS/EZBH4SNjhNOUPz75zkui6m
gu9sWM82f+nPdfNBs9OVbP6Vxmy51pZ6wX13FsE0UC2npDUdXCs2jH7q1c9XQDFwcTcArtssvtaM
ixdQd3/iwU4ziCYzoGAyRdkiYGjRCEN3xDqsaPAuGcA3refQJ77JWwigaEyT66ZQionaVPeiZrZ9
tU2WJBL2lThPA73hqjKXBQ1zHCfi+WQJOWVLoSoNfI1FB06obR8b1AlCSCa98Hv5fBLqhNT01Dbd
wQUYONkvt6A+tx9bTKQxJ40O7X8oOxX1MjmUfM6mh+Z/z0PRvdgwi9gR8mBR3Wx4HDy3Uxixwdox
r37t7ItJ5yastHqGSeNWUqIz39oLFxQCVnT6nYRWomeXdmT3tPXMbhQ5lxeIjjEd/zL0F53Dxema
AmAX+wkx23oPcD9gNA+vB54UFnlMpixNL+4AsLjQGgKEiuNhuOppdvt8ZYocYrG6QknQlgnJtg8Y
scXj2AvrHmkropxxnI+ZAclO/mjOeVtgqseg5PtTF4OKdTiIltiWevW039uGedrISp9RfhI9vf0i
E3ImRVeoUmpqJOQsybbWjCNoFKePX5KmWzbRk4GJVXvlJ9xNCXDnO5UVI50hDPTJiYlt8o/bGy7Z
1Dcg/aCO2YIaxbONnf9RZ8JcNWeCFEMMO8Mjz8trH49+/1rHS59akbWEsoY7x3urn46EhcfHCH/d
43HwUOwghojqlnkR2nodJtHgpKkZ6ERoA/qLfrrxqBhCPgW08i7wHOXrnfBRQ9LInXYbzNhGfySz
5SxTwUKnlpj0gElUHMfwJyEtbmrElJKRMKMVVtSlcFTqqSMv5xTMJj0M058igytSFqhlsHilgzgv
EWJZzvHbNSSVXo8DX7GyTgUKxHwmiI/j1XY+raCQuL4DfDyNKZ6vhtOH/8EZWB06plDRQPm5784m
UR3I8KW5xaa2CbGD7WGfdzO3LKViZi7/xyJB52KQp2jKvQng0bNWtBoWjH9r1afhpqDXsPdfo6ix
Uy7HWMe41tmCy3QIARsRlPrhn4bhrc1zh2MG8LI8TEdGeitsRhMKpfZr7P/3KjeZ4UgBZTRQoN9B
cutUXGjgeIlXKiwLHOTifcjCxwZ49dOEGwBnSbn+xYKy6C2F9RUVQlsKWhT8Xk2UhjvYstjIJmPz
ZSAtBLoBSPDXBSLM+MW81/iLmbCZL9JRB9H+5wRRGaOdQD3F58XcFYNIWkoU3UijDVkOfPFe1JTX
vwfStMI2m54sA1m7ZoLwON2fTHwt1+f/G68+xLcz3eppzZiUhV7va6g1uTlIc0qK14U96zHC3BNE
YWqFUFeB4qu8dQPVfipOKuHenXt/xeLJVZ/32JnuCYdSDCWA7BLwVCos/iL0eInU2xVSOnCmWU1M
fpNuEt8kvvAkEhabz2wFyfpz23DiymimRFgkPW5d3Cxq/BB373DdJ/VQFksLfCNEPgt9/LQCa35B
CfsWhBv//ABWuZQb3NjZjVaWKIDv3en5op49R3COxaR/zjoNsflZ/kgMHzkFQUKFFsPnAgE1qfZl
OacbtIx/7giCgVRjvWCp+oqI0ZvvOlskKwrmnJcM8SO6ulcAzbNdDbQx2iYcnvJC0VKK2LAiCsvq
gGLogUSx2SGqCyX7W6HqOhv18fe9XtSJmJ5yyQMoumk+tUPMIebUtMapJJRY1n99+QhXGRO/BBmw
qoIvRejlRWB6z9MqCLzvJtt1/uJlq1e5miCWDfdRW9oDnMuh7+tRi0A0Oxp5Gt7Ra5XVlHIoK25Q
TRrPbs8pMcbW6mQz87eh1cGs1VgXMeyxHBmKUTo5kW7DwzULyxLXauogy10giWM5uoNSrxOXRNEP
LzK2CxXe2lrHcRXEzFKBSdipJ4j4yjNHlRX/dqoScKUV0OTx7s5T8kr6QFVjTriTPaNm9jKv5rT1
aUmC2UClDI/L0GoLLjbgYDSfkN3L3c+A3y4REFnVXgeYRCNOK0drYuVUMG6CCOJl2zLFmYowkugZ
UQHgH9CMUvcS6LDpNqV1wIN/vNgjFghqL0s1GJkePi6TbVEtWa1lmUACbHywn5Y+IMQEo5bS3Ymt
usHTuJYn7mcrn2B3pifA6HCoRgh7ar+LUiekOr4GAX5xKnAU9gnUsbn7Qb25HseXO4vwxFdWrYCz
VIfkGvT7HcFqkAud933qVFDTv0LsGww2P7LS5UFqHMatPHK32xjRAXJII+kj/PoyzvNKFJ1AQFTH
VXl0pI6YggSpPP/sauovHXKkBBbTzBWPuMtisYx0WP+dCK1cKibf+/25aWhnspaZBydDagY5X2P0
Qj34AUV2wljfT5GiH0T8RxKJA4AnmM/QyrBd3UlrcPH15SrjGfM/eFtIgRCHDUS+afqd24896kQT
2ub8UsxZ75DbTW82RjiEr73qov/jOLd4sk3TXqn6MA/XaZ0aFuXVZbRN2R4f5lruHaZoPpJgiZka
xTUyM/jb/K62q9RqzaZzhKx6fiDqMrWcm0mNoPkrHcYabbmWiC0GFQH4U7At0rhDvgNKlhNpOYBE
DvUBAUVfmd+dC6l5FNVpNKLMbncgdnppZybXzcFCH9KvF1VhHmGUhIiCaF4rIx9VnN5b/JbF16dy
27JdSGgkcpkWmXhA45Gbv1osh8HZa/D5jsCRcdr6UBfl+k1bJGTDJnZ0tn2zmR7sRVRzyaxEyYqC
cTNVweW9sdGbKP1iIbNy64Jge8hcp4XTHMv0qO1UlzpFQBipKicvJBrdOjR6nqtnVtmr2G4CgT86
4fq/DfR4doF3qsUWRDjZeMBpwA5VE2zq2+O+MvF/j5+v1U0CNyPG8hpkO5bqknuUn6LbO0Pa8bdO
r30FpSStd3SaxnuJdRgHilJPqCmjL8400cBBptNw0CpxKOcvpB6Rd4abuePfs3kIRcYA1Y5+089H
Q1IovOoseatcXB6j5I9ia9kGAbavXKICARhIt4OxW1qXvyjL4tWXGyMO+0xbVyue/rVR3jRzqCeX
RBNvFoCB/Uu5G2EXLiVaKM+hFy9fR14PsCeKXU9qbANOQfpI3zzzUVOg3ySJ7dSQ5uFU+P8D98Ox
T7lAW5aGDRY5O9QVjSHeX6AwP+wBDQ1+klZJSPZfwIR8UCHEEI80mhoSX10JV6RoqgDDBwCh6Oa0
JxnInPwWRemVdaUXAPho4VGGLRzgIi5hnBZs872aKdipLeehuYe7fQv3YMMkWSDp5TUeSsYISx1y
YFNd9KlMT9NdBMxSATfMig1Lpp/eSE4uWnsxBPx7CeQ94dg8f/YRSbU57JVMimn3xCHy7lho8eOB
3Rslqmucawn5ByJQjcZvCezWHioFKCfoWjzLASnSaiNVC5e4e3GyQQiXRH7Zni/IAx9J9/SHWIhq
C/Nhtk4z22nvBpKD6RaO5XGasephFXtiQBLB7lsZ2ARxVZXsBrcOA325PZ5EvjOU7H6M5nlCJ1BX
D1DlgduEEnNY9sInjnELAV3JQvzhom5ZAyxIwdtpVF+upbjtWZVasg2Etumhya/AawahpU6/KlB3
40kT9WBqoVgr3my2JL1V4MbBZ2O6O9uQJQO4cHV256eXuQ7y39nsWOXyYn1N9GkrY9YcG1dMGkhL
m3x21XWdmBtTBVPmXM1boRsxsMm9B8OB6mfOKY4t2UHA1S1tjgkOn5UjfqtF/NvCsz7eEaCp+S/g
n4Y8mUIOsmQFSd6lh5zdTmvwdmKMEj2IlV2OwbeHAGU+t13Y1X/RsFfiX0tmMONOsOu7EPSTb2Lb
4vmeeL2Z00nD85RcCTvu0TVmoGxyIHeDRRdY1zFSmvHSlaspT1pGEegiAl2TnsDgWP6G6WywhjIQ
ihfeGvtShrEjhft7VzUhkxl+R4G6fxqlmtSQrmbn/1EPDCN07QXtGlrbtdhgcAmo+KhS0AYMNt/V
IgyzSAcKcxrOJBhK81zSMFaSfoNi5s4qfy2yIfXR12FKkWw3ZAhKDGVr92YGODg7CVp9WvLoQjEe
HfwEHXv4RhPI9FE2302r91QaLSwqRSZ9RyY44YlbG+QPxdOtxfI64SnZAKLROa5m41elpOpB1X8q
MvZxRAr1VNzggv4Ibbi0jP+P4y+VzMrmB+fxWIDALP1itQhiCBRjfEfWzMjU50Cbn6+VgwR5RvNi
A/panPJHpDidZBok/8q4ZvvY25s4pNJASCuz+ILXYe66JqLltMTSd+QDkzUo00xhSqfI0O6frqFn
KLe073XYOHmnLuEqR6nsNVVoviftdZhV/00WZ2pEIVyhQ9Dan7oa0gNi3eY2J4KfBhddOHQ097zy
8R+sLuCcw4tbaWf6lkIM25OVI5uC30lnchIhZtZhDVdofho0M8kY1fGkOMBZn/u8RUk8n7Mi/Plg
2gWXE82TzhESK7CA6YtgTN/uQNlOCHGvidSbClHSjAez2AroG8Ug6zpyVfzv3BCyNw0WSzp1qd4Y
fUbrpmStOJZKQOdCPGwajRImL5bZ5yeRUDACIi2H29gYY5vmlbbPs6X001ZAGYgLEiRnHSyr+3hd
nvo4bE8o9tWhJZlq1AtpauvtZzk8hCtBbxa0ejYW6lb/7VQGqGH9UrCGDItRmgj6oRKhKdLjDVZ+
p260zqQyANXkLkrSjhbsFo4bGa+kQb1FxMsYNgWx1iyfEkHRmeW6RWn7OyS9DhJXJAVISoGJZC1m
KJLfuMOj7k5zSbjfcsx5vepy1bvJqrEjzr4Kqf2LAbdeFZ0BLAxOA8tvoQSM2rpnDu2/MkymyFKA
qLozZcHbPZincRuInB+CfUiIXh+1SVK76QcDUKQzaAr3lpJeNpbTtQAIsWUqNYBIGUyuhDQxNRl7
OFUDXVO7+omV3Nl9w2FIqXgENcnKrkQIiDdwNAPdnN/avjyyg3yZX0kukD208RBAz/avrDQzq6S9
DaFSXex4U7nrd2oGe60R4svmPSsrCAP31WQuSVG4u5vdD+KHJ6BJpnE+m1g4WyQ0bD7cJrEtTWcf
pZzQLPaOnLN0p8ib0FIELCOsI2jHjW+3R5oSqtu+rCKS8dI6v4tMe3E+VAjOsHJmf/d4rGNXoUzS
SxhwZBAYszidtEZgFOSxeNrKmdgdu6/wUEHAS9VMQCd0Qrut99D6jOQ0wtz6vbGsaSyu3hAES+VD
30Hr56qUV0rRmmgL+WUEiB6bfISar5WgBk95SsCsseki6beBokNJ78d83P97YtStyCupIhZ9qwxF
PtZY7AgD1wHgB6C28jJgaXSY8dVvw0eLlmfmLD3gQhJamgLgt+9wbJu+n8T09qDFIf6Bv4iv0NAF
wZH7hNZV5ca6cqlpVBNgUcMKJ7Jb3rosbhJMb3gELL4LpzcyNWeof+Xu9vYrOFtyNUwGBbjH4zpw
AYe67BV1ulD4QYLt10a0HLsajXwJg1rsMKAPGEFAsylm2Uuz+fqic/FCNaW76EMDYMwjURLX2TOy
gMkYniAXorHTTyTIX+rYe8mD6UcVo8WcjzGOBvdQTwYvrBiPdDAObd9N+RA0lqQBWvfUhSztk+xH
2hagi2YNmG0doIwEFBGOu9djL8wz3xAM7pavOlPPd6sxWUlOV0K10dfs0dogARfdV/blkn+0fG2U
pG38GeENmeC7XCrOmv/oN1/C/pXtWInpWXdrzlUNlpGtFgLl7903cef55SU7Dpn0eibwei1gZSeB
u8xz4yMJdCzywgpNw+ypqn+zp9LPQlXSyjrFJ63wml5ZdxqPo+mXCoBjnAiRT9lulcAXUm9u2T5n
PLmp/wBqRotsEdWAlJ5Wnibal2SIr6DOAAzIr4YJvK/hg3dI+02CLaFH2AfOT+WypZ6R08oJL7GN
HfcVBKIsNJx+Sv1v+RU57k2WKfqM8f1wOAcZICBxWDwpTWYiH62I27jzDZljxT/uaRXa/IIoZqFk
0K6KoTUsfHbWh0bQwceU06k+9zVkTrQlpZgO/uFFl482NqMfTKFE8WrQG1PPudursL3TLM3QKqJP
ZQgDK52/hbGnZCnG3ZC/r5tFwxYj11r23hb6lm8A/x0if1+bIS5GMtJu2KEAsBzY/P+1FL4/x5KL
5K4x9LKhN3sF2+cm0ZatD38npF6KgasHTZjWVwzRfoyP0DLOYRM3jTC4WbsHJB+kUiOgUxWhpmZQ
3tkTVgjCtWp8J1VDWlwgxbJ6zY2I7+8i4dpBIYT5Z8aB92dba/5KUj2z30kkMqiGebcttcPEAtBW
rXjEpkO92SIbdx7ce5hOg4fSSymLSeMmJ1TdMQOQ5ACOwfVswCpzi+W5vi+p7dHrfaVH5ZECQ6Jw
nUWYIZrOvLzmqeWA81xxQLCUWPRkBugZR3K0Quud1wsuCIvyHHxdfXE/YHhHVFGFODM7/KJLK4YK
61naBtwXzf/zUZzRUMTL+zRf9EI9Rz4C34BjrGVDpy/K5jWYkAXQfBp3oqr7ZuaZCsf0dzCgFbV1
qfWUUcrJ6G4XahC4AdHBSyLcZ7LDzszyDVfHDJmiJNL9uFTCoQK/v9Be4j3WSszjCNvQF9gS4DQw
pSUZcpJdzck5UPdCSEjm0rtqjLWgIfZk8zvYq+v/Q/uK6oyECBEyBUuwtVeSYB8xWSDa8u+QGFOD
sDUN0C6hoyiwFW66IY5JmiUKnywSn9N8kzia5tn2QEIXSSMWcgIh62IPCTJf+TE9wbKlVeNi/ZI+
DOVyXKH0+RqVTVaS397NPC2G4FZL1q98Ky//bIlI/ZQhxmUMWqrwStSwfrnLk3PkvzIxNRlXxHlM
kJJdMtjIBJ/GfznN0589+AmPTlUmjg5IVGxE59fdng0wF0Tl51icRrUW27juaFiREAEbXllDSsg0
SqStaniHiDt4t2reG4zwVtDMInjlqUD5Y5bs6Krw56ssla2OkAmO77n+qrOADhl98ZYW/ayoaY6t
wj09UL0b2eDZ83rgVVtnVZYw6PeC3tN6p8atfitnCEUrAmMJvIrpVMwsIwMzPL28/PN+YWwlIs6o
KBwN4HK5/qnjvMPN625yUf+Y1weZXx/M9Cl7UDXc8RFabtTGIIsLUYR3LfxUMk7FvK1PWcBdPDAk
YQr2O2nj79xs0txHSZq3CORgE4AQHfnMsqJUnzoSxAqMbyvwFEShG7R++QJOhndeG5hkUc0yDW3c
OJrcQld7i9qG1awj9SxSg9sgEA6mtopBy25qRj/schMpn9focG7DmUgIfXsweKxXX6JGwNQQxKVI
JEPPJYAWRkTHlU+RXmXUJXI5v0g5AtChVntaFhlaxYOgLDUqvwGKw7lB7Xn3xzn3c6l02CeklbTt
Ffmdc6FT7/zXmJBBYf3wFQxGjLENQ9hz05gi5++N5b20y/nHC/nMN4MEvjqKdWrwf2WwgmSdegL2
rkRiRc4KcPuje33g/0pBq8t8mcloEMbtX298uz8ve35/bSzthSBCRtuF1iF0zfG7ySH1ovMIpRnc
+xBXD6MxuehhSTLBI+q9NqkEqCGF5blaKhDEBNRDE9X3y4r4h1qe8E0dbqWdatsK5xky4Xs12pX8
fenoZZ+6GsfkSptDitU1hB1BV4DtxtXLju4RVk3OnSzQlc1LOXxzTG16U3GmuLGN03g8SMEfiteG
dQKdEE5nttUql5B3GPQh//wCiG0Ldl2KJmUlpnP3KVneq4fFaCmLZcwC5KImTV9G4s5ib33c8vxS
piauoS0vptRV02CHtMO/fZsQX09Q4RmcdIT4swWrqec2a15JL0z+GEz5ARHZJdo2UAgJiveXDsT0
jicV4L9Q829WesgIOTTgzsoP5pExwmlo3YpmWBKRhxzDneSzVbYXKDQdFCRxDsSaVdUhYjIVjCix
B/ZPqTAkYYVm/4fNqLt36PtjeE4ON8BNB5wb9dvw2eJAcaxhn2tnxiTdg/YxhqTZzyvYHVSaqIxe
xw6Y+D6xQkA+6GpdXAQIc/pcKghrw1LOLj+l6N4knYXOQGfA79ET7MZVa5k9zqMpHbjBgc9nVWO7
keghSqAzhwh97NMA94cwko9tmQY5fS/qYeLvboWwnEhBeSz3jKjBoj2EOHI+O+4t5XwG1YWSsCct
Toq/VqqB/bBOznVyxdXTWGcRHM73WBpkOLVAmSJ1cDWn4z5H+Ni/Dx/qNDiw/laNzGqrcpghXhNY
pucYmhrjroG8S1TRxiYS8uqh2fuHwWkx0oTsr3mnwweKgmwePI5nN9UJIucJ7MmVPlmcb98ezyWO
EURNMqL7TOkcWVUoYusGRY687wBHrrOHkQuV7WE2qtW4ofLbU8iSHABIxOabV4BtfVRsSI/Tj+yA
dtTMBpTHqSIELy/HhDDaz8JcgF8QGoFZ+yoBd2mDHi1TLKU3zUMOlk4H/E+GcYk98Taq1qUlr2F7
VrxIdMuenMt2XuUePAeoZfm7bK99wykkQUu83oWuTVZyL5+Nvfq6eEMHMRSk1Z9Z8/ay4Y5vIAGd
Mw3G5enbuW2tKCcW3Gi3wgU/k4uPyhj7GwMoEEH03grbYx25+4i7tDjJ7DOsjA2Lx1qkljHfYJmc
SZ5TvJRd97kJs8ptcGozWsuyx5gMT+1UrHVZu0Cx8STzDjIFJcQEUbYC9RssuvHWu410OHLcnIMb
Ys0+Bb0xaDYCdrPQpEJNsxWxKkXHcntsiSpeOcoD/T7PT8iXZn8eK9kt0zz2BNyMD52/b9GpUy4M
wAp3edfyXza+lETKTdy9LK9nPzB4JKhnKU2xtR/zchVpMBjlk2Er0JfIF8j8l9tdgEZicXXmUL5n
D6PPQcqVGp7rG9xTrAo3VsN2ijZUduiMwM5qHLKM0G8bY22t0+aGlUrVN1iqKCJRbW2N/rUrzenN
4EUwO3b+EBHHSjV9dYn3nRI4zgCxCH3M2R1a90kJYGb58R1/+AoLG52AGT58J4mP+WUrhBasu5T3
tNNYjnQLnWYSCAu7wqoLfIknyZTW3kM9unSXcvHnDcTH+QMmOKWhaNOMxbLRTRBV5hz8DctCTCOh
0jUFkdkRzFdYJXEePR01tnJEZQoNGoGP/m92n23Ep/TpgPSiIPJGT2hI5oVevjE9za6Zx4wMdEif
YUy3mY3f8M6jTJuRJstRhQeJqByJDnRxyBHoa1D2ZEH5ovpM8AUPItmgEPNkJnY1/WSgLQx49uVg
1mf6i7x8Q5lt17n263Kq60Ywhik88fwZkBJki42vi1/jSR1wdS0F0KWSL4iOs0xEgzau7WHIP+eg
pCv0hGnWWiyZlUxdty0CZzVGr9LiNDsH2QJdwl5gQLy1/NXTdsEDWQAauGKeYHvQo4SThdArWFDF
PaJrY0WIjGJyLLmJjKyn1Ekl5Y9qJTsXGS+/I2BawMU3of4FZbg4H1RpyworhXU1278M9lVaWx/b
VUWoUWKeZRaM8BaHqUNqhmvZ0G5/NLL8+PUOFuIZ0RJ81Rba9GayHuaAknxtsKJcyh7uH0z0+fDP
UB7z1WbhVeImCgfHrJgTKTVfigHqdBPEtaxIzRNH9PqIVhpWwL/eqg3hxO/PH36kvzgAHrRw8sbT
f/3kHw3Mo62iGr2y8boVwNll9Tc2K6k+24D9uCYciJBuM4wbSnIVfxSb9kkGxU6EYir1GV1BaBEI
C5DzZIBCpBrazc4fALvPPwpadlnVgyyeNc3c77LG5I4BTPirGcWeKhbZ3g0xPqODSvYYGIaKNM8H
J4VdWQMGSLdqLa0B4ZzQNc/X2e3T4D9MNraTMbs7Baowah05GWGwlWUtytEhnm3zzqU11DxA967V
+orCQEHOurwCMoB6+Bdjp13AQT9EAYbszjiC1Hnuwmw3zztF6SJgqaDf7/eIVL4v33zbZ+3/nYPk
rElXuxQC7wuM2cIY0/kBsKmKzmSr+XFUmS4DOD9WJQ0ukFU0mpaU+gAMwHHbnu8LDL12Wea0IE52
+LS92V4nhPwFN8cD4g/0fkKp41yyhjR4ZGuOGzkNX5jYIPGfy6yDKLj0c2Be63ZshzaQ8xSyYkJA
80Yvb2eV/ZmwmUqslLQ/iGygk4MJYUXchZXYm0ycjrbTJLSAkApzmHKl9ltqH+5GJ/b6d4EUGUeX
Qq0Q9Nsl/2gNP1+afX2M0YWOlE7rAQk3p6ccCZLesMVF/AFeUayKXm8UxGuFDA0n45EtRGG8iyqQ
R3kcgJMbYTOwR0aQSWEd1e2wXbJxYhxfYAO5+Xw+mfK6r/sLV78sgXbKUQKVzVnLHndXCZ3Z+hsA
4XCr3wsYljs/WfjQMEzjbBP0Y1wtbhLMoF5slo7ZoVNPIF8uDZUgdB/w52rLZ0KtqqMINGBPP3F0
l8oM9OPjDLkdiOuM7LPfqHki+givwSC/nZQ+y1qyY+FMG2W79jFSuYXkNCjU6jqYVfr9ihL2HOq9
ZSARwnLbYYlhxfTXT4u6VqiP5/z0hqQa337ZLoeQhA8seDq6rPJQsh+bkKYd2CjYVrwKnJQoFnE6
6GBlVdttOmmlu2gZcyGxpxctv1zrsbJm2mFSi6FML+iqmHKnbp3Q1lJTgQaGGL+GWL/ZaJwPp07l
rT2ncKIH+QgwT6QGZDgRlNxb3Hn/EYPvjyL2Z3Nl9j0WZJQDybQ23m8OvmDOn75wEamgAzIjNike
sYFOPfQhbjyeNMYOuxKqyKau/Q82hSb61UnEUeQv6FhBPtMF/EHQS5zOL8MMqh7LvY8pvHL2tMja
pMKV7HPHPifF0wSlwZDLqTNEfm4P50dAT1bN9Gcd+sSSEoMAr5i8r5gnaBLJiYPIM9fposyS0T7Z
6F0/MY5Yk64AqRI/K3ydFhzQxs8FT4J4hQj3KgH95kERupMctJ+WbyLh5o/R420GKPgFozfTMyy5
79zNMkG99a94Q/xNc8ByorF6R+LRynxwUkZt0HHrqh4QAplhiCtucc97QgqDtb/xhZKu7DwfJ2ya
xAqyXaUy+q6VgpAA9/fmGolcjdOXHxO4EvM9MSOLcsxK2mu6XFSLts/RI9etnA3pXdlUlp9+CfNl
Zt8ySyaeVcW1lQGtLAMEWZPThvjGhYC9NZ9qZ2UulBmP/M+mxGj/Tfg79ao1JD0FA3psRNnMq5ky
a5VcOdx6fan6wvsXyp4A0DmpR50X4Z1387DhZZ1QunYV/CxL5qbizxitj40UhVVbqU6Egw8rAv/s
mG5WN/hpa9s6PCgFLGwg85UNoWWPJQyBxFGM+sgiofn/0/a5+DahivDSJPEd3IJ9zr8mE6VL9WQj
OrL4ZfN/F6z/9amGHdIPo7vukijPWhNh4MG+gWjYWNap4/cALPtcso6isayahX9Wed4qpHwnQqZr
iYmDg6RGLdC5HUCk+M7xkKwhXvD/nRGHejBwVlp2lSs2wLob/Q7GwHpsp/4l7GXIZ6UaU29PwSEP
1UcBXRUWCjOBRCNAp/GvWN63mK0CTMiwSRwFJy7fdX40HDLwQO/S7ez5p3By/80BAVM44F2QRn1/
282yqwt3oyGjE84lFYFUbv/YfoAd7Quf9Mtd2dl4zJFg6TiP3vk2unRWg++eqjCkZpIYtpqa3S6V
Dhv7kwFRMWwyeci8QT28OX88wTVtEvo+V5sy/ZlySJ2RIIcrCdx4xjK7rdubLZPV+Pqpa0GlT2YC
gods3vzDY16lKsW0pUmwTsGBRSBtSxdT2wWI9aNxC/SzGuLTh8YzvUx8Pn6DIf7Wb0/kzZPK7zIe
oj95Z0hUEmulHz3NLIqPs4hcDzHfWao5WUnDFK08xEY7e0Rj4tUM3e/TSOIbi26lUKYZaDU4Ap5+
6CxwAUJwRFFZ2DfPAduAPhhToUw+uaJIOIo9091lN5wLt5NkTkBOkREtlefiZ4TlG954amI8m/CY
aCIi7lOYItPAQy/6YTGiBXBXC4nuLBEbzYxwCvLolSYDdUIwKwxGGJpk1L5jMoMUrtEdh1G6cmaL
jNz94PakPG6nPTWfW59D/Fh3i5XgOEPOkZrpF2LSpM8Ih6qPrPP45bxpRlDWv7S+KUfnYNEE6JAC
QbSoSIbQ/d18/AT3mFmgZOq1BuyuZH8ILQRmyY3MpslcNGmE1tCH0ZKT7dwo+ioP6ok8brhxDXdT
iiBc6kVjVacQ1snXlggoS5oj1IAK/YHJ34FhSnK705JxwF0uPgomCTmsWYvu99fx+bBZri/grytw
H2EC1dkSyyMv4RchzK390KqAK3yzH7rabjH+MnOokUrlEkQ074ki944lkidkHrlQ3yNG4SrMz9sN
7VTfoSup39l81e7SVaf6h+aGiszq2ywtVr+IS1sKOpGKD7umxGskzzye/Mjrs7m0GYslrGeFajfN
4VH0WeMyROk845SNlOHOOc+6iRNJ3SxCsp9F3oslE/5MyilSWzr+byMDpnAPtmOkxiF5I9PdlEnn
kdnspGbJiXcaGJ/1ofnE9WSrZVBwruQ0fO73Yg+PzTMPEn0EOJi4hg0IcKJKZYZNNYyNu7Q4hfvj
e17gRQ9wtkLo8PEZPQKH2DDvrntBCRP3XMxszONuMVAs5SWvzKUIKR8j5tOT1xz4EkxZT/oxVDgy
wFN/vcspa9pLZMGSWoo8fnNr16e7/zj0r254tpY3B0bxpaVOce94bpCKJhoOvoHVJa62LI2kPVHt
E62AgLpW1+Tg/7rg8tk0hpIpTKmNR5j1SYq0hL414XgB0zeARwOQ7EpkVBcmcBzrxH5B5iZiEjM0
u+ZRYXI9e2OaAHNewTxdm/YZJN9pcqOeORgl1AbqqFH2DYrQY68FlHZMhnJdsuUkdGJzxfb3Sji5
XUHc04SiudB3II5pOsrqS/G6GBCz/J0FDIDHAWGsNAnODF7bkckC/rusLF6gsvBUziDYZLBJ26kK
OIz4rzgY5Hjy8lUgHcF2I5gahcNKuseblXYG79u6FIs3UTjaq7g72kEvAmv7hJ2FC5d32VH7dOOb
c964VIF1Fmc0ibBzLwdwDMva37C1G2c01ulyCYpzWRxg2wQVG4V3tvT4gJXCRAv0xNGcpRoQpC9i
dEfzsH+h8g1UUA9HQN+9/IWJUeXne/MINXBK6ebFbVduDKMTtmsP1uxhXCxmoqFx5t6XwI+iztdt
ZW3sZKZkHnPdr9txue4C85EQKJAxqMGlHsUNqlO5ZDDJsDzgNO06JQlD8GVU59S/rs/zj7x3U6mB
VRk5q/1Br3ta7qUke6Ofu9DeG/cBssIFV50oezCEK+sdPz9ZfzoO86pVwEY2MEJlE6NvrYMDw3IO
qigta16sNtkRuE4UIpAI0LzITtuYppQsCrWDpbOZ5R0/AsTO6hdkjwMpHca6sRpNM5K8BmCsgoPF
6kIezY70ljGqeRnfA3cq7c3FXwb/X2XWb6vG3RvNUUivC1PvZuaIIBYHTm8UJZB3lSkxP2Di2IXe
aQzNP5riyFlxrgVjYPmSrT3M8UqweK0+30lkud32GpS8TWtcxUuhZgIlkbNQOtp/cph7LOY13Us0
LTNCs0HfsnQzwvGNv3y4DSrjlZUBzU9M6Ti8YPh9lwbXgnfdVzFybuEFMr4u9ksi9iGPPUZVZYVY
APOIOvs/tCLq7hzj5hfTmRHZQZDrUMgZhtdqqM1Cs7EDxxcUcz4chkfpE1aELrPkEKuTEhjKJhyz
hA1sfty5V62+Q21WYxAtmXG85LnlA9NyFuaCFbStwWlBIHzYfYgRgR3O5iJGVLt4SKPw5LYwvJwh
29Jk8tcbkL8PhiLZycCE/jQi0XW0e4ZotLaBItEuB6nifVw0WKpP9SculdFNFtw7tzqP6KBtPF+J
kUgxQqI9whXCVrCXSyUA+uVp2lFhgtJ9bOjvwTkoYaNAbx07P02Cry22wIRpGptc9lDgomwAZFgv
nRzDKH7C4uLoF05r83NsD105lz078LTwnF26LoeWNsIzgoiM+Al8ihRuE5qxSjiCWSvc3Vffb83M
Rf5vl8fpQtheoOaEFIzvTXabfn45mg5uJb2//sFf1dKS+1RrxhFGLje7k9A+ouAJU/9GAfTpXZL/
pb7H5ODbXZIxJX2M04mACpZiHyp40kweuCzvGQEcJJueAaXkWFHLXP11dxHsfH09HjweFhr63vRH
Gbj+hpHNCeBriBq2Br3jv3U1Y1bOKIPoKZaeG54VKhxcKPbbDNMTkmFK1/czfQVblFwQ9/OCljUn
jGVFknbWuRjSpEwKegzkTb2xyVGr+y0hY5hsN7L9EXG+NYmb3twlEYiiuXkep01Nm5sM5OIMI5Gx
p1nUZBxCDj+2REd9MoR8L6hRgj35ZUKhiW5JoTyWsk0C/SjZjLg+NRGfV2+nnCY9I8C2i5mrY4ny
KECWVgn3Ii1SFM0Iv6++CRjNu5dGX9Zlc/RvsrlN0aDvGcfnVbnx8BlEjM6EhVuUDSStv92sPO4e
+Xd1ClBr6knHteOZinOrD+RGjaFjbSn9CKRi/yFLsVHxOfIeISyh/NTagubH+SKjhvf/chIe3aKI
uImZECm7nKJ14pP9N/flxf0uIBiL3bvrWD81gc5LeBhNhI6yBJU731Chblptt709lpnE6atYafju
9ErtUI5ta3NWUyiwXamEdIObiWKveGtbapnxrT8b1TPloJcMssihGgkuwXiaAaXDmd5g1ZFdfFAj
Oteafc+FS23hLPsRspgkfGhnnvxRjHtnO24KuXtozrTzZF0vMf7cYgwvC5Ez+nih2Pa4LolBZgkr
uCwOTvu1ctHVityi87IQoBkTotWqrmMzJw9FfFPnLqR2i5QAdlLcvO0td7CNidCqgsNDD+GrWLGM
AiekzvBJyvz+jfXNmhxpG2fCioy3Wfo4DuPWcRKF5cIjo+pY5NCV2hUrbQWF1eMFjuiLWmQUCjiW
RrIci/DumNweU3TtgreyztfjzXLr2MgFc6SgdlesjqNMDvfGLhDQUMrJl7NlEXFQ6JI+AAe1q9jQ
7YssHzvkpnZOnnUZs9nviFuXjkaEb/xyCWZxwqbnM5cweLT55UcMj/LLfTP1IuKuN8j3PbrKILO5
vud+Qm/KA8UbcRZ9nBPu1SV2vlefd1xkzaKPCmzDo4t0a5PvO7AtQhTdZ44inyUCFupZ2praJbaW
Wg9miRgZUulRWbl1b9ev9Az68F5fyXaQwNLoMgr9vD/c6MTz9cb9T284a9SpyfIWtaiADV3YbuC8
mslCQJlgKgFYSC+DbC6O7MNnLCoW4cu1j7KRA07SJg34C2cIzCzxw0yefx/IlQUN6nnGyJcjWVHJ
8pe/tG3Xk1iuIO3DVtk/ZnXNtup88AYP3AwXqauynsS7E0QNc+/HslQxrZhEFj9Pz160ety6dyig
1huuk/GEpTshjBt7AG30qt3HjN0VXsztrVvF39rmqtnCmzT109ayAL/xOOA6i8/mZBm/seB56wyH
S7zbfWhQk3b1eW4/P5hsYXEeBRmDMQ02pKCjG1mHP3ZXF5wsExX7DIaiZbehUAr8+R1kJUQnCAts
N2Sw2XqyEdNWqRHVgcFrTClRgCQmHuVyw4FCkeaQk9dopicIxG6SMRQ+dampwZlHBzzGP5sqCzSw
7vZHBRYqMjlSMadt6pNTr4Tftn9w/8nUDv2U8NEVlhXc71d/0gAelvV5erM44fzTJ6U+Ow4xVjHu
2iHttebEVIgmD/h1advmWVOsrv7pnDW8cwO4aSQVa0bBXu1fZRHKrLWO4wpXqRd7BaRALDNqF/TE
Yii2b51StZibCvQaN7ET64uA28eIu6Ne9zBXuXCcrbaVlkmFDaSGM3bm0+k+0sxExCDivfjZWJ23
lStHI06QXBh9gchLtdj2Wq/J8p7urJVBnXMawILUyjDK0GFkhyPVEUJ1jJftpZWZ/oLFW/IFy4Dn
vFp+05LzMYX6lgUF7mDeckqcxD0azENAgYRJYU7oVbCUKzBDrSRM1KRAorU9gaFIXuxlG42dMmr6
TBYqiOaHcZjSZw4G7l0vnwxjPxSmWjcvFIRMJcXBnGEteBLhV1IEtmCzXmePk9BGMkuie4xE6G8G
o4CA4peTCIj770AvL5dMdUapaiS/QAGMZaWeFkqyFfR6dXIv6P7d0VbH9zUEZbps9uHNhQLVCFmr
N6u+prQs+HkfM6KykZIjb3p6CnWz27WRLg2Bd4JUySMi8fW6FntFBbZfvQT5DWS3yibU24TtpI01
HM/0NBU+K6BtiIdc2AYL9K8SL30H/MOoQ0luCxDlGMVkF6jaMMKL+F6KnbtA1cx364MbTTN5DNBH
haiDcVY9FEAp0lFHGogxsCSru9m25VG2OZFazwuR0Z84psQBgaZiX3TUbrscOZ6gyAW+JXTKpcP6
x13ITXJaKS8vSiuFWq/pkJrdMPCeWr1oALj+pCxZBALw/64Jf6L1cELnc6u12KtNlJ08SqsERG7a
iFWFKRNCiawn08o7ISD6xFNoqBdz/IlXhzycjE1Z3h91dcN8oOSoah77RHTkYxpQR5vxLRmOSqsT
TW5AkggD6UmFT/FHmrm0vxr9KbEAWMe0ese2dA9x2TkqTsJkOhcP0vUeAr+Zi97TmcBLVY9QdO9a
mrboAaHR2V2jXbJMkxaCB0Ex9AuBpn7P4pLMNvqK3QP6hqYLT6q3sXpJfxE9pRCXmUrnfrIoXMDP
swdckZjw6BdY52NyEfkzgerl+VelZPIVJ+/v8x8R/LpgZRPC7zIinqYf6IvpMRoaSTAbK626qSOC
1H6PnCUSRznxvzcDHZQgapW4hMvI+2UgoQCl64gPMgHWdggZyvMqD9v2D5onbKQDxOz6qRZ1ahbr
AptlasX7p1ffIOxa/SeguEfCa8CAMJkRG0BLMfxgx5c6gOEyIWOJ2YIYCXIGSt9hYx4dkuWe57gX
Mg4QMwOBIsY9fCbeHpSxVugPKy+uaIf0Coc6dGAbJyEsTZZO8hJlPMlW8NUbeK8HXaan2vGKeKGJ
HTLdm/DCisElj4iumo68bIho4YZ1n3IxQHllpLUXCFdJvsM/6VR0c2WaGJGCfj61BWe/boWVviWW
lsayjLZuw5wm8MCSt5FTdxOamfAOfhtou+lGMk7+G5mKxgfO0sk4Dsk2ZIUU0vgUvXow0RHcO+3p
d21CDvGYjw1B4JdRMQMpp3+/YFaEWjgbo6Gi88PDY8MUYhS+SD1verwnqkcHMVE46BUz/3mwrIuV
y/uIJdWrJHH9GUX4gAXON/7s8zaSZoaS5gY0kkavHcVqTAFNmhVc/5y0NmpO/U/tJk+T+FzISaRR
qupfMvI0xEkESyZoKvEj82Vmka9RLTBGm3EvCCozluQ+3OELxMimYZ1Ss/djFZ+E29nc9z8MRE70
WRCC7Do9sVepxP5n2AYC6nYh1MgPcbUpbI2uXAS38RL/xyyOqtWjUauXVTg/TbOzfhXPkNC8EB+4
/5BBkLJ/m3Eej6GDP+K+6K1Ptoqi7al19eXFJY1xelUAlm3nMt7dDrbRMdHDva9h8L/plAhHOr1k
w/C/A0CVawY+pyG6jMybqxvbUy55fsYl/n1wU9ud4j69GAR7u1rk7/ZaOJEoYNc3YYT1bYg9yJRC
rLcooQzA6gFevijYwOvLd0EitiuP/IPCydLwUSClfXVpGHHP/P5HRPjmwXvNnHJYJEF4ifMK9vAw
sl3yNS97DaOwYDB75fSsJ6vDEjZsUB38mrOUKCOywAbIv1SOzvioOcY4v7O8uUZ251ts/dmSgTlD
c1i2AkeHAY2EUDLAvBXnyZwnwhX8Ar01BZTEp/Ao8zT5gfYKFes8jqpmTCMkx6VaiJv/JJZQOopm
9Anjz6xQawXb2NC77swkS983VuDmtJsm9ic2kIDrM3UlFH/aplMEBd/Fxm6tfSowojsfqZ2zxvh3
epr16OG76bOLatILLtNA9ODSNk4HCiiki2/+gIISBBLNcsovhM/VqZWNuwQxuCkPSekNh+JBrpMS
KHzZG2nKMS83EmePE4ZcKpmj2TVY6YhywJ/DBI/xwFBaAc8iKb2w95+UeBhIIJ3bysS7irAEw3ue
c9lHQrirMq0JBR26fEQrRkTuQS/W4pqoFioZTLekp2rdx0WozEUZEotj9f6DBMqLlIV1nu/PC/bD
rTedRrsQJoMOyR+G6DQuEXpXvpdWCGUeg4JMwPIsBB3+X03/wnZ7q51ovu5JZWinCnHxl4BMzlsI
1Y7nyp796NUhEjUIyQWq4FMgw7dh8B0PFWRkvIxu9NiVpSBh1X5LIdXvx0TGPdjMoxCRKzcWAyay
OqBOZRR+VZd38bNGvLSCvaQc55nrEA+NvwKizaWzZQw2LelkOpi/K7JGNb9iUbvhlwCTSdmQK8zW
XTXUKHmwEMX4yFbtjcjQiHJVYWAVPT+SUwy6sFkBc331gad21w1tep8Pdl/zAjRmk/kWu8F4legy
XVJ7fkF66qdpEnkucNxxK0/u6QAI1/QurWezpMIWHidRcml2NJudozzyotevbe7hGJ8yBkzpCByY
BUpdfnXyROTY2/iiTgW+FEnFlTo5RM/NRfssuLO5/ZwcTWctiGqYQ7vDTp/uTpXUo+OFrF7OeUMP
zWw5g8Ip13UFAxb+jRg77cl187PQyzLVsQQYzQlfZnCFfQB3n1EzLEHo49Mjg1O1ywztcD41nadt
McRbI8HvWSCbvYcniSdgasaH5mM5ubr47ghWxShw4yZbzPBSBIJxEqLIEdpnQ5LeZWNQTCL/tFMI
FEHLyL3pCOo8udmmLJTgUv8pvJKp4IOLTOTwGZ8BYBwI9V3W4yG6tUDo2JAKmmDD6FIkoRkVMEFz
JMCwVV2ryfFN2FV/YjHsoqKstO6+j3VN3BJOyvINiSmNKLYKvNKfd1gwTaSl9JEbWOgJ/dojutim
2FbxlzCO1eZLBJMekYdi5RHhZx8W4WIXeLzcxa2o5OhYL+nMYEzOngV4jhxomSNct4tGpKJnTFc0
kjiYgyE2NtJ03y6+7zdxj1o178Nb+4/dpPurw6jpc06OUoncO4pzC53BxUSThJJBquHQZGbOST0d
zcJl1CvvQoKDowSQWUG8HKADQC/tKqeXL5yXVVVOmJ5nREfYyMUnj7k+lCqq/O6CtzGuQQL9ENKq
6H5kfgo+FGvXbdX91F9Gtc4K0haQ96sNrOW7kJO0WGLKUiMg2N5tn85HR5beWk25LuaOUx8cDyKe
v+oaVG7L0MNt2LmYMQXUVXkM0BwYBtvPqRYTQbkkYW1obV5xC1K+gYlu1el804Ym1YYYb/ro9tIa
s46nEnFdtlikMLaKIrVhkF0ZYMquBpdKaP7y69JUi0/AkVGcyTpsG+S4VQdor0bDc7RwyXo111cd
QdVCx6YHhHng2RwlVQ0bfwuSgX3v2AzVQi2VamR+tAVy3uu+sZM0GVQD2T7QRmhLxJKHLDAlYfKz
A7ewzmS5b/No7Q9/l8iInPUKQLyRxCY+OEgj/LUyQy+91xkwyR1L796WtLe1/EcAST0uV+2YYj6K
aqYOVHLDjMv7NyhywpksUQQlkFBw1BeQBtIPewgt/Z2bwRKz9LMBVRUFx2UyHlIHcA/VlvAw5biK
ofN3NyYyAjNFJt/nuj4sGPy0Q3acJkQ/oop7qXeDwLLjnl89pWsEqo3mkYbd6G3G27/BES1nH5Bx
LkqJsQUvFgPTy/VX+AIEYBrx/3X1EvYFmw4/5pp0aEM3KZpa581DRQ3lRyfHJlD/Krz0XkT+gQcf
J5Zw3IE6VP9tn8gklWs7CRslVJLik5DUEOHY6CJK8MTjAAB6DVzCXyKQ7DalDFKwMKjHkR5wwS34
tAqOOxU3jBK35S2qgFZA3qf6EBOlZ3IM0U1oyIXb7JK8YYnLbeFZ6j81lVN+7gr8ggQegD1QLqQO
v6+GrazqaT7+SzY6Gl86gbSZLsGjxaSXLgSFNYizMYZLkoOF8jjapi67ho95VinE2Ev0Fq42N4af
XFKzH+1qjQh7GFxR8XhTqnDwMv6Z2OzABs1AMRMFWDMX/qM0LMy5JN9YUtpo29gSEVvediFbrDly
T1P2IPtiLCd3UyJwyyG9YSDXoahOm9Jtc43uhKxr1QmHc6TCyxY72GAhyTsNNNFZLU1h8XfNXtB/
0wxt32iazyeRxYNQ30RTRgpwjlYFoJ/HO/srI/AgujsDj4aLCAlBixXJQKh7GRkcPgNKTvuyrkwd
1Aie6q7AD6klgSO4TSUs2kujEiJDi6OJh36fIQXzEVTJ6jgmavlx02eLnpJ0FnETXW3wA4JO5oWf
OskTJrwzZcXDwi7C2TKZKjcvZ4rDoc+eOX1aqzfnHxTDhi/ZoM7/2qA/nb9EfPp2UbhrzTcKogcp
O+T4K3dDqBW3bie8pk8UfGtRVIpJOfG1lV2OmYJVZvx/IdvHovF+VuRe9iHn08RJAUMGk2I5VXfW
3R8irfTRrS3GNye4d8M08zq1AhW3mVXMnjK+t+bu0nf677KvhsZkmBDUI2qJENnLLVAEZrcMtJ6e
pBnN7DjjY+HXPja6eBOFJ1atDSopWJaawpoom3611LsnnFQtUi5e7PicWHc3wCshn3gUfCO3hT4B
7sb7639oYkyUjhHsxbRAXON0/T5SK4HBv2o2/gFHfKmKUD6HisQ+rPA8Qkyi1968inM5xrEeILwX
0Jy+7761JViyDW9Ox3whS3i8RPMvN6j7i/ELc5VKtxyvEqvUv0R+lDfKaJ3hz32Sc3PIV2hG9tZ/
C6H3ZTLyldQyj2e8YS8oezZKijyKVVOoMqLnxttftfAmyt0YFZT+bh6UaNia2jS+URWNv6qKzB0n
WaFXDVSE+rtFOpCKQRaGOe45bEiSyBC/n/UJxvsvXxxlh77TGE+X8vzYMbamgeghe61nfDil3VGa
v6nEnAQwwaZDYkHJG7CDSHpO99qaXVOGlK7TEy9WnrqobSqpsHUzC+ViUKB0iSGbVsN5LsystSFk
XqP1Xd6MRqhg8WLzMr9ZDS6AAhuKIQaBHqMU8KhFQOo6TAnCfR1xlGrQYLoHejKXhVgQKggPGUsX
7hvq+QBb5zAzuAK29L7V7cj8B4Un4V2UG6aqQNsuagYic1K6asdc8rMdv4+jsVYhWjQc+81vsXAz
iyEViN2dlXMeLX2O8Ru9iqtUWjkBp5EuZzqXcB76PN/0VqlQRVY6ctMThu7Pyk9bmMbAWx5yxHb/
u/ns/Q9Y/XVaZ91V2W13DPN8Gyz+Ic245s/TdYG/p7UXCPIa+AurXYdNHkby40dQTZ0VqtnNCypB
vce3zLQGnJvVhTWeYxJ0LzPk5e1RwMqrwftLtiNTgtbr6b2XCVv6KlhKWGBmuxu+IX1fZyuaUtp8
ZMC/3+KsK0b4ydBHaxetjHOZolhD8kh3iaDr++6f6t30bpIIds5LqpNXB756wn4dgyBMB2T/ymkM
pa8ZZhV+l41rk4GGB1LnVXpqLPQa82O+LPj5kLe4PcPSqsLvaB9+/g2CbrTavWSx54srbM7c81kb
h/gPMk2CY2I4/jsdmJxU5xeJ9xREgclYHftuUQc7cyTcz/fIZIhBWpZb04S0ocUy+w86JWeDC8pg
t911b4wR7Sr3U2bFUfowahfxP9OYhUZIoWu8VQ/EYtP1RHVEIXjY8gtHQcwDgLPPz3FevGPmEmXm
pv+TaBR0GATeE+zRVKIMF0N1duckpo/e73YtVlO/bzKy5dIKbdgtavW1Tqgsr8XXUs5oCyj8DYr0
fDqSJ8PlHSppMKuyLN0N9i/ZQ8VgvgRGP6hCqPEHp4iiN5oR76jnDYcsK/ApkOFlVsSzIlKZWTlP
DNq/lyXi81OApHq2yYZXtihJmuoz09yLd88CxtKXYua18tt0CYwPOcyQQkJ61x9LGvTFIurz1X2g
iR0xscROICYteVcED4nS5ja9ciXU2MQd9UWtcLjXRMFlXJ8w591G4mgts2OOOS4xq3x0PSXpIr1g
BA66STTwEeHln2HRgjOwXBW6KyOS9PFnr/LTfsPHdPpDgh+t4Q82FQcE19cc/NpfakejK+5Z9T5Q
yOgRaSqElzIhULq3ElDSvsjmBVIu9eOqsj/jTdPb9N4uLCOH44CCGC35XZwSJeV+pssSO2bkiw6Z
ku5gQdJhCBrM3B8tNqzDx6LlqdDZUps4BB2CeaRe2sqBqCpPOuBj9e3DNUaEcS6q87gqOAq6hyDW
WlQXn7vYL6Bq/Ff0Vzct0oANYyE2FsNFcvJ81beyEdbSHFPP7AY1EVVL/Qj3S59avNFhHliiils0
OcUKqyE0ckyZRufKdJClzPRkD36W8jr2X3fqLHhU5yIUSuk9REkIyaasW1SfDoiZ7p8fpUUt5xS4
3XnlPVTjzS2gyZVvDLkP20BapSg6J1VPNTdKhg5YciOOt1PisLe5TtH+zbgwrFCMz2tG6BeX4/xL
36kFcBwIeb3XCsLjLBrfNyEnCvWQke2nX6yp/sAzqBnsyHkby9VkLaahi99bYaKyeNYa6DsgwVX7
MBaYHv5yM8dG4NetS8Vcc5mQkTNQppb9CSKVeIcTAy2LdacsSJpXOMeYAuuvHdEstjQDxSqwIJku
l0gIbtyKVjAk/cDgayTDq66oioQBC/baSIYZulKFdg5fJ1RS38fH8tZ3W5a/b/2U4qQRP/SJu5RI
VETogAefIrGt6OEN/ltjcQLc9Q77+98J9wEMmUnsKgMHkhZektZpGCAD4DEO1IIqPpPBwv5ltduE
Er+tz+aHGlhg24HSN2N5nBjTIIUDeWBemlt+5mrUlntFqJM1OFmC/tIIBffMhvaHpkh6cDLe+hT+
rdTT4tQBng7KHIdkeI6g4eD1wiYMJ1feThBU217k31Y0hhuOWnmHUqaTxDiXDDkTxYBHwfV/0p3r
A1PO12Mvy2FWv1WZBgl1VQ/d69ftAXk9o60sPz9nNXw4kzbhwEGn+/1/50f12WkebsxGzjThuCA8
4swqiWEPmWe+jcLNwsA/WrekwU1MeS6V+9GuW3Z2aV6LgSuoa5rWBjQa2LQkbfN0ZFomj90XJb83
HaF22SpNusFWvTLiXaYfSbchIKIHPfYBIplTvnnoMds3hb3Suf3LpZL28VZMGgf682is4WAeHVeg
KkYaZoBuhd0apk3nj7JdzkoVC0v6QTmXm193l1BGIQvxLiauJsnwLBu1FBmq+JsrGyibSspqtXz+
uppmnC6yEjuUlQN+8jiJTxJUeF2RqL0kTHGlySLjhR1ZwHfbeMD4G9eQGlz254m5r4OuiFB1EwPJ
SavZObXcYW/FHIOVmi8iTWgGWeGHEuGThkvpCcm5tVd9JKKLpb55aU97507zs6hYZnQ7Gtj0WLoL
QbA5hZasY3vqt8ZA6ovQGs2k12bnClcFejlpU3/VmVXGvlT0/W78M1XRjoUCSPaJMDGxgKn8c5JT
ZFfkEf6koHjTjlUr+G+R4BwTOGGetbI7igr1YnxSpNK4y/Vr/fb9X/7rU5GZdpfAuFPV+JnSa8wi
YXQAvYBXGjHYNz2VPeFaHXTGDLF9fwqaHWYdkyi76tMxD7aCJad974lvvIXvMvLNIJrwJd609scZ
5IqFVvfXuiDBaajF+4S3C70tZiUg/UIE0pdd8Mrc3hAEQPHY7a/Qm6zPZZ4YhPvav79LVkKftQsw
RnvDHw0Emf7K/X16gU8wt2E0iWSs82N54BaZSO/vtBYnrXP5N+H1wguGdSAKOfTZZ0PyjIY+GteR
5YtbHWPUHcPLOwnPbHIOxV8TU44SVhvD+Ydx4ZfzFqf+jPBw+fzUx90QuENwTz3uNwe+azokBE68
ZhWLfDyRqzaaHojaFNuazXM8KyPGE95xJIqzd9I4Tpn3V2QdvWwsUbECJf4XkJwOWJudOWjPz+cq
e6hKm3IR5/KinGWNwWi4EJT3VrgEG9HBJQk0JSbEXWCzpyeKzt8rnl0gZgvCjmqQx6z4cKZ2FM8K
/tkkzALmEIkGG/1qriYIHb/Rm6vcd/M1vQOp3h61+BhsvkcBp52rD5nguK5mZDMkma/iXFVOFPft
eLug/LYLWTVBO1aTTdeSuj4L7+AzA2PeB7HS+RQgx83Uu6dBC3JoaJzG6tvScc9UzDA9536+pmE4
JuTAkYTpk7F+sHUMlRGzNhNRq42hdz1dPcuTua370o3l9Nu44ooh/euAA5OCQXjaZYW5Eqwb+qJ0
89ANi24tXSFS71L23fVE1lt+5DNaecbEVFtb3j8bS9MUOC5ehIjhNXVhx9PME9r1LrL3Xqd1f+/n
rIIGthDr7v4jfxXd8RhNwDB25CWFOR28NpezDLI7yZJA15w2Ys39jqKKTOHFP8JApNeGn8lgGgyG
9ItRL7R9urYxfweF0j1o5tEayTLei//5+SOGgT02pM4gxwtQvFUj87nQoUy4P5UikBLADtTTMc9r
zFt6AoE63ftk5ERTmrXvh7jQtTml8utmT9C9wfFLzMMsuE0lPG7IfHwvd3JWTz1ogr+Wy5B11UeS
r7uznwycwcG+wuRChjDAJkgHbqmX56w90Nqbpk1ffyahYJmlkP10nSJjSaiDzm14hkGvZ/6f69Yt
D0dB4JdSmm62HDo2QsOvdVlI4yvSXb/n/mSJrrC+w88VLYweDY7VNXlKbADV6CQjP1q0cAPq5NL2
Rpnsg1YsdhkN8c7bVH8OAWVA4v1bYElrJrRfcXgNoxD4ITf6/w/4KbWm4ZhUHnMXzwABj42V+Lrv
HBMTawHrr0eNMeBDL+XXuz3HnwEvYbo9V16eK8/xGSvBbV1+BFc6JrKz+51457BqaXtNm+KU9Kck
miLT6mXZuereBu5uREfpuQiaRidHmdGgYhJpWFMLF0SEsw4bnTl99Nncb5l/qMDDli1WdbkI1gq8
cNjwcn9JtfJkz1C2v7tXrAb+NSwaBEfNG3l18aGDrWLgXlHLOWBBH9pVqQrC+kSE1lyNmHtH8qZI
b0T8yr59bcIeCnQg3AG4ik21HC7Uj00PtKvdb0vJ+EHfDVO69DXODD1hXqNUExr/deuI9Pbi7ODt
taNDZIKB3oiacaaJA3UicUEd+9iGlOL5ikPN7kOkRe4o2+GIIaWwRH78Nbm9h6sMC+AJukgCtvuH
9C+QBNxalBB36Xf7rDpcQ1NZ4YsWtDol+lTHcN0rE8mE8wdJIlpKOaMmXiZE6xJtlyPRi+iUDjmf
Ig1rd9AfO+dpgXI0b7CJf8mV+jF672QlGMotWurSwoZBnRjL4A9vx+KFD8QrDsrUZ4HQQGyALDwW
ELfaZsHsPvAKQqphHQkOpwRBEEa7c9Zo5QlC710LZocUXfHi1OIJrqfgc3NEnIweeKx04VUtH06j
4W6LTlVPp5p19mMPADOxwgW/NKmhWIRu6k5hx2Awed7Aq1FpwfuEJ4PGRkfSUafK+dYlVXc7Ya/j
1HiYhSoFsxGwIbITRbcwPrxBwJRUejJmac/gt9BUGIRTS6DCVk9fPfULNR7EPhZLCELAny+sQMz5
undeoc51aF/6yLh/MfY6j5B4gC0UDgRWJgkmbIoyKKy+/cZa80cfVw6jEQziDn9TuI9i1G40gTZy
S6Y4midLwgZsOkzVwrtwmg5WZAITbB/7mhUU/AKgkUdAojaPhc+O1gs168MlSgYDbXXveMy603Op
uCmHJs1Vk1eZL/fLqUQpkOydCVfDDf2m9zD7VAwcBpzNZuHAqdQ/TnmmoN2vna5Ky7LidRrCop+t
g/XiRZPfDRd2+Qhm4UM3cKzmuBSNP/C1vc93qVfdPi9bctoVrUn9K0/RB2pdT5xEmiwnhsJEYT/h
r9i/6f71RGIQm1IusFa9eHQ4VuhVAW+RqVB9mci+l1KC8U3lIpI6GYe0663ZZ0tBUY6oGvUwk5fs
h3AaazjTDtdLK759V6jGDz2OFTBTaf3+Mrye1ITfnEOYA+XBnog7RQpxfgg+vW0AhbrPCX/cbhJu
bOhxinefg7XcUfig5mXhW5IduiQzk1DWN5xuCrbWkRNR16Y68w46xsNxMjwHXmMS/fwhwqqEj1g/
m9c5V3znW6Y0BC1/96Arx/EvB3C5hXR8HtTwBlN2Y+49pVTh+tEh7FQTbPnPKuc09nsH6JvC0bOU
bxGB4EDTvo6EJROQNXL2GyUna6V4Y2SyDQ9evL3h2NE370PtD1ba/in0OiZ7XhpiJ6UWUUcrAhkG
QB8U1s6WYLAjLaFWV0BC4roHXVmAoSBRtSX67q1JyZ8PjQsGlYgUAn89WFSgQAzsrY8yMoGR4CQH
S+8NvUEpbZoRkqgbehv/2ORwr1NRwELJUVW8QfTCP8uXJDI5Jv7PmMvCy2cAu/4AFslZu/BBvLJ2
Be6JmNGc9cHFofN/2AG0FC0cFMQV3e9Nh5DqfjLv1UfBXNGke/b2QbJE3Bn3z/rpB9yGmEmC4uO4
Sxmr+ly5b0FyA1ucy79cawIrJKN65ysKjOQEIKCC8rxxPJDisoI4ijR8ZLAbYRXE0JQwSNJjPwhC
bq8kxDWWpy4GpyjrcKaEBEvphVUObuX3ZoUX04whYX5vz1IGLGW3hOgdPO4ADyUXkrlAtYl6/4Pa
4OFUaPTyvNcZLPpgq7zS6Xkm+SNV4DKIFCEyZSOB9mSdr7nHPof2RKLQN6bZ35mYslPxPlWsPbgr
+/q2enObn2h+LLDyDQhrN8QBu2K0Vhsg58Gl3cUbahsnNOmvrMxWK9DIjJLSL4R0Vh1futJYmKnV
QTSxyJ0Cl4dcCOD7/bbNjnKMcnG853x3m02XR44Cnx90tjgKh7LIssVp0P6t0RssEOWQ7ji7Ed9H
SPwTXEV8ufpEEgZHiq2Fzal9Eod/jd8HbTXHh6q3skxkiS2alwFlgwTFUqm7HEguXy684Cg/qMdB
Jipsyzwj6drXKxmidyGxuMDOevGbHNQ++9qMuko2WWww/0wocVm6pDxvC6tDxhYGDuejE+0dd4OS
OZ/o2YpQmxUzY2Yg/9+icOxpTWCY/FFKlDPIauXZaPu4wtzShaWwzXKXDDkFZw0M/drOcV8ckc/K
COpP9A40XXM0bbaYNQAzstfLK2ltSlmWdk+BdtIUmA05gHpaS367cgBmo16KqAR6KaxUHGU8uJfn
k5kb9ntu6AxbVBcUGIbrMqVVIKofTLhCh9MrCQWWiWlp2JJ8GQSCfB0Kn6lnPNi8WkdtwVjwMbAy
4kLLotOEegM9W/SuLVrk1lwJb/LAesWvDcugOOGh9QZeNpVNo5i+e1Bn4roq17tGEg+OpEtzh9Jo
4Ec/oiYAf0WuF8ahpDQp/DU2r9RwuHBOwRJVnJSFlwX+kGyrKsOuFnQ7GngMx6lb5jCQXa5v5XB2
lKtkoBP0IugZkB+0jKiEgld9GG5JXZKqapqsYluSg1MmnC/jitMwPgIR/YV9+AUPqvLKYb0Pn+IE
ioYodkK+7YQwyq/Jof0q5d9M/HFxJPyQuC1js/3FfhRd4Zijwh2DjzJiqgAhx1sn70kXbQulYIn9
5gMyhZbPW76Fc46X7Jixi92+b8d15yoLoL3lhx+bDhlzd+O8ijhujOAPqUx5FYTHgLPSMkL8NVgJ
4ewPPPn6TmJMp5kzVZuzvv+sr7cuqD/HtxrIiKHR+G+qtjSTr+WIV+6trdkwAdxKfrHtTVDqcFwr
svuXpsRw9Yd+mw3YD60NnEvHVOCUagzkIILoi6ahdS59D1ATYPaAcbsNEwMqWWF+RuN9G3Y2V4uY
PIQcZctt1elF/cAYZPUC3TpgMEJcEsFNK+ola4zS/NNaIGinKgYG8R6FA1/dukuBtcfgD/43GfwN
tWDN+KyaGdZCkImokFRnc6gWpo7NjpC4oCsYt+/3seyii3ViCDDXs+vNNTuiacIhFdOyDT06oxLF
5y98+D2/MHYC/Abf6J469ojBkpRKZEeNrH5ksKRFIW+aSd8bfXbTg+2tFcTEGhqlk/ABYVnAwt2B
oRN7NFSS32XXVGmayVGvmvI0QyQcPW1gtATqSTQIMK6vL3SvRN8WrjdZK/MyLUz/2J6YcE+2Tf0z
KLjvoyIugkHV2A4VNU7w4SrODxRQs7nnTPE9NDXpCeJvbsCrtHag2fO7svnIKJuGayFr7OG/a/Te
WCsvZ2FIAeaspPePR/VUPpIRbq4FaahKNoUSGhH4QPw9Nkt3jOsDeeWSehTM4qWewkUaWhw6+3Dp
5eSnSGKC5f/WbF/cvSKF3k8qYD16RU7XABDVK7iKHT/55fz73cDg53OjmiKy/K+GhLKg1M8c49SH
SXYW6JLg3zd5BNcnFPH3kDr+pfwk5PwXjAuA35i4hOCoZi5RRvE2ZgbBUkB8KY8yoWXRSAprONOU
cQUU75qDHpmxAC6aGMVWpiM48XnFdZEuuDhZGgW7AGL/FfDnB9YV35gTPGHDp5PZODBLBerjPQxa
h3CKWT6labGIQLexWUNdNL3lGVl88mfXG9X46iTmT+hpEMgKxE/Pl88DGc0GwycZVCON648JHvn1
0Fia+MR5k84PQ31dvyOZ0TFyJut+AULjlpakxL/tupmBQMlidXWVaoHnMAYx0OA30hDAyysv1hjK
BiiANA+dqcaLW2DE1CplOl/peEpEqxPqN1dwgAU6/a1jkw0EGNmB298rO4sqY8xobWMdvZRLRWgA
z5a+dOJcUnxJQouZYHKqDDnM+ZNWd9TicysBqT51w06sqCdrW09TuwBtTvpiyagFL62DrqtgVIhu
27Bxn7UGsICj7NLbEyjMGixsM52LClsyhmMAsGPi1kkefeaTYB+6QAvj73wXw4XkZWIKCYYy/5Kl
RDk0XDXcocizkaD0IA4VCgHSGheOemvkU1z57O4mvf3yB1ItIB327tvbqFA6Sp6ioNuDGJ4tTwYl
asg+2B9xrwIYbcTji6Bfs2CPY0r46txdIK1qbsqXNcC1RstScpVYlJQOoL0zQ3CvHaTYtW3/T1oV
vFhOIiCLpU/h+XTk7cQYB4bE5Os8GHgg/G/shZsK5a+i/KqJvAVc/uvLA5gY7g19x1lY6/g1nv22
+PF83jCU+ZBZZ9OUTJZByb4RiMq5rz0Z8sBJrGbKkYGeA7X7E/VSPj6z2xyT5MfYEGNKyL1RgzOK
vi9d6hR/ccUmMRCqDgC9mX3piyVAZenJQOmvDmQ3DWCNFjYG2MYuIFSCY4B/DWK5DchcYrJpHeZG
ooNWhik2x30hOkIj4DbmE8yn+iFsHvkxigyBDfJwmkAZAKdQcM9KgXUsfU3sPoEOpBTcrJ/dAlEn
mOjTbSkm0IcYWyhFdcXxyUAPWt/sp3aoPCo83A35GQa81IiJ0BWB2n9klxKb+356EECMR6xjoPwJ
NDKu8mlX5fD176cmB98vg0K1eJT1mucTTT+UL1rsUwAJPWo2cLUh4Xr9jPUYwi2aeyDcU4kSJbO/
qprycgv1FHcQlrph2H2mK2osvmiEts+yKULE/2r0u38eUfA7SzMhIyJWo2xXUOx+ZYQVkDhA+HL+
ctsqzgfQKgPQBTIgvLX2ycjH01yH6xljdSQfx0qMNAd2C6UxCDo1L4vLynZTb8gKUFRfEr4LJibI
LzmOuiIsFNp5xoNirHyrT3DwD3BVOEKVMtsh+x5SfnTFvOATrJ2UPurw8Y46PUd84eP0R3uk0yVz
Kt0Ajy3dnYtHc2qwnLFO3SZYhM/uEmQiOTEISpl2TG5ARjfY+/QpM3ek4LkeRbjSJyXhXMHY6m7c
X0AEdMwG+wH3n/0biH9ctBLkzC41j/Tq2qRlE7hDlcSHNJnli9QmDVgVi8NF3OrIsWR34uoHAKHm
kfNJv6WjtITYSanC0WofUnfthdlaDFomAH0OY/e1zeuEh1esFP3rGJqd47tKa8RX2dtZUwuaIw04
lFRYV3ptOsDsKSkHNkQvmwIPX8P7aOJ5mrJ6KZvOFoB1gHwmX6NzuOO2Iy7F0ADzs89SaHLBB4y0
wDZSTZZiw22p7XFi8H02Z6DOhvusdhHdmgry4Jz+XkLkVY+A2O4jBx986l/0Bj4f9k6q1Fq9w/5/
lxEplfHFpUaiJefiImWA1V9wAMFB/9ysKfSnolviqHioVUtqnZzervW4R1dqd6hMclpS623IGvVA
NrOigyZKyP9QYcpIsYSvra86Z0PGP7PBCfqrJX4IVaDfBq6i0Jc67qoy3xzfhrXjjtT2zwWRKziL
p0VA9mmfIOiXorkvLgs5dqcU1w7uq3/IdxlycUoVll510OrH8vL7wX5amSuLqdWMXJ2YSkTNXjlV
drDA0jWXCrdtsF++Y5vNtTxxxTYigQzH9E/wCcgugraaSoxpw0ZurQ+GFRYmzQT4LT1BbMGZ5Fa2
MmSK4NSTdVHsETTmpARmYPVdiySH5b5AQjZiZxXwv1pfP+5R1kNobk6wSpAeU8YFilxTyQZ6JbIT
5br4d5uoSk+CE/Wqnn00lWHBORatYnc64vDeM3W94bcQJH0xcnRBcxjjGwh8JU7LFabciRMl3pWg
3+omn/6wZ8EjIJCDALOG1fmS5C1NrN734y5az71Q9CE7gqiNKZ19P1WdMhZNs2D2qb7yGNdaB2sX
YCg6RhkPlJWWITqPntUXBGAGllqS0opnFy4pCc5ZSOFWf+uVSN0feSdKuB/X66nak5edh59oc7yZ
yoCAs5MKF2/i5/BlUs5KUb/Dd/MrM84l0MEsQ6tloEGsMuEj2AYXi0yR3z7Zv6l2I5uIfbGpHkIw
/GJHDH6Yjhv8gWOAQc36tV35G32IhzqvGp0fW2IKW6IWtWujtW4oixlMM9whPzsPl7NsLB35LA8R
/9zE9UP22vIc54+d7h3Zn5bIqqMncQF5pbSw0S3NqRHe4S1HLR9yQGO1+mW9eaeCUDCoBSz3iHBY
Pc8bHzUIGEkLmKzqsc3N/4+2p7T4qXLW6rdCZeFm11USzz4GwLcuOpn6MOz5wrdBlS8tdRTbqxzr
9ox3Bz5JlxSZSOh9B1KMLjyHTADTLyGaq8lUYoxnxyOPGVvujPy98OhIoyJ86/FeWxm84odbo1U/
di1zmEXVAjWfJf6dM1tJJ+0+dgAZWmTmARniqOHsEyj/ah/qcuGFxUDUxwPKDGa8udZ6t7WrAutT
Wstx9op/7RT/v5Sjjwj+aK7YmB6JYzbq79EqGdviHM+NTAbE0vLbFvG/zPEYl5uckG/0N74JcpuU
spQR0R6x+Y1KQRFBv7K1HLZbSu6teZffg6QYM3VyNyQ+v9UMYveNbAdTJC20YtmjxhfICk+McaRv
bFFSDeNQAAVh84FP5+47nxs2BsoMCfZGqypZ0iOqNy0x6KnGk3EbDjLwuFUVQAp50YkfIGMuPAKZ
gxMsFaLLWERfMi9FdAfjSKEi7nALFBkczeteOQDZu+e8QGoBozYRIQ5YqbAWZCSDFxSn1Jc8Ahof
DnO2UWF2MtsqEKP0oyUmQ1Ywwfcqxps0jSa5BgU0XFUEKIuVr+5VzmR0yGvWbEhwG4sm81vPFbmJ
iPP7rkmtKzbe0EUJ6noF3ukTqYLuIU/zIXlAZXi4XdyzGbQVLKUS1gy1z9Op+7qogpF9WdDRPIH/
yXJUZzXBGKU+hSoCh2qDiklS36B/uiF+QcIvScKYM+ddt6Pa+LDu7ddY9fHw9aE5wSJLhOzgc+QB
WXaJB5q2HObA7tFBq4OJNBhshJnsBZoRKrzRiRxfaCV0apvpye6Z7wWx7zHva3qXMQ2QP2bUIpjS
KrwJJNvvwSz/cbOX3QjxWKrkQxiKJddCOZWrZ/2wTYGta4ik2YjCTljiIxtQ9Y9B+FBgCyl7PPGc
UiDJJChl6y6IUi/9zJxfAMR2aImVMaFS5GqDVlUK/KBtFfWGNlhuyUo9Uyr7e+AjaWCDgbXJuyNS
T6w921HD4gNi5YN+IfsxRTzKp0k89kYDRtBdege9BHkm3Nj9XlAaj4dFcP847sLK3xn8kY+cUY/d
eY046obn71/ue83eR1xCTvPO/SRE7V8B1EPHKwPpnyQPPsysPzmE174n/eTzcQPixCXvaP3NoU16
WUqC2Kaulk5w2PDJLlpv3XR1QyXewfIthqiCjK/6NknYYvBAUUU9PlszK+3G0NiFMO1A1/3Tm6fe
4/DHUkY9ve/n9FsCVXJcKN1RbXbSaCzgoBC+SWWxhbMQgyy96FTjn0JTZA7/tceEPgXDshc4MNNS
4l2wZnl0HlmNa5tNNU+B8nJH6Aag2xa0oBdPyHphMszq5u3fXxkWDWVX9Kb5igaMjWHW4VNFfV9/
BaauY2jngDDYU5v4HKs6SPvpS6JpKWOWRO72uFe7O/BPXqOvRb1lTNxXikVkbHnij46PyAspGXXP
51hic9KTjkhNOpvaNtc4xGzOp1SO+w4h7mJF5Q+4kqPQT4k/gjwlYExLSV3T3nM7Ho/NqZqKJ9dV
K8NS/Dg6HF0OzbVNcTmRpyM+P1o9j6S9bXbGkbvp21W1AKf84m64f1tq/DCTcgObRpyqKlImVlX9
Cx44f04ZiOf+PCa2oxYgavxUbqKwx8n/qZAuDVGF7VAMTUZv7NLzWeItyxalmgGyFbIr/TTWDz9j
dkc3gkWyOusJye1lToK4c7y98J9/DcsVjOGuia0sHkD5DKgZ0P9jRiIkTPeuOd6mlL46pC+1vwbm
ihx43UkVkg2UfGDiK4BesjV+ZaOxw67R0mxxgZI11uEBSGtYIxcl9lUPlCEkVqQOr2igxwnQYHmr
99RLjTVzSCzqzf0DoFIAaCb4X7B33hDF+07jsQEQ0hYFQHFZX+Rbyj9XD86BSTcAVyrB0ZNUh1zA
87c1Hrlq+XOwPluKK3BATTj+0OWpXVi7xdIQywm+27hAEkaXRu/IMJxgZdvaPwyFgjxn4KwA6XNC
ZVh3xjMaA0PshR0KhKPAIw9evtb7haoVCj3i7fTLgKmBBEce6YQZjMf0X8q3SYw5K+vO4FrAny2i
lGfivihAV74QTaNDQEMwSVyaBJoeeUjv1RtVsMoHpOGBDqX4F6A9wy3RfLqhnZxRKVcRk7g8Tdpa
/HjmPorEjanuaai3kJxVPeZpmhCNhrlFqt97ohjkG+Y0nmbWmRFV6FloNPxuFi8NkPOMT+EQrx1m
R5oFWhacjp/yCZKJDDMdlgHP+gSnu0jSGLDUTArjtjIJEciQb/n+R2i6UIHb3YqIWuZyTiGVM3JQ
UVtp8Ksg7r66wrR0FdcxYGWXarjvysyrp/NEWm9CURz1+ZGAlT3eZtWF5mxU2PcuxeIFWklXdnPE
4rdGvuymdskNoC6kvldg+7FKT/nD8yDoVeepVBxM30jwluK6OBsA8dX8me2L/4ck1V7M9+0THZj6
UzQLezSli3o//iV9ZyO8qlyelknRcif4dp8L19XboSE6auWgPmOmV4zIM6+zvBFgNtUORXA9/cUZ
fvNbm+wEsRMwJIRP0RaDdZ6aXlzyyX3VOOMCJjbGkIoQf+ODLW6kdsjqbitmJkFjFYe04xFxN48I
JkhFC2JSOq3vk0Gs6PnKctehlCkChxmbCaouC+xpbQ4gOKSJ62D9w4Sk1ut/57Mi4NHXWB/Z4d68
Mdw8s6WmeYCaJpe62DpW684FKUT0mYmxuw1S1R3+TsUDM0U/RzhlrgtbS45u8eLXhodE4O+ksx0E
6zUwoFB41FG5sxbGq06+vYK4NhlvtrPLlY4jI5tBSCiAMvLsv+vtAFsrhMyDwyhnyDS1Ro0H8T6s
7U16ivWKJm+z/jor8W9wXgn9/ny50SS14SI1n0UYivKOSGEqCmjQKACBnHzw/zXi/7YycIMGw+Go
TTmekNbcQWK8T3DMotCqrwOFBXyBUuXRgtdYzkAg4GW9v3erK1W1Ap/bcYEAO23nzGuKSydPVkmp
alu/ZCKxaFkw2Ey36MiS2uY3uSDQBkwAYZeld9ESzKTbMxRvEHl5qyTsEBrGXPIR2NXiHPx44tHn
uhJHwu4H6fcrIg8a9S5usc14S/IZyAAY3sM0NaAAetxC3RDwaMR9D/5wPJIPYaYxH0GTuSv5LA5x
S8Ziej1dNzgnvJ/SWNL7KYqgSWuqjD1lpBcu87t0om4+miIfteRZAN/Hh+HM5EdvVhIv9QB8OCh3
LE1oZCWNtyqSgVFx2f+P4PFNLd8SPGFcS8IHZfhht5zYtGQDFKTYzKxukWwdbaznIpNo8QTGpRDx
MRTKPoOuMNS7TTrmiJyPWH3jqJpQ3Z/p/Eb4D/i9A1+75mCXRIJjSSUC44MQZv10r752BSU/GQvi
qOwBQe08+lCT/go2GlQlDpmY4S1nvzFVnfF8eNyDl3z7Nszcq57xKTdEkGgbVDPfpHm+qElOh0x6
8xD02WjH0diAwacN4jgdwb8fgGu4/CICqAq4hU9/IYe9d+O5z4EZzb+y/hAD78aooNzHrT7HfK9B
rhI/olBZWDoe3VzftdegQsx1/Xvg9RSH/2dxhMv1wttRAZ5decHtU6wO0dysGbe7l7tgGIDvFyri
eVY4e4dDKDm1gzZB193EOtN4yNxEZgK8sYdJPwrxWZloCMaUFEAw+TuRzBgqP94vXDqbO5Pg5buD
L5nm3SJU7rZXHstFvalJaxHjggtTg/cWv7OqcA0hSGyWSLF+t6wB5bpvdBwqyJwzlztTeR8waLVb
P88UIkvci3nSbCitO7bN1CxrEtkg0E7eqOpPAjRk1nw5rweKihgr+L9R/axqkyhwUH1bg5M1KuK4
E4G45T1LUBvAWnSTmnbe61mCFbOErrMriASF7Ank1y9eC3gGoVdvTYGn227EC7i6ZGFmItFI1E0i
zC8EIzFg95l6ctRpmET+DWPgWoABL74zJXsudDL2KwwWngbPfCQf/LvWY772NN+RDLzAtNP/7DYv
9UkVaupkycW7zUQKVxoKv5zYKB9KaCod0DzQ9lumy0RDpCsE/J/uO16lZwG5nvkGSxRoZ6pY2XIu
789CvQaHpaN4Yg80ufa5PNBY8Y8Ne+eld0YqHHHny2A34f4FIV3WGIjCOrfOT4dKluZ4rUlAtMtJ
NEUTT0ZLjjY90U7DHJTTjlch84AidZkaLMUnETV00A+Ltfny5JTrXi2/9HpoCI1qGn8sGrk/L1+S
YjpDMFASlFzVqdCyW6+k+OH14sek6Bp+LXlKpE7GN9GSahHaV+HFt9HizrP+MNWjuwL0boOKslUM
umafXi3Mjs66rJpnD1ITaNZFZKmiEbtRjj0YUXemojyRcmcgVWCxlQAQjRVRmAmu+wAqLkCf/2lI
QNfhTmLo1gHyrKeRqrh+6wqcsnQ5WiNfNhv+ANloFNmhm31k497Zyv7afeT0nFDbJflvJuQg6woA
oO7FynUCU/GFHKU3cr3ArxEdBPiuX+7Aj0skPULGlQrW1dTGXkqnWEzXbcwKAaZGQfMdexmbABgp
tzUPwNHWAhf7aizHoWw6dEc248E1fXwrOKX19uIe3KduoKCO0TW+jqOUrkGBmcUUgQuXQ7J5VOPk
+pxGFoIDAmCje6d29DPl1+tp9krPJIz9x2vhR+Kiaqj35UGsQmMIHqndz6v9GPORvRW50zlUCvzI
2aSJO7lW6RS/wCcRzeoIlMpSxEPS832R2UFW0k4JrZ/GLu2pakGVAdEoDoKr0PAiEQoE8akc+SF/
sV204z/PYC6KtFMVxrI+YF+omx9htOEYt84Q92fbNvhGEmuJzkxVhqhIklRzjWGRurpgEU7x8c6+
Kbg9er+B2+cff9oshKKmgDhntqL3Ev3L6ePdJ/6sXDI1tjKKnDr1L7r2gEGqUET71yAEl40rTXtM
tZUoOUZsrWWHg0oS05Gwggkgt6FTK/iz0fy4Df7rqmPl8CPvtEVSrCDbHczbns7SmFVkzIipYSFN
iEYnvpmjCXPPWSMetpQUpid7naO9dhqUpPn21tIA0eGcATZX1fiaQP5CQjTQ+t9DL2Q/onsuz7R2
eRoLvdhMppMXTj/oFHIP15TGJhRe+b1dz9HYBCwEqIEegNAfToS09K05MeN+GuyRnD/N4fy7S3fy
zwinDBpr/1Y4H4nAm6eqtzAEhVv8NfKRJqqDrw4xzUqYqMrWIAN9wlJOj0pM1XqCyG7ubYhqW5Ky
rCHMUZtgdHHgxhsflJMNCuVsXJZk77CmqoMbijqFb+DEsTS7vkp4wZmDPW2MdSzq9i/pdpgKG+lK
GTSVDYSe/v/l7iDCKRp2Zv8t14MliGvohE0LwAauXR1yXfIbRx2av1YjKEYtDBIPQdhdRqqglrZC
+RzqEvXoPzEAH2wl481OowrP4XsImMoy+kfspK1GMmG1lvuL53QB5SxZ/nFFBOg41vv7a9lcd+xF
JehFNMsRNE+lVh9IXaHSwlB0FTn6XLOjwfBUO4RrK2qkDK+ZBuTmHABpdH4enOwSaMq8NgyhMi+N
2ugIFDnbZ1W4oXtA0hpw27JgXoo266C8PMcQZF6MgiB6H/IO/tzW1JeysbUT1N3qwOF1/+LvLE4G
tPBYioId2BEg9tXngdoZO4l1I0rxfflCSfvfpOtbz+82/U6He5ClnXkGvT6jC6su36Sp8wmOInyb
gTO3i09nWAS10DMc2wFKkcd/QWaOPrJaAj8UTjvFECPQ26beLw5tiWLAiaki/rgOaM3G2B38o47c
Adifw8rQdw9sB1EZHG+fI3s5i2knmr/qMWK4D1DHN9Vx4Y2xtHxEp71Hac/ei1F+3cR6GIaHGf0o
mUQImeWi4VhP+HWefG7q9nH3hI3PnaKbQ0wdZPFbCOiF449eO3iGzO2RVLW2m8It2ynPX7yB+GlB
e17GhPa3udQ/5Gj9vPYSSHu0FoTzEkQ9zO71R6YDKX8uufzZHI9fIvqEMezQxuImuUTzH17J8yf/
VQo0mYSVIvxYGUqn9bSjijEEN2BEScvcm+ibEYaS5zuV9hUpagKHlzGMfhxIOvgAQgSLoTfRyF1M
XvrV/deOCiHbezcV4gzyJzuJgdM1hBF4oMerOKeJx9O15rBcizlbEEfl64nJs/ba/5dwiWXvFZPa
w84ltPG3zFXEX1Hu5AYNBRRBhTXvKRRrLWZV0n/qYo5TyXpBC61aDo8XHPalucRJiI5Q0UHCU9k/
JJRpjyQLi0m5tAJl+HOTnom8Sfab6o+/3zQb+38BEnUNzmsjLPVAI+YV53XLc3T5QS5+mD1IonA6
3IWlddp9Xj1ZFKGI6ZibqaSlPIhoEZwU6Vx8g5WPQisYvgO7oMevy0vkHQRj0BBSosPoLnBF4OAa
Tm7ZTrLthAml3h0oPn050aUOqWJ/oX6bn0mYGf01YinAg4pj85yknSW7o/AdQkiwzBmQxz0mlCnS
0b8JCGXss3TVvHAApb3cRqTP0f4hg4l5sR9AXGH0dbN3cr7ff51phl3M5F+nF2ms/OE9F4KuIpJ+
rKbJHmjlmNI+8zL9Prd/OO9QP/FNNIS/J24nZTgICHfXSB2ICvQz8Azes6OOJvaI70siVmDeAM7E
wsoEx4jLRWOtqpN0vVeK8wQ2LhS0+R9iDbPnBFTC1vE0XDbmyzTU0mfeQQZuQs1eZToB/vGMptHb
stN02suwfNr1nWtni0NjdAu7ed3lNeayHJjLTXv6BRfo5a6QSdphk+Kooxp8mXJqUg6y1QLj6edc
JZsFUIPz4CLIGg41axjYIrJBkcTdS1vQ/NELN7AEXsv0jfkzX1YAEdRYesMG71y5TUKqx3joAhHp
qHRExG2VMzQfm488h32zewLk9T4m6QzGiI9jXxeX2nHOuyg0ufavy4ueclgqqDjk8tlNzPa9QRBY
P2UYwmu2aImCJuYcNKGObCj1m1U6FrgwzZApZQfmLYKxCOsgLiXaZXvonsPLFvHhMCLsZE5a52zj
vCoAbGObliMxxBFZEgHzLLg2MpCDf3cg5dpucKl4vywvib0MLHEB+t2kv7ke4dsNhNJX87Bf9zec
A5xIn/Z9DIolU8cIc55Cy9MixliER2YrXArhwcjSlgbQGtl2/SCcXfNZpH/uOdw9qmYsY/W7qpui
FRCUJXDPNS0NUN2Fgn6WZMF/41g2hX+HWE1UMsYLU3fwLxiA7QPdIDd6mL5XVx1Q4JpisWNZRYjX
NeWCqzpDnDkNpq8BpODqtGOkSyvwzIUhzNr5SbGciBlsEjas0VYjTK2RlJF9XA6HYCW2ZvSYfGe6
wpYhvp8eY2nSV3O15WX3aYNz6ivQNIJKYFGNudPyAx7V+HCvVK/zCqNz8I/Pf+QqMd9Wlh1ZwLFD
VYh9RnVZPWpEvJ9A0/ZM63B2SPWe0Uu0a0N9qrymNgbgsyhCF8cSJG5i34XsWdOFEVjdhoiQYDzV
6fj5CxMo1zHC+2J70WEHBxnaKMbg8QS03G9qWfYq8/u+pyA9E6JUjjrn4jGl315yzMRsIlkx7BvP
MLQsnUfV9/yJBH0vweH763P3mgh72gVK2MsWzQy72/jgXHZEaT7Q29fFT5jjpJYzqOIuIAJx6lHs
ZwZ5GDDg4wh4ThZsameDQ3J6B9fbIhb6ctH/otSCqFtt+Zu2gcJMVZlTA9px8fa4KbVUpVJEnEhZ
L5CJiVbFRRM5E80KOuodKwGh30a39psKHgnvWOrIzPILVFk9bwgBjpo8Oimh7630B7nrbhNvA8xS
e60U0j7A74V0a8pgN+M6AjCeEYR1XhnYK2Nf0JooimbpvNQMYajqV+Kt2OSFiPO6prNdmaY9jMmp
cIlpeJiZD0O9kUC79YFbR+DltfBv57UGVOrZw/b235Ig5V3sU/0NToc1Gr88uxJvRRBSFbONQz1q
tDdxwalpYWfQTgb1Bro0E+5MbcEIcm+hyUzzySzlqYszyWdEnprmeaVgAFLUWGj2y3VYyZdn6SZO
g4HQ79L+CEOAvB6cTJik/v9au6tO+65/F0uxZEku3KXIETJZnNrl3DYV4H3h2LjVXzxSPG+JXVLB
33ViQklqL75MsPafm7+tgEwLIrvRXWEQXQFSlh3IC41/2aIoT2Gsy8EWQ5sp6LF3B1QoP7yuj6pj
jzFZR3fs/vxQ0OXQsRfB7G0uGilLnfkkdeX/h4gqKGnxt3Nda54r6R6E5UUrt0ZG8BXBk2sl/PI1
Afj40GBHWeSIf6uaJ7F1T2tfNcdQO38+Jhxt8C0O79nP3P/29wmwdq5OSCqZNPNOwSb7vpRtSGH4
b/LBjKaHsz70ssH0XktCwBaeGq9rLV5/bE+stCL14XdPPQQHcr6DYqXjI+kv3lPcDHViB/A51vbG
ngMhXEXoxLxAMuwKxNG05hQFUhX8jsxvl0BZuQDNiyxSg3QUCpEnrUoz1JLxIa7wpRej1fvGXBmS
ZyZeYeQo++LAgFwCiimrlV5ti9j3wQe/CwIB4RdEE7ir7Jd+W2kLfKmHyr25fgEoIZ6wONEHQiDR
DLJkEOi2xAbnpiO4HHFtd3Kun49Tt6RVfZ2PG/0VfdKGfECpelyYq5hqTCHZwbdQYHJ54eSHsKWF
OgcuEZzF+sfElLQIY02SuCfBGVTX2OQJkbrWfmFRstC2dTvmp9fNlRJLerObtS7tfCqFK1RFeDD5
JFIRmEvo+WyNob7EVXOpcIpqwFophNqA4xUVA+XUevY4qOGh87qihA+5V0j8vEOnU9ogBHWWeLmK
nKYALp2Ir6N+ABFesbR0XLRy4zv74KegYKuaYIeE+XSWzU1L5u1FlPqpNvkXXgS4hipOyjeXgx5u
TL8XPQTBoJTQ6WTyuB6ghfACz8/v4NFm+Secagb0nRIMT/lunKsE9iLU+MnKn6CfJy/OwINn8LmQ
TQyVSMTTZN3nBcG4t+Tz4jUvHPISbdpvg32x3Xgqqj4HopRC/YzamVAztVp+EE97EkdkoTGkzDH5
O1yoFf7f3LVfg+WL+ZOha2XLqOJ5BPUeaszEwYu+GjL10f5ZID4jrz5/SqyKZcESLxQk12JaUTCJ
GTs2X30he1vn8lkewMUHQlsyw6+gEIUyYm5ioHoURM2nARxKbW6YKTump2oH1pOQy+kSzXyWwOHw
EMzVzvYROtpfqfw7CCBLgjxMh7Q6Qd+x3cAwOLCM0eH5+Iqynj44wm7HyU/DSAJ3ytllEiUH5Rxe
KKu6fvwCKoAS3IutJ/xX70frkUBUx+C1W8O25c7bjvs/j/G2jK1Ak3SYVgQ5Pml0aCKMxUMU1DYA
l5a7TsXaz5kyqkXnDmc+Qe5VRmYHs2DDrAutX10FivL4qeW3IZZ7BrRgbX/XgRFbPWFUr+bizuUI
5SEFsQtc50nWadZj3s15msjRfxOLg0+ObK6W+1uSDz6liTmc3zd9NlBDqhWJOtqmotWM4BRVJuUk
j3GUQ1DXq8iSIG8RRiQQa4lVElslhr3QFkRUhHOWpDtN1iwSQrh+Ie5TCrDD6bVAciQZVnEl2SXK
d6LDDOha7POke6PM8Twby+AVcWJDJZyqtRu/MEGmyFdfXeDTReRTYck/Z7rp21b2/9RAW0iA1fq4
YhJWLlfgPN/53Q73bskpWnJvYNhk+4W8Nit8OpNp/NZJAiwx4qINJ03vbbMVI9pxjtX4/QtgI+YC
zZvb/jXF7XSKFV5XT8JDSwRZ2PAaWnJoeFFC/rxPaOcjTQtdCPCW/amd265Q9u/47qnQfOxm+3d+
OWBvuyVZcZP8NT9zUrgZFp3IQVvywBqCl48KOdX1DW/7Sl0HJsAWOISuMd0MoQgN6Gwhpe2VWwcd
L6LbZLz7muTVgYQL06B51yFKxLJfOkUmOlJdv3wfobFYtqVPuTmnV67WlgaO+ekDydtEtzKa/wFE
oG1xkCLs24rBtam/Clk4AicHFwUgNdkBn1qvIXRP7HpggCTWO8FhesZbyKeOlYoBoPztLyzXG3iX
zJgMjyde7rkudVNa3m7aoKAX4i8P6m4Sm+DRus9PWTA6mHn7mj1P7lbMqrEflH4kxoLzbhuD3rRc
LuvWkAHA6GF9tEMjv7gn7j52WHl4meirn1WIGHEakbnbRIGDr7+LpSw9pNdbON86jDoJ5wnPmA/Y
2/6zBooju9SGTWyXdha1xSzG66Zci2OOEKd+9AoPxEd9Sf9VPR2xMznQXhPgBYZajoKnwKyTAmIs
rQKwarIXe67pIFyCdIC8HZPReHAhnyHSJJnaTN9uwxTJ608U9ktl1WipXFCHpp4tHfNnOCuaY5kk
ijyqi3nxsUeuAiq2/eSnxlopueukaMvxHcHrnID5PfI0VxsgALuk/TUDbCvTQXbjEy21/0AuA5lj
1qDwaa0V8AkXSPcMlpYykCLWrZZUaLJ10kKFCMI1xDgzBVFcZKJ71OOAgRwfC5xsAwlCcHsVrugO
WL3XRrEyJN7ywAUL6dK9goEPAawjy84ndBuBv0sBg9TI7Q8MiPwVnfHQg6UfhqNhvoTMxjjxAjP+
skoegqTxoYa0G7MsBGj501a4pJn18UnJ5R3Be5sELcXD6gqgsK6s2h5/tbd1EecLmHEddwKdNs5S
aEuNZ5gxApZarWX3PO6Qdcq2EAQvAL9JbaCbtuVPU/oKOUU7h+zJuKCRSLr7p9PMYwl55v9wywla
Y3+Lf2pl8C2tQmyHB/QN39+RnBMksRh3R77lTSI0x60ENDmGDhiDcX8DpiSyFdKtpF8i7KwQwZFB
6W7Te7lHvs/yGlzIwcr6OcO5vxUCt+Yf8C87q/p6Ism8IQDtI22Kik3R0j33ypjuQhnBkPB8qNjl
ZbtHx/+Nxs0/McIzjbky+JU5jnt9EMlqcqvAjWWUToz/JfvfF3PRt4Nul1OzEzku8/Er3zdus22a
saqyyFJN1kJ0ghR2S15nkuFuuLXJgcf7GHNMzqynDtxrntI3Ayehn58zhxSPV+EnvkCPW7YME4Nz
owxlOJhoRuJsTBtVr9XVIM0Ftd7a7khAHAZzdczU5OL6ZleoJk4DrIEIxFAWkH4UaPEGBxWpusKn
NMJqP0TcmMdiPs0KsZem9DYZpBhIrrXPADc6WtjFVUs4KkWZ3QanuJm3ZtYgfO5tFO6YjPdXhdMF
opkRdjsKg1F2lGfJ4vaAUZTH1ryyBJZWhTK4Q2Zr6YhoL+5MB/VHzcoYZjeLaTrwdcnVgp424N+y
UyhX6JNZBqLmUuQCPYZ6vPp9EFCIEbaQkRIfZ9Exu2WNY87GWqxp8inGIjVpduPF3svLTB/VZJ//
2ijO8YcwDrR/ReStAaDdNQChmUh/m+sjLDW2iWzZW1iDzT88WmSlWoZfSj24WvaIJTYM0Cp9UeDU
gNoXMKvU+KLKfHv8+rnzvRH9LEtqH7tDtFRSUqUD2S7i3ZJrkVIvuhyG4M6P3VtKDcqcrqU9fBcl
PAjWxNrXWDwR8WNBjpNY4sueWQ+wQ/rIlyfnHYkG+vF0+1rsevhcTj6bsTxMQLgdUXZPkdtM/SOp
207F21arrJRGY8ZKatlXueFUDZcQsIF5yiDDkNOqcNZ7f1+bazTUDRhaXXrC3yNvbm9tslFDBmC3
164uK+1XRkRgIDMIUEtz37p76NglcYIalbWvFiiWihIaOzJamk91r8Z4NcCGSMuoeAX0YQWo0q7A
hCb2wnWTC/q7TxXDfQnWc+DRTwuyth23ADQomoVklRr1Ao0ijclQIqi8s13g4V58tlyMCGsX6Nm2
8PhU5wMrSilqD+kSGhj5PuSzbOMbD3iIQTOsEeWpYBg3aW3fk+odAUDzNAVSR+HrxJGuuv992Ya/
lBLpVechkzL/krrDExDo5QhRsPJftpjRdP/3sg9VMK3yqet/HXfM4iUWp0Ynk9Xj2lJ10ucKEU90
jCxPj3aHhSmh6zK1/whWftY8jpI664eXHY1+TkaZRmegJCY7LZ2l9Zmsl2JwJ+6fZNnj2SdInjxX
Ar0CB8ie/Bb+MVYAOzEOtoZ2GN1VTuE4yDykc6YPOFxOvM6IGPGiX3s0M999Tgq5JfYlmB/jD4Wo
+lw7lDuQMkdbTI6y2+x8PpIiEJXtf8K2hvI/scQupMYsVsd1+oFLyuWp8LfEyYWSGRYX5WdNRGCQ
D67KbrhLHQrfH0M3orHM04FUWRP6Rk9VdEibLXSuqw+Fyaj8DYyMiciwFC9QQVNnQkjI1TTcjkWm
iUCVsHSaimMLnKpbwWOjzwljpz7rtBX0Re4GVJTveJJt9Cqx22H/RzThPJeOBEX5w1QeJt2WHC3K
RQiLmgS+EdGbnj8GrXA3bQei/gmSuOJd2C0LYi2+m0cZj41m/mTT6G6oSxpIoKw03y+eQWlDcgMo
7/vegeJlQrRH/+XT71gVlJH5Z5ZV8nbDhksjPRLVySnvSkLG/4lxCar/n6T9B+RMnBPx2UV/B0X2
B8egFlRrpj2xJ4cvk9GDhbNxFoo+cIYIJwIbOAxh7IonGwhkqDocB9uR3TA4mwxqDLqi6drrupXz
VNZP4Oah83Y3wCCug8lhMmrkN0UUpDLcSt+9/85QiwQXiy4F9ybriUSs30G6mgTKOz/wYaYt9zub
tH+5WBSEz059BGA+JEUXjWtz+goV0jhMTmJEUTuTWQz5fPRQuhpOoRU+qvhK963WzJhxfu2rmege
LuGQKbLccm6ePJBeQwVq/iVFuiuqQ0xwX3dkIuqlt1kqgwv+rQ8Q8eAeRtne1LrZZv6c84WVAnrl
ibeIdmKwjsoXK0GZCyt6y/wDIlcvPOWzO7Fz1xvYOJm+vDEEngOkkDByrzM9XrnJi8qreegh3YKh
+WPm3E5SPkaZa/MP0SCW3iYpOCXmHO2ulLkAFNPC1QtxlxErCF1/Dh9OFeMA6DKW7U0RxL0qg7Ei
O6Bd3ftyodpluUpx5YzON8umXXSQnge0FyIKe5sSaVywnPumbZIRuYLrKwtFP2RjN4LMMPmVCLU7
C90+7gHTvY3qi0lUDyVnpTV5HVaGrLq8kSmf9rMQqWt3qKf7QmQAMTcn2js0MtPAOT/qJI5iWWh1
9IcKm9cEB9hKKRemSP8eeGlTuBvM1BWvMbHs3FYmK9YFsXzU8c1OwMIO5oZ8DajQ+CWXpBrD1O4Z
1HX8N5WPBbnYC/GzqFQktGUanlDE2nnRTnWD0FV9ELPt2ctPvOGEVSNF10tvaf1sXTPpV8TGnbIe
Sz/3qMDxZzTVEdkf9xbu3HlzYyi6o3A9MN1Q1DC3tcMseJowRMOqlj+kZEXmkZmiTtAlrBcFOF5w
esBW3WwymNPLI3ESoO1D+c2SvEEP730uqo1XokZitK8Gmikkuh9FZe0F5Vy+NkKyPTfDr9P5ZmAk
PuAYrPi54JoyOMb3WtDXOIZm7mdscE/V/qaUtjpTEsdK/uXyMf0R1bDbdWqpqnWY7hsGkiGmIfa2
aBtu32j/Q3hkbP8YwIksXrNt6oNomDwOpOPJ8TK2qLTQBj4abN2h4NU8vvoBXHpM8evUHB7QEIzm
E5GKUr8QAz/wKk/v/yAnTqkJpurGNeBq62PL3xE3DRKvre4Ie02stHrb+8qCLgPOgpVYYpU/93NG
JNVyY0SMFkQK0JM7CewdP1IUBzEHP4K0SvlNANiYZKq7kqZHUKmeRTmnKR3trcKJ5LTcbJOJNkLX
SKtAHfJ1RD/DUrcXwaeXNoBFVS4KWQGByKUWUdI/3k7S2X4FV6s5DpdEfl3iFlxtU6JtcZa5J9uf
WfIsS2EYvAZcm3yM6J/XFf0e7wll3tcETE3eg1eY3bwP4fNchQyKrMozcIdTu9vuxc7jrVY6dWnL
FSWo5Zxs+oOflkY1qdRiODoN+BaRjwTCflz3v3yFrcmJRViXYqOrK/PU9LpTiDExXLZ+/StvGLIz
r7RHYSL8C0NTlY50nNjrM7Oco58cMBRtr5ovQWilbNy4T5GxQBwt6GFU3lvG9hzYytWb+Gf0DNby
8R0dbDOxS4AsZOXqV3UDeiE/ff3dSxxpyOgVQT6Ei21wLDg2qSIJHqr+wWaNSs3Epq2ngC6WJFWz
XacsWVsXk5I9TFcnMBK54KDdQd+w3uzESPSbnPvBDEFQAihOifhpFCyKq3kOtQHJMlM7usLpuknW
WbNhZnOrk7FvbLSOTBf9vjl/YdBp16/8gp6qshRuxo2cJtRWlWflIrXCsfl+SmPc7Gx54hU6HmGW
rquHiLhwfuk/JNV+cpW7IxtUC0744eXzsXhGqfFmijK00dU6evOdLPrk2dXd/n7stD0fuG40+EPI
fxtWc6T7/0UdlhuYTh+vvuBlM+/sxdew0EXxd6lKzBC3/v3KiP0DDwbwbNO6a44O/OqwRwcvmXak
lvGoIao1md8UI+5DQGuJPKmGJBG30UR/GiI3WA19HVBf9lliIvc9V6HqDNC0isZYGNVdXqcoCo48
/7QSazxYccAwF763jCIW5W851T/qCSA6OA54s4CD1wOn8h+/BCBw7WTRwmYREeZmO970NPZ40XU+
kWM7xMuJSuh9DfcHwD4A57HVALcnypKwaMnW3ZllMAPq4BO1mu8wN9tJv2iZUC2LNro8+7D+l5jw
Ehz5mIa2vZwng1SyJ2WNTQWCO39fKU5MWGXfYzd5vFQxiFsIgEM4AhdUKO72lZUBbhtVhR+WZRBA
2TWY2tKx68vFdDDYF4pU8ovPvZQ41PmApspbW5YWhASWrdR9ntX28pFGr8refTDKMpFcWMXYb+At
cY8o5DK13JG2UqN+K2FgXrexB/qwpLsO5ROMxzVzMOQeh8Ty8WEq7U2/06OJidhjpGOwL0cHriO6
AE5bIee/2RczESOGFZB0QrbLVhKHUEk3lrHVv4pXgb352JHbkHxLSfC/ZdVTwy5XH0A/Nc5Y4Yzc
MYx4tNLIpG26khmSdCIrL/Jg4VLx0LmjAlubhKd+SnDOv2+ZrZhvHRJysSkQSkpaqnH6KPd2V8qO
KEGft8QGqbngwi3aUADl4XE/pdb+k3HEGe5uSqAbh8UEkMOvgRKqpc+SsMzvsIGeVRokC24uHK0R
Rmf5T60PLnxEgHcL6ODop8RRGcqN1/zG3NmfcOiYNqK6gOKqD8LT+rbH6zHNvF8rvrBsHaHJ/uf+
HMWq6fKCIxH91q3EkodU9cvRaFvS3pclPOQWhvpugyAUe+hRZbLFrp/zTaf5OBxLF0MKNFXjn9q5
S6u4KgJpjSYFsTvUyVNU0bzpxMqrPBa+kyK5tyxKN+nnn0ZF01d89AFbSnEfqECPbakld6h5BUyy
apauEg1JzhXq02K1jLDP8XrNbHcwYPQUcFVEPS0OexsMGLciFNe7RIQu79KrQ2Ap74qW6rBGU1Ma
ZfiycSo/Ge+SggG8HlSo6s1RKVeAje2LkPJTleYZ+lt+UirEs0o4fBMkYtqrHrdA+AYm+Jg4ky1Z
MHcb1UqmD/NY/YBo4oVtFz3tnQr+SvhBCQR0MTtAkSwRR+3b0QI7aXXXk161E12nWhoRp+zBzfJP
/g9r646GPS9W9CYtuW26kmrEuOg1z+1lXcduiGIJUuH9ERPZ35ma1e7IXSUXl+0gdwCz3xXNarV5
va6CZR2NyxePmmtxUNzDFiydMKydo5SaoXAe/5OBnS2L+o1tjlE5izWtga5JxAu3+sLTVgKO5lDF
IKYv7z1Qnq8oqwvX3pgD5McYBOIRRchIID0Mw/rh6nHno7LSj9Qvcwi4RE6wK9NJmRahp7/pR7gV
PDV4BRbIauiyrGM6VhKP13KO37EyM2+WeLWgr2H7lyXVpm7u3QKBHPNOE7uy6j5buQaakpMeCtxT
7SXYr265smi/E56wC3T4/V7hTSFwjvWge0CsJvwu6CQ8i1Nx/KUCisyl9PNwi/1Z0f4TicmE3a45
Hm6qhRKloMSQ/IWl8dV1LCKzGCfRHxYXQQqDxCRDagzoMVVX0MmSsM18/5LxZp1JMa1riPy+Uib4
p/SLzDlhD1L+OkTc8IM5EoTo6ErO3+uMcQ0t8HzFCHNl5G/lSCFpKt4IBGzPlkcuLffw2d5AZpE1
vnkb3priEV4M5QLHGXtkvKdg/8Dr/BFjJTadbjcZGJHZ8vwFQL91H8nfGf7Nj8yM9ECit+SghPOK
wirMMxtjGI+edqQ0086BW6P92052vxb7HLr9EfsG5QcLgz2W6J/4OgKCOrmkhzo5iuuVzeu6Zjhe
E5zzF2T9auznaovGaw1Wp7I4ZqRJ8Frdtd2hWXVnalLbHCmvh55LmoZmGlDj+xUAbExrv/Ym0/PP
WmmZYHcRjg3Gjt1WTjxh8kycyPqUuWs6rJ/P7ZrMgN5XoW2NjAwPbI5greZAPo/xShz77/VBlTPF
Qf5n+hwTUp1KWx07+yq53ZursVR64Je/CffVyz9tYVF+IN0lqmeePHobDrhYT42rQKXJ4jLtd3FD
WC496brWMRiOAfYtsUI0fedaiwb3edApHygh06L4D+8Eg99SBszE5QhySXq0/zk6VNLWk3hQ33Hj
iyVkFJtGgxfGtZrltpvu3o6w5ORS3o9y58wwqKcm8KA6qLnctzZvQSk9IoO5kj8xpH7l3UCHV/ys
UTyuQGajGzoeV7JIrExJFG4dt11/cFCqDAAAmDu2p6AyrZn9ZVanjFlIa+iZIAdO0mzG1CAW8NYi
TENLL98Kr63aYaIx+GuPVV0WsZ3L3oJ80JIubhX4A7htF5++Xxy0fup9fXcyBDbsfg+2Nlwn3QeD
DPtjQsAPN2DayIVzPTzTBYl1Tb/KfP7lwdihOc37DZFe4BdtNiH1u2sHffk9WpaFTxCJ+Ghs8EsG
Em25XSVJC0aR0rjGyqouP/0MRy+bRI8VJlqd1xVuz9WxihTodHRQpBfXtxGW2+8MgAWRTxiftqGl
g8oPdqhrZYWs3IrzMdpn61w4l7pGkUktZHoTVMXc7/mofUaS//aaUGWFpJ24XEFcG1LyL8QJvjXH
r0/3jeZy7tAam0iKb5ppe5QsFUh/sqw9Op9dRn40v6T43HSc6zPC45Pjexp/j7VvQx+4oD5SqFe+
YSoEpni6RziyJ6D/H86T5sgiqwkZ8ey9TUh/9ZGN6HtYMcHqOwoWx+/2PK+EkIbcuBYWq+GN+eDs
Qz1krI8Bj0LnSNNR4v4LKi8vYzwnRTpelnvK8tBEH8gBxayWFuwT0TbZ8VypLYE3XvXSlW2Hb1lf
0iW+MYsAl5SkvBe0+o3YfyEwIouJPTcK1gAR+USx88bUrr981Gn+rTohflgio6qAT0+GryWCP98g
xZanBx9O1hq2Opv18JZLLPVEnM9Ghnpx7WWngCS3WDJndbVENHUsJqKTUzP2LnmF4AsqzQFuWqOX
B+og7gjS7rOLfhDf3y70TGjWXMmYLZljC2fPhPChbSY6oXOMZXmPa5DxaJeXKjNhpdMnYVP3HbJK
oSw1/whDJvPuxEU0/ipt2Eu1vKOYSH7/j9K4JLQCLNAGbiGOQbT6aFOgcwayGSX0A3/B92GuEz/H
sRxeubcak0dPeV/4+tLzESeB9LqeXfPlC2qLC5LGLABDmTAM0b0IBarT7qvBNuRBqmv38bQnuDFW
Eyp3SNwT1oE7Re7in1M6yqkZuStU0Fah2BBT5sXyxcZ4oe4AFUc6y6U10K8h8xuVFHq0M4aT9hcD
xMt7RicyYQXmGjh/Bkvm0MxMC4oIUuhVZ8KVGbQmG+ka7B+AswlaqSDo1svhsFs83YUdCkG8NJu3
yu5t+9F7h2IMDYItf+K6VLwvJIMQYX27yGgBY4Iuck3M9a/Neb3/VRFl6Ihh4awyR5JHRfoqegRm
eXbYUXQBvhM0hgdsIodW7ukvGylYb9whhKvNhR9/qtshx5pyVQgvyzVBlv5k5v1avaSN+XCtTiZo
Zn3doEvbl4JTv0CmY8/GTTxs/ubISqMI4yQms1+3kD2RUu/oGKhqrCbZ95r6K0Oib5x+RqxyXySh
5zBtmbkXbGupohJEQcGJtkEjLoiTC45nz9pOCelPC+Efd5RG6wkI+MYbdQ9teLgr9S+5C8cWrxmj
/I7As5E1nJ3riqr6yZfqYJVqIYEEqUKBEcQK04PbgrKckEgVyh7oem+Oe/eUqYDAdwUmJRsnKrqX
Fh73m8MOB6hPFKiqbhlDaIPe2a2lrcb9bQSJdr0fHxywZkhIQUNcQDNfkKs5O4UOv4MEu0Ziy99b
fEiAREiMWCM/3Uu5Ev91REO7OBTlfjQjjxrvVpqJUF1+48E4JsASKbJW/fYxdhezY0oNd+3EAKUU
U3FGXrOvJfS1CThskIpF2ucuIGNuh81YpBQn7Js3GfZ91/nKzsM4q08VLyngHbQNUWuGmnheL5eo
Xoy6Pey1MGBA+UulSeAfi2SqamapZ5aV/OyRYt7z3MxEcNQgjfDlsxKsFqU/7/8lmuKJLB2VF2wI
mB8242NeS9pwhosLR3EMI02RTN3DHXcAeApMgZ0jCxmPw/vMdouihXA0TYGCkMU+oy0DPtt5ZvTp
dOuIkqg/+JhuK/akHIt4H/yj6bdxw5wtJ7oB7QWi5YjfDuA2Qm5SCWCiu0gKfeH/GlZNDfwvGVtb
37UGGUKc86WWYkCecF3M0XFnYOmgyOAfA0QLW6JWycd8r1t2Rh2ek0OjxxPq6xlanJZuo2rh4bol
YtpUJljV5XyFHQwlTY47WtD3XLreJGyFVxLkk8yuPLTAIaGtmImHpfjZAC2xSv9sf6FMsOaAxm7i
yfCsIQP9BeRAYGSJOX0nsVp2ZI6vdgWpRr3lJVBOLuz6TiGL8YzjppJ0NrOc2HxsUfmzQl0MZRl3
amXpeIox9yb3ljumm9AZmhCdKrT/sTKb2qiF/fda091PrV7SwUt9n6dj6TgJ2NhCjI/HJb+Z34o/
8heeNyZC8JV3Co9KH63WAENaBT/Z30zBdiCLxIz8ivqOl774HbEqgZUahU/JKhqpjzByxlWf0vVX
NZGVt1CeG9wggAcQBDZeT0PGMagYTAZt+mbu3YLhhrkHRcwUXhizYxKqADiYzWZlBc+u+cIqaOz4
jPWrx8B68QEvrS3x80UIzQoMpMdBPbhPKexILpx42WOaegMKELyWzYhXHPr5OEAc3fxgFoCSPFP+
pWZIUALDOwIb7hkrKgUk6Ri2hmLgrHgEbZ5TruHEkOCEoMvfM3dHU8D8oxgjXK3CXNC6RhrxOTso
yIyweL8Zl1LQ0kDyHg4CGT2Y4PCgjHmJ7K9Yzew+fj+LQTXmxFisl0Zxh/S8onzMzG2y7vIZ5F3F
oe2GGA2NXDP+nkyiJqj8b5+H9zFVHN/T3qglQD8jLPA44kt3T+HlXKrdm1/o1mYCI3SlzpsLgdDT
HiLgeuQQbb9Ia7A6aIOV2OPE7sW07doPSxa13HHqFnlIbH1izn+oZaRIHaMqlnVvmqNgnAfeRy5t
/iLcDjiWN43HX55diy08UcR1g4LyGbBQAXn+qUwO7oj8yTIoLiDvaIW6PiExe4dfI/AZKV9JS5kV
49YK9gOlSUhUJjM+THR2LIu3LCgclvZgCFUZUb0W5D3qdtLp8TsZUajEwUv01DnCS/BjINC/5bzl
nfSHLkinApKz8EMHYGwDQzeeUyKGh3luO+4cypvwWQtfL9zvKZ348CRe+D9H+R+4vnMcA7zSj6+r
SObIAM2HlkerGXwJ/AGyYxeNoYe8Ffw8/bw81IcVwyxjeEc+9JBgYMBu8maCR7+im5PxRjCU6aN2
Fox9QG3eRuXx6pm7VlfHNxCEBeYFaXrSlTwIzI02KrcwSeb6HsYauH9mI4xI1GgnrmpDudqgEB4p
H5XOJ11Xxc1l3wXDJc0FMW6YoUYznhsOoq58ap7KH21Ix/UPCc6z4D00XtXaaz89cbePrZD/hrG6
T+dxyWdUwoelFOiE2/z0UzNjJvM3+iF6jwVhccdZqNmj0TsWCILOyGdxPlxlZnU22qmC+GWNixMC
EplNBiNK07HVNwKULAz3YQt1iPVKRbcsnlovvicg7RRTc0F+kQOSESRClPdkIPGwvZGB1k8xyNdv
CzuvlE7BDKJBwKYdY1k89U1waSqjrZIxC1KVQMH/xoIs1UKnBx++TlWNXYr7HrHFviX8/VMTHs6Y
KF9OdhvnKF1KUVJBXqOkwC0h+a5f5IlI0S2M5XjRoPrtZK4ELwwH7exad7ohnNZEQT0/t7djHSkR
HkEKEkp8WuTvNi58Di+h8UzSxM/qWFMmk+DkPBgDSdQBAawudPVShqaJ9ArAecSFGXcgJwfpwF05
XO4dkiN0MlRuvK9fFMPtMZirkhKfKHbEcr4hQ4GSgwK/KcMi5MU9IRA0o4CD3RD9I8QYm7YlEX5p
HkAIT0oaHZeu0lL1hJ2Krui/arFClo23+C/PJDsHsszdO0v1F4lL9FvdZ3zccklJqH517d6Gqp5w
8s51loWV1UW3syS+DjfjILs4X/r0HSKEUWQH+yLyPYTwUbGFZt/eoNIt/aotU9zG7JQgU26EfesN
YJzhJHsXoNTw2PiuQ2w0kuEiu65zHLXyZAABxq3AhprOtCiibXBtvHMoUC1opCNbKnBooqfVf0z5
BccqEfJLSyHpHERJgebZlD9CSVIgagk5J0eB1IPZlQsZtyiXEg9CAQ939m70c5mYIsC3m69TE39S
Ub3vLBQC1IQ72RymdxrcBpl9fs1oM58Ial5WkwnmlYxLzYYVcuRYrMqEC2AQu4ed+G0l2nvJbU2g
ZWwzAg6OPruhrDd7rKp4tA+U8BTce7xsQXoWZTdx4KB5Ie6L9Pm432MTBbkogVh17/Jc+FtDzMF6
y6u4DUhXiiQXRGxerlBzvSdvaLP2O+TAi4lO0K2sjTDEC6NIB2T4RvdVa/cooupAWR/Lt3zopApa
760wJGdGSy1ta66r4sv4Tf9arg+1qfacPP9iy62YF0tMAoEYC8mzoxN5+SDz47CxyyaYHKnz0TM6
roablhw15jaAx+jv5mTmiPCgKdQSN2ArCivLtUzOvgNZdx/hnfIL61Er0zo8z4I4MWIZ41vDwiiU
rN1XPvxM0Crcl/n6gDZlJPno6LEbA/iMV7bj1/a6tZxw8Y3caepikamm+C6DZosCHadl73uvwnMa
TPMaSz0o/wlBTMg96CeAcHBKMhjxQyzqoZLuR9m34uTPBGefu9Lds87vQXgcQwI01yeGkAcj3TBc
LLz8iYbIg4stPU+aGnR4bdtG0xWDCe4JXd9UzXmWtG/dynhaXMtdMEv30JwMzQYw+rva5wo4D3cn
6SgjgYAj47fTHlTcq3WABK8vDGX0+oucdkn4ELFpCUXlKRgamWSuZeW7q/6W8Js/T+neUeuJzhkQ
L70EpP4KJ81RzosU838tk2wvPF2qI8B26FRHDNxl7WLpnxC1P70ERQC+mRc/SYD1NACXI5gGNhqB
k5Y2/WGIlVi+zBsDZEbsH7AfxdOUhjXAldxV83FxVaKZUdcKIKObeCxzkAg9jxZlcQWJ8RN3vqiu
+Oqa4ysZrv3lcni8RL3KZ2bKMIcAIOdMG7QBbzZE09hTJrGLvjsdvT8rtpG4Mqec8t1fF3mXDyg8
BFng+l+qQsfgReWuE81KRukAkdbbGkGD/dmXcdO6sgTk8UXP6st4uNv7juSMHGlwi+DmHDRGfvpO
RLsfqxoUugBii1Q9WtF5Df6Awy+Kx+oxLF7lU5pV053Eo346CQJtuii6cqm5oB08n5mDMdC676XH
ZmOB2Aa8LXzBKnWgKMbyo2tLLALePx/kzUw/O4W4vaHf2tb5H5/eT2pHDjDGli9SD6DtwoKFRZnZ
fCTdwWTxh01jbWsviuHukr7cs5YQ0P5Sd4UdHfdGUfVntwqAj7O7E9EtkJpTV7x2baHn8LVByVej
u1EbauIA6CFc3Piu60Q81XJHR2xOP11tfLoKKoVXUkmpIdB31znat2FNCHuqX65NALqS3eq1Uc+A
Nn8afdLcGbiPf2/P42KvjRNmSeENuumDRLZsHAyJuVHIryagrseQx4TYdOIm6jPiNKW8gVh2qtuC
ASYat42MThufwZ0Mi8gPTp1uuzBjdc53jDRvVghhPhCBD41V4oj2VObeBkwHaGH1t6Gxhf9uMWNz
omZ86Rmrme9Bmo3brHszBmXLE5Atbeu6aoZkiAMickpUXjkx2UQnhY0MZq5sJJ4uE+oLs4ho3woC
HOBQLC2K06gU4+vWEwPWo68dmRa5t5oK5d1x/yaf3JrNFgUjgBDSPyobQiPzfrXkU8jyWbMSNEpI
5RcVlm1OVBWT/yjB/ecIdHE9r73lovrS/EoX2xRzV8+JYiPnZ8eJZ36EVnWQ+Mpq33mpcJgDkGnf
6uyU0cDSv3qxZ1DqpDofQRDZ+nqZN933CRqW/ecpaiKnyQjmomg5Q7i+LPHhouloxglYz+orwe+8
2rBARMqLK1OiznAB+2w8o8Hfl6O1nYO+us4/5i403oH09Jo2Ac7AyrsWAd+BZsMJw1zl+xcFuHCn
9g5aqUnz62xZ2g4KYG5ZNXmWUBEzYwM1ZKcBAUVpWjcWoidk19+8WXaS9XeiNLQpKUUR4jNFbAA6
bRtg6TKK/OIe4UelIVWur5u7srghiVRrmot22VA3ekzFtYhAQjWNYSUxAQpuKTBnBRhm+sAEAfqU
tDycGkGzAh8k0ajOVJMwwAFllcnJ58XrZP+NVlnbqBXwqRo0eL++TAayLzJXuyuyIoEjDL6XIdQr
JHY1LRTGAQF5zjd6GRKdU3YI8LUiWaYhBrDJ5LJDUEQNsXH9QeStT4eYAwJgeRA7nfS4UCYYfUMo
Apch6akpZkgZU2ElEdIkXjM9FIZqDQPut1coOaO+sAFAwCIy7KhAiWv8vHzFdcdazuE0d//8uqPy
NyGH6AWfoNFiYrk+72BHvoOSqjwWd4Z4zgqS4c4PBZ+HGdxhG+dXrlRlrwZBLr9GlvAStMd3UyYZ
M4omZEVurl0080Y2DcgtrcYDIyiIzzfqqvvmn224rte3dI/IrsOnF6ZfYQYYsOOE/CfEkiOEOejx
dXCI+jDqmG7Mn7geG21kFklMcsZs0u0kIC6WQsIFnW2kOoHPZ74MibRtRlTGCIqiarafgT+tV68j
rAWe1StM//sKiYfZb5N8SNAfUD3uhoC6MKAXQMEly2F89iqBrlDrt4GEiuhV+WvbibtDSZZ0Ki4W
KkkTTDmNkXLYCQaHmMm8lpsMY3R5+5lyNvjtl/vK22G7+kJq9cmZbBPn9XBu+ANt8YnADFxxwVCe
QdodjnW6PRNqEClpyMLZH+WvOKgNSnf4EydFuWpY8FuMG8RS3YdPv4dUy3zyHo4h14YeYMZtxKxk
I174kbKd4ddjDtiJ6ARJCa/pdlMzyJSCS9CtRSi4nSADIe2HTmRyB6U/7kTAJipgJvmlfoDVXO2+
aFXXfa+YfY1Otq3khxz4WplQiVLbhvBpgETQUinYCVrdzh0UYtQMSzmbmv2eNPAIGWpAJqSJ1VWQ
mhTOkLIa2od5K9DXm9cEp0Fjhppuzr2iRFgRLyodE/wutvSXhySqqBY24yEqyjSn9CoT7xzn5aly
N8me8c2WW6AUOAvDXke/rvr2tsy8HIxqTQ987cq6EEEO7qot6IDeeHxqKLBBL1bgbxdEyfE5ihQ6
W4S4gMERaKn8YzhxtQSV9h4RzB+w7XMOiVlO4rqIjV/tDzBE4xTwYyCTCEHWUHWD2CBl6kIGy+cN
uy/EnWqmyrSLQmmr745XpmsKMW5W8JSgbSoi1DVYsDMdbDyaVh1vZCd1o/W3/v6XmkGeM3pse5Wc
ADAIUiKq5ATBD7/lZP1uQGgg5QQbb9JBlwPlbLwC33Cq1F1O7zcoeNGVvI8oH/kJnh+yVWsjtfkC
nf4ZojotzOCAtuStOqAedUgD3JdhxwSXwTXfK3ebD2uM1CJ0fOi9TqRkfKv4kGXSsTjSCiAp9edb
YpIEPLzoPZKHQL0uYT0V/s3TI+FwACD3xRbJb6iqNvXYgbjJlunLyafOiBIN+ookVHgYV3qumRDm
F98qpqEsY7Qler8w2BcxbFpkjZ6ZlOgsX972qGAlgYx172SgeRGeWg/R5cznsFT5RBbAAvkfCXFR
4F5MwR+bb8cUrygC+irasI+CGRdPH7kN1vZxI+jwA6Hbwi4hjhcVTqxVrTVcfowG7wz8YFmWP6Is
nTKPbywEYg9SBjgPIh3Vl+yXVfsJgV32DssGp8KudD5YLsRYmnk5ZrQvytywNKXBhUtnuTMNoIg7
f135ey5Wz4Vyq1IXjkyjjT535LTyQnbPO+FitKBjGjqvTQZb1Kqvpzru9HP8i1yUus2Uidcs6ALF
lMityhZ27AiR+10xfTa8VOssDjPGVlsRSnRozEC5xQigBAoSzrpKY+ryKeahdPse1TOZEeh3ZhaG
dJnEDzKJnSDqbg4KmKPbsl218hpd/jmICrGMv4K7VOXBLq9nSx1NDKfu+JhD1nFcbTRjNDj3fwxI
mCTUYf0XyUG9iQK0V7XSOC47M+MHc2ZVSQ4T0RSi0HlmykjTZ3Rtznd/2sB3orEoApIxVeLl2X8W
ebgIHXGmNlJFwj8ceYqbbVozi9elgYCnUzvocFnTdpMNt766tw96HVrU4TFPZ1zYxaxdyRpjoCnr
7GrVeK8k1hIQO5ZwDQmSuS/HPAc+H4kret5Fd7P9O1lrxRy0L51ri+MNhnw4NTDm2VQ37aT0kXyZ
sU2WDPZYQqwq5jq1EbFCrBkdKeLY+tIXKcLaagdVTNYxK1j/HE1wBAVvgjx7J7/hrEDcmisE38D6
+mttnTZwQT0QRFpNolY6DxIhWJTbagzR56uRk1ww2GYdNAB4ro3KyGpHs9p4ftw5rXoFR2GHUywt
YLhsafqnb/Ct6Ka0JBe5IqTcgKELhWrS2alaXg7oo8lSyKz3MMchUbM5jqlBg39FnFUaUvY4vSha
YZJZ/ro003Wx7akWTm9aXo6E7dYLDYJypP3ob15bkwsxT2wT9GbyzhjWANkPCFP7Iuq2/J5W2TRR
Qhtj+uvxK6/JODhH4WJV6lMOHga7iMDNGjepQvTKPC1k/PW7E6BVTndGJf73VSZ+08a6WBzSlErj
SDOaq62AGiOqZgEZoIk2xfWFEmTOQ3hTRfSWh4hPnOz4RXSLMInqQfgoVCCxIDS/ecuJcS1JuZVm
FyWkjui43WYhsLCDzpnjPXo767lZ+95fZPzzhUu9+F7tIntU9wz+rjF5l1zKWzghx8fZmeaEvbbL
jaFEFc8z5J6oH7CwhKyk2sR0hJvdrm2tJCLPodcC5mIjhQ5Tn1oD8NqzKvva2rLSE1zGaL1uUIB7
psJqfgOkRVmHEuBUzcz7KihIK4rQHje8o/Ik5T/LbxiNkOAV5lPP3Bd7Qka/lHVb/qlSvp/V80wb
+gep76SKy54dzUxO/cJUuWIHXGZnwUKXn6IO4lBp3+bEnR2rSrbBSIMBEOH6vaq4tq9rq0MmIIZx
Xsbut/6Y38fMp0Fuozg7BpBAyFVK/GIWSbdarvINpAU4FAnsb4eGnVwHp8WOBrFm1qFD9jg0E0yK
duaXSDBf1Ehi7ngOPBlmO5lMsJ6q9Hds2sHbJx+zD6yN9/+2ufjjavJQ5qO0ST7N3BWhetwB9FPP
PUwxfjkv654CVTQiJT93zk9MoqJIGd1aJiiCsop3Q4xffvlLnCLKGP4qrCiX+W3JnpX6WJwcJKYU
l5ZOFF5q3GfyZ35DvWJjd8acCmEVnqGgM+zQlrq0ewJ0ri8UuNehHbYIp1lO2ItabU/qLnCrZRG0
defYodmTwPXjPPOpsVbyuhKM8LYaKsgeJhsrzPE8wk/o/QobGYC+N4DxWUjjymtERbREJnCrHB8u
nfBbPicDPn+hq2McAHrhuoY7/7c901oillDpGJ9eNQxBlcMZdiCC16LsMhf3s7PuD+7jX3z/11mh
yTtSFhz976YLz8ea9gEVmCHPmoiirHR+r48cGBk6z8j0PtYqJGVTYHxYhmqQ8EubcVY18XPGcW+k
WR2bv7L49XrEoC4KBN/943589ZRK5886bTPV1Gf0zUmI+6AOUGNCsjASwEgI2tJVn6BCUh3QUX9b
jAE3zCsye2t2JBhAcGX6lrRfWHTkfKrHvDRW/UE5cXbvVMwyO4IJkA5gpx2HqpqTAoAyOUoWSVOw
732k8r/ExjGqgeaTJcggRcKt4MIy+M8/bGJaDGPRE+uxfZEFL94ckx+eEnwfTWdY4lDzJafoBXU7
xYNDd/j+J7XM9o9DAgrcsqySPPYEj5Qol/9eJ/MGTMQJ+huID5n8BIVDPZnzZ0K7K7AdfAj63FLt
dShXbgj56Hb2dZZDqfNK4fF0OqEgUl8sF/Ycg2pj9afHKyjaX4nvOCe5PjoUU77ZSzDL0/7qGJ2b
lLGsmp1jDe0tVljmYogVhHzbYcW3iWOMbnxoTWyx3HrQh7IXRSS6QS3/5NO5aBftNGhksdCzyZCK
ZBTd70pepjWDy6XxAl0Npbul5326nNap39WTKchRgFwnLFFlFKvzzxoLLRgSxZc/S6IDUvv6NFm8
vNhRkpKQeHUldL95dL3wQ0C6lk4wQ2+6doN3Lyp1mLJ7Lw4GGj+y1uGGnGlm5ZFJJS90zh2PwH7m
j78Majs31CLF2FUqAwiuUxlsXwQmGz+tZOmqYJVhBg8ayNaN39Z5HJxw3CUe50aFuAS4xyHRvFWO
SI/8sEYwRj8sVD0Ov9uwQ9egmNlt9M7d31FZKUc9MrRzbKVmVrYWljAma6+YQB76y13NrkmuXWIy
mwgYbPpgBopao9BSIJk5Sr+bCjM8qyzAZH9mxXnqTOsyP7dGDx6LUO9zPAUI7gIV4FUXh3SHu9uD
g64fSn9lblijTXZkvX5joQjuvhQ01xQ6e9bi+dIm7R2mCioC9ptYNrjU/2Noy/CuI7t3x8uTtI7A
ECb8/51NiYtmNs42ce+Q32V2C7lsiq/V5trsN96QoFckeG/k5c97CjzWJ+eP/1NXFlgtMOf4zKCK
sa8wnbPQbBG/LTawC1d11EyXVfB3jfxccw4tLGeYKqmIYYP244+3byZBF2G1Kyk3M0zxuzAvpLiD
g+D2uHYDgP++eYJFCLG2blb0f2mQ8mvJO8oKgdC++3knqX/72iKwccCAYbKVz+a7JcgQpacqb7M/
HuexMHpMFqVxsj6GtnVk9aZa1ZWE9SCg+QwFb/ybjx0COT6nmmWY14Kzk9G7AZmQm4ocDIpfg2TE
FgHbfe4PuHbgS54J5E3lceT59ivS3nsDFa/87T0WgnAuy0iRN+BFhysG9LZZlu/4ff1C6xWWXXp7
bmoi58CUU3mPpAVkw3OpRsWis5w18Pu6VfTLF2AlNd17hVIHU5E7UwqanK56DS10hLCUG2uJj7I3
RoiWVUahHNW/ESGMv6MumSUSi9Zd+bbcoJJW2HcXr9xZP4xnaUwTV3gWJofQYzNx5IkWxBbEMDPC
/VMyPFNCkPuRw39OXpoxp+H2XmN0HLpw6lRJvdpRNAtFpoMNUxwAY0ZNMR6g5kt1BWjzCfABk8WK
KFhrmGR9NvjPxrcq0KthbTIjbzc9RKSSuNGekuKhiGTDY82JwykF7euqKJuVyBY4Ixd25EwVqV//
b3a6rZAXjXQTq33jAgi5Oh6MtP2aPx2npn0hDMbtVv2CbLmFI3z5GoeRLWTOnpfSfsGmrWk/UuPD
GNJOF3G5AXtEBHM5TLI3BxoTQ5NKAcxF1w0Hz3O+8/gSbwNeoXGCL7wD0Nb3rM8Z6uWKtUeBPTHS
uTZgvVmbA786iEj+wsQwgbi8cI/mu4qKLWUMdizXJoglkQoa8DE7tN+rgp2zBPsEW9CFkNAC/NCK
dGaBotTGw6ME6GYAux8dCuf2+prolcuS2B/0QNVOT0pLVrZa/CDL4SzMiWjWB6dyjHxr4hIl7Peq
m06tVtz7CSfIVAFyp1J+d6hEVEJriubra/garZHqssIRBTZXhYgMW1UPDCRppwctHard51UZZrTy
tMU7sBUlxA22BzN+ILVLuc7HVXy+K4wbDaOOtZqPv9B7mWxjmoJOJKPWLC1Gorj7YBagdwfpnRJv
ejZ1t7LZlb+cSTv6yPixPH/6HNbTcb1ev7TnE3U1DTgU7Id8EXLbnSvTLSARESA+F/x9kZN9OY9R
AWvlXVNQ2cwMjO8c0gvTrfn/SSlVsQ4oN5uwzU/lJ3b1I6Q7/lDfOrKDkyo9mMH2pXU6aYpMYy0H
eezrBMV+S71Ovax65lxGHSwvZZUnu0GtosXdRT7RV+HS3uoVHCf0DEoU99/kWakyZCxtTh5VL7d4
RKqF+nLQz3J02OK2KMZAMv9GjyWBDQXlzL/xXph9B/5jhBjEF9aAp/yXTnYpwLm393HQHWSrI2Wb
SLPZH6t5WmQI0OTql1HVpMzzk8+szeL/KDoVUdvvXm5uiC149JcltZCdAZowJkfdn2aFcL6h3MZi
l761izXyZ0mG1x3tko6MRuO/N4A82p/06e7QumdPwjJrFtwsj2xTsWBoov7Wg2Ce3rzS/xSautSB
erTIde9LMceEjyXtIcvOj2NnNHm3ydyjfTgjeeOovT5U06SdOUOiJT5rwAHyTQC+iSEssf+0Bg9r
vs6bgnQ0TC4focm+v7XzxWcfjbWnN44aR6dyJO2GBRHIkc2sh9/DlOzvVlM5BDYZHfYupZaU2I2R
6NlyAYF5HubzkBQTPyrkVHWwmKvmFB2SIVpR0cd5d4gjsBFi1fHYfIbjk4tY66q4Axgk98LReoYb
3NqNl4Ev24n52i9ddUn8igYPLZ55SK53mz2nEL/cUOPVu2S3rt/qe3M5cYj2P3uO6eMdg5ZBuC0O
mqEc5w+yjcYuN5UqBrDfH3j6pxN5E8LW6EobJ3cTS0EnHBgxkKVsJpqXxDF/gBEc7nu7d2uEmZhj
SmVo1BwqpBwVMPNXChKXK3AzRKBb2314sjoTXPFn4Eaxt10r5DrKb13C/FW6Hr+UrEYcqEYYYUvs
/pBKNT+IZ80rxN+BVSlOLkShbb0MZuZMnL6oOfaVXlyFabI7firlDstSnb2+kwGr6us6Bd+GYpVx
eGooULGeZxWGQnkYbi/wyebeYPqjR94awT+9Rf3NiOkX1/qlBIuzynCjVmXb68b7iWjoP7VdGkp6
KLyS402TXEsdvzM+IijALAGOrDfeoX6gsh39XG2Gg/hQ5AoaEi7GEkCLhEmVL6hI80HoSWxOS96m
5v2pBKxGemTvAInEmrW0JiPdRfUYdXkyy5Hiax9i9/5Kl+gVZiP8KndXN1C5j5baVvHLJ+17omc7
qVkJnS99P+U8lBBGjJ4e++Ws/IPCZRlZRRomq65L/MW+F+rQVLh8nbkYAUKPFWyUEm7g+YO8CiFk
/JANqhQLedT9smzB6ekSE62Wd+8zHqHkT/aDPEUCok7uOLX+znoIcYjrEqTc8L+9RPnrcS5S6j4V
0w1ExwB5TfCOAGdcsUX4Qpd6u8MyUzml4gBsnXcjmVK7QedO3WKkbenvn9jjBeIqYPmDGgVcmfHM
tWun7Da4JJYpLVe8ZpIqZPJmEQmaZnDOhSfKXvyEhCKxXMVsJFzvJWhA1ihbazSpI8k6AM219wYu
hDO1Dg08S/nj4uOMCYN0wjveUpcL/fM3PU8U6d1Niqh2CjaRu/fzyJd00YuHsfHqngakSw2nPqm1
Zo1qnHvY4bhtDbxsYXGkMuaAEvLcHOysIllih53S8aoSDoLpANA6apweRCCCYLGKSyErzo6Sh2LM
1rXo5C4SkUij2OwrBnQQCaPqKIXtF2mBB+JMXsSLwofwqWiA2PfhsDaTXgR4L4wxhuN1USB1Li1p
LP633WusIEBjNeR1U7AOHJyATW5YOubBIt1XheVi+RZ/EyR6hOn4rm3svOXbeOHVXNiYd4pFAN4x
a0COz92/MAOgG/om0jQEx/jw6UnzFWKnb6xXrmNRXjGumwrlObZqar6cHq4py1UxBPPjIRvEcBae
HUrFUblg81vnU776ZLjRXAJiY4aLR5AmZ4czribnQKIWmQMzrnggV7tUGMtDX9gPhfe87npzK0xq
mknM+5kgUbHJpimjnO3hhlVNhCbJe/90f//qOITSVXulG1p7Ak9qZKN59I9QBHiq61HglI8Vftk7
8LAFEZCQMlVF+d/TxCxNOiswAz2S5V77pU3gV80DIGQCypXI6ib9cnlumZQO8WDuz36ER7RGF5JA
EnvPk0gzPOs0uhLdHIKC6RzqIskAVKy9jnt4/YcVnds2PwRAN7Mwg71FaCB+PQZ6gppScUL4HA6i
gfESyBd1jWRwmAUrugfTpWMq0r/ul5L4RufoVnzV2Z0YjiYaLjVG2IhmTLSjnvr64+UKnhpghn2T
3FZxmymkD15Q9EfP/wITOXiDuIWriVcxH1wlKGoeT9LDIl88nNMkda17NebxiG0Qwz+Qwpki/RQ7
mLRRlY6AUqSSVGPKJFZ+QwesdioXb2JeNVUlF7o0whc/udGqLif2PAsoDSb0PbXk7Kh8UhWy+mxg
+N9Mo6/PTyCBywsMwYLzNf4FKJ2xKg9Cyc4bfd/unF3dSqIQluofZm67dPL0juMJNQNXFkkaB/vK
9yTSQ/5/nNkq9p+yNRHwli+9gVpVnECT504E9ZxqnGgdhDP4+5Xm6BvdU0BIXU57yIzqNGxecmrX
RuWZ7k0Z0jk+lWAathJwB/nH0FMxrjyjA3vcucoYBlLPvxAslOSNHl7PRxalYcvjsodfrjdjavdA
C8dJfnU0VDCBHpzwhw/RtKxjFhOV1W5/cB2ae8nur4t717YFJwq0ZYPBPCpahbLX9HrMSx3vXWNi
FixL5MvtSxflJnhLSObsVKOzY1wStYC2iYAi1RF9zdoUGKUrq70YVDJUwGMAx3LS8gHGR+Ovpm0P
VIML9aHpDob3GMW3IFPaUtESARRukuA3DOGeC7vSTuaT+rRdWX8XHyMqQd0oI+oxwzPzhWB0jn1e
/vWYix4vPxOk406Apily6tVC+PiNtir9Nj364N7UurHy8J6HJJyGm3yoggvPQ9gylEAK4jY+LyBX
2KsR9ezMxiOl9obdNn0lIVdQnZ1lPjdv7oQohQdl3NcwlpReD2Mq/9we7lUOMdTyMCALEsXLN48x
lduvdZorTS8XfeV6RsAy+bDovcY7koMM44ygp8W4VbZqlbhsyYdoHWX2jfC7EcPF/GLvKdMD51Sq
Nc2m3+BPxMKr1RuaUlWBPrqSMI/XyBiVrXr9gjO5Ikf21XlECUiPeSKCUNwr9KIezE9i9q1hr4A6
9NEYvaSdvBt2Wq/kt2d3cBg01NyhcbN3YPOSPL6fOlZu9D+v1Sd56ETkO6YvN1I4cOh6Bb00+q9L
YFB9Ne4NYuY78ZkuVjrPqac+jRj5sL/qcVLShLx7vjJfHe6u2vRjudOdhK9LTGLLlg2jT5GpUXuJ
k9Y0qz4E0FNF/yL6LXI1iYkyBvyG3jmyjzsh+L/b4k6hRwSflO7SAmglPnww7anHgS7NNk7cGBLL
TxbDYbl/55yEGT0rBX2rgEH+yd3Q1SJLy9ztOaKpnGpcT6PeD6byPaHb5Ods51VtisZjUvPMOb9s
od4U5PHUS2yc9CnOnDnN6+39N/k6vesZNi7bisODVNJgEG/uGCKzqu/SdVaVMPXSxDl1IMZGaUcR
IiIvl9BJkaZRu6IpB3DDT9uls1efMAVTTre4DPFbQEBifis/BQEYQccvP3sORK+4L+At3Lx2MLRp
YeG2Gc0E2vEwiQQJY7sEBkaJj2Vhu9Jly4vdyqajfPXlJBeGOYEO21rim8n6BlPNrk9jNrVXJkiK
Va0BEi/bSlbejcENBRZO8ha4Y+ONg9idTN59lASBoLPmF5syjk1TyoDC8eaPh6CmM9a1Kkms5XW/
BCYB/oACkHP2X7SQrLhgYn9r7UJsL87UPYVFPEIsNz3MLl0Qp4y/sevX42q2ji6uLZB2A+lSOAB5
roVO9LLMnWiWL9Eg3ogzuhd2n1g0HpTc3RH1b2cvHKAiLM+JvShpmdHiOJ4MV9GHQacsKbpevRJx
5sycdqU614Vm8VIPBpvIs5B+svhl2S5k1OrmJ/apuAb5pjLsR4lBs/bNGPGgwW/Nd/ghGk+wk0PD
Imo8EmgafDlVpT5SgUFqDKH+Tnc3nvbGMwktLygne1/NMyr69/p2TmBRI//RiAewkEaC2r53vLVR
nDjou0Au4sKkhXtJuIZVaI20X9FPBN95tKsFviZfp05o9wLebXps+pFKPiA6iyrLyRX+bADFqIc5
Pzv8fO0OERkmicLo+yj8I5b/5T/1lfTBw4lSsWb5yNT9I8wvkC1xsIdDK3SmCr+fa87Ot1Kfmh5b
jl07ICqxi76p0uX0CD03K4Wh/bspiFhKIFgO+LQc/Sa8yo1kemt3qdgwXsGYTTcpPhwfrQjM8UNE
vfoj8Kaocxed3Mnq1tqLLHADHG2K52bs8okJF5rx8e0dfdHwVPOZ50LjKNaAn6w+Q1jGaSiuinT+
g6CHe2GlUBrpeYFLOD94z0fWXZ+8l7NV7mWDnA3JQBpXATe8KZaZSwOCI63OfOzmDd9Q7srVBY9l
pV4bsSUcyD1y8s8l5YWzhI0xonCVPHA+XyPbvZV26mx9fYPr+Ut6xXnreJ2639zfflBig8fa7uyc
v3mhYMjmqNst3F1rd7FMOXCmQsD7df1wqwyHITyKcFnh+7NjYqUMotu5qVAp2CeFO5umoHEf/4hp
TJqYdoRLgoiwGz81ld4PbxSBp+n5e86M098lJqi3DBbyqv5KdKvP9EaVEZWkBkTIeEURDRt8xa1J
QAxqeAHr6YamDGTbsmAkrLX7NKFMAfnoVckhf07ZKc1QuT3WWEZQQLCzTk1D8iewv5UxbbJ0IMH0
g7qC30WQo0xql+yRiQqx+FI231oswufaE0e+WRYFqq57dGfU38Oa3jOef/aRte0PC+GxyQV9zB91
ltQkCWiVgz2e30fmt/dPbqrCDCGzQuKxxK6vOpYMKPfDKBZtCoHSEvMIBRwz5HWak7t6E4b1/VCP
1d8VbyWzpEbGQ+Ehc+aPNh/+SL4Py27vtUjg9HxBCNlJAWJFwgsAT5y+quP6vblLQArtDyezj37V
YuQ4WnXyeMo+Mf/lpl6cy2HrqrFp58DdMI3MRTo11p/GunauBTscuq/wiqrH/IrIUFhOyFwmMSHy
ZFWmPeVH6KazxJHYhBrxJvQz/FfIgevWW5fam0I8ltkLwyVwPPmRIBVzHEduCRxGxH0jfukrNAoq
7o6t36VUZPQ9Tf9lMqAo4VuVky4BSf1FUEVZ96JcUAkDMVYpGxfUMZa8UB/w6E2093DKjLStJU3o
S3Ccusd41DW65wF5CnCYugFtpT0fvfWLDd4MAQYYkM2QLjF4iInRh5X64VjXSJBRzxCymOpoNRp9
7ho6yNZmH7xoSSQ0VuUKBR4Xh+yqGbKKutNBCM5t1j21XPYnCh+n2DcsluF4/2TqJpf2q7U9Sreb
P+dVphNyk8cV3Dw+873PVPAnJGL7kjyeulOFak+lwrqaIT90eOEinc94FCmJ3Qjxp9V6a1lPyLI5
JXUXsm/qmpHCY0SW/kyXFaeRwv6n7Cch/4sw/SYaFJ9QQtUMAoVN4Z2v0U+bq+1iO/b85fhSAEvU
4BwqI/MzAxIGLI00nKdFCpl/wuFXVO8eEfoMtAUgQULq7AG6MDrrSOZ1WIAuJDLWJDugVTv0XgS3
jhYOhPbVnBdhfuoeV2+lKLjgnJh0yVjRT/YCL6elLNafZ4uiCE8Qbab1AuJkAAseZbGBoNdeZCAm
jeq7UauvJluvMWl+f0q/xRtrMDHP5o8d6po9u3xexkAvTOaEHhzxg0CHMydKGh9nvimWSs7Pao8E
p8GhhQpkrTpwV2TvqBgyaWvAWuaw7nacNGj/Zm0CJhH5uFChFET/+d0JumS1wNGhac7ziYIrJvtk
R7w49Q9xIQGvf1rNp4sTMA0i9vAH5GNRORwv4YbbXrL4KUHsNFFp/qYs+CHAO7MeBp1zBBc/WU/R
I3BCQZa/hQvHkuiK9kfamyhEW5h7O3Nrg+5NbZDP7bOn37h3hkivG/YUcdQWGeCE9M4Pn5SQzWhu
TjA8fRz31oVJ3EloXHTWoNurEZ6dUQmaZ8PXNCY0kaJWAzA1neLSGX6bPMKU8zOcBG278pwJUA3r
Tvb/G7lFUbTzV0v/qYk+YzhGhSLQzUoxzaHvAfGJm7VnWGg9PRv7CmwQB3N52vfoKgo7KU3sI8sL
uH2iyRMQdK8bAlK8kdvlcRSRDvLEYu7jfWMwckYQL+Vk9I/6gQLn8IlAfPkkaWESJsk+FltTt3pC
st+gHDS0X9UUX/7qUzLUxB+uAalzA5RBbgO7YmgPdgGVAC9RVpnMuvFFTb3UJ7P6mJkHSE31yd/A
8Q4vanB/WosjaMYAto05gVOdRa3LSdUEfFKwi0GiFzJ4b4tjoe5s47a2x5AzNjypUuzHAzTCMLk4
98YidOCg6pRVm/IYWstbW9Yox5fL8SBtEByApCjIKVb/FnUQOHH/LewNGFZO9z5Xdacui1pDoZB8
NK7ny9j56XMTVgCDrY37ZwrLZOomJsJnk6iNBa1LxEw2OfTPnP33BXgTifbOtxR9d6xkUsWmX5j4
dh+aQ0BE2mHDKe0dB7Skln0HUPxmsrpzl3xjr4fH50rm9xdUmGMFC/ISCNjipmZKWPRNYYw8Ma49
ecR3WxaqRGJnx3fsDXKlPXm/HLF5bZAmTs4+2utfNBv0txtkK+SVwhx8Low+9KHXMbkjKVLz5mUx
3SgiVi4+q4aZMo0U1yI/ADz3+wxuHiUbCqnEnDkd+Q3/x5wL92EFRjSC3bQG2k95Ep8v4KLmKbJT
kgteK/xRzv5UPkd6wCc/8hkDfH8nJ+ZnzFhIq+VXCJhQ4k//X8fvJaB9otBXnFs8KaHGN9uyzsI2
V8/AVsufReR+3W65KA7RT7E4F0jGBU/OWg5Ncmtw1xLif2Wbxo/cdFgMrOq1oUP/43pdBshCPtNS
W7Ptdk/KD3ydk6i1vHdo3FNWsMY87bZkqioXxUzM409z+LvosqLFBAWvRQvPxdiR1ECKZetdNuGZ
4nvCLMQJMgY4eqSMkYC1OUGTtyMN1AWRzoyyxgTFE1wi4Gx0qm6NyDDpFLng9Da6BwAfBZ5rNXoF
Voa6MHtPYUvLZNIaDRcSodU31gbwvovTray6a1L9gCww0WVUGp2iGUyn7JFxxsixHtUj6EsNM+Z/
3OMJMXK3vT5AOzdJFhv7mzOqXbSYIQaK0ahNlrWzte5/GIAItVS9ZeUYafCa8wdQN5FTmsAXrpeT
7iX+zWSqPPzwhixmW6q38Ys8mfIjU11wSbu26hd5mQHcLwHOGf7syDYcdg5Jsm6h4mtR/2VnLvbM
w1lYdT1ycCD2GGuhkFsO4z7H5HQJW+8+rL2pkB678WS5Deb9BAFalSs14oO8bewoNbHaOXh7NrZu
M/864jTib8jGMyxZQqDHQwd9pxkPmXYBcbEKlrOabUe+JRC99ALs99C/SLejxVaTAUT0YXA65QDQ
K2otxLzFgf+1EF2uMS8wIpFPwHXM/7w+OEf5iqR4jqbKPM6Q/CG025PQ3oSBmkxKfR1P3fZRySi9
GdDe48Nfc8FhwizQovZw6pr2eoCAujt2ofYjO2qt8UTAMsA2navqBNm8SfrFedmrYjzrClzY4ego
xMnJS2Ln+2K1btp0yigcXF4qGBl5Ir9p8mzIlvd+uJJUvcKH3vIoCrNaFdwCO9xCdAPfiEwor64M
yDUolsla+PZPUXn1L/jYU8Vx4ldm0fUmSubCKHLhrZiOJ3SB4kbcD4ROlUg4zot1LgLl/TveaHNr
5JMPQMxxkYocMd4tsunsDgdzBlWWfjKw0tQ51I53kIK0krASScZ7bA4DkCDq+V01dCqVuXy3efn8
NFjmOlqQf9L7LaZU0ipTXzazxQTWpocZEReQME9bLRJHsZUUiGmb+yTAYQUseDw+iw1R59CxRNSz
Di8/g1wljiFEZSmxl/16ik/iO5kdCQW5lWkvxPKwnY2lVFpTYL3oTwsxnSHlWE9//rWPQf+LPkcs
Q2PSpMFzRI95ae73K2hd8+zjedbA/LeyMd2DLCh7g4s5185A1iaZWA0QekXSPJGQQdx+VQ/ldTMd
B+9ONH4WOszCpYHVD8TMUpFwj+Cew2ezgwxfs74DwMyHPpUm8M5Ed1VpAjyqzXUKZfnufN/+IWe6
vC69IwwyZPUQPZW+9EnVcUXWP6EYPi9mttA6BjLQq0nXVq3IMR5RTbE+ogo4o/a3/T4LUzQh69GC
ib8KfdwoCSil/EuM45C/jZWad1n+L0NSX139RZNY/FGtol2RfpbQXqg+CRO0sGhhG5KaW6iHN9+P
ULbaLyRdtykK1nwcG6R+/u/Xoyh5owPZvc3QH+QqHVDiS2NG6NW/3IWIfSV3LQZHPnEcs/lvCHRy
1FkUdQ9qIlJ5QrunrkWqd+t12RZCtX4GDFTOQwysCKnr+pIVtqv/nUv3tscemiatGr0r6Kc1ywzq
CYF7anOiICQZaHHaky0a88kAFqFa7zxrfONe8QCpV+3aLyG3G34cRdl1BwZsivof6yy5sOJg/f8S
NOReyvt69L6oSVxJ2w/AsUmiwfhXkeMbO23FTXOVmduTqzs3A5/ad2LL3a48RTouLyq9P3awiE3P
G3cNGZke7PdLCz/0uha8ZiXGX2KqgqdBgF5kcxJX3Oqek9RzyraL3E1QfKOCcvQwpy+valXZiut7
VfI1kKis44lEjHt5IWw4m5YdkSjg/JiLt4quZWl76QefLpdH7JWa+Z/5/XxKo7IUSaaIJe7M0k0i
uDRpDzJZhdcA0Ed39bTSEYYQXkNQ3i/NBIHvryDgh2ZYjr3be0KX6ZDfskcYGjDF60mSb/AsuAMM
6GYhm8swsktLNvecOQr21uqQLm9xVYa/uJPo4cNHxmsou7COL01QfBxCt8MN8170hQYXwUn0tbse
K+8/8yjiNOJEAmEwWPSdnFW6VkxQY4KU3vi+FkEn5OlOtUVi+v9MOeLE2GjtEiKo4ovTrTBQADNu
iVuU0LG3gT2Q/2W3f5A8fIX8QIjSuh+Fzwes49nawnJQztvhK6R4jnN87YOGed4qITMvL8BdLIRC
ENmRtDeigun0IHS4AvpBFgwetlNdmtrAaRXn6nDrj0fGYxLwYdobwTan1eaN/365uycPsL9kTZLv
hUS+2FmsjUvtw/3QwHL/EFgzbrOgEnOmxvE4OFdrvSN0Za5MAU3qkd4Ii3ErFcIhJhqkdY9jpOTX
vsQk3STzlCpbFnhqxedU9qdykdW74SA5qWG82dTb/TCM053SOE0Whe5HAxSxOmi27dx5qjk/SuiP
iC6DZieeF1YQrJTlT2rQ44SaUHmAGbrwK52w0wEUbV7VEXfWZPoWJQw0zCycYSceJNypE6fvt4OG
sifQhpxpdEReWtHrjvnJWD7o2xSUOVuOV63+1JlaWg5Ogh1iO9OjeiacuU6MEEcDMqwe87wWiRzh
kIRbM3S5v/c4fM6xP8Mwm452ck3jr3zQ2+Dr3UbSZ+wLIvjsqKEEuVcPv9vZ/OsBb+j98S55I4HB
EZxQtEfwgV2HulFn244mFHstKXxMsKSC8D/VudAw9cU5HFp0gHM1t9RHEqUznb7txtZUDBnl1eKv
4xZzNPBp0YFC5+piUiNJvt9CFjvINMhhb4mYSBvmRvHTRM2pmCJJ6L72VsyH0G5C4I11uce1G93K
SrzrWXCERMzUzpjgqikde1N1qyyb0unc9m3YxlkblAH5zS6meVo7spHvIi5mwhnSDESgOizlLHb9
njphS/ynkQXU5lZIqeVd+KHyv1LsPmsJEdZJPw+iSeGrBa+N04PGGm5oOo4yhIMwLYTsa9DayPPh
wdbpcDiyOQ5/WcceUiZpTTXx56Lej9T6a2CIeQ03JFJ906I2H5X0lcBJE27hmeDl7gl6ICd/Td0l
r8M8YourWp0Ivk4oLfoAHYrXgdOMcEHqbe073jGQXEgmJ4xb5HWfzgbYnE5w8xyET0ExplpSyjHL
9L8v2T9tizApwNY8GbvVRTCJxM64bCHgOLAYQQCYzNcmURzMCBMXnpjeug0E5crZ+r2/Ar3NAKYR
4xTV6YuTWYwwwpbCmBv0i18hksRbsSl+Zt9QOBavNzL8Q2iNSOfuf0W7aT3LKXlo88Yyx0oChNuR
q516nRqSVo940DdY5vLGiwCKdhk2vDA4ARUWVRgRegG2UIyNcvl5Elae005NgTR4ILfQ38/u2PX4
9JMTuzMXPuGAgGi1upeGbGIOrhPcIi9mhjY6HwF9KxbnjdnGItKUPD9l9Xtu1zxZ+T6JITdWLKUc
wYFqMD7rF8lvLBVHUvFToflypSXue94+uapqxbXaRrjjdW55vpg2uHdUAaO4QaNJyUT6Dn+C86ea
GA9YkRHwzt1FToBpswsfDHGTWTL2eaMuhjGIxK8QSo2dLZq5W77F04PCyGIM409IOUSdcunx9mxM
LPcNGhFbbC5Aw5nS5F9x8ZFdx96xzT3tt0b+8MhmNLVqySU7F0vEQbKVkbrRrGtB4hjA8BJjO5y1
tO1Bs4uujJeQaRcXkK9HFduIq3zrkdb6u5UbKkuEmxw98A/FRkL8f+a0jNZz5ppxDht5CBxQuNRF
1QKtQPkmn8FgysBi6BYgtT203GjVcyQsI2sziqZRnZrBhNa/+C0bXYAv47UAKionKGYLEDbMHdi9
h/wK5xtAs32plCh/C9ELc6ZUH3wBTAKMIb6n6P3r5SOqk1rxNQBM4kN8pE7uEjhA+qFOEyNkOvQv
NKgsgMtNVDHufBz35NJGRbYhkbMch4agN5qGnxJT9EP75lNG6sTaIKpX2XvwYMX2srLNsBYYiDFD
2vWikvZWZwyUeO1yUzftFr2ku9YeaMcKUgKZyOEoj0jRK2+FA0isXbVJCYgKNXm6pV5tK1rXe7qo
TPsmPfJNovHs8fuS/oqSUAAUtzdmOJ+M9+J1onWtaR4uOXr5tBGWEBGRuKOlK8cER9bJtox0nTqz
jdH3ym7PMeJOqs9vMQVqnJ7Lv56+0RhnzXzosj7nEezizoXkP6dvw5E5kNF1CYT0AO+efE2L1J+i
QhlHDQ6rH0/7z9Jy+ENzhpS3QAa0BqzeT2oe6nGZQ3jTsrcJJ/wFIkSUgzDxnA3NMuBkr7lDRtUi
beRPacAo2ixokUDtlT9/AW6P9U9PJZqyGxxOM/+SZ1mirI9ZvX9cQy5iUAtzdMTwUTVJzSlkPmXA
ZC3P83YWAel26yHZ8r9sk/FHSYWRlmO4wpey+u6n2OJElLEl4bthisrWYU8Gt5MxvOy8mlB9mWib
qJGr+iyMJS6NsBMyy6Q4kbFv5wPiMqzrSgL2lsCVuH5reC9DCT6BHtMdlZJtTduVHoVbhHnusmv4
ZtVq97GEau94DxJuYgORpGEKR9nPg5k8VFLecKdjsFfAvFPzSudt5lFaXQ+2zQ2CWDUyK/ISYwGU
bqtwqtv43xbreH4YBPsjKDmeyPuyXfDqbNCZlRAEn2uFZ7xwU5WLSaZblVYQXtPW5c5c15Dk4AJl
YicWb2A5CwnLyd6am4ed1HLEAsdNQh6e0rA0qx3yZK73It4OqoxG1gU6sL7TZP4J3X+H2QZWec5L
09Y+LL0HagHKlx0zisQrBNHD/WawHkM3hJKjaUIxkx7c0l6PmqI9lll0JXyeyQzfA6ykiqPmWRo5
iLCzggLM/5jMj761GT7FC6ojW8XCYeQaiB9rXdzFB+zCoB0mc4oMyQumoOTARIZRwnBSw/qdOD4w
caSXSwGrcHbpwEAPyzQAge8fDwSMM9tOdZPgXIEjGP615/EiKA7G599cZKBI+F3tVB9E0wIXfYPf
bu9y5eqtii4iscb/Z/d+xc4FLG8mxW14xB16W0n4NY9HumzjO44rtdX4TiNSq3HK1kXXP+rO+Cuu
kYb7CgYSNbfztXl7EEaETqvN/v2e3dgEGvxzK/ogCu4VU+jvVoR0zGietECl0+pZPQe/sRaEYz3G
8LPA/28Dsee3DWDjkh9LTt3dEZkjJOmJNa0Xd8zj0hlSUPeYeV2iU7ylkjXJEmaWjw4OU5dC8nrz
Wkoxi/boBp9lTIQ/2SijxATE4ZO9ODwLb59paJyJuezrxSXuefF0nnE6A8dD7XH7GtL1OYam48bK
pmLmaqokYiWKpnY8IsCDAG06KlDDNt5m+uG1PRpk5gZehn1BHE46MJKI2TBiVW3QRSW1EfhkHBiw
MjpR64cVRlZkxr43U7yD8Rq2Dh7VOxIa3WsPilX4m/VHzmI13YhaOngp3bYyyhAeRF8g8sd8TxHg
5wD8iTVvl4nJGVfiU3nmlLE0LLbg7GGqPB+5eOq7vVMLyDysfvpE4wYTdeeaq7ARaVjQRmqIbxpM
zHywn2ysfTVK8MDLmUZ4+P5vMPauMGGP4Ac6qF61ukZDJ+aE8AYsduVLgqhbdnzVIJG8fLdLMSRH
dRP2maah98qcUrUSPebmJg6MNH1wDu7R1C14itKvR5wjaGuyLfDQX+WqXod4f10uwBB9NuuFnfz7
FMR3XoIGQv6tFja/WR/JWEPzrlyTv3112msfyhFA8sAMbOBE8OCxvpcKhIsCQfnYoc6u1M7k4Qb4
D+G10vJdnmAGCKy12BrMtvX4vJFBbAYdoJL21D1xeAAamKkTsOzw36+GD9NC+EHNJx12ZhZvPULC
TNU/aIjNDItX6Hei91SeQhVcT2Aad2SH5sXt//w5YSV88Sr0vFQrSrOF6c6jOkQMKWTFxNhh7gV0
ryozmQbwYL/85KvgevnyefDNvz1qGIhAwmdfUPeTFQqBj8Hzs3YgfsLOGIfC0Cs4J4vJh+0bMt7d
usM2rX6W12eD3M4iCEC5EYAy4jgDKxi6KSES6EPLFRNkprFzVhY9HcOA1337vRVEHWqEGo5QVz8w
y6FiP39Z8mPl8mTjbpXXP0ENOELskltstgLNJtoyupUitGZd08Ov9Q2wCqmfGGHszbU/IyQ9it2e
ZY0XFBzQflUwHtHO2UD0yEa+kyoHzlf8kJnywmHBm2cU/ShlKKdUvZYM6FwJSpOCGCQ0RtyGNyzM
PMe6Tcgz9Q2Wl8EWUOdl3/6k6hf+MLOkIM5T+KWx/e1Pm13eZ1mpyRDtQxyfVkqsk6TjxegNx197
iGdJk+qWdwnGIIIvVCzrKJXtx74kGLaUyU9Ks+MYhfeOkgmqKvmDEM0uLMXtJXwSKTwxVVobCL1P
ll33AiG1/ngAjyQKfwcYz6eA61kerF3B/oSf1KMRlJxMcvdBzv+BSIXf2HV824zh6/WT3REAzDZc
C7z1CGoHH9/sf4EY2PP3JsqZjBErZRwbggmySranSfNjBUJAtNmS+cVvX3N1NzIV9Biu4Ap0K9gn
EUhIEMT3n5Mpdt0ugNvMIl4jySmqEjtZdeJ7lkT4ipkec7o2eo1S6EwjlLjADhtVNjVOUw3YMnI3
QUhJZUh6VzcvewY4rq7c9uUBPbRRApBq0+JsZARZ6ll3Qs4104k/tLgnN+8JbG035vSqck95FQe0
fJudyRLdCJy95qzd6ZrA3tPqd18TLuPV3wlPdyKM/CdIhPodqLEuVDX+wWKli+PjGI5YPusDekwj
WbWLXj6CDqyiK5iETxlScJawoB8puFlSCMnCkT0S6udpYealljp+MGf78c0Lo+CqkFkv6VdbUNsf
DiJM9XLXbEf9/12mAUfpgZaFHAzgx9AQmu14hAIMrLpbDsqFLDgPMDz6AXNZPnGBwNuH2yMoawvz
6ygRlBTZF1BE7ocIggHV6HM1pbUn47ClFdKPx9EVCJqQhPRLWsNIItXicbR+EF4K7W9OGnCAIS7c
GslKGir78SgaE4EjcNIRV8fuy7LXG/6KCmpbsGHyIsoxkD7D8+T81zNXm0V6b7kE1YzXvS3rJtfM
ch92G0UU5srjjFj2jBelucDSnMmGRs7SKSIx8sjD1eVq851ge6QXyTDGuSN/OpYGNnbQ5N+NlJHH
38tKjexHxYD15In0bmwEHeAe3vLft9newNLOosd9rrlMOwzANv9EVHkoKrrmJGaa99g+TS/bADwV
cTTyvCjs+n8ask273HBJ4TYqRfD1nOCJraSXffF7N4pYgR+ve75Yj+MVhoX1hwmfD5Rcvx1MV4G6
E4QKtRnsVYPcsl4SHykg5ZjO5N7huVmo9wnH/RdselVOvnQgs5RwiVBXSbPUM1FySX5MKkeRfpgy
I370jpGLOMCZoaeihAYF70FjuJ5BL3Pd3sf4yC+t3TCxSte0P4GQ3SvgTSl0JpERroklmUVzydPT
NPGngrgVUqazyYoTayH4dujDbE/XlaoD4ygRK6y2WUslVaYB+k8jV2eIlDDU7uhhR6ZbSe+z6k9y
6dfyuRNjiXZsTcP2zixJVSE6Pf1b0rce4Mj/Vk31/OGIUkwQL8rq1Ku9NxS9YuDRMkA92wTIL+jl
2VWO7PHuXj93QN7q3ry5mvWmEpSmznJFiP8UOhJgCtkJam5QNJmtry71SkmZAUjdS/aogkVzzToD
cOWFotA97bMay4WceSFDivwAWLUaRI5jdHoXuXXtt0D264J8DGg/+KnHdTWEBneNrfJwy8Wz08Kj
iXxdVXMqDUMKz7A+qQftprlZihVcBSfTvt7fTjqqwyNb3Ull48U9oqi+/H1D88Z3UddzS6Ly3oDu
Jb4r7plTd0c71UqBhCQWqFV640dOEr5nNjj8yqH631Wlzr1bc1gUFwzkLuY9BR4rALZYqlkdtQkg
XWYEpdN5PeQ8o9kve2qYt14EXipTfKNOw4YPwlIWVnMGoBf10drQA6O4NhIydSIbuOUfcqpuqFrE
KivggAKhLk+MIm7dxLb8R9Q+nvyFLQ6apLEzGrs7rA28J3GIPvflEH6yCYnKOhZzC5RaEXI9p4te
USOBKO6P+KZDS8u3ExXAcpSd2QQ+Qckd9SRvzXsFYlaEDox9VhAEnSiMDjsteNAF64CMD1GNre1q
iVE0FjxkRu/x26ojQZE8ynAOg+7oJCUWvxzTYIeznkfrl7gPjoDb6mCB6oNstSSBwyDJzCPdMqnj
zDVHm/QuczXy8NjN0jBzTUo9AKTSaMf+c7x9oWmYUXWkwc4ELsyAaiw6nX5ZehTJeY5ZnVJBhqbn
FBzVNazLfX41FtlrpxPbZCd7M1O2VAdbvD6KOsH+Jk6tAgJJPYJtbv8VqEmOHSe2fl3ZtT8GIVRU
06b1TbdY/igYEFqKvUg3WS37WKKCKwHdzqRmVhf9e28pxw2TnzUnp2iXO5brriMMK0+YzkhiWAzs
tlGcxFlYV7iDnelyZAIvOb0krS4T7c1Tsq5I9Ln4bQB1A3dqctnBdaOuTgaWcRCRz7JyWvGgy5aV
ntF+2y4qgglOwRw/aDMmgBeviKdcViy2KlnLyNqzApo/fAggTmLTqfuor14mbdMNmfX6UkE1N3iY
OSyWMA/ebzA4dsX6PBke+1UI3WVs6but4sTlQFg+umSw1xZTJZ7uDvAL/JJM6ZuXORc0KH62JqpJ
Zhwblk/QzdEFsvK8q+AxUbEq1iwfT5K0eIFmxWn8w7femX8Az7EImJvMoasOzrT33by85UjI+C2V
QtbbyVHlpDKkEZavojb+F22kay36WPNeCWAHlVTZRz146SbRkqkNGJ20FforwaMHStbUNJ/Twf2Z
1L5dtFBGGFA30SaCOzGWAkaWMplNAQEGBZkVMuCLxGz7GKbG2fkQ6O8EvZNuqtXtXoPEHx7P4q4K
Me/cWZVq3/IP6iyMvIBKhTx9DR+bsoNOpClpJijs/MHY9Fig25GuVeJP0wiCZr+7gXJKe8MOFaoK
GGUGNk7hDCy8ekA9ywqKg06D5kOYA3axia4PS7mqgy2OXwKOftwtsfHaBa+7nC8+vtPDGhTtNGx/
kLuao4yAHmq9SmovaaRAPLsXMOqa4/xCr7D2DD40b6YY1uih1WTMSK8J7RndNrBO8e0DOUdPU84o
AKAeyNi16LfExLYlMVHiA6ORNoH8VEwCnBIm9qhNxi4SRb98R3BKe6vARXNz0bslxvfMXjyghWSG
UBAfYhFUU1wKCUXicCC2HvIkaVZlhBQWJdGFdKmOFJpyouv19gem3xRf8GD39KR8nAFk4HLDaTrs
Kfpy8N3byimmB+2w6URzQnJX3qw0KrUAEc4cW3TMWhMp8/8NPV/3bMKiCR4mT/vTcmFqRMNYUPLs
JeHE+z1arWM4Tq2g18GyvldWY8+dSWT4OKX8k7NWrWr73hH2VzCquEuKI3uu2UZI8+LOHrXSW+sm
SQp+LboTyYikvsQbycZfN+u5BoSuAoWEFC+PSWAIpFgnLelMrL4t4G+RtRu3eveVyYD8cAYrHnk+
Yj1iaOAbONoB8f64hwmTC5/F/z6mg4Zng0c/Ts/qrp7zY/5ekEuzETYX4t7eYl3vi3LSQU42FlAA
RuCsZTgtz2VWn4zOkrHNeSaKuN2/VcMD2pcOE/iit9389Z4aLN3DSFA57pOnLex1tRzN73l7avyO
ARwGf4t3XHNSIsOMfD6paW61lMxYSlpveskhxqoj21bqZP0qUYTDfd3l0V10tSircqY4CrZw5EiF
y5d+hrUpVSwzbZMXAvyLB/QLwR0lSnzeeGW6tly16PDG+XiZ16shKD8C+2DgiNipyXwRWEGvGIom
7TF4rXBSieqpCa+md0EckQmPmsMHcOO4MU81aYlywQgDw2Mk3zTeDknjfLxFq6haOg/CKpzmInRo
BcozzNma9xe2xBqnG3MyOOktM66/va4DYVxXNlJTM/LRGaxzD7tAdrqFC2XM4cE/C+7LSEumnZD8
O2VQPjjeidjDWhLHHA2EQgUo5YjOwicu5h2uOEEx71Bo1/3FUK3QDyShpB1C2ws1W0pV8Nvkpcm7
MVe/Tp76aJn1nUeXty0wnNj4Y6JK+PSWl7BDPsxysqr8bhscE3WfZJiMSg7xbFYu9q6cg+awMwKp
UXhcxFEH4GuiewkW3pCMKFsrmvp0366iTVtt1vYNbBDzPHvHEpbyLPP6e2svbUbhdGUdOEMMrNbi
yTqB4hxitWHPhhycpDFM/gEqQZujh/D8v/a7WG527vxgR3BBx/HREuSV8we3QDl02dsUXROo3jbI
RA8CzV/OOMcfBUVPatYIRL6ehOxsHj1rTsDk3x/3vRJRve9iKtuRkEi/EOrIRi+s55GnFHCyR8Ub
hdQ+0kEWllLh80gxG/G6Q2iBPGXRUM/BFGbIjMqfYTdYEClqPuaG0OHMRZIi0ecn7IAt7mWiZz5W
9K18/qkd3DhUUUT3BtzD1PQMIExPb4aN0VW3MInX2souf+vDnk5W+L/lYdHXlyna72xX4HcERxFE
ngp2x/WU/a9vXd2rPpORBXSpRAHAEmFNuuj9fob4AxCcaPCogr12lx8JKpL0OtQkvJWe+gajkSW4
/MzMbSYSxfFR2084akj3bCVQ2ddUnTcZS0TzdsfoQJ5/sUeRBINeoSc6+lG3yVjX6uXFHHRd8Fld
dqq0MKzCQSZJFj1099XlTIBOLWBHP2HRtVZNmU/47DZkJ98/iZQdJAj76O1h7ryDdOzx2wX+uf1B
IUH8tthP9xHwpY5ImPh7kDIv1RV7gRKzB56SQuIECvtJWK/BBreMiKxL8uBU5w33KpjxhRe01HzP
CPh+DsGdVsfV7ExOnUd9rYTYHbxnFA7gQLYybWTSh/n8bHtV6cU+2wFya23o4yL8+qqWTnU12Sya
gUTDT5Qk9fGro+JUSdCQDKpTx4asPgvuGOmI2Qklz5P72uUMxMX5oWWdkXA1dgNz7J8zEeECNc56
/7DaLKpuBEHbVL+WRFkHSbwFGYMfYw28RVz5tDzHPntz9G2OKothMmfBgxAb+tikGhCl9Hz3GPNa
Fm6XIclvaxEEY4RGXkLaH09wwukkBYQgtg8c0TLo4nmdL02jMSQOHPGRl6pVlAgn5ai4nyM81Rpe
ijOzJJpw0DpFXfyF4W/jogu17Qgz6PlaEodJRboFGINg2pT/XU7Lzp6iuy7nnVRkWP+9NiWnkfY3
Anx3gYoWdT0LAWi0WNNh77Y+NnlWCJXzNXIzK/YbH52AdVI4LP+rGC9R4gvcMVWDqii6CCL2aav/
LSM0r00TboFAuW0iHe0pDdpaK9e/0rpo61Ki7JE2IKuAlidR60nZZfsysF++1UAgbiE5xoTg1Dha
gs5Vp0gQDGLUADAGnSOkPvrQE4tX1/WZB7pA5Z/xi/BxErWD5dnpsuk0O3IV6HY7F9BrSe+jlTtY
jAQSBn1M1fmJrpTWkSZUTUTaA6BscoF6zuWhcRLO/nXl/5XRPcllRPzBOvnSkvTpSjBOzatTb9IY
zwqOiqFjmx/8OQr9woASveKi0i7o7coS3IiYyRm9SXtdZ9Qd0NrV4wCddZAh8/p6zt06E4Ja7NaD
icX56ovCqdyK5avocqjfm68hoDUdrcVMYKcmnjiGX+VYgwLlI/OHrhPmPod7xs7cAW9aLM/1qjGV
eaUX+jFQZImNrDYE/rOCm7pl2BYqnf+5e7VnT02Ff6L9lOp/n0gG0CI6xAdIAwjwOEpXope8mjZM
tElLiQEGooxcqukC8pEOwdy3+iGz736V7LY5GZN7xMcFGw8vrQV9ALnNKfTfTlCpBRqj/6RDguE0
qcKwGQdmOWt1QVETtA6UwtsZ5S09j5EhBCS1XK/bfq3kPdC9R0CkfV1PGDZ1afDDFFmYVFDvynh3
otJPAEkA7HIIPCE2PtFMYnOf8hZxWa0kBINfxUIkOyYCpz1IgVSuSN3EvXKEA73mMf4lzWRqRfjf
AcUkwz2rRFxaF6iKIjdEnDgzhWSgEMMEPbUsFIJWDpuqSLv1BG4zCLJ0lAh8gFe6rqWv9sh121lT
IvzrgbCPV2twW5XLW8inmpfMrwQVb6qX+XKRuKJWDhur1KoZ5BCbfNwP14fvW8E3klDH6pPEdoaC
vEVpXwB+Q6Az6Cm7llL+WDNqfrqp4vt2RXYr17fTzgVB8o0vZ5jbXNlE/Eymhy6YYeRi/L6UQ2R7
QIJYdRvZwI7RivCKVx93PbDpk+u/Ge17mlTVjSLosMzoFFg6o9zaA1kCh5Xz5NZX6Od75+gszV/x
b7yCrxxlPzn8driiN8nYCiKMDKm+QqTjTA1XfZyQY9ZTaL7u16crdhfGsNTKEuDGSyGr9oeam+hW
9GobDmZlI+k0Il3lSCnm9BpBZXEE09gtzpr0KTDemRiQg4Ii8FGeTD3w1SeR+Yn3baVL5h7BXdrp
4djrkwYTZB1OXzExSvfm+6DMoxvlbygzflkciNmURmAP0UFaMLS8upouaGMDS+3nysd84z9huvwF
BM9GZDOGyt/3K2iCCR5T3Fi4tcKxShTZDtuFXhubr1EP1k9q1rTz8okj91N6nZi+03DWG2OvsPqV
aNMsrx/mEUECdjGfSisbVD/66u6rRb3TMQERwsmWRzuY+yjiX3PDZqc0OxGyYdhbXmAg2C+Km6Ff
jZ06LSN4eCJly2nRZk6PlPeWokRIEfJE6S1TY6fZUXN8SeWcjrUYuSXL6UOFElflfyRVDtzl7OK1
TNlFPkVG0sxoN24FhAmiqO7kqErqiNean2Yydl6cmMvCRbfPHCuiIKm/v4f/zQRMhTmjkwWgNx8a
mdzE+VkXLPLdRfZS8S6Tw7qxuejouiCCJWzfjpQXri3wILTC/g1IH/HR+JdzTCmK7EAy1impiRDk
1wgltuvSNlYMeBlYAWUHMvCN0q8xo6yOXMCv+SRrtj7+JZw5k0xuflAAjkJ5ewjXAT+Jc0XZqCQ9
0/zesfYMZqGmA4dmY9Vz3JSZ1Cqpgah2hgoC0+wIjK7UvrGmbYA7Km5BG8feCmGbhYMTGP+i3ZfE
//0/VnyVqjRL91wI/2R1XbaKkzRsQ+jdOhFxgveMZTGbpVuqrNqvvyPQiWOayN5Z8NYtYdu8l36t
g0zxMM0g8uPe3oiuOK+aDtgMKNkmV8HJmYioTgUnZRYA7JRQGaHHTLC6YMj2ZJRcAGeb0vgavXLd
J2NAuvEdRCN5Y8+770CLxHQgt9gHsl4fynKd4zXdyMzegk0AlSO7iLuy8O6yzVfJU6U0hj6GN5S5
VhpnB7wsiwQUCvd45ZYgYGYeuHTP2FJ8kBbSaYaIvG1wCtnWpVr4P0P1W4T9mcVBaApozgluQmVE
sDAJZ4MgBMkLlUwGf9E99yPuwZGtDca/8ILznb6osrdxLlCIxuYZrxglIV0kjC6gq5kCy/7xnOUF
BvmRuiHzfWMakmIPCNm7QlnsCDR2jGgLK1044PLdPyQqPDZXYQ7N4Xlvpw7tKuS7NhTImYKRKfiY
Rw/r7/O6MZhOdJU2qSvrNUKJnEbqK5SJXEDOiAMPdpH9LohpdnQiQw28SE61IzrBjMwUdscRcVou
aEEFSUnzha7sWIIFYKPknSLVnNMw1lImGO2RISrU8ySGihZzoL5heheub4Q13G8VKF2kxVRykwlb
JbmsMYw3hdHjQIHdONr/fr/VtKshapn4MRH8VcKBw09tszanrwGay4cFdjr1u2DI2Pc1DQwAD+oT
TDwfMyGsoSJlbLPrfquS/plhUC0bIacrBH0oniMFWvZAWQcyf3QwTzwczdC7DKK7pozZJs/OSC8B
Jovktn3RUHSKuvv+YxkEwW5LoqWpYO/MTdY+sQTLekxt+CmAdkP1uW/sdZMtBRcqm5WEjx6a9b2T
pOkIxm7U3Q4I+F+rxk2MNx1reJMnyp66sc3PHRaIILkyZb9fHQxtou0qj7UO9cY9sbWhLAMOcHn8
QcQb9vX1yYv+fj5bCZg4cuB0htfozTa1yPjjI9JTXMW5eic0li7sGi0lCJy9NFFnldyEFGeEbaQS
z0OBv4d+SDpJe2M5g4fv+zY+6WzpnBgfAHbdMotkPEQzLSH790Ge8BADam5+pE8GSOZQyRhCryAz
pLP8ZWewHOB808rMZWmyHo0O9KJ4x3VNtLYA66nfA+qoSLehvSBnMcdlJIiNDtCYIh//p5Q4tTtJ
Udrj0arCWROM2aUFJDkyQLHHHuNIOfUI/8bGAP/DTThjDVe5Rm7QlJcLvYC81pHLDOIu0o4svX7y
O9BGcAPWRrx2U7ZWSFGq2tXQDvCF57GrOPowBm+ij9HftRGuehCR/ep8KK9zI1eG2rcq8OTvcC2D
45/wtwcRnjys0ni0O965vKYMt8QVpcr7CHjrbF3Z6ndKV0SOz3eoB67bf13HVbpgpM6uBe1tCwy9
INCKoO7PSOR35uexcm/lBEI+o3+YqmzLzeTEAEt2dOUiLdZhCIRuixaHhIEaNrGDMCvYZItzhIgA
j5+itG9/EF1l2BFVzdThZ1lZSDJBNCixupk5dxbaa/lxmGuSvemgoCTix6d+/MM78x0VOPxoPZ4s
YtGLK8a1hchp7PDwoddw1QndZ1qLXbGZn34LCoF6WE/RwQpgpMvezmQxJger9adESjwKD6jK5Mn9
L5GUNWk0fnkRACyQR6415rAvpzllU4z6jZWRAX1wu7fJroj0RH6bmTjbiX7JR63hAtgwK6+OXb1A
JHC7fngxw6ELz65QYjE6QywHRUzSjimdC2kb2IPz6Qxzpe7dlfkeF/SQPU6uNRmz0DlT5rmky5ns
E3iOI+m5z0CPDWtJhgAjrW0iRkWgdwjrO2/ujCccvYnkujsbWQCQpVEo+F/CJjsTpnxneMlwPNY4
8Uf8ftTPVHOBRGAdkDsLyFzrqxumq/BO8XxIVjIRltQqQ8ctwOWt7pdXdso2zllmar4Vu9rDgHg4
BvIykN2/IA3OAzO9YEwvQ7Ee7O0HoLGKxwSsZYAt5o156EjPySqC0oSBBXRBE9W8zBM3Xp+iwycM
gzvNAQyrKt7bhYdHZg3Wvr778OQgjZZcy7p9J/1ZTBE4U83VCD6u82K+bmTNw8l64m2IVilyIOiT
mEVOsLQt+pKy/wqY
`protect end_protected

