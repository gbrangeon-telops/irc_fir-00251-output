

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
FAkw7gRmEwDx0cT0lLfFXgH94E+u7pXWs5ahSt/pzljIAtlVd5PhOu9ztNGUELVfoO4Gol+zPLUh
TN9yRctY4Q==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
OsI56UKE4Z4O4++RpLw+Gr7y1Sd3eUkdDGmGZYBu0aWjoj+iDwzKGBcBG0rF5D+4LwCAgnpAGiys
xLyYTz/ObATK7L0zNe+Mx/H+/j5j5SXpNvpcXkGCWx3Mtg6EpqxneRyrD34svh6fn9QBg9AkFvdb
eTcam3dZU+Gacfm2Ivg=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
qc1VB803xD7sVBXVT5KuCy+daGAjeSNtMgViDKH2bpJoW4aexvjdVOFa9Cn3ZQUudsfzbRtbOfND
3qwRkfwGKGa/rWJp/b4u168LG7R497q3mKgxz4wZrw5VVWth06zATVCPkvVwwcP1aVCYV0wxe3+F
BcZo/LoE5dzRftELWM1hbxUlZMlSl/apI9c5DLD1ZPtssPXqyfH8yGBCJ6IwpqThHkCcKlxPWOFY
XBErOYYrcO+fou4DBovYWIgQB0ZKOhCR4cvN3q6rg5XOYT99xP70Y8jdZqXKRq3PuDDZEya4uwav
9zgp9xA7sRjUN5/fcIvFMcfDutvNPIc7IvkzWQ==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
xeydwtnivo2IBZhciZFfy3r1qoKk43zuwlyfDAWr7E6QmSwqVQF5VHmc7oNu8/L6oqsi8CW2guof
n3LQZ6J8fPLN7CBNStOEImWoOU09vnECk8Bwe5gJEo2CSwnqojJJlM/jtH5jKtWnMb5YecjpsAkT
3bnS2U0oIgAvNLFItdk=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
QglgmN/aSMz0M17AlWb9oRKStkdBh5nVOwe4/WnjlbCHuTNXWcMIzqLlv5JcAmIdzL/13EAMS4W+
LbXaFXFMcWHAzC/5AZxX+CZbwE46qfB6uGUmUBTFEckk+Ba1aO38uKX6EDual9TqDkiz6OPrjmC5
MifvdDzh7mlaB+rYqb5sjxUWUfJCpXIOgO6lavL3535AS2e2hAYpmi1PB/ejGTuva2r1NRmDkiUk
Uq0oiyBI4sQwmU7gFF9pADJRyzpgRQuSICfI5NAGRTR3by64/5TeOArBdjuY9arezL4gMGXoOIu4
E5vrAQOLZikLF7X3/wpaihrUarYdJnuPPVXNaA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 48992)
`protect data_block
Wwlls9FU/jOC09LpzLfp64uoGMXxXBycSfuTlv2x/scpYP+9BNWiMLnuvsXXVgrrh/VSAep8/Owc
44s+fXsou+GnZ322+dqdAGG4jXpI04egrzNgtHySbPkmWKfwSKCet3FW6yECnyB3rd75Gi/2z1yW
aACyfG2CjE6qiidoJAyQXrLN3f82983Mas7Hg5tIvlM6OlB5roD4S+l3v6JqRto7FUU08Cbxsi4N
H8CD+Tzzxrk5bEeQZqUipF1dNw3jLzbD1+4/SmXevDe6SYDLG7X/So3YDL3Dyxl2G4oGq1Sj838I
7XXPLnBKIKNquDHyLUzBMHkexwWd9hwlY+gNGq4rWKZG/eCtgUOL8A1XOYlTk8w9/q0jraNIPT3/
/kxeQURBEE7itm0MA7W6PBC/3CIThc40CAROUea2OoHRiY20sCrlgbhGi2rGrYWBSLbqDTVpgVKz
57H3kz8WIhmdRaf+vjYIXZhd1YyloO5CNvZi1kp/+aEq6P0fNYrgNj2RtObAcGrQVipQeZDRh69x
ABjJtbyaPuwAuJpcDW4x5ZIMIqYuJkLwxuIZllUnimpI/wr25zriPm8LMy5Sx6OAOLaWKt9z8x2m
Ge7OLnkhZQGIqVy/5i1EDTK4FticMM9OpH0v3REusyVVkuSHKtHsruoF/vy3l+2b3FgSSJ/S9ZIz
vsJQBY+zkj83UBvixOM/6kS+FwMpyqXv+qWX+hKuUTC6LVk4ZAqa/WcLIu0Z9ub8EvgH4kIARENC
Nir813VEPWWYTiwyK3IovFYi4xeLazoeluu6AHT4j0NGM8jo17UrvKc5bARzYGhZmLKIFZm8J6TL
2O8EioS2zftL4oL6HEDxbtHbMTr3KICCgFrTUsTdVEhnmViSw23/B6LV/Hsh7TtBKnT/+l96eG/W
xKjbPcdVgvW3d38tpPcc9AWutpeQ1SdhM5T5eA71GVKTJFLszta6VLywbfv16cpzeqnKg1iof3m7
EJt1KBeR1wbyoYSEI3b3HBd0rm6tF8IhD73wW1Id/xUdMm8O+zsdRSF8eIPiSUtINLQKPZL8nNxR
4EUeD/zQlGhM63ECJoap/DyYFWxSGp9Ck7cG9u6rrR5ZCUlj42MqcjgN9/l7Q6fQYpv5NfLxBDVO
ItX+vJ2yFM20wkTIERkA1hgfzG94OKNdVc1c4yen7nklcdoSZlIkE7an5z6ZUe7QBuQmmOnaFMjR
K5B2tMJXrIKumofbKgYMdvRCCZ68vQApe0LbFfDpBCz1MZt1KhqF0WX7qiGPMZnXc5/1QIDluUsW
2nLQol2TSAAyqh4lWJ6775kLkbjnB8TfkDDxhcbGclAUgqxeaVhxE98GnNX76ulNZ48+nFdHE8OP
cGfa5Y69oCZqQHeExYixn26XL2LrS0R/BPzWTJAs/XfvLU49ddISP2MHJ81x6zjPvl7N0SgQiw4E
oFwW+7Lu/mSlj1OOCPvFNFhkqTGSbjiQR7uPal0IH83PDNQU8mGNpWQvlVb3mFMUjuGRSnAKKv3w
ie/yrlpjm2HKdMY94VDW5i3SgAW+RSpYpzy+oBmTV+VjLGbCZT2i73juUUTz7Rwwy43l0wvAMAeQ
Mqu1kcJt7uMLCFFx/iV5aITlfZzOQ6/YjaGUoQMHN4E2Qlh5dF0l4HCZMydzVjOeHPn+5lY2lC4g
QY+HDZR8ph8iqJqnIJ7xfhRaLG0mvgXNVO7f8om1iTrmgsrQLYCJWbqgO2yR2fFbF2dZBqrut52t
k/SGCCbtL4o6Kd7892qz3j7sMhBynPQRJx3G2h0lXTAwtuLzzW/fc+DYvoYGbZ3fgQTHLHIl/wCL
3TAX1EwOpFeQm5aWLoHO9DKTY8N9D5MUiwEDysfJoSBfJZ2IAubdayeBgN+fy+gzMfJJv//H10vd
yBl/pMq42K1KKDK1cacWNq3fvBY6GyDMjgqQUXibArlkrz3q2K+MZWG9l2gZELb6Tq3RqLOulLcP
iCw/peXnoG+R5B9Cmi+PpSxzpfFtijIh2iWZrqIg5qSbaySFugFC5NkL5W3IfZ00sac4JNe7Tayt
L8PXh6wSK4CSoSZGkbZClCiQ9Xend6q5xCnjwP4euSHdSR1fkOI7X0vrtEMtO5v7WrFTVLyI4MBy
TbywtF4Rm/VVnafCyAdZcgYqnvNQGRrcrv56RWnK860SZOOOaDscq0TWSnSwl7RPL63XdKIGa+Ks
dfcaW/BBbFLXYYn3/t5+uj6ML5+2R6mg3RfclnadC/pjVcnrydEzPkEKx7FcPtOwPr4a2YNEUr31
euIBXgx1W5BIXvnZUJUlvG+chkj4y9+1YBJWeCom78KjBRgec/pr1ybU+7O5cFeP3Mu/iactmOMP
04Tx3UEYcllltD0h72YggQ0onYPHN2NRVP7HnPu4H58N1ejthVu47A4BP6OJkr6nPpzzkKQDXNTN
vzqUwp3+hHAc4hp9KpGoaHeP3R43fkXUYeTogoUYFhHAnYzhAj4dSiv3wWgFMEuV5cQVTl1RYdjv
Lt3YSgprGRP7wikJuYKKCqroaAkv95U/UBjI+h2mBpDe/UsaBsN3dx27IvlO8F4ip1DqZEg+4JLw
MLl6NFkkBxaCaOGZZIHV/kvLOrt2TDamogvMi6Q+8goN/UkfRqaOvP0KMT6UX8PreRbGj5ruC4mY
NIDTxf4F+HrNHp3jApel3DezJeLsNmFbk8kYBkQIuhxQI7nT2V/Ok/PCif09tzAZ4Yb2iKGw+hhT
9yEbKaDpT1LCCDjDyPHBfWRFWjVOQpRfWqve5ULkANFAzliHg4H+3UjhtQSTcGJiHv8PBM3ccfmk
JzXgE+A42DVIFB+06QaPrDNo5L3QcokUsNeVoP4vjTBEQOW0ySzC2EWP/RUQmg3eAnJL/oYCMmXB
q8U9dvqNmooDgzTwLiZUewOVGHvWI+vmTF9JCxzT7L5H/ctnC0yrrHjguva0JaKBSSC5RyNn1gQa
hTJEIL2VdJh2Tzobh6de4+Y8FsAYzuyFYoUghwLXJDVAmkArqYtnL+eN9NRc7vlyujdgQorxjjOn
D3kKl6R83Us5RHYyiAld2pzLuu6ZS4aCtHG/Qtnpkd3Kq1g2t5IFBR3JKi1sKYTJtF+fmsNkGXXH
SAawGtywB4+k42nEHW9SzhC04n75GTrnl+Yyfgv5lWKwENN20GXqR8od+NxJKIqmsomIruqynjgu
phH/IHvsxb4sKHMbF41IZX7uOFzQTYnIgBZnNj2H1m+L2jZgVs/PphivMnGkdn4OGnqdxI/gTwfK
zK4CMLboTkpRgNpZm/FljYtF2uM6nTeD/4bpi49ZwAXDx0vy1F9wseAnLoIXHPqiaorkEu8ff464
K0yp4wwHxrhtrqeqXRQce9+P6rJQKztfYnpGCjHVa6Idj1znh3BbcgkTDLlwC5Wq0UBiAggaRnwt
As8/ClXp6+2tPRiS7BJxQb0mZ0VgPDIICtS+zTVbW4NeI/Rz/Z/j0zu5GBoP1pyfyT+2SSQqWe/J
xeXHLLYHSCFui0y7gNjoWAHfBbbn/KIGG5ptj1FP34guTYf0C8ZnPWPbqq9fWUr1UPFUKtl3rzk4
h9hs3q8g4Om26s7BDoLeFb0bo5A2Vo7j8nNCYwKNeJxB9Pw/Dmhri3ceQzmdFbD2NEG8d7Uqr7zn
ffw9yZ+zAH8Yk2NYcVjigc942Y4q4lF7YpZUUjSEzLp7K2z0XgXZJkdyVJVix5NeJGkyZ5pbLje/
t/RMEaBxFbUyEklpafs9nYzUSlAKisPXj3ErjUMfgTr8XPSMT0kLoBJ2L5mxd2q+Hqy0XflxEe6W
8LDXb1sOK07AX36w8loqeDdgrm9uefiQDsNyMnDW9G8QpQ2QGyanUqmLXWqfSZ++6AgMG7H9U+zP
QkAUm8bSiWJ5dQvH8zNPpxXi9YxNH6I0LwzhtSjlkaBcHg50hOFKcYH/Z0QiBItEqp/4iqBYrg8L
LwZgOiwSJgB2/EVZODsLTJzn4W0I+Xgir0vO0f7apzMIipg8sC0bJyl8muWcJCPkH2/NOQENBbLY
S6rii5LWRTVlhM/ODFNTZkJgXhLXaTiqdxfRDOJXvBmCmQUSCQKHqD0JcpSt1NnpB8ROdGzXcKaP
DXqk7l5sm/jMhVdjCe6Mwma93uZrfELCvGJuwC/hhwLRNdvgnYSt2WYqYI8jrfwAJdfCclKbSsgF
zcMPdcChwP72nZQrLxjFkDJuRHLKvPwu2xMCfIheB3WZBz9cTkbMaM9QpKdDk56cAMY94gbF0ods
hDcOqhfBDNvqlI1V4V5RdpnFfGgFwZd3COXF/DDmG+IgE16F8dsW+udaSlZ1dY1ut7Btl3XNE+lK
ITsloSk7/NkafooM9qRraaZQaeGAqO0UCyAhfINhFoBVYGyYCXV9jNAqm6oKcEneSc49vgoH9aTT
S9aohp9qk+i3fKcaBMB+bae21Dh4YIZTNmW462l70BPnlCpCMErkShGTC8qNFTLrBif0qK2JfLeV
QXV1D6+dav2MXHeRuClEN8bg3Vnf7x5KXGMXn8c3aAe7ugtf5zeCTYP9dC/+7nGqjpqIQllS3Yme
iLjHsGASoo6hSHTVAPPVKU2EJz3cxzoeRqqiFqxbP0OarlqAcI69pfPcn539CHIRmN2YLzQzOxBy
KY4rIV/rY32RWNIlqD2YANlJ37Ww22muc6nyGb2UERA+RxijHwgHzdQR60fswbYdGmNZq9pJNEi2
Kpj3yyG/yCSboHK0SHXCg9qsJvUpIb2URPpyUbx/SuAxCn86VBFEQpx25XknyyVI/QYgE8yNVtcp
D/Y8AyC1UXDTEwgFPXmhI3n7c1jh3RGWQVNibSORlApmvayFY1PJX9dseiBOEHpbo8iUXq9yj3Yj
T2xxGqahwbPFBomD86IB5YZyRl5aCiZTIXsaBPIefUD0fmoNe5xAUlUUMe4DKXsIBPUUJNRsHQdo
xoXHpkIL7saZYvt+FqeJKE4vb2FKgV+9wlkL1+pgBfs6C1/LTOAhwnxNEl/yvuEzGaYPXvuCjjfw
7WJ6IWDa1C69yx3PMjySQZBDkhvpz3mkqD73YgQwss//xBkuckXCx/Pc+dwmlVLC5QC7ePbf9/jv
twqYKOa4MNdK5ISN6luKGVR09SBK1zXjoebf4WvNUuemhh8lNAjVjHdlFbhH8lhHZg1C0V3Tz9M6
Mxo1A5TS1SLyD4HjaEnAyU/JV9wqRUXOzsRHDFFtrAxhJQ02hFhcyRbdKO/3N1wrKeiW7Wzob8bm
Zo/Rv1mVy7hlEraz1xV8Lv+vfMPdCChm6tsaEgpYOV2MdCV5EW1uXNiEvh5imn+tOut2abo4qUOL
yVkLr8CbrTJ53TIYhRPBWlOsGU+3DGPnlGJJ2bciwfE35hcwBXFtHduoxKnrrY7uhe54RgET5c7c
QLRPwCc/cbnEcNM0HmKKepczJOMHunzALgYjdSRltf8+dKcxVkP8bXFu9jm3pOA6GEU8ZcPx0yeZ
7pBPhyHr6Vorr0q+lJuVj/qwVEgGT/5gbi85bZo63dJPHbP0sd/mLpzOUHHitFNCns1enE9slXaI
xTOwhHlNGP3Exi0fvajiGLNG4EY90nn1MDGdI9jkaZUpqWxLhXP1C1o/4yKNwZZ29PWqVMyZXOXG
ExKtQNgU4TjqwXWcAhmKR4nwFSGCvtDv9E3DLYBarWlTUmWAher3rQc8Mv0g2vNwlMUcaZl/2kC6
RlnTs1I5UyP4MCc6j81KSbCEUKRSzI8uwx88H0iJQYVTvd+htICNH09p+TsQNVCEWat+O2rmbJaW
K/WtX7Accxhv9G6c+jqAi2D6eYpBUbXjOz7TyHie71aDXOqWIiMWIx2wazdojPSKejsKWAlyhxr8
/olT7gur1acTVIy8mCkvX5Mi8C7YAW9XKOvhJT/Wyt3xsn7eQoQLhN43NKyld+/5tTCjRqVGvNAK
/Wz0qiePgPPxkcwKhkjOsFAuGLqY9RJShONGn6rUmy2B0b3Us4vWfJDeEOXewSUQew3lj5xR20Wl
IAAQ5SvDysiPLnY9nm7boRhr5XwB62gAKg5wimeqwEGUZhFX0jB7g5yCbGbSXeWxKHEUCD+yJzJL
+r8trqJ7XyKwIzl/aQUxL0K1HzSs+VDD/QEJlHMztQagtfj5/CorehqXDxxIma6/b9md+8aZ9K6d
C7edkoKbLnSHjie6CTqh/OnncKEZfJAyy3xEqcDdDOGCBsGgUj4Rh9rp/bfaknmJWTzOK7upzyMT
92wVQxHYAIz14pIoTtkd1Up6SGPE9Xflm/Bo2B5purPJtws41IGAqlbo5S+FRkNNo+uwNvSUIGBN
otqVSm4EMerdhegrLSdby1QfRl9eKbU4QNte7zlR1FUuPktuxHcA0lYkf7xiI0B+prMy2tOdl5Cb
Al2yrl2Ab43/yDlvWyzkv6pgr6oaXZjji8AbLSTDElbBRiYm3HT6IMOsRoDUAGXtpaA1JIYnHOCb
vj81yTzi/yYosOxBJOrpJq6MYu4ICXN4jE2bAJ/h8iTx083MCvWIbADd9bR8dh3i3nHcP4hPUfq/
7kKkv/ihS1/TmktAgIpzHwnT+YwrOjB/kMra5VWmEnq9fTWkyUspKIi85X+6lCl25dgX6PUiNB+w
SDHXQUxc64bL7BZ+FY8e9wroKqX3FuZvOi6WlaDBgsHBFtma9XOSlw5JIO6TK1cTyg81dzauv+uG
7unLaLd2ipF23ZnJ1G248NdpianA6ocCBDFnXO/Gv29hFHjzApGLva/4Cgv/hz8nzUi7KHzCsYiZ
YQwYaAs3BtzkiPnHQ497JrQp0C9s3kFRNX13zy7XFjlTmoxeO35Pl9HfqNGmcgNiBP3wkHimG2+d
KoJk0HgrCFcc3OjZNPtZVcWgu3TjjZS/Ye2/hX6tpdC+rL9PTlWSNAFB3LVKqkzzR7LDJ/Abr+pv
YmKx9PCT+HvkZCJ2M7gTPuNKqfM34kOsuTJchQN5G9pjavtsYvtiYlNQAcWmjoWrB6PN/E8DlRRL
T/igZZMu8RqluSlXmikLxl4IOuKiG3K/mTbRw8L1dcPYxLE8Qz1ozMD0tP2kQKdnFNQaSQGKdTvQ
4jDnLd3DpHbEwu1ziS0PLwg3A1AdcR8DdE6ilDfCBvshMSvo8+v8A23Zzz7Wby71S7v1qohx2Lyk
Abpw3jP67F98WObFxhlctzldiP51unt50N00VyA9toI2Ic5NasZWb9pk2lIOqFT3GM6ZIGQTbgoL
4eqY6JdFK/nb68cuA3j/mWuxN4U2fBo/3dXzUzuuDlI0BEILV/xtxSdkj6Wt1Rk+IEEG79nIAEz4
dqbtfa31+F6hJFRE1FPd94sHQKs3e96g5dbKs8WgiZMRJsOWP/qU7DX0byTW3vPI6/xKZKyJBBJk
KfG3hZlTIQmn8Mow9G5eym4+YWmdcKxzyBlsXfAL8mCZtylM3kgbldlRy+ztUZHyCxgWhm3dAoRY
15+VQ5thKdXnXFnfVMA/RwD1j74xfOH25t191PAxZW6fcqUkpVzMFH+pbDDWR/kInY7RTgPHO2be
dIUF6z1g79nbYrF6IIFDFxelllNS0Ewl76Rq0lVti9PcQI5VwIK7Rx77kvryLm77kMVTbX7fzvFI
C1mZLpjeceou8Biu/DvQAvLvmlv45BhUgBuMlIaBHOtAal9rx2QDmvQdi7bW/xwXjC1Y6iD7JT+B
LMdZ6LCeOmXc8YbnrpyD6lY842YEzxqHUvTsgyvQJaF4pKKA2vfy/3/CeBrJVQxDtl9ZfHzZCKz1
0CIlVDXlvI7IYoFZX2HXAMm/kjNNpV9Q+qZ+ZROTeMPDPBYE1v/B5UeZ2WxDJ5czwsmioH48SWy2
TUtbfSuUY7QfJVuR+Vo0R76MonvA1JrfaX7KaMp//sautCHfHiAgzqHBgG+9PxFJ2jZrAq/Z95o3
EOXPlOMlu1jKORlk2Cryywigqpzdq6G4S8EDJSDQAzcV9LnYHQBpaKEuILf6wKzvaMhzHCP6hQpA
GFZGu21fXb7ZqZLIXbvnPAF1t2R1EQYHnb+ZrscA0CAp5iCd8Drmrge4jvboAzem032rMS0CDaDh
Gt2CMM2cezGovuTSyEcMPCZf/UiwX3tSltViUFtVrW9DbVq6LA7zmqmyeT4u+ktBQXKJmG5qiEZT
R6M94XSkhMU6XN8j5ddectObrI68eYuH8jXOj8s+8RhaoJ24AmwJ8XeNOIgTyFyeDVF6A+JqbRhY
/acy4XasjjXCiI235ZA5lPJoZKYcQHysbuD9ParyBLiQui6e6GrG5qQXngJ2qk1QZIcMoAI7k423
UAzmVU3WaldFv86E+Io7O6DMCIpuqPbIhh14ndWuGUKzPRRCBXtxmdTziipsgm1Kel+RLkHpOpRH
F061HK+oTBMc5qTBELbGKpG0vc0vSUO7Bw5tI50AABsfj2AtuqR9e9MHjIBWlEibwY4dHJt86NzQ
OkCipfVe6ILosfvMlfryYEvo4jfSvs1k6bOt7TpvMKEa3A/yc3x8UvkYKn9qjBR9MZV4AeexdHnJ
7Eg3Rr50tV2IXa1dbC0H3nnFN1nHRQHrm/rrnd0qUOH78XTkzYzaFIh0b3+plW3dU7z8Umr4vnlt
f+NcQxLZ38tpvEaoDDdR9L4TaNtOOLj4Q925dUhTJ/bn+oMLEtnyAO+llBkumHoS3itPIH8yXt/8
4fRuduCaatltlLuoAmb9WJ/1n7y7DlFb7x0IQVZEdxuTEdxCPbclPVOjs4xOlqrKhzWS42Gsr0aT
AUVwojSQOdlnfJYQ3MIOd5TPoc+Kl3CiEqlSGa4PC9X3i8VFzxVG4hRxQKEYkDfGprnliL1/D6oU
NSZ+2oxDD5ddUf7RZQkaJoqFCxn3ZCnWCHrrwKVnTnjn24ISIl/mmNBokDg4Ln2xdjKBi2kxwKBD
eIVv8BHv3AknvyCvCLSk9dJKbZM4LHwN7LOB7VAx4XXeWqZHsIJZetmC5+24oFIU3O0t2ri68TAu
gBRGLc04OyzJLHmPbAIeNgugoS/ms1rfQfgYeUgV/C78HtrrLawC0NC9QQOTIpm5gdwh7tyIDQDC
gnpEK6UHDJeoGBwxnl5OlaapFYDZ3ySgSOtnP31/AdKALYlpI6ILTg7JFzIU6yGS791fyD2WEQTT
uFGyO2/DVsw82d66J+RFEl+EkDuJ4J2AL/WTIEsdkqI4NrNdAYn/IgyjTGMewbM/GT7/mw3fqYsJ
NfHlBbsReNPzABigRSXtygpoSThd+eh9RCka1CmV4jZfemQvIwx07NkbJYdBNfMRIvQMS9U8mSSk
H1tN7CWDMtsfNr/CI4HtCApX+u6tpkXkG07B6MXB4dIAqEI8yc+2TY2rh/ThRLxiXqnSKu6nLeob
OlaHTV7iHr8ww5e3BNoALAah2Z/BZhv/sidM805NM81Yk98kq67ZUxbCLOuwjv2PQDUswW6h3zTT
iT64gODCN7c0nc9195Ji/82t2XFo2d4I+2UeatzAXmdinzTpFXwLfhY9TTo1XVa3WxBnTmFaQISZ
SeYMOYLT3oFp8lDVHXvxbqTuQhDFPH6awcG2VdN6YDNb2fwVPQ25GNIXyKHbHDdy6OQEIJwsC3nS
MNQ2Lo5QGLXrR10KUocE8+gzdfz75tHgq9rWBxO5wDS+b9n4EGhoTD8RsytdM/YWmBn8AB4cOEL8
LauqfetT3oKK7C/LZZlRCxtfTTZ4sbZKwvay/2eSlLETXlGmhEkQuYThP1LizCCZ59TGGvfgcPN8
V5+Brch2YFZzbaNXOdVRF/qudmFBDb0+acoucwZJsd/fcYcVy5obf7xUW1pbw5F5ne137NGS23wq
Bm8qoM2hAN4362oz+12JaLEW5OqfeaCydVeFSbeWLlAJL+9mDwqx0EuPK2FuEqbnCP0GV6RaCYDJ
YI28RPtQ0AL8zD3wBEEfPHE8ApSrkbT8YX8TjeWBUyu6NkU3uwqyR7NDkQoxUC7bbS7O7HaCpWm1
hbiOj0+T0MGx+WNzQcv88yGNFxQUKl7s5h9XLleoxw3FfNqUTgBEMdzF7ztIWaZ9zejBYjRDsIjI
lQxuz+Kj+GmA71QbBvzN39rDJwAOd9jYtxAPgGVKwaFuzMBLMg1TCQm62nweW4M+Np7LkoaDC2NL
X1+Dwl7dTJuQoquvSQw7JDROLsYFjfZxPftIWLsvq8pB72gaMekkajA1YKPejSvifbmb1fWK4oc+
Jp622C0DCj2eYEzdicmeUtWjspni/iLw5ZvdrFHdOq/vTnfbC3c1ZGJwu3RX/txepPu2y94+0HeH
ReFDq+0aFpueYIGgNob9N3o8+SmuejR6Z4OSevzguxeG7cUi73A1n3y1XYD1U/tEHQmQlExYLvwd
/ne4hGD8/dAw3HTCW6BHjRCLwRlUn8PZhDoE1UlmJji8FmmQ5oKE8Hp06VTsaO/R/NYg8uppY6Mk
lFNMdkfAboFn8O30R7qG01jdzVqx5x12QctyieFs34BAoxz+/6D9FQ0PU/wxyE4qGOjzBW3Cg6Hi
42ehXX8826e/E2P44W/cd0ukDdJN0m/vBl40s6qMS1JbU6iv7Ed/OaxrXoJoly4Z++J/s/TBkYkd
pXuMiAMfBJUiJwuvF0wu4aR2J2eYfXV5cJuCiMJvWgzO9O8CG/BYZFkKVnb5vSg6mM/bRIgkJoJ6
RJOPqauaxTh8YHjSmHdvKbIRspe+Vgy8ztT0oxXjXTwmLt8e7bbAu9j32pjFNkHPZD/WY5gy+vEL
B4mp1QkM3C3+HLikqEEnvStnTS1YeqlAIKgAQ8cXdtG78db305PHys4OPyyXGjljnC+Ui/mgtD7h
zg6TjhLuT931F/+e1slDg6Om/KLwm8JmWMn3e5h7FCmTTlVGI7nZhr6rshWJJf1NS5hPhmdvPof4
5312/NmyguYt3radfBY9xdnkjRf/tz99qsghc1q59bC90sxx065vEp0I9gaU8Ea4069uTd9ZtsQH
ad469lY2IEo8Ct9+z2kO2VHjivW/0AIf6Bug+w/k+rkcVQ2Sri0C5SdDQNt0OLRubKuR1rP/wOwT
qmPL4fhfxPM90vGvQ1FaevJgqBOmMVytNEwagwENHDxNC+ZGkBBZHiu7u9ibJCXgzx2On7I6OLc+
MxDdCFKQqKufK8dzNBMqJYbfhhnTcL5KcqR+72D2svDJ08Dk4q8lAeT3I2383qtyH5NWuKvehZRx
VruW9Qay+qYwTD6YrGE+giTMJt002Y2QOLcuHGkKkzEvwH1e9a4f5bG0O4fmqR4xLLZZc9JTLyOM
EU+wsUmzG33xuj1X/BvfOqYvAkUsZNihJaI5xKB90iSj4wZai0UX+hFwWLndYGI7UvM1Yw1RiI7a
m1DQIKrZZXTMb+PUmHTVBVFXrz/cK9+1S4Bnx+CbX7Nxj+9x9S/RphDM3eoQSxG28BJEMkM04VYl
oahq3SyRSNOwnDSgXj6W10leilHyIZrhxAr1OKIZrzjoI69848Ul0TPDpgLeG6nHwVMD9dDLSrlt
tgvgHLECkjMqmaTgihtU03kmDsm2Iw90kZSIEKnXoyokl9+nFB/E9YmkW8rlwvYYOX8vZeXbFTnc
3w4mUVOmRhSOvDGNt86HxZ3AnhVerhjDvExElLi2dH48UtYVAXR1sUynJXV5+fXaWRJuT+wzWh3X
w6Z3PvpGjfaNbpJtKM07Y6Q8TZausuDCQu276Iy7Pg9SqZSKCJp75Hp87JYvatJ0zRYLNhjXZyk7
nNnIduA5jAGjVawMVlMvXAzoqDxZTfnKHdbrdhbk737j90tMlZr8WNykJYEmqwyOvSwgAvHEbsxr
Ls0DhtkYWNyHHW9L8+H55rEZUu5fTeT+Be8UkRGDKoafkwO4oerjduZ/QgdsJuiUAOghn8jLBd5K
CqCCPhuQH1rx5amKPPtpwjDPt/evn3xzG26XC0pDwDLFmGcYDs0RIwWmBn377fpf8KU+IlzPRN+g
9+wmcZi8w1AT9ewUYLZhY8yqFAJMFlzr77dsni56KAM+Ww1t4nBjTrkUhr1t+gDolbbJlbcvxn5F
TibeGMCaD1Vcx+99+gtNzRKEZIYDgZm82Ts0cFQa7iwxTz0sSt1AmMlqO+giBecA8WYZp6E8FHpn
/chkevN846l0uEK2bbyEztvzBXjnFBws7I8NB9pyx3ppSLBZ2AzhCowVEZwx872eS3vyfvJm+nq5
FZK/KhFV1jEhdlXh3C4VGYaUc00ngtk+jluiC/m00ITRWnkzV8yn7kvRPCM+0ZwIzhQFJRax7+NM
QjqyJ0DqxillQVyMl5KEJmwdZprXeR5R9MHhFUdGhnV9oYrlx0euUumwsdqmc9fGQvJXbdo44T56
fbnvNSnpyu5bcDjRKBv1YEvukONm4LcSHY2VJzyZzl5xHdk3G9/cEZNg/udPd6Tuvdf5VidBEzTm
uhhuse5UDnwKb1X1UFFZKbiSEhTotjMiTTzXi0oDwntjbo07QKaJcLWrx3q2xyNXd50FA3EjacxH
N4vjymewAJ5isw/nYzcbD9It1vG/OuLjWSIQtiWjP4qVU13tnP1kccrduG4N5P7YQKZOozsVm0mA
J7jEDR2qxUV9FwencXvWj6/kN/diFuoAMrIriXYasF9FdiQORN4jdlEPi1DLe98e3Tbu03LDzxt+
+RPHO7IAx6CMZT/tVzO4WFZ+04Sl4bm42j7lqZfLrO/P8m+uByZGv7YDAQ/N+l0n0jOQC93Kjwib
dpLc0Ny0vHXK+TT2trh91ZB2N0UWBTOPAGIwh9WThXt04O7gS4SN6+GpPd7Hi/tKhjZJFKaDNK8k
EGi5CmaBYlNseU7nxS1OwNvicwNqjFFg7QEbc/q3WYG+R8Di4A/euJsAq8yy6ZMFkGxf41vcFBGf
9Bv/EtykWVVCmsYJf7XdYY39393/yA3GJX5bf8wxckrzY0HNtZZaEnkpTfLWsjn1MV6iS2KBP13n
tyWufJTVzPUPem1PC2flnc9d5UsJNN9ZZpEhBY3kNvZzB4ueDLunA0/W6BovyBbb14cqbb2yGJEK
iG9m2O8Zh5BZUVC9vCWzCH/D+Vr0AXTdcWkV3az57hIHl912qboXe6orgnTLxb66+mq1jTnI1dWW
4ip+in0vJhi7pL9bzovvMqYMHkf9t1yBdNPaZkyObhSoiGdRXcC2aYLcfLtNgUUVtD9yEx2I3q3R
tDsFVvvGx7PLL2VPZaMHDLoKdqOoYiEsEByI2zz0LAds/EOIyeA1vXOgwHRo3ryocOtOHmez18Bj
sAHSbbEETWp6J07a8F12y6/qd4S28HLCzC99Le32wsOdxjlSuq6TRDS3tOaS/onlj9wJnENKjFKT
TkqUEijB7/8aBYegvKVFLlgP+alrpSmMGQw0gsNR5Epv6W8EJIIRrn6KYW2Vo5DcZdr7+Ij4C1E7
a6o1rrfyXncfLqDjdVMJs8CtWE60mw2idR2SURG2QRBM96w9yA5jqnt9qqF6RaCN/bBbEeyrkTeb
cXF356m7M7Hrbewy43Y8H6M9k1Qztl3GHli6c/eJEkaTg/HI7DB3AnkIZLzeQaSovpISws9sr3Qy
BLtflMwPfNAhhuKl2O3JoWmgqQNsDT1QyXMl8h9yH7n41VEtrWr/2sJdXmO6peH3P8BuSqg5j7zm
VDvp9keZB9drIyPuIC/3/+mRrO8gjN9BAXfJtKCqju/s9NtBQAz3YYMSOVFjJgqGj+toURyPM1Sv
EpAH6upswSObJan19hI63yzDAW2LjNLpa1sNv7v7flz0GukGXt1z1QGo/s33iAE53GDxoJ0s8TEU
hOsfFlPH0sAPILhi+knUNbQuCrYP2IC0gkBpTl5pMeLd62W+A5thzER7iOO0OGxkl2jivyWcvGGN
6fYDmlsvTl2+83NJAEs+oSs/jjIwjPkTqto+V4uaPxLKigspciJJz0dqGp3MXIoUD8OJr9EFfV3D
t+bf0yl+xuxxae6+mSR1nZH922gQ77ZJnCdiGulblZ2rqL6y7aEjNgI0WQqJnCs9wAMNsze++cEt
1nZfT9Z2coW7biPkymWJQexUmNv5Qx/RgMMssN2ZwuPawG54tZB+JnAkI4urJ3Z8N1eUYuH+tDlA
lQ+C64f4tLXyq4dQZf/HyZ6eid0OhfLmmJAYpHzrFXyS/15LCfx5gYzivZUzIcy1uPI1DiodKUFr
rYJYgvAznpzobTHarVXMWTHz0ObAOt0Hbo3OnwifyvIm/tSqHnLtlyZxMyN/2mGBYxT+8rcwOWOC
bF3IN2AYxUnHcNryvcoApreic3v0gLFsMNRZP8x3KM/h215q212f8PnPZfQSQy8PVvwNsHLa7Bhm
W0aWQIeis5Sd7pR+0OrC/BtaKEvE7is5h3e0SUjF5Hd2KCOAG4mB7ctrnhKMIg8cWg76SZ2alxSs
KGbA0yOo8r2idgkcU6Z7/IwLAZCLKjh9JO1QCJR15+8p27GuFDd3Cd6GXbWfDJJ7QKA+6hmNBxQZ
A4quQ3Q4//m4R7NUhw6TaMNgipqs3uQi3BmNrp0aJEWtIhYm9bGRqRCIhWq7f0suYa3+XiCT/3ai
iQ5qxajjU8mSeYBdm4XeNY88iKyUeEUlemu9+avLn4T9TcyKhnrt0hCuhaS7bEpx/4WHn5agE9hg
7UXK1KRbT2UaWvqDEA5Cvb1mPRXiOB3eOo88yuC+XtBp+Ubn65k5w680SFkqzFbUzj1rcNANyUIu
ZDpM7JEEkGxhu59J2WhRuRn4qkxr3K3/R3+P7q/Mgx9VCaeIrYiuW+4jOpu+wiwGhw02RdnWSn0H
3J5tKPti+fP2fTVDtq1Gc5DbmP4ioyCMu17aj2vezML4EvXGxTd1ZHvrUBY2NM4WKS39VooyvL/S
yTYYzUdP/Tf3Yo5JiOVdtZBGXzjQoghMi9VjHHhWYBmDAjgqG1HcgAvQYtt28qKUGzxUNIAW5EgI
QEHJ7GWBR66FaM9p1KCFTVJWBSGH7/NPowqHzuDAwL/1WHqGVxvdPcu+zEqvmARLRCuGlJXbUcGX
JLKV0+CEb69ge1hJggKdr94ldStD0BeLaDVeiltTtG5+dWNIJ5wm/Ehbi3AWAGCRPk3cVg2u0cs1
wPxLNjVfAV31dPUK/ktuX9sPa+Df3oWMtV0JTUIsLaN7UJDK/dgSpPLfLHKY2KW1mJEAMODBaZP9
6GA9eV7KFw7aB36Lu769Yf/JEaIOJyQh84eDzBYijDlGlnarr7sJLo7pmPZu8HU5tv+ICTdH+J3w
A7ijoGSFkmeDEWyxPEITibANlatCaWzp/7G+JhnhypWvmjNb+tg1iiMWlCJsSEADpgImq+RNb9rg
geaA2lVtosOFHbXmpzSAArocyBEIf2CS5zHysJgUObuVIZTa3wGzKeP8V8nE3ZroAPTOvpDoOxGN
VD6OghIAnCpbGuYP5hvZRkVMFSXPq8Bb8DHuo3UFPevQibEsVfxQNEF/YSFd44yD70whSA9MaWgi
TvxngauDeljJXDlLAIaUaNZ7TU3DXOaaVQxuxPo9Ej3VdHI7vqNlHWZY67D1B11GqdiLnSjSwM7y
lFZehlTf4wJxETugNj5cMVnQC8qyu19IUQdSC0mMhdOD13M8BExsj9zFVKDPHwMek1LQdm1h9FY3
KQcNSpee2E9jcdDWgSLm+aQUgoKPw+l3kcX6RTixi8N9ybQjzGpTMxHUBTVgFl/t/tyC3eqHB6H7
Az6K2V9e1yDT+ARZiPwt3ksUJQul7RIGTibsPT8YVM6ZJWZ6gZrlubKHZUyi+RCb1TWEZEtkAFHO
L69CEmpPaeoai/ubIN28iqgFrTapn659xgK+03hNwPPv7ujcqPg1PmABL+e+BSd944k1yTO9qHv8
0uNOPwojXK2T/OeGf9PlRCpLPCmTilq/Pr0/r6HT9x1LhKBkcbmNtQOlIoDktPfge7ED0FAqjESC
+3pTVTX/yBcEsed2lZ1eDw/J8HOVWO1vKeke5gho02inT45O/kgy3FRMdFvSCZEYSdSvxmdcMeFq
wTad7r1lNxEfRMPotHcrOS7nwUBlPmFWB4rD6EgBLTgE52TXqPR8O98ytz3D/MhDxV1V3hGgrI5+
PaEXQ4zKwKSghPhQNu27TVeLaGkzv6TgajjgImD20OY04wnMl3b4XzadnTVo6yQwtWjKKTxT3uiB
xigRLd1qLg3iXVyJ/bpwuOmVfOXGmKvvJxTW7vn/eOwHNfb3o0WFxWgxWNDS9MH0ynIZirHCCnfM
Dc0iOdaroP20EwhxWelGAnyZetRb3SSMnFwY4reGFMXNJlGpD0bK/FRUjx2yusH7UnoD2KAuHhmK
a7NQYql9AclsOf2zA1hme+Tnirnfnc006I9yYd8OIDmZXncuSp4LJBY0iIC+0oO4seA/Zw1w+XMh
xPWVLCsnRsyL+qoCXtf5E/6TS+nA68wX48/QC5Hu/l5iSR616xPTd5FjmkmsxeuvwU6yo7qO7WFI
gpZsFHBhXkPXXCBLaBbsXviT45U74tj1cHSSRFJcqc+Xt6E9Bs/9+/mKuWs2MTSYgLKiogIDr0V1
L+TnkF01tFk+VJxOeoefFnW+1ZHruDdohe/a0Nu9UbfXfzjjdfiRyaZeSl24cLnPOtAA5glzAZNA
xCgbPiBbl1FatpVmhV702f+sWaPz5hC5HagP+EbzwfPs5RJIJvZ47Bq6rQHotK5aNevDU+69NKEg
qU13wYZVuLAZ/UaTCDtvNlwRw7fB+cQjJ3S2Xwl4lXWzOeN9nJS9lb/VPuqxz44e2iqS/BQXvhrc
16Gqn4+J4FqY1b5HF3n6TgupNjtWXk91B01WP483zdNa8feaSqp4JeraDJqEPhRvIaYiaGSs/8Fk
2cz0YCk+kYA/nq/Vnfu3j4uUHkkkCLO9qMczjoQwjI9+w7PyiF+2T38zuRtr2RysmqrLgoFCRlSW
K4We/miDhaGasSsSMka6jPzYZKycSmyD8fHVYahBd4WhMb6GfkgemUtQd+9E+u6SaHaW23DrHTaV
JfTqwtUAbMDVooz2keONmYdi+2EegCxlk5DNCpIuqBDiVp7QxtlCRQExkw7Pkmz+aox6O2b3CumB
gvopnf9J2iw44Q3kaq0iyy8IWvPHfItjHfnGLnZqlL2oD7veRSwhDZTXoE1isPPNcPNp0MGUcOwU
B1DFPGKnnpDWPKqFIAtPEHIWXUcjMXUcZicZ30AoD6Al94fyOuK1naqVeUSEP16hw5s1IgqPFu1W
30SCLLCiir4ELDpFP6PW9lYhp5dBVNgUWE+xqrO5osmQf0lL7tdBV08UvdGJ88joC0L2//V/SsuF
XBvonZ9jfLfrwnnnoVaw+lrORCCtIoDRP7ruhy3tVrg6ISDIeOt6hQo4vQ2AMBSxSTnDDBpznDXQ
UWrT1LD17q18qV8HaulLyQLQ8SqI8j+pEgG30dy183GhxWlREIrYRTRj6NzAtaRfhNzKFY3fjFny
cVvPRPEew5QYKa163DR+nbI20WCoUQZjh57vWfOFxKCueGAcCtJJeGtMRShcBR6IN1IMk7Kf8Tmy
aciAgJtiPMQhqyn8KDXH1FWeGiI+tYJQzGAnxH1yFRivyKPPlhigJryjdqPkj2dPv93jQV72+Y01
m52pQOwoVEO/r7bXyHIxH9rrDjxBMBmtgpe+2fybJOUQLLEYCE6rEUUNL9USLt1C+VeZLmG/O/qT
cbOU2jSXvEh6J2X/p5egejqBiLXmSBX2KwqEFhTfZEk/oK46IGlBNbTBbgfMnpRhU+S8zO96iqSu
vPSIih0e4xXhNTb48VQH7cGPabwg0eIHbK5a/gJeuaOdHVH1BByyNsdv5Po3+9hkXkN6QWh5p1HC
x7SQPc6PfLqUBtmSjud5cB5VC6P4eV3UETtJVnjaKUhb4VXwCG63tW/8H/5Ym/l8vdnkK4U0H+aw
gtyu5/09N59hmQAJqmdfACS7A2YJ3yTcRkU/mxYvGA2kfrB9DgBAVtmrPDrLAWrn1ARgWg6eAUc6
DfWboOCBGHZlPIy7AdTGlhHO3LIaAvfuby/UhdTD8WPbxFU4goN5D2p6lzhluWLsWQBxezzfeb/7
eyCq8FWlfCDuc/2SzPG9zYMucuhU+o5tpDsnkSorSqX/3ZSBEBjHOR52yFR6NtBXadR4qKSwyBlk
KWjl/2L/+j//hRnJsJXhajS/gq6nTP5Ww8adJizi4FjcyeSSk6TIN+/CSXFbwmImLpuVvozdql5i
m+grm11Nuw5t6OCEZAo8GlGDr6gX2aw8bnh2Z/y20z7ckisZzysUUHTD4IwkXn9ZTr4o3jVvjo/q
9tVDTLs+DMBRNj8Y8OCqX4aSmBFJaY5V61pTXpH7wbM2tBsKwtoNeZB2kb3eVyXveu1PnjQB4x4L
zA7cQ813iha/GAz/f/OjJWCWz5ZNM8mIRNZDnZ9mtBkxUt0fH4RN8HJsc5m8BG9EyYtIDDNWemNf
FVsw53eVwSB22iGf42j/UG78sNtvliEBffxcSzBS7C+3l288BxdsfFmbjXFs00DMpDfsRPWXnVC0
Ofb2Tsi3I1rGUbrJeHu7PQ6vW7uINBGgYi8SgTTw47etju3iCNxhtg/NqaQy7TtBBg11k4opV9X/
6hkc5gAmkMa1jpFQ0MgPrxJrxZa7R7a+0dnw+6xnRG3Gxe9esgQopZENPeqQfDQ2sv0pDywghR42
ylZY7iMFCusruIBgmoeBEb165QwIjwy74Pntu+2Tw4xMc3gnlE5a2AZcw+P8FXx4cQ3ABVDGL07D
UMWRnaGDdmCX+0zbxrv85fecyZ0gPFV+OILB7EvPVzzPad65ejHmwMsaukPtShWVFrET+fpWkux4
L7de9XIXMHGmdkFAR4Yq8dC5z00vFgx3aao5mqNwykT+C1begogbXqfN8TPDppew4+gdapfVK3Og
MrcUtrrh5IDyWMxaqjKbO0A5jlp+ojnpNbGzd4PPnjY3lTiLGouemoIRPRLX8dFcvEbv0X7oTvpW
VtLjPq354QbIe6FiDTqh8zcgQgaxoIAAxWmzvn5L+YVvCWhsjm8eBZ4K+nS5Chf3dKjrd4UApVey
AX929XoZky5PfC8Wk5HJOrOArguBUPigQr9PAFc3yKUB0sN5Epwlg6reUiMJbpGa57F5ciR/VSt1
XmRvGB4kaQfrTXmmngxQaiSJkRNy+7xqqZDlRPoaN51sv862t8vcQ7bBHi1RlDj9BDRYk+E+T/tS
nVNxfuQF7G6VvPzRi+6L/ATLM8r7Y+NiRmmBo9TVLajAt5WQNkdpn2UX9QdoEUqUW/A6Re9g0AOq
gSHXbr1neDBRogkL0f3KyJHjbfBZnE0TafYvQ9EUL5jAZW+/cj1YswWqxJqDZ5GTEHizAeWvMAxC
qGBmhnjFHj5AceD8MX6bEETbZUOVY8QbZTKE17O3XxtxKSNfnWcxSZlsNW2aoc/OOU6tlm0lfURC
x9HOqCxL9GC7wcmtuPvEndG0Je1TKHia2Wi0oTrkIu14eUnG3z3jX43h/Y0JDlcxksG4b/+SfTeN
tyPM0wKYz5MNFFFVFSxzw8+GUjM1hYjTRaV8wA6KA0dZET1gjbhXr3qA4bFXu7LtRC9WdwDH/2sy
ksWzaXgHjVgB9376ypuDJWCZb1iGarXXQwbj0hgh32NiZm5uHQVOtbwQhRbGSwaoUA7UAMX58BvV
BeInVfNwy/nswXAzKKTVxhjO4IOIzYGCH/ZQVO1Ftsanb+AHJnMACTVC1ei4no54hp4wHXQRu4BH
QtNf+XyLtEmdeP8sfouYCNQpqn66En0580fSVAbscPk/6fSaPbUpOhm9tz71hkXExQd+msQosQe6
b0tCXwL5aww+BlG9LFfR1MSHbJ91o177BqWlEnJIrD7askRiPTXeNwbdQYSzy38AkeJzISdBkw3H
Rsw/xV+rfZ0JNkgW3sQQZJA+3NeBLviBknD+LWNFv8Iqwdqu7MVgpPgEvJWPUFixmYGp3M6ZLY4c
b4jB07iGkvaVgQhXcCGNpyzMV0H4gD94/0DWhRGoZPYY78PDP38eB21Jo8w74pSO7JDrCp1JsB8z
Bw/vmLlK9tSnXN7yisUJ9t5k9LZONq8HVDLs8OBwU5yAZWylVH4FrsU+wgTi+mtK5CoExWIoZFCT
y6rG4sVhd48efmAd+LpGBg6oE0Kflai0Im4hzWMZHWGn87Fu0H6OKVh87ZEe9Jq6Fms7Zgg7GLwy
IO9SPSC4oTY9NINKYkpEg9kby5uvGiQ1PgUfApLWcA7Nw38v7KVJmzKl7s4zMwdAKZsZaXijjCJt
5BRuKJ4p83SfUb942Ia3TNjDh08mMnJwT06lEeUwAtcNxTNEuwpi+24+Bqs3a87mnZttRluhd047
4FJuH6s/ZZ9rczXe5ezC0hCND9mcHklmtci5d9UUmDH/DEbtiX8q7PQ8epN8VUmwAaZZw1Q9R1c3
xB8HOKQOKRQ7TvNorMxM9M+W5jbsXL62s9robpCCzFz6LfrD2bxLAFp6fTOcVDhHZUpFU3L8ES2x
OFx2qpztvfjv9kaL1Ek6QP2JnRKq/4qiomgHnOZs8z/341VbdkIpwDWJVNrGXtwucg+SnsTOUUwF
6UBYogR17fH0lvOWYTVKhkeg3M3f2nXdKWn/0wtdmTXrtngtG9EMENkkfGtADmVme3MWzh3Vaom6
URjA3nkrnIpbMOKHoPHi4k7ATeROEKjD5QhbVsQ6p65k2XhAaRTRlJ9MTS5GHqfWBaAnmmWARj1v
6lktdIXYBKLtL/lPVqQbWlhm+IV40zSLCt1Z4FIFqs/SKUVf1CfYwgZIHWUVl7fs2dJk7LYE4pmH
U828ARcSjzqEaG5gwwp4IJ2TJstulgWcmBfJCypD970u3svKBzcO8z0O47iwidCDLdTlV8hlb3QX
4xxLM54T5TewO+s654M6hucnNajGKr8TBbfAyXIeLpBGCXFaPhEzN5Xn+2yy11hBzcG+LXwEWXkT
F5VklH7PyvkF++8WPV+FmQe8hkEypCZ3Lyax0FJ/4oHHDt4EV2kOxK3bj7U8xxOlwo77HEl2KE8B
oJRFKoOCSrVHYWqtj7HiWB5DvKXev5ABHK8rXwnVLPoPiBzQyyFmQpfhCQgR09tjcYVd89Pnv9xz
XNOMSBZezX5YSDzTieODI3VY7eQOg3auxLrs7WIVjyeGtQSV3oGSq2H/c1C1Em00VddI0yO410AC
Q7zmuA4ojezXrMDKr8PtNafy6TE8H/DYKisEOyp7Q6EY8HzSjUun90y16cX1B5uHee716Wv1BLTF
/5V3IAO5l4HhOUBMLb/4f60bbRHgPZXSpAWpRAXWzgH7cZk9cVdpbcJjm8mJ8JU1GvuwH+u/TxHw
cNi+haBfDH1MGTCqaHlb+qxFBxUbRn7Rb+hylpe6J8xYFxr6I0+bESbq2amwEROsdTd8JyPHGRE1
pXBHTzXM208PzGV4Zr1l9j+uusgIaLXJK7G8H/4oBhF9Q/h/G9rc7uqZF4KnEtOwTd69TmSs4qQj
Ffjbedfx4U3gQXlwY9599VNIj7aW6QrJi127NQyoEKUghrJyW98ySiY/aOQN7MaR9GoQPQOfbHQG
qS+dJoMgfvLCe3zDvaS6Q+c/zR+Rei04AStcOhkcm/TGpNyEb2e3m9aLPXzejtwY1utQL60ZMECx
BQTTQA4ufQ2+XRQn9/l4Xfz1i/2v6w705Y/wMkESRLIKuG4ZHir6on31W0EqQTHITdexjpcs+zA3
W8Q9ZO7mysYNUVu0WTGl/BI4b4akaONUQ1kWkD/e5U5CVM56lY+H4si6jpaWXperI97AsMIBrxqh
9D0ykzLIynyaw1DcIQruBCcbPtveozUqznAGdNBs3IODr7HQHwEKqIqQc3RsZ7PlkYIYJdpaBsZG
0FRyWm+ObEpfiKXAEDCMq73tpSCzWKgYTyTvWZmF3zraKhD4Rx7oY52LmLOJ+pJd/C28XMAVACtn
CAMfi0R5FmHksxdri1yLSavj+C9AunQ0jt5p3rVYqgt6YfOr5/ZU0GBUvh1Yc0Pd1OuS5WYzopQh
8MLY4/ti6BhfflO49lk9GnTwWV6M1CqpQEbGNQLMgveZ/T3KpZcupDp+1AUSUORGooyd6Y2WTPrb
w3h0AfnoSmyb+F9wQqMGIo+06NGbMj778PHv0iPjUnOgYnA/ZhwbkTZOsAntq12oQWdfa+DTHRqS
8wkXk5lDJKtrkIwnDN0jzgJ47Z0HgVzYhhPPK1QtmHfhaKSlKttTOTuMt2p+/6dBqRmvyCceLnzS
IPEctdRlmVrO0/Ppfi0cVQgoop09XUBZ01t0H6Irnid0zgYKc91O7Yn1mfZQ9eMpXikYLNOTuFMp
NpRxgp74LSGGRA36RDS6VF9iYD4znCk8uRNbaceLFzF0HsoxH4s5zol66J9BnKEhRytc6J41QQpo
iryrL153giufhYgULUF2crXeQjKAd7diSeee2Sfv2okGJwa4kGa+blK12nkb8y9ujKCvXpcacS7o
vr0BmBDgOZBLdLadStFfYI6aLJJDI7sXCv3sScGdcbek3RxcS74eGhI3pMdKSrbzXCxKFw4qxymy
Pm/9db6Yr3+OV8y5z2rShhUgZh7utsEJKD0addZHAsNSvLGe8rf0zwrscHheVxhVQvqEdhcjrPjE
uNuFFrVEvT8ITAhLnjqShTOmm8GlSeICYzLg+ShxqDwTadkVb8/0pffrKF+gzkiqFgLs0G7+KmqP
gQmwMyhkeJ3N1Z9z+yRYyzD90dpRnIQBUTOMInTXPYi/Ecp3YjT/kx4Caw0c5lC+PL1cCJlcjVTJ
cNf77tKu/Cse4vqRxC2Rxbj4uMr02YoXuLh52I0reWPSMzkhzxEObsWwxpl5EPbYJSxDgDuM4Qgj
ho5+X/dub/wJnvpsHKqAMHyUB9o18DOe4xkQodFW6MR+2epqjKe/zndozTcEBUaMp6ZIkZhh3iwc
z0AeI6A07+LwuubmMzd7KevAM4paTmdqsRbz6RdWb5o9sM+eKonL51BPkTdfKrN9xOEuXY9MGC3d
2XQGDH9stXFNu5yncFbUigeOqabjlvZQyWgf3A2dsF7E2w4mFsV34jUcjBz5/+S/ES1dIYR8jjm7
2J9CEp8oiKfR0UVEpn8pOFrwUAFF2hdtxujR0nM7LmLeFggvVMDRaguhD+Xd08Tx/XaIWLOt9GqF
ysGWSCMO5O4l/a0+hE5/mTx3ofJ7AJUau5bLthFozMJLpdq84tTj2E/bZ+WQ2/adDYOOP/mAHbnN
Z9mLZz8BnJj2nqwTGbpOUcetfayBocdma+koAZPJ3rGoqzNGKnxbYxj8ny9vPeN3f3dUa3PydsFx
ummJRTB0fmsnNK4zVnxWwcLKpwxL+w9QgVepdlrQmnArOLxDNjPnZb4QqE5RsaBPGGETwjAiqIyo
D2e7qtungwc6Y39r/0lK1OACnescNsftGnOv4kmiwO45JzA6xQeqDRbZhi9HumSqtv3BAQDDYHZ8
J6O0O5o8aZi1HmW+JdAI9JPXQ33sWwKY1XDtatGj/sqYwZAbM8cTQiSiyfWONRc57wlnfeq+MByw
naDQ0mDv1yxp8gFiNzzTZNSd89b4mRG8oYTZTXCvWp+jcb17dBZxhvrbKIYYuLkOrHc0vV75buZW
nqZgdVGrVxsgEh6ea1dGnMVlCMnWOYafPvPl84rVGTZeLpTeO2BtKCuhJmew4QlxeI1w3tv7yXDh
czxBtZtqYmckCbvgfHZy3e9Z0FMitGwMKbsK7CQeeM93cU99nyXhkXjFD6BJndty4XWwfpJzWlJ8
0A1ZpjNpselhMDO23cFhHllm0g3jsvn8l7m5RjKA86YY1t8jMH5t0zct7FfaU4NYDoujK9X5VnJu
Nc4ZRcKeeAxm2bO6A+dyprIynzQIdIJYE5tI6LshJco8CVrXhwQgV2Ky6pMFvkCPcnz52luE2Ydm
hZsPF6wBKdtsOk5UfSEcemG0dNLdI8HTPugA/RKbPhTVLEKTmCUEGZwfwCOkpX+t0qdi7orv9iRp
vKAB7preq7EkQ/xJXiaH51CibDfS4umid0gPp1sUa7e2kSbidyowui/Nn2qp5pUJSPJMRSqx6l+V
kdPqijGPOdpcU2wMeJWsPZkNhfMCB36pOkyJdulk76BHm7BUjRnGrx9hqZRBnzm51BuZo23TQ9ed
ShbBGfu8TeMVQAcA9mQN0VxOJMxUCR1hofR6RW4gXpYdmW8MiDpW4YgpMSFMeIfvhtSu8ucU5EdS
Pi6fnSK7+k2/Ymy03hMrniT3DtI+fwdy4G4rqv7SuxMoexcrf54QclOVjKfDaQa1/6/ztt+houSg
t3KDx+vIKTDHIdmN5Oyu5rJTft7pG4+mr6kSIWE8koYgm+vzmwENgjTBjcHWRacCQZ9X78bE7nKn
OZHgGMg4z82r+3k9zH5tTqwlnYz8Qg1t5zvm83F0L6HHKJKcFrxtyiYSx/4500O1IvM5ZGoso9KK
Y9CKPMEW4fNOf6XF5inaADkoIJ5BRa4nTUf8I9fcJdn7yi1XwYK5XSLw0pHORlO+K2NzMcvp2rPb
AH87CBhbn5j6P2q/6clT/t6TEJsEc013SmlGmyxbOlIwoG1P10G+gscnesVRF4IbIPKxnB1iB+Vg
zOpALBPF7ryZf2UP5rRI3zIWLUMlu9QwGxNG+xfl4MH4dgDY0AcI5LWcvHuNOI7tfQL4Od/yxVh/
oOzx8lC5VV9fQ9xWJqOxnPo5vpAtOb/gZzMvLj8KaA7CEXl5GWqKFFwaQs8wwnmEclqkyJGCEAja
+cGOcHO7lTPWNuQa7+IwM4as8sWWoSeEmu4c7CuIA5SggGyqDh2tPdLeC/OoH5UZIbrZdMzrQ7wC
ZfHxFcR1YvLNCEiW/ewALdbY70JLNmOmFlilN7dAedpueZj8qwLB6Um0EpC+2Jvcp969RI1yjkL4
DHp8lDlaAUGH3fKqgS6yHkfMyUVNYhBvP/n7NeqLYRNbYjKubLlY0Y+bOtRmAGsVSxDW+apzAmqc
pqZM5yN0yBewBwsogvZWAM1XV9wq7hfvI84amkswXBNBwYqTunMjnv8Vf9amUt0sPvDLFvwxduNO
xKp+qSBAJf9hC3u6l1xx3y75VDgzhQlbmPndjwDDjgjhRJ3QMfA4PsfP3S/uhrc0/tuelfUEdSMF
Nwtj9LpHYRc7Iz79YVb3KD90eWj42aKp46TR306SNUn7VaUIoACS9BEPJ21T+9BX8Wrz9h80OuUl
zgNvZMFFPk/fFIwzbRyaX36Rx5b568AUKQfD4bw8G3i2+xllMBf6FXjYcBb5QtwwfxmzawnIJ6VB
SU9GUFC0UUbVaO4tB5+HLu9qcF1tlHAt1s504NpsQSKp57duvauFRqDKsG5ixh5NxPoCKGiTW1kG
oFL3AZznh+XBUb0v8pQ7pi6OY2mVYuHGFKVEbBZesTfHn3YRH6ZDtsoyy0Y2FN/nFsbjWQFaJzFm
nx+yaH0RPs7FQE6FiqAg+3x9ocWrfAdOTzNJQ0Hqy6YwWOxNytoKh7y/XemQlpE/0/EqkclFPSWk
rV7itcMKPSgCnyfU0m8itEwMJj15RNsSV34q0hkqiMDlOLq62RSov0uZdfUl2bTibpKcey6GFup9
ZxgdOkIG/5sNqVpu5OXFkPtIXe/OK961DzGowAPqMnphIf/Mxf2h8MtvZ7gHKVqNOsuvtsKufI5C
qlIgeAG8vZb9zYx2px3l9MrmOwiD7zbS7pRK1xUsirggBdIe5NMtrTzO8PEsyjEaMcokQtzxju4f
iG/2pjDOB8wqFoKgqc/bCH8+Zal1C7S91KPodPQ+N6MlMcT9FIatQEiIyFpUjAFwpzEYjEB2tXjG
V+eneHuvw+qK+bZyFnMEupwbVMIgpoa1poqNmJEPpdl8O2p0b/7rO6qb2S/IcP7YRmE24n2PD4OQ
I43DJ8PqniLxcV1OaTa39LLT7hWfdFu1sXXukn7jefBB3PHaGHaCeRbfbEsxMAXRHqk19DgDPrSJ
z6ZR8mSfMuTg+sez97N6wyr43PpWD/Gqs/CHjK8UlrDLYPSs5TSAO1Ef7MI7bMxxlE6bMUxuAjzf
YJlSt16GRtWpAx8gowVHPPIcl1TRmovz3CLbTK4ckzgU5fkQCp/NHixtGIOXZKixlCbkcXBQTkCq
yvpXj+7nCA6tCCX6+UbC5I+TdSBVejO3ZfoHm0dv0TntVifvFF6002nBYjGIkKVykWn4NvzC1VwN
FwbjK9bxKAMrV7/tgMgn/jylZWLK3glFAB3VmJIvu5FMFmoKKjN8FUoNc/BSEwIwpHWkDy741e8z
GtVEPckej2pRmPukD+KpjcBl06XtJ/QYr/eMMbjYWArlIELtAib4XU+2Xw7b3C2/1I43SeqdOwbH
ZAuel6F+P/DrqaBisMRSJ3oof7S5yEr4xbqMVm+SnYS6SYiWGoECM82so3UmnR1lu8CMmU938GAD
BDff3PH+nhgn7wiUhzxgERz0KPWUa9Wsoh/Ha1osiuQse/xQzXQwdhLtEat8DKFseRUiY7b4zIzh
+CZQ0Yl9HMFyZtudxnFkDljyDtwbdTJMOvt4AEXh3tCdLcDVHc1gICsN5FlNz83nr0BomkYi/3Gl
jAWbRKzUA7TF5OVhce95ylEcLriEFfre8eLhdBYIJR09PHPKxf06vS/ltuNn0RSedya4aJTuWjRV
XVSrNXR/mD/7MWrTQ1e1cH+mxB5CMwst5wzxv9MGfKrRTafukDK1BDI2dDylSsl9qDBnPjaSemoi
CutEHkydMFQfgjobSeCgcYHKxrgPShW4bpCuG0Lv+evnmmgfe2yrcmRKWF2eXUKFcSKo5MCkGbPb
Iy2+HBlZ+hebUwzIMSTF4zj647tIFGZj6pUh6IUAgxu1P1qKjDDp8gb+5GRUxB117KfQ2ZECqz10
yK5MYOOsoUIWfm5Rnr3kj+hj3kcb5I73Dxm2KbakkzQ+5afRSZOGEagfnGbKj/a8Jc9+g/BfemVo
96Lk3ouRvQ/p0GqSjScg4l+EGpRXd1SkP+qO1qsjvgZ+GNhcFXzXBjhHGpSd/rNThAVYS425U4PP
qSGJOujFHYZKofKlbqtc3u90gzfEZjCb/y9GnAgL11N7QGPeX+Ok+7HWlqbGWqawqMHA+drXfkDW
pZAS54NizpH5EV9ykzfWxpLCztg2uYkmc/WZTMpwywqHtYYUzvOTn6FUfNV20bdi0q995L9z6M5N
Q5oqD/l03YcGMW5t2F3TnUDZZ1XjITJy+h//MhFTGwaHk9kKDQqWKbgvBJgRPG/nSjmLxzTG3/Rl
7boRPPBvg5VCgnQYMbbVDSDX6nB7zKsUAKS72aAeyFfj79HrBNnngvf6xpGzaFKAdF9Y6soK92lz
1pg5I/fBsH4FhiHMGBexp4PA+R2HfMoy9KtyCN5fu/+aMOnHdIXCXcbGCZuYD4nk37cmb5PABTSq
ytuEz1yPgCMUyfB/AjTzR+KJVzYbXUKPQqV/hrV5bCKCj1nS7O5RlTbbLgpO+9ufZNNy8PynoeQh
Pt6dfckljVvC2BHyGmlr/GHM9IRwOccRrJt9fnR2na7I+fBHxxQFsKzx0Ix6zr7Pkr9/oMphwuC/
+ewtNRinwheyX+8OOq2LG5nGvfszTmwAMKvCJndxWHyZ3H0zcS+wQH3BrtORFN3XdZ2Nrx9sYzJQ
ml3GUV8tlT6lhtvxOGcvhHKKUkcSxQkwjzn6BX6NUMmpRFDQyBJ22MKf4oPjy0jORhVdOOe6Mf1r
hOKPvdPCB1fxIomDC0igdxGdJoEuvawSXTVuttp6tdqzvIugRbyYV0tvo9Ojiu4UHisMhDo/yFL2
I2yocK7CUgMSZFF7u9ku6YTTnNm4Jjd1hKvvOsBKKTto+qhXvBB5hofuy7iOgITjgbdoZcVb8VYV
wMDl3Q3Advyx5SE0vwV9+c0ZHXp+d1a34aX7mDRWcxb9Y+ESk6O8c85cUjtyMxDum4mO+I+/SJbR
FboK54CHgV933HS46M3aelmRNx3aGxHA6inYHWCrqNBEHVzcD11im3kcIq9Q0OicoLMAfYoofFzC
4AdyeLCy7WvnHwjPmDFNF/tNqFY3JxZ7Vgv+whcYEM7gT5y0dtVoEgnbKYIKjAhD5D+sozt6O1pg
E1VSorlObgnPdp232DrIJ4xDkf4pF2iwNXKJA1aWElbjO1VzNzwdWnag8rzMlFMsZvO7ND+grPWZ
B6VP7whN0692td6ijy+dEPqwIn8bvFEJINgApcrgQ6CdCTPrS6MthiyNQRlAakufFy5jySGv6buR
nCE28phoa96rZ1AgvoGflEM/x1OoklYo8Wg36Iipt8vxiGd+iSgBIMtO1b5gtg9WKZE20hRwGOUs
SUGWzfTceEe5b3QWMcXF0Z21PbzHqDwE1znpSC2Unh8Vy1aCzsnyR9WnKz1Ijp7MrR+HdGHnycwZ
3tF0qugRwvIR8goRTeijCtc/3HD9a41XbBeMxbGxnTrW+tJfpGoaDHZ8NU3qQMGG4/lnY6j/pMD6
CiMNPrVAY2FUPIUPCDK0reHOIT0BcVD8yPrwCk6NGg+5zaoFrA6D6/qmK0Mxq/veH+05nXvtfBqG
dAYPFsK1IenG2VgYrRgE5Edvufu86/aKs0tqH10LFak/O9NmMBDDq4CXHfUcUMQg+sAvJZTtJF78
o0xmXFI6G2IPB6k53fgI83iPCM/o0pMVqxPwbmWx0ls0oibQ1wYckopxCka6slXsuF2gSK2IhgZP
Wv2t3t9GLZjhFj8PKYJDZwJHdNu1sXz0eX3Z6KLzfxjw0fHlbTP0SOi0LTFD8c5zPPr/S9hk4QHj
n2bSQ2LsyQ1GNcR12t4VBWxbu+a6LBKP9Y/B7hH4VG1b/6S/kFOv33+DGpf3cAqa74Y9V97It/40
memIuQZyRw/jq05aHwHMDjsTR/4NMrhvjUS0l+mogZEpGvcQm1fGS/xHYEzJkMDarqP0V2kYA87s
hb7UlIFxnIuwTYxCh75EZC2Hny9k4aP0bHQXFdsBA6sBUCNARGLpHAWouzMba36yAte8ka4gGEv4
Itlvf03NsvOKoKSIyovLfLBwa+AiZlx7BDR+eC3aPMooxqyqPq5YUD8iO6k1EH83RE7LmHejPGkZ
/N4sgfQ38ivQuMkZEbkDs5EFKF5fiSlzLF5rV93BQnBuGOdvf22TCheATmkqCc3KSz6WXRyRJ3Nt
g0plnQHuSfu4shRdhkeCyHjme3cRHUoyTf1ttsJ17H87NaQRFH/brczbQlmy6MJ1+beOzqZri/ZW
sU0rKq4bNCQnWDAqTvbazXXJx+FFehTZG6YCfe7hivqAb+vtPsq4ARLuwT6x98YsopTVDIO01iRq
13l9k0o4izE2JFLQzegXlhD3bNZthSbONKgKxUtRhgqpttcm9e3nH+ynN1MspBlurtMEnMDBatF8
I2E7imvvSutK47pgxJgRXyT7ztEczJNKAbCk26F94m13wH9XmDwHYM2JCZaYziPDkVr+DGs4CzfC
hSGLHa4hHUOSZ9W08VxbCpsXs/kPsO/7QlWeGvvp/rDwNYzpPdoGeVmvuac+NHUvT9eASdcwEOjt
7HbteRMNXwo5zX5HurLokk3GH2CQyLHyZiFbrjPoZp8TSD1cJBf03/EMNCFD+gyCD/WFHztzWjrf
7sgOVClRk82cINlWE/youymxjEClGa51fn4NjKU0eBUYZp2xr3aJLsFkd/kyXneiBgtcKQc3air7
0703KSP9fITEPmcl+zuVrOc+vCzs4EW2v8GnamiWLOIGozujnXNnBTsQTVUX4wq05G+fTMZz6Z7T
TVqCDUYHwzUdobedFJKp6weNrAI+DCoMDfaHysW7IbUg7toOAdnKCyBmwHPKn/OmcYbsADPPWjzR
GGnHPTR1yasTGu0aDbWVwVAObAuCzJ/pXgAWOSmL3RGYsO3h+gOTng13oN7yFNBGTQqGgeyri62f
Lz/bjwhVW6zGJCyX43/vfwTv5TMQwI8xU0ZyoEhnWdrTZaZ3U9FpoEvCFC0ECq4UxuaNBYqYu+q/
j4MwPM9+hBYhSgWRaBAvlR8QDqFArSjGKZMtwg+YJ/6KoDo4jCvJ5tr8g4dfheOtKRZu4OYVFhcX
3EqPSAv2p4EA6yEQVgdYFFC1mdGTnxo7A68WZw3Dxmw0baZz0bJfDDHE3vOUkTHOuEUF1ipgQqO/
BMfhXj3MZrqlNDr14fE92+HiBcdKEvGMW2Tp5HR9RB2H1Jmo7tu4Ntcmi19cohOaHi0oDGP8Y10z
fXAjG+zpyseN+trC+rOZ6Jpt/lrwyRE949YhZIX4uBBOYm8WCMrad2TpgdIYIzCOyjsDbAZ0BPBV
KfYEZISzPYBNZ5MSsEygfwj7AgxUNaiIK3jWmPnobhJ4l22LIIXW6tL45xheY9okH/bGJvVfQYb9
82Hj+ojdo8WkBK4/+O180SNSB0+lFCXr+UR92QyuuvWCpR+WsJRpUsX0KJsjNgNjfSzQ/cojAEDe
w0AHMJZdrjXmbRPi/V1Og9Xl3fPbyBQzPtP8EUgxap/YXlQFGKGXK4GfRar+L/58zCVgurwWo4EJ
ojtbn8YNg1/DKLfi5kfH76xWkISHyhYJVAyD3TNQsD5rvDTlYjzRu5UTvApDNtt8dm9ohA/Cclc9
e7v+yrPnpn9qGRb9Ak02dbAKWe0HBhWFmWI77PeCjnu+eFlSzQWBkaW1TKNm6GMtEPKATRirgjvF
tBoeQdkwlhmqk2b0i7ugEzc2LuKa8mZO4oQxC+tWdrtXTkQXnxhGCt2ubI0rtScY8u2AjQQv5ZcA
jHVNH3nNlRiVytHZBZEYPgjdwWRFV+YNAGicAJXEzkKu6wuaoILRUifjfMkr9kDtct2h3tKbHje2
tLSKVfnIL6bu+12ykZ6Ghz7v2CAa/DTvv8QSItClok0Lf9X3dSZd8QsD3JHAEeQyiKtOnjKhoE5R
7wS8zSYw0vxRty4Jo3ewFyt0TwHqUW9RcknDW+Ca2EOmHlAowGxRSj9MHdi/KIGL2kkFGMNV2FVi
Gzwn2BarJvt7UyErv/JqDteLZ3dEu4LA4LiW1C8sUxMH8ZDrZOKCX/P/tbC2fEkB3T3HhyT8XG0y
fUtr0FX7fn2EruN/gPuSAXZa7BBqKBrqmVSBQ2XNHoHR7h6kOg1VoyYQtbZl5RxfjdtpUYqTrxee
4UGOOiwWuOszcpj8qHJGVfn8Nps2aLRRiOXQgmTxQCA1Kb9kZipEtouTLQ8n+cecuFDsJ5Z5cUku
ssjWrA08vXrljwKb3GMMMzT+6s9K2z8UtsrmN/rD6/ovTfYX1s3hfgocOT63YOFJrGO4dMklCRBg
7Lqvte/OMGy6l8eckxOGrRI6K9WKA01EwBCPUWRCA22ZPvFNkmERFAJhQV1G70L2mdd6iNExHWN+
0bQo58sWfRGpgbI3n4qXSIVdDbDu+k4YsFM+o0c09PNnFttvAfvn6Axu9zfmQwxm60fW+m93Alm5
+EtVOiQFHebmOWmKGLs4kaxR6PC1l8BUsR8AUaG3+6G1GTB6kWVL3bub4vQYqHswNj84znZZjW4E
0mLROxnTIO7N8PuWs+wuIBqQ51F2FtO1s1FQ1DF3rqKEkY0/UHwx20msjt6YvYkvhsxUqpBcATrp
Mn9xpG/Bw4FZWBJ353V3bzd/2HYW1O9boVId/hPHG+9egY1Op414feHmw4z875WYVVzKLPOZRj5r
8p8qY4jRpI3oMklPzgRyFt3V4MtGB57yHRLlWEiZm6tqPiMTrDTIfxA93HL0pRyrM//XSAwVQwto
ERdAl2j3fQUBt/Q3I8sOf+F8Zx9ZFDW55oLUiFMMP08QqQn9Wq/4D/oNlaNLAl+wCertSLIcr237
rilFCjEbjSwX1T9Qr7Q5qTFdeL0PuvR6Qd9uHrOYlboxREdmYy8OEOg07Z+7DEsDcHdPmiL5ZeSt
Snz6m8nO16lQowyzxT/kRAIFllmRK9ivcOkICX+vAq0T0UqsmKXWFjLTAXryAQHCl6LgmyKF44Q1
v8YCiEQFyE6gBlPE1grF/kfO+bcG/MJjSf0hLQdP+T+ZuHRIVT7ogwajlsIvAH4mfgNd3hJ9qZf+
ZqC9re7UmDNhehBvZSxmcuh45HSftUozfE/teaLiDEv0sbWNj9RPUCqaQ3JfjtPh2MS5BMWOTm4X
QCFheR1wwLZpHazencjKZKtxjrBjlNbv9txQWrcuQIVVB/8gphE8afAD4z6wM4gIVRmsNoVkjVLo
keLOjyVOf4TNCj36OOfq61R3VKUr6F5z5OLOOQhzLnyXh5zQPMM0XW3seWnjPrHKpKCE1lgGNBzT
we6JVOSB8S3V9N48zHKNZMpIIrnLPi3mZogUKpriQh7HHdi/ryLHoH9rHCocSfQ/CNxY7KLs04e3
3QJ9MDixngXwt3+4EF0EF4XXQAI/Xn85kD2qIvGK+XYqkM0EAN6PJzUkOG8PQWUrUB6pODcSrcqu
TmcpuopAKuS6GbpXn56lrmsrByhRKeCXvM0iyDdzXVpBpxvYjjJvyrK8ctgtf0G8KWwSTrWAc8lE
EMtJ4ARByz6D/x8RQuy4CnS7EoAMqwts2PUWFb4m2WrQNjlRwWYitmQyPpocHEDY8OdVgK4Y8suj
qu/C/nzP5jihwebuOksxiDYjYjMfCJwOBlbBKG/b3mqday7j2h5xr6blzAROy9Egw5IyvsuqU8gP
NU1Sw+o+8Rrl1YnBmK2MAE1wYEuVKL2MzJtad+33Gv6jo1s7UHEUJM4vCB/kwh0qZFOha/61vHhs
JZBxPfBLsl1ocASPEKGi/1WprzkHje12rx6lX7xOd2fe5dx7xIdiuelHpxnjV/XEIO7lwOFhX4Uq
dfWkTcA4ez6phjwxCdwH3TGF7gj+L7CXUYWHfGRtSeB4vTbR8PsJMbBbqyuljN0fSzNOBlVbbyO9
rqqeUCVLGQy8PeGk1VVQuhTRGOqcyh963P76TgklAUhhYHW+7AMfYs9mW/SVjDIxO7XsFgPP1zoF
jegXfPKaajNwCwMx7qYXlaGJi5JQ8uqKGNLu2zbbvZGgdYHlOnE24B1gnLHFLXMdpQArMgcLQPE+
zkR7F3PJuIvgkcm/9xXfs5AzfO457v0MrXs4fi558zdA38EQ8YlTMPmRODWfWgBzG0BiUqOdPfYd
oWa5KyfgnRKkg2r5vVbnad05KkMdkbrPA8L6GV682KRg3hA95FYdLy/Y9fDly2ySk/SDRWUWYQPs
khDu/Yrw48ZM3JgQzCM834brjpDjXj2ufyBU+LElYRE1StkkxlBTyd6trFqXghLTUt9KgmIM9LVr
BPHL+cdMVRsi5zoHAlhxdkuLRo6nIV6LQArq1Ul9JuZ+2bBqhItT7/zgmXhtUZIWxgSyFEcLKQpz
Ab0QTAXIVFESpDhwov+4YlKNtnfruk+B0zmZKjqhTjTdWQX+SIoyRqjldcn9uW8LGfUPt9Ijs8pn
kNhCLn5S4QLa3CYd7UB4c7cAQ0XjtAPKNw03NJi5OFcoMiCgxaDqmpW4ft7B0do6ck/X/mhxuqMX
cPeq53Cr2rNm8Es3Y6Uo89q58b8rU3zElZG5hHe71JxieK1P/2T1NbVO2Q5eWkIbxnB6XNNT41bv
j2K0loX3x/J3LrPVoIoLpWGCrStbNxq/I4LX//EWtSFh/PL2Spf/tO9FvgEaAZBuIRMbHN6Cqf2X
R9fgS2lFHJyCbr5HAGNp0oFeSf8VE18i3zYngrsl9a88xbsMcjwhbQKr2ty2bvrz7nlUVzFv0gf2
nNmj8YwDV1a3ioywKkPiblfZVhUxeXquZxjnVJhGDHHskWcfTcO1ixPkT4X4GLVlhfNUwbR+H2c9
JQisSinPQINSKbLev1TqAgqwLO7zmosX50uYGyDlhticqwbFzFCsd+gCUtaiqSAPglUYCPuptMx/
q2sDDJ4x5GyvYRmZVNVToWvSGt8rYA/kWcNph+gqNbgAW0jmXbdwFOMKOrl9Pmez49AcUH53oi5G
gjzgJT9EK1uxAdmCnyFobC1feD6scc6ff54t6X1tg1JTWCvOcqn6knf8E9Sy/qZv9/6FY1I1zh+Y
xGhLbgoO89YIhfrlvdCKD2GW4u7r6BgDjHYMBbE9cFJEPxDkHHORIKYkUkclU5cgW3/Yz807P42o
zsppw+u8Ur9bLyDOMwQlhKgLEbFl/WPfLqbWm3xXhh9i1Kn06I3awPi7VAXop26qM+dvMn/zRR8Y
ACDs6ixm/jeT9hsdc/MQUPs7JE1Y5859e+A0d+BQZR8wNQnQjIg0GRsg34zft0iIw7G6dimkd4hI
UYz7Bj1b9nrtfC3dYsTO7MLpA255ilRKAVLP37BA/CoAlKG9my0qzvNfzdi+Tt3fsyLjtaNpiyyP
Axy1Pk5Wtq8KNjmCY9yRBojrMCyyPSK+YdYVP/zYRIr83A9bbDhBBEmPBKVlyHHlO+8+4MvrfuIi
Th5emw0xBM5iBvoF9gZy6Df7lZFt1YYj4S5T6ndnr6opxJRkOeYggh+AdsKqLlEBAVII0nzYGEbp
hjUMZ3WXhYc82+1HHZVhTPY+k4GzJ6sd3FYAePchXqu6NSeU8REzJ8IZYS9BIfpfOqpDnF8euztU
7uX87NfIhmbbjOT2t85aeo5j8nGuTxRyWpZv5GuWZ9xUG1vzgGgtdYtsSmtQ6ouKrqOiucK3hy2f
IazvVWJzLI69xtqNGc4b/BaEHlutu3wot/P0R4fAtKE2yimPNiTOgQZ5fpZQHCu3be4XS6KWFF/r
YRJ9hq7qF2fie7cUF5WmzmPkqrWa5o8QSomC6AoT78sdN432w1I+PgE8Jy8SLRwbUUyo6BcVqxaG
tAz6WEefED+ATZlWcS3sZ4VU/9k3LiX0UwTfC6FudEVvMYzLME/1qtdizQ8/U/kH0d/qzrZEkrVk
TKVJ2dnbmQUSMpCMH1oxHrst68oxK2XmaE5DZPilEtdbrKmK7LnK7yNPTclveKBrKkwbGUSJ7ADv
ukR0dT02zNSfkNTAHYKHofEV0zJlK/Gt+Z4oc6eSMJxZHIWTIS4REwCIER5dxRs68IjmBzTutIfQ
2hIg1wy0SAIwdQ9ZpJnI70AMuitld2A1GTlFyy3BxvpdCrjQdXd7mxrUeC8GYVWYwzVq7TRudIKt
dNpxft6tyHBSvFylQwmEYMesS96zchDSYjdAGVoHH9PpnlJme18WfiXHj+54JlGBqwylGkZT0qlL
E/ACS6xb5Ol3XxHtI67pmIKjXSGaXxWxBtE3k0fhog8Vi/eP/gZLOycHlzb6LZEt1uv5uUIihg5V
AcRiPN2RPjPJhaxzm51yvu22TbNqOZZkbYt3bQtecZBxCVyyJdu6jm1FiDowNhN4Is18nO4nbnQo
jPnTypR8Culz0/6txu24tf9sXU6GyAPV2iUOpdhnK99a5b/X1PPqfoqQNyoMDl0BsxPhyB4NE4aj
c0j8ZjKn8+YWpOlBbdzG7ml6xEcGlXeRaNaFLayNvPwYQYpRgdaRvCTYpjWmVgeV4zIEaH1vYCNZ
+kiROsKIzEY62y1p1PaBhdWnlLL9LhPr+wl/qXG87CARbzIIf7DwnEu6I82BlvZcCKZA19asFWWu
xKxnu+kO9LRgIVx2FcEdpgjIMIKuJargEzQTk+IEkYyfMJeF0R+8lwatvWkotFEI4x7uEZpZ1Hs3
ujRoX00T1Ihjb00d8yvxOxnAFZu0XYN97u46nQaBxPEBGcbVQE3Kyff487vyYGOrQTWPL7Gwm8NV
GXVPgS5yKlnstCFg5/QnaGUZJ8eOE+/w9sipB50dlqV5YcOLO/YOZN4MALxU0K7wRNGcKYjmCZld
IhJkjMAhfbLgIMMGhuV94kkMzZGjGiedyk+xQX6wfyKRosV12sUohLb98/s6e1dbnF9dLbcUBCFo
j0LY/aswVWivq5QDAiHYcOcNa6DmO8B1innnoo+IL6350ZGoa2Oiix0xEI7Gu6De4lA7wFccpsf/
u/hdiRQ/I0dTWRcTr+diGDTWSK2DlCRv+CPqOOpGpxAXOcNuXFsB/160ol7kufQj+2kRccsH8PcO
O+QtbbImRAWTnWseJ74iNJmjPEwq8nARWj8yxGLG/xjFKkkJigH1pw7ddvoa5pzKWpmqmS4e39+9
FwUXV3Jy/ct3hjxbdUEb8hy/J3mUJ13oXYuiqVxiSKlhILHZ+mtlw8cpUUuPnERY4mYxNW4vSGx5
Hh/TZeWyik8XF4qi2gF9N/A5hUkUreFQHM7rYoewl3u9+I5OjMJtp3RfMTv3J7j3fWPgKeZUCHp2
7hP9mN47I/Y+Ir8TbrHoZrUPPxjb1ht1ti601oXZDBZK8CYIrB3AL/n23ttr6RG/amro8wMR8EWW
Vack+g37W0fdFGsP/8wYbmf8+k2m15y8LmY/A8zB0eA2z9BCC2rlELWyDVA+S/X1GNjXvjXNjT/H
LJU9YS1OR85Ni8SN7C0XLEd3i7ApawcGKakPxzChRiFyllIfj3zmgUkEwuAPMt2AKIiiP8isRGR1
KMZrRhV5RaGfrl5mI/mPpRAyd5VKDED3Ma62xw3uZ2b7JctWLrIe7oMuq0ZXIY6NfkBvhzgxULwV
dJy2yPcQkFadnsDDzUJKDupoi6FFEpt42RLSud96EAp+siboZLALQT4GYpo1NOwVKNxeTpB0hgwk
8Q7cAmyV8rKT0oWbeoz4XEZ0fFCq+NVTaOa//dSurJ4nIBm4s5BoQxqDUN19/NvStJKCd2etBk33
tl/kPA+GUHjuZgrR/uJlnaQSZbNViPm8E/IFSC8cH8vSAN1udNYxif+FXLFgQAmbOmoyFvjOgJDk
ZJtBkLdWyXA/tGpnM1OSoraRspTlg6cqr5Lghna0Gvgbl6k067sc9CVu5ztzmb6W2etMt8Xaa9iI
wjqOsLOFMQfzwxE9JZ4jT5ck/43npweMHRo/S45Qx5RmZQzSclPxRxaAYrwkc4wJ7b/aLlVYTq+H
TBGvv6cDQAhRaLMEv/N2XUJxY0K625/FdfN8x4CvzpbXwHryyf3FJeTNZlA1Nu/JGVbeY0BjlpL+
vpkoWEvfj62uEz+K+jq7jaPzVwfs5ep4yeIn3WZ8sM8RDK8EVuK00MSO4f3Jsu4I015tovLe0yzc
z65ZWHW/ss6OubxA2GLutG6PVmv0Cxz8sXpROC3kvnFI4TDvoETDiJMIBVNRloA1Tfq1NPV0Pnw0
vF5wIT94PTdYynr/FZMMsZAXcpsvvCl2qfUuNCQ/PIaSqffy/MEc93e1SDu3r6l6Y0GdsPjc+Kiz
1vH+6gyHUepCYHs6EWZQFeRr/iktvekEtN5Xe1mCdqsmsuug9s6RL8hEr/oDVxAtTwFHNhzofdYD
HROi08cLLaPOeT//zlJ8dRicEs5zhFRulBXRHdO+21Act3mq7cd3+VMS4zox25poHVrxrZwsQJeY
cHBYt0FHDJ0QeSIJAblhWwPabqz/71oUm1Yxg9LTFwAckzowckJ8QfwVOHW5bNim4LnZU20iUXLj
5Wz25bo7cXCZusiL/tqCQDRk/w9kYwrtFNhA19eWLChOwyP+t9qri27Dm2qZ2U5qh8ryV0CtiLSC
Fs8RFpbX4IakNSKkzqEdVlNopOWx0TF1snEyB38QLrRClwfCmjDH0JrzyjofLE2zBwTT8kvllpmc
jDBZBE8N0FUfL9f3pHg6S7WQZeKaV0XzJXGfll5lpbO+1wfp9zpBUJhnxeUlCpRxjubLamTb5OWh
7ao+YmxXUvok9zs5fqJCodtKtJOUyFblBpx0HLiRIPQ4E5DIouHh/IpUUWK/L3B6ofiGknSGzwzU
QABpc12oiZkoVatJ9uQy4sbKQAY5tymul+sIZFp1K2na/uzk5tLyQKlvMFoSeELuz+Wa5UVyuWyz
tN9RZT1KAci8yuLQgqeXsEMxzH+aKLdiXZ+QdgOdBj7TG53+e/imY3GQRuBJyFx8zBBxesjO2Tz1
sy8M7f8cK9DhulvpwUMbLVJlCs+H4lbGqU9vzX4Zt7yFbsSE8u7xtSoM/WZ7yOACWr0PiYb6ry/S
vLUPioZ6hs2BNuk/LN03fbNk0T7l2uRxXwgzZX8AZR4s2kSOP280+/NkEoUCEKkSz5jU3Q76w22K
KPFALB4LmLlUHgdoCO3DIo80pfBVui4IdmW9VuBFD4ehSdswaOda3wzdgwYX+nItKBjmHpKdWxcM
dIm65yRdn/SHWTFGK0qHQuwZeB8L+jxruqduovD3hQcxuA9QdDqIW7g3LvhZlfrQuiNka3CSJ5zP
lslunK9rsBk9IbxvlMyoq1xcHgq3N5hE0b7uAPUOmeQr3BWPVP68HzWlsSq+IPuV37hCZ74dmwHZ
iEJ3T8RoG922StzLTrYYyo312sKgTRqxDZO69SQjd/XEH2JaRqqnXm88OjGBBGh9RqKwMr6cd0xU
dpptjt+fHMWpBhOJjS1vcw5M44D8x4Z0KdIrP/kN8cZVsSoKWtKpMT3emYrl7m8EkfmCOKU5gVjm
8aF1kT7Fc2a5Q9qEU82a3Hb/9eJ8z9C34ww2TcIOXXeupu9wSrk4elHE707+7fZTqh0wbI9uxQQw
XLwHb5Fy5RK3jZBcz4ukKGcBqx+F8R98oBoPl6JaRlROLd8tJba4A+KN8HTL0VPiR32BqvF8nc64
P9j8zK/cGpp3uRUyazZDpDGFQ3Qfhy2VrOjScaHqCgvQMANvSIPov2i5eAsUb6MbFu/AGie1Nzc4
BlkaJmmq1J09h58VDmtzh7+tmC/p8sqk/+jJQZiMiu0dqBeRwZhMYBEcMCMZu5dKOKZfBcUdmaBT
NFd8sZf4nmdrZXfVKaBXAQOTBMFuai+GkA6k3/CQ4rBNff4idITDjjuuTIdGYG1pZPO2Nbg3MK17
FB/P1FlZYZGkkpOqgDkaqoOMy/RCRrfXtmmGM4HHuOX7dwCBmyGOt4sj1HfpTZWLGJ9kMPe1blqB
wMpv1fgvTN3zzYvt8MzsN58qeDp4VA2oC/TDeSuGt5ENydrRou4Qk3zg62u2msCde3Hfz+KmGlqg
5hIfkjKB6Ma7z6BkjFNSygtArVBk/F+B/TYA0orRd/l/yWmhrwjPy8lwZ+W05xHtX3XQgUZOUosh
CUltwqBf3mFDbG5xjn0hMwi08y/lWJRjH4OyMC6r8JlniuPppnEHkW8x+4KiPzAWNeXwSkodax+A
/0Su4W6SpuDRtw5OQbAVfl0AehBelCuuWunflyxMeCUVaWDWlor4picwhGWlt8gvba0V+2hZM3kG
Rs8rV4QErFrpzlPwFZQpX5yM7yNKwPcQq2ESWHJOFWNGaXRHoaIyeUf4610pSJuOsXFkaIz0g1R+
D69llz3Fy/it0mjAZG9H85hFW7vidMOqrUVsmdmMy6a0BOdYwhRgl97EmzWxpF1WWVztvdLva10S
xrgBL/4G0rOPME8Blqsty8hfUWky37g1ytNA8AqjWIH8AL6dRq5znTl3XwihdCOA/bvXW/LzCAW2
T+aQ/4BG1RtThQRhksdHJBL2TRiAxKlTwrvN8T0yBALAs39e4XqLSc6HBlEniEGF9ydFfDioF58f
LYdv/4ZNAp/T29QthMwbe8LE5MsBGjrYHVzYLC6AhEEVWmOFxbR9m6AFsCkZsiFwXUuklY4ZvTYg
knfw0xnuSRJkUMH/+WLMLK5Yng73CwyeenEBO6tQLVb69ixgkNDhT/zjd6o69l5TRJ6iVP34G88O
ppwj1eIdagegXuq1oFdbBL0N20n+TT5EHgrTpGnoMdf1RzNTBYNN2y19rk7l0FdKjJxbykq4Saq2
5iFMdOuCyf2Du1rKpkU1u6ZNfcyTVOO847LHJjAUOBSoJWRBcl91RdzfI37Ms7Y+Y+RyPh/ziCjr
X35BOw6glsKF/h/XBLqcMzIfCR18eFyhgYN9XQWHoPjzYSjFwtq9GRxpVDocArdTMvKl/c4tHrgO
melPYwVR+lbFJTENIPMcHvODxFuYM5Kh929Ycy0KNSKEmUV8ZrP2veqcAgK2tA+oVvUHp9xTYUrU
pElCPwwr1J4x9WzVEfhuqNL3fKOgaEnsswuqkOnv6gYqm2SBCpp7RUgjoVKK0rDZYZ+R7UHSZeqh
3NY8eyhPymzfF/a/ESHyb3YV+LX4ctKl0pKypXDIpVuFynU6bpwiXfC8XuAkcZtWkSG0QihC+ZIv
vU75jO33qjvhclTb1AUwnN2Bx+dG5poYRVAkSTlIJoNUn6D1IEaXT0LIALXoM54NyIHaTM1p7b5e
s35y2tc7d/LdLYoNb1hMt3vtle/fzSoPmXNKrBJG/bwH2LMNQHb85JsgxP9fuCCOouMv7IDZQBiJ
iZzmUcIiw19fZHGQ85C8m5kgdMSvOgRdIycjNUfKN0H6ut27JNc98vzaWSuajCkPdyEhw3+aVYzJ
q8iNObc/m6sdL5Aqs4kRjrjVuumxZocefe6Tp9HdE5+/5IYkWetFxo/xPaYxpc1ESIR2rtbrxwYe
VlJ6cUML/mkFP5E05FZOvlSL8soHTDyOzT9V7rgj2HnzI1trBIEH6dkq1StHEz56Ici+uxcUnNWH
Rke1DLOIS9C4XLAfv67IQOXg1xi9mFTkYLldd5NV77QLJdMZlLADb9cBnSLtqvYbIxS1GiEJp/Zt
QL3c/JP7MLNw8W6lg0b7Ikg3wHZrdpuP2pf5h9JKhGvJZ8vQRNY6ALHaf48CBsDTFz11jnERONYp
XjbsAUgWYAOAEuvaWulLeYuI4swT1CGV1CllNnGLqGcfHIgxr9UxuFkrHEkAzhvcAQ2WKwPaxDe9
NMU5FsXEl4AytrXAsjChdJHQqYkc0Asvlgi9mqNMU5ssWIJG85lZRTFL+2eo7dLLVF91U+WFpuyb
to0R3tlKH5tWd+57aFLZjPx4aSLfKE4zDJ3EnsboaVyyvz4Dq5Fj/2pxG9nr/IxthKYWtUuUHdpD
mvYj5eUV48Taq+34xdYPMf7FOTaZ6PgmsJEHGanlm0hihcwuhafv4CPtM+zx5o0Zv36pZ+nJebD0
IEaHM0ETR9oL3lxt9G10nU8VYHRSqWFQ+sUeh0D9fVmPv5n+DtpcUzrO2PkUKJbQAofujtiemohx
Eikg1aKNxnGLaCRUyc+uW62Zsm/05lGlq7CBr0/qSETvH6CAIIalLKEiESUzlglm2zMpM6z0wf3B
Li6/LG+d/bJWncL7ees2DerMbDPSPCcmxt4o4Yjvrv1YNd7UWgnTIfVkE05jsVZg4hcuJ88prQna
grIzwefcglv+J5sOgLIc6CTSPu9Bqt52a+r697Kli5pnxqteDOD6tDW1uSvHxpeq7ARfR5+FWdGI
p4EUc3jkk0Y+7Q5SIMsO1xCqFCx8ABJRiznMfznZd3Ur2ZPhbL9mAFYzK3EYI1NaD1xHusIxkHG1
Eu594IwtFEKuCHm8/nQR96JVTTLYF8m7mzkdjIwXE1t4YpxXuLiG1ndwxwFo7j2kbsyEwBNTpRUY
9lMZcCWW87/QDRz7Uh2hTBJH0w9+Rfa4iX0HrgbfYPC2b0gTjTZyr/nkJrSyZzlh+41jSGaH1XV2
pHiAEg1I2R905e2Ji+PnTmemLU5MaLF6zhcT48pAYfcNfAi2a5rwrV7nIZKw7rJTRmkUuc4eP3Gu
4FaW08PSuRrObDRiDbP+iHnyD0G3o0vgdCGbkJAVXwsKRkxVqqMnir2Xo/U1LCniMiYWkH57CIc2
ZczBLSE37aY4z4nc633M0/WWhW8ktTvnVRzsAXVIO4juOpOHdDNt6Shny95frG0CJjV2lera9qif
+6460sWlLEAJ0NupjcEtrxl6vaooZgnkfI6IagAqwhRew6Tc/NJsLqsbFdzukoK9mwKpd61d2Eml
THP3md7lw2cyRds61yOdHR+xWJRaDFWiPesyNup7S6StFauzdjItMemaCq96/zZ1gfUHSlkQK53w
CWwpOdSvGRQc4BTQ6D1V8IZcOX8S97djtRwHVkF6WGkcoJO9pZFaqPzA1dGnzxdNUBoDme51LhuV
l/6OPeJOST93baU8/yKiOeeyy2U8rWpsL4tPEmfamRQTxW2S6JwOYifn4/UO0x5AKbIrmns0kn4e
9WS8xVVMNPZuCFqPRTsF7KGKc+9T4rZcAdf6C9CYgAHImXhEcUw4dnIrvhEkQJTF8F1HK+TPxxr9
nBzt0xqddAjcR1o7nmBsWNIrCE8Y9lJ2NOkJQ+h60q+BXwCNrs89O5UcbH5XtdYrvP4baaRJ5K/k
T1ZbGrugNfaucNfTXEFSjc8wXWBfZEhQc7kl/xgC+AE25BWMqhEKRZnxM4hFqQHhWuPit/bdk1eT
/LThKgXDmuRyd6yJSks+MXvyGcuPhMHHdxizuCnGIXIdjeY32rfga71NlWo5M0PBdbBgVvylU2pD
5QCD+4NA3nXNxZCpLAS9gIqL2b3vp/upQl/3zz5TdKQczzzHTaNSRTEcgLs4NdajhSIR1RzQq1be
i302YAB3zuh4U+E7gXP6PHJ/dQvHID8eJattgCzlpIBCpFfr3kUzKcpC5U8CE3KpRorugvWjOhY1
JTq3z51b4Q9W4rWEsA4BIdKcOM+2yq8ztTyOgyhZypXTPp9+n+PuX30N9tzCtJhDrTofcks9ScKU
WoxNjF1vaHgSNIBjvIanOlX+fPErSbGuQ7hRcV9em42xcvLs2BM5dNFWNOGV3eh6+DXm3HS7nGYR
Nfd2KursMQ6Zl0z2C1IN8moSpk32hlh0roYUWQSBLerOD/oir3thAEeI7n3cPYrVNW94GErm407F
6tTyGwLtPYg5bXHUAniha3k3K97b463wPzJrKmFqVlPZvkFEjccbCurpcJt1RWjKtKir+QOQaHaY
IVNdXe5i8een3oUgJJFDpGNUgye/EpcTwwpiyYU+VKVbIjxutLT3UA/tBLn2ZNWBlVLiaQGgjoUn
is+RFJSRRl1ybqOnUnq7TdVBtzVsvY1qACuPDKW4CYKeD/9r8xcHFvOKEi/7Okqiaa2KxavfP1NQ
P4vJIM1zPV9edarjGjsw3GhRv0PmfJ2FAJ4OTd4lF2x3iFQ7RZDwfxpDgdio0DRkEgCiiBis3MKx
E5XQUtRRNyygmnkYIiwjIKTXXkOzdUSYT4y63PSfB+vlIbk4qIDkUDhO96OBlUFGhQ44Md/4Cs/X
sBdk8b4xyi0A3mPp1ewEtaOHc2M60hDTh4AUsVZJLuAL9h/gVnl3SBatgrE+G17gfU2+ddT1mKij
/CTB/G6lQVCitjOwZVTM351W/MLTPO9pm/t5QAzu/47CKR/ISOJUEZS6ZeQvplWgMkEe7IVRX7J/
mP+7/kdOTLeUt5cP6pbjVwtNHvhcQBrkrK4yOUOL7/WKHUprjIE9ONOor+x0rcDT86nZhPbjFBUN
3tb9AwzSGh/xs2TZl4kqPoO4X9mVXte26ofD4APGpmyD0R3YowJ4CbWvSubYpjfLsqA+/cfMTO9+
tS0YuNhdAn23dzTkAPMT22qTyjIMQMgcueqWG0sHOeFBjlR4whAwgf6aD+kmTMPV6z3u4WiO+mtG
2F48xxmUGkMmZzdzT8Je0t4f2K0wUAUdWHYi3F4j5devr7pCreob9h8NeQleYk88T6RdRAlakVjl
7/rEtbrqfztg2Bj2mBsqHsm5yS2r/80YaYhfBHnf/Tgv5Iuw0dn7ctOECp1FkzyNYP+f1L8YWub9
pVKGWwiPrVWHfTiC8XUAsTUGShmVx00FwKWcSpn/dauLW47zpEym406w32zFUOzljb94C3pDwWvG
zRar5WszqeD5j2EAmsRywhEuFbolPZqW8djsKTjBzvALMnfQgfKCNMcROeuAJvst6THIckzwYB62
+dCR0UFN24NZHzgS/p9UB0sHddk9JcVv3DLiUbz+IklZ0NqDWCqMuoVlHLpXstPSrW3wpGJhky+8
rqlylEoR8YldKP8nfurnGSpOgKsxGcWkq8BDu9qBqf4cRjG8sS+DMgntO1zTSddcuVSkS+H6Bmzp
kvmJlMcKzJaghVcTP60qFzJTiIdAvO1LXQ3HIaX1tAaKW5eB16X9gDe7RaDSITGeSQyDhzukP0Fm
FQGmE6m5NWk0unlnukqzGfGVmFbgY8SWFoDNPS5f9MtkQXiMI96DdlLjXMY97wnhamq0BdGPDfVO
GjHFLGMY3GE6hPnNz/wWhAdk62Yskq3QcbCbn1U4jyxP1baiGg5y+anMyy64KnTXPOHXTeA8OD9u
zedFI6govdBccXzxNQLHMbrwCSVd5s9RaqhRsBnhl5dF0DBOrDtl+NOp8B2shr4yIBNBsEw3Im1M
p0+nHIU1XA49NvdxZcfI2ZIBS4QUBk9wjnlts9zKarn1zX3aTVzcjk5w476fei8hGgxure1+1Z0A
iuG6Io6LvfADZjB2nfKzVKrwB4dCiucraBSaiM2LHhVoKtukd0MTmpcJVO0gGgBRDLrUGiWTstOw
NgV4zOPQSXimMJRNlt9umzTQXoG0+IMfboYHy/n1/ly7weV4OGs3hqUapmH3P5Ob0uufmUylIhR8
Zm2Ldm4HAd8xBJ7sed2FSEqmNVS+VI74QFCrJmwzH2HoVx9isDeNKOL9+zHoRtEiJF+F8wu2x78b
JG9tpWua5tIvav4UyXIg53GmbIsqK4Job6gEUCvtosQw/l71Mmdt7LmB9Gy2bol02yNOljw8SBfG
b9V7Mh+7O2medaxRsVPrWZmXbqTyCPenf9sh15mthw6dg4cq8H1iLJ+7zQYDFnit12pI42PKYNzI
ayGlmzuAXYZQ1n9W5kXN8XR1VLJjPAPaWCXFZ9MxQvEW9e89RYTe9/D+kPce+1uBeHi7V1E9vxLs
KJB6KZZdg97T0KJKXTVGbzFYLQ3dWFtIposdAI/CN2cv7dlPnuBy5Y3zIgzWselZ/Wy9mZ3qrcCy
Z1XOufR1e5n0jtSrWFK/e8ai/gx3V1AEwGjNUnj0eod/q9ybzhDmi5MVRVll9iu2QcNnd+kjSfJ5
LSaVqnsrnqQnjcvKjyhbv2ISZwI04b5m7C/oDzIuZoX+QmD62RxMKjoy3wwP3OiykMrlsCB9ltBk
Jt8pp9Msl49Qph1V4gZ8bEkGqkVg2HNkkRmknjHA+O7vXS5T/MJ3q2FGY8KiA+n5l7OmpfcRO82s
v7rNEdLFC71UEPu5Ps2oVCGiCzHLiyrCr3Fdletg8lf0tZvPJ7vQppI79o+hJ20xVG5V3AXelmli
q/1Y8IIATeLdhU4KBp/mm0HSiCXZZrkskzhWskryg6F5q7tEEg8IkMNJ7Dg+jBadz4Q35si6Ax2y
h/2kLTnySpi5/Xg1Ttq4yQARCE82I8biRZGWXeQ6djVch7bZq+NABMMtVyYrtDlutpwKFb0uXqpw
FqJt0t1NP02CBBOXmnsGr/ZveH+KfPORr2Gf/lKWXVA2qXTB3SSR6NOSRFFfo/8eVDZ6fHEZfJQC
Y+tjY7J923lCKOqJ6mTqhHscXaDINjBwxDg+Tthzn8B4quagwV6T9W8ThwWMaB6SLroq3fyioJ+F
6X+8Pf8ugHMR5bKawNOpIW6olqMeX9NATBJTsxsE43lFv0/aPFy23KZAhuT06TDc8PELT/RUpGke
v7k6x+7md2gdH6eOaWWMzfYRqj8PRcqmsVyyVwdV2XgNLSMIKNdF4Go2tIDINiP7HBayDITb3eVb
pow23V1t3I4CLzN7NK5enbTG/VsjlZbbkyMj4twDxLC3iYqzR1n2w7Gzg/SEcNNrpofcf8BjC2I/
6XgdUg+KRkERjpiZ+oDV308bEM//UD5hhD5rOp7xV0c78bgwaHs9sC2MFwzDN+A9H2Nq+L9vxS7q
s0bxZVxbS0/ORnmLGplvKb6ItYhHdRvZ45EnweElz9dcy/T2IxHgDEZfLagHj82S8p1AyvEQ51qp
NF9GRTVdDgHjP8V0906LBntSWiNZn95UKxG4q3OZd0kUfHnApFdFc4kJow/zhDquq9Bnux0ZJPef
w7OAP6ctgP5L5jaAg5mjP/eVk5zAr+9rRX6s6Jn28gHE/ljGEyLO+qUGiOW3vql+3OPTKkIjGnMe
tDN4s7jZlPlfpeILYmoy8GveWEqXfMoYiHrjUoo95pv0MQ1UHKAVeR2f0956uSjh9JOKwQB70I8R
vY8Ep07J18pE6fYD29+Bl98XSJAsfmdHhEpKb6NdYkulfPG7JGe+k1IFAxkmwR1OazLYZto0mXyV
C6TDpBqGzffSpWM+qWAqyd33c0OoD6TGadyZkSPyV3wKxHdsWsiMXG/4LkXlb4hbfrAQLn5Q0gVA
UBuyU2Zbl9/L5EJEJ9i8atUTk7LNOwirStBx3Mf47QIWMQRqPX/BrVag+QDOY8WuDbz+AtUypysD
MR+hYCZFxAFdYDz574F1Ambdut+mlY1C0x8BwyXYK8IKvji2Gmt5Yhyy09PVOjzK89fNDgFhumlu
QDve8j2o4eP3MS+oriH0EK7nZcCLeYYH0gYvkRK3FPuW6hJ0Yf9AfA1htV3YHMNjW5fhTQJNrpCg
XnKT9iQTQyuzCw01xNaaC8GqWTtilbRV9fl5/GuxIG1+QdiAbg/sCCblnTpshv+6E23IQ+NpLQ8r
wig8t14loo2xtxqwoOcOosaUN71pAj3g62x/BgFa0lVkfMzLzzznIg+hs9vVZIb72u1SEeI5XRIc
vUfL52gphTaww6ljw6nghgXb/BcB+V0yx8+j1QycsQaGlD4Prl0iwtskh//ciJPVjQgRYQxhmORN
TRM9fMdVXy0HbbdwUtPIBcN4hQxZ4kDY3zZziipN9NocMyZasTmacXTXu56Iefdz58RADRtbsS6C
/pGfREivPJqxu9QFnuYd+cIl7zYN4DBuevOgxWz30IAIkBGgC2vVoH9AVpZz6TMfVs37MiYrDGAM
1owiB4b9PDUwmbQh1z0wEk6WWk+ELE7t0jVeMCPC6w1BEJJqG+VZAPWB7V3s47tcCZsWpSX5eFNW
3ASkJeaHWcvLceQA9dP20lfMRNKiIHm37TRr7m8Inl8ChlOZS63GCWyq2uyaTMb+rYpBBrhy07Kl
78fykOLQrixazTx5EwpL8nlKN3gZ4hWCrlwDtvKeZCz6Rill7GAQk2RteTmaiJHqMxu7+nw6mSsZ
iTQ1kb59zk+vn2J97iamXU16A2eS+KJ0h4OO/KKogqS7qNipbIWvK/coLN38Y9wu66nrZ0uE50ti
EUzv1+X30+Wl36PzaENrR3yWYcWCZTWUAVKgBt+yaFDA2mVQg9zZ2zy7r+2JoI6ri1E6ZkTHMdU+
295NlBLBgHawMUHrIfPZOQCe+D6eIOeXbNmoqHYK7LfdeG1Vgm7K9nvn3FQd9I9SZNgFK8A4LyI+
+pY+Jt51ofSLmaQrnmNWDIuybMrkOzs4bgz/5t+Nu6OjCufNVXh9UdpcJaaO5iQCqcbtGOjLAUNG
Urjc5WLeu58gntjcrCiJEsFbBgRdPr9Cpi1cnxrZC396tiSKyDhj+n2NpwtF9MUM+59jnWa2vRS9
EROJzWsVtc0hf5qS/Uwnz8URKwPCuG4LufcGcYvpxjkcIs88+biy9FflazhK8TVVyJVBjy0ldLFM
b0j1Gkx8Rh0S0f1epK3JQaLUyRta5ls4Du008NmtwOM4/DW/7wwgS54PGQGwclLMnBOdtgbd/cSY
MrGFBsfwnFYDThpmKvxl3XmT7gq9yIf+oeBJ8tBjfIZNcnwinDCggnS8lyjeu8uh7OGeR4Uuvd1X
Ow/bG6EyCsuURikoDBl4uHEkmiJhdmZSmU2HLWITQTzNMwodKXVIBPX/37uW/Ow7nGIj7fD1MF7c
Eg/jakYI8A1Mddmd3ZaFITyhNcud5FH4Y45ltTKDY6eNe3onsob8K2nddotu+U1bpXUplugiyDeA
lOG++Lek9E4gXZyw2/Zl6CVuawskTMEDshKRShwaYYr1auXllG95FEEkoZ6K7Dmz39rno6A1lbd6
Fje/sX9jMlch5Iiy0yP7vEKOexledSDBizmJF6xEsxuS0fBz1yk4GsFUkSbq/+ZOtmdlsaciVLRI
EPTpCXHQNT5iCLfGF1nKeTvmiTzZfxxHpSgsx2Ww7vFuA6t0xY5/7pbmQmNS2oJ98LwcMq0kpQ4L
9ZGQk24gxF7pK7viC2vjjx1hEUGCj6WRToc/iEYl2Grbw7wJVTnjhkpb2//1Kzsfi+cqqrMiKQdT
g5PDIvV70u0hmbtPkh+WAkCPcQzBh1vNj2+4ajci08sx2VYfx/miU8Kl3tEBO7di5fQ5HpMza5t/
s45u2l4DUv4wHUkqL+Wmoc64/UgKENswLEsxGQ424Q9Tbuu+dlp0W2v8qBtlJvZbUJOEqcDPDuKY
1xghR5IKlhmVZKYCgLwWnTDCKhoNOfZALheCvzUeCXRxGEKEzovlDmI3ZaNt3h2LpGvTdMSyfD3i
DVO6jc32kXYsc9zo5EPLwLDOUVeEAsNNXEPlLnUCD7qh91iS0p1ut47VRPz7BmwpiNVSuOPGEzjT
EAG2ZIwLCsSEbVLQfF0aBjO06ohbSHltYyA6XOJCX76mkztM3WH6nvHjdgmOPDvOxqyxtHOhTFy1
MDKn4iCsFZXTcF7oCpPbFyGTGrKaprJM12Af10Tn/V9c2ab7G6cpJ3sLmawAOLhTP/8IktN5TDX0
c1Zf/duKnNLfe1e2OhButhys/iuT/7fw5hBX0uCKPuh7/NnqHS5yWz5LVX/Zl2zARsfgm1omN6md
yQiztZP3povJwk7BS2IYP7qv8cy8PAvlED4ODCbzJx88V+pccvME0EProRDkWjv0jyRcs6I2qU2L
JmcqzQW5RS1EZlZHqHGSXViQ4RUSI93BOLBapCFhBzjjcjRAtgPaIsFb6qv99a9V0H2qXhVXj+90
1Z+4uDj21hx0e9bVAQm3ivW8ISIlMziQzV+JUzKK8HvLRv+NHij/FFZJGCbbTLVKCtpwEEkh28zZ
mBBwKqz0vZ0l3iQN3bChKjMkFzQ1YsySaQNQFMWpYsS/YQhY4EEB0m2BXoBmLdjaxsgu1PUfJl8g
NlkOh69hCnue/YmdfqB1XJM6OHrLaJaxklPnBG/UZfKzrogGLPaKXUCF3NlGRHq/zweT6uVgoV0n
CS4VSkVng1TS5YqmS2xZeugMpfgwdJFjAsTTKIZ6VKTRw89L8kEc3OiX0jNnJx9aD/17CDeNkNcF
RPyrwjIs5U+Eai9DBkQqBrL0d12FQ4XtpiGLqx0cZ8dzFzhDPKuHT9D02eL9QQ9x2ggm2ytwget8
GTsbkVFsrS0Oql1EI1zZzGwwXDkcamsyPS7MXw4k+O4+zD7ccf/f2m5XAdUtnn3R8Dsug3UVrpQK
RjOZUKJbB/nls5c1HqcqIrtbvBxIYvPCSL8uc0D9eG59n7yqwNzEKTPCTa8u609umUikDQLlnmuk
iq0c08SKXqKDnmIiNGbFOO2beP58K9OJVubhxvyEgVVLnUK7w1K3E1CXYHWdrx3FbNMrRk/vg5j6
aPX7fvaQId+5N2H0blpr7tziVK1YHwXR+voiuw/iYR3sk+TdlbSV8AOvgPSj383bgL6ym27Fe1wq
iIrUsgHKA9gzg9uLG1CzGDsCOwhwgLPnWACSCykPYf3oiUBzbcyFKqgmQoLd2yZDrHrt3ypPNJSu
gQDtacd9YmjW3iomjmzq2qGpVhQik0ZZC1DjtzJVx9wQTKyTVz+QU69WbcezBL1Yjbb6s3yGJKba
nHBAAnJXJS0IQjvbQxc5NUYzYCnplpRLzN7SgYRDDQlfldVyNGa4OwkDVRCpEBzwFcwrzAp6QbgE
WaKwgzaSVfY8nYvSKAwwC59xKRZYyZ5sGpHCVoBmr28FnpJ1/qbo4Tsf7yYPmgqfyz3+S0UvOvZr
Lhifj9TdTOL6/VEBVMHRg+resNEfuBqTyl3Kvfz2eSWP+7ulbuyfy2XyT79NOJ77kacshINtM8Ej
t+KaVkVcTrHiLTpPIbKWYHFPqSu2G9dCzL42gN3/QamIIH8JjDUQnf4jlcrrdlm+I6VDFfMUMFwu
r9FZr9NERrPJAQ0fDUc6vGygOSCqsMNxlYvc4lzN70Umq6wqatxJ2Q5K8xAVpzvwroEPJuzgZT5E
i+TUC7OkqxOXPB1QTVibZD0uNIyV6MsvnMuE7V7lFWnh0dIexd6xrAnTx05UiiaoGYdkQ44XUIWa
T/J6/KEha7/X3u5mZ79LKMmI6qRQfN2BvYQ8orT+qK9fXW9+nouoURd+QNksomNzy9tph4qoH3EO
+QZ0+vTd3vaI8HppJVBbw8VQVoRH7CLM2XjWYsld9LVcqCZBR7MGmog83PNf4a7hGY/75JowHUQt
UcUpLVOM0fyRkywI13wIheq8EooPr4MPFRnIrPgGSvKK97kCmQByeujK61Ii8gnvLPl29mycRwx3
Wvrd2JtgWDelNk5ZpdH10pxgrW1M8kmjPj4G02Bebbg2NqnCMB8O4QzUUd7MTj2zonaGXBTCk2At
F8ReXuaFRKlLes0tH/fQPVVv1wnMrq4PnWVWmT2lZDV3dgYr/NEg/0ps8uj9W2u7cSD+UpIf4Tt2
Scsd7Lbyl3W+Z6DuHDwOI5TKdrgGmuttf+4jRATbQ3IcwztzoURhpKKV4xqzWXBqjNsjRFPzUfKQ
fAIWdLyvUX5y+sddr6MK45ipHPJOiRCCwylhOtiFXwQbBRgs8sv5SETtgLZMCCuSmPjQ07cMizFH
qCQd17yGPhIfPZvUTN9apcdQXsPhtsame37zxpAWZfI2keWRxvoPTuarSArpbLGZbRc3z/sGRQ+/
NbF7UC/iBtVrX4os+TUayNlbgRnh9XG/qbFJQhkqv8WxR3Ixg5B6P3dM616IxmDteCtBVLzTS/0w
Upj2IT9SzLCzxxEs+a+qNMXE5J5R+va3DeRBzZAwLBRGPqKSb5NEKG9QZWUwGpITYW2igwR0VY62
ssE+e6nH1TyF432SekLfPmfif9TnbTb+nRRcVxddLnrIAmgBpCZfLCtLodq+tLivjbSI7Cg+gihc
N8cOGVORSVIwqTGlRLfY9oq646l29EN8v8Kl9oLHaNsKtn0HjpP0lSYqqyai1/2RqXYHdAlrciX0
Iik7ZXAqCSq5o0yL1xP2xkrKjYVllCbomAG0hU9qMBVXXvPIIwl2U7HBqhO9FO+p4QCAhEHPYrCV
swq1y6l4JI8uFsLu2ialhnABssGHwDJ7tuRkNIKD/Jiw0lIfwxde9IsfH6MjXz3Fvbxa8XNokYJH
/w2DAw8xPB/HZX/jlnLnFa3Lyq0/734JogQu0YHJrdQd6AMhlorptBLr1f0hq2ysDZrrofm1c7II
bx9dXFTcWLwOUWtlgnkDNPN1jBw0QLB8jz0XNYhNi65bG7ByAs/+Pw1XMTeS4TM1H8+u5VNGTKKE
BGWM2cK+azCmyLv19Lc0tKkcMiqSq181JEmsfdK0C08NRcc3xhAVX56ldXhq84dhj8shfNQeLAks
FjRBQE8VGRVBhWlWD3k2urQ0hYsqk10KoGqkgASbk78T5wym+TB8qguBGXV/k5ep3FXEDxqgSiyU
t5DnJHLDnQ2y69tZ3LOz3H6RaR93DgT5H/0QciyWbtYpspKy75hJl30lbJvoNR2pOyxzN4qNnyQ1
3rt57bHg4CubqlgRMs3fym8iU8YMW1JyWN5Nj4w2hY5LsVlN6Ny49aKN3y8MxBwem5zIMlxycLJR
f2gmVt88Herl5ds4nCrkzZYNl/1hyxa5+6MNEqiGyyPRh6GxubHMZn/xRUhRflYRFhXvgycjTlCy
xiMZJYFjRv0USqpkbQtLxrcWBpe4KEkAr1D3I2pdv/mYHRTH5zw07BvKtE/intN7fgEAJHj4uHc/
8+S2SvA+WdkOt44aBuSrODniysjJo+CaCGSehRF8rse1H8XU5S0BWxFLJvJY/Fg1t+W3fRxZN2sb
p++Yshh3EAH8PrGeyv0Sg88epF2rgAYLKlJ73NgWWck6Ca2dJaoBqL96g2oIQJdD/+54zYwXGgmS
67Vb0QcD7eXFTV38sO/CrF3SLeN+wo8bU34JI4YYoHhnqIdTKS9wupFcPiliIL6LQxH598FdasMH
+eSOMSlAWixf5ZX1ZairBMoVY05BMqaaGzx1WB6MFBDr8bzQdHFoZA7Jheq78oQ7KJfuIIcVZPPw
2iJc6VHuh034e/I5A+Tm4OYhhQ4viFBksnojpLRFuKZL9AjpvKmiYWxpR4h8yXGu9nA4MRZiOloO
9KGGpiY7mGybNMtgvRLUiuuizS79AGb+YJuKjJ2O5a4ctuZkVvlB9SbFKAdtzK/LgfwUdmoNSRgf
SNLzDgMwwi7EMlFRhiqF4+/VrrMdwhggdiW/MPbh8VZ5lJ4KQsj5cXWX1bL3ViMA3lZPCZJaAUEK
tAduwm5bjp8Wbj2bPLpHvBODOhRDCjI2cmAMsuPA8JUXOg8BVyDD5W1VhToh6JQkbLL2qOlJS5W7
jFny4LS02sihBBCCHbS8ATwT/XLvoW7b/31NW1BdEv+MbpCPOq1RRmw1P29tP0neLOd8b7hA1qYT
21l8QUDVwQiYVHqbQXwkTqivzhevX7oL3aBvewCDZSHUj4szYaPItW5B3i5i34NJ+ojGOCEKvzaG
qPbx+yGVsc8FjNwIFeykFSeAuKmXOq9dk1/AMrWGlRowf59hSlQKKBBIPA9XJ93/KP8gJdhxvvM4
KYPsZKuYKlpaROsELYnnpcdSNIq7dbrO4rJ1JDVmUkj6UN/9Y/6qlpvxJ1TH9hl+OletHsyqE/oe
oQuZFVH/G2svzbCyAT/K8ooZNZXMN88NzZHgLwcceEHBMUnFKxdTaGfhPfj6PLYUPaXQp8oui25/
CxvgBTUbDuwQ+epOrE7gm3+HTafaebM+kkYsd3NSknYbxXR+Ra6w4YdAuS1YoyJsi+TQd5xoYyqS
5DrGsNCXjNVCuxE593+R/SBqMIphNjoLklTdAn7ILj367jc99MsWW//c89W43Rk08hl9M46n1gAn
XJT95fnOn2JXnd0bEs95UBCxp8lrADgIyNGqc3bFnaLjywdy4AdkYXy3aZOLMQktQ1FPyU4ganhv
0IWwBSHnFLIKA9wKH8k+6FPn0jHn1AEwKPW95ENnPouiKl6/4ML47eLvSUUCZf86ZTKt9WteFED6
YTF7/XZPjRNqzjrfUghvGLVmsaBTI3fiTie53S3E66j94ZLkap57yJ2DvwDdrKRBBrCmMX/w1NFV
Z4lOLxrWkaudeaUIqs648wH7T+Rnh3r4TaaCCTg8mrcGiKoEhn8krMkpyF0+DDOWqWMrQsH72sHI
UtqoZpI3yDMTbspJNH/3Rtm0IaHoXapxSqAX3rJndcmwVb468yPrCBIFFvUfwO5lGTUtX+AD/2DU
ZKqaGkw2I6Rus3Co9a8hCFsLUpzUXPMAfbGmc2Dk22Au/PHOEecDzwLzNFO28IMO7HWgJLxjkpDJ
0459q14RuA1+xVBrmk1qdO3XdPpbT/r4FimBf7BJwFJcY+cngnPp46r2OKLUQl6nZhE8q6hwjR67
Jm5LaZDx6rYN8exweeXEObNIQP1/3QOJWTHCp6J3CnocXxBfgtFteVG/NuV2ykf+GC3CjvJWMJnn
rprVZWlQ0Cd6FCPoHMQ4Ct2KKawjDsz53+DruE6I1SMLTkQUteiDS72sRhv5ToSAmG9n+3RnSY5Z
U9vnhsEGXbGl2EzY22Tf9oD6NINtxXvnblvSuDZ6uFyh5L0tis6ypd4YnrE8wPpc3d/ZlivXRbNJ
CInM4aOMZWIm9ngiC5ByctDgQQ0slz+DrGC67BsgeUig/GKVzp/lqLEeDpAiZPFcavMk/sxiE5Wu
rV+bnInB2P0HAxwVoVszqXsrZXzPH4HzdatMPZgojAX68D0p+gOB9ABkk8RqgjAYXVSrG09t6Nmn
z+id0uXM9sEmK5VYVnz7YyLWtpdZIvF6AstyGEVHuF0qeAdEShTUNHcMd+vaBAtoongNEM9SN12f
cj6Rs1XHfyFr9Xlhn4J8166F03XZqN7FdFGVvlIzGSwPuAcU/9IKVQMZcxhnUru4H8qMVIZI0r7h
eGW/dPVPg7fWfSA1LtrZRG6xsyJgAWZimkdfGWR6QYxKTtjlwetMR08bUIl0F9WZbvdGTjJTZR/J
fb0vUB6crKFA40a9lPDiHHD7KDgugfeP2Th8qeknIiutlRvBoMnrRgzGjESFo8/R63iwOU5PDUvw
5E4A0+7S2CBan4ZMUG+QX67+sRFDv8UnWHl4AEOO+BuimhWoReVkG2FTegdVZK+j3jz7EWMr88g4
JlCfdR+1mMzCMglCD5lLq6IHlzeJDEKIQekAEUvqCSvyRxPtmW5gtifOyNWONjgklw+L4mxfzpre
8G51D3NiRwX8em3omUzDBqOUYr8LLkBRDEq6swxMtBtYQK7DfTUijJWj6LfccjiVFgkV00y7d0fG
OWn+8sB/QfgEAqxBIue4S+quK2V1tGExCSUfroWOGv9HCd+yum/wt7b8YafltZa+ElCLx+MYF3HS
0QfKsmucQUSGSr0mGXnOF+wS0r4cPEcMkaXPphYF9JpkBmH6bA9Zms/xcMrlS4Ti5ORieJ/jFFs2
VCvzboQhQIDLgpMXHoBSFzSEqC6Nl2HS4do+LLfYdwV31YOEDIGhoU3Lz32vay4Rb/WgwvQ/xRTX
xTSWnkJgbp+FOuoEmd6ZiEbc0+liP0z2o+1pYgwhf628L884XX4l1/Ww+3vbh/7dtFs5sAJAfxBw
aFAQLDuN4LoHRHdwLR6VYvk/gBSIPs3j7t+yEapd1/lXwQS85fFWKIptcaaclDpgqBv9m3/xE/H2
UDCedme86Wz2m/6t8U/wmyfwapYPnOh9jahOotMhAkI97kCLhslzAEeGUcU8JOEFY/f6OtVtmWZm
pUDZpz5lynYQC2ge2t98gjP5R6AABI5/HtEqMUYvf//3Ad4CIpUaWK3WkUzNxw8bmIfiS0xdL437
RgTVSaSHg/DtaRtfzTfYDcmDSVh/OISVmGXHvHZz8jYQPucCXaTDJgOJu8AbFtXmLpK5es4RqLX9
oWaYCpkxfqbbGFfwI6vL4l0cyk/WiSsW1qM0fJap0HR/4866uQhBUqIK/gVYE7Jwh5102FT8AUIv
3reivL1MhzM7UEKBVjN5nKgTvhvafv95siNmFf6oT7mtyE/ccYZqLONAd3Z8hVnTZXcTYP7gzYSC
GfV77VJfMBv8yTHHqy7MEK6IhxTLqhkWye5IVvzqh5UN/4qolMIXKNtTIp0B+Gcf4SluAYMuhcm7
cPXm3fZCG/4DUZVpFtxyw7GNFam7TxNPVPg3OpgXyRU4rW36klhkNQwQOWvkPEYA59tSGuTrQM79
aP7TEGG+QB99xWdRLkhY24D1tj7bWwUQFzj8a6SIXsej8B/97/PV3TYGURyylUMD8TnQvL8RC1Lj
f+2Hd3He9ELV2qkkyJ8yTsdIPT+RyWKOvpNBAnLdw7qRy1NzbG990V8HXsWEpJPzAC5HDcvppbcI
bGpgAJEgJQFuspCE3A5VtcZ/eQTIPnZ+f6qgc3TbVgHKrVHrzQ6wMOr7d6/yz+lxfqD7gCkKMMDG
ALkK0Mfk6Vlk8VgAwRbKkPOyvpGILgqbK15pAEdUncEPZKcKvbJmhax/va4+x6LLJApYMERGDO8B
c34ESDcshNQAOVHyT8WDDvLL4w5353DfWSnO+Svd5XS7c2JBIj4H1tDux+nxsU5x9iQDC07Oo021
Ehue7iZV+b7xbegXFEYbzgT92/yMJ+ukNXJirYkfQKso+cTnU9nNpws//GTjv4g07nPwiAc+jUJs
p26STxFKpu8ZPtThb6UiHJnT0IahalF62qoEh1DXcgyqfkco3s86/nbdTpqugYwhIWA7GEqNr/dP
1cQY9yiQd9BBmWJ4ST1nvDPvWV3p1LYdmvpElMUVFQu0fMbzT29Krvycb6bFCgmiNpqoVDle1FyX
F2ogUlMQwCKA8LXwb4o8/ZDM7VrNg7Avzwt76MiXDNum423iy/eQN5ACZBp+ELS8uwdINuQbWzM+
cWy6b1RLSsgpPj/DooFGZqsrudPG3ndBE5UxleaYo/EOWtzYyxnzK2YrcXHBVUx83rMaPxi809EJ
9yJCDVaWaqP17DXq0UmMQvpVm1Ff1WHlTPUhTy6Vzy5FonCF/nfL/TEi0lRALc5kpY6Yo4dUYYsS
R+GmP7XG/V5WXEIO+dumsv9lAfTUfmNtfzs4cjt+z7NyNmqnXextiYgxjhEDhIXtBUBc70VsM4P8
rNXxLdsIYF3emZc2RdakjfCFEEGugsaS2DWdPzYEY9IoUgRKj87a4oTINut+N8fWoQQLQ7y7hrxZ
U6tXfZPd1OAIae0aJlXfa2Tm3Z8ccAFsIPfOvGo4L1sIPTE9OG9zxwbZdU2K9OQ77BQKWWzib3gE
mfJan8gfbEsz5eEExJth9864lDyKhSwLj//wBJpf7cWe1F+spTmWWPorchHdDgD7LG+HEI0l3D3y
XVhqKwrMdhGUG1CX/k9d/247kUd2xeOzYrVTZYGQJKTz/ZRsvqZ51x055SRDjf3mloEYwwiDaevT
d3N03gh7megK4IyppEpHgudsi71FRzRGRF39ecnf5VT1LLuh5pOZu1tG+yQlN7pySlzmlh+JXKlj
VY7by2vsEU4s/rswiQ116WvM2G+omkMQOUN+AJrZjWB2XkvKk7rwROE/QNj37eLuV1jIZ8SQ9mEu
h7RNqK4js9YIUgKAOr/KALLREfnZb0ArLBG78NnlLQP9rhvNERORLjrLI0VEc0kc3GNcj+TMX0or
snSxliCA4Sljd4CCc7c5AXcM1ikyWjfrQ4bbt5Uq8Nd5FhO+qwNXUkyvgpHclO454kvrlwOJ8OBS
sVK0ycDdTBdBkDhoXzQTGDyoya7GyZDOyhSPH8TqUsucUY6ZFXCK16/6sjwSNRJQWSatvlPE5mJO
5CEqYIRdTJ87PRr0JuPunbxuXVc+FEYMEzHEi8XojewAi12Pib0ZuE8YAWyN2qQgr4+klLLR1l0R
JQ0G/NtzyAUQB/S2/MAHrp1kGg/za9GwjrZxZiGctUfnaCO5BhwD62ajCJ32t/nj0h5H9EuauCf+
z0POE14m58bCWBgTDiooPe4rIC0fsNdTp/yzPFuUPjSgVIeRuqb3j4dgLiNeGCxCylJ/qos+PvI1
WxOSwWnGNgAEsbXdSEtRMTO2oNsZMYy1ZQ8DOngD3Zmuidv6s3+ztQr3RSDq3qD6C5hVARbrpZU8
mynfT6vYWmmouhjqTeJojDxv9yC0WSiqZHi3p9sLlE0AgisQuomd/2zsMLGRhZGS0pR9D3u0wOpd
bfVDeKeRZSA7QTcWGNYj1wXQo5IX+gpPsa+gTvdl7G92TzA4m/Jj2gCuxxEy/FhIYN2ACzb9QDWf
v/2V6kSPmmAmf1c/b2NWK2MBE3EWw9WekrOwvBjRqCVaTsh4SVFbK23mO7MJbBiS7FqwqWC80ht+
ozmG7ceKlXiOQl3UpQbK2S/bhn5UyDN+jBWOVF5jSKVkq2QVur7fPUAGyhXoy4DY4C0Zl+3vRoxz
HYCupk3hhbLgeXBvJvIBowOUaPNIlLvnStX31opLtcWlTIrjJO1QVbTxS8pIXUCiYhMQtEDO/Bvl
aH2EigB3hWV1MwbutRIVEVfms6Rn/stvt+Ylw9GmHbdeeKquKXvLcr9TPBK/TPAIZAnbfUQ+6wAl
+elYYV3sRZl5ZNLCP648XaEBdyXe9pY/yhMkZKUgSpn1DpDpNaB/pZ313L1pqBfI1kYYrVDAWEth
PHH6WGvS3VEDKpayE4y6n2jgCbTkqPF8DwHMA1tmZ7d8KvQIzAcn/hZSF+FqjtH88gxKm8Kr2mUh
oVYJqhfXMYD1b5qXGIt/LYTD0mnXoy7rmO5SKic17TSaXFwiC0IhODmWwV3PC7r+ynXAx5am2mhc
7l7saNlPW0HbQ4jQXFjqdxQC7bhrRPfnIUEc4KmrCv2CdzhnprsLrElfZo69h+A3KpUkAEmBn3EQ
AJAYkAWE544HdlNpld9R+h/ZFNQepQDf/wrcqj9t3UGKfY6kap4iQUDdqF/jvf29PLk2iTngiBbQ
kgmBzLa9C8m+Y1KXsFf7yLPb6L1lWFDeCHqt8HdHm9Oz7+7i94VPEPOW3HYk0SVVR0UXtuCESnQN
OmepRd5qohd0ona5bf++NlHkNm2L2TYn+VgtdQz0S4zgHC0858aXrKKvKBKgCeueII0ygSZ36RfZ
oOfvhDncdt9RlS2AJC+ixDviYDB/d3MKCtxcTA8WPqnAVXHmQt0QRReIpt8V427YsKHJprIoSq40
PHDrGxhiO5lLEQgjHbGJW/10evimrWvF5bACVGcb1e4cArMZUadB4OeTqDalwn4BNdxUtN8rFU7z
IZ//QJYZCtQd2l4RbCiNm8dkyCxQPum6zuMvmb+Agk55SB5qlCPGdlKiaPIRjipGDzp+oGXnhUem
b4qEBimnPviO2W82EYxVObNfH3o7Bq8czi/JsQDDoHJNZMMmvfNRpTt1PRAHWsTq2NBKQLCshtX6
GX9zCJKfKecbdoCflUKuDEobdEwEydKhI42PcJ1vSkoixLCYDhDuhhr+lmL5OUEUDtsWAAToAJte
KNP85GpwIQzdKxzuK+EF+RhPYxuel68PbAR2eOAUI3UuujiCx9dZxiZTsTFTrjWqi1aXLvjy9u3O
GdXPQUmezWHBkigMsm1hWIsPTPT0sUZ4Jm3JzXLebvx0VI78L1GTkVP4F6sZ19DnA+2oHgqp/r6P
t7oSqGP9+MnPRlzE4JM+xcQovqpDmlwITKapoL/qgkNU3FTw9kzP5epsp0o+E+dcLKHWfUhcEfKp
xqx0tq5xOtLA1oR/v4DPcLBA8MCcaD9QobCrea5tFIqwR0vNU9cZyNq1HdNklFrNrNhT5Ah1ndBz
mwLkNTCPcHm4bDBDXiz+eXPWGDpOoG/Ja5sOEOxm75cJYeAsEcP1YULLekIx2Q0CYd/nJEgRVOvW
p1MEfyxdtXKMGcSDb6xUlSdhYGbUDfVVK/vAyxcRzDwkYCB2BFNjZP/IgbjumEGFZHffIUrsQ3Yk
I8XU94n2xbaftIUyAYvtvGo5ZyjoTvxfqx3d3yZ8HwXQWg59lj7nFCShzMJKnXwr1XdArod8YExn
+NuY5UdLo8TI9E9DEk1C/OejFOzob8wI3tl0DvvQJJKTiValtZ91RMmzs0w1QEOZu+fEs3aAC+hB
lH5/Nycd2Db6jy5YitrhXRrCCRcQRy5cuTqTAxZnNXKKPPngIG18GRb6s4XPQEotzeXg7pUVdJLH
hBFokfvbUhw7R78OmWqZiQgSQ7JWd8d1Z7XBOfbQcsB+hNRK+4pC8jQi0q6voBWwJzuckjz4P556
Se1XGGXoCJtsJRuepElih2T1OamOjbAyUUZo4Fkmf8O7wz/nbjWaCttEfafjkQhmZ5G38h45SHNb
0goXnTfM7GNQ5xKE7C4Ab4A5QWl2gLIdMRjUY05fO3RW1xRICYZryJqzQRZxR+ThWd6k8ucSnVT8
XBaP0bxy56NjUudUzJI4Kq2jMjJ05VtGxNNp7JkhaaxbZNv+samlEsCEAILvrnE4GdSlWbRsJ1cP
B5A7aVVvkwJE2f/tlQwkvFYx2cBlsJ5B1cYv6U3KiRoe/rqq0S06pwY/DES7AtPOMhSuNCMnaPmN
7flEh0QFNkv7AzvMfCgLJg842kevlyWG4DO5wJdiKxMgGpykEHxzWAuekzcJXnH440mUvDS4r7jN
2o/GQqI3d8M2iniztukTq9ch//YJZVSGq1OR/Xg8t8WaX++2VA62Drqf5S7sfat1yZA4u0QyY1hn
0Pw4B0+4Yh9k364+S7GqO82kyjCQnsGwMAmTggVV4DVMHs2g3riUmJfrHBOgoO2+Q6dbgd13L/2r
5nknuZfdDCYOHbIv3Xe4q3A00eMlfNqLxPLrHv59fqBMfR9qaNe/NsczR8+MAeoCwNr/yJrEejHR
2Tj2jKo2B1GH8ahqRhiU5qgFHuNXB8nLoHp7uNE054K2J49V7fmjNDUtPjg+TrYHWqXBFhnKzQk/
lwEowtNxE9LEf9Z1YH1borHsU4BvM5QMsI1O4JKjgSWOKtj5oqqZxOSdNub3L8C0yJhCeJkbY1rV
G7yWbJn3pDrNrZ+4L5ZihmDo7lbdLoZSPaBzx/l2AIBmdGrt3Dlqv6yyjXyG4YgFfOEoQADwVERt
TMsgQqwKCJBquWl3QsZphByKvu1jJB2IxKdavuWfoGjaqQ5eNimVN2btB/FkvUDohfD2J2PRuUi4
6+Pc/+22IfgnFspjvkyXPKZ4kTJqGZpBq4tn9KDUYVLaYjo1mre2U3VQAV/BHRs9aTmvG+/lr/dD
rPEVtwHkTMKR6SvesiyNq82Xr0rRJ7iSey+Qp/5ckoNhKeR7b3t0PT2Yw299/mlnodvJORSP8t33
hQH3NPseJndZNPfIWXdw8IUoipLM79IyLIMFc3ng8+ldVI+UqOxdbYjp110nEBtxBnQk3HXhfEtK
bL+iDkF7HbX9f3GvoVJB6h1ir84EAbmmKMw3R065WRauHEL83L0hYC7Ebltewq0/hntquXJqr3xu
XMHVeVz38z+zwg8o/+bF3mzRXJmzeoT4Hsl9/8wNTpDoo9GvF+d3DOPzAZgHxv8gya056tl93VdH
BBkjfhl2vvXDxTpY87UmZ/fs4HxMPDddvXowBBLjDs0qxffu0x7OTXwrM9+1GW0GCbCHVghKmMnC
B5dlWLaY10LlxUaOfXVkqUi56XSstFrYstGvOsv86p0SOebCO14zbP4clgtKlYlijVYrjGUUOMC7
cvzmnuoU7A8g01FGsR9aiZ0l7Odgp/sAe7DP++nc6nL8w9p2LJ4o17eTJvR28dLM7aoGlgQXQPJN
Le0EvNYf1cvB2uUthHc5Mim50xTR2XM37QWFw40hI4Y7aTi8+LrmZzSlQ6KImL6iYDEBbrTkOeUR
VflDG2IVWFWRN3woKsPkGO0wMETVP1H2E5SfEu5NxJNroTfkk1r0wBoQZK8sB75Rae7antVcaWpG
Y7K379YKP1vO+w/GZaYeuh00vjOKXIacPWyK4sFz6QnAi65blv6BGFLCkEhzCC5ZxUK6Eh0ymfkq
YbjziMGhlyOv+dFIgF3p49gFOMZulEX7ObEFMarYmU5WNLuRCT7H5HniT9np65UqxhwuAKCg63Dn
cDw6foQ2JjyNcRUV3k6dpj0+kgsYDlKMik9Xx4umAZK/U+l3aSPBqRjv2LOYZlhUh4t/w18pJT8h
h4cV/KV5XrVTRPQ9rMou2ZGya+fAmHMOcwKYn2X1NVvXXGkrpoxJXc6xTq4Qg2pJAsvM3oypoizV
v/v/bNFW4qUP4lmLGJCvp6IGw8Tl+OIqEFRMz7Yjp+KjWWf3IUthF1zaKmHJM8q297nmxnxIpJMe
wk4UDrHrv5YTMSBAd0yuKpMIrFdSw+SUwDOXrBR0JCx88TVGos8A/STbb0hZVJXWermkGGAMO9XC
0yZ0XRFFC4oPizJ7nJ0QKhHkpokdcyPaC1xYiYqjp04xGO9KNbHO9MdEu53FKVPvjpWYLH4Jhjk+
IVGoKgfC5q5Clmny2wmrUHgnobhx1cAPur2HH6A1pU2B6eDTD0Gwp+CjXzA+IPkJxz1e/MxaGi5p
v4WuHH1WTpufcOG4Jv2c7VBumIbLvA0vUThRei4PLKXlf1pFk1p/OsSD7Eudn7QiH0UkjFA4pWXL
px3lnS17GT0Ke31tw021wsqmlucvDS05re68VFFSY4OoUJPMg5n9k5fPl0vyKqYvJf9JJiWekDmu
R3XHaMZlyqmJ/ZwhPb2Nl9n/wHt0E0+0yqksyvQ59hAaJ04SOL4fjkZInJyzUdEJ1VjGdM7y68SY
bbhqyjplKYVYRdhlCuHgywtDt5AjlS/54fHdm1mQdmh0sB+4afRcZXKJfqpH3CCiZZFT2yXnBfQR
n0gqh7gP4Z99NGX/mefEzcI9Qa6pisK8G0Ibbh1ePWkGtOgA2N50u4qKbIsVIx6NLPwiWvlUCdpD
xQ86QuLHhvpI8kY8YSOVECmJllZoYk2935zC/MXHopFMrMWRHxTDersymlVfzvImyp8FlW4Fu3eK
t0mwJcvX5NEZ9FgT0Qz9fbiXBWNl6OOk+Gi3omjn2/p6Gqi86SnTQ+jEwdvGYWrTFlYu9rQX/keb
Rc+Z0KjV07xlTxbffUtpywVrTr1NatjtMPnVF2k8PWcotB9bkNBX6OyFsSwo4wSJ8RCYQbivT2oZ
YckLToCZD9Ou/K0mdQ1VM+P0EZiHgkSoev8lRYocCV25DGjE2y6OpMRur/U6/dJ7DGOHGW/n1Xz1
LwRr9EvnNJbnE38ZysnLxRse2Di19dnt6Qfkjca5QTbdUsaf0Na3FtyhmJMVfvTZmp5dZJ7LBPjm
NS2XOjXYUNutZzKFMCWlP5nlOEBi9E3ftHjmKFfCmvJR0nQVkb1wGV9rT/YmEW+FGh5WLUqD31XK
9/tFr2llDqawwdVNnDhkPgARUAAYFixEQ7kAl2vp7pHZ0VPhM/dQXs4mTrTgf7Ee0gezJTYDfMWG
se1epich14gczE1yCoFlUlfdUlevcjS690zwgGWsScXY/3d/lV8yJ02wUV74/WJ3hO7KomYlIsPj
02pgDJC4z/xAzwDqbpzNeCA/ahjO01Br2cwn7I2tURkKxfDniFbEODb00aJGiU3vPxO9Fz+yZs3Q
0m7y5izNDYu0Mqn6IB+w2UKBryxpIVhLu2T7SVjY4aJyNaW/lWxpn6AiQbFwkixwqVxc3iQZhtL0
GKYUMLIOgfxHU/QsDvS78kkSEJruwtzOuvhubpb78lvhb+IzMnGMasUt2sQNzlK6FFM4TNyLZaT1
XzpGWv8TVP1vpynu91+Ey4Bzp97FPW8N7b3kuFJyNwiRLQV6vpkEF30uk7PcEh/MhIXsPv4u+M0c
ssGe4NQ7zJMQiDjBRBjOhsNRuSGG5bKd40w6RR/zETDjmkMvfyNz6cHCd8qA+W923jBlEefoJWv7
jl4oYyUpRjUXu2qX2uyG2bQYHJJYSLFXYY/5u5SeUCcx4ZNxbDfPgjC8aJiw1F+TfJuFVExEPN73
BtTFrwZImiVxJ9kGY/q7QpPmwUub5FZPttA7/eNwoAlH3W+ruu7FWYvubQa47+RFaR+CSB8hRIqB
IdZgg2Zdue6BTTCoDNvT76xFbBN16bbzKCwn8WqRPd3qbTUdwPIsx6sX4Wjb0X5g7elQk0HjoWgq
V/x9EcMCukfnVOZr/qbAcIGwsfM7DotkAEpmG3jDgUkyebb1GMlJ9Tuh/DoCaWxwVORYGQ3b1EV2
hr/cTcfXX3+6hXIRtt0CSyAjwzxlJxIer6iu/lvm1I0e7IzEpmOt5Vi8qUETi8U3M25esQEXGJ4p
hguRU/Vcxw7j7+56JsjhyfwgCgKErQDU8jqVeTsk/+CO1D8pZF7nCARG0gQKU6F6Yyd5bx4idf/t
IUrobufwz9MuyH4g5pqA1JSwfsB9k0Qte44DHHWP1yBZmHm2Oa5RKVejZ9Ld7zvyGTpyCEeUIJPq
2z4KJ/XKyoTjUOqJq65dP13OMJnLiLWYmJ/1IbG7U2DMVbwzvGUNzyYtRnbVdZLngleUh5D2nx5X
uP4MRZk38CspolviMxCVy6h9c3M7YvSYE3FLWB6q6zYZk52rhNgkHvNaKLdNolOSR2BHtQlqeiP8
e6POmyA0iRTkklUZsY1nCKArQlfZMbnEWZKNPF88Tkig7jZpOnZxYuEqNsqoiQqNzWxGpLlOx7M5
4AICOzwOcIYvI5697HZT7pZDXH8bLQXdN2aYY+hbUUsLACjqcutHQmP++QsyOORASzfddU79IyEo
wfEUqt3vsfX6Uw8649H3RlMfXNM2j3pd+sw8+/w/bInGa50MeO5oktz2WjFQCe1C6JJKAUnpiSnq
+jSfKlXmbhv0Dfod4kCryE/ST7FSueh4Mt8G3tHZMddfz41LD1tApjpB01e08nYqUZUPu9tLguk2
kDNQ2xne0P3awQmgPOXuKAdYVcHVzA154fQS5KodhmaJA1TfUjtc5q/iOusbCPhlIRsywIvNxFv1
DdQVkgwYtM2gO8D5A1zq5d/DK/fUy2o9qoSHH2rCNUw8Zsyhj81CMGdRdTse+umw4SN4vi8AfBtZ
29xWFkHgaG9t6NmbPEgFo25ODV47mA3BBqPB9taI4JKi2LCQH3EG8MT2432e3B9/EqTjrjY5X2W3
YWLtJH7CvAO6qYxoH7W5c77IZPRcfSTIiJ/iZc/2BNITEqS4KZXhv2A/wo8dFlBF/MDZO9ASgqg2
cMmvMRD2FMSILmfhzTQzQyc6B9DUU6ya7Mu+V7OyJv3PnfGmzrsY4aiMGF0F2Qzup9DNlZkLsPEy
FaPifXmOxkBptY3kgUb57CNnm+mA71hGHm0RM1eOSEMTt6smWqZ22TJIfbtSeyFKqfvg/h0QXJfT
yOqejN13/ycc9f1BPg/O9B/g0sNTN3J2gDBv14lIERiaXfj8187hxo0RSw3VboADPhs/eCiT8Hjt
FLECNEmYYuALz+SAsd1PUN5lO1WFzoVQA2bgCbY9O9F9vI5d3FAlwx3SzMKgCNV46ZafXDQl9JLw
q2uFExIFJgHKyn2HaXVwD+61zVQxjD30TwY/aYEd3lhN6xzzhwke2UVolBauzFiUT0jzDdHoxcjd
VEQ2lxIwZGZo+u+fdNq+WP+HzaVD3C+bTeZ+S2znj0sWF1N/4co6ZpToctFODpQj2NpPTwKuPuw/
Fa5ItcaqLk3dL/pP9KckadPtQAsraBoN4L+1yd9pk9612CmO9AfxOc68DQKH4w77ksZh8N7ApEAs
SrevKlz1bzqimmA1ML0vI6QYzywSrVim07OLxrYUzKTIUXneSS5EwAnMpmiNeBIlOdaLM43N5Ajs
m7NAokqRhXMNn7O0GeXHbLvkP1l2KWJTctjkBknuOfY6nF9aS1EHFQV9JK1hM352RoOvGqGBX3Mu
eeBqRgCQ99Z1So1L17FwfjP7y7US67Vg++36crE8ksn9M458KLcDKn0/NzG9+Q8gDPGbZ1CTd30n
VCyx0AYVqYkRTcjseRP9xA5RQMeO9DWlb3o5Hye6FlC+QYBFe6Em6B2ld+ZhziOZQqdZswVyy5BM
pgw2A0t3QGejGaKt5Xs+fey18jjVNw9HXKLkiwZwjxBtQJavMAW/+BcFrbhd7X03i/hZnZibzB8o
lmqLsxNe37ukSgyJIz89o8Q3c4m1Zp3xGjq9DJy27dYd1g7mfO3UuApMWQ4ZD96Zr90hZuJk3KQp
gM84rgQ72DVDirmJxDIv0IB3swbSyCe7c39Xzd+M/tZR/oSuxWKMAYQJdKo9f4hJRQAP8Pms+Rko
xdMy8T3MN8HUK7Qzy8OPX2DeYTKy30DvhFMrtzbYEYHL2rswBMuI4eXsQ8xBp+jff4UXmq6nYPWL
wAicocgY9w6XN02tXisMesmU7SZqVMVOQ8QZBGI=
`protect end_protected

