

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
EHhlU67zSXzve/de+KpY85nXXvMNuZL7tYgf9fn2xs2MMX6KZ+NkxxVYV7RC95SlNzgUt4DfQ4/9
3ul1mLnDjQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
UlAZFSxNoqgvPPKliBxVt5c0coSpd2sh9B8mE9L64FOLOsIE10QbDZBGLO1c2gEWIwuQ23M7QvQA
5NLCK/AU93Cer6u3Y5Kw85Zu7Q3cTJ6gtsPScNo+F/wtG37D/TBvZy9QIxLBvCRLOZx77GL+Y61M
X3HQ3kaL5tpBN9LRA7Y=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
BhywTGDm5IJZmP+63CSoL/TDCpGJVG3VkCIbV3f5gGTJ6iLDPwvtFhhY8681GBR+EoOyUSMbP3AZ
DMFHBgscpLa8vafzBYp5kDkIAp6zpVke5p8WT0T374mfT86d/rJV4lUvVArJtTXZ7Qb2BRu+oMwW
4NXsxCdhgqbldJw6uUCqk28aEPgcbivrgwKY8foWfBnTw+EKHyn/oWDvwghTokcxfEnmhIMsR0T3
yD/98FKNKviERlHfn1BhQ/aqkW51Vp/q5U9qrKs/+lZwoRMsy8lRZRggDQnNmQrFO+0t1Oq/DlpL
Pzgpskdyam5KjVkaaUDiD9LunE1mnunv1fkvkQ==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
M0G+I4o5qs/wY3cBNkJHuC5SdvD7yJrXn6vr03zDaDrjCzuSM2xSWnhAroxnc+rs8YiB5XG+kxRS
nfrpZghhDmt8SYAMsT5eb/ToWHwFcmxPkOwf0TCRf7UHox/rcVr0f6gppZYuBp8i/HMdTy7/9hVi
Jazk/jJ0qiENaXH3lhU=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
II8O6ksX/NQP2v4t19inJMyzBruYXofFp7EnZduWuRh3lmwU4/uZj2tsoMzEFI9GURJGr6OGMrIR
LHPoTtEBaHFBnPNcL2m+mOF2hh90g7CmgF4J8nr08oNvCPZORB5fd/Cj4ujbrC4saBHdapCX/nOt
W3mratI2AGAl+T3t7Q0k1PLokEpC1hOrn+eLqLqV9hKaNBlW7DfM0Swj9M60AbHp0kL8sQjj6PfO
zKNcq6Xvq1JnJLzZ115Py+hhtw8g3az1/vAI3s/sf20/ggZ0t1s4m7+wPif6Tf6IZJCySXPmKW47
LjAxEb+MGgXZe5eFDZ4nbVPt5Q03mtQWzOAzTQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 6240)
`protect data_block
8eM14QBsfQQ3kgqaNN2TZjCXifxbhrI+y9BZs5DzHavW8ZqlnfKXpatjGaSYFwgp0rxgjAuzWPsG
Tdbn3jiY+gYgLg/bdU02HrWos8vKBuGkNsO/nhidNYUdh0ZkI9EntjsszFRKI6krwacp5eibSInk
6aRYQITh3A4YtnoN6pEQxy/ngzJCnML9/8L+BwxG2FwzF8LcbFbQywlh23nEFt+aRQYVldAkrWxz
0qM+vbk7Ifd1dZcYh6e5L+A4swMyO1X1XGu6hnSFXFUheXnWX/ZJGxqg7UdrGwtYzHGMGPvwPetE
g2UhcdQe8L7iQGfV9r0dpxkAWWoGT2QTalxr/wmGiKnsO6X8xQmJZqRLAD3q74kxogHY8DYdbdyq
xvKbs0+G9gm3coyCarkh+BmAc3h3cfkkWfpZPzUuX+vPsTdVLEslu7eeSHXH1SOMXcw1N0lE88Q6
OLJO1vM/p6zNX9fsEkeZiJPV7aVfGYmhNayVTWp5imPNUfZpvePvSBgk7T18LGFgXQSI4ZuEu25R
zTIbVA2od23xoSprnWRY2hOBg4JCZkFm3ahfeFGCLhAja5olaNH50MifAPMub7BiHVm/5rrlTzLS
5CB3IxX+R7e/F9d0X8AcUUQOoNHVV80ZAjzvuu12DNOv0FMjmAiCmpQbltGzLYwFiJVDrrBrLPUy
YJgnpjR0pIuzJKTSAw04H3AQiRzCB3wYjRH89+b2QUE2lQ57UfSG4WdgBRlOgSU9o1C/2zZ4O4Sf
nV5tYldKSZ7fYJ6YoKTOSuR0vK7IeoQ/pkJcEzL049iTwSTOugJuVmHVzFiPAj3iL004wWaH29jM
1ahwYX26aUY9xxrUnbxyM5z7n3DsGSR45Dfzn/zknculOs9f2ojUgJxueHCxxIMg0NC26Il2EIBY
OeH60d8bRq/PoYOD5E5ubVtK6jJG3GIijbPU5jzF5TtPwQ/maBHHmd3ZySW7YjzF1Q3Ki+IpSgxT
tao9R8N5pgf1pZd/3+3AfoFBiLPi41wAUOh/4YXPpZnMk477/kf5f51Cj3mg4MUxs/XUrmZR8/t0
4O6xvJ4E+y+nAJ4D+oKRLVqalGQp61HSEx3xEObED69t4/aPMHguXAyyvNgIovzLk3jGOMa8yxGK
JoOOsQ2ZaqcpEqJ65YW2mHB4pmyh2JXBtw/93vHH5MdBqlrLa8aywiZ7ZAGrjZqFkRX/N7TAF0cH
qCPTC2FcYLq3dHlumyoQXAt2slm3CrbVruh3t/6l2XZVooaS8dyzOpjErPyAZpktvik+sVLE5PMA
QT7HDvMQ67v3JLD2PljuJ74CEaf8FPwkqBUNWwdEbzgamfB+QM1SaAF3DCAfjymbncZT++3EALuS
M0k37oy7oI3J6BQrrfaCx20rqd8WobTEkcxF+syip4q2QuUca9jQbjkt0ctjZnNsPHIn4vlRlnBw
odbZ2nSOBrsQfYg8leqFqmeAKTFvaeYJyRWOj55zIMpKPun8mXlmQgc9vSfoP6fPdMiFVpecz6a+
o1ZaEz0ofGqIlmESsmAt12uR80FEYL99dYvRxqP+be202ENebhOnHQlqbRu31BnuDxaM/SxXCMkR
OecR/tEmIZ5m9BwrcJcbUSy4SOQRdhxv9KHbao1NyIElVYcmUk1qp9vReYJv2/jpHRn+esQJhxta
IuOJo2Yk9Kxz/J480sCT0iZOtuHnOhXkJcF0c/zm77153axZ831CdFo1C2Q9wtobCVGUzkLev1dA
q+uBdSkBmCFdu8nBtZqvT1zXy9ZD6nF5qIstL7nU7qeT2EgRCyKaNSb051ug6Lujd9iEy9LinE8H
UVZVlG9v0xMkDYdSIt+sXfpX85YfZbl+5bScGc1s3igqNpltEOqiDsYGbDXTEVOgyKmEKoMOnPag
Xbx1pMs2Nz68JnP6OyCyM1n+fOllKzqOipOWf4a407l6G23/0bjk3lLXOsgror2hWkM7OEaVMd0f
2YKTzb6oWBwfJ/Wlw7J7Ql+6Ph7xWaoIXAiKHIWnb9zflEGi/W0faR41p/1j36KZ/yh4YgRraL/x
W+b4ABRj7K6wpkoHDbhY6kykRDJm3pbElvg+1xlUE/Gt4cKl7UPP27kbsO3j1x9SIAaKZD3RSlvQ
WkLJrZceCAw7StzrSlUc2fvrkvW1evBOVdudxFc9BgnEeGSOKT5B+J3g8S+GSIXV7ZW8GYi0WF60
4IXisjM1JScksm9u8xWLNA27NlvVrBjvWxgXHLU+ohHfYh7ZM+r4Wm8LHRyIx5MyUPWlI2K01xBc
ZKyPk5mERojFXJdcybPBDXKa5OeeMOepXZikZDwtA+bwF2JrQTCFqONnKdmNvulAnV0+IctzNHLX
32pHQCxZaF5Lt3NB2F4Kbyt0fLXaChtaudUh7ehJL37LGEQY2EcLB9qufTLKjZ0Ibf4oMJaAyiym
cOzOJYw2SbkZL57WAjtMufZ2vzP1svZ4IT9UMv5QtMutTlTmsGzVEW9z1MO5+k+PNOMJWqwzVjmH
JacSwwj4WBbaelxn70g9K7qIKIbTXDg6IQV528IVw9K+Qfc9BJRroPy5lprgncldc4LXDBjBPJKe
mXj/CdBEUxEYNipsheXPtbHXtDdmxb3Pf4djShLSQKn12hLv0msQneN2t1Af7G2+IxyBlVo3zIjf
tvYggLfmrnN75lkx4vCiMVAj7ATcHd2sutweKr7+TkBaGjWqOnPsbJrTjQKMn9EfGeLlL6iT1Y5J
MQxNEEoK6euLZdK+Ny6yhbBVRKIVQRXNWiM3Dt5c4t0AKyXN8nHcM7HMKk2EZ/lB0gd/G2Rt3MwE
G6MvyA7jh6VQCf07jGch5jpZgMjfjQaxCcMrv74EFVYxooQzQklNjrWo8apVXZx3hweSF1lCRgoR
0DXSWipw7Z3PKZatmIjVrAtd0fibheG44CN0sksr8T2QenA8BUtyfJfykwW5oug5cplKgQtSXCU1
wzwHLqEL2y6nOol3aZqbVCByLkYW9G/fGBEb3DavXjPfpakgiSfqJgKE3k35BI1SGBWOvIA5Eieh
sazWKCv5N6VgE9QkSNBC9+7vEtuVQR9LB10k2Hh2CrGdTKSF2qyICLQxj9nCm/EXh6gYcQhJZeKA
tVwJwZ6aQRHSEiKi4tnUaHO29RGd2paFZouOjryRbgfmnAfUUN24EQaIGR0jVvNhm9ou6iswp3Ho
B6IPgkA4pIsswfxM9QA+4EOj+QQfOAHiQwqy1emJA833Yz+UGOpKEaVa0+3QDbB43dZJc+7c4IhK
FPT0qiolxHJDPE2R/fSeQSM4/b6XUFUyA1uqX6xyj7lxe0WWJzwG8tPqVW1SyTlZiow765W6taeC
1x/9J+HdqawB568iZ+lp2oh4DIUF+bzFn3ntfsSOcARITwRkL1G7W+KvtsWp1PN2GSxineMRxhzZ
1UW/5/RxU+9wDEJqeY/sJkxGaVOQCBjwQ6dSnGo/xsMHWasnVpEa23focB8gvJvabckgcN1HkK8/
vHegIZiawIUBBFhsbVPVfJW01G0yO2YgVqCMpop+dbuyJ+h1Uh34TgmwjWngHstWO7E9yRCowKEa
mufqe0KuwmXHGl982YMXfXAMAJMVzGQS1Hlq6W69pJeUnF1PjBavsbGAq90nsT+mV+EQD/U7pBo2
/+4X/zjTsL2imfzdxL6zlWV7VJggFobyaHMvkO8X5928ll8D9T6ZntH621AJQ1HhfaNXzxny+0QT
GG479xo4RWig4m3/ofljhO2vpR1EX4wIpM5pTPMa4oq+vrdpmklk0SJp1LxlPCr8ardxJnXqPh3B
PhgzR2XRGMyo/ZXmyZSUzchbaCFpPyh6WEFxtSNXTijRQIrXjSesGSEt2U/E7AEssrST102f3k7I
QjKQty3gLfFRvhK2Oo4xhMEQeomrNBQL3f4OB2UkjUnjntWAaCdLRIvsMjpXf7sqBthaOqwkax8+
UdFWl/KjKwJQ/Az6kq1vACG92MjGBD//EMnhp5hmXUB49b+EXYtwg1lYJp8N1uDAkqxXMvZ7Ajmq
zTBQ6s7qBXS1nLYxuBGbZ6r1/EGWSOrlVJxxguyQ1DtCiGN05yL6tPuWSW8EtK0ybbyC+eaOVN0e
A6H/eFk3ayYP41CzQb9l3RnIHwqbxLJeXo0bQg7PT0kfvo3+mSIpJswQFCYySZMJOz6VEdNNh/V6
ApV4kh1XzpQNoMTuRbn6bRWtWXd1+p8oM+jF8Qknu3OEhI6io+LaTMMsrsQ3e5ZMKjszruAqkccm
ps7RHFdzLLNIo/SVuDWzSRKNwSlwUjOvfLGUMYWW/EzpOnssQhL6VtpCPqAjDCEhCnAEZV2CTbO0
71n8he6WLGAnY29dm7iG6r8XVkI7Tvcef+SkjS1WuX0EaQDyrLZ4WX6WIZ0nbo6+WqPfItMth2sW
3sAhOC7cizgVmJ75No5SApqShHnNhS9PgSHVSEQ97rUN3DGeqeakkOv2F3ojLol78fGIGqAbT9Wn
5VudptxcBhF+n7nv9WGIEFO/HKn5JcGveg9ujI0d5/QwJO2TQ6Q0Hqg5XZd7EV5U2jBXM8AGiEDm
pAuJtuM1M1uBZg5Bgp24YzVL312ECLEE/xpcPfx2VHwXc38fuQa1i/4N5591zh2dccjNOp8u/Hkx
jHvWzWxfS96cjcp9zCUY4+DKe1bklAp75dlZoGFvDpDkAGTKD9ge0XdoHX3GUujfQAt9cR2TEjIg
7N638mtTRyOlWAWheZ0OuIQq5/38hDV9mPP36PHbab6IkCApCS7OHid4pVyJWQ0+L78WfPqQ2wot
9bNbAfz1FagjJzIkIAuEVnZL38EYzfUYoWEi9KZLOGtp01a4BO778n1KDMKWfBnNk+ZgzaiK2rGr
kgIAX9CIjrUwaYLBK/4Mn3S/Zddy/MLSozLD8X5HNh6uOapnh5Dk1NZ/WKhks2l+i7fQKbiDR2YM
hoxZ7G8+00uIU3LUTXMNm5J4Og0AwsVztuO3Z82G+p2QVW7Ei6E45Ts800AsP5HMtwNHHxkQ2zPu
pwld7yp2PJ5w6WA3Hba8y1PFNyjARR3/hKorrzy2A9x8aJ+3izbVFlP4SyRtRlSYVKx2SbQDw+Df
jngcU3BHUOSX3xYxC/Xp4Vzz9s973hlHM5gn3jOBlunYlE4jiae44tHsIPuVGkhP5R0UCeP/eMOX
b5GcEE/PzCotMoHT7KM60UTQFl48dlO40V1qmifj9qKNeG9njqtUzDSvdLwpMyUl25atFMenDHJv
kT+n+kqR2nQttljd0gT6A3xpj+sJLn6tds3eHFynZ9ddrwG6lXYyd2+KQSrkS1P/kTCmWipGqF9T
3m785/a+2gkXWkieevVrAJUISM2F0K+/J8gcS3bLrUiS6X35+28ou1QRhpP72fy3fpyjf6BQnYhC
CX29Qo6QICs+JF9rmsO8IbHA6plH7md7w4vUbDj1RzitR15biaYd+f/vnou/BSbhS2hvS7uiREBJ
ey2wHvo85Rf6wd+X3oslJtT6YkWGLiGdKSGWvVleX3293m/ODJ7WsgejFK/L8sUvKd82lHjCSQdp
l+zSN5sKtBTNoVjnyQP63f4ysfXnJYadf7ycOZIxnr2/EsPcKpi0Mh1pGV+gt6m6KTNnP15gqr6z
iY0MiLy3Q/QQFiDrYrgYUcG5jGJ1kRxV1TkIHIcdR8rc3h2vmt6Ovn78nivGSlErBL7RmYTD2Xzz
+2X9e4P1mCRO4+vr8LnwsWdJuzrLiFxWvS2DbwFKdz65wJJyVhFUFK2qQj+DiZ/aYLRh9zp5Bfl2
v67YwEk/d1SgHTs0U8nIRHUSPm1jO8HRjJez43NvB33VAHWbwCgfscXtQX5Y9DM0/V4/rf4h8xBe
KEdUEbFiU5CliXjuiq9oLRGYYULWc8oD7vJNa/MvhlK0tGcaqIulB+RVDQ3idMdmbJJZIpdFv4Hq
w0MiZVGLJDfcvGfpw5IIrcX61cikrELc8dp51JYP0K1Aup2nD6xb71lGub6pLAHONZZ/0cFDrKu9
5dvkDSfKico6zvRD677tLCroTVsfGKKR2c4a8FtCd85/DM3g8bEEKGahxlc9pxeo9g1a60AW9Mem
KbaqLxwrNyJsycQx8mNuS+TpnTcaxJikt013ZXA3ih9bRtVqp3mnN84ZB1Rp38lFnYhO09nFc7L4
i/ce6q4fK6ekHY3FY0Fl2lMMd4QPZgWlHPsUprFaY4INFDpnaUyckR+PLNFXkpzOBVmHeQ3iqDq4
A9AZJIxOXYYOE6uU0IJ8WUjpdBqfYIgj7xqfBwCYgv09AO7igbdJ4IBDMyksBKU4GMVIE2rJ8FS4
gR6QSwGK+0haa8g24nb7UKabxqnbSimV8iRyqnrDaz6pvsGozQg2Weevehc9F436K/NGg6iZtbSS
dtm1Cbotg2UYyaTyAS1MZOZr7pt929tcBo+zNDYOyNz0J3USyHCak44dxA+CrF1jJjco00nJmZhr
O7Sh6+k0JJ7B2dzKMBv2qBuI4LtqpdIhEi/J992zitxg7Po9dHy8kVkQGwU/mhqoQ0/jsu2kNQWp
kGQDuzTq18gNm11sKzGAiP7y12w7WCKrvptxqXQC1j+XIUJzus4h8iuTJ2f2C2lsMTXfmApd24xp
on7euydAmK9O60GDK0y33vt4iUzZJ4stoLLRiv7JMH2U1c6Uzq3O7DWs6ICqLh29G17uyABRKPZB
i/jSnyzONxNdPyF/69Xu/Tr/UYHOV5//ChjZPMxy7hoQ3ic9hHkVOp0/2TM6/KNsYkt722c2Ij+X
Z35BcdkBA6iTpM3gAxYOz3WDtW4ZY3YHfEFpeknv5b2owELdKm637rjFgo1/0JUEZIPuLiNZJW29
5Nb+atRfNArsI+7vPpcc7s/MPq6ZVv9D56HKB/HhlluXbIG1W84zU0HIpwPywRVGeU1iX41Z8Dr9
GmzwMOp3ZBadp8Q2j/ruTtm7nApfo9gLcxjDXR86CcfG1rx+9kwz4GIUYlOPxVPbW+DWA5IzNwjN
oPBdTEyuthfEfQnu1T25igX4VPBibdEWJ2kenehU4Nx7HtnK1MIUdR7ls2C79bsSN76VSANcYRtt
mna9SaohSGqF1qEFGFedbxj6rpuQx0SZBfr8l6EMYillGVDorxir27ETPfAeajsrD7Iut2IDd8My
tCZG6pOxUSIl+lCMEaFcPSj6UjQxv5gB8zBWQjYmxsg08pxBT5DjGX7nfY3RQ24WhYleHXUQeT+i
eu+7A3befSxXSapYSV9c/L8OyjJib8MMVDs2Gw7eH7iJdfbeaErGrMypO5ifPL7tL7JyausueJ4a
VDr61jqFdJyomMREogSpZJd04qGiRjb1ZphFM5z4MT7PzMSajmv9wISbuVnGhCdOUhpgcmF6jm9n
mqN1EGfJLkUvAzPfc/2khRl/ygP+JTnFU+ey8bdERMqkwnNMV5RIjkDwyFprtGusq0Hl1PsMNo0J
Eg+TSDfRM31ZlZBSXANuxJWq+R2WPwAuVnwImDBV8ul52ogJ9q5vn7c5Aki8or4WuwYUE7/5Q9aL
FUNNQlnuzCOfDt7q2V6z9WJlV5/EL+4xz5fJ9NFYwF3hunspVPmKtuhfbmZc94v8nQ1yn8A86JB8
gbOobD7HcHZqHNDwFhscFr6eer7ktqTr/7KfaEErNcj2d05UJ/Et3BWnl/K76IStngPyZlRHvV42
jRpyCnIRVSKzQJiw5wkWrH/rKpV8oa1tAVbSfqjteNueVuwJJB4cz3y4hirVv3r5zAQFMs6ny4FC
ZpFETFfDGxV3PomkzS479iiRVmmQwg4kkfuKf8T9Y1q32oUU+3nFlkR/UBxiUYs67Djnd8N81ozo
ukTkrApNKPJsfvAiYbUwJI6GpQoqNBlTb3/TCgLzHwH3fUD9lgYKJ/4tcf1sEIRJ+86AjAxxh2LG
yAkKOvgZlDuRYi8yyjuJDHyMce4p9G+jy8xdRFy0ojFkPjkaTwNJSc0/cwUXOs/S/RzWVWwazvij
omynVYW4fKRRB3Lzb5MJdIGWMsHQq4toB1F/LYHTAc8vvbpWVSMFe7scR2JA6ANeXmv+Dmhi6Jr/
Z2Jzz8oF6iLM5ot+R4lwpsOMcV2jOGwOGt6JOinap/36AxeZ13NoCUhEJ9HnSc4q3OkfMd0kUne/
CRzEyhU2/s4OEKw/43qZMyRUuwlsC1I+13AvdzsfkD58TR56DzKcMcQmdjpON6y2vub7hFxw0ER4
xju7mXCLudVMd3XemXfjdrIsp6LfvcMW45z8omwsMK2TuoyvDoa5Gw0Pni3QRv+E7bnkd5xcGUgx
uKnPll+Bze+65horgTUwVfS5xwYuWexwH02q
`protect end_protected

