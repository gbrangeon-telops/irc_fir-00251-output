

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
SOOYAbmSVdMSmEhVcX6OANZAlRBhIeIgp+j8aWie5qMiZZfkKWRKGFlDj4dOK2MxGgpLi60kolAl
iwo8CvQQmg==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
XO8hvx7ayNrMYNs+QowHbS9oiS1GjnY7XWvxUBWvS8S0pBwgguPJgxI5Jawjx75IEBra9z6gur8D
+8bJ3wjB5uOzP0Op4TufbsYZTMy5/IRaR1m1haAiZDNWpnRaJY0iGIl1ZfXnFFB/FNm2d6rg/H7b
+K1wV2KmxNsYmhxGeUs=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
qrXPktUjITPZaeyYovMGSvjyrwEeWSEPCoXArB49zu0J+taotc50izauZkw4BvtuT10+TUqV3pWu
H2Y4+wBhbI0avNdhBTQ6WysNgxNkl4xSoIMSUDeWLPrThpvXqf5EM2xFWnYEsoSt1fOlTzsbNp4Z
xTF0/8eRzGcTqQK8goNirFS4li1yNxnvMyocM7UB0Hgwd4r1WhVfwqexmsE2F2aKD0WceDfUKvzW
BkaD/pggzoFKe9ZBj4krjm5QO6MJe6tmyETtklCe5Tp5KFVAoUG5SSUacYfOW5JRRQQN1B29KV6+
B/PXOjnEprmrDoW2/GvnZUOJ8iICUgvcDDx9Gw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
RfdpJMuL5lneUspdc3THLHWNRfMy7ZKvo7MAlgXNSeMyJ16shj6csIbQx7zWlYY0s5cmQ5qBeuky
S0nRybRR8cWMHwN/9rEo4V+uesao4mJ5GbtqRFTH0pGXUIW0hSA/qLXBAZCtANiThLFmTTovXGQx
QWChhP7QcQZsZBRuEUY=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
KfAPtRUOpYg8KaNj0Wxd1r4Bcs5Lt64mregrxrObBeYBNNIje2iGcuv2d5+PQzzomKwP4NoGlbzx
CSYz6XLlhFat5X0Kad65Lvso8ilyZLrxVgz/cQQVMyGtqJsflyi+jbqMWdWQzDlLboEzDolIGqLM
T16l7bjdTv+UHoBJFQNNpgCUB8RCwZwGjuOrDkNOQRBxFbXP4ewZBD1TITGRJ+9yag2oeIszJxFS
OnxOibAvqbpn5K7zetHoNiQFD0HLxODP6ACT7OZWy2QVwDRr6smLhIBBF+7E8S7up2WgvZZ778OW
7Swo175PkHbmEfmpa+y5XkNQNOq7GC6XNCURkg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 11344)
`protect data_block
pCg2khJc2+eFK4StR3v0GPHok0hRKm3UceOKF8wnM8fqktsI1TlQRJXall940vm/T14svvsGDGyr
Nr8/yuR6F8R2TbDPN8lW6x6TlrXtzuew22nDaNMdtDiqzxJXXA31ckB33SP14lycc8OXOjTg+Hbx
O46Nqqb9xGUyNrvIDG6YM2qvqA2BRo5uZCjXr0TY4ouFt/zi3CtrCpokQB42QJAErCgCJi4HO75o
EyEIX/5VGGFmxEaTfeeqqtvfHRA4/SAmdxIkMJo1osq1K6wUvCE2Amg2qLWXBmWFI/V7z/icuuAV
abjA9JNgxLsxHgz/h8wOKXItr8V2jVNy4Xx30cZPLeuOioHjIXziCbb5a8Xf2jaNbXWgzaVsfkJt
qn0MyWJ1cxZwyhVXZuTiDdgpKXJTJCYusu4kFS+ow73Rn42kksyzPNFvdAdYIQjgiAEVePmaRuvH
V1KIEEYaPiOoy/o6u2hzdEt+uhBHomfO870gBqYaXAEXtewKps+EvIMZ5IR8HI8Dhvp0d6X6/Uc+
6UyP6/rlHwCsUXAl4P+NDgbnwhVtBmcGxgLp80J7DVbhMzi67+Z+x92OgtcWKAti6ZQMmC/IhBWT
Y1Slh83YBBJTbak4rB7JwjEXPnTu0AB7nlPpUqdkzWZAs75ZwEWnNPn+bsicr1lXdSBVTAeYM1Yy
YRyDUR4eNvJmvpX/UtjeJ07zchod9GNmpGeAZ/GXZydWhe5VWPum1mR3Iq5bCc4PyZs3SdhdMZw4
EUvCf4waDPycVR+iB+NPGZCSW4DicoIN68RwAaVd+hGX8IM0IyeAkYIAv9WzmGVCUutkmLNZtmuq
qzfBGJ77pfNVhUSpO5WtjlWsIxYczJXrSedl1amqsLB9NMoNrvLmwKYNgow+3qi4VvU+Jb91eAGK
pVg6QSJHLetft64oh7+mNQqih0NtHKMIq/ljrI4rdpzG513QmP7bphV+Hpc8iSI9OA3BHXtBB6Ph
H/FarbNokq7uv+OwbZO7t6v48U7ZhB6QJLAlNvP0dMr4G/LKynSHZAMWFUrMkFoQC0IP3k1xaXy8
4jUCwaLrX8KQO9cFjWAIdCbbotFz+i9FVAdWNn+RdST0098P8+3bpZp0VUinD1+jf8ZxqDIRuuRD
vFd6Jo8o84157oRyAmZM40S6Iue3MpDKIk0zHqfyl7H88b0xJ1g+DLnOxyQ7lwEPHwIps3uWfvhb
eaYluvNDscoWxNO9FzjyOnozncX3QYEHFBIIzVtSnjDRVyPnTuwbdTXoGJWuxP/b1w8rHIuuP+Ge
49wCEiKeXS7zaUcctztQ8iQhdeGpM4nynTc6oWJddaDyFN4LchDlM2pfbv4OKcj66XYNpZb8h9MM
yp9fIGUpm9cvzUf7PFJTyKBT8gNoSHUuQnUSGsQMqLY+zQcjkAUKgVtt/foiObwFxPnfKWHfJ++G
Ny8ZdF9MrUZxIKnwBh6s767gK81mxhBDjP7Qpv6jDqbgiaCg3gkcTtHls7cEAvp0KxBKDtC2mDMV
kor6TZMuJKvK5A+cxrp0J0lNvEPxvoL61sQsFC1OftikWMtkgNYqV8APiXpTTod/YG553AufasvC
QEHqSpeyII1defMOoPKumHr2moEA9bMwbLBR/BDGf2+T5XVyUlW0Z/EESqGvjWerA8i9+ZqM+8pn
DxXCuSCaj2pRZT5s7Z73NJ0zb4bqf5SvNcUorh4IkcFuWDPAdYbmIotEiB8vu9BvIR2xyaAfd9rM
AmPL4oJETmENPg1156s4v16wq7cZaxi2RCJKLdibLqQTOMbqJpnUAz8DoDXcECoqnQp9lpmos5rt
HFryJPtxndp+3bZkiwUBvof424Akui2tWRCtql5qM6l7VHOSRCb1mLFOWywH39mXL3UlD6nMo6uD
aSzwbAmcbfI6Dq73prtuR3IkzPDI1JUNNMp973Y3n1irGbckJj0qlLAvmfKpc6jBp1hPjtGqOG2M
YF5/tM98HUSEJZ0EtCFFdoghEzRfpbLq7Gi59pV0ASscCk6X7C68rtrWrMUrbeZXnXec/ujWSw78
SXC1sGMbMxGdP6Lm7lnZIkoZjHGA9Pcvuq913GpSSI2YBs1pLmVQkYwg599aqEtlsFG56IdCJTNq
7Ar38VOcXsuofR0xHN6SHJq8QS18ZHr9Es+de48ntOJ9EEzN2i/nc2J4z9WfwhtgYb3ppijd8bmR
JXHoF1dniREoLGSd8cof/i63YsjuAVhXgL0OvZ5nhbPqYiU1PVCKNwAYTEi2OydoSV25vQGazGCF
hS4T1M3xJxYcHT2UOO0Stg/abGW0oQu0OFfGsOLAi0cEWZwcwKppIiqFMN54BR6aZBvYmIbiBvlj
ikUdadYnad0+nZcawnkyqqvhLZjx4kXDG+iQB6NqZVb9y0TcnY8DQ9rl9+aSOp5x6KI4oRHzB8ZV
3THjRM9uZ1LLfvg4+qy+FCbQQlTQ/WGp52T9xrwcE0c2OqCpniAWQOU0nzC7AEwgkvZn5mhDSq7d
rCA5cuvhKxODaA3uedNQCWpOe5Ml8yeRstZ6kxvGHlMlXyn4zv4aw1u/5ssbLLeLWKboWwEzbqMQ
EIYVcMshdvHXHJX765OhBx0kpP5oLQNf+aMZx8W2NR/MKcAI3Eemj9+9RFvTECHYSKYrfIRXiBGA
GegtZ52viVe4/6eSsuixbfyPXPIOXpVoBwrIZDdmBCYm7fCSJVflNbrlyoxtJpmGOX/85WVrlV/3
ns53zLV7UKx/r2Gu3qL6wm0fAt0qVcyR8IffhSFnHtqKV+t4zXz7GXBqaeh1Bv/O3KnlTRooBqye
SS+DZQclJF7PbHZXprTUAM6tOyYNOS4p70VPbGnRAilWPuVWVbna9Kr2FT4T0qB5bfTKantxMR/E
l7E+uNrSfdKiiZp88pQh+b5ojScSnKcch05QA9Kpuk7nEyxkl21SUHmoSgV/4HEZ+wxvkZ+zowcE
zMopZEYms+sXz6uRLN2lMSuPVW20MJJ0stWCElL3ncsQsgMPVWQrVZWxqMO9Gm1/qjGJeskoJGJl
GTdetkDjoHwR5xWKTbOnqA195nqF3V/vnKi7CjHoyO45rIMPlU5K80txgOm10FkWHitB0t9ZfVfY
vlMwfcSgKwC7b1U7V3LXFNMqpbenbsRClno/5aZ+VXOMnbjeDzkfR3X1vXSp0mzd05arDW0ul/p2
bhNUIobG1IoOYEweN2oclpSeRU3erSLXOs8SKntuQQumtrL7rNf9MtS38Mdx/+M5Pi/5aMr9rzIG
dp5NQf3kQUQ6XR59xj2mLtc0lJ+gQcAINWyG9jghJGEBPDTQK0yoLUYi4DMvssPJf7ScbYR2r0rl
WB1qUvdr6J5FHxem1kCTdz0wWnYozMNcsauxbEXJ9v+xLtF6U1T5k4JtXRB/JN86vDVWL0alWlHk
eA4S3fmOmpI1sIrTYF2sHTEwXoVAW7cHZX7u4TW7SVwuNRtBEh1pTMLH2x73HxPlJQpBKYRjV6mD
/RJ7qTs8mqAfPFxGeEcxPKMBUvZCZGyYXSvpzCaT8XdBIpHF4XADyVKegTS84Ab452ktl3qz+OXp
R+HQJtI9Iw8bqY3QcfPeGwn5OFltcaKKxys3F4NJheRkcJazu3Ez8E9fhyhUt5srxPEkzICqi58s
Ddae8ULY7pklikFiZO4rKYNmgdFsVPig/ceIE7jKT8i7B5iTaYlvPh81noKtZYFPtZCMUvhViA6s
SuIb/ffRph6/M0+TLf1lkydsNC7rJPD/0MYYxhm+a2rhMX7IxU9dmEImgM5iVH6N8c/iV7hx5nBE
JBTdGyELgdsdSM0n/A6j75HHBzz9uyQhdO4EnuxHhWbzrg3X3h20BdcuyQfeo7dutCJQ7qCSegEZ
DtKQAAekqwWusw7xQA8EFtH00U/F76DeRzTDc4TDii6B89uzcAPQp8C8zEMEyyF6dp06MGWe53y4
gdRL1AtgoCFivmy1/rm7/GmewqRK+/p3He5OS84GIZZuk3+rKs0u2M4QH7e4Nn6O9zL3IwEDbHCP
Z0uavjC3mOzFQqvRxWRyiu0FFC2txeAMyzx6MkfHSsPit2XB2wleAMSPuVUjRmdFnvl2lmV+76c5
kU90M5hxCSbspUSrcsISJolGDICxSdn1ki0DNnJwfvKTmeQ6bvoLj1cr/LuAJOlKlPFu+VRmcTr7
zUW7mczLOgXx4r7sh3UGdIICkZNxINAeu0w/HpRRqtjJnu1YIep21zMTcsLtwfGs4dEORUwHj2Vr
9V0cUBUGj/P4pbZb6HtKhDok34fhmAZ8u1wFcgNqWE3OW9Z4spqltqvQ+bWm59EeARdVrAfQKVIr
tV9pizKcNEpC+0+cDioPZCQXwsgui8uB6uniYL/LhO1RD0DRSNTsNjYFu1Plw6dkyVuyfZQu3F9D
HbaF1MC4lRPNR2nbixpM+2CMSZz/bbY54mXATiOFugVQXVnNtVRSAlJPqm8FQBvkrVA1C12p+d33
eNU5FzFlXWyBYFGsS/M/KRocSHnASWSXiRQVBsSI5wFqlHR2Jo/rMhVDTX9NvD6rOWA2HikEh+LV
EHF3vkICc1bNhq9KMy12dNODsTBXUf2D1k8IONGLC9TBLH4NqYL9Y5I8F8i7vVLYoNOpXET8gGOQ
+LyW3F/v0qwKSiuyIK0HvnKPyDe0HMDUT3k/s8FTJKQU13ZE6r5ipYusiLT8DMpfCQnEgEQbZ73T
hkItIvh5AEBG/pRo1kGlM5COQMSLVJ70sJoa3mUJ+L0vmsgDNFBj+yUeEX609dGdnEOh9Ft1fuyy
SAuuG371gRfEco3Zfu8xIF8zD0s5VRP8hXUPmw5oGOrOn60qvbpOABkJ/tgBEAvH3u/moONSrsRF
snraybhdp45ieWDqe6GP8IyRlSbCsQ7nWeBOiX1TtFN8GjIeqO/Bx7WZCEFLpQWs7SY38r0LFV8d
PpZCJ1ZJm/L1FG6Tlwwaz/F5lRB4qw+Lz/UTyxBX5JWu26JRm7SG8KgyLhTqC+QF0efSqnMkQXe7
dXZR9mTQCo7fwmR/Wqq+Ce19I3Z7EvYoyT2g6ESRydZsW5OevdDOHAmdgpbf9Yn5oEQu79NRGD6H
j8l8qprfT2sbfFSlW/+n/8pEsvnR/n8fhIoiRzr5JwhJWFG2BrbNJ8lODt83FRcVQxM2vU219szQ
aHmbSseuRSOpEIJDUF/+h4pycFE2k2UArL+HCvsC0n198AwsKg+NnsQjwaBvMv99eLD17GI3Bv1E
KK9BUncva3vJ1bvyUCY0A/mOq9FHKD8qRjlgl5oCZdW2MVpdxhzGp6mTcvIG5GFvCzNE06C6p4yZ
1lcMlKOI8mnBHwH/cMkw93aW8bJ6Ivtwskj9GnaaVqGOcROoum7OiMXrBFzo3JylA0OFD+lEeqIk
c7vKxPHkFv/j/hdnd9dKTSPN8v1VGsMZvZyRj9TpdyM9dvMr+Nd+Mc2wbxe2ZwrJr++8Mu6JjIDr
INcPtYcHNbYUQZzw9+xjuDSOB4yqQZpByGctGggg1MywTFgk1gOVQi0XS+s61HK4FzlB1hTn9AzD
tpV3AitwvIiS4EGnEGZqsfeNYYsP8fWz5yIHb0dpnD3TaiPxxrFJSpdI5EJKS4NQ512L9bCOkimP
zjat8l2dC0Li/vm1FAiOIuMuMvZaFQW16en1s/ug5Eqf+YFSVObk0B8qsY9IY0rOIW6+WYoeXNZe
skxd8UYl6vThvHiqtd/OQ4jdovigfV44vW4RKhZYzlSqr0OX5ApQKs2/2ihOCYasYLaXZVp/75H3
x7a4f6mTgjmhjWedhcsSppZbo/P91kv/eBrYejPqzBnWaARPfQysAoEVp/pNSoHMyKxjA9NDxR9R
UmAkibPpf8WCDwF87AjdZAdMjG1cuUIwPHmnK2WvyphzJY43uhdpz8knV1Y1TKmpJOkonJORX3cg
PNJGY46zsTBEJ3nsLFtzwZY6gJAkKIzs/sSqI7j2IxrX4aL+UkXOkdyFgjo8+WfeGx0VnAFBXd0S
zd1hCsh0gy/ZzFZYTDGRvYSJtqdKrrtB5CKem+mi4nmPO0yRllRfSyEjbX6tfz9AMtJSv+jLJi4o
yy8X1oPMqtmR/sI3+rLYMcOMYrxNNHlVdsUxEpIbTE/eTrBa9SCEA1AtvXf39Njwt8QPTY0NMGlK
U1+UPC3LL0/TGzJiF9NF7+uGVEqGPFmWGbiuFy1Ymbr0Qa+qKOJYUzkX/fwbOiZyYJUTvYnnFLB/
H2BjlCoym1n/VCQcxRLN7I9HXhBwn5EzLon5fjwGmn9N4oD39BGJAlnS7RH6M8QJDEy692DY4yrj
k/1Nc1B6f0CILJrTMTEDjJ3uInC2G/eWlGMuKv2iaX30PRsBQgghYdlqNIhGFw4J4H5mGNLd2JgY
z/FtgNVCtfVboxj8LOhgiydzKNeX1zE6SZ95HSI4lOpeUVRScB7cUTQHFdMFmVGrl3LP3WAqZNGP
OnyH7YYDBZxNjWl12gw9w0B7CkJdpimNXEvLYN5CyGblx6DZ+2K/fN/xKLgODJHund9qjaQJO5Wn
n5D35/nQ9tE56B08n6MwxRmsOH3Ior9mNwUhKp7ENwd6wFuvoKPeF1p0ZZUye1QjjM66byL+uz19
PRhTB7anQppKGeNPi9sAAGRks8NrrS5H1hjt2Aw8Qg7qrDX/1VrQYCvCKI+w3P/oLi6FujFYFuFr
qQaPasLrB62gdxmvbD83eMrviIPdnb0NQNiNVOLGEXvEDaqeh+l7BvbrEXrccqyVhTef0jBYWixs
0rcfECuMKtobhaWWfXyfNCM3c1DXqTrw71TOP9RR6YIWHgkBMQPKVQT4w69z4mWgTHsKyyrgfJrF
g8fmPS1j8pBZuALpxnpArmUjhoIvdaf3lrZoVCTVDCq6UQwiipTmSFeYvVbDxMofEfKM9/DB34bQ
oESOoWhKy+McJGP+Ogels4dU9KrFHk56trDFWeE5R1YqcjT/vMfS43GEEfli/NmM1lhnJNZ7Kups
eayA5/PneHdpBnh+iBwO02tcbgOtPpAuSY/jqtilMDU5kWnq6VhT3UCYwb/JqD3wrRVhFUgBjGT6
aDQVQ8th/sF/G3s6wEKDaQ7rMZCMWcMXZJ5SSpmDHex30PktStSCTjoP0Br5d8nlErTYRwUJNE1C
s89GNyN1IBO9M71/SEb943PwwMMYi9AVh3/nHG6J7dQ/OqT8f400+KxJra+OUGeeMOpCEpdu1qwa
2fpZ4IiH+uheLw41Gdo6VcjB/HlfqYKMKGSgLhbbTWllW2h1bCjdxgRHYED8fwZMVnAE4jpWXMfF
VelCITCtBLz5fVH1ra7y7P9KFIYUGHuOH11lNserdcnnRCbny+95YSQZZgt+3qnqpB0rxkbgTTqT
bez4Nv4AuGsKnXr55vbTDVSvhkFHvIp2ZCFUjceMw2feNm++hOEOYbKbwictpk3bGtCuXG66Cu5u
f5P694M7pP64qToMHtkwpwADeVh00993/1MERG0xdwquMA0/bYmg9wbZXUneEOk2CIJF/iV1QGir
ptJvy6eH+bLJSuJGbi69YJIS28zpnFpXW/xYOQglSjqltY5VGw7VffJhdYyxamLR369KgIJD+yNy
C3sGcEZCaa5BUsjnQnq1QWlwAh5kjE+RMJXOThjtl7Zm76N7nKHE/qwUBs2ydmTTh4Tvhee4iHyQ
qPlB7JpM3jEhx+0A33Q98U0Frxha+QmFwTUvPShKY5J//wF+dX1MRkIrTbbNXU5hGfl67p3iUnaM
k9zdAtml76eFwx2ojCjb8/sOlB7gq+cnNBYmGrVljtG2+rQPQR5/lxw5HRfg9GjcAaFn0AqiEYXK
2gS1eF3hG9dh8VEwC5e8u6mYti6siVjdtQwHku7FA8B7DuX9sXGAvG7CqUek6p+Zh09Iu0JBSm+K
TEb9qKGjpSqGgyTeYvRP4YqBz+Ju/q1w976gZTxjDNjHBuG2re0oqNVZ6fDgx9oNgjbKTXc8oBro
aAzsYoT3KlbxqAH0H84yWPFMfjmuqdD/FdJ62T74be0WUAfnL+NdtbNliSpq9z+axlyl2aVKibKa
Ioib+h6SOF9ASkJwuHk+/7HF3YIcRWKlyxKu0dj9DX63FwGdyqNpLaZwxIAeGR/PYwdLzLDxNKYw
SeKKhchsz3FjDQPXzHhNxB2a24cysZo/Gd+LB/ttWORTzRKoPSLoJ/Bx7R2Kd4MEUYjNsYwmMyzj
4jI1an3hDPg8tzGCv5/8jLqY6JG99+S7tz/9xECFZXr4MkLdn+XrYUe5ZqFbdBC9wF4HhaeoKcPn
R4XM+uIlU26JdrhReBW7zH84q7JvUY1nEmNos8A8y+Hb1Vb5+RxkvRpDcNJj+mMzJRARCZE03tfw
/9WBvKmE3Fy7V4MNKhUCSjQKfIl6jwv7/t9jctDmGHJJyqn2KTXgDiL+jxqsGO5OGhUERBCq9X8+
Ak5skXY/DuZNRTFlPp/HJ3UBkV4bz41o29LtnUFHpBUS6ZqgCzS3HIo2urfwBsiMW0+Ro2a62cy1
CPXl7R6466uMNWO0z9T8Iy1r69pTENYrfJ4ZiJNjZ4MwzaIJ8COgJ/4UN9310RibiKS5id0TwKNT
oR2BSdbGFTL6C8nLdrOz7u4vs5MaUxrlfKT6ESpjLnNSV707fIlvUczQS/MhJZ1PHa/6HU21anQz
/Uv1oqXSJ/7CBO5lTCuBWGBhpY3FhEa0zIR+qSwYQTFyWQ2ECBF9ObNSvP56WFA3FPz+qTTbzbzn
RY0yiEL7oDD9syq0mhuP/pVdv+a76CvzlEezW6YD8F4Q5URmDQ7GE0d5nLE3Mdq04dWusq1PEaZ4
SUYz07MaY6wsielrHpRHZ+HO8FLZX+XcUg5V9HivSmFC5r7F0Z9IWuRN7ardbvMrNaoTF5r/V+KR
EotcYLnery4R8IJaj3M7f8qK7BT1Iyr2gFAmUtJpH9jAZ584l88yA8iNt1MUzqskVUVo/XL7fyZO
f8IDcyYPeKJuud9BUOIK7J78sJyOUhJv0mnC8Wa83jmRBY/lOI3QvCsW2UpkMkFj6LG75FfPl8w+
dRb4/wsSap03Bl6r55b2vpI3az9aEP/09c55VPeyzUQRp9eIoUav7rMp35qX8SgLUlExMLhF3nAr
eIUngt/fML+o9vvw7mjjhzbdaqlcyFDBKeifDGwhRPxXmEo3qwexHyNizv6/bHsSEwzxY/U9cVi8
M41ngCliliieoixt6YZ4JCx0NiNowlUZCTTwCmB1/0GKDDA/sUa9fAQ95sWiPlGAMJ2kG9XTibMW
pQwkL7QyVNVx0NZEvX17vOm6wEZCyOuccxXlNH5J8gvd6ttr7JiVnFmTU7TimYsPqZlOZD2wyaJ2
l6MT1hI9Rji4u9asTrinq4Z3Xtk4nCyh9kRzFrFo0q+rW9yoasyJ/ErQEnVs1nWP+1PGIpQePVf+
+/opMkUxl7cx9fo3ILFgzxX0vj72tsLc9JZaI1dp93DMb2L7D0NqWZfEQ7R4NR7ukAFxoztX4d9g
h4gsftVPUDquojohrm8gNzIO6doFSIKvBbcrHGaeodEzJz4GDX86NOW267DNfR9iIKLQfn02iiGV
qvPLrJeRw3xfUnZaY+v1f5mU/pnp6TzmXtIKdXWZa1si6qKt3LRKdhYrljrl7wJIO/Bf9Dh+nSj/
6V+KD2cXHMeOBq4Mw1QFuzlexEuHPNlinKSatmc5nOuAlbBhq80V8GkaHgiNn2JhrRLlEzq5bm1t
G2g5cFj6WSOKoTw7CCksLuagEnhYiYJrXnCU9UJ0kG6tyuTEAZZL3WHTY4mKaVLsfCYOI57KAbpk
XwDTd3Qc4ym9RnmnmwSOq/FnV/M0PCtMVFD2eh7I3em23yEQ19JH2Owd55ZPOD+C2w1tjZeFrtPz
f5Z97b0J3HeOxoxALaVhgjh0xSoRGbIwQmrvn0RRyAGkREAxz0efb7FHM1BXV80C75k1pYk6QYDk
Y7Lo48YtfZJzCB/hdX16gxZk4JoYEGMVfCEDaKjdEHF9efwOsI2HYCBRrpxs3B4liUifujeVDi3L
vr/HRnSHceEK28kr9D+R4+Q2cTAYHGVUJB3N3GAs4Pv56gVMtWd+5ccFREybkw15Sp+1kHCGUWlb
Qe75PRBT7t4S/J6hvZ/95DHN6nM4wejgqw8c9sixQ3G0mdXGt+jP8spkMJBv7mrXpm6PC6QyVF6w
igYodXTNzzIS+CFvcXATUZ9MAWK8I1LMPOMH3VOYmBZlAWUAZHYZ/4lBhWNOMswa/fXQvUWBj6qk
e2v/a3O/iFobY5f2itH/dlKCpXeME/qCQUlVzHT3l+1UOQBjV5tmYw0bu/EB8CcL0pA2jshCDVcc
HQx+DQf1ZNHm8lCMrWtB74pcoh1n+F0RlCakUMiZRfTBnM6md5yjlT0VWqehasd6bkjpDzn4anXC
hrgoTtZNsN7OORZsILuBRxn3uPU89rW3rZF8Lf2dkIZhmyRJZGSeRf/msgsuKpWnCx2oiXnWYv6E
87Bu4+QLPiIWBoEy5P2K/BYcopN8WeAoNS5L4WCAjGUsVeY3PRLTIIEIQIiXL2enhTDElcmjIf5N
64h7BNl4dpXxRCYbi75XLUT3zPp0/RyRzy6U3KSP59urnHmOCPmpixK3107o0gIJ83Mj/AqNuQbC
KrT0dXRklpNQB5mNcSmruz7LuA/DHjPS4DRw7e5xZNR0LE5ti9hqCrBdN+lO5Fe/2SHVrANGUGqR
1s/oVG9bNIvIxGngqPqpLc4soXnCayn5GY3/RNoqtdkVvSg5yPDLdgtIOWPndKNJXOOeeg1323rd
Fw257GIySY778VS14+U+2pWht583PNzOytiNf3IBU6QN5iXmJjLVhIFc8+jXf3lWpXWW7uis/lnM
3qBGb0SY9VJ77BLmN6fL/Xnbwxyuv7d+Au6XclZKjfL6Np4i8RM95Khx01wVbOtsQkW/1Q4mk5I0
PbB08jS+CRU1uBm4Nm3ZADSxnXrZZTNva/sZMmKBrsowMZrKfCDK5axjeDGbDaLJmZbf06Ifzchy
D7oZqJ3vJrVy04WwU6+AL4cmvUnVK3+d8jIgqJQujp6AR2Fd8XDp4PRNSGiUrIX4i5CypaNpWGCc
RiyX5suqmfj2j+zyQlS7i9gcZ70U7Gc+Q47Ki4yQBc/vPjzFLICeAn6bdfhyYJ5uYSTPUEP+eBET
YVt6wjqbDjgay2oOqwjJNg5+kI0bXwHM/cNAHV3lLHWpfnyDBtC/OTurh3wdnjuIu/Ujf133HaU2
j4liDsluQGqV8e/4PqxQOyEY1fuC0KpGtvEmFsyosulUi1ybqr6e8ROlo62Law1N2gIzC1k3La8o
jy2RKAkk2piYNPuMZSs2N5xVSnTkENXYQO3Jdk+doLiLxV52fo46Yovj3j0EQTjhhAmVCH3ydGsY
jxFGqOITChJMtOQSUbOw9kkj59rtYXDzxDffCKXCuEJxFJRabqXeagvbtySyz22o+U7I9JVTcrl1
dJOzBnh+KIr3hUewEqr9HCLM4GTPNyBgy8BNQLTFLK49MLlA7T7gC+Aj0pEMJfTTsgOvL7BRDHzA
/aJMD/7YYgS7acXbJA0oLAKKRRlsXL75S/BLOo3rI8ONxI8LmXTd3H6ufwyKKVe6bJhd2PD6vHCE
HQvNvPrRauTRuv6mLJJfbGKALCle0XSwgaGF07FhlL9IQ3fb3+W2SDxWTti3/jZD7MW7CIi1bE1I
oTWow3BEgFbgDkagNGDIX5ucnA68JacLd1v7FgubRVgS/Zvh2xaljmNYHRU5xPqkdeVMVCx+R32R
1HujHKQ8iUpsyew4RcJx6MyG29S+wqkThRE0M038N+osfQnvy7H41gXdn16l7V6zhDMJpL0c+N2C
EUg81szLKL6R93MZeyuql++1DSFS8J8ftY+IOAlkWVqOGZGD8cJe17KSGJIvq0P9W5lsLsaigjwA
6wH8wu/Y+YVWjFJSDXY6Z2CfuK03mXkYA28mqkYQ/oUs/ts7aX2ZSz4w1+MiWHFjcpdC5+rscwTy
sejOV9lUlZwjZmkK4+kw6YaiclfEKJoebkivBoKccT4OkTXpXXk3rxy8Z9asOcmiPmcno/yxHK4n
pApoHdK7a2+mgWdX+VKSduSlrCS/A0k94OViKs2PyHKLw8JyrHF6/OH/UnPOGhZOvwv5lAOvD9r7
RmeGCh/R4g4aESBNQX+WmbsaPyRjNgfyDLHEElsxkzXoriOJGrn1QjRkHxvjnVYWtoNHzQdUlw5M
0CKBM43vIQk09gH1j9LV4FM84fiCdRD+iOCl5Hya0N4v542zAEr4Skjwl+lZHxp32k3T2xdMU3MH
G0KKgq6qO8NPLhGwTz5Q1jNtggtX/WVS2ooN1DlxJuEblTPDb0t1aimoZcug+DAfcmCrQez07V+A
kPDa3fJhu3fFZ9Yc6jNpS8TOgwPWywgsehxlSsLtlLvNORXfh7mze4ZnSn85GP0yiUQzvWWxdesw
PP5yrP3DZ7oQuRHh4ONsf1WAsFx5P2MBnK6mZt6CqkBVyxA1P5NxmBl13EVXoCbBZOgl5Kc3elTn
3xR/X/oFKzEDwhuqmdgl+dgZ4wUej8P/b+mNsQU5V8zjDiNvSFpjoT/XAvlkPq3PWiR935JutZSn
9w/EO31MJmoFZhJcg9V+Tr6Bv0sJIDuidNGLKDZg2oc/NBRz0DGHH1ArZQxrzt2XR2snF7l1QQin
LssDfchzgx0kMtrDNXz8oH8rp2nqQWmwXrrQaTA/3Dz3tFAaG1o8BEbup0YeKHUUf9E9OesMCHoq
/fRuOIZSE/2QbzhdtShPcd4uJfX/uPewWSNAstxIMMBMZMgjI8IYnPu9lRpUJXY3+/R6if5dP8ol
KU9jKBGVLs4QjopnvPeWMEMrF7jtYbrXboG9kv8YaBP64y2mZIc10o9NCuQilS7gFraQoyR7Ivbp
YTbHn9rLTanRbWBPOyrtk+gbGeinnuIXu6zwrq+6lz/RkG2H++HvABpxR1Dxqff8tK7TOZJO2RKi
L37yX0lkAKBJjm5r9YL5no9gDlLJp9ZZp/FocyYmHLA3OXwXfgBnU5F+EteU5m5Z6rj12+cOJM2b
LlRopA4qhRRTcj7SU4IM4AndTqDUjjhsuniu3wPVEigU0jtx06ScRHcdIyMiHJy44fDC0A60mAcH
/b9P33RSF4Q5Fvva77kGTlZABj14PAFZTQkflpsye89GiP+XQv9/a30P8KcVIAfMhnnH82aSLSEn
X/tRxcsiE43HJTt9mx16EOjWgeLzkxI/g6t2R/6mLWJj1Tbe4/LbTny7f02KR6Mxvt/hIGSkcdg5
PVD2lVwR7q7txEJLuYYnh8catFdcFAXKepv5f9wTwevwpvvLqHFnI0g6U7ka/RUT9TZrnn+lsiEx
M4sq3cRKgitfGQQV5TV9y0gpM8Lh7rE9Yw5S6nEA2K5KkkEG3a1VCnN8da8lBLUZ1ygza0vGWmlJ
bHyE3GVj4yeRJny+jNdIfTDxdJ5tbJo48OJgk2vjXyJC4I+tjK1Ep9iMYHkie+s4Zm/wAkt/Gdlr
UX5l6XvYofr/ki430paNwp+Tsfi6IyVO1UNR2ACAZ33DL0DpkFdd8Yq0NmJp7gPz30mAA1bab6Kq
2EfZpCarB3RXe/qzh3+yy7iugTGrh7p1l4StiJ4UcZfnXiruF/qpZ9l3+WV1Ft6/aLj7ieCssYgX
IE3fkJAGaf9S69uyFwcuMkiSY1U+/f/mDX/aVitptYVFWg4/fwc3zDIEE6EiysSQMeiGV9S4STeJ
om36sVY+xglqy5rmqAXrIKQPhy2mjoEOWb0lAeGK+Gkid3nOQ7AQ/I1kyFE6N2PT3FkjYOp673FH
lzFWOEjmcCMAIMmCeZMLAQSh3ybi9cpg6lLAgpVtmxygy93vgtg4prerQ9ggd1sHC2TanUvKSbaf
tNuWg8y8JhCzpX8fC896AQ9h2UBE3WNqHZKZytCtc0ZITa7pBCKf3yXJzGbE21xTSYHUTPkaPe4i
Le2PyBZSUfmu1ednkx8NF5gDfZNCwENqMZAuKRGw+uNOf83yADgH0JwPrXpG6xHsR4XAQLgXdWs0
1La9YDMHJrykR+VmqAlo63A4uMS6CqlF13NIJY5T8X6oI2wiywbyXs5s5/5O/2fxtNRl/yfKpDk2
WeUzyTlklNdUZGAWVSYqPZDr5WP+L7WEi48cvyPEZfqiTPn3oghAzxLfOILHsLbsZdKC4iinhXft
+2qWUrEALBVdoTIP1RX/Z+uyN/oZTMjGp3GML6xpRpkUyYKGG+ZsQUFBJHLzIyVJzZaw+INinNPz
zv0S3grxh14NctCCJw/bympsmwtBRThSscj6GxARKw+mT3dLLLOsuX0/BnyZ6FfgARtlfu/rpnc0
CgIaZTn3G7DvCco2ZeUCErdu+hbNDKazn+/kqps48kGYmKgrrAgAg6mtEDZp9waE2q6zPmxt+yTn
trRj2zuq4FRgfRAlutxWFJwQA4ObZgp9x0AY2AA4qfmBjz3nlhgj5VPYVApNVpjJQw/FT3vwSSqs
ko+/CN1TMumO4uT1MZRocWPbOyXNSlIX/dSH1hL82+CDpU8mDez7RUs7SPbFYEq9v0B0uyE38NVD
kIgDtCgJJgLJacDFIpsPlbjILBVyVo1554vKlYwyFjZKG984fUaabA6M1UhMm57WUIrPJI6iwsYC
1r1gegd12SwiDTRW4a4Hs++SWE8Z7Uw3kOrBUsUSbSs70rGp3UORbZfFUEyutwWchPAIu0OXd4jR
DIHd2H6Cl+ZdJNy6brZQYW4KmOGqrMo4JnlD0K+CJY/6wjNFN3dYIKtGg8L2Xc17a2IPByTOw7p5
kCHYRoEDNV2F3XYQMLIVHUrkvEMslm036lFW46ovTf2C75eulteVdZHE0llGIzMEhE2hXabi6ZaI
gYdlLd+MkT0XCktFvFlU70VERS9pJoeVuXURVAKMd9raAXU5AYp56vfqN1ErfP+AQEk3qvJ5dl9X
cb9qRhr4Noi2rIS0i8H1WPvWr52fRO/DkJU2w+H13cdfgdLwBxtfB+W67sCfiAo9SQ2GZpivFhk3
J3gH1oKJXJr7cKxxfKUlaYVpOo5D2Jphg339lqrs78Q5Ab/CUproI4hH1dmq3ZxvSYGI52X+i8tq
Lw==
`protect end_protected

