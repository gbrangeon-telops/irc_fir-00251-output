

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
PpoeUczC12+YQ6zcBW/hk7KVg+x7UTioMUTG7QSkaE8DKLm5OzMFnRnSP2RdM8C+WL55mLvLDYfA
5lOC4Ruqpw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
K3yZ7/h8XZC4VnxKqSX+X1dWQEKELq4EziAIjvSKKzex+MM5ch0NyAGabLWybM0VZcnyA2IuBQRw
LXtEZmU52Vw900CqGAC8j1ob1JJokunlfDgROKOp9VekmhrNu0zlywHl+eh6CQ/t5W76EWfCnLXS
TKcvUxKzMPqBkiVg3Y8=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
NSAGB2MTAPfuv2AfQtQrWIP89UNTneL4Bk6/B2TdOO+6mmG5j3iveazvIvg7qIHwAqHfCGACbbAp
fGS79Be+x6ilLMPgwgbPlwYl5oARsjb29GILZJJbq65kaBdWWJCFrRmIDIFHXq65c5qChGV/7EF5
BRY2p2sjUe67cd7MFOLVO0mKHurU5wiieT+wdpbGs9uEgt/pGFeQKlj4ch2XzN03R8Lg3KmqOC6w
j6pa6lYe8j+sQMdh+WMN3EmYurAN2aA01NOtdnD7EoaLrP3ByXrwCKFB06hQfAMKudCun+42nXbW
17uiY727vjm9PIB2xOmQazUdPEZbwz2Eeua7KQ==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
NPiHNhu2YI6wz7attBCDx15tEqFL81ie9/7cRUJzlr+aO842fU7+GGF/JOlqWsuQg2RB92onmIR9
gKmj6xIVPN77wRnezyej9aQsYy3bBfOSvbf7a7d2lZQT1pTZcYMfp3xveVQ5gTGk/1BN6rnnT8J4
QRALHC2oqPHhQZ427wg=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
aHttOHUQP+m+tZmSEhqIMk3Jbc86fWQ1/2LKPbbHBoOHb+XyETCjDqnDo9IWfpo+m+LC80obW4Zd
cXgM5NoQ9F1AYdG2ggcdGNXeaparpheOz+XWEe8nirOAN+Ks5VYo+yRWYwO3R0Y+0V6Yw8r7cd48
CXttfKVhu2QOlKTiKegYDKMRGhVyrdNkx/KDldRFk70rkBceBbiSjdBniOrozyhG2imBoMkKkCmI
8TwlLhPf5Ra+r8wceN6j4BjOnyQ3EtzJgw91ujnHo20MZFiaPiqLQIavDgBT1y7leXT7TIK9Z2uu
L3Oj5XHzPc1v3FMsMkjnu8xWqC9pP05Ha8xR1w==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 26736)
`protect data_block
Sqd558TAR64FHLhD2daBB+Fy9QVZqK4msqn2AqA1bkg8W9l87ColDQCdV4l6DOIgg2zrF3jYfZZQ
rEU8VjTcdAVl58y0jb3IV9oK0fmkoB2sTuteohcCMl4FUe1xA5My6G3oFjwd8LdT9redEs+ghp9d
y4LT4Xxk0pxoP1xZAi533QCSxie5cfiDe9Cqjihb7GVihiI8AVzq971QvGfdbufPjbKYCGxMLvFr
Bmln8SIR/kbQWsvD2M3DHKzeUJyj3I8I0nYNT3/8YOGvfRDb6hi2yZP4gcf3cjdU6GsNGyfvdQfe
Pdy+n/Pmdm3hqmz8PdHx9UT7OQZ8quR6R5Nzi8HM5fgvqoiRk38TyXLD1s+SoDGP/gLbqvqqauBW
043wL4mQcSa7hZwFTiOMc9wZNok/9q8kZIe86s+V4mMSz+uNfZEAftOwzAsrpPZJ44S7CsN/SEGl
QoqQytjuYdd3TPBFCdVfWdOV+r7bC+M9WlILm40jBIH1pwko7SagasBM9MUN5eCUi2p75MchNol/
ObYSE+LEKDPQlFeEpO1zDum3ACv1Yzbuyk7uXmuhn1MiQnYkfUcD0xBZsO8029WZS7lbRfpz6Dfx
VtuB5F5hvCK/OyrrNyQ8xGOkw57oVWkGG7BP9CAvshxWAo8PtLUI5R+O95B2/FWS+KlK0g/QhdZ5
F73SaLUYHjISmR/jUbWRKYmHBdrq7quNK7oWkIWNwUWYVX/iwYhKWyONybWE+VvQkRq/utib4XJk
/y0k83/4xTqxmVfIjsAKVY0YKZ9Q24/M1N3bDtAGbdwsoLFKLE3hvVFNMqjggDGe6Jd+LRZ8q182
NtbaQvpzFM1Wf21ekaMb28MP2LimBauXygWxZU8lMqCdJuIHSDtTbInugYQyKEjzSYzLpcj2eXPp
BDAMcchL1jRE3fdqZgezegcRW+oseCaM2dJMmIRjBggnQecixnSUKPIUCTALGNlzm2Awg239nDQU
q6g/cy7RMySe5M4OBzLgQtu79nvts+WpeGba6T/6RZMDl5FUVBbcJlHBzSy/C3OpXb3R6jZHcn3v
3EuO8oWK3nhams21/EFVhbwP2MQ9UXgw6vOOI8k3/cqZaAz5tC5m1iZ7rYTJpO6uaHKC61EdMVlY
sMfvBc83cq/oDQt8ytR6pGzxQFnFK10de9K6+hWK3eQ5/amGTma9xnNV6HTAyZDPdGP5YlPQ2Yb4
iUNwTyw0VtbClli3voUvV0tpTszk0Qnn3UZi5nE6Y6YGNJ0wUiGc9IvwVbA2fHrvmV0H5u2OPP/q
pusqEp6d0XiwOTjFiNMogo0VFpa29E1+qmqmfOV49wv+0uFCgggU3tkT05+vGkNzAIm+rGQdRnRO
lENz5f3eIaO39/blHm4B93IeW5kPjIp08WsmKHuTjtploHgrQSSGcB6mA4Mcu7KLFu5Drf1szwtr
SdxP4dwRCqoCKc0K/pX8+jTiOdm00riFwY7QxYRqRBLqYW6hbmb8I9/vXE1y2z3jpKsDq6IMqy6/
KSuX3MRwk6+4bOtQMlYBf+cILpGif80rLApR08o6Aw8K8cQj0HkfnLIXwYzsgZqQOlxx8Zr/ITOn
KVLHy/3PJG3/IQ1y0odKkig9JFe4jwfpG92dVEOJbrVwQiZRYmaVGM4SMKLze3j4mxOV2l5TR9ts
MiKwT+uKUrLsJp7DD9MFr0djUVQjaQzhvj2YwUgtWJ22ZayTSf3Irp3Zv/nJ8PsGAYFCoRkVsjfF
RrVt2UrQH1+EtWn5/PibWcHix6aGug0jzCSBdW5FnrguS3h6COUV3TaNJoGUAqWG0rZupckewM73
9DzQrZbyMH2+kJ+GCQ/Rvj5rsNb0bgWk6CbnTctHJ1fRYgNfoR53zEeqh4oRmV/htb+BiLEQsTm9
vnlKnvtxKWL/gQUwB3aUAWo7ie1tsR+aNDbYoWy61KtA/3Tv2ynVCplI43eWkFNv0UqFewLTnMEe
XIg23XiOLS07E1vvhGaCFA/93K35L5BJeZQsQfM+43evbsbsWhxbq2oiYK6NOJFucvriDaIv/J+j
DIiyCsa4tGnJ9mrvTTFPEuahxL3cD6iD0FjaaczeWWnEbHhJBccujqWD7wyI8w2XUoDe0C6ctA7n
ZCrIw9uVak60BeWpjFpobeEHMA3vy87+25wGmxLusgurziSJ39yMlLX8g8ElGd2ZvRPHScsnQu1e
VZY9DTX2XLDJSz/pcKcU63aTHGXR6PXDDLIOXHM9z2FiuYvhwrQiYaLGC9AnzXjwF4R/KIzwki7a
BwI4bZnkuqhX2GgnRWEc27Fa/GQxN7jOcBSJaUG9DKG18qJOkPpDt4NbJL2f/qNltqTFpzFm2Wb9
alL9WB5gkga+vwSbPvk9+a6mZEw4z+YfCAGNgjtOb5Hp5fSmTeullulUGcyFjGgT/elnR/uZcBWq
0L+LtMj2uSgR8RD1JQB0K2VcleZUxyRoFkkkHHaoCr5SWfEohaeMHBE4/vf/sv9Ox8N3eiEn/oor
W3Ov/MSwq7lurIAqNwE9CLULR6ZaY8K08Aq+MJTxbySmq05uEzb9n5D/n7m/3gtd+2VRphN8I8Hy
2eS78zaGzaLZtF3eRapSq6Ft48HVjf1/UPF4Ht2Wnmnh4Gs0A/xNlowsGKdwjU/shhAqEUHUBEm+
WL/bK0oJRmhi8052F8ixQ9G5jKhibeiJG2Vskyq5x9j37lAZaCxMrKaQfMJuBX1eqceiLbVgcmiZ
ngf52hGnzdaam4nQ07ObPd0q3ii7TSdDle5Ilrp5/y7n9R2wXZazF9YdvFZfGecRuiejQXEE24+N
5xWtNgICAF7zAb/mn3JQpKvSmIFSPgj1TFqUgEzcMR0ru0BYkJmUApHPkev54BiCvNx65piaJMLt
+KGL9s38nBA/7/f0cbsb+/Deqtz9PR0p7m9lBgZqij6KofPD4BuqHYKwjHKl6Wodk1t2R+9lZo7z
b3/WRjXkSCxUbRuc6JVGmaBjq25VxohRcUz2nZg9XEFyVPpp1ZBNEpJ5eS7S15eVjMGo2aGJh1Rr
T5BPLMQYZyjpWjrHnbkuFhzT4zORSn+ErVia2Yos0vOuYSP0j7HFtPmQz+GvnB1s4TCvckcB6+tN
e6oejXQm2OPaOXMbzrtlOFGKJtmL192lR3wVkIhMgISwnCfxIBwe0cZNLNDNbJ6ZB+i18lNNUOl9
FxMnv0iLrotGfvUiEDIiQtehgTgK8sqlkoXFrXsvusq7T2HGtEIlqOujpkW4LARUgUKy37yXobbn
dUycS6o27HDR4yJ3CMl9qgl0sYHu4RWVmaiTyqEWuKqcdZjqgTeuensltEilC6qK/fTKuxPD6Lo9
NYHFXg056C4vZvQik/momci1VRVyh+CN7OqvpwfwE3UhVHgyXJtBYvLc4ZafFI+TXZ7KfNSAb6US
GRh8+NJmkSTkrRcsnbd+wNNUpACMLcgXpSP/hL3LmJnKHpDEtCI03GYaMaqwIYH+Qz06yMekUmE4
n8IkfwqI59CpojRSnsiHASf6SrtMgTHQpSD5r40/3+f6sGhhh1pgN0XTot7W49ONxvXOH2Yw409k
e5KjGJZMIp8lXiTZlkxx2YNPuR9hiSC4ns8N1iWvnm8v/ID2h244K9FWDwJDYVbnmAaAq13T+9wa
9KsLmZ9MkcX/4qo1rShrFCNHCoa3NyzVp/N/K65+EtZHoExMbKhIF+IiQfbzX9bZV3IM5PIsqHKD
aiAJ6GcPEMrnJ5THitLu2itYBtDZHw97nBqWR99KnZnM9bbiXIDw+0x2purgWTEeKwqrTpi4VzFc
DkZhHg5afSVBM9Slg1t/YPh8+pKpy0OKyNmZzRjpLOXWXXPfW1iD2p4iB5w4WrCP9rFLrTjzyIt5
xpYm3ZoBI6VM5adqE0hdJHl2EY11gh1Was2CdvcBDLdUsjT0dY1yhB3/VG7kqsfkMb1M2/rpYvnL
UXZhQxScpNXfozaUoOwpCU9UMVfI/czdnnZlRl0OOJT+BhuYxJ2VW3UAa9Ifsm1sMFbYZ8bx9MAZ
jRwX1g88oruzaODXSstcc8gUn/ZCDP4Nkd4fv2TuzFpZ0ZEjUfLL6tVWCtDf8vm4pSDWh4SS5IVR
6pmCcYjR8C5TtpkKWSYH+AEska2Jx6t6b/uPCn/cZYSUvNEHaxSTqjdGX24xKeiBexz90TzFDp2X
+MScFqlK0M6hPgcFKImous6jt7qp4RR7GdBap/aB78pBCxOwuLeEQVYp97Wos7Yt252BJIu/IEe3
PsNMW9IPSX07c8HMkchhCxwTKhlj3iD3RsvqxKGBHy+NMsaWuu3QVK5ci/XOz7wj14fJHvMcxI7x
o6WJbBHDT5RnrE2yhqDlg9VkLnm3EOTsshqH1w7p6o3abDVwUQBcuTdj4oIXUzJTg656Vbuo8k4Q
xdz3LJo/dLjlZU00CxctRj0ZKPFhW+QabPHqGwYz6O639MfH9+KwAF7EeEteHEoKpnmHrt26YKcX
0Sov42eLe8DytujhaW3lfpgm/NKzMeYik9uyhZzrpPqVwV+AVBEXnoMKgERVtsrRDoW3KGvXft5m
qaY8bKsrllkoUoANSBwR7+WG39n4cD2tNbFRrhyWabAaK6ilfaUlrtKa1CN5SW6oWuj0gBPGPVp9
T3cW0vratoysYERVxTxV4pnzGA9/hzRKsmTWJl2X1kX0HKpRT1cc97Ikr87uoD4He0/UMvA7rsPi
6LAsdqSBVYcfeTrl7v/yZDarHPLTvFYbcdFVhOT/Xvz4vw//v7ccGTl+tHF1i6j4eZoxgOLz8vW7
LAdupku5P9+S1R/JmSNbwE7+BiuAR9nqHVN530dsfP5BRDIbkSnZm13snAbsSYhhwTIyQQ7h59RE
cQnJ8XeEV2NXaT0zDw5Jq0zZW0DwvbdVUiLi3FXGqfeuymnzhTIIaE8GLN/zUsWC2j7pkWXHd7w9
Cy0NNCGZ//zyNOjv/K7AlxJVfCkDX/U+rRelDYr1cOgNR1x6B9BxaEJ1YVZB/qyUMhPDq7IR5Y2U
O4nMP5hiJb/EWSAoaMwzX7JxsE0qxYXqsux/Pu6URaectXd6LFTqJlUrT9Extznlwhl9RlasmloM
Uac6qai/pULnfVAYwrVZvsmwbb7gvJIBU3JsVcfk9dXmOKlfxdDrFbCnDYL5mui1pyYNkmmpsTyp
3AyEBxX1FVBoWUJt5AZERuGBcIPjywkCdRZr1gH5cmiWg9Pd5eQHFaD3Pyt/TodAvb01/UPeK2UX
8/eI9gQWoV2UGdEb5q/lcW3fhcF1Tf+uPDKXwAeH/KGToJmENZdeXyLNitiWZYNsVl5ZC35XxxXr
fZE3eEA//3EdXNhEUeLOH71QNX+QFD2hLU0zcTQeLqbmZrPm9fqkgklIQnIpmbUAKfGuNG0ocU6L
55Wji82e53KAowLCS4DPf98xXPxxbvf+PFWjM0ATR4GGKIwn9w8qi7g/L0+gRRdQDvpaDfhfv1G0
y6/VNQQYkEq8IJ06aQDnKdUcTyvUubNclyBIeOgr+jaag/+o5O7t3bD+tlVfZ/pV/HbgfIV72hIT
pHiAJAmsyZawrtCOmQeDBRe3y/7XKk60jVXTtcpmhkjtW8VuRpIp3rK2AvYURhpdbw/y6/lBnbbt
zrLRhYzC2KIb/W9SDM/YAtTsEbykl0p/DTeHHziu43tH6I7NghWrdAAboeNtFJivUIfY86OOZiwU
31CnxkoHpJMIZQlzhuP4JTN8hH7SQiENHnGKspV+g1M3vBfZTKN6H4Sd2nINfneBDCwKIg7VBksX
JUC2Wcv+cYs6DngRoQHEQP7wVfWLfH2QyAkrEQLzJd1M+eX+kzFYB78fcWo4HQGihsr7cAvcZOBG
tPvNBdnOuTzaLhQPXxbFaSk9C9IGTAak+2MaHTuO0NsjR/F2SxFZyeems9ZXyzFjJJIfJbEqKAUv
BktOayYupxQf3TT9JI1wZEzJ14llGvi1ekzi4RhhuT7DDYYKPZmx+FtLjA8aadEBF97ZBRgmcIjM
k0dB1MFvy4ElvhAIeSzSUioWWfKomx/43GQAFvzjFrIhbCMJldtLN9R4Yw/CdfSlbMxBkfgQ77PC
NiWQs2aXnTVGbyax61ZxfvQ2O7Q244AQ1gSCk5eo3/vQKhJfMmEF4QWiq0IS2fxYZxTgRSbEXtjF
m3Ov/EdYEKposBviq/bNuwO02DN+7852kH+Hp95KYk/TW+ryWQeES27IOSdX8WFS690s6W+8gTmm
bG7EOKuRhMCqqNZX02oAosbE8mvmWEj284wUyA85cIoi0j+ImtiRPbMs+6BFjdLTK0bWpv29Vfwi
abnBqPk6Kywt2vayQUaheG2EeVzeJpbRZF5YR9AF9Sc9WUEdyYx69i8CFyTJ6PBR8g3bc/W2tDzc
2Rui3EuP1YjH2jjwzDtoI0U2lEvAPfjbuh1PsEX55u4bRvQJ30cvghO2UvLE94+XdaQr2wDZwpXq
jxSfbNeFexGS+lBV5LFl9tGvtvLAFpPMxWOQRN7fh45ll4Rec1fSgoC0inNjvbrf0yNrFyre4djX
XiN72i8g1JebMYLsuAroHgtkDtL9evEpYr3DqkZrWRtPleMMU8Rsqla/WRyp/ZEenYopepmIpgFD
gBumZweCAsXxJFo8ZyX5Bm6jUitSyrdtpn6S056vXFl3/gKavEMjQFQNdMOOHw3X0SfhcD5lu23R
ISRviV0WkLdPooaiRde9w3R1hBu9Zpk01yk8qdT5LXzrsCN16KhzBhPNVMEsUi2knDjKbTWc8r6/
ggYfPZcLCWONE3bxWudwBwfXE6SP9WQzgdOJwQVeQJZY2Dp6tGh1fHGEMKboPSOD88fM6WHfuKQO
BKsT5muP37wdmVGFDBaWZzxIUsShMJttTF7nzvn2lxA8QpjIemXm14TvCY01lBanBrRZ3IbcTXyA
pCQK310aLPPiK1QMeaYTOUqHurXTVRW8AJRyZYl5Ys/Rug+s3pKXyr1JFj1uIDtwWhNrBgxFaMSQ
3IunabZjScDZvDqIMMpW+sWu+5+ALr/Roxk2Wxt9Dr4UrDQKOQgt6ugbKAcLlRiso3nc9UNqigNO
G8Pj+4qV5CrO/+DaQi4MLOWrlR+UZEKb+N4EST2FJ8saJLe1gAJM/wvnTcnfh82P3Eueu57rZ7G0
5SQfjMC25uwK2K1pNCOzcwSj6kO7vIIi0EMVnUdMWVtDpaumJGTF5OShykKob3PTLNHzJ0GSKo5x
JpcEBOoHvTI0RiNivC4ZNmelP8MH6XTucvfc5Qh5wBzBheHccz1iyYj69WfdDmoToHcOnUWTBPFd
/HfBtOp8rIdtICeRAIebbhSkpho2QfSJ3QLa4ofUOQ0627iZeMnhEvjP7SrEDBpCZF5h4pt7Szhf
XDecrTMczE20SIuxKobD1TngYP1SA2spBlPD12F3rXfGFQw9UBET07WMvUyzREnUbDbzV+WgdHji
04rjCGrrDLnBBrt9w7uWhlYqURqDNZSTMQLTxLZNnlN6cCfwgMy7JWSgQ21mDKmUQ7+6H6cSR54M
ZKSwwH5nqFaQoHHF3xDSWgDbLESq6dkdVm+RCfpYUfTrKfll1NlE9DtQDuvGoZJrCRc8a3SUuXgX
3R4mGwbDcSvz6+rADbFegx+zYHz6cce0oawrD4ZMzcs/fLEB4HN8+Kg7Nc2w79NwJVaGH3GukD1J
gNkWzNqt+DZN8+/b/c3Jc5T2fycy6qE9+5KiXbSPDK6KjZ+YM9ORPL5rBWopMpMl+v6DdKV0SoTH
lNf+xRr4rurAW7Ho/IcN/gAR4P1leZEkVLk4/Dt7M5ybiQVjt3kmksVLJhSFpovSSzUKGRThi6FF
e5g+2Dc81TUj+T4FpjeCPOMxUNbTLouM80ZHGABsy77tCRd0abX3BNaAR4dQ6azztPm4c3jWXUdu
ttXLfvpt58g3hYmj9ps0cnxXIZuFBtZ43UN6mmBchwIO3OzH5NVynf6N29YSGTBYGUXx2KROFwAv
TUA5FAgWIUz1bUoW9oBhtLUutP6/uxIbfhPjaGFa+87tV0lZSzGndKNhB3sOryHk8Jilx8tkrtMI
q+Ycc/rMQZMDizGfqFg5LZNmAyKRnIChA8B97wb65sHpW20SelX9MKNb586OY2irQk6u10RT9I21
jW5b0wfR54xMfJ15Eg2xxeFgoA+e2FsxF7IlK+WWDE5GEoGPfK9F8wnGWRWg35DNBLUphT+NYfuK
MzNnHYwMAg9eOWlJX/lEQqgrZdexYGuMyoeDPfhM2p1GhlRarWeQ9730BWcZth/0QGJ4Xh/FFAd5
l+mdDZFnLh4e6VmIxC5UKNLOp3FLG0uPcEj75IMXq72eVYoDF6te3vtggDDpOlNeGCISfbZ+L0L5
B01zZaqzFxJlXDtZRarB5z0vymZTDWPPvvTM0gTc3yAGRjhExP2gU/dMNxilOJK/PVXYzXduoNd3
Q6snMBIFlXz019uUW1POlRgJnR0EpTsjLepu4yROlLdDh89A/iQul0ucx/9bdIk5nJMKZ7k6hIos
IHkNeruaHYwu21EW8bmACipuWEhKRtmKDhEcfk0ifmk3S8XQuyNv9bVYGlKxmwgJdbKYF7/IchmY
kFCWRETqDqX5qXVG9w3/qA8++9N15YJ1ya91gegXcx0TPvB1RzHmcbnVzvbUzlTE2q1B9DepN1qa
ahrIocPMh4pGdREIuvRG8lcatOWesglZ8V4zZupBX/G+e5Pg731w70PbJNMPvexOXD7UOfsOLQhM
zGn1BwFuJinuGYidKAG28Z0NzUbFpUElUE9O6moSEgPcH7K99+lJyejUJv0tCVZ8SeRRAD9n8Qs8
dYgzOzVm09VukpAHylX8o3EzgbrMG5yg345YdIkV+aan9yROo7knx2fXS+I3uYBBsh1JsFe2k0dw
2jpdJt0Meahhf3KXOVM6OQmqhAwWe5il06y8dAiJBOqNZ0sxY8APN3jAdmzQC8BnGABLZZVJ05h4
hvOM6T4u5O20dB2mQbkntVRrbffxRhyYM0c31KnF/YXq6/mE9VAHYi6//n2YsgmDpua9TtG8tbb2
QzmwuQiEVSs56WF5nQwtcUFXFS/Q7cdxC1FaA9Iudg6/oqaC2JfkWOvo7RIt1tAz8knbnJO3neRi
wJAK8Vl7f6+hZ7Z8dGRePoNRyMbOyUuN3rHMWKYgp2cnIEK9Bz2A08zLS52W96xyyoOSPAJq1ZOp
ufY/GnaVhDUZPmAXwkpXkDiY2GTdymi9p/i2dZgKoGaJWYSUAYEDcB7meDn1gZ42f+kH6MzRxqcT
n078BU2M8dWBvSdkI8g+x0wwh5zSdgxfmR8yUDYxRonkT/gc9lgYvjbF8p21JsXdKS+HgJ8A/wiK
L0kxT1UtUWS2XXGhK6eGOjHXd0xBQrWzVuzg3oe99pPDw4U0gO61KKklZjUh3zTNjgDPvpScBq0b
ZA4Cd3qXN1hsvRvkE8ITu8MKWw2/QBK6kuF/4KVcTg7iJCcPIpqioXdffQmnLjmpn3+bTj1tWYtZ
8Qq8kUr8cnKv4uLEXYtsWC533Q9npfxgzmCSc/7TFuSq7cj/d9a87y6FCIah33L0Fjk/F6KkA1P2
WZoBlJX9kFoDrBoKUKNMoVmGqURli3gKYb5IktRwte0pWkE0nxVjT9WcxWQNh40Eh54DQ9gveM+I
iJtcmfj/ZAd8Kie1ubtdFL4djsQ7vuKP/a9xm7Xvbkz4cpCeSlyPlI2IyT60WKMjX3/+oXM/q6zs
v3RH5SdMbWaoW2KNFHkaLjKSYRUncuG4+wM5tI/HBfSkqY3hGV5GOP++eTPw0PXhLMAQoLrMzpHa
UBtO5dRU7ybpI3Z5N2Ns5fWZUEvA6eeaeZpdavYDJ8/iKXaFcA11HbBesCAi/DCCW6gac4cphby9
TsQ5c7thIjNZztP+MawP21mn7GhjzcD/czXaC6vXpkf/8Rl1cyHh/8ca+yT/whb2QlCcyD3CdOBD
Dyz2iOgUktzHNg9+SuEz7J6agJlTJZ3KJSn9h8ZkqyIAntzRtd6XDWRimsRIHGyJgdCjgWjazA8r
IiUzleUiSA3+muMNgi74VwFbXk+K7qcIPZQw7AWiPSQKeX+jSrqZ6vKx3FQBF+pfHx1A1+sA6MQE
VdcyMPV4aE8sh3OFLud3mxMHa/2fk990CorAlzcZgZQDAy14ztMPId75czK7WGh5XnsBDL7p290S
7TtWq9pjiGWYMf87HjERpCYex1+4Myix9hTbAD/3p4JnOVJRptMz7ufuMlITP2Jgl3nep9uLkpTN
UIVLfbWHIKwO8EcMri4h2z+LKWTdCqCP+RLMGSAmf76jT+nkGCMSXueqLtwvJxiOxP8QMxi4M7mh
VKkZQjEbyTbVmvugrN7qF7a3sjloUx20U+IVvo+J4VCMZ7kZx7zID2FFwgu215ccpeLxYBSYerbb
CV+TYEnVWXoRojOy6hNNQs+94EAIdhLSa6Nb3a6Sqjk62YUvvQCWbJep/Rpz5W5sTKudvbOYxrqf
A4ehnYgeq5B+7G9QZTQPMlTTn3S3QBTMFN8pwHTz1rx/+zU4VqWviQMlL2PqWP9cp7CbhF9JUKTb
INOBh6kJIBdNCItf6rBtwnk0IkCjSA5HtmDc7Em4PqJBaB1z1pMd9tXb5wBEqhZrqDDMjdJsRW7W
z/ybc2gglvbv+Mc6UcE9W2TffKc5DD+7B6rEitWMzWxzRqmzxz7AUiNHWIQrbE+mjdvcghqjRGSF
xB5xVB7perIVlAIc7ZscZ7FoPAqltGP6gjUNQskyJkIwX9t+e0Wo25pnvrpSnNvcyJB/UrRSaaUv
2QUmoJqjw0ntS9tzpzmPoykQOb6ttHWwkKYVwRH2wb1Nz2DuN2wbnNGPhCF03LG4z2nUDDOTKrVd
SkM7p8qngJM28blEQ8IH50cqY/huprBsnvUicDdMlVSwKyhBOiV0/v3K21IM3lnli+5JrGxEXnBy
crbUUaAZe0+ErPeJe7RSPdiJ3Jz6dcbjTGp2CHHNi5exg6IhbOngZBln/2HA463O32T7Us8Ywa7N
vwH8hgqaODKS9qbeBoGyoDSEylC6EFVjUXqvn+QX+OdZqc+gnPPDzX0zH1XWTB0rB4epMcamMOoa
eJl4L2FdxaGUha4c1O9/febRNsh38HdJ/daczh8xNaKekfBicX+RHJVzWVZMrPwZcllNJQ/BaUlb
WsPmMtxN4yyFn4ssBCDZzWSS/KW03OmVIvtIRFLbkAN8iAxbGad6Dp0UR4Zsx0/9M4cSsVT/tzHL
Ub4/B1tKNQ24sHxQBYbVWYQPgqWFEIhyhQk2aNekyo3jkcnsxgja0RBczFJxHSUsaEQbOs8G6L6+
egqC69sD9ifF8cJbi/pAFALweoDTNBCdl5Ew008pfCTCXLR22JQNDTEydlyM7ObXLP/zvXSl6TXN
V/Lx3OE22JD+EzfT83Qh141DEIn4mq2MO5fxIVZ65TQoAVRH4/SXdlOqMaEEG+DhEg05MdYRTz0c
mSiuRUTPhu70WzKFfUdgTV585Mhn4mbsvhPBKa0686pL3QBzTpSr4nYOnJjABS5uPtij3Ymbd8I2
VqQlg38VYRDQt5BpAzWG49rZNXYufCb8RKqlNsaqiXzMo6JbwZzpDleVo8I/4jBzmQAyjrx0BAxH
WuaYflf0JDrM8bw/NG9BGD4SQ2WiIfHx3Z4F3Q47UoyEbqq0XxEESPXg7F9JeeIjEK3GB6TPCyl+
PggOifXRGVB/fI4+a4bqb10iwun76gI6+A8V0KuHf1WRJdeMsMLG5HFfuO1OAbqtkfRrwVLjNeYS
gmuZblmxqjv52JxbU2VWgqwv9u4L7y321DjK9ZjcawVApnu/5o8EzX0Z1juyPZDeMR6B6+XKV29d
RVIgf+qNM7kRYeqYheF/mBZr6yzwaAbIACjz043JKxcaKzTiwtIAqM1YE9JFmCs2/0UxezOIWPyc
7iInS/oX0ZABeKz6gnPPp8TdcdECBFRIm5Sn5MBQTdShPdX0JszrndW8YCaHBQb6ZbNQghzd23uQ
JOen+Bm5ddbLFdQaD8gmW8lQnXmp6ZnCG/NClOGT5cxmBLNSkoZOHxQ6EUj/k3dCV7WzMThe1trW
Nm2OwedZWV6X/D2Kgf8HDHyHz3/hdIO3S3AT6IYWi3B7oRHrGGUL3adcSAEXXkkyGsK0y5AF7dS5
h0Dls+oHPxleeBJxqmYk6UqfRoJdd8EA/S15sM4X4+xX3z8wt0BA+mCFfXvTdFYVhD2xZrbaOHea
eclNWlM2DzQL1ebBnS5O3ysBHgKQnVENLOuu3KOSAOU/bqxtK+zKSoe5KpGHRUH1QWZUhDh9TTq/
5dFm7gTeo+uoYLDPE8Ny7W0PitOPjroXOhXgAM4eugd6XTS3DS+1QyAWNbExIOiB9qQ1rF+3Nr2m
tZJWGA8GXomkhatduJufHEHTksDlJsT0Oeu2MPyR/1XhapYatZrh0tFoZmpdhTMdVKufmVN4PWx+
L+KGd8mnOX52krdk7Si5dlu5uvHd7f+yFShJ0M6XF4X5xf3hoxAK2CmizP7qvp2sSBLKKEE0Iu40
c08M68idi9EmlXE7Ey04OsxYLKvxcusFxK+wS/FrGM2k8jsXjJ11+S7AddUOfZmeIBidN5jKTlfm
sdplCM+E9Rez3UjR5uYY4eLEc0DElUl7eQkgiLbXzNDuwcfOqVeLKDmXXD9bra2vEsKJFh6RWBEC
PCuAyOSxiSDGQw1uusNo1JmJSiefvwQ6KO21yRZRfnFxTQMkx0nUPwb1tab4UgXJCRsRhUHuTHYY
LB421b4wMxassnW4TNMrdHV5vy2RhIcSvySNouzJh7/CdWFQ5xARSy+/byjTnGVvi4c4m5hvP1BA
mFpK/PiYVFQglmVvdP+UohCGgVhmfoopSgTFgI4R/WaX3//okUz3j69XAmmFdes/FpBYu2KqxGox
PTUN93LCtOsL9oaMeew/NzHPXuEta635SQ9vALg9AJzlejwr/k/JHzB7G0sfQI7AHdmTK+XWJv/1
MoZfsGcG8E2s1euhkTGgnwtrY+lLG/7hW2UWQheNfHc9zpUCUQPdZM05+CrKfjDYlq4LegXtepKX
iUtuHiSFsr+zvTggxSBXc9W3fd6va6Fx+lZR2AU6DA4zAaIT+TVC9CQUQeR2VCZtNoKoMN6NDSAJ
kcMFJVOSkq9bQJ0WuLDOcRbLhblhqcSGNkz6yvP702JK5SPScJfcbpMecfYMoyeo2tNwbcCIALJk
VxHvvQIqU0LSN2NqLIFP8WEr4KE3x/dPGBP2t/kQJzteZCz3XD3iJUDJqOIns+PibJq8I4XLE7UT
8l3wN1wwqRZ9OoR7OCVcL6usB8Zw9XHXd/Myl1Tk54GklnmkHbMBN4ca4+4Oe/4baNI/hJnOFmRw
z47fNrVe46GKJ9ELLTm2f2D9OvXp0hUZRS2sbkDrC4rr5FWMF3KKtm0SX1jRmcm6kCw97sIZ1beK
vwALgDjSFc/lglIbcWk1fjSwp5J1j0UAkeug0W9n75Tv/Bv0BNBQI4j8pEse6wKjvDJTEamHwnyb
pBgtt0Gv19xvoAMvI40KEGsQYdB01O3oWcoaW89mwIgQucMD+PFkEmmK2q02TLUhbwp5eggpNL0n
cPrFvP4eJQ3di59GblR8vBk7aQoI0BVfoz30BApc7evIS5UH2Op4nRW7w8CV3irWL4XwqZPMV/6g
w0Q8Wozu9dQ5hTdT3EjY/qRqSXxe7eZq3Xeb+WfcMzcMvsCt/Kzc8jAZvGzTm4jBeUQp2dDVjFdw
CS2nEZuY9MrNpYFD5kjaRQTkemYj7btWnXt1yzoARYzMvYgLOGN4gAuxE7eRDDe0pecLfCQG3TK9
BzJKiJZozQfKnt8AOE5mz55Md7gIajtKIsLZR7hNIEnW950/xun3TO0/9FFddpxOdtj/O9nVyCSy
hTn2CcsqCS3pX1z5rf2BeQzW0h4U8jmBrh2adQKEItgLtZekbZVMStMBmx6yOUCEN32EJvbmoYaa
aDjcep680zptg+CigsCHjMZ6uAvg52/jmoQ2g+gTeyCfY/tHTwP8CzGMSfFBEpD6dUQayQqVie6p
52DcbR5fH7LiNpQuRTWqw3ifArvNbRULwh4XSVywzjD/YsThVuIc0038BVFAP3JszaqnZXpik5gw
SQOibIkwaC4yVkjf8WRZdrPzIzypTh/lDKeC9eA0cb6e4KYbsPhkicukRYjm8BAVh7M8UguJqTjl
I6SCNfap/gJZ4ULY5N9SB5fxsoLTmOaw1/XPMA9i4EJrm5LDnQ3Lo5GgegjJaSehQpPy9UQ5tmTv
QgoIWK4RkMjPrAuFJWCNaSkTsdXUsHdzq47l5CXEbvgmvkCM6m7yBrK9kA+8MegNUizos6pkjKWd
nVJ/2UfX6ZUD0C1t2a7s2N1+77z1Io7F5ukLVvGiY4Pk5cfIolNBjzrwGD8//n4d0AYq1o9ME09A
f0Vav73NN3aS/nKtNpjpZPKWqMPjliiw4QOiq8FPum7GlNLawQloP8CIDbUI9Xfu8KV9tdpg+zt+
gZww4Kqs5kRSLDGWlVANiM42mma5OhDs7mrDVBvV21fka83Dxsc0hGw4nUBmyAt87Ago/lLAjL6Y
/dJSJQ2p/rVju6QDRyPKtwyE/3Z9zV2L2mgjmB/7Z5DlXfYy1IxWmKaGgtbirq3aM0uvA6xxM765
IeKnIz5CTiOZfheGptQjJQBFJcafUtRJQsWQSxFQP/N51IFqRV/q4GHg8H5QujN0sXW+KIbAHoUa
7khVJt6e37rSGf3G8CufQZdfQvVVe2HM9ytDm59CBMxSdsAeMV+sVwZ61cEAedUu+HL4RPpN+9cN
pi6yecvQxqk6z5kxwWF8v8Q2QHKoGqWZmmVEZxfnn6jdohVs27eP7HB6dv1ouciHlC6gzd7co/Er
+OIKHv1B+By2W9a4vTw4/6zIQ5BhzAhykwgEM8dETRVuBZ5PWCbsfFSINc/6uuI/9boOO/Nmc1ZC
8OpgMtjgd/31b8erStsnue7TBKhxGEkTqL/op/rdTRtIJCoTWE7O8GVHLmj0GNpJYsoFZyUVl2Kp
n4V7LTAqPJiJj+k1MiU+C2qLcgXj7xgwj8n/gB5qOxdw4slmyhP6XACMmBISLIxTLYS+ovpGh4L5
W/LZapylZO2dlhhXM5FVk2WtlyaMvASyO6rXzaZ4bgM4roIcXS2q4gG/aGSQ5Zm3vlg687EaFgyK
V7MlZZ21KB0uSud5091Yfd1M55QvkannHgQT5xo9HrbDWNh2UGsXJW3ajvTn7nMyhYkMTbjeeJcq
QrUtptEF932J1PWcjQW/y8SEaqg7gFlVtnmgKvz0ZbN3s8t2X5J87iH/hc4lis7vQJPs5KCwwVqf
02pAEkpBpNKpNYX3PngLf3AHkoAZ8eZRMCAZkBc/LpzV9OlLmFOBle2QQL5GCxYawgC26QcxNec0
/bxzFC7B2ZBDCcE11GELIdZy2S+8zNpqDwnK6Gb/kcw7pTV7/u7UDnvLynPepz1AWTg7K81YOzIZ
ab0RfAw5Rx8Y/3Deds1DiQ0K3VPj03bJz9k7GsNtchvwyy241eWSHFZ6Kv4KsBOZj3fPTLjhIEcd
3M8hjI2ALzWjhEgOdodlm32U+hFLhCDgxj/d6VvGX6ZVE2u6DPEOYFXPRpKWGiQ7PwiXTvZHwQsw
r3ivLLoR1vL/pHMDifyumQCrZ/oMAViJdkCey9cC+73hceflLZUHj3dBxFKp53QRdT8QHD54EUbi
8Yxnhcdrj/sYmgurbrOXgySliC+4jRj/26caXeXf5iaum9JrCBvkHGnzLfrjoMxZnhkvV9rHX01p
kVr7DEDddW9ZQ7BnybyCQXN6ifgVc/1HRQcy4MDs1KgTDnYcZ+a9nRrv500W16qflmAZpjGUkd38
YZ1XCjzU3glDWDN7N2HV1QuCn6qfNBXjuTGT/OcyRz3tR7Y8OBtqGF4L2h7so7d9XSGprFxd1oMi
zLitTsh5bt1yGaRSjw+pQBE1j6CMUS+LVtGz4rjglVFY35mpWZfj1DmiPkWvdzVippL3utc55QXq
EWK9wKV3ANQkUJ9b2aWFn1QokzUlfM0o3sQsrL4S94JD2/btzsUQE4AgmLWekfSdN/G/JvAV7W41
IdBcRVFpEOSGYfDTnnbL1esjTjoeBNNw6uL1L0gDv66KqdV8vknytT06WpphEvW38J+N7On65cz3
YC4m5yFoWEwxX2QfjVwzLVgipojcwdTIMLTKtDvBYLIGFLSOgyUux2PKL706027y/OdXRCOkL7Em
/d5QEukRsBd67asMV220ogw0/8Bw7lKHEps3+xLlI7b1VKN3SJ6Dvkm9fD1zml4CDJjCPwjZJNe+
MrPbEpGTfvuYozU1sBvU4WPPzhf9uVsWxTOJ+TUPq7lydaHzoRd/6Mxy+LZqVkhJ4l2uxiw2e15/
B8mwm1MZc3JYjIZwI81Nc6fIRU/Sy9KlJfmSqfOJLCg3sjxRmqWK3AGkhGOhAuyuhatJrRPJtjwY
aRWZPary19lwC9nTozBJr0XCKLEc9soHrJm+PfoBQ+cnh7FLnBMbZXFZnyTdekUAv0n1vYbhkta9
FJv+JYqj/+Z3gakmNzD06v561+fY1Orr3orFg5rWjN7EtrkOqKKWudqYayipOPPLXd9ONKnQFpiE
TrrHEeWrlDgt11Cj3N6ihetlePZ6GeyEN5rVnZrofYqbk9aArq5/kGKqeB7p6gz6ZUZrz43i5BNT
9Jihc/FpLgtg7EC05Fpzb3s7KCE8tyGSBWjCaTbAedBkEF1J5g9/eaF6OAuKPIMtaqw0RTzbjaHt
QMVbtIZB2oHEV35FIilgNUns5V5LYuAMtI1ElF/vJYdd2/W6tIDbXcR5rK37oPFY+LuZgZEUpgye
WlAUgrdvROUNvfK7BygKVDZqnJMKmhE9r7XzFoLDdRV3CR7pQWDJTFUzv+t05Hhhr3/GYNYX+RgS
fs1kmYjPcFyH+tlw6AkF6iEqXzBtTCIl7aQZ1W4HFaN8W8iskipXv/wGLoaLKeES4FP17LZkxD9i
RuaXBE/ggx9MIG89IhcFtmAIt1Z6ZTLxq8LUHXOSvtueaEWg+wUFX9qTBYKwXXPWNhR7GAQknXhq
SgU5k6q9hFv0z0anszcXocbn/KbEQdDgJznBmRWWXaDeWOujHVfESru4kxQvjkknozwC3voe9iTx
mGwmlE03ae0UqVUpedL1cFEVLQdSnmDxktS+Ug9iexzIHdlvD2+fQNL/qrvy/XsfjqnUFN8xNc3T
SYJYP+tdS/fKt6L3ZkWY4lwLFTdaz+XMcACH3AmdJTpc59BCIqmUx2XktQItcWPyVBM9M4q94CFq
D2LAgUXvVXniCxI7WJvGEiGYpG3VnTj0CdvdaEie5YQo+U0b5ooUz2tuhnyI5K1DPAGmcJLc2lIh
Waj1HH2ZgVW/dijxyjpNhoPXKQyp0LvbNQyh6CnRt6+mG9WiV0cS1xXWGQJTTvnKn6p0mLvExqnB
ATAGznx5pjXT1TKKy/25bN4sfNF4HARE5ChVvSfA/vFq2pTFSmDPFrhNn3tQCKtS0VjLm6+eyWGC
Pa8AdHpys9YE9pIL0sec+XATB1mQsO0oGCM+nOvLLvCDRoHHSljYOXiZzBcCw7wmxkGKehPocUzJ
G5XlRlT6GejkRNdAYWZTu9AA2TKP/R1RvGTKtEYQCJ0+MyALrCcCrORIgdmAWnPJnDTlFYaFXlzX
cyjvXV+nEVbDG/3O6TY+JuNHCsrstODy7tAoL0ArB74he/a/fIxZgWhPAkjDJ3Q1zQqU7/uIzNjj
MWezvr1+AzBS9tVPocQFGpjVX12QjHMHJj89dXiFAQwb8ZAp5OI7EbnFZP1w5iik9XSbCMULVpL9
hYUfoVmKphG5VDf+18gtkyT9IR/PNXRB+fMsdYu8eTiFSg6ZTAQHbHrcpRgNX3CKIDlMYEBUyQBk
7Ao2kVmWtpozlqUdevRIu2/e1WoT30oXcdnLO8XreWtyfr6NA4TP1JrlMJBYE4+9X3x8ovmuG2SG
7OaLXkOPIndf76dznontkcoAmykaxhLA84wiA1GoBXXd9q4DZfmyju+Cl69CwS129JGLIbE4NkJO
a5IvPzXKt2WETcpY4Ywt6wswB+FpZDz+pHarwzJ4IskntDPMoQgGN5pOP9MoXDBFQIos/f3s6ecp
fl2or64DtK8oySPS2/3ubFkr+4ULmIaPKH5WkBqDN5SM1uiociHk7yPvOvu00ufcWA7gIqSwsJCg
bPzh25ubh145OpgVXjjb9Mp4ICgLKJv8qKxMQ5pfRnooO5PeDOFYVkkPuqp4kM+K/MNFoe8Z5lHA
PxpVlIW28Oleww8J50fmLyGeEOU7TouJCpfZhGjoTMnOL6cujoztbiiYnRreGE6owmoSLoMG2Z08
wr4ZdS/O3J8obXBUY/L4u5/jr+ivebr/DG6C4JtFpFCpUGdO9lAoSnQi0kjrLFlPMd7hUUkuWJit
9f3X+/40Uyv+QXMDvB+1/02jqi22B8aCL7rJNJ5l7Y6TP72CdM8KpWkOi+o2+FL7+4vHpqiRcPb2
pLEB7lAVgtA7d24z5Vvkdrc2usBk0/G9bAUFAShDmJmcyboxCOObLqx07D+fem3aTyLqs3vBfmqD
0py6TAeOqO9ivWUPcM0DB+cou/2F5FozBOGHkcDwjhNe8wyTYaFeD+dPwKK4usJsM4ls0JdpRRea
b5y/7uVwZEleclNGzzD0J7EDvVe1aPZo1pWMrzDzjhrS7VznWDO5VyBOOQrp6IQXdFZ/k1ifL4FT
jQN+ragUJ+RhU64NtjIa+yF/l9iTkIYFlB04zAuN1FY5ImyVIMOmmowsRNTFjv1TdAtCYZdGbwMe
2pIV1bb/nc/D0y0f7pS+TqF/GLOvIIasQmFMkA/2fl5iTwjwLiREhSj1kBsQbD0bQtjzEun4sW9o
PtDB4dKA3yyILdfLWN3T84Vh86k55WcPkuJEKgxkcbWpsQuHLcW587Hllrxjz4AGIuj7s3aKYUFX
UbLvF9h0S1ALCkuHMHf8KGOaE5w07tgOCahVrsPNgObV0wpJBh8YYsLmOVsKhTg6rXrnDuCX5wwp
WvexP5jvIn8irOJ3MGx/Ghz6MnxBRV5ms/9pIgppGwzdW3g9bx2aneAs4ggLrzHpJ5eXF47R1QLg
btuJdta+1Hg5Fd7bPzD9ZgdDqI9hpm2eiNAncm7vFX3sbIHTsoNwX9MXRaJruhHWqCdqadz+GDp+
K0gRwySYmNm1dTyfiwNDTwnrWjPmLNudmvQFepz9o5kCglf9JxWsPkjnldH6E9wqsDTSwO29FYZF
C/OwngOVbKJqvonxhk3hjcZ11iwRf+tDqd9BpHKIRkhxHxz9wkjiX6qSSRO16r0fwYrNxmF6HWiT
Wt8NLMRN0DP9Qe/BpfKBDmIxa4IiJT+3TC6FW+SFQ6mmB0L8spZCNYndWPPUGAqumRsiUmGw7iwM
xac9x/MThqFerMTCQLDTpEIqzFH1B5s04mPYv/b4aNTkYptv/QqqPlon8mW2tLF98mPNWGh56/do
S8UMyXFjHf23SIw6jj5fqz18oXSsgWtj0o7s51y1zsF3JB5kYIBc336laOd/9CR+4D8AZcj3ARrj
gG1NqUmJpVTXaLuWN62EAQCD8tcNP/v7LRU1Q9nAwwPpEpQKGmhhYT4THeF4UhH/OY2oUKqAsj19
prD7mcNWpTuLWAXrxmtu58uXMQlW5q6UbKrQ8E/PPglIUxaOCwrJ4OER0rA+CDRcRFrU0HM8cQS0
YOYwk02eFNHgVHTkiKMfP3MpRhLJvBZuUip2ipodIegN8bUYHECn9fdQtC572HbZXZgH9S5NqJpF
i+zlTqlePtLDPx6GSCOFgnE/5cMkviCXDzPnsMmSsclf7/8+766+zzUKBRVB3YhomV50ZQQNkR0B
lFL6mGHlLSiBEamjnZW0g0U+E6yQPq2Ii7UHdrbOKmYMThkH/jn2ke0nakF/rZyq+adbVry4uUAG
pizUnCXOL2UQdnGxb79MCc1LuzN0uoVnAtcsaZ9j8U7csaF9JTMCh8hNs49XGibK3puc6ajJIjUG
mualGiCmg3EgEPVwseRvamAOzcjS25jSAJfkvRonyxSZOSI8unNkc68wF2uggCbJdM/YcSHv7dT3
1ZBrk0MeQuAbWkvtjzHX09SMA4T4kBUbIeEjf+ywGJdip6i8QafFC/IGg0FO95Ao9j7HrhGL2y+s
d97XVNpes3Wbt+90jrvMjTKyQ829iXm5f8FPLWvUnrIOLq2Fsi5j+sODq5OHlAh1pbvlhHBtv2S6
UF77iCGeIfCbhN0l3iM+iFWjGpKREYJrKzrvGNDGB3F3vQFx73tZJIyx8dGSPdPeXM589at9jZ73
8xMgjZU3KTF0d074o96AoXWf4zK3nfqdwaL1yxRwxnsJBLe1gbxo7zS3evQ2nIrER590izfPK2cc
BlLCRz6hikmIG3tE3lpX/XLwcBT2y2ha+4hCJ2P/YzUUEdqmGKKX+KbXNFMwI7AGHE6L+PI6EipV
xvlyC/y6jXHwOYc3oEx7ykAXzAsFpgkpoHyLnu/sGq47DQoL+eu2OmHpYv9hSLEt3zoqU0f/sGJi
bwBMfon4TLY5kZr/inoKK9sAnHeippYnWf+u2haix7iLVPMLzfBZHTZIFX3mONAn2lMr+QPpL4uO
97tBXRqUTqna0552lqsqw31rSJsUwgrE3YEovmM9PFTpRV3x01iz5/4o0scUhwYIOCx/616Oekr/
m6nJ94/cNGwqVo85w6RyhBklUY8etp4JW2NGpPzRpFZzq/U2BRaq+hSdkjj/FzFQqa44fYhz3mZi
Twwyj4qLnaQhApFzBQrs6EIH+W2t+/dp1/iMBhE1a41JzbUsiUSeFXKVQ1RNezZOPTydNyki7Cl+
8gi/lMHiSIjaXUwLHINgmmTMbQzEWY9jUEFlwt1XfyzMkvhXv4xO/o0wP5G5thRPugYo9y2is6LF
oCY7e1t+gifQbRlBCQedeXazQO6rO8zfMN7PeRMKxMqxyWXVRGYJiXbbdACEVRtz4iuhJ5CwJmjF
0p+WFRM5MkUF7kKvpf48WBq804cJpsgCpAOpF1xCusQ3y6SWvWCz3vVjLLNG/p0qIMwAczvajZ2x
hbM9JtS3lrSOo4rLyHoZuJ4VOXGuVnbMqHAxNYQRaNaXaT4Mi9IfwnAAejFnxn04vjNBiqAe/Qvz
whtvX01KjzkjqoqZXvrzIu20KRlU5jz0YQLjx774f7jSwE7yfd/e67r/R0BcQws85lfsK3u4yY3f
OZvTnUFpE74TW/roNuAJhbCLWgV0VP3Lu0hzSZo50TreQnNKnFQXqXCJszqCaaGEWyHHQbRJ6caT
gVd3xAGIprz+OVgtt85nVshNxuWJu6IaFYSz0z66xW5lvWDiDl4iOuVQMWptlr4eTiTjcamTvPXu
LFNAbB+jlGcp3vbFGLKCXAxqJC39frOQ6QnGjnl1iOMlOLBlbBZrDr0IXH/aPvHJaEgJ1SI+5hyM
1ZMbLA3c7vuGwN1OEh4qFi6f5LntDfvYWqrdEMg9V0jUGcZzh8GYjf9dR3jnBmt2RYHXJ6V0J6+Q
ogBnm/74vBICP9NfciygbawlPziYOn6WSo/ysQycm713ntCJjxi84ObSjgN7o8sk1yehX2XYe06O
02PH+O0IGhf0gqaRfSsDGv7pPpzX6RL8IGDb5Zk5EtoIfz9ZQaRJT2zp+vKvcmZ1oovBJtYA/eCu
9iGHTr3O1+QVJ5ryKrek+D0RhupW46zknV2pFcPmD3TE5DDUDiyMs/sUoDjI9QGA/j+rw/+wNfDV
JnTr4kQKgMGtSmpKHcX12OE0wbrXbJqyblOmJDbpCMnvPWQ3WdrkoASLFZlJbsKQPa/HTy7RYaB1
/gBXMK9Q/MS7Ttfcb5FPXlCfRXN/VO99HxdY0pcRd/Li2by+g7Qxbcp4pWVkudBUp8+YqZLCB492
BHkj29K3S95G9kHIZefMX+EdTCaWBpHrbhjfW/T8UUbi1/YgPqFfaT1xbUdMYPXWoliTSySHFoa7
QAlNMiEHMuMjU86QGCKWUzLtuLpVnH1lY/DkEYzbaSM0pqbVQURv38p0DuclOU5Q4An/TRfFnC7/
HLf3K4xgTtuHsFaUX16Psf7KklXDbpXEupUZMvkrSeF6fUwqZeVNh13sT4MEJFJ5AbuzMr6NOsFq
vlSU0Ubj2J/xhcAcRSBXjtYLsO/hbSbu2hyR9XXRQ8inJG0l3rUSIwT5ZcZTVNttGX2Nns6JQ+5u
zhUYinz5nfFZtgYeyItpTQ44zgFvY6taylypY0uVcQ0JTHVkWuoH1zFP5p6tyJVqtBsxMMX64pLT
Uql6JjsDKV7UfhRZlAm/39n9/kP9RQcLMNoivot3Matk9tk4P4obytyCrOIMiQfVXBOe2tWANUoL
LwuSVO/9X2Xq2htRobf6D/E3uYkRqQ+pAuLYrfhiPDK/o9y5+8a9VpI5Z7FpbofM2BVh2Wg3YnLN
g1aYo6cwqB8Z7/VfFi9dgcVTja6nZvrZRDjIbMTnp8Jf2rjy2x6OACC137QJNXcAbYRghgSDFjmM
16wBiaO3nGovJsaBw8BB2xB5dj5QKbso1Tztf5YeCotXFPVrMIxu8Det4Q7BO8kXk7n0Iu4K+P0x
+cAh+uio1oDlIkJKQD/kQoQ5htqLZoHFweU8MCaxbjhGUQykTF08etz7collThIbkuUY7+km8svF
/v8cEQcQIwmlw+rvbvr3p/fcUKdxk28H7n3Oua6UDtvt0R1j9YEweplq5vDZECJmN+MHCY2XHZUR
EyckO6YfYdkhPLf/H4cskdgNHcupvpKZRh5Vh7AN/wNFRDeleN8p1PVT0M12mt0ZXq2cdiP7wsUW
a4UvHYeOXeDDQDp/+TL2nTItxlyhSGY9MQzzICW9IsErVZ2uXJWFszznMge+h6USF1kfDDJN5Cb8
FGe2KJlHqIsH+wwNleTPJgaitCmtgYpAgLM2Q5YYmodvimvJQG2cztlMn5Enx0vFK4u8z2sCDYG5
wnalSWR83RqqcbmN90S6ZNs7w7gkT8NKQMiobEC1mk7NVGG5nrW6cObkQ3VfLte/DhoMmyhXpx5w
jkzn0nGMuLuLdtH3Lu/6QAnnDEhSrcdjCoSgCmUhppvNito8rJYD1lkG1zijCqyXEn3llIsv0Nz/
+iWqvShaXF1F1uorwDtYAhsecIF8QwRlemvhN5UXVaLHPoDZONmALuh+BaSHtr6SdXGwmlw0bZmR
rg12WUu0gb5GxwU+GhRWSzT2kVuE3z18kwNnuJT2PxVdLlhR4+U+mClma7kC87pa1yA7FdsuwSK0
/W9nP5inbqzKJVhr/uW2/CV4AHqNp/TCMtZrHnXGiBuzes8VH4Ia0zD3J8bNvAvoLgRBCHZi08KG
y634a28renYs14QxyisBCy7oRPYzF0LZV3xjXUcGncUS9bG9FEGRkpxb6gJhTH4XIWWIKGUmQ7GZ
A1YtNCQT86u1BTUNzwJLyFH7K5+zRbydR5n4EsaQa/02HRYtTHZaUPxrlO0daG3aA2xWmUcR1M6a
bCWNMC1FYsA9/UkEEZ0K6KJG1YuCu0gD8mZ+2hqKhNqWI1b2g1J2lgzRpfb7aFaXnT4uI59w7xRb
RFyUFpB9d9trLsJQMmNBz7nlWrOfcCHxBPuqGskzjnB1qwTZnC2xKv6nSaOrynb1SG/apSbz8xAS
LGBPaA8FnRxI0IKTNMBUh6Nx+sYl6COMTAKXY33cgJ/GlVVsw0zbs+S9fohQvSUDYXtsvf0h1Cl6
JdxhXv0LW3V+Ar06lxztpgCh4isMp5sJJlt3UbOUg1jiitvXttrwd9t8QAcZntQyVnclLH3qrY4g
jzkiKdTcIpuO4KGjPlw5hRWTU2lhqfL+mAdERNiTm1Z6s+RnCzVi7qhvj03qM/Wghp6uvLaUwEOa
uTo6m9uALLpMOVAM9yf8hrdkIOOTwMM1/fiP3hJv7IICWFhLemiWN2CRkNwI3fglqkNuzhW0kLUz
tApDT2ZdtjvhhsulY0h0L/1PANGxst5dCLR4Lf22/Iq8nLCAWhcI9rQ9wNLIb5o0sjO8N1zp7OyB
haciq+bYNUASCnEFj/3Z54FSWoeEdGfe4uXIDmLI7VyNNaYiD6/ar4SxJMDwmVmm6+UnlS0L7uEi
5rw0IxBU4VS9kkLtHHSpoXg0yKjpMGEj5SfgI2hHf5BWHRHvfGKms65DE3NAo8TahbbsbNunO5gq
cXjf1ZUTBgOA9VcjV0i8uDit8s8Na/VhThCl+y/WEJ9V8tpKjx3BsEvKpAST6j+YwL4sWfKAKAvp
fz2aXV9Vv1edjN4Oy1fAg74w1EwTbtzaF9/weLzvQwO/Bmg+xvgOpsY3ssTLwltuskkdCtpVqFc6
Ls2GDdb3yLcvG6bDfEKM7ymedVOIdGjWtyiI91GnlC9Q+b4E0qXL7tJcB5AlecbflUjXLZYIdsm6
VvR/Jmx/BnT8zBg4e+T7D2dIjH9CQmMha4wyauUmCWtm/iZSI3n/dPjUcUFbL88SoT13f0HVulTc
H7epYdTbnIMbAJrYpnzrXCqkIhoHONMUmxecyTZtVbblA7IqxL5PlyhDpKTehxQ9tmo0b1s0LIb1
YwcHSgySy3gU2XH7ZTIalKzj1Sq9n9xuIL65qER4gcBF5ojgk+duCS9w4ReTNo7FYH5fYcfTNz0M
6HdTmnvkn1hhRQIGj6C9IeeVCz8VU5AzvFaG5gCu2Kr+TtcDIYRA49Fasy/88IqpDyOXzlDR1/+u
6brEgrPBPXBuCS+ZO4TeP3dU11hm61I9dpqfYSEowaO4wTzesxIHItaL4CXtMBNA2WIXzj/d0DRG
TngIaBvYwO22uCNllJ77JXoLXdyAlFntV8KOtJBudv01/wYUl3vNjZXTlmE5dBc8fOwyw+46eaHE
0bo45NzNNtZw+n/75hBD5iyFeP8fhcnnzNtrq2qRMS08rfKrrsR0QWLcFsSewx/ZxG/YS2H0QpO/
AM2SV3SVYeIqCN0VyVKeG9LHf+h36UDzTJUPCotT8f4z+mald9s0KKwwTk/TLmWHM1edsTYloo42
vzRxGLWaDC3z1/iU9My5aIzKTCxa2dnw7uecd/E1q9csZtgr6CfWYL9yxMU8u0eSN278rj9jZL4i
ATmp+3z5ah85Op7g9W3SrO66xYQULtCIwDbOgU6T9FLdZJkZJ5BX6ez5BWYSKMH35BUEIJ+hINhW
hhypa0/quRmnT0AxlTThza3L101T9cjqWPlUftpi52Vb3RaqzFEoNglCnOsQmzr5WvQO/s2hSVBT
Fg4PiGgUMNqEuE7h9gcYV4qWjmp7hvGAEpdWtccCGyUeNrLiD4vxNZf8AQAahs0B69NBC/HaLUZF
eIQhlwmcVga9lQLTi9sKZuvLPp1b1GiH589NnJjcOR0heHwKN1wNYeriMHUBl3WBaU37XLNd3FHY
zyEJ9b9uffxawXv82+7+LaYy/bygIpErf6XwOJSyho+lM9TvCtzJwdPpeh0SP3aQZ5ygGy9JcuTP
YEuL3/LME5TDN09DktR/f0mVA1DpoN2P50AKC9ZXavV09hRkJ3p7SFGhN/D9H4wqCbB5Atj7bBdn
baQRY0TTZC9ErTvrFIvBKe8iMbsiZddiRdUPK6shPKjzp6j9lOxfU0JNhTQIkWbZVedVQhq75h+A
bubukaoW6By+CFdKu9aQrsc9ptR19jlHuKjm71/czHP0RHfcK2B0jREqeLYacciHndzJGEmgyePQ
mTdA3fKSbJ8F/OJmnOTrQmdISEz65IVlSMpJ2qWdPxvFfFcEWcXeiAGVTZ6b0Gb5kJqUxHSdaY2H
UthjG3RZczqWmQHTE/GH2+BuMliY3GIrucz/a06oiJ+ATWnaVEY08L66wHUUYIYkYUL8V6m5pprz
TDZa6+2mTunRjFbR2d1S5EbNGlKpN5dN7q3xabzxWVjNm+hFg6k6f+OeuhQZuhPtgcxhwDi/3M1K
rhRYC9V2I45N/xkLA4Yiizr+d5tL45tjF7jLbBn6e4a4X21t0eFCRDxVJeeoMBgSE3WJWiG2qsIC
WxbzYjxCE/bZvodPhjtcXz5KioqOElHuVJ+f9uuv1v2VxjsR0KPn5txAxoi4KY0BSh++ZKVhp8kw
GiC2OeHfw9RbaGSsoYFb+5udPimfY32hZHHpsv0NF2efG4k9ZcrU7c4F5NGK2WPn7r3MJe/M/DnA
TyLqkERJSGEYebNozZfP4ldXLNnWnnJGI3dC2DD7SjKRQbskFjXqi8MQ/udpsYtAJqwh+nxQWsXk
KH9xj6uB7DGhsTSL+oGxmUnZMbKJo9tzyN/Xn78ZduyzPOGM5U/R65ajnKx585KI9VPqltARG57k
Yi38zOE8vRkDfggfmVBF3xRdCD3ztPyIyEraf/6XFezYOD0V4PuobAd7v97cJ3bNheC9Nux/M4Dl
ukKxGbicLHDXcxprd5MTcYuFHngz8G5s3z73w3B1kAci4GzrqrYCYf32WvjNv8U2eQiEz/WuN56k
zU69rPHKA83z2xMjDXxppj0CBolKsPUOYys1n4yG/IVBk3Msibyavq6POHkIy9f9nzeoLs8bbEnB
knJP4A75zEZgLpvh90nQyaaoM+gfiUtN+gPtT74KRYZ9647S1CKDPyQjI54TMLlgt0/eItEwZT1x
V/YYSWVSuoLNz8r5+tYxIVwY85R43/9+lNO/r5z9Pq8kVDRVban8or3TBPVEr9vKAJBIYpltKfgd
BFOFAIaOEKNgwp/7MonkLvsAwLtguhdIv3tlc4mk8eEf8K1J5rtRV5g3QNzzGKKouafe5LDJu7wg
xRXDpyrbO+mctvctctVMqwO6HK0nmYUlrb4rlE/m950Hw8dgil2BVH03qNtpt3VSDS8JheqRv6Uh
JWorACz14HL+L+jeWdYdrVP2o9IqxJgiU/Na71IcOGhHh/IBeSfRyweoZ6kYo4vVZpm0KDqS/9Mv
Oo/ufvkbSltdfDav5rgbTLGt8uwRQfJK85+9cRdN/0/6BpWSTfn44lMI3dV9pqFHAsuQroqqpYQH
/kvNBzl3wB2/N15EtSdvCpoYLrcsKSXOiP8chk7YVoLMEDFKK8L/Vu0JPJmEV5Gljk6Og60Iknw7
ZTxAN1WDLLasaWOciRPNxmx1J0hDtfSR5udWgDzSiqxPgOpCRX9fanZtwxdxJ4R1H3CdptzaQR0M
QkNwAcjYXQxfn5STVqbMgYb5thWkf8Iy/bbnCFWormVmrNBuHmH9XajuuVtH3pGeYLw9KBHzj0S0
b3kHN6jadPyANcoL7Mboobg97r+MBOpIHg6EdhwFGwmYQdsh7wGkwjc/nixD5Ow5oPkqFSzu8A4K
9TkK+IBl40NRMFgMMeeku8Mmafy3mHB+0EyAekTfZjVYVCaOkc6UBd2cus1TrnKc635tjYjygE25
nrGRiM03Buop3L2hTP/xeISqzrJaZe90Mx+yEoKIyhYT2tgSohFJ4lCsnbjwy9Y74F4UGQbxkuvQ
g7w79UPf+Ju7+4Lnj8fTl0i6vQzYsbjTrFVh5uXT1Wgd8eMF3QdQnYgAjpaK8b1OlPIF8e5mU97G
FN3aUgS2cDU886/qYnbsEArs4YEDS4JDQ70qzMgZW9ZSLojek1EeSqv0bE2EUk5ds+xgcQ8CwZnj
CnTNMjHobMnWnrkVTAxWUrSYeCxoN9WO14NIklGnLwfdkxPia4dpBmIZDBDW3gXy/xqDdjtyNnqw
ADBra7DCe/n0C3h3nCaefpZLhHFF4daPVBDLy1q1OHYIvD66LLhpYf9ih99lU/PdSu4OnaG0xNyE
BbBBw/NBKm5ACck+T23O1Qhqi7UyLMrKdwqi2XUDzEJFp+Bk9ezcNpYyVgGvoKXlmXpscEj98iJq
XQdhwzb1PdsS2zKVC72P+cysFXvq5Cs4JQ5I6y/l+y8zZyJaviRxnVOnFRZ7TI46VD8X0GgEIXEC
I+YswJY6ijblTQmY3e8oURYzmmMRQfR8NgRlOhAbzwug8jZ5FxScgewtgmgOiv9Wxyvo1/wdHE7k
rauGWHkfSgP2WLv3GBpVRLEUzWuxDogwUEO4V0MKRh9arwZNp9JLJ7Jaze8sfIcS9+fmdZY94pzF
fg7nxl+5Ipuv/GbH3DBhP5tyYPEruTaBjOf1j+61Cs/k8U9sfZM0YAu68zqspGFBtN2TwJf8bDe5
ey7rQLtGStOpt8wnid65JQ45ZaYnyZu15aMsGAwmQAN3NF2FQhPPIDHhl6Bc2PtQ0eZLoOj4IhWK
c0Ys4KnrruYp+E1HpRy82rcoXdFPidAxaGskCyTFwRjgHZLD9C3bUUdxhNmtxqfL8bdlwdbkupyc
qZEXqEpa1TO3q65JUWM31LsD55Fh5bVyGWNVqCYyMbaJEesS6ke+PhEqyq8bLBoCPAsopY6Ggmw5
KIhpbUremYdy3jQCh52IReC2xDbMByEbp6MWgkBhlZ1Xl5qxiQWyDaKoqomyLXSgLCwK28jFm+nn
D1zeXepMWFYhcDZBEzZLyM0Il3sEXrTC/2Tn3fwOKE55IoSJutZ1ZEzB5jUBPEBpEV2XLuGudh+W
MdYMwqDnx9VrGYSX6ri6c+cGOy0KbAQmI+7D7RD9vlfkUapKvBeSyf7nnH22shyPSp6yPAIIiDcN
LQChInbuxL/Jj1jel58NQhd6ozrBNCtyDZbYxLV4erIiyhM8mZcLYB/9kOUssv41d6WZ2XWa28K3
ZVa39dPeCT8OWZdzfKYoltcfrzEJs/gBJds1QptdKQ2JM6E4xTjnv6EjNbRjHSKzFylQBMCrT4x1
nGaGVmTXUGvgIusYOhydJt44tJW3M7ZsW1zm5YJfxmGoQSIdkAcdlTvGPr4yRrKYbRXrWkkhqrNI
bV6BYckUffFJEi7s2MLK5ngN9+x2zeNh12NYUC44Dbootbdmu+DyGa1vqjL4kyEVq8GPnHkXil32
a0hEpLUfiivWH9Vx5ZVIAbR/n1dS9DpDed1yGPh+wJ7iNsJ9+ztvNYl/uHXuDPZSsevwjAs8DNlV
wmJEQ/h4nxEL0FdYFbGVuJ7o+cIFpPFrIOen/EZsbFQ1EVeGgbiQM8zbszqdtBZGIxZz9nWk2n6T
ozd/1Tnqwbc/sepzOgsOsHxSwBSZGSro//+k+WP5cyqVbYbMWKqBwO7AOesL2feuZKIwsuUV4vc6
rEDpLwmj2KdvS6ohB5CML4n83on1vaQjAGPVDQjv+xkZiZWuNOdvOzQeoxvlTMO6EVsLR6wpZxMr
AlKdYAHruMpUKW410sLlPT/eP7E0M0PPADcBH3H0cjtfpdUhsLz37dfYn+n/0nE/OEUfAggySHM5
Zjo3U/qHpNmaKD+hzME1QMXJoP9CZxi9fWsc2EeodQbZE+lh9vL7EX+NKFnQnN1GHZdeSKSlj8fN
8nfhXMyW7ofPBrekdAQL4EaH2B/HzdA8Ie0lonSE1ulECuui7v/HSJerAOeV3vkehycs5b6aroo8
xx1WWza547JsNjxBuCpD8aQjOhQWIGc96/M6bkzFYX1/CLmC1ic1Ppte4p01+//Y7IfZHUrRUkqQ
5CwhrpBELnNsXfpicfRFPCAOjbzmi5kMf34YM+fSgQciCSPBP9cmnN6Ug9Pj7TW5NqJiL8UnhpWI
1AyN0C7sKcLxyzy8osXXLiLVyJbz8/uY2MIEQsN7wBdHCJDqQIxVLDt4npdoRFLm/Gsxa5hZVaYC
ggij8W6kp4dvVTi5uBQ0N4PX4P71fEGSjcK9fZrvD8XBGdKyHXlwbR0kW47KZPbYin/hDbvqWWVe
vVwmc8udqvGJS2UgCSXlS7EhEmFWV3o9bjHghUjRq/h7mKsZk3GkAXSwC9l9rBO814bwm7pQmulF
JxCViXjvVtv+chmVkdzqrBtTHhKDDGRwEpo+u1ZlBrsCSlG4YSs4ykTylOoRbTCr96FiHKcljij3
y1C+QlrWPZRzsAk8HEOus5oIVCnCBSiaVANvXWE8V8sC/BcbqOp3Mfnc0pWfWgvOQtpl3j+iPgoS
cbR1iwJjUe1u1OAvhoc7f72kdHyh2Kf2NJTGXoKWuZ7WJe5nXYjRU2JxK7surBvcqHEpA9SkNFHD
SUy6y5QCQxHuYe54gEF6dwre3mQMgCuSReH9B6zygRUmysm6z5yDtSGvxQz6bO2pIl4Og08g+sNT
4Q3fWN9hXC1P/7chiXEPZuCg2aDB0c57hgiAnv+bIIxDiMc81XYrMGOq8T/Nr+YT4EBu+02rdk80
Y/vjgVb4qTRcauWS1fY/heltIzbovZozBYhfS7nm2JilbJ1+j0Gant2szE5nULABDLVssIuLPqjg
66qOPso1Njg9sX3zMXV06khld/KzRcdAvl3otwWAXP7BIgus7KhsE4tn0prgyAM7624nB0TzeMi/
R9TpJUe7kHALTk8HscxeKvPlz3AzagPDty12IOezotXVBwqK65X+fbpTUTEcZuiUFv5Iekc7gw4K
H/SI21JOwG/fYJ/PSPN2fqnWT33nr6yvNfjjANu0PVCmr1382yIV0ky9uYP4jyXHqw7jyAjSOvVW
/fJxLL3eD4kytqt+anINC3uedZPH+QI1GJ0lWLvwI4lT3ppr/YPMpzOf6EPsJErKPDjvmOm4WT1z
SNwAU0VYqrNY0ZeD4TpD3fVFe2VH2paEf00ALIFa5G2QG0stZtVwWPsiGtufV4F4bxlel2vr9lQu
nOsJRs6+FWxy6QmPWcPTAROItzhqh/dHx9Hgot1LLJz5zFmqpVCFsOzQEJypaWc40spvY8A63kAl
oHY9vkgERmec5L7aJI6tUJQQg81zJb9fj/dBc5OXEFSH3fvYMozMQjMCp/NVrPO8y4EUScZcV9mZ
rAoqX2VsJsxc/1uFUtZxVZFRpXGkytaV6yIInjSMusUkeFjoKQhhgk9IoBX2pIRPK9A+S9/4GXFc
UnfB5IdUA9Ab5uLEjM/g3Qsjh+onHNUOF3adYYEtWyRe+whgjJlPGXi0Qybe2vdd3aAdGf1dCPU3
HTKjRyzbwwvywMR+340wvSEhbcxpmjghLSBqGwJGJk7WKZtL9MgOJ3WpQ54yYGE102o7OvG3uXCt
Lat+MJteRbdmzmEi+k0FQuftwQIsQnQv76WbYdBodsLnWDtnrNqgYmLkaw0ohQ7TO+sjOwkW2DJ1
v6O9osg/gCrSalCYKPmCYUrSzcENfNkVMwWyB4fsBDXFjMxEa/6Dk0tLwKOswTVBQLos+HhqCbK/
08TH7AttB6dpuLHGFrHlesibvxCX6OMyHLwk0tYSJZN4h7Nf11CycAE+5VjVCc/7vZ/Q5t07y3Uy
32y9Gf60Mljn2KQP/stUdcwy/iSModWS+e/4W7sdTVWNOzjpR/TjxXB8Yp0dcPeym+rq4Dcr4DYE
iqnVEAQBEPyfY+9Oyyqg5DxQps1L5PV0zd27r5GDPYZMZHZkctKZ1ddPvhTvk3cvX8CPN21nR9EA
zHwdPKmDZ/0iW5sCPqN/J+B+4J5EKTFZo7EpXcLOToVJ2yOfCw0PhQv7D3etdryU88zrdBQqEyQA
pAOe8aKCNvs0BZskJW/OVp3Q6Zi93QGzuC4OrbG/Mk1XN5gwy2dSD1h/wZOt1kcm0H+nEVnpo32D
nDNvz58f8aTnTZ3EIomiL9lGSfQ58QbQqDfiOvdyzbbBLCPG266yXFiWdhf1Ow7teH1GV6mzn8Nr
vxXoTaiTo19rZRXMa2220C+nbCyxLD6SfI7Qxafu1lpoyhMTbm2tNr1xEEARyIJJT25GwZAAAJNz
y7OuJXT60k7EJbVyGEHwPrezcsbtNJLWEwpqOlxwyu83D+isBihS3XpWYh8Cf/di1KO587IghNI4
VH1KZW8av/2VMtIo/07w5cQV7EG+ty9HvrEIuCoocRho14IjomzhDrHSvIqpMxNzEwenQ3TGfVto
xaNARFjhmru4xCRVmuLYQwo2c/gL6nKNqIad28IKL1kQB4UvdsfzIzOfIFlWUyGiNVObf69+I0Mx
ioGydsofcf0TIlSm2oEGrHKqEoBSaevX3ZG5WhWHqiYi/nwjthpWJLkfqBoOIOMZdFIvx9wMpB+7
9Lo36D6N6tbXss2p8uElkDVVmJvG4lIjv9qEFS/WSfEH5+Eg/VKqrrPP6B7GrSlReD2Tz/H2+lrX
kZk8L91lBIvHBCF2O70wAw5x//Kszt4QIXwKTqj9oD0ECpjmwv4J5QGqN5Fx1Ctzl8TuQ/NfV7cd
aKRuuCYNjs+/AbWGZK2Wc8ARlMW9ynmophe5XpKs9ivrMFeZpNtcBpr4BE+sq5GE7SRvKCh5xh+h
ko4OJz41hFS7xIAnicwl3ae63FRxfGcJdwQQsCiCJVZp4E9o72MDdMT/OPzjz/yvfZZZcOZO464g
bbtUoam9DiI5/oxNVE44P/ioCJaDSBRssgCfp9YCnN3ElIu3Ty+IlbtTtUSyRW4b6ISEQjzKMdPv
8PO8NrT5KY5UBl/oiV52Rx+FhSIg2CwXifCPq7lLSbM6x23NSal3FWOJWjEUYcJlXOjdAakl58iA
ami4N530zE1//BwH7yJjZQrlrIMmoELW4l9PNIkCaT1A6JOex7YpO1oyGyuN77duUAppkLZrWh2o
b9YS1DyWit78bXjN2NVi+z6ddsSceLQkAUMf18dnZEY5ldsYlbGrUayei/5RU2GOBROafdeWQQyR
VeLaDpL2yb5zEdTNRM0SbL+BbRSbU2e5bCLfdbCX5mVWFErH+Xri19mapkqFp6zPX7BYoJ2rhLr4
M4DGbo1KJywaBU8K9RP1UJo9C6rJzOBXCz/MrH4Ho/mjZH/4lQJFxbxGMf38IN7bJKCQo6Kmh2SJ
X6uCTYe0PDwWG0GaUwi3Td6bR40OHC380OTA2DxZZZJIHK4pOpIHyYjA+3EJRpnyEaXq7T5+0JxG
WkOsCoyepmrgqOZ8SOKeRtGZS2r9CvvD3QU0efD8i77vYQgmV22cY5Jg9MDTavSIH9de28DkCLaa
HMXnnWNtPX5SsJmgewMkFlvayMDnhGgBUcWEq19j2ISKWRl9jj3aw/4A2Ol3ovhi0SqQeHHF97Dw
ZFNGT2A/00eIzVBFa9BaI878tpCzkMLT8W58KlsP+vqVo6o0VvfYwlFXcwxm1PJKK2jk3QHXCCdO
ckH0BLJl9OkF8rsxFEm0XBTgLRg+qIQamV0l8ZEHF6zmAhnVJt+b6tmoFb2vEQ2dmYhAs3UnF13c
Ll7ZcFWqYs9PHZPQghFGJiNfIHlgmmtX9NZVKS7G8Qa4JrlFwC/H+6DIQVEfrlUnBeJtuMJ6VuYG
vyB5I3AFqps/jM8Z4yhTdSAsBNcapn+lKepuLCuijkNAGk5liUv4YCa8Hs3FevbALW4OLOF8xMaX
a2xtmeWyStcJI8amwsMOS0vTObi+iYZkacf/IeL5oJQcjtojeKkUVkeqvXj80kGI8rgtNDuH3pLq
3nC5mpHEQVkautgMS0Fbrb7bsdEXgw3PFVrBh2QZwjFu7x7tezpk2w234RIGWz8D7FNh8LpqmxZx
EJ+JHSA+WRx06y8E7dicD2OfijrmKD7PfoEFZEOXvpquQhJO7ocLUtMK0xAKobbZJcH0P/1xxWBI
qZnk8I1L5PKitopJmeWuw6Km1hXdgKMFiikEqXCDrtUd6KpE+7ax6HZA2nLTE7/Kerq/cFF64U4D
fMho0A/e7MgcdUIijRHasyG2mk/0pWsCznMt3TjQa7ruCP06myUMFbRYFO78VbzgRPCOWpc4xgKG
cT+hVXTyCODy5EjHvcaZQZV/JkkQxRDm2FXy3jcTRK2EgMnOcvFwqbyD5SATJFXjO/ETXEoplPnJ
8gIM5USmrqacFibc327z/0cmf+jbiqu8mAx0TeMW+eelukN7RAeSr1xBp5qzmZAIQOE5qtIftb2h
kJHb1fp2ezpn1om/OQUs6d8kekUkvpd3y5+8GL+ffjm1rxRRhHWLrIRJov5Ps5Xy8mWimxmPUi7O
IL8NFWWjBVynOtNPQD/uAEY35Hrai459ykIKDjVOwMuaMBxOuLOORLSFg6LU3ah7LY1PKl/8/uid
MbvzPiLpwQb8cAqbz461wPMVCpih0rPc9pY3QMDCyk9f57/9xZlUd9MMJjzo7MKxTOaQdifylSo7
X29y82hHv/6QoKkbQAQWd7rdcq5nM31yXJW3j3YosJmqZTnZSOXRVr/ZBknBabCzLpcA80Vmjy1N
rYbIZYEHcY4K1JzJJMymfnGrKknmouA6RvA6gDWHAmYOfABcSZVwkM0ECtu+m4FX8667AOe2En6U
MYsZM1hDlZeZliZ1CrRBG3jLH63ccDF7rwccKSSJkNVjIQ9DEIjGbsqcvdrZhmubJ31CEEqyymQp
epjhFlmQdwPKhdfTwAVMf6/+ZDA8i2fKzEgLkHwVdWHdiX3j4BnTyCYWeYKHoTUX/fBqldnA6V2X
ANRUHR/HQTpX3S2WSclws1CU8dxeua5bSDOaAXXk0qVLfLUr7ITU20u9K/8lC38/vk9nnjRkTObg
wNgeEdx1Dd/6INnyUqRR1BWhcnNu3N4A6mnCoX2DEGSrXvJ8bCeFAjBbkT5ZNMDorDFMDqbVnA26
j2QsrV1kqjg7s586VgSDIOnG3/YKMdFkV29kT2LNyB30Vul1WERCejg2+4VxfYADSStKkDFgSooG
4Z/C9GwFDphKWAN6IoE6+sF28HA/CNapuAihtgik0gT0XSq7wDT5nf1/u2xAfub1RWWAUxkNSqWY
kGtQ2f7g03m1i3v2KUdXBJpLcrZNDEb7j0iJo8nL+t2L+ky8rwD4AYX8SP3/XF0uspJjqiYH+Q4L
77xqP5p9VaqreQ07SCheTTxgpHfovutjThTNB0NEVewOZ9MTqluToxn361Ti/meOvViF0tRtA65N
8ZS5NayT0Tb+st2hcqmcmkaVWUTekAKP1W/ybdXTRiFaJcexXMsROJN4QxOUWcI6CVswKRSKM4i3
J8Ruoz3f8jhXGNVvf1Ubswki2OB+QotS7RbIH/Ifx8tgGPcOE1Zb9IszF1HZRHjXkPqN86B10oI7
hSvVPC0AInATNetPDq6Ysa2yJFjqZT/aOKJK3n/ttN2diFuH13ym7N1TH6PKYh0+y6kB+2cD6a1r
BOchx1niO6tKxBFcPPz7BYkqPEOCdBQTp60oiBIj5cMyvC40K8/KrgIRTwLOTqrW6js2wSq1Mc+/
VSMPud5c130I80YkO8tY/1c0l4ZeOf06fES3XiKSPmeVYNWJhaqDPPr9EGMSrLKZQMfRXipDTwoO
0uULyqa0JSHOPGHL8+O7pYNy27vEWlG2ooOYd/b4NFeWIiJq2lG0J6mDGQRlTa1yuCLvZDCfueZZ
hEj44jv2vT/tU1EtjvhKXAXDYasXP5tDfAz71HUzYq1VzjHE5oD6Nah5UI/HZS+tKq1tOX9H0CFN
zqamGZCQfOl4XV9w+9sfIoPB13nKCe4hC/HDBJUor5COzEXKT1w59VTZL5SrI5Z1IS127rvnclga
1WBMRWviLmnUrXETIX+QWPjREXlmOhK3vCZGzSAiXq/OKLaLA6leja2R5X0qrEMXjc22A/Pd1Cu4
+IA2+Bj0ZeT+q9hpV6wfCsz1e1gR5ilBhVSE3hQll1jsEyYp6Eom8tMm3QgOi0ceoz7fkNWpto4v
g95p
`protect end_protected

