

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
pabZO1I/O5UlEfYaQEPwd4l9eUai0bqYoMxFZDUmBPXyS95K3GW98Ld97MzJKAXXnSlf1PewGW2v
0RIeWd32HQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
MnYS98CLv6GUlLtXXj0MDq/aXJWBamrEeFXZFkhzX7OjMU68I3JzEc2/1UN3CHInfTII6cQBis+f
MSPPkhHYfjWA/UnlZNCfIbUjCA7v4zzzEDOXLdUwHhey61M2PDbtjo4F0M+PSYsHQUE61FCJYZr6
+aBOwyo0CpKkCUVEbxg=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
qncW/Cwz6DQ02ZtEcvyp5WdAA4sItotGPpP0REUtLyqefQhCtJmFILcg4T0iyRUg7VuYEwIANO5+
QvHNNc39qIJv9lOesalgHBZQgvNRJnIdYWaRfS0GyacwI/2JQRwAkuAQstvDCp4RTc3l8lwP6/ls
9Kgq/wnF0FIDD2zIsqBFYPVau5gOg+E2Yv8daLhsLbgUNkGI+w4/OZjRbQGSUjwZLuzAjcC7dEzW
IiD8iCe2E3P5aTpTA2tXeuvseQy8KOwVCxJQuur+f/bmnE2QrPi5PPQMRcOyc4ok7k5U/64SCKlJ
oITfL/xIL/xwZa26tMPcLgkkx7p0G3RLvL/tVw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Dnf6vaqe/V3pNaiPDsCpL4mEkUhuRTF8jsptuAsYR5QlsF0hNdnCfK2+aKM5H69faCvd5mpbM0GP
Pqz+qhNmOYPHdckgaTUGR5o/7QyV8YKLvzwfyDMqTu2isTv6FP6Q6welH2CNBnmC1/h5T7i+fy/Q
rlaoXYJxfrB3B6n9clU=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
IMf8iBP4Q72XIQn7cHjsTbT2wNsnwrpqWy35OTpGthg9IgmIl2PQf4/c9imtaZPdkPVpIBywT+vW
p0seCgJeCim8uHSlCA4Yuvzi7NiJqnEZtjEX9xSzaDj4EflUudOJTsvuYMqv/3kxvUgkIK0AS+U7
CWRV3RwJIjyzXaV3SkeD5i2xf0d/bezTocOrvt7wO8hz1n7ziicW5bgdFMZpO18+84bLDi0MzKYQ
Ad5OLz8QJgoCqRTe+B2lLXuByvKd2+XBYArz50J0pDfy4RubYe7FYpZdW50ze6dgBWVP0HOw0tLX
Pt7eQrmsKxnIhjnIQBRBht+Bb5QLkHSbaJnGbg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 8352)
`protect data_block
ndZwnJNqARJv5/JMaSK40t13vAhd09FOqanitILnIlw8zFrQhgE7hOSP2RjGord6KqE9+mUCDQId
sx1a4WEjKywor7pQq8+pPboBxSwUsrEzORFJmxAbzOscwmcYKh8bs4haLy3CfoIuVIp1ISVRnvkU
P8cmRROVxOj4OPzebaF2KdjJu0bpxqEEbZCxY0feULRqufJnVzZeSOko3Zcz7zTiVkdjPiHwNce5
lCbhZJYhpcYREAY/EJiPXMGvyX+jiWCouZ2A60gsuV2MMt74ODlhm2UPN3pycu458D/1UStV4qfm
0T9f3zOhw4gfg/5DbrpAfzmU7zzTpGbw33DnqTNxmko0+SHewcXtolBgCM+SaIIOJRBuHtSuJeMi
6nfqD2lrf6hwT26eCfJKOgqBGnbXyViWEfwinxXMbBmOwAfm88PezI+RUzXsaQn4DEcWDfu8rpVK
Yppv3Xi0MTsFzfS7XJgTaMGaOftJZ77p8D+oTLuv2DoMBeGp9B7wBqvZzo2TPL4SlKJmSoJmhOq0
01kMieZZIeVRdh1XCjcW33SGM9wW3sic2IYFYR3/L/jiQpIHvaKNBBvD6rkJ/AY6kuBPsDU/fKbL
3kGm8UUnbbK+QiLLHpQl/6jPpFeOVeMqABuZNKgC66mD+tl+LMx7sEfMQDPjgQLL/n9BxFzFUYlV
+ETt26voPXsTogT1GKU+JRDwLj+QleSsnv6VkcRDeV2M1D0jNoPGDB13UoMrr+plQFUlWiu7ZOlT
gB38/S7uf3ken9Fp0YgDhssaCBvueMAOIeVX2aq1jP5j9tgUWIyQlHckMVWqDj4qxOsxtManliF0
so+bzA+QnSbjbpSiORK/8Jvq4CbkPj+L+zpgSkaakAJnZ+nwxyJ6PP+s4wWQPHS4S3TsEqyfTlo5
s/oM3MI5ckOIbB3OVwIihRSbH4Oh/OHnR9lLzdc/SMd6im8wtaZSxFlZJSgIIRRWqLrri6LRGAvq
oJ/4kgjEtVTYcx2wZn8Xdu3k7O1zpa/sv08ArXg47yp6qyzy96ywilh4YhBpGxV1dWdHGcyNDONY
rJf+S/JYxT14Dr5vEuyABwSAkI0RRtnIw1WMfC/6hGH2eF3/fZj2FL1Rc1sPJP+Ea7eQMvea+Iax
I/ooe7HhC7Yuh9SVlIwZvjrrS0DvsJo2j6Hja1GPCIJugeujbTY0FiPIcXYeRHD8hizT502yqW4F
YqrO4/wBgT1Xmaul74YHPBO/PxDQUAyVnMaTBJ40tfEWMEP3abDGvuQtrGJEDyfPonlVAz37w4SK
zUuvvEbex7dRzlyZEsBtHwqK2jC4NbkRLgwbTbaiWgk57fZjkiC21o82Yf3xGI8TujU02rwMMgrA
/YkzipZQSWIrCQlvC3z6FE0f+p6cPyNPLMqlEvLaaheGTwJa5Bmk4O+aaD4+xQkr72N8i4i433q0
5sBxSs19jF/lwSERX324bWL2b/KmfSced6jyCxcogxoLbLcLVw1dehPavJmwTEFyZNgGwFoFv41C
w+ad8hw4cSqF81MNRP4VQU4sMd8V2IiMIhUKszZCTM1hAR0Kwm8gW0zp3Ginw/FSSGoSu1NlnPDc
P9VsZOZxIxKqWiD/pusTfb5/rNuJo1b0eXSLw7Fd8NOtaweFXmt8jBixbiZ5bIA2hSzRbpvJ37hr
+masu1DNaYl2To18hqoCrZsctQYGd7E5lDs2SEXgAEvt9t2ewE7yBLKv6sq6qxEovW+zlRfv2e8w
EoxyR6Snyd5qmYjeu9lG58H9SzONChIYMBtrLp2vMx8YHOpRyz1mJeE9Fd49pYHNKouxG25NgqZG
nDoPxv8CGRCVnd6wZwDWcbon97LkFQixwyZfcBSsiceudSa+YiAy/UCWo2kCjb/klmmRgoC4tRPg
ijjcxl+RCcZpQufCt4/5PaK++HAEte8SyEm9YaHkliSOp69x7NAb42PXlNsvubprvtH2ijBLYFPL
r47kaUiy2lRpvi9m1QTiNpjj2s0oYPK1ERdb4N3UCTYUCZs1b51RKWo+p1gbUIWdj39Lbm6d+DsQ
x95iO2LHvbAElLiKQ+NwaJBJgmAxsAEWShOf46RIPbvBLuBHEnPL5A1FM4rJwpW9Wp8+OPyjinaZ
m7gVnHFRWNkJO8b69g+BlYhCmHkixsYl7iweppnfPCrO0K8ZKls3x72BdmN9/mk4oChJeF/1SRH1
cN2YTXlmc0pI6yl3JDqS5xKcUwc5NMAqrYU8czM/dGh95XcNhyjGOiJmX3Nm/DtBqNjB5hndfoQf
xlLnLAMwUyGz6k/wfxnMtu8nU6l2ozr4UyODTCjx07Yn07KC/b9BFBVpaWDvEPYldFblRfARA7Rj
nfYdU8T64dW4Cqujr1zgC6F2wVRdGfturjIezvpG3cCuyDuUZIo5thUtfcmVcSRF3AY1C54XVUr2
WLp1UNvbZvDbZJAF/0RFMFP3qE3ClAgM1etEee08SK9Yta3cfnP5kHVTfnz0Wz4H6icXnCDz9Fgn
X6zh3NS1w7DDj/fUwQjq3LzmargzKSMp4BwmHONiREjhiBMNpbW2dnfZHnly6roWxdjtbmY6L5yl
qQ5k1DEN9ow/DGqOmK7CppllUlkptPVGSN04OWqfUgauwyJDXTe9PprCOgD48xvZrmdjm16OxGE3
SOXj8zYBTen0p2hovWZ1ewFxYhpjZk36OKrGinrDxmS/KCVKL1h0UsICmXL/tkzu4PTEl+mFxBBq
JWeDN6t3ll+W6tC5wBZoYCTtzhFpz4Ycz6t9PfNfzUbg8oA1oSm7hdHpgUVZ+aEnOLJLddJkE5lb
P3BVFe9+iATeN7UlL4DhywR2ZUHjLuRXYZvGHn0aPbAkf9LrgfhTg7ZDp3o4ytcN+zn1Q3eHXMEY
KZRjMpNQnSODIFi8ydT9Qo/rpxopb3VwH/IbjwI3RlJh9Dt9tDNDl1xWA3xmKy+8vyo4d5xEYdz/
AZK39VP9OuD8EM7NgZWuv+sfrbR5Wuv0SUqoCE5VieYOtPix4V8jRsSAT38HjvjIfEx8+fKzO3JV
92pFdCSajd7WgssyaTG7+M7B/9JW1oRMLk90HstdrCob63fQzVS3TlJi6m99SeTFdB8P251TZUft
11w1fYT7AU2h3FfRHhV0y6yuHCdiNM2Ux5pRqcy/4hcmK4fUORnZ9/pwYdSRdP+NDdeDwtvYZrvU
pyOxk942EbV2J5pAMc9UbyszyKXZ98g94mbdgY2ftwBDMzut1TUFt/JYaqPYScZoY5QlaXXtCU70
/Ot3vlaZRkjqHaMJ3PjoJCEdSc1/PJChg6l8IyUWEhahX17VQsSxQtfM4vqfECncvSLif77vXpkB
J5KVjDuM8MwI425z2j91jyWfrvmak1pCBN7pglMJsdGBIjQ4I/Mq5qKjmW/azlIxsrVe+/p9f7f3
VFtCBbd2zkdA7To+n+x/OkVgl9Mn4ouMug+9XT/ni5swKlsEhIf2OiWz2/rFWg6vlDXPfJduL9Td
tRvLVtNCCM9VcGDQhlEjaIzOe/l3UpZY9Lx/D6VVbqlFQDfAn7pMmS6iPaTT0gQo0FAAJXIqBe27
RLdW5ldKoHxEuZUihlT/+cMuwj+lffDDZf08ZPBq7zg2vWLaDBUltl9utU/tkYn4x3/Z6LtFAmSc
fLvp9VXQiS7taW4nhhIF3aK8POA1FyXXV4oxIVZKUwGwGohHoBQW3cpVPsS5tayS9bxAF1WLX4oq
9gS61X+EivGTYKfvyz4iZHxmesL8uXODUGjdRveVVe1HCAwQK93VQeSiogNMqbbYKyKkhIwELxY4
ZKG2tYkYieDFA+8+cAOAgJw3uPl1Y3ymUCfK4O4ll4CF+DGRQG/ZGI+d2Y3MH+JoqHwvYwCa/YPY
Zoo1WIu+4puqLk5PEhKcP+yYHJwwItdy+3ViCV0/+H5o0A+AzeTm1vH1By8sI8OsUJZTEwhHA+vW
/PVbj5umHi6mKdMymZcgCAK6SLBV+Y2/zRwQ4LV7uQCr9tAs5IeDwzQ8sANV8447lFUQaXfVrpg1
QNQaOPj1QYuIkrmkuHawGF4zq9zvNQ2dTe+g8gzLn/NaNPy/W8CqKYL4lVQUWvQs2njLYcyfLOat
SJ9rXQWDZD3bZdkPNnrvJWJdQqe0RLYIIehVdmqWJ34tXOmEmo9bckXdrF+JiEBlEz+60g9r9GWf
JWXbxnpqV21SNo5qAv9nXLQwMAyCy7nnAXtYe6ZtPSXXmStll+jCHEYkMW1LcvDVbP6iRLplgqoT
GVUXvnbAzQ8FsHg8/muAyibZdpW7yNJeywGwYxm3xpwXvn7sG1FAV2cHcBqD7+tT9x81vFfjQSJQ
qL8kcXiMv2k2pZHZEtvgmHnYd9VhQ4rdFOxu3SbjTXYf/BXLgCsHf9EuLnhVCvyE3eWuXOzPloW+
v3v3FiXToue0hWG41yuzl0gdKPpqId+3iUlYqbNStLyxItyNOoaaOCOlwux4MZtuQ1YwhPM0nD0g
b/UPCwP+Lf0YuWOTCKhZdo5dtWI91fjyb55BzPqIHd7QCWyMRRbj3Mi0lBZ1CaYbV6dVDpl2m/K7
YtTzxsqeQmxuWcFw8eRkE8mqMrBTqHHKJikjzF81oSn+bPi9ahK81rFzblYDra+28y3P1g059S0l
BzHO27+9G5cK46mKlISBCO7lISX9zDcgH8nu/ODu6907tWFxlpLdlHAfoPGspYUMmQ0PvXg8hw06
mYAjaz6QEtQx7VCDMjTSWWYYKoQ6pUyy/94HVhXgMFyddOiH01CgVQA+Y/vTwCxg37WLrrQuKsVp
wRd4cP8nQJLDAxd+O0/IGtZqv6aEom3Qx+atT577FNTxZmBP1X/PGqYCr9J9M7TCJBBdqPbAEtlZ
IAA/2qELpSPk81qo8Nwsw/z3t3wJJP4eEFhV/BWH+KaKINASnmPM5gzU3g/fyk24HqSc07vxSC2D
hVsPiXcUw42RHf6BSBgRYHR/rsE6i43hxlNnUrWVJK5/lIBkhdQZHO6KIJt8qbTKAa4uFbKWevy3
eeIToL7v//XyUnSO54RIByjeDEWadorYuZbNPwHzwMbjx9hVCGwkVPRk1f8ZHmEyvuCxsGakGwfY
MEjpgKI3LaxN5GDVPeM+l8o8sTc/TVhwHclKRo/A/p/nmUSOFui+3RSIq5sq5F+XYdBhqOv8+kRJ
mLbjLMENcACKCCncWYCwCtEsSMUIl3iR6Bt/iSEih4b2cSjIOO9C4XlLwjDyJHFRmA4EVJKHy7NM
Z2s6jPcGyz+Ua8mU0KOu2/3wCweUw7flPnPqToZqs1zMcp1vyXs3ZJYTpkLUeWv8McahzLSa72u0
BsBB39qPbhm4BsCCsvS7p7uYGOrU0uqy0QgVwmpdZPzM4B6Nd13zeiJeQQedxQ+5fgtJIQs3LDkB
yghqLhiBh+hm8U4hmg497BFawb3t65wOC4ocM0LjCiOQNHDFAO7/fsx5Mo/x9jXHx4RzgF9uM6oz
xF/DfprKJDqLzHeEap0hmqLmiPOPMiIpOzl9Ffxh/cDTD6twVdFviOkeGdNSJcrDbpIbP3uOdd/b
J5ceh4o7jct9Zi32EN+1LcygpOc3FxFHejAYuQW6xr0UOekFCdxYqqH9MFFHC00d0pK3AS6etk0y
YuoRWt/OqSFoEvg+bwWVj9u/smd6bXlC53hQD3dPOZQ9Q+gpkZ1I7v44xjdCtliHSq8i/P9h07D1
b5KQjoRlEInrkLBCvVrvMmBttfMXt0dI9UurvBuugI6EAhZFvhvB8QxoESimJn6wYhwwCzhnhRmp
OvpgKTBk1c3stcyF2NglohDwP0GcL3AHVVZpcsySYLn7D3C9kdgPm8fz8dmrau7k+7Tymqw2nLOe
NIzUXEtW2foFgju1cSKCAUDZKv4izS2ot3JFKB4d61w99Tew8VyU5tfYmTpIFW9KTbRG71+T7Jec
41oFLJ12Pex0qZtA1Kx8qgw/IlyBKdHRHBuWNX5JUn1nJGNhxLUwkRL0FSm9j0jMbClMZhaF/THG
FBYtcFxdT490foZ7mOlD8q4o2pV6Zm22SwKwA7qSNnGJfQB9Bhc6YzoGcnxdUvr6BA7IJeWM9Kqf
oD57fYg5SUR0D3fZBsTcybpqfK3LZDkum9qngGftEvoFCZ5Ts63FB046HmQzBUjC5W6EDtPxdpUC
ffi/Z8s17flDtHLMP+/cmh4dWAlclJuLJNZ4ZRmmd+2EMFGASpSNAy+uxTDUAWrFyVx75vg3puJY
a72dB8WvEHu2fzbCvuSvRQVY3eTAdvGoD5RvNxhRmjuZAHxsrD/Ib01hvOVnblNoE4XBUYyVUOw1
aAhoTt5u9bzase7d1mDB6xGopvcQy3xRQxF+2/4mtkAUAxTRNN4ZpO7XDO+mB9q0WFtdkWqEvmhG
sV5kBax6XTsKSyJc/yQpNAxD1ZELh5iy0i5NzNDNsfVgrrdcr1bRUZ2PSMuE1RNdpPlVFEWAl2bu
6ulPRgyscrd7mg2xHBchvSnka5gQqm4kOoTQYsjXJfAFWofdwntK3kxUImo+aMSQ3BQQu2HgeAG5
IGGzalvOoVxQMyOfLx++/iZu9Ma5CgrHrlkcmJKX3BSrBdlAaiaI0XWxDgAfvWQQqMmcuxzfOMUN
L3kYwUPWqulVF0T8APSGSiIumuEYw0a2BG1umnx39F7x4RM2d2fT2tPXnUEn+ElWMkuk9gtf8x+x
FfuOBlufqOny3FaDatRA+LAH512d772K0bW6yovg5ma4AdQSAWxkh9/wON0vX2hor+JE/ovCDuVg
tcZtgHg96GnQe3xf8m3nmMG0TF6vDvK8q19PnwV67BScDOCvrBFl6zH4tKGWY1dNsf7UgrYogtRy
uH2FVsnHdjjT7cPtZy7HqLJoMrrJ+PLkBrTx18bhM0MVV3UrNuoaBCNKoDuEZHxxOewMEF0NjxOe
7+AItiFu6r3O88T4GQw21v3GkFNM+jmP+pzEFhLzk986DYMeOJ9bo5aWJZ1CRAb/Gn5WnntIjJge
Saf6+z/zPe/nd9nqvgbwBMM9MKzOrjl8CbkIpYO95LlMhgDuyEe0+Wpz9XxsXHYFsYSDmpiS1Q9j
PYouw8yIXZtV3VAsz9dhoo0tXp11wOo8QIwrt8vDfBoGO7oEKD4T12AcVAkEsjm8RmHRwMjzRR9L
n3XZbVE1/YFnzkDv2i2JOeP9+C0b1++eR57NJaRz0g4IZd10PGgrs4pStgS33PGmdqFkmtkldcwj
GuxcXCK/aQOCFMyzsmz8c/THn1fvk3+FfwzbX313CDPzpIpxt+O+TMLHJQvpKqOPwi5sherPqgZc
gr0M5xADgjAWX1vGy52OuwadFOhhaI1qeuQEtxenRVIG6jGjo2w0LGKHc6XgzfJb8WKrbf1XKMol
wDoBCVTfWddxhag141euibGHo33rd/P9Q3CFTpL54sDsiTfhie0ISJ3zv5aiV5IYzppBcedsoZra
oE8sHvths2JyHDN2YxjHpTaT7roYmgGo4dzklhWH3UFTJDyfMz1bltEimnYZ2MKNTyh5EkCUHHUO
2tJeSsH3ooyjQk4iwGr2nLB4mXJEHnlmE1Tf6NDX4iLyazVo7z8rNxOqWEEpKVOIyvjxgeC3dsMH
kKcfkiY8XxKC78DbfWt12pn4TLy0LU8dTHZIZwOnH5VJVmuIfMb1x5Gt5aQShQ1GjcQ8w4/AmWs+
9LPfj/RkDsmuqaq6YQVOO/uam7uJWnW0qv7hfDodBIUFDPy7ghle2vAaNPjnsJmqth9bcrUE2PIk
RwLANjS36uiceU9s1t8VjDyTqU2XFymXw5Prck5EA1m/Nt1dogKk2McEdTAGLwj184M+DCaD5i7r
vNzS/93h5dJSyEA0mUfX4O3w8YoPpGaLp4H5zlNL5rN3BJJx14uCYRI3im+ocS5uH1rvsp39/egN
9SYEEWg2ZXbFytels00usAyeS9myHepTFB8p00ldKtEsA732aMZmslS+x8ShopBf8u5ywoGFN/M7
s9wvUh91TtxALmLosXatinyr+AmLIsc+Tx7d0AIIQW930RBLloGS5tYLXIqu4LcRByATOCQsVcck
PvzyGgxg0zAEJ9MtnLyROvPJIEF5+V47myoNhgr18f66lOgEv8VZm2Q/wSvHndWpDsCGD5cDwXg6
L4Ca+Qx0vsDwj8UCZj7A6EkXu80/TLUqZNnV4QndkRQ+kPQ4QvtWUH5gXT2u2VhD1zD5AYF/iBjP
kj0q/u4+sTVcUOcgsVoKjlMO5lfX/WmsxtJlm0v9JsoCs2NT2b+5vXnGFiBZE+0gve50ErRV1oID
A+gkGdOs7l6u1kwNcaf/Qe2gIYtjY5s3ylTvPvAxauMLOliaDpoVrK9co9qOBjyYqM+vrz3Zm5Xf
h1I7R7qYETjOwIDJdS6BTuTj+bQXuDJJhjhOUKOS+4++C2HkMAi2HhPo4TAf8Q8bJgFtHGbj79P9
fSvYDRDpYbBetLLoeF1MPA7BLBLxpPFFW7cj1uarZWN9uYdfDQ7cSJlz+kBF/eFXV2riUsglp/cy
rEUwY+PD63B3x4jKb55to7/OMImOuVfgm8xO2Z7OaTlAHD1Q/7DQg0VkoqOWKvshRcx6sipX+m9H
4o9NeMH75pwSWRYhBotn9E0rGphyXNpkDfZXZV1YRKjv3efLlDGRfrcJkbic6cFpEy7W4MZ261Uz
eHbU49we3ghfEHrmgx+L7JkuLicXfl2qyo87Eb5lZqcdJZYlVX2ulPPlANdleyCHh/4jH6GuaQ7M
s381qhEzV6oQKNaZcG0fjYi2HJGNivh0Hf99WvlgA2kWkicTnh03OiTVeU0Vg4A3o3uWYIWjNH7K
Hf3mJ+g14syhyJMl/ZzLb5zVjV6JCAxExJWh87nB1q4uKsPtiMJBNrqJJfroJjuOYYLlLo7fw8DR
SsmA32l+WJmgGPrtf4RuJnd8adMVPe2OrnQsB8G5aCSBR4ugbN889XK4wL/hJi2n0PAaupyvykxC
1pG9BHhJNx098TCywQmIwu6ySQ1bAbXWksKDFUIreazYiN4tylqEXNN+y+2Vggx+KDpKmoJzpR4A
mFusMCJQoXOigEjd1Hf280a/0N+xaIkrU2aAfGwmEOJZXBYrdGeRaITY8f2+ftY7jbggLFZ1OKw5
4rFCeun3eNV8jyUIObk2K/H/QvsH/s/jz5QNLd4MejtQiyZBNMlbC7uaPUUCegoZBZmWZjuDrr0v
dhbEZ8wYnTJa0XjCHEYjCCqKH4xeS4PvZ88C0ixh40oEY4qO4TdaL4CqllhanNEwVhqZQWWC9Vjc
gA9KMJEcYfvmAGqWROaLk1jayKijlSMDEemhBTj/Jv8Tz8hjKATJKC6Wi99wajV8CnMahgfnXTdx
SQlX/sGTt+yHHmV0KnJNbnReIcyARuRPsPEA6FVhs2eeFPV6G7Y4OJWGeWGYyz/pnVqY72tZuwfD
MFzKD/DDpXtSCFXarH/F66FEetLBDpq23wRn+mVnw0eiJhmic8cH3y8sNxdnYo8dBLoV7gwPCH+/
OFa+9sMFotchOnJocVgVHDszE/2MKg6Ek5d5aGw+MRFJT8ON1rchieSC5DKzPy4LDyIHpdVnz0Ha
VoMKlffukeu/2lgtj5fO/UJSxWnls4bx/UGz7JmVC+MJMpt+O6ewWBxfPkNvtsispZJZfVqKNazz
zqOxIMcVSJqSOMZNHavWKs2tqWaJPb2W0f1g013125IsIauGItyeBriYoPgImm8h7nBGOxYGLe9b
0o36FH3ZTTf5FV1ZPT1zwsNiL6rgkxTmvb8spAwzc+w38I4ORslGUeUOQGrNDYW/gnjCmDN+Wj4h
gwohDic5rBhe31CQTTgSfPKePQf41FFJp0tJE6rTh53YutefYmzG7hytj8OCPSNmzZ3nw0azzoKd
Wigo1KZSOMV0cCT0w5iYNuCyKfmoz9DzSgsJdHMzko6E1UBNRu7AR/NAeN13W6dKRY8NCo6yhz0g
A65/p/Pa57lWFmVvpmZ//TT7W7W3EoO/NLLK9hShP1r0oL5qamolM5c9aTriWNzFurRoJner797I
E+yJh0UdnIF1FcyCDFd7XoNK9ucmY8uhzLgi9pPsJxm0M8UToKT5V+0YEPuLmD27372LwFHbjfdF
5UX8+Biwbh8ACUQ55HLDLw0VJsrW70lznVTfdx722H6NWLWs8/MJvqCBNktXB38T2r7AcB5Nx27h
JBcMkvGz/WXDR9P6rspW/8aIn1Rq1f3Vv/RlpdYLm9Cm4aWX7iLdB/Ks2tlKHIVOBbAE+kG3wAEP
74c2CT3pE7ovP7+5wuqDDVmnuRJi56ZqrYKGt2PtBdC1F57Qfij1ElVRG1CEYiBmqSbeTydjgDr2
99KTRtfUI1JxlMeAPrCU4c1As1pUVGY+1x/M19pGDglKAc7vbI+jiJYaiDU5Y7MPnCoHPXTvQnrx
RIFBuadjnJbhmLvopetvwQs/3853Xx3BtvLqoVpppNmIXD7bVHB9TQ4yER4ff+FJFRvN6MXTUDFO
yzrvXuUN6+TgseCqtmyGo3fLyiOxNjKZTCLFCrFWyOk3tKMoEpaKspilWlEt7stmcYFdnqi2nuBX
jZp67ofPsHMN6Y9YzWhWxRZCjXns9B3Fm/B5eozxFdUcr/cNY55pGVr88s0CwouOD2MsSZycjiL5
NkuZ60RMLVdX+j/g89DfG3lNVm2dFAuqGF2vxNQHJAR3IdZnpQjgr2nBuIEQuWFfcbLgUq+qUIDx
iUbyVE0ogsVb4joQ3LvWq4uyRwB1JFmCuiMDFaHtKR66SpEy+556cH0Pa+lc0XGPoM9R3ZCjRmhB
PKEprHFeiS4sz3OoOTuFVBQrOiXNk0iuN59qVONl8ITzdCFZJL1nh3WHRAt4iPgDGD1wywJknsiR
akyIGLODK0EaO7snjhQ1+YKjUAELmGk/KLEh0ewvpDv1tFLyme+uBV6KqvsP5LxAfwB6DIPZqwRs
2eFTcpuAe05dFA+/Uiq1EQE0ozBL0/fPDQDv/Sq2aBVSwyv1/IYA1rq89lWMMiZ6vo2ZQPn1JRB1
i/7GrmSO944czj6eJyoPZf7Mte4R8Qe3CM3na3gscZS1VfM6GQnztVES6mRycGQTmXPtrEwY+gnp
EYoLAROO9XEktyy5C/sxQnWJaTUXRmGcsMOcaynS
`protect end_protected

