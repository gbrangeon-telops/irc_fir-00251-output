

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
OJrNPv25gxVf6MOkMLDXm9qPvzcLiFn6cGPtPoJyX0DRSMUs1CiCHluul8VfoMGYUnRu9NzC2pDa
fD3Q+Cro6g==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
OO53+YxV1fz+fdQXiBafTL0TfU0s578DnGOkBDgcp0ZiS8qBHyL1R2PISafYfK37QZ2xP9F0gTav
+sG2DKzZYRShUhSDZBSgMOYpY7yZxYTXlswORtjPSorUAG9VDaJFPSJUqemfgu4AY+n/BsniNBx4
zqFaZSDmDQebEViRgn0=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Qtwd1yFLlmEutFKAPe2eqNz2v7W0I1lWfaUYyRoJyXavTq0FDRoJFjh1vw8Id+dlXsCh4QCKBOe5
q6ztRPULauE2vnffEDrTLD6uStkKikAcWpHaB5kHv8W/IU3+JNz65HQM8j8hOwGUzUSaTQzI6Edd
Kua78SuOo2L/RNS2CApKLh4UlLjlkL69KZuDAj8Ds+wPTUwjY2h3tf4V0N6PH8lPAy9xJk9S3EgQ
ni8vjkjW6lK8he+zqjEtOf7IEGhelGexSOLg0dP3NDhMEcaxfcI7Zo8kOCl3C+GMy2w3TEyTZkQr
3WrfN9WllC++Z6rNtRNAqHVgNVA7hObPvyuA/w==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Y5YBoFz+YhLFw0DE8aie27jXEk9zfvZg7zgS29dcVa80RbYJrtSDIAboa1ixJiDhfiME1gY5XfYR
MSxbx3I2ZAkTI/5DwNAjKseDEksXdqu1CBQcg+U5NxNg5wWuw+vr6DqkJMxvZoI9BhjAErRu+2EZ
DgyTp7XS17TjzQ/Lk3I=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
amEW+kSm8JLnUlmLoRCPt0pU7eCAirRawwzTZA3XEOaldjEiNg3FqPsvTGL5ScrzO4MhYsVv9max
1PQJ/lU1FLIUBgG3vy1UPm9QWkUIWp2rve3mDkSCfvDRku+GIP+/ziqovgiDyF46b73fS7Mrb40P
ha2QhSaORrSFucLp3v+D7rdh8lKmMq3YY+qxM1KZEpdfbausR1NP2yVxQP/t1g0w2pAjiWQM7wT5
6xmmRvYxl+7EuZQkxaCLozCO1ELg5LiuQuDVfKRWPdTIjtVbbBvnn/eTARAw8sh6+JXXfmhauCWF
cGkCTU9noi1D4Z3I/hvgJ8IXztgyejVNBMRBwQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 7392)
`protect data_block
bW9jHO9N8Rw5Pdh8JrEfx42kP+wP653PKBD9Hnv0a85HaidxxC3VRsT4PODpsmpzfgnxdPXeuVaQ
Qn5PvFVjpV2m8g+axXWFIOAZikG5c2ObIhiDh3b3iIImLNRJZULsEHGvtm5MSl3PJ/41TU8jUlY+
N9xYTJmow/bzzqcEJ8pztOuSBtYS1rYwukS/4EGhLy6vt7vXqq+nDqAVG60ZIZkGEF+rJqvcX9Y5
m5iLqxNKelUy91fC4jpHiM+lAkcGem1yyDP9BU15PvrUZ0BxfF8ANR8WfGRtDECO3jeTCldpHzoX
sLJSdtD4GgdWVCXYSWoFc+Y8QcBqKHck+yHt8meq/lbcLtMIWSn8Av/uswA/Oz90vhZlbbd2RS1j
bjpEJ2jXprcgd4LmLTdrk79Ir125PLsAoCgiqffUx6Ia3bbjFCOe5N9lxa/05uKtpbkAMIF7w7kL
EV3dfO6UROp4XzI97GD5IGhN1xM59DVPAjVByOlnOE3FM8wnfWPDIcv414QhyrQKt/5GsXKbJtrg
/6Wez4I9vnM7c//pkWJs14lj1cqAk7h9qhrWPCOC2qkDtH/uqyiUFWwOwd0HCvrWvTZg02zsX4BL
+us4KJgrBKvar/4ZU9cQJqaStMSrusYk2bQvN1caS4VEEYNktdMyKhFU2XJePIGqh91KG2SoQ19z
JOo9mNDkTaICHSjQPKJB2SWJMx2dEM9ARpQFPNRYp7P1Y0B6xHaFlQYVdF6C+LiC6Zjx/h9VRynt
jEEa1/lUE5g30SrYeCDUMr510P1GJpwTOIIa0a61o52INmVhhhYmkAM6y2cWlnC4RnQ2yiXsPYdQ
Pem6rNdj9ajkE98PpGkYXiLOmb8o3qTfG4zqosCaJdbU91HSPb4TOHckSnHs5IQK7fcg7PfPXEUv
YeDSgXjEEZoJVvtGir8Z9Bv2ZITR0W+BhlbzDboIFqHzmHr49xQ19tHKDAYEt2pfYeAyJKH1ja4e
3w/0enldbtV1b7Usxs1YTFh2eH7Eoy3e4bcrE3IiHYKvYv8YZY+C69SXucdLz5cXekfhBJ9i5evn
a1qcEQFgzFZrmZEESrWmTyb/hncpM0Iwut62K2r58TDgeGrFlAYlSSVOBGh29OnSSXvbc3BhRLrT
qW9JlOjW+7p0vy8/Np4cOZ+ht/L2DoTE7RTIp1poSbYJEoC8ILyWzIMUzSyKa90ZVksrVasK16vu
uL9o/N6MrOg3D/OQDXdWzvqqDLsVpAR5eNi4LgIDtVen+bfw1cVFRbWU4xNoLHleyhTh5wflViW2
IKyQvKpDs4+8CbbCv9bjje8o2askfjvLWiSNyjeWOLcZEtNgeARMgRpSsBG1ISMec1a29YPGAqZ7
zl8vDdUFYZK6OXtj3GEJzrsTm40jp+FGtLxhZ7pS021wz/yLEuCpe1H9dV9an28LDxnZY/Ynd4H/
ip0APJbEZa5eXHNhQoU4Y3ZG4OD4bBKS17U/vV7C7nq4Vj9Qb24k6ywP82JGF2FqSowWNhdMQeAL
ctftLAKF3eij76GGT+bJe0pbNUcxoZvmZYjmCrrWeTbS+vfL+/icKtjNCUb+cOr0H/Bn5ySIVILy
dftFFoh8lgdBXhW/5wVxqofEmvI/uE2pt2w0WkSkWpXa4PrXyt+/KFtTV/o3tywQ4qmdnWCcBL0w
/9ESssYa64/iKzaGt8Fcg5wWCPAa6Kueuslz5QLLnM4q9fAo9HLvscOIfMUcM8UNzrgzYEaufdJ+
Pypjn9rcN31QzcsRFXAJ0mJnk96NneaSFU2NKG+lKF093cJtVNwKGi9kcEpqLUfSxT8o/GD48eL9
IE73nZCuYk5xpaF74aKO/KtKi8MCljEOG1MvvOpLzu/67cX4SUx2mEqsVc/QwseYN8ddbqkHFA+K
o1x74RysBR0nTkvo7IPmxNeEpbX9Czmphy/15cCSejfwoFs9iA0bi0VmrV28jsPNb2U1tmy6/PU1
uTFYqOx3L9jtchSLWlllzQ4gpGoGjcHnkjRGVfvIcDxHxwSQv7w7c+SrUTaMGzM09E+SRtKFAtl+
XrlSezPaEsXZr1XoYP9cvF5aOz3rDMMBnSv1yVWoDvpFR8NgUMEVb+DKJ2xuf6gUZIo2Fx4JAX4E
6sFD4vlVlw5MxgDqkMw8Io4UDDISUYZexqCVVp/iT3PYGeQv/kvfFYn+ap66lPkcekqGk4BT8QyH
LYTodIhEhCRY9PIKnHj4W9zfp2PEYbjYJ1oDc8bJLRDQW9mK2Jp0mTxxqAwy+2U+4lBiQZ2meBDy
LwAjfpcnNTOKEatZugkdUvlEVPc8+b+604CiQJncJQx4xjrB9DiLiQh8+XtaNiF121kvdcJQ96PN
FiiMinxYjxX7QtAJiJHV/qhPB4STl6diheAbwOlQMzh1kwuG7dtdCCJhVrdUD3GvWJth4r3s05Y+
w/apxXFfYMZ4cdN7ozea6+LTPh+G29YySzGPI1dDcGTgAOZoIWdDNwxwcV5nap+IAZpNTQRoy+hy
umuX5f5WieKHgV8t0IrS/1xpyCKHj9iQNDskf1IVbgDnq5pXbx5+JrXDsf/fJnZTNAYMogGGveda
vAVB82q8GdKGj/yIY5IFYeKj6ADO0S2r2wRGfK6k6hubHHqGtI4+oIGo+riIoNs9WXXzkk2txUXV
w/zmLjpot6ouqnnZBOzM4oU3TfuAJp1jg1SGG9TY60iO45hq9H8AoC5xcTXwxpYmh9I+7MN7wq+A
NeAIeBKbak6ii1JQvkqSzqj546VRfIi9wBZglwzC2ZDYn4M0CvFODEHihJe1LJ9ajwSblcvI1tMm
9LrwIvyZY1LQ8OoPHh5FXRzW4aKb4WJprI4UnERgidWJeyCxRY9sLp8KOT590HAhlVEDZATj3PCL
tSE2o+YVYxrSx/AFpWZoKtV+rrDiTN8NLOUCM9o1uTF7ZAP3ZTIEZ9fQoMB4X+TrjZXA2MGpejNL
UtaPVkyRBAXCE2FQLQh8z+S5uxjgZVSRP4XfQ0lsbNZciIBttTQdIsZBGZDGrWbfbwkAUUv+34uz
wBr6q1OqZYxggVYjzqe6FyBqUnlI0zF62+3Ix/GD8t9qPLfAik2QoJDJAKmZA6JR055fUukm2r/r
QW9v3ROOqrFHUm8UM5bIX8QBtHd2oZnxVABRyj5fIuK3bsWmOGc8QwULgU45mub7c+7rxh2A3nyx
bpVefy9wKHptSmvzAlATqcpeqfvmksNhl5ts59slS3PLyY30zGgVkoPgrxHJTdIZ8jjxzmlrkk5t
t8oFWsWsIhQ+5R/fDjP86sM8UEEww4iPXi/ZoJuJGQvP+S4GumFoZcnrt26Qk7r1u35BYIlH0PEu
d25cw4CZB9Lz4enIR+RcnO7yF/BuQhEpnlwg7lc53YB1uzR+PN9qwXLfWdHlsOdXg6mLVl4LKrsS
8YcCyAvIVYSOMz+Lr7+suE8aLu5Mn6FMF0OK9F1hdlC/HiWOaVAcQTEsbIM9lRt9qattD0qoYp5G
bdHS5ufJ7Lfso0sXRygKHXDT+xWJ1K3YJ/QynRHC0qycrEkL1FfBx1swSZUageIK5h98qIKdR22N
Wdg+nFe/EbwXkLuy8rOEzUvRb5XkQRXePVNy/AjlU1tVTpl7OLx9F1Yh1YnCoNf4LsjAJG2PWO+V
8XEnKS7mJhuPM98y2z+LjvZm9kGp4798dseneT8v02Q6NAkdyWSgejbBuw/zrzsz+cDWNiA7JYDv
IRQ50wMhdYGvE4NftVcqbMQSVdZaDjXGJLWlmpjd0eN7UkP9L6Jjh1pj7EZmIKQYPgStFpfz9A3d
z9fNnuF7LrzDnWbbw9Q3nIW7wghc7lG2y56TFJm5ayhuU2GPM6k9zvo39666mOGQAfl98lzs6Gnu
7XlFSmYiasSzlNfkDf7SkeY4VqZ+4NGuUgly5zXYBwPiyxbzrc9dIcxqi78jlfqKv3l2Q3snMXax
WibQc5eRhlFbFfcr6awc5oCTW4WBylxYb26e11k07g5lwh3tmDt9Vs5zJcIXbu0FWuNo+99NYRte
SNLr+U3KDoV9AcR1o0BtiJG1m/3ya5KmzDQ3MQl2gAe7eP7w4g2wZxU9eTG+rhiO+frXe1FF84Yo
YSvkkGllzWLdmrn2h+gJ8S0lCDgW1rU5fCucxQrmpOGi1jrsTZnae1UB7ld8UWsJIUTU6WVwG2o2
YbimQa7ZNmANdfCBREeJS61c7NaNEA+MEOXsgs7RUgGs+uLwL1sT4CnDOOpauu+ZU6bVF4vxcvT8
T5gyelPy0bNNbDumcpD9ZeQ+439G6TKBeEntcmCTqTz9Xc7nKimQ+Y5CHoVGsOFgSiT2DbIpdesn
IeaAqRPU+cNkUHixitSWhIdL7TWmsFaUEDnxgfZc1NmSOF8BxyxERsRwETV/jcpuC9uwHFUfB0yF
E/eI2ngzkDiqw0VQZIlMppsJ5bPIB4kS7+hdIj32sQHqDQP7OcNJo+AkhaVmR/iDKUAqYkOV7kMa
5DSB2/OQdF9IdUQdPcuVRhlNbHksa3E0Y4MlixZWrA43RJZSTK5yZQn/MDd8gbvZgf8pL+tDnCjU
9mYfEByiUgGSSDCes5jLVvMyUUzhvF8Gnyk/Xc9WW2qZLsl/Y22XZYICWBSiEcOLMVfvoPABCryD
0SDsU0jAMwjPSkEf0VJDfyV7CQB5PVlid3LTHCJu00agW+IOy/o31VcISABd2PUdcdl574I+e7pc
KsiSrXKP/SIwaiXBebrU8yU7rWfBRZzWnlexe5JlqbcZ3xF9tgLikuiAi0JrWPbgYwM7dHe1CLsX
cDMSW3FAK2M456U5as88pE42LGIf/Pja8AHHFvSH6OqsZDRwcLJB7jjatcDsG+FgHMpkyQw7Q6B3
ZHayaGsx//sS3tHlXGt/D867eYyyNXcg0Du5/5JINrPGEgWDDJBfHz+8TkE52aYqhokDN6NrSFLU
FnRU2Dll71A2+nvtQR/X8yx0zJk4IHk9tTjPMRTl4flbDiFeQYY9z2dMziUkIUOJPDPzab5N5WcQ
CbI62GG9XSAh1wLtS8sQfTFrazSBwi2kfQb9BaHfLoeshnf8pE7LE5tLujmS36kO72M68QDKNHkc
/SfdrvvH2RZK65NHW6BTMj3Xeigw5JjuucU4Kl+2DOlvOAjQnIsWyTQGdzFpxSReD51DYrquEe7A
zjGvLNTXf3YWjIbT3qeJ0btpw2vFgm5dZRczTLJl0XQR8DKBtCwSXn3poPeuOUsdR+lTr4KwXnwF
DEhDKBE0p4/vuDKDTDA2Uf+8SlYgqxIMh6teSEr7m1bfgsixi1OrexYGd07SdLbOgJ7xK69x9ts4
pivz7YSAJUEB91nLesCDoHjXC28nMZtbE6Tl6jhP9BqfJaFVCM4J/0drwwjFrkYwH6JyD5Qh/ZcN
NKBQpQRdxzdtUEzhhXdYRsnP1PK1+WMByT+FCZA31b9rXkVIKAzdcZEieMHFcor1u8SN5QAvkEOn
DhLcaIpMYJE2xPkDc2VzeFVWhHbuPHH1E+R8N18SQU5Oxp10Nck/tu9HAys+IM8YdeaCk38+xWr0
J3SiXByC7P+EZSncdsrd3zTjNnLhLXMkcTEat0ofym8bQgpKDYNlNHUFT+hX1hmZENGeW3ErHLLm
U9xf7JXe6cSG3Cw++4G820rvRcuM2mUa7lT3+r37MVB0qr2Mrge4OzBW1QAlDbSQBTM9X81lmXKE
2fuw0NJeEXKNmWr366ElKJXn88USGeSkTpQCPf3rxs2zc4Njsj9SMdZP4KU2dhvBDFzYZrh1OMRg
ViHvWzd1KJa3OXC0EIkv7ggZH06YHzEzKqzBgmtHLLJ1tuu4F6YQjmjL1TCvM3s6wmcde5f/Bzq7
WIsZuA1lZWzM1Tx5z/AHsD/yjMbQooYfPBNfpbR8L49iTnFDKD8Lqigfao6YMww6kyH97GpPeOA2
/Ies1F/rHyRMiGWRoU01kgvundpWcZyP240mRt+KDEe7qCSBHmQNTmofpOomTKmV2waG5EWmpjGq
Bt06TyiFHUWCWJ/NqRXQLfzdygbqYfy9tLKQjY9yB+EjPboVsoNDvqQn3FDiURWR8tUWY9RPFcYi
Ws+SxZ1jHmfJMrH4GCsGjgdV5drOShQL7fgipWrPwQ6DGUjnukRLy/nFtTsuBEmsoEQt5asPBVGl
XEAMQ1wK+JuWLHLLXud/9KAiGtEIztrFV/FRt5r+A1KihhHOnkc4VKHgLyEgt84dWIDayXXgk+wP
kt8RRKj4EqE/3obc5E5cCOERuSPbdXKgZamy2LUfLs5jNnFMN3UmT9tT+3NSJYvS95tmJM87qOIv
vNEfVB5XeXDYYwg/cUiNHzU2HYB1njt0flW7R9N2ABTUEdftRRJVfZe5yYQddfFE8y9WVL2r6Kg+
kOk5A3IoOhbkPStmZhj/1TS1ooLo3ZN1f37pAcaUtt8cCK6f2aJ2Qo4C/m0ndHCAnhCENUekSGE3
wjkhmraYkzq5yizOurBuU3UrCaeX8w4vDhC4tWUdIifTymjPBfu+v5fPPW7FoPT9Y7uOpbV7nyuj
wkeipJDe502fXsqIGDFeagIj5cdqF67bnLqEh4M+H0okgwrN64GPLGRtgrQHKua6yqMLGoAwdq2X
ZDE6AYi0oQvAiYwCftoE08Lwls1afSJK2lYrrMSx68Yva/U6TjfXQlAPPXYAMdoeppHRNzB5mkvF
Uhi0p3O/u1GPeKcvcSidbWnAqXd2rydz2EPHMlCIqT72whr6kFKy3balgcKJbp7kjm5ESSCjxG9+
aP9qQe+SnDg7ZhI01ymDL3Cm3HcKzvwmZDe3J3k3Grt/pcD5NuAZykLUdeXZEpyiZGTHlHVCH8Oo
XRaMaA5bjgjb8XxzNXIWmp5m/NY+J0PR0U/I30zJjnegv6flD0+cuC2XfCVb+CH4VthIlDYUmGX8
SNEEb4d4LgAdsk2lwMhUF+fNb0JfMIAiEQXZLFrLXXdYXD8g7oG5u2TcMHuWg9VLcePDpoCRnZj6
7BC25xVV7JCPYBYPUkrYYVj9xr6rVh4y/tvz3WiIYCqmmpuNyNyNdArpvDm10cZqFR46ezrsobAU
iTh8E5XVXD/waRioIirlY/Kr1jXQEkaW7mTXnPF1XcTmmpwmbCUG1Pyc6DG1Aelo7ieDvLUB6+wv
IPYsR6ohlmZ4ybzR8bXCNhm1n1kaIoZqXUGBQN9Uu1AGUEWVxjKTKxyUtbn1iuUeOP5cnY4+ZTfN
UpROnFgWtdfMkUVEiTrTgcmo9AFR/Ag8tLX5MGu6PoyxJNp31cG1FFy5KHgdiOqTHq+5YKNDov/0
HnXU56ePgTjx5IM/KN6sO6YFI0xs6vfAjw0mkC4u/fIhFlgS7t2BduwIEqBnR9w/+uMtpq6fbnv4
l+iW400p2B6FVKI67QQnU/4KGjm+C7rblIB0Ptnzgz9XLoPOFsSTFMCQq4X6XfNcxaDxjNluN+Xq
1hn/mylVfgcmIzK38gICIJQRNGquvGPx2pEXjp/QU1ZMwMQY3fjgDIjU8VZNQnUY5Z7Njbsyl1Q+
y+QZytdxw+W2ce4Cd/3OctI6s35xcf6Y3jy+z0mpxBV9wRgqFohmnkB528mM/P/fJkt4B6e/9k0C
u6hzMuH3Izqh3djE9xIHzY5XOqiGp+FNpm6Pp9o1mdk93RgXn/k6ejknfv2DUQUcoAQT5Rfpdusx
7UHAkwB8YeQ4Or/yatbbAKKNUJ/xKtWRxoPOIE/mJGmulZy26lmQ+8MBN8ioqgrWJ9AG94AbgFpZ
Z3vtTkNoxfjkk1btqfd9DxoCqKC64lefOZ3a73QXHZUs3ubUXmkdb2o8Syuf9L3725uG/TtvyVnN
EWumr311G487SUWV8+j6frOmF9dg0LV5nNDNBNLVENP+HwPGMR0mMotuWS8trBceHIXowUs+WOTr
eD2bsKwOvwSclB8uosjhWdlE5IOS8uamZtT2JFagGehlu/hV6oOlKFFAh7qyE77Yhx5M/IbSJeCO
holl5bVzFtJrJKbgA94EvXyxPnovxB2YcUm/oogisUKAhdZwWqiSFEnhlIxFf52Fex8oC35BmAYm
C7mLgpb3CBpqvHJuj9qu3IrRO1vhyoHkEBqlywWuAT/Wm7z4v8yIhbJJgS0aqht1nD0vtrrZsaj2
JWisCvk9nov4QDGcs/kltHEK2SreUYKxkw3fDao0CeTEQu/W8qa0EQKQAf4LcWyv3P/P5Cvb58iA
/owiI+uXbnER6Te01eL8UjpeYn7OK/08gykwiqPEh7VtdmiA9O2YfEUJbDhBzaRVN3K6bGSOieFK
uEFMRJkGMHeOny4pG8W/z1SlXtIlYvtrAxVWGNrOrIugynBfHTS41B9Fw6CI1ci4QOLOIGsiuT3b
1TqnGmi3GFRMn5DlzzMPvqp9W4evt6vC6mRxxl6J4bbJNilqifW/m5Gfv8uYXO9FSJfKjrys6QQG
coJmURZCeQTy1giLXZVSeFuzBiBwYA5gBSJApFbQU1KSi/xCbDonE3Cz5KWjRZfLoQMHa0RUSDGZ
ZfuoT6dMaofBGUz+PTRPgfQa+29asxoicD5MUcjyOcVqHCa/GtztnrD14KeHJy2ZWWKGD/PkQuGu
mURh+Ci6xCmXYFEX0CDM7Lum8q0lxKosGVMQT99bDqTDZI93uyNEiGd+3oTP9+UPfjizd4jmEvtX
4IMtmOnYR3PYg83J3f/IDl3xcZ7IX5NiG5/9vfRMoDzYxndCxJyS/7xKjy4mZH5ksjo8HRO+7+Jw
E50fPFqoGxlTf6owL3f57JS6zrWx6BCkB3CST7WwfE2NBMZhxGyIdmGIyle7KdSFdZrehgW2KeuX
q7rHxRpEbvWZ8TefMdUBmWUttzWZvghtNueXsTMpnPymYBLU6yt/3sblHvF+9JdUPdSlFzei+8lb
RutlWGV8nGzZ3gPKXOImxM0BS91NEAU8Pu00yZt9xVcQaEGmm3rUiLlO47hriuDFuCpvZxZ+ZlKD
g7zrPPTscEuxLdXm+4ePcFrJp6yzuLki5kXYsk6s5ADdV76uD9RvdNIiE333/CmYTC3Mz8pXG5QU
Q/rpKRTelhquwdowIsU/giBh3RiMB+AudETrUsXFpd4bCuUb/STSZ2bJr/Wie4C3Y+qjniDmIQhK
nHv2anLDLQE2p9t/E0xZPwsF0ddK4YN7dtSwGBnX9pSJo6YuHmCqPfiBBxoJt/D7/DQkoP95FHN3
ikCi8wNWv8I4RSnLXvioCBVVxYLbht34qbMTOKDQRHFjUVj0SqyjLth+Wz94fLEsEuIYN4NR2sv3
zdhcl5RLJRCcrMhTfnM4tqJqtx6Vx3pgEY2ErX5N+kmp+qSfm3K20YN3O2wCeExyqujaazrQPRPD
f38N/R9ZV3QUqIhWN2Pp636MuDM7BBKonbKjC/gLo89UT+RkanV1UZDoWz5Zt5XqSw7qp5ry1Qmq
YiSuE/K+B02g3zsURSp3gZD01KXSohGtur9mEOWNoOsVUX3T19bWy8UPF6KOqxJXSbfdSNgwJJmf
zWsizKjtF2v/m9PANWrqXn8q61jt3Qbt2OerKolqBBiiuZeIItAgSXWVTQVpAnNzKryoClAOn4qT
gbriAPo/CF2j2r/eke8zPy0hSBN3wXoGKNWUcUPlYPJhRcwf7xIFTI8LrWdQjEg6zlL7VaV6i62D
+PXaLB4UB8mfmM8YjdsvP2zk1r3od9oDFcAWoVGOevT1NzIMVGiWzKn8523ai5XDY+YhFjdn8IVV
QgOxAvALUKcwx8yCR1wJMjiRi0YY3PvjN/+jQqy5iJOiSCKvrIOYARgkSwnwY788hcmG76suvfQm
C4M0QqDIQ/hh9ceqCDwYKCKvMWjfE6peBbID4k9zcn8a3r7ffncF
`protect end_protected

