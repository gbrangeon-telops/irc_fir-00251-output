

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
ccZ+VLNSpHtEulGuEKVDJLwcsmbh6zDXYYsSS4iGpirAhbXM3BP50jl4c3979n2YR8HDHLXE3QbX
SjQosk5Agw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
b11dY0owYoWaWqrEwg1RlK8C89M14CAO8cS5xZSZiTQ60prhJpRDDBFmDC0asd3vpmdy6xip59nG
z+R5fGAzPFXPwL2mdZ9u5u2h5M7NuqWsd4/PSQwIb2Zc37lWRpOZZLKl9FzYzSgF2YNv5/jfYnLz
E/n1SJLECqBWTvKh2d4=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
NDjOIJz/ezAa2sanfwA4cBF4MUjfAWwRdI3fhKW6WomA0dTdlLUaUk3d7HHvjRwYAFZbgsshlvRP
BFUgnI13aIFlirt9v75NS6zbC9iHo4+u43o4DjI7erTR/V7n1KuL02bh7njjYqFW2TM9DCTV7yyk
HpE/bHTEqhTIUHhN3s21EIF7fvF256QO+AgjOS/tV7UeysPdiXp6gUoJ4fZfor+WTfQVkJeKE9LJ
0zpHP6pDYIRgknpLIxX5LP5O6x+a+epaip1DIHLGwD6CJeBzPxV1RVmuuHt0FXHAwR75O/YbsdQ3
OLvEz7nBONr7GpqlRI7TlZBuj6FdMW9zmU7ONA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
23D8eH9xZzeJ+Ojv/tdSxXVchNNJmk24MJAcRI99YbyO8+bv8JOBxvZhz4Qlt9qTY0ExdOGGGFmU
aQ35HO0+71woQEgUY5FOSxt7Z+X3DhAwHoCaoUzrhIzpo/Vibci8Aq5CktZeDbbFyKqw4AG3L+HI
gLdEde8Lyo1jpmEidTc=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
MgM0EI48WvFKRy0diETe4cjudrS6vIt7158toM9vdseTaMD0TZIog1UmAGNvdE72kJ9RDo475e8B
1F5FJia14jZNw9OSBZ6rrUB6Tjk4EmqoYQgrN7x0TfSl9ybfwnnJEUbiXZrL/obnsUVUxuBuPHw9
KwRIU7YdWp4ONQdRCD9vZVkexu3R144yonCk7ZQbQol5voGa98xXkFS5wJ9AioaVUGfDCcHlVgYv
dd/x2xkSx6aLm3qbkMFW3ZMl2N86VVdkP+mRZE7JGaPyJ93l/kjtm21dSkDxSaPAALmdawaPAmzL
9Uhkk9hs8yLNZbslAd/6iUfM8JK7nIIDO1E/WQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 20464)
`protect data_block
KD8ReD1O3COZVQF8225jQ3VNMWJF7xONCNvXaOd3DlPHVtX1GivhmbVB5c5bvTgD4OqPJ21AwtHV
FQkNQgPRRa6RlYiweTw/PRQjShyDJ2ZN6kf1dzRslzVL5GBVduXL69KtMGTmjV4B8i1lEX/6M5K0
dEsyHOP5qRf9kxDvCLtm2iXEV2U/wWgaOTbrVe1Ii1/sj23cJTjm06BkXq3O8oIs22/p/6bJARla
23khqX3PYi6XiG5H5p9CKgjKQ8irgGztVG7JjuKLwVcKBZXj1gaaoNvoqKIZq7DI1Ba6xh+z4FHN
NCcV5EDCK7Yk7lXFjkkLEebw+bcRnZngaf4/IlAE6MHKzR0IyrQ5iZLkfmguUhMVbPq9fynyHbKw
HvcczDcJM270AuxWzNaB6v6KxY6LYHb6QqT87HNRljt/OG3xV8u4ULyTXdOmEimfbfeRtifxNtJE
UIObWi1IEqexi6VqDnfujtrLFVjdo1Yz5vFg3HLS9uYwmzhlOd++GQtg5KwJQ//09v2OrEeXexzR
CiOllcZ/npkX9GuQR/Cijps+mqfplVqeBEt+LxzLoQVz5Ao09wSPzIjrrBQ4r8tJGx4pg4rCKCxz
IuxeLsWsXm9hjHPkUk0Yq/FYKo1vESqX2qKHov7HTr5DWojsgw25CRVKbgOrC59W+JKf5idyoxQ9
S8p03r0XkZ+tbvHXaLxcYIsX667U590WNUVLBTh8evhjf6MPM82QDuuTaB2rZI8I1rezZofXfR4A
iSsrvdeXNJioouRE5iHv6dDR0BL6Clb0bszBwY8PD8grWi3ARVTXPBidFocgBcT9pit3RLyGvTi7
uEXquE80QWx2H0wMgwRgbAr82MByiYecVBltWFWIF2+DkoTgZVjpih6if81iOOCqYWySOhxmm1qn
t+Xs1ysIa/zQ8UHNthfLYtaJEJ73CwWvX8ZAZiAXUX5N4bnNpkJZ1eZ04LGhoZ6uTllp1i6H55/X
jigKigm3L1uxdMMMpWrJdhPJSAw3T8/uVovvQFtdNjSXc5GeQOWlgYRcTuv5kcQ6QcLWySlgj8U7
wguI7B4HsSVeAqFj/2es/DsAN6BQEjJcar05KPzBBpZRFn2cSL469ZS04RrxFW7yNuj6bREEQMUf
4071EPK94YfZD+25OneQ72ZdnziqPPSvy6DEP/glMQGIz3wZz0Y8ljWtyg8RYkxiYg3ViX/+PSw1
liKjLaSZJUOG712gCBukOAc+w8OIo8ARboolOZHYIFYkUoiDLu2fv2Y+WkDo99q3hgbMfSuryVLi
50whjlkHmsg8wCpoL4aBtN9LOr1/ggVGppITvisOwyJX4vhexw7dRw29AG91GjJzjZhW9BsymbSM
oJMjvZsnqM+qwAWcow19+jxnz0KlK1vM9TVxMXlQECG1FFtRGYTt/bjNvf9LEiB2Z09NmBFMknex
C9RVsYOyXQIkVSsew8/xB0pjfINhOLS7CvgLe09FOQ3m20Kle+SATUWWhUEY1RZpiRub5jpntxkz
3ZJHEtDUv2jwYs9/TBSutPvYHUwBcUxPT7QE3yzCHU6Osfd5hEMBWiaWGyEil81mUBurtGe4f2FC
UA8SZGLgGRQ/zRXCMR6d55TeyDtZ6ppMPv2Q/l8y9psMK27CTKod03OY4/HAkHCzo0x7Wllds37A
y3ZxmRemYOXhfXWi7OFdD15gMvps2uE5Wbv6Lvm31XdpgYCEub9Ygs1S53S3ChFtk2gsVH9O4E13
8aPMnViMuIrLjC+GRaMs8vK1f+mqMrp8i4F9HUrdBOvdBK90E9BtTXVIVFQtFtD9uEhqimA2itCY
e5T/6fTP+l6Xv9+1svqfeSPnrCjMcCL5ehpOxIHk+nD4KEGsBi4ShWrVFOu2zDZ6gzw52cEFZLIY
5Cfgk3K4nCWjKtTX+rMj4sSth5bcMwontXtaakNIu43kdc+7ZCTFdSxE6++zWmsFBB6eIXYkuzTH
2EHBfWhS3uodMJHjcAmfkqKMsDpFx30ZBD9FrziTL+DQSzc3Enjxzb1pxAs7vbZjKanGlNlm+Y5+
HkJGPuasfocPZh1+7Mxn2azJ7XQ4FRrISn/UJ9MkNOxH+mOBjgJbG6gEXHHY0BTWQZNgmJtgZo+o
rFS5BCGVSqfLhDAOVE7ccKU5HyHelIgmVYf6sAo5AsjzpnhSgbj3Rwr4GRhzzvfST99k7A7lE6Pv
RHn4+cEwHJpRIPStyXxOQCNN+PoLxvWYVaifhqFLS6mdd7V14lPJHNLw1KLUwOU1P0YQGdTYDxZd
xPQO2fxXtLsTewv0PChzR1NBKJkdqtjVFXHHVvVh4N5z/gS+HF4mBlHPVMcqPN1xSM747NzxnRaV
GU1bqo30k8ziAegz00+W99qasGjrXPG2sTD44OnTEX6qPLtM/w3H0dtGHIB/fHC6wQXvJPqlDOyl
sXEC6OOygLQ/oNpPTcogxh6911j5mOSjOKUwkufbWb3Ud9Z/bv5+o5P6h7oiHuoLS4TByn49JooG
Q4ywRtWYLzAAVS+ST1dPJp2VmHFT17Rv8+uzAaJH4sFWKuLGYI6RPukwAO/D7ONoiXckW8rj+uya
AizZDIUEPdkSqNU74LBa+rDHDXty0eIlJyhVZ+xJSwKJWP88eeu6Df4rC6SRv8olr6h78NH/FZ2W
2yjyNqAsJmxVOriuiaklpB3tCtsLOzPphCiuW1cAAVzaZu69Vc5TWdiYHg16F9nnfXVbXq0OuzLU
CHsbXNyNKogZNLg4yOkLabNqeml0ii0dxI83q+FTxT1zmOKLMFLeisWOTYpTGuSY3ezyF9wSW+E3
fESxoTjzyhbJpG22htdIXIxBQ4STky61GMaSt59thyLTGdmU5+C1kdpe8bXS+FH+JDP6dG424XHU
elr0wsq9LieyEWXBCNDPhnkpWctnvnTyKG99thraP6tgLSTkAtVrVP8bijR5UM2BZApcSjaFWNR6
ZrUqHEUNUUhCWS87R4TCRwFc7/FoMhhIPDC35ng3V8IjXm560wgKS6Wc3LYrR11UIcbHcuivcehI
Bmq0banLRfk8uwzAsFWzkLZG1iLra+sJPS7WuLDSGUchI+pjVgCxN2FOmutg0/kSJfJHfr5q/lLc
HGmNayu4BlQiT8un1m+vYjgpwEZMj4c6ocffI8jzBseggvivMv75NhyggCJSg+V8zMFk/oG4N7LE
Ci4Dju5lvDZzcF7/k2pLxtH91T8bz3wp+0ikARkvIj6RCxB10VlSJ+3pKDUwP+RczyqKPzlmUS/G
2gEk2bGwcrQyYVBziU43QaXbfPh7rHpTUgT3ZhQAZwBkG1gDlqHrDWTyFPATwdDNCIoPx5Dp0Ef0
gwFkzItry9DQ5FaISleUkPT8oy06jTM1aWeLFg0VJvF+YMFqmE01+F3hb2gfQN2J5WXalaEYYVyH
0bZijok7Se78EB5qBL5f1kVSfnZn1hJ8lpgCc1y6YyEJgaSsRE8jUQN7khBi/kYYof4PNmXkUCGm
D+qi67nydzVlV4G4fIXoNlIqyI4+OKdDQ6PTPxdqaEVJnuJuKzHvL5PsvQL1Vs2KtFG1CZl6X0g7
GBANVCbxXsu0R8RoKTKSd6Hn2mcLNCyPtExvCP0YqvsdItBcyuqJYgrDMBXGRaMcTIZO2IlXPE5+
k+7vzefnnqJs89/AAOVmnJ6butYCCJqmZXusV9Aty3JXqZMMD0T427hmCxrSi6UPsjo9ElWuPW7a
HjT/ZEOCk3bI6wQ7Feqcshrdndyv5WVl9OpNcLWI22k6oGV/bjmGpiE0AgK3jtkxCLc+2VRPdWki
6YzLfWz7UBuLD4RbdJOOWv4ta5z/4N+Tqlo+rJEChmSZSdE04XRe+xC757cfLG7PxpMmBSnhQ0JX
aonofPLlOxquKhA+0lNxiY5OVSyp4Zd/ifjc04LsBDvjeQVlObgyGCfdWzYGXQXMaV6e+xYajksL
rvTwP3IJ4IrSgHBxfasuTN4a5Wy44v9A1GG+GTxo6Wv8FR2PxhkKMzUcHjegtpRH8cFUxq2Q5z4C
BPEaynDohO2oM2UML7H+7s+BX8NhM1a3ZJ9gjULQRvg9DpSbAYbgMYkwkZkPeXKUUwS0FURsg3AP
W15+dQtJB7DGo2x95MGBxBzgZdB7+vON5ukoRd2UL+zVzQs2B+XUKk67vT9jPVieFZGINFqgkAwZ
Bp1rZkEDgmlW0NXAaHfxp6kdiOZObTD9o18ykxU5NUUmAe8hgFeek23j0hzcv0xXM89SIHX58XVk
NvwwR+THCNNJYXSAp22RdQXkFNZfbeipHnPaHpmHE8CWXZ7/Zlo2Pjr2BRAsjrtukFX9GcibzD2E
ETlS5Ac8oZ0LTudlW0QCPHD3pGTi96EKYa39CU1zFHukNfjZeyf98tfhU3apeZW9AbTlehi/cJ9E
m62G5u+VwIicxjve6F0zx4x6e/T0aUvTA4OWgk8oD1yXzOX3aQlxiKf1eXgZB9YQckzTbq5C5gBI
3hsugZkWyytxEgMH7ZR8VSfa/d3uuEBNuvipWqJydfgJ9fycNEB53HqX7wtGYny72FNy25wTZMA9
FJvoKdCOjZE0iodeyMMvW8cvNYjYoGJ/DOR2t5Agf2sQKY+7xNZVveCc4jgczgx9FJCKj4yP28nm
mKzNL8ugkRezw2FJpLjSuz/nFMWvSO8/34694pPVNSkhDp7pFjKPvX3UQi9bXhLBTCozmG8Gmskg
lLITSr6sx0OgTdL3OtYMrGFQa26vDOkGegvkp8HlWKfpof+dgiz40/cTanK82rQZd4StukTE5kWs
I1HZzodiBPRuz0AzkiFCcSHtSgRu0XulVz6x7XO8rcvrUuvNJ4gUXymmdG/u/M+5azhXldO6Dw5D
Q2IcNrGjw8mAbB4zWdL3ruXyjqnyndIKbuvIfPEOzWkNMET/wIkJ+D8/2p6zqjVM899GnJGooJEP
t+2o58u4SUkJL0FMBcCKKyZR8kqNDvhdjknkOvQ/bMrpQbYwMiEh2tqhz1frh0G7aqr21XYcL2kn
+PmsZQRo+/VMTDF0sQwW/0W9/pLHnd+pGu7bd9rWh/07wCm7266uLgxbRh42Z9eRadTcxVLowLi/
E1Oe1PCqFhJEWIdk9uy3yfF2nSAtAKYl4I7IdQl+q1Pco9XmKwn+Yv26abiFozIEj4zYxErXRzHT
O8gQNm8cNOpQtGyCce9vqBNkIqRY0Q9aYw/nc8wd/eS/tVHyu3g2DVJXnibqDsbaKGnyF6u0JAQD
XYbXyc+MKZp/Pb0YTJe8FCD4TnFvnp/NwwXn/mqTco51svWyGCZJuOOBy7pc/3sicXux1X7EkN1g
6Bte2w4PDNUjSjTkEMu9Hk+DNsOyMF7Z+f6MIH3t8gIIO9n7rvf/ZwmcYJ4wBTkTa30xUj+CxcBV
oN0G6CX+CGufTh/d2K/tundqpn89UXdUIa1J+OQNJDkd8MnS6xSZ6g726+UMOZGJvWxxsPIpfVpi
8UQpvuJneK/2VEoYlTGAsaJHl+bT+td61U8KfVxq24iU41msdTdGBVf1EAU8eirFlC/phiArwBED
g0CZXWdHQKXr81FhWAaaPeu4CWntwhBD1zlxbTwWbq2VGrfw2i4qfhWXx8AZsO+7XmNM5cLXZoCN
UE/THP1l3mvNHV36vV17Fk88P65P8mjYjhdpNjMOn3YAUoGx++Cyo5ZNlzUgr/tXbFV3wbRa0L6C
hXJWJ5UWUkCGCE1+WG6+3G6cadbV0JUEq8r1m57iFbPYesSTc6iwyyijVjoKcqaCXf8tlctMV06h
peVKdA0fQMuhNhiIqi4/9lNYOofQPCN9Sijva4xlViaBR46dm7CtlInH8bSH55EoUGnh0xLlMjqS
d3wCHCGMPidGwRzybjV0A+/5lC9fIltSpFP/VQ4mFIcU6IIkAS8TRKPkfEWJsn7HlAWv2InICl9a
XN09NnCAaoBPO02vqpBlv9YzDBvu2HyosFfveSQmH+bpJFRiIjqUVxuGv/IH8aQMdH2b60tIIxyj
SajwGwCmQVUM8ijNWrQ1uoSPk7qS4wDx1WvrajnBwg1v99RmS5CZqLNX4lVZEZ5kSvxa1J+H83to
rpi5qxYmRXEZNaHOSsnr7BbS/r/YkRKEwVgBGqlvSFTlXVCmPBT30KCp+ICSKGxDTNkyYA3nHT2R
Csh0FkgrXaJ1H1h1zISexSqhDj0jgDszr0OhiIpMp0fTWXCl/8N0Q58DYSlpTF/w/Fa+pbi6jP34
c4HyIF4cilyKuF1lpQfI3yz8QvhsHHsvNMpe0fSFwZcMIk1CkfpMWUzsROsgJadZimr3Fl4YmPLm
5OR6nBCZHu1vp050CWRGWfcLWnCIdCRYVJ31Lam+uiYQBDzsg1At5lo0eylh6tKSvhXSHIs6gkjb
ZiIIoEk0o3hzNn8rvoPwVaj7XDNf4+v1mfVvkxQRgQWeilp8VG8ozX0yqsPhc9e40OUWNFSW/ls/
/dvp+PY7/Wop4q080J+Njs757I6IMTJHKKAtm7XjNvLcZAp5s9w6iH/UXAGq5vkNHfEiB2E76GOS
ehVD+CAwC4M1kis5owj3N7yKw11KhEJaT1t3Z26KH/OBBpBL8XG0RjJ9ocs06xGeM+sZ/F2xBTuf
7goV/khnNJ4+N369CqknPF278Vqm51LrG2O+ka+n/C6yEye+6rhH97ZTLyZYbuRpI1cnFzsHMdCD
SFss7/+Q7XLNO4SiWdm0CWYli19wl/7JOVYrB5ISxwGuilHKOnLn8ePFmYX7C4vCZNHKiCpxtaOQ
JNT1ooch5i8wasi4N/ELzNgsxbHeHlgIiAbOKjuq9JG5/tvrlVCHvxL/mUslRcOjuZSrESKMV2pg
z3ViSWlYBtA0NgCxF0GWb/k5XamkOI18B+LcygfNKLp6jYRN3X9oTUH2uvf1M4IKblktQWbRVILU
Xk4So6SqRFvnKselLBic1MXWslzYD23hK5wawG2oOcnt0I+NH9UMAeVBweC6R1iv+CvM28KEUf3H
gy2njNFZEF4R1cyiS6qCPQiCzzl/Y27F4Y0Yf/5tnET3n0rsUV9mG5p2dg54UM0+gAIYVlnxJ9/I
KBvLegUWF+Tcj90/esIbhucY3KqGMgPhq1rQoY5VYGwBgu6RRnFRhuRgOgyIEC5TnNM3YpCP5BU+
jZ/JPTmRURPODwGDMHI5TsqheApW1teq7hjXwn9+iMt7fPBfg6KV3DvbAHzhkO3D4AqZUL1OjlaJ
Pk+95MuPEwIRxGR/dWhJcIMLeq32y/G17BqIgckSqmUQwBXPrnGyQGq8k9QxRF23n8IVXwtB/lv0
5wwY+yfSYkwZ5DlJ+3sfwVs0w/5S4JYVax/Skso+Dg0pJym7oJq2ILN9DwWxEZEPov5gnUn3IWou
kDbjIu2uIeDpHhJPsFLGtaS72TSPRyPzXYatJGu0z368tcrvThav3EQf5IXSO7AMPhBt4iFf/xwZ
c4RaUGggM/msUx/fY9MuXnbORlT/CRsdK/mQSXAYhv08paQJlmtSnbcIYIYjQST1K06Wk/cinJF7
WtAnfXTI0NqZJN6WVtbiyepENJXt4MXL75RvT8jwnxewNLbWX/QyG4OCb599jAcIo4OwriW/Ieqj
t7/s4EbF3Q7jezyL3cC0pk+2cV7+XdnIQLxsR+dZSFqiNd8ys3RK20AUqKEsDcD1RbZsMYn17HlQ
+rHZZL3LDjIM6qq9vtiXOXD4U2IYQY7qKV6Jq3Zk4gfwy+N1qcq+T2HfR09UDOnXOKCwi8AVWZLX
uN8EyPc9wvi3CfE4VuUMzISeX8li/jMJElH4YSpJ6Hq/YLxiYCDUUyVwCaaME590Rjd1FsIo65zD
aMvE8NxFJJweXB/1VN/fIj3/w3p4E5CrY7g20aoyd1pkW9cLdnrRyYkYy+lU8LFghdKA7CwDVrxJ
jlBtTPMCqDdKIZ9naQGxa4An9frulVq5m+aCWFHxNnSy/mFiHWxYSslhC2kXBWYU1i4M0l4PvMED
QORriFrcZTTAKMGEds8/UaWVdV0eBZyd5VvagUMcBWue1PyKsquoFlYM9exJTIpASky+wobaYSgz
oWCMqbmMhDiad2dhi50+ZXlwPDkgXA5ss4q86AxOQ6za6L/wy/u//7anODpTSM77NWEH82YCxQlH
RneoniYq14JZrbpLTqdmNGlIoOJ/Gwbqfp6ND3ydpfUJozrzonRBUfiNB50NmSxB5p8WBPW6mRJy
2jFdknpxTPpmqeheSl5xEeSjBo7n6qaxe7YwLP5bwFDHHsAR9FJc1WFwuOKTXM4dJtjJktuZaEO6
q+Zrr27qBiCTpwQGNkndYZmGUn8aHd/5aKE7ucgm3v4+kBnrdlrobpYoqAsS13CoK2gkXbzClr4G
XY3XJbQykqO93T/pakmFXnTKS8CmCa8EMEq3UD298F1KegJSpmEYGkqiJWsLpgMZCTgtjhuVT4mG
KsVPa2hCbWRzASDez0+k1n3OeZfEPuptdwiKRzb1v2NU3R162AMDmcpwVzCAIRvxzFgMEwcKp/vU
cZ9syUDY0fJjdHcot/yrXXabglDBlQ6pBGwlPZd1fSxQmiaekWGJsWFQM6vc5ttKMrLnnA9RxPlf
1Uyj4yjNbE5VBJjnQ5nXu6q25CvcnjMgYXgD4fnOQ/Fwv8M9uz2nMjfq6E6EWiQIbi0cpUG7mtOA
l4LUSafbtbBXLLOqrc/RyNfzhcibUMAOSkIPdkM+euLJWit65nbehMTZlZhRrSPXzpp2DIsoPjVb
G5tmurokxFUL2+3wd0WOOLDB1+fIxlkL0Eqtp8/d/uAuCnY4xmfqXRujhzqfrEqq6JZgmawRNS32
a2KIDmk60s55baH4nRbZE3Uf5v3+VJnl+58PWn4tSgscXhWENOWdWvuTPjdLo3FjoxesUR33W8Le
JX8sB1BW3vWuEuA7hQb19wK4ymXZZz9Ts60D+qT/iaagtNJ0qtaavBKhZvaQjnirGYispQT+PU+q
BG0K/g3esgE9EUKL37KsPzm6wkgIPYkisuZt9AoP2fXwHc+Lzq4KKXQf2GkK9dZI9/PWk9qfHFC7
noAzwSG87NKeYGzopn6M2SwFIt0ocjsLASNPWR28J7FNTHNoxLA4f2nbKKh74Sk3Qm/jA4nXbe0B
oG1IPzO5jTa91ctBfFKDVg+NNXW+nf8Z+G0wuCj3rQyTDRY/u2kb4IcglbBgUPTIZhaaxqksYDiy
iyKgj4UDGXLdkHYLhDgiWCRgKvN4JmTwZjj8nD7kNJNFiCyC+RVhcGhWDfSVKLOIACXv74MWptWa
j6ytbYmhutIVvL7Fjs7wVeqKAdhG4thW2WL8CdlR0V7H7ss6A4WjYVdreXaNgsrymwkC/BSu5n8h
S5+N5JbMEiNexQLsvgYF1cU/MAXXOc6BCDb9SyZTBsJRuPnL1Lnv/RpM5JNArQa4OS+5HUS5k0Ff
+rN5Ew916y8SeR3hYcLqzGsI2D89+34ecmWEvGa941ihBbOyQ/66f+TXHmrkDhtuFb72DCi2viSr
2DJXv5nI/k8JefKvvCeypWLBzjSdz4/75PLezYSZcUSJwb5BwQUTrMhfxqxDVGZz9sNpznbXwUpu
oTI7LBOLOR4eGvsVExeESdHZACWFVOJtKfblLQlfWvqv4MukMu7NdxKuzB1LL7RHoB+WsDUu/UeG
69bxnvzafbs2uptuu+XF8v+isISsgsK+aeA6134IhjbI69U2TzTEJ5m3cFMk5n3A4K5PJd0Wes6N
ql+FYlpL7hphpJLyidpNfTczoSohfm3XhosZ0tB6MOvS2Xvg6t7SjE1hBz+G8up4oHTNgUOijqm9
AKSGj2LiLP/bI2hJ+8TqZpGbH37SMbjBGKij2GLYb/vd23YBqoL9s+8WFzXivGeHKfOy7/uxzqCT
LLXG3MzhDejgg3FLZkZBjxRWgNstfcc/8ZzvSIlKs0OjcBovBuDEz21W0Yy4B8LYyQ7oes9VKU3U
RA+XvFLAKVhq8oA9i1tvAFDWz73EX0ZnrlGOEvdzWVkwlH4IzI+WQXG4PDWxZM79GAsEEfFoT0y5
mX36JY3sWoxttLxmNHbDQJyAyyU+t1XK+rEWkHxw3LVR4HgSBg3oPi7gcy/xJ5z9VoS4tIYxawjM
OYTLDtr5rpPMX+AZK80jjUYTSlkbLWRCP+EZe3PUdpXk/uJTttDX9niaghg91tCREu0m9vqjxHwF
06BPGhyFHOdFo3oOYUGU+5FSbRWRFYk87qesiF9dSm6jNq6HUYfjuvKIBa2LlcaTxFt76m8cM56Y
Z3VQPt+AWqGcJ/6lW3qikP3ZHFPkbOWUcUrhoQ/AzQlptAOhQvL5BW/MLZvgyHkeg+IfRSUjtpUP
DonYJg9vVHGOwVZVdU0v9yg5pKWeiAh4Qkgpd1XvN9hnGxNRrV+/m1oe8t6+JXS8ccByZeLKK9aj
cVj+yGrAp3A0rOKyLfHB4app3TLEBSE/HAvjUPix6299afLSZo90kUwOBY+z1F2y6ukEcXGPj0wB
OiCAJGRHXJ6z947Q68vDOPD2IHpKo6syFMRIQZFfpQmtO+OpJVn5I7Ai7qgwKEQRU+TeLhpsWqT1
Pbd+RK9gDMYVPa1qGb5cZkiX0xRLyX7Uif8/J7gcWwUOW2kebzHzuabpARoQMhlDrmxyURAcsBDL
gDIUd3WBhI7KXzHCqZZ+GtrGt3jAyVcOHu6XUg6gz5m0E2Zj5Fqym16+yMImH8ZLuufImvaLKure
Nc8R3m9bEYYz4a8PaPg1CUY1+s1vEnBj9lNqGLisKK1PxJev+5YAk+i2Amo7eYhPrQauZzdqRPpV
8KA21xuPuClrIsfxH4lYmwreBqRGhj094jTGl1QOr+E1cty9d6s1bT7FB4Yyzsk7tkD1775hBix0
BFOt6zmKa3nKvYuR0teoEszqDPVCBYsB4/4YivNRJmSGf/Uh+prV+MkmyhGT/xeyqvmJZh3UqURD
gWbIRMGGaJhP/Cg3O6N1OmtBz+GsP1tBPzWE6lxGz/xgr2TM0WqbRwy72YiEx0CKY1xvg9P6DSGH
h4tCJ+Xel+4UGelD8+CAklOxK0mVtH0vtzPxFd8v7T1RMU39YBCYxq3mzrCb0vYKVqHaZEtSLlMz
AedJhqjnHFqTKMcm9qq9vAD4bzzLnIl+dtTa7Zf8IOgQoAVUKDD//zRygxdepiMmTzWp7myGwl3d
WfLkpEKeDjU56AwboW/gTcz2rGXNcv5W+22dWSSR6CqK0YNWmvtL6yNHRuWs7aeeKHlEefXT6llL
Hc481YV9o2cywiyibvAOJlQ/PKmxFezlR+3cOKQycDM1PudP7n6zcvwQz9NRskjS9FzfBY8Bn7qL
TAs44TRBYbJxgssBQbu07k8v10APwk8ovH/2qzs5JQXIp0rZ8Y3It8/R7kZ6XLxYNi61e38P0jWd
C1WtqRK/fU7jLWOOyHb3fXB0wja+rPRI/4fNlPxgmi/vId0fBcfl7R01mhX4DjEwaQEhrpxQjciY
2/Ian62RPQBIT14ePlaUQJbXDbDYsSliwmMWn69Qc6mMoVxArHHqU9/lJUFVveU2CqYNjFe5bsNf
uNQZ5Q5MwEM9upK95qcamzAHAzpReca8A1uGxsxklS9LyqjM4ZzBYdK6Rx8M7hPiHI5pvL7VWhO7
iOhTHbp3VtVRRvchT9MZQGMKSCJX9KhMNitl+A7WveGAPghK14vdFNsAr6XCixX5G3oLImkIQUY0
+NzS3wd1K+WRs/7+N/zh7wSE4aDS2TYtbIwmUEGNv33CQ0GLF/8JsMIjabzw0LWD+EcHL8mwTKBt
OR7SfHzLKfS/tl1lVpubEUJpTTq+JSLfS4XhOnZszIN/lSSZ2ob2JUZgPQsjPUjwG0R4ErJjs4bT
qGS7zThduoLjOlV/T+bv5QPH31DOWBveT2Wrhv6Crhg7JXmWEDsdWcwtXPmsGzrNWW40qQInFEzE
7kuN60Y6Dm06unE4NMghgw5nH9WKhlifC5vZCX2EfE9/Bh5Rkq222LigUdgQexBD94rxCI0aWms9
iOgOJOWnMrQ6I5fL93Dg3T3oMp3OH2sXhfrf7czluhijW3qBy/49SwQeI60dCYpxM1maathahgSV
so/F22AmIN7f6IEG5f9ZUGeNymcu0XU+sGtjyp70A1BlWqJAFrXruO/Prc1SHqJG+kPQ4mgH2VmH
9nR9/rNi4/zCU1b3DrTV7b4Z0RhYXV1ZPePdMsexzgluwbLcUCc2bQazXkiVNBaAQI8nvaE+2FHM
JorEbPwaFORIWRtTOt1+cPkGXAiOcFJL9KCrsAQn0YH/5AE/N2brBj5xZRXYbPXf8tdnXeU1pBff
bZMe1PrtqyjdWdeS73MptrPiKsee9dgscggkAjJdV2VwhKIQuRb65E00x0uGFfJUZMwnN4sWWabN
2ELqxJglE9QuruEq3TgkaFjJVRsAI9mM2/AGKjP3KXrIFsHaHd3u4aBdKPGNpWx/ey2Uv7f9H9OA
lppCBhxOGJJzfe3NrAXk1M4fN3DMwdVBt2Bgs+T+gmGA9YHoA87DC5vGoPgcqqf3RPpn0aQcBQt4
wfrZJEz+vMxIBhceJT0RMy23Z1FrC+xgwGDGmJzy5kPPnsVj9Vu6/fkRMEJecOJXxfnupGm5ivDs
7UpMgZ1d2+4HF3PCUVO6VT5SQV3NQZ+aA0+A6AMxtn/78/wzAK9IsGlLbaiUN4XkaEkxjPkSJWVc
0PtxElEfLqdrgy0hgLBVpPU/55GcMBe4jabAs4gUs3FB3ksrdmfppEsCBNpss5b1BXg/zd1xMyMz
WZuxsOtewZgrzSZ1/XOxW/H7EA4/N+E3Lk2vXjLEBzy7vk9Dl9OXxT7jDriwp7d+hS9nQvDckpTk
eEAKgOSgIUH70gXeUFvp//eo6wT2AgBQyDStyif1QHC8KVD0Kc7es8xzkaHok04J6mi9ZpYqn4tx
l2NjKaIJH5v5QheUw14gAiRJRIwsB76/zSBsPFvwQrB0/8igj38J2jzDH2n5vbEBJrqPrvpEegmX
PabTdBkAhKVFM/XMcLU/3HUjVW5z5gy7SlEjoMG294kj54FkfduWqPdYO2rKmM1JnRED4kDUm+rg
fakpEYMrh6y2EWvvPbBMoS7Towd/MvHd78gSylmCRBy20yYMcdlenmM7KD2LQggZ6FCyTDyfyh8G
ljeRXhRIrFuZRVUHy/BKZnB995QUB9IkCZCbrTtZa9V4jD5iFkNnBw3FXJMq0JeAEP+X/y9TSILn
sdFRpKH0I6c03f01aAbuuEC6X9yCtWUEAG+Cf7wMaRHJ7nhgWPWQtF0iGjvQG0VXpgv7n1IV4qtl
9QG5H76WU85oGdDaFb/nYs1AcZEvWXRmWGzNZfI9t/Z9F+EeLCf8F8h/u7xhCQotwPs6RylUliYR
+2LR0bW9KusSRm3r5rysOfu62uvM5Rd3V8/9/mNI4JkLmo24XphFTYuAor700TGvkGaOaHdCVAzb
XSqS9ulVkn5nGMtQX/SYtY3fTpbO/BuFWFEt+mAF+8LvZaiYhiSFOFO9L74wLNGXf1mjyp1Dn06W
EEoHt6ld/QkduPQRvDVJc+SjJAaioHtn/dk+8ZimnqB/VXOs4f4wJehq/gnzMPVTRZpe4GjrSWUX
LAozgGnHwcszpwKFVWwIKcEPKUlwgA7CESju70HEkuc6AJmrMxTCRBINoC5pRX2oGygiiZb7yV3l
V7IfqkBFnVIyyO6lMDxz6WWAyLndUaJppj05ibIznWiQ/ec+PmEaUMgnDZfInfr6Hhp4ntmlzs8X
PhkxzJKsyM2PlDXmbp2MepaeD2CWn6eFZS6GAWZe5KU9ZYfy+R2rkZTa39sflVFPuuzIRLQp6ovv
nIYZHDInejb4i4b5Fzz8+iqcherpP0g3y9GUIMuBlzi+VP1pJjHivXt9jbqPaf2GkEb6vb3fUzy4
7Lv0XdyFbD5ub3HaJn/msz2w1Nw4+Q6aYJTgVR5V29/BDlqVi8IK6Ua/CzYKQWRKEAUpydT+pNSJ
+Fwvfp6bEvx/lJByTw6rLMjyAdUo05nIczcr01mUP6SNVJn+xzwKAe8XR5s6YXTHA1g3eoG7MGkE
F9eMnhy7dozqJgdO1U3/6EwDDxD/wmJGwosM+i72ciGeCRkQhhTc6L1+E2QtCXmy3QM6E8FJ6cnH
QAlNaXKS5wd3XJT9Y8XrJQeO5XCnZ9qYbJPgOLWLTokOKZpS7g8WfQa/ycGLPYBKj997P+50lX2T
EZureoI7jrDlWxcWOruAI916nBzXcow4ny6EhoEadeHN9qZRg5Bcubnvkq0y8ZmHN5Kb8NITGu3U
zOfNtXCx2tHF4f8FMnh8pWCvbA1PeplXvCO/afbXOxr5wR7jeOtpegV99R3R3yqCGX/njo+cOYai
PMo1QJuOpHONapo+0tRnvZgXwexAbIdRnDKmp5VLDAxCFFT/+/zqh1xs1qLFZagBGf+djbvQ7W7Q
qAaouS4CGWePjgIcLKWB9m3/CQ7qFN/KZc0ca7S0ClJdx06GGU9ZOs/GuBaQEBLL0QqH2P4p/1mD
P/oUexRYPL4nnsORFIxXwrxVOCYExKQxCwxLYpHTia/LY3wnwhK0Adwu78xarptY7Tdx2O3W3+eC
JL+B/odTWaQB7tPVi/iB0zcW6zkLwt3lExyYXZhvT8iW7/FEcIyDQDK37tObDZAUe+/YedfYs4dZ
fsiW7FPY+EE7JVAcfwbdzzj7Je3ftKp+Tq4sY02zRp4y5oeVAySJhEgNXyEjZ4wNsTg4rz1/DePj
dXX65POwk+Jj6sxWZW+sZd33H+uIjxOvpDeMsmH+uIh3TuGqsPOyDdvRKHwo6no+i+nD04wrxo1Q
zugDLlBv1CLAFtD1vWNaoNbZeKylUqG5YHlQ5sUi+xUw6/N0hqJxtj5ErsACCPsardlt2n5rgeoJ
RImgx9gShV/2UeOhDrQDSNOzWa1wv0lGPDQnhM85jg/Cd74pDduJQ5jAUX5RZipBoirCuxlbEYIf
N/f526PUqvMxa0nU/CwXNR9aYcOq7VRkDGJ+/HM2zB5iZKU72QpA27v9cyvnM1AwFNtnWfItrX1P
ahdRj68Ii3mtRtnHhWlq8NJ05oWJ726rESdUlzCRNSUbFZTZDoFz/FsFG0A0oVKo/KRdsx2xUWb8
2dTjjoXGtqTkimK8y2HreGGdK/rbRWR1+1K1EntANJQdQV41y4WH/FOxdYUoZXbuzzZcRuxsRzNU
zsbIH7u6AAwPbchnv8+QlW9l1Yyaq5V0rPixvSy/z13ZltTXc3mN2vHVlQM4beCi4PwCVTEN5TzS
yooR8iKXlbK7RYhG4M/dJdOxBBif0Rdwd39LS28bKwfzI/orXiCohbpc9Fnnq6sx8qatzC57f0ro
COFT7IQbmVCYU+q0+94oKnZr4TBLKGn1gD5RzoahQFkA2T7qQHBziOH7EPNuVbDo0FmIibS/RYku
ZaIdCiOpQ/HQX8c8/nng4PjOD43tUlVZ2N2hEGkRLH+vnIg2bv5kdQEyXd5A/Jy1MghlJrARBUxG
lc5pNpidzVR5UWXnz7q0yK2XP3E1fpnHX3/9nX+3JXB5UpufPBERFhXNlr82Fcqs/CdLJuGr1ty9
CqbNJSSMpZhzlzxR2oj60WkP0BE0dtbXUvU8pHi05ipkOOHDI9/B98KuLkYpJ8ttYXI2ZIt5fVhj
mYEBqdynYlscXVoBwsWevprNVDW6OfkexD37V0yfl0JO/p8XxlTlpZ2GHa5Ic64QqkXov5tjw0OB
P3aJfU+ZBwtHa8nxJx2tAqgvJCpx4WOpQpfYiFDG9cFMtLLSNDBh8IN3gHDJNRE3Je/zCmIMyzOP
9XjyqqTEMie3x6Vu5kIbt3ZD4bNOitXiwzqnUEsMWOpTdJrSBhj2sYhxT7WLPFkDi2FcpJc4fREK
skU4UKtUmSNLEDMZxtjyqD8GZYDQZYNb8mGRHDGg1GsvBJig8hkDcKlA8dn/RtL+WIA7UEegcQn4
DkSNIaqUnATNIL9LlTqbhyF19ZplvXbnJgejLD41c98d9iY73fGcbs3EFq1SYSgCUKF3Io3nuwwM
q8g2AzpgapzfspJc5CH2vYhhofCkx5rr9QssrP8hQeUGjt78f1oAG7/7RbtxEM8xkXAfRpY9OWx2
zE49GhiuQif9vKT6wzZuRicBXYiWN827WaONLn5Drzooe3v9rbLc2mlUrQxmFSApnlG22P5JWZ0z
7fLnKUj3tlJ35zV9TTBYwzbshhUeEglk0qUkY6kvpLPrN83l+u8zopf7Jh+N/rLDClMpbZ2PLFBK
d/2OdLGl056k93KTqRR8fUveEnIeQjH+Ed5OnrHEtCVBRIO481R2iovOSf1Xz73YAONe1X4Bc6/G
zJJtc/WyrzAuV5Di13lMPiWkofjnvUDELqZ4z80ujnsTDom04jXUTeO48UYfRX8OQJsq5XlNkf8m
1fLCByx2w6rgsnBzKxgXzahEwfNIW2epLo2aqheHQPKkGiqjCLiFCUXL5Iioz0bZgL7tiw9C9a9e
JI+636O1AwP+jf6KtNXToPpjo28gzLa7LAdCn0J7m8k/axabyhpWtGTwm0OkqdO0mkT4nbniFWm7
vjrvoNEav+hrrAfH1umD1Miwj9jFjvyMP5ZHQ33O3iAJf2RGCWC3sQSwmN1VBPb7z3lDqnolm3Jw
G2XEiXjMqxYLCorrxQDQ4UNJmLEuIbI6z0FKkt5IHeJxqk88OSPyNfuNN77vRwQJTjaYDDARjvyX
TIVoLeT1rINN+/0fueUf16s9MN1GYGxRl1xtoIp4APjmzDRE6rUNjWWDKCvpSU9Uu8NSEe/L6PuZ
bj9B1FWhPuzRanCyKR8rWpIN/sqCZhJ7uN6Gi9w0u+beW2UCRLkVxJjpGJ6s6wX4CXPSxkj/I7ud
nJDjnJDkurbqoh8KiImwwBcfZWcY4vvhDG4EulHD0YSi6iVxabbqNUZfb26QswOXRwT52smc6hwE
JU2PdM6MWrFepwg2SMPJkEUVfv0VhX/RkrW4Zh6ih7MBrlsscURxCyMy6W/GcAoZk0ZYMP5VvsD3
FnNRnhQcU9UDPsxFaEuT+aMNtgtRvzV62Vf0VOb31e3PkLCWE06O0c+kvgI/SkmYUt8PQD1DkVGt
0rUY/W9ItEc1GVqwmNm+a1FKpYb3hgm4k0m0YzL5EXuMAnw/gr7FPYTJE//qE4ip1xBUor3eKOTM
YDkXOd3gSaHd4Nf9tJaIXYIAVmfPNRjYWnm4PlBUsechIKMyX9zQtB3oOAKaLH2MUhQQ4kTsyDC/
xPUbMQjXO1oW4cZLUNFOUzJrE1ZD9EHLg+2YF3tFM+8IEiPqIHejCfoNpG5Go+LqNumtnL2/0rtX
zeCVyoElSKTQk6S+AYBq49qG8COgN+/I1SLmOp4Wcv7oS9FP5fE0j+8Mbf0bPh+DwyIKJNn9FsVN
r/voRczGyL3ulO93GyxvAxBZil9Z5o5aSwkO3SxkaFM2Z6/8NE6iEpzfrrfPo1nDlMU8+WiD+z1W
xxS1x8CIVGqC4t51A5T6oTath7eloCsblJFPL768xbaHiqkaA0/oaxdIXzvnygRMY8eIKDlhZuMl
d3XcN6784Ww4lInNbr7MSzVExx1M4SAGw3P7gQYOzCj6Lw3XqgpAqKj2lMJ0RQyd8Q4QzqN+TEFj
tXH0cwcdrHqhFUeehcqYGNOC69+tLJmNVG3Gw3yN+ESSzRTW/7JIDC03xjza3DBeFVyYSL9+CsNH
OEE7nrKVWi4MlZ2LXCYctjGUxo46cFABjdtj1Ch39eXxga/aJsdrjdeFUytbf0Mv7av5jkgnUy1n
69qNT7LKyTKO1twXg39KCaVt93b+TD3ZX8/0Ga7SkIQQi/40vxrfDiiVy8hakT2T5vejH7dPpbBU
Giik3l/PMI6hwInOqTbyc0dAAH+t+/8H2bYyCKp5/tQe5W5QQunyqD63EeoZdEm+vDOTX5P6IEp4
DBuni4MMXU/1OlCNz6/2gxc6Re4c2WP78BuGarcKiQm3tbNVZjPw3iHhkyT3WhmdWu39e0dsIl9X
D0uXjbqsnVZbPsQcfe9giG+HaSP3b6scH3A83jPk7KIiNCF2MHyPyx48036Am+MiT9nvMjwdm9ms
AOC3HerMdrYgwfrJJemzEgJHlCcMaWqMmvhu6c48ZkOGuZp5vJoxAjdjuGW0v03728hdA6R77HLQ
X32VBWpTUEUkp12YLRUwO911TGiDHO+vBaB2xjTeXrR2Cbv4E5t8rN1xuOc/RrZl1QnN97Fxvpeb
5Pzmcq1FCPsNZn00zc9A7j3mNVQU8siZcKvAwldURBymYNHFpuo3bNJbA/NnO7Viz90h3QRvW9JM
CMkuJyoaB30tsAwj4ckCqErF08xjcR7rc1if5Adhzeub4D244s5pHK1qCAcZijS8wSXLfe5NBTon
KQUUrJfUle8D7B6hQUzY+/WzQ5bhRHPMdjVUzEodf5ke2yggsiKVazTJYZEabQw9bSzmtwp27h4b
d2X1mnocw7/tYtMWtzEI7LkZeP5yMwN8Q7NgH4NSBXZc3NsbNseOgtJMLHF6ZzhTX5Em2JpjkI7+
i+VADJvSZqeScoxf0BBOvGc8jgtRJlPlonyzd9iuIJHbfH+jHF0P0Fudx1kG3PjA9dYC6xUSfO/h
g4RfAvObLP6/ptlIaB+YYZU+uh0N6jHYxRp4Kri5ujIO31I/E8Bqcy05Xq4rVn/DC34Tw0Id1rnO
Fo3OXAY8sCSYHWrvCQacwXZfGceQL3t9psd6f9LC0+x42MwJxTnYxfqsakCrEaj+UdCYfaKZY/Sc
SBMqv18cygMGbsmkAedV4eEG4ikHpJEZIQeA4M+3VkvIR2ijSafUg/rN4MBnmAdrjMQ8LQBhl5il
d2ew7Mcabr12yYM9uA57gL8QSZhUhi2FbUF4neHK1f9RC8t2zoKnYocgMUGriT4aU7QbI9v2nJlB
cv3nuWh+BEeeUUfn5sqduXt3zxSfDSDsr++7tJH4l7TqKVu9lK6R71W+tj1NnD4Nm2bjBDuWqxW4
S5FQlVTvAjlhNjZpj7aOKg/nY55jP3EGN9i4ZBpgQJ0Pt3XoaMA5NGAoIsUhkbcLJViZQe3jQ0qy
+jPd7N01T2AnjN5vLpF7juNXhKtyHSqoDiREXN3XTrJ6iac6nd7adYFA+LGRPrYWk+WpH+RTw6Gx
AXzIqbfEgFCB42jl1/mdNQjZS+1Ps7jkEbdfBl+0Ghm2XZeKJIqPYZCnMfNqpC9gvk3WBqaHZmvs
Z/2nUwKaQak2ZwDGolQ6vweS4GjMg/a3Vv8Zkz+QKTcTUenzaNjiQxf2jyVU4yNd5/pTMxmPnS2n
IfjyG7PCE8ImiWk4TIXqTIBMd05DoAQ5wRI6plWBk4Vm1hvIS3Mhtloed5tM5Yd8Nbu/iZMGKz0C
z9gKVd2QhGJAPZRqHupR6k5tsbfJ7TC/RGgS9dazxFW3gZAawyvGqiML+9y0ggJOH0HNuCqXekg0
LrV08st6OGb5Vt02j/ngG6NllHLDk1AUFlqQLdElLjlJFDyQsn5+zslRlfW5A39TWxI5GLF5U7eu
3pZJPgv4c0SubPi3IFOTtKc45D71tGnoKKUVLj9LXq8WvI7ipLUgkgzBOQcki2QPJPe0apHACYzQ
IR+xRdGW00jYFU/2Ka2tOWZONwlGXl07aSAwo/AWtP85+FxkWNzqie1hMr9mtbZ2enBWI7epORN+
lTI5BqwOY34FfMnpqFYgVmAvZ/C/i/+XAc8+fmIx31bvkHpARA9zI8V2r8/PkPwV0sA10Rg+Ehq7
0XZcil71UOk7J8dvIYaKLwk3ua/lcVdFSKGu4FaJIOhicZg1tvaBPZSi4LyYitswSyQGwis/hGzC
cJ1QSVr6akrUuB5f4J1jS/XaGyzMK4bEh1CceS/mcikINC6bz4E36P3cE+YY7Imlcn2TuF03mloU
Wls5UFVOZx2IlYJL+DSVTHAF+v9wV0yfsOFusSy5/lYAht7GmQLhmfs6IkGjiUwfQHvDSUc6u+4b
WzINQQHA8h9r32ehfzz0rDTBxmNMCDAhQflFJXrZGzXpzbwzhPS0oHNRvjxhMNWXlYfETETfsxW5
fR4gUazb9PPtNbOnL1Q14E4mfl2AZHFs5JL04GnKmPm6oleGa+vzZaDe+tKPHqrEoeRyStb0T9+5
krjn7AxFyXlCJrMWQC8XjwR3ulqhmFXtlb2Ui/tJZ9gOPGLz0UP2BJ8HyNGsHfGdLxzylZ3NWOaM
D3r4WatbdPf9oeVek/s8QNpStFl3OPjgEwOO0m+2mb0OlgcUl3qZjWw61eU95lVruzjTqFczylHE
sNEouE7HfcWds4+S6u6C0uxPIFqO4aY43NzwViih1jRqmDO8JYLrWiwNEDFWuzPWUc3bXzv+69+n
JMHo9dyIU2Yc3FzbVq2bGCfsdZLc4aKLeCs2zWi5V7Ynj+Vcaw+gd17fhSNza47jbSYzqDmzUq+K
7IOydKrPOzxNCzAopmPap7LQWCFrwpK8h7o6eEH095guxk6RZMhgb9Y8IZyGVtnp7UuvkKuloWfb
fZfsQm+QbuiKBN0yzDdrssStknOaKnomukKWsUzn9XrSxZ3+wD5gw1NniC4A7icT2MRL94PPZ2Lx
m7tzZRsOAArOHXx/crD7AUwbqpX+u/b0Dw6mJYgKePaf3kf7LNWHMl8knuNhfon1/aYuQV3Cb5r0
XB/McmqDYRy+3iq9OSNIgB86y6DTTXKMBAAvpIwZLTbaJzukfFdJ7gReoh8tmB0QX9ggeHLYExcc
plX+tyBJopDDstTp9jPlvTLcz5wntm7/j+me5Dskj05uN/NyvEm++u8XO2gSB5j3nTnw0NSMlXiE
N1NPlpI7Wby3NIpf1I1DakzopQQCGBH9inroJOx/Vwh6F0aFVj6Vs5tSsbRz+yrYycYmELVeTCCX
NmPdP83wjQqllAu1nX8wNwadDrKIH3RJ8vfnwc8g542Fmr4iLMwwQ3IGhyPUYv8cfKy4dlJSFP6C
R+2v8BKMvc83KGhKPtAF8Sj+ev1REaqsbqgSo9nwhfVkPchgDZ0G8APl70IIldI1rWtoj82iwIXR
gVM/qxpTUi2hpnjPV90XldEw2f+RUdz+QIDyodsc8QuyZBKR9zDfXl+6BiCpVLxXHZ46hspyo0Uv
v4XoziV+lY5g90bW9ogUU26gFVvFM5hUOtrsY5cZj5FPNXzvdPNlSSpNibMX2ubzb3NiA5FE6Vsd
xynQoybUOjRtZjSiU5a3znqhpgCK0DeD/t3UmLLgBvD4WTpknVm9FUadOA3kuzHOLvtMN43whmVl
HTF1CiHzjVxNd7hOnfybjZP4nBVyjicc7jgrRcYwmhunFNWxkQzqkG1Hj2aMXSdWwFhncMLHXViA
ncS9Yi389H8qAUVoTXWZXjzgicFJyDHVrNTtmWutzK83+FsekmEIZ+LsA/FYfA95W8W8laVXlGG2
hudtsR9wAkIOA8A063VtAyDH4u5jBv+Ofdt/ZwXNCfvO8HyccnrIjEJ3sBpBZFkISFM6filDv2DB
u695EUEwIo/1INcuD2KTszhkOWs4QHnoEV5805NqU40jNVgSco55/Nk8krL8+2q9RP9xHsaH87jR
Zdrf4mKL5pxfpGIPC0cOxQVzQuYn9itJ35H3/Rc17yCevf01YfOIgWsibv1xgJOVjvgwMSflptwK
JaVAH543mUCNsz3DaqytlLaugJK7j1DTCkusZxiKhT8D8jI82f3zjFjL9hWtVVSwH5FV1t2aF9Wa
BuOY9Iz9G4Lqt90DlIDT9j2ZloofcDJ/6NhMn25BCXlI5ERgpmFTekpcoPqQKaGHi2XQRWih3gCC
KftZ9KDe8MwvAHtwLT4hizP0/NW97CnTXtL4F4pZczjyZYr7zI44J5+XGLDaNErXb5X9UA2EfpqN
6ZS3EGwBMRykyDxSz/Fw22x5yMwlWFA/85esvbTjx+50NJFCJL+1U1vtlEl984HaqitllxekiBgb
NnEBsQrg6huvWgxLY/8bc8rjWGltLMvyYZ//9zkgYQ7vYNYijOOSGSWQzw97b/PfhqH2xhERwuDW
rPLd7hq4jvj2Vlc+Ci4+D23pKpDJ5FrZZbadwvkigYHBKTPkGtTrQrZ2ht00suWgmbq86iS+x3F9
knQD9j3iVaqny/NXJ2lJq2VBVw46BscUnmlhgg89mErLWhRs3638ZrqXRBSir+Uw+WNz8luA1iGc
7pRh2e07b+YyjKGt0uB47zHB2bQxh3I7Oir75jD4fm/+U3aJt+lD0/VmqADwbb33dC3mpsREWuVS
I4rL5jRSyh/riiLhOuGuUK5keRGoyPCc/7UC3g3VzQZdr6HtXGLr8QQWXRw+dGMh2gIhaycSMZ5a
3S5GT7WIzfnRAusn3OE0qbOxTH2Y3VmfkAdDtMLhCXuXOJogRR60+IvF1G1TbwERRTwolhI+CndR
USzz+91DIWvtv8It0z91jREs5GJ+LOcKf2rXdQkgc5ab9cSg5yjZzpS/YHdJw0qGOG5FuVj+3sHR
E7v4OYOZE9UOBMsOYxUlZit5Z9FoyGEBnGQmflL6IGL9Z16hS3mDAnIR6MwMDJsmDnATI2C7fKfU
L+BtNkYcllrsa4Qinsy5blDLq0sBW2SUYrIkng8w/Bzwk0K9zDg3IMsVjWqhBafiCRzT0hMEJlXr
uzRLGATaNO5yEBQYItFWOGf9kyhXlyRorBYN+92yO6zUtZpXNNe/aBicbClYU/u3AYwBymrL6ltc
bRp3GjA7Q2jqrZxcWcmd16OvjE2peFIeSL1URYw5LBHt1EgVLGhIj6NYT8aAK4pa7eM/z1B4dFgS
Zt9VR4H+Fj9raSqIN5NmNu3Y/w0iiJDAZ4vjPZrANG2LCJWJfBq3W9/4IlWpkLAZ0/8zv3KB8nk7
s1V/tWlrRxynhr/YxLA618Lto5dUp2EMCUbNIne9Sa0tiabdV/05BVF63mSTK9BHflKa3GCTIXVg
VflDvNUqhtL70PN03C/cmpBQDNwO+TPe41oxjZ/MT5fuYodUKV3Dj50ALu2xtp0EoRcR0cFC/gVR
4msXiZOuO2hetogHdXe+KMDfjP3vKF6qQ0Z+ZhfQq+C/rDKbDws1q7B6vyv5/Vf+o9b3RVOy16MJ
xmHJiUZIiyfvrggYT2MGBB/3R55IV+Im3f/ojdq59OuSGIaoTqPXuMRNV5FBOTW0q036ivApy5UR
ThYb25wthB5pAEBIknbTPYBb/6DXT9Vuhv/8+vdMOezAyVZMCjCBgczHHb6Q/NKDLYvuSvHKiQef
KAxez6fXd6zamnGS5DUhZSWdRFpeSeZIu+Zh1vLnykPPAhPPCfABX9M6eXd7lFoiA5uB7Tj93qD4
1MMy669mv4q66rmmNS/J++qm2AuBewvkcVpuFN2wQF5hMS96PDQOtkAxW2YAyPreqCZBw/BQg1fa
41Ul36WePWATfmB06sq+AvjDawMCbTT10ABrxu9FQ37kMFe/JOx/VXp7bV1lD814G44XgovfRMIb
FRphWWUFX9UC0R7IhssCGBDcZdpZ2vbF95KI2aez8yRO/PZZqfz9yfS4jxl+E3k6V4BhG3OgP8Xg
oTIduSsKfCIoPT5fUCmTfFlUp8hhm/B4LqfHdxz4+7KTGRwP7nL3aAiyTlnfgawflu5hVWhC86NK
IiaeKQg+vrtk8vl432Xz5DAJm5MY5sijsbQC+v6dhdiNXhRltKFm6XFGQpoBGDN26xpFNpqMPRb5
MtMNFLml2JOgmlW/1LzTQngo0ryvsyJw9H+DZdFGSCIdOO3/YZOh8HZ2f7P7Tou+Uct9A0RVBuLV
k3YJFPbr8oOLaQc+PTw7dnGxEWcXBJspXlzd/ysYpd18bhrc6tnr1Z/yzT9UpqQ2NOexlA3eAzG5
jz9kDaEzEcC4/8F6VkfuQoy22dR5ESa+tq2Sqje82ubDNd65d/VfZY+iSyTxN3QDrLtdOBCp/6nF
Q0JFLJJNn9V6Cg+l8Sdmur2ndh5EQm2qzWu/yjPe+PtM4Pk7Dl6JlNBfFluhAckU/pvWIGkmWsVU
hKRpw72bfnpt3rOHTtWQnzgh6CW+P6WrVegmLXs4GLv04YSysjWRgTtMpN4tjjPSRLQoZzBJQ/Ag
W9Yx/uMhXxJvWsV63oqlv7+GmlCt4evHcCHAdt5P3qkIU+82irU17cJsrHtJJcQyecnUYar0qu7X
J3ADcnieledwicr3XDRgGqQ/phPZBYqXlI544vSwlIMpcpLzsZxq2WcMfGoZe0EWmpbdKJJ06zji
VCtLRdRLrhbaTPiMLBU7251iQHcq9Wi3EZDa8OQG/y2l1AQiLAJVSdiGOoKak7NlosbSQTmLjv8a
tr9a6An/VfoNIgGtpPRdFZw/2s4ZCi1/+Ag7TgPl/MZ+Ih0wvqvm4muh8v1VOlqJGzK3IMO/Y0W8
4l7DhQv5LuKA4ozZlahO3KWPbJma5n5s7Gp0rq1jdn/zHNxytx7k3AhAOiOlMgwcAwsjR6eTH03w
OEcdOwiOyJNCBTrWdOwR+lw3M/4acECSWcEOiBD8msbp/BPsgtVbrsqKzSE2XEXNmVsYq5IxCYmi
C+ifWyl8TOSQ/yiT9VD53KMS7nPr+8mqe7/RYx/JGLotWw7wSoiCcpLedAFVIyPxr6IDyaLbtEzh
4jifa07O1Sfyw81rKOdBMs5+FepTG/GroaIYGq2lkUK9gnlhap+3cnpv3kHW3xsamldSYNvEZ92D
+K6kRkiKaTUO6uDUxw1PF9fpAwPaKTQc0UVVyjvJ4dwZsBOlDvGef2yc7t0ejfFNPyKdaFSBF33Y
B6HUrc7BznUvTSfC0FGpyCvjxQFeNpaJT/t0S1O7gmYT/U3hdQifgi/JmncEw3x8cL2k/JreXHHM
i+PvrCjTpnNO9RVF+GEWUr7TaIPkk2uSyF3RV9LnTJjLFekjPZ0C0S/jIJjT/BQqMsa1KVsQV3Au
he93/Ge29pI7VRKV4MHd3dAFPPcwTReF3LyJz++SajLznxcJgowFVH+Gqa5UmMCE1xTpG/W1Mq63
V1qb5QMTDVxMAsrwh8D0SEa1xwHXaU+qsDdcXznG0G+3GD6bq0OhdLHxUA/DhvJtIY6CbWG1VOnI
DPf2UJwsp9NSOpAzfhb+o8u7Eh2NjWBWjx9wtCyMyKbNtDLf2uH83ithUT9zsMrOp7NOE5tXrQrc
NtVt/u+ICLmoO4FrErVdOuRx5mffmdrwSPmmUupVBG4XRoXF3gxb8yoYho+8Qrxt6+iRvRGkzjjs
yKdvifuqU6c/nANpqJwb/77OpjnrrZBRTgHOv/1x/OCzwhajH3eEHEmYcIAK8cjI0IIdifmC6DLi
JnDbwceX+EK778w0GJLRDj0wW+HVeSJWxu2kumk3vOFCicAuu++j/x9mUfUaeAFVaqynOrNIugkC
FNWguVew0G+y6jkoyspvDyH5evAAZodq7AFVHfHnHvm0S1vmqbzFCaVP2atTcvl8IEEOnhZvHEUc
DWJD89lgah1OTXNw2wtpSnT+DlJwtbFHYO6PFBn1w5i1vZXY6LYtB9tWTRHsiBbY7DuSyE8yIMdB
FafnSZtlgy+yx3SDdJP5CFINCnrDcWXrmYmOPK2Up+YSySScmicp5ia+qiwZvYYgCfqVz3nmnaI3
KiDGBLKNGLSpRP+CPmpZVzLZd5qnc5AZWmGdSXwgzqjXf9P8A5oVZYZdJed6TBt2vpwWARMrkrjZ
120omj97KesVlgNKU4GMHIHX2ChqciFG4kcLml/K9W82oeJOk+kktcsBxmtJgMtSeM3g+43DF3Wa
3ZZeVF+55dVB90zeSZOzlcLb+Kuo/zcY2W80uD05KXk2fP+itvo73l3p2rz9g75OQd8f5usDAn4b
ZkFEFioeV8Ra2nrHf9AWxWCG5Zwiab9A8/8xVpmvQmUGjCot23W2U9SviPX4f5/FmOG+VYdsWyI3
8Unvd21vZ+bzpbYTlHxGQDVIuu13s8l/MeTmht/q15qPF4vf5CPDxIvzlB4q7fgPK5qrUoW1teal
nBRfIOPg6UCABk2QwSmYvh7xkr9Lo/kCwklSx6kvZreGbWT5q2f7FER52ytIgDkiLmOwL4Ax08un
jcTYX5Fa9jNkY89RoPmTg5K9HnozhgbqICmNKSstWup6LDFuXE+4g6DvctQKCOlzb1d/i/K15kOp
1izPSu7GIRIZwe0PjHyxSn8QiiWZEb2ZsIB2oVe9Ff7gQwQ+y/olIcmvuPjexFbL8vwQlyi8vYcE
h6h5nBI2AtAL5Ib4bLoffsGvGjTO65+17gDYSUWDrgBCT2ec3wQgFbqaucKeQ6RuHQ4SyQRrhekg
mPY7FO5gf/JSCSbxMZSJ3xrKQUhCOXe5yh9eWVad4VxQY+xUNKIegZObOsbgOaFtbGJhDVYjJOnG
g3f7b3dKesA+ilfmQlsaB/DFBKMD6LeZpN51UEc/E7GwWZJD5XXor9k2z/7t+LwhTAq1nV1JBiAQ
iKlCbhZp81v9bMse+1NACJYaCPHHSuWcf05SmMS+8bf2oKuvIPv5z2B0kyiMkhXeyxTO4Mz5LL9E
l8SkfWZ9utpVfVmdLcl/YSC19zHmKo6lHvf2PFsRNmiddWRcm35dknTOGwn7EOxhA40STnh1oK/z
RxhZ6hSAxTflQjP4SZ8Z/V1OcYK4R+fa2dEToCGabV/WNTwQi9LftQ5N5vTKNawTZqraqYcvZYSc
ZAjx8d4rKchdrgt9TKkPg5lsznB68+XyWhgmHa3zkIrELjsIiaXqw9P9bLwF6Q5LBMqYa7TOf0Bm
++s+O9G1lEYIqvYpVDM3qb/Sah1gnn2/tsa3cvZFKvyCz4oJGeKSBLPWYwjp8MdDEAKX0EUicIXU
Cm1vv980lbSCJbPnF0FwLoL2ltSaurGnXoV9Zo4Pq4iozyVOrIGV6XHIdC2smWgwM+FqaIZdgeoB
pSQuLTQjnV5QTCSORcsSN7Y4ChBTGiv9bpWPXAr1AVXysV6r8v1TdH8ad9xKD4PHC6Ub9xlQ7eDJ
oHj4rSbNvGfDRPmAkxq41+N1K/vV2PUMaBIyb3bpQ1aHYZueIjbwahK0ExeBmGXK//UHQZjd9KxF
zXBjo37kvG1rmon0M+wYBadcQRgPi6tt4V/MXJ5opdfFYjt/SuaIs3gowVZFJGZ4RIl0Pw6jncnS
oWG22JE2O4M6660BQZKBQ4JLhMMEpbP5rgLQdWdjpsCu5B1FMp6yzeN725WnDZEaC1l0hHTpnA7N
wMXls+eBRZdt5pW3Fy5lW7KolqZ6rx/b50OCmcMPxwxXt93wNRcOLL5tghsgiXCK6EtfL4aMluLj
RQ==
`protect end_protected

