

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
PFFltKdLY0A82yxFqahMaWdN+zxj5kThYAcsDyz3A2vhpKKQpGJvV8/AkpYYPyltKlIzJB6Md9uF
AN2ca05J0g==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
obdm7XtHPDQGZMrK3kNZKnRt8ypfk4aZ9VtSDpnSwNdbgwrFg4uylDkc4YjBW8BFR32vEdXmCKFe
3L1bSMhXRkPXZ88hMJlBty0IcmSYNatn3RV9VG9yYtXM73zMkJ4NIx7KoDtvOCnGQpHNAJTknAv6
BNEUXajqHzh/vB/QNBQ=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
nx2eU410BtrBCSzpvDl9pNpIplyp0nHGgzB9LvwnXgdhN5HNF/YNjnH8WXRfWZhIT380E9zFeNz1
cIYhUxogcuyFP2sgar0PDv645GG14wyLd7prd/d1E3Ur29iNukQkz59OjXTEIN/U9Gy3hPt+oLVA
TwpP0P8RgeQqCkJY93IlvPGfZ/yeDQHrxDZUMFMxHHI51HM/LG6Y5RjcVEJMkX5GTsC4gSd5fEHc
DWDREOSmqmG5Gmciy22xZEiB1SI044vcLqlJadcUhINRbAw0576LfZrf0pjCGq0s1+nEKeJm9MeA
baA5VHd6hhXLwLD9jRkKDvFp76mdZ8cpvFpcXw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
my8iGpxybuJuMik3+8MRqWVv3aAmCE4oY3Ij0YIUQTpme5jJv8e5DOlNoLmgXWhUlepBCUyZ1Ysj
JGlFKQ8MBs9R5aa1TLi8cCVfI579Nm4AO6VpackDfb6c5/BXCbiBb8XeC9Q6z0hKyH6xYDDC0Z7w
m1jdROr8ONcmGBJr57g=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
pEGUMbCVqav8XqUNf0y2o1L56804gb2pssAnfqbrEzVo5CXZ9MmyISfyPG7HY7huXkJ9tWIeWtYt
bUG1XTbOUAj3uDqhigkZ4KnTE/68izmD5rgLlGDQ1sI7w5GLUgtjCBINeZsiQZ8IbdNK2b2sCu2x
1k1tcyPPvRv3myvuFaOhmiYYyCNc8F9T3cW6mq34yHrMb8GcN1rGLFkL16mdIcoRSSN9znhYYcLe
21llq9uuuR5MD7mOGEYx4bKUQGVdPOHLC411Ms5bCd0IbhTC0qWispRkmO0D1uXT6TguY5Z6gKTw
vMvXdJYpwStmSqzikX3kYI1zljpfWHQ7HMzzTQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 66352)
`protect data_block
8YMARd8XZmvbGzMcd/FjHnf8A4CaLNiRzNqlAopMHBKXbdJ77faUYptjb6cP7uFfFZ0d7NpQMWPn
ye4O931zsw9k5iRLvVoJ9l4UPLfYnLzLVQpsKAV0OyHBh5fao+E91tABvKEqrJFUQk/YFmqcu4R9
ZFpGtbpaeSV2BQGBy60oRS2YQbXVEpwXhma4qLQxD3bQMLwHsQJQ6x2NFgA24NtJuHoCe8O/1C7Z
oOPfjFuTz/f3fIDHgwVA3bvjYWsHfwKVLyzxiz4HU5AHoRZg4pIS6aNLOKAAeWAyVwy0f7cQrbJt
QO9Ok0ReLWjxn5lUDbSGIl+Eeuno7dXzJoU5pBftqgE4yyn1jWAbp3fdoE5X0GNMWeL8Frf3O0Sm
dtAcKNsF8W1uTZP5JXvj5kwNIeA8eUmCt14oVU9E4j44Zo3ryMURvklyxHKKFkzHftc4RNuUIAPJ
hgDwy34Lj/ASAWaH9eo+JDv/LhyeRQhsbrxbsVj+2cDvcT9OqHAOcIHNPhciV9XYEkL5D9RcE8Ei
63vf1E3ttM54CpMFKCqK9OrUlgzOv1jyZ0Jb75yhxDNS8g1rpI5PKtu/6NpnZ2ppMcBCd7mGtGiz
4bPG4suCJoa2qUBwe8EbKjI0LQ1KVqSL8yfAA3V9GIHzxJ+baUVJcRvL0wOHzeQhDKhRQFJWx3Q+
644iojgIQYx9BC2kZCOcevS7geNM8hyKLyOoFSHhXV+aHPzeVydtsIBtxk5fesWh4nvL9zppB6Kh
Q7WK46r86MhYWtMRSdiKxMKBBVlxXdYKzRTsBVw13KyF0bcqawYEhZFB3GF882ZkOIf3hO6PmAOT
pgEEhuooFsRMuOR75OZOQaQLUf66A+i/Ux8uSxZQZNMahn18V/Y+91uFFKXqUwmTHycYg4P7BcHA
XDxuOHG1xUdM61iA4K6VS+xI9mqOddT+/VUNznKbD/XAfLN9eJNOMnWfv9rMimOyms2UNjmF+PIP
lYSihz34lSbcIvYDpUCP9JymjYUVX5w0Zo5U48LBZ8FUGHZhGb6DtdvTx5SW5wlCKOGbTWPyNCVO
ykVfyDmZeKEbSD7QjL9kDOYyFV6HD3ZgjeyuB3Sl0gFcri7nowWsKdIjHd1UzmRYllc8HRna5dpD
0Je1i8D7q7VIzdUvYwzndzjqV8xCUcVezOdiBhoD1cLwej5M33vWSEs9FqE/rCKfrVRiMB2cXhOP
pBZ3C40bfqDRnZycrqEuTAQkKPSwCGdkHUaSU1tyoW5acWeSr62xajBxBP6N2/GGL2ZPGus1oGdg
NxEG+hZwH7lfDo2rHl7bHJcl1cK19YGQYBNAJmFltf0JDD67MkNGhHtHTjSP7nVEdH6EQo7d7Ge9
2TbwB7A14zSBlFtg1zVzz3TsBSQ1S2aVmr/2ep9hTKuhAmneo5078mhqMvhv0fDYj92DWCVGuUhk
kT9GeIHUKL/RlV02KzS7GBToyF/xar4gZGD3CQNWagjC5vVEQLdEK/JmY5ZrJnZPAo4b5HErDXBZ
NlJGDjSzgAX7btKT4LKlbzXCNSgxFxbDGie9rSvm0OGmTJgw2pU1+W8jkTcTOVpJtmBhLwF39Fa2
asuX8ASMhmpOI65pyUnAD2QG66tu7twf/6oGXGPwYYgPkWsJJf9R0u/GyY+YgYN924DYIYPO9y48
INrMANM1V8feenv5W7Y19eh0QWSwnDtkFaXoRvCOA/pIAT9BOo16ce8HBISvoEpECKJvWQa3j1ek
DhL4/dKSGWbL58Qv+dDWwo0B/FT8IFg/hFpGc96u7gqPjb98CzNCKqfUhenMLtf+UuA6SJHB6r28
vKmuc6YSEt00G5dSJvSw9YXJzqQj7OcDbG5ffBVxRJ7UIOIKDuhKqCoGxIOaQLrLIkvowSiw6PN4
IDp7dKv3lcuqtIy/Z/2SRUsWdbT5WcKKfncSqT1drGob+oOPSEt9HeMAIWzGnsPcrN3R508Q4m5t
69eCuynEfSmlfXtkkz+8hiIWUWxUVqJM54kxB2QdmLRGbpMzIfmkY5PkfrLzB375CcABCFKBfoPc
wEDzQb7d3xAdWACeJ9mhvvGQmK77uibORw8TQDa0jYOfNLyxUGXX+QWrgv4ujDGNIENJvdEK1WzY
S+6V/xpNcYhwmHTsZ2jRsHSZi46dr0JuFCoqw+XKzwz3SZ5gl6Zyi91QYGWHWUwCLeXHXIddSAVl
tRZJApFgz3sXwK/asdWZoQDt6k2ibfP0sONqdf78FphMCpLsugCxsl/ouLhWFtlEJbj4tMbXvD+F
yx3kOEaSdf1eYo5Kua9RPyyxCldx9dzmJ8IL6+ehWZIzM408Xo4wAEA33jNQS/vujs4nVCe4a4eR
4luuDc0Nj315G/IF48394q8Z3hp9WfS2+M6llKF8nhwKmWawZxOPUNuygW3fmIo5LupWb2EyeNxD
rjHl9zOyVKklYLsC3kYmsLpCFSxawst8pSOXb+UzqgwZsTUd40O3gIpDFiVVJlshxybGvfFkLAfc
/9q7FI55Nvns+RefB8SMAsbRlL6gh0u92kmhFouzDdWQqdqAe2oT/LRczAdW6cEO1CI9fX3iB4PC
AOR/V1CVYkTjWg2JPDrG7j7DhPIxTucAJIhKodkQ9iObFko5ejOdrJGWqntRGts5UFkRYVwi2op/
/LfRavt6PCZ3hVg2rbeNnKJ9pv2T3z2PLxJRzAh0rOxi3NK/bleKOvXcy8p0GSgylPl+bvq9cTCN
+idl+G7y4IUXLz+1zy7hza4+uPQuBtyS0TsqpP/oiXLVUaF/MB5pF2tkGq0sEX0+LHx6AlbrEmBi
aj93Z5GGngl4Vowlxxfi81oqxXaxuQFuNxG+DGgIk055/iD5HDIxqkHDAghB1eqhV6W/7wAF3RMB
43L4+mHV1NzCCv7AMyvZeNPrYwfS9rgHmjgiPJDFf/Iyuv3nI3/Zylt4JAvhMwALHiDpToBkhCZE
ufgfJrCnTa++zNCiuK9IGnajDYfuEBWgr7j8j/RfmaWanaN+O84VbkKFWIC9q3X+Oij27AsuCJSB
coX23/3HYU20bdJAFYshXZ61UXFO60uKHfYY6618ycgzqwIE3Oql4VibHHH6+q2cPrRaJVazmxuG
YIJH2vatzJ/MSy7EXl9jzdJAkDaqmASTHA3FdFQ9ItbB7Urur3zUC8BZPYOeVXQTjZ4ed8tzFooW
n68swXO4OeIV33/sGmk/AtZn9D/gmTaJslTDyeME/K+XDXtf8PRTjFLxUPH+L0RFWRWFJsLA+YaK
uj60Zgdj46MzT+dxVwb9RJdVa8BuGTz7s8K0eDpe68aUwPIIRgQ04dEbl5y6qRoM8AlTPEAJDnIX
tl+AVRA2VAj1ARkMBSH1NRr3AQKv2Ui53qDjwnteIgKCeuf8GmrbgC71OvlcThOrMAmKyiVWOavu
35OezEh0ffGag4u6NhKPdPdA89lIxcxfNEBUZG6xyamvHHgWaeHXeAGhp6Mw0HgCHidHebiA338X
tO564nqoF46Jqd/Se/0oPf4tVbMMnJUQmRtzq1isFKK3vYtFDVjXt4c8MJ62Pi+ylyTk7ydsbrDd
Agkc3xo2sT3IL31sozp/REhev5mrLJ7YqB9UZS2sfcOSOk0cIQrOR8R/SoYaSsJ2/m8tCMdIk6ii
x9MB/a2EmfExwmbJyelTr5TxG/juL9QrSl7W7K3MTTRZUeHsyWkE1HsBa1vXRrnc8DOzgpmDRf10
j+kaMuRi+4oeDH4KwvtFVbwIQwvkr2lkYqEjQjUO0IArnsbY+8dC6+iZdctAuaiKua+P5kONagoZ
Jb2J6LJqhZV63nBEDlUINkDsTtOL8VrVxwOpMXjSINxhP8tm4VQJFxbD7jZAKclc6HwvAFrrMV7K
Ro4sf6De7PsISpFk/LsG6vFANZHpkI+2DeThCN2mZ3yshMPhliNkT4gmJqnE+IplED4O3eqHQN66
xA12xzQlSqQseq6ZRU+XeizP7EUxl23fBj9qcY37SP7vHoW2EEDZntymcJQ77+rGxBRH5kZll3cz
i1CnpCXhj8RJQ91nScDrFWcB5GAWXY2gOWnv4Es98YF0S8mXhEB1Exkga51yqE3lethgp/VItwis
d4z1y5bDtFjf/SkPoPbskk9uK+nBYnFuO+qlEPEkixkYA99VzCGB9/2tIr1Km4LaYGH9MIi3bLpD
qjc/Q6RemLgB8d8DU1gusBMzFfiA3huHkFyPY4w6A9VK/t5IacP5eVPolBL6GnUp0NEij4c6CNyC
vLr57aZIWIwg7fQGZcsbUwo9ju4RLqF2VFnHk1qdrgAlY3cIkni/NORvlBP1MOAbZoc0Belyt7Cy
aqUGpLxMJLznYEteQczPOE2cTOVksX1RL4faY1+48y3UC/NlfZa37yKbMOiFo4k5/RAwxNx/P1Od
rxiSlOX7CPzSFW26hSP1eCDso/hvGCLF2OaDJKrjOqqK+s71fv7syYh09fVJ0kXjUQX3/2I+1xEJ
oWYMe/TPki+Qmeame9KsmtRWHNi68ZrI5g1wkoRA4KKzEfZCi7DCdqd/SyA0W31u5QrJLwoNRJWe
Q7yRHiD7Dz45JtBMxAZMWr8y5uXO2rVwFDwv2Uc+GNoRk/UbeHywSew9sljMPQNskIs/NAfuiTER
tA9KENM9LzMR68vaImPwWQD9dtsJqEvk0JYMDdKsd6EjQpWTKrrIoOQ9DirIupmfDh2ervlvjiDh
TVRSo15HQ9ol+UADcdPMwIB9Yucr5qULEnMizJPlZydbAmS7u2xMicA9giRXER894S+ZIRb2LTVm
NqI6ya3FUBMCk5iKyr9dAAgT9McykD/RetN88hICZWoHPkpBtu/QpXKsbwOsbge9XM+BOGRoI892
yPYyD4edRmEWh7ScIbeURkW3Ssj5UGgOi1ih4xgHjq2/udU1uf2vqVzFwaxdUGFJBGSuUMFigrmV
nsI95/KX//b2jnaS4OAwAG8bCEtCV9jbU5nsf8o9uIBNKPsJTA9fEQ/cD9miPvS/UtiKGBS4rUwI
iTwef/2njH7fQ+dqIst83604ONXa8P4TtyV3wKsXnqoN2dkHosC3INDhFOjr1oWgKjheG85chPt8
YwvTWBPzNL2w9UQYF9mIkbVYj9R17fbCdog1qLLVIppshCyWXdmgWLpwMFQEc8kiRSpvtcucJrr8
H4U4kdRmzbbcSVgHT+TwBhV/hEctio5mIU5K2d3Wt1EyASkp9L39xJjQePBWk1vVSFKi7zlTVaaj
RehzExZm2Zje/9Mhs7qBBt8y7AKTJaQHo9pIyaZXK2WyEdLpAeopI6PE+DzI/ieVPe5+HKxNa25o
mcxzrqKTLRNvvgSVXoPbRSimCu2JYHNlgyiWSLEE3zNGGrcxhKev/m0FQsMAJ0veSMGcCgss2yeG
goWagKnrTet8cczXOZrN/HXBhbG9lXKeOPvnnnjDeXl5qpbMAA87FjhJUqnLSWYPT0dKL/gD4STC
5kQ8O61L0VdEfnZ0G8CP4jFNv3QfdpKq/qxDrMjKJFyA2pJiPwJjWfWFVyqpUuo6jTrFin/UFDJR
xpFYn4/mHpgh3HHLOAqEG4QxBK+yDhiGHNfDli9iLq/fvE3y/ah3c7fdHwLUg9QzHsgv6aQ84fww
wqY8gVB1XNvgFrF8eIACtwu/BKDlsNP7g7Q4NN9IzyeSz7/7Z1zQoiknImqNnyOWNO0z8TkQTJtY
uC3TOS4ZJo1101FlTgwGwWhINkPjf+16UQeRGAZGSJP0WYoX67Ilra/dXqonfZZijRUo8w3DpdeH
D4MYhJROAzeCHTMNEgu5eyPyU10oh8ri4jHiu3mupG+8NehswyRGXJ5V5VpNQPtltvA0qcpL4bYD
SXrg/SRc5IeF4A5PbZX+L9zZZCarmUvm48Xdfgo0KhzYnSzj0a5tKvfkNyqILB96+q2EnCuAWLjE
TEpsLavLQEegV+Jyq7M9xw8n989i3WqiUYzB8XOJvVnFlwzawhEy7B7jg4O7mKPstvQy8hZh5ZQO
inBf7x4zLaQy6rmliy1aiPQnkRtFXBH7Zcq5r63C6odKqulCMTMBFmWpveZWaLf6aNLYdF+Jy8vG
pbeFhbtzChirF96EVzT43Y1JoJHpQyCqAizsamvzltJ/by92xPUROj+DkUDjSPZ9Y+w2IS4iSX2A
93AK2Da3tZHW7hyUMaLA5x+VfQv8gNvdYINE6lK6Jjpv5VCUaM//kAjhTM8SNmdk6xzy/NmR85C9
sPjTuem4ZgYntJOQI3hqsDyMkatquBmtYjVeEy0SlYNjSJ6jAEmnd2uQrv+5MAfUWgmc5BhkS69w
5UYC2pOYXyrky91YjagjWk9YF9dfqQPOPU5ZFVyvgVuTzn/ZT2FtEV/C42pk5s6hCQ0ybwUq9q1T
wpGKCFSeGrLOi3VyB4K8S3fLz7dPL+Nrm4iJXfLHsBxX6GfyOghTrXDfHygc2NRdrAhpTg2WPUk5
xqPKVtrivwgRv8U6dc1VbpB98OU+xaEFXtrAaMSOxKXcWj57CkQdXtYFY5rftvXmz2EdtJHZZa4J
VqLLCO2pKol/xDUlTPbeTLAVM1bJAXtQ/PHM4ELam1+5KMcFv/KDSziK/D6q/t0r57zvD2Xioh7y
uJY5C6nRHYheRyb3xrjiX6N/8AyGx1AN2Cv1iWrUEp+t+mvn6rAVTHzHAyuZ7vsHTumYqodkyjio
qgk+Tr5ZlmHsueDozbeQCCHIrWOAT8CYNUYduYxTiHkL5BJ5IxcZltDSJYOX3hrTITmy6HIwEaOn
5bx3oHmnYIJLV1ToZFS1BBktQSfIq1es1VuNXztqGGcREx6p10PBkYeRnvZowmio0Rq9mCeuq8T8
mpjm/AkgHRpc9Qv29Ps1iSnCias37lpxIYjTND4bwsXReJEsOZWBh6pssb6Z1L34HZdvAkNIYSux
1rrNlp6rrjd+P9XXgJ6Xtc5K6EKwSJ48/9CfWIdm1Py5Y5MQm7jo/tfs4EJsM2Xce/BAhtjd49a9
fcsau72vY7hBecRn9Nbg5CNAD0AxUhsFjTSbYs/ILZ8iC/6zZaWnBHwfSOp7DGnVt0skIogiYZJd
SLvhCPA0+Phks0T39pPH2J4/JglbhO/jJ0fIt8VKuP3E6yh+Vn5BWCpGlat5ccpokqamjHNe30M+
HBMMJX79J+aWwSwmR6ptGkDRaYbz2kbbmGP4l+gKqlOavK7F/fXQn7lTl521NnoZoe6WHKYcBl0l
OyQS/J3BxxrQ1vj+LL4b8x45BHJC6czKDBJd++C90XWN6p6F1c3eidNty31GO5EcuY/nRba+azh+
MxauvEYbaHmUFd8HcImDw/LIYQagxOLABQSpyBvZ3lejkTVdJOrIYOLLL03eX+yEpxT+Qt5o8iF2
F6vHh4fffEORyRg3UlVXKpn3ShP4AGqJSyCxq8izN2/UF0bqcyj96D4ELMoIEjI1DWCMXPDRcoZm
ASVNVdZ4oTJoTasCn4OfUJYpyMpZ72a0Gh7A3sC26X6EhsW74SWGBfLu5KUlXWheqV+BZ1DLRFfw
aQmkbOx846meTtCsXno0HEHG6K8leKOyVl8nfAUIBEWVVQWwaXvT9PFqAjzEBrr4urolWMupK5N2
LU0yWP+lfyU1wUHourf33VF7ZiL1/CfucSiYbbhIs2PQDJGGXyGGy39RsiatT20jQ4A7/04y1GU6
2+IlisbnsW8xeczXQlOX/1Hmn85TecGXv2a0T8i+6ziwXN2LTJW0WSyFkp/tNYGoPjBh7SIDV2K7
VC7KCf/+jSVSKgnuP7vDfJtkANxL6lkTJj/73G2QgGjzW0CIMvMefIh6i70zgkrpLEP7/YFz+Tvn
ln/KQLIyP3TfmT2kxuOkQzCXKZJB3Bptm6QMBJyqQXc+2TvgqeiFAus0hODnASRzwixDJFGKzCDt
KB/KLido8R6unkXMKyFV3dP2RXpYdj6dqpkjgS+nnk8Pb+WJlIiSaPPeFn+iEbpbrJOhtXg8xDa7
PLD0kUIqSMOEatwLawlwPFe+96hLu65LrBLOvt2KEzXLG+OPhGcpmTy0fRgEJOPUEASFunR8I5fu
RHyRkbCwkOPO5ek2Vr8qicS3MeW0QCh6VYiOlqZdpVBO81tTewfTzAkLgA6B+5QoTiNvtYdiWjSY
ginSZMIFWyu2o13aibwjMiNAvwBRzlqIly7AnDtxJ+AvcsjQchwqmw0oq8+A2DU6Y0/ixmmegXQo
WtSrdwIdPHshngSoqeXAWKGP8PUE0R+znTM22wpcR7TwNKwqWmyilJOwHX0aHsKD6xqtN6EVVzmx
ya37BDY5/RRg1gV+Lt1hFsLcPh75lL5aRsxthx5Jw9SdFqJvqlmntC8Qkod7FmoGXRTuszvmGDOg
QbLTYYTMJs2RxWyhW0OjyiEcmaLNvljtzp/g48uNdHEv694nHSoR5WGXEiYW0rSqjadpyXJT71tA
JZZsZoY08iVBRIWhHBfGK39NK1Jp5r3f2FsLypLU6UeAu0i7xrQNEw/xCs1ySw++Bu/SAsCLS7Tq
33yceXjXHSc6i1vJWG83XPIshp6ES63RIDGY/j+Cw6g04dNWLscFNRDzccOfuQhMmP8V0DA8SRR9
Br5iUx3GivaSnwWmB1l22AV3QynTZUvhHX63QJyaqazIClhMBBmr8oeUNXKxDUkuw3PPCL5NHXcw
ZWmXt3AX1zVqplBHe+s4MBBq6lgX/gu3se9WgGcg9poZMx1TEN1+zvb+bCL15kcFKbV8gluqYPil
LMpZBKv+VrJp9DkE9smblRIwFpkauJJbHTA0TZwnF/DivNYpB6WUwmR5c+41hIzMi17OMVUlitUD
S2L0qRJzE5c8+cO6lXlDFcQQ64MbsZC7dyLwHYlk1ysebZoTguT2UmjZvEPJiskur9TBpFT1I2Li
a45Q7RMOJVLAVOplMi46gLw0lYzgx+ezI14woNfq/G8pXcO2XTRbacqKXbchtmig6bM0SMWwNgxj
qLjUDtyYCgcRulL72oFcj8sbM4LzR5RMsML7C1w0WwnuCdhujChIejOLteLptkZlzQd/H1b4p2QK
/ChqJoKOWQh/HuCeOsjaY4LDhhIy954oyctpefjUJm3JfwH9Ww0815F1+z68Qsy2mGnP+PgtU2qT
ZIMUXVAfm+MpwksbrRz6LFVs9hEIPrMq0LcB9mTjYXQVFKwxJ/TsX3cXHLJ3+nspF43sgTRZtooY
fyCuT61S7Tqv51ZKVVjb8Y0DmgVuMWyIo+XJXRbuEWCn1VW38RHlbcunPtbglvSf9e5Hi4R5A+lf
bkIvR3mKjMogMqySqTDINWYD5+PJcXsdk6JEozyWlxz4d4/YLnJoE7htFGSHAaF7UEGZGL3nI7O8
16fsgGfKCeuiwseEAje265vteXdZHjJ6mYRDfIiMu6gedIoJk414L1ZRuSygK+VNOpt8Fe0RxN6z
Om6m6RWCQmMGsbm44aJSoCqioGrWk8bHQB+JkIetwhRdxygyctpZ/jUvwTM5PjmVwyredYnRR3pg
GmoHSh5prGMSyURXlQFIZfXb6yc4jnrQedEbq2YUN3jeU7W4EY4/g/WQK6MxPvHLata1B9riF044
jqNexCHmyPgNVXVxhKwulBKXTL0tyuou8uq5+j29bzMrFx7K0D6EsIMLisQvOXqXShHR6x2ByPdZ
iKbT+FlNIGd9F4yjez8xxjPTm9J2GoBvV92n8dEOWRL1pkUWDQm9B/OixnCOYpMtzF+WyVUbWR9w
StosPFDLkJW7zLizlw6KDJPfAkjUME+k23WEA96+GvoDcF4fvKo++0FdsaX2Zbmlw7zTsUZduElX
WdSq/9V0pDsBOHJG+zyDIqGS2I6B35mDbZmbqvWGq8kxVrp6rUN7qnPHEuF/gffrQZw0kDdVO570
r53xznQfoT7owJqUmoGnQ7APfioUvO4g8YR6pgYEOIp2ZXggkp18ex7fhAl5bJE3v1LEOQ5im0Gb
7oNr9q+4uw7BG1YQBfJ4Z/0vLcEklyw3IDRw391ek4+uXhgyoHHcNBMo2uy+50wwowMJ4kAfL0jP
uu2gYlfuD4VtceTS99gYXwNlNTj5/kpmAOrnZMrk2jIXiYK6IiCqwdQx1WutWrK1l83+iPu4VqXV
dLX+TvihP6AhLRSilBzI/AxH72FNq7oh+IEjjIjG70y+awbIXkn9EAkLUdFhR5g8Kt2l5tY9ubA5
0mXiYHij+lmdiCPnwMhbhEQHsODN2etVE/7L/tMwK6KqbjPMSVset/axF0PIPRMG5uVDeUYb8Smf
ssYPd59jwA8pefZAPY642qw5KWaQRV04eI1yNeMY4J12NyNgAge2a45/SQTSIk9K2+WDM3zO13d8
yc9SVjKi2iq12PJdExQ58P35A3bUOYoNY/xoNHLEg0BK6YeCOPZMBohE5A9HAWiYPCIFm0JIncT9
ZoVxClD+ziq2Hvg5pytY8Mb+3yVfZyrd3Iqf4EtrzVdFlFKYfowobn4rgh8LmFqaVVlCPTVxsuuV
aYEWMHrLh51GcpB1Oo1h6HR/jXAJ870gSOxwGsLi+5IKEiBitjeF+dHBbacDqmvB9zPus9ym7KXf
NdyS5i/BKiP8MnU8J+VVDI4wBThwYxYjktS92kx63S1mAjL3vbEyPR36Ga1OwsI3q5nG7hsDxsLr
jOzGGFxHDO6mFTdXNI5AlRYJyPoo4oRwI4WPYmcjiA+Fhr3KEuxsKhKQuO3oyoY8LbBJROg0Aizj
KfpF+wRGkkk7i6Kgsd5Ovgn0wdYY2epSHQ+DrR2fP2wcbr//xw0R6gHCo3cXwGZsMFixc9cMYcPj
AzllBs6pKqMhYgQj4z5Nd3OGmL9Pg0eT/O6TU7uXdYOx89yopFxNc+KgWaLKwyFjv/DXHOiukHdj
LtIdSrEgn5zOKC5jiKtHn80PLUzzRSQE+MWHiwApQJl7a7DzORvxFwG2Uu1/8NxhU3bZSR2Gjozr
/CyDjqJPIu4b9ge27+XvGrtFCpRUnmUH8G/t+nMhMeCqyGvXwKngBCXMBcYrA3+9AOta7OMSlKKz
JzSbmKnnS6e019/6CEV/95YFefdu4YTw0bbYKxysxsELzjon0nl025RvO2fa/fPZyaU1mSKT4t1l
CtaUMLcDzvjHjn89epS5m+p44jmZfwzw3a5DHssKEf9DorOKTPQHUiDF0Fdoqc00SXITf8bGre/9
q3suMkULTzty4WbBno5uTZX/lKGEGB05mBXLS02rKdQsx86NsCCnp4Uh9ckvTFw5FSlbiSyoItTX
oW9y8EaRF6ZYxGpsmH/tkmU64jHflsM/AFvYUEqc7cBdqVIM0omtCpg9UXeabMBEP0PlvuOJz6Ci
LbFYOu7xedAuDG80pWTrGaVAje4sFN2lmv+d3E3qMw1hyl3Pvn8445AABeeoU84wSUgvazwlUjb7
0QCY9wd6/gUNN4IphCq7nbzdG2iLAX0TlPiyVBgSmynjBD5s2MuKOMzgaRF8xU3wSO+xvZ15sgiG
vaYDygMhIcTAOJorSOJH8FPevDrWmzHxjKYv2WBIcxJihHTaY8LyAq9sdAA8HMUccq+vSsbb1egA
gjLcOVrLSuBk8ajUjP8CpgPK8zz0PkCH5DoA3Pn8D0IX6wi/dwbDgkCjSpSDXshEoLa6X027YDPi
yeoZTvsu5MsnqXYt06IEJborJmSwJ0OAySsCXSodhY3urw/ONdxdo57XiJSQJxm7JhXpDri1TO0b
OaZ0hBrIWCoIeMB8nvBbJoVC2ErNHtAmVejv3s6TIJGejwCOu8x4lv4qq+zHx2uoZ6ZtVtITPaSY
w9wzRGnfC6HKv2UTyVD71pAdE8DJ4zBt3V0VcCERvEvdYrK2AgSdiC3dWMPfJg4N7282uxEnhxnD
jcXvEQCFsMpky7fXuzlocxsIeoxKgqF8H6JzyJrMd4BHrtygaeRU0WUk3NOHQh2LIFQeV7nx9B5g
HGaZnIqJ521PVYsHcZYkiIaWNbbA6t1+cM1vK8gksnGKdnCkyaGmy+/93sF7MMGh17CKfIcYd0Aw
COPL3vi31C0hiNYAHRoKPXpgycFfRvc1TvkdquLGlZoLQrcG8cAtzvDWjO9djN1uIKQyxFa19o+y
l5u2yMT4YyNYGLUVNO4A6I/9atfzrZ/NF9hYgP8L1rbPwwwtXuJMJc+gUgJwoad6ebSHBpg1kVdA
YZrki1htifedAnoqhgEPMMK4ZTjxUI6u5iF+QG+ZTZ1Xd8tbz2IwKX4CVYAoP8+T6B2j5MCOz9Mt
pSKf6D7AAAPpdd7OPhBcue6c3yscUWklzZyhhYnDLGQ63H3llTxZOljUS298CMQwNfhX/RVPP7wS
iaOz+iNsIoibGMfCBjPVwuxwAcV7mfMvKmPia1RzSUINUNnrVsJEN6zK2MERSbrvcA2k04wILp31
bONWLXmVYwhphK3tc304URxnSmMJWlf3+Rs89ZGV6XCJGdoQJYnlDWgZaGIDxzT9nm5jchvzUa/T
7ThNZytB/nApg0fccUTFKUEnTztRyo+p7rC67ToVAFm+yLu6jFOt+JcjY8TaoWLkkVO6Aza3mSRa
78KZfNfgcA5oKndEw6AwA12qocnDklW0tEp/N4UxAjG9F4csldu4EntTea4uHKzxzKgeczZoVm7g
+BZKDSG7JDtWPOMZaLZzrS55Dmx+fvNM8Won2opjjnzVRtvumg1pCneTbOU5eMEhU/QlJtBEU4ku
gAevkPy9b8gfXE95ySYXh5YJ2vWnjulUmhk+Fk/2BfrwYkBlfMbrL9lDrzfa69lbn0agyJzKZPOv
KGqs2vM3FnsNZeDd71hCgBaO+xNfVewtRyLRmD3vKZ8MXK4NF/1CSfxGOzjjLGKogBLoMHjKK5kK
CjgHkf+U/I5Uc23+1fNaXEY5AttMUbTxjE9LWReazhEE5Qb/N54C9GSQ2fOiMk9EmQ+uEekDu+5m
PXtPR//qpN9v+faY+7mB41kAHhhshFqolhjftv/4l2NLF2sbF0SzzNDquy/WdVSAKWmNzYWpARwx
Xz7uQoet0jZK3zQIqwR0nOQOUrEot0yc19O74xYr8Pfd8I55b10iv34FUblKM1NXw9ViLcKNmFNy
7S4jfFj48MeENBQsMXCzDnKPJkSh39CF3W+EPL4AmB4nigb66xokycz/128qAWSPiHNI5UIdQHOD
N1lqzDMdbE8t2ATTCPmjgZmJBBDuUBz8UPocfeiaipHCL2lcuscglT77O9D106w+fiCvrwCr5Usi
7lBUu+J3yicPHdB/Y8OypnZeaeZX79AfcZWD8BbVPdBaxdREnxkUAOCY/d9HHFKCqNAjUTrp/YUU
uBZaGbMrH1jDBJQEYMoHDS8aclD2xB4dnIdZly/DXKHDKGbdzq3YMS+kQ4oleR5P+3WyGU2nCRPG
lcG77SgA9MsNnPEys/5hZF2UUdBGP5XWll5Zy9CJ3VGaHsQHejErPn20Q4JJrq5QlLih+pL4bH8I
Z9K0fKxuoMMMpnm3EnZkA890EzELjBIwmXsBS575oiq268fJzifyk+Po36SgKDpnVoNkfk++SXuZ
W0U5Pg1tMlhfZdy3R5VwuBFY9TaF8B7lN+2okG2YmCb9duSPt+/ZDcY0kPPFspti7LXKzxdnQF/X
qpzN4OvMyi1QlKUuLG4Ii7qUESMjEmuxAoDMcRVKK99FS2h8zSQfTeq93Vv6ESdWhcx1NDF6aeaO
rKyp4w9JdxIS2wMdz1pBztH2V3TWvmPM9wQvtSP85sCo/L16aVK7ZK1XV3jV6XtXIN6AigTjd62m
MMxO/KXdkb7av46fq336wlKsWJzmccxNZSynptjtcoIHoja5YXmqEZ8rv+/QpR4eaAVZuqEysohe
BOllln1ZyNB/6ySp7matiWdarMlj8DIyQyeVvzhSLUE5YJpr9h8pscw8PctM+Gw6PgmoYa0sMpQK
Odqlw00Gszwz6Vlf/YASxOHHqrb2TwzXXG8WYKsA+15SvLeSF0FUA8mXSb+maDgyFd6UfftYcjxH
TTekpDXUeodN8rfNd33QaD+i3YAOL4KTxm31vSKslyAA2KAffGAR6reb+7PqHt7t/z2H+twDMFXX
qIAoDlK7kyBF5ASAcHLhkED7Rbj8tQRBppdg+W6JiA6of5SZo3EJ8CXXpxk8d9nBkQ1HPomnDzIT
ArjQ6lD73sZZWHb4jpOMgSUUwkwG+hCfrpg6NzfcmgOmbWtq1OWltne+Dpeqll0h6RKpAK37ffkO
p34PJsaCu6hxyauc0MJa8cGpi0k1ARt9ifAcBDuJiWPJ6c6Qfh819Sp2+emBLAwfx6SxSz5dXJMb
j6cObZ3j0QzxlQytgFMfwoKmZ6ZJxXsV1e03QH9tLgqcu34IFLQMcfvOcZEepQ7O0U/izmbvNprn
OFaCnuypdxFsT52jtxzRk8QG+VKGu3M/VVm2isQMLkFqLLMJTO2WQr151+pm/pM0CVQqtZbDT7YV
CkPgAPvLpypIqHCSXOn+1QNdVcx2CJvyrkhAaTRdcZx1g0lBm//97m/z1c5O/z+b42AjRwYxfCih
qGYWK+0ciDFcdoFWxAcDext2bjdK3AKRNpvRFBkNdd6kIYUx9cMRpEcUJclydG5Tm81vFaaWaYqt
nu8XhlecW2sS5xUWi/fLFwM4VwUdWB2kwBmJIAUAm8mfHXM57XpwbkJwdXuPEmC/MLmIfue2nzkC
r3SWmqWyTlrzZCfwbypqQLTMxryv2IPt/Mxb4MOojUmAWKuy8JpRKSniEjy+9L4CNzAD1BFZA2nX
NNTo9dkz4ttHgP6HBdR8sUnRB2/zqdr1XDcMz6GJDu1TCFJW2+hY6a8RVA341ZpecfyEyfp4BqV7
v3V4zEbkYpU43YFtHke33TwgNGMAEOm9v1KThE+/QJKXlUttNmwpbEzReChVr+JXBLexHT+ycBSu
KDeNKJq4JR5dSs2AvwJShYRRNLJUevIx2TC4Xv7KFxDP1sDxmDieKPgTJiEGz/6GiuFdiFqWaquT
TElpYHbI1zbvuemflF3usuPH1TF4R4BBUYNbFHLYNJze54/YJz5m8jvQFVPAK4L0ZLCtxMh/49ZD
HvLlDzSEuUe5BDit69wo67SBt9rWoGGVWxzxa5A2ImIeOwyTj5iOPE/ck2aMjZT/3PC4i7q6H2bq
s3ttrZCswulCN4o5fV6SznP4i5tUfM8g+4+yRpw6r6yAEqA5r40RoWooCciaZN9WtvhcaOANCDDB
2D50XSuVPjhxZuQEf0ffVjus+4Pk1tEYyb97z61eLK7gO6R+BMF/7nDmewErvHeF/aYg9Hvl73uf
xPVRovc1dIi0f3F6/NFS6qxvssGfDz/hMbTvdzuYp0LskwHOMdwp+EhG7DRRvrpmdfgbuMJHRFUW
71rGeC6o6DC2D+ZvB/rBPJkdzIXfWvb0xN8MHxz3uxibT0PJeZfZ2hYAjpGQhRdQ95MPyWRCuv3G
EQjmia7+m+svrUqjgb2ZtQZoukb9hJc9sxCNVFyPVDbCe05x+1g+uhb8AIPe4YeDo2p4NUPp7dOI
E/YZJLZeHZmhpnPHXG4m/ZDDDXh/52HGXEU+vduI6IYwsLdic0qmtJt0JmcnrXEbvV30MrlfJzVh
MS8B37iUCm2r6pFdQqbMhtV2l4P+MIPKM0YtFiBkq6BR6SbXo11H+aUzbRncXPkiGUUbK+lmXHnP
DJIuyFx9TCz7jpjaEk++aCarUJqNcyOo9RymXHaBwdaGL+nMwBcrHfiJb0kJ9qp9sEKTBVJ+yOzE
SexmusqwzBzLMuciOIZIKjJGIEM9GetsTt3YmG5Z063gnNO055W/hHIGdGNDa8yC+XK0EmFi6km9
is2mCUV1bAe7sx0rUlSGVqXw9kW27VKApfjNIal872bEk+JbjrazcNRfQGSomeq0Uqhg2DL5NpIx
hDL+Zh5xQyC5XdU9hTGt9KPHOsiSAtbgJVgI7cV1NqiUYL2xnQvhysKLgMyKbLODq9X+WaLX2KAF
cmkeCAWehpcoR1fBp7VtKz+zeU+n4REphAs3ScG2LJZBg4Tj4AQ4zC7zqRz0dEi+ydodHEoMpyTE
y9IskiOE2VbhscdELtm1PG/wjFtaWpZ8h5ZmE3Nv0K/cUQPdE3UPZ5q1jGKxeaEVXzZazrDwJ+/l
XTG5QtoTcBCm8Yqgcg0Lzsc3ONzaCxkWWJywsuAQDDt84kW3lUP9BdyN+YuCRXNFqmSneg+Yco8P
yYqIAUZZFj2rZbU6stZdUvf93ONcC1QIvna/XO7zFKSnj197HhzhKfHf0/mreqR8DnSteWHLjKfJ
Kj4+LSWfLvC+dFaZhPjb+wU3v1q6iaBz+xRQeen2OtVpFpbtl1H2Z870rqqGS266cxYDnHxi3biW
/vbfaO1BQoWZikHEMbmBvbDK9+pijk0wcUYqn8sutlRoRnPzKuDKDdnIlKjj31LoR8Br4LEK9l55
DfhherBLPNFm2TnRaWjC05Yt0YN4IxwVWtMsPSoZcrZi35Nsv/ZVRvPev4Gfun/Qsc/sb7yNEP+0
NPg/wy7VT/8TgAI5JjTIgX8omvGigukHIgYA+FqKCNaWuxoE8Qf6GpTqXgCvja6NTeNff1igrHxM
ebcwp4GS61Zgp6QCD36DJBoCimcNds66a9oO4IBq39bJ443hXo6Z0u420jsSrtSrEZ9ZmGBiwJyr
coXenAOIRWzfhoPC7YTCmWWmAvrH9HpwZIyRm+nA6VYg/wZKXsxnanilF/JevmDdFo2y3DcZGnOy
F45mMkEeDizF+LEYoxlXJP+tvK96Cpny+FDlBsby5W8n/O/gbn2Y4PTihhPYd4FfOLZsezllK+AH
ah8loqyBB6qGlgfnMiuqoLfU5OVvVn2STbAMGbUsaPaZkSnhGIK4ETS9u/XkfMSspE7KLMPN33ft
M1HOUQr5F5IavwejBOmLoV2asE7yiaVwWKji8c3oBjAHmY+ChYDQyib4HdBOHl3pOUjN5yuRTydd
oEyBhVy4b3lTxT6OHsycQh4gBnkFsEQuGF4OpZEbdzBSsOqXb+mtuWTVPlXc8jvcoOlADwSWygwn
BCkfObt1NiAVcyMsuD73mxaZVPNKxwmELmpTfGRsL3/s1lRPXyzLFpappRtkiumP6CjP+DzVgmft
BrMJlj44lbitlixZoWUaSkYdl+h7kBLhGaM1xQV2CtPvqE4p2CZBvH8T+YoJiwoAXewUfLI5Jj/W
iVId0p+C64tzHCtcOnbMyOHNd+6lJa1GB5jYZfh8AlJWP2K4F4OhW7szJiujNXjP4+USG/3iatpE
c17PPa8qT39D+rb0V8RppaINZ4pBx3PocM5TsT6IVW1QpzGvuKbpXi2GcMNRKfC3Qy7Ni8yutQI8
CYkoDyEue2juke98pTnBHfARq2mnO7NAQL4ZwxvKfRRIzTdIhsaqxW2h+rGHQgzSpuvdk/6G903M
iUSh5r5cbFzwbeh6YQOnu8kBVZwX9n+JsUGsvnD4eexnXW3k0cSxEPytJfwpyeXC+PqUgUbdfQxk
Pt/kPFzCwAJGEE1x8uyz+VKac8dISmZAvWikYUqkcphqzzC54Ur+rqn4PDy/fmSgVtHDIn54FNJg
Jf7hzq0a57xmpapWrw/9Rvm7wJrfX5L0uJFpatOFH7m9dy4y8RBmonYkMmQxxCdQDA7F5xlReaXr
ts5dqFCp9OwCpmGK1+gqfFxM35w8yFUFQcau8U2KUXeT3CPFQ7IhZ4UlLQGrxC72GFtRYPwZ38CC
SQNRFblxYJ09vLhDy/Xed/x2doRHkQ9JNFWg3cS3W4iUet+FShXKC9EYrswvf1IXOiWqHoBOJ5Xm
fQR424lFvE44BLu0/fF1f/S5sDGpg+tcxJejxQj7giaJz5uVAGafd/qVLUMMy4JWUoK8n0DIcz9C
dA8gl6bVGQuUSMIFIhzBztQajbQwH7NnI94vuSgFgYwJiEK/BkqQ0jyaoix8BRfcCa8imnthk7Tv
eXhXpCFPL3SYbQM190XmJu/BKrqEgj/58PTDuwIaQv5+hqmwWesCzRZYAmFq6jjmNYAdYVLUxxlV
ZdFswM7SsP6F93BbW9GJQuOj1STqg+YxXa6PeFy4xJJ8qXGdD8qzuGvS89v/5VbtYY0kNBbnmYjy
/rFU3Y6hAFtfuM/bQXoNDoPMMUpcAQ62uVJgfp548XtpvdIuAustnt8CSzeDctaRpQiThu+NsD3s
Z1R4YJZyhqqTED9QfwI5hW+5CobMOjfxUIZEg3FbfiFw7gYV7lUFDJ0SqEGDpNoBdYUC4rke7s0H
ogG2zqaP2x5lpRP+bzztYJYABWXmqH1W9uMY8cQaB3SAJrB1N14T21fkaGER1QMRXt4wl1i0Nnub
nlQ+e3umJCsRjAAHunoixNpD5mvTe+iR+6FJh8zFzuunctkPDLiekQ0tpS58OYOVtDWAeyJy5EX0
LHtXcs/JdYa76+V0ykO9/eovQxlWRG1VboS3rh2bzFOz75jPtGUlqJLDkM0ut61oZsed9ttP6AQN
VYP4q8KJIi7Uau9F37IVk5/DaRDF0442h45gWd7r4wPd4kqtYeTE99XfAakfNOfCY3t3yjRTNC6I
Y9eiPGqSR8W67lZRfBYgXJC3BNEx67KZ4Yvee/EfBNO1lypTLhbd6thieDmb8tu7qL55yaWDrChT
0bcTWgjhKMtwUWyP08R6mbtvQmZg5epXgByKKFMkduOQoWMd+pp4USfjowQOqvYPQ3lS7KhN8gTH
82BLXDDoslo/9+ExtRDtoe5CSaRoY2Xo2+5v9es6tN1COKe3x0tnMtpGZiad8AGu8skzFsvu/Olu
jbCDDK1iopin2q/d38m8wGMHAxnoLn7sBvVtw9e1zVu5asTQ1O6LMIiOxXWWGpKWNzINtlOG2qIK
58yWrYIU4FosAuz/ETz8LVRIbyl9YQGap0OrlYa5X3c8HPoXNl28rvXng16dMPve4iT2TpP3rJrk
kn3w7diPWxsjhSvLsXfp9PDAtFQTxO/lgqudgQtb49DAYAlyK2hsYQemjoHedAzwD2dhVlekwq9F
7EIZ+JAd4IJ28A1WE32CPFmTmVuxBGl7cJBegOwCgh3dAcMyyc2LJHcyoijteeu2cajoitlVbSH9
sUv3O/srtVfDegQI0Gf8B5B0SBMcLATdKZ5facDYExZ7vrxs4sEag/r0ts3us7l9/VYIXoZlgdLZ
GRQ129D4IqD24tApdHA7N54smf8YdPn7o65toissSjvPpEy89KEH3SmPyjPm2N9Uv5zZLJ4Qrem9
FAXpyPLbAKwIR4ZtB+8lv6Zb09W7D5w8M78JQH71f+PO/Gu4SVEI0SoADASURBVY0/6u902+ghIo
Hf37jMN2sl8b98/LlLeWXbzKoZlTxKBmpsKri5Qzw7c/0VuSnVrpbzF2sF4cSMI2UT3z+6Rjzsl4
ua36DkzUPqvJktlduIAdyQ/wyoJYeaVLRQLXWyV07pB7hQKGN8Zz2N3z8BJFyL07rHFLeYaToHab
RDHqwZxrgukG4gr6TBItxlp16DV0+oj96jh0OMLs1xS04p9IfRXxMdLc8wiTPTARkXth+McbURo6
hOQrgF5M1LIp/SsPR6a6OSIIl7T9sEQurFVfdyaBks1fcU6KQyYiG2ROwkBPDaEKlGMTPdNiHcKm
4qe/lfKd29Y96OOdO1aq81lM7kYB+qmi8N9u6G56idhmtwhuEvMaTkVbNqnVf/hczUHsgZ2A0QM3
8Ndmeir/pV05qLCOVvJGUVqq1blF6F3fexnnWeRcculpan/aL8SuA8qCtfgyfvupctoZP7Ek2RTJ
jkkntANwwO4a4UFlB824j/DD4iQmCVQdqJmdAHMa7EzEUqDriUbie7DQtc5O1HardGL6LGlJpg9F
XroZpcUhd95KkoAYD/fC1TXeToXFa0V6QFn+yQdkAD0BTLlsH3vi5uoDZ0EBxx1SGbwZ93F0gv22
7bL55c6noedVOuZmvaIlJeuYX5RKI2AnWs0o5SuIyVSqV6E2YQJxA8RZJP2S1QHxxtLXzpTLEIMa
A6f2g7cgm4erwpsSQ3TrhPybn1KVmnpskEmHT5R9YkO6RCavMhW3iSVCmwLgOn1eAHGL/TKnMl21
q8QEhR1iYG/4LHJw/SFguUHYHqZiXstQPck7o3n6NnQZmWQLiVrFNalgaKYA2PoJoSYbPCMHlCQ+
38aOBm369lJnljTH65jIB2fkk3hn33vgR1As2b9DdKGgYvQ5ZIEkkg7Oj7TeN2Fyyh+tHQxOEcvO
5s8DMsJMzNt162xp10v9INpzfZGcKmOmuhqzkhSeGEEhMIgVujb5SQGrbNE558ZsPOmwVny9uyWW
u/sE6oGCDKrHYSSTFOjakRATHnMPp5vpsQus4Al7HCHZNdO/gkxGf1trhuozFgLqm3HM6+EkFp+z
NZrtTfRJjBETEsk3T1UlEv013cql+OWw0gzqc1Bfw7XqPQI5zkFoVXGSEtbNWWqHqPe90UVgTvxk
rbZUU1fW+TzrVRkWhzWzKh0CCs/NDvruHBxqx+dFy5yGTHu8S8j1P2H3UH+AevA/9nNF23i9Wwnw
LSsWB1C6aHPSF9kb0CsKk+AIhO2bpT4O+4O12bqLMHxMfC++q/3FHbBytjRmqTZYUu0wWloFa0cP
6IL0oXZpkLjARWWdXg5TsUdTtXHd7SswV03ehIWyKwqnfAVdmqaUDKJjx9hhvOY6NZY+SPw4c3c9
klyH6ZE1wImpFPzzOmmW47g417fwckO0CleibmolZfMkRDukO9DkZaNyYhap1Mib2Kty5hV3nFAH
3ovZm6zs/dv+IPUrGDNbdQD8XiZHWiDQM7S1PsfeyiradneNscEV0VkngtKgF5z1ktKhfCg/b4Kr
AGntI+Ca0SEsMVFTzXdfIG9jp3kdZoNGeGUsSsnKGjELFP1geXiANTCxd2ULoYFIKIc7I8yBD6Qb
QW/bw+44hiwXNl+qkyWmStHeUzjeQ5vEL82zuoCREdZM4Mg/ycrWJxohKuiZvAbtMxvkyCF6/vtD
W9nF6WNZYeLAfzqdJqsXSRQCa3s5E+I58DPZW23HwxCQ50fLjPChsoxOAdodeeHnlEZXhn98XmJf
DCTs/wuybSBtzav4Z2e2/LbWolztiQTi09Fr/CkW6AvJDuB3wJsoZ+JN+rcorC5acbok9yu32kmt
tzOQNU1uW18AnskSabmk+i0RFMi7RQhg8QCFAzFrE/cq+OpSE49DqtoLzQwdTheWKLV+W2hpt+cd
Eb19PqnwffrdYpRTdPV6qyc2yWAcqRsM3uWyzopHpV9e5Qpxyv80PZooh1sja3Vh5OamfOkgUPR+
Ng5G3fdK51OTyJhZXlx7V01y8p+S0gtKmtCp0FW4XvmnH6FNYAjPmMOmy2485fbYH6qGzeeiHrhf
p2zjoue9oe9v6TA4s4awe01Mua6GB/Yq/+DGlfMEyXXdWw3LTyER5W7T+36/R1HL/dnHssH1MMyD
MCKZlxuekB84p2KiCYn5EfkW/J9E5LN2/fQ/2ua6Oqg8U00cQJwbBfX5+NN3IEt/BZqFHOmy6HCh
LCRhSobwaHO7ujiT71I9h4o42H7BzeqYLVu1s4rtBfxmpdZdWWHhcAbtfA5pAFji1Go1Wv9Hf6DU
bWeKQChfViKoFjcM8weBfi42oNDtDCBieafOsVY1nKZBqKEeweN/wHykosqM/kQnOQEc3uhyFNTa
4WuZmR/LG+wl2LFWyjD505118V8gSl86dV8rCaLL504vWAIOLKc7L09pgvU6rSMPSmvm1zBTNfd7
iZGvTD3cmfC2YbE0qHVRvMT9bgU5ka2b3l4gnA49GuR2Wo67ct8P3XyX6TY7NfjVz0NhcyEp+tGk
lO/rTf6OR9wxF0Fx4FX+VvsrE5ToMq/jqqZpRBucnUT3Q31MU4d9yASM3iBSBDLLKHyxgraEVmC9
0XLmGfOPKssw5+3/Y2n2Wnnacj3bfUyT2j8JjUgUi+fzcNR+PKompZFhIsmGnhzU0JRls+2bugfM
X6eCzGvo2nBPtDnS/Er0+88QoH7iGPIhbqifUFXEW+R+WKZMYjqxYlx25D/cQuGP0HGQ2yoYWFHW
5jj8jAL+fGRcUkLs+AxqJZedM6Ak/b27vwwImm9WCpYVjzMPkYwECezf+xVJDe7miodQ/iZqBdSY
fwYWt0OmioVuKNlMrNsql5OtU1gnzl/aaol4JejyVbeBUF4/XF/MD1ydbI4yT1S4QLMBHs0BOFhM
ajfL9mQ/+NtQ9vHVMx71HKDBJIvXYE85iq0YkcV9LyM/mGHdWWLvJgIqIOEKLsVVMyErUs1tHigX
NOhpts2GevKQoo4JC3qn1RVk2rzvaH3AXF+iCbn4J8x2dQ5TgUEE4UhXqwS8Pg+uR6/0FnjLx6LT
VaLUW4z7NdN7S5KVCVDFLXsKicbrZxSJZMG3aYxvCw+mmtKmsPpR8ROQ1sCVSHVixpzlSteRoOXY
WY+gYuiexGHdgQVJuWjOx16hVgwP4tui5qgFQM5X13OG2vNQxqiN3UvR3CI+f05E9+491A1ZnoX+
wIZzTeRL6A7iQ+WcA7DVtnH+QFWkDZHUWYz0+yeFNCbxVYtOr1DgXp2Ku2M2/yJZLZK/UgCvABQZ
UHIasgHDjbBwcpwsP3xpi3hgQJoTjp2D623EY7sK7lBYYa8vF3pPoYCs70519ePcKvUxS803XNC/
Loa3ylMJD+3WBoJckHXadPvfCmz2Z2ePBJV/pPiKPAA4Ji44mtB8ut41RYH+ItepmIMpK1RwEuZg
2HpVVRnB1j3mU63ha3Sj/PSaSgDw1Nhb1+H4lqDoEDq5u/Ww/t1FBrY2SBBp1Hl/vJXSyLPaIj5Q
gSQp8W2MIxQKjlOT7PHzmFGo2sDBb3hVrKSifvIt0ceGB9nk9fVirXbJasGqFrA48MElOlDUKEVd
aTzH4qPXSnqRxINEE4/hcBppWqEERVq801Ek+ACxNwulRp1PphADwDw/F3zDTmFzPfhr5HjPhHEA
BVVKABmqc2l3o7ZSOxw/fdGCXH3AEeUg795buO7zarXei7lm9X/XdlLU828wycrMaZOyY+1FVnPi
y5ZV/T3AJU/Sv7JBlGGjoeXlMrOw2ASgVu3Mj2ijAV0n8KEJ3+rI2wUQg6qvFn5GcoVzf78k3jf1
xgFFSdA+GzUahBWof9vBxE9DInOM9RHHYa+nJh/GlHChbRezyZvov+gKh1AIZHfoSn9EnVn4BGGz
0e8tMHLwnioq5t4s4c1dl5d3aV/b9GcOdRxVu/zAvCk2P/6Gfe/E2kdFi9ymudSiGt4CprVHfGYw
k7x6C7feD7UL1VeD4MmyWYEWhfbPS5LFWfT2BvtBOHFsu6sXpQ2Zz6tQN0rZYQf8F2LjrakxChVI
3NrDeRalNGt5FJ+GHW72p4jH/o4wMSxpxFX4Lr1QykDagTO3Ai0uVfbsM4qk8Bnzpqrnkwkn9xx+
2+dXEUFsuayZThC2biCoKhldck+ypzRWuw09693YLbtxjtwWtKsqJoTL2KjiW4EMElZKl+8QVT8w
npcAyam+ieCYDzrWvBbi5AXlyAawwsixp7h0rooDjBWXwxpUEmqL2RgdNOTdBu6JpazeCAM6VPNi
qWJR3xSO4uWA96tOTF8JjSSsywh0+kWtwSD5UYwmFUwXGkwP69eTWcyZXYFEk74ft0Ml9k7eKsN9
ej3B5PD+ckxRfj1GoNQZBxDNJFHCtvDt6f7F2W2EY54ciLLBSs8AKNmMl5Z9dwf9tWmFB/3cDexl
6xnzEY+LKncmbTnX07Csx2YWaZGG0MoNjVxU9SjIRQjSO80f+VVuU5+mgjJpeHwNhuLm0OJs9n62
VmPz/R7Qsm2NPh9mSLKstS1J3G6R7JNk/Lwy2a9Eqc7Nlp97nqeDKeSSKGlv7qRFwK2q+fIfwIz4
qBfmO1cpY1kvotLqzKgSzkj6WUzSMQKtqFGqWMRGDpz4moUyP3eTGMXAPoz/1jBzFFfDpJMbWxoq
AonZKdWRpA34FiAbIR7P5QnoEYONLMqc4MwRFEWrMRYBdCc1bFTtvbLa2vtyf0b1ZsbigpxpFycJ
OaUKcV1IwSEkoGCCLrf8bXqWEi7aSfkJBK9SoZrKtGzH35VaMTIgs3lXucstYPs+/S82bAKy7+lT
hE3dFgL18OxOR05Y0bhQtFk3RPWQ2xvhiZgNQIKMEPWKt3PGrVGhYq6/xkdBMqHFgKXFON+7y4LA
E4fAqBRe9GH9ShQpSgO8VCkndAelZf6PqulIEynJaYnyoF9RdWUwRNzdy1LU8pFn0Qly24sigY78
xw5coI+oRHbKrcH1MAgsNWU1WkGiMiV9Yyj9pN8Ji/v2rlbjpegLLAcPOOxVqxj/J7s7bEI8F61I
F/wG5cK2qp4davcPMBjw4+adBvTVbTx+ExEyGF0HKW6RyknAU0q6VqZMWKgSgRYNCDhz6Yvbd/Bd
GH5W5Vs/apkLl/8J/5cLpIkbashE9U46Z+dn6DaJOSHiXdkqIz7lpQot4OvmWHYXiPQCmSQ9DraY
KX0CxgzrnPXmlFP3mIR7cboIWspJOynTm0KD/CF4HVQ8wJmE8ba8RVbE6NlNvxOFkkMF+ZmRVUmu
FRcdiJfDV1VL1iJAMRr9HHiFVw2LL81Lx8x7BcsyFW1TnZwIRNTs98gGdqJINjU6P05E49/lYYU5
5AyyKiNvm6TG7pqHM//gvJ76tYkTNIp/AZ8/0lL5agPVbmp0FsOtgukE4k2hMIWFitMeQxHG+/Nw
5nnl7xx3dxk4FAoKIGMyF8/ZK2noxLJ7LW0giA4xsm/QOmTiJKgqw1zG+VCRKw0aILiAPzNVS3RA
e4BKL7ky/CP5jzkjdw1ckaHgtdo+KCdcUtLhaagA61EOwWjvs0siG4ukij0LFOeV5cDk5QfQm/OX
aZK9H/FkULMNoYaN1Tn7sG+9XYOAT87nvKJ9zH9KJa4Lz0bGY8jKfS2c8QBf7wPICAT85SbUq3TZ
pK744awkab0KFjQrqLLh8/xMLYOVx67bR2+p9B2bthWHM3IBw/ac2rLO6tnr0gsRh29Bq+nsN6+X
iXcWqom3hXv3yeuun85SUm8CmtrcoTQor08E1/2UsYvKdGjTRJTwjUt8s7PH/sn6SoRLFnSEoYbn
yMDhAO9IhF0M8u2Rd61iHEUnG//EklQjeTltIhOd6keEmYQgbgUoZEkW6wsP2eycBjrlogTROrFI
ba6bW6n+c6P+MDxEYmh25YU3bYWSvwFwWnoJ49VD91ttVuVZyQrPNQ81HNOZBGHUd14lBHhZP3M+
UoYK5KQtDuuIYfQGbqAQiFKqupxosx4EUjsKh+fTURSACAU+pPiRBOWyueixdfC6h2/6RED8n8/+
KIQBDWK0SZY6xNZuKemFf60HlWHoaFBwNTFeiqx3hXgPc4HZTJjefCJOw2Mb4Sl6JcC+A7DgNfK9
IbIMXEy3baabpPHu2t9gwqu0HSA6bxzfhlGG3O+5eLrRhM5bjAPpTkVKihUEmWF/i07gp9Q96Td1
pXTNtO1SamS6JKXE6P5FXw4AL2SDa20V8dCPEjg6C/hHXq5uZSLMuWqn81Hr7DQf4OVKEIrM7wtc
yyEeqDFXBd+POtL7MOwPGwkTISrNNukVXNAD+b5/qSD6EsnbcriH5DqS9wZQBqQvhMulTrk5/Ueu
zzQ694z1qBTOEqqQPufPZClNwUh+aoFse6DfG1nvxaufefFI3znYSq3l+blYr/EvyPDKyOcfkKJI
f4VcfMdeFEOf3diAaMY8jqwza6cB3sfX7Ko+QRH8YBJeoMZeb3mz2tfh4fsVDhePQ+s1OohTGdRt
+Kou905o5Y0N2SiiWVWMgREqJoZXixBjKnMx3i9yv9DbizEZza1myJ3J7E4WPxSavl/JA1+xGHIY
JTi2R23tCacd/H3FWunyZZ9yE4fGnXcDJApYe6XBo8MKqxuSVw+phyR1Mw3+zko57Zh4wFXfRhRJ
Htvt0SAnT88JEwFw9DdD/ANuK0ryJdznpSwd7Ijp+1CTCkL+gXZGSG5AroyFBXa5tiss9D3T4Yhm
q1Bz04/QoYDyAWhxXTVWUot4bYvZV11DQxcZz0uASuMNsWAGDA6SxEs3N9rRGsRkTn4uXI4rI7Jk
tcDBJlEdYxYL/IL/yNpQswbF2bHDOwza1QVQ3cizmNU18xbpwwok8LqFB8boBPjkiRHj/LRYmIHm
9LGzGDV3xiITKU6cT4iPDxt15yS5V3GEislIqQ8PYxqgFChko+XgMFqA7XU237uC9oJgYijEavaz
cP+9ng131GT5lZOjdBVo76rdWbTp1eQEkO8J7o5XQwnXM6UTWw/dbb5L07rZf3aZUR6J0leHJ+fu
U7fFYntaRQE74bWFeKEvWsBw74KDw4UYFNqpSLGZfa8DQ7MHByRhy0jPMjDmUzZvIhQ4SoTfYfvg
V82aVQRHZJIxVuhK6cxWqM0p14jFKZVuf4YmeFybZHSgUOD/AEeq4IPIA6Lgge0cM62s11ihcA3x
SU9kXKM8wIsPZqUbBgMj/sZt4OEI361U8NbaNp9dfeXTxbDW8N4vlvbGp1dj2o/PJPl4Z3zk+YIa
k50qUBaCVCVRbtRQ2pLc1Lajt4/SamqyjagnbqRwOnVm/jfTZJuqRasx1q8qAj+3y4adJBK4DdpD
wOooMwd8nmFE5v58afmfIMZc1/m5CaGjtKAeIH+TJEh8riGirvYMxm4EdRCTUmWsjzoo4IPOYFME
BUPg92CrOB27WncNDbmmPx/Rlr2pYUwDYW2jxI2WH64EAxr/AVWBz0SXZECWq9Hj8LviZwfZKSX6
J1YpGEEH8ecgu2d/R752Jr7JRMibIIyJLylwS+mPowK8MdXuH1L3J9qqYMoLCNBWqGpCzS6eLvEs
v7PTYxSL+AvyCCSispdQ70VaP6CakQ0nlRt2NtD7xBeBBoqHbfGDrYvX/m0MfE2amvFOHErbLfdl
5vSDAh5xRYuRoaVasDBIRfOjkJWfD1u8m5KpYJNPIi91fedb4bKJ/vEaBz+vX+Y5a+2e7s/bD34p
/jEcNYctCCafJLRBU84vxREGvG9Gd7Cv2l4hWqF0SNXcd+hhZ5d+op8Rwh/rJqMIFCu0NPr54COG
nRAznwsIQX3yn8gIstR9/DDsX71uLFHffV7lQYt9BDirJKfBWDjMqIRM5HPXmAbQKzlQvl3e3C2D
q4fZ1CPHt7AR62Pi7c70S7diSkoicZrsyaylcKwipNLRfMFwRnqWqtlzgkBa7kV4BSWo2jwTFy1X
jJRKSK7a3vtZfL1vPk69Qdk70cBUL1fj9biz9jQ8vi3cDbs1gdxTwcSheuBlHBRpArN/MuFmAq0g
emig2BZqiXaHwg9rURvL4rpkseIkcof3TonPR2Iq8mXEvNrsXAbBvb09wSfzTQXQYli1noB+ZOKe
Mlu83PWABjgtK40+KF7msGwvJxhfLbbESpAoFsGuJCnfOiWkpGqSGkkLkyg6vQ4XqBBM22Vm5m65
zS4DtbTPTYNOD6jxso7aU9uHH6WROcf9jqTFbKkV6lew/DKxP3hPXwb4x3wFVnCxfEPtlCKt+TvR
Q2QQcZIRrJsWscv2lhsrxvPlf7vB1PfM4h8FZTS7R96JM8azvIMQgIOCpKG+bzI4mu9Ex3d76koq
iaa1BKPHaXS0OygGlXq7/59JnvTkRBqo+UtPRft038Ilqe+QuSFfilEqQSs2sBMTuli8ZPKXweUh
ImtLO9A9O4KmpXjIUJLp4NE3Wl5iS3zUjMjC6xL6nupaQ4wVtDSeeoPUczcm87YVVTf+5d02eRFZ
Oxwc6CWITPXA8IWN3lU8dcRYPwgOqiaDsPO5gUS0W3ZVa3KeJ8Ya7BuaBuASsPx5E4tiajcxPRZM
Siq0nPFra8WtRtkPueqeRJM/L4nG9/uGghnESxkpCugrSQmMiBTn6Qz8c6UHPqGcuNGKz1/X1zDm
H7HrMgVG2z9CLVk5Z8s/MCrV+RLyEITjkKryf70dzy2ir8HYvHfvaYA6oJJj1NtsaB4Vh08ycHXf
C9K1j3qGsLa1x0xeQ/zB+MlWyv5A9215esxRX2jpIvshqqUHndQKocOLgHx5iqv+UIdV0Mo2lQb2
uWTz6MQrvOSPC70jeSltZaxriljwxlriItA4j7nTXEzLz2QEwV00OOMi8gCPoNwFPsofZ3MmfI1m
PNjl9IGLumGG4vAa+cAAGmP865dBSKjLf3ojTZh6DnkNr8tql8kudbmwEW072EC/DkuCRtU+vV7l
DUXYBLaxPRuxHumBpWm2OiAR3WCzCE1e2WBhBxQKu6dl87o6GX/kK8YuiXwATUKsU3WVTiZtKC1Q
lBq5DK5cf0cJQrs//0Ln1/nAfxsYzruxTjKrG4iGmmTsA1bzR7JB8ohFclioUuufEXJoIhVR2nv8
H1U6SoI9he6cPU4QReGTO+rGrOHxbdpt8sDJ9osdJiUDQpKCuDwudKJqBJ1GT/ry42mdNj3UkLH4
NrmvH5FGoxIgOEwzy4m0AiwRMRVuX7kdvIVyNWhbVu1rgbZSgmEFuE7w9AsQ9EfnB1UTgMQJRK/W
ftN+Bsrp+MMAphq6dXar00EWLU8mMNjcQrbboy+NSx60c4ZXqMuM6bhj/eh78NBAkRFyL0xwyRGz
gsjVTYbfYv9hyQ3z8thEq/lRWuZ/ReCJiIaF9SjQXtW+j/tugZ9cOIfNBzvDRDGJF2D4P3a9yT/d
f20c/qrv/YiwBai7smZehMuCV/c5GxpyqjbzUWffGJ0xFsklNGiUkf1JmfphTekWXYskub+18YQ/
wtpCPb2j4C6Q9cCelB/YeIgOr5vgSSNLwBEnmsEYd0eY12Bz7Dss29orgbc3HpGJDqp4wnG/D+eT
kBfJvgPHlXHeEzJ6B8pF0vPZAcHMGvPSlqrApanhgQTsKwBxkL1NGDqCUw+ABzbKv9ci9xX8f0tL
bUaC4eJHRSgY2f2B8BqI6FqX1MeOki4H3rDNYQ9uPobeZaoHGqDeU4+LL1nihwqoi3YbmrmUAIsK
No3gpAYl8pYAyQq9kyDw2JZvJKZyCzk7IN7AJlLZeFrXs1KUldcGVL3YQAeHQuIYSy2tnLUgjvP0
5WIdSvvYX+PoN+dUZHU8j7mLmGYEWJ1ACUYCPZarVyiFe9AGHWRCqo8BIm+cB0SHMBGx1zti0tu1
8TiFXb/juhPB09r2DTzW+Y+JEhi/dEXtCxLuI3bCUMnendr/neNeIMTP6WJgVnEVX3GH/3M0WqrB
FjvDLIzu4D8e3vREIDoDPXzqLOhhjJZCRNzmZKoyTR8B6JekSkqHfW5fi9xDE4Bdcxcbs9BNifoz
n8K6mKBWjTrssUpL1GMQXnSpfzw7l8bHtpUkuPUJYvF4KjcDsfXX1uaBiXrOMWJxnTYbiuqslVt5
n0PqEEg96IjN7pPXtbnCanGENVLfKWzKzmSD0+WiIrAj2vw5kGcEFL+Gryo+GnzWGtD8H63hb8x9
O3PTF9PrRudUxu4cyWT20GoUGvUz3AVwTNVNzmSijlrFe9FtCJqMwwR32Q6b6tb1aB17w/9vNAlj
athfh09wTTSEW131h2aaoDiIO8SlnGcJ5Nwx98ght5FU47ivHVQYHP9kWXWxAe1lJGY9wq/4ssC9
a6DiAOXb+9SI7dr+tt3XapFvuB0sy3GsLqkL4ThCmZgrTFBfavK1uooP/bFsGDhpAcLLRorJJc/k
9YfT0whT4doOZ7WGTDDID5oKr0jXrZAsO2CoqCPmN4A4U9gOBN9goblFb96VAyfq9qMcsXlSfJql
Vmbr5rLs7gjvT4fBJ5/OtrbDFR6CplaJhFMUKawcdDG4umS2OOUU6a1vwKWXV58eMBOmClI96ykC
bfKMaBr3Yh3Z6KENi4YbiSsLU+pyMYEib/MDEdrC08nqFr6UmNcBllEqWxEpQPue8L8S6MyeiiT7
QMXQlHJX9hw4sQoXvTU7JrsaGJ8MKjOekSlkxQ10ShIj9Ivnt4e8z9n6rW6VIngqI1eBxeK9s/e2
RonPkJss23ULpbOEp+FKnYHXnnyvdl0m7Z/DZqEWQDPZFhI2llQxOnwNsiKZ5zSrb7QFy7iLBcyp
Vw73yevl6PLGnOXH+9vEoJFBE8lQ2aepkZUIaNBAffejFoPyBGm98Yr7Ak2mQ8brNeJcHknz8xS0
rbHW8D/ejggavYk1UH7WBPzuQBqZM1lQuhhp6kEJMLJf8XbX7f0Wi0XNZSrK7CgrYUpiLdQ4NuOd
GkBVaedQU7V+jRehbff/r1PtxJBd7az/KG/BkvTGL6/+400YXEuYO4PM5WpDcjQhT/ntN0C4RHCf
mbrIIVxMuctKiEV9i+vAoa44KAFfnRRpIXsNibijuqMwFJkhRgTb1vpuU+9Xgb+yTaAyyqir5q6r
IUwopyryykEet1bKb+QWEMLDtQ6u3CTwVuP5l0aZwxmifAeU2xrNxnummoWf9qmK42ASV9MJ2wHA
sIzKII6LwCxRPw9D2+1NKRntliiysi2C4priCTfcZ7l2wZifYAsEDUzwi0n7I1mG09I57K8PB0xt
KwCOVkys/7wCC51fshoUiy2Oa7XLgusvu1HqERyqvINDSsdQf+o+cSj1S/q191nqREvmU19+dfz5
nGeYP+alOWnYgCTDtOHpIixRVxIR/EMtef+GIQPQUNK4WXZqe/3Dbed+Nuel8J6no+N89Zbqdpo8
y57mW2/Z5mv8VyXcVyMtn3sG1dSFoVwJ6Gq8L5EGNFfoc6kNljKrmO98VUuUeLCWIqWCmhqq8fjn
OXr/cByBxruf16XvAttOjDinyRCjwarocPCLda1nUndu8d0pX+7sCj1i4OBKnx3K5fu5ascoZKkT
Ufc3x4rKAY1LitafCZfgoS0IaOgnDrYfJznYniQ0VsWsNibm1VkkRmyLzUdRQOQtIAqRkSv0A84P
gGS6RrlPBHsy1HzojqPURD+ogKqnHW7fhFPPDMnfqPfAGBEuKMSt6WFbTqB887gtHStbERXxAt63
LS3T3JU9v8ZfJ4AjKds5K6O2E76YvFgU3dGWGgOA9oXmSH9RrMUVz6BVyjuc+34o06qVNMEN77VH
/KLfXTE2a9xNKyOcmE0w67ZJbHh0BVQHZ8LtTYXOvGZjeUG82RqT4s7rBVvwHTfusFdPZnNh+HJB
USz4hZB2to1qtSdTzrUXOrew8AgcYaRvZr86dzjzi/ny87mibVJzdfOVnAvWZkZ2DzWqfyoyE8bT
WCQMsosKP8tSRtgsIGZLFXvra6lOcyUAGtbHJRhO2wU7GZ/XdH8gDc1/6SBcQ6nbj02vCJRc+pmX
whrbRnRw0pzT8gMoRfDSD0YsDgt2l3vwm+jGI9wDIzB1M6N+XmOR8ZvhrmGKfHvKgDeDmxo/+lUb
2+MLk8ubDjKzKm/aPcAYaqUFnl2uv+31hcWu05sfcERAEnd2gMA2xaCUG3+7oToA2pdFbcqF/acv
7fjIkQReQJ2C2eE330bN0Ed2Ebz/7j4PB1SorICSCu1iEpWugKfIhmxGh2Qza+KgpYNEqPyEEyyC
QhTqaww/GHhMvrOllFb6oQkjB7xniZw83UWukyhLasKNtB9NV0g1/YlaFukNNZRPFjMkTh5LZgP0
acEvQUNYDpFfgG7OmxOAswPe8vI2vMWfWM4hGwbeXGyAMz8FFoZQFhYn/FU3qOlTVe/3PSPg/L+c
E1eWNM5mcYAEmhgH8XzRf7VySxS8oRWQgeyFEMDDC9jZWEW+SoNZ0D9/UKM55JhoEW0FHxRV0C0I
dv6P+50KHsSE/j+MSiYQ5kq37Z34Zhc2a9h1/W5gL5/w0IVLwbwt2yBeBn3qQ+YCegGCb6J5Ovlh
/GVkzPxaGsy5xXwDexo2QgXC7wELxxZud3QUGiVl4TzdlWjeFzZIUEVttd6iZIDGih1vpRGLmndJ
Bg+kWTt200U9h20tWN6NPoXpJoPztvNDiHK4Sdo8HUG8AfFgq5W8HfwMLcpcupGj8Me8+8Cy11hV
xwU1AMCrijqpm5siR6d7Ve71dVMN1r4h6JjGdnQvqxnQBBVlsxOwSK+aWa3naQVwzjDBluBk28wi
brpkMUeJ4hwMKYGL/jOWkbt9N2XFmp2UdP++2cAU4HLkl1l4+iMIsFWhZ1lz7WCUW5+MbGVy8Piv
W5I8sstp8z8H4RjJ0kiGl0IuEGSnGcUPfjDaulOxpCGk+bIpsXTCMmMbs6IzIiSu/1KO/zk2yYzP
J3RiKPma/gkgNCSXW9+PGVBRSiUZySVyGNfQSTl1gy3dqxEMm6FHF1UBu5Dt/mSZt3UKF5JQvFHw
GjzDeJeDxYeMKiXQ6657IXz90PISHLnUvJs64W1H9SKMMD/oxwx7oFWOBD/fpck/Juml5mxIupCi
va5DYJI4oblXRcK6PbFeauCnPnhQPciXAnkiyMnWNnEZtOvI5RI+25RWc6Mzqc7FTUzayAuZDdLh
nB0UOE1QwwoFoN/kKbjKV/0GWtwFtgVsmU23EJ/YNDq28UZKHg0XBq+L3NFMsAZ7W0gpgcE99kTy
/u1Q6foRURYDHY7o5UwgaqsvEAdY5d7fFiGkN4zXIWLld/nutPtc07JEvkoryUpgGQuGQCjexVl9
llo05pRlBX/j51ANVQy61YO/HG24UarnGksYb/NPkf9g/bSl11acRqY323UNfs6rPb+J0dt2cA46
HoldR6pIv4Nsak1/v/BwUWhkn10mLR0TjihOdaS05aqW3Ygbd/UVSQNqiIKsEz19RJQ/KCK7tnqT
qJ+R83gan9G3TugN6nPk0hDiwuV0GBeBV9VM0VzErzsUlu1FNFt1zwz6v1aDqyhCljwqr7kx6Uyx
U7RYuvCFtixCqk/waOLvx47ILN+80OdD7G7LEvR1dW57cGeSJJoVBblzBF8Gn5JrLhYy1PfUj1oI
F3gWJBOvwM8MwfsWwg9RwkWiok0I2Gx2Kyn7RIg/8fZIMgGLjaxh/fk0SdMmyqnTkbBaWosoOk0I
szzBXJe4cHxtcN1CYnPCLRxf9sKwzVf7NJyt5wFOzOMFllQ3p6ySxGvpffoQnToGnlGJ8OQBhUg2
zEhEu6csNbtsgbb0OjYqS//UQLCn8vqmMpY2NTZz0neg5zTw415Q/700jBr6K9x8in6s8YXAFBWi
7dbOcVM4B5FaRdInBbjXXo2UdnOxgKqGoczZZIE7/CUwuzHqTPTJTggJ4I3XT5BiyA5Dt1cUMxHj
txTCoZR3kvejykUeJkwWBh1B35bIt8DezhUAZeGw0YjtAlIhI1z59K9KPR5WiRj88xbmAI2VCa9I
19ESqVwAl1bZwDDy1Q9Ld7Bn2WikiVsgz3kUqCsKSElJS6USVM7XkhU9GJhP+prsZkx8EbzXVZuN
TwFpeifloSmX28dKf+jNpKnMKCAs5WriiDbZu5yi0RhJSrHHJog3DzdGpk650gA/U6gZo81YVdER
J2P8/R7x72UUYBSrhFpYVKaQ/my+xzxD6XIfidMte4mn1C6I0lG94u1/6kkt9DX8ohbD3S86wIIN
RxcHTGMn+Q6jXJ1X0CpkIMPI3e9fNNT2Rc+9qXyXIEhnyWeD3VaVnOH63TAfrPcAPq5ObPhJdlrO
hdI8l1gwRKK+dxrIZ96ko4VKnK52zXSZy2Cbp4R1irbOuGAOYV6we7qDlCkP5clDWznTPSROC0vH
VtKnszMyzYencTTq7ok2ajhiac7M1abEE92f5acDWFZIuPd9AZ91RTIt5leEWMz+orCfGbj/qtD1
ON5N/GtVJLm6hAHRWs+IY3W3rXYFafqzDnIP6o/M+Gb+leYyfV6cscE9GHR2k9+Wen8yL8m8rE16
jYz6tPpdZeblHyjLKtlqgqe8jVnI+dx+b25SGuSKyTID0/KZPtIwofVi6FHxqaj+ZLOtM++UKAAN
NSNa0c0aDJ/FKR/KcN2SC7oz+g3VB7LRkbgb3Z4zpzOAlW5+1GAtrF8MCkhuD+cIRvCtvXsgwsca
BQha6k4f0Hnp2A8iJKlYjN738thfsJQJqycPHUe0OqrFRr3ukWBJYNGTvFxcXMX4jGIKiIMJv9em
N1qpEWvoDgAf7wjGFZ/YLPeMaQt0h8eY0t20IKlLG4uTDaqJcmOm4p/GjRJ722iCC5C2cik0Tdhz
FdH3Jw0oJQijANRPAIYZcLqngRWKkLVDJl06Y60mYyw/FtwJbRjUqYkr/CNdq/Xn82SJy7OQdQgy
vLUSqx/isXQyM3BBzNYiPZ6FO1cl8/zcKO39n27vs1SwCLa0/rfArc5V+f1C6HGU3f1LbZXNKTo+
iPwjyd9EVPrtM/xWrV1ECIrVhJLcrYeBhzGVXyaaNhOq8Y1w1pIx5Gv+Jxs3eYP7m4AaKZO2UgQw
K2YA76Y2BfZnp3ojVqMpHsFg0GvMk+Rw4V2RYtew3QnK0fJ3X8IioYkuzyN4VzCnWE8OKlYV9NVC
DmT4uAdlIpt9okBiJhShaSfcDkVyirYYnHOo3xakCjeIO6VkQuEiB49kua+NeWnXO3yfeMnMEewZ
GjOFj8FWxRF78ejXIwdX7bDmay5hNj6CPLavVxHB8dY9UN6mGxjUmn++ire5ldcW0yLFQnUOmkRH
NkoJdJrrURHWHuIG5jKKe2g1SVdV+x37RgOJkwmNbhb7kQhT2q+kCvqjYYAUGJWfDLWOEtyULAXv
usbADhTixdkQKbiuZN2dWShMVK9dNVkqr0tJd1WyChqe+GA18KIHoJpyPwyZu77t/U1ZmteS85XD
XQByYqgBCi/qbVWrOxA1n+WtbwuHvxBOIHsLUW7GgQpRn1joOyC6kovcg7wqK3srROEZHItOg1Z8
T8DyQR4WVCsCdJoxZoOEc9ugWHb72pvufkUFwm/K+TLXyiisTDahQgY/6HT/ObTjr7hIC48HhZ3t
wHh6AbxUgZMQ8Bcm2hpkJzCkb2ouiHyB8/SPlNUwiz6cXV9V+spmkwuWMAPCzyJvbsqKmdRKVfwi
tcmH6wcctyq0hWsxHQRYzNx96a82PQp8awlnIiOZrSQedrbJCY/ItG66QdojHPE6qDfB6AVmVMZP
u0GKvIzA8bNqb1/hSD/bTY9859tlGCiIcdxjMNrdgvYhfDMTz29DMnfZ3ij/2PXK11K4GvuvoDFG
DNn8sJiZeCl+KMDzejrjiX0waju70O1FmK7tLLWk66E8hC2nwONUr5HOo/rcZkfxfSZjM3lZtmhH
5YW5XP2QBxwnggplboj0S2ZvZxDtiGNmqr9wZ6UU1+YzM2kEeag/ZMFnn0qubfe3GouqHL09RV39
HoUME1Zf+DVAsmKD5JYeOuv3KBT0n82U9ePoUaR66WK9m34mWJvaGmq/3JoOvW6JpQD5NhGcahAE
VP/F12fOri/3AMRw8GAjuKneqwsNeC+ObkSgrQQK9C56dAsjEdNSRTlPYUeneKkrp9dTmo/7DMXw
lBCwCghimijYceSGW6jDUS8TxVcuYpoki9un0ECaWYaGlKoJhlk2wzc4HrNhX+sR/tw7Oy+lTth/
xpr54RAxrWFRqW4gN/4g5k3/nrftBx1K2JhaaQn3cKtZpbXvjzQLaklcVKwt7rbHa6XA1wF2Oi+v
t1jknbTPUO4Lbh2RywQ1W6XKOx+C3T5U+ISznsTPELwIMUSz9Wh3PJEC5F6rsDIKnJ9B/gaQv1sW
GhTiwOLQIg4/HhiQG6iCGXYSrs2ugQQHyEu20N/nG1Uxs++nC4ulC0kG42FD88+Mn4nfrJb0jQxR
quVt7dvqEOIek4YWRSa3yw1AbIy9QUuNyCmCH2nWVZ6/8IS0ryi2KdaPf47F2ZlouzZvNPjTkY75
RYbYvehH8J5vUZxGXU5QSjM8+fAodwpmJDfvLgwEexVi+r5frmKbsklWKqp5Ppx+XA9NkekX9wZr
EdaUqx133Mfbzm2IYt4NpFsu2O0NaqvcMAxMvd4P3sMgCqAtE0zjlW8kUPfZmwJdAykFaR0Lepk/
rKDA2k4tRVjtl2bf5rKt0+DrbuI0oJhAyH8byaHG1coZckNjiQceKnNy9TXf9hfJuqqUI/dTYdJ4
9FiDkCe1JWJvu4wsmyeDNxnmLBTLp8mSRsGK93hA12+IWi4O4b750dedHmVjE+Kq7+/omtbS8mnd
BsZc1u0NhmTY8jgHut5hQCXCxDHNNb62o5z6FOQbgm5ZibekfVhgO0XFSkjQM6IVSqSSgagMihAt
RQXlqfQ5owvmIORhm2AhHuXlHtpXIUjpBVTr0TU1tNhNlaCF4zFi+705DqIKJ6czYd/Cv28bLZCB
inAIZGGiwlOs/blmhgE6IbztFvWp+njNIKqAgruO/kdwYecT6d9ksvfm1MfkCVQ5vps7RtX7HxgG
XZ+WaWPi4wVV54tdru0NNvsOu8eQmQSFxw0w1G/Wea+xFYeQJ26DWzVGPw+91mo5cEL96582DseW
Tdl+/xXVkY07LWMPeq6oa19JdVrwTttYFz1D0iN3hqKgcPIbfkqQHaNVhoipcoNQSPsQ6W9I+ICx
mCRpetCDd3/bzGMP5FD85C0VWE//x3loe1RkcVmPU68fhH5U48gtHedxUaqElUoiX7pw6JEQkDyo
qFdyMF/Zo/Ze7/cX2DenXiLXEKEs2rc9FsV+8AqKqMWYLm8DpMC4HvTilZytlJrhQqef4ho0rF+P
xFj0zeJwzHILjxYZj+U1eyWLkHyAMwXAbeLWOyQHif/uEvSPaQshv2N2SduXa7aepnAinU6buO/9
zKSt6+ZjfuYZZsTlVZHKU8/5HiFkCjcAKD1rs7kBd+2Tqq0ZUR9tdhlCtJfMOQxBtjp1J8jDgJjx
QzFCn+IpUoKhqjDQeaKtIzD5nbKJsVor4yqyzB8HF2OSeFF1+z/uxBDektBFJiOlZkY0diLt09TG
oWPdsWsvugcHGkUKsEc3BU7UAYh0lMIw098WTdMtrCyvNPrx4Me1Ik49fe4WUjhichEL4MESdpwt
rc5SKAhEgtQK2CWvsGwHrrOt2JtbzWpzPdrQICd2u0/Gzx1t6dYfwmlhacqLzgFcpUnmmQEHBeeM
OB1zQjel6mgibCn2XCukczwn6EmlJyftESW72qVD2Lgsr6pCx+X04KaOEoOopciyrhPN1CAH2ApF
R0rMLX9iEgpgkCscXmsK8IF7rLxz/MNEzFVTXDGqF9ILcF3rvXuU6vjgFcONq1HWuPzmA9qScYg3
1AWAzUIZ4lIQija8G5qkeg2g9qeDSgb4NfatfeKeNfCpK1c7dzplZMoKEjtEQLmLKyzEawlRKuxV
4km9CnVL9sPEzNIymX3IA23Vop9t3hp5JWUlbCGMkR91lJGJLW/Uo84xxAPq8WYX9c8CBI/DhfRc
Hg7B5O56sYj73BSWIkMHdU2Jhxso9fbYr2fah9gpHIgKsXH7Yx3zmBXTF1RIno7xdrFxM5AXxxDy
J/crRDSmbGs2D3/IMEYCq8fW7/H0fhepv3GpgJfzMOBh0eAbvy9sHScyXc1ZUnvInEZKvsQZX6/+
S0qNl/QgvQ2ZDrhkm1Uh+ryC1rJGKoeyDlUAsyBckrGkeGIqS5g7eyrEU0oHsnGPO6iRZ/ZYsqPe
KN4kGID8Qw8RKt5U9UhGH5f6Wh3K4232UFBLaaXoDVf5Pn4nl0DlTz6M5NXMYj0UGYjfgA/VpG9y
R8HqogIUY3YaCGrJlx9vmBEF7VC1RM1e6masnKSuR0HCo8EateFiaOYBQmhckiqgONKSQ1C/qXo0
S1e4GU+0R3wpt8pmz1BM67VSTz01KfMScUM8miznkc7gFPGJa1jUbrvJDYWPFGSF6Jk1/Eksd94S
RNfFytPTzMUSP9yLVAONQtZELF/58Dj4+mWm6mB2C/SI1ztwlm0/A3svJWmp+qEMDSDq8acK7hGs
lnhKWS6WSYS+T3wki/AXCvgWGHSQ2CDyCm1HLuZMWjEf8xPH6dKDBor90A611h37+PoIJx1cfQf9
Ih1Kj+cINUcQTfsLbfkTC4wlY6VV1tY1iWZiYDPh+qOIIOp1MEptozhMFZtGauSiFPsj2mZvC/D7
uXzJbFGxVZ5AYkz0Klnwab/XnLxiUHVjLQo7QDBRv9zTOfaDHjgBzBbDUfZValMknLzSvflYPlkE
ponbDVKKfWdH9DdPmyHbcxj6Xdy9+zy0/O/EybZaKgDSk4glH7KP/D+45H0hPgywmPtMOWX7FAXP
i1u1anwmCgm8WjciuWKBmvxcgVQVff9ZfCb7Bjjv90YDONcNtX7G+qgZwb2WLVylOAdfzh4WTHNd
7+YjwNmkIVX4DedytWqwfL6SFl5miZqRrnqNAP56yfJThvuhbpNJs9zlCgPlwbVDjg/P/+t0yUyG
lju/6mw/KDVD26LjhyXkhYj0Lh4d5V3BxHkXCW6SaJaNqdwh/ZxXmzRRod3RiK2pdG67JzxYrvQA
DC3HxfQKN+MDo2HGouZRAMP9Av4UJq3VYsKlkrThHynrVOFtHf+anJNDo8+Y2eUs89x6gzPYfrEQ
JRGRBg++F3W922sjNb172QMrasAjDV16Tvog2u/0jwsKQGkcTD7l1+4nXYgGA+SnVfMNW9rZvPkB
kMWq4elbhont0BMK/Du6eeEYZMNKYrH1pnntqW7HLhGz9iJYnWY8FSaKOrcjz5XyXJ6QweBdDHd9
51b0viyffQbZyNyNE5NoooGxhGLCV3s8HrwmGCUzech1kurXMyWMBTnjIcmZFWMXoUz9o2siLD+B
o6E7o1ACRc9/NYNqwPrfXTHBMD8eIco9o9lAuH6cOaTkn336TSo5VKOXYr+laPytmQ4QpPPShmT0
8hkoMo66h8pOJobH6dD63OyNu8NvNnXG6o7tI4817fR5mUjY8gL5BVOd1Q4StVSlrLRCAsxgMmlS
u6WtisPeZzRKdp1bs+qIDvhWXcjJtbpiiv7euBRPGkPKa1jO4pTaqISam9c3PP5q4ScdZ4EE5D4x
U0AJWNtuen3pRcLvm0QU/EW/pEg3CdLaFb1SLycR1DXkOnNd2PVubIc4xXKvJeRXLn44sV8NjJMl
67yZKtlvaU7lMHqvkHCk3aH1D0q87iZBeT5mtx9V5nLiZf2LMPus19+xFfNn/b3SFE+H46SZGvE7
zMmM28ln0WtXdOJjif0b0z8IwRAsTG/fC8x6iEqmOtdWoxnuPqJEbZOOXcPW37LE42ZfYhg2+9q5
UgLdoh46Ehf0oMTRNNxR43XwpfRfRNcmgUlWP5zLkI9GPKfMUoKuozHUMIcxKDja1wfyf19kyDDp
QQhKXVB6YLOIerLB5EfGQs7It3uDJ+AbDN5S3wat4cchzK1y9I4ynxTIlotkx91VTTA9gCtxrqlo
KxSmcSNrCjckd0p9QbuFtSZP9WYiV/RVPsKcgQxiw91gH7OcBwNCobughOp07s/2LBSRXvO3UeKo
9k0rkG1v3CmtnpyLl6NIkrGeIUySVqHfAUR/aeY20LunFpRWAa8OZWdMcKedt81hj7K5ezh/3vsh
RjyWbB/pXrtNxf4MFM5zPlCKe3olKjOQBNHWwOOmm0I3BMAU5vdoFo+RANfGD0SEh8XtrHrTTfcc
uWQ3af32Um7VsTn3bMfdLsnoeHuwpDWxIe7yLAnM4SqKm9AaiYQJSmh7v+YgZrdzFGCTPA8lgxBo
xNCYbsNoezyRtUte+M3C9jE//XMNeVa46saeMlk34ejtDQjJxBeudlxHPkhqHbAWPNDYmeGmw8/X
p24dVLFpGHJvtFv0TWQZu+6Clfuvzbf1EExR1FyfFDDswx7gWVk15TOkN/REHHJuLxM4fi8YLUtf
zoBvET7y28hvaHgznLnkN95UEXcdQUEEEqjDON/1a4XLpAknXGjGVtXUsroZVDLc6xFnyxKESF7u
W80lPNHfs1W+cgx2MCHmYq6RzzBda0NsUQ+P6/m7vkWasCiXC8A3/DxjzlAw7A1PU5z+CVyvUjY9
QsA+AZxcqrLjB5c2lRuqNaXJOyIzSHz67+LFCE1XgRv5MXdRckNTVJ3r/3MjnX620l+tsdDYeod8
NU03Llgr3gdFBKON7UcqRc6VJ6MotYL08HEniaFmA/xK3MCtTNoBhw+27nuppQdRwtwqEys9JUY3
kO5m4nKC8w7impAjwT0Yf9FDMpI8T9tMW9TUorZIePBtEM/cXJ0aKBl4E39DKASXv0WS/cmHoxPl
A3bNIfCXLLhMM7KPJPkfw39DrlSY7VDX+/CORJhZwvzCv9CIkFnK4Hs1g9PdfpmV68AN0bcnxhwD
ss+T+UKVa4vZahE7Zjykcsrfw4R6V7D5Qm9ZOb8D7NIKsGRD4qu9S5DaVnv7xXAbeNqt3VQPBs8W
KwIz98WXqFsuddFtNyg/DtKL5YJPWN4w9bIOcKnQz7OXltKsy53Lf4xY9vI4G+/Oo/otxwXlEJGL
Hsyf5qN0FpQNIBqUp6IgtScaJBvbVUFzje8g672BcN0BP8UI5lbBxbWqsGFoMA4eoa4WodaA8eRi
sWFVHy4JU3DY9dPyKsprGn9xdCzCr+jRsYSKSpsic4u2LvXiCGR58q6Tp7b2S+0PAkYuwUdpg0Tb
mBstifbPmqn0GgEQjBDsdAw/WPCsuBg9Y0YEWiAtujzlVAe58u+rup2q3XXyHIUkAMdlQK9YxtIN
FIQIaRYz/wu+tTgdtfpWGKIItuL+Fn/YGqwE1N79acjeR1Dm6yl7nQSjQ2RlsoO5PX0uzFM71usA
xfRZBkJzUgnYa7rsJZmFCHQH1MarNKvYeBGH8KNYDOl8Cvs+BxVqUQKLwIBpewRGKOCianotsXc/
hBZIKxpeV3gBr9HJ0Q8uY4G8VfLPK4Vhe2khs1UYccRJmloiQotwgS7F6LFunaRanupFg2SUpM+3
VXjSfuXJ3Qcgt5xY45SSjq+TsE40LvkYp45dg0GWVV/UfLCxHoJuKJ1SfhW2TwZfsVT9Oxm3Rpge
R/Kqe+bW5PbzkM8tDV7zGdmETeaE436lB75Z8dahYCKcpPgDO9+eqzV0il4teU9AsdWiEGt0R2rQ
yKXZBCi7AwjlTwsnt4Mdwt8Cmb1oqWlbgTxdg8fKHoBn83jYdSfm2JQwZvyVauvoOsEbURU2INIE
JDe21xNZLnCLa4h39h7PVOgFhE4tnzmrXCarx2UOoj5y3zU1RI+rl2r5aijTdMrD06QRcTWG2RM5
epfLmHiSg8MZc65lp/tJVBriGEuBr0MC+40JniC1ENWw2jRI0jDjq598P2+CIpIsSgnKZGIVPT4a
R1wq1rbJARZutIROsJiLuQy/Pex0Bn3/2wSxxvwPoNABM4g6xwHKSnvzuLGmwEJJ+8zAQvvHucyi
Da6leqXt3s9+nle/BEVPn9EE4mxWKD6sfGh8ycMxr7QSDfm2r8c29+s+wA6nyD//BJo4jIKHCAjH
gGhJOv7OXskU8y/uyUabGwkW9znW1DUz/d9bljTSYvA3932K7FvAPjZx8MvXjwcmdKnbauNprzQ4
HWHv8nyzTlF3TO8bRi0bIc/Gt6ZDtEQcjDXRgSgypm7P16O3TAaOiJnsb3B7cqxQ06zNrqAPDMtq
k3NRa8Quo7FgTGak2coowYZ/nwvF4E+9e/EmNjuVOZ1vsUbF5L7YhV15Aidh3yZY9xix8uCNvFZK
kfrNKzez5vLphtvaqmlr1Qhvyhc7Cpau5Dv2DIZ8DvG0d4JPlDxs76JapbfQRu2owM2qzYWaLnd6
ELKNhX6YfiLXMRJ3Kob8EV2htzLHPntY8Z4oRXuYyeq0FuF+v3tzuDRyOIa9IG19yJNrkk1o42GK
VQ6DaOG2B6hIww7Wf/xMvYh43PsKbzOv1Z0YkC7sA6OBgNX9EIcttYANfSko+4C8S/KAZecMlOxG
o1VcuGG/+I3t2I0Coi5lK6z5SZl3EM4LmL+6lwsTYkgIy6h6rLyFxHizSyvQHL0Wj4RVqkyYZylZ
oa0APX0ji6DVzoFqtaXFn+b46OUTgOROVyvgk2MT/0lmH3JozrOlrEDl1OrJUv15jgRTO/VGn0H3
Rx4rT5DOrDQocWEfmHKIEZJpy0lHpJ4nsm8UzjupyxCKWR+8XhtoNjk4Efsmd0P2WqinVkx49hlc
ZZhy6Rv9JZB+WEPLK13ioeQJjMLp65KvM9Tv9CXN2/dlHQmHiCzrExjt1qIH0ouUMnCuU4XLrb7r
ouNHh4xGCSDVmyukR+p27/GBDPA5Dbwl/yO1ubewsw6vv/OedKtAc4v57ifbq2u0VB4LlIZpMDyt
a433Z1C4piy5SKelSKPyAFn/d4btTxS2S/NrM/T+YjMuXcc8iplmTo3Z4p9GYt1pNDrAda+D8TCn
0ZUP1+cPazcp/m1iwLa7PlnketmNZeF8tBWFvGbpYK6ymeOiyBw7/TbDLETEZobzRoCYMH6Der3/
Lm0+gzV0I0MMib/cDWignyLHCBAiJrp/M88GX/dQtdSqvpZ35pzQgi298oTqr62lgtAeSaPS/Gf5
tNRQk8aY7KLm8XZwCK0PIl+wCuCzhWgTHOXXFVvm2RoNfK/gZOhc1M0TlBFwXwjzdCdloYdN3cb+
tdGWuURLO9TztxT5pybeMze8G+MUJbXS7cnqDshrVegXO5kpcIePJy3U+uEQDmQSqyE97YOfha3h
k9LKoHo9S0lwoa8osCN846pwJ4TZlM6Ab1d4uVTgL/sX1B7qsS+go9pPkOB2efs3SLZRLpLTyJXu
0UQE10N2IejSqMwaItoKBnaXp3fPTKc7Gmnv+uePnJV53BtMP7/arcaiv0KwqZF143i3PUxR9mOR
PWEPnYwEZw8blfwp2zEN13aPh3o0rJ+oq9xQC+2twRjqQjRFjFFuobxR3DtfKtE1d+CiFznmZozw
MFmpVXsW5J5pe4Xavw4fUQLS1e254b1Njhcol50MWljYJr7icxVlolXmYcgLYLyl8wF+BjcxTHHp
TUBGMrnUi1y/nMrqThi2h2D2OjgLjKnStpmTNbZmsBNxJNdBPc22EwPggGZIWHgl0Bc9q3wfbK6l
Ur/F3zwonAEMOJM7G7/XrZg/yxmHJuDr8DUxRzBg8IW6hIZBbdhBnWO+d0Et6tdiXbnMD6xow9A5
fn+aV1f+T+Gsd21a2jBlteQTyO+1HJzw0yT1U5hLnhIX+/7ZW/iC6NAIIlzyQ9NLxehHB6sRRGja
Xr1bAJtLBlMpRHVm0IDvCn1MFr7tiz1BnnR2mfRatSUzelhFyB4Oye+yZawQUwXQBrGlrfh1AIcE
KlQpX4g9WMtUJhdOkinZqM0pLh0v03BaoodA2/SVlU2OhEJbmiXztugcuUy3wo/8Y3CUAzCxfglz
7st1NpNUsoQXM4g2ncVZigFlPVNpBALq2QI5SNpb5xR6BgyTsxg5vKPikCHmLAXw1/YBGTMrMMYC
YCnci/Kv2hSoktPumKDmc6hXARiInZPGKJHJ3vjgg0a8atelYWf3knrdlYKZ7M1Wn9flH6YhULlQ
2u3Cj0VybTUfVxONnz2HI+TYJy6gIYzB5hgwjQDaI7EtD+Zwg43RjAx/C+zPxYYWLvbnqMbODXxV
EmQVKNJhXN+4bKdi2NLd2wkSpSulNAZygOTL79TRLbRYGosPO1L5YVao68BLwPRYtRgb46ItE+9t
pWCsBmUSBsBwah1xCEBcSwD0qtS3lTOGezR7vmC9Qpj013CjAqCr7ziFJ24bkI1tIj664AJXFAHJ
Wa377rjtm/4R7vXjFXR99J7nHx8GvQ4DvwXq6bAJryP5ygw6YfbjHuTqQFJdQJ7CoTraO1U0fSsr
b5I/7vhgzDWzWbUmwTW0yH9v6PIuZp87SjATgoBaobyOl3uvD7ITG0V3NwyWa1KLewY8D7v5OKp5
xtFFs+q1+WbDNyg8qMuwZc/9YIS+bo3vNV0dr5y5P1sYWwAMBpQHWsoS/EUPCY5tNktlHNctmvt7
rAVftoWNgF+Zn4kypIoXG+rJAepiWatHQeEWQuZmGND5WhBFqvtrmvwedICPRpsl587wnu+3anYt
uMxAIHqUB6O7D6F+99CmTmkqKg4R6j1/uz25nnr8kS5yXjXMdYsUCJmeSYCNTqkLfqQdF9IpPTGd
aMbyi5EOhgA0x4qaqfUZrn3kkZWF5klPxlSLgIWjlAa5w5Zs1+MlhCNbcUAmI3ZjuVHXre2vPrrS
kbfGxQLfQ/njuu612rfBd8xbvganpIlkKmFPyOoPBKz+CMM3KfqmYn2Zg3H6X4K3Fn0/I0eFeXYe
QjBB77MPDz3sALo/S4ygPQ+3zVDAjOC2Drh2ggUEPOkRLqRWjU852G97tccBAK43v1VKIgpBp4cb
Ar98YpSYr4OBjSS7879a6R/x+0pqimnlNMJMUezYCzpTZ+s0MDDMfyU+q2WeqAWpHS2VeqnPbzvf
mH+CuANtqRTgS2h8F7MMsQYYEon6M2LFZ1Z3CAWESLN90FmSX2e9LlcGR9JMxoSbI4hsYyxyr02n
HCkkMbxGAdw+gzkrGS5ekOQC1E0r/8JStt5Jzhms1NT9ZD03LKx0JEGTvU0qL00X2DkG7BO2pGsZ
SR6VFXmp9RIG7iTZrMVJRSlHuGf+b8VYaRBcwa3UoDLvrpsQwcL5enUASjiM1PQEFY7mIlYLRmU1
P73W8tDOw+XZAmpL7jZIQ91crfaUG6iCFYOZsEHr05/p5v+2YwESsJ1wgD+7X9r60FuWCBnt8mDR
3z4B6YRWw3pTHQUsJXWQ9sU5BCp3fcmdKwK4v2YkPVN3e8xOoGHMNUS+juSF7FV7Q0jSQQG5/pzm
7h7sru1NuTYaHjGdORGVcnWpHOUqLnfc4Dt9tot0n/g1uxitL+s8mpQ+45qTJSJ1tbeccUP3Y7d9
2tLSwhL8T/8NZCtueSL8OkTymbdccbo0WxMr8vDdgd6Hzgfw1amSLxHISMwK+tcZ2E2TncRk+jQa
xKukJX0+pS9EItcxtgTZLcoux2rGd75dA+KGLXdTg6FACQxoD7ljPVjwpMANqpf25UeXlQDadBDd
eRE9D7Vf8j2pmLgol9LiUxPibVZ1l9NEAexhyeFKqL9keE3hBFYLKWvNZGaIBj5/YsD4tgngyz9m
6uy16T69KUgtk/5gEjtfA+7HnlVUxzFinsY+BOgUftufvCLOfcgzB515+yZ2cZ5E2ndjnpLg0SVf
PartwFR3Ha+sGW2qutGWD7JDf6ZocE+doLGoFuQWt8UejfJyjEgnAE8q5qRb20G8ui1yvjGEU44y
KoYhkbIArcPrccQDPAWvh8d6/uKZFJYnkm4PhnYtEgBccWMCQBNZA6ptVeNHcFR4ZH6626TrDkmc
WXFD++EFs8n5bEjCbFJCyqaQEuEOPQDIgezv/EfZMxdpJ2iKrh7xMDm6cICQ6sQksWrX06ABfaWE
wuf0bCUAxObyhKaqykT+resaetxgLavzk5enpcX0GqiI0j4+GWBOjT5vqjFl8M95oz2JdvEbi190
719sh0lu82tJEmIy2VL7ke8ppDDEzkrGbUjnxsn7RcnlWf1Jvazohtqd9EBnqWxXPASyWAloNGJM
o1NZg8XluSO9WRM9VKteTxRiaPb+gywNGfUdXWYO8IkNWCYq4wQd7S5frkN6QUv98AzIik+iuiVX
PL8Ej1kLkLZCrBYnmT1S2r68dSkFiVTYM/F+rAGxSN+MA2e/j7GmE90EyHeKTmmBcLNheHqzpQJW
nymWN/lbllzEceZ5o9FACcngimW3a27eSOBKX3/22hEUuELkaP5W/MSqlH0hoG/F0EQmPmTFe88w
uEZkZ0WGDmKnG7wqKw2pUtB5o9XXbodTBpqIeVE7rsYWJYoPG6QyqTO/KtYUV5ON2wzyy5f5GflE
86kGd/xbOfmvC4jSY4/LlkmTEzrkwq9qJoiPHI0GogyB+b/ESqdK2ys6tgca4AEJbVFm/+Vbj9zk
hcGxStCm1E0BgOs3wXchr8sjIlG5zHkOf0fZhw5Z5o9gHjHsLl0g8FiHPEFLsOfpAjM+qKhNxnUD
oEEl3CS9+OUbe8lZPgL7zsWn77tKsSnZ76HKi5QM+Yj9o90Nc27a4Eyp2tdL3Tlj1IjJZoeGfl+A
RwY1oe2u+mN2w9977cGtgD5eDVqWyzW/smBVSk0kb3uUZzgn1WpWKZrYybTMfbI58lK4uwUKHV3F
7IVGhEKHC6GZX3H9RF0+JIUvymKHJh3vqQz3SN0Xb65sKapHYUy9xDgSDLRozrZqprxB9DX8yoOY
QTzFIXFm2OFzFUwOibJeuZZh+R9+7r9Nba89lKRFgF5xgwjm8nGEOiWsfMoXNnYfpBjeAZYSD5cR
Bgy2UzqnLEx+OO+nNncL30TyanUkyvkKRNIW2O+km2B3OjuZhFlxcka1TVzMBvdgg6gMBsTvMN7S
+u3hCRZm5U66KHoW1fS5xn9JB/D0eHlnajelsgE5VyEMW86qfUIPIJ/v6TXc2oxIAyvK1iUZ7sh2
wMKfAVqUNL/4MieO1duGv38h88dSGn80QYY9RmCZy7JRf5BLHqG0odyA3fr1zmxrSvXlQFjIBazs
wEqDV7p7xjiXt1ycn1ZDJqPyMvDaGp1OWEh0xEoe4xSyzO0kYxcxAXTrwZ4pqEU8A/Nexrd6Zad8
DTl5gctuQZ5SnyRTH3ZXxUVXKzCEhwb8Tue6L6uHGjK6Vo9FoR2TloR5cY2c9UuLOmmdjWIyxzZR
DaU1/I3A0FrI23LvJ80xl4kWxBcQuMhlw7+NGgOWEwMwZn7x1Mo8qDjHNk3Ja/jttzuMboCtynF7
MxBrixfN+aqVZbEF4dGgm1OzM5PBH8onoBVuaC/kQ+nTR3yngh8DPhAyJncbceP4J64t7mA1hG5l
amrB5PxIjKejtpnSQ81csA65eXEnAXv1G9yFcv0KUMOP3lbrbGw9MMlh2QJ9zzyRbptSnCREPVvZ
CJBpiM0r/9CIxVrQ+d+kvdo/3O83KLD1sSb78PeMWxErmYQaL4wFBa8gHmrL3YieeekHKoOvyJvT
nunivMBheyqv7QIv7SfB/oP8oDTO+gnNLwt3CZMhkycPMKf4LCy/KlO/XHG3++oC5nS7vE3JXKRS
OgtJPG+3B3R9RCqxSETQMf2tR8pOMq3VF4in7Db8nvYEo/ix0sy+5oZm5FLFojijcX5YPBfz2NI9
Iutne8prJWXU7MeppKjVpWeRpPF72p/7vof+PFZ681xHFHWSR+awtJIze1g5qA+L7PVIBUuJS+HS
pK1SLs69P++nX2GrGRSFj27frZLiE/fO7Fkby8mN1v+U/7h+Y9/HT1rWrGJm16EQ92sdCMumxN+u
zwvbQcWt5tqdQZvUCtkAh1kl2hTO6aNOaZvsY5Ahj+04P5P2MauuCDmPL7AMyAIHl+Ocli2tszmO
r+sClQnMy+9HHqjm6m+jriEgdo+ZMzHgyNXV+frrer4xf6m0/9Erz7cajbpZCBvkD5TN7nyzdnY3
WZru2dkhi/dpE26GjO18mzM4fiBHw3SZtTWiEmpn+Omu4sJ+oiBi9V2Y1dhjOCLiD5H2mnwn/i32
Zvw2ElbD3h3qXFRewoI06ubk5LDRLX+Tr5KjDHvByO1lLF83es7b7Fnll1GsAf+AIjh3/9Asf8zL
HNqco516fFcT8W1W1KFxT7WS1BS53iT1sL1AyzOzB5B51sSX8G0EyHUPjlzpd0oehOieyx99mEzf
1TydqkeYLhu1aejaWd2iKs9+tGEHhfQZENyNegxrY/6iJv60lRb1ea/aNOGU7W5EaY0KZQw4lcKa
l9EUGrRBGxPVoTYIejuCKiobVO8CN62M3MNTRAqr6PX66JC4+Ix6yx71eYfGPoeC2/IMCdTlZryU
TX726RWjTIBAxW56QsSvORxJymJ0oEFWyjKxndCns70iqxvE5W9nfB1e4XP9uGvbD6kPg8x7KmBV
xlTlqH8rg68LddT2oFZPSVLECeqWRcw7Oj6+1Qq5tZD2b5Q6K7GKVHETBqblHpAPK0gA9a1cBtuI
3pKdY0gO/frDjiHhgaHSDvAkmCUwuvHmSt29+DYd/NUG6pme76hUoBYH4ck1h/EeHgfAQe/JS3Nq
scrOq1M8NxhyibxXEXfjAvRztHuMM/HRUpmb567++IysNEdjeeeAtjQSKhMoY7IsDJQFaPwh4EGb
5/NvnwwP2IewTCqlWtImXy31AAS3hWJWgortH9s/UGzJrk6NH/bTGBUjNrq6kH48nZ9tittxnyL7
WlghglyaYPVuESeACn5uL1WGANkHDgqdklBZS1eH5H0LCgXahHJheoOcbWss1kqlyeTzgAClzje/
+h8YHY3DsFwKanCaQSUKCqxBdcjsUjxUl17NnnJeZsuuxxLr70QX11SYHVXm+43LFmuxDs635G52
laMySgtqelmbHJBnOXP7n373hEpmfdZ8MGNmuV6KAzCqmlecmN/d1kzjoDzRqJZcXzncLCjZ4VYr
O4OgArJVItonkUe/QSNmUy0mSLSFjRK70kLsqDII1k2im797Vx8WAGuOIUBtW18biSveu7TkdfpV
rexzqoVk47btygeOWegxfafQiLTY8ApTWTlBl5MQWVcTnsDpzU4psRvCV26ROaVeiIAaW6P/DJd3
sWyF7+NT0EInd7zlq1XzR3A+qcQc0r94o1g0yHpdxwLighB4qRxQCvKeSmKeCwcfmb8xvNnHG2jK
LwAJIKkFMqP5X4yywMpdxKpMwz8/j/6527RpP1AuegFKhqzGBEXscTp8TaTqTSoqz8TSs4Lmuv4c
Dtu77zSjQC13s5Ik1QotC+WgbLHj9WXybqwER7E3C4XN1C7vG4cpw7olVm5vQVx/4yif6HBOqiup
FYNcoJSOhloDSWcBIBZd8y/ydmlP92YfCaURzy+srpng6SL3HjxSRwNnP/ZErAST7VymB59p351V
JI0b8WEUmUc/Lw9UbcGYZg2oH3TLSbLtcAQVasofU2XPwGz3ts+NvfRVmMDcBGS8hGaXHIKVkXN3
dMtFlZNYlAysxdq54gJm8d8jP2K/B6hYyY9pd1096lc6KVR2jZQZO6jj/lEg2Ps0j2mrEdPNBSbo
8sTxqVitGJjZGgEZCrxUzHt09zdAA6xJyEYwNYrdyIOb/Cg2aAexa6DUERLyz5vqVAQhlnP9KMPf
G0CVyrJF6VOtwhW+JoyV//rZdvSZTFLJB0smt9YLRqo1FeZOl3XAg2aNkz1OTdbb718/BuTA7Jkn
EZtL2m2XjrictEW/NQM5bK/XoUcVPHb/kQtixuaK8FA3z3MQreDpd5h/MSQYBaUeD2hxd6OvjwX+
otqaYFIkGy3wNb0fK9kQ70Z4cmbV19dfmRQdTslaaPRozDHMY6RjBsEqAcGLeukYHCZD7RWqbsid
aEQ4+vhQlXrjtl8vkRZPwaXYluMlwFUWBt7TCy0Ew8mh+od9f36I2mKEVy9yPc3sE43uXpIMQ5um
OwfPulQvo0bqZBZe6k8m2ItYINp9FDNdPQlMvb99NJ3WirE2VIWnxcDxGoNs4EMcf6yTx0LzFFVo
OHVljLwtiF4Lvm5TSHGSGp4SjR2k+vx7Hi5zbDf2ELl2UihdewLovLwf0gBjC80Hq02PTvIgVOpb
qUvROxK9r+HYBaMSv/uyID8yOIb1qCLN+E9aXXfnY9ho1O6W6B9KQ6BBQWzkyJ8kEB4XRgZZJUbz
0L/KxrOJrHgo8GqPxBgaZSrg258aLOIKmwkhAqm+0a1syg9V+KcOoUvXx3vM3gIn7UuD1/yXnypa
mVaGEZrNBGGMjh4TKms6tk75kLae/cEdtEaKB/SxM/kMH3oiYpFRJxAoctab0XggfuzBfxaEs7lG
+actr9Ua+9/sEFDoWK02/DqgEI6Z72EKJiKqfP8ePjjtOnwF96V+ZL/wj2gJWWkG9lkiFDBoFgKU
iJqj5o3mI326e2VkShBCfyhMgOpw8cZ+t74OT+gB3t08JuvLGcE0R/yGBu2Sl8O/QyWn1mpq3YsF
bvzCrdeNKISRcpntrfWBPyWdPetPjsVIykgNTdAuGSL93p8N6wrA6BkgWcw/N/Wp+XaC7YwvQlx3
ooq8k93zLmLYXuBYPJNLEHCE+oHy6NjmcxjkTaZSNyh25EsefiNVoDyCNsQrDkOPlCFX9DqkUQuQ
zKRa3MSy4EaTemy+dp7cwjaf2IOx+qW+6dwEe0GT1MFkwid/OxLOXKKXoN17lp/0oTgm3oFFBQiJ
a3PlGeHAr/QibzG4j/CXGJmpWhHGJIOxeYxJ8GzNHyl1iXTtVPy2aE/Yvk9j9PHf+JIeexwpG395
W3gU4LTAfeIS8hPEkQ+Xl1W0wkWg8XWiUn/EnYohDfVkIyNNj9bHwblJff7Pbt5CVzFg0Sn4grBa
ZClnZbWHqjdmVTRXwKGA7d/ogll9Cd2B3/HCUQcQdekx4+pTq9uQYDOzulmaNo+1kGydvJxBe8dV
LeoEySOH9yTThUJy6BBv2CetPAcqW8L8M4/NGJ6SsuRpz4S21im7QkkW7pgBhqWkk2Zrod+e7TPN
mWOL9uVuxrhE8IO6WyXp+SMLFMyr9xkGF/uJBkBGqSJ5h8YT9DoLZqs7dfkTaR5UhIrPqPnRNJYS
FHDXbcXO2ixVx6YDxylk2Z0h2LQNncyr0IrljLHfyrr86OwsOj3vJt9oJnROGRItW/lok1BoPMBU
lUOMFwyppaveJhrHKufovEg3Qyu+tigx8exSq67UM3yJWVQ3bxwm2dcdVKyIXzjnMesUuObND4bs
rxkfKONVbfjqr5YAaJKX8lLWyzoMs6fs/bv1m+6DShSYVZjwOSQ22u/A8U8DWx+QdpcU65NWfHSu
SLYxw4kQY5frzo7ComD58rmWb7rAeQkhEoeYKvfg2ZfVqu+2ZMOxZVOU/yfQTYocv6ZcWj+dxBb6
4R6M2GhMsgWkacEUF2LwxGZLfBXBiHSE+9v0j5/4xrlwaeVTLGDF0JBIgxurW+CuFb26f/TasJTy
Zg7ur9FGnQfCVm1ySe74ZbSV3bXDhsOc+myfIVi+fmvHWyeI/1Ax5ZvXKzbkscmZIeoA/0EK/OTz
xTFy4rTmtqHJRPRQkYpHxCr3IVftUNUDr6g7AXkFoWYnvtmwHP+qbMy1i1kVIG+i8PqJUxshYBtq
LoHuu2vIW73PSweKOmU1JlX4KEsN6DT62EPGImli9Nw3BU6Tw5poDy7Lo9vBBPw8sehIprbYK40l
dlcTdOlT9IChwI44yq/cXUZJVb7GyPoQv3IKCB3BhemYXFdPxGJRbvbcvuGKwjcc8NUypQpbDLtA
2lYD8xBcH9nAjJEVJxtEEEE00q45JP/T3StxCV9qE4cw2DFIpGINLRXH1aX+KN33NhrL4nUXXo1Z
LcWX7sumu6Tgi93E3FQvHXrWmayoDVg0Ny+HiC5AQ9tXPMejEsJa7tNp99Bhc+iTgkqysvCjW+MB
jUQhUuqBjpujlGoqGfZaOnIE1J/TetBBUgJJwj/5rJed7gsmI1UcUxwXrvQoUrBMm+Pk/6aVVmLE
mJxfxM7UpCYYv05KnENyL+Kz/94bfEiO7MwtgPsWohgOJEJbOE1gxVs/pIccxlcZv8u74Ok8dfEF
VgLd9tgyJeWPPKGwylnhwUy3n1k6gfb5FE2qMmf8BMoBp7ndfv0Mo+EQoVaveMQCrCM7kF6WX6ys
sOmcwIj+X8GtFIReMEHax2CXOmQ3Xqd6lAtGviACB7swkLwTX0+FUZ2FXGh/n0hdhh1l2dMeI4TK
dulN0240O9v8k9AWhrbDxiiY5YDmbysI6Uz6jEGWBZwGMIBE7Ca3bB0KhvueHYMtLLp9AicGbC2R
jmTFePDSLQw41kuuBTCwIa2W4Vp44pX668TH8r2GB4smbMmxrchjA+U6UNX4XMUU/osy+hEd38ji
2yuASOMjrME37wWwkuF6rJhebkI/mQjdRDr4xT+iJGoFVLGPVeoY7JZVK1eLmMiAIxsGUpTFijHX
5Obv0uzdo6XSdVK5lmqV/YFB3Kacej/vjAIzO5knOwlvq1yWjKzLOfm6a9zc9Rr/Uq/U1BCVZWOb
ymS57t/DixflcUr7+4eNJkUEiocNKfmT5hB1SOHcPoOtMDLGMswfT4WTOarLW6Y2ubg0HgNRFIPO
lA0iBmaBu8bOPxRxL5U8TT1jqwGtvQbwYhcDEy8NJI2ANAIW4t7fEdpnr3oVKvhQiyiJ6kfZ8dy+
I4Ife2vMW5Ogaj3CFDNflav9gj5MH6yzzlEKYhXV2pXF3dE+pyhVqEzyW2F7vKf6q7gqe3l/icF0
Z2KNEvysYF/PNSPv96B2kYEwEmUOGHyjIciDX1j9xo7ewVKg5q+1JInq7BODnUg5ASqtzEr8ZEzz
eDHmG+sSfbKZbi7DDpt1TmDLxp5pu5K6jW9Bol2/e2pCmdFzhWmoiZEEvlNZEld2GW66PwBbO7VW
rNMJRU6SIcK0P8J1FuwHuGTvvd01/jrIo/JVUYR22k2E5SedHg8W0pY7lSPVL7jvGp8D78Z7OtSU
gzkz9e3dkMvG2fXB9V4o8h2s7OQoEse0F6kXxQhY5xlKfoPa7Kpp1fyPDAsQ4TIWn7UYK81YagAr
/Ht+C1Ou2QGpuJ21DmCqL0fYubinyiPMEQVJaSAE/qdjuD/vWq55DbXcXediXGjIXpUumbxzbpO7
nk7ra3MoBXLrIUr5nnhDjGBG2QvoBIR2E2U+eHN00CMCAHeLJ7tUhc5IgQ1qjIU6MyXZ+UE+xgTe
1fWw0/7k3sz5pW1OJ2UqoxH36ZTtil+eQnoNKgp2+39kvpcqkW8Lop5qcFvOGCG8j1ZdvkKnlRIM
xsZmatTCPlqKLpKsAgSLrMnxTMWxpkdvvDOQxe9aPSdxSH58UvxAk/2LbIMSbjQNcLEWn9RInmm7
FdvWsRilImKoorNtKRkxGwyY1WJMylyyfB0dykmDhgD9++SAGIjN8jYPiDkNhdPJt3mJgkWuMxgZ
W/wQN9Opn96VANJjnLNXCuRvI89hYc44Z4dtQTstr31BMJcqB6zccUgCG2qvTumOY/9US8+y9VqX
z2qBQqcFbrEfh8WCEhZiksEfcFGIUZry7Vp/5IwoKq3HCy77K+KMIPWemP0n9ABYiMvmoL2PnIvX
wU/yPdcdXmfwUU3X5e9XM06uSFPjO5SND8tColsTrIxIDlHPza/n4GT/cQPvE1s24z9kjby5a5jc
oKGPC3pvLsJvxLsk3vkLGQ5KfByWPyjCaF5uk+5X6rfT3mIduYTAwFDbczbTYxZ8/Er7rFuFVZD1
QzmRf2zekp37mMr6Q1rSVlKstMczczrN/GauTZ+2+u3T0zQ9MIfymDp6O84C9SXId97JRQ5BYP3N
Lzeuj0CVWXAdIJ6Fd2Tx1gR/jZ4netHSvcqzp7Fs6o0PKMInR4a8YuMd90+v+WbSc4cxsxJ6yPhw
1GRKKqjSFVcNWsXvedIEXktYg9Egq5xOo6nQUibLyrJROaRRaNb9WFVYPAcuTPPOYAsXlW4Px6QI
BuZjm4zaEzSgKuJtNUkphr/igg8K56RmAebPhRiPSSAVpMF1mjpyJBAeEB3hdNSlss6+wshOF1z/
wtWjKRFros+uwjYQEOEGo1XG/EQdGUvCiPKYsBiEG4EkfeQpuhi2/BHoyxFxCKvsTLWbz3kOLL6O
xLmq8fPAfZUfsCBjAPNLcuX/Pk/f2zngdweBSd/njco64MXfRP2HzsqaUkeo5vvhA+HDT5HQ8oYG
8z/oo3chWpa7mJsAukKJIOGSaqN815MwV6FeJddSoDjtVa2qD2KYJ0xAHxUi7OSOmjon4yqneU4P
MccwFpuJi/X6M8gy0BW3KHq4SvO2tZ0qoD7/ZqXHnpcuhIxrsPSiJvufKf7Mtw458uH+kaf+bMkv
Nbw+hi0DgYYUC/zkz55V4gCIRW7peNpNzSYbhbRKLURVAZAB4ogys88YpooQpJbnZPalRpP4Lt+s
zbDhtiIReBE/M/1ZJBV7P6f8cyoz0OUj9Hou0ZwxpCbaTzMqpDXVDrSGRcbwjDvsx0RNU3Af8Zxx
hy6fsPk+jQPlc7nq8jF9sUCMbRE+53RTkO2MXg/2llkb1mlbRul2Rl1xYyW/7sx+Gh2gNgdM4G+K
aoHymwXXcVV8isfqsNKwwE0z/HY0Aw4DoQxeKPAsBc9PFx1JHLCA+P2GxWqiscLXqZ/X2BGeCUpE
EANAd/eC/4HYgTNj76eSbgJYOfe3rqCtMLSE1vsUqHDETRYihOZkrOPSduvfKt/vwHtWX8ynIahK
J94U+tGkX4pqDrFeHE+RGcozDHmebUFaZtnzyiNLTXybDAu0bHNoVIIpRAmfHGww63IZWLr3CtdT
nV6pf+DM0HtYlBqiSS1YGmdVkCYQ1jrNtsW0v5dt3bDndLH24iABu2LYRedGTDS6qEhA/wVmCsq2
ovttoVpiW483QlRW3GkWgf9jUDBuoay3WPxr6J1IS7z2IzzEE8CVq5vorwyM+40yIK9hMEAj2RsH
OrBA0jpkxQ3qKj7pNtwrQ5eqn5JxaRVelgeNV0p80/0Mxa3IKfbl7OgXht0oea7/5hJfANqTrdLv
C7ul8d7BhDUEYFyY6gBODUzndNkqVv/h51l5wSV9s4KZP2nfWSXdHIpG0fPza88tvefe8l9lkkFg
YN7z69TtBrXW+BpXIGgBexjyWhPN5+8ygY2UfxAqFuNtg5CM6sQ411D9Pes6UsKvkiMgrt7ISvqK
DA4wgVeM/7mSrD99NuERQmW4XohtdA/Z8q1x9gqy6Ye3bXv+rrQDjt07eoejpIobW3dRWpQD4ZJl
k1aS1H/xPidIMIOkxQx9q9F/BO4DJf04ecsTpCPE0DP8kYsTcQOBQk52r+27yBsXH1ZH5+4wg6Vz
/TE5UDzHlcWLIWUuzBbOu9Cd2pvMnpyXfB9leE5R+wvdumGA1one7pJZW4eHLUE7rGZZFSi5bTZf
/jfUgDzfRvVic6QeUkgzPTmRtZfXJW5MaO5DS2B/sTKWWyl7q0Li/gP4h3HAT5XSmq/0FxB605Ra
54uAOObMzt4xp+mIWykcykSglFlze4ou7B77+TtkSOZ7TFUPYCFGa1v8D6b1sEzhq4tAM1EogGeW
WYCqOsWdzs2deA+UXImfkStyQVKkAn9Sm1dRaTHpScO8upax0csZNWnUgAs2F0BAgwHf2mguHM4E
m9ljciXEn53Y4GCtY0h1mp9+R2JMY6M4h7wavKNurbycSi8SvYN5VkaZCyqPTmpimU1B7XuJbEOp
BW6BFHrJ8hqPcXxtSKJyMVv8FKsFTyRGNLjqfPOvwXOddRppeOC153L7pDS9eD/h7FJvamN+Wcoc
DqXB6DD2B/buZgh+vwpa6BeLnNDIUMln8Di+QkCkgx3l/3BKZzd7sbal0wfm44GMPv2+dBsp+iIl
m6LanWvEFZ1t0jk3SgM3GxtshoVqU+IkVOr2rGX2RNmdRPtYTvnUsPXZyabTmk6R99nHt/M6mKZG
VQ16dS+1T0O29yPunuAlj9XCKIhzwZTTIocFs5hMV3g4dYoQQRFBPJIfS2/hy0+3BF3MzBIpkK2e
S8iKw5EA/fVD8FfVjNyS1MQt1r8RTK3k2XIcYbqJSlGEDE991tVGL0l1Fp5DMMPK4qCSV9Z0DP6v
qJ6lYBa07KE1QK4KU1T1bat9XDLM73St/kAL5fzN7l6B07Os2ADQiv9aXg2NeVEvFu51Xi/X9aIh
v87SOLNBnUYWv0kBtOwHPTrJ2ZH+a+TZnstm8z+u4GZAR9UX0Ws0ft/VT2BQvC13UBNETmFvkOZi
RPX3LLqZyIQKljuXaylHoE8TZnzWPtC41WisNtBubDxDIi0vkvE627uMVD0GN33qrBTNXQkLwWNt
rWr+SfsxoDZufJ4IH1RXenopYrT7SwyLV6ev3qVYkejbaJmWzB5ws7MZgHi9XEv5h8X2WlWDQVVd
pKqL8jkL06sB0MLnwngYwR/l1cV/3jWtaX7tP35po7etoFcN+02reBbc79tgOurZGhK4rRfLhRxE
9efBf0MSYrCqFC143Sq1xGGC0mCyo1/l8sovqG4mUvIlpJOJFFZIQr7lbRMz7rtcD7zm5GASXxYT
hOcZpVYhRSDYz3XcIr4O1H3SdOK+O8WO2VNJLzPheR5dXtAclgdNs8IfnENHdA2Zv+oJ45lSS5GI
r9BmaLFvSlYwplKhqJFwoKJuzOz8YKU5RafCRe6Kw7Oamm9DGcA3ZHWlJWSPc/TIlEPzA94JLij7
8JhB7iQPIX5PXSOrIByuLpJlEnt+NpBXcqD9EbDBh0GfKfkLgPm9HxBKH+XLlPlvIUDSkRvJMsv9
KZfsNSPl6rPyREMJ1c3uR7omJ6/tzuGAebPpN80+Rszj3Ckt/Fd1KRldpuTR/71xHDiUTXM2RMKR
PrQq3twVlpt8smMg/ZKL2/ziXT0VXur1i7OQPEAtUes79lT2L4qsaosPlEZP0OuZp07whVH0fvaJ
UIPJpXrAMyX+70JjHqO0pfIhKaPAeRxo3lyNWfbGkmg4pNA9T8cY58TrouATq3aXGQVJ+DtDlLy/
MaSfnUXzw4e0h06eu/xBs4t1JB+qRON8p1WJZLFWyXEiLTe2ZgPQtMtXS0LgwRgd5b1b+xC8Y/QP
pnXJklGFBIKY0d3+7op3d5LSwplk3FwZCHNjjG+wC4T0DD0rHGUd7gy4tbJTCTLZCKeBOc8EsFMa
wbnXaZvFXXboaBoHussmac/7jNHn4WmNl7qUKZJUTAOjAEuNlJfXmwpuHISNmBrFanZeXzndK8WD
H+v+qj+KJg78wgq8ZYzPyC4k+/B3nhH2MWS8u4QVnXiozqKNl4SjCjrLN1rgnptX2x5+1p9DsxhJ
EqJvb8qju+66vdcDn8z4MrNGo9X1OlJF47Td68tCLSkus0Qb6Pmd7m5BxrgQBSe3HCdJdTZfIaod
LKZxtbOCDU5mrfmr/PB2CR6tx/1mGvG5ilTNX2Qn2qfoRRIgDI3t7IYTJ0R69MVCsLhUIGyCX3sA
+y2qJ9kWmAKeYV8eqocwS+Y83UqSw9O96vmtCW2rRA6akW6PnuBUClePLjqSQ8JkWjtJRY7cahQ1
HqtWC9i8/G7OBv3O76MSIhMv8CB0yOdpxCraM42rHzyFOvLLaYvEPfbtrdtbMb6T8c1PWQKmNw+z
Glv6M76Uc1XpVXzcxTzkQSL8v3avA1Fi8taRn89GaJjtRAAlwvW03V2p58fsc64lhYG+9dlgiuhN
FNd2Iz6+0vmPbGD5D2N28m1SO7bg1aaYVbHDOIkKAA4s9Ce95aLkXKqs2hBhBMnTfhERzidTqA9p
XrOn6+n5y575P43EOL/AnYB04+nQEJ2At0NBROIuctDgJat+dURdHHOTLPWPsYDX3z6+9JnAHwg5
QpOebsx+jZMe8grnY0LMOhYPyZY/BrTTSABoJOz+gxjLNIL8tRA73PVURIGxpMO/PmUhiNHp5IJr
mm1ducwS2t09ptUv3cdNVere0ekK97xrzOXnma7vfdb7FN12LT6WDbWh35dCUvla+WC8JQh47PNn
dygqtuFz36it0cXK6iPrVBoSLZcz5N6cMb0ELZVCGaH/Mra7Dt7SaHScoiqLBMcrszF+7xrCeSMu
F0srG5I1Zfzx7ouTLOEMr9IeWCW5Kk2n/4frLU3aGr3tBV8e8MnK4bUcTGiZ7tZeR9u7UAwuOw4I
3rIbTXbWGFnN2Iw45NnUF1Q1fgQT4lF6K+QqvRiBcv8qp4qmWnF8cLRsnrlhX62PgVL/S7TKRKEV
6DlYfjwZu+s9e4/CUK+eLpPGfLiOAxt9NzxjeYvTWTWH4kjZmBeO1W4kn16maI3bFRUVjBxzd40U
91XO8XVufIec4kSdw3Oe89Cpu0qD5802wcWzfkGZRYeRsLhb3VRE0k/L3/3Y/qEXfjvsuCEkZGMN
1Y/5utHbAkD87uIsdUuSatQZEBgAV0/uAlWeH2kxXQkv7zDloSPrykekKRj8IF6lRoVojz0mIL3Z
Rf6E+H9XsD3zTnjSDrbLAKfarm1xT3zOahgDUzBOmb93LM2z22YPhndfUu51k3GDC+yFEVwVwlBQ
2d3eCrN+gD0+vvI8Ng8vXgFmXopgZsPqCaC2EhwApozSNjhadMX+KfKF3Kp/k77vBNoTZXeXkffx
E3OUYiQ8SuEsW1kMjaY2DhmKsvYFC4p4pvoKHUEGTM7auWFYFy8anWjkmcCLoIOSs11w6EHHMJHn
T1e2m3XZFju0klsvsxl8EllmrvRv5wRfSMXePwqVLrSOUKWiYwwFBbGXvyXMP9VJga2xFTzv2FcO
pdiaIWfTYcAcctmV8dxS/MGWStQeXIqNzPiVINA90CsOIRpBMWcGghGRBfPUH/mmWr9kroOn8fn1
ofAeuofYDenAk/KLbgV362Ysd94uyLDp/h/zCPQJXRCl6yWB2VQV/76v99b0eND+aC6zmXtteWMa
denJ1LU8kjsptz7pk5YhAtqCNvtdtJz23gExsSxtfMakR1KXaxlrigk4YLYY+pJDDuDqb6GOkAYv
NsNvA3x8MsGthJb9HViw8o/8DzGiG7AtT1X0rSuvp8x44Id3/7gOO9QeHepI2NaoK6Ca6SfpyTfG
O3Bm34Bp4C6RbNnq3b0ARXveFfQ8RRmGjEhJ0AexdMUK4n4VIsFhD4eXfaPYNVqIVjIPLwWE3+hK
ZVRfNzLKvZK8j/Aki07Z5qJ5VwDKR1VsBbqtI7cN9drD7BO+RjL6NIWhFn7EGlim3HAsB890GDeN
ZbOR133QFr4rGGgJPxBZ8WUygo8AwsfcFzz+YvmrRhzw4Dt/Tg6UzXrCu2H+6xoPP6mXCjjA0KfE
zKzWScLiBmkoa4+gP+fv8k31TjTOWf4tK774eFrv9/IaGZIs+oO9kK/zuLFi9Mas0cWDZT7e1Arn
hLM8KYN2gisKeV3bVz4sRv7XmOsb8n3UH6z2ErLgSeACIFbJC2/yA0NuA6bNwdsD/9DLZFbB+Q9q
y/1LPzxJ+NOerBWj0GcqrSxRn0F1FWDckUyPZol0Eor3tmYDYzNQJLpY1EL7jt7cmIvTLKArTWn1
YBH0kmOmalROxuZd2Fi+giV6OS5K+6ImxxxFJ3jrBVb2JW3ZRrGs8Fi7QhP9aMvOaPiHii2CCzE/
VeSsX1RDjqOmr6Td1OhJVTf7FEtFpKp8MWvMVFql0TT0N3OJ0Cbjksj3RZwUs+qWW8mgiHu/mgeB
RhdVOYvlchJwq0Dscd/a1EAop5C5cosudyL5FnkT2RAOB6gK7iClDvZHyJR/9j2X3k36kmrcC7Br
g+lWwV/vG8BX23pneBmM+9jYcdqcXT7G0F045O+vKQdheUAqVJZuErKCy8JGL+PFhMsm/TP71BT3
UtPrBJD0gWt6AkpxNmpXTAudfTwV0nO538M0usDpkqM7YwTyVVc6Gljz2VgawU+XuIH0EBr5WYli
8en5T90C0tPVtc4j+I9yDb7yyZD5KKOmWDKLArbholL653nfq+82z9DHWiJhQKDjdzjy1e1onY8y
50xK4l3eBfFHEVK5wgL//BXo1PqZGVenIjvtjfoIXWzY9H03kmNO1lyWbdS2VCssI68q4ei6sVKi
IvfpkXTXw1hyG2IxXcvu8Fm1gYYkc/AYWu2GXH7pwrJQYLS0QmVwGhZpW5epedmOpVxWLCsNCcAS
Fc4fpOwOKfo5D2UQRYtwNl+3tBDLZUv3nZL31a2vCHZNVx8tq5xU6PQmllE6do23hBOmyrxU0oq+
YBu81QI8H7w50+0ajUYDUUClyCvs2+i19Yhi8NlR/NLdXEoSsgEWo0JmpnjQhGJy+vl5yew7MFJ7
hw/HrT1T3xUHEMR7GeAR5kHc9Higgel3C1BzLMb1Y1aYez6Jo6n74UnvUEDOwFgsp7877VuvZNZo
Y1inQduSgQrCdtO/ilCPACZLsNHJa2OWBUaLBYkc1IWL1vTES/0w1GRs7a2yIQOsRu3YSrUL+f0x
upkoczhR+DCJtI0FY4k8/QIPhn2u8Pg8Wqre+uyx/JZ8xGPuMb0983KF+hPNYH394We+77HnWjIN
omx7jcyTn+prJu4vDqg2skNNTRxv7GFoWW+cT/xjCzqy6SPChwIhFPSPu/TPpswEKKTW5V5cNXa1
ZVHRo62FXXv5klPB7RxnA8E+tNby44VoJrWRC++Mmi6tgW1LB7Acslsg0VS+Dnc8UHbmbx40FJ7J
ND1f3idsMSLoPCbMHsAj9SMA7HmUFliuIMSLsC/xckEXgMB1msJNhTqOY0/KMsQJiqJvtjwZkUn9
vSa9llGISRvmyHeEz7T2g2JP9+NssJTQaURibz6eWMiIN0M/hwUOiHFS3lVaknsEGSdKlYUrv0CK
R6VsAM+krH1jK/7fNSvSliIz7OSeW9iykN1EVh2bEnwgTJtkpK3Zpz2yKT36YOG3kdVamBKQ6vgI
nbX/y9RKPLaqG0jHThwST17P6wOUOsbYsiTPN/wb2EwFRTSHMqN1IYp0pHK/dRLTHtZFa18En9Hx
6kMIMYh1/NFLFwi1nDYNx/rAG67MVY1JTj16yrt+zTETbxEDiL+kv0EbwPolqXmKGp+xE235D3kV
Q5SyR1D24PZFZAzxioMlOfSoTj5E5chnfNlEpvA3MzxG+1/XMjG3q61goKYvIxnWoZxVlLYd4Djx
a0Jfj9HsCp5ygZLWs4LAlBipwSjCTwjBYs6wQZRT4rQmeroC4P7XnUwnD6FqbB8cY3LL6iMYyZqn
9WPX1MPOypnyHI8HCJYuK9fr7nmhrXQuglPh/HmnKQPy0KV3KWDGiDjatThus1dohjLVbwIqIax1
yPqyVK9JqpAbBViIhCVmZu1FBxCWodT6c5tIbe6LKGnowv9ZnYZCUBUFBTrsNpOfmLlL4HCiGazp
jLHi7cThvlGCDJCSWaLQtpB/oKv64CwhSqB1tFWvbqaRKFAyTTEvDONnCmTJBu/bK+DvcJcsfYCf
ELh9OkShWMeu0F/E4M4Bn7a+/p3xsHA2OFWNndPDwDuounAG77KEspl5dbwBSF+c3v0NnHggojkd
Ban3+b6X8376KyvDDfBc55xXBDqoUk2tDnTsfDOG4LVYPM5MBHo1Qekha47WgzQasjKzpzLpSlt4
C6RHMxr75X2zRRMH1haH9lXJqnTO9/3HTeHqX5m/2eSwq2uegIlq+EmH2mjA0fVHZOeHVRJvUObi
Al8yut2z/TA69s5HvfmUKQxqoDACCs8v3jRtj9qniILLBJbHWt1xrXXrOFtdXCYFnUEfBMK9WGka
aKZrw+LCHjgfoidR15pMKQeebHNlNeNo2do70ipChLQ1+1PUxHehILa3aSYQE+kO4dtNGuW1g7p/
IykFeHVnbXh8rpilP+DdlLqaWT1T/CUAymvz2UllvLXmVgJhJthjXK0YpiXY5qELdCK4fsme1qkF
vp7z+q+Tr+yTgC3S8lWxErQ+n5Oe53b+9FAfwP6NSRx/j74GLGtkiVSMt9vO3KAkgVehXQRGq98N
kklQxMaUnHPU7y7euuBqTz6Zg4dtlnUdeavNkUxzYMoeTcwAosuyTc9dkEIoq3vgb6x5rtrhFygD
cjgtqI376XOrkIs5CiO565Hi/BLpMr8grkFnFied6nB0METIfluGb+SF8ey8CyFfClQvY7xZa9E0
WAMBwCYmAdkLT+vWLr37lGmEGW3tOtGto8v41cVcV3WCfOS1mvBtyWFpviGF2xsUP0DWXJJRFXxE
Oh8rMg6ZCztabOosJgVlb4spObCTyeUrDAlXT4jXozDy8DOy86oB8LMFFl14IMdXGt8i/Cow4fJ8
gOmAUPb9vB1i4qvqQstAMxAN0mB/h1UmkIger8JdCniLwqiSTwF3O3Z+94lz9b3ssjqm4i6U3lLy
Xdz93YkJsKX0bODwvHtzjmtPUNQSs8YkXAZLtXXxYy7IpVnphNFrrlhqXSJUxMiPlIuw2PxpIbmV
y2HncQu/ikD7X766/AKF3mqYT12hEz0GJtruGWJ9l8L6Wpn9O0R9O53EklkWfMiCXxtZH85vc2dj
Edr50gBpPSvk1hLN6b9wts3A1d/oqvlo+5vbBUyxgDwEMN30rxG7aTwFdyKrfODuIh7jrH4a+pBN
r/i9B6WoqO1Z8xAt5pRm3aX6c7ktC1PQWHq1pptNBzE/xhs3HqDyb3SaMCKYc8FZToomDjUOLRyC
4mYNRIWD7BaukclRZE5/VuMM3CqmihyqB1nq8OerIbuZCA+rLL5dvKmHsVLJw6UX1BGzFVg84Ztv
epe2ez5kjx9x+gtovRNXbSiGk9NRH/fRwce99Ho1fdssEpCGjkzDGP9J7m5lVJtaqBPSAIuJUzsZ
/QtjUYMjKJ5RNc9iBG9eLmpHLtYnRG1/Oezxpnm0CexGdY+F2b6hHXosRbARX5uQvNi16OvIws4W
JgDlU9arCCQEZJRxuEniefW8gjoYfVNCa2seiZczTomXlH4nxSjg4JZpXs48hkoPwjP5SMRETqkh
xaAJYP4B0CzVdGL5rXPEa/FcslVcFLcCk/qUNSJm7De0sB4W3AGhmnhbU9T2un575qQBnDGYCPND
ec7a4e7GgajlWhaYGDCzI884hSozm432MepI/sQ4iMcnCtv4a3CeMHHn5AIMv5Nwb0mmCsSjHBq0
BTWq2ZQPHzCL7c0sXYvpfjdpuq7AOoqpnKXmqPZHMx542Peveq4JacDi2KUUPBETaZosr0G4XI9H
j7NsddG9XXAqRRqp0I6AJOUvuYc7ERkBmHlqRV1b4FM9Y3Zq+0rt+c7LnagZAdaGKo7MIOgPUJOv
JMrhnu+l26fgZYIz50t+mydrd2I987hVT2Dq2UhngrboEq37nz/llp5QKrFufPm7FgV9yFIhm/eX
OFbEjVKE9iAfw4T5mjEsgADgVMWiVrBLPn6Lf5FP6v4ntpd/l1KScBQuzuzOEVYZygl4tNk5wxCb
RcTSUzAkyNLoQNmuXxL9KqzTN3PbH8l6skskPGHgZdpo1swCuBS0H3Ff2NQa0F+nHqICO40n/f4C
gVZG+1QN4QOdPuqCQVpiXmlIkup4eIb+MlSg87lPLFHNym8Iel7R+37/nQSRyJ+cjxFh8eltyUi0
/9RH47KujiQ4MqJRLix+kZMEM5Y91/Yr/PqUmfUFeeXWaf5NoztOEtooQ/Wa2zq79T1Q1CgnWQw4
Z7Id+gVHgcPTOWIbFL63WlIZ3Tr8T62pl8r/mtm8iBw1ly054hQHvSeTrS66cUjDsU1k6UTtu13y
FPNCzcQICEEYlDW6TjJfER0YdzUW7uAmwjvRfXxIt5O92h4+wB7UgNAYlMfsEFZ1HN8hXU2G87fB
uuZSMHXbCg8YvjVlcoJpPjxaVGpMtZUL4vKkg/xKJrH9uzNvTZNQrK7B8UrWIB/eccVxrtv8jQ82
0STjgQUvByOnjsBaZmgF0UztOQb/SbeOLHf8zCovsMqxjMtDt0P99tJ/l+5EI7x4pXVD/qKl0Y8E
tFBDcGxPli2YmpV6AGU4ZtKkgaQIphKRykf8g/BX9Av/rJ0yIiBHUEB2pNwJtD3zUNBJDpP1SbIU
7ZNF5uN6rcFOiWrwbGbFMKbNsFwAzxxjQa1XsW28WC8y1inK565YeKfSHdtYLJTiH4wAULpuWQGC
KS7k1D1brpZIj9YefV6Re+32duRJtU5KsNqJWUhS2TKT0gxF3Gz4elYxitAYZM3K82jo7CDKloHE
zWVA3/tUma579AtbCgJjS9Brf08aBn+oxo440u5coAfAUq9gyXsqWaqtowL7cIlFS7bRkgrYTlpn
dHvP8tWjaXf2AAMkMVpCZ6m9aFaOsrNfzJS6YCyJ0IZhyb8Fjb/Ly2EdluGPD1Ipi59Ikl9jY7iY
b6rKCnxopuGswJnBsMnCFTzweRtPN2j1pWFsBgPdIh1khOv3BYdjm41d4v1iYYM96Ypsjsw8Pr7M
2gM32uaznXjw3xSZz6AATRXAQnLsiHujcLGCTGs2iVXhekmkkE9Kge7KL/UB6aldtStOusNxAdSV
F6H+XWOPZjwk+ijC1tnQLSDg+6PPo9abOL5b5LCsOip24S4AvAGdWELd51bbpvlQ3QVwieQXez4Q
bSNTG4pk9df/1vhuu+Ri+rc5IwEG2c7cX6XoFn2bRXYjIbpPdM3ymjxwII/yczyDKSe2RYHo47h+
NUjWbDObne42ijwg1zUVZc/vli6j/ZyW4aQFj1zFV66QvDASsAMGBizPmWDx+AeBZ8vy4lzUDak6
Fpv9TJfRkk4tA5JfvkLf8lu9A4XsY3Tn3KYOVKUJDAJFG65RVLK3Mkw16ft9ocAasnGz8ZZadAa7
1QCKCZ5xjk22bYK3AibnnAEyN3ygfUdLebPmRNETEM/kbzR/WpBlftUWSQBUlKAMnMxHzZ3gxgYz
Q4FDJR6xda2ZCccKa30/WiAUbOb5DdMTKAfrj8F9F2MJyrQRXOiRzrTyQUUGafwkyb5B6AetbDS9
7ymzR1YUCDwYiruUtAU46m/UvymLLWQXLh4se3TnmXdYsb8G9fDUebEPncKv9HMaAADK/QkZfxwP
2eU6J3cIj8yx7fz4qJk1ST7MdnFwD5xYygw+vn5sO1racd+VC3bbLAOt6sYCAydkHmq12u9n3ha0
WWVja6TsxNra92I/ezYINazzB9DR0QaP+Uhs5HQ6oVpl1Dz/hQoAvVdA01VasXEVOE+8KexccvVh
hpLuCNrfn0VoQ+d2fq3Jan/7zXKRfkdnX5OC//v5vnjKBOqAP7JKRL4a+OpXP/WChjlbC+SSHpMC
qXQ9ML93leoBMk0BFp+o88Y3KToPgX55xF2m1Pb7jcEWMIbVbofrsR8olpwfhEw82/6zt2M2ohIC
78brpR719OfjWyViBvn3t7exJGDWwVSPvLx9H4AwgsbOaKw2fptCpAtVnsDC3vAkF1c7Uwd/5c4x
xzmMJd9zpTwSKmyGZi77PAmGOFdRIt25v7U/Jrhmr/RcYgw8ZcfrdX69gz3NlJjAaN/RhEk0wbZ3
VDKWI9vRwfCYSQ/5ZyBZn8Mx48fBGW8Brrl8N17sDjuEGJ1LAZ0icDvUHBlJBdLMQav9rQSAog20
p1TcC2R84Xb5e5EOEoQhhGGUPHeTtomTGLKlnNwR/NJOg3JFqjWZNq+SoO713FAujk6hmHaFGnUT
z3/Buyw+Y3YHLoYsileAO81++hoG7Ka0ywt39luArw3J2ORmvx5MKXBoiPXU//Tr6bd4VU1ARDvK
51FmU9/FvRA5SmiM/Tvw7RUoTvHY7ZquSKmN/WL3H+qw16oOar63EwexMIa+6TxY1bKtLHvgMjqT
l8L6RIbl4N9wM39UvDSBgf92rmwBNNs0zSFdgSWAtmqG7ilWETxOg6z5cISAerTQSwQ6jC3d7h0+
1kLwftYhygPqkQkk8yqafbSuEhVtNCeGZYiGCx5bqLkAvQCy1XQGiCUvLVYwPgVqYDNvdLs/B1MV
fjvEETSBuwpWMkCP7eh0uktU94BTSsb2++FLtfJG7EC042QZS99/OpcWc8lxXjyPXWInieKveTnC
iU2ahVBpXxct2ieI1jrPOe30JLnRsFjkvc30xjU14+mP4v9ZWdRvoHbN8Mvvz4bXFdaNRCX80yCp
VSwtxS7ZEWsfDzi/EVwSieUif5ikENbfvBoYQ8CF1G3XHSUXuuRFUjpUOsU9wD+Pvn4htIyWKXMQ
VnQBEkFA+Fze3u33PTQesQO3bEx2tonjXub2EtkTtog/6eZjh+ZVK30Ogs8cBdZbU9L2u+tUQswR
nykJbaUBVKqF0red3kHwrhUpkxuaVgcD7XMKQUF1Yl7kUo/NqEeMbDP9IwJPrHmUzU9sVq8B8PjY
PY0wZ4+71jqVKVC7Ozj5qxrRiL/vTGFwNkVUyCe4MHGp+9ViBgm5QWaSu4WUchSYIjHr6/Iy2KSe
rz6p3H047MUDGeL8UCQjYhRT8brlwCDySKNGFJnJNcpoj4Gpt+Q8QAtJxhue7mQLHG0nh469uw8Z
ixshvHJ/73KWrKEWMu0NQ8djFuu4ZZVfTpJwvmlHWBWegWntgfZqrlOqi3d2eGhLzePts5x60WsL
/PhEi8XNKAws5QP++OP8wKRiJMXTdDoEAde6sMcC1vZwG937BJjFFdkeHXf5DlBBu6NCY6g1jZ7r
vZUPjLXe29kWogZQBJZbBvRhOOyr7yCzq/YsnDcJGTP9aQnvRBzlpBTna+L3bcKgAC4/GisJSD71
yqqIcqnA/Cdm49ghC6HbQLRfHt28bLurwL2nwFePFFHOvjxcNZIkVC/qWJHRCBP8eTtD1YqJU0Sp
LovFQ5+0S7RXPw/ZFhGJsRP912W63a3PKWyGEbB75IJdkYgDAJxG+8n5R/R4maTMSEVeFR4y1PUn
MkNU/UxyfwWJX0DQE+jWFMJ4ON/2nnSWTWMk+xX8HoRQRuo2Mocm7zjdxMn+QoukWEJctNmPmeBG
jiVSpQXCq+/Uwrd5Xt8CMsRq8ir4Ag4+/p2txV4hU7U8E6xXn48Uy9uP2RG453aMYAANU78tiCOY
4Qn4HvDfOa88oc8HldOussHR5951dWvmaMncCTjAsxvTaAgCuK7m7v3qyfPQSTRXq3hJJbGqgubS
RoJDatch8ai6eF8pNgW/7wdS2Zpvr/qbGDUfk484ll19vwj83qY8IASTjRvvikYAfF28uCK/4MbJ
sjSvRO69S7Fu5dgUPHYHo0Bw5cLgUUb/lRUhlxW0AXiZzyAzE85ms3Heiva/d3eG+mWrXA3CDiUL
OoBCEud7EiA7cCsI66hhlalbdraEqpSCZH4TIeWcNO1R5tJ5kpdo/vq9x1KrVFZuuSKnRJeqvAF0
etYMkOPeNO+kdoB7rXew1QgLIM23OHLjk+eb8E+uwI2XEYae3iMRmguWQ2UF1UkSUIwNZg/dbRw7
8/FocrTmntAXC0hbQjm+K8LkgC+O9XS88YHfDT45+5iYV7BYZo170jb+2Cw+BX5W0Sm9toiMxIdf
LpNO6Hpg3/p4gcb/om7dMHTEnsm2CXyrlORYnC6yySHAH15qDkkGsa3c5FfmAsoaE/MinUf3PU37
MVzZZhBijYfVhBiQyb5qFF20YG/F/70pooDYVaM1vIatvotdq0V0w4zlJkJoHFfLzeMhfGErreBU
DVyWS2FSQ/nhJdiFZYjJ3JzJdL34X/VAVSQSPKuKp+HwdDqUfR+DDrYUU8LCDxbjddgw5bs6BaSM
bdF1YC1NF9ZFlnSARrk4rrBB+64OAFXjTEhV7ZscSzmf0giP3ypUqDJW9CjFRURacsDy0L9ojcvC
rhaTl1EI7dEvPktiDTiEc69s/Ues50WOsBeXrFgTVUf+OHDk46U8acj3t63l5itNEeS69cSkiHYJ
hWfC8RDSY4Wow1ryI0SSNUuVDLuRXi2mg7nB2KFkFJa5PjEKwT86TovsRvNxZls0oYn0jbpceNxy
w6xR3nqwP3JmKtAkrE7gwrgg82zQUPTP5HcvExKR3xXhNQsSHJ2e8iZY+eXrgc4NO+Ly5dUo+s9A
yztEjs9HvDukn/b4ZQ21BJRp4lO5CYkP0lAHFmyq2RpiWXrx4xzDz3tO+Nz1SBqXj1dCSa2KrN5C
Y7r3TlQflpoQv5+fWOHLhJFXh5hGAkZodAa2DGATZgI38+YXj5ly8orO7cFMIRcEDpy/UiUrY7Ic
wFpB/SHxFHm+ZP9FpsiJwg6LazPobriaMctQju/mdw0HTDbUD1JsfjI0w/2JDmy9rQbgW+jrc91B
dWWbyjRZ8zyda5V0PQvJ3N/jfSbDt8oqmwFQrC69idsyom3t23lSs6TyRhVAq9j3wITuNJPv8xAa
f829FWmL85UhF91btnXDYD8/uj7IUawBXYn8X4Q7Xws0vlorfG/E6B8uuYJ1KjWaRrQCz6sWOynN
9b0sMQ+eWS0TErgeGIyXzYX2+sJ7rmZhowyXbm2TREVChRvHACgMDF3ZbMw6x3VNGndSPZ1VN025
OGdsDyUL04zuAgXLjVsRv9R4TwpK4l37mreKrflP/ocWSyla9/eg/krUQ7dABiitvDUgBnOkU1BC
p7eEPMfRiYqxxrXcgNS2Y+ldXi88Co9nBkSiyAMu6lmNgB/4yZAmrRO/aq1ZX/O7jBWMaAt7HfEQ
nQ453VW61PIZRrYs4QygQq56xhGxxOfY4hfu5Tlri6AGlpO4uLbrJNupXcA0povZknbYvvDQHhX1
wpUv35/qUn3OZ+LwLzgevcABZZv5Jkeqqf5HBqRy4z9J6twM8LUmHQVGsRUK+QNxqzpGDKvCsTf9
FtswusZ+Fbyd6qMYQVR3qCAd+D5C45PTJshJS3eQgii4eJ3ies9nGYENgp5ADLCdUo6gtFEDNrsw
hlgJxkEWloXwkeqb5cG0U1go+PK8Kljo2YvuiED3eJ5WdtrDAbkxvTsG2/HFycGl7hcqBtk5JThD
S58a85r8VMgWnHaLhP7RYxl+VdSn5mRwJteK1mxQ9eMzGQUDGacYdwym4wExxOVsy46t7ZDJHObj
7lj3C9YptO1RUSyPFJG6NbCXTfz14eeVA7YC941CafhwMxWp1p9Fcut3RIDtNsh92Ek8E9wNGO8v
Htzv7hSX2dD9FXZNYIm7EIzjgtGFLNsqvkoAmh8uWWisYqZoO1zoY4kRtCLfEwPjYllxMVWeStSB
oceIoOcFfOphLdgHVb3Jj/TWt0qQYP5wyxU56fr7X27mYMfY8tcikgSMkdxgVYfwX7mspwflYoLg
7DdnZBeQOdG+4vlOpzySPDfi4a4ocK8WRZUlX3Ba6BSizW6OcO0sQynRssimarHxwzZQiOJfW6TD
hOXKPnQQaiMwC3SWFU5UH1l3s9Ufq5xXGYYy56MfUb3Va6i6jxhf/yWK6eXdGnHam5mEVVpnXtqq
MPHaivb+3jQL93HJU2nY4Zuy1ilwz6hKxeS/pnNbJTYM3AwhBi/kOK5oD+dZJl9eL3xHNfYl2e2v
sS/RlGrDzgwir6cfaPXusAflVAJhDQerHLGo7aIYF8LvIriCzUbvg+7Tlg2L51kg6kc1M6/n78V4
AGN1GekVYFK/XwKkN/NzD6ysmaUGmnbIFHGURe6WECK7B+dgNYT9G3j4Bq7OUGmoJfN8uuvPOXHi
d1i0j0yP5jmfZqrL+ei4k5U1bis4mFQnFS16Jn8z2WSr+ytzH44lM2OaF2UYz8ogMtBdPFJNRQ0d
lGkk2r2XjUx1ju962ujRGsCLciWSTyO23c9H1fZ4QXsHyQHwPUCSkqBpjuPl0Q7BUBEf4aLBn+Yq
8iiQp6qEVls3XRvgwaW7x+OEzMpiRRJpt7783Rru0SE5kirLrQV1A+4yGA+kYZXDlvKP0FZhmlfp
bm5gzyTSmV8vU2+zARGU/oc7/jSwcvA66F/k7yOzKmFiITsRmG8zRCf0pzI1ILa7pUmc4XsN6jD4
mrhz/X7Qb1mwcP7hWp+y/Z7s6I7UnhMJrkC3MqnpPVqWFvmKnAitImXeoC67IitImDXqsldJ5BCb
KKgrJCL4B1XKhmxTKisDIeACUs6+whid764lAsEb623B6KzcqVwodxiXtuMSAyDJg+xYh9qMAM9v
2rU5TxdBvWf6um9v5lQhTtB6kwg18Of+1tziXxMsq0g0QxmaFVzk7A5iSwdwVXuQ48wcMKbBx1TE
MsrmJMZmXikfimx91GSd5Fs1hByn3Q27EGyuJ5/2rBT9vhJ6LOHaZKTUJH/X72GGaouPr9LYAYSs
4ybvuQ7n7Y+uXPfb/DDu/VhqL0JS8RJo6dluPXPJFdh8hd4dcwCu5+KkgUo6nDtZ9n1HsdlI0p8H
w7z1JS84yD6lFl+FG54w7uRsWjfSGbFevZZQ3aRV/2kVoyv6Y02ufT/9bDjFkMr3VkFEjxp+0Hm7
dWbQa8pa48PfI4ejS4tXy/OzFDQnBs3aBsy58mRV9aiMiOulOcTaTfmA0FXf4212QH4fm0g3LONX
FPUfavcUWZAfxCQwtuyNZoXamwFvj5FMwBMFPwRDHoKiGlp+Ruh7Vhv9Zgfb/+Y6kv/yFt7ArnQ7
XOuzafM9GWxgcJY0qV8v5f3C0d+tvtJfPx5JRG88zO6ZKhuk64Y18F4WEKRNtzawZCvujtqSZT5N
COgKOsKnZVxB3+VejP46nDf2n/UZ7SvNudvnHusz4nXq3zANf5dfdk5xuYiCTDkh7Of3kmGyBfjb
BaQ8wJ8OOH1EJpy4kwHRZaoNUYe9H6mmeUdXmV0u5UpvLfsbPQZbVsCqIrppDrpec2UmfcNVP/0D
pU2QIP9r8X52FkGF3g0xFIaVnhO8oZcqdyaeiUo0+DioIO8c9kzs0Cbq4PQRNJJeq9NpE72IxFjZ
DufzBWoJ0eNNqoQRhaXCUmoNs2VgVO9RJEJjeTqfXlAsDgnnRetPJvNVUSePB4fHHozZxLu+8w6O
4kUezdCskW1phX92y2sPVamK6IhASeVcS/aAYmUSLNlemhqkxX50M0QEmJnQJQDwpPPOHD7nt4HU
gfHPRumoAOQSv06Gp8JnkulYALvSk9g66AxBnktyhMwW9JGBDQTnsDATMSHdDHSKbm0JT+5iVyUi
hi+l3V7aWZGfYVcind1HzBtwE0cw5PtAG0/CBoIAc7gTTrkmlgggMw1T/OvOO6p6RSTk6TCrtFdq
s8/PFo87U3HLQpWm6SufdDlMrWKCVC0kofZp2f+sudGQGMkzxOG85vktx68E2tci7EDeEUeq/kQR
q5CjpLTcLcWJdHVfPhRHZ7XJngBDNhFsJzNHj5jP9ZdSmrLQsrdABTHyItGg8yqwrAuFz/G7SifD
UvhfSLuF0Fn7IRKU09xVjD6135V967hbXAY0klir6prSIRI+J7m7luL0jBpQoSblRcVk0+D5bU06
hqvDtccBF03Lgl8zt1Ya1jbCOVuWbJXT11LDAnXtgld9PKN7gy8wW5ZoP1x663McH/b3AG7VA0wH
JNq//dh/GYdGua1AqAUZDsniorsG4L6NCsVbiYeBHKDM//u1PtjVcjDucZ+SRejegqtPtvYqa8I/
GETMOXWp4mst0UrmoADOOQ4Ye1hmq37vhI9ZUTLYkgFkTlOSe9/ic0kPJX/Rgln0UshV28OYgrgE
QKyV52bQGrDXNIaFYKBxweNAofEWAzje2OFHbBDQctMvdOn0YkBVU6QSFyKnESlpP9aLQSQwg2y/
QvH/dPBMGUydp1msJRj76LUvAmxquVOpkmPkyYyOcvxTfqEhbC/CbAb072LmH1uWm2KJ0cWB2PEA
TtLdpW3exIJWc5mME2cZ4JcLzR9+ypN0agzZD7E6drqAXXNUfJ4kW5N+3BR7oiI8SL+Ms6fORjdr
xp05dccVl1mKThq2/JmX7gZV3KvrBzLF4GXkaqPt2Hs0ZzTj2vNJW1RwoKq/C7ohoJd0Vz61QUWy
/VzEK7E0fvL9x7Ip7Vn2WBmtvrrGf35dYQEZaEteaFSIEGz63SjMpuy4bSy/vsA7bydRhypD7CdX
8VX6oWg0pqL7LhO/arlT/fK3MSHxVuJOfMa1Y3X/72LUiZnec/Wq1jV1Vh1B1FGcm6b9ALQptB2g
KticnNn4MBovq8/8YEF8+iimjLq/610i+sbYe93tNQ4ewRwJ9Az0wF7bcMEQJqrRLCaFEE7NOakM
A2uqe+S2TLxtxRA40W/i1guEaGXAqEh3BJaFFjDpbOV+Z9l3ChVx7jcuVb0PM63lR5Paee1eFw28
w3Yk3JkBSkftyghZf1jZ9VrBOS4p9uGHeuSaYjyqaLWGPP96+9/wtkmTCI1WdpRlFw4ySMRJza8h
+jOhRajqUsabFyczKYcTjyp33qdRWOBWY/FZUly7JDC/dZ1lpQ8Ye+92AqmGMqKPVHes7L2Lq+eK
5K6ImJb4ifdGF7YKN5wd49O++CKqf1KCsp+xnTkJlkvSKr3CoQpNka1jeEjj++O39iuIaJ+a862S
W9NwAOvydBtoczGisnguNHRsS1FE+5eeMG3Tp8w1BOBv6pYn2fP8S/H6y30Xt6sRpoWzgqM+sFe+
45874m2vzHSwIGypFdc60LmC6KHJMqMVqGlIQOQuaMTtSZOpTYiz27BNOEFcMA6EU5BxHmtoWcav
LW3MwsBkzCrKmQtefh5/2brYVbEx0hUodg71ijYnJympUl1Wzt5EzoKAF5Mnw/LuSpoQcr+nhdlj
TZ06Vh0RiBL64wJt8B4P8LScv1W47iACzm/zGKJCbZL/f/am7eMtMiKbsnvrYY4x94XFzsXU+E55
1tOer8V1O7UJPnErMLBWSi4BZRtl0ATSkA6Vi3Ce7Ll/5G+KGwARFfNEZgnXKHlpJvPiZzS1hSKH
XLU0t2GFGVeD4jEko6fIbHfAnjDv3d+dYG270HSidRfcTADIekrfMcI7RyRQKbZjfl2a6ZYTrx41
VFjur4gwTMrAfo8QGC6HlAwdWARZoddyVBpIR6ssctxeZp16OsZo4qxhPkI+PcvH18FJGF+/FPyK
EcGkvuxTv5tEnzuswQ2dH8scNW+SNS3wHchhvYtFhxcgpQGZEwJNI9H5EKW8HIOyP5vQ98PuZSb2
V0YeQfbvlNNDjEGMjfrhpOMWdxeiDDuH2m+FtNBBgOM5PdzKz2m0NNYr5XxxCRI6F0gwOVdXmNAC
pjr5ZdOd9//xyT5olN7Loz9YwAqxUxoYG8prZ3bKWplbt3MCoylxYsjC1h0L1XfGrnQrtVujJHVE
lH9PV/xi7gtBVeX6HltzLPItLOABx8mNgrXWMFyQS1sxSXRKhjXT6jstkcrM/D9+f3uI7Gjzrhl/
M6w42NxqRnFWR98oJM1zKnON2dE49xBqf3/fetAI7FL6+ZlCggi8+j9/2Ftf4zN8vyyrz18rSwuB
yW170FmYkGnZLZOZdx923+6zJaMVaspirXmJej8nUoCrFh2I34Y05uPF3U3MAgJ+rWLeEXp64Ykr
VgK85a3KYb0pEV2YsABbUu5E3e9S8sDFHgHEjh6+eM0ppaiRzcTwPFufEQz9hEbBgDqM1Xefj09p
6EkZ2l/dz/b2HZM3Hc/IVQZCaLvNs333M0aFeiu2mz4kMaBC0WntqzYfsmOonE+kVkgdC3z7v2DX
18Nco6Svco4yyrY/E3eRd6inOQvRssXxqTFTNnQKx49BXdwshFE/uh9f/HqkGPr1i3W9ZuO/qc5y
FfvBIaog8U7vAXbbv7NcPWEZagV8L3vZCPr02lPA4DkpsCkFtHNuvL7EyapajqPblpjNRThgdSnw
Tnpe6X+VO1qcPybb+PJvHFVT9PGXx3gyEmP2rcqM6u+7LmZj3NWAwy9NJydnwIb7ZT1AMfR6pgSa
RdTrAgxz2RrdHB4C5FboLouMGMa1nBUHAvYDuSA3LVVa/W+s/xi7MVmgQu3JU8qG2nPPDkiZDM37
eer6tHcF5B2c2meVpQ8me/SgC0C6ZaGJYEJHJ3RecCcifj7wIYlkYzuDjcKMr38TR534plDTmLoa
BBEAtca1RLwILEj7T1hIFnbm/Xuo2EPJVIJ4fw8pOC+alZLibq9xbWyNKWZb4hNy7BFQr5vZZvhg
hH40pF9Wvj9EtlwAc8m3MAbinIc1UTjtRwaUlyZaiaOPS8i4aARGInQRmpy+anyz6d84wvK8LlA8
GYRN0uys8DdjJHSLK5nlQ5AEhkhe5HSt4BYUrNSrPWE/mvKpv3ISo6bNmpkqrb9UbvvqjbhMk/JF
3i0+GLIkLw2XUR1v6Jm5c55MVliB3fZW49YHM0i9dshiPcBiGjP2Q6qr2Rpg1z2nSyq63y9yX3TP
c0DY5eurRaG14z9+YdvCHN6bvi799Zt1ltabSUIvvZI1ZAzynDonzs7cTVpy05z0crg0sQ2Pesdl
eBltIe2k23EaXfA+IbXD2y14XQ7ouEqkfWBBbOs6X4nUxAYqu4aJYlweIDBjetsB3rZSA2vqSwMv
0Tx0hxTJPwmrF6e0i1OgtK8vFFvAen36/GWVQNtFqxqR272xDYqIoiq3LS5tZt2Sx8y55ayJt89i
No1DxIK2bqqEeP96kDb9uYTnAHJWBp4eOVXn6NBABGXeXWYKGVEo+7YaN5JP/vXrUdLw3FAfR2wV
XPqRtpp2O/ihs0fARIRMzuiBBuMjcFx3gT8LhASHZ2JMmfiLAB3HBu+chTnYM81OpDPvZtBHfF6t
FlF4gW0l4axl6dpUIcZe2W8OAVpMU6fpblpIWjQCCjwN7GAG9AFfw5QtU7u2BB+tOWpydFv2qtfi
O4CKh0Qw78y2W6y6rmn8eFyYJXBCOz6i4uatkBpktBETTnV/VxjVkQ/pPbW84Z9FYjVrhDEndJ/L
J+xJxL0Qrw8c5EJ1vWcszv8T1r0m1HFSytwUe05SHy/IMg0x0drZ30ABhZTiqqu40sFBMClq5fgd
/gZOYpoz4WsL2cNgKJpDzKs9vj1a5s0v5PB2hfTn9PaqV/SHp3cvWtNhCIGUZO5PgJik9lfbM2sw
XBeGCApD9h6hxIBwrmyGy+bQbVS7GcOCKsQ51tgpg2rHIB2q3LAMaIuObH7D50WehJ7gw6Ak8/s9
TVJX7NbUQx1upxWk706ZIkThjuQQuo5a/bEswjxyu4iw46ByxmT0+H3wc0By8CJCjiRR0TtCnUh1
YZxL/MyWQWinpCu71bqvoGjTQAdJ905idEEXuXlUp0vJAKr8Woo6F9J0Irg6ueeW0aJRcZxOm51H
8OpBkNYXc6l9QYnOmFDMqi0hq6arEwPenz16Wg6PU4uk1R7tTP9si2Ns/nhjB2IicJs6FZq1fQYL
kERB0MwrTB0R+n5vnYvJ4mTP6N0lZIK9xyW3vITQ4HFnFm/gSMclMnNj+Q9+mKporQiCdVMBiRzC
cUj/yrCr7gNFf9WwhF763Eqh1+MIJ7G3lKbyFQbd2zuTfateEHcKSlwIAPtjpJVL3BtnL4IMetbZ
hrjsnPZmEEKLy8shQudRt2/YMAzTFp45PDI22naJMnu6rTNu5DO6mOx7Bt3adWCJRa5IHzu7DzMH
jCKNMOIR0m6g1eVPynBxjdfX+YbXiedX730nczEFWmWy4ORppn5KTOFSwlta/vNWo0dh/btv0UrX
h+0MYyZudyMABtTL66j9EPG2cqXvZ3z52qdbrFp51xGf52AzTudCRNHa+nheb5h+2UjkMJz756jW
4uANj57KYya1DVXNTi/1afbvNr3OKuveWYlHXnDF78biRNNXzcZb3QTEZ11oU5xculuUu4EIw9fF
HSHvCKV40Go5muwQoWDUgRj7O5H/kFKYaCqyeQh1mL9j7q6PFgwLNPpbLxGbfm0quDvTb4D8RRpy
s/iJsLdIqKpiVac4NZjG9TO+3hRaB+tSIuGjm3uIuLHFcWIiBZz+c9dZ8Sb78MIueBCNbbP4tyS7
DXps4qPTiS8Rq6/AyOvGBf+/S6MbT301J6g8jntzrpsT73lkdOgCPanc8UYim+lyGOZeXMWLdUJJ
nzTGLt7nkLRNeQQ4YFH/nFk7/mipFlWfzagnYy45pkOfyzH+mOsOe4CQQAQpy7YMO4j++PgRQKa5
E2l54ykN9IqB6K8HO5X3T9kXtnuL4eV7XdDcetU6OeWqyN+k/C+Qi75sYP6lgczVUpPDua0a2aNU
Wu3GeOBHqm9UGUQh05exjHXzaRZzY1rm+oug3cd1QJ6rS85lb5eNHqJzqy9hBT/Jtjqx8L68CewI
5gwMN9XMpXXhBhcbipRwMc+J859JeSttZVwXYKdt/3ZopYhy50jdQRyXoIOVLpOrCNvxIJuwBcg9
IQK5f94nvhhTgERsrXTbZXPlvNE7IL/8mXgNOqfw3T64UzuggHRLE53rX8FoVMaM/xYJnVwo/yMC
IubXoLJ9pbHAmXzhn3g0t3rh74CAmWBVQuOcf20LYNtECdeWSJW4t+nBGdFl+kDVVlougmoyCCdj
vvxOnuJncJNbl/X+3L3SNowBPt59VaT+ysxaDFhXJPhf8y2esPdJUK0t1m2ZCsfJY8h1YjYh1Amq
tdtsd7j9tCwDc9N3a9Cx+F5eOLCDxXDF22n9BcvBvwnM3G91eccPhx86wUdMN1haBfU/g/VnBzpb
m0tYJSXpGlpGZ2qAI5MzwKWPiTNvNmkXImuduwGBT626wcioJOGYOq38IXy5JzV6K3s+n+QbK+yh
kDnzM4y3OrcyQpxz4Ck0vLLDlArkkl4jUNVFplBxEkPfYs8HVOcX1f1Iy62GoIhyB/8z3gJbFQ0k
1KGMeTbHzUN2BPp1UdMoAykQs/bf5yxJARWpuzffLuIYHBdNxcgLU1ds4FKqYXuDfGxFTwgHO+Y/
G2fqi80lL0gYGPh6CQg18KQFBGeR05rq+3sdLtMzWJrQLijpAv9YfdKp7LGTKm6pl3tS0qn/mWcV
jXgxjILf+O1EHMAv43fySa484H5Bh71f8IglMrWFNzWIrmx1aM4MrUNo/ngISwVYZI0WX4inyipJ
wkNG4kFQOKpNEjd8qpfYpXXgRP1LVPw92rHZmT+Z/JyOR7EDlpQoahteNyTaawe4sAHdt867pxB0
PcdOYRGY/Zvxsie7u9pTEgkFQ+cGIrgiD/9VOAiQnmvzIEzkxS+nZ8pytqb3U4csKkxF/eCuNIpS
0a7vOqA2JR/+r5EUZZseiX7jno+xoSJZpQ+OyccfTXReTTtCfbbmXCvOAw1inOjF4iSvX1xMZYZR
sGDUL9cMUZ5TPrePojmtOcBj/LAqdkSxhjCtg6CbpfcAjznVgbf9l14XrN0DlD/YKbpAqJnss8hZ
ZD8fcavbCGwdZ5pLURYZ72bBPZN0zEK9hxFENqTJV1qJiuXzARzBlAFdErSEoQdc0CAjcMvecB4W
ZVqM9cXZjUieGEp8HDui3apj/cTcfjHQUtgP7DZlSZxjl6T0tOPHSZspcoRLHssCRIHCrQL7Dg4Z
gIc2YvUvdF6vYCDoBOlMEyX7JAcNwagte37HpAPm+sE2LTp9sMzN+RpLjod8NwVgMyoZkkbI8mxH
uDjEKK990yk50psLcdTG2sBnYU1esZggJidb8X+d1Kd1ljTWrlV0esd6br4XuuZPfAmLLK9PZbiS
9K+oR0JliI40szDbhWO4y6hq4DlLoASjnWGXvACCtkMg8yDhGQdT4eDi5m9rNzHTR+4uKaISRwxe
Z7+XN5zRyQHfWZNcCVbUG9/9LGb8wXAloNtV1HMHCYQ8xJS/TwE5XbR7Ac2AD0KLT96ZbiQ340x/
yPwkkhCgUtSNsOJhl7Pct0sBHtnt3FUT4fmclm/4NggrBNPMvUX0s+bF9PPhd0IPBYVP+2Edv0+R
ZFyOoGKVh/vmOCSk/WBL7MHIbZf5slbkgoix9ND2WH+zA1q47g1FsHJ0HxJrh2ArQXnAu2Cmf7QL
Oa/n+bzcCIxN0O5tOat4haIiYDNnbeIUzxIMzjtvPOTfclLNcvPuwqFnrjNkoWn5tsCELwty1WeA
bj2N2StjC+NFgkcwaRLZNcKe9rP9VKuCyh1dihz/8lTlujIOrno+qCULVYJamY7uBXv6JroXevxj
PCyT1aYiGYs2GqGS/rA34gsQEryUuEqH0B6gfzJYjKn9CMKmOWr7ZPy+F1n3z1Xq4FA/i/Sz5Y+A
wqoUntYI55gKEa4Hy1dZMB7myyJNlRxPhi24+jVeUccfOVreX6yDyJQIFZ/kl4kXohUR0LXF+CsN
HH/KA9qUf9wLkDcIX8O9Gy+5RVoP98+rEtwsE3BG20OoqabisNYgajCaQ7+j3hvQQ1gXNB8Vbp1g
G6tVtOor+VvTfsROwnxdOUcfzDok/0dgFHNfprQhRUhe9omsazzf/rL429f/M98iFd5TQeUk7fcd
cXP5p8ftTfaLCEei8oYUz2ZWLPTP9nTvnfOHqkEUaJDWrC+N8E3pKrswUpfisUf3CpRXdCk7esVc
0rAjJnlSqZMA1clNQq2OePvgNSanZIK4icBMDRe4wREEf8dHeL9AJxfDjO4C+yJI1fnkqpSQibvN
nzaiXtLvtcgFh9liVom7lW6/6Jh06p9d+slx94EHAfvQKeFwOOEqNuEA97tp2h+nZJKhVgKH0k7y
0bHv6kxGuF4D9KSaw/cOmQYjP5SM9xqFkbaxCAE4CgU7xbp+X5mB47ARyUR5xkg7BnHhs7/RpJYm
xjFop+RbbHXZA7zypiH1FiAKYosMajUfsPV0C/1GNI53a4OX02oTeEIMV5wVJKjeWOAEemx1mSH5
Gz9w8FzOgGUBitOHrBPb+Za83CppD2M7fpF0fT8AVYbiFF9ARYjRj3jyEdJniZoSgdJ/Cwb5HZ7d
eKqLdPa4NKCFiNYrufBq6ttUAdEhLT0K5TkyZ/1OWeO0aFKzwvZ9qNR+De/z1ZlIw+mqMltvsJ2O
aZ1dlnP7TTg0GK+ZXwDsMJy4LJKK6mZ8Jn4fX8kXefbg4k0rTV1HLIYVDnPfYxuLT+D0l4HeiF4w
VVPlbmP84BGiBcx1TFXj8Rp5x5xsHM0zHVZBLnBwBrtuuJIaWhvrZgnYY13zBS74vepb4B8uk4wr
uNvuQTI6nAzfychSwgHm5RYqLhxTt9Ed/VGBMP31P3QAkfogjrImRPQ0hwl5huCjidsYp2QzQlZJ
Q4NVnU1Oo03vXf2wmcaWF00xV72ZKMKSdh1f4uR+1ick2vi5O3Nh04iHjvcKxQIpjZ7F1eM/YWmB
XgcWUZG0Etnq0kYACjk/wTS8YdFnquWgeOBBri8EYQ63mlzLgrv8GxienDOHSuWeUUrL+9tcLk9U
/FeKnhwdgQMmAbk3hSO2dweIE8e9Ot6hVYeWxvF92DUv2A9v3UVBTkRh4LXHJbDhjRCTTot1YLzz
/CZyeKBL7T8Ty0utuzm7b/ru6QzN53VwNx0ErrhT7EUggjrFdJtC5DNr1UoNvBNkWWwGotkbVe++
GDwAe0iu+rJcP3l1oaqA7skoZpLZyUhSIMj2J2ekNbfUgSLiyjr9X0FCFBVyS/K1amUJnTG9LEEM
QYbUnSrGgOdGI7MOF1vLD8FqZjf4vSI7Z2hQ9XJ5XLUz88E1TSouOjo8f2ksv3PqxBgk0/if6nj1
iIp7eLJyEVWEym5cHy7xWY4owQ0qaNYUgMpq1/wzSOP8B47pXhIs78AYs7HIcy8btlIv2dye2WYt
GoUIpG259wCZq+e0MJumimZcUjxbT2mGpQz0Y+aA4+foTKA5x8mcpcXHiIcwUM/6/pqqKEN7KJuI
lirWgvedvRd8omXqYtndpSOKFfsL722bthzWRZi8X55Aqf8h9GUibJXzDLkzYmvdRdQrXzPNro54
pMQXMJLUYhBn4CSfRb35Bo6+hCnBaVWiAtAJc66EGKy8FmA6meEzU89Ja9zAavBstwtTQ/SRja37
dsbMLELfBgJ3EBwsvp39mVmZr2S5c5ISCOLNkirQ7R98iswwcVGp1C8WgXihl8dLeD8Kugy3+adz
kRAlgmUH3uQc6helQ023Hp9XyQcl0VZ8o3IBBoV2prr0Qo3GQ3qhLbHbGcfh2HKhiHy1pZ/rnoIp
HaBNs5kuVbRTxIsGoEMQ0Zm8cmx00+yfew53cc8y+BT0c40F7VOiw5Eu9nzqg7Uai1NUsfiKRDkK
PVVmLylZBTCr3xNUhhvEfpg1yAqVJxIOMGa5iyeYybmug3SmiNjj3sRkLxGhESat8NjrAWjjzfOO
YnPgxlejKpCObCAfIcixTeEJqDxaET1Jj/POu2y5OjKtDd/u/iPVJxXtZ2Rblma9pltHYmI+Jcx1
AJ/Ep0MOEfj/TCtJW/vQmzV+9Hi8i3uE4huVvqo2ChsnJxvVtb95jcZoj4a9qySyXQ3/B5V9GXXo
eZG03ZnW0hnRuUKgivvBRqjPU58qzFGvdOOjAQo1k0vbV2TN9s9wAgwvxhCv5JOwgy/vdn5qSoSe
J7i/8NWbElmSGOPWIwH6vWqgYeNFHC3udSRJ1CjM9QDf5JP/lUfVDhG7JK9aRWe3YKel50rZfbQx
ryQoOt7XJADtr03stU3ZxWp184wnYeKwGVUlFzsqoY1wlWbrHRfE8grFZ/z4QoRSu9fs7IGdB5TX
iMYByJi1kH9zsePgj609YiTBlXfN3rAYoSbqPlAYvhpPH3nN/xF8OVsWxeQwq06ayRy2le6ykiqI
xYQUJJHMtWmE+rLowYqf10ls1k8Yd8ImwYDssNYsltqTkKDBeVPHIKRV+ftiuYWPZzmfx1k0841a
LctPNXwnDsCT0uqlJpLQqCJPoWaKfTTsG5zX92VrMhysrDbzRJib+LcLYkOQhpcgNQpQr1w0h7+/
291y/mjAQdb/45XckFEGHxfgMHEgauoTNjFVw+KXC1v0SbNlUJD/OIwgijPVbgO8gU2+WT605x3Y
otSGuK1licit6C9yOfyZbxcKwHYk8AAWgm9hmjfrJqtPUvuN3hgvee2qpq1Ywi0hpuzYZgJicZiG
rhOktNijhNnHUVz5fWtnALx18Vn5dro6T4HAxUv6Xi0KUuZKGWnz/L/lcvLv4gcjDaITZ2JJS7cs
IImGv3owNZ/iJRq7cJKSW9R0QBr9ZhE3Q+2SdQY5310liGHGpHjsog2gcR5Eapmz9RNjcBc0kASk
uSvCXWaHuYTXGrZIxOeU1000LkdozeyjA7dtsrewiH8O0bCC5tK0JI5pY2XNV5z1Mk7eISSVAVr0
ca0M9NmmPVdrnbYN8nM/dIuWCyYDvOI5evyVRi1MD/MaSaq+PNpMpXOl1FMnTM0AeMahNY8Lrq3E
DiXy2i9Y+Evl7ovKyi0TVRSuOcoppNofRs9lf4POVWKS/2Wi1vgs+vwE/l2V0OdusbY8yG3Ratw3
kqxkvzPO1zkrx5R2UDYJore+Ai+Iy4vcm27lGsketc2E5inOtCUsqgiwcWNkTedBRa5fTTei+KGL
1DUe5td6q07Cublr+Wn6S6qT0e56Z42AAEWiOwnd1FS2/qX+n/0d5SOrkrdY4DJIPafb5p1+puR5
IxdzVy3beV2Yp63dFN1ximmVnqhBIZzoCZL1uBkHpnWJqNyM66SPqKKKrBxU7kqVPhUltB3ir32B
RRQGDmtZ1LiNZg4Czq+jEGpUwww5Y2JvN6q0wF3Q2DhYAeuMyqIsOAh0U8iusq4w2ywpvusdes2a
WrU9R2+7L1StFS0Q/0v3C6okaIC3KNRrOH/6UTR+6dEwSSQNJn27+QRTlDn09FvwSLNiRECDl/4s
TSnwYyp1cLH1VmDaU+t82hcyJFtGi9QdSosP2XUqdcm9a1pS9RNU4Itt6beRD6mfpX1eyMen6Qvq
nG/OAuCExwC17QnJm4v4lbIZ8KnPHsiIMeIYYMwlRYtMNEUVRfNnyeJD+vTU54X/yZkZhS6OONQp
mfD0Oa41549EkVkZPyuAoV47lJ3658QHdrF2x1zuMHh+m4t0JU64jSm6UTr41G9XFkgvaMS75HYi
kU7TjySloTkiLua6idH+vIF9lWtxPisok/tHjgrD/gGL+jB7VO8ZJ3NUDOd9CX9G8LHxChmRWyHU
HKaacKlmFQrpBSK24hzA9TwIiSN9weu3vHFFC6g4uttWQTquLOC44Q/HnKWaiUvJyJvjQh3JxedA
Fk4/VKvNV9v7DBmV2YubYREKKiJINszy/B+kPPGJkAMJqtoqzj0wJ4SiuZA6TFTVV7WHs+K8ErzJ
3uCGENuUoxiuWXnjUPJgPUNx+tqewAJpAJcirqnVZ+uGEQLhh0d5eRVQpMOS1cT2gFqAvOPbi3be
R9WAia+u5Qfv80uNA/hrOVZ1unasKNZPaFFExckPQ0U+8umEWmD3HRbZtsURSMSpS6qzunbUrHMb
kZS7fAUF5Ryo1c+jqxVQiD9Ro4Ld0D5O5JNi4hAG9KwoPjmD7L/GJAGa2Z2feVe9UbHtUtyFO1df
2haSJjGUZFcI41xevRcuPuS9rXM386yWMG0feI71dspB+tA8Cy03d5KYyTgoHTqAqzjjYDaHuepr
jAjXHk2kqqdsU+RlX2i0KmI6ep9QZo6nVONXlxDkjBCqb4KCqCO8Jonvu0w190wpG4sdGejXwEpn
wvxbLT93psYca2a0cxdEoHPkqzdUHAjwvfJgm/ujaf5Y6Ky/Uv4alURV7fad1IX/ociHRRhA1V1y
fLzUYD0KK75ZpWofLLQJaxFnv0iIwXUfkk5l7tsG7xDTeArV+sVTDqY3GCOM8H8mFt1kUzrNtzO1
eNgKqNn64bbVYNpPgLAbC//qQlMpmfnh6AiIxmSclwpPFykqPWoaAJ9oTi+rqoQ8zK/n7aWLkEOq
kIvkc2zcyNXRw1b5EzSzzW0HZxnZGbgxMhdqEf4LWNaGUKxK15TpqT7kf+OfbBv0YkaGJWwg9BEP
4zgYigik+0YSZdg2zC5IuUb5QQm1NPepSLsb0uDEhyHi2zX7K5SY4WDqrhp5/lEf/NlDC1E70nvH
M6JsN4olbqB/NBHISEIqZ1lVfFHvjixTe1W/24PolpZj6Fd/3Vl/SIevx65ghWzH5ALYLQ/Z4Y/z
Zem6bxaFIgVsoCpjxgt7ziIQAsH/O5UjGIhtc+vnBbzSlgYVsQX4CJZTEZLLrtRM3EdlswM1HhRk
ssa/wWhxhvYq41QLhNB4LV/6XuV92oU1BUzOlDHXv+RELK1Zi74dW93PKS/5LrZFooK2kAu+PW9x
B0jRvBn8nB93eoRX5OBw1IzMLx7lM/YcO0RahIbSBBbPUCG9NCLsF2UspJFZhoVlj8AutRzI9Plc
pFNKMDjW0AdHiqzYIZ1WVkzjDtWD/FVMIm7GmgxKNkAA+t4BTWo2khR8yYDWGMw3n4jVKHrItTxt
v0t44QGzEoSdJE93FcLRju3UCB/WVZxFLpqZa15SNjrxHSM2gxXQqedzgGff0n/J9rE3Bu2d+MZw
WfFlTvQ/x/4GhSWw8aX7njNyPzBc0KjWgCumOrwihQYR4QNrab2/UyFkY3RxwUm59I1GwxbTMSHI
nR5QrF1gN7CnQYMfN2najQL4KYpdsNeUNCwIuwkrTqpFtQOTZTrO5wFM056b7bJKrRen15R4Fo37
w6OFAaf1DQsYn9f2P9iRBeLtNZRmUOgGGnrStmONDUmUTM2qoBgQ2xu5HdZuHnMFtljXRA5okg8u
MbtS9SEmRzI/x52R2o4Y5NGk4g5+3ei3WOfi65csyBwWVNB5w6YT+4T3Q+lWYAQuycFehrP/QcJ9
FxrppQFp67NzyMAyIaCYYLxCE95+cYadZKUQxRYTTRrtgFsQ6rYWl8opAW1BlGLMNLncnpq36doc
X7A6CSHODwk7csyeVvwEqe3Ekv1eNXgjy/E/oWPSDjp+SdCI7UZ5cU/0Cn4/NcC88ZQrqRKu6Zek
T8CnKuzLIespS70XVG46XabNhY00I0Y/tmtfOaFQGmHZ2vtyh7sXc9g3TK9hBdVvNeGLfnSF/GNL
PxxcXQGy1OhM+PpFHwehP6mnbYuRdQ8z674J/JBnnU8gJ46dGPSL723Ahfetkp3GYwguYgxO58DC
JFaEPVIyzTyQNT2AVJthjeyt6rDM0A0oncCj8Nu8cCkVeR10CXeeISnkr/WDUqB4c4jiOQ4oKfbO
EbNIdh9gIClvIoxcrFgzj0r4KC8takAoTOQa6rrDqBdV9nGxAjflT9ag5iWMkX41U6HdyDX37bDA
CXQ6X2cNZNK1uoTlavvD3FNR4ZxaZ8vCLNWrADpuNym259wrKhdPTljTpSZ+bqr5T1QZJxhnr10l
nh1iAQuPjze93dSKWbOmHzx/b6hpudAfZVLnP3mwQdbXLVxnBRi8CayLvdMSgIGtiQ/JHualH4h6
sHn8xo34RjtI+Wu4wBOYx/JGszsAHvcrNU8DeZG/z6LepsRBHZRR96K1FwLUZf0jXjM1eTmPFQ56
yUbzoHm7terfwCBPUfikpC23Soi35vYHwPjrHsRZ9Jrl05lM9X8Va89dDVd0mgkPFGvyvHDp6wCh
bbfbqGyVB/Xi7bVk1Vvfz3ObmoOSUFE5u50ioYXBCuUAUiXul8HeJES9EUwDA3/dyFDc0DZGIyCg
Jr4mBBuZ5HtmU74rjRohNhtw4og2vKTjcunLxDqJBecF4I6eonmfsjagUbDZ6Q267CNZ11f5rLQ8
VDFxK1InOG0dfxd1ZfSid0tRZLfKlIBuPFUVX4PWzoPLsmxoor1++D0kgB00r7fd/fq2IgfIMtOF
XrpakXEHCkV9jmFx2TxDzmkUOHMd+B+Ef8gj6tc4ZWmHXxGFb6CivI1ScksisRYV09ybB6rXXLQi
XIvOyosczI0LiFTe20QQmmQUjFU49cc6Qb9KJV/3I0NeHOtl8Tw8xqRR/v1V6pUEuXyh5N1rYjjp
uELL/R63QoUj1OSGdYlm924xv5GwHNWOBvqTtqANIieSvNyX4ijmINVe7RG7dMcjSBojqrdATRg+
cIAAvbArwVcOjKLDvVRbFy020DkEw+kNa4OrVGGUHPI6W13qIE2aWbXj2u4NdUBSCV3KetX6U439
bar1qlMUBBWev4zGf3DuWGEtsvTpAF6v/LJX2wiZMG+8FrBhek45JuVzwjkgz6L9bvQL7UG1vzIw
4zU0YOVAJU/Zbsomx19+S2Czz96X+NzjSU1KLnwSicGC6NiUJTDYSK7oHuSMeeZ68QqQWxGVWHdB
E6bYFz+lF10iA9LhaprYIsVJmTPT4vjpviu3NvrTORnwWayjMfG4QLFsVKXbs0CsOJjFGAoYOtvH
Dug5cR/lDGh81ugpKZqecTOxDghniJkV7zoASJQKB/WqziFcZn6BgJsulIoPHno+xipPjjn17ZmB
tx6uBpdCcJXceRgeOxhhll4AA1tMUaPeQz7eCAqs496IoJtLnZEtE46c4F0ojbVZ10ASHmIS7lC+
oUUExwjBUtb4JblfmTjcQsIL8un+ekGszSZfQw+v05VyD5h1RaHy9BiDO9Z2+czUCgc9lsjAW4jF
7S1KP09RpDYfKlXReOmJrIib5kay2gXuTkFL/dB/lf+/vqSEAV92auHX8WEv/MSCCClbX6ytI9SE
zpQnigLGZps6HmDKOh4x5UIAZuxEqup8voQyZtmZxwolO+AgEIKLgp3GUGI+iRgAjsisabfzHH4P
Z3q+WYupxUB8zVMA0V7dzph8HvW28Tlq1kbPAyIfV6BQClu0JTx1EEqw8dGiLumTohdoBQdHSO4i
smBabwIYXO8cqIOezPE6TSC6kmD3H6Ad4N13lgSa7sjtvIkkbMSqYanMaGeTvpbo94Rexhi9kYAu
Ei3sXTfjAK5aj4K5yvtUl1cYbSMGchnzEk8Qudu79GNzu3C0b4EIwHjicAuy/Nru11qSgsMOJ2Nd
5zpQvOz2jM8E7FY+ptvRM70/qcyzvivLrnP2XkWbx7rqg9pE2O2jCpAnDlTHOSMjeNAizcuu3sTB
tZvgIkBREhWdE7vqqfwNyEPhQ8vSSOTh5H6uE0B45F0GjMBWa1pbgT2qsOfaZd21zQM85WJQgF9M
tySWTe2z7hKrDujvTymyN/QpmTBdWo7KpGI8nqK6/p6+lnNFHO0wObPk5K4kuH/tKJ3rNtTApdyp
6q/Qf6f+E65l+u2jP1JEnMqL4wxjdQuw7VOos7wsz7BpRQGeQ7gJ+mYm4L45ilLtaMKvOKKHcWjD
HyuN9jJbJrGvsQRQI6YgOjaaE1g2trECbScFvQzOsCk08JtkkMwcqYE1OKto5kMH7anjAcWyBbX6
afOnQlYRlopEuK3ij8mv/QWHRaIAIYP8E2vBM8laHFxm3GCuq+ek0new03yNeHGOr1QffZSNZydK
dQsr//jCUiWM3OlaN5Ek4mIQHNOHaIfepncsq8iG2L41TrqDB4j0l43BuKM4VDSPlHCpK2wVjP+y
uKU+1vfwQFwdXfJhVUFuaG0tJwO1kGX8i70OvqjBWF4wPU6isA2dcosXbGDQfBAJ5j9fW7Cir9yQ
0WfWpBB81Hy32pjzqPlA2DsI8M94dI4CzhwxODdmELnckYM6yXEA8pChJ278pUzfgNLOpvSIwY9X
y875s53sATvA9mBjf80+pHyT4tO0OLBw3chgsUhE4ymVyA+BpoWyf6GMmt2zdwElIHEQCPujmv4M
O/6Vn++S7dAPdKt9ziSVSiIwLgNqHC40KxwjHT0bOyhUhopqcEEl7l0+Eba738mlSE/uGN7IUJpE
Qv4w1YURrXqWADhrrR282nUuOTwC5PCIbPom1jf0K7B6l/+9UJEHQB2G1daEzrthe7v2FXX+fehG
kdyZOJAdat4pzwnkstiO7J4NjR2xv/dI9uVJrmYuHAS2FcTzTXQs8/NgeGiQ8YxY7F0vWLxWSvx6
ylFf5K6TlWDPQWgX3nIIXdL27bPFw20RFeSBuGLpY9nwShho0D9/uL+o2QItvqCv0f66aMxctFLz
NO2g1KnYWCFlv9chx8truCZZzpA5pmGFS8wK9Sd7TdgGU7Aa8AiWb4UJ5OxI5i8GOudj9L5D2Rjx
lgciJNhgvFwSwJeb4o6Ws77cV6VjwSbJIscSap0vJ4X4G++tgmIStH4QcC7XNIUqoc2SZVoLxN3v
CP8YeR529SifpntCmxAtM/K+uJY4OFPzYM4SnnTEnjoHfB8s/wqBYG4XtrSzGsQcwlx4SW2X3ZRa
ohI68DaukNou3ZJpXbJtAzaiio7XssBQ6CLR99L7fd21BjIDm1OLYcuQy/oE8/OxmiMI32dvoTCl
9nmcy/kiXPRkV0j+bWp1NUvtzgxr4ax9f5AsRymHX0yy4AK4tAy5vwLK8HA/6pe5w/HUufkbOHku
7beYxpL56O5LjXN/iAQyT7rR5lUUOJizFs2kwQeCFRLn11I/o5DsORCJfN8t5WlUQ+qNhSVh/H8m
kkcETcdX/mThC/70KLLjssttA1hsjxurrI19O65MnQ5PK1zZHezmhualeBy0CBrBvkQBSo3LX+HR
Es+wkJw27n5v4eg6BW22Hx6b7gNzpyEatwuPZHV84zsBdxqI1DYw79DgqbanTJ/+y1C4efj2DBaS
t+LSWRUqvqBP7tbLTSV2BSEbcJAOYtVYu/BNfxPLYX2LSNOlYRSmo+Boc6etebBmrk/tfbhvTA54
J53C0fQNf2v69/60eLjkYfNd/ErO0gV1xV4Msp8sYWbm1Em262BF/8ZVyMD9u3Lz8uTMTAm9l+Di
Sz35OvAMKoXJA5Id3IiJRrUFsNhJoMJCiKf0PmPU6b5nw7nt44LirII2wD6kW2Ea39Ks9cF5sKP0
mOdEZYhbAqxLT+c2MIZT8tw0SZ4k2Z5PI7QcA+nFcVJ6LR9XzhYEHrk0CWHNlYouFo1Vz+xr+REH
n8UwvkZxYMTM/Fpe3YCkWhCuf2mtWwVmevZjA/Lp+rGxP6Ct6q+bDI2TYTf7TaPnmY22ap1aM5S/
Sy0GmKRiIkX0NE9JCv7A9eJz/nPj49CRIudSpOOLrMDFjvGCLV3QLLRldw3UyD/nYqqbuOPQGw/s
JOV6LzJ2/uYwXDPesVEzKqTnJHnySkCj1+jYfAIBPKgmduX8eGOK3pmPJOWyy6GnuUF6aBp3s+ka
IMY92lWpLA2kOdMi27x6kYoCcV1VQEU3ExNTmoE7gH36JAihybGuo4WPVCtGsa+jEThX9zW+tt3J
bmpIbLWsHpAmJvvOo3YIV56J2d9E69EuTPBu/bb3JTtUMys9mLrAe/t/K+alTpVm4uV+Ktab8iwT
dGvCUWLw07sQ0vtn5GvtueD1wYWgZJ97geK1PpQOl2n916qzn+F8JMTQPsjRJcUSY4bf7G9ieY2+
fxN9n4kU3as0fywfO1nDYPyaoH+6sD14MeZ1kC3BnpwomHBxRZXnzVqFZVvimu5QvbvnuDH6XeL6
P6DYFLR3Fy+nUH+x5gGeavxc6hAxzMNK7aLitsbz5gQLVYi4OkuIs8fwJpYiu3mme7yfPSJdv9Zl
Z29YH/urW44JeINiEo9hcgH2KwHAvfLFXpl0Iisp/AOIga8FWBhFsCvN63UJohdONpbEwa2R0dsF
pdMyyVsvF25hJeyMIiriTpDFEM7/pzyW680JLPlSWkkAyYI6XOryTjoOin5Zecm9roBmnGCLsL9S
EmI3x/8/5tk9X21RFxqU1Y++1nP0r4F6zoLkfY3u4tDsArPI3jv4VfIVTAa8hcvlMZy5soXX5dxg
HhFnr8hyEZVgnlg2TlbtmT3ZGR+uZu0fGqj/OESH/7JebdPir0uSmP3C7KpjgeVrkK9xqEvm+sWE
iUhhFVLnGZ94OaOUeSAPG0iU5Amkyy0TKfdgKcBpZ1njMvZS2t+bCBOniP6M0aYet4Ni13I9FoeH
Sd3CR6+bQgtprUxPiRkjTlAnnP3B2d53Z93gPdP5Koouj5FWMGGMiv5XSMom2esgup8Hk7DK5/U8
zSWfmXO44mi++RisN0X/f3MO+uZ1bDe3CsT3S06L4o01kfWSSLWF79oxVDbHRphJcZefAjxX4QSH
pC9FTzX64OmsU8LKsHIwcNXqPb3CGnAnZxLvAXrbCPOpKKD1zA/mfVienkEj9cN8e1Zt1ERHYV1I
yrOPCR1nd+Iw5wViyTGZdSxRvwBu2DImzxZ/z/5CIVCxJRXddCcBggB+QJcvKQTzNtXavdfq+oos
dlArF7NSkZjlk9LXnyYn9AAZ8JdCe7pEAAryxhUUElJ9NzxWVMe3wriLvVFDVXLoliRY6eZjyeTR
17aBr6lFhloWCafyUICkxnVXOaMyv7KX8G4Sk2s8NDq4plO8SMu8FjQ56Cj17HA2LzFCUSXb1HBu
qjZXyGF2XwSvfdbmanFK8tZVCrSTPOuHz2viy9TWi3N3IkYpWb1a71qz4GWqYD8b/nwwrUWS67EN
Gxf2Tg==
`protect end_protected

