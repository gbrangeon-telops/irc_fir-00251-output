

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
XZtM4bLmkglBewlWavfkobXOIMkrnElgJo+k4jE78ykb7oIZp/SGV6Fmfr/ogrusY/kHxxmgAde8
wVKEHfi+cw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Qj5OXRmuDbyb7tXOe/IIP9hVzpHdYEdnGFMGPum5TPAz9WJzfNr2HnR7yYGe719tx6wYAvdRlfH7
1KYaZqML4WollrpclochLq72pgPwbtC9iEEWlamVuKdvYSw0+IzNRBHdKqTykxKbBvXaQ7+UOUjw
UnhOWIyi6vA2XCWBMhs=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
wc/9BtL9LkvfKqZJg7KOk8nPkSL5jxvAGfC0RV814LDUHBZcOVMBTQdouKf45+uYbzuqQuzhrFia
FyTrOU0b+Dpp/D8a4O6aOPezhZlqDF7SuDaIsbNJNkVeEPTzKN3+pib+HJ+07zD5sgOQyBLQtobI
4fQy7ggQ0o0bOrWPzlXO7kD45yraaLu2CaLqYlQzcDjqnvaWtdvg8Q6aRiloz0plB7OdNZ9a1tRM
Nl6v3ocdKRatScwi+YnBgJn5ewXMvGYuuBOXAkUmcc+AFWML9u7RnCLEmrft5oAR19N3inWP9hTR
9sdW8LGJ406SdzZiv/gZpUV5t/AFjTB8Nihgew==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
RuHNUBMTP+a4VfkYIP3nKug+Q6Ygohn4DcPwrCybnrM/u1NLZNct3nJM51Ftp2uYn4LtBCAEFd4j
J1ykZQnUjNHc8Om8TkpAk8Xoe4lNd9c07VFQ/PdNEPsRZobFbRhtaTn5kYtwFZszGT2+NVjW60i2
zzHWmeNAYn4vMcnLRnc=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
M1UhZ+OMYDjkT/STr81dVx9PmVVG5A+2IqAmn0405vupx6bbRZIy5mB6w+gLHolhJXN5SjXXAhWo
hTPhhYqRE6WXBSt+aNme9SGwhhYQCQHfdP7l6de6Oriyjp0GyOVTMXW7th225i4gd1/MFzrJY7uC
eTxBA69zF+OCz0UpsBa0iiqA6SmkbUtST66y3rCQ2iRlo3MqgxqTXadwVQPjyKh+YrZv8hSoGQfZ
859BObwRsVOuARh2h2mJuicqAywYo8mWCsE9MJAhCYkJvjGEbdjUCSpq6KjZZuBtdg5UMkBgdSnW
7odTSYiZWcCz00u/B4xtOP+tFTZhOrGrUTKipA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 81744)
`protect data_block
kh6dcHG7LSstmrBbnV9bKEmFDuuowh3YYtpVpPcQw/CqYla+CZUQ7VzbaJ5B9Ue61ODuDxRBnuQc
LO+zCSfs8CRwsezRtoerPZYF8FQGxuoR/4MldUqPrA27X4xiFRYtx23+p2XlnSmsu0LDbtTbU7vZ
3B0zPnmhulFw0ccaZhTZhHNhA7qcwGCdaUpqYpcZCd93r6K4zLgmyR+YuQ9K6lXjIM7/W/H/drxy
PG85JggM3OYYvZrvOS4VbheTxcdkRPsib6BBKBdbVe59zXpEEiFJiKLeWXz+xFqTaX0pk7Jbp39h
8zAz+ge+xyNmws72f7oIR2x4dzLp+TLXJX19io4iJfp0JBNx0IRoGB8Y+o9bJ/bedKdJ7IpoPAlr
H7WQpMGm9W6waatIUV6ur7ySNrIeAIDzyl7uBwvqwSSO5eGWzkPr6K848eRn7e4NKSzcciIkdkrr
eZvqyGhhKp+J+4J0YxgwkNmMW8YLKlJJtUeJmcyKHadaZhojcIpVJZxxgLPFdrlzi8sbyJ/L+E4Y
g0LhlYYp+khCoxA/SPN+mBpCWagkpUgvWdq2l0TrfkAG7sAHi8boYi65Aa1ySJDMjB2V1qCWSsnU
XFrGkHMqg/BQyMssll6rFec1VWtG2ef7BCZlk5mYvumAmoEzy462lFSI62eyQyyKYj5hXhpYa3fJ
xkqVglCUeHcIXcozrK5E/j15meTDKFAeVULSHewylfCrkp/XFATY8e7txuE/jQ6ZboztjQTYwuIY
XAm5kLgx29C9zxdbyE67HDsNxMq2bq0UlvxhUz2RDsMwrEVvVmFQWTl7hraeqJoOzn0WGhz9MF4/
hQCXnjLGO6qOenXbk9WfGxIDU8l/RVV5K7KrMiXVDAd4naWpT9t4mG1f1OIJyfNljqFzq5YNDJBt
kInj6huTLpxJilbfMjmu3ieMv26eKEfO9IuY0Dl8tTEHl1eUUfDPyIpQVTQNaEaxPZhPd7KtliDZ
YTweW/Ang2rALrHPL0yyTb6/OkrLroBLzkKmSRlcam0/NZnOQm531tUGy2HR+5cYMAb2Y2FUWLGN
Vo+QRiXz2txsGeioCu1B91nru6adLcC7k/t5YdNusbh5CbAOeEdN5GFj1L37dsZgARmhxuGopiEC
ZVn97QFo/ElQnqzw0ocCaJP3Dwt5iVSZ3BOf4STEj5ImLy1uj7NEU4q6MZVXOABWL8YmOczxppLE
TEqPCW1+CEqkjFIjoMm9q0G7CYaA4eoLIQdg85KZpvIHA2rqdS7+ST7cP1m7BHe0ouodFfT4gXHC
tcVXCiGkrzod7j5TAvX3u/kCNPvvnIeqHdRYaT1c/evzEZpo4NUmfqGo4vfig/eTrg4cM+PuQ0q4
ORIPeci7vq9Px1kosutfh2sH4RDRalcEPXRL+fldPxmT6qYPDqo4Dsmi04II8EEWTUsk08r30f2E
XwY0nL4jn67Qm+tUpv0tyxi4OwKX6LlaSJcKnuuoLyGvKLJAqfY0FeQk9Tu4ZeK2C+JPb3IHPKRm
VtASqWU8O9H+7s7RXjTvkIl1KxycBdiLdI2AH2ek7L8mCcvF8Juz/hXNdsGFvnfZOs0tI6m3KbiG
a4MBi+aEq256oGhIzBL+H8mniDN0rvi1gITiM177v+m0gEEC9B5F5iP1zCVJUFmrwlT+Cm6reZp+
Ij6D6K8d1qz1wnv4IZdu9lH3XLNy1lY8qXbARjazqno4wzHLDvXSsfNPP3NxbrtpsMx0j7r+wXyK
Cj3RXjoMAdj9XS9t/5wf/iZJyBqyqeJdLy4yhyk47tH7jSB95Cwc9bq4JdgUtdflrEjx8m1d0BiJ
SzdS2S/3/r7FUAnNghgFsY9s1dcDlAKMJI/Q7i/GE5PoHC+X9yM7YC+TQveWXv92b/TSWkm/GZBU
Aco7AzA2rUjqSRYvAgDb5kYz2AkFjQjdE5CZKPDCt6zV8PcFes/4CMQlNN4mGzfNl0II7pwmEluH
uSzyuwTqLfZ17+E18lyrRIxY9gMucbMmmNFTqUZQBBrBeKhKHm905HfCUR9LnSh6/yvrCRGGsuWN
GEKMs8QGfRSQ6XU5M82Fib7d2bBIIJ8TvUy3UsXqJ9crsXB3bh2cLhMxOgQf6Fl+t29pnty6plFN
TX1kHr5spo2MCRajc9fqLZptiYZAwEueOSjhYWLZ184p+Sxax2+LHaGS7X4W6Xe9wTWOdF3RESst
P/BLWlRYtzGxUUds6fcoUw6/225zcijcobzk6pIC4JEpKSBt6sFDaodnlgfwVe27bd3R5hgeS6J9
ILt/FOUJZnYA0IAKYdGKY7Kk1nz+UC6P7wnbHqV4fjle0bbi9jncrt8LmvXg1sY8RRFOC/eObofo
tijpsGcFg6jpxiJPZ3Flx6GjBiGbxkjdYTu3XCJE7Xw0Xu9RYqoFMKYvnyXi81zuETc79BTLsN0w
h7XgVvsVjQxY51ZxCKSHFf477Xz7yMwSQ/pNvao7By5x+573tn7sutpe3+On5WnnKQRurS9feFGx
2iatI/fnAr6VkWRxswlYZviKZKxl82zuM7khxEwa3P65solVKPOSFX9Wx+J5sTZzKRsuoWcZFtQi
jw05XI7auSpo4kkwb3HrdlLjY+zNCmUcG1S134DL5jCtbT2sDb5leflQ2HQEaWwZe2MifB9w0ZMk
8nutpTJIsaP5b2eJ+lKhXA/ahtlrG7V9mBWIG6f4IfP91WN21BgXp7EvcF/Dkw5kszw8X2yD83Uw
nmpUx2t0zo7DTkjvNHbih2NyncR4rueX9nAbAvm814PH8uktSq6MRqyFVavKCzeFne008bqHt2Nj
SgnNKYG+Wb1OieGArGJCDpVboEo6Stah7G1AWA5K8x55Kc47nR00Y8DMaZGlIrPh1TNWbmHQ6SMq
XflrlP9uflRppowINOnzYCHEYNHeDOzeRBeCPf/X5rV+AuehnMZhdSh10GOLuzUOUMaZ4orIvrDN
65mluIjsMxxbWmbYWl/PxLEQmBuSeLdL4PYnHNIN9ZRh6vzeOeGXMkfUroTvuv2ipVAM3yqHOKEz
n5Mczk/a3oeYorrd9C8Sj8g9oXL+sXsSIStASDUP3zxgxtUsDK/6d+M19fPrfvAf+9t7EbOATtCN
HJSQGJpN7Y2CqOgzAIhCfGXAVC8Iw9dT4zM6H07L1ARhuetUisjwukLsLH5FoHzBq3M4pzB9foPH
4nOcsrlX1xV4Jax/I5GBw5Q4QuY22hqFb1HxPP+bMAS6sFLISGzVpoJJjWtfvnX27hkT/SkK+jqz
oL4sHpFpIufac+gXa3pXiy4p5FDlWGYUbcc4O9Tiqyw9+qHKZnx2jSUHhvd00TRXlFcwzmA5cGTs
Fmi/FfSBYHVgLQNAivFubgpN9wRWeCv7BEgZ3C7rG+OUHuukxas5Nz/y2MtN/Tui5zFCDexvoIAX
EkXy25j4cbYdRqnKSMsP/75+XAf5CDKMoylikGlmaKUYvrSdNIj7a3CyrGXSKdPulo6oIgUyPGXX
uREtKYexzg3e7fBu0HbBzEPHUL9/8JwZZwTLfmPv+ygOF6KdDm8iLAol9nPjcqUSs8lv2REDeATh
D56Wc3MGpJdY00z5kRofvHEJLLAzIpRzjRNDoOd4/4jKF/lOzDDyijGUvjjHFSJf36DK0+epJmDn
Mrxr79tcqSTqdxVW1qoVKF4QAVIFey1nUL6JYdxCzm2W7qK/cND4KgU2P2ZzCuNQy3I89kX2YDlT
TISgjaFyRc+p9LKJtftxoi20JWitMJ+7odSjGzl0PieS9WvqG9uhHprtBTOWmCMl7Ib/2JNoaUc+
xF5H1XoF9+lricm5xMdE9vBVXsaxqLrfk4bdxYJ7/IzoWr673yi+msvkNC0ZZt6nGJjd8PFN3l6w
s8ddOSjzM4mxYAyTA+7aiM42WUdRzSCDNlijBtN3a5OFXKqUFA4hFAmmWP3sJMyyuYcLgCLsLqJa
HKjLHrh5U1ITaKn1+G7Vfh9zb2KghuhH4s3d1PK/suEiMXUXpscCovag71rIRX1v7cJHpBIvCr7g
vgwfDt4N9z1KReb5QP62awVGWBUC9YPQDUjdG+ECbIxEewyS/dLwviZ2s2fnFhhkXzKzMTlhc3X8
5vZKBQrNFst3/0D7t2AEimVLleT2SlaXMUjiDaZ7SBqp/kBGZ/EC+CLKCpbALq+PcpTAbQiLyQyo
GCXn6imSX74fk/wxYlA0Q1rQvm1VIqxdQjnJMBELglr3LKPS37TYDexRjFWa1CfKqps/Pb5VwWvh
vP+Em2QoZiGhbUICxWVl1N52L2VSar1w6S+4YqBruPxKmcPzlAjOsbFJf9ibPjzv26KgRwZ/s/oI
9b8fLUvOgHA7lu9UcxqzIEV5Y4UbINhbnV4ZT/ZaoV20PSdPuAF0UYKwjYxyZh/wzbrzER9AKUR/
+/qWqgCs5h5xQH30v1rTYaGofPsCFOj+cxioAIcPbNrgsRu4kjTIoitkLPV+tIf/NuVh9+6SwVZi
oLc+xbaM2DiTwpVX+zIQS4T3surqeO+qKZlc87d/yUFQ8ypFcjrUI5bKVNmjVPMLKcMGW98Yr/nR
KneD/l7+nQ5qlVvh37NFoFHX3XDH2UGNgZSpaZdWWy5qmXdBGr93XxF4I1Fwm5fKSPwnT/ZhPdvV
5M3fPM+NMakLm9SYaA1rolSH/5fVISofWJ/0CapSP31RkLedIN+wMH7h9Ty/PnZE7fSeereJg+7F
uH1UzDeWsbDYcHOdVxW677hHqdLtpt4MKnqHQHjYy5Iz0wSq2Wpdn1alPJ+AbNpNlJR/e6T1yPwe
x3dQ8qPn1yiCHKNVHx+xEMGB6Ke89fKU/LnS/myly48Cso+8a2yr7ho4o8ONkDmcOgf022Nt+jbB
i+x7D7sFpMm/d+APkOMxuLOcVkZkSjlfynOJMmO6xM4F7SjMoSVJU8CIF4Mifj8Q6uQQUt+Oqeo6
3dCqXeHK4FpGqn76SMbaO2GQhI/YSxDTwsDHlPJlNerNpvzFUdg5ukMdc3v2MifUB05C73RE2czW
H+k/5l5f3J4o9fK158SZy2+zKWJMfUBdCjnuJHQjU65PDjAgULtaxhOaylStz3k2/y/f6kJPFlSr
5OeKVNFPQATIToeLPoOpdKL1QRELKTtuYK6S/iZXcD7LMedUrnDawHBPOybNlfRpDLifuNUEWSPz
q5yilV/Mo4PeJ+nFrOrk6eLm0G00pPIGBUVFm2pFVrjO5AKqBI1eBfYmvTeLO2G7CSS03MTDosKT
0dbJ8kO/g4MYqw/25mTMYH1hI/4EdjbTgeAZhF21utWR9t1cxVWeaITHxrVZOYCKUEIqCOp+OuBN
Hjp6QdrtB/W7KuuGiEVKcMViewqUkj6ci3c9Rrw6o82maFCge3R/ppwsYkD+BAUxLEnvLSYUc4R7
5BfT9/mjah9Pnq3t+Q56O0+JWHYHmPWJLMNAdBdui3GlwM9BlQMDsPDcVZ9Pp6xi380UPN3Im7Uj
k8UIU2GLrfQ7TPqRVLKfdQX0WrW1rTXlI1hBI24ufazibOWayOOXnUKmL5xB/MQUurHo2y4Su3qh
YUgF5VFGu4jKek85KESmrJa30qMHfREOQwW/A8AwcRMa6xEd+n8HJCpBnq584/vYFVbHNvjxagkf
F43Gje1RklRHhfIh5OMHvmTiNc8Eit6fVM0xAWl2Yi7R/Unvr/pVRi2vrX++Hfg+hPH8grnLga4S
GMZed3axMLDzYT4rSerbV+38Tv5uLlVcMjl1ldc96LxGANIPf3UIv2ax2yknW9yqFhEOXUlnxTqZ
TnHruzmT0VFGov+h2nY1P+GQpTJszjQUhWfsyGn1pbPIdtPNTgkr0XnKTvZgi17U+H4IeotsK5DB
D3t1WxuDjxo7s197WbgV1A6BYz1A1vFcQH6foE7jvytcKX0Lz7wqL7AhD7EOQREtenfefi5hON/l
h6ynUWsaQ2PrnWQ0KPDFQu9GjCTRtZn+rkfetcwNCCQQ7rP1QvQndrdMUXB9ekaUUc17V1/6+BKz
/SWEWVJsdSrlc1djR0ZHNUB5gqCWnz7ZkURYjuIlK4e1AhoPu7XBXF0j3yVvtnHCnAn8YqgfVoee
HMbGhcXVWAB/CPtKtcQHgtlKSEcpZatNbgT7CJgfVHS7hEGCv0mWQaJdAgVOLTKo2F617fqRX7cW
z9xeOmKUeV68tp6E9ac7Y9Lxr2YZXm1kh8oDDQjLh5BsVM1tM7FhPtlAqAMDTdGduAmMRsFpohap
x9F6UKBZzt+cG2u2HiiQm0MJinJkNa1ynQrAyAvtG6vyp+W+jfhxSLaB4fFDoPhIV3fQ/LZbsVUI
vPn6+j6W6xQu92tUpO/6aEvWZT441TgnQAGyB3TRwyOktPiTy91m3QhlwR9qLBqv3I7E+YJiQOHO
ZtHx4unu9+6wzusfIauqJ/7eCl20rveEXjnWplXmRlfqKyv5hqpZBWeUSdGhIZz2bisbgdm6qfWx
147qyn/qAqsQOKFPVAc6axD4tVJPZjJTrFuvSU8rMckOtHZQz4aO6vE/4nVWxuWS4ATovdrmCjzr
iqIgiD9jJUVPON3fR865dm0DL0qFZL5IR73EwRD6+SR7r8laPynu6zHYqMTNOG4LeGZFPbobcsR0
0aotZ2jYQNQZ42pKhNyOCoPzgdw2YET6uolcsdE473yxEsyH7MQSd2yD9O4aOfV6h547qSxX+WDq
B5iNyoKOLXiJuHOgHSzOn4XTXIHcWniKhdiyTz4LuGlcBWfhqeepyN1OmSp4j84WuZkezGW0JzGS
8otusGaLup3H1p9uVHOcTu7dqeyZZZr5OhjdhFClXF4oMgjJW+53GtmPsrtM25+tRGmNDHZUA5/r
EzG3d0deapY2ZEd0iFYngpsgJMKH67IcvpJ/MJGmKV8YdtX/RZFex7HdaNy0slCOab4OkWGqQFOn
sOLFmCnl1q6ndOj+vUFc2EOFtXBZRvrp4df0wDs1/0JH3EoQe+dPBrhr8mKPSvXotdB/m0IPhzn7
yfGn9uMnEGmq6zYXbJp0+7FtD7Bl7kTQplWanYKjBOQ064SIfeARc+NNCs1/oT9eGL5KBnjWP9vT
x6potAoAjqSgKox0EBsVI4/GP7i8g18DJB5jIyFjWBFiLWDTc4gaRSU2U2qrrCGkfDhDPfII4deC
uBHqpzxDV5+cxMmbd6aUA0c9lOMyuHsUxspjL5v6o1H09DcH3jktI+1EH1TQLsT9fjhdtrT/n6JU
4Fk4Ew6HnqY4Dm/xdXLHGJpMhQX67aydMPNoKKqW9RNcJdfvZVt62AUhMtwn3YeQFGt9IB+Ryuhn
50WcrX56UFhXvs+CLEePM9gol+kH0NuHxexjkhckIQFaJrKAXjG1xQYwtHkLocbUxMKiljXw21rG
X8n4emqhASvvZ1JF5clifxX39tdn4zNTcSRkMwwGiksCw+PaHLZ5pO3F9dDbx6TJ5AyZUVmIUTKJ
KAbshPt1qt3Ms40GdYJAP6HpLQOnIFkr/1eAcjwpbsZ8wtWEph7ZZUVnIYhNB4rXKs8dt6Ott3M4
/9xj3HiIiZsRKWwn1hOLKyLciwuGnp6/WseHtfUt1Hx6riRMYoz2t4qzyJFZkQaJvureXUG7+i0B
w64tpBnYxO+bMEaR2DOKrqmT3M2yqOsvk4lqsK9a+bqWEq5dhOejxNmgkBh5DUcbtNZUsptLt6Hz
vrKstFebHSdL89Inzb32M3qTikHLPdsdDkQ2cZOZXPV7nknjFfMIGGbqDruz/48qCExdt9ujp94F
oViBkU7Cd1BHUxBMfP5x+QL6gcqtSxZsbhgUDs27kDeokGg4OKjmVfpulCwdx+jhX8FxbQGB36Ar
4VunmcnmzVxYD7KE10voO+CAlXcVOqKPCln7cAtszeiSkwOzW202W3n5AAOIAw2WTu29TK9/VDbR
dj3brT3bbE0dXO5T+RPL/4FLJUdfrvMX9cUwUXn5hSAZBEBlcC2dztqz1t8EojZ7D9jIrnt0dd+P
++uWRj2cFpvyUKvvx20QveRAv6o3+9DxJ3k+c2Yc4037M0lV80TRhZvRv868qnXW9mK56S/NJRQm
E8zBULGnVFKJcRBM/HfWsKM+K5VhJ35KLmezzonW8eXGfkINXbK46D62PTJAM2uPfWlanHcuqsdY
baZMrVkkJQ6Y99ltoAy1ZrpXoTNdIr9wTvFFQIVz2BcXiRYonBV6v0S38OvOGLlcpuglvW/KHhW8
Uxv4Xn1gkm/CWKhjnToOuOul2JwrDYFClKIt2njhi21w0XhUbbvoQa3J04k0CJslaDJ0cw5Yl/l7
vyy+x7kewInlKlbe3OU38NgClwcb516Rb3djOrIH3lnss0sZxUC/8r2wDHYkYphXisPsXiDHo0ao
aOmq8zfC05vryFRnH8GIDXTRB43MaNGems4qIs1lNLRyzXCj0n159AMjqZwMACaEvqzA/Hj757ia
5myBp+IBA8D7jXOexXcx4R064BaeSanpnSzWz48EooUwXc4Y+52QZozTzVkvhte3vXvOByEadT3p
xCiep6SRwz5UsZEeUZcNh35akSef6PfoYypy5w7Uq59ZYE//x2jz756JA5KBM7AGOzmaXRtPb3Rs
mE+dCSTnlKoQ5x+imrAqF7/5rSCh5Q1spg/Nt0qKw30/9S/64MCYcMsyA8YM2s+wxt/hVb6XJNI3
XL7r02KEStIbKoPkUdSvqnZYLiVs/EVwbWVYHUIYLUAkxCDAGKahk3qM5cbSbIlxLiof+3+jPAoh
T0zS0HnQU0TqxoiPLNRpUaSbHJJ8FZ97MbOUu7v6K66Qp3gU937oMCs9YI+LfbjxpdZJFq/hGleK
x4fg+SBaSGbV3tbMiqhOW2JtDTjgvCfAE+/HUYTcoQSHNqmdsjBIqDtSyjW5JItlzIkZOnMroFJc
27QVb7l/2RJo0mGvn5pbquSeDOqsSTFMGpKrh8eD334dxiyBUdcj62EVUJru0ULeBF64dubeiIll
uTPfzABWRubY3qBlGf2c+t7p1bS+A4WKIMT7ZOaBg6QGC3Dnc8VSBALB8bF7gnuZtxJ8PHQMZcvm
DtQwVd3CgNQBcGfPs6j+l2hWwABImRcHuVbI5wGhIz3eyEoqdwIYte651RYje3mYN/JyU2HOpude
ux2xwzwKVQu9GZOwtuZ2mnkJTYu/uX08/FrLhP9eddZIRPXKbQIDxjC8H1xjqYAZrRpkAKvURw44
lL0TWCuTPUzcC2ePH/GDaon8mNL9LTXZgAi22g35zV3OQH+RDl1lpaq98mEQ600W3hEEt+Nl2qQO
d8Lw4drTpf+or9Nh2iRjbZG1ptQhSwEydjiFx5cfIf2v+j8sgUivB3kR1JnUtemHYak06GOy8ZGn
n9KOj+EWFAH+qJeKt8Jl3LvrAmqSJWBAmOOwijVQ19D54bc9T/eNSlGIJBB18FL+R1IDsdJ5LUlC
mm71jyeuVJZAvil0bYy4/cWSoAl5U3lPtJ+GGkNYD+B0qjLtfdyeiugWBYstl0jG6wkQmTK+m2ad
vUJNL0JPjvt2wiNdbSyK397HiH36Qnc2Ct2NZd6G0gCl392rWXd0urVwAP+45YHsClmurUFv7owf
bZUcKE1TrSYR8GrGAYBfz0HgmlglMfZpBrtKLQR/tZgwaDWNK0x2zr3OIIbiIYPCowEWDrRp1mDO
c5x4ySwXEJaRx1T7VdeKwWm5FjoUk9bP7E9jAsl+XPEuzvKrjnqluHiHXZcKbT9nJC9IU14ExJuz
BBbrEpsCPlWB4Tpl5LzDqIidqvpr59G7spGBUdB4+Du6DT9Q4FupH3acFrsy3UfezfGbXsRk0qHb
0xf07QNFkbBtyBEebtQG6mSad/F9wTen8TVEpKy/80xYvKvPAScWfQS9QcHt0ItKmtIbxbDhy3hH
5wCb+kfhlmAnEr74ytgyaxg+vVALBIWy0WW1lN1Q9p+8JAjYFCx3dpcPg4FvaKP43BmKWykSukQM
+QnM+hUSRuWh+DOdQ7aYZATqnY9bs3JT0Xw5YkzRK50fjlefGv7rwMn4KOTJmwD91Xpo86v3aDpd
sDBIF493NAR/e/9bZULMB/LU/heSd41mvLFY1dUimDvpphmVvZs5Dz60tRhRhOUTdKSgch35ohfJ
t9X5p8XdjT5NRzVRP5Dke13ak/iK1eBwsijg8gYfxMPKg5e+OZcrclkqy5i8bVV5mqPEi8xFR1z8
cCS+IuMT4UVYAla28UXbLW6ziG1H77Llsbz8ikFlptlBOE/CdVjMaxNHKTO8P0zWfWEGw/Ayxuyq
iIu68NW1GcO2/MTAFYClDB9/YUxWJfLM6XhRxExBxyVVHRCY09O/Hz55QthAtRFqp/GTzfZNlByO
dc3Lin2hta3p10oWsbz3Dv5dxxrX4pzwg4QRQDp4kd+T8p2v3kHa0GGlARucwrK1PfZCvcoOx9zA
AXPrK8MuRoTr3huIhu27gFndwKg5vaR2GZ2DBkr+ySsZpRJ/fCAWRClrz6aFxWGeEtWteAPPxOrf
J1LeCr+DOp7Dl245UEgJKebebo9UlcVvRKyHe9tQFNYra7RsWdcfL9Ih/QKFH1W5x0cLGEHzSXM0
a0d46VricTzqbLG2WTi1zpv3JXz6ReucAO3zqYntDO+mtmTc2nVeRJFyKnEA9BKUhECwPBf8PgGq
W5Bwdq6whBHyXtOq6fOW7zjSLjN4fjZU0yTPbRDWIpaNG9b+kMCdevvjtHH4D8Usyk7AGSAHeQMB
4g4lW1hibNJrcDvXKX4YeVu/7yNht3IbgtusGzz2YSWgne4j401AM+z06GtFXZLFNN9LdALx2IgT
66wndswEDIfx62WEfI2P6hEWpTbS5/HYXe9H3Sw+jN6/2m5n0+7WczWnH1ebmg7mb2etVhkhwlRr
KvOBbUK2y7frohjvx9DtTYt5o4uIijo4CANoe71c6c2QPgq8N8aLJWTnnxB1vnW82mYEDZ3RAL+6
YR8vHHr8goM2Utgqk0tdL8KjQ9pza8pNSw6N/pXpRKPFbO916DeK0r8FrsEa8Ztm9adNIkyuZfNe
0KDobN92g0Fw0BRkXmj8YJYF5MKw3irb1ZYB2y8nXXU1wWKMVkkAS6RvIWuvUV18dHnVinUQqzUX
eoSOQHIcwpPyb79vYBfpOQLf8mW2LLtD2KFXvt6CUCa8u8zcCPPA8E7+Aym7m+ahcgOHKb4Nk++k
wVt8CD6nLmWXThQmQVuIx/RyXMabn8V9NLGaGegKVPp/TuHeaH6U1CM6C9zCKunVJNrO0xW5KM2E
HzoIFEvk2rUfZBHYkpKNJGp4gVWmN0CEtT2vWM9vDKLu6uUDYkk1x+MqqUEDdvYujJfb7sO9Bz+K
L4JDDQqRP5QeNc2y4lpjGRRR45w7K4YqdPq77JXutBxlYeqqRCDoPrihcfh6tAxcXijL2/xDRopT
40+QCvxHPoCKQM/XExlg3F5r9aBBkoiqta7M7U7iMNCXODkJd8RMJO4UUsdOgTySbbVZ/fbWq0Ez
2XJ3puQBA3FyT8a1697l8i/CvHc8BLKNbFvYokstokAIu4MeWxBWfxZDN9SXU2YMJrT1xArQrVSb
xk3vkGHYQ0MY4bgdFyi74sJb/wkulA5btqBdI6uLJSmga4Eh1oPmWF83v5BNKeVNKxN+0UGIayGV
QLH5brD7D0/E4BLgwgKdv/xjCWntNFqVUOdNUvzUgJVe8DJ4RYgTXH61av46OSn2aTnNi37KkvQ6
DCPU0ogGA2Zo5iZUznWCX9YNbH4cWuMPN1POyEiKHdf9brwm6nm/XplRD204jDSqdb40q6UPuxVk
JZshrJ0kZd8lFYY8+eV8XRD06bJx2RDYJBU8fgJSDVa6T+2R5t2CNrOvmeXazsVbzpU6VXpuP1ca
SKZKlnexQPXw99nJY9bddAOUr2M00RmgnlXqSLWoLSBfHkqMgpEbEMkkJuCKYqVLsg2ApmAaW5vm
92ANRVoupzm7njdxXPTK6cP4cqyQVz4PYNeY4ce7H2IZ66QNzQKJXbBkxoHe2t7326ECXJJ46fIv
635PPGkDyk4Sj9wJVpBJDLF4p97XdasxdMDvuba6Ix0MwK2fu+3HyLlTIsdllL7lwpCtf21LXPxY
WCsZjaxMXqYt8ep7WRbeRscOtGfe6YP91L12bnniC8mnYezR6hhRMdFMV5T6qaWeEA9lQsnpR7it
zcuB2jIgQmoq4vgQqRmn894Y0PP+mNYmDlmAIu/l+d+fYVImeMmCylkfG8RDpVaa+2p4RV51X80U
I9bdBKudnm2xboKef0U3K2ErzFPh/su/Dn9cTPEElfQExIkzFhC604pVr8F1VXDL1ErP2EALKtnA
rhenqQNz//JRuAkjsKV6sODXe5LXtg6C4tssfiaqliJSl6nZvAgshc2HWLLyMJWo/HsPc3sgVIrs
L7/j6ZPaBp3fY41epeBlroAHZL/5yQ8KQCl+6uJSR4PakkTK8H7vVLoay3k1dztPTuntVBvng5gg
odBDoAd3XiS5HvNIYiwJtsg4Kl3vFg3RWib83fcUkJJzABtlG/e3GLimbU77PQbHQwA9VtjNFOWE
+PJWxZAchO4ELR9WxvRqSu/GJ2fHKB6Y6HIpRHUn360smgJoasNAuRrD2SqD0uXBfaDhvWtD4Sjm
gFCG7LHmpB2X2ruhq6nye5tS7N7SZemxSIR4sn8shDQgC3U1cgdVw91icE2p/pIjE4+iuZVzQlNR
QaxFNp74+UP3hvlJGBvOWtbCB8vc2U4Qr7pmNqB/sCjI74d1dhISnK3oisq4Ro58d+TJZQpjkmeQ
j2Dc3AdX2GV1NAxVPceLGzeVNuvTVvwzUGMbYSoN7agBB+Ysqjj/zTedZ4illr44JFMyjfFGJ2Eo
H0WpsghU1i19sK3Gv7J1ecjR10ja925NW4yghBcYPLK2WXikGr8tJtrRBA81W2rpVGbIDEfPI2lZ
jVBjT+jvGvZD6vHtGBAA2hsxRgPduM6KIRYSP6vL3MtNoVOC5SJ0kK20jNp/iJgudwGLJyTbRq6v
e/biwsW98bXXTZsuNb+8KrXzCUkWljwR6L/DLIoMlCozkg6jQ578QSrh1dT84etHC+6k71K9GArC
GpKBwd3tB7U2aIn4FpOx4Uli4sbY9TLZkc9ZH80y306gYBI60zUro9gTnBMT2UqskFmBmxlcKIVU
enDdNA6F9B5XlNaqmbNfmlDzRtYnQKMtI+NiIFRGshczzUL9KMyTJ1d9Pv7Fyel/L0N+cNAdQWtv
2h04ErxBKViriO2LHtjHFS7WhzmkAJBU1bT3eeGPSCSEugS2+h2R9eQNSttgeZTmv6jnvPxQhtBb
cHn/ZBY++gq2PdYnswZHPvCVP6A+hQG4Ccz0ff0C56ILc07rY6JrMrDuWgl4uFkwcL1HUuLJqBND
WK8w/0j/Vp2Ng7w+0yKc+HdAvnRkl+kgzBRuMsC1GGcmgMGFSGG5gmyKmF2ogSz5gJSKjjqk8Zy3
Yjn57Yvzfec947CA/P80wNrxGwa25+eNM0MJX7O9pU7iyq5mhas2EgCgl3AJFrs1bFK82DFaRYgf
LxDSOeB0TMUudKdbNWbAhfZVdMfpsj9IizzOZuB8eSfrDNBIDH+8Zqh+mBab/f2+wrm1Br03Jzr1
w5GQ8CALQQU+Wiw3IVneI1toPL3ryIIzTKYqOpviS0nip7HX/I26C6keju7yGfipI1KQMd/aHVST
Z0+C2tSGNWVxwumcdP8ev04gYn/7oaN5jLoC1tvQWH7q9FExi7g0vqtdHOjEPk184vnhyHwxsBIw
wiRE+YkIqTiFtKbM5au7mF25P8NABai2VRKFMTwm9zavmapcMfakku2Zs9bIOrvUntSyswOJZ9PK
ZkjNEtWXjjKLgyk318qxw1XxTqyxXM/tDeWJPfPQa76cVoC7MKyzPC1davNclFsbIOd/V87A/55Z
+c90iosz8bTCTEqTNMTDrfIQ9DzTZWUT+tJmrA7GttJKkd/pTNA+9zvvVVnZ8pge373tbw0OBnWm
XMhnpofqBgTYTZS1wkYkrRGLKXPSq2QuTlt7C+HbFQ6MbmJcZ8wg7KelioPEDuNkweup64YcKXu9
SR9/uXSd7hDDQ0vQwQWXlIiifCr5Q8gTr0Eh1/2NLAnGFtNuscwn+R2ZBHqvBJOiF4hP1hhJ7EkU
d19XcAPo+IP5Kc9dNUis362C0G0OzJ3bdZg3sxd18FJybbkaYKvgPakPZDhXaJD5hpcz42MWmysT
TkKus1AVfaMgdwb8JlBvzVZJcUb1HpsQNdQxSYGTXmGOpqABYa905qO0ZgOqX+tWWGZNrK0JUGib
20vDkoG8AlFpMeywUp2iC6NSD2JoF2AGMMrx9HX5PRWfe6YubhtnB0cZI9Tey5ar0bravntecPdJ
k5NUTc1tJX9XCAVu0rLXqqeDC7mVFgeBjDymU325ceGL+ECdeM5TqbYyV5U8t6sTdxTndlf64MfJ
khc6TlI5vvdS+8vge6e6PXrrPEcaJT15jEMzLd4v/BQYLTQESVlL2ArIK7CZgc6XLxc/JrxJPjUD
B7glOGY3ZWbn38f3J6tIZYDNpHZzC0dUlytmxIvl0WxYGcmCMf3CLZn8vJfKIA3bcBh4EWJpdbDi
MvwdCjiF0xzxKOsOfq1k6OKWJ6GeOnByWbg/6b7FF7yXfyAcmLpDl/1zXfnK02F3tgsVs7XTWjXo
QZBQdHH/qGwwCm7hJoe71tZgjmT8Gr4sC6f5dEl66EtQvakK9ScK4OipU7Lsd0naT2nZHq/MUBhq
mOz4J7YLFHwiZK3njbWPVOjJ7eZA1Y0PAMygS8+rQorEDM/xOVUO+8xh9AY2/AoT8QnqLDzC5641
oUZMhe4GZiRablpzi5MKzfF16cwF95hhrbjtEUFNKZVlv93gtij14WymwvGUaCVMaZqxbeHL38oE
LWuUULuNsAP1PZu99AbA20Y68yQ1MVm9aHchfewhMPDXwhGLqJhhif4iSHZOpH3P1x/HRk92c2vy
Z8UAhDwNeV7D3GnDjost4+3VPbmyfpJtXvplixwGhkXKAEfprVbD7PTGsuivg/itTkUbzUflTVUq
3LwrXFkZ2+JD2MfwWayQvCTkJAKLLSoeRyIXVLYx9n2UnbtFt09VX05T9ViEPljqpstZi0yz0Ip7
UQWyyn6JWjIVY+8mnc3SPG4CiuaZkybVq5xl08CS8xNaIGpphDER4XZuQC0iz48wCD4nN6CYsMmB
OYtW5FcvGLdZ/fHneuAoWfTkx17Bfi/RcULrfr0C/lQ9KDK3ISGpKUoqCX4NpuZPqEv++JKiPWFr
lx0Bqb6DQDtYQbHoPMGR8njIPpYv88IZgQCrVQwQARyLArPxaG0obrXAF6uOec5QVGYzD5iSPUfm
zBD25l6TfBVAO+XAN/ky314q50uFCSFb+XLmctpwXKeR57Nw6LkfdRkR7ZmPiewDyCl9GPB5PxLe
wsEqva7MdPj2QgWosKRq3O0K4/8wOpoSevcXXym31isJ4bU83CYFkfLzWyDZJ0TsQ+AeyjcJ/CMw
cTY25DE66BLhJPrLAUktt+wriSfsfioqNxZyRosFFuP9XJ4X0pFpR0qVVi1bWYEy8mWfOQLh7ble
X9rHXAK9UOqS/XOV/Dzm4s/7fEXlmSuSO22S/vxO/LwD8v5+jNCklBJifPfDpgw371+1okZCdCuU
rK7iT1G1QHvvgE0jhDdZUsOMD2pjpCEZFCS/VptXBodj8WdeEJWn+k9Em1f7LgNGbQGIwjpDV845
qZNG9MYcIEEqGo5ZKXVjQazEezdjg/qX7gauuQIW5kVumGlgaH1R9Hf5gX5iUZWixkr/ZbyglcGQ
Q4mZ4CO1MYOvQsKADfDqi5TEHOV6J+w07d4PjpfuPvaZhPZJlv8IgwSZEySFtKEgbXqhmYvdTqqu
Gshnl2JHnUC+UChGRuc2+zD2jFw8dPK3u/DPJssQ3Iyo1UFAuEHIDDDkGz/oaTd8i94+7KXUsr1d
7c5GUcNFnAu3raPiNEtspapZutqglLMlAhkFUoiRjuNPQ/Uz4seY45uELNGg7Je3Z9OhQs2MycfG
ZjBNRhCi5kUyCSQkcKM7dW1T6fHT/fxdQm3Ze9Hz/045gR2LYVf5UG04DiXYdVBPwrFyWyQ5PP2J
7V5tgTfZUO4pXtnphK4EAOlUcOo5p25nYRgTw4bEpwKBOutUaKcyrWKlT0+uXhU+b5bDbtPsscS+
5qnaruESZKfLja9/e0L6C5iu4jYr7z4VHd1zldYoSZAH5hJtHOricmu4MlRlPhYf6UtBffOEtR2R
GZkLSREHVD4qbywMLjgi5xiXcHUZAGL0UqttwV0Tb1/NDR+jTcBGU4vtnQxcpscKrzYrmizGXEtb
AD+VVGGa3cJxtlWdK07/bqTXkF4cLuiSH9Njugj8T0TwbQBLPNlFhzYGBtQ6Yz0mhqXrdr5zLFTy
DZL7xO10mutE177VveKN/+xuKjPdZoWXitOwd0g9K+Id8e71po5bKTJYUD52oBFrFFU4xg+82j52
B13fDDk616fhH8p5ncACGG7jn4a7D2QJI4mc8FtVLPNFra6ZCuDGJirPZ//agrDxTjb9w3WtG077
FRfaeKd6XRpuIUX3cKQvZRVU7JliEgW6x0pMz/1MWVggTVGWkC8+fT/Zbfej21pDJUMvLaELvbzI
I3NkKL+0TkfgreyY3HpteeSkG8U2bF/2ZbLQVqZtDtUi0sdsS+udV0x+3GK+2k0QAH7cuLj8keqT
d2IW56Yy53ulJfYzXFg8UANwcUTNWCRKWdKeHPRJompYv/w0HpCkFF83GC9Ym1NdPIB4QfD2Mcqs
fb08VK4LO8GFORwwBxP0lCa0KsoqtoV88N/oGUti2BCwHb2QWLHX0MY6MrYs0lhsIJsM6JIMNdw3
DuSFsj3j8N+VjJjTfWcmgVmbb+2tkk6bfjxgb+YnA/ZLbOIyUxsoTo4/2vsvsfqguEISgOJ7ICSO
nW0mXhH7IaBA1XOwI8kwMhJWBREE1nD1rRk/4ltiIMvmnnOriL8AXcTDGWcL9+JP3bU+LaoV0Qvr
XlUnhAZkUW4q6q/FRq0Ir16gM0a5LOz9sLkntDTolSBXnqc+zz2m5mEfnK1vcDmpyw9sCAe9wO2P
VNxnWQFmn6UukNiJQxBd1tGUDHp6WpFn+7YIy8veFokU1h8MIysiu1sxIvOX/uXyJVukm+R09BnV
ArQfmXDLkRuUjzwDPOrwZ8mddop+U9fPzbUjSUk448lEASp2cLPUy/p5nZlT+rcSvYlJPWCjgCov
VRXGAHZk+LhAS1X4LguEYh1mnoAhVYjIQ8wNGvugKKDn52absBZp8V1lqSZoms18KwsUdL7aJaDr
vQ4uW/Nzjjy+bQ4RxcUhd1eaV9zId2XE9ETx/Viw36z+7KLFBfrf2svzXL8IjaxSv23DQPTsn4cR
T9NHmcPeqlPHO+k19T/VxTC0ITXSw+Clp5ItJ/w8A5/VFFQDZGJoc9tc4xuu6ScwWWHwZn51q9uL
lrJZ5Hi7aSNId1XlMIZeI4JQG9A0EcHzYmkSaIpjhxdDoX+uOkoJWme0ny3jCLmxJHgH+Ll7qseC
LLma54bh230d00rERILLUccJU44a7fXU5gESlKT99MCIcUtlERDO1mn4RAG2K2r5XzXVPG09W58L
vrJb/bE+WKKQe5484K23X+lT7aKYMnbQQVaa51yvOfKSyiGvSKhhS3L0uFVOoW4nFaObISt3fZVP
Jm71W8r1YAtkGHnJmNI3WfFNPPJWwoUn1rDhwfUxBtQDghsg6W+HhMf6gI4olg025kT6EbrcRcou
MRFkzfI9sh/1Dq66tQaojK98SvORLmal/5Q8IFFSqUi5VX0nP3mXiixcgUmBLW0c6SSLYhQfyCxB
tWbZi/b81IiovejIUJvxJH7MxrZfGEzWPDDFLwm0wF68325CitR71IaDv8frZHgZLrihjw9sSNvB
7wu6dZmuz6RZNCdmRe5aBMmmixUCMOZgQGT5YrCO5Ax476VHLW8lCFxjUiSIuogPMw8Frj8oXvG8
XIxVkyBN7BpqDujkoV2bm2/N8CHbaeU4wTjEZGXwLWi+RiAuGqXbhcbeV/tDNtn/iIFls5DLpkI8
DH4RSUXlZ5p4mKzBfwY6TVP5/pn8quBZ0blMTeCXUAONCykRAI4NIx0PWMWNALLeWn2aL0/Nzovm
fbWrtHvrv1JIjTVPKbCD28kQhu+DNM920vGhyg7U28C5Lv2NEs2CQVMELMSOrU/RPE/49+FyaMmy
wP2PeST+ZNN21EMQ1nkVwvwYXSxQqbF3BhdSzP7t4rACew6gQeHP8k3yKeBv3j+wHtFyvclw5/FJ
g1GQg4gaZ6BtTI2qSSta/y0lA+0sc1vJeid/JLry0Unn2VkTcT85TlYEMQyph5S6DPuS3+lXGUBb
fBIr9GCVYXBhFC+xXC335raxSD+npUjH1JQ6JUzEosDvTg+gqawXWOuKBSKIPbZ0q4V31ALFpsu4
r85Wz/NfMiAxsVTYe1/g4UtRwFwTH9l90SPMlOE60Jzkw9la5EJDioGKsvSVE+bvdfjbtSmVGXsD
qUk0QgEt26kekk9ZTpX4zgFrolQfs8fnaGmSNLErGAWrnCPY7IcUa+zWyJ1mGRcXap/c9r6j9AGC
upE7+FuB7xJZxS8UC/UISdpyAuLZErSv7d521ezo5QSMyRARGGfivBI9gIK8/N5SVeC4cnY8Qh73
syX13xvuvIPrCDAJjNNA8VkW41xW0ALx0B76yBDlQkTO+hlMsd6HPnaIH6ntwFEemM8uqrk9Jn6O
eyesbxiwbRdqPb3GeSmVBEHIpcLYpyPM/Td1N/t2vZ174r7F9EoJpW6eiTfTk7XtsAGtUU6HJiwp
cbIdezJbz46On9VBAtekOR1D5VsmC6VnYxpLyhm4K62KTG/nvTtGF5SFxUj3JgEh3v7luhhTmnvZ
LALNbBlizKGcwdeV5egbu4yiSRwPVuzafnKOnkKahee+Pf6UM1ucvMQsH2Kf7I0KX+f1lLsLUNBD
5Xw6y2zGAt/nAuFoL5bv1WhQ5XGZtfo2fChYdUL9Wg1gMlUAi2gA5meKtQVniJBwt9mBMEhf0VLd
NRwfNYhDXV/K26Zt+SVrWzSDWG+W8gk2Mb85cjC7wh9ZhSFKn9TFhBZn8xYzBp3vaKobNkVKw9m+
R1AAS4j7ng3+caS1fj13NrZPHjl1n5u9dnZ6/af/sTxr9u7PSAg0US/C2n1Sl0rqpGEt39VYExO0
qzf3wKkOCzJxfkR1IQGBFsVBmdfyyW+oxRkRp5sgA32tbZh5+tV16BQUg/fqXeY5LS5LiQQpmOuO
aXC6dZgriRWeQOTK1Qpdc7GddGc4ixyUHdfeQHISCvbKFxO2umHYBH+ZJQ+1m5V41bx6qBEru9bb
XrP9N150leYNaYD92GtqXZCfa8wR3dSSkmbndT8ZQS8xN2bKFoPNLv8gkXFQR5JwRgjjvVQL4ajJ
R5jzWG9V7LUX8WB+8nk44ZYKKrpxRT6dStY4afvQLB7MUYwVARNz292adIX2ezpXnB4yQxkVF5Xb
yIp2atm9SojdmLDyqTt/+giB+T9PXwMwBmxLZd71j1d3LZM2+udml9MB9miWAbVVI9hcR1rXxanh
uner0CMhDIs0/CYFwkLSdF/svh60MJd21sBr94bXsK0s571TBQZJPnoNn6vgxsXue9yJNTW9fcjh
LMJBWlbvuOGn/U2Kd93NZjlaALHZb5zCxOlpJP8H1xNLASXVTi2x+y2QWxgUR5WwzsX9Txr3d3gT
bDVfjpPFdp/+cpU79dFDEU9kRpPmEQbZFmAhEFIHGMRKc8ioGZ7Ssr7URMQUPZdfU1whfYWJ81rg
32pe/8xbKRXRQFfiOTwJVPjwFXAJNrPe4ttagMgRd5ejSq5igpwgweS1GzMBUxuUZCggHESWRrRZ
+wQzpWrPejHTH1KgGfQIY6MFyhNCyNP8caxe0eDqNwshSKVmVph2xmZXH7KieetetlCuoAoWQ77i
KXodS9PreD4eexHEI2tsNVt8wzXrfuRr9syJB6wHhdZIle9YlO+4eJDpgqrW2zAVOf75RZGtL0ds
jn2W2zpib/R8g4P2nsomCUOZiK29ROAeYKGAEmTTjdWGv68qVThtElFxS21LQ/D8jcxiX5KGEGIW
U8mX5oZ6yGMQ/7Dpazuuh3jMVr5q02bwEjM1JtBscCCD9jQ/DqRBOhiKZ8o99mxtXmUWaVGkPRPm
m4o+lYzCEgbsIj4hpCJAtAsErfEvOvaLd9dcmg7gTgnVuTiWzB0u1xjwP4oPHYJ6Pe8hPPI0RB1F
hgPr41h08ooONtaryu3CVYH2to/6p8WmU3qkM+tUyxsN14Ojlub8+pDXoPTu4dUDIMOXXIAkpLu2
Z/Uusa3cuyreChL1Zb/smbqQjfO8HeaGlh+6dCVn7OJKSgkCv2yt/9eKkWCnfB+VDX16JGFRltWE
Z7FpMtY+5r4l0M6HpcQZ+Zo990++1AUJ7tWkmSmwTndE99Bhwh5KU9vKlc4Yq3B8Ok8gHu91uG1u
S2HMquwfSl9XsiEt/xZT6GKD5RYv3SbhyN9HpffXeK0+2AT9d7c0+zR68ozoWCTXlX/wlp9uUtUF
p+WSbWN/ck0fjpr9sdynLOnzhfUL8ItY/XK3awCxFm31juYDD5T1sKxpBH6WgoLRvxcsi9gHfH1Z
933clKr+MbK++I1sT7du+StbO6BYot+Fr3UYEmGDjyRUHsrWGsSWPymiIZKs6tZX3mkI8Qb0SpqS
nM9+LKHIA9PsVx3vtI0gHtDwQLbVpfc9LLTzC0wYqvp8vAc91cf/RroJjzpsM7gPEKcWBIc4I+Ot
x+i3K5Qp0Yaf5EHrH/VumX9m0pyFAnd4gtvOg9DywL4CI1GZzQm5fd+1/Hy2UINN4bKV1yEe/j3s
fRJxTIXz5jfJASm803sVARWfGw4Q1N87pWoat3hGVDuiGJGb3j6/bhc/Vym+XruDnGatWsYLTak8
DX5RKy77SibDarBDX3F9yfM89fpf6AiCsRVI5avMhaQWrPpeDYd086yeu10ztbzVq5BuMbE7m4Ij
EtJrN8hu/LIIz0uLJcJDbFebbf6NC5JkfjtWMqMJMLe54HcNajLXZdbHZZrO0vpNYmJH982/iOrQ
m60bTbZDtKnf1ewMDhWNNjW8EqhcPp4MuYoOSxy/r3hHSSzGlf3eoA+yBXbDPx1kNvEB6EDkeAcQ
3vS6Hjo4VIuGoUc4NFx+Umzw0BY6Shzc3iTnRhXQwkmqdR7lVbl4fOBX1hDafJcW4YAEyd1evPp7
smnPMvWqXYTAtvoAktZO0XYCoBO4Ak/f9Ku5u2w02FP54+Dpe+4ew6M0FlFc4KrBtxzd33Tsa2nM
ZLG6ue3Yqq/BC/eEo87ROik4aNTPvahVX7UCBKaTGGhWma/TQes3JwpeUUBbA6TA74CVFvxNzeeN
qX1S/x9v6DIWNWh3G89I1qOhanotgxHM/fxVxp3TfJQ1ilN2NLtxVgj9w+qe9dS71UWxT9GyC66j
9oKemms/9t8uzc7zxyf87vv3NEPLG4bzLbCuWwZ8jnIViEaphi9PEufsBvhEYTbMetl0esNxd+eN
CkIQPGygNvE8wQkgJfuAYkQHdz4ZjvGr0jfnNeGIiQH+ChqnrQz/d8a0Gx6mQh1a8kQyTXk28IkS
YoYK3dmxKLQ6vKmBNu0462A3DoNjdQkk/A4cifknKB/nGEWNXY3+zNXkFYh1qduI64aUHMaAVcIm
/VIoxY/Y6vmedXAyJ8EqNfqrbjKyaVmYVI55tKwZNEn160LBKV81erQdXrYJWzhHV/86gM8hXjst
uyYJymHOz6VzZ6U+jlzmsc0UHg4MYGxqPC7dS2FgccPaMjeDAk6LAwMcd6fCDJXDGUdGcg0Fkk/E
G+TnyCRvupnM7TAPpz41JY3qN5lLzluW3rH/G7PVM/bSCPxVg5nZz2zK88p9M3VzOQjE7JaDQvJa
vQQ3rct6QcEKjFW8dwkKX9h8d50prUV4x7HragzjbC74U2qEqEU6F7Onp1j7Sj73yOKsAbL6xnQt
WNbvLwzcTEcor8DgFBQ1/H0z5me6l2kM4X5lt2F4USVjQGaJLLgpxFbh2kHtP9PEbLq9VzDChqNW
+9VZmJsRVi7Mz9CfwwXQf+cqHQs1hCk4+OGpRQtdtFkAyfNifXhcWwcDjHlTOmjkBIP0jFdi9uvT
LsRNc2OM60KkWNhhC22S8cAU3Fmut/2xtT9p1haJ3lvlZvNVDW2AQ557sf4gqRPHV/nl7oa+KzFb
dSy6LWR2VYkm80FwtqUcalDB38Q1Hy+kLlyfZHSSzJflXZyUjf1EEStECFOT2z63Pi/cenXAD4Y9
ZGcW3ghjUyqcz/Lx2E9XkmB5AoittcVHMmTax05k+qPIY1buRlSbBynwY9BJdTblczz7++jOauz2
8BDoGkDD1fqi5l31Riyzel8yN5BpBP6eZd1RpuMprnVoT6Hsosk3PkO4/rVOv09cz1K2ugYLrFP0
Zuz4eoqSnkPGQRT/HX5Oa5VxJ3aGW2Ia/MBJMNGRliNa8yCd9B1MNegyQ4vamXvceRzN65aOG9r0
tdRC00LuJdjMZ3ekiNWvWQeZz/oBf2TLuXgEJHJQyjJe32//C77DKCIgK4pC8LrZouUOgYiHynKL
+nkV5l/NuAPu5UufhXNswHmuDkda8MvBF7Az2VYHN1DQBNnw+LYR8WCTlAF1qPlHuIYAiMPGerSm
jFl99k0FGY0uzUae5FDYflBkM1VRsD6tboYrrLwZjzcrdICimSSFQeexauMz0wFdJUqGv9xGllyQ
I/4pMFZMBFbq02zMLGzl848QSwK8VpwWHpigD1ppqfHGCsG53r8o55Tb32+jrS5vIJowxW5EXG50
HqJQ8emsAiGXSKK+cTogu2TAsNAGOhnPoAifKdNnLd/cEwCrjLvTDLMhq6FN5HC1y/oMAc93X8uY
f7saybawW/U8UZQGOqVorLYFGme9wN4y36em4ZPTGYEOrp/P59dXzrvH8u178zHThowRxykbQnxo
oYPN2KSdvBrWp03Wfa84gGQbZ9hRkqu8+9qNeDQRSQN66gkxSdU9u9Q5nX6dlqp78IEJ3azTUK6y
RYDJ8Gbpl90m1UnKMCfJQ3dZ8q13InvjmMSFzzkiLGEe7s1Xqa+XC0dBMNUTSXCLuxmYSuJsJr71
DL2aKoySuqcQa8jocdTY5B8tM3i5X2RPDTqGBCWl4XJpRIMwU1Ad/hLEfNPXIVBbWA+b0vKEkVYs
YVtWmUK79FWqj9l6EFKRK97rJYHkvNyOq/uc+T8Vo8QoLp4S4x+X6jrWH8gOn31yVHPhPErkBcuT
BsF6Ku1ml4KQj+GLV2PXd/WuNr4wzxE52ikIcFdyQs5RI+0aXWrNiDufn51Ry2fJPfPlxSg1iW9W
ZGZp0Ybrv0YeXCoA1BSaOuFt3cUzFeVeHhFnMWY1jnpeKSOswAnLF34paryks1xNVSdhoH+BdDwb
TxcfH/25KVLBmdnEJHiPla2m/ToegUSkUS1x5syw2Yjz5X499vDiI8oX42VK2/lq6fOfy1KU1vU/
Md1BL7PoQ4i2RHtHdbEaU6FdVe/JYfrQYkN3ZY0i6RQAVQqGiBvJoHWNUKx3Kxuw+ztUjaNiD75s
2qCjen4qZgj3xQQfo+5xqsluP8ts8rqGkaxkQ+Vnt+sjQqHbg0dP9v49AhjKCMC6d38j2GtQN3si
m2qh81bVh8gHbH+6FTyp1xUfkapMsI7LXjOPIamXMEqJYyliBLDFcHuyJHbS5z7mrpHN0CJkTPlN
SGfAWx/0nmHkXjbvr3DxtsJSiv8UmKtSM6aAymtJIwv9pVQF9oCTFqcduGdMyRCLeChBj1Z0KWJm
sFIVMK7K7/IZS2QR8HuFDH2ZE4LO+GXFXiaKdEeaqu/SIgUFoQyG6wsuA/RUYIwKaNRMF8SdBGW6
ggWLLGVU4BeoUpoErS00KHRdDlOAQrUvHkr49rT0EWXq1MngVJoTwsfqNgL2oBwu2vq+ccFr+Q9g
FM42aDAfux0TteHMhUBCQCObZjs6C4nXOPZeZtX82bZ4wwXtvmtY/dHGhPsu3heVYI2IomXXOJPe
Wp5VbIxs676slo/ZtUH/DOF7LG2VY7+/zTKqjM2YCzo4/Oxis7yyk2rTvUEmeFeZdnz6UaMvfaJF
43vjhXETI4GfZcTlAf0G/IBUWf5rK3qSK+WGv23vjlStuSt1xm9Sh30eEKmtVJLD9861zt19HTDU
YFJIgJJXQNXwusQM6xyL+k6EBJgonoj1IcdFSCTZ2q8YA/KJFijJxsJrlnsCrp7ewS2KlZBY10y4
MpX8Iw8+Cy4FDfoslEitgjKgAtjQcLkvWjjfqbBanRTTII2pRgwshpsk9YV2O46aqbq7NhpZv+78
+o+0ij6yzLpg+zMmrJXNjHEzivVyVqUD9Mhc3CVlCaPqvjrVex36Pqr70xVQs6Gf3A6act9sJvKZ
aHUXBgVls5LJaWmD9gmiOJ3aaZNhTVNlkzbJ463J+HEa5IzbUaWzzOighER8TcLwQnraXbLqo3Zl
uSC+zB3lEWJdgMWxsWg3bV2bCHnoah36MhwzU3f5YFXnur3zFz+20MvW5+f3eT6Cem18uMZnpHNS
islun2MmLtOSHn39et6Skk6bTk3P7ufM/0ecr2OTP1icZBO+azHzedChtpd4ntDrjyVpkQqTWeus
7wp51KdWu7SMCRtFIz7bqF1xXvi+G3hUSgM99/7IVtMi5uL7bSAI3J7qsn1cnAoRQSZ4bFRf3ggX
as8HaZ++Seucp4jAfCl0Xe9v9+BDXkbM6GxmCMhKVSg5BDNtnVYwqjaFAZ2fxxRAVUHLc4JMWhRh
RCblupx/YgzDCvE9Zo4m0WhvO3J512R9bLtqEIpxjY+L6lQggfethE0QBZIUfbsjPUETbGJk+DUa
JSWmWaVAm4VRQ74Ws6h/qTBs0YWqVcaEKpkCfl75WOzEkiapFy+dQQ/dJCN9CYwp5EydkJgJZ2qI
9q23DreKE0FpbEYuhuT8wxiQQ5TY2KIKljefF3YWckZbmU3NO/hClK+2BG2iTJCr3UsHtt66cLrj
WIaKt8mezHUOVI68AEq8lF9dannNJccb3ZFJfMa2OHW4eXHN3a9ESAe4gUfR7/2DE4JOXaNw0YXz
oUXjeAmaHRoLKY6DMwtp/ouv7fZGdQi33npwt1xedbY6ElQOSn1ij/TkfiV9OwHdiqkgHhmNWFtb
xdrSiUwa+HfqIW12fo1UMmvJWzsnD2C5AyGFQB2R57Cn48kJ7sdxAgEE9Rogn2IUtSsWhPCmPg7N
VxneTi4gXB+n2icdERuUEnhP7T1itTDgIb8OMzQdLTmND/+WYWTEvahtDBiysQhXtYL6Pbjm8OFS
c/Zjve1CilXShQbejYobC8UGaPeZhI3TW8fJs6FiXqR5auanfkkDMISrX/NEDRD/0hCMFDbEbpzn
yZGrBKTdH508vMvZ2fTa46GTuOIFroMasq2l+vDZvNqxOPjfY9EMks6c23BCmsU8C6YZhhvej7C9
aO1yqjmizFyIochZ+XJWxsI+zGUbdVepQVpqWNCZWOD1s1Y8A3mhIY9EVQ2RGjdsvv3NJVU4QbB/
6zB9rBkMPoe0GGBtPQ8vQ0jEux9xFRoCJMrB+SsVHpp3Ch29ez/gHM6vVnO0F1oyAq4ZH7u6aXkT
jGV0otZeC+wixwtlz1n0tfR+RfAFSVe7aAg643Vt+EeE85W2eyG4aFxVLli228G5VU3q6RuTGNGo
0RvbiEP3VjvHIWZ/vju2Ba5qj2GJtVblOkuvjDYx+yXPixzZ3Ri1xVAihsleUBGdBRvlbsPGrJTI
89omBfWKyiW0ZXdIRMKw5vqVIGNI3uFgfWbrAocohS4UW1MN8U0r6mnrcn5gV7B0CZtt4+AUhTi3
R544TThhiAFDTEhf41QKZU70hGkXT7Tbx4vQA3yt/8VJ2a+25tUl39tttPpE7MKn10wT159C6PpJ
VGcmkja8rNWhkGjqyHYOrkcpNusO3xOtm/8NMOlvITeV4efhtO1kJPNTlZ/i8QjQLNZ4ardUELaD
6CMjKouTXdygyF/eKPrwoo4ELTTmrQqvmrbwQIqxNs9Jm5+wF502G5aq038mX1sHbmm80aEemuqo
2VMbIN1FxLSNvp0yLXQM308wMihR6aEGQVWAN1sDqTwCiLzm5ohyPn1HJpW77cXKHj5mBo+Qw23w
HK9dM9+XiWjTXB6nMITq05PWUwOHB/cNeTANvD7n/1Jhu0IoIo040lZ1iCw2AKdyHu/RwsakXJtY
6j3wiwcqBbJ/QCeQSYp1u/cpW52XpqVhkKkMY9G+LHrvggm9LuuTsFxnvcA8MFbb5I+pdPK3aYJ9
K/8tbKSswnH6K3/ZFOIa9QpN8LWlctFNP0systo9qNE0yb+hhi09oZT1azXt+kczslEHbQAx1SLT
hP7/nuM7q9MHkyEPHp5fkh8j2/syc14BXGNt2tUE0/5ZrvRyoZoW9AMCjdsdB5SGGSiwqKfRFyra
Akhe784QkGJyoZhrMa4icfdeQEQVRcTl3a/7YzSUydWCig4uXeot/5b/CHqazt9flMLgLshnZcp4
z2ghK/5T+dqBy5hZWRAeb17AvpCJjmtGnAPRv0cBjQ7ZnaQxC9nX3UmkSRLu+UZxpKPAKLL4N/Om
YIlS9mwsiiLReco1BAJtOgyVJfkbxW9/MNNwqZSKpbNIY1Vl1oRsvoPCp1OB6Ke5/7DPnpwe+1hG
xy09UQJPmE1vXIUEYJ3DdOV330JPYmnSYYzbxWnn1Avk6duu9IT57sb/IK4H8RLWaVuNtWHAnXMm
ClQSJvB9EWwbdZAKY4nS5hjbRAxGo52iY0VfNmkUku7qC6bBDlfvj/4Q+r2z6aFoOa0HaWJdmA0d
CY9boSqCTXh8pWMC1gEjvQIErbfUrAcUVgdQBvnPg1O7nE4VripLFCZvVaRY2/m2jjkXZzer/k8n
JUm2GWa7mU9EBn3ETwzrW7dmiYgcJtZr4AjOIww2YspzsIv3/oRTd+xghhFtDmEzL73hCRgO77Y8
voWR5cxzxpaAx0TqbAbzUboJNlCF7cL05C7GiL/Dro6lfJ7k5szdwGrU6yvCG7fwHmQoxlFyQIhn
huYQjrCS/OGaFkmpFvjbTShA5y2EnPDWqy0VyjCRbkPhtAA8EvdwNsD9TAuxtZeLo0lzQEWdl/zc
EUZ8yUDeYs/KgOTjenhB6lQbT0j1WWsYSRM+Q8gUAhPqsUvjWtkdGBghs9uG0O1LJqryj61QdGjE
/QsTwvFbqFhXwW7ybmxMfrNZCJ4uPbBRZH1Iq5QHEVRoPXlMvRnSo7H1VpyDrePZFAygrkBMOx2U
yAfq2DBS0lyxhqltBZC8RRZfXxVTQbRt0ZBi+Rtz1u4ZZJkka6wfTRydtVguCmIKf0h4NpR35kjU
FfxAguM97zgbuP6/oLwJ9PsgdAROEMOtKBxdL7lPQ03jjP27XMqWq5P45fKrhX+F7oz4QqCG8o6s
2JjXwiq04rjvjefxl3Jd9hBo8CD/T4XEYwYGGo+nm/izbCjrkh/xcdzYtAGqetT6QdsxrOZ4u18l
hv2w5TdmQwbZ5urbeCPoNAN9yDZnVyu47F0xu2ULTfE86FP0vQWqCIbM3gxgEfB4ZmjXMt5mVij8
Y08cvYui2Oh2+jKMTFN3Uqfi4mxuwltIw0AOyKmZDEQrXDer2ls6kHiN2uiA5uINSCf/L4OzIIX3
Ci8tgye2qaMthLuiV9G5+fzUwJOoYDC64wKezJw4KHHUaJ/qM/TWVKM3ivD0DVOIkyFLKp+H+Hcl
aWNCy1TorutoJJFsYZx22Ww2N4tXuiS3xkDeh00vyvlM9IL8M5JLvrr/B964RQiy+zwEDSxOJHBT
rui8Ys4oo3N/+dSXi9ZjgwOP1ouf9E7fzS1K9MjPt751wB07rVrfgJ3PScnnx16mbJ1KyhoAId8F
RXWQ/BT9nbm43Tm1/m6e0HLu/bMXuYXzDYZP28AJ2zcnFK4FrGWDqt+6BbyB4GXiABZ1JXVMms7M
E1xwfWGATCcwJe9kAu9zxa1NklQVsHs6tfJ/vT/0w/7sEHkrBr9Z7h+LfLq++xqoTxwgvsLFIygy
qZzraQOoXq4d0Ne3EgtUg72iUF0Rvy/OhdXE/lhriodTRBqyDtc7PBLtUkPhQqiCVc+U/mKL+h4f
4l0E9bqnVVI9tsWYJebHDLEO1r9AUpg6BhahTbDPpO9PGQB1WKQ6sh/F+eEwcUGBJuV7rF4zeIqD
wmK2rTSXfGwbXYsBenKS7wQOJMgD4h7ckL74b0GMIlhDYiJJVWbG3OAKE2uVXXhWQhV1V5P2H6go
kNMfi8FAVAvSwEK/6tEe94jGttxiizpbBX3wtQ1suciKkL2jXiu70EDs4v5KKJnk/iwraTbRVgzW
l1biCpd3cFK6K22MP7x1+idUH1YKmnRoqQVeoXn1ECFteh/MOFgb6s1cwo2cRIcgFm1L4Lr48Jqt
tU4BRYh5Irhwu1yIn8F1DRZZaHH60vDGGJqFWU4HyBrjOmBFeGzCIjunqpTCN/RRrKsn0cpGIwXm
PQw9TvD5CXhdSJ1XkO0KTUAsgx+VEsA2bAfObxPGTLAvBpmm1Hl5/EsHFi8OGlLzv66A+jXa00JZ
r3Wt0rh7zaggSAxmLE2fZElXVASgxvSWmgCRBZ2qC7ATZxO+Hdfshb1Cc3EV/DyJdasbVGLRTXDk
DmDnvvprkCzReYuRHhNcFvNpvuXrOQ5Hey5dBbYNCpY5CApM6RnFnds37tftcryP2DLbNHFcPnUa
jUWpIra7yzyJfhQ9v8xV4Vgz3BbW/OA2GUWar0yG6VNVBJY/jPNVdk5ha1mpQHtjCWyY/OqkycG7
+DWDaZQO9v3tOrdzbZiou0VMFwR/dgf9ic1mWABKR2EttKnYk3/NRLAmAWzM1TO/7He6ieZG76O6
cB8mjHbeqgOkMlICGJtFVOHXv2iUE156wL/AEnVxgkwZKRo6lfV+VtsT49CL+gYK2LhIgUGQxOXH
FosLIzKLRayFr28MSm8c3hEprqxXZ4DDGpKymM/5cg+MhdXXbTuM4iitWmjsAoulbnfFnDtG+OMt
Dws1BfSrEaGnmA44d0qbeSx3RZaWK3o+A+Levu1UN5bdYqS2g2trFpDKVZHWMb+gP9uDP81ck0F3
oZtYSaS7DlKdjrzuArrQ8qx2A3Gucpsq1fa6UdNtPjFzgkrhRB0Q4i0n2BiDIvhdFuPFO+dEv/qw
Nn9jBzrqwT6fobNEpzO+EVCnPAf4p26EfvGtgMYjgXhcB/eRuqzyCivtdGlO3hMJBOqYxBlS8O3v
tTHAVHIpyVZtTG+gf0NWPN45F1lQmo9xg6UQZnLMa8ENV9ypoTYrQ/0ep488DIN60UbR91E8Jyfy
NnSQxprvPbo9rny8jHwf6o6jE9svrQmDKOGiTm3JO1VYLt0J7CUiDbSrSlRy3AOA0QyFSzVTno+7
nanC2KzuKPfM2U7sbjqdc49ER1MsrmATIa18JCuMjamNIeoUCBxzdS+er0iD82ZoeftF6Wq7xONZ
gt8cPvLTxj0Sss2CJxWBQztZA4/KzYAxEZUgktfftFYJvhZNdW+209/hkR7jTm15nsVv4JlMmui7
y5hEa8VTFn/fDc+BbU6qBWJ3zr11VB0fvoLLwz8HufK2bmS/Wb9/TG+DUsjHVdqXcYYCz+IotQr1
RweIJ/jYi/wu7lPSdy/ViKBW6KLm05BsgqsSY9PqlFeXAhMPS2MvgRFU9yQFzu+rVpQJclliyGZb
8HjcEpbeVeh7hNpiC13zMOMq8HD9RNFutPJIzJGncokSX8IKUwuaC6kbQqNF/15ru5MVMRu6t6xX
SDuvYXBIrLRhNjCCIEhCKd0v4N1YkO2T2h2KqGxpjdSnFdsahjqaXru6o3/ktBTaF35wACaj+7Gx
qfDvWWJ2ESCVuNf3cPF+uXB7x8unzWYXkCeSqlsJhRuZrZFSBqVh1gVl3uoAQ/0VlMbt7QMdhUvk
pPueTVhBK/GEA0oXGJ/cMor/5eUzazu+xUdoxYhb5ZFxYXa89V6Z2jyGgWDpG2wekn07fT+Gj4A9
lzRSeknfjtvhXIfAEg/+0oMBOufp/j2tCnSFkQLxXuRhv2nG6AuQwsHYg/B850b192vcRHQJFp0D
LBo0llC173MnqhlskZjfWS8y6ih7eJL9L+WUx+2ZMclWTUwEu3wWSWjnSFT6EHVbVA4gM6U7ZzDK
QMuQ3/wZPinwvGVuVBwJl99leoX5nlVRMJVHoZ6LmBbhXa39j/STL6i8u7LGaa0Xw5oKpKalBTWJ
sx0ZSjD1cTKD8HOu8qxDmCN+yRDxD++qrzWyFkKz/422Ua8fMFEfPv5IiO1CTQFVScLUsUVVeSRe
1+G4KrnTCoqCysJ5tr30LFSUhXXjDv6ZXjLAkcCpMwyFKDismTuI2nKOoZ1Xpv5nfO8w1vcZ0lje
uNA2MyOCVzRBt9Wi9W4mQ9BeWH6pK00mvOtXVbgBiVkZr+DWQmMTbD6rseuv4EH+hPV9co72r2nv
S/mfhvZvUsNlTNg37awvA4VVDIDNwwyM2BWKAcixsYxswGZB5+RycHDd44V9qR+SofroXCQUhkiE
SOVPv/1FC20+f+eZs7qc++HxXEWK3B4xeaZWYVlrjNZ0nKlyOjx9NW9vL/6pv/FI0+RBu5E/xBDA
wRot1qbObiZd5TBXKJH+DZyf2uGEiEXEDZbTm78r5e0XaniuRrAVsDwmoH7YBBXBUg6zwPsZNoCe
zHcMOdJGf6Or6mhXzpWbf5E808h569FQlRjOcEGh8a5sLxLzVJ9I7AmxXOoEKi7z34ZJYv7a3bhZ
RV1GWTnKvjxOxxXWRDu4lM68VFNgFW3TFWJBJou1Xs3cBtzZ+cCviISJtwiNotHAR8k05xPb01RG
mU4bE5FeyDLkb8TfHPMx0Lkx0yHi/AoTGLmTJ6LqbZ856gkn5yaEnJQqPALIGRi0eA7/I8KvBDej
TblkjtOK8YRjTXc6ByuF6z4mbHMWERmC/5z28nDpWZL80baFl716LgKIbQisTHCPbOCqDMXxUVrx
2usSbMCo/thKlKFll7kHx5xFNdYbtTtqYtSVcygIf5Lpbhkhh+/azvBT07DLG8OmazlDHaQiBrUT
QdhrtAaFAPh/CYVp1Ayfy4AiYYTUBWYLKxevXIGqYbobJ6bAPXVDf42sCVHJMEa881CLQ08jPg3e
6kPDzqigWi16/5c9O+ko7hJHxEJ820mE09HDUUHNr6b62k1AZEpsBuhmMTZ6SDoUkICNWK4fflRI
BLqTnYtIDDgsebR+E4fbniCS9PgW+efGu4M7rnk5OMhFVSl5SwBYzv2sc9kz4jRnKynkx84PBG+u
c3I6S9R5T928PlmqPGtsp/NQc/jLU8jW36fCG7pzmnVOGgleVCRVmtPQAgXJUYHVaIbnHsqWqeQC
J5ZdCafEmaSAmZDDl0dKru9KO0aC5lKmFU9h4HXM5Y7Uer9v8fSQbTF5UEPeqph/SwCBJoq+ozev
Qwibims9a294o7xuAHIXwl1XS0cIdcW2WPUhEMRjr/LfNdoeLrd+s5Y8tPPHr5hmmaqS+Ig4bq3C
Tba8A8RvGRrfPVqeB1NKgbDtdnI5iaHNXAVZb7v6jUAXlNNAr84bB0mNv+T7QMA5PgfBkHyFWbXu
WpzLFKo2qW/VFjU8IQhF5n9f4csqBuBWzTvltgVRY81PAEbV0rFwxWMqFIPVu+68bNxAcu8Vdwl7
UEhbuBNWBymu/yDoHAM7gnSCFYqVdfYqcwEIUuEFgsMsabJawnkcB7OTGk4xXmuY2UWWgex771JP
0R0ytapeT4N65psx6jSjMxsAX3Quy3qYgcjCueD2I29GqxMsapiPr7G/+mTCFfUap9StmOJLM+R8
fdMZ6wIpSF+vp/iDL9TsTLWJ2snA8rwJxz84pYqXV+bcfPkRt9KgwmVRAuvd2i2AwqCxbUgj8WK4
9skoMIZsCdgjAmKLBDTIYrJRKGkdvya1mDb2VkbNoaX4ME6yN28EEvl5rMhby28Hr5VGzXilDVrC
4IRiuQSxjx8+rqZh1B44horxLLXyIFuDxBQujV7as3QvrggqObsDGLHtAMrLrs1A17bAXNtbRxVl
Wb2/Bv/W6VtMnh25W8rE1X38zC2fXTTacQA10RkFGU9NR43T3HoQ8snl2I7j/uLGgjNX8zvKR3S8
imLDsN+3FFM+5O0KiXvxFHV9TGTiyX+6KnxzRDxXZK6NMt/m+bArENMzJqC5fPp5w1p7/2Q4WSaY
+YcWEOSJQMhhtrjh8xeg8wXfp7CFy7NHQjgjicVxgecSQ+GheKq5m3zF+x96yePGdrS/UMetUugQ
KkHIO5H9hevjA0IKu0nsxDkrNWzxd2yE7avs8KzXwYSU4WtlLMTokDU2CWEuFHIsGIjEWT3xbsj/
Zw+oGSdsRmQVTlYPHRQwz3Wk6VSP4PgCp1KjmHsWqG815WvezUjcFKkthcGSOPSQa+gfpTdOBXY9
NssvV0WDs/r+YrroKZoipya1o1p8RwuCbcsHVhM6iTtImrjFH40Z0JtzQTxOnaQPvxtwV/nKNXdv
z9BVLgE5l+Jr3HyT5qSh+9GeF5M+LdfPoTNICBbCoh7b9+d3NpuxVXymURTSfcGootL6MeDPi5gg
Et8024ji5YFXuWd9FaEqFNKBZqfdg/OhKyOV9XDxznNXMNrsHdCif1k4z1qtkOgvEWf2t7jCbmmg
qtkoo0j4mGmLdVcS0jLrs62unIy6j4+i33e/KyIQhUKfWq+6TreWHGPSVLzDd+OJyOrDho6MbziN
qMAC4JYmdSuItWYx0eeggSBwGBbXWE2HedzEUMFSbCNiSHiKrw+WjOHHRTlVWMiHv4gSWvpzqd3m
TO0k3h+AVXHz4qUb9tYp/vNtFN7Muqwl9O/tpMojACDFrUwCKpUCZfIIxLqsySFqpXrdblDwSZlT
lKTisS0G6X2A6JjG8U/AJPaipgKP5f9OL7sgwegZZDhndq6tYk6LLekuR4/QPWrIR7egAqhjJy6B
Y9VCWs5Ta262gBzgf84YvDHXjj7nXHBEr77Fw6q6zC8S7gsvlQ+tyULqq5FKIXAophUQOG5qkQME
UcraGUHLr6TyWd7o3qS7EE3aA9JC5ZzezdZxBs3JTOC8fbcApEMwYZTiQSUzR9fFtR6Zb1g8Fasj
9BFp9+Zrr/3PVjpSwPjTlyi/jiQ6OEoNHmW4L01gk+ZX/6p7H37ToLA6P9sxQCpurZJSSQBVebw6
RTUAaLJal8qIqdElDe/BN0DTnn3/nTN6T22f9dR0Pm5W2Umsa6zYzJbgKS62KCM7Rj0Z/J/DnZTx
Uao2MoZGJJKJLL5mVA99xEBluWWiqnTBVcfIdy91a9zcXwFhCkBPcO9BTjudgiFwi95OSol2s/Bq
31pPXSV1mwargyUOyOups53Xc6TCdwfM9dhlUImfvnlVUjACo8rwFkiVGzKd/GKNel8Xw5hLmNdr
liQHreerq5m2/5D3XhR1/zbn4IA6JHjjwxA628XhKCu1q1zQydZERgwlm5pa0VeYywqNemdK7GN+
RJuPxrkGme0ZfE1xIrPvKIAYxmbipuhp1uBgRox6XrvzVmIB7lRnaUfJmxd5jxew1XscmgnuEb+/
iwwFR8wUX4tBpIDbejgnlfAlPOauXiib9hp8QH3IMtXeAhkELiS9WIjR4uXx/RdBsuYR6z1DW8vu
9TtVuWwUh6brOBhAuaYcYGKuYqiO6P5Cw60gijvTEcRgt+iGexDlUyBqUcUKqSYZTIolyOr7bsd/
CcP5M53C/kF7fCEyUp6P/UDvfnrkq54KDNSzOXqGXfv57TOlsoUAVxqHvLO0pmVrmbYCGCJcHvn0
wBGmuXQhPpJOI+h+1VYTsnxraE+U9Xu1FdUuFuQktMWTpGMZG7tMiYZewNDujbDwi6iZicTUd42z
B9TSR9ajwLLTPlGL2MWeS+UF0S0fyJnIP2kSQOf+YFa/twu83VnGBbd2PCijB5wQ2zwboddJWmRZ
kKIXrgOARydI4tfMuy4CRUKG/0DWkJKfVYVAvTVwabWOJoUiJb9UnEoLQiYP3qfu1/8iZnUJ0+oF
aqkZWKBQP1ZuRQi6fLse/I4halGqpPS3UtshJig2hvGB3XUTxqfTIRCYNKJ1NcFcDQDgg8ij3VLe
kfbKAXjF1LM3GOX6xdprVQ4YSE6XNvdHA2T+56GZJTHoIVtJMeo5WkPfzJkvkWjVmiV5+BfQuWNK
EsTQ0XF6xKpBd8vtL2CzYoJqlmW1GTq91lyFxz0oPhyGsjxJR8T+LgJqVrvacSworXL+WiLI5lEp
Ar5N0CeBc+Pvr3kHmajz3c0Vzpew3mwR2enHSiePe1jCCKD2ENphDXk1/5rvy1LJojc6KWGFu799
OqY/PtJbsUJ+pz4F+crjFPAQChuDn8Cr2Yjr3tFkfoWGebudIEsHsRTYlPxlY0g7o7JsigH6DOgE
7zvg4eC0KWXZZpkNuShYdgnnABUfbGCdP/1dmRaSWzBZEsYU46E7alQJfaAq94a2IXYJFGKtv2tV
WgPet19BCplGG5+KgjXLoP8AikJzeS5OEaOg3L1uH5NCL9ECKPizSDTCG+7TfIEOHT/My1ZOFyFY
3cR1k/ShRMN0s0nmG4NI0IGcLJV4+tlXcd1FllffVMlB4f5DabPMK4oIJ4Y08oIklsdrZYhaIGO4
m4h6izRcG0mTApyBBzxEWTvSvy8FDPDqGCU43hZMpU4K1DGJnQ9wFUZlQ8FW8HL6ZHsrnthKnjsK
gT93FSZRbjyO1hAyTNBLLRfmUHb4T92o0Ow8bTNJqLCMxmQaZW/IYR4Ulc6jXWAbSfjX1C/fey2X
9GtFpNj4JyVqEw/Dc6X2GRA+QGyAQpBheVV69pwmNfA527JaV8bHZnhT/iSI9edjWqF+m10pbZbT
TkPcka5k3wzmR0H+tayQ1jBFUMsGmTavtAXPiQQuaJBegO7Rw03TJObwKmMugHQFA7PserUsBQIJ
88Olm33Hpy5BPkR6VAtjkoVcM0nw6H1hkmkqPwy0xEZDHQd1cPqJZiLqP9hYAjMIg21fnWz30pfd
fWyvFAnM6Q1JgWkbQW/55DLK3EMq0I8+3MtCpTzjWztYHxUNfvt33G8/Crffs7WoZYsSGJ96+ymz
hDweIhlePWolO6BfLyC/q4YODWJQyq7AMHpPpgoWcVM0Z4QK+5EoyOxsMK1WHg8Lk5QBPqDS8bZ1
/5uR4u1HSbSC4X9vD6sBXvJ/RITnBgrL/yzMwnuGuYqUAr3ZTWT5xxegPlH8dQQDT5rsYskDXSPn
L09d6QfH4aPBH44wqPnQTof21J2j42x9tS3hJTzr3OFh/ZGDNvNedE9JzyyF6ckAIlf4KqoVOKxe
zUkMIGUXnPNg2XfZnL61FjNP7B/b3lsUtEQDk1W07Eq8bGSa0zxGII+QjbJUcGHPxFlX+DvYXxxh
w5UyDPXYN0R9oqtZf8w+kOFOk6LnYbpNG65UX/9qgdY8i5wYcBvGI55m5jXlE56qNM/yL886VR82
13FS+gqBjc0/bC9sx7VzkOFU4ktHb0qvnOx/jbjWGncXq7QMFy42cOwN7aRqwioeJaxfUQnOBdrq
LsAaba0bx1TYd+IcV3ldjZ65Np7DrwJQpL6w+toVEedIeCaAb8U8gJw+z9oDgu/qKs0OHIOstUWe
Z3aR8/47safcpTj9iPcqreO4z13Zg3djeuuc/hfQ6snLEFBKep4+VgqjXC/RfBCiO4MhEYqOZkh0
aBidzwS3wBkIMzE9GKerUXJ0LvmGkZDVGvigQ8MzQvbRFuEaBjCsZOhvzV7t+cJ2mhNlVRwEEqN1
1KFOkClldjSqFlaBW91XIDCmd5ddkpULfXX7009g9Ft4R4DIqv796OMW3GdRewFj0Ro0Wqbmvt9S
n2135r9+U86YkBYVR3SBEuKaM1FfLZ5vb4nIZoZuDHwuCiXbv4HGEg9CfpO/o9E1mxOLCpgAHoDI
qiqAooRURxzSkwdCZAtUYksQoHphIuxdiuqp3I7DvAgWvbr0bqML2yyW2DzAWXezxs6aGS0f31LY
UKGlcjXUMfKLj0GeLweTfux1XESQgedayYl45zjSVP10Vu2Q3wolM4JPT3ayyefVhPmYK4jNJdj9
QbfXpRKw8W8RO/f/+HyheIUvZX51r2TZLzTaZcS4Qu3wqkRRx2lhy9p1OsbVsJOEb4QL25ASX1Cn
UcXZokWUiPX/b+5XOHk3AsqaqyibL/NmgUG0cZMbCO/b74R1E3sMfepnQUGrFmVl19XgxSZOIxSv
ft4stlcu61T5dMFwHGrVPghMRnEHX5+gdVnBLzqSxHi+zBI8WnvbSLXaRhPhaVKgGwh8KewqIeJ6
bfMnVoooED7CZ0U2TNMtZbKfdIg5h1cd3xw9ItzvFsyEkUJ1LkPN4JP6klJhjXoMTcUaYKDPFrBp
Q98N+9T+uM0AKv382LEZ6BRJQTa+0GtVor+hHwmXOD0q/k4ctxjgJs34jnjWqJGJNspBjODq4Lxo
KGJwYmEWwfFlUhsnBOprTEvmx5o0/30gEPHT38YwpDV5mlW1QtVv8NOWiXkba2FDMZzRMnhYxHPj
zTR6NPPP+nhT7LjaJUBSA50De7RxiqTZ8lt3lqoCgrZ3F8C6nhEcuFd4EsYomUgHmiV4tTwc8fGr
WUn8TPfUKyO02276u5CcRjrtJU4Ox+RMPbyDL39H3dX1GRGaDHa8WBEKQ4EhxkZimA357uoIbDqO
GdlepWY540yhvNUJRtN1PUny67GgFpNWi7aBgqBNZFRoQLeAK8VU6aoUIkKkj27BYvLCuSu6llIv
Q9ilJChanIcKhPp1KmeJdzLAufuBMoHOkUSZchSzTBZWbMZnM5lWcSWqfLSjoI2DU1Jf9HkGHkux
k54XFnDQqRXFf2B+WZA1N0b/69QYtjkPe1x4AKT5hpBsq++3aKB8Lb7U5vfCXVPFxafH5q3AVFnV
Sn+4g5JpiejbkCye3gK4iQUv07Zmwt1zRskVrdAEYhR7q07LixooV3RzWa0bIJbAneykT6F0Vg9v
7gE783pT3wP2wKIRpCg4xRxOnjfSCIqYJJCXr4L4HLWzbtSMG38XW2H7t4yQ1mlG9OICcJpv+W8U
eHxNJwWA0VUzi/269D4pCzXOXGNZYEFTw3weLV7brMi1UgMagmheKzfBj17sOOb4EwqWLL4QHN4K
4v7t+j4+wyHjTOwMBrqfcVCM7wyJExyeCDjuUDVWR39Gv4uDUySgo9VXEaJuBaf0n5MvBLM+Vhib
uq81i9O50pYKQk8HOBTHRvU8wtZHdo7GunilyMZgkQxQXDwhEac8iL5MkObL68X7+PPwGz8PN+tA
uIu008IQhbCl0RWApO+Sogm0u2cj9yQ8rEMGRL1Hggf+Lx7vn+3jHc36U0v/bN0iXlKLKEV3ZMIK
pDMqWYPeOM4lWfJlbiJVHWlKavFIC31+rUKG5WXAAjEfxNdST283PGLqIT3sqaGuLJ57llt/pXlg
N2/Hzsj9GntGIXwPuw9FQQW62CP7CWo9apHptcLa6G6UV9sCt8XgQBOQR5Zw0bZ7d9MIEhr4N8W4
TO57Pg9OAx6jXB5S8SvRThnLZErzw/yezzj9Nb10uAenB28KWe6bkjEyTU282ZiEi7sEIcWvCXKz
V0MZXw/NUxzQA0BgayeQvrQ6yCZOPrMqMKYK/RDs+CpxBJUcv6aEF39Oar2VMP1bvpP34daHbHmK
vBuF9MKfQQhMbw6y9QfGAhmoy3/+pIa+A52Fd+oWimd5wryiLAIGJEOjNp5fXTsfUpNp9gS28zTH
1W5WH67uC6knadepf6JE0AY9Pg09z78yOyol7oxYDgW3dWZrCFlgNNGUyvLK5TF2lvp3pg0cTXcz
8WCYCEM2QKqII5IKB6mYxj/Ao1B56ielk82jXS1tWRs51mTUmgmK8myMygTvzyqiIU8zOkSduw9s
/X28JgcoNnmx6kXu9OVegRmlJoVpqJiRAnnyr1uv4MBK450wlvLewnxj1WpWAUpuZSK4eI9/71m5
TAxMwvQCfdNkIwqL/h+Lj/WHt6F+R3+nA88ix/ZLqVsBRwrfCxLc6lCDoZg22HHRnOS+t6jY7prS
hEuO4F4rabhN/h+O9afybTr9MenqP5JluBXGvSpQnKx2ZK5b0OeJmgKFErP6eb8L4b0ERPMFR6PN
Q66Wg/BwfifW5nfvu8e3CGhq+juugFBOKN064SQHOCatTSTOGBENXK8zaywwmmYOcZtY3fnyFZGT
HbR/J3BOrG/+7gXDiReYLOncLIq+vQHdRcepMd813up99Wa3/EMMBfrbvzoQT11Dqzqc0uGv6pOi
UDpKn8z8f0B0HN4F6uZZVy72JEtudtmz1pCGBiKpxe/6ukpsZg3lUBitbsJdGZyS0AwXzwM8rwKB
/Z1xOT12Pg6K2ZlnQYhT8dFTqE3XIsB6cGHYgzA3rEYIN8VXaclp35ff+IyPc+ZNff5sFCbE5Hcz
xyf4OdWorsshFHTHxngdI6Gx4mBEH9vQzonq67GgG29CvBAn5SSUz/x7h2A8rvXXwzOH4UQJ2rD6
riam3cTDAoVksN0TF1V5LDATVmbhWDqV1dAxBWmelKinqKx0E7+pSMo9QHoXTQM/sPyHYfGG4XN+
Vz/VoelyaZQZwoQyZuXHbrmJnm+Sjobg5E/tBtsanBaMBz55YwKODwgQUbUSzUczngnK44uClFHJ
7cO2fyxMV9TF2Xw+A2ZiagPXBaRLWTBGrOzZnJr/cUJWL2PDFlB9lySDAnXDPxIN5dmq7oTJUaRK
HzqF3Kv3hGjnLPRR/qvWtIAuDjdbB9cGdtnLMi40XpdgysD2IfF/gpZhovWn5/sPBJrjF93GNJYr
dKQjVsBm3YVVs0RMEulsz4KoWj0mjXSjvilN6Bs5Ur5/scW6Jq+QZd2W5wwY6/UA/hC1toxA7QGy
zo0b7DJTaSXfeVtdy9AGbBowlUBSmkLJgO2t254P9ptQ3Saieqol9mATO+SZvd+AhAgChL7yaW1d
qSQj1oJRLnlNplOxzVLSDchcU60BFp+2Les0NkUTeESJ6MKQhwPNwCLSOdaXWC2urZ8Fblvki2nD
NNOCacf2eP1fKKPUFiMkOtpclBq/l4oyhLgcQWcaFFsJvZMly1WK3sTK72jxXzSeAQDY95SHBrh1
4MbFzIW1+5hDEw/8jka5L6kgyeCPjhZGkqfwrsu+/YrjnwCilMPjUSgHI24JlF0UM3Jqln5XQPRE
gFV77DSotECv6/4EbwouXOyz6c4dw/36zuVPUuMVJwLLasyn3LqLY0RvgrKtJSDOSv/+4uxoEYpb
t4tXF/b+QiCVeQQbMQNTSi6WeV+eqZRJCwngQtbfcoOacvpy/53lDw97rmMlJ+xeqEzgoyMiAHTW
mBq+GfQ/wZsu0BzGqD2nyef2bbCxpmzpO+SVgp/ogr5tPW98FsUwMvqZWBoVVAo8ZfDnWsmHxSRn
Uuz9mZlDJQStrwHxRDaq6D2oHazjUh+BKO7d/8biDN67QUse6w8M4ijZb5ydLMvnFjANgOU6EOHV
GRuKTYT4eDPvE1e1fPYMxLuN9yTfMUh+b2y+J0pXd1LxVkLXLbZs3k3bkwu7vclB6w2VG8TlJGtg
Q3zDqM8qmt/rlzYhuB0n/2FP4YOa18FzjTMkl7cqLFC/VeF6ZGGUIRAN150dK6as2LL7eIVZALGl
aZ4d7XCjvUuZeFT8MBCxXAByXAczSALMP10k+GlXhtRzQBlrTXnBDeKVH+96OTPm9Hk0b5klTwAV
smcTpIOXKX6zMxjSX57bjz+pcolJvHdXAjeWIJOjT8rR9iY7C3p3bGGge/+5v8ZKjHW/POAh0b/O
kxZJspEFKHrXljubNjeSuerGcmm4pIKqZU8aPgiWBOVGqq3qlwMKUGPgi1wp4QaA6lb1L3CmZlk4
arjps0E00h2vhZODi638tT2Hq6Tq2BL14mi/RHUwjKaJZsCHEAjFT9HxHmWI+IVBdCC8JlxkzYi1
L6cM+XvP5lrbW9Fay3Plvw0QBK2a8ph60Vs19dfpa87FjSyrARVrLjVavBqMme9QEA2v+N3OZIQp
BbvhAotWpFPIZj5V2yo0i580/gs45/8x3KuGsZFtjIDUvU63KttzVEWc89BpSdrtmRx4s0BCEL8n
7UzzUN7DVsi9PnWcpFoqRtNA+03UgnISSC6rP3OImPH2rw9TeB88n7ug1Hjz0at3Qmr1Bz/Twf/E
RtIrDCnj3AaFkRVOzzWrY+X4791HeA/dZgJ8o+bniYxgYONCbXReipBlUJsH9KajIu33tC05zDKa
mzBbleF2UaeOdZtlbEOhAfAH+/a/m/5ZUqNirikq2SRAvdd4jtjrhysTmWvrPw72Q8ekRvWFIPwK
FAhmZrGINKSrFAspv7ImqzpQLn5yv9T4lpPGe+AVY9YChEa2bkF/KPWoFV8BXpAqnU9WvmdiZy3l
Edg4rRoX0IX1KNvxTsIi1+cLOjTxha42n2g1diywe+JSp91OMlri5ligUbroS7nLHP9HShwejv5m
xHdwrRw49AXdibpyNT3mvKDv1zp/DpTY1OetqaS956Lbn2A7aJltXJM/t/XOgYyYvDMu3Kj2jdGG
IunP49A2xdOkn7/o3LVZu0HokRvnrxoSCRV411ziv2EEid4PoRtu6aa+3mVc3/21sPnkX9NqrwNR
z/g17H9wU5nl4UKXfoDgOiwuEnES0SiR6AdfT8oUaL9kQhTHzQOSNyLjTPXpKskfPoAxWtBT/p5N
9ZQQs45DCDmsSEypDF+3I/vHV8yGk3kCYji/4ev9S8/r4/GcWIbQ9ar+JA5+Yk6D4fglt/4mjz/d
TsehllC1SJSQhsF5ntFYUjPJVyoO6yZ8/0wKSm9OM8ic9gbUD5agNhXN+uNb5p8XHiqLspOWo+Zq
qcsJSWyZOXu7wuZhQP+zJ4K67pZUKtxbg2hAdC2DjxpwOWY/WG69BQ1z6XnQeLb8WdK61DremR+Z
Sdln1dMOGnVWxbfg3DKCZho8/y1WtF1BCxEUMoWS51lLHEn+VkXxvljHokpL1mcmz11efb0tuwSL
Npew99eB0DkpBOrN3fUm194KBPaui8yGS5V7UYw5RJQ5zncPYUQEHAGznEoFGgxCSqA3br2NZ6qz
onKWApHGaTIDfWmjIQTEYD0UdTbGctUHkFdX7WCnX+vvT4T+s1njdrFl9mr69LS3a8gD9bQU62fa
hLKql056M85hBdsJSJPZAligfulZPG0NFUHbeQhctMrshQPQrDHKNQCOl5Z0I5UHLTbq+MlM1y4c
vOAldJUMuLyMZxFCZlspjxaBrtB/x32KzTVrAoHE2JESJhcmuXAXzA3JeWSJ2W1Gm6GPiwEsu6+m
T54wy5dxj3yaKnTTe8Y3+hL4cfyB3hdt5C/IgQ4DrYsC6rDgFaPw15Uua1Kfmn0PJ2OCwcf6oh+K
L40pT3X4YtQjSIu4rKY6X4Aelx12/usmnq4ygE0zbI2eJHpC1cRNbYDwnCUofnOuNXtd+VihSFPP
/vLG/tg14+8Tt3i3RTjduQlbhBdiOxOGuzakc2domQ3dFZe4rBBtEAi2dxyLMgqOep2WbzQezUS0
qMJ0RvhYooSgI+1bVeqOUkV+l6BV+Zp61cza1E7fgDvHhCeFVdN3rr8QrWciYJOdjL82H7aTVqna
lhpUoyP1LYaG3v5B51haVxDeaLDPaKEmyGOOTVHRyIJmEuAB270yc34g/lsxkLv4GLp1TMQh9r0C
QlangP0OTLxYrc+3ydlY/INKv2ukrrluTD7dmOHVV2leCpuTKPzgmLsqcDklydeXu5LeWGq7RADB
LX30qfw2BRZReCjECs5ErXkJ4gWW28aPqepdzcyPYxmNDVccl0CBYky4WLy3D/gKGs2b4aA7Org5
PYJZxQoA18SBJ8TX8XDnzbChN2BkwqxRohb3hSHU8WCYqTqcZFTQyETcqBvabVJDS1lUK0iVwxGd
ZFHa72LU5ZWUPNJThjtbqDNI8Lnwj88SM8glX6GzjVW9hxssBq+wQA+hRnrxz9kpWfRpNqyyPByT
JSwwCUYchyUucwO4lCUdZujQ9aAPrEdf5WBNUG4JIJdst6YgjXbyFxIMusTRkKspPAKkHEBfpAjq
OWvX1p4UuCdsJiTNxBW51NGJ7U1zXw7/Zvj1r9N5qd5aPNV25ko07JFJk4qg8990l2nP2/h2m6UK
mhOG0oCay2uLPWqDmEokJ7qRZAmKqh7jBg22phaTUmtyJWoF9ED89wB+zSGMHfzMhSQjQmvClvJ6
PHhgKNzmwmBB2xG58nYoYLDj/kF82zl4DAEG1994FCpOWweWmgw+paRxBCbG8+PT52D9TLucaLEG
hi2JFCjeN3Bth43tvWJ0WBj4RaIN8GEmRWG2l1OiM//PZ3lyYsDmENxD3+Xi9shi0w4b8zXI0WW9
kh+hGFw3QI89/jzRFIvtJqu7f1M9Y2jkoXecjZUoh6VLp1a/X99vOHyl0iCNLVUXSLwCff6hsv9Z
2iMccidFYaCiKi/EVRx5P6HSeajCNIYcxbgZyibI8tbCD83KEc7vBb/aWzsEuXMSENWgcw517Quf
iR8+EeuKwMyNVga5Z0/SeZ73HPI+01wUNhfXAKdw4X17z2LY4TQ+AxkDuD+Z2fN3xjKXP7Ub7VlJ
niBrj2AdRrUrp/mNo/h0HyZW2ph5FzQftwS8P5yGXOve4rb1UXTRYz94ZNREf9L8oIWb79z7yQ2k
9SOdZoGEF8ASdCUb1iXFGXVZ9CJX6VFo0v80K9bBuoUMljpId/82wQVSIRkT2VD01JonrEibSOcT
hdTfJLV+nMU0LG+UNu10HMyUT0nD1IRpOsp2+6WaYaU5nJ8o/EL7SKvq+UYK29J6S84W9EbmFIe9
kJOweu+Riciw6DOr9drm+lCFxCmub5ndepG7PZDorlv+m4s4iLaJQqO2oBP9HpaTOPmocW97t9zU
VNAtX2EBMZmGEpRHP0sclsqKlcI2mAw+i7enqR+Z+P/EV6im51V0ra6O4+/j0FZgOnQgphHwbrjl
Akar+vdQaxbDCubkIodEq253bbZWxsAkMDmhyAIcn31Y4LhWAXvO1czXVj9W8q64ZbiXpvXG39ee
R3VBmNeedEXz0lE9bUF+/OGBdcuOQN0AOYAhMQ6dBQr1G0nYNZ7mbzw8MX+PNaNVqQYe7Pw7wSQD
V8JBGPBDGKLG9x9x2lrz/wOlomnRkvIwky8TkgC3a9mT1BI+EPfYWUkWviFboDcAhXerofcf2Wce
VURuOE91nt73S7ryBMmRWqWMqorfUjnHI9v1hVMTsSQbSCmZ37qiH5guoimYJpHanWnmQo8W6aU7
cXNYc0P1fegiMY/RqNtanwtGxaBq/5/uLM05nQ3JuqeJ+JwPvEN7NPSU+w3G6mrUqBS2tI6wOGEx
I4Ga/reOOgN1RU0a/Aig/+jwlNwlydrYrlwkWP03VJhPwlZP0uvGgfO1/SrWw1TfZ+hLtnk/LKmf
rMp2xBSsbMBQ9mcLGP4mfsohPBPqCc5nry5gxVYA3/Rj7HJvbjZmJGboaEc2iqYA9de1OCH3exqZ
H/nvHkL3Rdxg0HblgptvICkltpy6w7tNKf8BX0pWOWbYqINGtdVEl0W2wgvYsOqki6Tk2orcnGoR
+mHQrD2JneSep+O3uUeZTowbm8vDBY2fqrJmwvfQLM8+4g/Iqsbg1R8LFTutrgJC2sVIp/kI36sP
p6xfIza45xk793G6tRhJSNi2oez1kGk9v4W+zYwGkInABrDMrbMfrhb11rSQlpHjrLZFrhZ5Q59N
Kwiq9HC85L3RNuCcHsNqGyM8mUMkk4NN+WGLFtHjEd4VXw+2rbaDpvimyfdLtsvQh45evb5/QpEz
5XjAgjBAoxaRBn1Lif9C6xv5ioytel8C1oyvnKRrflDFNyE3MROYakkR5s8ED4Z1w1xiatL3EZs6
qyarEwdkIYw4C5Aa/zrAipfJ+SpTcJkjhCe5og+YGY9hd3GtAFdHWyYr5gYnntWMX/SaikzT4zMf
x6JAPz7IsNr6UeMotZqsp/fTfWdevLBm2zfWp8GvwpSQmFI9W6LAfuWlECXRw2Do2cT0ckzVavK1
/znigt7BO3p13pJdQaLPzHQ2mbClJNGdQqmRktMKPHiHLX0rMaQju70OXUMuvlD5P8YCKFtUXlYZ
KgxJES683Oz4Jl5qrsEhoFQskFuO9b7w6Y5iRgchCxb5cQ1Nk8OZUTLaS+AIKzNUNkTWV0mWCIp0
oFcnp1NVzvHd+3eEdGqPM61FNhCHdfU9gKen+byqgqN5uEmE/rgv3jIOZ/qc/aOMlf6NW7aqhcBw
lWPH/yec54j9w8yqnYf/IdonBbAHn0wmyuAc2tlPoxx1KFmA0RoaHB5IFWG0x8D7kfPrTP4ak2jC
BZza4RnrDdPHj020cZPrIR50E/P3llvVVAzLp28DNQMtjYpWA+K4jkL/Y9UzvzAegoEkKQDBwk20
uQrRIMy9R6uHOCbUgKTa5ZW47TaPiqvAjzsCvQigToP0mw7mYs1Qn/0qH+kNsLVrjnOpBcQGUW6V
kw+ntnqvqk+OWquxXpWQshWS+nqjX/skuVZlH+q8B/+Qt1Pmwf08q7jmLsvPzrVbN/f96DiVglBC
S/lP42eQqokoegidKn8Djq6p5FSCGAJadS0u/MhE7X0kaa/EW3shaXUrU8X3Fv1M1xxAtviUh3BZ
FCorBVPboiShlZN6NpmKkL0XbmGjGzsvYmMkKtYMQ6tZyocmgoAjidHNPnG+0XjwAsv6/uduXDhn
BQIbA/+OKmlfvUGI6eNBjzQvSGYTGq2IZFHvYpiVNONCSUujEKGyyJS+GxIb4MrWWp1GF3OeIKLM
7N8XOfGN7SDZS3pt0qI4JGfsT1EPWVAI6GSU0ET7JCRQYh6MZCPyhKQabcvIqhCbH/bOXEhvIG8j
/cmC9RaAkaKzH+4YooJYJbIJfWPg9AH0VlA+vvAi0vv/+C7k2OqEWabgxlFcoCwu8xKBsZlRrpdk
HZ+tHC07rdje0uPqK568BBERIbR+w0YGHU/wlj5RWOjUuG3/8XzD9W4jZUwzXkCVME9E3MLQifj3
E2OHwVWDDpmEstCke0aaQA/+Uz9kwW+TkWe0cUPQ1IwuSeFUP7l0A6obRhmsKARz/9Jl/3KaSX1t
dtiRW0L11EqR/iXVLOVaT8u0k0C+x2RM0N+urUjZ9qHXxmZid08A826gLxxRizbl5Z6z4EVVlZ7j
uUjlXmYJprZ8JO3UYOIXKd65nQVau2HZGG7/DxLpQ3DOz9mFaC4DTo/HuHXlZkLbn2iEgmXiuHms
eBWoa6JMJt73IxNCa7WAKAjM6l0S2+xF6cb2e9mEXOcoBfTIAdkGDABOdvDbHNvhWi4sK8VnhIJJ
Fvaj+0bwAAgTDDgdNI+9bmhiwTF+LbbJdv+BLgjZS5M0RY0UqzYbFTJidplVRaLJBKOcTKcWkx+v
vwItgv3S7tFhrxhz6zp9z+bHDky4mt5wnhkxBhIPPAMoH08UHOlkirSqlBZeJd6qlJ534Po4zOY6
BegCSywE4MnhOTaeZhTyP17TXXZGiqVjd8EW+m2taG7AOeQIuHbSCHUzoFgQPXA+k27M/AF7GvG1
Ytc2kM56Z/BQ/h3eEqx48AtFCAqYuqqyy6RA4emvUsmyPbfN4x2hAO7ZBFTNFrLITT9aMhJXB0U+
xClXgIPKFkOTcFjcchIHIHw9GPAmlRfb7uu2wiyr7zQE1z0thnWbkErx6ibNc3VVuIVQkIh5B0z+
ojk5AhDX53AQy3FCWDKt1jH7LAeRvF4S4Cb0upO9z4Ld7EpA+Sp67Np3DwSlFs8+D7iVkP0T5jmf
Yra+oMC3848BrdOsVR5xtMS6yVaWX7qAu9K5pIxJTRqrA7Q6cf8rGgoRKEEYOg2r4nplrdidT37l
eXzgL5pjlaEPP9WzGmCh3v5PKbRPkjp+CmI8BW6qEAFiWetjVzCRmGk3QwFrLSFC1Wc2Cs1tQP8A
CTPFeTRAIVyyw3O5xxCvpKs9Ux1bq7/QbfVloCN8JFJk9K8XiTcTdyRjAX/gMTKqo3YiPNRCnsZP
ZgAj0MGWE4BytNWtfG3dO8FeO/flTw3hnh0MUzMGrJcw0Edb+yOc2Dal2r8LADv0JubWLOVgBmxI
YKfw/VNwsbBOPwsmBr9cnstQJUvGOydZE2AF+Ro+hXKrp4N6jnT2zTgAity22zY/JOmANi5A7mrU
yEO+Zrqp7cggd6qgnqXi10yY26IfQApEHHaFzLGhg1k7YwKrHvXmzMYQrzu/dwGthE3FlMBEBAGK
7lMnyALGa5A5mpXfuTY2UYn0PEhOJLqp/hwCseVrtQ1/Y13hUNm7OevFUTXPhvJdmcIz+l+gpMCk
0P7tVGpLnC4e+T3MrzRQP4Q3jpbTMp5gp7/oj/mUwFncyZfYZ0q/jqcyDaeR5NQ+ECmUtjk9mAW9
A0Ka8pKQptDs1tTANcH1u0wHBUpWadi/gYyxreTFCbjHp0a5TxxOe1ohszLI77NwtQmwPlFlpKXG
IRfg7n/KNq4CHgIDWBHNw4ZvgwiQzOhvo39pRiba3xJUZi/iaAdHSe2iBS85Pq/En0xsDFi+KNmt
n2pvoLymFs3c+hE5z408A1SZJeJEzJebxAfDUyifdXlu+1QxDB7LtLLlgm+MlQo7QHBV+b8UCL0C
i9AyEU7HFDUAUiWvhgFgXMkuKPGVB960ZX2l0DTPTBeRicUp+OtThbMfxfgFovZBOx4/BcbGIvkN
RPlGMbrN4z1xqW42wd7nqPp+QSY5fwsoJXlzBqag37cRE6wcml0kIUQnSCxdvv//5TMVw6uRQDB5
RjO1yHx3XddZWneLhDQnf/KytXH2EwMjid6hdydnVjbvJdWnO4TvGD791Jz53D59JoPHPsI73nNE
7e2bDS9XTWCfP/u+p3AzPtlyocDwnVQpGW0eSzRi1zLfQZZV39F0rhA2N2EfW2RFupaLotV626G0
L6m9JsBPs8G9WFhZnqWDflepK0uqGEKidfcapblqXxw8o0HrT3ZqBAuOPUN9pQh7juVoFjVG2Sib
SR0g3m7/dm8dWl6q/jAzG76sjlaBfaAkyvBi5JmDZoR3zXjELoRgu82iNe5COqGWfZMBYeReDbOn
xsewcm1/fbeFEuxYn6WqBtX/mvv+pvNNsh7XXx61kN0TDq/R3LlAyEIDasejtozT2+XW2/ycG9UM
vYJMoBvg+9ywRV0EzIm0ThLOJnvoyEJaEyoez6cZmYxauxdBzYpH0ytOwsB1oyjdBGHErTfo/kXI
vnXEVwOrnv1ypEGVCV8klOkzjqHzPnQwfdlxE7VhL7tearSh+gbS8A+sPMS+F1IymGae2dqfyCJQ
S6WCesmyOr8qa9TEB/KG3mj02DRNJoSDLuqT2WJyqI1VoPXn+0//7zdm9JokhJmqFdFHvUoojYN4
dGEkLDvVb4DINZMRv022ojiwkaytRxN6i17aoAFuMGR3968JzqDDSu5M5G3Hs8VHftzdWdpE1+8p
nIJTDj7PnVuCcHSG16kR6PcRfxEd3bp+Qd3PHRIIGGlHIZqCBOTPOCt7MMIWdAk32yIlw56Xyxs2
d7TE19lUIF/oY3I5qGgwNP6UOylwP0iEBwG/YUf08GKCfbfj9MdXnuFPl+FC1nuz7qM6ww1zBbjE
7zelwfSQW1YJY+tjqhYBKz2T1uPdELYOVql7xlsHpJviNEabMk6F8m1JCCr9X5BP7pPcTv2vFm96
A13UG4ACsX4FgYvAjaR0ESBZNX7N1c7xl+ljo7ylRwlcOfIFFuSOHiwEY7u5y8cRFb0NPfVn+A58
hwTlbAzZxbNoZz9LBOF0kzZRT4fzVsaBvJSVQVps8a/YSuNMqjWh8Khoem7URFcyjYQ7f30KVrEM
zcwTWv1FZMC9cAQora9gkzVkAqtY7NC0XjWdbXY1bd4F7RUI7aYTJQu4zDwRxgkqn1W3Ejh8U3dS
Aev1apNysrKxi2Nj/NaOHIA94XXZ3Bol18LYEZjl/BxjLI1jDnR5L+NarxmfudQo8TX4V03sUFIc
DRXKxvLqr5C/9W+hot2tTIqf4z5Cy15J4ui9DV6t3JPYm1+ARftCgAOg2/N5dpLgB8rAx9BdaIVN
qlZs4pdqttioZp13MA3maJIMzpFwExuFvHDkwCquY/fvQSxmOWF9/8sR+nT0aR4RhmlSbvrH3NSb
OhiVfWWN4PV5r0pJBiO8N5ngB+kx47SpheDigUmsnGaJVq6DT3SKm1S7JGIwoTNeb3iwmQX+V+EH
lx3qpbTC8gcET0iRW9uIAo0NG4QOt/ZZgiFETk/KhNz/+9GI9nsPW9qPYvjhr7UUOVSC/OViSspv
yXVq9Z3cxR8tzT670bcFRZiAp4JKAu+PwMX4QcyWSVgJqQL2H2MmdY9Q3NK7xlSJD+VISqASw49Q
fJw4Y79Uv/iWJp8MDnNSMeGfPEK8cKoTwbI+zwTobvMFh1y0HTCCYgwdF20JO6NaD1hFnneI4tnP
q/mBR+VfaO2n57BA4/qF1/O2UDK+UGVGSnh4jEeZjT8sJyhx5FIrRyaW0HSxsQJa30wK/uck4rrA
nIJ2WDCdPYMOAK7P7RjNqeC+PD7vTd89t3QWLjspq+b4gz1KHLiwSv7uitB+xajOot9HxWKI+lEW
RgdBKEF+2zwdU1Jwhy68uqSufojnKbWtzyIPzA8gQztEB3e5qnxqhgjU+FHmSl1hPs9dv0Po4G5f
wc8+waBbHUmo5aRmQXAtva8zcsUEAsobafHsdIGvPA52TVMzCGZbHSsCMaYiNCrtLJy2NuK3QQ1z
SDwN+wv9uBGm3EpqorXZB/Io75XbwKdfPDs0LegyrESN8curXRNpyyZaohieCpGyXHYLeSpaxOId
J85y65ovcqfNis0m769oCc68382lrbhw+7qJNyIIe88G+6wonRMRj4H7Y8UWWAwRqioeiTIlAAZa
S0Hr7/lx9qFysoHEQkUIXO0Fs0SzC+mMdEyC5tm3c2xgLp8PycfsNBISsR88UlGlpDHLEHB4Pw9T
rbILaQYrWcvL5NoGwOENVBzwf2O/RYkdjKiiktQ4qHYX6HCsFDD/nlsC74hBAxW3HoHIiCXtiavJ
06pyQjoY57WkvETQsw5sExl/gOXQLt9W3qqWK21eCdchIKLqY5LlPEBJQGbyHcfIUD6cI2Si5Fxv
+5bM0l55rt0Lh4eRAzARWwu9gqflkb94BbQCBjWGqFgOvh6YsdoQoMXM5+M6AajFsDyDDqAXoiyy
Ub2+gfhGIkSBZFLmV7BnTdto3IurPpbvD6c2XlpODh1eQVKKufMvgXp7AaOvLE97qYkdQf04PrfV
ZB7bNPoGtDY53lGTsjSrMlrr39EqaBqzeXVQfnu8p34sLOLzIK+iKZikW474LaBBgocoW3Zj3WpI
9gZPVx5uOv3pZQwtPHzMRdRNtXH8FOtrsU3Bm80bdTGCLzJeBlH+vtJg3xikul0paxQp+ukeuZCu
P22KW5p3xUc28GHU6KW1wAn29RN6advRTsisEc2PKi7fSbWEaBgY5O7WJ0aS/dw6UKW89h6aBLDk
9AwSy6jn7g0cRid/3Nkz6LjXQwpqZtw0frz8SdeB6lMrVZSm/NsF7SPj/8HXQIsYCyyKVKdP1baF
w8L74Jvd+o9xEfA80sMyYgUir6yFMgOA7ZsJdHGmVfe2IMnw87YNjYdg845iSpxXJXcagk5OGX2F
Tnl1/CI/qFyh6GQ+FzpuYyhLUA3MSDKmmk/Dj1A7Guzrngx7rARiN+dGZtzNm9nB68EnDAy/KTv4
oRA2ysu4hr3yRZCQV6pNm1vMWU6Jd7CBG8uCfFonVJGlLBqIKyYUgSljMqiHipjVqLao2GB7byDh
Iy7BRUwGjlG/7kwCiSrJGdx7NsubuhELQYcflqk7MDeq4dmEtKujJo+jWIjKifpk1B7inmjXa9S2
Cl8qXRBmsA9k2B6pKY5qB/uoOwMKlkjgonRPZUcuwa/Z9kmIAR29OtBgfdWr/DQcLjY6h3SNQCKg
3LxqftsY57fA0lsVUcZSbxmsd8n+KgQoTboHHCmJNEDou9QvRdSRRrs18ipXoHwTuMunK91eASHd
K0gUV8GPrkpWuOK0LCNWsqXLlEKU0LNUOf680iDrSz/wooiEArl8ghoh3Mt3zWMiIZO7pyscjz1w
XDw2DuxWSlF3FnoTAKLI9dupwVKIPwCPvGd8+3pwV3pjQXezqa+aDxV2b4ujGBBVFUEdLAVxqZQo
qwg7l7s+3mUVt1ISh20jTlnjfksuCx5hlnES1VNPvmYO3W28wCkpT04KuenO+Gk7TJoUscpJvCbE
JN/mARXfjHQ7/IhBh2cnkA5iGpwt6ZqAOIGKPd7cxCcrV+KrFy3iZtTQYX4zhZ7yUG/+v60deDV5
z863OazR+HFwzyd5VTr00auT+yWGMRDbPjPOeTf+C8U77ANoi+Nqau4wgx8wU9T6nCqnOmXELZ6Y
a5UzCPIjq5Flc51lxbEDZDokL8eDxYlm4yaQNGCGSMg/iXSakgrHS8BC1Sz1e42AMEd6zp5dW86e
9foKMOgWHd9CDfYIlvCrlBmUPKQQIVA27Z0asKheZlJF5L1O7tEheuxPSUGd+1ZHeYLiyMnbZV7g
5/8ZDoiEDp9N+QyOFBXNmubZI7bkGSl8Vh08Q6lYPSL0mwYT70X7OaI+CzA64c2eZh2HXm5Q9OYr
vjyAqeOgEY3k7rUh9eUQZ2OfBTMAOHaLVdG72ySUMuqHxYQEGiBDeE+6b4p8M3qHT2Q8f0poe5Jh
jE0WV0xZYX3S+4fdHWTFmAUHUrCuSn9hyyZkCRVRhZvJqq+DXyVvcubkX63Ab1CdbfCyi5cbwcnS
OyAXttXQYkJo5N1JmzyS+ea2XymK6b6VIBBTHeHlMPRQMIOd9RYfmU4owxDk5E9dln91LL12q9hA
4XwOpqRnFHS4f+R9DfhxZKnb/svAT+QEkK75c+vlaq8eEl/6GCQ2lgeMgE33tFK482k93Dcg6TeJ
wdQn76GW6aAevbPULLb2tEbTHeRkbfN03lOygjPEBYvDZdBaiug1d3XDvGsN4xfvouZcVorG6UgD
JNjIbSbonxJL6bVpiPwvq+FQ3KxQMT+4AXGlcUbbd045qFCMaWdtpXgLyIsCeer+PWJLnI9dblxX
Ow9rlVcXV1qXmr3hY/7/rvJRiNeH6yIsfd5QgAxn2aNH1A048LivBMur8Xj5lE1jYkkUgjz/mPaQ
tFoHdJM/NFfKVCsS7rcyCEZLk8phdPcIwLjizbLapMlbEcSderS3oKZ+f/aL2KzQOlHyyMguopA0
pyRhTcAcWdO8hM/O9fqAOcvYzVsG02q3ObHY5Uwq1qSTY5wRgNpki2aCCHBIL0f/b8sQbOI66f8a
FghmE3yunC0Y5W8NprjEMNpnxvLQBjogZpKqRZDBbm9HUghpO/Agofx8kPgdL2kiWoVcpGMINt0S
ELN3n50f1Yafgf4wc7z0u3xTO7F5RHEJbMypAh0jBCqZknh4wMprZBwJacsdLeVIRQTEMPJpwX54
AhRrrDyNQsNMDURLJUGaEJm1QnXhRTtiP3xOlFVC2Tpm6RxmVQMRY6/TK/FvjXAd7OULTewo65pF
zdiakrUN/6+XxIAvd3+6cVLxD3ACoJ98abKeG+WcUZuPJG2/5E5d6vdiGcz8pPtbZgUxcNIZtYv5
ly3eUU0bF0nQUBiZrR4C5tKsgFnyajUA9JlT3y29HYEkjKB0HtfKaNxnY1FLJAIdaOEtoCejc7h8
KFIU1SlgPrd7SWklMSWENthv5lefkQYkQeNt3VohhFppDegzZWBLjYKFiPi1ZI3/Tqg0AmbhPUp1
AlpUIzOOfZRuZ79GFL2MVubpucyab3B91RZUGGTKojgCZf3VZDUYeVtLaST9XIZDwG8ITa5e67ZR
MSLrq37ADY+HGy7Rm31RfKC7NpdcrOQVQ7wwmhihBFfi1Szh3g1QNfOfE0xjcg76nfopwZsoez7D
T0uvXTkuZtMzUbBypXD8U5b41dsEe8bId8cpRLnGSDR/0vFmeFXa1tSeQ7XkOI4kKe9e71YQxd7U
MU6XILz/sw7CW1sTWlb6/NZ3FSD2j3skSNXuTODbWHcaVxwKs81E40w28cMN/C3hzEZLD08VE+Ck
rYi9eRxNUug3m7K9a6FWOPt7Myk9tZ1sDito4/kcD9jE1ylCU/kwXo3Af/i6LTqIeAOYfjcxwJKJ
Ez/ZAJXXn+S835RMPLjlcFb5h/cFVtCPIRHrK3vrXx/4GWhv1nbFFb1FiCKCw8Qj3Q0LQd5TzPN0
e4o2x/M9GA9saqnkvquSsqae1ChZUQaYxEzHm9/R6oFwWS5V9/+iVy7VFSk7+dw1YdDpjTA1CgAZ
zyD0EbjgOsZNKmHKYT58ft6L9jpIdq5E1O8oRds4CGtLaW/wd9qEywp2jet9LSJCirAkI70BlSAt
VbBawWFMxnS2ajJ4tnI1mTy+qLClIuv0IcLzdjd4tLLhqs+TcwY1eb8x9zZ2I4U1ICCaz+h/xPCj
49ZJUT+A8TAJrc5NOeux8cK5uM/7Bg/JIYpeRfctB54phl8dtOBnFGuwzRj70XDiZ3pOOAa5Dk+A
PUGrZ5xto9zRwPlpbCL8PoXDYN0fBpdZRoQmp3q+g3odkR8W+ETGCawZIouIPvnsEcXdAwXhB+tn
G74rD9nuEwGM/kQj7iFVa5UIaxFxPvUJ2WwRfnRYkX5bKbDqYmU7GIz4WQ+pWiZjDjiZlrR6Zwbm
NRTmVRxF9a2z6s5PKEB2aOiut69nDrk7TyUR/l1MJVVDo/ZcXxjtCIoGW5wVLvc94NSyFmhcZwnm
ZfPjHetKVoWHwhJ2CzJG0G0tPUyuHxWYmOrh4yvgZYQK6NDVGvRCvHUiMnZ2vVzuoM/oEfhz/60Y
i6tlw14RQE6FvkCTmA0dIE3GIllMfUc+GTrZAt9TY+8EVz1EJ76UnX9BsoiXHeWVZbQX9IFFGcKq
sp2sWd1vPNWFxp5H1hlANjALjBrE+OA/OA+Pwuetg3hWNzcyuY8vOcfKYYH31JWIdHeJGaTKLvf0
2OgmqWrfHRS0XbsLI6NqiK8nNbEG1+vCNhOQgSH9MNUH1jcyOsUIS+nFyeKXc5wdaFMugD5E3xMR
386eg+m8XHJF0Qx34kN0lYrAiS/pLE3Qv5zShrgdeSlwIZb5NkCezN4poj0YiqiAxwK7fvsBLbsZ
ikkg+WbAue/134RHHfPEx3qAiMUdi237sLUyYLXoaFWL+hJ/0fjqHUP4Mi2D8mMIRFkl+Iv5155e
ii0I1jYdg6dzq8ZfUiPH9t2ncbos7kvYo0GAJQ8RCNUc9SHumje9dmMU5kfnAdpifF3CXC6aw5nc
4BVxiyku/n+jEfJtJA1Z0fu5EKlE53wRDGvWm/d2fdJc33Wk37Dtznfm2WrAaYzt/zy8JkcBIU80
Y5x26DmkyQjz6dewWNIpjN2SioRtdmGe9BXkJ+p9GGTFqZFpSA5ehQjp2UdoqXQtmMvtQJg4ipl1
7HnGHJQwKiAse7tUtRcoi0dljZBck805x9Cpy/F52jglh8MmxYhch1ZoLpkf26xhbUCCtMy+U/b9
Et/WMLU6d+Obv3+USGOOWnC/K+tU8Pl1dyC6seNQg10noXiGr0ZCv+2bsEyfyaUKXrTxhEc+ZCmJ
Hc3kqqv8rXC5yJwNPB2CyYPt7+TTCnSOQ1grm18Dcju2zMag4vHkvxlGDvs/7/YCCPCbFFai27t7
U1Qy6Ec0br5V14qscXDTJK9frRen05uUPX2NV3sdsecSzY2MMeV9WzLzg9HfqL5dh1qV4kT2hD64
64gzB+iivfCU7yVuhqgbhDAtQae+RNtDQ/oekPU/qFgs4hCKvdgBevj7YEwDDo0o55I/X+R3OjVJ
NtHvcGBCe0InfGhHN8zuDRVIiSOgDE/5Kv7PCRU3yH8O9eyPmZx/uURkYWqv3O9S921/ze0AeEoI
0ZwtezkrKJVAbRw5Cl7FnXmeBdu8twSvILVBxHYbuOWBekbrKT4oGU+Vd27D1kwPhLufD/wrhYnc
V63AiQ6dqCF12/FhkqFX2Fl/iK9sVX/A6tHnqHVLkK193R3YaHlsFi15AugysOoAz1QWGtSUlX4v
QbcaicNcdwQS4KzK5u05j4gyLH4/lWDqgcgdO4rZSqL6Hm5G2QjlfF1teAJN8PnxdACtZMaVwzzd
jZeI7NTV4rKCr2p8QvRK0jbJuH4+C3Q94MLTKuEELLKpnxHtuxy/yzLTUMovZHHk/knSh3gEwOoF
mYOQ0gzhvRkuTKZL7gWuwM2EYo2Oiy7S2oGiaP9qqQSjkYK2DkAKPvy653CTkpBoeMws4PvlEEh8
JBvIGs0sXVvgrFgR/wOPqY6t/1oIzYwY7SAHp6J2/Ga+J/Cnkl2nHoeqTIF65BpFRgj0wEuhY0W2
uWc/Bat8/i4eRgWF7l6pNsYNkxCTPqXO45ilNcvsT0XZgXhdUXW/NXlrrLn/Niupedgdal4S/zox
TqMRIwyNMFi5Rex9rGgkfgCwkng5MW9dSB62SMjwWpa5pY7qPRaozXCrTVbiRSyQgA1O/tauKOUp
qU7Y0GZhtAasLR0jTcXvK15n+FhVaZlWOVFDdZg+bQ0c/EpR96njYe+z4fqU2uPVRQBgeSTiRUAK
MKf3I5O8ejlGD7WY02161VJ8SMSW7tSjmYpYEAf2aR5nPUQ5leSZBCPX3FghSdbzjn+gvHjgiIJ1
n2LYDVT4iKV4iot2Gvt0ju1MY+2ASqqfGxorhpbY2kGGvrhkcKRyw9MblufuI/wYhx8Z/FWygH1E
gTerJp6244DnOUFQBm26yzjl0JAHIM+NP1ETsWQxlPNy9FEmu4q0kN5e7I+pII6Xvp7DLmJdc2Dl
YhN1cnr5IOJGN6bLHJBSgrpkmEkp1ohlg3BXeAJynWniJIaR079pX9/IQZJPt+sQ7sR0G4q/Wrrn
QxPLlblS6vdUbOU4Kb7Gim80sC3wtGmad2gLrfCj604VEpFJ+mH4R6Bg0r2rL9t2aY5WXSStkz45
cKPMrfDehViHVQ2nwQ7hHzDXND04GYvjTHwmzF2jbQrlRT7tEzrsKNXnUPiWaaa3uzyTm6ExElPa
teRB4fufUARW8zoOXaSCi8X2I/9ACUjMRjrHjqT6zebY4hl5IbCZi5x5LmihFq++Pw0InuEu9hyp
7db2ANGpD41f7f32IZWrpUWufkD/lzf7T6CyUSrjV3H3AS/HNFDeUOe7TTJykJWw91wFB4fxpSkc
aAHizt+uforQP/Cjkr25wmLDcskBK1N03qHjcCcJAv0eu9+1Bh2OUF0lQRcdTcaFHtQAxpPdsiXS
zP3C2zM4cJ0mIQ+xEZmMTsMT8Ou+SsMpbC6PJN4N3UjAPRZKCu14QBTpxebYz2Z7Mgb67rWRi8G4
+S3QBV4LxuLC3NNbehoLYyKpKF9BIlY5FLl1eU0bZ30tFi5SZbif5zo6Kd2BMF22QSvfyIjMNaJC
drAfHPfFE/uq45B27BSG0QeVGoHAZE1EJGfYe8rE5YuZdk1u4ib+cOR8Pij10EvC48VKqSh1KUWQ
1EJtjUB3CF866o3DwppJ4SW3xQ9Z+pc4S6bsiy9qbgfoiMIBcld7hOfxMHdzcEUgjY6mjP/SImXf
jPy38VAwaVoiB+UJX2433eh7m/M6+m6o8E2pq7qa2yBLDhmAasQlcbAHjLBCQzIi9SMFaVr6MrlY
pqUH+KYu7Pe1fyPd9Uu8Ddx33it9CljUXDozhLUUZ8Laz49U92CCH/Y42qOopVtKw66J7/Cyf8xa
m3vOkD3FYapwUL/i33TxFMCcd+7hMEYhMO891qbfyLtBRzRrv/xg8a5MuOS1jLuqQyUh9qSwNcFM
3YYYd/xhGVSut/84pLS0xmIhUQ+CgqaMwGjayA0Ow3iNH8k8hNoFxCoD/BUbY9x6sp5ZOxxmrszK
u7ryVS51jReUAzT1nCpMyjsFgk+VMcuD1OHqmO0jGGm9wAOajGUiGNj7CMSYPhjVvrWZO73Hmubz
zyluc5YEBAlOtC6m/OqRZ+2MaiVPkoNqLUcKk2wvTFGPpb7tf8VIkG4Vr8gxLNk1wC9iyM6R1Pca
Kvzr8/Kk+oGIvgnQ7hx0gUxDrY+a6j2uEEpvjOCYHf2IgsQK6+iL5mo3IpMPuHvTI/i771ErBM67
uzzAu/NRgf1A5oCiPAdIbWZNG9J+BWhGNsFhbTi5YS6R7EkPRiE3JKX0wTfgFm1sIcIOFC+K6K+R
ik607DUkTbBlInP5rSB2Ki68wsezNsP/RBGByK27fUx6TsaQwu6GaoUkYyNTifYnwwMurKIOcS1t
MagrFmU6KiHezqwQHBe7uGDxiPZ6Op/6qiX3pc2UWhbaR8KqOBapub5+hWZjivhl3ZNzi17S+9BD
PlF5+s/JTgUnSWUUppFsuvyzdbJIYFCG2ZiMVtAJtyo6gYrEF0McMJUAKZsamGurzaT7mv/iLg8i
dD2/NtobeSgrz5Dy8K3ewHf4iWI/XQ/J3MzNVmTQNmWBhRJDVGRT//hboJzpVhsdr058iPSD1Nec
z8J5JkyZAQW8TQ/XQQkSsbIs04/y93+9yyYlSHgV/C/J25UBAVClwtQ3FGYXtb12tGGInyNSI3UL
FfC4T5S/lO4EhDVcSZgcP2Z/HxUZMPmdKDP8oLoXcaMk62S3QW5UjMTu4ND88f3h3VNP38/YhPYn
JddhsrylljEjlkNNohMK5ME+z4E2gEi3AnBJTdt2VdgxlJtkAZFuJILSc8Or4rYQBUwCclq1ytcL
RjVq/vOh2vi2YyL5Hnlrrcm1CBFBgQN9dhuR8KIbSNWDJPG/aU42+MklFDjzBuOZIBeojEqzRRk7
86BNnBk825jMUbbknMPWwzq5xik2GBPR7SNi6WgTgl4+E4q4HSkhfl5SStXAXOLpAIZBe3CXCm4D
61TiyhKZsrN1KCmQTEfcpe0wF6lLIEvRxuGEGZF5Ja+OkU/dBVdw9tX15EcJXf5rp2gvc3KYwWNo
aImJTneBRLccO+ydFzYVfYmvTh09mRBVNOl7erJxmXAcSRgapDfAhtHa0eEW1V1vG7h2ZIdOE784
1IKe12Pov+fYmBZdEf2Z74eU3Wvd/OBUUp5qXL3ZUwo5XcbyREy3XVLHZt9X9twoxmxTM9zTuu9D
v4tyzp4UYv48zg/DqP1ly1bmXXgUeT2qj88m9zxUFmKkywEra0idlPxPAbsvg5Wimzqh5dWcqvhW
PENZVC6FdHq+tooxG4EZ5yqlqkJyIFTGzsljz1ix8hfLdOXTZwft+2rr7idly5OZUqKxdZ+U1Nk1
5gz49clDeoWMPVfF1S6KGJ8xeoV1WLndlS2bS4UlmAovpWFvVTJZZcD5LY+oRXsMznpI/s7C5u6Q
t+jfBu05Geqa8ShUEqwYKYszo9dxMwNctDIvOY0Ke0hHdNSAewfrVJSOu9mwz4R2VOSuljAwdmte
QtC9tFgEYhk4Uhn8x72JXO7e+JHQrUA+Fvl5VdhbEEj3uieRxIhrzNDCbKtqdvoSQpPcEn3H7E4V
Ry6oC3N1LyTzZ1B8QHgSnOMD3iNlFJ8xizv+ErHuvhZBiMhE0ETkIBbGHgbWsogREuCE/hF2FkCq
p88/WzYoG1iK6az0h/MMkK7zdwfEg94aMiLzC/vFX+tb/Xu9MiAjHz9zTdr1JumPAetwYrb8+UpI
m/rqtUR4Y8AKe2M8nPRNuqSybOaZI3hhZyFgGJFM9roxQAxlInydbsTEpbmhgFdLp8noOAcG4QL0
wgDLAKhhvSoYCBHmcp6LbATrrVM+2keudjt4uk07G4DSy04C6FK2KZx35JggRtw3Qw4LKSHDDGLv
yeSaXZ8PYdNGjBeMpKEiZdf6LyNjV4Vre3/J9Qd32upytgK6t/T7e62BPtETolnfeTtmMjA65bhq
dLqjnN7+v0FS6yaWsloQCXjutVz4stBJQTpFNMPHLYMzbeS1nTw5MLFJ/LQxw4M+sXWrkFEfu0aI
i/k4edHva0/Loh7X/dsn38cXaOkEDKbzZr50mMcD6AwF/H3gwQ2riobVxJOGe+PrcvE/5Gt4TYhE
G9MbMH4NxycvC7snuyDvH95zodoyD6xkIaVCcynm+nlFI66SJCQ3f31gv6N+BMQWxKH5qcLK1E/4
2guRIw5ctMhhn0cY4CQTWFX07TOdZfGdJWwnmTJuWINCNkmFzkRKRlALtPZn47KUjcpfXpz50efn
pFUzY5cFQadoEHsuuE7TQ/J9DJJTSdPHjY85qsY4qHeJ45CpFugdthB4gr6pjxGIj7fx3UkLwjXg
fsZx/Dkpn7VwUBn0MITxXzzTMz7LABcDgwLe1/kC07VekTevynmVfXAtK6aMH/Emq7+1BNfBMdgZ
f+mwkh3EWPzwuHt6oIVgx5K5o6VKrR3cILjy8OEFoewSwmFM5kCZgGXytBbbWTpBk/zImQxqQMJK
ZLAQpziP3TySqeMj1JmolMu9xBgvwvSnRcXcRE44znYBMWEtO2R0D+8KtYjUfEDTc1kS67HKM/w1
dbF4UP+BB1t4ddu2whILJXvVG4PeZqidbEUOWOCwkcgdTWrUWc/hAns3iCWGRa5QJI0gpyWGtEcY
ooNXhgiTyqYrbLoz88apISp+E3sHN82to08dYbWI7OyNoh7N+rJmwwn1izivtqWJQTazbNqG1EgP
sH1qVtMf22dbG/XAzYZRdR0d1qa11AixCULWIU41diI5YBAMb4EC9ZRM8oKnG55lCs2omzEyE4DD
yPjLoKJYMv4HSKVZZouN9ooKK6jb7fyuqyKKr1m3GiJep3+j7A5ew+X46O1UXccC5XJtwFV/AE15
AhyHiKOGaTTIl/mKswLK9gsYkwb6FdsPieqJsKJBVKrQ4I5Lw8B3Z75Bm/aUiuXFwi/UHOn7R9zS
gNHiCL8PJ7vDu5QdfhZ+gA09zySUTcCTMB8g+p+9CGaQTPisgbkPDWjOKMtXbim4CYhs2NrHlCfl
AvpfH/wNE0cOWmheScLbI9kJnMMZrv+NL0n2net+lKqwKcsfBMtSZUJ3PVOyfqj4uJ5EO6pp0QaU
G+q7JxgilXae6ltJYIP3Ht/byT53LCTitj7NV21Jkz3LPYI05RstTf60m/hsWXmUjpqorKeAkYDk
BNNUxef7FXdx27qh3dhHuOotmr/O0nuQL9mvRy5m9OvqQkcfZjdtqxFOMkChs2H+nXHwhIRsXqaM
+kVhNFV70Yif3QsErSqK3Sph/9Dn2MC2CqZKHU5QRwaZxP7fLh6LgEkcxTACiTYHxLc4XRboAREW
bwnc9nLQE8OX4Y7ccnOjTXdKbm/MQGgxNcKzLG0VkwEupH/FzKXJDANBSsycibPfOqHzVpALPvyr
KrPAc1EXxXFHC561hL8GMNYGA/0VlI8yybG80e0w4onr9DRyJu0N5Ip2i8cJiGOJ4fqeJM+gBrjD
96q/058jCRjzDKY+8a+FfOdYDNnDVj6BZMiRR1kFcw324B31797tTcxFDPTQvv4bYpZTM8j2p87r
dhoadm97CDzft5F1USFiwEyeReTD3sNyyrwCSQqVJcxRE1wY27HSKV0I5x1TLFtksIVCc81LTDmw
THXILOCRtudWyN6qsTqJNohHgKhVQRPDwHpg8CGe6mtIvdyPCYDtHTJUK6Dn/894FJGp5ZmiVycA
jjBhBbHsaGDV2SN5qmQD+e+26OaI6gjPekQIpjyyJXAqUiOSsZxGaWTJ5yd0YD0E56b9bok0RuDR
nUth0o9RWH6/R4t6LcZVrz5kFGAgFIfd/oIAy3biDwFAQo3JE8osYVh2rqJugWmR47YMjvJGl7qu
nbFsBOjMidbI7UvwYzGgSUs47X7M4gLQQpEg4oObiSHwV89+bfrbcVxAtaCb9hUHdKinzCwevs6j
Xiubw4jX/xRT+89/ANsQGqTtPuV1VROTtb8CDslv2k2NxBm7NM7wADG5TarCAy7apzNSxzrryoMC
rNleXw+/ndrxPjdhDZlMeqRpO2snRIlWknTeYlBaIOstRLAXiyZRxkT16/TZ5YN/SJF9GoBkwZYQ
6i7ZrY9QHXaqEg/320WJ7ujnzDYCaw0/mBH7kfXSRprCzlY1ygXZaA4GwMdlnih7tC1eqZc+oAS4
QCYEoWA9rNZg+7J8bErFnlUJAxkN3PXKEkbLcCzkdZYzKgV06QQYsDcEPc4/Px7Z8SGW1lsWecnL
OzqnPwxq7SNd7XR00eg0/bOZBqWJ/p9m/xbBUKlbh5J7/BMERKyw7x0TNOlAc7i67Cuyu5y2eMmR
1ogfkbzhUI8nFO5PTmFwdLo/3i/tc9zyep88stl6JwOx3y5Ho7u1CLyqGRvXOLq4VLoqRXzgIMsJ
diS8GvgpHpuIQY/m3Cb111YYu45eig8lqVeb6bT8EQww/IUkpp3gYRenlcuYGvg2dx29HGpJ9byW
VY61fMw281DFuAZ38yOX0ajb3UPl/cZpMR0i2+oBpjvuzAIMnB/veZ7yIcLshlJs4oP3TrqgIb40
2nQqhCLhqMuEqxXoFW9LlH2V8wBem/HcdAPAHbhLECW8TWy0MTgrQsNjHmiQYYczg0TV5sOZJSdB
9ADE7zTi8+oka+DV/UNoKNSUU3GhbnRJEPqUHiLIKssdDZSpsT9TSo/qlb9PqqLpc17FzNDiCe8p
Gk8zZIZ/AxCqudLomyyq4IgS6c3YaLD1MCmqLPLncgJYx59q7r7xElCStQGbh+D57pL2qIzCT4PY
0qtTo76Zm3RM/wEatXK3Zl0ksolm4kkFGD3dtHz/11hQ1h5b3BSuJh40tvDYnP9JwzUNkk1yc/s4
OVMA/OCzJWU2K19RIm9sBvhh5wTlnM4nM3uzXrIzkTs4qlLBdJkNIGqgSM7bpQY2NkPxFVbHAkHI
49ThvBMLkOaXw/8sjbHiXyrmRjQ4wWWxwN89JpqGY8dYwerb6PPDJ9drEqtgUAKF6OUBvveGZSi0
BpjM0Co5VDnzmjYAtJm79bDF+oDfAN26LG373ZDT/GumP/Wrt1usTdenECx9H4hFZIdmz/VBqvKI
tshD4CDgBA6ujctBxub826kkNdikl6tM8BCK/MF4Ou1EV1MdhuHanNXYEqABuAHyXqbUeLKoQywq
kBRDv8c/JRTAVkSqwFQAI/0sH59kAbVpy6uvy85KBJCOv22tX3Rv7SjXNj/lKWx9raVC20kLWJox
etEJTh6AfO+S9Rz9ebNFZCEVCpywjOVCZd6ljQ/mc9TiV9p3UxZ7L8MaRf7rSf9KKm1aXcrhfjNM
GvLqr9toesplXnbXdWF4YN8pOqGvhkpThGCfDUonoNoe447CmSp79fNFJj2ufnOHi9lF0q0nT3XX
KGbRD2PWIESbfvdXXRoNSxe/6A/58CRC+C6lHD+TXP8IlgJ085AU6vyOjxtvarLS6k+mzk4N7M2B
TVc2lWko/MjvpDLrmKSn7pczkGPIzKoaZ6OeZ7Topxl9yLQh6EUVSu7F95Fxb/dZoTh5SpZkHtsV
Ui+H49+iakmvn/itLP1s8K2/Xk8Wmxu+AwhzdY4/OAII4TxP7zlTQIQy0/ra4U7AZTGyw0/YTlY6
ShyAcnNh7ChGc9nxn854PEX674NWQ/wqrH4Ga3AMnEd/1MdAm/XEJQvhmdI8lDuUncDi2oRXNT3a
pWJVE33hthrurLcCPZmKRIx1mMlCkKzqeeN7UDV0TXZeUoHRz3ef9//9TPO5E6KA38ul9lQxYnwx
1bdjrBcdr/QJax/DaNKoTGlwPC3xdc8ExP8qfCIDWx3kMqRH4ck0upopFdhLUob1GkQJ7/PGSMXA
XxfsTs//gdQDUe4vBcKJVf+TyTC0dvoNJYX/WzXu1VVr8+Lt4frKm/Vk6H6nwzqDs6XL9dwAZJ14
nBDvziaTQilDm6i+i9W+3BfG8n9e/LhvkltIjjvV5OpD1ZB8JTFp7QhhFs1oMzHz/cT2Ts3k8NWI
mX59ganq+mC/BEIH7lmV7UBXXzYcKiXJCew63NNwGE5JFmr2V6g1sSm20Km8eXnkOZoFhRSJed7R
z7qZ4ZAofgKM69l0vrpQggPMPp/pTVYxcpjnub3wtojsP2b7OVmS9045q/Kkx/tZ1VNnx1xSFGVu
PQiyt80MI7FAQp/RxpgvIa04SmA4uVv0tQi2ocpvuuFHuQQF51rye/W/a1Jh8m65n5gpD99b3iCX
RKpmBhoL8xHcZoNgVL40e5rPBvOQD094vyOz62BUH3+BBQ2A3VPJD+fSIYUQvnvCEv/4dwrwxdn0
uECvr9/OwVYLAIDEHyOOvIBDCIh7IRSnkVOz/JSxogYSEHolSWI1DiRKnfUsgoJ9wY+iIbqPyrs9
ZGErtLc/FgrxbhGp3vWTQEO/LI9p80ww1a8Dab+c8BcwvrujGDI3lk26rOt3VFGxoY2h67lXi5jp
Y3dRzFhsyuru09MiDRv+xNA/aPe0EFi6Qeji/podHyasuWe7wlAdEv62Qi+rdoq6SNI/cgDJeWf8
zwFp+ctCwNHbuf4nFhJYWoScop6LmqOFLtaYXdLMuvjNelYx2PhJMF+Og+BpEY2jy+RRl0d/MN5w
gb52mr3vlCRnfgDy6q1INb6plzGbryawZxwx2cLPvi4vnoRCqSPfRs4cGWKmcCGAd/WkgfjZKfvg
whnIOjC2DXpBwdGiXG8KG4nmEhtGlwhL3MB+uY/UKKh4DkTCXbbWsvFjb5tdifdMylO3vPH4ePDf
QkiPCm306i0dz3ovTHGTQNAApVdCzofmr2x8sU0LvGyO0cVECPRQUHlBtnD43LkVY1rGyvRRr9jU
YgUuYwh0h5ylY+6AWAP2I52GevHZN6+62SLLjtjQU4TEiU9iTmw1JUmZszqsImmJDm44+gJJeSA1
a116v039B1DolD5zspkolsb6Y5rs8+Es6PVC9W7oQz2iB7cOdfcRF+AB1tGo1Ah5uFoC124a/VBo
EMNvGy3lIE7vFAu/38UvwQkelaQvbSC4Or8xav0ONv+2y5QXyrQnSzizsjTpJXzUyleMpQJXQp64
ojyKwZJ3wTtK6A5333UrB3sk/7yu76qVpsUhI8LiYzEAggp1kzZ16LipOuvQGEISBRJEeaiYVX0o
S3+ih1/V2a6oHZ+hfld4UebKR/sTuv0jEOlpkQSZw8PxeyVV8rQ8Jj+w0/IgXOmTtL0avye7bx9X
EFWWnpuXScun6X3K2MaNzGSsjg8mFUQbrTw91UW6ryK1hp8hILS74cp0d8gPWLLy/6Z3LJgtJuT2
W2CWyyVE8K+RJSyNZFkn5XGJ7GLuDBHd8t05UKlrTMByY7B6uKV3eij1I2TEv4ZSJwwobnGKpIYz
4S44IfMiD8fnDyWa+7ov1XA4xZSRaeF0CunYS0FQgH8DEwbr1wNQH9UgpJamV1lfiRE1+k3rbV3s
2OGeP1reLSwE21VEFim9bBJUxy7d/3nt9hBvD9jt2jG6JeHL6qyxPQDrO5SSRzZreDk7k3WVYL6z
ONj0eOgwrt+ee+jWHauZJgqxA2lYFfOmamzAFjDEUQDKHgUvrPRxRSKBRSbe/HaSMPtc/Obi5n4M
yCjzp4rf7kgl/LC2v+9fbBHSsrtmL7JnyVkdEHbMJT/fH+U5QbBcgYEL5l67SGFsMMAApOuXJsH3
iX2SKcX+d+FQwMsTfsM4D2hML/b7cdsV5x2NkrUx3HLvQII+e3NG7GYWYFTuBejWrSlmjGp/bIwA
FiFitB8LKw+6Yxs1Z3+npeS3cHl+oJHusPQMOH/i3sCn31EYvAKOODwH9DuiArKlj/Sbs8sVBkeG
YFvE0bJMDfeBDDRZxUcBfoY+CxYMHEoyNYtH9ZIlbGuLMILyhimKoPZJYZu+ITrj5daZVMPWwdGy
oaG14KphuJvqXQcN+slvKe684+N1Yt6lPrfszqrjXoFPtyOtSaBytkfO4zQzlHYHDJYsPt9TD+4K
kMH72RpRKm4U6/fI5o2xX0I19rTChHNKocDuDXm3qbT2hjRTb1WDq60sSAlF1aegRIJUomr4Acuf
nD1z6RjWptamH6Rf7ITAUbq+6EWynXWdp3UG0i5RwtWzQxVGCPKNvceXOJThZWyidgOUyQFqrc6J
ZkMiHA/e1b3axZxjVy/BhNdQFe//mX2TtHE+H7UhyQ/Iq9AmLqK9pUPgUWDcxgBnm0zEtdYfwA6t
h25KOCxWUHPMBE9PRr7nEutT7w5uUuqmEQ9UedB/FVcZqJ8NX8PP+11PhN2dHY5kk4J/L6Q7HVlH
faqcojhEybWo9i0dhw4BT1pQ3mGdMg7b1y9Y+sH99MqN9CuBL8YVXgORAgB7Wz28rlIG2gjEyOnq
TA0v83Pme1k5F8p2yllm4vmsv8uZZQtut6WymHBn4d3jVoLVcKY9AwUUTwRRBdqVwc5kkE1SI1vS
PG+y+vW4evoaz24sSk7FAji4Z/ojUnsb1iEsVYzaP0lUJqIrJ0q609U4rU8kFsJyL273Z8gZQHyg
mF1CzdqgRZ+HVcIAOh4w6y52jz0LpiS9YwhpX0sfMEzdQ27Rpfy2TMrLBicshtz4g7wxiSIkD5UP
nFGUPI0V9T5fZUrv5T5e/xvjNyBUCUmzYlQY6EPSwauZz0n9YahlQvD/JvqLObEhMwms0SJntnUI
jxoL29x8qi/eY5lPctgkptbnIpTmgy2r6ax8XQ5ENNYflEWFGTPbWwkEpJMmUSURAxfJtPiPJP1n
d30Fd4wN0PEK5f9kT2Z/1thxTZrQk/JtIsiOGvKFLA/voiJs9jH1tfgOXVpOp48BuRdwYXvm2riu
sdTWvjcYFNQnPqiS2l3bNm6QxL6o41b/1z5/HI/RjtYqUqFmBBQnYNDVGlVdnSrKPys9LQ4YyqFI
UNskwFQo7x0vqDWRD+xDqv4xREyD5haDATU+hRteRdlTVHi+Duc0bWYiFrrJjZ7ZEF9y0H7jEihx
ecr2R1sT4bxrsEAjXM4rc8/22J/cq1bjf3QABdII7sCxnqdTB4LmMosjcTxXS8rchEwMIibcxeP8
45RjngOGsXuwgXdT+oJWmwTy5KE3VANyI27S+35Vn2BwkNecM3cb0AmtQKFqCWHpCsOJ96x+PJVC
O8lhlUCdo6OuvLF0k30cumriFHy2pkeg2HmWEpQmgBZVceXLKMN1rgBe2E10XN11W1nilikvcD+p
1PUgWkb687lpdERbLTf/jBHYLSxZ2RCvfDhGD+JzpG9NcjwnPVPgrlUIx2eSp6OxAQMq/FfiZheP
h5V6rtG5Du+0fyVb0ZcxjvQ+9H6ja64kR36Xm722ZTS46UJp5/54gdIqL+uZETjmWyo+iwEQNx/A
/EdAgss2opJmAj0ApVtdGQPNAsfi2NnGAXYcZDh3DQ1+UXs9feR5Z2zW8hZ/8jgB34YiyQT3yyLw
JHkjLtvkOc/ZOA4kiGIUkM0rtgSDsmbM+uUtWQ6778IWj2RRJGKqjzrtJOP/wk/IhCaEWqwb2TIR
TFq0906O8DFOf4FXsh7h+Hv/WRBq3r+oDIPl4iFcWkjRUko4S7ra71w2N3vRq4Csfoh+9porQLh8
QnB5/3mb8s94HuVhYLGgHT25EnKj3auE4OHVqQuREurjl8Ul0DFNJ3QFn/nWcDyh+3qrYweYOd4t
mKcb5cjCz+29BlZ9p82XL1aOwETUXVtZ2bwGHOLFK/iVhcVhEce33/hCZvgKCMxcABUaxkHnLcyj
2THCODQgEuyFMBadUyrNXMXsddY26mMlkMFCQzv1f1jhmugDp5pq+yXcaHfjyBorcFUtvBlOaeBi
ABIG3AgiBnmxRSyTHFkrL31ZvOprSBjdl4lFOz7SnPcTOSn/w7PzJrh81eWUvv5HuBxxM1Sf0hLt
NGvySIjPuOQfcJo08JFd3NTeVM7QqSHGco8eo6lFrNVEjsy0Yed5TCAgBwKH/IDkLckVbK12GSCI
Gvj+ArZJjBSbxsOeHJ2HFJ35VO0DZjE7AcOHD3SLLdi4AGG3YeOfFQjbVL+IwvAu5woD1octDwDu
O26u6Kaw5+0W5JKf3Mfw+DazW22TNzwUWSaM2nfTykiPw22YGNb7u7CEDN3xnfXOreQrcdNwSp2P
dyLHCWkNRffOGELiWJBMGsXhDF45HyDYk0GlDrfzjTv4A+M8sN4j8GNjkbGiZq3EWWCel7FtW/60
qsmhosvWzxQDSlaRn3i26supqQ1HNQG/aVwBFbOhbGpb8zuMGi/czPD39kEFG76bylgrwL+9udz0
UG3nzRWeqrVRPz1ZX4v4GrcWR7QmV1XxwtkDEIp8fAfmEgOYdgwW3YPYIvQozP7l0MumtUtTewzU
gO8qo24t/gSJGKzVm9dzSgt2839SuMgG53eDzUm21GckAPwlX1iNjnu5BveKhxuDIBLE8llVlryM
ef4dt0OGEHwKjvjSte6v/cUCvTRg3rrOAOkz2qsf39y9afZer3go5Gg4qW2Em/tU69tSnnexV36Z
G70+Tt1cQfPb/EknhtEsKNfPWwCxBz5VL1f1l23ZRe8ScVyXkDehNCruq+uSxflqQTvV28AxBuY4
/dgCUtFK6rsfHdy4+ZpGfcDyxg300AuhM/nJfiV5qfE00Gu3egKOWz1ckmR8GIFLGaPe2ywmTi5j
7PIxUqK2TLTsoBItFQcMx9mDeCyfhroGWDrLY9WbCCoTDYv04zoWcRHVUT6yx7LewVg/hizPxGGe
OQ0pd43GAXEmNB5wpXV7brcw2slybubniGI76rPGtCdl48ctFv98v6FSFxtp7exGwn7W5TUEcER1
rE5wArvyDwQ7hXXhQmf+Xw5rUCulGTv8luLTULLN0QQ5w4xzYp1M5giqMoVU+FhadGFP7BBKVedb
ru2PLPSAI/+eiVuxL3wh3uzLxmN8RuY0tRs8HBuPUivTLJQt57Z4VJe48T0V/7uzpsWgntC0Y4ZF
Q8LQ5baHOv1r4AceiAID9h5JO+5fNhm33nbqPe7uL57UbtHwqEboLhATcNOgfq3Ls8dEbLdi6dNb
MfrU+HS77T5A8N9bS0601GtMFUAb4GKOxR+BaxKp9P7EwP1O/1wbjlVLkp857JT/CPtS5zovg+PQ
rLewdp41/0vXN6DC2+zlcZYYh058+etu7DvTfNXV1W5aBBv7fPJ16D6AyCBoSdKwAU4H9LNixw2h
QJZceQEx9FPNFjtZEELxOe+F1nnkEnkyK2W67vEcy5csaOE8nyvU9ztwzLF2Rc++CVNTsdNpLuEW
Cz5aFt0jgkdgWxTxLA+pH+i5vqfjY/6Vg65e6fUEu60K0aIwIwYGscZBIH9w2+B/+7zDHSgj+jqL
tytnbanpihIF7fCZ9pWVwcgkNFbrfS8WEmqgmCjlRRu0ivvunyqnThBs2S+hynMf5e9IMqT/F/W7
UN/K2rrVPrTCaHBU3XzsGmtWNBE+MoYHTvUm9L/tw10l47cjthGNBBn3lVDLXvj64iRb/rrwgBqD
aPc3l0TrQKoIiZezvrM1Fo9sX+cunOE3FWb2LoxJs5HIEM5McQROwtlzzE3wiGwXGeCzTmJgKkiG
kgguOR1dftugJBYra+EG/bIyfy0ctZJeXqEPeq9hKDQ1xsC49KRv1ttpxsLsCP1iKvCmgPJ4dZXf
MG87VWlDd5+WM/JsTjZ0nYS7xLL6IHZ4VSEdV3lNa11+JL/6oSceuZtEORBWsj6tzLbk10YgZfQH
DlsQfgyhk3NQw4MNLf0DTBWBbUMM9Yr0mCVVcKDff4xk9dxAvxWFyLAmMSR2xP59YDHhN0tagaF/
NbSGJy8pNl7sIu1gxBLC4s8+dvmB2eqHAMmOUHug/GYL4pzbkbkdOx2H1iQY6XUfl/NFaj9kyn9L
KRooa414YneL9gRMsKBhrAg85ZMPHX9NvzdoiuipnWd0fnJ5OC230sKOCZXPXnrVWQQtrWP9g+W9
5UzAJgAKpiDrwcbw6wvOgHuqE0V7MareSsvX0m+9qvxhdggMGU2BN+rthu9MHYAjqm2Irbo9qZ3T
UegiorzN7iUaMKQJD0XBizZNtzB+lvuHuFxFCUqeRlh6DdogL9gbyU7iuxO11NfcHz/MzWEsGy+H
hXuKFlWp6hpAMjfnRc3Uhm/lRPEfnYZQMiYZRkuQukqzlglFMx/60t40OZoD7dUWCg2hK5pLF0TC
AEz4A2rJKJNTleajMqI5HccXQhYyJGojhH/X54xzmBfcrOJ1kQolR1q4WUGYJ4KTpBvxa3nYnwbZ
VXhqEptXYipXbX8qi5fqCbf1v4As2DWTuShnFttMlY7LzrPNbZTbrh8bxf4qxA4wxhg9pXqUeCLW
UJbnckMZBSCLXpDZqdcXmyYRpb75nrSVammeRKTVY+um4GVJt2G9xZWkRuKhjYErlKWuWOjuDeVB
nGXZ5gFOGZAMuHcO+iDMvrVc/zN1yIZyzkbJ0yA0TsslY+lk3zq/3ow2D1Smppuwe0AbLwzp3+NQ
SVwZvetuIGzs1ow1WcQxT6JyeX9QXB6YgozH5y5cPjRIl9zI0N4gC0lFL6vbhj0BeGmYdkOaxrFM
NXFZeHrO21CbeerGx3za4wXz1DTtWx8717/Pu6TrWCq5ZXBsZYJQ9ljj1CGpBecIjscKE7180xFX
uoH4kFtx76dfC4w/S2vfPzHg8P9nfu2b07YIKQB+CiXcy6Eg+DQYV5tIphMbpbSFvCxcbZlF3arc
zT1Agp353yLkIDFoFsRFf97Z3YMlLJcCt1G6eunWBWPczoxLz+w+QC7MwtMg8jbA0qs9ZEnrUib5
VJrVFE8k+K2k9BNEwDzbzIHoZ/RrDXDOaKgZclRg0dwLAkm8J60mv9yTH1aBZsh/3Ffmi3DaaX4d
/jBqtNQnpqN954OkcpljXR+7khQ49jWt5ZRndqLgxXmUHkHtGWuQr7bpu0u7Oa6av2/0WIqXu/8q
Qi8VjRU9NA5NXExp9PNpLIu9+m7tGvCASFXKHy3dpxtB7l+C0VH2mFpvruhHdOdhV51UdH/pRHDD
rvLYzJ9XMdkCEDPIJcNf2EenNIdCa95/aky/cveQlrCOwBl62SUOFyHSdWXsp8vvf3pjK886M6aP
3v+jt+QO0Cr3mIOEpsCIyZmcsuHePgMe57B4eovnrCsK3vHv5+vr9c2hHyy2vzHWKVLYEVLFhtnK
ebUg/zD1jSCE8yu8Tnzkhw/mlbG9nlxx3611mShFCknz4+OSV7/I7vt4sRIIgg9Xq1/unscY6g9o
ZUy0kT2u2grCRWEYkSMt48irZIT65QQNb6ULvhn+rVcek9nznLkZW+63dNdu3IAEc0zkulhAe3q4
0LNSnWkXMZukZbyx6N7hxwKLsPdv9CnSTpZzxfTYUUiEZ01MGRXYZ+eNBvC3m0OmWsv6urd3e4ZX
Q8bKo65uMqUAWgYTjhQxHu1RNgDqdxEN22vJ3RmKdOheCoOLo5Nyn8lOmMvU1QpiYGjCWNm/irMI
fl+O5OEYQJvYSbGpg99W46LiqSljWIl7qLRHHeTqs5DYpTKAlHSMeMujN7on0b5pLxprS+Zd3tOu
CtZVTlZiT+y4qtr2zyWM9xWJy5UFLC+lnmIdTbpiQwikq/nqvkFu/hsv+LDJpZLaV7komjgBaS6l
rTfImBqftpMyPE7abf9p58yThXdK+6VH/4l2x6X5ooVFJp9nbukei1sh0z/dvSrdjb92YrcMxAYX
dM88T9Zb3IJhfSPGtG8y3bTTLcQHlV4Iw0KqBJzWub0lvhB5leM908npH0NDJnMtjpdWa1klcHZK
hSS0Q4RjP/AaUfcBFVr06Isgp3ihwBzM4BWvkQqO/HpEK3Rbcu/L7hTctjzWU/MzGJLz+NnsuipG
JvlcjjKrq/Ee8YaV2crS8q5LLRDrr6oMvMjQTUaimN5hN6Ykiz5hJydU8pkGr5eaW8XQWJxAF5ok
x36sX9PBJTZpxzWlbPAbfmY3JM2pRLXYbnoV8EukWNrMY8kpqDt/HWxzXTVLdQrbVPdxaqiGBGb7
z6fDogN1zR+5jSq3HW3dksDIZUQcZn3hl7XfXRWxLO87etHlXug3rNxwSgtITJimPSTnXfYM4bqM
/YOaOXdadCyrK6mR9XrMAJsxzAG357yKsCTF5rdLlrYZLmDPCuITlvyyRctkvCiY0g3d6d1RBb6t
HzH+14ESglBH79eqWjMVX/1rruewcmWTBHwm1lDref2WUXyhV5EBsc0gF8wzOLeP5erDS2lZ4MDY
3/i+pjjcg3Y35tvhPiMjCvutAyuQcFfxmamlQ+lq5GNHL2769ZLOo6jCQeKe3ju2C925eDfCCVto
zJjpPBwrczURkxWMjWcy/oVk9w0UNqqfMzENqdodoMnmwxwFqrMH6FIqSnQFrvEeKF3NG2+Ez4rc
UR+k0ajyy0M0OjRlgL9M/I+PR69pov3UrSbxkDCEYXrHltygLF/5LMy8eARxuIDKiwBmR3NNnSSt
3JBsG2vxfwa7h+KPaVJywwUbmfIEY7Bgs73dG9XtuuLr9JtAcdaxq62MH8gu8yiarx1YaPQ53bh3
HVjdRTSS8swaUzIYZwwUCUWwf4wV6tOkH452JfWNegghzv479TA0S8qsjrhLS5Pzq8NOuIEOGPBK
sBAR49kbqxeoKXl9Q7ZbbzHej01sscM8l3AzEKdQp88u/ek8uRHGvdVB/TOLLBkjWEzoBtf9WqN4
vI44sYTYxSFnlP45XcGMfjMfnPmEm/Ffl//y/BxdZ1w6gw1e2U0zThdQ9iiHJn9gzXp5/GYx4A9x
1nqDJuTSlHfzwKT6u0QlSVqJkvZ0x2ts8a60C8nQc0tWGEBDQWhQza1K+UlPWDQXC43uJ544gGKS
ex/fB7Pjf4P1u5mqQhkNVwOT7+yzqi8FRf7PEvCGSyRXTv2lAKkIcNiTF0FbyU6WjYef6fUD1XL/
gELvCh118079oc1BGyPs19XJnuh/2QfUSKcRJTRKLjfjNIGLc2cSlHVfyCKtV+wb1nWwNskg+Pwb
fIBspe+96j7WaxrsHEVvjDgNQu2Cmb8hMwkNVMyXDbhXAq3Is3q4to50ci+IdRKG4is8Z0328XeD
T5OjzrqqqU1JCOKZBFlG1Gh5Jiy8Tt/TbEdWpMmPgocYCtjRGOxSdV1xt1CpgVQQ5zLCIZSwdktg
cKfcFcMQEXWCMK4kGz312i36euSz2G9qwJguQltEtBLCfVel9DtvMvTI8ssqfKHCcq7VMifWkD/O
KL5XjeUWLYLPxM7wWb3rfpJsymubirvHHHVQVaU6qobPexLPipevS4iNS2GGEZMhQBizoIWmPGsG
8dVDCjm0JvoTG0ZVC1KZ30AJdeIOKjnRVBIlWVZOiAdqEStdhoZJCqM3FX0235Cxx7ruL43QjzoC
DYhYNHwhUihqvdnVj4a7B1SHL4RVnwp11V+Kbakc/w4///6ga0Jy3g63F1/+fbyhZykJY+/r8G/0
ILLxvBZ3TuJVPpvq95z0Rd83aUYx5VJykOmtbJBaWA4uP5wrwkNoe+YifacCRY0tCDpyQa499/2i
JzXd5It0oWjLnsNgoxHjUwzQthc4QKN6ElvrqzcrEp67V9eL1xsoZhAq3Dbo0UYDjaIhKn7mIVql
GaIjW+f76bvafJCgWP+HdZSSFaGEFMK2MK4jIP0dbKBmhqF5+tkRC0lvY78E6/BLni/WBPwnz7Pd
tho54lSEnDeMpKbwJX5O0uZvnEC9fMkS6MU1MWiqjAyCSHAmntE1TU/yKiIj4+u1jUfBn7jKCxTj
oOynupfx537sMoccgl2fOd+ZiPePJJvz4ah/4P2gLxsZOV0iMwSaxUcMCpwVuxVRv9mZLp77URFP
a82719t0mJVE2XnfWlinDTtZthLq45GvUnXdpXzRH0nE924rF+kuM8+5y7GNyNT7GWevomf+1kNx
EN6bTOyPSV5CESQuLsH2V/+akPriCyCy5G6gLPVH305TfUrg3IImShZoM0DF5GJ3bGSVexoM38t8
O5tJjqkpHchWTpckHVQgM7e5xnjx62Bx+i/LFcC5y0ibTJmDV1LHrjHGV8gFYl2rvfwGNVgvWsn0
/fo/Rmv0J8TWF66nIXq3eZ5+M+lzMvs2fTxRt5G8mLjGSEtZDwlxgLfIfAj8yN08TizmVAz7TvAp
bccdaqkCFzWZXpPvkpcZbXFGzRoc0GgOejsbb6l3hSjADpt20sABxD68C4DVZG4lY95RkDYJHWzC
r33Mm5y1NC6x7AGPKMxwhLc4d6NeKqKAPOEKUBOvRViJi4NFQMSvCxltRSPomnxPorXrk0ddfy81
+mF3kvktzjkQIPq8swWVKHIArKAP7pCVuB+UDghPFFeGykV/fOvHY99WmqfLiskYiH9l+4bPor9C
yuwC/r798zg7QT0CvyMSub1FouxheKROmk7B9JNDNwnDM5GIVdh86qNwSQzMW4Icj6ZMJ3KB/9X2
357ZOUO+Xewv6ZMME0oMsODEzCdPQBN+PjKF8LNK8psXZ/PIoIOeN4tRSDGYg8hPX1263jPIumDk
XCrEORdncL3xnhQSqVKbeP02M6Zu4Mo+Rw+wO7TX1eFybCYRBGBl8PgQwpKzmRyRIboOg8NNCFDV
U1ug9mw1ljxrupSGJhmylYQoSC2QFH4hUqmhSUCedp5Cov8ZJzJnDVaM2Fla0UDpRt1EsOaGMZUq
TRwab9EiOPNI32lAfsZfyBBb/XFsXRpLZtn+9qEc+ca9VbwckosggJ2XkWRzhWlg+CIIBiy7LO0d
2cKxksEHNCToj1Hlci8uRujTNpg1Nrb2F+Vr9FsVHIRvQldm/0UB1ySD+8l9CjSPDkUgl5LYakgO
yQQnNgDG6DZcosBtDjvwSqZelbNKgtk1RR8DuP5/sRlqqBPNlJfJZx6Q7qnJh8/0YFg6JzAK0yp4
sB77+w+7xGT3i/W1xLxX/T8+aPLvWs9UNHoCWQrZoCw9nInqxGafzoWNfSVU1sHlA3Jkt9KIkBHe
1D2G0LHoa4dT28ttpRWcSnsZmYxKZSarUQbg4BYlCiHmxqO0x7SdfbN1wYIIJYMbRESGsqTw3Npa
MUsodlHaERdfCj1WaKIAKAXUgz0itTsmyiftRfXawV+ruyyHNd2npeUpvfgXNvDvK48okjh80JyE
DpwznyUhZ/c4ILyWobAimwnvOUmkEVEjdU5HqgKralPHrJ21rt6BQhicXhvgfGDpQM9X1TFFdxor
dTJK6ocQnGPtp6u6dv7YEs/gum2ZOISdb+8TrVDB1vM83+GHzWnz9g6IKroHInzwp2NnRcv7DSPQ
yUTS037Wihy1iBUV/fY5Dbl2wS6TQYlgjsvChE5byMbvB0MMVIy/H5I1VFmy48y2GJzXpt1xHXBi
JwzRBw7DpmZevmEkUOUG6Cpaor9bTERGvyhoImQYBrRmTqwJ8CauLgHQkhV1gZCnjf9uLQj7xqoD
HHGX9U+1JMyAZfHljHB/2zImMHLmpqVpZ57RTHZE8G+sG0mGtCRTyvUb6urd8mi71XaeqIFXU3I5
kX/1LCeNnKYZrYB0dXf+Uutj7Yx5JEEIUZp9qhF3/K8EUHTo6WFzOaqnrL0Def5j2bRafstx96Ed
WsSKWUqOtW+lMEmgn9qmDIA60E9C0GW6LO9rrKlAJfEjStkpZxUszJdNCOUawhocOe/Pn7u+Uq+k
KGWgPiMzB7RMgVOfFoJQVFaKrTWswwAC/smkxhb69ASJI+8ih1aG9cd2jx7eTVowZ3+7XRx3Xo3p
PLC3G3ibOc6vwwZE0cPK4A5ryjl8BD46WBiIuC94r/pZ6zl388kbDFeWDDEFS6IW2Lnp3F9u9mx9
cR4IQfKQB+wP80AOGrNqq/31IiGXA1HfTdBTWS2gPHnfV9YAUgNx7KRtvnwKJSmauKZvm7cY7mTU
gC1BuH3t3GnBDn56nSCq6XEf2nkIeJvSKg0/aCuopFh4T+DCb3ZMJTk0s6urMnuD71QuUFN3LiPe
heFSEFbWOYXiKxYsLtK1iqo+6TZ81LzflWamvOhnPT+pvAXzirHxNKUI4+X9CS27NhMcFTBEkcoQ
dE1DrEW91vDC5K6G7wx6ZxPYeIca7c39R5z7oz94mDF27tEMuqjlRBjYxizHz3IbEuBcZ1al2oFR
LrH4oJ/QPLM5vUPLkmpkVY4ZbfhM4trPkpK3eLiZTiCfIV3sJSam+IAQZe8CGDl4G7EG2P+R8c0k
y7vhXCc0VvHq9C0jEyiRT37LytNM5K9XScBbFc2ntzw8hu0Q7X9A4orMqUIhs1DEn7g1qetqrGBu
9SH9pegEwNGnq8rB3UAZDbh+b759q1shTdPMkDrDTtgUmJYobmHDrNXD4MQyD52rgld5qvtX4U4z
mCNum5i3ci6P/2Mvv8uKONfWkTCrnhATu7yZQIdVxL3FhHItIU3JITMvuZ4dfj080QTTMiy9W7Km
hkZMWKgR134ODHkTZMriTnt3QoT7jXcDJnOrwMjPBmalPj7jQ+wM8R12T65yYDy0UHtfNCIoCuO2
TAf6LZsbz44X1idehPNtLqSdxdhCjC4nKLkw541HezRiHLT+sJITfp+ec+bdlQn33RzlRoTac+HT
QbyZ4uoD3z2Yrv0PR/aTrv07OVwldyC2warSjQmTZt/c1yLIlLxMaAeXub1YXqbMiOx/eCAxeLwx
qH/ffaglU28cU3L12azs9ycsP+EeGUNmEnwPeybYjmRT1pZIqDN+axbPUh5GNhk2sK7vbviRKNQk
wIpu33dxwHShqPiHkzVhkAc4udyN95h9QCywcv34v6cvkxCjvGyMtuwtE422IytqbYBgauLg/gnZ
eECBTqSDFHXJ+ycN2X9XLDBBlelg8kW32MqyLspYikYYWt6fx1+xUoyJz4S3cNeM8YlSnfKmfneM
M4GsUowhdASRM2Y6t7tt5tK4USjDIhlNtUgasqSS/A7H1VpfbU+zBUct1uVp9K6DQauJ5j1JKMjf
F+A12gYe/kizO1GYHjuxstpl/jtDOZyudVJ8qE8ACHjFqWhjGU4HaSNBUi0kELoj9ZTNfLySoEk6
m+KJQmG89Q5U3HBlDXOiRtPY9sAzPjBf0B65gvY07BJnnudGlGReeo3bMZJj/HP8Lw9ccJFRSYxz
QflQ6qkYQVpPg5a4Uw/EFqIIxP8tKydj4jNJO3kwFht9f4LFkJUJYDe/M1VdJfz15MA9aDzq79fr
iYlujK7oVUSQ9cCY2KNIifNkKuXhx3tEUWHY4nTYPTJhf3u2yB3sdk9lb1/m1O8B/DeJfeLvgWrP
SQe6tXhfSa9V7ErDnrEccZOflM8G1iR+j59vnBKn8dlK9TGcIuVmbp5RZ2+nY8PMvp+woI6b5xB6
G6R401gu9InmoHD2zCpTbN63zbhrylWvTGgC9g6Kz+8HMWDeObysrsl+i1sskoAbz8AQYeQVwiXu
3yX1ZjTVdCX7QkdA/IzgxmL7GUlafTZgrAh798JUA44FiiGiGIlkG+zoRyM6oL9OShs3L/dMG7ZF
JCCVGoXpcVC+ICaiO2BuuItacnJruUimTB+aXBJsAIyTbCu99lsdHD16bEH4E9901AImsI+7w7Ol
cuwAt6CaTJcl3qr4K39k1yJiZjcjbaqfj2FMY9prdDaHpf6RjZB0iSxjlfxyK/99BurEsnxjbHhT
k/aUwJ2xdJ+ZYGkmv3s42eX4b8+h7JoKUQV3olIypv5aJtw4K2gYtrxCbHoo1pnq6TT21vkoqciD
okac5p0mSUt+wcnxdf80ZE9QhU3RR5uEEKAtFqZrBucR0ShfEnhc/HQSx6RnkFFLQ3+pMrawt9mS
vrHoFqKlQXgqLMOld2pn1m7xS966QKMbDM3J9ha1nQhckBArPEsbJHmshu+NUJ+H3GT+M9cB3wPm
DUIvDMxC9cjzhwYCOF4xMOUwgTbnx4iCXtTfyQjjaFYdT6ifCQxGoVdaYFd+w8Z0d+QIlwq+yIHY
X5cnl336uTbKeHsVLgcqjY24PWPgCjqyp4X/gaM6zssf+kMt28wnLRZJOUn5QFeLXug7hyLbV4Xi
qGoFvahdFxPKlWRhfuuz8ECkIdOhGhYICUpYGYhoefQYQNamnVj2Ueaxtn9fwPNuAXk66IpkakII
xLu0KrNroVG0CS/GqsxUOGDYJ1CeipWmkSsrT5My+1oeSUQaZ9PiHMxt87odd8f26BBIkj8wBNOv
/Y6QfyYrGnp/7eHEkReyd45q+Cqlv8lvmExKqTIFOBaFCi52jLHVXiJxt/Csruxc6jd/NFpgO8wX
C8laOs0ejbWQxLDQWwvkZ3vtCE+TMQ3pGkWdjil12yWMxAUxm+6zeQVWhL217L6YB1P0iXsjmQ92
zHAcdgWcGDacFLe3nQSkwBrszGZH5snJTxfp/Jfz6SOoWBjVYnKxiGa120I7oYmDYKHS73pyJvMj
IpB0sia2nhD2AaYw+QBslwbUAU7dFB/wg96QN5mHk6w+anUgIZ499E9yotpZBNLZS955/W3J3jd1
stYIYbSLtIwowMlBhDmRT/1G+YydtGJE7QjOv5CjDuSnKsdjbjcwLWIP4WEXbSgEAQiC+FBSVDf7
fmKxMI6yf/fbQOo2v8p2MZGLqrOpjUSXQMya9Q+Bzi8DjaLtTZ5l4R1+XhxFAgFOc05C7OsYjv5t
nXji7MI5kqpUXocy2KS8m3hVwoUeJ3gXMi8Cm9G4Fg0zKzAkPRB71Wm9jPirA6yRckFBnRfyCvNB
LeuJuiC6vCWjHXd1FIAgxnC8nbY6qcfANCdzgc8X2vzEqIshyJ3Su1fpMwuGPViQc5ENMC9+TQFf
F08Brmwo9xCbtz2ETWzfZCtkMo/vW7qUxWqo3+/ZZxEBlPQAOjwC156/FLPI0fUwSsY9dyOkAaOi
hccs6FhyDuKEcK6MhrMdq0I1HbdLDTNnGvuU+f0+k5OS1HxRj7AnD+RHyvys9MKFOC+tAUDWjnTF
ELlZeywvzgV52jBamfEKt+tcdCffSTizhJlg1muy8KGIrqHrvUDem5Jusk/0TQUsw1lWZBqsOB+q
bZnVNl3BTf8yJsSAe566kIPsljQLQaQkQgjNBH/Kd15a27FIEpsgLdcQwK9PMHUeQN9CwwoWoWO/
ZbIitf6zEjJ3fkGwg2OmoFTGvFLu0aQvincK8B8d3Pi/xkZuzn2mJbaaNlpFuYGBdahSSynd/qtO
rofTnED9EsTCMutxaHWBQKtBqsp/2YLaf2T9mqVHdl7tJTSA+cB2BspAOvKSxlKXZ/GJgVCOrpki
52rmwYPCEl8k1Yn9CjvFsTADWJDUVkfOnbZ0FoGVSaQX4hsLHf3kgu1HpKbQcSHkDOEqtgnsKAt3
MydXEtNTINkCZoXcBdhTezUXKmgJGz800H6DC5WUSC0jfAAsOYu1MSiHv9ffiBHKJRhLzAUDbXjZ
l7+OPSFPjn01svY7ITjqWk5a1OvDdjCGFtk8sRNZxAKCLnOmcRW86LFueqw8bZFMNILd3Q6gmgCP
Nz9/EdaI13IaFuCyuQbyU8p7j8E5bR09XXcGZlTsHlbj5nEHLum5KBK4itQzot641UouSw3dmlst
PLXRTc8FEmB3ow0kr3C8/T/MUwJ+WASp1MhGNfsG2dBUjExBkScrUAcSwkhWenYzvhA2dTImiryy
eIPiEIT3o6qnomnfuZQK7VUafq76olVjIrRo/acrQP5XELUedxe+o9OeCKgfOMzM+HImqdftouC3
tahuIsJnK+H+mVJpdehNdv1WUVVZMxI3BJILOz045jD8S8K7D9hWZgXj7y9Z3+KdbtBlaGw2ylf2
rQdqMKsIAgkahVJr4SG8EeyrSLPUNTMZUfuV0LJE3jA0WVcgovhKBwFray6UKiAFpzjGPtxyOY8O
UrpbkgrTqq3Wb9v/6UnKUc7HhPOZYB9HuLXJsY9t+Iv7FRpqHUlILqNtj8eUkR3N+n5PilemaD/c
fgND6Wzv5784AsOiKBdQKRwtRbYsZOFr/8B2CMf9kxrLNbmqb4W1tS2IifoKHHBEHjSwXjv5zI4b
oRqAiiQug32ynHT/pTsVedMNL08a0VIqzCZyMYnN9AoVnebO9yUbyJlr7XBdnxMfHpof+yyYPIxh
L8i2SiNgJLZ446uJwBtb5Gnh60/OzQJljzqJ0I5c+neoCbif4t/qjNeVDC/dc4X+vEsNDmVOIAs8
uIMe5AefGI9hH10LULWThWdRcRUGvVboBuAz9V/fz5S0Eyrz9eMmeFHOVbMvb6bi9q3zfbGqOyOg
r2KRV0bvm3XkYn1MEVDZ3F8vkX6p+eCJLNINimx2d1eL3pJsnp+Jgvfd8ERPCYDVE2u9EWF7Xalt
oauxHiD3y1NdVjRcE1dxWH7Esis4OEXhNgCRUtvg+JERBjPy0NuZpkkDQKD7sOUBDwmmkYh0Xsqg
Df5bAz73Jo5tt51XAA9SDM5YHILSDkH+BcI4wtCjKmQ85xcydEiCn8Ux4U/c7psr9gCFm3ZazOu/
pgLEPGJAh/X1238WVBYezppLaTaZEzOiXF11dK2/CgDVc1J5LFC0WySTK+zSf3bvnl8YDAIcE3Xv
svmUk5n3SrtAubjlKQWDKI6zf6RhMdW9CIB/lCA/TWOagof16fOeQkQ+JVQap51Tlp8RsbmSrROo
XXiNfg+huHl72WTyAYgp2twV4qeDBLe/uIQUtF00ThMD5jVMpiqOCbET26lwzAwlao2wdOwho5Qh
kOQti5jc2xpfV4PyXxRIkTXD5jFbtOiGCFd/z6uWdQXHGmne4b1dmUtPusZc0ivpt8J8z2xyxAJ4
XcfUpgPfLXYmKZ/0zVX5YeEBSiOzM/M4YFjtZ8Tk+zPXALbL4DBKB3EFa1uNuYyJM6GYXi7zB96O
0713AlSbmhtY1l0Dz+c0+h8IdccFjBKfA84wvFKLYT4HzmBkz4UzuT3d5bgIVd2FYMV9vKtp8xq4
H6Gtyu/P07pUQqrT0mRVavaI9ZEeFl0YcUcV9QaGbGt0mnOLttAZiJShThCG4GQ+ZidCV+InKw+M
e+SFPxUBXh8fmTM8TrnrDCEJG2xzSlgc2lvt6KFiHnys6n7vl5S1rq2qiAZNpZoIKRJtKM0gV0v0
lsuXnG8EI/esLLo7IFDxK1I1TuHHcPcLvEx7PlO+f9SmuurKQA56zrlfW+ADt45+DAmqPZbBE4OT
UELs5J75t/9wAO5IbHx/D3bSufef6zSyh6G4A8jpda0dRadKykMArhhVNKC23WQu5lcXKygIZqz/
ilznnMQe+9NPWLphmPO/iqXwBuP9SfESHI5phqrBczfkz/oS+X0+FkljRWqOkJ2O90+uNgsR3SmY
rR2NJZm7JtKDyyky1IJv2OXkf6I/gYR4vkcmHCQltHERc2msluzMvDErotRJmqiEAN8UMFYUsRf+
DuDLV7BkyVaVen3ubkhZXo8apke89L1fib3Rgpr90vWVjU93Wsrk+HpiEz0FVOCKSVBcc5dbejIq
jVngq58gulvqj4jZpwi2XBwN5cjsIjG03+R8L4Py2xa02ch/fnY89IS58aYfnzDRAk6m7UNGj2Ym
kG3Z45injfTrJlgalCkUYW5iOgR6NZgdOFKlxep2FfNa7puXJmeBSyv5WvGzLZVJ6KYvsOPaL20q
87uGG08kbGV0juwVrO8doll1NWSbS1Pk1u71Lfw1uI7NQ2ItY05afqesHJaB3fsWQu+amlbsZr/G
BNhZx/e4+8edkWLPjbIC7aPClxf11VfFd+Jk433yDEFdYeTvJLlvMJ8se8UFiRxNpMjjazO7301Q
eCkO9rSLTNzsEaD0USnu9xiQijBgOfGka8pzGcPej+Yj5EYw10yTSVlTFoLEe2y/Sm95e14IPend
vrRMtxf7p/8aNYCXiD7YHuWl5ZZL2W+9nDOVWApKuW/w0hl08qreAlxWhC5uJDREI7TOFGPcmxrE
YMo26Xj/ac/B6vSk7l11cw6rca0miPiaJ5BufKk5IyEq15eJfqYqE3NBIYOSSItBuaDyiUuh5hwt
S/zvXrkhpjcFAECWyBTXyCpLQNZ77G/Lu3NHXkl/yJv0HS6pVBloaWyNeXEejLmt1n7KYT0a0Pxy
/l0zfVMmNHEnuRwS+mZYd5rGvIkdGSKVvyqPpO3MpIOY6hCFolEX6LncIULtC1y7SRCbtQBUhDI3
LPuP/jUpaxMYJq1I9co3UQ5hysbDJbEtVJ91GSpBovbQ7kD8cF6eXzL97rZqB/TaOOIW/MXheFNX
WF96Wrle5EYs2vr3i90R/v5vhAzsUDUHOLaCXDZRlWW5dmmfxpqxyhSTmHzLV3hUA7/qi8pS/LoB
5RsX4lsCptvbhop0luJ1N0hpFEm7GCrxQh+00BWlSDH0y2q2mYz1Lo8hLnk4vXjLvFkxGmLZCgci
zffySqxBNl1769xkKObMS9lH7dWsJ/44T9nlhKW87Nd4cgECyggRIb1HF8mwrDoBwrZyrTrD5iCd
C0dykWCZ751A9iF2XwiT+lNekCdW1NcTbgcljTSazeTsnAxSY934hshchX5E95C8tl+W2drx3f9W
oRnxsmDiDoZko8IJ+wDnnYWQ43X+zQe6H11CGorNozxebvA487MOrz5ZLGqgQ7ivWv4jLDclzVWQ
cV/qt3dJ6v4J7U/liOR2icjs7W4fVcj4WxaRGSNmI+qn0P+CuNaUBprb27eBOcfv8m4wasFLo/jt
nGk3DdqkU6qmwhMklCRXu3SwfhMLXNFFIyQTfAIDH5V2YjKI89LPKC/CN8nXRyUDd+jpNB9XrYDp
I5D0hz8lLvBgolUX763qvZKU2IMT23WUVNg6j0zKFuunaYfaA6f0k//7Vm2d6SIJfFc/WR7Nn97Q
EFpSa+xYYxpDzyRgpMoVjkLXvW5AKtw89+NPz2eQ2Vx4XUnrOaHXaNFlAXfWYYzBGxtdwFDOmLOu
/2lBaL+ytPziafMIfsv9RpuzsP48/27eKPwzAeT9rXbZe2VeMAF+dCFC9xKCAv17nYPPReyfp8A8
8HtoY/eqwEj9lyraxWm7d8h40amffC+worVhFnVzgXwuSuRKbarnEaoTV85BsPZGM0BRgEWJM+hH
1iSzAjn/3UuHRQUqkh/2xUioDxdvPv5pT4IJ+sRmHMW7ew7kM0VyxSqDs/htaisb2dL9Jp/PxLmI
iEzUU9KqUGvfud7PUChZzbzXIaqC2/tzv8bwfN/trIXiLruNw1Ft/Xl6WTPto90lqJZb0j39eQZF
7kqnEUNUMYPdpgJc29TcsWlXPedKY8YcwKH/GU3IK5RRNV1c922DVfAw1AUR/TCnrme8+nuPlRna
mvj3BRhD2TNadnB3aC8nU2hdzJoCQ2YvydiekA7gJSDwpI32BYQgkqUwwxFKp7Bkuk3VwuZkj9nL
1eSNpqkr+AwYs58JAkvQoMzsGql4W56m0DBBlKlgHA1weI7OTKu2xZX1f2paluS0ubWzr2+EqxGn
u6EpOj5Uz+UhMYAShsbh6bA4t21jeUSHG7guB5L+3UTpC5+8sBCrH0pVFVkvW+icRUuoVGspz1Ft
t5hwJbLclAsqqQo8zLvzEgR3PxpcopUD7tZ2X0rrQ8/7vDowvF+ctNODiqpwmy14GWz1MBijawed
wbAbt5LblWE1KTyMHHi2manT3TIKa5LMiYPu005XDXOoSqPHP5m4rcOk886GF5O411y2GCAAMwVQ
0SmBKnScyzrjMpc3NXfH708Z4lHzGdfN87MuF972gpF0Mg4UkLkWEqrt+aG0foLz7NWEiuqVW3Jq
zAbeiEtaXbUGd+EethaDZncfk1+Ap5EA8N6Dnt6OdqNGptQtrOtl5hMDVQe/tlTZLlY+80pebDHr
ihqj+kh5e2joL/2DOSf/hdgKsLfCiDJEQwNGwctZX/1hzPz89sUKablB1wgjfkAnqkw/RAfL+vsp
pF8A6iewDtztEUGWaEvwgR87FamksjBuf6PRos7S2pBscky0yojDbJV2AY1viiZEPSZ1nKlR9kmp
D3qi0Lg4UEP+V5vu1VQkjYSBld83WKP+EfM4UE7bqd7ghEIkGgNwwPru/+eb/SJ0s29rsAovohTX
I7jsDlCRzyU81NA73Z5srsRogkHuNTEZiRqjp/4AYAFR6jBA409V9BEEW1ZaQsz/6Wip9cQtSpDN
H2mOZS/ho+4YECIZemJf0EM9YFY/F2/+dPLJicvYu9yJqXUK7Z4QHnyVXIEp6c4B4TvI5s+yDCoh
fN4xJKvDfHZPDaVBXb4kR/jNNiDqHPPM1BrmNYurXuiL71SlYWkkDLjwa/2JUr+AmNZ+e5gTK9I/
SKOH7B0MyIIFgXTGBLWitbfRv0uiTuQ/leojKuo9mqW55fNcLBIAZq4LgKTMbPLfBOWhzJuVUgCN
Y2tSud7IwujBL8Fm77A4WdB7MMItzn3afgtHu3hxJRttGUlOWZiyYpZEtzLAcx8aOE1S23uZul5K
DIVLx12s8LM8dnSrR8tc32GPezY1nf6zxR5uxB68LOjCpHWoVrOC1Xe74l4SJtZJKNcTm3x692X3
NQOzs/4hnls3GYumAN7KWIA/x6ky6jAxHdfLzzefQc58OIC2Ag6TX1xEHBRWp7TZ+b3jahV3BRyC
7tfOBO0dGsDKRvQEbHDo80FN7SmCNk/DFl91iPZaF7v8Y9qWCjbZ5NhSCqocDHe6W6e/L3NXUWcF
gVK1ibq6Gxfbtey4i1eSWJgjU3FtnGx478qf/3fCRP3A9zOul90E2HyCTSTU9T2e/S9OSbEhqV11
gJbXH0791IWNkKABx7hvdQw5SsyZTWVs0X52NHFKGRlzS0v60gNzh6BeBJfxAzC2b9Ex15gaTEeM
41i00KZRks2ubIkfiCvoiB3xQHzLKsfJ1yHndKK0sgJ64cdTYlOPZYjTR10V9eSRARbCjC28rrFp
jywF+TzT3w6RwTNyxM8JkqJHpQMMq1+pVk68chSJ3ZNDCQmZXX6k2s3Nx+sjbjasOBX07I1MS78q
Ex+WNSkLCeLvNJ7aFkpZ5r4V3zvBIJUgtEq+4A/C7eqUp7oEy9gzwrb6r4M5tezReiQyErYGBMAC
Ok7PWQ0ZS/fFWObnSHxjtGqjbSp2P51EI7b9E1ShDULQw4ZGVIoGGZc24QYveFmlTGUmzKXpAyNh
fMB1QcMFk9A+YJaKYlByLoyKpZ1MLwq1H3/Cl60qyhg/QZsYcTK3U3lY4+YsUGLBP8FCCsij8S5B
TiCqExQR5TwfcTCQLE2O2gXbRhwmLUywOEUtzN+tqoAD1PRtK/Zno6JQ5mVzb3abZKPGQquTulua
8OljkQp0nd39ZaMo6HSHuNLKKWwEzPJ30iksrR89EL69BsNJIucCYWpc9Bc0aBSBmsZ0aKKhfYJH
4CnEexIMQyuk/9Y53hdIbkcIUSilEhtSdIuG7mgDHB2SRFI7uCuNlA+wKKvVxXwlhvt2F0MY9RSC
rVbSTEmuhrpPl7T7Kiyh8ByqKNjK0zMhUfJ23nL34CdSAmedgmIfZh3jazciGYZNxSXfCDBTQeFF
SiqB3o5PE72/kPW4HRJZi1TQQhLzFq0IFprSyFsXw31RjZKTkz9KHR+P2D/AJkg4cG6GfygkqD8s
JCbBhRQ1RFyRAqF7+/XAV/gjR/pGGEhQZXipYloOVnSxszbhQmhSwVKbWiEBsioZ+daGu5CEHjPb
FAEbvtdeDVUsLRnO667cwuHVrHbc0ZuYGS67dAUse+zrDBkKA5UrMksaj/EcD+HKkMdYHPtuvy2N
9zoL5Z+gdUYeCD/bu1TL9cLZTbXQiXv1KSPsz+bfeQau1k9/kY8YZehXie6fpuDAoOrpDLW8eUew
rN/whKpZNeUP+AQF9cppDEWzofxqLq28zuihDdHC2Y8qj2GEQQiy2dosrb6K7a4k3aQ0nnVQGhVk
l09ZyDNkvUG2C/MPVr2VoVEmNKaDKyqcvZKwJsdYjAAc1qVtSOLHNxIR9qKXAVRVlznYMLuA9/dz
2Dr4bPFPzcK6HhFiGzBBzzK2jAVNh9EH0PTMSf40qtaxUbwxduv8tOZ9vDHU3tYXYymg8XNNZA4f
Nljzn8ilO64weQTvaDeiKgZHkTsJThRpVY++y1TA7T1cOsGnxKPBeE4dhLK+eAz4hdQYNR8Ydl9J
p0mQogw40IP+jgbvfuP4ao6FSwV1vc9OmNHep80UaZ8GEWsR/2thUVnSZOwRmjBy3wksaq46kCYP
X5Ouf9qqSz63uIxjYV6HLuhcdpzIqFBpy4lnqlworhshOvx8dd9lpDmcpgAP3hmQYU/d8rVJMPMv
bFBmtTAq08+Kcx5KXwGz7L+sEeBaeYr6mSGZqVoUd8sb9wBtttsydrFZn0HGJ86dNG9X8BuURZDL
Fi1kazpnZuGCh+88Q0eI7xnwuqWFPn1sw+AMKYkq3pH/J4etisORQYHq3C2+aWh/PqXs6cZ5Jh14
1wAXl+1/3kk8uTQpEx8dhTbb6N9tewdETpARhSfdsrVm/hlepv4OHGL0rNs3PxUUKsKMLMrSXFwp
9B+r3vpAN+NBXd9IqPcNv2zqelEBHjbgeEsPbT9OHqR/Q3by8y5vOIAsJR0bWHy7NIFTr4XeLM+R
gSURrVxUxdngakmXK/ZC9jS3bymFMy7Mx0KQc7NRWv2ZBN9bT7oFqPF21Egh7v1y/Vh6ciM3vAtS
oqLS7d9Ke8PBxC9aZkceYoa+KgUcqGt1XUAsOUYAygO2vKIHPAt9WtVvmvjwDx5XUtTunGyD1PBR
QTd4cnAlpGYM1AptJguPgolNc4VcA+iYe/HLeumU0bPWhn+mDXVIVA+6j7rSw1PbeSD/xIGEgcCj
qrr7aDZUsegUnDhWEgTo3+I/l0sEGfxCzO1ZsosguwuesiC4i2kWlw283nRHOE7ikQyfnFxdqBfn
DeOIjqSYqCvdVf3wAD3T7nQNaF5i8OXcVrzlw6LnFxPvRsV63k6zXZoawCeIrCWPtlFgSdR4r7mz
HTUg9jNUhbcIwRhZ4XdBPVKDbRVzBkMM6CDF6YUkQrjlGsEPQM6V+l0gE4kGuiDkABvur9FhzZJ1
DIAb94ji+FS1jWfF1RBVzmUmAw9fNJz/JeZLPMTfhPYs/o25XJJhj/PwiMx2JGPYrbj5j/yOSesR
rsz5O7WwJo4pLSK1blm0y8K3uj3uK6K9N3+0sHt3kJRnr7dH414KGoKPXCDhcF0QRs5aEhyoUp3Q
EBVEFD6ufyZ9AN0nvaqj17QOA2ccM0l6BDPSfKXZ0DqY9riy5hrw5l+enjxEgGN1myxnXo6blGYv
WiivFWmnPDdp43lPX9HCKhwNmfCT4Cq4pij2woIeRPWFuEde9vjeZJYeAQnpVQdWTb7h+gRmCgLu
mM8pAaNfpvvWyF6wdDxmSPMynADji3Zcy50up1YZMuNYvgs//Whbw+qPnTCkNSefbwKfgxjBFuWw
4diq6RScGy7nwPYeaeRZpQPBodS+Y++xG0CvqdtpjS6wO7IzM426Ig7OTydEDP4pLj0hwxuAu9FN
KZ6cLwBvKMGZGEQKdzVTkzR26Xk4PLjGaSMb6Cab+uVmF42xor8pVDyNJqKpYStO/gpFsD2N5DsZ
qm0epdpOXAKxv3+izJaJvWRmLJkrB6famWzxw6ZlcKdBW/X+0TpB9wE//owTywFo5Z6C+yq1rMLM
edJe4FV6drtA5MXidsPnRxYPgcbeDmWTNHHUIwquBl6W0mopg22y5+XuKIEDdjIMiOWctArVWLs6
KGAioFNbdq+2KR3rkZ3DoziYFXmlEPiThhBX4buXSl7kQdotcZT4/Ax9IGlzP+seGdCyn2EctqEs
3vdZadUh40B7yVEYyW/UOjvnqBduenWnWad44QSbc1mrI201wESJSJzdpOtDCfE2iPoNUX378Sm+
dFUy6H7X0Pu8JoMbW8EInEHwPB2OEmtLiBwC1UoZVtIJW890e0w1jfP67YpFLIXNZBpfPocCU8r2
LxIXthyqYsdpygibDLzxb3K6Dd1w8dWqXR6bAksiuzu7b/c3ZfnekRBh2xPQo966EIZkOBSDnD/D
qAocusvFTrRUq8C2ZC2/O0tDizjzrjeOPQsSant02XHhxMo4tIJt18ZwjiA42TNa9plwQvhvsmzr
Y8msuCvrd/iHdLzlTxW35xhWUzLfurIeC+dffR6edMJM0vPrMRW2kHLcKQAbmxtCAk6jip0SPF1f
2Qky6liO9kZHmryB9KdLysDjT70ADPghjLEXmhHhhk2rMWh9hRIMCUVFuHytc7DP8gbGAkVHi7sI
6zDeHp4Pswo2o4XD3fuMb5fAnHChnOSRm5PhbKSH9KaJ2hQkQ+fmpNA20zUHH2GOWSrSlKuYSRRt
ylWBXlZaKutc2xCRK5+MJO/dRAYWDnZvh22LAaEmvE/9tTL0kK9YKReJrCDQH0q0LXdx7k0IzDIY
/vxb0RBo3C3z0sV0s0C4qMN6ngPMkDFw+SHKah0q/xzox1PRVmYmNYbzGzfJjY4NQMELEvBVt73h
YYcVZPGeJlnM793bX4hDNV7Ob6nKNjJgn6ME5v63nnWESfw8fe7YKdAi8t0dZHi2p809Kfxxuh8s
xFdyiO4X57j9DJTrckl/ha21+7u397P0RMB6a8KajUkjageeSoVDly/SE05LnwgG+ULpPf8Jf+vF
Lj/QER8kjGgrX0TqfHVsoaSXJoI8oMApPHXuGtXYR4nJOemXl79NMf+brbBHF8aHV6SopOipPjcM
cal1unLVuv9hqtEBCsoGX3HICqa82EGLk5yVF4paM8eOwGHkB2uSdGQrTVia8gD1bEim8slwvvC5
reNVtX3HrpzdOdlyniT5/DH+3ej51dbl7iWr+IlHuVanjjU52rc3pxPUwdA5iSwKihpc4O83Mz6u
Q6hp7lqSBtAPGz7wWRBfujAbLeRB7uEF6QRAxME2mNsSFh74GNAio8Tp2fjtEy9UeVaLgMeFocdZ
PrchrCrQp2XhG8B8VceOrV6zzLvmvrbxOZy1OfV/lffJRiO+lOMjJr2GsqudbXm46dT7c9gZNHOU
sVY76vmynOL5LUJum8vbZuQYLnj/XWmoGFYO80cifuup6tLSKADsTliVQezEjVFYjsRWGzh0aFaQ
/K/jx54LulbuPK034r/PzBxibQ2haXJQyBK2JXMZXLCGYknMb7nARfRwx/J/hsUZ54E7d+4jtuJr
Ig8ewIHHfOFBWRzFrsoXJCNq57GYt8jpsV4QVUTciHtpVCG9m2bJ0FPrO5TaC83aHnSFq/co2t8Q
WeMuknXND63YAV2Kv7NQLhfagVmnNxZl+YIskErILVyfegUlqiD/IejdrWqhRwtTaRxElPxMl55J
YWXHJILIT8cOmEki4s3uHxI9NOgEAKVBIkO+FIRe3HgmXwPFRYyPwE1SeaPcgvFnh02nMPeAn004
9wkL4kXANAxuBk5BlbSUy3FuTFbFISOeilJ1XtJx1Q5B/aoOaboblp79YZTvgD8t4z0JarLVK6ca
lcK6XgXtDNM1kr0yrXzOoLQh/dSSuW9gqOJ9N5HxpVRrh+KCfBF2Dfb8eMnmpp6/gO01ChmA4LU5
ABfZP6DaZ9a9/Lwg8PYMBn0YvCAU9JfaPCDj7O3q3T9ZTpYg/XMf7rgPTOc2ZgwmR9LVJDczVYuO
0igLMZGcm3FbQfunPZhWLf65ABp5yRX52uSOva6XwK6Mz1RKUwMS90QT1py0HAN2vx0bn4D2eHzS
hiw4tjOiN5gexkb0kICKCcru8fPy08H8ikt+5digHsV6srqbDWcb+jmVqj3AkhQ38gRMO5RoEp95
lMfnc94KxZrx8gphNYrXZKHusedRdm77GEA7oTnTjLmOsVfwvHKJvLERayCFkdeA6IIW9/Poiaeb
xtSOtKH4iR3dFUp/rputSAjaJV87HKV8gT0P0bgSczGf9EZK9V+HE9UmEHnZCAGoJtshF+8t9drt
Z9jPCljKIoBJFo56sHjofZw6f00/mCWgmUo1AmNzPtiGQuCxjyVUf8D3eu0GxuZ6HdlEnSPVEdcP
edB04dIVvEIVe3i8cD90Nns7bLU2y+M0a+liU/wcxpgJe5ZtbW07RNx4VSfH6yoglxKyjcas9aNX
1AIP47sQB34KXB1EFSX/LBe/d3fGc19jo4QsFYlotVhCqHoNAZ+vBSQMqnp0b/2KYM7K9SqqsMTX
reTQZ1ZTnq0YppS2AfHtiwmJEnzvqRB2l3JQNhzrOijQqRvUNdTzrKDwxgw5uU4luqZrXgAYZk28
iZdU5lJkSDTfYmI8+rZrk8BB/w5ThY7PXvuillDIFS+on1w8aki2Zq/YYRi2hu0TQKOU4GjyQZWT
G8IA8vJFG0rvclIDbnj8zRY5+XwxXX0FL9mhS+J1UwrKu9/hqYajDuQL22rXiCHGBR66/j7rQpCq
/6EuUuf/o8W/p3YPbEQjVSK/mIcJ4oahWJjIOzURmY0ypsdFcSt2hcBm8AImQn1BLfN7nfLbekD+
xUVaPHWKBRcg5Glmp3kR13QU6ofhRexLx6ayj5nNni9/j9cO5lgC4f4/a1YHBhJelyX1VU7Q02b9
CryqJTrUEZTabKTWDuTcwH4uI28cgAwTM2k/SNjZjSuUASHlAhCrPF96yacy71fntcEsBOuTqdjN
18O1VQmLGOCT8M9i9PV8EYLGFNlcLurrXSHbB+yDocH5h7bUj9inSuJ/wYOmziiqI2TNqSWAPH5s
Du+EGTB76guMJ9zNGS9beLXW9OIgdfgchGluxsWV2dNKjmhaQsi4Ae15jPG0Y89zPwojUDizBNc1
M5p8ooSyY5cP1lzcyFbxciIMVms3AdVC8/aLSJqoqWZSddILgt6L7WHBmRzLA83kTqIyUtglfWBd
nJD7fhWejn24ROScH+IW57GGluOwEUFzzFjwiRfHg5cUunvKe3Rn8JPS0RtVCiGodihtmNQsXVke
Z+VVjxCPBtWZ0sMCVL8a08g5cK16kujsCJeV6Mloj+igIBuo4OIYUNoACncgDb6pm9jmAnzf5OBd
bqSTZ8iWbuGQ0GUW6TlbwrxsXs+5AtAHiFQ0HGq3AJvQvXnJWqVcq/B/o2EfG8mEu/jTmkJYfyiU
x+joqkLF+i0dYnEWhmvj207N9tXQCHemzPQIKOExk+u03adA06OylBkXMv17eGQ+7pX+2X6mzolw
tS5H/5q/boP1HzFs4zuInU3Ls68Q0IPEh8pJ6d7b1nczLx5todb5L0WUm8SIGQfd6Q6GBQGQOUB6
3+19w+UlPmzvqqDICV0DdRSerL+mKhdNveiNR7LLMOXSJyblJYp4yXJa7rioUw59tE2tk25lTRws
IX+6y0s7bVFz7qcigXcwWtQh7tXfY45nLrF04N50e9Q9G1GYAxIbhCDKHHVEz4vLVrwGLqzo4+Mn
wSKfM0ZehsCZ+hln4QM7AiKs7VPnl9uLIU3vJc8Zzgvxmtx9OEfsvIPPrf9/ra5hKRHMSDn2D+T8
QgbzdRRMDkYILuQU6tiZzA8kb1vUvrh0V+k9Tx8dsYRlbfO9s1Re7Dlkw8T1s6EPWO42smD1Pc74
mtguQf62Cc/KLZfwyqJSui8Pz81p50wLPxHdnwid8Um0xYkxHqdR2aHINdUI70F3byv/tzzshhTK
JXgC5N50JUSoE9K7ZwdpEFKQAZo+BfFUujGK3wtBP0dvvSMvqirta8AfjyaLXQr4zVzj+NtgQjs0
hAZ7N+0E+7QTt9s07vaqWfawVEJP/6pZ4DElSaMuGmLUS6amcT8BnTXLmzztws28H9qEznKK5+ef
glXqMJHU+jxI89dj42WUOZEGLosvAPEjgvgO4D71wL9bmEsJPCKkdug1J7UJdN9ot1VdAqAoScoK
gKVtGk02n86Ug+8o/GN92UvQlfTfEf1BX+skCYy7QVfye312DAoDNZ3xRzD20IIVxXmjkx8h5BhS
dftLgq52sTg3IVqo6qps93hKdq9zU0uLrRWbTkfiP4fRXpE0zUncrdF0RLAMwGXjJpEbgm4bWCv1
1bA/uOSIaEeURZKbt3u366/FKZzonCTw8OpI/VyFbP5252U5uKlxKxdS2uqxvFfWR0jQnbJCDedF
hMHAFQUn5ITDWybM6O0YpwxHEvQuOevr+jyIuz8hJBV6hgIm7lgq/jiU4x2mNVpGar4Thde+NQac
v4Z9rW0RcC+VbZxoV7HZYGpeA0e1VAUl8RQ63IpUtTkz2KhqcFhiedFmJtedrjvP3CDQTkC7yu31
m/264J2lFdUCExwvvmSKzY45kGsmym08iTPVY6E69HXcZANn3j6ZgbeFD0Kn1GMZkrVhPfNgH4dA
BKOZG4FtW8JgI9uB2t1Fno9jL4DK4ElLsL1TOTNHISs88QZ6YmEFr4jLJ49LVAK51VcKW21/uxKv
qEf3i99Lm7d0swPEbQAWt1qRhgWwmmI633bEbtllY0tTADD0dz8DCxAY8cZaNpsM5if6+XTHhAcj
IzHkpd2e/Z1DrBpXA3i/9xzH1r+0Fwyj/YM7uf7blLHrhZtQ2K13iU5mDIpCiBPBdFUgfIpqP8d0
R+pYhmLLS27e14UvvYiwhY0qm3IdKQYjmGu8ZGysyJh74AMRkLDrAgDDhjd+Ae0CHd8VdVxSNTVy
/H2vgeBNV+XC1EsvFcelf67JlF/TotL0+HlBb3HYYz9fwp+jUMlsTqjDk7ebNkmsQSURgnkN5bOU
2RkpvfDFhE4dArZFv/OJtNhaDvshmn6zPNZDoYJU7zWpNjAXBu1aG0a7THNK6XgNaiyufrbCn0uB
3jJcB5K3SvFhcCjNzRNZG/C9rksseIDSl4RkIxFrH0NoXd/bp0WQDF7bmpvVa7A1ZaJJIRJTLIf6
Ij1b332UqNRgA984vA7Mr3AxPFgrg0zV8qeoNC4NsyiabndXSoFyQcpYiC5btqTSqK67KAfEp5be
kdBQEnoOVX0cplNTE0QsUDEESlIPtBChIPQ/vIcNhMTBNbU7n1OSDL64xhRIoDx+R8DJwtF2O2Rm
liDtEXnSWT/n2gXnZSmKSxYnw6TW3qewSdXkVXYiGG5a6nNyEcujdYZ+VyZCqVVXW/miAI8rxYm7
CKdXQR2bugXBdQg8Xb95S7HduNenx6FpP8usxjo8mjDrev3AiQOkh5Xd6cDjflsFyyQgvTynEKuB
ayOzs/a6qz3i+eaRSx8Nrcat8un0o/TIKd82GaDZPBqjml6Uym94JJL6B98Xvb3fjDcDoU4BJhhM
IFXsGesCLGJCVWt7YcScTRRHO2EsDO04VaSQ1rzKgkUWbYaI7593qvIqHpRVTe4qTBpt2P7t0Y7f
0U2/Vs7NhAAuvzhw+2mBcHEW/7mRKK75WYf/8cKivltlfzwvJxStgGRyZ9T5y/edYoUxCFNAyo6l
G4Ekv//ipJqGFCFRpb0j9oK4gTFO3zrBpQT0QAoCoN5xsQgYPFEDlpjhcFQpmy/a/TaXA2eUlKYl
MyDP5H0Q068EVEpoWpYJGibFwnyDvVsFGu7/YRdzw+pIboJ4FFLKKfDrWFpD5ektEWkFa5X+Ykt+
ZyaigLRmgajSwcyUNx75n5NyPBtW8/yDKMw+K+URFdu/ubTIsJ9Tc60bV1h8XlOanbCGKVyBfY7C
7rnUXpmlUt7UNRfcidV08OZCkm5XO0PkGXsOUk7HRE/SQlTmtxv1lctGBaCQLTaRPAoSV3TSkUZr
6lCFx09h3Am9Pb6deN9cGmx3IGml21viLmxEN24NNCGZlEmBV5rjCfrHTrlsgHkTD6bO1gIm/jZw
zqzR6BxyDPafVdpnMXmVPVTeUq9cFpOXtoLw4DqAy2XFZCDSFxty01X0W8PqyeNGj4F8rgDyTgEm
x6tWqzTXTJttfohjCb4K/h5BFwsg4oMw5xnsBZzkygajFNfZY4jHo7bzrMr8vcjGU8kJrVUDBLTf
p2+anoje5v6xteDbB/6xKzA5cUBbmJz6i0ZhYAqrfa7I2e0SDgaVWCYaMwpQWkoBfXfpY0rz8iE1
rclG8LnUgPz+SefuJJRaolIiyRo7zdsZQ4lmAPhz2nhbG/BQ5H/fRTXjW/baNYGl/GXn71j8nVcr
30lYiYHrUcBZr7GMkwwSiio6iEV6gw7H3soDzvlh3tTB6RU6peWu56B8LTFeEsOBv+oNLIYGBuNJ
R2s0MBKtQHDDBZGnsPIW1Al63qqA2EXl9aEmlh82URe5S54D9+0HBI7h6CnGuMBCuDxWJi6ymZb4
70qxW1cBY2tL8uhSJAA4QixZf+KHN0xDb7JLL8ShT2FOVEKegJiKiHZRSHRY0nLUGbji3b3E41P8
Ul+7fLvYZd08aCoAoU0MsTMELkgG/Bo9ostT1S0mVeX6rgewfOQT9kC3N1Iwul3DbdrhCbHiSyE7
9bmxrr+5BygJ9bcWZkWQJcnZMvs+FE34j2Mpq4cGJgJ6nQ9OmqcE4YiTfzlw7rzMmowTTFmEMt2C
2u35SCOFVmNHNbIOTSTUZ4DG8VDVOXoEFKuizIrGO399zD4q0g/Q5iDda1haUe7PfSZXpZdwXxyI
BSNSASa+HnecA4L3PQBs2QfhgFWAY9IYf1tSHZQEeuvbk9hbFhQzF68dN36gdowtf2qgr+R1/y+P
Lah6jSQlsr2gPkoSZsT+Q8gWqaRHCS4fBopPJ90FHt+NzhEcSUqjMmVQTk+wPwuCMUmL2xTOAnhE
fOOCSAkQ+5v/UDQuTUBRO0yVbsveY4txVQuTkUQX/b1WfCn1vwI1u+uGdyUHliTEgwHJh220hP9x
pWWlwiUiJ477a4+8gekxYWsVLDYULadSLvzeMLh8+fDS3HHi5ygLbfq00Jes5+EEoj8NJS7Ltp3b
khXQ+VHn4h0VDJe1KF5uqdVowi0gqQzZgp4y2bYkKvNgT+vLs/O1dNyRzaGWHxh6TD5cOzznl6Bs
8CaEj8NGlKnupmghwi5seDXcwAOul30o5NmUUuT/iKqkluSJcg17BN9bf9/54AfWIfLpf2/smcQ2
ILLbSsVz5HcHKHq9c1tPHXNnCFzExA+Gg34cJhk8tMF0F5865LKMeIMsPqn4ljc3u23Pau5w0IBV
saqfV3uYucSvwlDni3qThrqorWFHOvSZ9YSrjhR9OJs8HtmusCoknzM1VSNayPm4uGgnpfktiqsk
DQOhrMYnHSVcB3WRWz1DlhSYjPlQTkLGgeG3KNyDTgkuejgJJER7s0gjMmCQVsoxxZhSOiMdACjk
WBnMyiXv/mWWKLwZFEqeMuD986e4Mrbmv5aHUeJ6AGtFlu6SGW6/aC4tL8IwM3EjmbeE9qAJ74+O
xPlW3qFxctegnw7p6LFuop+IABQg0ViCuNIHbq4UcJAJRppFfaXSAKcPVq+EtvuqmxqlvvA0UgkT
6/vRss6NpU1IojALsVNKF+z0eiLjwTywC02PVZsO/wXZFZqYkcgU2PB/tNBgUPu7ClmOItfA+ChE
wp4CAnS2wAp68UFEYZRZ70R4raKC4my2f9vL+GHSi5yLiW0TDSDNOXdiks8pwCo50u8ZPLB8AyZz
RzoLN0f1YLEi4N7ZunLfmSc29UKp+9m3zrea3XAcRUVztGRUQEl2G2KT7krUGyMZaIF3S5/e2cuc
CVHRrfyWh0H1RXVydFiKQsfLdHy7dFxZDqJzmVVFU4/+fwlpUlX7myrSSoP3oHgPovgcEcKemlMa
sxlEfn00Xw9TjXMShbIgXNld/R2ftzfvLHBRzoaP9zPJH7iL7TsiAVtVB2uoz9TY7c+lM0Bwp2wQ
/5QjPicg/ODB8nD12MbeZYvyTsw1mI7vxgB6qtp+d9HewxBsiAm64t1p3cTdQsOK87/sIW5j6RqQ
rjiPhdqebxk02yH9b0T+4IMkC3gjiJ/elxqa429Mo6xjV7Vq4aFSIzOPo9AAfTbzUdCPEmCcGu2X
yDJiLH7CbmE066XhQRBIgoi0Z4WPW1r5WNT8ZmXenBolrqQ3F2y9osbQbpr+18YsNZWQjZCT8Hkq
Zo5I8KVLMrNU9qMBHzR36tK7kUw52NZkX633GbwtXg/H1oXSjNbrUUs83hu/hFdILu4TLUsSCIc7
6bAugEVGaInH+fKqcURnklgRKnRCVIQK6nuiT1BSzU10xK4uke2WODSj646kMxFQTgUKMbEwNGCX
K2a8J8Xhn+9aZXsQ+qgYTTyvVQlFvqM1HLz9dDhk3bkVmsV+NRF6Oh9WRmJCoa22MXfTBO5qn641
84/Mfy9W7P0RzwUuVd3gZ1fJ9yOnYwCPwpwfUSWdNPT7dg2nQjm5V6m2jneROWmc0+KNR+9j4cO3
ifCEDZet1ntxGTQ2Bq+EtlEiCLLBdtxf0n0fCduu09iT2bKWJXvpYZRwv87E0scay7jzVe0+QPeo
xSZqM9tsnUpUMDJMCchlmNMOgviYVlPFZWfs3bnYtNG6pkNZKd1Wyo9wt1F8CA3xRWJaXF8rgZX8
/KBl7qXOtNSa9gPit024URfW6QZ/p61+wyEEflOEW239BZwFM6QeLpCl+4DvgJNkH+cq2zPbNYoz
9TGptvWHGZdud8dNUX3mMtxGcOBzHes5Wi6AD0QMlI8sIyROCAPL8QAYYXoTCSZFgdB/V5zVzulN
qiGuhxgIUaqxWbq0vtZjWd22fr+rzNNTw07fGOf07K+LBZGEAhIgOtD/JJNqYcpWEJ7VLgW9oFYS
UuF0GAuIGlotT1Y653nbe7CvpVUYUkohBX4BdHcXJz3FUv6QmSYFZ6EsjkjWUMYcwPukvAbcpJoS
hKgfsDHbScg9AlbVUv46dt/A0xb1nCWHY50sj6H3oaDwYebeZxFGO3taJs1Z0BHCUXJu8GD7lf+q
ZzKAZ+IMKY311KzylpNBOxAV0U7teiiJ6U2IQxYvPmXTJvXClKKSl6LfYrGHl7qiHI82anyBdxhR
jqTOdDplFEALw9EnWFquAA0l04xH2vZIhpqW2MxH52r7k8U79OyZ1EirmtR9ffoMaTVohTAjRmdu
XVZNT13l3WkF5xIn9hoQrDJxslqvI6U6QTozvLdQq3tkGmJ4f6GLVs6IkHS9/Ckc2nrFLzNO31os
uc6BTZF3dgUpIH5vnXsHLrJKM1Jo75y9ZX/q4dn17mei3r11PjiHEKW2JK17WKOHcEn4LH9AJEoz
yKOOBk/ZYaW0xRvaTpmQm95IrRGmMJ4/RV/e03O0d03qsT27AXDtDbGx92ITdNxYWpGOV6kCuTUG
PgzjqTZlal76mi1iRdrNoQz3kRx8L4OJuM0FDwj8RKmNSRAONMaJuvHvbzCfJhZiCnBgtvkOz8V6
gZ1X0TRqe7RjTAIifJa38XSbRiDJ+S10F8FdX6SqQRuXvh1lx3BPU1mfx3DxoqGP67mTooNsy+y0
f+H8kM0FYC8CHnbUEWoHjuhqUFIIwq41LlAGAhsiI1hHiB1NglVsGl5kz7qg6bEcOBhsIiEd+c9X
xPc5/Q95HxcLXO4M7/HYjRg7V4ELabQAckOsb6KCdAzMPdxYYvJOwjBp5QQ6d78ZlbuTUp4nYHjd
XRs0q11zjZHt1F6jy/jaZoKdMxowCeLYdAxhkU4G4UYC0ZumY3prRip8dTubXOQ+a0FXe73KKAme
YimRDOAMZvLn6fgPS5os2lJQDou2Jzg5peEXc2/mfUMBm9w8GSpLtBv41jI1tixFxlxer/r7IoVd
tOxigOjnH4wO8SXzW/DggdB3Dn+yJpb1td0VUWMLajaKznjXC2y9ny4RfaAtMLrdBNsbjxOvTeQ/
bcqbpk3HBaqXmSCaQlfYpRmlGJQyeuK1gpT/DgvWSxNheA01evdbYMm4ZO04XxCB8VDhDQDjYhPr
ZM6Pk8Trl0aHD5ZEXnwwcW7cEh5TTIjegY3VvhToBafMiM1rPJzAzcBtTG/wNyXdrmpEOj1psnVe
93KMFOW3iJeBsCUT0QHFiJnsFy0XOCI55epRArVHm6x1vYpVScTlwbC8ohzh8hfJ+/ilWxd610B3
PMYn26V1Js0oN0eTFQCM3UFT3FeIrp5qCLRCKzscG71ou7OA8TOVrujnveHlaBJxoUFvHrFZFkYt
q/jyAnZqd/0QpLa/ucC1/Gi0e/nS4UFppdLm0ie2y4Hr4qf2QvhtPVaa9joEPnzin1d2WfBFa34M
8ExhFlxVLu3VMJ9562junUtY9HAC102GIrABHgA0vgGBBE0nszDw+Y8ygYPJTLhadd64WvcKHXGh
xPH0EEnn06MtIW0NazpQLm5+ZRisyHudV/rGOvNLX9paa8H8+oQC+eP+PT6Klq1OztLNfB8OWETv
C0PeJ+9Yev2iMTb3sXplBWkf/kA5jbfcVLE4TOiKAcRaG8ImOjLQEOdAgva7hEII7am+yjp7NcS7
ispUz27cfF+e9QHiBhsObbTVJV6pjZWogeij+2yvrRMWMVFY7gU9Ep9+sWXl3ZlEBidfeW6wFDih
s+4HcMAZigHXjoc1D7lqE0TTWH1+zUF1k7iAwLGDswnlZ9I35B4O9VM8UbIKj3Z7nC8Er2P2zDgT
4+9FjC9GPNGKAT4RdZdNMJhJ9TYlakLiNttGM4jx1/xy1X2WZ88n+MguPmRTDIQKAnAcuvPpKW/4
JM2dSyGmhCRjAoCFzeTZ+B5o12sk/UlYnMaTpEufLjQ8dq4853TwexwaLqO2+CCMbaansQV5Ziu1
EYS153/C4ZhfPmFg06xn+Bf/9pmzUKA6/j75tsqAQnq5Q7NBA6bUlQla43J4vlRqDqA9Z21S3fOh
NqbX6vYGPiYEFe5M66VfUw2f52DBOnIBNyTrfc2O238OhTmH6bxXgbAo730liCgpc9jbsRM6Efx+
ssm1UblCTC1wpjKRriItPHrLRo9owblx8LS6eVgJF10tyhgdC8fwm75kzsaAFyTqLXKhzC/URjpc
so4jE3a0saDlX/Ov6bR8LzBMe0W7awkdSoQhQib1fO5JrJVB5IjMtJKT7DPXdXe8cZluC6LWkCsG
0ZYhbxhiRTB1+Jpa/X/aUGlU+iStsTR/Io3MuCs0fI3zZga8pex8m6VQ9MHx4kF4SfX63rk0Uf0o
24ZFDpjv+kptcfjTfnPjRNTUmI9l6haPUDEC8c6sGNf39SKWSr9FvT/9vwgvMhm2fB3M3DeGvMeP
9JcDStu6xJd2Ho0LwJ/96UW3DYUnWzJH8fMylthodIxTp/U07uwnQq/PE9kWTyZ6a4qXV91ozEW4
YVIipS6bKA37GCry8c+Z4coaywUXelystWMpfCBYhRYIneVSseM1NVJScsXNcYmP35IyLIB7UuVy
ATOjHdfbWjq2Tkqs06BbB1uuqtpYuuLFQwXvbPLKd8r8LxjcN0OQBLnDnWe36zCVnuQd94uAiJvy
YGDFVhnktwwcdbLLBpG6YWmCgG9kt96h2Onolr3FLiYFxgJX2ClqeCS2gcu4nd6KRZBFhclEE0Sj
jSeMfXQ15v+Obqs2DG/x/Zy+buCzSmd0J9oypzyjeV4IuGnBOiWdu77yLj6wC3oop2dKFpPHgLew
7OktypHqzIY49i0uEF9gS6/ThLLdmWSwh51gIbezNtW/KckZEH39nIyNocT8Tg1ti4Gnx2ob4Cx5
0rkIOk/N2xqpDi+YzZhwGxelGzshWbcd2bl2MSPyBEPGxFLXoy0IgvwGp2cmFpKM543StyehR5FP
BR0BPScfrUGKxFn+oDl/wS2xB75DStHir4otDQKv72yRdh6KNGoIdrV8izM5WHJUiVM+EJgFyQ8q
F8hZJDHTH6EJQRWgvtocMOuToM0VlMrBajDGHN1FYTqn4havMW8bTMOlPtnLDijUsX6BF3Icdbkh
KeyXvW2dC/+OL0ZyVWV3mwPZwm1UluNR5KdxhD/WG0vvPXzoxK89u/PGZbzD4QtR5ChEVGSLSlYm
6Ay2NZwAR6uwUB/ZeWkioHkHzsXszZlUUJK8bkfyyeOKePsCSVKWXNVPViutkPbcBIkTotgc2uTs
tpdIkwxrL4xE/V89J0ux8g6z9xG/97ExH6gakZCsoDPHm0jHhbkv4edp3SXuGEc18cw1wHihgQxC
+fnSgJOoWMtODPEkhq+7YNg2J1WFObS0tjOVJ4VWQyhaKfXMD9F9V2Ee9G5WQKhIuLe61ylEOccl
xS20LW5Adbx7VjhQj5tLQuyJQWvmdUnHVHHJbTGnGeN7E4ybhx/jgkIta03JyCMz7v5SWyMhgWBn
LmDNnHzhr5Q08u1ycK3FRO5lzwnOOajNCKxKpQUaf+f3qDQ77u6paQc56GMwNm0xdEsVhBApPVIA
4XvsCa8aA0W9QBAF4F2/JxxmW99W6qU4z01NpKgrqDFoERgoRckjNWt7SCoWXrPaUAFfst/BlQhr
bIBPWV+Qqc3KDmRYAyTlIizUkUiiSus7jZTHyL9dtjhRMHYufcnuAu1RPP/GjIqJHPexKSRRVpMI
kVLm8NVy49D2ZjcoWELuRlNwQGPcWFSLn1waiRKbhbtStBVPOlxNxerSSo1foZkPelfxEVeArgqw
RzoF8BPtp+1FkpK0lOplGa/3Dotp14f2kCWYxdRudYTZj00RRj4xs29iIcunTvPPSuuqgyjPA6k2
Z48u84dL01IrhbY9Lngt3la9MVLFMmPnWTYQIzKgn8H1obOo8Pfd8+svetx5KpE769F/vagNo88x
LVXCQwwr+Cb00xKCOakA0mGphdMx8vYIhw0HajRsTgSdYQqQFTzX+f3hpPpyCXOC3vNQeIQp+hne
f8rjyMk4AHUwBp0rszUQhws/IwckYdUUweQ5xLvIVEzOUWa/3XamV1pXsLyugALezgWxBL3ga6t4
/428id/0xTabtqKvOaE725zvxQ4B+MFQdSI1dW5lLM5Dm+1yy2Pt4eiT+gEoYGD6cFdNPKmoIZB4
+cbsuyImisn/saZFV3JneyX5KmT520WdYVE98INcqFjPRe06gspdw8cEM2exZsRVgm2OT6+St9oN
zqxtwilQYHeoohfGORe4RpkrT526ttpedLd43IbNhmzdJ+vqAjiRq8WOUAhX8B41OOEpZ6vOI+o9
3E/5DgfNnlsp8GnQeMdMuGG+oVxmjcXiG72MK/ARg9I0K2yJ3HN2D5dph7Ne/YePPeFNiUShjbho
x+GhnLP2Y2vb/E1SQUlaDrDpnJcwkDhfQDY2w5Ewm9EmALdVxpgOr2bLeB9AC6SmUwu0OP/dl/8Y
iL5CMTOmIAIFKtDvVeFqQLyr599di72fZnt5PYjUvJ3K1oWJ17Pp0HcwlLuYiZ3/pN0SUoYY+wrS
wd4jYP3Z7lggYi+nM6+kkXI4Jfxgb7C1CjTk5ypGCuI7CABxlCnOcM3T53O6AsJs+OzgNbtfWKRI
33hEeyfqfVF+qJr21wLcpVJguNXjHpAX+X4mFk8GUFDZVQA0/1P7pvQyCGCvGI5OlmdxGT+JerX6
hP8sSh5fgBZvIz9AyScIa+5sjZF1o+KKRzfbU65MCnvDbUPArA6web9V4j4WGkH7yH0Kh5aHWoON
983IsyWa7oomGVcxcpClPbN1XoJDkDCpZ2N5/GZyig/mgFbhkAUFPsMq/RKZdYatOal4gwsPLBkZ
5DKNaUrqQGbBijYj5E9m6/3MDdF/GtZnRmrpwX/CgzCRIrM9qN/T/pF7kuexih/rVNDw3BeN6TBg
mIzhQnEnVZaAuOoR20htGmgdxxlKQOyldg7F6xMqZfom27BMEpycgnzOzF6bZ2D51/4djCeim9e6
JvZXTEDEZhy1/pow0TqiVzCS3ZqbOOjZmPDszIWWp2QEp1lse1Jg3AR/ERRTM+GEDwkb812nvo3N
1KOTwfsefYAVn9KtxJY381mgaDVKPNHJ87EVN32o1FixoHTimN2y7FI5WDwhjcwgWCPo+DKuhO/X
fGVceF8xSmxexAL44fSebdD8OczWZZoWbdmk6poRZAw06H4VZWdvZXLAKSjg7D/4G+YCrd3RGJNc
brv3yjfaUAlKAP9SzyhQEtsHs/oQ5YQsBghSffw7+66v1SKIKc8M8M3I05OhoSbahrwJPRT9FV4N
1EsLLCfLx5ui+Kdo2cVAe/DfxGXnVNT5fFED1cb7PGDSz/xBvWgHuM08c88dNCwFufULCMA9tUUZ
z9odeh9xxIEZUqqfe6pJg93TN0stakwApsL92QIT8rPmvPWuxyErvTxdRK4Urlw4Ab4P7sttWk2i
g4uu/ZqZWEo4B7GZN0JiHW9BRjYinV8BjHdMkgMJ5P2fhPbUglkfDpzt/SizK/D9AGR0Lal23LNC
tnoxM79sXp0ahlhV4XeeAgeWqbRcz3wjdprG3S4BTpl347V9Gq0WbSygnSMPKSjtAtGKtC1O/gyR
kDEL/MShoX+8ErQ1tsOGYYGNHnOolXSEODgqFzjJ9bKvtbc84mfV3mAvi9T2PMz4JLqTkX078cox
+X120SJPJ55TY3gDkybZcNOys1HxLr+0E5zcIm35tyCIJgWVtEpr3VsbK/tMbgSfeOkqqZi+6wWO
43+u4xupb4D0/RhMNEzG5f5mM4vJ/ZQd0t4YcAU44ym+/422LaKZF1q/8k3BCZtE5T5e7gqsQaaW
q9wd5vnVhj0sr33vg8q+m5g0qg65OaIXe/j22LlNbPQAn5x9etK2PyoqoCMweC5aBEyOfnVkvP9i
A26W2lVSWQOCOv5boPjgyaHZyYKNBOS07P62z6pYzhUsOE+AdmchTqXhRWhC44derb5B0Id8+QNo
+viprQJknE3OAvzmBmLD7IvXSx6jhksu08k+h+CNlft3Ka6/CyFA28wG8kUey79eiVbA51s1KXxv
gLkvsYdEtE6X+oL/wCoidEh+FFf5SOdOB3vaPg4OWCViCNijzAAA8CiUlWnHZL6U3dRbax7ojNIX
9Ynb1lJ3D6nX6OyABsPFFpVpEH1J/2waRvmO1taPCSb/ljC7cyrsMdVQM/lhyvAm2s+3oQ4+USAj
0qRVGQR+dCNElNbmSVDCRRjYbSLm1XNtix1M60u/kFarekhaKw7t5yNUEep9h/b5Nkgqo1pMCBVr
eew3CF/yrN/ieoZAAl8VyA51avES6jctgMmcURhJ28z8LWiswSyZQ0GOZtiVEA949OX8fkXVKnym
dzeIERtJ5C88kH3seT27HM95Zv5LO1AJtPV7g6EafUiuKGd/+qsREm2ecWYEPwAq9rv1/4HfmsGg
DULRwQxcqbds40cI9lHDXV+RaXPxcZ7x67OvO5r+ThH4pX6r0lu5xfKAov3lYBpm95oGtqx8UqCZ
GWi0Fi9Nlx83Gl+p8X7kQpY17RgHz3EyJMvVFpuyRJI1wQHh0+tnxuC3YndMe3jUblTlemR63MPo
hNs2wGULQTieQHJUKk6PYClkI8OXxAkM23hywSlrozXm3qz432fRTge9zltPRO4zgSdp0I4RC3Sf
pY2H26tX6Q7piF3L3wwPrHtgW92R3ed720mp3HvJ0ri3HNOPRXNVC5kMg3PhCYNmS1zp/TD1q0rq
xu0n+GiUh82Z7P4RmYQhnCea0ND739c4VZsmNDJAWKACY789bcIYdL6hv2YDyJlTPZ/mvCqeh0IS
hC525zTzmaStnZnSp3hBEyqWYhBez5fRhCgtLZT7UPNhBGRV08KGFq70B5sSfEVR2Li+WJd+ZleW
vwr7uWMKTROlGUsNZjZCshnKgkrtFJ3AkIqES52pCrE3dksYyRUkW9Jg5XbhBc6tNsBsCKz2carO
ptPfmfn9XvTQyq7+XYdpvG1gz5NLyd6CewZkZtxiGk5B6uzZSasu7Qlpd9J2qTyu/jHQRU3zLlzJ
7RHrW/BlAAooNiUnV1+AUR2oHpQaz/ZaQ9/pmw0dgzStb4On6clHrtthz64AGGSYwv7a9NalZ50J
7naaYTlaY25+Uaym8lcj8MKzGdwCf6MHzxnvjGe5FhHYvmJ+jbhygVkSoFXaY21XGfaL1aEynIWt
VNfP0SE4qLCrCPrD4uJ6BVWtrR7KI+8YyHd1+qzoBqK7pF9XJ7DVmQKaeG2FR8xMPY0JeSYHvf1v
v7jMtRM77k9mczqsHgVA9HZD1T38ONDCbcn9WrJx8TSbALKe81plNTmwEFvPSUuCvw4R0jFPRT/N
zcnEG/kMRvu+iVUE9qMC+JvSAleXf60olj6Lqdnp7PEVgIMPGljJyPoypkTfquUju8GTnilKHoil
Oe0QizXtxKcv/JQxr5KbZ0WifGs9dyUWI8agKsWWouRjrYrg6HnNuVfKy+hZgC50nqxQ7JdKYVQK
MKUS9TMoPEocaHEa0G//qdDbxhL4VRP2GFYc81Q/XmUO2u1MFRzuIW+gvwDKepizT4xSBUO9KMti
o33hnLke/bBwwvoyrhrjVqFkVcTMj8YkEfD7wsc04TqCHAikGH8dqXDBirsNyMvM7+Bljs5HqSBp
V83O5BxoMqDqo2qTZsAbbj5k7najVYRT/OpkClbetOh/ucwMhN6EAV+UUxAYWrIPBAmvIxcovrMv
4sTaKKzANLsFVhVPTNKCchhuDaeJFkiCfybk9wyD06oAXpb1//guINfAWAqeR9oQMnlcsBQUvQsw
QQfGRpEC/y0AUqR2Fgn6S8HTyFzticU3GHP1AkZebqGlJFsdN/yUjUpn03q2aRIrymNin5vgchcD
ar9Fwx4bgkrShnPAHvzpqpZf1cVMPlTcljfj4IhW0m24WrP9b9cBRpx/p7vdqPOErSotlaX7w84S
EzQHcHEmGsVa8uv/sy5eDV97ZHIaF1MKfbsmK5/IPxhsmOQIQtEGe9l/dwoBPc+LRlAZCqGUnvIx
sQzn94ETyNq3/lZnzC5gydpznrhmJAifr+7v85Pccrl8uvx/BsRcCeqvTssrSZgP4HicCpivmToK
FdfUGVVRRP9yEqwkb0Yjo8Wwsp8W0OcZVivuNGp/lEkcL6Mqy2so5PmdgfV2fnYj88X4boFD1Mnu
SJGlpLqk6R5MfG2ps92AqyVN0A6Kq4ODkvyGYC5rpB/s4JqlHayaFL0JKrrNXpfYOVaFp+eE1ckA
esMniLMadmD3+IN921Y3KVTT3KIVFc3pozXXHudL0+SfzxKYzxHgHflBeO4cb8Nd5lCsTolDNvTS
tx5589Us5aCGM9l3ypgXWVvrCJm5xilY8x0yKac4cTdAeaVT4TqPYSSyDcmyCh3BDqlclLZkmh2Z
A5BNHqA6yvuGw9BLqwXaL5A4vNt453F377GFqlhslMxRNVhWkr9NXngc5wnK9EyfcX91nnQkbIin
c6G+x390sj5WHAr6SGq/fPt8E/eI4zuyT4K/OxKDkhB2XuoLCqDGrD093KSarlY8aoRMYU2nVUqR
vriGzOmgPUQRKlxmRPRLNnjTVaLGFsbVQOOUNPCfxAvrPAJN5RR5c3OpwP44UnzUeJFpo6FRb+JQ
b+jiuk7LROUsrsDjIbYnx0ygZbDyKuJ5+8hREIi7JJUMkmqBMQc+NMWJwH/IxUauFC+6fEHPpd4J
TsCtHSgEDur2/A67qBJ7PGQIr8xAQHVWGj5CaSWo/VvyMh+D6g8fMRQj/ESjdB4fnie0TZ8CU4Ow
ja2FRwojc9rZzUZaYzbGQJMekre7NdMDjcrOd2WJi3et9Qw9OgpiBWwST8TjEbNG1RVllSeSCFfz
0s6jmmA10ffAYYwpvWkuirOQn5+YqKTEGR2+CAQvFBxgYxDq91vaVp03VtzBdrwvPjY+vJ43oPkG
SNQJvf4DkRUn2IL8HcQj1DsDzx9aYvVzajINdfWhi1geUotT9G+WXPB9cCShuxAkJN3YG1bZnRLA
8709XfsnFeNzc/rZwCLaxAx2Ce3ePEFlz77RKogJpEfJ5e5cqJfLp1Lv1pGSIg7+MzY1Y/Y1NCPZ
JdpScwhBSMxPxbIDjj1tkNRuSJxgMSfRcEYq96pC2Wq3PF4SJOQ0NCQftvQ2ORDZn75tU2rZG9do
9MbiWh4JWjtkMDMwIrCy7SrCfHrIyiuENoQfDfRzS0vAsTZz5MbSp7T2wuWNEKYk4Cd4wQ1egye1
6tIeqwEAqOllJDnzP5U4vcKUYhWWtBEy8QpMk/pBy3ipbeHcwKk5CI5Aobbrte/WskmmHyRXv6CM
Uy9c1T4fD7ekm6KsjNqD1VGiKqs8tW8rGuzisxbyvrvlbUWr/TdAd3PDjUq9mYI6llCfAb9QSZR8
VQMmHAUR1nEYVbHUnnvr9PJBuoE3RG7nQPvwWkqgf31kiQVm8bKrq4W2l4qAoYsdT6U2K5rzGsLz
U4EAGzmIJqQmVD+DBhd58b9KI3zN2ZSNXP2W2uvEa75sThzTp4pWt/H6RNH98IJIzQEhTX0xeI/Q
LqnFBAOgJ15DOd4lVOQu0lwtrsUcrD4C+bfA+c3fh3ThzuQXbrce+Oo9ChHidbS7+21LRASqc1w6
JOLXenAiPmQy0X5nD1jhsk5LBD5OtAUp0DBzIxZAZxjFfn1hDNNpDT0JsgnSDEsJPpbskpj7G6Hk
IT2c64DJjIEPInN9/rR5q8uvqIXb7NA6Ov6GiOXRyFcdgImK5b+uF/9MPL/dzHswUDWrEWjD66Hj
PYgsqxzYi2t0Fkt05GA6nvG289ceiyOXIB0utZ3b7zaRG4LmdnZ5dgVNDr6QQRTSuWmvp+T8tafU
xEZSEaE2GFu79emoznsujFBTwwd+Geaaxx3FIlLsjhuFIs0yXNK36lA9ODCw5Qvh4qOTdP0nRt1B
T/K0hZ2g7pAO4+devHHj2R1M0AZYPDJY/TWS4V/Qtv2E5JCP5DCBURDhr8hCs/ruRWoG1kuPKgYU
CYoofgsE8Np9789C6qefROiwwlMd0mksu+rJncqRXxoTEOkBNhTs6wbr8R923dF/rPdI1nTrhVsy
zPnJQnbHShPp0r58CD6p0WMX9qW9GL6NBwPBcl70zoWNceoxoqqca3KDbBPR4g3c1iRtugzXQJhu
ZFCCvSABzjYQOVozzkzj5IVV38zDv2ZvR03AFtjqwLDwgNhR/dyJa5g3FxGZxvcPdMjMi+6Vj4vp
iPlv9lRoftqjiAAH2QzBxWy16nH3jOOErGZeQ7giUxz4YT0hptvGe4Jk6vh5P+pdPj8tOSw7MasS
ZYVU0MFEzp3mfoSmFR8jMw5daE2Ah0fsmRhXMX+xswsjebF7V2S5UQRXZFNFTPDF+OYu+p12jtrs
O8c3Bgopd7wW6UZZOT4KZMOU3AETwiGHR8LiETTlUzuM2411LlLXKAJVruSW0B2gYlkXPjnUf4XW
oxT7ly6ESn8XNXq49++XmH5pT7c26/4C34PxBlUr8IgniNbbkmDRWvAibcH+L0Uc3i/Ldd4Ke8AC
3HbWnT7+PknktwzL+8ntu82NEzLF/bqWgW2U9I4gFHvZxPCzM2aubQ84tI8VkaQLCtIvnomj0k+X
nN0HzMM5dRZ5DaxXtN7H8gWWOilvDNgMPZuUVeZjJLdeIvK6m75mwSICjy+NyW9kP/bp9A7dssX0
2xU5+m1jU1HVUEsXSzKLaxbsCXjfYlMvacRNzwNX897H+C4Dvi4aTo2Mj4nfAPTIWJd6IhwCWvAv
1/8Eshx/UYZL92nPzSIq9kwfprrVF1a8Ml/SwQo+Pr31EP+K5Haasb/Dr6Q6s5HjNcLStf4NnVQH
inwMpOA6Kqj3cLBgyWPyukFS4AMIsLgK+NuKoTmYH/TcmvQaenbDO1w+40OxdB0VDLKeJIFKr3KE
PRiDqReDnesWCAodlD4vKKoepZqMwXrx/JivU859WWOnhxzzKOs2T4tqbm1YXazw6QdAHtDgiUHi
9HPjKjfRCUFq+Ns2vT+I38diNPn9bmRb4wGNTN8YdAtR/zoZveTomO1rse7SDuCk/vFL5YSw51/a
ea8J5UHMUcM1I3kVUnKWzROrNZ9yk+8cLAhRH6iQPoxI45vDqIBAYgsfY3RkZ9hr6+vhLE1MTfWC
5GU8AM1gCPBSTsJkpjZf7sO0j04y62Z7QZZwsUoULVViH6N/Bu3EkKlHA//A1m91M4DO18AxyxeY
maYQMFMbsavr8HuzlYv0IkkTLFC4zJ8Q2fLR98woYX5w/rmTlGVJYz/UGZi//71qsWBoA4mDNVri
ISo6Eqju6LI3K0t0iqWWZbNLNI7rtpwPa+tRjElYK/VVGdb1M6KJRLjPBMtqDyTrEti7o3MXts3F
8PlMQHVGimCQPNLi14U4vWfnwFGXiDW6WtgQ7mt5H4ylX7R2uyP96J9ftFj7v48CvyJI272KCA6J
HJIqTzJVF2tmbHSEh5DS9B21Gky0h2j8KBwi4cXqe4rwQfIEJAQV8dJwkRDoJCNIjFyw+9FDGJA+
KUXRHKb9w7/tQYj41YIW3yFWW7pS0AAWDkUV8wAyXSEHBTO5afijGpE48CJSu4tORiopYbJ2Cke4
wcJDOUSDphFn8LJOGThEd24qUc4LftXlkJ5TMeU1J7nhJFf+PKe9Fb2QMR8fUOtNHy8sZvDTxh7T
2s9z/7nUKHGEeTjbRyREMs9vXGDAOKw2Q2YFU7B1yKT0o63nDfhhcSQhtDIxQrmDv2rLVA7fnJpx
26Pf3Ub810C12Bn+FY4eXnQjdOmbr/2uqPl0gRDxiChtojBpcNjDTtgxPAj4JXBvFE2pvD7LdmWE
ghKdqadVxfQTEjuKsgJUhAizjyF8bPEArlH5d04rvNbHK2df7RfELa0yLVTn1Y4ZXLPXX7/VyBxG
qYhIeIqyRfrtDehPgjHEeQUsG3wMuVQNN6kZ6MtIfnRu8lVVOj2hC/+/LbFe8FHdYh2gxC4KqaY9
v3/lxJmSwQvaEvfhw+xwn3AOHL4tIPW5INdbqiQUjByDDvL6S5GWidRjWE8JgLhdNm/nMPV/MjnH
enh1O3W7teJapNYpnYgAN6UgR/yc+iPEcTnCaV4dKWsvqo1yA62fIPtEG/ZBPbJd1nYPsa9uVSL1
Ck0s90tE/a9bYQkfy1djxAU/N2JbU+YUeMfRPEhH6zHXkCWhaGdKbR+8TlAf4rgLBLHP0VNxNthO
GHng/kk9LQVB5YhDhc4IwY3DeNCSBCno6UOS2CBq5JUqjR73xHmTU/0Xx2Fn1HD21xPG53ie9Yvo
+CE9htpUd8p/EGzSG9JCjbtkyT2Z656QbRttXBf3gKu/fq5TC15nMF1HTy3SSQ8Of+gi48LSW1FA
RdBLX1E3AJaMb3QxoGsfLQauiMQpC9VdOA6N7DqI4njndJQDRYNdsphcGZYnE14Pvv+p9RtshZIY
SpDQwXTTGLZvWeJIREXSfYWDbQUyeo3ravPfhYvuHMOz1AOrwdkq268WDFaXDPngFdBdiUJPmYu+
5198KGtjcJ6PZ/RSlYDdnWMUfmJR1NrN5My19/jfPLp9URFvMSdweaRs+Hci2zj93FW3TCBUa6O/
ugEyMAg2yA85IdRpGSksFpxk03weLgq7iEE7f7fIiD736hSZNevTOhIhQzDOWBJD3npYYtUGc4rA
ZGkFuFn9/66XFOpRzxgFmz0nn9wJY69wMZu53pu9yHjyJ1M0AXoxoeL3rnfC/UK+OIORqzz2GXrU
txnog4py3agLohUyQmwb26Ln8NvOlsFdQaDHxrOmLL+TnYGR1rSfPEkMqiqKSSo2heIo/8Ka+Fos
EOVsgGQBpjTCe9JnHuOEu8GY3lskWGWuZ3hDOXRHxI8Y08xC4jy6CfZdPKTHsTbopdAB3jJ6Dxup
txgs4hfoFLsKxTKzvlHEmZk33NayA8gWBFjMrf12ih5boRa1Of+VqYljnyPA8TRhIMAib/MRbt/a
ankVgQXEBfF86PdSJa/vuDG/JLsOz4Q4vpn12ocdXzfi1/ZO2Sb8Ha1JMCbln8ls4iYXhljBt9p6
rsr93AVly/HJnCp2Tz/YYDZ4ZgSMo4u2IBbUvIC/VTKPe+8Mgac69DXe+sE+wR8/mzUhuF8j99zL
UvgTGO6gJW3QoyrjDKz/OYJfRgIiWwgVXdT4NrwXnpY1Xy7KC4jZM9YLsZbmest2z4YsMpBiWnlW
YzoFJCchCCx17BBQJRDHuBLPaCez00diGOUjGmZMZCoyTunCrXDAS6cSt9b4zOudbWX0hO/xlwRw
ldXzg6JPrB3fTZeIPOftKPxv6z6ChiGaStku0dlV3Lc4u6CVrFkXW2RFxyqwz+lx5+Kw6SbIIMRk
f3y+e4ik3e9j/zwLJywKk6f8LHUjBP3KFvtW2z4IdEljRHfRKaP77rjXgoBrpBZ/O0ZvSh0jYZJ2
Hgw/oxOKI8eNrwtoCELIVK3GPla3EQRCA68lMuRvhHqsiFOrAlHlodO+HUVTVa8STPVPBOskFjSb
CVoB6XfUR6tV5gvoI01jz8mMLoqixIk/j1ZXe1kXxq/O+21KEyYJrRVIs3OhmyKT7ZA0CMXQo18z
8szE7sS1OE1RHUHl6bp2x9JJIrO51kW79kSfRXN61i+lZUmlCOUMnVdtvzULSHkmEGDoaa/EIDrQ
h0JYqT/qGMQ4gyqYOM+c7EDGi8jIcHQXRLUKmFdF3CSmsRvA99cXqidyBuEkpb8WdRHC6Jt1iF70
PgyoupPhvqdw/JlQSubN6HDjIW0LKuNn3nW4wWBbTXOjkC7md1bdcjS7btLlnhPIwXAly0Vw7VhD
cQZ4ZjAZvGuKvvkmOAXaRdVMMQ/dl+UkA/o87Buz+miHEQVrdHhrouwzYCC4zSEoqUh/ZxNK7mTF
O1FswQvwO+32LAvoaNmJcoC8Cu4xdprDGkPqOh9E2zEHXiduOVSnwg2J1KJVy33hTt5mvV240Ng6
iHIhh5c/cvz1CBiXkpSuKJT55mmQmW7YLjDfURdAyPrWXhkG+w6Qt2Zl40UkVPKGMkp+Lur4eqkQ
u+y7FWJ9la9uRSTj4K3aG8/CmxcP2Rs1OxbCP8CxrJTWjgaqZTcYPMjY7t9kfGxdLRD6sQnVL3kd
1ThEAbMGefbqsgWIjzJBYBs/Dnw7OapIAKqvHXttz4R/8EsuGixJ1FiPLoi2i16g96DQKQQh52/q
GMYGJ2bmcjfh+tTFM7HPw3GCeNb+UdZ0eHiJy9F7vmzbuTbIvDkexOL6ze3+bPeDkAnjCCfEgSeT
AP2BOn5C1KuB66/NEKvgT30pCcAXfYCapqUYx8nsSdvpxEdoOHildWOsaTg8Xub7JLVmAqF20g7D
P4v9sIDzAt1MVkEHuihI3P9oNZ5WGin9GmTbzp4M/mN0PwqFcooR90w280YrxvUibjCZ6w2zt648
o/xZwMZM
`protect end_protected

