

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
kNSODHF2BA8phv8L5aZNyOOK56HCcQ5lgKBxF8hcTzwkWRF6WnOKZaH0cAk+oZsvi02J9SlLLySq
oKFSyBG2Dw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
df+BuhfNWqGLyuHwX48C4kdWet0FAm6osy35ZO6nvLm9LeYvgiC7d+QWQpEp/leK8jaqvimQleVB
qNUNsNTBZzVm+VZnT/+N9fzr+Kn5brl7DACKZQsJ/J0EK++GrIymGQB1+7LWFg6RjvqxHctXSERU
pIxXjKUtzcqAwrR0kd8=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
j4klfuw/RrSoDKuTiN/Si4GPF3r+1zWV61wAeT879HAyso4ajbQGVJETjBzL4XBayVtdsViewbVc
n3EWjppKn7DU95ziVUsafFQrG5PCVJ8TPZUJisZwRf1u8N8ojLSjd7Gi7vpDvGySyTXx9aoOQ69U
XzJmTqPAeaivz/FLFyjHWzMuc078i+06EYa3j0uxrNsDH6/IL5syM3QcJV3812LlPGSBhRN9Wynk
J5AcITSvkzy/dqcKICGyxp5ubBr16BEoG7l6F/VEXvTJm/kJnHW75YZ8OAQ3I6icKjHkLZysnDlK
KEU2K5X/pkwYnpID2ogdwsEuEQr/xxo42oEmKw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
AG9C2Ti5ZMi5neBsWpJ1qwXbrUaWpaRO8Qn1fL70JVZk4SiqmPlFkL5Hz8GrFfE4eBlngUFZoung
TTZ2IeyMWjxhdHHDVda6+BqJtPiX+FBQnaCzRd4VBLDnB8KUn52eheU5F9XtqqkHq+oJV3U19TRZ
Rq+NhUtknFhYrHlVXfM=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
TuUXpu2xk+duDJnZONHfYiEzeCuzIA9y6Ut5Y0LAE72Cfiq+aIEHs4lmSaypPxj5+E8SKfd42Iqd
iKQPBy7GWczcAr4hdHMLEortigKfhxQvyiAB00CsQyuj949i0l26Eh+7iirhYh907kSXNLc4JeDy
uXkHZzsX9mKBsIZLMO2TtO0R4ECsHQbqo/hSpi0B8kY4ucdqtZfLpEsAJ7G3XH1L+CD4o7on7UAz
BPPpoVV+VIZR6heT9EgSZTHhg3uYl38G0Ezv8g8s1cbXnSuowx0B9mx89vkctBzRxFOLnzsFdBr8
DIKQCrHZfdOhrNHz4ZkgOrKjCDpwEkMA4ATVfA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 26464)
`protect data_block
fDuRH4YlNnBt57OeMbg//diTrcGT+SBhlb+fOY2IgXh5fFRMMyIgYrZjsPZK4vQNz1PId5Y4koZ2
K5Ao7jopx6FuzbfVeHGeErmHfIUjSzytncAHPkaLrXUK/NfvK1X9xoFW5TWxk3iyWpAt7g89J7B6
lJlgyeQdX7tGhE/F2D/jTfnAEYr96zPdwgZ47Yrpro6p6BQdQZ3nPUr1gUf20eBqfGTa6DjdZBMF
pf7+GacPqjtPyk8JzUL/aIhNULXc5MSONxneoDZVKXfn0z88Nl07644HYs/7ZoYuHQQ9ypF7zf99
1z9VQpvmKpVjGifmiCeoEkpKfO5KjOP7C2y8lXtOwfb+eks5J8BDAVHDqPUKDb8NKNDXRrHsJnId
71R/5ZfaNfgINyPrUdpGNo8elkBXNg6tHSJ+vAv7HVuxDthNHN9V+pO2oL2dniVCp6D0SlGzhEKf
XXW6teBfIdJyX0AZ9v2MKi6lsPq2DW+RaH2Ya82bhwXnShGrzmRET3tdSJWIbwKIkEQHN+iw8npW
/hR9lsRLZsrN5CwLQhJiWyGI3Rtmur/wPGR8y8nDa4p0KUTwcB/QPEGICNXKMy30Oqeno6DcAzqs
YSN28vb0Oeh+oFWKi4pjY/Kl8gUACNalyYRNYRXGOYu1+AR/RmNsZmdBtPqs3WLXXVdovBucnYsf
urCAB7CmQj++l32zs4QzljErTTVhcjkwlpsvh5bAHzoCtHhnOX+L1ti2sgrCARx9STO3pSqCl7ke
kz+0poFs7HgfB5kkIJMuIUocXZtoB0sW7Y9RVF+dIOoi85vIGQViXKHWyYMIfdrfNrsWPEZ60luJ
32zO4UPlbrwzQ4AgLJiYylkSya4ADnypr+g9QBJjIil3n1BtWlTEwBrc1iz7m9G2X8hsSVB+V6A5
WV4Ua0twC1PHvPGKR3TwBezus1Bb+Q97rpyPBq5BlXh7JRR22YsvkeOW6AHhlMKssgGCbBg+mT8/
gKWdzJO6PdZmqIUJgTRz4lmsIDFEPaK9msMZG1COnzhkD8XO0hAfTMaIc4sAG9spmw0uLuSS5oaf
d0mrYAJIAzTVJyS2zWJIw2ZdgzNcNvdxhKRW+NVIbEwXpJg25YFDARyhAAazBHvJXcdDG72Bv1YI
Fwc1+jDbbDaEe1jheClu9Je6L7wyg+5AckhAkCEMA0S2o/VEZPpCHo6z1fjbliSW6ULRTGGLOo99
1ziS9XH0GMVOt3c6vwX1k4u35SyuVQaWiI/i9OPpE3j9WH0zCmKPLi8WH5jYxc/1FYBt73JcsRLe
roWemj3nTcqTu4GVH5DhfLaIMiyk9grcFDeIMIMDfmN7KgV9IZOeAgZd5tqK1qxZxd1+xPGuX1bz
U5yaVWlaMAuO+8LwNf4wkYbec7yMkX/YLjYebtn9IPGMU6tsJHBjp7E/EeG04s1JzUFK6+H7lKtz
xONGdBI2JoS2CU025WJPAyxa61ns2CLYGe2ug5kc/Fe8gSWnVRg9xiMcKL4jo1H7aOv7cYEmj4sd
8F+C0ixGS/VKesM+v9bYTvtRGP5jJN6HtXZa1wqzFxq5kIV7bW2C4GdH5kuLNy2gXXUY9YvFRZum
fFJAw7NfSOhjo1n2bG9LpYfj9vK7btiP5YDfhxlePCkeVdYrOmNSkNjXnBB0e7RzEAYXNxlAJx/p
hZw9AaWGPSoglKfX1nDd7oIGIqUcXJM+BSlnTdXuCZT7utAOHiyeux5BO/KSV4nhakaPINfmfd29
PlEhFShFsusWEFgsJcpElmFqOoGovw+58OvI045LuwYeqddWLeDFl8iYzjMNR4RPcBTmUqsJfyt9
wP+CHZ0a/JtLkiQp+aVMdEw6PLqaBIgyTqth6xQwiNWJxTDFkXK58pkDNa5VM/OIP5IukHlYGnIp
TLxWTcfaiY3o5UizDwDJ4gquzhnkkZ08XIul/mZxft0jHL3MEEZWG3G4+FNU6Jbh4qx8apERS3zY
m69wzCWEgB65rKuJjLSJ2sFqDoZ6mu0+jbRg/NfvEaCAQu7d8Q5LOxFHMYFuF7qXpcrypBOpjsPG
JCjwIXb+nTLXl2TzkLSoM0rwTCrJB6TtbWFNPmiiIZvfnn+SbObNyVQ9O2C18J2Q8l+mD/Q9vtal
D+ddUUh+AS4xJeddifU8PxwsTPheqMC+jwv3ABTCuBS2EX23Zz77/mQPIbiP4LIekUbEleLruZqC
jXfE9i2D+vOOyvr/ZzS2/hcdzRTftlErNp0e5yqDSNwa8k7a7DhOpcVHSgAJJp84MqETqJNO7XOG
pAPxU3+LSP60nqUIq/kBMXTTdeSTi9WP5uuajDPTUnyPeFptV+215HsGSx2+UkTonA7+0BZ94U5r
y95+UpOf6exy43Pv48nP9RvXbupX8vhCZVwxUl+IwMB8zz1LvEnyRsetppl3R1bciGrkMyPCXQPL
X961JW89c0/1+vEA6bitKz+gE3RW+59jBez7w856+iEoGq1ZR3KgxcSq4ZLkwdNwhErBkXyEi6n9
5gTYYLAuudorZqx8lGDn84xw0/Gw6E7mB++XaUTPq4nK045hTeTfKD3KuHatTUtf9Z1TJM2KKakV
luwKE2UyFDgUueYjrQCcXPxId76VzlIyczzOBlUgCc3XiroGUZD48lx1E4vYaU+0YPbhyOgel47g
zgUo7RiEnwPeAgO0QBHorvf9Pzjz76O/SWM7tjBbdLA+8dBgEI7MWhpIt9xD44xUrCxPXwhLZH92
nwSrMRByrT7wiMfkCDrdhS6cbK/NtVduFPg8zQfGApRiPDrTvPO7M7Hean/jtsxJAka2du4xK/KD
QBltXRckhqmfHT2gWkjlkTY+9uB0ekcO/aleQHR0RQEd3kron/qANhvd975BNSt51cyW6gKNxKoE
0nMJYJSsQcWZELJpKptSRjfhPx3bWh5ZAmJov7D0VrZhv7lcQUZDtU6IxblRrKnbLUZ2qiG2VV4/
rL3+2R77M1mvyaLQSlmY1MqxNnh2+f9RYtZ98CJFpV7GHkONvtfcrQZmR5Ga0Pkhon5QT1jrBKbd
ZGFOOh1GE3m4v1MlgoJ/lEiPYevAxmsk5x0oYiJtADH3ZvuSt65SP0W9aeVqM1y8NSwmCOUia9mh
W/eoRE3QlBDjNar90WJqu8Gzg10+SKYXVUSfwis050cdJeaCm5BI5icoBFpoHVRhF2RCzWlP/zPl
EhsBR47//nqCddZj0UHY4C2zzkhc4VYJOkdHbvdIDc2Y1KneB1MiamnThxVMOA+UXJ+jfr+hYf64
37emhlVVpNUPWeq9Ux/TppdEtByua3UhDHi1C40g6rOUYrfWrdrUe0Hdh3wujK5yzPVlIPMW/FvH
J7YZiI9XVgBXEzyBl6TxFlKW8kwdauD65caYNwUz3F2HPfnGE3gedhxL8ghR63oSyBlupH0MFDah
vLOkWWlQxnwTzZSjut5N/3PQ9nLNMqGzExmsFsj8PxhSi67jkKhi2b4U19JZvi7eS81VEjqRGJlo
rHw+c3f3ka5GhxrgGnS/TDTgq+UV5F4YAD3sJim+5QsK8f45/1JX5nVpDpbjOq6uU+PSFeFc9NDw
2mlAdAViAlI7Z68Jtb89oGBoHPHPqmQ85RNdEldd70vKBieTO9LbYHIT77/CZ/VwBK+M2McBaFux
6flNZZHiPXj9D9fcSBrgHpJdbyZWfbcRRiCzHQXTIkoYWBxPabJg6qDtrAsPvfd9V+RdRHav8BDO
V7XB8ewp43GcAwoDZUKa82lZF8AlGBPMk+yTL31v1QyjV3D+uFWjdPWyh9I9yeKtFFx0HpdsBSJJ
iwgQPKM9s16yQCbFL9rRpKRd97zN4syFr7eAfFq++rSRYg7pOh/VkD44WJqWfsM4fae5QbyFVagi
ZMnkoMOQMEM+NIjwGI22eJMpVoMFB/rEQ+INoxMwOW/5+bRUhYQ2JvZr08PHevFO9qDqRmswfxUc
cJa819+QmahN7ksnsveS9OAVzUpaIRtBM9a45qFhelhd9tUcwOppKe5HfGf6yDrgFqFzbYIScJCU
SUCtKwNalGjut+OkjM7UxOyVfOXmHMyU27ySGK7EQz2f/souwFPQLltJM7mmv5sOAIHYunWEv2n0
d8U+Q8JvEdSFCBMZPLpqLTq2w3ZHz6ENQ1aooQXB0/rn/QzuXx9uXHUSecZwypObWR8CXY9D88zr
evbNGbh8RZWLnWEV85qRySQXNiajAtFU7JtbgDfY0bgO7frro/72UGLXhl7PA/3PA3AvsMUFq66c
/33e64UGOxTrkLnyqDAu+vQuMDZkqQwhM5rNGc4sH+W6a3uUO6GTyZojTWkDKmuN1F7bRZIVDCv5
v1ImQ9Z6wahZl860JttQy5i7bF9hQvxBPXmlC8Ll0bfFDDoaqdAs0NwK2y/5eCn7iKszrkyL6wVB
4YiA/k4oY5X4/WVOIGaa7Yvoeu0Cr9LX8rhhyOz6+Ian6og/CDFO2MgyxN1nODtyoIWMe9lC8N78
ttPJPfe3zRnFH/6mPXDGuDnJ/srtPFPMEWkj8rFsMDwmC61aWOZgFRTx+54YOqC66BpsSgCK4hes
C8T35Rujostl271xJUPQIEp0cxE+FsmHmRRDYjZePJywQ0FthaspdAFRVeU2McXnwcUm/QwWUhiZ
7CZXBfbmk88IrcFhJXzy2agkYCa0llljgdciNtrzB5eVG5DfdCtFbTZWW3fNYSzVIBLFup3UgnOQ
gsW+iSvGFS1B/Zbo1ERPiEGEGDeQIZtm5Olg3Y6J7mntVXHYIf5dAYmy6+T8AD9+f0Gbpg1VA3cE
IwLvyVZBlms3pXzcB4V9csCAmfFAQ3c6kR6Uoz9MDo5/uDlWGFamnYkjFXUls2NNInuUpCFIODvq
w2/w5j30XaYInG4j3sGSi7GjoXa+k+DCKfeR3RQVvwDPL2bu2NWQAHEz4b28073RCDTZUznm5yWR
5/XZOAf0xhtSgrpYhCQIz/jLZBYlf0m/saulVVYy93V0kmt+ko+eskFzz0a/B4jEf8YLKP26YY4e
VrwRXDTacV5EhJgwzpnE0P4UN675FKmqoTE01a5qG7OFzaKuNk5tf2UA8t32uSo/9ePolwCr/4hQ
YeGp1nnhk3FngnogWK/XKOBf//kz3DdBnll+2OSddb/J/dT5H0gcKF+w9aFOKYziPlRPAjCXSQbs
8jY7cKA8Cf0c2H8Nvf0+f+JSVU59LwrTJvRl2R/ai0yFJ+oxdr9Yfz0XdRt92l3Y2NOLbMONsMlg
tpA2uGOQSVcTavcjFChMlUft8K2XbblzB75GV5jHnenttJI2+XdHDFvaAB9BCYautX/hkz7i9rNv
c5fcGCzAbnpPsKX7NOvHhqieD4+tWmo8S9qgiSZpkJEPCRlkLteavd85Vz3BjkMp7wVpaKPevgVh
EuKW687Mt9Fi6HhfBQwp1s+OEjQaXWJASmRjk42xrE+5AIcCwqpvRiWpukfUwK3onpssVjuCZ8Ru
cvIy8UX60z7A1P4PHi8uqUxly/MkuH53lIsARbH5L1iM6OoGuG8WGjAUymqW1Y6hWaIBEiOfkcnl
nKvjSZMRjp7uQ/Fuo8eN2d869NXaD6aSVBtttBf75Fm/nfEcJwYhORL9OQjx1iTKu5+EJJNIwaoA
sGxnoeJkbGUGB/6Aztmilcn4fXPifKgsemGw94aZkSAVKIbksGTtKdxY85+MYLcQCAHH6DOUU8ox
3/YrhxS+rKOC65isujdzx0Pfq+E3j4Um0pOovGyM/jY50aQZJ2pE0ql7rhomF8APM08CuXfZxyDA
0bYuHuqWRGCmt68tDoXXyz8QZdzhVmjXliraf9I0FH9CSAj25gKLFlJ7sbyUVUwVhfsqC7FcrQlA
hFnqUbkbsLxdrUO/OjaK0IRjusjZ8d1eYhtYV446YyyWGN+2M1Zz0RYXKmKkuss7zm/WR9OoTeGv
xawKycSaE9Lpsi1f6WdX5Ytc8Vk+9540rVoAfyscRh6xN8A8aPLIJrtvV18+NRXqLRsIf9V6hnZB
ceZFQDUZimC9oJ0scARz3zXQu3VNzgLxup/NKWRltX6EYqJvn1S3mtJIQ/N0oWYHz5s0itTVfKJy
NnTI95hkBES/iCKUoxaC5EA2eBo5xPLuhdTwTmGb4FIitNpV42XS4okpGRBeyV6+mQnj3qamVwAW
qAjUNLTecdSq94GmN+y+5wnYnWyxwrNQSFvVGZJINclaTof7GqDXsffddzK3xYG3gd+rV40jLQLd
zw50jKdtSvb5AUEblBu5Ns3V0nLqZjDkVWpr2Ir29SSryDrMPc1B0YWvfZMVms2w40NqH/M+5KhZ
PBv0/veVBFREur7WSf4fCT8PDIy5zJ7Hc5WbJnIUJzy+V+0Q7r+QWuRK3c+cPm3cpShTacNZWvkr
9YqxP4KxSeJNgWmG1ybydXSmZ+b0/SZWxsArFiCl9rJnb8DS8zgZT3mUUuNF75TqKh5Q+d4+Menk
hZwCZgYHkd4oxvAQwwZXfJ/15lGo/UHYOTMosUwHAJuDPBKIIEB/vg2TMDyHGoZy56skQDyhsJ+n
Z7dUS/LbgWQl1gdKsV3xlqY2RjMM8SStW/FceHtFGC/XdUV2s4a7gWyr6OBwTmKpS3yj6zodgfCK
92Df/gfVTWXqqKY+lfI/cn797ZOpxBl5aD/c1C+wtSVrfi5B/cfiwmy4DQe+p8kbESaPSCiX9mJR
xGbT67xskw2eaMB1cAe1WVIYUthibo5mXylD0km/ENq2FoB1vV4y5TmHf7MKkd7bqywQ1gio9gTW
wZfSYlrqAzIkQWaP3rMuEFQuDiQPiTZlSI+WKGdRhMi/U10q5qPmkiT6MDQolppnG9g430s5VGtZ
8QIHVWJ2lAIFjEXi9+MBrCjEFXVWd5N+s8Zat2TYZ2XkPIdOc9Vyx7VGsmy2fDvJ1Gi1HKvLnLnd
rGcSwM0EEdY1IZlOUzY7AIFe2xB3bOp/VqfL/df1hKYXh3X29+b/Zf5nOJ9skuYRnelLbwLNOrMZ
e39glMmHtv0A9x1c8IvIhUd3n8ODXAkaDlIKlRkU0jDBF1sKZvC/mp5Lof4Ly63tO9KIp2o8IILR
y93JrWm7/Yp6qPWJ1007BAzzlimyuMSZtH0oK4B7XPZ8TkY2p7EWySzgubkDrMFCd2+w1iN5OYy+
A7SvvT9luqF4OwOKnk8XArH3Dnrmlq3E7Sd75zsc/ctNki6zfGHmXDzqfB7y3ZTF0l34GvTzSr+p
DN0vkQl8C5mqOMkzM2MMpmsVXwg5I+sCezhxpyIRt3Ms+5z75sfVsf6o41MnL4ihF2csGl7MvI4o
WxylOCBHZwhFbZtfmF/iLUanaPZQWQKG1ajPUkcNKyygwstqORZy86aWA59RsvI2iBzhjQWAg6wq
tb6zHPOg/Q/Ci1JLnp4uF6/UboUyMONtHrbchSuh1daY2wbTenJsnoCGV4Si+jLhCMWwSCq7H5wy
7p6AlWvzwc2pXEmcoq3qmWwdoAqth2gCxsBRarmoGHWgW5di2eqZAsOiOMKunctyoetFqUQcU1y8
bumI4YqExIwslNoJVVXEr/KHMGU2282lPeFQqCGtjc5CTe+3TRKrfpG0gY2c3Mx6ydilJZ/P87f/
KxUb5UiS6Ia/tfYRqJJhI1fZ7B18pHFgsyROjz95ZInASZaFyrxyaFapyyC2nOAQC7K98n/PDYyD
9WFLtwosz5R8/FxF/gi4CHdUYjI0W6P6DGVTVfaS2itYbCBivbQf5oF1h07gLRmPK1pOCsw1B9ma
XiL6EnPqHsQFw8EusdFDV387UslZqocQ3nDwv92g6tv0Tfg5HBSa27Uo6VvnZEFOzSUtbQ+TFXau
FMU2N9qZ1/4hCDGzb5MSPt6T0/ZHTdzjCAeFtCcxlMl0GafDuMGtsJp1RYbLwXeyTgSRl41egCEB
zilhBIW/H1Q+Z/g78EUz48UvUuI8HjqLlrRx+9rphddltsq5z+6E63G2NJX38E4s/ZxSwTWQGpRp
H5c7IO1RkYCyQ1+27DOlPlp2xjH4XPLTQMMmNmNrtsIKrw2fpgikk3lhtOfv+Csd+Z57uUMGZnH/
gEkKGuRTocq7BRgIm6+na/psouKAiRPq4VvPmB6qk2Cn7B09lhLoTi8IvaL1EAshLSK2/LpR1Hi1
O4Yj0kaMDgQBMv22HGJjihEJkEGx4vUHCwzQ0J7Q3oNpoG8zvejCoK8aeJJqlxbqTwCK3cht7Kt6
tbjiyI0Skved41L+U4OvFCyVRc10DVTCVW/PsMwVvLx4sz9/U2qHT7mCWWuitfbnS/kb5mmhXeWq
NWGPameAFv3ma9F6yQ3/FEsQSZrW9szYbWZdnTWTv5cJCGAZYEVVbZ9WWKGuA4bYe7aZasrM7+ua
2YB66MazxJ0AOj8ql50nZsAwzhJpph6L/xedEREEBQX7/4BmYrzPkapQdwlox3jiUkmDLD08gIPD
5er7BMtd2E8rl/EbvWNPzKjrDK1Y2AjY0XHiI3WVtA0dixPfS1R+FJ4Kt6Xh187ELjP4W/4aM1mx
xF5tNQTcQ9OjKgvWNN9TJY4R4iknGs+rzzX740gB7qaVaz4lp/l7Tjaw1qJlzlY+7SevEEvZiTJH
EK8g3G5vqWxbB1axXL2QdUkIy71KaH4mc8qM4CSguZFgRLbx+Sx92Dl9EPPkbS/iKOFRwxc7hhYV
+ttbJ4pUOShcM+ll1Vs6/N7Y2541JPGSmeuF409Sp8BdSTpiXnWN5R/ZyED1D20ZCUGjPjYxZAk4
9oq91wFywumF6oJa0q7B2AR0zTNIdkwmU8Wh4D/7B8YjEf73S4r7MoMjPk7M9XzG5vkXlc/aKx2k
lKY+zQrpvGOmpnsl10lgkq1pB6pOK+3j0bGrQ0sJrHReZwIRJnVLWzGNmi4jtmTg6X19/XPU9p9L
6O+bV2RND8YhoT287i7yiUp2i48vS222h6zOGXrLAcE3PshKRSJMlaU1IDARHhc9Ix3njYPeNmqk
imB2IKmv35gmC0WVu1WSJpLsZHlH1a2/jCSBOX5t3Ehy/7EO10eAXhpCOJbAfB1M8GIRjzQ82CPN
B5bjYU/ydcH+vq+fQ082MDHTnl6UbrdPw6NgSZdkSfaEO+OsWUemA+pNB9ai8xfdDxOBcywERSTI
xRhsMDdrm/nDNSo1pRtCN2ziwKjQ8qP7hhRWxEAj/XMaChLsYk/u6io0UbuMbn+wJhbYcuipQnMl
cDxGJAoB0ryARYO1TYO4Lm7DiABgWgDurwceZD96d7Pj490QilvSp2jmPTufOeTsjVMCVHsTNQ3A
sYTJgIkJzS2ymJywKyZR8cnc+TfNHpyGBNi2hPrgXVrqaQie/mHsBYxj9tBaoTDJkOd6kxZFcXQB
5Tos/CvnUpmj8x2YanXdwXH42QsL48L4nTcYRuQqPTW0hzmua3LnzXmEGaBPjhzjsJWa2/+Kic+w
h2HKYJ/f0q5+EZ3Cf/kgkHVYLmUte+DFRFvoPcpnQkV0N1qoigNE0b65lhg7DqsCUhMtWfHWe8CX
hm2+V8ab/+/VWWYtGyW2usz4q6Qxft62GQYXIiQcC7P85l3BXHRxO9+Ct/5yNyZvNe+PAiA9V1L1
UoYl5RRArSZLjbQtFnAzV1KyH0rro8px/1ikTjA1fJhe4boLZ2wXCfgQkG7r6DVggwdfY9bk8N+8
9JzIDHJUU8ak2MCQ1qVTQRUBO/Mtq/IC2PVu3gjl0WznGoExtMKHkVI2FOdGbE0wC0QJfdyXvCbj
Sey1DYAE86yy/Hgpv0qCAwI0C5P87Aha4fseBflAtuXwwGRDvtkFfUnh53WXKFaCBbQYYX1EI6xH
GTO/2m6ZMed23BxADBfVOM+P3Hk8Gne+bFUMSBUU+2AqAcOjTocigcq6vndCur75Rq26TRGCjzEf
eS4Q1WrvaWFq8qEGddQf7XZrzI4E5QzKt2bmZAljV7z6RLcxixEgRyhujTL3h1Fd2mtDwE11sssp
EFMDXJAM9ok8JPQrNei+d/f/UhHk7xAk0VlGuz9K3FockeEm48wUMMcq3fXCUj/HWPqIme50LsL6
t0oJ5m5atSqndzB/tjED5LBTKx8wizumW7rDiUUCv1sL4qaQUzrBDphYWCysh/Z8WiXjk7ZlA+tH
/cnh6IdbjJL0P1t625gFmSlIXbUG1GKjB5waii5Rj5rezeIVaLYDPigox0nOClX1FXn3vu9w3neC
fnpEhQ7D8nx8q2RD+dpuCFAqCxwomhdcnUIPguNvTXD6KNUbIMMeb0pXOr5EMqltdaLHqs2eQsgf
zfALcyPbQYSpGZ8LVTU7garoxhRsrjhO5rMWeDFfPIRAGC6JdpLAjoBRaBQm0BallZy1OJ3xV7UB
gQljJqvOwmV4LQM3aXyEZDRJNHmWp3W+PdYx9nEAPqd7YTAWPo/M5xa4bEtwJ1nIt6KhzKP/YdwI
vjCcvkB3IXIMTJqJg1LJDmQ5t6pKIyqra/kuaHdEMP0tnfzgsBRQwdfbSwFuZr4Gq/By+EVqpdEV
zZqd6arYK0U5CUX3BOIBM+iSDU3R69f5NhGn2kIV9sRqorH/yAzP84FAAbATOppBdUkR/p3nRHzg
Nz7/ZhSxU8ODRWdTxO7jwchHGbtgXKkF8D+d/8VqbQuuKUgDTuQHdAK6hWm+eafSco9BPaghpFKg
Wj9Knx6UTUsBbyTUwsfbfUXaKZeZvqeAuEmVj8+B2DxomYIdAXpCmRI17br/pNE2+HAvxUUiULVK
bucUn8b0R8hmHd7UPEMZrSfCxGIjUfgN+oWwdemcQVwK82YunTVkwnrG7xHb4yG+9YLxmhXzQxnC
ypSHWkR4ia+ThEBG898pEpPoxgfBXVDrvrRxyoFPFXnqV86q59qDeb/TRn3O0CBaNnsbr0mL86BB
boXysIA1R9LiKYNrZfMCSkeE2vxeu5ow3JiImMu7BEQPdEgIokX3M/QZ1yRAJKKRfjgYgd2g4gLJ
e/dV59woFTThPGWuKfg+6dhSy+jjd+BJjvwpu/4tTgBCp9y2T8zLVyEdpv/pnTxDrMzAhmVj/9mh
EMNcpuZSyo2wbhS9obRuzCodooGvu9YYEb97OotppS8C5mpzWwokCjVREa+8wJeVAFs7lG2/FPAY
6/fCymyhFI83DqhW5Y9JnNfFMq/fR5VqR4U62CyEa5dQB2S7T3GmWo1WSPwQUgTvcxkpvUJON/ce
eeqyXFT1clM2mn+w7D6/czEUAFYR2SjD13xRVzOQllbUjVi0tMDItfSUfsQb1xDhlZyFWlw4z4r5
l3yKbmATk3fwKut0n6s7441PpQ7egCPOzKj+8PNwnhVbqiPX0dyH5fBuJZRd/uUIfATMLzTqElo/
dggP7tan0LQZAH3ICgDp4+hUU//62ovfJ2w2pN5HU5yFlL86bo6cQauYqBrkeTRLOHB4yRXnMfan
mhy5aX47fVZI7nRxz2wcC/YDhssQ15ptpOaQ4Lyi0LLc0p6708gay3BY30Tw+e46Vnmtmq5es/lb
NzPTJKogJB5RdpdervHNhsr8VZl6FzofejBMF6YTfLJ1ETM9lLCwOLqdx0jCNzRCaENYM1zxJA39
QD1uiNpbtMCltFgJKxah+F1KYoAZJkY8XU801as2mke8jvToa7qPnZZw7WJuQqUSuh4+HzSJNV43
csUArOLDf0duBdQk7GFdQJdrmwe0jv6dOWF9Q4LBP4RMIbRZ5CktuxVwkeUa/3CHAt54cmpro6K0
H+g7AQXptYIWZDI7j0kSYovLfUWgyeJklzk0SLEJKRuSH6wliO4IiVDe34IPxHR9PC6PI9nG40BS
5oE5NPIFA4Ip658ZjU9EOaUhFXsV0eWC1WsbBRFNkDWmcc9aAmdLQu4kiHGLudeM+DOvBN8djfY/
1TWkkjpXnccQ+RUJWXmFmhgEaPkI5qP/UEnX3iv9du+cPJuCtVYStwPCxi652phQMPUasuB4bCth
slgM4qoSwuPwf/409LTro6VzI5TAJNyTYVCIP4PuQmOw+eKXYDrSh16TioG96nC6j+b/kziFX5pZ
5k0teL9i5o9h17GvyGKYGGI94ylUWQleC/GZjPGjFqC1rlbh+ID/OC0pk2v1a1H5bymTRq8owGb6
GS26kPrruQjaDC1Ia3yb5E4q/8mch99LryMeEptVgaFszjaWyDbAaNPxim0JqBmiGM4H7Y4hNBx+
ypwj/njliEhGUDsEk96ytipUa03dbyozkFmumaDPK23CddxZlI8QEFJEIz9D8P6k+qc1R+vr4g30
gY9xAaTwNB96RSDiVW9/DGR75NuAbWa4RMpdhWQXULAt6d3zUD9bqbqLCayihqjOIf+O0fLdPHZJ
zoKK1zUx6PEav1w+H9JgCZkz1SXjtLMArWyuB+6bMcjwUjAaQJysUhgoFvDzS0ULF+VvfRZ0OkAj
C2+/UGR0w31iu6j+mYPyr78j2HPeFBMKdb9IxLI/HRn4phUoy14rcEc/wiO+NNjcorDWtD0RJ9he
DJZJwdKdhbpbQNt8UylqSwh6cDpqKj33LBQv95VqcnyIPcQWvwlzYMuBbQC61N9jJN1RctwdHBq/
SsRaIZtj+dMNZjoYCi25cQbW7MNT8QiGmZVSm8pyHyfdN9L4h/ftjAj8fRzG0Kn4BXnAY5ZgSEAA
V+E2328cGfX9zr3ZZBGuEWcrrpjnoo5fvQJFfX9SyC2oMvG0IKLYr7DyX9t/FGdMFb+1jKQGNVJe
9Zz6WFARFwFQzmKarMZpq9s/4aBtK/+xgI8gp5FyRuXGmpU2Z8LSfQHuu+r8CpKrylmSz5PpEWnT
9f/Zs2h0VY8OqJqGXfWlDcWk1ohhyCkHG0nqwLPFDJ3Z3P8nsLfDU2IbYbaT7P72/8y7wKhYyHgU
TrxjVm/ogT/S2BwzwOhgijxod2oqomS7cLt7iFErfjIgM5W4x0M10e2v7bCCR7V+DlatVz5Xe5aA
A6HTJ4EfQ3qaeEAvZ0QvRH0Yq3U/iJYg+u6add5sAA4muQY7mqIjjYJs4kqM2nR6Q+v6vpd5TGQ5
0ek8srFLhUf2sF5T7UukykiBEoxN9ehpohlpQFTxkDMqu5eFPTFd2PN2WC/xkybLzdzKsQyu9E4S
cstshsXg+cPAlATso5VUKyPvHSDImmdylVHFBqKOEbvIJgC772rBVD4DkMDCSFwhWQuwZL0v4Nq9
xvg2VlS4nCbv7c8OuNMTUqCUFUtdUbyWAbG6lN926GzUNKYtIziK6ozrGbxjLhdwBFbSEFknjH5t
bAV546kAeXtarESXykV+miQGeSqsDKcze/lgrezk1Eki3ojsWwXIcQZLIpBHfsUl5T40PGlaVWZh
tD2lIpsveyzKmV2Tydfbc1N+JRLX/ZIsSZUtyuH1gbMRI7HcwmBRdx3pwzgKZxPprMKXo27VUzaD
MRSm3SIr4LgcYaaSA7jL+kZhHLvL96IdZrhWe12N3XKsyKxKvMA+yv9HKaYVD1vcwtTWdH4WGSO3
WTvnl6n0BtL7BXCbkFe2NZCuMkOXB6oNncRmxVLRlDXHKoHIP1ujwGa/5bksWQpT7grk27bC47G8
NCcrfOntJ8g0cJS98zV6cwdhXe/9mF2XBT7Z93bWnxCdz6Xq/YvvDPKmC0S0advIfocYut5LHNns
BohJnCb7m911yZzhTOH06BIUvh1C760hMUB3De1rtuCb4h+MxuBZNDuWikdj0ohX1Je84nKyQRsp
5x4cYFaVenV3dVR1rNyjcYMeGlwBXQdWA2zOrF7aI1VMY68Jm7V+0ypFaHS5CHQOlnmV/IxGg8Lz
e1+llapiB7V7BNxjB043loEalQStQ44WPXKz5fiTG/6NWBUw7HFT+DjEccNLx7cucLVHsv60+3Lx
3mBzLr+9KCbUsmKb5vwsVd2qRWdx5qdRsl4XSgxgVJ7x24UW4IQe4YlOCvLtM/UqTdW4T59Qrsrb
/gNW7M9iMfmiNB+7HhVn3ySL71B+Nhc4sTMv3nE2Xd1QfbZmvPuwwd8cBecTmKHY5d1WfZvcbRal
kYdJWRRWpcbLvIgKdrUTRVgqidfyt+F5uRE78FqV/3URmItdPoztQRXBd8KiiovDgbyDnNMwKAhC
Xv0qxHbFFy+K7xiiox3VMnpOzy2M9IRzc1wH+zsjXNG81e4vqblMUpM5l92xsxorOpW9wEjIYrVx
y1QJhSZhE5Dd9s0tSpG3N7MOhP8rcf5BCl3QxL50MOWsTDHv2uy7EX/pXpgWCbruGWbF6shvzySF
T9QeM0nn62lWfVvGJxIu0lSmCbQJfxyS3IKUBDd0MZgisyfqBhEs6vu3AEEK/vsqeCsqwWzY6T3Q
pJwC9qzxuLET+B3SmTWoUivwB36vzwNoMnRsjipr0y1yrRhnSUQHk3q0lJfQ1NwjP8SUnB+NhWDt
TCU0NCfiuZZBCPc1GkvuCqrB0m3OhsiJTPxSNcT2aU6zpdnDQYFH/X1xWiXFR7kw6pLb/IaGBV+w
h3cCUk7PF24kcuWOeKhyywtkac+Mynkg86afjudPEH2r01DRU70QoxKzMW7u3LJPNnsDXOvN+YvJ
l+Fj3/HTcHXCGHTomvKwiWL9IChEgeg3sPHYGVjnGjhbJQXurwyoLNeIVlPL6PcPNZDL7NV+r8XY
X+JTd61340iPzCn5gcpfYzD2rmT49hOJwNRDHKCfPcnEukQu9WDHEi8UGLUShMFVxOG1zs6Ewuj9
izWGbj8oT/QRQDHJONH02236taUxzxJtChL4mJy7itbt34/EOOLDvVcH1+rkMnYQ1O2eCpISsy02
HhwewGLU0JEdNqpUPoLE3vYvGqOSe21L4Vyk6tEkDftZKOmSFSEH6DJ/k2rmEa3cEPc79DGRgQ7a
nyklaJa4Jij1RVBnAOTRQzs/nvUZLAwkfcVBsXzw7InZPCCdz5G/sN4uS35XkXd5d7S3l2S4oJZM
3njkGvafRZU5FAe0tKQzS6PyDr+SUkNFFbbZyVuOys9wyduV4Kfh4qe6ZJH1X0JgX9ADwF+JwNWl
8eNqcpimMeh8IDwEsO9Otmv/1fBOUEN087uzxLsm//4TQmb4yFrE6PB1p8HubFfSxkHKgDYX3az0
kRco+7jdeJ+A5KFp0m6sOQMPIqzd1BYOBLEsL6XsbrmE2m45Hgjc7xWM0dVDgjtR0BsisS0Y9JnV
+8ZXxMh6hYvJZmdIiFh7THxq1nTPDKbyzUNMpNo0lhICvxPcNuKbYj+ChnFbfsRpwU29RP1WLEjq
HkT6X0rUcy8SFYuRMjsRnema0HOpMyouW/kDmQ48VCX6eZ4sDE5Zy7jgcAFfellOlaNHlNEWaNpT
pVFSdP/NyU2Qc2wLCOPFTOn6A/C6KjzQhcYp7hNuftnS6lSzES9kqv8YOxqujpjkyCubbE/lXR1K
0wOLNCftcHuUaE/S5mwnAY5Mc3IbwuyhkTtBWJtyU5L36CEzjcLRJcFybk+FFhd6eEq+R2H89fYW
KfuLceU50G7wBrxtxLSH+kExiGLfQXj4AVKJA2hBPED0nZKTJTevMw5sg5oWAme/QI1756sF614b
sJ4+oIvhAfpBkHnUma0WzVPCXrxRHetyTIR+bMTwueJPs0Z05ypgiLA5dilfKqsg/F5H40thG/BV
S6vUsZUerJkJMSH4luGzZyJMh3ncR0jjO5J88U3LjY8ABJzCBe3Bu9PWQYHvKKLllbQuxBJ2W9pr
hayKfJTfpEbefyq/NV+vpMc8E4xwN4YPgz0rxDLdktPNOBChCBGvSPeakdkAcgGRz2+5f2ng+BSS
FWLZ0fZXQd3WtHbch2lAQ6QaLvTl95B/IZI968Bq3kKXGb8v8gH/5Q+1LmqhS4fyPvXRhIJC6nnp
u7SkE+C5uNOiJMCrGiWcLJSdkt0OWoF6PpP58WYS5udj7P2uZpPbEpn7RHEjzbcBlEbH1GduBqo1
s0A0ESIkRKk1yEtjHgohmEpkuRyzsRjbNlJaMvMUQj4Rqo3C+1/6K6h0/jmbAgxalecZ2Fhz1iYD
6lhjOrz4t8TZRJqMMJJDJ6IxweKtgPbUnvPJpLLtgYiNbRG8zNo+zAv22zGR1wuNuoXX6HMrll6J
tZdZs5QcBOZOxFeO4lIxgPvecHw7680w2Tu/z54ZEdzCezdYQKALj5jcsK20XjT34i0cGUdTzjkw
GnJFsLmMuzstpCG1kKmA99WtcAxTyVx9Ifq68LzwGwMY2D94MKQk8wqYul696ZGyRTzmhyUXAojo
tNdv6daTfZoPI8rCZkbqzjsuP8eaDCBfYR/ARBOnf027HpG6qyWtOrtkTH1kYIkuqneqHgr8cMn7
t/FuUqH27FgAP9/TRNbDYiIfIG5kvhQ4FmGjyD7ccMk8Xh/VUo/9vmM97mtdf9S6SF3th8aeuXsp
Bltlq7ScLv7Q1y8ffhFex5/9PXPLMh1GtkcqY2ZBkK82xfUeodCWh26SvAHs0dOZdDomC3zSeidQ
9x0yh8p6viMJoSeYnZ91lcLprNTaplOtma95wiota86AuQ80UvvrATyImyKGPKwuYI34S+9FbpJL
lquWip1MR4pcWcE3bLJ3/PcPC1fQKSgy0yDQs7PnQ7WlIDXpUihBzGbljHe+ARfMc4APqoQrg1QK
KGnkI8CQuFyR6FzMw07PsTgxIi0od7uGB9AZkGf5JR0EirzXP7oL+mc4c4mqvdJQUid1cMAvrH3I
zdRJkoXUbVsQCSoxzNmXz7TgDE5/KeX79T2/r+V49pWUqu4yeq8P+2phicqnDd0Pvc9CeENekt/R
si1DEIAyq42MhwdPHbzzVIEwBmD6Bc7e5mymtrAt4FNzFfZNmwnQuB6sd51pkhEqbnG3HKgsD/90
B4ef0IRprYGBZ3Uno918rarIH4wMinpNdDayPDqfB51bpxuJFJGkM9IcocsOvZZlitUHuYgNhe5P
xyBjxNKEiCCSHpKkqz5HNVMZ3DCbmakJYRSosuoLBbkpNSNsVEhdIHeXI7Gk+Wkk1D2yg+W8RCdh
j9491KxzqGUFmuQEewxiVoaP5j4hBqnvMPtDVnjmW/alwQrG3AuSVkE+5V/2pUUdW8hNviQ4DJWO
JOMoPOXUsuiYoYvNds1ADS61i8xhx0Sa+FG/qrM7G7Nqnea4oBQ4dtLVffBdt6rK/trthuGQCe2C
+2IQ+3bHvnBEc9RBG3Y4nG0E+0Ph18CuY+lQ92qW8AwIx6uvCiRbIwKAMXbZv+EAGPTCBYCfGaif
a8V9GCn4bd4bfpJay3b24gr8aFkrAA3VBd72WVUg6RDnDyL+ToC8JygPF17ci5kbnX5Bav7DUmaV
nw6BcxNgIEC9BDhK9IBa2/W5zG09O3A175loa8iASAMDbu8557EAUHMWJq6diLbd4pGv7VIG6yXK
jrfxu1T4Q8RFjzOIHOhkXsj+IBcjuDPX8/z5J2u+FZjgkT87bzo+JHuinHKfC7fMzcu139A54GEV
HkpWQiZMrW/GYCfdSMCouL5BCkvtMkPA0UlfxsJvz2dj/s9A93C0Go4jlZgtpXOEh+7lMkm5mVU6
Z+twrrYigxixCcFwmW2FQQS1Bxx5SYO/IWApN6eZk3Aw8bSv5uO6l9kFI58G4NfBHS7L4HQE90YD
LywqdBY4loLvc414fhGbXVE0sjE1tHTrsZJ8aJSBKBfhUQxAJNOLmDxORMTZg1FlCRVxNTgxBXKh
yR7pieRSed8iW+22874sLOtc1Evtbuimay11Wyol6kZuZr1d1OflGZ/pNnkLMVapL4m5QdvjNwUj
IKnYMgfBiLSYxk8csYN97jM01hw/IDDobOVi6Aw2BaJN+x7VZrhmJB5Ixhb5UAEdaBx3miGZW8Ga
n0uBR9POHWFKUjhLN1VcCZHP6yRPJczmFwqFkrKOX+HMy6ZNdfL1n4hG/meRmzxIrWWUInIG56Oy
VnyZpeFucRdMlBsIuk16CFAnTCCYSxSn4Yq4RL64G38ibce62xNuqfu3jP7M+TjwvenA4g+gcMOv
Y+vRUo9TDE25WeS0m17iPWTXH6ekgHIIeTiU61Tdkv2ZITecx3PIb4WLN/hnsKcjlBwAVzP1jiil
mhfJf0QJ1XDzOpTKM2Oyascsd+waWR0cZXVB+VJN8OeD7Qvpp1eu1kqphXllQigfzLMchZK8ZT+/
+1jJUhm4g0xgzxDDmtMDu/ufF/e8jM1wRgQtMkDUN8Y+zD7tZOZuWoD9Sf8tJ/GWuKDLlXv1k01h
2T/i6quV7PzNyRYMJSYC/JwnTMa8XWC5If2j6V5QrM0VD/TvToL/114YNshPlQT1nEKL6DczaeDB
QVzePdrrNA0XGl5YdVB9CsdDUSjVs4ZVquk7FQNiaZHOKGhqGKq/nkLlDEhN3PWksveWZs8QWEty
hE0r3k/d7ZO51su0HSWYkS3gq6AtBcMy25U/qMwM0Hk4gawiXcuV24jzqQnT2AEy7qOhFVhM0+q8
RxHyI7Sdrp9ETXzqdQz0MuBjiKkIcNzKdfzlzrlCtyrpJSTNIXOr5zevnhKEI+u3ORzi7J4ENj3E
ztpT7Mmuvk6FwKzwjmbPx1jkOVjRKUwNbqqEsZAQ2KmVJSYG9v5WQkQKwiXqafCz4blz7pTluCT7
jWjZxvXtjjt09uSYpaesghYcp08iShU5+hytPNmxovtg1vJ45zbShsEfKuQP+qlFHoKPQdsGGCA6
8Yjte+o244/ZJ/igt23y+aaXvcSCnEJBozqfu4vmZMHH8yyWAOWqttvLiH5IEWcl2ZtUCtFsKn2J
R2ra0FLqFdbMe+8DUMGT2bX5b93wWINL5rSRUgN00Dmg2M269h/TRriY+mitUBJJpjNMeUlspins
/lhOC1YOoYWVQ+CjI9iOt0x/KqfNOJl+rYd4QYhuq1BnCfTzoKwOmVuClGm4L6pd50LL7Y+hNt3o
UqBj9xZcElDxJXua1A9H8GWGYfGzHe2Bg2QFkO/7LxWz+RWWL5mPWF/lJE6HvpkmjxI1NaM/LMJC
2wSg6J+i6UwqCRND0Ac0wk1vYtiuBSEQZJSslMpliq8s3m345ud/a9LR9BfOJgaPg3rSQyaRK5cC
eTxQSSU9Nd7x/DbA+PETWY1ctNap8t5uluN4pPqUiKbI3WygiczY5TeINt07eb62kPtWcrVvJSu+
G3KTRONwr/IMP1Tyef0dw6JHRDiPUYqeqJxCUrA4r9xrNx57FZPWOhxynX3PpTP9rdg6WawbhXNu
6AdJnzNtTuyYlRDRks/J4HHLaviXDYyXqk+5e5BVsAW9gskojnyibW3DP1dl94dT9jA+A8A6HhYM
r7d+glihpqPzvCyeuRQ7BGhqTXLsAaLy8RkTMOFcLSRPhLN4e0QqbTY6ddlfodDgflep8I22qCXn
fHEDXqgC9gwxrxQWaQvWkhxFFTbpT5yRPkyBRz+InV5gBU+tKwMsku+6KEjrJFQSDTeBLs3R2uip
q6WP0ayXnjQE4IA4Sl14G4BE6aI34R/oKN5Q+iTSF6qTlWVSKc2YjLQ6ZLjIB/ONB5M7+LTxzIQj
m+xJZYdUw1CJ7khy5X+2EJXMOf4jkDqGzmdmVnCkrzbwmbsOIM5Yed3rwcB/SuqzK31/1Ekx3r9H
wJhE97otIHGRwq/6DKeB3ANjF260emKad/JSLo2WDoEnLmUqbV9Vu5orAGEbRqpsyZokgK+PGGQJ
eK+DcFKTFP87oQjBRu8cikz3wR1j2G4vKgImhpe9U/0KaaeE014XjKxo8dvV9EmNmzcOL3penNOj
bZXepmz+1luOgjgRDKKFghlRijhrJooC4t4rN7K98sjqtPdgW1Pj/3ZijTjLnC9lBTCs5WfjUMr/
YcK/qMWOJssiiSTi1E/YBUJuA25XFz+8MEHCVr1YJu9BjiTp9iShLKakN6NAcgsdhC1g9I/knREN
g2KVaXAsU4MaO6kDc4hLOP1pQSsMZ8kqIDwB1GJQlgd6Pl2+s8iJsCXxu3H/Bc7qQzK01S7j4CcE
En3JKHqqWR4VKbU4GoeY911cLJMmTgCl5LyOfukBq8+nKzagQAqIPE1g2cfcoAT40I0gmIj2JuPo
zsoYnHjidio5Hgc/hNjpg+/51/wU3LbaW/kAO0eWTIeB4fI8LIkWx1ikwPx73S9ihCuT1w9UvF+T
eH3D8uBSjfTr4tU8857q46EfjjEF1tl4gQ3BPgli3PxJ4LNxzfVZesUQtG3TNSfYpyrtPCRWxTsF
eacg5klSqaEfiduQweLwZBPdZ+Ohkzr05peZz4+/gs1PxxYD38CBKwgLtRi5ayZ1dp4u3bbBxZGS
W0JQtIf00ndpXRowdN5v/thuKh4CU1M7eKs4KHQCqJRu4FasN7rqjCcl1gWzr/xPJxNh9JVn8Rie
sP5d/RtmWakoPyGegvUyz1CjvA6fOvuqZlj8zT8Ei/P1jD+I2UNkR6ok5VIAXiWdox+Bkvu77jRu
swbJZGfGBETrZD0M6DXjOcRZxUD5gQ6Lh0E/Nk8+dxW5A++PxWEz7dt6mHqkrknck07++fztj3i2
XCkDi+vfBje0VMZYr+qtkevFSyXHUt0CxmQEhYX1uILD93KsQoPrvN8XFjXsTvrhEUX3Wzqi2TFL
RU7VeqXJXtIwcjo03FVxK1L49gXVH91fW4aw2IMoejwrlLjyG0Od83ZzfD3fMCOlSmXa3ylGxXzO
VoCyCvFjyKNJxj6ZOkyfGFKL2MmMmN7OLzpHX86GgrBe/xuf96zdzSsXKLrrXK4AnK+su3uZCEMm
bgvbyTESqNRVD17ETHKvHfmBDX1T5eQPV7fbQegRBapRaHPwoh1kv+qJfLe45Mdtlp8YMjXLb8Ki
+bUeZoRrk3KP1RKVt+1HtH6WuqqyIkglE6wrwWZLBt+ITCwfC+NTVWdaMfzqaOkBzx4LR1B0hGe5
81YqkEQcNIBSCqsSZ+AdxTvHuVMoYOjmM8K2SFhZ2Beodk7nV1FjJ7yn/tu9slsa1S8LU7F+XwTl
JphfgmFDf+7BPi6Z8+TQDt+aZmjYuDbKe2BtLeOSMlymDY+BQq+9L66s9qnlszt6jtzbtufQrqaO
YkLKetpW3LSBWQE/PsawR1b0kBs4XlBkd2use5JYBfjnF1vI7Sy3ygjZEckrsFUfzwq/t0PEOeuV
z9+9VAxFhO8swwH5GCXdRVmn3FiSJZN/W3fpNKozkjRdQe4XZGlcYQI2avmVuOxQfLvpvwcXKajf
+B9iwp9S7JQ7Lz1t69sFxehAtOj1q1k8ZVUn69BneICCUtRbIYOHxtqAjzOce77YyeRlnkxOHux+
F7Uw5dBkV2buJVtnY9EVpSZKBVVJi6vdVbHhZ349BV8zKUlklD+8JgQhuQEODkTLK3jjUdqw+g5O
t7LnBvcNqriY0GWPBOTapKg/v/N1VidQTHA8yyOMHihB0JNLfWI2BkhAZiD/lkdit7pVZ7yiRZdN
Y8cqXLb+/6awtxLta4iN040JECC2F6eyxTzINSgRGtpnm7cb/1GWv08lGh/lL1jRBicggpk2R6Fr
A8HhG42GEUTh9ndBm5bx30Vow/kWQNz97d+9bvAkSClF2I5Hd2YfFSobyzQXqbPLQmNotnZowljk
jf9X7gbM7YQEJToo5+Ls+iGUPBZi9LvxbgslCW2TUM5H02BZlNb92Qj5cC3pdn+19+iKv3JmSzml
bPkvB4ScQo3UwKZD+6zon3+1JVqAA+yPKjaCwPKIN8WXwXWmGmAaw3ltKnoHrDNbDbItf867odRK
3d9Bgh1X1li+mQxF2D/ClE45LsbSBCO87qFIaEfeV/yYNbHGpBwkhSKq9F4FmBM0hK9t9lW7mhtA
fNFQLTFRdiUgbFHxxbe76Y3kHlm92BEEcp1h5RuQyjdo+udLuz0LCW1phfcsuESd4AIWr52TaGq0
AJKRJrsnyLIu5sqLrd9T/KlBmlxH9crt600RaN6ZLLdFwKXMWGr6lwJIaSD5qELj6VVNfhuzgOdU
RZVE5rIPmQ2fF8nRSJqEtBE+6F3E9XrHx4VzOvBmmFLezdXm00WDWGqiV4A/gzBBithBvNQO66XL
rWYK71+XkZsnsxKxWBa5HvMGYiAH3beVxP9sQIAkqWvX+br1vOmUBYrFNytvxE6BuUulzaTnsVQN
GbMgo02rKGzslWxBOH5TojlOYuBdFjG8KiKwSWaifb/bbR8Ug0vqV7zv8uIgJAzuueKVdmyrst4l
R99MSfuNs9BJcuZR6AsHruAkrBSGgBAxmsGHaqxB6uYyPYqzOX6hOOYz4/FkPte5uabUYWk9HvIb
KFv5UfiektB7UGPHU4T+BgyJMgpM81CHKDLnJuWpT0OtKoc0EoKydS8Wjp15tNpfafQVToxOw332
0CsZW9kEjDvjNkyTULSI/oxv7OLrv7x4CUMqmGn5EAYOmD1R2X6jEb9fBfM8yddMVWy3773RmXYh
9ldz7fS1LoLpzTwJeKlSHVXQ+wg3dfQP+ch0CoBmzMpTJQBe3qXKWROrL38fp3wclxc6Kml51Brj
XMzf6zPw3H2f1h0Vuo8p0AesvST1un2KwXxPtmbOrEx4pmgRBi8+3Pevql8GARijcRFKVw4QvpZd
pNWmxcv59hdHy1RB81ikhHKSIvmfi7D1sKCta7yW5ZNHEyLu3JrRJlMqiexvPlMD6WTQU1RnoNfd
nfDjJlEw5Cmua8AtHQJtyjkLKg4c85ZaJCWqdAIntv540ruFUdv6m3efCiS0crZpxs8bjRIUQ+cl
CToevNCMrD64RX9MCsnjivAaifVeirdI6b098/BB105v1g/J+XtaOC0OKd6Mt9vm3qAiqUTEG7rM
0ovN/8EV83zSnYb6YkdbYpDsIdGtx1JSP55DRy2Bdgk4FDe08rePbp8Vrw8Kw85TO5iSzng5gg0o
2nrEbI3vTTd/pCg+tLE9Xzi+bL6uRuqrVNqSaWA2LrCb/WIbPYbuZzxUC+nEnV3f2vfrgssPvxRB
xmgR43c6csgEf4bAvHme00+B7rqOHbufwXGZ9KdlWZ5rCag565ZZBskr1BxsCcyjlund/TidpRb9
D6N6fFWzqkhZY8EcMCw1XJvgcZy8CfQh5A8UurpdUQ/xegCGmOnqPNvh6Q7+xPIDRuAZ146RpR4Q
Z1vo8KcEtSzslpZR42C4wzI75r97O24+FTgsSAwpztlU17zWFQiBskbVOw+X57tQhFr/jYqMDTPD
MfEh90IkdaZqBHSDVQ+1EYmVX7Kz/6q5lTL9q1PpXQ19JL3e/qnmecxehFyCYGKALUKVyqOnE1KI
eRXSKTcgSsvrjn/5f05Q5TuFRl9yk55U09fOuDmYvyl0x4Ey8rxN09ZKEsQItZAXsgkkr+osG45/
mWI7u9yUjAFkRx6P7rx4dZwVOYPWZ3swD/SAOtxwn310AU7GBRNM+hFGb9mpyZGiiZN+HBKhFl1S
VxBcQLWyF3BykpUlWhfW2DrpUmPLVYSScKlb9zcZvV4TXtGQ3LI2bmr6jHqtwfcTlL9OvpEY0k6Z
5nBLmF/dDAqyn2Xp5qtdhQLC0s25prNFVFtqfsX534UuQNQ2M3a0eVA+HqynossW9DB55+qjJsTe
1xlHajye4EeRLJApN9gIRkNiozh6kgf8aZixr57MUbB4UICDg08K3Tu9Kqv2jFFFeBo9xkknanF7
AlmoODHV5Zz1B3/WKHSin4XyLdECGuWYs9z8Fl9SLB+CKKXjkY7VxgBF51aDCykldlm7I9Xo2B/K
mpUmL7tiv3G1RK6mxSDLyilF/UelTe0gfUdjfibR6wdkvccneDZt1aO7nnoSsG8LFZe89wr6mcxb
eCr3N7v4VHrdDIdEzc9Nc5wxo4lqfnRjhkoPzqAEtr56YUsBpThhb6pJbcIxsVqsTesLwejJBnvz
tj8m0VKpMEc7ubeJnX9HYkG3VxCEokuhUCVs4bSUsiXyoP2sMunVBwXcRHKbwzbG0hdesCn6+BuR
qQILM/A8+PqJnl4RWmOpOupg3SN0m/bO7u6p9G+GBdGy4FHiqFhGc01ckrZ7GK6OgVi0+6qRBpAQ
oZAmz6lC/nHsSG9ioHKaPOvmS0zPWb0Co/ivJPRi4VgLtIJoHGwB7cjTeyrxTyVCHix2Xyn88tBj
L4nz6fp/TQnER4nSWJt2RMWGY8fPOjXfPquy5iuzL9JW3BGFXcbpPzcTqmqmwuzZaer4aW5BMwqb
FDyzn4oQxb3qsriPuFpfS3AjIZbjJmcXX1uK15hNF2nzOHnBiAP5Bo1DqeaKG6LMth2DI6Lux/H+
eU8fK7bmpj1LDkM3715bnfWjgL7ybWloA63z5K9GbtUljno7Tl9bLIN5qKLfOw/tGIUn3AYHkeT/
83AbsHk70R5dUFFqggz5gBP95/ynuJJd3n4aFfav81RW0DSV37Luv2X5LfrZ/boTP1teFmeombdW
CpxqU/rizyk2AlVrdWxVgvbRCengeDtNXVTI7wLlgsXOkQGIpTbBpqzhHbQeFEFPY2JgBKBl5HfS
rFI5xu1p5gLuHDwqH4es+eQ+Qf3B+cqxH2l9k807WJoRm2fgxMKYcbiKTJHdJ546+hm1kQ6qRwdW
apzCAB+oWPw56RvZLxJKLZgZih2FCBIOSbWGsdj7QT4w9D0GLCF+mdOVyqdS7kW/A34ZvDOxgpKJ
act2Q0UO9JWGe3tK0BPTSUE+uly0uCHatAfmeGL90FkxfVBog2HlOZYVr7jnUYpHOKTeDAGQLskW
VMmsIFnZH56glz04UVuzCoKaNRCmFbXTs0LbNcSwKKrir/orDePnsw5UB/b5pPwosbv1e7vUcZYX
dcpzSFpscsxte6sDtm5JIdNDVmwxVUAWuNMEn3j7nDNyMSOFjRWGaWgwVHbaqO4cdTk4DQR+RQ/u
CiqKyWS++9sZosO/byt+mzjxNKzMi9fhwTZeVE7DQMssbK9OAt400tH9T1sFovqXnEvHyG14vRJr
Dq7i+wXwmNXGVBG2N2cTBPZDKH9HsecAVwHvRn61UBdkFxuMkBjzRD/ezdEAXFaL9zVI9SXDO7/C
/W8KxWEf290ZI5anXUp7Cd3rk0TCh7QHfGKoUfKi9+Hh+mNxV2jvcN4qY7DmqOWh3UbF/iF0zDZZ
ExjWq1s7fAM4oFztXZ4rqTKadfLLwagfCuCW2d4Sc0C60vgujbzcTH2RJwOkeMCrBsmmvGtY5pb7
uGWzreTuxJsjLRZCXA99ICDFCzG9rcCaKi7vX5w0G9VjC1B4/e2FWbLLWJTAeLkRdbeJ98PNsbJB
lUog0u7UiL/WPXPjonLnrbhoudY7G3OImBgtNgZiXj2OmioNQP+E6XXkcUuCYu16Ujftyee61Ls+
BPDHyzBD4Ye0xjVV85GO5x1r/p0PyVwVXXk7mbVpbIRJg8dgo3L1M8wsw6WulLu1ijNxUGlrMtAF
OI11tBQq/k4ebPjOsxvipC+Zbr0NnQ7H8Ohlh+BZfo1cBOM6M0JBEwTruGOxpZDedhbji0WX+AAg
Xnztvw1j4Jd4Jx66CXJIIGEhNJQaIfLmSLnmWrusIIqxnA10CiIMymzQriB03dHsw1v4XMc7krZA
xBD06htS2acRGSIrxrLax7WbBqVHyeGE+AlrOWX0eErNRjRHU+3x0Qp+cbeHvePopmxQ8plTqJwW
8APzmBo8xyu6kFdl25nL4zdCccxp2CKdHsy/Nl7qlo6bsApkIXI2RGDbkGyFK40SOuszgq0RkC9j
ny3tPcx9GFTaCTBHkmsSwVPRNkawHVRQ4HcmmTxAzYeyDCpTCwhfZGwm7ZOhLb1sU3yEmoRaAUOM
EI+T/RWk0wEp37vmdHX0mo1UT34dByvZKduzqJQK01f7hLUGSEaaaQ/kBGLhubm3RyPuyIpf8K0h
4l/CU0MfhnaNiS7DHdfSEnJ/IciQbKtsXQ+odEQEwidHwBB2/Cn5jfEmJRAcMdbHMcFm8PZ8WciN
ufyFislohblbWq9PjSkg3o4ufi7ABRF7pv0J9oV2v9YGu/6tS1iELE58qvaj3+A1DSBwTsrXrgxz
3aNt0zNSOd/3kD38eZKYuPxrKb52mHWXrbRtauURpLgyMPBhSxMsfkzFCTIGh6i6qu9k7Y180Cmy
1f++N3Xj90MDLqEPTX1DYAGJqEiwekyiyNEf04304w/R2H1zDdWrIRUJsTIV7tNcGrPk5ilhXWVV
FWFxEwGnLV5sfZXSEF6vAKpiTODqlHFOV5F/UOrnq/QwJvflfZlXVrN3QqiQpU6GipJZzsQiEMLf
Z3uBGZi8JDDdNSJvYyVrByJ50et5L991Ou91Xkalc+f00zEK7LryOXLQE7KxzhtlFBIpbZQjV5wg
el4/vHXjOGri5ZcCodJUmdSgDS36PuqEUt2IP8Am8iMUWJ+AX6CSUhRrOroZzaDDGdxPSGY+Xn7s
kEs0Vr15KoaeZp097kKRz3PltJDhH01x3tcLxKvYukrnxJ0hJYb9YW5slhph2QkVjDYN2GJ57H2G
tQ5DbiqUvVc6PTXmTaMMqTx6FbQnvov/20ag7/rcaKwS2xE+0+lWDh2lxYf5F4QmKiSd/WYkYeSK
Gd4+luaclcVmifO7EzqnKpiTw92byCUtgwqA7RoAwgTr5X2gDRxV/5CLv1iw6GAFOR+xIJAfbqTW
AjUU57Prb0ssdmuItKz8A/tvs6nMTgkbGq4upS7gjz2zviAZXwGYNj/v97QwM6GTa+InTZkV4qLG
L/0GtteSRbjrsgVzESrSDUBZg5nXEX2p6C7ZghYIs93UyvsMvKvvnqcStw5H4t0x2xpTRnTSzdHP
zhoiyiL+b0obG3O0MPkdGzi2iAnE13seLGv5CrxPhO1lyVfZL8nh0ReIiG0WjWJeZIfkrovo1dQK
5MwUyQc72RybVjbXAmJT3E+d4Z/bJf+KpvMT520PbnTEowihl7xkWxtmz5UMEcmiRjHs6CN6jeVp
lNFsKwNsWfmDw/lxd2wV2Hn4snu0gWoIvdB920wcfuZCRYh/YHc3u4GsZ1oXLrG+ustGAeOwpm1v
S7nZaB38ItCtzCtnPRaNVb5w0fcmzeqeoLhzWdrA76xcb8HliZZfH2eKabD/MgI1J2xegrg/zwDw
ZXXIsBJfYx+YOXIuowZXhS5GrPV9NPMuY/2U7/gWGbk9zn2gqjdmAA7rl6ZSJm77uiEMIvGxwDVh
umyRipipesNavSqOfMaAObGFiSNApM1gzpX8HFzdKISEBUYwkID7jn8w8o55euqOX+8H20Tks2sM
zkfCRaS9EZENhOwBZjHWm2LyzTMsC8U5O3OoJoO35aBktUf92ZJH/maIyfLZuxo7hQuoUPqd0TGe
0TETtAm2M5AYh8A9lA83pV60sn/UdDNczuMVl/DspsswFIoUOtmZDnfGEYNokY2tXnrGBcRdwfKU
xifyWQnzk1N6XrGVNjJJd9+SdephjB7BmSSUyCwigAH1uhdxl2KXp59ePrfxjrw7m+puhv+3Mtk/
O5yu3yw4QBLu2ypGVSWOB414kDn9X+F1rebSmw2aj6mxKK+2CAY/qjjU88/czR++SfwyjLWhZ+XC
Jymn/w0JzMdEiIZQ9HiGbHC9ZfAmzzdakmLOBU25ssg+HiymmaaU67iOwqFYBL/nPAstNqd3IN/x
KAmzSMHaRuz+Yd+RG2sCEUQrabWPO5g/bHRqrlrVM0R0LmaWlZzwlXZBl7WSYMgCjRgLlNxPweTJ
DVTRnC8scOhRYubxWpu1ppyuGfLDImdyWyhymjyfSpPGDnud0p1J2nuy+B3emgl76vKZlIOl91u3
ASBCwqx32l8+RKF/fSmFaBdXp/nRFh4l0bpQ+W35gLoH+sOKrRb06xzRvdKoYHnhrqHe52RgO1Op
d0cXDmMQfAhj0QxNZEvsI2j2/6dp8JRYC0HGRvQAUjdDj9XNXDrRXvfBuPzyS5XE0bfrZjO5YIKH
FSaUu7tIv5aSWay9+cDav1yst3a7pLG4ZNsitgmKN5dKZwxNrsGZI8IflxKL1RQtl0TwDXSQtObE
7QmcTtU/Vf0QtYnux2wmiyheeEAw5ESLfgUummeN+R/YvW03gF5z0AWCeERYLVavoEKp3YZqBzoD
Z12EDKY+55LBHY04sSpuoKF+ZLDNey4U5B6N+bFgyhktgOSZzwXj2itWrbRf6QooutoIB5ppGENh
npg+ch9zbt+YNBWVLU4KXSnHu+C7xKEJldFQdvB5EUdFDqswzf6U758m9iGlKT+G8t3Dtne6iPn5
/Q0zVFComi/MYS3YmX9k8HAdGyvx2F8nLBAwSX+gD8iFEYjqu6cVwCv6SJ39apJ5yDfz6JMbmWb6
PCLwGDKFk7NYwnDc06IISA85dFDszXwNb38g2F+nHHqBSLV8iv7VBfQ/O+Y9gKmxJPcUi4rMRlgY
B3RUO4D0PtRZXhoZx1+DTc2IMjHbq81DMYULVq/m5hSYrdh9CriCvmQ4qYZ0XU2271c26BgeAUUQ
zBmwPQrexEbgYp6Q4L8vPWHYKq6Rv0mr3CAwxqOx9mwZPU9iuhiLbulkekGZu6SiKLCQBZMUhoqj
B4f57WF0cUM0KTE8OXz29BvVtu/lL5NGDNnkpemDRj+SqNAWkyxnAYla4ojYYM3aBAeh+K8HIrnS
g9G9se2n8ec2zKx1wBTyQRPE3cvWA+lVzJxic33Qo+KEqUanaJ0TBim/uC2aCuJ7shDDdufGNJM4
pZKyehutiC87fTXM2XtSQH8HyFtGDrsbdGv8/Pp0wQAVZs2uY5zbOmxyRDOMLTXKiwMjbocM5kQt
faA/0p5Ke88cC3fU9p1hHxxTTzU8ZlJr+PrKhgnWjq58U1ucfJox7P6Scp5u1pCvu1khVjHHdDQr
FthsPBwUzfaQAzdFVl+tUJMFEPGeQdWBoWNrw/jsp4BM0gt1PQbg5PTcbUhF2j5cNQd8Wo69q5n0
M/xMk1628fv0MEhidQVh3C5fuHIC9NS81d8E0V5oyhKuh0s9D+48BWSazSbvyjhRjaD+e2po66PD
0KrH+FUSeK26i5dcxK1n/oOvsm51JrnS7O3vxXNi/E6eVKlyWVbwhG0FB7pK3VUAOXgFzgzm9qYE
lwAgAp7vtV80a+SSqQiaeohV7n9N1WbCteD1yGZpqORo3B1EUyIYwIa2RhqQav1jNTSZdCk4HOeV
BO/wKedG5bX5o8PHrrIR8RwuTn4/PtDxu+xU3CT5UNfSvQG0esYcAhwswZ29Cql/7OsH0dnE8b80
WS+zibxBpX+LnsZ/24/2FLJ71H10mezEH1BlFPXYh/xQCDMfqZrTjQ4bDrWE4Aq1Hh/wBg4xFI0s
RwykvaaWDJUNWnbWAxO6x/wSyF5du/hwSIsj2NNA31XzEqQB0cePEcvEKdqkkSuYbaR7b1XRfuZv
29u4AtwBEGQp9j7SAVriZFScde1lxvRx2rRb5FrMQ9HP0hNBiCfWAbcwZjCEa49BFmgvQTllG8rL
XlnkvY9rCOQPGwnai2y6eEkt0hv5K+oP+o3EkJHwv3xdOH/HzTMVjP52OQJAHlkt925iuXAH2WsC
mOMvepNSQkvfc4wsMkNOJeTklg8pzYSNIaaSi1ZCtHOeJm5eV1smkqeKDUQwQDZWyAfXF/y9pJEs
DyPX+Sp9A4cs8jU/tUKQiU2vMiS5C0jkD18sYlSScL9n2QmpVN5tfxMtC7uLJbDkryLkKawJYC9j
ot/EMWqu1DecKQGDyNeSVcJFYr/+lcw/7bFr8NvfhnftXxkmThL036NIOksVhBft4TWnBJdaHREq
wb/JFA+EwMNoUMegDZNpevLAGBUIpN4wbpzneu6Bxfk5wxGuSEpxp38Xh/0Qc7yKxG+3wo0+uPkI
mVwdTpFdLTIttVLcW0PmHNK1yPNfJAYVPk4s+fOV/rXE4jaYL5MnGcFqGhm7O07JI65QOLR5tU6L
dOq7eycR6OeBFwV9Icb1XqsD20SLrzxVHGMP+Ld1+ib5YM3WHDpph3RH38B1TC8d6Od/xEJ6vwot
vl+FRLdYBj1bOAj6lZukYCctQwhsP1CPTWEaXX+g9ghcYNbq4vCFYblTMS4cBJ6nELih/A8xL7eI
6Rp0EPQKBh8w9vZFhgvxgflm41WqvUaFgFfWOpf3JH/9T9ttXaJs2iLW6zAPrlTyPzLc6qRvx9kj
RMtW9YGwNq4h4Dd/PKCJybnJ69MCTUDNS7gcqV1FRVGiG/+Mu8LqI3KkS24HOlRv4G/D9FJEyXl5
ssHXo3MBNbqYZUfx7mSs4h8szzdrxcR1Ry19HdnREkzqmTqgs4TYI8a0YuXjFMIwbB2t5jltlfRQ
32q+IHVz28sQKrswdKwDV6yzVUnrRU6sbx8/tJ8TSSQpMMzTAvOXDgXXJmhepv/Mb4RaFt2gG/7H
XZyMEzPr74icxfLpP4PxxrCjLhtwmLO707qCNo+Uk+jIA5ZDBrcj19kF5ReIwzDbzskZ8mb+MiGT
RS6Bwig3ennGhZsxTT1s5vK3OMJFlrQiNy05m6miEIlA3HJCGlYYZXlSJhUZEyL1tocDf1j9StjM
D8HTwBdMCR3dBPg+ClGhwhyll2jzM2lc2KiyOnzhqGBjc2JhDDP1B4E4dXChdrQx5Lym4QJ5ywdz
3Z9xsFP10hPsjBB2HcSB4nNj7N1viYqTvPXH9MFyx58wreQdyohC2Y0Yp65QDKv/PLnpeNgXDpve
arPINXrUG9vFpCNxj+98RgBTlEGs8+WULwa/Z3abcKsNyp7z1ZsE3bB04I1j8CnYpvrzH9BwqAAq
qjEi15GbE1RfVmN0aVYZKysosyWZ7uvDUaeg0V7AJKhZ9+jN57HE114KumyoVcqe/zU8ioW+e3kB
J1h0pMlJj853noRne72QAM0x3czb44Fyg9fSoDZyrUasGiiSLnu3yI9qEeBEjRRUfoxzdzjaMAp+
FGXM0aadZCuK8rfFS0FvzBXIh5I1wHmF3ZkJJRW86wSerNj/yCr1D6caaJamHShtCMlpai07j+hl
47tpgy4yhxM0k8Nb4TzwAArtHRvh23bzqMcIKKuDLZn5QSfhCKx+80HvN4i7z6xlIUM5MtISC/Dm
e9JxYRx8xsuipE90JXMfzsqTzgJ8az419YGfrWn6tEcP3PT9itrgqgCvDO+jnimmE4FkZj5IPX89
/mvTDdl1JnW8nbdyLzBF8r0qG1mJT63GMiiT5q+jhUNkIWHJeqSitZTyv2t5DoAQUpU5On1o3DHK
LExVOHM8QxSnBnxRkYY7itzeOeFDpZJ50XvEOf8aO6HytgxCA7oDOeihD9S0kN+5ZvYFhS7mKdCN
HsK0kOgpIsN9t+UyQX7w9olqHOD8/HErBANYH9pxk2THu86EgmRDi3Mh9cM3KX83eqznsqZTtmr4
1zIKG3/8eq5ukwbcWncJ80cDXJpeFDVr8d3AFMIuV0FXUxxguv/OaM5AxlljTf3UKBOspReu1TST
3Tk68kHC7zIdz8P46gMpD+7xCL6YwqW14+M+0YLWQUrg2u6bWO/1QVDnLtqEZxrKRI0/kQd3j/sN
TP40LjyMIhA4lyM64kNqUFxX+Y0v46dVRwZGcsMuHpqTwiad2PdY606GFYulGF8IqaGMAzQLs/c3
y/n0uYxxRbXRgW7fRUJ1N/djMOU6LFekx5kafO4MBRz+4wB4Rm63mdNPrwLHw+sZNq75YUrYq2v2
AZF3Vnq8c2XfKoxURJh6bVPBuiyFvIf6vkOUfFd0+PB7s+oN2oIVjSOAAAKz2UCe21qE6atgyyYy
9YZct5VXBrEgN7Y6LjtNcagjupVFSo5rhKzSuWeIgFMnyZrJLi7QNTwEYDibFcjSB7RrQVMKkuJ+
UYXkSIxAUFqrIsWHEESXVlKRzYLheej1xY9vCHNiNdJYm/Sx+Oy1PmKZCpAKcJwxklLORE5BiCER
8MIYjSQ5b+lXH9HpddLd3l0GfZe4NhDoh4uLcBrIHOtL/YN2i0AdX0I3uRNPSd12ugma1F+61/lm
X2r0JQ70L1Qn/Frhv9/vmVANorhhFWF+sYKakJZvE92Svjh2GfUPdmSRaW99wOP8+YbwcyH+9MmW
aq4tCxSbtQZwOjeCetD+eEbNDro3sgLHRjzukgoDr95qHaB4bMJQTRrDQQ890yik1DDeHlM/c5E7
P60IY6mMDVjcHevt/aYqk/Jmt4K8JUUvvLky5k3AVu2Pd1CiLw0xcW4dD07L5Wa89KVBvW2AdxkX
PQGbFi9hSceohLUjSrKWbFhmOd2gIKU2Ee2TPmo+mxy1UObbUraT5YAwOv04FThARjqu2rNASUyK
Lb78tXRhx/OddqcT5a8WxuA9yE4wVg4QunOsoQOXvWxgWmjgDOpUj9cXD0E/grix2BvMmweHapAC
ZRa09sluGwkl9v401jULpiRIvVjyFKifZJYa8qZF1LsN3Qkmo4aioYvIXTXqx2dE2mEpGymw+7hS
32Hi9ji19FyNoXgOlgE9OC8+zntgnYAUh+EW5eG/rryhE0bNSp7ygextQF90ju0Z+im1TPCfPOol
GH3E7ovu+va9t3kaKmRxVMx0QZDaDp642tKkCb/6G6gzCcw//LS/NB2IjGLEAoAmlA88Ck86OAj/
AHEtuUP/w71toKkZUhWyVr6NaA1fn87ua3L9JbvAENKg3OgBubzg6mppFtmbwMReKfOnGlSA3Hni
Vh5BiL6fcwsvajIm/5gWN8O6YR6uOKxWAeyejb0rhN7AToibKMjki3+uH3ZIQcBgg6PS7nT15wEH
chDGmwF+68zRsKx9jxmgE2kKL6SeSFz/jPUfcmz5rD/WzwKSL0wdOdull9aj6PeRh3N+OCRtq9Qn
oHm6j7nY+OXNGU//dbD5THDoq/DI9vYu3iuyUes1pNmDYuOgvwEZH2PndlnIvs31umjb6pAf2g4R
qShpEHeqEiQkjTRKKI8g7IUwhRjQwBBCgAWmT3VI6cJxxMeGqA6LEbSn0JeFpLOvERkdPzykaTKl
sMp/4qGOo+1EdU0Xkjch7jjwxfhK2Qe12bpS0PkFwZJrJO17HrkjqjZqN/0CvZHCkA73WDFpFIK9
vdm1cagX6/dUmrqv6qsSK2EGqTMSY/7EE8KkaE+CKw3xkyrJ5AfNxJcuXUkXlSYkEeSwo0MmSaZG
vCWvQEVEzxljqt+cH34RyCp+gZxClgYmX7T60C++5JNnjrsABxiHwg18TNDIpDvX09UJWIRm86mR
PjDjj36DFleTZWKeCf5vWJdxU9Bz2BIXKMGEAngaDkzTkRvB6z/g28ail6BZiLCpt2xldQ6IXsYN
tLBhzVK/lVga1p7TPoUtoKwVORFIytphtFktfvLo0rY/Ny4fV9dVsYUs/R5OuZlsjR1ygx2lYVrt
WVbFIYrvpqmgIQv9Sw5+4ltNSC/ByDwWq38QXfWc6mjJWReVUmtp49H8dMP9Q52SyA/v7Byitwfq
Lqg0M6Udpoc3IIGN6EggKBjYbvbmJdHtKuJfu6zhrYN2qTreTRtGk8QqTdj9fT6Y7srkHL+x9iPQ
9JhN/4eFU8Is//DWzOyIW6ERJCZtB3/d4yk/ykB0vg0xcGJkCrzjr6O4mlhXJlkh+STwUf8YMEbC
LkbEq8CILdZq5IDfIWjAx83p94dgcdXaJ3gJujQg9sPErVynCBDWBb2ymj1u6R4AUMrbwGX9XfWH
bZU57P08bP3ml5mTK1CaxkIYQbq4gMHQi1Fc9gyRlebvLYYvBnpMZro86p7aTyKXBO8FuyKwBlCe
YZeJ7WdSJpZn/C9K79eMfswPxwAPa2R5UzmA4wtue4qNkcVnmoLpX3pHv8x7syg5qomeosjUUExX
oqDY2HXt1IjNXB/NWzwRGzl0ULjHvTv/qy5jk2LJb/R+41WdJzdP9eDC97EBGgTq9q9BJVrQ9sYA
d0hQ9EVHhTWO35XbuoU7hlRPaLD81qWGO24jiN14HZsuCuzjqdt/dDJY4hRvrX1MNfRb+v7nNy6s
R0cT5LAuQNQWBgShq+yd2GTv1sefSBIRFE57LJOiTImpzeehnhyMCiysm1i0DhngMPnZQxG3dVn6
kv4wQhkoyoLBNe1EjzeqRRlRuze76FT2JX5rUAKV7hPz60ueJhDl8ue0oZfjfMkPOZDNQoaBg4Vm
W46YGMqEGKaQofzOu1bxCvoRToRwTYQQwG5+xwqsrSmFUb4EcnOfWb3uP0BbWyssZ0CAfqDGd62f
ir+IP0UYCuWG1DMLFhqnJbfU34oWdmjMInHUYnFRb0WxwLJ9tGh6x03qUSftU3rnLr0ZrT0pqkqP
1yUTpbqpPeGe9JATpHe6GPyVrG0AxprB2LTa0EpP2wzg/8VTdv/B5WfQutHWEg54nhew8jkVFMyW
UuxPyAM1WPk5DwOGDZCLJWjFzsNukvYCsTxkWHaZsHZO4QL8mtqS5wcmTf6Vn+lHj9xcOwjw41Xi
Xy6XEiM8HZ0496LgRivwSLq4/4PrnDItqBnCf4qzcs8JKlLzBTLS3P99MQp97oulhLXYcQ+i06Gg
0m+/HbnbtflTtrRpuDsDBV6TvT1jmWJvJFzztNckQJZY6UBtwkVjOTjgLFIJCaCauqsgVW/kxiuk
GsAfe7HjFuQiRzzXFCB04vcvT/mIDJVwD1wyYxIWxnNFI6c3KP+Sk3SDae2RwrQTOzpyanUQQztv
xHuPt4gskOO66cup2eK6NsOHnLthvSv6k+KIA6j8T41d/7AGMq8xX6KuEIBSgRlAolv9pA46JalW
AoWBlDm05KPyDy9mp8h4UwkwqE/diVgEHPpBPXmj/o9izIYjcFpJKxULoonCilML6MY/jBZDq+xy
dbESokdRUSOQQbO3+PuWM38N4sA2juYnB4iNI3KuRJmE2kWoF5Dom1i4lnfJxYI30Ofj7/J1GcVM
VWCPUGmPyZByzOgOBSmLTwKHS4vxRPkDhzWR7WebAaU44qtsGMtxo4reKtkL0vMMCY/L+u1OHnbZ
uvk3LEmPuLulmEQgNZIP2dEZmpdMbyfwhpMPiVXGh6YWBgB4918pK6hWMPkuuF5DFHBsVjOFHwsk
ExHpcRxZOnZKuk/aGa5pxUChSALN8nJ4dn8KBxFC0C8xxUIWm1PCEA/7UDdCl5mErSIss2qFNotp
fmpqhNuiQah0nLwUyGng+UA3naMH6FUsJn4I3FOVWi68ZpUhQ5r9aSXkMzxVozu7k7U5J0wBDwoF
QXF5pPwbkCyfnOTEcwJaVPn2pzRhx4ihZOG7TxUgWOmrRyd46w87xnlw3cKypLVd2IqJzPBERDGJ
iLHAv3xPPxbTw/ttCYmZXZ5Ev0ZWdPx2UZyt3xtFrc1DpGHUYrVTCVPXMRUUT1ZRC5d0dGoW7Pcg
iT3Wp6eHV4La2V+XgkR/UjSYQI9aIgFqsSmAYX61SYvnL6yyT6IQ3mvh7VZNIEf/A4BGxhrdCRhR
ZQkNNnEsZk4CODVOR06fSA==
`protect end_protected

