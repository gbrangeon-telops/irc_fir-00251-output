

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
UXXDHK9d3YtwspCksVg3cn1OQkWFk3QQ1bnN8kcpv130B5dMgVD8+qx+9EwjTR0JFb8FYrcL/7dg
lIwdmlKGHQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
lGlirTrah5ntgtsTqcFN8kWYeCxRHbehSLZqyiEvescJE+ORKShYIOu42/ExCc8hSawNVl9qCirT
UlThiM+Fc1evKMQYzaFIzbKiio/Xw8rjRfhTJKjaxdK3T87LnrHcsuSrci+tl+anpBCM3X47tPxD
oNmgZzATBY/NVtZsbvA=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
UAOAU0ylQuQrszr15mLZsCg4shnqFlxQBAKcqwUoJfM+lTESkAcOosPqKsRH4IbbLlaKiP2HCFU1
aKEFZccPWIgd9WlvneNU3oFbpPCOyV9eZTCX4e5jNTf/7OwRRATKc0mjpd4lxBL9xFrSwNaUKgs1
3vjH77tdesEDAIn5GZ1C/7l3wjwnB4tAiaRNqLY90lB834tlc4mPcP6x8L3rhv5EXfqU4jyJC8B1
4zsO/vH5+VVa1595cRZ3xWXEGVMvmWhY+6TDUJCMhztjp+p4kbQ87UqJz9ddvZWB4hRfjo99Os6I
PqyD9P7zikHIa7jafFMtZu0Vj7u4HDelVYnPyw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
qRFhWXCy25iIpt8SG9Mt+xW3HRp/MFye1jJpn72azeuP+g/A4uHCFxvcKVhzcuE8lYDqFZ9IBM4P
ZjcyPOhURivBaWk0KosUyfzbkORd8yS5XcayTSj5/d+90PPk5PXVCLjTrcMbg0+NO3tiyKtPpLQJ
f+Ih38e2az80fHBgiqo=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
tjh0p4bhQQ++Enuq/zxHJnIk+bY5nNzFWlWKnTVXUtnLIlVGko6ShpeQRaCrGzeMC58aHThmj0Rv
eUmPmT2uqc307TRbbuUeFDYMANj1kcC6Ygs+bdXnSkWnOQFu5reSEq5SE7OMIvzdCIaR/FDvSj26
cuj56WGV7WVTg7EZvTcQQsjBPGe7MBQPj6gVbjkHGUTFOQ09cS9h1BaC9UWWfJNQjyJE48PH9w0J
tqmbE8H5AkyiSVZzE1dyYA/E3WjYX0ib/4FRIxCW96Qs02ypuSbfnvJpIyeRwyQL7ko2qezd2p0h
VgIw3omrmALcnzzjpdcOgkkF7sgouCeIApSqBQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 51440)
`protect data_block
ddV+NGq31GAGZDdfmzqgol5eQQPEAfeJ+w30fL4MCepdAgJ+JLYJQ2sR8ReVveJc6mFnPR+s30NF
Y9Ev1g00zTfHV6MY57QLYELFXFnDG7uRsSIXIoNqR32m1C41eFIUxM5r4tGSed3sB7Tgu67XV1Lk
CWvzNM8yinhURj2lAx4mcc8Yu9N1cF5Ot7Mreqhp3MxvjOcB07xTnnYBEQSbUFQIPgkGLPhhdwRx
eOUzVoTGChflVRMbDUu9dj7yEFenwgI+wDDaimzxcqYbb1kgx6FY2FKjdHZeR6gepqGNVtFLHfI1
itjy3IssK7jJIwWXFmM/MgNzohXdmRMRmd9JsYrzOor3LRV6KuWXivxkjDPIMF+XVs114y4c6lDT
gIzviD1pfdvML46fpXpSd45LnNHiDsrfoi9hfEC3X6TC8X8l7LnD3jQm1l6XvWWIh4VsSir3HFY7
nLccK32E9TtwKfOEqGP5UliEvWQ2tA2wuYejq1B1iolkawYVzidIMqYBCtayxvUyoRilQDt14n0a
yp5jrYo1YPgQpsu3OxFYVxhOQjnw07Bli20nPxB4nJWMFF99NWvtgg1LvZ2sMKJ3ebJXXu+dDjjO
qOd91G7gzny5ZlfTAz7FOB9jc6lB1J+3iHS0txB6rv/4/7u5lMa3NNy4PU0xrRZ+wzYnqQOqPh43
2CZyEv4PQQ9ncC+5kUpoKjNLRmDM1fbFhwW9SvR6uHPtyagxk6BFCWNZiOQCkDpILRSkHUtubyZn
h8a1kAcB0Ic6L/adymQ0o8BInoH/35nDLhyYbA5i/kN6qlU4+jy8kMfuy4ubAtqY4QnBIj4AFwZD
h6ufkg0LBUF24g4zl0sZBXPEYncjUkAXkULT5496w2RYveqbfbKYdgmGHe7EfhEqg4OT5uM6NknF
VDPdVwV/vA5p52bl7cQLfwsuNNRKa49Ap6+/QEu3NBKput3FopwufyrOzf2T3a9J15ELi8Nb9RVd
puNEsITS77v7xH9CrbdGm7oc2HwZyMizuleCtmjvXQM/e3RcZgS+g0XqdfjYARAEVo8sidneowTW
o24nsjr7LkfySr4whpKxcuOlYC8mm7du0rPRJIdM5TXcUBe1BvNZvi2D1H8B2FJBNCfc+y6kT1ea
mE0ssx9heH4QsgmyZhrPlcDaP00/+K5cCtDX7Manx6F1u6alM6eTqZz6vITk/s9GnP5K8i3mpYJt
qfdIY9ayzyrTAea3wNyG68977V2wSmuf3Sg325lkiZUxFco8juA3TUcRvj4EP6My/lZv9gCOULTS
Mh+V/FkxfwASMqx7zCmNOMMa0w8sbcpL1aQhwUcne7UlKj3pQ2O8cQ+Mk1CiPzWDEYZWbUav28DF
rY/Cn7cAwjXM9uY4Bj3PeU813OPjYNA1IdNInpDS299wgUXqME81mOQ4l58T6VZJQ36nFx6jc3Ld
pJvoLgDQ7jmtY94ZScov5nwuHOtqU3CzFSF7xDT2lCRJDGuKIDck4ySH5go4xenSkJHZfG3P7EzZ
nYnc5ut8YU+kdBoAna3+5VhDg4V6Nd3JDGTGY0qAlbiN8H3B1vYhKqFbwmtmj34+k5WWw0AnUX2A
wZ7A8hAfrXhVRkXcEx/gO3mBNekipCv2Zd+eep2GWvBqqwf5ZbSN3NBsAZf0j5qgOcHbFpb5lnCF
MwWdY9xKBd37GO497hioaoop72OcTv94ZsLQl7X1495wf9M/MxvJrX8lK1ZsL/Y6X9r/gpDcgLhF
o3FuvnAjuIMhuvcEE/njwCkhWcqKDbA8sEIqkHJSHrbQ9NcuHxAlJdrnIj16cSrcxUGOcIt85efX
HvTaQPaWgcfXQenPuSW/R/1IE+SN7xY0F5WBfK6eD0Z1wAUQ4B8bzKBqKdd8opme2VIZRtKZ42Xu
SbGmvyNnYU89tLnQP9xtIUX/7w+Z7VOvbmgzRRDqqzTe/7QFnDYM9xZDxlLodXdxOhl7kvQay9b2
gYofgTCyuUc5JQPdoaA+2p9TsKHTBRwohKwV2+qL5EGylw/c6OSuit21yjLPVvpUQ2IXcArJ1/p9
eS3ybVBM1lNyZ280ycVmo8RCy3xZYJcbfayaRLkjQ1VOmYxQO18DX306wi2aAKON+h7vXLIschR/
l9Elj3YSiG8fyGA4IqUKSKETqXcZbKuVZmpQy+wY5pCfk4MvCnEHAIgdTpZZsvm3Jm/YWjvBM7nv
i7PNFuxmS524yznR0hsI1xNEdkiqVB4N+nnp0rnmdAXqxprDInSSRdmzs5wvs10zKLqNURzi/EHX
9IzyY7iCaI2e+cfAMjBkhai9hsoidB66thQo76sDgKPWga40DSBdSNN1dDxTDk80DlWGxPSnmjGa
BJgwdh7nO3lj/li/yfgfg1aVmfvdTlfMLjXXJEdZjoFYRWqHS/9e6T2BPynQJJV1bzp0NpcKhnqd
gHSBdgxisLzVzYYpLd5r4bQ8BSl6A6TmUkwjuzUwYn0L07SJz3YwvXq09XW5NppQHxRDm5epj/zc
ArJhvsprCEc9YOv/79pCD5+aR2kwebUp/6pqdnTvBsATMibeVuA9wXU1oFj1fu7uVJ488bAB7tB+
evc8PK16DPpc1AVtjsZGlibkuZSOiW4LRvG3mIiPdhUslbDPaGbJdwe9ATbiV1FPJzEhQsYm7rb8
MBZqWZF+f7mmvw5jTlwW2QX88Dv/5pgJHi+SUElFwxev0y5bEjT0NEtayNy9R05dAk1ItWBsZLo5
4C3BFioOAWNrRp/+Oee08RQ8Uymq70QQI04Nb+aq43m2WeAAS0V+ndLwKzeIGAk3l1WionkHOVnC
0BfB7drbrRhEIghqjWsH6mnlyaWAR58X9FWz75WRKhZZFrHeU4Z3fy+DFy1QfrwyLB4VtWCS4UbF
1hghSfVvOzJvb0PE9p3xmgeYcSHhRmu012EuW5VDrhw2dczQZeRcU4saKDiK01VpP3ACNQolfpzQ
GhelK/SRd1VjWgVaHuPotjDFAgCy4YXOrcmCy7IRAZpuFyLMsoxspURjErzVUYihyY0vVclIiXaB
9S8bWoqP7dNbxJEoXDcHh7tCeT+nOosBmypMPhdsTeHwLiqpLYQdMlUYEfGHB+sH9LIpWFfLId+n
nGNZsrgrN/2J4c5CM2Z/oar2wbjzh6lYTWxQXr5wIH2EXGaOJ3InkygYv2zusGHnvzkrE8phnVv3
0/2m6SUpSv3RYZwvKL+3DknNKxccmRzS3SKQ72jXpHO9Zzd7GndVaSDOHP9xISoH6vLYp+XxV8tu
lQyudImgF8ztk7XeplVAqtBB1wgzX3FxCGxnT0nrA2Odca01LMvjVs0gX9h2yC1uGDi18uE2q8O7
LOH4zDW9KUbwLuPBP+Bv7SREfoyx+Uo+1FNV+aavD2TovYf/9G6UMp0IRhVk+lIvJePGEYrSEInM
cYFOxQqhB7ud58GUqNcV/IMTlpiONuPkWIVcwwpcqjbVWO0Ds1oph/zfLnB8fyxgomNE5If1F7vB
oi2YIjlGuSj/dxae+XGT97jwMG2ncWPbFfQjMRYM/trIbAqqpD/WSFRqvFcS5Ttxpancutv3+6P6
42XG2FpeV+F8/jPk2vX5NsQkHBT4z/lqFnyo40YW6zhExA8CO6R78hLziwHWu6RWwtxos/LhkdHc
ChZWI2xE0+72631C+9p65CwA59mF0aihNThYGTlw26sxL0lkTtZIoc9+xacOotmoQOQ8hDK9RkKw
XVb7adzMXu/rnlKA4srAO1wYT1TsIbRjIU+IlFXREt3EwSWUeqYDdey4QoCH8TB1Y12tl4Sxfiml
5/hOrEsgFao3qUKxF3Q2w0Y3DbmrCLPhDC62H0Bb3eFh/N6cU5UOLBHJfc5D1wLeWps5PEAFvHoE
TwIQqGqyQIQ9y5Dgk/z8M6kvhxAjaByGVz+I30+P8XbNfab0qq7/VxJKI4JrH2B5aS7uV+ZFXiDO
6WWH6iyCpjsIeS/4UEZeFcKvqfMmECsmw6RcEYqbzi+d3lxsx8su3f2Sst4z2ZtujSof7zTOacKF
qnLnlVFrmkF24QIk0W3zJ5lfZE9f4XaLQLPE3YLLeAElocp4ieHByInUbwTVJJpOeBPdPUtT2DQB
idIfgTwQ2D9g5cWKeCBzO2q+bv7yNEffWUS0ROt9i1Ey3mbbyc02cQ1ekhpv3aisk30Me2Z+SMS7
v12EZiAOV0GkRt/Cb3yAfVFJ5gDy30c9UK7hBdfXUSg/1UpYCWUbBDQMT/CPTz7j95ht4A3uC9fT
s6+GVznNNaCY8Ttay4y3ni8Q4yXGhCCq+J4AqFJ9jgLVfxjKl0tEex8tQz1X6DcaDI+azJjpLZ16
0PaMnOZHsFAj8vBONqkvdY0zsH+ImFI6pnvvO1/Pxjs4u1L1lD05FEt9qZUm0NpyEWcph25Bfzd2
hznzm5soei3rVt8NEQ10D43Wjrzg+XjCSKdOblCj2XI4Mc6xCydu5WWmB0pKNM5Tbk+Nja0WFudN
gx7O2swM6zYW5XkcmBK0fPvR9J8GgYJRmrnqfuJ3GwTvhX3Dgrf1no1VE9d20Fj+wIkRC+Bz2Wd8
xRAfVLnrH/IdEZBPp9yvkaOqPdKCs/RMlSR2RWRMhdL+9O0du9hDH3Mf8R7hCV+H8chHorWg6f+J
aOggnpuBd1NuMDmAziHLEX1XvqykIV8uF6fj7m8eV5IGqazuTxTo0/oF7gTdAa6ONYGX7iBjIrJe
3+5YdAG7Z86hAmPF1QryMfHuZmAHXavbELKEOsek4TNCwiPwdVRUsOX3LqU3NcFNCbisBEAimN94
5dYE3/hgIk7OS9RhQI/pHfFj+9zIs7qQv0KtMrde+dNPcqQfNJdWwH3TSgsS87y92jkHcqewR2W/
g82epq5hqiJXs7VPh1pSztYihQwbcJpiYRJlaL3F+fXcDyg2G8tx18BY19RfIn0JeflmIGH1MQp1
Wab4p77NK0sokgrnoU18Ly9wEDchTwio+9zRNiCH4IfFxUku1ePZjo2JS3HlfNepghYNyphW8sca
pfSfqXBbsk+ADsyPuH+hm6+KBtqiU2+BRBMGylZS5DywUbXQFLE2rvyT/tjSDwjAq9kgr6/J2rLI
qLvfdIxYVUwGLUiE1NUIizLqFIJ7o6/xFjhAXgbGoAxHExPdhIKb9Yh66DXsPovDVknnz03vZXwV
pw40n5AimRy0DCPrHBbq2G3G/KCJN4n2HINXtWhqgVHI0TNwckKf7a5c822OvmKJ1x9OgU+rTJHL
HbJrNCqd3+Ev7gj2RYtwA7f7exTg7/5JHR0Bz59zqjV81LQME1Jxmpx8PNbeDm9UmAvTy+cKlGZv
KAnULybN+0gW5K4SUrOUzF3VL+nnrl35UpRoBsxUsOEg0jTg3eBLibqmySMBWCxtcZwxK0o0qSsD
UlMDfIHfsf7Z496jO2CiMTkf5/67zalMuHBvOYR1TQMDcYuMGEdwUBr2WWxPp2DHDPso5BimdIvB
rrl0PR3ixd2DIomy9eqxqKKKY/JVhovm6rClz6VgaInmjRLdPBmtZHVuKUHL0md9aRhUZbCQyO52
YXlqxaxW0X/lAVpoftresKY5m56NtDEubFRcrWKTO5YAmQwHk7wbrMT/xkV8g1+1tOnpoVmkNaOk
hhkppy6TU6Ta5ZyzJxcr6TU6rvZLWP3O6x70UV1trQqX7yNRMRC4S96sf/a00D+Z222D1DtqdOzj
e0Y3DfAGemZqASDszWuwdmi7QbcBK/M0Il0bsrIf+50L1JiLDipSa0Zuc54fUPwlNyL5q4PBLYlH
OpZv9bXW6Kg8hPcq0hciq3jrZ7ZVw3vguseEnPCVI4FQWdtNXwz2jJD6igS/WdQ9GpqXKHZ648BK
E6QOk41cDt63vwf6oNRcAsXIsU7+xRYjQJsjRmuk4hzhvC4dCqXSIeVjEywqkJ0rdXA10QhCNpd1
Dw8ag3OQyFOKDvGDJgIaOaL6ymziG0LCzRMoDhOOqDGbk240od08zECVNuAR6/dMEdOSFMY0+Cnf
T64zW4kiTA3L2NHf9CWvL4OdG4/4PYSX62LnVYOuCU1pVc6Ch6FsIW41LT1ftjFQaeiePndoX+PB
4xhhxWUQI4/1yTk+cGD2xwKWRRdr+dOkbgQjIcoQUUaODfQ1NLXvjacWS31KoJDVDmw/RT8Pv7Ji
/u/SlWBe+LkX+O52f7Zy+jscQ18VxyyZnx0ymhbn1aU3iUXsLPScgUVeEJTG76YrckagWgw7xN2K
5jaDBvEWz6TEPFIslKylRxTYwgqYnh5/bHBJiMzuA+SdxSKUM/IsFrsiq4E1eXi7G2e9y/Z8bNFc
C4A7TNAc5lwuPAKcWT36x6AjeJ7o7k80g4AiJ/zQ3ufEIQpaC2ghWr89qLB0QFxKmqIWWKRPOfpv
gE71iG8dXYGZ0AZopg6GZ0MD1QlUSThdxYfvLrsOt4LoUZU3zIebToGvTG3zaGYFWQfcz5Xcxo+e
2CTiwyVKD+8rFOTU1Xrq5GAqvivdp0lY+cSqJVM7sar2r2buwVYnacwMIsHGvVQVN+X/u6XnB2e2
Y4E1ZmOhe7RkLdhCvualugZ11wfQoBzagI5R2t8iPBM6FyeqWxk8A9ZzTvO52cCC0IuJqKteib1W
AZmdD836yg4ZW/0B6fv8ZjfNj9dvK5lYaK8q6nSVDvc2sdvTwnecoXLpePR+0ZQJbHwIq1lWrELD
EnY0rQZvm4bdilpG9LKOpi0UFaCmUFHJewrA/Ox5NHqGVWvaTnnCFN14Uco+wEYFYX753lBOVZ/5
wDBgU4m2uPLKYur1NXkvy3JViVMTPaBq1gbqK8t09UyLpH9oE+TdWS5UGClLQ6utrW3gJ11TQUD7
31kMZRCwyuW5eGUb+qeh9g0OHQ6+mYU9q+GDDwwcVwXO5QohJZuZTglXyuDD9niukE4u+CniEtdO
TnlNvkDl2McNvgTFEHPHBCHVWJWynarFdS3xUK6PZkIMtarNrqZrw70nVIO5fd+ctF11/QdN27Hu
vSIGomOS0513lmacLWKne9ockQCyMytau/chvfqzODFq2tYRLlma6jWWbJdvMFRNldr+EdwVnxo+
MLwpexCPJW+czkzYy9MMSLJMxFZBfpcYr1WAnH+/DRQoGUlF+ylsSJcmJgKQykU+wAc7u4E78ns/
YKa0qG5UdoJth7HW5afHcVpFm0cauuK55LLJOm7t+H6/xMzuH7A5ToLuZhJyj+EcKETkSEqAW/8p
bZELgDXaWB5RQqTp+nmezykszQGUtjBF354yIuXepG+Y21WxTzcKufF5d1Nn4o2EHJU3B8/d3CIY
4Y/lK1lbY6CSw6G5TP2Sr79RfWANhzCJ4fQ9AitT6zn24F+kSevIj7m59dW/CGwWKihhWn070Ljc
qYkYGEDL0/RYIlVJwJsMzoD3GIseoIJrd+ICPYJXVRdley3U7+kUu5KoZPGsKYriqD9gmRHluhw8
pyyYAxRL+Vs0Q5OiTmV16TyEISHvyu2tTZl2PzKqkeRTF3hQW+soxGj2/f1ff4KZ8w5IeN6Mo/d0
cbKtXyxbcIGEmzC+68onUct7JLy9TiB3TZYrFUYI+3IsZM97fEYl1qr+OFxzO9Zy3DU+iKpxqM0Q
T3kC8u+vUGWGjyqPMi0mE4NnOe3M6EbaPFa29ZIX3fjSeokCdohOs3YexFgayt0ewZAQz7Bp0b/2
DS4r9Yl05Silfts3RNIpS8+inDyT0dcD6QNIDu6gXSpkKXfarXgmmR7aRz901U9lUtfNAuEQAyiU
UFhABQ5Xn1tthw2d5Tou2FqnrYKQR5laqoFq7yIsHkkIfASzdi+lHxMai9ts3S3YfWGk+NdAhGvB
SiNCa4vfRZkxCtqnrFOenP0Ci4g9FzgWYOI+B1fCq8KMBuCLkQxNNvrmUfSBSQa4tWUeMcOHg9jt
tZ5B2IeXRl4NkurQYgpCjGN3JBGJgKnZ+chatwSstZUkNBtlLH+320OOsrN6vls/Rz1drjBtOgrn
06DSvaG9QezO7MSjd3yxNXsYxdmyT38xlclfh0W59t2leY4mHhq30Ds2UOFtSBmg+o4WU5InWtb2
vZF5IRsnozt/oI6/aMf/UKuvSTIsx31r3bHfmBNBTkeCQ6DW9SwLQnEjdVZ0i7THm3s8iIA/uwhA
U7T5prbJylG2vMlEoeo1N8ghDOtLOmc5JphaljWsmmkEZpswwP8PUIAyzp7/fiTfDGVdONoMhzSR
7/FEfWs0HKZ/hbrsBuLlZ+LxnSBSg60Rtg78aWVsSUj/EtDB83FpX6uIccl1qRr40Eo37xZVu04U
NWuebSTQABZwp59F8V0K88FaQeB8o1lViNBKwHTgJnAWB/lwOK14ljtxgjaoh9kGabQcYT9qTOqF
SstSNEIU/OVHTf0p/WKe/oL8YKkBJXEP4t50bc8eskqzUw7k7ElmeMmpeiGOWFMdDupXIelC7UYa
5TQvimixdS60y9dKtVqHdEfu5ekWT//FKpfcItPKq376uPkWA3AlwAmGpAgg4p2i111LMeRCBr63
MEO/mFKi/YRRvyi11NNOXxU/chAvqNMzJkF5vi98E5sw3C65NqJd+sseUTJRtVgn9xNWzf9aTdiP
NtX5HEgOzRQkmPqAvgcZbxDCoZQHgYQSPIhvz1xevd5gH04XXDRWnR5DBOkTIYFGXtoTCPiIVTL7
quFeN5Tp6BwTNB0ucG4nJWlPrMxg/ClyYQbaq4Z9GPBquNIyFhhz9lNdfco+ie/T6H7Ij+Pp+9f/
n6jG3pO3/uoQ6VSXLrT2nP9iFV6W9uthyPP9vdHn2po+b9d1eU0ZBrkKcoKhKlzFukiXcAyFdYaY
M9Z2CkRILK2KR5DhqVwVVC+475CEFbI3hfpT8vyfMoD7/zJ5ec0sNg71cFwF0QBcAsCmPDa2xL5g
Wh385OE4++Z01OlNBtqEHiHu/kTl9jVfkfJcQN/c3YQYT2NoOdvw3axDE4IlryZ9w9JB6sanZiVc
1ZpllQ08mdThfz917tYD7i9nFEQV0RCZqE+s9z9gKtqmAThkZJXUJr7WlVGld7cc/VZjQsMM+7Oc
2uJHubvyBpSKCjX0kH/jGrlHxApCQvD4NSQK+f0bwEsgj76G5dOIj+4ETVV0TR7RzCUP3sp03Oua
XFHYAJuOWrY+sgAwNrTBGs+Zel6xZg64JeO98QwChNBc8VGXdqR9dcudAUJr4XgPVH7nMNDjTXNX
a9e1D9t6br6rUbAO27JPTesUmCIGDmfEnqXOK3sw5EHXx5jwAljLEQYDzyg+UZ4LzfZhD/sxQ5HG
gIcc7MqYsDUXpSm9Afgj69GvDDcMtM9vhsmNQYG/7vqsxl2V0/MoOK+pSHHIHYCNwiGEDztVtsjX
4tI1VjjJ3QdQo3YigcLs00vLjGUpxv1i61iulcXD+zREs3tUGKxxNP9xXvAR+WnU4HFkvmn/ADqf
P25BtIyeNA/8csxSER6PcQGIHM/2HN8KgjiH0n+aFKbaoWgB3LJynM5OZ4lSS/3EfqJvLjjfzt+n
gWdtccgDGifEJP4qeO89l4S8M6R/HvDTAqdeFziept5c5llJo0tepHhjooBKzwCuXtkfWrXwM/fZ
ZQ3UegtrjlBX8RbeAFt4Vsf9GLC9+1oE84PLP4PdA8fNvj7NjHoNB1T/yHKfwNYdm971NOrvBTPb
v2lq1xbzWH1D6vE/VSMMLFUM0dV/3Kf5DZvF4Vi9zd3sRmeHR2YALAKyxcWLdh9M5g963rHajRqY
vSDCFuQZVNepKVXsf6DkbkkyyM+lq7Kn+P4sLgo04M3IafBBsyH7/sZg9XAcJ27VEf2/p8udT14Q
W4d2gtBZafYvX3TJpizsYXiMMkp+kD5+pQb57OgWqIYfZ6CrKGk6zlbPFt6Huch19GyRpi4Tns1B
HrfE+qr0TcETgSTjCK23JPUATzdmjlJbW8Q117M3Tk7Fjf7CqAm06c5ahnaog0hOmedgi4dZO+cP
8Eh0GwoyMkfBtw2HJon4X7WaOy3iIYVT1I13h1OTJDWWn7XXAK8j04K4i78d2sW3p10nNTqTpn9s
/6KpFSPIZGHQoTY4IYzcK2ogTqA119GJSP2iY/LGvvze4qHcNT/yefTW4n/KJ9EXdV9l/FDUCnIt
hsl0LcbbjYWqBDSmar5UH1V5MoQ/Vt9YUWb497mw2e7rV5G4pcQriMgOKFiMQWTzH8aIfaltSffB
PILJ9tt82KjN0JklIIFK2OgCbEhze/0tiRfLENDaV8PDS4ABXEF6SXmr/GOfWG4slnxBs6JwbmW6
YUZEY40JZHXqy8ns/595njcIPFtjqrOibVtrxSaVs3YQN4iM3V8rNE8jKp1n2QNnGVxMygmtf1ZP
8Oy2/1e1cbaqW5ppcSu4b2b4ZpJGBpN1ZmKZ8HMKqnH7psO8eLMeVwG5WjfYa154HhH/kM46+L82
3bIq5Q/gFW1qwa2XhiF11XfV5Ieu9ndkXXORMbPIK2yM7imWK9djnBtIRDxf270tVw9lRcF4kfHE
YK8njU+ee8rsMzZb6s4achG6Bq7tQeo/eTxT2pri5HJAeEltDfVYa4FMSz3mKu9Azbf0nEe30loR
lXhsog3gSqVyDvSsdJ+bgnOdvvRUHaScf6uQXL6dxjiZa+SHYEqnZPkgwDm4xfVeNiEn1yPmpbWt
gNvqonbrShm1sm4bjFan5fWQoA0+asGuQycvSrUwU4ixVMOixS52jn6URrPsel7teWgHXbxZu9ii
X5OUqqRc/1yrrkX/cv4X2NmZBs0+3gOhBFyBk8Ktf6HSLGC/pvEmaFvqig7fiaDXY1ZbvMtvipB8
b+GQKJJnY4vsAP0jJfPMn/7D7y1XBvPxJTOo9OOXNG6fmCAjAdMvMByvWOrtQs1+ELqM+WVMJfGL
M8Aoksh9LwSEzbyPqB1b+OHErrEenEjnltopKzDAla7Ysc7tmJ7y66VMNwCFIJuoxylK2xQ01Opo
ksA8iShiYoSweZe7wjUhnDRac6TKmVRzvwnt9iSc6WCRmnVgViDTvhkxSZdKHFBawPYIXA07zL3Q
lMa7rxhPNFJlhFXco3GXAaSIPk2lV/Q0JzNV981jbmA9h5bBDkR4tkCtcRRiQvZBzY/GIa24eqLC
wbyKDKW0MKMqnIcNA4/Qpt5r5UnMBjnonlSMyZmbMpWNjEzzX24HqU+DHWdbshd0HyGBwP8KF94R
q4xA4f0Cszry3uHranCgM0te5goaxF65mO2FP813cosZFGNiWYANXeLW19QbD3CuA/ystoZR0Gq3
04xyzicVC0PUNkcjOnfNvbs7ZncQ7lo7OYPV9zr8BakWRaGKC1TSzI/X+pgShOivEF/BKXFBZD8S
Xhm7UyphanYf/xxDlt0Gmg/YEPj5lsE8hu9EbTEHd+/Pa4G5JaCI6eAiSeW2cg+4ObRK2k471S3P
3F+jwPDDsIKw3CqVx1zOj5tPXRcID0H/PVlwKzLASoEEjoeHB58FM3quTsCaN+uLJOzRP05Z6s03
1NHn2qMPYBz6NjuK/X21P4JQErFBneHjRQJ7aqQBEDpp3udXIE0kSVqBdpf6XTFm+QhaTJnxmeZd
0IrT3aQb5JnZ5ZzuwebPamnP3JwqJm0BG1Zv6QQxHDs0eozbPIRynbmTwqV9WYdsel1feNBDKICR
dtDqdb30qNhe1fOQt7zY60B0Knhj3iIksSKqF+KAEeeDvv3YOp3DP+m4yLLTQ+BETlzvf7r2eAkp
09l8p9BbAOzOGkN3E4A72RIeajxLsADvyZ0Xwa7vmhur0DFwGu4Pj8A7jNp5nIwASrnxtgQzeVqL
rn3ld20bF+XCD/LYCU+A8H4vQBya+diNF2io2tMe9PyAinShSJ63tyoPQ6cHtms6D+w66YjJSYAz
2/XpZsrOY65Z+A0q9q6kTvxArbCro8bGcwPYp3SOU7EhWdo8XaFcCs4iH8SJP17oDmdmsMkM9WAk
xMHTF4I3rqynT49EFCHVPt8T0jMRN4O7tFViA4biLV0GscZgmWrDhLjGciHDt/zHeqIechzIymVs
hCc5DxerPHz9bpYfG0sRznzK4As5AIwGwaRC0Y4xf4fJprmQdSRCwdZLStdBGkjt/iQixszThF72
h8Z3/O4mGwJyHprFg3l1tY+1zQasDDjMuNqwY0OU2GwRpw+IEoWVIfS/tSXS5ynzNSt/6fHEQtAR
t3YTbj20AquLV9qfnQPhdo345RTFlUJ+Q93U9CqbPkcwPUVty4pprqvbhLmlSF2P/Gzn0+ymR42O
+2Tgqg4q1yCR6ArsDN3unzlVTH5CvKvhO498CVP6qUMHIzZXT4Fzt75AUaFf8caZ3MMn7HTLwlj6
KiRqdhxWxGtbLuoPttmGes5Yi3J2dNm7K7SYygER3UeLSUZfKjg3khbI54+hBhaNGGYJb/87bQQb
d+Mt4KlQOHodiNHvAgEgO+li/oJMS+Vl8NEqVEMuu+wHlOC6Z5BvzU7d2o9b1EBxcG3pJKIeZGci
iigPwEkzkUM/K1pyVR6qLKAmeMjWITg6uBWBVWJBX26lHhvwC+gOvJLbvKpUOB24biv0tihQ2bBa
OX5ZeoTCZ7CkH5eWvXplZ0yCbNEcvBPJXgzoYCHH1kL+6UT0yVOd3spiLXv+iAQE0csMAzPQ+yyD
TL0JNS6fh99EDFDzE6xJCfc0KWSKLWPbbHHMpkhPH1dNYwVpUnh/XjtfGpvJp2S6VZwJ2xPgIvix
xUoACmo6NfSa9aFgO/Y4iNmv4A+JCdaseghvZ1717QmyJF76hwlvQTwFl0kaZNcMf6u6TcsgcUVE
FWpTszODl/uaEt59437SaDTYy8jlwnzzTSiz5ojrZ3/zkYDXiXDBOhfbsEbVIJyN/aFNF1typMLT
N16j2xFqV7yWoyAZS7iH+Z1hqdWlMwlYEegHLw1pNjgHUSTtyj34Pkw4+lagdCw5XTSLkNZnlmCE
jHpGYd+1NuB9fIxQ59LBuJehJiFElNfljbvWn2Q6KMJ6VUuS+ksd3cfQwtga+9QYgpa9L+/iQex1
AFi8je5gp45T9r8VkH+X4QEAlwO40rhJ5CWXn+7STUYJKukP1NSDUed0CN49y6i/+loT62LqKU5c
ul/m9XaBvuixiGKDhiFgOCP9BXnv+DCHeV2y7PIu9601twpytdKxHwoX+U3X5wIEHTTsz2y+qOsn
gBnlYGxJyYwvYTOsZRQzKHhBwsjKzdg3kVg05Wr10AKwzXgqIQE+4V1uxrfQxBLCFLA/YorHLwU1
qPa9JsMnJapygJtVa4WFw41eeQN7wajTCNoken0UVaH2P1GYi9iyn9R1r8lHBSX7svHzQwmpJY21
im/1hu7DBKFMRvcj5usLtGx1L5LCbmzFyMLp3pu6dee4J/euynXFlSUxUcU70BuLE/VWfh+a9VQo
C7keLIIed/T8XXIfJjPqy31N8y+9RTMLYiBAoJOb/+3bhaRgXiIZZmyuQZeOc6yWjx3v0W9mnx/Y
oq4tKv+8cvxjEXSFQvpf0bdDkeBcGSb8wIwCkpIvrcdUQQTC3wvCq18Lr7M0uLardkd4jLExeRnS
RNhKqBXV/SYiqcJ1RkNC8JPX5T28ZJ9cZFdP/GyEYYD+oFlkHI2sHiJ9Xn0SqWqkb9ysCR3cBBtW
WWDYqRgDLwvgSRnhBhFGIllLtHD7fDvwm7IQOPObQY2mCKkGQYE+8O4MNB1+/5fORz2hRauH+tR8
P1OL6c4ZkI8Zihod5rm3sRkON/BWOa8bQEt1DHbk7+uSy9+yfEiGJP/wK2XTCYqJIvEoMrb9mNyu
kv9RsTo0T1t3u8vvQGDJ3545/4Wz/HjnU1qivicev9pGRysPNHYNnv2gtOs3i1cgd6BnAU9RKNWV
di5lTfp0+7Kx6bIelWlAQeNuU30lDuXFfarZgSljl3/X2LMUMJ06I0GRTq3eBHf9GFq7FxCPAt/D
a8sDzLoKdKPCEnBjRYp96UG++Wk0JolssPpZF5BWq1lTSH1bVWavDnD3BOUcL5qb49b59b8BIqwP
dGAKLGaRnLpL9Ac3oWXQHqM2Xt+AOq/ZlALkXzAxxq+vmybdnbXU7yU8RcIA1KYPjk1uD2OaxLrL
6gGjVWrHCwYwA4CLVWLSOHIqt0xJUYR2D3u/dHSa0dTMB6X2NvUSr8xeEFC6n8YV0PeFO5T34Gwq
kevTakOOJbLnxo++sepdVodgWmceOn8g6wEB+xZo0BhgcziiwhXblTimdgWy0aSegNvXxSBglO2F
4m+v1ZlidGfjK377HZXhpDghB1pNJFy5gujD7hJJ5UYXiVGH9KWVI+NJlM4ISTvVeBpUiqocmcdA
qthN2ochHKxjgYNC0JRTOKOSKqUzdE2ssagY84lVpZ3ELD4wxTiBQzcbxoxzsrSGXaSsPbw00rC/
/tWSMBVYAcfaFJfbDKq0w20XseBV6QZ1BOCgzGmc1WozxWBaAbgAZlquGzrh3t9cj4kUYYB/bqAu
BaeXtu0mW1wc7DlbDOBT4B/GKmGRP3FJg/MaCOdWt+rb04Yq/PlnJk3uBJrAjo+WsUOJfw4BiTkP
f5deEIHIZTf/aBKvsnBkIDUzhgcCvmXxr6j3zvhWfGHIOeB601r94Qewn+xp6PwM6IRzzPSSrnIf
LfWv1daViUjyqkCbNZSQPU7zabUvxouqO7+sTiStzjpre5f+7g1rxqtMcCgLw8ON34BJJoOZSDwI
LfiT+LVBbHTGHPOvOD1gAAm+97i67zRMZ02xTyP3DZGu8I71C3q5gz7q7BOdpUbd9L+5uqV7LSMV
opxtCVWvKD14NKZ4dtDP2pVwhi6f49ETaoYZ1+7CVndB2yytKVvaAt6/0YGme+udk1PtdPDlRMym
CwyDPAmnxUd2ip+3V/YTomDS3QrdTM1AACh+vruS3KFLfvHzz/PF+WHv+umlJKdR+W3Xq2vZcRl+
TUV24RNwKnrGsyc26cmTMPsB+6o/ajHKnsDsZaS+YkKkjKLEDclZJz5Aa4penGN48fTZ2ZE5J/Np
U3vBx2WY3Hj6nFepEbaf4os1x6tQ4D+IVAmVXLgyaEomNVL1o3jzXCLY1VDwyymb+5YfK5VTNhNb
+Qnsw0Pv5f1HznALh1L/DbRwt/mqXVbvm1IoTakXSmn0sEuaVn6y9+8vW1YUHCePMXmbwZQ4oZVo
i93uYDVKnhSCrHh5Bduc+goOF1lNy7l/H1Avq1ILYP2N0pFUbryx0o0vH45TdTmJCBqIYpi/xbBt
A8nSw8Xw+adsTtkCwFTHQp9wCJdBILrY4YZigfNgmM5v9/WpUcaVq62k6iDKmEbWLhICixzM2xc6
6NSNMOJza7XCKRfO6JR8dJnsM9ZXvrrvichU7XLi8ZV/q5G4KufPFId7P0e6lzS2eXhlxDWvopCW
gnpOmvHmAS/7GOco7rYA57w40r4fQVIyHGIqM3+SclMdn83WHtjIsDxItj4jZoRzaPnx0NJdhgva
FqAGWMaIkw+Z+mu4nUI2kYssB2vj5PbWmoihLOOuhweN27BqpTG9ktL0Gsdb1UQ6Y7I2QChgT45G
TeOXQQjnci9ElUyAceMU0TP+z+nR7hq8fXx0IUlmTa4KAdwbuoueqsMPJpHh6t3b9SfdPT4aVdZd
zmA9WMihmrAcgRNnJCGaenTShi5sBKEorsbUJiC0JIGasR7zSiUaeDw+63MZva2brKZjzerRy2PP
dlSyd7KM4O/LUwGB/c8bnWy4cZJOtw8vK3g6DqkASntj3ZQB+SCdTYTBtOjnVDfoGYDtdglCT6vo
B4cJG9kFTl4psnxXc6moy5unjoGmVE0I4mTGpcYSgtpMcdWVg0pgt7pDIlZofH0SpTdaDuYCCNi4
J2ENIvXStxdyn7KE3O00LnvL1coI/W5os73S3dCgqrGs2nPcklpqnxDPX3ygzdW+HOPDyLSm35Tz
W37qEQa25bMTtapsmA1MuCGp7d3G3YqyuR58APuC2PfBTBX1sktkP1IS2GvwULxDKo89vgCkoWk/
uoTsRnVs2j7fxdJkp/LwS9vPhXZ2mbUJGzXWPw++knZF0XJ7x7YNBaGJ3MsgxlrhezfnmurUrP4R
vonmoIW82JnC4DKVs3e96SvpwsZOyKngf61d6avJ77To0LUq13Wki7b9b9WZ2uKJATBNiZ3oBs2M
TU7V0HPQVn+/r5fUw87HpZZ0EDfLzmlv3CGRhk9WnxqaO7t2xk74DFQ5WKi5iigGComMdr/hzL2i
e38O95htq9xIyLehOdnYrMdv6HJ3uIVtO4R02GLw1ksel2z5l0ovbIO6QSpOLvJ4uZM9LcQjfXrR
U+xF5/c4QaH7rgq/a5dlD1UEMXs+huM2m9aD5OUi4e36yTeyiDrTMUhT0kmV0rQykBTIuZNiuVP1
azJYQ41CpizI2f8cGiY51vPnGqyJiseBg86FoX9+0BlKTiHTFoIWzeNRskFI6jtoYnTKx+uEMM3Y
dedyGBcfb7qVeMq2i3se41zc+lrwwt2onOOpDygqy8dGnvFVT8CR3lsEsJYxhWQLsfD1/it0Syx9
Yd6ZQlJj9otvqNxaJBlnvDe/017fVY/cPalsQnnnWPhq+ugxyOcd4/VZM8NZDl+dVwVYdi8iG10e
FBpgl5R5m99Ss13rYyyFYAP01Iwlgk6iWrYvYyIURDbsHmbdnPcnNPS+zEIhXjOT6ydf9Zo2/NkH
jmRQJ4R49J7l9kEX4UQqtH+8T+wfp3tVGPacqWKNgrlLe3Kgt174plVuvBy9Nz/9Vz/ifCUX1GOv
Cu9p9JMYH0DpfRDRbi7ZV+xk0pe2mhVrUwTGv+8yem9qD9oR106zOkDAffOKZaOBQQ/PxnTJ0MSn
i5XUMiGKP6mA+T6gROlnog1/dhNNAh9U0fBtH8yXMr0A+DZdMnH0bTFBI+96t0J9ODaq3Qd5x2Tv
beGECXinkbBeVYXCfyf6XKno60cKxOoEuFaS39IvwanY9PBc7iZzy/norytbBsUXRipLmS/arMcl
GHfyEp54M7Jm3qXmKs8IE6HnscitN8i3Mm2t83LC4g4TFn5eEg5t77nWG/VBQxvLIxIpGypOC/gH
dW0WWq5Q8nXuSZ7w5LtgrFOHtMyiPLa1COFruet41C9ViAzUhli+agRFJLWxMAJf6+8ZFs2MXZ7N
h0ZHjFfDGYySgobA5fxlRy4k1RiiKqUz5V5bpXmHs6gJV5GgAgrFPgWr5VmKVrJFM85kjyQbkS7t
7bAy+WVjmj1j36OKFiG/JwkKLWmmcsdn8NecEi1bh9BfOkJ97ufeB2alsCzI3xsHCkqwrcCQcc0c
UI6sjU2RntuZqJxSUOKucKEWLSUMxyEcFN3hjspEi0l/a8I/P6n+Auy7WiESlzsKsNrJ6VZAZuq2
FUsBdZL4XmgGHhztOdf7WsZEQFCaFNE+i3jTWhFvga/RUZWIklp0o6WW0V8OHJMq34uOxvLwy6/9
yC0JaPBz3DpOwreP7fpWn3nC7GXuAyP3thDpMTNZ2XD6hRyrDZT8bWozdokJ3IV0VIagf25/rC3/
S9SgJaCEyt7PDF1piJX8arVc9qVxrkKgrUhdlqrdsbNtmbTXOgm9AHATnOQEy1RMuLM9IcRxz4xI
yqP5kRo7em967W90d0XbVMav97NMic0AG8Bl+pLc/mCCMOT8rJvmtehXjIdNEz+CNCW4jAI3Mzc6
jktseJbzcI2vqDi2uodrSmthGknaFKUckyC14TmvM8C7PJpq4g2aD/36Hb+fPrm12S+/OEDYkRz7
gNGqOjVC/sV2vhthPZoNE/Dxm6prQ5wa15Wh9Wzn7AMuLptOTL8kri1zKpkla8+P+2QvyNd8cXFi
taK0C1ovQlXMf7wcUHsQtScpq2CmfoGc5SCTxhO+0rpU5f/RgSRlfWSygFmnphec3W1ajbtqTbAm
w5Xxd6raOHnR5alPc0WPRUMJOu/laW49QtUa4cJqFXTOPGDD/olHJg9eGw7gGCZ+YJ8qFmGHIcgl
HaRkT4G9QKsdxrSbbCWVARF3H5IeGd01P2LkuICwp8GHmVdRoPw6tO0RT02p5/rfAOtM8rQaeuGM
N/TM+je821jQix80lByb9ucH5y93IJlFRpbJpHrQ5yBFNztYp11t7c/HTUNgc9tcgYlWJLZ9z2Ot
v5Qp8OqBXHT2OKBnfOC9uoT+9IL/7uiLsPsd92YYqgZ+rBBQ+3Lz14nNqrnrI6/55WNa9p21/W5q
sN96bMFa2qpxAoBZOh2xi31pxd00urMenixlf+0bxT1Wk09xk3RMWr9+MpMxJlH4nVixI+h+v2Fz
NarbedDPOsDS2jvy9i9zRWpOXUzgdBWbN1D7A9hozwc5LbMz89uTvBH47MuGjbxavh6BbN8i7DdC
QiEcn5FOUaC3nMHk/jICHvYpaGcj6oAxeLoRvhHvJrUXghCKb5wdqpNg8ZEgkRV6JTh7Mo99RF5T
v/LwCcsuGVqAm3lkbTJxxERUjo7qEa+zxy9DomHhWivulw8VfmUhUh4Ufo0M+APSevgKAnpRPJOz
De9uR/7ayBppzDIlC1p52nOrIMeZA0aOMUxG/LkVa3g5f09UkqpqAeyhIHlwaXYFSE/obt1R7R9R
td+z9SG1ZSEU11p+6L/3NY5Tr3beeKfyMNSG9T5AHwC0AWA4EiZ1MwCwG/A4tBmYLck8kdNHQNM9
AcDYC+ct+3slN5Szy8YQ/wkCX107rKZUyofbUU6wynS1/pPV1DfAKC9bjRpW3ykJxQ6mTfbAtxJM
rI2hWqtUWFEIFofgN5Ns1RdeBL/d0YfFWCqVjBA+HoM4OwpS56jTUfVnzwCEoQrjW1fNMa7ikN/1
hGkaiIIz6XMBzSv+S8Fb5D7IQaQEgdW7ecKZx8twju+89qnvIiTA4aWyzv5G9qS76hHMul7aSJHy
1+jNMWBvuSZajTfsW8FovWziKqwq9f9YcDBCDGL82dHFQc7e8Ocu7mdRvv+3HGRt+1f2I6iJsY8a
3AgOiA/nKkoDShmpTv24VkXZ4un2CK3PpglnNIxoSmvW0jw0Hi2NX01b8aI88vrOPqIIa3FNv8Ah
QnHUhwSIucZK9DFGN5YkWCceslkAC/hXWA2zCQdrstmiXhZrItIm9O/gxRZ1h8yeoeKrxLvxRRAF
5eD9WT6bDpaPPYdhjwr+qFo9ek0hZEiaM4RfxclN370XMjCJWa6dglfKZkmKZL3CfcYDrtcIp9W+
yCdN+z6cPJ+4vCLg3RzZUK8phoshJyV4959fLXPKrEVBKQiXt3WNCqU4F6X4twlgmLZondXIhqvu
5dbUuAhywOoJPKn05HqXogUItK2DVsZeZWURow3fqIwRJVAOZKXf6IUWOYNDqi+OKD0aaC5pYapE
1Ee9CAu6vOeVCUS+dEVeBQ65qhSQxi6BL5Y2H4PTZYUueRzeQX9TIs6hX7iUDW0plbyYW8epfX7H
Dz5wNIUsnN6rrZV0C91UDP7YClShyd8SleD6/Q4XGiYt0N5j7Wr/cFF1AYxyPsxdENUnn4rrESeC
fXO+PWdhBRK+sf2A01nPK+mTvzp4ZOoSwuKkow4eqkY64CQ5DfLW3qF12zsKRK/iZC1mVaCpi6oA
6k2meadB5am7gpYyZLd3zEInk4kXaBd2yAEiSx2oBKpo76gH0RJ+ol9d6cNm3ga8zrbgS8KzKMSv
e2ZD1/7aQT8xDSu0WipnBML7HwhT+LgwpKKtY7qSzyg8Z1xewiggJFofEkRqnJZlX3fJvIqPiRbl
WAcJGwnZxQmba2djigV0Vtfci0SHuVxlWZKNsRZNqobPPFfVZg4MbfEdgFdrCwlDaG9rO/zt1qt4
jYd9lyADMywq4KHQAz96VMVg957c80DxZR9U3R9yEJ57C7ONql3WYLSm221jnxLm5T3EtuZQH47S
PsYb9IrHT3CvU0TXXq8tm3tjdTGAyihvvehr8VTByenvC2smDuFFUl3EFSxqKnifVxMxnJphr6Ow
97dGBTzx1FiAcYLHNFAasI37kg0Lm12BL976eybmtuZrG0XS970G5PX5p4QdWTM7uG/O1KUXiJKy
hNixay1rq86afRFwmmxLfiZRu5so2McBnScTjgB6ZqUgAWvXwTYOVDzTe9UzwfpVR3+oV4a8ZA+A
e9LeKuXKXUC2pXX5VgipDlskHx0EcbZWHgbM+aU/C1tpEkS3w8Hl74nU2so/9BOLjhlxr1YMpX0q
e51JYwI3FcHQ2Z9CwHpaRhDLjN/7jrELE1obSMwUeOhDsEBqrTD6mRBgJfN1CD1txZbJ3YQYQ+f3
/p/3CxGt7TDcTrp4u02MV4agMVTfoeg7tSHmTrluDRBKvkp6CdhLfWIIZoZr6FyyDhH/fx6I6WIe
KakJkuA1C1T2Apwb9FBDU+Y6LVuC+NzKt995Q2dwssbCRvmJII6kCLXOZBAWNk88PYck16PvPdCK
TZv+QyhqIgDY0+W5XvxIF+CMYAK7QEOHrDj15ZswE8oiSDTGOtljGPa11nfpNqVSNbQ0QWoelZko
MTp/Jjix4LrHFHL2X0HgGeiwcmmzND3ar/enCavOncNuka/FQ7iyrP8UUShgONX+EztlF4J4r2pv
QKRVX60uCXAxZozieCJWBzSJgr81xxn8aCYjHEVT98ZX3B1sgV4io/622sT/aMKvyBW+mWNryiwC
icuLYLRQi6wQtw6sU6OihG1RsNf3sxsI2VUmhos/SoGuihwsf+aij18IZFKFXUZzWA93aHHP62Ux
oE08M2F6u4P393loUOcP3Ffvca8tBc6XLpkymzbIAuoyUPwPvbTr8nhGfIsDd6MMYo6y3szz7KWO
EYXdvEXKAPUYPSkyZU7ijEviuEfxZLNFbQP+MqM6gC7TxeGn4OX0vfmOdvplpmCTFnzaHC5ZVAVC
6Rpjo+82D3psKlco0lKmceyM0jfb4cosOY/cKQcE7Yx5LqHoLyj4j1pq+AcWdiHJ3iUG0LnPyKrH
ys3u/ks7aCbbdo+RzZCCSSh8H/JK+6I1PIIPhZACVJn1RIWqxboHItCssnsqwNGO8VYL/K8TxRhg
nDymNGefuICJUQjrfQ2hp2WkR3AOHICI6YuigntcgnB1QCmq1A//c6B0KC1g9adhDGkffDPiMN5J
JmvMaHNvAs+KqmSiiqV5Qb7zYNIoc8fwAeVIG5WKF7T3BqXwxzJkPa5iZISg25xVm6RecYCw59lC
1x1tXdg32ld97/WupzXt0XdZXa41jCgoxaF9AAunkvBuCk9rEnYi0WdHlAKTnwSAR27bV/kaCAs5
7nmKqOESLOMXNkFUyksAhCPxXjPXoHJSxewTOgbE7UlXGGQGrFktNT01dFD2fFodxBx7oKJRgyac
snhU93tW3iAFtt4Wk8kCqCxSIWhrvxQrs6BVAQTpIRVm2eDZevDmZO86CQAC5Q5svloJv2gwXQUA
ILaoJSVYbd6hvYCrOgVeDJEbI4M0xhHCTxiUBMOU6cvebbmi1SpRh+QSmubxPAXQZja1FgCSDXMI
KKxW4V9eIZn9slrVgZ3puio1uxwOQSoIgs/DII7gIq6hWdvXmdzXycymp7WwZSp6H3iuibKwJQZd
jNygA42kns2NzkbfmwMZ8wluM56+eWl45FuUQrh3QQx6QseA4CzlL2baQ/ygsKp142c6ekNANFOR
jOJqYx5VruhCR4uFnjP5t/7iDc8oAt0uIISVl0koByDud2hLUi4ACPII0XSF/5rTyVehvtozUpwh
+z+gBY5Nh1XPSOQM1TO1hnhMDzGYljwgLXel89oI8EfBXN6j1MfF3Qknajk2ND8N0+DP075YUYPk
PyRMasT1RISP9uYbGZj+jeGNir88pJ872Ot99hvJCNxX7ygkXCiyQO8e2lcWSBvYt5tP3Fqts5x0
tjrIck57CPNlUYCSMlaDVVWoYPq2kUn9OKqB2adqvd4zv+wlPbAP/qMDbM75NbvHPwrqib2hgywc
o5tsHifj8ATiXAnu+ckBE4ntzjU+n4Hr1eaVZ5MnLjUxAyvJzfXCrG01l/zaFLGOm5JLQA1Cy9VY
RvK5NzJ+Sdh0KhnWGjhJKaC6CsOpp7bVBf08GjIh2LAEKY9sbKbQFG9Mz2iyAJrbXQKlGLb6nQfg
RDlaH6jegrxyDdvjXeh71ib7HuhKl5JKD/CSpyQ0leT1t2MF8MB/Dl0r5g+iFYb33U98vVkkQV73
ztcM4zZkElm8PjMajxo+TX7UwRnUXeQfpsZ7L6c2XT711oCc5RFv95JOTUh4BNUPf5HKpPFbwDU8
4EcmRAyO2XskpQQBZxl+QtH1qQaWw5q9tr5P4cXlkG8IkdyTGfqblifplCx1iaCbFof94sNi/LvO
02d96gJ/quiC7oI2Wf4BWE1BsCfZNF7sI1hBVyq2UcXwrT9NmG1nM4RyjP3ffgIOb2hlTPHbiIvZ
C/jwBBh+r0HPW8ho6M/zsq7mRjH+zdVODbsdRESVo548X6pHRKce9szYOamVeSqfso9YxdzT9MBb
OgJ/Ky8DgdUo3LYL8Eby4n7hnIBr5VE8Q6P+T/uMPgxTPAN+SYJ9GddKTBe5pBX4+/JSIQnRF7Zv
r6321bZOGsk321xpgZai3IaIJT0Xni0aPVYjgh4m4RSntk6wGOK9XlKgqbifYCFMQmsx9o77GfLI
/UjCmJ+M/jEsHXfDTbMnQwjOdmFCn6/ImZ4BXFZEizNvHkwhr/dgw6lz8ob1ajpUOmhS/QIU77sd
aEe97LCSnF5FlQ0nBxGojIL/l040Z7shnd7UJfenGceeuGkc/jOI5/9/4ZP+30RQoJDGLFS76w6V
9CrPb/zJJApKUbDit5KSKFiOr+2wDkESVxxIybODiglUQs4qB0UUQ8TkMqT3movA0ebv2PXfoNit
sfLdfXk4h7P9NAGDIGgiRueZ6Qg++PB27t0xeXNU4El2d6yHvXlgLAIPQv/HYWc1vfjXovEWhiCo
axxphONyv2q9LZSW7GY1HcWFTV5e52/pn/+mCchQBMMVIsZnc1OD/Okx5KvMssmQCIoYqJKMpbxj
0GlfKyIdGAa9soawhG2PUeTk+qWzodjFzzxiahnDzG/dgTIONkXaemdoOlwNBJ539BZzxaLkP7N5
okolLmjA40DdKVeVdTO+BAjYh9J+oKPMBnAegntxnp64Vb6YdUEIf4G60k7jxN8DN/C51yZcciv9
OOl5iNlthwpGV4su+rQ2lquNzIjrrFQRgd74n1G1aXDUmNzIEe7f2pDEnay4zax9Z5doYWqBw3O7
1nf5FTLbXXdc3djqGrNTFTyAxE21EaHWGM+oQ6Nqzf+iy/zj7DqBmVxa2MfshtH+267eH1yGhYxc
QZAkJjXUxlcoPDhpvOUUDR78Zqhi4Y8gUSmgc0fr057aJgDVJ6cxVnOAv3nGijISUMq/oZZob4nB
m5tFFQP/RX1EIggTLoJQhqT5eEdUTNkncNAAnkwNR1ayBEu8iW+8exYQyO8EdXKkuI0c71QPa76q
ljn4kr4ORe8M28Bs+Krt6shnCqd0vRAnn3CYtI3ZkDevS1FHAGIyp9LYVA+o0jan+6y5TJsfx9VQ
2dwF1D/7wU9UtBrlMcHHS7MKjJ/NG1/93V7XW2EFkG0zfJQd6MwGOYxCAoYRP4wQ8Ei4KfEcEUQg
49pnK8XFkFFf3IgxjOIzZQ3QVR2/824K2/mCDnvEUkHafTZcfYlUYsCcJrY/2zkHSDBQSDxlLOmm
DvqM6Y/4zs5Gkc5iEQoKZI1SCvKZnsluhayQWjENRaE9RPxXOPptVcP7mmJzj8uMB5IPLYA39gb2
0eaMQBfZyI0izsTwAT1NCW5fhgTmWWMhuaQ9YtZirqAFh7JKpg+peXHwfY0sQJp4C99hn0Ko/ruz
cweFkrv9O6wO7KJ9/qA1Plpa4MBNN11hPaYGfco1tOoly7x505lJYLpODGqqfL8ZOLiCkOeZQuzW
sTqg/PqbrSYcEa3fXnRMRY1wuaq3IzynB2CmiIjW2rcPT+815gFduGJB7g2Bp38OiwAi75jvJoG+
nhqYm5q5I14CCkiIAeq9t+rh9ey+AxTshLgagCEx4M+uFktIIuv12J/hS7WeSqRg8zydCPjjC9we
xRMxxOtKb+mFldp0QHzR7MO79f+AwzH8X8aDJA2L4zSVv8cyrHt243852rPyRgh2jr/ByFjhMNuO
mL2EjwngkxtXD9oqNSYOCD0MoSMkOWlUoVL8W+rMI9VIlTUNtQSr9nojcc+Ukm8aOwJ9q/Ielwsz
jX/9X+fXiP3E+taBKK01g4MK722ZsMhFt8BuOzFH43zMEP+lj4BnTlFB4mTXlRExxA5XlVcBgh5i
LmaF+QvrJ22WREeATE4y8zznH/lU6PQlbxUl5jpNpXT2OQZmz4vjrp7BrTpTNdHlkWRt+WV8mAuo
FCBJhMkSxZgUNtlEJwSaZbDryYT1aAHamwz/cXc214SY5OJ53pvk6SYNSSKZp7GdfA7k9rVhreZH
2V29HFuD4KXMAeFM/+EA9VNIuBytp1fYMUOMBM2hrjZeH5co9Fe1ebch2yEKgg4bq40dU0+/oVC/
dMS6887TqgZ4vbfTp35YzzY5lzmTihRR1f9ZqCVZmZt8pijvxCxiBnbOhvff8JnNe0fWoE9cPTnx
058B+0aYo9hk7JbY934jswlXgz8PzIOs/qoQVSyY42UkoIeVgYy5i0PeyYevph0JpypXTkrEQSF/
wbAZsi1GKDoWlqp5aF+obwHZaii4NRDrYx1Yo5ozNHtHegGSuTA/WHQ2umkkIcNu4qgQzlR2fldO
hVCBQophvXHb2Mnu6TjgKC9z3C/zIOszyXGcug/b7z5JJ2bKAdq+ZKC9t4FB1YakoaARpqJhPNpP
vq9NW8+qT/wlWezLhKpX3Oxt+x7DmjjjGzlmoIJBnTFcikbmPTHTjXVOLMsbamfOEIJ7wzMuM8Z/
RQun0FsRcZ1JESKyK1ZtorWn1Mdh1RfPNgrMq1AyvHyBbLoPk7ykI9kJP+Y4AOhaN+qeXsuGmGbJ
jVL+H8nWNYx2E3nMX+fE2yiH6TE8O/4sH4sg3mD2zpuZyzmZ+0Va7EoEwkYXDrjKBuwPnzvXvfp5
EmKpPp3j2wCrm3FnG5CzzdV3Iy+3/00OVdbuMcSwOUwfggbesdZCRfOzQ5xtBcf7Z86wkSKvHrB1
ENLtODtqZ0siX4QsHxSXy1KexYxVrBZSlU+lwdP334DKrM0vudUfqa5VmsPHrRlRnsgMqT1ssLuN
qEDEgzQs3nCSeHIi64hdboYJt83KCsCl27CxtFp3rSeEpAqDfHwm3wWtY5HHtGvedTj+qoPM8auc
rZZvxrrDx6a0hKRa0l7047D+b5sVjltWt3onCQOh/uufFAqQaxKeADr4OIKZVBG6g2+QPSYE1QJ+
3NgRl8q2RTZ55VNuyPMoFKd2uZIgtD468D0SgdOreq19WC9gZZ4px7awEwDQv4/rxtZMmr+EDOnS
ajOAaAshAbUDuFq0TtwquvBidOIdDBbuxbGdpHvYnJVBjI/ZKkAu+f5oxfDebGhsqrX8j3y4nHt9
nw3jl/gqxwt2qn2L79UVawASmu5STZPMAQpHqjmTddXkXIvbwyhUm256Nnmh4n8U5brdkcCFRcZ8
bZDV4G1cSpZ781+L4aQMsn5IaETmeIeR1gf9liVX0y8JmR750DGjg4GUABGaTMuYBDvb6rj74brd
8Yxna3uoEuvaHgmca38mLf4ekVtJ/kM+8P7xjSrppvbe2GbuDelRH2mCHGxutR01M27DsMGlkdIJ
hLV4APudZc3r9u4PvNmFkD1xJMUmsyeLm3REG9BzuiLyxSl66obmfQze9hlVgS5Ir3DB4/GKWwtM
gY+/QOGo7tpdKloLC13wAvsS8ui0ajEV3q46QJaHA33qTWuGsmxcufY0vpR7QllXEQM3oT7+UgiW
D7XdCqEfVkTjXdGsngrxfSgZbKBfuc0+6odpbNS+fU0NuMZivUx1A7MT+zec9t5upl5JnfSUiYZp
I93xJ0eklOVd//oQihYW3dijijVX+At0Wp/3fA5NRie82ab1GkZpmdluggq4TUHIfOrZ/xYIsez+
B6zfOIU+LCOEa9uv5hYdIZK9w1edrSMXE3y4WqmwniGHG7bMRAg1UTm0O2Voul2wg3vY3+yX/Xf+
HPCtfr8MAoboewDGSBHNLbNwk4eTWNvenPetH2Ut+kWWdMxs8PJYhO1phDV+ThP1C/WdNxkqAZVg
jbkmRfSbgMlFj5z3VkA2sxSj/u5jfD7h3mkkJdgviKKjC4FJ5gVPv8cR6BUz/ard9tr+6Xj+Euj7
JSdxyq4TvYdv29At7ThNgubNGwVlSi2zQl432364uMcpDgi2iPESIaEPaM6tuAtkgodRTEx5kaFw
aMArnGrBDAnv8ACsb91KKDPnCb1atSD+Xjb7hdZ8pFlAoKccmEzsOl6o9zRvT8h+d22KI6bVqwgc
pracb9pgdYe+gaa/LLTh4uRLU+lrVHN0y0zhtnRhELqG/GEa6qzrXhpNnegjqvawRnlQeeN+BtS5
KvBDVcMMOMBlNExK618mImzu0Gh2PAP5+usQe+qxBA7dTklI2Y02wJ6Nnv6Xw4pqKStlkTt4ji+j
UCf6a/CoJznrv3fRPPlBn1cyniADuRDEVQuSzP279CoIflXARzCYbO6+fdFI2itR+Tp5zukdzw6z
XgbSi1WLYv6n7i0h85s4gU9pWuS+J2h+abaycQ2zGXE4iXjLQzZs6keyDbdGMrf4eJihoAcm+kyG
PlcnFZlmlBXPfYef++sEN47gd2Kox+bNq87qDIdeobRIrmFNr+NQsvmcXBe6UbEGuaqCBcMRUhL9
fEF+88I1AmIGyyGT5tlefAN0U5gjZ3WFrBNxzadGdiprs5D5ZLazDV8rZGWj0xfg+SwAD34EdnES
IMAflgCa6Ix0o1r0Y/t8ElBN/kBv3yHjWDKkV2K4FRu+BhLK1yqonrfCcWRB6eY7vd+bXcPFxtrt
ndrac6vjPKxOpI8dMkgcfYrtaSCf16honlHRKgaZpAYtDYwrLpMHkMrFAelCWbnU/2mC3APPNAHu
j/eK07LOn8h5n9JDZMicI34h2YZ95+OGUCW6wceveZIrjAP/Lxcp222zEhyK5nZby3nP8o1QzMjZ
mIbZMyZphxYuiEBUR9LM42VWSwRlCegt/P4++g4ZAkS8IcTVPlhmVPNrX9Q3rimHLvaBWptNkMiO
wWkF08jha5C0z2ZR/RXiDR9dzCiV30lmX1KNp5Jcg0v5EUvLT9aR4wM2Jeri0AmV+ukJzsc64GvS
UamnCvMAJn70YZ63+H0tYcQg3uWE+qco0iwkIETx9KPo3lkmqWefsyHlLDch7WX8Yfb1GMe4BBbI
xzAuTEASgI2JJQGI5r5rM19EeJ55AHfCoqJsqaJx5vl2gXvhnn4W7GvgU2xLelEbYHuH92UsYNEk
es4HzEZa/W3kzVSvOo/UViFF+5ifQzTsHnC7pOxw/O5BM5ToF/pNl1EGlFlxysE3Erz8Ppa6QqLE
ksK69sasX5btmf1Z1Hi36cXz+Tn4gJuLHf1igRAdiVL3bkiQ3Frb4zrPlQKdcEK+uOI1PGMaTPJP
hLJurSmzkagbYvknUEwJ07jlagLVJHQ2v+igYyfg6xWnTrEgwyWzOpluonq3dFRlV7NvCP3541qu
R093xOTW+WaVjjWGfy4ZIGGZVwK1+CwZAJbqMr/IY1dGxHLUcp2rhQaIB2d7L6/7rG49KmrSWI87
qYiZJEYU5f5d08VF2ISR7CGpERm+7d59CQ35tr/ii0P/dpVAFefJox3a996X5FIGTQ73xB3GoGl/
7eyidkGAyuyB9TZ/XA+AjMs3Z/NdvjOB4WYwKGz/7jxgcYhBzdkcBfXTgNWhJCXz5GnTK5pOUzdb
OIZcBEQImrIHRdJjFxaxhCLO6rqQ48FFatWqlHM7E9I9k5S901KPyHY41XbHhUY0+H5eKMdJYH2s
rtRtf/gykdKCqtIjcvj348vko8Bd6DG1MTU8/VZ5E3WVw30z0azKU5/1KCr3oqIjk4tUaawemBqK
YHloeOzEIEbTLp7EXzn+l0uxRNWH5ZjIKu3ww8Qv6VR/KUYQz44oqgfoP5ydJPSTNniV0rzQwadt
NBXnvWD4b1ectg9tYr1HJcFj4h0uf7KPh5iNqbAk7k4RJGWJIGX/Uj9XoJKAugKkYTM4Nxfshi/2
vqOM4cZ9GCZqD3jeqeKvUzVBcKT7SiMBrfS7TViQ0HiYro6yhnCilHfRkvtQ+liiZR1AJ9bjeU7Z
sl2N7DorUZ6hMwuHe0sI7eMFbS8DT4fyT9iWB5LP7UHhIs08LaQKiyTsU2bGIEm6/yz3nSgt+G1S
sfc0RwvtQK/0sAQEV0XSjd1r3k0ojd6yZm+zXvwAcLTZwGMyl33vYWDbKuTsuz1v/pdUmPGzQOpa
LWt54xLqP8IZFlEXQZVX0Eo2cDnAOBK1RXNh2Patrwnq2nfqaIfvvfmNgJAyJhAooMfR+UDM1/Uc
V4lFwkjxUoU+4ChmkMYiSagU31UELp9SzfljPadeMtXs76C3pmS6j0Citc8GLsG+3nJGvoaQbJzw
GObUP+9Anm7qy9ZQaiv/2nKK1WxJ2xhVxqtxzJxz+UPKRqSEXJ6ohxFnHZo+QQ1mPUhoaMw2IYG0
/Am93oWjWkkstLgVjM/oJq2HjzJrjWiDteRTxFEizVuOmFl+AonjFCOb1dEQ4A0NEM+85WPJ/Q1+
wsMHUI6T8dKL6Pt7yqGFfFP44yBaaxP6ztqweMrWwsfE9Ni9/ecr5QJKbTItXXaEZmGE3Xtw+TWF
4T9lRUGLfsh5V7SmdMOtO2JaWTqjs47XcAr7i15guNRTwDFhvgYCuxyormu/Ga7LL5hfUBxpDjwZ
pN+s+6LtombG5DUcvHszi+BilQiYb/41hQf5EXY9H1zIujiYCa6IguC6OfVKuNUQBqpvRnBivqTc
jDDDUsHjs4t9vaEWiO/ye4MUGXTq1XtOeiaynHcPxusv5Er0pXkMrLBX9fvU7DoBU1ou/AI8Bckv
gl484X5Py+EU8kwYexdKgZwQA83W7kG5k9wrB5wtF/QZRdYZmyWJCqHuNTeOFBt0q1vinHTFYlLV
zr3epr8ixxPKTxLvlAN7Fh+SGDxvMDCliqZHzg92UJSQ2uK86JM9WsURncxPgpxzbxrqM1AibxXZ
NGt4aZXKE+a7h6FMn7dcmBtwWU/vjZxC6XSsnQu7vloWjvXKvl7hCBvZbkc/S06CPozwb+Szmz2s
k243+IpQeWSKH+rzdMRTx05wVUWF9ZemuQZqiTAM3/P/Tp1G3T/t3IEBimE7rDBuZwa5Er3OV9bD
+7c+0ofUXVSLNwS0pGVTW9g2I/ScEiClqQ+QAh0Qpyd00Npv9axsVLLzTgxWef/y+fP8H0aLqOdC
1GJLvgyb31qLZANPVxr9qFlOuNDRO77GcTxw7wVcm/rx3QOR7j6KJhc0i7dSsM4EK7WxXksQBcmY
NBf3/eYkXmHTxX3+hB9X85ei9DBYi4n55d+ATwe4e0ZwHHqXo8Y2ZsH0BUTl07oIV3dXn/18X05P
95miaLOJLHX9YerqjUiyUVvZsoZ9H2GJKe4K34xwzvvmdLHb8NTTL8yNnDXRxj742A8GyAhQGE/5
2eRXxeTZdv6tiE/+V4t61SL740LgTJxHjoCzP3jJWjPqtkwAf3b4YzTH8j54enK2TiymyC3nkVEg
s9otVApMXKFznn+9mvfawNnfWq849AkNGqE/etNSgh2Sjy7b5q9XZlvfEBmTgVJPMjW7cioROSET
S33936IrzhsYTifqWqOdZChspTThuRTwo9hSR7pXHkb4beZmen6dooKp3GoqK0tzTf8GG4vHI1sX
VF/NApcoS7ZJx3qQqm56LsOQF4DZ1z3Jejhao+gKokIFga441sIWBdaTfx3zZK8hebIwxLqkJBvi
IyqXqmYQVeVawLze2+ikao1buudQ8p6/2CFX/bIH4oM0A3s16UHV7gOE8rqTKNNke1Fhf17VNDv1
fPF7g/rrZQDOZtVNm1zz3HaAnVN4fxCwKzo27tnmxob6Gu4huNEC7I1AMxX7rJHL2wvLOH7tYAb3
4u/+WAyCFjH/ykpSopUEV0LxlKp1RElydoN83F6QyxzyW8H4/DnT0izETLfM4U9BXOuqz2QCWSNk
bIGdDGRSedF8UOg7sPqEQ7/8b1QHAUI7WovGsGwS4cRxI1g+Y/HmzwJ77cIZLrsLSXq7Rboc0ItW
JtFZcVunxpNUC7XKe1U69pMdWfGatjknstvkxIwd+cjToM9rOcyUSXS8c1MhwhPxJHhscazs/KV/
a+IAeEJTyGpZqUYFRLlj9x2OSpA2KpNtATlDukamOI+OJ6cTTF39Jgt460u3oLADYiSZaX61tw6y
Vqg/gxZlsjHFCXpEg/Vvk6BDYi92T4/u7g81phRKp3yyA18oVQp9IkHwhv+k8WQHJxu3kbbCcyWN
AluX0T7BuCaWcht5OMgf1NW/OynHBJARoeTswAeVHmpovxtKzholzE/GeBDH0/JFrdVrS7cJfgng
FHeclP+1Bf5Y5TJa9/ZsVAvlGfaZvkytjeSU1GJXOMw9Be4IHOr+3p7qShEiGfES62ER32ZhZUV8
zxrQvPaApR4sXi9g/iuLzKgJERUUi32GJBWBt6fXuLvxp15mA8G3XsaL9LFD7e0C+I6EA75fN7w8
ju40CeVq5wcWO0jLW5zdYPV+bkWxapUqfVjguKOO7eS/2GDSjmjkvCR3o5jQMDvxwogwe7xBk9fa
6+GXa7nc12qnMWJ88gc6rR56u1862aLrQanGSb9tGUyxLKbTSFMVA05gGswqsq9dnWMzFCfU09mk
bcexbY/iRHQHwbIqn/hPzlympEY3n7U0BxfymaxUwjiYRX6U2ApCbmceBLEP+WLXvHOZJgtn49IZ
0XnLuG4RsLvHACsdyRRaCvB4kEnmMuEHmyjfOnmfXJBtR/v8u8VRB+h7spDPUUbWbx2GkwnrFr4/
xZjY97IoxxK6BGWh/VZhVnV4eDIgWBQci/bq6k4MxMqQIoLsMTPJCO6k/cYrAvUw0e160o4iYxfu
wDf5+TsGj2tsAoy2hWUs2F/yTJIxNEZMNX8onnG8VUVaXvSKk6MNcGg9YUF+WShuIH+J3BV7zkR/
PyhCcUIiBa0DC/m3vGtWJ3JQ1FzXL2SA2xfPZOvBHj6l1j+ootQMjnk6XTohTc4nu5SWnQ5bESqC
e7hm2FJA+DyfiQ8M119lrK6icVH8fo2nuNIKHIHlKRpaLcRfQHeAMRMEyMwh8FiHrU/YewrvRBJd
J8T1a8W4vBsAHXBVHlRlIXDLOTzw5bff78kFb37Jpk3BGaUCoJ1N3YCHY7j6h1VRSshFXatiDIuC
iUFJx/Ah/+JwXFs2Vvw1FFe2bdlQGZG9cOTkEASKqWzvQwCJRsobD/IugrQCi9cQ2y4kxsVvPwGO
FkdqOflLSuOs7rgurFqt7msacduTb5ZVxhpEytKT4r+7NUVBl05/NKqEC65jaYTiG795QzoIjlIy
wG2+ek6JzRr/3tEGki0Fv059vvC6xWSYkbFh619reQGJHRyW1S67FsyBGIna+c/2Jq+WDEpMGY49
yOzjQHGvBHDTKB+R7ZKiQJaz2GR7P/1ZxXenrzYIbyYladZLwlOJsvTimR2qYWUErBGin5D2UgNR
QTGQUa+2JVN2XN5O4otQmGZEtymjoCiM/Nbiw2K/gEqVNKTTvHZllu56QFP0M9IILBNKxjrAJyOa
4s6OQNWtJ5gG7eZPy1f1udfTAfdlYoTW8BTeEdMreBmtQf7FCIgwP8TUr4AQTxfizwNIFFlE4RDT
WycSw4VgTTgl++eHrUQnDvJRmdZhnyiKg9rzIdfw+xBsxmcswAY+90XQ3F2GenxQqLa41kffOT5W
EotA+CNiTVr9g5a/ydbZFd6JlwF4UXbP8yy7/AdHG6cd3vG1ZXRXL75v7RkRVjybgXtGCl49BlRy
9y5ui5r4AZ9luIuH6kwwENFkEg5NjF+IEB+5UOdo4EGOH7XISAy/e7JQY94pZZhX9biGDW0T4+lz
tZ7zbNDDR60xu8Ucbbe5AbVEPn1OdLP3Vj83oTiQDAV19bnur/lJ20hExMI8v/u9VgcQyk/KywPl
3DK3ewJhuTrddfXp+/+O+tbJfZ4exzVTOfIaLdm27T6wM2ozyzBBHoquf+n2KZxjqEjW7BwQhXYr
1Og1KmHU9dAyRWmghk0NoslusH4x1O+mp/ILV8Q0Yk4ARXV+LpCqC2+6V7LxKJdDBeAFB7UXHTMc
NjfEIT0rkZjUu2aHMTFu9lYQdGwEO9DaJ9ze2Jf0qLAB71MIuFJcZauH+1toz+2W3HymXogtl/HE
/K9Pw1Cr+dWJxOoeR2+zIEoljp+6XbT0t6WdvZ0o9WddWlgbmc6oUiAsVm6u8vyQ7FzbVdpS1Pl9
uQ18wfZmnMWvI96fPe9ejhWb14gFYi0lQJh7G2rXUYlt78HyXXCrIqlgmvbYkoFj4RbMRVaw3/43
MyLWbL3bwpDTWyInd8LIn719n3L0UYB3FVAyy8QRJC6VSPl7URGQ/RWTZEMcqlxXfTfelKWnyJ7L
lF6jbwXjgSvkkAA0zI2Z3SZO2f8dZJCjXi9rHf8NPFe45FreJ6S1gSZcCwCKbc/nFLTHdBZ0QPlf
GrNw2IlXBw7AUeAkr7fu6uVW6l2YVdBCjLq23RAH8653FsmkSEAZotnrc6pzJy6zi8+YBgeIywae
t5FD5GhL0/+4F39u3J4oGDvSIT5Ec77oxGLaw9DOSW3MwP0Gg4bNtse6Vu8Tr/TOhSA4HlHSGlul
WDZrpm/nVw7YQaAlVs+i1o5x3YohdNb4Cca9NbTAtI1HDlLS22ZxyRwG2utqFXbQYgjzuf2lRWlw
c7ZnLksbvcNoUVsUSyIaZFrxleo8ucamPWrGcMRY0o16GeFmziO4nUVcPcsx201q3qijkc7baCHG
UC4u9gpZcsXOEWuRpr1IAHzTvDc+r9kJN08b1ZVfPFEAH1WiwbUEOFHwhyJRZerAwzebPNGdXocy
qOhZl13/QCnt7Oh6EpIjowhTttpELCT8R5fypxLi3Ps3XNxhMhf9SPTTrzJDbaRRoG8K2xdayD9Q
+N7Q0CIAYTFgQ9UODX2ZFq+/zQo9RGXsl2iesTT/HDNbcU4/IZxrir/EDuAkeITtR23KB2SSNmq8
5e50ilFEphOexbw+k9hwaytYxHmmmCKVqY6n/kIwykOFaPPiEH0xYgQba8PiS8iuj8lg1rvdI/pg
lJQWTfdFCZl956kNpIV6u+zkImzOHJp69QJGB4uRO51vk9jwwILS09BVtB4QxpM9bmLFKzw3EXp8
aH7rI3wW39vkWSvUibhbILNeu8z29gxaTU3DUS4JusalOoKWQwC7aqiOxZ9u20Slz6L3GaVxJAIc
jxduliHx1+GrM1gnxMNXuHiRKv0vy8sp+ryq/WThqr17spLHJ91poOAzHkXCvGTLjBngFHIxmg+1
/SxENCiwHErWRt6TBVpN+YFMyuDbylQjo0H4zIdpZAE3/zkKlDFfgqoQnOJVlojW53lQn2YP0vK0
aiV/0lo3b8m5xkxPEkJhCcJXLuUe0b6yIegZ0yNw+OxYcIL539OiGly2I7aOWIaKpWCGd+5d31in
PZMGgiFEw1eZhB2xg92ygBjZdkm8ZVjT05LxmvMxh85jggsymB1kw3C39hpCEqo489qsZy/cKXTe
9/cXQnY4Y+Y/TxlBCjKkzY7dsuiUxLB3snXTHnLApnogJeYqCCOW1GB+OE2FProOTi6ytbOcct73
fWHw0YerUgKXcjYGsQZq8Y6XNAF+AolHbQI0KS/aGALRI67UGilANlWL//nRy1aAIA8BA3jzMA7o
BEcQ4NyYbn2jHV7XTAcZYdbdgkGxE38ZMBIyhEzCSgpsdPYvyS7WGqFez+ARKXX/bvX4CXxxDiF9
FDrkXz8kzBJW9XU90qTFdjB1cSp3fgxKKZe1bILppMYLZFQn2ynXfKmkVOUlidVE63sYC2pLyzHA
vjcvGXzvutqU2U4YPddqs19BV8cL+e2YLMFBA2oj7ZCc3uCbm5AMSKbK7Kqldod0bD5Jcbs3z8VG
jWo/iWCWRG4IQhm3xWvz0e+2VlqRbFHDM+6/EgbU5ZHZaQ0tM5F4OOCCrinCREKT7tWu4wsSlWc9
9xF5ITq5XcFRGvIonwjsCmEEVGkVscWAXzNNllgRx9KdFWtRxsk/ncEu+eWzyvWgjd2o879eujh3
oTOkewdX9OQ7ST1DCcUxKFwpHq03EYX1/TXERZZ/JAEuFe0DBrbVHb4bHChqCGbl5n7H39CkEHJH
EOLSS6BF0d64UBfOAARFiaDjzHRVtnjpyQ/I2cbQ54VdVPNnAHwpegPj2asoD2akPYg2whU0dI14
0aF3EbJufRTlH7vyx/ajDJ6gryeocDubA8AyxY9hYrTxGbVlayfNUqoyhU0sXS/nJZ8JyCUFeH3G
wCNVuk6jHe2s2Hepp937kpmIyvfEcmCP35nBRzTFHtlkH2OCekRK7syIJ0TWyyM/E6k+Wei0amMC
5L39ny8tF+BRakWSn8tHHBbttv+qYWLVO7zdeL6oEs6e/zR0L2M8o60mUgFI8d6wJH3HsZN/BPM9
2YV4eyZPh5rC98s5LwrUAw4UKOvwvCKV82iYRJVzS6Styh9meplYbcHx6nTUGg90yRL09RAjaC2Z
tQn2MmGkLNwR82E7Kg51laDb8Q7gfSKXWTcJlXFaL9Th39ARRqCK6IkRKJKFhjSSn8BZZnki8YvV
92n6/EB++g9BMKrX0DKsbDmrNz4v2H+lQTsIRt+KZB20/8b278yj21beXe/TY+zcwlU/q6zuVQYw
9cYLxLrXleLQaTDnLMNS8MJV5nDe5DY90AoMshDYk9ISvP0nUd6p9Bv5GFcZ/BDgXnnyZavQY2KJ
7DXAiosZOwau26gMKu/VGmORactnx86n+4agUGtmpvUWx8E3OfP8T6kK9y1pmtC/NqwlPdv+PvZW
qCDacxXF47TneowkrTaGiccso21ww8/q3zVJ1txr4oX9oxaRt/yjNy6yV0cm+ZOEpXctPaK6LxqN
QjQ8i31dKTvFpr0k/LfFZ8YgZoNL4M5fIY+8vTUJ3bJ26+TYAUXQyi76DBojsgbgAbgbes5up+5y
IqzfWtVHXEiiQOxSLWJdTxKUvSRITxLhnEmXJ372p73QTTrT9c9mTh+zthG7GZK8gZCkX1OM2iz4
phMEHhaFLUCPUpeAUl8IpT1SNnYgz+bqzYMxt4DsuVqBgMVeeJVeIIK9VetiRU/3nquOA+Vcfr/D
wu2HBbSNpAUMKKP7MOmVI+IK32NC1b0kl5iAgsi1cA3qAbCgaUPCCf/gCHhIP1fQtcHmIvJOtYYq
A31vXtumQca7BKXZ/c88YwcrpjVWtXHPaqtIbCTzb3y4m6ZFLG8I5fUCWv8Zq9hPRmhcF2I+VxNL
zbOOP1+MwvZYIPp8s1n1Ujvmcv/SHhkeVEKdUMFeDXrdxFJaufRqysyt8GoHfTLBFc8LWmr0E164
KHSJsNB6t71nU8ydSkwdFyVNof+KG1mdE6eFcHMzPPDn53Riw4Qoqw0QiTjioL1I8a1fh7r5Bhdl
8UzqcpNqsgG0UK8yyVtRjU7x8ZwUsIhyJgGdUU2UKC0OF3b06oCK+GzhNMBMVzhDKkp2PmQrT9yc
QQKqDo0BD+FrHnEcwKyZmLcztGaGsh1EHGwYcyUqdNE2hNfXHvC0L29r5UTDcJhgRE+D3AjhVyD/
zSSz3TYAwIL7sTxZ0H0kC+/I7QzKe4kbgGX2nOyIbbhK9xuG4an2nlHD4KMH/TNfBCS5vZaq5dBl
j73Ug2RnfapatkYfYcScBFZUplxZL2JlRg+nCufjd7J2h1yeeRi/GIkHoWUbqW04JwVmT95LsGgS
DTkdLC27+C67ebApdeVi+yVYJr8M7oOBdH+OYZs5x5Zd8JoL1UAFI4QH2QHOAeAV32P1AMqtgnIo
kXSxw3ioo60FqH8Cp+ExuZYX+KzAuRdsr+shZftpPMdI4Q5W8TO7zl2U+3d82p+xOr8kR+IJMpv0
eIWOT651RH62ltp2O5Ck641MZSCFB0eTfw901VuJwBmPxq7J1tQDskIc+XBYwu6Vlfhi0s66urCU
50Z2zm3Okt+p5aK08EuAevoJyKXMjXO4lShAH7H+uywKPbW0t9YisGTU1BIdQdd6uFFbph3WS4xk
dcvwp0B4nfL4fTTYjscDNV323urfYWsBL+e61C7W/M3SEzrQNCPDYKMQFjx8eaWRNCmY+1Q2bjG4
aj7ILKurIfIDZMac8ZyYd7dlBE1DqOdqoefDqANAtil4VxdX3abes2yW7R5zrFSIdt9f/dhjljgT
kkZ2H8oGg6JSiSbmEXbtVJC7xfnyeHUPu6QzDrwYezKFhTapGAJdZ1gjtVO7MPYPptzBJpCu7SnY
lmf53uTeyHwm5BFwsKlvd8D6hNjNMsWiKJpxm42u2OeriOLnJmIBMi0+eGausHli2yV7EjjR4uZQ
uKzQpebQChBoRbILEYSwAm5s3aomAoolpDkJhubB12TNRRxrPGjxAAUgXIIhoU00oCjjLYuImVHW
RxsQ108N1eg73Jxwshud4IWY1x08SAJ3L+RHCeKbT/7O22TsBWpqP5m/JWSzhIjSozflKcm6vWo+
jYgPcKqh092SgwwRgP8FDJYVxbNuoJC4i5LPfdxhU+lXA5lVuJCWqfDSkACbC81SZ7mxkKJsTc+Y
59mIAvE63HL1DD5ayUKw391XcZCCDrEk0YLFfezGDn52T8DgzqBB36+URJhdYtR+MDh5xRrlxmtV
AZYCDNC5sUK2aTTNc/OBn3BDsxR4+QkxBcAw4PNu8WF5l2AYgCLP9gM9CtFL+CSdMdXDuhxiTM5y
k3PTEc+hTPnD5BVMprHcFvWQ0Eab84Dn1Kan+xRJalZLvrrAn8e1x8Z6/jXuJCS6CN0CESPR2GhA
QCelfuqhe3hQxqw3oMFTlIkKZ2p1dSqZiX7opl/dRg5LhOkGB81qcWftAJmZk5BmHs0nQiouUKDT
EkGqVK6XrJho+5o7axhTRhSpdOCywn1whgLbfO3dADF6Xf6KdCW0AG0h5ybuTL1ZPtdae0Q6bI9y
bZFizItpdUlbQ5CmuDcLEovzsdmf1hHepkI2Y82B83OO/y7MobiwUncXltHbjeGepkOsApeTrQIg
SxettJMN2Tcliu3iPCuWKLXOBmlp+Hf0Ds6ow2FO+Nkfv/ejULCDyoYSOpIMMauOL378MkH0TkzE
v6wC+Hsm1kQBCsfcYf+hSH+Rb4/1VTy4AopzaKnpJP41gBd7iEjNdUfP2ERiPBOWhhVIHuZWCQ0p
h/SkcTrHm3KPIRBkFy7A0tsrR8DMhsKy04QMesNiJ9o5TFfpf2bq0eJ7w/2ULnk/RUCOgIlhuWu2
4Q2aqLYioVdVCMOrji/6xb0ahIc2ltUgaYjJkfq3bXLJV7ZSfB8o0wTq3IJnYfRGksnZ8amt64Cd
lXcu+jGw5IFHVb6oPO77Gwm73j616g2sLemSeEZOKukGz2qABsw5Q9u3uN2Wz+wcscVcdzA68CXt
D12OEA3W9HQ0sYdEYTQNBUeadPj6nYnIiODkmr/vwq8T7HQQtUbGOpvHZlgm8QoaY4LqIXokFt/Z
CVxTyzlXtO07NCSIxwJcMLb4QSV8zzy8aO8GCLbjrcPKpcuRE1DMszXZF7wUUCSkohJSeLPJNE4/
JyaGfk9y3v72Lqgqy/Mmkf4WBwJjhWj4GtB9wK1pAJan+GgkmA0olfvTAthguf7vtOOi3jq7NaME
O3nw6pvuXRIQYmxCU2Hbs/WPmr44DJtBoaPF/tIa5EneuLUD/lltaQzhSsCjCyQeugTpvbbmFFL0
fuAp68hMWTOOAbQZ7O2V4nyWKXKTz59vvucRSH0kO5wX9AoP0xh7URPCF1qTU5M2EKS4fTm0x6QE
VqcH2nMBxIpmNZ7Uhl/+QTEIgRnkrdtPc5P7CArLakeIAvNzHun8RyTv8ccDqyH0tT0fUVzulBr8
RaR/S3XzxUPR5WJJ+Sh8Vj5evhfxhRvlxYjtcVwbOIbsKnUXqCLTXzBjKYSQWf5phW6h0DOSHVM7
fEUusMHWuLGON8futfiesV+dG2EKqEtNi1uugnqLW4czbtYBbP4W7iFskGOvjeyBP7ouRN9BiU8y
d7lPV6s74GEnKIJ45bOJzfCJi/saUnAvS9xvGmvMIgu0O8YinWEN77FLZdWoQngLe5PL4NuE+p5i
wJjoTe46FFW/0DmlEsvPMPsrBk9wodKw3gxQN3NxvI80i2Jr9sy0NVnivy1XniaSQiqnilNdTPNa
KPQgTAIWyMnlmSnMGuOvYS4WzNFyNp05i0luHR9+mnF1I7eNn1Qe2BkqzuaPBrqMonHPLMvWLrTB
+S+S6BuHkaUTMAjrkSNvZTADvV7rGpMUzYfJZ8h8fkeDNSmHuLl+j+sKHPyToFvYLcLW5/1eL2Xt
6kvcG5nZFH43K727manIhdlc3Nqy+hZyu/up4XUO1seglruw5bL1R34p+/7iTSpSvnudro2mJpTQ
MqDBACTlwDF2RApAslYrMMr4WihmSG14tV12DOgm2g5oCdVdsu9Eao0Y6ZHqN+qSTI7U2oPI3jd7
ZEwyE0EAQrPELm6YVmu5nfUVCtduBeb4cpW2S4YxMa0CkhspnhszHzWNFRMnrj1DRIjNxrDgUmBu
GG5KFfE3ffZVBuqa3CH0oJSLj4D8S26vzHm3QqPHM1nRO/q+Z3eK3AvATyX81UeSjxrcDkIhMw3n
1usznJ/8gFXKYtyO0U4scZGW3xyfen98oEzOKkxqpzZuZ6dmMePolHSaVxwTVXbK+BPavhbIz7Mi
I8s4cLYBafuFXw9QFMXNWwznwFexVmIuIJspcZ00jeIHQqRVOjbQRg/W/Bi0sKf08Hrd6Vgy3n3X
zCZb6LcsfpUpmI1AG8u3+mluXm71ziKLG/gIo3SQclu5I3agJDQGeRIvU/yAEJmGA4B6YMppxamO
tYPkhjC9Vx39CkwPwgQTSYrQG0zOU++xtqqQk9+EV+RzeTzzW2YM43ZT1M/SBnydlzXGoseeFISY
lPcuHlKEya/PrvKGoSvvHIvkBTxZw3K0J3VvgoIldjGSRCirAaPIQY6u723mNL4svKmt5AHYwhix
FfWAhpZupZqKA0U8qEVbjVR+9qQTKlGz0uQ0WWWEDjls/csSZ14+IWq2eFZUk2kjNO5Jlf4x+5fQ
4tCmfwgiALJqb5W71zz4u6Wm7yuQt5wVaj8HblRqSTSb6JM7UEFHhcNZGKSMdIWuZkLtyZa2Okl+
2J9Yup0mlEJfh89lSodo31EMqY1jvxhBU7I6AEg5tVi9uAp6skKbqxqwRirUZHw2CjEkBSdbZ9WG
1kb4f9dvv97deBoBcvDXiaBriwDsptQAybwndSwzh81Ae8SpPy/lgrgOxdpPn9d6LsROl7vYLa0M
51mafIsUC6Bc5hx54MtuKnDbPKvHDryfF5FV0cc+9170SQMOgy/Yhl84K9vD5F0T/9xKoBhy4cih
+7WkEyb8HuqtCJ18CuuusVnIG1edRhiGp2kr6P0s4tUSXjcLfoTBV+PnOOhviW+IxNRyzjGtZKEn
mwD3PYGXg89jhnKNt2Zcu3xSrCR0MvN/+vJx7xop56zn1EZs6xzM86IOCxaxX05KIGNeZmlyujRF
rsI60k9onz+6enJ8bxi4vJxRUX7a/N+dfwO9nj7qZGt5NVi7yNmHuwD/Mu7muqeQ7rLltFlPGmTv
eNWlynxGmMEO2E895t+AgZqAtBKyUiQo16WYxrV6NXOIUDyGgHJk4PoNm0BRsro7PqvUa00kZGse
oeLV4jxIk/ocT4PC7q3asJt2tgGqsghWLBN4TqKo49HuhFl2apUR0cIbiaQyd9yM0OGDqwEeLfu0
59wW3snS4EECKYqeg1soaHVp7VBSc6bu+vK5KYY45SpPG3PZBLe1iAXSLZ5A55zpbWCzdsap+Qet
Y6gUZSu/Kjo4O2tEy5hfn2c6adoWKo55Udr2BBep9WI+PmKZJwHT3uS7ms0qgf1O8nWZcGxyxxD4
AwYnHale9VlE/p18bPjBqJnsQyRAYPt4s04WmtY6NH5msCH7vCPhzx3UuVLV8uhGvB2PKVso7qGf
gklmPshfE2z5MD8/CDplGOhop6zNAY9wtyw2hK1Y+kDA5WvtlSw+kXZgtk+llK3bHYrxC54FmOzT
+ZkCIQa5pQtOKp1kn09JZUkbFzRGhE9CWszkjkrMkh8+ZdKoOrrz5myRHhCYO8Fhli1URVVkGGw7
T5GHWGVhcbeklRhcIItPLwJ6Gjxi0mw3gtqIFMHOvESjr7M/siyoYpjb4oHV0mIZvAff0G2s6csg
mdlt8v69eBFXCjoLiRsJpHxs1NCB8VaaZqWOZ3cnfxBagAT1Jpe2i5mRxmdpckunUJ07iJCq/KOL
VrknicS+bplixMCCSZJWh3VKxDYx8y+t/Sru1yMz5D0jQAa0bgye7YUqBR2pvygF9zzsSP0cH3Ic
js1mDNVYmCMyfYsbVX5dkVuIiMjBaPaCoHTVklXfuutJAQZa6ByQoH6i1PeyOE5c4UTMQFgzwuW/
DHbLaD41Wbvs7tpoMZ3b+INZ0mJ7fhoJvUZmTPlQMl6OLKVfsyoZqwTsGi9OfRfvLkAcIohjavtS
ITg/CW6mGfcrohY1T2gDjmKWBVQ9zmT1Ju5jNRqMnfld6H79GAtG8vfXQgTac7FFajHr+MExwUYC
1OowLnRMysF1ZfqZrzXCZYz6+O+nAdhiGK45Wq+HZmN4+5k2sY5/7T0gpAWlX+JgFmtrVs0Ez6ca
mCiHM+EorO37+CVI458FxNLJ08E4u0f1dTeCBAdvhcWCjTVMKKnAig5SaGPQRm4EI7BfXmpWaYc4
0sjaCrkU80IrjNV4kDzjGMsiKi1ApB2vgzjGpFJxDHbooLV0jXrG7vCBLNCB3b3TSyAE7eSJ8X5C
6dOhuC7Z0KV3Nkc46xwtJkrBrOJYPd7JGdyOW4EXlP4Be50iKEp5yzP2IZdcOimGImXkbGRwZoT9
K8DEVN3fkH+b9uP93JgodQJan5wMFjFAgaCtmoYNeFiUQPyRGcsc+UI17VgL3QenUNFvgucvPZ0n
ChpVK8v3yfq8kJxMnoCePHP74Zz0cbSyvnXkclUUKMBx39PQ0Fg+oBUrRwjIaLAbALMGJ2o9Yype
BZLCtti4+puB83TP3EBfBqhqtOZfSla5id1V9RBEbMgYCJPMsYsBaAv8mmntTFeAiWZ1d/7aQzL9
eusPsKU/tgwAoBF8lGHWaIXVS59JXVgVlVgsE+l2CdqFN33SeFcS5zzxdMJB7f8EimAcmyqoho3H
pI5vq0hVEWcDHMBX8Zi/c8Z62dj3xL2rDx0BgZKhXJW/B20JGF0M7y4JLFLhKXsejzO/kbp+DTwa
8imEDl3td0+4SR+HzK74uR4nOXNxzODD49D7kwZurRNUSh0iQpQDJ+DNaPQOX+RqVA1y1eFa7oah
BGFqqq+N65CXuD93EHbn01V6JpT/q/NEnUBw0H0QVE3DV5R/oCp4MS9yUJmbuto8aueD/yCp0hpZ
lYFt1AtdBeuVN5/1g8tot1506+p4W7KXHk1zSv6CdAumIQOzWhlkDfq4WbCHSpB0SAj2cd9HwtdQ
afv/OAjxhb2wORJdG+HZo8jqv6HZDTbzmljmww0554S5pgUOc7xH5aWyzNMsxZ6Psjk0SWR4Jead
D07pFRIFmlnMC3IO+mcb5YrzTzDicHNatS9u/g86sc0iwMk0U6CSk5FLSDrJ4wq68f7//+Vr2/Ki
A5kA3iFyv3osv2hFYxFEZ7PhtlYWc75mAA8Imqdtfq0i7ZC0Btg5fzTox/qW5lkL2jFw9quQ20il
3QbdPjmAyDTqg/wvHuptX7kSZI0SX2hOXOjZbteBAWqhdaAQXOVaR+xgr2+K8WpF8WK8D3QTT/92
sluxZzlAW3UThfiWAvJM7GsxnEhr20jOHJEDuIti0uLNMl3Hxh3pIV8b9ZzFxSpB1S9pMwC80vPx
KFNpwr1D/sVdGta4+Vb/PrNxCaCgL8YVUELZZscg93M0/zV95xCPAMR9UXStD88Mg1aNnRc92e5p
ZseolKmijZGu/4xmTj+mWL0/gqd36NoZ+UUKxf0nav4oADtkh5K4rjc0CBKpYM9ecGCcQe72u0G8
/yMZgUqX5Ui2j8A9sOmA3bdNHCJtjiO9Lhm/VqLjXe56XHn0wQu6JitTXoaVe/PJacZ23sob9X/q
Ey3ZDsM0VkQ6PAf+JCSiNsEvCnP+QtGTu+ure9robiBkTzIAlHAIGB9TYLdtq3Bxgy24UaW1JAJS
O1ridBTk6X/XWEz/cdmp6VuN3l3DFCXyEkZGFIhEQ35miUvprUVI/+oToiEzniyC6OpAB7ZQx6/x
jhEiZT29hy5/Vy9z6x2CEx98mAM3nNVeGAYI4u/SJ3zNNF6LwwfPBNvLFlqh1qvf7Wglq2u+xT96
gCBnOutdBZ7PNRnxtfeRNeqRwe0umoBkNUYz9p/J2uXawr8KWxmhiPM0N/h7+e2kgv4QoXRHjwpe
ITAYN3Hk/9+FVhbcCRu3FSRCrb5SDl9tctLRUPljpkHfYCE1rhaaTs+EI/7AttJpp4JZ7OCUiNtx
T9dYMRPBFE2mP7vG2/8QnefjrzqdSWBWkpx1m/LBLbgQwnlG5a/W922Qa+zqukMS0FqBcKVR1ksc
hQOXn7QLdxKcfyniKZ7s4Nqz1dYe11LIZPUt+PU7pmWFnxDXXKCuLxzLQB1O1Z7Mkbr5C6j6tqWZ
GnB8SViTbEQ9CxGyOUP7xPgo/mf9wquU43lcFNgsWJR5ykwaJXhwOpt1bcFft4nnPjYqM5cLFji1
KGyLxxLb4u5F1yAX1/pJtfoWq1mq6r9t+zbKJltR21fMzvBQoqBffusXE2/6FDh3VZg8DNfqeUw8
knh69Z6q1GqMc37GW2JI4kzmoFb2PG4xWksvAeWfYjxaUM1LRvzqMTh5j+d6n7jfEfNlKqmICAcQ
5YUQYDpSjB0WjYDFtOuq/Ldap3wL6J47LxpZjnx1oKIDVNcG0qDSZQzG3QDzvd7RrlZC8Bp90uNM
TacAxfIFZot3zEXzYuFft51EuHQDXSI5uHMRO3PtJy527vaLJwnQa/KkDM42/fvzXlSaCVnqB3AV
iU+hdxOZC99bI8P6Ezses4Utw6aXSQmv+WemV8+KBESIEKpZwfG5mA3cT8nkWjMDcCipktfA4cgX
JAuFSe4WRXaH4mCzI22UapbdeN0l4QhvQjFQ8xwupi9eliR1noshGdP4lzE+kzCKFovTrkfk4rAw
LEn0TOvkx2xOjP07uvqDESwZCGuaG2/mWHMuJTBQNv0bv6KTJOS+kzlrl0aFjOL130UyMELCWarn
61wHe4vnBqtrxMNPfskespZw4s+pF7GOI7YlW7r6JXRISU3qleyli/WSYaOtSy3xF7kSzbBQzZBN
BNfP5FuhWodfd7rrBJFezpPjggHiePhsJvWTG+HSrHHMQAZ6ApOb4JeijAzUi2MB1v5ksVkTH83k
XZOJxg99e0ks+y2yZkwQi6ynDcmRScwPxMr6vPSvhBWTd7qpupaF57RoEYuQ16SIJk5RoI7zc3HP
gMkm4IfC5qcldT1+vrUPlOY9DLPlyDhR7LTx5EdM5Ev+IsyJ+pD33p5kWju4/whYuLcF6N6QeSgo
kraO6vw069mic8hCD3vl0araobxtS77XnnPqs+3wE2rgfs8xxIWcFLc7opH8L75v5SQvTxrCwhLQ
IPJgryx3bWJRZTR+qvZXmdRPJ6xnoJxQuRKCnOF+4/LoTiV81Tbc1T0FgZXGQ73PlCxSEJ9Q+rbg
j75vfoKLm4+LnQFXNtcyPvAYXPUkqfg1JBifVlga6DkWfqjjwsdyLj2Iv2W9msLZfD6FbMds/tbH
ylLwZ2oHnqtodlQoYpK+gBkjtHGuPoD0nnrYZZOdGbevWueImScD0vJFKp0Z14sWUsKqN1SUsUTU
soRycDVSAMln+WTaEKuJnXmnBCf1u2qCe+fEFAj0mvm2+F8NHeC0ZIV4E34bv9QoTwHr6NmNQSRZ
L5NwxelVWkia2ggiK7s1KwtmkBQilZ7BEpx6NzrUoSFIIbE6jgOyk5ZD3UuzFZaBmOPJgbFh03Jy
3sDFDI1ubxH5YD0f6u9Q1X9DGpFuZnv2CqRbH7LzRKDGaC587XUtX3iXc6m7yDZwp/lf9k949+2o
lkx9ulykvSGz/Rc5VhT2glAn7o1fHKIQUl2dJBWgyeQOa3pMjGs582aiNvVy+XCUOlM3KJz/NAnA
LBNe6aD4PGMb89Kzuq98289eEMbQrwqeA1M6TBJWQa84Yh1/NPQxbuB4nxVCVbxDIjzXkwDPzXwM
YWLSNEZCSBES1vQyX1AEkjS5qEWQDqaZOu8R2yUzbsToSAi1mCiA2zuc+48+tcuGzvXnMgDl+IAF
iuI0K8BgWvojgbgH+d4AGe53zxu/JlyO55MPJWMwL2Tc27OhIzKEsb8CimBF2DNRSsmvgr1a/Fol
rWNdoIfHdyF1AqCh4HCfqUvjkoFBlmWNZfDu2ktNYqxQQUlWPHRqlYwLrttK2i2Xko/6rnfCXncU
tTT+KJvD/X1c9btNFtspaJMMUiqEtRQJlARTPM3oCb8bmNbdQJE/aNrcAV76OozBNrL3SkNntKP5
1yK79OSNdZeeLSoKnMyywchv9ZL24xEahmarpBdnCrvSyympuqpSHbzl886NW6l9aa9Dl6niASqW
MJG9c7gwdTBK/BG8UkAmiqvrIBIjuH0sAs8EUfSt5elwmIQh8lH3qfFLamdq+U5pq2wYqTxkvXC9
s4zqKsWZ/JlYDv+/rYNCVissfFAZwqXvumGE34a0PwmTIjD1c+ihUwTzCevw/d8Mq+8WBHDO0rx6
Qs8BXRMWLtM2cUVbpn27ZL3obOboWeKsZc7/0CxgrP3uHZ4kkA5czpBD8VGee4vkX/iKBhvYYnGb
izlHPEbfpYsMP5HrPqAIGk81+wftkIvd4Srxr3TgYnKDl+fQxMOkQdpEN/i5OgzADS83DBK4AN8s
xOIX5qEXcmXxdpz/TKErjoLMjEqkG0BSQup7SHVVWywsdwJf1PUGaFq5nFzt5AnFQ3l6fGJo8QEs
i2ln4saE4jyHbCk+r92+oA6Fs5NGKx46GS5J1cjHvJPtOJ6ed97EMpmbgG29S4G3R08QLhwdBE9U
ZMpyFvGhWh4IBChQECCJjRTINP4aArcQifoyhBadT35QDOnVJFd+6NxeoNNvaCGC3jDbtbcLVoPh
Wx6+eqtJPxTBiamUxnI+vIHwG9jSRvMfT7Jh/GV1Pn8qLqktEw0yWoOEqB767n/ftceGw74TF/yW
eqVnknQ1pU88stI0wmC/S/KYKE5fllFOedtXiO7Qy/IUv7l1zFgr1EgKnPfOk9o/Yuna2SSAqmxk
0jNNdeaKGVgW5MOl3CFAV4YHKiAPLr4rm9BOy9bFMDyHYG467FBq6GzZdpwxKKyEoATNwopRZJ5n
tljthlxJ3jGCgUcRrqQSRO0sM5EWtvEDjhaYG/UAl6Wh2226RYN8Jy5fZxi1kaREEtcW41tIiAz8
Xve9sJBK21lL7Mpp9d9F0JEgqYatmiHgYWz4c2BgBYAPk4TRh7XNkF1jAvOjuS4bVAe21wzHCM9L
3bPppwrmSIpwoNnBAcxU6Udw/ITHDavYVfkaCQQEAPk0lr8r9vAgg+ZlE3wOualbuPwrcWLNiX4n
FSi/5EExMfe1wrxSL0HcdzRQKSRZdDvP4z6/iDWcYPm5NU6Js4E4vfmuy6I8y9sAmoYnF1huLY6V
vK4FsyEM3P/vYbZfK6U0rJwG4X4rwR+6MSr4kFOjZmPV/RLB4QmkJyK8Iq9nd3CTY14JMa5yTCDS
u06ff99GUZ3utgiPadU+a5XaXFaF6X1Qf+PERT2PBHMW6fZCzy3Bk2ksoN3JYTP9Z0PdFxs5UsZf
5owTFwhENpWlFhxEuyyKqIBZRbgMaZNid34n00sgZOHVIgQSjin6TZCPxISd472qRXkdERqki20h
9eeXWbzPsudN+lqcLDrTstQTETTQkaSWGqgIoAXbwVi2PQR6rQ96m1Ag/JGPix9iQBHviqVeQ8FR
xmCqRUWNJrQrE2txrgrFNs+CLRYgDYgLxC7ToHEHvbLVc7RMOBveSUEsyPsz7OJg6WsNPBD7YQq1
7CI+n8GHNbYfU+xIDtdwxpaVdRUdcctJm1RwSkE81A3PX+inDfNJA5lEiWo95MgtLd7hK0Vzu0+Z
kM5s6GtG593ig+lcS9czWnGnXewKB69H8/Afm12uRu9YGJAhbkAyCmVxA4aE01FX42OOALkImYFP
41XtcQrC8Ko6vjNmxyeYW3a7o63RU605UHYOpPRP234N0NRJwUZwAep8kayK3HYTe4BeI6W0vZf3
EQCaDzFHod+KdAcF8jJRo2WkANG24kObcRfqkSJlZ8WFUtBDna0xK4EJRrVLXmPFT0UlEhpeC+z1
0uHutJKRtvjSHYrIJ1RH1j/FMJSe/B+fqu2Itn9Qwfb03Wh7sJxJT11FgRJcAAACoznsHX1+iibt
pr7oVFTj9C7uQCG+3DhDj9UX4U0jfyD4Ps5ZznT10BqFPS9PynncawsiW3TRgXk4p1DyqzK/9FVj
7hJ/wOZbX2ik6GriGZxlJArWVsld4FlwWiOo91H3H97BqVPY3GXXt3sUOm21wgbXb4uFs2PEmLp2
vkBsBmHYOkfJPxkETMb8lIPFinWHhilyyuKXKNsntwwdwmE1l46r8ezCS71fthL+OhRQbi1hCtu3
foeeFqXIrEbEHbjEvLgYwpWGy+kCoGNMQuZ3IDJ6IosrpvQjFyXpaZ9q6PyOkStjU/kBAXCzAuuT
iXPkngeCF4FudC78L7wqWU1xUgwLoqMmCrhUlNvMf1YsFwSEkqs0M6Hf/qfegA/qIlgfPLzwkD4P
Xn4eriiPyGxsRJisNIDYOJlWnXF/qtS+n0pdxwa36/0CjZGKeW/pHdqyvXIhFjGd/08LptpfFhas
CmBGhTXT9WPgNHk+GkJ76jyqLA3LUdCnR5o0VjosOkVhdrg8GzpLCbtEf5rD2Hwih9vnuccAjYEy
svjHn2uuuA5EK7CtZMEId6kBORVmGhaJOqoA40N+NBidPyK4NWqCNrUs3Tz1LzgwkH5+P3Z8q+p6
oSltOjIK4v1tQLEo5S5tN/1jhp3+wYydJfsmMEyZQT4KqG8mgbRLHcwWltalDsraqIRHlJzGeUM3
kFzYht/4etUp98vEg7LkJx5gNT3HiHokySZFqdZeX/GH7EbajSA7lFel9ld/kB6V9A/Vr4fxOASA
cuQfk8gqLEVVWqiYvvIfZoZepXnFSesD7f9bwbFF9mpsjX7iHi9v/8TtaW/DQWt24XTnQXrt8NOk
V5o9k8itCgdOwEuA32j9GKSQB9A5DuMelMO9dURdVqJSBE42Ei1HfVd3l0Pe2US++wJCeSnCEmSE
qOApTn7YVQtdkjJCFJNqBnZMspTJ9dZAazbyR2G5xKZ8AMSJqcO38r8aNjnHSfKxX7b5RUd5Zur2
+1BGrn5Ko/zZJK7a+PTMsjI5Lb6CIUIgq5ghBfng6zkB+szvu5eVCNOT/0iJwgJTgvDPhaK+Itg9
SrQ1gww7q1kdX5NwNU3ySLlU/LW7UbUumf5/9jEcfAHARvgl7FHbAhv+MZbtrD/KAAH1KNd00JOb
TBHh7dW8lk28sgkhda8b46gyGmaZV8xbTBvPhO1fk63Wt4IYIl0ktDrhMoIOVGSWDwz7AN4ZJg3b
1rjyq6XXIP2k13sJP38241izVocFb6a6rOUfyyGYTCYqHDa+JpcMntSw1R4ljT4tdD37vxo3sHZr
Jar+WA08+pP77AP1O0eFjio+C4F956gfyxW5cfgIg/YIQVwaMfozCvAAFlZHcUFQm7UrpQNhtJO6
l9DI80rkLBFsNWXNB+qD8eEVhjfEgU04y3aMUe6Pn65hdtAdfwc/XIMorgG1XmfBr5rZ4xgLidPK
js06kLQn4qbCFzclx3TwJXOqIiCSJsXQzclpgN0a9428vmdjL94aeWNYdlrGQvB1Qhc+niGx+09O
hHcdfpZQG4KP9XXkDEO48UL6xXdWJCDlsilKthMsSel6/BqjESGVWLl7qFtz5M9WDK61XfDxmb19
gm7CPHPM85sA2CdroiS0wRqB/xsPlaF8ArPx1omEa7kri1KgEL/M91pZ+oUJgu4mhboG9CHNsUHN
QVa7018YhHDFrgbnemmaaMbjxD32ig4BtKg6DP+P2QwTFYF0bCDmJ2ralN39NICJoPuxtrfJnjPI
/3aJWSrXncpQbDzM9do4dDtzvRevHu271z+o2ZUnkEQqB+c9H7za0A3SR/WshDJXqfWxxAFKFx6R
CLIlB5BCGL0vovV0S7HM+14H/vXBLuhFW171wJfdr6GibeWNPFiM0ndxEJGDPu0QL7Sace76ZDy9
NrzfUmC21hMaWlTpXeGf/0PmllnpPkSzShGF6fjalHFAMsqNj00063TEXGpePjyLMporZCfnzZxd
hQjisYCfo7H5T635aw+8KOB8yOjrSoiE/TeyfBHtZgPYW5XJb6M7m2517gKSalUcaUIaMyJ1L5Tz
dvV11d5sp4LwRUHMBBs0e2Tvf5w8PA0AfklmGg0F0gLRPpBrYZekDL80OBCNITBnTURDYy8h6m9V
oHE7uwZl+4bFeQqBGALTSykHyL5Va6ydnNUeugOjg0AhRt7AZZB0sKMqKRKtaK4psWidiwjdRhe3
VgJQcpSeLVTb0XCzWsxaHm0uIhbz1ghS1lt6ihJOIseVWSQcbqnr0DDCyvsLkmu6YuDChlplzGyS
XKK4paRxm7Z6W1/cEQJ/U4gyok3ILGQ9QMmCz1X7cBKxUi5jdZawVwRDWTNv7mZNeRIF+POf5dul
fJ3wEe99Aux/072RUNVUCx81AGXg/UFXrN9mZmczM59yv1XaJl9nYk4UTqpdXBVbq5mHmq6uSj8W
pAeHYmjgdV3eR/Bpzkgv5tR25iUAQI8gkI4dVlVewkKLjtu5I2bDVBwF277h+L0Y2y+5ePlYrp98
J77wdRtqarpNi3vRhhJML4UTBIkqfGN7f7HbK2BlStbwNqNaC8paj5BrSh6PnyFtWqScorxW9CiU
YaZEmgHmzfVa6mjz/3jKWbHQBEr3YMPuULd95RZM0ZawauDvLnT0I5rpW1DFYXePC6DxlXliDhCN
GKYFnklQBipeYKh9xWrga/RyPopuN2WyybiGtu8NNvJBoYgIcXMEhULg8vBRYscH1/rMrjSVhiDQ
EGyLnG2P8b87oJEsdoMh44l9C+j6lgcSq2Ef7Z8PoWcnmWrpFBqtqWWVhitbV+Zin2jCVviSALQY
e5Jz9qicfMjGwJCHhWdHXzBy1vEjbjD50u+4n3zR7wdQnGZXlzVMRfYqUwuMrbQ07eXOCE8skPw7
dgJluu7c7w9J5U4dupoqTrqYZFwMEZ/NaxL8c0y1bZvzJuwTiaFHEENePJ16GuJ5VeEPGuF1f67k
EoEpIf97yC5d63jCLCR/5piXBRbc8FnqrUgH2A0yGriVyuHtIMzzawRWyFhkE+B5+6HojahtbTie
gfzdpXZNDqOv/k2cDhjjPFVY2aNubOzo8a9D7tjXfZTmcAsV4X+s0oA9Zuo+AReekaRDCncLP+uF
b+T0i11k8zoqNEseis4aG7Z7CSmUHl1PK320yvmdLiuulmbvCowACGzwUwlcp2J/rTbwQm6QPkSO
b6F09oEm9+7bnEYesLUBU3z3wjBdNviy4aAKdPm9Th0JtZ11U3RodykMDAFxLifMwiNK85j7oBG1
CMxJZ7J15p7YLpHuw94a+uobbxCIiuT/a3FKRK/t9YL8sxXhGxIoM7pIK0pkvLv2E17kNSLqDMAf
G9s59/zvA8Ynre1tWwsBWGtM8HP+8ln10bfa8xT6qJ3GWcREtLzU1EP9/lEA+14nhinUw3by9GQ7
crU82xZmODyKUEUEE8oyJ3NrvJ5F598JRaGgQkxEQLqP07IGll886j6YTPTtG2lnf3VjtoROsz/g
gWjUTBoihd0Mm9vD79CoItdKUNl6fjAGfDYMmXXqIBKAVPjSzk4b1hkVGEf3qbyCrTRre2PXhHVn
12lQpXuLpg7UngDgFem6n8qss4gPtdf46+Pmxi7EkOjN4a/p08glfO8U9fczUi69qma/MVOBBQPv
pHBOgXw8oY8C81B7GWvsuToBEVoR/yIYy9N7wj+2knYmhFpRYBgIQC+5cMPnveEX44e2KbxSI7OW
p7w0GpZixqKxqUvAIvbKuD631lMr/ofTYOEKyszoGjnyuid/7pAUacmCsOPpili88lKQurZ5UmEh
ilG1BwLI3luRFk7BtMRS+vswiGsjMDSppWRv6jrlOQ1UWeLrSnNK25pGD2BnXvX3VLZ45JzKap3X
qYbNE4GH2Nusvhc7GsZ6TioHR89VfQ3ZwnxXcKgYc4V3JntaiY+HgeJ1uQjgazdZ8hcFjpkBYrR9
VyzhNwETS8x/r3VYrsaBqOFtelKHWsijE54tdrv/dsZ5r2vZ4tOP6cMwEIzyV6cEi5fR3DeiGA0r
6bA40K8ChwNE6HmDjpEykxpOm+Fg2gk+/9O4KyKCS+zwnsuFB1GBQACQ1l2T3RqtuBZ7hpBaJKHy
YVoGMubZDa7S1KHOQ0F/R2hSThFGOxXBtevZwZvn7R3UQYNdBM8ANcj+tfZxexmtJD0lSaJcRaJx
2kWubjr0iCtzkq/DlXar2ED2B8Ui9nkD6fT1tAPa+nOlcPoM61/ZtfRYs0iPXbhvBPoGMzWyxAHD
j1FfIbwwbOMX9Yn3NRGxYh93dBgjXtIgyiupbbopvkPrQe1p6xJjdJ5//VlSHYtbm+QHMXUAPW1V
o2xBy8pD7/nd9GZEpk3pAmWTtK2wi369zfwWOkfG9Lgdk5tmzU4jP0dEMXbyGf2ZBve7vPzf4Jit
dAlzzTv657s9TpfBCnl3Zt9IPG0RCQH9vK1HMG72cMH3ciV4ZCVLE/D8eiEGrb7lA9ZuLkftrI9t
/bQXEuXVRRSjzZOIIUL2qtDGkv0jhUj3Axrh7/zLN50oJdLC0qlpI5XqbiqraLW/vgLEtylD6Wn4
5PeJOo5w4TjRh7ovJvnyOY607J2l8/FrbbLfDj66OcMpA9KHOwS97renGPkw7x1sGZ2F5pdSGUf0
IClo3fdp0ebAmpoxymbaO/bTXOm7HzeGPLVAOkrAN1KGybVHgXPMvo4esMkQyiCATbaBnHmmQU04
3VEITXrNVHa7aruezTeKYfjfzJB+WCFaglZMDoYv3AJCQPZvqk1lYL3UtlxGvwds88WKJxembyn4
8iPASOM+zMVcysgtILLrUVSbBrmR1i7R4pM379mO3ohObdIco51L0DlDoeFNnWviSXVYIwrR8i0q
C+rrl3+UDL1xqG0Tf1i+QvIyHic7N76MKpPrV1VxdnHFkdyUliZDrJJl/unM7hrne0ALIpxaYo8k
7APB8am1cGenNKBN1bCOoeCfyvRuUWzJsbmNKg/j1BesoGp4cvOPfn4KezIw1LRuqvVLEqufW3hT
6Vx11E4ZTMzYGgWv/gjLl0p52NW1l5jI0jYmpEHbUOdOTwygW8JRKm4BoEC+fGotRdGKELyOrvn8
LqEmtz3gp4iaeVyjx3XSwXlCqUEcLtBeMlCfVhqRVR6qo4/iMbOJhih2D3Rj8OuWEIFm4eUeWQGj
jn/tp1SMNiIQ5Y7zYPa6TcB9cFJFEDJdKdFxOWmoS0p1CoGI1277opRpJf67bxgQhWCKBjjhuwvs
q2MCcDFt1agriICWMnYGoPXvxMt2GFBqZaBiBSWy4Yaee+o9g0NDP4sHvXFKOZMXKFK79oMfWPlu
nw7l4+Rpi1ODZMU2b/IDXlRSl0wSR9/Si6SgLDKJt1Rv2sPh9f0R7c/NU07rI5IJKRfAHP2mGarv
3HcOOSzbrzU9hSqCnpPooQUVR6HoLqCuBcj61r8OFBBLKB2UZLtkxKxWzxGTEfZ05DkXTM2WFgGv
GFFTSdhbvF00F4FA3xcIROH1wK6fki7pftUvgZsV/RLwzflEy+nRZwF04MTKQllCFm1oNmpEZ715
HI8YH3EKbw9NbWdPW3H6IVXec/QotoqNJ6yuoD6ZqOAfXEY3jZJDO1WK1XA8S3RahThejX1jXRl/
i7QTnuQbC3qaZvuKEaoNcdtlOJ5vqSR7xbY+1wXayKqK+WuM4znZiNRuvNXUEiEJCs8wc/6BRPgT
1keZVj3sXCF6UqUAeI76ITHWY+9j03zHibQHWPJlrz4GcOvAdzDG7+qWvfWIICn+si5uIwuEt6jT
YcLZSEI/wGIdqh/vx+z+lb1lupHLY2PhvNyjmcP0q0NWlabI3l4nwWmiqGJKcl0rrGQcSKSaI6E2
NO9kbV1keVQfmZDPCrDix2CdJ+QEDPfXfjzIe3VqCpgnJYMa43RtXHYyMKDRp2Euv+WDxUEt11Zt
T3UnytlGtpFiKHN/pTFIHaCCCu85v+qKxGa7dJvOU9Erzfc5qDLuLJVkWfnI+T18bAiiuTUWcX95
VbXmGSVqTENpH7qndvPIY6LrrAkylh6xytrsUyCYYKO2KPGVVw8TARc+dDHlikn3563mAoVO8/IQ
kn45fPemaY7rfctCwD5RPLM2gQ8s45BGc9ogJ9N46q0bnEcku6B6YGr6rCjmF0eK8fwWNX8nsq0J
+S3ECFgj7FgB6kUvhDNMYFRIELUq13OjppRuBa5RmRg5AzqXEgXGc0UWKY/6qmOhv0JPH8bG8gpv
K9VkblD9FplAi3vUiAURBfNrS8Epmgoe/xJaAk6GEhUEJx4/wQvdahLxxdV2zJu58hTUqmH5/dUu
26mg/BCjxjy3XECWo1Os0Q61JS/+gA9tNhdY93wZL/4ytyVvC/tqm4J8ExD32IEIO27D/gkfWSRA
65/NVh3rexFOmIHWItvZU2liJ3BL67Bp9bqZYx7571aoWoyooHjfjuaMcLRlk6X+ofok7I+9NejG
6RgcZlVjsQjl0oig5+B0bfDrPg2JqgX+HUagFWH8TNclRd/rtepac1JlJfwJbQhHpkrFPgGzqmSz
xfbCgmU+c7BW9A7AKbOKuD1/ZL/OHQHwcbR0HpMCnfSPZg7GzXFw2xDhqEEpnrRKNB/xL3KYsogb
WvKsVMufFPjH0hehab9A8QESLHGewZpZELkttDv1pjyzzFYSNOWKaDL7fM/6s466Mf+RbHKjPYiI
qZo64wQakFwIERFSUkQ2o3LbpUCotDLoKcev369I5AGt/CN+YYRR87POs5Mto32o2PKtOtyGjh67
yrAaqd3wugckwZBOc2vro0q874sIRuZKaH2PKrK1aT1UOQlWiHfz8NsK3TbLRQx81BVYCkhG3jO9
sFmTKPrxmzOu8UmsRhvzVQ4CUR0LLSoESpsW1wObWUvekpr4M7hkJmZHq9M+QRvRiRdFBv9UdsKE
tFcecEjKaLktc54yJizA2df3CgiLUZMSW0sdj7v9XijhbzuGQIoWPIcft4ny9/bZCiboYlJLzM6c
1uK/BxjtVVb0vpzd4vhi9FgT1RHrl2mv51R2Q8aJ5Dgb0VKUWD5iybigL6VUGPYRYH8ZuBaUjKQw
WkqA1XBmwSJswnRtSlx7cEb0dY7a98bTWSHGOfbSCmOBEODJEP0QpLYrYMvJC5daAWYQuJoYRNQV
abx+BKGvLQOfeCZGCvney+9fGI0NxoqFII6D1P+L+iiYr1ug7qlwsD7QM4d7UuEPIM/IIDq9PV5D
OpqphfSIwyW56zU4Zf6zwSctIKoxWOc8z6bmJsB2lY84QspoPG1yveNlgy2aUquKniIRoxfsSZam
JLHV8Z9lsfavbCmkm7Cjn6KW0LZX7B7uRQfvs/nphBX9bd5nOKamnenKTDawmVghd82B8Lc/JQJp
dQDOQNwiSZIIeqf0csTQfottD6fY8bgnmYUOP+gS1ZQqRVs0rbHXG4LZg+hRHRQ7FE5xFPcgWNGi
u1BvGx+61Dp9JHTmksrnrCbApJxh7IVmPXds5Q7Jx2TbSSnr51CN6A02bHOVSIojS/nH1xPLrQXj
j3l6XD52aNAzVN3em2rZpgSmpKqV54wojwulpM4sJ7sbrHzmTianyrUpRM4PJR9QBq1aEaqxVTtr
39SMnbeoSnsaYkKdVz1x47W/df9qaJ2LDvtJmY7h+rGd8a4RkZywEUN3aY4E31ROWgL5sJ9tpsoM
R+2JL5Nt/xIX4FK+r/AkH/14aA401zpInL+ErEkCRWK9YwHrWjLoLGEW4wxlUTfIl5DE9c0zoNAz
D8nXOWOiiYtO6SwwTjdsPWymAYDyVVJ6H+i2cpAIK0V789pzOTx+5+9EZS83NxpLa0nU7n+tFv0q
LOprDKRUd4ssUHxSnkLC9iETy52jXaV6BvmZkRDNtETBSy77WBJXpm1ev5X3xiCvGhvwaDvCuszs
ZdJUz10G7lv6dH+TCyYwTW2+Cw0Dm+TKL665hd2lruPgHTfPNfDi2+3/UpiSkHP3KJlsZtKnJo55
xMk3Js6tdsDCiNvrDHObZBKOGTf2Nrex5VLxT82lISQfr2hq8AHnUwTLyGZgQ3lJ6XLSAClTpnWY
tlJUODBPdLagvHSV9mraiDobX83UgQ0D6M7rbo6CQrdnYRNr9IpqxTUzvc13sgq3XQHbuY7K5m8n
T48YvR5lYlI3pdrHu0teW9COIS35eTOK17EFP6tpw0/jCsVhDCxLfhfkETVzxLtdBT6O2O3gh8dU
TEG3igkNReCjDwNTMW2fHEvXJswMjSVw63yYQQZZGQkgid0Taj2S0fAqoQCxgE9c7qArF5DM8kQt
AbMwEe/HQCsVJL8aIKM87AXAt81kutw9Cs9XgljnKxYJ1NokS+5hG5aomyN//B3mbocFvDjs6Edy
Snn2zRNh1qLVDWqEGD4XAx/tWr2JpoSzMHKsLszFe4qUtVU6IYo0iFSEiz9gSradlMJGLE+3lqpO
sd2Wk+5kgH0e7suVW+k3k1IPft0shu77pG77ysenfCf6YnnEoz7MrYgQhDNXDC0GyiAJbaR9iymr
fDXiS5GsxL4ZdzvCJPBAYUwTZCeyPNbFxdPO+VcE+e2v4Nt8TtBcFX2ve7j/jOLz2bY9Oj2CH6MB
UJ5zsIG++qlpoR9f4ANJaN9H5pSJjnkn8c3umixEUXNF8M+LDGs2P6bvXta8M2NoldaFwQVC9a49
KK6djtgx8ZAjvaeF1FvAJJmxyzbNm1guNewEqMSiJqYrjw842FTZaWVHG8RbTvtye+/qusEyDrA7
2wyfBm5Nj9fMvjeclPa5XYL9RK7ReKLrh50eP2wmCxnhETkwJr8yl+00m0sPHaT8wiMg3vihZL7v
AHHxkzrfK0xwqB7ebB0BPV4gY6NV3OQZVyBgYd1qsqpQK2GJZPtGvsD8AbD+W4urWocZN7SZ6hv8
aYH/6keMrT4H9VJJ2/TxZ/6/Tu/dQ+cIgbHC9kQW/Wg2icTbKIBWjDicAu0ye5qUMOBkJjv6rbCn
oqMz1oUUHe6whsy63FJDIwzL4/dYrRS6SJ9ba+O09cTaf+YzQmeYrJnKJ1NE0dw9FoG2TdA/oZNS
zVwEraY4Ik07GinrnVs/kMd8J0NDFm09+l+ReqXkE5BHZ3VLC8PXk4mT8+VhyyUeZWjbJuYb9xB+
JvbERuaG8zlTCuOkAAk4qGVXnieqic60f3cm/vH5uIemCe8f2b1PD+FZAUSV7XPyVZZW3jOH/IRw
2YEmfMUqg5Sgf5msH7nJw1nYjGJZyd+Vv+wkkc6+jy0PNbblMVo2UI3rd7b+Uaj37tygMCeAPcR8
YKlh5AkHHLDxz9HBHyyiYAEYF9ya6v2oiD9YeRVt3fQurtJ+CK6BFvpm5wQ/jKFOHuSwHr6KeAy2
KF3aW05/eQJdlsPPyjoqGI6QTgFfPVVCOgiXj5mAUBqIB3YspLh15Z/uHB0E/bZLJ4Nvbs8jLJbK
nvw6s77uLHhGoO92llVlAJPo/Ui2BL1MIF1QBrSlRRNYvQsg8B1tDZCAlOugdkeqjdlvOyd9PS4n
cMjfBEwZ87NQmN76uTeS6mU3bWwLMpcW7L2ZYc8VuXiwXER4hqRdzw07gP4Yy5iGhN/297PnTlz7
qcrDBpwShB9wIUBUm1sasOIz8mx2unKV/PZVbrDhoseBTcR9ovKsaRYtL+432UckP2vFONbF+X3u
qrSICwUyDphFWgUbv9kqC94PvGv5XBqr94JNamFyFMXJMHblyOMJqt6PJCKJ5QdD6k9gddyYGqBF
/K7XA0t9msx9O+ukiSXadGouvYMVVpd6TMlVcDhCGDatOKyxpmoHCMZrpmcux6wOvDDcq9jNOq7Y
gSUtT5w8AOzNIZem/qIgHhy2evYmQfvxw3YsF8UsD1C7pfISM5YsevYmfVU5JilCEfuICNr0G1OV
4B45Vs78etGmYi15hrNHj1Bpgn0ePFU2TGbQ5hSf1pLOKJkwmny7LixJcspfYwqofczpurkk6/96
lYnTm9qgVWICsSGlC5uedh3ttJgip4eyv9g+eKIWreX3JL2dYnVmmUDy727kNNejm/apktPdanmp
LlcIjF+GILyaZX5npfMEhUHAn+kFGWZGZMa/wE1ilryeUxC7Vvr4mQRbJHE/ICBnqxWLlRTboTZT
MQl4zUKheEhYphJWBwIOClv0dffOrJT2b420QLYJI9v1hXXBOigwAelBQ/c+yFFi2CBIp05ll6Af
rg+vAyAdQ0pFEu7ExThq0w3tc+V9JZr25zlbdOPgj3o+5ngt/2K6MmSsqd2L7asdaFlkksxfnWdX
lLXLDIi88o5HH6BG5XtoTP6+jdVZbNPTsjUujL5Bg57xqkdj9Xn1Ir7hmQGirJmyBA3MHXtEScpu
AKqtoBTUVPMVCeKKjnwNtyZi0s2v6BT8Xyu8+3+Y0SDza3gwMB9cTfO2graWpkmW0nVEBcJbUYXF
99cHcGwLIIJ0SdSGbVPMgv0pW6MCe5pO7B3cJlpocMe1/glgAuwf45Sa7z7YEaN2MeYXK+s4q+oB
hLItecUA9CMh6e4kqbHUeO+R4oM4qTnfEEeR//D3KQMIuMkD2lxpL5gg87NI1XnnJTBu20xvxUYq
6AiHztN3lhNwS7wDktPeKLJbB44vdxinC6FMlLFasgNWIas2eqg+8qgrwy6CmMZbysB091gUDx52
jZhKcqp+ce/M66zhRJc5azteMow9tMfiWM5K9iJB+PjUdC0f3fI04yE9mtBimsRYTjUpluBC7zrI
0GibZ/got0GczTkouYqTmV9GmtE+qOIYsdgOh32lFOJKY6cDCiXNWOZA94XFonCoQ4GihMWFd6xK
Kna6iR5RwN/JI26zif4o7C2qHnF0Sbw/tQz/jTkotmzbRI8i+gZnwVmoCLFbxZUfB1JRYKpFAWiB
FuruN01Vm6IC+tS7Og/qEErstiILG7FIIOpFRldgMhgktjzSh8NtcgEjrqa7J0AViVZ9HVSvfePf
q0yT+qHUNwuNcYdxyDPEN+8xHN8dTYioQrIFayXq+G9LkE/HJd6iLv/DaMfPA27eemCVu0KRhHUK
VmwJLEr7WdHmo7ClAG1PQ1xjumrnWRDN19InPzCfclzr2YhXgr1T1O/E1da4nowM+jdfcoyEWOwd
N4nkx4Xoz18i4U1JYU0GWfA9xTVWf2OhnUFAraVjAvmqW3R1NxXj32Vq7Jl8Gj+sqOGbSwM41rtg
X1QnIjY17lGtPRfgtILn0MyTdD6A9e7W8EdBWeRupqM5pcHw3He2VT5Ttc2Ysch0teTIp4YmJVE0
9Tq+dRTiX4112Fqw+s13K0fSGqM7/8FyujeVz8urhAffHcwThmyPV22EDxdS0LAIBLlzRPxBIaW4
hjWKNUMbSa3hYhO83Bzxa0Vb12qmNAjUK7aNEiArQLjR2pbbAEnQED55T5FlQvD9sISXJW3fA+ok
2pDC8/Rdy8rDISrgoHlhUTrKZYY50t/eMNHHdONhzfkHVfFidIQfUWKnhMuyq7WH8BTP7a2fdvdx
Xwn3V3UJzqv471veOFUsepnkUBvyvlJpqYAL1P8/JR6bh7dzZTaCozzV+i5FCdH5rtl0d2IjMKp9
g+HsZJCLYoPm4HwYOmdP+sFdrhjEKWoTvsrWz3flsMiLCsmrzJviBgLWcUr90/cJMWhEx/LvUqHI
tvv2nbf9ApSWzvBv1xxHIN3i2N8C1naBzhFLcZc4hVj4uLJB4UFn9uMeBJtPmsIlS9qJz/N9u4Bi
cXc/wNQrl3bhASLHCduvTYSUn2cHiLBhyVa0xtSiyAcJrdf/oeKCNPl3M0euOMT5CDjHsE/AjYSR
FtEYHa/sbbfZmieQTca17aTsS4gnwCc10vNUeWqwAZ1CqMlLnNAYc33+Vb2Bk/8k9VDGL769SGVY
dUx0FxXLHZxH5XVDLFsjMd2FKiyoj7U1FrWknaqo1r/LRg77MNay9eYHEm08bI5urAG21fLHqWBi
GD3dV2H68OdUWRTLjrMAbKM6Rv0g1sxcxg9DqTsYwCvG2F0kPeMSpl8LRuboQHn0U9Q3rz65JqHu
2wODV1e7H7rjtQp/zW95octZD/1QuehDeLVPZRKf6hZ5H4B4B73qAWfiWhjCLER4J6yfcnG6CIdu
jNUagqJfFF1Whbv4eJuGUnVmTDPuDA+98TLEpKeswQl459gMkb4sFHs6knPFZjYaI0HASJZJzF9G
3p9Nux+CMbj7dPLL7nIw7L9Vg5sXVmLJcpKplNj5u9R00/2fcgxQY2NeG+yu4reMfnb83IvHfgbH
CFeOPy5wqFJ5RLgaZeWK7nQUrJ29wquwWOMiv6N/A42jOYxUH5bVKGa0oDq0aKbgUJ+VLXv/NTWf
u+fOpXA5kg7Y06SQRUnEaNgp6oAlwJkwFwq8iy71pKSXiCOOSMobnWbOJFd3rM7Vinka7S49pXda
LhsmydSumDpG7ZNTRhVI/pdvzToHSadOZlSn23X/ACUW3h9UEfuRkFV7GGFOe0xnr1yEOYhmYo4+
T0S3CjSFpATPW5Hs+NHCHPEdjKDN4U81bdhvG2auqEM/woQbfJd131pS5Gu12nKPXKtxztgsNLg6
Z0OBG8a/e+mmTkqdiewXot78aGwUFOBjNxZYjoCYwMI26Or0XPhRe6xwXBhyKFhFPr6eVIfAMViz
pO0OTFt9+zXx3y7PPyGa82zfKyF7CnDYMWzZrzW4O/dfS4/h3PxTxrvKQ4NTemhFJqVNS2Ndydxp
RjFl3Hx3Bt9rv2u+Z8WasmY5+iVU2hiE6QYupnCXBMUE3yK8f3bHNiulhNJuInuIAEFlA4w8yDu/
f5D+lyn7nocqpMc08X6s9QF35rBcfDhfTFWAFiQT7qP9VqpUXNBJDeyBNYwRyoZlSSbUORDlVCqe
gO2SJQScimrVPG+7NPGKm2c1IthB0ZviyK4OPyL/bjre33sN6L5z+GUpUMvfxe4eXDN047PXUA9K
vVeFXkz8TMbn3ntacffAaSNNYm8KFflFfBslgJ1SkbPmMnLbYvczeqCsvD/KoWF3vyWoyO9MlE0F
vfp6V4I5v/TWH04NVZdrmNa17YGBSpvmYD4VcyPD6Ke4/sF4Gqjiva+BrC2acSL00sjTSrgO/r0Z
vzD+Ho/9GDZEPpp/sWoBlFsFPHDa9WspvMHLw9tDL701KtM11dLC0XdkgNX2vmcNTGKYO5Lu7f4P
EMeDMf1UPCoDsG/3g4GIH+eGxzdWXDzda2cM8epu7yzHsrgKwrQunznZnGLe2LbN3PPukS+qqJLF
bis0ni4kNYYKkHJcKKagRAX1m8j4o31DjbnsOC9yxxhunM6lX5rMD3TcZGAwUsi3HdlgziG8mt71
sE48rOhdpR18kQCjRcon4Dj4/LfjZ0tqKv6pc49uPsUe1bxT5XkGIps6M1hE6Z0WYx1+KfKhnOYN
CFKioxLeZ0j+qxf/3Burty3LTKYmvVUxKakF1EwdVaRkOp9BzYLeLIqPa8BWaZXaIE92JHA4Ki74
xmK6peK87nxz92s1/107rMyCqkRJrYIhTaovraZlI/yYuuuQkO3E50B81AoNMyIOgt406oRkwx0T
kN9UuFK/SRAnoPTnyh6mWquJWMiCnGfKnhW6qDYjbtPbgirWttu0symR1e+tbcDNtjQQ4Bb5Ks0O
vVA4Hgl4uujX9Rei6+wmLy1GT8Lz9Hf3m/or7cRnIDJ9CjMShk4jQul6dGq55X61myPaI124GFyc
nvyYYGAru3gt/wVl4NkCdURpiJ+gQC9JISzfP8BmX5j0dR9mh0qp6uOyUj6+5aQzSkp6qViDbsMw
G6YpOMuRhngLUpfQoG4nX1/ekis7vW7D2oV+Ebyz8ZDDFnU/g7x+4K88XtXyKaZySKbQ2fNbZByx
opPxe5bT9rJ40+5JrTVByAB8kBZL1Ev39tg1DXxW0+y7muKZwx9sTOazKwLdEc/IjUAjjqZWqmzx
AbERfgcVbmlKcrr7XBHF/aswcZxxI3nafARcyXyYMFYcPr1QqiLuKw0NP6GmHT9q2orOpT4hpK4a
ZqOa8UjGgfNP1unVY9veNl2uY8Fb8UyVW7bXPjH0buKiM+49DmvQ0adrodJzw869V6sZ35dvfghF
/Q/fcxKFFb0JDZuyNfCu6VcsOnqpJa3YrCz5Y8wPp0QkyR2BvpETg3UNY1aw9eFufDR2r2vRehvm
dbVME2Ujjj+XYhaEteAs/HUcuTnOecSpLY2ZoCVn77J/8tz+BU1TAFCYqgQUsdkkve+GSw5HYwRv
eR/gPY1W1MuT7DwC9j4LydTbbRGf5YDlxT4S7DkXs4iS/9vt9tg1/4B1dzBGVJQbpgFq1oCVBU8K
ftpr3vsRKFxrjl6R2ZjWWaX6DHgKtVAKg83fWQ2iM/B1KxOfJNF6/gO4k6qi9gyksWhuBOIoDv6k
QtnDwox4cV35ZJjZyzv8wvVv4KBjd0qfNW03XwUpfucVdd8xBfLb6xI0UrOasPB+eIAXhq5wKcDX
QwBY+HEHrlfCwYp7T0Xp7d53sCC0vPAbbJEvkIua2+k1Ac/qaVQS9O5Z23D/lkcbIJ7mClrut7fh
Pln2fL1onspLRRvM0j+HanuF52BUmQ1nViYbtWZLaZR4riKBBSWGltA8PHopdmPRVeSJatysGzum
1HGd5vGWP1GmpyR6Ja/3e4ZUfxTnw7wb3JR9xUZ7wL2T+SiAq4qG91bzadQBRTmEIFO9zq56uAX4
jyuMl5+z8+BNOhrgl0+jSxkMy0/R8zl0q0T+qL7Y/Yg3Ei++cYkiyTmApYM9CFa2aWB99pZ6Hilr
Sgkf9kM0wVHw3sxngvQuQKmHBRUIEllCSfuiyHvLawqSC2EVkuunjhLewCTXdjL4I6N8Ihki3Em5
GHusX8w046MUu7MNNah6JGAk2I8kbNmDXTEjTI8TOqothjCESotjiZ0F9cymdQLFCheua+Vr0W0v
xSMNelsaooit3W7RkAdzv7Im2F8wPkiXY29QJHimCx81Rz27VNFCG6rtb0e+KKRuvmrJv98gYjOG
P3D83SF2IPjesrfqIirB0IGZ/soByEDNzY8O0/TWsWJsyjXD3pMoDecQiUPRogPs6IRZLnwBicJh
oWtL3WjSqnshx0fSDz8fa2c8LYosEjSm6vmo8JoWKUmq9JzZXIkick9CypsBtKv7UJUNK56jRvIO
0RdxdN1eDN8NpCetKzQQt0PODeY38B70qgmPQXLqF14X8zZlI2ej9M9tAhIGhD0dYBno8diP2jyy
zp2p+TfHIlC+Rq6/Fxfvd1bE1j3NSsEiNt++qA0ziBTN0HF/RKXOyckFY7KQg5OLLMRTwMbHn73x
jP57mQZgsFNps0B+rrJbdVT0XaQpOPhvTb+J+vgvpsaFKxWn1eCBNMkapHEXEtU0gYpphy3roDvb
a/Eqa/trPbYonWK1ZBMV20ni+VEHNIYXOmF9cFbAhSpSzsKFlo4FH7OJi6IJAJvd9qPD866khW5v
y0JP99SYTqH4WPYAegFd62E7USNqsxK9ABOJH//8ENsG2HhqBtGiM/bqqdhlhAsJF0rrJekEcGDY
9Jj16/uK5mPWyfc+zMWNIR62EndhgDiXEQx4WfzvA6lqA0yCvAsDcOCeSl2EkIDzW30lRxambsOn
G6bS6lCr/lSoTtVsop922ZccmBdYnsY8nH9Ws78R4fBBXvCKwKnCiwX9Q/okJ0P00MyUvN/BrnDt
RF+RsXEwqHoJfsUHxS21IOnpN/NBiLlqCk5q64cB0ry8Q/Z2aIXMuNjPGhwv9fEtWdEq113Gjrxz
qX8RQztBi3UjT9h2hZ+vsvP2+Ah3w8pJ6xxDpmnZc1sPtwhlutLmlpntK+KAlt74LBaYq9JuGcSr
aLhYSDGFioYzZZbrfjzP89ELc3l9xSMuyLGarNYSScz/3T1VkspI/syqE3V3Ly4PIzX+JBYnObTi
7Slat7XXMKlKZmgErPw9ZE3+uq7/jHmdjfX0cCJLwbHteuhmva0W/0mpXzrLZEMyZimZWN9DpLd5
heSUNNAeAentobzAbt2qXhOWyZn3Hr+3xY3nIdB6cBXILf4IH+c3nvz9sf/HzZHmNcn4vVxBT1yY
/hWEW409WefsIIEyHMcWPgYN3WxxLJ/xyeAhDbrKEfBky8WnC+5wNb73f43L/gZFgZcskGS3Sc3J
BQdVSaOczWvMwwfbEZCFrzdZJFKwUU1oeWQyZxAiIO9bjakV6btuIm9cBPHVeaGdTJXWpNS7xc65
N1q5Q623soaiai+IEydhe1Y/WtyJgnNgpBjfHTDkUdqrbEAbG7DWRdaVhKhl1bfg7ENwk+vpfax7
dtMiCINVqlWnqdVRGIYyPqpuFQz5+n242dgT7ak0G/beIKuPRGokJrs9uY3WGyHHZZLG4djDz205
pZL6idFcqsQbEVMtQX06JNfBNFxCFngJ6Nl3tqJZXaK0WnNnDS9ugV36Tn4Y/+u/stcbIgZtLZd1
YyUQDRElXeQaKJm8VnlX9LtVmgHAWRz8J/wLaOGi4XckE1WBL1x8Lf6dzNk7bZWQtEWWwlVEQV6Y
Ol1Ee/WTyJAnYxx1UNoEXK/6Jfuk1FVsvuYvKZ4duXDpzGsEGxu2n3Dbzk4ItJaclxPh7zQsF6oI
VuM7EysSpkRNQscFjZl/J0iinKRfYIc035uudmi7Esw1jvsbECEeRX4YALc9RNGUuBpB04nde7gF
CBRbsr3IsldVUTZJ2VlwtvgcLXfFDN/+GIKHHcfVpqcqXdp/f58lEv4h3gC3TmBy9VTl1XOqaKtd
rrUTSMnQuJ1RWy2pVWgmgEo9C8qqB/DIrm6thqqE4WEc6qxZSi0BUkjty63A35nn8i/VfrJIgaV3
F8sOJcEYWqWgITvuaMPQktoafGKGVebtv+9YLDxAhvVCbTX6fCL6LcvuGXAnsMX8YyXdUpTLAokT
BdEI3Ntu6/OeTLZIhRuNNNMzlsdlxBll7fTbHpRu/sLxhV2HV1NhO4MjKQq4OXCWucPbR0r+ovv/
AomtrxmbFXSyRoJ7cqHMufRQd1hjsTf6TVcsquZB6z/fM3FXuE1emhHUNtZ4DQymTUhnzGd44hbC
6J2TygonGbXmrlvrwNEoyCZKj9bXXsYWoMGyU2OUlGTQ0tm/svgbwlcxNsN9vm/pw1eojGr6SWsn
t5vCZNzMTQkb3aK70T2albi7sqM5ykVNJTHju69gG22CkA4BBioIHy/Q/Y751U2FqL3AU9hyMjqZ
E8hwCcQ0kdTKgb/GWdI80KjgqUTgUmJa3DCKRdEnht+2YA8zzwkT8tI66fus6zPbyWljx2i5AM9B
WT7n4u6Jyatr60EnVNTtGHeogJz6fjpR72bcArbyBgiqVRqQsVKyxEKhzn8L0mcqJXqoERjkNboR
h/x2uQK36LlE8G+9XaADIa2Lbg8d01jfnAeamidT258SiGNtiPRYXjXLGyZvInV5rY4plZlsMYLz
a1X1lbJh8cSIpAk3UE6LATz7/LV97YQlfmxzPbkW9m1jq/VgZHICVcOvgaoB8blFHc1FrIOm6LrK
pvwPuT6zYOTuPCu4IegqWsWzUn2LTBpfqi3JPHIVY1HiUbETPCLgILSkmUirp8XUa9TCQmIdotEm
Xeco03zBy5aVzlvU1c4mQAxODyznvrLs7VAo3Y31BANPDFBj/Sj66oYizgiLp9tlixCv7tyy4isF
CTRK+olRUCMbKNTpH1GK08b+pNfR9+oP23jlMt59WOgQAlcYK9aOzw5PAD4U5d6RL/CRrVyJga88
5cNX7ThB4o/K9A3LLDzMF4AIQYh9v1mvf+3mvFBAyjtrCfXyAf1tB63eiTQbfnvdNfkzpLtC6vsG
MRYHvGKyUBP8nBeipfc/3TBJva8+9WlNZMPGB6ppoEBdqVnsI+uzT9zbwsKosRVPrBPp+MV+LKRS
LsTSFHz9fF7c6qWi36Q7rA09ShIEPoa28l2EH0YFfLr/WxEQmb0io0QeyrZsrnMO67MMWuKvwgTE
plinjYKtPwJ6s+BorNz2nlz5P9pH10Vjkj2tGIHYhRL2kztwGnkMeI5XclbkAZJYNvgbv1Nwn7tH
K78BQSqfHCoFMUE0vw/3rC+2FS38DBjuP1Cq0z3TTUnIcMXtX0k9dKdrijixGhcoMyu+Clq1gxRm
pJLNZ8MKsirUYWtgVrhlRM64j9jvpL04cNvmwfBNlFWJbZfG6DD0CDYiVsZ64WmGkJ9WbyuatGui
6NtXqiuvOwUuoNxTsdKZuEamyQ/m0pIgqZFQlN4zD/3io91PUyKNeBK1vRf2eqEYeChAEnHVV0J5
v3MCgG2rlDti4I1TMMqNco64ZmlcGIOYcMJsy5bXA/RB0qsRcZpt5eUmwEEhSURtVEbaUl0IEgWR
ug++Rail+V/rbI2oe+Jwquwbt47HxPforEWpJweFvPATZ3+O1EMBEiLQX1ECBcoy5/BplGE53DsW
4Ew83NWLCXu2BZif+/ZqHvR4JaySQHKSDdiV03uhlrf1uuIQqOotIRBajYvVOKLJr/tWbcdB/5SG
1buCouFm8qdfH2y0V7e9AsQicEFeqbpIMF/cC+E8032LNwthYMXvP6o2RXI7kjg2r3nfds/FKpi0
s3LKf91AtO55q9Ppsu/V+jFQXmGJ8anVBpXKNBSW6ehr1LAbj/xtKHif9Jrslsxux7ycBGLrJdnH
G283AAKIhahp+AG9SJxm3wQxU3y/pvZbWv7TGTQcTnPXZn6D7tIHAVPT3hKu/ejLLm95jTADaEKV
L2YkHwXRXMw03LiN2jJkyFHcJ0LNGoBax2r7cgFKOJwXi5uJVNcfXopY2IdvIh4GYIUTSWZY8/qT
tf+58ubf1sCK4xUhdJzGX/2gyzrhnrs09bJYPK1i9YFBAKhCe1QqhmpW4QP7gOpt2hD0oyKC80pt
9uMo06VAAuvSXPhxAqaC2SBGabC+lu7uoVInjrr/Ca4bHSiNMY8Z8D8MJa0BhyxeN6fMJeWkqY2x
9gjWWgi3TeotQsmNiqRKfWyGRajVDqvgt/hXhEDNSQKLBQxaVtO/bG0MrcDgG5n2ADN64Qo1oVkO
oy1v7f66R6uA0mgrx/kwEBUS1p9vTu/8XMzahhYnKjuNHQz2Qe5pL0wbPsZ2xkHvosCL+yg5eoPv
dmAMYzs5GILD0fm3m8Z9fuI0BGvt17khrk4mwr6Eltqx7PsyuL1zFY33bylc6v9hz0Sl2vJG3sZ+
Jdzkyqny+p4ZQrXD1wJs66OYbXS3wUfOYkoh0YfP3wGboyV5JgYZ2ik0C9gPXyGYZA6+fDaVFm45
kNwTJvRdEZYUWBAVw3bV0icWsJjXT/7IF5347HA9C9udn00fty2JtIr5HA0ViKsK9rXxQbx2TzC0
yneXWmYezHLCVWg5cAIkhHs9AHh0iXD16p4U9qUa5MmOSyQjN0meECnYOXEM+yyJ0i3bgusah2zb
Ibx2Pid6N2Pg5RDAZpMRiFQsZBpUW4MlJzeFINqCpan5bFJlSkLzAs4bQ0+dBFUlX/CviKDUq6pd
QEN7j8OWD+KK2jsEjnW0tR/gHfePeXNxOu47BzLq9o+91ftViA9PBe5J4CzmJD0HpesgK81pxNQn
q4TDhEP9kv14m8J2l+ciFY70UDrrH90HD8yC3zqGeAQpsNJuN8neEbjEN45AHITcdhMW9kIDC+D4
y3tV4xdqt3FrGLjn359GMmNslXvO/I7lMPGapiXzMRz1wRBmG1xTnd98g+YOKRk/DtACfNYIVQub
KfbRwJ6QaSHwTYsHkWcjPppUl7ywmTsNQEo0G+Nk95XNyWyDky+vBpknA/TlcvJ8+V1FxIvezj8Y
1XZhsfV3iQtcDzerjNoSUF1o2qD4AJNZsxXKVYKOrtUQbnLNFxaX818A7j0cMHwhEySY1a19ELHv
5rvnr7VBy2t2Zyq7o2jDFmluiyau2oTb2tfGI8GXrJl5zOzmcJkmAhp5hw7ioTiYpASeE9EcHr6U
v09R3F+1g8Iv0Rp3clCsP1CCxjGAb6kWcR8Vvpo0fvnjpCZDNYijZoUSvFcjzshuLLctVAHiqL1r
2pvDdfv/J36pBCWoPd5twZCOLr0PDzADcfFCEWmeDsnxw7hDAEuwNnuoEWEIBH0LW3Zw+TOfqDK6
I3JSIM+QhlRitaq7EoRZtjj3h0/cP4oiHeq38dTF41RMNU68UtGqi3TYzDbaUBHiMJ5BttemFMLg
/O4OgefoqANiF3iWPB2EpZNTlDbQFfPV58d4HLMvV0dAUN5m+8CEdV//WfNsLCiuwEs0UESrpmu6
M/cPaJ5qvgKpkhjeJ+Cazw3uPPD6CKKH7e8K8u7DhFbtgFwzA3xAt0xBVO5vPeLKXYObo0eOkchi
NjUMMZHu965HJ/ulBguS7a9L0oMuZg7F1x/iETywwk8iL5ysTTwjpNH/QcYwo0BZxmO9h4p8IL8c
TXtTAogPtAqQXPLpwzG0WYnSsm+FohoAFvFtDv0KuYC5rzzkqHhyD320V3IZm7wj4u3aFcJXet8W
nZ5L2zJG0T6CcYX6NLLhW7cyzcuTuYCu5ru138Xl9Etb5ZkHWLZMeFpJdLgWrDsKyFhbSuog9KAK
qDkHfSVTSs7WCei8jGYsj23e+Zn1M/zctfjMSZrVVmfg+7o1A3Jie4WwegruB+ost0sPNMAeY3QC
p35zdExvT4LAv2cSm9kgdakuSdgHatAHDBmTZWleipDdRUUeb+RxPYNRUfefb4BuoumjTqDB2uPe
dB9oMQNM7Wjlg7Uky0ewDGW93Q8ANb1+yy0FRtBepfcr42kKbfW7QFKMtWOjZLZqgqXbLgg4BL2j
SrLO5BKQA/x60JT0S63eYk4eBvAUpHpZDAeu3b9m/i/LXTZLdhYp56y+xYhtbX/klT0hIMycRmM1
fQyr5sYu6msaMPDLtnPY3CsV2v3kVVm6Id3ye7BAySBk6mWmOGG1zA2NJG0wA9bk+vsIzEuFvwW3
g9q8KrTrV62WAEZVK32CCCn24XYCOriwPeR/g2lrL9e6g5YuDV8/+VnCFCmmP7PNfG2AhFX6+t5I
DucFmg7V8/ALl2/N04KR0LwNK9TOANONKuFTbmYBDjvt9Vt4IgxobfY5FpQyHs98dnIFKt1NhxEU
fxR/1CwavEljNr4lnwgAT6aj7nEiY11j0oFk3oV+Y9MUY1MdvWvR6nPBcTblvDJGzHjJM/WjP59T
R0f8gyipgUe3MgLhISSMn12KhCC2c01pvA2DEnoYB1QtLkXYv5llaqrt4mfQKVs43/tzU6YETd31
60Zm4OnqKwjplFnkmPSFIhhQkr0cx7Kfj1Wg2nTGHV8iOWoXD303TXcU69EHfl4Tp8T1M0Q97pNi
RfgI5q7JmriHHLIK+WdtLSxHwH06xvJy9ShV5BHyLB/JGkaRZ0URwbKO07CfRpq6EPq8OzAHFGFK
eg6R1TO706ZnmE9NC2nw/NdC5ylwlPMv622Q08xTmAAzIbka0OsIPNnGAeUMqFCpfXsIyCScT8yN
GYU9AoUrMpvpjqBpsQ6TzF6pVR3IGJUOnx018cdNUNFPoHy4pv5k70YqWYBuIoSQCFvh6vBGqXVP
+5WwUZrlcitPeLmCgtzS6aR8yi9M4F8rq7HugxcO1Mfp2KNUb33aQVomC/go777bI18Qzf2j4i5r
iUnaC3CuBYCSBaLyGrYgYPcwq6Jx3HDfo63MYnYkDgpJFXtpQJpWDv7hjWOu2mRdYel2T0/WDS8r
pElQ0VA8CN4v78Gi0KoagueH7zB8KqSnw2cl3MyEEIaKAJNm/T0tYv7pbv7QgjUCyg7rIQS0yGui
13motnVSdJm7i1HZ86Qvbl4lPlXdzU3wBZCTQTygbeadAWpMLQgNoF6ldwnLHjG/Zj+EhcjYXleW
oLwxX4l/Jkt2T+eYMGygq7wee9/7N1DBd6rp8+/+SN8A7frACdx3apSEJq7jae836Mdcggs2qHhC
C6ULjH7qFKHkChA/WU9oIjVVpywSSl3hhqCHmFbuiQh1Y1wqRkhJS5yjYiAcSq8HyptPXCA9Jmwo
Tg76bP6FcHgkwtYhI7N36oHtP3xpxmd5Izg=
`protect end_protected

