

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
L9EbKuxxzV/09pnAb0OGW9DxPQ+o+m/MvX4x5f3JCiR63+KWt2eYB17k+9mGgVY+K1VLxoYz0z6V
YvlDefublw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
gJD53XIM6IXGcoGao7b+pChhlJwhGxOuVwSTI1iU+aaEVIG37JelabzUSiGlwgboK2Zv8N9/EzBK
Y9pDSGcMvhlTABOa75VEGmta9QvVzRVMjXtd0b/jrdUkZar600zvkPbB8+QESNshxT7B96klkdIo
XvMdlDR/SEQxmh4Mkpk=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
uMh613zg14bfl9MaiMXKdALr5q+gvlBiCCfJpnudkmj/VEzNaqE3gABSgWbIJEk6l3XEblsHwoSZ
2eueijgOoGBjZq9eDXqLeir52M0Z4RoybrJFqX7YgYE+2quggoW8XJjUPK7bExWH1Wd6un6XRwZo
+XQ53VUhkTgctFKNHRr7bEqxJa0qk8dm+fTRKVmCc1Tr5X6rd28yRrr4koH3+liBwEPKquwcMKJL
zK5B0g+bSiHJvGXlQQpKzQNF3+4MebcveUUQPOYG2FAjfRJs1t60dgE73q6y3I1DMI/3MguCuvoX
78TA3nOFRYGLkISVFXDX28xYA0EnciH3BlzGiA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
2ADp5V47yVkwRII2+UsRY3zvclviExupZdil2h787eVOjYg5odQlZCOMnldkarIbxDBoj52vjMGc
rG04pAKa/Z3oDUnDkDe8ZMmBI29kynugqgc8aGxYPVKp3KD8EvhnicB6/4Tt66g9A8WsjHtxXLuC
0ImlGHU3T8u48JygeUs=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
s5k0DDcwk1Yhkk6mc4rW2ITc+jBCojX0QPFrzARjmvIjcmc9EJT8pAYSdJK1ykoSIGmT8u4U6vaF
5pchZ1NWV4+0T78Lu7ir0M6lHPYDFRgXZTR6CNdPGqAe+Si56W7NnXEM0Yylf/w4tAQ0u+05yvCg
wK+mPCq/91Em5ZiPcvKOHOdJBSTTkSYC7/n0QNniR1mBmd7+dgsFr5yshClYY/q8HngDDE/aNYfx
P9AT4ECjL+OzARXCnbTA6RjbHEjVx1ewIc83WIXkwbZjUYAzp9rYNjFdx68zjq8U1XW92RXAEXCc
AYKv676uVGq/WAryucxGApaihL/izu2+HGUsYA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 30640)
`protect data_block
6uwM7pdOL8FOy/3Eop62YbeD4PQeAmAf+W88yPyWlIOlazcmoeArt//RHYarMAmDlKF5ETgIwNlV
/Csv3x4kB67Nq5a9I6rH0OAcIPgSYTaJVhjtWMYKhMeuEyIHcAsG7PD60iwt9fENLO7kYlTgnSLP
/WvIx1reYSsKNL/hFaQ2GX5whDtCcsF3CuBeG/Q/bEDHygTVv94VLAgvHxNK9rj9W3p4FzhTwjUu
xW7fX4+l+W8aKUO41J2aLWP9AYrbs3nZyHMjKl6JaT5mtH8Evi2FI/s/k+UnTaa3O0eAva/oYRkv
BiuJkPNCPJ2C6MizC+WGzlgbEQ4I3b+rG2GrMQRQeBWJwDzYwjaCeww2RrHTDI7BeTIxUkrEc4cA
1sMOEHW9rlYKeCHcyQZ01SoWBnBYsojYp8hf0ZoGdQEtzuj293q+dnmg42+k5/u36IQ0dkqgYhX/
bo8shFpqlD7SAGcLWdJE9hBaftMHP2JhkHuyrUF076SvgoX7RIp1EBSkr6cnne9RcOcQr9vObtFq
Ua/SGUMPtXOjF10e4EEGliyuoLBCDBe6LevQPO5KX4U83oXxYlCY6zfrjUq9gKmrxga2VYBvyrNH
zkLQbHXMMZ9wrOU0UATi5uWeVwmJeadZ42QP4qZQ0chOl6CzIjKpnN45eJheKzE4Smm5dkOMsc9X
hBS4FeCX7Zhz5UVHkKPbnpo5Y9lTS3R9mZm8Ez4IyEtmUqZgiTyUyQ0JG/oYXDcBVvFSnMBqr6Je
eO/SZpXVP+HQ7JofgEQJtrhYrw4k+zg6MZCI5UK6o1yKIY0F0dDTAmbSvVwKvs3SCBJvhwBopQ4E
LNYzJX+IYxyyBIF+7K7Q0QwHHOC9ji2LIjVejsx8n4PJZHTjMy9V3w9OL2NdqWG/u0il9FpBfVDa
wTWWfbbd0oSsnHxvm2aidN9xvRsYeja2Ar47jUiQ36Feht766K/ldlVUH2wCtbb2FXcHZiR2FQyH
64mFPcJY1DlKd2EsHhCC6Dd/UB0BzuXZyZwtG2OgHttBb4ZiHMe2/YfofSu/b4LE3bK+h/5Ct3EO
+BhDCTHRcw4j4gq6TTGBQ47Pz8smqouV1ZrCN4ePjDvBMmF7lSHqzJkjvaXEDVGW+dqAgMU8hfiu
qxbinZAl3x4/OtPl5LvsvFtsOppB6Y8Bb6d9ejPkNAjPpPZJU09qEd8Lyc5EFKzNkb0hZq2WwYd+
eis9LYyk4O4XV6zZFhsHj8o9EP4hCwVn4Pt3qA61wY6Nz9LLHy36Qoq65XN3PQJBxLZzHW7KEg11
SmxVx1gN6BlQy1Ky7pzL8GHc8MzVezZQ0eLycthAIW5Ovv1nocVgV0inutrPZiPjDwtpMUf/fI4/
77QqWZAAYJcesvy8gH+wc/JqBRUo7+GlodmdkMv08J9YJwNvHn4TgexXeyAXyO6J6nh1icSkBDQo
PIodVu1PSa5fzvR9MVZQXfq48TRb63mu1tBPFTosPviRbQii5OXyikEeRFcpK8EoDQrct6eaDKY4
QmGwr9076Urj/668AlItyyGbGwqhQ/iLIhKuqwqMKAaR4zxfbdYRQbBp6xy8spZcISz7Xqi/d64p
CujHHIuJmZyvw4n9jvj1wZl5UvX+3B7OhSFwseGNpkE2w+2RqaG4qC7vaVNDyEsb9mEPjxXWsHzK
9JdaYLpmpOYET2axxw8sS/rkGq9mHkznAjItf+LPaqhSaeq34WkBd6qoWWMZCovcKDCREHuJn1/E
bYUub/Y+8QAC6hWJb6vBv2SfsxS76Iukblzi6Q0tedA7qVEr4b0fi4QBbGSRdJ06Dkyd4z1VDW1J
NqEhENRmdbmCUrp9I3yV6KIwKQv9zs+CP9AuZ0GBotzc7viXiyV6KtUxxDeS48HLTjKrSG/YDgl5
SDAQAXL78YQIGUCWM5CtFT2SV3C91gTq0+ozWdUaEQjzCoFuGr2eXQWsEC9kWvPD1DMHJR1FchX1
Wiw7FUAyV6/tSIX7FA+1R+BN5cdDmqeAvp7qcF8+nevaf/yl6Sijg0T7YUiLqK+jaihEiPnf4KrD
tn1fpTMFO7KUh/MLbphINuWTiwHRAe/QhLTHh4w+STNTUQMaWMck6VLGq37eZavxUl7qph4iF6vU
OinP3Pz/bfvRpvfjVvgUKWTNiJH36oAJlFYNhYmz/ycPmVrdHiZbyYyyJIWoGPm6k3I4sn2HKHtn
Zh0N5Enz9d3GaQOg3Jz3ZG8eQ5dePo3sdPX4kNKFfz0UjqoGrF0DR8YmQm2PGBa8F/oDjt6rMP4U
MhTuLGlBK7HzhatGcM5vmPd5xoh9wgY9YYQuRFe7kNEuyW1Lr07weM8Hmz0IeYHzQOT5sBUk+UBS
Po9j+yOOQ8rI18gqm0aOHGUYW6x788bkpIEAyuXvV0aeGRCRSJc7uXLQZEQLedLPr+akhaCsOJIA
9J7609QsPO9Mhs0C7RMZAo8GWdnOd0coLxIL55zHkuS3YIw2vvfjU6Kb6YbaUz0nH2VoZ0pxVL0A
2iY85jY4q/PyYgiit0/C8G/2hgtg1BTsH/bptg7GG0zUPdPN1MNlHykZ8yfmWGkTeyqcDln0iYti
sqw607eIaaZt1quQXhWhBrY+ZXuePOTGE5qTlS/3kDw2WluXxsei6hzVKbjCZpxVftShRFtvpruB
t1G3wGhjSW/uIRa/OX73Rw4UE4kaTddVyuksFxp2O+V/Z6Wgln+saTn8I0ynoE82JbrcfR4PpvxT
ZqMln9UmHmybeEh+3uUtc8SI6OX3EFwICs7WOGnIntMywx+KHXaWK1XqegQep9y9+OTNYvXqN0Vt
2gQOZvdHBCZ/cJXPEBXFBTevhyvQTcjHS6mIShGNAHKu/VGRP0nSJD9GzObTF/EszR/rioonkpUm
k6U44BQRptwiPowfE6wOE6AHMijGogZAKLrLTUuFl2MezxlLz5Y/O669Ji7horwnUF+ZKYs1GOvH
q1nY20GhWi8ufzm5NMkwbD6eikD2FQmyhZPv4AjQ0gQj5DG6A6QDqBlyd+fIN/Ogs+lLUh7NX9Vn
EqDGhJNAektGCunfUnZsGx+dBKegXMh3TepiYe7kqOkbk0o0T2af/oQlw3INueP9YQ0Ev1De5krV
Kxg+Dso9amlwh88y0ydIu77Foe3l0xV85K2Gbsl7lVRjz/coz4riR6R8+0o/54/15IB8Mb2rONnh
KxLH3xn0xxADvr2HeCJUZWeCtmw/7YsmPe8x726QfyNu3+96nhHAZBukRuzdrHW0R5WFFfiA6mPQ
YQqPIQythkBPnPRhSUg6NUeuWsSSELhFl+Fu+Fa9PS9P0mX5RvpU3UR9CPOcO0IJgEz6MiQ4R74E
LyeN1qeJdtOYd8y1X/5UHaVQ8fxXSZ65xxLQwswOdpeEdTP5AyhshiN74673mZR9Xb8lMwRw8LrJ
sYZ9QiG6C8s7MaQYS+S5ROVDXPnDub0VAnFYCzLjMwo1OeUA8Sc6K/AwWd6DVxJghKPUyXz7ii2V
84druj5CIIHSZeETpR+i+rPJWODPE8W7Re1pXmz64FFyAJFlxk2Onxr7SLFZ3qhDipQxs86dc72b
D2A4fJU46aKwO+YwEL0i74X5bLHoZlCEOeiLU+Gq/Ij5Wecs553MOoGFQcVoCDijcgdiB00WxYFT
7CKuiTqDZwBRfvnzo3Kx+JoexoMzOGdK1KuU5Gb/eTXoDJgYh/OHFs95OZAZ5JYa+bQfukP1BXFE
RV1BdmJdLs8Q3kLx4U0v1fQJDhaalgTpTRp04pHwuSSqHMBr1xAhFx6VhEHy1Ys0hIT/0maFx63L
Tn5iNZfaGv4vhnPgc/g6P8Id/dFQ6FwTywoXcGF48ZK+Bs54o9Ya7kBoNUHde9vnWi2Nix9PmYld
dDqXGWr3KIM7+M45/HtB6mBgPZHn9qCtJMjvhXv7NoNbAiFp+X2jZUeEx0h1Y/Du7CNiOoW3o5hI
GzzIw2p3liogotFL6BKD/se6OgDWwMyGoUZPh9VEG9uBxDHceUd6WIG/TQVbrC46CHImX7VnY+JE
ejM1ltmS3vcqHeuM2wHAGuwJfvbp6bCI1Xk6dQfxQBnl1lQUalsRwIi2pe2LPyQ0IL0Ty5WgutVw
8DwlcIT3TGVdoFMXYMmfGg/yMNlFLxbbEqldOE1CWqbZUOreda0eCFCINxC4ljFXhlh65uloIhto
EIXHfXj6pl8hT4T75pqChsEOmI/754COZF1iixQJLFDqOFeiAqbwo+QY31LvBmFQB9O0LLCFxW5H
NbCey0fflilnqOamIuEVBphln/HNvo/aBnMezN+obg64s4J7PY7d9bHII0ZBxKIp0QpKiFTU+ay5
HO1JTLAoaMmP2NoRL7sB2k6BxyC0TVrd1nHTwkSgygjGwlOg/89x6IcYAnch1HiZZZ6VoFpjo8gI
7WhTostURxbBu4ZTBwOReY1ACcEtmc3rS9l+1HvbyZRc/9nE/hqVY79erdhPP5TlzQJ7bzyo2lVr
wODdrv8ujr1Rt3ZoDpiMoHPtqBx7AhK90shWxaOlt1Dcyjvh6Azz4Nizky6ekpNLqVZHCqwF6fQ8
9OBNyXmYCxUvTNNVe9f5qq/iFRgEa93LWJsykbJl4mHPYcQBbWIStKI2r/UOW2hgBOrsX3m1/7Ly
a/tI7Q/+qXq8GdjzXCF816wlF7G1Ph5EpRaNjMBAL9YgmxlW60KUmsI8bgvwkb3f2OE09p7MKZGx
keezaxrIQ4XmV4KcM+Lm6Gx4iBnbD86T7VniItw/rehMdcWBBWkrIsGOSfmCyIqPTWoCmMXN4iOx
ZhVolt7xv8QAqpwR2DDsEwAWrMep377XsGmXQm3E01XS0FPiLxJHYGq6EBTMEGZ0d+r36nPN/t7j
90Lu1SngufipeflR4nK6q+Scqy4mMfdc0QOm4VhWvHzPcJDKzjec+jUTt3FalOXA4WkWOSgtcQEc
X8Xf4uQdDcu0kJG69UZ9ynQLF77bKsz3rpeNRzUZ7zP9gduhCCufWdmROPLzF+0YDOsW2aK3ZFGR
DYSUogGy2qQqYyVTb2hpaQ61ATXddn/VLLxRLXTMx3vdglwcYSmsdthr10piPfmygVHuNEw9s0uJ
65OZ9feQnGAGCXg1tbOANDhF17/V0il+inaWIJDPMxsw7qZuJol1MqP4GXtxGZ3xUUtmfaBc6u4E
+ZdlePvMoCPcAKWECsqKJltdeEypn+TeuCs9LCUeaDpASc3mIcQQmla4J9cGygtBgSLaDwIuD0P2
bompOcoUtsBElKogE85gbhQm81xNJnPmmQt/JzvzHvpKJobqPiEKn1Rnt8wjTVtH1GVeVuTGFI11
qQNIPCupqyk7+orEoBZPMdtm9XWTp/ya+4HuAZ3pA0CYqlpvCitxZ38/vCqES/r54YcvEQbiDY76
XaWp7AAgEHzGUP3Ll0kxDknnu2xt0I7t/WWLfnL96It7qaKv1eEex7x2Cui0BZekkzjfMxjLCOVG
E0TNSMQydc6cXyp/khuVeA/N4xeeHAvzgDnnI9+FBEbHEC8fVWCA8kQmErZXqqSE7Dkr7E+pt8NX
45SILFpWFyMUljG7FHsfQi0iNcoesGZCfANd9m7dEOZNwHzrQ7AQ4iCgm4SW0XSU3Y7bTTX2pS0d
gzTazxkj0wXbo4N0vJL3TpPRkSKJiQvtoY7Svm4plDLKzi8o8UGw+aSBlcfwH9HsV0v/r6Co6DtE
Gde0vBuQ9vGMjy9JqCiS1gfRXUGmmaZ9FUwEXdqoe1ES9+AuesCUVaHCQTP0IuT2PgaQ56PR0MK2
fnKsnxYDlTDnw8+QJOu0kon/t+TA+7gHLhGcBgKIh2Ql7L2q50p9A8Lsm9S/L0xNK4D5+rd8sjK3
KajWuVeQYBz5zNP62GSdd24lFo330ytdTwLsA4CTABh6shOqVqjiKT8B6bvanon4CePnB0XMBbKA
G7+uCq/3G6thbF4r1EQXRwY5bgZUduvuLNBO3+r60InfmgLpsVP13epDzWsTk3WzmsU4noYTzH3i
4FOfKY5EqwThlg4FkTJgnKOsVd77Pb8noUj/VQ6wIAQHvZUiu9MhwFpym2dMKCmQ5t4xzBTUBrfT
Xpij7oJ6kVTPOVp7RKAlTfvipw1r5oIui9ZZho3kkyE1A6B0SiEmGca83HXhBPrXeieLzFg9HfqG
Mt8LdrLm6rWw8ReFxa0bwlV350/TYxdb7AAhGyUZwEjz/tTq3WPwxaeR7P9jv5nl/dhjADtAe71z
2X4AsiwEkjlFK/0iNdCww5maEk6Q8W19h0hqLehVCJgqJj4T/FnSk4+Ja+0ZVyPHCrUuv1QfWobH
DOREOIwnIc9CHv4Yfi/E5nvQkRRvU/bUepeTKZLbHW4gcNJ25F1AZW8seabl4j/jdCips/HFvU5F
gf2YTKKA1OrTytIWzu7XkVZEWMsRdjU931Zc7d28TsaEJttYJ1JGPDlv0tFXCwf6T7TpRkg37zBt
teKsiMOO3sCj2YIJ7wpKDX10KdIUjSEuntTaD3waYEQxZAsD4uvwIs1eUfUXxi0ss0IVFzcaQkw5
QpPpZiLjSr/u2ohU4MKckI7Xn+jxHJuKSZZ+w3UQQ9y/8Hatlo2PfdEJzlOX0T33a0RiDZX4Jsap
/e1ZHKmIDpCWOFSGVQf8HUHZaOs958c0UYh7GzRjo0RwjlgMstgo+GtS5LCRsEqY+aUqh7gbFoXy
kUyrVaJaoTzsTDGi33sQV/1HQyiTWMMZaVyYpIM/ttOTGi4Rabl1mWvsZ+L4VJhVyn5L8/gN+MPw
gk9g+9+KQNeRrXo4XAS9DOL2YIX0tKttMj4QxtFNbWQpYsab/Q/L7SzHB3SYmO1dUTsyAWUqdW+r
m6JG0RSIQVAHvLa9nK1ixwuLsejEWuvx7eA2dbFX8EUCORNQMFVKnA5MOkm9bjzDAo3cs9sucsIQ
CPz2s9np2//58mLh17zjXf+Qr4LQEu0cXxIRGrXprPk82QvJjnrduFBGSc0VG0Bjvx9GxRdLblKA
dWoeTZZkd0ZVbgox3LK8wlKSgHjEq8//X6ks7kWg43H4h4l5wPRy9weoumbrRhQsWYrAyJxn+1xQ
Oz7KwnbmTagOumcglqN24mQxE1kl82rdsOqsL6gq6wswpdHeFpebS3XWmwLhRGTzffjdzxwWu/Zm
Tf5jHoMHc2eTj0AVOwgjhzPauAglyJO65RpUpPfwLkcLrnKv7CPEAJlTIAlBV+p+F3Eb23A50guQ
ywhb9MjCWQRhRGHn1a0+FOXqpDYfbhKpxy7Gl6my0zdBaeVe7AhAyA0pm6oa6yU8EKSgzWfwZOgf
lZRpAVb9V59k576T71QAFE2s25DqKEhdfZVlIoQ1B/90p+2QU5gD+RihgF+fxcdmX1kLz1m3HjHR
d2F9yI3R+UYwZosI13eBm+62jlONElDYKPjibXBPUifbyQVc2f58jY1hwqc/nb+L000ErLA6/dLI
eOgJEf6RGutOs8ZLIHJV6wyHEC/J+IgvMvK7zSJyMwB7B0m5OQG4LOm7rs/QBLHF23kGnjFai2sD
/CJpE7D/fTFXqhEOQMsou+zCd9IKi+Qxl0zLJj2YlK5L1pXaEJHGtJr2ox2j33nEscs6Y8Xj2zna
fGPLBsOgPO2bN9wGRNzqpUCT9Du/Q2+EOSP5Y4tg7qcTsIOfmnAQNqk/rbNnM7q0uORoaMXughFe
9yNdgK5U8qedGt2nETDAop7nJAdWDSNU2gZ0d3zRAUbntWlF/qvu7/iNMB0YSOUNw3XQlodRfvKk
etjo+SZhhx/5KfE33bQABT3+YQlr+4964NA3z55kx41d+vsmSXtGB18LFBVLQHbRTumzAiBhZTPC
s63hATzDWw4tAmMJDQgCQQjwOA9yhuJAAI7O+R90XOjRp8V4uhkEfEeBK/+RzOolsC0F8L9+zRKU
WfU08X/wTH99WWp98QkUQuaYlDnluT+oAmFctuNHaxZkZByS4cUOV5eSpkT0JpF4X2RdC1QdvxGU
O/cklAzmTx8zTF1+8MFdTbIsTtAk4JDaeoZMalzd53sUUjIkVGt+PAyKJu53xT/wkb+ET4z4YMcx
WDlEmMJddLvFZooVH1aGeNPvuH+Z2qhXwxuy8zJzaeyDUo8CR0qIqhL+G93apJoTWC9jODBWe/CJ
hj7qWdA3hjIDbO9WD6yQJH/ooK1jTBlrVPH59BDsUzQofTYbpFLyqCZtxjgk/Obbho2unnRPpA4H
OehZ2sn69WEM1ITMcl2NfmBEFhcSHjzzxM3E1Scqnfok58WVB4PaccXc7t7IZNAaX1qSFNaeLuuq
DQ1e9ofKkUu3a9B6kG/vhcc5rv7VwaJEj+021m02oiIygArTG9THVtbIq4PBLjku5j3OAT5uLZ6L
X66Z6f27+INAGUzuodFCgx127nrNQ54wJw4e/i+pQL41eWBBFWA8Zzchk3RTBKjoy8+hR7BFuI1G
tncwxgm65SvdQyKAqq+iokfwK8HujG5i/9tXlsAK2gux6QPdvcmerd3dhXtBuJqFwd2R/GzCtsjF
rHAKCJbjC09yIyaorI/uBfQgXd2+dOVSbF3iRX1xEyif2vJjprjViax7YlZSpa01Kw7r6qoiNfxK
5tDnP8godKNtIl8JupTOJirvICz6glfW+aChRgAeQNv+fnEQvF7Kkjz/WWA++gLG5VlYGU6wFhdo
FQLzd/JQ6W1a3IGOqnorFJdH4zq6A4hK27kexg2adyie4n/BpOU/k2lzi9gHi6JEZmuaLtNr1fOx
g0sx+xRgC4HsPDJeJtDPTSR/a0ImgPiQHgguWNETMoEVwa3+GUT3W0nEuFquizeKg8WgtnLcsc8y
iqaVf58Y/9sGp9yt5uIQTLrPF5JX8x4fOiYHUPrNzSGF2qnSQ6RQy6+FyQZqdIhVCrw+7WBPg0xb
Y+2g2lbqRQQZ9YrZLW5FlOcEt7LcN8nuhcZA9qmyd32j+lPILcI4sPjMpMnB9I8UeYqR9soVi2sQ
b3FByQWDohIkCMoijELHlhJkGFkSY9UHbbJc2SDiROQLf8/2y75zhTzrkfGnspI8wD5BxC57UO8z
2iMTnCEZ1wzEP4iQrXIIV9obXE2oOCHVj3Ek6QvJTADSSjJe11TX66/TwxCmXHm9ABuJGQXActnM
cu7xqGrM49Jo9K6eXZelFniKy0kNeNIwPY3szeQSg0HP6uE2R6s1+m976ph4+rZCVYrUhyo6fB7f
/2sC+7G2d301HT7b+pX7PcgcUjkVp517FLpPc7BOHJpG2XnaEMD4RuaQeEwF3fECloACR/gWTFdH
BKpIPeTl07XisuG6vJxrtRd7E27sqmJ+6L7yFewV/VfeZMRDj8Vk73O3ROcxBP8dIVtuUjle+EOP
YF6YM6qVbfKio+/EpAL+k1l6s2gMo57dFVnk3OYlAg9+yQLJSXwahYWbphWeveGgDwvutyWpF1lF
QMKnEgLaaJ275RkzHiWRovOegDwNrSjVa3g3KVnc0EbgnI0Z55f50tFQk3FwzFwv161oy8TGA6A8
YXfXQfy0susRSm6yk78F3jiINasmHuARlaosidQAeUef36Rmo8FZC6Rj7DfoMIASN6jhrOu76BpM
OE7USgGwxUnaA/GRO7UconyFRMODUcjfbKS1DYo7PlbpyI6OP6gl8uqrQkwtY2UeugEZc9z7LqH6
PFIa2eSsMhsxFTW+71EAmnBoGdDWtYyiZbwebg6QD+5mFr6VGb48M7fgYMXCbAFOtI3wkSYOfdDm
Mb9TN4d60uljvbTxa661RV4Xl3gN9myfII5eIUFtZQkj9dgDZ10oVITx9pOJnzXm4fHjE2ptriyo
es5aqtR/bC1ZVspmd5aDpzWu/YNJ6cJmM4L8UoWpR2onRzTAqFKR1HQSMGVaYlf5OZfvEtobbR13
Y/UR4fq6TTUkN4coxWvcbNOcnnaC4az6Jwx/zThDt9vCKdWN3zv1sDqFdgg4kWaH6cPq3aOBRSIn
U7XVxDZVNZTQrOALREycLInZbW5zEh1OSAlVj3fIvVfdarR8yMuKnzp+/O24Fg03fV+tH2mm2uFJ
FOCyu42i+/m5uISv/0dkRb4TGzZ3lyKNx6/l+okU+nPAdQslhCJuQaADD7qIR+lOHCWyykYeEHZw
lS0ubs3QIetNk+zoWDBk4Q5s5xEZ81qFFVAj8k4zN6nDJAhLbjtmapdNQYlkmytEqip+OQyZRnea
+zY5LZi/MIyIPIeSAgymwGt8Ch37MVmDi8nH23l/1mAzd5Lw7q4eYpFvuygxofRYyXVJfJn6b6eE
ZuoNpw7Um7rE6PT0kUaJktmiM/OKJSt5WWnc9LBYuxS5o3etJYP4y3cGqD12/l0SeH5BCauVfDQ3
ifsqk0YAsEnzXe+n+Ku+c8YiQHW9gP1kfnN260WvzxdWAePPOjvdUB2e/BrSAEsXqnuuUtTlaoRQ
TSAKLHVLbMbHoVlPsP2HbGVOSkEyOqvCpv9HFilT0I1KNBMSLjRQS5J1YKffedrLx2N7u2+xSdd+
B45B+SzNIFIx8pG1OtZjq1DXPFKoN82tHYv1R3TkoHcbwfbaNWPE/RLi5ds0kp7Vj+/VYsI0TT8q
4oEmODf334etutiKQnDWlhGInQdW5ghiMNd5Hl1lix0P7N5BaX1EnYRWuk7pjI+K3IkMaSWQyuDy
DX0akIFntABg2HWa6cu/Ee+aoFb8vBSEQbIucGCaUl1RVCqXvOwNerXddwGezQU+SmWPRoFdLHDv
tjnknZmpRSuNR5Dl/2wp3TDVUI8PRdadU/DEaVzGZSgV+f6nV8CB9a26rQUlQy40udEG4U70wMoP
DGAqPJr3Al822eZmV4igoREr8yTb2Uy9/+yxmb7hVNmdifToLP7O+jc5l50dKH9kKOVsTolwNCd+
kwwtS9JawqYHnWSQ1f0Jh3EVpiYl+TbcNwLuBatt1XuHmi++8rqkzyGUOm8V+FJytIdaPJgEWCg8
ESUqsotgaHA8NulpOOXcR26f4OgLLqgyjeQLSY01noQKpwnS9DfQP/zvswT0yU52yXEIo8ZKOrRU
MxLUHzBhS0b7kSMAqGxHJ0cNtQiUvEjkr0I0AFvF6mgrMZ6xEiC0N7kEH9TDeunjoXWViBo5dUZU
0BQ4ynJV4eaSnJzkPlU3QHFdxUtvYtOXZ6c61PW7qHqikjAu6kR0fKh6IMvIcnK1Bkqepd3PfECO
6tBJRP2x8N2zszV3H+4vOrTBmSHgH3nXYbLkos2mH2XGdYyk3/h60X+ufoKY/ChgJpDtJAPp1eux
vIk9eRmh6pmX0vQe4yzIqpR5CkWrh1qtN2T36vnq7XILmeGrQgf/QBEPxoei2oG4Pf5tSiFDwjxK
Vj15v7qXJBvpNTpbbDH25xG/WhrLalCJLK7yiGcjkAGYs/CdqGocxTQVdzuDJ4lNJhhNt1ml/jvw
P/YKZIyl0jL4EQotQrPU8nmp4f28n+qYk4AuJ5nhhBDbmprT5iUviSo2g3f5gf98P27/tiv5zRwr
D/kA5CuF2+cx5bcG4Twsb63nLqNiezJjXTMZgGg4pMwJSafb9zXwoCDHCVNhaOgAnuaZyrwKW4CW
RLUilqQByL8opoQccnqWi1S4VOHyJroJcDGJe0tK9X66C5fIBnn4XyKfGMD/KuaTp606jWknS7Qo
hqFU3zcuWXCelt2hkBAL/wl3CPz+21E4pSb1jiKJLjpRhvPj6mTO6BkUEu+FeNcc3zFrMiIRWjb1
TjO80JyBV4/h7UAkDzSWCuEGbZdBScGcsi5b5BeCGV4jX1rO+Lo2KhHYZko32U1WbLdxXUP8oTmD
JlTkX1MbbUsBZP6hS0JmJULJ7ne9r2mzZvidT4u+16CtijmyNOdI/x3Jvf6o3+Qx5KlcLf5/06It
iwAjw+vLdmNIZ0mzy5V+qOHDAfohTIrSM+vm8ytOs1LDEqsdnAEfdFcVqK6c2MEaTjImBa/myi6s
zEN/E76THevNvCGMkSaGXKAQBootC8X+FMBIjFcuToB1F0oeFkqUZS+xA3vM0LZp3czAt6duuIaF
hMIi6NKRU5g6rVZalzF6UUh9Zliv718sbnVo+SzppUMVVSBguXUuwhfl7PBM7koEFqBAGmtmk6bV
ILTBzCMyfSiB72yTrW6qn8CpRc64Y0u3wvvaf2Td6uqheb6UeuHfE/AZm5xlXVBsPRQU2YqQGqAA
EqlAk9/Nd6xTDhbf7sqjM0ZFeAC67oQfLR0YNdAsi6gImL6CrluyTqgH1AXkfYkYpXpKMdFPy/27
NOYXjCatdzkQOwMNYdz+CbsAcqO204Y8A6CmeXCPwqI3DebMPg0VPR0A5o+m97K03X5CJvByJrqr
fAZKchCbiQH4Zjg4prQ78d+vZ6hYy8cwxpRh3t8byFlGrx8WfYSZWg5V1kSgDq+LeHQjuw5d9Mhl
qVSqoSsUhSuWYnhnUAlPOwxebGMz18j5AZxw31xiGTjtfrI1vCipHfBqaHim5Af2n8i66eJJMhVb
aJdpYj86Uhcy9NaWnqAiC5WU8lG3U6vP1TUNhJbVncL2y8+FJqeh/BESPYXwoJF6c35CHbfF0fs9
LGJpad5mgT3BfBfpDPvb5IwpsKa1DtyzZi/iCmSYT3V6PibKruNKJ4cwTRKz6SRK7/g6Q/hg4DYq
tO8QF5gPhGG1gWe6WHberYnzK4kRSUvmgBlHtj47Nj9TsH/5cmccG0DLnC4BngbS2HU1pEmKeGIv
XEYTbsFq76BPpQYJUHzqRmN3pPnzBJTqbouAVcBVAnX1J0VScu98X7Rx3VI1M8AzPgzMnJ1BYFAk
sKMMHZDEroBxsqJg5iTOvp6YOjQ2AtVXEiUX4qa9jgCzmD9fI8X8QEhw1ZlYSj0dQjkVm36ilpAj
poyFHZol82hIHFrKts5hYniCwRH//9Ve8GI6aizu9+Y5o8BNKq/f54FZ4qgU0R/qIQKSB1pWuU2l
hkrYYVjq2rZRIwEyJ4z8w1CYth0eh2lJpS6zkD/oBnFVc5+DWn4q0XED8vjvdHn6x6JSlI8enRA3
A26PVUwzfQUEUHAxyND0xrvNab90aTb1jISW5iL2fj7gY1SQW5a3ifmsemHBwhsZGZIpP/k61ef6
3//j1QLx6CtBb3lOn4zr76QtnN6gRZmjdAiE6DgVYByHyoHh4qroIiN4ScPNJmgLKQDu7X6H1S8U
Se1jnSo5IECKokOi2ym3aVysmUQLOIFQvWhMYqDRuhWfZk6TjJ3YaFQ/bVcnNlPCnQBCI2tWbhjF
DdZbxOBT6siMES6gneNfsMzJ+tubHLIVda/qgwfGd8Kc+QmT/qf4yfvLHSxnuLvplAreNfOjlcZh
2F3okm1yscbbYijGX3L1VMum55szx1pwb1fsrOYBpFlL3PkhzldUiVN5pnfrkDqZfY0hAYkzoMxG
48yezcjz8Yg/mJ4VkFFA7bGA9FEIICb41TnrdabBrkNiVGV60frAblDXt7NoOwN4psdlNBt0hSFc
uM7ML+mD+8s8SmXbcioW1ABSu0Qq1Ysu4JFdH1EcJPvTh7aRBtC0A4DagZJknBFwHixO+jrWJtLq
ipG0l/zxxPrBitrGmx8mabp3H3/xFZrvwbogK+YTrcznlKZBxYXJyrl1ANGACMrVCr5epxYv82/C
TQtQuTUnNHzQY4/af+nc9+5DM1kFtoKrQL+BlAKuJbUJ5C3s33oFDI2zDx+L+tBQYS239NbrIDHv
V33ii4qbxANe5q7yZMvmCNo/nAUs9pMz0j+lvxaHj/9hBsNFS+28ensLTuEtxkjSoLBneIdar8U3
ZJCbNNPyRBAT6tOZkR0BGOPrjQbcYnVR9IYMd089GX0nvNUF0sYrrtKFuCNgYenxKL4YSAaTNLxD
jF5klq6W1xqVfGBJf135FgsQVN6TdRQx7FS0yus+jMm1cs6pqXHbJORj+UNT0D28dJtAvtq+NTUy
t6HDblWqPKaDxi+jG1DOwzR7mlkkHnnR1GaOX65mQxynJxM2iZ0K7b97ryqFSQNjEaUTth+1j/XV
RUB1lqF6WE+JIa7hYscvwSBEb5zEU6cMshdrVxUUC1T62/o3Xq7HkuaGcPwmuraCPEjeOCdx56gR
PDcN4nCywhbZs08ASQ6E5zwsWXSfdddxKT7MMysD3eFMVWCMz7g0Hd2CKMRKoJ6gyeKv/SBfd1jc
GNhmz0QiU3HNesqU9UnNN8iTT86+uPGmitfRGXqLMKDRHHzyUQ44NTDr3xnIA2Z0FrxYviZ2w8vm
5b40ZurGECSUAsRBndvS8qiryQikugq9J9tgFHTmej03Kc+vttLzjOVn5LYs+G0k5MZpSkP5fNWb
lL4o6rYNlp7tPMgt+DMincz4oZ8yRKGMh0P/fyn9SMAOzjR94G2lnA7EQcpu9sJCR72A8+Ig+/QG
noT2N8u0OOJIbQCfgmISSjqvfCLuctgBFNwZSAwoZYULe9CeLldyZzALfm4qvFL7TDlw5AOSMadm
XQqlED9qO/cDR3sg8AEOGSA4veZ4q7L4czz7DykoMRDrQodF806/ROmbwVGDJ5I04Zbadb0phqWY
cSBIP/ImgdQi/U28+oQpGxmCKhX3hJW8/psbATWj5MqrVlK4bI1512r8g5CsPFJRiGy2rSvKXGyJ
HxE+COKRCvgbaB/dTjNHlcdv+2vyLUvvwO1ssaZ1Gd0fDoPGFBkGSYXh17XJxTOAApR2KmESuay+
bYyZPOSEGt2ALPIcTN3fnote3x6YGLnGM1VCRxOdfjh/k+VAzccpf4k2tl+8m0oxIV2mSIUfHBQI
alc2X5P7kVEcMUFh5aormikkIRRWLL1Pw5Za7r2A29cMNhlKE+zZntjcX6sd/rha/VtCKSCXDj1/
ku4VKFXgiQVU16lYaVUF1LJlJysofXzp+rAGhGjnIA69/rjuMM8tiRxKzOfyAZzn4FmfgFfYGFXP
Zi+GMLLImyZ+Y4WBaXIcmzo+Euvrw378E2TmkI3tIICJQ6omA/fUZzQy5a8/pQdeKIJYvHgMsHPK
gXS3Inq6xsZyxS3LTAMeUWdPYzGIRzX6rdmMXShKFjrXRYkXP612WjG3mCJ/DMwx8fsmTTpKUaAn
6rRBxqHvQDwJBRgiXsktU2+OUxwzD5PSUvY0ewejhpZ26TsGeVFAt0XGePoHsLLE+JwPdE2ClkVh
IHSeDEIlAhPvxxJaUu0aM2iDAtJSl5Uu+4rG6sVQz3IoKodAq1jic8qe0XT8UVveaLiNsBfUigwr
E5bVBmQAwPQOhxAuYTp2sedQjd46PIYJtjDHUJ/SUxqzdF8x1phEKZbWriQDMl0dvo04uxIuy90g
WTipH3GoJIxUJVKRyCE18pDRtxPqluO++RlRKq6eqsDer0FPfdkjOpe9jNa9/V8QfJFZB+xgVvjd
gQX9UVTjxU35uLq3XX+pIt2vmuU0f0yBhcvOzxUWOxLTGmIggNAec80E3MSpfi5NhQPZuJEniRaH
MV1/iWLNV5rAEGbSVMVnIOWPKOusVhxxrgqIrTcCoJeRY1UdK65Y/6eTjb9r8YFULFoGgdQWb/aH
aLrVnVB2U7FjRLV7KnJ3rySd3sn/3ODi2hPLNs6Id4qk6S4lTlvv2Fisf99Uh9gPIYVL9LymUWIP
6K8NZnrOfdba+6j+5cNDRCqTs9uw6V6Ac+iGLhSUhHSBtwZor+g+I3oOBWwLQ/CFFLDSRL1Q2p8K
JrrZMgTurrmA8v7zaSmJEvZp47rz8fiK5S8EKs2E4JxAxIbh/VaqhT2so0gk8T076M2BrFq6nps8
Uv5t69/3ol8abN0q9192T4L2RH5kQSUcX6SYIAWQGj+qGMTC6RIyqWszCJ9B4MjlBkM4qc5ScBrp
coRsrTvDa7cyDwP8AgcdoXBnHjf79w0tWaef4vCKtdkesHjj8ohURP7IZeXc7qaVm5ZVnx0NfD77
cBGiqvk6e8faNi/gcS+kzGzyFx1HlYBjV9GO7SfFvmb9TgbMm3vjmSPyA/bbNS7dAECaJA6QZ4Cx
Cf3nSZjpLWsy7jLD4J0+aRZRrtU9zv0chB0qrlKViTY5O1ZvbtiQywkM+Wcr65VTHdQVGcZGCRH4
MAdpI/fFUNWDciIleiHRZ3NOY9rNvwn/iwQU4yVl2rJIzjgCmot24EDMzEFmUy47cIjrL/TXqRHj
rn4VHEGfVBxPKZb0KaiKb0Kqy5pVq568VEnvapxl5me0gySnTRUBJF3Kt4GI8YF3cqZSFT21orRD
i3rFtN1pTiHWNCdLXN3cf/fZ79NFf8x6lPrq8oBjmd9b99J4XqskW7mJ7xnwahffud9R2nTV6PKT
kxPUWd/+ARGJS2nbEjhDJZz7AqDnOREpgcB58IKfHDeYHyunnfnFXx79xq5AymSVvdmbiyqXeE2F
13bpukX8B0W7O/43d2p5adyY5mNIeCpmnbIw1prRnJZnFT3/bND7DruA2w4OerGeNgCLGRnhXWUf
XrEaqn/YHZx/yBHUoD1f+XXv9yOfVAJoB8nj7mgiBWQH5nsIyu5eEpRTqseJE1KBP13OQfkMxM5l
sXR1SLeXS2FXJZk+iNHkOqILe135kD+PX2lIyeGa3UH/gHccB+RwzYReqT/H2/4yRaUiH/cVeopy
GXL/1loEFK7z/5xLJ5fUmuZLpxgd8JV1IkOA50P1Qwf0ibWlClRmyxH5KckumOFIBELnoJDC9toZ
DxTIP1KEwWiZIg2JF9zLKqNNSOur9ZrQuVvKhotfKkRpLJdY64S9H94qcs25hou4yF9s8hu0dhky
SMGFF5EsZSyLk59kkY7DML0kNsosTOJSrAk1y5xriQO14ClOaIwzvHX81nMF/00X11VSY9shHf6g
E+qtSRNCevhzsvtgjsnd0R2Kr35uBLdigM267aMPQeculhbWxxntxWBGb5B/0gN5V9Ad8s6tidbH
YIna5awyLmkFSinM5+mGN1r0auCt+2sfNxZ94ct/6HFwMJnkO6u7CNrT6xewFYuDZknDy3j4P5nH
78Z/YXO1HAdROnBbq4f+uZ9o+4fJOFXyXRfp2fgtSciMdKJ1w9K+5YAlKzgqRV5AgT8Vvpcz0zcs
QgCQIMvClGgYvErxTFo3TkEWSZPo6y2iPCz6qIKRJJWsRb9ViZAd1cEBjsOvZIhQW2lni2Yoz6b9
wCzJNN33bc/EFPmQdzNflLkPeWsLP+ROGb/lvIsqNwI9kgwgBAHqNjydNZerM9MIlarxdOl1bXai
jN8FnRxW4qHxqpCh684ZoCHsPucbEHAp0Kvrnsb7a8ITlh+tGSXOzLaPr82e/3Qnd/jMzS74NYFa
YfG+aMR80SiFTNShOz//7Bzd2lWXKVWiUgKhBTMOzIOkZ5K9UWFHGfMRW+FPZV2mgCIH+IUpR7Mi
1hhcCr8i3VUV/kImBWtlgOo9uY/NHOof+jd+M229LFIOpFENDqWHQ77jffeVKpFf/2iy5ZK/fKlw
0YknPW+JmvfFx/XftXxG2oz5jSBSSh/+p/YYP6GhBY0NzFqVN2NJ+CYYndUiher9hToFCTdc/jjK
Go6IWdx6KXrnBC+RUBCEHsgVxtDPHE6wJr9gjVgQX5scjNr2ctwSdxK2fTHbe3oW4wmC+/Aoeoad
MIPPWGYKajguB93cB9uupFruflIsTjZ2XK+2f2mziAR46c9IMel7dfG7A4TXO4Rz4YkhZKbZ9kby
55th0iTSOJ0EexpucjKFcFO7VxOmYGscUXXNv3NQJ1TuZxvoTukTyDsPEj+5dBgNbVT/ftHihYj8
nHEiYmoIDTmfijj5BGXv+4Dt9YKCxtiGXePTyYu8zeIrudD91wyv79YtRTI7bylTgSWlrt0Nr8Pz
2kaIXE/UU48jhzYue9m+LRlmW57CF2DbeiN4eIlU6HaXnD6/gtFvRo8ByX9v16wGXKBIuWcU8N0d
ngXiuST9R3iCo5GTMf+WZajQL1XutD2J1JYe590O8Oam0LIvYrNcev44k/Y0BTXFlI/etZCqQ8RD
zxDQ+PZBdZowSJXS+c6sUocLc/XpnIM0Vt3nH6ZvFKXA5T/Ww9LtmhNqOvlPkM53St49iV0fi+gp
KVK4QQ8NU+n1h7WCUmFjGPhL2XiTJ8st1tlrkouOR13rtXoHFF74e3k0g6qGIsMqxg6RsV0Ub2gC
0JUbySNJ4chvQckAIVnwLh7NHI3X1GgMXAfr9D1rBF3gXXOvw6DiI1BMDL3Lv2pNtg5AJPuqSAgv
p/L2cvIuVCBroAi60TQZkbyaopbRpwNjz2GzK4Gf/B2ByQ9d1gs6p7Ouou11w+1x5j8vaT8cZOXx
zEScz+twZK3uOWqQ1hvVFexkjxXeivftQoofd8ajqgH1NN0IiATelalCEyZSoT7neqUdVBvnwMhO
klAvrk+FqqasGnmZeVqn3v1VgLUTc+4dWHto8oMGx+e9IokbvZvLOBUS+OjC65MXqvn821DJ6X+1
D/wnxIXCPbZ7tVTEgga68/R6KxUKndleBRtPumtmr53Kwz3/doI91TztLCJ4JVY4McwN/mmP+awS
VuYPE3m5/SoulbAsARSUPdB2/KWEzMheQo7383iK4BUpNb2f5FOTnhW265eUOKGEkZGIGclDHx20
grgTBe6LeOxED7O33/sG2oVi01f2XRkRtBfb0emh3AdEfDz/o3UnUQGEygIUo4VxUHV7P6QByzl9
PAbBgNpzPZyU2qO6XBzCO75XsKOy1EJ8pauqXxGjSz0BxIm63T7ZnAxZWIypmgkXxcuH+YA+fWgF
dQS1YgqFK2BJx7IjooVni4UB9ofKGhpii8mHL5HP9FNAlgVDuERl6zYjA5f0uaK3/SEjRS5GZF0T
zKLMcPb52diNl+8s4P1/OOX4ecptoGQvEgxuRDC5eUqQIH/CBs8JXT74aimPtLJjrgi6k4qibtsd
pP21rxg9PsIgzXUQio8StEgLFXxutIhMBlBKZ9f8ZglJvxZ7jvuoMpgvTls9JUQkdYEO87Bym3qK
Xh2JzS7BZYsl75715hD/n+XDVu2l1fauLT3Tx3VA7jJV5GDkPI9Ji+z4EgOc1p+uUHB3xre6+Y0M
/wxuEw5HaGAm2dXnsF9FZ1EDYigoell3rjTx9Lr+tf+hAPiVHKn1t3lBFmjbPjlUgeLgXj5X93DC
dO32DT8kq3Rei6FsYCOUpuWUAkG7FgjidL0zhQniMYt0ki0MRtWyQqWUce6TUn+DX+97qcGYO6Di
OGI2kQEBsnklnGJviuDJ0ANzcqrJrng3x1hNsuJs4jgdFtPrPEyFKCUbS1EYn0NMLI/RZUw7ieRy
w148psEBC8DQTE2hnh5qCY84omaI5QnNkPLBG+nubPTkXdhm+WpAK/GK/p8VJODP5qNFfQxQ0FO9
EQ8evEmMd5Dx+0d91fpl0pN6XAYZpczHFfvwiSiZtRPipsI6Yk4Vk1cwhY+hENqX9MjPSQfSZXxt
WfEZhguOzdhqtM0OZEUen2a4XumYDOtzz558fVGuklHqupfuyYij2zx5jrYJSxMp4NzmQfQDjqZ9
mPukPiKrC0oNUzzJaPGb0pU0LIBtZaFuOL9Am84jFSaq+h5JuuiKXnNvtrnolijbFQoaXfQpdB0n
6AtH59gd29AbeGIeMBJ7PR5tsnexnGmwMR8T5gVVtgDMg11w3ns9AVzJIfqALW/4vLAhROXlv6aj
c/byRy4uVKJj9XMlsEkPBvwXybUzHb20y6tC0kJETMbXaDvgDrcCHaFQT3Wa/IcdefE/y21BJ49O
Z9ZX9yMf82Xtj3d4q7Vc9YrKFVBzimhBsSH6xYcEF13GT6IY+vlv0uGjgma6oPmvP6qH3O6Dvzy3
vClB0MP18inQByv/NEn45UkxMP2VtCXhiLgpTINFCy0Eran1PWWhOpt4WQdvl/o2PFqNYGQ286PU
87VfS7Kfxcxpga0c3SmB/3FiiBasRMFbaYk5kT/LzgoSedkp1+1lAV8K/oV7HKdw4EUue5sAq7sF
I6YhH4xa4ykW8KBzmFPr8igCZRYzkHD3xgpq2/AQ6nSXh63GWTFeDdyl/QI5F62xRT8AIa3JgKIo
Mrsay+HabJlgND81dKKl2x+PaHJ9mDdpWzB5K3d5Mg0FuxUSPoJBkMhbCiF5JAtT0pSQFiVsbsDY
7/Ky4Y/AX24KMLYQ5ztcwKopEkYk0u+ZK22/jCvHlto/R1RQsoXHyYKj06OpZnBw87mc0Vvvk2p2
kUadRy8VAKHs1EZ5txUrq266/cUY8oiecwJVy+ijlJWUgWKBOSzKBmQu6YxdjPs17sfWYkYXWMKc
YSDdx8i7vHIFfSogwW3DzjQVjKDBOKgw7X2M3Z49evVCg8+8IM6aPZDhIgqzi1OInjwXxy/aKI8t
JDqhP5JH9i6qpnvhVbLBDmO0+qqYd0bUgEDC5IZf0gjGMIWmUZU6VWKj6mZzOFCcxj/w/3QlUy82
lvS+rKqlKMUgZ8DzYBspC0TTGotWJtuqpDdqc1vMvzN1v7ORSMegqAKxb0l2NCdBYe/olvgL4R2t
fMc7TSE8S8YlqphqtT24kVc+Qo5esxH43O9pkpyeghEPwkFN7zsiHKgEF2+wceCcHtoZtfhOdVov
vxf10tmGeHaJyZY0hZ3eIUhzLOP11BuLmx8axVrOssge1cSiOr6OdeidUvQKqYmCrybU2ymMWfIL
cuu6LhINebLmpyernTv4C+LbbnhMYdKDPSz+PV1hmIu5PojWN59hA7UW57JwVC5ijo8QUhlAaycb
mZ+SlMCpyznQBj1x4QiyXKSharc4HiSigsRLUSvtODSQjixeTnvQpvmRmYTp641o6UsjtQpW1u8Y
406SHfungLSc4xwWu5jU/8h0ajaMW1C3Sl9vuNbh2+WIKzejnJuftmSkuibY7mVe51gvc/kFf+2g
tPxdPH3eBTTTi1lZilKZsgxTIg9Zxql68hJpRR+jTUkarra6JaQxMK07ytiOEQg3t0/G4q22xf0b
3KtTE6Cclj0+SxQPEohg9Paz1lmSbuweJopBxgO/jM8YlMerA8ZmHYPqB+rgHjMdtsHJUO/t3Jf9
lltSkKGTQ3xooHs6jsH5ZMCnCbCzom3WNPBEN7cuQvK+fkjcyqYjS80qhGnYFy10kL2/sDgDM0i3
mJnioq60l1Jwkq/Ihz36gJMDVlD/+NQOIH/IRNBTMXvku+XhHBep2jjhDH3+aQwN4Q6BQWSu8FdZ
9jbbhbGiTuhXyjIE5NvvNTATIR6gu2Qv1RbiXlQ4KoZ6piKsTnq4CiNq9kUfrDoyaZgJG51pF6H9
y4HGfslK3jqeyzOl7n43BsmVmwMJMTScjTq6XBn0wZfNAgI4SSJ1XYmQnLQ+lMh0q48AfHzxFuk6
hI8OYx2TILg6h460zudXNeR9VkCG5KPgvu9rxJ+17slLIJHfZ6HG848QzP84vlu7bnknKDxpC9w+
CRnI/GNrSUbktmX5PIndUzNDxv7u3tDgG4rsbNTof7Od2J2Rnsu3AQ5E0etIY+yL7ar1TpcL5Hfh
rCT1ODth/krSsBQ+3MWqhtjoM0Af2jyZfZWTNrJ3emPsPdSlbShygBnzkmOm3DdGfXnCGh01SWRP
ofB6+ZabHfUGzcVCb7gxwgQhEK0+RAdgE5V/rFMKXepuyRrIwj/jPQcofpGlh3LMO9wv/545mgVC
fR1tHIkzvx7nlOpwInIlP3V/SMQY6iYiCECqt5d3f5Yl+eL8kVYeZ9jjEBzq+xBW/LcwY2XpJIiU
nmYRzG45AjsrFXatf7TKxKfFqz5ocq/37anO0H+URWmWmam1JE/3QpZg9UAHmMyDsIoZL3HigtVf
kYFNoxaHxoqZpbRKzi06nTKOSOUmL5mors5RGXvoKbikpb4DbslLs+ioLONRukULBVSADxtiboDI
Up0XZfXhrzDssxeDvmNhqfuJKeZ4/zXgZpNYaYFjaylwAdVeuMzq2sxlspNot94rEkRykNJrluhh
jOgK5iILkp96A4nU4eMP3R9cAxG+hvSz5Gvl0sEXeGcjM6wCRuwMVK0MVgXxDrfIlJ70nwNsOsio
7J9sZPoRvgenXFFTN5gOtRUNeMx37z6k59hEfkKC0ewhqn+uhPRZm0z57lug3ZZ4JN7sI2lS3o5d
oYd9SQOL4RghkCP5CTbkxWa/JVAvuyqCPUALeWRn9QzGUwUYGmYAA2glLVW6eOOwZfDUKlSSaJAO
zVjZrK8JaVpiaAKElTCH1IFztlL7McxoWhdr7cKKJPjluH+jEYl+6816HbwJwebznzYkW3R5jXWX
nhnT+Eo4ZQHx2hRfiQ6fvRZzCB/s0w/EwvjLsVXcDQyXFmIfW0JaFZcu255c16xLUhVFhjciuq5O
lJxfV4v2BpCV0OIANhrs+DJMUFJwk7Dq+6VnDm2255Jmwv5zKRd52qWxuwb76VAh17R56pAEyvLr
kQBMFnqsy4kaO+mJdGELrRVp2ADoEn4R1I08HVrhbo9+hiEXykzwD4bqpLnQXb5zPHUhflyMe+5U
Oua9paKXwdL/VIbTkkeswFG9SyaFqX/BBBxSwc7a5KIOW/Azruy32UrQkl8UZaHynHhfbaCqYkVz
PcGfWwlNq9qk4nkWPHzfkZ4w1IUYXpf73sGK9OGtsM7MH1R54ExfrQozui4Ig0EaZWqbLW00yc08
WBz/+4iSh+hNtLazCG9t4y64H4RyMUZVKVJl4W8Ls2hRe0hzYyH7l9d5wErs104NSBF7LVrd2iah
xwmPIuVCsFEiLE1v9VL1nmZCLO+tfyMKt5g/9JOPthu+3t+QfOjOWex2arHllfu/8e5tcvmpGzq4
YnrRlVcAPBn+sE8tlOQfNc0+GSbZztcQMqdUqc6q75CiumUsdMFgK1eLpFUy3jCLxVI8pO7/hBC5
dEP/cbeVfXAkXhVLoc6vpltrJLB3gP877THrzhQlYSMoYrIbMKik9l4+GYQVpALPN0ZhZ9iJ5j/C
0gEWjeDIaUyMzqMqsuC+6/+mBAMEgR5JerpNSEFzXyGyhH+nDcLrgj7eYeXnbTaMhpVs/XadbA26
iEUWLZrI2fG/TWOybqOIatf8tKaK96XdBY2Gm/KdwUdr5snNjejtdTU/bTNiENqFFFeGHMIidFdX
HJZsLorhWgnFbXgcsLaZsMZbQV+a6pif6xKGspVAcfCxne/3BaJjjkyabcQJWhZ0oS+kZ4NCQNLC
//SqTxi4QrDI/iym7/m/k0olvsiCQljLhHkP9WUbmYoFo3SqcGApg6SzHAEYtLiO5Zi47iRUnU4m
msVaX3r6Jonk5fezhDfyKSiYZiDCT7FFaELArVpExD7OHoa/DdMOqDOKiqjQpjbaJNLWJVeEF7pw
ItzFMl3LJDA/g4njwlCrPiJrSkcfQrgWCAw64CJfW+n+wuRagpUfZ4wctW6v25ncud/wB7k66icY
36RWnLYOG9hEGvh8IaYf78zC8SKqgdf4AJTKyrwu97oBb653fzwxR5b9b0YpOx5JfIuV3cgS7FtF
SFsQ8uzzRVvXkzhkUlH/vQ7z4XlNKj6aek4zvdZLqI0MobFd2yIHujRpUFlcqYHmXLwNeTu4wGB3
bzgP+tRxLaHiWZzESsw/kT1KAXTYRBGYau3oxS+bAQ5EgOFb0EvqKT9dfTbXYOgyM8QTj8Fxz3X5
qe/bvy6ncfaV7rX+IuW3xvdFV5ke3zpeH71cbqN1RPL5aTPD5C6jOkSBYfj8rn0Bzu2wu+4jLww+
DUq9LB2AEPSTqDKRmI95yj+oEF4pLFwm9sRY5cX/EcfJul/06kbXnHpW0OI+1o7C9aH1t6Bt1Piq
B/CSq+4jobrv0B5hOi2W9aGqsDU5ruR306COCphgkn6Y2RHKTSxI9IYjwqHmnOdynda3BmgFt5io
xcMExlsLdkg2OnmzzjXV9yAn2kPQly5lG0duPmty0pTEWVf/hHKEX9j6PjYi8tnD/fiOo1g0EQ8k
rfDdsVZuQ/kzEykzRPTuObbKfAivBCvefsRUTp30Zf44yfFr2ZyylMPWbTwm7nAm3Bkyya0ntOJT
Teu1jZywYdUwvHseJGwqI/KPYyDO5uAdupY5S0GfVjVo/tIIVNaodcSZsrCov/fUNYqTP2ABHxDz
hYSprtUEU+aN/j0bW6i0BZHgsoGEGGq0REUM3Oa7iTg9Q2q78lAeC886c4P+s+RB6vqMVegKlWsj
etngPq1e2RxZHySa/7zoewUjn7n3nSBoKV20ss54AB8FdF0KwiLrb4m3JZr3h9wNE2egtzOK92vp
aLnFjTtxpISO8BrWNeD6E77iX/IyFI3EheXSR5Tzy+X4zd3wnJaZ4DaUQP8nj8ZEsZQ5eH1YIP5W
18plaOYALWJWowa/GLDhJLCOiYomKwftfPtS9O84/88z8OAZztz6NOrPnug+E+rl1y0x/S/t4bSZ
rAQcSSX0nLFpB6QAYPBZIsHK/an348ET4I2oYM6VC2uEnxgnu2fhOgJIcOajCE6EaroGr65eTjkY
N9vHmh7BdeJy7bA1eldTVJWb82CD98WthBj29rkA96jI10/N0pmQkjTM6cuUqezRS5O5Ydbp1iTx
DjbW3/Fb/nk9JrMAUIq4k+hS/oxYsSM/aRfbVeGjc/Cz6/on3fHHDmgIEN722N8IYDL0oNo+SlY9
lIu/rsWSKpR6KOZP8F55mn1nQDOClzyOst1OZ1YXLGDTkbdtPHAjPnpFXpBHh0GX79cYv/FR9SBJ
DDai0eYLhReDQuO7iMq0p8F2Vq/kNKYmiDWENLPByE0aAqVANB25BRpyjpHE5NYRCoNQXhHlbVa6
dhy+b0csnmJF9aaZ1HsJwBOspHlfvRLgQOG/eawMaKG6VwWOfcjX+iTFQl7WYkCZCYjIXCP+Ivfz
U3JRtHt29+Q3l6LFJPU+Kcl4tFOGLaU3heWxKHyIzpJGGOIgOkLgVfRyRd7oy5wnyuMzEtcnP4+J
qE3qyf7Qfl/AAKTOxsqpsN54u6xQtf/lQtvpDr2ZPZnPoU5nh16DXnlL+COZhJDoq73F/SgtDMsu
8IvIh984h4JgfJ3fz43RV8CLKVUkWIbGuWe/LgfawTYS5pDq9f8K8lfiChARqIb5atE4GV/mH7Il
MVE8ip3Nn5F+KFbViYd0DiSxWoKEJS9h467HWBbN0RJjQnR4IYSjftJPXQBNhv6v4f3ksx+OXha/
TOgbug7V0SF2RUYpnuRY13xFVe3umz7Q2hHxGXia/ZpB64zEd/RuRXgBXFT3bmVQqSRzS2suMKBH
ZkD7uQ/eHGgCufBt773uNPsYDcOMtM3p8/hfb3STzhMGn3g8mNmEWtB15k1BH9+NJj5Pa3x353B6
7tTSqtHUiWAXTVsMIlPqS35EueIwwE/Rbhf0LAdg/M6n4hF1SQtgQ1gnHyE/Rf3nhFqCWQACYKgj
HdAEv/NqALZ1gQwz//RlYpQwlqyQiQdco0oYeQwb/+kQ9uW51zxaaaBuS5cydqmjsaaIf5aEnvpX
SKovGJzrjBQaYEWYMaN8Inab6eSz9yrkFtQfIKFxVHHSKCYljcN+sP2pbc8wixTEG6YMGg/RLf+W
OM+45k5TihG1ghKiPNcAYc5kUAYv0no6/vmAy+C+2H4mEpDvG8V/pOy5phhKTTkTJt/ekDoG8PO8
LLtKgZ184RxNRCne68B32qXeB3OT87rIIfACpumrbO3ZKQYb5TbOSRfzx4Eapd4f4Tpg1p5BDMCe
YqQpURAkB6goYdpv0jj1GPwc+rpdi8W83sq3UUTwBPJMjthCAebE6n2Xt0lJJnXEbDG3AVzPmdwl
tQ7sPXmwjtIrhq43tEHxzLEEze1DbQZGtPw9iXdU6RSa29kNZRdOUtpJ80oAnGoEc6VxuRCkiUQe
GxffGmCUsKyHVHBlNrq1i60jPPVAmxmO3rNbr+zJhX0Hf4rBefhtq+cx5w6KzW98k/d64I+yCYM9
o3dxBR2QaEnfnOq7RlR++jg/CoVY6N2bMybWx9Kq8faLqhwgQSAmqmdoDDjYBklvoWeb6fr9DoeD
GM5NasmB90XovuXLYGihOECxCNqWStBrJz6ky7Z7pehTpSmob4x9/C94A9zRkOxuQYAo9eVyruwL
t+1jYntvGpNfqnwLItcou9dgdDhvJtWDN5XWSs0xaALFXoD2OEagQQFexcmGU+itbwInflYXDen/
8OKWinA0jN0DcMpUKJCJF9KGxbaq5ls99q+iPsN5HIBTnW7uLER5efMaGEmhuxwAs49Q7O37ymAW
9PfS845sT5Ae1biv90TLUi6hIJiS/qifZuuIDC8zwL9WoX0P4wTQ8PCxksL00MxNQD739rshWKx3
qtWxmg6JSM0qwNofnhWAMsGUfRdtqqIvW38hVDbJzpUbieXGNK/F2XPS8WhsG31rXYN5AcLkckn9
V5loXbUHwLnlTn+O4G3YmC06OFe4+00p7+PY3031bqReH1xFkY9XAXqVR1zwETw7HmGo5I6GuVdp
+3N6ag6qQequiFMOkqzakQzq7g1LmxnADzD+JPTljRs3vBOGifxBjMI1FalbyiRytbd1mtE4oi5C
AnGjijKqDN6KewuW0m+UYGsoyFMgaMWrTx4ElhdGr8/2BCD+eMU4SHidTLdQ0TgG5OLxV9A+9WgJ
PXCSGA01BiuKY0+ZM7Z7naHW0CKJ9/CeLwSl4SFqPoFXN9UVdqg7uRAXjXE6wA5Vip1QB+udZiTM
6I9BrmHi0iUylP9CDAFyHF+/TL/gWOR9r0jihC8UyqpU25UjMHQ3RSW0kum+n0luKiGqUWJ/y17c
aHg7Zkwzutz+++Oe9FyICV9YBX0/s8HGLyVxLO4Bo4eUo4+lXCxYQetF9iWXcF9HfzZQXCPsiLOt
pWNHUmcLVgeAU7Ac8GJ6SuZFRKQ52GR9/g2kM9k2GOzzqBI02xoSFWpM0CyPCAzsy3XvytM7xOXB
4f2EsrQCrUYdl6X+vu1ksxD1lppDx/B/D6vbSaOCirOY4XIKwHZeUJRgqGbHK3YlvVItD34PF9wY
3crLpYTT+xldWd319PQkTvCa232Jff4kaBGtO74nuTaYa+enNQjyaeYaTj0FjwECEu/oVQJvWyhl
PT92oV+l98pg+jCj5AVuEZmjHRmGbvU05sMiZroeWjn78uR/NVwcj++ReWxE2Td4jUuqce3RgMwe
ONynJ66ri2x0d2DGkwvpzc/4NVx0oo7hj+F9huhqzgDSGIdyGe4wgxE1cYe4OCda4XUfNgBNnV2t
z7h4X4xn4jRILrfXD1haaVNJTqS7CUlDaYzXQMoifKOg+pAUZg9iL40dh1MuBsGMl47e/fHGMtzC
P7fp15j6ujE//BVEFAccNQ2cKfYr4D5DJc1Gbq0C5Hi4yjLQErvDDDLirmKuhLU8rn8xsKuYd7kx
hVzD82GFJ84ulJ9pSKQ5kopM+DwIrHfar3jQhx0YMyzYphcRWB94omT/W5GWMNrGlciYqRd5AvGL
pXZdUaVdN3zSojxfo2pdQLtG3r3nqjUjq7mNqD9s4egP0y7bxQDzFpWBN3jeMWpq5ot/fg/SgA/H
jryPpCfSrhzeYe6kGexi2T4XmQVXN5ytTqqSORtSisq+PDrqzUDeM4qUgftbHeqr+wpyGxDW9zQM
1qbU8eeGBPWSS7ptb6AXPtUMQ9DRL4fOwS5Lf8CZ0Wb+ARw2b4s/Bot+0O8a1TUpRBLQiqsJRQgY
/svZ+rEfes3O0tl3np5uT748P93tlsxsi4I/2uUVl6bIIpxlJCiASG15HTNwouE1brtNYTwhrahx
fxmkhjp7GLhWAbEMqec3oPmo+sRegfWqmmikcjyriHJenekEZPEsCUHcGUuzxf5ko3zJ8/lKwpy/
cbnLEXGC7rpqnW1tV0PFY73fUNmqvDDuUjfAqB9KwEG5vtHeCQiaXoGt/eQ+UByG5SsLoi43MnoF
JXplzHPhsifm/P5QSftAamGlMci5lsEk3YlNIE/vR2Pc6aezk11hk8qDHzIc0Rj2drpPnuSdrPdW
CfpC+s0Xb/xJTAPefzJkpvfEHjPS4FeFkaXIIF+k48yLH3VauNvM6dn/kAP7LgssE4mrfLQLgjtH
cb0p2BD9WE/XJIcsxS25KV1cbSXPnTGLwjvsV6DC9Z68c7GoWFQ5CkgbQBBuCOTJr+mqk0nLSNSp
w7zqQ8CYXw85dlQAK5euHRc/8X70nyaybxwVXIH4nIR/xI51yvnFUNJGwvOgz3+flPgBe8ZnUnx7
fDIm2ljTcBDOuXWtj2Fx+3JxpQBLviIESHNn4d3c9y0T2TK4howjQX+kvbNFmNUyabsTYuSom5XI
FPhubmOgUA9H+OycNX3QxWLDyA2/BSbZhr6RqxexL62/YTwcw0C8x7+WPgEQCYxYP+cA3WAXLORC
M7MGysBo04Xt6vE9c89CeBiBmn6T+Onsg0pv3ExJdLdK4B1hNoAntlSrYcaQzhnkrknVw2sPuYNJ
0bg4Z2AF2xKcbIhcc4np8znz5Tu2lm8GDa3wBvskl8M/ZF1BLgu0Pa1m4LjoOOWvnKr/28LEQZ+A
PeYPzK22iwGnmNKDRK9qKQGwnu2k+lu4vUO9HPdnC6UlxyH/srC423N7g7/9edz/ohyXTdBYmWm9
mNn3q+Nr/d3AAN5upeU9KFObLf+KBm2HmwQ3omL36J5gXnhpDjwgbJxZLRZUcbFoYKLDFV7tF6U7
9D9XzbkumGSlaANuqZ2ph9Li/K4X5K7ntVsMMSCjrCgiT2/+9vJnL5lvgSTaIZLYiT0L2JFxpGBs
OXotPfpstjs0elp8UEgyLRbAL42zsFEhEn6z2FLJoWKn2kPyyqHPHIlsyYtKLkD0Izhub98lom7n
0BljS32Evzuy+reNeybyEzqpTSWxmMZYjbDOJGA3tz5KIuRYiLy9IDylLRbTWz9qsHRMgGn21Q89
4QkWOXQKlU7AAYwEmDGDnCe9LUKLu1rSH5ZxKVt9WSgAm6cO9f3SViXdaq1u8s0qxj6K/bZbXRwr
f2FMRUdslUPsQEcoYQ0cOd86N7J2p9nMd9pDDv73N74ThOtFHWjP26INtv9Yo1BX51R9lR/Y/muT
DoenD+jzKJKcCeoq4zL0xFrcF7Vw8cDNPSup2FqTVciZVmWJzC/FCVsMU/F5TOYADgW+ESzuceuv
L0AgZqDibGYg8omEmcSzKGASwgitHZPr1+OpwiNHyiUIwCjXlozlwjbgAFlHejNPTIBYk38mNAb/
GLs0VCWy+gcdavrCwO8E8UZP2pIP/NIgct6voIQlVSe9rC+CP2HQnrT7n5LBvAHBml62Numrxcvh
TcNiXlYf2ljgajjnzNK9uprp85kj6SWUtYpvhIUT78YjZTHvTGvKYzQdFl0YbIGCCyqvthRHRXLC
PSpOzaP9iqaQyT2UgyPqKd/VaA/WlesfgcCO8/L9xy3wteIQvcFV8eCv2PwRmck0ko7k8w9Lpo0R
BOiGTD5dbapLiihPCW66ZojIM89GIvbPIHfiEBpAAw0o5ZPmy+5NKkKmWSBo/Q2LmjZbfFI3i+3T
9i+wKCiPGiyBNdhjv0ILOjxB11vhXYg4mBiMl9Ol+bQzplsiq46NAeBLpg8LGTYLm23ubBpdP2OG
OwSwbBOWltPvBhqY6ElMWXXVHIbJZROi6NqAslLhSIROC5LGs4fY79NEJ/qYlN7TLUd0wbNsCvf+
oTGIdPJogBBZqLpEdD1Tpefhv0K/OXu3dVbyUbtTsHJUFLcwoz6nGxXCeiy7uqE/kSMtKcjEDqdD
zCXNwgkMOEzMqEct3a2z1uyw+V3VPZmFqiWu3SVT/a9zx4SD9eiNPT/OGWWnVHEYvT1+NNX30naY
1oyExrurMRNN20c7010+kbbsUZjhWw2Fstmla9xvN3KQBhmfphiJplr1k46xWG2SwBAse+g6WfL1
lv9Pzl9T5kf69h9M5Ym2QiiJmd2ttoLGectBmgSO7TzlwVWtoKTl05Ya++PXMnSeBvFB7XW5VSHE
RZ2JOMDOWTvJ6zBKlYTqV4yp4cmGUwhYPrLrXCF5iaTTObwD3Du2aKIz+KUZuzD2cZxF0jexUV/G
QLQIUaJuvzfzbgidHF01TqvbhXueHV+Sx/AAamxd/E7rMKEolkoqh/CxTYFkI09eSsgov0qT/BA0
x2lBei1ndZN4OSMgMpz3ImQI9+Zb34KS41EUC+f7J18S4MYK+Ko68mzpysiHttDqE0RlNUzVhG/A
3TOcB170M453qiiC9zKMEK6bkQfHtjN1oaf8NRPDpf4sFMj3Ldg0cIDHXF++FDMtHQsGGTjbdx0s
mI0gFk7UsB3Y6gSg/kVhYmq40UMPOZCgKVg2qxd+XRjsGRoGHONX6hhOVsL1Q3czdGpx+iqo8FuX
BNOlGsexJA5IC3B1dasv5yDfm6/oYVb0mUoUlmL0lkalq/glrHTj1FyLKsxfjYSuy7mDGjbkkCtB
FyST/tmVZWZe8JjubGCCPEThhK/ITS46KX5XKxRWXW0ORtDxcJaeO4vzX1df1R10ghaiAI1m7cZC
xkzpjSx210Pn2b/EG3V0HBLMOcu4cxnuVD6PNbFYce1ySUrsvtPx7Bm7Sp+DbDzdgKrGBe/LLIB4
s0Bwnb7MCMtcioPcw8PphXLqhGovxJrLO90EObfgA4tepaeZ//7uVkD3lN3mZxQq76uVhHZcYcKR
FKREQdPJ2vnVOUz2n1ozd9fE49uRy0rdUb1ymymEzsHAPy7AXRJWnENvZa50RqimTqYGDjjd7HmJ
Lc5yN9B2qZUn9raXJ3zBwMjqEQME9Omv8UdgfQ553AE9bxnEe1c/evb3yq1pjjEUhAh+GdlGyqz5
MasV+oI9Y7qP1cYXXwHpqadDZwLECR2dckKDimOQFHuTi+xTUERV0LiciCEz/yXi9Jn8oKCnJ2CR
dUEzUxBSOhvKgVilRGw/Vo0TMGJkeecDdfsWU2BOIXOz6ScMNNyuAQ7V9+Oe0Mt0nFZGiIlwu6pV
URspvENkpTMmLuCBvBOr8mEaNFQS92+OkMM5KKuN8kRvDx9MpIEGtER3Xxb9PYq2YfSAuzIp0RZV
Hx9v4kyms3Jhuf3J2fbI5G2hfCWzfO4BCKzIAmznrc7N1Gi64DuT+KAGLbHzcnIKVmTmCCwUFNPq
Wg2+LOqGN4D6W0y54QXPZFOB1y7mkfjs3t7xU9i+/gypww5X79rMbANDfjn+Uha5SsM0iDCSJFfc
U+7OSTRU8OnAoL9RsNHr8ajOenLPUDfCHrHdrBy3+ghgleGXfBcAoNf2CWZDoeuCozvLo0xoH0PM
DctYa3k4sKH4MInqak1I30XwuGmuxzT8uq2ZzdHErhVO8YZ2CbBmkYqBg/DLb/UQKrn4L2y45K4D
wRWcGYE6M2URUNohPgh+Ep9jSL2vUz4oXCKxKMEhL0fIYQCO34drUGxqA76iW8Qk9ovOQlhRFTd5
syn7wURc0uWaWOAqQFFMfRUGrcZBFxCeFf/EbpnOwE5MkWJcv9iR9g3/hRNKZhMRn1/rA5rlgpEg
6OhyRkQM3KAwgwMO2wkRt6efpzALfAbP7kd6cWd/jwwkU1pf3EiB8XT4Yf+C4nfgRjldu6BA85K3
vDmOzx+burLtIygr3ESDIDJt2kGqnJWoKTWSFY1eo9e4CSjC/Fz2cNo8rI41aBuetD6i3WkQxcu3
MF166M02iBxmVLYIR8wWYs+79MpclylX+YFbDKsja+DYETiQ+9HMdTwARRMdxx2V2mk1IlDqMSdS
xvr1CTwrBEW0fXoMCa1TtMY+uXobhrtft3Gkmv6YR7vmVvQJKi88gh0R6Y9PAwvQTwbb05E2cYsF
nfXBJX0nd3lzuTAw/Z6+X2LnrEJE7xvsAwj0Nrd/WCRhrqIJeEvYr+wNpBvSq7gR9QBPh2qV7eCH
fXT5PIH4488pbfSV1C0AnKJNxbyLLf9O9IjlxlNMjUlAngRbUzLBSkNxfx7F5Q+2ig9nZ9RajOhq
GARZEMgu+HJhN1F2/JIw/Vw2N3zlxOxaOho48N/g/nKSbcEqozNNJ3IgmyAh1qR6sqFdNpopZVfv
xPmoZY0OvJ+nzf10+GKw11PNpmPJEj/MaF7U2Ht1mRUw/7bv0Rllc2eRUtvrRJUmjqpwooYiikFb
1cLnzbWBh9ZmesJvgeR3HXGhXqHLgXJTEINToojo2z4uy3gfFel+1B1Sez5WtrR67catbH8px/oT
+5M+7ONJSjHlysnaR1UuyAFe7g0uhetWBlkQ7nEmmTcns1a+YXv3M7wSUBnHP38m4b4MxOt/xv0Z
3o8TqKFaoOuAWWmp7NiX9govemKpSynX09QC5M7Kp+pM5wX/zVdpaC0HkafeILlpSKdesOWJ4xIG
c+vgt5iDZ+wGKXGJ8us6VbbrerSgeMIcmlFIJ/7NobcFGBMdPTPrdknqOEb6eDauGzabSo/wpK1X
ueyE9oRc6EOioI2IxcTPGk8tCjBf6FnnSUotopRNDE3Du4LpPvSrtU8nvN0o6BNP+J27DNmrjU0V
EU2LKYDqqeUIrIeo4pn/cMN7gHpDQT7oSfV32rn3qhyeC700ljV4mxR04TszRcuTIAvLG3hkvZ+S
1AmYWpwOW3t8Xczc+CYhFs81aVQd7JPYPEgd7mFuXQ0zDv96hCV9QVnFDIx4Z8HW42m8uhdGzy7s
iJf96JD7HuSzllzOMWCWSNEtILNH+wuxoYCA3z54pyuIR6NXnV/iVbQMq/MMgNFos4ZDGu7mKgr3
KZLK6eZA6uR3m2mVZ5qFjp7bz0ADArKGr62OHv9MHKQXCrc4elOaPU0RnLmLpHMXw0nAcpWfynlI
10JfVoCve4l2XnjaCmtPBACJtf4pHsoWnf9DAolyRuNIeFpRvpreboVJBl756ARl1vIIyMhHfu98
EADISZabLxXRv+rd0tMmo7vK7bOD3CVgpFXuIbLtZH90s/ze8bOzGEAxiY1iarRkdKfTFzyVJbko
8MozkK2X7+gHqWqWvHcePr5hYwDd3AjDBUqG1dJR9a+uWsC+5UVDzmx/kGhK5rhEehTPT87aYOTS
TLtDMKf3sFtMMoxeW0E8JD2S4EKaWZV5JfCkTBo4Xl1bfAZVN69bjzQE6zyFqZ3SVG6Rv9waiF+4
2glmk3/cE0DETEwzdtrMW9cfsZR3XPsYdaMXVo6pmWYbj3f3eduhVF+WS0rpjenCy0z4wFmde6Lb
RSqVi4Yn64tcuELGWaV5Tu7yxuzT4bNav8m5Zm2gjQx3jpQzoGRUIz+F6h6NXhTCwl5H1KKtxzQD
eJZGV8/FBVS4rcYhdoF/VL+CKnUVoTpdoViXUwq+nC24ClGZsDIfh/GriI59lY9zhz8umO6jWnGp
CKTDVyAxiAzfW8DMTOfGjttlymQWhBToYrhTko4j+JbcUj7QFRxXFgbYgzxhopltAccdGnERaFCP
vIX/i50O4hDkseRh0H8kWTi2a1eHGRRL/JuBeZMhDzmvqWbzT28CgUwtXi29iJa/PJdRbALsFv54
bLOYjQn3ZR7hMQAK6msgo4JwqUSi9AmPz0d0o7FspKdbixa0n7g2HGB7sqWKv6HXeC7NhYwwp9D/
xcDp7gwT3QecBpny/Exrw3TXauZ5czRjKiLV8FJ32dRDoGAj1INn5srjq0w+sSgLKa3c9byHXlfn
ExBg+Yqx7kJ9kXvjfQqP9wmMuKqRhWUvd907oCanzWA9060tQqcgxeK5iaK3O62kd3Qliw/TJYHw
45BQoWZUNESemwRYXAFyJ/t5ZL1MSwxwgwlz6w5bWgpRVXdvnocs18id4i8BxxIwm2gCC7tw+e6F
eVdREN+xxQRfsWUP4kZ6ulcyllYiyK1hyitHim847wBbHL6Zzhoaul0GtIyX+2YD8zQvOl841/wI
+FWvW+8w8u0qSUkYp3Iypym76yefHJiPpwvp5+zAdvLQkEMhoY5ydAe6e1mR2c0MaNaMOKq8FCML
Z0h93Kiy37m2pgKLa2aCV0XMmJ0jiCLsflx3iUbowToUiAbIiF4Wwf0CinBbT0TNC9vyO3IIcJUy
YYPYY4bOhNRX/sre0/JP6PyMXLd3KLE41/no2MpcL4+7xbscOGCQI/rqIjYFBy075qcsos3jNDio
WPLk+Ptuf8x+Lm7Z8D3L0dM5o6/uzTukXe31TdeYWvRusdhrRNlJXsONK5aCKvxsgrhwvK1HM4/6
42mYUyd0Q73aOJ4lGEI8IqjFtSX0DwPDr8D7KWBr6BNLuxumE3NtEPhMLS/fQl00+hxqMM7aTeSN
WXMrqYoFJdOD3dDU2yO2TWj5B2IKMIRhG4KYsqSbZkKE75TBcmW4MO3ZdT6MZwmUZMCL7URmvr6r
Ainy3wnNlDLBjIhHzTXj7Zk8Bm1LuQ8BDM++WBlOgcn0jiby6bARxoCYqnoPteDnv6vM5BPWGfW1
I6tvsCmGgT3tubmUD1/MCtaEm9ha9Zm+nzHaRnDH+Mxy0tPWn1+N321YOokPRQyeTI44PZ+7Chwt
a4OPZOXwwFkAmblyAeTS7a1frjdpn9S+6UZ/RSUolvW+bM/Ud6qdiLkwcEHfnoYARDzEUa1DqKoX
j7P/SHU4JZ9K4RA3p7nZBcIufduDx68QF9UsgcEQYdhajUPQLtaABht455T+uOGKDcMqNbiOKg/C
lpykj6gstp/7yslihZBK854x8R+pF2tIlFs3lz8NQQ5nNeG0M2TPtghT82peQ5ZOpcyKROh1yosT
5NZoT6bDT/xjlY5mcFzHiWBCaoygoNvgI8cOEgj9MbWqRRd2JS193VlbgPL9BGDjUj1yA/68y2Gp
FKNUp48MzdU4JDBkwXJ9OHasqv4f5raGLJHmmHk0k4POgWlg1FtAfG3y15dy6h0IOdYro6ts+rbI
e71T41oiS87xWeXSMGOii8GNxUl0GYOtMurYAUEMpttnEa+VrJwfzyqdWXlehuokppA5tblFUKb1
85b2+m514nBG5urAHQV+VQDj3UmH8vnXcsMXZhc7PwCIIZVp5sWczg/GRK71QLKo+c2I8ZM7Z4/W
N8xD/ZHNEOAe25OCPYhGv/TEiZ4Dc9Bhxhj53ssKEO5eGDG0C+TyGn9dy0wtgUVx8nY+f1ICIVby
RsHmqWbIK/KW+Mi81LkA0JAxaIx2ZdwMmtJpYNgsZflp6Xjy5fy9FtRzRvHVUes1wOzuSoykLg4e
Co+x8Smg99So4Z4N3dcU73kky5f/iAg/AymeUvk2Lkt9G1CERBLV2PZ2lEHcsy+LTYGjy6te0k27
E0R0iV946oULXV+ImcqxHqYE8bIURqQTKdmSItDZnprqeERkN6bXADASCmqZ8ail5/GFJJ6Hvi65
XtnisiLMHrJvjqq8bWlcmCGKtxsXXoDJDIw1CMkBmruacDsttkVUmiwEI2/+CRXPirgrEv/0/YHJ
JmBdJN7QXixKGWMoIr8JFO6+vGor39nPGvR1SPuFW5+2bUfy5UZuOaiNJdNmgtbmmnfjRVpIy1pv
1KnFFrxG72wJJaiS9/yfXTpts/LroripZKKmMJ/QdhN4RDYWJ8CR8IWvpSkpWApX7prcKWHEg4Py
seshNg5dG7ZCpPbX1qoaD6tPVEoh4k8AwuXg3CiD53c9mjsX6YjIjdREV3tImt8xJd01tyQEADHO
Lo3jIyrfB8yAFAR1vftR/I0UeaqjXDEcY76CtGMXhKN/liFJyYO1c9UZtE3KDYmRJ6DYV1uf3ofx
bs6IQKjwN6NMWctjjepjGih2mjy8Ok68VBUfHywxSvoLBlOe/26362qgde/qCem6KLMcv/8hJX5m
DOH5KqV/9L6tgohArMiEbQcj3aIiKopq3ToIKYhC4QjV/LXzniIFUwvHnf6CRNLBqxhxzcoSUyJ2
jYGnBV7gTx+hdLPqzPLZkrfe1/bEEulFPoWNUsXjUxidpAcuebRrZ+wbXXlIksFoSHVdmyHbj7os
xfCA3SKGud3kMNdmDwDSRGHkEDJq3BHHyt4aSSfS2t6qmTZytj+7dxQpJsagBEGjdRXsAArUR5My
3GZ2BGWmN3lmZN79CF0LqI7Xpuqfj7RVe6Jbxrup0Pj2JtrrAz/NL3/50vPJm2jBlnUxBvSxNV+w
hm6K3KQdP6jskJGiuqZwiHhsuDEv4VB17+gyAvd9gmPUktDJFUycyT0/kqlFLgn3wxkaBFC94DNC
VB+eQnsQKWI0MpKUwDjp0gY6H9fhDoxPw4DEBP4h+NvuW88kU86ZsooWyQnAVTIP1UCMKlcP3Sfd
xG/jwPvuMmvrR2pkGipAQLNo8lhfzFtc9ujeq0bd60QlWOGB1WL37UGoh5fzbVTJF8rvUmdIvhx0
RXgvqYwp161gwzs9r6LgHvJBeDEef0Bmwn65AkR6mqaJuZT1zJmO0RdwgsgXN5tcehnL+OgvhlAc
2LEmOUBMvaPI3C0qcFLMneu2w2PKuX2/1OgrEWU7MKAJBj/fLh8Lbsh1dljz9o/n71u/zPtoqh2h
bUVlSLen6Y5EhdpkWvudqfZhXfInzemyTJc/CB/Hhx18BkE1jucZm+qjVYsLVqx/iVpJLqIlxhKu
NXUsII3EZmQAucSxq7uRqCJAdtxGqwe2ecoLNkfbLbJZLOZb1j03TJIA/BfvX6xMmNQRSdBdzfuJ
ui/O6gtJOdheW2G+5Iy4GdgXLPRbinymRaul4bd+8ZfBrKuo8l7O14fWFeJ9Q8/fA6oI+WJn0KeR
FPG+g9eNJy/PtzWJAnhav7hHlTe4L1oFNG8cHGt7ioY9ZOtpICJnL8DJWPKxfDZoyNG+LUaze+he
V1I4cUbdPrSx9m8NcP26KQWhc/oyuqw2DfZ9W/PjpoU7gvIIiOkZ/had9CQhuMvA7wcCtizIzeFM
nzkKtI7CEOvYlVTEzWWCFpEj2O+N/O+KefltiPhGF2glmVAO5jkwE3I9asdlKSOUHRUZX6WoyGhx
4g4/1FdwwKUI/KSTAP7E+ETqx8doPWzZ2HtIpyccI52gLHS5OpKYJW3rrNU/G/b2ZfLFk/m/2d91
UXUGkCFChnNZ98lvHP5+VAi6O1EQ4n0CyELxrIrPCtgZpe1qk+e8efKB4oYQ+ncrSnKpK7/hQVn5
fwOeCxmSiWV6O1pqSNdEcRbLMUpx0KSRmvq2Rl+QQVrXVOdAf832ZK2cOXnuKnyFAcmhpK+wkvS4
RudS9v+B43Cdbk4FhZfhKNGHYT7RiSqjkgxusium6/vwjsWST5PfCGDqC6+6D5tZKte7af6f8f57
XfSnZoKrJaMbIFHLgymVkDg9nk1gJ4EfIDC3Uzg8f6s49U3mfPz9eX8HQY0JqagH1vdCW7XV0k0M
UtY4IIxMcsLgJOyg98UH/P9iBJ1tTYPUXk2N+qW9HufLnUooEOgNcV0GJdNlP4wjSAba2YiPhx6a
8V4BcOtPc0d4hcfncORaX8Yp+Nur6RMwMQvGvTLS43y4oGGHAYrQWwfIsW8LONqma3mnRBOrEPoo
AKF/yfhpmvMHjD7UTi7XianKawCBbLnXm8TGRdqBMpsWOJq4wgLaIP+5IPS3UzBJ+E5jHt/DNOsz
MtRhn4Rn0SiE+lK/w/pfEezWptFQahN2icvyPI1EHqyHo2zP0fFrHMdYaZFejFFQ3h/+fgvBNmbx
vGSFVeBuAadpr0pkXMN1rgH9ivWBqOMDFZUXaYDtPrdfbc/1RQ/Ypm9blUT2uTdQr0DI2U+tO7qV
iQGBN/wp1faB7Qvy6WYuVFeOEkJ3eVs70lc9pGhO/wL0op0PJ6XP0W8iNnGhoe+DHbFJMm3V9Qtd
2MzjcfcBwPGV3unxx704yb+xbg4AiCXT5zGAL2xZhCpM15LJ26IYizzufq6VVGeil1BzpIDw6fJ2
S2z1OZCeObY18pZxgr3Y5me4ihaMu1lCLjJlEsasuLtsnVi+oEeF0t0k5fgSoUvoG8tjU6Z68+ai
Q4eov2BFN3bfhBl+GFt3TPj2vc/VSHQB3hewoHbQ59fT0PMT3FqHe0JhqRpnPZbQqAR8qvNdkU9I
2SSPWUbnHhuD28MqLOJwIGTlnPeDi4yPjCavVPr270heYdDMAjHyTfkl0FjEF36MCxOKfjjuukUF
dax6SE+luicv3UD+zyQvm7Wv+BSG6it+iVW0Q5LEv8oTslNoYc+dScypEKWHBD0qWK1MJ793EXTF
Dz5LOpcvh8XlGj8WhgNyIFFnevQoXlSeEimAmOVuUYc2T7Fika8V+9zzJt7aZpAe+KMSU5sdT5WA
4HWaYd6+me+9X6/gt4g38TG7QFuWJUxPhZWztp7IcjlXX5U73VNktbjObKaF8r8G1434fvOXp6qz
rk2YZcIDFIbAUvYhoQKXxRso4U2qVVChSTyuPfa3e5m0GokU7eY1XUGBHJSsF4TE3vcaZROi7H/a
PXQ8o5b7YtJu9rnmYjcgOCqCtVHv8jpgrFioRvmnMHcq3U3ficxkQoTuz7CztnchWW0Wo27N85Bs
nW8WzR9B6EEuSayZn5cfjiC9E8Pk0YmwJLM8h2GXj3KybQxo5Z8N9h6iGtO8d+iVM+nHRcB5pC6C
Dpj6PcCccZ6j8piaP7yvgPu/n4RbTn1jFWiXyinZplXVSS6htEOVabURB2x46XOOQuGU+qs1pdmu
MGuhDJQFcKu0cY/10wtoRZNSDVaw70i1HGtFNaajuL5axpUNCKbSrS/8+DViC851L72ZYKjw31lw
EfptmO84ae1p6+d6oUtT3jsZ1lbILIMtu0r4tDdpZeqeGc1Gp8lBHKhWB1cY2I99MWHg+hT3Y9Jb
2zbXvhb8Mp8oEFUs8ggBV017zbMasC7X7ej+rfR2DNdFA4Hi2s3w1LdTZLM/i46ELTtqPXDFFTSH
dhgDD+eFHOjtuiNSIZhSXHeVwEK/xMKy6xLyRAHLwYnuoKtxuWUv+BZYEhQcgt/uieGn+sL0R6Ls
NzyNr/7mmxz1IKVoMB9IvOiSRI1OWEtdjWfu9Xr6DMmVdi0kyJ+mRWiIEUZ6Qhua9O3oUKvdjmnt
fhIFMib8Kxc8c2GzvBiKHfS1vnCD/gQ3rgflIJQ97R59alu4SATD4ij61DHJ8kejMQSONB+4ySgp
P8dR8tCt7eRjp67dNvHu8yC3+jznZJyNwb6UJC6rebzj8wx7KY+2vplVwVGWFX4Vx0Rs7At0/H+E
snNlqFAdpezsYKnyPSxUqPcxlzX49BElAOr0Mn+4m9it4EiI3CxE7ZWY+qXf8oubzmVneK7cxJ+I
ByH74r88LQhRpT07goVf7rRIyAu6Veo5feAlHSq0zz+H3Y0AXIhczMLWweQImVMCcegv7Xs6fm1h
XR21nkofv3O9koZZI5NbbXTtT1k/Y1cyNZHlPLslaM3/+jr6reA+St5bF8TwQv6pW0OCvlKU1COq
X8I444/p8nbKq+B0VqFgzjp2NQSSQMjlBkKnKZrgLPusb6qhhQdDo/bjlN8mNPhmu4mk/17J2YK+
nZvFHwhKIvCSsnPdU6IY/Y3S9r65a1cLcagocxIQDBTluAyGNTun0MRMSrNGP/A8127hOgq8vL0u
C0AG805vw4IdCibzJy9y+7mOxYWO8ZSIqk6PcjpweQgj7QqaRCo5bkpodHMxj0qdxUFHf8LsUGgJ
1OC736eZic6U8VemfaxFL4Yy0JgUz6adLGMBCcEY8i5L498fI5HLT8qLknTvFLK9T974RBMua3xB
wDVbAPymE/0UlvNBxgEAm+sFj8os97NoPF2iT+k60h4KEfWUYC+gd8oG+VOQpXanOKignjV+C3HO
m14+s61OJ5AzyOvz/cIXahBjgFHBM/JJQzyNP3YZKqEpnemf3Ju5cpuvqrjiU+awOUevfuucmMaI
6JNn/VHJqkRIMpXchOE22fHllDP6W5dGWbcWTAoBIxSyGObOSKV+NmmZHj0C912kgCiw1gSc7SCw
UV48JksKFFFh2rXRTNga/esNV/MK+mD3ZeZFYFyHnmuydm/YEsFSgya8yRYBqFXdtq3IXkZLmo1Z
QENkFg8ZlAj986fGfLoE29OjI9ddrwuEU5C8fRfSj2pHYSNdB6j0x717Uc/TDO2HaqSFWPmyxC7L
NYNSIDYVVNsltrCXJBBb739PzgeUTN9Fp2RHaR5PX2R0CQBZVbxiUGNrt/rNokaqoySHk2f8Vqco
PkGMoNtBdhXPa6AfMcJ+V6fDnpbYHniDS63gWNzDad3btb2C/RBq/0hsOyoab3Ny8+iHLlfEI5AE
0SPpwXkf6OiBNloja7oI/cGhIfnw1Ngtv7VyqinMUYciVmBxyVhLHC+yigt8by35QnS16HWAsitK
Vj9wC5BMDzVnagbtIkamUmdqLmYWCPaHTanSlG8zZB9GlLIlQ83//VgeB4RoXxn8aqUcrVVGVsZR
7ocvPSuVGKtjAHl33PHb1T1hqKC4EuQmzD3FPJzkyCCFnuOZw5PsLKnzNRjIrGF4RfXTezGYOGFC
MPCG5KV5jvZwVBxMktSRTOeXfeFL8MF/mu/jjTybRRSEPZ5a+QTLOvG+D9POanbDyWHtbglPe/Pi
rebbQMi+KKkqCaDmWuwHwmMP4KVOCyhCs6E/tNaxkTrOYqA7mSlmjP2SznSRWDbKLvAcAxhk0b0X
00t/l8yht50xaxHrqVMCl5Q6kfeglMpuFdyvbpqv522d7ZGNHb3Ct7tq2xr0hEKV4t7icb/FFivj
gSPvlrR5Qw/wriiYnyQdZZPSqFecLEMxwV0Ok92VTX6gzLgjDrbezpWXpsSjeRRhKvwK6N0C784r
7GuFeJ/uFI7n2WquGmRWwdj5FyMTN41ugFQaZ/X0lrKzSl5gl+eX9RVfq2AtaEfoQMxw1gmho7Xp
v4ObQf5w3Lu+et83qsx0324Ap+ebJtD5sQ/8RD+hOkFgLr3ik8d+2WC8QlK/A/8ZsyafPe/GkrD7
QGk8H954ORg5FeU4FpYlhdrQ++65LG1qomNd119eY0yCMctXJJAYaqgBdloEfEk7lKCy1ebjX930
QTdHBHIEjYxhUu77tfHFQJDr/3EV8wiDFosGjlwY+A==
`protect end_protected

