

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
YdpNuWNv5ANxG6sesr+pii9y21Kx+NVDp0WoJ8gKKxKHNSppxy07GkwBsVP2aDgHIw9l2ULLZTNZ
WthaAb5amQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
kEIsWLqGmgOl8w9T2kPb2uPP5XenCQ9kpxljFoCEGisg/vUEuVE5EQlDS3+mxviS53p6zH5m8hA5
bszDfKwHD76EbEoDDpJWL09MvEqH4hbAV7G0A9Qe7ZciYDi8os/DYZvhR8zjbLils1MINgQgL32T
+DXtGPXNuzJTAMDKzws=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
NxGGOrhc83L0V7+Qmwb6+Gi21+qsbQ+hA/5/9jysqY4QYAqiXfCrWB3N0NrVsGWuuTvZXoFNcxot
Izvlkgh5KOucyz0ezFvnhsYziU+FkvqQYf1g82Syrsz8zvyVWXqii6aXcF/WSMwXtiDjm4MiGpFm
yTcu8CcJgBMXYGVZx6nj+IgO08YgHCC4sfTqmgIgkxkmBrOsiH76g2hPxvXPgVWaBlJF0bS/hLIS
Glmsy0cU+pqQlcfbTEV79W+sXQ5Q3KPQFXj7AhMrHHD9esRm2Isg/tuzcRVk1cq3LsMUN//vGrfM
OKoYOozZxl1/IflxrtIzbjclaBUaFr5bvZYMTQ==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
dIJ+Oh/ID0KokdCrmxnp1QfFJ5QZBtIG4FQx5Pan4DTwhUxDWY/BQobSBBDXzWh1TT07UPg0V7Ui
zobKMfHgBNkMD8/PoD0AIDWLDLeXLvIJje8mGtE07uncec5mJ2eGa/WSy5sFj4M/Vdtk7C/Ab9LC
9qAaWZZ72ZUoEHuysZg=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
VglxNkzPd+guDL8DGRWVtgWGTdJbzbKKn0hBXJRIK4IuLrtOeezNwjLTIb0FIMSJGqYYwUrPN3z3
TVnjDJDaG+HA47egpMvivRkbnfO2/EAJtU7n0hK18OztWFzW+yXOUsOuQnFS20EGjEAN6HCMCAXS
ralqFAJsvMtY2y3dJNuE6ytT3WYkXmZUpTrJPPJOu2l9mCOnHkBU0dRG7RNYXf1tEMPaZrHSYyvp
XKWW5CTowIM6jJQxDVSVfwprGmWFUVJFtAmp+65D3ADXiHMcwre5cI/ty7nYS3euq41mrkrZyEF4
iH4/gU0xN9mM3aF9hBPzu3xQrdML35ONnUZTzw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 13184)
`protect data_block
5Ff7XIc/914rleBPkyDxnAzT9Unca7rCG3c6gwovn19/ypbWqnfGdyBXKtnrl4OV01/MSFzg+agf
z9tYQusBHGZBEA2oxAeoymGYryKQMBMjHcR9Z5eivTEzb6ledU3W1b6djSXrv3zVDFn32L8iKtAW
PADjz4sfXDSIMawElcmtz5OqvULSO5PMoWlTmPYyON7UgtFannY3ZUfPFtXWF9cgLcvpJlnz3Iav
kj96fpQKO6fE7G/AI5j+quDYuUNPKoswY9kKULLwHd87ffWhnd5E6XAcbDUGpwaIEJjpx95dL9n2
h8XhffyVIW4yWGC5DJMLbbGfty5Egd73DnMMnXNT1bNnzY8ZiKdcG04uY78ulaxbXOs2VVoxvB2T
uuk9gUBkHs1rBofp2GO342ldrEYNeZ/cgQUFSOP9i0SQdqmzfWW+xHBHuumg8nHwTcLAywQ24naz
jvADvmr9YzW6wWz5HTOYa+fiQnPAuSk4KhhjxMljbAZxjUXBeZs/39maRVuR6ifuN4HMAXR/5NcT
fxzrOCwXeoWP5Yff3QqrDs5xXh51BjOnlew2ivyN6Cr6nEvfHOXdz9JlNeqC29V3+BnSmr04qmV2
93qIW2BGMQmTNa0dHCg2r/j594fwD8n1Cw91+5NT36hs9ViYvpuRAYLjo1Bc33DG01j1DvNVgyXN
SKPQhRhycWBvfYV9Q7768EK5DgzPkdEeMh0/8Ph5JKcfJpkwgtpiG+wOg7VUVrUB5HhPUt0kcL3U
xd/OPcTKCwFSATQ8Dab32P1GmhwNsCxahVUlVm7fL2XwPykqVhu1oifFv92L7kkFuZmXJ46quQM7
Bpidd22aP2ZQ5ZKYLtjPiT3HDqWpevjX0HPrEg17JEATbVetwvdW1fWIX5gqO6CotJ9D4TgOq0fR
n197LT1CdkcRHiRAHUW3YBSMbwmguQ5eWEPhl7t60NSp0sUPTko/GkUvw9+NjtYSQ31GkFr6DuxZ
VjahilhjvoPIa8Nc84a099lRUalHi9TH2x78nC7bLs0d+yEHKHtnnnOXWoREcwh4SQeVVATYzLny
X++8cedZdil/JGiQrVWOe6UR6JN4cHK/GV1YEfAASMRU3BH4w+NehN2Yepb3WyzDfERpVpDDEi+I
p/oUOPq3TVtfMq8jEJ2c43vH14p4edqQr6Cc1HCk+0Z5A4z6vrOuYXGOrfo9JZGixLqpfeCD63v2
6sz83Nueg3XlbDEYchUUXwYlTJzOsj3r807azlwyhUQt8ypdpQ1xlNFdkzndCNCgJLoF2oq2Siq/
zK6FTnpYuHqJKpZi6LCZBHqfIZEp7y6fZclq0U1pPzPPtGzrmWG4v6mdCMp1UxX9/zLWdxTh509T
APgnl9uH3hhAq/jcSY2a2sPDk+FTbV1arR05fdwwK6El2RQ6Mn3kR6ROkSUsZHfF4aUpv5L8g4Zj
iGWg0wnW+JJLGPYXzQpT4yUzkRw5WfUE3UTMZQ2N5zH0J7HS0RvCngm8aGQW7a7HTxfy+gNhPFHS
RmNKPc1oBAz7DoP5+EeOoNom3T/hSJZU7gOc8a4Oc6Z264QKl3hfC2NQ3RSyUdZkIYEujnBv1udt
tUZ9gpNVMt4a014OIIeQ5Cxf+7+Qj5uXEUhBK9dUCBfzoMEGzyJEeqbPf2yAr/YrgGm0/tl62Zjx
6RHvAPb7v3irSn5fqkCr5l6Dm3aBJkqv1PhDs13bp30ravWKwLSI4U+oteabDmSrJFfr726vkohc
IprjE3T2JmJ6TKLskzjraZ9vbK+W4hRir9AJ5PoyPy+tmNug4env6kUByOm19J8TsS9+QtocsJis
Fdc5EXvR2A0InH02PUDHDieEbJuhn8PNSeyUiXOs6fa4u5gRQjIjZLdfn7dNuvjZYd6kCEFviiNx
CtETufSSdGp1Gf8ZZfOesaBGDLyeJqKso8buZjytGlbv1/nCfiaK/3mccU8CnSqA6ikSaoKnhcQ0
LHPRZ6QrZn4J0NuMa8EyOcYK31p99kjKq3v40rnWqp7urpxRW6ly1bywx2CveJIjm0618INjkUwx
hmKngAey7ld5RhQ/+erme2G8p8XR71hbnlUbCZU5zF97WMPPDgcOtsSUjJmYhAXB0Ppf+edXX3et
pu47ygz9Yo1/RmC1opTpR1CDeGz45LgpupJCp8ZyPe+ydNSNxjWl3wrFjkLdizQ2+kIyCSa1xCyW
+30mD6ellYFuXPqaeJyRDEG8RPEi1Jr9TJBrs5CUAEdTO+7Kq/dNMCW0B8pmoxyTtcDMiWbsEHZa
CyjlfCzKKtF4YKAgRS5dumtClu5RnDsYnBgHsGYKYkJdPvb2/xIwLOq4YzvUK5a1J8As7uPCjpVi
xF/DAmQpjpX7zfHAlhL6LKUYJ/Bqreji/uSh91ebQ9ffDDiBrJt36fDZojToRA2huMRJ3aGX3ju/
KW+5QuicSwnNIkgDR/jxx68f9H9xyDrRXu3RppjggSSFrIwW977I7qyBe6R4/JF7dUO83y17qADJ
QSdjBp5D2NJBEvXCy0XcJn4AjDP8Dms3t1MF8Th+901fWq0wMQnYl+4/UKqD4aMSV2YadLXbmqTf
+A7sCrArQwBN5vN0hVJ5IbMPJH5rPeAEYtUvaiP6PbAkKHsQM+WMxkAM7gzEqUNZUuLjHIe/9sv9
Fl0GCzNgizA4whLoxLv5ajRq86NTJB0J2kTNA8LEnrF5yad4I776jj01VJ45dxRuIH6DxTHGc6KF
uCPkjyJm4W/nzjKxluNOj2MYK8kBahZLowE/NVRL/ourynM6XnERPJwwwk/udXawXQLaOBkY5LlS
T02lc/+A5QVGwlVtn2b2tL/a4Sr4mvek3TAg8rz94MZvlsbm6M2JVokUHSP0wEixn0dxVCsUVUET
qZkDNN/hlOei8zJdT5V0lhqYlB4i9z0d+IRzTMtsPdvLrJT5OuwQWi7pQoOGGU21y5qo72kkiYnI
lKdfNvsyoGB1VAuX6iZueEkCwMyZBFlAW5YIInQ5yZWr/r5LT/Oh212oziZ/CW0ZRDRWejyZl0ZM
waZRntZNykjJ+7ibXlJ4+21pjH4X83zS9CcNvR2+iIiZxCyt0eVm2OuhGzw4HDZXX3iRXM1hrWMA
7k3FJ8kJgdMGJsRCzJZ1O+IMWkkq+qt1g5C9VRdKlIBTz8mRrONDndv/PIts/AcZBP85jqEennqb
UK3KjS5Ghq4NHQvLNwMjrcuz8ahF+VftSpGc9tL2cWttEMRduhhIFkLr0zS8PgXyS9z7L6DE6vmm
eaztkujmvCOZPOvKRnIK4OQw/jSFddycfwfdALuHnl8jqI7NOKXSSrYjH1lGFKcWrr4c8qfE03ct
hVhgLD69KFqoVLxb0GXlN/dnkZfY3P7901FStxaPS6Kjo7z2xbGSZPvXIe9JS/cXcFGDjqy3+Aco
MpAdQct5Kz4aavlyfoOrJu5Ks3QAC0ONTBuz0wB2Yw6K2TsUIiWsq2pLRG188kKpTqb2EtR1A6PF
lyA2KHyjwE1IE8vxYa2xXViryp0hR9fla8fspuakaiku6ksKPzM5n71qROG3CXFo4prE6GZZl71d
dL+H5bBKjYVlYhbW/MPJmyqJvwTImcX91N+agWUIsuTLGru8hC7UNH5rNn+0+9gcHadRcG7iknj1
9MJALZOjiN60SFHBVGM0+ZzO0n1SInCrU+Cjl5UalXY7F/0Vl01PcynC+MFk+DfNU9uNc09iTxSL
IuRfIVsSiCi2dlJulZNsYgVlUSi10MDILFbLybnSNOBdwYLxe+hylNgO82ZgBDedx/pVDght1TFU
u/KhCLiE7BkMjP5TohgjVo+P+tP18Nu5cnc1HHt1x+aOTApsMhnsE7fnwCEUgHqGsf89CDF7rgOU
7IJmSxdT4OEvbWrqgasn5ORRb6Ydy34IjZdxlBA6FSdhp9zTfJSCoMPwlDmNwFk+OAbOhCa6x8Xf
gGgTH00BimW1FnFpNHFks9YrWte2xEvfDZNlIhZNYo6dyyVGGYYqhfvalW74GdSu3v2b+8+8ES3H
M9msnc97kYaMutqtXsn1p1ZFMxCqa8yxVdFshnl8icnsmDArXhV1/VGkeNujkq0zyeAMudH3ufO+
Isee9Sjc2G52gZlmtLM70L7UAFsC+5IJ5NItNSVfEghxAw4hT+SWvgUL/DvGLgJztLk09mrw7wng
Nl0iV/FaNOHjaSIoGoxzkgopP4y7H2bj8xnamc7dC1cVP6lQyPiroD9daNZJY7W5N9T+k+PIkA0F
5GVJXxzAvsP7iAlG2tUmlN+jTSeb0av8QGjs1SGuRFJzioMD5qyUyVJgiMLuIJ1OHE5t9duCthIJ
J9cXCbajNCH0qxM0/nnvAjkLSXPPkAr/gW8amgRWPLK3fYGwi3nLquMzmlnvzoT6i9tg4sFr/KRD
i6Vw3sGXu1ChbMaboD9A6QOZsVDVaI73RTZCfJupgs00K0p/dQDwu0bba0uRMVVztLkvTfhROgQo
HCV36vjdGVGFvY9Rtoy9nRPhkj8PEQBIlIo8NoyNjynOyOELKc1H1KFYKZbZ7YVh6RfcLTWw/8UI
gDDaxP5mo7i46jSTB6pdUoHXRYq7cIfAOqCeysvVzwWck65SHPrflzd2lLLFvyRB0iltd4XFtH+p
apJMvIMxogKi9MVqmLas6veG3l6wLdkwvZcFwOrOrLNnDFxPGoOP3HKdtJlQoWqJSh9cBXv7c/ai
EQ0vn6S4CkN8y71DnyuS0ekeGpyDVOY6jKISLAU82hcpwgIHgYAlsxWuZSHa7fWs2dVYgIHTgoz0
PzH+5tZ8JFAAq8jxcDc+HS+MFc1KLmV5kJJYv+SYz9pBwI1oJhB82tr2L6fxpVxB27d1wHOtMXhI
nrujq4hv6cMJc9sMHeE6Hcjqm7jZNtA1NO6dCwlxXxfbVpAJ8S/CGV7qU6ZAKDJuJZNO8HeXO42z
wVrO6z5/ApcXlpa3/Has9smiuxGMq02cJblH0WNvuMvsDhEcwDEnfi5H5FP4O+BVgVu7Ne2T1FqH
6zRg/bSGLmBJzxSYJ6AgZ/eOx8x86WdLnA45DMeruDiaw0o+exoz6JQ6Ds8CirmXHBOtpAAWb0qt
nr1zCwiywQmpe452F44ordxUiIyTpm1/nUupU8y1ChzFTMtFbXJoyUcwmCiNLvu+mcVDTkixuVXl
GKGubApL9xUAi+qpoY4Cyh7xsBsKc16KtrfSHnWccajRIWKWDsKL1fpP2U6rYnK5QVZ9YwWAehmQ
uaYqiaZSYpWNMyViNPsmoHqu3m+53rit8ttf/2133kC1HdmJTVlvnvnaiPtL+HlP8tUHgdTUkLM6
aEXVmlu7c8wJgmNH2zh2J3lP1Q/rNAJIWV1qxTzJS8vPC+kk4nc5idwuBOYtkehn2yI+dpqzwG3I
zVR6b/2Yw+cckrOr9oPanGLzy77PwyDvL/M1J/XkdsM5TSD9SaFg6+JTpS6AmsfT6L1Edy+ej15f
ZHindI+5usDxKwroFdUIS8w5B/cq8Y5mws7/mHVCA2iTIR+I3xLcgwzbHUR4A1N5vXLhG/dNggfH
Qh23xOaJEyZJt//oMAsbUv4+e3vT2i6M0fmlBCvUbLe2+8ceBUuCCCQK6oAFhYK6PDH99GxZoIjU
9JSTQsg3rbUJwFlE8RMhm+VnMfV18x1bfoH0XmTZ1KyYeTv1YaGZdIqV7yGUlziytKpOdwap9rBT
Zp8Q7DgurNgzKCnO5tU4lpPczQVnClDXyEr9mFB0xH83A/wm8rMD3cAjwTNA3RkjehPhAke9q49s
5aezYAu+VAX+QFeOwKJFuSXLzAVYGF7/9H7YDapPnVX8fb6cGxiEMjpRElqc4iUoybrEIhHXLyz6
c034POhOdJj3gwVynw/M0VJ00fN3E3CFCHyYQCTyWHmqfjb8l2C1t00TnVZw+g3eDsFB5lmTYELe
VLzpO/YknIcaH4YorWEmX2GioDzK6AaGtFnbW0Cq/G6IJtwEsqp60r7h+8PYacC8vGIGuezz4Jmn
rEakcP/T6XCqqom6WatYwUS98m6M3t9j+QT/+69w2tCbQrspJphGZGIY4UeZjwMFJSVv3WqjNglG
BdLLrJnRIX9jQm+QTradVZwJb68gXYm+ZldREvHbHIWLjye5TZsJyqBPAzNBMiimoH5vSfkUQalu
XR6d+3v1QEeI3XN8X3QbC+uGGI5AuwR2I4p9ls6u5JrPa0pfQWu3C8YpHj2aSPz1bMOz1KNCJ3ZW
hhHpk2r9VVhAaZJaKVwLmFdaV+yDZfnEumCGZP1XuhqgvuugB2Dr+qa7GNU2L5Ccw+LqPRWV0e94
QmuuiDDFxieB55Csz13e/9Jfl+y77Eto+Cafy8E84wNCS4SuwVEGckATnHZ9MIjqd6qnRyGmMctn
EC6uXLjPy0EzKVGPcB2196Jd68mbqZN9G2WQ9NKgoeUvD+Hc3E2R8mXz+5Fnh00jwAe/xb+bcpWS
H3/+7s2k6oVwrAi99nRJPuhCn0tuD2mFKNxOd4z6Nv8OalLzc9bxxRmaYxAV4aOu68j8w8nHH7am
r4OrSVJ9CoMrRuK0p3ghpZ7RvgOZjSrkYseywbQdpbMIyXri3mXKp2rCzW55SlNF19bGOZejaTSc
a6Nv+0MLeW8WyuwJrrbD5+lZ7gJlJI2P9OVZY0yml0N6z1VjQ8rLiA6U0pQvK9N5cV0AlJKoQDfK
aNbl9Vuxt5bJszsKrUFlUqhVsg5O6uu4FwnJ08O5IYNg5Mq9Iazv7fVxerWDj5y/YJHYhUf2h38V
68V5rXBPwXW5Den/jt9ZJ+FdZD0bNDcynMr8mcGTAkVwQPCkDmdnmQlFBUZwFMtmjbwtIDt4mWkS
3R6AdoIy1nlPXx4KXjwoRh5pOTd7iC1Uelzj11nFF7EDmrxEkGJsckNeO5g2e15Yd+vbWE9lMT3W
3LAaO6+iFZwGYTvKEVHpwH2+sFoLfYxDSmAAZYspDblmNec3k2M5rbSRmXNwEiGnh/TZ2PZkF7GI
Ttb4f8JWN3XdmneCTlJBoev7j2gzHurcIrP5lM2jhZEsJBHn1ACbx4jtmn2NjtYRfA5McA54rzP1
A0b/C9nwDi6B8OpBt68H/KaajKBiNuNu2ZNyh9VGqVoq3+MtbeGIWA/PoU8na++eaS50S9PB9j0x
rd1yzjRirLKRbq82uBGhkCn0sKPCJxaf67iAU2xRKgeGP9OQgzSh75j6ga72+rrHundeU/+pwadD
F2rNVRU6GvdXfO93HeA5JGMKr9Ts4Ve4Melw1hxmlFDYpq+zQ/v7wMhUQOY7mKj8/cOCfhsnbxfU
O6ufOkDt0WDPNkBh+DheT17OwzpsJYB9bpWVu4p+54+/n0SDJ5scG7GBcYSqn1FEVx5KP+QAlx1P
9UaLm1iEl8d5JKa2f51bS44zbpOVaxKcZumCGv74N/6YuEK+ACs9jCy016yEfp+TB71Kp6AlYloi
xOzLPoW05CAjHJxcOZrnzyoITPUKonvJ0sDC8mJKyRdFeXPC7GdJ7fIvF6ZI4zJgEoimgVVQ/qRE
TJ4Oufgdh5fdXKa2NU4GX2XdrxJEvgcK543Ns4ZglfDM5u+Vx2x+BgBAbODr5e3+Ga/ErjPAQLKL
UjXLeFUlw0f/ulSX6lvLUtDMZ+3KdAoc1uBBcFTk5kwWGjaam+EAIsTbXJY766UPcS+WYgiE5M7Y
uGEGRf+e1s6Jxg9kZRKLXY1oceac4CZJyIZIEfoCz5re+wK6fGV0fOCxXv38xX85qF/eqtcOjk7W
1g/z5VW62LqKg5mk3gs2RALEzkoetpC6+e8W6YdfUxHACvk3HQ3x6U59ktXExUTTwpW0f0Vvg8C8
BYJWZxk1itk4guXqdbRGhLq2m2TwIdTcWkejSNQw7fXkrHb1w/yh32brBKFjpfvf3N72y3DkMHap
6+Km+K0TjI70pEM3zyujaCWyvIhl3UGZmabcotOuKcIqtVGFBNR63Axl0kEP2N3Hjx2m64hXg4KO
eKgmg6DmFqpvXTwCZBwKhagPdP5NYf+wcDSetuygf9Zk9u+V9xa0ceb/nC4mCgelriWQ1aDx5dyJ
mlc+YPBb1KmtlvItxnXmxXjJf33AblTpIyRvW6a9pKLsH2SsDwd6o5mo9WkYT6Zznpy97s7zNwEz
O669R7Ziz8SExUhY5CvdeSU7TWCq5uWr3Kdxg5KB4Gf1PHQIAkaxO1dsbAvn2TdabAwX0OMeYNo3
ZqoNoCWmDj05DQExAr6f3JiwbmoOcFkh8d2Sl6C9vSObh7IR0qjt9SIE2H1RFy2D4CLynfu5d/EX
vUP5VNBIHh6rPm1Jj7Sg0UDzSdj8fW5COgv3JFRr2/omUx1XT9ySeoHHcdYGTEvR0BYBSpyR9/X1
3axClgJKMd0+9RTR7sgiz4U9ESTvZGQWb6hbPyB6fxbeZreOIH+nNyMCDrt1tXeqnbPrK+fjkYBn
CgVJC8qUu5i9XLfdeUfjC1hRZUnQEP7vgXbGg/qkx91UyhSvelU/+/u4af9+cgjbcY0ajxubK5WI
ZZ/rB7cGWEpuvE2bL/s9MbvuQ450eAn0dKFUmOL1MuMsJenFcDl3u6muoZlE2Mx5n5uMl8ktnujX
zuJeldIz+gekQYqW6w/AJhcv7Xkxu8/L7aUR1IKJEKHhOJALYdkIsgUFo69szSTkH0j3c+LcO/5M
FxJBb4c2R7a3CWJcHMYkR6/rAn1asyVg/S29OEMBqjthhGVX1NjoJVqDyrOY27j4tlP3tZHHA5ma
YJDDxPZ12S33lS98mINahf5N2s+JpM6/eryE93/kGLaC5wk/ISrRPh43LSeGhj75JbMjfi+zyhLn
k3Y7goC1KCQUEjrT/fs2hCQMu6HgiO3RDoRvBRqXylm44ECeDKQieL7KFALXShKinmB6e4j/Czis
qgsUdFqgqKyGfdFfd8iHhFU6Km+OEBXq1BNd3BB2nBUjl1AKbYhdvF7MAYPwb4V1gYO1ibo5EPYa
UVKrKsK0RK6Pk2/ELivzIOluv+d9AZi3KxniPgNAoJg+3Ju+bSVWbB1TElTgggPw+NvrH2iUW5LL
YQHiA4SxSbDGGe65dGOD6S6i29lo8udJHlDfgKBIWt0RUL+2RcZVx/od6VA8PRHgga3cS6hY3brp
FMXrcGriNz5zxk1V+0EfLovobx4GZvHPp4k+uJNPVSW8LtJe/AwV+MB9+IaR1rl++LAm8ykifyLQ
7BJgmtaTbaIC1ajWSA4s6aBNPY+QaWBTtU4hvvAxJoQ8ca37/4h13RSHrxbDbJfhc6jzFIUEGorc
7W/KJWYi5wDS9cytJGuH47APqirvmkq5qODnIf7aRRL1FN+upbzCX0mLo1R1rN4VYwdVFZ8kyBkz
bbNERcL47SohduEP8UeXeD/+Z7HKgVKDnsfHuD/DNSgmesFZyU7mrIFP53QRxrbPShj3sU+b5CsD
UWpm+bqobZEfOm0EuY3KL+vDhHP2VR8ZEMnX6qiitIKqpewq0xFtuaFUPjubOy0Ftu6VOEd4cpsw
nxZ2EMBMi/7u9WcY/JJw2yZZxjq2Wk1lNG9lwDnh5v39hqha2Dj6NWI3h1xNfL8IQf1JORt7Vx3P
sQ6m/AA0p1dhMoKSp8Tv/9VIGmzqn/giTcIU2KRroYT9AJ/YoxXsh8uoj8uX/3RKxQ0IlF1NE4EF
TIKFPXH+tD4pM3SYRqiY8p5pKppK5PadbK5gaZAQ3V62PgWxRodDTrhxpPK/7Z/c4QjKkviIGrQe
L65IenT+A0/h9CXaY92KJcj/e+LrfJNdnsnNBsDupKAgQzS4d0DOclWUdoefxP3T4wRuC22rw1B0
QDW6zc7h76lIENIKiParP86V72Qgjl9aBtrug/N7S2MuTTQSuNZSkRPNYq1mXdWE//spd1HjuXlS
MjPS6drSDBexLi1rUIGeqa1njREaE90ksL4Z7phQfRIoOlVjuZUmxpuKb5L18LMYSzxinJOnh3T3
2KiwBGbeFkqk/GbUlo6jYuR401mGMc/qk4o7V+dyDs7jl2llmhEWU3EXsrEKJz2rwRPOs/8K2DdP
OU6Gdz8U/E+PS2BO1DjMgUb6LglsrNGGjGrYjKwhwdyn0lGE9mg8iYz6n1sGfQ3A34vgeo117mZo
WP4EBEJIerLREXKSWINMGCMZKq4fBB9GhhnJ95KgCE3iQC7EQVswbM0K4bsUZQFxE9Nz0s+ibWgi
LRymVLhIoTyoxzgrU6KcL10f7O0RAcP0SBuvlckG/TZFVe3OaQreKomZVP6VyEgvB/B3Q8ClB6i7
LH9mouAtssQO7yEwC+UP4PKB7R7SRxKPIlRxYDvwq8F+UoCbePIeHdsHx1+k0DHj9aZk8oSMXEj4
WTt3WjVxlxSap/F2vKMgc0/lFu1zxCzcT67VaodFlClbPMtg+usYZuiiTsWyUc8OaQ5Nx2k0V3ht
jDNIge5NRIbNG/8SSfWqKKobQf/om+N4CjgMCiQdm/BaVHaZrFgAL6zjvo7ZqG4QsIi00ziiPOAC
vxip+6dyQlRSCjcR6TajziIvTE0adXa6cePZ2hGTdiFaGLrdK8QQ6EWdS0+AlH12BNYBAcNNX73D
dNPPl/tfVt72JDhKJkgZDYfqlp34hYMTkpXTxktMNtMxXeq/2dsZAt6IF4McM84A4iscMDrVp2VI
t7ROgits220Emx5DPFS2Yg9VMHeYF0iVaT8O8iyICEVMKKpRstM+UTmk0aKbHdJ9sYxZM83rTsvl
FUGsGvw7JKkoEDK22NxNc3IcD7PlgAOlKa3ev8OLY7ZSaFGU1Cki6pWlh0/mQ57kwwdp7bsCJLkd
td2lvNFxNzjy8XvD6CvEL6zR034As6nx0WHLWtlbP6Kkyl/8uMEteUWhV4ZUXLWzKv7AO2JRzHiF
VhAl4FDpqVxJuqjixT99XS+pBww9FoP2yVGGQ6+WbufvqxF6qlfyTMu5ZMBM2trOyd1HAXnP7hvD
uLmVO5NSFy6UHRz9rAQfw5OzzWEMNS37g22Ony1qYN0GT5aJBenkWQ7KKoEj+b735UfuZlLymm7r
pzW5D/FJt3pktsol4cOXpGjvh8TU1xvLQq5+Nton/WXMkiBIk4Km/0OlkIuK1pWRFex/6Ur8l/0m
jhpiqIfDwGRWp/pbwM6lrqu2fDAhBpvOApfLKoOLIRTEk7Qg/kxDLHlF5p+5pPCL1koZCMcp5C6/
dhBq3t6qgUn5YQ8TSRRKZYc9iF7AGtzQOWPk2Bxo28BPhww8V59kYzaDP3FStJ9dtHko1Ra1K58V
ZO2lV4Fvk2INjILEJIfc7bqiDlEJbfYMa6mRSI6vj06EesXqhfjo108Rlg3RubZtqK3s+Vc6e+hL
cEJP5kCHzn6ZTGtIoTSZ/h1rBrygvYIOBJP37G/YckZDPCe54bHDt7IzK+grm0hnA20HaPafn6+L
5hIBjcGgeDacLPJgDKnfBik5KLmyL1IlpcM4Ii2+KUGesaNybEIZ9yFkePm9xzyw/a6SB1dr1V4k
IHc2hqVTFrGUDfqR/NBFCLCZrdtruD5rnGK5zL7mG5ScQ9e+kEY7NA0njCC0wbCzXtyPhXDO7zE4
b1pdCI5CIEYIo/A7FSB4sIb577g95FuQjJY68mFjftjP4AND3l5O1MxDEjlEYbj7BpVJb9Z/lLgM
iw9o9XYVUv0+jEhFoBeIpG5gjDX7bPTSJAMNU56JtmcLoFAEBqnJtxccFDI47m+bg0Bv2xbkn6dm
O9me2IWjK8YE2eUdLQGH0ZT7RnawuAP0jUNg5nzKq23aqShNtnxXPN593z97UxMmfLC3703be6V0
2A4NY8LKlegUmFG4x79ZpV3lB8kd0va4kQDtS1l37reV1DNcjjUHzJhlpmpKmxyY2QNFzf+X3P1K
2NZzFpD7kzVZtJccKKN1/1gJia02sarcqyJfxXBbSRpSyQX4rJ+zzdFlyuPZ5OmPpHug68lnqL3j
kiyugxr1pnkIjDbJQ91AHi6269tEpTXqtHB/paurWT+XXC1yn47LzTKXdD1oBRcs+6rX9NqR3XRl
AYHo0D+otu8M9JbigiFxfD2W7ei1tGEvY504H0iKDoudEzSGFtGVWC6NoKUpW7QOsSA+8dbvZH5P
jEE9zw24gj4H1TDzTCTMjFciMyudHXv0fNVZzXAKkdsEmdPHm0nTHSZtH2HryYd63d1pU3isw0Ha
8YORuIN1g7jW2JUM60qEsC8E7hopkFs1mP5GnB4X30TCAko9dw3U+mzqa9uBVzhSaDdQlOHy8kYf
5UUxhbBAqCW545yXSGaCZ7BxNUetkHoGZoUUAcxvGcTpWknWgDs5BzqiOVAlaSowe4g/CtLxKa6c
su95R8YW7pAZRFJjhaPF5vA2XmF2D+nmMnL9kds6E2DPv82UC3kJGpE4HQxuF5X+Df18JclbeDmk
9cDTIIcQ0WMgMm6/GGM5Zb02Ox0pxOVGnD2XLzeFNZIL9ra0An878cxBocCCwSppTvebhCZdTU/s
tBQFbQexxGUsYsDHX+ZzGRTudo/iyQA2Nm1FWANuLIjLP70254PdLuh92/X3WHSUSPvzLYeeV3RU
TM+s9ieiesXfN4YhoNGD8j5hKFvP7Gvi64gEFOl/EAaUBpeCaYV9+gJeUcWrX7HeCaVGiGyFmDIa
5V8gKiMadi8b8jugvWJI4TpN4AQw41G3A21wnYyfvXDjRFOPkcgTTEdtAp5SOtRtlE5XXUng3lf7
4v/kcvHGuiITO2Pnj+EG6nUoumbbZdw1RUlOhLIYKEUbHAVjmvRfHHqcyUZSVGC4e8FwQWanW55u
r+tZCa0DeV4JkFOt794C/RveEuCkX3DKsQA96E58kuv9Pc+NWdGWmE2TzIzgAahmLVkiDLUCJ1Jf
dMyKal1EbmkYxOQoKWqaAbChVOnr7vpkNclbnTYPurs8bMXiYHwPLIp4hhJZPrZblVId+fdvWJIO
Aoj7VWjVGP2enMbrTOCX+zlUATAtsS+skX2XQ802/d9V4qn8D+f2w5+3ld3JMaUT5t70LLv26NgJ
43y04naHKX4d7cO7J8wzi3NJy8/zHJOoA3kc4hP+pjlPcYC4kigE1B7Zwk77WyApOOyBuOPW4522
jYSVh0OPzNfZjWUnQal3CTXC1H9K6jAbQvPXo0Hg1f/qx092JAWdtNCNlO6VmghTT98TAwD72d2h
rvbQxDFBjLdOVPx2nVQhDT42ywVnku/MFIx1rWG9eb4euueEhf2nGeTm4/EawBChFj30RxgVvPPD
C2FufdPoPnPM7VQW/vVOvbft2iWWNyh4KTJB+ZNwnBnuZJEjhpyvfqlhBWU+EuGww98pxp2z5K+5
7ND1vOjRLMWlTTpqWhb5F8TX00QI/qJtr3w3ARn5fWyIW3xbirso2IqSJ8CsC46LgfhJ4+23dq/K
H7idt2F+qwGqT5OvWBiQjkaBtzdI9NEAaqbfrvlM9KIX7PbM6ZbskJoFLGkiJo5h0HIZrEjDJ9AK
2OmLXbqgpOjN4Ou1Rq1RJZGF2MgbKeac46SY4bNc653tTAAnjQVS3MJ6BnW0wyWG68idjCT2+DjR
2t1m3j9kOy45gUQYyZCPOpJGlrwj6iSB7QCoY43zwFCEuPZQG3uyVGCmx7BJjh+vhe+rMIN/TYWQ
yD1boUjVK4HgGJfrCI9TIybxk3gMm8FBwwKwLDupD/Sd8AO3MqFSvuX5nN0oQb9sNppMvDAyHK8l
8M0fBMtAjGk8LVcYR5w5zmdQUqx2KHziZPYXD9QtvbApOFePUkZcoauZJEqEnXmJ9yvzwLazhQPC
rlYWF1Z6+XkyIBsxNXKhAtSMUPVaN/BNBDWdjtmu2OivELkJfTl5+5nLYivFuXXtJkmbdN5M6vKp
ypEQ9UY65tIjcNUKaajE07vN2n1m/HxQMMpRFrPqyGIFf3Wr660/xOyLkCLf/enIMlfhkyow0dhp
Ves1rZobrBqbrEbZdvIRPEwrWUuJ29g+TBfa6qEAQp1Zxp4OB/L+0QCuU03Fx2tc0T2te66IJn32
0iaaNzHgO/Ce+5hSzhUMMcZVSB2lzN9/k7RUMxh3oGHqC25ZfPlawKEwhxyPQD+F79rxl9wBehfk
vRHAddauA1h58EPxC7IHEXakQ57vD3IZP0Sj7kFoXkF/WkC7pU7pcUB6vIeEVNP2Ch3qU6Oy1U9c
u5BQk4rbEfUpysPhKnDngCvyNVs4ZkP6476cV5PXWfwhZreHHMBGczqCDdWRjUJik8zvj8r2dEF7
O2xb5P95Sd+3KzE4Di8zqPrDRfZi1V3sXiYaeUk2qphlKROjjTUSr//p/5RpyWjJp5V2y9PzroM8
y+JI+Wce9S9l286C+YtUT1zlDGYqZqQCQ4DVjJpeSDR9HAwDQ5XSmT5hcNB1zml/qFeZFg4egO70
GbVO2Xb+Jz48GKt41qT31JVxrC/2c/Not1WgzDnQlAlMJqpc7P+5PbLp2XmKKYrn3Zz+fVwtdCzC
lVPgvgaxaq6JZsdtvdbg27fXDoycRQsHiniTdxjhpN7WQNJ4zcuzSbLGWlaFG67nrnaC2NRxdVqn
8aj4PLVQn5YeTs3QJjfuQdIvg/bjQ8pTagTJu2yvRJb3vXbpW1dgbNI7o8mF8eDrHsLm0GNdiOZI
i8lgiUJrAuXp2itJBQ8lB6rnG9520Hzzua4pNP5d7nCpN08TCRjh1LA8qwtV0QBSsXCZmjW4PyVa
FGWyfS0pbwfPwlWlEah5pdh4jkmKgi7vmZNf2nXSVvakTsKsTWcHPqF+w2tWbhu8xfXXhyWJ5Zvr
t9JWO5ia7+w/H68IPA6iZs8k1jYw4vBwwPACbfif/MRrDe8/tMFShGY+Jm1HH2GgAVs8NNuTypwI
e7jKE46TGmV0XsjOATu21trXRjM1YvcWkPrTNbt7ejap8A5xZan4X4tozqXuKQ/nG54HAwBPsy+h
U5g5s3bJmS0ebXM2MUiUoANgsVta395I8j4NveoQ17VYCztuszwIQeJ78faVwWWRyQgWfWY0pYQh
Gozx1HoOEnceaTnqUYt3odPmvD6aJbwXQ6sUe5tEc2EE8/p58lZgYqfh3E5c4YY65Bt52zO2ZbV5
zZLfDHeSvTtVnfjNfqdGMDNMGwigJVK6Zcjw9lp+geEYXCdtI+YD7L+7oYXrRnytdfLFwTIRt2vn
RabQMS63oQYX5uc/St2B2+aXDd2PbNfwce539Cq640LsQeNEWYHNHwG68UluHjdCkaMZhR0VBLN/
3IMvtzHBJPGYZsDrG6YvTBk1oCuLVA8nDOtdR9hgFu1U0bvVN12JSaP56wEKPOAmzY8PpE11/Qdn
vmlHHhg8rXYO5TrnSV6xoH6A/IDcxvXLXR2Qb3DXjFQ7ZrJVaQIJvzp7OMr2YZTHPyIWaUp2ROpp
C92z2sCyfUDwAjhsCug+DM2CvbtUiKU3D9Fv7X0hm0AREUuspHG1h6+Ket85h2OcyNLwppaQFtnt
Yzjqlk+N+7RQGriHlYNbHlQnaS+JF9dhuXdzMW8mp9cPIS+RfT09Lxrxb9DXbq4r9DF3Blh7dQwW
QU5h/CT9Vp8yabXCtzJUx4m5VaOF1+5ABbS2mEUOzGtSpg1tmS6JFkfWBlenfY5rD7zC/oh7NvP3
OpIDmi722yyr9N3Mme8upHyQ63Tz3VBdS/d/bBGs2LwtNgaLvmmDJdMyCeECQndoZ8wPFqght3lN
VjOAWoZX0Ow4JrXejw0XNodHGpBVJB5nFHJuzhS0+/jGQL6TIAjxia9Bh5xByoPAynkPy2x3sKiF
pgOIZ07+SFbQAo9x8qsKQGNniDVqhM89U/Sbf1v2shOwU6ZozLS2sIhWZj79HbVj3gZNzGefRe5F
wAbXSbC7q0LM/8h1+Dce6QbUUSPR6xV47C48Nj2I1EWP0fG2RiouaqTHmjuDfSwVHoJKgyoD1UYA
KuCFGEYg6UGNDgTYhbUoi2JzCe8OCK9rbWwcm0nz6bq8cSBqn78zDLRQs9ntBRkm0yl/NBmvCI6z
4ySq0glo/Dnvb0wdHqN2ETuutVyQhAG0JEhvQZnTb96jur+sqWllKVLtf5+ikxacX0kksz4fvXJ6
aU+A0zFA3x9stX3hcv1y42RvUAPP66ubyrDUxMKk3bgQISpYAUvaUW3rM7p2fQjQuXdW6WSGjChI
o+TObIQgCsHUota94s6NIb17oX5bzx80KRnybFTLpMp+1QHVrbFXbDRxhcgLQ1uW/tPcZmhpWlYU
GTNhxzymWxo53c7nrSxDcMfmo31G8DPXmFpO5Xtj6SHaZAgAds4CzFt8uBfJPTD5XBhDMucLQUyZ
BCe+c3QiaDS6Fk3FM3SBOIkkiLssZPrvrEMD6jhstZe2wdCQXkjSBlwnkEUHewXJwk2p7GBJHya+
m35L9CCKeGbn5LF5ZKPjFk7Cjd0RhbkJ+d/6MQl3e3eFgW/M6gKK/6aJSEbJGEmhf5qh0/O/cjcM
qTFMSYfnsGd+3dRwAbE3I68J/9xpbR3HH7QSNfK0Att7vsR+wTC4xbMEwsdd4GL3/tU4o5jImv0d
uqfk/TuZdV9IQuFrypcKoGfyKYiBVnlYcYI73v+r7xSFrj9KXc4Nze+IFgJovf7Yrkzl6hiYjbIU
8cFIBrNVjxys6Gkdy2FnOR72lFQ9TkwbdZliyzu4VDFh838oZEgYaMAQg04n3Fes+Z6KxjtefEOT
giP1Z9A4KmTz9F6Zh2Bbllf8JHSnJigURI5CbS6UBfPBhKK4TEDPuGo5mmO5bgIFdrE+cTJx7hF+
oC01whqVR7AvT46KfuerPOEYHHUZv9+tKRq/BdES3lsJNw4imGXWGu4kCdzAdpgEuW6h1t0q3O6l
Ww31DwqC68HnEjgG6iaxh9gMFLDHnYd4SxrPFX5D7YJCw88PXyMBvJ1ntB+JOZIfjv62718tOAHN
geoiy53C1NYArqANFn+FEcwJUyQte/3aHwFHT/9TOSuGJ/YO6o1zgW6SHY2uFXf3kbkqF5HUUFJR
LBxOlOQjYWWewNIqVtFXgdnw8KEwkPbFVVzvtlg3w3Jwi/WdjsVGB82Wuq4N5/Pefg+msGMqp/qP
C0mflip7t32hgBxcmJF4fZF66r5pNwn55xz5fwHprqozcbKh4aUiuDTAvf6SL9ou+oCdcSdrcNMG
sAHMlECz2KDpyBoF1CZsSYqfCke9YxwF3UYcWeD4HFS3IJFviLB+SLBjhGFbkDMUZM6usc8N+7Pn
Rsk+vdvVYsa+nHyXB8Vuzv7wfcSBFDLfsgQAzrKfmU2P3Jw2I8z6B7AuRT1/4VTbhtEpIZ/PYiBW
RxJhIi0WEID3HvDTgQ3MAQOyLCfw3xEgFBqkKDcJukLy6lboWlMzNV9j9EWkzYY6cBS6mfir8I0o
iBNpBvsEI8izrDQXq1V9jp38+0JdIKc48Kb1mUp/0h6pUgAJnIUY2siW08WRwwh4T2f5WEVigana
5aWQrt2U3hUKsEc3AJrQHzm9gPQausfX2Sjjp+ntpz0P9oogjhij7g2BuC1ShXWqrE9VKkEJVbRQ
7eIwHqVa+4bATHDa1cO05gv1h3i5WosVosAb71Hl2k/tV8ufsV7g2isjS6Vu5J/4T5+q+jaWFJpl
y4jU0z7hiVD8gzHjg40GlyE=
`protect end_protected

