

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
AAcalZ8o/jQY7YVFFozBN2W4CJ7dtDMmc4qCXcw+X1HsQOWsjlnqJ0ExLq/9HwwPaBdBtHuX8sNt
9MbzT1NoZw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
eb9fumGdx5oOSTot8dVQVSjhrvPnjy5/uUjD/aIEqv1QEwLJo5EU+m6JllUu7ONkl4q2pMcv3yUD
DaaWMJ5SKNM9IQtYV21pAAxck+unqu58lsMHcSYeRXYcYP0huhB41kbacBO7fQsq8URHfGRa6NSF
6GxQzFgW9OWA+QBW/NU=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
EWQNTRM+yXYG4PYEP5SycD9fkQkTTfcM6sgjpG7m3z8pRk88pPYs5UwluFbB09hVSCMPYEKLENX1
JIPX6A6AjJm02cmQD/SZk/c9uIP6nVMvhv4HT2PqiJbMwRsRLnp0RV8WJNl5IwtzQhAltPQm5tcZ
c9/ABn7qb82RSMRxfzibhF2Uc1QWD8PnV1j6nVmyG5zwtPXyKG+iY84QCANIn7Soa/s6m+bpOho3
0pAI7CU0STIdsIAbeZ3h93cun/ow5TnTga8aw0A3DbHVrLc+5xM9M4rs1eiVbJSSdL5Fc7sYK0UO
cAQhBC40rZd53OFEkTfLRVfwRFeSU8VoPsBCag==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
EUZqFPEsLcyFBckZdNISKg5E9SpkAkJYhYdYkwRh/xgSz3PN8kMAAO+ttVMn672EPHPSTTeJWt1p
AvumrJCguaLVBM7NIXSVbD3Ckha5a0glBfzxCIJFFOPOOxZ1B+rxQ2W+YUfoLzcw9DE42G8bHsgh
CvpFN0Szn2edsSc6Ou8=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
OK0W/E9mRq/arn5PVxkw4+3w3BGYpl3KNYb/ZgKXRQbbZBHdfBtfu0H1VHCuj27qhD0QdkPpdnd6
gHcvGTEag6clv0PLJ5PHHHzcIl4hIp/MStOr0nGLUPNhqZtLAZRqiy0IB5ktSoIvGu4wUrWu3P7t
D9RQYPlFcbj3tpqdazX+5GhWSHnpe6FaCtaWmer4ZDmYZIG1oGk2h3p7ggKQ3amLtCrg9RLkGQQj
yEO/bz1jhZ65yzQA9tlLPbVh4inksrXMkvmJzspRm61mhZF1ey8gENJN2v1TzCuN2XD/gXtMbo1u
8igS7KocN9wbd7hsHdkLAK4mTBcgTG5pa81agg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 998320)
`protect data_block
NRXSH7m1PPMKOIViGVFUum1NOBkj0PJ62hEQLQE+fMYpsFuyVsZfE2sTJ9vQfyYlzqSSZNoYQwdo
8tqJpf8fXc7675c0S7p5c0RQnniTdxsoT6oFAnpQxIKWBoNRenanVZl0r0iJLUMObPXfpIuF4vFS
MX6KAHHCEpKERo/y4efH6v54gZ3VQ0FmeyCV+0i2E/1yh06JiPr6DHamoduze5go3+B1iKky3fnW
3O7yc6vR/KdnKr3vAXkXmnZidUwlzF9iegLNTmd0LmOnWlzMx/h2hrEGSFKApeBKeby2ne7fo2Dv
YzIEoMOG/WL9Bkxs0QrO6hBNZ27CAcYD+pHhZ3Qf1VioP0Wl6FVdhnqe9Cf1DfNXpWX3jaA6NJYR
10tpCyEadkrQ5aL8XeNcGCIydGcVshDfFl+j1VLBu1Qn6L/2h3ON+ChfEKtPFkrevOmESRlp4dlx
FQ3OgqSd9yAqj69YVvojt2Tf9Zgtg7DMYbC2hgOSRIzkUY30m3psSU3+I1ike5qEuI/lp8Nn5I69
CKGwVheN6622nrlz3pwtttZc8fObQOhg+wdS8qRB7vMMKaXIoFZ66OHaX00TZE+2AHt+qOGcOU4w
m81JNL0U/YnBVF3nRnMryqm8vxQP6scoKV5t1gOFua2RzgSocOExe6FP9MLcr5d6rv7/iS4IxVIM
0tnVqUIkDT+Jc1xGWqgRHDLxowcdeRiJ5oetsFsOzyj5J1LE/90lPzEXJa95OQ67XahX7Nrd6q+v
Vs07i9KngDyZemmdnrAqu85VG60JiQT4jYnsUhozZioNBgrLWJwSkxrHGubuAahyCbk9sYWgSrzj
9+nEcfcHA0pLuTWvOI4k6PB8NCo3+m6xpNvyWazrteoryQqnTRb0eTAykQJQl2aVjkJgatnYD/GM
eqJ7t1AzVQeEtrMjO6nYE5mgdyH92k89gQQFJA/BZ7er28ZUvkQPPU/B1A7bpLxf0W+vuqZxLvPz
EFBjxXfug3HbN3r0lBR/WjADWdsPbTCaQiksmYAEIg55j8rANc5wqOrtAdJN8SIm+awDAkVmFKNt
Vfj1f9IKeKicGvv4otdWWqMSqA2qavHm/rQptHlX1vehtD5MNAz29DmozdyhTo6NglY18n/RE0O5
TTGTBCV+hjE7oAu+ZHn2d6zzzrtuToouDnOQA9NbweHy3KRR3YMISVs68s2fORpYYZNDgr7n2dPm
Fjll3qiKuCESDlNCu/wxoodfW7FvXOxhlC6UuzZy3dYY9hDd2aiYjGk4YUF4K7guqo1/23wQSqx5
6NbsAX+yGudR5J9h4y3RWrZmVBTqpaqML8xN2uKsekHqem+aA5HLuwCxz1KiE7BSrD4WbxEK9PT4
Nu35YJcygpMEP7F+s5Klw19XyOKde9n6W2axg+Kcg0PjlIbC8XAQzQx5o+5vJAnMG+EizhNUV5RI
SqR1GUi8qvrrFFXiaVwEZLerNNBFd/7+tl3/sSZAUaXlmlIubo3OM80MeWG8bHPK/nA42FsDyteU
tspl0tH4Y+e7sQdLvk2rM6bn2F1/qAeptA6U80uCW1x4fAPs6r00xpsVs2siuumcvWfPxUgXF+pA
3XuJQtmnA7C1dGzLzrv8Hedy0MvMxrPH0cbfMDM75nhPZ6bLTHObO0j1wmzAULCpLBunzsB4A/J4
8ZyQy1ekgBrmA4AYqHl8S2uEvLloCPeg80GlQPz4g66MOqeR/79TTt5svMI/07VkWZXDAVQ595ZX
Nl0+vSoIR4CYWBNpJgatt46Jsa+MKt1kzd6kfDP1rCm9CdUlnf7bymG86yP1ruZhnusEWBVOWAy7
mGgeiq3N5Yuth6PsFtmm7skqrn9vXUDy2lFHctaaVBPK6bF1EHJE8vtuHkBSJ905LvJCbt+zaAzl
DSOVYulTQJQ5H7bRwGi1bxomtwNeHbYfmuFYMtKN3/Dq6tTv3QKoWGeuw+3JtQANSF50LHvl2KC1
olXc/C/lQfxR8pDda/YrjT4zJeyHhDqakMi06bqI32N3hc6btKU3mrFUtcwWMhH9gLj0H3bZuhIC
vvWSNz7doFmSdFataXmcDzh1BksTdR+uP/zZ1hGLhMyurDRwb1bcj7bGwRMSe9Mw540rpfEsDekj
5AkIWi74Yn2WBMyaVH/ArTNOrzoAQhLvpv1e2QJi15c5GP6xrioWhWXNfk6wLZAJ/W8O/AyhjxPJ
AritR3kCvTaX3ionqZyJXC6Fq1liq8mqbHBTctu85jYZEUv3GorCtPLHL7O9kzHfWOkKmljE3F/g
w67Zqt/iqSWQQ61vZQkFALLgSyeOuUIFCaQVL39DOLH3+dRD107g4VJ8/llNlBocLa6x3omoJmJE
g+frL/4S7R8r+dUs9E2Gcdwxb/Sw4t6n5TCXcH6QNgLP3jtusqCvTBRkWwKiwZLAMojZBXfq5Tmh
WvVBx+4tE2YsUPFqKC3FCYFetPd3Xl8OhPnlCBtKNSQ8H0J2Iqke5Qd1RT/WoBgGB8GIQDaalX5T
ysVtmuJKDNwJYOiGbpqsETceosLvQaosYHyDcYjeDwoxrhdcJZHS0LF3ufbYfoFfHklKu/pbeeCE
1knnWJ9jpG36skpqoZkLbNZRiBRA2wuyJu/EE/P/0RWV0y4gfHpaEngslpQGj2ReYJgytEeELBEb
9lbhryqGKDEW405kt27RnEog7syCTkU6pFv6veyT3MecosRkX7A+BTivWz3jy+MFO5kBtJ0LWzh5
mMF56kSIxlrvkqP226nAp3MbWWNEz1Uh2wPlYwtgiZM/ixLdiX4/e7ZbRGwb1Ps8O5mHlN4P4D4l
2qtjI7ZZd9s/xUpqIF4csXELxNqzKXR98xx6epPbiPNjk+3jtvcNfUlXP9Ih1eYuPOFmyjFiSp5r
VPyXPNoQ7sjMK3ifJ0pRyppdJfs7n9BBbxq8wAJkW3B+wOcT+k8t72gCdLq6Uy66K67KKpgETP9r
zJdsVe3aQI7MO7b/nZVOsi286X0Oz+y6HcQSBNWfy7iSHUd5RlJAeoRe2rbQzZyq9P3K6NtuiZIZ
c1g31Nr3MaLRHZ6PFXKYw6KsjCr4vyD7vSLk9+qMc2HjlYA/KrjWnnkPKFzRbesrFarZtXzhYCe1
1ZW90/Tlzg0KpbI2RSyJgznh/eRDAhBf9EUFVAnpqJReX4INBNnM8UQzbVusk07mNcJ3uYeeRmBN
6ocF5lcikwqgvjqt5+zwR8MeicIM65ej1rhCk2f4qscKqtV2JlYppjaY1ZwIn/alwj+1aLCduJp7
Oxdo0Z2ISv07rhHqnLPGINCyKH+BuHeng7Cn28nwWRAK1iWR4v86uiUbQG1mNrsjs3Gcns1zrorC
a0eYcAdsc1VfQ8fLm9UPxef+dv5R0JFtVcEXzGOkMKk9Z41bRmfdQVr3wuRkGwxfqrH5uh0jn9Mj
1DUPQ/Sw/rxrqCqM4yUeDQ9uXyCbR+dX3+GdbExkrNlhcL7d6GE2BB0idiC+UpGTmfy1bnrYvsTd
MuIEntJc1SjQHYxvmHcaVRTN79ildPY7qdNyehL6SFgpBQ34lvbOz6RJraDmSRV5SUPYWdVDlgHj
fgeRZGdEeJfg4OxXyVQTAbqbHTxaFZC7BG+TAZIUSa6GnSF3LSQD+0i1QfVb2AOBaY6FBbW/5U5k
j351wElaRWTOr4qmfVc7JEMhCdlwMU6zmnw3CpbmfnFtqfcAxbCVW3J5zZWEbtqnZokCJZL4HhME
PKGpLr/hQLcJ3GDnRvPEBF7kCxl6xKkFbQrxDFNiS8iUrZ/SHS1LAVm+w+GrEHPDAmgqK+niwMLn
k/Xptk46zN6ajHR96L/JxStuk1RUuAIOI2U3o4Bm8dilGddtwOr7zzVcKvrD3J48tiWBr7xdBpO8
0HPxhNXzdjGWUA77cWtTHLvBVW+rpJVEy0wIDavgsEf4DQCU6zs+Rej/vUt+5HUiAN5ZNbb8W16T
hr0tUK+fEsHOKD5uhb2ulIWNLYhPTBJsyqwnjqXLuwlJwStDY+8ndx66DZ9brJf7kUz6mgdqe2jZ
DD+JRFVf2V/OA3jPvnXy7wnKwB9MiitA9eDOwyNeMaLs47m/XKDZn09uYMlYVGuH+U6QODv1CVIg
AiPMfwr2ZIHO6cadHrqNDHHedTQgoAT0aMQJy0aIDfHJRaljleteJEfnJbhTY/PQsniBsWrSqXPl
AsQQCCcQHMli8WXZgt2aKIYDTSCrrnu8h86Vpnvz51JJ423un28+Fa13dbd5kmNm3MJM6dkTGUIo
+ZQ8bZRM6rIZwKFsJqQ248zwz42oqTDDpJ3VWLrcpSZQF+Afhyrlz6Hmxg1G5THjHzTSTsyR7G0w
6ceL+FdjOCIlJbeDcYKhine+56L8kcznpyeiljBgpAI2vfWD58RGmBBB8nqm4Gx5IVOvCDdu6AkF
rLZmeujqfsSqgeA2wdGwQlvImGOfvS5QJmG+uBehAUMV+61ZbcOiD0Y3aW1n0CdmOo5E3lDjhmPX
mvXEAuBd1ZQyMHHbNOSu1O+/dWf9ITR1B9/heewqtABNAeGoNFg1f9ZPK6JOz9Js28giTmy0jKHh
LynOePrEyqcPULJ8Otpfm15N2sJDlCtNpc8qKE6is9+hwRlgl5PbmQnobMeCJNbooV08jM3g/5pP
Fti+DIaSF4rYak1u42g0YvKx+6z6epyeZaoGVWTgUsZPIC/EQAZsmAJzIrxYoGOc88OW2K1hy6Cr
s3MV5aLBLungODsPdik+joJTwdwi6TPIg8hAvM8Rny6F/Z+cjStdDBRkO/DfYoQOqIJ69NjvraVm
ZkSfS0CJ2Fb36nd+M92LU+JIRe+ySKrsUhj/Kpa4//2EG+AiWa01qWudnThn3aZQbM1H6seSgSgg
T1iIYcty/Bih673w3wPa+QaUVH8wkbLKXP6fDw5AIqxWcsy1VARZhcQU0WN8pkkaUGzrm1I+so/8
p1/Hf7iy+bu3uPn6UDbpS10U2Y6/cZ8DlzZec3oeV8gfBSxETeRflgCMPoOHNXOFqRVVTyd4aMUe
zx76ffNRjq8bFglBRhJhtBB5rqxpbc9eE0ooNw3jQRkGEmn8d3hFqWf6RTwMjyOGHKqNLAR0Gd65
LLUfLNLxuE6M3WAGZ2jNDmvjjaqaxW9G5IaXi/TPdLVzHpZi0mvsilcKTg2P0pzUxKlJi+/Me/Yf
kSzmZNi5h3Sa329O4Nqh2SOXBnbfY90GedJ5zGlD8ZG+lWGI9BXisruxnbCoMpVn2byN4GXcQvE1
VdWpLJjctcFBmtkxNREqufJiIo16fj6m6yUmn4VOD8jhYwS2y79a89ElN/VspIw3uuQawCZ7+rSq
5qgvo2EXvgEMHow6ZvMv5EsY5WS2m2Ap2B5V0UZtqulkP+iQ4bvQcvoAt+KRXNiF95f0Vfv8DxxT
mbY/K0RHcCRekiWl0Tdl6JxFs2UVO1xYBZBICb62/S0fa74LbiVfe2VI9crp1/Uti3r1pF3V6Xiq
F1Izb9R1AqAtqJetyDaT7A+0oKmzk0JHDJbIgbCOMxnzz1FWy8GT0uvyZv9J1Y/ibedlhQ+vLK0g
Yvh5xbbUBrjzswOC6JD4rgMNgCLbz+9B9NO1TMbapStooAm/yRweI8I3JJwfWf1xqSpRE+3imRXP
DHkbrA+sT8GeukZ6snUPhwQFok4i5XJ6e3z/IaEtT2pFdUlNA12GzZrnDzOqDk8EwWIqsOgg7ZTi
rc6jJmYQs1Ahq9vK3CxgAxgFG3qsrkdWOc0ArkIE4uEwr7NnTeYF/Bh/VMyPgAK7IAXeNYAxenHT
NnP05OHwx1dQLEpEGl++Cc95aUWNAQKutPO86CYf/fNBEO5YKhpkTLXdZfV7O49AH2qu0fa0uEBo
bdIoYpkYens6N3STpcWwd2ri4pwrbnwfTMu69hg646Ezp0Wk1KkRVLxdb4eeS0iX016W/dhIMK1z
TuAS4YG6cr4tmhImwK4tcFBmTYoD9XEbhU+FIvWWMNF+sZXAH6gRodO1lNH7AZ3MtyTfW+sCmUPV
hvnm0iszfIToupwLxgxaKrgeoiKzFlf31DHAGYXBJ8on7VWux1oJT28iG/oKnoSQpHT0exTR+fF3
9q8xapYOODlqqQBVNbVT7PznRYvOq/bN8jSzYz8SEezLnKghVGvSx5Q4hbz1AopNP12R06N4Lf3A
2Zp+lCrOmIOvElYYdzvj7a2WusvMpBqDpVXyz+LcJOrDJQGFDi81apMirwzRcvOUnnd9ubgIVQFJ
HYJV0bEmW0uBFJEk5ZbOeDO61MjcMznF2zcVr7oJ3MMq3CtkgI6Vatb+qdUWJS47pMkFDaEhyTZ7
EPm/rDC6W+aDxsbF6sky3Uu6CGIgH6YHkec9o80aKSeknYiSaUInR7VxW68JPTwH2pZ/A5QIW5Qe
ox2YDvTxXae5C2tDLulDqV0fW+/jdNKmn47OoxHMZkAz9Iv5Cw82hOuS3DTEqTe7DVVUTC8TuXpT
q2GPJmJKAvw2RMe3guxuU0MSto1RJnryeMnTEESmnwlaeySCpsxiuK+4QHQDp/69dkYnwwfCCfes
EUwiJYFCSuKCojhRDgRt4f8bsanjV21XrsZRM/XJRmsqzTiJlsTlS74BNOwZR5598yByUn5a+WXm
Mnqld6P457uc/d201w43fERRkIsSeja7EnADms5W0YLmXAWy0bklT8rLTKtMgKtb+36qSKh82Bx1
LVgC8T+hMnSQ/QXv6LbcsLqUtWxos++kGTPtmFwBsT1kOG7q0Jt2XeyXmIoIEORu43d+q77ILUJE
ERp9D+666n6VulF69ln1rKmzRy7c4bDpK/yIixH+Hwd9NdGAv8FO3nG/sciufcwoQ1EMb78Atc9O
mA7hQEMxbu8am4rUCfrf1OGpmVohTxRL9+7WZ8c/nxUj73ljZelHSRL1PQ1Wog73Rf7Q3Y6rLBIh
+ImtcSRO8ssSj5kEa3v11LOfCGWt4NEHqjck/eegFi4TO+lcjLmyimwd/I+2AFPnuqrZxGAy/vCj
LQEIpikQchipYBWuXuM+mRTcLOG6TsOVf+bVbTEeYGcHsOVtKH+ReD8mj+wFU6oJkhk2SZ+91uGW
bPAl/rBwrJfJxa8iy68T7yYeQNzGCln5PZa1wBCOy+NruQUJUFWrvde7LmjxXigJAbOCAsUw7RpH
lxpjbwHV1DYaQG2GuIc6jJweE6gEXy7or0bA0iDiBt2rbEyGaftbSuWqzu2ZjQtG8pRhyI0uR5D8
6WelNxU49gOD9eS1jtkJiVRWGaS4x5Dc0zQCAUcEN3tXA7sZ+mJSBIhYcc6XWNLcmAbZV2bde0V6
bH69GOckJVKzvKR94tJnjOfwmpmg4BwQDwoLVYJOfMJ6O8uD4Qwk8TeslD14r25rqZZ+Tug/G+k+
Sx9zgJUFWFUKFJMJbXXe5gveGlxB3TZsrniNt1H1dbq3b6mWj/JhxTfTf0L1+mIZNaNu0PKDFiJC
ViTd/D38t6Deo60q1LQf4oE7fxZi90/Oolm2qw/wvZVyq+1/v1BSDUYDAuos41c41xOf5LaCCv5k
1zmfh75UOpOXtF2GPyK9kXt0Ksz08izAdn3L1PZlqz0QPpvapQlA9C9K+GdBHJ9vTMQDroRDHeaN
MON4FOFvilb2WL0f1MDCB0gJ2VZJOjJ4M1tMbwzGFs9WcI9DwGNi6USP+sdZtDLXUE7oYbPTfGGm
Rqoyg8C/EAJ+XJ7iasjUQzfPgxz7UiVlXWsxXimwYw3a3YHqp1dTzGh0zWQ9AJ9EzXsl9aFBmMX7
MXI6/uU2xfSuqf5HqOFUclHrMfifOjPurN+6QoojhrM5cDD0HHUyskFjrpaIrTRzbkoegKN1KYFG
XTNEMmiauWa/IY+Um5/MLWqWM+hpZIUvoSMiEWGrvJQWAnOWZgZQlM+P1ALlsn/5hVIzHdXdC0lV
nxK7ofuTDDOQkpfthMJdthu7wctfd2cYTIexvh92jDxKmZsch7PZl8MOjZuqXhtH6biUeHq/ixjM
EEIS/T/VaLTsvoMQXZUV56XdRHGd/sQzbb00jxogDGyk9nJMBnniRZi9+tEVND30tAeywfQK3FT7
1p7CgHRqyy49z9Y0DD+aJVP2Il3jIM+vLX8/z/1yfM4/YYDh1jGwfct7MQEJDnX+sslN9L11H/Bu
7rTDf29jy4pLXZB6HwlbgrgYafYXWp2DJL7pwOOW42XVRXB8PEOyyJX/Ps5u1ibCufUtCQD4nwab
dbQt+u05Gvy1Trn7/YEkOhrKf19s+2/nv3jDnmGQu48AicEjxvczkOQZsYDr/OV6bJQb7cCm0ecK
YVYpHXUvXH193WsLqVS0OYvfwwkLySz1UZSIn9jVCPDu/d5Giv3Vi+HqzgY5koOgqkjDthbpP5X0
CTCq6mdzBOEBrqT8pZmEWCSsKPL1TRyH0YX+dKBlLYtz8ZVXFk6Dcz0Kud0LI7/2Tl+WDJ08+YWU
i/2ouQJquKJ4IZNzCabPyX55ZhKiE3tQPa5PREf2vJQ9UTzduBW1e8VwCzIAk2nBrS+j9pyBY104
DPAz9g6BzQ+ggRMf6FVerjRMDjDuRMvq/UGz2jSBMivO64yt//0CIC73IxYWdipSYSvs0JSIQPHu
NKIZsNqpwfN/disCns1Pf1KC+FL1AFjhFlJnBlBAS79SdMdLVFcAAnXWRA2ZeNNqnEfvKBvFo62N
iV/KsjW3r217i2ptpyVht3F6IU1dSONIr7tzKOipAsPPTLh2Ok92kYKuWVYZ7Nfw0VzzL/7FcL//
LLKPr9vE8ZZudiXHEX4JkCnLdsCOUsROUNjRyyIbJ0ECaeP3LoeLe6pLdjhk0/RD7qhumKYe0Pd2
ht+CADMz3uBb01NrVHilmPUOw1XQVjmZNg3V2yJ0HoTII5IocOsNf+KynBUkA/EZw1LUrVBaCH4G
9H/y4rJlRL6IDGcV87IRRSOQ3ehb2S5ulN/qpUM6rLPFftYrvBW3MfvgJCQKdjLAcnU8yD5rzw65
4PKl2CsU44AB/Q2k5N3HPZAoJs/bXunNs9zWGda6PH6FR4NB7R5gCYDeYIGMeHRkimtwo7b0OmSm
wYmEVBaDjSWvgPVbFmdbnZjTgdUvE2HtQClLNAd7JM/1DteAnfm8q79Ed14jh3fWntD3i701VQp0
UQVnEu5XIvuBJztHIP6tbQNCTT5ZBkLAZBPZwFoQ5uP4A41u7JFTqrhf8+NGYNWxypyZUVyzJq7B
PCJfyvC5hu/q0ZNmt4mAT30WWoRXuCdZw6vHq7s2/GSSdlaZSIz65R7zx4rTovXjhBFk4WT5PTaB
7SvRj5yJCPS0znIBdBipZHAbLU3OI3YNAnxbLsFg6pdmOV398VzUwGnByVZklydyHmN0xFAmwSp5
4EYaL5AkYTHrUpKoM8WyZvg4Ek1gOlptv9JqV8awXjpaM2RFbdpD2JcUc2eJC9gkO/16RJuIhV4B
jmHniovTgijzo/3x3ZI0AmoBAZiENyirzG1CKR4UrJcPaMhBz6+9AAJFO65/0AoReUDGJsX5qJpR
XtxXMxjI9vKjY9Gt8hFdpI9jq4oSA8lu7I1CShzihsFR7XFi8edHMavqjhspFdC7amc4T8YSZ/10
LECfJ+6f9J2a8mvZRJVpxXkW1dAQ7Cct3BxloR7WH9+ktI19mgktxA3QBGIhtTlMrQB/mH9WWNTl
235FiPZhS/05tQiaXOv8HJd90J5KEEsz65VPeI9hpvdekcptNhELGDN00cVEn11GaVp9qdH7buD3
gHnQsCDhMo9AdL8IKSJKj22rGD8OJNWv/kbfbG126qSjidwOEz0IO3sddDLFVxc0JXykOtwZlFZY
pmB7vgxNf6DjCse39MLI0V8eQ+C1cDFKfZuv+EbexPACdIKL+RSs8bK/GAD+XGwTy/MeUC3a+JpL
R2Mv5ceaI0mhh/0czEV6W8A9gfRridSSOvpzCGFypZvFUM8rvNmyfOF6uIe8RPwsDuzToOEtOct/
OvJQO4cE33co6KZzwTHBJWzFpn9VRPDKekiFuEUijpKwSy1Z2uq52fC4dzzsdW1sCPGKdSR3NjaK
LkVGBB4wqc+lv7dnANeAOsXxqfdO+b2DVPgT7OZ/c2eyJlafDzAsFDddXjDhUjpM0IknDa2s+qRm
I1eUcS6kXjivdgG6R5udUJXO4ODwqATZ48B4YyNnPV7r19yQJvt694KB9MLvbixKx8kFF9tJsWip
BHJsu69gYFvORxo0iBZHcjAX3UHpqJiERVRMsD2aIe62ftKAzHTJTR14z8GHzE42g+fZY+y2qvV+
+fCSHLMt7e/TaF9gq1Qm6E+2FNk2P0qBSH3LqQkh97yBiU9iHCOQBHsv1h1oUXKUF5x16uuifdHb
Bb9xw3bqBp9yhIj3Iq6UezRLJQBGVk0bw/8vDpQshGduLx5dUj6DODGQ7wJjSptQAn2rGEWeiwOO
NZHBQt0tUACn4Xh0OomzV7rwmLQAp18ZiqjJEH+BjzFMFPpaIyZf/kSUfv7lLEdxRdq3GYjrLtjX
lvZWOFGqNeAWXnVUJd/CUpSVRPFbQiPVxlVh6/ars9BHC0fSenQErO24imZB5SgcDCqzcBlmrC9Z
n1el7whQUL2li6TiLfsmKxtR0Ni/B2mIDw4JzYntu1G08cdma1Ac9XXPxAKMB+U1DYWp4Y6EbN6m
YxUsvvG9Y7/8iP2e8ivnC+axcVqc3OWlIaG6/cX5tCMcItY75NbUQo5w5amqmgf3jg5mnf2ehAVg
wIkWTKoahHOi90PnwCznF3gSYVoyAV0bzDbkuqfVxO6KEn/CLfFXuFlmZB9puDTl5jetb3ZNQKoZ
jN570v9oM4yuEDZw9ZY/4DN1Uv2oD3VCLAd+DPzk3E3ooHpEiUqA8L55gnd6y1kae6pHwZM5ulhK
5qEGKVJ7hgn2Lmp6u8NW3zO8xm+XGAbRaYtiSTt4VVkdGTsAdKnwKaK+QjqrLPgxOxDUhoYNLqjm
fvNeuP55/UrYygNYXWkD9hNZYjRPSoKn3ETI2M6wm0i1g1gcxTieUpbH1Gqm0iH5zPIUJL381otf
YQWDMrO0FNZqlP40eBIJFuVI1T6oQGEWPajuzNFKc8Z7AlCIo3M/8dZOTKA2ZJ3uZu+4vVCNqwoL
cdrT4+icOhI015P6O7tKAeECU1px0OpBbggGeIEHqFMGpzd22vKRSKCxsZkyc1n+FkJ/HkPsX6Mu
PHW5J59MIyNa7ZPraQryGTWOS9MThITsEIHMqiYKkHEo9xK9xCZFVjhiRL5M5Uffp8IS+IqPKIEE
JRNbCcXTf0dIdGkxgMRiNdmrTzDdmXUvGNn82AV5nnqefTtqgDQyKmPylX0dOY4KtL62+K0aC0ut
RNpIrCDPmEs4qutNH/Pa/XwRALZwJYdz/XMA7XAMFVuPyjOBRsPKgUJXRpVL/f06CF8dh/dRzQRv
WAWG5rw+iWtXIEqrkKgoiWKkH+TEkO3bPp0pfj4WMgTi11TsQqYFh4DoLSw/WrlURJc22QTkl9f3
diDlbUcUHhSSbQA7fdzU3pzvh7DlKjcDj8ejiz5hxOf/Zj3FJiG2jn2Eudsa5NBMlAFzaj2kLe0B
kF+XYcvcx5z9LNz7c4oohipsx7kf9WP+3TO8YvMt0wNth3gyO63siD0ZJ/QKD5+XchraMROzmoOs
op4QFOk34gENkJYOjqltvfZYAO4GybTwMoVBuM5qThFTy58sPvrXyv8unUEBtVsWf3f93i/mQqUq
l6rjWoAG7CLurBTWHhNrVHHQv3Ot9IROJbhN7sS8GGyOmjBeFCbUyqKDGq/j/li3W7ir1iu333Kt
Kg7SktMpXC67+8PjOw9I3y3CPxbu3HVw+4WCiJFQpQpM8YPGczDPpMnoURtr4kKVhSEIpLqxv5ff
/RXSOHCY7//Kj5j81Uug3MCRRMLCLSJajY96DNw3rmCEWlq2IzYgbkKwp5hRxL0ticnysu5FUuuh
5pi/fV94hVCqOkg0++v+zYDHMULWJzTP9vuwN6F49AbuQf5rAvcwckCel9E0dGDzLJw/ewrTTNIj
Af4Rb0FASM8kL6xYdFcN1KlLdzcNe+mni672TG5AsY56RhpJwEeB183cmzquMBz5J8RLXpbPl7kb
NPUHtLxAyMeE3mdLOKwPOGnCtsnAX+oMXD0DDE8n7gLhQI4E429HsRPxx8giGPe1qFmsLmEssi5a
JTwL6tnFIkJ+uk6FcQSpoYUjbbId0px6KOqR1a1JQ8+Aa9WSAiE4F7v2qxShshlb4ALgmD1hQzlb
stSDqrf+KwVsIgY3c3Yjy5cWr6JPTLq6gnbCOfJVlbJIguL/u4/Awi5TFuc5W8XDXnwmId0o17ro
l4FawC9orzsH97W9gx7N+gQHYFbdIr/KBqcT8QM8nQv3UzAZnwSQsTViO5mnWE3gFyE9YghKuTF9
g2rmCVQLwfnx+PTcXozP+/5mYuvECa+jiaRx0VdKHL+qk4cqAWlUVZeSQpPausS1LIldHTENZh7A
G3DjKTJsXOw956PlCKGea4fasEJTsjqOj4FeuMGmnry7JKtkaI3xKFknaDF6DN6+N3tYrmwvlVoY
kvdH659NuhK7f8egVEJhiMpYoHE9gbunPqmOSkmvQ/zENFWiSQJwv+OZC6J4+e4KjbByHvSVr7WQ
k/WcGUsgZF/pIujNMXrjx66v16wsgRvOLcGY00mr4JlVcbac23AH/3+aZpioslCb+HHtM0LNWo/e
PbgwgjwvfVwi3ceAaRl8xj1I3+rEW62B74hu4v1AXnZejdKfVVjPl55u8yN9fY/AtLOx7XM5blV5
+bYrnUtRygY/aPJDraDBP8Q0z4Vgw1iZNRwHqvg54LzI/uChHQNS6qWUAu1KH7LgAFc9YHrHgUlI
+adRzUGYaTSkOKmpRRvG8qB9nNq4kv5bDJheLCOMqkgM9sHHJz6U2x4xrXJrz1nsy9W/FTa+UrSn
1vvOy1NTyWmsAWnk8fQIhTuqC7ca4cZx5q2L+cGqp5HKmw65DPG3J08uz46NCzifgAuTgiOa/Ffx
iryL9NU5PLbiRTJip37ziaitSRNp3cOywgQ/vodaVBIyK7Gx0rUJL5fEIk6bzPZ3fy+HCwz33hHk
Jr0uosnsoUaChcLNHfXyGgycDnlcsaZh1XLWl3Bolhg17IWpeg1hoyWZN6RlwBJ+zIxjyVFM4kt/
BXOKktYh2QA1jwB6wwSgqZ3AZtFtdbS9TBYSkhrPiPLAEFE5+QYbfUBZxsMrMtaBoz7pTjXPl8Hr
PbWNNUg0tdGZMNaEqfLqCgBM5RHYkkcTQv23l2JN1V19hPE71IJhSJ2ZYftpOCsOjjF9oeacqrhB
OQWsuW8MLzsQFYnaSFKVmb0zJ40Cko2EmjDv2jzYygKalCnJl2l6mNApmRpOdtLWobEHjTMP5Pm7
OGRUGPQ5pfzh+StK44XYq3hE0woBfTPR+TJ9l0A0rHHpORs9qaVD07K0jxuudug9TEaehniXor2r
+etAvrmadB0xWZjPtkSr5epoiQKLsXsucuuW9HKddT8kLDJ9KV11a2vQcr5FteZw1Vt1ukUBo13+
HbZu/kmbfqpsXk0do5cKQ+TVdShNlRST7xj9PGFbA/JBblXKof+VX30TtSYY39m7ytngtuhTrkT0
LWMQtQMKXS/mSCBcLq69l+PbfgATCrMXIIFqfk6mFlugDLTfZCFpw0g3lUdxuYQkVisPd1Nh53Cj
dELPedniU05QP6BvnrD5oOZguc0nlh5rOjx6EaKzQ+CXmsdE0lJbP0+feEX3+UiiqhMy0fRCB6n4
QJijALsgAqGuvQg2h0oUNLGaJ/hgLptPZJn6u6WESO3YevoHPM8HWXqluDsadgPgzzFycmO+OMVX
rurrwRddI5QJcbut1k15eSC8WWYQBspCpfNWpJWMAfXslmwnX3MsvCCX8R6QkuHAMFQdBKb4BRhH
YdJegs53oGsJaOfdHnID9p5bz8xexh1qLgciopIBpDKRz1B9oOxw6+sh+f2U2rUnLljSN1T4k9DV
AbeYRa08MVECVvxBD/LjNIv1vdjh5XBNeo2/xL2GYdn586HI4z4g/0Zkr3walSq6mwGxKTrY+mMg
eqiY1aELiXfh7Umm2gz2S4ocNxEduk1oezizUlSJtJYeOBm6yB043InQzegYJwQOsFH447pLR+Ux
saB5s/Rm2as/7Kcaxt7Ji83uy5VmZa3EopgkyIJ5NmFQ8vsLluMDOk2Wg4VAT6TwYV/ZksA305Rr
JwOO/dVr6heLDxN3kfo4xsbltXFza3MxIha3TpUhXWGwKpXqdAZ0a/ps79A7MHCWFm3Ulm6eoiSS
lWG8BgRfAV/NLGGpsijGBUaeFaDBt8UqXdwwEOORRZcnXg+AWoAZJPsMPfFutI6qXecOTdgIbCcf
obIxIUrv5sMydcDBfxvhqXu7I9UlFesZcSMG552OmhJ7hQz4sLe1pU2XQgcVz5mDcTjfp/zCWqIw
rasRB8jt3fDVCtC/01paNjIxqkwYrahyfb8pM2niJ5dHqEc8SHd3V7o6ufUhh/8yanfQfaih3sA+
NBzl8mtg9DqGUGe/TXxPMUBZCJdb3fEUYDdKCbdUwy1NKuu0VNIXSLcBY3vY2UZu8AqgDExfU12h
f9oTL7fLgzeM9kfyLYKQKyyKO+KaDDEte0BDkdChYU3zymnUuHG/kJOG8cC7khY2PbQg5DVi+qNP
qbmaF4vAYjiQNoM8ZeKQyEYNk2K/aQV1cNaxjbZqCt7NRzOBswFXAgahgieEFV6PaFhPXmD9kHo8
qkEUtm+4ZS1FFZl/UIfn5wsCWtF9rkqKGttaz7VSnYQO8qzIx5Y4+cHEgqEIqlEeH31KzYuwC/8j
+YsUyj9sNnqgbbfu8EU9+uwsgP8jjNlhMvvu0abKK/ZsAtdLZ7kb5v8hXLvMk3qfvnn3rwWeVBFZ
mlbCqETN4UgWaf8SB5JyTWEAK4z7VdsBpLFa9h/6vTGboYnhPiwFV0wP/HV/JgFsIDNNqZNPaXUY
LrRbl/3pKtc8DKkNZCnOjUTNZzG12rSZQtroeXkQMEAXdQus/67BXexPZ1NzyrH7+1ZdRl7T7P+w
u9goxr6/ioyvUM56ZKZhvJMa+PrOIbJ+nhEzOJMeoNJn3TmhuvWRMi7Zw6iEp5ienCXfeZY9toGY
2wWmXyR68hjFkqsGryxQhil3tAeIleh5BJigss86u6+FK3okxeyZOspbZF0mV2VwSGFoP139BTD7
767Bz3uEeGq57YnxuIA7YjtWQiaQNI1jS3ANhm7J8aHULieSLH8dI1sblK9ShwbSTVBPTH+Vy+xf
tMMPCXu04QUJGaacBbiOkIl6lBgz4cGpAmYADeEbujJ+0fEHGbxLGwpGDSzinIvFhqYETWPbejKW
1GX4N/NdFtteTs0nAM8dsV6fSq6ZdRKCwvh7xfBs/fmOjWS04/xp0Ts/TTlL7U+9d82YDqo7NDsR
uMQYc1JYFR4IcXtRywOSbQBw7Ha+Qfs0UKliwhy25eAU9yJRLp16OA4tjiT0v6ZCGa36UQc1Zp82
WEqG4v3HfMjyxkQgcmB9pyI9pYQqtWs+hwbi4FAA0tA1yzBqATGG8iAOAdQr+44rgnSbGYnuCgkz
uhhduFo442CVEkFbaALL/DN1RsZ4VFTCGeqPvjqhzUcXDqiSk6K6ykalu+VkE4XlCMIFIgHogWtf
Y2Wfk6U1K1CnQqWrziWzFA7av8RscczSrg1DPNT0kkHNVsUXOcp8HSxb97uCizW1Kgn3OnL7SPma
eecyaYRtfibhE2TNs4IIJq1ZExWTxpcDBIEgYei/pl/lkCxTCKYoVOhxlXfqKqvEWW1qIVLa4UGz
Gw9dRUIC0Tn0hLFsFvppp+b7xoCX4PYMircWvLByEdR0ay3FEQGPnY6Q1N8ilo0I0VlyBMWadvOK
hY3T+WnUSBwYM4oywETXmbiNnmnastPAahL4pN4E72MPG/FUIrPHSAL5IZVV6U5zlDF/qQ4nO8SI
QGGdmh2rmIiVZa1/+Xd78e1V1MpeSW3k/vOx/hBBPm/PcurPmV8WSX6M49tSSzRZLmQe5gN7BNYZ
cv9dfPnupVrN2va8YAikkI0OUJJm4WugfWvzwETh231GC+DT9gQVyHL572PdLpgRqbNKue4gwXvA
woVerbFrjpuTyvPYeBuKdvHKNQxRn4hfmIn+BGOD4l/+3G9oqb2ev2cEAHwtGxCFxXaAXA13duvd
ueS79fcBIQQSw6DIZZURfqXnQ40zXFHvvA7JCLgaEfvyjxG6xiME4pwJm91PM/sfDjkg6+k0JMob
RxK2j4TDZGF3YDbsFLADC6NE8c1ChtMgHc2o/Of35fSxEEfdffBS470/Syw4yrP4FQGakeU9YKhZ
oU1v8JT6rcVV3oxhPlpii5DwRuwMhMX3tQ1hOZr0Bc6ZtNLCVf+3IK8+0Mbsmrzwokyrg1xBe4sB
ybXMEHshXn17R9mQdN9y4gHvN5kT98NAkNHmExtPHT5I41ldymuTCk951LqSZYps0nHvsosDRiRq
waYXDTCc4Odjie/ZxrXxBtJhJqTGDBdkXC5UMvAH5/auGM2AXGBXlQNLSOcOZ0m2stEfpV4X5QoD
6RHikvYm3MzXAnsVau+cSqjkDlw65KDmJa91rU+s08wg6kPX4JS22DxSlNIvtTe7ytJVtLB27RYF
F0m/97B9kilDfaNUyowtT0LcdrWLH6/X0h6NCfw+6LNHUiLu/ZY8Xy43TcGfFBMhjzRAjp2q5yEl
yOr/qvT8PqJyhwK1eIBS8qED9U8fyO6hz5s++VAxBPGc8GnQ9CTailsZovz8QcWz3ZbYkuENS6XF
oFPU8CebyKyFdar7CFTbjgvpYH5qg5rkreZ2uf5631CSdgTqn07l+yDaY5D7gHIoqqvz/ZthOmQh
ToboTFYJyz8qV4bGRxDTZq2U3cMXwLpn/bPpX3PZKrXzlXn0X0vsPnPb07WgXmx4AyULf4x7YuV+
KOCi5ouVdubHVJWuQTJCxAF5LmkjKPiGcEjee/xr2Jv9aVs+bndlhLMZhLrLFF+7A08YX2BOQWZN
bEqBxd5oJ2eSvAbHxD/6M/1biRGVWUd1u6RSDuB9sEq5M3CuRTbi3vQhxh8+Zkaaap+mJp6iU6as
Kb+6SAQ97JnyNgG0rBdNWMvPmewccdjpUu4qLHuOl/LmCXbnqESXBG9MIOKGobYP3sQE8GBFeUVA
c9Fkjn8nxJDfOgIkRoIBMfep5LNAzRM9XQzRLgsRy5OnQ8zBtfSFh1Sqt7fy14bLx3KI19de096h
DoBQC97kT1skEfstYYaDz0lPFPwHfU4qePRFDo2EByoxkPl63zW+bSuFHdbCInZ41gSJIKogAqwx
eaIj1jvQTgp+BdUS6H76gFA1bTQPJSOK/mGGqCyGIWteVbKw8dH6NPLvypc366ia3PaXMpc9xlCM
WcwmmYMgrgHKi5+q3kc/gBFrSmYKa74evrj0nRwUBosgTzeFKXGlWwc+w6BP1tcqm3gBT3bavX1J
k7nWVbkOvAxyG0VxVSa6dC+2oSenz6TOKpv1qapde1MIl2EXcX+Cp6PHxasYYOkLLIl6+RnxyMu6
Q8WirBn/txJ6Bd9GXfmXmrvpkLhJ0qSFp/pFDvGPzmOk1SG3Tzb22U0JQGdBIfk9nPr04lAg1zK4
3Ytq4Hsi8uQI/9r08lO0FubKc8txCQc8n8zi02QoFPYmJUBhIcFxL3WUZsC4R85l/RwLIlzjX4vG
5695afCKlK3rhNjnXYiVKOiA4dxY1pCIwvXksjv0+CAC3VD0wqfZUJcm0D00t4/Wq6ntX6GWVUlQ
H1QMoJeEjJ4tcdeg8inPeTyjyKergaFageEEoQf317zAOqzleww1rHiWYNVPm2RS79E3uHviplTI
zs7y+HbfZyXxlL1mHfFFXeRTLZgQpTqk/RPnxdbAZ1NuzPzlppLDuQ/64J5VhVNL8frqywp3RJj+
GlCoBunymk9SiavU0k+mO3cj3xpEYcBPTGdgtoNlF1haA6jrJ/pANzCZG4klsqtUXmdQ7jGgM2cc
y7iJbc5IcLYw6/U1rhE3QxkevqLt11XqSCWfWuDe2ZVadfwRLVK/P3VQgYDZwDKwT8mb03AzN/Ei
Lm/wtphxF4EXKJd22GYnzJupK/X7DiJVHRQm8eaIW6BG1F1aUqyS6gw4r00xZQ/dzNUSSM7wfGBD
jf3DyzZZHKdKlijYzh2YDP8tvag004FHfmyVblwhcSBuJllW2/c/k9ODjPiobD8PtYvfhjQ6Qbr5
yJU4aGft1Q7rRnuGyuk+EREnrXyBTyQcleIKCappGu0TwOUKN/U0RinHlYHvoNQlokgYPFdpTa9N
IeRCgxu18zb7tTthqN3AUn3Voyo+m3+Q6HdxggLrFyojiHWs0xRXAvCMXo3X8BsYAxIWs+2agIXv
VEaB0wqcbKvc8M2ezXIPq0Gh4F2wXWUkBd7q3rgGWZvDu7cVyq5rrL2Oh7ZeZFtI1lfPY3Ybzu9K
GFRi1OhVKgM0NC2Yzo2qikwsnXpp1vQj/63mrSa3UoEypgM/EPqQT9SFJi3xzuUoCivoipbMj6Jp
LncxMX6+bmcsi9h6kH3AxuZk7UCXX4wm8ndJjoZUmkisV7lHLCVXQayGjAZVZv0zVKuWWcmCRPov
EAWfoYAICMB+0xEw/xezfR+n3DDcpA1WbKRqI0AOOVVkSuCn0lAb8NIxykntDxaHi2NMGHHINxzd
HfbjsxuGCJaJeWo4wbFVI9rlM88f467Xk3dshQHA2DKMwhZ7Mtok+3FQXZwrIfDsk04ckumTBwmY
kBrBnRMGMBzxzB9ZDu99aeM40OUdN4xzIYwvrRHLCC9U9tQKOUh4d9vSqA91X5sRurWiPeA0rLb6
NqvxPK+yLUCrm9InZlAT5y1d/gxzGpRn16G+4inoKY+D9/4j/HM/0IaVKPkfr88KOLgM+az4DxXb
J4pE32sDLFvHQozzzj0XnAph7wJmNFEk1OrNZzOoqVUAwUhymxvkfqO+gOZPRJzWezviCrW+b8e4
D3yrmktxaaKIwjZYakKjoguRxEBWFn8JxHvUPOoN9rX19nk8BuR7Jnoz3OarTZI2ROdJdXewc0ba
ReIF0d/csT56lw4kgZvaitxh1Jas0vZOj91tc061MmxegEQBgS/D3zr5JOHRaULNrMRqMBe0CTjh
j9dM/FLdkjPLYftL4OzOr21WXo7iPm7OAfPMaVAWanVrJGblYjCY+20fe5DiJCIkax9paKKqA9+c
VdcdPFOOJv4W0c/GxbZfSckf78lnRCkPVuMZBsdCGpKsixvnDvG6y+aR7Gjqrh/tIK8xuStNf67Z
85CXi22OLFhq8wxscW/TlCy1oCW/LPBsTEYdiyFzCAvdWBFcXmwIOXEpmWrxZCYGk4AJCobQpp2P
IxTOjP0jbGg7B8jfqJOnGnQHffDO7RDEX5ACN3A8owfmTgPseZVDMf/fExpHZXQe3JeGw1AoiJSH
meTdiEs+zHWy+arAQ5Ga2AnA+U5bZT1jWENlI3WbrkcrE0P9OsgatVJ5/TSxaZztF3LAs/eeNHtJ
kX3BGS8j7YCJxn1It1oPhkEWQsNCYH8ifLXwMxakDCFEqg8PQ3NLcHK5s7b1qtSWyd+JXrmXKEBW
qJ3H27amNZ5U6OBcd/3tyEk3PLlq63rc9KML3s2XZD63yTJJ0Ol+RrisxE1P69umr2gQOI0ADASb
ttHwktK+JEP+PIoxD9H+jpMWoAk2dVso23ntJAZ72yiN+n2ei/XZ8EvtLZNmh4UitlwPvGJKU6yi
1atWU0Iu1+e7qvgAxAWsgEqZVDZ6dumNfYGMwOBxWAyeezgpBRn4UdTnEpIVI4TCUmqse9mK69kW
9atkVSXD8rUIauKvBpRw+H+M1b1JktlkTIwbE5efkWsLYmiaDlX1/Tqtss2FVY/NyX5M30R84hCn
BPWGV2Tw0RDlkLloYiOI9GDqrv1f9+z8AhwrREm9aS1FoWbyHUdmuam3z681STPUkr1O8VWNrirs
8CWZoQv56uJK5jALLhU98FZOLbZ8m8W9z9FDGhUrJc3TIegEIkL+17JD4BAi9U6TRLQoRWJ28gDq
rTx8H9peFXBL2Atb10MYKdOZNKVIUYwpkGnd9cgLSDWKal92qGmB5i191W0Ph7sCodex0+jSNzWy
jG4fE5i15v6gTnNhFCvXaVRMi+0zRp7RAErbR4t4f5KhakcqV+P7RFwwCHDKeHU8xlwdRXc+tAta
xnYMlsvbEeviRfaavD6t01mK38NRavVVskRh7j4/z1Oz2xsvdme/OZt4vGVt03n4pneGatn97/oY
GN+pRRtlsZk4I2F86tRntmM9Cjrp9BjpvUQ8Mfl7+aNbupqRz3fdUEaREAZl4UBs9JDctxf1oBf/
Ej+1RXiAY200mT+WtVDqs0i8h0pmkNq6E9EWasLb5kQFJSExZzgZ6gza/llEeZMwiEA+EQeiSe17
bzZVwhYTvk4RmD4oX4nxRw+8mIMxofbtw0Vdx3iudYNfwcCySeH4p5zsWah5rqTMgNNViYjRQR+r
XHZEe/P2umoqRs7fOAyItFWLSJwDA4bFuw5iYAzAMsUalkoRc4eULEhl+rS68aurtkYvc2w2TgTE
KGnH0VDpHRIzUvUiBEA3ttvKCdjqmRNy8FIEtIK88FgS1u1sJI48p93IWgFNJaeWwzxI//gu1fCm
Z3cJL0fk5ubIqvix2lIsYs2vWq37SnY6TsZvD0QizmiE979V0G2LCAE4yIJnFol2kulEcSa3bwOV
rey1HIw6N1JZZCy261qNy59+PidV0EU7kC+MrrQ3U8a2oRmkY1WRNLXicMgmzYSZCDXkbJ7bpZA2
rV9Rj/fBjKUDXEtf/HHgUXQKV8dkeP4TGXXxdv5nf1h6yV97jnFm31iyTztQxkB/yMvJA4d+9CNP
bLgbb9dYeewx8zT2RqAFMA2mzy+dyLO1S5IkL7IicJ8fJOK+2f/vYwyRqdK2ZsGi7z0IWymyTpWP
Sg4GJ/pLKHoPPy1HYQQkG60aK2lnpo4cBj1cGE8gJsTy1LszOp7u1QCTYcoGZstlkX1zEbj3Wr/x
donMCV/WxKlni5yWfs5CEqI8vwXIPWfnlkZwnd0/8LLgXDMG0dgLNV2jPaEw6SB7YVtLUu+A0RWN
vvHEa3exlNhWnu73DIvgbO5ef5PR2Gv4VVGeB/Nz8L9bDaz/2183lCt2ZynkrxsEznSLBVmNzeSC
xKWroVn2mHaP+zhkBdhjvJ89/m/My9EntJ6MsQ4/bCenxEUF2pUznB2cBbEfs8w8MJ6bmvrGo+OH
ouIzwT3VG3zrW15joRQxKFJf76gnrfahH/7TTeYVzILDLcqxyZCjv/qIj3rz+kNgUgG5B+dOkByN
AdraN66m9anENiBUsWDaWNRv2l0bpW2k/ElFCJHHDpU9XlbJI5o0inzk9esyW6sEoGmwW4JH4ZqM
1ylgEEvz59/OSgF8I/QoBx2IokLB/l1pWFYbnciwIrfYTSjKrrEAXSRyyP5Cp7Z4nZRjqu6//fdH
h4ulS5AqJa5lrQVr6FoBM+0DYc7h0PTuJcB3/JnhZKS1/UEtjes+eGAJvv1ob67vYc8NqkreFr4B
F/6eYbrC87bia2SS2znUMmA70l8zptQuh6qBnJ7inhH8FZ/AZZpc9/SOtMDds6QHlkuTbmaAJ0PD
O6Kjwv5xBXuEDk9879+SCNDAkdmgdeKYVIT37U/q3RtYbjmPKslcBsZnDYWqFG9D9afilOAx16xP
s3zAli5pMS9GiFIw+cPQKCDx0uYL6gOezZccHWkSRXa7ete8ckMYAHM9w80BEfwt26cgZZ3Hhj0o
LsmO75WAliLtOwVmVk3GRUzd3IQ70gw/asc2FJXfaSzCLfdEwNFIt0r5edk0sa/JFxYwSJ1+uwvy
fjJTr/+7joEl5q2OML1Hj+Cg6Xe/aphNOLR3Kpnzik0fbBiyDpY2fKkkG+kQlHechxf5HZFyX9xC
ClRGnYwderbyuheQibhuBlgqC6u6L3VA2EAi5iftNV9ObZCMUNGMhdF9027zUcoS2sZ6UIZDLU4I
U4UVV7T8N8/yv9/eU8dNjeq4QBXyFpiMpPZxYSsVSCeplePVzJxZk56SE4NmWA/ACsCPjQt2QqvW
eUKuuLvu6B2982a034MlxHJlx4WCbziYCHVNLFU86dgeo4e00B2/6rS1zDDypeIG4ZdbQ0jIXkyj
R5/xYech5PNfASeVUN9uQggw4IpGnd0Q33cWZsa193GzbxlHaak1RfY9Y/HSwS6codW5dsqz3Ag+
NKNUkN/wSTylwTvMSsYhoPWz34SmqJdgTkpXOoljahUShV9HzuPqVDqdpVosdezjrKX3FweM83dn
dQJl69oEhWMNSyuxsQhcAF15XvHFc9M65PyG2bjK61bLav6OPK3azByHwuQUIvexQ7uktMPsdSb9
4g6uvifhcU2FeElzQOlP8cIVaYMgEaVU1mVx9fdHfQkbyxHR8T28JUDfJmaKh+8HO3DwmsZI4KIU
njZkKvhvmxkh/2+79VK30VcLm2nn+t5HFfDDo4h/2tfBCHHOv2qnuArAQvNq+UHv3BLry783O/7a
JADn624XYhCSHFrBjj3djOxtwD8t4RbkLtjzSF3ijqScluOgk7vhhvTEGobC+nBLtlMP32g5bhmN
OeNHjMx/iGsbj0nvxfms0pcZLeNeS07Kzf67b22khgkphI9BukEjWjeAAJaxiqs9YNbXnVU/w78W
5uKnjm6u3Jt52mXUN8MeDZS00yvL/H8hxcC3/5CmJfRnPZ3xWhdZJxJyN7NsXCVRjZBnJI60ftwL
2cKSk8FpyW8ifVO5sY2PNvIJEeNRQMzqmvXsMKvfTA01cRIduXA3NVL+dieNlDF9UL44KV6VfmN5
MnDG5f+YbiqEdIVPslVXENUmV4AHS5QiyB8bXhdSyeSPDfBrFfNBf6bItWUbMfoF7/f5d9Qb3M2f
YyeZ8XKRIUg+98pCyLnhGw3vnWs+aK4oArCDrA0xNk1zCwUm3pZ1O6VoPNlXAqMcbigJjwpLqGF+
OnrBJ/8enNGeg0zszK33uPpZ0uW5HuXBgXiztHG0GU3NeZ05OoICPqepZZIGdK6DhkTQva2Zpe2u
vUXlpOsgWUkUPv/2/t5smI3c5BJRF3UGFmdSdxT2FwHLuD5knuvY29oPKk7qWhpq9BFHEuclmnck
xK1ld4s1x4APqpTCC3MuHV26+ok+eQEWWht6dOpnyiQ32qRt6wlFLwYBG8sb4WmKLAjdLPOgU3bM
KnDP2oX8rvOWhr1w8zBqEoJ2kLjZTbNhU7RPSIjCmM2LMkd1mH3DpGGOcufYz9yMbchlANz/2CM1
82yeIpALmBxmujphmrvECDMZ1ASxXEoaTzHUDjEyLsF6IrDjo8WAhlQaXLte8rI7Zk3RbcN2Hdj0
BUaxAHXdXPK5URzBZyEAD6hvo6ndnnLtbeRjQM4OrmmPP0fiRumvGz9EG7KJCcFlxdXJBVTZ6N8d
WmJFcctKLmWRyhEiyq4BZCtxd/rNG5L4YJ0LKFUheWAov3Avlv/lQdw8zWRPgxjupHXX1EpMUXv9
RfrsTaQqTWfx4+9gXIe2uL/tSY+N/pwOcXc/mJe1iQzEiAywBU6WHygnBY3J6PVj/DOAEETmB7K3
SSvoCJQKf/FXYyoD18TmEkeqeQim/yflwy5em7R2CdII2BRQjp7PX6PAe9v6q6Pb1iJAitfA/gfh
+BOnHXlHX2Ln2esV5ZVLfz8EtljJKI9pM7o8WRjKB1PJc4vCPoAvQ8UWPxj8xrfAgrRgorYe7ww/
C1q1Rc0RjNmVDgxyTCaQ3BWUqnrEYqnSvE8WTSsi1jVj8TF3wpeKWi62YhIxY/06sevpFrIq/dw+
nTzOMi++3NYjot+ZW1tkgxlBxVMUS2Vh+391xkmN3pwrTMufSvikLpe5rw7YQxJT1T5fp/dL776/
+Q3XNU8hfDYRPxO+oTKiDFXYxQkve6JfGDd+sQiidjMTfzTSiebk1kRRq9Tak0eXSZXkztET+MTT
7E+eunHM7EiLwAhL+QhwcbpsJEXfGpXWrmUk37vj4yycKuAsmcJfDvp2arASa8nj1MzehLcC/43z
vyUT1k6VEvB7Xb66SsdoLnMWxgfvXlrhu0oez2YlyCzYRviYTpRnDQdJ78KhQpqv6G+dlrFtAbd1
diA26nbyk6kPLj0ox2KIGWoiiUf6znqE975DLxTDUeKLrOwNU33moKNj3enNVBM3CjxrUCLqrGF0
QQ+xs0DKlD+zNPD/QoU3wvlVpGWJieyGF9EcgK4jEpjUqcvNGFBDbIcrSU3E2oEw8wqQyFdQjMDL
wl+rQ4TMUzX6vmWigdhAhQ0O9bhso3yVNSEarq3IEXAX3zfIjMiJ+xOF1CanduZ3kgnYRvJOyapw
TMg0r7DcGMUhj9OwVAJzcCS1RmRk9vsSD7rIYGeJWTqtNkGBZZYmc0iMH1yNtvTlw1m7wEXtnpA1
nAg1p5khI+HCqfk6c675XcrYO9b8XDpK/0H32/4IMr/gBBT5Gi1PDnG5Tw3GLY71dhPq24eJrv3C
Ptr9ml9HFlMZDrUU6LsllDIxk9MozDikUmobPUfR/JqlUqg33kltdf0RE9bPHDLg13/tlU2aY0aq
GPUzr9CN/4CmE5ZuCm+tII+qhtWxKQoJ4hqglWRqCoLju8QdcEnVzoPHv8EzamSoQfsLoic4pJ5m
y1CKLkQmebM9f/yZfTMOTGzsH2J9fZCIoxMTOwE5R3/racKpg1VWJ44INW3FxmAfdAcL0ApkTZhA
CDBXOsPqv5BLHt6wyvv7Iew5ozYjXhPNlmO5dbn/udQgUGYkgUrZgDoXp0rlPzBELZyrg1jJiFtH
d6S4Ue6VLsy7qoxFQdYSdLqDnF9auAD2tFiqSz9tN7WGhfIYCol51IGpxFk9V+tsXm049ThG2ms2
y7KN8DdKIvu14xxHD03fofHPSY5kzUJ2e8aGpMJugFlj0E/oVCAY9Mj89pBNu+OC64W7bcg4YpVr
WmcuT602VeS8e7sfjakpefiJ2B8z9hmmpgcN20sRUupEyEh5O8zgJneykij1idLdlOrYyDKRROO8
yyA6Q9/V+u84ixseIT90EqPXKG4r3W6fwamS3EKAbpvky0oAq3tBiSdKYin00fxtcvFxYJDQkUfK
ZucR7m9pvlTGjer0XL1q8vkbNH9xN2nBGmrL758iTmp+G+qYa+mFLLm2Yx7Z+k9QJhoLrQPVuOEG
UV4s6Jn8UyINF1l9S0zXu5SK545puRm0qzA97xZRT/TFsjwjaITCnPaFEF6Voqw5kY50eDTi5vmy
jEo6w99HlNWZoPZ9C/e3iYRMg4c5KWZHUpYg5b7/uDJ5dtJdTATdOkoMRWzUnKO53hHR9Ro08ANg
zb/sjwoscBXEREJss5uNPYZ96N4jvhqcv6Ch30vqMgYdQ77I9CQ9TQOyr0M5shM3TaWsjDFIOTE9
8AO0b+OwzDu5xFtNSV+bsJz0Ja2xTG6dgwMz7M83bMZ9/J0he/iPheLJ6eZr5/F8FCG8wdwY57le
HfnFc7wRBSQLQNzeqIDF/0F2uOTtJp9sIJdB7LbCdGDxE2bSa61FL+kxkGY7jK/G/R/xsK0tP5Mz
tYSWcnHtxpR3Ij8aDSGMm252i16VXFnBEj218HOpHN6UAgiU3D7VN+DkJcIg4z9D+GRigxu3yBxK
9NDIJ9q+nvye9ph2PwflD1Lzbfm1uRYKgGw3Avd9wzXm0JYwtMIAhygTSvGfzuqTO4WUXUDSuAYj
9TKuRCOAy07yOsXH58Z6VDj+iul8aSgKOY1APjUqKLFKKQRlcdOvdpmqTI1/weoT5quPkOdqNwSe
a3HowJDmbri+7n5TJe7DUu3rCc7lcRbZ/X6UPx9Wo4zcIo/qSl2r0+ag+gKzmNfzV+sec83CydkS
pXgXpZCrGcxynWwuJmwvhKuUxWtPAtubp/SQfXo0qKns4nPRyfkNIruHIoTFGZuewAgeAHtL7Not
/YchfZptxUo8RILSa83+TGqbXLbZCW9wV5Bvo9pqZQrQgoiE5AJKOaAvnzWnBKx0nRFajyJEdBbw
C52NPGhrd9NiVjUKs9i9QcyQDvfhZxvYOzRAX1W5DUQ5pZsdVSYO8UnxRiYdc7d7+1cxZbg5optS
0azr7NqhkRoEOtYoDE4Qhm+Wq4E9tW0OfZRMLbmLUoJOvO+oriey0O0igYUKouKHJwwdRZgJub4g
OetI2QsOMsWjRZXcwqmP/pc++94/3/BHuRgtGKK/55HRQQfPyOg0D/Mdj/eOqlU+hG5fSqjisfXS
4p4QFt9lvTeFzzO5m6wKvw0E3GE6ts2n/ofpAgzjmw+XI9NlXHDfuJmOPyI75fjF5s6BV2T+x5wO
0M0YnTbNcd3ChA9NHdIhdK/noUi3MDh+Gs8TvvaWDujhEoLGa/Q2lmJsnE4L8mt28XjOXn0pyemM
G75RKXLIQ+/oxkpOgPKrZ+2JfWzJnJyd+EGucmfadH59mZslq85cU8ZYdKsa6o7uQkrUpZwO/vfs
1G6EVl0nWxrA6wg9bl5N3cvZs+68Z5J/lcYPaA0e/E3FNcdWgTsoq9+mVf2eO66inZx+sEjV7xtr
5HBluoqlNfZjduwwFeAg+ebho3BUhToplhpg4Ti0uKDGSmNORnGf9vnNF5N7CuN+PNdeLr6Zm0bE
Xk7Sx1wRRhbhDJ5d73hRWSWOJp1LpM1jlM5PsBSwZxKqQyyasnbct22g40a7sWeiwKPXrpiqHO8E
EYdRLJ2VN0eslV8jbsU3RcCCrY0KcKu1Sj7ZkihOvY/AuPvd1cG0IhqthbcxWcB2tzCZ5cV5BJrX
tduEH8x58R1Um+syq14jpoFCNf6hF5LBcRx1VI4gr2PyLSy9GDDteXFQvhK117qYrT20T0xKUgNY
c+fB9prtRA46uAR/oLTAN4XHYRGxMLPaafps9VqIyf0P3kOx3gOLLOIa6tf4cANA/rexSY+chDr3
f1MvIEWV7FBhsX7LSUk/fMQWUBZe9JjZASrQH6TZe9mmIh/YWEA9unWdqga3ZNme5nengnLVDtxG
roly7+Oh2fYjPi4R5Qop8hM+lGCJOs4eP6d9x5u1KA0UK84nOGMveMqbHi36+yz0o8Hh9pfgThvm
sqpEt+LqkcIBjxgtDYKJH2vk5rm1ZyRqwlw/HCUA1Okp3CJIskMvyftvlXjyeKdx3LwfGM57DdzG
M0O72B/PMqqpm08KJPZa0C20w5tGdx5OvaVZlRRJnT7U6vbFJHbjgSiR3+yAy78rpI8GQPP68Q3u
u5wCIqJ47d03cDVddEKKCUNy1CU4UdEGSlTvwYRgZzP8Py/wHq2OFOkRP93Oqy/wSkn9QI7gHXHj
xhPiQcj9wVnu6qUGWWL3Sw6HBC0G073hhWrX7Mf6fpUCEZtXHWSIxWAPnpEdUQo3WytP6reuoB9N
7J918NqwfZ2eSF2zO24gGcsefnMIJQ4fTQwRB2if6rIGTBY9TvpmqSPlC5rMl5UBjZPuWBYm+JDp
0eNOKmQrFAcRTyY77RHwufi74cL26lR4rCCfmNmRidWOP3LbdezJnoEaD8LHswn23FsSjMzDu4oq
dUnYxGUIX6yKUH9ZiK44BU44UYE1tzeHzrvLgJOSsx1kPBL0NiOIIAkJjAYyYrhqekX0OY/WbAgr
PomCS3c/yy6VsXxPe0CpKkJVWSam0VJI2+ZV+Mp4ta6MEju9iUEIlAYL4xy+AqPJm6gLp8YPmISa
k7loLLp7VXybvbHVruQPkje9R/ILf5twk1bkgQnlfwogCQlX/24hGGHGUrDy/TOBp8PE85WjMuws
6skEIurI4lldB/G5S52rdrwGDqDvoXV8mLEqCsO8Je4wAN631aaH+b/3dWlAy58CMH3Nwglz+0i4
pzYHy3bRMEOXSflXB1MGU3sKhAKRHevayDPwlD3b0+X52L3uDWTScs4ERYeUBrlIls7iG2NkjeRQ
477m4r3/vo0QDI5svfsbxg47Fr2QmEAk/w7TqUHgp6N1pcyp48B/0thXeSxPmAE+paf+6UZwtAF9
Sr0dZ6pE5L8ULzLNzwaesEV8YVjyVRBNwanhAfdHpiZaJX9fGQHytbVtrXink5OuUF8Vjprqo8PX
xAjqTpWTch3YZb8shWy61F9uw92a3S/xif/P0NUiDaFqJycD16s5IEMLE7cTef2oWh0QPiLtGRlf
z6YAHn834iRtArDRd1d2gaiulpNcaG7uY3t++fyEmqg6e5DtXEam4d+N25cvyobwFu48U6XUP80a
quGMRfOZ2Dw1AX1ERWP72diL3nG72lDx7Sb9ymNdswrjCsTyRg5K+dzD2iq5+lYl9OgV5zhRvU7D
sjhiUE0CX2S4sA9Fiu1he9pa/4sjmuKtO9dbjH0TM3eahLOIrpEMcrw9bZNX4sYdKSz1k04U9hZb
uDiYljP5BJVCQXIiPPlTHmCgIeb0tU5/d/6kk22inPTTMIbp800/afJEios21sG5QFuRuAUTdFF6
2qYT9rrCY38f1p/wtsfPgy7QEpUVAATHi+xqGYuljdqAj3NMdBO6xv0ei4pZ1zqRe8mBk9XlXdKd
tApGob6l8waorwwql2mgHN7NQHIQY2RNZsYJNvnn5mI+MVs5tNoFcX8A0EfY4AjvLgKcXl5/yjCt
BobMMRrWu6HWPeW0XN0jFG4Prx9Sx/S8n3BU8VXgawrayEpJk9+OLsmnE2U526U562objKwR2C12
9HBjNoD4AHbwGyfRuVvPNqhtxXwVPaDwpn+DWD6Ac1OSTGU82wNnvr58V76ajXRl4wkIGqF/2G1x
pgD7yMwye6zK8SP93N9M7Jlf2jpxQzomRkfbWk5ZxF1G+z55ydo/XyuK4XIwbxKcCd6cdPnMslru
jBD1cFjT28EBpqaoCgcVEqxVnHpeOt5UdBoGMqsoJc/9wiI/y70SqLvRJvZe4ycq32Bo+6VfEoCv
MRcPbuFdVKXot+jlxsYlJP82c1i8AGv7ZEg5O4oyjdx+qjfpYw4ac1HkOZXwpzdzz5F28TJZxmlA
pb7uat3wVer6vdRVvylN8TNa+Vn9JdHWfEdFFm1q5oHJf6wg2U7/x6Gz+JIZXbIH5aLyB++GHe3F
6htLKYLieLtbn/K6iasZ7YmwRaC558JqdLNYZTNAsXHD5pY6c6Kri1/LH/nyXQ7DmWbaqgFyv+lX
b4o0B1gwQ7ccs/PsKVi8Zri7/ljS3yyQb8bfBvGBh8E92N+j6X47Pu6KOSLnC1LV3i62yQD/meXk
P3OrZTSAgiSkp9lRGTIEiNhkFuJgPFqxA5hUNxRrSzilplcXJ8H7X+v+OcslLwG0igZJfWiLHfck
enH2vMziZxWWTr/BYBedjHIclTOqDIUgSHkBKZ21R4H8zqrk/vpF7/c/O+biXSlLks4jw2rhV73J
FyzcdO7zrBYMtLBhtIhdhzvzfnO50XggbRNYBRhWLwIqBkxkmU0p0sDZF+h7clF2JkcI5uENdFEx
E94p5muVNqrhRj9GOew2K4tzmelLhZarEzqzRwZb72OpBK2NnpiZW2v7aczG4Lf4sl/nKAxX4V8M
AsJrT/QVehehokxUESlVzsdC45v6kUmOJ1ZxmTEkR2kHCK8OddLrUDOyDp0YB7Z2OG96/CTvBCgR
e87dIySouYkp2cgeI5f8mfT/ajo/IfJ079eIs8ByY4lcxHLdpKM7G/zrCmYQyx84j6ywRi3efU8Q
ZHhz2b9PHRvWcp2vEj9vSi5Qp+2576YKbPMANwC3a6h50XpcK5WetbdyGacIcaSs9yfYJkDISr2b
+VOnayPH03uhjMHgDHUMKezm0ZsPx7IfQHBd88BwpPPCnkwL0xU3lACZC3IhC2MqimN4Gk6g0dB5
IvTCiOgsNV2kMINcl18T8JNkSN4O8haDPJKDjpiW5HyRUaAE/g+fIrRagPgxCYQr7O9i+A/WdY1W
DI1KgtYx7bDgiRTLCpeJlPwNnN8A/xvG5UQCZAET2lBZOVQlJpha5VBszZ7bqKoDEnTtJ1Q29b+m
k/WxH7w/Ys0pKGZYULFKTmsMyIamg5AvlBQNdyYL0rv+fQEvDyBJpo/zGyXV4YG3jftunn1AlH0i
kOwdCsBfhDvY/4o155mJjZjLNeLnTrWcC1ugctSqWqkTDwAR0Vq88Zz4hiGc+MWGMBX7+HYBMNbo
85N830J9KJmWZEa3qVBKklxlWgsWNtodSESfsY83TgwG9lcDRYFx0vtzy3xzCbXwmILiOhldlxMp
NHn+UVIpXDO02NKP0uho5XdVd9pjXE9yMl30oSfIexruOKwKk3gt+sSrFkUuBmFdODwmb2vkBsmC
yAOAFcm70l2TRL1BhQRxnBG0D9KOP4AnJSJUUQjcz4jQd2qqmJJ/Th/hH6HgNpN8nWd1m6syUaRQ
9W3lrJCZuUBv0mI9mmSNFsSVUwzGXVT6/wWgPALAntOxw3wKUE+mPsVdX7WFbaO0A0JViwvv8tXq
8Ggq0/gvZVUZ77QbIcixHanhO03VAi/edZEnQoj3myHZ/mWEnuj0D1B5Jbl8Tz7FLSiOvF6b8iIC
Bw9GBau39eefASxvBAWxLlUzJ144HTeg21s1+EaeQ+UnKD0flhWH4kfaC9Oqy6UqC11S5GZnbVWZ
orC0DzI8Yy5C5KrRDAv8AJxtffSo3Kahfbiem7OHnCYwznRT5lje9deYDtaytZHs3D0CcKDN9v22
5TxIP6Cx3PBRTAp9PP3YyREHen26WEaYhXrFwqIRWWZw6fdiduGZNBAhpgoArazCuE68Fo6GNmFM
v5UEbjJsK64pcpvJaPdtpp/aTU04TZe3YYZ35JZKrOqqOH5TuRnbwZO7GcMruiODrBr4qAwWRgMw
CkkiY2IjLaxcZcIGX+yMo1lrMEweAlRwQ1nid0ugh3UmWev9mDpHpXIbbZqrKeUfvcQPbilFFfpU
l4Ai40kEWfsdKCk2uPMp0Ceb/Y3zQrsYc18PmN1Irp3WDPqecoFwxZVUrgK8jGdxjMrtUVxu05zM
7XtJibYomwbAt9FnWvZwL9bbBs2sqDTueSZ+B3VSLn1nN8r5lW7X7pet1W6LieWD8ZtrN+eMWBNi
fDZM50mshjyv/6k/0EgTCY4JzUjVDhYax1L7K5lkHJ5rQaTvBrIN/mp6/dtyiKMOxudrtxTAV3xw
cxqXzt2kuzPzWJYWCckYmuSzyuJdbsPo20pMh0hceU5gv7TRw1yTZ/W+sCd1dnFU1BDXkUnfloT7
0VpLH5usomyWB7Q2pzUsBvM37oOHFWgj7NRTai54WPRztf8okB+o+1rwG7wznI9uDXLVjXG/sO3t
ssB+AF1WVfeBtRyGVERCkIgUm5sgYfpo4utUN9hxSVp/7R1VVsrYi4H55fIloGzDLB66+pHfoqHd
GXOZLcRGo+8C6rwid57AU9TQpPCkTewE9vpskaFKAAzWHnWOynZcTV9qdXR9PD2YsCoNu4kWDJce
hY2boh7iXjrkGZmctGjdACEGeRJGwAcjn2+Dt6wV4WkPX3lxO2gNTnUrt3zxd3hJ9dGEWQLfEQEC
giAjUyATwbmJM03h2eDV8m/d0E77G3K2ZWVZ37Y5CyBSui1fmGWKR9US9I20UY7RiyS/U1Xplprf
jl6dX9RrazUoMRsPtnWQRtwLuLhmQRU+kTe51FcM7wyZfs8QTUnt9LdGizWRwSv5ZqJPApzIpRYC
fOHx68s+JKHlLAlfGsC6CSNNHHp+5XsiijTwo2ZDKj5/PGfDskXtcXh2N6oGhk7zDd252y7jIO3Y
JOhQZ+5YtEOKgucbvTa6oCavlI592sNqczE8rfhzi4RmvAfD/K3Z9SjOXb7XzP49a2AyysEPZ6jR
GnpVcxPaFqgHLNDS+f8Mz8pFYhJsRq8YwhOONTJLdjeQdw897iZ3WcNimr2uhVmzg8DLese/NQGk
1BbZ9iDjIoVnGLmOY/PWhTKrwNVZlbGNMXRX9/27S2+M1p59fSVmV1TUNQVfCINCYI11zD9hrt51
5XO08HABAA+X5GG29Djqw0TaTamqOpj0whddI4v3+6fQDqUEHGoI9rW7C8EQrBfUynT0AQI2SkYe
o8SpnkaQhd9ALCJSTEk3gBlwtn/t9Y99PclT1fQB/ffaGGo8hr91jbgvbuHT9nf+23abotW2LujH
Zgk5cqJDUB+q/N9LRsm3A7e9Do4bsrdBzwzTJidtJGsinVYU+k/9GIk9tzoUFXCzTwP1GuR+p9Ft
cWWbQqjdADnWJXryy1zIHBaYPvNW4KRbW6Aj3CbbxBV6Q2Wc6pRMXcOfLZnbjgWfxn4XNpuL44OJ
WjTnUTogB6Fd2RUkqHKYdf23jqW4GOiax+3yW/nPJ40mnTIHGk2So4L8ml/k1xmpTEYIhummeT+x
wrvKwAkiJ0aA/cLsvAvZKmiZ1rdA6XZC8JmPMzU3xq4wZ/4zjujNW529KwSACKNR051iREfS3vHV
ileTIiLL1xl3/aq69lcyPAFr1X09bt0GIzOUHNueDaHEIpU2YcF5dONupmIPodHU5BlWoU8xjXkD
0n3rqSR0jb+9pI2Ii3D0lkoya2oTGbWWLI1fXd9D7Bj5pps6obUP4zzNxos2f4km+G4sqFJBnmyK
MPy8Pdh84ZdTKTIQ/SYuKofZ4wmNsFkzF76qo60jGSsYCKgG17jtnNT0U63gOrQiUJdt/bn1H7TE
LWHi++aNHZBILyqD3V5jtfjBzi8qjgHWC5/RkfFE4YzJhcxnxkuzH9SDE7i4kBqQ4dnShFoZNRyG
jVynYbcJW1VNyisu8stRZY12S9uP3pgzFJvRaE14FUljfFEX0ELBDVZeHziAu+jnIvdb38Efn4/7
IR4s84JoN1+hIjRV0auFTkyBD41kBf/SrK/Ht6VhBFTd6OwlKt7KU4rMmyxamI+54ZjP32ovHKRj
ndNAtALbgCgzzT982TKikFvdhbguBF6oo2OUUZ61pKRyHOAsEG/A0yiiE2Eal/g/HvsPZWD/Rmu8
cz61+24p8f/WOYgqTnSsPars6bEC92IqaryMp25vmtepTydieh0w+RT0Zyr/Rz9A0odrpwTwkKie
/tVZnycL2AwynzU2pxxc9Qsx6Sw6fZquEBDVrpTf54O84MkEMPPZ+JGtbj5mkLQo2+TLRRUaiH1M
p1LoJwlJFS1sR7UqTHWkNTc+oHZ5EmSCWwIcpsCC2f7R/BCA/ItBaV2sTnvj+ncMUN9dJWTEwfVd
vmPtfmHM4HKHrtb5kPsfr0AZoMdHAvsq/7uYszAxqFTcnOxeC33GkY/F70M+G0Og3qaxUEWcx3a/
Mdf+VoG3Pap0guTH/X4VJHh5GXW5NKH06IUHaYByWpYQ9zLrFaAYgRR07Ksd+yyfbTGOtqvU3tpq
juctZ/ecc/cly1WI+NIXUxjk7Bc2ZFUzvLTaglO+RPDax5UGJr1gh1W7heucRaXhmUjhCgfWGiMH
gFnFUVvlvddBMqd2sB3DjpVDD0Pc+mMQ8JGOvEvtbVg5xXIwbo6wPuLc3JC6mitWw58cAzqBp0fP
zK2aXbbhDAXm11ZNYQMnLaNjXiNNgyDvppAYAUxrpGxdiJFdXmusXgzR1b1zQrsEMKHG0oLk0ZtG
nan2PIudxGlR+QsGXma7+EQvhNjqqtYhR8kjC2be98LRXttaVICVIocxZQVCWDowBKxQRXkuQnPU
Thkgoh69NylKiRqKlcgBtZBCfUcR7lkX69hOSdj6jrRfyJ16JmGTBKIgbeE0NMaXpvCxtN5GK60/
FPXlQNkPrEA9Pf+X/56dPRRX3PIQrX7eJaBqYQAgJFg+mSg2I8UcbSE2o5SZyumEwieImNrPpgNx
ZalJHnPGgdpqt5a1qvOYjvRuorlCerexAnoIg4dwCIV36NrhVhV4XaO1ugthjg9CecDMMjIkEK/+
H7cYsiQHGc8UQmzwpFrFGJK6XVCrHlprlhCErBcDwLQ76h+uhL8UdpsDkZkNh0v87qudgTNKdmZn
EXeyLfVyVI436cPWjYAHvl65ee+mDg0nPw22HOgB+eu1bOESoFV9Jq0zUEWC+y+KEc16mfFPP81X
VeXDU2OXfDBnzCBUk978UsyerT1zwCyJk2jlhxj8B8vs2cRS3iHNghyrI2IM5OccnohlBlCRaxUu
2iNcGFqvMPRYBLk0YB8sq6coYdlUFs5RArdPQtecXCXCrNSFUyLKVLwKRz67KOdrYOn1jAvifOG/
YNmB4txWdyvmLXiaWg13pS4bknlnMD8Gpxhlc86aVzyMhi0bejSrswWpU+Rrzsj3MX2bMF/7H3KL
q1/w3tqwG1nRFgFiL+yTdipMe6BMoTGTn539jVIh6tnVSYLTlmfOWAzI538HImMs4jJtTaXra36P
tOM2pwBu18NHkqS31P3a7MOfIiBsQwQggXGTB1c2pv0pyM/Vd0ektCIx6pmP0hF1Dla/13QRZqX1
MC+MBPb1YGeFxNdmhJV3owToZOXyd1ZjTnAiGT+cPqOC/6Q/TNRSTumSkXue5MRCamRNat4wgaOR
vy/fZwB7YSTXUlNScl1BNP8ehlJ22w7jcnXt8xJAfQinUcheKnpfEkdl3KAR8FX/+eCV2t4psQmg
GO+/0L1qyAgkZ6k9ZMDbSm7fkV4idnJJfJ6StdY2+TcJdy2MvoK1QfD0uLct9wBxmKPqHI4t750h
A/k6A5V9Qgip4rsVy+0EzlF9iEHZxlTE85zxX0Nm3RZ9uNSQTAVpw12lHudUte19trpVuB96QJUZ
CUgqIsaORpnoqdHc+XKMlMZOJapM7QL7uTTXXCN9lgBvoa63ARpZCJDMCQLaYrqfmr9/WPF5r4vS
Y+ddqtr3L6sk5xaiqe1puDTkZivt4kl+cfdgmvx2Q0kn1FROSYkfIcTk8pDJMmLERB8fdEerEcH9
1X6xYV1a2yZMjCzHI/qrPJ09YbqMjfJaScf3isvH39oqCtSEWm1R71N5PIjZ2GEtMfxOr0BCgEYY
F/sGGrn7Muttu/NDLSkyRAzUpVaX7rHC9J0zgnIMorVh3CHzlf1wGst9kCM9vLGMIzzwFQey8UC2
8KiHDgDSWKy45vrY/BMAY8hD7TT/vyN7Q6YsnTLVZ9+a/1oq7SPkoXEgxX4JOPeX7K5rEqXhUqy6
RkNWAk0biaPbo6GSCWZ5ZngXjZ2IUzewQAg1F0ZeK+a1gu9iC3IZGUNNIw2N/w7x793+A7SKGdSZ
fjkdui/AJFiXczlF/Kb50tLQGJwprnkjgH1anaI8V/qYi5nvgcprpMkEuVywpc7iZw8r5DKz+zps
keuPh3Z5SxXsCOiPUK8of1SOphdEwnTRy99FrIGcc26sILLZf7nbHmi/4RHEyaka/FtUyT7RtX9V
l8YWHUlMFWO/oP2QWcm9oFiiY0B5Do1RYK3cwGfOARYUu7AvuUYxYGNlDbqXndvtmq6VYCtwwJHs
bdF7qiA+cQ2Twx1rtxjlIqKRlE1OFA/uro/iabgonIXO9ZQGyc+UlNvzGj94CeANjT2qrGuLm15z
zj14ob8G3rL5Qgk9e++cew5iR5pJbvV39u9GSeKs62TUXCNXcCxrzaqX9K6g9sBf2hCSNVonsSId
pY/eX0uPgcCyie/xFN/77WIKIpkWpAp9DXW7XsQLN+BxKc+PfvCOimOiErurwdlqM8ZE2W6v0jEJ
4mn6eg/or7jskG1fVAbsx6AmR+cEKUtTk2L1ECdHSGGXBmrjapYHhIbC3QKZEOLl91QgTY/nAyhO
kOeN1lxTkXeKJGQ7mFaGcskP6JcNHi8u6WjzkidjISslsnB9gH+oz2I0TQTNOQ6IHrIecigMu0ly
N01xdTP1J+HulsbhycWTvZfewnepelA0Fn8YqvNccpPsGnKBB7MTPPNZR5MBafCxqxptV8qJmMUJ
VXXO8bC6RJTfZeo4m/OybBCa77aPOQGI/Nyjh9jcMQS7KxdnwNY8bR/A6T/xfYK6AIdg5ue7CUdX
daVSNWv1bk7Cihm+7UTtijyVY7vozZwmIw9XpQCqQaLXINDU2f23KTTXLr3Sk3A8dYwamq6gAUeJ
5/Sr+eAevJGdMSgYGwYKEF1swWs1D4GgLyICCckpMybmXvWe+5Q18NQpQRJLyNu0of3nXrtgx7Dy
eMLjkKaefnuxGF5RDrjb9cTewIz2alPVBJe98rRPFBpMsNSN/mQrSCKpaQwZmcfVtrxdlq5HJfXa
83xgTiBSVvxwSl/l+5P7MhXXmWFUQJXioSWfAzQlK6dAg4y+UZz/wIBICEFcpbaH2CPUEph0S5YX
KGzbYLWa2fMjB9pN7Tf6Mykl78bCAUe1teS6tiIfDKO5QnRGhbm0I2ypsEBvCXjB5HsKTu4ukcjS
zHQuFGkUvzHIL6TIMxpPx9Iovtwt9z4wzXdByRde+tC+gKWj5ZraYKE0RE7jPXVdRiSPgZCBsOA2
DwlOHkdRqGNpiWfeKBaLXAYIVVWT94vrAZ12XwXmX/+CQYBM4zzNMSBWZ6NMw/XZQnnTmNe3J0wd
f7lOgWWWRRKRL3rZ+jNfmP6PK5ZLo1N7lgBmHgdOweJb77Be+2jZjLqjJO2ZdLTicaQfwVCMZfHV
DZmDz8SkRjzxBTfYK1irNurTU7+Wq+RDpQoSBJQWumC1rHDszo9SqPCTXRjkmQoVjZN7Ym0sUEMC
/yDH4tjTM7PjAm5qqoyrEktY9JOuCku11T/3BRKJDL4sVaFSffVj0VmklVXWWI4fOJLxDtVHKo3o
hoARb7tRaSi/z1Ny5QvPdPcD8usOUKUbyXq/QC1OoN4x69kTp2jM8Qm6T/RtQvzBAMcpBoxu5EcD
I/f2nW5IROkQsWjOVOchi7reYVoftKHhb+ZkCmJzbY7erDST1Q47cHANKrJTjHXxDsBZXSB5ab+r
dXTZRCOUoy6IfEgA7BexsjHw88NOYK8YFXlAhy2NP7lweJchS0lt+Fubgtm27uS7Xra4XBjZKn5V
NxrQa7oMlYhZ2fKnr8wkY8OLNYYLj0+XsubODd9Jwl/xh+MKyJtYwaPRmQrie5AilfK0nJ9mv3gx
TH5P9PDTv5D0Vd55MsoJQ5K4U5w/NS/fvq41eF6R66fiXihmNXXVyxtCx05FEgzZcj0RuGMwM9mt
LgH+A2SgMojLwwtOLs9pnn2Ga3m+6J/OxxveUEFwolBFy0S290oebpHL/tJY8XgDWRXIbUo+UUES
udxYyRcOD5PbdBRrQQFbIYCmDF6E5QyD9IxfAB4D7tNsb3bHIs/7ju2vNhwcA7de8C5Eezwsw+t5
JFq1WPShUkl8u6JnNRkCTqTYRYAKMLTQqkxKVVejk4v0sxq/n1g5Lyt2r943oTbXZsKD68pga0e8
Iyu9Lv4nK9mEfJTm2QWtDCDVsRX++C0bNNf4n/NlSAvq39zjCAR9BA38Shwrcrb1EEpai3scvfhh
MdZWKRHTYXtR4EFNW/N0zs3ieBl7KET0OYyuqIvuga1fIvqfoUsWkTlPGO4UdaUOZFj6VH2e1aww
F8DWgPS/FVL2D0s4jbH7TKhOhmtXVkAHMXCe8BMLPRVuteU7hGOdzJj5pDRybU9kGZiN5yEjxdAT
Yy88U7VpAoCKkH5G/QIvPinWxB4UTA+qY20WrkfWb26VTfqEFZ1eh7RuXQ20pHN2E4p0akNARI5w
Y8PUItbuOmVcije07WM+xAXqxUs6y8V2cIJCApY+fiwOmXl5kHlVu7ByaRuDNn/scAUfRUPneW9N
8IGov5/G/RTZk9sThDlecL8pPipw+vBxXFF52ual25dnCJdbk2x3kXnuoEsN/AHh6DaOaFajKMm7
OJ4eSBe9EgpWwQK8hT4hQc2xlOgXxgMHGOH94cRyXtbqUZf/a395DJYKusDNMPRaJbr/4upuY9kw
FnHIWcaAEEMFVqSSkUj6EQZihloPInI5wQh7Jz8Ev+gVq2LIixYlHIQZISKexx9HTKYihnMVU83z
wtZyBL0nt7NM7Q7GGlEdeIpb7g6nyl0frSSaepftPflyAGlso9IDX6mIIUrN8ujejCiPOVIiGdi/
OxmhREvPGBK9Dg+aBLiVI7vcMnRt025Xw3KQDm6M4F4LuBfRJ6rdxEJ5Y9aX6cO14pPSaPaOPXo3
MGxXkCfpfG6Wb21elo5lw4V9QTGyfhjZX6YuMHttpANKvjI+eZyd5tmukr4mjgCTfg4249geuIIv
Hm61pyhcqX0i7Mz/6IntfSB8VlK3H0I8SotrTDsReuxnbT3yx25Dwt4GpiiXNfAkn6Dt20f5UAEW
igICGpCxMbqpkyKy+cULdAHxMsGg061XC9Uf48ITc+bpWSyO16fxjY4U8a/xskjFF8VytpTNda0I
ccmm/NEbY0xK0Uq/kQUfiLkQ/vQ73EY+6TcjDhicgZI7mNz7uy0RUmaDZNEAIqQjLXTRPKe2iu4W
2tDg9gCymWp4VbCZDt9JJfICkJbeb3TrzVB7oRGFk+VEcc2lLpOluDaw8BH7P654lvfHsUTBWpWk
swVgP5J0mQ68KfJLQT4zkG4EGNyjTrFkbCi+1RDyE20Q+xsEirHQVMKoOpGREP6wb4KxzPjYIhro
u1ZFhSkWAkR0FKhn+kHftokVUd7uSZGleUnF0VCFFVhleSXoJTUA3juVO1SVn3ffin9S9zOI2ShX
iwnvkdc7fE++bXrF7/HULYF1o9Q1P6NRIWoZwTDK36ta07Ow3ZFX7WjS+CSddPCxDIGYyyc1/ZY+
eO7GF4Zo4t+SuEgWy0KOhtD8B0NH1AZ4mpM8gZV12eqsmq1XCDBPPH5FC1KVWQwXfpFbreQIPUMi
Vwa8rH4JiKda3eyKSOqui8KY2QzS13KP3LQejwGDp/RuZMCmPQLlTvZ6MMXEWAYILdK7Laf0EYBH
sByOx/uhz283YPdLoTyh5vc4ry0VvbNxFdvGzBp8TbJGnQe5n22xRr9nOddbAPdSwmSWvBV983D5
tAXNsjAbaa//lzvan+hTK/TSyOHrfL0rYjSbkqbj45b3jk8QfxSGlgtHYp6e4LnS89XIkdeiM7WJ
aq8KcVSO7qSqq7phCRVwTV2d8NwIwEDvJGIkosYHnPdM6fslWZCCUiM3kmhQFmmzXS2vbIcdcUAS
hCZCzt1Z/g/bexhGLaI87YaVYwpjlwqC57zsKbZo2+wD7eeY1h1Ecr/+K+VMC2TDSpuGTqRnloT0
LQVCUNAxMBwI0R9G4tTL13ODaH6Ytf15IFkqaH4vVZ301JxUk47mGMVlWOE6PI7O6MfkuQrzwEe3
DSPG+be9pdEUU2htR9c4UhsWgeWaCYkg0/n9VaSrbYuulVWOWXtQh1Xh9QN1G1g9lACWq/o7TGqR
cRB6USP91zpzeHc6yhajjTJx/fwCfs+M7aOAyUZqLVhASvYMoUXMpkcacRrfecb32ai3A/5c5qGd
pUJzFwFFNmbVtT/gUZUyjBDPSSBOpRQKsBL3sbfeD5stxqLGRvfzP0jH4HSxrYE7ZKNVXnKlDo++
AKZDnBejP+B36WhUgJgu6R+kJQll/o+bxuov8GcYmxT1rk9xJQNKc1Z+CLJBnSq7Yse0px5bxuBv
HUIySxOlFEhmaBa6V8y4hrEyXVskKhJI1ukkuoPTNiTJ7UmiwNYQFECTTokOhkx3J8MDhMhKWw0W
fkH9AQExZpbzVcSyFkp0VnRonHaRdeK0ys+xWioThCwKvq37+LEGAAMkA6TcynbLVUDAn0e4gIbK
25S+AZ7J+l/vRrGW5x8f2M7XgRno39/x565qw77Z75UI4ORbLmJaFKqpgkw9cEqcGsiXPv7sk5NO
POAGFvI76S5K+iM408WR6X+uI1dl/9y9YCxW1uYNgYF66QqX8RptfWae8KB1RgpGMNqqyUdAYI6f
u/TLq8i4KHn3lspPu4NkW8jYUwupHZKVbSvR2mPXxoOYLjpl6Dt112HpeTjgGHdaFpsCeruJw1YU
yTDuvrbMSx0moTroc+QuZmGw0VBfwanoPanuDOkm8uTQn5UuMECThZtV9/jottygJ38LTxjtZ3Ac
/hch/IsMf+sc9nh4YHfpDCyxA8eMi4WjvD1UN3mP0PBULyxeFC6x/32xqLnF36k8DkDJxSSbWCit
KrH0m/XPzgFy5LEEu4ymJdr10GKjGo5+m8OgxTgZ/xZD5/YIEZGdSyq1OE5dDDCNKOgY3Q59mJxp
reyqHatIbq8b22cyP74iQ0GxL9RqOxr/wgoRGdvLd+PtoWoDuLeuLAHaH4k66GR0CY3whMZzAtzQ
vnMoC5wZi7lyDJ54nEG7ZTn/31V4Kby+v9vWIpy+1tCOddK5ItgNrvpSO/DId9Mi77vm4RnU/HUn
dewbd68eXuiC+fyNZ1MOkPXxPq1a1DioIOIcvVePPzx0lTAE2H6Unf0Ly6OBFfkG5OucRWl30toP
9qx/AgyXehcHW+FwyB8lLlJm83HmKb12WFxhdnX/XOsM+0pnX+sQCaMHukv2iajzCnJP6lj1hlps
joh9gCLCuxY0p5Uu3TM3d13GK+eoJTB9EQkilSIuBahhvCSB/Ts6EwSFMFqL3Onwj9wrhMfanQdw
f6jBWuRfZKJBjSKBdGV1boRZXiOi4w+5RLNJzp2zJBJTns11UOMagd5eE+NkK+XTqjFEnpG7jGA4
tLaR7tRmX7lQuZ/P4frLHdnWiSUDgNIgsiG5vGnQvjNxAEo2LuCZTupBSX8n5+TqMC4T+oeze67K
Q9kZoHgTvUHs0OVpED2gXLsA6lAYlA8SUrPXjn/HMTK+cxM568Llzc3iYD3sCTMFFzjf/YFqvLqC
pAhUQFormcJDkVzD2eK7eo5OUKdSO+yLUhqh3NbibIHS+WELynyTBoZJ3jct9z3s4N2LY3kIFlKS
vyvLkVHlNNaU/+zuWAH+ion1Xjh0VQDAOMGfzeyd1LwGwrOIIZJ7GUPGyY57R5evQWZ+Jij421pr
asZqb5qTBTbT9xqxrUc89DYyfLgZApdprbPuVSdYDjf4PCpSCtuPaHBws+anVJkT3c0MT6bRkCWv
YAkoaSPPgscr/0h5MRb58RNoO2SE6S4+ZrsmGcmSABVl05R7VHxpniiSwvVcewGglPWtGe7905S5
uMncu2VnJh+E72iV9GXzBR6AsYtWX157Si2ttzPcms2HYKLaBW13wfSmrpE14b5UzjhbZupQ5FWY
JWBLSsU+pLcxryAfvX+wu9ye5Xl/CLWrLRwLjrhS9sBsXEkXqsOSKM2zsOyVVTtEU6oGGtqhI45u
gKJdOYS+pEescd9R6L1Y0ivqZZeBNg5lz6E1kROaLxhLfxph+BE+JyJR0PbBIODQQkfR9hiDGUTF
KEYYqhMj1ispCb8YNJg5nfPSzWUcJ9Q9dZdipRejReMzF4rN0ywcunHlxynppBq7MouqD5HliXJU
rXe2rjfKP8TCyI9koryF0gK3G8OGilRIW0z2tze8oEQOiY2gg1r+KUyl0HSm7UjgrSBc+PYQIY6b
JUa4jBvlVrDyiKzMocIvxfHpJZUbVrJQL/Pz947Cgql1eFkNyRJjaVvtfaBcohn8R1UbD7e0kBwm
GyC0vSa28WZj3E09aFDwdDMIevkZrD/NCeAxzMrQ05EMr2IlfjLmU8hJ2asy015zDbJZaRjbOvEc
ClSWvJKza9pe5tYLzr6GcUB44wBHOXi2erm6FfIvj93WVAxnC14Wu+HpDe5YJiBTXOwtNY4AxU56
wYXRNL70SZ4gLET+ksIhWw1TMe16VWfnoe+EzvNcN5Ex91Cuto9vPHA5S4sK56g4p2TO4S3pLAGf
kibQ88YQ3ivnbcfM0nfCrcc1uCr37RDK1aCvuRdeL/IhuVMlOtnV/CjSFn/Om/4jj4LLLfQNkuG0
TCBrpsWnlckbLU6gig0zkXEja4UIQ1X1TKBWRsP3LNP3COaTi3IvKbJw6iSz+V/DcNPM9dt1qI+A
J2Co9RNS5fuywavovpBvq+0VWhvsXNJlxRJBjMR/LEemOd68gnV1+pjwDLKeVJmhgFRjZwMsTwuz
rQqSUv/JEqw69wEmTF6nkzBQ6O1JTX7rMTdVFge349tmOUFbNQ8AcqUrQCIq33TajMGBL5JdNABN
eNC0JtKUZFuumFh8jmazR8RXeuW35sgfP8BQDwtv0JY7YS0XSvpUuigHPh6djtuxFdHU1l5/91iB
Ex3P0ZQBx0DIKALx/Z+1skAOp3+0EG4CdW8hX4hn019i4E98tfPrYrG+5Lvgj2qd6PPb9yAGxiFS
9ZGE5lFwzJKug4G9QsBxvW9bgntTo147uS1hK0jcb9P6/g2SA6bzKB+ndNh2cBqMTQOjByqlTszS
rvTWCwQ7SySg94FYpykdsQ+J3SoeM8kHb3D0L5KBUDxHefD9OQ391z1l83Yt4akCkGqZqEGOqEpl
rwrfKZdd+v7oWH4QaS7IuXkh6Gv9WhnOk8+GWNShy0+eY+vzCcMC/SFLdxR0BiNDV0MIc7FTRlkr
MLzvAUmKe41m7GgCPswvTVIzq3sWPu/gE3Zl2LuYWswTX9sGN+5V0Wz+HaYfCTCZdXaP+8faPixY
eueOoKgKDoOm8WpLNgf/yutI7fYkN0lLldjo93AwlkeqQAJabAcAz0wOKazB0wpchOZaq0q0df4q
2kqQvXGk6SXYnoVDjzVKgEOrJtEy7ddbCTwgeZSWMctlOoRGwDFQBO5E4VlSC1Cef+fOQxzl+C2D
kpLB9H2GY7yVtD/G/x6O7wVayYL/HbGIeXyvCKRD01mxEG4I+NRXRV2McGZ3fFnXgqkubUfTpOGB
gfP8TX6xZWm4LdWRjaypD3KM7+2pgLFd4ABO1xphWcJ9G+0LK84x7F5kV4TbMYeoRQWzw6K8JUMx
Z4VZh10Y27bjWFSxcqkkZ0btkNZmZ8vjfFY/9Tef46OQXSb00egtNIamvIKZWK6xMGbqS/IocV+2
Gt8cN8GpFMD6uOISb7YIKB1Zn9rRg524xXljWtwGRXnG/VV0MTHTCrer7QW0Crjwztuklnxksby7
mOS5k+MQ+qClR4FzyvprXcoRUAKD4RjLPS+1asbfznhIiynNuNVauFNta0cg/ZUjofp3ag7Oj/yd
TmSgGC9wg9tUFm+iTYEJm940NePAaeSKD5KG7r5haEp+7Kn/EdSiLI6iVP2U0TV1mbn4wocgLTUn
xB3cEwpcttzWzuWkwy3Qn5PAgQHH9o9I3ZvrHjtECnxldkosTPpUTH709RRaZ7NGh2W/l4tpS9jf
EpH2ANYWq2aLfTaxr/v5fShFHDeBjq08CRAH3geghlM5gRoHcQMPmeYWmkitTnwC8o0FNwgLYhUh
m2RGPmz0NDlg8nDQ65UM4dZxUwUfOmOJDGbvXxJlKuKrsKKwG/dfY7kc//0MeAwCh1V+pY+VI9Kx
xoXwH4ajFdiWe0WtVv2ZcB/eZrtINKvBVRH/fLB/l8CGgeeCsDa4jnuqkD8hKz3NQJpP/hIKFuKJ
ouDChmG1Ujmi509VJorzgiNRDAjNK0JbwS3WzbC2VOvd/QELT2bABQJs7gyp1SGXlXcvHWeLnDDx
DT4ko8QaDSYLHpt0M3/K3943zHtuPZBNWPbHHsnXASVjP7VFA9ZbTfA/9PxQtThAb4xFyljG0zbT
GPsY40zVbloZ1mDd1mthqj9i9v/VGJakpYbd6jDK7wMTdqZoaLgCrJUa8OYcA67jKPCjX5BdfbFq
Zl+qbd1Xvpf9VpP/cbZXB4SXcyaX/04DQLYTBrKp4YcIq3Bf7+mu3vZLzH0H8/jJQ98toZGFS65p
zID5LhrbriieNCOx9jV50wxFULOdCnnguMfw3d53nHTvcAkbNI8jGbF+vl7p5PpZ7vjunzjvvC+c
VebBhvF3WOAfKBjG1grCs1Y8ufvCShGOcAx7a58yHXC4CHIQ883u2vMu4itvFQyLBTSPgiMd+tSb
pixSAZ0RxLZlfSohvlVr5U9HMyGed9aLu+bgCIFdDj8WZGz1f8hzNp6Np+Pb88nQx5/g/SWoTDXk
j5j3N00krHB3gwu0Buc/6yz4LfC3aNBqdYhHSgD9UVpWQY9n2UG34H3Tka8TRKYwesL/8z7Cgs2v
w7PYXHTkIuxgn86hidlw92LlJbe1oPL/WSnKW1t1wqVgDp1BWZilMZK14+E/hbYNLgd0vr/tsWI8
2QKK0gn6NL4T+PeR3Mb/m4yOZCfJKp16ocUvpBlnMIPOYwIZYmDpH3+RycDQ4h9TcK88i1jWtCAd
DzNjCi3MDjG5QzRjCVuCw8eIbNT8NGN/Xpna9k7pdIaIhP25rz8g4L3o0iBZiPR9RUNDMFgi5K4m
fRmgD/R8hC6cv9Izi3hbENuXVKlnjJcZN2Gic+503+IqaPIYxYSVegjB4GbHPSPOKY2RDyCLjU37
tH0QtNGQ8/6xI62VE4I5YkQL8L9r9paH/r8gl0ojNgvnFr961LTDshr2J+NoObS0JV7znpPPPy78
wpxxFPVaPjrgiwEOcl2SaNAo7478GxCjC1cwfMXxH6VPk2OBJ7gdYknK4nswVF2Hqy+lqTTbi3If
18nGkR1HGaJ2I7NZfOpJ974Rn4o4X3TzGkU5k4SjiUf8QdTxIsIoYzVOg9yKR2vKFq5zEZiCOeNG
j62z+PGd2OijQ/jtrSS1UJqKX7d1/s9R8pPFNoq8l9tsteV6ocaCb4sC3tyV502d462DkpG+cjpn
UVKBhZ8zG9+xZNRUqTjM8FlaNqSHPmf3+MEwebxQfSWcQ6Vc41TRX4OcG74U3SEutXt20fi7Jr3x
skkX3OP8gA39CIQavjYBr2MjEXbSxWg85AfiarWKZk/F1YWpk6I2N1d9xJIVQvpH28+hNwxYRoJk
CQSCXU0m/EV5jKpr1OXsm9l8GP4QjYP/+4+L6NM4qkqJofG7sOqTCXh0nH/azjW5cO82zmkExaNi
Vxr6PHA9u1FnfRwiBMzWwhMqwyFJkKYOO5eHOn3F6vcLdaEUUzL2FH9T3/r1x+jCackKUzSDB+DP
hcaA+Cmn8f/MKDtJmjtxLwfzGtQ9Wwxbs//8MJl5B8JC7IoDKwz4gIMeBKxX6PSNuLaULjZNp0na
zWXCI3dQT+soWk5HMrvq8W8kqQccIIpG/BetdHW3Vcoap8O769ZJyfU5L41iP5Vs6c/a8KUqRGyN
5HUfYdTQOmfzse6Bd8uHHoTVCe+Xdire/Rdit4Myl3Q/p7ONXoC7UaU9VrGRHDPIfRd7Fug2p6Zq
MEZbuIDdMBH4yHma54JjIYdVD6R239DHLx2pz7oI2tWlR6M0+MtRBw3TbpR0lftlx8G6HJb+WjKr
halApM64XBsk6CBx2LQ/SfiRyaSRlzIrV7RbMWD4jYJQb0/LUcWqT5gVRNsv0eBZfE9gXB+APfoJ
Rzq+Ju2vtmI/gV4S57bG7YNjFcXK2gl2wNwDdUYCiU52r2qYWauvUFdH20Avbprsu/csiddvsfsx
e5/COx10lAi1r8j9dcQ0FYxO74ZOXijoN03k6hSTSywqNJTVc5eK2Uu78p61d3tLo6mIe6jItsnw
kSIXjGTQKqmN6hK66t7FxQR5bvS0KNY9jrAwnxkDGPi+BVD8tglvSraE8685L23sG5TifHeWDfNl
XKT+8k4gTheyFM+VP3bH2rDrkDA1x+peCOLvdMMl7aHDnd69bwvQ9UfVJO2PbMTqaTxvdgmskSp4
y3kkoPpNvQ3tEcz2INcMCbTQ89LAzmQkOc6do80VLuiAsJNRam0i/3ATVi0EYXanBC20mLYSJnDv
JBxWpw63Cz71+4phA8l6HL3IU5eB2XpbCUaZTtZhzSyB/8y7ITFI4gMOKRDlpAwkPU1ENk7NLJg9
AYiuSvB1IJBNE+MuGavgOza50eJp1HFUl/nDwQa+b66JGoOj+75Wa21i23StRWOLf/bKDgpKeRMw
Ms2WWVeGZ0inu1OZzvROZxP5h2huhPW2HswIFduzyJJLgsOzfNdgInP9YFQrbPtS5+fQNQsCvsa+
a0WQBti+1IQKeqUAOSXcc6+fZWIq1ApdxZuEQlvPxE1mx/CXzTSnlmR48LrnEKlY46Lv4PkmBJfA
G0Eu7cmUQ25Zz/2j3lWAC5Djyb1fTGX2m5eGTfIDhZHLgTPEhQYPN/aKPOIRuvLUX1lwEjwRhepT
MIgmHCKsCPPNlv5UHgVtbdzOG2bW9D0fPylg/cVpklsPluHER8ij/QPAi0R5GajW21MrGjMneXNM
caXU5uyHkCsvCgE8Pl9OzLFQ0vwxBRe8uC5+v7WcuKazy0QndYVKGLYFjS4D6zLKGTQvphGE717S
EQBcSNtnZ/NNgONQazDeBa6IErBGT508mMwlO4jHKwMj4eVZZ9vYmO/g6dfKW8InerS6m2FKFmTv
XFg42dl2aWuSug8dGe9CLSZ06WZWtCHjIWRrD7xLUTOMk2Bpx8tp1hc+sVt/poF4/3I3sEEx8fGK
hWOVaCY0u6quYxW4YGphslNzUzZ59jBUYWPkh8SO0aG+Aho2svET55ZNqJ8uRf/6RgoXquCVEWnc
jZoYuAI71K8zrKcJ5eJ+ug/mMQNn1cFiaw3SMItekyCC9SKEjhZvPf3fwIogFIgW34ZBHM1Eq4eE
SaSGr5settmr3/tKg3DonIgcbedlU8qeQwv67o4FURhMoLi9t1uXQKUGgx1o/dio1qYjovZN2ck7
Y+WjGAMzdHYietYV2WroEzFUSYvFy5CWqbqhzFbCfUc5pXm8UEZX/MfPGbWOQqtBZqjxMx1wFeiU
9ai5yyRMBA+YuKm2S2snYuuwP2jebE1Lo3Dgt+G9fUdygDbcg21TkMB+i8Oi10aoWMNjtgViaEPf
y9EjzEeJm5Nc2i0EPMh7icyNm/vnPJqrRKMPsG9K/DYu3rWhCJvsBExzvZDEjcVwm+lMLhZcMGcT
+1Od/NUyi6FxQpUROxQgXewcleI7Dzp5fySTeXtECJEo+/+t75jEbrd79yIdTO+INJ1JcKXWvRLp
UdXCWZULMbXJd6sLnTAiE9adHshb9HeTcBEf3/Xulb0awnFGEgy89guiDil6wAy/F/GATTeZiCV0
q+TM/hgjwj64bVZvRauoqUIulLaO7+nFSDriZYGGbN7Ub7nwmmgfqliPO80qC7+m+VoU3lmHw+41
jO+7oLUmsFtoZBTwKzm4XgmJgX0OHBwzFl0OLwzbGoe5MTls9u2tkYlA8g8QIKa4Y2/xSBthRzx+
GnNcfZr+kRofgS7rqrsNyd+MAY1+ItiorVslucRTjuqwL5hyJCEVZTPlYFxU6fnGy1e4fXlUP6sC
5Gt8BKdug8hULboCU+Fyh+kzYQftTXgRlt+1RAXErHFxO7upBpom1T5ZFIHe4xpjLm7twDr4FFio
B+kIfwlfcjn8rQbrYI4s2u5YmpoZa23Sr5Ngyo+fFdzUNZX3jsX23OPSiw333ZHzM3nWe5IOCLN/
yTse8ODyizBZeaIXCVGJsRpKmgHEW4/lLcDkkNQ/0bUiSyaPsRklPO21RvK1c25HPwA6rnkaJLKD
iA97DrqSY9UHZCo4BEl2jJDSYNh8fOeyzd7uMeSJadNIwXK6WLuX5mgfRiT7Zrns0Z8RLku1f/sZ
kl/INUdKrp5lGGJm19hmLZ70IWqDI5omQqTW29KRSqhS2sPsK4YnQRyCNVHR+vXfejNZuuksr0WE
J4K+gO/JKsr4aH+F3lqQYm7CNBAjY9dwrTu+Jgkn++cr2te68wlTN+MfPdvO2JXLPPc/NVZs2FZr
CYVstskS8whrtvCztkznC9+4P+JxlY+MqpLfxf/Q7cPLfC/uS6ro2YqhxCGLcPoJjA3K7xmsIbI1
MjutPLZAGKFNxcruVu8bHNmsCbec25oqwHML4HRlKi8SiQVUOX/yMOSekj7NrY0P5nUCfCsqm1Hn
ZyWefYxjeNTi3BVeenRCp+6Mlu0TanRoosrk7gdqb9CFic+7nQ3dDXmBy3Dy4GkDQDrTY3rN0KND
4A/eszJs0/pFHtc5B0MFxsM2HjkFCdBHh393bqnDJzgHXebBlqbbiYUQGZDZflUkGdzCjXJY/48f
RXpzZYKsViZQW4UlBDTJ9ZxUx0nYOEgcXcF1iSXocxO1Bq4MDIuShs4lpuVK5hs+9I9utCOL9EFv
ye8b1Zvd0YSZ9p7jR1q/IGfHpdMLftUo1BEEc+Mv/EZIEnblDkBzZ2oWbgBzApdUsOx4SQ9XqZJU
YXINQDrSUbJaieJgqEiu7MptxIIqifD/KP6cXYFjBOm9fKTE+qWwFAUbD44RCTEQDwpJGCn8veU2
EuRLKj8EmmGslcYut964VV/65tfspNvnakG2AyXk1/EXCTm+wM57iLppzZfR78Zbx+trZr17FNII
6GMMfFPh8/XpVw7SKCm7P/UthanKrbpgTV+oT9+ySLHgTux+NdVO9t2XQDTYNUCYZ7nMuwoItX0Q
ddfdAwpxOKcizGi137v7KLE2phaWYf9Z7WFTIto3OCSHJi8xj3L9dPylBrVH54W2spojSkE/uYvJ
2ERzz/CcB+890gCBxLac7rUMDs9Kaw17gLBy3sSXT6BBlvWyauB7TxicQ8PT4Pma1Kgga4P0EZex
Srd1syBRXalypLIR9huvziDHle4lYoutROwGSv8MDM/3bMNU1+t0sDMqhhBh2D5J3dilTmDA9yui
kUjy18fk4jE0hfty5TldEDTmXh3VAPGImY0MIFSCPgr2q5PRtnujA6alssoiHBWyfUEyAof2lxFi
6q39MS0gADfNgVDiW5Q/E/TMUfzbh+uiulSaXWyYfu7LyinIo0hjjBiHvfhrSXbs2jXACXDk6qZT
CKswmmMt56WOWKPmD5IBOfuSrwNbgwBWA46LcYbqFB3rV7pkD/eHf0kjr5wQOhKOaFeOH16ri8jo
FU2l4KmeC8W8B8VkwcafHp0riGQS/Xi3I2/qePIuwmAy76OHCW4fuit0W2L9Xhx22N+i6sPBtCDd
xraMzCWhy17Re9g3UptY6wdyI4iCUqQ1Nx10UagxQdW7aZYf9UcHxM4XbLqWv8X7og26mr3sVz2a
sktblj5FC81eoOWb90hCaVCPHT0W0abiMgmve8fmEBBG7WXustwfVz0Wq2BkEGzaJOu6J4DAIOVh
IsE3KmTEtHMjv97rhoVhfpGPw1QqWpqkZ5gAbobilMUCNfjqm/Uh+d4VqjvkUeHJAXC0tB9jQVbY
UGt75L2p4XswZ9dBbUHGXr4O+skZdg3pjJzahsbYGRNLCL69oXYoFEOoadj5onAjal+2ZsJOcYSA
Tht4z+kLOb0rn072RVNXwNZwJLZ01Pgba01wXovO4fNAdKZ4mpOPU2Pmwxp42M/cP7bacKslXobk
sxCYC0bsBna8lK7pM4hSKIiXwW2pcIpDLW9hLmECorYu3XSrEJFUw8UDrCl9joO+ksj9mp0CsQfc
yozm2zbLZ5rkD2xck1K7kJsGzm5H4FIHys++Bh2pZHgf+2NBGHDWxKG/JEYbU2qOWrtxGoKxb0QD
To/vEAEWCMpYIpSE+pc9JLmLWOE8E6G8yLyoA4IWoYdfJHD1BC6LRKDV/LBa5wTmfGi7b6Uoi917
PqmhEf0aQPupPq7bOByvtGK1QUpw15CoVBlT19A/FFUpMEoG9XONLZtUMOv0MuMQaVOeGVYQdDk7
cPPhpqvIqArKN1QLKB7zbtqTEtzK6wf7IHVM0gRtzO0LY1o0KLl2zhUQY6liPp4iN/3DGe1vauwS
Qw0ojJhrq92LN2WisunMXkKbT3Tt88KqlOfjEvuRibnOkTvmGmzt1kE1lci235INSjJPBbG8DN+V
ZPRJDMkkdHIle7zahhF/nGOoVv/Pc6bMi+N1YMD2Q9HtGzzMKedxnS90q3yVnn+TLYTQrf4tCF2A
MTKTLt//wJUKThPdxuHKW2Db+vbGNjeSTbH3RPfHtd2Ej/aufpvEKdWYN717gDaF5aidHjjRHob1
CrLIaOc4LcV09rEuz4pzq+212tCcRAIys5+VIZqbkAM3B93dIRHQf4wJ47XPb0NeWE7+GjU0J/hs
ru+Lr0KAMHMspGxMxLyoiObEP9VMSDHdRkx2CKtyVpkO8Agm7kn38mb5k9RmzQSLbpeio01NDpdw
J3N2M0BcnzcJV8vVaTlQ9eb1UAjs7Ukkxws9LJEJXJ5vIJjfa6q018DXZRd+q2SbYwv9hnA8Ylns
yophzEnrl7WDjKaHDelBu3O7J+xd9itWEUaODjZgqKB/cCvSLgex8Mgez7fWrsvUuivQTFdnaNiI
nq4VbocirGXMXMwahnfFnSFVj/WhtHQNUvYINIfk+mL46ep6QTvLvThTvT0CPzFelUEn0qyWe0fG
w1sE5nqvv0ngePaZfEbD5dzM6ewCSbt0O3g5YP9/m0e7Vslb5xs8yCYeMrXCerBT4HXU2zJM8pVl
20D62nrw54d7LL6nWHL8qaKC2S9QkYjctkx9DU+zPFw5SqiV/Pbt1c0IPCouHNxy9mpZLLLnQHeU
L2tZM2uRrIx1+JRvP2xcfKvsZcWXYZw31Lr6YrbUHLRsodXed4/c3XswTcTEjR2EcPufTGOSnlU2
heKe70+QgLa0tBAPw8Hyjk44+pn9ZWWE+k972fEj4Gp+AcUrUk6g87FCmgymSDUgps3JVbxdwIWI
XIoTTJLRbp3R3wZCEi+oKXZTtn7/VEMj9PhM+szq0aeHRT7leBoEpOQtFQP6HcCCAQUN4amrMbH3
m0JLPvSRGMxjFDmeK8vm60ExFcqoQ3RL4J1O2trS+Ru5DftmzGLITBW+oFqbo5eK0saRZUwffkIe
TTTpRQcs4bT8WiN19oJj9vo5t1nbpuGdPKiwVHUb/lAlS8QdSgUGCQa7a6fLdj5kV0Qn+vIst8M8
pkV56cAoyoZ5Opd/5gA9WsvQhZHzZmv4YawEA2aef6FkRkwRkSld7H+he/zjBYBzWenIl5H0rIAL
01VwZXFXoZh4U7TXYa2dhAaq2pormlzBLaR42ba/amWPZRBVdogQZQFbrFBaPmSNgPBPRdYGq+OY
rLiFK5Xg/TW5Y20gA+egUlLzUvJm0RiBU7dHrmyjmUogqO3Dm5aGbMs5yOf75WGm0+v293+WnY0b
bcLiRTgGMUxwUtVqYccoheABg6BEffeNUwUGA4BthwzLwOOpPH2saT8v5PeB39oeHxEPr9m6dqf5
REtAM/65UqIsyejW7OBji64YqUUG9M2OaRgr6xlv3iYwVN265LvESFTsXys+u0oOrh4tV8TFEfqG
CjYHG+q2WHpe8B6MNYvEjTvmN5O4iax4LUfLL5QaQIa8h+CTmDvuTGbygsROwsXE265VLt2tkvK2
1fBelFSjLrTU4T8Vo+RdT8TZi8u18RQU3IA2ne3W1wKCHKkFitw8CSrXC3yJ4Ike8F312yxJS6em
XQyZp2cv99Tcqq5vtTItRzF/cTTEhoA+qOOn4mUl4Agi1pibgtFPPi9JfQPBatyfjwRnXnn8bMcJ
P2/pToNfrAy9LNldNVTlyJJFyrgGI4743agaDUQpqTEKLlfBFDtNy+lIDCKdb4jgwOEAyby5s7mL
S5ikSLkD3QbC5IzTlXMEfrOoQAbmqRA4F7V5wU+Sr8W/7yhglClAnfzIwmSHih0NjvPREGUadAYV
/sil92MDQnkhIuiplCu60Qy3N+DMGd0+IoRkAOox+ZkCccQ5tCQLJDWSRZkwnB94pVT5E3xWtUyA
ZVv7YeJ4ChHUx3B7XqU2A3m7xU3gYVBbT7U6ZG3Ipicn/Sb+PHkPoOpoF1k5wbAEe2qpl2L1KP3G
K/JgCXkkMjS/mKRs+YM0RlhjAgRhqb1cEMBZRbbcH8kMDVRW7e51Sob66eLO2ZlBWaz6EUATfmGm
n+XeX2MX4+2iYhICXuDamTKCJ2ue/93L9oMJah7TBKe2Ik25lBmbpqR3lVMy5og60p8YKzgySLOB
fynev31VbEo2vTCB2HHu2ViYcN3DeY5W/OVYEfEXvVbGN3BSTYx1eOq5BlND03Lqr5phSXR3eCNg
upHcypwETf4OT9mEU3YTxvb1Ai10HyFepvhUeDDRLSnbPt2taf2ucFVYdwvF9421y7jD+tCo6DBx
qhce4GMJC2O5TL4pQLAFGs6bwlpuEVbryoWki/+yQpXnG1RroRTuI37wqpm5IEi+sDUlmsNa/266
kmPaRHu6su75J5O8GEAdFNT2+8sOsDKjjB9P06WRCfS66R5T93UbVf7pHoNP684GRzIreq8aCI7X
djN7Z92h8n2H3kheidFAJbwyPpU7j/XgWkzUCklZosQ18KWzURE5BijT2vC6zuEQrKDnqdbGJgTW
lVNPQv8EZKwSV90/tk5Q1Bwjog+yMVJZl6VVB3kfM9XSbBZJtEgmRZQcaBNJ58pf3kSdkHCMWPP4
CEM+p2C9jCGCHj3Dn9wbgJC4ccMIshDxhnXMEbObknfV0CGl6M7QGxNr3vls8vo3hOKmikWzR8XE
m5CmASRaJHc9pL6/hEInoK6sfwHFOm7f8nG9eoRpqW1Qnlf1uh8bQQC9Wl/qSsqrSDsfdSv7PqPP
kPYt5ixLPLXf20iqcTPqgSN6/b2Akffx/FMvJ+rlYNypUAJIYTcvfvE8KPYDLIwFWrmrv3BXt83l
FzByPpVSvWwH+3otYkkJ64xQPSowkRT/vjg/ouP4sZohLTwEJo4dQkN+oUMA+aQCD3wN63/0G9QH
OkEOyeuw6DmS2FWetCN3bTNRpzjLzNCiZxg0rriQSsEGnNJAtqJJ48BcFnn4dUKqJGj+97JRsuaE
trwgROsfncXOB0Pbe7zYxHNOf9x/BLvtu5jhMxs5NzIpJtIVD7Bkj4Pq6zFoKQAAW4mzUPAsePY5
BCXwGOEjf6wf6/bsIY9kzkTEsOPXIrV5KbCb/wNwDkigLkFK5lALORMZeQLlrZKznggPuF6wyCo5
h5KnbbGPZWWZoFDXlWAt6UXCU0liZ4Lmyhvygb1eJgF6Y7YUgpQfshJDEHex3pyNwEiyMRVjlBVm
SqybRqjtydUqHunoMEJYKfEt3nZlDHY6X9uOulnaJvTXKxvVcspzwhQZtRtZUXb6MMSHvmL/EMUF
GQ+lQzAmhfP1J7PmhUm2dstYWH+2LlXujd7M3LBX+Y2eYcHgc6YUmGNCDsDcf21BoGyHPHT4KSMQ
h3GMCLtcJpfumdF6Wgrt88FEoxXS0I6OtQ7G+oyFT4pGt0dXY4mROap9zlqmRP4QJWGM1Ed+zE/m
7BWyitWan36m34Cvr9n20U04Zp8OIJBNhdHi0GmUe+yC4XqPSJCpbNXh3MhY38yjHYKeX1CNOQyQ
UTjQBUj4TcIif8nHaaTzx9StAlPpxGswOsUwUKMZZfuBLfeVIkX5tWEh35kENnXyDCHQRS0DR2R+
XF6pj4FylTZV64ivYn/wk854tMbe7LCHqR1gNod5fE6YUAu8EIvjKva7fZum3tkIHwNr2DuYP3Kj
IcULoJGp5DLWOEGqoE3epRGXzmHwoONd4p31B+PxTDUl6R/lOKLupegJO8o7Y6gqH8RWXtCkxc5L
Br3knfcjsCFpmfIZtuWxq0NfRMH6ceXCKsojjwh0AIOLtbAQikFLnutl80BjODcd3t5Cqy530ZC+
dCPOY7Xo6xQV8/e/ckfAB2pfZfy3vJ5KHHGIrBVGpb0IVBqD+GW1TeFa0VJXGd5j+/C73z+wqYJi
E7OzX7hivy/dF73ZPfjjVOZtefToi4s9pkkzYRPUbpStva6QiIvmfSKyzmNupxGMFwb7vSX+TWpz
8c3SGosVBB7lHQoSYRh6q6wubLP5CO+dIuDUTrUAq4EwuZVbvldhXAxITMj/JPZ4TZUVsiXF97US
WtGf8mn8naeetoJvO4Kx8Nvbm1IkQVXLvXsFr3MTDIJyNnuRxMpR+xNqIcpFlEke/ANgn2UTg1Fa
SqgLFPEnsoLztT/B/E4Ry3NHY+5XuCBu6SClkAgYA0yppnqRG6Es0kUgJ8rUIPfTQqx6yB5L/kEr
lnYp4MZoOwSyCKBRdD99/JsWO5aLKu72F/C65oDg91OdDhGm6FseN5r+35Bdkzsr0sSyNxaY9HU9
jYRDYRNTdSVNLvjn/wxbOIusbafUaYddUeUlrKgOzSihyAvU0LWGWN/W50Ea8RhOQFuKPMyGvjAW
R5TIxrnPXZ8xOaHborjDsGIbjEIYXV6Ymwu39gnm+G15UylpbLFVQCqxMDgKVOcM+R/aRWDgXvkg
TXVU4tk3iUwSHK3nfWZDzms9hgwWPm0t342CtMUTzs6n4EDvu7uSQW7fsbzfe/L0h2zuTTwlb+3j
2yBy8Kx/uvSf7CpELlFv4SKM+6uV0BZI7u5PeTYVtz82v/g/9oVFtV94PpzYaSmHyXyKqZpAfUNf
TDhBnOYoIV8QP863sLiya10fnNDD9f+6O8idxeryIQdzAO3pcvt6Y4hcPzIjCiBYF4qVhFuFzBr4
r3lSd2PoGkPOMVS3cw5xeEO6FSUXYCJU2xwj++oTOMcHq/BsLBUz1sPpIGvDyP6IxO9XgfH9u3nZ
8fbPFy+0sGX3idrNnE/zhEyL65R4oSGBLQZB5yRP7kLotAOrGjmTsasjEQcE1vXiDFxKA+Pmz9Zo
kaUJvmbGg/BTnlIQYSaa8bI5o+Wsodh2Gc/r7cuss7uT1lTexeJFGf8kNHJRRvmFiivFHPq2bd1P
OyC4Dn8g8CboumbAD8En8v++b0FzLu2lOp/j3z4wmgWnkatliq+gzePoG6a8pvHSBar77xilvEbE
LLky1vJHJ5idMjF8CLCtR2a8DqYrPqrCZ28ZS3jI+NtSnTKk3/otux6CmzWojBobstuumWXSUS1A
HDOd2HMzgSTmluxL98awfvGuc5v8GJccnoQ/PzGv/2bW1rzDr06gbTH2gfjXfw6SPkmkwvmlq3Ri
XcoQ9Fw6JWqa1Sv5w2+NwUbFKJBOz7xjKSeaALTL4l3YLARSHT4G2dCzbagUNPkGoH1W76kRaMv4
SqvFS0fJK+V/I/oYZAifW9moX8qAXMryAPprkE57iDFjyz6Uou4Z/xV0ATzZTU+8KlylUipCdEdm
KNf6JeOgOehBoeM0GDMzQFcDCnFhtW0lXwi63VJaCfxJht4oyhP2i0Cb/HXHjvXSIDzEFaongmc6
BhscCi+m8x4v1S57G71PcZLh1uQYv9chlbnPbPinmm3rqeAfjn1U/XV8PkVIH6jneFxwbT8It/Tp
siG/YVj7AP3kMO04Th41KvSN9Se2BJR1/OrGzJeMqCszAA5NGUTmUnynHuIru8UmRKbGDlJLaQUU
TPTjklsBwiCd5Ji8g3NTq1XtwdEiT5Smg01Q8h1lLQQ11EPZ1fii19gSsSl9mMcTdUF8LVwlzXPv
9C1MSdFSlbeBNbGXhHG1Ruhq5Lw1aNzwnZaVmMNEVEVAT/Zg7M+HlcCWlr5MfJSanjI1HF61LNuS
IHMutEEXoGtwxOwEeaEA5EQ6p5ijgmW6wVNcf6bCb9DKPKXXcehlFgIMWq6acARrxsw3hvTNBAng
AOIRKhIFpRYmaS8qTZHGoW7+w1Fpk74GBYRZ4FsblgcdjPrvD27M00YDrfhisDH8M3t2BBXjGmS6
JGGvHf5gG53UamRZtBddKENPK9vtIIEzcGZnwVWN63VATlUfXDiZJ2pFkkhu8faIuZk4XatAyEdf
B5NMgGNVCSmzNJiNhEt2Hhz4nehpuY+GRvPwFcyJQaCljujQvxJrnZfmw9fy7x4qtd0oQq2f5+Q3
WQ6xMRkRW6edLmMMeUXnQ3JQMbmwUMWeYmYeXDcV0MUk22Xqg9MZDEClnOIMyPiYsPPNbXAbLo8x
5s8m7YEg//1A1sFybQ4LvOm9yYlHqGrERX7+7zHkJp3Ue60i9DoS6tp61MZ4l0ClTsWB7h/uSnbi
azZxm0oPhspDp2u75OUT/01Gq1pec1Ir90oHBA6pgZ2yGLQU1Vf8l5if+qHE7JnFMenq6AUhH1pf
IZJ1YGwkOatHPr9kUHPdDsTvlsLQFHwMd4cz+rjwq+5JlgucmIzl2jnnkCSsUpQot9wLS78VkH4v
W7NibK0FeiWE5w92rvNgcl6mr4WH7X+G1duEoKEwSaicaHLUtlUD0Tf3e/vZ61y3IkrJj8ek+tq9
Ovyaa/L2y/LN49pq3Bk2odaCtxYJC59zHmEa6yXy85+Nz9gA848jGuP6B8csSj+F1Pgnf8FCBUZL
jAqRllgw5B00+Y6G4D9f3O9BA/EbUFbY1dLOUsuDTdK5PdTB/FdIGy+Wnv57yTEgRRSOvh76pezA
FS4tk6FQzFhnJr00JlsxM1m2aTBNOZHNIPIDPgQJjyf/4EODHgiyuQu7uYF9Y7GOBB5cuNTv5xzI
pwTvMr4ohCTE1Um0YJOFVMfDW6/O94rghrxVwG2cWZi4zbIq6qzXfOp4SWSnm1pARGBZaCLnJNxo
lPP6MYcM3cdnKV9yjvoF4T3v//NuK8oIHUZAkxV01skCyW+wWpPPoVUPkV910HMnlOct92gXU+i6
E7B/Uq60M4UzhxzGZhPNLt5d4PR+gG5gvvErG+mM4bM8QzTT5yb7ycIxnVlT50Y8nSHYFsuI41eZ
m6vwGceuAES/s0pAvND+m5E4jo6y70pDjpbwmmax2jJIQyKI3JWNQDAvBBKFsYJ2wJy1Tfez1x8I
yo+I57fpLyqdUZusSfGVuuOIbL1u7zZxjzvthSP85i9ee0+sznfCk1viKrI+wNu+d5Gx1j5HpJ+V
ZPUyNVm4M7Og5p9Us8pijfxIsKQ/8xjVDjsPGfiF9L+DloB0XDgdrK9PZkLlcZvDfkeGJQ+9NDZB
dc6kkNaly3IEyQ/qYarRZpcX5qKXoCKSmDMYwbjbenJN2aVBDz7Qclhyx1M1VlrANSSeAGc98lxq
+LRSScHBQhRzWuoahJ4mN3fxALNX7aPCeQeJ/7EcHPa09q3jOha51R8K5eQGn/71rV5hDe4iXyFv
O9dZ3dYDwp8JDGlNeFaoegGgOboQE+lWCYafbw3Sj4VgzDo9j9qaZ1+yIVsIzTERj+gWJ7HhmfPP
CIK5eDzjPmu/+k7p+bKTVdd49indmSiDuRoCw17H5C8adSd27khoMZ7S0U9OO2w3LrzUsnVhfYoO
5Idhx0WTPFlvMAAXa/AcOvowyS2eEZPxv96ek5kLigrN/jwM5sxYRsjFGsGHhUTrNuptMwt5f0Hr
zhE7w6o7SP97soBilLL4aVu/CjLpDwS5VjaAzbcZFRjt3exwYgjiEHc8oylBG7jaEkRFW4LeLrEb
34guItAKGcR9jLG9eykl6j6fiO8tKYbSZqERjt1zQY7Kcm25BFth5UWmn/TWJnkWahe1snxVc/tU
NiFxEIKxv3tVxHuORrVOuZJyzZBegnJwsVSOQeiWoDYlkCTerThVgaZ8EtvBj0qFVi6MHLIoYO1H
TLETKeh6rFl+JMrf62OS+v6JwecT8WdGWLWwWXy+xDuh6e1NpWBD34Um+/EzJneI8YKXnlC1AorU
+UNA5khdjDYn35opT3vvKt+xXVw8ncSmfkUIQyPodgLCkrbigVLkTjwWuEkKGy8dF3Hlk7JdRa/+
31Vcbrdml5QPZS8e2UAPNN7lv9kT+zKv2owRXVDfdGrjt4HVwfDjsFcQVDJXmjvsI2SSiIYYecQM
3zMfYgZ/9k6Vyec+U+lF5gw820O0DvR6lVqrzevftdqiRMAiQDlgI5MXh+BboGvZI9ov5tzNiwC/
TKF+O+MjTTYEnq3eQe1XtFt+wuOOBavbXKQ4ulBALb37PyO4WNp7p7dfbiVyxkv8VQ9j4FHbFGWe
bmMAha3B6zWyiux65+Z388P3ZqoyNr8BO+VmMb/INui9ZwtZH4+lK8OGQ+OTwAVvSkHkUqP939Ot
NV5ONaxSLVaanaYBtpReQP6NaP05AgMOTvmWj5FzucstekF/v0/gMBhXlj11P3IAtHYNUaXeOx4f
D7G6i+R78i2nB7+9owvCHVQlhWGCvj8dkQKafRxnNziNkkk16VK35Z8Wekae9uVdbQo4c5C6/5WD
yEPML6N8TD95V7SCKMV71lM14lGcP/MMLb27m12aHJ/sOC+2Kq1IfhEW60zBok6KalP9rCBkKEsv
sZAGhq2tpUVxdbHfR37fgaYD+lKD+loovMgxzlGJ2KRgiLMPwDcmNkE4KRjMWcB5BJw6yQYKvnfl
9zjvwk2FA6odt8GvYF9YTV7jWjjb7NPyyudWovUUWFrScIjvPkPay4hmyxPpOVsb0moayyamPDNx
SgTkfbFruD2CFUVlfDapQ5nmipNqy7ZDUbGdmXZO+uXDWvOi0K2yWC1kKCCXsRbuhMvbLTjQF9GE
7oQxLo3xaFVT3jdwfbzCiJucfCPfLNteIaoyYc7wAtyuFw6rEHomSf8Yvsd4/dJ1k+VeG60BACkk
Z51x/MuPcWgvkEZ7ZZF4NiB16OIGhYP2cWuXkHl8ZLKKsVbnVWCKduy8U1jrHF72p/q/NMEUHnlk
T0YD3MXLz8NyRKKWoTKM9IZQ9basbWiePLmpEGH0D7t2h8tgLGh0GJOSNTOgITH3bO+uQlybNjtR
GE6kL5NkTogFpFKaR1HMH3ml52NH6DgDrMzTc5Vr+b4DZwGh6WlhmO4BLR3k17xIkRgR0GQb6StZ
mK3ohNmGYlwI5MpkvFIMFvYuja2+fzPhHcEp2ibfiqhiVVcDJwzkmxmz61nV/cS7jVt+R2r4d/BX
B1PJ5rvZJMHyFrOYbya1Rd92HhpMe9ByOfEniPSoqe07YOV6AtFIRCLfG8eEpdFRS2vJAu945BpH
Em+iwxez1bn8ZY2czNrLdzD3AuJ6y0ER8fc7FzMaD5cTieWUZsyoh2IPn6sbi02ZF1MgxDUT6Ioh
WV5JCbitKTR++HexkXY6Y6YYJMt0NIt4yzTgVfZhC+OYFyx7t2pzm9EQ4yoKb4lgXGk2pDBkVHHR
FIsTi9L3WsZsDmp8xDMeER3M4Ud2pN31HgntZXSy4Q6AyReCVncyo/XnQLPzVylwBw+0rQmpK//8
FHj3S+suO/jxf82BPKEQS+f+lOcS05dkP95Ab0cSCvAopad0V6QVmdbwbrDsOuq62WWN8w+UQUdp
Eph2xbA7USKzObgj7PjlpOehECMamMm0MH+sPXonoHm8jwUCR69D8OWiC3syaNv1KF5rzEVEqSBQ
lpF6M+vu2iZEcljQtkiyIHchoUigPPF/hqritCP/WWPLnnBnjwyKCUuUTnph9GA2LaphET8bw9RH
IyhZWWyLFK25nfLdE6mR/14Xwmq1Q0nI2apMDc+Cmf4iC6xb/zywHyuASFPbAvxhO8AcoAQOauwV
xrtRDXp8rXZpmMPrIVfInD5K31MGEsXLkTcAJ+D5HMMyE4nI2WvbjvEvuRCVtKVxLjxjRzRTmkEI
aqQkh7OrrR+e5l+Vz7QrCL8dJIFMx6EJ/0JXpUQmMvmeCaDfIubBHC5YR8vPspjUgUHWXBrKvSkf
Zy1y/dkrFYuhVmmlo9r8OQcX+HU4OD5ErP9EOhf2oOd2nRdm3WcJBQsTBhlnXVRN/g22itvtQ7fS
keroKRbQAazXSTizWh5f/R2WF/xur8aaQfu87xZjHYRR007RRHAaONModFPLIqKAlwwUNQ1KBwR5
tcYAydD9j3P+Kk1FJTbODA6A3qdMDgHCri5lCrRhSMt9DfiqWxfnF3pJwMjUkJsqN5N8Rg5TW03A
52q15VJ+lZuFdYXyDrkPAfd/8qiyR4r+dmVl9+Hax5dgxDYjVYbD8rKwvtDwdwwtQ+xEKImTuY4y
+QQ4Jp9ImK7jVVlSl+ibeddVjd4SHaniAnxJqsYnDCPQCiN2oxhfV7QlcgQ4Njerlj622bPVAsBE
ojj+M7DwPaDE8yOn13xwRmzYwUv0Qf7zyCRFT4lJ70oEEgpoQniN5qcTwcwLsGBbRRRZH1Aq6Cq7
w0LNbiblABLgMMYFWFbkrWPmYs43KLa6TcSu4xJu5EjAKISj2zj44W9m56kRkqZY4vuLuJVpOyrd
oKN6xuAGLTauNY4UHxmHVmkDyfhQIMEKDKOmrf3ROW1DvgqpTzF/65TEKhwYbv3tHpuANBWCZ2B0
TcZbsz8yRO/ktQNLeRWtiv0zUPCAEV1KN6NZBfBOYmB1KTqAGIM2IiAK1tItroihI0kIIB3Vz0Ka
BKAzXecEa9c5wXxVwPFjpAXyK9JcKsibZCiUInLLFjYBLC+35IUfiiugdswk4jZ9YI380QcufVaL
zI8k3lp3kCzS8RzN6lpmxOgX76K2k5OBgoq/y7viTE/M9C0JS8EdHSrdqaBxdLUxtdRUHwYzOQ2o
ZaDjXRZ/vPgJP6Ja6clRB+IptD8ST4QM+JDigfxt3LAzoT5FAtBHWszBXbvQ8yvDJi1IIx0Ky3/Q
swzZpPpTAD7tonAE9X62rtKLLuuLX/I8dpAovvTZaVHJ4MNVqvUTjgzQ+8NHmDEnGnedifhJpPCq
PNb6whFFPSjaGCRjXDgHSDSlVuOMQqtIxc52WVo2TWVZ9klw/CQAaiOwDe3temJz36TmJlQcEFlD
pXr7uxsDlfb4tNLyDdaQZhrcsOCgiau+En/iecQgoPxTCaJik5ad1l4rfLGkOPPSZOjIZgGMJdcN
iFNGeO+rOR+FXJg0NifUlcq5l8PymAxAqRGPdoX7gWVKo9ZaLv4qxs8vrwzQbR2gu6F/MJeJOLD+
8Kx9gLZIbQmtHCqzmB1GGn2Gb6zuINopUY2hR3oX+mBFUoL5L7rrudRuE//6cYXkn7RxrJbgh1rz
vrwYt6JABOmGO9/wmOmVDbhe3FL+uYG6hKdexdklw2+C/N2rtCW2JuYniN3Aiu2RahS5hU9H9fPV
Z+HDVP12wx4aZ6/wEHshKaOdJM0hWUfwyDxCMSu4mJnNjfRxXhOVYNp78BSoE7QMHQe1ebfTc99z
7/bp0eJCJMzmlLWwqiBnzWZGO+u6vd+jq5t8SaaHqBQpHAfxwc05QSClrDYOqvgLsZjEl7RI4EqK
A/nGZyXYcmaLWgfXVGC6bfohn7GfttgQKcJAzukuBNADa4LnuDKH8WtcG/g2ALvQQ6igXdQ2MQTs
JkG17y/CBT8RGPm+BG+27R3qzo4x0p98HFsMPdE+PAPyBiYRnnZ64ou4x4NuMjmsSBhw23nauQmK
DrI/2Y4AU7fFx3dqYnTm9jXn9DwcPBb8WJGe2Ex4Jaut/NyhcXUkFwyY3H55mVYgEBepg4/sKUWO
RTTQEi/EcTJom2rigC0iFNN4hZao3Dwsubh0aIBfi/dfAh1hUUHmh5yVOa5wPh0Dng6vitFJPu5x
4ZjK8Z6UEgKZV8KipI5PTIDlGMDuA0ukTCXCTa5qmm50VJh1l1bN7xzwLCEDtD2MUQsBCjFcAc09
h8NAoy4+JFQ8hPmkWL8N8JECDEkauX/6QD8Rp9xkoWKu9B5SigxO+hB0prx4hN2uwFUq5fc1SxkZ
qjPOF9iwZDWopBan/EsvnQRWWd+6pmsIiM3jb62lEDEqLHfcu1JDKL3nMmt2yxLR+NZwdLe3lxKy
ZhvB9S1wTtDe7KIZYnpfHIETsOhpAZqKTgKr7OWVA+4UOz/n156tLxZJfiB1SpUI+CZCAgQf6gZF
ndQMDd07ZH/P7cCVbHd43H5uHGLGFcnmvR+Nrj+Lav4B+YzFjRJ7jdrr6IxpVn0p9aifzrXxrEgF
vf/N19dLqukfdB9XHOVYlHTGaGE388k/gzPwuz2QHGAs1rgESOwPyJgYSRcFpG2c3jPQl7YnumC5
StfhSsQJ4XHWWQ0jxevCeLmlm+hKUa5gRD6A8csTgCn7K/BZTe1a7d+veD0II0p1F/O8F92R7F+a
OwNGGJcMvWAImX7zhC5CQShd9Jljth5Q8xOMV9VIO17mZW/ihPnGL53FSOH2A5mgRYBkbiijIIFw
gHpdTP58yvGHJNj8t3l2+WIfcLuP6HPlLWTqZxshRg7NS/vjP6eg7Ff+SbHBV2R7cbqs4h4SENEo
YIoscvSh08q2ZtBN3087uP+8TNQMKQ8SGgpQ+i65YhDFHLv0OLTh0kCFoWPuJEBbdLHjkD2sSzor
ma/M161SX0hBmEKhs81zeaAvsOal6kztjTHrVu5cCoGiqDEpwCOpT2QQqor7/e0EH7m2/KXGUWsy
ja1+cRzqQTq+Rzciqq8uVSdtNCQm1RlmxlYPRW2Oor8LEBEJWCQtkhgTwhaCMtSykqXJD1/z0ZKo
H9pNFlmysV+//HPniahLM3IiXjNfrdBcoPPYlZ4GrBDCJCAR/Hdp3Hf2qyCxtbLWLOonMPNN441K
7WOLrMXOD36+HG0/O4AXl/pCeCC3Tucr3Gbxa8QMYUJJoXr98AaaG8SfjDdZLYJArcRObjk2riFU
WIjofP9tcHFDi4t5RrQKF8RnfjClimmfmOX5DGN+++0pxQzRXYRYU07O/99mNREbcCl6G81XSvbI
RByUuZNL0XrXx87dh2QzNaZl4wqoOU+UjAB5Zs84WDnbVpql3sCEwdRvk39xS+2VK0MkfaiTTy3r
iwHll2BgSfi4tA+hYsBVC+HtSVab7yMp/Nw0WaJRngwLljdQnMa60/RPS9QV9jW+KvZchUKDsVI5
Hjg4QoTnVKcO0+dda24Hfb+r3Domeh04QMwUjBzRnraZagBprXI534h6TJRvC28llZeJ8+ATv8av
53LGSiBrCt4XoAEMxElhdEyY22Q4uCpqq2Y8mVP8B6nMCwxhjW7ZckXovWY6prKxbh7VwnB17YH+
/LCB0Jr60oKNLKzy0+s2eb4Z2j9uUp2KiWtVpN4bJo0mdMNlHQWnl4rpxdVc8q+qLApwZXM4qah4
+BYhgkKNdvKVYGfT77GMpieLCBZeaVT6YMfq6fcM5qKR/5E0zD1++qcTO7bz3rvxzRf020zaATwG
1AXkobHkrmVchNGb4s5O6tKegbK3Q1A9k5pTMv4dBI5QG2qWNkwwuWTAcY/7O2MgRdGGGObAxCBj
0ZLte1+Q9F77IzLjxr/AwdX7pXHWTtRic+1bKF/NQnIa/tkeA6ce+D/2JooDbi51M0ue3RtXhocG
12y9ijj5wKlm91m4sjnb8LjlhU0j+63fSIZT4QiguQbvlVhdC7PsOZjEnZm3EqJgD0cOYaXNKhqv
CW0cfUm0PWH10EH/HC8pcwEKik5bCZD6ghBrRlnLRvGh5wXaxv2gd5SnDaWzoe6AiyPMXmTmIo2J
bWnReMYYkiPzwPKFq0tBHCAmWEKT0Dq6FwjFNeT0VOKahbaJMx/YIClOKhTkCYLo9Y7/EddLq5EY
JCqFTuhR4mUOaljvFVM1KbADPNP3KVaidmlcmha1SccCfNp8gmolBscQmxj/qPa3Q/Flf7w+GNhd
/3X+ZQSLZ1SLuMWflACINXugsMCY5yWXDQtSL/nCdCGhVgObW5Wj2SO25IMXAIdRWSYsAXm1otuc
Te0EUFBcYY+pqqdFZ4cuRiEaR2bmDxp8wCHkmJJi3OpMl5RMVhEZ2e5v7PpLV4F1IcjpCYNaDsji
NtOYC7FNpElsv+Sg4v802h+mDJITybwGH1MPnDNy89prJ+SLZGOjmFgLlcmsd0YDQ/53z6nRlI+R
9Qe97Ecb7FcVnWhi3ACjAYNWfiycrzw4nNOPilW+UI33qN007XqVMZadYdhn5cjhjitvpAUTNkda
7N3VnNf/K8LFNOor40/homBS3vZ8NeUm6Bckv3OSygfa4Og0MRU/LEqpf/7ajkxdVzL7fY/bqrDR
WbqQvcoUaLSUTVEKuwNLwA0ULnSKw5q9OLAC9KUtvBCLFaFbynB1Q+wfuxGdYqzrnD23fAd0g3Gf
4Z6btf+JomR1qaecZIgLFj+pxTbTsnqAAm/YGS2M+2Jq5bQJegOs8QFEZa6+BJVGRTM/YIXIKBBB
cEQVCex/aa5+82DIQ2l7CLceGFJNFa5Juch+RO1IrLTIQpSOHVt/5RHP2BvbijUbb65gHyonv2o/
khF2BShXAHAlymQAVTN9GD6cwhVnmMBJ9rljrH591HpN/S4zkHTzwU2RAxuzFR/S0XGj9J9Byly0
LLECPvZjL/j9wldhtO7mGqyXX7AsxhvM0kGwzoawLX0HfJA997UeR9BWvd4RT4Qu51EoEBDedao3
0abPXgSi2sjo1BkQMtGNCiGM0rXBhCTrnbP0GLNtjaV1hrPhbBKZZiS12cMYfjpIg53m7AY22f/N
Xcgt3AIXQyWNzV05xU+9IcRxA+IuGyFgbEb6X3LtyP5IpTmIOTmSx9GEHHfB8zMHLjevCOZEzfKb
AII73+dIv6FejpDSN7i5umi0w4GldxsAzx0pOAwMs/ZvC8DHv/L8xxxblyvD9NWJCgfyJW2WDFvF
DaS/Ko6w6aROF18oklAmrd+dizOF+96p3mzWKxASbQaeT6qRn9jKJrtybUj+Jc9Hy615lnI8etPO
wX/Wv/Sg2AQEH5hPG96EkVQNFXQa5Ldw4b3c0FiB/WwcV+of0qryu4r6xRh6aVrjSvo5Vez+ZSBi
xmG2gJZ7g3xD8aWXxMo9phPIa8q9O4U58OapeetZ3uV892NUZywryl+sZUuMq7OXxkLdUNe9LwpE
3oGi4v+cBH7LEOUsoxoYSVynwZGk0URN4Xy9Fj3pJpVgYLbiEFJIfFlMPdzeyx/AYYur831iPA6i
42el0XfRHQ53/xLEaJqmRp+Q9aGzohR+HzTvXeNJAXIgzCImicPudy1bkyfFWvoVICyENy3uAX8T
3qbwms0XZDOSUnTjgnUn3Uhh9P6LkQ/n+6she80nkjCSnwolXNhWg1Ron01XB6Mt+UN9ym5Byukx
cniQGlqjfvT6kAJK5XrPS3L1/hNX8YV/xiRgTaPZxj8NxvBrBB89qvgx7YZ+2TJ+YmNZ/jgWyZQ+
ZK9ecgI4U6QBrwazgSnT4+34Z3JudDE9ai1Df6QE7rJBMxn91x/qd9h33CPPKBdyGPD4d1GqPByC
h4yHBVrkWbaQzsx90tDzy97MFxsi05SQg4yp5DP6YDCh+Z9ob+1SlxHiJCGS/nu+/OIi0DcTLWdW
RWULafIz+PTHSrRmRAC1dI/6pHIcssXfefiADKy+4b9RJkaeLe/WakArRUxLcfzByKWOpGtI/+Za
IpQC6HlB1/M7YsquoqfQFgiZnwxUfUJS2WE1mXSHjbfQHdt0h2aiwNhg+LeismWKaRGhCuS3EUc1
SSKqxTJmSqhhbTCjUbMQl1ijW5/cHZoKr4UIfI+M0A8V0ifmlhclaKsQC2amepzUN8pmvzr52PFP
B9p3O9mxYY7lGczPSUzCbs1qz/5r7rSHsQ/VmkRSffigvVyDBop0czqAvWRnze7Gu7AOT5b2Ay6U
XsIrybhppq8mFuMEgoeA5v01LEa/9IxONN4I7nhJPnmQ7lE890ZyyOzwy8vMRKXK61O1B7dgQ4Ys
EyCD/dL0+Xed8q53RdCrn+rHzx04Vn1kDHWrELlx7ibZ7oaoNrfh+UJxbIWhIxKXBPQR77DBWQr+
1jUIAqbkTOlXjQxKRau6d1utGqd1AafDcxxF//XNNrMwGMbBW/VO6P6J4dHmJav+hYPIyE1b5d2d
/DR8EHWC+K5VJ8ZwF6otbm5RZQ57eMIP1l7artU616iyUxYpatfKdlHiycO993HPk3hgCAJJ8YiI
+KG7lvVh3YvISmx8HZWKyJO6V8etw92hJZ+sAqfkhmJr9RHKXbrw0GEw0r/wodwOuFHGzvq0PFJi
qW+Hi5f10MbRg3lC0SoVXDHFtkqeNymOELajok25jO5MzgmFrn/kHTldc6vewGYqtD4+BaqOMzD8
WI3/tlEByzrXrf/IJGnaq12Q2uvVifTkiwH3uG4Klj2nVLI4Qscm9agStZu2pa23h0DQ9q4JtmUV
pQ4RIyNou8PUWrvlB6OrFGrfRFmwGxL7/CJE83ONCNIzN4Qtn2/eBlY+CVDjuAoaeVQpdZt6P27y
J2TjQBRDFPKZy+CG01knIhluDDaTHli4hY9DOfckkoyZ17UVm+8HJEGOHMTnOTQ9jepBgN+eBp+3
qfn5SVJlFaq6Y8AJ5Txp378dSN1QHqy3XLJlarrg/deAvWlAzKEWz8oszihKzCUG82HztNSmC5Dj
0uMtN90N3cW6MA3QkjU1fBI16CZU4PH4VPCBBMyQStHlfhqEAtT0d4GrCLhecLKLMOT73KVvEmiG
/7C6H3oCz4idEfjHjsq7VElpGM+mv6h0enZXNdcg0oClbR3DjdRHG7Px25jg4JzRwBZwEIPith6r
JZERYGV5LtJUHPDBafTf0UzWcT+VL8ZGdtf4bel5hyjBmei8NJ2faVg7EF4GVW8LPjvZCCuV85XH
oIZgKBiGIHy2QXbKTQ7rzvrcYPYoQePRHK+lkEvzb+kWSXoMV9xvJESiiH7GzDHxIeqeHlJ9g9Wn
D877NLZsXzng3iZKbUAF1Ob/BYrczDqMe+Woc/rC+XK4e66as/lk9sCgof+i/wrvHb/SayLoM6X0
8XNF9SrPPspRQOzvyjS8LotSbeJ7GEfQWglVusaHcHVmy3jWqW1/Ld8kjzeOKvgbnChIB74N9H5e
6TCZbZvGJqCMw7TK3nIppNVbwnze1Uky8pGVRgbKes/to9wkw5RHIMXr32cZlQ4QGa66yiV7FHNX
ihq2Zv6CMXdI9/5KuA2cRdEdYlvegxDGaro/y15qEfzCsGPBy+u50J/HIQsXJCAAwy8SJ8YMXlvt
9dkFjkWpwqxrxtKtcnzexPYKA0ocl72I04R+0lnGPt5S4JHDiFYzw6DGzl8QIQlIyXaFqIZM9cqc
zM/ikKX9R5nwZuFUHo1ZjdMPBHW04BeBIfUWIZj4OCRuLZGw25DKcishVShrZbqb61wL3cuzjmz9
BSO1EhcyV1myDOWpizlIH1NF09NgeH40XC+p2iyNz18k93qSsGX8rxCthF6969E5l9u40VcvwRVY
PQmwguyJ6Jzaj6W1bl4UVYP5aHIWVgAauH6AhIHlZcwGgarqn6V52sXp24+OnmNRiykvVVSlQnLQ
GQVj9b4haer6NElhtacjb6RrQ5dJYbkicp3vAVOVEMZvY/eBG+YBDeZGjgaFA32xok7tdk0SbBMn
nfdnSpLeOg8jpVnxRJv/HaGHTlLmC0AvWB2gzT6V87Z8pkaLDlEikCEITu9e9sSaYeG2glfzInL3
+xRpu8t3+vYs13cr2Xz4m+Y9vvzL3EMwLu++jdrIo9JqRM2+WwnuWfYSidkMdZschEHlH8dpPX8A
SCDA9ZyGD++NEMheARXyopbtcxp1T9VHCQMmj4QD2rBS8xKp6ADpYwBNsorqTQyc1UV9VjPEcHz2
iJUgieuTa2+3fwinDQO8g03Czn7hsuSO9hzFJFtTCJb8n6Ktop5z+ICVWhRBne9ctWaprY8jFkOp
0zS9ZuIucVRGZM1docUepWUBinjA0Prver309HQ6vbJu8ZvBWtwXoqj7DCEUuN0f+Wh/YwNzKXAV
fofUdLlVrGpp0jyhtlCK6swg0pJahu1Wmk62gejEgI22F/ah1wfTlvAbrph93m7ppyEu1x3O4+q+
m2AYv10GVy4tkEzSrK5IAQnpPoWMzUzJRtwB4IF60Rc+L7dEY2kcLNQKEBb5uSJfMqokBy3XNT6v
Z351NFK7AAYjp4Ha0hmk+UnXS3sbUicN7Wu9QJv6DM6cSRv5ikP7qrMXwwowZHQ9zwtc0vDyQ/Zw
iWJsISm9oAi2elOLZDe3KVyPEKeaJdLev54w2bO5Yc+f7t0ePjPfhLu/CR1P74IA+xBOEhYH/0Gb
QfJh2FDF1HyoSx4yGV0oZoV8j3amiMafe4qvYqkS+GjF+nHrrUpCMbWM0v4yVid7CAIMbOWiS5OB
apxCpSPFX6K0fvFsvdMc/hwaihI2FtN387bXK5U5aN0Mlx7GXsY/R9YBqI+T94cQGJx+Kr7hyTpw
QeZxWWcKwLR0O1v/ocX4ZmPHtW8VCkT5PvHp3oyOzVYPo54U+sBUfBSZ6VXIocYzUBxlZN/ePHes
gHjAM3c/Y9u3ex/hnXg7M0abgddP7kA4ZGitxptrJ5N3ieAZ2qdBOMRdIUQG4riAys5FEECvlyYf
ralkJ6ELkYjn2v73seR/iFiIsp3Z9wxTdC3+XOZeDE5qolQ6hfhBXby3xwAtjU+eObPs6H9Fhv3F
9A+OkSFdSdENF9inIvsxolNe4MXZjtPSZIA0Am1jn/CWH98g9M4D7m5L0YVRFGAwjd78N9YsUfPT
ncpqizwv7yfmyL+wovXKHGXoMvB5K+XpVsVV0D0q2JEm9LkpYYG1bG7X4PN/ah5YvdKEYAW4kwT/
mhqHRDGFM24rdRL73DdCmL/wHUBRjzLHfr+X1NtBNwrtQBYGKFWkGLYao6KrhvMsHBxlhVzMMsPt
7ph147EgumgQJQvfCJROlyjJALPoJrdR4NgRcJlmjycd4vifQS16USSU5uLktgULG7e3wfgjYygs
0f8oFuhwdOgx278dTbo0DNm1NzyKHWfvgFZMiVFKSGPUEwQQ4zaMc4HDdMg3zj2RVTNdXYLn01fi
RW6A5X/iHQT81+I9Az7p8nw57oekVwtP0QDLhvkm5Wb7c/d8U7z7Sa1w+K9KeRlRtMvuIdIjyV2K
dSQobyApp8JzZFq7XdF67yzgLN5S1N7g6ZnaZE3nxyM8QIvAcWqitLCnQhKZ1j8rHhC6O5P8qPiv
4fDyxyHkiNTNdMb+Bn/gfOCvUFQgVCFlTyiQ7sjON9Yp5/ZVY6HDWZC0bbQtc78hV8Ls84xpM/KL
pCwYXHNXdv+XbsF2lQ/YFhUbBF8N52cRJuP/wB8klHE9WMnULNSnDqSo1i2JO19alkbiYjb9ErwB
EYPEMIUcN1YyhBrW3QTSUVlCsVw5+nPO5RYmJDj88NG8qQ6ecgSqQXx4mLuWhcouqu7PDPh69qPA
H9cIFzk+1D45C4bNXLbE6srZaOdNzG32wf9bsIfz4JQX23XkwwHboJO+chSmuNn9+wYVBS2t9UNY
+PHlaOs9fbw9whbUYdyqGiSCAQAOTAX6ixOmQsubd1zOv+LCFI8UK6HWjFJ7HFnlVhQJOkTWPX9z
I/o01BIYmdFS4HavjmOYUi855BFPzYvPOWmGz4yrzzevtGYPrVCbuHV9AasJl/fZJ12ZqSo1IS+T
ZUlEBGw6YVXnxKgIFtKLF0tKxVIwCJpaFbFbC/PC4VkMokCwm7shsedpG4U1nH0JredzODmwMiLh
5o3rv7zMTgQe30mSq8zZA0JKexIPDRB5aeICaqaIMeUFJKA0Dz0yIXLSVJICsX7lPzee2REtK/yQ
knTEAlmXlnGolAW1Tr3xwHpElKDBpwL0Pp3SwtI7qSAvUl03rdI9kG1A/QUjZX79z/zoaaEKx1ou
Hu/rkRpBuD6KaJ8+QgtKwVY7WjZVMLPnGurzrMlLlZFRfm3ygFvHgW83r5zc0r6QqRBeAkEFZKa8
aoF11BLZEcW2wunHd5bd/tfvevYNdDpHMIoHoVFKS36VPoHuVXBfxvUTPAZv6McqtyWW4FcQrDNl
nurw8zbYxflgLF3yL1ftL8ZXGowhpqdtq/IjZRX4pPXxsXM8VJjJFThpfrWwTz/Qdds6xwIGPHDa
u5Yr3bqkef6I5DstpWG2Kxir18cMiJtDBzCK7tc6EC7vbxT2pbmJvM+77jOmU7Ln/yV9ce8FsJLK
a/g5mspCFYHnlk/r5aPc4VJnJ/3wgrIJRQ35dyPirXF/kmxY1kIfKxgNHePAaV5dJs4ipqDWyLPZ
+w1CHP4aEfO8WNfgkFG9imB9DxzkLwVYVp7Dl32u98jLRiQdup5Yaz6b9BiUw0BPMAO8sO/lQkq1
C1jGSKmYwHxl2zms3VV4v6fz3PFyH21dcQZYQY/oBFz+CwzSpWCa3C5Cyiwn738Ib4Aiqiv1p0i2
uGxGfM0AAW79mWFhDNZHvg881Lr6HalqQko9PWtEY2GWTgqM22NvbfPekvFCvZK2copSN4ZjueVp
GBY7btRLDMafGzIn13jyJtoIE0jCePGuK+sAP7WCYLWhNa4e+/o1Aq/Y+D56Nz6jzVgUMfzEgmy9
V67gaq+CQjkAh+3LX3e4FHwWxHErGYMbSXlNxIeohYGiYMog4dqqffVNLMbGdrDIXVTpBPxPuPtB
UW8BgPzHjGdM6yEasglk5Rwf7BB3jdWNM0pmMO/hIEFRfhDXSax7QMA6cbBr3RqmxG70d2dtOy5Q
CuhS/wdfU7JTAta5Wyf45fb4BtUNukaamR9Q8htxkEr7H2TAnplFuECTjT7cuwhtaKRe/0YcxXbC
l/TjhZz3U0Mee7Kj/dSLSSKV8SMRwuUICJ1jf3oVNSpd/94ICBFjM7qp1QNmHyqfDSqWNm2jqY1l
k+tblu44pQNqg3QgFgQE+bp9VkFRyBU90WUH6+ZRRU0MYL+hWSiJiTRRQaKsxLNPVBOQwi2dbBMM
vZmlwi3Vc96YKGVpr/rr9omrsa7B5uEoT5yhG8DJj91QGhCyCjn8ZpgeNbr4GJBYHH9ffkyvuF3j
r8JXf1BrW34Rh71vjxa+LVxhwpl+rb2PVYoMfUXcRRNvryd1ojiC0VR+8hjq/XICnKNAYrPw8eZk
DuGl2MyZVjkg2zzWNMEKBuW+VMl7FnsedZ3rvMhcqkn6eEe3E/+4aLkci0Bxw5TPUgop2gUoaSLh
tpvcrpwLjhFFV1oa2Q+UAA6f71UIyQLsXJAkOELgksJidrOpBE5cF1dB3+ogfNEmA54OersD0G9l
LkPnvfllNS/VgTv9mSc99xYk0WMl2J/l7KFFSfZgHfmsBJpX8SASaqfJeQHfIYfO0s6FbWBdau04
Jv7q888VplSlJnnE/VtAH2taP4SVvpwa8oRlcuTEqgKYlE4ubB7zJAsGpqTSU3lyuxmj2+HiCJ2b
BaXRW3NkPBqDgADuTTWwC1Ymce9eDv8m5H8m2hOy1MFovFC++5LXyctKHrsPeauLHVDcqNMUUIOw
kLy3WDKp8axbAcOIcNXHRTgQiU9/3kYTKnJkFkBlS2hQ1SOzqdTaH1wa3T72N6MUIOAGgcj6P1Xl
IwtcTSj7bkM0YiAdN9K6+jK6f8TzX17kn+7sscYU1+62yASjipF2fkVIQWshuPk3HAu775wsEX+J
fuzN1DexjlUQn8QY9k2rmlBaQGNbkgH2/WZGZ4HodS192XHKpcOpm74UcsWQ8D8eixTCmNS9AcP0
ZMULWgI6FEo8fYgo4TPVGi0KrMJvQ7F4MjdQbFTzAqyOSCCd2vYtn9LV/e7tVwneNypu2iXVJqyh
EpAlpqlYPRydcA5k9ZYfNXJa1DXoVg+i/60/6PcjwyhUIOCTZ9n9E5gCeOCsir7mQq/Bn+f/5y2e
H+2TlBwdQAUhzn1L7SvuR0TnQPvoeEklzU3S4poxR28HmVkc8duIZ0y8mWThKe0BXX9/wrngEUMI
dIuiaBYwp+cpMAZ5EdOUq2oMrDCv3LVAmooKGtlosXKBVSKWsmiS5a8nhjAQcAU1qvfbvWGSPnia
yP9P/K13zzg0gy6kF7RAeenqHZODIjfJSQY8vNdrKynQ2ulVx1fV3OjvGXFLQbvsNzDN826TXbw+
49DEODTbHRwAHxjKOkTKmwDtNBvCXvVbKa9HpUoe0DncoZRk7fNIlKAPKfkhpaoep5OYtPirdwi6
4BFNqs/3cmdbmS4l3YRoK1tS8pkeZSvCFruh55B9gnyB3/Xvq8ot83TsOWjhueMgCFmc1wbSIT59
fhYHqdMxjtHIbWOzRwCQzKCultpf1k1Ec7jLxpsFSlr/fcwCj6HWvkjnhJpiJuMlTXG8bd7eBdci
BQNqGEWvOcKXLoLiblUjfLJHwj93A+K1prOI6kH/g8KRjy8WsRhc91LD+gM1YHVvdRuaGe2m6WSI
dEogJIlgNFLIGJGaE7asvdQVJMxABfHVpMZtCxy4rtc9U7vFeg5URv/zxQ1aQ4J427aVwtjOoIMo
piUR7qk5LCk3eijUiivJ6qMlzBZhTR7GvYsU0pL7xkfwcELF9ns5hxMe5Gr4ZCAKadNzNjGtXDqp
N9qLqulDjdX3tC+wKfziXBsrcVfxfwdC04+ZorolJkGM5DN0MoqiRaAJaTn7TQ4kYgVZsTLT7Yij
Mhpz5lon4h9gjt4IYIU/ZlkV2xkk1fm6Zc6hejuODJNjvX/Ag4Z4hb/qQ/gUiz/A3jwfa2zGDkeW
B2gwWPLsbJqUUrY8NOaVrOYvp37mK6FDiZRFL/LQ2RnTSgKzq+AyRZ7WLX/t4pzCd1tkyAUA0K8b
w9AthhGriztY4KaLIRBjXy46GRPMnDJCFCt0cXUR6Z89kI7Jm/XDmuwhxBdh5g04SdoH+kWC0Buo
GP5G4y7Cc73fAnKmcmjSVgy/vIOEi5u7TQEkTzw+FG+iPHMKBBz6ntN2SN7JasJG1uU7nYrbMW+j
/dtHoG6zyJQYlUH2NGTXnjNdrPbp52+egmjybNtjWXG/znAFRFkSid/wXbet1/8U+7qTCoDqt/Xi
Cgt4xFrjQ51b8pcKHKjvUdGV2uoWyIQlB1hrlZmlOy+g/VCbVyh1COgixCIgVPZwi9/CMx279f7t
5j7dLZsDHEOMtJa4aMOWVhnJUXxRslKYeXLmLhQdG9BFVtFNOPUyBkzspzdlq3OBvdz6f9e29FU4
OaD2AaeNJvxPKG347EWIGtKBTZeiD0MBHHQFEIG/tC36XgqNX5h+Xsa7s+yjdD33jugwzvSVBWaI
+bU+tqgLje9YtVq6ydKorgWRBWj8RJkmYWPrJVSENlM6YLTuUKmov+DV72vNg9e7rWYz0/vGpIR5
d8Y4qkHyFPlohndeumicyS1Ir1TJECVAe0jp6Pib+/ZZoQMZo8AQaHkRQFJtvI956KuoOVEfGR6m
w+vC+vObl2zFiRw2zJmEoC/JwoGSJ7QuMM9P5G47G1kToe/WrLKJgrCYTVSUB+dIen/kk/DYPE4y
N8fMmDBzPDcsA8BsdInEF+3EBhY2M2xyVOyZSQgwzJrmST0kcopZZ2wQPZPk2Q6gSuSJXSGoYWkr
MjsRd4SsQvJueGJ4QNwZPCtBtxhJ9kqPDtVXdpLJKUi97t0zZ4BhH25JNbEl0mEP0upkg5wO7EGx
VaK45mryUPz9DdxzPADG1+J9s9JCJfMb+tVnjKocKoaYB2gGujTgBTtOj7uVcL9PsW3/5wo+ma0D
BuSQyd44T02IZNsGHKlx9HlU8PwK4DKcWdYw2F8jdc0hvE/Kyu5AFeh/5KnsxqN5wI5CsahzGnQn
cmt0TYxJfQ511wZPtxiPZNrUQ+BAQlXrdUvS4LILkgd7pCGjjCAG8b/fvVfno1aEaNVsrADmO/pf
tZgbNBTtJv/V35Kq8/ge3BjG5Cbj/lrJxkB8L/n0Gvp0OjHnS8m31OscrJdW25Vj6ESEOYC1otLG
tVwtcoWhUZh0HmwxyuWZgPhomoh31cAYkgCgYmuFwqflssvJJUKL/q+LlqwyE6us3goBzZLKdYDo
rmudSutQPx+nwFpkgZ7VQt1zELM796VYAC0fpti0ylPEb9h4ItRnVUL4kSABl4vTEB31h/M77LtQ
mj9C8xaumLlwiXGe2ySQfNijysh00yDdmyrWNXTmsRTR4mauChnlQ6AJEIWlMohPmJAUHsWv5dE4
F2ctkr//FabKG3Mh4ZxxdqGaW72UrP+64kyYqqpK7dcS4vKQzRoJCviDus84v6s+cjCyEVQsByNN
uoplddSbMS2boUmGYZ+jN3TdsXuMhT/T/sDqzEq/ws68AIUdUqQ9DDd8PZjJGlkpkWiSl65THw5s
ho2QFQuTnuQUufzoOmiDS8mE6TBLhWPWBVUd09glJq1wJ3vWoWJoB10U0uRys47I8RXBh2tfYgZ3
WPcRMUeclfb02jI3nMje+tqJHZDsZl1Dy3aWjvoQytrPrp74MRuWDmAVJwzf+NOTf1Lg00hDHPZr
ooMgjW2RNL+rHJPRhS6ZMWZ0oWdsPNvO7jo5vXdUAaE0Wnob0rayZNm8rusdClw2i6UdiuR0tuOT
7eNc7E6HEkHza83AmO+j+93fQk65HG4/TX7pWXeJ48Grr6jiPl3t7YOEbPOZ86zh8Cv1nmEZ2Myo
RjCaV7XCAsWXHyrCO7urj+P0KSR39jiFkxJlycr3TLvvenkravPpmfofFPFYPU+qp+MfwUjutFZj
vQ0YQ0xTYGkvFL/Ek/z/+XLKlJCIYlbeuF60YLKuxmG4GwSk4oXfSGywv7yNQHzgEqGQ/vLMxh6Q
tCbCX+Q+ZHVVVWl7DfdQdxl2lkPDEgf/j6F3c3uFLltktRsTqFVYU/4zm9Eb3fShGdGdQGKUXGts
jTySpOGGtTDZLHpCwkh/uHGntOPrHKZsGP2SoQkqcSQ2Za7sM/xXRYkJ5ohlwig8Pg2mdv8fGd4G
6EsL4M9gnV/CcowUl8WG+GzYhFz1Sw6dTKdrR5AJLSCb0f09P8+M8kn1JaxQKbCxe9+Ji/MvHVgy
gJ+6Hx13wXUxLZfXzbN3ZPfMR3wptM116BTmRHMYDxOLBj+/Mvr4MP+ZbojNVzpMH1BeunSLfXsk
MykrzwuF14LdrTzVWTlU6G+Rj5GpCqrHERCki+yZGTEREiWToH/BIIY6CuPfH8zEBKxq+zJzEfna
KF/5T8jCVuonJhEhrUzmlQAx5iKkEnhUavDjx3WX0t/AS69hM2cVRTLE+ug5F0KYjgDh+N/0mAVc
kiZPDcvfo0Fic3yoQNuwHtf1LkD4KBlFY0hKymcPaTCCeYaMW8t7E8TWyJYQWLJQJfQkk4ImTWMv
QavDQvGS3DJaniWCQ60VPJrd9L6YSzqTEVHeYQPWBLakJocjPNKhx6S+u3KIUuM40NX9i9zcv/P6
7mITpWmslvm+Ne/Xxtsax1BHDVju+i+ttOI8EUrO8DMndsWlULbsh2fmz2Hrc/KCaRVPFwU4Otcu
4/GRw7Uew3BTY71mSHMttsppe5nnGFlZ9c42+VuwkvZhbW59ANhizW4yQazmMRoN2mBl9pmtPcet
0WwLAkMk1XfkxzKhJsgNB3QLrOYoDRFKAFM4SzK0Q+5Kd+kdx24idESh4VWbyHDC3t50K6VYhLXC
WmfctfDptsmjxoUFSR/3tXP4SfiPSWGnt6BiXMQNmQjD5/fqP9SU/ok3lATwAm0uhdKLIy8A4Xao
AzOVgGxTnFw9vLMZEmf6YK5MjNHSi6CP0rqggEa1mtc/laikD6plAvhEQhQYdibyI+J37OaBoPU0
ItsK7Fl8mPb5i53JjdCNOBslakcYjf8MVKdzYKpNXn0O78ICt5aizRz2dP7k6vhwkx3ett+5hEU6
FoKrQY9hVuAslWJOTx0ItwSIy+tpOIGDO8+H4EX6VEcE9UmolYwRztnEb+OU/UuVz93wyRotEopO
css8q0qJnQuTHpDxlJgyweM0CoAvMVNp8y5rvBGx/p8trKk5R45PLHxacRSujPitKCs9LsMN7IsD
0cZDefyHSulYvEAFmhH7I9NraL+d/f8ABJt7uI6+JMbHwuN0bdpQ0u89jWFP1I1e5+bFBG3kG9wG
ozoXQg4c2nuDqQ3Dh6mLjvT/b0U0GaqCUE/fdKUozNsnENYVsLa+NegPggiT6fciIrWpmihp0ENL
9jhFrArudn/2/Uz2rV/AgQ89rdRAGwnZrTM3K1OgGOKUWDfSYgys2jB05Qq7PII02SPKYa4v+Xbw
JsXEcGFer2HCfPE5l0PT3hOl2RZUJrMKZhx+3fdwdZ6e20r/DnzmIfMVTjqsf6LDnTKC/T48u/qz
FMRiBO029uFbRPLvVjvp77d8JTyLDop1nPMh66Bu5MyGxELeda/vTm45qBR342GvfcZpLCSkmY1/
qOkWbFsE6ffFrFn1rZAR1L0cMtmvmHdP/l9BezAkTyOoIyOWltkgmyRuFj5Wks/iBtN4RDclDrca
A+FbnbWpx6R5eOZtTDH0XbiF1OcW5h4t0nW+eZRgrPrfL+gkttHspkdPaR+gqvRXsrZcu/CcKhT6
b+CqQk5CtLWqlVyStDCNFcvinArFcomTYjU+oQ3dN8pxpCO+kWtfcoBW5Ux1W3bJZwoPcVjNPgDP
JY4hEZY+oCLCaOQv0YZtFMx1fonBJx7riimDG6cX/qGBc4W2AHxDfjuhhkinl5QUFk3JcpdTgsl9
jWOuQj6Y130HJ3shYirxP1N0lsJ3XkN41+GloJCSvxioQNino2JXLCa32nwhH2oJ7+NO1oQvCK5G
DmN0BQY8vyg++dBqlAHb6OoZ6PH99hBHGwjrpUQptv1hTgA9Zw1Fn+zMYxf3+f/WzqA8NZ4ahDOm
dgWPvOxaazRgLdxQL6kihcfc25dtJZCNSQ52u2vl0DbH+UFURpZ3QT3Fsgvaahf1pUl1GvfH00em
ggFqdT2pIcCoqsOs6a1SwcBvStMLF2qTiROS+4cCQQQ3wktYH7p7X0+1X4vTNOlbxjotfB0uaKiY
/jKRB4aVCs2Wc5q/VAR/XS2PUckkAV/ma099/lq8NhLnpfZPbWg8P0rxYrSOoBejTD1VcpTGZRz9
uWfjrqlUr8H+sEtD4JuRGCmtFgV8fab/UPQI62vLUZWb2kRVNWDgUthk3b1yvVwg046A3gCKct56
fAMLtZgXHT17cEa01DujXBe38NZCG9LLz4K2G38C31rsQ2HgMZ4NHP5eDL9Bpoex11SUZ/9Ry96Y
XJnIfXOjVYoAThoNfIxDZvhkNK3tNDSNjwkdzgmw6yeveaCpiZqxceUNP5fjNz7AIE8Nuo10sYLv
n3um1VhY0s2AgqNqjlp+pOsYzna1ureUcM9SjDQljjWpFTeJ4T1zmBNILf6tF+kE1HhwjvyAtNaj
3gOO5icAYbUfVkQ360G+3aNzvCdLDC46w0axUec+vupgxu8VrzZJrYspi6BoTad894z3q+2cR+qT
VzcykTSZnlivtA0FDEk+dhbj4YEPVyMNCDYZA56RaUf66Y4ZUq0xF7S4p1ltntd9rArZYyyFgDCZ
Iwbh30DERIjugMLP7IyJpc4UzoV33k80xWnV7J0ObDhUnmgCX3OAryw6Zlj540FihlsmSWV82YUd
H3oFZpTb3cNHFd5Gu/gWgbDwuNk1ITL3Kf5YsLzkkU+ydYRL2cMKloU/IwzsrbKzAq6Ge6sdX8cy
Q+YS2YyMWyuyYGFe2TTY/hyRojBKZv0v+rDXW6/AXzejAzSB/Tp7nHSv+QKIVx1GJ7wVHQs+kduc
8qcowL0JwXqypRUWAZVyUqQOHHhKaOD5VVpcOn6SHVYDCyFFGorGPaZ98/L8NWJhJQHlAv4uH2p4
4rz93ZEPxn4ZYXrtQnYBC1QclY8+weupHKbu/SgcVuuxqAm9EwbYTmFMHbPNKUSSocIS3XpRpma3
Y00t2nusn1EbpO9oWLLIsvEEgUdv/7QyvNFNimLsdOedx6PN6t8JkuNOfAMM4lGzIGgKEWiOOosl
LDy74zUhKhJjnMEunZsAxLBZ/Lh6lhnAeEFIbZ54Vfx9dz32xInxYoosQJv+9G8fSM0HsY5IrfkE
bDgpyMRQPDVXxQJAuMNFt5YzAc+MIxi8cGEkAyeKkGe8dJOMzJvyGw0Jg4Ag3vfEeNxLig3fBzxx
5ZfKo2po1Ynkg4v+gBDOTvwDkfVWlBAjy7sSISNi1GQiTktHDYbK+4eIWdv5Ylm4AbBI8LecGBuI
Z4P9niFMLM0BOnLGp/OCTQ0Kgk5azClDXZTmnX9fwiEgOQTy8VtJlYxFBddnQUtuGYOZPqf46ROQ
gIFp+T/Asvo3iYB5HwyS6L2WdSZ4hudwuZdL5oLpkujJmdfHDdms4ZhlwfHxDLg4ucz2WNXwH2K5
0qV/qR9TWFlkcjXMnelG1Aeh/PPIGj7fkRKLwXr9cxiakY229FVbsCQFioKVOEQttyzLAhF6xcVk
PuMyzF921U9pabtgdEpQLh8SaCX5OsQ5ux/KzqkSFYl+k+tjQ/CSTKmqopVtduOrOe0ddVZUp7sb
pj+ZR7jH67FwLTGqBPMO97uZehYMM7EuqOqDiUOoZ1VyHlLfnTBnrr2QpZyjQbz/dhATidRLXoxN
HEirRYna78kUHfCEqy63hSCxfaOhrALp3/9acgLVwpfwcnVyp5JD5A4zlqvtdvfFc5s6cqunoddX
funqA+yOq388TsCtdEyUGYs/Rbpzh58jg3Wy2ZE0oLjO3cPnzQJBEwYunjmNlC4jp7MVDTy043A7
/cTB0KdoI+URSFOR8F+yLzMyisg11LdhwIe1kjrIgh1E0seYWAZ9YOG7kRCjXWFQ4MqEpvY3jrJ5
re5/oqsWo4Y2Z1vRs2P5wujew61uZulso0KhH+/eCUYIK3VCfzVqWiWdoNNBVK7G+54iq+jvagVX
FyFUk5x8kCx3v0x1cgx7pqSbPjy3s4U7Wh5i+7kkjF3NfbrwhWo8/o1CuGkhjS1jWHBERJRPDvyb
rqrgZeUJeA7rx4SHzvXIzi8Ol4XVA2TR9Gyg98yy68gqjaxxxfMZR/MB+MnZPer+NCbUZSJtScbQ
1dLs0wb7REfRcB+hmDo3gCHb+wEI5c/HlmAK7zyJ0kV7DX8iq6fGXqWD9aGoPTCbOmMsiKv6A6ap
1lxYN4lT4PMUuUuiKIGvNV6rGPxfGveorJVKbk1z4lZWgZM9TQ3NG34MIPmVLn4XIrmVlCvVvGkU
7D9/VBk+jYQIlw5r8zU2u/2n6Dgs9+TvjQa7h2OkhLyjyAViUyuKRjCkMrqWIX0Qmu8WmFP8eut0
bJTfEhUlcDvA6TMlMz66mhRdclxG9lMp8i3jr/534APcG8ybVYQ7gTmKvyVCcfzDdmZPk/LRdrVL
7eTwFaBfRpwHUrVXzeNZZUhu00jyesFneUJg02ffSo9naIL/fEU/EdN8ZjbDlAV06KweYyGlb+qH
V1/Ldy1d5Ofnl96/IGoOrbFsVG8vjCVYOvGgwjO9ETAmmj7I5Ii7L9pEx7kPjnTXpFH9bAvc+o6D
B+bQDq4uPztTCROe7z23xFYeVHZ0KTuFERkzUSovkqdEZg4L3glc7HCIZQbdsgDyXJlukjMeVhEv
oBZgrKWQnEnC4rF/dDT0dIUIoyc3g29xg+cZhFQyQidwCSiMXUuTpKAdRI3vhMPYa+nfxtjOlXE7
E4Bo+pyirk4ngiyMEDtpsoZ7iblAjYHP31I1dIEyD94k2OBnRZBDUx15DFkdbwXjmtQyGJkbk3yF
7R6EU4uXhvWRNsNonbhw147RzKUITaTG/8AxJxUmQznf8THfbIEnKBFCz62c9yNSnstuky7/9uyw
ik8VzvusY5qnoWKuyKRu2S0eSpY4YUXgewgOjiJYXtSLcNi5G2TlIWx+tegYYcAMXEBohVJ8he3s
6g7Ab7jqM4khgUVVcsMsXPf5zBA2IQtkiE5CrOC5dX+lvdfwh5ZPaBzJFZokp2U4gFCTItuzC3UB
4wUZB717L98y1gd1YaAxCjBR0mh/nOuYOW9Rb2EK2Q6JWEXqoHf+agQg9YddvIWtaHodSmCewPnG
aTiNBEn0lS4/Zf/kceRVfuOHv7wQNx7eUgAw9dZPEuaGgLZnyuVifunQGpaOYUs6td+NeYmkCgGb
trfGzx9YbqfkpptY0RBTQiFPjoKjFWZp9iGk2Hxlx+XVOFuzI0EsaaaTdc//YkZICQvdWATu+tB0
GbGkMahuXLvQgpobjxUBUmqj76Vn6UvnGeugKAcPcCTOx1QvYmTGOGtfr6UcEhzDpMupNKpYeVLY
QTrxFzNlMxTH0Me+x2Rcp3YhZS9dXddqYlHQZ/HXPT+JcVqfT3+vFQpsb+CwgJiPpxqH17MXRju7
tPDlOYYXJwLssgKsQdylRgEtSvZXDW5SGt7AeJDRMrowjH3t6b7fPqjFMYd2Y5m8Ez3vc5Nb+gFJ
QA7PEhLw4WrESiDeyhfTNOJX/5q0wUopHuypbcnMoCU0mUF2lEywxUqw2jjSqZISLqi29zQOQ6/U
I6Z8cj7/+OuSOUmk8087la/3TyLiC34XhIzrYUWNr5RLluJcUoiRxJXwpZ9i3I+nU6niuuC5PZj6
hAgnRFXEkX6WtNPsCsQ22clHvwH0roQCbYQtQT/w6eCD9YArekSKv3M0cN3GpatHaKZc651O/oAT
Bjl7vcJcPAjbmq47114xQRGCmohRsK89AB0XjBowh+KJ69WaboYYBOuibwC/Ng6vI8lb5yNJON6X
dG7+PoZgsMf5gAsjHKbhXRnnM07cMF0GA2XKfv0BQZR6vZUv9fhGEd+AdfzzHhLUTr6OFebt5dAL
S1LX11X997ntkce0DWmvj2RuQFDREjiWkLKyd8SrguNHvPW57/jDRLqS3DLueO3MoSG09XIlQpob
3TIZprzzbJYBawLHn947imsf4UTaAAelIJAhIW51AaBQdAgPPRHSfNoHdGSqSrFUNNFRGgAUEGV5
8HNUK0L1lTcyVjJ434C/WtnQ4q3sSLwwXpdgrtr9SnQ6LY2EAWMNrB6u9/tX0i6+wqpnQM/fAxnY
ZltbWErJLKfQQ1kOZ41Nbe7Fv3yEgIBgY6PehA/uBFC6E/USir31k288tKH57sP081mqEhZRWcqv
Qe5vrtkRKX35tVstITY4XpUvUoQqYkRNr2uIAq8Y1r4HXzj14cJlma25GneIhdYXs+XDUxORA9Qt
VJkCNAfRV4Fy1snoDIbz4QsaM/v3FHCtUQRhGuOVwc6tDyY1U6xy5LDxtxGQDNpwnVUUj+aqyuGx
roikkAsNH9mAFiN6/IcsjnWTvjwB2MN3zkHRcT0o/HAMrRycBV/gx0nus/U6Biaya2TZI7EuTV+U
GdOSv2+VSv2FCj0DAsLvoFXE/KBpDPl98Q7uma4cL7xkO9vJWd5VFzDibJgfItTOa/GxLuPMAPkU
BSAhtBv66s1ddIInxqalzglEFzRgk680LEWlUYbb4JjoJF1W9ejMC291geQDD3jOMCPAenbWlZ2n
2fdXN24clbPXp5Qdk3eBf4DAWsJVzSx1aKq7+yDPqtMucTQm0IU4zdE5uQPls4GUaNyzvweFGTMv
O6fsVpw9W0iv7lOwdcF3ENyOsxjOpudMzG1ViVG912eQQESiMkLZXguoY3zXwPH70EC42IuiR9lh
0jn6h37Can+nV/PZy0s8wlaLGPvvlu7rRwh8TWx3I1gDS3VCgnI9twykwsrm3+vHS3bVYiOBLmGy
5SyriPdRl4lpaNct8pRLKO4wWZj1MnKU4HG1ysWRyV5Lc19QAXnF10ldRd25gwCODeDWTbWGfRQo
wNMGmIM+w0QdSh8UD3JnvJA+KAZEk0eBmHM62qEpvOcR9shgGdu4Bnds4SbafaX+/TFZoJiE2J5J
DKMapEM2ekN7luqosgI22Lrp7czcR9tl2s/bFaKmKVf1GnX0bFhjizkdpCWiJpsPb+UqIQi+o4vA
l1npwpzILd354vRI1dXrsvpbecal6BKCVppUkbl5QB93rB3uAJkmDcEn44hDnsUl0OGM9cqny1Br
JYYtEnyueVAa8nolJlr/xaSxxnnbURPDyb5E7qdtfxo0G2G37nx8XB0VxxtuE2C449YJdApyK16z
lrhfsnDNfhb4DVV0DjW2vJGV/qJb2F0e9TLcyo6QnlLzjYuK8mpLrnPg4Po4kulTVm76tLsN4wdj
2cAuAxMa7Sitjuzgf3IZvwqOKL6c88yERu3mB6HBLXYva0z00437J2pe3IrOUsUdgYWH+PBhMTX9
M4GKLtIwNL7T3/Vv1KH9BgLw/PC1ln5SOHk3JQCKdzf5kfH9We/a9KpFbeocRhPxD+WNIbdtDB7X
elB2Gjpu4u1hg9Uvn2GztHxa392CHQfdGkTE60cevF0NQ858iM2o4MRCziW+d5MiTxQ8s9fz7JWZ
fRWTeKhb5ZMtKO06FibGpA65AzqX+RKs5Qc+pT31+9IkUNEBw2XfJdfee42F0yHgoYiYnaJexO+n
pKp5IOtd9HvonrAzDNm9Z7tGRJJ2/lOWmNgOaoMc0C2xkkTLK3IeG9PKldvDzo48/eYTtdsjIlE3
cwnMOFNNZTZKcJl6Dr3PV0ysinkEgMmprEvn9M3uwhBrm9Q5vTYlYldqTT92OufCXahTEivSsMew
0az2YSHKKy1KrALnwdxd/yE5JVh/uxBp71n9k/wfGF6pNzNpfm19ZUaSAW1SB8/lJ7mFS6NTSHgp
Z/8OIkQe0pxHdciaIpPxZjJ4+GMw5bpDhBklVbQbWSXYdv7uzmTroBimwDch2v2fOuQMrA/tgZ9Q
LD7nX/5s9MfENAkw2D2JGKvhKT20gUxY/l9t5zxygY+A1m6+c6Ppe/ndbdVBeoxR7wyiR+NdX90z
jiLyfX/KNkTNHDbQ2pMdQ5lhtgsHmzTWXwXfnNM0beCksRjSgk9Hw5tDbbDlVyRgp8LKqcR/r71H
3BPoF+20HDQfHKfisJCXlZvOv1KkbZsbEEtk51Ew5naVKOSzhe0vJTD3zpOkfXzaZsMU5VO+jDfM
ItWBWS7kVDW/3G5XSf0A6XZPt1kdhHT7hhLfkLycjwtPdFjdE+OR4IbcpDpRf9C+rHHGs9IAAD9q
Mfx1WclUloA2rAs2qy0zI2hVePOAFGKgcJPqx/anMxgdkxliA6Ddkx9Inq4RcZdNl19u0jYvo55/
uyY/z1fAqR8Mjl11Lu8STe36G6FdkKI2glNNIiE747DA5MrP9/EqLoIqJPod3NNCsknXVrJhYbPn
wlK1Z1kCfOWMRjgEtroBk2qyBn85uRZkeXn93nh2YYzZt5B2ZN54L64XjJDRxYCh+nl96oHmImKx
AIcVXYWZnhROvFficWdsOJuuereq2OXBxylx7iG+jPg9gArbI3D0uMNDjMEOzWiDdT9whMjMLqBM
wCdzLtVNJV9TVYNO5rt0btyOyY9FR6gAh/Q2DXnZ/f61vKMXwEOLtZK/6mYiTT8z/Wkbny3X67WO
5NXk4ndVxpdHG/UoGaIPxv/ypBnHOBFs1blmvqWcpJknVw79FLdyiCcn2njzPwmVXz3fYu0bFC99
Jnc6ZM5njKoqZYX/f0ZEAB9cWyTfyWCEvH+M7aN/Q0X+aOdSrIWpSpA1mHBOG+7n1ZgO4pnZacLK
9WH6hHFCPX2fEqcPEdiJcXg3QEVpfm0sCXk/kZVWSvnkGFa86I+n0hM/Rhljb83sz+Tk3su+lOcr
Y0gezOf5DIpywMwk2/htxmpURVHR24yt+Y7SorNVjV6dt8DZm6WXtw9CDyQRQfmpTZLINYc7OXjO
V2OmsQ45KX6O2MVitQNBE2w6t/xDjwW3Kz7fYssMWaH6rdaPua5CzMbR2CNyyyawdy6efd5Q9yh6
AtAUiHjB7nxq14DJQzJ5DkRIBf87wxjyg/w68n+HpVyfTjWtq9YsJl7Kq3xRTFjOfC1O1UpTV5RC
M6qvTvva5WvX6KgAhA8eGbkf25KizW/W4iaox+SWIlk6lc4brJjitj87TRmT85xiJb61vkYmxqtu
JgjVUzulROz1m3+1NrnJMBYMsj65mZf+9epyhFqr/0gPkbZgmP4AzG25vPhxdEHC4JhD1edEfbQR
9W0cY5qWdi7UBSMCVOawvk0ThZ8m3QTg6wVEQKEx785ys1wmyL3FhFChZYozqWhl6CXWxi93Bv43
/dJ2iRDYAKCx7pOJPlb95DKCcwBx0BFMijWVFOJ9c3d88NfnHWVmtfUfoOn0hb+n43BTTCIzs45U
VmiR9Y7oPUdwi0pWbDHg3gEQyoPU8fRyctL4+m1v3s0UWE2uhgvVSQHtSXWo0N5RhTSVHk+zqURG
d65BRjLarabKPN4Rml5CYw5h9VojDZCbIji55q7BvRN4W9mO9TcQro17LQwv4pw1drsYSZO4H5/P
boTnSqVwKR8xNWsTQfqp5Gna025w6uPJ7kagtBXpmMjEtmQ63+TkiwVuibR9JxMTv+WyHH6bdX52
ocynMxHC1g8a+4HCGCm0k6V+9dIJVgGiE723gV1Acm8KYxbWeVW7kKVQSmljlkWRH2jrELNepv5S
CTwX/KVjXPY6aEtlPlctF+p5d4NJpbceP848VrFuKJ9Ira0eNAk6Xwy8DxtB37aCCwLId6i3uWsw
X71yqQu1g8U4ssxS8n7xcsGTO75prtoDfc/Z88W7iEZUliFaJkNQyksokeHal2JgbzijPx4R+3k/
8JLqaypL0oR3vNAaFEcRrxQHwATbjzmkUILkSAcoXDhdqTZxBuW6KSjgmhkMBqcosZNHASpnKWA2
CEzI44js1ytEyiAtFsioocPYKCX1S2p6kGeuFhCCr1YwZcIPLE7lkUH+THE4pFVkNrMnJmojc3by
WQOJaLQipkrY/QDKBh5kqyk02pJ8BdTY6pHtoVwbooCB++WeWhRigw/cg78uEvTKYxX9TaWGWvLh
y6H8mOczDsNNLyu20awkEn5pEczZJtAmTRpVl/4pm+FML5hv/sUTec8qCh9HX99xl+xd2cFqET7t
KSNje8d+roml9KGJe4BhJZ3gW0EvvGHBY8CnqIqMKtsyhThLUUmq3wf+ckEirCYcuOPMvtFktOr/
CjvRzd8jt/2/isJHYr8xpKiAM1XJIdXaH2O7k+NVRyQYsXLzZVgc8Hcqkhu9u7WlrWq+CPWqsF6S
YC3iRusp7dGfxWKy6XdqOMLx8u5Kq+xLp8Q3/VnFcLQ9yIIHDOvHdI20NUlKmey8ksBj7GCfRtDX
PuAnTtr8kFmbX96x5gjmPlB9pz3uEhx32YvUAKc1RroWjs1+QJyrJqFcl65i3TNWLtot5ppuBMph
UC+U0Tn8s1m1DBdZ4lzMP65cGrxyWpCf0kGdMgnR6Mow+iPMo8px023auXurVuLYT4TE1vQJeNBA
EWmWcSxgGdhwltadogzeEk+w7k+mPVXxX/j9fxUbiR0P+u/uHGtAK9nlL7gjlN/U8pqZybOur2CR
mV5FO5x9rwyJP0l1avzI+nYIFx1/LJKJqhLmWWOdVIC+nzi+jXbeZ/nUT/wHP/UY6jJCoT7Qsgiq
rX6kAc7lqvKDhj8EYGDQKDPGUcmY/9k1FvvEZzrxFvUoxQJNG+QHwfhvwoSgZVNZ8axjzasgZJkv
8c9nmkbhOQFgUC951bqKaUXKHq9J1ZC5kjXyrqHi11pHKv0uSENntoEUcbuJr4BUp7sOxlKFFAQf
XGi3AoBHeMdLrD+ofLdrdT8VUCp4n+nDpTbdRrV/VIsL3XCZA/FJT2tq3n1x8lialyo4OI3j1Ntw
pFiCnNDjybGn9tujNMAzXyU+MHBdFILfGBk5lz1WZCkguTW2v7BYVZw/8OcvX/wQPGiUGJbbdf1u
uh2dJCSLRhiTd2VPYle8Y21fIBWEI6vVHqyWh6ykNfxvfnpSQzduIpWlkxZ3H+Dgi7Ey/ilu+c58
IpO4UD/jEUH9nZPk8/5laUUaVD7vXm7Q+tB1K1NC4GbTHinZnhrrijdaxAvCpFA1CKPtQu/WPS3N
X9uaE09xYI79Bs1KA61k3o7gcGhP5kAlBVdnrJfATB/wm8gXvq6lfXQu3k1sPcJqc0ivxePpHvJY
/QCayHjRVJlv7uZjAWRCKeRFRO3d0oyh5yEibHmtqHAdoI+ccYOjwaHSQxIy1uq5wo33bbxV98/N
UMD81DhAu6YhKZmS0KvZkh+Gp3FyxA6Yh09IMDdC7hmuIQ2TtAnsA/AszI7Y5omALlHLO/ITD1HR
8Tf41BswhJ92jJErhC7ImFqKa9yiv3RCVUc6k54EJXgtx0J7jzIIAQnOCvRtlsyOTl1W96HNrIkE
XfFhISZjp+tXQoPolQmBI5DPm+3UwW1Q2yR5zNdD3b6tReJKYq65HO8CAMO01baWudpKuOtNpivM
CLOxE1PTcwzoMFC/JOjkdJRcSyEf+mnl8+T7SwmCqzpHa2dB3CKKwqyx2Vtt2CpzzgKmsmR18vtS
HnVljcRgI9X608lFEiTTAI0foZ2M/mSyGr9Br9fbR+lCWf0VBWwxR6h4/k6a5CNGDJ5hV5X6uVwT
YS6rcRSDyZPCVHKZSd3/jvdhsok25TDx8o19Ngojrj/YqnHxsOSW6Q0/lM4mTeB32Ne77g7P5HVf
IXagat4yNJFxS3V0t6P5K9JajJ3Zh8iWMcTv4oKjY6qwozSLurty+9qoja9k5xdGDH07gRBawJb3
TGs9YcQ7ZBnZocC3WzTQE6wbo/9ceZmRdSPLmtQjrH4pr7kDnBbwTzNQmYz/Hbw2HIWsFyn2TLAR
zchbrAqXmUgwrncOWG2Y+8WxssQlbAxDdE/1brQ+hVlb8vW0Quv/ycydj+0GixOvRxpYgFOUNGEa
w2uk0nc4Vr14e/EZu9wPcA5S95w0j9rSMv3o73PrBKae3lPvOTqqbQuFacnHpi2X/6ytaTeNaecX
VHuNvlG+/L2XOKO3DwuSKqxgfraRi6ma+UM16MgVgPRNwSmWaxQxeb2p7vt3zY+9vBj6mrrGlORT
YqJjEdtu/Rx6ptEQTHcwKLdafmJ8QhIuYYBlkuKzsyKpt7qcOxp4IZr2AbbTxpv7WFu2sy2D7QIQ
HooqlEC8lLAwT63obE81c4Bejlu3f9brzmmWJC3J1KDHYhegdWg83iP7pBPpQfIAt/xf4OdEh+CR
g16WsIbJwAxkhbCXq+HcZ9qv5qkV8s8yH6Xc62pDiqLx6rmzDslzirMFOJV+G0+SuO0Gz+0+cMYk
UKpxV8Qt+LmMolmgxtoPhJfAtY/NZh7eqA38Is6MbanPXPyD0BKwX1xWr8jcVhspcp18DVxQzh0I
DVXpUZErq65xkPs55fWWh+eqZ5HN6LA2RaaYIrZFP+qQhOKVCobMhFsosGCp2AiA0wuUeTjw05iR
wQm9Q+1hC7+DZfxdmZa5sxABxR16SHczPq0ZXrdNBiq8jqguLo5OXVRkYAM1Mm8XWXFgwegIv1XG
4VpIxrTwGM04ppkXqWhjduqSB7Tr1TVntdRrSU5EZIIkZ0idjsWHLkei5Bomvtem8sryIDw/yBvq
w/SdUn7lDpHbSudber11MWNP/Gbc8/EPZmaiiMhH+kM/gZ+sG/Sgl2D/QCEOtQAFzHi6+GD5RMw7
09/yowumhGnYG6OxEjGof8kTrouuZtmTp7ZMEnH4GQUoEE3dfY3vsP4IkG9NScRHa9Gty16JH5iA
ctOK8p1x/mxnEM6D8mSi3cWZOyrUlr4vfesclsAnvlYp3b0eaSzZyO0hB40qksPD4eINi/iEsV0c
kvXWGV0uYMDtO+S1yYdmckk6t1Dh61Y1OMr8eS5WiYzZcyIH0832haTrviNc95G86rhmB1PV3ord
jnmx8TBkh1pxr7z6lT567TUh/bIVf3R1McLafPmhoJ8skemo5WxWbEEPf0hiv14sM7R0LKuaKxAZ
du/ISZirlv4d+qml8IJT8yeGryeCSzHwrLBfEcfCJ5Ny8czGBe3UEQdjeeCOV1+bQV+X3myb8BPl
gMj1jf0oD7TSC7IjIl5HWlc1QGcDS9H513kv3tg49Q55mfR9wxPXHilo/Vpy7FutGVGPFxZ0dknt
YDOXuhBaMIfDe+3e3uz2KOWZ+fw4YKf5oTKOrcChPPWbk9cd5Ts8JV847JdjvOZoK2h3bmHQ5K+w
binxly3jMuTuIF2tU3VFnoU6B6K/DUEcGDE2sNY6IoVCca9xgmIsvWzU/g9Upav0zm2UJl7V8bZV
jr3AMt5KjDFzgg+0pM7xNOFao2CJl1USqsX0zBhcQXXhIqYMJhdfO+3ZS07PJ8srqK97UX6aBVse
ofAietG90m1CAr7g2jINMtB8KJbByTTTjXmBX7gIb/1gVD+460w9S9BtVhR2cDHNClB2CtM9A35l
ugtKvt1VxIEQZuXpH34EOVdGQyEkdLX43/DmOqq2gFJ/HYz00l4p2Z4Wp0CeVr7qXsR1xyQEJ8iF
Zg0tE51Kv31xKVSy5k6J5YEbc30K9q5vLgL0J4A8J2Sg/U8msv7RBkLK5q1UINnfAacnyQGj7U0c
yfKimjybgulBAa/hKrLZ5PEAbCZnfkUrvg66Zxyp0wfeaX/+pOOSIaPazycFwzTnpNyRZOq7RmYm
PbsILCvVaNk34LTVtwaQMUsMQ6nQXJk5niMkxe+TfH6X1C/WMq2dsg5XAqQiDIdCIy4lsMBBtNCR
/yWUmJ5T2d4w35U8abc5QEPuEclb2aEMT3o6+fVUOpIXZ+IXAwBiCowVRknBpPEMigyx1IKfMjkf
Zv4PUPyTt0GWk/8nVBqtT/IpdqA9azP9DygOU67yMg0ecKtFFNmLbAC84dAahaKon2DICXWsLO6u
phg3ZlcJ6NOOmtipEnnBMgCTP7SkcRm76ckqRGc3KAKkH9F+4mvxnrOGzEeCkLL/ReNGaEYNOskF
af2svwxk0nYreKgsTUIB8e0XfyXzG3EIn+aPjYexbhe+pFjwh5LdM1B8DfvHoNTqa1oD4HpG7aS8
sdu0ZGV1rK/pkDQtkwsBt0aMYwoegbQXQaPilAl7MDhYAnmhXZlHK6r4B/CbzyuJ0e+vZcN9O9rI
e4c3N73bYTNQ6cgF40TMwSx9ZOYi+PmMmdJ5eRiJSrCEU8LelDf39IpqXeV128q2cH1bQT9Zz6RA
PrYUSs8CUmfwQSDX/WKUjiD3ijmpIb5AX7eWuSHdIcO81sRIPD8xni44HxFKuYv0yg+5IAXC7knk
kHe51PZEHIhbWUzBwgTX6HK+rzCftvMMLqNpdBoLNbeSbXr7dpdKF4BN9obrm1rGuoUTeNfeOwaK
QL22XU0Eb/rVYo8W2SH2QtveDd/RZ5uss/9vtsWvWuHnhy3iLQc2Ia+w0Eaf4rAbem37TVGmytyr
1VDdTLcZPy+RIoJKWx5PFwvJlQ9w+uynHZOkx298tuT2ejyBOkvK2Z9x+Ql+fo72TL2reBRjGwoW
m2A660MoDWvLyWSjKjfQ8jYZk3a6ZHB/vh8avdwL1MJF7R2WvQa2mIt5rQtA61uxIy94CzJEX45x
FRRJLKwLqnpih1p1tFmS16khpt1Tyun8L9N/yeWU5ypMZflgT86eeSGHw9a1U2ydSPxFMPJdpK0A
36mj98h8jjHK9b8U1EuZFzMX+2gGz8H41i5XFVBjYqXIqjMaM9GvNmsnnLrKSZSz2rYKFB/GNo8j
4bSVRIJKy09jxUKBp1SSZdwjbybUZrLRl5eKcAbAjuQifXc7Uj5qOIe4pRU46dkZGFLvHG7RVeWN
ah8k8TxmbrtsIijYPX6cxGYGJW3+qkbIggnD9/0HjgV7TydI6FtQUPkwY+Dj4KkDkvBORi1zYd1d
JdZqL9o+VUi3JQC75zVDN3kYJ55pmdcj+fcke/chy47S0e0cRYni61IDoTxqiHL4VMAB7ON2U304
38kds5fAnzacjZqfvJK7TRMe7UcUvWgmkUiFXxGtmXNlgMSHb3ouBtW7Ptq2KK/D43BVkC3zquuf
iTcElaHqxif/dp9LySVUbb1UHjgbyvbFXkVdIR5FJPGIkHO7V8E5LMHYT7TpDqbR7jcTboBCMvsH
TuV6KxIJ7n8ThjMAAh9ZkTdErkkYu3iY+m0x29Bftz1wAzpvdpEHLirqjx00Hk755MJlWuhAS7hO
nMHXDotJUA0SXm2Ncra7i0mGnefc9Oc/iUpa8xTe9KqC+fzf07cFdGvWUf1YKObCDD5lNd450PYm
r0CWEesCUIhLwB07hXKYyFgLysg+MB2VIEiGwdDVIrQCBGToRpWUq+qrLWFy946K2MJZhZ/nP+8E
rZ/lmZHyGuUPPiQVBORm/xguYKzhr6QJ3YXBlr07dVk3uEOGLdg1zXdCoW3hZa5cOrzGuHkJUKow
Wqu8AUhHaoZ4KZUL8mvfGHyz4b/6ji/d8PEj9SC4JzOpw3Z98N8Ssp0gX4CzY3CcOyBtAdpjjk83
+9xwOamxpn5B0UoO+FIspCvWLNJTOxuaqYaAUKquzhWHsMhM6NX4O5/BNPu90WfeE9cnx0aSdOWo
gD8SHpe3wdadPLmV6cbnQc5Dva6h7XyXgVh6G7N5Xl/Z9tehamrJgyB7AP9RD1kjwY9ZOyS2KaF6
254jxPyTujodsL4Lfj51AJR+bERewEHUv1snOxrsJ83kmbraNTH1XpEZpIMrFcBwJn4VZ7gfpqcz
ir3CazZDfS/FCXnwkFtqQTdpu6tiY8rIaIeFSbUqbLDd1VTVXeZ/7AnXPun3Wiwb1ONFAkud9wh4
F7V+pbx8Ql1LhYwYDiykKEDK04hIf1dDwRoofE5p0yoDFR3NjGGEmMalU6vL07hr7xFlJI7GHguM
8VjkrKL3K/H6w/Oybjw1Olbjm9lAv+w9mxnXkROEIKNrD+TRMgIoMBrUd5Pc0DXC9tROzEgi4xHE
w3B60BMe/DbbXT2VtqC/ncNzSgYN1vwYlBiejDCycu6HYkPDr6QNe7otovGP57Bfw7gUTmS/mhpU
P7M8+cnvudkfaQHxzDj5ce3Gyly5v4tceMLSkRihG4gFC+pylaEDbIbMirxkoIHVJJAYKZ8gv5Cz
W0+qj6ZYJNZPk5bk2/s1w0jtmdlmAmtj1yXJEGOkwr27aCjLkSVJU2TOQaoy8JfF4neL+97Pxajb
SnuLWdoB0VuoMLSsPdgf/KisDDbyKGqN1YhfGTiPA25MkBtxNRnopBkGM/0Ud0PqAhQFgPyIaCJX
v4dnMYhvMwy1LtIB7UXQs7lLnMOCdvw8XOpBrsgxzWk4gp5RQrufglSnYl52rrP3af6As7edY+R1
ASHuo7c7iEI7KRaJGCiitOFhXu7vRhm5LwzLE8dbfAmgiTlpdVSX7gUsamdN+Yr0VrfpJFfd+R+V
jSL3ih9JATc8TQC4pZbxi5n+RYiN3brf20YRtNocXjaPvvPTTS8YyUbeKdnWkHNgch2ERqBzljKJ
g69XYvJAz7r6IImHKpsV2hDGLlsZAtPGwd9jUh3CSSBx7t5QXtuzZTM4Ty6zwc/zhbLU8xiXzMUU
W/xdbXvtu6pDHJDENe4IHe56iKU3w+9KNQ+bHy1FGe0/2WdKKM9QbnVfxMc6GB3LQR4l97553+JN
c1O/bCfEKZQtQY1D9WcVzCxdVn2+g15StTcKlohhyH93s04jK63ETlG38ih3kbBRnry6FUFQa1HI
jvIxduBUkSBTHSrrBhLq7obV+cLJvkuGOwInunHG8VsY6tqGc2N57qfCOkf6/7OCo/IpRaIDvUuv
DWr2OsI1XOJvF3m6+pkUlr3Ne2MWwphPaRPTBG4801onvTJvHQRNjv9poKOzXksqIqDRpMm9Stmb
1sHh5lhXpq7319+7igUnk9nkh2JyfT7HDUJ+O9QAyW2M7WkTeDMuceMKgZgYYGdsRSIfdRfEO6yY
yL53W9rfxuK6IJXchE4hyIOb0WD19B4cUDYqMh3agNnS1Db4hNqaCtDmbjINH7NzbUW8W8BCYX0Z
pqEKu2toZCeekUqyTWM1fF3UZto3EygUNtXMC4BsxIKFGosxbu/A3cCQK0zs+RY17Qq4Co/ALTOe
/PuTlw/S+t3E2Vlxm++lJ/lXFk48aGWvOn1jRF3dj5ocuX7Vag+PMnVa3569rZrnf0cvFQRYBUFc
HP3mE7BWAKUcapVPdLO7zno8zGaLp+2fnVk2b8s9dT4PtehoUaDnlFkslBIkPMn5xsmfjLshoTNP
Ed1jCnjb/Bat4RnhoGETUy4ZDy7pKU+tjNJlWALuyZwFWbGwSbMSn4VcKOcMmuPEIHa4YAu2Heuj
fiTjvE3C5e7zTFjD0IcTIioyXYtofUcJUhAhn3fNjSFgbmS934dQ88r5D0FCA55E8O3a8E0HVw6Q
4rcls/KR/6jiFMwYFUip6nKouox82B/xdtk/quD7GqHklk1HmionYyF0RMgE5vdHTmRZvTr+Wig/
6NnCvbZ8O8A2Nqz6oGxJyQB+1eexmiCnRsCo2WHBjQE/vQdbcackVz9P+hCuxqW/oGcAaBGEIf/3
9BlDCxPSSizMA1CW+6l/xq3mB1s2iVfOqDcBaFjgmf9DwWBHAtgBBGIpeDq9j8qf/BDKbcQqVj9H
s9ViW6bAE+nW6m3/2TFHSp/vWtL6afqjLPV0y+0WuYgUzmYoaw76y8XNts+aE4q00Pl8z+GsNlai
Ze964ovl0VWeYztdwPsWVzGXtLaD0j8x0OA63dww/5nzQIrxsTF3DU/9cOnrXyAsHJqttC/hkiCw
7aGq7I1GE9yt+jtPChsxbF4i+HFiCIcUZVGimkfdYaEyQFpPpneUNdd1LSIJCokup/FDLpGQNUJG
rmn25AEwTTp3iirIbPxODbKxyNJyekIA54UlIHP/biIs7Yhip1I8OQm6qd22EAgU6YNtoiHQO0Vn
CkZOuoUJABsClLjpzvvs7WRgdP9+qUGXH/QjmlI+Z4Unw+oQ6GbSvQUnwCVnRY3SS5Wt2I7Ub8Jx
G7q4zNZX/iYyBEBrA7xjuMGCDZXfgbpAOGSEva+2kJmKPCzB9j6gqhYSUmv0eB+QSIuvA0VYO2hc
w8xlN6rMO5imaz0Icsfkt1Gsk5RJuF08YDXj8NQUATwWfEJ3+P2eZ2U6cLq7VIUWpSyCXammGO0E
8HnNULxQ4VQVFkpFSlXMjd2QcnVw+bkAQyqBI8wNkFx04J6XHVAfGFwEPbjZioKoMbsFa8PRo3/S
dmuP8gMYHLdG9HjeKRGA1TtUSHDxSkdfFQPdy0nyzudHlKT/KmSJgGPM7WqcY8B5mTn67yIjPiGG
el9FINRydOY51PLC3Mqi++Rk0oxrz51H4YG5oaZYvCUUvoN/NtjlPjfF62HqRkjloJ1xJOgxzh4/
KB8s5OW0p2NBs2nRpdPCGM9VoGaRajG16rcHzukzfHICBx7RGblxKhvl6yhy0CKXcZaghHvW4qRF
lpofzRte/HpNSNI8ykkyxuO1OozGBAZ9lGHtKNyIUeZpIAwgjnCVAAVdrygxY7bc6kUBZb25soxr
BUXVPTJcuIwmTtX0fmX0GkqFSRL+ZOxaJbPnrd3Chcjufd3r0Bcz2r5YiFFsS96jfZo2cMfoOtof
Ymtp/w+ilfvyaON79JKja6Bv+DSPEPDkLHtlGMrODAMf/Xi9ZkY6/chSW7ZY1KH3OLgveR4OuD0r
UYOyW9xId9ZvVlDKHpLQ7TDICTYlj8CrM2aDh1dHZSnjJGQLgVPx+cR615/qrJRu0PBMZOihK1dV
rSAW3533X7wLU5i2O1CNMVmOjEzl0uH5z7Psm7GsXQfDqN6QRN1Zr14vUSPAX9+0EPkdIGEJnCb5
iLMUlgYROQTz3MB8ENqL0dihcqMGQWmKiqrYAAU4NJaArRWxyPdTdMSAzm1k2D8dJCCWDINxFokW
c2vpUg8BfJpJyJBcznTyRQg6cuT79wDXvuPAditE4TeSyKJ6XU3LuUqGMImdpLhNsTOVcv4dY6kg
vFGtU6oSTOT2TuhjUvvAgYvYUBiUUSPETrQaYQ+Y8VSOK2L3zwJPG2wJB8VD8Y0vXLFJciofH2Z+
gBdCvon88l8MKSIksK8ONNzRFDGeH9arpKoG4KyzHUlrA/4Gr+8GNdtazNDviCa7D6PJDFVNjOgw
ixWbxqaXe4MaPI91y/VXISVO1JgHFjPeAwVM6zKP5ow+LM1nnsZAHYQL01yl18poGLmZpgWgYj+V
hbxja2QcbyfDnEs9RUYFh2QZoVWN60tabPD25Ttt8+2jTWKfDNEgLfLRFKL+Vjg9NXz7MtzeI42x
ADgHm25M3IWWhKSywbMvxNojxNJKzG5TDGeXFJRSduYrSy8vEqaXwq8z5wX45TMskheep4C8n3A7
H4xTtcA+7v/UzXWFeRvRCbKAaPk1k8moSXC08jwntN81DTkBgFiGpAE6vbuze79k4SFIJtdkisyP
9hmBGgye82EFkyyDhs9Y0PzSH8jq77Bx1ZTE1R5eY8LaReUG9n5jpiNln0nuo4mHZVzNzGmpZ42B
goBo2WwtJ85h/7v9Y9X3Z4bfYnA0DyqnR9CbG+5e+wjXhF7xPqB0QHjSHG1esblRn63hPaN3t82c
naUHJJDwNt23B/xWlC7AhF6D1r/m/1umASXkmve9gbpB1r8tkCPeuxPUr8plrshyKNXNZg6cpm1N
zZ4SbTlvsBheN+0No5tB9JY3nv2b/B9sj7ZSqTLizvKNmgJ38MpIJApzO1tS9yfuPImZKbLJQEDu
5fXYyJsYs8tsaaarNFFDLy05fJiJh926lsNz1S4fsTIKJ1JHGlY66vPCPEu7eQAJ6Kxg14mOZFPm
V8ydBAgl9yNUMMJ7+F2Au4a3sEQchrO2UJz7A7vN+2Xsd0b1p07kLk6/30aRyJDljXiNzEqcyE5U
gKE9tzJmJOAgBxydv8vv28z+DrjxZF/WkHmf/W4sRdctIvYmfPZcovCnrfPqd4W/rsRkHlb1w8wR
G7ObJDVBF8uHZ3pVUWssCc4VhQVLZLtz9/uVwMLVt4SYKEfMA7p+ctArMg7udtSBhEd/R9HAdQUJ
7hoMBhT0EkYuVlrwg4kDP/vaivn6BgNTkWWCJze5uugKUOGMIrD7AtE1vrap8398rNQzzD77eShT
7F5CtNkuxvCTIKqB0NLstco5JzT5JAm3q95fxj7mXcjfnZWImRfW/ePGUrh8XBLLixxOK3qzNRsC
spQAc/eUFh4MspkoJ5PSBaamdIdBr2NpGYH+AMdUTJeBM4W/+iX8SlXJoL3yXl1lMtVYDqc3gfts
ze3fdrfjqa83rTnEQBJzH0SjgKD/vgS5819HT08u4CJhOAcd27mhF5WgUWaOJJ5TarKOhdW3W2Xu
OCG0N9SJBIuERrgfgCxDu2kTREo0i15F5pZfSufePWRBbNTLwpvtkNrW0ZQxHUskp6JUQdKXJb+a
3nSbNX4LJX0HyCBFnUbSV8fCPtfUU0X0Oam4CrQeNumbXPaEO2spBTKgX8BRke67iz25IgxZPupn
YpmcMXK8d4OBKBPsJOGOnvLbbsaBfKBF5KTUDUBMMNq7rD3IlF+E5ABbOdozKfkAaqYOjvIPO7Ws
D/GnMDnFaRkvRkr2QeKZuBXm4Ets1IahvV1mmxsddfVK1PRaOGwqaZdxQuhPuUUqR8lbHZsRhzh3
GsawMMkswD5oPTm4F5VA5RbhUEsd2Exqs6UGZr4ZUT16qe++NsBMvtWj99e9sDNUWP+019qhIdRP
zNogLKVQfcVJN4hdepnr5VFwWxuHCIvP5j26c5OHB+UqfkKRcYw5ojNJxktZHX533YQVk1FkS52c
cCN3gDJXPwk6S5gtNk4uNX2PqaGrrt+5gaeqwkSlL7amYn31Qks3IaBbNuOwb0L/zc8YuLqMMUGo
vTUxK1HC+04Fqq97GrkTejTQpxg216m17B0BGHkpifZxAcIOb39qUTmWAUWIwo/72I43VSjPQ4Zh
eXjBkkELbRE0lbWdTpVetsDaosWKvhuPcIeOgqL6wRDd+1k1efJ65Xtw2QqjLVwuYWP2NpzlK3bf
PMijMgIL/+U/HDlRdRHMAbNPmt4Wo01ml/HJL+/sCr7Dv/iX9CMyiN55C0extiE1KkDqEJsdqGvY
6mfBHYpwMTSvHcOUJn56jlQn+YeO9NpICMyH5kI+PLp819ikR7ZeCsIbVv/h37l6tU2dw6b2OyQT
ZIsLVQ3A5jWLpSsM6v6TseGeYtDJBrluh6HekcGIvLmLUPfmfLerV/V/YaEl6K89aKYxQTnjCPkX
+kafrClHHXGUuqQxGo+yJiW5/n9CxhXZLcOH/Y6eKbwrebgIdX9iEprQCm5kL0NKcocHCKS/gZtq
kMwGtarRA2WX3c83KP0qpzBJYMCEk9pijkItRMRTGX+V/7H5oucvLOyO556SvWh5zEIlgCzTzABc
8rGelzWBAbhJz+YIhAPnRCRBAvo/cpW75Dfvl9pyO/q9JC0bELaM4hTB0pCKwxP/6gqPlDkteBxF
wlOCBjzhqmCkPV/wyajqUF7rqlUYO18dk4lToLnRpKJzUxkyFXxKpV0skqCVsTSTcQi1a+SedbJT
wXOTM0u5TXesH/OAQM1pFNOODZYoU3jDc/IuOvFwK5x9KIC/KLii6YfQoSXRj8d82+wHlZGrNNiM
NaXpR7f9OCza1yhlj8DMWP69AKEsl04Tc1mREFrcAm2d0l4G2RXc6CXIn3/Z7MdIJpnyma8ZnQaU
g7QNKb8EqXT2cU653cqNl18haby4H/3OdN2NmXrex9xnn0OATVpLvMSOJab/8qvEP5J01fEfKTva
cST4JiUdt2hOptTn9hKkF/tOx4EAIR2P6+W/YSgP9x1oAZQaEiWTd5jkE504iHpDfIxnU82FG8Po
lJoZ+pPhiDSM9OBlNHVtYUzfaBNjkEXxs77AtzcR1NrCV5Iby+AF5iHwltYjSy/P/yGAgPRr/YVR
rlVXj+tsE97BQcpnQHxmOEpbQquzCepe600/vlhi1Zi4cgTJ4sdaMqIKjx2dO37ZzczwSeSbbzZ3
mBdR7Ba696Re2flQgmVIV1pJ/jdlAubvdveIVO8yh24roaOUCKNdd+EiRBvkuVP/+B5tZaUEpkfz
gNGWaIWKbgE/BB6nbPpnN/Ukc6xTgK47jEzfu2KxmldTVcMWmDW2rNzPOFrRZ2Muny8lHwC+aV6+
+tpc3KSpmEaGhOnx78vMiDrJ2WeJ8JiBWo9C+bI1GEv8ZKVUT3+CZQ4Tf8SBAXyJJ4Bz5NKx2MT6
bVcZaq2cg/587UMC7w258SjMH1MwFN0bV/iEvNJYVXA5Ivu632y/jVNhgQE4YU4lR6n0I4iswjJ5
RYF+ui6o5ztWoGVlmkNKK2DSHHeA85Kv19mchihLqtbOu3Phc2t0I01v0alkrN3SgM3m+sEpHXVR
6u+lubhOsvsx91TIZgP9qLi2DpI5+WGzbFjbsbdzNFxwugSV9zgnjbLuIRRzMMnmSanj7u+IW1Nw
b/Um3HaddazeCyZ5pciEseeL2eg/EsWYGaf6bBG+4KchxxrjDsaiy3+RRhhV0Fq4VjrRihq7r3MR
ZSoKwUj+ONs4mxTW8+E760wWljgqFWOgun0H5ydcoKMIYc5DBVWMXhoe32C5UNiB8Oui6DtYbHaW
NE/IP5FhD+g0aZjBhvb2GDgdAALAqe3BtnBbKHlzh/PEt3qGp/ZalVeW+rdS3NvTnDw8npYESGt5
nJbUy0JrY0VH1oDnDGBR93dpb7siBxw5yxBe5tcSznJeVx2KrliOQ9H3yqVAO1cuk00gVldY0vEt
0pCeMxPdda1ScxOyZxE1M5tQlS1SbtTob7kZwIXgoAUhggFdT2zhTyYWD0KsnFRxw0r4+UhyfNBa
gR0kJ5F/LXMJWdhND7T0McdTvdAizW93pVAOZ+C9zRku6BItxdeMUwizctd1TIuBpRecC/mO431w
IHH+3aRDqaws6GLr3XPO+QbyYWmxVwqlgPzfvFmJo+cUj+UuH05U2uU9UaB7BweO4UFvEVUd9ftn
jW5o/GvHtSfe8bM7MOMLVYSTAZk+EDTAEIduSu+YSDDWvuq0YZbBDF2YvN3AgdZ6WNz427lQj8PL
4IzY1CTtQWS9yT053Hzhsr2dRxgQD3Q5zmP1MFsbzJ1bON4ki2CHvgFSuTpSAZkech46N2ZlQbhe
At03DxJlel9I9wcDnWWBGyv9jQEkCOlAbdcuGAllj1Ao351CX9W3UimSr6OtdjTnGlL8slXfv4md
2e2A1EKByFqsDcHpLB5sGboQCPnB/eV0MnhAHMGLZBO30UDzrnRsh7CkYupyWefb8Z7J3RLGIkf2
nqK2xu9BKm8beazsVydUt4Zs0oJsu2askwEE/nl/4sgXEi+gD0DckQemxQF3E5GKCJOfkTGvHqfb
qgpBGTrEVJTlGfZBcJUATRNUUKWTDva+fsf7w5+0QvHifdgimdmNjK5nPhbHMflEyOnrLZ0r9aZO
CqUs6R9U9aHrvjgJBKXmVAY7+y4Es9+4yVNjoeW0BNz3m5kCyh0m2wqalqd18SEZLsdcCDtzHRDA
ZtWB/fqN73D1+Gm4WGi50XYPr8w4JNRKTs4ivCgg5sTKhDOj67OmrhL9Za7ebrbsx50gFY4OHIt8
7FkcwqVOv5+uXpLEVZ13xXJNf6if59j2kiVTAfcTrdYWfcR1WIguZmQ3oUxhdwLqlhle5uQuJC+0
iptwCRdEzR2xj9zPj2JGMIH9VkwsPZehG6PD825Pwyuc2rNxES9C2NIkGik6v73bGpXBnU5pMjAv
gKezQMqMSxXoyUXVr+cNFBlcLeH44tFrJ+KCAf93UybSEpeECBAh2mZWV5TlMXsyNw4MZLBjJhfz
ip9r1zjleGTcSqkpCTesK6adyF0VNju1Fmqmg9nSf4nI98yih+4Oy3VPT1hSvWZUQxy3DdTZq/qB
aEbJXEcxojmYKqvfOTP2bTuC/HgkV7aFo58DwMSoSzfi0X7CfMUXjPuGvfrzX/V86/POY+HMjtSZ
tyFXCw/AmWegMsR26nvhraBJ+qoKs8TV/6Yv2KDV4vn8XszS18vcZp32GWmv6tqQEPVdfp6k3bZM
dUOWz2805yhCH+9Cwg+AOIwi9ktDlIYKkn/RdO6sNJgb19To8CCrXxSc71YSSdXHTUFE6aSttoXX
lSYLexBT9OPo/nXn969BvYbU72zyuCgNIXqRTugnMNEtfWMaOmVVLRxkLC1WssDKpPoEx0/bQD4N
NS0AXject75Eenrn50wiTc1f5Z7uiTa8GXEYxV5wJuiwsCOAmmrt/rzmlWUIqwnVOJcwDblHz+BY
0Q4muQarTuLw/nQq6vQQNSiughlfYaS0aUaBEcAqTfdJHrEA0QTgY0F/S1HrrDeDyu26o69WQjqb
+O8yDpGNBrUKuQkwF6brS6XstYlIOKMkffAamoFZq4+GILOAbXnVRf5GHla/6rFnCdigpsh5IGfV
dM6RVtUZ/tXEm/p0QM5k3K2m0nx+csJvHuwF52Q33dvzkEinZRREQn9CX8OIuxp45qculpTOB3PC
5euRzUsCu2x6mQAlpeBk/Xx+HnT2wDL7N7LAFexmX7unHjZFi2yZ+b5u2Wm0TYYxwEfO83p0JtQl
6KLp5SxbW1WoNXenxVpIYMXRWboXKlGmS3e/aP1XnEjQ9AnxRjddQiqUq6bGWMowVvlEe0p4zHoZ
Pgacu0PANlM75GwBby0WzmQHKAqPppsdutMqpdXveMz5ovXpoAzfLTSFSekuqVL4IdJiVi8bGiDU
T+pu1l3SP8+NrCFnLshXPm4C5iW3fGlfxgFqn+/z9U/pc58NA31bjXQN0+9y2HJWUJsc/ra/YluT
A/UQgB3D3nXpk7w3OLDggbGqFs81uKG4+z/Yptkx0abw1kJ/J11J1+PXbnmx/AtyppvVkzzU2pYl
AFEXL+o/hWFH03sT6iXKcncpaLZeA/wKNnTpCBug6Kj90+4Zmk2BpxdoNLscLq4lzEOeL0Y7zepf
TsIhdyERh/jHJZYPWWDVCd19jPqUnMOJLZ3qFUkNHeS04VlXcagHNb4F/YJr0YbZHj+KznFCkFtf
ksuxCFm46i7gl0gqKdxRrQRYpJitjbX42QXeEtGyUi8MpZSNE05y/V9nrSTjmHVzaxfvsbdRUYL0
vSFQujyWFFU3usaQJDBeE2Y5qAZYX5DIQYZ1omoOKOquiCisFnQIMukQLFMQoHMoYvDWkPqNFfAz
DHSdc81N2R1xMhYnO90QqeZDzw9zmtEA6QvqIy2b7QbL4P1wRVZm3M8ds25utsbs/FWAt9l13Weg
zNfrcNUf+xyF8hw9+28OMCUR9qgWzVrQCXFj0GkMhiH+u5AhgH8IzLa7QLhFpOTV73tSMXyQERUp
3nBLdfIR8ahR0J0/BlFMlyrdWh93eICA7HlYN6SmF++1J4eCboxSgbwI3aKcQUkyGSi2+rFcm4gc
Ls/Q7VqqFF/cFJtE5wFkRxGuHJ4KMLn979LWC/XqvS7mqfF4SllCgaiYHbNd2omWqWW1UWLnHCQT
we1Rqs4etof7vQ1e9Sz/T0nzVGfSoMT4FddwGZNEYrB3j3NzwKrEzNrjK1oFiIbJVjfvE17NDSo9
VoN/GMv1abQJd8yGbFp9z6Q8nEK5X2IhN/KcKWuwSxQgViBb5oX2/6FVSE15H083pz8QlJUtheAD
VW6mmVntg3O6n0kwu+94vsEUx00nlyvRr+/Siolxvh+0MAKNODcwIE0VpUOvZJ/SSuawKk8bu97W
EyU2V1YtD7+0BuNRZU5mvhCqf2dudTzFdDDvc6ugFucArELoSXcAmmf3zV7n1yy01Z+0XvZ+gJgw
lQ3N9kBUX6I1m42pR0cHrg4tHNlnMPon4isnx/LvrwFNUGmQ2BSh/AjGD/gVPTXbxF5bV+5/nfss
jITeu7h6SC8BSomkWlrUC1lND2T5Zww6TJ1Lw+05ME0viAVfuXugq6rvRvf5GruVUzX/zKSadFD6
u6FAePS9/fC0OaaT5jANjejGwbYJt7qetfFB611gp7rSVw/b4QOAr/qY6jqJTa/ZX+aKeo+RG3W5
0rLOlgxEuUPB89IZSFR96EW3D/27iQl00xli+uWCQzGf0Jx1DBVJLInV+tEk5biy2NmIahwSpGOb
wI8Grvtr55pmpS/SyT4xKj4opbGKpDkIBp3Z1DzSf3QFTD3sB8FFgS3stRpOUtJgWysuUHKHI1QA
CbHgdo1J4ULylhyX8JpUOy+YNycZ6QDCO/eeFmmjBmhXRctQZJ05I7LIZPWWHQ8xAC2xuvnAQqvb
P2bQo3Djjqa3TXtyUNsg+FCSpA3LqAYSv7ih5Ma0cF81Xq2TGvgXl90ElZ48m/19y2LyGEu2tyM2
EqBH6jXyAaCa6f8b6b6BhYwFRw0DUalWON9BsbC6RY0hm5QVnmqezq7cvI4/D62q9H+FxM5u/cHL
0oDDxDM4QBfy36i3Ss3g2tNPA0EBizCU9QpT1p80yGfYDrt+Vl16Ny324puWvxVzyhMrc3P4bOfe
vNQyhr6Va+cu+W+4IbfXgOvBJSRfoWmKE0qXzEUh55l9U51yPshv3Jw3yp856c58WYxEpgekuxlK
RgIM8Lg+SKtrbvOAO6RzVKt4RKGREbxa2KaX1EkrZJL5zy3VQtG5bSfDp2nWDUG0eaQ+OhCz6bKn
WSozWcQgkxpFDA5LF7JTtPMKrt/eoIHjYVN45IsB/lJ4CJn3EBk75o/8VjY+XZsZeeLXuyfaKy39
idKLlFIprb76NczQ745w3ATRJPY2r8cJE5h4cw0RXZ1je34VmTDPguCwckpstRN809w7F7uLtRgh
0C4uMq3HThtq6nCrR6oUxrE3fG5bmVJQRZdpLhJTDD6JFpTOcWdR2OP0S70cQVUC2MqFu44rMhy4
7cb353qdk0LV5jntJYRUUUnvcdI8u+HOMpc6YXiML+jUKkYvFxCvsgBzE2ZvqTSLFnld4wT9jE5X
YB6q7hTyc/u2UnYpTbMdfG/ed/6bdAl0Kry0kAwLcbqAcfdGtoSsCjnw2nyNSROurNDf8w6Jwv9x
C+SV2P+RrgSuB68Pb9gb56PSUpNwgN0+e6qF1DArCWF/b2xTlzyxMWQcGF07OFoJrGzyS6OT1HSx
0pLFP/PRWX/Ems5ZXY1wReWRfR1JRlTKMWBAzLx0o39xrYdCr2UEMpFI1ud3QYabvUIRIOgrUzCR
z2nHz2m5KKs3bMqBqPW92X2AfO60o7LNJSpBM4QY4ubaQS4nYalNEeVe1plRTy/Sb/u+xn7o3+lr
5veuEU7xLU/hj26oPyqEttDCTDXa5h5w6Klo4kOSqxwsoYU4HaPeKfXgBSRH6yk//+4UDtgfuFxx
yFmhJs/TMTgjIWTjdc6UnW12oQk2ARrcW6JGmo/RE0dG3nKd0zwD4UBl/pZhUgb0cKxBrFP9JCKi
34Rl0E+5htCzTcSCzQXdqRUPt5wGDPJyI+LwSwzG/U2MHQVkPgviJ8vQL9zsFkSul9CFl7mc0TLV
wV3oe2Li2eCdpiMZkqfcdQOf3e9Y+ELquRRFOS6kKJLLCXzJ61SgixthkilPVHfD9xAFIqBZcz72
VAAccEQ99ZvqtGweBXhdn3XStHWZ+aRETuU5rOy2Y2FKJYRRFGZI6shrkxO6K/YIQAfiPk6LPovc
LikgFmM5ff8QoTzirrFaWibJKatr3/n45ro/2wM89KN9vU9aUnE3jAs2Ti3yI6BArKG6MaKeTDj6
wnwWaMDltYCEhGNflJBouMnvURdcM9ZKiRtSO8M5jQcH25+aqM9eIdYfpTnpwopSXv0/JEV3hlF3
IRbHYtRanuut/E5PQ5MZr02KeNPwTrpen1FB+5ywc45g7rfRwgWmMrMd84lw/h32xUepSklw4ShA
GmOwVFlLpybNCn8p/Xu/d2+H6SBp+AUI21YIw5ZowYvhdhomAa5W4MJJoFSo6pJWItn5Mm6YU5Ez
m2rY44xeApBvTkSIWvR8VWzehu4SbyMSb1DxZzHT5cMkuliKGrSPw5MJ12zjJM7OE4nJY1YgNfz2
PbjN5JthNP6mlmYILgPyLFGxYqG99HRAZVWpPlQCURHotA3vZxlKr33UKWomz2wN6dgsHOKL/8sQ
T31+nR79siDw6hwa0qRzpeAl5+SK3qUVJM+lRuo6BXQEq8G0HKg0XVdHvREJFgqfbLWQkZ3EH0S9
XjOAofRXhZfJxN83nEFPea8IGQdkBCiLjPO5AlDf/Ro/GPM2UWRa6LbwxIf4bVJdsIUEWM5+OHso
MCAOWfrWRiblsPLnbB8Qya/LqXO0qmQZfjT2lbu+lniymG/l1KIpH8rfkFWha6D8PEoOaUufknx0
AVQpxiz1pUKDZ/ajU+Z4dDiDK4F8tX1y+5nHNvFae/zD3CJ3qhKe5bo8JdUShgLf1TNbDQPzldGw
Xy7ikp3tfhSqxeTJuAdU8T7pZkCqzzis2ZOZylQbwex/E7xJjqTXW/MQg/5U4SLqeXWre9IZGWPZ
R3/f6pmnGwpEuwlA2DsnlLhTHUww+5tRwRjna5Z+/xP6gvHLrosdM5g1oERtNFwZJfvy9JoKZgh2
je0DXFoUKbGUBOV/pzN8VFghkJIr0Ktopnfi8EwELk1hkW+FVE1oe/fP+5Ya668T1NfHSr27xkk+
bVso4lD8kllz+0RdHhAYrjjWF7NU19CF4upotM1Fy4alEh+sEoOBWhyb2WjdHwnHOTda5gRbmpmk
rcqy+zVbKrvXcfj77B+vpN6tthufUtwPIVHBoBynrRUSsVOf1lKyqhdRtKvNmZA3GX7VbbnSJ1d9
0f7DXIsahhbicqtktxzHKhWPzu9wMxVAhgHCJPTIZPtN+Igo9F6c0YqFSIA8d9g9OEfd69ogy9il
N/imUmakG40iUmZ5yfgQixBsRbKof6u5Y8VAu9X7DoxaRrlqWHu8O94Jzdf+8C1faYhycg4OJqUU
mHczlVbw0ER+VgUl/wqfQSaSXn8kH3PtGZzp9ziH+R+yRuH6TjYK2ZBuMd6DI5SRNmI1byxVe8Sb
V/n9bW5E4O0B7h9bzm3BBvwtDKFtYBHod8ETgulkhele2wx2eR49F63EXL1/DhOdSx+2M9HfENdI
vThqg2bE4AO+YgqTXijKpIGywIjDk8uXR457H8jqaeJn8hRa6Ip51ZyevbtgWZj133pjXLp4dPrQ
MMnI1H4IVkY++FRSunNVIioKnP98K3fgPyWfxKdHgobP9VRBunpwjFAEbI5nB2DYfxKBP9A8EX7C
q8PR7ms+/ixT28gpGUZBC9EcFQnPXEMBF4EHiB+6A6SpnGOb8tabzjx3u0EwD2inAafr7pbr9oU4
1CGqyKENQWzuaGm7bSEa0mIs1LTfBluCwYhBmIrssM1oUa4XrXlAEBH9XRn05icBo45+mLYepYpI
l5ZacVRI9Ghtgs5wc1+EQlxt03LHQT/irkXMV2pMW0cn16fBVAK97+eh4znWq0CNFQi0FpXl74Ja
G9j9ug5gAX5O8M17mCGGezSLQHbRAnYQ0xf1DxoMQbHCOpW5zWzvlKgevlnd52F5Trx5fy3ckKmU
XsMZCadxLe8u8m7OqlMq+37a4+rD+VSrziMflVM7tDt1bRIOHUUr/SzMsPdYSN1gh1yIkpPs/USn
DjhvZf0QunAecMLFKEQCqJqqDz+WjyRu1M4KahAugWvzoNC8e54th5GbBxqmKVZui/CI2hRBtXEx
udzEWoRCyb+T9QIOXYWuEsds1QXUhvm1BmaUAx/7xY2GO7E4Bg1bZvEejja6dLKTitJa2pv7le2E
m+Q1cmHeupHY3N31UFMR66ZgKEHnfHRXfuqYRVU5Ur3i1pJ1EB9hTFnIghNUbcH4UqoOG1BH4cY8
wyvx0SdiaDTj2pnJtIDM8fDvp5m0j0cDnMnfZjN5x0JraCS3u53ESIkojDuV66ao7IC5z85X31Rc
U1OWjrFM8ZQ/bTUtNb17kYB3NY/LWUbWLp+9UlhR3D/1dbUK+YxkvOlHDQgcOprDCX98q4J69lrX
cEJsYwfrGeXHoCU0qw1bmDw70tVhSVq5oHiR0wKi0oqpsqFnoxfUvuXK2P+wLBmJyngtwaroR6yT
u/I1zD+Cjvly7aFCBUnGtePUEGH+bQzlXKvooBkgnkUgtR5st5+vbA0A5qTf3kdQmnbOE7KhAAO6
3oJ/rzbg/tYy9tCereJ4N0ImYuIvYSTK4W7DaoNpQ8N5mfhLim0RX7p2r7OKKWxVaTBF9qXxkaOi
5XdVFFyUTLqmsJFM6lG9MYJij92afIdXydtI+eWQdUza9b/Yf4BLiSDikefCrqgFe+XCKMGIMPR+
3T2IpmVeoIypP6aftVGYWnTTYoErVLxoxR3+Ct3/UHY4Ty2rLTwEibRLNkMxnyFn0VRn7EnuI/Mp
C6bZf2CEOcEtO1CO7sCPobvv0HoZSK4ArEcovmXGvaNGl2I8SnYaPOqY5/XwsVmSD2uxFF1uvn7v
5clFEpG3Sxz+frcdTA8cCosHEU7SONWajyGs8WlVEAgmGsmQQBmhkbSpkv3BdU9k3Y05kDwv8jwV
XWccfbQdHr4v6SUP28RhNUJhraeQxgFv/a/PprIoUINjTOeDCQasX7q8gUA0rF+U+XpGhZAV5aY7
j5Uaen51PX1GnGZbfqsFz3mEPpYA4g6/0K1ZdrLT6L7RW1Bf3S8mRJLxaxKEB5RPY9MOlBqoqnIO
3vO98UUwKvXJO+GE/c1YvfFAhdD7kLHLwG3aORtQWJ3YFrQEEaGF5/+Hyi8qDPUS3MBIDR1Bt4Xd
1y3GlZOx7IK/ncEh6xki1ai8lE10KyLyKlOFA/PSWU9kLamc/Gm18dGph3faFqErKT59fa2pdRL/
clZGbaV8BLw0PhW7zBTmlDSpxv/mnF2xkodVQGKN5lo1xCc5AEWkIoeAnI7e0riwSzDm11ojJaae
rbvifwwxfd4HnHaOhm4AxW4fGzyMt7dHXwubhXMVP+u/xHm6/WMXvjUPJ/lRtGUglxuJgl8uko8a
Bw4QDHijmG6NwRc3I8ZqPwZxt0Dr7naBjLvxDCCECoyrRBA2HSAd2e94F/zZLTOx2UDebzh5xHPh
keuqYLjm4c1dAhHMShkaRBp+6ebO89z+MMOZH08NMCI5q3y8Do3XIY5Ta02jVp6hgIlPzXJJsMmp
CilQdsHgx4TeUGAqWgBcxlP6f9aGV8Y5mTqlYOuc3ZiXb20KNwjbjof3zjshzjCUu3w17bv/SDpI
f4Jwzqhc5xSrHZQT65uCtW4Mda3ZKM5a2ffoSez65znCDr18S3ieSMFmrZykzEdhsWNvzkd8VSap
EeFsfOQaMFlruLvKJdKjvVd+d13UtND5d2CBPcBnZV2VFdVZyvslAbezeyRLN7Tyb1dCArlEVI3b
tTtJPLPCeZbK/Evp0JZPITrh1Kg2dB4FKDyH3IWT+YmMiwhBJ1qfgO2DTwnjT/+qi7oP3s/sQ2PU
76ij4RBtLdGJVlkTIgpEt5nxdnEbnf1UL+zjsWmfVmMgFNvDWDRI3tYJKm3oH29MBvwKfYs9al97
jtlKatmekoFjiLTpYQA6Qj8fsDvhGYbipxssw4brD3zsA44wcoObBg8IHy5O4mOkHnoovwO2MAJo
Dr/uT2valiGb3HIDs0xM3w9zWZj0ydEQJpmkJ1pZZzwTUrn+XaxUU/PcQoBFIAl4jBTH5HNFZyhm
ODd1Szx1ncn1FN8nKcsOrlgBSqb+LOOIT/KgSAC2JtC+PfhQ+5Xd/F7CavQTtIBCpRFNd/kSH6rj
XuaZlqSUQh5xhjpDmURH8gQBpcgtL5PLKPi+jlpSFBe292WHK2bcU19zwrE7zw526gqOiFsPtFAz
pku7EJc+KKE4PN+Z5TY1wvQdzpI3VDS8OTxMIAUyjVvWjXeV75g+3WiOr9Iic73A7ExE7maF6zPu
F1HjPZXYYXt6RHWpQsPRGBs/2pr0tr+SoanXhM7F7q7BYjKJCYYG714ZTkj4b5jc6PsbWAKyZRDs
DP3nmex4kUMjqaGiRkMaJxk7WicYC7f9WImDjNoFQi34WGViSicYbodkTT73cyUcL64mqwFtAS27
k26gEZXZuEVgwiZV05GQyy7ucObWgJe1J3R6NmBHwPqe9f3FJHSoDZLgoWuJhANIyTD5hyfcn1Ag
/HLsEpS7daaRXTRFceDFRBAld2Xtr9eEXpmJRtTMvlO41qUjKi+XBSB2+aCHWq+JMKuyCBgoFs+n
rDe8Ni2w34CTbNQWtPccLSBFAUgdoaw+l/BbqK3KYl2+lA/T0h1NdvuDb95XMLQG62R6cCbDsJbv
26AHrJ526IHcOA9hLX0sC9YZWeXmXSA4YMsOsPzcEoGtNTVEwcq0YgmvuyWDNXwAda2FCrj9ACFY
KeaT1a9CGLG7TKGnUh5CcRsCwZmjyhedW6vbM1OIexOMpT5iO5a0t+H+N5ofG3n6ClyCmsxjzzPl
6sJfH94s/FnLjBzDX4G91+Lrbks1ct45lWb/8ptTrX25gE6BkwR8OtDKjK3LHJ7BucakcxuF1tj9
CqsP+KnS0zxhcD13v/4QsC7lMmNzZgLvPEtHwrJV9sKyPSb8rNt4Yu4H28K2czAWcZ7kYfxljXO4
88WeIEReuLrlPdxLz95eGHFtEaMJ3T09tjBubOiHSf5kfOIEVZxPSv5T//4Q8zLrXWE1a74d5oFC
QVRcR9cxMOEMXi7aybIA3pyIphspbOMcXA5ENSqWOOzFGwBzXTyzvvCt5BLX4GmpM38LMVPnKxfe
ErFo5NS1Q+kn6xzhzoCrx1d+AvaR9g9tWp2GaXiiy2yY+gZZg7B0UK/8gqO63u3AGFPuhmI1U4zt
FxBZ/5s74uTrmPJlOyYa3VKAtxBWtK4NHFY530AetFzOUG3ldz0V0FtcHplBx6SSIE6np4jFXrks
D5FI516u8iwrHrR5VSybxZGUou0vZw2V68AjLCsixFvHGj8FXKjAMcr2wBC4mnbyxU7Q8dpwlpj/
FVIISYyC5Pv3ucj7n+IRk4AD7h/CknX8TBILPK5omq7KjmMnmHrcFzFrnVGS3HGG5qjTcGcoU8F3
gmziO3p3eeGQceVEeOdDS5rSJDmowkDJmrt2VqYmlr6f0XYbGrzjFmxnewK2JEnM+/arc+KUiE7X
EPx0p/Gdn2xMP8aKeyfQou8xJTTh/eMDs4CZoorQV0VIeplEcTYe1bF/gmR3b2G9JgAk8lTXB6kY
MrdTKNlf8K/jKA5puG+2opxRHsRU3iIw+lA7Fp8F8H2LGaVzPNv0rEaCNQ1elNbHxlOszE41SbIQ
BOd212RfsWn/qRHtq0uLRuW0/xb4BKAD/x4AzHzfQPHx9IBzc6Eqtsw9l7bLfvGEz7abTYNlnoDv
E/uBtAD3sXuo+LlzPOG96JCTmpNmKl8EJzdF3ooHtIxc2MEzHMm0xRsqdiu2b6Bj3A1B8GZtLk2n
dQq5EP6tVm03T6XuQ0F+pTF5vJ2hbIcOVvOrAeSnwJOZzhdH6U1r82866KbFDAzxyD5na3AKTICy
SzU2BYBGYkQjEgpdijJs/MM7ZscwOlPIHNpPSdQ3qcpwbyb4+iIfOkdix2TtmyQi3qgvphgEdazT
M2Ma5Sk7QjERW7R0kmN0SjPkiyxfqwB9fyC88MXE4ETlx5pltuDDzKhc2eSJDdVScCoa1Xr/SswY
7nKVQMWj12QJpng2II4nlB6OXHVbkhRFYQQBs03/usT27pIUUMnTPUSJTeTFEUgMQby/xUWuV/sx
GE4326w2ljzpKww1l8JXRIsD2w28JshHSpipGMhpiXCCyHla3MEyxjHkIXndVZjfNg1Wxg65/Z0r
iQvLrIrmEI+FBPttDOgj3qP5iQf6lDMCZ31Kxsz0eM7A1g96d753NbTF4aoKgZujk1Ee2LPdsTfd
SGBszBfuSPzeXnMbX8fYL/jWs+UBB19pBjCLW+wafuZRXWU6Fe2+bOLPhHb4eDTTcbvFtw9yXdAt
mssMKo90+p24y4dfAytVXd8XIV7fKvbHaMOLiECyp+zb046js7kkmylETjn1CWjxns1E55cm4l71
bHFiX/2qkj+6qYHtQhVGf2e84bM47fPN1kXfs4ypCLk+ppsGyCkIiR1m+FY0W2EK/VIgG2bFloss
fYjo8TLDANP+wwSzlEoe1e7ZaSKM4C2P81ZqvcDWVWeu1TaqqkItsF6aL7nPqQXFMLaFEzJ+IcM1
NOMgdD0MvPFxCtQ6gB9HRfmYddKwG5TTmDj35TODH/+Ad9PS9T+L1f9DhnsX8tOV19b98WVoOsSQ
WlrDLRabcglE2Crl0R40/3paIfl1OnTuvKq+Mc3RuFcQH7kxyDjZLZ9aSdLrZ9AlgJLT2rVQYNqT
eTBJs7sJcibhm9H6uTUux3gzK1+WsonwLQaEseF3AyGsoCl/G3M6ZI+5WGwJeDhm9TCutuqWJbdy
g4C2jGxa8i5unI9kLJu+rQLTZVH5RR55SpwxiUAeFLN7pTHYHKiaYNV7FcT5vMzRJRKgGlJYWAA3
oU9RQlqePQ9yoxs/iXzqJ4FMNkqLh0PSdZgq+eai4w/oxhkte4LeRHgHoofscKGh4KeA19X7cjlD
3tESAt+TGAu/XmxjwEOAyBFvWS/+m++znmeXnFGjpJOz371J/QdkADn0d94Wvyt2Kih37P5YTA/j
KerK4jaMtDAbv8RdemXjDUvXtjCpxCs+ayPvc/XMYw9gHMhciWVv8RT1WtGK4kP8kUbPMP1NhLVr
sngXgH2ALKGW+vrxVD71az2CPRK97Pi6dvyFthkHYiHEnN02k8kKRlfXiY/MvON9cNd16vf/9EbJ
DEFTFJ+P3SaznwdUWkcP3IQ/RmRQzvc56IonJUdemIATH622Yh111xBOYW/kLFqIi+wcGinF1ueM
J2DfEFbHcBY7nAfEvNoLxbTJ2n5qUBj7bvcbdSWweu7wTZcCvK3q0Q+yXW8Xz3H1wJXBcJdgfPiq
DXLisKSk0VSqAq55X40GQIF9bHBd9VccTvID/S5tFgR6uzgJwdnh60L4/9NAZnDo8k1Hv81O63lD
n+Hhdk3XMjAW1aynjaGAu27d8xENwzuOFOxFmTkrFKCWG4c82U3nf5+ysE4Ro/y0X3jxhPYAAyB2
Ymp/ZmPhZs6ncHEB3o3TPFArIXv2uoeZo5r4Pc/KggEGoZLpKChOvC+V49csfDSYplOfSGeY68jX
ixjlxKPZNHHG2lI0Q9S70M/xMLUxeBVyZpnMehubPXxbJfCYbR6infZlFoYmjuxPtjO5CnfAuDn1
3d4m4XlOvifo2LemA0t1Njs9EgnCIQIPevsmeXLpT00Axk72gasNc6WbaMLc5B8dG0Zl+BwL8gX8
dXi1aMUND61fuG9S5yytzYPAKp8jujSvYO51aWaHjQT3JMoMBI+67GQ6BkJ/7/Vzqvvek1xwbrpI
k2Cvt9fucQ0GJ+PCxv3HhkESmnPWA0+7nDMeEj8+bgWbTKoYDvSocune/RF3Np6JVrVswDXsPJ1T
sbmQfc/sPeb/eTVbtNdgLjJQEceHCIJ/aDkBbnC/5c3uYgpUQvrLT9avrV/XhV5Cv+0qdIYjA9Ew
nirVUbTk5EC04lACcqOcZlemtl0lBLEZouBrFZ8Crd2ClLtZlsCtGMkTLek4/hwaz3UdvCUBN/m4
f5CWkceHPkYtZIxBOX+yIedy4onGyyx4kgQxUnYakLZYaXwCHQR7XpdbYwrCpy8AnxCkX8GpOLhe
7K89jJrFOJbKx6f6GWGy2+LltAPrPRRaMR3gLRWxKJnuB44TFUeOuc0k4X6ZCFNdKTTKH8yxJ+oU
Zs1oaSEPoUL/mbeefmaLpLQqnQPGr4SywU2C37asGpZbkcFeqEXcnK2vZ8mhgVCsrFlSzw++14n3
tOIgvgzp4JyTaGHUOj42hDMivDqnKfBZ1/kOtxt41sTp7xmrPqh3vrms+HUjKV/G03G/Qn3YbfKe
epOnuJVkgxszmGSIQ0/zIXx1EYToY9/3s1LZBA61DRM0RnRWtHWrRfAxujJPulCD/MEMTFd6Vizz
3tIRw5sXoM7laMi6cUUUr/9Z6qPKZEa0yAI2NpWG7WxKjFcddkl5vIiMBxPmzqz4E4Nqp55rlTpg
j7lUrq9EnwR7RP8cliiPzRdxjhqAUGDARABTotIk0Pqs3wCGFs+bB6xcYbM25Gtx79LbrwWTDNU8
qPGkFM9Llgf6xV3oH7oj4S8XqSVQoe1g/Dd9xCyDfqIfM8KdG/wjp5NN/ohpVmbw5fmrLVzp1vi7
AMniSy/KPTNbnlf1quXzMO1nO+xSOlklt0VYRC2dOpMtXuBUWFs6FDw5tk/oy0sS/AiW9KGAj7C0
ACg20tsYIvQy2kCAEj6mbtJY+BSPHTl8ZCEgtbCvOSLnghuDPZQCin3nETicJlQE6QoOWCS1JVFM
1MaQX0+5PAQ9Y90923YeqRzGjfhsGLTrHBsei7VcZuAWlZn0l2fo1DtYtM9QatJqKzP2F0P6l4J6
GQu0bLCSvQy+EyJdd3c30XyZ3Vh+J+8I+1getdG+k0rZO6rG8QK4wDanUu5N2oeJ1ulenjDZOCp/
tSojBUS09H617KpM7RpwjJRmEauuB7attBe9oTFfddXbUEKuBwvkKTZZDWCLIGhS0aFs0KCDws1x
UYoQuX1mKxC3Da+p7xdk8h6Fg2nlLunBogjTTA+Qwr7rovS2Rpfoed4xZAHMwR+lI1elFwbVk5ps
bdKM1/wZzgfa01McFPit2ykQZlgRxrMhiBceKCUUwPlEKepb18SK7W4v4t5YEpch8XnfUZwYmdiQ
vblsEPBCMIwHNv8X8zi2VIHMRQguCE6sw29NVcI8oVTF3aneEm3j6xLTZ3lcP6i4H7MjDq9VO//w
cXy0rhdDMedimsjgygBPqw/VtKjCibG7VN6Vkr3sDRuxoVbLIFtuYb6n6bXTxToy59tnJdzSMHD5
llSe1wJHG/J4AoOCpnP+xf7uTiYa+sjdwMBZg5GGIfrPrICBdJW5rPBbtYcW/MhppqADTCOhbI0O
2aO6PuQL6xDgIRtFj++nGmy/Pw6mzp/NIlQScyVWHfEOM05R6GGYFZUcjFrObsme/uesREiYblO4
GbTeswURan3QWo8APezqALA90MClBz/yQjGbz7VXLA/mN3DWWFmBlaJT7DiBkXvGzCaPzOKUC6dN
8PmzMpHB2MuyzLzInnUYCAXYHDUOULiFHG5K+VPBbW1Hg39Gbz8wQuvAOgPewlboLbrkbxv8Ydty
BrmX9prSwTRjIffKa/HMYMX/bzsi/3U9WMcKVj506Sabp1UAO1i0PWZBpnRwtgt0XTiRrEokNpjR
mLp6pqqz8V2W0Mu6+G3OhOHOCz4GQXOgJI51qd3MC3oUVo5Ssjo6Js87IPU44NyYBRVHla1W+KAN
zY6qLF+rEYQD80HzwS0Lt5cwms7hH3WlZUqzs0zOKrz/DAQwYZjTBOdYZq1Aj1BdWpPSqu0jnulL
fuGgh+ddz/pmivPU+pvftjwYElV7jc3w5nFsKqCezUWKK13d/8B7mHVPjF/AHicJRpof6vORkMtZ
JHeiAMhYt9RPRjn8g+pno+gTLzey7UzPTMgE9n+bZxgzqM0c0M8Wa4H5+u1F1Os5Xi2LtZ5VpUK1
dPheKnBAJLHsNk9ZCze8N+tL+z/gf0uEThgkcmEPNQxZKBn2FEcmvczCtincVwgYuXdYX6qwS+LH
KfLsE2rW1Bzs2qnSGqkJD9IhGGLBVZ0woSwuitkJghxjRAJFXrLs5YP5n3P4BJhBaG+HQpRax+gC
JqagcSMeLQDAQLaNmZnw9hWHVe9DpeKEUAKU9RT//UO+WhSb7ZxLp25gVq5GVfLbr1UKYWU5Wsbv
xX2HlA6EYKPkx5AMuLE/QMy9rnyB+a72E2UFKfmczkxbtncye7IcMjr44zdPoIGvRsINb7YIPWVu
poiHte8CBAAJVH4vvA7KH6vK5kNQPtG9Ho+5kHeKGgzqPA3ILj9UbJDdSPpXZ4WKr4UVvKDU5+S2
THqD90ad8ZLqrmCOyEMZU2Rj/X+Zfutk+cGXXuM9MwCp4gtj0kzyPPuMosDsgrolPSs/xvNlGYae
CyVPuH8AfhXODsQ9DO+aghtC9IHQadQLMkg1NgUGhWXo0hHBUBL5tnVpGbcfTNvOCmwQDp5sEonZ
NAsVGeQMrMHMTi8sE0SPoq8jzM3eMomlTeHXi7kw08xPSBmgLoKyHwmhqi32MQiGuxdLvbZ7jdwk
ZxtaX/jSxxnCH75tv9a00HQa45EJK+Kb2ax9wZZb4poc6Ylr31B/h8EpA60WwTnocsbjDpRBVwLK
lENZFlyraHRT7V1I/4KUEVblIVZp0wNgA8vmEUXHyzR80h21LQxQhkC+gRVHwzjog7KdblCWhwlE
wJuYrXQ8uI37e0Als8YKAOXD1WI6ooxDfsKFVOEmUMqGaqgelFwSolF1sOCzYQsHY9zHDchaXEnw
ao/XVZgloPdeNAopXtn1iHIWDjH6xDv0REVvH+oc/pE9reaagsT30EQReY3Nk6ao+fQqhu7w7fQE
jdz0chob2es2c9uEK+4gLM7TXoXEG6xQvvFOldEowOa3u/tCb/6QBfRvb+L17LbKEaOyC90ke2Ob
FyaMtBYe0rpkVKOB554dC/92EiCmLh42QVPYgZJNldwjlwz5WAAqlbv87Ohz2VUAkjO3Pb7RP1CB
kOpM27cvWIQnZRa5zNuub+s3He1mqoUEovEu5KHQxpYPMt/LmsX1YGQOgMI5GCBe186vomuDVAJr
n6tOOj2mOt4Fvz+zcytZDNnbM0pZOeTQhcq7cDJXzEMWoowECyRntjejpHj7Y6nlKbNymrhvkrIt
udcTXufjo8/wY4vkehO7E3XLARkwJHUL0ojiIE6E1tvYBrhf5OWuQiBhapbpEWNnyFcva28eu7YE
wYYJr0jhJtVZrowXUIunyetT+y76GX11B88va4qs+u6exzXFJ27CLqlrWygl9siuP2Xa7vuuPStI
2aXNXuSBpYq2X4G9WMLYCAVDGxsFiaX7DqHRzwMhBHhSMq9ZtxwGXyXNjlqsoKM1kPhJZRR2FNXV
jDDRMB4sTHvVPXgYMgXIc1FDIfCFyvG7ZxLrQwIDK0PoGQLaO5ZuROziCVXsutvDkZbrDX/nxCI0
lBDjNyy390/6wagw6IlTttDbw1DPvPH1Gb962fxAFLI3Er5AVTfU9bBCnMumA+iabhkzrbUzWp/N
mDOpnBiEEh3BeqXF4VeQrR61/DyDbu1k3QtSSoE3x8Ixr51A3p6lS0WzusvXiqO1P3dtNed/FHIM
W4cYm+vw+PfROpxgQxPurPrMYwDyYk33NVwnM4k33q5bK+z3fn4l0zZJfLLsVZMxHVCJo1XLcJvR
2uGDRyffKhotQObUHLL0AA+bzPOFk0Hg5Cg9PWFdhkdCAZaI/qYhqpqJnlkJVsv58g4i7V4y3kUx
KpEZbT6/qPPeodmstBNn4zIhiYWtlFi6DfbCBNUu9R7jEgVhbKeAWh5oyLfb7VktoZ8Smf95FCmZ
kzrAgK8l1dd0r16Px2MKBNfvmnUFgPEY978gcpGPqyb+GQEhjBmfL+o65T2h6lxYO3UxCwG1CNSw
az5sC/9TBmPzWUzl69umyjeUeg0KpO/NxkgZjJYToVXEIAkeaRJODPnCNl8qu5ywq9RcAx0GzLZk
281aYxmZN2xg3RKJKm6kWc8Qxbk302usArYXrUI7Kl73DdoiYnu9ymkbP3Lyx3xfyf8M0F395dqF
3nFkRjsHhF4G/yNCwFwlHBBzrS5lzTjwBeDlb5VVfjHev8kznzF73wpGRWdWpiZ15dJRg4PzqQKn
1DO/ESyCw2pqU0h9v053uEbbPN2vaNJDZVK+xgN2yAE22OpV/rcnDj5jqsl7yAHKSw7BBeWD7m6j
rredpfYEB6J7dC8bbb1ubcwEgcpgdkxQlhxgTRBKJUe3hnsZ0zL2UqDBS6S9svABdjGmixDgZsT8
KyYriP1IRetORLpslCDht4g/fiP6xIx14o4JFuXXVHNwCiQa2dHf0k8OflakhhjXpqp0crqEtDok
jsVrAXrO5Djlu0pN54I2vSeJiVC5AeYtlt0ZHJDvGrUjsxc18sV+FdlnBqlgLp7bKWGfddhTBm4t
za0MHD8JbH4Xpdfz1Ooo1cXkN3949AVHhcN056xXjtK7Wxz0kjftGkhD5UBw1MRDx3Mb7K9GczVX
8S/CnOarQ62PtOhXPexmbKV8lJE7xEhoCS6LhfTtCxdW/5+FNF/W/5ZQQ69TNJ0Pj2/1jN4tr/xE
qQuMonbCA8E1BwNhcdc7IXbHC6mqQ1TcLsvylZa0mK/ZI/lUIDeaEmBnL4Y3Tr7fhhLQ32+5u3au
+gVU1yUqh4dggiIe1vNk0Pyn7UPgGpkSyquE6fr1AZBbFSjFJyEg11NP7zLeZJBRIw+Ym6Lh42Ts
EMdUyyb6luxJOzLfjtMPf4T0vz23tStKM+2WgK9Esrv/hjufvIhXGstqV656zLYe4i68tBX94buk
SUCi7ePqyfYi6UMDsEPrijWmUYoNlzsuv5rIPci3VtH+Rf1MmX2DIyR/nEchmMpz4RbsGXao5tUp
bB9jehegvHCGh3k63fu7Q2FAC28MayQU4hu6Rh19qiDqxkoS+SBIkGicqbhZeNYOL6xA6jzwsKwK
bg4M+kEusxeFAl40Rv6DYiJVcPj5X+45sgVM0HyHkWj0r+klso7XJDA2J32appZH92LvtHYFzhPE
xEcSBnm1UBgQg9fQkk0czVRngZ3tD6XGvp83si5giw29o71oDA9mcz0qwSq1wvuO/+BhFFbE1++D
dZcwMarIt0YRUwsEYy63Y6eByHn0S0Ua+eGjASocV/R5TVOPe/CWMb3axA/uSGM66/dx2EeqH/r1
EJzcDBtT4e3ZNOFmz62plsMK/MPjggdhUGyV/EIH7EK7NHTQ7sF49xalzKAp0v2RTw6N75Ru5zL0
rJ2pFQXEZ0b51znAXK24rcQ0yZFLnTBaZobAXaKgqheEbWBWgU2z2XKAoxjy27Sz9WdJ3LtaqNeY
FiDfC18AbQIMEz4anhs7z6LUHJ//Q1/K+e0ndp0gE0hqwHAurl+HAJBz8FHBSRRW4FLoD6uphoOX
f7L9pvPWaFE5utuur+P4uHYEl+/I60r+fMT+vPEe6ikPe/4wWQxdOIUwGC4pbgEhbEmELpH7KvBD
73CXto4Gat9ZpMpCe3P65TlLqrDCPy+ZNdkCUynFzCG5cjm0N4vLvtma05+OvYQP+mM5lWkZxl0F
K5MMZ0hARVNCVsmqbT/CmD4jgl108Sz/V7vGhq76H4wXkcQ+iz16kuLrw4OErKycOZfUP4QnuIT9
sNHqYrUzR764mHxmUuBJB7zlL1OMmFphkCZVKfXQKX2r175IaI4YLEgA024zfhYEneHqNeIJuN5Q
16bOXHPog58a+XXqHoNgK90vo8mdJqXqCUqblgdusP4Nd9sEHi3D4yg7DcGFtlpndAYIsTRqdHJd
MMpSIkTSuaQqmhlzn1r3m+dkd2VMXed3NFT4lj0x5tyxjLA6OSsOANPY/x6580354Dr6GHGbnT5O
i6DPzKYV0L4jNzwHYlcZZS44/jwm5FUe+FrjnqYudjLkWSU+jTH7D9njtmA0uVdvO/YTRlbP2fka
Ro0D4xKHsTA6mNi1Ly0XhJl6WXrBzw9muxu/DuCpEBVjFqCVP32sw6TI6jAbeC8Bu3pk0yiMo4tz
0J0SlJh6scMEyaIsEsGxergIo7NAo/aovitm3PPLrQ3jAGVMwEBQ0qE7FUdwWcI+NtYBIq2h3lWi
+gFlABf1lNpMjexe62ZR6xdUbM06VE4NF8ThHDL6axyRvmh4cXkhhoaz+iagS9O22zN48m1/ZtZ6
/EyJPojHFoAAJJRalFY9HxR9WUiHqWGiv/kHxJkp0TJvmchLi81ss0znNccqepxOASV9ouh+wgdS
/EcR915h5i5N4dp4NQLs29AB2hHhSHLBR0/DPCdQALlGLdMxEqQXQiO8njETLp0DawNVDoTH0waT
hHv3/SjSbCEbyeBbY1eOoy+euo9u83+TkQrqT+8Ao0ftgk5B99T2ptr8/x76tWu4AH9k8puGOyU3
bT76J/+2SRK17IHFQeGO3fiP2ehfhSq6HqI3/ZldH2E7zuQXQPNjo8soFHZ0nM/XAimdAGEoPfqw
xq7FClgOxcsWRFiYmNOvtE3U7WKYPnT0Zrab5tkpGjImhya8E/kUimwfmQY9fy3yUl+erWdJSDCa
OU5SUaOuYwtHZElDdM2EEID6lL/MFVPtfcCQApMfc8dZjvj8wNgZVs1YJhlbiCz3qPCbzgXdeA0B
VIAKNreir1337F1B54xHiQs7x7/bosoI+Fy9FW0ZozJgOUPTZLUafbijlHbor7cH4o/4z2cChyt1
brRy0pkFR/SXMEPDslXgYN+pE7gYISPK3HAAB1n3GWbRaa4R/8SKCyc5Y3qJD7l4aPBrwAySZfpU
NJEvxAjoc6S5e9YmL/RsFukze3U0rj0YUBGJnVu3cdsEoUk9w6DjUcHK84qd3Wox9K47D6igL9bQ
349CtP/24cLhMeXCECTq+1M5lH9LnXrRP8eCdf6FWG6BKtJVn5uz4cGLL9kZ/QLssI77xT0UVqk2
TRyz9leJsCaOHF7ka6J4PzXel/Zoo+DDGTGtvfgUtpkzV3r8zauwvaKGqUcsNtcAo7yyF3aBB8HT
IWldkp9ygvn0FVJip5nw72o7ym9+Tpem6OUGLfhjRquIaDN+NGgAhGMqcESL/DS/zU2m5g072YXm
gCCO9TRWJ8duvyf9Tp1sIR1FeEvTvLeGH70SRe8KJ7UJ7diJzpIQXZa4MXJ4ydbEg7KfNUs0Ocv7
BmTKrSaPpdEjfelauLE6oJoQxwGbe0pa5C4oSsKjgP7F7A8RillJNOy4Ay166nN7BDXUXwRy+Q/B
ZWv+56/oh0ltgIiXpgVX7AMtIjqzGrmoZ9K/3oF/oaCcq8ESM4xFjGnBz6A2rs8Q2PnEv4A+jk+l
gp3zro1JzsaRe6woDcd12UKrrjdyyhlogZ7+eZkwpUrr3T2nhk39PrOdbZ+LIwDRM3b5H/QDtojc
fzq57dT+oDAMsmyfv6CEp7wE/ho+5bx+JN5x6iFmL15K7NYpJC4RVT0Bs9pSDSH75Qnx7RM1AvCk
ABL2YTiLg2g7ITk7PKhMdIcLAkpwexveYnGU2xIYufz2vl0+i/onG3Hqg6cb2egcAvNS0mlCUScR
9bihjLGM2KHWKzRA2sgHbfHYijWkuvz8T/vDStmgjn/cSLjvy0wRmbyAnTB5PHDaWGX/9KQIBK8Y
nSh26QoyxzTet8g/q15pg1j2pj2GcAp1CyVNkzX9JEFfyxPFsWyp41POOUGLHgYmvF1IuW4LxIZM
F/gCZ4aTZaWOG/nmts7cuw5LkWYisMScdDT0zZoPhf9jeC/PUBTzG4Q2IIzHFcDL86z8f6QqG9zx
wWUYbhuO9zUYTehPv0IF/GLrV+RbHJ+TSc7w4SCgRW2K8wi7ISrQvwIcOIxQCSVb3Fk+85+8DjWg
pC+kWrODLSTi1zlI0mHVuMFA8y3DCI6AMxpMitcGjulSLV3m/JoGe8LknoLiSKA0B+ce3F6Kc0Ht
KCUj7RfvVKphIm/OpPmt3pRyb1RBhiL+IO/RGlaUNMSF8sZ2PclVMBQeOoxWjSTGJOat9ShjKa6t
V7jFLw60D48irkzPpSIXvEVcx58WUnZ9xq5FJ3Pbtj1YIoOM1RDS+N13myIzrBfqHsth0/iOks/b
Bq7/sPcYKaBFIaP82NKIJl2YY0BozDsAr8ot0b+P+uGwC5KmqJWngZ6rTff7mBzRhaBeiT0HBMli
sCcV7spYajgiaa12AgyOX6Q7REWcAmDULMvfSLMC4i4A4IsiRHuvOVgNkQNbVPpO0FPeNlPEkP0K
wnqp5SZcMiAQ0z9SN+qkM7+H/FKKUFMk9eAIDzdYdzabDkU6PJbAKnQFPrzyXsjQU+LI2IR0wZH5
NYL68tTfr/tYcaoKgPq5ID3he9bSyNhSb7zXiSqdoIYIrtNFW0bvCexwMCPGhP+ZTCeF/aBD0rba
Aq63YrnS7KqTWfiumJfTUTnmSqE7oshlzrVL4QgrrHRt7F6PuQnsGSC7fr8sgze/x52LGi1bgNv1
8Lj5G6sE0+tCIEmI55L5/TzeLNBQZm0dfHqq6wiQWxFKyA6KnaY/F8xep3zDq/S1wGOWFKDvRBE+
JFTMSanZKWjbkKIs3h277mr/5SkVHdEDMKRpA+ut6rECoAtRDAoUQFrQ1WTIfLDi6il/XcML4EvG
5G0nj6D1CrT4OTGIV/ay7ZtQBcwxA6PnDcQNhgZuMmJQl0rqBqAMxPoMu8sDb1Uczqpx4h4QR38T
LTs02bLnBirbMrQpAQxtyUbjYH+TxTNB31UjSZ/BaIN2pMkyliYOR06sUct0WGJeVb4sdfbpRNiC
u42hb28FvPmhRCvDrjybTVtTCFsS7df29YmqO5YrFx93QoWKf6npEA4utkJzVy2ZmCr+gxlvFFwC
7bTeguYg2Q2pAjqMcBwCAQybdYFd8T9+2n/e42n8+dm7cvHUJ0yzYyAA4n01hGyTYt6S4sjL6BOz
//iBll3iS/F1o5JOjAji8AOJMvkeB48/b5MHHynlYVCGYlubaI0rJmu+CBAgMt79Ldj/4aF5K4is
YJqfY5NMDMbi7jEKVR5q17oBsr83d79syyaA7GycPW6zuzaEyobgMtOq4nMWCF28xLW+/lle20Ir
H7wk87kBtY/OSiRXxsjfp1U9rwOONSsRTwI6CMydYeWVnOp0E8TaQzS1/cgPK+NzGt1z04zNMK3i
5NR019QG8Y9Vob4k/8zJcxZl8M5fxkP/O4q0mlU+aFBYh52/z1qV5Oyw6lowHjStQXPkFQPvLtHx
xtdVjHQDCYO4hVWuPfBNla2gP8KZ5ktc27UVL8f+c8N/TNSnm4Hcku3XMi4CQa4uqMHjiCNjWG2y
qv1LGfFxAhXGDmh1QSLSAQZiyyhW1/yyQcJHmyJLKAwDvGxj9WWkNL6bZ31T5j+57RxvU5dMYe/1
c/x9ksbXNuxWBOKSPxCYrvRU45YniaSUew4/wPU7bp4Ohbr2Z22JuYpJhHRNbUkvdTyDmrJ/esZP
jhgvArk/TpepwBAA/MMoEZUrReGberTT8jA6YDaTs+6zZyoeO+VGHdQMGJZkKLQoz6pVM4HVzvFK
RDRLrRfZkiwu4LvGFAqNBaQQc3X6fd6UJ3gXV+rRSaGeoUmGD6sgY4cZNrUqDaSw3iumzX+il+OO
8qSUcusIIDU6d06OdVyosXvnE8R3mlBmb7HKlnm5hRdTL4tgxaARtWf0aOqcJGten3XRr0yvX+Ka
XrlcjvGEfMX8fQKEL9zg58EqVKYmUBjZq37dd/J6biPmc/7+R/E/+9qRjTEopm37BmvljTQkiFdA
5R0m8s7bKK9IWX5NlvCeO6lflEEYF8X+a7Rgwtq1hZXUW23Zplmokenn7UK4tkW1RADn2H7fSyQb
ERDgxQPE8yQ5V4hGAoHGAlTzBmgAcmDyIn2c+MGq2U8/qReAEDToc9rOxElVOKvqyUmAnD/IwMxD
IlKqaR7ZHIrX+/kUE4Px/V1xCCBpIG5+wy7g4/OoJy8mrdlyo32J6r5Mk20sLesUpxfiBsRpe8d+
kouWffV+jgAvLm5Mmyku9u62pRF9rYjZaRxZ2i74koBBaAkVl+lWed+Vt+h1xW5yhvSDvVmVHhj4
zm/tmAAUFh2Xhgx3arhlGpo6TRBJYNPxzHFcAymNP3Vo6QKFMD1+nuen5ctm+/c7+zLQYpiR2+F/
k3nIybYePtaw71RTGczBXy4i1UTXpgYZfXvHu18RSKa/Fdh52Yqrh2Qp7JfBYg7D97NbRjK1lk5j
1mWxu0o7+IMgb2BJuyt3TGDleFSRGEIqluy6AEAfO9VKFvJmlOQW3WNSMfWz8Fr5kSExP773PLyl
v9S1i1rwuKBPBobZ9FuR4xYPo/b26yGUetTjy/XPm5R5zqHeIr/Pd8UYrcZlM3BK9w3TQ97q8KmU
MZ1HZSdnxl6wyZOLukvX87pNXlDPPAPaL997+ozFTTI+TznMdOUUN/Latbk5OgvYxEGZsAAEVzvK
zplkIUVaLqzkHLtFiXKaMg9b77M4K8oW62nyRjuUevK+/k+LuaAmCBo90nDEQ2goW6XL34Lu3MXs
Ba/2ujANTuvrjG2pzFsBXZptEmRpboXhnusNyjjTE5DaWhlyEZKiaMVLwuHcSfN6qyrSUzO5pLfy
IWLLVSaeUFf0V9hGEgpKAR0j/lVIeMiEb5ZUFWrsMpCVa4dAvZrnWOM2eRaXraYMdk5vLmNzjH22
sWm8FU3AeaPya85nXC9QbcNaJDlkMh2ZT0EUVaiNg6idPuP1sh1x0oNDp4TEfrq9o92jaFpFuto8
cf5D8zmHd9i4qlKU2LuVoPrkZCpiDpVYtYoWitqFwMPN1UVD5lRMrEdhZVBQoaql12fOwFlILZYo
Pc/sa4tkG0liUXtKXPuazuF3NkoUm7nXFFr8zw91cIY1b7KiInkI6DcKVJDXTzGsGjSDko2ZfNoh
kk8oTRadhaK43zvjZLHzp9v0GcuX6o1YD5Zg38t3oJWwhjFxwBFQwbslK8+cE19qK/yjUsmxAdRB
Ns5FQ1O85as0ybPsqwIYVvOYNDYQFB6uRVBaNU5XkkTEscYbafYbK1WiPLi4pULAEYA3euWRaDjJ
/Vr7bPt59o1caV3/y0ADtWLmhCITMr4ltVrPHPOP5GFYIH3LDO9hsSOPrWCCojGXO78KL4wSLyMC
FY+iATO+EDNjDLSI8vKdwc4Eonr/dSBr3zRGJy0tPAuydJqzPeGhnMEDpXWYoTy2NFhzfo5X53f7
RIz1AJMmEn7Bndy5L75SWe+Y4znOtAQg/Ve4Yt5T3NPXG6cXFgRc6ve1LTDBqNHvu7yXvrWyPbEE
J2WxyQ0Yk8uFIHe12yxWcUKMensg329sWnGlhl2jPVxIms/+5obwirdyeBXibo+4Tqa9zg3XgP/h
/XbwB9N4X4Y1zCI2+SNgWFOsPZfjy9d3/+v8a0+3sLTKnI1oYmPqFNEZiiKTrsG7eFOVAmBKOLX3
YJvlDrp4xAhn10pvFuvQJctNETjKCitKdjzPTasOchXTqp+5KJJNxRB4+/x/bouelJxdcv7KwQYE
OItyqXE0Xi7dRWCSqUaQVG/10CQ4WzoKAEtJdDA17tJeuAq7QxrBIOn7lPo/ajBuCF9zU1GOUMv8
L17EmlGn7AY4FCPx+idKiF4ucV1LfwX+19F7i/1BLJDa6lBur9S8RRYx1EdvLFPdhmuGzo5UWYEl
eT39umdiWzO/Kszrux5+d8GZfUXuClcCGz4K/838rEpMB6P8TbJQ4ykhw1qkc6n5GOc61HwG8QU8
Lfx59oBR5Nb+BLO6PQ89HYoSxnPAP9If4BI2SJcsphQz7H5HIYTq97qE9F8r+vGXGVYCw4BMZtDa
vEDuBr7J9g2L/9+RVeu7WqISPlHzn1IWQuH5yAr3YLzE63zOvJBuSuDJaV89eHhjBTsxprkj+I6X
3/6MU+FIMo5eMC9XiB/MJCrSeuWMBDmZLYc8Op9CqNjMqZnn6WFEsc2YshMfRHgoVU39H2+hfIyX
I6muyQdQyNvKufY2Hm6ABJ1B9WFYnNCD41H+iHPbqA7Ywu2ZA9vKBslSJiVfY40SHOW1EJpy8uO5
xeflsuXX2WjAofEgf6rJFEh6kN2CXN+eAHYCsfib3eZ2ob6IIqfTqsdZ5Ut5D75INx96qshBG7l4
zs7n9sbzB6pZvE0gL8h9QhQZc9kuVCtHWszJCgxLeThoVB9GgQzwLS188PCtX9SQ0nvLemdDbzvE
ofW6vdnLdjAUimsYhNNh8ziydsmNWKbBimTlT3L2B6Pi1y2wWVb05ipOcjYkYEkMBPsHfLV9kJKb
n6WrQpEkW3D9jlgPy75TkYzxCIK1q5OybEvaE9AfOyL/w3+Hy9h/3XmW8OTCPG/u3XP0CjPQPrUj
C0IFiANQDuG4qjR3DbYPrTYfygwfGpGuLV8NOTZk9iJKVzrOOfn5AtnUnXBK2yfgfIcEv4+zF1+3
GLL/gPHXvs3QtjM1Pke3ONevoUyqUJ7UhfeqglM+l+Edl1Cxg050zaNAftONhWCYOCjgRGWu63Pz
FB7iLnHvYV2y3xFF2KnKnmQUM8T3UqETEDkWjdZGIkWclWWZjVtCofp5JaoOJTwBojZauSD5R0Fr
bS3bzjW4RfH9On9UbXI+ql2KAKUAvJS4DEoBGPPvTnnHYty1AmjoQnhpLRqrR4FOxQkylNwlEXX9
VtwtqhcDYhcZTGT2v+wuXg7Pw97ylrsN9xOQnpf+1EyZkwpWsO2Q0TFIHTdZ4hAbNVv//iKCcBR+
QVtdU9gO3kAQLZItIdZL0CTriNn56+yRCWuHTUzYSukq6AMdTBOtjZeKgvO88+P3ijrv4KMJTyN9
WQYqagAzB36yRmCn3bLvsqhs69Xc3UzWgCzeDF+AtJJ5cPh+S3OpT+QVqYFACDXuIoRrZGf8gCi2
HoOiYUwhb/DhJe5JtQqLi5LWaNN/zPlPNJ2YGTAAe+J+qvSWfHw77OiyjIfylkzRaNT0NYZLSjJ7
Y25y9y/2lH5yFqjWfqkZiZcMhFI0pfO9CoQUDaWDUD+d4uD60UHGaodA6OBMnLrmoW7KIwE9YDgM
3ijh8hQ154yCY5HldRFwY9wUBgZylitT2EcKDs66mjzX4VYPkjKTTGNtAml2diWHIOs/8k8L+AsZ
rfkiLBPIOH18aVszktshwqKbQRmz9vJzq5vq/+DJ5fSZ1EHlQCAfJxH9XfiyxiaKAN4bJ4HepOCZ
rfdo7BwSlZo7FyxCB4um5h7GRVaYUnfin4yFGgO2+zLfC2S2PqNWSu5WbtOMcImNk/DfLsKJZixL
4QmBlXHy6zx3y54Cr9YBlh/nx4JRJi7Ukgi5hgxKRfQsuOwFuCRl78Gx8khYS0LHu3JIamZT5nAx
IlGAMqx66rnexxZW/TZAgh7W+3X6x7FWyX8V48JEfx3qhMM68lsueR0Lx6/ZKeZ+4xwuZpP4+Zgf
eWBy11lD9ykPC8c1UhNNX0L29oW/S+1/s1tV2cpayS0OyuLDzyVwMFCpVy4/Xoh07y383wqdK31u
/HATEUJu2zEUY6ylABD//Q3cSRWx22ct0jK9jFFpWa8FWv/S/8GnsCC5gTp4X1efevGffNyusYgq
rWl1AUFCB+SjNYV/IOIH+wFGuOUZk5XkWjUK6W10mILPMT3ty7oya0LMgLXtxr8JX1rib3dUHvPH
/vuodP2fmJvOlc6zmsluAfPht0dKKsGSxGM+e9RyxGfPJcG4oJ+KvfhXT9eSfBPgpU4MMCwuhOoD
s/A8YfDTz2gp35B4aOSA15HWORqzhglR3Yp6QmKSmorsuuMHNg9hJicNITvvjJ5qxLwoQ6a3jCZz
AA8WwTOOTiMsYxevtCK24bu3IdIprBZtIzsorJAN+Apl+RSol08sLnJ2SC2SFMl6TcUp4fHoETHg
aM6e0Ujjw7rrc8AUwVkC7FVecNfmIKrdKLxeXVkX+cmgUZwPt7UofBSo2JdCtoSZSRX4nqKMWkKt
R1Zk0eSQx+KhlX9MNySHllHhN5n58H566NcnD6ybikbsTiZseXpHNjmkzV1br/Lc0hIG0OB75r+2
6D3UgLTnvcgzIfSIKXeNU1+lVYl51IHs022XAIyFSjHHSP14W0E/tvwJzZwsAwisr4VbWkHTUamz
yWLUJE5yg0N9uV2OUEPIEfbGYygjhFZfZbjUvAwKt7pMQ960Xy1Xg92xYKzmsC9RSoQOkIDpDMbN
yr9FLzRb+clp4WkZqQDIXzfac2w860VTbFzdKjmhOzmttcZdeTmN6dbdS86D9UlK+T4QnRJOMOWB
PaqBMjYpx78a0LMxi84ij9MUKHPW81vhXvA+DlUFOvMgeYwM21JzYr+VIVNAFD0PmeSfnFvwd36E
MCcjUekuixgb1ggUmJb51ASw0A4YySkXfwQVMyZeW0syg7kKNs/53XZ5k3JxHFHWey3x/a1jCLss
CWs/eTJNCr8+cLpyPvG9Q6nKvXlXVxFrlo5jGGNt2W4F5E0lWjpAmj4xBaWtkL6GXGt3H3v1VIY1
9ohjn/BJoCnNQSs9C7jrlqraR/64JgKuDVW3Vd+iZA6bLKRsDXwtgAo6r/rxvfwuIVDbJmHXCkKx
hbv4rBgfnN/LAKhV3VjwXM6yDc+a15dp8WV9Mft3opDndUsCLBCInrNQu/5oEtXnuSrAGEl8PmEo
C6Z40ughyD73f3pGSEeorjgYpPqoxd/WZDIWUJK4nl1m2QePWIHD4lXL6Jhdba9OIVp+vrutvi91
UoFfxeit6IpQk16M1FlBuCkQ/TrpiTpDJZw4nZbNnkw/81JNTTpI6tbfpWdLEENLpaj+i9RzfQMH
HMl24mGM70PtSN1xKjrYFyASQ/p110ua3JofcVXnIf5era8l20OlZNbT4wJ3axu8+95S+1LMibPj
aeU37V2YQzyVwmjETI9hoh7xOwbFvFBLBqydHt7qMOaMywWSNhleLzpiiCo5KCQhcL4Z6/xsPZ9S
TnITklG5lgRjCDlAcbn1W1LyFRyoPdkrbiR0a8pSFOXL6DPBkxyKYizz/n3NP3x6zE3A0t4MzZP4
zPTNe3TZHHkJE62tVK/5Euo6tvlzwd4s+L0nkgYuB62W3LvAGqIMJOD9L3JxoxZsuhzy4pDPAngw
27/69VhX/CZh5ZIoAGMDE6QETrsh5McWicJenVxWbjR8OfQAlvwfpbxytGVrOJ6HBrGZ9J7N85MI
XjRwSchWllIvHragOoqbu6no/0xrHDEAmzAtLV1gBe3Iy4wL5RVvvsVtuW5oufBG/vDNknwCI4wz
3zr/xqFa/6xtggE+hE9M4kio6mPWtXr2ZJEA+T7JzJlpOfC5f42+pM9I9cLJH5yQ/3piqKRNF8pt
p0aFOJlpl28/Xw4WMG8BMnhMWRXHP0how/3yrBCM+nWo4333zY8tpMIe9PUYTzgFeqTZtrzBVKel
n5rj6ykGiGIYlQKX4/mdOQEAmD+by8IX2F0vbSiakSCWtn7aRv/Y5Dx13fcDuxlso6P6XH3Rr1sh
ogisyvWdv3Fpijxv2OcfgVUtUZZR8bOnronKVgN5ywwSx9SvY5SIobDEEyexRTlTN3YaJ647r00L
omVJJsB5+q5G3cu5oPQyx86lJYwlRd4KVcKIiNgIv8JXxIS77nlppmc4NiK/D0FRIOKvx5Eib6WY
ijzQU6eBM1HWgK63RLKvglmn5dqeiHksl9V+AgfX9T4olVJIkrk7wJG3DGyqSTpCtSPKv9EasPx0
ljqDWlpoZhxlZwXir4ZTG7+/lPcfxXstwWbMGmE2hHwQpHwFaWpJmFnr/EFwFlAQISxh438nkj60
/n2ss25veNxoz4MLuWns7BZ13YnCobTzXv4SyCMgEdW+gJ3s4a/4Pf+qeYQbI8oRTHHpWRahkauX
OZKjoc55VLrGxIGBd5agqFQyrtmYqV3Hlmu84ziQ0uhuv29dg8pDbFlsG7Mp3pBzR2xdPsQa19Dv
CYR1fg1QIndkrDcqEkhaZhbp/RKhXVDPKM7XoLIeUJ1fDJy3LYuvDaRYWg7GVmRJKjsk3J3IywRE
uL3I7dDQDTvzFBC78zjVvUgKIgpiFqDFE956BypObbTruWta3vduyw9ohgyg94MgSssq8jgbesju
gqGEoYTLCeYLvqZcgi46VOw7VAb6+ev7KoWR2We+yW5sBttT+QmVoWQHZAS4S+cvqMBTiZRJV/BP
MdUIQ4Z2RQRGUypXGt9w/7rtK/aO8XgxcP/0w5kYRTgcla3sV8W/FCHrBx3OpDWzGmW/uLTdc4fm
yyCrc8h2RMySlL0KLzdDavy2PAQr2+FMdLzG7fNcMrVSFNLL5XW4XHBsjNZOfKLcEQPY2fX8ha6c
n43YpoR3cL20gGH0PaWI9XpvSxpGsrD63ts4EVbL/scccOIEmB/ZUHwtYLO4hkZ9H3PGPrBN8UmS
nH0cl26v12r/GASmDp7drt0IqIJT8u2gcKQr5YboUA+ybqjnAWigxC5CenxjebqsN1pw25anps6Z
ItIutX4qi9ENbpAB/ydbwW0YaS6i+u1EnfCGeML/LvEDMYDFDDkXQSbOuaX8CixtiRvVgVo+ak24
47ERPTu9B9YTg+sLmD3hiXGnzN6AnRmr9c2okQtK6BUvFPq2T1lJG/VCWN2HdAiJvmPqjMVvFqbW
8xKnZkpTXXkg6W3WqAwMHuC8nSExyx7uIJn5q4y+hKkytNfkD2Pm3/r3qwBGepKRF6AD0lTNuNiy
kfmbevWuu5wsfvNZ81A3P/QfxYuliyY1QuBsQGUYB1IsC3uVTe6KLqen1l/7T3ggPBaozanw0kkX
kXjARqU9bW6qvX3uDFfbVo6CV6b8XNGEIpeLDALlYMox6YaEIIct93dv/R7esLpIVw2ZdjpmpNBh
RnqF9BOdqcCxfhaHiC9Z+X6B+VoNGfIBpD5j45EgaYm5k4Icboz2cHN5APM1IeUgXxqQeIwGea31
clOcyF+aStbYTRHRcWqUDJOKy80KQ5pQrcRBNrSYOdnWU49aEoDLitKn4+9daI6bQXrlmdvlX3Ms
YzPUN4AEdg6Abz9eYU363RoIzKBNvHNenwaKKwe/uUQ+Cm1PeoBAY3+eumIieLiG3cWyWrXPchA3
knewyODYIchQ6+ylibvGxo2ziMaL4rsV8mjU718pkwvvVoCmd0voAlY4bSBOTQTsxPz+smqNW7YY
Ql2eS1wB6awcgYz8X5P1vz7HqnDqkL2yT3d1Hd5effQRdrYj54bBgPx31skXdTvbo1k4ZkGxH2wX
0sIR1xEHpMpCmPPh9rBGb+Z5JzXL7tkX9FRBgvs3N4hFQVxe1HOk90Ez57ixs3dFjm/9+jP2kQAx
8gM/KGLjIFl5DuV29wulWCftKLygIUccTtpuv3iuFiz+kE4Jayl2Z1eHSHK15gseHO3Zzoau5GKI
HDeLJhjZYYgbFGt6Ffoj5iClt9nHVf1eqBDTa/DLm7qoC4afoy9VAVYvWQZVVRE+xsFzZFKdWh7T
NKgZrJfOJwxELUdb/E1TEWJDn3Ju/QVlgcF968ox3SCWJy0/v6oJtsOiWPtKKrlwCOHFXBvf5O3Y
+8i3qEb+2QFNI/Ah2Vqyix37przi9CwzLZmvB0j4Hpd1vy6ef/aZp72iMSk1OjF6SxztUwjkQkkU
qVO8chxdSSzFiXZ6HkxBcz1QsuJrDrT6LX7PlAB314iDDV3sCcmXKD5a4RmATinkCrG7qMpZf39z
WUaNV7VKVPdgVre24Fi4ACRZCua3rym7LGruAkTYEn5UTEK0o+ykOQJgp8O89J+AXUgG+Ip5vwjt
eRnL3gaD1HBBiRZ27y1ZJNu+hwQ5De71SvNKv0sILk6xIqzHvuBKuFX+UHa0JkmTxrl/5vyFox6z
Fh/C3mwVivL+/J5GSFX35WAlMdkSKwTctKQ94ye/P7RI9IZ5Fv2RUwvu0bFjEHi13T6j3Yltif+1
ATM+ikBUhDliSP/DpRlkVRuQVWhYPZEj+e9tI6g9F0MhTWGaowaKTQpvRf4xBo+pJRpD4pySVFVN
8BdbyJy/Clr/0tYwiqYB9jxQaOv3BuxuUP2FP3+16EoZNRi/fY7EwcM+kLFJUhUoF5a0w34fTTnm
i0A0yZxmZj8aL6TsgGRkJZslqo8D3RPK5ByQbVD5AeMjBWQBCxsKerOy/36tGD3UZJ9fg7mEIyqy
6hNkawH6KnMoXdnGVHYs9/2WewfT1IJVwBuwV5LvbkAAC2+167zO8zlntgFiyBibNP7zOdEpEgJp
b2X4jEAh+qtEoyllEUkIjEtsceoCCJMyT3SDjXgezVeoUBw/C4j6lcCSM8grvf3EHpwsfiIf30zu
fiETrTt5dlVrwZAQPjDuIUVwMG7j/rXn68LK9n5X8pjFnD/LOQqgqEpf9cdAe7Aoai+nM97sWlbi
+O1r+AexsogLGTnxlygolXUYXAgK2YatZCrkymQT6x8rU+vVCgGZb8Z0VP1VL9tm/HSORDr3BQux
U3E5j5g7MILYZL/IQtqx16eDYFpegwGpupvz1ZNvjpCyVuVo/Heh9FTvV01RWX3MaXCrh71QM4jl
zbZHEk5K/DzkcdAESylXCMprdCIdQUdNkkSzQS74MVo0iuFAJs5QFrUEGPjlYFwZrtEnCukIF7dC
ERwTtfGhyCkzTZtBZe7usCv523CP7kjDSuMRAzUOUSftTJ/IROI5ofnygFSB0NZkXvXrXPf1d+uw
5hyz6Cxng6V15v1ACPhyAPHy+LtB/KruBJm1yCHe5nUzXVse4N2qMgiYrE7D/r5HLGl5IdnW7B58
9Z6Mc7TKAznyJM6hP6JDNph1BxUD3axjVxj7xOI+kxNRBaxfTu9xA0tiovTqpKDQ7XTiG+skhFZR
9nicmjgfvcErbQnY3IWdRJ0NcU/1JSg2bzeyCBwHiJpZQrzT3bcya0SCRrrKs3lN9dnWnjBG6nnC
la5NUV1U2JxQKjx4O2Mvtl8+vxWHnlgxJl/UvVipjAI/NispMFwHC6EtS0BAK89QYQs+SA+mfzN+
Gjh9gOChuCVlBTXSyFSOAq2SxhB8+pKCgeus8cHhf+lGROdWTAsGi5w5pDd29K2wbNSaTryX79Fh
laOQmgy1LBU+YwzQphIlQOa9ZNh3J0b0NcVX25raB56goRKh6LF7d7KF/MBXGu7YYaLgZeDStDJM
vQrOfEYCIGpJt7XMjLOc2aA8sRimqNb+JbrscocuP5cQZI0eOqzH4yxKF/J0UUpolWoe4P92iiyt
m5t1d71EH0G533eJGHa6XPpXcoEmS0oRneMS0w56ZsaOSumOMv7l7HPs35ufltqMDhDn6Wh/BySC
/ee/knn9Mk37w7BYh/NkXgx3nYUN71oJv6ROY/kh7hb1VQxIkQ+igXzOBvVza9JIqDFYlLGXS7ki
P2X3J5PVlbV2Ax6/vxmVxU5bB7AC/vbdXjVKjhbBaeJDI8+Bvdf95xCPq5BM6qK7HmZY1j3Ivdkw
8GzOBQMnuTWYam8IewJebhU3g8h23PfKkYUCOuJmm+yDCxVgGaJuwQPdrG8G1Od1Na/CK4sIMAfJ
ZwITfMHEd4ToUIYHl8ZiwVIfFwD+MrBKIAsF6boGK2d27qeBOsuyoRtRtVvSZMaPZWyv7VgQC+wd
GAvaR8d8UVGRD6ET01Qo2CXynIhX+q9jFUk1TSLqBEZAmIDjnJ6K5s13BJoyi3KfYKwSgciGeoPz
S4OrJEgjBiu2Nu/3CcsddyMWTkDagn25q/xuNbmmskpyQM+Ogp2KqCk9Z6rQaEr9h44s6DSVuZy8
aHn8Snqe2cxG3pfFxmK+yeVxUXYwfVWYtcwBUgSYCgOmTwdkkrKFx5ELsUgI2qmGqnp8iw9xZZ/Y
xGOtYdcxpfKMoqieQPbGBEBuETjLCR63yzv7FiJAV9QYSl11jyQ3QrS6o+rVPtZbJigQTZJi5X7T
jACYui45VKClzfP0ogdk70KesVMgRgSL3C3SkgZ/8RRpLqeAoGHWaYj3t1GuB4EA7xREsJ3Oazha
umw1+YpxtwbVGn9WQxa756c4TFgc9O0yzynE0T0gXmULCcWaqgCpnfktBhTOA1Khvg1OthNgw6AV
gXAwecYdCKfGRxDqiMktL6UCKkgyCD+vez5B+cMxy3MP/7NDjFLz1rXryWNju5rdxww/2+je/Z80
J9wEX8Ed14vW7r+Ru6sr3Pdvo2MLUeLd/MqyZi08UNelVywYPQf8fNOEN2jiCBIkQzRRgT5CPrd6
UhuiXxoNg0mQtjDMPKAUoDFrS1ymGQTk0nYVijFZ8m6Qfgbo4M96Ueg2m47IbKVTbIzBsTvC7GQr
7OLT0krdNX57JLEV91t/ntQ5AaQ4vqQjPu2Q7iZSm+W4K/d8m4A7FRpuSqqyoQkF9PxMUEJq9NMT
Ps4GOUTYVgCui0p72MPZjDwX/8PvRilTit53wLjWoZgXa9X0C4+v4WPFWip9wc7VXICE8sZKUgAd
9Wx54OLF3+/OzspxtaI9s1aXTTqhCK8jhHO6dx0m+lWF0wDvd7tbliCkuAU2TbGvbSCLvvvZPvhx
1Wa52r0uFwqRsoqGouP5atY0eLuEOhPHrcMZdXwopmYOG2rMZZB+EoG8bOlAsLxEZYnWhZHKMWsR
bvHBI2mixeita/kgEQ2lCOgfsGgQYjbk3/vCqVHpn5l3bv7GF0JsOs7zx1tqex+bqY48ERI378lP
wLKTalzXv+GXXkibUVYbOgxjg8Yb5+uKo+kmJXBpgOFIVqnN71D8S1G8R2ZD0SPvSz2wOeeseWy1
nNqeNssmwezxkJxPdcXo4MrzMUBLnusFk6xsP/K4rEUwDdU2O0uPNEwpBG0cgOofuGmh+1X5d/6W
sVH/L47lFWhqFY891Tz8S6s0gRE/ItpHu/FZdFkHuB3mUHvYGEz2Pf9WT3fskB3H0mOhhEYMC+Gu
e/szg44aKCe7DEJO/rLi+xwl1mRsRWuKNsQf3ceg4a7iybs395QqLr0NO4lYkkdk0Ecn0RpL6xro
MMse1FWhtvqZXcEG/QftLmzTmM+RUL73QguV0htq9fjsmz07xdtEYxkJvKtrOQ7NlcGIf/AGoyqK
txORFJ5XQYSzIMwC7UYyrj/gak02xCGfNQIFWsWHxnuiw6Zz8HIRAqCWWpGEVnG/kcyh1M35fYPp
+2xR24poTd7pi0MGy7OzImz+76pg56HRK19io8sx3qKDRvPAztZR+36SWrSzEHIWQ+PIbzjqqmmm
m2TACMA6KQCIXvNI4KBeqEqFKBAIu9GOjZ2J8/+la6MpKRusF2Pyvzrb7Mb5RmZ34CAXxXkkMSNH
ImawPPkbzV6V0Z0IQK6BI+T39yTa27XEi6h5s19iYeUOk3SODuQEisIfY1vCamJqT2i89RzQz22C
fUFsN3IQQggIX5xoC7Xy8lHEpjaLo77zKo8NgZw5s49YiK13SHrqujTArmm1iMCOgwRQ9DSt2ant
l79fdlJO+IXSZ72Y8Shknd9+XgNFO+tjI1d0xfx+FE5nGS7frKohNOd+yVPnWguaYmCw9HiznS5M
v3D8Y9iT0BWoRXg6A8Z0lqSNzmU/uLNSyexdK7gF1r4NPpcYwuGx4fhdLWRp75dlZG4iw6i3ZovM
Sz+Z76x6FoapQEDhdYU2LK2hqFXt+brDC5bdT74bae9Q31ys3fcKBfeiyGteVLdE4hW/uID4dfvL
Bo9eZq+LfU5OEnFqedmMD67MT+0EIsK/C1QFFA9E72aRpuFjUB+8eQPuZ1aNXCRksGIRsbihRF8L
r7YVehlRYEclFQHzhffn5VwEnENMGQ3FmI7Nhe2lBX8ID62n/BLwFQNYuV6g6ZXv8PixsEIWBAhJ
o4o2lCXvS412arhTMICC5Mgu6YrOeaVN6gPS3IheI/MysW7WNadc+RquS1H8DD214KV9/NYgsdTo
retjp/j5FiS40BX7lEy3yvTg8x49Tuat7hQ+TXcsA0g0H5eOZLtRqzegD68pHybB2GjYNtsu8zHn
8wAY1u30AXPcU8b8LcoR7MQDKX3+KHhcPArtRRpYpS74BHY4qwdtUxu14wKWUIvzp+O27nPHkw/H
OmuoRGx1H3OEsajXwMLMZb2jQHMS+vIoYRDb/HgpDDTH6XMYjY3r9mlnwaHZew5dJe461lXq15gu
//myuvZKwW1FUiji6RNqkfmiYay/ND6EhTekquUPQHzp0sEP2MPxd11boxOpN53dBvB3NOo7xaKg
7ou7taDbTyaj1ljJ1fyoVqWh8RINJKm43BL4DOdLE8C9L83Q++lsCHegqhGnKsWeSUFoZH6UTbJR
4nHT65Su1Y7vAVh8etLaahGLLma+lWWwNC48IewqZdtyk/Dj7m/2J4iom+dcKuvOA77Og1TaQzot
JSWAku8BkgsoMA7abIiCGyU1//bYVa2rUD94A3FlVrznmWZFeB9BKFGrcGFsMgcGfqdK3rQHVfGF
BiOc4sFoXaJKA1fIGuLMCntYoKlzHvYg5QDyRGmTHznwPKwHjPH+hrgpzYhXqkl3Wo3Ub62bk88b
24D6nNnbCgDF8VaxDmR03OAiZk3Epc+nwXAVyhnqMy1gymnAqBycUe5usqBVtQLm9eDO6cNog1Cd
h9aSqAJedjchXki1DZ3ykJtbB7UDLOwCwIXOkyF2apY5iQGOTDqwbjpqpBEqvwk9tEfFNKWVKk10
yOGen6ZH/EShuyEILerECGSd3mRctmTv3gnJJGY89eLPwKX2QsUPI/UMO+nUZwpgIUdZXvhAuCGf
RFOdDiAoHNxtOajazbzvsTEI0AZhha/6uUq3y5czuNSZti3i7WW4zxiCFxw5raWBTgAFtGn1BFED
9d7JMwVsMYX4Ae24macu6zEzTUY+eRV6rLntSAQqcEc6bX9r0LJneuVWsZbS09SZsNx7OPuIcGS+
YTixQmHc8nEZtVktPkFtAFBa05aoeYw74creWnBULZfR5XDWah2ZXg9Jxa4VqyXdcGGlker36UR+
k7uB0o313pF5ySq+gTd3zTG2atnPkJZzpNgr4LXD4mxMyauZrM/w82J4zcDUy6GhvuW4BHkIYIJm
pO02gz7AuQDj+VlXLkM22JNKXIld4/xfOSXtEL7PJSNsmVbVtU88c1jc2ZIMbE91ZN4B1DiQMgPz
0/2FUwCwByiwZEFR5NoqArqQzXLpKRBPdkmERUTUfus7L8rVfPFWXq/M0WpondnWaVk7ZyxGzDr4
+1QgiHpeFfs19wonvMUyZ84wPaghoKGPD665YAoNRBq6H+/5ws3ctU1b7qyBK/29KcuGIEMe2ncg
insRp9p/3J9UbFiQIjPzlPnvJGeap+I44DrDXwDEmJ8aEnpUsYCsXW/j+Cu+VRPQ9yO06C/vKuaz
Vf5Xw3UkSo5OvXFT+gO79yOydK/MXdPFCI+MgFCDq0qAExs6UUFWQ+EmrRUxnCbdFxZBOofLl3Q0
se4pYPtPIdFRJfZpV6wKxc+vVygwIGlbW0lrbTxANsRAzzkAZ5CIXMG8HlV+PJ/LIFxhnOSRjBNX
i8tcI2DrQlct3VzwgualEx/p4F5dx5hsRUwSJQTPYZWxa8pGFbb15TA7DHmJufkhYG2aS38ugbDV
tGrA7AMZMtUGB1TVQNqCcu9dEKDDgeWug9TLV94i/GWRz7W004wgud/zQjIAmAJFAl0hjfhkVizq
dhjRMA4MJx0EM1H7TTPvgA8R1DdgujYPMvfEBQ3GfH2xL+UxMpbfNHOMAjFeW0Ze7SrMRT40T62l
4V/Hve4bpCs0Ewz1nSO4yUdR7s3bGUhm6L1onp82rgC9/VYaM87jaJafXlLBgpZ0+FsrNomgJq3b
zrUaXTDZkVHJWpSHQA+xRouiihgI7YjiZHTl3ekHW//StTWX7/7BUrJFeQRsP7uA+vaEX8wlKUWw
rBwPNL9ZrOQZ8530wtGqCC9n/NYhBuPRX2/oFhlpICe3OE4z/09F+1fgalfKJ6gKaq7qvUc56+ZS
fmccY9fojDioeI9ohwUlY6zRJswMQg+nD0tG+S0h80nNF+BvzhzDiOe5qr2bjuHGHL5DKFAb7dje
BnhrZpvcY77G3UhhxmwCyY3eLobOz4807tgwxMZ5E4rfxEGwzPEUs1pcfGcY9NoMpatEiJklbKu9
O5V2gqWa4owhsXQ/MtwUu1VZcn5aKHbksHtYga8BBxpuqK2lz3UvfxuiM0cnngL6eQPXkvTV0J9E
Dj/ilRbwOSRH6pKIpAiVxK03PVgcu9RJwM3zAs/+AJ88MIVGzU/0ZwVnEW9YX43f48XFjvMXn4MY
Pft4GX84ZGHv4ZYLoiY8NCtgXen49JdQ0TyadWa63QRIab+LkYvuhpNIvQUTkxVWG7dTb3ETRWsB
h7uKrOSeq8CM/hSFlSvCJlTm9YBcPrZCFJjyvMPt2lys48DyzLJDMrMb5QJ9I8M/bj/FBEq1Q2jc
Nr5MN6QY5ELWu0bx3I6OG26ZgYl6/BzAY9tgki/qculXZS1d+kXbxHX7PE5WPCwFL+bOe4RPkd8w
yfuY3XvNW74OCNxWPFJbZKN+MNn4Ry8PpyHUPIrHJx2MXjzChQ0atP6QTtEcE8YyRWxm6ljIsYXM
V/BMHkIom+6X0uGySwMsHBpRTFPHURZ2ZUotaG2OV+UEJnpqqL6pv5wMODgblfzVpeem7P0JtzND
PskzEmDeNOodLh3CZ6pOvoc2aE5C8Y3XypJechTVKEm1SNxz3bspCj5duPlmdoUt4x1QBjYiQYBp
va1Y34G3R+1BYLGyqE3yuVJnlJrRB9652ELbVj85HGWrmuJ44IohjtLLUCOIoIRfH3AAAAw2tDlt
LLxN2zx9pPQYjnLJZpF2+hUPHBVAuMyS9rSeV/AA5fhcDkoP4OMIXKSvMsIhrUm9ozQXUBsl/800
IdUCtHebss9Eb4+76rnE/FuMF+QMoo4uDCEwf4kyWZfwuRjQ1bwNA61V8z830BSF8BKEBhW3Gn3M
tq+UaH7fA6eagMuJyCIyyGeKpnXIj8JnaMF8CTIunMLa7aVOmyYI+F//PXrXxmeyVLwMyU2kQMQP
hpQ9PVFKwwOkO8fZFR1zKPLhX4GRF8dpuP8jArpTb2YiDffrJZaXggXlx0ZEe62zxCS819v+czkK
ee7sqFOf0Ngyi/W7a3cxgNDMlHmYwBsn3qJdsh7aVx+iv+vPxJR0GBlMACCvjqNqqJxgs8dD0sU2
AWcYqcXLyhyMyH5gebUwdnGzUU6FsVJL6yUY1HTKLsh2+0S2N3St0BK+NnX7QhHcAFaC2BU0vAKd
HVwWUrIdiUH9xpPRKRVyc28tpJaV9rgKR6hUX+laJsLcVoWfqZWdwGFTgWmO7jY7ffMmHWnDxFlL
SVl5/5CvitJQu0l1xZBhN0jWRm0WEBg5R4+r20Daq7Rx3c34Tgh0VEbr+QwikCWIpbXh0jm5gIrY
sA5QIOnmEZNqiXNKZ885eNWc/8Yt3UoDP1ETJlCjb4cSxpbP+ZCVhRigCBZcni+Dj3V2Y2NiljKQ
oIMV3eMHnOw7pOVuOokqEhNUYK/528UBVj5nZToQeZ32PwNBqX8X2a4ESQ+sTSQI3fACfJApedTd
IteN9X8RmmftpDUwvIm7FM2OGHfj9d659U9DHQVZze2wQ2n6nadgQS+UMeK5nvGwb+iZGIEh6GAw
5z+qgRpkYSGo/VSqbp+pzGTsSMhYRaN62d9XYBg21BM4WmSjoWvhEZzR02fXmpBFM1yBOUB0gPSX
PVfOPGVWiz7g+WiGS+KxvT3xZXjQSzlqBl0uJJUeuotLFBGk5Q//RsJWo93MJkEJIBazQu0Pwkka
qAuCL8tl+bWbYVmt4D43mSuxonrWwDA6qRQMQ9vngLegS24bF1wEkW9bm6nIfLW3N9y4iGeQso2P
oCY1eAarWCKOJoCDwIPSZU27QPNrnu9N30k49Kzf3pMpHgOOkcuiUqGWLMPIFLM7S/7ia2OLrClN
395e699Q388aqeCNEaGvQ4BHrKZfbOxrhnnOsGaYIiEnh0YnDOzJb9cHT/8DvZEX3qohSdB34gwn
x4g3v0nsYzT7DpBP/4/BfQ0E306LzUMdY5JIe/IBO75T3PhFJcGB2wlrPl7DfFoSQ9XhhYbw5Br3
pCr0u15cUGRSnvdLWsbiFUnLhoPrF75RwipeLwbj1PqelZveyMJoG9AmI8jEyrFS+wRu3BjR4LMo
AyXb1zqrC6z4AJhGI86czBU1n01p6D+Q+wCNA8jzycqLYjO3T8MtaXHA1dd4P+dPJswP25A71ja+
xrlH2TZA2ohcIbNwacXGaRF0ovAARzAbVgxZchZD5WjWktdbE5V3ladR8C//A/E6uVn8zozq5vDe
5aITVsskg02NeIm6t4dYGv0Tnlw9phSLfFKL1/pPnYCgczsagsJft02nLC+ydNVRANUxn37YZira
q1Yz8N5y8at74yTkg+VCac+uFIAnj78ngyFpjQL0b51w2N8zjBc2BbBHXb+KDhlwvn3CcJZoabCK
GGkGAXsQWa5mU+BxEZ9sIkw3WCWwYmdjtdZOrYg2fPtYdpKg06RSPMotVfvimYu3oC2CViMvvAf2
DNoO/1CkBpT/rhVSMIp6CK3Ws0LTbxV2wpHb91ccUIjYQnEtZOmO3Fv/lVj6rW7TzaMBM9vHdbEJ
m45cWKjJ3KS20RQ+gA133ERDTEJRfEUjMRQs5YtXwnSez8PrZ4A/TXGeg0wKuViijlBORyZVkelo
GkRQ1VxqvES7WMZKyoYbO6HTsBPl2T7hwszLGWR6k19I1kfEBVP4sbhR13DMIlFTjVTt70rQRoU5
utzghD/xR5oPEgYXLUQy1+PP1GBVUhS0tFKJZLharskHg7Gye4S6vRkb6+JMOoPwW3WsKc+nwlYE
X6rP4XGyAPqkSzcMIUEAX8jAK8+UJ4bVXYvgjuQL74l8av4zEvOfxHqzpQ7h0jyMiSTs7H3szatC
RYJK30vLOu9TiGqfLT+/s0LGA95hmWVgyO1TA7D/zU0FXrP1HDwL8askhop1Lc3gZADd01YABkqe
U4ajgSNukacNS8mjHBB/dpapcvWYIXt77lucqYxMaT4k3ll6YJ64dWRaS3P5BAdcGKNsX9es4r16
42lq3QEezH0tiLRIl1dz8iD1Xx4ZVenl7WbaNmTTl02h0x4R0G5TbQoR3z6os4mXmlWd2JRQQeNc
R2yFAm4RFl968wj1T59sZqdbZKy2tjC3AO5KQa+Dg9VT1kE/eLe68rHdZVBIRyD4Lgzv3nGWFJ8R
5wODtfBA1cVYq+BK/G7wnWueuFWFURhi8L5NwBFbss0JlP6tVlrrR9n6ezN421cJU24n4hJ/+lTm
wiWWilvMEf0/9pA88umUl/wndh0LhF3Ml+TNwQfGLuuizWF+yMMGYCQO0c5oSOiWWx2Avmh9JHvV
iKVrKboBKLQ8tXnsPFvj6/B+xGalWs6DGG+RTJyneTHVXxUqPsbGuOr89Rs16jk8+ingeoYDjqiP
+808QO8L6C+M5KI0dRCJqaAUIYiv6LxJb/R20GAWMXAy3BweZGpulUc3nHrUXKAKGNNT3N8walTh
ww5ut1PQzbo6BnzRjadKoPMKim4dtu5NLHVVWIOt0ACfv2HMF1QQJODFyT6fdEqTJCi+D9RjVnr0
OYVAWUkFsGkH/Ia4RNUXLSD4AskDoCSE1hwk0K/e0bcHrhBDwMFgAVtK5wjY9cIoQ15/tM+pDkNO
1Av+K5h72TIpx/23QYaFja4Og9NQ3ySHey9Of7ArIitaMxpO3R2qm8NVk7IcOb9XD/3VqpvXgyQ1
JtSZiSAghrvY+JBBom74f1p/Cq5Sy73uMOW1t/FVlcK75z3S2bzccFrnB/zI0Ym+h7CphhRW61Ma
UJaZiDpPpIMoZo5Zl3g6c1fbSYD3i5dgpuu9+cQIpixhXinW5xLn7Cy+BOEez0m9Sv3CY1VfmGU4
gdVkHdlMVSMkXcl9xfNfx1VF+53PohhpOnsAOHQ53DppfBwFK1N8XAE9eBcC6LODdyamsKqK0mZ3
5eb7UFhwjq0dGgNwpHej2dCeYgWFRA9xDezq+Pb9q0SI7OSy0MQ2tMyqAKYzVj8kIgPSMJtH9Ojb
AvJw4ltFJIdFTT4z84vSMZ+JRMHiSkb51hsTsTkqt7+RxQ60OCB9XZbPRf1hNDiLZJn3RMU9WJRi
KKKcJZjXCVPCUHhghBn+rgFOXpM/gJoWvfBTM6rEaK/I6APpbiewjoxqvbOGU5E7TsLVkjCabnsv
wAz1HITDFXA46wYPXiwi1elWJFa5jFuGjkshy9eiDlzGbdVCMkqk3DpMn63qhIMnxZ1fOHX5NrNF
tM0N8GWXsAB/WigascZ/J2RjhQWrLWlktRD73ExVGhtBHObVaEse6zfk19qWHfUUiJkvQMix/KAs
TjF4FM7ops1uB2GYc4EiG93RzzmYGHrNmriwvMYHLPg4k6GPbpPX/KV9jg2O06xpaKp7en//bOJc
W85nSkKmGjOLYG3SFFkCee6OVGqukbdLBjHFQVMf8KR4eAYvMda1ILgQodTYXOXPymwfFSocjVAe
siEQUY8sfVk0n3DeOa/FugvsF943G1ODDe05rVS8riVMeIXF+nNx24moTUkQOigNTofm27f1j8N/
VwOGHnDXWifHExVjkrmsYcBVZgWbS+hJYfv+FDZkI5h61RjXcKCfrLwQLjYsaknmPHYWf4D5bIPw
XqE+GSeazuFYP57IrC2V5fczEHb2VoVQjlwPpahlDMnEzjHlt5zmZokQ7g0ShpIPNO6qYxQLUrfg
nrfdRhnU+5TznaSpyO2vo+UvuVJsaN/BTsCThbwrjNMK6JgJlGL3hnLmac3zItAG0vo1MLPlKfv6
x0rfwyMyr0zrtE6ibcSJfP23JGPS/9e9hhDRrPdrcAKWs/FWWAUif5lPpdFT93MJQU1hO6S2XMAv
/2tcFP8SZYGt/jRj8LGmcspofko3jxodyHUYwk0pWtNyKNNklRcmbbpIqFyD0hcOODUOVPcKTpx1
Khprn1m8ax5tgbps5L88K4gfpr/XR4UhIU13Gt8gnl2/kcfozHCShm1lC+rZgOR4V3J1+IzwglYG
bD3lvjjeYiPETG+s16PCehCt1EzSBcSsro1PJRbQvMkSR8Vhmq1xrmCkQZur72ZGGV/swXGc+9o4
WCQkKcb/LunpdTN/1oKTbwAyjmbI5yJBm3jRLBDeXEi/G8eky35eyO+16Emt3Ce67Eo5VXNFUnwq
QLl29ba66PlrPR22QeEyuR3RQkiAfLgoOYgKhVt15NL8yVOOmIZmlbhoiAdCxkcYXcadSnwh+NdY
mXzNg5EyQwTvAM3hGV0HezzZmlB3npeInF27PeJJCyhWF/ouGx30v1y+00JyQd8bRzYzLYl2vp8c
lawNp8u/9NiEUNXM+TyAscz5+e8vPwBctTaqNcQREfnipm3GOspF4rQipONhhOPyeZa/RFw/mBeo
XbSyj8tzFE2GpjxgP/nL26cenaaIJ1bd5rgJ7WqbFuRKdjR7E2LIsmF2zgI7QezZruWjfE15hx85
8DZS5mUp0JXH4uqbPfYbK58inK4dodQcw9tp1KcvQpJW4z7+Icny2OC61l2kRA/fGmSuJnEOId2w
Tpfion5reMr5d5EcqmGVlYoY3KeYkMlx4VBpVHsyBv6qWpP/vLgznWCQ0eZv9o6v1wtdyMxDlzGk
fVsiyyoW+wg/DdoaB5it6tZY5BzXdmzfxJ34Jfsn4yLZoXDydrTok9zarJOSvFH644+Y2fdBJydL
3Zz8q7G06rH8+HcL38CXeYM0I7SU5Rr8mmZAYi7oFr7oQVuIiIMC2l1CvCm3uejo8kkXbSO3Ahnx
rzWQhscECte0zrzijxPEIp6BNZ1zD8X4UAHfJQIMFdFh7q+ZAKQpJJwVNzQHv7IoR/vh0MKMvq01
BrHvfxruSeFW7JjSt1dYtQ58FftQNPPz/Z4XdflOlsnP97H5wU2pMwIfeSOJj0nBGjXmMWnjpKxY
vK4SuUCpo+7izYWLO9IQQ3cJ7YfV+cyqLvj+gJ1dufGuA1wdGxvlUgF6hP9cF2OiHRVu+h6k3eQG
qsslMTB1prEXIFWbLyEc9pYLOaDUDhBU3KdcSNa5E22cM/C7OgKlXP8DMaQqo2tsz7dgBGR7Gi8m
6Y3SogX+jmhH6iBO7ElMkjVmzVqBbpyUpLg4F4CIVYjegREPvcHR8PMifS9xaiIESBNVMOV5OZgj
Qcs2S/DZXeJEh69BssMKYKTcmzG//tl96e3iYpriw8L/4kLrP43jdsZ4PDMmK0bceugC2pZ3mC6z
yNtbfHh3pl7X4lylFdub/G0CY2KXf0MmSO7x0lwFGJ/fSuLXh0K0yldaxsmhTgVL9NvlkoJsb1Dz
jOqUWzwqAfYUN6mLcTKiQiJNGQhMhk9QzfeoghdthJaoIVum711jEtfdg1fn325ZdHgqwNJjd7sI
6G5S7nP3rbu/dM3r7kCQBJMX5x7GA5JxAC70n49xiFTCwrIqHThmTrP7Yk30YQvVaIykF5ygohJ4
FAhwKLnO+lDV3uCP5BfYjbG8vlilfkUgfiZbsqV2ln2564HQVyhSKxTfYAcyhLVMOCCiYKDqeU2z
ccGNUYGRoFaI2wua1preZZFZCltYAP1/6wICFSEo1eb0K4Zw6pJw77o0kfnWtQOpkgmKaIy0yru+
iClAUnNBMTYFHFHxJxegpMnRlOlK4mXDRZFJsPAu7e4H93XYvAQKTPEYLY+tPlyLIlWSUDMDow0v
DDPQSc81MmOckGUJzB6WLcs3ROPjCeEwBu22vzOzc+CuawusAuB8/WC0xsx6Z2N8jiVifE76cUap
fxWv5vuxdklfSxVc5yI3j6xdD5CMldsjxgPHUGG9uym58tx1uJT+P6qEkD9LXeSf+rzmuRC2nffT
12Rm+q6fAh2q+aesZyRhyuSZfQ80vOvdjx/Xx3VS/+boY+jDJ6EA00EhVGmzJAHDrTYo2dN7yu94
msfhfttKxTFe65pp+jx1Ke1KmLlgcQY174S8aGMEbuO+Ze+R3K/kB4UnG5fr83Y8Tj6PJd6OAUSa
G0Qq3REkz147p2Mn0GiYLc05DCuYZuUhmNNXiyK6sKaBYMJr14lNZ1lYlJMEC+sp3TN4v7SNCf9e
ToTqAtdUo/UfR6uto0SXT+niv5dfBFMdGi34DEURlfHaIoWsZHp7UNaktyzNnlit4SdSdY/b0IWD
lUKwMJhnjRwd9UOOqlMpSWSnygbuEPqLyCjy0iw5Orz62uEblMaHb7nwxCNmHbjE4WORV84gIyoO
/4YdToGxprnCByCcB9PBPGtSLk4lzVMs8XXO3BRBDaisEkn9CMuc+CuJM/cskE+K/EOanaVgjDVP
v+4EHTC3y08CGgVPvdbH3VUWvajkTr+J/FCnOA4oXFjbS/E3pOVNHjG+bn96ReqgcUO80+ZCanfd
eQD9YS7xq3GJJohFlwrv+wVKBoBUUMuGm4+zSIwrxOD1c5O+w7n/VGuETfRF/aJHj/mKo+kYkOp9
E4XgC7G63QZ685IloBpIsE8siS8jtoukHlpbRZKY2M/t6jMXgX5EX+2RT6c69GwDlw9MG7bWCRm4
aEhID0jYA6M+SIf+ibrP7KfJoTZevfq+VVuhCtMx5cQ1TRvGIN96fwD+cty1kUNRjkHQxObaIKdb
hlC21UuPMRpmiFGPNtE+LbdxdTtGoG3keq9F6t5tyyC1AuZezN0vA6B9165SQOr2iqU9ZVI/Maj3
CKu5sLvAas2qrgYh5AySMvWPC03T8yZu4I7n0vA2+pLJrpKIgnlj9kkhDqTQLKCI4tXdOmLhIlg6
O5apa7PJRGj/seBToRdceAJzTrcyKGtbWaRXS0Bd7+JGOD5dTxkuirE3Aq7RY5+8DX69+C0s0nTo
UMTnfz/sxKFLVsjTCmI/25QrK3F5iZlDQbFSWETYnqN6MSagAp25eNTedZCTewy5MdZhpAigq5p0
HDRr4NHn476RjJPD13NliIdp9kcrQWqLy7gMWy/0nttODEanEiKRIREYiLzLJ4J/G5vp0eSYFjEr
A5LdGDHyxsaehEAZiat/53nK2cHu3R6Vt2iMlxw4fl5ywMFAr+tp1VMWDl+N07L2K/xAj4PmlRs9
bGw7wiaW1Lye0Y2grs56xdETW2Lr3vlCTmn0pae4zPWq7310TNhGWXvtHhXu2drxgwFdiYyICINd
LWcgVjpPT0InFoGkZfLlf4cXBM0AKYctvX5IK1vDv1FdZ8lDg1mulYUi2OuSvxAATCoX8WcEiycq
BMO6qSYUx2hclLXX/eJXl/8pNk7rrWL0kvCvSxsNxrJKG6C/JI6XPmLdkqM8AYPNYdY0PJa0GZ5W
CXP3n7BJzXmgBSVVbHm0zNcjddatAGy4L8DsqCRrJn3lH2rbF0OCy8Fq4uCSCYjZOBs4N/BsnGQi
ieIeA+22vg93f0jTiKTBq0OGuutaCruWoU3/BqtyfA9VFl9oRwY3s/aNhOrqRUYY8ocqDWnI0Nge
MbhZ/EgRpjhO+YZaXhsoVKONpYu9jqrjcE9gCtseso4lNfsnOY8zhhskKnBoBB9GPNbC0Bwqxcvm
UrfgPJ6c0Df+TC9snSqxg0ZIRXFNt49jOYb+Hl9kFUogZmTXRjuWJR5D6Y15bgLem0v5IrAEYuVU
tS+ReBPAZth9LT5A/vSDfYDH0riR9afSRGGiPuBQwFjntWPTytw2BJDfN0mezJb4q7HR8bNqFfl5
xLRQuwpulU87C3mSGed0Ym2jo8s8F+dzNPsUGq/N9FlktP0C84IJ0BX3tKwyjX4BOCTRwvWHEJvf
z0Sj+rPGw5fU/ChLrq+7dPPfSkB+Fvce2CNABO0N3Hj+k9U0tWThGkxGNDrPXDIESFEPIGoZCmXn
M++fHd6H5SWWPhHT/ySkcALKKBCo4Jv/bDvykNW8G5vsoVDLPVvye8HrsfVhyymrU8OqDCwQcSe1
W61CGhXiBzyFn7kFcz+wToYkjwPXtU4dP4FJXsi0tZaocbjWeIvU5bP1KiE/clHGlpc6ZYv3++RN
sQCuQkxUKNATcvP+Slh9i17yNBlAYYgn6QvQxoxeJjbkwo0r3KvHX8btbmwPkwEa8jzcY/tFXMxR
sgCDqkbSy+64pBp8GpWxN1K/FlpiaVZy27ythtdpDnJI7FZT23iCQvfRodO7Iezd409y1tLzB6OB
ho4sPg8jbuLaajW6jEOH3yqsjuYiyNbtlTPCo0jxogUZ0pFqqdMCa2jHv6oKaDJL0Ny9XXn0d4bt
igZxrzICfhwb2i7mpHZDzsi08/ZfPSaKSLUs3d1rW3gioFJOaoUK8CRhnIJXzag0kG83c6+8UXJl
J3r9XTuuYDYtQjVyB8u8TNKRHqnT8BG/nqTtcHeKYTylGQPkp3MpPSzgZ/7TuXE3obckQJUncBDc
Vpj0n9u4we4hjaI4qAdpuNL+sXI3yW8ATh90w3Wbnoekl6mS90YyguWKvPN1sZl9VNyHybp7UICu
rbnhxPhS9WTGc56Hl8DSqpPVA0gd9anwurMx/ED2EHOrSLBHa4iJ1tkQAF6TAwrL782SlD97MTNh
TxNmAHAZFDDJJFso/39pFtgKjgdbHvhJIgGdrF0kUZS1k7y3PeV1yWUyTyDMF8ENe8JshKFi4SU1
9jvUUTwep8g4bSAyZsNC3ojlF4u2C5yucD5hKvun6D5w3TZIfsX5o/UUsnnBNT2q7rCMm6vnB13N
Hokp+5VccpqQLMXxhC3x1ORFskealZaRFOdm1JzJD4mQNhVkYx8oBW4owDBa1WCCQPxfAA2GwzP8
/BGo16aBxu/hTuXJcqQsR0ML/syB40Cgj9GHCqOI5l24tCBPpuuyWIPsKIscSbZv72bYBENh1RLN
fYqkkiFMTqp0SLFRdm6LwBX1na0UQA1zg3Y8l8E2vBiRV+VZDUzkHcOK7S20+VRTY2qbGu7saSap
VCZJaI2QcWFvupPJnj6cUd6qMFjmlijLKqGcuiKXfXCwOfaZr7oO9XUDBTbcfhCLaqwkX2A+Q5C5
gBYQLUEhweYg+Z7OFNpjRk6A7R20b2QHeuLI11y8WUMtKKJP5g16yVzNtVBBwNUsj/Fkp79xoU5H
twx9xHYa/qr4BeI9sTsMyhO9WbxkKp6SEltywdkVhsNf8unaeYUl8FkAG7pLXwTzuYvw1WjL3/Q3
5u05xwLmFaTh+9hrr18g0ihxO5shs3j5/aZ1f7jXq/QYlxzEWqpgGa/l1ep4doAy7tbrFYRLaVg+
s3zVIo0eWRssdQPnx8NGEBVfQ4F9/zHDzMjVSJYWZJc6Y6ouxbKKeJpPUxsph/haZT+liGP5+gFB
Yu/kFdUd/I5XDoHoCGvfSLiZEFG3nksCNxiHIXBgIiIJogE7le2aaTu5djNREHQ61zCEHA5K9hw6
6jMzJGtRVi3WGQw2ygzncwRljWvEBUq0RRibj1p9aTxgmhRRg1JxCDeqWdfCqowgKh+3NbVqKous
WTvrwEVJK1jo5ci9SwUTzd4VaTZnWAkjv9mhn9MciglDQtfyIFBxAMYTsLtNY+B29BxFj7BcTRgl
WLO4BNPa9TtuF81ZxDqS9pRrEzPqd5sajfc+qK9S4g7aX3oxDHw3ITprAH/awAVRBxg6F8W6cLrw
/ahkPgwZk/hRoInMebrPhOskNRUqXvj2HrM3uMbl9qaKqOocP0D2Rg1pUlLQj1oqBwpqLSnmyeN+
JG7cRNXk15VQ8VfQHUue7LP6a0tvPKZ8/UIY1mj3Xp9bLSRwaZ5V3kSU8Xo6vhgqSJvM88bbXBpP
bTx3CwZkhcNWSpPLkEN7CxQHAoPoMm716xWgHhJIKZCZTHEOO80b1gHnvhKsiXqEHsAGthvy0WJH
+oyi58tBhZCXyWaBmwMYOaEBjunRlThWly3anUW13AXm/5PqcskipVG7b75Upy8/ZwJ4EcIcrDj/
y/vFYQUD7EFMB2/tZbZQ6SbzqgY/2/HpITQ5djzzIa8t+0Vi2b8uGz244P4HGIREdUz0fRVktMPS
D7ggRJPWkujYJjG1VZ9uMMy/9YveFcdsAj1cf1qbCzqdagK/gHOXPyKPG6SGNB5ru7sEH0J4fs3o
6nOTw24UqcW2RECRDSMWIEvhcI3b/cGKAO6AgGR4iStwoZMI3a+r7ET9DTR58OCyPT8H/L4OWd7a
+u8vcPaM3+Xn2g6qQ4ynjN1tquUJsmhM2onZnvDj9O74yfuiWpUpgNcnGwN5pAYTUBxI19KW823F
V4pStabMR7e9AQOA/OZwa3xzvS01cg2R991fAi53FjFV2OVmo4YMDRzYLL7JE0rb8VU12Ht68Rx1
Xpftblc7aQNDZFvnNWKYXbyYTSReITU83w/7uvY+If4YhJO++u29ajNDnbXtYPtAc4NjAvVDkyfc
QXWY4qXuFdtEoRSg6YYZcwZLfrsUEcH/abxcFWwGkgDqz8Wvnl43fBl0j8OYzefn2vxmQDjvKQAL
+WqmlORk+XywQfHmUxSuz31XWzraNZ1g44vxg7rcNQCYOOFgfJomINDvxVHphc3r93eLKmEtV8MJ
jQaH4qL9W6fHZ4pfKrwXoChSTtV0DKev6FyO5NxhPqHexQjTZgAoLYYh0nbIDb5zlh03Cw1sqRxK
dM3JeUv67NHgnh3r6qhgACAvotP9WOf8x62nxh8uS7xKEyEe6GP0rZk3rEpIHwP8hbZJ9uxY/NUg
hXJgnSz7n3+Ic2ITJjq2/m8w4CUVdBMv4RzaHiFGsgvXG7IFC+1aAjVl6d1TEjUOvtDGcMjR0JJa
XZz8avrgwt2P5y3fOEzsDaEI938BUB391uTjn9a/vzzSGeNqvuO7x3k125ttK5NfJbo/OdXaNMnu
AzYURSF+2pJuNo4mSjGYAXleUwBeH5pSS2U7ZjJNJOcv8CYLzI5HVDO8nUfEGLfMh532WY4r7Ksk
oR62flaqP+reQuiWIXHxpiS+EhQ9m7OzJF18lKwVFXANA9RPxeEuk4vAmVMuUkO+tI6MPEmRYRUo
jPDCH3wzNvvk4NVi/15ey+7KiaPeDtPz9yXYquN/7npHDH5/U9AsBAFZP9DT56qFpbqftlWHlBkl
pzYrBEluXJx1UXNMEqOWGJJUC9umOMKIDK8wDHEjjCFeHCQc05tWanCk4ww8LurmyAR0IlY8prjz
b1vG3JUrBfasy7a8gSzLOmFTfQyz8+YjLeRJEreTAVPa4bnjsHwStzbaRreceyto6Hr1fyejlyNR
jj1NUaDo5Tn7thSvJGvxMVveelf+Jaz9oUX8FQH81uzAUdYJeQEzHZA1I16OuuBgyvzuN5NoxAqQ
MvV6M+U/QFJiJq5JNQ40lat8ctE/Ifh4Mvm7vnkIXqhxgrSGrj85pzq2ARp9r48ABA3hbt1R4xsE
c6t4XUOZToBgp/drxpazX54I5Dn1625pPdjUVdYHRsKNGP5aaAhjWgX2GUvf/TCPc94m12VW9vdt
UBj8adc86ZzgmwKaqaN4f9HiXk1P0VRyBRR7Zn7m4lYzZ6owe1+ru9XFKAxKISzGZrf7v1V8Npw9
QjGLql1hPyNDvVbP6475ewK58t7YV9Q8oGAVfdLZDHklyFNpGtfBQeFXrjtr6O3givzl6mAaqITp
R5y/KB70Hi7pex1/3Bt5MZbEN3DOgRz5P/oChmZgiYQ0scSXNK4eT872Y6Xxe833rW02pzs9QOby
cJmrhBSST0JVCfs4EIwtgnb4Yot+AEzKJiGwHmLdi97tG75n0OPFPPIcQlFSW91vi3PAMal9HJxO
VQ9AHg5KLz6x5GszthvKry/h8bBMN3AVNk5SzfCFrzJflj8Y5TZrSdzMdxapTrWiv/UKdTBCRLSz
9rcYzoulIYgpoRJCx7Q4pQ7YsTGsB8LeyttUfRvMYu8J4T4ixU6X1eZ9MqH0aiHCoPMqgSS1xkWY
XGrcYakXcHV5fv21EgzXa2V3Gq3c8+jMRy8V1Cn5T4ZYi5OpF7dklaaHcWWgXTtJHVTglYiyezpZ
8dbQR88gwNhwNieC+IpxboJVZ1VaiLzYE6b2UjRjsQXX18n3z1WLdKFzg1TCoV0USRUkX9O/N971
yzsWjqcGK5ktXWvkNgzYuu9B3AWgWCUQMwx/30CL/s6TgzCSxgGA0qyDQm5vYObWsGG/dU+aK8nz
h2pISRToi/VG+Vz2B3Ga5zq/7OJjF0PAMc8p9NBrGkpd7IMd72YNx04fwa0dCeAMcf/kzSribtSB
efoNSeGn/h3yzj6LcETyAEoFByuhzPRxOD6zLf340PKcHDjcCcOOrg4ApU+G8GLAepECla0ExG+z
SXMaTifXG6neqMbBGriHrZ30v9CQrAzBhxiKcbHkX/2fVLrvVECuhcFoVFRCYtj67Z7MYoeHVsqM
eStOaqBMwWywZXZYpa4dwF5tHzIJjggkLtrSVXfYgKXUHEyxbvvVBGpW7qsOl21brux/tDzHXd9w
pSGi9TRzZ9sxywjHS+r6H/NaLpOHN13L0NJgEd+frqVGA86H/v0n1z3cPBwP8Wkno5/7XvlcPadB
kDQlezdh6/BzLd2A2KyrxO21JhsebGYil9thXsG1cjlocCe9W+nfg3g+SN/f+PdR9JRdbNFNUzbo
y/2xcoV7kjv0n6577550ot8I2lsyZY9ysRzI2ogZYs/cJ/XSyL2JTsUbmLbwV0NVLKLDj1NQ4NV5
wupSJcRSCavZgoYfys5QRmdHdfYfZl8qpPE/1+HPwF7cJ5zoNoFkuB1qM/L6h9iyByyNgC43rUwU
e3cXeYRA8bJdUYzCYNIolAGTD6+IP3upPQbXo7FYYyt+Sti6baJdnJN1AkDpKGYQmiMdRmuPbtyM
qYtadI3zFa+PRwEcLLckHqm39P3YbenVtionqf+aTd989Nz2ci4F2f5CMoQkhJ2mDGysBfZOiZqW
QN0YykwxgCJF8K4815lsSTIaZ/jm3kxkpC3BsADNnkUiSMmgcCWq5dV53yyKxL1UU5C+/3eXjCG/
nisul1cOl/iEWnPJnDfnhjFo3pf61eygX669smvjVfsnaLA/yQMdCgIUWlLVKIr64v0hL1lo0LHu
214lbRKo084AsmGt8PET735NN6VnobM7L6QUuffLp+57JUmRfis28UUpmRHwJ7XAGirrW2ViNNdp
e2mjjT7IxEv08TNWnE6NOb7TuCiNK59YCuoC1Dm47tVo08YrnOmPX7jlOI4vXJIHV+k/js0fi4Ns
Nbl8p6rp0tW4sEhWzoK1vK42knuyv14YWGHO6J0jPoHX15aisMHw5yGXsPTF8jqJVQXmswSDf+wg
1DkJ8POBwWuhruKtR9lwVRyPYcg+0bdn10zlz2JVPnkggb9v2h1FxWnl5T7kibNBe6OzyxLG/Qmi
F1W+VLGwKacyfcymPXotBEBS6JeE3VsjUpjdUPGjX3q6V/sk75890nwQV14F7Sad6H7KUPUHOg4k
IL4P7LcBE+hy1jSxKdCVp+bJGvma4hqpYThhNbBW0Ou+uzVihj+jlpSLJLU+2ZoktWHsZ321/Wdj
i9DNGFG59QvCcnexCh4gYn/4QsNUBqCjc7ufmoOuY+OyoE04BgyKE88RhLErArXQIWJArlQWW3G0
1NzngB/dlrF21iHwpJ2mNBwDyP4pKrgLQ5GlHIbz3/soL3z10rSbPeXz2EdEweKS+iPhhr0+IZVJ
GTya9tcWH/PrS5MSRINK6LW4YEPzVBSaY1XtjA4r2L9ypRqC/wTVjExfcbW/YsLP5tgdG/nh/oyt
mmbsCNP2BFT8I9RAcHpG5tlqEP/lxe4gg8dvZqI+IGG4+J/TbDppplQ5l+ocWKOA9wCHu2QUIcBE
Elx1Vcj9DzF6gwWt1KHpJmc8SvlISksg+vD1cPhwFz+Hei0fa7AoYqcey4xfTU82SlpydPkU+gdt
q5e5kVuohBQSsvYIMtzRFhuZsmAR0x/ak3y8dc1a9bJI1Q1ZMEU/ETVl+jcRESFwugp7HHGe2Mnf
ADn+x36r1O2tnwkYsGUdm5Ig1+m4jAWMV5lgXtkL2D9zZnThJpQu1WggV7N3mJCTro4SpyCBuFdp
LKXwtPzUDHRxCNpoHza8/Ds9EUulbwKUyoi1kSctJOl9gSEu9kfSrsV0UxVjqTh8u/jE49VfMVqm
/G0DoGaND9BmrbWJ0c/TOzvIKjvkbalZlfCYwS/nHCMm3KKJ2cWBkfg5w2VwFZmriY7iVikldk/2
RT25h2YONBuybiQ42IGFYsEA15qbbRHGIJ8lFPc1akkd9wrz2+WcI7VCj6i5RQLPkuUomRYEKVx9
+sYMRKvI5VpdM3E3MK3nUdLXiXQmfRChew8w7ueuzLkEJKO30Y7QXUr/iCHa+VzKzr06sxRy8BoA
5XSalyCfIbLVPnBMGMX6nQbmEysT3N3lpJYQEEHRZGAc+hdctKKek4rqXoUbIMK1MQTAxmmA5Xb7
M1FF9lNch8c61XfcUPoeQPjB8ZOYdL4qkfj/A3Tt9vUVT5f9gxcHCvAUw8Z0ok3+53QqXO5aIiyW
wpiSVUctbQZen31CHicGKxE4rlNpk38KXZI4Oul7sqMRyPb1NgYED7DzXmnFGPobudR+xqJoxWqb
aC8SXMGrazZjLr6r0jXsEfeKeIlk8YkpbJZCE0mxJ85S1lOGvJFxfbIWZPHOEHcbP07Xn6vS7Am0
iMn86Y3IP0JYzC6nqY4p1Q8YuT/9qu6Je+r/BQ7Bz9ETvAQTKYCCwNnTuUYCa/zN+OgwVk9tDhTT
gXa8QrWWVcl3tA/lunMkYjBY6E5E2KFLWjDLdQrVi2Vapvvj6U/u49gsTCz2+KmJqs0l7Thm6ge+
g4VKQMpoI8x+JqBbq80W6uQEvRG+dekDsCV+WlB2JWHLcX9DD8StuH8if6i4iPf+0AnhlscD+rv9
/u0Hq+me6XHEPXBkmK18A+kZmPLNJpxLZMbRAtkcuTqFdbLmUajUlMSH5CY/PZf+Toc0/4JWZwVj
yLFOfT4UPi1XC3jU9bwNV/xpwzfgtQIstdqsYC7Md5Yunki5sBPGdr5acg5HYTpOVEq43EtO01BW
AStqzMQMYdYkS2pgy68ZBhPAP5QhnTaqomR1HDFHMcE34HEmzSeL0JH2Jk+ie9nVNkWVvbqEYgXA
dmQ7Ch0b9ls6ABhY4ap2DLwR0/v/UNzYlz3CEz6aFicfQuTA4BYL4GoHlAOcQBh8M6SgpN+lHbnR
Tzv/7b4/N5NUsX0Ud++P6qpIi34MAZqhjZaT6q2Q5ELHGOMQmuHnxF7Gvr4ts/v2E3td7pJNSQFM
8aAsQureneTIhO19aFTHVMPqrapz1XptbuateEUx/AB0ZEwdYTG6Oq6+KoSBXjhLUMKWRpl9+gwu
5BuM04TCgfw8tJtAL76/c1h2yQ87xp0IXICh58jyyEpT0ig+1dxHjn+3u3hGe7dbl1E7vpWcpqwb
qMLG9hvlA/V2X8zw4MGD9MlFqwMZ36LHtEhaEZp7yHiuf/qkxe2Qclyj3NbzRNsqBDTOK5pYPrWF
lKn1U7uEnM8rKqjG0hbqENZ5NPU5qeAnYSnaedM6LQplpMnLJ7lMz6bf7e4gvYt6nbxVVTps36+l
p8zzWzdZCFdq8eU6sSZjPigP7b7dOp/J8GsgEgafRvFMh0yJFBK22DSzlCJaXfELW5BbWWnfiyrL
pWmFGD8Sd0EyJEVJb1aSwcMZEuuJ+zE4ljXMKqcKjdZ2E3VQqMHgyg+y4jcOJ6jxbkd7y4Jq8brn
h+YrgIn6AtFYNzUek8+Evdnd23bmmnEuedMJhPa15YuMPEgaYW+WIf/ah0xMNJ5kk6vr1POciFPk
fa/yF0kEY/3fwLRz5igKwJIb4Zx/MIpQUD6Lf1obVIbX4dGJdikk1XFflY5zL9mUHPw/XPVIwhwX
LrfWF3b1mpWm788+MFKjMYKbIRrE9FfjKhc7i3o3BWoG8h4Z25CeSiJOCm/9fK34iG07tNhAVsCV
cSSUCgsd4jx/LdnP8sZM795vpXLZe9Hjxj4wq3KIeQtwgD/c9JqpFKuO/HmMAsd83jo2xmDFUbgZ
V7y9L0hHopiSxJNVGOidXaaASRQd9jPLYaTRyf6FSEZBYO8xHAERfnnMmJx1bhkv9KL5n3379PGN
ci1S/zFoHg4QxBTNKfsfpFkCFD0RFU5MX7eTlZiuRrrlEMlOa8w0f3pAyFcPaySwEn2RMPWzZdI9
0TaOCVsiuwhUxuwwQAwS9mWliP4YhL8jc5KSPLa4fVa61leTJsNK9cVgV9ydV2jEYosEdy+wzK47
kTtn93v0kQe3kX/Z2pWhSLB7XxH2Dm3d9fq7BygYuBbP9LVl3gM+epwKYTNaQOli3WrVnBUOt3iA
kqh1svzL8JR0keLiSWhpvhV39RiSOnIavKeLB4Efx64HEAdjIxJEdZYMmzVoXyBdmhxlPubZo8Lv
Z78pJ6YtyJEiKxrZqsC0MSEve5enAFpng/zgBtHVsRbGRXDFxEPbp6Kir/GqlIKb/RnhtlH4mRUf
G8PgSKb6Ajxm9bMTRpI/qa8rQtDHViyoE2zflmcS9LdqdnOkxZA/jLqTAS+NaWacP1zl6CDtuba0
BjvDaE5a52XfU1FdqYZclkBbO/WmqwG6NR6uMWJL/LE0xtDIHOahyNPPdvvjukk5ZGXdXQdEC46C
3klxWLyfVAlXtrJbOll/exHZTSKmSoLbg/AvI7/TjItXXROwcFrW1BHyWMpDhHNHXR1Q/5C0jWRH
sUne5sU9EAHNU/kTxyOiAr8h0MJ9Kmo2D4M4LIyddK/IAfhflFI2WmrRYo/JoWXqI4WfrDY3jacM
xy+UvYymg4fusB5fbdX3ph8q1cHPAauMiIG4YToaPBnIEgcetl3gtnpF7Cv1Qx0M3CGRFsg2t/GM
sOxMz3zWHCHfXL63SJTbWZJu4lakR6Esw2R64deAXSKgkCWldyJfwSla1JpmThxQYdyRxr83QvIn
SS1VB+zHhvzl4WLRad1D8DSqZf+EAz1hxvH5pvrJImnzqcqIAySvD3j82xcvd5EBRh6d4k3GI1b4
sd2zTG0XNyRSzDZWnaB4bAHnWL4fjV0NW5DjMl0BzOIuIRG/MOVnctmL7Q/p32fksZViVUG8XAMo
v3drrEBhbnW+Fvn33erVaKQ6OMho4nEUJsn+NH5H2M13ZLXu8q/xZBgYKt/jT84EqLpqBZjrfhlp
FkSxtEVLWes9r5AsIbuI3sdQMLx4LQC9nITUEqTc8WCtj8jnutjRe7AhDx+NskVkUX88L0Ua8GeY
XSqoufsOnkrCjL3+mohGGrUQb4uXcK9kiwi7aViP85ykoAYuKUlGYYO/1oArSDRE7rPTjeDgicpn
ORonedxS7YRlWTQwMdzHDVB0zW0dFu6msFZ0bj49Wf+I9G1wYr0ShcWfmneztFOwZUtape9ozCRz
4+O7OpLt51diD/7rFS5ADYD0+3wrh4qc3r4od4Ac+c5tZ2VOysYSgL33Vl7vsOsT6MEvW+CCjKoC
MekFk4gvH9dLnME4lHLV9QmH2U/9j2FEyBdFxKw6ZmO371hL82LaOwx6HQ2VZTm+fDvyU1+sod4U
BBBtldQQHDwlR/o2rEF5V55AbB1LWlYxukiqd1h7St2UOmp5G01XgaNZW7Bt6PHf1RNtmJnUDXh3
gHOOOm9RgEROHsZa2plaMTsTyqIXDtdQx1TeU/cHySpnaYoAymSgdXoSX41h9KyER1cmPS8YRqkv
6Gr8/I3j60emUhW8xKj8DqWEW7fJWvpuGSEdER5rLaQVWxeNfxWQ9K6HFPtg2IDyOb+FQRzXrWBA
rX1gmHVksFrrLuAtlq+mSMqmYtEZjwi16VqfdiMKZA+4oeCc01rq8thintX/Ofw5NZQqlJM8IDtn
CG3Te4MOkviY+N+UIRYPP0Svl36/bt4iiINbgiUox9aipA3bmVJOR7jL4D2ZCu9ud4d2Er2fV9VM
W/y0mTZuwljthZnqeOtGGm12IdFo1a3nfU2sRGZNZCH1XIvuUs6ercBkUInKGeX9GF8a+yGB4FKE
Vgk20RP8NeNmT9yZWimEvuihIerRrWXI3p9gx2JHrpNAGmSAlHr1Bwmoax+w8wnmK66TheDhLnpT
DYVGuZPrioIp2CRHSl0PfsguG4m40oEPBXrcL5PgttH/+1w+ei+DHgg9uDOzYUHpMUsIWHSBbqOw
N5ZUNoNn8gy5d7WkRu5S7K2v2QNasaCJ+7uM12MQjaUE/noqHBT501BzsOYsFgN2rDh/fBf59NB4
rVLsJtyRPXZdolucw99+i0PE4ImKOoLEUpis3vazl748SE0hJYeFczYCye60Wy399Q1+I+Yu0tho
2Ai+W6rc8SYI11T2TJ79T7gzRd/unIcpFt8J1bYJUVjaTRy9rdhnJ8cluw+hDdvoyYr+CRwTzEuP
oBITeJNo8ll0abT6vk0ltow2+iZKclqvCIvbvZvVjulyph5xRJXDwr/QnBeqrOwjS4yyOUY+ZQLm
J1K944MdXIodGkugdmGtnxSR+9u+FzqWpVy3JndBAsX6oUGF+fOvgOdQ2Vevyy/MLOuB5Bdi0QwH
vUkhwz4XvFMcx+mtI7+DO9lFHe2ZGY4ShkiMPBegtPQ3md0MtbIYbafyG/7SoTgIzM7cU8cZNYTS
vJXxZmxSnGzRuUO8Euf6qwC+6xsTDgJymA6dVWfYRktriU3n5JMhfgA/DJOODkwe3Xo1JsglJy+8
1v6wB/AthX3ewHpqDV7cfBzxDgIPMNj3Yd1GgGOVq5XF3waXlgxLWYQOI9yGVewG/MpV89QC+3k4
X1bdCS4Ncnm0e5aRoUq8H5kuUHIcTUnORaKv0HAqRlk10EVWpmaIrERXQBgLiHOi+kLe3BIhtVGC
pTw+enga37lO7XWjrHq0ZVKRYd9rrt4ICProxH8bEm1DIzmcbwAWb1stEkpEYXSkCxEMBC0+tNor
0c9oMrXXxYlCTnR6K0BziDmjX9GcOBViGStT9qggxAHbHe4U8cJMMi3Gpg6OumiQjbAWlllo2QSF
xLTtGS5foGa8Tl2a+UWokrjxhemVkVdlHmj2zol0HLiPhKPSZbv9IMyV4eqtmYkDTo7IfC4Er9dQ
s9LyIfDZK7V/bxvmmRRB24TG6wNkXE+uUMDhSikIyncCqQr8L8hj/iheo8GYgWQuH/tNe26ea1FA
EIbq8Rpvfpt8psjz3ilW3nZDAaacDW7cBumvl2XrCp6VNh6doxpMyGVXsDL3YrMKHfYhvIROeIYW
XgwKJ11jLznUdzDXERmhkPn9W4/I2nfjO9+n5kJ72AodhMm0drHY4HgOWgxw8Fgxp1Z8d+dFqSbd
mfzEMApKqIKB/02YKhncB6sLOp/0gmM6Kx4IOpERRQ/JdDdhcvPo1qow3lVYGjWS0nOggJanvAJ8
cRZIU+NSFUNDfOVjJU9nWf+trq7OPUKuy+fplz35V2h7/PPdzJcGYkXUVPT5e1MuV5KgZCyfRpRQ
wqIiDGpzKMepJyJ6/Hl7r9AlbRYWeHbnowZkh03vXxBbRy/CsgFrkQZ0xkwRsSDIViJqWcYzaFap
G8Yp7Tv0LqCJsAFTgXafheLp2lCA+wz46fEFxTomUVc9iV+mstNujPqoBcRHyS6UJ+uAYRcgNvNi
Jnb2CGiIz5SfVDvAWshIKxELGwcZhAofgfdRcrYgiNhc9DDozvG1klq6f+eWxwhsXVPG2WGJzJ1c
6NevOITEF5k5+qYU1MIM3oJNmhjrosumqlepWLveijDy5RN2XSwgquVYOJa4eqTPDk7R49ehLDa/
QsBmekJNwAQHWvpxcdn6edQvmxbFRmMt7jwQXet2FSjOT3ieeDPx3WeEqXB9EJvFXZN3+NRwjR60
0tvkf8TMSH9N5aGxG5236nJ/xhT6Dy2dbY8fHg7Gnc7ugipE0HDs7f3Odpt1iPY+bfTO7djWoLsJ
Lu3hPpRN+1s9Ull24R6KEX9Z1f4ZGzsptSLDrMnl1gEoN0EO5XvizT1gCBQ+2QhZsV3oJJ2P7DAi
44JQlAeeB5x+0yZb/YAbWxMcpVA6ctwqi1gL5Dc1n191sOvPq6u26UhERl4CFIsG7OCEsaKpYYzm
SuqNlOvjYHZnliklbnAB1LTDpzie8NB3KIpc4ZobaBcuTK9ypX+kIGf/qdMqqYtTpkoPhkOmx27i
F4IWqN3/icDs2tcCYM43lVPz/75rIA5YUr1lOJd8cAOkLh3kvTg81mENTA6ElLUSMcgBskPAY7P3
KT+3dx1KS2WdARp8NF19JwwtQYEeO1NLYpgH9UNdeTmD67q5eJYjwrxF6jpI8LhfMmz77yJdR9Nb
q5OzcF9wJaSb/PIIUODz5Ohsxw+SfP3LMXMZDlVV3kkV3DqcIGfasILmCB4/GNJbO1/vOsJM6/1Y
A0M9fQPQqhp60QJlLXGuMhJwHaMb6WDXRqLjryJZZ2DrSQP3qfPI6IRClqJT0HHOMTsuRO1674RX
DGwQvgX05J8h7D9JR0mS7muetXBb6wkCtWOPXXOjMhpZrQQDhCUZH7yHmQoUzjXXhGQRHJ1bXHQI
wzRF8ChrrdxRP75lWvx923tiJkA2UKDWSB4uC3D88ENvVOwlpx4LguPsYhwRRX+ELY+q+wYt42xI
MkUKr3o32X86OOf4xbYC3vHW01FLs5i48XsKOUWMPduESNHtGM0atUZ0ROQFM3do/jyshMr14cdz
pYa3r+J9p4fY+iNzgJwWHRpc3CeCUH2Y3pcx7qJ3ZeZ0p/rgihmeRn5qCZijE4no+/QzU95FvBN3
NqnJQ90n0WI7s7glPUCpYhmHjMVL8j0s8pXKxRLInNU5vs7BDTzdbKvNhNuYOQD6oni6Qw93zkNA
ArEbtvQa2plHy1tzOkxV4wcXQNtXbIDQiIWtlK/TD+32AF8i0Bocs4vq6g4Lmg8yoqgh0qrTZl1f
cnadDHwV+AKEHsZeVDpPkI5r5BZn9/Ts0XuKw0sUUm5d/bX5/Vx0DQQBvs5zeIFmpUbCpmlEE7Dv
f227rALSxu2gjqfBlh+hvb6qWYjltbgUYpdJd6OZP0VfIkIF8TKLh2t9zweznDI3y2azhM+xOqEj
T52InV8Q+hZBJaKVwHrXeMaYUlyUHpr17Zv9IgE7xOWwmhOaguaiaNGQhp3Xzr/bWa/zcPl+qQ62
jPeVN/pMU5XZqgqEepcydw4rIbGV1IpVwDJtizCs2jw4qnsohU2PPrGUaA2yS9MYM3EE/6S/76oW
zCiRHoJdd0AqYJmrhj6FN7y/sA3ROLQoQ8gI8lM6V1MqlYKu/XL4pxEHhEANJBBvnwNldyobx8FJ
IdPWWeGp9bbFCJrkW3DCz6NWXEX4vzVfmr6J1AyVYgt6sktaA7Z8Aunlw7oQES8bvMFYKs5O3XhT
vtLN5r4G2Yv7kpvfnBi2a/9eJZQAzavp0kkwaJX4tCfp4ORHkkBeU0dd8FybW34lS+VcHrTvnFPa
Y9ZhviLTjRlTVErCGQL9bzhgcHdfP0M4+bnAEM3vemELIvV+bULiwdHvEkoZEOLfZs2pAHHBt7O3
p4vDfWB2D6nxNXnP2nPzAw+1/cTlDAuNkZL0N9Q6HOjS48sANJIgIacgGrqK27Q4r/nI7tZYceLz
8fY3oXg1CX1VIxB3nqVYCzQCRweOJWqaBUFFPcNod57CibccYXC8JRM0PvoCnophE3t34V8mOxsA
2N9ZSrhAmIxMosvNA7tS1kmSE6OuomsGOuOTHJx1sErhf5X7ZgfNAcVlYaOVNePxmbvCW9wgS3fD
3yt7MlJc4OBOMT4WCZbFY5bTzY6wc++tTA9OKoz8GhHLSvgNKv4rgNGh0l3X0utCmDOh1c1NpdUO
E8xWw26q4VWv1ke6dZIJOkH66rNFb3FKjZxiZvhUGsFsGhGPl14MGoA/oAmi5iB3FtyvwsDVQ9uo
oCmLzyUvaI8L2CQH62Pus8bJx6y686YnJwkao2/maakT+So2Pl8wjOOlX/x0K4SN5EdWKfFASN4l
BLOWwp4z49eZMsCTZWscbTs68jvBgLk+gSzvje8Fjx2JFNPjUhjNsV+MWzFIagxsZrj3IEsW+5/C
mQpOqs8/2mbBEkoL9eo0ydagsxtSxZvZNf7DUouMuWnH5fQMOldJB+WQ4H4zMQRObmW5xjiCj5PJ
nclqUgLqyOHd9nWNYU3jqzxhYOGvGOP4Q5nPKRHJ5LZnAt4vGKZ134YYeymCTqpMsBSAeVBSpIle
j46ePzy+sYw8fsowoECkOHJGlwj/D6iJJt5ZiuPgx85pjVPnfP/ulD/a9X3bxCJ18oN+DOBo1/M4
nr39sFwUmuY0x/ZcaBJkJvnaLDiwq9mnHlfbpEV6y/R+Oo9ObQ2Od4q+5lPvLY3RYpAdz853wop+
Xm+WZaPXFDucmaqshYGx6GxK2yiqRlXIFrWmhjzZ1VvzIxbI1xHcIQtyY82IDlkqcRZaebmuWxgq
nWdOzPP3pfh7cuWynj4KspLmYyKcaVJM/4PRakDd15WsReZ8JRLlqHtix3AxIYzLydt1msxYw9Gx
s5pAkMC+HtWfksqQzlG7OUy5LMBaqtNGB3JHOBSGDqatiDM0EqHJ38oX/XppNUIp/+ULmmUc/NSx
UC7Cgrebk7U+zL0+GuVsv/iw8kqpKS8AK3jfeNWczLh8YyL/R3PJ/lTV4BdqlXwEJGjQHW4mE0af
e7n6io8IZw0ul/ZhLVRMTD/opkvGHWjLQZsC/+lY+ycu+oPHRY6gTQ1YvFdzu7bS7qVXwYHmTWOU
12rVtZNbyG+p/RCvE0GrDXITZuA7ap8xPctHgfPPLd1El3Evf0KGtkFHbyARALEVrb4/q1gHWmCY
4FJ6E8N1HL+Dh+yU3CAEP29ElbNXCwt3MpP8YoZ8xE8AZCBQk7YbxL4lxnI8cfBFmbKBjWaSGG5n
JSMaFuT2u65n/a8Gb7cXNCTYHREefhmjByNX5rcuIauoIOIecwzGyV1F6n9vYbZoDyspJ0fuEgXG
n7q/nsSV7OszirJrt2B/X2wJ8FSm3tyA1s6qOSxghotAc1nHDX38sTH+9LzUeULjvP7Q6eBgFhSb
W3OWVEbwcWePK+5PIqAygFx3IKjrJWyfVTdXJEhF6Atdx9PF4buhHHJsEjUtOoC92lffOQSc7rt4
Pa5jPLQMk4JQIgJE8219TMrg9P3e8G7WSoNhO7LFmew8BwVU7Y1T3oytNqzE8HqIAORefXrIYq5E
thJuEcd/hoMMQekGrFuaT8oMCqYZeey6eCP2qelsSIAErcNAA3iwP/VO3Ifs7RwyrGdDo4J4QABt
pl7pXSNhBfNecPxka010qtS7eaGIE1hCvtnjPbCkGiBDyVBLWHeKvexrs/rHIWkDrcMlY1VF3URV
RapKlPBo6b2VXJziPoeBUngCXyp2CgS8WAreqB5G/J5YfcthYJGc3OAm4yKkhnpCmr5n0zBXu4nb
OiSv9+sKTkYW2GLQWe/InEtB5kZuSEifTprDcSCbu6+r4yk2foiTFu8YGCR1MqSLfwpb/6n2CSrx
qiHlOHIvcvNPaf4qdNkKqMIWTFae/59crhwPhTHMhF8b8raFHgxzsKr2Du1y5TBsvhO9It25MeDt
NqY9OdpFAlGs8NrqksCyYr4BzAYM7coHlV0Vd1AspkfCNYwnxPu/TYlm6xGPW8PoJYtutTGr9JFy
tRHPXEB/QE4dTXXb9i4AeYXlQ/J3Kb2WtOcY0rfjYOIh0HDkHjjdDQdinJY2j3g/hCowDBu3pL0E
0qHZNEnX9IIGocMBnEIV0cgI2o6OQEykatTCMlgPRVqluc4mckIEpQgZvuVi/xj2zbTNQpV9+S/i
cidxccNEJciwpP3yTE37Dne+zVClX4iibKuqHxiETMgii9Ic1WjUu4HSGcHCA3wLkxaI1o1idcJP
Arzi/rTdO5Dfr/iSocWeR0wor7j9J0114wV9POePkYGKEI7+CjfpiqAUGrtdzb6XK1EwxAIZDZoZ
solP5QhyxTFm1l4RgexXN8jOvW43sfw8B2SLH4fIh7+GjWV0yxzKY1zy67qqsTiUYwiarbh/iuSz
NB81c79N+5i1agJYzQWxWG6RjRiJ9tzkK3IrkQb0cqflXylobBBdt5QoMeERZIFyHBpD6zrETVPS
iMo3KBwKFyXF8WU9HOW4cD5Is3k8VIHvjLy+DU3Htj1LIyJ88MOdLj+I6IF8sd9d3JrigMg1UR44
mDqVnzcnQLPBRZo1QPI/+HeQOeUw0ZkibS2KDnOkLF6XkroECSvltZ1f+HCbiC7nHyMzhBQoIH9g
JJ1EEYyNrd9OW6g2/oOVhCkZtIBNoeyD+pP/ZrGLFotpatJLHTLQsZ66IgKhNKk4jx0cq3oZr1pG
UMR2JZNxi+3IzQIVuRmuVx8s4LGUOA/WwWZQhzvSYvkcAqe1788VUqm5IRw6w7h66utYj/VoPFnU
/kgzsY10zacN0GQUE8iPo440iWRE5Jm2xQ8aoxu6qBATSXUGhSuvQV0vXyy+4to25CxdRccCpHlr
TeJwntR+2vKfo7Uq1slk5hnAKCkLCeEnK2zxshM6ZL85B7fE3Cr4o9A2YN0NRFRljNgJ6naAQTCJ
aSHHyf0cWH/iy8L0WL/HdAgcpT1vXL4WVo4fTrO0W8rTCDNhmKwgsb9G2wADAxA96Il7O1+6c3+L
Ki/VWnm5G8hIh7eAJCftls6Hs4/c4pq+vosyR987qZd7Wvx8adzhThwf7X49dWv68+hYvF+T3k05
Cpc5EyP2ioQp6DachU+aRoYKQigsgguxQLWUklQCZm0BpS9icY2Zxy9FZxTw1im5OlmURbywA3O0
RvqTt8blOHuBMKSRuafI6atIb2aAyxECqO266z2qmuzvGLoMGj2Fhqg3FOKhjvwHVDfHovw/t5R5
hUQ09Yyt9DFCWRhJ6V46eZ9VUO/a1NcrPvVngZkzVca+ScjBiwaV8JJsiKFlXk0UYPNg1f3XeV/C
HfJgJi6pQFHsRBzYPJc1O8IXR5vGykbSwtstsbJdqR8fHMbaWLK1Di13KmBzORkfNlsiyYoxFXf4
XvmVgGcWxiTAvzUEgmkc4Z/BY5h6xj6EUFal14TJLn2FCljlG5BdDfiViRpQ2+i/vuL0JT899kvQ
pWgaty3E/HxcWNQNAdLm29Tb4eF0SuxdiX1a1e/ALsg+oG3uozfvoVAU9s4pcsuilK8paQAxZuGv
6Vb+5aeRvPSr+uHWuJDvnhlKd2YCQMrqIEvWAxzuf1XlMCTf/tVvEdRoJLp8W4Q/9P0TrwgcKHYk
zrVjRfZt+ZthnjJFGCbt3FH4vbCy2T/wPDzDJnS9sQoCEhACodSPQsesJ9KiQZfv9dxtO/+ZPxGO
jkIaAVUSIYXMo9e/bMMgpOUbboWWXTRAoFve3Ffw/qIvkPoF05Yqez7ziIR8XtX9PsTMcNQLJtoU
kp/kX7P636bgKKFfbGY2nN/wI+XThDeEAXXKmxhGzIcetM2BeDkcDWPJtgOmLPt2fXYUZG5PU4QM
wrVENq57Zl2sIc6AU+4l92T04HHR3bNdxBaZ2ne7xFxzVCHOQHX5f1gW+pRp9dF4bAHvfPSRsK1F
uwRSI3GdT/e5tTAWk63z0hhBXMd+hQ8rVP4D83ESN7x+uut8ijixEj02CCOWajsEBXgREvHmvAWP
aQDGyzOm+TqH4oxwLm3WByE5FiRZUEyJ7rBCQOBA6PU9OKzQ1/AXcLQMVn2PbV35yDXE2p/jAPix
xPnKy4FNAmNIp0dxPnZFg/vPVQL+PgvoeuR9/RBUkfDUMtWmeY18tkrbjEzIdaYR9d0rBUVST7NP
VG7iO1Z+wSc3L4UXY6DNURvK5b4KM7ghDhsErE3Nu0/Akmq6G9jo4EMUCavK7+osR0PyfBZIhZh3
NpLyjAwS0JHgrqFdPIi3WDRgR5LlVzkOcqdRT/UjgXHinUb+z47XLXIROeKTXNdCKAeeu9bYSPrL
LqoFMMxkt07GxU52747gZNFBpFWTLeVyrqqqMlkXWLt8qQAOPtVT2JGQLGWMUOl+E7ZXC33n8xv1
wWeqeIMGSYEftRCDfd5aP5hQfJo+jXCOQHH4chqK7/tlwRi3qFEUHzg2ZObbFjqabEqkU2z9rMLL
/SDIL37i7/IsTvWG0pz067OV7LkO7CwhNyjeJYOW8kqDuaxBGFUFKL9fCS4KSNzrJHNQYmeAQNwN
OI7fSDGxbkTDj29J3wt4sHwJLgEJaSOBMr7UxEsviTwNZjY5zp5p31Ol/yVSkdymkZPh8ywOCOua
YJpRiSiRCsJtphmItcTb8MYqkmdyXZlfmcQOXapjusK/WEKKzZLFhUX08MgM+y/u64mncyKI1oHz
20Ks8zDfTQkfbU8E+yt/BaCa5yWQ+0FvL6NjIUOXbEtIlti+ft80iVFKo2QPCipfzReuWxod/hJI
oqIfEHd6qmaOJrNCosZRId+k0ud0U28R0EHZa1clF3aWHdZXtZt4WfpZaiT99/KjGL2Kd0HyKe28
5lLhf2bf0uOWkb8QtPYyxVpfnDqLTIhAl/FE416FuDmJ6gL9grH81G9lL+hURo0LKb0z6f6Hi4lG
8GuBi9J3CH639cIUukXbtqneYURV+RDbU73ITLx23z0Jl5rfizGa/fKAigc5gf/Bk2y+mqie/DyN
bNBSIyhuQ3dNq5F56EU3DngqZE4RmzRYQkB3yNOAjBvxPlch3TWnjgio0jEtp6Q6jgwc8AvC/STT
uzYioK397bafR7JIVuN6PLc8YgkSvJM+pGbQU1tE+g9zUJ9lQS4NGZ5mzCCHH32Do9PXEEuD4GFK
GbcgRJCOTWVyg87ZbZ+Pfi/LrRl2NxLY8P6nXHZk+mbViYj3n2cbbC56ztf6jPu/jOjtCHvJ9zbQ
3ss2jEC4SN4YxL9OqsnjjgE4D8iKQ4jmTrMt10xF2/870cdD7hG0NqRAN0FTb4Y7emUDzfuiV7RL
lW7EHRGhCp/WNZUuGLbAUrSvCR4dfoV6vcYEsjV0L6mREGzaLuEErA12+48LrZ46EQtg9yN+/kXV
okFlShYR7pWwm2gh++V/mWOhQoIPrUHjQ2DTQejay+bZrtx0ZIBkc9/cRc3LuFhXT9TR7XnmNjyu
OPo5nRNDm/9Rnf1K5/IsPx8etS/yV1yD4Hqyk1JDGR8+IFlqVYZwHGTq8DJ1I/uzbmmAfyt6KMgB
IR0PQgKQaLSSyXa032/u+fZ16K2GapOarteHWnuKNapqTXr8ZR97pRDolMXiOJeD0hq5FsBMuEDC
8pfngXE32+F2k6WF101+44P3Tb07fm1B8us8hZF3T/y7stwJRKrszG69iAUcPC9ub6RGcQVEkBOt
FFBxXmVjIaR8U3Y8MrW63BFw1jXHvLqPlQl64o5nWSLzPh3WlCPM7sw187hpAlJXDigqTk04MkL/
dulj9tBnIKShpN95Y0hdqyYHxFeh9FwTGFWBxESt5BKO0CGgxI7sdQkdb2t9UBwbe29KY57/Uarg
oGe6pltCSJSJgWqgP37O4a8TL+C+wfsmF83LtwXPZRHCNqdNz8jzgezb9u/Goep75STyCTETHIuk
7F8l0hNy/q6YwPSqyqWnon79WR+0ZkU8w9TwUZmu2iYY3Ju4JHMfX/s4pelt/HrKcxHEFLVNOt8c
X/bkZs2Ac3jvrGX8RFgIXPBQMpXwdKg1m7xroqkpnzP9aG08MeMXk5TvHw1100tH5IoP0oHYoSH8
J2RwyUm5q+zenzPMBL+KHUvLVYrVci4dKVBbqDzOltlKDuO73mJChk/06WdDdwQNA/qyNZzhjNPd
2L12grACc//H7zYlXy7PWrM/m4i30IrcaUVOIxaEg02bVOmydTxEBEPPMHwC1sxy2wjzKqXugBK5
wr4ub/8LY5KbTTcCqmdb9jmL4WNwAStnuGC58CPLdtZYT41nfnl9kqdfQs9TkPw5Yj11uxQow9ZF
gl1NxVz/IDcEUMxXpxNm9rjIHXHwg/4Q6oxuLgbkjZFGUJfpsIapRmYZxgTua2/CRfviU64dQpL2
kgsEHGL8FptSmNrCSAk7ThclDwyg+dWZFxx9ODDlecEVWdZDPSFMN7Hb1o9Kn0R0LVryVl1IJoJp
sCFGYYTWqE3pF5xgPqVuiXiJRGc8IDjfT2rIv1qFGXBdBzX4n49OdvRYeu2rluHgl+4A/WOi3m4D
TOuaZ/6QAPidztlxjEeVm9FE3Y/jadL8F1sMR/QF3CdyT4CFiafcqZ7Ds30oi9gFwI2nju77yFXw
PvKWgNsFQgqScqv8mSvAfhh2H35k0/0LkNiNFcMuZJXHE1csplPO1y6SNAaWvFZwCpah5M1ETWj+
nBWYAtOfO18oFJkyiqmMweQDvHtFWxiyfVn6dnbG/vFKkjv/FAfSUSlhBSxrk6xNfQ4uDLOl0hh+
VRtgvXp9c1s5LfFftNRIQHU30R/OxrM8O6siMjm0LNr/HxpfR55O10LC0HsTWPOc71DqcEf9uuQE
W4/bTDBQbY75uepk16XMTrzCGMKVZKEygquyU3vpphryTda9ZQUwYoxd8Qg9Ux8caBBEhiiVWYyn
geaPlSbbVpynvx6ETN0Ky+ivBgrk6SectBy+CkeoBT4sftvDKKmGdBcZ1mAt2jUF2wtaUB0wKyl9
yD3p8Og+lzWiqXceNbv5DUH01Cjucd9pCGmuwH8Fn7kaXMFJ72tNFHKqvgf7/gtz7OAi1NWOn2L9
8vd76UoeKdMEgEv9XVN4g3VuE+jBfMf7SnBbeYbivVOMz4iCYoU/zKTLeoTIQLwOHcrkjEVSv5HK
fZdUCgXIre21UnWvQxQn47qojOiCHTY9xGOZEXaroj/aW99HNKrTjsDVh3mBlIaF9nxqMxFWriOn
+fdVj3teEqU9s2em4rIG5fLhKI4rkkp6XjXsveyKJq/DORhyZsE3JrYFcxG4DQ8yRJ278sofzaF6
ZIwotkPHPeEelpSiBVrGwGlMe1lG5P5qol/SMdoLYiZRGLjBOHKuo//DVN/04OBiAELYSr30sl5P
j2kWe5eDRb9A3yMhDUN0POJMw82gG6/KqF4YJ4mJbpmVb6Vo1kboyEKsyt1dL0U1Skr2vOt3WrWd
3hdw6SpRPYaMA49n+nsXoCU8dfXlWIttvJuGhQB5Qb30jXmZGEYH02hwFFXSeDOtllDQoTg0uj92
vG/t0mkvzkVwCjHKh5QMJwZPQe5UuS28UkbCIzxUaZ0iywFZTrQBOyA/e4jECFGM5MKlzosAC6Ac
lBCaHMq9ZidgF0bST7eyrG99oyZ+s1JBJaNHuTB1P4hDej1pUEetvj9OQ8S/8JJhSTMXZy++sYLP
Y/Ri4vHBrBKDtvTBYPqPjakYgpCu/cHg9zyS3QELxNlCAu1UfgnkzkgP0p5nbGHBbRiZcn+wAkiL
Nufi0iC1QJH1g72hJaCbG/oALUIHv8MoywmZj867GYfK6iJ0rwiTIc69GJYOgIxafsPOITaIiZGz
blpKGZj745WK7BqsoWp1NH3ClKn9mePpsHpZVUe560NwSRf5UwVDFMgAUXK55aZuuF/KR0hMQ69y
S0WfmJXyZY0QphUy1dPiS4GCQD9TTGD2eei17cj5dgd7nm3A+4KWk+FbRyQQuoUUboQFEN4VVdxx
XsYHloIt1W/8GTFdcvpx9wZ4cG3Fl0aXr9Tuqyyvybn+tG6qaU4GLnMCr9vdrws2B4gp1fkmpXLc
lmnluQ8dV2oWw2KvEuqKj4ZE5YMnp+4Uk1pNJ8TO9XU5fSdwZFzSpebCcXHsb/Ht5x+nanIYpu6g
L9YSZa42DDQFxDJHydicMe+Bwis2ihr3lPR1PhnTR/V7rCdqyGMN0x4/1LUNcLlg8YNhSdvgl/qZ
dSMptx/r00IbpWigbky6TrZ0+1QL4nal0TVZIMb9fjYETPK4LNVS50FcpV8hdj0FY+oHhVr2CMLM
+VbZh/1tSVQ+ahzfj42hPIL/jcr/JkCRWbtsURUvC0szqyzBWCsm1TbaF4iN86+BnRwD3zs48/kH
OLCusvBo7Ylcl7Rmdh9HgsBrev9jUof+GCBESnfwpCCIDBYgL/SSWaKsp2kQaX2YLnqIPpIf+mVD
2adX06YCEaldM03qbZ1ubwoBV4YsWkkv6efkYIMleg6R58HNJjvB8xU4TVjF4NQcxEUdG9cLVrjh
W+zIgUdXszkrdziKiL865AR7P/qMAFUlrARkK0qRerEQiXvuCoO/1C3/JqN0dL9g6Nc/sMn8iV+F
ldYXseSetNNuv81IO/JXto1OaKJrv+fMvcFzPZypeTAPo2BxPXV68LReIOr9kaIbkCNIfJUpe9xg
lX3HiLekZv4P5tMUG4m3k0HGbulHjrQyP/rwAx1cmiE40ispMVG9Ol1/hufgaogiASFbTXVlLJyI
qThpS8rX/a7hufEPGJMq95F3c76vY6tC/kEdFhdW5cNPV0q2/GB3NUk2XezxXA7XnAF6ChSVv1/j
QU49GdoPfeNXGFPWPDvNgmxUBd9yrhDLLUJc382YAvsNYIMzIgySHlnrL+Je5JPsOPr6uNeijsC6
SQWMEdHSU6uXl2jEDchdQ4feRPuu0+4G8vCjhzKWK8WgZ5XzMurykrxYqdme9jGJVyd/PopI3EE6
RSntTsVMbHuQIFgPRGGf7prcN5aZRiQqMU9531F3q6GP59SWeXrpzulyJZ7EMTowL6nQ5uSW/D6e
0HqnntHrbxfNvZErZXNlEGp50V+4e/le3KhK8KBeQfR6jKsu5khXQYbUI1HQ4LwN9Qz45ebjqcBd
8/ImfDL5OcPY7g+KOam5NjtghM9iT0H4prxrSy64t+tmIxCHtoTat+EePdHZidc63cHFXwYCp+9+
EXDT5N4bS+dBjjdFKCJB3aNUGhqaaOeCsbBJNKTSXF75XZEZij6yGuYx+FLxWsOswdUxG8MlEYU+
RdVv6Jzx+bnEKA/tmmieYxxDbRU892/T77EU1Zk98EDYmU9TQ/1DqCQL7QZ66jzs43Hxs+1iUkMh
0Cl+jY82RxkcXQQLqODpKNbod0rRxPWRChG2x5JbWbuJ4Ca6CQuLVLtfD7tkzf+/24xnnDu2fEyw
Ier7kripZji4EhuZy5ou3SdZcQ/TCWOIgRO8rD+USsyoux6kp/IbMvJygKFbin9ddwESEhrJON1s
QshAw9oz1Q8ErWbDyxAgIKRBtqDsU4l5l0TbBIClYJjkSwJvM5tt9JkXTdP4zCdh5THRIEFFpgIq
kmPbPGTvznIw7RkIV9MS45ExReGkSZ8i2ByNfkJOTIDAR05XZpQ9Tc+fj+sILMQbh190+A4TP4vS
HbWUeZM+wRc99VJ93FHAiD2YysK+cLmtqJFYGdI0uepIo01leors4QbhEchzU8BAbTHD4osWS8db
CmDzbOLhJ2jezUu00lkHRz7eEYbHajZxBbC3FFFHFtTGL2m9s6nG7gPvuA2itH7M3wwH1DkUkUAE
dxw/5ptgmXRts/S3zdcLMSwqgpZYo9rULalqAcuH8h/1S61Us1XS5LHXOOAY+u/MYOMyzS4Ky9BZ
AVAvyu1aQ0JN4MYzthyXYzb+8j6cU64OWD5VaWpoSwtBsey9VMZCH1iZbeBnkUIbHJ9PY9yIkAYP
MTaeWdfCsLJS5DEKhifzQxMbcVItL6+rbB+FKB7ARmgnFXDn5xhuufEcKD8IiWworkuBfibBOvdp
Tztm2FFOfj8DFxviJopLsNBhK64IoMGqvp+DugPGp4H3Ip0XeabCJ0pjfwHF6Dg/+lkRi4tnQTst
ZtZV/MaUkaoEa+w4SlwFbe5SGoULeZMOzAQ5hXNmF9miDvATLcn/piS+/Pyc7sxHUHOiiCKSXinP
Yeq+nr3FZ843q9mHK10QRcwxxWyF0VAd8/8ICYh+/XEWgcHd9XWc4zZcWagkMqmCXNGwGgnzfkLk
8nUSOxD5Mjupvm6ih4Gmp7S6b8Or4ov8O0civZ34x7Y0wKwhPVQXdk9tQgrJ4sCMBPz3FKSSlMVf
3zEh1Fe6N8ztVJwW14wbxopVe/5iW7ob65hwV9tSCNJXjgI4rFpY+PoQ96hWvc7cD6exFpsccV5L
uTkqaBzgnWqe5UNBEw2zOF6pxh+BJkhnERqCJdGrCG5Ap51wSJK1RsvZukJf3Kfvbjpv6tJ6ykt8
oPQpTe2v4GiOgU84eXRIGCSJF6t+7V6zgbgeRYMejybOtnGg41rNm0OASpxFtQNUTphr9KZQwSv+
vco927TaWq+RwYrCE9tzSjBU4yo4etol/GKrepVw17iXqaxo5c8wkEY/3VH3FodlEphXKM8vY80s
ifal0EGPTGKGRHUWnxE8gUrdzQA5vAj6+emviZZ4As7xGHDU/LSTv0uSjvnPRDg9V9968Iad6zv3
un0A2wKRbAY1TbKGsy1nKxDHAjmdRK/YmrFEnlhMmzYASBE/Zb/WpNeshExtPYKDHaQeKifVG5hu
wwKrx0VitVXyZI7TPuf8YR/RiXh3uvqRHKVj0xR13EjFrFSa94up8iLfkIHCIBQSS7qdWxC4l7P3
Vocq+87XiDIYyAHkUcA3pIi9n1fgBhuXOR2MJ5+7qIm7UwdRD8+R2HUgn0OXMEm78I39HEc5trOk
9+IXZR7J6I5TEyVDaMFxYmcnEW3Wte3w+cSAJnZXFP5XmRakRquZR/kPTqbB+kQhkel2Iw7QGz7x
DG7X1NCmNgaMiHV6VQbA3mOKH6a/lN5D4FVdkiHUU2wkLNLlYMEvEpRpWhGwjbSyxi21xa5FjJ0t
9cyDmVDBxuWqAnB/TJbEF94KNzquAxfqIDKA9qtozEEXiKBOoii9Bm9S6KsAp6wFYBG479AHMkju
OdO9vgUyZg/kyuoypaNVLBCsmk/PZ0S7phtb9MqvksrtXEXr5TEtI34rfWwXbHJl7SFPTuvqiiqK
DauA2XxaKqOHMhvlWmS/+51zXyVYP2/wbHW0YK35XfEvz+gLJoyiAaQDXEYkayNuVBuyW4uNEyNH
RyHDDCdBrHpcs0ivaPh5q1xnaC+gsl6CW9a2h5y+d07uuCvSHG3jf+KEo3Vj7hpAaFzYcI6go7/j
n6bs1Q956/AcfKl+0KGwAR06rEErjU0wNAorhLdDlHWPDmjpuLfKvcWEJjYkbbTZvdPzYneKggfa
ne2/HMXx1OGpaLsZFaRL1cryefGYM+hfH6oJOPEWfp10Rni7zSGJCga5gSrPvWxxmclJJgGgWxDt
nOLvA1/2AV7PBay/MGmsuBq2/KHO8wLDDRT8twPaBCVnEdN6pu13jFhtWxf13Ed+2JbfotRotfg5
MCrUrmB6eN1Zq3+/aQoGT2DptiT1Umh/yGzWqWiAQwghuDivpFpsOBcL5APTb2RGGdXwm1sXXEug
3gWd8DcHMDSMtMmBuPJudYRX6pT16X5/XlCFaCqPFV7wKIAfRUW3QQNFXzLkOWn0lO+6A0/LZ5TL
9ikUW6W3Q85G9S2HIK8B6rCGAQCii+kOyDz1nVYMNAP3HyMm5QVz9hAd83IWPB+LhKhnm+IMPN1e
WJA18FZvhg9TbyulH0f+z7y/RiYPYxT+1X6nOtIvoEbXXH0j8d3XfBrUS6oFObO9LQMu5OekWDQJ
VD944Vx7MAiAqGWo3SBgjnCI9QJe2/Z2bKjz1bgJlhis8bL3HnTbX8gyB26Q+5xyPBnl9QLKWBYd
8LK8iln3XviPxs4vK8m6MkAhX9srAFWq1usaWzHoU+3VabgzEiFp3/QJqo3CkRNHSZfdBd8RwF3F
GD8hoCxYkO36ZKp1ksx7Ze6y/QzeKve0z24P2xJWyPTuX7Rfcw5nDgec4Bt3EMBR2Nn7GT1XjELX
o+8+gQlBS5781yyyWu5UkqKvxxbuXiIoh7be6tIGV1ktQ7iXrkJMCyb8R25E6p46ITsvrv/EkEVs
eqL2CuufuExCCNyykdfBQOdEkb3ZXM1Pfy4Govf/+mQfERkPGSfctpYxQK9Miu5uS+jveAi1ttdK
xRz6JEZbugLgoJvoXGc/0lr/994Tf5WYf6YaOEZbU0fUbHxUpqmJUME1iKSctAz9GxBkNZRaaqra
1T2sh5g7LzACL3IhXBl0wiNaUQa4DeD9AOPrB1xAmP4ji6SnnLoCobWuwPqKIBqM6/EDhKQk3jFR
7VCiKBQro5OUEkhCApnblNm8MXss8+ldyoSZOCUsba5RhQe/lSGteekxq5jiR5FlcDHyGL/jPYi9
SQaYmcYwv/VwbSaRQSc2DyQgOu/Rw2R4Qr9xWuJ+HKHxmhlkKkQj1iJofoQfMV8tgghKSBKpDxXf
fSIcKwduo6zP+Ohn7mPM9WUpTp+ACXxhkkcykm0uPguYqu6hFZTsTGEIG2lRP3H7o1ujlDLOj4r3
WnNX2GWkpmhGSBeHqcM3rn0FmXT8CQ9ndAfdolHe5nbl0inXByb0Mf+iTf9MVCqPl+Bh9fxqk+7u
Tcfdy6Qcb8Nuv3reFjCmdUAlHUq55V8cbx/0/LE43zdrZlIeyOji7UT3rsbOXO6PzsILnLVTLI3U
JqJ3K1lanho2BI9REJpNDAOUxgJL7FtmtmrPkE7I+Pl0RIEB32FPXf/76lSEclhis1hFhUZNktJs
0zDdnfqxBUr4MQPZeyE4+7RX1ddgoAXwBzRcfaKghVaYMRZJoYAk7UAT/7tfgLwceImMvS3L6Op4
IWRrXGR2WubaEYg1JzKUJTJa62O1geyFDT7MJNV+rDKdAi5J2nJWXDSFEGaLo/T8Wb/Sc/fxbNeb
Wc4vB2u8Otg3S+fSIOU0pwOWYqKvFDvjPV/TOSY3t/k7PmAMa4cxVnO/wkC9IYNxYdUr7U0A5GOP
DvQmLeSUwFi6++WCnncMCdbOWWGkbhpxzQU8oDrkSJMjpVAIrfRSbTqksi9OwWxgF3AXABMmB9wZ
88jlN9WaSQeu238plDlTzLz3lDkLzdAdgx+dBhU+r+dmuKJ6PVusqIa6FzHB8f9e+zfASb5JrYZ0
DW1xGAjszyTIiWuY7sOpz2WqRL5VMoOfvuy+wSL84PFg63P1fa2eD+FTolSjHyLkhaZjwyKPcTmR
3NT0vBZM02X2/LTdK9Ev6U7Ny6wy7qM3RDlaUk8u31SM1rVml4rxke668QPu2cYr4bszUBpYmTp3
tXK+BIYGoYOWEF4nSo0aRWHqmLXW8TPxfI07Md1baDxAsa/2dZhkpdWb9kancQGn6pMCg1CyMPpe
hs8nB68w2reuYotEMRZAyGfIdZlAJM7sRoDuplGtUMR9ANN0VanRRSmzG7dkA750C0gtLafNIV71
WyhF1mq204L68kxBLSZIC2c1cSJAIPuZlPsZtaFmD9veZjsGkQwWst1EA/Rc1VHE4HeRc9TGZ4VN
sxwQJ/A59ub228vu+bGuwQNSlfZYnhWfaG9+Ah8wuzOOHFmO8f/qkwBaCmf7NtztXQKi7hzWdQ5e
groWSGQfvc1yjDsB9QkfvhwEIGWqPsCNEtDwXVUBt4RU1V8wU6kD7L85eefAJYhAPRnmKgYHYvRZ
bXkpuR6YgdClTkaEpdgPBQd0x6j/BINdlpSCB+Zctit1O2UbH7W/tTKAduwl7lwWJGxupII1qJvN
Thbtj28azjcQ2wQeGHLefbalJjkk1wWER0Z5ZOmiIcOPfe0ocsEOjjHpBC3K1rWNwifuueIvxKaX
BtNMbtTyayPXzEdB4oDCgUv0mlQGp3GGhQH5DYinWbWKrC3XGUv/A0fkYZbBDzYIchmSMIfPLEyR
1wItof8fMUXnGtE9kLWv9aZV486blF1JW/pYb79urEwZKQenqpvvA+w6rf9TlzeSSwK7MIaMrVrI
Q/H6jdUtyIp5np7p14x3qRpnUAw8duQVqcMB8itdzMjDcklssQZgD7Ty61ddCZHu/sydoaOfCz4o
B7X4oYLLjXBIuG1F+opjmZfkjtXeoyh6e8BfCPkctqkTbVI/akAiOmwDrC4FlzZrn0gbcP8Vj4mp
0BnyCa76xGobq0pjx7ipus2XmgM+jI2h0vElQoAay9Pw/EQk1ntb9BWOwR+4PdrkXpQT7XuvUQvi
uCcxb1cGVQN92ByDD+f6n7TEtK27TFb+xhCYkGTOCCB6L+DB/FMr/qOOAf3CaWs9o0EweXVhK+zS
/+lqurFAMtkXXUEkVkH+Me/mSOmIH7R79bGIU2QE+FzRDKTIibLeQrM4myKmE5VHbWQXA2HqIdur
XnvXf2lB4C6us6YjFV4rHoJegu5oOYa5/sHooQkJ1Ndnu6mEieYpSrNbSjUF8Wn8SdOKOMHKYxr6
+IOlAeT/qQGD8GtBn3rr8IzVeI7rDapNPbH7sPhdHOfqz6K2TjoopQztaf27ihWG2bDZWbNn2gJ0
25m36BDKTKSPgMgxXxfIxZ5Fc5JNjc+x6k8+cB3oIy5NT8Pq99TjC34WRW5QsagFHsRZQeL8qEf2
g19TOIA3BCjHdixw+gq/iZe3vxQhb0f2qwERce2wTKsZVWbg417J4rKfRze4jVx9jzagPn+j/CnY
yQZVKn/djxI5hV9h+UHDrzrxFp7Y+4O2hW+jSvhsuw6EhO18Q5De3Z6HIY9NiEesC7EZK6NVj9QG
HtiKVeW7J3N7Ekr43H6HyUdrl6iRxH8YfmUI3xcpC+7E99cfFoo8eJqLhkeCc4/FELOSRKxPqEdX
ZGYRuwWrPNoGcYj+VkaKm9+MxRxXhkeBW/z6Fuhx2BAxEWV8NCrazHJCv3m+Zl8aZ93KyZkGbwKE
3MR1Iba+lqirxXpjp0MRCCGJeTE9toe61RbBV0p3aWBrfphKN4NVFcBheqYu+Sp39PuxnRDB8AST
fCfo9BJUejZGiTfKoz5mrVi98bhpl6yHFahpQITNEwF6KyCBlI/bSfYvxME3/hpwI4+1kypfmqi/
epgw2YWhRsMMRihKE0Z5Hkr/cW/OcOdAuka3KDTgALJxI3HTLGBLK26A+uoSKuG2EGsnJfy3wHjv
jIOoxFmNDpothQiREbdMBe9SCiBHqGuzcUlF4U+9dDa64AXrgRBmUksOPN3qwuF2ksFhTNQzOKFB
B7zs0qu3+0vkak+RzAd8QWMJMeVTEXhep2KdEQwhbihIr6PbcTSYV/3zxcPLKuFUVpexH0buDBgd
Gv6Ct9yANxkH/YDRMivAd7wxXtul60ytCPdIzbZra3rRa41xotCpFJsW2bsKONgIIvwyJLhrXE8c
fU40A2T/Z3FZjakuATyu0LZvjK2xlMeXLpB7LMaOY6TrGv6el3MzA3IdcFqLrmqOyScLi5XWVXc4
OjjJ1BblLY1DcdpK/TJQSYaiv62PukAfg3MyFhbXMncQ/p+8ttv+3YYSq107shi3q3svtqnpvVg/
WnvK3nJ7YFAZp3NOdKHw40vklNokR1b2LGOyeljv9cfLtg6UJfK55mgcQLROAAotuPsf9tMWfP3G
m20n9jaIJhpk6U2E9tYsVLzTGKh9PpCHE9i0yZ1vvR8HWLmyQ0F9GQCnfwoc4M8hLbEbQH3moKCa
+2XGel0/0JeB5KTja++la8OHQdYzp9x3dRXj3HXDP8qMdu2LHs4b/6PSoG7w1EkdpdJzXtRIKN6k
aUW1oC7+N00aql5ziCZS7cv7t/SWLU23T2yxSfrN4c62nM5X62QVNCwhY96X39IzxFijRjKy7Q50
JOzPfSbuMdXHLq3dD0qtIMNd7HQTzYMKS7dhhc9gs3RBEfXjPT8VhWILr61T3ECrbFPXv4fiFXIj
6wMRDZJRZ/ksLA/inZQYnkiFZKZ8QTfZO8fcScWEmlAwplnNe2q01w2Xkwcn91NHaGQaIiE5dKKm
oYiD0Faloq1KqRabFtk1JqI1+PNco3J+NBQOxXlh5bQFtMe9MLsoW2++3URfm/aR927OkviktMjL
8oWZviLYEDyb7cQC4C0Ui+QaakRZV0i+tmAGcDwF6cw44QKC6Z4S3ZDSRdKtqTsmbXby6qFlnQZW
rh1Ox4feagENWO6Pxkh6P8umE2dOHBrccVoDfCl4+6SVPXmIhR6/KJ9+icd1Mc4NCBP87oagfRwc
QGcUgjCQc/OGxzpLEc4BYT4oBXwMJIx40cQ5D3iu4L3Z5XcSrYkIZgMojmaxVl3nZVP1Uj+8u1pa
ajL4rlx6fL7aCvmDQMPpPeqhE24UemYswEnJi43DL0BCWLabjFO+cKsVjU8O/mpEW5UTn+Bqma7v
Bf6akkCZmFxcF6qYta+g/rnh256EBCqDBg+l1TrLrABcqpzi6ronlJiDcEmR5Ko6mV5kNpMtJ+HA
esdTIz/MiJgiVvrnN/dLC/0GNovvVWd9/Wd3Jbpkox6OXN0fo5M2cTzBczJrnexLZSi4QekLFG0s
//FrQXAn6XXMLuZoC9057rZsXnh43XPhcdWZQ0NWLPM2KTcTq4YHiB1VHt/yYPyJ0pxuDBWSfYYB
5QKt4Y6tPqylrYqnzXzKpa97SgvWI+VmJuqJICzHRWpZihVTzWaaKOaBrnkP60k6mOsAcypxaTkV
gspOS5pr+5jJikrU4cD72z+7pASmm7FwgWhXrrWl+fLJCkGuuaXHyddvspsUFgQmW6L4Nde2FlZJ
D7K0uEAfZ/1CvZbCKn8N0OjQhb5u0oRuKwDiJ9wkANSTzIY4ZxdcnNxz3TesBUovFyc/45cxRqeR
oGyrYUqH0MGpHVJNvsyXTSTX7+RImaXUVpi8ZZQMpu1KhTZfy65pBYJittT9Nlw8D7XJBVmD45C2
QzTIRP2XDAuhAFz7I3Ms3RMrx56Afhehx6hPEudU1Mfkaq6cnOmUdBV3lZne+chFrd4d5UnQ11LF
Qv8M5iKvXI0v2Lb49+Y7q2Ma0IaKWQmFYhsnJGuMjAvBciFd7k0YxBCg9RxGdHmHNq4VjjoPih2t
8qdOE193zqkEpOcGDrewzMB1lOig0jpp4uCi71FRFUciFndYOeIGa0MDhxv/E/3zvCNMOlX1/2Cf
xgKFwCDXU8+Fm+2Az+oB8u6UFAGC93DlMMqhOKwNpqyq9WOX77lJx0/KcZNWKHS3toIOllANQUnN
HFwQ7xD9Hg7myHOhylZRdt5Ud1fQMHKSrPNgyw1QhvtWugRxGGpsZcF90t3qV4ZE+kVZnu7mTLxV
MSZshHMgwAdcK444cBMfsuPR5lmnptPsIPhtR86JHVigKAjoKzNpa7jdbe0fFkOUCn4lZHpxdSGD
1Q1ao8HoC1DBNXxVeJHvetfq2Q52UOG4h2APpIaORuGFdwCv1MaHYngbxMw8xITkcGea1VseJy5P
F/smaxJ+Lvhfi+vq/wz3xRfXNY/vKBofTN1IrxsjFQrpn3j6hmxBQYfguMsKs0aACMso2ogmQS9y
VfJwSKgs1NbXpQltymoMH9SSj/djHa5yOU2gILZ3z3NnDm3lWY2TnmEl225gV/nsCohkgp9qiRaC
xhjlMPrVSq8wsd2PPpcUgJfcKYWRvxQ94bWJb4CLzCx5RM7GaK8hARcEcy7Tmv2hZSbriJT3akfL
1sVZSmwHw0h7awCgR6Tts+35NQ3duJ+SgBKO4iYgWwdluO7onfPN+KcBgse+V0UMqU5KuNMpnr31
hQMuFnx1nl9fpzM+5YHvDPidqjOJOha5so6DQ3cXFG7gJRl9UDw6QvmyS3mSmoW5BKRmTj883vrs
OAuQDTKG8XLHNssYJhbzcHu2kWZOVvIp/MXY4td5PewGU+iQUVk3tQ6f/KKjluKnFWadY6DGvrqZ
AsLYxUM09nItI8xt94Kg497mmntk2j05RPNvhA2UygwDfSoz1OaUTMwCSk+jjnbDvf+t45Ea+r3R
zE2OXTG5fUcpWrtAb59BdO+CQ97NpN363LpzgWBVOTUNqZkfz9D9GBY2uLzeuZtUuYGrI4RBwoVp
B/6mfoUfVqluYdqTOt/vj1VKd8XTe1fAPBs36NrcoczZFaBf+Y2nWSJdIXmfeIPv3cpbG9I9XL85
NnEZVmix2C640LX3mQPyibpZj6CNWtLFitmAZ5/YZoHEbRe3329DSlvhhZ9j0YUQDTu8hR40NYq7
+ndKIuXA66cNW6Qt8Sm11nThKlYm+EtYu84PVkVl5L53Dllh9LTYRvEJ5z62+enLPTnrNENrL78Z
gbc7YivqwLOsELRd5R3QazSwC3rKGXgqqRdk9ru1SSD2ek5bE7wF3ctMiB88Bo78MGw9kd65aRke
Q2WvXCeBUiYlLxVSHAk75pj+m7SULfn1lM1wn1hb/PcopsxwG+SncIGKtYawxPMDnsiZIIBook6G
7TsaARB2vTz5uYYz4JVE1en3pZOS+edB+dT/NbP2VvKsLARHZcNUguRfowaBsLHnf0T9M05ewkc+
DdJI1hk1c6+CjN2pLiGqDAxA+s+/oXjDC1LOMCZt+RZ91LQOLKk0mpycGFtNDxz4NW/wQIvOh+f0
vL3lK0bZALOc/DlUhaa9Sc+ouEi42yRP4fn8gO5eOubaZW4hZAty6l6vOTZtdGTgUwT9E+UZZ4OD
zq1dCBUAd5D9j8LVCQsqXilFAfLv4WtBdKiWZWvAuswk/JjVWU9tUMemSyjez03/SGpwlEbCLcVj
9pkCcMo+zlCRJB/kMsWbNn65Qyk4LEE/i8A24i5O+i7b7DGtmFLIb5i/q6RJFEKAn7Sf7BMIT9IK
T5jn/hmG0eEp66YsZqFccnrRxPZtpiw6sIYGVys7ajn4EcZm9Paf3HadFBDy6J0WRrrrcWSmoI0E
2F765oPvM4Y2jGnBzshSWSY9z7HBZyuCdzoZKemAhzjVp6BaF2yq32xXa9jocpsEZ76rfut8RFwL
IrRW7PiRCTApAbxUlHF6VjWtbF/YiRh7j4JPAm++Yrxz5T5uf5qLzU3Zai/owOwBa+d32drxNr/t
Gi9LTLEjW84RMU8gEK81KTSn69AUSskdICFw/eUZOT5V6Aj3kKBUCbF22NSHzR2rW1jvBYNMTzwe
JTZsOT9N3TB0tyFbKPjfkBPVsM6rN4OVi6yQMz5VWPuDttwK+ro6OBjc+YvwnUKKooOtPmbG6/mD
lOWxXJ2lPXC4Wdr3+cYYNB6KVXex1xNuZDBZd4uXTjqtGpR3aCviZryeKlDi5jmFm5t8G45PoQox
0mohLDdiO5mDWgwFneALr+cgEdjNHDLhCRtSpCGBebLd7PETmVn+TZ5fjZ0P4XQ+XGZN/ADlJERn
L6KlRUr9HwREaa2cCcxsuyuA5waH7EGryEfXgO3kSkUtBNMSHrtE1Ics+4Ei5nfG7LgAeCoVmik0
DaUVgKgzyWljXL5HRZJb1iXI5Ct4s4CKILRCuO++pVSOfyHT1h/bX1/VWicMA38afH+9DF/C1qNu
qfqnbHnzRPrbURk/9kOcuDPQZCce3oz4yiq/2NTmAB4GUyNMW4lrRojILx0fe0Pykf9Yp2PoTUUP
JE2XIRu0ST4qoMVQzJEBcGZJQbrQwQ+g64eRQUKjSSDS1jnd1CyxSBL2UtNdhThtyAGZmuZCmpSa
DorNUc4FTaZv7YBHj+l8goJhUqIkk6TIZVTJkiFA86xdm3DmO3Si/mTllSAMjgOC6++2hEvhH6Bp
V1XSm4hKlhxwjTrgOBTK4wGQ3FHAg8oKsd6oLsA5KCBZeOel7oP4+lThx5XajqHGupeNMDdw22rR
b7BJkoXdeRaATZe7dRj+KsIt+ATUL+IQ088uZwmooigpFs8kP/hzpuyjOLoW9dOkzDZsWTMzZVhS
5jMt1gT1JvobAiqmnQtamqdLeh8G4dJDlZf7aYbbejOEuOIpRTnyQXhlwNNIEKL9PpHZk7p+fkpo
57MNZ3xhkw09bsSFuyPigCprTrlbP7nzqHHZLE5NmGdFJozH/dtMXYdn3vxoiPP0REJsssho70mk
9r6f3GvvfFTr/KmiZdPRXhIvuH+6juAuR06WWDQwBHtGD+gwMXDHocQFsXU5BtD6N/pXrcjaq3cs
AZsG7WMHfXTdGs1Zd+foFWM+DPWAi9s02gd1pdt22NiSjlayZBvviMxQgjhzPtBRi485y4Jjps/6
+D/dvlnenJ6VVoiWKNrxe4jf2BO6RUcF4vP0sKJRDLLsstqL1k78Um1MVSCaK0QBhtDdWrfXpmDY
gCh41vsIS2+FzXNRZ0lfdkx0/MDz476q3WPXWlCwOWb+xbQl0xg8bGyhiaERt8Ud1/CPYKwcCqYY
vg94mrKc2+g2QoiC8JAU9c1p6xM/tK7UDceWXS886u1/+jnF1y6Zk8Z3nxoVUqlFwWhxfKT78t0X
sdUs3gocSj0m5C7bXCT+vDxVjsEe/YxprJ//0TS/e7WS+gzQOhsjI9eAnApmCKPTUkf29awFxsOM
SGNfeVpCPVLR8tbx5ek3aBqaghnH+7hUSVXHR5MWhW5hOTFQv6ZFjn2Mu9kwnYR4VEIzGhQ7ztjm
f0xfomlVfjZ/mv7/yTDLFUOTX3JOTEplzJDegzOXrMZ48AmE0MoLrBxkTDEFGiGp6JcyAI+1QVxL
xbueqyddFm+x03/UD44ZlHPAH2ldCM2rsKRTSPyD0aZRMuE2uNyDbjgPzj/oZODchszvCJXW0jvw
Hs7TviOl4nhSWtqNcYRCXXsg8d4sJ58ByKG+HJwRZQVp1B5nYVIu/RiJiG9QS9e3Gb6fUWrUKTSu
H2+Vt88q+8mRZjfZudcpLu5iOhCBJ+O/TMS53Y7Fc/0Wyej2Mgs3f5riYc6VFhDH4qO8+lB+XCF9
Bx/wm7m2vG2U5A+L+VumqiWeoMSHwaQFxoYaFlMk2ESnlz64SOyhZI90VD+ndZl2vbuUi8MbKT9r
ASOC+PNHeLynfhDTk8DSuq1ipYangbct8sBTL9TWHWmVvVt7iyQyP0hKQ/fFuYf6IVEQlIRWE0g4
pvYgYq7+1G4dA9ITETU1Yi4cJR8zsFXGJpmiU7PpUlg+7jrwL0diMUAN94X2znHMPiE5T9M7nqDC
pGiytNHoCBmAFM1dQaH3MbPepZQWcGM71Xa3pUTEgVLY/fu8GZCScnaOVuz1gA0GHbIq7s44b78C
G0hHWV4QG01v1UBZzlTi+ZcBo2EZAKsHIJY6DZDuqPKEuxoLRed+0/vexX0reF/hnWXST1vD0ZEh
dvx84biZqEuiuPrUw9IdOpT/u/mqih22B2n8G3T3KtphPoJ+E/oVmCIosTouLKL2Q3DQF7aM6Xjj
B1t08IIvL4h5+DoNzbjBztc3mBSHow1Th16TM8FYjbgtGpqDLEJcnbB0R40k5P8hrI7G1Rjuy4Kf
hAz+G6JKLjBmq6EYMgcYj73AcPtbiJGfTbPBsfP/O5WFgnodPc+5NzJtON4idhPpAWnn1kaTfkrx
eDIFNutMWo1LOGBt0ORCkLS2OR4e1xEvDTIBxwrATxR1dQ3t19tIRYV/sz8uEDZhr66LPPPdApyb
q9+XiKOqoSR1qCA5DhJA3tG00gZE6T1EA5IUnGVcjX/trW9Z7GxpJXlGzZe+sXxEuybbkDnrvEdH
Uq1/Cu6fjnlJUkai6ochvNS/K+g2yL9Jddt7b7xyr0h56I18vowOtFFbAs4LV2dViRq8bfwIJE4k
HBD+oDSVm+ct4qNRpS1ZsgBFNiik4arqESPUTa9qaGvt63Xw2vfzoi6gqk8bfhUzNTiQmSjW5FsR
wdGKK6p0CuQ+D3SOc26798XtxOg9pLrVLME1Sk+Thrf0DSQFHJTOmGBtBACB+C7OUpRTUootyz2h
gnm6lsXimrDcEv2+MNns42QYOyQHxBr/BzAQE6FwWVGPVuo7aww6Y4tvnk4mmccAe0CaEvKCIqC/
c/LzZlijHdtg+ygrh26S+Bk87t/8a0AveA+j0Ziuj3tW3LWgn6QjFEXzXNeYkLuiWabAKT+K+zfu
UVbn/k/PM4d/srHCzEnEeZFPD1Qcutt2PoPG4Ehwa5eb5P4Tk/+X7UqoDqudWuArHhDMHSJyuG4t
aDjvVFvyEP247MPGwl6eLN7GpLTfb+CvXOgn+OUPEOIqPBipINyS2dDjKz1fJESeCXCLUaLmPpMf
gJbmGPB2ZsqSS39EWduLQFD61naZYU1N4P9WDLqFTR9l1X76FlBgwJgXhi9ShJ6J/PsBuFTKPUnN
onGtOtcR9+AhPvi4M566U1jWGwoylA8O4z3CY1akJir8bvx5XgstnJvvuwjpvp9RaUY5sUREbsjq
3o8Jc6/fd6PsDAS0FLYk9L2yud8Si9JG7GqZfP4XKVj76UD0p5/lcocoSbHK2F4iDWX+kVBymW/E
/T1r6ROOztQyrkYrfWfNeDVRGbPocWZYxhlCUmukuqdBoRFkpwfsgL4e2C+1y0GHigWPqn9QSLU1
YPGDQVH9iqr1GE63ZVwATA/msA2oO4KUyJOpRVveL2eY2CIs5lbGioVJ3jpyKG2I2slOM/Oq9gUM
jLfPOmPTHPh7W/wleVrSWn5A7OmgFHD5vV0/J4RAyOriCBBoTBrn4pgB3RjuCr6IUpua3YokNbhn
Tlen8Zbu4jdkHSChr165oJY2FI3cPiuRORoCocuAkNMFyHz9gGA2UDqVSF16wSK4BHzJDPm2wFG7
FU2MhYlH9oIhaAnKTMB42mLMVc5uec8cw1Cn9FXWRLFP3LMlHoPLM+nENeKUf61UQF9vMV3+nWRp
wlX5Jad3FUvqwEFcDrIC1RUoj1WWWFE/j5aUdREzkVhVxX6zZ2wHASqRnyQ/qIMM/1Z7VE6FL+04
oemWg/+YkIe3DoagZ/471Vi0unoK75ZYCINYgA5zNrpqlncRUCe2/vFmEnd2a0lbcytnfca63+L2
HOoqhK7Jwt/lv8LPEuKo81CZ13mXkDsKQa74Fym9uebhtiDJt6HIF2g2AjToPgK97V+N4fN9fj3k
O3DVeXKnd5jnC4KOenO2mfwYu1BWMQhWrsngCnhnt9CVmptJiyaD3v1v5eKOPFIU0G8RTt/50u7v
lIv5oEWerDK8ERNE/ebfDZCzy3QBMiliM/jttmrt/z6DaMwB5/hUU3lZuBYSefdK2i/a9H0ZnXO9
0KReYoOMYcahTKWV7G20sI/kff9y+HpqrHVrn1jat0n3l35KZGwW9CevlboJjpOERo/oXUa/McIq
t0xnI97NzAQAA2E4j6ORq7FDZJgoTYjpnNFuQv5txuNw3fDQlBJH/wE2Q1EPSJ+9wpxQ9lEX3YXi
JGf0iuAYKdLCJ10lh1YicZv10LB/HEBqA8jKyYFKs7JT+ZI2F6KFiyIP+2jC38Uv1P2i40buxjdH
lcIv8jwLW0bcp3fBEihaSy/qM4w8UPypQ+epLEUX4BGQsBrphPA60qd4XRX9UAVereIKplNEZt4s
63p/hGGY/Wypiqqhjl9iweNYjMtOkiE9AC1b5AhWp1BKPD6oUhV2w1CwSYoBP6Ox8jXQX/1sNuvt
FrbSuaIzKzLAXNcv1AIZkHdyFntYi7VlWrEHEJLu3BHkiRawxwSBIPhw73qyiNf9RbFcq6F7ZZVO
rCRbNTyzuTXKlh/mRf6OAuAmJqhD8mAGhHzHgpTJKqcndlC+8Bfy/PZ7MxQQxrhl0X/RmVv+uJlt
p+G/JWa0FQqgy1j0IwYrSeYevF9hZGxTVO556PwA1qwI/KIuNDtSqfTgMVEyOh9pj35kC76bUgVm
TddQLgRpTej+EUc54X3end7z6Y+uVpJQacF/0ZGCSQIDi5xreIa2NHJF1QC6v1AyQoe1mIfcPV6g
HBjEIRPScWiYKR/TRzCvL0xhY8juEFbuTF6GJZltSw4uVyugvMcePvqh8ajxnKyaWe2qNrNfsftg
zh6ZHHq1p2rZXxDJrJak59/X87nGh/+MOsVossAPD7V1icHa7yP3QRbIv5YkZaOa4z+bZPGvZFdE
H05RX+LO53dP3WsWBH5xNsv3u1G1C/pgSbTDCyOWPr6sYEv/FGRtyZ2DWWnKm96GG6iGO8L6kGjL
vn+DmfdFzQivvlXCC58z6lO39ZgbUGdElEiR1IVGMuCLxxYoAQ+2fDOX/tayJxNY8PRH8XWZdQKT
oUCgfO0JGMAsjAbhjrCBm0BqthKFsLWYaXczJzgy188Tx/YaX06GnJVGnVJIEZGq3DfyDx6tZdlF
hqxTj8buu4l+sKXBGCD1/3CZewx4cvprYb71v9DwU0ewH1IcI5jdf2Rk+tVOv0MX0CsFnQS6s/3u
jdnuIrPqrOztSxUhvNwCSEOA/dfmyyzYhz8U3peh/hAI+U3xD/4oGI0a0A936FH+iMry9XbCaEaj
iiLFeqgPp5eZFZQK7AVBEkpIU34ee/PSUJ5YcXIRojHzGZoOBk53dO1G+Ir9ieoSBm0Fch2ioHwr
aJM3GzzNjJk4d8b78qQ6EXFAZnUeLQiwU9Qm0BU2hB2d7b1MrguNpIu5Zi1/ij2Z+YlJg4W0IuDj
qPfEMedhnKP1RPlrZ8RPCjexMQz9IqJ2rqXmfJU+r2XE5zmHoghLBIvnfgNsWb7Eoh4Nq/s3/Ucc
pjpyVCRzfaRJij1jqeUdgirug6+eqYsXAjLcvM+eSgiQXAUEXAK+ZgAoV18u3bQYHyiZg/o3cib2
74KsQoIGEH60w8nllK97qIqqRQaxWwz+rsIK1srR9S9wmy8ogBTnM+Oh+ym4KagEyay6sOIvaMZ8
oQ/pl9gR9I253zU/GyzNvSQN4QmSdqIsoi4D6yCC9xcAl/vy16ck48s81QD20F693qWBaa4qTpZP
y3vN86ZjPlByHrDNt2rre5U4V6ajmAe95z7kazgTxyIjnBcXUu0+t2ao/6tmKFSCFDAIDIQ1NNV2
JXSoyLas4NGmYQXhSbq/OFt+Li05ggPkT748Wm9urW32Y125pIbhLYu3DsWN4resYgoxwP9on0sf
DZHL4lU4n3H+xru2KaLOTFTRmzhE4/Xj/hJ8kSCKjARHbne72AC5Yqdbbzl6urpN/fh7Masg0+2e
D682g642DisIlhBnAGey9dIjtOzXpXSjm+gFVgunG7Ogs5oIY4B5qpWY/qQI86Ebj36rPlj3iEmz
75N2YlC7yKhi8X8dd+6OSPX0ZeR8YlEtwF5umcLbIy4/25Y1yxrfFsAQaxS+XzWnhosIVF1Prgy6
rfeN31I4HTAuwo3mDk5O+uevv+Zuyz4w/UPgsvwNHPQbYo5Bx7ypq+Q4ZwnkLpsueijFpiEqzbx6
4YY6wAjvjuTc9+28G3vZhtmzKdJTGmYbiIDpuPtdzesi6/EeQrXJCIbEHX2yKsNyZX3rF5jM/8fH
C8FGb+EQoFio5akrt7W8/+qV4AqcQRRmUn8UNj1eoZgxSFScYUWyeenX90DzHNJkm+S5uaUtaxAD
UZ116M7ZKO/uvw5M1pO1Oaq+kPdptypNimMqPPlTpNjUvygl61d4MeEuk0JgSlzXQLu8pUvTKZSl
aXv++VCuxL53xcuvHTDFQSU+q6qSJOpZiN7XgGPaHZJn5B6tjT3d9f5ju8ypRHfaWM0l+nPSliLP
bCdysuDSdO27PCDyuN/W07BsACBoui0YpwCaYjaYbl4TBO8oCmmj6yX7QoJypLnPKf2FoIUn0VYL
BqOy4ZWF6N8aR4PFIp/Nv8QAdtGZQW8KefabyEmU6bjIGPbL4idDI6Xxskz9UPM+TvKVe1ZQERr2
Q5ZHPYyqeIGt2Jp8ypZIiBKLQfuBT5KHaNf/zPvC7mJ/lTKduBi6evXOBpgdj0CIXN2mqgA64uNG
qDdaGYoaaANKTXMsaT456wrgMMDs9dB3WD1VmzcTb+mFP06XH1mnzotzErhv1HyQw43ddMwShq9i
m8C4z7BtaxLD94KV3wtLUP/31hqa5cQb2ZKGc5gjUKvz8VJ5MPicw05dG5VrsTCK5BBCLqNFDYnH
ILljmd/5wN6gMlXJ9vPnj8kGys4qgchmVSH7QFX2a+a0FjYYdW/ZAPft7fnMgccq/En/u3fzl84s
5k1l86HfqCOU2E3p0GHp8sZQWyAZ7vamnen/ugM15nFrdQinDZ87shL0jVuRLtsksJ6fIDR9uvmt
YyvQCL0T4oGV/vXYOVd9qESS9A9tXtbH7HKpxLDG1m2gx5GOAOKCuLOAvx024FWedJ+oHlGIfAWe
l7DjvoA5+YkhvcLWWRYbxg0LqZ9zsupvit3YZdf4M4KEZrTXmz5EekmTk8NT9UJ6+b+sx/Zv29AK
wiSxOXJRIDqVbGqInGEqEIdfxbwHz/sXNHeeGynRYMMqmuoLhpI9egZLa5Il2Y7bpvYEOSdfFLAr
wL43EcLXgePRfrr/h3LDr27oliWV2jyW5Lmmu0J4QdcwnhTya+wmlY6ckhATK3ILzosvB7S5zEKf
5cnSiD7vhc9cSiqWbu5aZ1eS9f6E65pWe0RDN4lcnXD6gLyzJwuX1FtC2uGYyXrVbB2T1PX3KE6V
HSHelb8PuwBJc2l53me4jNnLq/4w2WKWnYHB+h91x1w92fORwJSrNsMWu+7bjk8wPZCzGbqw8CUc
ggC8FGGOHmL9swKXDUDBnQmihMZOf6/CPixz2uAZM/06OcgyuYCSU1z6ne2o7rzgUucZm03zdOq1
II4iHeQe7Ch07+bM5NQg3RqmxvWOeg2uUmMSifs/dyb02nxe1O8eUOgHjLKdDj+gP97mWX+GXaqX
L2xR+498DZ+NIM3Jk03vuL45SOGBFpsbXK2zDKdAsq/K6RBDFm28o3xcvqDOWr8gKGGIpRb6T/tP
7+LMAkKpvXnt/QTgbovHH+68n+Qa32AUbTcqdZUd2KqCz3oUaXj4DyD3FzeAb6fJSmHyW6eX3v+U
twLP8iTxfnhioWGDvERZa9oVY458D9b2cBB76chTjFvqP40CnT1DoIgOHt/qy5Fd+T9SkOP3wQSI
qjSMJOLl96K+q3l/vKLD2dd6G9BUhQhelJ9z9HM3Zw4anpqz/6v3PYGSuUesLQmdpcPDCIASP/Sw
Ym2XnoMeHBgQs6h9cfJ92bL2QnTVCfHwsfEiq4dK+QrDAQuEoVfymPh0Mneo/JvucHpn/ZA/dKhE
Mmi3oldSxQbhPPMLOvLTpWQkjyRkGswDcrtPiN/FZg8JSSl0/7NA6SEJzdFoXNPQ3Kuv7RKBw7mh
v/6d8a9WfcskX3uyCQ5DWe+nGd0uKsk6D/IkJGwLjwvO+uwoAYjKpj5HIUp0AQba71ffBIlF5eoH
vQahUlfceunttZ7/L5CgntuI/Z+KDgry+3FuCgJu61skqRlifu1ee+w4wsqRRLdD0V2A0OFErkAS
uI02pdHJalV4fLA33omG/5PGMesiTsv4S9GNKxPUaiJlCfjWpirhHqrix8p0ugnMmZ6azgwCOF1a
oRS/B8WSC2OZvyRxxI2xkcRiT3umlBl6+5CZroeNeSPJIsv1uB/LXbA9/07sshwA+YEb3rl1iETZ
PS4Y+3XVwmvAmiV6jbwPp6qT4mop8EbPhdCYa/enzFwAGHNcwjiaouEQhqqxcg9ff2SxVkJ9jCBO
U/aAuN4C5yjoJY/iG4mKi6LXC2e0xkNOFUTxnA03ROv9iYMAd3J2wDJUnT590AySG2QozSkmDbQ9
q5eVsbYpabiVRO12YFMecFpZ0mHMusMntmn5n1jTEN91TFlprHXmZ4AzZvLcPqzfgB7AK3IS3Apz
gjqb7ZhJYRP/Fk1DdxU6CkgL8GVyJnaabfxMvD8BnNnSVsmiqcX/vpH9ruxwvLJhZ7QHdHAsGN1d
Hbbg6u9k/4P/VJ006imcctLCl03TwUc11zJ/MkDOYWwzeIX1R6MNVhZ486KDWMf8Plw7N/OdH3MB
ANQHDgx5E0LosWYeMe2PcGDS+FYpS90OuR0jFcx8uEO1uXZMLJ35IR3ERK266IqUlglYGtQlARjM
PaWntKcl0qds7xHhapfCUth47RTRYq8pTuiIZ4G0Q+0AVTqZp3wn1xuMvf3hlGrW2W/rzhdyUjdY
YoXtH0IRzi4Y4yYtA55AkaC999jhSO3z3UfPK7mACfUETwuYmcgtJQXV+jE4mDGdE9TYd/vVUXVs
v9G+6EcWxWXFPhEfJthdDBkyT9DjfjcaHJjxtOcUkEMLWUTL7xR+M9GsUj0Jh+pNIM5Q8Zzs7r+X
r81rcuvOH6MT3bAveUs06v3PL/QM8lTaZZEAHUELlLCXCOR5BXIO1yzAYVENQLuW0zYa+bp9FuWX
hmpdhj2jQLV5s88eam0wQcis1BkEeFCzeH2CKzkLOo7trraEW2RVVptpgKqn98NyC8JNHcaCtIth
d0R2ej+GF3KdRbXeC+oEwCn7XS1S1Q/ePW4xL7/kPX28SMf+hssHGNM2Ur3gvYE6uPzb1bcjYnEx
Qj6anMJlnFxQUKWYnRkBVeFueB+kfmHZzCFsoLdKp3DKRETCxTN0cVq+iNGOoamUG6x9oyX+SwZH
s/DJcrHY7QOnTCsD3Vny4wwprahH/6sVYrxtYLCr+7fDEcA3X6N/WEPfyU5ENFLKnb2y+3y2rPwP
DkPxMkZbBkFu77U0Zsz8hn1paM+f9nmMET215zWNwEEE+7/lrA8/lcLA0D+uS87nJuhhbLLhPpxB
H7rCMxld4QtlouVm7nJY2n4jDMWVV2SGSkFVkbsbbe7Aa92hE1cMCtPYm+j2j40jeCJ1liEhW7Wm
usNcpglDQrwx4w83QoaZvM1xtiudeG6NY3scbX6Aryjm5fvQS2m7AgjewAVBubDYDAwGvjusT+OH
2rH6npZhLHwyAwronKG5Z3pF75slWs5YG9T+75abeNQzQRDt2KVrYANOhB6Z1xyDIVv/mjjm2DDQ
mK68DS5u1MRK96if4ZraJVjOMX4rPRPR0280nQmG43ITFVGFTEJaDsAGeE61xnzMiN4dsmLhffyu
VNrG4cfagKo+ILgheMktGbHcj0swtHn1MBeAYiNJ0Bc0p9+EnUELQ+mnYEIXRDl7P4oSmFW0s7Dr
Fdxujw4E7VOYlnRul42RfmtBiEWqN9fT4mkmHtDsk/yW+LEpWrIYvi8XhwW3eXRzQmRlOHdA8jd6
Yr+BlhW7gBywk0fYlt1joQU3xQuTQDq1Pq/ReavW8+dRqJSytbiDHMQVbuSwYcCvL/pSfm6h71hy
Xc/QufAnudpeVZ6jlX5Yud0SlXtTd6f3/pqltoLB6WF6dlYorJtNdy7DVN3bUfOJEzYKPsa9Nz3z
GpNV4vT7PlEqO2hFg4xU4vauUId9gMGzv0VH4Vdy8XjexZwlbU5MuiA4PwJKbykk8gyT5gg3He7E
y6p0qwc9CPqVLdPjIqXmd8Q7nxoPTP/s7dvTHAKR/jJRhRsyzyyAKHhwZhgO/CiDUID+B2uU1UoR
vU7ecg7r32gyOmta2QFqJJ4n3HkErjZhnnbI94iE4DU9UfwSTAYaljW+aBEoPVCXV4277oXUqsly
XxQfN4qErnFy0K4BbCt92x4O1joqQ8N6dn5lZuSvueZ7iUTqskb7zhxhqva8+j+fiUExgBiYQ0ua
95jXWXtOxi0JK4bS1aoJBteH8AYQ0h9qvX0BfLDNJvm8QcUwSrQqy8vDgkUzF37afvZvn6v/13bB
E/sJSlKQ4znuk+Mv9ZK8KrIOvlqXAD2WffwDaPrTv/K3uGhVYSdENSZ0traPRn/R2fiVyQwMetvR
WSZxTC+KjqDxj2XS0tAo9O4gg5sgMaNx8beMs0v33S0cFh6O0TzApWe0p03VbK9b1OM25tdCrU5K
jsmEbLfrE2x2MAaNx8a3ORzEoymhCTJWPEZfXplRNpylqV+HiqmfP3uKO/h+AmSdlAO+5Adc9rLc
dbeKbbUbrisdcOWv6dCZh+4Yf6fyyqqts+OykOKGTVSPhubgfJPDDq924kt8JFQYvsWHEP0jaU6X
D+uNAy2SF85Ollw3yAPAVKEgHf3irTv3GQOk0UpFTIyDmfRCxORD95TooYcXzoVvZIDYpUyzJSsV
XpCw/7oUPLf1+k8b0zgFxNRWOEhSVGxMFMxY2/9sx0CBRbkf6ELQpBQtUn2NLfc/7esyL/niokBe
SWtFnfRoZJnq46ciz5oNHowgexwecgef51NeeDeQ3aTCfYcurUQckJAmcWJ4zD7nNoqITDlPDqRc
7LruI0gi15zxDCldRHGZKefIaD4psHWn0vS8ouwkbJEpNdaiobeJNkx+tMaNIFQRVtCp4E/eqcKJ
hrndeMb/z0sXEmDc+rXXPkBwmal/a/8FeXIEgAn8kbz6rs/AEuUadtRg0UnibcQ/bTv3ocge65k4
PIFsZhDwNgF/PpMJX6qQc8CFsM6RDoZvHks1avzyZsynmJoeU/MUcFWLdyXDiv1CIOXx9k8ASBtw
HkqRBcDYw+VWU4wrqfUO1KNTgglqUYiXV5opRssS+Z6qc/ApdDuRODEVjtEpdGmW/42hkWYqLDSG
3++il6qBXAXpX6SAJ93u0FQ11ivUAe+3NK3STCCEa7HmHaCJWTXLb9MbyAqsjHJg3+J8LU5xqxVb
DGo1W/n0fBeXXsk9Qt6+u9LUJgGYxG3KRHx0hEhk7vyeSp7nXRISmPUVY/9PPRV6g1Pp0/BlFU6Y
cL/xu0fvlJTCXCtEaf0k1frwYfVHFVWtW9wCtWIY+uhOoM0AEkOSGiA7VINdc2sAC74PXWpVyIow
VZde/pXqZfcSg6lbKxyHQ0NI3frA4iNChzc4R025GgM+NkPcd99EZCkbN5heNnrsaUjYu1i0f2eD
ziKf5xV7Q9aAMHhvaKFrDqpbDSkoam0CdI7CVcowzMAt5IaoVSBo1ozmhNzsvIc2LDY3+BvYguWc
FZmzXZMpk5R5WAgi0ADJhmWhMue0UbMZyyjshGn3xvq0OkxynvraCA5kueB+uZomRkrtL2dcQvpB
EIoy6E3si0l2BREFsr7uAq87m34XtZaIlFSlok/CoB3ELzUGjxchk7Hf/sx6gAZxeARkC/0/VboF
cwm4XqgW0vGnuiCD0S6JjY76CDQNSBIu/6CSISY8lUz91PGIHcgf08yaosHqgPPxoGvBAG71Sw0j
PEv5/B/HDctnieU6YS64T3pZrSHDb5XApx9P2NIT4AwNCKRTmhQPG9vCoKw6I7tGFhLxPLzIbJ7w
LlPOtCv7mgA5D9uB7uLNEKYg7Jzy6TU88n34C1UwK7joVnPSl6pQLMZm+etBYvyFMbRGSpQBGjhg
qYcdB5OfEW3uq3OOUSapFT72W/q5T3Mlc/DHB5P3iF7GlSgtf1IvcmMTMSRa+sUY8iTKvKjzpaV9
dfRi6s1J8kCRyGB7UBbGbnJngsabGQR8NqWDIr3k9aRnT7FXBvkSlxE5Xt/J/c/ShFQmPqanqdr5
pqRnIvIcqsBPoYOm3BUQHHXE2BLRxiW6Bdj4ZIc4DyGykX/3S5vvmTNkXA3HHonHaZNGVe3tp3Ar
JQCCpt6OD5UD9QwwBpvGMZNAJMWlnZpr7SmFk14Q9ju00WG45rAj81ue4iif8U2fVUH/SoH+LC/q
CbLT8qInNIcysJmjHcPQMWI75apLyLFJZmkwfze5ouFcRNBzVPDhR+u0/w+FxRhHsHD4Gs2HGOTz
XvcIOj2k3na/tl6DHMFxCEP9BQHgTY+/i2kqfKldqymajOxD+uLmUzWAW1ZjaZNAqN5KPCtD5m4R
Nb5pPAt+Cn+p9eZIE71111y4X6LHHUUADzokl+fdbNtGDjOwA2H6k/Lu1DnWf0B/m3Ez7j5h3Rs4
QB2ywkeHWyHTGiLpVf7QoyksYoqF+8dvTuEN6S1qivA6wpnwjSlYeyic8IoVcBSXnoL7TmL34H58
FlgbmTCOGHJZzP9Z0j++XIsWRJCa2enAqHOFOCL9iByz98WlgVBOa4Uw+jwLL+o4tVPSCTRO/n34
A92cJ0merlfGz2ca8NlHhTIu8JWTpOflBHLSKLP3egtIAGSWwIy/7P4S3rY4rC5ULZgOhxsxKETq
RfkLeOJcITScFMVRTf+6SSSJFd9L7P9h3rnfH9OB/5FuwvjQZIWjIU7yi3KVAlV0ESO8TS6U37Cc
dNDI4TJHE45dwQ6zD/HqYu3X3d76+p9F1ogKNpoFt1bbyf5KwhdY046L68tPr6Yd8H9/i0P1y+H3
23jXD96b0PuPGpcCiFjTqybrgXG27YRN/P7mKDYi/bm2OTY7JljeoqPg0QekrhrpYx7oWWoP73pU
UpxPPU1C18s1+jJWk70QWjf6RFh8yhwli3uA2O15FEQJOehNjCsqn6O/xvSDmeUidls80IpLe7W1
XSVaxQbYfYkUwdNJjHi0fooqSMyey5MUFDd5oXSofx/d4JOIBsY7o/wiNA7MtVP6r4Bya5UY8b0u
obE3HhHDdc6iJbrl8I6GlLSS/kJt1jHsmaKhol3Jo8nrb45TgplWSX38jtt2mtH86Ye+jfGiIRUY
1LbpSkmdCTOvv2eDx623N7/1btmb9jFQy5IcPG7+yEyKq853KEd2sLa10xcPlBa59glG52/iztc+
wrXaw63j+v7pztHYB+3MQK35NMUkwEwDeevPfsvnQ1w3SARwWhzKNS6Ws54Q4OChT1qF6fCIVjnu
beO4pjoBV3M2mwKSB6q62h/ratfnF/F2BbjnDwSnG0qN/OH9D1f3sreXQ1wv06Iz/eEzR+44zNxV
IK7PDcGsILmHAGDSaGqgG61kDOa+s2dPXDULg8TptNltIVk6hLKaF8GmKzmRyZgs/+77EU6De+S9
uJE8ejE67CgCYBaXGNUIGVIpXD7k5zAZ/1+z78caf72oVG/91OvEJOmWDcTG/5y0fSq4Rcf1pXJw
BlFLCQ04vuFEvp7dEW6EQccEEsRP7lHSiWBdLGvInljY/gaAB3Hctongdkh0bcbE3yxMW0Mb147d
QP8xYDZQONo0Q/zOS/wLF1R5pWWGlLRioK+mgduSZtO5ieM4VIGCAs6fuDu1YIjkFhypwdlJnO6v
Gn2jgc010G/ts+WpYpG8JCc04cy5sgkgXqskA2HbrfjH1t8oheng1E/NCPlUelN3K9Wg44Kauz8D
X90c0/ZxRKXxDTrrHzTqSAAPT7bVox2CryytvuIagYZucKTzvytHO0x/stpZxSlazpvov9SxPmA2
2pWD9L35tXcrZAk6RY+x+Q3VEwT9WrI5gT7zGrDxjvE5ur7QdUUhckPqmU6ElTDIKoylxPgHq6RI
Bvj6JNii1PNXMuA4VF9l1Tlzxrw1uK+MZgt0AX61rXjsyj0m9bCIiGEzRhcTEBJY5cDd5Li7eZO1
hhoMwoE3mdReyJ/BDr45yWaFnSLsAjIcKMpimigsVWr3XmLNCNCMmJAFAe1IlZewcB9woXn9P61B
wNHnSYH8XUUU7cPj/9vGaqlhaPtenRf2bvjSlnA31U2W6gwboSCPE7E+CgIkGkW/mMLWlRbSKc9a
Aa8plcn0HSlieZx4m6cGLWv1HKxPFS1xzhq5g7oWLcjZsFDFjdfbC1PsdxWAJq7xBJOKEDXl2MLP
Wgcqc60SzUtH+ErLFK1Yqfnpw0u1+wWy5eawWsbrn+UmxosZt6UxMFW5u3VYFZXPhjsAHeLF7HPQ
HyAOYSjxYzciRZ7/sIFcCvsfa/OLwtaSEFIB4xrwgrXKEC/y7IMiy43rE4WDOjYSA653BaXRa3gg
nHI5zgCtxi/bA5LsV5KwV4t7aa1pJUDBXTWQQISIMT+spE5m1rei7dfHWYXVKJUr5eOOceEzuKRw
OK6i/xgC7/lpPCZ850QSCHwoykkq2roKO4d5gc8maaUAWipl3PA6MQ3oWq3DTOfjgmrFf8nc47OZ
Ji9JpNuanS8kZTRrB7bIgSsL+U27tA5HCPuJ6qHo3IGCCnHC1dslC9yQAlK2aGLAlBTEuHi7xUo9
naB+K/Chl6t5YMeIdGCGQGiBeQ4tJU9+B2fRkGN/Sbj3/S9cyRLK4emdbCT8dQDKMYGhQ4WoU2XL
vsHf8wmhE7YEG7ZkvgBKjTMHQ1gvs2X4Q+Z+3ri+qz5MKHKAeXfTKOIVDxWhNE8DssCDH1WTJY6s
nDH06nBCR9da4LMZ43bkmWIOQhjcY5kPBFt/semXU81qTB4vs2B9Ul7VLOtK5HkbFL9/c+0M0uvS
n80UmQIqtcgNrxoZppbgDo3rtDdip/Db2o3Lq9ZDZAeEN7Pc+Wi5VsLJZ5KkxWr2tsE8UxEfNSBQ
SrTTWs+8vP8+6Z4ZtPHkeJt/m/AdXQKdDg9PT0NLO6SpFM4v7hF/CG/yhc07Dudt8d6JFBzSiHKi
DY1JDh6VFyQLInQI7sohKMGi1pwkzr8AMaIDoF+tu/a+7u+TUp+S+yRgKsvoIEN0nyokvGz87Jk5
ct9bknWG3Djelc6zCHQLGP7XZDAmIUG2USZbqZlDLg63bKc4WksyVhQyOF1nkwg6ajkRFhE0NX5x
UlYj3CZgbarnaMlWYM+f3CHY9JKaIstpoHpVouLWg7Qrs9ystMwVOZc1VgDtMQhi2ptqDZj9mZ5C
fGKtkh0keF5pGLfu4+byNfN1i5cu20quoTWQampngMSUnib1eqHP5HWFIw1GyBJ+OHL2PmzI2lDh
WOChKXUY7/81DWiqxCv+fR2xV66TRskrKWeFp/RUtaSLqpAImrxmu1Cpkm92OoVYHKQmn+Q6UrnR
taQRQFvUh15W2dbrM91Zk6aqIVejK3LZTHJBsTjWUtmPF9wvScl7gYTXuMeVt9Kb/S5WPb7KKyRd
dyIFpf1G3OZMsb4pbdSXeeBljiBXvpKCtwQC1NL/Iiock3yqHsw9u4J5ysF5C7Gn+6FUAwCKj8zP
QDaYUxI0YVRqpJW2lqsQ+6Kd7S+6qQKIJLtptUWcaHoOlzQoC/BwDmISMztbaQ6xKUD+OX+ZOEtM
M+9pnsBtgNpnBafCVTd5BJyMGj0CvJOpBAkGa0oazfRib1GQ1o8+Vol4LFt5qa75FVzvFdN7mr/A
om8x49+8d5++8L9xfic/fAKszVbKRVFB2iYD0lKHacmSypi4M8SmkqOLqSKtTYA9tgGLJkqIUxXk
MTzNFjQCNHUqjxJo7DeJx9yl0ZtgGzoKXozbgqjzo6nevvoxtHMecR6htTQADIvFGqeE3D5W0yuw
e2SrO6D8otGjRPwh4iraZi7E9OIDa4aMEXHJ/fAhCYZSandVauhfV1OvtJUwz1xaSBfbzX1kR0Fw
usMkX70R8c+GEwj0DecW6WAZ7oY4t/Iub/wl4B2d28v20P3qro0s4YW1BeLl7StO7itxL42LEqq7
zPbjzdQAi+XtwqAS/yLfuDyblDAGb4qasrIU5yyYRXrum4Bg0gfXhLuV8mJg4xld+EcfBOAShx1Z
1NKZtY7MOpPB/GD1ZL4QfwOZERP6tqM+nXuazsD0N1kr/29kEGjfDdF1rvtdBi1aJCcKle16uiJ2
L9CVRElyr4GB70ciy3sfOeaHQCQCujzjSb9IksqpUdfBrgHfU0EbL8YH9My7l9nvb8CdMC2FS5cl
3jrhCyK2ZM7n04CSclbJypRzqBufW0ftNt3AzYGaF4y4GGDAyDV7/2DSu+fibNW36VIa2VtYFJwJ
61omygUs4JV/kkzEM4IZli2r6zAHG3U/+sM6TyEibmMe2Luu+3l7O4ETrYEWs4pF5DDlk1y1HChC
8wM5ITACVhDejX2GGdGs89rX0um72dW9lwE6vjPyvMj6BJZqGbRDcyhFIpSkZkrTW4mP2qMeuDYf
/AUPNbJBd74A4AXBzkW0mGnMkxsK0cqTkzK5oT6JvcGtwMgmFd92CQjPAx1uPANMu8/oRYYtDKFr
7BDFzTmXv5XUEa4yIPaJdh6y/ou6/1daHOZX6JRArNRLDYdAaVP6vX71C8XdK+jLG7IhD4V8fiRQ
DzAW3jaTwZssaLr+Ew6jt0grpu9zNG9ZFxDcxW4LcHRuKVAo4t8ustJki/rsN7JYYf9d0Vwobx+D
DwPAsL5Phmfr8s5ws5nNewzaVdcEOrvi6dUwUIfM0EGtFTcsXZ2C/7CXYgAIiwKqy2OO9PM2YPEl
3Ym32r2nWz3hQb04n1NU6GRiY9bbT/aNpLvkSbXbL4PuliwAbYNEa8a0LXyyjn8PNiOwZilKUDpM
BonmcHJHT+ajmr1Xpd2tejsNqG/cyot/sQ1mCEhhWK+wVYUyw5wXjUBEaV4+YawdKCxyK2jJB85e
GG8v5vYt3yBmw2pKFZRnPpJdYbR76ZlwCQ4jDTsy/uNv3sgCRLd0y7+i2r+rEmAg4GGN87I1e5ss
RaMDE+oMs7g2PWt9cTaWeVLfiWHB6l/SD6rdlFwRW+HLxgsDjzSVsAdTmEtRpltBpyfDIfS+6hkK
IjwwAU8oz8A4GkOIdm4cIpC5KaqNvYRFKA6KjuRoKd6o+OD6kt4LBrtkOihdACvMhwOWsGRBbcgA
kvy+ML4Wy1fVrGaq6XxhKufe32tng1Sqk8N2IH7PGm/x6N56HjkZnM4k0F74PpNaRMmvN+tTXiQF
Th6t78IoGD3n++JiWFeQuGxcGNF4KzG5dWT28UG1kpNAwMOKs+4fNEKEv/IN9W0dmjyJXfIaB6RT
ZM4tU+SMYqKb2H0NRC241NSyAk5EoFVpFJ/cY6VJmDjLdbsZdbZUTrlHgJXiNilKSQhJlbXOKAfg
apH+rctBZsawZZeguF2Z6wr8M385XCv8gOZqkUiwv+A+LZOD8u/XD7asKo2jYFhCTOcEBm7ThhXh
ku9LGyKuFfJJHT4qlYuoYEWZyUU73XgUKjFhebaK8xWLDdqeLPPfPycXhEMXUu4GKrcsqXxKVb/H
Mph6yYg6skZ+CrefAHjW8V+5KYUfs9P6bqF3ddAkg+EhIk3OWnGqNAqLwTlPb1if5wpbsq+dYyJq
HNWYn2Eaf0/02llelO7vrI1i0fUTNlZ/IPEfL+sabJnq8+6bnK64++xUpssB/OwxTvQmk4i/PkkJ
TL6kkpLs1jXXGmoUgdTMHMj+Xl2jFecWnZ/e8Mqu1WNI/v8u2Jg7cckG0c/Qy7p5YKUsoHhy9kLC
Vr2TvjFGJbcyyIJAwPRvv/fUAsNcwVBkg5vNHv0uOlbPoFC+EAu8j9ps62tEN6TLXVTsRFuqOvQ2
vjVGMOL5GRhgTGw4QKvAIVzNM6LkWN/msMJedvuEO8spjGrxyrsYT2qdD9LxfTNeoW9HAjW/cpoS
wFlniNh2lrOdwBq7Ebgp5xyn7IYr8sjrChqgdTSsUzR8FvRf9ShNHGn7ciJZE6ycUlSg02koy1zk
01rUDMptOHhAzkx9cJYx0wMJgEJ5JM/fOe/i331w6qICN56xN/x9aMA0jvge6tA1PiifnOWVBbjt
gE3Gt0HvalAt+bYP/GG7BvTHT4MK1T+VSBgf+CsThr8EU4tGbN4igb49U96S5lJ7VXkrGo+jZUr5
bgt+80++/dFHaEgtBX30iIZywf0BYWVSp9M36AOe7fVM/H+Pvv66C3QELGDBigBNcNj1m0k7z56o
tFVUIxztF/EuS9RsCXhV4V0rPNtn745RUT87SiHSALdtkeJqNVmv2Wl1vQQCHdWhzQhWTmZFF2Bf
QuHDnXWYN1HIaOPsBYuIfbNoQBJ6rdInHbMnufxIjKkJPGcYY1gM9XezJ7QYm+18U/MQcUoqMZsY
W8naOldDBRh+B9wSBcVGPqAmhlYf6LQbS0Wn+3+NltUAcsRYfFuOpZNz3LXHW72wfLYqSfOS+bgg
eqNn6fMzyFAFVjHxTjvCYeUAN9lX++ztPrECZ4/dBNppsoCtfmiPjv+PjOHHe2aG42c/cqUtTR8x
oEW1w/bHHur6X2NVWOj7gIOV4zPKixCjQ3PZMdbjwp+NINtYUXxHW4xKolrNTY8/zST5dNG2eCJD
Q+aZwfO+fKV5cLNrQyauPcTVHUMOie6krsMtGXv3adl/3ezYa2fTvjPidhCmD00eu802OpVErSxe
p3E7ZRKTL4qrsWdNN/pO99dqoP8IpIpcT8hlYK6qn0FSebMlHyvBYBRr1NtYjrH27rFEf/HmHVna
ZWzfNhK7gpGg6eXx5vagy1BGSsSTNu3YiPgECKatO1Nq/8GdiXsGP8aZcQFB52UwE3ae0+aWDAxz
+h5s6ly60rRZpfKXlvUrYx72pTYfDtkowM1zpAQLT0fiKuGKXDwjPwzA2C9M1d2g45nYDakvMKeh
g3CqRRjXK818FlRvpwxB22JOmvljAMjgALHFXSef9CIIldgdGZ9/ezBXMoLV9A9+uWWk1CkP2vi5
q+ntiSWFt2pt3FaohpPEotRKGPIrXZWASOrXhQdiUglaciZau0hB9wuGlf/j6pDri17J9yhDldrN
gt4mH1PDsvtBeW+LmO35wqy1IWsVVBLf1fFZ1/UA98L1H5qL2sk9YEfmWxi/UNYGBf2Vw2enEYCp
rkjdQXWxNfAKx+0uE0BDbNS8dxq+nv8DoQn6vBU23s2liwQyGFWAsc0+Y1G7SbzpaVQIDLY96oFQ
25jqH/jTvF821DnXBrrxQP9MH+igy4RyMRZ6/1FUqqsthUVENb3/ZyI19jTsqmzuCt+uxstxONUd
qk4V5HCbK2Cg0Ke7oqgN52DfK0rvIMrvctS1Cz3mUk1t2JcaGzZi8GskZOBrPrdl99gHbmybI2PR
fiQl5YvNkjiBZLeMLp0Sa7Er4mxgaaTKW0PD/Em8R+fiq0n/HselVaPoeeAlxuCPbIg0ncocmNI6
DKzSpm66p5FUxLGILPwAisOQEJu2gfqFzOxzSS8HjZAPeILBQF58aEyH/WdqcOTYgmjfq1dojCEp
sfSmqcrl5MX1ZF7mpB+E6WuU9meQ3X+EAq1XnOW7MbMbRqGtC4GpAsa4p3BuP377i1+LTof++qOp
IDB5mpgk1M7/gerhah87sR6rmUEj/2Z6xQd5WIlFFHAo5SHbPGrlLT0FwExjL4kyD/3hm97vj0ln
k3bSuIUrya2O9V6KbxdnerVsqixeoChqwULL6OhkKtuJAAIWbxtpZIlSSsBl0xURk/WRGBXNeK8G
GgSFfbEDYJl513qY32Xsk3F3mqHBFR6YSo4RB4i9gWyt7lLQGkQcm4kJ2uMfAf9g7T3G4SsiBGzR
fAoo3HjfJbshOAQNHsXwdy7SERcZkcGSOXerPDSS4QIHhu4RQLGjaNLCY9Ri0gdvXWzMxH+0FHeb
Iq0XQrnAogX5S/B3tVhyjq+ilzKbfOLV2wHhrz4G65zNXGpKS4mdiDjDlF6FDD2iG8Npz1dI64Lc
qKuEJzzanlCRXfwaFCiinbiWs9F/ssbhUm/dUBsIsdwfXegDsMHfvgpw7z1v5WDZKY/+2aHsiqs6
Hxwt8Cdeb40kEWWQ3f7WV8J+WAErDXtwzk1wKO1tXX+qwFSeFqaqncXdSa6ydBomeyDsuZw982cx
hCSNq+7cN0+7Atwo0Q8KvRJJciXRzKnmBgeNHHfrRqIabUJ6qkMiscUw8gJrYnpBXKmnR6uOLpae
Bn5Tad+Zxpl/I+0mnOTHxoeTASTtoLn+K8FOvPyG6Lgfu34FxJlt8fNvc/drOfJqYi0UUCPnUAUt
VertegzJLSlQVq02UsQoajA8dpZyR/MDC/rdcvk7N+qXM8Zs3R6TMT/608ti+WLq6jacIGfu9TJL
LDK7EvfqILpF5vj6Z9Kx1YAZdQouMVcl5+j345EBMFHvQ/dhOVBR6/EHLqkHPNDRm27bMulADBAf
HqsuX1u9ePru/aU45nif+05kbaI8ZvYFY1FGWuFC7f5leK86v4Wx865aFMYbbdEhxXJZgSs8py4R
kJ57Sc8cmjhidB4E3cvdw7euDsvT/uIG4IFEYRj/gDkRICjatV7p6UxEJFC7Sf5i1hjHvBKHfik0
BiZyifWGiIODHOTPzK3UuQ5YODiXffpCl+B+DvL5AuySKCXTcNhCJmKXeM3hdbIYXdSLNreQwkSh
FJpY//ZpqAwY+eBV7kNx4SdLtQrMLLC5fguXEY7d/2I6WBrpMeWIHvefCBdmOGYZIe/u2/cTM74M
3etwSkb0TJ+O09zVzS1KlyA4WPb1RJY44fsXGct0t/Qn6hdJ9FNv9KIl9IfMLTQBZ5wa33/QGmD7
tN0Pv+mcIYDsVzUsUmT19GPFtuoYamGZq19CzX/6C9YZYfbPp85AJAIHc1hXfwiCQU16VyAvxdro
rMQmJFAkY1GqYpKBOoJKG9n+iEvz8CS5hkDvpgZo9FGUEz8+FqgX8lpc5bmrujwq1lFubaKjfg5J
sLyVXvpRJ1t5mmGnjxGo9Ud34lklaUa+WlmnEwEKNi7K8I1DIfSC7FH+//XTVKJQgE0+AHx/O2E+
VPmqPjuEMm9mue/MqYt8AmOx5fbT+pv2KUTJbijfmR5u6cBxjCrK/GbYsUwzOb9Yd5zKgafnbwCV
WS/b2EOduUpAOApBTRPqzgMGn3S0+szuLui0g+mUj7sc0GSX/itohysNDq6MFZThnJuvmdKBXZos
Rza9OkDVrVMJipTQXEHqMANgZXez0nqgUMJORThUuy9Uf6RlSx6quylxTfLFvj9a7o/kwgRi1Bk3
g+FcV+hetQ3KkzUXgvotVwuVQotNPFxXMHuybctcx8VOisjvc+FpW4V660b00MtRtXPOn8IDyej/
/FRsp+WGNdf1lbhGQJ88ApeDAUogETdB5EzufGEgqyjEPcKLZiYOeLzuje7/3aKH/f+vV0IZG+mu
53wuzQ33xEHXQlISt6oSnVR8GcLRLz6Qtdfx1hY8E9+iTVpU7GIkjHfTTonufgwVyvSt9KD143a5
wL48upUnHKX1M61qW49dXZpuKGfOhpciBEr2J1nAOKBYLFl6IWj4k7hS6VuqrjWgjh3pQ+gJBcB+
TgZFO1K/bj1iSzR9ygrWiqWHCq7W+MChZ9dZB6Rd1krik3Qeq3Dxha9Jc+1Sq0iCdJ2qKOpJJth4
zzBajrH3goMCa8mBi5fAewSmECB+Kt9w31A6Vlts7DQLmcwnYPIHaBUC9ZsysSjOBfQed1HrwYxr
ThAhetQZ9DAtLvdl7mN7rCbc3Mds20bw1pcTA3eBXYfdiDExI1326EuB4Fh84tfSrp3sl8ztU5dE
dCh7g33K/aZVPf9LpK9ZnyCGP0AxFRVxD7NuScjdNK/Y5AhaEs0azeRkaR3Gb6EU6Ioz6jPc+Xmu
4uuLRgpPs5r/grGmnaOpDcFJiB6wM0UZJEYA6SuVEkO5uSa400v9k6eMu6M2tOfPf04JQBqCAHxi
8HjotPh4Z3MQ9XUBikcxX0PpeNBcx+olUUt/NEcVrZSuLOAtoFYxIOkxBPQjqTaBgPbA+LURgNSv
eGWlfInOSPpqE44fDlFcRvCA3XZQSOAcKeC2tPj8U0ssRDblKjGpVi4TxdIdt3AUfJ64vE1mZEOE
+sMFk3tLdQyqLkQJ6k3LFBK1n+Kqy5uOBg5Z5m6lVfA9gLSgEAFz6vsDOsHw8Q4qADayfLZDPqXv
M+IYMsf16vAwbXiQbwGN7CHnFFlea6Hqbw1oi9QeystvSbUUOENhu09swJlvi+F5wG7dG6coZbAR
1WDAa24xpaEFxR4+dX4TWNLRUGWWPM9I9U99PzypiCDbbk3PILz/tNeLd4aFaJ5FSkLDc+HFk6+k
tkEK59mgfKlUi/qcMZNCJRvRmzbQkg9+Y7WRQ/ak/q6ci9q0bUCC2rs4jA1Ma2kZkQju/gF5UqMc
7nrN5v8q5BPoz7IKhr7o6V+0Zj7kL9pFfCzGiXXDWILDfd1IhHzWNCjXX55GXch5I2mOBsFp//ll
vyYsMDBUZ+U8cSzwQGGIXRz5j065EUIFiRsSRDZuPb+bK8U5ygkNCNalALJMfAxbBgkRvvSmf0Ce
DUYNt2LQu+xB7tx4HTEu5ct7Y/e0abO6xIIjPL71yE3SVwqlMzbrxmWFinXICtGkujQk3Fzu3UC8
DjT04zeqMr742Nv6wCYTnETu/CZtgD7fIRqs0AOGKiPcGk98HwQ/f2ka1prjnyfxBe0QHjDVjsIM
SrlZTUBcWC2tDaVzrZf/JjqVaz7vrlEdGPK5uoA5vvwYaTLYV9Eq4wdQteXuIdU3ZY3iDTTIc+y9
zxCDLyEgOaSyAbSjvdYIqT+Wo7L8s4r5RVMxzmUBD2NnM8ZnzodcQYDVQrAJSnA+v1aFpwzeGst/
1daFiOc72Del8p8Thq5INCcO2k47ZWudsg92lpO1y3V4DOwvhdbTaJKM94ruMXWUDhChLTNeqX0H
P3f989joW7gd9v+tZwSH+/C0DsoZU96/FCCmTZwbYyzhW01Y+FmPb4EvJ7Lr2UkxGaLMSGjCpt+2
1h+IuLheyLDwXj46uGcZHR5v5q0eHRkTFNrSmyBpc/17+VgsFKNnyJ1BEy8J5T07QxNmRz6xA2xv
bjNcABbd+z8PyOYIvdwMVwb5Jz7v6GGPeJMuUXG18BRhZ5dGRwCtawosoF+mNFqnfzwYPzd0vwnw
uTDrEEIncBvm4yWXXEBnVhqzvlIzZIhthC8kZTbJzJ8neRo2rvxa7ZvHsEUEHnQcrvI5maMk/7lx
bew86cTIatjwVlNdcS0pElgkdXGkY+eYGyBRv37AHwxVnz36HnzSO61vTvpEjUKoC00Tb6RIVWy6
yCvhd7vfMCMyQ6a+RWOAglxnQvNX544v8TZioEfGxcNjEzQa+WyrUdFKO6ugXT2a3IXUkvXq/zAP
e2lV8BJkn8D93X2LTPQNMlYOMSJunLzt9rlo+Zi2UFaKHsqRx+RGB9zJ+aXzdX8N1VpDiSYzrQWE
lyJwj7UwwKLiW1wrmVW+5HGpzbBp258y9rmyuTVAMFgWfBiMhIIQtNkqOo6D56x/Qt4APWfmlNVM
t4g4NYrq4+3f7HfSGUSL3kApZhDdGxwVRf2FEzNa2ZCmghKsJNClm91/b6goEFjmss5nMh1Mgv8A
Pf9eeUadr7fKPl8bqB36GKD2S55FcnMwd31FcBH563XDVnVnh4f2E2TACjWSdCj18nl/sR2P6KwT
tP3fWnfLOiEePLIWC4efXz2tGfEnUxJafu1nmdpYBJ/pbKCdxedR9YUHu8XFRt7hcsdfr6KJlyyE
uPBnjD0OYYC1JsXOHi/AxDFNZDF+Ebwfc9XDTROYmMO6XN7aH4EF6LrldOwwbKMfeG2+lHJo+U0C
UcUbYfKblwdj89d0zkVI2/hIpoL9qvhHKHdPqJ/k20G7OI+jQ+bmSUJMCWpL7U2gpp041w9Pgg0R
a1qzMJrQtRWawp435JVEY2wi6j/t4xNr3P8caYb4L9XGh10jHs/u17cjMSQomoMHC7rfWjfwxklk
gOPtonlg3eDwvyrk/ojyWbDCr6G56MgrPOrXkih48WXZtdDyXQWutjfxaE9fBjNVY/uu7BZL0JlT
NthbEzLEabEK3ot6MUWEI7cqn64hUcdQRIiTOLA/nCee91ETBiYO0b9Y1E+UxyXlZ6zbIK45MAcV
fw6kPkhMctr+3Rmn+o8SA+4AXcH5mld+jn8vvXs2lgy0H7+462ejhfw8MmQBMScMb37gdzq+/Tad
8C0fPZqFvEH3kkY7N2c8fzDR0IGBXRXVPo03NX1lW1pzQpcVcrPhVYScYnM7/EyETkgN23001rfG
3Hltm1CFOt2r4+55gO7NV+AZBNFP18FGo1yKyo8E8pXNt24vDIwU1mpN5U673u9d8lZ6R/Ar327u
HMKPASrfcAwT4RyxSqK5EtOWUHMYt1iODWzMCcVtviTATixfMtVRDYtOqxAD4ggeflq8FcFvquzY
phR21O+eGF3JkeAhcVfQ2byDx4O6JJEF5enllB2o56u/pNQM5NHglgLSt3sA5GC2XDpUBJroynxn
vXGtk7omMvGHzFbDXX+viv7h6e4/6tPoOwi5ideDjFs1UDTuFX8LBgJ0fTRt9hsYteiMZwvOml3n
P/qjYVRMB/m70uFCva6SfjmYdXIDRkUvKM5gAYDAUs8dp0V2TrUUitEcAxVUqLo0Ef5PXUkCdN18
95eAgGQ5DCjwpf2LcxSJlkzwaO9qmkyc+0Bqr5hEiIIbAr5vEVByEClKjhxNLNcmTSJElQtyyohl
YMmuhoZEKxpSYY+0CE1X2YTnCl1u0sbv7YhV62qQBWOrOhhQEMv8NtmTOYJmRbNcF5/C9sC1ytfx
um16vsbEurXaQvQtgS8BVXBU3ZYG1IkAHljXDDqaAST9v311k72MLi4ATOplwlVKrkXhOMB4f9K3
7YSz2ocf1INsoVuy9XiCdy2wyi1wOpN42WsNWkw4IDYdwzqAaXNN7+E5ozhT+y/WhqAOFyWxij7C
gmYRmwK7NSG7ajq0Qc9jS+xX/IxWhZNNjpZrqfZZH7fcrioNIKTco5l/jWr3DBLhQHGzTdjurZyO
YFjzz35sBopInnPeePZba22VSlrulBCYJpyJ/TiXiEH7kho6Xcv2bPI18Ooc6uDvls8hF9aPKWuE
BFlEzvFHRGS6jXcOv9uY1cNFhfdf2MpWpXZebfCCtVYSP5+A4lOM1br3r5xt7j2g/yGPlzSywLw3
GRDSzoJ4xyhTZZX9JZvI77Jnxg/CDTNK82h9BP2S9CGZNChjyTFe5Bl/ZbofvaN7vl69InWC0vnE
hvB23ClLbr8JUpnS48eJRYm6aShcjilF4W6e7DWOobF0C41Lfm+DOTJ5EHsLVgXm8Rj28JZXQw21
CioN6hFwDWszEz+DqOrihtdC7C5UIb3a4mdhvW3Vogpi26KyauL9UsJqH36qdtZ7xHD8hfLcfpe1
27aau1Bcas2qnHolBwDMxj3Uy/EYL9fXDUVaejV90kD03V0rY3qfWv8ovJZ0FMWiNNxrDikh2Hur
4jgsFhgKxQ8vw2wDSH3se9gAD/UrYUMo9KPBhg7bfVgWYuxYEcV5JmUJ+dWGvMPU7J96gmp5SvB/
YGlugPljPTr8tJzDGyMsYxG8h9588jEpro+KHYNqCkzOcm5Bq/26GosxROBxze6Wyxz8tDPUHXAU
sSFBchQPtqr3qkwZhNg1moFSiD6j88+bWRFondtuQXbd+8IjYNULW3SuzkeHgRogZQwUSZwILMa0
HhA8/+hFcZzyaL43F+fJAgDlGGdB6Ic6/6xhDpoVdiS90MtOiu4o7hudngfRdiUVa/85yOR5bBwW
q0/Zr32FujQaBFlLKn8pyZfB02JvD6u1zQvsgFbj9ziGZvVSu2H/tjX8zm3YH9lrEY/WI5vNiV4K
wOsEJlFj81hqjFxIA2N02mdvkeXsrnKB/miNbbc4OkJpPYouIuxLqB0iEEtt8Tu5sPYsm7tqQH+J
I1ofMYCZahs0N0vu3ny3LHEV4j+usZOXGfXhbzkB8UIR/Bi0GET+8nINmyhnHzuKK1yCj8ZLzcv8
hIC3lnRgoG7DEnQxj0Rli/A1SJJM+wsJ2rnkD/rlqkgTPG8B85QFDW3mAAHTSXSzQ5+io2vGo8wn
fhhWIsj1/zHW7tS7Koxeo6Lt+hz9VZyFuy2WDBHvpGJ5cLjJOVpMhX/qEbmRc75Hs7Vey5cjT/8I
vBygW9VGK4HlrcmAJuH1fwGQw2uuUnGmX1XQQld6+PpPSrJucwpLoXAfDYzWj0fKm2dXHlV6ydWg
m4PIvjN7aaifZiTqnP2qZHAx8jvUgypqpwru3hnfH+VnUEvkbOVOBB4JjnjJ94A8/qeVUuQf1tT3
JE0KNAxE+CD8TFA/rxFO8ZE9NMH1l5AAo0+C/vy4iyFz6xAo+smrM9SXIH4jy0HRin1+MZabcZsk
0nbZiz6plwkhGDHf414tvuwDrJm/sRFuAS/7sN5EjZ5ld7g0vm0f+1dOEHTUzSI+p4U7D35mg97a
wSAjwGNkUeV7iCCuHGUFW2v7MLHu42fnS4PE4MThaKOWD4xoa/xfvkGrTbVJYB4ciPxfa/8Yoh0o
WXlcQH3iqkw+41tLrDbW7uEpbFkwYR3GRoh8/yBBCTsLcokthxmcBPTD/HFtH/aLn0oaEdib+EfT
4wyKRgmI2ry9p7vIZMmAOaw+iXDqyOslhvDVM/ytNcJMXCZi9J/59wTSQBOH5sBMcVYcnkPPYwIG
yHKbMZ4mYhhj51pnAzu0iGDaXrjACnSq2KPbGm6uY0jCVJw4IixOlsBFQZA3PP3Fm/Uk/lxEiF15
aUFYyJCLptwk9FNhielgc75rlUORceeCjGu27yzP3k3qu2sgNyduYy3XAsDIt0UvAQHbiSmxLkwJ
1H/ZENezpUpu9YFcstGjuyIbECOxYQOkKawfhpA9HHVac7pmv4AbV3xZ6rG+WNZi2OmlZwU9eBiv
McO/BVUKo3PIm4LSinPYrBcFmk+Qizwq5B0fl/SmNUSiOmIjqjUvMT6WxLqUnf9oqwz41VD5MF1J
Oflj1Unm76+zUSHfIp02Yq4pjRa/tDS5o2T7yEX98JEDX76a07o98aa++w45woeLr72a40bYqqbp
yZxBFUEyQVRCSOuLB7qVaLkwkHzHo8HsppAfQRkuPsK2pUoPX0C9KgzeX5ckf8Pcj4CM9ULWu40g
itCOAar5TmXeF1Ns799Yv9D4rA9tB7wigifhYaMffbtO8gIEp/1YqQXFmfxVdmnbLwe+F7EVn4oE
nmx40L0F0+x6/CtbcDllGrIBSVlO2K67gN4wt9h0u2ZHm+Qxr71DocvTEt+UZKl5KoJrcbsq7wx3
AtDey4wUR4pCjNvstU9kBUlQ3CtK/ocv+ETmQWTiTmkPimiNU5dTKP+0FwgILpqbOt/6MEtzxI35
Sn7ErysxZUNzeguhKEEAKUzIw8csFP8a1RSBhQuNTodyAtvmtSkadVMw/mhQzeNz0dw7+HL2Q3o0
uHfYAkUoOnUagfgIAoJI7R7Ehf5Ccs5sdnYEhlzVorpnk+0zy52iYRfTZjXOMdL22Xgi5vnGxe8W
wS9NR6Ztzp/2T1uuDDsEJMDS/pi1ZXMLL+T3QmK/66CUPgglt/JT344rVAg9mvIxsS2AWUZjblQM
2NX3qHjDXkDWIfosnnGRU5G7PeYYDP3SYBz7kfS+B7qv2lb6rLm9WkPP7TPKgwIcVbQ8rjrB0vxE
mljf3TklChLqJlp2wXQAXX2OG6Few+O4gTPyGYZrRrlSOX1EQ9b6n8yW9+y5cQy3+q6S4+qOogmQ
9j7SFXui7S0JSmdD1wlBdwWB7aNCHzai0HfBzK5TyIpaN3iOE0Ubk+0u2DchEYoS67O4d9nAWiqT
LIrwFH717X6SFhxROHkWCL34FDyZe+aZbApsGjGVouyD4I46xcosTs17miQfavOFJ66fZ7S4oxq4
oy7o3Vpp7FRkroO9cuYSHFdRlyngN8yRxcSgZHAHZRpU67M83pyANLj2azRuqREvjHSgC/5nf+dy
niLHORlG5H0WLfgkso2XTRD6WG6/OZXDFGEtV1XhDZaf1QSHdxc3HnDKzPw1jZtuPdEoVtlypag/
KEL52Ks5KzW0zbQJuIMGYWBqed/xJysum5YDmLm1Il2fDYOV2dBH/sK993FPuk9xoQAM5DnAmxQb
ijf4ykBROUkWCRl2LaolBd49gzLPnKV93ZG5DQoRQ97P/ri3/TaOh1LiEGmM+YsG1/zWzzrE932G
2xnqiMx1rirU4Nd7Zpxd1KBlrpwbVEcPatnERIxihwfAQEkN5PBBpKER5WKKR1kpbSQJspHti/pw
KtlNCElxkVUCsyl0UjpVao+j64PPWsLiQDyVoQ99jEALlq+1rdGnhrisIXwTzEJG77mZWdVRJLB1
QaTx81TfHdINBmoC/eo5KK/1bheuUoUyxonR0eoe9akYpKMmxez5FYEn7jKwwyw1voKIVMJm6/ew
RLH5MRp9me/iv5PvCcFDVrY2F8aL0NYQufIrDWy8Owv+yagOnooO/nJn1BK5puPtHw5o3mjPidiB
rkl90nlY5tETJxi+vtnOZTVBJSuMEQDwkI+jDcWuP77XZsCN4Xya3P6UJamueAtgguCegKsVHoSp
jdZZ7hIvzp17W/reLb/d9uGw5U6Bce0jJKkdA3/pmz2F+bD52U94egFlKyZ9Co5YfXSr0ftvShhb
M90jWpZtvp3EV4J4hyYg5KXfn2b27znHs3NE2Smp+4RJq5Z0FpmYBOEEl7AbI22cQLylRl/0CFHw
aDMyMvFML+X2PTqZ5Yt6TVXvYFH8U4fNFPC7MqcORpkQXh1lL7W0WzGd8SEP8jAe5M6/gCghCdHu
abM0fMIPe9r6pYUUmyFToOEn5buP80Vxx0wZptFoYklrly8+mv5pRviC+1PRU7Bc+4zIeOUdqCVK
K9Djzi0UoJji2hb6l78TMCdowjaeQKv2Vj/xs58tb8RqCvcBTMVsBeQ/ZaP+vDb2l3npIJ4+mNTi
zYUuXOpmucdsdFk+v7YNyAvBzZngZ/mL0ul0SGJmi/IgpP1yYWhuGsFBcPkRgUX10QAw/c5hFZi5
vngNRT4DM8ORf18CEnQjv9N3UoZQJPuT5KfFC14+DhFstwdKZAIMmEz7jHGUDS6ny+hppuZApdzn
sxhhnA2tWjrJ0aYKrh2L3MQQEe1UzpMzi3H80BKgPArlW7m6wNKxHNpCeDu6iWVshV0N6urtqOEO
Gdh1m852sAWjYsqxOiH6zwHrhUAuOIQmpiIyvGPfzDuVS9MBKpfFum54mvxJCO62BiUh63/WmmiS
boh5IwO1L95zsgxejhz8OgZWfEu2Umbn1xYSfn3AHSWgoSM2YXVp67daGyggGDQP52rJJ6+p2iol
4qy24+rtlDg29aOHH4c/hi8EN6ysbfzCpEZeY3EyHfVYQg07ZyU0vBxf/JKErD7a9r+h7pFo6qiD
pvT8/Fmr6ZCZC1Lwp90DIeEPBBOZtPcXD+zONE5pm1nWVLUF3wRN2u0JL7Q6U1mn53sUTeX74aOt
0ZogBdGORP6lZ7CT8abfALvPIlzW4u20i00pnz7IMbCMhJ+OHquSk0RTqczNkOHjljg4dWBGwft2
DPYZ9diztVWZ8LN2fxd3VsX0bF8jbjmQwLVNdF/RSXcYTu1EerO4PGFIu2E0cAwiLzd5EoMoWsuO
Q6eg/XRvtaY1pmDaiGzChpntwlDGFP8DQxmm/9hg8lkDp6fhjklQe88pjRrAK0e18C+nl5N5vMuZ
iBIZR++6NMrv+mF6u2yexNMFSb6UeWKhFLYRW8oycwJ9BFKguMiorRelr+jBezLLlXUViKj5AQ0t
7oXn5Rl36S9dtsG5VqoYkrMtyL1CgoMD/Zs1JGVIroRvrRIddwfsa85avIJXKISyQYrYyLTYdm+h
aQ+5QfffFRYdqh0WYa5PDjD8cTMLElNmvZUoGCXQmFs3prdyepMlrMz5daPZidca10HqPWssIKJl
fDpWXabu3u2lOwiEkROlWZYlZ01a+5mJDgZkEcXm2GICC03BmxFnc6BXKMbUzgv2tY6yDtgrHmRG
VZaKmSGwRupCm8cp+9oeTZk+dm2mBJfQ/dhpJbpMTZOG/ZdnEAt6mJ37C6267JLZxAz/fpaArxxl
u4+vgiB7mX7XFGkBcfcHs0fEK5ZHXQZ2EAE9UUv3YgKjcwttCLpMiAgT0mmouQfYUyUimITSGP/j
45tT7XwruczrXYuVh1xwfmKZ8eJMsFv0isS93cvvAFAhof6OYYKD1dxd5lJZjnP1j05qi+ZlikQc
3OYGoXBiBphXFIyk1uiQpFDad5XA9O+QisDg0GEkea/1mjVZfWnxtVlZWSkHdlD90io8WqdD+kvO
+5hBwTzQG3PS6qNgLE7T3Ih6IhJH/cHgLNvBvQ6Vato8mUdl3EKPJDHBM87wBa8GHadhnNTr0Rvr
Q0ymfSIqKTaWMSj3O9VPasm2HwUdM6eBXeiZkkqjCDHXMehJqhwh9NvW6DVpEkq77CNuqrizYz2I
CFZybPQxN4u2eAorpGaERGrTPuAxdy+XsGI5I7gynctl3jz4vTkElKISeDYYT9+VGzhwtSZ4KRRb
JltVOzKEM7BjXzFNM3nsMFOrx2/+06ctVk6TXAv3Ju7UeZvtHob7MmxAXntcAartzlcr+b4kzBk9
+2UYGTrLcPrLJtcxF9S53mw0mLTFsBSEqFwuodERxXrVpY0I3ngZp5c4ovHXuHFZdXddb2snZlOW
s1QNpoFhe8y88zlM+7US9dDL7613RkSQPS2+wSodiHm3w1EgRxPdf59xn5nmmRGhMseI1ijBa+K6
I5SOa5c6msf0t3Ltsk2+3vjNLIC6PtGTpaO3bkxKJsjd9LwyosI6Pkl0bxm/o9Cm5Ka7Fj8bkUn+
9gABZVi3SYpE6wZuJcLzKVljlnVPya+g95bBdT85DK83lcartHpu59DF9GFTwXEiV6esrPhEZRBl
psAYLPB2GZqZIvX2XMOnt4T+ljuyKL35ROn+6okU3FY05FIKixe61dCTAvsWCQMNRfLLDYGoe183
v/IO0Z6vNYJwzGQV/x3SVz9KXDwfd8vCytGWbX7s4a28pxSXYYYhEm1Lf7xf1veR61f0mUD9sMC+
Y1DBVsxRWMQSBz1cNUxl2ht13WogYt17hHG4BU6UoUCYnF9c1qSsU9C92OC1VvUFoKAw6QwboSk0
WFDR4kGEKvfQoWlr5qdJR8TwpND8bYr2XQrQvaIEPc+q9+b/HTo3xXuQuWs/38+veX/4/xmk0qKb
NKHrwSEUuz80GryMANlujhxUgJxVwbreJmsokrTNZUBcFEDPcxDfMI1VBmJ/y0eLWWdIurrHN8fp
z0zG6U8A7HUCGvWxKY+yW176DkElGi8S7hK2+kHJCMsfiPfxVIun37Yw4OwHWyOAGeQT6Y1bfewE
5cuGgI+BZINgt0xVZtI0Rb94Y9ARk2r4ZAAVn1ZKR7TdqUwO391GdEvlQIQraOpAsuMzVA7hIwZI
HyPG51g29Ri/zpDsIjKwZ7lN/qloUefKDkTJccBJEnOs2gsKgbMR0CZGzuMrfqaes2atR6zvEWKp
P5OKcdDe/gm6kvvhqkeAnuqtEnEgbtc8KuYJIk6WvHXj+Nf9FyJb1KUSvW4VKF1aC+ap9LGlxvRj
QC60gvGg8p4lETOWrzkBXkL+kaiK37H1xstMShw8D9+1qyFtdhanaZlXAMWMpbSr3BziD0k+kW3R
R1dW2bCn8tcZYqiOOtL9Ge3sARAugG0vvB/IyZff5tcTmNj9Q+wXMdp4KXkTRHX8U/uXpo2UZY8n
ojLc2Kbn4wrdedDp6pwqUQ/Ra/+qxo8CM/1gEQj/gCruRqFkAnSeQE5CRv2NZUGl0OvPhlFg7DlQ
+ie8dUxkMmqiZYrlroHm6tEOviJWVIczPwEWzbS9BCtOVUuqXYDOr3JV4YWrzaQ7CU4o2f+fz+1K
e1+QFBX3Ljh9S9gQUSnCShiAU0xmssgGi8GNLAiUJaQKPa+sROE8TdutwuMmAjz+8m1M8C4dvPVb
Wo+Ky6CUNOPKkItRhu6tP43iCglL0eSkPVAHGcvpC/UvUs3KZXA/5K3pLmWWHJzTlJL6+Ou8HLRM
6ke2va4b5CSVpEZyWwLNFff6K2Qh273kBS9Sk1YHceDRnlye13iJVrnqpGP41X4+0HI2Cvjse/ip
6hionl1xl3d61avenf80aSvs19xaOkOB5s4DeJxSD+7RSepvwB915LD6pRHIndLXgqgsa5Gk2Rl5
UwEEQK1ySobhn6P//PbKuBE6i6YtBb7dmaiL4qrTmIjzCJJPcZBr8b4hFpm+sqT1acfkjKyKBYtg
d4gwbauGD25j5Anmq99HQJyo9+fqImB5v38yPaLNc3tTb/onVklnyO9+F5fBYRnNJGptOAqYs0wZ
LmiN+Hzdrh8oWX/dJhDAzbvNMpO3H83CGG0zw14ndl9kKDaVf2IaUDGWZDq1QMVlqfK158NL6AXS
USQgOoC4bCwrUmE9eGiNkLAYMdU4vaTBD8p7fHeARzawgSRf/volbeEUq647FIPmV34sQhVsy3WA
UU544c3LZY9V1KKWI+We1SEpDwSehPuIjpVvKj5JhP4fbdy5FcpgMiStJ12Mv3pXj3sno8o8jNgb
RJbp2Uq9Bbty82H2TZodd0PewTdZ0Y4qGtd1iLh1rh/PMscntvMP2Cr+U+hlhmctOIxQ6W5WDGsI
wHpCCmJd514xosxxsFQkP3/aWH2CMTkrk38yFAf0Cf9LexSrXJ4ZPJK6qalSw0dmfkAVUXqvJD38
3++dhs9bPDeqhA8vPjXYIs3hH8cJJiJ+/xFRc/TfeZsmvaids5rlrik4jQi15ze1j6vk5Zi40VxI
zS2vZwGrojvJC0sYeWzgL2v2t/3ipJXqkohm3JkgWTUvOa14VbT7dmDw4nZP3DdRrDnAqoY0WJt4
Rs8EdBR5DTNTuv6FrZV4vinvwSzR1QJRzM8PnKFtfxTAk1vHhRpcwRR2OkAqIoRGus0jWkC33LEu
gIR4pf+oTNDSmlMks8VLD9RTBROhUTTzANUrmPsYQ9WOcrIZ6JKKcHga/Qe2xWMqdZg6mo1NlSfl
fjeTrfPfHJEOI0dLslxxoCWMOxPqAkkQ6AJQ3xfmkcXD/mVkwO1+WIP6nm8O/99XTICTRWb3hnhT
5Ecdmba5LTu5mnqehGpMdsi2EGKKEZsA56WOIecFhw7nps75DdF9Z3KGzwbvkMDF5ppoBH1ijIO5
Owj5dYpjJU7+99A62aTWKquPXHMQMQIuij7rd6+QyqEJrfnhVJRcn8gmSw0ciya1TJ12VjgdF65X
SYFLuIHu/E/tucQsE1RS5E58Gb21NexnSlpmXthdq45sxQx3CQil8MXhI7nR8TdxZs0VRUGocXTj
xN4TJ8i5k8zBDFmDNtf1ywTAtlibT7YeDbatUCp63/Y323Sz5A3BitMrLTe2UiRH32ikVGk8zQql
tsqYkSqD2FfWzt9t4K2VyDc5yIGsx299cjI0XHF6GPw/Q9zBCEx/EIKAHLYbYychSb/o4VnngxTn
z9KpKCV/hexHbx+1p6S+PtBzIO0V0cL4MYYApusLzxK+iPUK72+bWtigkFJpPxQMlDIGj2WDK2dg
PyIxLrLdLN1xINUAbnI8ECBy7IECMoZzhngDeeBTiFy5OeY3gQElD1+6bi3KvU8Nt18Z1PycVpYR
ZndzGloSb+KtPfYpDmvh+Pe9ggOf9Y1jFYm+uYnuJbGdNcIp6bR6No546xCkOF69/M9zzJOZh70/
kIBcYOuTSwbaF1FncSCUuKLG2pdlQXuYQgdGLW7VgRHBmqe9C8l174maMKa+wUrV0sPs8xUFtbw7
7ZXkvs/9bhyj5U32ryn6ILielKWQbnvKkF9YlAiUvuyMr3UeoFNozmM+Qnte7+QSOXioZ++KQ1B5
EpJLCdeaa9uiI5B9zonMR+bplaZzGEAK26Z9lulpfuHm0HNeGlXOjNkV0BhPDrof81tcFt9MN+Oq
BFVs8TNujffUmO5Rvn2f+yEgdjuur9ai3CAgR0NVRpxVjVz95GVRPoXyonDInvZqhlvMpdinavl7
lAnlQ/LRkDgVur7Ki8SsTsLCvnNR5gOwiplgrjPEHj8qPAgQplkkFoVomrZF9MifV3Rl6Zm8XeHW
omK6xDgEtzAlYMn5YyNefuumLI5MjO1YDn+GBgAjF/wWUnSzcQf4EudKnYH3KOGTa+vv5Am9MnFS
KJZCa5RGOoFg9OANj+1H2tn7OVOtvKBj8crAVQ5zo4CIJFgu33HnSdByuPUwQFaSkGByqf1gEPcl
jrD9zI/edpI0gDHGIldsBb17FoxoAefuHJyOPkCi0aMJPqafYyn84M5n76idK/m6Sqqa9ckvquzK
aUMpExOPbAvKEhzh8spizRw79wjbIdmmOsUwR4rXuzZQEcMKicpN9S6QkxU2L5apKBMHLSffVrVy
4QtOWH9tFmEPg0QbOLjrAh1nxpPbXTnoEDFJBRA0BC1aZxVCjA7KQplCP6N5p6cS+pL6kKfpKgiu
0TsQdyidhXD5mabsY8Sb7qvoCYT24dg/tIayNV3qLOtDIkLEd8IAFcu1IaWvE0LD/4yrPtqn3rxI
Ke+6Cj5l5GhmYNfNwg0So8+RPXYtaasPfJoLRFBecpuaxuZqc232FN6L9uHH7KT996+WwFbJ+kA+
+RTygPcQi2YJ1IMvef4eERi96l4oCQWhjbNtHesxb/edGERt63POhP5xcHSxE2gKY7wK/RfwI/DZ
IcQO5PDE2HZscjjqEG0C76hrBgIHqPZKTWMOUiCIrMfNSv10Z6f4zVm7xtA3Jezaa8QZpnha4AGt
TqDdhFhjE40hBkkH4S1KGcCtBHJpwxsCzcdtXapnwOfqQLvv447x23nvaaX+i7q6U7R5XkraGYJe
iHx8yv76XaAX0UvE9nK6yMTmYHL/La5Mys+BspN3oDbgj171ZVf2wjZn09HJ+sIHfPuh/YbfWys+
kOLesfTCRYct2kkj19rSdy/ZkO6FB24vqRDXsS8kX1Qn/NlNbcuHr6exozl4iKLUYmRw/CK8Pbfv
0MYL4GNSmNbniccJ5wu/0ggc9Xe908EVYXFPPs1DmYRT+qui0Ad7w/w8qjIoJ8OwKfEKeb6WdLMA
l5Qx5iiAykf+2h1h/sfv4rJ09EVD/u+YMbHRcOLishaOJt/BAfzQ6cpMpqGi0pGX1Ns7JuZeShPH
waMConoFceCsjizYm1zW+48Nl7EX0QykrWskbFlvUzlS5oK3EZmqU+NBFbu7EOBG8SUPld5mS09j
iOxwhFzidw0dlgI5M5IZ8dlgoULnOGME/d1uyDlnZQ47wr/KqK14afhI3E+1/KN9TL/LjBc9hzaK
a44Mh/cV7/pvNfxauyAUGr9gGq2Mu3yKNCz9sPfagyXmYUP0tdYApIxm2k7fmkHMkocVvLKtPWcH
UH4WZSrneDJQQV/gr+8Jbh4ypaB5TFttrUjBURrSm6ioa/quiloJNng592qqYQGz03s8yLJ2mNxS
ZEHh8Au60b59lq1ClhjRXDuUbqDlcs7wXtX5hmDpnKzR2LzLvnD6fKkI4BR45xW34dwR29aqVivx
HmBoNKsf/BXTZnovuOs5QhjYHZExdTKPUGn5x+ciElCQ8mxHgddkKaktykVN0PKgmRRJdzE4B4EF
0FRHrtozR8Bsv+r6OA6oxDV6HKW5nOowoSHDjEQSUFa1pfjYJrLCLhMIIZzOPt8J4VQzpYE9I9O1
MzttG+UaW0sYq224wnIpksCfYIc9f8PrufiUlC9n0kifxY3+YIWSeJSYjs7BjBUhKM2elX8n9eVA
YJafEHdvhgIWZ7Aw8CSRnsqenCfkNBtwHmh5jJSjYapr/UC+rzUYNiGNIyV9bfcpR6GR5WOdLcjb
vzKJO/J7gRYmhm4qTLSuKpjAzRxS4SOvZZi+g5q5rYDDQ+qceupmcNU71H22Hw8r5RgM0MH0pZH/
F0eqCfcqPhv4ajljuCiAYSDWvTipRqHL8HCtH9bnvoZN9hPs/zeTwYfcOCEyYxTKg4dhqw1cJ7oy
13ReBO30rUsfDj1qEbZet6GBLTUJpGlypykhvZNsYNAYYBjTCLe/N6CZQNeBBSNiZCeF0/qMRb94
WxDcki/w3q9w94NnFZhlxxHGvxduNrulFdR33uc8P2XY1UAOiPlq/Z+B1FPMC027HCxipEOjJMkk
+F5NpCpoGM/++MsJud3GZBaOZg21SvJZiHhSeu3hkUtJIsvzwBjaV4um1Va/remvCSppcWPLnW8a
6iHx4ofVwhExfshEQINfByaGp4no7JcKVHQ35PzGP/mWTNr6GU5h5ZTCRZaWmuNmcMbPdrJw6V5+
1ozbVENHCPqzCCWhYMc3HvlrLTeGfE4hARxrUqt6h3MCykMLuOeoEvORxfnV0/QtgCnS6Dxake0B
KQWmmkxVurjFbYqI3JtNw8sUU+/kcmq2ChxFIfoeFgCRouX4IjwtbRLkHf0e1zu+6qMp4TKNrqga
D2i2YcUvnTeRozZWCwT5zL3O1yXW7z33716OludVBUssDwE7ZwO7zXg1sq3yEQpdgx+QG+yH35oq
pq+ZwmNmXERAg8kX3ifCkeu4netNR3XDm0vUZ+vUG7WNCrmVUlQ+gnNHAMHrjF9aXR1glUqxsymW
z3GHvO7KAGV75X4Fyy3HuQRzE/k08qvk0uPVHv5RtwsY+t4S4HdEJol1ufJ02B1blToKrT6jUyTO
PldJ01AJYbUWJIxgqyN7xspU4buYCrUs07WyxjZE/8F8ai+jvYgwR1SToIzv3WGEHauJx9xDqauQ
KyXI2eB1cYseiq5nw5q946xy0ykpWc9XRaZlF3olIhtGLpvj+NhXgqClQ2tfUDkIldAHUatTwYpI
fP6Yz4xKG0SGDd0WT7vNC+/qHQmzzWkazzUlpzOmOferzAFPTsChle6S+rQMBWJCb73iI9t/p+61
QzDIAPm2GnZh2DC2bHUkfMLxfzw39Mo8r4RxWedb6W2tdG7Gt5Qytdds++FzyoPI5eowmtzkv06U
bA2bLunuc0OHRnC9k2M+b1autDISEAgnwSiSk66E8jnr/H86U7y8vocHeOvAuWEDgoMNyM7imL3j
od3493ZL4hLripxfwFBKITz3fH2qJzMoftS5JxsaMKy/+RE5LBmEq56IwLNPkCH7hCVzLJId3ed2
cPhDY9MAq/yHe4E4SkLI7h1ICsVd4j9m3Oxx6cth93Z4vl2+7NtVWGpHmA5eYdsFLBLbeob7Qsf+
Z0u46pJEZ00gM2ahcFZFMEffXHMGjup6IItq48kcYVUxnxAWM0FnvR+yCADmC4YECFMRFfZlieQs
Qlz2VRhKPVywmbQ3E6zW3REN+uQnEOH0KTcMAImfINbmu+KDI/HM8jZwTmSgkWwKmBCMcI92JsFO
Umaw0oMZDCHWTTLQpI75A8bvJ/zj9Bywnl4D0L/cZb2Wbufb5p7jZA1DlxdslNLUOa6Ss3vB81Dj
jXE9jMzVhcJFBfG+xKRuSy5/rutDcPVb0PfOeViasLgpEWD8pdSz3S6KMt3+8Hs02DY77sRvdfai
k5Sf0v7QnogEKVaTXEdkNJ5EFDp+HUvvTS7vZ7gqMC2rrVLu9+qBPI7YIBRWM7J4ofaaeu/XQVZI
QxMnUJEdAOY3FgWF+EISQ616oMtu8axfALs8+EbwAehOW+3mjjiH/yOHVyarXLfsOraqGfT6UHgG
zNJd1POS0pz+YmXV+zdVtBJXMXHdEwBm//fDgFA2xMkmclgKZJgPnggIaCD6vBGMA7Vl5CaWNYde
c9jPa8Y2kNFwOGsJKMQGmHCcCe3aZyLoXdJyTbJpvInWex6RDqIGgW3KAg0CThIMj0pzgwssGL9l
q5w47nD8zBF1nN2x/5/noWioFElaBbP6wWnbh3WlvZkw2OXAJfDY1F0vTIJ7OUm7UAJAN5UKfVrT
EaXpGSNLsOgQX3VZTPslOK5RGyTIs7llcaxdqppdSnhQK1wjw0+34SSM7RjpmuY8Awhz4C3Ty0fP
XVHPvH0LvB+AXz2J0/8gElEyoLeZl3W0V5flRKUssvEma4sF93yu8jEVfY9gstUVSI6w/uJCNSHg
CtKsYHBgwBRGBPXCysYTQ/yHHzJ6S18IEy99bu20cDEU80J3iE0Rr7GnTEBvoRIChgpNef/YpNuX
bqp6fopZMpkJ5x8Zg0r55BwMIEpt9Igg4yNbrnapsWAIeIeIb2Bxb3pfh5/4PVro3PNniP/WFx0D
NV9TejlgsiJDQ1rZZN4x4FAImX6QWjumhh6kuH/wYjuL60LaiDrIA2YQM9vJbjTQhk2/8U7xWXq7
8w1YgGMwxvrAF4z7Ohlh4DVClQzD4gbAuTJ4diodtbtt/8h5UIN5WuAmrWpj1ii4ymtUpJ/q5o2S
2N6EUwjq+4WBrGH03tpm1mdzOvywH6EuSXPlHJSPg416BkrB8mvNjGYcm3U3FAhVNGBtA3KU8ddD
BjMOqtj4K/yoT72VAGwUPT0qJzdYWIhB6tEeLVZgIqq3vraivYYIlsLX5J3SMomOsysZiG+wpYSC
9yWjr5XFW9FT20YOr7IzkFevK0x2398BCxos6f3+qkK0X1yp10UiFH1p1Bt8ZsD4DsnWWuBf/cDb
bAdnhOGQHTpLdyGlQloP4p66R4X/l10iBvw001PHpWUiYWkiEJ5CYEPnH9iZSkB6wegnUahihjfP
6pYaUqQ89hw4+QWJ26ba0tWRHmurT01MB8iiEsEmPq6b92GcKHmrdBGiY+lSiE6SRak4p0w6CByM
uzXbKqzJyk4pdNhlI/8i+ySBxjxDvG1CQ8FPDihIo5hRazikET+fJcpK0Se1DoURZ8dDidQXv0IR
VdN/wUnCngcXWzlVNCAlW2W1GNuZMc8ErEiLXXQCiIHtIsRqC3S+NHKf3JGJId2RTIB4oF+rTw5F
Nbd6+aLeDvfgknPnbALkwsC8zETA1NZVl/GN9qrzLkLQy5/fJq6fkUyIvmukJT/c6jQxV2gnli9k
l7ukvxHVlBcs8QxPpov9gYmFkE/JaGL/Mnm29SARq69qY+WUwHQncg9JPWn+A1iOcMtUftJtOLSk
d27D0NrK3A+GcDpkSgDqXBIaTTvNdr0RLIgO10k+ugXJDbinwvgzqD3RR6grZqozoCLQqk3x02OO
d2g/rx2fIs4ma7pOe/5a1mLH+o58I5sqmZvi999MMEELTTg1ice06bcYKtxQEc6+1knSM9OHmdke
aukvAUZDGaJ60oEIdqYNgk/y3+XwmCq2cRqcWmFKdN9gTr+IMGFqdMiDSXqiIxJE+fjry0bdoHtm
cPaEu5aRBSnVo74dgdBa68Dki2ALshcn/1en+Xx77gT2Un0qAINtLlQxPtaK1QYc6ANqdqkFdWlV
aH92qBsXd1eDCaLcr1E0C12moC3ld/XQymrILfFSzhmF/93rjmfhlarKj/PM9Ts3W8Bd/VkkFeaT
4LY8M8QOXCH5dkT8/IIb1qHk/594P8kg0xsS/5atGEy+l1CI9vquF3vwTZmp2V9yJjiuInhBsI6a
UGtGzzOEO5GXtirXMX/k5/CJ/dEtJkWFFJ4f5gbPbtOiVocwxv1IBFVM0TxEs07TOPIWlsyeUx7T
g4GfM/wtRCNkHpZcGdYWvZqn38TsiP6zP/06xd/kycm2JHsfNb8l0wS0sB9brJLnFik84kUqjLQq
GIkuhUAn2T37f4z2UPfgglA9zSpPjClHFmjkEicSZASre7lFg2iLzWK05n/Zu/sVlq4HBEiW93u6
iY4VMzrNzYCwxe235tOoBhPs/BS7o2l6gZavVBLMzbUsv6arKD10MMPhhmOXUmKTzscyDONXjNsP
wKKdeB3f6sXMphtfLxxJth0ODmyE2Jib8YfeFfGWvxISJjRf7jGg76qIORZi1D/qo6zPLBMEYy7Y
kGAsLCfivd6nGSQ9eWLWT6C9N50Wgeh58WFFMKHoj0XO5Dr8ZaOUsPiiYqkUrXqriEg+X+3UI9EO
ss26JZFZblJw3KFYWdCx2bCwmTFqQoni9NBQ+HIbRtKF1U1xkY+aPjzNC8QN4uw3b2I2tSmyhYb5
bVBe5DqkPmb9aymE3ELhpnwi6XbMfuywz1use7mhyZ51Oy54n2v6cYbe3l34oSqITomdavbgYdXS
fOAL5FM/jYzyG0d312Ss4+mb9BeGKFn4r7BgFuejSzN0QU+uzfC/MNVL8rOjsL3r+t9biU9xYBTr
1n4ZXuvDhosNzp7ZFQgSop3w9wscs1+fsRA39a52gYPhYVe52NdeIPwstx9aUzmcp/p10BQV9IIb
+ezMrDSX1mPf+RSF52C7JD8hbMVsCN+fJaYWQC5EkuUXsdHxjOtruyNC12oO8Kr4gePIvuK0u4zl
tOiHcIcqt0BYjbXoEfJHFTvN8sqoaluOpS+cyBh/I2w5zWC2KCdcS3c+6FfkITuGKhCKIr6iA4iP
CDJCfdjq1wo1Rmwc6pyUdA2Mq0wVe/O/y7sIm7JVQaXf9qx2hQfbcwhsnajcpwCqKHKIVJFmj5aA
SoB7skXrtB1knHKEhh7PqjTVWWqZW/c3waemHjioDdyMHbLqjDWUQlVX+q4FoCk7VUThmv7OGhAh
qAO/eh9r25dHYnM9DJqh7yHQ1ZbGbZODxfUv7Gzf6IixaCkGk1w3bEf5I+1jzMWRPWTB5xXZHIiO
vvn9coHlMeiAieJimUbV6r1yC46sscAu7pfl/2abfRNG5Cl6RpPd/bMVHBI2ooSD1B62JhUVG3Gc
SUEyrcfzEjIN6ym1MdJWFuVSCTFvZpge16RTcIuWxcY6nYTKbo1D7N/I+qmomoy2WoEHYSsYRDvb
Rdchf/eycjDTHhCxbLtu8mUNbGBF54TT+KnLpcXujHIhdD++vi5B1xfLC66v0oa+qXYUmw7DxZgr
Hxm6yL09rMANiEDFfRTxfH5C95SGC3A44y//nsm+8vxDmKsppt6JcpsEBfO1h5XnGnXjT1kidlho
pNRpYPwkAjmd20wp4kOmq0BekOEHmQ7lTVOE8oXNqZdWZd0WVD8p5/kA6xQ+9Mr4MVm26S5qA+da
6MfC22DZ3sJ0R7t6rJT9EooDztmcsb7Y4LX8Y/FJzLU3TUY/YjQ9cUNNLgf1nQoMkSHmEBZpv7W5
7zVh5CUxWtSCLAezdTc6mjz6NaVx3wq2n+LINxnx5AGCVJ6Itqi7qBNadEcbl/xkYC4RXKlvdEFf
OyoN5ykmOnMGQTE8YA6m+CZ5NrSN2F4b8ZQagAMah4KMjGUn1mgxho5yu+OUO/u2BKiPtn0Nd8Uz
EemHWvQPQYXxWTi0ajusxemFAIiDjqntESRqBgLJMinKjvxLwX1FD+hnXrr89l9he+v9kBV1+cwJ
Tkr6kMZsBd5ZrAfjotiM6Z008li9YyM3EQxqaEDwAcO7KL001Eg+cqgYpQcO1vEraONDsokg1pFO
Y+rTxH6isqjIrwB/DEk3bGjk3o7oHCY27w8nbL+X2yMazoQijZKfFlFLVSZu5b1Yq1pamMRs8I/P
BHA4Iy00GYPf1k8ztK9qA120u1DAskzOhl6WbUjuWAdeJNtuC/VBMKT6TcsfcCzZ0oMG2+xKKrN+
7Ls9LaGovMKJ68XsMVX2Ehuj16vYD2LekqzzVq9d+d0Z8G1gjjFnz9eC4nuVpS0u3KRs+4EIMv0V
faN9bgRMwKKEakTThO8n2brzkHLRL9aeL3cTf9rIVHzcJChx+cOQbWCejEER+GOMNgtTXcukhLuG
P0rJrxvjulcJRq3yqIobOCP39ZvhUGqxdT+zBCN2fQ5aeCJSqBmayjp3fYYQXVTIcGtvdYRh0z29
KhKFQaZjLpzgeBkKEuQcnO0XaS83R52f8Q+FuzYAO3x2h+h3ObvdjfFVUqQm7azRUxvesF+99/wC
1r+H/LM3Tolm9Nhb2vRBaLk9rtnuR3dfDqW3UiEmN9rrCBJTKuWvoHEIgLjXliJ/1vP4OFcXZBXi
UgjVKz4MwuXoXOZ7fmFsbHepsdNteqMHtxvFClYh/cSuPzUI9avsGxMr6hjHd2O7lAhXntsgxj1K
trGBnzWz1O8xRBd5Fr83uLs3tsh52GQTyLgPWvq0BIZpWXcPp6B26OkBDbw/Uf1M2hE5hDecBgF9
VrUv0Xi3xC8Se3HedvfpkKqI+xQOqbCchdYwLcAByi1W2pvlGMwkr7R6Wk2yd6m1lRUWfKX/nPqk
h2bsQ96LhSFwQL+dB8MVxzhmAfbBje+33wrXLj1wMotPOS6WgJIaoU64qoWuOfceRsfzG7rU4Cz/
liAlRdYCVr9kUiGc6yr8Qw2NuPzQP3iFp6jz7Yw/pQy23NDAGUTJMJdLNlj9+DPRGFNcx99wPPXJ
XJqesErTENn4tVTX/225gykUjX/teIi7hVnZGhfJhYJH+kVBUSLOh2E6SodlAUIvfZRYRQ5p1b8K
BiR9+1tU5J5pIoxxfeipb1xmmQbrfO2NOA4JqBWsde6UC9Z+TIFb+VWQbcTm3Nca8fPZ3CuCjPVR
oVXZo08LyQ0TUCm03CWT1Ihf8SCrie+g9DUOV8aZJ1Vs1Tf7jZ+ejhZsXzuWk4M8UyQLm6G+L7H3
cmBrZ93T/JAM2DBMJJFaW/1H+4k1nSRhYs07tytX6+9vZLgiYQp95yfk3vcZNJOujZZcYn49pjuH
CT9D88zKT8PVyQqctSKo7Pw/wnyjabQyJP5zBkOgRrQj3lhC1vqQ2T+C4+9oPHEGGz6XQuBVdZ+q
cJpyZiEoL2HCpUKVjLbd2KBfMqnQydhPU+AH3f+6rfyJEV1+RftwMF3KPjYUHr6Qb3PhEJIuyx/P
IriaeCvIKdU60jp2CZFNaY8Ea0ZXoE52aU8Z6pOZcmyDjVbsLU1N+ogEg7On0rQW2c587HwiJBjx
DoFJNk9vuNCpijZ5HDWl7kNzVe5vyUk6BGN/w+tp1Ctj+Z9WUtB0SxLLkCngEnfd+SYH5xoAZ5zL
TzuxYeGr/N790t2S6jzACvdn4SGJHhVIqfzway3jBbo9D4As0NhLQARgIFJFxiYOWDlXC/RUrXIy
o5i14Qj6osUDw7744Wa4KhVJu7JamHdp6ONyOitXng5xkJtjvy1vuabGrVmICkYeuQALDMeTuGXI
M31mfYyA8GEcEoTkfRIRLZWncCVStwfA6aJ8D6sX3itf1dgYxjyfxION8Vt9WF15AUCvx2SeJMx2
+M/gTam1PloaXXUhuzyCC6vR/F7s5FxlqZByi2GC4Kmf8FWPi0ZP66I8aI+Ut2qXFLMuvUwAGWYN
iQl+iNQU6djYkhRv0bF1wP0Fl2I3SD2uxMOirGW4Ei8N5+9KD7qJiqC7uQLxnr3uTPAvI1koGUE+
fQ+dEQh+SvjAIh9Vhr4Ja/TQaJvt8c5ItmxEJv4r7SPZMFVWWL/FMoAQuOJRbSkS9gCODvf862P5
I9iC6G32vZqSiKhYTAApkWtlwexX+MUMhQjo+xULjoI/C67egXpmWRt1LZbqaZ+CRaIjq/ICDazL
TDL4U4Z8c7CPpEbG323EUlh0Wd/Hb0xXR+qJvHgFvjqRv69YtUBvldcquWamUJ71/FzxxFkNPHmj
clBsNrO58ZqHczpNrFa6trplZLleH/H1ADstR5v3X3+Hk5BbjGRQohgHmMSHsLfZxOXX4ttpBY8d
/OgmUh2YPFJS3jJ6taEaseXnwqfdZzANIJ8/R7Fql2miUPvqpu7605unD3LnIFRZWFnpELRnUafE
GVYw+oVadX9AuaFAcvmgCKCzxBALZsb4BgB8OITPYR3kyrCWg0RrgpJbisyMuwJZEUAQhLwKOaeD
ZFuRE0BVKWVMt/ecGBOfpKuEilF1d4uruslgCVCEAd11AZqs9iWOXTAQjyaEZk58F87iLA48aT7G
tC+qwSZCRV49W9NrVoeon4hq6cwyVzHBtZMFfaqWzR+f92K+Qr8AfbXPI4jJq4oADEcCIpPoulO8
2LfPH8qclp0HRMw2xr0qIdbiFcE19ylKb1WgUGLM+OLrJWCiarWZMyoalJAS50Bzj8e4c/XGs/+b
zCrX3nB23wTS1wdP238DLM8l5R+GalhSf7PoLEGOvdvy4Rzt41GtXTYtdKfDPvnDj7dOn0r0PwWg
XjzWGPmAzVbBJ6m6z+c8XaOOoPwdJ6C6SxmLoxUec7GlqRQe2QMveGi1L+0i6r/Vl2sIyfp42BnV
Vn3Mg3n16lor3mpsynH8ceKqGO66hfMzRc5WvJuV6ZseROHoNejBl6gl65LxBxioGYXkEBDVmiyg
Laa5jCunZFTx6v+lzZHYbMXkvJ+cQHNzFWQFgP9tMsrJo9xoONiZlrjUr2IjLLD/HuCnvpAnq4TZ
9H0fPtiHfkdyVtGS+l86NjUGy4L6VQSj7HTOEQUOYli5qi11EqTBIDPtMlFhG7fNd5OpZLJl2FTo
pA3610oKsdb0K344+0P7tqpe9d1AYff65gmgZ6MswV4Y4Eh0/KRElODwueLZgUKMCu/ZN8j3Ikhe
2p4pzGb8f41R+ey3h20Peqx4FdPmVdu4E0eVBGI+LWQ7DGSqTB5tR0RmSOym8vbjmkHGqUGHPeaF
77gC8s5IlO/IpW4g65Q7aBhLjg/2I4QnIq8vpWQ1idOHtrOwaVbOo8wOuXhxGQSpPtHxrNZW8uKS
A8IXmNRQCWC5EXkpsHcrCa1zvhC22tzuXRoiJxojqv5l/4c2mKPRxBYMFMDFoswugS+CtJq1CmGt
I/zvk1SR8MGucJhTiflZOee+aIQeOBcNm/Cmag8DGdoqV1ziBf4hT/KcEM+1iZCEDlyBaFZvJ2mi
irEszxB8W0q6WLZervOuNxPvRSNdnpoQRp/BYIhBXNHJYtXtRR6bS2nm299GVkFHb1Ni8+aFeqhX
PrdzhyKXgtj5mjDKqMTA5Y8jnpz6gpDae3PdGASJDp2kqI+HRewv3dKGn9Lqepve175qJ2+5l5ZQ
OK30JfcQjUbmrqRY3/fDWpbB5rJkRedkdc3rc6c7Yq5WiQGPdUym15NYkWAH5rloQ09+vgwgIVB0
dcEG5SdmnZ3WjcgyJj7lFrLaJjM1zmTrGQ5rGXArl+eEMQi4+9TpMNp2TGNevH0sF5RogDtmIwWQ
bUuBfRLjzjj1xw0jSTcrHw1zLYjFZKXmD8kQf66ZOtN+xWuuN7T9IutPtnrgMmRGNN7OADxc4Akf
5JjRlISrTPvRxG18Q6ZyTQAY2WkCzgd6o1k6HdR28qJxsqg5B3UWm7bkQ6YmqQr0CXRkd3mtMiG3
qohbthacgKltQhAz9+dAh4i/R/XqfvOf892ZVQVc+5KUURT0kxY34WbKpXOFhDTk12e+3Dy3akg4
ubo7X5c6t5Kz6xQiMwMBNVl/NUs7KDnMuULvaY3D18LYu559uRTUMnvTSnPvu7lG2BDVepfUsbXO
Uwhhy5FNDhlewvI/dc1TB7tJrWEs0nPtU7FuSCj60RWnPbNhakpegSEBhAcSlftjSTisMzA4C30p
DTXG6kCOLTb4ct6wTVzPEetC6fuMSZZX+msgqi6j9CgskZnsXR2pKjKDe90ytU5wLbz2mAtjEyKU
mTVD3771Bu3RQmbdt6hdb9gVg7/B8zB72toX9dru/czD7P0JRjGwYul+Qm3v/67b5qoHINKHgpaW
H6d6+BojjvjPLB0sl242MVvARPXOMyslfE3fixjgSDI3P5xKmUfdHoPId+T9AMrxgRPl2PxONvLx
cfm8PWDp0howrpbB4/+5tKHCeoUgAxh+7HQ+cWp3JldoxWu+t9iWDUdiVhw/5Kd/VmRi0+ZMYD+8
V6RHet3k1tW/+VTgfuzwv8ojAOYJv3uBGhNAqPh2YOMYlkjwMkYh/aJeB2wHyaFIYeGbqk20wHcI
zL3DjZbm976183cdnuMz3IETQSUw7TEMrrroZL2Nbyuy7+9sco/xeFo7LKBImCRMiTUBLjZCyzSV
72/mgIIFEaYjTJ15XBV6y7T8ACyEOj4sGaIvWYXRidCXI4OogTUj4QlSyYEs5tDYp4rXElc6pvyN
G1ad2rPYUwrBHcgEf1iJasibbDARjjq9iXFweNX6dSnRGtzKOQ9F7CEERyYJhK3ockEbv9KJ7RN1
iP4vypWjbAOkSloFpFujCVtQoj8y1O+F+X4CgkLISa64Y8CDk+igh+gZFiowS8+rHjlH0SaRK2kG
FLW91d4Ne7DIWcYFrUbjAXfRlVQFikfGGZ0Rub/R/0OUOMPO6dICOizKrOl4a/rWm4bSrMcxjYiy
bzDzlQE0Dn8XEG5IbsGw74VsK3kw/9gmelZkql/NVw9OuoDU47AWIGXph4I/PjW1em3eDT72YRAR
yy4qmGkhNfJ6heG2QldHOyWUK9xuBWTDNlVQezLNmdiG5CvwcZwWTx6Z0yUYoqH+QlWxvW0HjY1R
NW+SAZYlPBRaj2xycKwRWINIxK8KeXbcl8ccY8LeY+Nxez5mL6rf3dYZYGBMNm3cWFblVZw+qSRt
Jhd9AMd6XnT0ydr+KM+78iw0Yk31Qw3laDsV/y+w/vxJ7/PDzN1nb2D4TGDW6i0rb/mu5T/nOYfT
w8OgGWohTKAE1R97rWOLnJ4wRRDUayk1Z9LMv3sX+NidgCA0NXZzhhVYh+VHXycjEGXTXMaYPjeF
9c2I4rkpk6aZpKcXhAUcWRlPNjhlrI1DXBewb8HEA4TzaD3RpKTbJwWSMWUezWjk4wC69AqF/+B4
mIZqHRNsMjamsf/pDexpR332mT4JhnSp4I97zBD8W6U4iXyv/K8LNlROBLQKzznTL8yEooXXFM+D
BITcVjuqUIyAHWsb417oGWKsho1x1PJsxkJuNSl1ZSOKZueIoQ7vLwpXemk9Mw+PDSqlRvUDrkou
uhF/C5d20Q1gPIljEa/pjpn/TNOvVvsdL1s5DWbxoANNsVamiypu44onxeZG2nva3LGlXyiO6WQT
wupH346kXkvcRwt6eykIByFAvNIZpymQ1vFEeroaUnJ0wBbbj1LjsJJDhgWJoSoQ/P4aJMoY10VX
lQ3r3g2nceZCZY2saHLQWzY6A6yrlFqNg+bG5YH9o6Nye+f9DlMXe8YKwTpzivxS5E8ydST99WKZ
LmxVkvV33kYQQv+rnINr2pnW0s0k4ziQLlVgVBi0PpWzhUmnCKuRilvA7NLZkIbTVF4USXeQknTQ
4Ggc6MGy3PQiA2ilLp7yelhvpZf//2yLoJEeMvbyxEvC0DYOnBofIIPT0865989mNRPpgMgbvgf/
miKMfkvlNdHCJy2SS6QNurCz+j7DT7HZs7Mwaa1GvXvVZpBwa+c0biyCTS90acYkzRVH61deaHFb
X/ypbeLlZ0QkBkt33pvxHn8FXwfokh6K0lCGccL/yJyiElNw1niXw3cMeLbLXNyUQh0NaIKfVfdR
5VfzTu6bKdzDgRMQRKiadnsYIPUzBQ6mxF0PDSwvrzsvW3j90wiUNB9f1JvRcuLziNa/LRHJPXYU
AHG2tOMpqWFcR2csOigKCW1PmHA5da4VcW9kh2tZTz2NSL4AyrEKqlPkMe0c7JcicjDPe8a1I0Yz
F/FLuXMD82RwBjeKLUt8fJ1zrbBsBhqqs2mRtWgiOfq2dDam0UOwPEVgoVb/1C/xN5y2y8yMWQgM
klUdMlRQ6/1NcPM8NPre/1riauEwpNJ4ztox36TKbgRTy89bga6p94jm3sk1nyd6nmbUTCdkUL6P
+5Nztg9cslc6VUMdadmi2krPtXu2pyobsKS9qnk9HPq987RjKzyd7QeT+S0ezHQ0sPpLKTXwNxtw
Wlei4QKSUceaN4ckD5QeSXw+2Q821WYQxHheXp4OYqeZakzmemlTIzukyhrODcyrUTZ3VQX/ZoJ5
mgwmOwcLobQ0qDE41uEBBYkK9OQKQJa32Cw+HrqHhoHmbodcTwhnKYlUAhS0AQKkf9uWuu9V3SHw
bWhGd7mCingz+1mwwx20OkTaCe0Ny6mbp7cwff4I/68TQBFz+Z/ZvcieBHQzBkFDavzt4fhowTDg
WQCXxbnJrZHdnY+HoRNShziPY+igZkUwC3KxnvYckWawN5gabinhKm/AFsWZ2AAM7aYLvLSK5pVn
j3GclT/94sBOWxvDpx+XLnjTp6ehtt29Q+vv9RkKF5ddACWscmT61krbR1c+M+QvGUOblZ4eQsnc
OWG8IJEYaEh76fyXho7hLQZ9t6F9xzAi1YkuoJ4IR7vIiusP86KDI+v6mnl0wk7P/4XtC7eI0Yes
2RZSkzpgr3SoNWNLtStrcCFSZ8gYr7ZPJmRoFztfjVbg/pk2+F1Ub03qP1Bw0koqfkku4/16GxuK
3fE6EiVq67oIUu5OjJNyAybULl37NaAeo3Wx7C+0m2SReTKiFeDK7OJQ26OszCjnLjWdWPg51w2A
5pPVp5UAcx5tIKN4wCnbXO87gKF9l4kKVhS8b3SS94VcGMmtej0p5CP0J+psABHu7Kuy4aJ7NXzA
fivPfj7h+EJOmTHXlL75mdQOI9YL9aFxSkgRlqeekSHaGDKLjMe3nFOggTZCQGXIjgtYkI5HxJYj
RorJiBk7YkzE8dSx9weUdbJ4hsdrdzdna7z63bGx1K7HB5OdrDS/9hWG0mb/Ftjru5ApPVxg1g3F
b61u3e3ytWBb6kI2ozBMuoHmK36I6SUhep+yTw3QJTI2WosUbhy81yWueJceWZww4dQSsPUccq3n
9BP9qvqut5zBCdhn1bAQ17B4CQdfwe2MPHdSbktXhsP+ZlPuAl/fzmp1k7o9iuhF58IgFfnPXuv1
wka7JQpQn8mRCk+xFnTTAelbEnsxiegRMRp7Jq8qBlRkoboGvDOX13fStt0HK9XYqUmGeP732uQk
fL2MhLtA/fgOUr8VtRPYyngcWOI/Pq5BFvv/W1hgyTQucFJTovB/tHTNNUMFZfekkcuA0YgZ8ZD+
+Zu51Jw1c6FjAUEmosHgCO9BhD586CGhC9U202JrDgABe/B4mRagon+OogUIkQar5Nt3pvdY4ZqZ
7rEi9hNPvK+N/6rVbo+B57gN5stH/8U+POaHwjo5nG3Tad32i+zg+JAfHBUnLGx2AmzcqyN73r0s
ovbP4oj3PJ2ujVbBV7miTqL1Qrb/hs3JZpho0c76YDswccKantIFNFnMRP13FEqrcV5LBlPwKhqn
KZmntliy5SJOTog9ObjWY2rfIqmSJIk2V4icFqBW7puGKOCykxn2nkDLfqA9psUyTo8W/wFxUO6+
ZHTcl6gPjuIVETcsIROuKUX67R+oqHQjxNaWmCeV9NW32239qBpKL52MjCnJvULurXr9XlDc1IBd
JO7AwTYveMrNRPy9ZjxbHmTDOfxL3L9oi9ek/5LEKV5j+hLoKNgbpB/3Eq4S3AhtkU5cmfeCmNIf
mnpS3g34v2WZCvFxdbX5TiLlMNtUU0H6FsWT7Smk1anHeFPqu80wWsXoJ/jtumS0hR+oKPidH1H2
Yqr47vNwG1fgm/qEnL4qi9DwRcNjzN6jZ3rDmTnjppK2tp5DgPLgJbn/KFa3sXAxjz/QELrh0o7p
u2fxoC8g6QkXrDY9lXTm4YM0pMZuJV2OUIvHaFek5cGJiiCM6c4AOHv7Eo0lg8/wU+HZNo7DE5Dv
aJ/jeXYhXzdpT6P5Mmu3TYBy7f7sDYdQPdftiVvxiEHnW4V1+xUJ/KeC3eFyhlUj5dT3JbaN+C1z
iu5Jv5VScSnWCxh2b034GDNJPwiCg9e3cW/OwbIuSNPEfd8cZO58PcAbgYF3Cm9CsfA8bVpiDrGt
4fFw48jIQPnG9d/W1Uwk7AwCVgpYstnCg7EvMuem7uHxO0gTBdFWA/KhojS4OO4bdc+aFzRsSTY/
TpZgzWiiXiPKwOp8WHD7DItxApxsA4V1w+s4R9mK9EPdiJ90Ybvxq6Ofw05aN/2HhGVIbJq7ZTO7
hnPpVFoWeG+iyEMp60EVH0s56pN5aTAv/1C3g0q+vLwfx16FvyWIjD2Iamka20nuAq6D2ctEnfWf
Gr7B29D8KNbOoWXBk+gTgYcAjMyTuIY/+1gbs9m7xDg4vAhkQu8ikbs4Q1BbGv34L3LjobfsuFRA
xsaAbg9eEiJsIeitfobkUKwDe2N5XSCW8I6OAdYIfVrA+Nbvh4M+MAoS2vhW6UugFu9tiDySt0ws
7ppGwfTjZ6UHBuammuGZRufDDDk5Z1C4TNv/rBTaLTa5YjIF5LYV5yCDI6is3SGfEE72eABUX+Fp
m/GTuKuXleXe5MscGWMtQfA0O7PGuQOurQPlH+akwD/wKYOrEN960iycnej0HZgMMfp7DUC4OgZl
PcGkXF3opxPqYmqtHFRc4b8Zc1mjswKCV8GlsqEIMxr1t7SIpMj1O0p8YOKv722Hd0QRHjYne1JE
SfL8bWBUkzTow0f1a1mj1GMMMLvOUDo3ahOc6+qWGOUx1NN2mWvxMazo2+v1sNpaXZnI9mW32TbX
fJwzRRm5QI+O0uPsL2g466pMQBjzYu0HumYeTFSURl9qjr7CRI/XWGQde/1nCkQJoa3mTdeW+V/+
lX5iMBA21jOJmIzSGmZn+6e+++O9IwJs+LVap50H+dJtUhJCVdOmp626NFB9rxc229LDoWzFSA+C
e02+06G6lwuy3vp3bislFUr6AYbu4TOf97/Ul8kVZXeHrWWH3ECVhFOPMP2kfz60N90gB9b02Tlu
TckvDA4TctKeZGSzn/eJp4/lchhJPSw2oyphN7iah84KtEeA6ftKH+ohIS5hg2XaN/zpZMJ+6SE+
6llDms65L2DhnMoS7xw+oi49PXImGvOVD47qYGEr5Rf/nUOlsEANj8k4B/9UNJf6UB7/siqejhGV
GOinrCz18bOe61BgwK5O8D/se53g2DYXXrI0ikQvd6K1+u9pgbiKqjvpxjK8Ti737C3sEg3zGoCv
awAqsPKPsOQe+O7herjQ1VRg+PEvXMtSPXoVlB8QYDn90FXqz4+LMJKj4tNLcksZ5/zy3991DTi2
Si5bWmDW0v4aaCVyuLL8kEG+uZ19983yYZuY7d77TBOo3WlZbuzuTHLQmeUq0L48ZGrQnxMFqKeg
dvZucxLMObV56jwyYzQzHBK9SZAD3xvSE6xe1dZZfDtbgwOd9e/wwimUOQbPXH4CBXZASZDeCtKp
slqTnQF3XOemWmWW8ATQRH2yvtahWAbU5S/grSsT57GTmwHmcTa5LfAuE4cm/atKHut/J7SFt1Rs
NkiWKQmfXzhmnV9Sf+Z9QYzYiOOF3/k9FugNmpgTtwUAaxObbYybHnRBm2JERfQF/9rVzLTnEBqg
YjmVaafEjuut90hFE1Q+U63q1TJ9X1pJPWEquSKJzcUp9CRqiCsdNhMljqcM7UPwjCIW6WABRYv5
PmDdjdwcvEckyF8I5E/plqmyesz+pjSdi8M4xkEAW470Fz4xn+vCKk1pZBMHqYkTDsmYNZPpJLb/
fC5vu5dXVgnrAPKVxKTrzGZ2YmnQjTkZXmmVSLbGGGVRbumYwQilzMN8I41gGFW9jm9pdmbG/Drw
tSxk70JYgSQu1GB5RuMKhFlZkCw62lPcgXqHZx8BzXH8LUrC/cIdjBMG2iJ8pQylGKYCOIgzBBkZ
3QcK/UmOcKVLiNXYf5F22SIAsbYQzuGCvLbIbcswFOa2CBDV+9o5+ImCU1NDUuPF4lMvxNi1gg1z
GBaN5Xv9O79SwR4wmQh6aMxdEi2kxOurvfrpssKtJKqtIn5+qAhgNzS5HymoResSm8w1iNBmo9Op
3SevwqlRzZw3GuZZQAtVfCdkCtVPgS73gbMs1/arMQgfp22Hna9aSCmBfi1FCkB3B+LH/VQIvb7N
Uj4tYtHAaUOHvsEcrsaTrFTKlTkpLH5RhRhoiYlsywN1mpsJTqXNsFbAeTHEmQfemd3yXIzE/FOI
DpznRdV8bua4SheW3hBd0f3jD0kkTKeTMRM43Oi4MPc34LgepvV97Pd3DLqNAJ/uDNQqY6UpaKlV
Zc99ESEXhNqZELOEVtdU91v3ITBBc1PwBWxsVLm04nDvix+7M/XzuBJNAeV1x7bsUE/0cDWbEAmO
dk+8qHeWATm3pme8qLzWx86qUKPOu2qePH0Mdd+rrD6Gq77byCc2vcNL9bRpOFKHRdTovyeToq1n
mWcGv44uXRj5INdp8Pm1i8vgy62ZBf5jUXAN23wGI0aQ2FTwiOk3/gHLTSTSlmFMoJiUdNy1w0yZ
JEfw7YahLm1HfRPNWwJ1aDUIEOlIcGOtCmy8uWMmmOLyKCmTEIksUT5m38vFSSGoy2+S9t8WzSid
2LsCse1g6P4LFdd0yKL0E1k0ot0qyCyZcTmHNlPnozaJSXImAvm7DBl4e/cxe2AXkLTQEoc8zgzX
7nXGiENDJAROM0QJCfq8SW71mu1hngEqHK0MO8xfL/a3Pes1EDgPVtbFnJZgBxyANFAHQyZ/pzUy
1xaCTy2bdchhFD8YGewZoGB5xx8SdkIl2GbAga9LA0gJP3NY/1Pp7ok0/G6H4v9egDHUzELRhMJa
fYC768CINZV1wcnynJEssNmGY/xlAc1wVIAwVns/Z6PETvuOTTWU8m1FLsLtX9YaW96MuRDvOf+E
GqjPC/Zq8wgX7kC1BbRyveTvC4fJkm/m12lZ8vC1isrML/MAB/nsplLYS99ZjtJV34d2anwo+N9E
Co2TE8RYRIp9SaGhxKD/2/sHo1p6KX96wPC+YfB32NTBUMzUqdVZjs64Vojf5EOxxDfKSmHzjcYn
ed5U2nrNvBr0OypScfCBjoP70g02o9kGWv0jarTt6cBiIaJ7CAzJrXmhr0Vh+3fILQ3AhwgDArPa
Ds9ImUSryzwSIPOQ7bCy2acIkd44AqXH7UtT0Zn85L6fwcxOYTbBhj+OrpXTr07lREnOwUo37zBF
hVzTbOTK1HtUn2q1kzKVFOZXHYPTEeMKNQUJmvpzW9pzon+zI84PiUd+Q2wj9CCFSHVOz65u7ATD
QQ7fmBPWyfQYYOViPZE65L94pIufT+SqE6eZ5PHDO7f0xk4KdEWVd5nv7JkPf+oidwsSxwLJxD4a
T/MjnMt0V+zPTibNHhpJQRSBvCTUqbJ4TtY53o7PIv3Z1Wq/R/KGI2QcXs7NCZBOoduMADhBB5en
zVdcl6DTvH3touKpau9HhlqackFwmgImnHFabcfJiYUO+Hd8VYoEYEAg9sEXddyQUmiI2LGd/5MM
PR8dq8wA7TlxOCGhZo5bDRQ3cO8C7iZYjIgigeD8XK7zDXALcPiPMCsqdxiYdXoB0SIQWah/0vp/
7WFj4G+bxHEpoyjqR8WIOfmIRWnovph3426MV1lHOhZLWoqRqwIUetk6Lmo0QxJ9xnervyw0SN3K
nex2AUZ9CvXad/+5e5BcIQbkxmW3fDeaCstlhfC9f7yR57iQGO/yBrpBHcHxI+GB2vXWXjlqypeO
9hg2wmWOAaBCBjBdE6m9iqRSK0u5v1JwnF6sCqv8TBl2Lg5xB+sqnreseeWgenLKtxxgpAyeESVv
nSI7uucZzUM0XjXMr0g0YaXiKgiypWjP2qULwrZaMmTUGmsa3JQxsVqRNtLIu7CwWdjpF/sWzDR1
1DtUj3mMFLFdJhmra3YTI5jh/4BcwqjDGWRv+BUCZ3B1W7mBd7jdLzpPRdESSlaw05+Ue1LhEuXs
S27imYFQNFDFiH6nklvqBuPeoW3auYgenh1lUrxXMaXNcJ83fSb5AK3Quocoss8l2J+KKo2XNnQB
kDN2geHpL0jFt6D9V2Vem6A3LDGNX520HRETCEpHu6e7Mp9FNaKpHm992AWHW6sZbmpm8JfPFZRc
i2w+8qh7NVTukjSi6PEm5WGHS2DajV4TcBy0MpYBe6dZFmXvUcZussdP07R7L865XJt1MRk+z/F0
fWmqiUG+jY/cHb8djxQ25T+xWmD4ilvIwWhFcHiliA7sUoDPBDxMlhTEpg6RTB9RVVNl6/8BgCA0
ZzV/U3SASYA5uGg5yml1NBDomZr1mry4IiBOdnmqwPfdSfKqhfFJb8i3P+41wakcbZjLPsJudzpG
0Apt/EIpwDVZgKnEd1JftzSkIlvAAg+sdVXOgaoUIO20Rvg11cjt+h20Mmmn14mF0ftw1rFwIb96
YqBawA8M5sW6w72UlUsPqeifOXYkqubtBQeYV94UInKWmZgzdocCjF8XK9x0cJHg8M077DO4KYy0
Y432CVqxtAXxXoiMde/SYaFweT/YUCl3RuIFM/4iGD2eW4dHwPOYiijUhMtflWbJaWJzyKS1D5FW
oBqZJN50Kj6BmK4iN3rGbb3HoPUUlwrn9H7SoZ6H+3IHRKHhuIWyvWdGP9fOWcIFFRPRblOIgZdL
z85E7Yr17gmEAMeTGQ+56Lum4WulZqDKoES84kqsGiEr7wcN48i5xtVGwf5ee/Dm9s8MMib8o/L5
epUQ3exSLysCkXH73t2yWYFhLO30XR0E2R/5HgVeXKQwqa0mjhuwNNeeQLinRMXG07gvyz4YIM0V
VbF0UV9BvSxAEWUjqbU3UK67iE0xe6djeorwUY70rdFPgXOskj/J8efpP6bM2AjPigIWr572GJaK
qs4DJLL53Oigv53wgUVLGLLZKs1ywXg1LnwqxbSTrHqgQtlTzWa7S5t5FQ81nfal8MP8sG3vcu44
UWbitkCOTBRi7SczHXU6gGEjoBg0VtJRHKTFxBbv5gucHy++H4kA/qrwbBf3FT2uO6Mfn4YwfDUQ
QFJkgCsNzotyH3770cWWcTF+d3JAYFh89+3j2n+zr3wK4urORsdSRsJv9fXSABJ5gRLcgpgjjP7z
PEWdZcE12Z7ubX1Fpa9a8DNSmmqQvL8m0+rRmsui3emOk4zF5thfNH6SYKi3YfaDoT0IH1TaTMY0
RT5nzefCWnoUIgk86V2M0GSytFpt+S0NKF76lBKRPo+5E3S3ST38kQQJHSCLRWO60YLsyG50xrF2
BOiimTChDj3WOM9aKNWsK0IYy2KgFPjDQd357sIO/bYvr1SfOyJJ0ncaLQeidz+00FbjeujcBMG2
N52gBzlTIrdpQI4F3laNQusSWQ+4nxqzmAoOmKE9OiEOlrW3zWKKSgV/Bjki6SKGQ9kwrSS6KqWV
D/AlHQNBEHf/vutd7UqVCz4rTtmm4v5KG6vg3xPgqGwgdck/xSJQRYCRgQ7Oh+CyJQ0F5htvLclz
ruBqTtbFg38wqqf7Wv2xuOr3RMKggVvFNZ2M7p06SgMgKMNtyeygzEVLaHWBs1ISye0cig1tXCny
AtNRZUXCYtU787CcWmUjUBjapofm1rwKWazYzm4/RUQoMVE5ygdEGL+S63tERuvIVzrtAFxJ6OxD
JztT8PkC2CbHQwetmfECMt80AQKtk1whTwthn+85vp6FtixUeQU9K6mWm70MqpLzaYjnsw+nehda
Sezq9KYqZXVd46nQPLYhtO0D1i9azX0c4g1oz+4Ae3IOJy8WBhcnYlmR361SeR3YKVumd9CH4fDN
3ZVf9eYSp03pEA+lDsSFNwDg3BaxUah1g1RRxiIffwDHkDiSCsSj6p3A2SsIzzOD7lTmqiJcgvOn
45UO0DJu/xDCXmULhCRv2/HjDdLI4SQ7h+RfljdTo0pcivMm6VeXbZlOh12XqO4Jm98OWJYqXOLd
jztefOWdDP76UjcApD0PHIP9U8BtA6damI5j9E4KPxIWqJxtG/5/Vbe9BI5ZZNoDZS2Qm3k6pEVP
THLsvXXX6OmOQ05e3UWt6G7rmbhupmwpo4/DbkXWn38sm7mBO02rJT/RhvdzAyoSczqNPMzHOmPo
DMviCcUSUY2qxp0t6kC8USVb6Uu2BinhNTW3FuAwXObWtUy2tbGtnHUOLWdo2PP36X7iCc5NIP5F
o3EpJyyAs1lXPPk5zPrIVIwRBDZWwyAt5QlzLDJ2UZfz8RGjGrT063GEEVAcdcxVJinpT+OASDvw
UZK9FjadkNFhRh+wiiMFbaSxPRP4zaLE9J7v/EvY0eF78YcmlxcjkbH9yL2rTeEeUifLLrF/IeGU
u2fc3Ijpwy54idIESlO4UOwbzOhHZnm5HWPDw/51oPQrOUJzKhvG/6i3bp6mMYzPaKJIhOdBIhyx
5LBU4TkIx80jHcy6A9a+Lk2EfaQI9yQHdBq6xq4j3r78TRr36FX6tO0vvDS2/omfAaKOLyTCd6le
DXkuCOl9OQzz/wxP6JixB5WKEDVUTT41AxTNkath8AF+/L08zXazk/392pYg6ahDHqQMwHfxz6UN
ydUNceQeET6c+Dn+fmzPwqAvNH1yD4xnIQ4Y+kwutpVBkNhN56Lr3iWUG4kYH74O0lS3ZiE6bc6/
x4TcAnAm+2aB8TvClPlqivEqT97lj2jviU/SzD7LnrW7LG5wkgu4RBIqhhvaNNQTjHl/bkvfyfHH
K1yzd/RHbeFqu1hmi0LFYl3DeGAiwT6gk6NPKI5Z4hWYRWqrUwg0oEAnwNDuhrs6TQFT1kgIg7ZG
8dfWG6AReq46OKvxW1Tt/9Gh7MLymV/53lQx+D1r+3XXT6gwHldIsnLKJb+m+FdKg7am0Qq7OZtr
xtIIgBEnPHtSJC7mZnaQiTlE6/45qd7bq/TKFqPArx1SBn2AcXpVgljb8vnEndLyuyybEEYkup8s
LcTYaqk1JDsH0fqRBTKqnJpiG4+1UgtGY6EbNgTFiIBPb2qp5lTBVvrCOpDgm5OB5poM6XuvwSc0
JFkQhDi1YeXbz/kAgPqG0cRkX8zJoqwVEMmjbIfzy+xarEM0EH8lQ+s30oCsZ3tdzobpuSd5y1dJ
16dGOqm7Ohxmt3OhC2znwEXQNJv3KD5kBgHlf8QCpkoStCfWlOdxaNpQYASzlf9ymH3ILGmghbHJ
QKJFegNUNf3oxsztkTmLpPCwEH2V5oz38ASW2FUWcwq9GYou3DnoaFxRPjvgFAEsknROxlFzgI/0
OLVlFXMQq9/RyYze9nfNK6eCMPLAktfdvqB+PcJb+S8QmwULQn+MPv+lfju16XrTdADOkD9e28XN
hdncbOQebYndRoRqVjq0D//S1c2vH6snOfw8jSSF4geMy3IVdl1iV2/soWFObulI70/tRuPKd9Kd
IM7AFkRAxdaqfjvKPFvNF3IwgqDO/JLOZEgaDhPRgCO8i1XkqdQYFzkuCfKV6g1RaW6I2gIy3kd8
4BoQ1C8IVzL+yrRA5b9gxeLdEdHGZnjnzUr5GzUHMwXGngVEA+Qj55fCc6h+Qns/9Jc9uAOUybeK
YeVTrglC0lLtsmHrSOEoYEcBFb1YaHA3GoqqyetKR323QumO1HOVkhLbCxTS8oS+zEoAcCf+OjPI
F+4hU40sVwwvkjREW8qksamiutQtXLLv2OPm1tDr6D9L1KMW9Ks2KTaVxV8ZfYJZXzaMuZqZ5VI7
/CsAp1y/zSRmd0OG10En5akdxCsbKGjXOIW3rzxlga+IUj8UoglvuCH9hFLYxJbVpckW+ebliXfc
0dCeqRziPVcFSugeuBBG7RuUwRWYFZOCHlZPXxXW2mHOWMWiFFQxywIKIlbJCuqOG07yD+iBv6uM
7ZX06UzadDTLyfkCjGlp5ZQTmIlN4SVKdwdFP9ULoJCpOlJfeOT0IqdmL0mOetoLLEGbM2cs0oVq
xsWmo0TZ7ELUHHaXrDvynGM6e4P5IfslfMKrIM/xK6ERXNrMbkpRY1XDx/X3W7t3tBDW9TOhgc6o
kQJqHNdfGWWWLtWEjkjVU7NVrFpZzLZcYb9WuL7UuAS7yuebgI5U1Jcd2sOcmkSWcfAUICXKZjKt
5g5mkFXkjQinPBL296hVN2j2zrQlYQQOqX0Fm+6Ah7oXKQdeNXDOV7VoL0xg7SidY1lhMZYZPsUe
M1ckla/pzfy/BxgAZCgw9MxbO/iOtgchcmFyP6UT3qiXrKB7yECp5CmCMd04p1Ulx5/nUb6PbM2R
aagdhCfhJOTBqNvsGXotPtuFbvytE07hIenbAQVFYVRcZNbobiGROuFilkPuTbaaImFWOTNO895K
HzXFeIMlrAWD3kxoirLumA3/I/8T9sHsBFuiV42s3Nv28rpMYquN+9vNznfveJcuPviNLOzaHhK8
CKIMnUIltbTYV7AdHyl7YEOVKsZhjVqMPtadHVLRVnVWKVr6SXDzc72PXBcGJHdOr9YjuXptPY4t
9u1wRq50mFiUMYnipqjMEqGCuhiJ86egWIW65jJwVqvLcxBv6PZviJWcUK/K2hhsaiMs0RHZtZ9r
EwaO47xqyS4zAVBGX/f1hIwtiGKejVG+xiZ0Av/VyxL6qYMyToAcgceTAlgmxMr2OYLjMRPrqzTx
xFRid+o163Cc3uffU5FT5l2e4tAQDIHf3qd1DH3SRd86rT8poFyqXU9ZfKAr244IrkidbGHLzaEx
rYkac3YthIP9PoHgcrmjaKYTcYvdkMxGTw9jruWGw3oDr7y+y6c0kFw6arzylDZrGa/SUJE/qP27
r68wx6/NPIIwxX4WxeYbwPJ3Hm4QN1fGxcyx1LE97SZuqx8i8GvzeVXUjAzpcYMda3W3xzclZ+eJ
Xl+acDAfJtqXnltDhwCLv7dSrYvvGJD1x1REajMM+OPNOvSMZ0sn0A1Vxplo2YrvsRkZFvOdrHS+
nyWDqQHTCVexr7nnk7EAyBPf+POtq1Qo7+3x34yOCZJojGtkuElUUSRncSo7QJW2NhfWF5MUFd1L
H44kaZStJ0Fd6vkuEhHs1vj3FBaXDTwJne6gw/x9RUyqs3rAX/23Ave+QCLkFG2zXTUvGioOYQfO
QOr0crud1Z3qDCCWM6ObGlB4msg3j1nLOefzG9ucIZsnpp0/53Uuipc70M6/K5DmNy2RiT4g0vHa
J5jBjqLPdPoeD4mP7dxib6lHGLCDHefAdPBnNCCvW3t42GD2nEtPQCyvwjTopMVT5QKCZPmBpJs6
6JgXleVk7udpH2R0KeYtp3mF4RIzXzlmt07zgGZigPdwmWhpZdK1enzJtqSPGZvEmsZ67+JSWLde
j8oPb3IYCjfmzymIFEDRSV1PMCTeCFMmmtTCHVIrqa5LO/eMZtarB7gWv44kU0Swtq07U8aRe/bA
i7/MvvlALZFpIAGpKjneue2t1TyI1C98yl62pc0VPxOKs1rb+2SezkXIfF/ObOcv2HlODn7HM46v
5jTWJqwSWyeqWQU/KT6xKicZNMSV/zgZ1+68uLJP222hMqTZ4dZcfLhEGuKcs14UNkyCAiX9/Nmm
DAktp79L11LToVuwM4KSdwdklZrhMrJJXQVNXb9QCmNdZ+nip8ifi3Lk0Wff5cu+TLvtXoGeLDjl
J6GKGMcnT69UUaAF+nm15KXrH6sY1kBqhfRLoWPYBSwfpdY5WBJS6O5LmqEXQ2szy7AbA+PCgOHA
a3dcsA6hqerqpCHq/nHsR2M2AWEPbU6uygKFRNaDfz7Tvb9woAf6Fdcq2p+hjQbim7V3lACB0oLZ
NDkgfYPFUojnlQddvlwJ6xpzlLGECakGU7PR32sPHTlbdrLR4BdK9HXrzivxW0H10MytbSxJxG2Y
SCFK1U4i9EZxvfoF4a+8SOb8IeUIq1kDnWrUQT3qQ3Lb4ueQaLca6YJ0Fq+Efc7xHjACpn14cwqI
rkJfiLDSQNgFiuYRI1MI/7xmue+RTHJ9a/Wzo+3rD2mszkbbOhOexXhubdzZ8u7qB/RmnglQ1gfo
fAYGzybKYzOOchhfi+ZL0D+/Uqz+g58c8RsPxIZto0xHILgWQ8FXHVj9EdlQJpTCoR8EJFapiXfL
2Jujsd2Nn9oMRSNQ+yU6hxTc4PJIYcuzmi3BfC7pz0O3XtHOjRJ8AzLfmKj7wE8WvpGkrC1eql5W
20BeA0RP8sjhPh0iWdaJ7C1ekzQ8W3F7ke0kWpE1QMv6MXwcq0SuWi4GyrmhlWyO5xhH1EgF9AWU
moiGWrnwR4nWDnmFIWQuZQkP/KJnoXeVdGu6Y1gKe9NWYK5gmb60eC+5d2GhdVUX5J+6yo92PpDd
aWyJz5HmbIn8EJK0tvX0r41IjnM559qck6qD293iRkH2aHxk6S1LrRFgKpBnFqaOWmg5pw3r+vCU
VIMi0hFLrnSXlioP82kMd7iG93EXo9a1fPycIFNLhzqsPagkh8rulVZB3C+4+s4ooGnp9bVwNVWX
lE7gN7BFfTsSZ+PtdZXq6pJi2kTtwdjygNrdTDZBM4/Sf7C9quGdNfe6wV9rQ9GieTqkxt8hPZOy
UrxIUz8NDNchLTDQRakzkLHV7WBIYk+r1t+0EzdC+tylNxpmCUI/HEE4N2soHkEBP8G2n/nzStDu
qb5Gh/SLYwgD/+XNpdd+OCQ2SGvoSH0LJsfnmtdMO5fZ26HIgXaIz7GXGGy0SAO2LyoqcX0HFtKq
LgJ7d3WxD7IcV3M63AuMSjrZ0/oH8FkOXtYQy/I1HW/tiUlkq8EWaw4fVGJmuzK4ylW4at96ouHQ
IKo5OcRYUrXF3LHKTOOA6Aav1C1od0ZvLQE6fYlu2QuNdsdEpWCjZilXCEoKX52QEJYlM/Ap3TlA
Dsu/ZxwFzvXhb+wnQR1k5y9EOhH4E2eeAULsZckZkBCCDujve7Xkzq7qt8ElhmSRKQaoFGnaCjnl
JVq0HlE9WwqKZNpdNbaFqzjqY9g2BLbRwxAeriHPVY3hoafCUBQlQejJ3oj8aji3Fe8/U81rKydT
SskFZbtIPexRrlPbMHzwFALxHS/jdWm5HV6cUAoP3DEYas6aW9qwHJgz7n30VAbImem5iv6u81GS
1v6fUMMZLb5jR81YIq2+4Fwty8KdjOo1jg0Oapvbgo5ox7+Htw3LYTe6G/n+59x+Mem/BFc0s37V
R/wBAsSrbzXOddOWFKlgRbZw0jTpoRsXM++BGQmsvByezOvqvcXra8gBcCO+iy+oHSO7hnmENfql
aWVFgnEhRMp+uUcC+Il2cOGkFvVAqh5ZnB1IlEjHAEJjtjAlj2FP+EiyVeObqOgM27pXIRd/1hrd
fB39a68V7NKqahkau+Zk3I+uUgCiabx+ewqfXUNpHlJ8UZ1+4TC5Je29PT2fufy2taihKuWs5DB1
RZr4vKb+eE4KO94g9bqjOQmDPaCcZXfCXNuvslO+elYKsLPFGCN1Q9ymSV6KGqbsGdt+wjz4oJ9m
lVY8wqhr5ZQ6sm0sze3UGC+z2pl3noZApr9ND2MsuY+p78l2wJEdvUdUz7UTnyyDK9bn4/sVTH8R
gHq5IvaiRcRnOCMHX84VXsdmNBxWbaEDNGaQ1SQm4Etv/ONPE6SuwUgZmBCqTGgBClZOX3Ad+aLh
gUGuZWKfcVPfKglz59Imb7FlbZ22w0XUmjRFFLyXbc3Vi7RGwEA3mGwhxN/CO+UHuQeUU8JyaAjj
1GkuNzg7JnIm1411ulaAuhsEXUFNpCJMTcs4nelBXnnxkDlLyN+UPz6vc8HYZOirSHGul0fC4aJC
+QaQSZpBVvNPNP9Vp0MR+BC71/vvAKpaB8Lg3YoGmbn7Qxe+hDRA8dz8eqNunaMvul10/A/EKeAb
ozuIQVJ+awhkUhS7mTgYPq20pL350CycjwH8/MhhKZNQP6Hi2AmOUKjr87G3wGmHF5NyaPvkvjJ4
Bc2DWpDII1PW2fzIUf9SHTpVaeTaTWU0aHWjBbAdAbJP13Bx/loiowmeOYBsCK3m8ajrny760h9S
iBRGBpJQhRNCej4t3e/+kGUJ4ZjGtX1hD8bmTPw4cdZpmQdDIPRH90V6wXVHXj96YLHMQv/mgKIm
Y+27xAPc2Y4VXvk7Tv2ayOItGUkC4pq9V7tsiLzqgyfIONB2k763o8qwrvhfBSdpyKd/UAXGu9tw
T/BM2DGpIcwKFuSv1WfOHAToAba0tNq69Suj/XgniXEEXWTYA9rM7cJ7dlPjbJPgGdOHsL3gATpC
b6q/sYEAzJMmcqTOaVjahWDidb6z8jJMxa+pZB8Ie2BV8KCGSjn2AQzGDerMrRpTqiVCWaU3Xipw
AU6vyz6KfOqWeF9oL9jhzV59Jr1Qbukt+Yb79+8Z2bSmgT6ge/xhOK4v6jGoD+jFyR6ffTFmf2Xp
vygFQcJQuqv58G5XOkJq4rrN/MGLGI3vfR5LkuECojL/hw27Q/vh0IajGt5tuw7RJcvQ46Af2nmo
5Nswiu7TA+dWx+xWHibjys0NZZqcWCcpRjfHdyR4bUSZ/RLjSrGkF/9G6r4szyVdUQKDRtbr8Ia6
nbcAD/HccRJRAwLch/vhLSYNL0vpLGQcSDOJnh+V2RPYejGN9BYXVHk1S8WD7+CcRUiR6IaOQcSA
zVwjFSf40S7kh5qH7dl7LjUIzKDIkpFfJqeH5IBbAUp/fPFaVoowoyHQOV1zCuSyxYGftF7/lbnp
+TLrCYXXLXvnjI5gmrBiY62Fz2gLTTDp64S+E8GN3ztsfXw1NQduMexrnmiLfebxj9jR1ewS3z7D
Iuty1fUdJrzCvzBbpZTjvSkWm+CoP9YDxMRrvOcVK01ulTe34kKqRKff1+Xv/H6+f7nDjO+Nblj7
DmG0kAxMGOof4gMXxfZza6SaTaikbleZngEZkWIfng54Qi/NDEPG7TZjlwxiqgXwnqnZYYWLx3Jb
cX6rru+oSoG+JY8ORXF7dZCngWLS1//ptst8FQJBETJdQEVaiDhVBFKacKUrk74T3vZz1YMrz4fp
XUx9F28sSDgBPeGMMegRhvKUI08OBUXmNEGFfZOvKB/dhBjhdVPBUmkhQc9qtmWbsYnOfy50gM4D
WTh9wTvR2byffuZcz8S+LyHoJy94g5fcy2KLFG4DjdyNAo+M0myymTWPmH1JQnkvVB0Rm8IVTmHO
PaFtZokLT3aRfAL+noJlJS1NXt89iDRAlLiWhXE3r8CYrGgABrg/JF740xkedKdoErZnxI6eAxJu
BdCfomk7rtaSvzzwLevPY821CpM9vI0R9glYZHp/NKCRvR25EuwIF1p8z3wInuMT5jUkGnGupWzj
UMs3t5e59ta4Sv8P467C/XliMWhyOwwz56F28tA4VUWe+eN1Amo/jYH/KpJqgekzOaQ2f7vLb7S4
vWCd+u9VcHQdG7wv7Njd59cqExhWbW5CnfFMp8A1CzpEjuGRTTTZcIbFKDbeY/+bqICE5krhPWJJ
oeOry8XLjfcQ9T1lhtdrxb6PiHZKQRH9coZDjdejdTFf/b4O+jSx6E1krrqSRZzU5OKp1YgpxX7U
R25vvYbR/yxg54Njop4uzzu5YCoFABmUR7c5gXSqqutIhTlMbx/YW8UnisDTQXodLoFl8cRXmwOu
MHSDHL75Ca+/5EVvxxiANADJ18Gsvk7Dmtub+Odccs7LtTrBRnfHn7OyK8iHwjvkf0uU0sQ1jukh
ltMCSzly3JQl+5LaQnR5J4fkhsvY3rzHjZxColBk7FeXEBkQWYZI/lHMjIJO3av3TwDWT/+MAv+9
19jL3ljfdYCKWmUM62kG0DVwUXHp20KGs57CxpDUWAEtvWQGTcwp/doWzlctV0VwDqoVmZkpqhlZ
EgrgAo0Ryjw9pZ93bMpi2whklN+IgKrCW0PxBLS5gMdiCOEAd6+WM+98988HsDTPLhUT3KWkBR7x
DwTHymkWPEu6Qq9o9P9zkTZLESZQYQLKGB9b5U6eHsKFFd5Vtp7wQOjdDuNQ1rjpvx3dAVyV+Uk8
BjTphgB4i2aA2nGDbt3B/yYn3KKTo8qs/0AtYu7yryfXSJD71o9ROdkY55vzwGutMlBC+Y/9oWvI
6lcN2zd0Ybq5GNaEuUBL6TUKSdacvk9wiIBV59nBd9Ul2++ZW/+RPFeJrtEfDu2TRsV+nziYd6BD
q+rn5iahGBzvA8o2KpFPYjsk/pyjXPVHSO5PHkNDUL0TzW/xi7bNvtvFUIcipfip18tW06tfpDaQ
GJRU5biBUYRtJynkpwRdmQdK5EbtAjkTxrTG2wPIqqJX+MOUHv0FtbM9x5AJAnq6MNU331ibAaVq
gj0+mSvAYcHHSgw7EZqLeowoTukEgRf8N8NCvQWzZrfbSZuqr/GCgfmGIN5pF9WRRM0TZvNcP6Dz
oSd+wWPsnCfskf/3gtrWt6q41+ZANDGos0B22bdkySzdYXYI//yfDpgBvFxrj2vp+sSP1lTcoEKO
JdVuGHRY7ebz0pW/5IWgMm6d+wb52nMTFSs09JpunZ5EWzVbsLvWNPrwKN5PnlC4QxYH+VJratGq
9XQGSrcUC+Gr9MG3V1FRa7b5/SIcYkZGgyMRRSK7lcI++j22k1tvSB5RhcHBxlclscz+h+y62tMs
qIgJDV/f86tDxLWLszHzxMF2cO490wZemFb+rdeNwP80LVukgbBzuCExWl6VYmR0iGJTJ5T3epsG
r/A9M8fiOIIfTLtyTUpa/zpPNzl1R2F7/GqCXe2HW4yiMps24TREa+0W9pCpT62pIkwZy7W6zcze
PbErUcYl1BL7ztgB3lMgJAdV8E56lj0UDlayk+Qs5jUK+ZP1k67S/QoHkD47VbGadY5xOkd8nNj4
A/l3SfpIKvPAgbGRROIrzO7NxkbtTUXexii4fSDjHKDsDa6cVrKcwe9aNrToDWYNWzEy5Rzk1wI9
WlKmjI8CTS1wOsK9HqRU1CdjvUoB1gU0dejdYKUmreu4wkefdiJHWCL3va7Nn7BeSkvp3f2odUKa
Hi60UUQ1Jkup51Ri+gBDkjeJYcnZDHRMwH0kiWX2mEWpMrf7z5eHDgHsS7ZdU9IfB03vkAFmCOqU
k/fBmHRBpwiRUzBtPQ8bMtrJ5KFeefa+QlnqZoLOac+MXMZV6vzqPNUOGR26GZqgDtgC86PLmo+P
yFpSbLPCnTDCjck97F6MtC+a+VyA/KGhSj2HkAqZBh7AxOHy2A9DRF2fbxTGLbYNbJZ1vTvNCHlg
xKSYiyv2cUmcwyB+Bo8lY5fP8eN+2G5afULFEtvtxFvJT7PVs0w5qdG4/jHxb54JhBGpY5kg5UZ+
4vwm+ZVVPkfEAip/6Wsk0F5D8lXTXcJjrTfnVBJchyAFxx+gvvpGrMVeYA6W01Xz735+d5MWlEfL
E8ZXgWa3pZlKC/7OtLR/JJ/L6WKbHJYFBBbQK4keStqKElPTeldCyyFlHh79+M/pMMUgj9C52zEO
RsK1SRHhAmBQOEqVqDRDVJw0pDy6FehUdTUprVPXgjnG6c6KWShGwf7RKE2+aI3Sk4DXHIU7uyNJ
sz+Hl3gelk1t8SecYOgqrQd2beSx0kRb1fWeZkUtnff6/ufkB1qrugnA4L8ma7eCsQSvI+sqDWp4
Ky7ZFZWW9Bx5dM+4hxd+li3QChkepaAOpwc/VxoF/yRpXbLZ/e+X1SZfYRstZDQGiKXJMY7YaQzZ
1BiHvcoRoX9VmkgVSLdEm/S3uxEBsJ1/5TzgYBYHxcNRI8FSr2pW70xVS5Nh7QJTSYAlD/S8Zv9K
/maz/OZMD8twgHCH2vbq4luK3ZzMovhcJsXB49UhOZ3omX65LHY2+26N3aWwkFiPFawQkUD6+hDB
9A3SGEvW6y4vURCVnyeKY8lW4dYx6GYwz2DJ4sXSFQ7V9QsqdaQ9k7om4ojiOEdu5nIpB7ld8QpG
XyRAzv77Aiu7hiYJre2QeKkPgsFP+HDZttRNdoMz1oty0Sb4Bki4lbhcDl4eAgP9RoDFHELPIXDn
keRDoIHjjjSqDDM3/L5eu7Jq1YwD6y/Ip+fs/464uVl/zkPAm+GJgyaHFJ9Q6eIT2Yg40ht8hnka
B1rh6Oo7XdMH2pJj8Mak+wCmwrx2FEsb4mBUBkhcuh748jdXsRIHgrTxU87C+LESVqFmspNGUBNe
LAYFtNrJwN4K4oKFLppeNnT8H9qHRZJyECvqI4pRYIFKZE/1e/DhIsoLWpN3uLohNySI3Qxv7WgF
XQxgoGHPNYEEx7VOeYdtek2ci8WqlGD78Zli6IgnKPIEyNuJiY4besLyjZOTTMnE84IDk15BDFfv
PTNltu9n1PrvhWj1ofj/t1waVIUt1Y2boIFOcAhtDXtaOU7mZM7xki12DvbWV/8N8a7jUIZucxtB
u6IEgGAQHLMa2hn9Q58zvlDFl/di3HBqU6RY9UQPrXeh6L2Uwr/n5vyy6fmFJHKen7PH82YH+Esd
sBIUMk1vSyLmHiOtaikG0vc2K2Fy+QE+raePEd3y7UJHaH/PNqdxTzQ9x72Xw250KHz7gI1YT9WP
Wp0xZBEa3nEAjPoJ7icpbXISF3Cui4VSFUjKg8hEIPpMsG+lBJMm8xdRFUJ8x2MxljkoNe4fITwR
FttYGuSr0B0Fque1MMM6jxIPov5aew4AKPEUFabdGPx7lvn8pXvQ7GuIRhD++7QSbPohSZcpd6qq
roAeSZrNDMf6u+71M7V7LooQ35suXVbM8mzoMqtTAemLB9cmvgVg+9bjE0ijZNWone4OKDhQv9dy
G2yMIzdnrpuPXOYh+PllU6vqbYCF85PEDfHBHUqBzZTRF4UVUZm+w1V/BSqKOKmEcUvF21ErdE6V
+CK26SYnwb2ouNmJoWMLGPnDwNtako7CbjgaQJ+qeanp0c4WjrjyxS2YxxyUKRtnQ2L7qe1JUA+0
N7Za33NEYCQSQS0PwvSjx2btc3B1H3GqRHU/W/QbeUOAUq3tj26e2fi21BTwTTg0hZQ20aZKnkoC
F9ikMSY6URgjZfmuGpHnhhNeANVR2+BsAjlmS3yJ1+GERaS/xRIFE6/nYqrwqtqCdIa7QkRvlrX2
a64qJl2ZuQK6+H9TFmpFwZpAJ3lBjMANBxFtbB07MoUXsMnA8JlzZgyN3WyR1apuuSipFFkAXdfc
aJl8uHr9w8q8ZkADr6byjxG6ImOa9WUcj9TFI8Jqb4ZoEsbJgYeQ2TXFOD+pJEzOaHu1dD+AYKui
WYYjElIUGaNoY3g/GZEXE+nAAkT+c0eiEAMYXGKdUoPiAYwmkydT34fBWAr4wu1cl2rLd/nQLq+a
xMTu5f3IzVa1yvDL50InU1CU4if872pf4diCqeKeMa8iVhNW8xuEYamtslXrTNaeK/UK5/+hWCJH
OAjqI8dpMNow8n3eFNRfIYx2eiimiys9RH4zDctg9+etfrAStNRG2BBeK0IlxJLcQ4BnVha9RLyi
Mtyu3hyZP8UsJau8D4B0PXrkVCsA1Q3L7mOeLcaBDPM1wrix8u20WNzs787vRVbETQbfb5whnM/F
aGteodzjokToS5e31rjCEYuthUbzWOGBoNUioP7UaAaAonapf86Euneby5fD950zXVO0/AtoPcqb
Kz8t0bh2fekuj2YXRcJKnZONrmKwaTbnCUKrBR5jK7VQUdQ3CVq6WemuvVXSReeFr3YzeybpLDiC
yw5e7aKXzRB1ervbX4StfkRDOf2wTMSZRUEWosllnDU57CIg+h5isemSM55hkcght0ANcGF+DONU
FROUO5ETj5VmrQ8kjFZ2MNiOgLS4z+Wnrng+7karpwLSt2aWOIeLA1Oo0gbm83W5qbWkURmjucMz
da1bD6hD7myDAWklhWUiq5crsxg5PMXeCzFcd+n5k8Dk/PD/dGwbTQdrAk4D17m6BHvqoC/TopI2
3gxV+8YkWVVSqLyjs5NInyOZBqtk9VZ01pUdP4TNCrUo1trp6rXyD5vhpA6IdlMef2XzWtahpUXH
isgzz496jZ56tudHPdjh6TSWFUl8SMfOYf3dYuAOUAuCDz5zSbyzYNETsh/icO3LYfY6j29vBNhK
NqfTWBcsyVXKg6HoUc4cc6+7fKYPhgubBAPfJQjqqnWmczM8bjXPXCQRj6FIztbOng4yh03LWWzB
UNMYz1TqM8j2aqyFvvih8a86gmW8AqLB9EPdNhC/y5yNHbW84PNFU/tILq4I1TTq1lCKTDforAdy
1hcIgMCsZ8lFelW6u6YNholIezNgDwkgqH+BiXfnO2fSFlD5lQDSSZLH05Fr99vQuoF4gZhNXlUy
PUU2wJddyAmdAG28iufs7/FM1DI1FDlcGg5YJMMQI62lbINlHQj5zP2k/lJv3tPM8TF1jfWnqGZy
aXpuSactqhQOG8U0gwoA4ESEKIlBPsliJGqqwtqZ/5DFsfV8k+zv8Hh0R6fNcHe3r8B8MtZzb8xC
/NmGOFIOM1crFfLXD7l0XDk4utHaCCgvCfxX8MPImI/wnSjhifht2bkF+EIX1Wo4Fr/m/84Md6ta
KxfcmDXVUVyFdzFUkFsFapSEGbgQqnQQxWwHFygbiY9NC1C4bGNE/QR3DAMFL2Jk93ID7CRnqaOR
Bed1d2SbdLKyHytFZ7V4F8dwJdciEdVpu/U4IZXOc2XtrpgLI3Dsf2sxvesarLGApAY/HsUNIjCT
QBXB3VDU7Wl4Hb55T3zsgqt2OhiSHiz0CukIqMuGzQuBsQj4qTxAIO/mCpWld8LPNiuguoEvcctj
fBT4kuMN4FePCCs8J4p/yIq7jyWVwseKViTF92UIytA0Y8Hx5kG7dbCR6nHWYHyFp+zIPtYKCVXa
IEmhRMDB+EZkfsv6wS4TKUYDe4jqYkHqVlbGk+NH1zygJFsVGe+A3dzveMH/GThI063q2eG5UNbE
PhVWuc+VC3lHA8v7xF9M6w1ncx/D8KusQVgs5XUqT7AOt3WGBbXPSbei5osQCzzd+7vzShaIyu8B
iRmAdILFAcO+rKVMM5tSBjuGIpUXQW8TZhpfiuoqVDs+pb5k2jt93ShWSQ4sYSKGAfM/IAC0HMeJ
7IEQXg3eK9KO61XDBVLurb5aCs2o4aVWfqGP1WlNnZP0xxHgEyC92NGnCRXZL3FmcaQd3XcwoeZ2
8EvAhZdrT+nnLSBDY6cymtihod3xvpDXZWTFqrUMaUaf6ZiQu+PjzvjjiOBxOW+/auwBlEqtzHOJ
0BdIzlZob55z1I3clJowXyFo0gsGL+lc48j1uyti2i0kHH3nPSTJDNpZFyS2t/loNw5/zhq4p9kK
SQ2XWrvdzH4NbfSAHKqEo9fjhZD7HKXxE0hTiYNcl1jCcW7fXdV7VL7yIbsaki14zaNQ5vvPo1VC
CbbEBTCEUdJoNA0fGG/fSUsofMtXF4Aae5osyvPc1thT9VadxQtXnq5jWU99laGiBkQoa8OGyeCX
zYVMa1oamk9nwbAgUCqR/qGp08RCS7AiesuxeAfgaJKZCKYjmTupredgTQjQl9rJh6rLjhkWwgQ6
KDp9dnmC44YPlhAdrAHcvWo+V2VIolr0cVcngjJ5dEDReKUG2KWEggqPS9yfJOu/HSx4Ohcnmndp
Pvky6anvnSI6BCbVWreWnQXsTqTXQj1PmrfdgNlq8TNLJ7quMEBLxFlVltyBqbJ0h43tBbSQR4tK
gZu8cJnXUYUtPdZFW3Al8TkNMH1ez7GxC+r7IaG0avX6iw7FifLVwOuCR90s/y0cviR11OsnSKBy
RY7Epe1yI8G6Z5MUf+5A1f5nscdizhXlYo0hnKqctp9W5SLRiGNFPfGoAFM0jchFERPb1lm4L+CU
ELjy7Ih0epCFsCTjhpW+YnOIJIlDc/J6oJOGjLPZuz8beK6z1VXHOMeTquiIhItVP+0XvQwgPgEU
wB37TO6RZyGibQeBy3T5hYhgbw2Ow0I+rvaY8SLWIiUiCb15pk/qXPZSFlIcd1f5bevL/YpbhcIz
+7dpj++Wyq02Li1CvAslnSMoaWk+kmlNDbD8NBkNG0KyhEgPZQWAtJmpB7y3XeAcCVbOl9gU1kDh
7ON2bYCXePQfPXfbvcWbhTZs6ag7xLeSVX3QqXfwZC1uCz3i6WFNThcEYdTH9zj3J6UpBl09IPsS
J/zFMYk3+YVLi5rScchEsUsvZDFw1M8ihEMH6VvcYMpdthlTdLINQK7H7/FSTURQaucbUH7YABM5
GHG9rHc8jCjHtyV3i/qf6I8tO12MUB63edClL31y6VTMhV5X98O21Nz66lvJpJ6zGGxRXKraEJwK
g8F8YGevaPo5kgRHi1BCj1xm2/tu+uYb2aRWGTRjFs7seSpb4QCYKV3tNDXHNKVNPM4sWBJArpFQ
d/Eukq+8CWw9s8HUqj5ASSYZl/pjPiMXq7gb1rTnVBq7GOM9lRR4soWgUZhT/WuxPTMm24GBVLph
kyXDJ3v9U3iWHeybyomlYbLXFiDTwj0sovKBMxLvJ7VU07yUoAFiFvFHl5xYj7Y6a6+OfJif9lV/
UdOGew9Sq++n9bexqzKzle2hV5cIZ+DprqoPUEf6GDaYDkVTmQcCArAD+Ov1XcKuqrypwHVYR0RB
gZba0JduWu68FbSe3JJzsIxC8n7ZScAxKumXDk+9rOMp6rzG+vIk+0TK9AOLx16jKo3y7BAM1CQG
0CTbz6tFegNxSM1IVtRpiZRkWvNJdMRhqNt1ziGEnNYmKrXpbGnY8q49c/wWfgdhQuRDUw6Mj5Aj
UUycxv3i2T68Mvjv3i5Etd/6j79rcrIfNDhjTbjfFRIg42yEA8t/SQGHaWsJV7/jcf9LS1LQPDz8
xtUx9bZR4HdVsEmLU6txIq+mwJBwnIkwOgXZ/J4bRobMQA+fuDrFyT2PtjkVMMj7Xl99abbQwWh3
sG9Ky4cDi1+bYu7xz1NS5j/95ZL8LTvXzGU8R5M1A5PxptHkHSm1LkXpxofuIXQDUZHbS084JelT
FM48VC8/JiAoCyKGag0meqvL2MY/JDt7XarTIGV0ckwReco6TO4yfPz2s8lGxw/8rkH8OOHrIvGT
KfODdUn6fjnSkNv5erT4oPh3PDq1xYh8y3P7AIlHgVk5nf9JBeHFMevCrCLbfpODMOApfbgYaEhs
532v+G2FPL8IMp6iZVq2L1FfIr9WZ3tD7uc6jUe3TpE6yWnDc4lVPEwL4eGWTeJZ5AFcKAiCiYDJ
mNrwbJCLFQSKPZdOv+J/wMhxnh1xobCWiARfa+R5YDYJs9nXff09mN3+jEclu3MvVXhYit7v90gg
7AM78BBkvOtzYiSnHbcutV4I3uqPrgXmiDVyH8ONuHhLOCcNAzDJ+rZzTVAS/rZ06qXc/KVobJyT
xvELH9TFMbRW3FOkmyYt3EKb+4vzBBZWxauLlIdnDMPk2Ux0x+EFmAn5udjIoINmLrsYj2BooQHb
toauKJ+FIFhAtxqC0DLHlfm4lZ+9pUaaw590BcpT2sySfy7KyDgUqohR+N8VoVPn/YKcseP3a6lm
/t0z5WFv7BplCVpxbNmHhkWr88RpzSzJNf1KM3pQGlKuTMhqGh4O3VPm30hD7P/XNQM8fDe7Mhf7
SqOWmzOU7160dNyQWJU/kZDjpIwfKMPrApPTqXmj5TzcDFmjJ2RGdkB5QRgpqcekqdBPIqH9IAVU
1ZoEBfg/QN60YJNrrlNiBnMITi6tBjS/wwx1CRMP7duWF4Xm+dtxua8aQ46jrWE6fIAc2z1yVKNC
gUPUulOkuoqLMAPTAhh2rEDb6ubyMC2sXgtLydL1ocAnL1WtdJ9MKNDsKND7krERF3pkJNA/7oYs
Sr4NmFzp0ZIxoD9o5HaKODZGd3jdhj88WShIRN0tTt8bjpF2yXtW/vDQdOqEHr0pUWNHfEMHmoLJ
AwoIs5fGMm629YcZdM5NWNvtGgYYXB0p07JuH3NB66E3eMyW0IAxuZJppAvF1QHeyMfc7XgYDeL7
/C4ji1RDJNIXyUx31RH57BY7SKniB4A7kEhNLX8c1vibm1M0TplyVFjzI18UjcmccLzJ8Lat43iX
Nu0t/lLdsRWEVQtZKZTM/T6ZZ9ZjkJWqhkpLTdsdDBeGY8Nm6ZTCxX36myfOPOOhKaVuVEvPIF7F
w76hBYau191nu+CyLxLdGhM3XlZSmqkExy3DDTIBBzq89GOUEVRu8EOuNjpdPO3vulfLeNyrO8xG
zSlik5bwD2wZPVkRRJbfli+eKbFoybj0R8ENFpj9XZrO9ewE6SaA0vyFAhRKgNtaX57Pf+PQ8Wm2
zYyaQNRBpbU+AayPcJzS1+qc0wV1zJ95Rk0Kkhuc6jEvybw8SyA7XpfNxXGF5N3lqT8tgnnpJMVn
6vaASDtoIqL8hNIUkxo03Wl//B4MmG2MG7lfxL+ylmM6oJ+KlpZ9n0rsuYwZCpmaCDiYWEIZwSD8
hl1VnK8pQGq6AYzkDgyTCgxlNh3TvovdTsP0IbXWnnOoRQH/k4Vckw1LFhGiRhncx7OfrDZL+40C
OJqkdDhvvnz2JhIrEvdx6Rd611vZu8YP0kvFD40EcsL4ihHk8gURZFHN2DTP0uHnuZih/6kPA1eg
tDwGUlfNB+ATVUA1jxoCuynXsfWXVzJApQUCM1Qm9qoZHLsCmLS6EdaRU0l8ygZO95cvvnnQ9h+w
nMv2qxJ+FqzISgPH1Hke9hKihZNKomgTKP8jgda6eyhArYP+TQetM3E2QM1tGjK/+imseCGELEKA
jzb6tQsIRqZcBq1Oz1P+K4rl64EOMxfLfcHYZibFgek1SEEwavX6jEJXHiVc018g6LP4he69N5nv
lj5TPzXdhninrb5NOQNdPI7l/IOtLmNG0OYV42i7MgN4r2+jYABNbFpnaQ81HhWaN+xGszrixa/I
RuEP3e82auKu8f5SrGCQNvtqY7VQT3iPSAN/4vFgLsJf2HYlH0N6k+WHO6IznELfj7vj/picXV2q
Zgwst97CHX88xkmIEtZXUA3G/3KezYaMCXllxnbMslqPvLBzxzpp7W8RpOfqfU7kDMlv6PqkVDxs
6mop7GpmrrGTq3XsevHm3fFSbtl61Fx0Q9t6YA2YX32TPhioOEIwm7BYFK1I3zpCxv1EIL0Bk7Sw
Ez+WyCGm6IIu2I8on6ATPTszu+6EqM0G5u9kGCyVJHsFGiCesQI7UIxVeK9gvzuTXQY6O/pbChH8
EWs7ekkbNFu7hVfVDIF7acQhFp+RFJXkh7UGKy5hACx1F1W2rRodypWeZDmqXynezHvvRSwaV0N4
NwNe1QhcMTvDfCjitOMq7RT2n/5Rx5rid5VpHkTY/GJKg7f6JEK1ET/DGutU1AK0kIG/aFoSuOzq
Qhd6pvuXBHzSAEZcYlg4Bs/MxpgbzoAT94UobwFB46GFvm+yZjgFIZ+Jrreui2F61nBuSfSY5roI
jBIDj9chVM8HdAgXA0oTuAF3f1Kal/U8BUYEG/b9QG3qz/MTrJYoj02usSp1/bLsfmW6TtIxsuH2
0pE4nJeLkZWJUNTBQ4FoGYY8qP0xF25Y/Dm/Fl18u//lZxJXSkYijLTn3JE9JTb9rlns2Y8PQE9r
WErucyYIyrSOXv08ltkWLYEw/5BsSQjBZzpsgm6M7Mu/12dKtYWZ0y17DED8Psef11PmiH3WKkhI
y8L9lXaix/V+wYeOXtj6NhlM201IhhIFh0TFm9/FePsTaL9QS4D6aCxHTItcVbnfK72i8r4xOByv
DcFlF9JJSb40D1vw0cSoOx1muYOuDD4GwicySVIa+7rJ9mqZc5IW5UtwYMvVLj9tLFHKVD8ij8ru
4VRYrjgPTGIQgWXXsuBQkPB9jVwpdFSAE4kuU6ldt5QqWrrJo3TimHFbpi8Q00hG82tmmxCKyrmJ
xP8LPm88KRLNFibhVZBWQqyVDZmWvkT2yRcyL6J6meqK3fkKJKEhzpiqzV39xs2GKPaRyBtXiiWS
jmApwjtY90i9umfJoIC7lMaufQkGH57vcRHG4qPaSeuoRp8cQ9YqYLAlz8NNzuxAYYxsJFzGX5E4
UEfQWb7FVTSp1lJthAg8tFcdmSK/Ovr6PavISkdFFSn2VXOrQuEZDAewsDivfR+cLbDgnDU8XarD
mtm3qRaDYq4jhqXcW/0YFloB0hs3x/xa3ljpagd9oGohoYWTXE0yi0eB/TMqyaKvFPRKTJpyMh5r
k5/CH1T494aRrgtTwRnCgTjHrKKT2GD7AU5vieMlsZOCx9mX20CzYoA187G3MDy4eRj1seZwlLlY
XJ0JC1kMjRhSldp3tHNIQt3wI7F5EMpIw9Nv4mawjmdt4WR0tnqdq3gLxwylRL8izipu1KcezSU5
D9ufTNnzwf4l/SFBUC6YM+fYSMdY3+c8XHC+X9e18xAqMJofKza2vhjV4UdDi35wQbo+n2OhfiLm
BMV/3efE5oTHseA2yCQWZDuLeDrGMzCagbYrG4294aAfZpf3x5ghmQdgaem7gLjFfu9e9/w9HCkU
2SMUvKuUMdUlR6F4jHYJmFs+Koyb+Cl/0tCarTwLVa300UgI/m8HD1+2SToE47X6fggw5L6kOzvc
RbA21eo3ZMhsUa7jTv64d0ZMhyH1g4BJuEuVG7MunWAECuMlK0p6rSK5H5g2WvecQN0tsjCVGACt
U1u68jVNNR6FyixXUn7X09eqC+tE04ECt61ujhaoYFRnIOitS5MfY6JxLRQaen35em3epj1TJWqh
kYhT3sbPsmZJIIvGwjvnMF6bt/5DY74bwQtkKRxeFD+ZN3N5N7E4TSkZnrJSx4/R+Vog6N4nWQ1K
S9BDXH5MGaZ3bD+QruUQG2qmCOsOdBuhWkjChOhWYW8yFYQIjmvAjyrGxKNQoGiAW2tvkCkOjILv
muK5H3TXUrLyAlrJwgX7H8QKjED1ourOWDxuyVjhJV0LGfzUHRdj+Ug2pwdK4fkZEwnuNL6HZeFO
UWp5kZii4bFcTiTZJpEgZvjJcJQgtzNTpvF3r8Um2PpOK2noA2uxeph0r3ioj8JXF8R+5IGmAnHV
6rTZitDUIbC6yj+aSjRAFaxxXFW+kK+AvdEAMI4F2UBVWV4EU+Z30pLXTFDCBJZokXms0KkXPKq2
6YAV8rfxMybmMXN56aFBwqnBJ4AdUaYpr6+VuaykVkV//Huuiik0rHqbBah6PFsu502O6qRBDff0
UcuDUY/dRN9I0+irjQPqwUtTJU9YrCSfQsY4W7C4hBG1pZcCcN2VAPP6EFszD4RTMbrO3TDugg8/
/SPh8vdQ4DhI3asJ3xkkNexVrRHL1GDQJafqDUpVHJsqHG5+aeLTJ5vbQjW+/OWjMM8k5FrL95Sl
SWV5Ug3eSsQowaxtHRlMGvgsqa1KyDF15dX35tfbytI7/jqPW2l9Pt9Q+gS6nIL/9lWg7IoOPx81
d2UtlXpWn9m0I6eUDHzfE8wEiAV2IU/CD3OPHJ1MwM4obIQ2LA8CJjTcGiXQrNrxUjzhlCpny/e7
D8rGxDb/IOlTznMcNSK1p2vvvaPlvIcPyGjAv1soLsBZqLv+KTBYEv3JBQW6QT6m9UKDU5ToWkMl
KInXKMbrk2K27ytxD4gCljbRdGMCgTYq13PedZV9F/QCLa4+nsHKEm7QYo4pzlH2nxBBd7Bfrtna
YNaLf3y0AWITO8EpNrauwLIPhcl/U9Ix7PdGOGTzoIN0x++fQ0xdw5GTgSk6UqmTRLjqos0A/TRq
EsbTmzOj4doPTM57yEYMWNe5QMiOSZ9J7yKU1nFlsTNRY0kUpOr6WYAuh2xG1ucc0fh0ZX13pHDq
pQXutj4bPbT5AXjLTVB1fuHChR7GxngsjTAOc4h0J3h+J8RktYHUsuZwr8uMT/bKudPpa8gB29zS
sfzLWHv/zk++ldK2JA05HvHz3Vxb2YAVm5XfG3YEoMCcZljR4TVGRvKk/eYc4HH2qZCgKD8gpwfk
G5CrJajvWEREE/qSqxjTeywq6PYxdshj551XjfHijVAHjttMBmxpAohglwwISVOJSUld8TL6/dp7
lwoEW8qarkusPFcP46K729CXkgC4RorTvC7tZSL0h7cj61IW4HjZlG+tvZxhpbtDyIe56QMng4vJ
hqJUMzFyoPdvbEeGsebE3F4SyPrppRQOrRmIZHElaVEpUmq3VAPv5x3RjaNRYyNq3UwZp55b7TLa
ZihHKMowQ5YBo/Mkf7ix/pInsJkW1A5XPmpu+NLkYXf9t+0a3x+FFtLqEVkKn9r4qbsqMfZ+8r/v
W2qJvbObU2fxQUd+KV2y5QJAtcz0cD04dgeXXfCOT6X565QQwu34qgKK1k4yHSSeD3WCoo4XX3ln
qupVx/+29RYIYw681HjVcMtHrRepBTllbnfzxw/vG9Pgocjyg1Deu7RyMwSZWeT+fNG/c6lAbDgc
sFNZ7yX3Q/equ/SBo4iM/BEuy7qo82ZUc5GHJsEpd9/0QHEQXLmsTUYpDjhOA8B0iS/ObU4gqTR4
g/g2019eGOWiRKpdltr4+ESYgPgJ0XL2CxM79HB4I4gEzxby7AaW4aV1alBy2+pt6f0W02HwOmiE
DfVHDiJlzcrR/reEHiyQa6rS7RADITp19Oo1Vu9DeaD1kHclfdAfQqhfjrtHxzja9rsYBuRLDSO8
JxjvTSfnpzoLo2ovzEGOjZ0jE5fOzpl4bxx3KOmkS7pAl4+a1albTAxvX7NMxivkv07WY2Oa9dqz
gWcXFC3hnYcCK/TIFTMUwq6zDtNrt3CFf5nKiT62Rmf093PSamUUA5APFPkxKZR8P3cHA9S0O7Y3
ILahgB5mByu9tANP88f0i5kX6zVBHa079J+b3oE2CFOXyB5SflD77tyw81LZZ2NcRgm7yrQR0i9+
/SDZazeaKTrrOSoIPNyOIYIH1NyjWN6BJbwUjxf0AD/rdSJweiFqy5eviiGuG9fBxHhSE7pofB9l
dBQrbqqhOxFECNhVIPcj93/kq54zATNc0YTv9fhS94IZtqR2X1Qwt9D1xQ25sBU5fyyQqo1x/d+P
uHFeK1zRTTNFzwMS/fWzqUTONhPtK86jucOErzHT79eepIxbLhBOl2nMGs5ibIwxyVm4NkIHiPI1
LXepkFOzi4oyztNvIud2toJ+k/ZWTIsG0MVGzANeF/gkvPxfMi1Hqjtz4qXVkd3bjZeMyBu+Hy3z
xdNP7t+w06aGi+ZoUTSZ0e2lZ7zYRvjF4FLcl2xlfofaP7zi2SMp4c5LoQ7Z0A3aDEyU91qiJa/A
021II75wEUrA+HLtInAQQpvBomc3gd7LRtUmZMYThRGmYBKddMQIyLSD9/9w9/7jRg9jWvgrl5Aw
TD4COWZoE1dSXMyiE6tFvI5RyWr7Bs7touaYro291N56ltU9MCs2TvdZ4Pg0m9v6cxc1RWeBBe0g
A/KsEtZfhc2FKOevQDEvXD89Bfo54Y5OUQObVjZ4rDcSbFm/sV2sjV9E23LY5x+5Nq2mNqz4dtNr
b+fRP9IfNOZslpG1giVGgKBSbRGDwKh1lUQbUcf2HZ6atH0ZvGEk5aD3lSsDpC3Zw3ylDV17p1MQ
lhbKxwrBBrP5gaH6Jpj3frxAbRA0sxdkU1vSn06svZU5RT/Qj7dUHli720vGkkbZn+POjuejoifl
McO8QXv7Masb9B3jVAX6DOcgeMgwXl1Csdi1ZGvKMICttSClBKbQpDOyVLo8FUlBMLGb3x0yNf6M
OLhuelkbd7RfU48t8WvFWhvPuFpLC2YolEKppz6wsxvxz5fG4yy8qytsi8AqpuXsj83WgEj+6hhC
l5dB98HPukXWgY5nwWmk8E4CVjX+nrIEbO+s+6ehgY66QFLRwlM7nVrIxzgrJkW+1QD5D9/FU3us
Uca13Da8szt/hbvvNpL6j+2+gi9j4Uvf+jUcuhaoihtQQpNWMa6rOHRoavix7Y2JJHhy32tI/Sju
wan37ZAq8PPPTYcFzevyyuvhMASFb34uI/86s3yKDIFo8D2NFm2vNN0zgvwr5HOJ9VBqu8Q80ufN
wMVKplqV3o3lisy2aO9ccrFFWCGHUijdC/H01hauzq8ZYRA3TaM2+ERVT926swd3AwNN72BykMA5
Ms10MH2d1OWbDRCFmIReG7wFI6bFXzcvYfe1mOQxNcdASH2CtEZdeB7rdxLSSyUpgQYLg4aAlJ00
nB37hcj6CdmC+9pC3enOPtqM6SWsDTtSAumBOwoAa1y6PEuV0yhOu/Nwjw9Vt0ch+wTjgOijsCjS
KgQDjc4sELLKyLhcBDGJ+FUiRnB7YjUiH9dP3H29xNDblcH9hqXPlMfrxHcNfiP7oGsrxbSBMvru
cM2VORGfgoGeg1ZpvBoRfMSAz8Kazfpvyp88PxPRu0ran6X30pleckEzTO35RYtVMifB/kCNkwPD
SO2tFpRny4I9kGrPv7ucAiC2UDnHZvXyRZMqZGLWkRcDKbdVS22w67+461oyevqM3kIwVrsEiFVE
Ser/2B/cOBEqf610rzgD2+7QDrkiZpwot+wNRDsrfdV84lB0INpg0qVFZKClzIU0WNLM3beKeFWc
5irHAiKuPIB2AggIhjoFS5a3Zf9cOsWTzPmhfzrR7l/0UfiklV150OoqxDIBFHTsdpL+YZMAE/uG
VVhtfBZIJyDeBZc8XgdzuEveGuwOU6TS7yKkQQxSHkRV5GOin2rFHuMC69JATaVmgkZ0gBe6RgRm
Ny/ghJWov71Etb1Cpz07lZeKqzMr8WZ7OU2ezP4uS/GxnCTAx117JH0qa3EvLe93Uva9ePerB6Jl
X+yw7fMPtAoxE7l9FKmkxebJXt1kHCOLZaK7zRNuosJ9rFPcrbEbLH5KAj9KnVIqvOcp18iEciwm
7bBB72ELG7cCBkU5d3mx7gcSHIqd1eTB4nwT9Pxu+Bm/rUHu1UDdEmqeFvSWUj8JxOazGQ81q7cT
GZTg0L1mO0TkyyKvTa9aEGioFZWm59bc80yOWHjIpvmNivp6JPmN1TdWdf9IBbRBnxGo3W7X6eV7
HEHkIh1ZR6jSTLWf4hXGuwWRHzprOae31IG6Sen6gYiRaOXu5iw+TeUagYTHUSKJINVdYo3Rr2PW
r+gThBiaBoeJsoFpKiyi/3y2++JBDqTzE3p6se1DSVz85TUe42pLR4uCF4KLvVZeqQ1/EEKAcquO
rfIe0Un3bWNK3FHpLr8h65IwGSLwMQO5cYaW4mkP80Y7UsIAd87ciCmK1tK10ZR71jH03fo5C1C+
PSfQwke47h3aLrPW6+9MjEm8LWXMxKbKuizR0paqMUDqRc22rcsNYLx6ccZ70Unlbe87kcj+K1yU
fAbQJM1IX2BzL3zKGKiP0z4ABQneNYvmHRvRnqHTSWrnRfRx8HcNyk0v/vXVbpkVWADhieAikRxr
igAMJfug9w42ZfT8Y8+nJEweK0x/edXCyKfXjYFingDFBmQkN/0oEHa1qaDrInwfj1vpIIkxsUW9
1zLlWa3bSOfvq4AJDeshhr8i11fC5D73/sGhKX4AjUDIoo6OAAdWyO2ZKChhB9VC8FbtXDiNGl9e
vyF+IeEsn8zUC42I/kA5DJpfAGwdRowLWgPuI1gskpMv70C4mRn3ufUzTkMNoGX7dZyIPcQS76Rv
ZIFkFxkj4sEDXqUk5HT0JK4qwZjDbuEndYLsYjtKp1HLUIfxZ2mJq/X5b4WcrLZINN5GURrlefqi
lh1WNpf709FW6nNvRbNo/modXyW47SxOp5ZulUV6fvNVofyY/T5wUisB5WZDBIggAcmGvIKYkKSM
tMNV+zNp0nuft4rdYGF91JJgYSB4P1jU4myEokAmJqY1N9yKr99AnGtw4mEUtGDQCP0zE61BSzRu
TMF2Dlrb+Wns5Q1ojWdJbOe397z7Vy7uCyWPDQxAHADokhlyOulQEsAsLFg5yRBKm7yfvFIzm5KT
McGokJXNWt1+a5xzCi/vdtD3iRARxdI9x+CaWOVT3I2XfgQbMc9ZyabxQUTqjQNTVUROyczqDGM0
xh3Ko93tGxnFNU4efqn1Ki/xrZbOo8I2ft+rTv9UNJw597Rwk+Q3aJTD97cVaoFG4ZYRppfbCjdk
JUoJdr4f1lgITxIxLo+6Z11NifI7TcyMPVZXtSkiHLqfaO52Fqak/CBepqkZR1Qw871arGXh0tNa
iPwVO6425/Ch2Th5MKLgHU5beAtQ0iz+Zm8Ir/JhNqlxZKlN6vBrbsfsxa5BA1IrhZfjso+rrlxu
uZ2sZYEzcfI4k2WJThRIKnmEV5+61XGdz6qFltKerveABgxIZKF8660gBS1Hl6EviL+cs2NtWE3b
BiIfyPQnFFr9Wx6JejvJx8Z4XEAbbGh28DycIJOsvBuPbfcLxpJ/Uww3ChEWTO+ZWTQJRX7WPQRv
O799BO0D2UntEHaY4z5/YMxwMI4v1oAUpJAJl4hCmCZxPU9Xh7ZkDzi4bebnKSf1ghTfws6Avrh6
JRLtI7n2btz2bVUWzacF/U/1vVxDIkglnWJWpxqqdcK3UPE8UK+EKdraendjn4k+KEta1aPs1xWe
6LyrY5rrtzmshcN6DxC1aoFCPHLfvAluizdNTO9QORRm5zl8cmg1DWqWCnlhgQUdn06D8j5WCJoL
vTB028kNoApYxQsRoXCGM8sPut9OylSuEE2Va4kjOhiLrEl3fW3KyZaTzH0Pk+qqsK9Qs7xhOUc3
ocP+NwBPu0DFb/xYntdTspkazz/mVYi4iXwpbWWFTgAdjSLs0P4vQ1OxiqGYpGQWikObWGHTfWaD
FiWhNLQsVdjrvcjXp/jFKIqqkh5HAQMnjdXsmrOiLZJXOxfPujaM5dskX2Rqlwm2WhxXL82+brKB
1a6Y2/9IhPgYNWEcOUbLzdSIMCcvEOsuGKO6V5V4pn2BCAw1w8+s6Da5s3UuQ+/1OC3RkBqxX8sU
Skz79RB3K8bhaQSZoGAQbaLJSvsQoyjHs5DKKgUyKmDftQkgk4dQfKfUg44UDKwwy+TW9U+l3nSF
rrZKh7rgHMKv4d2GqzEQTfz9+kMtoyL+iy0kApP3vrBFB4xCsAj80lBDszrdJlDcP8SvH/dAwIAR
KC9DXc+nbPmUH/7LYhdbRVfovOEK26MmcWb0aA8SHfRXBLFmy6FxTAlyA/EtzCBohL8KopOr4RsK
zl7m7UbgHqTHeBJHxYNG4q91eBDg4B8NJAOBokM7x6bOXPDFyWAxPvA3Py8ApSIxlGE7+A3Tyb0X
bTnAyi13zLr05WKZWK9Ac6IQy85mg+VsTySYpwG448I+PeGg8yfCkuz90qAkphz7dMC+AbxnXR5W
unQa3Vxg4V1A/cnYoKMuUxPLBN+MajgJ65UcKwx6mHVsr1OW7GHDKkMpZiuc6v/JL9c4LvQHQK6y
+uYVyuu5itKINP0VB6BGOYAZKmkl3+M5ZwtKr6/oVOpzPrWmJWmGQ1cinyY+e5dsfKdbioeKjIJd
t06PdA/wiWiYoTn2O+Q1UiPijIWvwqMXoqKXH+wk2oHU/aedfA6AJhMYj4ULxeVU5ukB52CJs4J3
KTiaC4qxzRgp/gzXvIVsoWSvB/UlvPzziKcQcE5MicrNGKLEPCvWQp0OZOwSwBMH2zshVSh6N0T9
8KFgWt/FopWf+ZMDpkW1mOEF9RGeF2cpQnHzzNp9nGtFbDw+Wmgd+tX8t4Oyb/LF5axOADp5Zewx
5FY3Ar9dg/OuMKw4BkcBOeUaR/Kp/QXX5v9zuvIW3pIVrqJGHXFbSQzxKG/jSlbRBw3NB8KK5usM
w2w3Pw27rPJMdQEzUOdnKvlsA0okoBGdyf3txkiYo6T6e0Z0i6AMuXgBmNSb91sY/uECQmJhWODo
GCd/qACtP9RaBPtqq/Si1i/cV//fVsl8Ja58zOjsW0M5OX6bVpw3TfJtmH94AaNVOxeVMP0UIqDL
5s2EbGZT1xGBuEgkBNB6hJVX6ksMkXGDaPABMvWuZBvLp/oGic8NSmWtfX57abIoTtd2EM44Gip8
eCaglPBHmLz/yzcbC1wHJsOXePECdq6oAjhwqpz2zDN9AkQpuXK3J+C8ojYvAAbfTm+3PPvQ/lPR
GivT8ISmYd1FOl06ZEtsLyDQKriKpFkx3BPw4oeMyiOpme+dji6AfZ31bI4mQHLl2n1yBRDK3JZO
1kb4tB57NrMHVvWru11E4dUbInx//6hl0yd6Sr/Y454XbeU43kXWCjj1TPkiLBhnJtp8aorR1Td/
5HnSKEyEJWmi4Zajz01BWQVChRnh1p4lvptMFftAkOkEnHxGe6Qp4yc/FlaYX9Kf5ntZi1fbsGoN
Q2BuhDoZ31vg70bz6XxTqPCCN47yMgprQ6AoZPDcaRDlIH8QQ9++t5uKhbnFjvdfZCxJnJb5GR7F
3y9xzbZsiTW6Wl6hWkHfqbguaJh7kki2e/CLIyr6daOmY5BEzpjBN1RYeVa8x5QoBllr5bD5bKy0
pbd1cNx3jlMDY9c8oZj/j7VtGXcjYvep9qRnuGpStPNemlINRnwQsH3h9o048Fev+pE7E/vNXqsI
RmqVrU9ezyNr7tTOSTzk+Uo+RVmA4uA73/C9ka3nfmGA6DWrTtLw+mFkK6wldzotDdxlOyoAmh9y
9Lx7qliZ1wkS4dJ5A/AO4RYVWyGYVrExC9NRVN3yNr980Z52Q+R3vdc4N6OQoElqHdoJ1GXRuaah
7kX3WqBTTmvzyQbqXSDoMlbDrwCBqFKGgA3ZKz1TDu4SVPmrm9FrnhIQuoPdn9XHNI+FmTqbpJby
0UGiEER6TdMZZC9YHN1MqfP+gkU1OHWWdTIk5ZawA1ri/TuiekjuVT0Bu93bU9s9oV5FcJV8SYM9
LPF+vm9sxYGzrIRh+v5+ozmrrogaoLzpzYZslwV7YE/YSlX9LKz7hTOGqEoxpvBLabnhjg9RF5n4
C0gpfWBaNTwNQV80OGBun7Ig+zHNooJAbuNGqzreU/1vHIlwq/tld87VjiGZKBlPDniCTezUf1qa
x67tsMrgy4dSYZOq+6agWt1MerrE/zJF8B48zQvdm6F8X68GKhzi1DHdc89USYLDAYSQaLWfkC09
uu8z8u0r64rrrThVGyGpnx9BZ8NXiYABMYMQdqPoltja4Qo15aWYwv0CtTNuucmw+wQ53CJBYm7K
WrN5HMKbn/lJAT7gE26taI4jIQrORETI833wA3UaX2UP5hjl4bZqPM9Vv8+JoWM6hfKDEGvq+H+5
I//uSKc/FBxWd5bgB66tJUYM+ghoZRuA42bR0nJY/7roHhsNWdc4tpYsoN1JlDsfxtwlBFSW4t7K
H41otRxnjP1B004tF6JwVH8PxlsLIVpYEy8drCrARZ6c8d7Prxa2dD7OWlsk8aY7HI+JNFhZhqx7
BlatuBHYRrijbNjvv03Xg1IeKGyPOQ4fN35XNnUn/aslDeOnWITP8PeFFD8pOerFOYLPyiUwZL4y
xicM+0NP8pUr6yc9ToZJoT+l/5tuUFIilji/wcVeu24vZBev+fDJAbGiyy1QyHzgPX/owp61RBJ5
d2eIOJtdxw5a5sMrEGVfFEBnZxHXbnqlbhXTu9Dlv4VOanET4nt6Xe699UY8PR4JUEWdEibq+XMP
wqJSish0Tcyq54c6TgH1d5gfBgn0ZeDziJiZeRwcj2yKoZI74rnsZ9z4mHKkK7U+tLylvYOQUSR6
sNdKCYNz7/fVONGUy8/AFiUlJDkQaYBXhaSu6SpPmfBzbTD7NstNZxwOPr3Hi+B19bFthuH9pPfe
V/SgHOcUzG+IaGB7X0dVx+UZbEXKnmdWKQJlv/0NvYWZ2yj6v2nTqlZi06RT85HOcGLlsKySRJHU
QTcNv6CHjXldm1RGOCFJlZoc61cC+l3GdKkCYz+RVb+bQF1ATyk4HDjB8mxDyU1902OARFOrEtnw
xJzE20Zb6PrscpCoa7zxXJyCNr5BMOwl2Zm3tNg9wk+6EQMiZooCt+icSdEo86apb2e+BvJ0TzYY
6Gsu2zPqAqkfgGAfQEgENy4JR++W1jnR+Xl5OsOtWTIA6ACYBHi3FcSuD+oA2JUGWc21ekvigioS
0etdPkGvLTZWYWjYs0WSocvqm+ZoX1D7ilbpKMi/uDGNuA/Irm63hTW2eAexBtqCjcsh4VvUDcVx
NZ5csJCvbelwPUzez69K7Rnldhf+KmmAwH4aJEa8tjnIU4/O69FlCUmMSdyJKquke+N08GXMmK4N
9MdCXmTjwoKnuTZzaV0EcDyAaiC4SLq43ZlqtgTs8yyspLNI8UFgYvOjRChM4FH0sWzLQWFmZm64
8Rti9dCkYtIOMfeU0w9Ozb1EL62uHK7+QeXz6LugKHAk0tDT5SszwGFm7Cw0hDSdWDUHvQY2cLK1
X7AHFLp3lx8k1MZkKVWZbbYH0MJ9Qg+8LRkzE1pJG8Y1c0GLkmp+gtMjop82W4nuAy3qrhMroTt9
n7d9aWBOuY/6ITs5KLbtmE0rdo8SFrXF8kjed32D5rUUAmEilc6+3jtDAVS7LIxQuiAUsEGr27ue
wI8rWuLyDxMBEDrCJJVlQPdBgr9uilZYvyXICjP0/Ir5KyhbvLNnKS0XsMGaxBEm+7NDGOlUbPCA
m1MYagwnnHZ9YtIa/WGBx/NoxPI23Q2McnD4l5ElUkEn+0JeL1KRJwMcHAfeX958JYRe42Drzs30
LwRec3PdOw4kFV8rKAaym5SbrmOIy2/XWg+uNw2w4vTktuXk0j6DlPId5UMO5jY5tl7r4QJBIRjJ
6MRf8RI4UOL9XeRTushM6JbQ1xowTcj7V/4DI+xJr4et1TsnEkCvkWzEyGPzik8x5/AqxpTDnQPs
PGwvFcs2UjwtEMvahcZJyM6NbnEpLMTz3/XNYX9T1PWO3oLe4b5je68uSktAW8G0xKaSFQnqC8KF
qQF1/7vYDynR7aS++/v7wdaY02rGGMZbz4wkv7jOAOsMYh+lcR+JWLi5lOsOm1B5bLHHd0UJvbIT
rD10DlC0914krEFY0DuamN3okik98TNjjBgC+8tLmJR0hG14NplyJEWpEnHuXpr2fHxtjLBqD2KS
c3Nsj6MUcJQEWVGZmWQ4R4JuKL+c6rsMObpuhdsUBsh4GytxEgkps/JqPpd6NKOU0AaLJ9Ymkqpt
X+68csFKxHnOsvgOPZ4lsz9T2XhUGvTNFuEo4Hjq/Wu2loShKONEf3KTxPuZx9J+CxAO+fgnSugH
kPRj2WeMREWd7PLF9JWa5ceEJyXoRHSAu6R0r4Rbeg0eWlEN8I/LiV2cxvpRs3mGWA//3yODXtlp
o08fKVHHeuIxUOc3gA6jPtG/03Ar3YIxpJukPhPQIJWmVjakBx6vfnHMowZyEMOtyTPm6cyQ952T
JoBl1V9QqklUqbLW2XSB+1mW/5xbV/GqMKmU21jVmT5rSqq6b0LilHeMtKPk9kR+vZV2t7ErBmM4
4XAXtPuG1dq9172YcPohz+mf7bl0qcZ7l6FWHB8ffY0SK6Hll3waCvH6Xc126sYr64ObBukks/mq
2TYuDFFgrT8P2uBUM8y3jfgEERaCnhpgVaYCYL6zXt9IMPlMBYl+RWodfzJn9QMBSGiep2Pi7RxM
/PUltle09usZedyzjwbgA0Rctu3lnGDHDgGGOTIy0RfezZwQd1ICTy3xeKgtNwhLX0vZBO4hvQUh
O2JEIh90lfAuJBrhiQ3r07omBGBhdyKUlcHNORuNoURPYdzrOPdJUtSKJb3DDBbhCpg3pu7jeMvi
OYRPiSmi2VNnD4sQSDZUfSA7wPB0yJDY/bEgYjN5Y1o7AvdKiBnqxBSfkYHJVrc1vuPaPI+lyPPl
wTQXBAhfo3A45rjr2k6mskNbKDu4UauDUmZZQoALQWP59OQAjV+PqAWm+o2gJdexdbpyktjIvuyQ
orkSWQ/pvKLFY+bh6dHjPvXT41suTvVlRrUwV0higZqyurpE66atLmF+VyCfSESFHK/1cMQhtqPI
bwznzdrq/ucvdmKEgFnaMYbBR1PVXFNq0JlTzTVcJWdGHK+b9illMN8YN4jakyek23LXA75XbfQi
Qpf0ILxuMzxGdu3uZXYew5zgCAV4s/D0Oz4Rukz66wtnBkChBFosboJg0D5n2uUULNMuF7q6VxhS
qqhxOOG700dWmPCtoJOP/mRgbNgkPMFYvcgWtFkPZcPaaDyFwivqSmC0cuihiS6bBUU2+FUENu+o
sjvZYfyznvtYG7DOpBYwJFNk9zezeLNA+nqQGfg/vNjX6pXJcRgO8BUtnycO8wFBI5Mt6UdAePM0
hWL7SVrAFRGpP0QInVYJk8+nR4ZurQ6legAVUTBMWsJf6Yrpva+bhcw3YXqWctWqJdlHWyHiIvZy
Cl+UrhmbXRyDKic0ABGLFeXzXKt6lO/ZJ0Nh3fq4kpugg8qvOYnNvjARB8zlgbVT6YzKdr5loIQY
KuWApjScBYBE08ITnYPkbcMxCTj/ab6zl9tfo1CgiZufiCsyKZG4nzlhDKP5IjeX632uB7wGBCIS
hYrxUp2Eh8TvXqhkAzlZ8GeyNhnw7aJzWdjlvIOWPBsALRLhoe2ogKyLou5T5aT+5/v/jhAq6Ys+
GOYF7G5iuMOL9aRjBMQF1SvaChgpcga3n8+qBZImUoUdr02dqjewk18jcjFKOBWNP37O0pWwrzqa
24H9xb+cdURJ2PToxQzt3oub8B2H5zW5WyjVIe7EmYFaH5G1COaXCAT/lxoj0OvdtEWxEZ4QyypP
dcoqqnmDynjqirsIn+lozvrzrgEhfVhyqm7bmbeDjEuTCxpMVIUsLZ0faWV84DSbBC4uYM7R3EUz
AJnIPV3V6kyS/fhWSadpw4ZsAYNCXXiDjvX7tDwcWqSxioe+j3NNGwVguuaWHlQh3YBJULJV96w7
HgQOrfhV2L+6O+qXMSHVBb3+Rvp4vTTzg9iIe23JCnEyywSVjWBrRnAnvnX9R9cC3pWE8Exyrd/P
xl51VGyvQ0ITSQkH+3PgybidZbvleqBquhFRvOl6YxClKOHJ6EMmYUNbdAcS4+8T7yZ4HmW3uUrp
cUOiRKPwFVd7oxsUTqqLhmouGDdtMeT18zvMZpzvNTyXi1o8/DfIdVT/RqrK5ovXTokhdFqEOtwU
jP7uxoL/MOTPFAX2n9FyN1DD/dszoshO46OkSZsgis5A22Hs68SR7kishQUJ6Do8ukGathHsmgQu
Z60sUnaZRGgZdJQNjvzvFQaranmLo67pbk+q6FtfWANUO1qzyA8wdehXMah4g/ysuOqantNkgvXh
egAZ2p0SEL/XC+X/ynFCm022phqUUc83M07SE+MvaacKUTVdOpyA2ifcmu7ykRLj4k939TEa9xnq
HSdXVmI/agecKRJ0NBY+DQ773hPsqtZcaLi0v0oGk/UzYidrc5IBRo7/lAA8h1Q0tV59nt7mRRr2
rJKS4emJv20NAY/6bWQhzmfxMQLRE+w1z9v+DrBQRtEXtQqwCSaQPPm0RJoVb7qwN4E8izq6N6b1
GExmKohKSl1Ih+99n526bwPe/tSQJXkBv/m0EYYi2vG+N3TI/zZt5Lg2Pr5tSKE92RQgHpHcQ3SU
NgR4vkW50Sbv+3fllHvDPPTvHJQW4qC3YR2SG4EODhQRMqW/aTAhGU61AItZeTurLnawce+cgz3F
pE4NOPOmi6bbk5F3PWuKZfnnaZDzLElA0IC9HSP25lnYwu18BfBvKDMUnq1Ekz0P/jEiViSJXSy3
Vjs2/YOFQUdvhOyvVZIT48bRMEQQtWCtoBtYfjANIYxIwwhtdhDQinWlHxiGA4g8kuMA6rjku4AW
x+Dd6Tptl3q/Fi8ArZlUwTYYfMXyyaDl2kQzu9UyOIqVELRvVoM8jbpwhuTJhtmMEJunwZTTDYHn
pl92lls8TYd+bHNkV+bATaLzBgb1mjan/jV0VANDZZ4pgHj6WUq6IRBm+DStHMbklhrU+AOfCSzl
ril/DzAaEpGc5CYZ8RQ0aslLKFSmibOSINLuXtu61YMSJwfrSARnOCE0bvdfwnSotvOrl07wuUID
4FNclFGafdF/ilaiWt1mh9Bbod3i/utrhEZxStx+VHBoUWhjVVsIAjZRvZt9J62eb75dhHDA+/4d
nD5hbQ7WCAU1mANPFzw75wlVHE4wdhB9UPce2TMLptOeiSxz64qxmgGQV6IFjPRC33xRoBBDY2lP
WGzHTMLNzwJ2kjCORR/Hd+Sf6x2F85yPFvUx+KXsKHbeE5ZJrWTc9mzpZS5U/OTcQi15iMTRl5QB
8LooUUnBu4WGgjoedhxn+Mbi64gbarnS2WX5rLqqxl7HWKjNx+s4cynke9ZlHtec/wuTIiZ3P+ER
1hLIjueVSiPfRu8YAJUVYEjeUF3iLG7Xfpdn0PBqqGvriVMG7YAvYNQ1l3BXV0tABldi7FHiUZyY
qOANGW/jRAnlaSJZyuh141dwVO0T70zVCmhbNG5E+OdFAtwLF9gDveUZ81YngWjZ8q6wszKqtOwn
KthSYQJOFN9KI2pSHwlXhH8wjaaYcU84+94KgA2naRn/jtZVukfLWOARLas9IqcW6SeihpHHTgn4
uDdUnVVg7VC7xsP8k+Owev9VIvc3HMrn6dwAitzXdGG/CMbNGRPOu1ZRxo1bFubHHQP6OHa1k3Mg
s2ldgjUMqd4+t8qwNTYSv58wBVHG2smJ+D2KcJGUrvlx5P7xCcxBnO8R+mHLsSkN9szmo1nO5KVu
UKxFqd+K7T5oGSjiOpcZ+Y306KLq2JdbHOihNQRi2nFlH4F81iMhaAIFUWmQIEVCuQnW8IH6cuVw
5jv9/Mgy7XvXd7QzZ55sECKlxtTLED3TTeeXcb6Gu8bvaYLdEaZhTHaeulMSVM8i2yq4khud7b1n
rwcjHayWg9RMhpY7toasSNcKmVNNGcUVFk0HBCJZQJ0KOLwEpo3KOkF+wgzNFqroiMzMK9I5xz5x
fKOo2UCbMpSAXuO5HjKbG2Mr8w3WMrOX9fSYD19H7Gpie/8xErwQUWiFP6eIj5Uf8e1iOR2QXUsE
PuGNVnUEmDq6dxUJ72AfBdiiTSgEKNIiY8SEBIGKrV4UZnwpXt14xogm//ZqCHzIEmXCl7+VAB/z
BYiyYrSmuHJmJTN8P0lHfan13G0o3Zne46bEMtxT9bkmsq7paCR/YnXVQ8fWtwNoG6QZ8g3LcfQu
yhf6z9ku6PUghohMBeGzlIxQMjet4agi0mhnSQ7i+6cKAj0ZNkTJt5h8WI0MCroFeZ9pPwvKAT57
tiFv1TLLK4KzQjMtJdbMsLdlA57YzS4EBP6HBNlP2k+XadkoEQECMBWKowaMZ3E+Rdp+fbv8K11Q
EzPmvhtQ8XmDxgvV0qdXxE3XW0kwyZEUBihPKYZTRucLmdIP1rTFVTNJoYW3x3GzYVTHRjLJSyDC
PSGd9pQKM7UngrZrWfahacnoYxGfenahsEqb0g6lQCP1DCjfbirMUQX0ZN4t4Q3qhkAvIAOVS2sB
lbTkR5LnTyTNUE0IMvk1200RF4CbQWulrdDgjheHoPbW7CGMSHD9lZnclMrnNIOPDej/L3ekODpR
S9Y57yeqnqCs39e2341krqZqGXtp4cA8nfsdjVKBMGP+yRpwd/iCxyzrxjZchHVhUCR5mKV0a8Wm
cX6a9FC1cQpoK//X3djNWTgpiCZofEqy+V+ocgBM4dvWVjpzUrZyYhvWvl+ujpY2XI6rZTRRaVFT
p9Z1FRsD56DXOWn9Y2F4L9Xh9cIgCLtpL0uIusBryMhMHhRj4Rhhjsab2yeQnGoOvWJ/0w73UetC
BFX4Ke55EmAnU+PYS87wf3Yzby8QtJ6Dc1eAcMAvFWHG6TdEm3E6HIxzaN+DrkeuGGBBHhOsn6Xe
6RvGV6F9vnmuCZ8IAh0t9r4d4ocXGpIzIAjR1B+A5lXcalByAGGQEnxb9fQDRSqXs3O3pzwrUGcC
5KbNryGZImQDNz9RNtOjermqZwE4U0RrUs2xwpP9Q3zeAkF7Utqixuuaa2bKFD2ioQ4A0BLUCeOu
SMhOqe0tlWIu1FW0SXr4+O5TiqbgptTeOAPiBHMwcM+4XT9dwfKjaQWeBG4grUd3He5SRimskLQT
aYACtTDicbaPY0T29Lh53BBCxkDJwudgD7SqqVzF6EbxVN0fUZ9JR9zMuQd6DkWNi+ZN5WzlQh1X
3227qPq8lNPjPGm2+Fh/wjHydfz4E6OkwYXZS1DHvpkWQhIJKtmhbYw+sTQ0E8Zh/sfxWA5SNDOg
a/Bz0CacYCoRHZ5WEMCbYmFHuZ50p1weoR3316cN92Obsl1l04+33ogOt+PVibNaQzW0SfHH+iE+
lMfh1FKM5DTI4yEmolU/7k/LkFLbDPFySK+3NRKEdo3YRtoWMj+OKipZUDofKf448dT3wKQfEPO+
vS7lDyIwGjQxTHL40A9yY3jdtKCDcxkxvFKWEA9zrmxj3zJVHzReKYmAFD/to7PiG/uTONVvSlsZ
NimDX4YK1MQ2YGArXw8TvGdgoj1ztg6j5ow1Zv65c2GgSjKdL1Eu2nRKVpdHtPwMNPaBEpSHGPHz
4Xz/4LGsvyHUk78weOKb5AtKbz1xDf7ftS/pxWhlq3TUfgS5Sq7XGTtmt6XJj5HRqd9K2cT7x4Sp
Bw0a6rgDUKNDAKLfVDz1GcoHMSZaG6+QplM80GcL8lxQMCDiMBgIIx8UnpFK8srE25cwKZgTxB8p
XVAxfHski4DW+8bz1TnOQejzMwwVTlRryEwqT0SzUelAKwBYa6ua2Y7fRCOxafM6hkOBbvCK3tU2
1hOiNGiVlbnef/sa7f+HQcFuiTwO5GsCKa1euFK9TPDKKx/OauZ3wWy9x5PtLurDSXMUNRepAmi7
RZ9W+Uhj32S5mBevjM42dOxVpowZwHLUSPNvEeQPkPPX5EGEjAZF8d23cLxlTmSjJl/6VhS4ZV9z
QUraCtuiO7s1UoLIguEsm/PI8U93Nx/3ujdGenaBPrrA5yvE5422ERWt8jOQd8WEnjWmefJKj7Ak
knkyFsaatyTXojIRJOfvJzgqPe6Dyjgi2qgBP32tgi4cMBVUX9I/ER1bM2gwyyn7S7n/NKPy5ddW
ngM40AWuecq5rL/ZP6kafX7Dxv2BYlXZVGmSMmHSl+ZY5jjK6+zVL1RoRHrO4jZYdI9U/RLGNhcv
DB6F1eDfY8mbUPnMDcMaAJ1dg6wYj3+tKc7cIwZDd3+diluomQqQ0cRI5vDBI7rCgk4lDlsJPQ7o
7Pe4vrMziYmJGzFXULpI2haRiMYaWoeSTPgg1RSbdPnUwQ7yCnsVPEfwuXQEA2CYFa4fC3V46ys/
wvkSbgzctr3GmXTAw3coNcTVBDn1VV4/dY4jzuP0XbVZWo2B0G/4gLqT8to1OPwaAUe16rziu0Gf
dKfFuC61RCnPZCGV3xrlVSlf/TcVpxl2EKJipl1K3IktHK1T+IcW/pYnL4us5lFXKl4L1aPsDj3M
FJAPBPl7GdciyBfGU3bPwraRtAV7OFfjJIDdDPgradZHgHDuk2mIO4RIFay8Oim7wq41cT4PqOTH
Pf7fdqVIZ3S9j755mlff6hVe0s0QngNpAczHNMHe9skNF6wjgSxaI0M8eof+dMxBH4wc4zxCVhwr
XF8pYYqShzlBex7mC32XlIywf8vpoxAEA8x/u17lofwnzDRtsvSUdP6P1/lCXQ8X+0VG08pRaZb9
j/iLpPNa6pjJgOZG0MrPp3AvJBwtnDwzzXqAzdluTwITa9Nrvbm28N/keX1GmUcYdy19/KPQ1NIh
l0Qi0XegjQtJlzMTMnyUS5NTyKtAGn+nusct4PaBXyHvc+mHmae9Qi0AfJW4jEyv1SWUFHrwPjzj
xy90sBaCQyTXnnn/PksCTJUwTZgqpteS/lz+xyjpDNCFZT7nS9Hk78ag9f0EEOxJoHs4FayA+Oe6
R8IsxUdP4ac66S7Lg3wNL9Nf9DWlF2RKthmPiTBKcKdN4MTu94UTNN/O7aA4MWEq3eFbQp8vAgxN
Z4xaFuqzA+QNkjmhWZHebKLVtZ1ZyF7BFS7kLRRnDV7nOlKXSp45CtywrINYezDHoq2Ro/XY3mB1
YDe/f4APJVXiCOloImh1ZY6+9c5ZQjr7Sg5EVm8IhurvonvoU9W2LEk1STWZKC43HFShbjFdf+/A
YkgDTpb4M/h4lnRgc3Jgd55gaiMfOsBvD9ZWst+1xLyNq+QgLcD62A+QnUeQqM/SDeMhQwjeeKz7
4oPj6vH0RIwd4xJwi10Mou0U+7TgbN1azTAQK3ugU+mzquV/Ka+SYOb0zrG5zn1rErhUNRH493xx
WsiksHqU2ogarVA7tDTfo3cPxZ918Lo4JPp2nCpif+RsF1QDH5OGD5vtiuQklURT7xmh41hROUfF
IDLZJOmOg0yvh0Mb4KjtU1aYduHvZmhk3UhT7xWBczS4OvCxZ1TrweoYU26Xf7CrkKN+5bHzIDgy
X7eHmgk9wqk3byYMYZv23FnjlFWIxozhKnECEQ/Nd2MtuMp2IkmTo/QVyo/qQE2ntOdsTrNm2CYr
+BllJ9w+nQyegLy5BqGU2VAy0veXPowpAwVyQ/kJbl+AQyrzRTYv0g6v7jS/4sIJENYlY19fzN6x
/e7heyLIhiQpt4RukbIp8abZV2jYZH07ZWpoEp0ieFYgXGMbUm5US11Ra+XXNCB8pJ2T90lNyOom
o5CvyRle3tEiLoQyxpDify3hMZMnI42EYZPUoVjfvoIi8y3cZVL9sWWs0tC/5HYT2IsdHfemf0ph
IpLkzC3Gr0nIlWrem5SxgIAvzjZaD8OzmH5DUXt+t/gL9bmISNShpXS7NvJWUS7j/i4Jshe2BRTU
8pmZA5Rj1Iq280BbODHsU/DVqeTLSDalGBaGWkVO8gCf97KK3Iyp5ZC3MeA/cc0YbmKC1nFlIwAH
ZXYslCdLoVWzrVdwwv93S6kXULTvO24GtRZP0BturnFjhtHzEm8K71gm6mZJuYGgwBE34BEml8fO
AO0CdK76mc9nF1KAskWPPvbhWBzmsupqC1WNuuaszNbg5y38V3N/GND8eE5cTwHYqSdJuv5IEWDm
x0XCkbTdo74KETEXNyiQ0K6ODf4yYIxoYNtu+CvKhUvf5p0NuggZp8NUOq+j3IKloP/EVQj2IEFC
EhmaVcZEEaLWzZPTOkLugoib8T79gtbht4hyqfHgLOGHmzJ5Qa3y1YkiCNnyymRBRRshkEKn7I+r
i++KBnItHRFmCAwnZYGiUmV5UlFB4/yOlwwB41GdmkhflWiDsApQd8ELHGIcrkBrbUArQwdws4TJ
TFkovXQhqfb4dt4IG7JqHEoB+JZjQ7H3QtTqgDe0636wl4NwAig1rTI6BIsnHOwk88Hff8E83LiA
Qd9geddw84YZCqxFGiWMZdwpvjnTUBKnYE6Pj29c6bPWXy80gYZvDaBHSsS7rquT/1JI6izMZcuN
C6yIA6DR0RtzQOJVJtOO3owNXM4yLr7BxGRRisCc9h/gkbTIVsi/RVdX2u5nUmAJwcvcz6TNx1Tv
7pXH8eOk6edGMPadeN76Vh4uDOEJIPor0caIvi8MFCisTnEPkqn5YzIna0whpIKcWqGjsWg+oOsJ
1QeuSN7xUTw79oxXphQVJntO5TBSWivOmwrgtaCMyhQcaWB9c904VM6dA+sbbxh/2YAS+TZctK7p
AZrGEfl5LAaiCUVehsV9wbyogqZfSE9kjfeGEEY7VlagMTlUni4FCXAJeZ0M22KPQxskObQa+A1Z
xHpFkFYsRb77eFGNRAgT22NgfzGdMEymQxPITEdIOv85IS9TRQWtW0QPHm/wvnwaj9sGvPwApkhT
za9Ovx5Nqm503HwWYjPKp4FA3twummiOrRJijyZ01S/ruRPXL3BbkgAGXqGBAJBWWUer0Tv55LkE
paMGjBFvjIbIUDdWwfumybwJofzMMLJseUKTaeLExBoaqmUC+hoztu7FigE7h8JK9tW1CMaWCreC
12ohuspUs+X8dAgKP/xmcibFgvIUHEz9beDe7JQkYKqu1ojXmQ3/B76dS1HXPF8FF7ODVy5OPi84
Nl+9Dkaqz6Mr7vMTRXQ4v1mDkSww+J6KpV7eC3PRUPOoSI5ihs0N+HQYS+KEUwyKakjldIOu+z5N
1wd0Bym1GQ6u3W+EOdB623LqxF1NuZ4pkYyJjRCjEimspucSQQW3F+bqiS9lYrx8+wcVWDqqD4YH
sZqk0A8ST/QJ+msJmSYZrh0RhsuDZF/I7N2doyYDwQ+FAkXj9kZPK9+paMRHmUdco+B5mLmJ0Uob
GXSEHox1/DutII86Ls6jkRAyzV8yCDiKetq2w/1y1HXVwaw9eobHfCd7bnY3f5MYzzPmsT9XiOUz
GidvXGgCKycHYZ7FbgntzI4rAcM94ZCkgtvHy7pUubrfWSjp2NBzg9ArTjjfupH3+JkAsU/1aLTl
2PGo33g+bnIy/dj3mPCW0mI6pqIA6BBi71NqGW9DJq8qg390EU1RfV+bbikJKolGZ+BLPl2KZHm6
1x2vpae0JwOfF9BEXGTCSgH8efxAh/wvzaFIR7P7hs4/YBWllZc6xqLq1Xu67UeGqgw9jSjBwOSV
gyZrxQiQa4CJ3p+KsVqbZUyTR83qb8lf1WiaeADghXG+y/AV+UF+awzZx0NONYNpWeE91Qnc8eFB
T87KmmRO8PbAE0g1p1uKaYnmVASGqHLC8cyGv6QYQOLXhvfUmxJJumt3xkiTtBXXOTQKpPVotR49
bTfNrTAPsInTEQZ+EVTtbAj5LxNPWwd/esHwrkd6auFeZILCtm2yQo9ICqObLtlsjnuph+wL2hF/
cLt+6BWPfr7GI6EpHRcOx+tqH7khX9/fcocG18Px7bpLDSEWEz30RyaT3qtjGVgrTJ1tybrat9GE
J2dhyGwU4tbQbN1u5udsBN/x56SsCY+FNyEUJpJSiY/Nr0RXFRUdAprYjbiG8EBEWrFjwwArtj8r
2BIehGEd+25iGI6OMafPUgLTVZOGDR+QPYzd2wPJWt/T+8xyVYydBplGSju/SBTy0KijkHCC+J35
8XvpnIKIA15/nG4Ft3JVIgjsDtQFg3/wd8/CcK6WfeC4z81QKo/rr3B5XruAPCRuRBuuTh/3IS9w
hNPXXfFSaR/kJTHCXnBUOKRbRqRorpF0H8CxvyZCth3hkh8INqjHx+Vo4ruGa/7l9z+S9DM78Jtj
CgONIAsxOTJDYmRZOAAzJME3f+CIccqxaSlJ6Y5OLFSDCOnn0s8gS2FiNiWk07tAoUZQJO5wxjdG
kccEkub+quznPkU1eV0AfcZ2NULnpYnvgJ0FgEVShI0Hy2e1sStuTP85KdYJQCRxz/bLgF3Qwmqn
tbKmzVqzyL1naCnkxlpOY/os6leoirSpFCvsanGQ9To5Q2QZCLZGvoqL0qL2uCmtIH2i2LsFIs38
TzJNTlTkPyrc/PnQfobvjkeKXd4k8toWaadwGJ7PaI+z5LzVO3oxjm0SWb82S3iFstFI2BM/Ey74
suwyw4AdirMLp68bAtRIhUj+wd2JhP50sfr2pIngmpFnNfTRou0ws/g2qtBM5Z4R4d9sg3KL8i9q
U2SWDP0pNXwN0D3dA52pX8K+foBBxKAgqymsdN27bvHEvkAt5/xxYz9SHnqwCWQJRnrGK6vKqK9/
74Z8MeCVaFGHcUFimOq6jqmWYz8hWSf8p6JRYmu1ZRNJZ4CHa9U9P8umnEHop72AZao11Eyvq8Pq
USaOBh7NwcFGFIaFGnVlWXTGT4cfak2G1PHi0Mif9dU29YgtuTi+X80n0Qf5hZotTzfx7wxWDGXc
06d9Vu8aKEYRCRKFYaDnQEFgYeIVtfvCnoqttJ3oYPJHkZ9mMr45P4R8VBrB5+WlqJzu0tnOju9b
uafiFAIcCqJqLPtEvLSuNrzWuVcGmYzrd4/+n8lKPBzTiEdMdX5/p9cscCeYAQcziKb5OAlPSPp5
H5zKKC0TO+c8gZMQOb62q/fjGS21FhDa/mmG1N6zNN8tx00nljZcsGMlncZmREVv44sP01yXHUdS
fHNn2R8aVra9iQfoCeSJPr5fM0VsPrFewGcJrkbBNvC9poPXvqwFkbC6z0Dnge1hwCPTtFX5FKVW
4xk18z4Aj8IgdhhbRdfx4l+Cuu1ZI0Qv+RiwFtIo31DHjIwxznPmO+4d1Wbj9O/BijR9/YcEUYKr
O4Zr1xUNk1GHNoSKB7J9v0CleKKszA7LFvS6v1x0/EFMAyA86VvMd1QrRbM4JwzYEFJHSWYnJI+1
6DZRaXqergbVisAqS7qu9sLb9NtFHhaCvnAmEZTTJp+nrZU+mal+UNi24jQQumbDu34xiyJcoxsL
C0+uQb3Bgtl8BegzJ3oGgku8Hk7wyLXjKZYbSRrvAvd1wF86aRbouTGybuX5dRuKrcFvpVanHMvA
l0TXAPs7yp2KGk3fqoXQxD7furJnNiZKPgNH1TzsDyuec0zB9LL0VahxhM0GNq6Y+o/2NXqGcqSs
H/tP7AFQOzcD8fi93vhTGeF8qTbNvjEprnZTFDEf5Mspx5uQyXgs7tg1j0Oktdl/QEYioWDT6sjc
UuIZVAxYstVUHzCbvArunlSBLItJdc5SBRhkBiNFtTbGDmrNed0BH5n1oLRTy49HWmJjGz9nn2Ue
MifuDVVL0c486H2RU9B9MWFaOOBWXZS2x1ZvYYQF0GHaiirEA7eSg00uGmIX05tnTrCHIOJUhpIg
vezP/S+jFzhaHQtW+23boBnGLYWhuYTYqiFoO0SmU70ERez3+YGj8Pw0GFX8Xz0sjEUF3dVDaMUc
wIbgerNwTTAVrwxMkV/BCS77XLBYya9mjcgsMfKH/mkneoRCuV5Naz0FhDkFhXeCLzYn5pLjTI6o
Ys0muNN2HlZeqTX1DjI6y76ptG0OK/lqeXp+aKDT1QdsdIceR1IXaSwLTe67ymfTjn4MAVl4i5MT
Llto4ga/cDkwN6vsqKW2ra7TkY2+DOZCCZPyzlSuEd9LowM8uNrgop1LoYDPE/8pd/hayowjlOp1
XeyPIqHqUGh778/3YlN6emWtwoMwq8NJKkSOdpNe+BCu4QcLVM4YuBVsULnlKBFYffMK9dRpVy3e
VcEjtmxM5RbdFfc0xkA4+IxuKuuL83jsC8ReMM6ttGMb0bCz84kmzB5cgsd42anga95X9sP09j8A
OOFumQoifGuwIa7s4zeSuQ5IGXvGL/EiVMIOx5ZdsPp5bA1GNQzq4w1fnnpmSs0NW5tL/E0fLEW8
eLA9skfbibT+3qsIvhSAY8LEqdm9FaDB7IfixjYjLsLnxb5f7sWhggG/L6GUAUyXAm9Kl+GFv4dM
nBb1pZq2W5QFPjceOle/T9d0EbEpIbIDGcojm7OTYAd0kmVmqDmBFWezFhTEd4BX1sTgCsOEWDgW
4hvVyOZFBQ7AIG5EWg+LkD1iLATglQqPuvFFskE83mlJN1lEj3Z2VltfwNkBS7zWDAgoJRJoCWzY
1P55dKslryq0+WhnmnSZFZKDvmrdC7HtaGMBvvv6s2u/gf0jMfhsS2cAlcFs8mla2RTtbeaPSxBc
riYSkZInm0rV8nL+49r7N+wqUWEh+8ktCNdIqIYT6RVKDdyd8vRMaJf4TyStROV+rzKY62/jK0SR
qK3mMDr+zYyBwHUV1f1Q5hriga+n5CU7ykpyZpUeh851B/co99C68fEYSdn0gfFB+EvwVpYlerfn
8j/2zJ8qpKY0/sRNYYybkK1mvVnqZ1f6StSOkPwGv8IMaD5x8KoGxxoVLGNc7ruqP9KMtprDN3RF
Q5W2av6avUDtqUixRdenngi5prX3li1AZ/dw506liXK7MYc6oXrnDxPjJIKUQx9tBrD6MD54oJ5W
8MfyhI446imbWtfHvXcE6/FgUX5Teti1tH8IApxpcE419vW+/NVm8vVB5R2J2LELYk6/dy0aGOw1
uMXGf5QiTRAXErbZbrrg+PkbECrvpVsZ6DXJM+AMDuDXJlqm+/zFDwsaM7l1g0AoADimjskJuJTa
wx/92FpWK8nogDHf1d2r/hDweT5OnpfLJ9nCowt8ZG1gY9pxYsL3zstXO4YlnG+Jh9A8p/qTRNjZ
FZTxLB79el7ZM+T/B8QkQvkSlvLoEh2h0X0KtHuCXFOsnDBFKbsYisc6li1WDwYxmXeCl/c6c9gm
JG6l0CIhze5luQCdvmMukXMe8jEUxsD01fsHXUx2jCeeT5R6B0CMMMF6mEG+eOsL8DFZYYoLbI04
PRUPJP06ZMSDLOB+bHIp0SCAx2kg3qG0x+Cbdnwmlc3id9WeJEaVXXxnW9Zlv2mnlRWxvBueaZS7
5FDYaAEm416XqWFeJYqnFcf5idu/b3FkLLDF3hx1dTzpicHNCf/7YjfEp0YWuCEaU3FJYM6V/GbW
vDStDVSy2qDHxkDn31koiVTlnmOjD2zDvoTI3a+dsE57Ov5ULutelVEsf80T/sYrlAZsNwKvPCkB
mrhnZb34hUdfrEenlJqtLaSNPaUnPArgnxlGQ/XgpvNcIUdUY6fkFQEOTSgFpVFIu7pVb5Uki9ER
C9FkIVDgHD67g9dpbBLEpZ4IDQZh8ethu4oB30jcjNEu/Aa9P0y3MLY/2yoSyMI+uCb+wmI1FCLq
sIjL3vfSlI6HITFM7EyzvJ4jORbYDbkNpJE9zCQslqCZ05ImZQH+abZg8Dwlk/5lpR7y8JMuW9Hs
qW43d5zhnC/jc6tEQAS+jxlEjnbdGtP9CI6SFBoo1vhtqB+9+4f16vTDf0rXSD3c4XhuWY+2SV2y
E/0gT9YAwSkVneDlxTokpwGeiy1gFgNKeUiMgorCCg4+MQHBqPv5RpeakMg3h1PnGuy8xY3aKeVi
+wDocJ21a4d9Lr/WlO1FvXyASAB6tFP2RRt04Nxs9gepcNsvU7uoyqxknSQlCK9mpAMuMIQkSITN
QsU8z41mBXB5l9dML7RqWdYO46NEjw90cG4xf1e2Z2m6YE+MhMWm4srRgtjWDHldw7o7KDzuh147
470pMh2Yx9xC2qe6TxjPF0jzKpPMuczdZ81dbSSEAkctbrAJq303/pXg/x+l3KEBHEp7HfPICStJ
p82ZHD+1nMwUc0IO2kPsuHEDq7Dshscz2aadeJfLx0rtC0M3LLD9MfeetplkcVhmOWj/TISoOxQ+
MTRWlfRVqJTr1+MfuaMd07+Ts7bx9QtrIvZGCzhgNPAPyIEwXU/UcZDc2WDeppox+rJ9a1kQ/ejP
W23zYKqvGUSEer1/ZhFHH94uHRrrlKRa8mNeXqD3i7+kfwUluQHtjJMWNUIWT0bVj5jQ0bna87RQ
5evxtgA0kQEB5Y2hO76pUiFC3gwr+Zs1VdSw1+d/6oNihGFiC7ei2uxdBb+s+RHC5brGXJ+Je1Yh
qfqppxetQtenMVV+fpzXAzzpTDMGPhmkHg3HjA7aP20kc/gHVmY+18Szz8gN7K4D5GfpsJigcdOj
rCYR5bmwq6fM5n/bUOVPB8YkBKYPN0KV1mfi7YD17QkzuaGIbHKnfnBfgWgfc6M2FpZzFjPayxME
v2s51ZiG8M3/mwArT167eYqJGz9gs2gjtUd2gQpZ/fHmKH6Ae2C4Ei362wxHMB9ZQyCxwPG5ROOH
nRjk1pJJRSPtQCxwExPDnNT+fdrFdeAzZRLlTBpnxAK9Xg/z3H10DKmG3LCy8XFw2LzbmL5/++uo
SSItcqHTXI5+k2DrxH/33kgIlKSKuQd6jWEHYv9rM9oVrkGtFg/+y9zJHzSYkp7m6nHHFM2Gv/2D
M6NGjcia5ASwiNdj8pQ0B59hAvtmJZaZo4MffW6hxhHviuykg6+F9jFv/MYhyDC7TOoHE9BOTOSR
jIOTERWZDaIbVuuv+hf/Zqxi1uBhSNRG2JwGMTlBlzzNxBOupdaYxE8IKLkjk9NkNNUepTEHEgNa
WL/WE2VR0aSaxSE+Xabp0J+ihMjE/eX9FC7JRK0/XZT503csVs1oqf14UckdUYc+t7qswI/u6oP9
/0ZgJtL0SUX7+nvvxdFTl4lNv9UL4iKWWFL+USenXE1ojF2OrPtQcOHl7EsIUoDJUksoihDl64qg
jk5XTwXE9rmOgzJ8lyY1mTjXY2vMa9F/+IFpHaavmHrDERxcGxXVEXX2tJ0987h+kcyn9JEIuRcc
o9J+8kkIS4l/UIqFIPP+V+yNdNkwnMuuVOh6fSQortOHiZ1RmZ3L1Vn/XY3Rx+5f6hOhbRzUmGef
jlR7F7W3O147I9yKZqSaWeFZqr0MBvuoqc1On7PMvor1epCjNAmLAxRa6MhkcHbazuOTMkvfchog
d0D/AZWEbcbUvAJzIpEIID37q7EliOu4tWHqbdzjZl+gHgdfLdIQy76yIIqbd+MpvWKxRxwvIwxJ
G2FFvJGJUiHqMP1B80sC3WDoIgw+rhosQ/QPwxRMGxhW2fGdu5bBUhOAaWmgk99T6ltNauj1v0ev
Y2id+OGj79Yxz24XIaBb2xkvaYCYOq/mR+CKVVSZnk6/d93mT9mMzD3LgcPXhcwO4ByHArR+ui5d
29un06A6fBBikPn5i1FRUjuRcRRfUFUawlsAuITURYfAg+z/L/h7yeXbgSGnsN6Mxhz9vg3NdcGh
ygggRtXf/anhTq6wXEaJ7CoAv6WeHPP4qpmGtScFGxsc+21423fNdXg3NAE49zejLxCLPRZf7WKn
WAFbq2QirA+0lUkURjAXYucCV+3xHSpr+K0pYfUHVqyxXJmImzBamxrTdzID0QU8g6J167SmcdDf
MYE1/PAkiXA9Hd9ygJ7sZC4UriEZqrDaQVzqrIKwWtrWDD4Oz3Egr4xO7tcenGtZS0+BfnC6EpBB
xnpI44qmiW0fY/SZDju/ED5SUAo9+9vbQ12Zzqi3CvSfNhY0DNtIPvrrKhNNKm9SH3Y7VilaCbja
xuLlSvJeHYFHwQT7/tbBbzKspkuVjTvA8sOkj+pvme7iglawU0thgL0jT5etyJtkae/yFHzSemYw
PmQlNy/3cBNGgezmUGrsc5SOYZiCdq9PTYiBlVOBugxOb8MCRIx5rUkIp6drW+aidPjo8B4720MI
RWX6b8iTQyHSQoXe/l/CmDk4dkVDNk3lEplO5UTJo5InQCfF7vBDzJ592WzwJqV+a22TXvX8sj31
kStP3j6etQNJVh8LQnCW5zXxn9GumMdqFxOJeGaWp5PG1hXv7QOumYpJm5qClLrRpxqwNVJoLPk6
X4Cy+YZdBytraptMqAfI7PE6KA+c7T3S7i41Xo4QUbDKtHA93oSvQ/awM/dvb21/ovwE6OCriRsh
FqdtI8kTFXlLPNRuF0zlbKc89Z/nO7gY1jm029Sz4PT/f3BRuOxPRY5/ajiV209EM0zHdr7DUAcp
ggNzFH/s1naM9fRU3kJJ8Z+FQKdx7XemIzBwH2EE7xRNcsQrNcBE1OFOwroCAbYwiTk6GSDWmq6g
Oa20v9q9W98+SMnwzic2CGJiCUJ7jA/ZQDnaz+9qcTB5F4sVMuF+sn+PruzmRSEaafJ+CuRT0sSC
bhvUfjfHw4SaAqfOW2IqY0jwc4yLnwl6wwUlIF7AoCCb03ko4eRW3BHTZ4KQbYkwtoREqyN3jhyW
oUB8YjnxOVMCHASKmNEZB27DN4RWCBy7RFj/a0Dt6ssNTZGqdGYpNw4nM9ohPXQs3HenuLhN3Ex6
4wiE+J6UUAMHIwp0xNwVTjoLKkdpKo1UHUUMnw3dKF04xqCYuPi118AWDi1ltE+E6d1k9suj3F4y
3BeGmyou+GkOFceFUAB3AlX4qaRkOl8ibuZN+hSvLnIFAxhpE3o8IoGAzSDmM6itwj29Tw0BOuOc
nVf4Jn9zULCsTG0Ia4/xK29HS8QZgWD60zwg6fKSWRmfCmvsf6taWxoOLElQ2EJypywrGZ+JRK8K
6HsYksp60qxADLCLVEMBOMFByxP/DzJ54GVQVEJGPV3xIcYfVziXP9OqfBDL2K1RHsVjD8jUcd+D
sHMylzH6MK10AqwOmQL8nuOpWTHtNnSEuxoLuNBjqeRKHuhg5IQcPXOth2A/3sYMw7HkdNyXAlLZ
TuRI4t4YG6xmQKqL2YVuLuGnnt2jPq9O19LBWGyZXx+ML383sxdMaeT0Vj7CMZmrDeeQDPtJw93a
XK11Ut8batHdMdOitKly4pocEzaHpMPIe+Jt0j1jq9JSGZB0oEvwD2LrB+3Y/RRIG8AYQJF1LNGP
Xr1g/gmxyq5kX1bxwxNTK9FmJEXYacu2/cWdZSBjhh0xwPykMqJPZsPrqEvmifNmaSX6ROggULH5
/RxsivBRgHseCOoHNjmsik3uoCGhQap/VrGWpfpwcUj8VtYRCgv9pXQY77Zry2B8FjG6a7Y6ToCP
ZxiH+eFHbqHeWDXrM/ofesWDZHaXuonvaz4X/bsTV8dnMyRPSq7DVfxlqbLV6iYfSKKqW5wfmYrL
W5yUIpKyMhL3tf/RAwwvWDK4sMI3w+tmKqcrlQhznp1tGUhNwr43MVqIMTvqZ+CbyfPjWoUgqvXG
AD+RZopXe3chH44OvUoekjGIaRMtfQASsUyXLj7QFsmW72lSWmXbEdOjsFD6cLVXh5f7Qr6Y67bC
07SvAzGX68zz2beMbDILALf/rRmDWHubF7giowbm9n63WofWSOpbAR9O4FGlO6Bq9nI8/i3Urz88
wtlkJ+TlXfISys8D6lOiX2nykvzLXEwdMwJoQTsO5w/QbTupvBPhELqiqNBWK6EhE3LFukGTvkby
ZYzwK9S5H5Y5vJ8Sl7IaBTuES7jbCqoprbTWMKVle4+rnLZ9saqvi4iLP26xq2fPXXJBRR/LjHsK
zODiMZzkrNthGz90Sd56heCsMv8lfA97XOfWvShvGAHtNx5tl7V35tfppX7bhDmWFeWaDuUSdPNS
W8zW7kOu2JuXWsjHAL4y49cowjM8amvVPscRQz2+uYDjRAtGDfy+ulXXnMtkGtBofeX4Uh1iBfu/
9ZytQT0ONXo9WdSDiR9Wxzlzj8XgI2WYN1GdNBPe6fGyBbRluweQD7NYOnFiXZ16c33ltH72Qvzy
RzlrDSja1ASQXibKXMWOXuPnrLbBFuLjlJRfGx56vl0NZBwminMBIlTYWvGSS96dMBAbNslv+pGo
7gkqUQewjQUDdHk6rBeX59n4LU3BGMzB5q8rD6gN18Rny/H0h6r3+BGatQ4B+lwAhCgl3tnycEGx
I9tUPb/hxiMQWiejdNiE9y8qTeH1q9hIUT0LbWGzEhVdaVq7VwPshrGKowqdTux+mmVtnzpp/0uF
NfgCmCnVJtqd/dMcFCHqnHTg8Tt5EuXvI0gT1OhwJ3LN2vllcwKjydnXMfdDq0WAmfe7ZacxK8f6
xJ70555UIoUcRsIn+2reXluSqTissZDTvnnd5kRsd7Q/HTETilGs8/LJAI0EoPty8/vxTM6KYlLu
uPrIwIlaPF+fE+MHjNhNQtFpjaNC/dRDFTTEwwKsAW2jHbcTswdKBE18Vg120ZgzbU/48tlh8CcH
tqE0J8bWL4C07z8LlMiVKrMzyLUj9MX7uzQ/S0Cd1LZa6duJtOBuV8KPHgF/dIP4UI0MzXo3K3Mw
NhLwjzpU5MAIA7wkh3FsbVptashVo15KHQCAsb8CrOvEh/vHDz8NuOHqEAEvAzI0/M6nvkFshmAT
oiRr1+3hGIJLfu2/h8gFpVnz/H1hEF9mfHzlTW5XOeQl/F1AwwBXRhT1/w+YU7cwbeWQYS5a3CPU
KO5z2zOMZJKGiSUGWBlBzTzPXALAPZdh+J6P0cfwTvMP0+DiiTK/5Am6tb3hdiSZD0VxoHM8GRNv
1BAjH5FUG8PaLarIkuUNy3vONklKontKYf+7SV6zOYKmYBIug9XeMqNKNeE6yf4x2b+lRFEwFq2Y
toakObB5sJKn56yfYIiwdnWkLu/07FqapW+6gN3Rocbz6yngPcAkKhoAYj7piTvLkF37S+rWyBs3
Ak5o40A2E40+BV0go0kRQbV9/e9jXlNXTHPE02ff26LDv01bOBOiDnvC9DAnFE8ST3My9TsTeDsG
3zu4J29QqqN8veQwTta+xEgpO9wYlNOZ1nHeCIrAZhGsSoM5c6q6FzOWLUlIDOlennbe7LmR9/C3
o1pAyqYZBaQwLzEJI3Oubmu96rWaQEfiFiNGgSNrjxrHbKKG0VDuYCoqNJal+v/dqAE4Zhmt7Vfl
9z5Ir1q1pD6dxibVFhh2piyipusQ2A+7J1EZbnnAjhSpxb04Id+ykcRu99Qj1rAVn2Le3Oz3dNws
0Rm9a5CPiemikhOv0LMkCI70VeOh3Hv6KMtXuA9jFhbVCyqK3/BOTbQCbxuqHywPRGpUhvXjyb6r
lMqIOwpK1b+stM9x/xQXwKeE6SR6DyrealDQZoqvqyZuF7M8ief+NBRXkNWEXY3ob/FRLg869P5H
Z4ibomxwoi9bp0qnP3JCs2wgFtIHSaC0rutcbaQV7eq2uEv8TmFib6L8iQrztMdrTEF1rCXFzjho
GLOWwxmxCLNNTUTXBEcMQtGxtn52gQFPGmdS+SShdMPDtkFAkZfUNhgiQPlu6df2LoPSD1zY9zaw
T43kWaHZ999BNCzAujK932yc23QpJpAOhKPYZYlyFFNECVM38VkaTGl+p1WVvEg/QtQwDclhT5XI
jOwITLfcSxUaGyIJmC5iAbx+kycSTab2S1M+/YfFo+qkf1FDJ/qfOTAKT7AgFnAhHfA8BxVKeBXQ
BetkA3ee2IcNEYcaIRzcCIGFNLwcxEtrJZI1MNBHGTc1omgsO48TxRZ/ENk3cYoOTRumMOIpzluI
9NRS6e2lZyQB0peiiL1vp19FErb1v9DHyGah+sj8EJu+pPFmTtzE9WkCOm7iEmRxaGj+B8aIB+IW
0tQcCmgXGw/7XgUx6LNErNLj8PvShYa9viP/C7e2UQQWIY+1D/6V8lvbZocbQ0i0M/UVFcNuK2Al
8Pca2c5Z8yAZNoEJ2Q9NfHQjYIClr/k4DB+xzOe9Z8AlFczlFDn0z5BtMsVdjW8eI+WsLfZj/gEd
+0mnMkqKA4ydyqk6mCgnwQ8QVrJiU49Xth9oRThNl948dviAczMikG0/TLcnCkkj05PEs4gpAvr+
n4I2btY0FVlwtImwZmUn6DC0KvwUaOPYACZKbP+qkHa8tNJZyJPRuS8s0e/7Pnw7KJgq46qEnVBn
ZMAZP/0Y8heG/x6iTv7GqrY6Iven+K6kF61wQURE94ckqxiY4j9s9wtEWyXVsmImTuNTsfW/nx0T
ALBwD25+jT67Y6jFwL2lnFqK2z7+ct+eM2sWF1YW1ENaqg4AiAuGAe2MfgcfmvQPIh/22LgQVTea
XTp5WmJ/bv8lXnjP1ZYh8BzsSR0mOBzFH0xNQQRvWVEnUdtjVLOYTVaiueBTMAAyQRIvLk+K04Ts
NBeTJGJzhgSQXK3ylMpkoF9mUk0WF6iBDir8jVIicy5teSxYSe5BcQ6e95YvVMwETmU8PJE3iXSr
Vz5K0wb1TVunHBhlNf3IEvXCFoviKqlJ2bF83nPtC42+UC9V8HkTGV4QFTj9d6rre3hZGgxZxfbs
Te0vSa411J7wlxFBnU2Mgn9ouNoZvkYJqEUWcEbP1q71qxkn3eBjUt5uiwDST8Wz6ThUmWbXwK1z
0Oa+W+Gl/wKJXbRF4wokFQoppcrc+xZBW50ugXvzBNHUf7/KdiIcSVxjacfi8zCMIOeQRcXBQrhx
MYlYWiEyWVjOYlR5ePj7cP6J8RuDr3XBxNSpmUip3iI9kWGOwpCV2iZy+P2y80YA4kCyNIjrMIHf
BxlIQLAnsAQlKjF+X7I+Fs2SHEKHsfrGBx2G7T+ffwUpKXIcjWMN8zZ3ZIgLlvoAn9YYYjrXc1T6
p4SA2b/fyr5V/i3c/RPOw7nW6T7R+PUPS7ZhZ8QL9CXf8/BxxDJKILmBlIp2EjUcQjA66eQOFs4C
7KqsrXEhnuY4b9A25YMh8QemjMW7G4B4RO6VtMWDI5L3yKgF12dsBequCaHadsMYUEJSlTmpQ8lE
VJTSJdDeH/HyziECB2dXbRYacr6poA7/HAJmcLApZi4v4Pcr1vzaT/phXIKyieVFmRLQzNGjHTOO
xNPRu1h2X+FxCr/XcNuPVl/FlOGPTex7UkKfuAFYyZvM/OABeQqy1JSkXMIxLLsap/0XNun272Pg
zno5ybOtsdZsl98RqYid+oxvLEH3spEOlY9XBYnSMz9AhS+rp/2Oi+la1nq3gpOQOknqaCsd7Fwm
SDE9Rd+EBYgyvYFGqxksl2hir3rVyNIOPJJwZNpPRRxrL+YzUfcDeX6ejSnyH7RtOPICV6ldo0jX
1hkQRLdcfoeE96s7D+AhcAz35enNQ6cCQMuY5Ci7P2DCOumvyfA3HSGs0gYnG5offoWDKuZnfAUk
35BxGRytG37n0DreGu3hoX6jCvKNrirrvLjDJrChBVm0WDUHF9v/2fkfSPxeoBg/A8135GMbSLEy
VF4Zojs7eskkV9rtStvDZmEcbCfjH80RXQSCz+GTSYBzfBvtlL4XN1x9EDt2GhBOTZbA2Q+9/8gP
BXBM3xEmW3TIepX6eu7LuXvWTbvWhcfzbIvxFYBrNvBsq0rmM3oerAVz75w/Le4XBk1W8XH73ktV
lVA9BqU7UJSpv4Z1Cwox68mqOrd5klS0HvF6ccBnTcNB5tbXUePAtSIhcPL7DnydYUlPiHFbj62I
YGPkeX4b5uc79haRrfuPLgSwxx/iIo4bpZVdhLRtNEVe1xITCQefiIwT+MKxY5dSkINsQvuNWrqj
JyU0O/B9rhgVYFqG9rzmzZNxHPppCcI32xxVOZlk3fHF0Hig3ghKtCmx8oQARYLQeRti3pr6DpuV
JA2g4+5Dh8hwWSTqFazf1/KIlFMhlRijaR0pt/NoGpr+kjaqu9YfjldjO6sX3pTRUf8HU2Smz9wy
iFPERrK7Ia1RqNsZzqSzUax5ii6KPg6Mri7qXIU6xzsU6VR4PuTyslN4f9X0VU/7rtLfgey8Yzkd
b6wl3ejVhnvvqbc8iCXlnweGoBoaMxBW9FqPKi1dpA257xoqtrOCI6C/MYgPL9C5K6AVtp37Ex41
sIsX+y2mrGXl6em2HeZn3II6lYVwzqUdXgio0xB50oTuippuPC0QGbXcT4m3xc890J0QoT5Dnvyd
PHOte4yvlrQGDlAavW8LHRu8+FYi4Ny8VxaeQu2zBNwudmICclxtTK1JW5QuP+g1kGkegUaF0OgX
rwMSvCVpy5VofBzLDU3fuy+BEcmAWM9iubqB3a4va4zwdM4lWu7MM1GUxhtt3nl3Z7dGCql9w3rc
DDrA79RHbquR5J1tmenE0rigFaClZO2EkNOouCW+eLOfVBMRLJd0QTuPV3Cwqino28e8M19FSpOk
Aq140OJnahxnUitOoGEtttV7nyZgp+JiXitHlgjXSf7aZkFqwH0xHUXBqbstS8Wr628T3GjNAgna
Zj0BFxWNdjjvjK8mDgtqRMccBbn8yntrfXuY+0QtZxByv1NMPLOP+/iHNX3umRqnFIQOdGF8Wso3
214u98PQqjQaAUYzNkwhn6w7OrtVIHgHf6iI7DdYImdtSJOzWOo27jpkxAM3vX3BlPj3sTB45Ak7
rtyVekiF/hS/OSabm01ioPRjUCEkVP2vran1GlCyECZIyE6PW7zu5G0yKYbZRtc0xekvrXQZbsNc
Gu5pJtSdei2F0vPDuLNeKgLzVm0iyNfKlv6LlAOrKfdUiSnBrRY1DdBXJuU2DkNpMC1HagGbch4p
XWXoXi7ljWcCL4qa48V6/b/T36rLQ0apZWP4nK6tl8FmDc+lMdn++iN5SjqAe8OAXOo+nj+oAUMz
ezWO+xLE5FFseBHxTD0rdG+uOjo54j6kA5CiGJV57PieyxT5KjicopWv7gzIOGNjPQOCxvA+QV+a
sDJUSRaCEv3ZD/L61TcuXHzVD76xzdxHiiRR63NA29/wjX51WtMUGCXj83frWvqplQMDi3BP5qXV
8LHLInDEtZ7sxOptUf2SqlwOmVdr6CLU5ZaGfB8zBQBT4phjm7lzB0DvHeYtDuoZZcDbbxTNpG3M
cNNHVt7nHjXkc0ZZ/6ISsxd6+EmUT9kFcGrVYCSCK4o055wNPWg3VZh6VE1/v6Z4B8pCaloXNlGN
zrePaK7so7Vtsa+CxiLhlfkPtI3Rgt+Gt5E+ANValZl8HPAc+y5nRHJ3AkCphpKU64L4bqXFalOO
Yxyzq0qVSqbz7QOaG4NWMbmWrht+Y9nU6gUe9HsJmbdnRklryQgLyfGckzNko4T2WO9OQ9laoAGw
8t01ChOAj1L/EzTPMxWpgoTmxwzkQEQsnlL3j5ppU+79e0oFZxJNw6pxZUE82E2nh10cVRI/GjaO
MxaRLitiDBrQHBxyDvCZ3b6A8aKuReP0wloI12twtUNTiUkX3DK8qc2HdekCForEtzcP0++LNwi7
rQlT/deKvWuB99jGz6Y+2cKBG3qyaf7sQdzgcwlHxP/+ntD9xHyUQ9XMlI3uari7Gji2gcr3p+Ha
QG5gI6NR9Rtn7/BGTkjxNsfBJ+/Eh+iAtnWY8tTTHd3ioGo2h9Cd4VBqRbohd2gT3Xa6PHG4T/Rh
RSoF1xuiXcBm8TRsHmZcNpyBNNu0F7OUQsWXjqPpZsZsDGm+2yLqg45mggOifQ9COjuRuyDF9Y5T
n2LEa774B1Dg98VHeIqV2xEkk5/aySG0+3Pv4Wv4egEJ58PLHwLw2m4vwtN/lyb3LPXGkJkRWp8U
1Q09vPrkMuOmuypvK36ljwpIOx6ggBO7htMnCuSGe5NGd0/VnJF7idHsQf13z6eecpLXYY1dFnGh
2xHBTWr9hmlK8TfwiKUIhZ3Nw17RmfSMQFN0jYp161ZvV69Uqj9hj9FZiJ1QIFv20lw+bBXPwJkI
bElbCmbufrg65CjGlC4IrkMdbEzNDHZRzpJOfdfFyyuL2t9SNKeKSuzSxXicYsDn9n7q9o2pJJRx
EmYFErecvTIfqWcZTynmSx/E+k8h6V1pLNGpdLQqmhORh6I3w7IqX1lvlPwVUOK/Bh5AdjbdsTiS
cR9Hl1awp2+ll9/U/TDs/Cq2JD1BgNEnVEdhWsZ+i+oEJlAfbIR8f7HtGzPl1/M809q4oKFv6Yrt
mVxCmjdTC3C/6NhpcU9VTp7FXX53cvWXbuYkNviA+8S9+fQa1MiCtYVGQqlfU9WZpe6xB7Z6blrU
9gsDajEUSuDT0lvr/uWpKWERegCmNgjtqrXf46xzNEoPbGhL4VHQaPR20cSeh9Spqe8fAeOfPLbU
sa1OyotRjPFs6m30kEljonasArDkAXEh/rvnH7/+3a2VUSIOTaKwORFcx6mlhXZc2Xir+NXFPZeJ
JlE6ObeOCuKyMEHQxeZD72Ynv3ejex69jSRr8Cb9tryNg8CKI01yi/NzzV37iM5U5RiA9xi6v7rI
1EhD83r2SXgRPyYy59Z9yIgXnYsnINXdQkqe2HZ9VDRbToaViNAzYmMaVam0pAXX85fbHQo/cY2v
pNXcta+ELJMTgKpNxY2Wfq6SQZroV9TnZ/NyrvodbUjFX2EYcjJarseEQVnvzFcS65D42fmu59HP
zoFGj/IEuoMKP/iib9XAWjXQNHdnWVnUsachiH+M0REBWDXErKzNrx5bcrmLnWCAArhGRK67a9YP
ofhzobstF2NhaT2Go9ZaS1buZIAMruLXDvMvWMB45mviZ3KdhJXle34jxb69QpcIkzhj/1sftCFC
MB6/zjf6f3ITlDp0q03WsHnhtB6r3weGrCQz0nZLmvyHpHco+i/VJ44uVqXzBoC1Fevsy8ETu3pu
14rl6alF4ysJMY1p+RN11Kol3Vxt3GQxDcPTDQ8sWfNupMnCTYXldVtd/+ghSUjCxnx8PSo6eiTy
H7UbG8oNmgsp2pE4aggVduXnSeaCg8mpVlWflF0phNO1IaGDxp0aUAQdc4rd34+SC+D/w8VWc70S
m1yDTb6ZW8WeZrYIiGQ7LnVKXO19d7NgvHVg1KxfkfBLpdDuPs/UVugaBQf50vcjfuB6DPTw5hnK
/IG72WEUuUdBXsTWGAey7TzsAUYXPROreiqkycDejqjgYib9Pi9t2bLfLUJLL9+9kdkbfaKX4f6C
B1Cw2PypNcGn/9cMDs8/Dces2hdWBl+BuT500Im/8u96Sv7toa34eD2/mbh9GZuXIGPnLtP1vuDx
2ll5V6AbcyCIOMqA29TyyG+3c9+5QNu1XzGCAi7ptlnGIHl7ua5Syow/+OPsiEJ3CXUXeja6VQxp
Ovk41Rqi3thHRBgWQc/vo5MKDUJM+4I9EW+GWKdtzRmYgWwdhjF93rTjhILbR042ZdAW6PoduWe2
CaDY75SOQDpUkSJOY15gj3u3rXiwb7fdcr7olxLDhfCIKCnvNHqR6Q6Wv10NLzrZl8pX+Pcbm01p
K1pp3kwy6LplU0ZSfYQywwDGtEk9tavRJtOncTT2ESc0bbZ6LZjz0Cr3wj3gORQeoQOvD1Ij2qFx
u1WpU4HgXYdW+YQntKF6hgxRy5BtGBogYyi79SH4LZVL4PpxYZeVTHKJZEknMp+SkYb48Mm0/dsT
EpcxvN740iIh2/mXSNs+t0HzqI0IfdxqgZsSrfFU/hAiYqRpuONJ0/np/Ux0lkw89cbDBp1F0eSx
nZKOHHqS6IX2hMFSLPnEqQFdjUL1fNpq0BKfJMfLtytuEDkbO9mpEsbfxokZgJTFk3dSNcu2Yfga
6i7K3X0BFSiToa8IWDwTeJohZ+ArPkbA47DYIcbRCfwrTlU/oue87VJtWkRMiLU2Q0UVmvCINQnI
1OIgVkC7rTipnVruEC/8ingYqY2QR855NReSzFTDlv1F4zEtPemSMT4dbkYbAFSdPa8TOVKZi71j
G9L/9abFrQAtezEI0eigwvk7hSQhltl70fDKe77DYDbqlJKsz5F23xny9QPO3hW7qkhHHG9hpQU7
RMcfzB6sxzBZKgs8EFodrR48lOIbABvCBwNwd6+Ds06WUXONzd37mFaV/HDjRTtm4qU8b1+eSOmJ
ckYQaoruNIDe1D+N4SrCp+DfBMDLE1jiWeV9Qa7AR8XQWbHb8fgKlPHIxfMIxu2a6F6QoeYamt6u
1V/bHEpwvEoqGnsSlCiteKy9x47oSx8ExWGUvlt9nlufugXkNGrIg5ooGpecmmZOCvvWsIYUmIBX
x1qb53Q+0/FHI/xZMubzJE1Hk1bqdrRbpksfvxI1o59ieUrJCkydL/mLDuEUO5DvmKpZDjJcENU+
j6N4pmfJACtuspzfkzSmfDAL2W8P0yufeOyCaVPzKKZYYxkF6r4JxYFPIWiha8RO58hy6dakZ0Ek
dGsXL2x3tt4AjatD8qANGDnS7h3EKtGMoGUO0PcXtlhsHmpmuXxhLXmH9uSOEmrhMLAFdZYOo/Y/
T0A9sZOQSBSUVpkb05qLEecOMl3rTAOZF5cY7r/i80ic0uLxBF/9DOXxY5yWlP+/ALl1gJad6oot
LGlg3K1KtHqgerkDN67K1c1mTV7cKTsTMpqUKlBbVLoxkUJY/u3Si2ew+hg6OuJnJwnU7psEbuyi
QsVVD+aNA9ADEoC87BVajh8zeH8AwpWnNS7Am5GMzAx+ksQcm2JFCVATTR7JGlYemIHMMQQ3l5mA
snNOSvsphqbk2/PWhZ+XhjwmciDMs0e4blhP5Qfcs+WprxWzPoChESh2gf3VlM/jCrmvzrPPVy8l
Q7enV27106ehpWLsYrbOXbwxrB8lpX9AzvGflIe13wo8BNvDFpfFNHoQ5CSJ+QlkHJ38CVMFPp74
xZ7KIkcJCNTxfDwCmf6PXlBnLwla7wWxkCBSKGzFWdKubGMhKq89bfejtGgyfHdN4Ed7Imdh8qFJ
QY22zUZhmrdPoID4j3b3aui80+CU+NVmY0c050BZ6FF1MxMSlN6Osh6jZnaoHzwHJOnAAPLh3txk
DU1ejojfaHO0NGgOopVD72hNRA8HI6E2dtQ2T4yJRBoBL6PfAX2glwG6dosia2vLgzBmErsdXUTe
/OAuolmNggOHhraYllhei+1BShGXq6wRTpE1/SZpukCMyPehUvKDT+JQWeoTF3mss0p0bbqbeMhf
m7I5t66VSeYuZQmWJoP7pgSMxlA6R87qpCCbprlx526+6KU9HlvuxirRNhFHRtV40jguBBRriluS
luYwgsoIn0EPjZcswIrlAA/teULac9bcVIlEq5xn6+vYI6N5L74YrOTAJo9gksmKDlcnQ90Zl2K6
fMESM0Onx9D3IesSoLQUIQX0EiuTRIJjIsqFwZcNYT0SslGRxl93Dzvw6HkWouerKRlU1ioVPCx4
EtzoXR7/GKqdjfkjlgOUFL4ry7rY5ZhU7+7MbtR2TbRnqtgZ5ameGTRO6fiTGrtExi0eC5Lv5vgB
wfKNXQARiLHmYoa5Mkr6t2//QZx/2lSieR+/FpCcgQSiDBoFtFLW5Kskla6yCD7snvDPwaoPFdmJ
5uiTW/YWY9Ytale3+aFgo+v+Hbyld1+JNmxuRaawyn17ytScbO92yDTl+fzN8I3ut9fso+tWGdVz
SLb0FZQyr18kV/E84Dh4nwYAHwxDIuKrTBVhb4FjIeYuLT7AjYYMTzVJUbtWnXpse9E35l4qUyS9
Tl0cQ+nlMVU5HaGhCsMZOoZ0yZOyjQScWN4HSKUH6ZWjCA/xxVk1K14PVZ0Lm7OfMHNJQF+5vtYw
lcEXW0fpevMJ2AW0S2cIyuVH2RrrRwZlz5eSagj8OOS9Wzz4/Lg/y6driVPOubaYihR2O2MkZPrG
oLhqihP+l/jFBZOKdCRRPtTqm2R+RAhL8SpbciEcJ57gJKNoh5JH+x2FPqXF3OHfSHqGPJU4Eu2b
S2DhzEKC7KenrnNBNDTYOGull7jXnNvgSQJRYu3ora25KHDMQT2E4oxo5sRTeSBUipysm2HCcjKK
RECOo90f/sWYrZlv6pgYIWUWf3I99K9uDi9QXYCfJOUiw5acFbj4+ChKYYEyVrxiVw1aQ1EUKimD
JDliW/52L9fNmcwP3nMG5fXwGZI1+X5WRGfI09QXVrkZ6lq9AfV1TebTc4e5+881J6WrE8ZuJ4pX
0YIj1gurGgCHk/sWN/WB1cFkROSywFeg380e8pq2FC4DjMHQ/NuYlyOikQE4jYfIM+mhmj7hEvJ0
4v0jsKcuw3XEwRyaWAzeG50GAoO1ZRyYZgxdbND6fKysP3XVGa8ZD/XBvv52f6Aj2GWNLZg0SDYP
GoZn8dLMrJ4f2iBoAj3McvYgOg4/ilch+VLwkR9Wy+P3nd/1e07kXhJ3rMfba1dOjfPAdx8HgmPQ
JS+qXA6ponyMUiIB6XaYg7N4b/PehxukjEfdTXRie1/thXRw+XCriF8ot8cDNVVVSk9osPPHw2OZ
h+nPT9rsKlT959y/kvzbARrAkWA4dS8pgaIjyL7UBI8UxasaJr0aVR20uqYCE3sS+d5GQ8mPgT5s
qFmnmLMA5tKRSHFMzYjKsoJXXqEYWj/XglEwT7eTljJlfcYqbFQXwP9Hk5XYP7/piFUdK+D8IUxx
saMJ0++LF/Si9QMRXXpLd47o46DcJ+jAKKS5joFVVG4EcUDN3gr9K8919pj3+WDq/INPXh6YpFaS
x1mRfs5u4WTZThQFCB5SHh9hdu6EaT5CFkikaPKSn7+0kgK6Bdl1/Xsf0HNQoWfmgP7G0ldhF806
Y99lr697oqhP1GF4h7/d59XzQ4rJvaZPSmeRIfb/TepbVmFNgjJvoYcBB7rSpl3k/MWRzp5aWpth
Vgok1FDBR5rVTzxAB8+lYU+3Rvd7s6H/gOGMp0WCqyd1t5dvttTwcwlcSz1MApneDe8BSaj/ERrU
3nAcLFonF+9p8ouKHgNfOfHFQpTi3origRBqX3ScGRXM71AN8JHEcygrqCnvdV5oGv3CkR/8ulu0
E3a8ngUz/4M9ZyEIgNZy2+y19G2t71Sj+H+is/jLIlnSiPcRRJv49FFyRKO9bHS9uCE3LV4U3Lzw
G6fRpXszgTpHIrlPjoEGEhssaOyPnoU+kS3qhY9o8G8FaONynN/Z4yLlnpbczkbHiAN6WIS7LC3m
pDquF6IbIOn7u5IdQutkjzjP4a2wOTly8YU4wZ5IeTZRT35OC49EmescGZy/FrSaOA6LY8d24DZZ
Acm2WM/+gX5+j8tF75327O9kCGwFHNi9XHn1nq0y5TKbNSLfbWDW3/PLtYpI+fVQS2eYHgA/bUmq
E5XRNY9uggeTvH4FY9hn5uckA5KOJ9ZmAh4hy6xUmcXkGvsTtipwVDik0njbkXoQAIHTZMOC5Jy/
GfHMp2edlSeoabMc10M7NBUoSxi6nhqdy48tsHYAjt25OAW4dWVHz02yV+ODAMMwQxUWoQwFftk5
tRPM9e+3TdQruIyIGi8veY+zsB2s9KtYF4MoJoBGfQNJQHialEbG/w4nMaZ/IVqYq0UEKgE2M3uc
NTX6tDelDtlEANJ+moGCcyWUh/WC7Xh97bYbug3v6wQh7Ukay8AIi5t3vEf5e2tFzBEQH+FCtxRA
pONSYxwy7d8kehrYFBPzVHaMWY8GYFKtSo1Z7992QUBXq8M0i1nR5mdM7jDK8Lq7ikPVn+DlroE6
JkErnqxNkEVy+n8Wx+n+00YsO8J+n+6qft8VGyB5H4rdrjzA8CumfQnRtFvn2V9VqF2gnc/7vjeq
GCoKSf4dCBUgCxqszXi25qXJ8Yfg+L8yVq+p2sljTPIv9x6dOxhhviKAus0b0xbwygLR+1c5weAJ
dsYb+2V/bbA44WS1BeMJqex+0dTFavPw7nsxvp9OABRaRVPLU8Hxp5vPAFw7PP3XOfMdHfw0ZBwb
GBb/TE5eHaoIOnDT0cQEsn68bcVL/puRmj+8dnMDDwlII5pFN8mw7qaOoz1RVqOWEn2WUoprIgci
N+Nz10TdFMSensOt/hQcW7AwQHcQ+34XOqHgNU+3iHDKzhucVxbZEZELlF2VWLfAWoayCUCGw9ZR
bv0z1OTIhz2uQLodY+OGoz5bc4bcZlnkwUBXVsDrELvm9BXkUnq+rsIUjj1o68gocaWw4rsXnSwv
YaG7eb2hKyxsGhuPZpjJsGCAYAJ4XXorwX1FTEvbrUAtzQpzCiQrocIbfmZ7wcnR/Dnv0h0Thr34
TDIIMkC23YVnZ1gIVoSBMzu+qohaeEK3f+j00ZgK7a8LWG7oO5KWlLCBjMidK/YFWs3fZzfVLRfI
mOuK/vEqSfgaxTVEAdJVaJpNU2vGgwT0OyzjE+VkgfbCZKtVrbLK33RaNjn00SoikFgmSzdqz6sx
FBnvlYD4OR6SkRSGGO9BbyzKmpg1bAuq/fp5iXOJQprRosyFzXEZx191QOwuD7Ue5uMDO6wDZU4O
e+DMk8/TwgMOFamN5VCGyPWx9yJCAKrnrHRNHUW/Xh1Cjq8sgjfzL5FUEyAvAKaVvhSZLyvsfMh4
TBiNkdCVeBpeWDl6TOD6fxzW7RQ50L91wlmKtJTs8/Mhuib5Ky197Z2730p2yD0X4LWrsJuttqMG
ZyE8LUDxoorz149y7otmOy//EZifc3pKBQeNeJza5GPK3rfKWMyJOi++NYhaee60dA4YJv+jy6XN
RiTmF59ceZy0wb/wYtEj046cLpl/4mpiwvZaZRL+dtEtZLX5hOnHtdvIqn54ugFE4KX/GXRCA/iq
tutoH6+XVAEctSr9xYeMRXxJkmxhri8L5UcXSXGEvq41RYjgBgm/9LyJ4BxgLDSEZCh7oAHRNc6V
Rfad476HyKps3Zdy1umGerIAJjO0Vb1wbZtGz7v3MNmo6mN1X9XNu2KqS35qqZuXh5WHvKQ65T0B
b4DxXetl0ZTMCo3zObmfU1FiM/krORBZFD/snEIbQH/8H2fissrsAYp3/UcKuO8TScgnWj49j3QN
3t+QNzKTG4eZEDRJO66c30hwnN4xBC3LKmQd5bt0VvxFRMQNL0sJATZ5EQFobsFWZjPVOaI+emUZ
HQNtbKxl4+OihPvd4GL7RV7zrVFjxNt0f3xVgOvvKjb2uFpYZaf8uDIa+rj54QlYwT9SAktr1c+H
RnQZItsfBiUSWuVsja0VJRkvvupJ1GZWEiqSgSVGSERJPdb0gpVccAQaXLHTwpeX+IHhn1q1CrrH
nUjt9uDCcJDI96VLjSE2TKvwVfosVG2zWnbZZkx9z/tCPC3M8sy+Yte+S2x0s+6UoOcWkY0ScWMR
IF912X1gxMABmAOSLQaN4F8I4MBgScx/PBaaZt82O5OrrgdSd1PJssTSm7Ris8fhq2VKl7ds9Yli
D6JKfrN1RKcnVUSOVqHlisGUSKCc4qUg86KKRDVCiiTkXlilzFEGqzBGtWy1lA1tlCPZqwApepaS
JGr/4EeaipzpVbRKYXb0sep1YCOZgiBm5eI28rvfaWIik/wzfanf7cMp7kOBCfauA7ILxGjfTNKT
oPWHPKe3RYBWACVlEIUwVupuEMlT5GmDOgnzNSaGpLG0jIdA7KWYeJe5YcrKk+tXzeY6SUqgMY4I
n03v3s656rk8tnxHLNnNmIHZtpGuvrlLbG6fZBiZpd9190jKbVCwQyDo8Jwz6tyuJ6TyodJOqcTZ
acUeX4SxF+XeQ349CLf0ZOhjqewTtXTss+Cb1YUgDLxdJ02cx/pc86/W328fgU54MQxIeeFZLE2u
xBzmPovk046PJsT5ExT+1MrxX5COJ/rNTDx4Ni/c4D00pfKW64jLxiWlY2qgsyWcOez2NRSJgJ8I
19/LGICI3JSlWozw/I1TF2ajgVBmh+jNY4mMX1t9rVy05ydFkVSyOsNemEl2QrqvaWv+p/CXShwr
1qSjHzowHZTFPH2oFl3JFncooDVgXuuAQEYT3w+JJ+suwfilfHkD4sHeWhjc2aw9vNSWtOqR2Al+
tXzZLznlqIUaanjyBrLWNCPaiKu24PPNbRnv3RhkYT/dTThJLuixdr17mK9ySNRyW6emgLADq6Uh
usz1HLL0aVnDWIoPYVgkW3/GslrjcAXlARG8tZHL98ulAasJVnKtZ+rKCdi//lUQqKPDLKBVhjh3
FeXx7NQBMy5VSW4aFZrEmrH/467YqW278t3SF+Smt/sSVmD9JmI6j+VCNoeWtIPmDlwM0CXdi/Qz
FCWN8JQAQdH7R3eCFH8jtokZBYXCn/BJqCBXQ5MfEtsUnb/Dw16YlJuN3yVWFxzr3Mainp7rr443
YuYcpVk7p3M6t/CdLHNuXJpnTnRnsIngmSz/kH71BZtq9iMjYC6xW4hdPiJpXojR3ZKRY7+DLRbb
NSVlBBgN2Hkj2qbUD1bhnDPRo7CROyzAV8p0VbUt28v3OSz6xtgC/YACDiy8PpkVKUC5P0yT16yB
2Wc9uWFrR9RwlS9sxminIpsPhOOYhWjxtIlHd5FnqeLsuKC/bDG5rI76VhIW06+GZgqsm2jzL1zj
zrQoVGjx9sdZgZDFI035O+XRIf8zLuVlZ6ZKybwKoyej4TPZ8eEF+rVpRPefsl2nBSzoiGoTR93v
Gq5L1Zu5jAKEP0VClDkyzmQ/fd1r6GrDPtd8jlQ1Aa3JKoMyxaC4FIAskCJhSa3emFUQf+pitp3u
o4rrNomAUJunhZg0kRZ4uLjNf9jKAGI3Al8M56owowSQPn+E40h7BbNabYBFPW1N2hql25QZImI5
UEdStQamZF4h7Ua4ti2gn6msuyLLksJayVxUamEBIxBo/pw6l2Jt5eJbWx6uJfb50RTqAc/u6D5F
/8brfBnum5weQ1jfddIApJ1m3SOtIiRLBEFnfqoKrhrUu/IpjjANKJaPZSXKf8J5bnpj5VtLbTAv
Go0Vqls8Vqgz3KdO8mhUlO+hXySL3ijyCAvKzxAT7J7sqEEFsn0BiKTd32wKDa78IXjA4NoWdukw
PAuhjhOehIrQxWbBE+7aNQwf+D+rSgqotIp5fi0vLlgcMLnto4aFIJKsu3DPSITSJwmI9ehVuXDF
PeCBigxsrADcofNfMHeZTGcZsFUse8dnap52rSj9s1GY54qPmjiLkAM00UMCQ9+FZwXxA6pqQ7fT
4C44+CTYlzGXWU+wghnPxuvjo/AZro1GsI7WFUMKmZc1SC4itoA7XotcuUR9ZL8I1N4/jyBzzfFR
DDB916x11BPRZ3cqm5ldc2B+ajRwHHuAd/sfGHWHTt28+xQa6VKLl5eALV5vpGVnI1/Pn32NKECJ
G8GHvFjbobPvEk63nuNPt0K4qw6CQBkUj0yp7cPmbq0g8+D4ZYLbfbpQCPXuDhydGbahh1bKe3Ci
Ct5+NW30jkf+YWyf6h0Yq07JlvmMolWgiEgdfSLEvXlhMgopKD7rKuQ6HFIcRNypzdgXTxq+Gc6A
u+6K6tNUZypzJXqszI7vCdwNsx/CnDV7pBwEAldpi0jB1CfEzvtZjk3D2FZfjxYE+dk4NDqS/Qww
cLVvPDPSE20hbo5ZP/+Owti944t6ygwExu5VJ5pZV8IL+WKgUq+CJdGcPdBX6HkW/hXsaooYWyAC
krm8EnFpU+oIIf+B+6IIe4HDuhXbIlJKJS5CelwD2uBlHsQ7oYIlm7SOlJyl3Iv5t8xXEE3W+66U
f3lKu2liIwT+GVb6PE3vzwwk0glk/Ph/82NUk4vpY2D40nI0oQEXkoPkHSnftHz4DXsBFKt6UBs4
a+6QWjAIbS5DME4bzqZHa0VSVV1nAYiUUsj8SBwE+vXtee3laY83RoWzRESb6JSY/OdLhkrsGDEU
3UuB2i1MGU8U/ygQRNQwac0+ob+e9DTmB9dxTL2/C6k0Np3vs5ocsuvE6goIjI8L2Sko0Eqre/BN
mM/eYXoucKmNkDdOZhogNCcx6NjkY494gn0Gdxc2kRTNoquvJE4RtFR/19BPFHZzmOyOrAU/ENVK
oHcU/wHTrDYRIU99iO9MEavWmCpx/W7N0OsV/XfPE/oNY+dfRaZ8aU7jXhaZlS6EwVYivx16G6cb
/ijxvh5VahyUe825ZjE/ns/WAaoSqrailz5UDi5vo41CjZtERHiujRJF4MmSOKxVkqph66+SifQ+
kEBktye8BTehsjLo6ns86DyU8j+TVMor0uC2IdBP2s1/G+Vwx0kvexbcTB1RJXXJuBTQieoFdRbM
NzAEt249aD1aYr6Ra9oLThnhHHEuz8pbYS3q7IFkGAAz3aW2NSc+aw5Wj3T5n80rflOGBLBZA4Qd
BnBaB73clatJiWr/i8tlNF49ZOrhY+MXNDKJwTWwPXy8UmFNZ+36RjDLquduArQd5Okn+wsH06rk
g8RivBrDF35A3ZuAUZiEtkxjtShFDdKUe+biyPRzrk7DoyMY0rfc1TnMOlAg2g9nJACfqr8nt5Vx
DI8DM51gvXg3m86WkRL0C/G7PdY7oSiNSz2G80kcVmWXy+YbFS2K7PXXnxRP3k+Suq8igRVupFvB
pYaNyAY10Q0bSSA19g3CWW9Enaha2OxQpP3+DGQoEn5RntKaDdiIOnxqz6Rx311kSMGZ114Zq62N
j0fnqFigGNp9/sPqjobWJ8Hed0MXyQlEylYwfiuPUzt6zazJMQdOnnlWthdu+pd4GpQ6sY/FJc4E
Iwawl47dzAQ9ZqtVYmXKJy73jGwrgn4nFl/vArhOpJt/Bx0Oc31MFfzZ3dc0RUz8hceTJu6H/2sg
izvvQvovMA37d5XhvxgFAeGOZdiXu9VWJ/CPAz6ZAGkDI6D7yV30d9q6g/8bIkk0CVKoaglee/SI
jZ0JNR9Yb9NECiTHHZAI+2d5oQYiC5x+wuwY4M8yKgM69yMrgO1qi64L93sytlJd6iCwQHkpi9h4
zXY6b8qDnPZqWeVQ+3UTtYCtpKEc0gZJjZJYWz4US0l42T74ZrXIrvfHt5Hejfvf+tN6pD+zLZw8
UO+Lh+cDh0zRQj29NuVld/HTwvaZTTpWHR78IRzc7QWxXajZ0azun+fIA574wkl7QJ0zbv3eg+46
CtTolDO7NqzfCCghyxq5uitbuddUW1O3veHe4u/wP5lQAcVZBtH2XdW3zpQdCO/DJ7mWFbiiEQiJ
Ftw8lIFWC8D5M6/hN2midS72InBP7fAq+L/+5z8sG2/unUHHhl8EkJwp3G/8yheYZVShpTGkPajl
t4UBC3PrX8UsF4WQO6b3O2vFNsqf3T+1JZ6dptrww7TbPCuFNPMrJt1fvxu/PeUPzzI23liYX5VR
fJe/N5wOVW/5iYa2fwBQrYzQJUv6ED0BFyjlhZhTylvYA2olOYze+Xb0PRjnDDsl1DjSj8167cow
6LGyhhBaIcpj8mvmWpzgAIBERbE6qbMXU5dZze9wSDhRdTZiXIhyfxojO6AaLnWY2n+uMMYGdNZi
NOA8rIN5MZshd6UeY6W3jMCP8tW6I65VVDDGDxNfNpy7bpKlidT5MntDVwU0Yd1DBg9qgkGtUr6L
15g+8VFnYBiQrn7lSps4bRBWrspjJhgdf6OY/8eVzI9Sa12czdEbBw/aWjDJ9gHdyAiyAfHJCcpR
K5vcJ1unwFquujqWw3LlG0X7ZqWgfA0YRPgT0rJ2w/VMZMG4uZwNHW9X0f4T7OZIjsGhY2pPDLki
0fYxBQ3lcd4o5cFVlmY8pLPfQbMQcH87RjfV3Xc10YWj5t1GhGFqzndb+qhEpw8i7TyTwYqbjU4V
9aHop1Jp1QZ5xPQ0GRd2TDjgO3fJlHpx+SRP6I26qJIMgjYt9RcPqS4wKwmmFq/t82vqX3sba45o
Urig/GZqviBV0zgE0qQcIoFOF+PA68Wq32D8j+/EayAWb1Dlcu7Pk6djz6UwjL4P1hF7vnsfpwtV
k+qBAMjTIBl8aOy8u2s5lcOi7rFFuy2dXS1d1yUM6r8ZXz0SJz+65Pt5smbytyy3Y9jGQ6FGkJbD
dmB6c4095zY2zFyoFDlmqEwxpRZ7xESME4Ou5dfUIsbVjatHuYkD5uxh2LH/m51YizpTdtD5UUVK
SOH9LkS/P3rkB0bXuIpBLL1qTOcRzCyU+l0rK5GKQ3K6W9NsImES16o+B4LnnQUM/mWg3SLsJNCY
7Hf8I5QD/4Pph5Ru8QvhIXT0algpWZuD79vzVo8XmbIQpp/yT0gYmlYbO7p7ecRJap/WWzVyw2xG
wpCWQc9vlNz9SP0hNpVN5izm0degSlpiLTG+sNOViswMH3JyXDkhumKfgyEEv6hDkRaeVbmrYda7
JBJ4hF2YMHzLruOdHY7hkkw2FjpEbo9IstUh7dzkRFn1VIfM/eQpyIDgAKI52i6/V0+KVk+sLthC
8Z0OD9/Xi1JFjH+oeOY9i/g377vLkY5QiQqPrYX8Wtp5zaZwdq/3rf6EKRecMQbN1IFwNX6GacvT
0cGkonNuRoGotb+YyplKwwiWHzn4Giabv+Pfe0jSR8++DAlwMvJiyBw0f3WCbRNu1IhnL4ufJoIA
jlJoFsEYLD8ZX4ZjGTR0HLa4BMlyFj6j9OFQPwQpmaKMMAU7J7Sy4JxgfSdO4oAwIyJsrFfb1KQF
i35kEP1Kdf/v8ekM0u4uF5LDBCJLyHJycWtCnYaO7keYkQNWZrHgG55fkNch19c9oHAsJTAFaYvI
JYWe3BMDvt+H/DOHlor76JHLN5IKAW+5xtpvOiNH1C+oi8LY9WLBc+uVHNfExVn1qjeYxLdEv57K
opafyEELtn3t5jVbY4pWpksapxuTbOXrC+PaWX5spnye3VFhKl8XWe4jyRXJ1AO9veA8pbNjyOQB
c/rXsp6CiwVQ9Sc8stddpE/CMIpUQb5co/quBpuW+BlzsZzGBPYQRxI5WX1T1OikglQazAcUxPiJ
tfkepoaMw3SO4WgxZ+UWVMqx/zJ9qwt2fvZmybKZTfY2eB/tkwQ1JdnVFe8/PmjvQzP2oGaVb2v5
BmDYEYpYhUJPi+5PJ21gA9whnyYZFGen4yfkTE+2Xu4RKpxvRA+Cp34qv7P/n4GTTJXeWbv0QSJR
/1/8JA314IdtwadYj6ibRWrU0rbyzlQln1aFpMvUeZU0L1YvOwh7DtPJp6ZPWjg+o8Mdu/6cZKge
LX7HpBOpuWyelmynAZwLDglXI3OWTCb4qCt/76CRp9AMHLWgvg5k1K5uGOvqxi6hQYPVXhjDlW5n
YlNpo0z31T4L71mvkg8tPNvlOsXq+TmHd2D4+c77Sh1IzwnLFKVQrTQ5AQhhJU6hTZn/xHcRUEfu
jKLf3O4+n6XAACMf2m4Oh2L4NEBFyrR4f9DfSV+hCP4Nsj69xRtZylb/Umx5CGVGLNuUC5nx7glL
ldiTlc28HW/SSZA4ZxR5axY5SIZT9C5OeOLvec3uoeECMc6lZ/VQiduuv07RUXwvhlr1BIZBWxf/
XBqwY5ITMUFe8ggiDfT53hs9or+AfI68jORlCIgYSYiyZri9XHi6oDqdOtvraVbgmGonV/bB/D/w
72+5LG8rc6bMpCxyDyN6pnyxP3HKtGi4W0eK0zXWmMcmApLufmUh5T9KhXnU+BBUOq8h4bTNXKw0
SzKBtB9WH9L5h3vQZ40/Sgz0MtSDWdWK9pAmiz8jvucNxULA58SoCVsNcy8Gkxi+WkjsivCT50GP
qLuJaLWVHKj3pz0UPDG0KrrlOi52QM/vf4Aa2P+5VPKdZhQ2Se+EDCnIkONbCVSFj9/hu7pX/397
1vrjdTXY8a4lKn2tFxXmssqnQTyOFs9zFD//2yUtlX+5lrUJI10x/kUwikN9erQnaYAhrz4SU8QV
rG49YFhSKQuvM2mQGTu2E2uj2VNT75nlcoaBteO9ADdY/r/s7I9jxuh7EWpSzSH4SGX9vNvbQyuh
/rrCo8SFMfFYfjo49oCw0LakLS8bn8VcfGCn2gz1qh27LeK/9gOtmVYC7Kpys2C0Dw2/1DU4HxVQ
zKVwwhPGtrcAd5861VP8CEE9JkWBH23LchTKg87M0nfvX4MW4H3ux+mltQFxAWmYcW28r2pADBeG
HP5Ej4P3Vt6DiwIOBcw407FfA79txPxr3Bsbs76BRiApT0e6hAOYcW2krsojMgiFKemUlb+iEbdS
i4+41nwtm7k1+PhdWM0nVrz/39TP6dllkIuN8DT8DGCtpv3iPDU2neRGUThS6zfhvFkt3vu9Wk+z
XJo76yUzDik2+reOuZlchBnYo26V7+630QvX/eGSCqVR9+zrhwZuqqPQo911EjgjlZRI+xM/P94Z
tJxio0iflodcEcvnYmCvNA0lmxl+vAEpTfJaqI+9IYg+/o+2TWdIws1xtBksBnbAs3M3Ut77KKiM
l5Crulffr0KKrVN3VfarGR3ggFoRQohY/L8XIsD2xoPETSGhjE4UP9Co63G9wZVFG5jD1SEWmzjH
k80HrV5ovlmLCJxzQtEhJHCIgDJtuPBZidpfmOIc6BtHDLAVK4Btmw+oJoSfZXRQGLogbl2tQUt6
sEmHrAYYWLSvdoMvba0GLhnc637V0TqRdKsO+9KR/Fcj/w2sbDdhyZNZKFfxTid6oKHJEuMOckCG
GwNvfvZ9fsRAlNT+O3LdF0CYOk3+31rUHZUxjXeJ7Rh5Url+QoV/AAlBiGPHL8G7YUkIb81rvnUm
iafi9LneueiPnOVb7wYuQ93Oz1ABIFlv9SaAGfWEAtBYoTn4gBLb6gpZdi6PiumAiSZZZm++e0me
3k9b99puOx1mR4UcpXRwJ1fkocSk/VLlVQoCXup06/GPsA2rJsT45/DBdx0raWRwA93nnXJ8DEZT
6ZXhTK4fO6wkQjiEySEjI7T4xRhGsEqK+X64FPRoN9Oa4YCZ/rD1zpquRf8j8ucTJDrLs8MQ08Nf
dVszanX/fkcD0Iyuqo7QGDJW9tbRoGrSI272JcslO0uPw/ipfVmqTOleMNV7ltmcDHamGQ+D7iF1
jvd0ah94AzDMTEyPodojJyt17vWdIsWypNsRdGypIEXXQx9DlCwUX/AbQzfhAyM5kgZXGWqswN6p
zRtbkQU84BF1YWlhAHkEtqPWU9L6QdbzBSpsxfomB3l639xfivCmXAmCGIpSAwVt6NJ1k/1u4JIB
7CcSRk7d7sBbZ+aFSOtoX8F2KZ2mrehqyLKVo0Yqbscn+69qoHPe8NySp5W0qOsqExEjzyWwU+5X
94mhIsa3kVIuDuS/cZPffmG6+8IbqEH8IHJxY8R3euXnVbHnjiOe/si8XJFJPL7Ar08iR+STtqgb
sTVobZ/fGnEnCbpcIIeE8DG70e/RJGPhJh/1ZNdKcVb7DvitejaIqRiu4qYVabI1wkQU4PrPoh2g
LfW7RIGgvBk67bIMs4pi9fj82Jp8cRJ7FgWQCpD7zlId/iHwmGlKiVtlnz4WP8kmSulv9uGqTEpa
aD44VITfNBmFHPfx90nDhBvDo0ll4KfE/D4h+I6tJhzaJsoziO+bYGJCCretdupn4gAchqq8S1bg
bbXHLjDLgn9NcBLdnLh33TZsQHEbR+JiYRB+uWJHXdwyzLBfkIMO0yTIdYU/4muQSAq4jXi0Q3by
Lw1/EPudc0/ai8WWPuEcIHZrp2uEPJaWF9TojpW1TNsu6V1aoX5wdFUcHOhU5k8TqtbjI1/Wr9DZ
2ia+YsA+zyhNBwfn/Tr9xVdPB9e0j/bdIUXeWg4UeLKJ2me3SAKJ1Lpal/WQ43zvX0fVneTi4ut1
LbOpAZ1LoaUUSXZtgId9PZ/zylWc3jBBnQ7F4l0GGJSwtaTRVN+e62/KEimWt8EKZchf2thanFfV
PWhKKW5nKIJ0nk+JrWZkfe1qbuVN7Dds4jai39gzRoXHkLEf7DL0eWxaJgFvhbxOuoqpwB72dOZu
Wvbuq73eGDkAz4hnRKB/rutUdWh5gQzIdssyhDrvMx5jFsbexezAeP8F/xDWCxkOWCHUqjeVFsjv
ig9oisqiqBo3ESrU6XyW8NbUU6jfyP6EqMcjfVNaatq3EgT1MEdPCUPVxM7YQbgzVdpG4mdT2gtJ
7r8ZoKzFWXkSjlcPamwRAO4E8SW7aqXKUzegs7Mftin5vkXFn3IGw5pPieLyUBFcSW1YX7FLPw5s
cqXLxVb2RgQ9eSuh0Nh7iEJnqDn9DqEhytbVDDBhq1ZKRBwwtJNQ1R+KbYzST/i0hofFgAZVr9pg
/Ae6myh++n8falLV+2CCOujGnz5Kyxfml7dog0o0ogo7cQeBBAqu7v9w2tyZ5X/X6rhRpg5A1olh
PEBL6ErkhFdgaoz4jgKObJSFZuOG14qpzWjNpaT2k2z5C8wSdqvuMM0L4MOv/JPcXjvVYh6YwPUj
M8CaYmqLClr+abgaYaUKhVeLvSFb72k5X7vvo0pLKf1rFmK9MmBRcxmUQECogOMI/Dx4l+NDayrE
wboSB19JevxhszZS+zuAOCj7jAbjTMP8oJX6uQeJNfypDp/RJWlkrGlubF802KESJwOMXJUaFelt
9lu7NaYlBCsA2DPiOeA0yHivLo2Gvd6INsARO1eu0N8/GGtBDqzL/bOV1yaCAtfBnkA6ONqJvVHb
NUp2FfwPe1E8LY1QoMCe3/9pQROGgEbF1sgE+bWHmfNeaqFI9j6QfkLWepgPFxtoEIefl+YQWamQ
S/VFq08XoVkd36yCfb5ZBuJ3rwnZN5Kv7KfEAeeLLBgQvv4tG1RB9AicE72nkvvSPWlz+DkpPy63
CFQOFR47gCEJB1ddWHyqY4sjyJ/IR/fPDtH3oBpJfgc/11ka/GXepkQnIHXQlK6BeUBBpSqHYeCB
pn+RoKw/1UdBSWBRbj91cQ1dh2HryeJvp3dLeXP4iMwd6cu3wSavelugU0PDWFcRLDfMUXJWCz50
gNQVAGvVy7UJqCYMQLRCSgxg4UmlDpy9hJiqwKIQv/Nj1GP4vBzEmKA/XFZcmmsqs4ukufy3Q/6N
MYlGSqlnR6WglDr0izyMx++jfh2TxtWOykA02abfCOxjZSjXLMy7q4H4IFHoDkHzhE+DPlYmJjW9
s1B2XyLr+NQR7UDskSES6tF0IiRhIi8VQYwguL1VG6/JEyIHokbDQAvjDAo/LZfKA5QLiMgYi7eg
ccIxL+9tKnQTPG2VUdjNN5Ma4CYQgwVaP2zIq/TrbbzUeaO9DiwWXKPlNPZsapQW2kr2Llb2WL9u
pZeYd+/VbcMkN202rVwUtIVHsdUeUEoURbmA39Nd3Nx2Ubg6AVDbvY8MXjY2Lh+lppL2eqKWPlQT
mYWT8OHqypysJ8Cb9DC+RYv6OWLB2cM8Oe9RIMwBJOJpb/UfEPrnPDp9UXn+olKFsyCZf55D9Hey
0cccFVzbUv+NcCyg9TiZZrZ4clR1uQJPKXNZA0GMywy0VtOkI0NT++5TyNAxtx6KhgudAGe2lPMm
0pycoXiMyD1AVsQF6Km1pp4krNF4hk3EJu35h1M/OXsij/87t55x+Civdmg5mczSbitFa07evIHG
e8YFXCd0MiSmBJEP4pHFnzjUqv0DnK3MLwm0bUQSdO5IJLTMCtfP9dBjhm7McsA03epfhY41Ousp
DB3cV4FHhZPVXgnMENGJNYB0oMqLjtgiMq6pEYQIwKd0NEBwMMgEPB7HkWRJv/kJzfpoNpOHHK88
UfJ7+hIwp6ySpDv4jZ9tScErYeq8wgqDsYy848Xr4cAhDB2og2JjZx2e5zrpZohoaBDSuoyhl1n4
2JR50VZXo7UI9asKAw2i5jL+LHThC0/NddD/EHbopm1Km2bIfJQjgBg44KBO0WaxgWq0P4llov3y
i3zasRpV7xXUQZQQcTVZMBjXt8nPkcT8MqgkqvgftE3S3eueOMrP3JxeIJV0INE56POSGil8+E8W
yBVzMihlnngViBoZ7arDXKpE7cSAw2MplTHYVBP+LZY/DtjoiMzSDeR6EjQlprZxgzQsyoodNKuD
43C+d00h93fUSMJQcnvTACKijUXbOdajWCeenpSn0WG5XFMwOu6OebeCCFsZZcgznw2Zpmb0zEJn
om/LbVNA4y+c6Oh/JhgKMtRMLPHyCgD2M3EmbhCTMDqirxA2VlBQk388/vDRpZZWE48v95xPQE0+
128Dirm+1AZ5tG1f0NvlUq1y42f4+jBlqlDQlbntwgFSCrHrO+fBnCU9Q98Sx/dm76JUuMuoN8dF
FKhSOfeGTKaMOwNcLcvJhS7bghlB7V49FsBbBWbF9VlhJbezLecdDABoXJUwKcS/yBnanprOjzZo
2WcAQEmyp+lB2aBkKggG+D03Qiy7PSJAqxPkpBScshJYzCtE8S3IRBSHmEqdn09evWRbZIvZmIru
ORkQAFF6sTkWYLnpkdH9E/jwSTte8M2aamjiUMVN6FZN3JC1jndmJNhQ+7Pk9Q00lZzaUsunpag7
3qwRr+7lTMWqrUhahwK9sTBPQpKfwtW+ojSfCp6j+UC5Zb6oXVxzzoqNr/xrbC/MhT7G5o0pLdtz
FwGcvDaaynvkXezvGY1FXhrCLGVcOK3r5+WMPn/ml781aVIZtXNGjVqu9PFGS6OKkocxVLiLT27r
eXoa+MZzpFJa6D/m1cyBsJaQw+69nAiEp07/y+MXynQi/GXudW2AlzeVeobAI5ghyftrEJSWg6eY
e6L2GzFzlebqSs+qszSv86kYnEA623EMxkQdydnD0ha9yHTSxBLJlsyGLLHUeR6SE2bjjPlsJL8S
mfNLac2LAQYg+GtxTU+OU9jpi5MV+KddhaV4BlsuD/1joossbBBggC6u6k5NtBiK7YQh2QKIGG+2
I0PaEE4UK+LOip8m/WvE+N/NSZ3hpdiYPUyKkwkW1lXhRGmRcNfchDuQlT2hRGk4ZwaGklAPxgS+
u9aD9OEp3UFHW/zszU6FHRkhGfvPVLIfv7Ewd97IHBrWAOVkWEendkti1BY6GrTHRHLvmPcr2Arh
aun7S181FPxkG5Qh/IQBTW3S2s8oVk/vLbzguMZJLO0+bDkzLo2xH4IakPs3WQeQiKYmGe1sF/bO
T1g3kSOXsej6gtarhT52QhR9GsxQ2/yXLR/9J1e4mDHdMffnotBnkBavRjJj0goWDm5uEW5ShIOL
ZHjM99NE2vTHmKthv7N014ska4OnJvclcwZ5YIjtLNGNl+ow1OlaYpnR/+AHeK3nJV3Gc+LoMuBS
9FDyxqvrjQ3yVDBMN400Ae9IplHSgmG6qdFVLGvyD4+Twq0J6MEj7zx/IBMytn0CVkzZe8IgozGg
9QVBK/ymX/BY1XL8708jI0vMtiY3tD9mhX6/Voc2Fhb/zEiEAlhV4FlubsPTFyHOrx1avoI2ydg/
UtOzj7OSEWMW46Yai4X3bilu+/rqATv33oK8qf7coqibOpJzMcSNCr/dnHHD9bszuuDOjevfU8te
xuM1ZeLqFutaS9GTlgdDLg8zRFK9q6wHLw5M1+bPW+sVM31VEn5cZ7WbaCDZLJCya9EES9uqisen
a6tPaCgziI8IU58u1a1C81wbqbeR3OHR1UzoGmStZMakF2j6GRMhg6Diex9ghOTITNAPItBjZqgY
2ygkFZc8DurvHlncw2VIemN8o/DBLn4UQ3xTnW499N6xxX2nAz59sWnNxqqxkx9vuCwhdWDTvhpY
8iqhqMI2ZGKELHFH9bvEf6+PjcegOtmo10OR67E3q0LJUCHdNU+ro1ziO13DaO5ctQeTIwBVHFES
FOM5AP2XDq6xhzo0ipLYFGMfmAQ9gR9gQ+FuqGnv2hIH7jaDeiN56xNwB5BI1GskfLis7EBDict5
wTDY4pb8X3B5v8mbk6wNqZTtYz2btOn1VH76Vqkx7k+jSa8MzE5s2Q/XIvYa/yqO6RaJlay7YqlS
rLD+cpb0bw8d1/dCk1vCV2QDM7WT6tiRsE/4LFXK4T7pWjLbrpS0foFxMkrevSTFc/bYtc9yDuT+
Hp9naVFRboRuK3r0iDjVoefjawWtCsiSDk5HT3LTp5IluPWERdao2rBOHbjEw949MlAueij7x699
BNVPNT8zhrbs/6rtuZU5MhXUghKR4NDkTf0HHhel0MATKv8QVuF5OVqYMwYE52Wy1WAEGzchS565
345tLaG3IWmBwIRhMwGl8f2n5LCAdo7fYhYkg2wzlfELuHxzeXafKb7WWyO0qvaYBF+qYt4gIkdD
UV95dzVKmJYtBDk3ucpsjYUclrTAA7ot7AzHnwmFwyznCwkg14926cUvZuDzJYBanyh/AjcLxfRz
4YcayYWQif5pJnYUnQw+UtjWHI8pm7YKiBe9GgJIaXequrGEg21o4VXo0iA/xA76/eZMdUk6P7Ox
ED144sIXy6Uv6eoqwGT3VTIcMsWjUO7pGFxuMgB1EQN2K7f2Z3Pmwcda1e9jktA7ziE9yd6o1N+t
yUTtfnpghq9yFb+l+2AYADtruAF/pDurS+EdlX8PPdNQcbDyful+8Zq+KhF8mKA0MywBP/e0K5yD
Fqr3vaVG0bp5pdTKOfBBi6VJV2KUHhoeBjlNyecz/1LPbYh0O9J/PKebRMeaqMQYcX62TMCHD//h
XLzGEkPVec69P+eay4jWmHIK1NL1ZXB4kkLjrOZ78+SFx3Z9rB49R8EgFJ7faDqqFfG2V0om03rH
ab/3YqK7vsKZlTxVp0Z28Qu2An0E96cdoa9nE36hWLmF1ph3Aods1l4ZNqwHiGQzqtr9NgosQMrh
6CMpdQpmZMEVziJmN+Ax8rnqAnHZLGHpkkhO329thODGuFwRzQ9QbKdNgjaAbZLV6eStTgU6v17T
22+N4qmAPhgd6Wet7mWNj6TJ3uibR3fHjOUXG+pWvxYNH2xfLuScPG1seMBV8qTAS3/uUqZNzIUv
8qlTH4hJWKAKWtIANfWIwFK5h+uxR40oXoEv/5h7RbcSRsh7yJZ1+7THwl0eX6Sgkef1ytJoeuQW
w5AAeBd2SIU7GXCDAUVkn+kq7cJwV8jowfNcem/z5YVn18FyaeaUJJJvx1Ge/C3ZGF51U2/Ra1ml
ToFVANv42ZQ0Wz1F8fh0VNwsi9ySUajC0S7NsfNVMoKfkehpXx8O7SqN1Z4SyORaWdwb8bU4lQOy
IzBpNLmZLEs9eMAMv6wQVrrw0CnFaNPhwMRBjyACz3gckyFTQfLFgJuiPkJ6WFbEViWhvnmk1VbP
4qbWg0YAplAFHArctT+apSZNH7jOSt3TkakEgF5+uf8Fmf6A1xlNwG68FCTrtRRy176DcEzvn7lr
EOhPkoxPzKiYqFi21QvNoD2XWiAxM6s4nJ1E0RKo+mfhLHTK0I4LedVPzs6AV0s+HPep4UWKjeHB
wBTTLyBYqY1dzeihfET40UEtkcP6ojGPU2P1J7zxbKZlZm4czIw8tZz6FI9vBf3oAMXKyX8bHlI+
UBsqqs3D3QjZuZLcEXKSiWRJAW24I8SOxLj2d5DPSugiwfhMcpneBRONiIVKHvA2gJTAW2SxdPrm
SC8O6Vp0WRsEL/Mq5GD58LgOYoeR3S2kMRo2DOgz7L7iWrNhU9gzexA8DGAkYyhXhRrevk++4Bxg
LT3Npxq81Qn1EAcdXOARC26z4ryqCUZLX77qhys9fO5MrlpKr4AegpBCJ6/oT7oZKgJewk1JGb+D
eDIvWy6xU9qHQ+vaEQ0k+zBKIfg/3Hdi+OY9ONJXhAENqCY+i1Dtu6QzGrai93K5UM6NVMXF13Yr
+FYnvLYxOGNLVVaHOGhzNLXojKs5M91e4hjUNATnpQMQL+Sdfd2nrn//eu/dXknNACUzwJKlHNg/
eKr+xM7KthvitQ8CyWZJzhszJ2kAgn2xwyDkwjHWBhYJznHYGn6hN0znHifyTRCMj54Hr34sG3u9
nV5t1KSVAFFw7RT0HY3B3PyGielfKv1XWTCN4meZs8Gn10xBZe1hoDJFlAwFMkoM1VVIIkmze3ms
Ne2jaMlQsGBm4mdXYVbFQqQjZfSeZbgnG+/gYpz8x7CporU2Tmz5G2QrI/YvUMx9k7DIiyAoPo8I
dhEx7GaYs+M3YbJgu7WKKFwg5+lRsoIN905kRoqkAG4Q4uyxr6lW5Uky9eqBjtVfZZ55kC1ck+8+
iOve6q7iB+PxltKT9mEohoEkUh8RZsAxXk4J6lswunwDTibgl/GDbft5sZNjY2NxYddcBP2GIyQT
Vh+tAq+DYnCvRborW7aWS6FHl+29GKxLF4aeud8/hLbluJygFTY+M2RpsQ2Tlu/Umj2fqsF/HM9H
Y/PwGax0rAtydl8xADGK46FOuOEETJuzCTQ1tH8Dm66s0Q92s+rsE9WUdV/MjblF9j21tuFLmgH8
Q/HQOLoQSo1eZNWqdvhoMKUHpG7oO0/5N3Ei6TB8aQVc52kr5MUDWvCv/RtSwGjyZwtqxHP1G07h
0MIQ/DTlwkbwgfHIXeGT2apIBx7Qpfgv7q4PHQTQto0UJsDb6/+VphtsRzAcKWrMz0ztMPcpheMm
BJzUHeI3u5m1h3Yf4MpU92OSAseGlSC8XWqwyR57fQBMBheNG3oWZfYHfNYSFCVVy7mrysi7dSve
4Yw8hhpmfCFnGbHnsMowqdWx5QiLsDRMskjqAayGojW/67gOzc9/gOw6efc2f9OZSHc9Qd0qsaAC
S1cgppFNosfgA6KIfH5YBiGBazXg4Bi6tNb0Jt8KTeluhazYg23aZLejZdawMxGhSU/XanKlyVkn
bVKBv2y/c3howwgvJYOyFghP6eU6pUamkV2KTGe6EDLeAVt9PH61dEk1jYqfz8/aITY+bkqKDyZz
TN5ZWN0lVCMHDJLQulNNXPBPtgQF3e1lFJm4my8mPsb7izWlaDsP8PuXCjZn/PobjdeaVLzTtWtp
sp16aIdpY32/t81XIY3EQTbpdVp3miBi9VwYkZq6/5E42h3nZN1J3MyPnnlcNBpNs4c7z6V/XiX6
b2jRg3DiQZqVWSe5b7ft7YeMNBir5vD72O+jhh7llUQmDdEsNJbKEh6yeTftfnw/ovXDlK5yQQ+V
tAtJYYdcWNHsiPhAiebQEGdrD7umn4tlZY3QiS8XSyZ6RJDiXo9jGvTulalt4+zGchUEwzNFLVMv
ZelYYbturRlHJCFOSam35PK6nT4Mc/IWQtqWgo/R+gWa6V6p6Iy9vh8ORvgOoibCvoT+HFDbobKs
f4+SzYvIScWB/h8bWhiwao76yV9U7/LUkQTmF2ds0WV8I8+V5MsyRwRs8TrC4n583heJvHiE4/E8
u0WnMf5dU0/Zz4JEHpc7rUA1QYahlE2PvLP1lBLiSJjH5/6g2uTS9h8KMSk+LyB1Z/gKCbHntE0k
+VRev7Y6zF5afXBMGr8RdfnN4XwUMbkLgXVKCo1X9bPp+hCpe6SaFo4iAnzhkSv4vJhMe4HAAToC
pxNl3RUO/rauEBfa44chNKsoyDH8HvbTGk7gWQVKTDFH2/g6AgCYs2PFedxCk1JJDMAjJk8TYQzi
TylMJusA1TDwzUWrKTUmlAPLgGJgJ2995Vhyjt4eRSIgGLNW6P2YtGCPPsdMxM/rbiH6XOAVvW0X
N4DYE3qaMtOOABVMHzp90krm1J43tPRaeWOXaWV3XfoGmeKLNGJg3wypxUOxCwsVSuCWFs1pvi9J
+NS6qeli53rlGv2tdVVQBz+XO8xByV2v0O7sbHl7VjKq9mPdZRYeIo+8yoxPbFLiHTWqcUvzo7AY
355OqCHMrjw4avdQNY5umHpJhGGr+BYULL9awBlN3yUD2djoxkQ+3tMoShaQ4FcbpgEUGehA5RKB
G8ItLHbH0rFed5RrwiCX8MSLmAIIlfXfwE4qG0TsjWNl2/XlmTdsJms5NOcJUP8M762cIpl9QLDd
8+OsOPJwl0SQNfDX10gHAVkr6oOA0WfuHKnC0tTXdMw8GZJ6vbUiSfotKZ+GnjIsHFthbiw06LBO
HE396TPPdctRnmpMATjmxQ/KtLfVJ+j/q5L076omL1E9VOpU8arjZhlGhm/d7Wwh4Gx7FGCwfkR0
6IC8RAr5KWT58ZKVqNzbcofXsACXrxiXD/eVjzWx4j8yuO4e+MhT01ZIh98Q87JQtIrUad9V9Z8f
8tkNWS1Kxe/4Q/pslXbnWoDPwf4wqgKUWGrF4y9x9ddJNcM60cYC7Sy9092bdos0xeWr5LP+4Dfg
qFI/m+EBMVFhmlljcFOo7DlFxtZBmbii2N/6bTogY+sfDPaNcAZ9jWKuyJrjulivRMmEc6lHXnhP
7xD/GAp1BfOfLGue9AQdHfpAMMFigK+MQtR1a97gKqxqEaQd054NRlpGLSz/H5YFWgJL5+DLWSs5
h2tM+NSJ66/bC/dr9YfKvsH/lNEruMn5mfHwShIkr17kiT5Q2ujI3DsVsuEhxD7hgJ5wIm8Fpz7j
Sq9sAaQlSTFShY1Bat9+MdYDQUhv6jpjkqRX5YGszSU2LxJNe8/tdkcLvSADHt8D3D+17CGwdlWJ
Lkc/G9EIrH/oT/XXMVfVK83N4RCGwedbfRzo2e0CF5sQ6wdn5b1p7FNGrUzbMwstnR7MUDqfszOb
b+XCaPG2td7WhPTPhd3sBn5Nu2Vk4wA0QUWxZQfiamNiD928pi72qFc5RdwmFc7eqQO3D+3T61At
OxzhmuRg/gInOdMyAl1amGAdKeObSZtqhGDjs6soT82czlrceDarVpPzvN1smPDZgMlIllIu0t6j
7OatuPU7ofk241+j6PoJAX7MdtHIOS8NWAtqMlMeciWeHCH/qGaMuMZ2Ne623udehoBWanURPV2g
GVZI9zuWY+0GHV1f4f/dltz39yGUTMnLZFbJp8WFCakMVvxTnSX4PaB3RiBGyY9ze7spUonYOtBC
yUa19xACx6FocbP9Qa5Iu36foT4lYS+qvHTIglvO0EdJsQdt2k+hSyGxcumHTqD7Y2DHDhton7Bn
KXyYMSPxXI3TPM1vvzCSgPmSRnTioUndtZgu2gGRwCFnQh0XeD0vuYS2As+dG5vyfcylJHNfKsBq
or1yOwb8zK2ytDb6L8M2a/d9+HRSNmIXPuWnGHoG0dRQQobYqXm1L3vvxFptAJyiUegH4fyRY/br
w5zsebQAMPJlc0V+awyztOeEitDmIQyep4otLCTQr2Txl1SCpXBbTe6ms89zvjJTYQGoUOVLYSoi
8B1hQtWrGPwMchj3ndaMlYA+9hUy9q6r0U8zTXGMgC7WS6NCWzQ1CAkvP24P6vHMzOUuJXyWO78M
pMeILB+fcU2pE5xQVccq3muztWjyJLAG1W/YD9dQh8go1sBWTzYzM/Myh/kOP0D2WP6m0UJk3HSm
fUrr6NetOKJP6kn8RZJ/9ELuHbr85OE2axfZ6fGPJVU43qRoV71fZMGcGGc2ZfYysltmoID5ugbF
JhTdm+z4Cy/hZersgW+CLL6ADzFTXGN+CAYU6BRl3/GP0wwXnjSwO9TFConWSsdTRjbkST4CE23i
mtH27DN/L9KuAOhJpe4Gecsnlb6GnY3qZp0WE9M6f7GRr/CvIrgUCt/x0Hz8R0PwPOrxwLwrLbUo
QCl7wiwaTD4ooZHYp/XoJhJHTRBe8XcIcA5qM0EbXceTY/6CnpLUhNGFs+sGzkUIiafYjvhISE7H
6rpB5iXJa/e0lyv8dze2Vfs/uw/DBgimVVvAJn2LPY3o6nhRAdATQ43KaOqS5kKRqE1DSnQF2Xe/
RDLnU/PP/4jAJ2Db0rLsJS9Vrd5YlkuBiRrQ9xqdCFkP5uv4lQ49No+38BuRPDcL3wgYIlIOorpY
N4e8O0YcnxkKwzMPkdZcf7LY6FHAvzKBxF11LAMsQh9F8JgLMrvW8ws4aMs4OrSswl1/NBm0DPzY
eYIOgqArllDEfvj75zNWf2gSQtVYEFo01Dpa7zNXfzFdywlw49YpDGtH3v73w06z3VCTXk9lYzF2
6U/xQdFn4u+rWnW5ClxNK5ir/AfHo5FH+edV017avsXe70KgECboUTtVSLTTYFuNPMtmdfN4E8Aw
3Uu2ELys5BOrik5EcKs6PQ+w1eTuhnOeEwaPaHitEEJOLyVeT64ir6hJPT2ZwAgPukcb9ZNSjxpJ
ilpYc+aiuxjtNHBK/dOrU3s9BdbUsUl24C58wptZPi+owIqtXcW8HWTO/8mbxtaZMzIupVUFTrDA
G1nABQqy3Je7zo4rNHAgS1779Ddq2WNik/2uZ4ghlMrKhnLhPdXoQN8TrebPJDQRgq9cPEvH4h7q
7cY+1S3U2MCF0q7qirrdOwqwyUD62f0BvL930eQPm4pY6/5VP6vThIViVnqHu2pOX7h5fbO0xkXE
K49+Y9g0koySLfVHY/MU4CSEI6gBEYqBfjvGHO83kg/5KfQihANSGjtFgRZh/fUUuTIIJs17ym3u
l5cyFelCEn/ud1RfGpH8+Yalz+4l9yE6afFnQK3hzDkWYco/5bTWNOYKAUJBdMkEJ0jD8fFtoE4r
WUU9QBy30eysP5/IozicR+WkDYzTyo6tiHZ/C1Nh7MgMj4Ix6w+Yk7X9cnZ4sIiAf2PPcifx0f6S
GoyJD1jXFYKe12stMv1leARXnjgbirQaTCOj9c85IFwg8Ajaz4qNavGXsjpE7OlvFkoTpKq8QbQq
a6XglkayohkboYlYBRWrNLL6lafRSR9d81ozAkEYrWTFBpzFNZ1lIqEzrEYtNM7H8XOkhgHoYuBq
g+pxvfTV9mvgYM4OQ2snPyWZZ8bfnVm2mn06bz8BsatlB3OoG4LDO+yVR+gZvxSlWmQVNVflmALD
DHUzb4lCett0+RCHjGZ7F8LNpYsEoS99DQSfNkQxOrc4yRdqTZiqORRTQG/md1hFYD4UTc/cGLgE
L+ZNZ/PSAW0IL/xW5sDVzhmwVrl1LgcIo2Oj1F+I25yG3fuUqVE3mOUMA1c6Jn5GeoLMsoIkkYn/
l4l/AthyR7vPw74hjgSowpBjw2Qfufr/SL5M2z2NiVAQlc3+Fg6Nvzvhu9v+YG8L00DwwIxuAgHQ
hFYCa9ivBpKyl3G9KEbkyIcX+CzUi/vYr7+guZbqtO2jFiEi6t8GbTU5TZ4w4kYUXfFMnNsEo9cF
WxJVIouyltjdGpFYMByWjqVEDgVdUGTss75bzby/bP6KqF9igKi4G8qC8t5pXtcLqDhjOsvkaGag
lZxPnvkj0D2cC6g7VKTn1VfV2kCjydrzXgQcBz5/WuEV2vnY7ikdh+ctF2tbrTWLITlGJjmVGthS
mJIZKwLFVGTN1WMq4HatNjuwlrMErKa9UxQ12NjjMCog5YQ5qWCn4Emkh3iHm7piSwZlE8KiAi1q
aquklA/PIUcyhPfZDAbIwVTW2wTb2ezyLFhAIeOJKTP1esss+eTVAJzssnkz9BJFsFrPq0g1nknY
k8TY8KlITdPF0a8ZsE2OZUzp/zmfQjFip9OV0vwv/5cVp2qUsik4LzuYjTGa7gvNA3TdMQ/8nAyH
CMdRGP0wW5hugDHh6uPdC7h7TK67UGENSfm0dSRC4cNfa4ZCDCamRzqwsE8WB2f+2FZiTqncqmwO
KHyADDZp7jEDM1sgcT+tP+5pMK+n9mirYyo6KeAtrqjZEXG6j/5rGxOj2ac9+D1iWzyGOLS/Kpp+
BR8a525hqXmyI6ozkWOF0yTLw2ZxMyF35HXFGziygI0O2LNxJncVHCSQGn2iSuAidBEJ9yUL+amW
vxe3WZCf7FCTfuXB+Gd7UL+LfsbtXv2n08f3PA+RwrVxWZ4R1ACdUHYWdQzEsj2YngyaaLv/nCu8
m7uBtT+LidN0nMcM+ool7e3r0AngbLEHQP/Z2LGZDy62TkK70t2CzevBNHnkI8ZS+pTXHCdv95JP
F6VbS1AIkl1vhhpnbXT22kT7MKwDeprDSjiAC8ud9GuhtnPekpbjYO1BROAxf99J98XJB4JcdFSx
HX0u2eGuNtxPu596Jeu6ScwHzlyY78KwUL2cZ9QQEpvO4D1ug+zgVq+wMu/7QTC+c43u2kbzSUrI
mlbuvjub8ub/nQvGBmpKp5hDDqTQxUOl6Cg6u8PQ1mNNFh9/5QqsQBIHoaHD+jAkQjNvoH07Gs+y
PnlVKk/WQ6tcVSV4ubYfcA6dd81O7C8MlQaIdF8Ed7mi/BrRhaDLPCLNgvAL/5y+cjCIQbq8SXjn
qDSqsP2Dorl8Q9SzHcfJyGMezUnwU28xt6jNJL+EC5Rxh6KjZnISwUBbVLZO2EA0v1d/MA2qW4N7
7vd3Ui+yexiB/Jd3HVO82unj1iaWqzATxFn12yDjOnhRhwhWVK/34tefT0m1qsGUWqUqhqsUK7aB
rUgnVPx6LYg5vaRgeqhNy03nZ9WPO9fsIc83EusSJnBef2Mi/oqGONDjfGi6S56xBfNRlU5L7gAf
JuYd/SJ6oXFUYBUb0PiMhzvvRDZVPh2AbWB804N9dnSV2uYbGwj5zBqsvudMaXTcZUr4FhtGT33G
PY+HgU88KrYNP6IzJJuC7G7UV/QvjykknaqxaDkNl3QKv0x4P63IFLsco6+ROUmq8+qIePwd4NCX
EjU24+9HFApVpzfpXRHbf1KxXn4wH31M4iH0ADB/uLRfoMj5fF97GaltGrpSih9v+ELylLv7Ug/G
KNL6wb8wbOmpHdgspzz4c2BKcO5qLuE+4gDUtoq7yjVU4+JqHLGyVf4JhhbSs4EoXBbuWBSWD3bu
25xKqDfGAGWJeD6tOPdcGcBMETZi88oPUpwsNtozsDF5x2TjuNthNIwzMNTkRQhTsJfjThIwz5bE
OQVZfSIdqEqDS8g+ehwpflz7Jmn2nBjG6TOQJzopOdx34fjpWYVXtH5FZt/wNQ1PQDoxh/zUE3cl
YX5OA/YJLNMy2+AmFq/OEjw6NsthUpnvqViFNsFknL+9KYO2dhib8eH05mRDUY8WfNjVdjsOomas
5RC2c9Zz9K+t419wVg5M5DjhHDO+GWQiD8GR9hVl+QdEb3civ5EhhOJ/mFyvPvykMbTVq4vo9uPv
Y5AJLKBzrLRwtPk8ZKUkrzKfAQE0TFIujl4mlpVO9RdnGHMnAEPKD69ow4Rk1U5pgZDDaQXKAiZp
nqfgCY8/bxG9v1k53DPMnseXd2ptPRkXDaOabHOUEtN1IcrbYbNw9IgmWuWC8MQdtxITVj3h5rme
XgX2zIw9gVeoXH42McjoANQ0xVRR6RFOJ8tS29S4KP4BWXPGyICm/s+JO1zOBLIrX7TaebPJo3Ip
9gevWWqwgGg/tqtH9c5R7RZIIqyToQozmYvGpJMbC7ZTdsgDFWz6BEOSxU/SDvSpv5wgk7J6aPnC
RfTEV66Q34w3gfDSJhRiNob11c26QyGEb/igV5Q+lMLjLua5D+4D8WrkdNvEGiDMR1iAJQ1/49dB
gmHgbDhz5+37mWCovkbrl0VCq/vIgGGCxof4kToZm+2kGBcAMJSvfHmD0EOir4H7vC81NbW7Fjo/
B0z1G5gjmSgQ3xwIAVfAZkjmBGEBzdfcNM30YnUMeOtSqEkdWK9zaqfzMlkJvdoVHm/pJLhyA5sj
sbko/S4qGqmlafewHuDpmKey2mvweuKGT6qGBrdoKAzm/aFhypV5fvJfPIO44AwQPsflDNHj8S+5
A5SCAXc4XX5QUIWDY4SsSXIBlW1dDJYHWhl0WlxiD8oIdk0N3lF4IbkXzSb1VHBHokQWqk+lMtEx
hFdCki+sIVyIw6qNEmWbrkn4KBR9+KQyOJFidKS7AukC52ttXJpKR2ExgxfpqkZRr+jd+d/TSYvJ
c3P2NpWUOb/hkZg94+M+yHDTamSczV0khQRhEEYph/S2cB4cu8mCfHztZ4MiwxNPZRcqzc6JbjRi
oaLbV/3b/MbCi/vYrBLZh3ENCq/5gFCicY7BWBjHKJqgfPIa407YSNkvlYXPjQsZU0qnGo7clCK/
vlBSrflGtucRn+pVf8+3snt67FXrcGFZ2NFDKSCU+VVW8g3g2hQaZzZ1TduqocqBlm7aOufSwnV7
MBc8MJNlJEOvU5ArHTY8kL729XSc1SLkWlJE7mNMn6PuxdEkNTIzRowdu3HkBYqOB2LKFB7e53wK
GUkpintDJA2cCjfA/c2eqsHdY2bu92Dj1Rz5cuk4k1KiGy8G96Ylm9qZ5WSlHo1eog7c6A1n55zg
6inCksacCVwWBleeplgVDYozCBosmwYuryXAyrEiM6XychbgGp24GKueo/faT77lFlrrhZylZGL3
Hqs178NYWU9sGfjoptG8v7PomRQxA6NE48m+tjYJiBw29kfxoZ4dfQsNV+NqLmnAGS/g+BfnCNsO
J/la0g/3oxL2EtVvKUOBYnvsPoWUt/SUEmsRNkP5GedXSnHUvhkAUnkjY1aTaVZVi90icd7TtDFZ
k/8v0+obSXXkgw+Jpp8wlPVgWKwKW8wVIoBCeZDigkHuBdXG6TRzbJEReTZ/03Iut5qWAFJSfJWR
NGjks7IDybs9tiu0BhKnzBeNkG7xsZ8Uq3cHlfzUBUVxF2w7iVMOQPi4iYjSYMpI3u0rA41OFp+g
vjat0PiIaoH8PQMUXIlhEaDRB70RDwrCsbsVnOLGIzKYKEnfpRSSnuQBq9N4bMPbPW+UUDZ7lqXG
axf8iFHr15cLBEGwdrvm09m/V0hxKsxeudrkE7SNfeOzIvSKQ9Md4jZNNOPQdVKbASx9TCZJUz+B
MkmdtBrZWzLeayPoGmGmIn+RBF188wIjx18N/hJSYnmGal0kaleCyI6t4zuvoYI1Ptqa2UarOEPH
xYyKL9n13A+yBOTHRhTMUORiSxuQ04yPZijZMk0eVr85a6eHd0tAUopVOeuaFnDrZ4hZbkCDiA+m
NwoGUdqKYRRFBr2d998Gdmqb8EKuz2K1Xe/8eVSoDiyr3VktaekRtpGm07v/vK37uUaS5VSdApIG
E0Q+72oM9Z6BMlUY9dOhwmQGPiBNu4GXF6W5NeNnpVecQylazVcULpaGfkdG8RdGsc5oqWM8TJlW
hBEpHfhtnWGDI03pBq+B/96s4hFWKS0poYgYxnPKnrpFPwHkhyBzMJAJIcveZw1KhprOS3pdQUF0
iOQM28yuR+eQF/AkR+ohK9yLb/kQUIuD5KbZiT5R3MHpGBN/r+9qLnEn9kdurdHqTBpFfyAdzKEe
XB2SxRiSIWTPasSd6Gdoo5PDQS++M3RBPHFQ3rYDic5rpETxHhnN5Y8YeI+TNNfQgA87/E5TdiOC
//vuH0W0+MIFjvUvfn2/b5YxTHekrFgNvIQjQuSQDOvBebSy6Kd77/Hx5dhw4LMWoWGiwkptGX5X
Ch7Jjiu+Xvd5wM9uW+ehLPQsfMzK3SwdTh3jkqeQD2OgUh1kTwgCr3qD9GbzzHloc0a1kbGUnWna
Ghb1OGoocjA4jCcJytFPq8zBrTRBcVowa7dW/OaipnNjUnk3joehWuTxirfNvj01JFVfFexPJFD3
6Ou543jNHPVRmySM7oUrJoGDpuFeosiQFf3tzIxhHuyoHAACWpD7NyxfCok9FsQ+E5Lw12Kdlr8T
wLMlznV4TfmaojK4rxAdnqgWf/0bdg+JU4Sz03YstdKZkHknAd6dPtSd011R5QGyGCtggIn2qD1z
kiV+pf6w0gmTVwiOJ8Fhevtr91mJ1OpvugzDj6+KZ8ag9Ogad+6vdDCWTN/EzI3tpYlBDlFKA++S
t4Nn23dAYDzAz8FygFjehVfYoAXehD2D5nwXYl3CbsUvQteJ87YLzQoR8ckjLQEfPXyjKpmUTSmG
fWqgfB0u+DLTZuCCN0mpFzLLpTEyGlMYE7JyWXDs18bpXslisgD45zsxyCL4C0vkqx7nwJJ5Su9x
Q52v4ubbzJ9l9j+7rf7AUmCS/bDxB2F5sVaYZUJy6BjEw5XD61cd9TTl3wK6qiLO7DvHx53Dgu9V
koZBqxBwnnQ21sfJYub0oM/y0dREf7VwkqSYaVkY+BfMg7vil3+V2MfMI7Xb6mTrGEjotvfEwjcx
bNKHzE2ZboKcIunNQ05QQwqyrW49FXMplILiKQbfW7QtPsM+oLbYSPQuUaSLk+vENr6YanVaWdGY
InCuBxALT0dKOzVK8C3eFLq6BLIzdBYMntzLfExsVHeVOSOO5hY8CZKd81bbMlKt/azk7qilpjM2
stEvwnDXdRCVISOARG4//QasuyLaQUsZtyVM9rkWtL//DHgzNQUBZdB7zQ2Sq+kXYlFMrsP4cT51
6dxSFhu/or6YHOE8sJ+uzUlURCGDOo9pbH0KFugKmd7ziDEzTNTg6hRUzTZRMNgvEY8zB5Zt1qXW
mh99BCwwsUWsZ6MXIQ5espBGmxAWXKQrh26RsCeCTSjrCi7FAWxi6eMlR4TgxXMQZ9yrZk5nGRGg
ZTisa0VGdEu1559pQEao9317rqzbxc8utZH6T8FmwELfWEl1wZcQcA6WoEvul3pHnrIY4KhgNorm
CAXK1Z1fili94L1Pp1JzUEfU7T2hulO9rTFGKO02d7ESSHIcPpsrARAGffZNvZznrdKc/Ue5fTmM
s0bvehh/MrvAANshoz2tuDf5TnwkJ125mi3du6ZbKhqhXHNjwiv4R4ezqlSD5E6UC9K04J7gY4IH
+m2oMHQ8GgbiW3c8ZoVmYTaebAI4ZvYtV80BrEyf6UW0YzQA3GgaSvUj2/f7s6CJCVQyw7QD1O4v
hEUEDkl9nTCXfwWkhwj0reJXXdsxKoVo6VJc0euG4HAcatAAox8KaB3KSmRfwQ9sXVjPswYyBjx5
OcM1lmkKxO5VwfKOjP32HRtLV5YiC74jsmwYwzINtxKy4NYk8XG+6mBYoBRf1c7FKzWvV+fnL5r5
W5JJyvdDqOowzOL/jkpvA2GQts/Rxqd+SeaOa6dk0vQLL88Du/8O9Mlx5fxadIch4oMbtgyFKpVt
K8mt0nL+61xU3qwrHlGdSTuhfOVh4EO+meCn2EcV0aeX6cj8F4i3GG/yPNQoC8L4SX2lemYUzjiq
L81F8LRK5+XQmxzA+JcKRReEaWF9DHejkLUSSYveZodjWoYFZakqDMVCl/5GjgleINj/QRXqhLwi
rttVRcA2sO3D/z86XPIER+acVYzcB99oVpDA4O5FDH8LmuDNGSiZCR6UjpCZnkAOIS87dHoLd6j1
jwHprB2UJfiz/+3tx0Zi6uSOe29CuGh7+eRNbWxhIrslZzXYIb17D6xe5J+iCjMykzpyaqto4/KO
80tm1W28HXugcZ/Q5Vrx8ZZVccWPejWOiqIK350Ly26ckPOU+EbWSGkQV034NlA87hxHySITukLa
ro/hVgsyMj7wsGBx4HpBJpLZv+sbZDZWGCSL0azTbf2UlrGxlQ1LV177AOf5+k+jc/OyQ+Eb6Fay
umP7spbIHAkbzAZjXgVTp205AMMjgeVEuQ1UB5gA331UrXWipvcaKTSlW8UCG2w98Nut9eQ/SN5Y
upNwBSteO6CGM41KhMT3qIlKcth46HGcMfqikAgsI414nD2KtysTG11BvUgbIV17axmnS2IDqE1u
WpnbHmZ2nAw2cYMwA96J4cQQnpz09XTBMe1w1IDhw8368CaDW7c2xCLAB4TFlbk5dw9QQtjVeCLb
mwn+CmPnFOMk+KKQdlE9HiRRR5ikLYiNs9oJZ+iI8z3UAo6oENvz+oqf95jBYbui63hZdvtgtLVZ
l1m/MU+VDnLvQys6Aav4gE5kPeT0jI9VS9W1WiHJL5p/zdlSg9nctZqVdTtNEVHtMcL3EUiWetNF
ykV865B62+8zBr3oogPTnim4J3z/eykyGV/4nwqstf3KP2miFl5OT2Okwb7WBa1JGJNZ49mjaxOf
BjalzQtlEMN2+USUBPIW5xqd5j6bziwC7/heSCVwwDTLt0cNOoh0m3Ygax1bq5zQV8Nj0vMUTHjv
7t1tZTN9Lusro32UQc2xb2YTEv1KvVjuKLZDz6wtssIu4Q7qUiRZclIgfMTslMDxC+/Mv6YYan6m
TplmAwAR2Mkq8sGQJXrY9sa5zn7iKo99TMoBch1tUmVE61ysryceX4DMFEx2Yrj8cJ/0FxjAFS86
MRwzK0hB3rsErk7ym9iihSI7N1JUeQCVFsKhD9j0n4RZfxl3qMdknI+6SePwkNIqSmaMsuSBB6sg
s/FvJ7dIf+sXUWKHdYBxURbAdRdLcVZltBRQ7gY/RUBs7Ho4bsGknms3Sa47v+s0Du7n8Xi8RaIT
JFQM41hEWolpfzS05kJtwYdmlz/f7LQw3EtqM6vxfxGEu5S1iqanMQy2w1oyxOQYG1k+8rdJqswL
sAaj6fDZx6CXHyXoUHZdmj06gbHZveVTCnAWnWAy74G3ZddvuVsqif/F6PU7FoJp+dUZg+0/p6he
n85XmqnSTMoqEX/8km8EDwaCMVCEl72ZGCNomPpPM6pJafY90J51Oz/6ccGpTggjj1Sx9+0pg0wl
w1i6Fe/gSRU851dBSiXpWw5beTgES4KhC15/F+62nFhMw2S/LesEfDFuLWrknEpNU+rmTGkQuVvQ
XRXogJHe3LCDD0e+mP+rKit9ifOFRHR0aH0aUlHi6ep1luIpZ18OMUOHH97LXNEoz/Z3MFVCU1EZ
fVJo3NRaIEZ+/bIqJcNSI/TnY04UesWgy6OYUmsUF1rLrC+DUR0svC0yQYArSxLPOSXWpqhJ5J0e
7nSzudUx0b3Q2SCmVvryw8avzguxoytUM6xnrfYdoTZCjdlOy7OOouR79/sIaPGxsL6fbGPokX7N
3RLhxLwIfdSKEkqzVC5CQerF1gqtX5lJ/IZBXhpaCM3aq+ujfUIPEGXLHdxuIDnLVjm5AkhK4CJD
TFa+97orkjqeyqHtTNlu/0hX4ukbwamgkPmOOII9n5wE6j3NMAiLio5HZA4xJGhiT4d2wW0ErDxY
qnp6/4mGUzOCKn6f1nG/7uOQohqyw3cxoN3ix1cmqzCWtopKK2n+X/LGFo8zpctxue/GROEbxwsc
fHa7dlEiYzlO7UA5aV2uLBRlH1J4WVkktAITuAHcGL2O9c7gs8c85HtgU8S6857L5epQ9H9Rm0Sl
SS+xPil2hk+A1BJPmMOgFyeENetSIlNMp/SA3DKqJVmPMNbU65tzFCtxG0fJ1QGtLZZVfnivzCgV
khl/Ogj50mAu1xoHZdry25bdEM1AX+LqhO/CKpNaSCw8AXk0LjQ0stj7nH1L+V+4oAZlrJNcNd0R
UAFLbPN9AubUsugEXVpu7gknI0++r4gl+m3LU6ZeKiH2x6uQhBWryIlhI5BpU6xg997aW1dmfB2e
L90jnZ3CcH2j00TrlXdsO6rCbO50O1PBv6gcRDRWWSji2KbA8GV9eCKtXX37JavRQMzdVnMo4F+R
8ECbPyaLA1kY9e87vzW3JXxbKehQc9f1gzZGTXmfuha1TO7WlWA1aA/RVHAo59F0NqPqojTpy57f
W+PqPKuQ1UzbLnI/vsXJNcN4MZVuxAQ1asmrXEGObKZfxR0jLUfW1QOwNjiXXCKS3zEatwe90UAB
EUP5IoEQowgoi75Qbpaa3n4GsxkEeH+dRUdFdDo7KXovXsSVtxHLJqU/EO+nxWu90X94TTLqWu2+
q3JhV8UE42KrftM1htXceHCiG5wWUpe2S2afJco8/OrCNhQaESqlxFfGdcXH+kK9vPUx7mg3k4X0
oFuPG0WEarLe4Y9JEoL7Gt15Z7D4HosdibESrOHvWja1idgSTVEFpfeCII7eQssi6aeEtjlms+cc
Oa5ERvSQyLAGPBQMMMi8iB2pG5BdTLp/E1Gtp53ztAYn9GcA91tXe6XEjEEeZOxAhoKxd/5KISFZ
wXh4BR2QYnWTjqkuylspfDEBcHpmVY62pciIBRSh2+B4nUBELGq9pgG8ZRFJ9YiGXus8l+7lDEAn
kGGacjFJEEbjEeaz98c6GIGUOUL7wIQP3Zt6dxDrf8SF2Xq9CiMP8zB04m3Qsx+HB/2iWPAlIasz
Xdq46Zyrvfh5K5vkudoGBN1qsg5hfVZ+fK0eO6REf29yvBjBxgOTWjmVgAsgQU6GCKsgNAZLwg+N
l22MoVwo0pXeUyqcJcfICVM5bRm1RFh7ce7APBX0Rmh8bLK3RPrin7YM0pu2MuL6vk+iZokV+YxP
vdJBLIAQfxb31921kRG58KqvdoQ8XkVA/+Q5kPb5rebhLpVIt5AHYpCYdH7/hbv1RPxZrrHHc4he
0CYYQV++d/cpd9d/wuDjIjAQqQRHJuM3MIabD6Yr/golOP2VgeN70JdRoDjrgACKE/Y4MRTASJ29
Ms6i1cBybnMli789bY1XF9eH4F3UHEEIT8JDZqxPDSvgIPGIDcXNao8f5C1I63xQxcXgKT/CrZsT
F1rCyfya+0uQdSuX35vzrsOZ9qnrNppdlnccAZgbl3yt56XNkK1npwTJEYdskRe+LkuoLh5TGO52
OO9GniaNydC9v7mX9kNhj4i3A16/KPvtfn7gd6YzbKVkh95V4hMLWAcbj3jF3+BPpaLjZ9moRRSJ
aQ2Bvk4Heroe+RpaYXETavz/dCezV9aAD0kaEILukr/3Fy5G5ZyGeXZkDzFziafV9yyV1i0nN/4p
PX5Fn0GDA9yML46LJq44igc7dOVjfisr/p/tHvPPLTT4bxIkZYTYcXm8zsEofE7P2lrh1p0pXC15
PwyhdxUtmQp9MmmA2Ruv5rxL5fKv8JSzRBe+sqRv3nz6rNUf5aY/m3R4tsirpr3LK2PlfaxFVwEa
EKhGgVkSZ+rDk2pqGES/+sqfT6SOnFQ93Tikm4HKsqt+0o6Cfb2u+Z3OCiJXp4O3wfdC+8ytbXK8
Pek1+Rz61hyjvVKlmr9nv8Dm2Xsu5doNe3zqEbdKI2CN6rI/MkMZ4rRsdWNHY+G4w8PJlSJnxz2F
uLqfGmuykWOse4q6zK2dUYKmCkE0BjHxMZbVK6gallmgb1U7UY9fvrPIv7OJnjBclj7wjH5GtRM9
jqX6lI0QgRRbelECRv2ZAZ7EPfBEqOl9MroIN2VisFnU56uOCilzrgksUTDIlpDCyCHAN5MNTmhX
itGdPSLbfgKUBglJqRqSJzOTjKRa1lBh6Rqp2uAfVp5NdwdIikyAv8/atHFirj/1REg7cEWu4un3
+0Hq3KlBTYCauSK3f1tjkBgNbjoxyVGDbD/u9rNqWQSYDwcf/hFPN6t079hGT+HeZ4vJhUAZbgTx
0Cr9eRK62j4gYoyUhQmw27MLFDFX/2PKnUDSAiHrokqQE35Fjp+y1hOzPkf4/Ko9c6+EKsaujrrz
fNzUil+2EjG9+oP+VqcZlhWXMsZ/50baLok/naaFDWl96DgizAQanUxXQOEH2UElWwA5vLaNnPql
DiGWclvkFuVz+UN34frIf9WeaAkP2s5NJCkcYrlSfrzsqlS/V3keQ5jWFKeZBhGWOlg6MabyhQHG
nMmPdpPBdABoK1ObueCErG7Qo7ndhO8cYjigvxqNUtswi0JV3t2OrTNk1flOWPQmmk/BEmnoWVGn
gP5jdss+RcxwRod8WRRkBW+5FFA4U41+wyAQwUift2h7evxE81/pnrlDcZpZzQYf8e9TTNL8G2R4
uc/tIONjeIamcn49ixlfxuA69uVNDMgzBcpvc0OJWwk5LcXNsxbpPhSWITJSYapdvBn1myNrTHFQ
H0DtCuybTzJgHFrOeZp/mOBIXkcziOxG3oVqwDlPNQvBn96A0OlAx1y9MKmJia3dLaHoP87JSSoz
NS4YiIHbb8CDhm7Uc0xW+ERLQtvgsRccuSLH6LklxamiOdigFMcfFXLwaCea1wEr9PHVgxoLW04c
B9R8Q/GYBBiMmS0sQ+5BDmOiWKYnrjut/UNe940GkoMn/l8WjVOKTOsqipFmCmqEYQXHwtAyn655
gzl6dJMX14XOUkxQO6vToisbRrQM6rqaXyGARVCn/5rsdBwLtCw3Z8xPWOLpSudbiywRUlLmQ0S9
95zC3e9GeasrtB21iDGlHqNsXRAlzSeW+WKg2DGVFi8cS8gff75xtjitgpdp14g9DAWia44XZIRq
63i+QHsE15dvC+ms3bkSqRfWpDS0P0v1NiBJ7RD6MIeXJI6/ZOtTujqcDgvT6+A5EcDzZFJ8uMmm
Mff68a+3JzEAMdfjNg5y9t8O6VhFnyGZ4AxATMtFo7F89UnkBurBm2aNVH8XvQkE6VMz8fXQ0B7S
m/8ngtmwVRt334/pYTVsXyvoM8zy0dEoUan8LzHiIiUrSzYkuNb8Ew/8hcVuGQkEQohM+/U3WxHq
jV5I/xzlv1/58f15P/KjF9ZOgCJEmJGZC2ipsyBgs8n/hM7PyUxf/CYdqBtBTG1/E6scKy0SZSOr
u7kpgESutQQd5cd6zmol1IgVQrYmpOo4mE2HL0IM47GOxmAEHA41tKhu6U1N5OP6cc11YQ2JF5r+
ih+2MXdsHp1HBuUiqgR0RLpdKvOK6DL7KyshH3UkabZX/MFLSoTiKkX68sbBV1eHq6bsAAMXjyYa
6DOYgTmT//xFB0twoWBfedE8+MP94kO2X/sWYWuIJ055hN6M46FuWFqLsfw+F0xNflTaLMb6EQb5
56W6nrkfYvzApDdtfqAK2SI9Sm7yb+iKDb5Bbg1aZj2TI82TVwYSR4iVi2vSNIMs9zQ6VGbEF17T
PkNsOpi4WNIGL1d4sacoCMneODS0CGDznLm7+suZmIFri6J/ddkHYYxqZ9ZdTca1Pzva2mLfEteb
DNlTmRsMrJ1wCGEkJMwhIU0+BmrdQAyH1av5zPZijWOsRsUEL7cx0lu0et/GhAiejp3Is0RB2nFI
k2sXUPr2E70CVKe1edGuFjmzDHHaaLLqYJS0jby8+Yr3SwtmpuBXQ3HPRHAiXKgnrSSPVRiu2cEf
oBTUo4+n0PRT8PIBtxVc1cWCdL2eHnVGRFr9PvA1uChzfaWOBvFkS0DLy9a/wmGU68o9OL+Pb2Y2
Phgbse7jD03IxhUsupt/jYSRqgXOE2gtU8mh517G66yUET9WCqArGq1Y2hHec5I9E/snBrnMX92/
dpx768j9pfIdGHfoyG3+5XXhpvYcVy772UkugWygPfZX9NZOdbc/HLdSrZrpXqU7JQQV0I9vHBag
n1WFqsjU7n26zb+F7lyHHtznQtrwwpkIPNsq44q/ZOiTrt1JwAP5IQwEnD+hC3qVMZB2uGWYAuUx
JjoWBj+jxyf904JvpWyDz7kvduvcmeN4glIJ5mbYoJwOSULONyfYIJmfdNmMjiJIWwEswencmM4v
ljw56lM2LQ1g3qYoHa8LejE9mM6pCJOjHANtKMGYZyaIbo6BrbH4nVztf5uNaQdpaBOELCJH4/qk
aoqeerfbSYn9UrcnyLRzMGezFEz5lCCLy4riIiylCERNK+azdRBVz9rde2c0vDon39lVJpyUCICT
EMhZxt+lVM9LaEf6+PVT4QxGAQxrHUF+XQTokxnEWyIdWcHg0yheBsqeWshiTTcj/Fw0EVhzsK2n
PEoeQvaCIhmc5oB6nbpY8//8FnA80PeeFzmispA0oi91MbzxnGHZVXqmjwDRCMY6nb+mE7xnlh3v
YZ6S1qPe4se8DiZUiYsPwfG8AC7C4lQhE08cQrDfuCBKu+gNhxVCk5jXkipVOTQ0DlNtuCqIo7Un
/L9/QF8j0UzfE8saZWF0QgRwv+xtbI9G8PcIQUQ0adHqm8av3r9eAb0+jDeVqXTYH5YiF5it1Zxx
01lt30zP2gGfl/pmyhRRoOcf3uiX0MGtIIhx1zmyLeqioixIwJQ0Y4YoYQeYy7mhKtPuiXBOn0Rt
f1z/vIeIN/AHz5Z6LpMasGH0drGNWJmgr8MfX6JlVJOqlGdAUX9j+sn36vSL43P5dvumoYyaKTUM
y0+Y6zWrdgsFtuL9v3U5h4GkrJaP+6kKL9iCGG8TDOZGwdx4CFBTfkl0oNns3/0MP+Ma/1k109LT
HDagnI4oKsBISc7YFYvvNJxtFec1nLbsp/m2ZW3l49GfexplDbYVfN94pKHWRwIsSv1nPfUJmYx0
QT7xS5ddnABnFaIBQj9x01yNwmvPVHJqKYYlo8M13EwusyzD67ijLbXjiTl7hadOOmJD+YkZh06d
Uu/XKjt/m+1ILLbCi3iys8RCQo9vP3mFxUEk+1R250hTpGB8rzxvE2Pz4VX/PiaNvaOMjo1rHpEX
F5JRlJHO3+gfc+Qied+xwdTt0ScvnKXBU8SYYCSslYrt0aFeupshCi9uxtHEOyENUo/ynH6HE6kV
rzwSqe1pECk4R7q+sQawDO07ct1zne313Wl6ZHNFIFrYV9QHUxJzM4SEnNLUS2JRbcBM0nCvh9wj
Ag0FRtVCQxk9Jl4VFqqYSH1aB05qrD6wbKsZi6FqSoI6vVenlZvrdSWFCOr9K4QLVwpxRBIRKkZf
LE88mRCi8ECmBp3GPdJ+dap4IQY0m7oY3avfqRoHpDsnZ8nDcWJ/JmoxIMbCCkt900T0qQ2Obn6r
Z2JZqGHeJthLOPRBcT6UAXA7a1mJRSn+TIv3DPN1WzHjNwW+mrsIdUhWjODBFqa29vPQQOJxxIrR
HmLnjlev6uh0/mNJEXd9sqDgRksR6MuOIXwUHmkYdj3ApLX9A5Hb64XKeXelkhLgulwOKUQeL21d
tn9s/4JJb5QjN8iliXeUFNlC6Vea7o5I/zPcEc2ATkQNxjZuLaoLiAhi8MgCuG7oP6yAMQ92WWxd
48lt5lbT12CaSZ6fxuSkZOf8tpP0K04nTtwTXKOchyMm+hT06R0fVJTK8MUqJfDcCoUnwpbfFlEK
8HNjqdbr9FSzmjIAPYzH+qV7e11nPQjZ2/qeQzsRq3wsI0fa/UDvvURpnIVhDNC4J6D9Nwpn1R1v
g8RozFccFOMhqSGrNnMsN7ezBEzQunqHtiUyO2TwQ2lI1Zu86BtQM3kMZZkXZz9TgeKeyMd8lfkQ
U0rjUaBdQQNFUx1DQ43Fx35TwcPdBKeKDbFUxU/Rwt70KlJAxDgX2iAC/TA0JQFS+ruUlC26HuNy
qLv4U49oWSKcfq2M75WMD3j+2zgRsUcakXzU4eF/Gj32vWWp779sRGb8HPB5jbiu6ZGOBse6HsC9
7Tq4UEqnP0j/AMxlgUbmeytWDTvodgURoBWAnplxM54exkdzGPHBaXN7ZltGp2z2kq6d5MCJw5DR
iKhy9+a3sJKm99pyj9t2r3dSMj1t+A8Db4qglwEnk2/ftdXLvq4aDEW5X/MK4ArSBbOgpOK8ZQeN
4y8OFch76UgZRhiKTrYRWGwXLdDr2KJjcJUOgWAlMnm0xfS9Zk/ZcVNdBkHAKEO3LI+/2wE8jlXM
XtAvB4cXBx20PjoKkufGrI2s1OqTV6UE8mzeAdEiqeNbBBy8BmzDH76T7wXm3qP+yPRYw7rvF7VM
7wT4BJzFDJ3JsNAn7NXLswfbhJJXIulHuUfX+vhStFoOpm1ZVHPmjr33EJSXJ3XAHCKozFgKR7ix
mwS1+/4Y2JFCtG5DcyUwIzbUK07iRjZbYFe7mtP1FPsCQZjABxgJaUETtJ2FORyOVgW5ZYdGlCrN
UlMeZQsQArKa46R1oBIjL5pwZbMRCmh2a9BHkfPiZT80oV+uqsVEGgTU1ufHZS0Kz5DfvAfIYRhb
M+tngKy+tNhj7zuD/n8PzrGAmSZgUWtMU/JX5McKC0MI8hP8/Soge9cGJP+GIR4IzwSqrpI7CmN7
48Z7JtPj+dmUrfnsYoK4jPkGT217YBacjLUp8XaoA9ZLyiLkghkfNkQnkarw+nJXFBqzlg9CnLUl
D4eGYbxA2feygws78CGwDdWNhHc9wDcpI8AqU737N9SvJkQtnC5Gn1d5Fp30NRtTywkFQhUgvg4H
DErR/i8kmFBJhbqrsuHOW11UGhK2yRYYy5U3VJtr4wa3iDyluXDvQjOEZ8QQ4Cumu+DvDeGUAjhI
Hugc1fNFdWs36yRM6rGsZ7vjz2q8dH+u8glpRm60ehh10A3CnHzL2PbyGWzVUFWisrTsyO9ylFpv
n6CyYx6+YRNvTuVPkBOYF1q6kWgT+OxnkgFLAGzd4CA5dJXH1INUVfTiIx5Z1Cf3n0FXW1a/NWGa
2GYbOlfS+9Rkr1Ty3RTdkrg/1jXhMgy9y+JNURb9FKH1AhqMPxGWo7eMrrbj3UiMAHNuVUNb5arj
McHkaxaFc5CypO63L0WuG0rkNphVvJ1gbzDTSsOXKvOAefWs7wYWefCXaFilSQ+dBuQ/rqPLt3Fy
GBafbT0UvfczmavsBMGempfFQ26nSgJejtRPilsvXoxIA9Z3sWdrd9E2GkXJHEKij9hntB5vbK+n
hM7M9ZP+zEMFSdtaKyFKFrBNEXZmZ5E8Y14Dgx1Wi5r3pbUdgyyuLtYHCuEqYaeH1GJQE1uQsGsP
tDZQ6vHb7+WiUhDEhC4zWLlezc8NFVeB/l3gHVu9eRHLMwtglPYn0e+Nd8xX7iHRxbithvc4ZQnk
p7RVRRcxtPbwkmNGB81EWE0X0N3L0Jy1pTewvfhaLfunJb/XTnF6BOefp+06axPeSRlo4p5r58EL
ud8BOGoFnflyCd+YOT9dCcYO3wZ3QaWB/TTM3/uX9ZwCsDZm5TodDzIOczzQ5cegVx5PWoDK8uNc
EPKg++17Wt/qdIORbMGA6vmauR+ZejEiewMx50po7ynwU0BAzbvhJBmumoTmF36fN9Icyi6ikDSK
VdWpw3xvkaDQs2rw5WSzyKKKr41dYO/08foswN90mJNet9HTFpxmFp0T2xHzk9SAjn0Tv799wws3
/9wMWpIwYgRNCtu+qqCVl9PTvy8LpLMp76D32I9+pwE+INF7P1PY0XINistRvrG8MnBecp6bsHMe
MC8e44zl1dj5K5dGsy11hKpB9VIpram+QhL4NsbPBQHnW4wxRfYM9zMcpqrKoy47irPtarnX1VZU
lmupeIcrcU6IAB6OmbTFK0ei6EeXtgEDnc5pcRBq6SFS7zr+4HB4n7mAL8+rc+6QKwiNhYDUtFgB
dZoxhrkDGaTEg+Kn77bsaDNxosPO63+lfnbmE8f+VNuRWJDn2unscjNKBwiicmidDlzk1ed8/WKL
kIG11l8dsEeKCPUbvOLvm6O66bntFZ6aimg8bZjm6oMADq12jPEfDganhoBJ9tJIIKPWnK4I+F1d
im7qC0pRVdhwLcqN+Hs1cMjrJcsq8jGOz8i+LFbSUyVqM4bHv5YZl66NXPh/m6Z/I5nLqN9ep3Ud
lni/WRyH4yrdGaxLce3PPkLXkkRthBbn4zlOW1EMpdAexq3935K2QAL6aGpKOwLnbBjG6uPeJwLs
dDTGUOacCiVg6012j3k0FhTGr5uaXnm/L3NZxdkF/T7mRJKWh6cc0glpIznh7mJ6HJCxDipMhqNt
TaCL3InKxmOfSefDl3YzR1CiWyTUQ4cc30E+v5IkDQIMMMaAy/DMkHFzQQS61vGUhNdLy7XeKZn5
/amxbVshHndepK36wPP9/foQ5n6Q9Tm73F7JiqfIgZqSiY+pNfMY4nXxpJ2BK0sbBgEGlEY989n0
QotUoD98lsbmBhpzZgXH+YYWxFcNzqPID9bNcz/a7ABV7ouzg7oFIRcWkkct3QvyMuIIZrNdmBwb
x5aYBIKenUsG/gRWxLXnAF7MvuzCSuysLwEQGCZkampVMcI5TUecQAJ423iebV7YeXhIXivcpfm4
FtMpw71+VCSle6S0yEwy3qgCtMNodW5Sb6ijOfEehC7C6sB9HazAdumtR65iwWkIo7ji4lK9Wd60
hJHCRb/PjYTSx4QzCXF16G+6wThmOhXEwVACweQa7V3FqTSrCI0hTplAP60byWcoOgaT0qzt07CK
jp5Tg9iPdn9g+TAsng5MBGohtKj2vKCqSpnhOaVrTNyNkLqwc2CxKhLRk+zGihl7HSq/DfSvccdA
kFM00NVEneFeE6q4WrQCghlHcuEFBrOtJ43aht1p0nnxu3/umt+kE8VA7ol9AM/VPL3E4kQ1bwPq
LMiD0trBTshhuesQchiY3om41xu14Wfp2cARNtPMnxE4DBpV21gLvwHgK7NUeiaw6ZCUK5Xz7Pqs
cKM+LGK3ziNphUsrFwMaYfq1372zcWIYeHD6Pq3xlTmg0t5W1/xg4hsxJA/gyYchhAz7AvelLE+j
h2SoyJ2ZjvtV2B0fyN146sXodyw8d3s3Xc/lCye1TAE2DIbUI3OmVP9Va46AcDaaTqhvFKWoehZ7
twksvqIx0xmErJ2q5a4ZkrmPQOOumCc6aMDtNTZzvxnPr4j8TEP076WVtzOcprap+0blH3OE9CfT
5zgkEPVjIvrmHZm0QSWZSWhQ6tvZfYHHQwBsoJ47KWX1j3Q0ImW8s7BjTV6GHvjpq5i3z3nWGc8J
ldqEVPK+CuLn3qynqvPDo4bD3iYzM8S5DTme6n2F2dS3mn79w6UmCy6eafZyeO37T37toLf5VZW/
MB5QAZfCYKFJcwkBVIysJsaBLJHOd2jZRVSMez3Hf21dvhSAuv2bgs1vFc1hN1+lMEZd6P88/y5M
zVXEm86xp6ArPvMl5pt4tuy6Qp2lnj/ZUWo3VTPvSNk8vP+wEUL/GqUHt9OD5fhVQ/2CpIuYanYm
53ZnWAn1hmfYag/euZ+uBMbmbHPOJBh0Pczx1a+hQb18B3OHExGG/0vdaLQSZ+RGXSUvnKc/y719
2J+QLUv74La+BWokANca4cFeSBM53fgvukwnVR1mRI485wtL3Ru+chrG84T9wMxSVAnPOyPpCx4N
cL1HmmJj0jdDeEKWY7Q1pTCwvV2nROzjn409YtOrCUIvv0xVjRu6lXKUPHpowzOa3QUAzSYq1Aa3
kUln8abEhwSHrODj0dmCRnL12ZY4KWUu4/AwtM7EiXDQv9BhwyvgdTPyYawVDZ6lSRxylCKB7rTn
z5AJpPlGAuZhhj2IYCOCjNhQWk+O4M7YSVE1plUfcfCZYBa4sKJZa4vE2cDR7FRCpCRWxG+8YdNz
nHEKpFrLstGScLhclyc82VZ7X77F9abPBjEKHpE44AfxKGZYMWVtL6Iw8mpSALWh/w2/AqrwDSIt
ZTT6zHGv8jFiNZaNgqt4RvyDlGgAxeX5ZKK45C/9ydgWRit8OdaRaLOeaZcCdS2VPIx4zwh+qFyW
I7w7ODXaFE2Auta1LqVwpFsYT/P0eccHMo8Ov0AOClGEzKCODF9FN0RqihjMjgWN7VhiqVEWQpjq
iIMnJITEpsNC/4XkUTTAzn/2i7Z6vhTmO9kdzEP3+OiZ6C9hMgBRXxPKwSD0SXOgzL4u1EQGTS7u
G3KP6z13k+nGuHcdctKCqNScIKm3GoMeAMaxGZxhroHtnGbw3WJhbNdAx6N/BbTs7VID1zO1w5rF
4+lJNLrTTHOM14Fkq3m5VetBi9yrau9dEDav7wMJVncxYDPy1IhCjN/n/flV+Yx6FbdAg6PCtUKb
ovVrQ4WBb3Ejr6lwWWexiSSJptfQ6dzBVVxUqb3Q4AX3btKhG+t9q9CPuNrG1i0v4BJcUBo4FpiE
dRT850o4dpc8bEkMuCThaO73aA3yjtSd+DZJLfP8c1PtxHm0O0wCe9qw4eeOtralzvCQy1BwTKqK
qsPESPwqnPszTR5XThRnVJbwkX1tFd8C9/ItjjpvOza49eyN/VfFIXbYJ9EWGnrhbXRDDeSa8cQQ
oIJYHsNnq2W5HuygzqUMca/kbh9wu9yy9+dSERK/HyFRoGJjgO40ENvzI8ri0GBD6fDmGWBFrSDu
uBvV7d7V/fVKSmrsJe8IoOt06yYfvzppryC74NQ3hPAbTsHT2R06yqB1+/9d8yVwdmXIjIxaGtd/
fWsKxEpqDdj2hj6NzDail86RHtTT06eWFXRdU6w5F0k882jJdNjYbEGXjppE9K8+HpPUrY8Eczef
ySKS3kdTFkbDOK42l3HHunmrQplwXidUL+HEGro2WEVNm7EPTe5kQtA1CX7rpslqX2H+4koDt7TJ
gTScR4t72NWSraFCagX0Qf1PwIFCo6YzwWwTqDbbTVVC5/GJ/OOFlR3Un7vUepgT5u0V5Z3a/wM+
UznydSvI/H04FqqBHTxQ5CD0uYszOHWuZGG/VZI6avfa4mFihrJKLa8qi1VlLpIMAwwDOabAySPx
kPCkw+b4Vf7K7Pvl9LATLJGhHxtkzugpi6X7rUu6jh7Ft2SrqlJDSyGgGe1y/Z3uOgEVXsFbCE8h
3Tq0FNwffFlvLoFDVfnCGQFFu68dDZ+Zl8OWzUI51WcQ+DlOboefe4kBwLrpNLX1hKhDESagastq
MeTQjnWn0KA1jGBeD8F4QxmjVyCV/MmpyYpSwj1eBV7IDYojzkxcFQCR9sOPV9ImswurTQxtIX67
DgVhNKYbOqKU44SBeMbACrnmDyCUFSFNPcMmvNAhPOHbqhcAV5E7Zb2IWVHz85KheFB2eo8GZu0N
oT2QZmieDXP4rXZlE5yfbgricyTQL26ecqPWEfvqGnf4L7nFe43FuMxv/0OruPHvENBnMkHlyaJ1
H7682cKSzZBQyj7vZMN6FRiBl/M1qiPBmrMGOv1PDtzm7SL/iOOVBpCwBLfd4H9Bu17hEpcgAcg8
dfgxOB6bsMZlkA95jhLW75VBdDKvqF4l9A8bv67LWzJiBN8SELakO4HFlZHzWgWMKtxznwPNsfCQ
THTbYfrlgV5rTi3+AJpM+oh70uTbYjoq954bErh8fBbDeJ4zIMilR/2VkG1fi1QC7j9KST5ImSZO
jAzzG/DlDN8vlB5f34MsYvuc3XVtxcyMQaeAm32p4ozr3KNXJfyDYxiDYqzYSdvU10dyle9RvZFC
xmuGWHnW9B0xDUubp0hYBqNOKEq4gk2vrgczmFZrxMNwXO4Kloxe4FXUDfhLnSlg/mexbwJvZD3r
MD1Zmv1h00Gc0cTYgB3LaAff3aysvUj9AFkDMPRr56jeeObrKvBOMxjFKE7tmwCWW8vLW5gf6IsA
LqliAHzt0chtGOC5HQj7N9N7z7b5gwyz3E/r5oWbPEnIPxSnbQ1wJ/nn0UpYBuN7oNOUuh9uptZe
bGpvIi7jKFMYuFh1fPfcBx4hQlvE5zDNI2ohSuVbOPaqOCmNHfIVLe6syRSqEoAN1+IRnvxCTZkm
+t/oY2nrvAWXQjH57QyMAkP43iXv8vkFgyHzcFgf9jbiohVu2LZnosWVU+911PXsx6LJS/k8pGMm
vnCNnqJVusbe4rhDF9f3WFIeNLIAyXtB0vNGPOgIR4FZ2qkNIZ5opv8qbQK2g2cvMrPU1jRIqV7w
jF3sCiZ8n4IZIuQkls6ONmGp4Su7WQWMbVHqyaUYgvHgPqIOVm+0m7Kf4PZlLWiXEVW1Zh6zWIKK
zZDTcTMNuYPirIpBShlj/nO4h4s6YrnSAOhtkmeaAiyGzQcTdnP4HsByGTQ7mzAn7AGO5XYLUkeb
fJCAqY9lJK9glZhb/1QY0DDIo8N+KSP59GLT4NSBAcM8M/iM+45ARgB9NGRXbOjCzO1gGGdRpq+L
GyrCXNljmgb4vQ3rY7W8y0+69kqC+PtdEfOHRfn5z/xwH5EqMaYf8k0KSmXE/j+Oii0KExjnz5mj
pZ1ZepzuK8kzUKgj7rbv5g6aU2wlEQzwrfH6ZG8Acojoq3+Jk+p9AGSZ1ogPDmC73YfmsMTe9KzV
TT4WSnElljH78DTAq+Tl59HrIQ3mP8G1CAykM0wqNBKqoEqdld1KOyKtbxFKsSbc84B7cHnZHLx7
G/dtgeoEHUFCDvoZk53QPV5NnSWkDIxa9hYA8zapOi6BItIMY5XDtTltGBPHLC0gcJNQkDL0LTfc
iJQ1ihpVweTXdvz4I4orH+eUMDU1OcLFkAD7EN6/fi7S2A9lc2+7nLsyHBUKxoSLiInIuEwygU6E
U73ipUS4Vm+lPNJFfnK0ZCjkrWZAVZkANR4uHV21Y0KqjqfNXKy//amV9mpfxKqUYjvsltyrEzA3
tQAt/WdjW+3co7e4tBiauwyx7byIM5c/JtF0iPFbpoDc4IqnHBr/ttZ19MzGfaQfng/DSalPsUjP
VlI4RBkpnUyavJsNfk7BM53QvhGFdPqQQVsx4QAu4pLM0EghGTmqbqy9wjEvw76IY8X8LKo5W3FK
XSf25LfFzXXPXQbSZVxQZLiMprHFzEo8WkNyubUb+CmY0im45bsCF9KB1or7oOCH3dN633o18SOq
dzupOb44WQmJykc1MgiVtcYeDB/pKWPQQtKzcHGS7MP/z4oPMuN14WMYQKlJMT7q1hSln5fk7vY4
2RFZ1HLPCSknsz/vWAdUWWOj0+NrJRM1SxnmzYGbNKpyri8nhdKjysSm39/Nwg+U9XmB7aoapVMV
2G0q/d+whhhKxLpBBIOPQTGn9CSsroLKHG57SGSXdZ9lCIACRLI+9JJOUpq++Vdb3lbG3HslsjPF
k4dzJOnUMQB3MHCn3UitU+1LYLwRF92TuB+YYuDDE+dfbGyJ6KUas/XJPglFS5vn41kKPDgTgW3R
bM0CO1MOt8O54/xy37bS5SQ6WGgZt505IlifqBmUB7y9UACmG6r2HSnKMf3QiNnqvHHCxS9paWwv
GY3e1GKrb4WIsdsg6WytlgXRnNwnibhcKx90FoiEdjoijHLGF/Ge97x85JY27Wn6BEmWpDwYDaMQ
eWvPWbfFZUZ0ymlUOgJFlAA5QFBHKpcLibSL7YyptVhwsLw73twB8R7ay1y1T6mcDdDY7WD6cVpJ
W5/B0wMVkEdfzSFAYxj58FEGZXrnY3x7SRandC+XbokL4nfv2T4Vk5g5ti+yiSzJ/HcsMVzZAAet
tGuB33K+bS3gfk+xOt26Eb8Un8H+ao5bBEUfbBy0GjQ94o3PdU8gIJZx7s67uBhw+PjwLEk9ucy4
9+oM1Of0AcaORWU0i5vZYfG1SECgjiUE8iIJPFv7ydFziyHG5WcQPV3QF900vvOPqbrWiPW5bxV7
IGCVczl7CHPHb0g4x4hTfiuYakMRfEOMAVq99ko3qOxzJzJBaCNl+u92ZYrWXv5sJMDvStRBWuL7
rtp4OXh/fR3BZ2bzMyfUyMQ2YP/SkJIyEQbf+1kXo5qEkfTN2FxmLwr58/11iJ32Hw5vMZGgUY+g
Ci2W/xFzQWfV4NDGpG7rqNlqsUoqH4ptQ5K5KXdHbQzaOIyPmwkv849JvhgNef2yBLwBVwtsa94T
9MzHDW6T3E7nwdDO4KI6IcHmC8ay8iXON+JDCiWuC7IKHLjECx1r+jo55gV7A1tvyOuzWCWdqjOL
QJvNWotp42hM0BQeLjYcDcG3CLkxxaqGyeYoTQciKPH1pjiMZ2jRVELysrOH/pbsE2hkMUZ336PC
qU2CmvuvfVwKGhQ0k4pTEfa16Eff6bHGbB+Vy0EMCu87VOQD4zGyO4II6D4D8xhEGFA/MvfFh/1C
C596qd6irwa64FS9Chtib4fYGoQql1ypsCr8MeQ1JcJ+/rybbRbekvHc9JHUsKLhPMS+EqEsVNEm
T33Ewss8fJX/nVcZivOw2pHBHhTyb65Kt+/tohSTZGCcjpMeh9+3nw4iZ23vMoRx0bzXf+S/v2bi
AZoNy7seLB5jpVvmiR33gyzlFb3GLTBsvnHLapIDQQKfsPMg7f/BE83sSPML4J7/5akFyWd8bN6B
fBTUfqzZmvOzoWh2Etm+Gv529k6JxRCDG2v0iTX82d7QhNb/ZN5/M5bcqt8hld6zpwQ+F4zKIhZ6
xgIc7QgtnMcFfQvHHauSrD4yE2EgfY2KN57czMCYLX5Rkvzqej59O+LvfpIrIlr7JJh2waLX7VcE
6X/ocLEpkN7xwydZ0JvT5t2t+panKFTDe3rSdWN/rcd+iRtxJD6QFosI9lg9jF8/u0s80XtnjcXY
82zx+kPoYUDZkOFxJ/PJOpFp6uHn/TH0hneA5RzPaF/ne0/6aXn+ZWPLFY4v0VYLI7INGdEPy1Pb
FPMq+toERuZW15u5aA96hw1YuzhmEh+AhhO07iiE2yi3RJ0BoH22kDSQ1qtnvb4kwWe+iC0mK0O0
W4aTupXUBCeTtiMvWk970GW0uURj8/Jb4heR+Wcw2N9lHLM2+/zPvKr9XIq+4ivsGYZpuI8Cxry6
Mn6RmeXzMgrnXCA9b+R5TMwn5zoBqyhh5kLt6KRSr/FkZ8iGuyfA/axRp1rU5z6Mqnemx6krxAcy
GS040WAO+cQpsXCUOoS6sOeEtbmmHSVCGgfMTvCj2whsHVPPBAJXAMTqD6sEp6WNnV19gmKhySdL
GgjZK3ojLYYOKsbubnQVfCt7I80TCrGzLFSTT3woFvCEp4Nv0B9+97CTFXJ/jai4FyJ4cE1KNYnt
zszJPnpfN20gpmWpYywCRHXT9anK4U5AZzadFq/5W+QAGwlCrforcIIW5y6E7IU89z2d9J1X++3r
+pRLLAxlDzUiuef8vmJq7f+GhOjnCxHwjO3Nfyr2tnF0VmReq+mm0H+b3tKDolg6snLQNVOBttBa
B5uwCjaquk+jrCO/wlNvRY6mgiJr50rmsSKKhH1Lka8WT2eXllQeepDGSqXCw/l0yWSDheIAAiCq
3iPhppQ9zY4I3zae2DQ4USDILAx0sqTRtzuddA57e4mdw+WY5eeGGY2iszzI1xR29/HBHGna2mKE
GM0sDIJOcWZsRHrfXTOKig8Joaaac+aembsLvmYr1p8t8M7frcnHYm5lChN1wQ5T+7qCk3AOuqgY
4AEZ1Z/NpH+eZ89ZvLtd/lNDw/L2hn1HuXuLE+F2NtXtxzKBkWy7r0z6w5ddMx+ysbSOEx8twH6u
EUiNEDgBprt9wYwX44EladN03VSvTHtXcDreHV3j5BrKYZH6Z6xiuz09EP05LGLw6L506LoZvzqQ
Ets50qxLoKcnwp61bSHV2UMm26zFo1/k8EtOkV/lkzmVo9yA1ZAGQzo8XD2C3A3vquB43yB+KllJ
NxyGN4sFmLva/HQ8Hg3UXzhfV7jDKPRQHbRyO7pSaubU9Z9OCsHxMdXFmLU+CKllTR1DRwhtGMaH
0/ET7qv2nJdX5A0nBEkmvg9GbgL8Lvolwz07xs8dLuhZXf0/bLXzfbFgz8J49mDgJyF2YFSuwuu6
d/yzsIe6gfrFyhpyT6ATlkb7PDkycunUhqwnY1VQgZk94i5gkjcxeul2+SB1SnOOlq58HIhdOh43
6HRYSvn+gaM+/mJnO3IIvB5WoJQBnEIdaJZ7HozfkC+jaB7nrikC1hXlOTG9TzQhOLZA8oksBaRO
p4dLZE9c4YCVutxG95ZNdDvt67vMUMJGLHroqHYEx2w4QUUEY5fU3EDIaDFh1S7qWBRhwdMfHPxY
AoDhEt/+ES8ONAaQZIdO10mQ6rIJpiHflKgxqyiIFEA3OrWHgA58Md4jZUK40EbmM7CIKf54i4ZS
7t7BDbUWXVcRMD8SeZpQzggvEOwzwXiRFybU4/pxsrQM2U3eE4wwD0yg9kkchTZIgmPeLTHPgXvQ
FDgLrMoPestXTROuOUHzsfNy/m6tVP3DYFbKko3uWWzdkzZyWfqA8qmMsG4kO2X2lxBQj20iQG75
KMOfpXYWnb7uDBhQikdnzaPgja4YerwC33fmLjHdrXsWFohdlIBoxIZgxJrDawmAnPJ8Hu7d0/c2
HFKPoXwUs64C+VYEGZ5yEuapn3tuwfNlUocflSpTbxsdYrHHN0ob0kv1WSu5m7bCR2OM5hR3R722
YiI9/eFG8L+nq9o2V5s4XVOM8QKH3bL5RHDL7UiX6zWY4bAEngJr3Ad5HONUoQC6r32Wvx7dEuPg
nQOEvfSYcn0AlctI82uvtZdN+KXqSOie8NCPc0zwxYAYL1UfH6dtns9rh4bzDzBzBWm1nBDEaJcW
g78jVdhxyzpN8huGCUTFXYfrqq7yih/bTm/lIZG++vNnH3oAbE5uPOrLb+gRrbSO10ZiyqpRHf5z
h6kZAhV+34Ix20Y5d1Pcdj9B4nwPi6vBMhP/GyuI9kaPq/kDRxLkauGeIZXJ4n5x4DrUguHuoigI
QpbWYvhFn0fVhu+8YQo7wDFy97DHqS/tBW8jyhmGZRX5NMB2NmyCQvkQA0N/fjCGCh+mzit/9pz5
Tn1XzMnbalLCk1lstx+Y5gXgsWgrDu5208NHm4oH7GICXwS6XE2QQIWTEfphaIFWy6eAsbXYRSr3
M87TqwoROQnbWYrBJfy4PlLtbhyUAHZe5iseUKk5U1flcOOmNKqSktzeQx4SKCf01WzRnfJ2XDs+
vsohcjFQW4EBSrjXqyG28fF1b5krpZ8zW3+QUUi9TgmwXtsBh7BVmXo9P24/jfebCeCdqJA9NjmI
eNjHM+GF+/ImZPXGdNDm0I1L5forTCtz0MMhzhKO3Y6TprZYjqEEtl1QiZRUaoq8sD6F1S+ImrjS
ijl3AXBWf8Vmki0mxq3wlWo2fNFjFK48dxxHb/bKBdiKKvx39AJsTARHXAKkeCYa92rJInvyFJUh
hs4Sg5xMyLg9qJAIN2aQ6SabuhGrCyQC6+/1m1dhznLxnZKl6LLi1mpwgVn71l+acXL1wc3V/eeK
xGr47yraFQNpjn0cty2a0nPtT/tNIT5HO502ku0aZvLdoBNiGMSsXprXKq9Btmo9PiSqVfjEOz29
nWS41C5M/2f4X4aEgVZKnTj0+dJdzgq1Yr64IEOuirzi0MmivDSD3MN3Q2NBEplhaHXoEgt7VQU1
c1bVOqD4+Lbk4VkbHmMSQtw3CZTzB8TPXigr1viWyhTIHQA234Yb7s90JPX5E7AXuxgrTxP3B1x2
n9RRHtwebqMqAJQf+gRM/tGJLbaW65hQIQp4I479fknTT1U0v4KhWz+c+mXr4UfwBeExQbC8Yv/v
PdE9JyOKeQE10nDbrDdC/s3TCQacvuEBcFJYrl6bimFWccO1AXDzSWAUCxiEa1AjmQeXTYjI+yAN
WQKL9gTXZ+rC8qjH5ON4U1wUJsw99WoAgwFaX+XEhi+b5NpFDcL4DEZVjZ/VVXo3hi1rKUEMAPD7
8/uEutSBt4unCMi0jwk/kcvZ6S6sFQq5vuJBjXCDSQiV6o6F3yaJXp2L+2WGEvr+lO8wxbExgdX4
q2hn97ZVdSyb8P+i6CfD6LKRZ4X/K/lxtooZvSGanweuoTEFVNLN/LByyTLjcwn8P5l9NA3kFUpI
5hECMjncA9La9yT8LBPdo1B820zZrOJq9rcTSiKFviS3YL1cIFFHBbBs9oZaY7aVYE2/guT+Os4/
YcU6hJgUkdesYAYWevYntsAHF8CaTZGsmyXM5gf8GFNhW/3HYc6lzLwIM6ZOoLUfyE/mAx5ed5fv
XaJyVe2HuOuJgbhLvLSo5evGc3T5sZH5frHJCogQGE3tGO64st9D4Y9SAgIw6q1Frr5SKFOwQoHg
Za2zjYJ/r+28AXH4tLemWdZaxzo+G/jL4t7J+GVocvku5nAjbh5dbgOP/g1do9zD7X99zhkyYwAk
6p+WY97QVz3jLro43QnlgIVRf3QYV200zxAhjEJMq0Hy5MO40HMBF5j6UBKQBYX6ZcYsWux5YwRJ
U/dxJIjLfli8ZkL6RI/5AnU+nurpSiw+MaH2bvf4QX6sMVTBqEZJCI/p1sf6EZ5vAD7Z8GwWS1tv
g1tWFjI1Odb+g35iNrbjGeUTQsgf1lCqM5mQQa5ZhoINyeS+pNnKanK/GdEf87nr0/RGtqNniLN+
YQtKJkr0x1xHaYOvR5lfTAbYNM14uE38/oBx+zYmfwuhXuE11sGwxUJn871+uxjWyrZFCeJ9CXm6
pEuYlT7pBg66qQUx5VtIbfSDCNIaynpU1c1nixADNEnwzbfsddheR2la8dGAiQFcYxwOEs/zAcMx
evZBKrlRITz3K1LwfUbOls5AKAw+b1Dn6MGHmRwVrzZsXGeVUA1kW9heNslExmrWvBSq+LDErYmO
PnPypj4VjLXzxnKIcuiYZxxMFDOy7jb7U9N+onqGAzB0FEnu8nX54psm1T0XYbU92cK5Q8wHarKn
IDk7h6L7nxKBMJhSpE6BpxuHd001ztZ+YXCZB9u13a46EqfjUDP9OaLs6ATLtNKoe97Ytz+b/LvO
oDk4hUxISLEq4RWeGQwdOTVtsJV+UTe2fAkTZp2fJ7WRrUsGYNp+c18HZNPWOTXAX4BCyFcvnJjD
ZsTbN5gb7L/Np2LTHXXY/md69UvJf5iRL5uaM91NMfkLBlnVgxFdlMV5oliV6hOJt0Nk2lYeiEcu
afZgDW+vGNtkBZulX34af+Xkk9/pWipNuK92WZZHfuTa3c/UpD5QGnLbUMg5wIEtzaE/Q7exzZ1Y
Y67IAPS1mUpoYUYDkDxGcCV+RQi+8DVP9UffLLT4TOOJuKcjP2xvz82VpoEI1pgvidERuBbPQQye
XgPPsVFIlYpAHMaPBsHDEbxEzvEoYaZ5NI/OlX4vPp9TbHNTNCoUzRdajOigbuGfU1uzMCs+EDIp
n717sG/R854ImETBrMDVPPEjGSROX+o5Z4BXm4qrHmMvUUj8BpRSN8HkkD2zoCjWc670jlXDh3Uh
4HIHxKhsSq2+qupUaLLED6dNICgd+ga1W9wQQCUg+/scc84XflNfDd5a1nRmVhuoaBeuacuDrk37
0GJ9rFT4GH3mNmOVEh2bmL31sh/hsZnyKZzyNgQ6q3I/LS4Z1RTyWcdJZ3GJHGyHyJ8cfJQeqIKa
Pij45t1fjTwAUo7hZ9voSG9/xf2UKm0u7rFMlqBbN1vCRIdnSqRUy8vcYn0MY4jnmgCRacbk/Wny
u6T9zm7Al4iEpHA6R6LcgO0qsJB6IfrXvJtuno3vPZ2LipyoIzjf8SycdDwhPfRM0asoI79Dz+s5
KMZlSsC4DtprCgmUSCOk5Zke/Jkj9f0RsYcuWN7PO8lOWiNIrKyZ1NQ/vHkf4cUhcR3PgS20uaSP
TpFTgs0C+aKIdWoD/0yQe4LXRP0GkKUCbAA29K4JJylPNYQpt4yPf9etr2Y6981jOVg0Vqib3B0h
clphvASLLs3Se2jAj2fPWs/kL3uo9MpmYCXSrgqQGrcrvXT/p2tugSpwP2Ia0Phk4oT0E1PCt3hr
23x0pd5jwKqRvsXkV2vMiSq3M9KeT0zHqtNycILJ/COTpllqpqC13sMprHNK0jaEiBVmpRT9sgOf
j7XEANArWnfLcFzUzTDcKqMgq5GjvWOVAYR2oorlFWKyqq58UPEfl+89u9SxN15CeS7gY6+vW8RL
O2Ycc/q11GeciWi39na4L3n3hmc+PYvDTawU/KOaIvDpOm/wtVrDg5o39J/pujCPi5D3J3LCBEbF
VD8EBTPrbLoSMxzZ45kzYPGoTjKjs1RhmKDghCYLY+qFD9w0C4qPAf/BUSriS7HLjbf/Imc0PuAP
sfOqJsAYD/hS6W9q4JgKfRluCo4MUQBoGz03IHqiZCcm30robGrK7lSRm7fRo3I/M5Au5STdWstV
zIBARwvBeviGssK6VBFV6TPDKP/nNW9od/+sINtdewiEQOuUm8ph9XJ/J2KEUfrh+AvIHMy15y8p
JxBD6cClSWupFhCJUDRj7BTYXSwLSGxJeM5i0aBYeTXIMbXHzk3WhlyGi6mT19v5KT6N+Rv5wuGH
nRDbyEcbCkS4gFPEfEpWXK/cbZllXskJXm+QDnDAD3SoPpxsT5TcgyEL2GO39ZEMg64bhqPIVTXj
63cGlvPcj7mQ5fzpfs1z46X67Gc4TK7M+YguQvqDHtNCDHLdTcC3SlsDV/fLhzP0L8EsV9pejOYB
DiFh4C7uTDRtK7ZkwGyVNUKyt7Go1t+m1N+qJI3x0uIBo+PVdinU1DPC2kqXL+Ks36QtGimyV3H9
lFMFHEX590VZXi+dS6uvj/NBiwhf0jHZP9V8u50r/HQHCLqUg5xjryVpx74FuwaA0sHB7SWXL3om
WVCpoqN7imxe7t5+KD5Nq7cxqSkB051KOznU+Dx+w3Nkr3VXcbuGRz7FqqNCl/b1UHXt8SD+aod5
FoQBqxe54JrlfJKfpX2WTkCvcqXSC4Eh11wc1uKh4CXDiHieMjEVVG7xBnbcESw1ODn5ASzImrlJ
Cs2wycdWUsE16SVAQ7UASdCF1EDbXvfEzsaIzN9odsBHHmca3WUuYI5hJO9VB/lORa0aa9+HOiJW
ITdcDA5ugQI21K9/IU51faWAGGQR79nctusLCPNSPqag+ZgX0o9Cz8wL1+GyVOiX/qKur03Y9UPD
9GcYE7Bmq5BqVPSaOaK7rxBDOZQ1mY+9F2PZ/5nE/IuGazzsHCwb6+T2rXC0zy1fPbv2gwerWc6Y
L3mzdGIS4VayZTi6nQZvNHKudbx6UG4ubVqJNcB+HiiHsenH35KtLIwLtLKCEHtKD12I7EkhvXUx
dhQJz9kNXOFnBUe1bUpwsNXDUtI6qv7j7XePRhVFP/YC2cKaKQQYuBlGLpu4DhHTYdbzM3X5ROmC
DtdhK0qTdiBXBL5xwjqrMWrVxiOtYQtETZKGbPgwzlLpZrP5hZJnlYZ9F4aixhsRgFOA0C9hPqhy
gNL5ICxiwfowvqMNPKrRa7xUj1l3dY5r86vsdyJLSN90HAIX+Lxd6keHJ1XFuJDdSDtZK0D9ab6i
Gvm7THiQnTzkOBlekta12MGsJZqtl7mYXHMjrCZ4FrbPNpxy+0FYNmR5JUu2mNlJ426inAmtrEH4
zcltHrOBRIpq7lk5wPOHai3HAmWuaFQT8IQYNpxM9heDmGvS421UcaYOhEEQIXWz6xxKdabDLZ/4
/2dReDA9JnJZ5WCsqIBCzT0/eHfdyclMFJSM41VRT9RvJro9DaiGP8MGdeIwFtvA2ViQzKwFQXGN
x3DYc9Ly8Y6SecTEk3OhIAhVX54fA+Mu0aEu4jxt1jK/KtMIYZfOSJ9SbOCNfcg7WOVkWqF51+5I
AHz+M9LHvKTo2wZDsIVDtCOnJmlxJzck8pI5426k79qmTBocTLwMWtaSNx9eBQ9zeqQ7lvxlPxAw
P1IkZ6TS4FYAmCy7wc+b4oJLsbqxMNjLQuZ/wdWUzueLIHINbgwKnA+9qphRil6vJBrAkgE+iF/y
nX29Mw2MmKjGs6VTbPYlXBBDzKvj+hn7eCp/Z7cjW2P47axE/3KQCEguZSlz7CJcQOyWUlQSTCFq
oD4RldQtHxRIrJrpkD3Bastuw1re2bvVPf6h14nvoA+vq8JrZSdUjvq6dnJ8BjwMyz9NHkKIU5CM
iGMLpr5ORUWz//FjsrFx9/MwbcyfL8Vh5egKFHeK+8ithRagQwtgSMPrnuRhWycdIWr1tkAjfqJ/
ll+Ifh6sjQfUJZb88d7nvxiMLPeYsktZRG0u6+Do5e2Znth+4Zlw5t2Ml/F8oTNBsUqULt0vXvSC
SfbMcwFdonQZHins1KPt8Hv0k5MMpHTdQpdVcwbakTCJf/Lp6snpRXHXsPhUeNYdWyvDBRoH/WpN
MSATfN3wXzFSI7OgHUr9AV0zUTFy3KR10eQNquTmJrSOqPMxMV8was1WjdQR4GeMIkyT4DDVJxGH
IzV/OkQ5FAcavvOr7DjSDF8qeg1KKBMFkYXj0nhbAV904nMTxdT9iuqF5q7dWnVOu4DJyoZdUqzK
SRhjMkPMLvvIcF9yQNAAiw4SHg/DL0hPhynlKTrbbudno5MIcYwoZN1U4Cjsbshn3NsaB/HUlRNr
pZ+DEBNpXo5J/9m7IAa/Vdtaz8nUyLOwzzcXzvmxsTW1DYyXQxGf5SpFwOSS3d+/h3q5bAxVvpa1
Mt3UBDITrEdWv6lGsdXzKXL0UCLEgh/Sw22Q3I3EewgYiL9RSSUBU6m6dvqee9YhdCSFd5lbNdgL
qJDw9Hq7qyHn+DH17XTeXw5/famDU/SobD+m/nEXHatdNTiyI5I2nIASSuqTZL4fuSfhxmOVkeSV
rMpO7tx/c7oYQrXzT1y1oHNrQBTUOVzoV2ha32x153Mv8DWMgZ8J9QCY8646sKPzmlSRKUf3c7TX
qQc95ElK8zoWv3KvSJ9th028Jj9HZBI3RxsRoOf77MmmM/8q2PrhotI88fskEi7H08zij1ncE7MZ
Xh/LNZqUuO9bH/iKtp4AYJz/8wFhpmZw+olqrpKs7Q2No4+fvMiIaxlsrdlOPwf3pIvASNfvTUEY
CR9lcRJyXQcAYhP5699eJA3yOgp4Cn5aPQNxeMRVfQvd16slIakNHISghO+vtKU7bKCQmbUK7pjG
3Gcj3YDsiG7PGTrBXsIjy/iDIFL3/tuqo8tLYE0zz1PPHb8aJylAWVaMdaWsdTcbRVbL6pH9BJ4E
E8/RJCNMAJd6SU6wTbVjy1BUncrq3aN+YKGa2wefuOvcIsItB0G344hPxww7SoeVqHsb7JDnEgfr
o6es83AetO2y3ioksmlz/nzTYqoLQej9XWsuUvAnHWoK6UsUYeOAgnVAC1Wx6DzxMVzXwetC05zO
nSgqvCmLh7HG8grElH3N03juGDq9z5npigoFLVmkWYUE1ug5EPPtSenGUD/7PNK64P0A6Zc7Fwzk
/UR/xaiq9ZrYgxQRcSFjeElW3ldF+44On1muS75IOi4qmMbiKVJbvQ5s2/CXXCIWdaPBxdwGARC1
S1T14gGGiJR7/oy15SMBz8J9Hz1Tc/SxO0XiLv9w1WS97v+qY7ae2Cp3m9nJ/8On07f8lJc2qxMe
HfdIawHh0j9+zAjFdgEQEwrhP6HSwJQT5Sg8wGquCn2rEuABWDTzDdxJY7FwNB6O3YPJpjt4jbTj
lvLUEpVrapRPcOr7oRCo0uc0b9V5dB0uh2P8eUuNO4YeWKuKsbEKTpTuj0Mwd5GLLSOVesELXvIH
TRJ15lZP3os+vwsX3/UZbYppWt7chd+kY3t50jtIYNiJHYn6wEctYWYgzTFDBgPGFuN+C5h+BrVq
OQFTjjKqfApX+Dnly59tSSYBj29UaPAQsez1P/TwPIg0K7cL1GmSwQEjsdEcm1UyFnpRGdCUrcOW
X3iRscCuVUiAiF15kHpw3PGvixham0YD6fY+Se+l2HyXdGMhW1mwKCG49sxN9HB5UtZLxxWUEYwm
K3tKaJASlrwlstsBVwEZ3zkHcLUTxG8e4ctNgMMG5ipzsHsxVbqILirzF0NLj9utWCQFXGIQLMlQ
QZ6LBKcBw7IPpCMfy3YRFi8mgv38phkaD558/8NRqvyO0rB6d/4x3YIY3vPqkZoTDrEoAC/T18Pm
NU3rx7BIr8p+/1B9D4HSATJTiB0fQbo25fUrgAcUfwKdqkVkABRY2ip4Mmhu4WoaXnHhbOODi3ma
UqMZSrAxAvaOBq/A088pEEmiq3U92dKWu+CA5VqBz6DQJ8WNADd4cAkn4FK5h8Rfq5dfohiQtp5P
99flU0OHw6nLPZioxaxWWSqsQ52LDjtkqiLjxw9D/8Gr/Ze3rEiE+/P0okzWlqAFbbRMVFPAmvgy
6tU680RkjuD0aZscU5WrTFOXPOnof42HGx56bX1B6bg9A6Osx6sBkn+C9LXzdAuJJ2jR023vY1Oh
lql74oOPmc5z4f4y6aVq0JxC4vI+emTm8yLR6RoNJGtLW8jg5Bc+3Y4WdBGtQ8b1+QO/7+AkEiMQ
txELWIzTia+/eIWHvWIugEesuZeFqhiZq92vSJOFSLCoq4BxfP8QPctWw/M1eH7TIo/shURT+XOt
7HBKFJgTX5nbZZLOsv5emd7DGm+lrelYUtNnCYOzB6lFUr4ESxgAiZFTLZL2rlpshlxfmZExDFPr
EeRCiYXU/WAfmLJkwGSfNrJklALRIAfsIqgOhw8/J2nR6bjhi9toPTo9GTEnqIV/GsZl4xDbMdyb
7lzLaCrZFut8TE82mAJiQJ3quGDcP9NKmxxAl27OCj1s3RIyMdTxx2yxEXXPck6RW4isf7Bu3Q7G
hj7Zl9lbLatzZRMx4thbYb7epJ8MXIW4MAmmhz8KRumyEhcWU5juZIAgfVpF5HaIZTwB4D4N90yh
m+CZn+qeBUvChk4VaiaMLM+izTxDkLqS+XrNQBrNKgdsgCbjzGqe6UzHZokMh/GJ7rCy3rG/BMku
8zwPSFM4dngO1ZcXOiMKfjpumnmcr0uF8n6iaSRZbUCA0r2Ets34rGyvX823Sat+Q8MTKAyu9ZW5
EomNaaqhxC21NPBtCbD3iN4aApNgheWXamCLol1aE10gPhtoO3nQ2hiEgcS/S05WrGdIcjY+nw2Z
NHsso5Ixu2PgboAV4i47bcIDQC8Wqb18hauGDWqmcd2yQxw15Hk8Y1Y4iFv01oJP/kJyKj5Euo4y
rNzAqeEfIqGuvVz1hkbBSnV+xqfK5BNMOTms5JVbnLumNbc3HHbfjZV7TIwul5W1b2lKegxK87ht
lSSbrlUn55AZtSYACNSGtVEsiXwa8XuylmI8nmediGYXosGd/DDG5yQjVubFozVIIxjypnENiaiW
D4NW4oGTx7X7hhKXR5EkReQIc2l6dqiBEIW6PkkWi+/QC7JTa2xNd23rZXWbcAAMSwLr8A8DKrsw
4vfuUMaeJRgtrcvl4FvJ93UJffcdvpygg2qu7FXG6LFl6UoqQkpgC4nORlEofKMFu8+q1PNux1Tn
CnRbPl5Mrji7Q8K8A9ifkDJNgv+SuMvLiSIpzHSZJzrv0IQetvLZNkiWZl3O8CmXzeEB5n5z2qku
SR9NEcOd3E9SwioyLOz1Clcc9GVVYNcaoPbejBnbDmmNQVAf+8UPpXEPLc8rvmAcny/CB+mQlCjk
JBJWFWGNuCmAxxZAwWFJmogQUNFSUIRhL7ZWiZG1gQB89NSLVtCNUr9culA5NNUt8j5bxIJCEvRv
P2+MdHCviL40u3qo8sYXlZOIiXhytufxQpHCfoZfSaxW2BdTLfyI9/dKGXxiT3GjPvk2nq9c8lGu
FEqhaVDFotdhrm4+E6psUEIJ+Q2PCD/+50IQmXiU+wUq5z4kzf277NmaDxpB3zGSWUJUZEBAyECw
n+iMSXBvyaBwQpw7yZFkrTxLrKrf0AcorYFcpy9SDg1YOwbTPd/bf73Z3aINYralSSmbtXvgQdYe
/XapVsW1M4h5IkBiQxyXNF5x53wBvDBZU1SqOQRnFVefVHBWRI0dPQnv3rsrz53eN7HpactmZTRR
JZ+jFQE+WnEyaU4wz1F2FEWCB7xL5jaDb1FVKHer7t2O7nl5sRfY+IBmLz7F7apG/V7zKvpVRh0H
lUmVJJjEGLjRfr5JBh/wukZ4Nk4qmYqHJCEb6dmKBaiB4O3u5EcOdfukjFtrbePYXC7DWiz3s5tp
JmDpFKGJ3R5KiWuvK2uODWpLJ1JRxJ6ZENvHdEJy1mCv887SiGoWYBvRUdHxF7DzBFnapM+ddTcm
h1yf7NdLJ2rWQqqtp+PgWticMMqFA6PyZEbpTOBThNefM650csY6QVk/8debA1Hh6UVFasMw0y6G
U3z5pHCYcKy5qbsAv0tevtKB2i2OZvkew9UKESAX/jaSW304jGexrlXspaf89C6jB987Wm3mUxr5
7jSuZ4MVLKtyQFAl6OroiX8S4N/uo1M0P4U7aQfk5YSXWKORbnjHZPClEGQvziJ/HsPh0U2jRbJC
FiFXA6dY5FU4Kvi328SrvfEYoVU4OZu8/f7RabBDHPCn43vs5gJ+3ToAHbIJtkThOcFomcRm4K+Q
T4kz2tHj5g/Cj8OeYdFXTyfhc8EUZcCSAt2ZrFauoQg7Bv7qeOhA+YXyKe7sTo3NFD/muDJ6AROe
iHv1FvEsgt+Q3vGfdpMRRoa/PVx/1dpts42UPqKO3JquEbNAUBn4dTXevb9DE/uNFyh6KRP5fdt6
sLniErOGp13MVrl3YqoQ6YoSKUK9rKSgPGpV0l+fZhM0ATbUCDLJK5PkmjXZS7sSpVDhllsTqEQb
Z4CwF3GTapdUih7mXUW+IWX+7eSGcpg/Vnky98xqvSTYV4DIbGME59kA5mKMv6bk+eeryI8pwtpq
LuR8tD7og8hhBmZhrJd2gm46iD1JzAQ7kHQ5qc0RwEGVqtN5MAyY+XL9Ky+kBKICJQZb3E4nYcMb
X5fg0E5GEskp142DhlW8Ukg3mmB4WuRkfJhzlsi9cdYLGA5WIjALjCZyXzbKe6mrCeoj9r/n2Qit
D70jQ7Pz/Xp/r4PVwYadLItrTtQYfDNCjEjqv5vQSsn4y9Pe10m8A2UdM6EV/sPHGevcB8R8Qcmv
wftSXsuvhrXWEz/PKRBwl2i0jMSA6HFtMIdgYJBEp/05+ENd2RY1+cgUXFfbqQtg+pVj+ROYn92V
Hl2U+xd9t2gH7D46iJQXqgUePG26+E6i46abUty3CXy+zcOX3epILyjQTQbpGmoAv53aqAoZEu18
I9cSJRi1sJyk97Yw9j3djDM/ptjO5TtMB/dlRqXkessQbXh9Yd9WmalG+mkgkL6nGJDeFPN+r5Hg
joRWJI7sc1r21jcz8cUWX6zQmUoatNXkX+LHxsGjFx1AZqJAU3b47p45Trexhxhf8ZXEKej6sgR7
Ckqtd/v/Ket+FptMWJ5bzkBADyXczxY52UclGsFxdZSNX7YBamM8szjmUsUqgTFkPcOsVHukbvqy
bmyr66gQxC58VQnURTKjmpYeCxTqBBG8LgKNx8+814fCs+WZ/NUt/QYneVKZuW0/ST6hTfuc8lWQ
0SPq/5P7uRLcYU2TCsRH6ydEPVT0W01WklGSHWSlL69qOJ0inEcqgTwwJDFSTGkYx3Vrd/B2rkUC
w3/GzHmXTvBTk6+Tedc3hBjsn0LzchzgS6d2fam38dFCl19f2XFzgqKzEMo/dkpELLkqoofl2TEM
TYgLqhgUjUNQRi0K4CUCcfehm7n0bS4vriML7OnfsUJgOr01VoAEyuteyimIBL8ciuGA6Z76Bprw
arqrgIqqN6d/8gMuOs1f2llDRUTSBGgdtym8v63gkVQd6vmg8UIqZ5dvPginjEl7dNQNL7HvGVlP
hPw2a8DhFtZrMhSsN7L0re7DWjAkhAecckDlQRVVQuzqWRLVHBeTGhmrLCj3TZRXBnfqFmnSCeQD
eAXWvxtMx08oM7b8JY3ijNEvQrmHgoD0jxpZiAI6ISOg/zFVe7LzWauqOy5Rkd7Qx18aZjZ9scxu
S1m67k5APnTb4VMP5TXf3SOe9JpAh+pi+S45BbMdaKttRnfAtMIt9HGPgwh8fnOBa5FfmqSYFLsY
zH/KCL4G3veCMlpeon2lKPgrF/W6/qfky5gBaeYYoYuhBpRgIKjpwNDOigar9mu0O6vqDW1XGsNx
fog7jpa6UStwtAO/FTPRNUrnsL7RzZ64V6mu+K8Q9w/LuhrC9lY/tXOzdqbd45nywvnk1R8yfyFg
MgUFfOquVJ+7Ccge0kLUKQiSOSk/cv1zdOk6A4wi3BVJvDzCubAzyMI8JQ8n7jC1s9FSwMWzhqzI
d18FVf47+voHci6P/qYT5dl0ooBAePhwB+hN9TuqF+QIu1tQa/+uU6HR3XH/69lWdhdfGXRLBmcX
57TrVAXm12cbNN9I8emp18ZiVP6lLRa/6JeZMT17uyyr+j791t6UT83y0f5aE7UcXyQQsgmYhRcU
W1x5HkMD0B4DuSXA+tKvkHsnoWxzwUBbuu9Yx8sMifGa0PHqzPia2Rvuns+vdk6iOLunRU8XvWlQ
0q1wlyoOTlmKamhXBcufvJIhybQrcibdzBB4TuYEYuQPMIRm08ABv1i+fXG6RD1uO5OAeLz/bv7+
O5vfH74ePGXsprlkdK9JdhgdJRv9kcM+JfGbndTAvZHQG4+PH3kAu0nCmbT4CrcL8zWiz/4mpRP/
eu9V1CODnlpIAYlIlQympQI3/FDtQsg3Hyq5X35u40Z18qKeK0BSMnrk42C9pBNRQkS3i/XVjt5W
hsCHiHQDuF+cikEe5YvAyQnD1c2tLWqEEAyAywA8kjRT3d3BshKxlbSoC6czcflRL2f/Dtho+ugA
n0wN30BV0VfbDZvfYu1Ky9zdcqCTGY8RNXPR+Lvml3PkKrZc8HeGNoXcGklPUJRV0Vmnfn/kzXtm
xXOXZqMzP6pgmut3ClFtIddNweRHLkJHnM5HqFFJJ3Qzdq52n1oqqFAALJ1rtgbgjgIcludyfFNf
uIH/rXuHwULmzv173n1a79fQTNebjgKnTZ3V6mwhUV8vyxjSU8TviCSU2ITITHiXcVGXxjnD1yAK
3EgMvijxWAtRiet5AFYRjTUZrt0uRSFdlrpiL9s46K3W0JSexfiHLtHygYyXBR4MG+dhGB7xfws/
E2Erj4LtvWGtfVA2buzl2eiyxOdvVXcQa2yZA6Npg/H3d0NiDWn4i1+hIBx5hKZV3MGlH9gd08wZ
QEqxALma3WAskRCqqQQ/eadU1Es2Sk0moTnMFrOiZOS13CLBxmaN3eevLyLZvecwSbXsbZXzQFRl
tZmIvUtR8zYFtZ80PKWEIASEBXa+aqFXln5l8jv4pRjP9Gdj9IScSAeSc/TagMIMtIbmxH+UDIx+
7ZPKcR6nELbNFXza1S8Pl8cNNNqeClbDknsPEoygBdaJhxIx1xtn9XqmMCq+LCVcG+zlBFUjvj1a
DIGD/vqahr6xMwVJNc0vmK8RxmGkg97ec3q8QDwh7Lc1HimCuh8gbANyZPa1QRgbkRSvvXhN/UXv
I/SxVzmLdlfDS2c+mapbss05fBgPaRlRfmm/pkM4yI43nX6G/qCFp+RFTRt9beeY+t+/4IFNaV+3
8uE2TmKBJJdnrkEj9UJ0sBdTua4k+JCJJDK3LB3CbLRFwW4ZaVLm8PdtynmfGkt1180ToU9ZdXL+
PmO+ZMXRhz4QqUetEgTXiNBAnR3WXj7Rb6DEdqUo/K3L1pbKUXYYU1ik6g9cvDCtO+xUVUVd8NtF
Welfuid087xGCs7g8IOH7eJkP69yCUZsaUESQFSGO79PjRnuFhlXcuXZpXazwXDq93WVAT/sp88U
J2hxlU74R4FFSTVP+FuiDQ+R23uulCa6T5ffE5EIY+2AGboOG1w7AqcxbSWbxhgp5tMZjKGtp6v3
wIhfZi0bRJAvfdsC2lvts1ENxvf3mGvc3e5w1MCnya8dJ82/bXJ4aaH/C4H/JZlopBHtGbQWtyxw
5jxgBt/MBfbsGYIwykJG3CRu0L5W0i7K+gVnxjsuVMjhK+EbBrT5eobNf5OHk8lTW4Z3ytMkIUnU
sChOHKErsGoqaJRo1yoeRvjUxIc0Kns7tBHxrfawjR6+yaxX2Q8fBgWYiJd0IQoW83V4U67fmaLv
1liYdl0WLDphNECSXJLRTnD5BJf4FKX5d7OM0dDa/A7FHN6XcJiANBOT4zY4IgAqnfZDBa1TnWuH
7NAN8dRUP9St9EXwFwN1baJzkVWcyy4oP67bu08r/zJIe2kSG3e2CpRi0HxWgFKCBafIP8qjRnka
n/NJRax45p8+YIlojxUWRGtqXuxrrIzSeihmctexdezRRsQHVFHuGPufMkPk93EQKilytzYLh8ul
kYlxSSf8WHAr43LupFl99EW3ubPvJnAZSCsze+nvvaZZM38O5PrsnkcBFkP3FdlonHMoZjNHO269
ODD50nIP+twAsfE1d6Gh/f2duMkThD1Kf5dHyS+W8056yVQx4Nbn6IE2PtiUw78M7/R4jZMkbw5J
zXRzKLJ71Uo/HRT060pgWPO4B3vkO9RzUzEmtwYbddu+WI1ribVGnc+YrXJ0byzdQKxW7OAczTCH
qR16Ge+NjMnrjt41qxWZt2HgOWeU2JEUa+DypRdXgAJBgNJJbGM6dpTK/MOaAO9XeMgTzGmC6dFN
mWysBmn7fdlMBIEMSuDnjZHNio+9Rk+nEh8jcKkWzve6AwyAMt4pvwNsaVAou7p2xTu4C5ukPBMV
sR5ruzISExWyAbhvO2PXcSTr3BIAhGti7929Y+zaXxW41Dlv2/P+L9RprRT3ohi7TXda+YkSTTs6
cOi1Ov+QF2nV1kBBRQDAKM+JpbLeR4qC++wZU/ULKvI3mOajE8xjypZWw8JXZaDKDV0t/+9e1Wyk
Ji5dvys+eZI6SUNYEhkQzcodA1rlW+kdvVd8I0Wra1QJi+kFXXpWxS7QuOHLFiktLsJo/Wp11YOm
c7vjwaKqOgTluWXPH6L0Y2ISLVl0vxX7U+SiywAmdEoVCy/sWAyaSyva2JPjzmA4Gqq/TgELZhCo
Qe4is6WAyg1qglaJGLf2Dec/VVNvhrm3Bv7909iIBv8IsgpaEbINZwvckkxvjmxsmn4f1KZKzune
3eOqHgQ5+SfdqM7w8dSbIn1DFgsQqdZ5NbKCfA7xIzXzUoGCtf9QarS+946Q+LHFRGahoEjAmHIz
MYmtTxKcrXyL8jQBUxFl6KcRatZTQBozrQ3SwQnarIa29AQ2oHn4k6xeddcqTnIwmqzPMqr3QlTF
lFTwEYyI1n5iNEaNkoHVD3kak9mK7l2JqLbow4/MFsmnL2YUD4jwZuLVBhdykwzQ98y77IN870W3
l2dRIL05OP40F5bBURuLY6OiKw8qVSmvJmtTlBFnhUwpkU9smpxcZzbrMeCw2fabYGGg0HrJBNog
FZVZNQgwFIGjaFJUh5AoBOHLmtXuFFiw8XwW4KdNopfO0M867z6fy3baPqQ4ztMmxCKWUhiTUgjA
s58n9dN10pCIJE1ROGsGfEuLgwd8MF1DrK9/wCpthcom5V2aTzSMxmHKu2/8Cfiy7+aBI00yPGPw
h7/DTTWuruemDu57CRNRnrs/5N2Xaz9pxMOomCEr/rvlYPO/4Dvg3J4+jlcK0yHBxE9g3xMMvTo8
RJeyUdoAVvYp/T8sBaiiXuJNYmsFyAiGsxyRJ+lqLzm1r1UyMsJjzi8xNpbsdIPU8mnp1EXIpfqR
qvBWdHkEn2Sq0LXvgJ+wMUIUG7200GZnBRWQQ8iaLJzcvuFpCN2sP8iXL8oqYAEzfzq7Njtf71cm
0iondbfREZSOzi8/D6pd3DWv7e0PAec2X7s/eUlLVT17+yJLdd87r8/viDLxoGwvqLChsh0a/a4w
WFp7ihS+IvvoTA5veJheEvbfWhqbw0axRCRpXG1NlqPhaT90EGNB97oKMd/4XnOz3Y0xJQ5LMO3b
Ttlo1RAYBDaSGYTntPYxHNgMmunIbKAcwwhACqjm+uAac481Kr1gduUW1FZxmreolsVju5h2TFy3
yDxKKXiQREJ3ifAaga94iBZF7h7K0uZsLRqMbTEwiaW+bT1QPpBme8+DDyPBpRbtrjPO+6e1Dfin
ROgcFibiPRxqjM+ALJJz8dU6E/qdPAOQ6JzSSvUvbVVS+2iGpfbbjxdbisgRRxZYaQjUDCBgK368
ZjNLf7nfOTNRgzT32elLTKmT/0+ByajEiQ2SWz3KI3xM3NGhBs+x3yAzpW0aHqCNFQTL6ojua+8H
BL/dGSAmZt6DWG7pYKKHChpGQmA+LbfUi/BTmsUEkvgAybZ1lNEjo/eDICYPSB/aGB65e99fRpyL
Tl/4o2LpUk5M7xVREc4O669yd6jsUviYfqxMmSATGKXNYdJTugzJoeRNmaVszoeowMQiBS9ACMP/
jEXe74GxC8N5BbqEN4hbPGAiNtE4dzQx/zNUOVbeCp3SQsbQh0zp7dPkHNnlYMmiizvcHLW8OUml
g/GX3OvDHY1YPtWfAFO4n9JocWc2l3cyp+p4MdX4lX91xMnO/tKDw/mfhLJIjkvgoOU9E+7rF4tp
/QKAGvsieFUsw9ocLYsGnr+/7R45bMAMpSj4ADidClIrNGlaFQq/fT7rmzb8VI6FU0+4Lg/KS016
uosI6jAzz8hu7oM+PwdQj/LdIYOXllfqnXgzmCzGOcAKGIp0eSlJTqCE1UasWn2XrZJCGre6FHu8
EWSXOu7pESo5UqWVCAFhvFVI5a/cuV2bYaSHN7tTK4/RPMcdMvrU5WSmm2kvFndU5Tv8U53djoTZ
XYctVeUZ3GafLQW4uXr5DR4wNjeQbRjNBAcF5wfkrVz6CNjT5+L9pWx25hQF4jOkgeXYOVuXbrcS
X1A/UOieh5mJ4sSbeZ9qRuUz0uEriJOTgqwe2Gh9GOV9cXa5/G22tf+tDbFfCSmXdAI4XZ15U4bu
vT9PzceV1REAuw95PUan38EOCIkBqCV2igmRx5peNz++L1M3XCY54DE9q84HvnRDuHJK1zcWqCNf
h5RZxB/qOPxD41lSOzk1795BGkvQ6tx1l/BZHCZXn0Kb6CGw+behaZo9HpacRw3UMucFBxY/CN/g
4kKllGCkslsX9NVu92Hpcd7taoV4JUNemm1EiFiXhtFZOXEI/yfTs4bIi/I7yCPjlH5+H2yaYxTV
/IkUnwacswBtkHfxruhpA60PYKIxL0G1Irl4CdMBdY1F98+Wtb87Bt6DGxFXKwe3KepwWBS/m2Ea
VhghHkeOglskQGVj6nu+fTVnWhOLwCxvlgF+NQveLKnSUH3gs+bT2s01AG5xvli0NiFMjkqL+rN3
px1WAKJkcJosKJf2YrsHDuFQw93Dl9znCxfhkgN4yZqqw70kkhKI043V0dSibPQACfVWkllRNVV6
8PaEK5BJ5XiXsvogG4DhOIXirYyAQ2ik1jFz15n4cZxibT2iy6z+EZuEBg4UTfdpNF1ur0EfcS7M
8Yuuukx0JlrtBAnu+hMsENXRYgnHNEElK5zpim3Jbh8WC1H8wRwNBy9qDB/SZEk8z2iukgnoPOC6
uf7cl/TbNamv8ylGVJPfAP6Pj/wyj/KVTtMBbul513f6M06xGyz8eOF4cr5gH2QYlBAj/lfJNTKt
zmge9TFxAMMDZje8nldKO62vmdi2FzKSmNb7pxypAQi0HE9gO7IC+zoGGQMMJDG84ANfmF+j/gm6
X5hFDew3GsCd0bRqgxms6fLoO40ffxDKLZ9KHRFQeQrBUiH3ZmZq1SXGQelv2o2DaWSwBnd0TMin
2mjv4wMPGoqlRVzc5kK1R7UM4tZDHiAE38gtS3Svb2j7ROW+vAPtJ/q7MTG7stlNxF0nZ9fB0ty/
fYpy89Y+7Q6/ZMUiObMGjvEcUTm4FGdPCtDvbfEBBRAltT+cSUa9KtKyBULKXM/J9lOuXX5NI/8i
qHOuGXe7P5T0wgNibZToPIlxLMwcFVx8AyHruSK37dhcBzw1CN86ycS4REaXg2Qg8hQ6t3HODA64
QEZwUBdnUnNnC39PKrDRISiSfVRGR8iDBtNLOpSfJiDWMCWXkI7aBekGULKKPs29FC3Owf7ykqg9
Qmgo7+QoGf9W2TH+cRu0EyZKCiVbd71ZNiEEWodWGCxAa+DCNRBUu2hfhQwUxZjdvbw0EYH3k7Gd
jB4HvNPL+AxZVK3QNbsqkTbQwRerGH4qZGwPv+/M06qki51i7CYl3WQFM+7FojN3bSp/b+cFhhxY
AkAjMbw2Fp8evlU3LsiWdcgfXwbXmKwmwttBUTa7IgjYhvSW9h1P8ztV9lvDL5vIimvJCgH7i+OJ
sE4qIKhQ9+6QRs36LUc/9qmIpv9VjuWEtVsN2dERJe+UwAlyMQt8AP+pD96uX0EyT2vDwvjlJEr+
QK/pWqBBZzVT7P4OrmGtx9DLTFm4j1as0jiPzIt3m//8VKkr70KHcNf4pbFjk8W7jBB66CR7EZAd
jh+lRqhxzNJfqFrydqwdgWFmi7iQF6EVU9DsWNkDmvDgdydTZNCvxReD7/NB+bHgl63MQp8DhImX
/DnPcpttSMyQy6mxX1alBFAwiSTwY2clHmCkvWZ/dVHcQAER+HiDeyX5lXRSm7lgKaKLbeciwhmS
k9BGkO7nJgjfP669iVFmCWTUAMxTTNDmaDKhG9ztvYFRc8Kuu3fHodZUsg/bDxcgv8+sTqcqrSXD
qb/Cf7xVrwlHB/qiWrboCZanxEPqNhgiGV63skxZUX3qrgjOdIWyTPAleiH3edj/rTU+R+DQ1FC/
Ko0S6Z9O6T+OSTRW5eMJcxI2S6keg/bxKpHeeMLcW9uZxQ5k/Zdi0U0hAFBlfMK9tRBHty54uiaa
R1mlJFSv7BE5UhcJ1VFeFItkg4Zpy+cWR2SMTV7YXpUE1a1QQP75WqbrBz269CLpqGwVKAEsO6ES
ZchMtnLEBO49CHstGsvgWjx44dRXi0kkuiQv9SGyM2EXFbXYg/zZ7Z9EPgoI5Al+N53AhauOJbf4
OmQrcIEjCjT+o8bW8q4R7dF8idSTKLJImhPRHJsJvMkYoWTu+1/6YkuKLRliCEEJaQG1Bt5zrnyq
pb1gURz/SnEJPCcnBygYnQuIEph0fUnnkjcSst7711/HUGJmc4amS5nkw7dgIkuX9hv62O+F+H+m
xtfSQf2HxsCKboVk/ghNcoLUPhaSbsQZSe2Gnmqu/2E9NdrDp5FPoG9yrHMWX6x/Bxam1fDI0yJb
cqm81+X7BQbwl9HULUuucIImy2Xmmx9Y0kN6gEGbPZwIU1+2rM9CNcC1LwUo/vXB0uY6dcU/93EL
mzGBUpazrxnsWAKlGIYOLHWHzLLl51H/8ASikNVhOcL8i4dKu29lazTnVYx2Gjmln/huaXy7hr02
SogP3/MIdDgqfLLWQxn41QfVBAjCGXqO70ywFgIepF/cYZBweM3QZsEKRJ9V9JgJIhV8/p70XnZS
IFZJaC2jp0W2A6ucnAofbmas9jMY4tj02dUJIR+9QzEgesRFnbH3LdJOg7/XNXWi1y3e3f2f0x/Y
WQ0bioFmBmq/TUWlG6LFmaHr9mxmx/ngDxskbXDyszLLDEH87kNmU7xcTBksii41zZEvVZsUQnAl
LzaDxiF+hRBI0OigQaitiI6NG8MvxAUGpoMH4VB3HorqGgMEvnu6Vs1AQH+sT/IiCjBv+vuRBF5n
uBOUYZanWX1bgud4+bHt5zsl8Y4o2J61gdorMDLlLsr3Cwm99FJ+mq41oLOa4R0dkQCVJ++59ZHe
3v04VkUdDPInQ59ulK8A939hhC7UDHE940ZU6PELs0+AF4zEW5GHsW4Szhw0oOrFdYxQah3D0aDa
L5KjkmksqzmIQ/xvE9YXJYFsngDmrCASq+f9U6bhW6u5fdy6JSexiRKwpSaONxzNEmPZ2WA+fsCR
V1Ye68RElu/NHTtbokNatSLjiqeNM8QSKp6RDspZfOEVvoauZU5lL8Qzum1CWesPzJfx20fWo5oM
IP/cJgRFkF9Hh95AyQ8wwh01bqaSxgr4G5d+xzGScKiJCHMbpDV+EWNvX2IVsc6zdQtpe5qMJybg
aNrvQrO0AutGyE6bUyO7Q8xVqbo/2i6fpnRxh7tFeoACwXCoFOKqx5O3v8xiO/XMc6EH0kDTaWB1
u6hPKGezOK8LzCKjkngxzuvxsbBTZ3TsXHOAgukkBmgJT1RQYmwcevjR3HAn60UBc4nYEMHrYRxE
oyzkQcdK1akipjTsr9XGrr+8HLhZoLMnvV3aTU06wTfIHNbHxTgH1OTx+rWx+OOGMrxYwoFEdYI2
8ZnINpBeWkE0MdFVqNXC75ltuR/BSE2QNLUezlItCrbpa5cvEwvAd8FzoPaa6uWVIIzPGw9bMnUa
cR+n7APvpLcizro715aNcj+RLAwAMhn0voo2TtF7XltyhJ1/v4V+Q7VbwcHIBwDv1aexeYD9jFi5
iCJOFwT3xPrt1NhBBpJvDceI93Ac3VaHbQfEaRn+FOOwU33mPHxTvQQnweoZsCBYk0msw/mfBRhj
mYHs+dcJ+wKuKnl8o4UY5FD0Yp2HtMso5wiwY3AKP/N0wkZh4C1NVQnALnnJT4l1zPWsfu8AZaQa
KDcWlZbBsBfzuFPBQQPSD9yuNlSYKcdluR6xpZr3qGPseN2Af8kqFfCP4yjZgyfAzJQPxDIug8Mz
KzBLSqjqZKYRC6zMgxKXzqhV6bQIGfcbwjQHFtgboiWiancUrBFTjWkV6NsSVw/F7IW9du4UdxD7
ZmntnG0xHeSOlFaPM/SEbZo0oTEhxQme2hIQRf0pQbdKqj6MemtURa+w98OqIn0ggupEgMe/13MY
Y0QMthKEbnMvVr5PEQUVCrlPd/vHNf71KAatezT5BqHgzhw8LL3DsP60J68Rs2UNWbuzWVIdkLEg
uTXV0cOn6941zkxRr3KI0VbXf6C0+OC95bauMuDD52SY7ffDeLfuCw6B+helS7nSxDR944RZhtW5
3tsuY6O6HqTXGpl27/KoRsXEyqiWKW4jix/FJ8A9D0f9Gm4QR+UFST4M2dzbk+7O7LIWeigGtkKO
M1eI98xBvy9VmNuf4p8vVs2mjMSg7OI3iSmMpDAh8awOuY+JOgirnQIgBoAoMMV7p4YhtYijzmn5
lbWuywUGUZzILN5p6qPhHeFVwLsVMUcxHpr7okP+IySzLKJlTZf0yQaAHDKT91Hx+m86V8550MHd
IIYq3qYKtTaKA0fxtSlCUeUCgpl3/iyFBGuF4dI0yCLmZXWbnb5avf4XnRcfBa5fGtSBFhxOK8a+
CUMJa1ehPZkFw0Nk922UVSTTZQ56Wn0cUrEVGmpVHvm6QaN9bjOSeT/hy8u+XmquRM3R0mjqKSnU
WjONMbR95T1zmlk602JrJoQSG9q9K+XF8Q5poLP1M2TseIjAFFKMmVsz6tgGHeRkvc3+NQFArQ74
PKAVUMJKWiz/iOiryTqQUnw5fS40nagO9Ukf4s89zmAITNyIuGbRXExpPvlJhNURT/QjJ6co+uwZ
98n6znFeK9BNBlPxceRJ3p4Y40gqWQ1ZGlaAStGYn7Eqdlz9SKEa40Qi9h4QTE1D/HvCFI6NgMpX
bUBlPKugl7KTeFgTbq46VX3D2TV00cKVhFT5bvGJGb++kmQupR2effnaI/GqQq05GOwWW4CFWaVP
Iind8cOARIe6ZkuUgXW95zufkOjgdK14LB/vnxQ9DmZFObonfxXgJKS5BEpAZnTEHJSFhruzFayt
xZunf7hdtGxnUOufDdmGnv3EQhNwC2/Zx0mW4+Q8LmzDuND/cXiy5LEoYGNVEG+KzMhUrbllI7ua
nEaQmLuNTQ7PKRNyVwKivqaM2q4eF5l+ErccqLRZ/54TBGbU5ilcy8Abs7UTihdF9sMb5XXTlUUz
wflWY0xdADtfuKu0ltHSstMyhuQFtVDOFSdUTPCabdij7eVcwj36ZKP3rihDqNdPxpWHvUJNfqUF
EUos7b4gWSM/Ma2SIwKbIrdcQ09Hy86vsGQ+LxyfBskr2T/QV1SxfCU3QuizcA6jdjQk4C3oeH8p
NWnCIzJWRFNCfne7vJW+Sk1/14tqaX7ne89SEUY7aCvgD8kXqXH2+9C01pFJGPeNFYRqZixNYweo
x21CsWKmfi8PSVgHDjScB5gn4zotdcX0qNPlZu2WKwac4/xJUuP/2T3azh0Fyuy5rpyU9qMhy2Nt
McGfaTytKkmFCDd6DzBKregTt1qQIndleNxX5AA90Zab/IhKfg+p/Wlzu7mIvaXukJjfIWUvLcFY
gTePtZ3PSCgC3wXL1dySPZCrGYKDLMNOwX3GejgPwXNoNulxERcsqwzyjBLeZmaoj23cRuUDc8zb
NH3Zb+ONAFb41n5It1N7mqmv8XRlOzyfhDvbBg3Ac7P8lOqnpGZgcBY45QLYTbihgbXow1/X8sc/
bfQETwcSIq9JkQJE2aVlK7JWq3+004KzzhrRtEw/0V7LRkoW/1Y06IVfOZCfvH7VRoC6v9KlETBp
pwfS6sABsawbJzj6lULVJ5y7xExEL7h+pPTu1A1cePsQ2W9STih3eM/RZiL3HlSZ1KbsPEpp0a+/
Hpi7qAmgcG4D6ZqetG3kw9GniPWBGr8PaHNCy5uZp4hTLSWQ2RPymd1U7h+RPJoFwCT1rXH7UAgx
AzYGNObMie0nLf5+q1+U5Ra1jgcpyNbjINneShh2RRkxkn2DCHC/+m7KH5k7jAr86LeJcQiEtuZn
YcVYtPCpawIsjNqZ+iMIlohs3huhC0/LkeCL3B56l+Mim2gh3jsIims+Cj3Y6ovUrLSbO9AXj7UM
51sROUSqDNE+avemMfUxV1r8aeBP73adetMb0xq/n4inTwosR3lHVo0jNHnofFQQdy60WZFQiMK8
2QtTOTQkXB2s01snMRZnw/8+S01jsIQ+BsF3MeRcTF7lrxkCrES+3t9SrdD7wpoxtQLIOnznnIOX
0UaJmmlvrSw08lkbbyfPRhGR3Si24YKlX7mKK81RSxsolqP4+RKYigf/SY25VP7TaXptonVFTCta
87CnMA0Fnx+wGvvONfThgKMgU5pJXJGmSnIGfscW3dNhnJ6gVedBuslScG7P5hrrguNkqnBbpWXp
/ppvQGsjNrYSuzNTixMvJPJnjGI5DCCdXzBjIOA8Gn9P38yzt69YdgU6f3VucDewN66baOwuuGVy
6nth3lmPrDyNGWMDT+1fT9H4Bq06obSfIVS+ES6ttFGlqo1y41mcMJHFY3YXZbo0igGz4C3CobeU
nPajLC9481i3K7dF2r+AhmNCiuurDZ8jdLmVfMQYnfgM15VPxa/ZSsQ2L03Ku3nfHsKtDAJOmtA8
139zbYU7v7xNm8PHRHihFdeMxbl9t6WjzEjPcsTzXkMPV2Dtc0XR9srV9k7CLbuIkMJAFNUYDPRA
6IRUsAwfoK97ERkSaZXfzROFcoFDUvUoS4x+vUVejfok5Pzl6Bvnubf2yEfe4rXRbpzvfqBGsbSZ
mtuXoFedMxxXvDt0D35dErC/QYKyiDvlzO6WfDN+KLSm6HbiNi2v2B43D4K+4zsK9gS57P1du0bx
nODZ/b4edPL5xai8ZADt8YAY5ZPklU0740hgGp5MJB+Kv76tEpz2xl1fI6wM21fEcrYSrUIjZnw7
uQWNDloVPweHivOFZSIKYaeE2g17mISH9/wrroRO72oqpPr09KCnIxX5c9tc0kIAmnFtxuCjeDQR
9f3aRsONtaq6sycpsI6YHO0M/pn89Ol+JMI7DggywKfFWuHy4QFsYTTvJGWTYbUxvdMnA3lTHbk3
pcPfnCXyxijJEEe41UFkiX4ZBaPkJQzTPQBt/2GTOIazv6OjY/JOc+kYytBAlL99FP6zqkkf68Dj
EU6u1i8CJEjeqNA0UpXt1D9eYFCMlRPG+SUTbyVHjf5EHsAqP6ZAmJrE6VIdnp+w0EUyn8vARiII
xA8EyNczxLizitElKonNwQFkpvVzatjW58/btH+wkbnMmlGl5Y+REflrjUGiqUbUQSwykPXEt+jk
i6kUXcrBC7KU2m6K2wp4trX5ju+ieeiXjBG+riIKpNswXQBSKpCRJNuGnFU2/F/uGFeitOH+TnaH
IxBrsMGwU03W3KzbH/6KyQMU+X/Y86hJfsTO6w0Az8bPrZfARuduA0e/gHs62EGhT6ATB1W6NFBD
p7AM3UaKjX9frauuCWgvtxDUr0/WwJAccntOZr+C6gQFD5K2edWtusE9w0ubIYD8GBdNB6nV2Zn2
4Yeil0eLkTH10xS+3g2hSMcIITVocprvnUFzcYy3acvhwolFGO32uHCfUXTQUOtLUZ7KVRPaQiGC
glOps1vtQ9ELedRFLPJcS9aRQpvFLgSzDjb1qFLeqzmxer6I+gjKZlaQGDla0PzS8jD64ETcMYFa
14Vjp19rdY1DzQT1Y0G5Rbij7B4XHh9IPhPTp1evRLWKXSFAH4kZ8MvSF5oQ8sZUGghpWZoMH1hR
jjdBglKHyay6XbeB9kZs78cvOUjpYQJt37Y6l4CkPpdLF54RdDQJTaMB0nhVOhhRAa/i11c2XU30
s/eTxTQAVKbigQV6BocEGkJesVREHf+3Zs0RjwfZ835ZnZcJckLTF6ZrKShLF+biaAvOiqIdAShS
f/egdG8k3yYOeAMxt4PPv9VnsQoEmMhMs59XiERan6aRmIdZie7XuuY3r9ComHkdkgXC6S5eh2kc
3XxJNzeIdY70CNtbBe1xxe2MnNZ39w0NQQL4ISxxck76HgSeoE+2U/cjQ7QViZXZL6wQdNr4AuDl
akIuf6BUKDwuAXQKsxhc14xmqJAo0j+/zyGDWmnDDE/siMjBSpTEsSfaSnAVlNScuLISTrADlqQQ
9EPOVgiHFyMvXVtLW+8QNcgjVWio3irO0sCkDiA9ezP+nMHWLuUmOc+C46h7ZJeko72pQqDQSW0R
ASLLZk9if0YGf9bzbovan/RDJMnKmek8N6D8HE7pVzfj9bJmY9NkbK5DsG4ohAb3jaZCS7gqqWP8
sH0hSvIjXp306VrF56jLB3nAJDI+MOG7garzxAtXTbJeSgXIcsyApy8ir+VYojK8Eowqnys19tqX
sOBbPYcqLRvsL/cMDMk4PtJ5Yffunv6SEBJG4cEPIIXIf37RzKZm78I0SwoiLfEfU7UrA5U83QRY
RpFMfy5zkwKho1gTVSk5qbBRaFIUAJWcNBGICIR+EhVT3h+vxaTVzggK/fAoTD0P0rgwn/hJO86w
TJF8iGuq6jRPMm3H5s0hlK5TlQaGkxq2+i2XQHM0PP7ZfCKA2PbtPaaTMj9sCvNiLzXRLy+N9nKA
0X2a3IURfK8FVPfpsvos/tr5q9cdIkzUc4cRw2ePPl3OlePJv46APc7MiIWP+7a7uI/uwxVSk1K6
g6csl14aFefIUENZWTa5HL0Hhi+lyjhCJuJlZsdP2bkfEBXai1INX3eOGorqiTBxAQZ2gGc2TkR/
G383gQKpXD5tVzggk3UrDHUafffMZmIGbK6dVWIq7rGBL3PcnBmo0Ims8kzK3SWsbs8HWHbZvBNJ
Xik4hoMz4JlryaLoALDr4gj0Rn8r7mKaDbJTwC36WdrTS9NWaMUP0vd9g32yHKwoqlixMbx+Iqkv
iaxIdsRzxfCvT4RvkPoSi4owIWde9mhmjZHSFtZI7Exi1jpyGmA/ZuxyTO3sBI11/DgbJx0Xfwfz
Dmqzp7DMaRX4fwVOMex3pgOr+h1jHhYh2WHAgBnO5m2JFJte6NSajpAE+hqycVj8f0QzLHLv9s73
zFkZysDL0k+oyrgGk1NKMB8x5gBo6RDD+/gG40BPDZp3Q9ZqY/DEAYyttmC+ZUl+VEhD/ayKN9Cn
DvBXbABZOSxejBuoLUmNtMNE/sNsJtQMmUoVdh9/6PZgobFBDzgnOg/sEn3SlqoEN8vevQRkW8zC
+Zb4mdwfOB1ZVfNqY0oRvIAtCapV3y0I1XNy4HGbmPot9ynqoCMiCM4H1ghToFBwTC5bMsCidZyA
s28v3fklBxiYxyAGzP8gEOSeqXJ8kdKFMHN0kGP/eB4HNQZUJYLfsKEkWmgTMNeOPSGtz1jCk7no
7/IXlM+OiiY+3WoIR9WUtktg8KUyFQ9xEjBK4YloTMjFwXBPMao5+oMyE/iLNW4tCRvdVaasCD3z
EtF4I1K/PRjMqDesPwaQ62hYfOM5vf7bv3kuIEodk4TuQKdRXyoridBkAgbt6GRxklB3nrU1KXpA
oBlg7t9/cBPlD4qvU+zt3OmPTlqv+FnF1rCNhoNeTbioiLRy6zHMaSTSnQB3Q7832TutBn/RjWpS
ivXeidTgsybUrbF2Qwi9VjzxjFU3vDFxkP1MTUpL8yhumw7kno7nvrKqICGk/ovQ6jWnfQkEERZ/
sA1lrXaJKrFPhNteghuWA5cKZtbEva9+2JiRJBgBE2LuZtcJm/okqw/8ZBm/zmZJ9KzUhICEh9Fn
HmSxHoMcSIbBS38aoYIc59lF6OyVI6oaPncjN6PbvQLGMI52z3O5cojUugNj1k+M3bABYMZLxb/y
UwEaVqjRdtFAuiEbhVBK6xXmWrgX42R0EhMeAzT0Ed56CRd0yNe2y+lU0o/XGHLe3oKjRypNfVR9
KxQFposxf6meqiN191qZNZZNDGi4g+q3FAi6RWDj7bbPZwkvtP4Gcu7sjTMVTUXCf7pb9rYhib/3
sZuyHWEO4c4cEOnv7pJq1RMn5rcMJF6uI7RDaRVCrSFfa45O+ipBbf6Iy0YG9lfJ5WD0/XIhk86R
89/KxZ1Dg1qAwAZREEe51kAHpP82+NJKvCtqbYkf0JznN0eJj4db8dexDEjGRlLInhI1QFNFnofc
4wpFnqkEOpgSs4XABYltqA9r0wjN7msshHvqWKLnlQCI7q0YhYSooOy4EyeAOpOesJ46pHEZgEDg
8e9+rEdkPeJtxrrylO/7+fYR4CIilfwuniMQN90gkMrHBfdyxFEZbvP1UfpfUk8RISvUr2Ymzkdd
4xl0nH2nDbOuAm8v0YWV2jHMoinr7R/8tmVVkwaYeAQM+ju4DeMCERwJmi6QcTevl5ETEgYIUspW
BzWO5HJURZJEvtc/JBEkLdcepeDQyspxxEYi+NJwmXzlvX9fofRs5N+emzscnBa/dAPSdGYH897s
qBUUU79Yansq7kPVZZiyleo6mXuAR/pdkb3VX0Gjpi8nIAufRFLhzptE9HLbVeE+wpZkE2UsIelW
CWS+s2SAtk4Zq9tFC9iAvZfw1QCauhaCeonQ+E6rGeGWL+UxbSuvyHjRBj/MHd0eabaULRWLXRUN
47DfdWHNCAH0AATl9TMN1AxHTBVBWaFqCcncDXxiXBfE+1ZIJruV4QQFX+0qJTYO8Dk0x5b5Ruvn
EHEXQJzardWFq0idrh07ZrgKqLjPZlFkGF1m3tAysFN/IdWtEVItbmBkpGU9J710vp4TNKxSqy/w
T2dtzM/TiqGyVWjJKaU4KRomskpFD95J5QqeaM3eewmy/pYkPmdUXLANNdYfkbNzbQqBNaRmGqO6
fs/ah6GWDELWVfChn1OUqymPKfdH4jE48JJox9rnM6mPzMzFjmrIQlUGnPk4s09/eLLVg+RY7153
KzkuneyvH/MreU+eY0yGX8IZPw7m4Y4z1xI21dYpD8vCYLwndpgUF+/Rxt+MZb7yRoWU74C4urqe
SofnebaNzo2MtSOHjfmc9k29W3N7emVqYeBYqjbwQPfAe8OXRAup0n0NPVHHJ0tBsKvG97V5nvYL
zDRw2OMwcMk7Q5nPlwfah8DJx99nBg+ysFzbxxWjbstEqK0gjSdKCggzL+IKRXp6ILTGdGdBZr60
4ToapRuWK6xjY98zgd2dkjRKpJ7GyO66hrOsu/eShcEx0jqJ+S3dy74lEnHpzw/KQDDhBFFOkbK+
7tapSajWnA5FuOuKMyAvm/sPZJXH+6+KW+ZlPTcTMNKU0bvS+eNJm5qisKWBP4vE8WivtSDhKQh5
ury3a6LQQXZ1MxfiQT3bH0BdoVDj8Vgx9rBkOHnbyvB0HFyHtum/h+sjqRphb+pJcZ0LlvcHov5A
9Hwbfaj+Bk9e3i0myZUalB62qMT78xfjYg6NPZB+HSwSZMXnUjdCFIKSh2AYpXAeHM/Xnn92U+65
w+qMLXlv5jWLMoEQpkHAzxNq3ndhjhatG71RFk5lAgUXonwNP8tcOIDlzyRK0EFxpTEooNUiIvAp
yhRfw8+gHvKSNl6KVbHXotdypBkxjHGa2jtyg1c4kzxM7EVR3aY+K01V9i1S06IWmn33hA8qm50P
eph9G5pjeBj/04uVUao0D8MeLquq9y1bvv4hNWTr6NAFqJxDeQC/WR/PePjMSDPzCUNHVI8qJyp5
hcs5i89Q+nVrIMwYzZooBamLzIbqIcz3YT76BJYrJpDTfImQrlsCFrACGFSp05A6NZCfUgDEPNR2
TwoUzBrnm4wdmR5HwUUtKnqyvMOxPMMDeH61wQBtmsEeERBaArIiLeXfL62xV96zMtfNTA9yT8im
hNyPDM/9Qw3wGPMWG866yJeRq09CuC1nFgemch8GH4d66wKWvKvm87+TC8wEk1uS8YsJwwHWK1xl
+ZI+o1XIp5go7xG238w/ubxiYZb6ygbiN+5Zh36QEzP72vx0c8L71SAxDUywlk/lU5SwKJEl3UmC
HjAmzX4ndwDeFPhwIyXssvYWxm7FqdZKfetJTsCBtgSTIDU66ypDouLiZVV3bt6EvZFBRAQ+MI3f
S1ztxPOtECPUy0WLSaW8TZiqvTKQgMCU6iBWaUJwK7r+3PJZTz7H1K3FfwlWe/+vzlKz2j/ar/Iq
yj+37RJt7H81NEtBbfefn7B0guG8TH1R8wK4vLDe9+LbIrm9fhU8NuyDIAFcGzGb+ioEaklnlQUs
jClvbBJCd6L1keCsv1mqaAjuI4Na5rlPWiia9yETG35GqKWDgnX6N1BTLxORAeQVeSb2gVqCJMN6
iWKr9vAC6VAUqpmcFNymV22isTLFv0NKHLX8vEcbhrU191TSRCxZQOmQnZlUBI1VmHmqQZ9IfD4S
QwYgeDnlFCD4a9mbbPUXigHV0D6kQpFa5VVWnsze6RzAE3jGEPifD1ztLDw6EudFTxzrHH90w74z
wjso5rdWO+eAE8H4kP4YJxzsOFPiT80ZIYh8Tp8TPzVMcQvM5ZkhaY2JxuGRCdwyFmvKqa/lo/o9
/XLo2hme5a4M47EvGXlx7jejQR0zmDiXTfVeLebf2TaD5ij95qAzqXpntbClWieBq5KlBwL8pOkg
0sRx9a2EHwDeEx3f0bs6mc6IXBUVYpCbQV1MOWlCRhENuo0X3Ehw2komqeI8jQ+gkPJ++7SKesHR
KzQL0fD0QXX9zYjLy1GraEa+Gfq34NWHj9Br1wZcwxv9Y8tX8ZZtTI83w83WdOojcHFGr1kQAWZC
0n38TYZDzhqPDNmbQS/tUTUQ2TuBp5GSDkS3rNg7fTYiO/gWUA0VjthYxdsuJbaeN6ft6qzzf9vk
jJFwmRsicJ7wySMN8kdL87IKQRGVd7Dp3bNBjm48DsV7cktprDFbUC9zXzj16mcqCJjqxNAASI4e
LNyyM7Ac3HTQIDyY0VJVoVUmintfzNUsCSMJYjyW67pve9RGbp91tbux7uTLWvKlHnSU10l5Dauy
HGHcuvm+G/Db1PbhJlGLp79sFegRXdikX3dgijlWe48T6rIp+7Nc57dukr4ndSHPCnMwmnWmWlXN
bfBEQlGoj4Btm40ICw0GkTZ833M+b1mC5aw7Ht8ESTxom8jSMVbQho9sGIpjlPL2sC2G8bf5JGYR
7db5Mb7VpE/ge5XG0ROGJKqXnmn2B0ndoVwouBZ6YB+Q2kdnEC2T/hCEdEgrq7MO0g6418aMxqcI
0CJvuzOjSnyQswIzfbv1VLe5fq1fqbd2nFI0xsRQ75MMVMWJ/d01znTAeyDHh4DFr854YfSiZtA1
9jziol2aQPSzMkrPSyCFay8YCNttuBtLdx55/98uLAFC0mdPjOBw1sXsGdiHs7PvL7oVF3CjqRWr
vfY7XbutAAtk7XoXI+g/BVBYMF9RG4ojNzmo59XFZBu8kSTVjkEggtkpBAqjR/MPVDVTZidzz+f2
OJx8sl551KT4/Xl0fGwZ5AO2rEnBkjHyWWNQUrbFAZA8ojIhXG/wqIaXlINSMwgLDOAqHUNpgU+u
gLstRmGy9ECrdKyaKjxmeMRRvSlSSXy7L2GzXT12XvnI9waUphIsfKeRZJ6XJbPiX1VX4YxrV82b
Wr/heyzUxMeJWTqkuJ5pI6QUnYNHiIHA0H6I1apyxAWloliyVAKypOVqkPwQkD8oS+AEya8p1/di
jIsoibbnXpX2pXg9XLH0WixIYUQheOoZ/1AKAEgKv7ngW31sC++KyOXHXL9ehK3/DLnkwpzlDKFh
jpa3+N70WhyP9gU4J5v4xVZImmEjTzpm5fUAqJvl5HEeDq42KOm+MI37PsdiZ1qEjl0QEJaeCWkN
PiD9FAku4NwlFLKzGY7FXZ92CnpiTAD18dbZOzPecavOb3kRlqXA0FftaxIwOtus3dgg1cJeGT7F
3BcPM8vACzZjXWNfM1Z5cw5rp0BK0Qn/ryK+rwte7B8yKxwNN+HrSQEqItFPUBPz+8W0gB0T0qMK
oumk1mfZjP1/vlu9NCnpsaDXuJ/mrBWRPaCme89qtx9bAwf3jbDsn/ohlyrggzbnrc9C4YhS5x/R
RU8WbaU2zxGjR0RX+qOd8Kf3GUuQvjhzFNGS8clEjwuS6+d2HkDK7D/xllE1JhjOVnKisgbvVWXS
/tzoYZb1ub3HZRIBksj74l87T/6lZ7XyFfTi/jvhoJWoHvtctWnHd2VFY5JM2y5NgATRZFgC2CGQ
GPuIzkRk5Zk8hIMLju+QWE68+wQJ4SBoPPyKQSXjQPJdmFeU2DaKv+9VOIPMg6Oa18Bivw4Q7OmA
fY0ROEJ2aXEuXVeeYlwocYuzjDsel+73ZIsWNw4g01JkFQLcj1k9mNJMcTv9wT3wlrmt8QLydtha
byYOyYJkrPLvjP3uhVj4BvgEA3/tsXFwWlhvczs+w7iCS6415T47LmihklIk8nnwZkeFFcFb5qxZ
WOdeiSvNmWjaWPCQvk5O544Q+TEueDqJ1zUWG+uw/pZ2YW5cdGr0PfGvhEmJucXFm9cjgJbbWOx5
hVSfq1uRjni2l/5sZze7gltA87IYXJ08yx7Shqqg+ok4PiO5niQyjAcykrivfkx3YmcGlkAwwEoE
quclbvdaRx2NMFRb2VUDQkZoI7KLDHfloxCKIe0CzVAsaxFVLQgrzJvPqb5FKAEEWz7JlOxqtBjv
KuzH6HJW/sJZHd1q7bGMkrBH3q/JBUUKJFdbBV3VNWQka6SMdpgsIGLRoLyuQCa/0Y7vOIJvqUfo
rHo6xUX/frM4scNhira4gsTI6VG4VGwnVF9WKQLvGPeBz6q54WPic+6tZXfUCM6J55lRuQ28RJ0J
ZzWZ5nxr7HFV0vbOXp0Tp8qP5Iag6WetK9EHwqIXoeRQ6imAX+RQnAY8ZKrK06Y9m12j+btq7nKE
VG/74f0vwS33UjE6UzzN//Ki2cP9+8+smb1T6WL4X3bVpza3j6XYX/GdNhIdqxENUtT/rt/Pb1lG
fV2WbbetYKyA2hcDKx7Jj4eO6kiR53YUzLOS78ujEqrdQJfkGLdPL6JtelHtHs4daIvD19iLkTsc
FvyU4HcT4MIaFu/RdSqu14e4mjLncfZygqCbmTQJ+D4fVCycjeQUiiqEof2hEnxhMsqMRrpccE21
kvMrc9MxhTXtqJrfGW04oobQoVFp2BBQgLrKo6KlSCSNN2UsDn0gTOBHXvJKDCDuo5KG/pKg3ygs
pNqqBctFue+1n2YvGtd7WHhnTxBbiaUKIkZJLlBSaU5qdU5Traksh5IKkgYe/dE9nVD2HtrOqqg9
7LAYhj4Z2dZAIKaHYIJmfcoUsvcFzIOOBasLRpsKTNpLoDIn2VV6RJL7Q8TmekP5sS4Vt9w9f1Gf
IYhK1adrsKN1PjR4AUs3GIE8EPmGzaWuw+JRwvCeT0wxyg+JGYEmSa1vArXf9heaBg3DeLuSPOaP
HdRCkkMjaaQ1E8igYfeReYZX3e7H7w09XifW0tZhI6S69n+9a9ttQkBvAPGwhtfM3Q9KyaTR0YyQ
7Dwr+zOeaBHAIcfWB/5QEp87V+RpGVCQy/6PevOrgNMMxPUX9gTpArl/+7JGluRx7rY1tGhZ56ac
gOifhwIJKP6VIar1Yg17SXSqOsUpC2O5wklFPCWaci9DaTP15wPYl35nGNFheD/IkOGw9vJSchGT
whyBHuUI9OMWwZXcv3CZYRcJtzfw8Vh1bROFZ12u7gtUst1p04iSE6Z9SV9EES9QCuxoJQfJE4hs
ZSrdEjny9DHoz5GZ2kMe4XobHMvtt4f0PPED5cVpiJTRCeqor2WOui2Y+ajbJ23pE85QwKq4Z0Kf
zXTmu45zc4oVyLIC3mlBsKSYBcPsOUsBvdWnstoKq3/vUBE+CUnFILK1hLkKJg11r7NNGZrd44ts
oNU01s62hfGqDmTBWbiks5qxk8OIoXPUy8tETbW/4bCOE5huOFfvO/f2fBnzVRs8aZS91d+h4BDW
9vAMzK5PzAX0OT1s+gwy+13phjRm3525lz1rtr1WR5aY18Nn4EBY6o+mNHO1JU3WNuRFxDa/qxSt
kqaXV2QxRApyMFxG26c4kjHjqQagnBy9FDGN9dkOeEXmjI7ym++ZnJFWvrqOR01/cUFcumRSZlVF
duOERjNmwTzCVtFW82vxijdQKXTAN+sMWBJ07KTwmaQbsArSwLv8HpqXnkexQNgOjB8sHWhgMF9H
aqd2imjgSH3n2sGaLlUmakiCOb02j2ZNDfUvZ1SZOzdBb1DJhdgGT0wUJCw6DRVhotEvLXQTAGGu
YSbW8X8wpO+SZeB8TdHGU5Z4iAYW9WfDQSAViY+zXxbdCHSbeM3U9BlMWW7o8N88atzFBD+gBAqs
pdRKZSJCKgPsQHU1zmaW9v54srXlFBY1C3enxyZhw7j+NYFokjEnlb0mPwHCN1NIv65ghCPHS22i
4+wgjc3skP2yxQmh1iiqnwokd1DBn/9eYKHgG1mf/F6HUEYilKcgFjics0oqEf85adRmAw9JkFvv
bmptLlMXMkDa6ViAafci6uvsyG/r8se4Aoa39kljv7ynRlSEvCUG03AC4ckKXONer8xWrZDhNgSI
fN1KWjCsl0UQCcBs+Trz9O6EdNAHX9vw4tfyA3muDO5+GVPp2ASiboIrBYMuLo//0BEdlXF0zBQC
hBM8mWuVlDM27+qOS4pWPrEAKAFvKCWEa1oqLtXPVQdSnVW9XIIBRILvldAMHUGpDPYGp4rqgoKh
YngJlLQwmD9W+9Tl/4k4YO8x4ESEDuGydy8V5+UdAVRVCvmk/PKp+0DWfEZH/5h73bxcdjq/Xu6A
JPtxSAxFurNbFWS3Rn9z1/GJn/DiKDikC+aGCkEIqf9SZ94DLSq3O7jP2d8wbR/v7Se9JFIVR1kQ
aYvXxQHEt6RUG4vJtvoNL9yyqqj7g71GtSYwNqpxfsMZ0S1WKi3/lO7H4mhjnH884tG2E9HbM3+s
p5IQbsMepjbTxV46aiZup3sZg9UBHbDLLkVuYreb5oURVU/Oo1N2vl9fYDyUTp6iXyuWSwQ9m7b2
WCzt5pRym7mTWmGEI8U6EDE4IDQf64MN5uICNCfu1+z9EnQ49M5pLGd6Z8EoiuXpz5z7zkqbnSB0
rFolwbj/GTBLR50DEgXV8law6SUzlEejudQGmckFSxd1fQeOZqk058B+wuyzbq9mjGrEmN1dbPnO
uEgtKi6BOPwLo+ALWXAsfsU7F5QYKKdb+r/w3kIHzE4MKC6fSWplO5Sl7fGlnUICqAd3fWtl6Enz
y8ojQ+J4YosdDTfdin4qY75yMClBE7ulswuJiBmuIpMZh5tsXSfwIIr57PTcq+VDX7vYMt76wPHq
2Rr5qtAGGI4NbFsjQjijD9+sudP6Ny7lo5jDI7XZNZyWf5PV0vk6ci5k5LCxhpFgARdXL+++pTUO
87TYVkTk7DbRd1Xju0C3jFIDYnEbfHVT4/nK/UsCIpnoeP4pmZgfEDqWHhRTTG8HNNo6+5KD/4qL
fG1yu98bgB1n/yslNY4pgtdCgoSmcDOefgCJCqgXL3nh+uSnaDJF6PFDypwO2OAGR1Htig69/TFM
t/DpU4mxUBsCWE5J2GXGf3EMtvke+dkCddhXFekqSt0u4zT0C+X3639HIQNoz8HluTQ6nMuRTxHR
fkS8lpQTfOFhdaqjmpQDTmrRD3AfndoJmcsvpf6ooJgFxeu5d5mRh5NNYkuY9i3yjDfaFCCyd7Fe
eCgJUjRG4IHZnvvzI3l8TMMNzUsGsVYeZ7fprAlTGT8E0259dC2vqD49UATkLOHlqKtQQBWpU8fK
pWRpUhqG+Xc7RzY++LA/axzlvxDnzCCuhh1xOWseNzUzpcilmwfXHdlGvyKScYzF6mg377bEbtXv
AnA1L31kjilNgMqn3abbVw4tpXIr8vBVheXNzEDi5I0y9YGQq6sGgYb0eLaHXgh6wOAfNiMVtuiW
mzLvnZPnohDcuikWqKXxw/LCkZDthsTAsG9TLUgoSIY6JJD06EyHUAUwOKqDjkLMii3WUMYmP0YL
8mJWCt9jRKDMRk9cV6LKWMQ+yrBg/gLDib5jTRMW4YhwxrIqbfOGIQCl1Xm/n1a0L+2nw3Lkh6+b
T8ZnQ/cX6IwcP1pbD186QgzNBCYiW0GqQHHCqscGUOer2660b5P6Z9BtF4fHhV2lWFTZx8nHRqyk
G5mekVVvjsF9I3DlcvS4kd/9mphA/94y1Je3s+OVEPOASq9sujNu6jb4naeBIpEy+8hV9EB7eZon
VlnEFcFGz10FL5o8lmog/IFlJ2y5zhhw707DR47h6oZaoWUKOltE/EORxgKVnw4ZnrS7VIDFrnhB
AwyjXWEbVK7udIb7fSnVDZKc+m0fDuYAEANvabTt20uwiaGEXf/in/cSWAVkzkOMQqmByREqpKSX
2vKdLxPHrNkbKlyvRGm/X1mHogVpJAKPQzwHC52sCLnXwFVLghm9IWTD8nlrrcv9yIz4VpWKb6Sw
sfXmJ0e/WNa3PdXfIRiBu4fnnTg0wg9MvDV7i53VEURePe4jUA1Vemp4ndZPbCgfQSFr3PjpJ0T/
pSv2Ris9YN3P4dFDpzxVRnu+c9zCyH2N529Jcj2y/s53e0So/GQ1mxrFHGVyyY9H30cICeOaxvGc
hEkF36lIR0KdcChlSV4FmBmvbkXvBijLZQ5sx+KV6U6WEmeELoCZgpx2zU/A3O7+D2cPG4a5GDej
f9+HKnd/hn+2qfO3tM9Z0eKmsAoWB99F1uPK9PzrZ1Qd1+m/UnNmTWmUlhc4hNaus+YjD7aALkEo
9jZmGDpEjO2ArX0FxfBJq9ZlN3eVHZaaelWvDiMW9ecGNw+ooQCLbMfR/D3at9tKbl74lnp/LVeX
xl3mu6EYdHGPapeGi67iE8veqJzC1ELV6rfDAafg2MA2caTtKYNVRVWRkAt9bw9z0S/GerMoDLiV
69ddR5C7BmlOCH1ySTI91ibidQ8Shb9DgnKMOG7ZQ8u0SBJ/o5RJrL1n2J1C2hI5vTWLZeEo40an
/oW051zYH+Q9oY/l0Isa4devkII+5ks0Vj44liFXHchsR7b/ik72NEIHQXbA86jl96Wfb+8Xbly7
yGypzY6oo6TeCNmzbxKWwNTIh6J4/7aBcPuJrRTgG3q2sPmGwo26L4XPDCv9b/UknFmcE8coYyCf
kdoBlnj1urO8dslJoHxaztBjcA3zVZvVcQbfme3+Rynyc8EbqATGLVxPtQtV49gj0nTB72z+I73G
9EcnTHvUwi66hNqUXLg2oOvx43i8V5inPEuyfpgOQe3YpDk4Rf7k5VxkxK6urDLkzo632ZM/HuF3
dKpa3yrE2zhPFnCE4qsts7/Nq1F+vfyz4MsubXq/WVjNpozqbRjyPTkYJ4OVlcKx6unOlslhI9XP
ZdH7gf6bl7A27sEdRKvnAu7KU5sfywpBqs9SvL2BYYwOj0S18yA+7iFCX70AN/+44ffeAYs72YJ1
oV5tr9yYcsYiWi1pRiyKtCI/6D3lrj3zvCOeDPxo0yPU7x8d2QtFEzpSwpftulxmZyVWaYyrjLTx
LyPixcYSlQTurq8aOD4Ew/Nk+KkWgLAa9SA77j5cWVzX95/Ozlr1WMhTkoggUTHfA/g/tSmwUlj9
22NK53PJVLLPttsDW6YGOfvoksqyPiOo+4JmlW1AJ89Dw58Ebi6ZcsePlzW6AUHGgkfXJLwJwtB9
IbNC2ukeyloLZY/zG0VKHv2g97L0hw09jmvnJAdYeFkgzWnPwqZRov360Rk+VeVrAvY5+v02VRuj
HWr26ovG+hjDYbrNVoviDJ4q1dLHv2E76Vlrr+4GqnUbNfl0iQ1emK9ApO9JupUjko6WGD1s/GFR
LlQ3zUzsUOwsu71Rag6kzOY49S2gIZe+vTcpNJutzGLqEaPvtcRj6OjHbsZLIk5wMTMT1JQPwSlU
0my/gunII7TwqBj79E0rJ8J+gAhIdTuwVjSiXz1W0+sGN6zK8B+KSd1f0Y4ZoiFLSkkkIEcL6ijp
Mku2ysA8yDQJqkeOp5grbGyNISnfz9xoYTmD5iIPaZuwvABwh+gEObMptWZoIH5oHXq06YCZElwA
C0hHVubxLJh7FZl9XFabK6hbjO+2DW2HmdeG2v0bqCg7V+ERpiVYn+zqCNBo1U3TbvlLIME4m0WT
c/qj/t1XkvEdMBnhfs4fKytfpP4I0jMbk50yLBBDEi/+yilAdNC6lJvst6WG6mDjZ5b+CkKZLpkz
hFoETD2PzD5DQ2HXqESy0yeJWt1B6sy+EOdo7QI9bMVO/Re2ecyALm10uCVMNQWB4j8VGp9Qfep0
gpbfN80mFatN0njRCNfWBwYCLeLbhu9AwBSbqMbLNIhQ5dZ84CsUAdBuQM0nN+8jR4xJTOhmpp9t
LG9SmcdGjZQDxFN2BuoV+muGcF+XiWwUScRA8hGNNYr2oO1mGXWJa+rEgeDvGs5+S61JEsLlGJKg
LpnOvPmvhHu1+0PByOwp1bD5tOTGZ/bSS5KEZDhiwcKTp/ISm6msNvMr7j6RmbKglgY4kTL3HdZC
ai4TvJESFKUmx8h5XuH7wSeCq4/8fYsgm7T/JF+yo0P0LpChiKIvcyXxWZtcRqH12cc+8SyCxh1y
uj3wJOCx6lAIBN9/u1eb6GPOR6dBFOQe5rJ9vwpcNkTKldNkigmgX8eIDnVFlHahGdAwpX17+EoP
q9RSoKRJHofS0jUfrxNN2ehdZYuw/MLsA9RgvshQEgUaXu7HUtq3OXMfK4Cs08g6ETWfDn46gXHT
QlsBxFpJ33wTnpV3zSEMkNfeRHUB1iyLuMvsIOIR67RX5d+bMQRKUhVLenENeIPmpRSBXEr01Iz1
RkBV3SJmuUvosViom6mGAzW0vBJpZkgZ+XCnEaAnil8j2lzm5vZrCzCwu9N0eDnJeuDGWK1ybVLl
6TVPsjnBpRGnx3g+sEdSdiRcMcXL0OOx5UqD+ZabgaCy5yf9i3kxxIH8aaxKRPLN7ckmGindtRPs
ZTCGafWoXGYM0xLEdPqVRAYYl+HDknf2Axdy6YYla0M/2H7EMD4qqaGs5XJ5nku2BTii52hb/x4X
1mJG0RLRss6o8u69dsNfvJlAE9lDo1f16HdUQuTKtUe3UCcv7SiSLlRIBIukvcsLzPOrjH2yY55f
CQdZX+m0QqKphTl3YiCFwLjLjDb2rfvNo/XI/dY7ePNnr2kwQiKQR9fsDxTb3yq805r7U4FLKzvd
8yX7QfDGqtQ2gduY3ukfErFX8sUWG9k66tD7gwsiIiNFfyNFA62RPwX/I/DiUW6LG0fJroQSJy1a
ToiW0vciY0KNSG9hl/3ZHkxUieiZ5VPUiOAuRYb7IUm3R4SvPRWxwXaEyqJxYEe164L/dZZhY02U
ZG3eW0v5q3K6Zk3xB2bqArNMyMuwz/n5pGXjDau1fh942ngVRV0+Vwnxduqtyt4rNfF66bT52EFO
0QZlpWise5u2I4ygjBAHwRiICm02wUuVXHWx7ad56ozHjFk5yyZoOZFOO2VthFVfqEcYgJWOpqck
EMGi80JLCrC/7cFC4EQF4OTP+bSTpRDmAjJsnMrgBtw0aNiqIyAuaUiUMFwvNUkrtAqMbyIBsanW
Fl1T8VSAkD+7uz3xDWfBDCni9N00ZQ3HyEzutrDutcfMjP28LCFmuN3EEgkXouPH+Tvth9fDgUJI
ztrzkVNBzAIpcsjVDVfwwqCZkbOuNGlGztYXs4boQRg852UKdeIFU+o8KBIK2FkxOzOqUXRaoayV
MoZIxSXnlQzMG3iLlXG/Og3gI7Nvfh9+Ib4jrj7Tm77F1FGo8zlQG2tZyNdJ6rokPx36oiKUA4wx
w3DPziEyaWqBxv5kqtKwdFFHfCpwCTbezhFZKAZReMIMZUrpz35rzaW+tANjWUN15MV4sACd4Fv2
uhddOaheC/bWGSQ3bfm0gS7yri1EwrQJA1BeRT9jz6Mdmb6NTq7I6bK9vgVfAgeAdZ4e8RAnzQDl
lf92bhgGyUrm6WvNELLEaYjzNEwJr9G7SXxVtvJLz5kOYrM9qG4ITBrXfUlp7ydPxOXL4t55+2Vb
jY7Qyf8LxFnJFtRguiH6JQKluiKoxJSZvahR7dgwF10ktngJwQByJPzy+K9WaXYKZ1+DEyGKcfMu
KExLGBWtT6wf80NAR7/Pp/Smp6+baojjqsfGX/YL6dyaoSHIYtWw4Q8A6CPZ+ilq6x1SbrCX9Kqs
aKjpEYQnONVrDVDe6G1oIT1mUsDOM6Ac8v6czzJDVRWz0/acevF9x8nhtUYHt1gtAPjJRidVfxOE
Vqvx/b9QOECLkMolmZHYAZdmWzzgG7nE8LYn6CfygX2JIbZUhVPXATyHx8VkTwsl5sdDPJU44uYB
tQ1KVMfeb9ZV5tO4B4VdaXQY+LCkDqSCzBSGwFQZm1UQ65TBxXXK9pAec2ipxJf4PN59WHvHgbWe
AqCCIzjYxyvQ7pa+oOywzOxhmRVO9US+YP71Js3cjjIRPsVZu0xrd+Fut78w+eMFurp1K4eSsa/8
AV64Qx9fF24HtO4YeoAj0KuG7fww/7w2DHu0jPjPCdf2u/97tcO7nn68YDuNdTp/eQVEz6crRFVO
sl+nrdxX67J9LsOsribeCcDHYRxbOzaigl2IF3hBHw682qYehlDgMgB+doMu/IYynjgW/eFrY0hA
PQJRUMFtkfub28iOaDcKoQnKeyZ2L77aGhCq6huRpNC4ztXARCq6wTeSVyXmybjAkP09ivUjKyBv
3EBzqDNpJB5SrIYXCUfWyJPKDEV28j/VIVj1rV4rLiGnvy0XGbvK7lN1R4zPT/KNohhl0zyuexbW
Vj/rf8qEu6Btbjz96gNX9bvM8kxkqBfvJh6xzGW4WcjaS9kTb2n8iJJsu3ddXgenqt9tAChuPoP5
biHl16Yu7MvZ2IYqOjJxPW+G7kDW6nn4yFq967FYQNC+LVNfvxwnSkPds0YLpTuBDH5NU4594vop
Af440sqgzBRvjcFwjnIcvA0Sgo7kEYfpOsar/tNtbJdl3/rNBH2Y2WjnMarYASH1s1tknaFzJZa8
WNe5Old76ilBmGoQjAQUVCjuIGUMS+KRt/JI6UxQRo22lVj3y8gbOotfPThMoY4ZXxuyPmpyz0Qf
IFdPKVRmv7zfHw2w3mfYIgIOB9HpiGPFwviUZYMFDpg5bcirbhgeKcMaaFg8Ce2IJ9IRZhxO5w7b
w7Mmgfe1Uu+Yl8/BEhh7GhhOSyRxTI/iXosnWQb/lygFQ22iDgFM5Gt2C+uST/1cRKjgClziCdfo
M76PPHW1+FVtQk7vwImWTuKAWYNTyv7vUVDVKqoY7mkMmE9HBxuHA6kjKnQhRP+d1cf35Bo3ylRS
r2PsH8rppiFiAOLII8E+E2KSHszhEUrVVVX8in9aqdJ2GuKXzpRzwPQzq6lgxm4Du9UJ4YBKL0MB
7EXBNV5L2McTP8P7IXlRSZZRNvq4ImdBBey6st3iEkPxa3xdsXVCxiX8+QGO0yami2oTNBKelbue
dkizUD0tUD8oN3de2UCuWcOFLBVYPED0nF2U4vz0CxXPF3UItO/twn2IaYHexQP4XL6WWQJ8pGwC
2v72Y8DQ9qC6iNsGZOmdy2FGCCXDIWYxVePo6YAtff/6brvnFo1Iovn6O347EAlDb1cZj3dFl8Cz
LY2bA6AS369uWoSAPgnk4LvuR8lT/SZt+D2AqLD/AjnWqYW7l06r7jJnSLQgz3ia3NSxhwfjKZJk
BQb2rKQXJlRuh0Orev1eTdN1b4hDZINu6rAyozlYymnsniPdD8e2QTYqeXheQWU6sbRSB+CR7JUr
FKI07hdIlfXcj7V7Vjhgq5LSgaFOTTVwwlrqcEKPGvRAx3t5wEwgrLnx/yqHKspiUW5SjZyzvjBT
lxPzwmrzSKkxHax3CAbmP3NROdEAPmyNCwv2rO18GWqVGWdcsq2VeIxb00HtFIY9btWoSJDi3qAQ
bDf33mfnH1pdHk775A9e5j2Ckr7TswLGlCHh9TwZrusDVWDlrt/5d2ZWBPDlFMzlinFpRh3Kyd8c
rqWS0OA23D1HIgZIFbHxoOIf0+zz4TDgVx1GZb+5CJ3bQ3b6D9fLezEmuSPBGbaXRF8Gc+FNjkvf
Z8nhOZgAFW5EjomH4PtGrsmxPhx6a9bP6pgZK3op+r+mSBs753eQ+F+6H+6ZAB9Xw2g+FIFT+YGp
XKQeOhrym7tJKjgmBYZFHrwc35EdCs/qdm6ek5/UirukHHPDVAN2DxCTRG0p/ZSfX9l4/ySFCNnT
cPrlHjoT6J7XG8fPI1BEjESABM6BOpWE1bm+7fPh9O0ybeddLzUjuJOzUgChkn3Oo2dwMOYJeaE6
sossdRjEj3pG8nyba3rPo0hw4jXPqp2H/WC07yxC/y7K7QFfPXEqgNeUhQ9JIrdgxY32SZNnR7Wi
lGGnHIInPPcfLBUkLPYNcfT1umANc/HDZx/OS2mjWfcnfe3c5JVN3QUeHHFleiqICpw2webJeMku
KaMZxNBbvAqSQNM858/JZwcIxC4WGPYMpZV+NgeY9zbtyEK2vySNf5I1GQ37AekFjJJR8PWFQLhj
qTJjx4yhtcErg2ez/IzVjiPkGjUD4lU9egzuQe4ntFLyvrWhvw1YTeG5gZv4DAupH9cL80uVVa5O
SaCdvMan19Uv2G5rVDrabHx0QLPp369UhV92PitvxYP2PeEsAyixWsi0ZwiP1XDDXo0CS87EyL+Z
qb02x9x97ejaxa1vQH/L6Jt6S382b8s/zDdGOGUNlE2t+p47gMjrDDb4HTBWArMs1HKOfch+YUAi
ldB4uV1JbZzp5sSw3wr0vN53htYXBwX5HCExTlrnxVaDmvLQf9E5FyQzPhDzxEDBnDdx6iErGku1
MR+xYFtupzDQuXfWvAOXJll35JdTN3sadRJTaKoLPuHJjVuLUXZIFAKwsZg0GUpXA0qrW5nE/N77
ZvL8Zz6Xy5769TKvFslXUkUR03V9KL59bBfdQkrL/ik6nALNZP/z7FnTMIsQqIFO0f2KbOOxOuKw
MG2cvxH6W/wAqHqUiWcRIjAjgmIDvaYeHfP6MeRUme2GGkInUl/pKFm1TKktjodgtmPEatJToEVA
FDtZrIDcTUmSmjZRGrmFt4nZjWdfphcYZ+/HTO3pNF9/zVR03L4PW3eojvEOPqy8t4Sa4Vp/nBAl
pr76klQSZVEhJV1XaaQ1fsQGBRleJTHTTCVtHtB4x3c1WxjUo9ZBLpBySF2cAQz0Im8qpZXASaPG
T4OwwV4Ta0J/rsoBZoMPqjxASmVAfGuefM8ak5bWvhk2qHcZG+xBk9L5IlU+PADhUXmLo9I7rTlW
rRtcIr3TiPPJrsUOGqzP2k0nDH24rHCiFwUkCvFDlqgdSm0oqZ0m7QGqqYVrV/Rl3/1kwmHYVeHe
y+2A+F9X49E+32HSAj+lCwi7f+OadIyO2PE+smCqfwhRGCZJwGfPmjRVXt7GEiCi1fXj0XmwHnH6
AwOT/cOMcUrAanRoeSA8PnbhpE3c/triRQsp2nUU7zdFoIcTcdMF2HQ1G9pC6XWcT07M1L6Snedy
UCjo8YfYZIaXgPKBO6JiPmk7mI5iJaLE/G5v6nED1uVjKzG8wRprwsI664SrKx5Jw2/OjS3Z3Rkb
J2uji5y9pV6aZUYb/A1X+oKzuDa2kJSsNmp+uv3Aec0GWuU5LOItx1+RXZCbCRiMJkXx694UNbcx
q+NBoyflQEW8qL/ANVT8JU81NHraDsnXiNINCQCUokeGHjSBpWmgDsNbwYjnxkvlyQiGQKyUyDKF
zwYk3XhiMIsvCeoUqm2WSYCSpLlejEv4dmdVqmtOmyRvf2A0RbUWTBMTV9N63D7p/YOVaPpAs6TD
0AfI4+xpLNuBAzqZEyVpDxG3kmav+YPHnirS0rWcPRgaW11PsDMlycvJV7YZknc67Bw69f+P3hzM
F+G59nTJmrc2qBA4pmiujZMzqVH+AwM5/3BrgryxyrpP30VzRQU1kDIxoQBiZzLFYr46nUPYGAUx
DgsBuk0vfRRnnwJ2A4xA38w1wopLiQ2QmltAc3LhLoT/yYUlMLgYIWQ+6cnxgOVzrYu9rLu+DGqn
ecYeQh0q/iLGCyh5srd0gAKF8vZm0hPuzq/KJiWVY/mX/9UyRVKm3sUqoE8OPXtvHkdzL+XFWOSf
uvboy2CmPRTEGwhJ6f+Uit5sfAWX9ajHq2uPrx59oCN4nogDXlbBO6eomutLMXvXXD64H+N1TmiX
urXsR3mNz5dfwlaf9HZ0Sj0vMu9t7RViJ5pTEITU+/VyHGplCTbbPannNPUNzEHrheaEsQta/FTi
B3FLrX0fzQWeCpJYLkk/4TBcFMqSNXYWa/9RSuRkf5+HpmWm4p3upAwqDK6Yz9w2L8jbHoRnK2II
BaCzzeIdw76/SspqUEs5CUUGozb9DoMziXGazFTxhSitgMKjY3YQCgLeZ+ixrGqeR141Pay0ehVi
/s/UZQ0RSAX5sSdGdjY8jbsvgmxtt4z6tXyQh4RvJ/g0UJeQODQuHKk4WrGcAx1HePYB8nSiTtua
r9x+6Z7hVcI7AnUfmyUDP9GDHMyH5/0i+x49O+5KWwk9Nj6yQR81xdyjHyRc364mj70IS9tVcNkc
ENARZymz5lFMq4HAUtyVuax4zUqiT9OzydST6KUxc5D+5NxOKEBX+xCsymXthawISrY83v/q5BFn
r+cSY+ZKtslKhWDdl3gZoRj+rd82uEySH2pgevF5QzlpmXNd7KezgS59/kUCPliRv67iYKtClAIh
gMc+mWuu2MsTqgcM2bRS/wsfjIi1CV1iPKGSvDS931f9bdcuRYB1NP+QxQbLP45piEBsl89n75Tw
AjVeMDDtgsKFzbXOuJYdynl04A1oLMxoD0KQBBGy1Ydn10pUtcuwv9ZidLM5W0hYCbFAGZOQC+7O
heFKCtr9kPAZ1PoBRnVDhXqtpNewRPISSa9qieuHuaYZlbQ7przFsP2/dP8uk8SCF7ADdYkG7NVZ
tV07zjPgQ2DNF6ilnUDZTPbFfl5ZmOYWtckrgPvylwZiRzYGqLoaBIV/Jq1QPGJpJZX5AY2C3x6S
r+0jI//19z/Alzm945XHO67qGHzRxV9eXslTtKobbswuWzm1fLhQGfuDvBtoS9ewX4K9jD3AEzCK
h8C5AYTpR7xSPrp6Ttqswh7oXBjR72EnVxfu+RiO9f6D/4x5B9dUVymWeY3ishvM0p0hhzz3TZTx
83324JMajUhpX3MZB0SXRzX0V/V4NcbhBd4NzYpHastzmrkLoxcEaZgM5Op/elqhA9eTqTC6M9HE
CygqWjwx19rw3Q9GvhExch+J7NslqrxAw4chg8Gka+kqkRaEJHpLkuJKac4eW+k5ONBb62UzSC79
1tl45HRRmvsVZGkl1dKdHdE9KUBv5I028kWZ1kb6IFHBnLqwTONVbyVuXXn3fK/E/cXMhbHVFgGo
vbrSkrnuZUeLjTVNHVxXBrfMFQ3qgPHMH5Vq9NM6WYzCkZeVqB46ncS8nUX+LmS2A+6yQiFi4eEN
iFkVvQXwiLVkgO/49kGxRtdd1n8cMK92WUOGnynauie3fsy7rR764lR6eI38SFpWGB4c4vDvg47C
PdnX8pdQUoahtjP+W8BCicDm3XmNfkfI1fuyo9JI59ggNxdtcKqSF1zSLiDRJ2Qo+XahrYnNtv8O
DocollIl/8PcXFqGQH6kpsij7dl/zCV58vUzP6cISQYyod3cvVUrfLDXndUizx9M9CXxircuju8Q
rfAjVI03yVXz9axa7XgetK+wBomyP0iYdxpHSIyY3O9UMyAON0ZWrL8zIF4kK/AUqR/Ptt+VhP1/
9Rkt/q+umImTrK95D4PXZQh980p7XzxBH/LZfjCZfYxzBQHFGEjrkLCi71q0OmFI4lOi2j4kIsky
d62aFOcz6UGw+ZQRi6Kc2JO5Kj9PR4XeZFZa7rJbQZnxhgOBmnlScQPMfroLCSqtEOB0QBMJfokU
80Sz3v+KcW6ZfeP183d/FFBQqQ5Gk//4ScEIEjhZQvnIjhWNFtTmLfHqf23Fs/XM+ojr2oCFRwPs
9Q48oNJtW35xcRUc5DNb/3f09N0euq72Mo7EuoKXeyOM0ywZZwR3J51e/o8xldFLRFV92z3R9uKg
wVDtNIhKMvGgsbARgAr2+iIinX/o0/DTU8FTmHmXcoaKFV3QrbGxKttHFYq5RDGTZKG5f3zryzz9
mQtQIajxvThmXtT7HHwe0ofmTQT1tvyZiAiBFaHzbbP0FL/XlanO5Um3/uSY9R6QHp/3pPDSHzJz
XWcTjz2tjg5A9bR2MSnWMs8dzi9Obz1I7kk3vjJbY1necJQ1CACBpFROhP7nJb7mVd637GhdvKWy
gHdKc6m+0Rw96cCjMrJrlmvVN8a856t7IKv1sC70UjvekEUAkqrKscMQaz+X5nTwNdUCd/RrLd+w
vZKyuYJ1NKRm6p1x405Hf1otmhCF0hCnJ07Fvr9+E/akgCDjHN+4ZSsJtBzFr5zsZCaPBnRX4xGv
HY1VG7ChQrv5uadJ51TXLt4xY1vO8W1WXi1VjdnMp4KoHff9UA3SAwLV2WrV6Qye85t3hotPGV0h
LNB2ChsJ+ODYOK4GTc8SaOc7YbG7rfmT4Kuu6I7eG2AfkntbTEzmb0lvJTZk66NEWaS3cUAn3/Mv
pGp9YR3usJDIxXZIP4p5KivcH5RDkPAPKYnyLy4tIkAo8TomiGBooxoG+Hz/SOsUFtVphJWa2DrR
6xhm7ag839dSSlbBsh+0MQN+wscbTyMh63xrD53bkkjo3Evlu2My9n4BIsKdSPJbWyG4gdCWd6Ed
yRGCs/tZW8qw5dlHfKAL1WHEEtf83u+MQa7j/E75eUCdHEh64knhXJQg5y2Zb/MT55rjsBwjM+sU
4vkQwexAMg3EusfXQrsN229G3l+zINtBt3zrxQWwvmLaPjkbrhScTuRLyJ9QC+EMzoPEX0IKu3wu
ZsyktZtoNC1l6b1eS4fUTFYhVxReKaRw5g6nN6ozL6wJS8utqCxI3z3nqdSXH0kPMcTrDyOUNp74
1JqF67CFzm/msDjtSaY45ymwMv9KtVxr5Tdv2BFA5xjywXBrAlnHzXpK/dHPKE56lBp4mXi1t27c
KyAacxxd29xew+JGshaOrc4pybeQJS62azp87fxq4wbvSR+iH1nyBBAeF4BXbpR3meoyIl9gUQ2v
fsPU+0HoIFEt4NIC3nVs0irFVmGE9NFC50bkLk1JDMO3faFhlA9ewIYV5T+VJQz5Oxz00sDzySs3
rB2uNZzU04V8hX04NcVK7d+UL51aXKYup0I1+tVEp/FPWRuiIVAH5uoVWocPAOeq8klIxrZaX5je
Ml5pQ3ceEl722o/rehCuqDJrcYlu4b0a0e3N5XzFKdGlO9BkiHkFmmIgg5JSo/ODGbLcYel5ybwr
FMGBlSv9tIdJQpjx4nZzjfQGaIefkUArqNRyGyW0oSC9pbCW5T1laZApwL/OeJSj3idrgqbgQJe1
yGQPTy0Osrm49PCg+/ip70/ZMGcskxRAn5g5jvrCT8TZDFliklA5eAZ1aEQcNn74NSn/ygLGq/bN
Y4Xff400Wv2GJOhtlHjlCIBXCKriz5AT7AMn+zbnj8zb/A8+C2H14VIp8xTM/0XpQz3ES02+xN2G
y+idmntVixTy4UARM94dYggO810ICZAb/xNWKQGkBl8IyOTRMeWcTuvTJrA3VYYemfkritySON9y
ohZsVFuSzv3e/IbXH0zTPx3jxhoY+GVqSFIY84CigHxeODpEV4xjOTnZMfI59jgFJdesom02CVdo
F9EDGTOs75YK9wYiG+kmEhaIpYzmAr9Zy/mjbixoGXJUDfGpP5QrbxzZd/KTSf5KN5sXLvWCYWGP
d2Dlan2Kc1tMdW20Exc0zuSRVEoXaZoJviz8xv+xpiaEPTDug7q434cYpLimW+EG6DZh/DtrP+z+
IkgKBBeJSfMeqWd/oh46vuea2PIiLMmE8NQFiN/nM4SC4ieKX8IYH4rhsEYx9XOYmV4hs325db9h
r3tZnvBG/M+U6iDuMrByBy2793eOvXWjaaxGua1fCbYJNDULax0nGnbp2mxN6m8gc8GDgkzRPKOj
e1lVBugEMhnXXqz420x1WKI1NlP2aqTnDRFIsLc3pAOZHfrznMZon0RDCXXuepKXCAz5V9mmGjPa
38Yq21GbZyTuKYfPR0kBwAc0uA5M8Fewca76oq5bHpaKcCwpiuWmMlbJKelHDRllzj/BG4UBcSXt
DX1Z4PFTO0ed5AsYP5s7QvdJw6C4yD3dhIjB40GTrt5OC1ey+7E3e8GD4YcbkjINpjj23maAKmAl
1DVY+f2j/v9qQkpIQSQeuxaDJvf7/NmUiAZ8EOlhMfFSEPUpvinnOmtpt+qjuiAH2hCEbI96tB/v
4sBK9p/R9mwJchRuBLacFyTTjzRC9769in1Yvco03x5TqHUqiT9C65i0tDNAt/ntX/k5eckCxt05
QbX7SXjvAxESdmyiErZaXUJsh9x7LQvU5/jLb5zJV6B9v8l6cmYcEu1AGACBk5+q5zTT4X/OrohA
wNZXik+JSsUgA+WExp/j8Q9ADguPBjDTljXnYNoqp5VEylDfpt4sj+dhJ31dwx2OnA4b3CCTS84b
lUqJu87tEXdP5AKcR+mV4OlrVA950qQleZVGpHcwJSKm25alsPZkErFBJlTrhB7UDi4OTConlv9l
alLQxkMCmRd7EyKh8hi6SPu0v+FRUYPb4jyBmRcs5lypkp98k4n3B/d/xYqC/X0rU08SQg5bYmsG
WzLGrud1f8M0D4wewSwxxuPzAI0jl/wB2T/IQoDKh8lU3LaTlpKZGVvQN+LlZpKY90COUq1b9KPl
h9M0fmJKczTEsAYSHK6FObMhFPnslyuHRUHEY0F8AgJjuckiiLBhN+Obn5H1WAhNnG7NkIaeQEKQ
GPpOdbU/yU0OlPiBviKesQfVPVA9aJ2pg/zE+GZizCm5p0cgenPvTXv/lelhjdcQJZYW7iz+cuSX
CLnEzkMCTIAOd9BebkOlXlbro+osX6/RGXTZr3JY4AdmeLaSSlHtbQOV1EKwTCboD5J6Li4orSut
ZRQbMdH4dbR2D77Qiukp/I7hc95t8Qonod+P0QDz2uKqPYqyEwOknfMRLQZrndVcT7qibcc0SI+U
uzFZg2cqcTRDCtA8pm+p6/mPrXmX5R8J2eWrO6/Pgs4jGvXEZEINJCQiflH4CthQdBy7RfkaRONP
UCNOFWJyGcY3Bk3lsAOnAh/q4WTOV4hGq+jDUQE080uyixb17hFhILtx5D3YBs80uKYj1ENLy6CD
B0X+1CDutq3OYLOlZLmkf+86zSsImnj2mFb63VodI1WDSUZZCHDo3qlmSZw/a5FSM2ux6HYTvIIV
5Dsziuu3DljVLWkgiyJF9+dGCC0YEFLCU7o48xJxxuAIcplhExth6lshZXIRunKIvemwffrg2zrV
/nctsxiPtODXTW2jN5mCXBXh0Od4f3GWfB2WebSDKOE0KQWCTEydaPf5AKIxIMxBXeA+1GAgtlYs
i+Z9+Gr8XotWvA/4OITHg5u9JSyC2AWOFRBLtdYAwE6fIz+VrBARy574EGNaB58NMM7Ek9AVCgKY
B/LhiePmLkOUhfL6FF/ceF3RmwM1ZHnZurHTIyjOeTjSuNGvRK1QT/Wnu5OMlsv/+Cdlc6RR6e/e
JmwH4MOwda9DxFeUbch5iPqViKkqYHKM/p/C4K8w/4qsqaQEy9L89zXltbNivqM4DrK80RwdOFLY
E7L+ORcEQC18NCTWpNbaWLw+csulMyQPNxCFC2dWI2iowRETrwgrqz1WsQP/6P3wL3l2KrW+7Y6h
+dBhOcILw2eMBYvTE9OEF2OILdyYHYUljeSH4CZaTZ4GNg2uglOSzp+NusnFuDOZ8LhvoprF8Dmh
OECDZVgc6oRxLyXibxaCzfNWYYs/AueHvB0fkCgn1W9gTty1kuhPb2pJ16yI7h2e7VcO4PgzwLn9
jyqPrI3XIFGlSoje/ZaoWJfOrJS9+ih2arq143r1AEbsNqmpASuaVj2Xd7tdCvU3Uy7luSee/cR9
/IU1tyazsNDQ10Jc8oCDs8eBjP36j94qh6ByHqS1/sIyrpc8Xl7ZJnb55Z8xWTGkSbWxrw5OjjRW
fMvPfLGvf+DKZfSlqD9pIK/QPss5jZ/55enuPSfRQqcDdQdRw36V1tY4J+zTSdPb52zIEKtGaTv1
lM2jz6aL6psYoC9F02h4UKeLZh9qfkJ3vDSY6kO3Ct94Fe3k+7hPVT6q9dqvN99lnpeqcgvHvwms
5jvpLRlPNukM1WeGDdBSnyCdULZCEQj3nsft8Se9LgUT8RatiANNXCrbj7WIBPne9wGfkbv7xi8d
mPxv9T9EAqM0LWyl8tzPcqzl/AH4YRbtpsT3urqzCBWxbd7/KBrPlczJgHBKKZGYt3zKlSp+l8Zk
Ryx4WgaFq2UuwDBhywkG24OzDidFno/s6TySYzun2Du+Ia/cxBNfKXfNHKV3UkLwCdv6dNl4fq6E
A2k8jjJ+ke7yub67wqGb+NMAoTjFHscfnzQ44+ccDeoz6S/333tSpykmBsDyCS8dHOhz+tfJWtiP
kwUcESSJSVx7mNdytNJWd6xdPE9y99Lmm1nsAJmuNttuiL99sHvuQH/+JrfdCjPwB3Fi6t/l3cDK
SJHXGwcNHYciEhPc7DAMci0/KypCcOTaaXnZGRaVGVjbdIInLYPSRLmoe/iW5Y0DE12RkPFjRF82
peIz4MdvxFyYeOl2KPm3t4tPN6ahp47ND1dRgb+BhLuVIVp5PLM0HEkcfj/1ija0/8TNRLK7QOWP
QiRq/zVXEu4mJjvlG17EXGb4OJrOcpmGEX729VSQT8KI3eCEiPvKPltPv8dWqm8JxPetnGH0xVOP
nWuwrR/9LVPjXobz3NWuzl0dmFRMSnXZN2xyGHGRtweGoM4xw4SKYiXQ1UGHVtdDYkcyQiTTmjpa
ZynUFaGIr/WQwxgb8GI6oxdwyBFBxlG5E0sRHuu0Knypb6K7Vqgy/m/8IbgdBKDrD6ylKHWfQp+7
lDHaz1MVMCXu1cu5j9eJAFnvsBbz8YvTazOYbjXjr4OMKPgqO1dFMpyWiWvyE18yjRf3UvPh6Qi/
kTeD2FLJIAgTpIEpRcGa7SUreVZInX5VdbGt1J6yoYGdgl38bCvLHCG6r0QmA1wL1h4HxFSPZufl
wuioCTykM+Js3S6bBzldaMJuL59UXl1i4HRzH2FNuOBGELC69qo+ygvxHOWdKTJ9dB3e0ZMYBuBT
o8M9kgxHJXjTtjGAHA1p1dvLKvJvSlvFE0pPvTQBQJo4g7nxWS1S3XxB5cqdL5OzFzG1jJJj39so
igU09+3MSMQOtSvzUqBPzggbve9+0iiopCLgaN2j5nssh0WSl4bnyZPp84gu7UcVxJWELcz+ZSnC
UTPqTx99SEzmOfgw3EEvJx8914mrgU8v87zd1mjI7afJbNtRevz2/lhoWUxoNSa5/rWXG9jbsy1r
qEDYee4TMMuPdVaHS8XxBNkpzc2iLKEhnVcZn1RxoYGe5lb3ShCpx8a+ELJprXpF20y9/6Nf0i+x
s+/95WYcT9w4ZN7dBPtGlT37Fns0la1TEWFlSsv/2Ho2f4ou0ce8xThmDraGxsLs/FYysVmj3JiP
EdNGhRb/s+S+fSdcD5e0c+kl6QVPfbJL3QKubgNRmRp4UkeaW/hHiqpGGvdmwEmwVkSNciUA0ZBb
YIVVEBKnb/OpZxmE4urY0GstI4AWX4o4MLxKYB87m1BlTPyKXlRpUIcHKPrv0v2AuiQWmVyRH8xr
/Byo4LIH2W79zwHkzsFspfYTFNHG59MSuT7aqIbAfpLofUTHP9CqTEJAUq+AfGWmjv90wpSoNrOX
OloEV9m2mvBJyl3KfbWP4NPD7FiTMtxEUZB5pCPDlnpM3y1T1XALgluY0j7xbeX1iLfq05VRZKcl
DUYdoqdN0Cds3SaxouoQF0vhAdrwRw+7UhD6IisaarkTxGpXw4WJNa9GQkGjz+4tK4mfn1fdifby
R7svLDSHakJ7l3yD5bPCBirgwx97cHKaCMaTwKyHY6pkCXE4RqPtMoUbA9PFi+fiBY9xpcgjcVEY
wLFuiRQ5HXdCOCdADiJiiVNn7WZFNr/MydRUgCTgLna/SfJDE7GcmxOa5DTMA4EBNiBP4HV+DVn3
N2tfI0wA2nh/d6zXmtHfQbX2iL3mIS35UYqCXj3Ihg4t4IwlbL2T+AwY1RbWBwPYdiD1elH0xfPx
2z27pYw9AEfaAqluMsWTnu2k98pJeaqoU4Hpio4Z+GdlFMo0xElxUDgGwwNYqjAvjnXrjj1HSIjH
T9TFtzV2GVpRTYqLGaBpFkrquc4qitT5/k7wX+PGUPvk2uvU8AYsgKF9F9BTpyuVqZDAOcWFoccP
kxxIiejTDOiyMAK8HmtEyjFZW7lSQ4esHRyzx/U7lEWk8WQv7ilEj3p8yZlnf71A1jxnxBZn/hug
CBDuTED3CUgfI80qQY/6hfpnRJJvReRLZNbyfdtCrG9A7FwdZxw9V0uROzPk5A10t3l8o1tynXuu
oTSlxpEWTcFly5Bz0ONgLyFYR6IqY4/QXjl5knSCkaPT1yFz+N8GP5lnzPQw7BaWNlhvvGv0LjYv
PuUo59JC0lZUcTa1G60PfLe0sjuNldIQU0Qe8aNe/Am8wx6wMQXBXJ5O/GPp1Oz5olQq27Jn6pKF
EzOgv0ggQk9hifQOTM+76J3Ca6Ck+Ge98eBmmSNB3WcdRW/5Cfr4ViqoLRgBXv44AVBZInh+6sjk
p3IZGXYftH4ZID/JZFTtTHXeJ9CSsMg4mFo6js2KvsJDWjCzTAlfuiKxgEapdC0nDTOHoceywXBt
lOdi5YU+fSF2mhhMVoRebjLY6u+ii2zH56kH6CjB1I9ExOL3S1ZRZWMZSFsjFOlC5lS/GW75tcLH
3pABfiRL7xObOodAC2p5XaJ2CnJsLmVX0tWQ4dQZ7IFNbJTkseZjkj7u08Xs80yEhgkEua3gsJ6n
Dv5/7YPsaWeBGkMv9wrxd2DKn7Fs1ByhfUqbkdHWMNmLC/2/zUa3AsB7jdwdR/ozukKhIGSSB5w3
eBn82DtE1UEspcDBM2dsMmmMIwsfs1sb/lXheHHl/EG5yX5kXj4ZEs9Bb0xB3PGK35HId6feAWBH
56U4xDAsZKe79ZQbpd3y9VmLForpD3x23TrG30lXfYzWdCA/LUshcPrgDFZCi2TUX80EAsb5NgfE
5sJMlRVXQbnYVMiQH6coPFXQUSZTtZzPnga+2FiSEjtWwksxhspc8lebDuxYbdMiAYUd/whiHto5
ijpgX2AdLGALHH/N1p5KWpvPZzRvQicvOQ6g8y718/TThmGKpt6SW/AECEJpxmApljJaVZtpGklf
aBrRWhxshsr2YG0Zs25af0L/bgIS41mRtatCU+RCMY1Y+06vJX5FiTiwrQPNwsx8XRYbXXSyAKpm
jokgNxMaEuAxVN/4aqLmP/FPmC2FCVZx/ceb4p2X7CbyOUqND2gGrERsbcUW5kThfUucR1ilULI0
NgqA//r0i17xFDz48wCI7eqsjvoAcpEmEiXahxx7nL+KkqHC+OyI3wYDlTYU8RE4bcJmHzkc0esr
XzRJ9yTa+CxeaAlOsU394SIzHvEZVvgcbf8a0WSrh1PGvogZq2otemY0bJmykCBOCWEEhI0F6cQA
1OETk3q64VBjirVn9/W0nBWP3bR36ntUmWqr96oQa/PzBIKkvb56mf8CofGbyDeAUWD60KhvqgpQ
lXQNmsMwv0sJIAfDLrKcShNjJe/5I05R6oWegPeh+AarqrkUmdVrAGfB/RBgNx3idrQkjw3kTfC6
ApnV150rSJOsrVJpruSo080p/JpYOLjwA+8GhzU0kiaXAjI6o6RwStZ4I6BZ9EtNuYk1FI3ey78I
wfCioXJoHuJSQl+xSei8rk9lhHRGkZO5VPbChLXK15j9OeIqpD7LtpJUMqRHlMd28DJvT/9GmnON
F8wyT23LvScU4RFVMijE8A8Nq70Z54yIXJncUWLkUe4IVHAqh+73DduqnDOLnYoetHolUTsnD8tk
rWNpeWIsJa2UxS8hIy8FCXVRAWEcLGNUPQ3oFu1j3rG6v74SWltkjM6lnwWTHOnz3Q/kKMD3cxbp
MY3awu8EUio2l4F+bvyzx6rcNyRqdct3ExvTMPRSmZKuXXCYRrlntqsZewU8r+pnLKVyRQ3zXcHb
1qjL0oMu22PXlmsVaYblLAaxn+2jNbyF9+BqsCRh2ZNi8ZEU5VRNQCX/Ci+fW/OzBOq7fMS34XNh
F7+eTBGVwSz96tEm9683G9KQ2FXlBFRp+yBATRrapgI66OJlZJVaG3VlQytICFS1TGK6KhF7J47O
I3UMbtlLTuTneUxIsCvSGET8MQsWqeNKUwZDU+1FkL91FG5bxk5e0bNOlWQFyIuTZAXlzrFarmO2
GNVejQPN2KghKXkD9rXKEu9RQByurBm7xJ0+uEYA2FpvHS5l6XebkFdR+vjpbe/4rWRvfink6zst
Pzt5qqwxkkOf9VzXZVyd5KSo/AZMmisw7K2oFthD78Gcwr4Iri+PkoLBf/Awk9fO9NlGlUL9/trH
Z6XEr6Mgjh+reWib3RhhbHhiryPZrcLkm1tzBGyfDN8LbAckJIFHZaMxB+5D9saoxq8BYgQPRkLO
9AaeMu73CAVEKzQ3ZB3WR4LXmuhOn+NVWADOsGp+4QeK6d/HSwvsemDyr1ZFqD0yik1f5KgFFiLO
V+jPlvcwR7muLzUkJ6zzW3Gupb8jX5gnUePfEBxz+R8/25rKEq9m5vM3qZaO2MZ51hKYKObXeisZ
m57B8HOtd/3FZUBxOJaPGjJS/ukOeWRoPLH38p5J3B4GN8sbV8gQfzI+U3LxkKe8TNAxUO8yoY/f
fFL73JBo0DacnlMy/XSobfMIjViVJpFY2JwptjNwSX0fIz9w5bj0HZ1oOsvqZwMs9ia2avbxPs8S
tWqDrnLeVcrKutN+3tntIW/UKRSCcxEE5ivFCvl5TnnWISAwju/7gOF7MHspHkkIvG1IFs+RJU+X
Y+WTi7R+kaeKx5kBaDXw/JgO/TrlHJ/EZfVG7w5udB53BnyufEpv7++5VBMEI2v6E/wtUc7cr4DK
HWgu44ws1Wfe3/hGXhwwu6ZW/oJKbjNk4ko54AHaVKmNjoYAbUQS1ssO9BzbaLBwU98d5+pWVUZf
NbYosyRqMp2CHdo10qjPrx0pQ5VmSlAtvglBicc8mDZfjIDENu40JMDVCDIda0pzcbFshe/hdhAP
vATOkjh69eW3c0/ivMPnxrUEprGwhh/NlCRofok2Qcc4POMbRANiATM3s71f4Q/lk21jRvDF5wZ+
dwl3o+VhXpvz/5ThoOh+24IAO5xu6RfaZ0TPrfOwTjt5wMXhn05GYsJdan4N/ZeyLKWrU20OY4I4
UjJXyLpwriiFN8S78r5R1iBf0v2LudJNxCZ2r3g20Zus0MIA49+XGZbFCbGf0Qvl5ZlDIiiyW1Ar
3bdOzxpRqJNB9iv9xXIbSHFkLAbzAENZF0UWuUKxA6mVMW9NDX4oRAE1fjzalNd3I5FKaTWZLaWq
Sr817Oh24Yd5T326G+yfEHz0t71zyHDv2mYAkUI8tM8caMZd3V+5Gtg4W2hFpRbTqV01JqKbgWlv
WVZcJkidDP1CQA6+b6AIAcq6GdUNfu4twAJCtEry7E05owru+h9lBXjRUuNRTk6/GrOKbIGCzDXH
lcwYeUqzen9LO8bLx6Lj1DJ3Nz+d79p4fRyROL8cP6J2g0mKCzbo3CjvrM6/npuZvXANPwvtaGnJ
yAN/AvDIXk74MvB1HVE5prY7FqEz4G1ukwjWbAdu8eKcsCMBvk4dRtic+fqOWfQwRElJPPVY9wmu
vbCU0CO3dkth6RTNAtsfziFgphZlLQW7tDRUb9b1YxEgGnArzM+w1Wgx9cR2ZjOS2UCpGaHidrF0
zn6ojuuUunFa5CObezULMS7IHa4cL4MpgvVm2l1YzEygOIimYs+f07AmozPUtg+JVL+NeEtsgmf1
mDcRvBClt3+iZDpeEOB9MEWdVoKPkW5raINX6yavA0euwRbmg5+5oMc0Aq6JNAdlya5ApfMP+5AS
mLHf7euK39tpSS6ps+Z/c5yNZspho/Rf/91fbJCgUVOdczl8cOpTa5ij78KxNExdJY4lIR6ulxo8
/lS6q3qG2FUSyDDHoDFQMvNBnBVC1EdFULjQRCu5m1Bof8rVGU0GGkJOgI+z+CBGjMQ2vSx0Uo00
9ii9SHHxR2HOd2bEOx4HF49WzPiX7sp76yQHziH5xZ4lFolhVRlE5BdHvDZyhZEncG2Q6o0cC5Aj
WOGGyXsUiknETyu6eK7DuN3mAedCqeA+4Qgz02P/Slxn6Ds9xjvjZh3f+iKlXw7VckrIar20GfPQ
aXEoB0ZwiAM5fP8VfWWX9/8qQ/zVmiRdYLHnu+BOyRdR3JTFwmjV7k7mVSbM6FatO6xW/gMvEGqc
+gWLiqXQC+c/EVtn9N6fFz4CKSaaeOQ59XKRnfgIbI9amuRnrGoxwEob5HXILUbzEVmcI+lfhCpN
/j9Nk32HioHL3bY3hv3L+ZbJUlJUKIm3kOlVpAqoI5AnJl7r7KfForX87nuK2waASszKOPYErK1r
tRtTauIUG3zDg4tM+sOZ0f1yQbYbEl86Vw7S78LsmoQW58fB7TP2kCJiE0Rr8PSCtuzl/zDo9gTH
Kh15TdtM4bi7OKYaTv91N05XeBcHwsrVGIhWQjAQfPEyC9PjXAgKtNY9ZYHXqDB6+pzw66XrADyB
e14lHVHAeaBN7YlyQBlZ5fTrww4LT/s6ZEW/h2cmMTYqGpn5L81FUywW6OmbAd+61iCSz6oxOkv8
S/wdvUXKlJ0RvRddQ/EJyFdXNJucdSSrax+Y2VlfWR+kDHG0TwJVbz0eQlw4iljCzTRzYZjpoo0V
PRL7IsyaJFQVW5XtoegqEa8f237RnzYibsefNGMlglQxxdc2Ip1huySFR4n3gPUmcvgoQ+YbqP6K
piDwGl8F+/QwY4DtKPkikKxXXxaFp93NzRPO5i9ka8+AUo/lLhXhZkc5Hk/hfn+6hpoAVJEI07HF
obAdwVVYb82eE/MtYy2J4VSB8F5AO4KterNR1oyQYJ+3MUS1UrTmEkDOiHpWGllY+AvDnzcmic7N
Q1l2HuQUoFoI7UydOCsMQKdHVXR0O5wcleStCO5jIBMCOLKzxGmI/OtOAzbEbERC07Q7WXkHTHe9
VLhq2a72tMNDdzqeb7njdaovmRucjvLLJTUrOK+NZ2rDq4+mwiQWaPsQqJnLX+0dQy6DVwBDCnTw
N/OCuY7iFEIxFifKIMgGum3mEM3ttuyw/ptRwBs+Xd/wGmAjC17Sdryox/TkcegJ/TCqSZaZuWRT
1EkOvQ8fO9VjL+ePoel29+5PqdNUc1KaX1F/9m+ysCNAargqSOTto83V8UOIR/urLz5aHw6+kK3K
PqggT2Ha1pPXC2a7+gPydGnp4fN6RqYU8iyhtpG3+NL7VD087UCX4lnepYnIsrcO86yVeD16iFtQ
8sexJspUZXALkG/1jzzRMBJppLmeyeSKAkv/Dizfwa5pzcQGPQogpb2pFDuUOfRp3rzbPK0ZeRGJ
6nNZtpofek2CHtWFu1GoK3X/QUEAoSfz1ufROD+PHfGr3r3qckClovyrC9Vfi8uOQhdXnUBBlopj
69WfyNOQ7swT8mTj8iNjeDG1OeMksTZNWHcRKzg0wW+HIN1BjivCRLszZyMx1cF3t9d8ly6Qh1Bw
NtjpQbvUdp2CrArzs6A2DrIKDR4B6CSz0eIDrp0mpHn02haOKMnUSlQ5xzAwbE/9EKedvENUUGnL
z4GT8Jawmjfq3o2gNcuETq7Vt5rCFURLJY89/nVH15D/m9S32u2LK2krVb8p6lxTI55ZK/HvkJAT
qg5VS68qkWCiWf7fnKN/SFMEyPKHyHQt128xQh6sbSWpcPfQpDgplyNo3V7kyywnHZKrFUZZP8Os
DntPAM1Ja1m932vhD/VctOhgXp6yQvPWAqdbjXGbRiY8aedpRGr/940095/P47al6VK6IX49qUnl
YBZywKowvGVGgiORMu9XxlstpH2QDfIXsp/FuzXrB+6B3XJOHdaxHdBsXsrWLmK+/0DfntPhFEmf
VA9vpdlUQvpm4DiiYerTqJeqXTsaiWdHM7RHbeKIXTMQQJgXcT7i0f/tIXcXWxz2hVfKQcXCSaol
8wapcruov2+wRTzHldibLTjzo6/qQ7vFmIfD5UAnz0csRmVILKrovsvXYM3n0XH1bktahksqAWdL
DVwhEav8hZ8GBTN4+rCHhofaQGqkqRhc+Vdy3OrYZvJk533rb6unJ77E3SX1JoJYaYA0ouUO0qyP
77JwS62ppFU4DivOjYiRO0tPIv4V/tAZ+yU0N/jmfWWJePrs/0YFnWouc/QdeepEHV0pmW/WUvOE
tjaafeSBvzkE0BiLAYfJQig+ZaQQ3ECdCuKs/0LHSJTy49+utEamKg5lBhtjYFpwxUst77tTfBZH
4c8DrxhXaMZoz8ursy1eDtGuoIMDbTIM4XcZl3mZ2DCM9GP0flFhPbLJWodYlPYBWHUYzIsFV9iq
kAVPVTQ10F1BHbaickYgZoEqNHi76W7x80NdQQo/zE+8vbYDNeaSFHRV+X+zwhlKhM06IYViwBZg
aDCWlVllvZ1GZbvlJCq8Sx47CkEd/WV7F6axGOQXHjy1hNdPQjkeDfXi1ZfGUjQ3mjunymZ1SD7O
g2guuhCZwm+MfGflOEmkiSo/t0H3voE6wtb5ExQke7Dzq+m+rUM9zcEzEa5xf5vk4F/QzO5YZIpL
4OtidXsvieoeeiidBhoFpDSaokU0tr0xmkLYDc/IzrNtWMH9n3WXW/Bb3F5TKO9E1c62nbzTE+CH
oPuke7eKxOuiX/6pdqBOAJ3hO/7bx/xsyrRHFuf6cPabxlp1kQSDB34/Kn1tO+OptCMXiYzIiDYr
nrv902T2KEp202sWZsw0mNRK4OAfbQVvsFDCuAbGrt71+n5V1aN3dS4fvVjmXXKsxIJppdSXs7e1
X1jc8v3JWe5zPrwmz3ipvFFH3kAFmY8Bnqp+ZnahXJHEeQH3Rb0tTKVst/S2obvjo3POIDC6UZ1r
6N+vlUikDZ3AXgbR0p00wyL10k57Z/g5IMGmdu3xO1RCoBUDrW6Ynyot/Ovdpp7Udh8g6KQ/tRL2
9egCjJE2xUR30BlZyN/aGEuVACIAn4z+xUt/dnFw7c6tayPctcL9nXWu/ujFhkPhNftf1BA9TGa/
xZv9m4QKPD9vtbzny+L+hXeoprtK6VZY4FK5F5w/mP0pfKOeWu5uRomqx0TjKlGNLnhMYz3Fo2LK
UHa2v4Iz5rYyUVU0cgeM0k3c7vDHIZF647C3PBCxjQJRKUjm5R1v9kYo+KBVlBW5wZp0i2rwG6dv
/ZAUgoHLMvCxuLdhwd4cMaDej8oA+nFiPGXBqP347C3T64GaKfeEhcTuYK9z7MvD4xL0ZjghRlx8
6tE3PJNr5JUudGRGUAtYq+NA+9fJ32PZUyz5tMVDpBIG30UISuLXiqQsvfAE16x6TDz/aqWYbi/H
k+Qy9R5xLiMrEj/gDJ4wGQLXFYxt3IMEkU7fqXILwpPAiAP57I/oBTidQAdAt6gCLzsnw/0LLrkl
/27I8AFYX3vWQPJo3PyHejlbjv5cHed7MxHXqbwUim2JZuVTSs9imqPMvG6s2ti60kjhCCWN5A01
XPR8PCO1+8e257GrDZZ+GJPmAVw5S5zRRgpc9RhxP9v0JiIWwRwAay4Oekd2iX2PGYwR5OMKYgu5
d7YspxJH/6IvBWTyOfm0p6ory6lsrP7y8SRzp20zOiF+6kcb2jLSgmPWytLg74MWbdu/fxBJWy+V
S1RNgoU7viXEHQbnMxp2uVmBoXEHNeyzqDKoNYxqpfpM13d66+w/TiMcSbDlUb9IHgq9o/QuBF02
nGUlrs3Fe2WMwai32RtzdsoJaO2e3ISSJlK2yqMKzgJ63yOdO1H+ER8oZJyfPiZjJTfElgbhIDWT
4LytOzkEJhQy+UlM9J8lLTxW2Z3uU2sJH/FvqJVVBtEl9E3VVSpDt9+4nI99gIN7ihlM35UcoG98
8a8fpV69C1hJIUvEaAyHOL1xW45TSuwRXoDdQoTL2lhPP5CxZ02CKXhdLk7WmWVaiY7/gG/zvIjf
wG1G/zVKE5Tg6usyviYcgE1CQApSLwgVr1H34OSTclKhkXLla8+d33d4isMlEEDqocvxb/X5WCES
4QWOJmjjSFCjxgY6K9iqdWQDix72W3nh/BGwlEnWVKR0nXINLgimvOpxv6IKphBAtxwxZC6QnnMV
WAXxxiWDguvAn3DnmXai7ShZ7O0PDgCOOYatm+tcVANwlzUYbAlnwj6szI4LrhoqBmxogPYwP3B9
q1S6BcVRO96J8eLfC6eAttD17kaTrIEsYY2BkpX5Go1krVs9Arom+Dti5+EQi2A62Sbau7WAi5ZI
AKdSuWn55xQtXoCOTFySEDLo5qY6U/UmYpT7V8V3O0ITORwNOcnfj0zdPytcvHqvNqVsbM4U+Y7e
4C648N7E2pLaSP3osGafqA5xYek+vM+ubvVYLxpOg0gFtOgkgUDWhVZp8ARswng32vzY96kaM+he
1SUPhFROwWUOamsX87324oDijJc7G/JCj0JBsId36NZ3ebgEx3nBxttEryXz4e/kEno1OYRVy6pk
5dV88UeUCZolJD6FpZ7rKH3BJGxRFtaHkReEOhs4ww9n444N/9BekkZg1xeyoTZXstMI/kFfV7Cc
JIjBX1Wg9CWZVTUajGXO3MMJmewHfIaFaU82XYcuLe5/cDF7Vw6Js+uNWNHnR7OWvy69HmBoETq+
3k+lTUZYwkE9MWwWZ89PZUQ44W16oBTgu+u12cOyGYPgNLFhvUeABxDNm4q0V7QTan/qfXxoadLT
Yhftd01wB2Alc9KdJtQ4451DV5of0q5HkLLMZnOQxe6vhvBVtl4f3zha9n8VmyMMkPRuGxUxopMd
lKEqkNZMPU7WWs8kqRI3Dlszq/73siOBBkVvazjRaHBQ/D+3nFqI1HBwDxTzTGcOh8EDwFTlgT4/
9ra61jGQ7CDF0MTMD2yan054OPb5WIgURpksRdyw0QkC1YloK/peV2O9iDwqEAVV/gz8xEXB2PzD
fhiNzq9tBe3DgVQ5ysnrqMsWWxPcPAejCeJQHfYDDi80Rsb+74ImKt1cgm7kK4cnfasagqbz7e8p
fonNIFJD0xjnT1gQ45zOPkrDGeDR5A4v59guobOGGQt3/1wzZiBUfYLU8pTtAaHyM9VkXf4pHyIu
2vkLpYRqj+Pnwa6BO2d7RAAqttNx/+fDSLB7G7k2zF7dMY+gCSiCs4/Oz05ZX0LpQxLU+b1JAdc7
g6y+oladvws/TEldQupJ250DnHKQiOGmPhg7BaDyA9sTfFOVNeg+UmMxGPsaZBHMmaNf7TNYpyPO
JS4FTnJVlpgXOmKI22be6SrEAq75UKT6kOnqAtSIBSU+Q+KCyuv8K0BPqQhdpiZ6H43Rk7gjmJnI
dRO6ob+xmc+FyoHzQkQn/kSC3BIgbSm8s+dcx+xykvwBRdq7yP+utREOVb/OAVJBVFMoCI+uIbS1
squxVeK3ppO0Kyqmscy6m3W3xFaL/lnInx3NfqvglZGndfQNYdFWlNE9iV/rvnViblh6KeUg4tcl
5KxC5zag4WTifM5GzDdlI4r8CaFXcAjVegkFy4HwRThzBdIfx90vUzrQV72CKLRI/R6VXNPlj+cd
8ksANLv6PVpcp4PsOmxMLmdiyZR1hxTtlEMEmXRyJWt4OeKyIh9WOCzincFtvQLs11iyQrR37nIs
skIYoWgSrBnbHOVCohNVQ1TRdbfGlaE2jOex9mRn39MLNdl2QZjgerW1O4X5LdlZYdczu7JMubfX
D+D/HTEKvTSpJZyLhIArDbxjHvRoWvVe0SbMc08qU8RK1z9WEdZWUFtgH2EIyh6c4aPIUoaVNrt0
7BkyZ06cVIlTU7kcb3HjwCVA6tH8JTUkzRbhYp9/XurbwEebA3lxCSUvzOS756jKELA1l9+BtmLd
1GOUeeRqw5rlCKAbKVcGUsXbZkqpuI7g0wg73jXMcZPQ8riCrF4xMRNqhbCI15pP9P2GmotyehD0
Pg8xWoezDQzZ1qIvaX6Q/jUsPNV1oBKyS+UaqIZawK9TPymahI1Ib79snptG8w9OrUlQb29AOYPu
G1xdxk61B3VfDOUc0+xN8of5AdXMzkM2q+P6KZFQCxt1kyZa00d4CrZqT7WQxUyLn+e1XJyju7rr
HxGzOtt0RbTdrNdK0rNtIen+N+iTyKv8IP8Up6uADJQEk9AWnInVktq3GRXmDkD1s3egAGXoeyr+
4rmnufZVDCSpLVUk1wNfAzcqfFPz28WbStOPbvNtUTId7cDr97bh/uMNLAqpZrhR1mUcJJOOigW9
Uzr+O8q8Lq4/rfcm7eVMdNrJhbnuJ/MzO6jYIlFfUeQzOfGZdd+JDvM+kM91R1zBB+TXDuGRm4xZ
XjxP7CNDXmv+ayJYZe1L7sM4fhKmG1M937swB+miRbAETtopelVulLa7CmOp3PeFWoElg4kEcs4V
ouH+mnAKOATHz578hMPnvpuMzQIMrXXhhQEUMH6dqVGOzxNvG1KxAii+bUbxsJeb39eEoeaN1YuW
U7+J+ARpz2DM38K1gXM8j4XCeRuiJ/7sXOOs1lOo2GMStwkwjS9ufLRt3s9J8fimVjXS3DkogmDB
KtSDHZLQ7g9/w8Hra0JZjzXBInCa6bnNpdmdTOfnKkMxj+15qq3eS6FcM9/HIGkr/+UuieLtHqCe
30e+deWIGfXxUrP7UrVWk18rmXODRhM2mkRO6ZULECOMvj7ry2FTKg1qBSepHItcUQOrx7mUwMo7
SSljdKfRsRxbRqUasllbbwajoXwGAV6t25TPRxCXqAs3ZY6yGSHpV9/1NDJCfjp6ZH1PokSmUBPu
IuasF327I3wWeWLlWJLPCVlHGhliLB+KrqJE9M0jHtFkovJQ2pIyghGzgfoB36OD9s5gLBYiJjIb
gbGv+LwswvhlSQ9VTyBEZC8k5anewRVhRNpL6Bg5I5yuFqeIX6j/xIcKCFVd+C4apw8y0LyCyL5s
5RWExRmfQjj2hGGhCrplxpTh9VuE9W0HqasPQJYTtl53z/EdTjJPRXDnOjzxkVumczqW8o5DNcgQ
z+YH5lmDebLATnW3smjq6HS71iiH+OkcNXLBk3M7K1A4XGz+4UeWCGxq8cmbrQELpBHWuDN7fIzL
cIkHksmcMT3Y1TtSbRYEnXm8/CB8hF7c+b9PKNq5n3tmBl264eCfO+uqKUNpUYPZAIlXcNkEb3ol
k4PUEvx/qGBcI7x0/81n06Me4eJxN/EublH5ALKLJyibaVkF2jS/NdwSepYJRdU+Xjg4SQFTvQee
p8FnBUk1tLg3l7LT68vUWwCUdZpDHuc24XR47FidFWFvhL24ACsj44WNs5dLR7grVvtgvohbe3tz
2YkiHStH9hKqhd2yHiUyQi2qCevp9N0YV02WfqdoX7YcRa29tBEjmOM5PLayEiQbtz/Pqgzkjz/x
u//UubE+60sLI3Chvg8fAU77ja8gNqpAD7qf8rTgN9GLkbhu1fPRkCi21fAyfzjLhvNZ+9Xpl9uB
H3hjgCKicU0vanO2hJLLWGcjUUPNhefEdCSnN1AqjBbmuJviWZaJ2lLxTxlY1vi4zqMqf7qOcvyQ
yMlD0DuJCcXBLv5abz4iWms6hdGsepLZRBhm85uTjREM5kgU3SaiAaE878+QU0v23DgyaFq4/6ek
3wJtLhknSJKe353GQtulEkL3+nyQP1qrmzdjAGtu7bnq1t0cQ/PuFJr7OLPgckKRnCTJSeBPnTgl
z1K1gQlvBxuCGgO2zzDlSETFN3yUXgK9YKSvi4JnwaEIns8wST4fmkmqgPvD/fjQqdSzAKaS6jH8
TKGFY/YxpfXW1Utd/s634yzllIPCpAUdoQmeo0CTcfrYOhrxhOhC/MeSZxtnrJDFK+NzTdzmzfDp
K0Cbnt0X58R1B+NFRKO4KQ5Li+IDgzySjtgtDs3c54UrTRw0YEkn0ZgfSzWNVA7T8aO7nOn+RfeN
9bNEiXSWLmn5oEFncE9z8D5X5AA94SHCPxA+Lhoa8FdeO9+oi4Jv4JNNFf0zH7w0ZC1MiD+QcLEh
+LBw6en6EseWcp+PDEJdgUH8JGrceOKUOyUoodSyiZ0zoWM8CR1H4L70smoYm9Bahba9kzFAjnuk
G3kOYl1DABU4T7Qm6B5T/VD8gj0jL07+3HhLtWosHOGuq/j3FTrko+FhsvKqaGTVGYPrnlXtSJUK
Kfg50krsrX87kIa09COpDaZ4o89OEvblO/jaAuu4YkERcM0OhkEZyDvyjL4dVEX74+5TG5ZJW2mG
3lKPe4G7rpixZgJhFcaE9F2MOu4mR9UMWm+j+feVR4CxZLZbzEmnqpr7SDF81080U5DTxIMO0bBF
ssYE6GXU5cA86YrtoZF9nWONk4QTXpcGK4fLAtgmPaZjedc0y5NeDS6vkeAFLSWREdyNRH02V/ig
DjhzkuBPgNf4VB1LLz7NeE3/NUBJd1pUmT4181siBDuA7qlDGe4lCNslDMBC+G0Z0pQUcqi5Bllj
7Zgny6Zd+mFgqdT+T3s0DBDvSv6keJLL6qB4ukcEOqaBMECLmh/8HkbG4hqfxVmuGctXvN0si+Us
QerOwYw19iMBww/bSmlDey2FUbbVYPrKrVMNKDHv9xqEAsQjvVq3xd5nv0WYafyXju2244siX/5W
xB0QXa34y89MPQ55xC3ylHBY4ygDL96EzPEKs+kxbcnxTqSgp/Rr902d9a8AKTPbcktrAm0dSJ+q
e2ymqm9DZekVK3NjqmJZjmGHn5KV8e+gwiUZqYvb500DeUWQCKH9ka6yxWBBEEAbdUeQfnRdX5oi
aqud8u+CThSiIHqNcLXglhW5LJnlZwoI1m3joOy8VgXzIDEzeRB5Z6Y2NME0thkZiMZ7eoiq8ZeF
0HE1zejs31jYvTw5jtmI33iyutQL15AHhvZEuWxQfgNFTgAUCEoEQp9g0OO1EibHSGDKMA4Pw6b8
O9ap9SfrlBf+whTqLVqQ2gLAUAkfM8LMSR8hgwEjoCl7L7aybLeu417SsAX4ZqYsYk1TwwDvcwAW
aEKmy/6Qvmt8ob5qoS6jY2DLnVWUs5a3G9b2eagR/5XOXqvPCEmilcLHQ9xTOOuLoMlsa+9HmlzJ
+FURRSPDPl0SAfEHdQA90KOWX/+gEyDER8SQH5D0ZMho6Z3OCOojCcpKLKKoYQg+25Hl68Fkk6Z0
AB9ug1d1KtfXgW4a4EeExkc7Sd6SxKhlU/iB9X2ZAiuMDU5Glx7sQ/Cr0H50FOnKjl72tBJvrrD2
b+CvNFOLVIhYVNuLnDO1etO0DKTuN7seJM+VpOUfxDcF9Fk549TDyeYU3Tw7Sj+hY7vvSdDjeOxp
B7uVbcJZaOQ0AbrW4CMUA45xVqjh3wrBZdd30i6TcZobMuaBXb1q9x98SDcHgsiyIrjlyY6sQnIT
ksZ/aSGn3myKB4KHyaXtrUBU2xe/HXTUob21DNHbmXN4JfUizScE/a1B6qmcjEwC6Z7YisD5z1dJ
bCLoEnwkHtcbf7NDslzuu21KcZ8zP/sPOwhxe5IWYtOLAZmw0LRfA2lh7PcF0yIy6mpHSgZILQQj
s6mAkWWYicxdsyKDzO7hmhTDETvqcRCLFEwDH3paiLiRgvXOM1fgirH38xcQzajq3z8v15g5Ty1r
kDaBUOQvVYtqVfoG57IXP1gtru2mHAk+HQSd/PpINIXqdCu7G7DCKS5gVjkBbC+On+ZdQCASWxLR
w4h2x8AIJdX7GRixeJWHuljOBKfM5U93vgKAzHByh62iD+UBdvrpqIWRUSrtpwO3FsbB942KXjxf
t/Ajl/wHvVx7E5Ys0hy8BxCCEE2HQAScwSx6R/2XFhknptLXeI6Z8+ka4wyxOFbmvyXv0gWjYTVm
+6dXDMZW/13izLpNndkkIwVEv2VmJ6MqNlQDv1aPqqyowhBBW+A6pSi0+9UJRBuwEKrlj2PvoLq0
EJT9UhTREVe873vDofNIqErcaSMI1vib/xR3xOCqeqP18GqNJUFf/yxDaxqK5p9R2CUhp1hgpVz+
YaQoxRBaK3Sx4IPAT5PKiLdmTCZmnAwsnXHMMcvI8CCD6Aoy71/LtbiA5AcY4ZxEw/1BeWw+gpAu
Jy1jIKSf/ecCs+MNvhowolPoCpg6FP49q7j+a5SK0iv0THA6JCD5ofmUR0K5/rU/VSXjGxS3sHJW
KV+Sky5HIYcZBmq+wSVbm8xEesV/bgwRQyYCVvScrXpKLHUF7Gh2A425zNxxeVQYOAR9Qf8xfPPT
GRFpW6NfzElCuevPAUaUpsfJnYkFGyiMYhqMau1A+XEaS9jdHZ3IxvPydXyoihiF0RzMrGEH9jQ8
PIQ07FaiJMUSxBrMx2n1W1Ktm8OiFm5nm2LLbBC5RR0o4zRtJGRGciCdGv/wFz6E2F7ogIvpvRh4
7hkm8JtoU+PQwrdcrFIcN65LbDnz2IIM+pzwO3/n1Kp10b9trYRvjrI9m86Cihd+V37Oc048S6LP
+BN9kmJiB6a6yF+8hH5s8wy4jBOOTM26CMgeAOTZUwGQLCTut5v1plhNxRAlfSSbGpzUuxoo2qMz
cdbbyxvXE0phtyptT+VxDszpKhy9zBptUEjwOJG9VX14x3yZgVEeiU81OX37A/y5FI9TKeAw5c/k
LzFmeFsrhUYTUMPq8EB62XAL2/srHQyNMP1+V14RJZoYApqMAm0PbA6I+qzdaHV8PSZaAZAUMhPS
bGN+YfWamoz/0sRCKX04MFR1PrsCgGUeEFILLLeF83eXJ7VvBAO//gakfBvOaMlSdMSngmgrVLwP
P3HuabRXzVIbVGGlSY0BlQDNohUy02lEbVZYks8mQvrS/NBB+sFFKl29Ij9xBNbiFYe1BIywO6To
8wpiZtI4qOL0UcFWCkEcGZOZe+rD7XLnzOR6h6zzcCKLaRLNf9Y9bGLcU6acnQdUJKpevbNWKjFO
3ORTQnG4rsJrd8E7KP5c83RSTpfZx2ktmmr4LYfLkUQZ/HKNKX7UoUpzSDHAv8AdF5OgWnywGTT1
lZR2CkQ+pP5Ep1ICGXvYxB+bAaJfj1rC5/4OMlmxorlv0+2mpujtXTmv6aJCneVRG2L1BJBXc1/N
Uxp4tmXST0ADkIyINNTM626pWTDhPeGoEcbeFrt5WgTvbS0yTUKI4m+zKUAEkG059coCJygzm9wO
nwSiJbvJsLL/03D5a3tvZUwX3atW3PA71kPgmqIzaeH2Jwaic77rQ6lHlq9xnyvge//DTjkmQEp4
wR+781Ql7KdY1cVoKuZoaf84QzKesafCgjVoHxCmOkASS8QJNmlyN3MmoNJSeuMVYszRJQtXqoA2
ZOwIfMrvOpx5+ipeCkVFrgIPv/TEzFDOAJjDVOx8M6Lo912RljXrC1IKGjA5OESpai2UtZSey1tk
iPA/OKMaw+KSzk9tS0Y0Hn/dkZwBbULNl1QTRVSq4r62kCwU6TFopwbrJokv7SJjJsfmroQplt+a
x8Pm1F7Cl7xONlcbJAAvgHrTn82ZmTCEmXzoANGBcNgZ2c0n3Gh3unrf5yyNwXREJt7K/TtuVa3F
oL2/dhXDylW+0ERPq0HlBYi3EaF0/c7anCfhi4PcluEbqZS0Fp0WBraNYpEoGc9yqDiaVa3LVAZe
VJ2CNufrJnbwwMhHuCu07njwIyTXuI51BsMfVe5viGTdIHDNo2Nk9ZrO5F6+c14NHV+OA9gKfMA2
GhDV+WPhp9R3s03gRfDcN+8MVlp3vzzCHue/mqQIkxIo1AEAdUiexm4oArtx0CEOTmfoO55Csvs7
ZTmGZf6XsfsFlXDlVdno3v1DD+dZsp8kjZUXLutq1XWkimUxfGm5jrwOdSos0/mxiVBvwjHCI+uR
gDee7nSBHKqIhPQO2ZT4jrdr0sXLC2ZNvfMMujaZ6StX0k9xGuyEtEXnG5pa8dtdBeukT9dI8Gjo
pEFXER35Nz++4Hw8y6wSHFJInpyj2re+038EzLyy3lW+Jc/Z9E5SI0Rr/VVfCkUtcbBAcr5uA92l
8wNbz37E0Zykv0pWnN30x3uefZadN3LrBlCujama8CmCkRnOfsGkuBaX/WVlpc4A4hVw6k8s1Ho9
fpI4FZ1bUzXuRLE1EU7m/Py/Aox8eEqzn4MBwDqTKLeTWDQC34//gfgSIAQD1ZK5oS3Rq3a2SArl
p+PuPnaWpr6/GSGq+P9wigUZQEcNTl3OO8EDyk2pGyp0KgYPJ+wS+A8seTLxo4qycR8L2F/wJ4jl
1sUAwgI3yQ6u58p/Aw2s1mCpWEhRSMzUIBeeibje5iNwlO6gQeal2/iFA5eOXA29I/74wOIk4Fae
GDNDbDUoIw6hqGjYmaKuF+Bik4qedoG6/AaZWxcNbZYCNne23hE09jjJ88E0OYA75/oVe3XBMrSO
BLCQURspcv0dzt1jRnw2o3c66rPmX7ZJBTgf6upEOvam3YrQKWwyvX0JUEbL/imXDSsGdpC+gJLO
2dmtb/gfQF7I5n7WUCdXKkwRhrLOHiAVkzM8RESMqaAuQNdCUKJYI0ojDBdL/SgudmDj+qLhehVu
ek6mlPCi5Z/b6eOXorA9c3k8m+uvf85/LVRyV7SZZug8HSvrC7B6KUs+HWzzlx3YYrOyu/+SSOtF
SdEkzseddhcaQRXP1MSDXDw7Mhe/9Z2c3OZYi/a0ffoIh84itVfKmBSP9n9qmXniFB8ZE/0fEQQd
+sF1fDul+GR8AAgJjNVzGt8IApCLawVNE6Xl260qhN0gsu/LXICR6FSGO++K/9cTrty5mJPyUXod
rWG27L3yxIQVUxcHs5m4nxPJiOcJx6jzjyb3QHALI3rGZ0cw51JZrh6mV/P4GjW/rjbB+UN4/vn5
KAKVBOA57CJPyaVF/i7TWLc6loNC76LBAWRn3Oton1GQa8kNPPMkLjXFP7oY85C3U1LhqMk3r2+0
z8evZb8oR+5GrLJFsgQIOwvRvfB7YnwEDnJGzMDo5y7G3Glv03SJoLp5Mj0x3CTmRg0gfZjKWYM5
izy6ORze2Udu43zR7yDpg0cNLxg8vptOrgJ4mPiwDcwGr9PA2HsIVjJGIzscdU+70YB2GDeoFcXC
Y6RJ8Bw5BOAbKmsnhCUmIJVbNLdp3njvuAHSx1dPjI/xcFBjFYdjSbZA8Q8GPzFqenk9ijFAt1O8
t9pWQa4pCsr/vytXIq+l0juaOPEMQTfoL73EDIGmBAekk3SDNpVKL65gAiqVQUPWfipNS6aGrOZF
pO/YB4F5Ae6ezIM9feDJkpJrQEp7JGbKLRlNXa/3HAh6VjiEJ3yFTRkMWCnvNVCIHpB/JlpspX0y
7jG9CxvFk4A+RKGew1MEb82YS2x5jClqKJu5uR9v7q2jP98PT/Nm+bYfLBxOajZgwM0Cf+IBR5ia
d8u8jniYnK5Xx9rbmeH99Ri1pEicVPiwztNgdtC9Un6XTRjRKfdnWLKhpUOsLEqCJf5SE/O7F+Nq
kAm7AvgcFiDwXnycjYi3VNecHKTdcQC42I4pquE/jK4/ZHuFL0dRICXoWGrtOKRlqCMJM65S/N98
ErDXsyLSAxXwtny7q1YrMaGadsAoLxAu8fBHUY9ZgDEkfox3tqJX889HxHKNquGpblPFD6ZJgdf0
6WwOHvbyU89nF3nXKwv2gSYEFHCByh6yoV3upzftt6nqlVX8+jNxS8GIBaGoYfdCnOIjfBthlrqr
QBuK5eptjJysrPNu0jU9IlENxJjZT0oMBfHLCKcLOEn+3DcpND4Y668jTLdP6DBkINy36HlE48TC
tomhiFi8zwphThZRt+MPH5r+TwYL3VLJQ0P0J8vkGma30w9Sdz4tKMRaQKUDOM+Vyf9RtOCIUedq
pv0WDy9+rrr5oLJzQU6oVexedYcyR//n7lIsWhiuzUpIVZCirYIDH+1qlYHgIIFQIvYmMz5+c2N6
mJlpWtIM55LwwF7x5F9xI9v6W+Uv9nF1HfedbGsJrO/7OmsBbRq+f4p61FR504Erp1LPYyS/NLhS
8YE6Ta949K7HPrsVWakuodssdn1CnpEyfKQbzs0eXOyMX+ql40cjmOuO1Qpw9RNx4N03TXze3GN4
VyOau4j/GKrBYoUhS/WOgX8MkCGRbxFHsWWL2Kz7u7h6qNrO4bKXXNjPhZQewER2abmks2ObNVmv
i23rftcz0hMbYbzQzOhOMAlUpPnUM2IIphnOkXxdoGHpeOW2Gv5B7moXntJG0Pga9qBq1aXZXh36
3CnEfQDXPJ0ARy8DKP8KxRRo+IdVlqGlPmWOjAT9JWS8dhEHv0YDmf+Mikmf9gCX6xHRPl7P4gL0
Wcokz0uBXvzN0mvuINWUmr7ioMV2Ea7TMJJ//ZSpOfQGJ/s6s9NeysKis0FsVeWcdr3ft1uR2yOW
aRQukBsEignQS7u28wRS2cYKsVUnPCALSh/cFmN5a9xd5g1jFjX64BVznF3kJmZwFuwzIfcP9KxK
ra7tOJSrBGM5ZGDvebrFKdY7949NjJDmb4hf3++PmJGO/6Gtb4H75scCMgW5jFJc0iYB8fXPDkCP
LWBpb7/SVlSPL60QaAuXfT2OAg/4UWHKu9UMo6jPgmqzd9hk+fwMfA35YPjdw0SVrGkbJUbgpU32
fgu0J/tjmOHeLmrDPdGGiTzlW/QDsEhjs0n8+omxCns6o820/66wm9bYeYc3utWv99rzk19Comg6
eROZ51hZggWwDx8aAJf3KLLTvG+REMcXLxhn7FjaMxCSZ0kxX4sjrkjNxTQYn0PYelXwEg8HqkXZ
OJ4opzcTmNqH5cRrbM29pfouU0kbpvSygxCRd82RJ9Sj77hoofzQi/XyJfvVUq7kx2CucdQgDMRO
e2CIJ4Oqq40Dk0bxDo0D0RX8JGJC+Bvjxhu01sTl1zrzfnkoHHItLB5BZ4ZJGcJwU+TEfk+qf7Iq
WWVwxP5fXVVR/z6EhVunl3fnSJfh/+pPv1/9XbvNhMN/WxbgwvK5y4Uts5C5JeAg7mKlKItT1uef
ila6tKIZHgp4gBDc8LcE+6m7jws+9wlqjZrFZ/9opIilCcAKKEh0DZQylPgiL40xTroJTabL1viA
1X/VFnfNlp7RdZeTGNjY3Xx77se3CksGXTf4KdWVMXHzQN8iWrSIbf/vceG3pL+SEcHMG/8lADKS
GqVTjIXxiBGyskmZHrET4FrrlLWvfq6Cj/mqlZTSaJag9JCIL0Gn7LiQEugVq8BJGO4rqY3AubbA
QfFlnA52DmMjglXjxOKYwVOweGK01CTWYaDBelvRSDmMybgXEI6SF4PkT/j3tmTk6C86L80EF93p
maFNhETI39slhqDwXnQD+NPJ8g3BYOXDnBxptYFQQaKS867KzZacWpIDzBR8Dh3va4hBuVHS5imd
wAp+6h/EXb2MQSfdN+q1nytcN3D9HoSweydt2DVuhQ7l2/YiDQSb3qg0dMbrASVm3EdHtuUE4mFr
fYVkc/3fF+hSBWfoBJQQr1qY6Eun7mBe41SkmjAk76yjKeHWSbfR2TMt1nN3XZxqv0PCjzGwlahF
m1IFNTNyvV1SrBF79aePF7XY8PKopEgFG0FuWMIkgfJ01LoYJKMK7ejWcGxEERaHHGM9ydJ5L71+
Y6ylqnj7y34Y2zgE9qr+h8me4QDtCayiSAoCh+tCXzqz+xQHjw0F6nczEaSe3iwineCC+NWQuLWT
t3x4rdTxBM5Ks05cjh1XqMnDJ+2kv/CK3qXH4dE6oeyabI7lESJ3Z1oeWhnaPeI2npH89Cu3eHxi
521jBBTOoIt+EMgxeW1qt/QT/pz4WR8+2HBSGjFCRw0m3yKAfIewZUHj2OdkY7fkt04Q9rNCLZQK
/DmBkCyKjbAbTj1Bmo4GL5eN159PWwLrcGJn5er4PM9lPqiliBp/P15noOmKUaeDUP7TiJR8Aych
BuPykLhx0QmdRw5VatJJuetPq0v0Uw84w3S/BAThsI2JCZQVbJnPXkKifWgTms+bUQCK3xAvgFug
Kot1zKIYkNv97vmwJEBCUCgaxEc83A9W5r4UtXEtg7pJX+ngi3KLEeCUl4SAopo/gapnsYgT9axi
zSNmXpKOWQOoPk1Cqyqqn6CM/gho6K22RCuLSLlZ7nqWHCaxjZlgZo4Klo1ggu/VEbw9o9u2Hwjs
79+Uc1c1mWXgTIZhwfdnq3WMN+3/TK/Qv7CQFOIN8HVeLmkAzbp2F2pIxajJo+LbshZhdUTqWUWT
7XzP0k3c4emCftMzgeu+4TM1ICnfhhBkXCSmY8YvkOlN0G5K8IRI8csOCy54YmWf6El1wO83DJEg
dJDYa3awVdHfUYi3LFZTOUM4axwd8TCPbQgAZiE2hXIHVM6YERDQKB+s51pB/Kq8D8AaJTSCKADQ
fDhuOYoXJbMiHFHbY/CuHMCKyz2DktxMYDqNZCVenNZrbetWvb16gWtuIX0v3MdXdnpJlnbiR1i7
QsOb1dCWqwylUxCU2vqOOmEWA93jnHDyObtox7dA4nl8rjHAzFaCXMfq0c6F1D3VeoGk6SXqTF9G
jItvhQGKtqxufGIwRqgmnrS6yLpQPRaSE1BeOfeNpPyGIafsaeXj7ibAyTcTVKXB8G1xb+qwSeGv
Fnd6WKyEro9yiJVUChsgWzKrSCqkEph4xJ28Ujn3AbqHjaMa6aaD2o00PJkKDVv4jJhwH0BqhAeB
Bk3mp3lo2giJPseq5e1YZZlwca8dVL5oF0yIShgUpj4LEpea+OCdadpSOuqtizMluz57PIipSS6b
cpPnqdgmRtG5dffgXeBcOp8IRuJRuNFgjGSAX2xD0uItDZeB87vYMj5wKXiQvFep/0N1fHhOmIlN
fN+wtjY7lvasesBooaHplvypqC2zhsQNmdXoemKbLZQTUYaL614NZaClfpHReiNtNocXJKE3J4nu
YiPKW+XrmWEkXfA0HljYxYCz5APYiovyRrR/gVbrGPGz5n1pZq7Wj+LiP+GifOCNG1BmhginnVyE
96YDZnMp8bkWa/R4kipQQV9hQFYvXbhXCm5kQDYHDhyL++2/BXZ13APkYKmOAshqbbGPy/G/Do/0
tZhSYxSF0xRWulGFNnmOxcbZcHxK9FNNEzWhDLquapY8kyQU54PFltfesBPWQIdDKfq/c6DlKeiJ
NyxWFSBI+KvNpJIHu3qA0Xkl0VighkTLwA3jtDIECNy1bHerU/zV9LSWipPSjzf4tK6/fBkrU4kI
0zbHnBgMsF/pb/rXMELZsa1UjwfdW7VgMYaK9fbLUbtUprUtm+3TdvkEpF6B6jVUQzmcpkLI6p+H
vOtNnFsyMwLmsPE3mcildZ5K914srtdxxC3sd968SDxgyLE4kw3nAs5QXtE8gQV24mAsQHSE1zFp
qwkj1D27ZEYyqNumonxZx15qYW2XjH8qlGNem7XBnjOIXvsLmh3hE7unWIc3wyVJd+icid1SbhHZ
cztmZG6Rf/5A+chZDmSv5754qAQ7vTbevmRO/lV2sNZc1+LyY953r2z+QYxBXcx11Dgkv+WToMbn
pJJ3c9aeFYb0oAkol273q5D4aQ1ayiQv42hu5elNKklRCWtja9ogn1iVLvxJ63iYiYMA4n4DKe02
cVr00LMh8K9RB0VYJ7Ni6enPL0B0hLSHOrdK4Pr3oKwIRE4E+2RDadBUKSLYMal/IAfelungPg1P
gbX6GuEII6vuLVVPWTfuTLvP3fLhkWN/ElJd1dQxzwmH+W+2+Lj/saPMzve9GmL1d35Utu9UzHy7
6ZEHhbhY0mFZ3uR99hDJdbUNneK9LYKufgtOudOIpMAD93pYaRQQu2AMUb/paw9EXWhHH6v5l6Ho
NctePOiW8iYMcc9L2pZGFkVXVYYvgwrkkDuRYhcJgEWwUdBGzfbHGmwq9FIkspDJrci8Zxp9PU6Q
o0siQ8wIjp+PYhbT/LElQTc4oAao1ryB2NvDS4E8Q0mV9noNvDtjjzPz13e785xEn7dZ+4IaU+8/
mpvrfUHv0PQO2mRisincM/LybDmINChk8STrMLXod/tYBg7IGIwuTRK1lSinl9dT2ObQEwjPL2R+
si/Ban26PyrnGoBfniclNkVyTcAtzmdOshlZFePMQNbdZhttl/Yz1Dr82qiVKtW//nepv0Q8Tie3
8NQ6fpGIahO4LHPUal9XRjSTsXCEPZcJtqBPZKo1tUzdOepMTSj6gg8noO25yXm88gUEVr6sek7+
47k7l1xzKim2n16GJcdzfdBs034CZx6k7AFlfKdUy0lHItnk8+1NNvLhN4LPhuK523nBX5Vme+dF
GneqE9sE4Bsy5SuWg+RD0iL1ZsgTWTOs21oxRXyIIIlMgCrQmjcz9NxVFC8RBiBQExbpFDmcZetg
E8s0qebsaHRYn0oehloa6iy58+WrWa97Vfb4SOrTZEgg0ITmwHR/vCekQbXR4mdjqQT0bnnNNq5k
AgwYiJAlgwmafTiV93hdyx9Q/PJeQHyF2ajeUJ93hW8YKAck8FhmeQ0ui1xZ1idTahyyl6BClx7U
ZoMY0+F+gT0KVJey0I1kqE7WfgCotbQ1RWBBnT11V94Cn+ZyWLgTG2dkvjJ2oWhKpjhBgARA20Yo
F4tddbWic2kLCYrDmMXMLdqyJymPlBY4jrik4yLRhjw+/NmOS15ejHXGW/NLku0BOFE9oB9gQmFi
SPeo++dIhH6+N3shAnqF8K5Gdj0L09pUiTbL1g3uJZxbKK5UF+P935EWVZYFLweiwGYK7nXlbXd1
CE3QaYXaEXOs1NWI7MjcY8sM0haAdeVgK7LsDEGiplQQp5B/t4lF3TARmPK4p6ayFy8SalvCO08E
dLLU/wiwJoOSfoy1bd+X/mERW2UWurHakVB6vvX8YvuB44ZXhhZ8u/weG1O/U8gBDBVEjPBsoD+O
Z5yMAvcA3HT4kyUflJCGURh3gdOpog7CPIui0XI97+Szxh9KjyDHA8dPs/QG5Uiq+oZfMll0gUcu
ergioyIpGyBak91m9sdZRiInilnrlaBowz5ektCJCr6Pt6QNzNjD/7/dTT5oJDSqGaKm+amOjAqg
UA/ypzppW6j1jKBV65P3u78EC3/AbnlFJguyyHWwBdge8UwO2hVgW84jmpIAEUnL/HU4ZPvoWfN/
x2IE2a/k+vEvohoHSabLp0jOx62voPmaKI/oGltRwmZyr20jEXmfKJbkdVhRAmc3ltUyzxmJmD7P
dMVqVtydhl+Zn/Op4EK9CqMhHeXGjnvnBujfJa0OglCKvCpwNN1QTCdrOo1y6B1r0TmWEGSnZ0ae
ilwuyDLJHDKtKiHlOahrkX1FT12feUcyp2HjZdb8RNOjIuBo1ifr8CwYLotBsaD1rcGPYpl+2um3
sxKVChOSfsxHt0wo9m0se3602DRf1izYnkdycOBwhmaV6WpvmxoW6/hYk6MhaZtxIqWNWmB/Gsqf
ZDjSRl6tPmY7CWehF2ooD2HN5sGtTTJMTPnbl/wOFP6RDvoMR0P84jWUqcaDl3Z1vzvUG/uVDC8T
v/qNtk2VeGtZMZbOfBIzgcTfUzCowIQ1BdpaqROVf0aIU9ystxMaYBdJ5ns9IVEgVn/sNBJuX5J+
HNK5OWyuyh4JTM388/z/xtNNxzBpeJJLbnggGJDnsbUM9uQ51K3G0YPVbu3CXCK/ZNWv05roSuDg
KT+LyNBwRaofUEWM2G0ywmzPO6z+42eZPPyKmt0kvkFTHS0mVjPWyKS9N6kmalifgeCFwzNZo7UW
Kx6IJIMZ0f+EgyKqqt2O/F0GmS6u/00wNTgt9Qczwlq+3eeTnci13j+J6JY0Cz4TQkqWlqoCAB6U
EaAEqgL1O6HNBCbHhCkHyygL/BVptWH2WWvn5dESdLGq1eT8THleePlgVS/s70kCgl3vCi2PjSln
raSzcUVtRYWA7kz0pFlrPJRwFLLBmI4wLJ8YuBT+9n9aW10lppuA4a9uAeSrpwkYigwA/9eAcxcF
BjdwH4ERFc5DNO8zHrTquSYq/tLt6F/1fG5LdzUoPGXiUyntJYl9QPu+arccB3W4O9WAXerLhNpo
0WYfCUDIOoFUkA/KDi5nPbRVtBajUDtKi9aAQt1JSWeEUE0uySMpYDIHtZnuRT/zV0CbKOxJfZcd
HSLpJkgThXNKg30IF6yXGW5ScaqYbkF73mhAzUKxECcC4d83ISekymHcN9AdDS6hTX4wHi4K919b
/N9bZKEfDUOq9Sm776OHRghPBcAMNH/vxA2+noqCw58m9JzUG0IEU87MqqLZwJUrZrnUi6HWDEDQ
l1c74D3JjqZ/+FyN0f4sKm5TKmrp7UWNLOfoU/1fGteSdbjKfd+qkkIfdqCf47xp7MTrWuKpAzJI
Rcff/EyuoDCY/v+U570Hu4fR4ls9RaDwAiGeg6vz8ryUK1m1RlA7paK33bFKBfLn1QzSnDBPXQxh
LF/14f6LABEZ+yXtUlaw0F75TCD71DD+A2vAgipRNlyIfJQNc+5+umH8W/h/kwC98+2eJgCmPVX+
RfigtFGfrEP2AQV7XnkAkIdX4clQDgnD0XAK4ERPGbWnvqD9ArBkZFwFW5pUOCpngPuYD6LyLz50
0F01wlMjZY25nL1c8i0Tr0yuwoi80X6sNsSwlP2+rKH4rDmDoB7Um/Ycoj+DvMqTxZiMt3GD+OKw
R6PaSabKIN8zM/5zggwJfzuViZV0iaGWsW2SH7Py5Of8Ha16qjn4UQEto3X1IGgnO4q1vYUtmbCV
yTVrNFyAhOyvv6/Bb1vmQl8fRgt0YkYqrQf8YHkHFbDjpHzbdIIoAUzDCD3MmN3jBPXHxHBOr0an
8kI//W8c6SZFQTic9mfD+9jt7MQMFzbXYptFdDnACA9O8TstnYWk00prCAjCx2e/S9mtqv5WSpH+
laZPpSxMW6NCqFTy9aTVIwgWeVhU+YoPFz86cbBGapKcuZthRTxHmbxI7CNi6ZqSn1Sij+FUPOL1
G91qC5BFImdoBc163ZIX/c7aqT1n3XOuzWg2Z6Se6CGG5DC6h1A+KC8oqQwFjrxdqXzF7jrUYCWK
DJagclDo1Mwr6V4CVt18dZxtncc8BvZWtmHOIQEoygoS8/FAnCTRdjcQM2e/zo7O3U1VFo2FRCKU
BLARaFKiLoeVITMqrEDfcj2btI5SGVz3Q8iaaskxChFI+LDyfADlu/Uvy5Y790AAXXxhpNK0jRQq
BdYZkGmhcS9BTS3AJN8VR9PA140T8EPRtQfBWTX5TzlBu0sqJZR4l7fScez+EhqqsVtgaklApS0F
ntAHcYUqfuNnPgLSUyCg4QL4rsXRbbeRMqxt3PsH5PwjevUVpuFBoKvwQNGryowuPQwuoftvyZFE
O2m/yRqfo+fR+aM/pTvHDkWsRrU2uN1BOmGen/XJNfJ5iQiF77U2Pi1IJmyb0L0xpXXC3m/cwZl8
EIsOB87VwK+sgYvj8bbubPc2W922q+DkxOFcq9Lk0UoBmW/szZwiJHpCY8zaofSPPN25n6IPSmzM
Mt5hOhGIfTZoFnVAH16p+2BKjLfJx1wA6ULPu7C9dvP88hSKXphMj2M91yPRKe3ton+EFASYnYy/
bBlA6PdoqOw9sJOVhC97uLtH40q0XEuPLb0lbT4lnVqmUzSm5kYu2D75smEl3FSoOssBwnrvxX/S
o2DiBwUprCXxtEoN8tflWMO3AGLCskQ0DDPm10N5H8/g7BOjhvA/jlH3k12kZuODRuxFSLrzzJGw
2i/psSy+mJ7qvgCaCXcCfL/RhuMDdSKStx1OqLaUR7kxGHTmi0En930FDVuqSDRRIcUktGD8yJ4U
byVeTPXyaYQOK8dP2BXjywEIGqQTp3u3NYKChLmDH8FeIPiC0kW/edCrFrOeq37mIupHUaLKKe08
sRqQKo8UJYXq5Rkk3Pjp10KcU7fFXikX8fgNVDxbCz+Rx2xzldTJc80T5T6pj5A5ZVw5MIuqCFiK
+rKHq9XsfTfD89WVxL1BPJNAO8K6eZHOUXCN2kcDXPh3HNsO6CuGFpZ4BmWUdiRlGiF+FdIgfvt9
x+9upApYyf1T8iirbSFr5MrtNfxQ7yN1r1Kg/cAl0GPWtJwZk01HD4FHh0LRoEPgfDRU21jmCrxZ
2tLD5RGDOMuS516bGAjTzdMsFXDDFOSh8ANaeMRLcarPdKcLS6ivjkcLPO6Ev1orZrxY4Q1E3OrF
vD0f4RZmy1ZV1DHnk2DkAg67yD91XFlqcci3tBqDzhSQsEnfMK96Q0noqylWzi4O9AO2iSxj1uln
gdoNktgE+Yk7lVkiCzZiO67+f6NxT10U/c7MVnOc51gWoVpCDhY+ru7zcuH3RpLKQ7TmawDOuCsm
DAwO0LKRTyC4Lr3hB4TAXJkeTT3ksptiBczxhhua0HBQ/eF4hJugKhV2ydM5fCh369lS9sl+SmfS
cLuoPoiNKu0uWPJllZGsPaiZrSoSvWDykMe0SFJFMNmXYBhOUXxolK94GgvlOXSjGJWFXZ/feGO1
hULaFFKNwSy6y8WUEnBkdFxeXy7rOSC/9YKV4ZbHO8AEDu5GpHo+bcDzuRHPh3GnZfXTUDnoi+J1
TEgjT/OWIxC+deljZIAiPjtbVKfF+/5rnNWPmahqmG1nATEoQmV910KGVqf+fpLAb6aOTrcKr8dv
RujK4xS8bwY+1ffbYndPeVaCpAffG8q+rhos+8hzjf47QBgLfz0kCEGEKSrfUhmLwFFWsQQL5qo9
cqNIo8+VvtSTvTw3P8YI12ICZGzb5h2E3v85b26l0ce+TE8NtTEYXNgiihSRrWLVYWP3PJcXXwS8
9IYXooEE1dKKzOxbiNL9hwl17p2EKGOUFts7MICqrhEUT/FjRlSd+tMj+wWixLw9LRCHpobGFFUW
ju6G27j96ZqYzY/rEfz3+GNTTg8p43LxdtMyoMp6Yi7f2aD5Ixuyb67GNoRncseUle8YGIbrQv4b
pgvO4sJkrU8NXe2IT2du5uQTzn1MbTHRB0iHF9Zo3xG7y0/j5Jgz4XQyIrLtdm+mR6mKjwfIxruI
j9shjBSsFSCKENxSfLnqd5tQeJLYe6w+MMuZJXA29qmNSC0PBzLgKuV3LTFHtNuWtmYtSTQUAcHf
yqo9s836fG7fIu94piAfI0Th1gNlxDZe9p/G1PrQBLeO+bNeInJ8d9xUvew4pgtdKfiXaI7VKrFD
kPCQYm+7y/mO4unU6aB5BpTcgp35ma+GcMBsoqzNY/dHmfmKcYZcYxI6zAl6aHMr7t1df98hnk0W
C+LLUb8ymAvPgxmKf91h+jzIitO8epW3ZrfG/UjsjZrYkgfxnniDm+PGMQJ81GqjozL2zkOlNEQn
fhW6Rv+a9U3Fxa7+/cNxnmjCn6uhzk1lvRCYFelt7Pbo/ZZqxOdjMva0hC4o4lEHC09TsdZ19ifd
3dZeYPpSAVsW6l5tTQh1Bvc5AJE1iBbAEuxTO/1sL9N2W0geX4F/cEX+LjVzwsR+lsFvyXJDctbA
9x4XlAfcLmLQQXDJ7XdOtRv2tsXmE8N6qnVtQqHWcL0JXhOwWDQZG20c1u4oJ2+jlr9znxPiwYi1
Zqg0Jf2jcXFb+C5QyZa5A+yz/JiFDsCzfQ8IDRHteYDku2bv2Sr0FdHk91YpxnlSOxNi8UFkHiif
iVQS67aNi/ICgCzPTNaeQedcLdJH1DvHHbNpcb7V1uGS9UYoCNcVE47x1qhM+yTP3zMwDV8idzds
gpuThz/aJpVeyEYS5+KDTzueqnw53rdUciAqEKz5J/l4PNxI58m0UB5gmbggmqrph+KjBjje1D7+
iTKjaVimmhfCb5JYmWKRklt5u6pb5knn18OKUBYy/ReLNjWB2GhF4FquQ9U73dnfYSMkR8Vkaocd
3OWizv40kmmyLqKdpCPFDRO4GFVpPCYM7vDAHzC0qtDs9z+0Xo8a5Jwk1C/W+86xgbnIb0zq3oaH
ifp29A7pqOHKIeJSXKs+6fJdJt4SDrOPugB9u3OEJYNmvx4O1Z5OE8XId5aw4E5QdqVRLsA0kYCm
zTVl+IFGredJV937ETBULQwx9OeXbKRoRVPuwrWVO0OxR5Yzx9e0saPkNlYXLevzcvhqXtphrqoE
wDQMDl6b/sXi2B6Cx/9lS99hjIH9OWyodEN9C0xDnhMOr5oN2W1H1P5BI7zp2Q6rrjlMDUjIytJ/
NyZRubPJDrmqyQZKGUFjfTu+eRo8lz29S5G3Qz6kqdas41AtTLYLpj10K42ZW3bium3EB4j/MuCl
eqDvlYdrwt0Eo+dsPPBuVylArxtVpeQyZzCm6sBOESG0Fs05Bgi4B5gUi7r4sa9RtBcZJ63jMLfg
w8XyX0HfLpMKM8XUepLCb23XPVfLkrAcOkPQLVMMSWcX9STQZyxGVn9xjj//v++z95W2Bb/S5KhE
SyP1yN6j0TFWbn7Bp62g7vMDN3ARQJS3mb3m2fvGY6Qpjm7b3IyakYw9+396q2XP60hHQqTsPpG8
uhsOnTEnSQkfHnX9I9bkSMB8Cp+vajAdjxfwxGJ9WaSl1FS9GDgI51KGkDnSHE9DhnQy6Mql6Lnt
GdAlIog4hwb6Ch2WHvw0iXuo43vQnj49o9wq2ovlSdsryNFqorrBu/SlMQBqfqcABSxFVQNssUhy
N3KOM7gBevRvfnuECoqbuvoahcx+oKkXUILvEkTU9U8tLyvrHcgRebsC3PPBBjLnKPHLOl2CsOT2
1Iek+xBCFbHcw/pCw/2dTXWUFHfMk7y5A6InKP8SRDELwzE91R7HmhjZ5WOlvp3Q/oV0cV4JfTmd
NLmtZM/9d5b/ADrzaHD0BMjPYSibQpJZWc4BWfj1I59MVKAMmjsMCUnFv1vUVzR04MmF0I5q9lGl
GRZJZv6AYNrSeaJWDF4q9LtTeJLv95rncDY37iVSU+gXW8jL7p9V35CkpzBG9E8VJTFUfOwzMKdm
kFRQEQ24hDkUU0tWEdfH4K3YShaUUSHFfsn2HvYFHEu64iLfuYCy/yZzun1W62RC2H3qXtWPXnQA
bW7fuxev4K5TEFRVEYjqJmVoCAc9/wb6vLmPwzsioLqcy8U8f8AFvo1luF3CYhGzi7z54ezvQ6rP
zXCF8ShCwa31VU22xVaTqKJM6mpf5FNzxXuhvxEqybeCi1A6YpnDqVB5IrLwaxpRQykQsWRMMaJg
h0vBTYqU/EhDC56ZlROS096xDLWASlmJkTUEIW/QenAPBxCL4XlSjS/hRVsIAc6+8lcNsGbgweUb
WJRPQXCKY2rElQWMGGtm99wb2wHxDsk/m7PaPrl/b2egHxdt0+zGcsbZsFj8S0G6TxEBQdyQWw7X
BUmY1wgwXF8+2Bcoy7IZHvC/+3MWLKuYHA0t/9uZ/UsFxBwplUse01ACMe06TL9JApsfnG4Zw2Md
2yhQvkAhHRyrPvIzfm6qEKePJVTAHr1qeDDf0RztUJcr1GdyiX5cZGQBJyRxx3S9eJENHl7sqyve
yy6vBiZCA4GqFpwyz67LqHdI/+BYg5ZkcsbKQthr3L43GZagDAVO+cpZWlNRybEqJxk2K9Rqji9J
YizEcS2ejnAWmLjaj71SHdVMrZFk3uO/laBzm9TN8Dw37PPTwk4EeF/pem19F8BCjsszMuEz7uZq
3tCEXNzORxkW+DCnBdNAlT3x/nNPmOgZgLrZbN4Crpa/ywHcuM6zqLinrCl6RFOmF+5hnKf/HSDL
8sxDf1M0VzAYsIAcNXoNCiKGdi9pSgDl8PUNCIYjXurRyEpp8cR0peApD5IJO5Iig7Bdwv9akL6S
BfRxfZaf8Ny2T6c40h2wh492ldNayIxM2fjtQyXBIOs0xXXsYm3gjFH0vRBU0IMd6iOh8iHCSay5
Jnf596ZwytEWWEkcD1Te/BjumaUoUiGQbLa6e4boPydmtwPQoOD4tzQTPfbD2VvRZQCzaZFYF7RR
0SK4DDyACrumhHqc8yGkZjTQcevSImLDdYRSgGlPIP+rFoQFBNizXFLT6GYZj4fz0J4BJvDRPFJH
vWWbPCYRurSPbfC6X0V5LUShfvOc2bX7B+mtx+PBhedaviiZK+KKC6QKL7EUG6kMZDmK4QYwPnNu
u/xj0iHwMvgObj0P6Y4GbgggAsRT+V/XF2KHHMDwVDp4XnBUiUyV81kU6rC+tvFsbFKWpprswvOC
ZJHX+x/sUB6ABfD/D6/z6abVRD7dHnUulYYXP6y9bgzaf8V8BFdb5zDqTSkiaLxagUWWgp9KPXGa
Y/eKptgUuXICc2QMI04yoM4HAPhYnvMSCfZrGsW33lCStBoFXbTlu2gvIM7UY3IjZaiLfoJiuX7H
JOIcPRZvSJ1K2Eg6li3URIaGXF0ICOtmH67yInAeFLPQDg7fhw+dk+XZ8XMcHJheKNMTTE1eQoSm
7qvvueHOCzLhFnzW8M2RXIgdGWhJYpV+mXF3htno8pCcLfqj6ahohauxkWIt8SBBqEyLTiC8yPLv
FIqHSFYLQC5d9stf2izzu6TGbQpfE39EJ4gHgKNr214rTS5UAhVENebfxy+4biB78G4Iw5KR6Dki
c8qS4iKGqxpD7/uKfqLIFK2ogVzndwnLsZAJGr+jmyqlmlAkDlAywQZ5sKNW7hgcDkVtx0sWbsym
6EYI3PYpbEpPkSwA6p424flWUMfuFLgqDAGVsxa6gxjoxE0MSYHtim2DeeQRiE8HVfbQ6FNSWNdM
zVFJHYLWt0moRRgOl8dnsXsKStLHWfoZ6QWJMiTzm/vl0GMsZl55aqIWHMe8IhaEYn/P3RuBxKX3
zido+BeD+nLSoSc6FN95aRsJxdjO8NOEfKNf9eWaddx7iJnQr4FbQEn13KQ7sCCk1nGZwsXtHehU
1NxbyYPhJs8jnqBf3b4Ofk2KytTwWDDpfMq3upcWEYoSa2FDnohqaPbAYexUyAPhmZUZ278mPLni
DziTzUVWeKuuRcJ6Rq06AIAToKiAI1oADt0ysG9MnxJsW9Q+/+AFNzzRryAKzPDkpkTw7HL4eFvY
36DP9/ekl6dJkAubl8nB3RDQmb7iyljPibpI8Lc8lpTsSR65byPLyg5zEX/+IDqES9mrDZSsCVl7
LNx2k80MkHIuzLiHcroGyYd9qlRjenNYlqYnATfDsw8NgR9G0FBp4bGz0V7UrSuM+oWBbid3fehI
HB3sPt2ojF7xRmY9z8yGNmvl5eXgG1CwXcSS5oTUXzjXeoEfLHTSsBmJs+l9tth8tbccMxJWDEfL
rRvQBGr3bEAYs8GQ9AkR5ZDMWR3bSjuk4DCbCDUiTUH0FDduOgKb45nVkW4+dx5EmUWrd+igQBgJ
ru1xZO9Q9rM9mgbF9J/RZM/3WErDp1l/bXP6ir+gDoOIzuEml9qA2DBF3MxctmEqu53NKHTsb/00
CnG8Gl5sz4BaI6Ucr2L6SCLFvfC8epoLDXYfnRiUlngVgMYSpTCmw+sqYt/XTVqw5+d1uxUsXwYd
oUwJTc+KD0i1wHhxcRo0GeMzUpthX3Z1LN+fH3QKqNO1zPNS4fUTsvWQWh29MtJtei3IuyftXdPl
8JcpmNe6c+lxlaMm5Ez4CpWsjZDv1ESLvyNyGEgYv7vKc000c2EqMoMZTvwwzzFQhvFheK1Qsg/h
wKjHzYLWEqum3oKT9H408ugf06uQdrl8nG4yeNV4r1HG03k2a8LWMvujBU1AvN4UaAgpcvVNWDsT
hcz4HNkcE79lwvsyG3wHFxDbnIlL8/2owsFiYmgPbTcM62s80wjLCWHBaJio9Zi0xnAK0cA3hl2m
+v49G+nFBdRUzMt91lD92uMrP6GWWKcDuhDow9urrabsB19CUoVSVHsFJl/mUAEmkQ5PqCIZ5hWc
9D2k7fcIRg7zB8tmizNvdoBIWY9aXnaPszwUt7pxGqt5hB4yvk63Qo5fCt7dT4i0mpqzZsCnx8Su
n4Pyv5KQCYSvWBGpb5hQAnpkyhtv3xCVIRjmLxyN6LGfz41GO3SnnFYoM+zGyVNuqvV1o9ksZFGp
KDtasforTyeHwMSoqWcZnv++fypGxFJY3sC1c54PwqayG/AlMcRLUB8KnKXbwVBk8TV5wjPDnAiI
+PppjZ5js8gTWVz72J4a1qCpO5BfJP5lYY/yi2FryKY6liyKdVcEJIJujFKJZxt+zkGyLMxYwCkA
3Lobi1DNCRj8fDXQyJVanAyj5K3iHOwRn3tQBlCY62+YFBMUMPIt6jLseaL6lNYmLElA1SD7jwS1
iVwHBHTs0LpTlZ4ZyLr9jgZnFxANzeoy73cQvlEmGnsUIeATsWZ9MfQcSwGr6g/0FJIaaiGt6LEK
Zjo1Vvm1RRoCls7JGm+R3yUI5XbM/UOWHNiwXeZ090Djy8hbK69f69QtgSP13LHZjkCV3+pKoXaO
QUQg3IdZ+KKcrteBLte++qUXK2H5k6F92urYImuuuocFmcQSGBsYnwVxmggEq8cacTWU0G1SRO9p
xLfj44HooKSO88foeGV6dxCXFPUVyqNefwczMw8Vg6KhEz0v3KW01QMJGmB23LCkPHQ8e+1DMpj8
qSp12CgGleIqtDE4UyidJciuJqL7m0TuKMq3F9rOXiGZ9K8n1GLLYzQ/dTARWLhGE3G22ARLsBJG
W1D379jjToLcAfATtQsA8CVeIQtn/Mq3GyFwoY+9Igs9KhlJa43LAfKJ6oCdolPIWKM5z5ftquG5
D94bDVV/BwqZ9b5dr55v+pwa+Pd7tXZGeGr2ih7r8KTszredsWuJrJp240VlrfduAs5TjzbtbQ1P
EbDdqFGIHUniytdFsFkuFxL8rbKa0rSFdCpyqHDlEmO5zz3NZXyaf8d5QgTmvh3smY43M+hND6Jx
D1RJmFzqviPl2OAOgrKbADdd4dD/4nHMSB6G3TnCShqXBahE7ZthFrY3DpGH3xAOayQ9V/nx6Hzm
FcrnBuH+OThvU403+uj5+5l9930aEJMpV9RpSZeu/a+aNQA9vbVjiKqE4t9mGAtblnp+gv3VXxKH
m+y00t6cOiuv9Yvpq3kgqCEcukAJNOYca69PCwu2jAguvzn+mSOJ/W2bZl9Tp32DKg6MUvahlx52
EaFy8QQQAOmkpvkF0FdAYpKlDlxi6q3yBpZPJU1IkS7chHjHPqecOSr9hv0ww6Z6k4NO0Vf7bZ4K
ZCWxpawSA/E/lNAI67gH88uIlWLsOgkFp8yHKhixVBpRVYe77qMMFib5oZYf2uKM8Cq8PPrjG95b
Bx1EpyK4NrtKThnFkDBnhQkE+pII4V+78x21pdJVVtq7hPV3FTJS1AugluD+a5uZJL4p9TZVhiQI
lz49po6sa0fBPfoQ0vDZLCMliLKD9p1O1HfwqAjl8coPNel9V8Wa8m72Pnlm12pG8kmX7MbMDRo2
+2bU9KREWhJF/ZnpBzfpcWi/1Ir0WclJRvFgewInHhZJvZ4Arjq/JWf5FBGok47mvEIq9SKBKXZa
UT0EckFZjsPmCMhWJls6dGVHXzs0J/mJn4W8oMDHVEjJUm8D7ttHLakHXfX7l0mnKYUa40Z5BeHd
eigw/n/H6BNayI/H6BdOD/qB3JuUaZb+vEYZMR+F77+Qz+mnbygTZTTqXSbYC71NqMctmbPnLh+H
YLSnG/Tsb0ioQamKMPGu52OaZ4BU1hW1xXaTeq2BVLy00+WnauyGBbxu6xnCA7525lhIK3w1MOss
SMyvm8UefqwwEpfqRM1lDcpyCL7P/5dlF7O4F/QSXtjBdAyHxaetjSRfaF8DtucimdiGk12Vh7p9
nlEK95UDJJmpnOOwbfdK04gQT9iQKVSlOwd4rvP7idp6njG+TdSkx2xRnivOk1pf0M90D/9vFsZe
X+QwLSYkKPoEfXqtWaoEu4jIL3bW7Jj/WA+7mdTrEsnXZIlDc52oFKxVHoMUg0YT8TTsmrWh47Lv
m3OCeGZ0RuQV1cMNxyK7qls7MTBeNU5Bo+/gYldz+ug/8ipmytcYWE54KLGt7P111ci7WjHxzgQq
kh9bC9GvFQRg77j8CX9WPpcaolNIJ9JReIMxsAP73tuooYctE/wS5cNZoaXJj2banuZY7Vb71Lju
m+fc0YFFUKrcqT+Z/5Fsn/+4uEkTHYoYdgrTvyeNFN69lgMj6G6df228HIm//+wszhdEjYDSgNdj
s8xw9WJuHhUpWbWlz77IczDBY7J1/SN4YpUqCLFNbbUG3vRVRUlz1A//xTE5ssu/hQCSeJca21cI
0MivaBP7EVbtu1sMmMXGUmZEiP3CExqXM/Y7csT3oUDSUUKnUxoxtc0bd7GjQV/3miW0VxLBOYWK
KyNMII0EUt9gOk0UoWEJUjMTewO5EiyMJj8k0qP7z2vXj3jmnSJ7ycEYiAeByq/wU2DdNM6kFd7W
z9Fu8lxvWvhy2eVomuLJkZINFx60/p46cokBvGbFkKAn64MZj2+7fV1sqIq5sQtfcAZmddyPtaxP
Z4j8ClFKMRJt83o21ckxDbniFgxYAD3FPomF9JdUXVpz4SoGGlRpYOkp1iRYyNEFOqE0X/TwNF0d
B1WiBOR9cWF/wz3dchR88jT0usmE566ZWkkRkHHTH3DhziswI+Ya4w9WD/Svme5jwWzKBeSomVsA
Mmg5kolqr7kwKzxA+Xa/CBUm0FkteE3Xeh+N/kn5QdDLDv+afXWk/UD+lhW2VxPpgCSEGhuD9NAJ
eB1b5PDHk1y0PEEWQdb0Wi2B/PpLqehCK05i3lVNeKOFu2vyUxa6jDIxn+hNpWbTpC4J0BWjXoYd
QSdStSQQFChKMxRZd1Pd+gdPp0hvlP2yccdUNcMAY/ngpCuWTlIgEqcDWjfDSK/YzCIrgTUYzpEs
+nwYRvTDuK8gxgQbb22zWyJIrfYmX7znRgGcd31Wc/wThCvukhPHuWsQyhCtnGGXKQ4V1y1eg65g
rvr/t8GDDpsjxTZH8vAWPfJke0Uq+qLwtgZQXlx8HrDkQIzMKHwIGor/31QBe6X88Jwz5qIwQx7Z
m5KGP3o+JI9GKTtGIuasluf+Ef003P+k5LuhFXHNQSn/zGov2QGaikxGWN7QeTKPxhAG/HCxdVle
4FzcwOkxDTRMA5Obak0TlGXZrjKM7VMNQQnk/Hxtbtj4gfZNYOf2OIYhk48YFra5JdSOhBLGecqE
l4HOyuKXg6a3TqFR9S2AaJFuSgNMINTLdS5/RfE3c39Yf2T7XQkbodPg0Q6pxBsqWV73+5XkzaQ3
wQj+uduUIveKLGvJYrZE7NZj/N6KLaTcK3k2yasDOS4gbjFqor8Y7fnmKwheZgen/Bn0eaDFPY/s
V0MMf2ODzvCynM49/R/C3tzzoic6YMJON7+cW0M8tsvOAO0z4tCQuvIMeJQ/06YLqsPtPH/MEU4P
ef87TWQPkAdSX8J/fukfmWQVzT3O2hmKX4lxinJ0DIuw5wVqijuM9oiTOFrweNyc2lp9VX3Gt4pD
XBBNApfhFk/sBOim3dc01IrGl1BZ004O2ONncIIhbDv6nsPlfr9GgegiXXLVTpJpxbCm0FbShZnJ
fLkGin7W7RGMYzw2i3NhxMVm1S5rNtmpDE3YXxzTICwFxT764e2TcGSnCb8WqiVniUtWiuAcAKzi
fA/R0RXuq79nvDFr0ZAM2B6p0XbFdbFIxUL8i/fYo75RmCS1oznFZu2HvPzPMsRs24QEThemOwR9
pRT1ya7rJ4Zo8dcmtcH6OQEZXXU09osq38SetJt4sDvLXy+WK46pKVa2S+atjMh1NiNvWRm0V6Qb
v73+Vl3NNW3e6K0Aev9wvChsD3aQwuo1zm/UM/2oIDRLHRA2USZIhgfBtQY1xs/TZ8QwBmLnD2l9
AJURO0YjKxFaAqmJ2t42czuFvCbEgHA4ekw7WpjkDwa/TuF7Oell37ijGA6eswXoLFLg2fy3CBaM
48rBxR35LhWmH+/XakJwHuGoJbbByr16GCzndVYPBvq1SS5eR/KarbiOGgALJAB34uvHgdx6jyz7
XbbXKO3x5LODAGEFyYviLcXpWPVKDSKe6DEETfEzKt2rowGpUrAEdX0FuazelGH56FsnypBwyZCq
5Cs0Ri44XOmTsLmUHk05LELwx3EYcV0dQA6qnPaSvEYzmz1SqMIfgX2oB/PhMjlgeNSx/7BSONBm
/sicS3NkoG0CEqDCqRVVQdl30rYFwdX6d3vK5esDcOR4Y/d93dTvheB8fjXYEujhJaV6aFXOpF9J
SSCNA+s0JTRCzdcbbaIFBRC8OB+yXPIdYVf2T17gXRzql1HfS0jmzaP230oNm29ht9CCAs/+9zSV
ex+VAH+h3YEmKH/wpY894S4H/Oh0AsqcbxJ2WfQD9Er4h2hwwecZ2fZhqCLLstCctSQoem1H1PdX
rvGALwoOzg0RDa41bnN1q8XtdNLU5/Nxu31wlErl9ekVwmWzCkrnFFd12PQ4h03+zhwGemXLGKyI
DEzpeeSa6XFsTxzJqIZVqEuwBX7vz2bbRB+q9ZnOWjuLzbzitPSbLTw2p+pv7YoOlMticYiboIjZ
k3pljBO+5J8MgqRHV72eGsfTZxwKOhiCOxO7q0Bd4poHdrduVRbVKofN6zBVIal3P+07Jc4ANkXq
yZn3danhdDUjh9YCwBqeCGuPesSt1eeSJKgdhmGX6eXpmuE9N6aazTXZP+HbND2phLPpHUTqm1/U
TtIfEv1wbJpOZCH2uxMHU0R6T8eaQ74o1iUth2HR1aAWv5yWP5fRRNfYie2p/+CDTQbkBTMmcVJy
lZNEFXF2TzYgNYEPwivB/G0GTCxQJlG8sJpk6YSVfP7hhBuayM5l7v5zTItiA9nSr1sof/kat4Mk
0y3vbky89D9KKJwLdfSW5YHbbtJA7Yr0eXpbk7KCwVcU7Tq48MZdpPoyvnG1kFOOabUkJ5zPjHgC
dRsBtpZn3qWMi8iBc/FulhDTWY46LF2ElqiLa1RuWSEyHGIfQKY53jeFqi9J/VAL9Tn6twce8a26
kaDzqbQ/LHnGLDajqV51U9KhbcL2Wy48yEss0PiIhdnDrEC88DUdJvLxt2Fv8A3DIgmup11M9GNO
1UBN/eNTIMr46O9CjNZz/lv31/bDmrlNRUe2t/iKCVnUgv+acxzLkhYa86PnPslootDnJPeWJD2m
v1TRHpSEgJ6FHMKvnSzBAfP483ttXK6RX5vYBQd1X+FTIifql15J40nhIeWEW+5cc/3N29urNFPS
KLypzhmHEH4Mk6MH8T3gj14s/kXIf9SyCzJBKXmVxRMLlOarDdmC91NYAoyXpvwr9x6XNNn3dRO2
+GjNbJeJk3aPiHDErjtuXo4L0ijxw7nYHoNwj8Ptj8zAKZ5ZB35C5tzP+245Gh/J8Qsx/aUOpBN1
9UN7aIlYvnFU9maktq/i6beKB2OjecYHMgLAzW6NS1BCAkaqaGs9ov/AYsacvtD8jujoscyUHHWh
wLoCSxFnbu69Xl/Mk8TBb97qnd2o1gXxJ+o5WafrcR6oOilux4y7pg6WFumw4BRoe5wr42yr3VPJ
oNKNuK+7ajORjSaDz9QAKtg/BTXhUuhU8m0LWkwiKMSlObFx2gyPg+Xi8y6BBf15PsbevPVXEXEn
HtzonFhG6BMDxRDoBluw13hWNruR6cq93iqpW/0WfCYABnD29Mj3GlbRz6t2ucMZoaa1FNtszaQt
7UPU0Cr9kqFyZC0MgfYU/dI80AnGAAtTC02geljYmKG2CzjZDCe/nvxHNPLowAu+78NRr/EAqrAn
ZegCQhMKNUDsODFlpC/Zk0g78mJr35WN3nt+9yi0c9PaHQkqy1TtaUIUvhH1KhYF9R2yBvYIPDER
pfuy5/OgGkESPorN2066A1iIHyG3Z3bdwThbfSkNmY3mbKi2AvnekDLnKlV+BWucgNQLuSQS1RMn
niPg9kDa5BUmsGD6/bXTS4dZhO71tD+T8/rk7XpH45wwb78ELSdBncxcTSHmRTIoDj2gbeDs+bbE
VfyFGc5ad6AUZPudV5ojlmvrGRsEak8VPuvO2XuDj5xPIUybfsBUYGeyRrP37PR4kMxjYKSK6kFC
YQii/I1OUL/1YM2StyeLJW60cV6BiXmsXYNOm/ZGCa8stajLDzVgtpBCi3WgUTHcWfaUnA94JXi7
Roc/t5mklMP0cBTfNGGxIQmDe+2qFCEClRSX/8vUnS05xPBjdGQI9e9oc7H8H9pn/ai+/Tl23duY
PzR1UABgVVQeMIKUgsMLl066xZJurt9kkwWNT1hlExQvSxRCgXDN8RqzWGCYNQrob8QtCe8sDPwt
OXrCRQ3OEe0w1ElbMYSZUZk1lL+50oVgIUWS+tfOPfPA6TcracWx8JiCzMW3JTPBFiorH9YZ3HeD
BdPpnS16x33/sRDWcrKkQt2LgCLMYx+y3C2z0XsYGAokcd4Lz8GUSXS+phcR0+YI9+c68hAvNbt7
vz2c+prjLyyEVgjy5ByUqHkG4AMgHlp62dmtUvWBBEMJvAT1xFckXCkfE1zWIVDxc4iXhDfYIpI7
kkwplTev3yxRlq+JCdIwC6AiyJzL99njrf0bi6/5u9U6Jp0Zlmcop29XFD18dpcMzg1ne9rDQUMK
CbkXfN+XWeT/xKMTC2mBzkTFjL5ki9iwH+WtwO9CNaY9+4ygdVsiscK+JaX3bW2K5KB7Nwm2Jo8W
RN6o75FlmSuw9YsV+TaW5ozY63wqltaXrAoPfFhecVcyI6JTNVAiBfa3moCl9jliYnhXvATwYw5/
COJ645Tz/LarEcQ6Syp6q89ESSZEmf0QKjZ62b47FS/oBnee25fWMnQ4BxotsErA9K2y6PaLfFCx
surkd7z83eXjuoAiB1I7aEwapawyVYRla9k1hQByJ8VtFaGsIVXEPr5TLvoiP31ydUc65Q8+TY++
T8KLW1txf28GblO6Q2bl6yF/W9xaJtULcvPZd7x2XDc87LoEYHR9PkW5MT3V6lLnf6uj8ULvmr3O
/d4OxWMkq5rSTE3qgjblB6gjxYCdd6I2jEcr0dPxjbClOf1CLEWpLJrSdht0JTNsNMGIlCnZNJEL
iZihteHKa8Sj5q6cTwQChpiOljT14R7wWbh9hmM7/9L05cP27ZIMV5m57qf/02F8ccTy+p+PG//b
5LNlGz4uvhzkB57tvPE21l1Uy7cOvtVmTBL5zT5RnLE/AMrIQTFEq2UY9Hu3qTerWHlpUZiF5DaI
xZFht8UHMzsuZI7h4jxIFM+p87ltv5t1VmtEjimhDrjjbNg0SmnY79nqtz4SDN4zOCVjeY99jCfz
t1t+yV0mYE6TmW66scTBIjBaDjufKY+Qv4Fx0Jfycwfw/t2a7pcUNhw4bh1kFD7GsrpiKSp3bFtP
fTTzOGklYwCVQMmd3U26Xj2KbiBiFmgzOYNAeUjxQ9VqNx90id5gxXpR7pTfZn6JGANKPA3pdSn9
HHsspkAbcwGpS1UKvZi32eV52+BWDk/+oqizwyb6oYIndPIlIvT6NhCaI7wn0cfU9rj40zH1cCLG
riRddktWZs86ztFef1QSoHmgO9hxQNTnBhJuo7HOn9eW+WlPMA4UpmbIiuQKC7EnMaPYHxkpB3eS
mHiSgZj5XNWHKfJ/CZ0P3KnNHoj2iU0BcMvbt0kG1Ry9wNuvKz8l631++GqwTqLLfomEGpWDHO4N
jOyQBoU8CTBzuHh8VRfvGzJqHjFa7hPs+NN0V3kubDJ0408jh17hFRmQ9VB2jPZv5PWPGTv/NFZj
PQzKp1i2EkdM9BKSWMP2HTZ77lFZsTE9tlw3966mDc5tvp6LLjBFSEk6Bd3a1h2E8OjSb1KgTTf7
vY1N8x0fFoma7U0+hHo11ngrPIT+/soTLpfZUJJ5q80FdF/Q9HHlo/uQql+kC7S65vesgK+lum7n
ljGulo8dKZv37K+DJ1Qopzn95ayDRBEamJPL/liesbxrXyfATvRqyTb8QZFdj9k137Oepq4/VFO2
uu1fjoodDiNcZVovGogRq3Fe3SoCDtuqJMXS/OVOCHIxM5ZG9lwmbuWu8oi9U2/y1qdhDWTVSrLi
R456cp6GAR3+gu3S9ylHmDhSSBGV/dxhtOk4xIF4iU5rQs2GBJl1gYH/OyYIAJDORGo001+fpEJ8
45mhCWXXsDxZt0radAmTOym1X5QBsZWoIEVUh8ZRR4LFTnxN6ueeeuiCBBP8qa7A1DBxX5Gk/SMm
05oEtGQzo2TucUoatvrPml1nyXIau/Rp2hdAijkEDBlkh/RgKBrAjYgszDuYRH8liJIuX4OM6LAU
ytX1XaMSZ7BGYRNy8UPlP7kw7+4DxPPOiP6YgyEDd3jtA7ADmIMJEtr1e4TUsBP6jOWKFjFFIOAj
AXQZKrpsfkC6WgemKov0RihkR4XbWj9ZBw4DAFcd4WhwKKiPdSsNbPjhyHWLqVOP93UcjZsYumS1
XIzrzyV+D5vtnzt7QDDEdIQRdyMfrd6fNuu049iGEsMIcQm+sbm6duRJ9/7EaLN5ZHk33/PkcLWU
01N9j3maernMH3BQfIXR6EKluaxIx5y0XsJZXVHTyLbMc1XfgcDMgn0Qtl5PWKc8bDqrYGAa9iIk
zcSHU8A8+9o5q9s/oeYlE8znX1xJfLlg2bmujqOwjOKXb7ebK4acU85dpWZVmrNz6flHD8QuiujH
V+J/P5ADHBFN4ZLmVSAoZ64SYcWWDvajiySPdgUXXW3rBQiCdUr32QOblYOqtf5Q6a985a6ZYYng
Wt+tJwB3/igPW9iJBFyug+94oM7TqScdP6U26kP/LNamlOkv/J4nPJvjTZSx8lFTkBHbI+x1uwnW
4Fb5BMX4sXZbe2uLklKlxdS4DdnZZZNXqjWzdD/L/pd5QREnrC/3l1cu+Ajp3zPcYyoPa7NN0LEM
pT9UM2CrD+Hendypw1dqFamQL2NK2iqeEHoi9TXkMVo0kizh1y1oCv4VLEi3xja84vgxbLbVxhsY
j0QpXvimWT8vt0jRaFbyzzaRTurmHgfqkEAxQ7qxWyzKjJmwrM5urQV/ylnPk5CwwWaXAh0VfSW6
vl9+5sFAz0jFcgjCcNaFSDsxOw5ER4zSKiRocSsvJc6u2f5/H6tHUtHALmOtN2Z9QMQRBJEG8sup
njUoi0EakKKLpRw88LLql3ByMdXmB988fmTqwYSHB6TKtUcMAECTwGcAXLE2sbS2or0VPAGom8XW
p+5eekPO2At2CtaIr7tCZG6AOFg92THRZqQhABKYth1dHuhH/9AGXHcz5bJ2PIQVCXSME6kyXwgT
zWuLc+VcK6m021JiVxLP8z/EccX9BwwjQkmql0UPOHPi9keuDdFoiVGYk7Cqkp0MMn/kbToTaY8W
wWz+Slln5v8A0mMDvruQgkH1hzTJyw3AUsdH5tzlJLunUfH+EX6f+aQSLBTaeecguS/RIZ4t/DbT
E1hWS1VrVqpuVqHkAMeAgK9bU/ADUSiloVPMh4xa5OGwYJ3l1WhOIlk1ALbZdXbDvmNnxJYyIB+6
9n9s/hFFZJGy8SPhl3wfwSzYUqWOmv7ke8iJMDSDr/YM6f1wHiaJpDkQjjFY0jDy7k4xnrI6i3AA
Kx67hZEaNjIE2nJj4/H9C/c4KxYf/lXZHP+kmgJS+2VvdSgAvbasCBsJh3+qAT89DfFX8ehC15Fj
IocnX6oC3O5XYQ8Mwyy/8iXSBGzLcgpbrzWt+oAig/6MJ4CF5skNjSP2+rCfE2mjv4OF3qQrWJfK
WJUmK2CQjTMAmWTkPbgR41AiXrllbPZFOV3xJslF8gaKlF5ve1WrVLeqQcqdovhrqn9ktWBObU5B
BIDxiMCIGVUD3SvL561JmZPEneGaO9/A/w3rna+q6U32KipyiTPXqcvK1/Ni22lAtUjO28LrJztW
uJPKDUodHqAmtYU+iXc/o3w1GH0iInTR10JjJVPXHxUTJwtYUu0IJZORv0vR4DEM5oRHYKYyy9Dn
dzioMR4tUnxUML49cDBaNRuGy5o/aqDidb7+8zpKpDlt4ZL49tS9LEswh1/w4iiEG5/ospGcVRVS
komC6V/0LbRTWnL6U8l3EgXhHeaq88t4/K+FVvaJpxOHh1sIhQrc6rmODUFePRkLcoHzSILwsSC7
a7R2L/nI+2+fbk9KIb0iuERtglzTu6mHrvugcTXwN6b/8725+shmHoDER/A/DfSavkya1GpcZ8Hz
wxBbvj/Z9xw4BmFcGu39bExCC9rKJSZtcF+AWgw/irATnw2VDosE/NyRRaguaz6/fgYBr//ONek0
X3TMtaqxHpF7mwhyxKr4BPbOYbkAWJ9pHKufSDWsOYV+XTnrm6ZGV16rVeN3oUxMEp+DB6rt83/T
AcrPPbYty2FEzXXtbIiAANqDfFJioZjTlUkoAYHAerxtWgLTXvbdgkXsrCE7cxLcW0GEtLxJVapN
9so+Mg8ii7Hmci7l9UHMQQdxW8aKC3pF2/+UMKTUsT7WSDqF5XSC5ZleBkbliuRgG4H45Lw41YLG
hm+ewhqLIey6l4XcauNX/8OiIfSB2D8T85K0SC29TFxYHh41bBHtjLrHrhkCZH4sCPVjlZf/JKB3
cS/SYSENoItKXeYd8CBW58cC4grL2pCtoh1AwA2H4pOYyCh5wTmFK/JWAyri1oIIdcGcPjJbk3pM
zojHq5VIpA6JhcZXjDF5H/55YzAsFg+qqQlNA/1Ek6nWK10T2z2RFwWAh58p8AQ6y8xv/r5mZiDu
ChqHlrieUBzYdEB+WXycnNE17CnrDNxOwO9lCNjNuHyhss/XSDrmA3Z5q4CSGMDXTsHc7blRB1cN
HcIPPHhpGb/WmYxIeIBbj7fHu9fzjPEvLlQ/f2XE13TNVQhxWBcstrN/+U2ZdFZVS1JAj4jPLOkA
WOD1hqbHVJEdQj5QAcC6n0nA7vekMkzICmLWc4CgQS/hDYaDME/S8541W0zpLitrzkxZbJmbxhj+
52sXpgnllvoOxM5IqGJV5F/D/HNqXNFytCMIw9pqDbDoGIG80wKj+n/zetdwVNk3ZuAlEcA3Fnm6
/ZA4zOEFFymK1mLNMhdfCBYCWQHiwF1mNikahUuGPb5WKaA+A+I6N3MvO5h0OPW8u+uywQaAXU4t
q6igflL+0jUpagBjL8oSFu2Zk4vr/wIGTfIfnGRLx3carNeB8xln3K5N0xbN9BNTBN5YUbPvrPA+
p+TqjXRTuierVTgQcxVjCSTh/G9Z18/WlF+OQW6DezH+yu9tQFb/jEYQSQejyAw/lT54tBuNV2D9
ko0F3T0eBL95/7jBgOOTax8uWJ1YkDLuChLoYO5uQ+dTRwWF60LXLrV1Ly75BxZpR9Jc7+CSU6/6
zTsdvfkoIlwCAHBFD/IH7PupIKysaAB6HS+O3p6oiwSD0NHAmmVuJz+FS9QT//fzmjwpW9hkNucL
dBp8uaoVSG3caTjwECyHnU2htDNJyCDPiWOcOGE3A6S8P4t6xVh8pfqyFlsqV7dTje8Aatgu6ruz
BwoYWs/GM8vhK8nmOSeukFYkpVS+ysBrTdpZg8oiX/kJqpYLACJkWRo4T2p4dLDLIE+lsXFtUbrF
p8q4zEQSseg7lqdy4iPcKIaY/I9HIZa9dMN6Twu54ZIzFaOJujOeVnr26m2yOtwoNmqBRE+f4xHR
63r6H7KYUXGrz3tvFGZtVqOIxXVr8Vpfq40+3lTtfXhxdXXBdOUQNx45UpyQQIG4GtgFdlisqHa/
86wxZq0jGX4UdRNvzy9Y1OeUKuUcMCVTdB2BP3IUD4WsArcl2MU8iiErCki3iDq36ouIWDj/DQY+
pQABTvKlyKUjxG53gNOSOEZKbr6bfiIY2OHKAskBUrVmLTQ+G/TUFqbiIMfJJqciA09rw+J/ryMS
wVE5gFq6Xki5C1uFaEauuX2pcU4Cjc/J4VphVyha63vocBjFqGTHea7Ygq5x8RKzWdBw3CHWkEf4
uZZjJqR/+3T7TvC0EBg7C5Q56I9Xn0bDo1Cou5CiBb5V71PKf7P7IHMU4m2pPmlXjJq941/458X2
dX9Z2TKRLYfh0a/Tm9RDapnW1Dh/KQzHi/xKOcXgmZpsdu2YXK4M9L9RUNvrKHtOR3Ha4fc0DLwL
Nz6dF3vL16SJiH+wbsbtoe8HdyQm5e/l0HVnKvYT2WA/JoTuRNQzhYS36S/fFXMBgmJKZxlptlYa
kqGsf6wM+mBOCoadUX2esZun5/e0VbchR7Hp2wv0c8QXB0u4/Flz66PyJmI6SPkjHnHcHtzUur8E
fnVor6gFzItlpqwu99cktnF0WTNCTqTOVBSe9xAZfT5wdRlSexEiFmJMT9o6oPWx4iKorhNbm4mg
YRnWgegZtwTc+yyt49AOhdUzzWbCz52S0/j0plhODQcKg+ZaSw9yAoPH9vPsP7jp0qQ0jCZHHqJr
tk4f92Btvd+/2yNFHI7Z51rPIJNIZjyp/hjKlmwsSrQ3/URf1SJM6Tf1kSbAmcX8RdDiWewVZ4oz
/y7NUyjetokabJnxt3VndEzzJy9rCc6IrUSfvKb2Dh5uzeoK7V1GYbFIRy8oSN7sptkOazn0zEgJ
Mb1sc1BXjpM0wRAYj6tthkI9CssFHU3mGVtNUupZkTOeI36vsByvGr5zFYcuIhCnSEEsqpCJg8yT
exDdevEEBmQJ/87t5N31Hns/IA00AwNneKkNvMaIzMhH0sRIp8RMJOUSCjq3xY02YR6hVnDJ/3vo
Zi1qDlDmOMlCY+70B0KRSQXG9quxhDq1awKgXzgVf6YzeaWE3RMonCDw2oeYms7GqcVEK9Xk7RQ4
mV+Vpz6WXziOAS6ZowDMHsOIHxkFm87WdB10dgj2VHAI1qftnYs86S+cGxTY50+Y4IrWsjS6F3yh
EEnvCwQw3BGS6QpNHnjqJQ03IqOs4IY8kUWSM2PXammC4lw30vRkYU1Le95zRbN7QSOFo3UXvTKr
7EoZd7Yj+s+QJytw7hYa/AQOA4hPlJGdwuwoy9THoeP1EHWUQeyWdjdKjiztIN1Q+X6YOa6Nlzlg
FbkU2HjkzvcQM/hp/NMz9M95NWPz8sBi2AsSx+o03IlFyhLuz7q7DC63GFPUfE3dUsQs4S3OdRE7
GO+mblJ0GTuh9BYOyCOiaTvELQdYEQjvOZ+yjWbd+DD0mI37IcXfZd9HBT3J2CqN0JTvCrlN02wa
2j6NOvFwPS37upCYuQVBIcCCLUKECKoMC96Et7eZNiK69Z3jfsHD2e4FYaLi9J2JU3g2C5mwPdQ2
EDS+UzY4tOEY+ah5r9vXy5S3WH7AWZNMIblOyAQP8a3sTHzAk+5pzcGN6N9i8p30lvryBE+H9Qc5
sDtuDOt/RS09AspHmSwFdglM3RPudRxGo0vXtrBqC8y0kgq4s5kTp+hNnROXE+3U0+MH22OfaOch
mpEl79EnAWNRoFEXsh37iM+EYYxvM3gA/HF9jDZG8xu1WDxO3cskQDfEJ/OUA3I87fVFuSKncDjl
yzJNCN9yIqQN15A2S9GEQTlzyKLWyEZGZLERN8qqg+v4YON4YgvNsC5kB6l81kRpShdFZvukYBmp
7AdK1JUHdreOC8k5lKMVie2eIHDA+1AI2Q15q9XkJGhxRCZcUM2hdsUfzqOL6petNchC3fySyd4L
+bqAIahay3/2+OaW3VGSubgpOBsvJjBcKRSORmCCDP93JJBIpW+Lo5FgFUXpfNOzZtlTXN41sXuL
3WSbWRqmxHAI3ovYWHkUJtab8zbPhifzVAQYL3WUk01VXsiLXhYkj24Yrb5+TD+ZkCa+oJwWBgcV
q7JSExhdAQ0YqcETpj9A799Rh2L66Ra5n9K6JZYPO5NxFC+/AVtWCO5DJZ4dpjhIKdUH4q9lF46m
qMNyL9V6Dss3JcaRIFfgQf/45AnetA3bzCvoZRyu7GsuTsVAuuUt23d2SkfESaF5tQoSX6Cx2Yqr
B5Qwde0Xt/UR+VfXzqAexUaEfmh2dWGByEfmYcaXdE54+PsyaLsQ7l9qCsSRVW8qW78WwoA44s8Z
1ETcKD3aeKPP8i3toJ0+eVDppl48SZ+YtvDlXQqMWMcwmH2ZuQ3BX3LZglJhBCPRtMqWJMddAWjA
hGzfYigB+pSf4TPBL8Wi2vOYodJ2ED9u5jeC16qdUjTuehl0LnFio7mQ9SR/mbTmkcgvYTVT4Ds6
7fEi7grR3PQLU/p2BlG31csaJO6LMQ0bTsy7Sy4Rr4j9seFhteG28ZQ/sE6mB34X8dBt6U2IZDFk
cgxjEKYydsL6fkRGZnqwU+Z7Sg9j+o3far9s7NJjYPQzs3f/PxKrZQ6yNgOx5q2UmGGbXdGptK3n
lsv7NDRELFZD/8KHLznP106rToJTs7cN4nZZNUsclZfJ23Y3DcFQfo1XKSY3Jx8VO58zb50PT8l9
43xRgBTmZu2IF7iYVIIBMuE8ZDoebyPYncM8X1FiFLutQ5UHszfQRLQUT46P09PpCssy3XC0FzbX
I8lljGx1I3GVwWp/XsGVbizoIhfiFWGFV/wdLLobvOIa2PXQ0SkSXP1EBf8MKwEXvawuvGqpmlD2
Fu9kXqu1VtceV1KW6GtsUe5U9n2TLbFM5xc9mtd9EsdQfEBY/mEa7Lt+8zw4iN+LbKq9w6xKmXeX
jYcZUP6WWl35Q8vsPU9uuVKt5olVsDABItBQef08eB2+n81Ur/Qurk0btUxYBLVrSvdMCDs4E0Zw
cy6IqDXAZBEu1MLVvpeFot3xxPUwoG2yq3tgdBhBNC2Ixuh/l7LezFlXGjY5iA7cUjWFaKdg791f
fKSApu7wkf8IjSt5nKP208TcHeTj67raP3lqifzGu4FmwsDPa4CxYkg6uM5KLCxT6FT7gsy7LEhE
8fKa66wvxqPpZS2XZbd/6CRSaR0UbUchndINSVEfAenqRhKG+joBO/RDn+TgUQWpTNFrswM42E5T
WuoPw9g05PrK29Gc/PLI8xqX6IuMq7mLxMbqXGs6FdMPHoN+baz3qVEpMQVhyT0RRLNBNaEmweUl
A7FWuHRYo9L9I7WbEn6j/ABTtNmFgGN/6kZ2TQkezIWeU/z6yg4oc2nL4Ett/3W4T6DDTaIb0ITy
5vhVhL+6GRXwn0lSy1JTj/Sj6dtGgAdqZIBbh0gzRRgs1dElqFqbvO9gzj0M28VBy1k5AEvM1Jvs
pXVaMRnrMuKzIEycfSPbQorngAHoTWLZYUlhRHpp+Cobb3QpcHBZy83Nq58pG74xtPnHWqm+ucJ7
X1vRWUqpTkaPnQub3D+7r8MkySSNZne+nbKziGpVmkNNxIwt/xgP74Dg+sz0caXTl518k3wiIDag
NZkngN0r13xS736AbRbxyOv2CODp+K0DXcYv4wK0hS2yBO/KYryHkl7iQbtqv8ltKFvOaWJ7JOLw
LZPtEKQAZvJTd4FeZ1Iidu5ALkG9LvZcdGAdtgjpu9f4nY02lyBe70BdcINj8pVR7QJTnwJodUwl
NurY/IRUIO8st6SfyuPa2o3o2Soo+eBl287NAcUjhk7qREGEnTcUFq9RnyuFTBf/80ozDHGTekwe
nvsgX1R2C9elR8l1Jgs0ZS3m+ZVmOkcYd0ZMzmeX7ARHJN0eJfnApFoidbPDp3hQE4lLbLl13xGg
NNUSEdynoIb61sZpkbDB50RN555AmTC0OQdeu9ybCftEzXYkIT3t9v8kG7uSzDkhwZx30B9ypOzl
dIRYddsOwzX92QdbIkDgtCmhQ0rWpY5R5a/qCsCwxbhnBFk46OFaLo5gFm0v7vgLviSYDwLKzYm6
MZphNlT3vHC2AaVZatVKMQrSw3zasua+3N3epYgH664BJc9bwED+KSR5QdK4g77zidjfbHyWXosm
EBqkWgZ/Nosz7lxN1midNLDIxn5Hqf0UZRHsg0oUfSWxd63Vfq0gY7jS16b+DoBAABn4IBhIbQCK
eyGRW+88fhHner0XpLJ6A4ADjQLVCstf68rT2+92lQf+VE7zvkmBVAu5/GHYEsMpyhpW0TLYdsA8
EpIr1LXvqQo2iFwDa8I9eBst4a8+U/eKM6Ju2mcnI2a91x7fxmjw5C2BKO2CKQqA4yjR99J8HyVk
OdR/ADUiy7hzXV36y01c8TZkKURYczSfxMCg727aNf7RPD0Fj5PvIhpiKyPH6Z8e9SE2/wp+yGEW
/lewEhso6ZxqAHpMm7vrVEgWrOFeu3WiCUg6e3+yAyXFuRVe6T3CFrwxZ3uAaI8JGZuqkIxtgOez
RKodhgZEYqSt19vsaQLkcmaSTu0gAOGxFf6BBqVaGcPDCl86jJMb4/VDBx2zShy3tBD0Oj4FVHnU
NaQR3yRceM9LKd5vMpGrnLN5Ob3H7pB8+TTWm/BJzlQ56A8CtPbgvPj7Kvu2bKRas+o8NHRVF8bq
jJ0tkf/meMJAKlZ0IKP8nFPEW2GaKqph2QsmiNDiLmQfVNfWvl8hLTzKcIEPa/PC1Q8/abbtU0eO
2nIn6F1qErJy+IfQuJk1/txawq/yRY6B6Hm8NhxqYCE0N5I0dyzthVADjOJQ9NOM36H69irIyo1l
onCdvLV38TV/uEAHNVDXV54A837SDxsTWoWIGOlX2xX9FY9KSrGMqFGxUh2KU+D+pPiJGovSDZzx
oJjl03kc7SsSZPuaA9dHrHqwHKyi0zcCT4OCHueC2TqqH+H+qgN9wLCspCgx8UfVDN7Zt55rLl0O
VXhd7HfpVK4Y9XD+HdaGIvBusQup2K6+89h4BAQupC+1Lesj/JQ7NYMIJPg2TfaJUR89xviBQe5M
yPBnbQSEo9aT/xXzsgMxq4QXqJwyHFVsuVvliMaC4S8hmnF1tyKFjbihKBADPVRatjX9yGu7A1GN
2AAAXtnWGavQokhxn/T8TlS4DnBQbS4fZviN1rDqu0tgR3CUkWt3ipSClVWre78fyZ7uy3P5TQbj
vIaY/DdnTgcr9uQaekkTTslp0NzvltwyhGa/moOoFxqyF5AuBWByjy7MiDtGtHacUlIH8dExGVfU
DB/anIyH6fVvH2Ix/ohN5mjWVeDyaym+Vd5huTO2hfx99WVGNNDhHdj2e0NUjvS/m0jhQwZvFwJj
l5T7WIgjEbJCcm/fUoV97WAEFzkgncQlwbmG5uNJDpDD8JpOP6YL6swS/a8XyJeT2pgQDvEKEytG
1DXqFSX1AXiZde4v+hPKYVYmTMKAohCa14S4E4eZ/KRIjKBlwKTH4ZeZ3Cs3QjIJyEWyybjf4eJJ
HBKGCzbwqSX5qzeeFWJYN6NFzUJWLieL8EFDJ/q1Szs4Q9MzFIhCrsqa9l3KBESm/+MVA9lqTOdc
cB7qBaMch7hHpGpTKz1Ncop5SPQB5gN3iY9TC4glBYmDuLhFAqqPDdmgX/CeqGHRut5EqDmq+vxt
QZ0OtosiJP3PFgnUwws/EzoKG8Pc6Nw6s+JUFtqOy/WP81aV4pi1qnrLW0f2zYO7wF+BBG92vsxX
aM7RiLXD6KcaSgOfojRYl8XtaexBPlD8Z9jqwmxYTcRpcvRdvL0Wcn97/X024ewr3+qQ0ubU6Qti
9qRL6xRZ+zQn6vMjKllNf7Y54qYfSczMf56C6qmEwnvm5EsqpYt9JbNMVQR21+CjhT1qlnP5Hxc/
y86woR+Mnk0rHOi8J3qpynqjLFp23TUnkN6mmFjHdIqkuQK7q2hXWmkCQ0Lxc0CnjOio6HutI601
ivgZPWPHkriPoifHCnarBSb97yJfU3UtCvOPF2XKuu2wyVDssBfHwbYwE4gtF9mkEcQy9UMZ56US
wfBJ/to0BlpQm43hU4+TIYt2EVpixjSMQYMHUJh34PMBzC+YgGfqpCajmqzjN9a1GvrHVtJwroQX
cqOPHf8B2zQVb4qxMbF/sU4Hqkt+VQ4E6kCTGDnrtiQdJnMhqYpJykETu+bdVEdq/JQ6GcjuhZs6
eHKOgpa+IjEhL0xSz3yfK14PRcxQT6UnvnQjCMd2AhYDFYC0o0vRbPZQUnOIAGNmNqRHVhz2R7o7
HB4aiJd5n2+VqnilXq1lXJ1+3VUy1X6/QAGD45p4RfVIN9VPDkGBM945SqrYW9k6+kbQReHQLqwv
CErdH4/+vjQVfzs6AHZWpwkEUJguJMUM48pO2U0A8MJNMYtJPfGcHg/+lf0N2FyWXVqvPzJjQqnD
NOlNk0aY09ylsLpm+0n41v4aS0+nZDCQAcXmyCk6wvBYJ95YKu7v/aP7B98NA96jC2eJUDeglWRQ
7pn/M/v5PdDkS2VC8Z8cRXjug6aBphbhraE5WuVeOFseK4+qvtemBvS1gyJg+ux5YjBrur7fMKYz
sRXRBjCtijMafeG/pGMTqEzlh40RaRvP2RpsI+MIL+xojfMQ+4A8/gr2bJ5DAHhrN/q9B3KBDvA8
gtnfYQYjVMlXGnQrT0zR409N794UG7B/kLKxiSK9YG6mDpdTylJ0KNXWJpCPbr6pdRjzkzZL9i/+
witVwZtv+oxXBD/mo7YE4wySzlwUGulUP0XRgmba1bLRlxmjYPz8FAauSQ9fDeBEhXEoYa8Lv1p0
+wUv3o6ajg7z7kSVEPFntKAOIYGFICvIiQRycrkYoJAzEns+RlfNsmz8uF7LcUlnItKIDIlynlBr
crMSh3te1yoFgJRSIDwqYNOOCFAlRmzWyEcV7PUtiN2KXK3X5V5f/7OKLiTg9wts7IBXoVs3ep+7
6FgopbzLebgkkeQQVirxVyXkwvYmHqurzzhHcxRmhbzkGgWvyhSRQ/tdI4bvnvv9HzW961CihnQM
zd33AkfHyL+5qm+I9zfPIladpDrc7k698yxDheBWdIf+Dk/tMS8MkYVsSsYocbfksVox0stTVqG7
PNc40Man7j6OWwWvDurXPvnBNQHjbRFnkZPGEGkgEiXBYxoqYqENoTBKnqqbqv6S7RD/B/0H+379
BHXE2tCFGV2Lozjo2CFO9Zn8HzqCwa99CYpaqfCypPb5DNfNvC02uEw77jdgyC7fjsKul5romN7+
m+MqaWkRxxX9nAxE69wxvFZlrwER5LtCHcFt14msNFE/LKzIGsZOf313Kjgkb7clz92BAQOHK/o1
hGsEY+xNY0r3svyd2q8xVzXvs3JmdQd8UwfGUCaxW6UQ/ocA+i7yEAYM+dRsmR3sBeB7CJnLKJCn
bzqm9nWat3uTxVgHiFWaHYJ/7JUNDHqOHp4ylYOtsWb8/Aql2TyA/daa6Rn+49luD5XRdVtOsSuN
F6aemiDTEolXiB94fctvu2Uinl+6T3FmsCBfdvR6ypf9YzR5s1NO5muvPuXmUBVhYJua970gDiPY
SPjLz7ivJ8KShD8p/6uezzYWIOamROTxi096+Qoo8IfrOBSElDrFTngOnplutVroq6bFpnCt2XJw
FVbawuM0+PQuJJuGyGDqZmyuiHCQNH/zsqJLmDh7fbiXwDsDPNWIjX+REawZSZLFC6w+aZV0Xaay
DV9zVEWFJ6qK/cV+ByMf8sMcef42DSxoN58sBNkh46t9Ji0Bx0SOa7TcvB5FCRoPA2vsb+7NHq1g
80YcNCVSXGo1HtodzGIlvxA8T9l4enbwe/cyCocxmCiGTaShHiK2zH5zCeJDXSCXkdO02YPEFQbG
7b4ZtAlwo8jSwH5JW4F7pULt3BRUZqYU7cq/9rFNkrNFO3C74rY9QhEg4eynTABhj671/y+VeGZx
rIwgyWBCuzmwUZCibhnD2Ij81/MUkTmzCZPiH3v9tt6Rr6d0nvEkdPnL0rtFP8SmV9vuZSZtsnXB
Ky+RIF0VVq0jwpPdUAnqDDXcigBR1GoYFESClUXj/fKWNGi5xjrYaezQC+VTN8N++lePuD+vM9HG
/hHtQKGEiZeawlbNW1dLn1fib4l05t0Bsn60FYq/w1uVZLn5dGDeGFwtZA1kYIWSmR5Z5bzmsCsd
WEhORNGeCpNAfj7vVC8Ediwv5NwXRbGXWVw9v15l5gNk10e/LIy8KDmbiG278M/GI1R0zGHnUbqF
R9X0yMrnoDgHo4fAtONQRwZsvJDu6/yFhTu3SWDIcsdjOD7pm/BNVGRmFPnYSF3YGAvDpmLBaIAg
1dOSP4x31HbCI9OwQTdWXRld9+x30Klr081PwDxP6YrDFntCJYy6EBmFQUkBWfCHWpcnejFTsvh2
oLwsNKaMj5A3VvRSoRKT1CMVYA2EKmPGMpNAqV8js5s4onxJ+buU4rDAcCo2kBD/TuTkaGNhW3x1
9+CQjQFXNzeSNHvLScL+as4Wf8fuAkn/4haoqXASCFooQFZiBQ+njf1x75rWIJwN8NR8e1llRwo3
vlwNgC+L4eja6eZdTFyVSD8eFD05wdHNi5rLteCS2Zlh3IfyJ8BsY/RGAo8OvpcoPBiqYvu7AGLT
24EExd+6beW3M1l807/3c4/o8k+Mll9qlJgCg9rF7dqcVuI0fLB7lYh861Q6Yn9GVBtOmG8aiYZP
pFJYJ3ZNORnkFlHVa/zHEL90qG5mxI5Fi4siYoTvs9F3Vyu0ihkfPcUuZ3RP6JoRqsdR0IhTgWrg
v+PDbulEyJECLCStRaLRpJciJFQWlPx1KqxKRVu0cqSI1YxKTdX0PlEx8gttgwZp+I6+pn1qQTDA
uVt3as9I4cECFMpVBkJgzBNS5pv48NDEuK3yDbOrIiTOVpN6XTYysjlsgtT500RfLsJ1YGqpFzn7
Mho/MldgiL4Le5obp9a3pzMJv85lw+BdRm4VEUDRC6GIeTNHMKjFFWnrWV/5WOTy/u9COarRQ8ty
+h3w4vxj68z06M219EWqIgwLbQNfHEYbatjrvc7nFGRHwQVCKc0Yr4DNDT9w83sBQ2vJU2bAfNyd
HCLl+MCbrMkVnGTlGz3eMlSs+PPPn14euytbgvOEm0hWo7AEXHPXD6J2lk3XCZB1YZZq7OXA7vmF
eF9aj255alzcP/1h/nzZmmHN5BW51X17wYuUs3qS2gTLlCS/ZwwM1We3OH8qUiHGGaIc+IhlO6CR
4AFXTyIh3RKQ/T6r6kG60t721i29+G8nqa5ou7fFpkT8p6mc2799zF6Ltph56mLroi0Ps2/hbYRY
/Hjw8rqJkc7qbOKwxghs51tQpSFY8P4Of5SIVEMtpBWhDA+9+qnIOZ0lE1KSuxwolyAJFtOIUQqN
6/aZzqcZq0nqxJWLO6IN2VbHlpaIFDCPb7wVuGNn4KEEeuTl9Z/3KKrdtB282SskghHMTKMcCtyL
eJEVEHaFmkLqxfw4ET2uGZkItjeNa7ULUkmaVj81Q836dUWulqMna2coHqZMApE1lvj4wlf+0o/H
J7Bqm3UkqMtQ1Odw8j4T7S2Zcbr83TbbVHs2ebte8t2LxP1sUACL3ZkSAPAdatIDZY8r2JlQbVx7
JPTgZlToj51gi97pRnTigZQQg8k7ZemR1k4rzWsWwC9D/uN34512Db+gUN0iW9yl9FhwOfSlmtGe
rgcUcAUxN62V2eYexcss5eR/9gXbgoatW1lQzfnIUxGFKGFW7z86+j4l4f1NWWSvqyO0aAijGVF8
zACSUr80gK2ze4NhneSpIHUF8XoYLyWfjKvpri6WLRdUwuv0FcAb62+4EtmVnCn6b9rchihx4iUv
VJjZVjSPqgqmsnVDQ/U+nqI3tUDBqV8pxtAtm5JPd0djE42hMokx05DO57BN7XVRhkWYqsX4cnc5
tc7rWGK/HBwTxoxMSy1y1QvUH+jbN9feIrhWE/OvQ4INdvKO+Cs3p1hRBK2Rap9nbZBftMKHnslY
W8HQnY/T99IuWBJ9Flj/WLIBRca5f1vkQVKzyZjP1n6Lf4QGcCzYxg5sTqnKRDUkUQ6ec+isuvpp
IaekMFaM4wNZ0ggeL9bsH7VObw5S1uYhJBw3ep6I1SMAudXfynylFxUE94uyCt3wlrC9zSDg9YfF
lntABf8CdV/51mpMUFfamFdQcFMz6DJUj+RPj1rkXoHrJwL0soTi4OWuu9kTAsQLUHTD3fD1NEEh
yvX4/dsJ0n11NJgUEBqR/051ZUv3RbQ10iQTTmNMX4R6pC7S9HMbWolMDP2FZCAECY26GiFx415Y
sGbR80RFfn6MZ5V0+3LoYk1dw06IcPSwx8MSbCp5sHG+pxeIQAZfn+P+cW5jtVOyg7vP3XN6bCJy
oUmjLbLy+TlskGDEL+ZpuCAlThnHJq4O9cEBDScZqjgLey05oTv1dxu7qOI8aZcz7lyhRYL2d/sV
ewSnSLmHxGvy6Q4f+jtLRf9Szd9FRLOPUDRS6RCdPexym+I0LX/T9EwwryRwRGmfnnMWsDa7qzHS
8KCXjYiN0np+Yx01QnNVU2iASUuxolMs7pNUh0fRm4PDWBCrEpXnjhQhPd2IGKHYbDiilmWNZfKK
Mcrd2VSzzKLshr5rQXESxMbZ0neJ6LyExlh2X8a31l9oKoDuL2JF1MzcHQFdWMP2CqNDYTOmaGC9
MzRDmim46W5BmPqcTYXFJkdShrzYo8Id2S+u6bMyDiGNUy68Y4hLr/z6Sid7HO1VjLyCvzRN8/Wa
ZDcAbGUGCLquaSH2/UAXSb14DvqTj0fCskLdK+2MZ9ebcU57qoYtdQEmoCk/x0BmtBzT9KeYPyvh
O4m7o1aH55H4AF+jpQM1KKnk7IoQrH25nHxAWENhBQ78TUdtGOH0utBdo4TF3OLeDI/3RiNBmoUv
MMhpBKIx2RIimViYDC5HbwOrzw5SF4Q4ZWkvPSPT9lGtRnKzyM51jZL2IhXLHnGMtY4Cpmojc7KK
lIOUeYl4T3qmh1ZbC+x1dlDbHsf/rObk5R4VEh16MG1UV7sKh6GPrk3TmgbL4MR86eCQ9oRIKc/v
3XzdmXqEQs6b43jB1ve6FvWrq43qf2KvOkR6dUUYFpmDkGOeH+8c35ku9F3Yle10VjKkoT6EpdLJ
eFi8Bh8G2d9vxwHKXVVFVFGXrh2EV71PIMSGxJE2BlhHtiRWenkrphz9LLXmwsuLUNEZIktJDsPz
fxF15ORPUc+u9CCf+s1Sn/7Ym2C2tJGbEPfMUP2SrLvmeaE0GY6Q6qTChmzwFvNNEXy7bXFLsYeZ
H6DliclvVJQI/9pw2Aq1pXtshRf+v7lKImJ3x5VkkNt2fL57UNeXlbwhwvK/aImPalVxVImtsita
hN00qBNRM05hJp4VHvqqtJIQDa7RLW3T7LX7Wz8HjOlGcZ53UKThkZj7/BCD3HRLLGceHI7Alnf8
q1NJRc+rN8G2vG2rKBEVEIjKcddSVrdWIL+0Y5lkJaQPlI2Zoz4KRJgIiGgqllAq1FKaTyavwl9d
QVNXrmmiglyTq12/TmmwZ2+UX6lYF18ChHN4kRDmz+e/Eej2o+2SOrMuzZfwZtOIh2yhHZoUVBiu
Wvzi+mVeM6imLsZsNsYozaYWXnAn3Ydjn2d4K/GveUEoDH9GLn7sWYDQkeGCuyiiXIlaTYKM9q0b
TY1sFaU+MDzt96imfrn1MiBfJBn+bnhVLmgHcxBDcAcsuhKdw+NdftiphSlHHEBuW/v/fNWBXNEc
Il6oPRN6ZENlfn2XwsYHp68uJ9wUoGt35lOZZNzJPPkxZp+6FUIQ1xFskDxKNF/WbRdfVkZ1wUua
1YuuY5pweU8J3N432trHFZ/3zsu0BCQbX00e6CftBchafASaGWy+vXl4rxW/I6C06vLCiaNoTHrq
rhbv7qNcNHM+xxe+YmKiEY0A0oW3e5ZXzMjzkxiRBVrv/E/h1BoHj4QzyCcH3HkSU9bkK29Y8fDc
RKNWcgQivc+twnbt3eyGzevpSOOUTn7yUaBnDF5Dqz0r1ZnosueXrG+jAfcA5IxD5GCEzunSvTgw
/t3SlqMkQCEF3t6TwQPHt9RtAOOlBmnuC2fUgzlHekeJd2xnqEDyktnvq9d4sx09XGKXOB9/aHOG
+K67rFX+TZKr9VV4/zRVPsaIrMoF+1UVr3AVWTLG+sU1tqEEluNaSwjNtY89r1xc7PFN4b/jSKJu
sRXYtrOlD9XFaCn5LRFoRny3T3Dw74pLXcVg89Gjdg/tc4+Isi9x3VOvU2KL5QXVEAzi+i2dO4UC
lOe3s8n1nrYPsvoH0J8aE3napUNW+pGO1GupJcd5kOFKpx5jWRGv4snbCLJ4Kk38t1xui1USP4xQ
cayCaygMHAtzn6lSMi/ajxfJy/UGh6iEFs56m01pyf1NfsdMoJNtBGIx0WecdYSeyY9kfSqLI2ue
jRA3ogh92ww1owKfaXSaYc5KHbdnlfhQZ8s1OZMwpKLUsjlTkSz074lakOQ8PpoyyAr+ID007l+Z
0gMCvVziSjk4YijRZiMjITgsoNZO8sboN50K+X0KSrGRiljUwzklROAwN9EGpiYCd8JRNsjXYztY
5FEg2oQd5gbV/D45XZmnsTnr3/Bj2vEEzcmg7yCvOhy/bwcc1FM+DzNUpuPuwBQYF5CDlQRvdO4/
8vS4Bt2dpCVgMLe4opZKd1W0nO/3lLcyrUS8n7V0b0E2aLxXUTzEdgfl7niwwk3Rb7pzvYNbDXiE
qDZqcIXx11RtrRQDYBs5kVkbzh5XYGsoF7Lzug+47zwkyGNUOvXWr6LWXGIsjftXySW2/J6SjIyr
fTMUcAni26TA1UlNVCL8j9Rjol5pdsP+pNMUz+O9gaj+VzcCP6bWsu5/oP/2RyVLjvbt0q5CGjnF
naiu9Svu56ajdSlArTX4c408mkRrvo9gvq1ja96fB+STJFc4xmTXkqnxf+iwBU1IRdVZBx8AvQDg
RKK4x/TGC1Vpea2Ki54x2GRyI8SkoFON0OVT3bOb2nhzy2hIhcqiYc0mIna9zrwwiXG2MSR1SVtY
x8Q5QdBZ+jkuqvQj7r0qdNu8RtYCcAw7ve6va+UoHe9DIBueddnCoyc4aVFq0l/8Woa2/TcYwiaT
d568TOJVnVx2KI6dpzi1haKwLVVGRLNQRDw/Y3uBleFa+X/f1S6TyOq6tF/5ou33KRR0n9AXb/Kl
JQXQAVQGiGfHXDsPZj/hl/qDcpmqnFVM7s80d7yCQgFREND+fu+oGejAGN/oZvRvERzE75gEmq7W
Jkfyn88u9sIW1zZzrWaAon7vSQMR9MyywvUoabunXdjkYDlUbkuCSM0hDgoPkEQVEyuCppxWCsXk
29XoIebDFoSHMtp8PJXn8wPVWVwfvn+ulfyHTYSJ3JaNaF6uWme5duB8luN/22Vc3C/04QMfuKZU
hqMlUhflZVw2z06n9SE1fsYw3YxkCk0XXB61Q2qWMdADnhJwRxyY7ORNkhPEfCsDEfrr9JuU2zhl
LlM4pYpBRFOgXreXUIWxtQ7N82sCsUSMrwx4Ky/bFJyuFx5u5mo/hJ3KJdweV0oY3yu7+gTHRBwy
KEi3N/U/xwanYTTOxHHkWetawKmKTGwlw5kimk3KdWlYMvUa1sQxCZ/E2niJT8wCAq4I+Vw7enQW
tgDzxhqi8oaqUqOtW/sXKbEX8ZScrssYVqm2L+vd2bBKIP7i+7jH6Fd1H4iaV17hJzQL/Ra7DoWH
l1u2TwwzIIncMclmLLMT7EGT9o4Uj10iTZfSXC5tT258fGs+hMM9/4mqaRH/2NlEyCh6ZdlRts2f
sJBvWQotKKrtDMa89YSXBYq8Gz6yq96wdWvU8ttoVxhsg83WFjl+BE+7EEZOWPSJGh2sRJ9ZWOBc
sn/Dxw/0xvmi6OY/RNddXfRGYkzqzF0gR4ehWeXb+nzXrvlRRH1iENX94E7eKGF2Xx1S6F0GrqDo
f7Nsn6Lm+Dtuo8KU4RRzVldyf1qY5zDDqLiP4eTLuU8nFJj125fn/sH9T3RYjEol4xx4Hrp/t6yK
GPTx0BFfFQPoaTRiSteb5ZucRBqAzsDEF225KD4I5QitGWOHbDeCvtPy6B2+0J7LHyvbexnAoDQt
qf79DHNQ3HPxoPZZuVjtI2pcL/U1PP0VQeJm2ZF5u6fIVNIbDiTH3eBWZDe/mYjG/atVt3sGXfL0
D5Eg7aW4ekoe/huL2pMAy5WbAVn+P+AOTVHmOb1YNF21k1q8VjifHN7HVq0yri7FIrEyh7PyMppn
HoQrF5TAl3RSkanjZq0nw71QrLORiFQXzufl4HNkK6iMKL0zQGQ8aLOJBjH62sTawU9mO/DBBAIf
xbSEvz3Xx+T0c1GQ2qgcciauNpPTQFPQbO0QN7BtHGSfWyaeuc99MM3QZRqQ6EvJ+BdR4NyFQiA4
GGwwydNeKBR5BNjlIA48LevOA6Dmjx0v4lL43Wx8TnimOyLwBmHJclOM50UAoV0teR68UaMRvYNc
9d2CV5MAeCr0VuezLtrxqDE07puHeCld0+ZK8qDXcFvpfgHU4PMPq/kWc56nNnw0vR/uUY0Udwdx
YUG9EiqqMWs5b2pkfs0DW1w6l8bAMY6ItWP4qnUycpVbvnMlXKG4R23yK6k+Ox8TeKB/9/cOYYYw
Ioe1EqFjR+fgywFBXUcC5baAvnJxi6PYYnkI10Hqj+Pf6JB6yFHm6bfdCX461OdFTUbE9JUaf63w
6j213s/QrcwOu8Uui8ESFhYxbtjsWgCtE48lq0xx0tAhQl8LRdDHDfdewmvk7msELt1Bn4yDtbXF
pY0TxHKUBBgiNhLsjVGp/g5G1/HuwTut+s3fO/II4vkkdYxJoazVoz/Tvr9ByZMxh4L1loEjh9Hz
mxNKv2Pwt6e7zfM62swWqhWV0nyWLEIYBvo0anTzvGDcYYZGQxTWSe6257762h5WAX1yHHZHiaR1
AMpZj/NzrkDmpJqZwZI3mjdN6dOSAYG5rtoOfjvgKEMcbFAsAAqEnHy5wmJJ2Z+stFxnMuNBEtBd
rE5tOWc7XFINhI/DcW9mr00HjVd1pBrYk5wMXcCcpnNMp5Vn4b6OhnhCiKbYUV00PeLxwZIJs1I/
UKmgwgNG+A4JIt+Mza1HoX0LNzIBBKIM8I+h0691lKxswrnIB2wBsBJEtjwClMeNU1ji3TWiNk/i
q2EMoAu1exRntf2PB0j9SYVy+A2j/QtiV7STuknWx+tltGX/a/5aOrWfiSBJ3hZEPm0TYJ2jdJ+e
74k5+KYRMjKGqUH/zcweAFiMDITx+VjTtn913YTVa9R5fYH87CMxBnhHymsVXNB9WuFwpLsaKYak
h6ei12HNSVNrIYmUYDe/8ChIfXPpvD3UfA7W8DGAbG0YMlOCdfysvXfnhP+9xxO44psUldokTE0q
rZa9CydrBH6WP6D4B6MKfcUjChrrClczwaSFbwNSHbtCiAQ+O0RrWQaKFhiUeUdwRaylViWR3i9k
g7wmoeXpDn9d7i4C968VxBfWPHSD+fCECXnlHgP3kY5KQ3B/SQRZ6+zfGLQJ02E6hYkxV+EGpMZY
r0soQRD/sno9STczNyriSXu/amx9QQdoymgKcoglB/Tk+MZEMZzOoY1rnWh3A/1lcqm6xS3PoJR3
MDI40VCtb/LMx6+3SYt0Zxs6cHOKzvzZmbHO8M2UjS6KAKJSplzlkJEW5jlDRcUubW3A7nWEr0Gq
67TVDqt19ohL41qsw0R80QCjfRpnEQC5gVuEZuGsF75YuJxquzfdjQh5cQo0+wgV2YgPp6NbFb4c
KH76/+zfK7LxDJNXOEb8I7XOmuChvOum156emprOtBv2/ejQrrWrzKEYetDmr9lsUlbKiIRDvYur
2vm64K9LW5VWFjr40wdfdkL5qCVKWXX5WFZMmPtmlA2x6m+pwigopw+Iv2QVvr9lCLVK/iWWIDrf
fN1ZrWTsB/HNf/XJMqwfXpNIYM9o1VsG/Sl0PyBuxusz+q/CjuvPz8MCUro3hun1c4YZ4XfJ/lnd
ms4jJgnSx+/gLjjRzzhTJWwVus9MTBXn15FScTbqWIuelIwXkS/SMHahvpB5OnnblGTFgmVj8EyP
38M5amyyQk4PxQuWfw/14+3lp8hZHxilKjyYaPOkVvswoXECAgFhjuULvTUiofYqVNoAaAnCE3ab
0zrJnzuOF0lCefRdlfescxbdGBKE10ms+YARSlQm12vYK+ajiUjEMBX8PgsHfeq4XlkPi4ibElFq
m3j7ywueCzRNl0IGvlvHrNFySW/e8OKveYWb6oTAwegQH4caH6I0Qe79Dna9ThLIiO8uaKXZcMt7
2S2tBZUVKWDeSqKOg/ohmNW9nA00RUkwJy689IsaZ6tvzLI3jSgfQD3ctm1u5EhDEMJR6zw8v51N
mWs5/Sn6hch7HhB02kmz8ITcXUi7nFNshWiIzmwIThnZP+uLQgn7OqgC/KFcLJatLNing7cILLtA
6tDCqDXtTWgXBPYox/9yBaFiN/Hn0Im6H7vQNw6DvN32pOqVm0bBWuufeV5y38qPtXc+ob4sBEU4
Dc/btVBWt+xaJCWwWfTxfO8zxQC1WRq+mmkiYmvImMn3g3Jb1PKnNoOLBtAAeF0B2m5q4QXci8hc
fouCKovUHYU/ijOJyVljnFcXTX3sra1s3laMJkBPdVD4UIPwYU6FyxyrB2zsUNImkLsU50leAKaY
a8XIxxWB5BEhJai8ynzr6gUsrKb7g/VqQD3bCKSwcJUiAgPtCPxtds9qum1UHs4StcW6dJwJw48V
rtQDMgH0nzVMv0zO2M6jzyAaNn/R8Leus1NUwTCrmRzCv7sxjbaXi/yEtHnRm3BalniS5TCsoHAz
BmHY0YBm2C24qwD1IY7PKJQu3c3byoh4ysg16uNDVQvGVri9CXPv5Zx/xpcOZY3kQHHHCA3POM+a
wsEYkfyAMt07Rch1oMXBkTooL9pjFfpdQOfBTJVNl0dlPhc7vJoD8HUTyPzS6bVAd6Wb+/us8/SF
GaDLrJq7yWi1lysrJzf9J7WPGkvV1WoYbtz8C88SJnvn+pZbY3Lpwm5ydp8yy/XKxmm9Z44+izNp
QpnD+YFIstS6GWX18sKvtEucvmHlkxwRB7CyFIjaZDZ+so4Ih7mF+Zu06RNzZ3rIKie2CNp+K9+s
G9AxGp1W1V9K7kbzADvNRM+b3KG4u/P53Qc/stgn803Fkj7NwnyBFuYmrVUZA472qJTOlrNnwmNd
ScguLF3R/dLserfOBI5KwtXdo4L5QWsF6ogqUvE+K0TVQ5PlRH+X70e+XguZKVzIC/pQpFVpNwn/
QLNWW0kQK30qzqKUy6lHCWJ/IpH3+KMaTsl0HWJDrLZ3a+wIjDHVpB3oItOh4OmWT1Vd2ysCuOvB
YXBVIPO/huWKyT0XJ8eEjBN4UauuAz9ib0OC9i1MWe5oDUVjqzdJ6Gyuew/92IpWV7ORjkIR1EkS
6oYY8giNAmGR5V5NVSTzkA9U5FpDQOHtTezzQ1VjFxb0/FIzWIW3wX28G43WQPbnoAQJmVc46Fd1
DFy/OSQyIamtbXnnmgtHLCzmx22m0BS7P7v+7lhZbyhSjWaIbOjcHKqajkdCoGXRr+aZYt2vvYho
pA2qNmN99hb0rg5x/4yo50o97YCfX5dEVHeTiEO0IP8/NNpu4tl0k8Vv6sbxSNvVYD6qy/PiOWBj
1CQ7xFIE08jVOc4D2jfQ8RuU1gU4sZC01YEgYDbpikfy62tgorErv8yR1p5MaMsp+kA/2a+FehIp
9IimUTYjAQ1at98nTmyqxGNLn7B3b+w4ucuWNG/guOBq+LEVL8BMGpg+7Xowx6BY+ntV4UUV4TpX
yAovdP06xD7ZNqmOUj6t9oZVl1cmP3v63ovuPHVacpFtKzc3/zMHEqkoF+gPldUJ1csH/vVbQOXy
LZwEvH1eiKkFowEuLoUqtfKrA3PDN8D4pOyn7HD5GRGkTc9bXhWr5npmMZCVLBOY+EX9hOStj0Xp
JfLfptLdzFoaFf3MIeRE/X/Qpc1i2guOi48fJOxozXzpEWh6J9w4+iVb4xHo0TeQvBaXb2LET3XB
Dv9tWmGZuVKugtWbIkoI8hu/CgdZa+5xLYC3IWkug2vMFpaufbYLMc0lFhX6eBmFsPrC4a/HiVFP
fPziibxr3lMe6Y9kNL5owG4gxwVfvBgsjWaq3WH+Rn6WAIYJT5z7nvpdoM2BhN7PkF0teW7Y6erY
+g2md4fDHn6LpTcyxLVTnn++QN1+pGxIvLQ74lXc/DV0mjYAinYbNFpN88HJjTARei8brDbY6s9a
//atvYW9pl130gYJrcnLM1YUw7YlnhhJxIBsJusS21jrTi1wr6P+lF2qyEEeovTT0mZRUfm4zD5I
EF9IkxKYs941Bs1drU5q4fhE0vSOPMLtamKaIv6k0b24AEH+T5wA6tgX5I14JNncv8Xx6yFiJ5AP
DBwoDutMpgKxINxvyStrgnEGMEp4EnTHApZbFMRJ0fonxZesekQj8CeLC/FnRQPaUp6UouLs07re
PHmpydAt64E3jw2ald1k8VK7u9+RDSUqFIOyKYOtrbkrIqZWiPyHXbAQRuhDuu5uEU7hJZkGyYCU
ndqUyav0oc/+dtT/u5qCsDOp21tVtXE+IHH8a0O5PigYOOVu9u5YuuK1KD7K3x8UZjVKvX8oE7ln
JpbL137HPuuEuv/rhYj4bmgjzz+30q3hliU88x94EUPwqryfXCkVytD2BBOfZjFrXTo3JktcxtbH
Ju4eZDWOQV1K82GI4hQSmiuushFQc/Kj+o/kp3quPkSy5fko5juD1lgQYb6wp7QVbxbJp3HXSIss
cQ8WtnItcLJ+pdxQ5+YA22mGDvd7+FBspNK0jGkF1b4fW58RlATEQ3u0OaDXomZAv1qe85XRnET1
q8KaQo54a0aiaaU3zle1E2Id+inpOYtfYGmviKAInP12uHxq1cgwzzFHJOaXPm0gsU1vOXHfxcIt
3JtmyaVrAb85hu7mjLwUv5g/e8p051DE552U0HGhT516/qROFyy7OepQHzVmZOdOih4RZj5nktW6
L3I7oOiRFvVFjJMHua9VmL3CRpn2gfpZSVpZdyl5jhg48FGqFcMTgQNWF4CfLVOT9A25BLL5sifE
kwpor83q/u0TXWPQtIQ2U2vJuPt4hhZoWWv2FfzY1Sa/l129cxNV1NN1ffK+omG7EPGAai8kGUYH
P6JcyHYMB+UwzCXAQZy4DdEchBiXsgyDxuPj0kEmkEKsHTYE6qTedGNG2qEZ9nACF0MyeQ/Rffl8
kvO3EvpXU4tLWEAL97heW/p5w57cUxaoLwKBFvV9c2WJa6j6QKCY3ze3QwURbKXU73iRcYMjTNtQ
GPDqR3JRjzNi261WMbEha3iDnxZ9prdv/Vkl6Lalhgz0JJk+xMJ4Hbe3CtVrbtzzw+pA5cx3vrpw
3lqgj7QCOwHcOD6bJqGKakgs3sSzudxVmI+j/V6A7TXTwK8a0b1HWt5L81J+QDVQTSG5naFaaKkW
4xOwjh5B8iJDMQ/5YR3K/t2g3Dj34f6Z33UV7weO92480SuhDucgojwEbqH7r1Qyodz2YjtgO3FK
l1NjA4/AoGJcL/xk8zPGLoTDIxp4ZIkvoGYQtUxNiBa8GTDpY5eYBK9HhsOxs30SrZazc4vTwvjQ
61DYQq3HON+n6haFpt1QaIuPCt6jFZG693pnpc6jUA5uuCtYwCrrSM8ttdi+cqq6WtsS5gSRHtcl
rvLk33s0sSXJxWfUK0KPmWgSa1pvyNZ5aUlvk9nCXxzMU0nyimeF5YEdvjtJ7rYhswD+uKU+Em0L
3DLA5Oa2jCUqJQ0lViGbXo9p5fe9Rlj1YU5vkvJElzjYSmss0IpTVj6LAppJfogdu4987UlQHijo
txbu9lIRrZDSdb8RM0FbD2fy5D69uPVJb5yiCzvG0HTO9wzxnV8PflW3GFXpgsN57+sjzjnhvwct
Of4za27uC4tfUBfGOVFPVYNL9f0IbNRbezlrbm83aHllZ1jdEUFYanCHpNJQ0QcqNqRnYt6QlQQ3
phQrTNbr6MfbRNdGivfS/reV7fx1GXdWPoNUZUDk9AMuFrBu3EoKhh2kxUq3gWdDiDCGDNjaoXxf
ICdB6W+h1BZTVSGPA+9P96x1tNfFH14Lcf1kLgOSf13ipCv8zDrs4fY9bDk0oRm0cjQ7ceP9Fgvj
DRlhum0q+rvyW34kmltNC2vCJqdUKb8cna+Xdo/XXYgJL7ADgUROIaQVRSnCezSiPLN82SpLPRNr
IcXymdpWUUUSrhtVpjsTWN8AE+uLNbsg82W9C/ymzal9WFUp5vnH+3GExXHXuPWlTRNAp3fztUlI
sfXf/1CBCxfFmwx49jacR0a/LZIADG8n3NxHqoG8yoe5UgYU6s5cxGA21Vz9VQeg2/FCIeya8ymy
MHSNu1omIJ1GI0vT5pkv0oogmGcP2ZJQQ/1Nm3tXAUcbcZP3z+tH8hmM+wPKCpnx0lR0WFeXIIQv
G+1z4BHXlFh0gUJP6qXHJi2m9iwCrxXlyRokHSVdu70r2pUKOQ1OsjB9yu9iFbnfqEoCRkPM5rvp
L2SiAklEiWzVoaatE9BkxiIBvJn4/xJMqm3JfAXUubmsmX/xnTqW9e8gPcKPEKRBnOmxmSTYUFrv
3yOnV2twvPNcItQpo0Hhvkc2qTTB9NU6UtbodZtrIxuya+C7a7py9xXJCmUk+GohKCU+CDZOjJFu
t/LLDuN+x2c6GBliAcpGFX9yAijuYC7MWQLGCn1VEqGElgkdPZLWVc/FCsfOO2UhmaMP/XDAfna2
TEUhp9T7L90AQH30gGfocAa2drqMGvM4AL9dAMHdD4j3Rej0GZI19rCOhtW9rf7QHTJ5Wz7+OU6L
ZV6/PCXZDVp0uwvAGXhfKjOmvWwfTI9eS/YvdcW8uHJz3szvKQ1J18vzsY8sI601Ww91sD9F/yKQ
VJrfJQne2Vx8z9hg5jjKV4HVyRprCqFvm+wmvZc4lACOQIkMceUDm5FSPPc3SqKHk/duZIhnpbfc
AbgFzo0XrYgDISM7nqCIWU1ROTFEerpJdiDfE11a9eAkD7TM8v7nBCWWIPE9cYeybvQJk+3wiA1V
ASf8My6S8HRdNt/NcyhmbI0FjwDyvxvMCqFvbw7P50Q77jQJMPx0RTNzj4giyE28R7Cb+EiOKzIr
v3Bn7doYlPjjN5Fe6DwXeE3sb1WxaAm4i9DRQOutMVkvXBg4Ivow8nvkJ+OcQlkCJZnKp/jVQxD3
a3tUYOK2WcwIEjTpO4i3cwfcZ1U1+bfOCH+LJKXjQbvBV/xGdCN8RP4h4GKjBC/hggUsz23jezIQ
wYTqSxxjXKMII9L2i7/JsAfdCEDXPblkMKIvjlPr7z09aOE0PHsy8jS//aKo5jDSZMCfRQgNZ9H4
TMGJTyPjS1r85Q5xGqCk8pzbG2TjtjT/qSOzRyc16FspjJE9qbjBkGPj2awq4ieb7unssjQPCV/c
nheN3ueshgGquW3PN6lyqAOJyjAy7CBzHD3cn38EnAQypmkdV0ntdSHlHLnHWfk2k8Qqr0uRoVLx
cxF+vkxtAC5L8PTDWj4Vh+FGViLwEC2y5H+TJFOZww0J6QPN9HKj1i4nhUejSP+izC0bUOUUwFBi
8DAOFotdViDJBDEh/LtNvtC4d3AZxRoZgETJ10V63EQw9XxhAk+5wgaury6ZuUcrZP9/OH9nNcLJ
wdll7ZnmVH+/fEpBelQP/q2mn4yJRcOQOZd9Vgk+bT03abKco+MYmkj7LXEEA+1ZelXXwKwvAPAK
E2OOtzR+IG3IoXhpgOCK4K6ws5jthWy3uXIHj6w/VeZAyO3DdywABkHBYYIBacklYxRevlxSMi/O
yKKNj5ym8imMovtO54wFt7JzMkB/VSazhtv1+fSBGnK0ahVE4kafMZsTnxkLkN64hoz4uq4gX0Je
ZlVnMwpaO55kgtJKywOGToWdP+w/bD2TBNy9FMdjQERXrVPp4VSd1e1PRs/MqxenJC1GZUDVAnKu
LWPffEEMjRABOyfRJmdbWH7AWxZEHX2BvVAQNS7TvQJ1LsZwJu7mfKFtfeZ8H7aS33AQ6q8tfdrD
0vFpPyEnzs2cM31bh3cB88WBxvYdviIyfnFzAyDVjYVDjWzmsf80Eq6g3Ps/SrmjtsKkeAqGfnvs
vlzk7QuymEQsxKkL4mjXeMcaA2fHZZz8O+DTRimuhtoxJy2EF7sxZzZy/nokS2e8vDMKJiDPK5BP
F+ttFAkgBVd1v3/j5Z1Qia+bhCglxBxwGDCZ+jZOxwjiFXUl8BLElKylmPOZ2s9DVXoX+LVn4MNu
jOhcMiAPjr3avnEWJimr1UZkfsKC+jrAYqttDz9/YMDi3CYyIywzRc8/EkLliY103A6BqQX5I2t4
X3/+ixbMR79zA4mFI4Y2GqMFYFzQSU/EZqIs7xn6nMnDsLEALnH6qm30enpxBhpLop2ZiOjERNH/
PolOlPcCDN4KPX03p3CRBnCNvz/6AnWQfygubs6Z+VS4WRpyOWAVRh2zjYeJQHfDWoaoC+Nlr9AL
ZzmJnpCoRiai6na3gWhz7ugnzidDwfka0oePKqhVK9z95SdGMogsbF1+NCO4znP/f4vd5DUAvskW
BHtXOr7NexXwAdjMgk6YC8v5e7cZApPrnGwwGQGXfamFsiwBfnMF0r41I/o64iHX95XsWpGTbC0X
tHlwn3oZZiG1bJUPNoM+yvPfROJyYd+60TL9PBAoyUuDytqRpZxB+B5x0CwvwAfd6i3mFuhUoGHX
J2rJIaYNrak4NramHKYy/LvlUvGZSHa1CLGID2WFQXECZES4f8dLPe+zwIctp1Y2ONE9E4rogp8D
ekBketzjQ0CKpg2UZGdX5YJks5BP0CT4LYgLnTsaMccG4UYDJTP5upLvvHNNHn7uHYd8FehMJgO9
o/3XGVG40Wu94kKoU1PPi+TRRBPYYrCOsFSi4MU/FR3jpbiC9rr09XwRKZgDWA21t4fiafCgr4Fc
oOQwrkprUYy3Xkivj0SuN9dFQW+PioHQ4EDjQ2XtvL2YVn/U60FfR/Xs/pX7AM5aB/0t/NVy+jDZ
gGyj0yrMxAzTy3FLjadk12JiQ0ubIoN3l+KmPrizr+B8/2pzz1i1vBdd8LIGnmf93Gr8MknDlWzP
fS4k5Za1JaneH4kT8V9IEsAp1pqVSj1Jmr6ROfEs28ZSyw9UXbEdHXKqQA5Yy2FBmZ/sS3iCBvi9
D3ZH5qZXbWuj4H1TmbvLEFGfoKEbN2YDKacIvGCAh8r7kmw4b3YAUDakYouMl36iuOt+aTLGoaOy
YMEAkCzPZ0CAcCvgtvP74+X7xAe5CBtutoHz4/s89xoVfEIapPAPOnwmD0rc5dXR9x/EG+FRdBCC
gWGAqrhpHkL7axmBS7u4WXMYXJCtGwTIj5TXpzUjx2tHokI7ENCh3r2Pjej6LUJ3+0erDz2/VaMr
0SlNeHwGMYhiPhrnRKkwfKmNw/XHgCVxr2V0VXVikTBXItbTyhlIYbPB7tRteNl27qerycqMJgf0
6l45H3Dugov4gEO0jeaCBJjYZJWTN9r20yo2D+Xa3uO8+saxIZNrc8XTNKCTvpzqAquhuOXjNe++
yJDSk3YnVhy1WkKbNj5OhLEiIK1YuSc3hzvKeiKUg5cTEvhqRnNO+mVMFuQcDQAmrHvyyqxABp81
uID34BdM7a1bNMQ1zMJ0N2T6o8CVNqSFu6W2qpyGoU3fELnnga7HrG1aiiYYOsOidj4JdebP7fh1
0Yk0cLQIT9i4TOo2JZuLyBugALN+joMGjmYk5b9oP1Ftyc0zP4qcQBITSutkKZsksqMKaDGg+c+o
pqoLWZNh2hfkLTg1ERizxJ3l8FJeXAjrO2J53HwuU1SYjK452Y3z8ijlKFdGfqa2X+KrMvL2x6O9
+GLAx9Nb60qAR2eVARHLYKcxbW7EyVLcYppV4q/XXmuwxYErkmpAcp25/5wiZg8m/TxC6UKzugPA
Gp5jtkwnM57cchqhuZXVNIKCLrMMgNYDBGRhBlKwdld+UWpoxcLGxRU5jQe2V8OHpscq1sEKRdWI
ub6oWsFMVLOYKs5aljZKLXOSWWSPjSvmOA/L0ci2FCg3YdD/jc2srkJ5uShEAAs0btgM54HHh4mh
BT7Jcz31jGQ2QDq5Jw+6a5QZrxcO3houJn/T4XxQ0DMh+BDO1qA1P/hNDxJRLSJ0T6T4aV8Oy4ww
cz21eqhK8AecE4s4Y7E6OHXmZxvcsQbaE2LdRoO3tzOBdd9sfXqmRE89NDKscYym8S3NJ8ygLSW6
qPnDzEn8HvI5LLiVHAJV2OmUiUIwGCBWCC3rdTBb8G/FfLba+/pHK7K9fx/gYjTpP28Dym9pyQ/C
BAsYuVAR/TRVEq4Orlw4+JhWzLBFWOuLcaIUYGkf7NFRjC/cA7DVpM8tVyhu+gD24hDmc8sgC8MU
gNaFui7ckbC3oOuOHVoyvOmFIKwkMNj45xDKY8BEC4caIcgflM8NwrS9TQ3Cj/+rpV4j7nHCSW2S
hsxq1nx3yeyi3WzyUi/D+AFR2SnBwaRndyAMZejn2vyKy2WNvYpk84QkDz3Tlqn+YPpSar4EM0ws
Z2YLry0BfWKmhFEkjJ8sTRD/pfALsOSfrDGzoOdgFwYrOSNPlVOqjSJoo1/dqQeH7D49IVxCXoMf
LWkSFd1igRnX63GET4rxSCBz5VR7i6WiZAn+UPsBPyHfV78QGQcibD2OBJ+zY7PaZyUb+fK8/GwP
0z17Yrx41zPr2CZ+rupHjMaQ7Ey8FYnJfINWniyePrrJv0kfH1KSYc6O38nHm8ELzIEjWALrUlbG
K/fiyiOAu2fTV/Q7ZztPA0P8+1zjLG0vvxspReiC0X+oxFlKwhJiNSyVe4qVyMh2y5A+RQUbQfZj
hPLk2OV7QwdeRLkWPlb0eZ60igGVPsmF4Cp6JpRlebNFJHxVBZiePxYHAqFvOx5E1qYNqI59mSF+
dHm2vBvozQCJy02UKfi73TVbWJZcA+72PZ3qPc32h9t/+C/Zz/1Fba1f9xphrUXLhSL+zjIbIaK6
301LfrBujPy4IrP1NyNTiXDH7XqXejQ4YlYpfuZ5Bx/XnDYs7OO2otpgkNqazbYi0XNuOZY7c1Q8
FnSr9Hbsrr09m1rZ4QuqS6PA7FXCs/VsBXwacUObTewZMngv8VHTjAJ5tS3IrfRDTRze63A4k87o
qCb7zM3/oYqJzL85Zck6DPG+hY9WwUJcr5CbtsmDKDIfRIJJp6Mp/D4HCnpfLoo7A8+nk/DfyCMK
gTeDbMoi8BX93P8y8RWiGglb3OCDeFRdvgs/4QhcjvxMWnCh6MUqYobsvmS+h0wMCAfehyqgmqbw
8LtEknMNpS0e3s1HY9X78U+QlfwH/hSnSdXarrkOkwoD2a//LmlOTyHFnG5kpjB8WApcp4aUi3iR
Hr2lqiVuxo4Jqktwl4+W7dHT8vXLtD89vlWOph/QQyLgKgxYfjYOWkJTk+WjnxPLAk12Ycn51Z5a
9xMfDo2P0qOKgIfUGhIdghG4aMPF3Rw51c1SqeotNWad+Y4cQ3epRNESRRBbnr34f/Cc4iQqoWXg
ycUBT8r0N9CgnWZTv2jLfLK7LBI+OheFobstaqZPlIxGPecDJjd3qYuwPk9ksLXHFUxA6FuTKo3l
RrPiSWyBSA5gTh1JzPMrmuovTwDQGgl89AuJZnejN+9x2wqRypTvxJWd688DeKg2Nfgymt4um/eU
LBnD1swgLPEn8AStV4kEuXkcy87o/NFkOLzG5gqdATT+8gb8njdd9QAPUzFWFPVdkN/21Ge6nQh8
G+HeBzPzU7X+G7/d2nX9rpfzSCoYwzM/2SqxKA6RAGMxsFWy/DAzP90sgoTcYBwvtQ9CREdcwrz0
1ZgyoHehRGQteOYV1aUP8ACVgR/6PzF8GdD0Tug+DrXA72h8ZIwuJecIBPG1WQB23tnU/Ky//QUb
WJbO1QnCLyZxNC2all9MD7Ew4KBoZoEgdkiDQrgSoeoOimI1cpvSpLoay5V0Wpe/WG2Qe+WhnDlQ
J83LPInEudo54aAkQcVjYS4psHp6Ei+p23/Q5ed1VEdttRLlLAGQ2mwPu9V5KGFmA+x8xpcUmhH5
IWXwNM8IL2CaVdU7HtOWORhPxIT+DA08M+/Mtp0Wq3/qdrG+SF1dMagjzqW/m8QIEOftXTmXugGV
qtZACvljols/VQEl6T9/D+2DQkAbNBEb7ip+WFm7ON023f1DzLmtWLwqOn8+SdBFyVYV1sQBBJS6
5a+kx+ds9+sgSyv348ItKZzUIqMj3zqu896hmCl2Lh1szNtVEfCJc+tA6TaqVGMxXD5TwuJX+cT4
fVOzsBV5LQZ9wYNUy+bb66n/JQJhp2qXexVghh5EsIskaMquWEkoEtHxXZ3ruam7mt6hjSJNI+LJ
eCTAhHWwx8QaXDDwGgcBW7uUPdUIxla13arWwwTfYrilt06YyytHjmtcQwIlkhqngQVpX9aV9tNO
cEk6hxaxRn51fwTweBGba79//6lvKPwfYVNXi8jlL012Z1H5V/yQ6+XAR4W3B+oSKrqAbf471S/i
4VVq12sKh/7tmRliFR1v0BpecYWzhAqRNbNrOYHXLaWK/DPOU7ScOLZhZCFDDC316LyhG2aOHWTD
B/NoocVrFz2JzXkTDWssOJoympHVq29hLshsS66fCIsvhXbEJSmyjw7UqoxIL2YXgSoS0kqubhv3
TzT9gQf+BKBVsud6iKlhwUnd5B8HTJf4nfst7wbwM4iGCcj5Vc6aDSDVQcE+Z2FdyO5MFuQlTGu3
2AciDxSad0D+dHU62fb6EDskXrtZXPKoEjBeTuQpmvq6wUdyiW29eu5sWW0VrbRDxF1W0Kz4jsaS
7wi7kIWq0WIZ6B4CJ/DmOJcK+rEy8nWYllot0FHHVOwAl2KJedMS2leeyjjJQKTrF+Ea8daXfyBq
llu1NckIi69GbvleNkxUzhbvl5ayj2d31CJrVyO4H/8nDD2akuOAwUo+CMCIeHaljmOj19t63Dxe
Rp2wIFkr9zywrpexquYT8y6tmZeQc8ZO2ypbfO3LijYuvKMSm8ATNitF28bqbXKwq3PGo4Yyu2kG
5CVYbNo25nt19GWuOE/ZeRlmElg4zLy6NJlJO+Wg9J9D/tsW9+c5b25ySSYJKr7Nej2hrpd2BvFi
ImJH85VTtX7RCvTuavETpf6TMMYdxuDHix1wcD/bBPaWVQioWgx/Sc7Y8lx7VHSQEG3FB3HwYBUU
+c0o0+Z4ki9iyRb4hJP1SFc7BDZmw5jxcZMqqR0DbdzN2myuAZHMaITGQyKtQ6AzB+n6uudR/Ez3
exyrA23cJSEppn5qbiWN1htgV0x/kkT07JWRGpVjbMibjs14TophqLF81gkEdnHGXfwZSwuSgTl2
M0iS8JBglpDcULV/ubrhgpx5z/fSlapgIT43tRYY+BTwTD4iOWRiBkq3GQ9rPmbi2AVRHcRStUoh
ExR3sPhMPu7OZm2IbXydQyqzGx3CTF8Too4tqxRQ0ZKnwo2O/mkkdG1noEuOJ2VRq8wqm0GkzfCF
UTewsJwW2j0Ja6bZ87RU/4+CrAGFDj0CUzQu0njUYmE0n7Br89U/HLI8QuIeumvdcfzNmrv0mcVN
/nYtDvN18Q7KnEExymTRuO0hhtCjhljxg9T+QVsQ5ybgzddBbMpIF2y/ipK3sFA6qguUZAvqsh6I
/taVVUpD5laMjhXpMMcM6S7y94Asq4Abi7cVZFc13rKycr/KS7w6edcVI35cTozZiervYF1aS28x
WsAv1PxNtsf5xen9lWRt+5JT5+uSCsBA2CpmuYJ+U4Y9rDRuPi/ip/qlmOrfD+Sd/NX6vqPeJDGI
NhQPGPfZYDqc7vzBGsdqLa5n45PWdM8Nns54A4wFGU2alhgINYODWYdUxHbf1192Q42O33D5f5L6
ZJBUJIIq1WP3r0Kyoxoa1gMIBHeHzRGoJmxpKAHViPfddX8n5OXlAA/hW4D/EdJoQTEYbcwHJsnN
GFkMc/0DvCWRj7aWrjG83sSgaLUrq9pIgWpq4mqWjbaesRNjeB25hUCrN7gyEETgq2DoSS359Euw
X2trQklEx4b0P817NuXkh5CIYjsa4D8MlkYHPRQdSjKCn4p/4eRymPSwexO9gA9rYWiT8xd5O9dQ
E1DD/drqQUQD3egoDtugVaL98ytP6cLylWvnMVUHjv+wtcjbJYYRErcod4UHuWnQ1m+Z8XUxVPU2
mgChVkIOVXs7mwH7M39uwn9aK5YgFBleFMTHVUed3gsFsg9bQOqe+s0pJElMp+9Ppo9VGbFP8pDf
wWq2PUZ07s9YwvANxQQv38R2Af+/hX1Bj2NVWBolAyRW3Bv8jLTZq69/W4wShNg4x1YEqCi0F9zb
yt16ZNshki9xCmF+A5c2qJTYEWCgzvio/cTb7n6Mo21kOXxRZXrSwxHE/nvNDRhE4X53gtgvsO1M
P5r01PwRcuDAMsPSgjHrzujkSKKL3+3CZj7EtpQlavDsua6r5ZLv8drOzwrxaSYCbYa9my59SDmF
79MSSRUCKVQTqpRJC6qDN4gxUZqLoXVy/m0fkv2p0CdW4BEgEHmTnQYjNSO5GauNKP8NiukSZN2E
fGgmwJ/IUMqJPxi0YynbUjNEIfHpX3wOJA3vjnM43nv0qZzKHvbo6KRl8olbt+IDxLe/qVFHgRfP
/g9X/R5KAJ+A8mNeRWvSthymctTe53CnyU4rbtjjLVnIbL1DDLSezN8cgMjmoj4BKGKOTRidLdPU
s13KbYt2ARWEG/35bEHaAoOtrw0AwGlMVwrRMN5AK0hd7YWOZk0PI4eO2Wzx2M4xes37Nf8Yx5wn
csU0BozD+e2F5spXWmxJ3xn+cw3m5/1sn/QRCg+ENLIHTHe2OQ1b8wgMPzGPZpLVg46BHtl+4z7e
yTZLZklI2PtcFpTMhL+99zatD8pTuIt87fUPjWIeo7h1uI7aMXRnm79TAWsHGqVKQlwf2DciN4/E
OFPCKW5BGTZhi8c1WbdmsYrgDbjksReLCFIMVzHB+Z5h8wXaw9KbWcgM+Gx8ZRgG4dPSwUgrMqut
lI52l1QiZ3mTOKJC9BwSEEGz1EmXC0UzVur8fT3AcvxCG3fVKKqQ5wg3SuXjNu7YkJvMvD7/ZT+5
q/5S37oowFTieHrlfmqUSsGZ/x1CAziOuIIH0NIVbUrVkg3cM/cl2W+Tuk61KTHFJ+FwHAcwzild
lpd2gOq0Ufz8AW4cJGIvPVMvu2YvLQO7wnM3lzCj9tKvIiW5e4ehiUDnoFgGZEEF+iNpBRhQEwtg
kCoMHZIlynTZM06VE4ravdKZGnvV+5E2PJMsCmZ/UTX8bkML0mjWzLFk60+j2ruzJvXqizF+PEwD
1YWUj+Gmcni7cQ26EDsocV5ZtRJvX3md86PekAD5c8fjlus5DG/U27h7oknNXXWlZG0jKoRW2OVo
ZupPVke8xPAn4mYZwMjUqOor29EKZeKz8rLJhV3GOiZp0NrGRsfWGZEIJrza5i5gVYqyUEEva5c8
6vbBOMWvhx9ytRpbU4QmgzXMToaZ4vUjhW51ytOHIXnlc1L0TxKOxLVABTkVBGQ4z5tieXdSXvmB
aD0kMr7bp0s1X3CZN0ZoaZnFyRIONEAyPqHHwl4jkEP+2sp7PlLCvqBCChzZIfB89ICBkpvupeFG
J6fkmwnHLGwI5uqwgToOT6P7mJSg8jj4+fAjMpjOVMhzD9olpBl8BEfAyHxhB+xpOHAFSnwZ2P+F
Qzz91spJt3S81vD1bWZ3AhTsmTdIWmzHYgsI6QzhAgQTh3cDYEXBrh36gu19zf1EWiCAAk0pKJDU
dMZpevakayOjRXVsYup1+4D5tZEOppYriE9JIdvjWFvHIqDBPn3EA1LmW37FeND0G41pAqmLjy5k
vgSkNFcG3v2Bo5ei1N0/4Q7OIULrxoQ2mgn8sS3DpENH3Ldk3VGthfZf11K+HW86D8uwLTnp+0XS
T6ap4MyBlqR13c64aLzaOG4u+qKN9RjOZgeGBXgvRz8kMR3XIiGbT3i+Gd5HYmxQ2rysgOqmctAR
VhspGANCsAhH54pxwRaLlEnKEltblHAIiSJshkekioDnS++2pPdLZ+yoJJm35YR1zRFwLD8o/Bmr
WGLdc4K9aoZeL+CSlbOWMDBpm/NGXcl7Q9cE2aCSVP4eyLKH9bjS/2xoKYJXIrlERDmEBSgfJn6e
hVDYy16OGwDdkmEeZcV4q2zKhhFvOzmT1NY2ogQd2Q4uD0Unr950Psteoulz3tKK/d62B3PGnlAH
CpscqctIz0eoWy7L++wtXOZp4x/6vZJmSKaMo90g5ZDEAjBwsIFiY5i4KHTMxzS6kEXxerEW0Y6H
InDLQnMYFOIJCElolHYPWdFvHBPhM6zE1qC8jK6KBW61PJXU5dJB6epZbxc9q2RmwUx6MTzgBF7F
X2KNfMoYecz310kkX9H+Z87oprsgePX0ZlCY7IwMFTS7TxGaI80IC9prZ5zQVIROxoCGz6tM6ypQ
ifMD58SYeZLaA5bJEoj29Q4OuovIhZ2iR2zBfSj6kaae+YFl1AToEuFToqCvg2KNrrBZKFZZvucU
UZDml7fKtq74xn1GwjNRBkF7x2+1qTI/RRZJ3OvtRu0S02WLTaaJwVfV+3FQsSTuCi9cELiyHvAu
8KLjMhe3Jiy9DrxFp/NNNS0LyhpBLCqYu10LUn03dPJZAYa8RSAQTljR41EvUYGe8e3LGA6toFX+
AKW/193TdJlVgfyVQVbYVgvZB5CDfos+vmDwj4ZjV/XWb3KXWLn5b0HxogEwgpumyWxhBJaH735w
EtXGorKES6+nMFN5FCSM7LlrnZzaJQT9Ny3SgcM9Wkyhxsp3BPi+yhe6sarWwqbvKKk+R///YNb0
S3sBVLVF1OZ1ohWRFpKoNhlLGDVuFbOaK1OI6vBgwLXh9zLAtmVrh68+JQg0uMKoZznxeTGSlAHI
DmH9EqRfdqQSg4vt8QwoYowf5hKtcrfVk/9BWweDsxGDACoPDDGU4NQuTnWMrjjxnWn1Pie/lpCM
hLN6Gz7jsYl1NJBCEj1yCr+SMEClo+By8+HU4i+vaE3Sm6FPKWii1es4hQwLLne+AICsRHvROicd
lhpngiMfiBWPAzFUISd3+SLyWoOnE8Y2nr2tMruWKHXWhYXr6AQ4EMpMMUs5HdaTb6HYQpRCV3bo
9QGjL0TeFIFcl/a4DuR91E9aNI34oZGEhyC8rS4s9iuzvESAYsaTQjCKZnVvN3fTOtkgD1L1Omzi
4/BlnTNHmUl/6ctdn9STM+TBIokRs3M202HzbcVOkAV7hCpdmZ6CWfIeDy8QEh9mgYKlTVnLiSGV
QSjK9OCDF1UpohMoJ7Ks9vH1sSLz1UyeFNKBTL38H38tOQgcDWuykxn/taiYOYmrH0xj/N7uLyws
4NLhIH2lRN9w7SApI9rwKqfReqoX8w/U8YkR1hZXldAX4dFdaFJUc3xsCpwXuYLIPLdPf6mQ4/Fi
48juwXfIK8DXrR+9tbjR2QQNpI4n2WLVJLmURvTHh2+BMIHVX3OoE0cey7oyBQ4sNxw0XIZ/76BI
ndpB5qylOgAkp1m65kWW9J6/v/c27orDujMGkyg0y3k3FxnZ8HQQJQj/lmbH1WkLjWBo3vtCPfzd
uTupgU4J30KI/wAM0zGNWDGDswgDE9WwaAWmuLOlcjBcM0bgy2hoah4MaNLKgX9Y2+3PkuO/aHrL
PIm89POKVtMoR60HXVrV5smnI7K/dysIxdGRaarJrc9OCRoKII/Dni51F6RBfchV6L5wDBpeQS7w
iKgu/rd9KidomS6+7vQDXHLrwGbiyZ56kjk0i4U0FQSRd+0twuucsWpTQN8EF8qWlOUhfzZmKyFb
yzkGTheN23/HKoUmeY/JS5YHnhX+6CZWwv8inTkAj+Ina6pDqckMYvpJvE5MSPFzfvXx1PDMdK3h
NWPvxKBx2gIew8NzT4TqWNSO5pkgJK/F6PAVzJ44vdU9qDdBUHryGPduIry1uFKG2wqvWXH6B5tT
6A82BM3WdH+xdSaJTDiHHmM2R8B73K/qhWgCcAmERCOtEPt+hPdLX+EfsjHhdox9h4jH18c7pkO/
jGDUo1wHNTJ4ToK+3IjbokUr2A4UkYIqoLPcsj364TVRBL46Kww0K9n0lqW/YTHsuKc82yHQGOzu
XghGHw4S/V7Ph6+qWBvSIbpc2OK2WTHcSNf8f4OCnAcei29mr6f/0zoYywV2CigJrkl+OrNWCnz2
zT0G4xNyqydPGu4maTB74HMFWJTg3B2wL6mwrag5a7YB+MsrbOz+7SF3087hiieDEl7nYaIJ8vF5
BO3qEjbTVfhGLdwaYWBdhv2v6fJCsADLuPQ1Kx+Z6Y3waPrT5sYdq6zDdDdhZFlKpLlymdPxFl9g
oOCRkavVeI3DhfePP+rqt97DKos2XSkuFIz4nxmHFGLv0mHI7eTN8+LZsAeVa7eTjhYqL5EXlZmF
VxkFpyZqEV4FOPMEA49B47LDnOPfNGwR7dyuYpevFARz3qwcy51dUUixjIjdpXBmE6jAW/EQC8XB
SPRYYIKQL7YC5LD4amTfArfKbRM9YNDC54Qm6jfes4EyyM8a88TmsT4xA/pxwp4QZYJpe2maIglL
HqSB4GfvU0NG+gxHQyJcBM/0rSHX/Btjz1dhZaRurZABemEJV+xALnv8YB4tuJddDGZeMJtbUT7m
IEbn8W8G5g7JnrC3BZiow0ACcTp+N15FetpvhCFz6L2fiFrtTcirTdzmXlNLkw55G0BqLKrxNj83
YviA2hzKpdkE4tFtaf6HxRRNKUtW5QfdZM3lykmx5YIPWw8rcLQH54cE9O730I6Lj16AUmump2YL
ISnIaxi6OSU7qWOAOEWjR+aBvxbBMfWS20AaCdWlKURhGeIaAt+JaV1p1fKYfRe7pSorK9SLzEq/
uxnGSDIJyJCs3Zn/Z5+4Y0EQIJv+QPsUSr53SZNXCKqH78+MHwOAGLgni3R0cZImc/t+y2rGex+w
6OKDM9qXYXgGDI7KrFY0UFA/eSTlzmPALfDDqYNxbSYdmCHRZx+pprXZ5uE7qX5re+pEF8lDOBnM
P2WGlJWCu0Dh/dguy/1dpHZ+tD4Gg0EDpe+QPM9Q+NFOERUuT4x6BFibgvOK6nMt6HVoHDVMV2wv
ZAXHrzuXBNNK8U/JMRqfZDHNTL405r7e0BHJ1fA+eD0rtzi+8CvYJ05pk3s4k6bxhv31/9qq44Qd
bDuQc6iGSWphK6NMTScuz+Dfcr0CW9B62ZcMgMvb6yiTYiDCV37VhHGLYDDnPrKOKjRX5vJkn6Kt
DSSh4MZPP1TyT7FhHWMwk9BcecZrx5aLmPYqQ7wcsVj5fRghNUY5m/QwD/MoFBWL+57WOuQBmy4s
RVdqeGHc2FTIWH7yzIMvqEEfTMAme2Ju32EyfRb1vx2hZ2sx+Sbccv552wtcmb8aFBArcGTWyd9c
Qc7w7SQHU94XHgVBqUhMTdwvLdVU1BY+DtK0ts+D+pSRu9GzF4YQeMDbX5SvptQlILWSJZkNdzBM
eh+5kM165HV/wE/rCIJ6B+p1k5TNS2iumb6HpKrQ4QGDwQ6qJVIH4XQPehQNKSwwINEnMsSg853w
k2TFvw8Pw8x5RAsLUVgi0EWQR8OimCsn3cyFMo71KYL893umXkuInK5vRV5ayT090AF8jpM8UlIp
GGAP4eV4TuaI4ybEVcKJFTE4etDntWzsUAOPOUzuBG7x5KWud3LPsleiuqcMviSMWfLvZngKg2cs
WmbSEU8Vnwp7mpw7L2cKcZkrx60U6J3XzdNucs0dUTo/bu5FHGu4kkK9yCbGlqLvSb6G/s5X/j+s
qXe6fMa3LX3WPzxsIaji6jJlRLXOqtSlyRypcjNZumulvyYQsiJCyfkF1gJtx332Xo61szUzflNL
Hj6wRSQbEONU0fdtRrwL+HQ48aah43Xihat3TiZ+G2yhyyPCs6dopTtsybA4x6A87yzb4pY1aHHq
189tuVBv3IfnvUPjElQwFBHmmRZe1P1NsG3dZUxgviUUsiWEK9ayK7dMPPVw28gAmLl7bOcEZIvy
NNtSOrK6z4V7wNoEFla5FvJWdVmwD0qrS/+NcKA06BOUJBE/CMsUAeynaUv79dZxIV3i9hD4uUZR
5KIa0aUAAQA8xPaavZ7N7tNv1HmpssuC8c8oeKYaokdahP7IyQPxENSrLq8+d1KeKsNRMdS10b6O
9QVp0/HJonGhgWr3QS1dTBVtIlOR5QB03ZIFecbm0M5Ce/YLZE7NqSczVbTZHekmLy+02vkKCGpW
CYNxhVHj/eEF4ZgY2ZpbTqpgi5HjOo7kBpOdQEJNZBLQYZgVZKgTdmB6YR1ZYVXyD0N3tQPcJX0Y
fPI9tG/3lsUTwFjsD6nCET8nkuNhgYj1ZR4/rQ3adn/CZG1FR2dmdSwrAkVc+pzTDDIGKRVRYRH3
vhfSx4UZWCSrIJr6a29J9vxyCrlTnpM1QNs85XgrserAq0TSqDp1x2jDCrns9h5+3HeOBk6a94Hm
JXioaFwwtwZq6IQePwwcMKZbD3oZVo4pdZ90q6+alRIISKZtaUGA+6Y0YflfAypOt7NXwTYK25ZA
8rigaB8MhbcPoXDzHrDsCfFJfQ/sPp7mmzZvUAwi9/D4rllRu62w5+29a9tL9Tqqi65yHBoW4RLW
zlc8xvZNc92EmhTYpI0YeFdW0AJ0mahzz8rhnb31pPJS6ffvOn4ypWJhJKxjIwTWmd/mqHM0pc9+
KscjYmPc244n5iUElOE2Osgzb1AGGPQEgiIiERd99Kwg/wUGllLqr3WmHl18CUcr/vKsaDUuwGxF
7X6kkvF3ZnEJY66xxJAPGQUJ//eTHRClY5X96eJfkIlY0Z9D583Q13Z/ndM2WNUtgg1qwxZ94sYt
N5z/tJL0Ef9PyyACZbGzYNQksu3MMILX2XGH4OTBZ1E5rwC8DwC345sDWGHxaNVxnJJhLrS16OUz
0ZcRxJUKEUg4P+VTmU9UT1A+mMbcR2NgLO0S0EcBtr3OtwvtOs9NbjECXFUsvSJIeWJ3jL6LYZDR
/koqV/Y0V9DD5AKo+xsGS7iHxBlbQhzA/d+CR3c2UDmYIqnN+z8uEovlrjFUGGtODIj+KqDwn4oF
/ku0ElWhJm8r39USXtu7XJKet2n+fek36HTk0ohDpPOAKmvuHTvYVxeFet85kEN0ecRm7ZJtd8NC
8dep0WPCQrEj7A18BEyMhN+nQvmtJYTh+SDzKugri5c2PSvLK1IT1RFDA6N6+qXUjrgAACdJOc9r
d56QQimn4nOVcVEB1B7rq3CgzAfSkt/iXmOYPDmhO9Cxs5Vy2gm8pz74apZ6INRU09PQpsoq4RoH
MpQ6LHdSTdwSsDp3L2KsCBRhv+3lqY3rT3iMsbi1md83oZ0yYOFSzOmj3rQdzXJ8mZbs2csxGVwE
iCerg8FkNWtN04ewR/V5N9qQmdR453SZNq4pOIfJTgvIG0WjjGFSG48yuqhcyp/tCHLXULTKKoK1
z0itnE0ffDaUWekjXuVZBMNF+1PcyeBbV1cbv8z+BKbyXDZAcIK2bQyHG7xV6eASDLzXFEkgbOv+
gwJ4rp4eMZ0n4eOd7+mJwxX/OP914A5afAB5rG9pg7grcDKpc7FMTcvarWF5DiqBPTgzKP7ZrZGQ
guaQFQqwLSfgeeUEkCUQcODGSDavjN4C7jJCwK3VQgQO6MrbTg9870DOo6iReV0ijnumHvBbkmY0
VJZlTUSX6Xdkqtugnher3LKS4xUcsQdD0ZhgeqB0vb3KgNdxhiv5IabptjvXN1fqZxkrbzzvhW5f
rsPQwyAn2pAhsPX6+q/91ffSP4N0/ODt2gIvlG6PV9NCd3APw1QRY3Q4EBos+6S9ZcFyLN2p11nR
2FP+yR1kHOpsLlwLSiWLQDPEsb21fA0gjBCAne4uNC7ytAf2qg9I3ckeUV9BLOshjfQClfFWIE89
DLP4lt09SfXczqDOVHJ0WGGlH7DNj22Bi+Qe2TW61G6GRpMEeRxEXAeTctyT2UUQjMIPXSZO6AFl
NMYbzMTEDPMba1X+5VBVUFet+taIdEb3+BIj7I84fvjCJiYKnB4Ia3AFzSvp3ahGkF5bh/D2BeKA
jXazfPUY+Ne6kBXTtLTeYmtPpHbzmCkULQX1LSWGJTWviXFZM1+4eQyK7GMW68L2/TyaNojw1tmI
C4tCbzCV+Rc02kJSWaxntPH8FLFVCytkfDSJUBfCVLxNF3glwU4UniENIXI1lsWN2rldqrKjAPUc
Ok9IPsi8UvT6iwtKruJ1Aod/Pp/AfJV+HaaTd1kv1ZsjtK6FhoO4PSCks1Vi1fvpup+4gfW6vMpG
l3qimZTJPf9A/wqXMszqQFXYnBkDS9TM8elKytI2ehs5IGQOfGvsVPOnhUDKbf5nlxnfOh38LOla
tLkKnp5lzTp9yoaPvt1xcMnc0yLhz9BKjyGCHxw3g8kBDb4n3srhyVopsiL5SRxCdlA5LPLh5x1u
p4Iv7lGJaq/PBJkNQw7o7ZOFAR3UantvN/afpD0wk5S770wxCQtCE5HUC5uIRnirGRs5PSNCJu2d
fKvWdDMymtAG7XfiNYckMvG3iCbSkilO0kyt1DsAesVbh5QWgE2yjzK671AeVbnoWq6a5Y2cE8cU
3No+8Wmaatmea2w4zf6iV2qUxkl3eq3HG39hTYWkC48ze/0aJ43ufGtr9RYfVpNEbz0OB5rhJSEY
HFy7BIZPOwz5TAZNRsf+7WKQIb3k9+7JsRXusU+cuL0Uaz4pJCZVOwKawIzX+0S6JugYde/hcQpC
KxEcyVq4/vucOdEWQSM8hWEeJ2Yr8lnCGjXYoOxIlgth6etmdABLX0UmMNbXG8RdurS0wnNRes6C
zlq1G8GLeMwzaez0yAYd2wuKiN4JLSrOp5OFjloFz92XaxLwecRHRaf/6I2+wAToK0Ww7/lw/tKt
FhbBzG9p0hOSgEOAwvkfgsWPuRRK4bn79Yg61AdDjeW1vOLoCqLLfcVIfveIb3szN83jeuYT6rzC
oyvBbpYAxbJ84VnjwFek3W1L8L3LCLEN9CeHps0Ia080C9YmRLarz7FyBM8L4VbRNKRfCpzc79q0
A3UnViQvQ47+bU+yF1RwhiDsdU+joGwRbK45CCHQOvum63IkQLFUPhJ9V3SSxIqlmn3xEwufGZ0I
ARTqTcPRg9snA2+L3+Fr0nATdCr36Iv+ETJ+n46KygIuZmdhOlNGpqYK0T25yzl4dhCVEPuUl8SY
fmPbb6mFtZH36Pg9+rk9FSVHMTSqAGYYPZ46VjC/LgrIidgfC48rLwk5JymoK2X4RTbNTgTGHamh
PSFl928a9FdaXr/VIKH8pHBMW76xJQ8Hr1RHHMmmu/XlL+ovCYWindfu9SDh64QmkjhPYWeQg9Wo
yEzAbop1acis/OWeSbaZ4ED9jV2dwlclns+Ef6Tqu3Xo89XXqeNuJXLISjZdThBWkwITUhViqSqJ
58Doqv5hOgvNMjj2MeesznDG9IjaH2assYfdxYq2V5UbuVpn1YUlSZaUMxuvYmlK9faEN60LuW27
K42JLYQIcmOlPPPz5pWMMJ0DInVr+pd0D+qVD3jQrzYznf1vKri/jLUMRCAPjLuzdYvEKIyusX8P
yL3kLqZAVV2ifyYOz0viUUsJEDtNGfKjUZOJN8VWdSeohTPOV5qBVSJemMqp8fkC3Keu4THzI0yT
1yR+GsqyjLG4pTFSc2anOpuKFHV93hTyNzPIIH7qWZoW7mbB4SddzY4DwNt4eVa6mx/jnl6kJCcb
WhgmVAiSkyLV9xMxOOnWT4AAD9dSzX5Sa8qZwHCBkda33JcODBuf8cHqhOgzV92dE7VVs8JiXQlQ
1hfvNTHRrtHgtgo7mlt5WXffhzyD0CLa0YmIq5xOCPlNt5DZUTZMQPmm9IuFb40yKVV6irkvAIe9
ftiLu3/H1+70n+Jln4799iwX1sGZ3YOPhjNDY0R+mq6RFZKAK3UByPiTzcDWe6SfFt7Z3nuzHIjY
2cVEAlNkbirg8xbhXlPX1L7Ux+LPWyaC2ryE1a8ALI/SJuo5yhItbySqyRl7TebOd5jTKQsjFqJB
Hihy2w+eiAwexP/RKSVKM+UkCEpKosKgwzx3U5mecr4rTPyO+xIl7YuQwErKQVNNTegBkG03zgA7
d+9Nfxtw1rhmF8ShriUqf47kWTl+7hM8XMzFAG1p8fzbfNoukXkCZSurY/VvV+oHqt0JREigrR8A
i2duetlkxAoCcRtoKhW4x5mKDwQ8q/1Jp+EpEJzb7i8rDgQUqgBdrp77YqtNFwLfwjhRZHB0tQNg
TnoGCw1y1WJnwmMoaUHwxP09UJD+r/MEQpqvroWOWtbQZsD+Y5O4xwm6b1K+aWVNnekCR6LF2iRe
4P6Qcru5cDz6UN14hZL7SWr3U42ChASN0zKQXsONXr47w0gsHUM1h/T5F5vmzVP3TuUcqeCkEz76
LdxFIL+Y41bWEQvkjNDz5wDa+GmdEv1vqcKbWJTf682pgsPmUj2q3V+Uk/h2uEAbPshxyjJZ3CFP
cTgavO5XSlVdrSJe8KfETkGcIEcXkBkqpsxwDpMBcCiGkwKZqlKl1Jz0+v3tRZLRFF88QA5R7wJH
R3lB1WbSa2Iz6DV5i/ikvMPjpLpfk+JVYUWAaQVFslbbJMpjkszmF1GfvSG4T1C2ekfGgtN49zbh
flOZ5wGxCoLhYDgzhJXG817njYohprQiPAyMRtmYrxr/5+SUxinY4FE9hW/OH48wrJf8uQ+aWXkV
yT2QqfjG/GV43EIf7zbvjx1Wy0OAAAGD+LmN9C66S+PdZ32ej3n91rQ2/OgA0WLaDAUVt6008XC7
yE7J36plJnKrMby5PB4JC2bEUXCdPEpXbfKSJBP+NHLlIKNckn5zZIwItX4JWEzXPKQ3uHIVs16r
InZfpAP//LYHGe9h0EIsROcKODy1Yuz4swbcrS9WHP3oP0XJjN93nuC2oIG9Or+SSk1nY0AdzSU3
Xgr3t25eYD97pH16KN5HHB+C82raXkWviRt951mo6nz0TbI22S32e4+LqUTSSBOw85f5Tl1s/UdY
puTKaUiUTqOUJ4XIYRumaymwtMENoVroCExs3iA7IJ2RNVB8OZ3a4rPjjEKxX9kLmn/cedzJxHuB
6Vz7f/qEN3cL8dCqDnWoUu5UcL0NvUTy9CLaSDl1YELhqlQilB4RJxU4s/+lxe1Heymg5mePXS3F
RrlNijwWLcv/zh7IKlerEL9c0Utf5XUZU1TAGXI9a8YdaUt22zPZv5KWvM5wcR46LU6l1OonWjPn
DZkLPyy34uV3BZqaYJTSV3mWZPVgLTz7yPHBd81yM0VsHEdYTY5dn3y6hlupCKoI2WeZyLVv1JWv
hTgJ3RCO3SHho6tqbY9idoLYtbB9USKITEpOsxhCh/8tCd4fxBv0cgvcCGE9Wt4Knqmk9yqYpd9n
MqqG2xzkq5aQ6FWIOEI0tKd5vbPufpmeQCSGtQ52lSRwuXgBI6s5ACKZ9j072WAvtqzWlJN2almd
f9ZgOlcYI4Ws5bkIWx5L9lC/wJAVGygjrPd8DG82nTa7GICZ3MkNk1M0eYJ5g5sND/OhjVRggWG+
FT7xjQgbiRIE+PkQIy0BzYMt+pLbG51E6Qqxzs14bUp0lEvTFhMV0eGp/DRx8+l0ZerG6RbKeCYs
n8DB2BurSYHi7DzpPpgIQ7mcLuoqeDfEp+gjUQxI1q/3DMACNX2pxRF7VzK9UskWmc1KUnz5YthW
EnZbomHTV/z2BEP+S5WS5JaZc/U0nDvW3xGv9nSqkBUzmWDgzJCIyXhD3dw8BpsMAx5pl4MgbfXV
wfsw19iJXDHWtyMu6RKdY7DpcKMJ0k/jouA4zHUE1ZAlAtgMcPd1q0f2+SAFMR9ITtPfNtOVJtxG
/wMKNicgwQr3xNg6/6fxuJcuECmzUm1rwUqcSw/Y8b3Cs9Uv09sYdK+8ZlLy2y88BQ+kJgInDAed
t8BP/aw2l6OKlvyqokvFJO8xiKIzGC3WksNVdXN0eHpX6UTIt2Xz7i/ubsR00qFHhTTo2dn0eW2k
xTgCTxmTx5ZKgcWUZQhCow6Tb3n+OhSHygKT4KOmQumYz8ncxm9p0gujJaXd6yf0RRezruOJM0j4
TcsDYepeYZGbnDPO8bwJinF3YcwTngDOVzs1XxXrHVz8tDNAmoKppl7gNTKaRjxoF0LM0vcoTZdf
lbDl0Z/to4wCqZYV07EifLdPdHfJaiCf0RNbTiJc+7+MpZ5J9hJ/o+haXWxy5EHY9pziwqyzOMUq
jCOtyexI/5Ty3y/7p8HgiZVi0kpikqhOaUC/lMqPaa7NejqBBf3mIR8GfjQSKPck8zYOicX4z3ql
8dEfGqDwuh72vyeMEVMPAF1BzG1Ub594ErRFx3byk5Tch3BzRqRNdZbvMb4aZyja6xDYhrldKT9f
y1rHwMkn9qrpgC7+qy5FCNUFxOjlVv7ygK1ckzo1i8ieK1qolQv4ejIBLsLn8LS2bHuRjH7G0HJ5
nWZM4l37lWvj56mtBQnqJLIJAbaLqq9n0jqkZjBy4zY1kKijWEvcJrLY8d82KnFeli7zhnKa6fXX
Jrb6ZaU2H4280Tt3R2Ga4dy+ck2PhkYzH8RUbc2VJYWPgbwpx2alT7SIMWV3BV+26Muxb8yl2/qW
PvbjUaVA2+VXxVmI/6EmiFqoqJ1h0TdVmY0spVuMi2i2HfU/cnweCQWX+jDpk+E9Y3pUD8kwXdEg
rt37xWjZeLNdlSR4jfS1vTvdFHJ+p+ZG13L4JvOzvLlX7+tvGCU2LTtyNzCoJDsNIm6mEKANOU6B
EMV4QSR+2/OYAFLcA/nYfqNL9TjnRokKa3eIrt7lIxXmPV2BhBn+Ut4flW3UwYIJd4F4iRXtCkq5
Y4L4vBfF0I/PIZ+XyjZtQsZgsXFX21VccwJ3KFJAJyN7XFvPorbq6CoObziAXyLv0brYS3m64f5R
AqYjN5M5XvAou3viY95mlpSVeAQkY7mrLjYSMTtfOL52D15shkAXU5qCZL+rvoeaIMyk0XkPFsQ8
uyM7daxuhaN4Im3wlcOR5GPwgLYhqIQ608PEOE7M7V8UC3x1gAa4a7MTol1Q2oRgO7D62Hy0GWVH
L8nkGR7+Xdy/7ADBIVxwXueUQErKOENceeymsN0YnbPrGgXFGIEei9vvTZWXQBCAwELW54lo3dDn
lSY6sPNmujSM7cbmDeTSivTfFiGFisrlidxGCDRSZGKX1Ozh0Rn9a5VRanNiQHm0hNxtlLNqrOQO
oL+lBBalu7OoDEpp6WLQAh8RbpoGuva2bij2yqnZIAUWWIfcIlsKDBD2UF70k5W4slIgZYWrehuV
bJanUR2YkUZVLk/GlktUq5J0bta5k7eqhp8usxftvcMMbxn0JtNeJKMVg7dPUBVtRax69ANHUz1c
MhpvJErBurEl5T+rmO/nptOgdSuEVcUG1CHjv7xUAS915JIO/LU8tEkQqpqpi52EIGj6OfrvUeEc
FFwWuUFSdX0VZNrHMjNzIVPDjBTW9uQ5Lft7Rmk3hbCCEC4AlWEc+3Cc0cLJiBZx7QwkOZ/7QrM/
z4ons1y8GrwhtgaQTYq3dlMnCPdVFc5nBGHrNOH46uLJzfSO0hvLdNUsndQHQaPWCAis5poxb+WM
MuHXg/zhbI6pYuxhcgSw9WZ4XCYtNBk/WteQt8ZVP+a9V9I8PcoKXHXD7XpqGiLQuobPfdUwyxea
D5gN/8uyC9gNXXn87tqPsi2cEKagajBxePyrg7TJTomNjSBELoX+an2zQq6rmb8N7VXfBc8CaeYV
qz+tTUaLNxqKtdIjQrOVFxRr0j+HwThS+5EmfWA2bdifQe6q/9KI5si464igdRnz2riU4a5ruPo0
EQrAaaKZ6rGtmimtFTCMWqzXPuSkbR0q/NWwrtJ3bKGKG4oLJCRt8A3gISmPfvi31APE/uEIjRiM
u50p0TZSRqlxGMkXnRMo9RJHK5CTLCJNqF3kq6lc21EN0Zonhe0X6J9dPDMsi+U0r89mtjSf0w3q
gFOE9RwCsZ4ZVYKyTi6DUo90njFAgV3mszWx0epym0gqfCaG4X6+y+vDRUgfa7atZBBaQ8LYaHys
tPAq4wAgi9QhVigvfwg31WBvZFLh3BIrruUG5cGlRj1oVkSo3tUo88PYbhEoAMUCuoNwIYNoVjmm
efxun3b2xAJj5zdkZWjX401TCodNPHKiiK3wq+qWXh8mEWzMIZ+94COQubDMU0LRZ6SYqIGsgad5
TEe0XYJxtEdUup90Vt/B92xTCf2mH6yi5RlYmjWaERZk0W+pSyTjtW3DLUHskINUW4hhusWF73tk
3EXU+4ofvVI+RVQx3qnDhV8YJkrPBPRxkb2ZPcPYVdVvsI77uKbHIKCgpdoZ5VFR25rmQgtmcfMl
9QFrx8LtKuCpKxEMGT78oE83p/RjpQayuCzI/yZbGrLjF5f9vico+Sm9YUXqgAfjcaUc3eVt0b4+
xm+OHsSibS4W3pfUgQsedStRG01jYgt19VRFs0GDiO2MjNmUkq+CwFUok42cfzyts9/BazRcBgcs
bXskV/ugu66L95RMkluyfFMvnmwYpSaS/9bE5G5JtwHL81yy5e5CvCfE2zIwSbZHmcQgEEIHgwjP
9+9Q+kQURCvC8hk+uMs4FAJp9kPKEdLktmx5hdPRcV1zY2vyoXjv+vNwv71UOL2Ts3dWloY7bRZo
2OuvQN/clP/xGT0tuMxqHyQziccYZfmsEx+Plw/39Eiquxo/zDddZgEfwLSLOl/LksY1JrjVJM8W
X3OBbmG5iExBpqpV8IEUWjQd/9qOUJ/Z74RVh0tkLFmOeLa/MPjrGZ6H/hABUnOd+PYK6zOUJAyz
/hGW8g5On8/nH2MCiuNkIsGgt3eAiLIUlQqHAVkXj3xocXd203z/JcuJHeR7iRNsqxMh7QjsMjHX
6gbdc5j6OSpOdyNTsTpvQR8Swwk7PTo8bi0rZbfZUszzWPT6Gm+wvjmf4E5SSfeil6VT7bau6Ss7
4IwlVxyMgk43s26G8ldhK5Tlhfk6QoCgyh3abdISkXiFYwNHcN1JWrhQ+zlg7WS8UpHK3Q07bMI9
8pIYh2T/cet7WqOelJ+yG1Ua73s1MdvT68yfhNlK/eMiNQyOHi+DnD/QEQXhNm9XROKPiznO57SJ
mR9jubFY04dl/5VM/7P91/b/0fwkS79UuCmV0fxAGgDvhMMa/mJdCVYx/6n7mjMlLmlXQLRhff6d
ZDPNPeFVeSkkntwXm7z08WcSkLvQt5Rys/IQV22S04cvdGBVOVpJ1zbUQOMWveVpsJQQyqr4FNRI
JPlcJ2yg2FobpN38Bnz/NjzXyg81nEqCg5orEBDQt/TtcVvRExozg/1BTpFhmxiZ6FuSZxF0+gjN
kSOpN5JUORSxDiU/dRt0FfvQ5dVggc8kiya8jFufri/HJKyjBJRAIT/Bs2gn5UYTE/RVd8acc80M
Fmjx3XokMI5yzijqwFw83BpKv9WBNTWoRov6ZGlycNnYai7ZHMh7BSEJ8V6rMmQBKEA4VOO83GPh
NKqvC8xZwsiev/p/ueoKWRQRHNbhH3o1yFgFZIWwj55u7iyFbeGbEmJwubvXt2t7x9L6g+E1L809
Ds3+1yeVu310gkc8I8fOaiv/rCtOn4YH5nGYsybUJzz1+HQdUwsViSxVafND9MjKSz5CUPk7ASyn
ebRc/CIoPHLl0AmQAsfE6zRqnHlnHNKBhY1dox4hVbdT/OMck12W5p6UHBOINwVJoeOAFticd3nr
T/9iU6ootLA0bZwYhvPQ6uD65HFq47lVfUwvAcs6aLx26/08dwGEUHxRmj2jae5hjKghpKrsnReB
7TqS6FDRBvFKYPjdFETumyS2BGq8dU4cmy4MLUTeA7xk0e1ev3VsSLV2z/bnfPxNejkwHjK4S5qZ
NW6XatNnOF1rs6qK2zmi7v+nZGHPxya/Z9JdGr2zFAPXsitCAbGeUzdDkXRbjpGgctxDkcfjoCOs
EzYgukZsTUuMlahY5IUnfitcJex8TzSj/Aaza3pYhh5vSc2rl5RHnKl1+wbCdVgRufhRcNB6v3yt
UaDLhU9G6suvhwOf/4TdZaryMvjtDZvz3+AYbmyKKCzIVQtOLtq84p0rivpzQBbVAdRjCzhqbgWX
y6k1O5alHZ2KRCA9g4UMb84TSJyIAqDYFBpx42zRZm6DyLOrSKfYikAZK4GvzXSv3bunsOnAGblW
GSiu6529zpMmJ6NoJ8WUkkMvljt6dN2WR9+d3izCCqB+sCwIxP0AhPmnwEK+9397UlTn8KXkkLTd
gpY4dZlb48ecO1ltvYhSGYMkBXVH2sG15JuR8+dRaZ/ULFXnZX3Wt8E53BbjTzJN87LhHmQYiPKX
9dUhUE1Zi9Z9obxGsn+zTx7vvhnvXKILvDqe7l4XLIWACcrI4jd6A9o1ADS8lX+R2KkVzEsF5EEm
Kgqi5xowgBrQ/ym/NJcPZzPQEOrsTY/HSfIDGWFEOM4dVO/Yz0PVA9dvHsEqgMg25KudvOV7h/Vl
w/Lj6RE0ti1QBNGW9atE4rEBj1dGdWMsAe+auggU6Yno89rvS/LgmH0uB6tQTu01Vt7aTKNO9j6a
mm0ukA5Jwqil8PO6ZebpgobzAq8Wb8v/Fb8EOZQ8zwpet5VZm9sABGuu8bxfvf4REvAsegxpyZuF
vK56dIkCCvk4DVZhKo5yvyvT8T67Cd+BgRCszjtBrbdh4+LphYYuTFip8MT0xzbuKAMZYU4vNBMG
fd6PB+CMEAv7zvHr/euxyYCPlSLYMMjlnMlf5SWB/OLgHMY/6QvySCVZgqS5hpYDHn6TiQbJLXAc
4cBESlE7b25zvNwSaNp0OFQObwXGu96zu0n328aeX123JHf413NJWOrQ0tVFFsOe+74xAistgc/K
NEPfdYqJbswyymx6YJFZrgTE3NjIdW8TbT8UGLyoMJxfYMrlDEMLg4w0NwBJgbfjBd7CuW97pi5A
DpaIpakn22LVEtvzFzTsKEeoXu21tLVvFMSFaQheamzLBuxQBx8Zzsg+GPyWYzxSP5YAtAxCmKzn
uJplfnfXdc6H37jwWRMgZOS6k9L2hCyPoHRvTRR1J1e1blO/DkDGyOwCvBlhrokDT9nWJANfzVPm
sNh3w9uSTgEtFHlOGKCeTdsobqidqBan8QxmSxpkVoItHO31gW3geJbMbuFLQ2YfQo5L4gcEDjCU
Ut/Y9JtqYzA7LkjXjNgtzct1xUvA5NQgTxooWwsz9msV8ZEwni7M+/BzmLf680cibUs9Kt4Nq02f
lhhD5fx5rnP9+fo1S50XLZCQjB3diM4MbKso7NVQw37qTxSiMWxIY8NItNbk7R4oNidm0YbXl87n
6GkV0ark6cGn74QpotaJ5dMkLfjG6p8XkUUtu4Fbq1hlg2klGc7wAP8UpaHlj/w8HlNQZmaJj5W4
uAEys/zG+PJZkkVC+FlJK2WoAD7+9+rmH6HnqU5AKTIeBu8a9mXtBttZdpEBCg9cwqMPNuoGkKnT
VU/nM1w9afE7x6V1HTR+v680culDzv67DCgfwMY8TwUocCjZy6noWfmW6BPBT4Hy5S9gq4OsbymR
ymhSAMhb5z+AXkgn+oWHmisw4itYvjedLJGbyhaeaeY/boNONdk7zYP2XOFUCW1Fzw7IPERFcP91
phS3YXv4/mw0676SnYR+jP5f+ziH1+i7fA/Uavfwtk7YOgxtI/UlmjfHHlvD68kcqYFliK6NYaA1
mp0Ghg089yJll8Ab63vsa4XcSMnBs5qLZHiXDuCeONLNqCKkYpnvYZFGlCqaPNrJP1yHzDJKl1EY
YJy3JOEqTitezm4psMQ/lcB7cGLTZ53X5BCSbcMsf+DY5D147CIbXpe1niZIe5mhC/nDrlBi41Tx
sKZ/EN4kdU42buhDko0sW9rPOKf+vKu4jC8LPLd4nK3sO+bWOGJAZG0qvquaT6YW5UWrorCcl/hV
JYxcdbZixTDml+BaR63sRODJwMWuONjIouM4yVZ2TSXpwpGCW3y0c2BrMem/WKPQRdVSaG2bSl1V
+aXu7SEf94midJGO/HcOYYX/4ON89NzhWELKEZF2dBZ61pS/m28Ab0Yh9ogmcVgYBBgcoYBQA5Nq
Uj4xonRkLcGGCkT2WckU7SOGOyO0Bz1is/zd4GrTR+lXGmu0bgBoZ48WgoZHpRmLsys6JaE3K+CJ
OkusskNGHmEPBvemxhzrcD+xeIWG/aMOyUD9x4+xEFYvboNWqCo5Ib1t3barwNNLUNLynjajfVwp
c53BZbNvyJbfMiwcauPkZ7qlzKWBFuoC2vA1EyK2Te73QAaEI7RVv+3XagVw0CEBDzHrfNwA6UeB
eu5L+APcCmdg37FE5i39FtDqTk2eBcmqB0kbCK2/Hpf+WzsZ+Zr8/jHhmXVTfZFBNZD6JruDUnho
tHE5k5c2dDlv+x7LVRwZLezD16L0fUX1Z/xdvjINvMroYiuvnJl/h5LM8foXzmTbJXyL9UxgpWsA
471g8KCSBZ1g+8oWzbgW6Hol0iIpchnD69Hzy4xw8M4VkTv2W8YVLHC53xdsbBP8otU1ayLTKhYP
bWRrQ1pDYng5HaGNzLJrZ5oNkl9BbjIeRBJZkcsEj7A0CEHmRxqzN7f9LSHW6QMZUUL/xf845M4U
gfw4Ffk72OnuKPo/I5UdU3rHSCOLRJIj6ZG7pvZQvHyzzQGxRH/WRft8w1WW9y7f25kHj85o5M3d
UTO1/2CXEp+ENZVsavsQQrUD/OCiv+ePCr0GnwylCqUK8v9JzpyA6K0DriRS7CdsAe5YyHqTgVGw
Xm0KHTzn9ig+xhCarQBSkVYwkc7P41Pb+7HM5yeM34iH2B8wFL4fCKCd6CtVBjEStxUQhcZqYMzY
hgaVGUxCBmG/pc3P4Xs452DXfSUoyjgMfDcmGnLRyKDP6tM1C2IUSyX9eq0R0v6Ugp0V72jJ7IZp
EQXslqQQWHsGDZOoimTWDs/4G6IemnvLQeORulMDfyYw9vDFn771UOMtZK/KGWt7sfmKDS5jYEBc
FrKBNfWzBe5Ev2kYRPnXRMQ6T6w2/2x+XCK0mbM1vsTtOo2XdEUQgcXRI6kgbDXSpzb6ilLWiAFm
iDHJD3xfTjiYUxqNn6clc+OR0So8h3OPfQlcEkY/wJVJC/g7jFg9b+JtY1hktWHY2NpweVFAw6Yl
0oZFHDuK5z0HIQ4MSZijep2NRKQDaXvnMrv9yk2mcMUDPsZQZo84zC4VpPniYShaVd3hMYybATQi
mdJYGHhW7mVyMQud9HPGDWSfoJ5FyVHbkzwMECGZdxx4sBjzgSZFMpBU1aeTiJ9f9Kg04iWSXapH
w0LMR4WlzNBVUBn3RJt34w4WZ2Z89yoaHiks5Py2JOvgtpVGFCTpmfjaoZ7tJtrIzdWAw/cf6lPa
ozi483eLiX0lWDDbTxd3iRemAlg39h6z/THjrvM29tqaKqJ/bnSERhOmcZvm+NmcqxRZDep1Y0kr
tqLr3aSgdA387nu9rvtmxCNf1otfiZ13Yznq5qxJxEFCT9aS3ggPKo8riLiukAZOSCekpcMEyAVM
wG8J6JYwYBZzTOdPPZe6VfH7VUY8hDvMn+qK3nb5u8rRg/IVuy6JJnYR7lsZB3tHT1tuvew03Ut1
rcbWhCsmsbgnU5Jb31uqRHHZbzU9DLZD628TwItcDYJ1wdw4Sjhg8TXuMgVGyF+a//fFOBCD1Qch
ThFzIy4E53OP1fTJF3eef5TA4+qcI8oYze6DjtjZZnmoA9RP9HxnVqMPzypE/8r1pkR6H4sRo6Rd
CaJ7BEtyjeTxHTIQchVxn39LT3bbYorBzBszMUgtxFFpy4T/HGBTPS3HHWTcEq1d8+/IZS15uL+j
a13h9+AQytWMdINh8M7U4y2+zBd1xoyV+CYxRHNuSUGkJykl8GHsWqwMfm7UP+vvROuz3iotUExr
wl3tMFRyzIuUZG02OGnQnu/lpIa8IY3vnyrQpQO++fYtwarxtJm3nWs/abkqgvhU09C33Iej/nLp
WOQW+tqK6tMrGhaQoOTiYjYLozqXpATSQDZ3HjzpLMH7Zp9Yi30pQF3nT8xGwZ7Va6aot+95pFqS
FVoCx1l5MNXTNcGdrv2a3pYV7ejwPSOs4BqIwpomY6eZK1A+fDXb3sLYZI/Y+vCR4Ws3l3nEOf6c
gdsIqkMsxU51UmHp/B0GCvfLtsYes0BIrcMjlc9g2o+ZiGDqgV2pqbt1KHtWnFL5247KMxwlb9U3
w+hOK2n8v9ofu/DbsE1dPFV2bo/r0t4bOdmt8gI8X4hFTEppyM3iFGQwCDadthn57M7XzbD4BNGE
SN79eSuKvIJlwo3vU7MCnwrOxu8D46NJPROqZu4bABzALyb04U3ypc5eL1Bgzq8zKRZUs952y9aD
BuqfuEpw5q4HXUuc2L+YHqLVgDxdhp8pjMrQz4dDSClolwT9NkD3Byw3FZUH3SvyCKdy/dYocvUA
zD4gEz9ohg1XRI7Co4LKr7OcPN1eYUbAlig+dqhXfFAd0WTqbT/caM6kqBoAX+gDKJZ+Bm5a0r+W
yEPfu15TqSt14XkPpLfiu7AP+A9eWaZA8ZaFTgiCvHMuU3jyNGmLBT2kYLLMPDV2bBY9MrlC/gM1
FwdEli8N7dD85f3EWU5aufVmLVF/7pbGMp0TmT6x47kgC3IbuxJYH967nKJN+NlzD5CgGAKRuZgX
5EizC6mAti9iaeRyuHDQ5x3w2xaMwG6ciahG3mc0kmhNXBNqihGYwwWv+mTXACK/zMn4JfhDgRGf
XyYSXfYYXe8jfGg3Zu/5RSaW19yGj/zEUzK/AFmvb4lVHP9xa5e2Y1S8q25+tdsgdZDNUjkVyty3
VHAcnd03YC2VO3TQZTzPyC2YHn+1e+sxp4EY/TD81Gjr8ToVMMsb7ztj8T/82WKouJ9XLDs5lLPA
Tt3TKzvPIa0PqhY4DAF8bLDjzPkRIzSwjSL/BgO2FADT5d796R2iPfb3Rzhf/Q3EGpqZhy95vkbZ
5pCFUKO75gIFP5dvIusAxQS1uZuVQ1qiwdukObx1vonNAU07ORSu//ePi/5voiSNg6sCGxlefklZ
Ib/PsCEc1qA2bPhckhyTohq0rzX6j1fXzubIcXZOg9UCBgwoRSIIewjlU3PFKdguvwS0JNvDZSsT
T1jr0PNqXjhte1YG6Hc6VBTdsUBsFNFvd7tZ/P5VvWsA9tf5KO+x8HW6lIIFzjNvKb/Kf7SnyplV
mwViE5+Voz6XZtIGY4yEHRJ8wLLoGVGdtjjmWaJg3b4B0veDdVHQMpo06RsVa+2jUgxy+kmy8lOv
61isb2HV/HXvVnZWSj5OYL3g+RWNpnWJnLE46xjhL+tSDDj3BHgU5ghVe/0NTtRgl5m29FHSjKeO
Td50s//b6L6Tq0DG3SlIRWO1hfSzfET1Z0eJPRNUaLfu0mkTJWAxaM1IqDVoYliSZppzxMYaRONA
Jc/LegneaMVkp+Z1xAuhhW2GLvbwXc4px8jakkUPmrr9kxSY+FBqxgw/M1ok+QabwXl6qHN+c0Po
qU2KWmtjab5g/uZD3EkCTJxs7eERjxIwFXOepv2fmWPGBbn68MXRj8UqLlJzRkK2Xr5miHm4TX5D
RP0X3yhneP2UpDeAZi09WPD8IkLx66U3pocwjpSfEo8yXaN+0nULZL10b6Pun7thDXf2wl0STwsl
mqMyIJq0U5VK81dvdpwT9qCo7QgTEN0oWujLtEHxgrQWXhGNbGWlJbmbzOThYrCkKce48QMOrj9i
J1N6dVztETjoOTdZCuAsCpooMwTl3nPFafF1zCizjZi1ICmGaarIIpdRR2zbfmvY1OmkxcIVI7TO
6JZT7jF69uWV1CXtWJDhJalC8R1/e0UcidHl1HaJPfc7QrLmc5JOvyf3pb99/Bnll7MLKvIG3Mze
GCWEPC+sosY7dngKLOIgnzXjuQD+T4STjfdUHUXCNr/UXfFUCBRIfj1woHwI5+tY9vT6Sl7QWefB
ojagMP4uQD1F1bQfJyA48uhC5tehqsJP4wXI97CgEVsje3w2L9WUtO0nNWa2gp1lrf7h+LfRUClg
bvV+R9T3wqlXrEyLm/UvjHzU3AEE5rVD41139qnTIlUW04XeJKHGNV0wE8D+dNFGP2YoNn4Wj8Lt
uvgdwGfzDRxdjAjfkIy3WOWcXfS0ERfw2naCUcSMETvLId7wno2VkBmWmV8VjmGeuP1BAYBJSxry
4pJW97YpFLO/uCPypqFgIj5UqUP1V6OLVrHi1hxzMgF6tMZ2a921id08Py0J+++uBKJsaI0Qjv+W
pw68RkQz2BFXjhvw1Du4gax9FbhDGvg79lRzMrBoEEv0ca2fjF8M3+eSXfKJp9kBq1DnOIlLyO8W
zZ6qoyek/WfyLphkPKtpr+NglQy0UgFcpyHMKruhYqTf8kmDGVZ9UeQmWfF/H9RH7VIapIq+RiUU
wLBIdfliS7kWG2Nfto160Tw1feHc0wdc0ZLsPj+L31mFsYqRgFJpb3KmQTvng7ZXeBg653NKCyru
sgweFoYHGSKlb3ppAJfTf0d4G898Ie3h91PBgY7uw1fKoiGND5SuJodATInJgPmiMIFV/QUtgQNT
+6wQ2XiRQSvoIHTZCFIj5NAXsKdw1qyJY5wviyaET36I9WKozNONIlmnTAdlvrK40VDGhxIjntzt
tDsMSCUL6/UZ/F6fKMbdxfOQw5TF3LKcTqub6jwsCNiSQxW0CcdDTq7Sv9WFREHsY4TdsgUcgsf7
EeoOEEjwKNaP7uTLdiTxHplkzkocYO8nr4/klQlRC4ITIbzEsejn5J51KfmD5ZWmTJZB1cU/zRbf
hn240aoO5lA44B6JKyCVS1usDjcYAPIffBQm6Z4kbDG8ec6sbEYwAx+1iBqYns5wSLzh47twGthk
jGQqi9GeVdf05AXjwrNaW7T+gXaoapel5IoXgsUwNVn3acPZU189ORXfbHa7TSXC2X0FZaAHJqA6
JkYPgkFIawHkOZjow9uUE7DCqbas1v1q/KnFozxCK1V4iZEzkovLwBnNztdLuSM4Ye0S46UnyyS0
LcITO5Ayq+FvwNKOiELRoWDFl+350xmX4OkbhDLOG+Tpyz0yaYQea0ewldWPLp7sL7inCUOrK9HK
v7h50iE+rsaIC1w0JgodwIyzbaytxz9XYqDmJgxeuE6pQ8I71OpuGujYSCrjlXzHYjXUpDfHlAza
VsAqSjzaF3tOM5O/uaazwxXLCrz7i5mz5Ar9b86gddUhhJqzuSM4ZjugPbFt8DAEfqpcnSopkVlv
Xc8y5jye1f8FSpfPztdguHECL1aKAC4r7Vh2ywZcI3CTtfKRJgIhXm+VmvVwannOpoSLPb4B+0mz
8QeeLsAoa5D7jcClNgokoyAEqbN1JNUEMhY1CqkNqSjrNU0iswdE/t0+geJHDnyyRVQHwkR6xQgv
veisPSkWb5BoiQbpf3A7DNMod8sLnj9x2E7pLo4jOxT1ekvvMLEfl0uT86fxWzlwnYPGWEwnuAVv
SuNL3s/ch3z3AaLlg+WqBMRvXctSXQ68TxtXy/JFUPurnq9EIJa0xYBhzim61NhRKjaFtXesIrPM
L9hKHLt/2ipYHtszsSKmHeGUux6DbEU5TATt08Q02pnoz8Yv6glEdH32vwHfOXN82Wki3huwbRTU
+dggi9TkhSE7A6WQAye+mkJAF7icGvIxSzM7cHg88pN/Nm3gBRWKS/fmI63MVR8XrapGp4iQQ3g4
lMIPJhz1XcNViVBoAGKx+s/9Vvg0Kf1d/LdtSKNxV+atiyIeWIgVvvmuGQWtF1fEWWq91bSnPTCl
fHH21zVqcOE8jbMvQISdm2WHzRZDlfRRLoHGs/L9QpW4yyHtVs3nDw1SlvntyoC2Yjt+xuxWa6vn
vm1kpPuSeMXNsqmc3WTqUYytNvZyAg2Ruj3uU1zIHkfI/T+BB0qS+n1XM4npJFc6bi28QQ8yYIrw
23DNyPGzfi6cZUaUCgjV9pjwua8poCcpWeU6qkyIsde57sVDAR/RfTz1TcEg2NjNBj+0Fq3f+CBz
4OVD/xq/Jd6Bh95yVm8Q6jVtBN2Nu/uWJwWWjmv5anHEJUvkh+Q1UOjDN6TKGFnDNzfn0v2PhgW0
IK+FAy9vPX3ffc6Umd8U0cnY9SIzs3Im7Nyqb+j8xODw3Ofd9bbJ6uh0qYbkDkmcu0vyYh+3/zhQ
DawL77jv2VVnS4CDHF0gjAJ3a/LLHreQRBrowDu9nn54Z8yIWlCNF7JOaIq2RHq2ThsOPM4qzXww
e4qvcymhk6ro1lS8a9W6g5hid2AmTY5ABOJQl/dtvfs4mTZLFNQBPBTypGv67Fnvi9hRirZ9r3zm
t+uXNmd6fg1CdEF+QEBX7A7b/zyTmpaZ11pP17Y1HdPGj05Qc18gRK6VszMn+4P+MsFzv7FtRUck
zqs2Nax05MnKk5l49A3bQX0FWzL3LwkDbCAyquvjErAL+UFZe0y7K/TrKJZo0fCNkTFz7bSWx6ZK
xJ/YMGniODNpafY6yOt6UIhjmv68dsgctCIhkoMdhtxuDe8qd0Z96LLIuD6LE14SiLsI1H03eMPL
eNy2ZeFsw7iqO/SkP1Jdn6vp6/k/+2FwmqBsDBMwwp0uPnQtg16NVB97+FNzqqgFQfNR80qVTP7I
jrBy16/TK4X+C6rsFYoVwAFyDk4/t28iiMg1+/IQGvOH24xVAOLjn+DomTj1MrncZeJ2hLOPAONw
njKaj2eEjLOrmPbpDZm7zw9p+ILo9OMXd+7WpftYhbgdbpVxswsBAQkHBfR2l/6+6nuWU3gdgXYI
pqrL8epBOEILbgqXdvqgRtZJT2U31lvjZeqFgJ2r0IpNM+B1zzrRcnWxMTwSV/leppraLU7scPrA
9G8ee1Xq6EtXn4W5VZXZVQrjeLy1H60K8WYxOMag66Vs1eNBSNUFruvm8senvs41qut/lgggKupA
+EsGC2xXqxfAXLZpssBbfazBz9floW+UlN113vdYT9naEjt6lFHBQEdIZi9FUKReI/+SNhrA4fBQ
sMYjk5iF1oxnhW/U+ZUPQz4HrEDPcWx5vp3NZz2iZS/p00iP6ZMMZVPBzRT9GAa9sO3lzS20BnaH
td7L21Wwp1+afor+5ZyEExSY0jAZwAe8hd5FsnewCbXO0Eqw56O5kM8H5zvZ/xyQMbwj8j/B6y40
s+cJfWz+6Mtm74bD1JRz8Brpk+pGLvKjsT54lm146TCc2O7XDgr9G5vB6Fp1QPgwzaBL8awJPydn
I3PLdmvkIjRbeTgHpKYawG9L+ypQDDcLyFBvO69f0f3aoqVXiYivVcPACuQ/dT2GoKR9WmcWOV8m
4fXJGqQqR1AN1/+cMBXlXQKxfNLTopzysc1tdUGTyhJ+IRVZokW9TEXiG+iI+pw8cKc4Aw23l6DG
sZg3+rpAct1U81YCTQ8wjW8vlh8ZCviEU9t8dOFY03ojGLZzclCUQBB0RYgBQl/Yg0/+l1SfP0p5
A6amBK2PxlQ6ZFyfbZMOw5AvSMZu38KpelHRVRA48+aWiCXUpTG8QzQJ+CLfswNoIVOmfcnzwyyi
8SuHXUeQ+Ghx+BsqGkwWN9nAB6XJ3/aXYZOLPl5DFhJT0u9s3Oh7yGIZnonLv5e/ReH1pkSy4fuN
uJZ7sVNV4cdj1EXk/RjEJkyK9mNEMPAa4nw1pHoYegRMudZ/NzBQqj4VlMNecPpUlEGRP/Q/fwK6
vvoqQ6oN/8HHHSRK+DlmIbUnwfqfsCQgGiyYgiRXTI8gNR/4aE237OoT+px4pjhxqAuvR1QwH9La
j++86CwvEssDcyGxWxd32IR8QjBKyXmBQlk+QBYZ0AQ3opBxCPDhgs1fk8sYZUtnM8CJUa7cdaXt
Al0nOjUqqDgcjCemARAnM2hGxBbNGcLvB0OJHvIjLiZ5u7Z6l4ueQr8C7uEEKVfddR+vQpwxTblg
YANScHSKd5IVXHEweBpssxQQ2nztAVO/cCzh7+7UmXjhshLwLHI1syUoPolUBxB3OAkF3Oy8adaA
ZgBTJCxsB3m7Iuq7MMKPz238Xqt04k/DbdhP412xpLatn6/WeUk1s+UwdfWiCgm0d4GC5Qb5tEmW
R1voJvFRwT58TMSB1JCc593965rzyXAyb05Ka4UoZfIhNBVF9FD8D8HqqATZRW1IK9ex22oOwHxt
L+JgkbGJ8t8HAjBGA5pUOhNxrbQgAtRKIdSyZ+sRWsUGzbUIRZwnDfJdyxpxbkl1f5b1vRoYSGCT
o2xxmLZJ7jDsoElcN3xRUWxchPcvWjoNEWi/WxVA5GT6SURY6311wkfkPN+LtOzsw+ECXaWtn7Vb
zGXciGqabyLwE9GYWIk4JGcoAjoITiLiMTw92ufMmisFuK7mtDkluvOoiAx62EZAfzkcfotANUv4
S+HwYmgDqkEOi+63kFxIMbWEh2BnyhXJ+MlCXkxZ2AXmeeTwL9L81vc4d6qBL/x1db6xE4Gtcdpc
B+S0R7KSw5npQEcjuftrLZr/QRV908mEt49ApoaU+zVz0542dS29J4bGKVHtHYC7/E+sMXt3M5Ph
FyfjQCDAkdQxx+ie2LlRReu76hp2R3fVEarw9SkJ6WdXKyEZABlrZge1MidCV2rYIwKDm80VMcX9
tugXtCeFHlshCQ71GcF6lWYM+M2ad9If9PYTtZcu06w7koh1oQx8mpCN7I7JtvBTNh9tVZoffXsL
Fp/MoihUdo1E1CLXriRfCDavViP8rtRvYiAfcClW3cJ+gLQ2SBGeOgT5JUYtr0PPCCqcnm0NQmpC
pvTRL8jFOdN9CrzPqKou26VInMqvCZ2pYomXEtvi5eBaI2siPpHSi8157SS8/5bVdkj2ywnLEyND
25bkjVi8c8UXfFYupNkjfvfz7MjBoF/efWpk9OH4RtHGMkKvaWuPa8cYWfLspdy2pRqO9T/Kwcpt
u22GbwY6oAl3WoRKmcJwy8jiG7zFpVPXXSaWuM7TvQ06BqiSFAMkWyBoBEAwlqiGOUiJ5IDK5Dp7
/xprTJ3hJcQYGaUi5xlrv9UWRlNdhaqfJj5NTL4qTD0ETcQS7epM3y4BCgahjA2ksfnfGjF3M7Ab
xMZiqkgJngeo4RjqZOhtb5Jk+nwiMgjIh491l+iXhJFTEtkY5D16sh5spHcffx7INK1s3OJBJOqo
GsnLq6m/12zcn1ZtsNVVsqIDjGswoR9cL54CaBDL9vxFmVQ4IxLDZxKAzPKQ4UwUDqe0x2Z1Y57P
AvtqIHa8FZsbMagzVjRg/h+X/YJCYWJxq8nw5zksvvkeBYP227ETPTrlooJg4zdgY1PHgpt7Cs7Q
l+GB866sS0vhrY5Rd0a2Hf7SMR3sApSlcpMOBs05+FkcAtRTWJvTo5b339DjM2yKvBr+fF7Sydqe
K023uzsFHDCgqR/xplbnev0AhuHzhvnpcbb+DLLu916SKulim4o7F23BiLFhaxI+aeLFFen7YfYx
6U+5uy4TOvetGgEFNtBZasOwj6H5lkEX/fdn+b30w+SMD+NbSRlxBLcmZQskRKG3zzEIRxPnZH1R
ekj6Bw8fYax++NbsDNxd8RjdnLvOGjXvq62Ev78RwriMbwGq/46+isdQAsifdpCyZIolyFYRP6Av
xz05vMeIHJDKOf3ehYGqgzcfBaQK549yvXS5d5JYMyHy3uw+QbuhCQ5K7P2Hxo90FQKRONBpOOyR
9b8eacVGq469tN+ImI9/4iI0ej6DalHjBF6MyVXfy1wh24vzmkD3bnT34pRIjBVDvEvigLnaC5QD
g052mWbo+qJO8c1LeQdPUd5e0UY6Cyd7WU4HtvMuCnUE0DnN3VCZ95mGpmTlYxKW0WcGfuClL7bY
TJOnelIbiLypBG1ij1J/SIwhdwLWPcsYAf6mFycuUmhwXciLi+/YuEg9O9c2diAQuJR+6I4QQgAu
hmZdGTB4J2JjfOWnguekpqwsS4SLMFxZcTKWszj5iy3RCVeD8kt55U+UeoTWuaTkZj0dRsb5aBJV
Lh5b0rRaN+i/f8RLDd2fl4uXWb9T64PoibzxBkyYvfK7xu7AtvRjcTcLgBTCqGHnRj1+a8nf5lyH
T0YVux6985fxQ8JHLawNIilHsZre1IxvCzf8NXyoeVyZqwTkdV3jkrLY901CNvxYRDhnxq1Fo1Ss
BIc8hgYEqAAxy/RMdoD8V0QRTyP6MWK5egAbFiCToNVDu22HD2jtnnbcBuDFuBesRwbIxA3yv0df
8yLN/CxlsOx2MMd76rAfQJOmcrSizpqtCtkFYjteYcRvZ4EWe62+HL++Y2xsfsK0t+UCmoI67yix
M20pqtaRmmQn9JJuYcPX+epvcNe4TCLn9xWgHKWyc/eYkGZ3lBfaeh5Pow1VpWDB6uLhaKkrHc27
POhE0u0hAxTaIQBaD7UhBWOkZFUYkg1ekIYE5KiEXAVEK/0r3QyMeRLvEnLTu5ks+9LxhnjktwdW
xSFZqBoyKOasXvOBbwx4LIrfoD4issPl4qqoKFHv5p0XZkn2dQMsapQh+f2pced/A+FQeQrjscDU
24DaXCnH60edjYXy+qC2y58yAiLSq3KNpw/m0/QUBjngfCVAY4SNOhbz3abfhKQc5psrEsebI6W3
3ozwfp4mNvVnRFEb1qeZnGaix2xE7rk5Dblx/PQba8/pbWjTc2C7rOBpEIUBKM9xrszyeHsv6XT+
CttK+op6lrTnpR5drd7/z3BEpDbGA7yS1SC29rPzfhLwQyo8I8ygDvDgsJMKD3emZJ/ZrpyPUpFg
Oh4zOxrzNaI4m1PcRdSq7jSFE299O4DGBM/YLUjQjszdu0rEeJlfVgGrMU+TBF7AOhViodtp6A6e
M3lbG8/3UWEeawQZfjvk537NR6Hqg3PELxhUFi5GXzkgpVzAYEhnjDgvzn4X7DMek8K+6oxHKVdm
rf17gDiHsToYMXJQHsJND8jH+wLND2erC8Akgdw1YMEnZW9vOaO0WAdoYHfPSP2V1IhfFNc7ZvQ7
3gj2au7nw11Db8fOkI28MwXLfZxgKyCrndXhwsYtMjSyZvUoDrkLeQq6UGUiLPqEJjXQ0PVe8j/m
IXJ0hmXpXVDmZrHjBE8w+XBCIsk94Oa/dPSoErC3s69d6lJfXdKzxngNdtqvztwsZYOz+eUat6fN
NL+9yUwxzx6vuYevY014AxB7KM6jkrKtr0UNXA0hnDRJqnIsJMwSD0fYRDPW03yhKmPjRjyLPksg
9SYRGF2X9FdfZCa9Faf7stV/c9ssTD9pyHLwjeeg1kGI5SaAZmv+C9KBm8i9vAzy2UtuvhO6yRdD
SMlCvkqm56OlDzqrtZaJP6IvH+CbwfttYc49kLQFwaF9M3uFd2zWe4Bvnu5CSiJrka7WaqPd7pEJ
J/zS6wXohhxxEzWdKN1gckiZbp+t5qtesxYTygWbGZMz/VpkA+0bSIMqB7emNdHRaZnFPi4APbh4
iXYzyPuzof+37PbtFfoqvzRoT6AKLWuFFoHP+mB80CenkQ8bKhelDeggMUqvN3QSry7EB0kbRCpk
Hmag9GZVkcP9BIfxPz4gqXC4angVcC+QzcIhKe1awI0LMh+3pqGsIflJYq3B5Uso1hyAB9ZCuEsm
mwx1jggTHMjHipAF/EYpfAyCq32rY6QLt5/DcSxzEAAjHLqvdvAnHDEh2ISnejBhneRtETL0/Jym
r2/9UrAoRKyrCY6gnKCH5A5klTFG3tq96xtnE1G6/2g+2WX7or29CkIYJnXvnvckgRXMbuqQBnWu
beVY/3cdHeW+4EjLUKKzmBun/8k/kfUY79IQ4cm24444ao5EBUBcK5A2+Ia0Ws5Fmgzta+4TARXF
qZqkwKdYf68CL6tHutf11l3PenbEEhp4XphJa7TQiueqHPmqo3//QVNLCFD6Nz06ho3urdmKdIQN
ELwFVJ/vPFPWvF9isK0zgQvyxG4OaeqRldPY+qOuXjkRw/PCD0BJ62pDiTklBUFVPwMzW135U850
YTBEG4hGTH7ELOZkDbnplXVG2DbJfqXcY+e8n8VB6mtPCv8ky8TK93mCZn69CjtKgRTzrHgtk4Wd
z4LO+sFoClmWI7M1gKJuqtczum3bKnnVM7/onxS+Lbv7V2gjfss6f08VgKKlBAfufl2m4UUj01Zl
9JuQ52W8MKDE0vr3TsLJIfJ+CGiyGhICMbMqq4neOH7+zRAef9s6Of5v35tlAKjG+K9Uby9XeeIU
Ddex3lVb1VY7dqWPQWlHIcnLQ+6//tac5R1wjJIkFaHf5neWKfa5JUuQuE+AkpXPCg4YWoWfAvXQ
7EMUzkBHmL0Qjv06Fod3YrHwgFVjxqco5YCu6kVgG9AmZssAXWsI5DATDe88O4cL5Ko3mPbt2P+X
dxJntB1Cv9AOEVcUihAEkEdbwr+Xjz4NPUDpRGD9KPpgZriE1cKzCCxeLk90b5/u7uloa2obYbrR
adIpRUzGueiiMmkCfH/BNAsFWCBLRLzFSKS6pxy7UbRfQCqRxB7l2+zfwWXI/SlVVVYlwtPlUywU
r8sOd4fULvd/BlriMIVVgAlSnefVP/JsRkb9RA+fswT2rIpd+rBM7ayr/LrJWsKOG0mHJROf0gAo
mJc6HYe+7h3HhhfZHtYHHEqgiSwpilzNWgg34mdttgMbTsvYY1rn3eGwvBNeP4ysWJTC++gWa31b
b9U+w43CwzqzjCJf27NlB0677w/eXZB4CsjnYX2UnOpHJaSE0/bQ+cKp3YSHmNKgkvO613L6uf+H
CQbaI+IVX6AZsoOQWzJtFUvZLNswj+hUdNm2UPenu5MzaHEbWxvmawnQ8ni+tlWEeKQ88BKJZFUF
c1AdntQO54MULTU6cpF6UB0+EkwbPZoTpdnSxlGkVgX5aDPTld/wS1FVzXRmVUezkucuwCJqJRFe
oYc3n1bkWKSmSrbqnTxzWD6ckuWOrm6PCN05qNXm/Ew8JMPPDSpaZauxlBubduZI2bxfCg/b5Zly
pr4dOd8x5qQGKe4v+dehP7XzDgr4JcJYSsVYb4zn0loKVS7TAPSZoTPZkT6KysxSRujSkVrNGK42
3vH+UgxJWTE63mCrAwyGnqKHqoKUtm3k9Uuwrp59nLZfwcr8gIFrtaFfvPiZAtKNhgcv63xONWU+
d74dkQnXfzBI35sJd0xX1VPtYnK1fU7fOCxjHq80sRtOVcSnuivUqNJe6TiMrmQy9LIBKelm+ku1
ZwRJypCp5AHvIfa4d2i1db1HW22vXbyA7PZ9VENbUc/ynW1CueMYyje/8FCL41U3h0VStl36MOAB
xq6Sv1yv3loQyuspeCNr2bjmLyB2itwNdRMRlCF1wfCBdN5z19ayBQuUwj047t2Gzf1gfa8WuU6t
KjQXtUZIWYlCqrBPie/CSaznO9QH+e4kb5G2QzzaYBVCdcbY3qGRXoTXfLa8QKNTS5zm7v2xA6tP
frm132oiQVBIkBp7PaojeOWi0R95YMewpREarGAgzt2XCg9jD0RhHlB4KdJWde+JLR76fwgxdctD
BNi8fmjOXubMLxtjcHrLpGr9H0eOIq5cRcvVruAFcyF8Yz7z3YeR9dDr1TLnHoBFHYysg47VII31
NV/ktTbKM+WhE2CR6rKtc1wc83poltC39bbqquHmLEwpNuu4QCB8kAkccA07SLIuOBFMyrezTR4x
An+N2i869xu7bHFR1bcU4qf6B1oBfHofHscT4W/RM//emLDnNW8+mSemHX3oEUP1BiSncUP3VjDr
nwxTbisoQsZJDcUaX2rf8gQ/ZLOMOv8YC39LkZF5zYpbaq8Cbv8FAqbKjGVbWzUo+G9+rXZWxNBG
CWD7d64IN22J/HjCkjDNvzpjsbj/akF667yoqKsrm0xEJUeY+kan02454k5+cFix5bnfxFpn3GLE
ww79MJTx2GVmaJQDfc7Wl3eQjBKjGYcEaAoU9FAtPTPIlIddIhrDuCsSoWrcBSV1khCQVtUdnmS2
8+rP1WKi5B+qWm+pgXacvG7QWNWz9yfjtvwsUp3enOyu72YTke3nKTjtm9vN8fGwSG5IyMFT9wwu
3fPf44iwSPGa1h72AJbx3iqiTCsRETuFZcKvuGYCorBlO3OhTmH2+Z4WKEY6WWeG7DX4zZ7k2R/8
57QSy94aQ/YUHQHH/1M1oR0C/eb85BIJ3L+JHKo43gYUxQkt07NtKj0Z3eHARafoR3qbcQz/Mt/S
81KdrNP2kptp9AUIlMc6oEd/cqZc6lO0VTv4WeH2MAjSfAfcG4HN7UZh3OkvVQsd2qA5Cb66curS
db1s4PXY7gJsVJZfXtX29qPHWzSO8zlUoIFwiy1spf8nyCXN12F+Y0ZmxRt4v5Dm66H9T1t1blf3
J/tJe+fBJ82WcatkiHzIpkn8U7x5ncXPY0vG6TL8KegP0ouez6lhv4aqcaF7wzGXKI5t1imweBrI
5jpiSs7nmritAhmpatBugTQnpP/9j00aKkT1Jp9OfFrLUv2IJGvDL/H8K1946YzUCEbBfbFRy3wV
Xw1SZOFPx2nSJzEJuAT0LOTGad9E7b/zVUxNcMNqb94KSY2ZF6CxkdUHEbGqiSO6chbOqFfNmfKP
KXuRdWuPnois+uYPlVBr50uU4aHZshc4IL96niW/tn/9dfhfcZ9Ypdtt2dbtj7revykTTU3hR14m
wOpFYAKDCvBAfDmc/sehVRHIbMXrZf+Czoy7eZb2OjacPkolQDTdLunE/ODoxq/S03DYCb/W657J
YtvFbAtpGkh5UJSmAoPm+77pATi5r5UFqXUlUG2SKs9s674BMuiHQ+DgwvNYaBscZydeu4zIaCZw
j48MC0ZLi8V79Y65oE6V3O81nSi+M1bsyrUJX//ai/ue7IkB32x1AvEz2xrFQALfBXchoiOOiTwR
WFAGdGfMTsKkWfqUN9i1oBgflUQ1GOTNPsfYzxeogwPvYESJBAFJzXS5M3gVsz42wAXNm1esVyif
Qo1ujUmVLT2gnJG+ZmuepXYAfqbR7hzp2/rZZUQRHwQ/JrFMpP75ogZ8DXwgaaTQdjfjjKqW3WN5
BY7Qax4xSxLlLIRq8jDV1C/fd3px9xBRe8Mbjsu4SNIkds7X9keik9UdOYU1rdP7SDY7ft8bmJ3K
vPUPDBBLlcQyfi4hJ/alfCCyVRv3JMuYzfnUTRW2f48xXN6Q3Ya4Ra+nP0kmL3zD7Q3ZQLWyFLdV
3fo2Tr7x98nHAvwYyxlujKvyBA5LY7jivvP0l5EfJgiIAyYL4bTYwcc6qyQHg2iF/vGhzjLBqr/y
xxdpKy3o66RI2Z7gua+HbzUIT+L5RPLJWsopm38+oyUhrQFam5JDTkxnLQ6HXimiZBQBihuxpmTJ
uvXDiQNROoZBqeK9daneqs5h5LNi5hzKLMqHzfrs6mjM/COZ9AB0oCOPa95lfPQVfucoZZXhdPBe
CIuf4Lk0OiNTE3yYAacCm5Dz5sW2Md6itaZ+qfoe5dTwl2BQW+w6/6gnMk7cls4PogKLhoKukHri
/Wconjrw4jpMsiVGUDvOPiVzM+k5cHUyetdtgIL5HXIJRXODN5E8GonHMVpXashvZuZwdxiRu+uQ
QWVk48R87pKv+955UOBE23a/+M0wqAoBn/A6NH9H8y6Oz7x7zHTKoFfB06T+6zSA3GRFr0qCIQDO
+w2wu+hCpKx6yp2RjJMPPmWwlmmRcU83W+Uh/MXErEdkmTpP0COBYio8SFvhFN3lIHckQuRWFO23
OXkT3MRs7V0rj88EpFbSO7A60AbtwMkof6umSPYvqnhh6ZZhJtI6pi/g/8JoED8qxiWpaV3f/cLD
2zE71WDIE0h+Ec+Xiqj4lGRKoPlm06+vX7PotzEWnLlycLZPfpSFuuFcVkYM7Tlb4/E7KfuTjI7u
MLjMPRStsXrP6HKb9jeIQFsZxMZkT5fVeltFJS08zmeehb3bp2DbCdRHMrzj9T+YLFu6foGjlKR8
lncs5p3cEuknQRlObwHGDT2+wZGEsjPkJ7zLCwXK4L/a3dpcPx4GK4KTsMWlbjB44Wdc/MZa1ZvO
qegYnSj+f+pSuVgqNs8sy8ipYgFtIp+QVbFtr+uHGt98vcWG8C9rp33QmgTf1Nw8iBftVkP3jiny
XnCOXVzugJKhJwnsLoNOjpl/FL3XvWe65ONfOb3B4MYyQKlpwTgVnyzMqVHvLbiQANcevRXhFXsm
MKxl+HoDVG1jWx3fuItU5ummvQfS83+Ayu9qV+Hh/Y7KMafXNcZOnmolANEYcHu44Hnm+1hBCJUH
3/gy5O+tBLvg3AbXpXN40e/Igq5O9XoXVIftRmXmuhDIohytjLwF6OLTKksYwJ/oEX9mBjdzTZ3Q
cNz2a4qulddTB/ZZegoUPh+d6QSjGM74K/MRHIWN9LVg0tTEWRBZm6P3b67CaidnBTAQpR7eYRE8
Ng19QdSVPkwyNNP4KFKoTec6ElM4OYF/nLjc/AbtE0VElWNfHIvbV4N+bramQoPgfahS9qlMrss5
kusyGLB368RfZl8IHT7k8DALPHI8CXwuELbd3UJt//nUZkvzpxTKCcXM5U2IfsgQFiCkqZS9yL9R
4fQnVdqsE+5nxLZvvfWEY/JLf+sZIb9DwnIPqdjje51WG7g9IA6dCUrmB0/tsCNtvVSCH0h8sYM1
BRd5wzv61C6K2hJjxeU5p1AIg1reG3T27kwA5cim7FH3eOHCepaOSqR2+RAZ/FxTugY209phaIZS
QWltIkeEFkuhwYjWQn22KqWKOxr3S9mcZmeNYCbSp2XfEgayFkwOHPRYoPgLik4dN748jUPG1Rqx
mSp83krSjjekI5hMIMISWm5mrsQ376swNvzFi7vFF0jBXawzqCarMgp8UbEgvRG/6oH87Mf50R5d
js8gIPgi413Hm4GKO0+gN2Q3nZtaG/EE1yylV5kDpg/qfj87HyHAPo3EKBPX6jS2jVtnIVF1lD0l
TWu/66/oBuNXJsjXcvFGbK3gcUW1NGIT4sFJiE7bB0A2JVfwAc9lGyeb4WVLxOlj3nj54Cz8XTA5
7SGWFaSwYPUHYHjL8mYV4v44Lj6YxaGt2FuwwLoUdSxHgl8fo7bIUVGbODIG8l9CxeEkcqvJcj3w
OWg1QMp6q5gqdxMCGI++NBQ4gvDOzPylTv9Q4UMqmIE1Udh812L+anGDx2MxnCaHcwk55R5/fCIx
ttGzt7W5B3OTKRGcf0eBjxb8Wf1xorrYls1CBBIemNsNxEZ7Qv+aiizGShpg7aWhKFI2VnLmblU0
Yy2/nR0HMDJCMwtSGP6uvDUwx2W8h2dcbTFY175dmHwFR57FjxqgeFFDSbLzusXFDRS+nfezgR8/
3Dr5ZRLkt6evZWeuPhQJdhrDI+chtLjpcZ0lHVUB5hezyNBUUmJ/wUGiYOj44TAejx59edEmQ7oi
v2BXGjWNDHx7UWsLFdQlvo5VLOUqRdYn8JMu7wSuEfAOKzD7vTc9NZu7SJkZJdJgxN6YDL1pliCX
wswwSIJgMN7epTKU+JmYx+X7gLmugHVw7DlpwCoI7jJYEYbthZLLMiTlVohIePxdrA1uTUdijjTd
tg9L4fj4VHW12re+rTaY2Kg+ksS4hoMFVo8OW6diPuzKBgls1X6nkyhpGh1gxfMST0eUb7YQqh6n
35Xm3oBCYh12WH2fIPgXYvFimswqe/kE6RoIF38W8ZlPvYffLZr1SAHiSl1hvrYqGKIWLRXfHA6W
vYH7kt3HJhL7MmESqUnXl1LgRnKgzjORGbjR79E5yhxGZG0p3o4s7YSSdylBLiDov6IAvI1PzdYy
hyoZZaD3AHeWC5W4i1rBet3nQngPfRcsN3CIx4Jz+gPHQNylvE+hr1OQr4OUTu7oUbvpGPtsocxc
oogT0X4c35VvmfUqgXM2G/F7+zZGpaLgpvWzb8LMVXhdRlYdoMkWhhGeqwqo2RHmAw8RZNvn5st8
MlynGNU9iPj6lLu8KGf/kgSHAt4jihzuO+gyRT/QOeAGAHLHwi7BL/jkMerxyTLISHZsJE18QYa1
ZUw1WEhcg/w9HTHHVrYDyliuusDcDUyZijm/X83PjDRBqDGuF91mpJZv16AeNUmVZVOXiONj13sq
yjP9/rUFJZ3u5e/4dJzQjp2QelcI2PdBJOJt/rCuL8f1FIh3qjMBlai/faOTjycOgxoknbnne66n
rRuLDXrYIsyAEHDEn2t+CyoNlpbOscyKgJMgsKmOlEXKiiHCmCUQ+1LDNqxAiQYU+aKAaEBMAfyT
WK5r4curWzVBClDQvDBvt4kewBdZ/57zmbymxk9uR0uVL5bf012a/m5OeTqMPIrUNX/F0mbyxsGX
yyuWTfmGcSAKX34aenlsL9mgrGoV9OMJuReZdftwXSOlAcjKMiwFyv93UAT1EwIPUUpeYw4xcXpF
iq06ymm3l1tZDYK183wX5ZoW4hyDJKG/4Odj7wf89TPZxGC4/XMdm1gha9dlH2l8G17Un7Do/iOE
om8PyId0WF2iYff0cqpi2Qm9SP5YIpw1zy1EOWRmfcs9hkt9+cchgdvodC2PajIOju+A+B+j64lB
WG3N+ySRf55H3c0GxDb+PI2OValJ911QRfRvERw6qNI0W5pDUeQ30ketkDNKc4DyxWcdf5vSd6Wc
vs0jJ0/LObO+2P7slZ25qITA5NwBBfBcjCym62z/zlAjxrHhmtKlE0kYq5ghPWewX0Jbi3ohDCQt
0VNi2J6TrTgd/t6CLNDil5/7pmtPVPyw8aCKTz0eWFiWkBcAvZB48TQedu6/nNq2HlOc6GklPKZ6
zID13iXvdqM1NuAW4aQIUIGoxK3CiTsH1Ditc/l+r1E2ba/YGOkuiU5ofpEUTrCHwFFjwfngZozw
f9kIO55prfO38hyzbMep8agklT7xRIrEPjAHj6mNFZuX0vG6etjCuFBewgR/Lf8+ZAEQhjBwkHxT
aESGzODKSedgc1BB+Xv00psSh8im5zsZSJmVtfGMchqbcLc6IY3PWF8TD9KLsFagcTKkw5SiKB1/
dBgAmKE/UkWnafhA3NsSizoY0tgth7AJ3ywa42uPBsjZtg/JxzlymNVaZOBuVinZmRIFVy6ebW5t
kQly+lSiEco0Nh2wqE3vGgm9LGxsjPFZGYAQ2lMhR1+OyA0TYKZo33u2HJFba28GIRnpmM0qaJZ1
wA8yEcSodtDDQayT6MetMSe1cJ1rHd7O7QxTrI6PbDsrJt4JrYTM3qoJV2JT1rO5iKMUgtha4aV5
/ie2VLCYFG8Em90lDF4XNyLmSiI1g7NIQrI3+G+KqBZvbrJs21G+AzWJqoAIvCZHWKHn8JhW56nc
G/HvBGhqJzob3x6qJgdSjFkwaa8fgPPN8icMIUqgYXHZ/sPeopBxyGShJu/msiQoT9g2Umx2AWjU
0XjM3vEywpgb7BVg7yMOg717xJOtciBIT4wru8hZpBXTd5vs8NPQc4ofqOpRzj3VbmGNma/DV3bs
LMvRvUMuElpAdw/MSk27Xg0P3IkrstImYLldXfujS3vYQSzBZgulijv+aBtutHgVU9cl8l1gMhew
PN3xzkK/kCNzUN9/p9P1kFykIW+CjKvEpR6kAD6NW9nltha57J3LiBkXagRLZEUGh9nmqUnrUGDo
JtN/xaYDIVbM52IHjbH1R+AjKpxOAggNuQZiziVutcfXzxtXzg9l0Kq/wtvxV0NdqDHBzZoKrtku
JM9Cp0nFkU1NooUmb0M6kyew9J8B6htBwp2a1Pzn5T4Hh8ZrqQhl6zaxD/SHZUEjn/JQUsKzzxn/
myGHCETOfD//c+Wfj2/sQXg2YjBu110XMc4uMgrXVsjisK+jwqYGEmrnBFjp+I4krf33qrAz6QLV
QafC1U1I8dN8NmJpFqrgMrSGpPapXm5pxPTLWgoLmO4wETWwFKfXgus5FM3/BwNdxbSn9APK3roA
dVLMzVgPMt6p1Z5NVgnQrhnOOFOPRj+TAPizZzd6hTl22OjaCRNPwLvW17K/RFpnISTx/ZtIhAC8
o30H1eqcA3+t4W+JBf/My0ksyWocWOmkQFXsxuCGcdLQrulA9M4vVNGmz6CWmuO153KcV9GgCbQv
dfMFK7CkGTvSiYMAWoG0a2DqwGKGlSmf7rB+8Z4IObtaKboKrnuvKvDarypHkmjGw9eSxSQhhYmG
AMAeXqLLMYvSqnV7g4bdazdGwFVa8nk1igITpYX1seczGBOEr16W0HHSYr5siybbCcbmuD0A4E3C
/yq8RBcM0XrZDg/bu5HwYOK37+7TXTUZTAR3DJXPu9W85o7bI8f+2+3azCwxVOi3FGCFSn5TZqAC
YFtv8Dbi3yS0PopwbmbYYh8+FC2LOabiMhVLgfJWkFT55oV/qst2MGhQoAjomIuXwaQBywrP3Vzf
jy2XdmZQVLuz0KtWG0KM75NLbM5fdoaApkKV+3mLx7mQ6I39bwxyqVJsUDe4TJj2bJh7Q6p7n6x+
t7E0O4SVqsLZutkC9EeXA+HZiSN3lC8Qs038Zrh6qEktMBRFqCY36Au09je0igg0Hw0Eoilby3un
sEMWL4/M3YmNXQGUlmGkdj/CvUUmlJCHuLBqBs4rmRb7GG5HKpQ0JeOOXJgSOIb1Evj5JX4y4LfZ
6VR6PhKfjqbLYF+L+nwpfqyaYnioVCs2BgMsKD7GKD/MDOMifWhD9XlYDKExMqNyTWphFMBSqIIH
JKN2QQY5saW28a3nYpBYDNDYn+PortQL0u4cv0t+lATZ1NGBXCjfl57kMsRBWP5bmKPNHzVFJ1TI
30jQlrutoUBPtSY56mpsb87CN8I0MW5fllGnC7X5AIJvAULVBht0I0Ju8vS504eWpArlA54MQO7T
jYQlG79OY4QFRisk/9rZDu1MheDuqzmK5YQIFqUrqeCfyeMP25f7XUF+VCd6fgQ6YzD7Rzn8Fotb
P9Ce6dO23R3NRokHupVLc3CWC1mjkMGEVLC7dQPoauBeAC/kuS1o12DKHqAr22icTw/BPa3WMQL/
5WIWlk7TyUrlKDo/1v25F8jH4IERqcL2pgacOFs7OontVO00M69SP0aywdlq9uI+mFOTPqWeY6sV
tmuN86Ryf5SyqtnagXAxmyCNFcVxJc80Jotf5XckrIhDXnpkYYb5OuVvzVlpD/iUKuCSIAiWLCV+
MOpFdEdrWvndaKY5mJT73AK8Bn7iqilGCNei9wveiB8PvbT5GYsG7uPzTA82N5DuHFjdYrUZpUL5
oAQQY08wwFOL/dtWuh9OH7/vhPyEjJ/1r7LzLxOKoJwg7akrFqyJdR3jUjlerxv9bgLjUMU/lJ1U
3kkw7e5tqsrGPwC9JrYqW706hOaMgOL16YH9BTLk6dRyqEwS+/E49IMxEcvHfwSA3dzgWcictiID
ffcNPqcqPLv8WIZuB/ukGYgLqzYudTAQl52LDTBXd+tLMPhCP3jOoTLDKTEb9RRfUwX4MYppRicF
WI8mrl+z97n+4mkU7D0Qgi3rsVu6USLE6zLuxRxrC7rX7AmuQLIMYUOWUE0PW16d6y16ZdDtjfK9
m5zVddgO8ag+tEvgU68hfTasaG4ebbx19PtiBJqKSZAOmIiKqGrNnPxJyrmAKdT2LrvO9pAQcDxf
0FXBoHVaBKQf3DyqZ+5NQEJ4NPD92jTX13S74drUqp3gT6skRzx/DEWz633JIrJA6AnhdGOoqJp3
XPgRO+xFkRUh1AjSUgybljoH0W1evEzwnC8SDzsukT8pjqpoGb//q4ii8KqzYdfTwNEGHbBuIbYg
GKfB6WhQVM6LMhAYweNvA/vtk1E/jkbXSsm2Z4rAvoYXbGBisuiPERlBEtRbXbzGYdYZtfRDI9jn
hCtlR0V2f4kDaP5cH9sn0fs4RpK5+weebXeRZYWB0DPyfTMXkKJloMgUL665WeDooNhrLY8HtiPC
oc3+PdYjHj3g5PO8aGcwLgJd1ctWmnndRY/SuURMSB5pW9jtSaN2p3RSW1kF7JRT8pc/Rt46ryCx
n6TYTl8PM07E3l5zUCMqCCrzypiWWZnykPilbVF+r6LhM+90xHNZHL6seSQRDKgvH/wcVhcbIef4
rrWHzmzS9cQXb7xKOAl+N4bxxcFpnpq0TBsoU+1RY08BLhu62wDKwxsvLRYBxWwFcNn4aqdAb9dI
9gsgDDuF8barlvGR2o9vdQp/4t3jOf54mAIgwYiJpJgheD0gvTPYYLreD0KbcYQ0Dp5umq6ricYi
z1Iil5pWkhFcUMfXb2Tx8lr92DK6UY3QnB+wXwGvwIJloSuRoIiDTj5Uiv39EwfV3uFg9+mYGHa6
cu+vzgjbrkKmrdC4+tFX9zQd5eTnsXz652ddbCYIOQ92LQsnVpvCoHArkYJNi7OTFNWFB5SSzKDm
XRs9lDfAHaoy9ZyA/QP5VuqvHjRE7T/Yd8+3s8W2KDkWmdwRMte13K9QaGMUeJiK/KTEB0oISzb8
rmXqCTbxXsQE7J0JphEaQXfg4NKM2JZdkVF/d5T6J9DLfRUeNRztL4icp6OZI59TvuknVXPgk46+
KFr/5jABtDF3XoQfbaJHHwzLRkItm54V4y0HpBWt9nmDO56WNkIJzhQDYarQd9Kq5ck0qFsg317M
TZhejgZxveEshei1ktu1uzoD+C5LV1YE3Bmx0uDZPnE05YLCgIPesBi6ibdCblzkyDHWvFlStD2W
Fnq8EVGSM3MZ0jbffnOjiNpQxNoTfFMg54uWAGyMt+XNkxmZfAe7C+V7OKFLkeA86WMqVW+TpOpM
Z05LcvnetQgkfK69BGJ5aCLFIhe/GkRFR3u5qMxcN1Bw7gvkQPZB/gF/IBAPqYmd/LXwpwu8zYpZ
gCrZBlfXuceHCy4hLw08UEGDLzvuzRSNGHrobr7+wldABreIFIhbJb5bwhOSeKP+Ivu2jW2y8+8H
SG162mkJq1yTMeKu+LlETS3caPSxPp0vc+zfS7wHlwXQW7di4882oQWdEk4Cag86THJfSzkyyB+4
v0T4GVEjR78OhNjA5J8XQq52WnGqJlXBjXrCqDvoTEBlScxrdKDDrgx+/ycDkEjdFj7Q/kgscpNk
wTzSiaIYYNepKy6aVYNPvClVkmdLM3UEf2/wU2JZyBXEMeuIVSR+KdC9J06iel/aYrD4odExvz0f
vx45WlrEWx8AZGm/ko1YZnpPCsOtWdjhCOYaZXBPBGICdkosoP3vzaERqieXBLj28+ry1K+mx2A4
UPOWt6WZ1tV9yJEBIC2MqXSklXjqFOylRWpOHf6IqR35M+Efbt64i2TNh24tbD7MONJxiXZJsa7A
nnDISFufeXVTHzhZp7hXZ45jdn+jvlDVN2EDmHwuOwHBJsncRZPzMPhea+swUUotaHM2GQ6BBtNX
aIQec8Eo1n02TM545hukoFMfhSVBBnqIzOiApiXxPT+RxuNDGkifIrjtiLf0fXUf8BTcZ+N2tO+C
vdAqEQpIwjgLJgqF1FOJBWxP1fvLyW+QB7LJlhjyxOvEu5wKtymtIdHscuxkfXiHqbxJ7LnfPALB
MB1T33EqYmgtKBTK+lqAdP28dsZC3G/ND2qJbVcbIpvGjnkvcfPVq2VSN9s1Wt3wrhb48/9w6M+M
UHfAPgsTS5uk3/T+CwtoN44zuSVeD+z4boxwiAS0k5hfR+cNH4byNNuUYFhbGN+K1jo0D5mb1ImT
vgZq0y4ZNeEkvTa7j/lVuG4EDz1A+3p9GnH+zVOYwxpd++ApdyipJCasP8OWANvmrbaVfeNaBgux
rQB5gu9RSBxPKRxTta/kr5xk7VujvmEnd2/5xjNOVVxxVsXjywcrISpOo/KoD60fwrh8CsFVFUja
bYSJTRDN92SJeZcwn571eE8Okb1EEhJccRcF0HXH4KV93opWio98k9EbAPj4WqDLo2TDdd61DhQw
QYQaEGvQsT7tk42U4trxOwuHuzhS/Oh2pfg1qAtXNj/5BudbPcu5JspJ9hSjy7oJ+Uty6wXa0EmP
5cSc9G6+6UhjbkbYNwo9nVz0weadI6Ce55/O0mFAY7TKR7KSuBLnn1ikt5Xujj/DzxkN48Xe5xRn
dc7n6G0L2GH4q+hExoP63ctf1C2WJg66QH0PewaFcVuF8q9gYSmgSIueNr+RK5qkMqLVtl98bScZ
w/NmGUk7wQV+PmyaXnMZauy/WQsZvTjMOSWXhEgfFxIcUdLX/OuExGMTThBXHn6UTmSNJklXuxco
8I9MRdrSYbcZT5EzWX9Kp8Yw62ffvJWVahvdYOE8kiF3lVHXuv5tVxsvIMCqIDftetZnm8byDG5L
SzK6TB/JA6RQjLs0LZIKr6yodNnLd6GpaQWxHxSeWdlvfhTprmr+Md59cczdvcwktNwVVlfAX3pv
Vmat9+Fdme7pUwc2pwEqOANe//4lG35hstiWsonpYeiiNAeg5Hy999ciqrWzvcgT8/HnutFLklyB
5SMcgr0yezVMEBAXjSqaGMcq1wZU4357RtNM7bpGioKnKa89nzB4Wiro2uaKZtvTEDZzLqRw6h2U
u/OG/cLfZeWFzpr9rCwzwg3fEBwwHiL1DZj7wFy8Wb43UQQknjAAKvTtP8aVPKV1h0s+NWXvkJPa
gGyNhJ4Jhxit6+aFREyHtoQEmDvYkL0bSSw+K2ZD8OnmtgAETu+Po3ZwTHSMbJcAWqLd3rLYQjMS
cJiIYhbb19LBCMY6UTknCzV6kAg/PtVxkbDbPqkQwTAoLo17+u2cbjZa7NZ3hl+lc8AtEGczx1hI
gdZtm5NRxDome35EO5LnPNIppQfFMfMYfIRK8juo6kkeCOA4KMzMDe6xjNwWpTnMVAwJl8tCxnqv
nUuO23J/+ZKzTfEgYLcDAeKp7D2ZsWcAjJvQkoT3yuFZLqxrdj+s0Wi//Q3BgcJvpz4Lx6rqKXBK
rGbFzGe/HgzmEC+Efb721+OfGBc8rpGujC1LVEOQKuObflN9QWKlSm2eE2326yx1oFKqYKQI9kEu
qSCELv6YrFVvKE4dOoy+bDYEWBBCwZVdOEj+1eaRb6N/f3ypQV8PD5Irq3XuLQfE+Wj7SeSkU5CY
jhrSTE7k+qB2ICkD7t2zyLbLcdAUXKeisbAmTHWDcYg9Zjb1hjg0PstlrUO5emK3p3dP/hFxplRe
NN97ISTQM2yh5OTvkagAQRUlUQCUk7npmLZSaKXV49LFSIRqQWaEtymc5j38IkfhN91/HIyFGYhx
qxkiZSDdZ3c2FCLLcGD4ABZ+oojHMNhiyArvpYbUNIwMT1sorZxfUfFw5Nll1+fZYIjoJ0+l8uqI
EvScdpbGl8iDlhd/PuhSiO//1osXggB3A3p8KiG55MNsIdo1p9RSuICqe2SDIk3cEGsh4UvxDmUA
ggdG4+y3b0NOLkKx08JMiFZ0zDeOkMxJb9bnNjfhxfMxZ02BSgJkV2mujHspcx6mcQioIlPp0sas
v4NJTJPo9CJKGYjB6PmJ6yvviqqXcDD4awipR/n5gxUgyh5BIl/Xj0f1RQNHWdUJAyJNGPr7NxCE
QAvfGzZzWOtAK4FkwopUMiQu5Y5t6LaiZ/LOXIo0oorBMC7VR3L4qgJ3dqA2ThgZdkTA4UkgBvKn
XRLcKOY2W2Kr182851JNach3SVnG3DEgPQaLL4Kg8VTUCPtM14BOu0ecp3Bz3v94Hl3RjecuBQva
coFkmnqRkyP4iOTjtpq+tQOhJ3ox/rECAiii4d3V5xaRNfYbPW6nuCG9qPiIq571SLtT7EU6wfgY
WAy0MxZAsU1Qq29BdZSA2vDz3SD1DUoNGppKjjqPC1mFvJiRMHL+wliAJtMpL8GmlDIoFH661WKX
+iZPiSYEkV+ZZ60SXvU4eFDMdpcX8rf3yl9xP/+ojp3EdTNLBF5d+MKYznpIkxQ5XlQP6IRtkDXq
xuoKx4RBNXzO1IeZORq17lHV4wGkn07xhbxCbiNXALIg/EOAoFyiaTtstuTrsdH/db1nmQf6UrE5
rNx53+wKSvEXMZ6lru51xKrla/lE9nO9YYIaBA9rJsrkBrQjLgstAtHDYpjo7QWdmNxy4UH3nbaR
DD7gHMn7i/YbGnbxjUjcUiIi/0ZesZoUoZdPBToARp0eVSYrDO0vZptwsowBaCwDI1uklI/vnJL+
yirQn6KsZd/psJ+oaXtHGyUrK/s6AeADLcMH98earDmaRc//bzYlM4T/BQAruJZVjFyMMEiV/FJU
fhEUKGPEAdD3qrTKPDk2hR2W0iiF6JnFNh8T9wR4i7ky+I0Izhr7LWEMFmVwwFv+0ljYdZApSGSd
5I3rteRWRUsC9qgQqcwzWv7X9Aim4uM7jJsVeyvs53oceUF82Z6Mh0v2QCofDzkvv0A7q22zoLLE
15QO3ixc7syJTOA8rKyhbpzCiAhGV4OzAyV1lnMCBKmS1rpTRPEIHzEKKKt/ZPYOEEdbThM6w4Ui
+9eiwsXF0iE3OC46S85Z6byWftofpGPj0D+9Ode20DFJnvngoofCCamsH6YO+H5QZFIszVhYc99d
5yoEyXVOuJMzhVomryad0MilpiDcu/hB0QgxTJYvzVFNNyuTe/uDtGNNC7DfXdwwtBIQbTVzuZHu
kRnvzIgrxqNWx9/F6EgXkPVqWRaGmFLup32G8jC9gJTeRjEtijz94AnVsruLZ7qst5gnhnGZM+ld
+9Vj4uucwi/MmNNr9YwyS1Tni0Zr0+1Q+BS7iIz+zZAjLKWQDCXEbKgnIPC73+N71wmmrhtpOIhq
quQFL61x3BZVPPi4HY44aKYXTNXnC2quBqhakRd3qTNdgpVJPAZqpZj8DChP/410AnbglIl73ClG
lcaOY5jjAXx3kbU6Y7gXRrDf8dLQ/ZMN7owOflsCYDvvNf02znXMwF3ig8hS6pq+ZIlvqNY+42cE
gbk3jHtI8UHo72W6dLfwUofsZkEnZRFy9fbH40ia8xFIvydTRpZnJK4a6WMjYbQFu6OZWCFzz4r+
IQfYgIjfIt5IHMFfP/5gAX2RWCfTOcd+9SS4hWYWlbbBqV5epCJYHAdm6Pi1JP2pq3jiaYIpNA3w
K9AoCuYqrIESWtXyNo82RQLp15t6PQBG8YQxAg3V1B2ul0pT7eRTycBIrltM7msfLLU5jtnf53/3
fPFGccFlJKSL5NyDL7Giuk0EJkzOykT86ElgaWJSRPkRsH6pmeYSH8jg4Z8WjjT5rnxRNmfyY1Ag
N6YOS2YCJv93Ru/DVKSZqOi+MJdIMpjxU7NWyiO4n1QpPcJ4/uyp/4dgfT17w6jXOS4lZMtUjqM9
n4nFEVNK/CKp5PhInfqtQIr7ppxi3V4eQ5IgD9Bmi7068q3dN0r1nDTQi7qnussgHBHBMTJ6UeSm
VCFIz435RXpNbKi/XPtdKXWXflv/Cig4F2s47GLYiOaAo0lmcsM3dbWXG/rCo9anjyeIDDLCRiZf
vX0su2pII/5sLassCFzm1esPE1+MElCl0Z54iAQU9+2787PKbcPId3n7anjfHs0tSK4l3KlN7jUb
SeyKzAbW31YxDU/At7OjpI7nT58e7/C9gFu8QWFjjK3bw58By9OxeBcLpjl9kuxfKwbn/LVH6+uT
g1yXJ9pmZ2j8S6HueSmW0bcgJSr1dZdJGNyjYr+wPUAF/AD9EjGBwW8mY2nngJxQ1AhyG4u7djc0
5BmOSO47JDPiHUYnYM/0yOeL5FcIqPeOxVuSWimRPi/mnv3LwaoV+uWvPCTqJqONl5ihmFvTFokO
GXS3AaPQbZSpKF4VQLvXGTFqJIpYmGH2rT5yFScLXGW/hyIZ2k4ylXHNYVucAsTL9E5K484nHYkw
6XASr3y8rRrKab7Thjp5Ao8ztlDs5SLTP10hGMJvcYWbTJWnileGhuXdBR2L4L0XPW5Hpbl3XtVd
9ns7KKEp2TQXlJmyh7PvwefhN5kp2xEyHTh02Q2e3htamIxegqPkqhtrC4Xdv4bL0yGJEH+bBy01
RyVF05vUCIIFwBMYuPHuv4kdsBBi6DDjPSXVPERYHwIAtKUx9yJS0QRTwW9fIAR2FT0eBeCbQg4c
DLbt5Iw5MzJrzky+OxSuYBhe3K86sXoOQwdHzYjmryaTkoUTP7bSSWLlqVzj1wlz0uE5aux4uKC7
mYFLPEE+15XSaDDiOh8p36Yfqr3yFxdwZt0cgYYn15gIf6wE4VF3ABb/Vbp/H9Tf5YUp+jiGqtHC
X+WkwM1eGPTm15BfLU/2i6K9EePmuPAfxpSOd76QzzenGnnQgq5B37U5y2jP51mCIa+8SzHsprm5
A7/HyofE8hvKNIoR6vFOjycInNCDuIaN3kIjOAcWstaFspxjU2mOeDDc+FbLiKKCuXBsMij5PiKQ
7z6dzMAknTBoxmqQygoBOUO+kcxA2u7/CscAnWQD6gk54nlsWcUJ+9UkQvuc8lKhYvUv4kyw5kq0
U4Y+ooqMMkD0dvbxt97Rolvyg9tGPxaEi34pduxI5QtflRpNK+5oVf3XNUZtq4rcMZFVajgL0dLN
p7aoVxCySPwVOUbMRnhwdHO6CIKf6yaCxuXoLfuF2YIAvia8uKoRsvvzFbHEGbsosTEupkg2leEL
CcG4COHUd/3J5TQizWV4PINobaXw4Uaui7SEEUlIrSt2LDSbjDOzvWXVdNiTnYF/+MVmlhzmglbv
QpE3VG69NjsBtDRCp0VhSm9RyExiP+T9XjU5Ot118Flc987LTARt1E8QU8R+yvbaTYJtfg8zMeIT
vn6mSpJKw6i21Q8Yz//Z20PEVjHe7HPv3sYxAh4Et/E0YaH5O1H3NHduqIZuYf0JKGZRhY4Uv+Ss
EPs/jhBRdnMc4PLhY6os1kgISbhLj/p9XQXFi4tOVvenwIarcUFBGKKWcrqFit+ZoSbB3XbCaShh
/4FMrfT0IEBWITkRHAQKDtDRVc86Y+7A5VHXhtHhPzY/RFfcAK2mI91bIU9BqRl7pDFYCvM7Ntwf
gtztAaEsRU3US8vyK/xkqtYfnViiEI+7zE/H14fUWYde0hO9qmedseyjV5bR5BgKGvOkb9jRMV6X
S4Z7LR2/TlDqy8agDp8O46l7FcqrWmkFwrjFwTolXz0llAvJN0D6Qjf9I8ojFV0ifFFuTNLsXA20
ZuzWhmdMtice4rHk1Rdpj9fZ+43MhQ7O7RxUTLBVY0hj4EPefMH2zRJ5WRyP6rGRK7ds44amnpZ/
1JgDjLMOAXwYJ5Uu16Df0hfTxlZBINiOvmsemK95O9zQ551kjDebwleBwH+5ZfSLZaJMXsbACyHL
YXCIXZTuaRIvFtAhfP7kHyPsosE/IGPcCW4cF/l8NRPBLLrpQMa//E23bYAeO6/Dc0NRo3yyqLlv
dJttVCUy2Jc6vW0Fs2rWRKNBNKhRqxrHE+jwWYbzg/2tFajhOVtQ71tU4jpUEnwL92mVrHVfhaIh
qoqP17dNcXUmWX4llfe+fPHon8O12PmSrhzWy2VBZ5B7506Xs3n6q8Akt7rw5ImpeUK940bCtpqO
msDFRM/734BU6s8HxxAGq0NFcQqUJnf6mPPnCA/B5DlxNKtK+J3MxItgUvUunEmOHHUu0AFjTxTA
AIBO4MkrQSYhAENMT3aj9uHsY212Yoc91y7Pu5pzqOkSQWUoqseOzGndp8po6xKvf/pNHrgMB2sn
5tSZqPip/VCzDS400rC4oJw78YjLdKxto4Jt9ZGJRph8V4Y5c+lqt/+kO420su4qowKbi0LWeJGQ
VpEC7MdItAHkbLeO5+lMQeJpDbE8p0iRyLxY5KnQqB3JHqI63J6yTyG6ijoqjW/skg+3YXPp1z5L
hwH9Ud8/OLGTMNQb43FDvLGti9Cq6HCmJ38cY/2v6NW1SXaRKO917ixZ7WGYtz7Z/YViN5n3voJ3
znZB9BIPqUEDSi/9WomMFalYq5c+8rWXIYPHEIqrAF3hihO6G+8QKZXisTYh2Uk8wqt5Ccf618kq
CATxpMXGqt5mODGp8rdiMG8xwVfNjc2bXF9RnPPELxSrq2tN9fSdoK7KiGKoLdKXyhJj7iyYvVjZ
RNFADpzJVJf05HWv5sPQyyW+XrmDF33BHqOf8QEtLz3qDgpdQRsXziqn1yOqY2fcQG8n0o+hle3w
NXKJyLSTHO3aDcwmk/l7XtFnG7+UIPupmISBCsXOwT3yVLxnraGTiWZCgbIbtqSrfS18NVEx6w62
9B/NfomPJXt1PTGPNE+x3ML295SGnL2If1Vs9ODFDSP/4n5ut3q/jfD1WY5zMms1hMLCLAjDkd23
yL3tnvSm+ng6cYavtfdHmRR15fxFql8fTw2qoQrEYFcBnR8Ns84nAlcvajEAqTpGldG+93TKFW/Z
p/6SkNm1wqSJo/zrh5Wr0sR/wj9+RZlL8YbOUF1tQVJp+UJJmOIHTRQbD9EaapoqGRvRJx4n7NW3
OSzSEWIfCXR8dJBdjgoKf6Qt5oZYxZ9wNsT6WmWa92nhlCvmgKL9737jn0lmgGQi39OH9X0l7mKe
6XxCFgn4B6367GwFhJChWHGmpX913dEiw7OPmeT7z2iNoG1Ws1oqvC51MHZeBOuJjTIG0N0jm51o
YLWgalw5SB4NAlzVEyJ9Ypm46fByPVAvhLpFiVk9g768aAIivNkkrViRFAAJkES9McRr3Vy/KW/h
3CVe55URMG5I86D4mjlRf8xoiHN8PxyWMvsAVfTtBfIct1DecjTxJ+Hp/AZJAVIr/YWaDxjbRuqh
7SDk6rU8hXUm66ujpqWjoorlWslaRg+ohS8+kPkFijpM0LWFKCLf69MgX4fK49kBL3Znclag927y
lBqWbiJt+Y0BlOsI1m25vmj5oi+i3rif86tjxHF9R7CFIl2b9Qi6WJer2rxX02XDUnqth7O4nwR/
0Y4HOrUR8RtoHsqEA9/P85TTzD/sv0HmR40c/4IYTxCwJiLvwF6vfPxKyDeeFxYaPsh7d8gG7xzf
FT4l6Dgab4dhPJeeWLfS64ePgtLAwGLzOxIEZfwJZxx8HMncw9kY0UzX3sQ1CkQJyIR/yvgzFM1k
OkkU1OYSoxwVxjiPHyGzFVFdLrsLRzGjF73Wb5k0SUJJKfNvBNhjZ0jEPK6cvSrSJY77DBSA65ME
yzDPvWqHNYC7LSSsnmu7/m3WrqBhY8fU2GCLtHg3k6RmZMi4rGhe9fgFI3YiXtroobbcq2pkFLME
dJfgGNw9tuUkE0XGccm8mstEn5NDWoS13dUQ+7+DBZXDQMPlmtOZ6HSPzjrWmJ1foVTunWcpuydl
nfao9QkyFtUfkZxlxwsws2bepmpAiQnIozkoZTTc8XHJdJho0Qhrjk+wYV4pqJn0A+6RfXLpyvIW
KeBku+1x6BoZSffaywaKcf64lWg0NTDewIQLJd442hBBPPvuzzXKzYKP4aSxYgMUXaX8T4nA+DVd
WBOqE1br80YAAW2PsIqXnsilSqY68vZuNP9OcRZuMBKC/SCHWI1xDj4csjSlCBqsPMHi2KM/w89D
vOm59EOw8Qp7bik6IDfPmG1FlwOakGWfeorTP5cD22wDh0rlzB2YD0IUSB0jlc4WuCjabAatpexU
PGwGDyVnmFGOEbBHX61wj/XtKlUuDdCogmuk/JefC7NfGBYdVRdVCLUjng+ugLMHCEdCqmrjG8w9
tfAwpyyEc2LZslvBoZJWIIBokzJ4IW3OlkrUT91sA1te6cdjJMkTycuLAlaXJYHPkoO0NqpV+k77
nKB7EAJ6MGoQIWJwCKn65LFSuCqPaWvDYCyJWq7go2f2xfMcI5NzcPPUt5Ll87g7qLe5zx9obbry
GjH+PNbzIuqvPO+4eu2HeajS9lTIifqGRo3y/EB6HImidd8vlyV/S5k1g4tGIU3LCwqgg6vntG//
CCnaq0sdLqgXqttU3vwDjH0madVFpVg6JAbcQ6+pC1DM2C/OqsnNeoDoOON+hLt5VLa1G13TIiLu
sVo8QelPobHxVIS62mfVOYWKCTp3T7q5F0tpJNhql5AykBP9ChE7p1yHzhv8wQojDxziP9Pf0ctL
FfGIhrphKczNciq4sdPmjhxIk46gI3zBgpaqMXSMXmbdTbAoVcGdUHpbZXZvjPTOmGw0wkhU8Cd3
sId0xBMswMXDroc/mBQhwrZpOROSZ/2vx5UTdJS/JmubTbYAV2kDUdPI4+nNdz3ZXteqiHkxre7k
uipeGYeNTP3ZJPS77mhzZCvBED9JeyLg68v9BIumkHZRdsdnaoE8V45pUjSQ6cGZcshTYTJad3gP
bMx80srP3IGVqKGKwlYXRZEbiM1grKKBJw85SX6IDYoecGLd6MDlB3lry+Fb7BgDtPso10lEJ6Vl
ZhJXZ0YhDdfSP3/ZTWBl7YEfZQzKLHZ+PL1P8CmSIbzeUlf/pM+32JThbCj9xowulrypX6nXEvy0
UxVx21/Q7m7L7I+tKRxJjtFtkHT1aJIard3IAGnVKAT05G9EibrhMYimjsrI7WontNHH2rywIUTP
NhHriDCL6kR+m3wOUAJ/xQgbAxy26x/IzN2gr7uGQCfLFDdhBZ1Ycev4YRWBdXpkhg9pcZBwabZT
j7MTAAVjFX9gAY2pPodFn0RaIgUWy8nA2xcQqkvve//heM9JhF7z0vXs6DgmuqX0iw95ATxoOaMK
dMZU+SnxbvoBsAiwn4QX4QLsGpdiGe0+mbqkFh5CziYpLnSsg/hD4A3FoRQKDGPwVqabTclXWh7q
bPP4yxukO3tnAEm+QGAEFkVPxXm4hCLQWOabqsDIfdKRch1go0XCanWjRkk3KHpNN8QjA94TLqTn
e4SaufJ+HxOSkFpyfnWanrFE4XfwKag/UUuYZWDWSld3nmUAzXkZuT5NQXygaHjGs6xNHXdQbWQw
Iw0ZulE9exh4ehPQIogwWd10xRmfQWkjwsoVae/tp2626r7h6Gy7R2kn5uyylETLmk9eZsqa0Xvl
iVoJ7cBCq4ni+/lrE90i2qBzMpHH/xmb0eC7lz6RtoB+hRS0gVfOeETSVfmrvIqonIIlxzPCcJnl
5Z9afhJkrsvfnIZGh5lJYpfEUe/KBawZqYAJJGxKnLrCGi5Ze+9kimDqCB5QRQLavo3XHy2A09gL
ERFqo+sNkdERDktOTKjuFlNUwZ5le6jZZsMBUHiCBZZdTNQk0XHDmWmTVrQqnOwhGsw5ZJsIF+zL
0/dtbWkjNK6QPPFGC7rjm0iLkh8rc4somKmLcRbJhm0BaHHnh+oa2UcPgsjWIuIpH4lOo8jNDMSZ
lN/Z+H1NCz2UFpWSsT5qG/NXhDxSBELs/hVVEV6AhX/XvHbV/s8WvUYXbtPeuKkyN6dJ744GynOM
ipYTSl/8GgzJ42Xb0u9Blq7Rj39YoKoqsCcv17VGExln8qFKIdkU9MajopTHFxS1OjjUt0DkuTzX
xzshikw04dYyPdpnwPzCquuCVvLWM0/6DzHlNBayEL4KDfD3ALqlGR2nSKaxgyocRogkW48rJIKm
OxDkTflGj/B88fhat3w+KOTMJHP4IZhw58H2P/5cix6z6l7a/7uWWuoOnmOcSoftLCjVb7DHbjjC
fXj3FLvSwHtEr3zZJRJg4HE5RK5sfCd94vy86md/hDnmVUXITNXUwyUr44IbItSgZQF1xc62An+b
FPqcd2M8kHI9z2VKpc+CfOquMNCzYzx7e1CqDduFinhIGNLJol4pTdX48ZUya8DD6I8hdkQ2I1f3
Lr+TBnAtS75ltpodOjEFXvfoRyPCG8ZtfEva/FWatNSzYS2og9ZiXU1Niy0zdWABgcCmNwNCEGrZ
byR6FeKLXaV0hkzhICax/odcRqWXVU+Z93WCCZt300rUIO+5y4GEe+10PXdNG7CuuvA9fFUiN8YU
0VXs7/T+NqvMtPiYCcbiUYdJ1D80LHexhR37zhCStiI33uZR7Ce22XsCzaOkrsoeIXgzH+YRzdWd
SIOw2xkkFa+MTeRHqbfuoeqBKgGzcP4kKvU+9XnpVHBrOFRsRwJhN7VAsnFXpWP+XRrAgxpEpApy
pd/L3HEj3/x3se3wmrGCgSBDEd6m6+WitZVX0dGwzjfOzA4lzNAybNzjYedSw4d2LfPudSNdVVI9
lvy4UGBA6Th3rZ8dDmwaVDDK5GlI6L1DUjwFLcA2pGAkrvjnrZs1yM/IjVXDH63HLHUgo+jy14In
CgooVwyDPK+9OaMHr4eopTX8L9cyN1zl+EYhnTamq6v2fji+v96seTeuFDobi+A+7tZw0QHYHjfI
Zn59HBIfZYwAe5qFr2X5evYK/h3SvSBHiTStHBpdcFB02pXooZkMQd0/dqIYLkdZOW6lQzXcFurR
2eIQVobFPatxX+vDKnB3Vmcb7LZmGrO1Lx4MmNrI6eb9gWUU4DEbG0bDSrR1+XBeWvXtgfz2je0+
crjrj1T+cMqZexHN+UbjvJGI7kepYUJCg16TZRp2XRY1g3yhFED26MLci4E/9kg7Pq5T3fY32zMt
8UlS3+k0nx0XlrMYxQvLPuTQIqeDN0e8eyYxguPGfRP7bjTOr37bQAD+wXJBWEUQxKgTBEyEerQi
wW7dokCUcP+kJ/z3vXiVq5BTHtWMOsLhe2gafIolBeA028kGtp7urims0HwB8Gc/8n6BvAXpvXvh
zUbS3g+bFWZmHZeN3cZYQw59yUUdgSYEKyDLCif9TmsgPiCACIl/9Wzde0nhGG7wdcxNJusEjCFp
Qyp4AI63t3eLXnIURV0rAU93zZqflIRbf5D9sgSPF2zLj2xSr1xtt4dnpclvzr9fe6v6fnrCmAe/
Q6dmfJOgIdebPdSRfTqZCcCgxkW+AlyBWoi+ld6zXtCd5fo3YUa0mdRGDNwC2oAIH56TgTaDDvH9
A4R7aJ1k1wakkC4CVN7UtRq6au29LQwzAT/R56zq3PYxQ0afOz+HaNkZToH6NV8IGlPIof8W88J8
4C75EkEkgm60uLX+Fmyyjq+4WlPMWMit5v4l8n/WAXYmZXMvjQTTcD9GMTKryCpVnhdSsVv/3NxI
FjifQiY3WOh+V3ppsoCs1Zv4Fz0XYAbUpCUtLFLBR2YB0vtkEL3Psnc+MlYiVK7+v6Fghs7X7+gm
o8fyOE9cvswoIacuMmQIkFm6MT4qJDBLvtWzfFCcr8Vx6tjsBE5F1c6/Vw0MHRKcPv3yMEdJvsK1
Q3HfGD7B2PPHSr6prLJSPMFkOsXvz0p9fnbibLdgPOjEXKJSkgJnqwHHnnsYgnvy0sRv3/NtSdHJ
AvVzm+GGG48L6boGjcSGGpiw4NKJvFckzFs6JjfqZs5/a6NyRrDAiQYh390RKkoDrcHcFVmGlpIJ
oCgq0vpu2JikJIrr4gqnF8iLbpNgKg8mWyeyvr3eVidzz7ZPSQTthT5RrsBMHmBVt7jIiCIl1G9A
RnsRRInUJUkA1cn9ewizciGb0Xd2v7ZK2Zkb0OCHpZC0EkpKkwwruAJkHh/d1z0m8mb1ZyqtPcBq
BCC1SHLiZStdsGgIz81/7yefdQ27ezWPoCoNOiYBFL43SKsM3DzBNjHIcazOqRvwE6DHqm37levV
MmsxxM7ZeV1lXpB0W8jD2K0cRWpmkOk0EXkYiid/2WuUM9Zr9GIXtxdwlYt5/4ByTO9id9CtibyC
E0ibi2J74Rd9wa2RE0JD8Sg9gynDlWdsIq6L4rQM+WDwfUGhiPGT/7JYbzc6+SzVz1xdFwfkHZoa
TDTVF4WqlIYNuQSPNrLlM1OaI/Y44lzSd/hhSqoYopqMWKWAIYgv8nZfcBBx3PQckLN0knUmfhLS
ShxRi7T9GRsRqXWxZVeXJuTHh6is9iWvZILU2lSYVlSiWkAUe0eVOxUjZydzMwNDUQjtFzHyw7B3
Y2L8+Tb0r2+hZ/gbuxYsCcXeQO1HAu+AoXgVhECkJsd+UYb6oHyCrsRxdZb/Z93qRDghsgBpu4as
Xpqj8xpTGrCoT9MVVk29B1GtotIJP2gE5D5v98BSD3k7gCDi1o0XFrfwXcCaPke8xcj4SY3qvKrA
2Uvs7hljOr45mPAKnjJu9cayjlvsr/GmonZLkh9gxiF6eZ1/nHbNY6Wjb1+x2PYwoEPimizdsaVc
p0Nvo8iKggts27ttXWwYSyb/DfxOJhWrQ8KdceiBbsJqDNlcVfQGMdA7wZi82GkpRzPruIDjZ7hB
nAvJ46pVG7UxakDF+jFn1+9ftR46ILP/zlGatRNSR1drbNG3Y7VZNNNEwHM51Q70V6tFgzpS5DhE
ts7DKO+X4n/qU1cBncCAoFrPcI/Cu/4ee2Fvr2dB5wAUVfvlLihdaw/h6pbZA7FnWN7nlS3Z4tn/
6mn4UZnHZkHfJIwVdWBWXWNhgy9M7t7MToOhzdyxVTdsdHd4L3tFpNMjnvHtztNqc7dBKUk6iscF
wvT0QwP2MmO7C0agM5FgmSQ2zriFwTo/sR/jZJUHhsYdCVH4wE0wRD84aEPkNLonk+AeRXtIAZtX
//Gu9Mv69JFwwiGgMa6anD98lxWY6z+9Ef8oI1d0Tt7TdVpaQQQ15i5AGDnzF/8b51//NbMm4UB8
3mq58QVaJYZ6M22NOnVmJDJ7gEezc3q+hW3y6wEUTMBWFyXYmQ5Nyoy0NpAEU0d+uoHL7VWj+thg
X/dHdfKJHzlANItULKbrrs3GRW2dGxVphWgLD6QHbMDd6xPOaxA5PubPDxfbSiLQzY/Mf7VoKLVo
O0JfcRI450A9HuzXeedP4L4fnRv1hTmt73c1dkQObRCg/p1/+cRAxlSJn4kpXBrWGCcfHHxZC2a4
Muk3rxMOe0rWpajPbVZJZtquJAE1xkaYpjFpZhZorw338IdY3hO3aqPVQy+eDpM8ksSmRqJc5m4/
rLqoSxV1BymwhIYY7oNrHghTdQxupopoxU/YbPZXmpzaXWP4hK0CU+q0MKJ0zlE0le9EDzzTh208
36wor2dejxueupMWwiJcspI64y+1bI8j7cLaabxbcTdd29cBW2fQx2vFio9jQZIh/zRBoh20meqR
60fGR3qxSpwrTzaUV3MdqEXvZTS/6NaNXyco+/BF1YK+YsUqqvOpBNVEGWMiIDT2RgqUTEZ1Sgty
uGZKgcnq9GIBSFn9V6wTHSZKqScwM52JoinfLAB+eYQqTS/ix/fk/AYTga+uRsGMZMBPg0d7CRIc
VCFN2Ag+zzd85PVk46LlSFQZnCwjWtTDygwanBHOhGqlKwKaIJuqnm3q1bYsu1HVZuhOaYp63eEO
z8+Yp0gVUzX0jwbSaW6lO8M9XJZBaK6DT1dBX1a1rIOzTP79L4m7BntfzPSBh9mxgZ7Y1DoqNEWv
1UBtiomxh41KTarAscEY66iVEk6xVRaY6pYwH61KNg+7F3HRLzKSe6uKezw+cSc4NUCumveNEmSw
l18Isr1xVex5BPjN6J2XzuU1acmzQ4/AScd9/4TVUHPqxcqOTxTJ57fGB3xvNl67IOYip9XPxrGL
XTUBAIsnDuohYX1TeFHO3i7zel9TbIwENEW99+aWhqar79bx4SWTIsQEkUbcrG5rigkB/GTiMTK+
jCrJYa5zneXCU1mwKbcYuylqz6GzzZ1XlvdCycN5hDo0A/7KhjHc9Fi+G0bXU4X5KT0sM5bJBECe
C9LBuyVIyk88IzxaBWIr8Q1NXf0IrS/xk72VdzDiqRs7wibUJCziT3koqvp/mEujdvykiFeZXPXB
EgC6oSp/6ZZAVP6/rUUa0EgTi8A/HiVwxR+/f9OHM2aBMV/Fuc+c1Rei/rnrnlHoRunbEANXwGy7
4mxDvi75h1t0Iz20mhVtk/mbMjZ5a1MLaqNtWmCqohyiYKoQLPlS+pbFJFCi1IEUdQaEBJhj9pz1
9VHcGeDxyBcoDo2qkZARzAdGrE6XIzcYLH3BlL2aZLa6WU8Eo1M16doRf66D/UOtX1Oj3vMh+Efl
gqrg+z193DCWeJzltjz1Izfo9nqah3qNw9oFdI6hsGhz1yrxivvXrGT3Xd4c+3ZE5rFBDMa/c22V
op8ObiJyj66QdYpEHiq3wvTGkUTDgAa3pGSIbj0dM/nJVlwnQOfaPzfXuvf8XlejPhCqXx9G0np4
t+3SjK20x0jesoukJMPutb1GpPXLpEVL2C/tMHmYST7C1Wje07t7+t5yinGnMN5yspKJzxNLRt4a
X2e7rYyJ963ge9m40uSR9C8+x5TiSTFrxnv9BUc4gcOlFGk++SvZmb3xF6omweEhCASW7/9/z60I
lap8fLBwdhhX/er0J3cgtGv0oiqOlDOkU4203Vlo7Mq1U2iV0Tx+wKzLhAKLqqIimf0L1yTYJBGF
nXtHbeGr9DNmsI+LE4JoI53ZTBs9B2omEpAF3EoC/pTaDnpqJFElFYt5cMdVkMblXE629yq+No4A
hK8P3oqVuAXR9Ah5M5ZRm5+16AVcLeY8IZSUXOV1msn2puaT3XYH0014wBHO8c0rywZ0EuBemdeP
HIyv0nqbhHD3R26hS7rxdiWXfLXOF2x8LYtTwbulQk29Ctwtd/6QeAesHW0TjTJjgOosbajW0129
knQmYSeb3BB2PxosjiACPJswmaDAbaCaCmotoxuP3vEHS3PxDkDPJPWt/cLHCtxBYyZSZX6h/I4E
FJfYbFIZK9qiCzjtgfKk9pHqnDoW84iaV3oj6MCqN1QqGMcLjw2pO3n4SKLuh2fFx1rzn1SqxyOD
LAnOU2cfFUCxRjBf664wp3vS4ChfFSD7andZqHPCr9u51p0DhlnQyAMlr1QQprTNwY2+lCGZmiaV
eoQLgXQw+j/UR2oMDUstA/9Gcnhp6tP7Vnboi6I5/x6dsl7z5GPEZ0HHVnHt8jCookBWrij9uAZ/
ghR9mc04hc62COoEmO4scoVKLXhRGpqazc1qvtPU/pLVTIjRZ0/4jcMtDQpFjuhdxRcCLqEB6tM4
kyGxxKlDD9RqmYRNGAeE81jZ6PnBTqhZo+4m9/bmiSNVXLJmx3ZUz0ndCKoz0oQj47XK2NrLDnlB
0EVF90np2AVELQdw0F3aAynUi9c/KYckKrcaKfo1MaEvv0IXqpHJfsXI4o+sz3ShVtZzOFDsqv9y
vD5vAtgWytzfERLKd0d1jj3wpoqY8ZOqE2SQw5Zs94JrZ24xA8KnZSGxRNZLq8JqUk7yaFO0/ESl
yNn9DDlZmicjmKCgc2n/zgB5vzasntp9QNfGOoV4K2UWa8IbaAfHrUvf/ZFyDlp3eY+T+r+8dPiz
LfQGNfw68ckBP6teZJyFY+XL6Jt4aYYTSzdNw6XruxKlb4i4VO8kjjlaGjYdl7D8oZKQU3w7Axov
KMCJz4mBnjqmeQEGwTbjWx+Z3Z21+2BcLgYMac84/uZ0TajPCY/1oep12ZQMfkCHjyerYdtdk61G
xjdojpXYMY5XKPwfoTnasZY9zXzmneEnErRSvsyepEK7IT469qqxFlp7C1FilQTBW/tUv0VibCD0
vLn6SmFXBGXPV3RK7B87rRWTDv2v+py1h1afh4MMno22+DLX2w+MWSmNwmohzsFLBWMni8ALvn/K
38yWb2o2yFVpVK3HVHqi+nkyqTPFA7uFyjt97MpkdHG8KbZBUOMRcDfZ2ZNzvcijv85hA1FrPTLz
wtVIlf7tXObFbhe1AgJSnh4KAS9ucARcB/CPpMUIW63gImLI8gSJzegRIJjxcecb55xjjHuvS0eE
59Q3EG7NkIb97B1zmmFoA1uIp+w7RDLQNBWseSwnF7QmYXfFm9eAizjFCAPAfsvxOuXjAvbFL/aq
hYCvLl1CdUUkgPQnqsoPhC73mQBErGxzyYguIpicOKl7EPMxpjPqpeY9HtsVJH8HoWOON5/Db/j/
hbBV3Ud7Almrjyvz27tIK+m9nCQ8QffO3LxxDryhCvZVKVUVIXkcLj+NdZSYBhx47aSAS9FgDv9m
6DKDjrwKp9vqjTG4XiA+sYpvY8tfEFKuEsS8Q7UeeDranY5kjlyfgS5sPwqquC3U0CZn5I076B1m
i8usWZCROa5XK5jznzTVPpzvRZBO3wJ4LoSESyH4abWChTyrCPs+Ev+cFma3vn2WPQ/T/7LoQZ72
Mt+iMjImh1BXY9yPpS+z+jY4jAOyvvmmOxK9fpWCq1YWpwwNE5k/6ls7dzbEEJQR/GJZUvVYXTt2
WiJpU4Xq3rsZrQbSTtBdF9cgYENcZbJYXhw7MR6iw0sG890Hv5CijUle9qWBimXjnR67zK+NJQIv
DaJHGnOkucqWFOpJFFFfcN8dPrxWynEUhWkG1Fa0HjHZbljfPHa56pHjWekGcVp8BSgzohSqZge+
5suN9jTU1LJHpXtH7rtqa6doZg09PEyLcLxIQARBH71Zv30RGAdHM4nFfRHrn3uZD5f80DFDYeAa
v+ixA8wGNIuQc0m4iJbsbfnrvDLg2y6fU5AL5EPXYbOhc1yg2X9tsmSevClHogC0L+wiCDBd7XUl
nF+uOSKEEl+yoiDExCNxptCBxIU8UVCi2bZ/v6HN2YWGyBtlsnEaFdQFv0fdRYfKU+urVejhrf8O
WKkVt8dedEPVb0XiXnnz6uXk6ZJ0rzyoa7i9Z3zBeg3kOp4+R4O82vZ99h5ig+X/MyrXOqad9xpD
1pu7hGHRFzTTd7Zv78GROw7/667I0xPFDVxg6Xb5I4ezrTktIg07wcCYK27R0/jHUyxRuUXFJ5ph
ksMq1856JbbpBmRL7YVpee2Q7tTMHGS1JvLiH9A70mBPu45nvATj022fCGlBpkhPy5JGohMeFl81
T/zsaw95zO67fRAM9wNC5Wlb5DqhR3kLufPr/k+VaIMkjbn9deJeDF2U0GvhgU5pu7+N4Hxrw/RS
FYiZF+WKF4SLeRAVKgYm1TSj382Nc+/ISRk9MqRB2moZF6XOXRyEG4OEAvgugsQoIfLJwdcT5es8
fOdHvp9L0NIQJRc9EIfLHgbWJwk8kt+kROU+iRmHbtWvFCeMRQP8YOd5SBsZJbBhHi5BLXBj1SWx
lEU5eVbW723IKcnTXYHLDB5fnTCcAoSbV7SHUruRB/oDoVSjXYXkrMOUBru5yjnqHnaAdQmVKaQm
+ABWoWtqVK7WKciOqJCnmuN0Y6I9GXANulXr/KTBYw12bhzZ8ldu7DZyof9wVlsFuumrC++eb+lr
0tnaHir7qvB5SvPoIgYPFsL2cojmYlEco7wPwhZ/mY+7IU5NFBUoImNYfJQZhy9YagS+xZJg9TmM
KX/5u5aOJ079aoq/Wt02uhqHg0odzY/kKfZ8voF4RGMRhYhEKRya7DerEzdatEJdVy01O5ObjS/3
smyajatxNGlfDKaFBYe+DVy0MQptMjBbnQf1vEuHcw1yxHAbllIgU2uj3UUtW1hk5Ak1xKlTleFw
yKx7z3gcgeYfWRvoKJEsIoTse3JOfitTrHAsmUHIVu6v9MW1iZmo2Gmr02GbmZV6VO7EzmMApL8Z
6/4ViIJY1ifI4yolNZ9Wthv4jIGR07vQ6b8aaGTKiJueq3k3qZ46r0F8+Cl9HVGBSYjBtqr2Z+Ga
dlZ6M9W7+cJgu7hFy2dkHmjVkzHdf9tm5yhlZPzg3ZcCn7RFSJoL4oG2ruY2ohnrMNb+xsS4n8n6
uLJNhGyjqvMNV7j88JKDzi4T/gBo+vL2HZuWWar9ad7pOnAGr2wUTBOIvfAsdYCgmca5ETSl6T0H
cqITL0V0sQ9f7SLZmC/immVTxnMsiqTIOSdVR052syRGZMWmYGF7tF/MSd1LZoEDvUetSXmKBiwD
cbcNf42MdPiEHo31v+NBs7GpWTbHQkHsH/WAwGG6JiPWQnWsexAVhoyjniqURDv5vBCx1la/RBQ/
7yCC9v9nZMyrNFmFlghmsOv5uzBwWwpcVTpXBOOXo6Ld1F0WVIdR21q7E0OktqW3oPMLE6An5Ft3
ciMVy/Q05Fwcn+1ikfLgJO1Wco3HaAj1d+zSoRWsFRzrv9LSOBdovjcAFdckuFYPn4NRPJ+0yOqi
s6Hcq6qQbQx4S76lMh5fZ+wQrnyyQd2e1ewI6+BquiaxYv8hjxV41eT4Gcqqy8uaUyK7uPxKLj8H
rpAZ43mApTYjGX5a0CW37w5SrK353pTVTu0WEjAIaGxb3OVaV5IpViwG68QD/Kw8tBIAeL669IzL
QJPcFWTkkA+fYD9IJYm35yKomxjPRXD9EUkP/AGg6YIZkE0Y6LpXECZ1/jcuU9Dg6MwS8PD0sEIy
jK+pky9xV7JlHr5XbsZgIzWJA2oBASyz3yEilpaT/eoyJQJkCi4oGg9yxNgKombs1waVfUxWuv7E
vZmWExMYmODwIg/i90gLUOGio8/Q4GhvrcdCNeCpISmPuVQsKmjCVfrnyC9GWsxHnSZ5ai/FNjnn
4owRsbPqdZEb7WadR1DG+8o5j9Kd4ZInUEGojaEBwjsMDNE3rz3T0VXlOSX1mCXqCFLcQgIxgrgV
Oz+z3PizGFRW5lK8SqxrmBuscCt5vA4ogg0JrIrEp0DGd7lcKrzXQ44+rnT7mJ5BoiruV0jENDbq
XVTAhXiZHdnbXcGL4aoCw27/wAjkji10NH3il9dh2Gpudeq4Kx3sIy6NpDBa7EUTsA9jPB6h2asy
6Ih9e2UlFWAijgDtJvBdLPjcxFcXUJ0Hlvf/p3hpPP9zbRCq2D1BZRWskgHAhXxwffAiCa+7Ic8i
LWHG9LpWcYE6dLne2xplGauBL5V+zn3ICrxA220+ssGp4kbVA9zU2hz73WnD+yqBmucm++wuQubG
TQ89j5h4s6z5umEOzqOPK41yhNtQoMWtC6NPmNHs7x6KxZRAlxncCNJ/PfUqar1EK6ufiBW7Pdwf
3a9iIV9H3cLBgn7610MgGgIpsI5PddL3iN5FGzSHm3Rci0aSy9LEhdW7On9pUt7Id34J583tJtsK
iBlgGwlbpW92matr5QXedjI3fbCcmKRcyY1E0zz5SyMz+w8UqB3zbmrKPRcziUy9/guVAtcOwoyq
vjogCl7LxozdmIbLpm2VoyDzpq4sCP+G+PxY9TjeRBlNMdbgLJt10qppOwpJIOPXtjSCFAOfiYPE
EjHXnHq76DixcibT1acp0MJ0qWM7oHynOwqvWIBQ2EK4c6a4MLAsdIo6Y69mUky7jR24/fJ/IT7y
05N/HrnegJPZEKl0Idb519cLNqhV02m1WtkPn0L18RJ52xpmRQI3YRh/WXRBV/d8JNzkul4OB2/z
hV2otjW/qbQfveahq5PsarCDpflC7VI4mqdn+3MO1YJSbCIH9UB9ne5qr2krPQ4FlY1xX7caH+pV
2QochticEK4BgzIrl5XeIwLrRQDqX8y3LM8+v7uO2ndgQfNYhXr9A52MzUVy6prxQeL9FPERMdtS
m0+c6TwyQCjha41iUbvtWXZRvPnBsLamy2fNXm6n7g9Hwo3A8EHhbMU82mZjXvz0HJKgKLp8xyTa
LWCZ1WI6PsE8hX/Y5ppTHxziIQr+kuWPz1jQyx8nWt0D5z0WZaVRxS5FIFLVv0mrdvVPx9HNwZoL
52JEw3gOAyM/qZEu4JPlxGoKs4KdZ/5PPl9G471s2QxE/V9N5mnsXydmLWwdihyAQ7S89lLmmIno
T4w2vKsmizfKwUTdVtjj2Lnp2i8zUHNIraECBQYqis2qTobnudx8iB9PSNekZ6W4bTXycDQdbmom
4SYBbI7Nm13R3riWqPksNDlZy2r7gXHoUPeTxXXhC4zK3O0/N/q7pesYIjrHlPq2OAVJ+r6Bbg5M
iW+M2EBZe6ln+fvf0S4bTzxZR1hLxfd4jTH7MAze8EkF2rvVLs1ekRWCZasZ7tTY5zCBXy0D84jp
GyauGzUY1+EWUKdDB1cikvVSGcoRJyAoi+J9OfEkkRSI/jQjaRd4n5Ne2gz0lRLceh9Bbprf16+B
iQmB1LLc54FyrKCK8VDa626Ar/MemssrOIFCJ6aCJkLIv2T30NAVmEhdm3yqiW7f9pcGYjEzxxuG
h2q72PhlScjbxBBApDWLWzPKJaF/7QFbOZodoUg0Km1iWqhnN1CtQHxci3e53IEDvA+27hhF9GYy
SM4zdhaDlMXmPgDmkbez2k5+TT3rUzV9b6J72Ep46O9w5Y1bKC4Lsq1r7tMiY5HDCaGIwVJDXW14
gl8Ru/GH1P9GsjtHeCw/hi+9fyw0wA2O/AHf3J57QKhPedIbAf/S7tZa+JOwv9n0Qgw672UIaEjT
fqqMPbK+cXvYrAxlXMwUu5d+ntCdS0fumeO/EaYrhWXz76bNZ3/2oK4ANMrJyhuyWnCVzwiN2u54
8MaemEBT8z5jpzKESsyD/D6K1BL1Tpr9YGJay1Ru3Vn8BXXQbOeG5bbheAYPtZRFBDjSTFFvylG9
NIh7EE6erQtn6hfCUHJH1pqlxR5gqNKdlSQ9fd7epnLL4KkuevdVvhmLplQuVkHIPj4SdfmY2sUs
TL6e2TqIuogO7Z+GLoyHNHHaGwc9bEZi+Ydfyu84YB5ckpGvCJSkWPFqSsURV0ILHjTV7Q05B6M5
yObfywtJk086fntrn0OaiD1OTwWW+4E9aQns5JtkdsO61Kep6viOQckCXmNy4QjK7sTs579INXYx
Z7rbmDheT8mhsI7bOtkCS/A4noWBtIRWx+MaNk2a6NAaiV46V12fSrPtxxLHvqt+zWP8VZXZEz9V
xVVdjuttL8BPlItzPYId/08m53RAiECFYBUQC4bq86e0gG1khXY3B/B3a7b+1kvbk2pgjlp8FNJF
XWho+PemKsmP3VPNVEf5vz/GYO1tIs07hjZJAeAVpsN8tMTj6vUxHTsqrxoSvq2zxdPDkldrwnVV
5aSi1RGbhrEIE4cN78YR1IbXc6qGVm0Z6x4Ea183eWxvDjhCKX5mHNmF09OWak2F6mw4WTpTl2mE
hdgAKICYy6klDIH/VcAlskeaK2uyICSe2B/SNs3VzGFVS6lSONWkEOzGODDdxK6uzn0iX4uEr8cW
QeOaPNoz/x7d4vvbrzYPTl3IF1a8VwG6IeIzDqpLVy1DUIwrdceCdZPz5WnXZw1K/8qi7UtJrIqR
BazUb2Zg6AKQMOo1i8/Zoy7YQSC4MYJ0J9ehW3XhgMd/3WcQ7U7XEP8MMJMpHDMtBoXPgZ8n8A/Q
1MUbj12GnlllBp59eSYje4bV6kgXfP1yjvXw1xHyee6wa6RG+2Cc96tP+kvrWyKWorhti8nQ1wXW
tg1kUYkDLRJYSij/d6xPnPumJjfAojrSmN8BCCxe0VJBm9M7jAxhWPdqFsVdZSaJBBLv4HAgmOOv
eD1fz9cz24sNKqtloGoqzv02l/9rfYMOcSpGInGdBVgxN9Xu2rAtrUP4wYm0CmJWt8OUBCFomKR8
PlQwcI3d0PgJv8Q2DXOfOIAa+Iizv+wDHQNKGm4okXg47neVVO9lpk11KOIuBOxc9dhAQ0N53UVH
5b7eZsVpvlMlIMbMfPeDDkHeolynw6nRSrtBKwfve+FgN4OWPTILS0vIjMSCONlcJKWyq8LinTjJ
bJEtfnYNsEH0JdMuKP2LaAdYIpgWCBv/AqbeY13+zb09Og0ZFcxEbBQgnLFcESYv/k+dT8dXTFEr
eWIi1YbhwEnCit/A2MDSPsWwDVfRBNXTm1mxozJsY0EOu3ri6zf/eCbMZEoLYB5GKCdYnHuJdsbo
3Ionn/smDN/GON1XkpudU0gsTLJE9rI+cxXdTIUVr0TjtLezeYySyVPJzpfUE4Bv1YmSM2Hx/VDB
7kGajztJkcPKcIN+ox4GqyTHwQOFgEuYAS4+Wk4PqlIdIQASqgpqUPsNCuEPPov7Dyxqvtw/prKO
dK2w8XZejLYK8IYAFbEbcQl5FMLyKStbMikfhMXY373hLvFFbd4wyYwg6tzzVYONHS4/y78Knfiw
0tKyftFNa/MgeImRCJDE11dfTRTLmatBG2vbbxx+J651Wqos9ybgM1aKR9f2NFQRk6BLsX7cmr9U
2bwTPDOD7ABV/bcjI7oh2FjvZZEBTpgCY7Kj8LSjVhty3WYXHCr6ynOJVhSTt/NCJL9GyMtxxuEq
Cx3DjLxG+AKJOcCh1qn0pyxkRlRAnEVdQtoXYTPrt82Bg/8gPqR4S03SxYqvgiw/G5QilDtHu1rP
em0IcncOYV54ANYN2V4yYZEEsdFbp8d2dPfPJXVdyXW2Urp3LaWX83flxDmTrv7VylKNiKjJwCM1
/MDOPnyu4w56BoX0Nk8WBu7TZYQRJVy4cWh/xRMR3C9GHqd7rjxd4rdNh5+omKQgJsyswNM120gl
Ws5oMlN5+w5GJVATHRntT/rT9DyCgCH7v859SBN/P8vHzTKMrl4371T2sPFH/gjw1stfdThUVtFC
6y8q0fX/vPmjjEWwGlKpczxzu00Fw3oUXfKxEyDHkEGnaTIXnDOitXOgasSK3lhkSfq9rD2vNllP
ik1DtMBfK+O7W3+w6EepW6Vde7gSUwDaAv9BsCyPlabJcdZ8gyxm9mVMUPBoUXHrVHtq0heumz+D
HkiJG3gDlChPf8ztLrLFA/ZxdvogsFEVV0Nfdzm07WYGEMetCtFz9C5hySbMNnofKRvJhm4maShg
QFiNc6qlW20Ae9Jb/aInQ6CyhsZCVQDMRxAZ6OzarjV0XlBlglnNe9aVUN7IUgtw+uMu9lziiKot
R1Yz5n4yuYre7oN1CVgMXSan0jIDZlbdQyuQVW0Mwwgx2PL0oUNCSd6+u55I+WEEYAGoupand1Rl
+pRPHa78IpkdAqeK14gvNTnMMl2p8AmuvPBsHCEJn03bgJicqFNgz+v9UXIw/SU/KjMk4BWHbzX1
uc3hqxIg9WRBIoWPogiUxbtN0c3YeL5mjYb2gyRRhbq3ha1WisSTOQum99TK7/JlcqXzkgGnotYk
kcYIpNIkD7IDN+D33TvBgevADhwJU/cDcaSypkF67c8Wxm8THzHJKx+5zxN7MvbzgUIp+UDfmL1v
3hbJBEaiXGEeMpNks4WmlQcdvOzKKkNUC2qGrYSlmROQianVnMsJ4NPXlIQXdv+Lnjb1PFVdZiB0
5aIUzHi0AEjZGo6SXCBMLVKsWY4fDA67xXVHD2x06uSOjTTbrHBm0QuWeIVdx5exyDnvlfirII7v
oK8TXvG3xXfZByklYS02OqCHFe23ZONygM9ScymMY/wwaGhpzT6hFhnGLiUnrBvQ3Oy+UV6U2IJc
lYv/RUzWIcjuSG0jkUQyatyogNiAH6zCvamx6wOMIFYwO3q5NsQrQZykx4zolan9lb4XkcQFXvGM
cv1yNxh6Xnx45wyUj70wRoUlpoIABcBaba9L6cc7Mf+t5uMi5zMxBG35WBLZJrjaq0c0EB0h+7/Z
lziqA0s3SzlNtgLu4NB6gnSdA73pyX1YefJKvBLYeswwSxaanXoHievmzJ3Jnj/9s3XH/+Syt2oN
L3dwMfX65UqrAMhBgNi4mftcTe3DsvQw4DBOllPBv7ccU1Y90RMNryjhGy2LGSQkxRn8N24W12DG
6DiLCfDytpMBLYYdd/2Mr78J8ILA2e9/75M1pyZrrSNDib5fFlvb9zfSFvZN/VaJCYzYpPurbuqJ
y0j+UY1N7P+HSN7S0XbHiAX8zDsRRxDa1KrwMqvcvFEDdEI7qSld9wbyR9Vc5OfB5WcABfeczyGK
QfwtpUj9AmLrxDW1a08od35EL4Xdfn2PIDrjitr1nAKm6FIdNL7VJUcYFuURt2+N6KI4puZRGeON
J1YcYMGAjlIQMDF3B7I3QKweF3nStbLRKC+ytpX5HDXZu+it/MxdsZYGSzvMGjfo7a5CBFvezj0z
QsGM3QaJDWF62VvrOS90xt6a3hHgWhnTPnaKkC5ulcw7qQAQ+MH8nTwFLcMy8tIxGovdiVE1rLtd
RHgM5/UqB/cvwFtolidnwoBfheoEE105HZOAv4SKuKOjvNQ+H8b+vL6cqH/k2ZDu2w1yzQmthSC3
mjdPSi5VJEv1oZ/1Px2i/6XYZn0GugEkysAVcVYwS6pl+d4pBIJ4M3FCNQaTwM5mIqU67U2/GzcN
WeA2pMUFFLX50UbUgMSJ1YbKYzefIsvBlDPDZm3BAsK9+HMhCxYl8eBc0KzlcAcNw1SsG1j7OcUW
ZhzcWF99wi8MlI4ANfXPhpMikvJxH5yIWqldD5JBcVPyZ4A6X5yZiJD+iqVMg+9ZXnGvTLutB/q0
L1oJ1H1Wepk39hOS1haXOmcPERRiKlyHnQcDRn7LONip2QTsjUZ52n7k4dTV6jr3JczTHvFN/MXO
kYoTYd78ifrOnSqQK3EzGR6zDgAQGCcjnBqY1Y0iL4oDlcBf+y7PIvbl8kI1XOAQLayRDG9cVlgh
H1KT8RQYNcOtK8exJDGIem0TxTO8uH5gA/bQuCyKeopO0AX1zq1OvtxkI1Rv8rfK+kwvu0KS432J
5WJFzTgjSyjfL/P/v3If+eayIMSovayp99TKVKoe7EdpqRdJe5gIFQgBPOGyq9FMu75kEFESN4fo
Bt+bTh9pqJ2sjB/Onz4FUvJ9PDKXs3t9gm7cWWRimTepJ9N6aFD/++br9LuMhluu8XOmA/lokVTk
ZkuaUc4tsqTl9fCu5GDQU+cVXyKH4NxZhNNfcycqnLYCRlFZqseU3tJnRQ3asBCA57sHcFHD0UTP
zSB/AlR76OglRgQRCle0aP4Ol4WEfug4qu8ucoONVDQM0oOqZkDLL1o4kSHRPjpHCm0IiVy9SckB
9/AN2knkLDC/SfX9edJYK6YqvJ8Tf5rUaxcDJdV3m62KJr8fqV8EtUfl1HHDDWVBBBt+Dekas6uI
XVIo4a4r+US/vvzfht+d0fLomKyifIDOSiAI8dkfO+LI2/uDWnjyJlDHgucjoR8wsS5gD6jlEYX0
QVN3osdjMmWQ96Dsrw56kKvJ+5MOdkQNw0QrNe12ao//SLglt6QnUv5J+1vrQcLmiUk6rSXOxfwv
ajAjmptN3A70OdgdvLynn4ZieoFN4K5wG6VmErnqDCTs/bURx12at0jlljAFlcmiucdIwlkJgYXP
lt+tnA/Bbf6hzktAUSX2V7K7x2XhiHQjOogSKgN+McKgjbbmSsjbvF8A4KLdni2Msr1pNbotSHD8
8bQHCoa3MfbtX4rOCQhYjb0qrX94g78d//ZmL8Tw3B5J7DD3d0wiykU5vu5KtdjwVfEdKxOHGHZt
CaSWoenHclhm6yIc2HGEcAzqqC0daC5RRWT6+la8bdcNHjd3bYGbsP6u4l+Oh45eynGgHkzmLAHD
r8ryWwDFNB1eX1fNmxF0HYmc77Rcfv7k56YoJYLRt1GeCyRSchJkFCDOElaju4djUF7hXzceFC+v
0k/LOXjFI6wqD3G0aa9S6n+TMC1I6NC3GITRFkRM7NIsB/qeu61gd0LweiaHGIg3Ba78ZgAvBTL9
cUaz/9ZqbB6bSunurJvi9z8FpquW7rVhyQyQp7pLHo1FXYhWBvW/hWlZN/4XJjrY7RitgV0FtNu/
hZoxso/ozOblcICa+/qwb8wSw1zKB6cqgy4i1iwp9QssQr2PatcPvR6LtF9uv2531e7faHBLqZPN
UPd2UAoWhGsx4dqvCuhhDCWGHOCA38ApzhTxKCTqX0Etwc7lMQcTcggo+adC81dpUiPfsBVyOpq9
Iy6h2CwpQJPjzqyzHwwWgQBFITibKHg3Vr6XLkRFsXIHrbuc+H3PCycvDf00pRODNYjOBsWamybX
9l/6pTY3ZKpL4j0sgzbAVu5YoF7LwJ6de6eC6QZaKEosXmLIRxtzzc19BUTjZIYJQe00hPrBnInF
Q6HCBLPf5CsgHkEp5EY6lbglDXpAdsF4TTI+yM82kJZqq0znxYH54uqtcgwoeEbFWGWt7zmmPrMB
mKR5PuzkrG9SXhfne2mErYjhbrIPG5y7Kqj+lNb8+sn8TcLpFnXmOvbPW4EcxazO95eE2NRPMEvo
jtRTwZRGOUbIry9w0r3S0XDSy2A9AFAshQ3HnAE2fmRluuav6owq7kP09smTd26efvAO0Wx2HrXd
rzSJMoKP1D5tiHU4QfThff6Pdm5nIWm5hNBhOxymNyTvgugc7X6fhROi8uimygkaXoYwsZKdzRA7
bWTTmYuNsV7dWDcXkJb0DHpeKrzzha/gPeKZ2H964mer9hvdd19DN47OjpNA5BZ6apSilQQ2TcWu
mv4qNnThuL1VJ8UqvL7XaWayiIFy52rgDcpAUhDqKHMbTq1LVPB++jV4Fjx/GXa0xwg8H11j866X
V6kHB/C6yeL3IXMgCCSf67QNaV246w1L/LLdzKDaIwLT5mt3VG16CxvKVVAVydQNWMPoVRqx5flX
DAD0goROHQFUYXapWTkVtgLXiy4lT4q88fDf7+sovDkdVmCm7MDcanuG63TKNKEUxCqcCewluVPD
hFYaFwbsdniKj+q1/59BSq4BZogxuPlWC5TB0Vm+d/GvNcGT9dB8rQSn6FyokB/YcOljxFrO85mK
VIwGyWqhZGIXpbSiCOn+5MFoEYopX83mtF5bpgWZHWkYB7fw5eatuagPBVyMFxm5IFTbSSBc++QV
aZSA8e0A0qQ02psz6VsiL67l+EAk8sk/RzKWuN/5Jg7TQrUlooU5A3vOAof//TBFYT58JrlV+Kbt
FMoexJBZyvvM1iRISPg6Dp26gP1CkHPEEIPAngDsrzjcADK26celGuYgJXNmLw7PMwJei/wMiQUS
c9hWSROO3lhaD7lLNTqGJ7bdDWlyceDYfx1NL4ZpXsIH5AAdzBkRMzAPg7h+Jsk4OduYHKXwbTRe
hoTUv0nbvVaV6AGvD1Dw75cW3aA/KXiktGu/nhR7lzpUmJwX4NukUvjxtbZcxi5V8gEmQLVmFvIL
MoarYy5LV5W0fqOHb/ZWkugfb160+FSCsUeX9NB80D+eERFL0gNcj/2DVxu+J6+u+l/4dgNzSoti
G0P6fNQBrdGNAtkDA5OA8ZAWHYiso5aNx5M68RkP85Opmviw58lOgrVrxJdFrwjxNg3BpuXCEztd
jeVWc0d/U935GmfD8UT+ORPzJja7IVVCs759QTVlGfcQGWfVbAKXz1CVhQtSTF4v68j2hVnC1XdW
lwrXGqDUxwpzSKW7Yv0nSYWdlcF4JiHmO1DhHf9UrVetyzrdzm7ieROXJO9XObY5gWnwilwedV8Q
JoEhgFgLX7JvuPhSlO3WvHnR2qK9LRnvk+gK4l2Mit7WWgU3q1hA0JlzADsf9kg/9TtkWrvxKXMl
KXj+RMe0BrhaJgnMW15AihTghzhwCiCdjBLePb+Xjdn4fzWi9PDub+wi1iD6+UybhTfcgM5orLtu
cw2Dlvxi0CwJVTnaqa7pSVNfHnIKfOPJLwNACeVh8uJ5A7KNOuWS9mcF0lPUXwj9NFEeP9UqaWO4
VBOviCzKR8qqVopfhqxuG+57DGErwEBWqZsgyywxbyIVCofCMOkTG25fvsNDlTB5kf7GNvqx9S3T
WOp5jaPhgxIayQEyy9OH8PQF+6k+s7OnfYuuPQBq7+OTpPTzMbIYCGPm/FiH5Ky0SzrJmLYA+/Vy
TcLeUhQV5dSwEyQhcXHFqhGHpmIstNzjXUQZ7LcORMjAMLJX7osgQjqoPuJ8OaxCbzLGqiBo7EPX
Q9lp1QKTis5e9xkJsr2Zc7lMMJSUV5zp38F0zlVFM468R1tDqt/eS0AOM4Lz2mhc1xa+tqyh4n02
mgzSWp9MPwSW/wnIa9mHOtppsNJkYf7AJleqvj94quyPoX3n+HYuaKmljncTx7bt1GEktITJBbXV
9p+sZKCgyUf15tyw9r4FReAt082/Bsz0/Q2gNIm338iR78TL8Mn6BVTKZDW0emcgL+8iZOtHluUd
j+4TlZZYuaqtazLUkNGle+aX8xRyvPPxP4U0d6oJqjat3T3fmTd30wLGNZ+G58A6gsrr2WUoLm4+
nqsaERKiqCzfdNnGZfkj7sUefIjiiVw/b4hvuAHBVHTh/m9nTovoMY3Mhy77or88hRqdfypWAAX+
8lAQfYNEskssAX18UD3Q7Ga10HibZN/t4JRFxnE4iBU6p9NfqPt7w8FmY3D7AV9oQPJ6l/oVo0gI
yBK6JcMOTaTK/nCbaiwTschrWQlqYrVXIFGHv0CHNc+RR55TeiDhDYpM9Fnbk/x6hON2ctVjDfJQ
QQTHcodJZBNglRSvoJAy34hZXZ/MamgEcDkBn7H7UY7UQ6sUxzss+CaiYU0TAWfVt0Gsv1Kitodd
qBVa3Wkeeg+3kNBZsqae3+8qF5BrraUtc2E+kEQMg4PpiZ5ALuVOIUgYldQfysOH8qNnCjvmQxLK
oLlOVahHcEMxgU1/0jaV6oPMCSR0+6wCNoMPoVEI5GVgZl0cWqiZJW90tApxn8JxBblBTNiZ52En
+tAxIe3z8HZuS3ZBNnEaq7/YXreyG0c8h08OQtZa+Iom+1obuQmSDfJdCzJH/0QUDZSSEkgEx8s3
3HuoRzv1HX7OUVyp8Uh7gUawfzVGyuty96nzB1cr4is3ddc/uhAbqoNhlfO2umTz4OjYMvpDrL5F
CCCNTjnpuSmAhcsS9BcyGw+fTpKclC2yMD7yCRQMZC19ngcSHZuUwefyIjbB5uHokveMrfWXsjpz
tNoKuPbSdVIDCt3rC0tEmLsK3OWuyN7Uweu/NsSdt45rsRdmhCTrzACarh8Bhjvg7fR5t9gjH4L6
Bqg4XmycsCdTobWMWoVJWZbF+MAzAsLP+4mu+1slpema8Ah5afqi0JL8uadF4Qw9M8T8ayhinPzO
L0+bH9HUbfSv368gLtzVcCj+YT/quipt68O0jB6cBsH871fh2x656tatGy++gdMlnuY8S0tjJhdk
mvG/kvyycn/cs3knUUCzo0aaJdFg+LXaRV87kO8fVmL61XDsdpVMEpqFLKYem5eQDaYgZkmrDJtl
5qTEqrtCKikAZi8JWvy99BcUq/giypF0xzkV552cZwx6g/V36WBp5rzekZdPUs0/po6k2dJFpkFm
vSTGUSgWlceUorydMxUAQbduR62kA1TebPwBLOOvK6jc739E/4aDHrx5K8AzrBdBIZbPxokzfYAr
Jr+HlcYndbbxSQBq2e4lzK9olUZ6bMRT618rB8fwNaecX7h53VetTm7j3IYApa7Ukot74DmhYSHt
yw4UiNpXKGHDheFC6rZ9ETHMpTH2IRj7touXMV3udGzNRjIq4au4vhf3WlIxY2gllNPu4r+6UlYy
UJIYmGBTW8UecetbGu6q0lNTJo7NZG9ZDrEJYrAth3hl4trc6WXdQZ1k8MmZ5JrvMo4JIrhxoblV
OnHAYvVn4G1qsY6ZuQQW4Ai7abesZy5iJd1I8VLVYIbjHE1dpBeLuHVONhkz+pvJU8JngeObNrts
14FqaRRYnmSFQu/fJIWGP5qFNodXOQeDjuSfLAEFUUo5uetoFtZxuIogxg2HB1ujXEQc4KhZMWEz
upIJ+y5ereQqHhgDm5obaYpuAaMyJ/6mH9ERZAR1RqND3cZ5baPMw2cQPdgUtb2bxzFqjBiZgu+S
DKhqa7duNOsxHXs6g5OKRKMBfaHsd9nLZTgA2gxnAGOGu71/x6+Xer9GoJzSXqxwbh78kNJ7RHQu
INsGPZCSkX1QWeEPk24qymNIDbX4YoXQc5uklDKqM6gAQ9iZi+kESNVAPc/ho+mO4BZo3yOyUmpg
f0F6RTsRZi/6k9VSR1PrDxSI40u4fG/DvI6UfazBdwpkz8DRFJPGaaFDHjNoCXk/BhVCXXd05fMB
YMUEMG9MNJcaYg+b9ulCfJJUpx09/pXey+ON2X4PdfM4iMIrQkh4RjS3E5mzKeASfxEGBCxjYAv0
ci5XaaazoLYRXfX/mfJ/QYPGaCGKR4fVZd6wTe3pUbCzLhOAFAu+ooM7o3OoDroAI11TcBGMjI1w
YwUhNbUEeFLSSSJwEd7IzRcHqcmQMRKqREy5FojnKdinSG8u0emwvV384mbUo51sJNVgVt7Bb2Lb
R1BSfFAJn3O1+yvcX+5mzQC+NJFkHdNB2uFFPbdFdzLSR0bodMrFvLQyj4PY5YFrF+jIbmLZbTgg
v6kVLR2AL6WSzmjgXwsNFF7Iz/MMxJyHBy/0yhKn0yuFbwuMcDb1gzPgmLzVfspYbarmf+/R6wK5
RVzI+GwlPrBNhE3hFfpaimj/5F5BnEFDrL+dXXoRu18eG8hh83XAjgJ/yJTWMZl99TSeTRFtrLXH
XZA0FRRnJCPsZfGRGVQGS5NgV0gIS3EWXzp/MkKDOWJWYgyGRud66SaF4DucgEFnQj+usvFbBJ9E
4/AJpJJAiGTAXjxnsc6r/qyckZWGCFP0nzsiuv4NdRdWggTz62IZQ3RE9nRUX3NwXzbRGZd0us0P
+tIdDv3hmA4lj366qg24GxNmXvCVO0GFqkB3D5sB3hcH8G+wcu3XyuKKsR7jfcPyhLZ0bC2u7RIw
oiyPQRtY6sAp+TLvEYkflLxGS+ht0i+iB7oqP7cjH2OLTrxQPufzANsr3eENGg+Xz2PTdZjYiu1a
TJYYPrsuP3mvHAdEZAETHWlleUJZ7WhDRbE4rnDgmlfH/mRRlaCmQycyW5LvuJMK60FAlCqL6q4X
3oay9dBXjUHnoAOVIo1dqATIq9nYoNNzmbhwIauW+vDr7GfpUsGjPAb70fZFhvAPC7LH/3yPGODX
WEORW++ndfkiXX0ZUh1CIFXxMlKAMBb38IIYIAe4g67RPHRXwk+6161d784JPNUmB9CbCdncZwcU
a4uNkHA6lOkwc3YjssRt5JtNwmVKfiAIwCLq4B+zPQq1qtWlyU3IYXqokJDjdvSrlvChF4L0sn0x
zYN2VdD5oXTBkm4bKk71x1s7QjBRrDglLyKhwcxZWjHCJYhpoDMCsoWfR4qBn96G/YNC3NjKEVxR
cVrW0IFJ4qY7dm23eFW/G0y72xPPo05i+Xoh/xh6W4XzeUvzkRmKn25b/Qr+8r7FDkhMuI9PwQ1T
9adk5E+PJHHXalM2tUng8fkOIz2ib/nRYv/K/M4mp3nJO3RY1xHhrq07LwV1cRLSHiTeXacuvfEm
X5x4IKSpB7v7v+DkCdmGjrq6FnEn83HjxdnjRsVxzDi5ACI5nm4VSB6EMUXOfgXW348GZxHu61l/
q/98fUgg0QMSoCzlEEWByRU+fS0TVmGf1ZaRTM9yoNfnQmAu6O2gGrF5hQOgXJysTNfSGjwBSLYz
DfUhZE+0dkRG+IsvBfhpjcvao6Xajm9O3vI27FMfDnBe1sYSBqdU6+mFueYXrF7ixqgldhdUhJWc
wvfawIA0SQ3dD4fgQg7Mo0I/MXEyfYWdyKSbRCBd5zROhGB01AAJrYpJqGwGdkeubZb3ZLXYH8h7
44W7ouZbmsGVFCm91/k529PXYWVp9HWX5eqPvQ4X5YI847Cf/60E05Zb72ycGLKcMjkt1bZt775z
/RxfrJwhOivrI2yHAc4b9tOzraNnvaUWAPXiGz+OWQTEt+9xkr15vQuMS/hSryLvIeX+kbSEzLSU
tDgAhAhJDx4xPJgYCP9RVJMElWmTiW300xP46vni4bx/cz3IqcHuC/2blJjuTkjc2IQxqjAWO1/v
XDlnhfsClYZh9Xq3YkSBLt57QHcqgeYQASvp9516lzK4NYALswjH1/Anmv5by906w0rBPd1lmvha
BtbOJuk+rb6cSnBvg7y0e16bZ0rKuoha136lpAE5mkeTNHtUh0paZAYUYol+oTMqru7yLEDfWn7D
w8tFuS2XRBWwuVBaF4Y74+7mhyx8M0+Bignw+Hurm1+SB3DMLSrzZ+NfvOspgnEVO99U7CbHGhZH
YRe5RBIyxEsBdIwZsA+tqrsyf7XQSR0IDEuqoC/b/QZ0J+Jt4nLq/UCJMR2vbPsGmM3Sb4t/Q3xq
2W0V86tAm36ZGk6q2GrDmBn0QGcYpvHJH+Ncl18vBk9GtmLVbGNWQO0FOOkN6E5RIZzrk0LwQQM5
S+4E5MQL2y92PhYziezPCTP+Ik/B0XZITNZqUyHY08rkzXz5p12iMxIJXa1Kdd6LqAJmPg/NhWxJ
aVnTpdBCL2RvD3pLewqYWFcJwT5Zit1D0wOP2fLOIpVigdXMEbIJoYt+hg4VmaG/T/UXwFi3pJQ2
htqB53+sEdejFO0YENmNMNjyFKFbsIodY9n5F+Ifs/GEY/dKNlGEkNiVsmdGPrAjypncLP+y2Ieb
krIjeDtCOJYebrTN8+k/OSP3ojl7jHxUMEgpg2xI2aKBjLOYTor0mQzjds2y18bLDCXimUB858Zx
NDN3SnKVLEdQaHng0DgLHdoX49NvbVswZkR9TXIYaXYro8BBox/J7CWXuowjznOmB5U1rEHkPiWZ
PMaAJoQgG8mUlDQmf13mlsfcBYGPANZ/fMJw9s/7rwb3I3aUpZI0whDe2RrvB6fxqL5iisl6Bbg4
5g6msBPzo/7yu42YXA4+SrvTClKJ93n+3kM9P2ZpHIB3D56fLkgevOS3c/VpXaXKC9ihB+63RpgA
ijE1zjpsLup37PN+sXPJleXXWeObgtMRwTTY8EcqpHfQ4j/hDhHhTDZHYdDs9CBbRRiSDRlx4Z6p
WH88uVZfTAuTqu1+0L//RsNHuMGevnv31DBCKfNM9quaxyVZF8Jj0xQlm5Dnxm6roC6HTqoYFca1
tgEhY3zrJYwSVtIh3GXQRfr6Er7vR8dJVadIWX01eBmXwNkn5gRLklxed+6tLZDcsxkf798SBQF2
qsLx0RWCJpos43tdg1OvoD1n4PGbA5eOoB3BgznCEzx3oCM5B6MLj0FRXTEmCTF3Vx9tGyAmdoq8
T6Dz8isrY5FYk7WRSVPBVG/lMYXBL1XWD9gOWGt8nVIskIxxOWWnhMTRXzC7J7bchMWeNC4hSfMC
Ju5wX2Q1RF3GKN1fvIT9lBrt7nAwl6p4u71pmmvP80EbDET+FeWGGfrL9DOhNDxrMSY4DGFoocj4
Grudps9vtVG2gW6y6kOynV+66ua9b88z9DnMoiTLaVtK3/M/+a4vR+iO1EfQMDdNy8c20ecPD6Hl
7ELpukgHwuSASQ/Lp5vdePUqsgy3LN8URPYsmdJBMQOEpve5FqUkTNK5TiV62m0Yl0N/Dg9z1uq4
aI1WNVKRP1cUFcRj1VBBW/o018pUww9zuZSrjJvNMpbCLuKrBNnSL41hQ7mX9FeNKaPDIG15NbSj
L8blCSfBOKKnYWu8ZcF2ni3mD4aCCRmf9fZcHCYtoXkunmMQ/zByfm/t4RvNWUi7tO2uS68T3u0Q
phO28k5gxrVSQMzwlUdULMdcLDJ8cOPRQWqadcJaOwY4bPk9sYTaNh+PwT9O9C2pzYoMqL7ZxRAE
qSWu1PHiFYXuw8EOxpzqBPq9NSe7lsY/oC8V/E1+7fIqcmdGjivGysGONPWUjdFGL0t/cuoZk4Gc
e84Ckm0u/qXmURV1ioH1LMpnyyHUxl0v61DphHAilmGyX2nJGrdREuy5hSUTAMNK2+dauWi3mf7Q
DWplEQxMxyzRoxvrd26vj5KEUB13xhH9hBW/MKgtmwmo/dp6w8XBZy9mAeSloKENSBQjs6TIeJfN
vqF/ChfG7xM/cnUxoceQL44MELSOBBuUu0OhR5T+VwzLM0q2hPXMAYaibyj8HM0nE8m7MdRXyfXT
E76GCSa1FITp7dkRBOgBPv13WWeTCRVHc0tCHIWotu6817x63HEZPUzmw5NPWJuM4QNqd8pgWHeN
oPYdcKx8Ad6eTtlCDLAkTBdC4NHYcFdRWSPgp099iVedcUFJWDhDpvnKUgx90+X7Siz3fuoalyeT
OiGGZtgliKe6lNEdKFByHSDOPKcebXU2srcOrjftfyWI/ziVQKOZYK0R4lpbWNHFnUpHHFWcNYMy
L5CkCqZak/qOEvkKvbnFH98Z0K3Ss0yo4IcFdhOsyFZt3J7WBazKBiW4rYnzDJiVzEztFq4K0bz/
fct0VHt25GskfPAFCvUk4Hjt55QF+pkae4lhCETP+KXVLim4o0DUyPV56P29J/+DJ5WBnelJL1Kq
tCPDVfsQyT0Y/s77MtwrEZoz6d0iN04CMYvxldwtfrSqrqReJwkUCXzM0WmY0cDiAkbC1uPxlgJU
ho/OfEvDD7NMNe+KU4+wsosU7v8R21wZyWAluLAmVVTRb8ha2xfFNAJ30deXk1TJnTvuwBsxDg7j
WjfzvaLngE2/pe4efayFSRQieNiYVDjweIuFpWgtZ3qbTRHKcTmFRux4oozO0zUMSgxGVOSea0xv
IPp/qG0EKzXBBM97g8G7LOE2J4beTyYIdo14quPP6qIoqGB7r7cMotSKYnERngn2fi+QM5TBOJaw
zrlpoa0szaIcJqZhc49LXjL/yeD+Fhi/LU3GO1/zyD8sFGEIvrfOFnKXuG8/PQo06UU5vZJiJOQx
aQll5gHFNuqaJW/eISGU0TBesMWJVkKWmPSNT9PnDP5s3uWmDhbB2fiZE/HJQiaAME9XU+vW28UC
0mqIP51XzhSSZfgFhNsOg3kHLJtlasYQiZzVOAXUGn0mKDK9HIgUpOO1dVxTtxD2cYvQ2P3oh+jY
pk83z0Zsc3Z+JI59yw5B0083abFDegzkJxRr15eFTNajw+aXvzpm7t3WFOLor7GL+6iCHHASdjoi
yX9d/dpJ5W4SonFx2tW80q8BhjSuKJqiADPxFnvqCqP5vJdQwalfVwtfZH+TdxjbnCub99JJk6ga
Z7VOO+8UDE82okq+VVoqIXGFPQvgIi3qlDG7Z6hLnaxb2SP/LEU7R14wJN24RyIb8GDrcra9sYTc
RpmFAVk429vsAkwRGkGNUQqELPA167USqMMvv+CfkmXTOpgGsgjhEdqNvIxqMNBOutifxc/CW1dm
fNlue7Y7xecCcxY+SbAULEK5MVTlLy2/eXFmedILmYuh9gpcIe553w0+rkI9Vxlc2N5PooSytUAM
xo4KntbrcC91U6A9FPL2Me0Yy1oPlUH7I+E+ckOYn7+MprugKc1F/IVYGQCkiOKha2rcUXw5pyBM
n/A6zIV7B4+xz4mq25RLg5zvOUkOY0AtDI9dt794TlXTYYrqG23XULhvs0GzSUchsKUM/f1Cy/3T
d+NT5FcFIN7hU+xTn90CE8As14QoX7xdmbmAxSFJZlLJc9RSl44cO919dIt+6daOGB6TiZF7aZJj
MqLZBjbs0HnnHxrQusMjWoANC2t94hWoOVByLx0PCpalCcTRkHMt0akflFEzKC6voBNO9/60GToS
84gIpe2nh2yKXBD0ySi0GWdRwNgG8K+3qx2Tc5PsuplzEiO7uIomc3oHPB7irAfA1LNciBySN3nL
0PzXlBgvkBDlFewlkLWzKHIrx4VtwzUhNuAcGqBUPR30EMlx8ZMbmmEI+yvC4kyRGcUnL8LRl2e7
73yYfVrQ+g56yIG+jbM5dwW1hjPc+QH8tQF3lHOLW++XF5VQY4VRO3wd8IoW4WYvDlbtBn9OZdAT
t4wkPmbKPbrM+fPMJtI0jWcT2pi8Bd8GKTNLy5GDggY/VD0R6JWe9n4ZpyJMcvQgIFlOgukmb6Ki
D52OF/1JZLXXMaxl4GNxy/OevP+s3D8W/38l8qmH9gztZCAo5RK9q2Ybsm8gKRM5Vj3kbbqKFxwb
6uEJPSTnVSM1ShwW7iCauLvO4r1EAZNn6pWRHvpH28BEv2Urhq0PM+PRd+3VyFfxUEZpT6n1B+yx
U0zpZfWGCWYQQlA6Z74PNTg6KzV7nTUvNK+hQfDDozH20okkWzS1Aq8BtnNQlIofPvA40BMlix2G
Af5kBw5yM1JkR8951BA1EbQeGGi+0hpJex251H4SuAqcB9hiBqzv+o7iwEfm1S2NjkvbDmqfyw6S
xsUxCkGSplCf57iKTTmO5G8IUj8F1u6nhZPy1UdOdBuRGXwaTVWBb80J+neM6WSevJd6cr3Z+jSS
6kGLNmQvOWxBqvK03oReEQYsML6i3cIs9UnGwZhhWWfLErj3hoLzY3zzYd6c/89Tf0JWo7iBxXdb
BXPsB3RLWhykm97vCM/jDVj1ZUiUTbVYmr+LKu3KtCmUTT+Poy7yQSYWqbu2TuMLtY1u1/TkmkNb
IHUX87mWgSqpvH7PjtCKsNe4n3XZqV/WJIyfiDCUG63+ZKiTPFfM/YI/m/YQ5g187Ol+l2oNUSz3
beMzu0xv95wW3chPzhPS01DIFqNCuUNUN/noa6AHrzwwUQHjLiSGAL5tRQxc4Oh/8JhJorhOYDZO
7DEPSiSRSmaIfg6KqgfhdFK39sGUB+xVDDtISc9XRYghPg6EEwh385rwwpj/jnxMztx5FVnIdftu
eY9nvVK2uHwiQxhGcgys/SP4bkHbUx6MKOcZnGcfcmELwO5OaGFCM1B+0XRr78EQXJFIlu/8agt5
ZbqwxI7kpw2ueW+TN/qhAF9D0oiHaHPsp0ojBy90ojjEVjvuSFts+dGOqqwuQ/9+cKr7E9P3saIr
47y3HdEcEIGy50/bIYq8KE7D8YtDihRMKITzkCmd+Wx1GqklUphGB8992kT6To45fxiLXHM7XKYG
wOmDAGvfARwe2E+RkmS3Db7tyOTPSpKrJBU2Ryh7xB6znQ+6jqD1/PUGf9avyqenMW7QyN5W/UYH
idK7U5f0p+Cbl4fMPKxMVJOyg/U3u2FriXv1DpFaL7wgGGC0EQ9otK1DEjqBWBFTAZoyixiOlRkV
SKIDB3xwVDlvu59yu4v2JJWJ8tjq4UETGZiLVbKOqQK5bgyzuyaW/luxVrO1OIQ1C+skBh4h8FBj
9iZ6yyLq2bzN3okzyIoCXE4UhUjhGJnvgrL1/Jh7hMLxcXzlSEkP6NpJQMsFx7hCX7ZGuqkqvoqr
fHjVZ8hGWzP/ujMVF242XqOPy5XhJx8fAZelWPDZVdaF3OPwe282aGXyw7AiqkSAfWxf38xSkH4O
t5+2+eJQfNjltpUcg99Pj9+5/YqZBAEqoyFT9FJepcn2YEfVgvvWpiw/lutrDVGv3pd/KE2SCkAO
FK/mnBKJ4ntCP6w6kU7kugba1bNpQ60+HgRbdyCqq2+ojH1kXg/PfOqphxVl169UPgOh4IafGR58
oIayBRzLJLF4J2uSTqsNC7GUm8iiwkInH6n52nmQcDB4zzXGaWGhCj1EpfylBAUWAOHTHhJhr9Zu
5+QV32pKyZkZTFrae/k31leDnMXa9OALK8BvJA/Sv2McSFFe1+2mCxWiqEBlgxHg61EXjwDjZM8w
2GR0U2C7SuezjN3RSC4TiFPCKTcGe8sE6UcrMWzVK5w/x4rbv5+Ec9eUozl8t2I/vWqnMggbDGFK
5tB6NOpz4iAN6QKVQdcRFT6DTTXeRMxrsFz8mKwlTrpBbEKBFbw/7X4rf6UFzOcoft4juh7DW6BE
hxyuhVHlcqDMazrPa3MdV+3ldiGegHi4LMAp3zVIah8fTvITGAK0ygyOmkM/zTEkg98Zn0nUz8cQ
6n4WBoSDvQ8GpBpyS9EOue2p2NizNgAlAoop/DuUnAnmh5rM7tOOfdzL3PQKOh9nJzweA0UiivGu
e3HwOLDrsMQOWzFnTQqgSMD1NksRPFbBGpk21kukRmUY4IhKoh1UFarl1fgzQc5kJrqCeB1GG/31
Ya8VnFGneOYz+m3VC/qBRhscQhA8nfaLVQepWpAXhEHMYMPc0e6FvZS+rRGSSqqh8lU1YNta1/pK
0M53HuxtAnFMTjLtjGTNAeq2DPDffPc2H1xNTbA+4aLI6gYro8VsjrCmKcVwvMGDaDoWUfS7Rju9
Zw8rbFJbObNWYYaypuwHlSjcrtK0W2Jm6pR9PUhy4rPJal3eiNhj9qzx6fxf7BLinsf0AhiO8LxK
6xsh42uK3rdueDOHU/JvQ9Z4W1hvNoalrHCWTEMWgoUJJnnwB1j0xzrl08R3vPdUNH/Psq2Trgst
UP48AC55+laIzF00uI0QwAM04GdDuUbFB7fNgRwULso4uu4HwunV4OQeBe0fgf2+4lOyjZvjFD8Z
aHZCwau/csEuWU2MmoL7yJQGHlSXaIn2veShUMagJLQbLXSPYwJ9rDkhdoNQpCw3nqTH0ZYWTd5I
dBd4C/AJ3b0LNHhG8kn9WRyYceqNaB4kGBkIv+sDEsJD6bEGSZKywD27MHfC0OVHf4k5jJ9TYy/n
cpyfkQ9Nk/8Uj2MFMq9ShvxKxaSHruEOnJXYlwgRD0EMAlWlTtbNcjl6bGUAxms0uB/cW3HFm2fX
P4N3U52b0Wf/FuQLoSoUjweIGc4ouHoSp+y9plqunT5UgBzFMnlnkvzh+k7YpbWiF4Iy2h2hx7mq
g7SAMEp0FL9+OVHVtGTQ4cm0q4ZIc7oT+0yLVhESkcZlnaip8TGJujWmbVVNHFFHmpiYPtgBVytB
88J3uAmBLvCJG0dt890XtL5y9C09FjavEl6MHeumaOv1YQTB3zYzmsdQOdfOjoUzkP/k2e3H+KD4
X6M+7+O7A2JcZzlrNU5Mk68hx3ZnnlaNv9Km/Ru3TzBUhsOJeSDEJMJt1FpJIaAFvSzIVatW8PrE
D4+6OcFwTqEPcLUcYgxpM2tb4Y/NzTwISYAFkZInDo9RCrSTT9V8ytWRIkOFKuxPp40Z7B+hH14O
ulgPZlhAg5C7WKmcv0o81H25NJsMO0GF4vtSl/Zt+w3DZWFf6v/mZ/RI36/DsDk5+U0oMYPq9w59
s7Nw9OHxXay0kGQ26ewEnUT7H+/QdEONh5cGtnutvM/1p+mtVshxNguMOkBLqeQ6SKMoKNecewLH
9uew6IDTpQ8b5AZ+SwD59+yyws5uYMs0gDmHbPW3soUFYn7KjM32tDQ31v8odPWH1QT6frq6MW1c
aX+CzUTq715HJpc9zTnmWsNC3+++OlyoZZ+wNcI1d2PWaz8hpMl0QjRN3RXqmh/aBEwetPv2NOFy
gyWeRjGLLI9XmORi6niAAdw3ewRnG7EcXGO+GG39EaB4fQsRAfDrAFKKEQ7q3JVg38D94CiV6j7F
wY4ijJDCwZyzDTPi6ihD3WAb9A2jVtqR3fHEoGxWFWDD3ebXS45ILP/7adUNAV8RCKydU3iKt6/F
C7AykugHvHUhscbY7MJOA40kPoNn1/eqTNk9YD5Cwnzn81bq1lLspEpXpQPg7FSdraFYy2Mu3Pz6
cCLeZvBhcShLLudhe4sb+1EGJiJpvDvoYboYZUBG+W8EG1QZrmVwneLExUllSgmmQFN+t3kb7G1N
aAknL5lL7vWd3OJWFEPMSoUJJF6jCJuslWiGdAbI6wLavUR7XHhAdJ7lXOFf65ZL63iG75Lp/hli
REOrFZWJum/5PMyirJ421RD3ixAlQGa+EjpgBkw+60XR3/DDoq2pE+H8XjrrFo8dlgKL7hdZuALJ
PL4MkuMRdToq3ujftxYjB4o2Fnb8exuB63TkZCW9mBvROzLipIUymUO2SNq3WXgIsSmfDnKRCJWQ
OV3PdVlM+ByZa50QOBX4Q831WVfiif06SnAYB5QQxk76wXtXJCO3vh9fJZnYUGnqksuwyuwxeGUZ
SFyFplfnci1C9oGiDaAczQv4fwihgpdi9UNKCOLwEPfCN80oA7mPJy7XWAmjBr5lJzFBGfXR0SBt
QjAetcOlNSvDLWF2+lmKhHBAkBpL8KSUoTA4eOUf2tqaNKuwk8k2sz67yvmHME3zuyNux23VQl/C
OWRTi2Gxc6Zwh5pNkzHfWo1Id8JBZso1E16XK8gPXFydbOQapVqyYrjpPvyd3ZWDMuZdOfZntY+j
gSycOc86Pd0wx01dRAP1Lp8skTfWKv0ajZnzMHFcVI4Q4cicTuB0XrrVRVFe4Tvg7btBvk+3d1GF
Icgj1cVKbEN3saUl6x8al+ws0NQ2E7rssOZCQ+GeIho9XUDBTVajjhRVjBpbqb4Cmt0REBqpmOAP
8D5iecrEsFXg9CIQb6SiT09TuDC3kUqYVqKS4yNLULAO4JF7qIFHkc3wU1dNBLsRP/e2U+XbbMrS
UUwLG1a5b9/GbxJrulnSO1hQ8EygwARKDS+qRNB23UxH9Q+aENEroXn6j3T5RK38AeM8Ait99I/L
l3PvwdOpl7ZajQrCoTCe1dwcfOpzyUx18e0qOoBEvbKc6U/Gfyl84BrpxgYISqBXm+WQtjhq2bAx
zhb4GPpUJao8vbAlSU84+TMx1TqFADwu0+aVpTv/KQ2KDUm8XN0f7E8dl517yfbbCyUDpR59EY1t
vc3NbM4o00MCvu4arG7KQ92hwOHP2qQaIRR8lnZQk0tLwAQ6GhfUhtsxha5Z7Cmh9nDBilTvCff2
v/SJl0Iwb+6lA61oLjTl6Oi8qh9eGmJli4stuROZPBVWwZ7WXA5fYrQXt04BaUH3J7hwBX83FyTx
PAJmcuTKMUplww088J5mA77N0MUeZFGnl5t7CW6avS41zVPfDL8Xg6zAiYmv/QjZgEQa3zBBoNRB
4AmmFs23b60bTINPzqXVEk/A/MXldEeFiR9r851cIyxvps/48SE270QgxzSqSuw2eJKwWm49eAiT
vMhPJ0AGS63qr1yGmt3ZytGs/78WeusFK66NcQsiDRtTcNC6CkyMcCX9B7Xqwxsg83rAGDdXu2+C
SUKUATHEhghURIElPR+d1GjhwyYOZWeWneJIsC1oa696gD/YqR40fy2lNbwVNQuQ6xub0yIDSX5h
8OyBgxY9w2aqFxvNX2EIsgLdCzyJQgL7z5jaIfYg+0UG5gbZ+4CB/sk7YQqI1ircXF0RMI9mNh3q
oraNO3pB8CYzpGehuGUoMGFOXwcFJY4o/XF0Ml2oZ65Dufn5pbT3Bp4yigRcum25JhlYOP/tiF6d
wlEsZnsVcBPA2k2oK0MwWVLz1ZI/Y3s9E6Iyvxi1AF6kcwOJE3UR7gviyyYg2uAduKmWYFlQskIo
Y0LL6oqoO1HhJypFmvvIo49BzmB4FRxvZgGjBQwFDJLkLatt/F1mGsJHkwzmZx0/OCJ3RiX5IJ1N
CD/mCjEAuIHbOaCeQD1zzi/5fHuj5fkiu5ttvZhkgNwUnD+GPo9XtlUsWqvcLuRCsdJEVZ1r/BTL
GdQ7AL3g51Z3JfpHGv/U0WET1Uvpq0mwLBNiAF0ozQ5rQeKiVAYE/02MGVYinijLIKJsH17fkGMH
FDQcitz9a4sB8+5j69FPFknZuK21ytx9l6u+3IuOx5yqwW8V2QG3okh5YL4y9IdvOGq78k6a6uSx
LQcwqxGfBaZi9ZQtG+5UE5IZRcx6pq1kmGZWaespbEtKZcwm8xvi8g69DtW2sZvnuFtVHzSyXeh7
DBUVNSDKU+I+g/c4cm1yDfvmZykUvKa7fc0yhlFZ4I0CR6JUOKBAa+gbF/YWvUwvt4sHqAO9poek
nSkGRYTfZQPvJmNwEpjsVrCEqn4rgmZrgHSyzkztU2alW/u7IC80ea1qVcNfJ/oHM2hna+R73gDx
amumBEFhJAMoQibgCgQ85Ry0FTjV304VR//Eg7O5b4vNtnkbTZDr3l/Q3osqGL316F0LG7351MiX
4O+VGc8eI6NF5pi2Axfx+SAFVn+8kmuUZFSeq+q4icGRH2YHPpuCHVlYsoQV+AP0BX9NF6kCHpPU
FkR8JzQ8hMSmjrTnzEnECqYelD9yhq7fXuXKGy68Pedp5yNGIPKgWd4IF8U7t1X0jyNbzllMpEbY
N646pNRi0xIDEvvfecnpy1PuhEn5rQ2JZDlgqRN5Q262/NnD1XMEodhUutbbM6NdMy7goq+1lZ+G
G1bdDght/2FoASg7znDtgI0m2WHayFPS+KKbdwUOrsld5FvfxQBE078qt0ht7mZsGLAv9pTXi86w
lBmOhkqSjcWQsNUjzpe/4Cojn5iXSOLLCl3RUZiqwZ7J8NJt+XbPX2cln8MSoFnfTW9yR7ylC6tP
6idhOPARhDYitDgsi10nROPh14IQPj933atlw8TGTaQBbtwtXRiFpiFAugMnv2OXduBY9d7/jXPZ
VUiO3EdRGEZs39mKw8LKybSg5tl/quv0Y9lNCrZIbQvkO8CPqpga3Pk1YywcpBKGZ+bHja8MIOiz
m0L+oYq+TQfgLj/8A38zvQCf21fKxcINub2kQR9HpiuQIBeqz53rtDeXJNSCNvvxgBbufnrepj1v
dj776PKPD23a4EsgX1D0JT9HatWjmglcxWkYc4TgAA2SGoH+5g+wLNa5hzI8REwpTlva5BZO/BUJ
Cq7M8yWMug+Vh8g+7X4QszWf5tP2+LYBqGxiH/UGGMFvWFwRhyl/V/8zPXoEoAGdCMF7fypWn+u6
2EUZhXh2RZVOQUCStfxYp2+12/QAIgu/6B7I7C9VbaVKnVqQVDTm64hmO8kdhO2/M7gAwB7QTEjN
GqmO78DFnGTVgvpDSg62O8z/UxUsr1Smt2tkOGKUuYHUq3pjTMY5GDelFSWxKo508o7PU/3Nsc03
dqGGRcHp/kUfvok6BFeOagokO279Pjmiz2ASvP881KbYJfXQGTWIUsHTmcR7aiEqfUm3YAHhVUgq
mf2U27TRQsRJY3iB/zb1wIRDTYzKjjg/S+VKVYxhW9D7VId/hqEpJy9vZCQrBBpT9q0lSeUWSG6G
z2IsjxaspFbHy+AnvS1GbugnFiNQn5fOi3fmTw4XDmGy/VIWbt3uBn+LddDcVHX/acWy0Z+497vX
VoJ2K58KA1KNknVC7k+a7nyycyyFYOhGIFMsu/8Q7NTC2LsGKNjXe+2iWZEAFm8LywQyDaFXgZbq
VZtOypZW2DJmT9m42VOrVWVYLmWZ9YGVc3yffF2jLUzyw+yyR8VxCKlGCHpaZ6kJ5WyyWm4zxlsP
vdHuWChxTT+vYbxG/eI8C8s7mQ9UJ/easn6hSEUvHFmqzqr+vBjfyVkoubfGCB4jnpKciBt77QHb
UzxTQ8mSDwCzss4pWFOjzzhUqY6BviHYPsM9yAPfkFSz0KwCf5PR5ubs0bAcSE/rEWoZbhTLHKvp
TVxx+8RBtM6PUy/Xx535hJ4/yjmXpE0T2vg1mRPbAabDaWwG4lPYSv4Y3ZpwHxYEz1T6ie634rS0
qiMZ0RNn9VGCn38O0KZLq9OYYglKZcoDcqGb0zVZD3mVD+4kmdKA4EjfBC0QS8W7pH57Mgymj1nS
3aJjxefyAX07Ks4fDlQ92A0g/ggogfdm0f2Vl+a36GSSnlisU6r05/a3HvXXmy5QhdqFsNbF87eS
GDejw/dQMLqGMXGAoxrmtkdTCW0vVNa5G92k2KI4rzbNo5kptssinVZ/hxkaMoynE/lHz2kdV2j/
59TP4d2EdkgVC50e9ODj4qNHeDvbyLP7B38FMmMdj+a4Uvl46r3/2Iz1EJ9T/x+7xUD5g8UlcOWL
6E0/Z2IU90g/yQUQps1ollqBAaQLVfS3LD2n0p5nSRYX+ybeMKuxYlFS5PnChOutByCnls4alvC7
7qHlbkIgu/di21IDQ2vrZYCggf1oY8clBvQvtGzWci1JriiTWCKDIqby2+I/p8zhYglVVU7shHYc
rHEURpNLM5w4zW/jt2iMVRFb58N9yc6IX20AcB9HhYMjqFy/Q3wPLds37/9KQ+Tpg4jkpNTfqx1Y
4Ci7gkOgrjzbF2ncPsHuHpx5BqmmD6jblPAUDhlmUoev5ghDDAn0UuMIITJhOeh2w/6kLkhg4IVw
FnwwC3x37BzmiWyvh8Olp6h0KcH5sgF9Mih6A8UuQXM0YRnrohig2QybpJ86Y7JjhNDPCbILab8U
0P7Si9xhla76RQf1yPdjkfDWxObsY+Pkq/iKIc+LLald1iEz0Sy47SLzSo0B9K+x7NewPAMt5PQh
pM7j/bPO/UtKIiNhUDHbtyIer70hWSkQWR1xBPWPnLMvxe9/nnve155uF2qNzwHrWoAuc3PTwInM
5K2dYyy1x9TtkOrnJvqk32vneJ2GF5uaf6y0HjPDPUWYFj4VcHYS4d8CcAzG2uibuJBh5Ex03rhu
wDB1cHJ44L5ECrEv4Fp3kYOgr1+Zrnjl93v8gUjHn/78M9OuI8hWJCYEXQATEcOtj0ZDgBegcyxr
4GYqNs2UJ/UiZE5cVxOtyTXH36NTTQvb5gS64PnspPW6fJTWbgMnzOk8stTF1Ekwmmqq0ouKojso
MbtnwTvRZZkskPb/aKBpx4SVO4E1xKpePe1d+1kde7J+qMMkYsW21zwyQkgG9+28XMsDpov/Y/vI
/rWH4EKcxuDZzJtiEI3q19RCMnLySCPACd1+XcONwkn9ffvvpfTTg8psbunwDlpXZNn8xYiRFiEv
cSxMnZexc6mklVRmGobc4GqIyhnaOVLSkWRAEWxgGDQ85Wi7GIT/cqqMRtG9aCpW0gBRoqo5aXQA
g8R/fDZjyZ0R7+F3qaVtAOehzNZ+oFysDz/oI7OC8aVRmvIdX1W06xTFmDl/HKyXPN1j/tHNY4PU
P6NM5b2XsNVbgExqYzyH/hgPvYRrrgXkITog7LkE5WIfOkpvACF0tqNPwbxRNemsBF3aRb28/98d
zTs1y682VAadGfdXlGAv/T+cDS5s8Rex87FdyHkvg585Y7SuyyFaah4Gftfx1pDfQ/JvoyiWu4a+
uJiL1GWIkZfBSroIK2Ayymkt6ZcWNBCRcuREga5qo0i/X6rY5m0AhA+x7cgfcL60/Kr/yif/7zuV
RSKYpGAuFfyVfhJTQ6ZDcU/tVbkPhvKqeunCahbnkcQlfdm2Dm6Tai/LUXCbwKHj7pOOsAh05S3D
ejCTUq+wXg+zhUq4GzYPYNiT+kqLrKoqTjifM0WEtlvPukByYva81g70uHoTevhUhDwsLE5hVg59
9gDmWk/EcDpVPotKocZgBJwIR3QLgE3HH7V7gqArFlPJHoFPsK9rN0CQYLuuJvPHwZarY/b3z+JA
Rm732L7RoRWzCRaBCEyqoIzIGZHtPBOnP3sv8waZ0q9v42GXb8AX+TcA/JNtAabnlcinCA/HeyF0
ghPYOgB3FUE2ZBtIAiVfksS8wAtfup4+rmE6tC549NRmZf002RRH+cJfI0rXxE8wGhMxRV87ClhJ
m0+ZvkwQocPRnKEeiBGfp27D4NoX7jq28dC5+980e+8hEww2rA8uM1zvXJsVn0PpD1nvVjXQWWT8
/GIXHTCwnxgnaMiOR44+zod8fVuqTaaU7QO8OaDueBVIEv+J01l/dIeY3iO6uRZeTlA/6c+y2Wa8
RU1HyGouRZSJ2h4HqbsDtDY46fFXBszIKUBtBDJcW8eg/MSZWPMYnj/9WbIfoWwnlxdBnSz2bJI4
Aqm2lxN0HRJPk63GHTcjjF0qk0PiKebkydNiB9zWui8gBh6oLRYh1ABcjzpTcnlrfwcnUWAjXUAQ
/ZlKKvP4GSity72mm5LNFZ2VipikFwIqQoTtkBxqKXGlSa042wnzKHZgL4XA1MV5IAaRVBsvxMFK
Pip2TRw5ryk/kENmQcHn6Ngnl1BtmkwDJmKw3alYQD76lEerJbHVuJRFIzGXm8tYJhSfsQPQDByc
xn6JC20Jno28dhakDTp8UHieSUaM1fwo9NjUwePb7zQUHX6j9VZY++GYUYRHSYbtxmrsuptohgCZ
jmCE0/C6CP+YrLLsDEfxCJIxVxPEeZnBLTkXYfbtDkQzCpPu5XpqrRGjZmNk8svdxE72XVNmt8oQ
Q/7N9buhTnuqDcFih9WOBlKP4ZlrToyjljS8j+XFItZoKpqEAqkzZmWRMRP7bY81Edq2YJP8p0Kv
03KyfkDlge/zAACyHo9K3kcADCSVOBKXa+tMv1Vyaa3S17JTI0pglq3o/cgsG2fYjo8toU2wHTtR
ChWs4QJnU8CInKkawA3LRJLABLPBJXj9JxCATqfAaDMPiEPeft6aa32hWVsgJk02pL1c5LMzGygH
fUGnl/USGk7TJXxgsvxrpRxzP8rNPnuAzc2Q++tZKqT3CMpGsC6DNtOfrPcwLLgzcftz1c47/vte
ZejqckYgjoFME0Nnfjs0CT1Zh3n+n4xdz2lVj39lfHDikzXxngAzcTIuCinN/wJMyvvKcJrlRLDN
eL3TBMD+0ItXu/Spj/NE/s89Dmu8wXplmqiv75VH2taTgXL9zwk2v02BL/7+WMzYubgyc3WbBwFd
/JoZUMkTZoReUI3NA+S+VA+lgGBLlSSlObUmyA2RpIqB63tn4GhURFPM7htu+CEJZg4MyqY6ivEJ
KNSr5IKDepf3I0jPUZXwyINXbWYUAUANNz6KSYKd6J2LQ95ge7n+mNLuWe66mGWLrJTYr8GQaRrB
AC1jzVTW1NpR4RtLR1DhYttyQ+wYIqG1ZPeJkTxSBUVWpJKG7l5zAstMXzsSLzFBMzt4YxIZ6ZYn
bAzXYp/aqT9VrVDGqfTqptlKHd+ch4qBpXSQfb2R3BEMmNtXv8laTeWmUCenCxjx3if/DKsRMpxx
RGVKVnD2c6KVhr7PresxdaF8JBtm1uIo10c1FTzQ1HebZ5EixcqV2Gv9oDwL/AFsEOFFPNjWS7C1
NpSifrSQmqbFZRUcBLkKd963U3c84kEGBsBuMhKHSuO1lGvMmbKpR3+QpreXCF3uKgFwDZraCB80
kqwSGSznET2Rk1uUECtqetAs2EPHs2Vq1stXLulneb/84nJBB8tY7hVdA51xjBm2tNPtYaTynesl
LRVbO+fSvgHIws4fQdqa72ZBYo6FvXf/iV8uso0+cU9kcmBMGdQG37/57tyIs5HMH7huEKEr1EO3
oHOmmbftqwaeYip/PKBFB5xbSovmaOKh5rtWusaF8QPsUX+gLDtL0nCIyX5nBYFQfb9vVXLslE2I
nW+akZ3zCBUWRh0iRrlownuNOH3x3+d6oYhkSPUgx5HNDIP3xQJj29DYwLPMmfzllpBWZO3ouSmo
KML1VPP0QNWxgKZOx2XRFy1K3Fv+w1wg0cONY2bsVq+DTTSCocZTQyaQcqgZOzHim8PFMPVBN2Fq
XPtIQK0CkCkdVpVJrKGhJY2bJDPX+qRWBtTsLDCYoe+4ETP0PVUdvRcEDfMNLn+u5Gq7Wsvo7tIp
yW59qmZtgRqdmsxzcwoQOdBbOj4COwMZrzGAwzZgdQG5zUnFf7O2YlgdN055gBJ4QpBkkGzZnwWD
LPLcjimnqhGd+uYbUX6PPRMYkshMJL/A0NOtF3fAcibHURDZb2dvQX6d18PKk5RUWIbrk8OmfBzp
HABpkS/YLlnusxVMDYgt8Aqcl1v1W4xffVOimii7OOFadPHEnEImvORhwTcsty71Zfc3QTeINtmc
hN04iryO8E/9erNYScC/fl66zpWsyR0PnhQczByydEHBd6P6RP2+6xvDHYAydTTkey3FalhNhF7M
sX3Zxtg6Iz+CGOaoTm4Z5xu+Oo8q6I3eR81fLSYLj86spm7k2sVkMaNGxpVkce2p0sXM2W+DF/Uh
h5Aq6v2wwSr73DoSvzxVuohD9XHJRo9Cnu+/3YkU8HXozG/8aOM86MEJw2s3RsgEhTQC9z86cbp/
RC766FlMV+5AIFl9B2Daq0AqCja1WldLb6TxK4hfdyIBmyH/VhhYVnJfs1zVp7mTMlTleB0IFcI4
8Iul+XGrYChx/DsakSFw12wVNK1sdFpVCu3q23kKDKErmtY9hJyFTKm+WqaJAkJ5jhp44vdz/a1i
X5CujPvespuNxhGLtsTb52iYTvzO222/ZwQn+oyt6j9A8yvVgz1BV8pL55omI5sDNtUG7/48vKCZ
aOAodC8u98fYe78G5wf4WZMzd3SFMade+t0F1ko7IfK/iA4RF9cK5Zt9sM7ZtqLZOO08PLPA3uKY
f7PgqOjx6EmA3jGvmEaVx6EsLD6ZhK0m8oaXFgp5st86CAgMuGrXQWTvZZG/THEedTD8iJDl7fg9
eAmUTPqbs6eBNKI1E/Xc3GNHUXzwIm9EbGKgUtZfVLPyrJliFhuTzuGRNJGS2E9fhvGm9Y0rxl1N
abL1msuKH5FTreRWR2ixnr4FB/5hfmUICLAlWrsp+sgXThlXTMgxonmKxzok/W0KHSHaMTHEtzTm
+JGam76iqDeHpDaJ3tntWbxDGgptCJKj+lr1ii51pbd1Tg9mOtSn+n9zWxeyFJ+tokEKgqLsa/2B
NvJy8caAWPVCJ3d7KhMwJTWvYJAZW44fsxoWq2hmqeGbwApjfzy2X4o3G3mdfMqrruAss9yPIZmo
kAUK8HZyS0fNCcAOEzjUwCkeSgnSRM/ubvP5bcOGQ2oP0BDauTkuTqMcokY7TplTqmK+mu8ou260
P9IwL1W88hQzE0YjFJGkKHkDTfnF57BCeEnU35W+HhhvWPoZ8wRZqSCXRgOFLrhOYZNRoyjgA7UL
HsUp5IY6i4EiwvMNOwP3l6eoR76NaUQXjMJeywiB7BG0zVsBfHST+PBRMFrLb9M1q7lT2jOlfOpo
9IU8G+Le2nZJPlUu4kqVceBVyl/hAWHKhFi/2T++1+yzpHfKpXERvwcZUD+DknJU0ejuQjk9zhTm
WPcWcloPZwwjDniYBwRPXzh4NpX9t1pYOay4sa8BcZ2enOuvc7SETW/SAYPtPi90Q7p/FbW6lP3j
oPSMm2stFZf7EoZdBixKE3/6AbM22XsL0ESkcao7QF29T0ICiTAqL5S9Z1IVjHTlaAaaVFI1Kqoi
oyP1jYkhk/qLMYxR2riVDF3GuNADxAgW/Aa0F/uzCwch56PKZZUKahydT51n/Ri0vQcMTsVIoUxG
ZjNp9kA93/HYX4hsQQzp+66pQJfs4ZYo7wA15JHw3HMkJ9V2Agg4nG0T6zXPV494W8xdOnjDl5GE
9FDyrPsVJfXie49pcaZ0+J8WTZzOBK2ngkaZVwPNXeejl5UEZex3emuftXNEGO6FoQwOCqJ2Zsfq
4clANM8OF4RHUwtF/Akd5bR5W7qQAlUzNaAbyWOE0HtfacBiPVIeWr//TOBbol1rQCusisT28fI0
qk8BRTe4ivHosHH+xGh3InkNYWp6x0xprIL5vxgBDVSfX7moVYBfeFYa0qMi/71Gfr0DMLeQlAwa
HVlT/UGF6VJMwrTc+X8Wg+bZE4Xvo2BwiuK0Nnvy+fqK4NSnN/9wQxKTNTtDfmiYJ+oFFmg+F/PU
pdxeR2pm6JPzxE+nVze2S71CWdWw0q8I3vLQz+ZwEMuJQRB12Qa0BJxnxOk+kXbvOtb7AdtBqW7p
m02oMM/MgbZzcEQbyQVoq/th5Vv0o08rAEC5TXOUXpLN2Ld1zplXQFfTun36MZA3PWUhCfaUKiek
zulGyl7EBjrJMmsSyzHKXWMDZIQoxWSt1hPQX4wl0ARhh/sCcjD+T5v793lnwtNU94MvS5CzxmJm
SOwgDBJsjGIpLi57FohdvKlZMZbAvL92atC+ErT33/HcEeGkUg6h8L+B6aGRWoZA/AuwrDShTOxc
NRyrR7ZzXfEGBnpfmDZu933KwOPgqwE6ZGdKFvgF4PDTenpw6EYzxZd6/Nv047Yn33chHc/WNYdN
IFrWEkr/FIKQOf9YFZXG7SqZ4bn8cysk9Z7yWd7eTqfJ0kB/AJBVyuWGydkXeDlJKdvxtv7hZzp1
xDIxN5+Pt12H/O6cYt1Yx5AbmfU1pYlA8PC6T1j9ycpcM+Gi/xDweh4f+nEDhsDSjqG5iD7OVQ1Y
lZDtv54TvC1Bfvm4gPqIyKLI0+bln+57uibIpBLBu7UFukceI9apSIbfx/KmfW9omvc41d90j82I
6HHxdR9o7+oiV0D11IdDPSGWlS6S4DkArIo+KyHnN5X2fHjEfiFD2cr14y1Pq+nx61kk/eKm+2nP
KMTzgDF7zynzqJFpCVcQfRorkMq5b0c4hPDgEswHfttuUqNyRTftaYuVHCYnCgvfnbOwSHxH6Y0p
z9XJ7Z6QPvpCiHOPPX2Ag30pS/NH1mUHmKpNuj4Fqvbbec8ZiiN+XVObSLdTZGMKyHSu17pMdfkO
Q6s4Ozg4pAL8vupJe9exbPEMmVrSEOyPBBvBAy8Cp6l/hcvP+BFtWfIpGHZ37uhN53Zt+ZBFGlzy
dqhmNddJtmQit4uzf5X4NK8pM0KRrrhvxAHQNXLBQ2Jl0QbDHVKe8mfGwdhrwO6doC+39EkmX1D/
iZwZIS6a/qp4glcfYPEJ/65yL9C5j1j1g3+ctfnfZ5/HqKDL5zw6GPnE4poUKGxtRfLQGZp98sx+
QQBD7pPFZSD7qsb7EQ576VGJ9s9f18gA8tgUW40T/BI3K8FWDPCM7oF/SnLlMxw9aFKen8oauRbx
J4tqPNmsoku6tk1qewJWc9lOkumyJzJWZp5Coa6u92tUiGfhwrLeu/riX7a2xkF21jsWEbmeAv1D
I2EHRP3PxWyjcHlDmZywunPzr6DgJknQ6fjc4YJIP8J4tDMfv0q0L3qkOi9sbPdcBlE1JeNRlrQx
m4T7R1n2Xn59lYsY1DZw3vQQPatU3pzATU/da5y2jMxCrc9yeoDTfjA7wXd2p7rtT16sC/NSovJN
2UizQc9OHsd4ZPzP72SRMFePBx/zrYsOadE+BBKHizaxOPreQ+al4Me8KiDgmBC1E6J1+lCwTOp2
RQomNU7LParygX8WRx3eGmT2fFvgMe5BcLzX/nCDjvcRGAuP7CUnTVdo+BMPIWXgfuTZn2C+bwRn
2nQ4EkGPnHaz+Mg4sRwHFzzj4Umfgqu6j+gTAk3tle+qDC3YSmWePi8KsfjV8xp11aIK71AUsLc8
oND9yICR4yfNr3ai8P2y7sSM4kgm6mw5jxRARsXiy6+ssbfkhLkBmPcs8SovLrIUjMntEG0pvhKb
1ZGp2hK5ZlRfnDITr3oSflX3s7LzoT6aGN8zLPY4c/i/I6uRLTmDDiDYrfvwRho5x7eObyTGkkbT
5+hY+N+qsfvXW2OJdv6RaaJOO8Jv9oZxlmQoFlzAA/Um0Ad352gjCUlyOa/GBGh5l4IsfnmJEmrU
lbLAtqC+jA998H/9ZzPqw0y/vmd5fCFdzlXbdsqsKtIS2eaCHJUqWJ6THTcduCD0OYiFILTfysBk
BEDl4Kx1rQZt8grYBFbJQvTxyW0gWufH9XRfdih8YbJ7xZ6ZF9hxIeKN2YAi5Zsh4vGjeFe7uwYK
dp9hxXcG5gocLgn0JU9akcicPKT4RKZrJreHPEfUmigSceKBcVG7IcMGQcwz4gfHIQADlFyveoPy
0EA8+xJbuWKi1FSN9utpYENhJT4MjbgEwYp2o1NrTmv5J0pr0OFfs8AhK+nhetFx/H9n1ScSaTbI
xOGQ/MOnNWl7IlvAcSuIbotkkaItHm82F77BdKxuZL1ZCzuvZEK0fshHQGS7lE8oR2H7Y/4LYVUW
aYydoLW/IFD87ItRDNrT6+cEtrwLMIIZDapy5xgL4tkCHMd8dVG6gvN1MqxpyepT/3MA5Oy+TX61
wKTAtXclrb3c7zIMEzrLd5mAG5OsLMhh12j1xEYW45yOnodXWdSSFhIupOb1702oPNdo7cnj/85o
IPfapXZ5pUhCpDz6wlZ+f6AY6qbgS1J4fKnlpIOeaVvN8TiYH/OC7IawAsZLPTF+2K7cjedkeG5a
tamj/aLxXFkcYLEKgXg78s127IoU1nVlJWV/2KafWgbohFNfXcPNY87kKaPzmWluEeCQTLGmwKHn
0FC8EY0gGu3zWWDaagOV9mOoSdovrt4hgDgLbjBINVBd9kKUtGUCNjBtXhs4958sCOOUJG4gsF9f
edtyweYyFxEnaLmBd5SgcHl+339S1Du9Iqk79BG3gpz49DG0W/9d3hegilCIcOxpdA+uZnCHu31y
RpNeCiU6eyMkzQS32SUeD4EGUxCfalotd66bt/A4ZK3UFPdIZKbSmFuetyDYsGN/YDXNAtE01uSy
4h+0+VN3bAdwmAEiXEnzeZvcIpbKxm9BWfHgcWvg92QZ/3eKjoBj4ZSbLMUqp8As3YUCQAXIY590
axlvSgq8YmgLpQWl/hqwdtRGCigK4eo3ARTBMAlQYed0FIxjQWU7Co+JDUTNpsIw8UegRPjIr+rD
PUz54xfKmKbMzQd6INdzuLa7oUvR5tI3fJ4KFqjsjr/gv4Mr6YU/QO67XI4UEX1/CNNMfl0o8/gz
lt4M4uPFaw46bbOpzUtU1Y5nCNAdGCvgD4eyQjw4SOWIvLakmxBRBpkhG1dahIkTCjcIa9kN+Jo7
yTg2iOB4wIkbNAGJY1du1BSBT6ONNjKSQFSs0JCTvCfWhBYuHk2VQRARrzT9bOtmeB+YpZ7tZ8LA
/DCHkU66Wkv98v4l46gtvMFynPJ0HeZWnlfq6mo0YvAh0yfnbA28Dm8bQSuHtAXWDh7wBSPhhSlc
Nnj2MGKqn+6JQyM97tDmMg3DGusKcY66mp/93FHYIyzdamd13ujQ1ogMnspDhxhcADiTFX6KzJcb
oJ5C6NfQSqqy+qFbbt7dlZ87OZZb0SajPonRCOyVOUitoWZJLJ8CVpciW3QIH1yRCQLZp9ZMybds
22qvBl9VotokkfzHQAX5+2CE1veksAsEoqgodp5xa6EghLSzlx4P7YHUVCBY5z1/bx3RTq8ikrBl
G/9a7Ai9NRnDRs7f8ibAoj1pkJcT/fg+3Uksz212CqQr8Ww6K8Qp/rrQ9WLDunzT14yAuvdt4yGk
CAUu8os26/fybNVQU9zMb/cns2iHgdj4An8gsyPgwETyD5kkymvsyK9CvCAZVJ0K3jqzaHvKQsvV
lgpTHf/GH5pf+LimyZ6a5WiwCvMPYq0/LbEKqeZ9+VnUOjXRpDqkIcOle7cdwYrbnpG4lju/8TGA
Ovmy+fm0UDAIJWk2j3rrmkm7y5AFdRUqhZ9yyX5wu1NSV9owS4zSsWeyNm9HuxC5MKeFoBPR/z8x
EyT1N3K5aUAsXgi+MedFSa+FDcuzux4O61CzP1RCDNWEZieZkvYlKWzfDgeQN+Tw5zXuf4hDYVlg
Ba5CCrX2GsXBkPbmuT3P4JkoborEyjyIbLPq42U+Y0uFQ0hoOkRBtpwsys9FD1fsRk2aIYKj7SzG
cwyID0rHrrvrRcxyj65J6E4FY0q23/hTt4Pw7rALpR2MDT9M903vf6/nMtSJ0OQo8OXkBZc7Psk9
xNI2gBvoxi2nAMvVGiwx9LtFDP58jOmVWsG6/prJcH3Sdl86LwXL840OfFDze67JM8ZywsJI4LT/
U7gfJ6D/JJ0amxkYtYfJTb0XhvgOUIcovX3JWAPkIRIKYuyG/VhfZVbY2WZ6iOT72iorrhOlmzpF
9Hc3cuSKILOOyEtq09OKtrFhM+cfKv+Nb5AbznWVfhjnlJibwmbWXAyznD2Cg/VU5JVif1hkvO4I
/DEbpGVGCj7YTLIY0PRnl7QRVbFJaTxRiA5ohPQtWQgTqf4Iq06I3Lja2GCxywJs6OQ04zUccUlx
mxHE1Eam2jbkY1n7aBpMKepGlStJ95Se1pf2yByz9qRfy27Gt85ZOOuv+c9dQTKcllyomXlozfCV
6frXXy3YBRehFdRq+pTugo0NHPySG5zxmaE3HlA8A2kHL/DERZmUkyR9ogEywp0D/XiVTaMgGF12
DApjeVGXlfCHRvQhloeuzjHh2N9Bm3qA18MyjqlHzIQqzYScklyZ75aenO53ooGvAe/vh3bX6G0M
bBfsj/JpYuRqvsVEaV4+DgU0so73yvkGmTdBiKp9sCgZJvfJBx6bCRZI+vdnAl1bDaM8SvN/kpQ6
7o7KJKf5uODvjf/XEj2U0CB5v2GUzqXLjt5QaRaYA6lF8LPIKWOdICWI8FMTFyNIkE3zNjOlQvDx
48tfGmb/oi1PuY/bUn9rloCJ20XTodipkW6ot47oINRlZe7aq8SZyOHHIXRjNEkCuQvgwwDkg8oQ
95F56TanKr5QVW2zUaBG+JuDrsjUeCdzh3uRudo5m7PYjdDrYmm63DtjSuwnCfSlkqYCK92VBTuV
Oh70Me4gIoZyGo5sQW5PF/zKCCw/+WC/UPMGFTTDlLuSJsf4p3VO+myHX25ha4KBH0XM4nSiQFjf
7VxuWu0MBtUp1ixg9/HVJJSyobqL2OfJnxirQOuIVMUyiDFCMB7NF5pMLhU1v8E35jDN6B57MaQL
/sR4dvOkDT3RleK9MXZFR07RZz/eATV88WSlNareXFANkD0gQybUm4eEDkOkJYtyLBON4oSXlz9v
2TNlPAY8aCRXaluYuTXqydiVAKkwbjIfWFgjtR+xwEwNa24DIeJbcQQ0Reuj8NzqwrqvnSJslurK
uB9NUUET+0UetUqaIPwjIpEwnG4WDCfKENjZpZ4gA8iumGq+kCADEko65ezcVh3b0wcS+cEWjZFy
SzFto1yWcL+dVuK9MlGdG1LsPiPEA/dDT98wL/KUX4rGzal1NZal9wpn7W+j8gqW5hdpN4YYbxVs
+vg85PQhCn0lTGSVngzKg8qB8y/3iYlBoogGxElVZ6VtwhTbFQZiJPfApjJziAOf2tLAalLHI22G
su+J0xHfmCklwYEp60krK66Dv2zUDSisVHWwCg/KMxTqsvGnKKSHsgDuB0MSBovre1lYpf8x0yvN
IuyU64tXczOT3X78RyZkoceaFggavZ5+TtLq4E/MHvzmcjznIicZilPvOfp2NFOMgtsYcSe2/UYy
2yUPvPKZxNlG1dC+qi4jSN010Y4GX3Gz+mZXn1JwZLkpHSEd9QyXA3abxm7ReIpj+tgiUkBMKLCC
p0CWxB2enNNsHUJovTuoNx3O/0xIH/dAWuTQ4WzBTcwRs0WXDoT8aZj7Jn9puOUyZuz0OoaWT6RO
BZPmKH4bxJW7+35HXSncnPRWQe3v0p/Gra1XlmpGIzHatZzo4yJqeb8BQHyd3f3WZd3ZLT1o67x2
YI6wuZT+8USiWDfaZo7jbxxYOoFy+td8aFTX6PATK5Ab/QoU8oo06J93g0L6pwXOHk5XGIZx6Gl5
9/zU/jVRe7tLrd4BFj4Jwt10hFzinInlhyRtZacwKwzza8G3jGUzo2suKxMXwBXn5UgoYcVtDs4c
zUJeAdI5fLdv01NC1IiQ4sKb74UZND8SYKVWIebJdr7ge2PYzMueKoSNKS6JrGRvx8m4SzZ26Y/B
W3khUTSqSrbkfI6/OYJUed4Ebp2dvpkZyVDSyLjZSWWdb/RF3NkPxI4p99SFtkX2ypQaKJT0vUwW
h8HNjOK2kuwCKTfAGZdyQaip+tGC5Y6Q2zORZRJQyLPVT6gRG2f3rZu7Obz8OHQMuqfSAyQyqFw9
jNw0/ysfBoxCLjKkhiADrKZZ/RXSwkPj0lyPCmwXUr++BY3xkntuNO8ah11N49Ul2pifhOQw7VfO
cm3Q7Lk+Ocj4erJDZo5ATReAvykeHjHBO6naf13HG+4t2i6MEwpwMvrWpoSqFHGLAYCwjKarTvB1
K3ZiJDHx3eBhH4MM9OmHFPgb+Hc7kxNzDkVGfLUNp2sgpedoQhxbfZF/eePrDgb4EPPoR7eGmnV2
sVYE1wkimrDx9jHAl4iF/xlJgSlRDpTITRNc+sLJO7p13XHMmz7CHcQskBpzLMwjLy/eG6HBfdBQ
tZfIdIEO6fl9tdxnoyrlLFZbiJkQEruoraNI0LKUJeNodTY/dmA/Vc8jK2Kr2/P/OoFKcp1CdQdu
US+U1D6hHbNSAJS1MF4sZ2BfuqCxaWCHIjwXVOBRz7oKi3oF1zpEnlF7AF65srCSqvQOH1OFcCjc
VFgGeOnRvbZqLJFJj21PwDDvr+FViiGMw+ACa9JbseJd3yBcmF90iJ4tv08XXPyTRzI3TGIQAGzP
VoU0/dtUJkKCzvcckNLRqpbSYYu1d5uFISRjhnlh5SIn18xfjDj53rbY4qbAlGM3pLN5ztIoKO7m
Of8nYTJZzfXDAeoG36slCGgVxsO2dYWVKBX9UsGLcR6K2YMLdZk118ChEZkXSGH5mh+n/EeG2xmy
aRlhkIghooWKWyJKxb+Fxw37ooTAeDm4mC5gmgPwmdDCwkM8UZUDy6KAEuwwz3ufzqAUZAiFjPtC
b5SylS4nDZHK5i17xNmlWzdzaCX+qFrmtTyujzQRndq05rDD70q/O7tZxjWdzaXAufCHObdJA6i/
IIqQv7xOExcMletly9K0ZMFif0LyK1DW3NUtLcUbqFnK8LuGhJWo4XEGym1FwweEEiRGv2qUSVZM
38XKXg1f0jvehwJHGO/qEOHlVeUgegsXsEHTrACFfV36mwfkBsJWRFTAlFIuy7n0nKSSpI3+aIrC
w3fXLOLB/LiCvj5w0I12sfuVAGn7wlcpUoXOpqI2ZffCeRvjt8ojQBoluQoWS1E54K53KqQm1j77
tL6+kU0islTS5DY0i6xMIo4weQxZGnBkvElSjQ3EVhJVwj09etHuVbfNxTQdR3fCeWVBYYHwd/TN
kbk34y2pEMXvYzHxZAosXGLSIaYCKBsp7lXFBtNh2TbykQdzw+Wpi6/RwWfNcUb7qCK6ytT9z8d6
T4MxFg72k1TT92Ba2yQGNjPTG8DNMsxzdON3K91f7UMUiZ6g2zZN+xmkESIoXHf1MlQZshYL42mO
68ujUYoALviqh+5v8IKVIiipIr/f209NmkezoHciaFnRXbNzYPEFT0BzK/n+kRebxPRHMkt7YZQY
4L7SKCV0jZyunJQIKEC6FnZ+Y1/GVNwS6cTdsRk2E6ahCXKlnr89GB29o6XTmRRUewGgwWeIPfIm
gSlKYWEg/pxsaF9HoBlFFdKLWRqsAxXzW2LmTiIVUghprGwR95YNQbcLX7zFXBGPRwz3T3JJyaCs
Wf8HHso4Evgd52nZtLH/C4pZcJ4uI5BHXVfnUE3yk0rOvXb0XMlHQRToCHSgGnd8bau2RAloPPAS
L9jMl/QHqRYsqkBM3+KEcZh1PEOMFKn/JqT1a/sRzwzl7F8PHY2zGVHxixnA7elHMCjcOs95YzaX
AviGDu9FxVpEz7SKl1+h8+IPDI0MxdgFYB4URI6wx1ESWdbJkB4K6s3pVElQn7l0vvoYOWbrvZPq
AaYjr3F57OMlGnp5Dqlhlc3fOP5aRGFeINTVueGS6HTYepSKytzPW0aX9nxHDxh4S7+PbRwGQTb/
dldhiR2YZAiwHYbCUbfKCWlt1SV9lJgVV7suBVWXrjP9S55zpKYRaCC5+l34+FTKfcUxWb0dE9sc
MCQsy6c/WPAHUUMOdinKXSqIus/Ix3YQRMWAT8Fn1Xh7W8NfLgZKV1SHst2L2NdDiPEW9X8y5sXj
ZAJ9hxuAEofbYpzcOiRq0gliQDq2EuCFGFfMQGUT+LJAtEeyYKhOmvoOCkWjTr1UWSUyIW7NN/VH
h5kNPUcqQE7vwe61z+eMipi5SNsrqJMSXn9kDr2jtsF3uLXi9fKCGLWADDFLX+KDoGFtck/Juy+u
Us4q7d1v6SByapLE80HlPhFOkwH+uTXpc3M0unF5LQKTi8oKT7Z5G1I1+GvMB3WcTE7e60rclWqg
AYLbKTIbz+CWv951N9lC30l92VAujAN3536atEHRVNcl01BZdoE/A6F6p3PybrjdF2LS5oK9imBt
lAcMw7+/8X9hzrgjbK/tbICMniyrQb4hTIo52iniH/cNaui1YMT3x9Z0pOvsJLBUHY1SKDZ0ivN9
9a0Qis6vZ5qLFwTXNd/peAzO3bfj6NESUcHMTwzKnmZcN81ifcELuIUfRFN5rATTUphlS8dlYNvz
zFuDxo9io0W35c9mkXhy4RTuXECxT0yhuKFYfgbA/T9UTdt5BaZf8uVlh2oOeJtwtWE349OykYNp
3/SiPgMHOoJ/CVx77n63Dtm1Nvq9+kURgq2FkLTYanbhsWhbTJMPoJtOnAiEWeJJSe/J+pED3DVR
OSH4X7jRxsoz8pVAWClpvsnkPQ8wnhT8VV00jORCnTl2n4VRvIczD18af28MApXcUydXa5yJ5s8z
9VbPQ68y6J0j8EDodIIWTD9SMSxV/KVA0tXn244uR2JkfncwI+0Zms1BXtSOwHc5u8gYajZQLHHs
QlTJzYN1VBGMrqwENcvk11Fu78X07Bv3n+ACskNC6NhLXpB8hVrRHINlRg8J8WctIruuLhFu29g/
U8dUHo3Sqbl1DbRKMN8Ek2i5vDNbbY6p7yL4SKW6A3LYVqeLNO5WLhSsJ6iSM8mJYGKjusBT4+2L
zbzFKx9egAifweFF71/Pi8Q6eppnYV0eWO5hebga9MOR9kpIoJvNk8V1Bs4aypof3HGJXQNaQvzU
TGjr/9DhAaAuDbVrvHoX52wt8p8iI5fL/zXKXn8acx2+vQGxkac8QLvEhMaVQuy6bm6hrDsjSITq
0tJVlR5w1DXku7Xoacr8M0X/hdOlOFBFYCb2wYFD0i87XzMqIOue2r3yXgJRsODYVdshPDS1WeT6
KTUB7C5SUO2Mgoj9udZvCTuofDiGUZkGWD2Y0AQ9sg6YULXjNasq1klm3hWGlkN7LFqfbH7T0iFI
u8k6Dd6H2zCtd5EvHRYNS0IDn3Fp3JLOW64nFbjrFoozoFLvaNp7io9fG6alK0o99YAouBHIeENy
PuYvTlJtERM8fD/I5axo1fTGssLjChFQ40Ca7q4QDfvz1DQYfy28TDSqg408hqsVmOdKVhUIqNIS
0KVCdDo1oskUX7GuVYKNgYP2/Y1ZIkPkcJTUfWTUGJ36wDzXwmKe/JzUFEWY6drVqa1YZM3HkEFH
Nmnl9TUmTZ4a01U2wDJ+UBqns8PHGL7gvUqjKPLom6+Cw7oRw3QM6JGwbnDcEaYp8k9Tk6uJEwi/
foenHMCxeVbzmfcfQxXNUalQ/bCb997FSlpuzh1z8M13HNlxwnfXGAj75UItaakzrHqIiSERZoAF
z7+mqcXVSHOTWZswJqxz/vjtanYijdklU7/995gRO8uYNlXAaQx7gpVzFSuyYHr106QypdJNY35Q
ybSttTHrDKvVHJCQBSUUupRY1I+FSVgfkiH48VhHEqYhnF2gmtT0KY/wPjHpYb13ycbwtWTi1T2a
zrlBkTz80cPgbrRDVBBzu4dBvlJin7OcGCfYpe0V5OdR042009/EuehxZGyD/5w2IlPHfKClgmdt
Zum/77P879L4gftAMWV/T3iP5Gd4oH/BRrgulWN7RurVo1s15eoI2hz+2iLiX1uCPPBCJAgHkqa1
5mMDQUtdUvZPMwdy21rJ8N7ahE3dRU6q/eVQ6L6PsgibKkv6av4LJWVCx2ziNJAScd9eYwUwN1d/
RSNyb7oH6N+K+d4L1kzL3eFP9K5Lpli3wbAMzlyFtW2O4/uIA7ogr36KKVzOGqHxTU2QWghOOLfh
mj8WV3NevZuvnoFT7JOx8+ryZFTtY/+0ueT1KyrPEKvVYkWtZjO55BgUzAYMWOpQfxcrdKcNBusZ
3Oit5VYotOExaQ2pLcEawAJnOtEy+Ubh+Pjk7UE5OFnNM0kw1prrDyFkqBxSNrF/S1HVAbUYUkEa
yxmNwEfw9WeCJevibFnhjocqvr1yO0H4Lvm13rduBLeWT/LfVaudYt3Hc2fH0RFgTPL0C1X1GVNg
0lCE+1iB9lEopCPGPztyQATQGkMhE3YHDLp0Bg+F7j2fg1ejFBaEJPClXL6Hh8zdqghrYylZ/8ll
chE7vNYW63LgmmcFpEbftlGIvtM1UHBK8vIHPU10C1zvvxVM2z5F3zjfEj/eMhgf/5OY4SAyMxRl
XjzgkVmd4agZ4qcPzOZf8t2jSaH+Xg55jM6RQ2DNpg1UCs5vSXF1yAKIh9SrlI/9ne2SPVWkFjt4
5bYKuyOuQM0Xp43OS1jSdqOSenn5dPsjxiBSVFgO6Vgv3bj5pYUMurDpmE169jhZ6LBtBQSSDBkR
peGqdxmhWIsHzKw0iJu8aCQKr2f4jQ24bIHKteS0vFbjzMjOi+Sjvng5d6XSq7j6YO5UfCBmgM1s
3+3HgF5zeuhlwt+YT5PsSETTkkLnfgqhrnivHtFguk3PLzq+jaSvBmbPNzlEJJDLuO/Y7zqtMN8d
DSK5rbVC6qCsXRHV1xNbsDvJ5ZSavf4J2V/aNTsgVDIvQda4xrE8HhYZ1CXcPXCt3EmA81JB2gAF
6Tt3t+06nVMj1ShfzbTNBCJqLguiCvhxJQg3T/hIdX//+1SZKf80cTVP4JVes4dBpOIf7Z2ewVL7
xpEU3SwN2BgC3TDb+SonkVpkuMZgv2NKP2/nY0UAT9mRaJc/mZLR3pvtzU6B9vLHUA7qyhhfdIC/
RkVaa1ifgM8kJlXpzTpz0gyszvqZHpEUouDRKzSekKWoEf4STWIqxDknO2vTUk+c55whIIwSvslE
LEDK4gMBQ2i93fZZ7BW760PRmlF4kpzLvRpYp5rk73wjL4HJ8sdyqmU1eCBLp/FonocDpeNaEEi1
2JWawJms4jlm/jlkDbd4UEk80zTWOo8lauR/9x0IuOg2/UfCpHQyi9jQF93mx2W//ZtF5fwUM3lS
pXUsj8/7HRoWBZZePZOO67KvpFNO4PX8XxvLZYpcz1TViGzKt3QR1BIcMnTlL2ae+YSiOKXTydZX
n2LYrUnzboddTPp9CZV717RjOfVf8/2wz+2a+rz8ULjNMmDsDWrcWHe4yQyq7x2bVj5elWH/YPQr
lAQInqLow9D9nNFb8xbTEy+ueHJxry8lwmY9QtUqW3J6tgtG4PFXxUmT72WvJR+voYgECTMVGTCG
8yvO5OfMjPlQEqvilQNOnZhsesIP/VCiibgiVZ1yq7naRK3hs6/Q7Tu+3o9MggMI9uwLqnScKAeC
mLgYYtDUIpOKEzgipm6rSqYagpJw0ltROP7c17sxZPNLlh8MvbT2287CvXia/rtg3BVOW4Rj4d2x
4cIvBQqAL5WN3cpOslxzlI8Es+HtbqtZ/Zdh54mpRg8Ybzyxn/4X8m3IS4AQRGbFvGzgRb9XrF8f
GlE5GCi7is84JeZE50oc6AkaQS8fVbq3va+6edshb89YErsp7fnhtJ1N9OJefdmzT0IquzN7yh5F
QQus7+IHU5i6nQwhg5OTY/JFIMVK5KfDXb7jsjARW8LyD5/TYFfJMJ5xGuVK+Yg2zYwVjyFXdxQb
7xpuGrSV6573L5fZLwMAHcQBJ2AifOtsM33lr6Kdxn+CiIcT3+EjrHszQLa0BpiJyGP9oT7lEVzb
zRHZZ++wQ8hdwzvnVCEhJSuxpHN6lvNMnnIzwiZpYbjzc2oLLP9KG/rZAxnlV8vvktCqgPykrvPQ
kTPeP3uzHlfyn0JCE3W9LlWuM0eBsxlE1KJsDfoG+NmBRmdspklLMHg4NcKc4SgsG/VUVtqWeagW
W2VHkjrLbjwKrML4crm2dqal1arBWA90yDkT1qAXc6d5izWRMl1S5lvFvR5hfckvCg2QfJnRMYzc
TdhaleN0pf6X+tfP2JFtzR+SjOnktE2Pq0A8aVpy8o8lHu9opcLYwiGhyuRAbOBWSlm2WKc+DP+J
EEu85PxD2lpTF9IG7p8EHQvN5hn+Q9YywX2Nj5tJhQNnLJguYWt+5vFJnyrRpxgIrPzYisRL5inu
1RApY/beo/R9GBNQOX/6loFfRTkT5ae7xCemXjRs06bZqJ5Ef3BfyCva9N+Baq7kqMRFWocTS7jZ
ZKN8YZ3pJjD81hwBcys0uRpDIb8LmHB26XmBi4x4PB8j6FDTZa1USPf3H2dHDSADWIYBt16CD5hI
J+IaR/XXKTlmH7UFb8vx5JWSle6r8hY+YhDwJKYZxaEcXPOdLX+PXvO94U5Kbr12TwYYtpg8dc9b
KxSlL5Jsq/qh36IALfAb5qIHoVzF2eMDWi9AWx99oqXfualYdbSTzldhb6vfm5uCrlPgEmHqhkd7
zC7T71q+VTBxulAWtB/YrhJCKY+7wXhe9QC3bmNyonOLS8xPpo9WZdRfyOxRLJWnEunNG8eHY2Df
cvWitvryGfGLxI+zFG1hYsYeSAQNtjOkJ1AhG5YQtS8hRGOF1bOJX3kDg4A8H3xw2gwaJeYmwBUw
aVVy+HAR22kIauvGeiYqAJOPDbtBZpS6g0il9S7EGhGPrVvl0K3jn1ln7P5LFnDbodwgpZQLtfZt
qfTcGB/3UXnSuwUe8IQYLolKR4oE3k+kX9TZk+wzymAZ26LxIQYnx3go1qCp+CJNfTUqk5YIQKls
WDurRQMdaZ90xoFeZZGNcx/MhCk9E2U8JGCN+wRxCYcX/vUhX78TnsMixq+C9mIBjyxnxDEbgPTF
iLGAREuczrS7eFE7MAneXML5TIWEbmx0pRBjG0CN3liPqpVbAD3Z37J2pXdXArATySp8rQjChx8w
3HWJNEdMS2sbIpjliwlP3szVE9pDksp4sgz+mKVMkU9QH47zqJ5ZPlfmoS6C9pLFpiPurQTUC3+U
C+gVj6pMyADCAXZnIPsxVrQXArToT/JLINyxf7czA0RByFRO12UrETwSNWKIHW/GlpEScrCuoWr7
StGr4CpICJt8zktBzMThcs3SZFPGDIabkUrUvNx0f1GV/MZ1omHJaOQ8oOwlcIGI9B0ocvsr7bBy
IZlvzaOlBXXJHtKXLMUMFQ4hgMawyVI9LnIAVK+8kUgQilyEzcl/+z04tqRKllKVIawCPDwZb8fP
UNVZwW45PYY7CFt9ng0GO8UJzBoDEoEyPgbJcHq1ltASxXuT6PgOPLm0a9DFxHrzNgDwc6giZJwx
j0jRpNLgP1+QewKm5XJGZ1NzD0ZC/kXZjUR3T/RyxGrxiet9Y8rDwN1Ct31rQBpZG1EOZjFVT1hQ
G0nhqY3zd2YWgkFi/6RGSRMU+IXQVVvYngpNjc1wNsVSJcsgbe4CVZG5oghbEZ3QcJFk4fri3+/D
U9j//fhjTXVsG94jHzUczuy2AT6zL1LGpyObU0ZN55RpH6f+TBN0ULdhvBdn2Ja6xhu5agwfPEmn
RdT7UvNpNXcCYjMyNjva0c4+cFlikcBd2ikD52PmdYz9UR7ZaB1ufsZAobOy9QfP/cnS1PkLFHyL
JIXipnw1scScVmwxWAeOj623XwtwUis+C6W0pWIA7D2DC84DQVXw/Yo327DQddxLi3Pm8Tt2wUpF
IC/Z0rMBdP3DaRmHqpfSZ6H+/8EwNktDPZRJlG/nCIybxqjUQsJHhwl2JEUrJ7bx874kZypP5Jyn
q8IbnKq2LO+xYJ1kZfj6S2OrsYjU87n1WqD1HBhBmHsaNHpF0DndTJsnxH9IHRqJsbEJZRq9twDG
cnaVL6m52RIiOjdNu0nF+du3f1PVHrXTPFJskCJI6sYCXZvZbOv5qCe+jSHLQpQOHYgDlseG8MO1
MiV7H19slvO2uasnAmsGojtMUKVDBY5CQdV8+2Gn4Xg3y1WW+P865lmeTgZ//x34l1ez0Ajz4orb
KZGt1l21VTP4DGkb8S5srYm2Kaz5o7sU+Vh8j3+ttnOO65oFpiyMRfFGBWNlGyxgIpos1LV+ZdAx
nH5lGMZSRls+QN1E4HystYS7nFiobHlSGPMgUtRSzdTJlK78AD+5aHKp29Mk2AZyZDnT7BXgA5Nn
YuEf3lOPUaDShE6BfKhBYlvun447ZdviU6rXjAejL7VKbGaYNJWchKpvco5YLG9xREUuSRifjyp7
Y8rwxLjtSOYkVk+HAtGG602uljxPdliWVKvnAZCb7nwsNTvXfGx2GCKOLqVFgOe6+ZH8Ke69A7v3
p8h0ii/1eSSzrR+hZRvgmW8kpxsBS7qwmxZgfk0+1GnGzS4g4jtslS+r1gohYzkt3TtlBgTSeOR+
CUNVA0v2P6R5FMjHaIjVe1D4yYkBH4xx7G3OyBIjm7rTGSPUWBkEckE/8tNu4nB1UIvxdkCy/QDP
7S2ynyq/MrIcdJyodC4WeGuNKPIoBIKRF3J8gO7G3aDMCEm8MKHfN4zFnbN3XZX8olWpT2cmWd36
fY76zQWnuJgs0UE0pdlmxz1YOLxIqeYwPVGi78zy99EJxF+BUifs6DZbwAbdtx7a/Yqcjy4hIGuQ
UueJJQMrpCn8X8yf3p3pVkga87HM3DmsKRm0vLICpiUH8HcKLd4kG10wfabJRQxPdbYzaALMc8Fa
41Si/KTAjYQ3GDZT4rNb9xL9iPEYTE4ioKWvBgkBbykawDo52FpodDR1fFikhbcgL0f99MGLly3s
USBgFNpu2z5NUVxU/gj+joY3jFOFAMnGfqUQtDYT4Pl9YsGEJftmdOl1mP/G/AOp2UA7B9QJV/zk
26bcdslOmFxWOdR/QCXJjfhRrUUrBFfx2Gvn+3K/8/r1jYpU2jMkQzdSJRlYaAGAfbC9wAWurM2u
Ntk5MkosjAJSZyTMXExeyQ4/C12lsN3unJRBjMpxvbsBSjZguKpNejMGR/zBC9oWvWbKdEkshTjC
sLQ9kl4rS7jiDfnGB25nP8tEE4zX7DkaJyMTK3G83b55KZUkj/Bccwhpzs25DhiiTBTcDvTZWz7W
O9XRAyVzOQmZLf6wd1IaGwPctsJ0RVfNfKRjEuFIW2ZB3I0quB2yAzkYdUxkqlexEf0Y4e6T6DGp
VEPAtZIYw2c6lZeg1oiyl9es5XwVEGboclT/a2hPiKMI51evl06W1JR+uWrfbHYvUKNedQ1uNl0H
AqVPwkjjnFuDONTrpE7UPWSBbAPEoVrrTz5XJQjzw6lNBUIDlV+9aYee6bN/crltAexAlPF2WB/G
iNF34pLreUIX3riOrg4bJALIDueQmcBRriumLwQrOhpDcT/sfRT35BM8+MTAKdgRDIQ+/kBZYbcC
Nxb0l9dJrnbqZ883AqNTlCUQ3EP4RRAsTawc6Ye/B172hV/CvcqYCE3Ug8dJjL53rrmpfhvE1KUC
dCeqeXCllBWFYzicjBDzRUFJOSqVO6aetmlWZCkNgeXLkadNt+23W0Ju1Dy0Lv1ePN1PCUCDWtO7
xosEi56JnPMKXfE3mj2kX56/5WEujeQEzm3OwG5cX/PYlgnYAJURlh9deIx0mlJHP4R9/mY2Ptlr
iSXgza94QPU16mUP7Hdm/0/bWTY6pSM1zFj3Vr8YTPfc/whzUI6rsbcrqJ+pywoKQistZ03kX6LX
QuuC4uqHDbwJmDxKGoWD59tcEJDJ3mWKhBZZ3B0zgRNFnJk9dymsWUnTk0TJ93AkJxjlfLN9F1IX
SkSl8Pq2bRWICrEqZtH5WN7aq4/kD/Ojiou3Ez/4hfohT///y0RlRA67cFdu0/ZUx6kqVGsZD4Ny
IYsdOpP6jvl1lFpOV4njW/7Ng121DWIsFPZYEgHnb6ayNXVqzYWGuOOVSFzcOgac0UAqe9q8oVlF
TN31Y4ym6qnWi4U6rP0rx3HYF+1gMWSxRCZIRKkcgMGnAMdt7IVtP9xrbFOuiHzQQ7dYrU+ykl9I
KMQatnuR/V9Zxf2TKKraxsi2JDD6XgUDXcFSVoBhANBL6aPo8z31aQtJ+8Irx1nO60IcCGbt7Kyy
z2hnd9VBYqRGDY+Fmw6bdl/jXVZx7GcO+YLx8G9ncf2BzMjkUXi1CvNiRAVYJIQ8hP+uNP97WWEY
HKu613j30wbU57u7DtPJGb1cqbZON9Sz/JWoFQI6OjRk6adSGN7M274QiZQaIoqiN5+ka+RrkdKV
b6Vt6agWpEGjVuCwiJRndYlQa57NxgJji+4ovT9AeV0qa5eujxBqTZPxoX7gTJUCQ8yMagd4jHoY
Mx9gQliqGDtyM2LEiJP6LUfXyjUnD3A7D34EQermC4S9hCDbw3VcRNfasQYuhIIH2pK6PxOQJimx
d+3fDTYcqYlAVSk4tXL/+Dbvx2ARC+j0EUowNVTg5hDq+BO3RHu5nrRtw10h9+kZoAQKiU+42lny
V7vA0ceKTrMjWGoUEkY5WLediW5gwB06+8oU3T935UM8p8I1BwvJs7Q6IyCwXPyXgoU1EGAyITJk
sSOfNZspOSUWtN6Wl6xQ4/RguTdq2HwiPDDFwfUdez5nWn5P7BLbFGD7zxfAUdD3xDKlTAUcepRc
0HIpEbje0/FPaqOxdZoiB6NI1A+NQ7XOXjzE7b96N+r7c15n4zKDqPdLc9BneKHok7feqQw9nLRO
l0kbdvh+p5/zRSJoB48I+eEpB0KLu+g+YBLvG3HKJewHp0B5rZJLHs8PGjWps76duPhewzocAMub
+Alt8Xmbi7K5C89Km12+IvSVBqdPNEy3scDyOpLAOvTMWMOpMdXDpIKTc156WSmXZe8qkhMdl0yM
rHMOQyBYHRIPmWv/DCWSHF1SqNtRGZ9wMxAznQJqBUbkavbP6djhBWw+ytC6vklXA6XrjUVoJxrZ
0c7nl9Ncnw7O6hJVEag6jeMCUbFJEAg840fykohDe/Ax+8VH8VIFWySulHkMgZda+lkyl1HM0LCP
QlMpFkOCN+mNQfD1Czu8mJX/Wi7QYTpfPlhZ57aSRyfD0lDAkTK2qE1/oWnwghihHVpYLDN5ZvOA
KL6mzuxuEszZuh6yK8HvrWKDfW2SVaC1bwFAmbqF253LUnB8cqeOQXLFYMaAOCKIP8alH+TCgmA5
9dwXRbstSO5QDZlRVWckm8QMBBJi9fD/SdprPg5Vbt0RLJo8l8/OpKLqE2Nzb1gJdW0IX2MlFgLy
Ylc/xvcQ11R4U/0GZt7oHadlveUuaonAfOYZKKDvJqC3g2ConKKI6isUIxwOiDP59l56miYuxi+3
J9X4km1Xosi3KWEZkvTADlATi4riziJBTwa8kL+UlHCyKFa2zsbZJ6xyrXE+MdE0cAG5xONANzns
SC1oMAN6accVZMqWjqDfDcoBOt8pZzTE7UA0N+UYy7dEEvi9uu7HZV7mxfBPu1cLL5snHG3Fqbgu
Tj9Mrx9rCwkztD+74i9DoVMK6PWjk6LOie9Eh1Td9gfny7prxbh+t8zFd9ZtTWTiyM+jjdJK3ZRV
w86hN540cGY+nZpeCKSv3gp5s5/RCqTPRw7ZO6xvfZ6xce6Dsfxj+gb3RIV6DqOpK8S2zWauc8Jl
40ZUlqjoqVqO4RcXcUrTdJmZi+VluJF5oMlsE9pHheT/PWDr1NzLV0/Tjwh0BnPeDAbmyAK64L2j
0YvtM2QXwPDJIRU/3+Jx9u1lrXPOk7cA9C5mnumVrj37pG3vjeTVxRtjy1JNrKNf1h4m1vFnqUFt
p6xuUtNidohN1d9sKlagXNXgbXy6wEMI7hesKQQ1ZIL0oh4PGi+qEZ+s/ppJf5L9KYHd7HwO2Ajr
oN5aQiyWFNR1cGfKfxI9xWCP4uDnhylchYZOqx+uR+eJm2k6sLnGXkPNsgU+63KtYxu2RqPbP2xE
VMPCCVqqmll/3NDhkj4UZNoYfiP/71xwdFsadTmLxO67ki14F8Sker+67/ytEP9uGexRIx5dHs7U
ofLERIRZweMKMcMhMCBGs0HB0z6QkA3k/5Nd1HKdlQFfVTS672liTaSqhcCH5UejgOkdkyYAXaZr
3Wp7ye9ZJJ+rJ7aHb9sz3yeDCB03+tWYcUdb1tkB7F2oUIBlx7PqLT3V0/4iOQjkhEO3BRIY9jD9
nx6tgK2L+fON2AaiYQAOMdpsMTwgb0cDlslV7om+4RtdfFopN46JvZO9CWEIksCUoDFAcf4MHucm
ekzWxbUuN7gpsU/L08OvPTIzlktT3jcJYXAl25jVt2r6WVL1PTU3M0NmyYbdmVQoptMcIxu3RKJJ
2fUNyGyccITrW+ndncDwa1UW9VccCf33b8WkfVhMYJJdZAdw0ewd3Vj8ySH2/RlKxn7u1kLH/py5
2SAawzxqm3QdQV1T7ej42z85ZBSiBzqVCvm0oiBsKPGmPLG7R6AkRbIqFQnbmU7Q99gjOPIKUHbM
xzGdoQ/2W5wW658svmlPvkFx24guoQkr0E5Hm6dT1/taJPPCsvrauPNkgXMzX2q9mfekBj/nDrCS
tumq/6vlOimDPIF4UcRk91kEziCuyJPP6fE46vA9wiOn2WUkRPf6/+0JiPxQfX17CucC6fhmKQY7
TqJxWpeLmLWrIz/4NKKdf7d2KP2x2/AXV0zOJzyxQtB6eYw4UXfFj6/ecgzLpUeiCVIZU1QNV7Jq
kcZdKTt5SoRGMehCBkSgvRMFOAyp+iutsl9XM09HIaVTlquNtCLigTiINGhxkvMqwdYnwCrRkndZ
S3qSNNmEv2nVuDnRx4GmWyFRUEX7GaBTDtb4xDWzf04rnirOBp449t0Q3uMC6zOomRI3ofcOYgGb
/KXxKJx3DA+2Jl5CPTBXwHKuWd/FU1VL4h9veTb1e/rFfb1QsPfe90G7ZVXA/ulqhoIKxqB4ZC5o
vbM78wR0VlqE9kSsjEjTC2GvE+5iO5gKqB2cULYgrQv0erUL2KPrALkUjy4E45Kp6vdou9hNOiQj
Z+H4POHGvgaoEqFQIIWJU0xb+6HPI6Ku8083hAAYfbocvvOGoB4x3yRl5Z4aUTmzySdKJ0/JtRWa
RgaPhQg78dnOp/c1Uyqm8Wbvm9xvi2PJQbHledC6Zk6gNP8pizzH0C6xc4CjWe2jrzgnq/hMDwYm
DDeWFVBF/UZ8USomu2fCOgHMtU4yPStwEaJshTXpPTqs+nloKEWwtQmmwiWTsBXxx7bGuKoY0cwN
R2vMo7OmSVkW9eb/4i0HGqnVV3KDmmSqg0WVvDIjtawjSeUSEyeBduAQ6ZEQPv1QJAf43qvkO/ph
na5ahcUp98XrmvvhCASDqTfHNtQvoGs1Gxp9+/8dibpZARy0zFi744oItFRt9qI+S/32YAUYuWG6
WO8lm2O4b4Dz0uKXzjHXVGDAXvBNkRClGxIpculqsyzWeptgeZH2fOrcRMb0Y743Jk8RapMs0w2Y
UWionZPWbdtYsGvgDmOjGMWPy0pKfCqgACAVdfHQ/3RiwKO2HHAptFj3BaGfvVW4Fo+KUe7kxflK
yjjJPNG6PMc82GFtT76CFiD/ZU1jdC/W3OVeHjBuTVDM0T990HD3i7rMrGhUluKwH71vJLfnFwrw
+VbNZ4BXI8sMlp7hxIncWzRcgArmOC4IQHwANUSNIPC0aAny3c1w8SB60+wz0cwP0JrC8yl+cjUx
uYK3Pd52KbohUagf6DsYiiAHWoA2685WXcheRZVOYB+/Yz+dTlLpzkan0Yu7XncmnVwlSTuRzEs5
lOUPfln3O/+wh8g6hK3BXnghi40B2M3k+5Csuc2M417BdgmB8nBSrwWugfxKR5aguZF0rZTqUsjb
TBTKLpc3KH+SLoGaeWJeatOQr2dyKdaPcpeNfwIuLwbRqapOfDJ+3466fcT7hnfPOzbQk+eGWTQG
iTjpQOme16LoQlZ4BSyfz+Mzqk+yj7f1z5BLGH2Zf+EDXq6je9L3enubbdDTH6HFzXY0AQJpFxHD
j2CEKar5bpidakAfX7ko7oAAM2m04d/pPnpUXXKkdbIjfOs3XZKhGT0K5J/5RrtES8vza3hJ3Id5
XofNZ+qmu41mKB0DT0KIej90gjf78WhS5H2emM12x3DqX7kIxY0+ICssqQW9tn1+UXqhJg3ihF6B
pwEDM4lcPes8SE46mlY7n675HQyZ1ivyf0+7kbyXZSluCJ8RT0cEuLcl4GmtygXi8pUawXiJYnpn
cv+hMPYGftT0SR0/ZR5i/RV7uvLcwcqEc3U2wsBLFbMy/XFoY+grvn82tJHgm2hZe9cnAE9ASJDk
6Fwgvchj4C4QnhAOnEbeq3Nb913VvwYsZWZS3AlLdWaHciow+bRzWq5ozv/vA85xQkHeMM5YPzqq
9noSCHqlwgbjTTnemNMrh0ZlsX7TPQRdWShV4m/YCCKk+Tvp74WOOtxIWiXt416eXwRRGlJhiKfG
NccFkXcyZgOYUX2MjG8Fyu3HNaTIDC7KO/UOEvMMEsi0CojJskYGXKI6t4rvCcyaXWEB2EW5TjMT
5Ov48aMbMPtyQd0JK2D4KhceCP8Fod1iw1Myk3SAJo4Y2Lj50UvcHsajQqiiZ0Pk6G1yQPasYgys
gcJDcDluz/gGF99dQGRjvzty30pjaLPgnYiwIY/0xBgQP3OmDNP5MZ2Mxu7j3h2CSgIUtcuuvQX7
wwC4SpHwJkYMI/CisGiiWgvMRxUFqnPEqu89ODGjAExqQPPElUEnyhDFRh9NEnLqdkb06nVJZaaw
Re0UtXYCkBMklfCyyFENG+vgcDjfP0MEOQstaJQtG0MqB3SdqzElzDSvx/HBTZI0TTe6U89ZBYPP
1rEf+dpz67kBr0c9PEn2MjyAoV/LnY5//qawTrzeA0yqKVAPhjd0VmZ5JSnPV121XKitgeDsbiky
e1sN3RWVgh+b9GEb3jXFZU2XHqgNDz8ykJAHnfsTGKflCVgVrWoZEceKydkARltXshbR0lR0DlF0
MlZZ41rXHWS3LkI0znTUjkPV6q6qq29I8XskKdVBjR3RL/61A+2XWEAmTwJJ3lPXAtzetpeNf0gT
tcBYhoM+cZToFS4ANnIfzSxtxTgEwiOpW0uHcbXdESnUGLCt5R+oEJhxEcaO3Ci3Jq/rBg7YDiXN
zrJOdTnib6XuUZtzEsQqsUDGBiASkQ0qQJltApjYq+HGogt3lYlCMRQGcQSQZJkj0inQb7quvo7Y
HWySe8Ahb3WjSYF+zaoolGkcqhdTMpRYqNWFy3voRNfH3VJoYU3+vk6btojT2JzqnOVqHL5CNEkY
PkRJ4Hd+tebK8/jPDbYPKSpSQcH/rU60ngCe9v9EgCAHcVlh+aKdJcD5wuytqfbUls5+5KPIEyO9
12HPvIlplve3gGxpkWqd91JEsstTl3FENQkZhROU9CFswZI7jZVY7yiW5AyIUinN+iVYmvxZ7Krt
4J0IQDqAIZqjrJdCYq/4lQRn3TulYtcuo3GK9oBgiglyBoi2G7uv4EcANwMxdSgrJIkT9v13dafn
G9gXVdZbMY3WNnF7wSvqeg56KB2MRLxrLgYOk21QXxBk5qYqxVmQ2CgG67RrDp//zpEKhdHOEqja
y+wB0uQz+hkJoaqOLcjTvZ0sq+ysAsa7rQ25AXQoe+Erv0ZcMkiIzfL349Zh5hR07EjtwKahAeI3
ytdVvD9F8CKC1+gAc0+xtnSwgEsfUKFsD3yGOD8A9jqylyUgzMsVuG3TGrACZEi8MJ7T4VC9zXPh
WLUtC9QFalYEhrqbYqm9KzXgUMzxXH86sd5qwCvr1VurAnvAkn6nbEJioYj6lOYCNgkvipHmycYz
Etb+jbXp40vOqf4h0gr7KoQwlnNcYsOjj4k0bjb6ncoEJK6DMrVRIXuE+D/mcmNNAynrMBRUwQgS
DwSUSLH0QdPrwb08tl6vXTaUZglmGxRiifJ83r1LmyVBXnChjZTw5D0nfMNtFwrf8h/PcDV36HKM
2ztiZR6ngSSgLF0LZ3QwzpPbx4G5SZm/Z3RALIkGO+lGYkmn5ww7sfIF52EEsB+U8Cly3vmPTklH
wXXNaxFJRquB47kRtVYypoFu2FIu2yZwPb4p4WFIOYjxWSPF2qSfuriG7qOuJDnFb0hwtZyKg8Hg
WVHIZNoL0sLZlbsbLJ6mYwSTkMMtqK0F4R2wM0PT2tx+/eIFhWqpupDjnf+us8szy8i6iN3eSMro
XSEEMcVEOLirU4jSMPDgbAaXz9uxRibANSkcQaORDbBVf4d7IpxCuyQgJrYTin3TxiQbSN0Z7P42
UrKdkXCDlK4FV5JQWq/+3AV/iPmxsu74lRvavQjxsyFT+2DLsTv2fqhWcbc5DrUUTSTdjNOHk7mD
vO9QWeD6NTQdImFI4RJinSADHs867rOkbzZord6qvdECesyz6RMJiK6Dpwv+kz4mKjXQdUXXknV+
1RXNbLE/cGPDTES+2Fe5rN+Y6mFwzb51Yo1Nls/E+tE8rn/1ZLqcPbVe2VhUwKC9oQxzKj7Ld7GU
6yTSCYt0BsznuZqHsIJ1q8ybFZ0NPmfs5NKEllUcpNXQnTkFD3FyVfRGejkKVB/irhnqsYAK0lXr
EKlH8B/DcDSISU0+IrFlPEJFLa7P2ERNGZ63OV/E4Ce7B90drtOiJxuZr3IVIMqeSMp5zAXJvYMU
x7DE3meKbWh6CYO0rxcC/M8RR+L9hfdm3YyucKXfDqkX8zywrIyuv706KqNaEW8go2Hej9tw5kpM
o6mWF1IsumrGuKYbu4nQUG5hngrQ2psNe8u8Wugf+Fxa4ERDLtK9s5m10SXvSK/1AOM4qgDFQmL5
0IQxb1ZPygSI+gHIFq9Ef+rTS8hCwo6aE3rfaegbHyDeuf6rwUbNrUbGBjedgaE6SYpbyhV8+5AL
CBqdk2Bi+cLRn9jjmzcVilPiQ7PRJBAQoPIJoDPWKZPnh3RIVr6MCb/5S1vUeBdCCwzJrWUTMTT8
thj1QTjnVwSjLe5+w8We882D5UHLpAJH8mJXbt1nrb03XYvVlmTDdPIuyL6s14HRHNPotJsYVHiP
/i6ALAZO3snOpn5W1vxry+H4qv1dpqhk2K5mnNE4fUtQ87hGbgIKsMqEFCbPGF9J1bFJ/vo73UJQ
RiZK6xqwL3TL7pvLDZOKq/86t27oUrIsrk2sqIgQWi3IVOo1Gx91nhuuJpcaax/qMWOMO53mUybR
32587ZAtqroOz0ujfC4AwkPfNexwXmHQPQX5TdXbw38lrEYeIrvGpxMXXPZ5dkONubJmyMHnv306
00lhOwEjTi6PStmf4T3bPkBmBz7emrwF4bE2Rz0CuJ6HqYWR5uWViwny6FusE6lMvO/P4r1mciSV
7mkSKOACuo2gMKU0EOdIFLr5B/jADif6uC++TMKrjCQjXFUHKavJFsJtDZZZ/OLn9wcKC2x8GJGi
+DESm7b5h414mlbDDP+6jhLFHKHyGVKTnUXCBjXTWlv3KHX67WhryTunJN3iAM2ImU2C1acSNWhN
xRs7+Ndmz03Bx3xjJKzL6PEkRhqGIvPE7wwyKjhfFH5P+U7y2CsT4zEIOe2AcR6UuUl1idkcAHsk
It4k87N3tPLNn/waj4S/4pmQlUaiEnErUDnSjt8jPuEm9AlV9FK8cTGsSDcPE2fqW/La/I+y8+3y
/9L9faSqrReHJFk2GiPKUjx9lA7h14UedXDKw72wntEuFlDzGhc8l+ld0rCPz8JD973BGkHKJCCn
Ij1r0KYbV0nrv1lu8yUABKlT1SDezuOyc1Fm4Jdu5Pf0J1AowZdZ/kAPGYhxDV0KlWalX5PPQVHx
Zs3/TAV487CyyOsvt8YX16V9jVSo8vJG1BSwt8yiCpjO8lW2QWHG2xf6X7Pozd0NvKWo9wHfRDQg
vtNbd6nP47OatH604rCrQT6npciCRHv5WH2ehpwcnIcJ1G8noJHbyvo8kvaeFwSGsiCV341itWB6
4knwKJNwPnA4Ab6WGWnV/RMbvpde6hp2z0WczbB8v7C+ie2rDUg9VgHSV0mzzlIossgNNX0DDjr4
8hWNRqLTCGyFYzkyvMAX17yWNqZYtVucEKig4oD5DasF4ONcXzyDbM78ccqbe9zoeozkTSA0yfs6
9lvcRXryB+74FZMTQqh8/pDCqWB/uE6ym5JfmZ308lgeyshJ8pBg2WzgitUz0HrjoADcOkssZDLJ
JCvgYJMkuik7Q+OPZi332zV89lYCLZrpysdyiryLaOGMaVJWEy8otWhUcxkk5MlQAOhS8Y1gObHX
N0lpm1DHIYIiltNvfxVyKbNknJeHJCZREb6UnUW2gB5oByh2M4oQ61bKyUdapIrjEtxGm/8j+4Pt
dg6LDHgos0XitqeLhOnFxUiOo3PpPTP9XOzQq8zwiFjx2OOWRoGpytInxnGGcfa1zSX2/9q8ddXU
VAJ41laBxhE3cO6Nb+FWVaAppOtIhUjawTOSl+7t+7aHQlzDJEFUqUPEx/0jQ0sAAs7C4MAU6OGR
HUg+ij/+a/3tb520uQvF4kXAe/y4Lq/0ICTtSl1rjoPAu1UPC2g6AlJS+Lqo1nP784c9g+mm+t1a
f6LnpghRdQ4fw+glg7c9PKD+nHl6xnL+U4cx9+C+TtU1u8A7jUvA2X6gXQmPj0XRqmZdE/T9FRJv
75A3SqVmyNqu9LfQFiKF5qe1No9hml3pODrbDxo0bIuISJZ6QxgPeUn6q/OrAtjTnKvN3Jrbf+4J
eb7Md0L+fhnhJ3UE0+XJmdSjC9Oxw/NNn5Nl3ap3Vt63cpz4jgXHPNXKiq11qbDZvxbaCyUruZfv
9kv6xbkiCw/yC3TiN7VLszBmZ1DokMyo+B0d+mu9ruw0c4iyoMfxWHJ8D5VtRjlMoEnXuYWwlikm
mvcitE6EiM/xJTC5BNYPWJrE5bYxjdFtVbFufuDItXZuJY1e09N6OB5eYYMz06874FdkK/8Cvdvn
A14xss+Xnie38Z0MRWhTvwITPX3xswJBREsvaIapsGe8Hbpd1XHUTCuRxSIGufPJm82MnJ7gg5bs
IpvQki3zBUEoatS9yjHmP6BV9XW1EV7LT7xISMFauB9RpCUuXJXRVG17FO4fYcrpMeIyxvQlRw0f
zj/wIpNGTVD6DmCrzN0QN4MOBi/4kCAh1r1ODNDvFj4ei3gS9mXVEkomlqO7HcS5YAiMlFft8cSy
Rh4zt3puA8pziE+S8yjdr17VMzYbvqUO8tTKG7MpXRxL5lYkN78Z0rxmncSIZ5f6b2mrz8pKRfCo
ABpeJl0ZfAJhOl7boB0p7UTrOAzVBS6g7U9ZIFMJuJ9VX/IpwBb3fLr6TDqKK7pYbFE9BfXQoC2O
WqtAOZ6WNwkgjeOR8RrSJDxcK/ItxVECLG1Ds6qD0TtqzqRvYAcQOshV7pM708rk+ozuGS42jMAU
8rN035blCYpT7BIyoalOo64plAdC01yWHV7nb+PlxJ1MJLSG+lvQgQPYWwwQUmrsvhCm7mAN0UdI
mMVSFs2MNcM+KZEiF0h/ju6mopOWEPr3NWhuYFBvo5MhvSinfIpUBpAEqMiZw5rGxz7oXC2ZFSYA
GHTFVyg8nh0zHypJ6H7NoXFidEdE5dVdVhTjPdxgmXiDhzjxSfil6bLG4bV1lpztV039yHKBomke
HTBIM7PiigLuaOLLfkVsySvl1uFurGmOHbD9Zgj47fdKvxJtcMUQdWmWMawVp2QiOSlIGMKDclZ/
YH1AYQkMwuPrfPQfMywtR/VN5HEG0Sqs3M8QvuqfPw0LxCtl421oQkbc7FmM7HDTYSodSUTL6LUP
VJjUSzTQSkeGjxiViIz4K0XbLtxC+r3Nfl2u8pnyCfrcMfJr3Wg4HOw0hX23lSSkU1IjpCJ6puY2
wkaycBJe+SNvfQxRDtVEsz10jSl1pFscYFBfRX17i/0YSleAq5P6tFsxcHMysg3l/DdOe4CUEP9X
q/KjON76BzTYnLz3iZIpJdAT/aEBeCKIaAwq7elJ+aINXk63VIC5c8AnB52gPNTUMhPVt1BJ4CHb
jqCPF13rRuLS9paYw8CJvzLEUjVVwPm4ijZBGEgaCSWgGIwwc0nSzqVKuPTQfU1zVZ5EVrxMv5M4
IWh50tkGw/T8ZGpemzEgRJ0kgDd3lmezuKxAoqwFY1i7xA8LbEo4FwIZ68EkUxf9WzfMdG6ux3Do
3H4Ly2RE+Bpl1iggGxtzBEmZ43xe8nxz6GvEJJe64bHFCGNmmtcAsNyQxK7pxZvj3QiiHYy9TqZZ
Csf2Le7/eweuwzwNPOtxJiNSHZ8Nnj6D4omNFGWz9tUDnZJhDYlHuK8IAPojCqjITiXR9VX1Y6IJ
yiLUQqrV6QpgF6gVqUV/esamKo4sGdHvavD6qSkD2nQNKR+nURjRNtxvWKs00xwMAmn/ktcJqHh0
LlLpfylLpFd2JK0y3sZrym0VMjGfloYt2+Txo/vC9inSQbzywxqj3kHRpLH4G8jV/rx4+tVfHX9R
yDron9oi+yDeFdMBSp2eo8s3Pg7SIDT17dOdeKug/KEKCwWWH7cXP1KZtXi9E8ASO46HwuCmQl1x
x4AtmATqloDCoxrG9zB8UhXNthcSPh5lSxxUugCUuIv7GUADWswvjnZNHkeweb+rrx+yvvPatXE1
HYgSByx5+8YFXYbCy1KZZjGJKBbKif8d6oA/GnCJyrOl0B/gc4SVnhvHYwiV2LqfuFL5aMEIDfWq
ct2H+SNszRgPX1cPjWnEYRbOU5Q1kB3vAxUS+Okr1Bpusrdph+DDtsfj6i7tvzokPK4/0xW1xTrC
O0GugAg7C6/tq9Gk/ncfNrdqtEP2yUUZyTH9IF/WAOwAj4h7VVI5WYZJIBl7UU0nuL1pL1px03Ib
B0ybxMDl8oU5JaAwL6qat+260lzFsEfHN/TGPSf2CDhpM1lkP++WwIBC1igBiVpA9IqCD5rAZljk
mPFV+ae8Jp+1UwkSEZPTeWn+8g+pKsokuMj3IP2+GkS1cnqZ2Srx3i4ZyPsBzyPC+xaDBZWq3Pgd
ktIPSl99LGYa0xeHeBOyM3Clm8hwfWJK+k0X3bHYAMRgAT/HBqFBkVT9DCIFqaDnIvoth23G/m7W
7Hw8wUGoJq6S7vRHiZv47urGvZeu4ad6EPhyIoWkhlTcu9ax1bp5uQOeu10CcsWCYymOKKJz6dmh
VwLE83M0RCWXFM+PcD34eCgd1Pghm40hoOAFXq+M3HVAHoTaRh1Gg12Xvik1xqMYBpm+Ojdf1oJI
PeSSEP6S3HBg1xwfKDg7qSM+trIqgoWQkxe6SS0m+MRiJz5mz/I8wqWbE/WyqBOTCebbJthvclRs
Ud/sWHMy+S3aVEhx/r78cfCivjNOBwRDHFL40STDXF7AtpJGWPcYMIC0nsDZ4tkJAmrh7vL/hCeB
XamO2ruLmg6/5gV6zd0Nn/+9jeE+DY972wx+JfMMUOEvPqWma2TTUFeErmScApMKlMdYvXugzKBo
vxc9hZ6BWrSpDeaUhHHml4S+VZcfDKZ0Y442gl8wX/Hmmra4NRYDMhujfU01E45dmjG3AUeg5aVJ
U5Zln1jfHBxqWKvtSsEosEjsVdZQBxbLQimGk1XiCNIdIflsSgHo2klAuPFOARXvZsIS9gOlwFHq
nUJi5uJiO9gry1ytXR3JpI0mqfUqDKRzPqa4U8DZKMTTZTWSg4hSsh36zv3Gb+C7bHOGiDBCc/N2
KDBEt7PQaApSk/ayf5FqKJxPe9c3Fq7AtkTt9N9Yzzva++uY/Zhffwe8TktF4AOJLapk673EDJn2
waAcORG0+zyriS8TwpDnCkTBoVkr0/pA5uIpCPoG7vh1fjd9VWLlJgAAXkvbUNVEMYNxmnISEVgi
RqBqVgtCFQfD+Nvy24f8IMaRidDNOhUwHa4DNorGG1n/7FdGOA1VHLhaO8ZmRqNIqyBnCvIVvcyV
HkSxvswjiLGYlu65VpABZu+0ZNt6Rjofv7/2Pbo7VnCmacUC8DYkvx/p+F1N46F7DQphxuvUpTHU
IGCSmnh7gESbilERqOov8ZOL4UJSpzHhh20LF38hT09kxb/TyC8s26OMQBEuek7npP2foX56Gvcm
M+w84HTPJyZ0GVOWGpuSzoyMeRQZLGgnBV06RfvnAnhLe8SVlqZF18XAs+abgMSwcnaeFqO4hsVx
Enwq29rMjC7wh1JUGVEGWisBNvq7qJ4h5030A1pBVXRg13Y4tU+4GHZ7SrJsX9gRyI+j9oDkSSlj
drBQTpHcXgzgjVy6qCB1RAD0BPyrbyYvhdp4kU7O2qEqZArWTHachfWNoictQ0qCgKyBB8daxXp2
kgaT6rl3i4eaJP8WRb9jYHAhdVy5aFUsOomk6PrYssRs/nBi+myq6MHCBKKLBZpZd9qCvZTH2IkX
hWH7I8cntw2xJqRdC3MGkgwdA7aoEhPKbV78EiEqW2YDXNYgoEs/qAKECD7wg9bCTG2eXiu3wpqR
VNw9acOc3Z1R+p129gt1wp3ljIioHVeSisdxN0mrx7WJXm+OcEiqSZF6A6ggsrq9K93m52k6iEOY
O8wOZua7Oj2RvTLqpAx1Cp688NCNaYXUJwsbHdLXSOmmQ0ykEFWGLoYrJvSArfsynI7qfwBn96mF
MJBNMMkRk2c/fbForwXux4jwZ4TXV7n0PKKBquDAF8BD32fhnPG1//x/A1KwljHVdEa9Z43U8mJ2
/5dQiWPGLP6kYpnUJ97N0j+1qxXMtaFuP5C/UWq5LlpgD+ji0FQ8a9+M7DnjqB8ovd2Vg7xrwTBi
Evu8cKUUsLft0WZt2DEx5rP1dlOXJY2XpOPd6CRuXlyhzE7tDKqj5gyjIbBydII6pYj1/uCnz/9n
zFJq0EGgJWruFuN/QJ7AsEVF8x8C2IutrryJPGyIg7VwrQIdkem8YoyvJVUH6iIhl8jVWhektoE2
o31DdrP4GBN971ksZHE7Y8gb4c2pj1TRFiIvO524gEfeN37h1B9A6ECcqxhunRNgEr33y8KgQVcM
B2o99rdpCa95u5RvWS+Jqu9mGzL3C3leca/2m3xCudylYABX1rE5TAK0nw2Q4o1B5+L9Nh4MlteQ
GqxsZ/GOUpLb6vaZ4HEfr5O1vUbI8LedXNLsjm2dcxs2aIMh3IzcZPmPyl0WxlIOqJQ4ucVIxmdx
DCbTEBvNyt8Sn+aYyJjAPOdAFZ0iqOO2iOVgPTlsHL3Ojq8Yf9vmjKvMUoDKWg3+GWNKjli1GQb+
cZ3sMS8Mdg0ldVE7SpdFpKaEOXRs0vFreJlg+sAFzkbNLJOatUlQU5lvxOfVWrWZOogdyer5Qjd0
Q+LWBhLq8tkGpQ5XAp6IBgAZZcvJ5qifEpbxbaTJx6fjgb5sVK1QPypWDZzagXM8NfPAkfx3kfih
RGYUy/ZvAaN9oDp48m9fOD5ct5E9uGSZK8umPugd3i6Tq8eMRblVsPprmuz+a7cdyqRY9OLMyRhf
gHl3acZlnpQTB8PLEXxTnBCPBNcZrS4tuLgp8XQVz1COPxobsCa5rPlmPz2VG6LhiC5S9PA3AwjL
rtDJaWCagOCoSjs1AUifUbRD59VP1MwyoAwI2MnRkOqHti7p5I7b073Dqcxg3ppBzaPQ6rdMpR4b
2NGpi4etRMzwmgwzWD/FYCPXwLTU7UC1N4G9VZzmYkF0vSQBCVG+t/5bWy9+Wn7h0pLzO1AmDV9d
CHzjWw+cCRYPqeldLM08jYzyh/NQJ6RWQM9JAp6gWDkMSK2r0K/Zf6F4Ae1mdD4eJlzGyHe0saYS
PBmB9M3/Pv3kOvWVzDulOwEOvoq6kmFi4bmcs1D85OoIysoH1ePua85hsLf8gG0V1if27EDUNWif
2sVnAaHpsAWsnFODQhQYSxsmDOwJ4o60DvQGAOlOddsm07tSveFU/8bsQgqiugz5S0rssqd+85Ch
qp9hycwXMoM4wZ7KWamXyJ66H7iXzYjjxojTpY00f4l28+0xwJSWWAzicRK3ab3vBNOsaIz/SQgY
OJ4OtMk8NuVnbOPV6XhgHmBwc82MnCmZL9gUWWJJ0SNjy9q/uoXKfRV1DCe/jAz5RqVNDO+4TKUB
TgtzHfyiqhCdaoCzyegXflPj5IHiIpLTT4NTK4jQPOh2uNXF0RrrtToTvlC6Ei7tVj4bXzz/wt0j
mmJ+AoRK2rdBkcjs4Qb7GlqL7e1CDFWGRo+3hG3cIfIsu5ygF139MaX4nU1gwqSCUwS/kJpQqjGR
b9JvYr+nga9aQoWhN3RdCa510h2R9rtciwHiAObulCr4rWwyRQS0akzerMU17M0dkFioKEIQ3qq+
0hZfI6HbRl0P6tR65LzxyEnTBLdOSfENibwUsy9rQo4NPWvOOcqECr0sTn3TmzkQuneU8aH9dwXO
9qBq5wCpK4fCLOKrLd5Tz2zk6mU0fz6KD/Gh0LL3r4uD9RKDBWjesk1jmKfBFoo49xxxr/DUOPj6
2qaXGTgR85o1h6rPLpgRw00zXiiI3vLVQQB8bRwInUcFCk+3Ov213//q/3Q9lLcmg1/ONYZWLtmo
o/xx/Uypko0bnZk88X4fHetd65x8jqtIK13fCiuPShGyV6zFnUAhxjeTllEqH+hIdXcvew1n+Izt
60dWLE0fFiA1Ze5VHYbig58BP5n4OPxqMHxKpJbs+olFMRhlqKKNHZPkznE9UL6OKft2s0JKSdZi
L8VMV5fZIYYOL+CpLNaWOCk3hjdH4eFltwh7a5jVh3SNIq3eFEGbFcVO4PvHqTI9JCrbxFNuFok4
/+YVp3k8x6+xEBRQ6P65YrDxmY3UGHjAPLO20CGeBuSq5jWsZgY/oQlOXAWYI5W4mA0dyK/EcN7H
QiqHBuHogCOo/a/X4MywaQZ4obTpkytrfTZOd/UNj/JRSW5Eil7O4WvSZbCx48UdHla5osi0H8PS
JZ1/EV243xUNJqIxCycLmPrDcvxfmvKPjo1H0SGZg+IplmCQjbS1Sy/5aduq0fnfXqKfBsbyuB5i
kj8jbUCWgt7e5YVfLQxVdZJ3XtnWxqawymmPBj+xlYdhxYvaOJv8TS3SxZYWjyweRLJBDsKNEHL6
QrWnocNYPJroxP4222V7Gx2OIJeJ6Q8yVatfPApzbemNNSmMDvtdw0imHW33hAbWVjbyqqqd+aoN
RMUpD1sDjt8wkN2tMX/STUmpFssv1yDZVlMi73k9Pl346LH/aKMNFeueEytLKmhOadIS7+E25jy/
h3kU2j3etpSuAhGAOS+UnEz/wU/cErwutKfrc/+EDiCcC8TCg3w7kruf/HJdPKkDTMOWc765YvO9
dlJZbuW8Llxo2PhfU/+VD3X/rSbPUDrujeDYmevyILLx9l4XN3WluPqcO2GPYVCbgjw4b5eox5cr
XggfWHQXL5YiklBfy5b0Iys9YkpfJxonQchRV2wVHObLfrgMhaPLnuew5A78OhNxhbNFZiVNShUU
xJnyOClKbtPSk7pse+FWR2TXqLFwmDPliohA5VeP/a/PbP2uG9Sr8R/dvJ2ui8oqA0XXP2ZTG7qq
UMzVJQxUECIkCK6c9WOLfWX75RpV3ZWPg6JfpA2sgKK//oM9KqUckYrh9GFPZs/Y9NASy5AVmTD7
+6sUHufh6a2jnlNXXCJV4Y4Z3jOsL5Jr3jyddrZiuCf0UnePjWEex4nCejZwVOYrj2yKMqNtK5jd
clo94u30hn7Y6R4yV5lctw8llTU+441eu+rLwFK6NC940bp1W3wFI/r87Mrpdr4Etq2m6NWUHWph
/88NLGtDCoDg6DM52n5ExfAdpCUQmMbIccYNY8nwyIAIpECIVmiUU1lWR0KfSy1UnyYjxVtTbBXF
mNFRRxZZYuz4YfBI4CY5hUUe0RaekCig/YVGKd3y+TutUh6SvHnmDX2j21IjziUtqvZu7ZRmWy3n
qGWqACpIYXK5WxoDOkk21HyOySYOMBT27PYFEFiO+Bx1heGTsX+og7Q9dgPkeQuXLwIgBFIvR9Nx
za6u6r3JQ34/GwazpCJcCWXBzbKiYCyr3PiUFkX7+7+VYN9mjMI/nG1eRCfZL01SY9FLAPaSMBi4
U0QgqUd+Nnf9005iBBe+8gRD8rV2KksgBkC/xfcYV/aYL9T/83xiwBkKoX1fmxBZ4sgjxW8eFq7M
0QnlmBB9rmNilmKinQs8LX+GOCMY0kCZN0rr29rH200bjQS24wzDpayGgIpjbIwaOF7A69wxj8Fl
OVbQo/jxV55FJcafV+5uTdotMAcA826sYP1e6bB6nln+BDi4RbsZk0ZeppvcVu6ZuRcSxc4lWDz9
AqtrRx3QPbXCXjAMhJ4pZII9gcu+Ri0ArvEsDBMEz2j5LA2nU6gSJ4GOI0NRQEYiQZeq9krffy2+
LwzWMMnNUwNNzph+BOBshwHYDLFc+QeoY2fbW/UdWCNAh3+jK2ab0c7gH4SbYM/7WoMzimSryaSJ
wJhxLWjxp9c2RZGRelTlTtS6l83RrVV2Y6HgTqy8NsYrvmoElcJsDRtQP6XlRpBbZW+QOA6YEm/Y
xIvr4za4MauBrKTeH6kMc4Ug7eO95eQwIGN9TpWKfiFbiMM8CDi4WZ1v9jw8kZC+/riE5Bl2qgje
eEH4kAeLpCZpGB/+8sLSpaMxCKKfw1y22eQx+WU+yfhGc5zjxfHNZpXPKbAH97Ag1J2lPuUdeLc9
RlKPhNdXEHImAv1+3WJEVQ7NN7mYfVyguu9Pe+MavZArcaBTOXgBa+KcYYbWXrDEjZ0EVKOexFwQ
I29tUGuzTqpnfv+kgMA0INXyPdHtyTE1UWGqG2pqf4vTc9gHElCVwwC3rO6wvzqGSofJifclpGQA
hmPLXcvemgsO14JUcu3xo0OoCR63s+KKEFsvJ1clWVk+L1sx5y+DwGfJ8YNrAvB0DbYmG1SGjYP3
gDgLIvVzwkateV0SL6Xhj/6EZrX8NRU5RIfZg5LTB5Dk3GmZJRhdBkmbQdIkrUZwWOHgKWlogZe6
Sp4WFqPMWVhAGLqH4sXDv3NC92oqHFxgnUnnoRHFOPUMdZlPGDMNOgsLGP3uDKtM1J4Whn379Rep
JXvqpCWEqFP+V8DDkmoqb27JYyuLgg6MZL4z8ud6+jOO4CymiiqDGJUAMKNxf3OiT+9QIgObUyfK
1gvBAQTqVYxSfFn6qB5eAJWla7pxBSJGf6FHnfF/eQ+8FU4i3nolFi7WiT4BNMnuexfjyNHJdN1g
UyiNdZRDfnPdkNRKak8pF99AqcoJ/tzUi1aev0/7ie0g98fKwOkswWlmumMC6vh55/cQdd92tpUS
d9xeWZnfARu34EfG7BDT2qsD4iuwktYkuIB5PfA5U0+oxhLj0WmFqsJ3VXHCppNsGRiVsshI4ybt
cYQJ85QZ48XUZS/DBOa5Lt31W5pz2Uka6Mm7Wmz10hpbp+nKAJ3Q2j/VV07MvMUoYpSQjrgFZhC/
ZsN86S1t82WgLOLplcNdnELMxIk+qESt4K+g+6XGzmRpSH0vyw/GGFSdR+entRRbzgX+yCY82nK/
2lm4DErVzb/d4f/GhP/phx/B8JOtid6CeI7pyj2e+shxEjApiw99o5v6d45TyjpKOKUZGpuLxyce
CVSlMn2ox6cAbSeKKTxpTX5NPu8liy/YtbXgieTnM1UUIwVDzY8H3MIKB97jggk6sVxQiTa+2ygg
9OAuVcTgXMgzWYVun79+8cBdeekuOp+W9pazLX5F+iH0h3dzDjWRfsDTN7v+0tFLnwpIG8lkV3Po
9lKd0v1O1ghH22zdveoPM2USMvLbNbkaAukQGxv7/TlJR7X4SKpBiOhXd+6Sr2q3KWWxeOCWbjhS
bJYDfxTo2F1H5djn6lWYWVpy5IiLNdEiDsGIlMxAH+izhSA2Qn/JuPW0Z/Gi8hc2oBAhrtna81tI
+4HjM7QwekIEWBQn5d4AJJc9qLYsTCZJPPQn4P3K+zpsRY1j1YL6jKkplYqaQDCT6wwOYH1SWhCG
5LMWRwhCCw8QmvmM917gtzi+Y2en8pPn6dabibCXMie8HiAkwxEpXmkibYqyeMrM9WUtHSg3jFNC
XfPUgNiNxVbz+1D/4MS/ua5jd2rL9WPWN14pPwLvE1cbIdIgfmuXdWcX0qio+jvJMMLOq+BsqQkC
zKitZ2RO267Oylhf5E01QGlzyFDaqp4mYHhH9FQBFehlT6pbMiS/ss9kO8vnknOF/ryZsTadXRIN
ySaplk8hqzvd13ONb8GdVjalSF/G+7ToZV/G35ql7aDhoAQrCKWBKID25HHdcg1vdwJo2QG2IvJL
LoJJg9GjAKJ8lfReLyug1hDJ6ZGmm2vyzvmQK2gt39pLnGB9iXf8RApz7K2IcvLdAswQzWhfNAwK
1D+q/e59wY3gUuiQWH1vKwgh0DFbSHVNEYSXYJLIaD043VR/q98ygb6DRbZER7t0EiqYbUxACZTk
XjrqabSZcAAoG9Ok5LgEDdj2En1l2ou9LKUEl2BPOdkjy1JMWFNKC1+LX2dy+Li6l+uTsPLbGXPZ
v1YJB/ufa+7y9inB9h0YOBVS38+n/C1ixkMA6y8IT36ERRe9RSQJOZjf2nKiBuMSSQhuPww2XcZ2
cll/v5VX/4rGV2yjDL+gYW33KHD4TUNGRlUpH9PLzfWUMb9Ao9cJdAceg14I8BpcqbYYcSyypFTm
/Byxtkg2GSnNRnOgIj0D6HSjM/Cz6Hoa1RcjEIPZ0E33yfbpEcSrtNt61LeqzF6j60bQ2Jz715E/
oGsccnx7cG0b/Qnc3aYn0soNoiOwJf90fGHHsAqIX0IaQWTrBgqyWOI8g3NDk+R0CKl3UNB4FIYf
BCwYB8G3zY8hPSMAAqU08lXVjpuFsyyU2/W8geHqPIoEtn+vYF+3slzsrtFbkpQAD9BiMhfcCCFp
+SoyGgQj/k9NUQmS6bfXtTys9wWhYGejbFSx1pK8m88KZbPScMC3/CL4FJ+RiU//GEWG0h3sNwSf
Hhiguyj7lxFcwNnAP+g7EmcJHH2VxY4Fhfy8Jo4vXnR6g9e/vG4LbW4Sv2fl8rCjZOF2bybJ/xRG
+ybl+gxOYyiOaf090urAq2q6NSEFpkZjZkmqyiup2i2uPbpd7nWWRHwhZt6oW7OPviIuLH+YdPc+
/9JPTCO3X0LAzLEBoibJUCCudgvKn4umF8t0dCiTj+X+BZBi0AYICKrxLuKrl3w+ZxjnCqHx2wYy
9Ul1m7LNjeFjQpMtRJRDVK18lnfSVA6q1OUnzylcHRz2z0Bv41wt525cHDZiB9nvCK/Ohi/nhjJz
TtoQ4PHSLB6sauMAfuYluAYPZtnSrDIyIheaBvSPbFhoT7mUIyeCMvqvPfL7ZReFdAKbsxAhYcHN
wG2zrS/A4tunDh7FkTGrTn0dZfEHLOhDVXun12IglvUxalPUP5MQ2A//UtqVU/vc//DM9AJHge06
aekQC2/NGWMMk5xRDHVzqdbUIR9t8FFqEr1qMOHgGUy7ZLZpsBnF3mgTFMls2HaCP+8RKvYSQp/m
6fsTwLSxQeB8L68vmt3bO+m0DIEPa+DTk0dpwZf0i5ALXJeVpX8ckonKaUqSPjWA/gBnoFGxU4gm
yoHZ+4VS5d3NTHoYuOiUeICD/9WRhXLWaDlzFBiaNx+5COd/gwz9ntlM3nRuvzRgqqLiVWCKqdbM
WIbA0R4UTXeosPXlJnUviHB/2CgGnLxzLJpmLD1N64qlRWKpmt8CAP23eXYNlUSTn2qxhhgxRVLq
qQB/XRv1xvPf2drJXpgjzeqjnbyqaklKEQeHpyOBZQ3CAdjMf3aypeszGJ6lHmVdKSZ5iXzu4epO
3WJ3fB2I0H7BZ4/m7SSXNHbQCo/a1S1GU0sycH78sOnjrbIJZjueD1RDOUulFcLL1ITZL1baaOqy
8grSf5AHTJ9Q5PeYl32vAg8RUS9J5Ua9MlGdgnn8wes/DpHayFSita+t7SgSgo0SlDYPniJrAgXW
Pv6P65O9A1A6XWkVOe0mICAght4FhXbEtc+Jf3iTOx+N7Y74dhe/2NeOB0cg+brdUJXutEa+p/UP
ROWS5N6WrTKpKasrYWumrcZ6jGcvnw5w4yRLBjUk4euT0/qd1Mu6HyNs6Wf2UZxi/Oe9IwqeMiI0
61MBFcxWL2wV2wIB1FVA5VG5bFD4PP12u7CP+1wO5mJJess1WzRAny8yL3V+uNrcWt1CMCSqJfg6
/uwNFdOQfL8HHsojz+jARgBnjEeQj4+eJyqUBV+CHsx0bH+5Fj/ZiOt5DEr/TFqHzt5pYN2IiLkw
X0WMTKQEwgL8GFQ1/7ANMAvQqvW+9RJ9vb1y7RVZVn0t/buMJq/OF034M21lcGW0Qf6gLc30XF/K
L9VgYjLQLRBQH38Nnn7qELhb48dSq8HbNgFU7txA8JMV5Owpg8iHEOkDNng+m6QECPf45UNznycR
MLGb33HTTSVWmoDgwI/tsUBDkMqAF065bThf65zU96ULm9FiUjfuy0gh1YuIXsyZU6ufLTg7z77t
Ol/4c91eUOEkwqMPc4rSuIkQigdcoejxx1JiOeVkbR/5ko8wgO5QoadlzY1JzqmvbmTDRntvnQ4P
+4ihDxUh+pYZc/KaPyYV9ac/R0PfvuF9YIsdF4JrAK2X9gnZPvVkuzxrl33Q95SyU4kRAZ6DGjA7
hmWLEfzNHvnHdWAnoli9zq2r/LjfdAz/AwR5QsG8/GG91XFMLvCO2GETDVSkRWFHPM+u5BkDolqK
x9xqQPwiXrk/BzPSWGEgaQWTtXFAlOmAWWweH0hVJ0c+xYPTghVMSd7I+VaSBnX/SHkIMZGkbCVY
3s8KMmfmiwiGftnu+4QfX/DW7TNo52CeIga+H52fdtnLrjHta5lwGDIxkkrwVFEuuvm9jWJqBLFP
dDjcsIUA7S6eFDoY10kQGp8nVvi410ueu94ostzoDrJUuKtCBXajgJOg0mdQ4bK+qI2pNjBk5F8t
KC+trYx3OwG9tKzpA69XWjZ13+xe3y0kLjtzDaPZFRUXCOXiqPxR4YUrUaiJ5MwQCe4h56iheOZc
GVpllcZ8SFZMCe18Nf8yHSQqLFK/ajNOrT6TKu2Dej4FcXcmF/m8Xuy1LX4AAoaOnGMRaP3TqOsT
EHpBOwpOmMwasuECku1fRNsOMkAzDyInklu7m34Q8LuLIl/F6lN8r7FTk4xzj4cQvtWAXsLa2cpD
fxjidDgz0vJpFM4fWQUBcdbLHmM5AHoMXKI15poWCydrkc3oB0X42BIZ43MMzmfs8i1GuN0tXfaQ
VFJK0wP2Nca1imLHuvA1uyIOkGnVCHurqmjO/DB2oxeKnxIB7YTbANTTHkb77bCV1ldoEz3xiaVm
Q0yvBmETdgkIb9yBSYIqNO5f4sq2GIMKA15xZIu90lEWkGHvrDdCmkImSqg5pIdOksKoDmqLO3i/
edre8EaJGSeK4/nM/JhpV+2MvgR84S6r3aOEsUbkrmi5rYA3kma69mXoZsAOoa4Ze07hyjGDiA4f
LnxQuboWRmafHXAl47g3H2N6ghzHryd4E3vTOsvdTXMWL+jzIbKNqissR9kZ3KD1Yj1GL3M4czYQ
Q9w+1vpcTelbkMveV5rniXzNvPkrSxizzUjrDC/iwug9GtNgpE1SrTCNvYiCNr2wsHfWzeYryqg9
JypDJ26U7DLyd5jdIwD/qvECnYkU5BltYjKB5cHY6NeL362ReluOMz/5av1icsf0usn/05Szaefo
rQJsayqnSNxqrDbwhPGsYFpctFyk8wsDaD8BnRlbE/QvhnmRgsShRivodbMJSBVov1Xg9JEsirx5
c0dfC3K9Hb3VfzZ87Fot9REn2k1iGTT1I2avJJn1wADt6nHcyegtqD9N4I4XfXe0EHtl47J3M1GQ
N2UFbX3sQZyFfPcrSvap4xgMJvffAWOzrBNPVeRtX4QQIdCOPLUegIKn+nnFRSrHQH6g+lYL9z4v
ZGAOvLNH5WmpypzEDzdYRRO9AHUtHhq3OSTRGiwHOB1RqC5B+ntgW5dWFRJ1wzgZahcE3hN/qFRm
Q0MFHfCtcJzWd1zrqCylXGuMqfJWzPld3lW+PeJP7Dy0xV8Ih0rLrjXI7N+KR7XyxKKG52q7OTtx
xjmtauruU8pfwy2Etj0nVirNdU0AE9frbjkKzvSTevhuPrrjTJ6Fi9nbCh2z+hFe6xZyqMomacud
tOyvYO/O78PdeYPSXfN10BzMsrBIr+1ipSf1m7n3biWh18maaKRXaZbeHsGrv0Py29lItL28+X2m
nn5J8tmidz78crt3kGLHJZrDSZ0pRRsS0Y34TmvL1hTozorfe3TmPeIz5VD+fpCsY/un03tWnOFV
YDiAzA+63wYwDVTNSoYQfJ+nUQXob0+84JYT9ZBUeAtv83dtBPvETHXG9UPrJ1B6IQDb+Cq5Ojkq
xMbL/cBKG+dVlRzjMV4SF5gLYr3iOqbbqiWRKn2yMMvbYi/DFEjRBro3srzv/OX0VXxOugMHUXdE
5eS2Q+r+xK7ve/8F6UP9zgOcwoMiCAxVQsf0iqlY+06tpwnHRJhtKQ+nhK7WUzLX9q/BvfY7Tnc9
fnXeMTb6d4fqvTA2r7Fii2xWAm8gHx6gZPG8cKTpmn5QDbH5R2h/EytFZAWUbYeG6bh1F2/Jz73q
23CIgy0H8lh1ImJF44I/0JzzmMZiq4DBQoSLJ2gzBsjdvrTXuzclJ5zisbPpV3lCMW1si61MiChL
QuPkmF4PKwvA+CGHalKp77uwpCCCCQcyH4HgjvFlncr0HED7SMI83auLDH8ikCjmR8UzVfVDyNVN
gxDnJyj7JVo78ibmZr5wjJhMnqE9dwwM+Dk6v3H3/t59gPJICvxbiBxPl4ZiQ5+CJErRWRzMoFbd
gDtJDDdomZb5YUPGooNU3+wzFQswlCMcuGbwcp9ZHaXVkFsEQsVRZOthCRSvGS40L/5hT3Ybnxid
waZIOVGOiT/q5j4cHJ3T/03lauh4stO/tbK/am9X98sgD9AiF9G2mRVpPC69fJISqe+hraSecTta
ATGAWK2BqsB2onGnAofoU/cU/ohhL0LH1YyExCzYXnKtc0nSe3idm8v80aqej3A/6MCmogsJ2163
SpgUFgN/lDE5NyW20VwNonjN5a8KLJ41JPTaXKXTWYBQAbgYyItDoq87tTOmHwsrpOmqY9tBg7Zg
pp/anKf10dyR7qivHfu+oCbOOeM8g50zmfNWce8nMCnG2fv2gsjG/6FbPrV2KleNyRSjkNsY6tPR
YiJlGEHw5Nb2r7Ce1NWJhTrwqLV3zJzG6esq6LU3TZWkgjnI7LF5X10ECQeY+J8Gxk8o+d9z1E6B
Tm6NnrHjbx0VxbCZxqIxOJMeV4tOLufGd/HND5HiORwQQPVkm2n3jkYCFG7u7zLEpA7FrzzdsLB6
cXQmgCWhMaU0fdk7txNy6cKGmk8NMEuU0QMSLJkXufGfDklA2W3GZYXvBHIf8P2zk5YPY7iGnddH
+RdYZzAyPRfb+8avOr1e5WLidUMUTE/znkw5Mylt+F2oH6GOgqrjQysNnHmgk4ZRQmAz9hsMXA6I
6NoDguoorDnU2JNhSyGafMgKqVo2kwwITVJQh+fqkaMeRis+mKhEX2Npu99veZ6rsMJ1pjoluUd6
xBIeDeY9HVefFLpT8YJRQfOHHlhYhFuaLGMhunoSuyBBZSpKafrfhRdaPv8oAkr84RMMTewaMStx
P/TohvsPpJFg6H0VOVjL6RDT2PxLpnhKu9zPnpvKHyTLqi27stMWtpMD54SZ5OTW7bS4Voj/vMZR
WDGungLhFG6Fq8VXCtGN7MwzJK4CCxa23YwBeFmCLiAbUM01FICNhgRn+E3Tjp2saFgqtDNOaCzR
KF2A1qr6EtN7w6R/pzoqecUwumqxXf/h5A2pvJmezUubG2JYbjqCqioG7IutCWvofNiKC6PUvxg+
9h0/v9HnYjBNxj6EB3jAgJoylJFm2T3hi0dXDw41PHzGRWK1qQOuKWfnitigExi7UoQ/twn/+Qc/
g0C4wCF0btZgLWdVam+oX0chL9RsUxUVdJAuA7LYKRgk9p4BX/yJhIg/o4iullbNNHxwKLvVDrVn
YhcJpgDr4HaFuxfG5BZ6jPQYjbwMR72/n0oaQeeWnS3DpWUP7CGkTe0HmWioU8rjAknl4VoqrhKG
r/cYgUYmCEKCAXBXi6X50P6GaDugeQuh3lS2/DMCAVKQ5X+BLipOByDKNjCkGRBWkqPmDsOLm0mH
MUa6SK+eWknuEnrHBeQMav0tObLCUbjLU3iDlwKuHldl4o+Tr2798vBZt3xUUXanJWTTWIr4Bn1P
JHxIJLu/tXl3qPDqfikicSM/2yu5yHyeaIluGpU6gKml475ngwML+/y5xe6R6vf8fyqzZPOtWYsH
zTLHfYpCOETezOYDIT1OP+Zflego+CBf34zOlr6CIR8MLiHU+4S8Afg6GjRx9EfPzvFejdqSrAQg
gerpoyvi7EpB95cAACBlGnGYrFtjIEE1L5t3UUvGZiyw6J7lOosg4fTS0SY8IY2s6f6BTcoLqnRG
UmqCoCYVPoWrrnzg5rQ5NnML5L2iGrQktGudlh48k7GyQ1XD6w4+s4l03dLNdsPBltHR5e/xIhss
d+ISGi+KVUlJq9z9HYe25lQLGKv9gtALL+WyTGhhC3P6aCUtQ3i+d4Wob7MYxX/EC9VCpBIDLlHm
yYcFqWwKewcALOlmzE6y4olslBhWxE9Q6EVfUkiRV3gdkaYLnxk9BwKtOgMsYFf+rNOnIYXfTwE6
4+EjNF3ztdMaihct4u6QJnqC5Ynnz9j1cIBXN0gpBathgfaAHGZklzFBZC87P3Grvk/KjU6LoUeV
sEp9tkGfAYJOzN58FlWGTP1kKOWLnz2QQFkEbGVdAPs/IARO6jm31cSPcxyLAwHUOdNMIwUKL/tD
Mo6D878Xu2pyEoO9T6uSTj4NHY3bHfaNwetyCaLZrx6wUsJJ94+JGfvi1eYwHPLb5cF7hedQQJn2
u+4nARheGFJ3vsG8mVpv9MwEYY9tKGAfvgMbEUUN44HDrFQBsln1ZkK9eJl9C3N8pvRxRraDEyiq
XUl57zdgxsEpds46k+1BCuscQMVz1/OiACieNjiAOF+5/pRzS4w+Tas4dNMiUD0y5ikjbwrKdhBq
rdN15lVvFsWeqnmenSiPY9iOCSx1jKPEUBdcFk1GAKoEBewKnuxIeCUifj+kpf5SAPzFx9mvTByw
AcyNV2qbcPNaD8GxqsauL7wEG7EWkCnxuQLv8Iv5teE7wV+zyuCDPMnU584TSDIKvA/5p3Lyz9++
bagDmRSgEmx9zIRbuNihVPED7TD77SjFQg8j90LFK5QojSErrDwMxzPJxoPisCj73IOIl69Q8PgS
YrVCE7uwi0s5GQMJeapvTK07qcdTKkBRP1bYznIuZbCIAUz4nvQNX0ELZXPaUyLpzcY1RXtvXzeA
8ZKajIFnpKlE59Kd/0fib00QDCYcElZm4wWuK8YudkuV/WK10GKHVQmYjC0Z8dm59J+AMxd00kh2
xpvJP37o/lG14HcN/PGAm1veuz0A7qw/NUd97OrMTynn0m0Dja5z+rSAndg/QXnqAaB8TWQQc4Wv
e6OtEfXy3ekPam+v+qNLNgQH2xnXEFAeuyyKkikVa5QVGW1GjpXZp9LKp56cgKBqTekcedWg0ME6
XTtCzfv2hVJfoKt54DmQzJ0V7UASgKOzbOeVBTdDiuZQVMdWsGTLWYKcamQIJ3Zten0GKQb9IxJq
aAnbsFjEHEGbQ97Onaz2JP63Tptzw9p2+OBRU12UJ21jWBLkzA0x2zNSCO1i2BM1nxmN+6lnD5/e
6kKf/rruIBn/CxAaGADwQwqKz6Jots8K8msyn0GmnAwU+Vnsgs1BsVCzsO1nbQGhZv0tlYYGZbvq
s7kgRsAKzT7rpVvj6Wq4FfSK5uQ+sYY6Hxuld3aiwOaRhbi9+6YBRTCODXmtpx2AqNGFlpRBF0XL
MwQp063Nc6LFKMiitSVRaYc4BJPd+kYpl3y4dFW3fwkSuFCHZ9ogTtIPZubKhlB7CWjAVLuzLos4
n6q4aiJzjkPcojdT91WAhLcU1VjriiO/rhH8ssleW46vUzFDp7rODQrAg94uAb6ETaE9vFPR4Ouy
eUirbJk6S3z6cCRPm+7nuFhha13Oa0BFBMngdLvzHJ63H9nCrP4AYKN7ANtt7B2hM803YASC8WYs
Vhjth1vzdZejdDIvEG3hGdE+gVtESNSjpvtVlt9UHB9TNE+nVEeuPUo0fnZ1/rha7BB6AKwjl9qc
JAntu68lyzWDH6nqncY0f464qVo5FLYGMvfZuSxfyyCERlgdBi2eLjU/tOHIDTzeHAnCyrUMzzkP
StHuihYIAaBVOucbF4E5DTV9xdBYKNVu42stMpuE7ZKqvhKMn4pfashEXzS7jAYtpSwGQkAghP9v
JdDD0C7JmhTb5X+sUL3oL4/7BpPQMY5KJVS4R+QxTyvnCfzJIdprtFtxc2cFDOK/pmAMeNeIoep8
tey+GBHkpkiC7o75vGZ+bp2Ng2UeUyabok5yAc7HaZh68qUpvvtTxyhZEv+7Ow4LEAejIbiLJK9W
AAbhfpaRmpW1eFvYprwzcUdn6eKxNY//CE9pon8SyCAz2Vpe8tqzlayWdAoRvSYfKMqam2/7xABG
vtr8NiYiNLP9nqzrONrANyNAaV2jNqAmQusEJLD4DuVge8iyElBCU33bXXIEsIiT8TEkjXpYIwX9
ojMkb3WINiNww9T4aQ/W1dkqGmzCL0oo7m8Xm+RUou3qGaiIkX/vIr66njz+FTnMEzuvpL1+ix1p
BDY5KoLcqzb19GrJM370U7F/+y8+M7czUhREYnfeOIotXnPk5BU95n7tZDYWq+fQ5YYHpZ8+eCI+
nWwvVM/J0mSZvX0dJEqhaEh8gaNLOS7je7RpXO8LRgcLMYeLTXzWZ+VntS1zLw8G3Bk0EMucAKCJ
eZbgVT47MwEio1qIwzDQFJhSGyUOcmDn2FRacGwozYWZ5WShEF5lyL3wLQN0tTbV+Yf/iujg4cMK
GUKknvaXRKdvyeSIAG628wUtCXa7ZXVjkmz/bzBHXRoiWw/yLcWnoJO6TAFGzb5ivQqnH7UmzSpZ
rJQ/xpFKhtuVe8XQ/vtNgjmjrVYzGQgKIM1rvgTycWe+7FyC9o1cKJcQq+L18/33sFEOnCZsOYJL
2ZbGA3QQJc07T2qCsVmUgvyA/WYJwGAPndgYEMqWa7tqmshXC8jLlYWTlVtg3E8U+PGcenFooMv5
3jXA3pE+fzXv/anHtCzUVS9UWcqiY0tI8QMQGOik2wqofp6WNfOIJvIvciFmP3kSE+l8HsFxRuBc
oBBltqlHnhYTSumUI/qsvHpIVA3gFn9vqlRn2fJfmUE8APWhZQMvg6B4OAJfUMNu4agwMmel5TMq
LMZsL18m8YQxRCQ1wVCSlSzPUhpMF9vlK+7MDuAteZTyxx51f9dUV1soNEhkcWRa8K0tdWO+b1Jq
EFR0KJ6Qb4aKmokx+bGo8azJCscw8JI4NHMkvuiIKe+SwsAa5Xe7ZziF8BRnXOuWXb6Fo6QdmzE/
01w6RIuT3Cqnmyc7W5wg7atT5tvSyaBNxiSZypDAHFDFgNms6WVoLlUhsk5CCy5IMyiFYM3WguVU
2RdFarK0GRTlwp6D+kMdbpxawMvWokZaOOdEv1esbiqNGpXPrB5S3gqyvRXIi96PdETd66IHsG3l
2DHbi6XddCZgQkQA82QUV1AdC8oslBnRkHcbaTL5jwAxyIlizH2BXnv0+hBo/tkR33Gv70RLjbDP
QSSEtWC6tM9graIb3Aoejlglr1lSFAea9HpbKBEshOzYf+REZsWMgx3ocw2TjdIhdmXgwQzfoSZc
7HMjUgerJlgQHU7nJRzozIOuFZsjXeIAG0LaiHZj7873pKroopBXmMUjH5/sKqxKV8gHM39MZcFL
K54jApJ6TAUoquvweBT50Fpr+A4WR5zYufsDJIn6CYK+UpuDk0K4PpaHtbtMpDK5aot0kSTnGyt1
LDX26Z4LMRlXQUrJdaPjzQm7otuYM7M8gaYha4cr/HrwHUHdJTqdfv/CwwYDCf8Hsxmc75pTVVbW
mOzHs7lZfncJFa49SWk+ni4/KW1kfPq5dsbN6p0LCEiZoagS0zlfvHPlg5+vGeEWeIuLEfElttV/
hzmzCgiWMXBKVbEf6ZS6VF9nnDld0HrncgL5LDeh3aIWFtY5QILf+WsHUIf6nCwFQITbRM9TeEMw
DkFF2r28JAPepnvEYHBAitvuv4+D5ixJHpa/91RDgteRr0SoFZwWt5h6SdkuSohK6xPrEClMkWJB
1g7rKTOT3YuqpccsOh1EcVjkTjLJDh8fQn8UBY3ALJ/d0RumxBAbFY1+NaJAR1XT0iw1r01L7XmD
/37weEWXXAuL/1U8iP3Lf1CVPep9iBd0c79eKgpvJXR7pXJ+MFHz4jsYBWQ/CIPF2VemWbfQsCNO
k/nzrPubECkpxev5kv/AGK6/pd7GsFFeO9LhfvXLivBf2+PLhGqXeJT3PyW4uiBu4erJ+ygYq7xn
0m35ZbxacqXKdkg39kmt8ncp/UXg3M94dMup5ffdIeoUgEDnALNXcJUQfO1iI4bZfaqzcg9KBmjz
loQWiHpgifPqp+1bZ2NJkS/iW2tM2NkjIOc0mrmdv/elB1Ywy/RRVF5jLZ/WBsqDbET8E44Jbwpt
z/V12bsAhd6Huxk7APIbTKiUMs4I8B33qAoh5Npf5EEjv/2pvpcVRBexQLYcZZaB56y7g/vIayVO
53YNTW7/cpJrsfZhEw4FW7YvnEnV8puQ5wftDsVL7zaxxMjC1Bm1n6wd0zOP8zDRBY4W4PCBazwh
Km7itXmN00xrURdZid9yXXNVX3lPMGikf1HptQU9VePea7cZ1RrO0gNFSL8zR4Vvhk+OKHGleZtS
WJDcLE8T7BchgPt7ipkBJCj8n1q3Pg0TerJ9X0LsJwLAGDY1BWnv1SEYiyFZjj4pQ99B7G3Adrrb
CXPwLLkXfiXajmZzpKksduvnVhX6mg84xQy3hQfxkKUdxCCLTR1h8+i+pdWxaACrxVGWN5RT74kA
IyCEtmoTgn498nZ9+VA7H8enPVRI3YN2jWiATqUrNXD9E7aEMOEc1Vo1DuBIfNe+ef3qLd0M4mQk
vhpKjAMwRp4Rkk/nHECZ3BkRfgAgxN4L2lL4Toz9Ku6xJroQr7gK46f7mZXdi75DwSngWuDnpdzh
5Z4le+3H5SStcbNXYSXgqU/LMyy72WepiLsM2TOFZ2xuqAZmsILl0POt4M8wXrh+mAYMo4TLIP44
AdO7znJ7aCAMVCaeHWZxllKJEcYbUe1B1L9MG07tRmzq8/4rJSwcMLaZzqDrGg9H9S93uIH1A1Ud
TxEoI74Lt6M4JvQsqogzXD6BfGeZDnY9Xbgc8TsKFePyzS8SIlP1v7yXfTJ+HlVAYPKJfsLFFGN2
+DOIvei+vMo2qu1dio2iXH7TtrfNOUBtmP36Szwticx53NXNp2eAHVfihtsqwIHzqZwFdXYHJsOa
Pcp/sX0aFpjZzP5eQbbGEu47mQ8nsNtDEV5oR/zXfO2QEMaeD6Q8sI0ws3obRnB5axs0UmOfX6gu
y3B9m+yDt+dwGTjBstHX1rBWgWvgcTtrMmjG1YJYt1WpbMXyz81PMM4IM+kISiZiUfkE0yN4wupB
Y/QpooyoFXrB0nnA7OOHRtxZ6Q/GxC+00DhiRFBjDdVbDh44FeEOwN8bTZPPmKBXw7NcsweE2dsJ
jXHjT/v6Kh/sFg9Xj6I8Nj6EiXYbZCWgNebBKr14qkeLt4lt076hBJ85d3LOesx9k78UUj1gElFO
cCcUtUAYV6l/452Sk28JrziGV0fuy/BVIsTej/T9oY9dP0Ni5MhMOZGb6GApUMH6Qlo4Uh33o99p
FY7t+HrXgwoVQFGQAS2rwPduDeGdh2flIA/A+MBu4Lua39KHi/ykv8JoOFBKKEY0/TZYIrOkAN3Y
jCuZDUr4DKhQDQbVZG64pFK7sGTJ2ys6D+8FE2nlR2BGRK+7KG80kMnEUY6VIWIRG7RhKhgfXfX+
TNI/CK/OeCqvJRY9GJ2xQJazwb6PXHCSpcSrBbTf7D4h/9HViZ/DB+MvuehHoZRu8AS9irDoGUUX
upjInriaOBWttw34/QOwv5SCz+qfpSoerh/1X7XbkWtidj+kzTazV0oG4b1l4rB7hg4Nobqu14ds
d/eZG62dCxR+S2FuB3kXYqhHv/XA8kmIZ4rIXvQzE4g08o19qXehICDOBYDyi2rr0Vc65fNBuFUm
DIJvyRYtp0wFZ+0ktm0UsrBwbmDWaFm8clb5/wrqFq1SnS0f0ulcTD0j/ZeFj9vQhH0PpDNY70z/
wd9LKnIoDU1P/8+ZBYamXHRwdy/tV2HUFk52t60Noivsl3pw6uKWfXVzveP9H5EWMu61g0woHlXS
exvteW6pTJ1yH9Z+loYm4AQGQbk8EbupwwD8Yx34UDZzB/+iMMZTUqCuZtXH2Eg/323ifhxFxnSR
u8xjvWwa1rsTcx961SIbYyGtKFVmLOMSahdZOkw0kQG2K8/ygIxZBiIYOmTnrNHjq79u4W3Hc7Gs
HhngYNcw+wCKZWckA2wnKckTRSajBtMqLVLdBIBQ/JrJ/3ZyRi25bpTyB0q8n9e8ZudZc/EjtqeO
xpkb2f36JBcJrKsaGDlak8XZQD89N5rEGcU0kUWcp/wKHXvS4QioOMpp9XixfBRG4Tabo2hpqDrr
fsHYS2bYLSU3fKOQV0zCW9lyNXek6idCnvrJ4uLDgYuujlFr6i8K3mKM0fIxsGwhC7W6tVAQPciC
bH95CvHDkZz8PsNp+k8FKqLu2f3aIkfGN1s2LkGeuM1ktjTHXkLrvUfb73AGF4sn7FVbjzfsC4Mv
lhmwlXXfsW+OIjn9Dx6mYFNRiZ8dB5pIudfiaBlQuaaXJrYvgactmWimFOqCM5w6wNA0wFd2oGpE
7KhsKc47rb9QJ848WtRCV/WpgFarbdY3oGcWa/iUUtZsFhRJb09IjDGNIQ1wgQA66af2ssqfpB8o
J+MSMpMJKgrG+5JMCPRCPJiGBD+Xar/0sY/NLoadPEpE2eav9NO57AvOyxiuYmYGhlxqFsTF+U+0
QTo7uXb0YrnlPjK82zXrhJyWxgDqZ84B/kOF5uI1x58DNpDHnxTH4pw+A7rJV5GTXxIa3CS5RjEL
EDEIk3bHnOz5yBs6GwxVw2hBne4nBDlTL5WlafCIXSWH5Kkv7IXJcq0aKwGMz6NjnXvwTZSul/wt
7nQCn5VB2ZtUbEZvxqkGjJSDbqlZREYEi4aIK3h408f6We+Wwua5a/3mqoqaKMWDy8Aaaaj/fOyD
IYvzIGDSxLdV3SQZEkTdM63mbZgv0SledfPpBllB8O55+dOpZp4ABpQwqAvk9RHt4IaXsW6J3Fg+
c/mX8BJz2XcvN6B6oUKHVBLvDWxQkBFdxdz1pZ89H/D9oi7MURLsymfW8zUh+LUHj6jQ6TBOTEiO
wtY52mj40+apqB0iEb70B1i4nqFEoxF6n0Hk9Xu8G1YACMMWWClko0FTg2sZ1F/GxdkUBqDkAP6y
qChlE/kWXjnz0gBFKKy0XGB5NRm3tMySjguPty2ra9/ZV4cR7ifGMqVKhr3mnCOedqxyJRqfq+8B
khzS9FdGRIQoalgsTZbvwV3e1D97VDS+bg57M/a1cQ+HyTe4oJxKq4AZClmMK0cdNgHOIFfWwfLJ
rPZJT6VrNRbUJ5Dmr6n+tBX4uS2Un3obHFPS7j5Pfs16GbH5NctbD+W1xtMHT/rPamyakgjYaKlZ
T1jav/7j8GoTlRomY+hMnZIeYvdEsp1pBk5sNBy0LElmpWYtzwBL9l2+kSevPr+kT7opa3oIR/tW
6yPT7esyruRd+pAdghxXJjdFwNqyZkVofIRIG+BSQh/iwZTr2Uw+6/NSLg2kNi03zKGCGKbfugbm
aJ/zspZ+nn53OPO7piEYb6LoyWvzTdIu6Pt9CkFdBbecGs1ArHZGhPR1E5sd67AhxcYE+yOJGGQZ
uZ+QzpnT0OQ/A7AHyANKvZ4MTW30Umn6sp3a7q8mMyydkUb4WDtaRzAY1gw7UQeda4CArBvJU4Om
x0JSDnKvbkP9yg8hfQG85ELRluOe/62fCy/5Ft/3VhzC/RrzF2D6IofvnS8izCimdLmZp9rHLUtK
9TsEerascMW7KIfta6VnVHDcU41n0g8hoGDOVTIcjYRcd3oMvl6lkIitfWrjaQH2k4SXZ1Ikbolv
7VFgfca7dzKRm3d/L+8Z9RUKCbqC9fAO56e+ph5O3CioEopFHt3iJXG2ZRITpNjNFl88NH3er4yG
PGTVCyeF+xbSijo8rZJTTcl/jcnO9JWSHricnrYgyzJ4HB9oL0PCtBPxHSSUMZpFAAzfsfbPiSpM
PJSj8OrxP7LWnrP8WYJ0aWcYx957GuakHW3HEB8D9UpSU/rLQQc+i4RGz2UcrKmG6pChBCmahv5k
CAJvGPxfUiqZvWtYGcH2ut1DLDzMGwBlcK+bkfLgAzYhxpHI4AnVbjjJjC8OpeYWAdrJipFJtv7o
B8K/ILwpCRs2BOLTmU7fDVXPxuQERwvmt2zs6PNd+RCMRVYGDkhJF5XJ55BXyqYmmBptc5SsI2Bz
eWt3RxnqUZUz8zyFXhR+DcJISHM3cAdxiGkJLyU+3nO1VD5rLCkJdg1UMeabyAVWmU+j41KHR1o8
ev5OEzGR/IBV9AR91LmueQBLgtNmZOctRlVt0Je0aqb8d4BuH6CK6Q0bKwi26qHOeBtUukun44v7
DHnyE63WPFuKsNuMilGBXgXXXRa/AfXY43WT2/cd7/H4Hjno9D8x1ZymzuHDtl808SY24/RKG4e3
t74cuj3fs/4fCkzzDowtywkVDRx8JMQxn7PBmcpPgXk1oG4JhzARGqRTE/AhCtdDQgbq3Qz0xjYi
2hvYZSW5JyHpNe7Plh5UNZmcPfRUKukRbpPyzjB2FrSESovb2mUVEhftrOzNfc/cH6Ltm2tlb8A2
oYCzs56wXz5BHDBsg74cmJvsElrqdvI4+mc+FLTPl795wJ3xe5smMNcORdGtFhM+L28u7+05LrsL
cS68nCkVxDL628MfdAmrWhjJtr8PJiKbMXm49ieqTQX4K2Soq0FR280TPsQQSsgQI+W8Z/X5ffBh
KkvZqBhwuZxfBuVGmrZbXS7Q214v4Ek+f4FG5XjLswzHxg+KXnmS4vt9sT9Sc6STWCepQvGnHo46
5o/wt2afHlY5z83sbBuO+8Q3SErUE6A69hXRAhvCUoohyqGpbW3v35qzwVi5LiVJ8MJu5hIKXvVc
VivMqnzAGxYZTeYuFWb2PvRT9utBrC5ACDWCtHyyZ4lGq6SZMnw+OlE0s8OF2HpYWYrbclKOje+U
MmdkrgGRgzSN7ImdmYit23nKpZAkDMUXvanK9GvNscvhttYMNAQt4ke5f1+AcopVRaVLYmnLU266
SqIEKLvlks/T3C4ivUpXZ5OUnXO+1A8hVk177CpEFCJlOKfHLNFP0g1Ue7YpWnXETkgVhwV8Te5u
Uqtk1WsJCN25XVv8HXjGmu0/zbmodkVBplpLrnsZBIOyXT9CFM24Twg2LV/0WeZpsqxsA2Ar5Ffz
FJO7ngapXwCtWPP+a0i037CyFY7sSXsbvFyMUoVZFS97xmgQh01MusliNO+JZpwyg1De1b1e4rXG
u/9C7cEXzwrG3GIhlxySwkgK9qf7mHQZkcAKO4FmaBhl1qNfFtUPGOOkg85pOT+/aYFPXnyKW2mz
8k+Fo6PyH7muspbbQi/fcJRXUSi5F5WE06wA1/abzsVtg5uFzATnOJOWI8ee5khqRr1NzhXmJyRL
12S64x8xXzVTxgswrdFRsxNZpq2h1H0rGS3up+n/Ajzx+CN29soBUXpLtVA0ZiMsNkJsX2zqfF1K
GMkgHlu2t5Ye78flyWi6EuzU3GizZg1QZukxHMpip/nSmqTDvHfwN3xhLvzy4YcBuW6OFcmfe3Ic
onx2ghNep5rDCTu5BZXNEcl5dee2mgsoHKO1EfQPtH/xAAJCiLmY70opZxsYZAgZrCxTlk5wf4Ze
XmqGZ4zyxlNngz6zEQSONcg0WwayNKPH5KF0hrtfYzYhfFugipXfjtLw+gWCSmGP77sAxOVDSTtV
+GhgpXg/U6/koA6G+KTfCuj03IXhSzMqccJar1kDS8C46IR97JiaLyhrS00KanbY0JhJ+3B2tmw8
qMy6Rrw2podAq8YdoSr/ERD8+94lws75PGHFBXa/arnTJ3p2Y9cJyg1hL+sk3hpT83R31LNlZoo/
gCKNDYF0GaZVaOkGPP2+EGxDrCd9LOSXLv/7XHKrsGs8XbismCot1Nx/JBbMiYHlnE9V6QzB+uTF
o4yQWhzNs9y1XajLLyw0slgxYXIHCsvAB5E0TrqcSNy2Q7taO/Sk4snGxE5m/k29DgOQeJvKwhTE
XHSupleR8hV6l7HUjyRVVilv9jJa2LaoYVpofKImYTxd0CneoHhBRdNHzroG12lG1vk3DNIrQf7Z
XH6ZAjxlweXLUD3PifrOPrS3+8TSfoqmpwY/tyvfw9LXB1C664JwYOxHo4qsrkWR3zjjObH5mbU3
kQywxFuOEvOqQMx65SDu9GC/qsu7SgBVxR4RQTOBTkLcULifOSnDrdmZBMRpZpNSyqtL+7bELmfW
JPhBn8zX7e087UHsiNqocyxLgcvEodRQLz5tdC84ePgM4nrzLpkcEHJIL1EfzVxi0veNUpDQ/OTn
hPhTFJ+7WnL/zCpuM/k8lL3gD6xgUtw0c0xkWYtwMwvK0jiS4sAQQgRAjX4/HRrCU24B5T3Uwwth
HEx+V7VcNDZ+bMNBfjw/cn7P2akdsLFhlK5ry2xNsQN+2pX4nSGGvcdfxbJ8Gl+fdCd+JH5QIMQm
QtOWMV2DBqamSzs/Pq38uSfaos/aubsyd61cjIwVQOsHjxGycE0dZE+qihVJ/ig0qNZShKqAUuiJ
SYOJGqJNuDyif9tcF0Q4j9XoHG7pJGckvHvefe/EG2Ny+bBvFO9bTeUu8Y19Z/eckuABOllwpXB9
SOYi9LqpMOgbO/vB2etS3l3Sz8FmcJMyHbrfP1hLLfZgIy22ZZtorm3bHbzYNrzs7uE+UpWGzRJC
hY6Y8TKurJlaVTHsfstiDETJ3Xg4fN0BcpxahC2dVmj+h1KU7NUxHM2iB5VERqDGL51/WNpHqLHX
vr93tnBiFLHt0LfkcUlKM4dERLB22+Rr/lllnw544LtApUOr0QQcPPoVBhmA5w/QKwZvCfFrYOh9
M+2f78uP1NIEe5OgBmqQjxuWn67R43h5FY1U9KSTCzXsQT/O0Lp9Gcz/8t/TKNrszzUtcrnmpd3G
22/dgccPt+lE1BwJ7K3MMz1oJ4QJ9TTF35vcmt6VzDnyVsLgPBIiid+jDhBaWgs/m+F2SIKyXaPW
cbJi9J/o56S0+Cko9myNjnDwUklvy2A5/gmu38s84wwpUbNBeSpFuE9ItOo/SYEKHIBf0T2zN4U1
E3sivOzcUWeU7r0lEvAzLusXLspHMbISSASVD75sWUQWX/ZS6lEwokP4T3kPUEsCMf0etvCVN+sy
SFlqSDPYdITAbnVuc77bByDUr0TJJmrpH2K8RbEVypK4GHjjgG2yVdjdi0CxBKXmh0IYolfYK+l+
iyXcuZAZTyhD+u47VTOc1TKZ+gv8IV5fhQYMaVamVEhlWcc8cySzND/yIgWsZm/lk77zTIOsOIN6
OVKZ5eS/7UgR0/4ihABRD1ED2k9augl1JyaagzQNdWYgBsOY492gNK2r9f7YfsZb3cqbMSA70h4K
ASkRnKRopgzRNogutcEfUxYjlGrJFZZ2/3QmD9c3ejUEhL2aktBPtmwwm55gL0PX4K6LDw0IGcif
YU9H/y725c4QOYULdgThMweanfFe2b1LSRrrRvqcuM3h0cqYwyHbjdXK+olQHYdyJ0B76JchThgw
uJZcX1bXfcBWR8UDOgNUUQFg4LpsJb+mVNJxa8aO8zeLh8xgmS51NRJMRZ7TmkoUMRk0SM+bc/jd
ct36FAZlFuWKs5ydb6kPRLUFy4/JJ3Xfvgm4bEwhbJw0W57K9luRA443Go2dBFJPTirRwCAXmMiC
W5oHOdiflz8iJaNHz+1L3Gayg7r7KVQrMIb5+QXlqTdPhZCNy7lbo1XEWEKCXRtncxQxxQOAPg3h
WsBRoD8DJOTxumHTA7qMKZkwCvvihMWVycr7nCTDVVx5XeLO+PuF3xXqf1ntESMLhRw1CTd7yEO5
IAUuoSMa2QrZPicIKVxUxrbH0lHwLt+fc0sx5YpeSks4xWjtH08tAPZuSmW6YTZNLZC+ZkuQ7JUZ
DVLTgtJ2I4RqEAZLEL+dNdfWxNy4j5GV9Vq2GMn1J/Gc7xSKxMr7xdW8hXbIH0R/5jcuBIhK2kMN
taS8E2sk50g40UUqnd34G6msEijA58MP3Q2ur7+OLvqfNeWzAtT6ewMQMMozME0se+Tp/lNGyfIM
5+4Lb+rE5yEi7cfaF2gaex8DkBsLb+LP2RqKtmuBKadMOwB4KkpPl8MhVkVOxuh34l40aaAD4yFs
OGrkNrcEY9ii5S0PHswTZ3GyVFCoutOz31GlJs2UbXOaQXxTqBUNyc0TTwky7m5r6uI7Bk/yE/+/
gY6ZbVhnZeZA0Nv40X0D4+PwzSFIteCCP7EU2XRH7wStzKfp63sw36aYjGr9cFzYlOTCOJqxr15V
29NsdQ5ZTNLt+5BImucKGqhc8H5AeP15Hwuc8MofmLGWQ6PD3hZu808kDAKlTBe/1PRP1sqid4xd
kYMjbcRmVkhPOY9iC71JJc6/34+1s+0DPvPfEYy/kza3XtHB/2JRK4lDBjIPDwhhKcz/3+B/8myi
rKDm5DYFmFjsTNiUzSxUFTOlOyoasvokQVCWe4VCxuXUlC/YUXZTHHciPCFcdD1x0CrB/i+bIADe
R0UtIb4lvMJnUPp66pAvYEYcIPeQnLESYv2ol0ZQmORuONQ2Ykf0AwQGgcR/zq63sSP3lh4MygmD
GTiDtiy8JgaflsdeGmwkiFvqGnPdf661vmHY20Izw4X9SKvgI2Cy4nnCZcLFhDScdVv/B0lMhCyY
TNkCJ8qwgaaOJY1WXApLBEiIvsDeIypQ/txRdEE9haXB6jIHg/t/LOLf5/y7NhroeM1keMh5JjEn
CmdHz0KOyPCZ/J9mszFiFjWst/38Ja+EpKx2vxH66bh2majXN3wVOp3qkyIwAwEFpTnlsIZl9OX+
Rj6RfqxB6PTBGbJR0f4Ncmo7QCmX0aU70OCXq7nFXm5E2VJutc+8fEJe88ktgPxqyWRN5IayJFPJ
JFOZji9eQAl0Uj3GrthI2eGjWYJu19NZ7gBMYhiLw6o5RHznPIp4bPNVG4kvcn2mCBGGikyXxUgT
0GjwPJt9pru8PgAtO0U1S2Zd1TjWv6Zshxz+ursMOfKVctblGX8PkUhNIPVZn06N9ebHbueE4/TK
p0/1fNM29zKFRJYfWIsYgEX3dqXPsClwCI5eyvmIMt17zMJ7shqWCq8Cxst8/ELccA9yqna6xsSs
RColRrCe7BeRmi4CDwNfr9N6Vx5RWeuETydp2eDulBPe7rLVoSlJ1XbdDqeI4kndmnYR+U1gdFwT
wnnsCsg5hU85e6+7b7chr9WCOZsBllojJ7Wr2Dd3bSmIC0+sJ7vvCKp5OHNLZypt/V/CoyC5xpwC
yEbrjAClPIBcigHmsYoQQvAiS489JU025XTavzs9znCfNC198MCh3bSe779EfTIOjV5Xj4rpOFY/
C59WOjQyYn9EZYs9rvgEpqFKfzUp1kbk40jy0Q8kWj/xlKbMzcUWeCwQeG1zurdG7xuNJrFSY+6c
NdDGWm69NEYPdvrzSzsxAsW2To+++I3XCUkukQRPJz6/W+xyJhtvUq38ppfLU4r7K29C/UytuzUe
zrvQpOr+RC11StTQNLwYXJ7IXBnen6C9TPRcmOguwSEMMs/kR2z+vA5FoohGWxhSMsEI7ee6ckid
u0lR7CANYkB58edP180YSSM8BByuiycHaWnOjFindsFbAX++JCAaGkW7z4pLn3MxhRHimQ97lsu2
u6zZyDXDinojI2FSzKpGcmcHMAc+Hw/dAt1OBCUkuB/o5VLsUx5LsxxGUjlbWTv00Xs3Xr/NOrx7
UvVBM/KlUwT/yEZg2L2owVOkDg3qvJLbnLL5hr9C7zf+gVh8Hro2aOpBaN0nREvCpTZsnYCj0ow7
eDdVCiMa0scp/AA4MofZWWHOFcPoviU9fKykdbDq7ud/Ia6l9Q3kfpiP+My+oBZhSP0hIFPekkQ0
lNhE3deHJ2NYrygmGlpM5zj+B7/rO1D/iRMlrSzbqOEiuApYMFEaaBmE5auBi6ttNrb6q1z5na0c
cDZN70Dq8u5r9jz2BHcxLbEibtLbmLP/pJgcrggOGeFYE8xVNLbnuDABA0XBSUKkhdCU9aOkt/vK
WV8p5eJh7uZMusZUs+3J0Df/QCjtvxcTWF4BImwtDzs0e1AbIiyGtNIJ1RR/NnnQ2NZ/DQRuyU85
Yjpgmhdb9JzCKsUxu8Qcc98hCCcIHH18zbM7YyA/8CspBp2npR24zKR+Qtqiu/RFbo/asWl1eQB9
31rlDLVe/j/eMAA1ZKoGtWtenSgtM8I83kbDShAZs+jAhOblDwHhQrA70hPTuRk+TCV22bRS+BoD
HEhBBNmQYemuMXWPd3g1DxMwIBDiXdWFCQ0iKinoMr+2Cww1RybnT77KpbPqQwP6uSQ19YNV45TK
RcyI0FHA1NIRTPVFsUSvls3ksh+/CpMjUB4gGljnHNW0TGWqMtplxn0bsjztf/s+zKiJwNU4WNIW
WGvqfY7T0t5+TV7gmv8I6i+7/8mIHaofUNcGb4qJAQ4q61GdcB638WS87m6V9WOkYdJuPDiaFR1o
CxPGTiWQsQMjtQoyKCiq8GAMwm/n6hgfNSwtFITdQ3FNVd2j4Xvjwtnrq4u+AZ2xqVd4KCt70+kl
fIrxLc9jQoOMJb4rORXKQfQCeD0lZPiS9cS1uvPlOK+Cc9mRpbCOrFhp7uLc0DhUWWFkzSkWcjvl
kKAtW+SPQ9Kp8SVW5J2SvaG4tMOJMLL3MfG5YBmQ2w4aMFPzH6VCVh/KHpqG0A1itAS+X4/lza7K
OnmcgUjNl7YKfaAibjyOIQT4iGQNCd2UeysXWaIk03+VmJaAjioTfdGbRnXGyv+0hpGShhUR6f/a
ORB6R44caiaEB3LdcTHAgFwhgsRZ9qrJX/lhK+KEFNF4ZHW3DwfSkS/KO/A4LloFgN0DDjpwk/Lq
bwzo1MTzVqFSHJ5z6TFfYzHkhu8zpqJsOcSv6v9CmgliR+nYdTJ2/HwMM5/RTWSLVicdDWh3YF6E
VxV9A4uDQPOt+VpToh9VLwH0OCAgHWx/cmGAe45o94UXnTbCPyHSj1DXXMj8C7e6aMKfI/+urz5e
d6Wj26ntkoWCc0pOoSrhztlwN7Pnnz1/YYRCocnWrTizmzUD9qcM8CcoyJbHvHAuMVdRF5BCChXP
YOfBj+s7UBorayv4thN6lwhtu8HVXS5R0oic99ANsevAlOSn380lHFsnHhrmlYSxMX/GPgTbVTpj
KJoSuBxc+lPZZpCIPogKPrZCIHb8fWxoAITa7sDwSEwpwJ+gXRBxGrcadmQUgxno06o9L2uduEvE
Lz20/q/kvSBtdPERU8NaeTpno6OJq+0FKOZoQ6LOGXOnNnGrHDbcpFrCDQxjDtO0LSK47EKMt/2Q
1YeclKZsRHgc2uXKL83fjWGzliI6oMgLD0tNmgc6NpGY9X0b+0Y7WKLAO7muqYibO/PI8LHsn/gb
5LpsYS0ED37DP2PETMFceqKt13rZo98okL4rB+cS2NAKd48GLRcNRPw/gfCvhG0VLOiuR8cH6Y1L
obnEuDx3HvPRvv3+3PbW8SytM1eMpqAviIQqHbnly1N+dKBKvyEiVzeBh0CYRn0hCRLt7/paVXuW
MDzON2Ns/+RMHMBEIKLl0Kx2Rp0OizvUexLNa3SdTWAIuxReKoqYjR1Ga53a6u4S1YlH9YpC0NpB
jGD35XoS7Eca4LdlOQpVQIz4efukiLxfiQmKkd04yPMIFAXHxJwvxZrSJeB7jYyGbT+c+f1mU5iF
yIRTnbwqb9DQA9IkdM2nFEZSTC6WHWa9HHweyBjmVep/1SBvL5TBn1sCX+pLBndtI+haLOGPYAGp
uIlt6Asjcn1I77XsuXHS5N8VHuAVP5jZII3KkR9+XCX51h2TvKKuwtG+80gT+9+x6H4ddQlZJYUt
Z6kPkzSPuOb6ygkOGkmtJyBDqkpMzxZdge3HdVDZajCwP0zdnn8bJn5d1BL80RyMM0kl0QlLl75C
mZx5XGThZwdfLv+yG20RfOfQSAal296b9TCxdnpwKs+BUkgIzZRgYCb+4vF1ZnCLPw2hpyfrNw5o
J1MVg9iT79BX1N912L1wl8Lqg6UmynJ2zLO/IHqeNE7JedBsi+dJ4tvmq9tdFDrVsV+RU8V/0+6P
C2MrT2t8kmOdxXh+8swf19iWFrGFz+npZlJbleEbXEnG3nef3Rxrqdw0ejV7XjPyZtnWMcqv2mvs
dF5x6m8XE6BUebUpOHR+k+yGpp6kiP+OAKDwBIlHnpc4EL0Zto9/9K02kXZI8xAZz3qTfV3qRhEj
jGZ4fDe2WZGePcFLBhSLf1Y2GmgM7zhEO5qwopP6qQr69amCOCQJh+R5SrPfuITTu97zjYW1cuWs
//7meDKj+zBmZBqzBpGxPs/hx2+JekqmgVHs2yPUpghBDintJnpcYx/FZUdViEX8et292iRVyzpx
4YP711Skwf8vhCFL7ABw2NI3rOTaZmry6Y6p0ICCfR2/Bi9cPrOnE3JuBNTZfAdEby2UMva6ise/
3xA1VM1UXV+EVefewK8UHq3G/guxN3uNYo58zIgFCFMmUd3MPwSP1nuschqVrNOnbtYNO2UQbPgl
Y+rRUsCiQmBQ/3fNrx3WCts8M0gDJkOGzfyg+BU6S1o3X5pqjKIK6N6XrwzNUsEqshATh2++aGuH
ID654RBXEZxTQOKaVhGo6h9nBEOKNTrtQNoEMGLoTh4PFIgiFR271poV6Pr+//oVgJfEfzyzNL6L
YfFP1jyVqlPoalPV7hwzMCXsbe/hYaOGtf8JEjeu9u73x1QrvdJKyBbJj1sZUgtMcVMroevLlDHs
hWYCDCzZJuvMh4dEqedrYpFRREs7jg6G6SJ2cnVwHnnTE6Fdt4a8rPJ/AY8MMCifQZ6suHIufRfv
ZRGorcseYbTCNPbA9JAsHAiyR8DcgvIHJv+5QEULZe6GCrjz0X76W3bUCrtA2XojLc622kAaXI3b
ZjdRJKkum/BRfGq/8HRXgNZFhOZzwUGq2N2yOFHcWeoZ2/0DwMl6iGD973j+4z5pHfJu1zwo4rYI
QAqGsXxhqQOaVWCG5OKUJm+sq7g+XuQGy1h485JrF0cQQnhRASERY1FIx1M3up3hamOxnrMX+zoh
0iJYRbzOcEbrF7aAi6N3JlgbCTRnQzfV3rbLWywspqFVPNoxgtHQM4bzBGJ4FTgnPKiQlzufFPqa
dzM5g+ovLNxGr9IdrwU44o3SfVaBuFQSuYX/690Y5N1smmY+qr0qdw3PcfmnY4NYtCrqsxHflaCd
OO0lCq0MNhxUjjQXZqQULkSp1DOf6xwLizBFpafESUyStiYMIdhPFenxJFjmEZkPMSaywlfbqi4p
lkCwQgH6TI2cZLdaqbXM+5yYpqNFFW74b9GvKPNR3ZJRJ7oIrg0cCW2PJfArS1MkrO7UysZb8Qqs
rW5TD4EM+Czr38xrO4v6i2Rmczq1q2hNH7pku/aOzyHtMhfBBkV0R2b95+vu6MojUWrXaaOj2C0r
XxxzMgKx2UqGf5GYneRTdN0GbxDiee1cduGqvehlu6tJA7Pq6+DygmrlFlB7bBjyYCq6PblXesLr
AS68kDyZsnDwobewdDkREW1RuyCXUkhvhkSgefp8BGdMmrv6CxO5Fk4++CAD2rCfr5n1CvmJ4j0U
UhK5RuhQy673jqj1DllxWihF+piMbs6r6NFGiXXKfHblCxRXSg4EDtA1T0WTfYSH8p4QR0P6kkge
UarqkCf9qtizLmSj4bimxTsP+An9bLApbRX/ICKOhYGQlfEa9yxw8uoMTYVCqK7PYP4d8i8zGPJb
nFSj0dmVlM5OflP0Iz99TCYKVp+LZKtFAjiwI4Qd0uJ7ktJgaLfaq9H0gnIeZhIgqdylJPUtTgzw
2xThCt615YoHppRCiq7R3EzdQ/aN1ANrHBKHLXU7ayM9mSiswC/bi0Nd5Th+FJe3l9M1645Jrzaw
vhSj7Xmo1zS1XtGQa0LuvIgLqQi6RehoDjcTor3aJ3rAsLS4lyYpQI2mhiYJyEOE4xZ+hA3Uxz06
iyO9Qh7F9lJVFcKWXkxcKW0Cj1WABLo1lzSuZvwv7gIHsKPdKZLLPX/PittVC9jrVKZPBL0/VLk9
M4oWR5fIrC1kKVzEfMqZr+qBOGsLRtKKeOuXLK9XjOkbN+ZJyz7wyI3Yw/G+AUIV7WgJApzhfu4/
Z+OJnhKcvNmqFmiLbw2e41BVkkD89w2CF6GE/zF9t7IMJ2Fe1+g//mYSxLQDR/y5d5v/npr+BcZD
cjR+abxJxFoQjKoLqCuoOjisJem2MaJ4NneoiJUcApDHSPYAKrhiHIMo5GoYi/lKqIA665lmVkCk
8auP/cR3mylD75eTw6vOuT+9+XHpSsrOEViHLgpCaSgR0hHmZJ0jv9pLpl5tBko1kl6cEX30ajRf
Um1mKFaUytlx8JnltoV5xI1x/YzTafRkdo5J7s/5B3INL8rQR3AOGh2yjewqJ6Aonp5bP+MPH8uw
matFdel8QX37GRyORPtqVsHfQEgfa8m/kEYoZJHKXOjyw1QuJh24xRXX8Dg4egiQk9NZMhGrPb3h
MBlvVa5jhp0in7688fR7XhdgoGPd9B05vZtAdixk21wXLrPJHtgPWUybAej6VLD8TnU2c9/IU4tW
LTZkroST6FTcHkDrettDMYggPWLgx77/E8OLM38P0eLkI1Klhzv1rDRXe0ttJFOFiPvEPj4XhtaX
m/DDxETGQQ2MrAOf0q87B3qRkSVoX+TNTfPHfFWobFUlWsNhTtghOUPtlcnvjrXlJxy1fmETx3Pd
YJ6ejZGo50gEXOhmat+YbLtRPq09y6dHSWwA+JqmwOCiEoy6+Q2oAxBC5hiJwWgO3Jmi4yEm7LVw
B63zMxm/OPB/9CqhYduUqkaSR7Ze9t+agMHY9SUUEgnEXjN+g+VHWO9EwZWtalTjO/Dv5fQ3i5Zr
g/wvewLrdd/9kGRw+X1pyUmoo4IquzSX/VCygB2YHTNdR8tlYGuMpt4Dh8gQ3FBS+vedL4MGg5Cd
k6jLlSaPwgfaIVHUmCD6OdyQRWq7H1Qqe5T6Hp3ERWSdfpRg5/EmbdRaF4oexpbziLv6CNn97lpL
PfVyl8ap2CwSrkFBOWoRxnSsZIgiDzKmSpRUd+SdyTzKsWVeNjY2pWtKli4vuyR4T41LpTfzeNES
Wi3C9ZjZpDQIpppo7A82P9dYdhGW1G1nCFgZsbp7+nNX8FsDXPNU5qrINUZEFF7FUyOigjwHb54F
cV6Mwq26KiW6VaFUNThxLDAVtxwb8316qxvJCw65YBTL3BC962ED2+GR8CeO3uVumgiH7i9S4atU
my+ICyTEDWoRtVOuhG9j90+KaP5WOY4k9b/0J2qMf30qbvOJDZYd+rGyERj4i0IicPVI0OGUjfZe
XkodvwMgTGla+lilg9YsnHfnhq1uNLUqWLDyplA4i/kSD/BNPoua5uVJ/8E45W4mRdyD8/vAKSEm
U3nela0avoRlai90TxnJPvGjt4pYBbsWJMAKsV+2yeL99qAL9/QYfSu1thLSJVQR01QBd+v+HkRm
4xKwS2a2cyy6y9c2nwMZdCXaaSwDLNwKqshHiht6GxXGa+N2xKEA1gI5QvRRGIcsjrxtIrbPxiAH
vs3odfsehCloV1JQjuPOFlwqNCmxduXyHjT0m81BBibHbyeTeyoMuOncMfhnnGQ1gHqkDB4vPpa0
CfcIriYzq7KAxFf70csiBf8Bw7V1kLwzaY9XJNLN0opAsaU9hlz4BOhlJCamDe9Z2RUOgVIgivlG
XkgYO8yEsEuwYCOXf6wP0nXij6B2raq3sur9BbMUcdlME6ERlB2MtCMyxHK5KLaNM/IWwWexJLZE
BLuvq14jyltmf3wBX5m7HcsVPpLicZJ2InbQxmJsPcMSSuptngLvwn+HC9FFqMupm+ii1ZwdKDXl
D1OOiYaWUc7uM7fbnsaCeIOyiLJZK2w3Rf3QZtxZidnIyQeGArH/UfW/VxUk1YtNVRYNSw6YPtmO
5pxWQBfz6adHQshptxfrf3c1cmKXjccyunFdByMKDNexADjCDoTTxUpJSAWzhnmtTo3gMzseBgZQ
1BHfg8nJZf1ZImzMRNAEN7GJQJaQNVvtMCm4azSYIU7LHZc1GIPwe+MVHpMfNAqj6LOb9SDrDDQm
rhjF7SFPi9vWB7AovyiFhjns9UgLrDsdUXog/8r5+10OntWrcyxY/VpY2Ec2HbB2vzhqlCxKGxx8
qNfhzXbleqPFBbNMfCNZSqL2aaJBlRij9CyWRfdrxrv97WI7bhgyL0MNsQNUxDCOkwGGaQjVBuMS
Cqfi5Mem/LLzJNVwemAEYHTiTgVcIZyjQN/nNoDQhPRkwjvHOXaMbtxvtDUV4GeUltb/vrn9iQwg
Q7SMd2sblRAKI/yH9f+8qCKEltaAs6lW2qP8KdE+RWqqSKn18PsT7iwraLpqve3CCRR8GGDYdbWM
VTVYkSsE06stSaeofV4e+isMI6aFMRO3tg8vPWAMVQSBxZxYLEIt/z1CNLGZyuZVfkWmX1WBdHXr
BzyFc8aRhVmBvhGQKr6GrXoDgO9jYgALWAe5h73AzbtPMuQp/Wd2sm1oaExNaFAW/QMxVVyUehF0
b9Lny3qSbvlyhd32cXJMII9L7wI7p+sMj6rAgayz57jQg4A+RclvWhZQqZmh/nupHBQxJq++CTsy
BzGfiGC1KB0jERrGFW4KRZ4ZOqFp7DFvwEVB9aMHxkt07l+Hs9Bk2WqW5xM2ciEYQ7iavR8uiAOV
vYw0K6wsWdFTqgUfB4cLSkdP8WbEgK7WgqNtmjVd7xxhPHyGZAiLCaRcUJH9ADoyC+U7bwc8y7AC
4yGk5tyybHsWWNzx4qoJxYfd+YKKKJR/N/rPokRUs3/lEM/xdWIOXJKab73TDhsybMxLzt2a76h+
r/FdNUg0vVhcO4sHs8xy66oIFeEhnjJyzNRYiawmsbPOwYUThHkugQK7KtSI4wLhKBpWMuN5Wjbr
3TDbVL7pQfnr3j/pEm1GvaG0Cy2R1oZcAdIRrVYTi1iG4FX3e30Q+NGGfSrP8YK6HYGDgKUlRcfx
AvCFVzx9PpVqIWLlXKGFnm9hTJl6YcYFNYnVSwESTL+u0wmKaUDe2PrxFGZdhftmI8Gs888R5z2s
08qtJ5nQ9+5nzoKwT6AFm1FUitKXSxyO6k6mocGHUVFmOtBI73nF4DWLJR/Ae8ex8aXhzVzZIdwX
KvyLGFM0aDcpfFIy6LcAHBg5K7B5FEP+53nR37XOzZXf6AFJOS48PULSIBh/rRLAMe30YY0R17ht
15KQzw1btQ2/zbAktRY7Z//8uFYuUJ7K6HVB4V6Kb6uIv5wGEhdqV6CmroJ144jgO3JZH6RrmzFW
k2Hk5Cj+NCGdnxIJZIun0HVJ87ye4ZNQg1nGc2qwUarrquRhl9fuLDPjY8tFSiyO6jYSACZiqvsb
1GVltsnt19xUWA5VL+6pKSYm+J2TWcSo5DsqkmEMUBeWuEICLa46xZj5BjN44CqoYLwkBZAMZzoV
F/yzYSaG486aSZhFo6IZEK+L64xMgARY/ykKf0+QwX4bzTP4g4w10SMWrnT+oWGGLr1jeGILNsKR
71U7IC/An7WHKZ09hV8aoT89rJj9Qc7j3nw4+cKqPVSL/vyy2/fn4Pl68y8jab3cQObjI+wXAyiV
MDER+OgnbnYmzlc7eZ1jFXk/A8O7UoKJpNtq2vgYIBH6Umxop9PV9exvsfkU4iK6xFSG8e32zYkz
XRmzhy5ZdzZO8qj/c97Qk/pYTKcRPENpmWRbos2AEqQHpUFStt7mjZJ9NyFmZEuSX7ejJPLXnRre
s11XrP0/mOoc5UdS+FkcAVwsaXRez8/abmj2uCbq7ph4QpykXvbQJtqirFojLvV2ZJ4Y13bFdRrV
y3NFQ3dADdzxzEC3QtHQIWHL9cZNtQEyPhxk9p1zPOvxt7D8Qn1cYE8YiOBxCDj1++9Yai//U1Wo
oVTpwfZmuKzNBzSa0ZrKd/lcNbSNMniRCSLPLvDRbIjvWU+IwIlHi78vVZ04T6MjN9/Fgl2qJTuD
Gd5tiP9J/AG3ikAmn6671Rg5I9edhajE9uPL+D7XgiqIxlw/6anKGMt/f8k57wmg3+fEuJEBRjsi
xAwEXvmpnGpQ0QLrYVxv6hCknxyEFCNwwiqh5sN+hgm9DHFijGXsP5LVzDges3DuzL2Rq7sg6NCR
9ciATAtlYYrYNxERcOf77YB78p6kiLavdIDY4C7BQRYasGo31BpFPcILiRFaHGAtfy0GLzEhbXMR
LxNx084+rhP6g1VN4XXUh3+hipI3dHAaA+7gdgUSNbbhub/9ewRs1T2wfqDHi7NLSxrhAs5jJ9MN
d4STLhp06FlxdXpkMoVSs7Kc3e87loTNpWdBr2mB9KQMx5e9BK2SgsEEHBSqrIR23eMzHKOSRQ26
i/7BhQ8PydJ4WPg5ufH4Pw2fpUtz+5Di/IJX+IUhvgCn/6JokYqnJkbgY+u+nQ7VjBYFOCDNE8aB
PIFXVaKuE7d+lnkG6fIe293IgSUqJIegWEjGUCDIu7v3Mb7bpL+p4BM9TqxbWe7KROmxAi7yhbar
taO0jMR+4nX0u3jP8TfJknB0cGnt/WSOyqlsOsu/wPhTjqozwYMabWIVGTRS1vAW2HipLu9HjB1A
IbllCRxfOIHJM3/e/9C5wbGWrsD73qoWVvvtR08eB3dlgmYtXN97rLUp9AOs3l/CBp+PEQCk8eGv
A+0IDORlQIWE8ecGxHCYw7FyMii8ztPDOrNmPXO4w5WP32sTeljvQqcVu/XNfvR8Rzk4PHOvJBh2
VONBpZierXYbAzS/7RsifbxNOdE9EP4pszFVBT6XGd+eAG+UFwcgcG3/lYMBLe9s9oOPvFQlSddO
UGsUVGcKsgq0Gx7KHKYJzzSO3/ATgH5TVwjA77ec5bUatsf+fd8q6sR91usjWTQgphE9aaBhbb11
PyJp2JuFaPIyhL2RFzNciuOkVx9gTCVupsHeFsSqdaFJ5ZYqhwVbzVBXWqAlAMM5A2TifgKOrzp/
Y/gL3NQgRJ4g2JIE+PTJXD/yj4WOSjS7+akee+08rs4AWdE7ponqBbe8SViKuHnDB9aCxFlS9Z/e
FIkpB4oE9JxUZRYdHKQ7/8yoUyGDlal6UkqfkmljBQrIkktkm8U70e8LhSqdu0u+b7cDwk1ACSQD
HjO7wH8DSZu+iTWbGm06e+09kjHbWGjwZtxQoJaO6NzT7FxR+2uC0OZYEHIvRq+DOOtrubAbZ2Ig
m46RAZle3DuwF/oERSJsB/2alv13NqT3cfjg32BzxJX8UoiVAhk5USf7kpQ2HgDjTYjTljv0shTY
NVroOviLSCnFlAbPIIVcyajYEgOHxNDhZ24FuXBe5lTF9XXnKysdkBvUHUjVzoZf8Vbk2X5eQ56k
JTLXlS746IS2piZUL6fgndbwGxMuHIGL2SIjFE68OsHPgtbAbl/LTF0DL7c/PQOxhIOWFBZPajAq
ejtSMv4DVucJxWoEOgulxGYyy/z0fp5We4sZsTfqSLknMtj5VI0gfhNnTQaVwiNHjdQZPAwIX9Z6
suHiExhhM1ySTCUbF68nrj9afOR1CieWsXQJ3scIQQeRcsddLyz31xLmXg2HNVfHA7kXTeR3WWBs
OeZHB4lymSETUx7joF9WPttDmdhtcQ3D5XQ/rsP7KsWYDOWCrHIlxTgID6tNiSoShq25uHF1nAs+
eLBcFGRgpcFY6b4Vh0/Dyibx4onFFYNIG/HT0UQ5gSQJbIBikBZk44zBYQv5+9JJN4WgEAdMMbS5
jgRziO7szmAV8ds6iHLeNmk5aPq8v4G0IkpWKOM3Bsfw5IX/9jBpcinf3RBRHsdwhiYIBkeGAaJH
rMOXPysn6n1Opz51WW4osm0bKSVPBWAXmNV2UBZTkyMwBWoxlZAd8hS5jhAnYJheqo+ooiaKtEef
E12JjcaQcJk35n2xZ0LeP8GT1ULwpxU/KqZa2zjvio/gTsF+KqrJdgv7t4/WF48DqxFe8adfqlFD
HDkr7YnhSAvxXlBLCX9V+ushWhcqvM44Vpc/TJwgWSowpmU9i0NN6/N9KBsdSjjy1+r78kg3zGKS
yZ3MgAJhrhJlKb3Oo17GIxTZuclwtzsZ7/cTMUJmcSXQh8MVQgAghzyBJns7UJZPfJ7rPBacNz77
py1Gy2/wQLZO+cp9fJhKH7lpbUtRAvmv5aeleRI0IcG/89bzZ4jiPllvgMDPpzpSRJh1IrBfcJTs
SG0xhYL9k/cPhnuogWKcERkO1h53ocJ1D315/fCWLAszkOMEWaxOF3jUOxrCHMH2YJj0wf3hLEY0
Kc95y4q4/1/oJTJZADT9oxifj3o+Eacx1lkJrzFUAHncmwyfxORLrP8bbDny60LJcpxBgvKKNfv5
l+ldmPHn6q1wpI4GmF1gj3uyruPxm3qaCq/lMALN4+hLUZgWXH5XyfcCSPeZ1diYRuPKoBr3e9hX
3diFXkfvXbF3EpLOJ9txkoEbXk6CO5Cd10LB/pOmXyVOJ/SaYn7Agt7X2k6MQNEZwV1ci9Yly0DL
pMx6LmlPiP9094jfgSTm1MlPS+lemNLdTTESrSHIZ2dGLSQg7jyF/2xhsVdx0ztEsHgZYHdAO2Nf
+bdfgYbvipkZN8DjrGh/MG8SGcB3pJs/VutVZo8uLLm6W0uDfnSb98LdApg+mTrnslu6K+pdBjBo
0RHLmIrLi8oJiqSBMcBiXCV4+Sa2CqDcCHHBwBbRemfQzMlBMx//Obxgf+Cje0kKW3JfBn9Nv3qq
Nv2nd2U3K3sw05Mput3piGil+kFUFVR9IdBlVQyybNr0QBq54DxcYIFDcnKG43A401FmGN1qvige
W95Kxsvn8BNP0S6ITrDMvJlDxZpLkORkaD12vr4xvYj9JyIecLJ3Qp3up79ooGfBIkRnPivEB/W/
hpyALgWA5ycvwvyTahb1MQHuf+pAiQ3Ie1yE1xf+Qv5EmuFEOMTDQozGombxEP0bJI3/2uzlUKid
4nFxog1J8Y+++jD9s5UU9IOlFokH9tbSfCDqGICiMLLiDy4jxHKexDduU0BA3IQ8NZ8JXeUEYbMW
c1Cfk7ymRlghd0YXHo+4vdM2xUH0QWv8PYlabyFiUYiC0iimEcj6X1Qp2BQTMF0v+xd1XeS05RxG
ybgbY2vwiTSkF0rweZNmW4M4hBq8wIslQvO0hm/YKWSSxV/SvbCgo4UML6882dwB0kuqcdSj214k
WfSfKuK0B6aZZZ7nNPORBLOIxq/kdSN0ITwxY0RpX9OMfbqYKSOMqRgbv00eLu5JgsqFaLdn38fl
QPwNSlFU0PFbIu0j/43suwYcu7rlp2eUQUauvGoiswehXlPnis517SZqHSA1Im/tdxBuya0HLIGY
zpbI2pC+bVh7nrywjjfiORctqe/U6me6GqnbSHANau0Pdogh28z5t2H77DHllnLFqPhVHBqH4GNv
QPEA2XLz0CVknE2BQ400Q4aj1ORXdD2uPxj//OEgvVMFDDN/nkOFMjkSBZGPA91VKIk9gHZJXG9M
E6sYFpfG+gVqE1utuO1xcWT9l44P5J+jWhXfe7XgEAX+nBFvrgZC346iSPi0CrdIkMseiYzgzmaU
DmSIJAaSeu4Zt1PesqKnlf7mHbyWdRqkTkA4DrD8ykyFA8n+Zhe1WDsw/eoM+mFQk7ecxAOHG3FL
0dXBdcAaHYq4pjwA6wLad/IE5yt/7RpbHFel/OL3e46p1AwfyKt/yDZL3ycwbdpMUUw0fVW0SSTu
aNYw5YaLA8nj/pWsAkbRxs7c4e7u94XRMUpCAxFc7M5Iw/WR5XOpZLZgkRkbjmwPd+5BT9mg/5Oo
Zm1pysC0ufTyOuep1fusNMYF4p8kmELJHbo1GBD7j+iUG2lC8O+SeuwjEFilI5FPVTesR2AI2LMz
KZ3n+DMvKvKnJ1WwhrMRgVogoTKJZa65hjwSyagHBeqqONP0qQQiKoHiOHYLlGeOqWNaw5/QL32N
24XRI9issEP93QxBWIwIawPOWcbH9jqvaL7YLhHUzn+vhCzuR97u8FWEeMgDaDhLLCYJ+Ocd448v
I7lgkXaREYFFwLFzzBWF7SBjGvONJUQTkajfbxOqNg0YVpuMPkAvNfkRla7pcrPoOsQGyVb7txx2
f7WO4HJDGflkM2i3C5fcq0JPJv+2zVzVHiVHXi1f7ByNVRx+UPeUhKRNeovqFuwI444DZsVp9TBR
ETZaKXdC22IukR9iDTbyofFmefdQzNSFIlwzY10pOijpCbXNaJLj7emBIFbXt99LVddsQjnJEFBE
luqrCLSJvBD4/uQtPuE8JFtQFdQXb0Xg8NrrrVzNEDTzLIU5cGRBJIHogS9sTn0P7z4a3J74hcSX
NdnCjkTNhUW1VjY/psMLtTQyj1i/i/5oCdYVOmr5YFTENnzIFsa2VNyStR7AHCKbzbx/yU+m6O0u
zYWZmc4PDXx4oBf/AfjGek3bd8ngZflluKzZoAW/LMKCHXZrJ5k+43OiB8xxn+1ksjDpCOZHqRzY
7EWvxCPZaa9DNNOrgEcMObTWfdVgWHP9gqdpXGJq0hvRmAHl75XfIqDCWQV1bedyWCAdf7mWbov8
lCOd8hJ61OSdkqRxswIXa8aCxs5JWoIkPW7TG9e+cHuLAFdOG28tHAwrhd0zj9T/QZ4rBrviw+Qq
RuPXNm8C24gFy99mInsd3aWGLuaQbq65q6aQUhE9S9Frg9+qgIOhME+Ud7h7yhwtNwsCUNolrKAP
bg5HYv8Xu+OmRwXejypirHq2NbdO5I/Ejm1ay5RmUCjp6qP5wI65YGkZmCu6I4o0jZO1DCa/ZpMs
dauxxIh885y+7zc4+nsVMMg91cbuC/VGGu5k68QESKcGei9UysTmJRBFxsNiXVERS8h6w4LSnGtB
ZXYTqiWtAFbNidacCfKMONX4UYR7Q9DYVinrjFO10ftgM/gFUbMxH9qRGQ5WqezrutUVsi1EQcju
scfYcoM65phCikpDIJJOhcegC6SjWqh75BCBOS2qcEL8xEZBvszUPGwRT7YvG80xO0UQRM6PQ1w8
NQp38sP1qyZ5m/Kv5rZpUy3UOzhrQlnfPH5/IsaCyI6uJGumnbzFHQdM2R0TQkESYtJbY+ZkGoi9
w8xcOq+/s4z2uGEhM+Zv8BW5w48BM5/tyeEIMde7YFYU8lISSlPyOwi2SoTOABg+fs3izxmFMNVY
jVM2xESHeyk8j4CiLkNMAc3M9i4viVSd9/ZpmFJ1+JigqzfStRIuCZnvSLbS9gwu2eCIqLqOnFpM
0CS8Lk2Y/wsBWUsC7FpNe6vUPN1fO0aAxNzvMo1wa5UE4kfzJJTT7dYeTOJyoWQvxeuB6m7w1WBP
lpVpIyUT6tJqpwXSbS45X/uu6W134D5T+FHnmOy05WPFJhMnYdXhcOpwcFKXPI6zkYmbyrhVQDAS
JF7SoKxCbfLMhAWFm3zbhfd4yZpt3GxWWUYbrGLr8AeHhjlG4AQACZHB0kd6rc6nQJs03purvPlg
EvweAo0nX8mv69ZucuHy6Sw1R6zjLRDUxjGvFEs3IzBtHQazLqB1/midsqYCeSvr0ucI01JLMq9I
uOndPPncLnnZUE5oyvqL8zgkFRLy8sqFDty1qnPcya6p+wXO6E8Z7LxGqJ4SkUSpXfw2RcdaWwBI
AZUsLqO1iVNLP7PQfId8zCxoKP8f/Cjopaq+aUlRvLrJFv+0aqEOrhuXK/Zng52QCVb3DmOpELJn
KwcH4cE0Bj6sMxi6fHsJB6yLdFBVZoXZdUyCNTPHx+EF/e5FyUI8OaEUqSvJa3MixKbBtffao4Hl
9gHGJGl8pLuMpkf3ldK07u9QA1m19DKdk67FNAs9tm5F+9pFE+w4co2OwwCYrxMpMt5uCm3lGqAJ
oEsKK9mSXAYrV7BIZfS/IzCd/INHuc/2b3ck/fgPEcWi+ibQmpfzElO9CdWYuWmUbeXKQbU3RRfw
TCAFzI77YuowIqwjDrukQYlrs2e9VB2EWK7a559kVVRzrTeI7fwx5v6vGEaR92jQ0Autw51QG0jH
i4Rh+9MhPjuksvX99NaC8WspKChpwi3C8ei6lv/wx3DAN53ZGZLJGgBJ56xv98vo0gj0YTcCrVv9
AWCeKtZTSmIB1qtZvjPZOwBtIkcrOr+6+bWi0IE2DiEphtFXlxWx5ZvC+h8sp3XVyJ2Uz7cAvKlv
3uycnspcgBP8tsLJYGon3qMoVeJqUKhlglxYKDnNaiTOvnbRwH5XglPcSiaJlP3F2qbQG5NCyKLe
lJ6BHW7r72icfIYe62FnMOwTz1R0EbEOLM7kMqedgYJH4Cb72lwvthX2xWL/3GsVr6VumLXjsFB1
630M3PVVTUJV6z0h3CShmTxTZe06ElQbNZeKNbW9vB0hTVLmZ1KwfDNlb9a8t3Q2J//jj0IcEQd1
VD7stGdIFL47Qq8N7fH9rcXtKAmIcq0fcPwY79j06BRx5i28Vq860+CCr4L0pJvOKT7VeiIe5p59
Y28hRRIRO7bEuG3HLbDcYaYp24FKzt6EVuaU/sPzX6PlgKwMGcJ/rYoHGJ1ai82mMFN3qj9CH2dt
zE49zeICtJPybuJTZ+9hOS5IkztBer5VQg+zgmtkW4lL6VFg6JTiQiTE02Rc5O121FU2/31jUVnV
bVMMP1Jxq0Bq4cs4gzVZUalE7W2MVbJoluW3bDm0vZMKsmf17QEjhVQ5QDF/lzgXEYqXEwt5GBjs
jcJRq8s+whmwV12ioaWE+JBNlGX1AhMPY6I+sSPtb/Z4obcEkRnTME5D23j8/gLT7HFDs5Wm14RO
xBnm/fwVSbUuKa6V81xqQg9vZUEBOg04VD59e31QWKlC0S3Qld8y/Cy1VoyeOLvc3Mh404iXiZG7
nITnWN58V+iXooS8M543ADcjRgwMlQld2DHMoadygYh78B3gnZcv+1y61SJuzQU1iWv+E1JKwx5j
fxfybcEv++B5sCetCRTn5XCs5fMR4nXhQTz6KUJQgG1KI8JNQVnrOt+WOoWTa4ykv4A5IFbMqxN5
7pULf+waKMCNuL6U2wbzE0owR4SNgYieDB6+yZIozAPnWSB0PGY9hoY7H2nG0BJNhYeFgLoxFbMJ
OZ1DJgM7tN/HhDmC/D8gxOSWU1+iRVVd5PTN+XzLeKxP8Vlw3Qm69/VugqjhqodLEfbLREAsv2rG
WaOhlG4H142jZPvzrBrjX+D/wh72ApNced3l250Oq4K9i76yuYzjftAqu+rT/4uxx229Ug9/jrGA
7ZK3e0IGdqjfSmb7dQnw2o2+Yq4Fuwg3P0b6Aay6pxBNhZ4KXER1h241qv0VpQZi/zIC/WRYJ386
oMdT3NxC2CSoriPF8KpEvIxLHkliCQoko3UkVFVpPiMlT0NZZ8tbm7owt1AXDond3yHJsgtYeuZl
KtzhEhwAMptsEyNL/MCe7zKQYY4jxWFrfqUJHid4sh3HXTcioADGzredW1QLPIevMVioMfoihZLl
7JJPDn0nrvABPDGcEcBkPHFkEJspj2hwxnvZOppEbdsmwGQQkIBrytjLoJYAMV4KHK9Dqe81rWqM
4vIHVci/I4PQX9H2oCfpqFHdHoXFVESnfU8GcRr8x9AHtReu+OFjOOpytp+Hp+gaCtdpAgRqDZVq
UdQXCNDNqL1NPGkwe83UxmFBZ5iWP/1YcQX4wD2c9p6E1SqocgtY+xCKJEH2+8LETYCbfUN3Sfh6
nhpJVGOUn3JhNl9N08I0HEGCCZBYq5AAvt08Xd2hpa7P8W7Jrs4ZrgSKO7wuboV93X5gYlAQPcbb
tlkDqSYJR/mzhizB703l6iRpXLgYcPM2ng6lD9hLMLPhMFUgmVU0dHG1d2w6i2o4K6HdmBnBq4uB
exdFiUFKBZ5CyduRizqjQspR2BqbIZvJjUZ8j/Qkxv87REsHvsKlm9XIJsCABbRVP3I+pwAGmds7
y+aY74MZN0qjfUwmdsHM3pmgv0ZwAx/PQNV6+Dgjm1yS01v/lxje5Qja+s53c1KuKfZ+MTkwl3oe
H4El39YBv/Eg3oZZyXmlA9SP9ulK+FFuiwareXtTnhCHc1xMY+w9Wf34/sAt6JOJoxn2Dwz5BhS4
hFze6NVbcS9ubptOQPaeVh4zLrbDUO3rn1p6L7sOF7Ns0S0qvNgYCW50/26+9v7+fu0f7Hrckp7D
MAB7loqhq1VdlcZs5CEW0ixGI8jAcuzmErmOUxXgpL7yERF1YNlCr5juRNVTt5rF2W9oVVdCiGvm
Wh+/Qw3DLLy9RGZ3Wo9zIgqYSsWt2DF/jomT791NFimHVsqHAVBXy/YAS5t3O2FhYu8lRM0OnSXC
vYo0Lql5S8VOADdeLfL+D+JPZ3x0WvtiynK9fsjkb9iAYTKNw8qyKTK4OoNOSC7o7z8TT9NS0pPA
tuoPqlOhcJ5NEmLvjXWp0okDSG8UsypEUp+AQVPnsotfm7B9ZAuC4S2xRDkPQUtPAxnVicpHMxr/
TKXSgwo5X36/MTplk0qcb8Rp0bw2VVxMXPaZOf4j61v9vYN8g2prU/xzCO72z+hnMTMOpCaIt+Qw
iVZrGfHt2a4OmM//p+Oa+0Un2dnbV2hNcjnGkxo7LeYwBuqIWEhWiH9CGJvJYcl5DI6qWw8pBKrw
I+laGNe+luedD1woEBbUxGBQ3QwoD1GLSFptjOqZiy1hyjU/U5E5SzQO+uotPTKohW3o3UpUNG9J
Xexj1A+8w0GV9vbtMKryKl90S7blWuYApAqm6r212y/PCVtJKV3Qg6PMHiiQ9FBS0gGFgwU3+ETw
oWCn6G/xKs24TJb7xR/UaxxZ3+2X0jf5pMA6ulvKlQv/gRlE0J5QOf70lE9VqgBkDHOVABf7Po7X
fFtNHT1Df4MeQSTFX4FOXYbeCXNfGi2fJMXIibVHSsD2F8eaROhy1mooRxth2TuAUBufwXxfo2E6
LPjIYqWOit8SnvjaZfl+sLO7ZKNVuyW8KUYZ4eadKVg1siPO/hAmPMUQ7hc6AE/WhW9wrycMghUA
NnkRsoTSHg6iZu5/pKuwnz3YMw0RVg0lzp0aAiMJnbh9xYnGc6qn8UQVMArUnkc5g4dIlyLCTGW8
8dcF1TC+thZGiydL9t0E+0yUImRu9QE9BqGnxItc87mJXShjekh9nEY8v/EcOKo9LTB+okYibkBN
e7oPmGo1Obic+zGtUBIphXoEUAykqM4dVHqG/n7HzyT6nYgiKGQn9hGgeQ2NhntKpU+RxM0t3GQs
KE1WAH49iE93Po+A4lp2ZDWjtKaG9Comh5M4j1m8tXl+/DQ8r0YiuGEqcn4SIkRpuTKKrM8fksgr
nloBqJ2WRgEL+JDTlpyux69AxlXyCYyLm1xzPOdFc1wX4v7tasR1+i6XhYtSRoiv42hqf6uKAmx1
SaDP7PkD5vPFI5VZNcNaezUs6cMSBwuYIRLQMkAzcpgt4T+DgQNw4gPeKTR96lE8QYYzJk9mTojl
VZlUkpzkYDo6ZkUcBqayN4UftTag3vwHdjRSLO5yFQSCAI6N9GtXQq0QtEGOhuqt2kOaTll4mvU3
mFcQOxnRetzDfmo0NanXnohYDhkpcAoSzz8Ttc3QUoGDGFssfmWKsAstplZpPgv8vaDuWZG6+tPw
E26JBIekcegwo3Vq+U0inU59cTCoktJcxVS63M4WZWw1E7wSHAOQ6Q9oBczqrsW/kxVLUO4yDBqO
Q43dxqI0Z4uppvt/Fusu8QA0ygnGXQJ42dL+vgNAifcQ73m8zII89i5SI/ykYwmOVy71GrN3dUfJ
bWOQkhi1v/oeZFt6Nd2lggfxlbgTsbqcvBRqnFz7VfDMPGY0SgTTJQWcG60OJEJNw6l8ALVPn5yx
zm55jymYkTK24MfjNNZeA3+31tA96+HWST9b2czGCL5XHo/ve8Hv4azfRrBJ6739fWaFnYLSziRO
grnYNdyB+XGzaoagwQcf5Xbc0Sr9XzDfZHJzzuwNVJm4E2aM7atF+3yWvXjHepxFbIMkkgxD6+aK
fBeASS/v0R6pdf+MTv6QdkHaEd0f+1YhzzUe8gs77SdU6fjE6C4UvOOJ0RNr6W3wBuSQgE+qTCnj
PVvjUn2Ce0t9H7ABsUiwA5MoC0fglfrPPqKfN5dvBqdNdCsYZb5KmGRAP/LVrfBmoa2bxup+73v0
vwyKA9qmI/9KrJ/k4RYTibTpbehw3M1QEguY0fRD/I48jRFKPNr3kKNgGYW48l8V3vTuU+EfV0SL
HTEo7CI3RP5Ri0n0n6rlhL/ItbrFStd7TgQJBDUmoYUAoAMJaSkMSKsTzoWono451UU+d0gsadnq
41izxIS6X4KtjVHlgHzVP0Qcm8M4HjA22wvwMY1mwmGgVbbHGUgO6uQ9M4+mwY+FlhXOCpDsy8Ya
Q6eKT7SLPcPQaSv3kYl4dqphug90l3uWzB5Epld0F97ePaJQrWZAnfJKZha/9gFgeH39htvR/5gQ
HfLoxdfEDT0PBbx9i0xi0OUFfrUj2bn2N5uBAvVmJN1lhjviyGd3/EuEK/uFBOayE6yQ/ArU9Tv9
qurAw+v8dAG5itOOoFl8C4GdpoygX/QV61/rXZMpld1tGGUBsKoYp/znctq6xDtB8Z8qRTon3LAm
k1+GHG82tYYPZLVreCLtrv+vB0KpYzxXoKlo+eqWr4A7wrpne732yMf+IoXuHTilNT5fjnV0wE7O
QGM7z71s4dN+NvyAgTe0t2cYStYe5cfT5YAgxrrvu70KxA7qlgoGnlXuVxMmySni5D8Pmbrgmx5B
Yl4Y2GljnqL7sQaC+TUDzXSIqzlHBB8z9U72brQnhNTfCc2nOlcwznnXu/ulqsS+y/Zrnn87UiWl
dCtUS/eD6Ju8zv02q4ehDsX902At/L9jwyq0ZxBfVrzq5CfAtv3y4FAW2T72Infqz3QhYW8oSd50
Wk7P6bDukc7JhUOp2XwXJlsA0qW4zNfYU37Ia1rvVtIHMW3tjYeCtN6HNoNU5LYliAL/pMkfhGMB
EfetAwfVA+ugXW5bSJDUG65uUtyZPMObujxZFWgm2GaqfPNbSrchhCi59zA5cnOSfhTeS8sE4PTR
huM1aTB4RoNo/GWPN7atiqTAP7LVc2bXakQ2ZrahDUzVsKUChSQj3tp40NjEnIPrhL+Y/p8/aOTo
3fLlHF8MVcHqqSZNamI5JY7r0GR241zjgM/u9pjbrlrqIjCu/llDR46kOnwBquaM8qIi5Crv6wpC
8YMcrSUTMFosa45WPUqlGLuHULw+lh/G9sgK2kcUjK/OmtL1EM1XGkUOYzVMKdcC174+2xeo6STL
3q2PHYaq+rWc8KOn/ZyrIQdcYMSjxJBmtIytoC/nmo4Itg4sz8Y2ptFfE2bd296xF3EAuH72W3/p
COaNum/+3x43jmmFncQE+1p3r92U3gGWNHuv7ZdO2J0XjhuE7HqusgiHZVSvQ7Y+OepPo0szjt6J
XEvE98hdKW27/VJt/r+mQOZyYTsm8HPgl9UEqC2HJOsbngcWPq45M5h7XXxZB0QZLOAOptFcTMzx
CwX3btiL8tyOT/gh5qac4ZkyZqfsZ4GOnHuecC7mRSaAQTfWdbQcglGaaK4hdaeae6725RNz2Pjt
E+Srg3H7/w/M4T8ukF2viVTykb7pGAtAUMNrCug0kBzh6gVFoB3uOuoLbdaIFAXYRzpi2q2Oouap
1STcgmOp9Ij7rGCDL3JfQrKw7Q97rOo/CI6oTM0PEI+d0Rn0BRu5+jZDjUc3EO24BWApsKwtWFul
g3JPOXwt7jF31J3v2h+0ISRe2W2sVoUoED9PWQI2c7p44WxwZqur2g/W0N+7o4orxXJl5l32ZNKz
YdJcJljHRYrmM/KFzFS9LUSiconKb2VP3eiQZgcQDP6IVuezTx4XcleDn2rtFcJE84IZlLzNUf8Z
QucpOmxxD9eKk0QpRLfkBXogTg5gnJFQAE3rwMx1FxuO7sWkMH6u5KuCZk/9fahqupROXoy4wza7
7ZfZPyet0aXUWY8o6X+N5nN4if+QqQuGCiof/SVbq62elhYnwVRZn9wHn4lTaQiGnxkL8GhNgF2P
bGaAN5p7zxIBKrj3nhrghq3XgIfeTfuaiiuvrGXRh//HmnxPfoBMcy4x4Bf3n/Im+eIpg4bNkbFp
WT1epkN5dFo7cE/fGME35E/XrHBHXAOeFsmeXqnNWsmtmGQ/VugUErO4yW9Ntdq1ZRUW5KAsbatJ
zR2UIL7/q4ONn6S1Peps/NRy0WcMsqi8zAvPsTbvyHs9wDmhj1EhmjU2bTjL8yeDB+3jKr2rfC4s
OH/Rjvy7JofhNNjNLHwFlkDcIP6nShS4POQg+2+X5YJe9yXzXPSrELqXbj7aFnwlPe1rTPM5FGa/
9MQJnLUeacv+BqzYlOfylS5P4/jgeRv2r2pOjbA17UhUIRee/u8KpMGv20+evjhzEg9HP09ISO37
CtEBWpR6Kvx9CN6dWq/xzH2nQwtBJwyMG0mPmXKcJ6zvyq3A4CpxnlCHDuACawK8EhYuOiYHUKXH
ckbJ630+3pEE9zy5zyGDYp5Ab4z179av7u5vELplztQC6fF6GNgk3Earc0yzxhlZULj9VeMdZFWr
ifLR7LvlVIlS8sn6xuUhGM7Ov9bliwJpJOBX2FHbeHtSRVmjfE9fry+wQ0UCqxaxJimjmkPs4Dkr
rHRG2OecxgwbD95NdSB5yBt9mHk5IeoiCxOrX6t1dPkTB/BWj0QhlvxCoVs0pzuGpyRaFEbPjwx+
T5/HhG+JZKeQGYZMLwHYIOfZu/DyIR6EFlmIRfn3mTMGH+yIHOx549p7cQFte5iwbajG4T5TKtJp
0gLFOp5XE8RjR6Vj1y826lZlFdSJjExaY5b82Mj2JlUZvmjL6PX1jQzKNqwhk49j7qMLPPfppDXk
gDZp+1h7FpZVG+uCz3LfwsmWh5aiikK3CJTVlxoN4ADXKn0fenOnQXUjbAKyZE5+cTSLPyc/LpEi
0yeYIr2CcjM6oPcch/j5GgS75OdC1SErLIDwDoEbovV8bv+AoSY3yfil4ajJs2+7Rl59Adn3Vg4V
D9GIc3vxWFInrQPeV8jLWe31SGEFuOMbdh1DBLDD1aWLah5ihr2rrnS7d13muBXdDZEJkQLL1Gw2
fbID0ABvpOzN8F5VN98S8D2nnmOcOdQwf6lhB4PFsPjffpKaMqT4YAnOg4+aVdMvEkfoiNTnXK4O
tI+Uefky5BWspiADu/yFG18k0p109UGYS1ex4zlh5rMCAZ8UsLXxQ5vN0ku/zEMQLzK2rrT7XAcN
4zeTYMutYt4cfqCak2+cR70pgjPbPHlWSXaQejeJC6epYqpE/mYEwk+07f4jFyGcW6FvjiQL3Jra
LoVAUoY2NpCsflrig9K8yWX6o1+8/so6yl7fhdIbEJbeaci6L1URC7pSoXb7rz18v3XlvwLsKz19
1842ZgbKwLfcvsYTb1LXKQZpb9OmEoFL1iZjDlXy8+CvhvT63CZvxd1npaLCRui4DnlZspweJyNe
8xfKTTwsoA1k3Rw4KiOnfrY9I7rJv5irb2UDG/airoYHp+YdHcbQNDUWZTa3nw9CaarEDQWCqUyl
5uk927lAX64uR6kY9bA+iW3VF6WtjeuaSytCTIuqZS0dAgVmBwv9ZHCbTPLSdkYP1mGwEf0MbSOC
YnJyrQ9Q3AmDIi1xScEmEatMyH7C1+OTvQLjKAA8mHzt79JyCy0zAxiBqv0ScSX2rkzuz+LWmzIM
q3gluHNyolxlXLE/AnGilFacSI/uddQOyULgui1AcT0lhe98oijwnVOz3Abnv/a/bLVB8dVKvfdo
MfMIlWsa05HvVoEe8J8zoGTcPISB7LPLjNsvWkn3ULgkgJ7NdBREanev4b9XZIgStXsXzO2nXifH
btw7KO+mBPJkyZaoFB3lJudEI81pCCM4mXZxM3qaSF3+0WM8yZUVGAHPA5M9U6Rx3OVBKD98Ch1V
GdUbD5FtYXsjL4lGCVcOK/gXBq05gZsMl/W6guWmqeet8/mxV+VGwHqpmNr9K7t/sg9XsE6L91qQ
tcpsMhl245O5ISilmtT5kjTmQe6UCYtTMiwNxJC2JFzkMY7IZimgusYOA6oCCJ+ZW/ogiA1dAVad
l2CSS+O+/lftGC5uymAlXpVftQ1XMQaZaB89tUMUHg5cOGt7G6vxSbD1xpInbgbrfGL5tyU06pFw
K0AHbVXe+nOFF9it2312mgaSuay0qN9jSeY31BNsCW78pHLPCIf7pJXZNaqFIesJdKDEc8AP/4os
dta2p1dcmO/3zzigrJhK8zPe+NFNl8D5vvd8omQiAyLpvuyreP4Ozl7kjfwpblkqQD2XrMnLqp2a
m0V7d2cLx5zR0sr2BR8JDnWDinPl1jo0bVWj+oOwazpAyRaS4j005M+KgzEihWAzPkXaCUdME7uJ
kaH3CUMIXGSWcxbAPfP4cDSo1F0NZTubQvP48cvLDA9nM6EAJ7Qvx+5BzdEtr7HbRHWdrVNc2GCe
pE+HqBh4DsfUZ/NhStug6xNCv+yrXvh8DVJz+4WIN6ad3pDwOTwmmKiyr/dBJGsvVSVDxmr9ylGr
PpytvCXpO873f3Sz2nQyTqzZEHnU/X2ZS2fIkxNRzbf/YoWwvXELdC4j3ciiPcYKxa1ouIHv/3v8
j8xcH6y4gHEjiOAz+TegqahDJJxbvHvou6E/sjbCen4x2CMyw/+DQWb1spVd6IqiXg26hakod4y1
P6w+ww/C/pMnUC6SmZq3N8kT6RkBMfZaMKrioJhjNBzkXMkVXOrRvy13M9DSEQuGMnOM48aluZvm
Kd1gXkyCANeBYZbm4hkADLZa8WTlJLYjm4j1XqXvb6yXs/nZC7ZlMNDTBVJfbnNYWnFpvSUPgAEe
Nm9g0lc3F06AJ8CagpKgrAWifvjjZMiiIRF158J6vqZWAzYL9WR/GxEK2h9AOxTpBN6LaofmivWT
b/NgqOcsjJ4qBXRPRIOg8rfpAlVTGdJ2pfzW4EU3AhxXoDsJZByJ2/6/au9na1I/FwtD1XGiJI95
5mndg4kWpXZmPzcmasvy2/IXxRVOmlAN3U0mLC+zQQQ7bXitqNrdqPWPPdRNwRDguoLthHUwFIum
ALAhg0Erg0rZzcUuQyry/HzzHMl+h3IeS6muB8WUXnW74EZdY4xD+VtaVKGFs7oYYEVvoAh74Z1t
ryZPbhfu1iD1IxmQ5w/8arpPO59EQzhrmrl6hAqtEqtj+3w5cfwQyYvNyoZimdTMVUPe47CtNeOu
6LgErX5ubPtdC7nkD/R4hFHbHqM6+otQ5Fn5SmmEalrlJCnHNTUNoxaJSwkrGSutZIhIwB/CDuu0
WT8sb2Th5wqft2oE7gUJfvBT5BpNpfVt/Qi5Izmen0SKakYnLyriBhqbMwu9Dlug77YaQ25FQMh2
fF0IC9xvrU/N71WEJiqIbX+DM5C3GwGU/P63WgmRSqUm7KCwHXmcDwqdnXFaMpo4rqV48EE5braC
ZWa9sbYUrJY+SBS9wNjHgnKlF6qwvE7gPZJ4Mb0MBgdkr0KCleHjWnbJWRxXtPg1KwiPIMoT5cOx
Oprap8jIPsEvqEB3cvtWeEBqZSv0AaGsnovzqNNixKlP8ueRwNxx0kqXPK5K+zi69IFHPcVmK520
fm/+lp82Tf+Uff4tAJmzqSP9NUKvyLRUoU4PSqTdK1OT/PdNpXplGL3ePF8SM4tJHzrjf4daN7t9
ZKAxK52GaOOIkDIUrwW/m62O5DkhQuyvCsPtp+tAxTfK9xFM0tn+3YlZyobqLtJJrmoLTyVrmkab
lsfPd1W7ulndRH4SGya9Z1RXMkX3ejLijQ9toYfqgoJKBCpvecLfyL+NIksRqe/LE/CxhKBXkaDL
nQ8+c66yzvLI+RcgjjX/Pwz1mFnr9q0SWDE/iBp3Uf9KJ+ScZ+dyHia71Had7CtJvTu5HJCPsEsB
kcIWxRQLSpQyih8Oii7PhnF3ksdOhc60mYul7wYPeq64bFQ7ksZhzWcbhwg5e3Oc00v5bgDPwGLl
vk8LkekscVSU4nkzmKWJ8Bkre0mgHKQLNFo476oUNqhyr6uBm0diO6hqM49J4rVE/95hS2tgv1mb
o9FlYYV962ZrtjBRCy0OkFY09i+aSIFDIo1aT3ThSmTBw5TTdIWtzj+ZxjxCekuPu1TCIhhC9RtM
Y7gi/FrY9TRZ4jWMJNDg9UcQOkGAb6fmg7eSyqxCTVk1Gz8u6C2LNxY6F4bFhg91fUiBVdeiBOQ/
K8Uj9Aoh5ge79+luU/n6UqQ2SxT/OKCwbH90Q2/4wdy+IbvylXloE2xWXe3YZGAP5VqxkZ3Dghil
jF6RA3l7pJCm/oDgZkNPwm6Hbr7vrlue8tICMhAzWWDIZFl0aGJBWehv0Lur2h4iyOx7PfAThkTZ
+Xep/SRdLOwWlSzH7Xiti7uXAjoJEZaoZwrIRx+bNcr4H92KmJbbxJfFdkeHPgY7VvPn5zM5nq95
76EeKCx1tZ8lqaM0YYKQswnGcduDaslZqKe2UpNi86Ov9gDNbf2E2oU4YfioYtH5FpeiEfuvjbFF
KSd3HABw0y7Gv/Yl6ooVsczyjoCj8ZbxKyTh5Lg7HEmo6wCbbfLbsoiiG9Y2Di8m6TsbZHdOFtvB
5jcF718HlGAJVooDcgSKMetSGg2wbyifcFSWlYfiggaN8kpyf7GP42tE/3b0HNk3PLHC9qZuqkk+
uS59po9xKahB5CCwnldMs4/+OnxTvgCTCao9hiu9YmvbagIbXXsmTBeQK169p2US1z89k0weFo0y
pdHh92X3Va21JqK0C78DIzo4qsE/XxtPPXUmZRSbt1exkdrZlHxD0q9QUmrp5iCljVAppsu5gPjr
44n3pixii0l1sUD31s+LT6H6dmQD4fheNEUAQ4vysWu13Bjw0riidLY68yNCtesrzvz3j7gTpkPJ
GsFh6Yz7gDrW6fzgz5y7HOMzwcVHG5irfYWADZ0eQoZERuRA1krop20W/Rl/UT/Jc4dK1hwAQFF+
FBsxbZChVXw+YxWA61h9GUZaW96zLG477OjDLyTKdeSIFW0UoqmWuBZ5BNGupieAxJxxFLok7Qd7
fauxFSD4tMmtph9PDwKdo6Fy7ssnpKTzeGSCW3qPDyC7DRw/PFocL21Mz0QUwcg4ff3Bcd5OHQAh
EVFzLQNt5ygF2WsRLuYyA4rJNMFNkQY1cpaKyXXiTDvALMbnFgyJ8OWb+ESt/IlmzQjoQmnJPjIF
8paiUSnokrmKF77zl0Leh89sW/EZ22azBxHUIPb+cNG21m7Nx/+r6Stau60aiKMb4vQm089g07mn
OiPz6DI2YkyppZ6Q5wokqG5tsgmSL+HnlMzVahYEwnZx40tSuyQEpq2Q7Mnjn6cltwKm6w4QbRM9
u4HMLYuu14q+eJaOQr7x6s8KQ/hXwVGQ0IJHrDJL8ht18kddA28s8PNaODT5omfurvz23syN0sam
9Ox2a7Sy5o9NDhNA1JksXT8dRbpAgS4Xek7/r/4/t2w7mn/C/lUCLXFaXn4nB/EyQPJ/9GEa63U+
lzcugxTOSeerzS+RBT/7e+zuiOBtuImeDrSbcOHl2NmqQ+JniOQ92AVvAQbUSnCaG17hyXWIVV6G
m8wpmrzWtr3wru2EEgb4FTlre/3yWx+dRZqvOCxk/SKrgkS78lZWnU1zao6hU3f5fSrqQk6dWVGL
u2zhoeX+KD4xoctG7pUcdvJa1UBgcxHXyhO9KE58hyPOYCM2kgJeQMM6NO5isWIo3vITHCTv373i
/KPvDO3yl+B34adKtH2UdgxwCmpp1Ys01p10mnna41/LIAwXeStvuLDXnQK4v8bLlO951PS/7AoL
ujWRvhY9S/GLQgKoIFI0SpA3GvwwrwQMUJvZzUaHEXOibu6Iz8uVaEjLUUSrgLOd4rpCFQHZE5r/
22GYnOIskAFMr5gB2cyurDTRNuoV608UlA/V9diKUEsw7RLzWBXg5StrmrHsCACtRcPbxNOP1Sq7
4lrmh1uwy5G1lol1WGB/g/5AUPGRgadOmKCnckyfjC8sKXjsgfUQRjEaBoB0mpeWMcDyjEsOqXYM
VZ/vdhrYjYr0SjygDZWcDQzdOvbdwmy+VMfdPBswJKmmWT42TxEyjDNLpNSTefCQZu5awfPsozQM
nLv0VVSxdkXvrzoW8T5WfRxGaEwbSac2pG61B01OdXU6wqII59eQ1BL6yoPxFOYkjDeAYTFbVRjd
AVUOGbSuBiPJ09lWQoUVnBR2R9bQwCJSlThE75fz/Hh0ChlrR7yheXPLxUTP8++nUm+LRE5eFbG+
vfYyxuN04uW0+wCmezIFE2jLzeVU+xNIvvqsWtaFSJywVH7vEYHczMSqJphzUY/U9+Bsp105WzpU
S32v/WHv5VJB2BAGAWgQAtqJkq8u1PXtEE/JNqxh0g0tdJSk0kkmcTK0ltmAnRU+Pw/3vELg1Z9t
1b2j++omOe7oJCoh9IjKzUnpNVPdTUOXs9Tr1Vk10PnXUpvaScG2tLJmmdcrLGDV5vl19g/adfPQ
EAh5EPCu/gksB6qtk8XflAzWKQ7z5XlWKvsDPYTNtIeV+9qWDoMlWvt5dUzSVRAe7JT5Jiy657tP
rlTzetlSRsR1obGN1bDInAqGCnm/fp8CGKiL3cY8s9avJWzapz7texhB3BNHej4N3ueOFJWZZNOy
OLShCetB8EVorwz4X2Yx00CselXbDRp2Wxf92kTQ70zQT6S1dZ8LEVJ7/lcczgOKD/CSlKjrp3YQ
PtFYIm3C1igglLt2LBEwiNnZRdLLcl++12F8e7CTDq84xNI9frZXJjSsj4J8o5cBd5p1QCfSUY1i
YeD0+TfiItRM/fSCFmOGCnSob2GptFQnpc7EUdi0q0BQb4YLTJUbUEbZmA/Huxm6zkbMHJBkj+M6
fSvR91o8q6CbanRutjxpI1nl4nm+7T9pz0LhWzxfFAfBOnqei6Bq4tl3TSsxpebXRUiVunWO3gmL
ZdPL5O5f8aVOQ2vKrk9xF1m0pdR3bi2Ai63PUgGTvg2Tyt5O4x+rtoRgu4s6sV5YjIiBpMelXcFK
C1NeEgJxkGKcvaoRdPSjDz2sQzEUthECzuy9taXBDBHgycUQtwcyl3Vlcv4yV+w3GOKdQ5h/GLBL
5URSkRPH7Ls/5xXghS66refcRoO6iz3uniPu7QjWMQgotXj1XFpRxdW23e5Vw6pCvPA1XXlRPEbq
u3RHv4R7K/DrJuwGYwt7e65XoklmZsxzO8IUEnSL07FJwl20FdKM7IhQ+cGLr1iReBmboOYiGMqD
AQBkKF5DAJ/ck0GMSdEjLn+OO/xWn1cdgG9qSffQzZSUMdHWdPE+WbCBjWTPx4vKgcJodybmz/6g
YYY/nCXOt+Z8dn3tsaiT2mUoUS+AxrwncoGGR8wUZCa3Xavpe6XCj4uR5gHaLkqe+2SIH7/CZmgy
r76RR6Gyr0cE5NMDCSsfcTqajqZ/vPjebI6VaAmNH14Z6pvE830qHE9PoQwSfiMMPopBhlOz2f91
qIhLV9RxiUNr6gdDuGpmBvVcuD+vRQ75sbiM9AE0erSydJMT4GEClGy+M+j5bBPoZ+YnRMHgu9t6
W6ETg9/wofI5y0zGpWaZF5c0I6Fy/t9Q2VjXvF9HXG81mmOzzwBf5QAkw1I1FTFxA9Gv7Bqx9ueD
Zt0oCzAdPcDA6wgyfb6+GSFZG82Bn8DKcs5lksD4+Roya0+EyBZmlcfw0Mip+MwXtn/s4bThhR4V
a7tnSGQRLnB/PYLDA58CdUKrIJqoUcj+9gqNuzM1P1elOTicK5noE1U2nKR0BwxXFHDD1uuOJrE4
Vlk2awqf8oYrDCKCHBVjse5bJR1Q5bhewVzqihBw5T84nl5EyeRfLDPwMN0iB4J7rAPtsj9rBFHs
DCsQSufBiWmQog5rWe68KOtJcHSJFFFzOGE+z6vHp49ueDg+wXbOUSeMzixYaVWYzt+mUKptyCqP
d6MnI469ldn8iaBN1Rcp3B84+aitx70XB0NgXOXNhkoCeLccvkf8rGkQYa7BVkQk/WB/sIW93QwM
PgFVlz0jCXFLmHyAeBdnrO28+x54RID/LpQ2CuvBoI2pL/BUdYwDVCWA8GFtGmIQT4TWhHwRGEyV
Kkj5lLiexPgi2Vj6FZzfAQQ6GOaIdKZ7sff541o2ZE5sKhAOXA5cSrswrcfsGWonZsiLr/H1qOOp
nKeKFSp74zOe6leLMgsi95+Gm27Tw2Qbm0HdghGJ4G0X5rXslvDG1tjXac5xW7GtKTrwJyxjEAwi
ssV1w7WqA8D5qv2JQ1hQvMLXQ4iDEM8NnMNOB4qbzFqKUol8h8Ip1GoB3RM+de/9fpagsurDRqg3
jjyQbDFCOx30cMxmM3BB/kB48uL7uUO5c8X2MKrNqORMCxzEHqXm2QSTsEEfHZr7+yHfJhYORumZ
lJnzRzfZXBpYNgT13ImlaaFceKBNRak88QAZjujUa1VvICX1hXJS7Xva2ucRVGazPLbN3yaYpjco
0GQfukRyka2Bd8VMzdOJToZx+1r9RbJ7FcXkT/nFMVYij35TFaHmpzwll9l8LNddusmiWjg3ZvyP
22p+nxjUktLXFssZTRPP9swU0Hwz6zsyymaqfc8N5mnGuzvgy0zrX/y+Ib2BZBYppnD2MlrxWpdK
9XSDwQKXr/S/pRXzUp+Afpp0OFzb49adLJgr2S60sjUVtRdntsNwwo6pvsh9KY67XO63eM0gQLp2
BzS/DwTs8gSgYqkorZSbmAAdbyMt1WZZMlxPgtsGfyHkdZFO0+BxyDtjJ0zVwjB5ouSsDEQzBB7Q
5d/Pi0Re9nupS/m4DJSoBmc5gKEU/TRLSznv6nPt+ThWt4shLJ6755eyZVNAZbsTwjJ3Fv9M9Jpz
5bNO5+Megw9Rq3eSsvPnxMU/WoIEkxgff2iCdhCMFF4ODXBnvoUSSEG+4KTLO3fEofk+gWVCv/cH
/0LEv3j1NlxN3MSi5K23H9M/pCYdECW2aDL93+9g9rsMB+GBJcL6DUiduuUpbzPB8wbaNkHlo5F5
WwB5xxM3XkWH64wjj007YtYbNVG4uN5unrCg5CqSGrranYG5g7gcuBJ+BlbrBGVIT9Ouf9bi/uU7
gDKDLWn71aGx0wdYmdKD8EcLmxa7sH3Bj47zNf+nsw761bZtvbn4SrtNsx8LbYfKD+gGrpkL+4UJ
YsF8jjFjuanM9E2GgMRCR3o+H6Dz1nfxp06zTgQffxKcFeu3AZenY5wF5aQtnWOtMsVKA4gdUFaP
Lka8kRWYtq3qZ6XxM4LuVx+Y/Q+gF6BlIpjBh0W7yY2icZl8hPl4UfZubbeXhz6GeINlUCfSDif+
W3xCl9wstBO8G2Nb18begf60CNkr+dwbuwtLmf6+dveGBMTLLmJQZ9rtXeMKR5Ndeii5KRPSUugf
87wshvD+BxSEOCqkB2rp3YTuluXGtR/l9OX5Cg/esBo1B91w4+jWCNIJRcIlyHeeduEfXAgZKS2i
Pb2TseJWFVXTCiXHhbb7nOdSIY1pz87GWR/wQx698lQ0PXTGio3JZ+0X6BsDrtqMuppNuz3tj+gS
NwA7Z4svP53T2EybLkg0fiZx1RLf66bgB95HSw57g9FBYpfPsKEyVR3bvAVOCiWHks+JFjE8Ktu4
xbxhbv3iHZMh/MXtCa9VgRXZu18Kc5WS/j6UFQlJcOc4uwqENCiPiI6W0Cte8TKevfk5ooXjUSND
LGqn0kVNPFdw8BsoUoIQVZs9LtpHiwZ4UOZhP5dyGUG8M35dKImBVn3S0gns/bsVIp4zKiSP7e8r
BNSFBdUpDzLTn6d5vy7QvKwdPqlru/GQ7vMyrEDRb7d8a1F3xZrbwJJExEI0iLp3TQCT74UIdeq+
aikDaRVU0A9MqwOYgXpGeFcI5MTkAYyM8uJ57sFNkT8RR2d9e1vVSz1xAxigfgrmaOwMtxYH4H6w
X3Jkv6EnJPud4LW5DDDqyloSOqq1GtU3cgYMLmShKjCoqdkQ0vwmc2M5ephSAWoObMjaorW1I0Gu
jPgg0f5kdwQXcQ9wVWvlDgUvgd2YzDkztq/9q+0CG7CmZASfPOCxkawOr8DwDN+qj30y95rZep1D
q/N/icX5ZnNQMnhDtvREYUAJoOKA3u9m4kJ9v8Wp2KFxnJyJH+IPApOMYPT8kQlTYcRoqkCuFDmw
PqR+ARPlUzUNDehlcbfc054WBSAI0Udw/pjX9gfaVKLqcv+b48Sl7GHmbZZOUQoJa2eJSiA5sTXJ
5L0fC5S/tRBDX+SYNx0OwZ0y5Gc5FQe4tG0yNf7CPQvujC2lpuBEh9Q0Nhd9PB6FXIOX8UWdQ4O3
sM5rXhkWmtX+vgKBWi4/EURQfFvZ6oubCH6UeDsywyrk+8NZ2lCdrkMdJkJo2jGm1eYpt5Kcypc/
/LtsJV4hyjRTjACjO1qXFO86tKdvewV+9C9FhjXgEfPNcRbwx6GWXell40aRAqZ6VgjlX46NGXaX
H/AfAyh5fZzLZw7MHuZTjBAwugDp9uXABlrYAPEoL0yE2+JQKvCC0ej52q4YzsSTXvZUpkOeAyHK
WgL85wk5QtBQ5iWrI5K/wWsnkuF//e9QcpUYtikayWaxKGOnTSAtFvEar0Jz8XOzfQ5J63Efff98
ZXi3tVmeF6A1zN8e2KlKr+6RZTPyfOd+lEjdjskSDTk0NRtvE8SPuf9EWpJNbHE1lGY+FtlmKE4h
iGMtGNN/lA8Vrzc86TEd+Gi7UM6brCPmYmXbhgmYWa05k4zJBl7D8otNqQ46tIYotQTfX9mFFJ4I
yAaQNInSOFHgqcDVs2dw/VUEmcLpeV1vd8uBGh9I04LYTmIvf5vacy0uGBKgcUXjsO3jtSh7xj6W
v+RPUtRI9rwz5J/DA7Q9yTwK4dBXTpGfe/BWxMvO1QL/PRbn5XMeVn/KPJSdb2yJPZ5pR2WNad6Z
UrdtKbxrSWsm9oaJCqxQHZrWjwOlUGeKBRvnvBHKaCnVbmiaT3CYGvc1ClJTwC6HrRjJD7Ri+Xnu
SoX4tNiCb0Slh3y/LJw5zAn8YOTbKOlmy0xIVFvqhdhJcXfTCLqaUy2OXPeOXE6UHlTkBvpGTdVd
6PWT+pJhUdYVls/XSXJdht/pkFU/klhpyDDENLt0rzD+kDapLhYqzp70MNb/0rPpXe9IT+LQqEFt
FOTixY16NOWZOa3sR8Ol4X9ApsBjmzQ//UWi2GpYFOSGoym9tBtIoVgmHfYiKnGlQN1HPEmXQ/rX
gtdZniDUx0tPltOxeA2drTGL+BtEat8gWwiw5n+hjjj3UZqf6odN1D2Vp227Ssi2/UwKR0/2Wt4X
ek6OtH3uqNk2YnufKKLuMfgbkH1lI3ImvThX2b4WH+TUYaJ8SEhGWTtD3xwSr7GcepCFJnvBWdx7
I3+m05zlfR2BcP2yz12t3QG2AGxtf4aowtdzHMz4Lg6QLNTo3lBY/hGeyJrd1YfSzBwsa9fTHUcl
lcK7DMl7WcgoqI6DQnHUkkYOZlmQMFCD7Ba5YjXh5NhTSEoPfzZDn/d1MpU7JqLFI6C5yevIgspq
sFcOytgnE23VberOeph1/8WsamfIoo4Fv+sb4BoxNgFnWDmLpYYdsGchVq870Xden+vBAGUG+1a2
Vhna38++mojv3zwNFTItUp2PVEBgkeE/WL63o20/3Na8Q429lJEDbsnCADF5g4Wsw/V/QjrdbhVi
vK+/fZZRKQDlUTlZrM4Q+4peTI06BcmT1hn21BJfgJjdoBrTsgMNb0zesorr2M/iuG89+bvySW+z
OexYlq3+L+128CQzCOuVtMXtmY42RfVbehiQXHYbRcuglTsTWgB8YzbgwFY1C6Q0ukc/9j1Xzdlk
PYTSeGoTDzrdz1lYRKpYgPJFPtJDlgmMzmFWBbyxbRmNiYe543S9Ttqm5tcR9WUGx1Rwig2LPS0u
q+fPWmOT8TYhOP/g5e/QFqCgJtf20yp7y0fg0BZD1LwCfNvjV/G2Ivvj3o1bXtD8VnBch/31HtdI
mhufPxgXrScygHgPmTAYropIjT0Ov4EhShL8rmZwqGPtwplu+/EoRu1+nRsxX6PAbodKzW8osQSv
avlMgrKA8UrcKUExaJyPJgJSWYlKP1Pu7jcrClXz2kw96evznged7b/p/gWtlGkTJUX/m+9u5IE9
790PKhcFRawVCuyAg11Op1x78ivoDmqrYOIV7a33i8FTUS1vNAKsy6WRJPUEOLhgoEIKzwIfCOpM
TmiPQe6WBJM7w0JWURKw7d35aykHeYrmchkgYi2LrmF5HH6OQQtCzPU2HDqCljJZcVhWUeiuYNYS
Lvl3yJOQ2l05HgRv802ufDaW0t8TNCDIGWVR0nuxpd3ewN3XQu3LSA4bGUQX7CDet1DvDWSS+bS5
wOhuzSbRgJwonzAFxVY/WzHZlfbkNfzwUcynsZeaGGgid0j2n2dwjphSyRkSByBejK/FJGgE+Z9u
TCRBb7PkETC+JjHIyD3P2p8zA8urFgHuaALt1UQKPDnzUGbgmbc3jjWvW6uUokkjjXUwW/dpSDcW
gH2lMJ9lmQhddOS1Zv2AJsX7jaAXwJHi/Fx9Wln/S9YAWv9n7uSgvEGkoobbf5tNOyPBCI8LL8+f
jerKsWnIe3NtNh11YnKJplNnL8emqxsZKGEm7j/wQ85brlivEyjHxrjjbJeIlxutY4LOct5GgfXN
/fpSvlfIsi47Wj6lnaUBF8XLcVxHPU1lNqb6HvqfRH8ACNnYG55qm4rsA9vS1/MbT2QNsgSEPyn4
syu6mEjYzkvNr2mqQBlfsKRj9i6h0w1qDn1R+WejuMbfswUTGBlkv8c9FDtjkiuyh2O0q1+x6dzy
gZSA8SnSholPlU2Hz7W3HuEypElNYoXEVlhpzmN7rr1Q1IPXJCkCl84Z0wpQwQzOnaR3WYcycqjI
Y8J1Z5DUq6f3pGgXpoD/lxiAV1122bllvo6Rj3FeuBqXilLhdm4EoGzyls7G1mxW78z9v5R7PStX
hd7XdTmQe7CO7LuVSJ1UXib9aBLQa3+tACEwV58TzBarAkaXJ64IKtSk9hq6B/896onTMm+s3cVV
0gAmxP7cpmF5I4kvUwFvPxZ4A9jue0qwH4wdo5B8tvOnIV1qQjR78y88A7QLOaODk4MTDP2uM5lq
N2p3ssG/ImkiwQEvj89zRV1KNgcEOdmtzV3fFcfJ0o0REF+r+rM7odNPr8Xl0Ru3kRewMQ4R3Gqo
awYuHEJrhCC428l6ih0jVD01US/xcLTSixLz86hYldHvudc11hJCN+zaZ6lYAnWU2z6X93Jb8S+X
ESrmhSXTAZr3GaWXVQ3LzzSDkSCaT4bnNxaJTvD+dQuwqW+KYVUWTVPNY4XKgTJHBzn67MsOyASq
+YTFgfrHUTT+quTH1sQ/K2HoV34Cg/22W6nhf/AtzuyPZZN+IzorC5gCM+nm+aCxkXCD1qxVNUo6
Cvrs0FwKYcsO4mGLSkrQsy8vS01MLqztoefuN7mvluiQ7sJm6VqEb/TQQ/Y77GL0LCjhfmiSBCCZ
p35Af8CrTHmQqcnBfmHkT7yK1Y84YL53/p6iIXayd7O4TEsd+p/oZnOst9PcXTPQvZqNs8ZHDO3m
KK7quYSs0qZECZJR9tdiMo1hPX4LUAWSHO8OFF2oJJcbXToOx9pMRkaXsV8CcgHTVGNDg5z6pWZg
TqFMcqMvQk/4FGDWBPpQtcWnEOaTV4Qh6CeETUspFp+KyE8FgcVUyRlFTheNj+W+t+JnshMT+ff8
SBo/P+ddlHy86UetHDFeKSGjQQCHWKNkqNSPvt9bFvDfygyd/EWN+xSC530J0TwTr6tbsf4IBN/z
0QzAwArR6vPQSaGqLy2K6trxh6+Q0mvendFjanbC0zRFOiBljExnVyVwWEjauG/uZZXGXf8oe6CV
brlTnOBDctpDvbjS8qiTV22etChpquMvJQcCBnaHFJPsBx8mmGuZl9oZ66qxkeUGUQ6lgylc9yiG
fMcmpq/k/yQAj1WTb3i/KTYzSDlbNzv6B6llKV1IJ4fOuFeK0f4uKDofH4noT0HCRsqWYzJer7CN
aTdvMFWcjp840jJu1UBaCJuWsEIwGj7v3/zOf7H1FRCDqYPzihrU2YsbRerwaQjxokdG1G/dzItw
eaheVGId0oPvtaDptchNVTZ73qIFXWsRVWZ3DmY2PcE7WrAb/bL1Z0wA+BnlRoVbfGjmy8nWIoWq
UhpA9zDb3e6oDN1BMgryPlIevriMPZf27rmlsri0p6P49VVaZlxzHE3ZmZJGmVK1+nlRQakVTUjd
4g0FIyIUV//3bmGaRXaQD8tTPFjkn/UwV16+uYeklDLIwuCBXOjNsX/OYaYpd7c3DD+w/JUPwtaB
V3ROzt/2ZfhMx9WmLvAzr6xIa2lDnGJ6vGswn/krx/95DhIgUOAQaNEsB45bdWt8UiKjOIR1oisE
aSKPXnSbOQxqLQyp2SnS2TcmfC3xXRMKqJhusHlhEu4MExT1Rj156gUbMlwj/+PB/SEgcjC5Vl2J
PBxrA/UCFOV4VR2AueTPHSqO3Ne2xQt+beNaQiVi3IlCweiouK4HD+ju0kWTWhUcB7bBwdE1ilLl
UgOw3PZWhZa5MVPHkFVQOFlE07v03AXXNLL2ohRtSjG5wXMVerThRVAmb8/mCO1xUGwPWDGSiNIn
L2KJvOlFRDGn+HQmc6KU4a2H51wkVaJlDkA9BHZDCwNEkmgA5zW6BfhgFyUAjQ9AzfTVUVvkGxvI
pbQy05apDZe+eWEDjC6lsCsD5gVhesZnR4QM+YkMxuk+GUoIr1oanWIiYqM/UOKJfKwf8Vtkm0ut
mPfWTu54qsngWRCLDI5b3tjXoWpsnAoWxMojtk5cAAixwr2YmjkXqP7E0hcD47fhx2lW+5O7vtjO
ZfQh1fHhn6TXSXqF6vtf95BHzt0Y2/3PWzrhHZfBLUbDHjfk7MWeefsvQwcCffZgAMUZnbHoy2bC
N+3ombP7sfILfyBhYCoPuPdstPJBxIf75/j95ezdreIwFZ5uo8LuGBvlIsQ1BLTrCAfprvfY1wIM
znaC5DqP2UTD5K8d1b9zYTzK8moKC4ThHxvtg6RylGAO7ro2ZNCgpQIiP9ua4aioNHeuOPVwRZ/I
+yjdB72Q2+23aoo0x6pRGKgHt671a294ldHfV8WPZraMP5wJzfb08IrBSdKvqFZFTfTg4SI9UC0O
Zv5v6BSAgg/0QjTad7i36I33bFqRRQ6COQjrtXCnLAKDsNb3V5owmhyHkBULoRp9p28ePl73gOiR
zLfdR8DYibtFVnKNPPSAOq71BTYjsilZl3M1m9vroZmG2sCcnY8QcDKpUW1nOIAkceyb36sXTguP
Y66GFnkyToS0NkkaDiVP97JZpt4/SfKOIzezkbr4gQGJPx+pdJWlVcMbtGlE3KTt+pOWckVIcCs+
CJ9JFHCE7jtjAc0I3Vrginf1OpSDTC3QllBchLrOlq5aCsZopqF/CaSLLL1h4I8/QQDjuizJPN3K
uwV1RybGccAINWAXyds1S2QwGeD/cvKZBcBgPq59Ym4UQJwvGi0Q3DUQsYYovOrwBDRU3XondsYL
7MDRs56mGX7wA5bsgZXna+B9xjchyKEibHaw0eCiWUHRwQ2yK5ZthjABxorOGPhpR2JHTWDOhiF5
gC3HukBd3I8F3gtcenLdjrrWNK/fY/pHrBUYvszfBIKFCwdW1BW8IiCRDDAdUwLh8gjDBINM1KgR
WV6epxZfrw3iuto95EI5Zr6PexEywBAKKAb5511evFuk7KYdaofe8oS2YaOQTe6x6VPLljfezfx2
KdA1oBVxwOIuUSrY5tq4wvr+/MdIDZViYLF29svDkrXGqYB172qi4MlEtnvl0zRPe0/VE1FbvOXh
+OaP48EJVFx3L5GoUMQI+vtrfapdtS5ny99vYG4TaEvGhQSkcRa3iwVneXz7aB40yUm9uPPmc2Oc
58YnLJTZ8058Y0Ff8MMVqf0dXJVgK7wKC746ux9ZqjXHdOdUUR4pi4EcBJQNtqYCRbNh8cL/8ejR
9xqIoWcMbrVic1fHuVxF1KnWC7B9W2jvqLL52Z5DdnH6RJWNZmKvPNGdgLr3jEsQwAzw2uiBxL2X
Vuq1NTcaUWB1OpRXibQJau37XT3nAys43/4Uk1+fh8gFLp75xC270VuIVloAO8kMg5YQ9il3a/ib
koIurFZwRsPn3aC3fqd9i7j+kSex1+aZNaCLIGEd9D3sfGuqUB41Vn9kqEVs8pkcbtsy3I/tkb94
u1+1ZcmywDwK0/+jykbTBmFYyfvlZToG+5zJH8lmiqxxFVxrMRqlCLx+CJJcgIGIBNy1oDtMOxas
YIFjPdlvMhnwEX6mBNyDjbqIx3CAv6knIt2VpO1iwOHCiYEcZ24HU/FOkFiaiV/9Y4eAgPtumYSN
mpkD/PcHSg05tKTYqTDRe2+VoIeLJ4rlCnDJaqYtAZ3DRRtG94HwrXKH5gAKBkm8yRytQcmqcWYh
yPDwbkdJLWoKtlnkCUfDuQCt01+bx0JSv6arVqav5tF+iZV3qcaTabUSxi67lq5vVWAWsRi0Y/pj
afuS/ukZ55AUFI0xW3s1md/skHdY3Q7MIKxxYF9vhJmikVRCm7ppis/nHWhZ3M90tJvH17+2/F+m
ixcF9/al43pEN7OCOPbXMQIjd8aRPQIK1HS+broS2cJairP5qu4zULhZIGFAp5MpQHDiJuENzE38
KDhoiSwz9+oFmStYh5K/AP73tsvoBSFk0Tg5rOKuYhSJNE5n+4oyozHPBAkB5y75UuJrCi/shfLW
Y+hSYACGYH7red21tEzKBoQL9jH6RFVtphAJFPgWhd41l12X/eck0XD5EtYXmdQXvZTlFrKcrmdq
O5ub4a4IXXuRsl0g3BHzNS34S7DQ7sXlqmFS1py4MUXB5a2gwYOKO7acATUPrE0SDGZaXOdGianV
fcmPRGtzPHmA41TqrrGz1/4lscqvrWBrTYMhCXtl2cgzno+QzV3207oDgIrNhwUaAYTcD4qqMIoD
tPCDAJAtjFfk5KFkSmZxn98EbueSObIkDHjLyNX1aGVT7AGtx6uOz9gJSJTUFwt/BCg21Jynahep
DgoV7uwfuuCqAn5LtDLQplSkuXrsJHkW/Gb80hNK0A00H1p2yzLd5vCDuDpA7SMq6lPG+dDxsj1U
yljWh9k+FEv3QW1IBgnKEBKMYk9RzUMdl5zgI8QF0kQTrtFPe/dnw9WjfpcrdLCOM7be1KqMdN6K
Sers+Hhm81Qefh+5yd/4aTSrQOb6OPuBb47QZDTi4Ijr77hHb4NPv87nbXTr3/p7N9OE6SzwGzNf
wyglXk0bW3VNPf6uOYXJFEp/nm+KqoCm/Sw9atw3iA4+IrWqLeC2FWFzGdDlr03OSPFefHpxUfqK
kcvp8SjIhYc311x0XzxjqSnlJmnf5ouD6HnBxIrOYGCz+opLJNoxI6Rym5qx8pXeDYP5e+hB/Z+T
1k5VXIwEajqpre7ABHBX90dOpqHXVQApaWizM9QLeIddq3TAR5MHT8L3f/bp1GY953QcCetsXnXQ
CjdVgcCsWocwlVo1/OEr4QjmIVd6HtaavIvfz/KWc14AfPnBhdVNqOF2hp/v3kr9lmoiOyo09Ses
ujvwto03aKP3HMhBx4uUwYpjC6usuaXiRGj6Ivo6x8kWvBao/FhYNdPkzwNJ3VukabQ7ld7UXF6/
C66wqsPdU95WQuwUdfQCOOgesFJ7tR8NYxPrxmkXIK27c7AUabK52P2ch/Q3lKcNeDd8B8BE9I/3
HVCi8vUPqr9SjItwgXUdbUxHxEXE9IldLdlTiM+MI1pHOlWigrZGpF3AggUJoL+khjO55Av0ts9O
XKusFVa9gxkr11ehAOkMe9TBX9TuAfCmmAqO7pj++QHtzvjHqiAki5dbc1+aHKLGzO4tOdbYG7FZ
Cd8PYrMbRHPsmkRbx53aBfzgfVo8NlfF38WQbzWPeE0UaQlo6REw74gtqzZmoNxHJVG8kLSrLs3e
iB2rnq/efe7744H2lTUUyA64EsPiv+IGJF9uE++HD8XidvZH0Kmh+uwCbYirM2hjpGAcflhtN8gT
e8cYv318QqqXCDQXVQi6mkDdcNzQjmS0v/yEhLi4vEY/0H7zUvKTpmCOXHahAr0cVsjA8MN1T/+C
HA4Xv8ErWa8qZcz7eNSRuUM2gUdEy8PGXjVDN81LAIqe+0vqo9oX0oBP4iTtAANt5b32agAKB/cd
JEKDcl1Ya9/j0nqthQIyw+5C4+4Lu1dIG2DesnhV7R6rXUd8Ah9+hiDa2rukP5yJd3YMFIap0zvc
zziAWmfpJ8/F1czY/Yw26y0N0CzsZ6iFS5KiRYsaTOnUygx/aSbHL/9Gfz42H+r8TMn9cwC+bu6c
ncMwWBigM8L1/QVhyc2/RuX/ND/7Mwe3i3gWUscsQHgyBeYaSFEEZMSx3z/gHux8QEPz3a2Ba6dH
721x6qd6eC9O/jKIc8jRXQ8oJTPGGxtTxQcJpAi1pQhKfNjNKEOuNrDU4tFdPQfEZSbyG58v0x74
O18iyauapDM7q6k7IgbBLvArvX2NK4MFGxaRSR351+DKlFMSKFIIX9RVbUnXA5pLX4M53kfzyuP8
5Ms5NhU4XtyvqFvRnZXCGyQs/LmkNcteWdEFsMMG/4knPgZAeUc4ZQvUHwbZ2iS7wFTtSDvM2SD5
GQiutXLC2Jym/3vntp5aJxkUp1uoY6l5Bl0KLz9BMventD0SJQiu3qwSfJyxL7fn7xBcQ43Snagh
nqRuAlTjzsKhyzOmaabZJjpLfUxf5job2jODWllZiMrjtNbz1NrIXd1XQ7KGjoS+PQeWGt3U5UfD
7dpe4yc042P+BMhIBIThBVQ0ueeD/+441cjDUYlvs4CQmq0tNVukDG64Ta2jIjqM9kIAYpQwwBs/
3wc3GT0aceOG+WeDE5B9rgaH927d95uUbQbhr6vxqkhu+CWeRC66v7SsG5MmMGuhbGNlaeWmydeG
0RRKCFdfKdxha1M5zoAUwLCFcmEMM2lgUvfMeqM78Sj/PngOxZrfHJcbo4QprIjkOzpQg0zDXz49
/mZiz3DJAG7VhaqMQt2f6qaFhfInzEtNlSFsRuZ3fU2PMq+Lxy3X4RS+pnR+jwxqiohjr0/wa2GV
icAee9oaqmds8nJOBPKQzbQ5J6VxXzDDL9KP4u4oGMkPqX5c3ns0Jks9XEDDYAzIqTAgzRxi96k6
NcddL0EX+GUGqIvF3/JJDRtdCbEOwR/okxZjEHY3mnebu/n2R31G6f1qBASPQCVlaLbjWoNCaBfc
JDmrh+1S0rMlU5mCJ38vjRWnNcDwa2KMMTTxE6btHQnmE09ct3Hjqx7egvyzH0VhpDJVOzDsaXhV
LLaG3sDPtBaDLvWapHIzKiV+TlepdP5g3P2WB4MYrbgJJn+MKHQCx1ykFzJQaWp2FIQwaNznd/01
6SIXgRbJMjcl5o0NG1S43F2NvQv2sR632ujhJTR4w/emj/9DOw+cB/BdIDzEmTJ+1jU5Ox8h3drx
i55ZzX+b0JzCGqNalZ/6A/XSrSemi9fi/IQ3B1s+Xy183LkA/zJfK6OKYj7rMwDgCpAvJp4ait3T
YxkptJgDY0byWEhU1yEABlV/fLXDvAjRrxuAcrbtIJlYoKQw75XRZk4ylGXZgHgKpt/2mhw1vKZZ
DSFBjCY39PdK2tLfBTpWMX0u2cbgqjhfTCsQAd0O2XFV3JoAG7mHaKkrW40OwEuwE+fKjiRfnRaV
jKtpp9viRJqB8i3zYwyUybd0Qmw+cIqI3b1Ya4zX7YpU3edVGV7x16dUJG3GA+l+wSBRYZu5Hot9
gN7x76yGp0dQrS4sg/7ByJ4xcvxsCVokUtXB1iYSF4Gm892mbuTQUExAgTr3Sn94vNaON0LMGvhu
3Rh1ytpA6f4YCAI+XONpGyOArHehAin1NWdMLcYUur0gKiWZAbKpu6+w305d+q38rWjPzhWDqJJa
BaHXMzGBhfzzG2K71j1AjoZ6FPs+JZTFlCg8/N0lFqbBzkO1Z95hXpcpMue4dgmaXF+Us8Jwasw7
xvxvbkkHa0rbf8ShICc3Eo8pnWXYch8PPy3ddjispG/le2l0i1iHV70JarKyl4aRVFtyTDT+ZZDK
VgBIockAKa1/gszsBscOUuZFMDCSQwKwBPIyQHhiF0uluiRa3rXjKKrpzY3wW9WMiby6N/nf2BIZ
HJRYxr3bxsDMfv0MXj/4+9ahTTFnPgyBN9CNZwM8npVgOooByF4xs4Xp7Ax8Yhuq/FC7XjcLQd5h
i2+A2ttod0PThQNflwBxXgcpM1hUZwk1FIku4mIs36IdGi6Ug8+9SLcua+eqQnDtAtoYZm/oscXS
6o6FurDaQKJLTLH2IotHWurE1wY8Xmo+QF8Sx7mh3sZLN/1R+/KXA1V5qiipFdYUsYfJY16J459+
cPdBhsu7o0ijRlwFZJhuxnFt5CK05DpKHlij4QotfpE5ErZANBNlknIwpU/CBV9aX1HuImcypD7V
8eLDp2SWtDCBC/TLQO7BzMlv2opJWZ87R7J1VsDMz1OeDvo3Cd7IBJ5sBzWWD7JH5qCL2Ff1v3O2
oAHUZyIAFzEs3m9TWOfth6YpPlF1QuhOaK4laK5xOnQeKvY58+86oh+xUt5HJIZPsR994OmOSnNO
7UL5sCiF3/ZmdG779NcM+Rv00Eq/FQZqbwUKPP/BAiQiIUSb7GMZdBGWWFgQkf14WLpyuxDs2iRh
aNTOhk83PlaQMZjJVPdWyfyzDFqdG+PxUQk0hip9WxTuK6HSP7gyDXD5+XGROlo5N94yywI4MSDm
ClEGr5QnY/2gCwnspMk/PoD9g1IpKocP/E48AJjPi5KSl80ZoKQaXLUsz4UEmZMQ3CdvPKCp924X
S2RufGZu9Ad7XGI4i6xYlEfK55cEvDjJ+kF1VQE5VWYkNAMLrKN0rkqcWB7zzOTQsQmFv36F5q5b
1kXjf7IjB8FpWCX2aXh4npH8L+XOfgCPC99HWvc/3T2NrmjX/f8xms8+P6gg8FB/nMOQaARyh9Xg
jnRJZ1shYFt38CGh/60KkC8/E4p7VcAwoBSWxMNP2JTLpnSsTX5RxLKCWFGDGHVk3ef6on6ACoId
GJQxF0WX3Mo468WT8bIaHRwwD5RJqQEkEDA20hq+iHJR/XOgxapNfbWVMcwIElcMHibgZEq9kQK1
WNpqSBjPsbM/MCUeEs7t//nR2YRuub3rBOZMAtjxG1b4+jYf/w1Kxj+wVUg6kkcO6APTY+QykeMy
bNt1GuuMA0Xr0KFZmLHUBGuU4hlf8hkGmh8TJnjYQWY3ESuNgApoWp31wQw4N8lclAG2eVbhZhVt
vflH4WqQpRNYQPtm/iYF6xS7l6AXbmAg7JQ4akW8FcoZqilrpxYWBMXuWGxnWhkV7EGvm7a5aHqS
ZBfo2r8+fUCEA1ibmHi0Txs8XGKedd5Dq7Xn3VtT2mlVhlnVDC0hiLMXozZORA98A9ScIpRrstiY
yV1VY2k+f80CiVxypNPyWnU3pcVuWaDHs+M/jiN82nmAk6MoivF6uimR4ZduTThCbGY0TEiYvLLy
ifBxjfGKX9vNCQcnl16uTd599PsI/55BWJX6VCURGCgWEdI5JNYByiK133tFreUoB4jDdEI/K21w
Bpnfv8oUQoA+EzeUSIjvfE/GuK91xExDiB906XMv4ubLA4oiB3rnudORMIuGJvI4OLUh1l7asH/Q
w6oG6MnOlalNlNgMn8PDAUh6jWqqvM0qx6mJoZ35OOoIrE4M0nLj7bNe74/h27Zc5q+7pjjfnGZn
d5spNTr9/igYG4pRSCw5R0A3Ol76pmqfmkgV/vwAnvOrxpDWexlrk5z0aS4wP8i2eq/i14s4eAfg
Hf5AFdGEw/e/WxT4yIqGrZK7L3IbawT86ATqgA/6dtlO76AfjjL5aLKpfKY7iU5F3DsTLBlO57BK
LMuEZQjd7Dogx8KpJOVFiQZdEgnK2s1BlYfCRXU3R4/ab53/MiKugo4E3onImmgJyqADiEGhW0To
m3ZtxRaefq7xs4c+3cEACKPTk8PahBgEITNBpNmE+wXnvU4PSwAMbW1LKcFGpdoybeuJSPYaalAH
PGQteaUpiGLn2cnD48XHwofrVMw/d3FCwkdFOGh2bjzVeds+VoiRzU58+oUwmqx3dEFycCj1gqDN
z4JBKA2lV/wXy20kq1ipTWlUBew/p5Pvac1pm3dsN+9GyImWOVM2bpzKu2/tJGJklxgHIoncbyto
xWp1/DS9m4iMVSQUXTw17kYZYnzhn9bPIgTbK0qy+MmTh7YIqnpSYwjpl6jSnBiDBAGAXiySKb5F
s/PtdDp6N/6/zs50wX4dcH8zWG2AukYU7n9TbDUUDCxtdDZx0OZPug37QHzEQuWIyO2VQaaYVa/S
SCATNeTO9uotEsPZijc8mwXPo/zdeANvPU6KagWtbYLaszsp+OIcSrgOyHy+lvx8HJpkO0BNGA6v
lgnnwnpKnnSyZhh42qbhGr1yDVz7n8MaKl4kapQR65TUT2p05x1RSa2bFrH/vtuBM/AqoU/fZRLV
j+l3TVTK70oLyxb9PIWQ/SrcNCrMb7uVeJLqSw/46j+m6lmVlOnXxTbF9r0aJ+Q9kUurxeVwFo93
ksWydvibU9kO+4+/xJWk6SvphkfdKVU3wKVcXFasq5yjgHl4FDec45M2v4sRF6gUARA9nlE8gG1i
IXQxq4zsoXEwX2NVl93O8gKD9hF/fLRURc4e5igfqRJvcL47khfc7+sAPmaXUs4dkRzoKdzl9pkX
/2JxTvR49/gAiehPY81IiNO1/qD4dBHA9wZg6/Nu5CgKUqcNlvJJHI6uaHVyM/8fAzodg+Y+av0z
JC7CC6+VVgvpDvz4FmCvOGXRMMDhtLeXugpuo1uqCopaih4Wugd4eSAI1rY11mTpf09E9GZe+JVi
OkzpueV2BnXQdrXgo7w9/RZ7Xt5yyhnxi3RPpzH9gnQN6ecYqiw4vBNyGEghFLpM8Tm/pU5aMloR
B+pnTdX2nBZBxaMdDFFgiO7HK8I904T/3JNXIz3RVb/RP8Jz6WOQlTwFUYwe3CLyFQWUcBrf2UDq
u2fZ9J7FYEkPfvOumAzBUi97nOebL4pJNKPEozSlsjh3h7bwKs09uPtZL6yu2dLSusMlOBgOG+e5
OH7Fcqm/5G8CBnzth9iEEDUgRQEBR0z5bMrhu+Ss13sN/sc3cWj3ovaYE8kFel3J3d9QFp2f87f9
ZpGIlm8c8tIvyinMJvP+j2wDMtMjKQHruPeOkJ/JPjMSoF2fqoVCAeKtEdBB3hEQn508z9iIf1gA
mjrvsX6YC9uNfp0/ofpxw7H7GLV32vew75HKJbXAJcYqQE67gQL4bbKzKdYBbBxih+8ndl2dJULN
UQMFWZ1UxU8IpWukgW1Epah7Av5d7DjkYLj2rhpGPTmloEGdjFNjjnRYtyCs/8RUEgvvN2mtIQT6
+kY627ixygYWCX8o3R9f5ORPdWetnuT/cyTseh9u1z8dAbK36DREw/tTD2/TPeiEbM7qQE/ihY9c
UcHKHbcSKZMbBNs3USkIlCclJaP5PWw+TtBnYFCygJoYvvf+aoNbEbiPWkSDgwOzs8pOC9e0LzGj
6sSoKszgZuSgMrm8hFUjzXCyINpYe4n+jNnCdHHNIrEDn1K33tKLUytAJTC+sDBjsA/anDEzif/6
Q6EOV+jqJ8pDrKzpDBX8ZGhxEP9CjLzrLWcvNK52ktdfF7RMLZdgqCp6Yalkt0OvspB3lPI4k/uj
//PiZvhbsujm3rK8ltZvkWg0LLwy7dX7fZlvuNwbNu2sQDEe77Bq4fGNe+je2sD9aqWHzVlWLREK
1yC1POnJXeXmbLIx7GnP/O6IG3kq0YAMODTdD8dBBDqlJnwiULxkEt6STdXTk8R6jWHqPhM+rs5/
yqEkzpBzGPIkeZZJr6ndENjjYcWOoGfRFgUq+pOSkL/AyQ63nKXuYhOIhWbcgCa/qPN2dvhB5ZvF
KCAbm7X+sNzWJ2ZI62slZnj9NebkEhcvabolHpz2oBrY+4Tu2d4iNKAJOhXzQo8QGTMPQlNkdlVV
P2RgtfcqfFtyZQzpEoXLHk6MZ434DfuPb/JSJkyQgs+1+k8Ykg56p/wzPkzbIaJwyFOvJ+vj7Zti
9RYCaPBKAHYavVi4invpNrF3YR9TS7ZAn7v4QcTtN+5OlWK5NDd2I49Y5sKflH9ynF3kB9HURDa4
4sNVBaKOXQGFDd02UBdPX9FDqjzhUSYj2HWdtBi56HCDlpIvk6aG+f5Acpp7NsaK9bMjFP+8MihL
jJIXRDjW9fEwValGGOLsyYUFaMEPwFtF8458BdgN22u+8J5JLKDy+lTF1l3eInl0MR4wxSHeUu5b
YBANCwhJViPtLmX5zcqPRfHS5314pQ9QpTqrQl4ytTZ0f8SrTes/RjtwCgVjTborb1zZz/bU+4y/
RJwmc/DT7rvODcyAxX0ZB2nLE5NZRGbhySLZjH21P8n/MjlVh6o2efqcjeoDJIqXT9LvqPM4kbA1
imRDdzoNN2JGMIyaYc5JBzsY9em92m3cLQUIUupvaeK/rM40s4YNVDPaHI9DVBet14YJsQEbMXtn
j080HM57NWSJtSuYxR63K684Wga7HVUtjlBaObFSkHE6JbdNvWqLF9dDRYdzDCt9fJjfHEFuip1K
z4Nf1hSJGwea4dESSTHdJIJgw0UZKZwK3yRact971z31V+YNXJpo48r1o/suS5abZfdEWF6IRNP9
EfDIeltLudnEuqdA6jxQJ3B58cMA9uoCSkzbhCUy1ApXuWh2bEnjddvROjcOzunDNxS78jJ86/sx
IuoK+tUMG+qBV43wPbjIF9lOKTPon1eez8OkSSED9oIul2L51xTnOXbw4beVE+Yk/WAJUHSoHaH0
FlV7rSY+xjh8gMKcp9U2Tss5N7NMiITy+XBLJHHYJ11JQhELL0uA2VapUZi3w+m/VUEUQvV5aeTK
N2JzyE/tR2C8IKoUnsVW+9dQI1W+i4QXx/e1mwfiOXrwCCczg/ydQ5iJ1h896bgPv89lp6q9SgLW
Nn3ZCwSwVa6DwxMnK13dHBnyMf/J5jjMvFX1Zyxtnaxy7/zkwwnufzVHZoaOVgXDLiT0frU0csRO
Q+HoAH3r4YcbzBeo2a0KcESzwoElc+4TmWRnfLqgUAIpQNSexu46/pr8sLE7mqySfBN9tQd3Ayrf
ApP87MQ60OKvm7D5z2qLWYiIz+mLchxMLRBKEzS+gMmTkVcdUfFnvoztIEGO9HYFnWP6LzXs+Squ
CvVvSBzc222F3L5PSAB646XxEhDE+FJVWmMAnnVIRyKJW5PI/OUHJ+fuN/BvXRxzfcrmBrs+xL4V
jch3P2DJnpqa0PfT01yO6siD7g4DhmO1e9Lbm1mwajhkvTEm2802SGm7LvT3i6bbkLXmY9eNy7/h
lstvqyyj1cHe+AT8dgy/TUI1p4aQM0zf3b4J761aMLjA35QlsIjAwU4PtWDwnq1MLjMCBsXm2NbQ
6ORBnjThTF84QXn0N/g0GNwSSP0GAOSH9hOGIfThq/1osNkspQ/b+ChwZCdRt1WRe9cB5V6KV5it
Mh7cjfvaIGSUojHwB8SbogmAdsq5SEBet2+b+gCwiLEFitVZ1DywONPa11LtwLvuuK0/SPbufvKM
yBtWYFNghBYT9WkUXyIrce+yncQMDDGpZpZPpJdW+HoxEnd6cycmyTWxGIwjGRZZSd70WPDN8bmP
GOhUc1xe071OkC3WXI1TbuFPHYu5wduiFb9TGqu9HBVeSOAG88zdozvDqp/vTt1ywyBjKvK/RWYo
yIZoOjl/5R98WhP6DgFJklAKA9SkoZxQt2Q2ZAQRpkDUaYX3srNdW96RdLPTktkSlCrbtcvXzXmJ
m3BRC/vF/K52EqbyUD103GIu/15JeSB7qC41Hj9civ2LQ8kk4F5TTY+aX0qUme6scmfUww7Stijs
6G1K7TcrsN8EPJMHyWxg0ejGUvqN037lnCZmGRH+draUbEz74rXhaKCn90vnj8m/9PR0DJ8iIfJ0
/RULXjDK342MUtgbkmyIgO1IQZYAOVlpSIqtOx3OxgKNGhaV5nJnDCQwrxANfIdl5ve5UpacnCUd
Pr0vFZUrVUfsB46+AXm6EBGB+fd11bq5fKfLr3PGRTJvuYmxtLb7ac4mPxB+yC0kMSKm52V9ZQAQ
2FRrksiIsLPnIGNoXx+vjdpfd9ETDGBtuZksqZDLWsJO8uTaS7ard9FSJJmu1JEW0pYkQLTZdHGC
plwpxHs7lxvzSDjhsR2rrmlwprMnYZJCuhE/OWgDFfDmtaW4dMxR9B/3lDRgPeAWQRjtY5PNxKhN
uKuiciQ1P0dF3BkSxWTO1ujjfYKzGJsTnGahE/fjTtYAj6fyS0T6upTU7z8+BEIbI09A+Jb3HK/Q
LiqUqh1UiGGXXSkZhsCvPPkjqXg87N0u6c9Q7ksdZStWFzWS6TXzDKxqWGubzKfwLwG7PvTp5fFm
v+O8CgvgOtrqFPAOyBYW7UetgpiwslQACSwIdmB/3x17wJKK4smvaFssbVJRDcaCjGgPFza1H80t
V9cz3ooyOlZ+GLSqXfhEPLvcQZdStSaRg56Nh5N7gsh4InLbz1kfyOD/Rj66G6OVD8RGD3cAcg/d
2yDCWi5aNaXJJsKr/zt3X/oGgYkRflcaMe5woZcIzlRCpffBP0Se/nvm34kmqV9i12Fz4fQ5I8hZ
wXL1r9hneajLI5Ka+bLupoCBLOyHDe6n7j1SQ8Y9HKT2ikJCotqI5Ex0pAcGn2YmzloocLawk8Zi
Bvn0nHbSY6cqM2QipScWJ06iEso4S/apyQsus9VDskSjnhgg2kyPEN265NIVJpWm2B54Pa267xVi
ni5m8FSRTjV14/0VyWVXo2yZ3cev4+mgaAr8g1cJV47ESYKjN36ifHZCBQ7X647kkdOfoJvA5Rh+
SQh9D+0I4DJf3WUdtGsOJhIVzAuNOQ3wMYPpgACiN/rFHK/81FRHA5py2QpGnizmBNZ9qnABchry
5pZhsx/oGJOMFgJi4rlhCQeFKmXJC7Jt2CQJzZQ3v+1QFrMbSaW2WmXyfJ4NngtHjpABOPgFVf8o
dQUKrFXBlm+ZNLdvbBxmQ1dZYr4MqioGOzDBOUiAPxNI8fY9CUdYJcgJBSKN9bcLjl/sKAH+KcjN
9FUnIkkOFmXT5LAx3hSi+Ep9g5FFGSfBCj1+CDPKnE9uybGRyrJCGQmhB61pdrLq5aHJxfR3z7Tj
t/OmUYs2PIkt6T9fWrri+LSN/V7goRwYIu8KFzoAKFWUxnOCO/HTWs1oOKWqcHHbylI93cNYxHOH
f/NsRWKk92ARqyytZuGzTuFrX7Thwbv0FQuQfyFQKbw5bxwtDwiwfaHFZ16XE+Fs/H0x5uIBSsFh
Rw2st/arO8bomb6PmQvM5sQEXdpKAoFFaAU2GT6j9rZFeALmANbGrC7Dm4ca0Z/9vYqUsqWdpsnB
eq/DT4Mx1WvOtz4QQ5DmUWe7Uwz+U3kKE9ha1fnF9pDtjm57NKyXb+jCpJy2dH2CcGy8ky0HJ2Ks
gMQpm+/3XPT2LElSF5EMJ6HJtBeE48GHMX8I7KUckNLrVSmyOoEjVDjkUdBRr6dkZpr/lAdClZYr
h7OB1T1hTZtwSkI1x4Heb05sj7H+WVydJ8n4xS4cSSy5u1rGQlF4gmTJXrHQJC+icrjA2gwPgZT2
I/3A0FL7X7qKWQWef4ogo3YKhklPQlHE0Iiub4km19wyudF26booDTkSM5lFJIEnVFIST0sIa+0K
X3840TAixt6Ww+tjHzpMpkhPk8YfcY8G8SzXX8GtNEGpSc8FpvAktOW3qhn1iUI3rFfMjwijQSCW
znipxBvW7hq2eMMpJX3pidL58YZWXS1zARGrFoYRzS4/ENh0842r1Y6kY86grfTk4ORP8oLVfiS2
YuuZT7GMKd+NmSOq6ZmGs5uDBoGPIfTk91QIC3bPUeVagr/z3MUq2RxVASEktzlMPi97rq87h/VD
6CgQ8NeMmoByn2lVtQVE0xsvgRYdymwQ6ycPdWcYAToF67HSMdL5xXsJQu/VqMliF0PNRSoVuiL2
43PmegY5jZ2xO6lUtctbACiLpsKCJLIsDLGSB2ACtvrYmBhN5jsEfdVBpTo7GPTcYkdwXB3Z7W1H
CnX/vhcgBRbELDYmVcO9vySdVefVo4+Z0SVynGJKdj6L+uDDoyaEQX50y0K/33Ck2QDg1uFqCuD9
CsHYRbPEE9hMFtEI9b10+sB/YUizQdk1QzPlVTYz1XHtDFC6ilRXRd8/jut/asl4vwXObSrm1339
MnDllsowv+3J/9hsdbVvm3RYxW0NcqkLcAKz4MNzeig79A0GmXlzK6EwxtlL5BzJKueocvLqkPGN
QfRMiaj0IKCkdcoanqIkVv9Sio03m8LNRIt6HLwiNJe9kgVd+BqFAPUircGC0OF1/fLs3bSW02Mk
WekwfixTeqM6kj0zG8vOMyWuR0VR9NS42SeJAZbXQnwZhVc0hWjqY9qJVH22Hq/wUnWnYEort26p
qePeB131F5D1HJ9VeZKINRUWX51N5JuyqPxgOENsXIbU5Un58VTPJ9MpeUmteqWS6kwjNFIgjyiQ
DHQGr2p0pz2Of+nDzp0OLCe/ryt+V4/V2uotdAaZ4Vo+xm6hTjdZhdEZNOOfCJDZCYYCuS70w6H/
GC6dpo5b4fruF74EClie1UZKszYMdP09yT2mDLMT5rApIJ4oO02x5ktMfOZCZlgKFgpMt1GjDQwK
qUJiP/bvseHClbiyJ1yADfNu6gVDlAmUFvdtUsRPSqveNX5n+l9CrLQDUM/p2cCiwORN+Bzd7msq
ohck8EY8MV3N5HcKSssXm/2drrIgTTHapNWMx+JYl4scjDgDlUPofOa0y37Jbsp70itcoz93lXs2
Btub6LPhp4XCKtYfFEsY1n5TSZwvwptlX6n2XVoxbumsmV/M4OSDoo5PK35+aiyzUbb5oXh74caz
n+gDQJgokgUpz4/agZqffDJAzW+07yup4vvMjZyHFshqo/X6layZ9l2RWTIPkMNvjOCtXNQb5/WF
7VoH5o3o0WCLfLfTmKA682fA9vTN8NzEgNSRIhCVA/1DorKVngZDmjLHKfyiqfVJgx1KVqyxIj42
wVl17ZpMwNAfALWKTKpjZp8UHq4QuXgUm+jY9SmHhkWzfuZCN2sX8YDbHBddu+kUi+TIL8GZ6jqM
z6xqwsoJLGb0Waiq5ZA2tPX3BFcEQjGoNfZI1i8ZE7HtZyajL6maDNF27aIySjq6ZYptNYfdMevn
gQhplhU1yRKG4M95D6h195mQ3m+9PYqGWYvQPKr/xSGV14xxBMHR1S9bCvnxb8SFrWb0Qt05o4E4
9UOUQDRoZ3W74K2UF6S8C4GDECJX0o1uwrNWc/9ywG2pvcvY0ztmgeQFw5zzjF7iWZHOVWpL7dS3
MYdo195ZL62URXz37vGTJqRB1Ey3+WITjMVlGyFAEBR8AjiL6+wokkkOw9yhnkB09SArVdHxcQNg
DESwxa9ZROuZaYqDNKqw8D3/1c39UNPWJTfFnSelLjEltIR3ZrrH5h64Sl66eGJ+wSStXGlP/L9i
skSGGZ/qL1gyMxaLvG8mG1l0Iylt9YaAN7vE5610GacWdOXO136hnu6v3r4fkuOEo/imBcKmZYWv
3gT2LIRgXirnPScAIGYXH4khTjcuXXI8eq6Uih3xxlwuLv+/OKGEFrEW0weyOepwrkLbtGIBoxrv
yGYOcsR6H4XugCtgQRLvUBb67aC3nQlzzO3sEt+mc1gtZSQEdtNRIjHhjqRpXLgzcoB4pXNNN0op
A9HENRYhZWBaTipTn/kSBIx2w1G5mkiNEnDP1M0Np+XnUCoRo8iTopgY9IZsU6tBVkVoXweIdg0i
1LWVetLh0SLrUT9kpyD+Z3YA33A2+ZzHdfUwZIpd5wLSLV+NBptjhal6so9kCN3Dcxe7rb0PuLOz
z3uD7RJgLfeDRetxl219ubqWMoU1ex8Srh4F3f9bDaYxQvFsk/l7ywQ8tjlJzT+vtu3xX186N8Gy
oTL3oFijA/WkLNiqV8U1KIeNBnpddlmbGEabM0kygdJEKRpOx9qfwJWVs+ONBLKqVVhdJt7BhL3O
lhIcS2b2l6VEwEqUVFW9mXxAeMPBM5+Wb1iibE8+kezScvGi1TZDbE98L4gEDLssKjG0Phr6XpLf
2JqzYzbZw9kiwRwOZ5y6vCuvWgoZxyfXOtRX/Lj8rBjOJ8sYivnUd07ZY/eb63VmthiZEZyrT0Kr
fXoLZD3UrvyXAI9vrnmITS+CkS3LtP57/tBcCk+SZHhC2I81OVo1Skzm5um5dfXr068KSvFhS23V
/I/LgGbr8I6Pz4HJdYczELUMf6r9ZsrkZb72DIHnU/9pKM7A/TCb53eT8N58nQLF9BzGxkY3aKxu
XwwGOEM8K7pW+ly2FFGP/kpT5ISqm+T56aV5W9W/ZYz/WbROLaJO24gkfuHxD+UD9Qm7/aHVULu9
rcWGqF1TU7dlU13kMcAfvuHegEJ0XVb3LoK7xMGBVOoPP0ys+HEKRToS9UwWAYlD+ITSHhsMwfaM
EZ7+Ietnl8AMUVRssxSLBratxzsztC2pDLAIa+tzSoWxzhNCbFMOy3vVoOlJfVBNspgLwIaiFkvz
KRivAxvEiA9iRrtJOMf290RP4HXsOJ1mWjJehjZs8mdF2+qJXiCFDPuGuhUQbdzfMX1banMXN1Cx
MBu51vQefkOuhmNzlAr6pi0qagflYmftcEjl0M0I9IJPMxZ32NtZBe+Tkb48/3Fi8SiiCohR5HPn
fsKbHSfxOoo368PDhn6rXdCgPTD98CYd5QcuspSQ6WgYh/Z6Ymgei5hs5RsTt9AOlLpAr7J+m7Cq
5CVJBHQKXYAYP7LBaQUALx7IREKpC26KARWJpib3xX0r7vlsp+mZk632AdpAyA3iQsgHrpiNoS8p
HQDasJH6ysq7t6ETUT2R6NoZQDDfvV9rNvx+TpOBoHAogRdHQsJXylBiTkHrMuypEoZWQ6gEtGXP
6MAOIdfQgigcQxV9P2AYHxDUWvsFZM0BlEs2+4EmAbD7MCgjHC0oYOc8aeRERLsTI0/9UffSkQIR
Hr5N0QMbevXJwv8Cb25sMGvytDe6cM6TLHsocalHn32ysINEXyz/WdsUo0TRhmSvXC4wo/hYPo/t
iM1hLeSnrlGV7aTvtAkVM05tVw/y+h8rYUT1L5KKfCcKqc1vJxdsY2MVWGy28Z6tbp1KjWNTnKDd
NBuVwLm5FqdMBZjyplq10yUr1WvIrt9x6pm3OF1MI/m11HreImjVwTNHIDZxE5+dB1z+DLfrx/eU
S7fFMYj1/XpTR3LLwvJruigjw2oiqgQcCIRrpMZlBBP676Pqo4KbhHc2YBU3LDIsEPgFNOErxzz0
JkEgHTv0adaUrEbtoAKTT7CmjYfeuaAxcMY8w/zhBjuhGkvqVRIfmYOiksaK/hik4aI7C0DH5nnF
SgB0dLerfsSVtUA8BxcQAoDjPrSiLnjhrF1Hrs8wzmqZ9RQYUm8ICkwWS1STRQY6pJeh9M8QiahN
14VxdTe5jJs024xnteCwFEFWcJnPfTAe8WcqzHd6V7GAMDO+K+PSbm1o5hQXGF54I13G4dIogMMi
1gsHwcJLKQDmW3678CJ+Maeh88ovj2f8lBIcs4Z2qAfuGN4g/h+LzuTJdI/HfB3DvVbmz2v3PVHB
+ynYkLz5mqzB3AViZJYsVAVgaPJnN/Pau2aRmL9o1aJF/6ivO7EDY5Np129rYJsaHB5RSI6zevig
AFk2dfhDaib3WLldg9TRnCNFv0ZB/n+RMWbkzf811sf4wIQMsdn+WLTfw1D2LvDersuq8BR3SqSJ
hMsOit9kVpletkiz2ctfU3BUcIZGkapQv5ak4IdER73HcI9wZx9UJWk+B1PsNWVCL0zZ9qNshMz+
flmN5v7uMSx18/GGnlBm4Toqa8XbtJ+DdipgDC+cmlr2bFuG8V8GQ/RgtVCHB2fEbZTgELKrkCta
v4wutPCO3CK3kERhS295Qfgq70Xm9zMo2aDgU7i9KHNoFZ3L7O6egncJJfqM+jOVi/FHgT+a3BOF
n1BEyutvwy+3bkvt1/L6el14boK/dURpbhe/XBOeZmKyVQ/an256Slze1qLhLdrPKl7dOpg1pSi3
kA95zDUTkZrthdfIrht5ixML9kIM5mwYEwiSI/9aTvE5iUk9VLvNdKRKxy28hppbPFjE5+0dnAj5
wyMv3op8G/ZyKmIqBcikqKarPbBtr1FYMsb4aArTszv9X7svKnV57XFyL8PwB5XGBs3W5J+Cnkwv
BBMbGqEP9oTh+h02YJd0SgDByvvrhL5QMxHk8I3vB58YE25hhJL4E+TrJnjSulDGprw+IxwloEpK
y3K3lPBndCzm4RECmGiJn80sh4PlmCJtKvROKn2FrCXAASgGq0FGmBnGq0laLoLnoq8WCaGKQH2L
Kuw4bnvM15NdgPSMRzKM6k7GLPTtOJlILznvyGm+mHaq0U7lpxSNiow8mWM8saQqTE3JnNu80ixN
7TCPlP/sG4I1Q3AlO11HJUx3sEKPBhVuczjDhK+hcHEN3cJCmTG/iSQGG9kMir0uvbMnnviv/Smk
LdWk60Pd44+59KtT86WsFiJsKqFWr49GYyQVAJ15GvXSREZKpE6uSMaSyAucCdSoknGWouuiBVZi
ixNzCSlL3Igq1PT3l/AOOE9jUMThQIq6tOCsxDNnocJ6nOEksSeiy90ZSugDJpN2Zx1pYGPYKt3I
QA28ZP38cditVjbDOQwzK+4j7stfZ85d9sQcE5iqZ6pBaQ9EbAqSa4pY+fKcynuZSj+hTseYaYjM
yy5n+8xgyO+lIM8OSyU+8FpLGcaJ9+7VVc6K0v7s7p6lFrn0pWWj3JtKkaYlbl2LxD6MyOvxpx/r
9qE9ivb8DFKfuuxXu675l0grNkXTUm/BznOa17xFqJJyapJJsXd3miS7f8WT+NrsemFszXOF+Eps
BtWnsVRNWQRFDeDMoYU99tDJ/jd2+mOPXN6M/tvdJvUlc18rnF/oI2SRHZnxUtgs4ebD7HwjIKcK
OFIg3/vdzE/pnYcA0KIvSZrky6kWT5iiWwBce1H1UlVHGT1mvobBnbWUkrYdYrDx3h07fhBixEpa
8JX8SwbxEpBIzWUIz+p2QYX5xVffRCmfNnSkJJEvn1k3sZI+y5Hj/VVK7p9n6jCjZ7CBUubPNGGK
4GZr8+ld3kxJExXNwhnhtcUZfaeKae223OszRufnIAZApM5s7lJ99iCFbFGWWQK2u1H7jEMJo5UW
Ie5EM2cSK4uq75TdGJhV7iV/N0xM7KtB2L6eW2mil0eZTMw6Zlv0pRgFhx9Es93D7Enj1slxgPyv
lRNND5BEf7YW/SKGoQgrTnZcwy1BgQtHbH/+SiM/mJcKO3H8BCEMALfXrHId1WnWWe8tvSJWEIhj
LqxR5f27cNizMlY9kHZEbVUv1Ig789y1kdUJNFB0nwDm/VChN8SqsC7JtIVyexWccWEHovPg/M8v
6FFn/0v3ucEEMZreHP2UJwKQlL5//Yv5aZ4ouNJa3Ce+Xt65k74wg5qBG5IhzomhxmEq45SGt3W1
kGtWLf2ghcvBtUdI5QOEMKHWOZ5VQnWYDRrjtxAUhtthWHkiNAsaDiAvVPvA/gsr+mxInCrSA28V
pt0YUgEuR0a950AmfDO4+G46XWSN9hebEuP1bGZ2i3S/oPIc6TlTDsQMrPn35QRFDRiRueUSToQn
IGJWEOWPdofL7t9QVQXnphqtDgWtR5E2CUpfT5NcmTSRhADlNdGSmnSpCWAZmxf/o5U02jZ9JVgm
o7DuT2PJ9VIsM5u1DB+asmg5zUUs8dGbvyprzQWr/kiJfRkdeMZynkNJx9zeFeO/e48lHy1JL5Uz
bt7HVM4G9ZUNAu/gM8gK800vqb295VRX15MizjLzvHGoXLIDi63NG9vUPB8leBEZzCvw4ArwCuCu
CaOdzK7t/vQoqsp5p82UyfuwMpW4kXmCtsR2+AjHcLF/LWCAesRzbXOkprFGPRnIlDjFwtMuW1KD
XhqwbV/ITGqhe0aSkGM4JjL3OT0KCekuQH5XLRTjU9emoPtrH/Bbza0XMCPUNU2Xk1MRGpdAfvaU
RmmgniXEgfzswiFHxqLrb/E549MQeYBgojMtldJp1dnxHuOAdCOI6A4UGwMusqgqJc7JUjGVx3Cl
qVQkSWLvFvg4JSJipjt0coOmNJ4t9Zn+c8fUpgEF9nyAgJVoG9NZ3fgqAcpObvbdq09y3CGRcVPR
ap3ifrFEpTnQJI4kLZUYzwWzV6umd+Qi5+v/y+trD43s58c/YPUppubj42SfCeBqcDvWjRtTn3N2
C/f+pK5EmUllbw0aqkStIBOFay2BTj5aTPZeVNNu+GeDVdIpoyra6zNwCsWKPWm7n2uns7IWljVW
Orh7Nl8h6BwBGLWJoukkhdNNq30FOaNx/T7XoIkIqIzxN3eu52IpW4AvQwqumur5pz8Z4msVjeFi
mDaL7XYxb1TEOia6xluSZTRdMl5p86FLA1DIJyvp8uoRV+h2sW+yJ5kx3DYglUccCfmvGfRVQS9m
bF9FWiAx2qbSYXp/qGcHj9Xoco4NqVLEwjDg4gVVloWfzDtvSPxsEjZJCIvaHQl6AQuyMcclV/XM
tXUbW2du4SOxLkbVF3fH2nLYz9gSk8yOSxV4tSAb/4J9Tn2bJQlbLxbA1DgseahsOV6yO6+xD70G
1Iv6Dbbbus604gya5suqpNIaMdkctiifEYe/e8IiLHjODJG/hL2FLYfvHaPJ+n3HbSTo4xlqD5bM
J1MccAX39V8+BROXqT2oyczMagN05hUN6KaN2EvBAp+aie/K0eeIZlKs8qmRUR8GAuLhQS9i82zY
Ao3H/viJY4b9QHluVpdwRUjKcETjbI5TLqrGHBdOV1sq+D2Y8LWkJjyUaATugjgBdqf/9ogWmkty
oPspHsMoGhukqax6mDI3dwsNqCpMOlv3MCzbp7C71jUPBH9Lp8U3lO/SKmF1mpA1GqfCCsqWr9UX
OALCUUSNEiDx4i1mdG0ypCcWmKMb+zofoaxTbjfBhO5Ahmywv8nbYFn7xpRfUA6gmG81N/eILjdj
6c5wExu9YhOwXaqjCCwLO9Ln4zKz8xcGaXnfTdHrLonHJxvVBQ8prOQXxjr+WQ0XrAnX0jrnBe+4
U/BLE+QUZppDo2rmu3AbHr7v0k4gBymijgm+G60XgR9O7M3NEsXoCQ3xOomlE5faSfa6PppIeW2X
1zFdj0XrCMH88X/DPQo7ng7zGTKmNnzZndlPIaaB/JSj8cvwl8L0jU43rGzEFUJ56RAFNPHhmHsC
vvrflRy1tibkNW6fjrYYs7RNtJ1EWxn9tVLLTXUt5V/Tbt6DllTVriVtGqPbRKmg2Z2/+iPbOk8h
jCc36Bg5LVKelopokxKW3MKEqCW2bDKQGIYcagmN28R1aJ8OpFZ36h6C9ECG7G0nhdnJ9c4GlVCF
3ubF+odqmyuv9G7Vyy9JYpMv4d5ygueFz+NHtiCEXLYF+ZanIfq049JTRhSn765F5je9f+L7aV88
SYbUVQIx5hku7rq8Kp/dD5SIqGo2Mxt7eBF7qL2YBDij8+f8d3EP2akrjJacTDu5H3W9ic4NHYUX
vKaR6edjTTFHCIoCCpe3pgAnTizPp6vM7VhR78GynFn5rUaUpU/2llLRC+V9V28Du4mtXfoA8T1Z
H/QEmUtjL9aEtl5tvrgy2PAFXoCeCvU3yn63AkmN9M1kmcWldRuVRmQ0wGM6ILSiQHxZMuKD+hhz
3Hpes5khFMW9ZhhpD5fFLmnmej2/Ovi42RlTb9XJv/e+PlPJxWKYu46nr5pdRruGQAhitVym9Cbv
Ex4YWhu7YUft4w2BO8+qEiRImiobMthBWiEXjAvj0rTx3EwjcRUrr2CPFSIE8eqK1KH5DtTBw1NW
uJ8xrkcrk1hG8fYvi4bZjUESha0ShjwpcaFjvUEkciYgQqq0MQildL3Fc/ofj1GW3aqJSKLYEJW4
D29Gw+mSQM3OIuIVNC2MdrYvk0ajxFmkkn/trM1ECpJAd4L6Ff1tWTZTFuGtF/ESQhYNfEqwVCrL
COMtlvC+QbSMlQLv/pIfnun0H9uMqYP8kOa9k+kUniImpR4xH/QbQxVHwm0nWPnyY16aE5m+OERQ
l77HPgGzWk5pxSwXD6Obgj9erk/XXschD+92stykOfKLl6A45SoVtG3ujNX/YN4GMCbJg5sv+mMP
wVpmUBPjZCAKv7QqKfKJcI+yrqxOi0DpbGiIbtlJG5MbScqoFBSuHTk2sC3CitAQY1HA2LEejJgk
G4rZ2qFZ15YqmMe1jCaRyEDRxU21XEeXIXv5CrRjTjpVv6Nhp4KoDfFQU1Ae0EMzv/cBOdKjataw
OXCOwi2IvamdSp70b7gaCVhC5t0UFelmd6ZLP+ZlJ0cRPoWA7/oqw/AqAKqOgwyz9eftAtzIIAG8
d3r4sErxaiOsiOLaITnDJPfs63HR5N0W8EwZ1KBET9UNvdnN90Yca4MSqdxflvy8sQGGXL154yMC
6JXG7rxflvw2w3XaaiQW7TcU4Ct5tlyFmhouzFaysDN/0irMXe53bTRDvqlMn9k6d1Y+VsibH9Qc
6ZhFOeRN1/U5G6NLjKECzKc8JeXJvh3cYreL1SDffG7TPbhdz9hZ47klUkv25v+UH0ZsFVpgy7Gs
Wfn1ZGp3yBdviESn4HTHh83FdxV5AmXAGHnYxWRwTPskCQdAfagbmXhVYGFq/ex1pfPn4zV1lMHC
8CFYhi9NFafnsfAJXyOCtT5L4LSOn/DGylvFtbcdA7bRLMQbd+3gj+6R5XThw94OSOI2779addGj
gzrLmT1EFf8ZkksA/um8o4TdAXFxYeaHexJlLjrA5Eo7H0bTXvk0O8+n1JC1XkvZiLB2TcIbddt1
tAk61owROQeHm7bm2zplIbuOw/ofkFhnyTfzfORmtGQSpTMRtBNMzp1otlHQ4P7YfcsIykld0hry
NHwR6uwPf+pZDvHV2MySW76avb+RgyyIbW2wowM0qH+FQmvHRGYdQ0nHq8yx1AC9QoSOhlEeEjDk
19wTtIry44hC+9OC3pgfUrlmvXDjmQMRrBJxD6Udi14HBAGTCixVECOK98heO4p/mRcTU/Y0xlWi
WwsdXoIeX0M/6a7O1b1j75pv+26uuNPlZU0WPPu5EmdNt9wSNVkLYHIpNyBOZh2lQ9ocXe39G81R
VFbEMSIfxHNl3Ww+LhpmxPWnT5N6vQnx2eDhzMDBanYbPGOwjvumhempV8rCmVq6oFVevoJypppC
1xO1yr3JwxDWPMtMIdxNcpU2uE0m0qXLB5KiZWbN3vqFJUwDWFhCbly46jhwkfOrRiZHuPF7Fqpe
5tSgu04VqHQDW/IrnJVQoiGlEkj5axNjQgUIPvG4Et/ZPIFoXYlc+EWCojQFYJwX130745EGwhOu
OvAWxEZNrumlcJvKJ/VAEHXCnifbtiRH03pPoEjv1TNxGgkZVFMHPBALfusy8cgBZvSiPkB1I7FG
J2hev3QbI53Z8yc6fgu62sjywfLyFEGstAW7sZ81KOulchIt8qKBReSCDV/zikISG8waVrW/F3Gv
2p0kmeTgkf44bJqqDGzSt9xuoTa7pPpwFH6CPUyz9t37rCWs/oXIA1JuQO4WyqikHrHfg/jyU9Az
uoHmxnE8Oi+ojWzhrbDAwRKYX+b3RSonxqqAwLJSkXsNXO5lyhzR79rre3BF6kNp04zN6jcAZa9V
ZqU+jYx7kMbGWYgU86ECq/VnZG2ru/TkhnvelB4F2K0kG2ct90qOfPc3OTqx7QYb6K/dev0cuFPf
YgCVreijAp54x+rrZniIe9ICJyoPWSWC+wqrUjojIU6d2ZwBP8lkdypbIrh2rSu0PXkaJtxjEbWJ
xs0eSN5VS5gIyNoHdg+vGiAStvMFXv8rt46htVbtLarEZHnWvIL990ELTcjSzYcO+R+PHSroJ3PW
6ZxN11XQtPwIQqCQQtvHJhdMWK445oXnawcWsJ1gU7EtLFMpOicRJOb0U+ryHe9+ylAvDNyH26Sv
g+UFCwKaCiQok6Ua2xFob1KJ8L3i1NbOHDxyttKtvzkrxW++Y45QysRU88/osMv+0eg7H9UppJAi
ok2Vp0qj4ZfoeHFWz4zWwdZ5+nk01mKqZTDDk4eXsGUM3cvC/9ONB38ottKdxNlcNCRXWUkGtEvG
G9E4TaFwm7oeBOH2qC6NH6rRASuakHRx9vRyuazezbaVHt3ZI2VUDZj/pDkfQ8lFeOnRCg294foZ
5UQhlrpAlzpOlU2xvnviQNZlJUyXlqY9bQZ+8ORpMvHln9+StK1QiudwYFMVpxltreVuMYTQKdhj
00P8tWtirD8zvxZrQZg96BSh+xaDQWvZC9kqLrLOGMSStEAqMgA/Osp9rSWsUN5UCQ+y2PkL0L+y
E/DSFr+oymrpgVWaaLZ/Isw0/3KoKhi4Q2G/z0lb7WjA1Gj+IptvZaKWPv5bzxWBXcc8Mixw5S8w
i0G3UcL89ToLLuf5mMXMyHKJalTmWYYzTGqb1blRAWni5B0EFoWuDVm//LvowBEOXgBcw6jwIzqf
dQpHofnspgSCTnkavcR0EQETzwyN+yGKL8hGKpIwJQp5ZLkge/f3CXw3rZBRztJa7dWXCIkHb1eU
6i7VTbJRsddigXc161oj1U4jv8jG+IlxBTDLVeXyxJZOs7z4jmx+zHRMvPRhEPQbnyyLRY2eFI3o
jCbwqV4ahyFWYAskKzSrL8MsP4iPWISMKMEOdVzeKruhV2mxZ/Fwy34Ntx0xIFSR9zoiAhDNA6dg
J2g29cFNwnfaZKyApDnqX27M2g5Icc8E4OMCsiebZ1pwOxziJJarwIPH3d37/zOx6HCZKQGf8wwE
enhvXtvJFoFAHMWHAHfpuDNDSJ+8sZBSvUGkNM/2qqKThq0g+cG7RG2hhD6wIIglaleZIkYaBHcq
3xug3uCla2DilaM7DaSKB98LFQ8VWtqlsI41FNnMcSHc71BmJ2Z2mgBeuhxTsag6+48ohlVZ5Rwi
K+MFw/ZHweYJi2zdO8dKjcBrejAW7HcnWqeodX9GT7ibqTaeOcOL58glLZwHw+9ZXOWmJvoFxWJp
uVpw9iY6U0YluqfoFokomUQsOjQkyE7mLAKPOCWFRBVCoWKFc/tcmVzjUnQxqCs9Lr9gf7URtjz7
E2zoKrmU/lWM3tHzmh8cn3c60FMAR6GmAZIHmc+9B9DMJ835CtiWb9Vs5p+T6eAotogwWlrART/q
dlzRBKkUFZDuDNpJoFE0qYn1OyYp4ulr9i38TbksBPjY2xpXCsCDIqft1TbUFQuN72iYiMSwgXz6
ZkXysKYbLTMPocwVGto5NCQNe0ehO2IPXSYiEgXD5k589V8JBCLGMHxyYC0eIl/lZfSLMDh5J+4X
K5jE+2ThGnxKsRMn1UOpsaNUTY6ZrMdZ+wJjfJt1ZUzNpYoWaUcHnU0VkoJaKINsSMLZQpSs+orW
BdMdXWmpL3DkO6OsT9Po3l09Kp9in1tyaDWvaprYoMny/SQlJE9St9ZJyqox0Zg0fkOr/eA2+wsp
uRNavgu+QgTSzx5w7LTKGVMkWFi7mn3ekW/7/swTJEkHkSHlBsRdJqA0oFUWqkQxPcpw8y7Y8PdV
UKB1NnK5vdUgjeOogrMyS70/0hwUzPNSzstIVpoor5M5qdGvD3MElz0+bAhld0f8VrTLvdSZehs+
pVgeg+3fwp7aAlC4KhAss8as4SjwuHB6qCytPIC2PeUg+sac11tCjN4JHbREzmnE8JS7uCcVC1Po
DDHAB32mjnJkpmLxqFetg2Lz3Kf7A11XQDLu5rhZ6gfPN+iJzqBNBEDb2OB97hlWxzM8lvKrhPML
zMr5KAD5Fm4B7bvh7r+8Dgqv1GiWGX+hgNjgba+w0zQWCbFY5UK/WL4iecwEyxtEGa8wKmURtRxT
Bp9Xp/IkJ03QL0s8E795BL2hCmbc1eq3e2WxrJKT2HDzmIDGMFqL3VUiN0jhY1UwCdyNAFm9632D
y8JdWD1ITdGBQBrhVFYA04QEHzgHmzaNcIIarHrDc0Cm62Cg2VcW9vnKcf0x4bhDmJUkdUHEjrWe
SMBzYb7fj7EknUBkKkCDKskJTb7od6ia1vJfvih/yB9hdP9+PcOvNNu2KT6pVJ3NPhmS7cXq6uiF
4wsKtnwQyJhFU/jGMkEPU0jRF6qItIPtZZtn82hOxfH6AXgmFb+Ng96G9uxItIhEM6FKPPLWu5je
eGcSVs/GVSfz/zD+d5LkhiXpSWdTjxKLSVtVdRO3jaQjFIZKhZk21ePqCGRASJMyaZP3f31d3pjQ
ycrpm6eWZ/5W1a1AlMeXiMy7P3kKLtm+sDiDQrzxOKtKyeCILW+A0Y0SFeQVrhRlAdkppGdr72Th
JhNGv1nUM/RYC2LotUMl/4L6QOZ6CM9qeD+4NK3U3irTpojD9oh92xgiVc8I3SEpRUvxSaA2Tmgt
NWEsvNRRo2aFBFnCG6JX3T++CElTNBoSBK5esEdiPYcAlFpFys9J+gV6tAYlnIz7o+dOo7Tg1VkO
J25HDV9/l6sPRaBP25m9i6t38qZFTfCbxmCzjcE5Zqa9EDDoJl+1LN9bDWNzfGWB1lsXVP7h29DQ
IlfM9kAW2dn/6i+hb/Sz8jGyRoUYU8WeQynkFfXN+hBArYRt9gO6q60Y9zPy1lqeQCHhutAGS7hL
Ftg3+CSuPcBe4FGWUo/ybKySDS66B7f4rse0Jz6zMYHuLUtqNWSQ2+w8GXw5g35TtZiXQv6XwGb2
tgL3tyXKoT6UWgR4ublDZv8fMNTnHH/Im5SKbhDzFmDvbMByNqnAGMIC2f0Kk/I/BQtXuvRCmxRM
85Osl4JIO4zTjBScTFdC/il41pIRafTkov1B90RDZyyyUKQVQNFaPSuuXaomnoTym9dNECpMPtL/
/rZxla3gf//mx1Ub8ISzIzuT70mmFmhjbSw5+6nRnBygJcCeOCP7IHse3Ulv2MSROK1VaKY8+qZa
aovoLeY5PHGe3zH+3EngmxorEEXjz4c4cHaB5Jc/4nU3QEb/HxHRjOBUoRhv5VFUAwPZtcfBP9fz
HqR558t+LsShjwI49yuk8OyTT54ByJXZPw3FlrvwIboPQjI1CVUS1+hmN/0Nw5TqUVhBcY4TVZmY
BrcKRCfs38FC6LIM2eNYnUBMjoV/wbaCyrCfe+pPKo5HI10ilTj6qxvEynUxMixcFyWl804V1ZBS
DBWFFCpfhgXuMDT7Na/Ve4cH3HN+rp0SJpa50dgM/ASRVjRtBUnrS2bFssrjB7vfqBfKXmSDmpr3
EqgG5NG8A3hMAzpcfMDMLR1eGTyIdr5bN9f6CAizp1WIOhHEUtMSFJuR9MfxodH4yjYCpZw2R77A
3JwJUB/mLBdyedzF8oAUP2D0KGf8RNxX5kCF8AdQKhwBQxzsh4s3jTs/uolD/qq9Exw66/CNJb+l
3A3GR6nmVeROfkoIgzF5KHaT3tH97ZpHSyQSpgb4i/LLyCxTT9UQZDQrvrTKh3HdDeVvB+c+RqSz
95kwLQvjvqW5CmcHTRXAHjKjztZSWXg3jBo5bC00giTob5Ej7ygp2/GI8/Nb6bYwpvbfj7nw/mjG
ypjNcyk3jK4TVBcMEVd07YqMo0yjx6Iqywk5gmGitiduzXokf0HQUSyTbjbmctvMGnwukL6rgdM5
udo5oFHVIcVDfF50O61xyTYREnXZe4CmmcHwlXqn36Nt4rzabSHGtAqaL1PBF2ppOpOsXFD9nD0i
io9D1f0hnxKCd6U1BVYzhdouxj54yxLurqzXmxjBrqDZkW3iX4H5Xtjzpv/xyte+B4symiuMJFP8
ebiQqjxsG0xCEIzC+V1AFfduLeylFO6FzqwK6U9HoB3guDVj2kscvKwcnRAvMR38aNiINUwT41G0
aKUBfSBPE775rY22DKndJ+Rc1TzfInsmplQgh2CxgMj4wUNFoW0ppqF4G5OFI+Kg/PABMgIkeO0f
Fy8DZc2yuLdwOHk0o7lmdrF7Hgau2YNRrqWeF0e6+7h3Ua7XH6cC489nofSMTy+e3X3gZu1xTc0u
Hc8WouwFWvGk508zTUUsOVVwM+09iV57J6SlLdzHzTwS59lqeLbJzeDQ2m+/YpVp60n2dCD3R8nV
LLshlZHr7q6KjykHJx8eJr/rVDBu6ypkxxCIrOuo43+GLGN/I9Z93ENRgmmdFuymCxi9wBKiJvOi
J+38P0TrGvmGA1lFQ45dp0hMRuKbuq69ejXRTlkYfWx6tGtGLOFAaf/m4HeSo89HLoUtnMdNGiQz
GtKn5uGbnSmWGHGlnE7jhNCv5KPxu/Xp/SVMLBwGnqQARwGy6DUH6CGlbcolB8CuuUIea4nzDCT0
VKlyz4y5cDu4PZYWG+j/AD6Asomtc9CucthoG9C52huPc0AOWH4G06KyWNEmHtWkyVSJlLKDyCvE
v87n8SkvXAjImiMEqJHE/A78atS2mECzdoq12eL5xuomObS/OiWRkNlx5Sq8FQFBkJNSLPjdwTc3
fgMBVy0jiKHMAsTf8k4xYSb/PlEQB39ihoE1q0172ZIF5g1Yhog60yITYWBfrAaPC76LZ7ioHYHi
eLYH5aLDSubxwDJfCQJLL//e/ueNqdbN0Oeco85D3Cv8JlE9AjVv/lTLoFuseTnnV6WIuCWRis1E
BkoLmeqjmrZ6nGrTff33dn6sA3D296pVPyhmZIJqAMKhKLdVNwe831lmY0EaRvP5aXfzq1ju0VV9
JpbxSdNQPEnL2oOlW92p9Vc8ef6hUnufl/kx6tqtJuk9k9YWkJkr50kHrAaAgU0CCCHtpGhPmEZ1
W9/UAugujvfBfZn6kg2oEQ/DtClirzBPm82g6s1lsrDxsvISR6TvJBaRSJJGc1TbF22GZASdGu/s
taYRDdJSyTpu0d2JutkwOKiLW4LLAU5hwaRM6mYlNFoGu4MH+ZH9vQD/GRg6HswI0f0koaVvFxxl
A7dnveh3rp1+nr5JRiz6PQHASXXd0cVttNJTNZL0adTo//Hf7hnwGsY7o01MmLVgSwMpSV2h9H+3
HeHkkOvn8IvxroTFUibSa5A2hhhz5pmJnE4oLhNX/Z6FVIC+WADxtXkZywhd8qjSTi4P1lcvH2zn
EQZwLcs0hEbvqD7UfE+mI5pOidtIObwO+pmw17ZqKLwiLgvhLmLlXKXndE0i1F1YOrDKYIOf9Xt3
FpFbOjrL5qQQJRbpjZXRVo4AgLHLCFIIPoZa11eRp+36G+kgVEbWa4571NSx7rZjOhYcyPTkfBIg
57kWjZuDpVt5yWpNG3GqG6Vkp/Tc8o8+KBccvRbXpUZd41rMs3FU/BHp/8zJ2QjsAHn+VmXiY8dC
9/4/m1Ys4yv5IofKdsRB8rYSebe6GqZUycIeNHkBiHojbDaP6iwRRmYmO4ybpH/dO8BJhEQN2hnU
EFaIAQJdUUUdn3CLHaHtd4sCsg+NoyKYWPesLMcZk3S4CrhOIsxAlFE+vTf/TsRxR5B2X2ac8GuV
MI+4XPYhRKycltC9ge2cugJyu/crmNFHT5OiDKdqEXEtuhYFmD5eN/gGW2FTkiAZyA1UA780hjCo
oYCazd1zdkERHGFeBd6qMWzpGM2xckurKRm2/H/j0qTDjAf+b8NNkp+6HWKY+sE1OoMTD/DakEgv
YFvD/0IGs4u3TeAy+nyUheDXjQnr84D39da1uuAoGDDHoc/U8/RKkGBKhOLcOQRzZRJXXLl1LMX4
bFYhTewAhe+qwgZqtAPYdrNQSm1EYtkyMzarjEmP7Se+cZmZ9RESLVyIKcIqPemeDHAiJf0XyaWv
DnvnH3onFHLBQaWGj7F4HBwV7S6mUixF5dY4WyN0nf5fJG6fFITVoJpKot42TpLKCnaEvF+ff96d
aKVXOjWVJ7QBdtAVCepWEioTsISG/nZ+pg/zXPgUYXSjnCfa7UnRgmGIoFfwd0s0y4jtgg3m+1tg
MIMwvK0oF6VwvV7D5oDtV4Fi72GtANm4R8UH6AVXk4LWbxsTfb0E5QdDnh+mazYsMaVOoRGNWaDQ
eI5Z00FnOjwD370B+Gy9II0cRAN2w3nkZnz2AtiQQDV+y17ZoiVYOWkTFnHThitY5OWgS+ETqqRC
U6HOEtelSdN5nRNhrNM9JzUKofF4QTWGKWC2b/TnxAQJGjkuyMRZ88meLHyqnISBPryr3tVKiCAW
uFpAufkM9bNGxMHdtdU46S6EGI3CNdzbPlSmlJXfLFbh+j+IL7qH9oiDCO7XZs4/Gp4hKull6iyz
PQk02ysydjUTsSatyjRc79lFLrTBOWvUHEgzi50VzXzQkwfvTwwZWpXBRG9t/oFIq/k0igzFKrbz
4LBoNSSw1px1QRsxYtDnhkVbLQqJOfZwcDHbc/a8W6nr0gplaiuGeTpOcH8QbdGWt0WkATSfiDHR
+0KGVw9bxoX2FpzuAdql1HvMiON/lAv0LlH0te0rjJiNNMkz3Rh3xXspre+CT8sf6NZVIrPh8AV1
DtCIj/ddS+QqZyKSQXYWh832NbUebiyjuigGxMHL0u6SX9UVvUR60tdD1NQUcU0X8+B+oQCF7bL7
w/nngjxjZtTbIMqSTaNGYIHmEW0AeXq+qJiEojFFMYFmMtOuM9nyFpcGIulqIhpSMl3Kdx+Op7px
5pVpbOZyBubDg+hXJ/5VkepXWL+TMIAnIkZoBcU8YWLo2urk0jOlLw7F6m7uSgIei/CwXxD6LOb4
WiB9iAUZ9chrqtLxNmG0MRGlNjtfUJWBUMhqcRbi7yY9sgMj6T7Zt9BHkOU7Yw5ObcaJfrSU842y
388+sKMMcRICwaK8fYXktCHd+si9AvpK2tI6eoQzQFq2W6M1Zn4QHWFoIC1e6OeCAdUvtqw5POUm
LmHWKCQE4t9KsIMh1eakZqBsSPDtTOQiNHgA/RcXmaMZi+yaIzbmH/ysdfFwBBz8fuD2wzEC14LQ
8SjFEAyVflRjrU5fqwC3xMyfinYTD4lBBZ9h3xRft4dANsLK+kQX6sN0WTX0ZlDN+OS0jHcvOd7Y
a0mKRdPIsGqDrtElHAqZkJnbNp5JKhh3I70LpR4yJaOIV40HPGxP3rZf9FtOyAI0a8/KtXRAbIsu
jQM5y0FYTvv3k4EStfrwUlpigZMupq1aitBVhfmlDCnFhHqoPjhngPaX4ahpgRucDYL8vJwMM/VG
TFl9mMPRuvsXY1aTeky6ml771qc+vxTnNBqQ3x2dG6MSzfiuY0OP9WWWOpcNo33DC/pcnJ+zlfW+
nu31a6gvgMWqwexk7SF+/HnAJVwYltGMy42hpCM6E7cHZNh+YUbgNbuEB2nIGygjqP+1jtrkAaT+
eeAu5YfMUKGojgBnNutAZxlYej6eCqpSJBLa65E6Z8iE5Xl5ftPqPH3S24YMI2yMJW5Eu84FcGeV
noon0m24iAavpLfFUU3fXDMFynYGAld7pn2o+aQytt5Unx3BBGhGb54LRK/yLD9BWsQbIPd7aQkn
1NpGrKm23mIX9R//Hb1nBRGTjiAY0Udj6QzdQM+UypiqbjfDwL9CUZ+C2ffgo/GYzuJKP0kinlN/
xp/B2AeenD0AlcwxlofVSuabESYs2SKDb2HoUWC75GqVLRkpBkIxZ3vj8Vi0xOA1CiSpwWDpQmoX
B/g+5F11+gmQi5zedr+1fvmrEOr0K3XWL5bibqyQj/bS0CtEoiZ8xOTi7R5uwbKxRAayYSoP66+Z
hkS6S64l8QMNzJ/jLZO0ZxKZ53lpnWjAJlErDMAvOj+TqJ7+GzdI2EWWMz38nXAnfOHI/6mCH9j7
dyuemnCmR08JiUcDG3gakoYlQF9NXbtU9oF8mp9jXDW/nVf40+MHf6AQQDp3c0UtiM3oqz8kggup
zgH2+F1Ci01eSfmULwz00DeLVanxA4F4GIl3i15vtvhJbwOR1+7M2GsElj5QmqO0zoDCJbz1o9je
OLk0tRWD4WHfcom7SYNx3f49GkO3j3DH6mFvmwQhjGFpNqbAQboNh1HDFjxA9HRIAE4TkkHl6gJR
J+cVEmmWfDwyzrmZmoydrZ5xgU8deZXnhIsmBeYRNUEIxq+xhGC4pl5ca1wav+U6lx3yYYa7omBW
DeZcGvyAc9qfjhpsxusRCZG/DRDUc4ggUP5bgls+Xj7IvZl5iDcJvUB6CKKC+MhBBv22Atg2H/v1
UjgSQ/qlLHOKrtVlF+y1tA5+N8wSeEFBsGrX5bi/33YdQhPJvC9vdSxZBcGBHsb/mDsXgma/Nhag
a/K+ZK82Zk65wBvTvY+HHGMqkTbMbpQBIwsrJu7P1XliIz+WsGqiOlQPjLHa0Lxoex/JmlZHwT+5
vcEWwhesHyKYwkFs+P8W8QhNWK71CDlvBR22GvZDvxrvunctRXgxvJYx1otX7+ySy6wnDChDGUJj
b6mRfdL8XkVu5iY8pp9tpw6KDTiTFAigBnhdrzx8ZbRh0l3ArbVDmqYCGfgn082xuotMxku6KqGx
UdbOJQLRLR2oaO2ViJk6oLrTZR/EIxTvxAda2USXJ0Tz0iYjiTSPaIkuieZ4b1GLKO7uvLoXnNtl
/1GhiVbaiynPGGhbgPxEhQ/9XaqKDxMb7JiuPWMZ/FPti46Fm8HqNx1WOez4W0J6hLT2sKLX+Lad
EcX/zB/KKWRZu832Ax1ttcze5QHR5ObHOWULqUCFo8T7wv8N0vkzMsedLzCRTS+MWHrtHJRsK3IN
fu7P1aER2EjYVNHUiS28NqE2mwHKhiu2pBaF6JZa8rzRQBKhQNHTlfZmQC3bud4SvNbnMZOW3z63
QF90z6LVowqzTZzgncbZ7+tG3DNlg1oGnONKQkuwW1eoY1716cRU5ErvjO05NuFEiSwDaMbtPu0u
awxypqrGhxDGzckCNOYg5FM0fZ0J6W/EaInuc3JNv04mo2Ixh9OO1TFrLm3FBNcyMOdY48NdMGf5
9dAX1FL+hN6kawuJc97W1qMhvl519ggYEOcu1rGCXCZndJe/UF0UXi0fdUwQOiwB40p2Tl087yCa
KBuk1qQvwXBq0E54YmCnC6VozFqzH7fZOnIF87FuqChNdAkaeT9t7JRNKpSraF5pV+7xafrIwPqU
23CR8ySypIc1477ETBfnT/JPEWtlIWfy8Td/5VCpfP8tqPPEoPd5pwS5rIwQ4LZF/ry+SJcfIoHq
3aASWACkL9Wsth4TDmnpg9UrBudJR8phP9H8+uTAra7W/Uq5M8udrhe3EyRB2MPY6POA3M5s3DSP
gkqDtWyk3C97BI1zAaN3GFFv3vZg0OMejrYWUdOkRzDWhGtr3xzrTIXXSxb2YsUrvd/gwc9vDqr4
G/cPkOgSJfMC2ePSkXGYfmQlLRUE0T42zY8p0bRLf8kd4ihZ1ZqxJ8kiVde09SnF3WM1cWJ90VbN
2IH9rvNDU4pbaRdp8BqLADeA5LvoUwURSoEWjw2Qt/IdEexhWy1FMGMyTV71xGq0QxEA9abTZ5Zx
F/QZ83c35c8Hb3G3BC+78fhgnAZiox4L60ST2snlvQ10K7oE7zdYcAOwsgio+kPDbR/5Rvfd9q+s
G6tAbNwAnSqpGQEZ6/Nr/KRcYRZ8oLK4BrQfqnm5U/yjWVGNLkmDXFz5VP17n1TxXjskz9B2sYNj
ZQvakGTm+7aSHa+Q9IEESQr8/B+knhSRBj0f57JJMVqANyuB//c84u6wcjaRy8RlVxl8u9X3M3y+
XSlKbOCaWak7tPYiqFOgOy8IdhlsCUDqx6Ab5cGHJ4z9NwWyfMJO5wrI15ZLdaTyjgn/ogcBn3+a
B3904j5ABNoHrw51xISOrbXOv/UETE/oMzQcwpXpovhS3JG6Njnxgj8AeaPMFFbm5tOeIh3RnfHP
++98iFyUctzX88/Aweo4EbyxwEGo4AzGx8zsSNAd3oYsy+3lWjTNHowVP30LEj5ULEBKDE6aMSjk
vva5JMy8zNKOkoOW4sJp11wYpyshsOoSpAi+D0KxEijNBNHi7hAu71Rt/5mJgRq4j3OaE4dSrSXG
15eUJtEob1NZfRUzq1fXQIsgZj6pqe+gZy6z1HJ/Af/VXFc9e3J1gTPillqNcYk5u9mQgPAo3dkF
qmgiJuzeiqWz0P6i/kAnrkgI3xit4mMBKy5Js1oSMk1gjwDSx0R+ooUSidrGHwKDvu9S7Q9aNYUK
a/oM8wzxcdf2u+EF1Kd9zhZNIj2y5yMOcurgxWSytg+jKrXZ6UIoNtt8kcED4poIsbMg0N3mPI0l
qehMtCQ3NMl2lNYl1JACOqSqCwEsziO8UPp9Q3Y170HD/4Ce5OtPi198WlWaOMpUP9NzZxQGPNg5
3BHuxPTn6VvOiJmaxNsms2+LsDdXSAXi0pwcpB9XGf6z1Qux7YF+EB356A8qwuy5Q22R4pnTAn+e
HdQ8lzBUYfHrNq9+1KjiBOqAC9zhaSiu0IZNHD4k5WUAYe/1Mwak3zs0LoGw803CTs436xQUB5va
/oLSV1M9tHR0UrmDN/iep0Nf0/VagD7K73tVThs2Wjid+xGB6SfcYHzM7FSpFuiEEfvAyc8IIEtr
o0ZHut2J0XNNGTgMtXOJlvz381DsoM7taagrhGyEzYiI0Mh0IeCZYhOI5eu7ykLMwEnNWzdC7pnd
w65HaCIX1TQbLdefg5n8oKXgqTrCZDiY8ti+Yegs9Fykie3Zhwfct4K33ChhLeRoAURO1mNmBAEg
vEj1v7ojoBW4NRKQBD6cv9mtdJSmtHXYpHkMTUGBI12qLg66dgwzJOlUndpAhqE2oFPMMqAZU5/j
+roOvzTJ4byla4Q6HBRwvnipZIJsENcuWsVp9rS+jRUEX+YEtOh3h49RL1C55jB7T+V4+yKstvEX
loVBCWTn+Bw0GkLy0z7CqDnW74UFAn8eLUUWeLpv7K6RnbqOsz6555CT4vPCKB2JbHgVH+l5PlMJ
rqlzYoHgePgQgLbDJP1U1sRkqig5LTOQ/sB6g07CyNzBCBokj0nohpFc5MkyohT8I5LTQnsbDuTS
cN9r8t9NaWlxBxtlfSPLsXyiUieMosVtnPcBRm9kH0797AS6xyafMZ7GaYbHPLN+ufgAbHplnpKZ
hSH53WWRWEsUjUHmmnjm1RJSRpcSsOV/S7zuhNTlbxx0pHRvO2e/8O4B1lj5jw1XM9TMSGFRZpf0
Px0grg+O6/I+Vc0gqJPNtQUvlffj9p5gI85CzoIfe4JbF7WnIK1/aIh6krka8zUwFOR0niRfY94m
bjYAv/S6CkOSrQsP/cRNxoGMwzzDnURIp7I04OA8/IFpVp95Nq4N/niNyyhXPy+wR31ZpTprUVja
lAEz8HR9oyzmbR5EIx72Cs1LME3yuWNdG1cnTWdxjq2jKJZNrP8FrgoaLCnbqKarYQtHE/LwBXlv
iEN4L6ECRV0P6laWFPwdhXNNWvs8uwC7PD11Z+P7DIaKGsr+td0hIXjgOtTcFfcw5Ex+851EjeC+
yrnJGm5Vpim6mKf7Vm1YP5O4BmGltfLy8qrFpclk8dzysc5l+tgqhjDuTjmFJB9Z/XETIfkcicUP
DuDeufZgEL1EhhfevAl9QxFJGBDvaNlJHl6a3mRAVtk6NH0Z9YKsvKHAOMOc0BbwvwzLQowisoiC
QwN2IJGpDS8exzLTrThBHAO+3Xatd2WBHl7+F7DUZcTgPd543PBAqEngm77lMrDbmEk2+S5g7aH/
LFW913OJkLRGaAkfTz/GsEHxk7eTJpEZttTirUbcm/arZiQ8E1uM+O678M8V4OHqHdKwK2HUNrSt
dIwaVv1npBCh1oo8CsQ/8l1Mh9B6mNPRvAPb0wA070S5KXIXisFPETVc6vz6f9crD+MgaL8l8wUm
xYv6Nm1NbcuEHaK3DnHl/ruAVhxW6b09IQSwWV5s433m5ZPiXlSm3jjOYSHz+AfVM66XM4vh8PY/
0VGOO6qVg4q5e2N4E52d7sFaVbo3Wtd4VmMNmyn9vwQydQztXy9ve9fI+34ChXpZrrUd6QzEJdKk
z9xSHwCCbZwmD1krQ69ihHEG4WoA0J5CSf4/w872/9JZoZHjwUg0kgaBkPuB0IYrzfkBICWEm/m3
mQgUPvwrdN4pGGMntKqGBlu9XL3VgS9VDxnmG95EaKYc9iXZHpZcBSu7KS4b0edy/1bJlVMi8fFW
jphp20ijqJMfyin39jp5q1a9zHfgMwTe2rcmqWsUv43moqJZ4lSxasGu5iCArU9UlP3GoBdkUnv8
z8A3nDCSVCHlGuD8yZZ60Jzly4cMMCxGDhdRXgrNuwhwIbRnqQGnZAtFI1MrP+9UBALr0Py4R/IC
ZOanodXoHmcf54AwjQLmk6mt6GRcBmPZy7lniguukqMRTwnhtPWgbxbjkWyr3WNtjzcAVzuYwN88
0NzpglFi9xgj3s69d9kpNtpCWvpeUp7+5vhMKX/vFpUuXnZUoVuVKCnkZ08dVZQ4tgJxZJkAdz1x
t4mpOYehsRg/ylN3dUEnseF2iisT9R07Rjz3gOTtHbT4F7060OISwTVE7X7DyE110DF+ITOzsNOX
RshwSm9gPZGIWQY7sCdahXq/ZchwZEwBK2ZJRsFzSWbsVuPK/g8QGHRWPGHOjVT6DShbFHcce8Wh
yWZByY1mktNk+EM0WRIkbGW08OzGl+YAd4uw/Kjv/JbZfFu6UrcJrUS1O1Ek6fBoQtZcz/y+Rcnd
iKyEFDm8p8HyHkanFbvAY31yD6qk2ASDG/p8gVd/WZBn+ZlIaDG+JWmxj5l16k51mGb6RSUkqx6n
cisr5fRJxFLJwbS5FOZ7jfyYqAQHTsqSO95G4oMqpDNMBIFIYYgInMRBUb9ne7UUoUmSibTbWzXh
dsI5qfMJ6tnnV89Q3+ZM5p8AO2kWuRRJA+GCY4bJ/IdQP1vdU4A4KmFuGo0qaUGivQv5y9c821/g
doNySnlDgUXweXGu7+gf5e0A8vZm/WecVbbtYTNLMoa7YcNcFzJwAdJzJQQ1WjEE7ZyEUeG0OOaE
e21rlgiwIdXRwhZ5m0KYo37oFe8Br4pg5HeZUTMKgPNS169E1rwrQLQdxDi9NW9Pv7VX4Qb08Xks
zEht2DcjdxBoQq3k7Tg3EbshaXQAO71s3cMGFWYB5fzvWWESo1IlbeP3WsWonZkBXQUhYHvvghmn
b4VPntEzBLBLrQPLSE3Ik3QtruxQm/hP6ztHouB4azXazO+Yp5S4jhYQC/OohA7bcPUZxK6NMX97
yRg3dIexc8rOCGmJecORQ5ZGGitVFW9WB0/nQ17LOS7LHfzV5ot8xjSUXJNXrsKZBS2oqppqWqFn
0jKimx/2OPDHCSEWSeJgqdNbCl+Grvfb1ACNRplaRV8S8ltFQO44x1CDn0GpzloMaQ1wMSNLAvss
wiPQmK5Q8lGjcVWY0e/WGaAQDy6xa73d94kdKcgSeCpYCSZ5+1Gq2ux/0KBC6oEsmZ1PgNcJwr+M
8koiVHIQ3XFDFwPcm10cGVESY8ZcUEixD/aiLI74k0eCMByoh6Ep47Dg4rUQQgwp6nKIPh48Wmfr
biTSxdnpwDSq419SGgj0LHCBv6wk47Ws4amqAmvHDcBUyx1DJoDhKFX/hhJLvaEyyzIwVt5+PdKh
PSxSEE4NRNItRYWriHw+gbkLn5aduSP7Pmm0l51ONpFFWyuFzqBpWDyU+gEXcgZkdU4idq3D4i3n
MmKZijrjYidbmFrGy1F+jtHLotw5Kk7BzBwMZrx8HH9SanO7kyYqx9U5GJd2JMJJ/pWgkNwf+geA
cgqJpX2V2AUpyQEEC9mL9PChdYrMEUeDBWfcuOou4dwLnh4dJ3bMybG+x0rD0BS37DslggAQiGzq
bAN1QvtGPT6wiJGBAe/DYhAdgbABzYbj78XzP4Be7nFgPAmNJZF+sVfANq++sFb4N6p8ePUvI+tA
LbbLYZcditMWTzr9dvl+ECuo+Jc+qTNomh7fhuX336s376M8LR+UNyJGQr/2BaM1IOk1T0O22Mu0
bgMJgIr4fAoRy+vljce4u8rn1+lL8Qrsgbq1qCvQ7KOwI/WOMKjUqPqyrspMN9MGyupicbfJ0C+d
3nxeNvEY2PhbmGrljtX73jGEolCShO8aAwGuhZlWWTj9uIsM/wM8idyMK5pZrDgndECc7/dWyhgr
kMZfG68FtFonlbxsxt2KL9N8RpGcV3YVBkedtdbMApqLdOdzcE581zvojH/NKE/QMM1DpIbfxnQS
/VvcHwKquAkrhARScR8PUCgbDbWjeNXeMPjuE53ulVD8HaOID3CzK40LBYVDfvutijvHEOErE143
0GGU9OUK9Prdye9YQceJE/+euGfjeGGxF6EGP2ISfo5wQUyablkH/yu2WETKa9Q6FrZO3pCm4Bbo
Lkha3TKczojNNbH6GiuyvAZuFSw74S1MS+0Iv6hpSlidrVfYcvT+8CtG6mUus9bphk0Q0R9NzruR
OYjwizSPru7eWxBLfAauBAsa6arRICJtPTcu8mXub0gTZvx7hxpap903ITtyuUQrUxvMNNzuIQ5c
9JOg2fG1E3OKJa7awvQ5TUEBF1d00FMynShtFOWaTJryqbUR+/LCWAyePaVShqBPwf9BErYcq/5I
cmg55bss9VjQOLJe+KEIhertZsKcJtL7w+sMfNo/zsnWKOvG23Luz2Fg61fkht03Kmt/6Sa1FMbw
c+qKjt8b6zEjwxhjKCsPgMdir+k6wEko5sNmbNXHLh9ZlZPIVgr14w9O4C9ArOxOhPjjpyZ9VxeH
+Dq6ysqoKjo/jnHmqwrUoYkGw6Yhmr9EECsX/8g1VubROc0Y5GTOM635yIRYepPUb2LDhYMmsaOo
Cx5JMy/Tu0V4FIvFKNsm0/8LbgbcNqdy3aCOOq50iXyG2NF5CVYxRWZXX6Qkli1h/WosvQqlqx3X
MgTJDXiaB4zB2Lp0nwGzAk8AMZTHuV9uGghnjrrZIPwdcHzKRJfHcVogwzfScIZiRxOuSlO6BKV/
nR5yHjgYaprq4mCZnQw/YAXOfaxT7fYrLwA/6bF4tImiaqSDR6G8RGBfl9Ep0GHgeRIXowAZouBI
K+FS9Il+WtO6kN4M9NnlfNk6yLA6pQ0P0XQ5JgbzbJDrXLtrH9VNZ3cB4qKb+FPhIx1g/H5ki74Q
ryRdRf7QP7y3iak183XByieAzrY2BjkGeJ4BMl3BRbVEVkG8DbNhfcVH6sPYTSk93Ojm+NYVj4nh
7SI1xypyxfFpUZugKQlUO4MNX0kztzFYFWXHPp9P6fnkxlptgxNOktEUatQFuHVUgwoDEacJOV2a
DBNPmNUkO2rieIA5IJxuy/KXwPVWsjXzSUbCdToQaOG3O0fv4QhvUzi1pNI+o9IHew/WNXPM0vKv
fFz94wJRySOSZ6ESJ83itkVpVnqMOopQMslhIn7Q7Awz43En0KThi3AxD7mnIKHC5VF5uamls0QB
0wIuqXnTA8Ef49Ja+F72wGa0jRWZ7qDDcWZ9EstSGnJDjeXAROHXeWs0d+pgHQpVpUTRwK+BN+Pr
cg5GP6OG1WDr2M2oOQ1p/OIaeAUOeGFUiWooThP5aFzcv1cWA+37n+vtG0tnbPRRIHRgrLQWnBqd
9WUVrALLhkcAsA05ZIGg5FmevnnkwGmGnCb34Fj3pMPsPe5Rjf0NpZW+/tnIsbCw5ATQavfubnpW
9bPWjw6kA1cQKuFsJcCK5f6wpFNyMG8vsOsrKcge/sq4dUEkJlAZ7Wf1t+P+9jxa1mb+/pHMmCBO
VOJENh94DrcjSgHkP6fsNK4QCYL3CYAhFIHKVU7yEeirEWX9q9blccTa7EwZ4cgLtTHiTaYbcGj7
9Jqhvdem31/QwK9ZaE7uTmt1WUH+kkG0HwABdnydm05SduPYeapKHxPUxbtwwSajg7SomxtK6XsH
iHj4HICHIgWLVkQFlVXpOyjMH1KGIHIwJWPepGitOyf8JO3lbvsatQ5h1UKjTLl3Y6RbfuDTH1xC
Oi8ejzpShruummjjxvZgQCoO6wGLonVhrdQ/elK3jTXmYEJCTf7hx/gcRjdNNKGvbD+eed2TcrK/
2nJrkLPf6Y6G1ocVAr4LonE35u2ZfGWovLYkg36c0kiXXIZQcHA/ls31psFJgFGFCJ0EoHyfg2qd
zTF3zEbuj7ogsQgEZU+W0/ga2G1wVz1PTZrSuTA4RMuBkgGdnMDAmu7Z6Ms+c63W2tnkoSxtgscB
OfhDFi+A7paKPtuLwN19l68VrrpxGwPU7wrV1CqrUejW9JxjB1LhxrXVEsTbuxTP6aQyYJfhEBAq
phpULSM+6HRBsx9eycpR0uQjnm09hWzpEkMwBLOWX/VLk0MKg1egu7riff7uKi9mKoTzZTBM0F6M
eRsTMOBeeUUbyzWEiJ06aq073iC79x+6FMxeiAx+ZrPxrjitXrHdDknhcBKkBU0UVd4sirQVbrrP
aIbiFy0HMJQHMzxRL1VxxuL3nVMZrGSI/kPqzolO37NN8ZPbZyT4AefP1/f0m5hiQHNEWQ3p2HMX
nk6luZSictOCAaP1ivcUwhGOryojKVECEQCto6V7FT/hl85H9trj8XxRmqb7cKlKfTGfhoRERqTv
ULs2hYCgchrLGo9sYf4jbca+ieyq/X4mwBDXUOKuudgqrnn3SCaRlTh02sgnUcRaCWMQKhdaJPNl
qNS5+0vI02vEtDhhyTxCJr1xMZjRuMce0yJ5DBS8jeJTZuBJrMiBIoSKeV6srb4sQpptqnmq0fEj
1sT0Ga7AsbEQGztCfhovxp8xGRKn4/EqjShQ3oQsa0Z+EJTuAGeiLykRIu4UMq6/0RiQ0hJczMLX
bUIOpU/bgBk9WqwEPI7nNUuCjtxmG8ITFVtB8ZYN4mvgyR6iv0AvFzHVr9QqgZxdCvM3FzK89BOX
Q3k5BtgXFDdpGF13YIZVNsypYfF5BFDgUapbh+Th3JYZZePEK2Xs4T8ETFvRI/wnC5khvAl9gCzb
aLHwP1/6oLGCMnfa9+wY6N024Emk9oW0dUeQlkSIIgu6OVlUG5f882W72wJmPEznhbsxzYmiykW9
8vDHv7q+s5CVehPbbH/y8+rCnhBvOFdqKHu1UOQ09OK8/+LypB2JxoskZ6rO3EFCCOZ+WXeVbOgq
Xc/DRyDkafMsBjUGfIYklzlmBC5pSZBf/e5e3fMphNl1a8BBfvvAAG725XqFshHiFOrLtnwkjoEj
+DliG0ZQYHhWIne7El71HKRAMPpbARzAE/rlz/g6VHD2yEXCSMMwYlpuwkmlyp2e7eZh698fI2D8
owgwdC1Q1P1kOP7lOO/Yf2vamMaHZ22X9eK900sk7LKXlgLaqoFq0+2cRbe5j1wbCJWR+F7IEeaJ
zDuVwoDCQskg5gE3akkb2fzoBmT5b/Yqp/fZNuzXgJ+tgV8D8tCscxtRJqqXirJ3v1f3xdg2X1QX
+OTFMF7+ueM9WHOwBqEyM/l4Ajii9xEhm7v1ey3J02E0TxwtGruxRmyBOPU7NjM1hiHmUNw42j1c
i/hbzf76rv4ZYsfKOpNtVUV0B1gHgunmutVaxgJvOhpSKDOi2rVoXyeFp18dOL1PJVXYshdh/D51
kzpBBXAKKQKpR5exFzTNH2wyPKEwkz27/Y62fwXXFroYyXvkIRxq81xZlcrZY4YbYifxR8/ZAhfg
qZ26LYflH6tpQNdc1XuVW8/bseP+u5iHTtisoh0kFjtAsNSgHM3rvYaKDjdwCzpqY3s39I1D0ni+
CuOLvAMcth+vn84wNzrjCyL3WjFM8OOxt5sOWXFZgKGA3dTcuVEjvv3xKrp6T5mrAvLFzkUMMiGp
7yZYtrs5JZGJZ6LAXz0zYuCbzkMwZMkxMH6jN2MUY5UAQpp1tat2hmO1WuqGaI1miKiefcLP25hy
OUd4lqFf7Vff+I6lk0CEftVKAYLkBFjmBylCfj5OvF/NzzSIpj3OTI2wCWUdS++27/vHnvuA0y6g
gZhodnNRBhOoPaUl6gULwdKCWbWhvzPOv9VEvbcYVlz7vrGcCvd1MwU8s5xf31vFoo4hz3RlJ6fp
BGnE10jjp6ZYU9YZProyEeZSxkK6Tpnx/AEsqKnTcGFjdX3tjxCM4efYFKPGxGc+8Fja4phSDtz3
bAtrSlCOSrW8u1gE83ovU+rGsW3APSmifKIQrFUOslgKXYV8CrmItcblxO4txezAtPtR4MdUFSbJ
PTuY3Fqz2q9LhxARjM2YcA3+MR9CSLrSo9eZBExZG1SoOV/1bzp9EwrtoxboNt4mhhl13ucioOHo
U9JK6Tg3No1DNDXsyWmU3KKlw/+Ttg0nBjTHrjgExftwNFNARsc/6d6ImqJQahGw1dPOR3GhWN3u
+BBAIWFw4h1pOhoRwHyNOfdZ4FAc3ImY95u6BF4aJI7JDxg4EzbrEX7E7f6YKcLLSKgxwYZrs1WC
geEPwmvy17JWSRxsElW5FG06Y3nS12FK3Qebtsw0HU0QIquPBQdTTBBol77xSYg7FhtxGEqGcDuj
9AwUNYbyKq7GHGhVSr8kvhkoNODMahatJ/jTea2mLQsCBEvKqCLHDKpm/miyVD0cSKpeYWFtLIVh
/4BTyNr8wX2k7FXPbWr9/sbThykJZ0hhCUlleIdmcgGQP8IUk14AWcdZeUyhXKwu9t/b9N6u7I1U
PtLz0j8yO/tUUSjFmUrvgz95mvFgeIgs7UZWRjPdpHcPRQrByhUJ7Uq2ZcX9+UM8kIAPyD5EWVY7
EhVBUXDl3CH9G4v2ilmUpF4v+m2lditFNLhmXeJv7CUo4rY157lesX8jpijmmWQQNuhjesLlhIhg
HCauEBKhGPEB/BLeMzREgYazZ4k5BZtORiZULGgVXn7parPSfTDXof12GqJMJljRetR63QCsQFn0
oxxFAfCzca23JumS/EG7iR4PthX4nc8GqLl2kpVdoS4VsBOC5wrhng6LMv7399Haah6tfPMBZ5qn
nZ5JMC0+QKacB5cvixihuMyVVdE9oeLWwT2r1/bLE+U5+jG1969nh3tF/VW2/ikdkvg10Qz5DhAw
7GshpKCp4Fv1m8scoFBfSK1oiDVy/9pWfizkKMm4ggKGoq1zGYT+21RkJzUlYRejCvyi2VGIkwdg
Vc/hP6RFr3FVPpSp9zJMYSsxhlZcd8PuEUE35EyXtSKo4tU8GNffsNTgJWVNQVpv2IioXKDJhZBu
KqCkZZgvR7MDkY6DN2nKly9h6ciyI6qmBiGCfO8X9QNd3jqKV/brfFlXJPKqLZv/eMXHx9eHzMNV
NsEPfW8kwOK5V+OH79hPmqPzZcJxdhybBXvpvxSL37grlg2qsEdIB1tVtk3W5HEHrPxqTgdoT6cB
r+i6WxORUGQatQJQaZRm1nSiJUZJ92qbb+mfEOcThFdk0AElo+VXphXrTip8JOlwJSJBNXbXPo9N
m/J0+F+tvSD4tr7q4FdoVXzHE0HhVf5Ij4sgxbX6DZ9tkzq3IKBSo9hEMCBrSjTRvWDxZgPqqIiO
1qhoTKCxn+EafsN53Kd9VrVHwbpUOfiJDQEjt3BCPx1q0qmedcNs3XKg8AzONwFnEJwVKIF4tnMH
0S2Wi67AAGJMlGK9pEi9Pq8/DHCkJC0xeNnFI+wBpJFxoE6l/AssR3292PxB26TiRb880OqY3wgz
DovEH/NpRSp+CenbTC5vVuas2s9BxFlVyhp1hQ8VWDsy0tVCR0t47u7ceeCXQFcP7oJo4WaBtePd
5J6wdD/IQjo+zijbWLL56weW9z8fgJwf+//gIpuTymIZvZ62TT4t4pF9BaSz4gdhziiriNQOz/zN
/2Xme02wliGU7PH18ognK1ArlbUISTEdC3ZgRR882URQ/QZmQkLmZro0WmqFCzmWaGwxC0hP0Xho
DSpeXcV5FXoX07555MZVhNBa5e+qlwRW2u6K93x+DlvRmG7EbCub/XxgNjEQADhhuHoWzc8+Ml7f
e7fjAPmUnj6KNYBRIegbd1ZVI0HnPHxAriekbvYcDpivQDzKLmLeR1KowC6FVkTeRCIQ69BfbopS
0tKlALwzTjLr4jZsfJ8GKxWtq6IPzh//aptBTuaIgHkgRK1no4CFy2VtzWpgHIMkDUZ6Tu4Dp9ih
/00sR7dYXdOOs8Jx5vtwzYmLmygdu5Oz46MNQIzCw7SP+hs6ZuhJw2aTlCpyj3hDiW6pi7uGSzuU
WuTm/UIv9ACHIPJ8pT+BX9rhLMlIYUyqcIm8uY1ymqjyEPPFnTths1nz5/Z0z22ndzPko+L2XLPe
wtCumdK7Fwy22oCv3AQONuEOwdykK43Tgwh8MSQEIngxU+B1J30X/TZXv/a3rRXUvg07juG0v8Qg
RrUKFsL9Z60o/LMNNv8YugtmtofhV/Q+LJSB4H9XNOnWGyqkVJefL3L7sYkEK4w4ZDu2AeWXBacN
a6n/ZAKewwlHI8wWeY/+HjaFn6BR6P8W3ezzaq+/2iuWa/j6nWJFCEZpKslbjJJT2z5HZ7oYv7aa
E6ITwMNViByrs2eL/u19xiHYbZxF8di2Z18J/nCyTyqmlpKfLWeey9MJD2nFVLVn1Ow4YYyYNfEg
TRsX/vLs9zL7lOUvajbAmSisGdfdQ27wvpF7De0bBrzddyNIeaw1a5MF7AVp/Z33kMFxNnHV1OnU
cO4l/cVhuMMeQuYNnLS59uiKu/M1R7YHoVFcPxB47UUhJN4OvXB7fx2NoJf//++fJSt4LyixSHDS
eqk6mnxxrkMEnnZMCQC39dNNE5bXUjQIekz3VA3PhlVuZRRF0mU0ReolfKXsMdWXsARcp91XmKiE
3458B7qfRFkLOigOympIeF63Kl2B/TBRoutwQwTodHXcaFo0funF/KROF/zBxQ+2e5dFOTUetI1v
YDoiVU8vxsof2cV1l4vsMlbP39mdyWrfUtszdI3vsXotHEO8Bi34qpRL5hh0MVLsJjIIgCwZ/v3A
hcdmaHThJeR5iufZxSQiothQ2O9TdIDn128XEx0FDeHMw2JNGWZQ/wxJeszwC20+97ybd2mkEZN0
1ScJTOnTW+W9P6orGCPOgsiEwtFr4X4KrSW9fMdHh1ab6xOp/2XKBGAh/UclTz64oe2bkLIYh+S2
9MJBW6XAOhpVEahO4s+grAMGqtFsrm5jS3NiyFSH7YTlebUEjD94jdmEslDXENY4TBEmHgDiVcoU
2lsU0xV/3LIbdXV5N6uAglVg+enbF1Wlcg7kxMjw1z2nLtWIwaQE4lwytUNWkR8NkxweNOYFmj5N
+GeEHnBwB8jX62cQhgn60P4VnXhVnj/WS7T7yo/ZXX21zY/OYluCqonRCxGZcyFGmwJlrlKSCtR/
JQIVBKXl51ln2xJYWELrlhtqqYhJwqt4vUq3cglHsX9v9yAXsztS0o+RS8EbYGDPUcpNtNtFS3EP
oZBW4HG2eKdc8RQL+bg1TSuNHOAMqeB2MfK+3jjBJssoxtWnPS0i9Wa6P3nSe3aJwE/Io6oT8H/u
jhxna+7YT2YWxb3BNVq3erFofoO5HP5vMhixg+3ijESeC2RFfcpr7csTTkRwMSBP8fEUj4K1NRfn
Lu9W4SkoBEs+zkwlW3XFrmhpI5kAqtbRxRg+tqcdYau03gEqheUxBpqOz4a+wo30dQu6hzapIU4L
sDj2+v6589LTRw5MHj7qwfu5OXJWTbLQGQqrHNLpGtwIlKkT+W1KDnFVx8dIu4LCIkwAnvRL8FIf
nUMl8I3QJ40efa40XTEhwW8Avx+QrrDY2C3TmgFYFcQZ1+GUrMKUn9Rv/g9MagCOxq/HfqyjnBCI
3dY5l1R0mFsHb2b68vNXEPv02ZmruiyJOjpXwP2w8rmdmNcbC9ZJAgvmN7FxCGZ4l13y3Gg53TGJ
RNIvC6X5XJPhsVtZz4qEBcJa4nISbpT2z8ReC6CN+spy/QxXclnlyJvdfb0Rf4O97VVidvqA4tPX
WmKCkMFUIjCKxD6AEz6B9twsu0jDoq4rB7agy9VQmvIygsdsg++jS+6aqEshXVXx335WsZG0K8Sx
ycScSna902lril0YKO4mfXHkBoQu4S1S2wm9frej9qJ9xNi+Dl6gpyS4amWDNo3dfXDXAKJuCQHZ
GfcuxT56PJzoGUs+chLYAd7+RgrABkdvIWLnNEM/1JpA6m8eyIsCr902/A0rNQXM3yWmIWMnKxuL
cJ++jpJJDkATK/KoNer7UXsu3kQUSpa3lrgkg7YGgzLne8nbui7H1IftRAXPiig9urHNpSGqcUom
Bdzt/prWYvbZ6sMr1y5CHnfpnvAxxLiMVCMck95zqgBGxUiZecsV83zk8ePC29gcEfXE/CiZlmVU
cwXeH6wA7p9KQ2YB0qO99/V8ck5MjfoFH4g9P0mzT8LXqpshfV0Jx4+iof4gMjKcWWEm7V9i3tDN
3fqpaX7MK9RDiwx7ZQ5CbkPiDVNTaziQOUgdyJ7/2UpcQwwt+p9vvUqen9F8Pa35jGI4FKJXsfto
S65wrJjvkKOz8PWBOZWtqkslOijHC6SUTYCtaKEH/pCiotMu/0mRJthckLMEufJci2Jjr2Ho/CMz
mePcdtqo1zyteOF/0o9bDqg/mFMhMPom9OwO/lBStj3ae1eXxOz3rhPsVb29S24o0J5fOh+iZrsP
alD8yK9GQ7fQ5KZLJLKUEAREaG7p6BLucBknJ8RemIhkH1uYq6aOb/9l5We6vto06F5iEJhnx3Qj
4FT5DBEnwIlsOJvbNbS1Bb6by30AgrLEoPgI9LQPvCqNJOZbVKhN1GXnFl0C+LZTRopjpU/njYr3
Gm0r/70FUxmmQLE8zBnhHQwXG5DUBJfw63ofC+3nQkNPuxI83Tudia/pT/VhsqF7YNqjAMHcpCk9
DY3EcEUQ1k9Ux0RwT+TVGQnsTNVZZuniqoB+wYzF049fhiaBatAo+gmpts6tQH6+QKfZyZvor59m
3JZA7HCUMT8VfKxATiiq0stgSsrBgpMigQGhj8wO30bEmmhuXWf1womezghyvil083aIl4PyUMqH
OJfnKLD2ElzDel8GpgZNf/nL/FbLAIGt/teYwKjwBRJ3zWfhxe0CGkQO4WZ6AL/WnN2F9LBp4fOo
XLsJBZij4f7imesCe0V8hscz4SI3Ie2AiU1uz7TssuM2ctQbEMgGizUJtlLI/YigqWUTQZHdoRWu
kEgyuhVhN1YAIvneFPgSzTDlCG7VROExOSI1uQzzpiCv1EtEfwhlmNJHIZuxTn7DjoD3hbUReevn
NsjmZfXNd/aQQl/IXFuRCehoSG8nqg71egvBgZI3IHDu3pZL41ZrRKT72Gc/dUlvPG5IcuvWHD5N
OdqYLUv5ChQsYEfjMWbYzG1omcZ2+dueIQt7PduzAmJ1NAYe72Z5LRNj4I1BViwGMHCd838jl0cj
TUkoJIk4cEqVHkb0tpoZrpSRH1D/DnzBcqCLmal/NykoeneENCTN1tsP/Amd0gPHYoMluN+dkVr9
FYA7mJys8eCLB5jzFSzx/fHosgll3A36CmztmUmbgVwta3tjHn85Rvt9dGZwHgU43rUu60EViE3m
W1GUinTyIj6t/u9tr+la6XwUFiRV6PlCHFHNbmI/URxr/JmHUkrD2UMJIaFYfFx7s35Or9EEFBrv
SEoBEvLaSMoS3sTL45OVIPjIMhP6ac7ThP6ep2oWFg0I0fxB8Uxms7s58GUz/NlsPuDqsLcbbB5d
MjyMUZ5dj0BcQdA+KIRdclKDfuIFxNXnjNlDhN3Xk1mvZ8ZPXQQf4os7GGTq2vDzrdyEABSdt113
4mTLyKum5/GJpDNxNlsSGG5luOBlR5HnrE1oX7eGFsdmP3qTp9sOtmplHF80oYKKmq/EwDrDHE9B
QPijfeBRpZ9NhQHabVFoyq4wBVtfkORYeyAXQm+gxy/tjP68WVZZalKbUrl8E8UOb9wtIY06ddwf
BTAYHrqxUnFcWYQQN9pBeBimgjspzRkRUbrqQ8hRaTueRRpB5MpiaXnyXZ8xLdBfr2+DXJcDO7Fr
rlpUYnNZChaVQO9aiZB4YfzXmejogvZBj9VHH1I9+ixA0BFTt805gAEnvx5Ee8+lph59OWQWIYIM
alGKH++gNGwGDaUXf9pTTTFxbdauzvO8ScQ+R6tF0sfzgZoT59uqz8J63jucqObSIPCEXloAvwbA
vudj2RZAhlzpapwIJ6nCR6jRbG+Cd8wZiejdDK9M9trHDep8k0SOIXhJl0Rsx/lyWEWgfyMXUJkV
Mjxrqf//QS2brhcYtfFFBfLrjzPg7m3TQVpiqhnw8u+Y2O5175exznBk2QTwBmPWizWmh0+w5jdD
CeVKrVzgqbI+b817iyYTYDkXkOOdIJh+xUKwW4m9U0mbKqLBYZ3xAIkx2UBsjKjNeHAS23xccdRF
27Lhb5MV1PqMPwlW34Tm51TRoFyoCTkNerG5ybqmaFw/td3h2mehMgiy6IKvthxmu7biB1dFhVGW
+kJ1urx8Z+ZKnsykrdnB1HOYzH9zymfZxCMhlJDJCJmXjWBvqlSCEuS9tFI3HPfNccfC9wv1E9T3
44y7Q9EHdzySXtvcPkFc8yslW0i7F+8tAjL6DwqMQRaZIUyNXyQFCnO4ZVngXZbVft3O5jpx7rtx
fllnXNG9jMUWddBy4u5f68VTd6Q61ILMHEKw65R05W5CQuuVk+7tbpaMsrngLT8giOibgW4cYahX
coCavLirnFRuMoG5ZOqE8gchG/BcFw7NrnY93wsuo8SZvkWU4MWHUTJAQNNKa03NeCL9ZhVbgtP6
Mr+rNBq/Jlr+DUzqQIalBd1bZ+WKNCHwtReXmUKr5S/R40EwdlGQeAXBP14joTGWav1U9IlWOu1A
GrBXfFmmXExoovjBjSDsrAIXuj5z8UP4D8JLg1sV9S5F63CG9vpJZirw4MfJsTcvllOCDZdGy1yE
XWJuVxrOTW3pdWFwGkYh6KvL38TKuI/aUIMW2k6E5QWdJxYNvLIrlV1EGtL6QTHOIh7Y+AlGaD8x
xJHReO+SMF5KBQXhEIJ3cQ4g961VMLujbAmJJ+3SjtgEy3MQrAfoQdA/wrwXlBGOpXnURW4pFz9o
bqdG/9xdt9gnAm9J5vD3OND9GxAtGB6SJt/SUDGjmaiQ1ZPN3aMvffYauZ32Ucl9TyJKwT6Z0hKY
hHYKRU5lOPbZLl+PJuk3AXW8tmlt9g6JizObvYXXVeZcd3ougQPKwTCFcL0AayrFEUDu0ndoPeSG
kB8MoJGfFbMAZlp3120a6yKQFg/4KLEUfy1jDttirUwPSndrNk219c8QqlF+1lqeUg5LGJGcMA9Y
qzsWTKPECxij7d4MHgP5KzxkESlefMMgP5zymECylcyt48UROzHqfIZoolYrVYWl5WyvSMWLFpfm
2abEcl79g7+khN2HomxuvQFZFfzsUepyNNPdUyoHQsDx1q1q3WI93In2Yl9BhqUAqlDypcirSH8m
M3wNgTS9DNigFSq3SiIr2/2usNckDoGuSMu7JqwHwI8OrsE/WtL3rXCSuQ+/2GQawUsMSiQdrit+
HN57f66qEAoQjePN1EjxqeJHA96ptG38hnQE8Jrpn9IVE0pIsFmMs/go0mYbkVrJwO0V8zDVT+Gc
g0S6g4w2JulRBd23KGg5a1w2T6Ah3mvPRaCzmlpIIUPCj9bego0mwIMpJ9FacSM+ENcvji6pWi/R
jFNMaZnhQNRVxzubhpzhTmDiMUb3XaiqtzjiSwSm/RUy2id8PRW3xH/mNYETkWitzayrmb5C/4dr
5XllUfH4zj3v2RVnouMmJ2jA1Bf1R0ZMO1GAColGaLP1GEfbGVqLtpwR1vHDQxSjIaUi/lqa4fc3
iIrZqmb0X1tv8O9+qYN95O6e3tlcZC9SyzWB3cViwr4V7rmnAZsnRB3Qxvf6+HSd1bIgCYmXgBfc
cBSrrtrIkNbaF/JqZbeiUpmWADwsCdoD0gcexLkJoG45hhG2W1T+zr7xAmTHA5+GXKq27zIbjTlu
32E8Wq4qSGurhc8VNNXmUs6pBK3SvtB2GgsQIOntd8/NOCK9i6h1+yXdS82YhejjI/yfHheMGL9/
+RCpckpuaz8TeyNz598CAoglC6VqPUcWvY+gGkPN1LjCYJcZ3dnx/dSrNZVVe3vFR1r5X35kH6T5
HUJqIJttjGEctMVWiiTiZlTbPyNkz5IKfJefPikItnJHvhqrYoy1cXCO7d0lqMRw3iuSrWrClkLw
6RuWQjn4UlBICeVPL8mxntA+c1T1pg2jp1OxN7X+LwuCJ4btKPuk/pm/gbCWVLu6gHgsi0kuTwhk
sPHjCJ0oA1zTPy5DTtfMQ85XEPwbjupv265V/wOdfpQIpSn9rwoEdc6eMAmBeA0nK2XFt6gQd7N1
eaICdPvGJXZdrn2BtvwutO/gUf6IP/7i7fxonJneckJntXWhaEjbpIT5agh7DYAKGH/LGFn7GtB0
MmhchxtROdgjWPvA1Bem53u9dasuu56U+LlMPZL9vlRnXFM0G4G5NWTqgcB6vUrWAp7/6AcRUxKa
Dw06uEsT50YXYXrzuPJ2WbYqwrKKrop/xmOc2lh5XL85PDte4uvqAp2Yfde4/WsOs8JLzNqc44QH
13adLCTg3wTQCYgrT45v/6/XlFfC//NXc7fGBDCu3Q+LonnVPcYzAeWKt87FeB4UsWRozqDVdM0m
fjfeHakrYOzDkUWVSAau+YGSjtvd8iOgl9rpwca4rkRABhE/yXxuG0tkojY6x6UOqy7U9MkTtdyn
lrzcL0bxW8jUxB15H5teI/LJqCUuDClD55G/wnrGVxHUhZeD8jA9z3TT1ZK+1DBo+KuVCyW5K6CV
yoAl0in3TyntZ8omRc+MfNIkSV421i+P2oHgRR+tZTxhoKGNEUHrQVK2Zz7FyLnaPOgMAeen0C2N
/iGdQ6fo4m/P1bMGJESGujHGVDgYUF4k4uTP/zccvVKi/Vcw4ybxPWlKiWhmuhD2ztBq7hk7Sykx
qIQQ9yMiNJ0eRv0SwDalTN/fiwWKWnh5pM8JkBuJm04dndvWwbQJv3Pd68P2gt2nYcYM4pp/2nNb
GQzvvmVimTs2ViWBLPcVnhzi9427ZG9D01SGcfu6PRVgZvV1kVHyfP1GvgywdJkEHrCWslVU2qC5
4qUgIkRj+16bdOdmhF9M1WwthZdn5UCAonr7txexBorjJOApXJCHQq6OuECPAd/MrSEyAyGD7+P4
8gJ1HsgQHIo/9MVnPeQBADXQCT23f555c7hOP0gAtzwo5TyTk0JEjy97JlSAUYiqDS5RM3Cr59Bt
/QMVq/r5CDFu7CcrJq5AIb81UYcLGxIKdUXUz9DDh+1gkQi4FLxmswY4QcCPWlVIUI8z/b0tgY6c
xpnQktyb8TJctD/n7BR89OFPJz8P33FPxUM5mjnq6IpU6TBGWj6I0zkura8rVepgmpaOdZpnzXZQ
aMz2glATqnpbc4MHu/vYPgl0LCqYlPCDi9T8URSGPhP+1OIUDD4hYKTjftTSjJW9/gBk8zXTNrHV
86W6xSqaRLi/oTDbsXxXil1ToLefnBcV6pCNv39AoTwI/JyCoTbmxGBLNKIUFBqBW/UgbM8qVNf7
RXD84UZobAxAaUfbBKQPcKJYKAhZWVNCqxajxsUuHojuUa0p8N2ivFQueW7YCgpTRZFSuRjFY/1c
aiei4WxLEtTLhYlExg6xNpMCRhUtIQqk6uXUyVBnPlwy9Hlk9limBq0yzeYnP3Py7DXVN2QLDlRV
OOBPk6Jt4+GxBGc545uZfJcfrBO74x7mnf3x54EMqtWX9rMfUT6TwewDJkqwhMqwg0zRi90WDDjU
EHIrMkKTjfGxT3hTvlqkVj60oT6Hk6LB3l9pGUwiThe3ThzQFgVq+Yxb5UG+taItY3FJkI3S1q9W
xHL9pf/A2vOAwT4bvkMwjwZoo5YiCHUbrRQAV0HNb9zxDixUDGF/IQLfeZnpXPZQsquIOguxcFMN
Q2yfLnej5NjSU4MIOjs0SYa+OXCCBaQZnqk1OCiaopqI/qKftv8RbKA2OO2tlod1xB6tnv1qwEyv
GS6z6nDl4UOee75Uo9CyWOTfN4dp3+BlwCOPuXe5LR9FgfyU/IxE8FdSJxXkJEuFZiHwlk8x2aYR
DduoyCDo42TK5VbbG57oryhMzEqboqa5FNjwZ1Z5+h5G/FUugJEltyTGpXlimIaj11a52eZSlEm1
qkv5QdNcprY24G+4HllBuAgZGupEF/Ks6L+z+ZVHAobU6+aNeVlqjgVxWvEccm9SQ4mdNR4euEh2
U9FxmtQrZUbJWsIy6h8rQm2AfbeoAyXW/4vjGZuLsUw987QoSHBc1Z2ss0npfoyIqsBKb4G/ejjF
f7MSSyJsIeyNBL+giPl1UWureaPBwbpGCVyjA2ZreySVFjl9Xxp+67VVRTKzNl3k5qN0ocy8p+Uc
kJ48ENZRfYrv+Bw5s/DiTmqLczCRZXOSxohtfJ6oGiJYA3P6aD5umEsJh0j5ygrfbf59U4XWRPiz
6MT9nrZQYIxU8ykgct2p9HSUzhrsoVeKDxBevpeCeToGEuSmZEy+vH1anhLcz0d8egi8QadrgFXW
IchG7gEhd9+sGi7eljv+vxo0B0plxO4UQvBhcN+fc/FIyWrZ0T0s5iw0380T7kteEc0GQ9M0ochH
YkgP5G66o+2i6HEd4Zf1UBD7ACtMJaHqP8z9m7Lg27iFQujgonbw+dHEwxaZD795eGia6paA9Wo/
StQnymI4hXVqzZMgpeAFs48R19jbMAS7r9NSIkhl4CHhn3OUlR5jtkGDliH83a4863V3WY+igbwm
jVb7phnBeSUohbTAe5bcLsruxp/NzjgOMCsAKu5MTqo2oHhGcVQBlZW9SXrie+PZq9StllGKfjmw
6/63l7PPuSjPsy66QeqTZW23sSZwiy1nBUXX/Tsm4ABo8qnBZjseEsp4nRDENO8PJE3fTFXA8Hwu
iAUsWxAFO79yEslbDgDKYKM7Z3D7gIIHmJOCRmJq5rGGtdUQelvAO3MFfPY0fwJQC5oAJmPKP/PP
piWVcR+MP7PwqeekZgZ0dYfQdekRVygxfVwjoS9jFdV+Y95c3k3vQywx0WcMZxm0BcfZf3DcdktP
qu6tP81Le4Cq7TVBpdIIkb9nEmVEMLeHdHiosegZh+mM+aPqnHqQg2zGsubRlw735Qgg8uyfejIn
2kg9bCj+u1DfG5CqjfLSe8s8A1hKhE84tWtYoN08iU92bqI8znOGjPMJAb5u8wS2HS3H0uPB31Yg
ZLveWkv2iYkdgMWC1pd7nQMkLjd5qAPqgeuEVFccoZsNwptUPrewPSPJ1CC2Lgj0E1/BqyX1RNQ2
SGPJnPcgmFS5mD/gHMq9OKLAikxKgZJxmdz9TUF1hGerymmk3QUpgIFN0a0GxXPpbcyUkpLHa+Pp
3Y6xc/+zUO5mjOnYHXv1JCPSKUKy8cDZxwCEF/Ph32gqibyuVDmhD5Aqe95oOz0W1sGRG8kXfANa
kCjjifrZ39Cl9tNERaGgPjuKnCHFtchsPZX0xs5Lpxn3GokFu0z7BvbG26iqDLy8sHARzTaLt7ad
qLqKUkoLN184dina5L0b3r4FRDLZNt37qrlgQdRFNSyFtVMp1zm1RKkChtN4gh/ih5claJavSuEK
CooKXFInyD9bxuY03irxvvi+YXkbSyA2F+1Ch1rsaA/XYmZXPqEMctaazbtQXg3MPJ4zvjTEu8Qr
oBj+NrJCBY5HMoad1jWv05Wl/3OT3DFhgF8zBkyaIsdw/WDC6UpP0QWsMnGX6UPFUdGdsF2PeRhd
StQaIQTq3kvg5mQfVrwrxz4y0gSBTeGqClIgAczZzYIAeaDamxXHRJIZ1J1soorR3B5PpIIhBCSR
mCVIbNYT+0m8RaP7yZGQ144dww9+jDPr5XkVY50MHl6qtxI2QxCuzYilAB/Gm+79C9GErfa6dl2d
lyno3VZr//Ko22XHT2COnNSZ8JHgmhivKJ5xx+h7Dn4aSt3Fib2RT7TZDQeN001L1NA3es1NTqfH
72iLtnSUvbiRuiP0wD5/2YjQ4rhJuDRypA4qsdZB8R8YsoZQ1BHoFf+CUtb7t88uWTsUn7oanh+H
o0m6Cjc1ye3HdS1g4ywmApmxBSXDhxAt2KMJ+vAp4MgUBrM9aj8zwFz1aJpFnrCZRLnEum5/61kV
7FYt8nc6Y+AkIg8NXgGxICqvc3q67JWJ42TwmKnBVoYPyZWXobrD0n1rJFPAj1C5JbXDh/lOaG8a
p4LYsLdgNRxxeW1RPMJ22yeZvzILeOUEoUYE1KiqvDe49zaRbgsD3HSb/M61vPoGCTLdVwnUMLHd
Ur0kksIrD/UNZja3wTqchDN1ng1a2ilmdaAd1LKZK/EZKwM0NYXZzQDmxQEJ1yfW0/kq9J5W61dW
m8MnFlPt9ILPRIhS6/+0fqeipTbUm1q8b08WQgXNF3KD+GuWd4EZbxesS8eDXOGAo3CrGx0OGhDH
x9IwTuGe6Uu2B/vAH+KzaQ1f025BVSjzdClqD0vzxfSuZkzYrN97tXm2cRdZ/AfczXqOf8azyoqR
KFHk+nK9ziyufUX4Gck6gfRWlN6QFHs98ZC4leKDhlMwcPbNSGuCXRkvP71rC7igmlVuUeZry/1p
/UY0F0cEvjs2HXtp3znMpZx6XVMkgUW1670YuJPjU+Y4A/c/rA6KD/dQTzdmjfW85vSKedUvqTtH
fWSswFso+gUaCun5Rcj2PzSa2NRe1Y1pi8LO9wKnifncmZAwtWyIaylas6UMc4jto2A0Z9C4phWI
QaUOIA2MqqwHdv1MqJRx/4QlLyduKB7fAoGZETM/r2iLW97elge1GMSpT7RkWw0YDfWjS8D3sXkR
8Kgoqc5Oigw2KrH6b7M966WcW1o0oBOq/o57Hfs67d1RczOjq+/EyIK13omFR6DlkQ2LQsDbttqZ
9VaibZXuTXi9pBNF3J6bkW5bRqDkN4jCvpWva+WoXV+CwzJdxaIsOxIN+UtlQZiqhwvE8jzFj8x4
r1GvuACoszjlMusmrrThJLfXjgAXaVivhKLGvfHWoakncFm5iEn6tJBgjGsnRV7BdAC0lFfUcV6J
WhXJhx9sZuhbb3HETw8/kLNSh6ayOIVCyyJjTJcxg0T3R/8VEwIm6J22Jbv+tZq3ZatEGEppB1jV
TtD5Bb67Z8kozXK+uV4a2Rc4YUO/2wklK8q4glXzvNHa6m+6n3ko1J3B3XBTO92zTXwjPzAD2fqp
SzK4G9VHfdIrJ1/AgJqTsDh5CVb+2Tdi2lUnFu1sd4w7vfeTR7B6vPlFdHYv2NpdafbrVcPpsB7g
fD045hlJHmB3tlJ2Z+soM24WSfH73fObwf+4x50v/mvoYwCinzKOaNHUTwCW4E1fDG+oDcPOMi/w
qWCCbv4vXliemMfsQAo42cMiFVnRpqL93MSrXzd14ipwvBns5u6HtYLmcgjrbZbPbDlfZsQxWhP4
VdqrNkKVQejCAFT8tb3IQqoVSfxAJnMJM7jFe5KQOZFMtj7B7I3Eb1wQ0ps5M8d/gSGi/JDqDAgt
VDgqIrG0WuLFXCC7IHl2mZH4/YaujbmnaLZbL7gOvjMx4Cd46VTrVoWWjd7hZWUJigFktvcV9VCD
C8ZldbVMdZl0jDHyThZJ88l9aObdB3FULkP+EO2t8cH54YPHHLMlzGNlFqxUnMCliQZETsMaRhZN
b+djwRm/5iyM2R56rGB+DST4dO/MPdYQcyhrWRKvLb0eBahuR5mXQojmD6CaGrjWIaoYJw+WBOyn
4/V8iNUesrGEGUMghiqNZ8Bu8IczGnLEp1DrngmvQpUHf+sKqnN/Ac7PjLp8o869x9FCgey2Hyq7
ac/DAMqvS0OafupNjr1YWEsuVSdm2QMmV4BS2Zxp+qEdbbWV6fVP6ZqcmT9mgGk1eJvkvWN3kOYz
BDqdAOMJidkdNknYZM5CCJci8Oo+7hVLsQTKszkIoLWyHWJUG/otO6qmDCxOUOL4ERU3REDCHb66
VeJJDemQeDaFO6esVih5wxZfBC+7NeMIAyF65CPg3gPE/hCW2V0hVNFcLj0EUhKRr7TSLzF/tI+Q
90AILEBrHsPwaaLgKEVWjYGCoaEYCds8CCj0Gs9+Jb3oT9keD+gK3wGay0RnQlmbUaW7ZwZnf7Oc
Vsl9NZ1W81hIftr/5y4hzb2njs591CsYrqeMr4Wm4dRrnT3KPRHCAJMVg2kqjKrqa4H5oeBhuw73
PoqqkYJGYJ3npEIhftr9XIsyrURiDd1gJsF3q1T3JThGLFQUy/yVYDg39HK5nKYZVBAHV0UHZmaU
RP/KIlHycmYK1XVW48ZFds5TswOiUBGN683JpovArF3PWc0ghGewdwmVuQHP5kBuOTVZGUCxDGXY
2Rr95EU/aIxh9vte7v5k6XE9NUT4ApqLMs3WGrXj0/ZrOyzSVbhlq5gwKAeDaJ+s1iA5D4UcY34s
ZOjYKVvL34hfHatcuYY4Bfs5jh/+/wDMuZbSYH66uzHU4hiFYihT/rshyF1flUWzhnZxbVC2R95x
28ukMjXTFlG/YEnx3iDlTVeonpkAXprR48hi5eVXfO3uRGdfQB4suTC+bw/QZJsX1uh3Xr5ymEjm
wVoc0xYo69SRtL4k3WwRwDmWOwQ56TQxhmTZsoSL8TcOSktqNlggpakXXic0HAQikNy2yQ0Cu2Wj
xxH9izfUVs1jwKwzCaY5dnnYvOLb5ePzc0pbgc1vSi4jdIlAJ4eDFl8VzCNFrQNzRJ4MilvmNL02
az9MIz8xlk9gM1NpuUqIS6C8VMg60wNB9+Nf/cwpMsr8gR7HKSaV8P0LQCPPWuD5Jn6/1D7hgq7q
dEvEdoC2sXlGXF9pThXU6n9fGB6xKr99Bhe8Yb8x+BQfIp240VLmbypmdiYqU2gM7UI35GZhQF6e
g8bpq7pVGJ/cB14ocIU0uIQNo1XPPnB0ArfqqS68JNmECmmX50tbIOjBaFhB+Cu247XEFTPfcyYt
7OsGfSgYtUkq+BIr6lCbHWE1QxGC7aWmKNaCN7/LNyzo1iYwDfvvUtNwO9dVtHXcpUj4nBu2BE/k
UILkc6CI7iPDrev55EuC4iY33yNHw10aVIch89vwsLAiDA2jDjIEf3ZuFi4lU9alTItRZR+UWs72
JshXomZMpM0LukGv5lKJIPKxZf62k0JJbyDKI+binP0QzAolo/pk8JkFFkZMWcqTausNApUvMZ5A
IRU+/uknRNBgbHbA3VAKehsjbqy/8wIPkuW6t2moWechf05hL9JX4EyccNHXGRozuhCXZgi8MI31
oqmzD9laG89LYKoEQgBpz0tPtLW04ZJy0u/iKUgK4HePv01EICqeG1g/1YQ6ExwbH7eNWMAdmWm0
C31zDDnCpz4IX3G8yvxA6vxRd9KLltczFcVnNlkgLZAfESR8kTlC6ktrjiLQliOB15I+7zis6SNo
ejrYyUYfae2XKFtCMhT+YnC4JL1RL2nUGJwB/phsGvn3I0N4MUv0kRX1DUSCn0AmMDFS9nuUTBfz
35g8Tb+SjuyrsrcubwSqu79Bqs9Kc+mgStl8EED7nAiGK/WgSg5MBpOpVPbBXzjiNHqWiJC7L4c/
XulFmsH4gbTMc0LP80qT3SRR94cGnKp1R0Hp4BYGE582k2tZOW+ZDvFPaxCX2PlTvWMWzIhH1c0N
cjcOLgUwR/Hf9aTcEL2hjPBUUeyUk3HpEIdoVdRYmyF3VIQzD6yKfxSGf7fdlX69RNdzxfYlXROF
HPEJBtG0tvzzLq5oNg0uOvfLaRN25cLKLl8UYotsk+sTFLs7WDnsu/+aZSjoaGX7wW0b3k5OA/m2
iI/FKKrE3Dh1l6dLknmaBnlaK7byY3p3lzmnQy0bPXiXqa3yNUm3ZKJUPXXWnblmKpuSnXM945Sz
FWnjbirFksrQzrm57G5HSVPhCdnd5X+CSayMEd8tFbdAj1agx8KKGQrbWwKsbCN9NgZUSfu7fBTl
fOOM2NJ3Cs2cC7CM0llYrkZEZx86r2+KiN9fEGZJEhek+Tlg6XCkFpj0oGSBrh7wzEeYEDvPX279
W9zaYGa9bzGuV24axR8TLrcvaOp/MDANhAKuupl+tcYZ5pbjtlZ0KVNRqamH+eS0Op8zAVO8ZuJs
y34i/r/yjPgZId0NWkpF84fAYSOjne3OG5Jd2hknhmExy7ICu1yMLe/9zlfxuyYFBb6yy6ekeKDb
q1cEnQPVKoQE8ORsnMmY0Qf64W6+pU1Mw6Pw6co7EC1TnFvnI/86kpwZvFH5Jf+h3BYwiQfdCqzl
bEGulKUXlbe3NR5jasOixSLiArWfpx+yUvTzMbAxqOersIXZm29Retshu6sAU+8P8f6ienpYp256
d75sLfYRy5uoUyLEGPMwUgljdaylF6l3i2RlMTCYcVRomeyKzt4aeTYxgwqdwgyqwlfoZ9lkCGXO
EAQMLhh2FIag07NcyzEffLi+ZlsElqJyd6sGoBtq1mSoUiFIQCxaBB5gHj20uhUSMI/djvtlslWL
/jDQfSxrUCznEkCJ8+2107Z93XQ/OrbFTQM4Sv4p6cq/SEsvH28OHM38byx1Gqpu7g7ImupzgCuP
eAjLdex1OTIX0yWZLJE54lDlvQYESztTDAYALLRlJSKiST3v+lsPkuzW5lVxDhtMQwlKlp+0e32Z
B+BzUq6ToAfROZsiRYnQdm02zgchOxdEvGZ/o2uaC5pPRZ9zSW6MRM7B3XMQzMaB8Vcxjc0LmxPa
EAlj24BnROZ0igjZq9+Qm4qr01Il31mk97f1dj/mmLoANkAAEpUS52ShaiyLOnRxEC5raUzH3But
xbL04g7U2laQQX43Z5ehTStXn0521uZJWqP66643U4UafG5md/vehv0uKh/3x+dKsKYe47gnW787
mFdjWd79gOJQygqYi9lKQIYnVk4Eoumv+MOrKFT06+GILjCSmAP1TNV1KLYMlyKr0eVnFIFETJFD
5yEoqEC3HFRTlbeQd3RxTQDNLMEQJ4CWKu8N8+yXziy3I8Wz3vRKn7wKhOvbdKvWydlXd+QthxjY
xhx/e05T+zEmfv1eXCimLf9vm7HrkeWYyOML+K+zc2DJ73TjUbUgLvG4D9GNdPuGxR21V+3z1fia
GxSIUnpRstOBLL9ia2hKjsf85QE3Qb/XxL9aFMVFcLl42VQTxV7STRrySOjGfPXuDFHp9BA5PNCp
DIXJpFw9hBl9on7c2Q2i5DD+s+i2b/b1ENvjnp/gJ/y5dyIUweI19RJahYVvUQXD7vGviiM2LUtv
HeQ4Rn/NyoXjaRhCvgf0TMHCQsgLcnlzOEhifwgwBQ5oCDIKFmvPcMuS3qSDm+SO+hxMtcDP4LTu
Snd2z8bXiNDYr2UKdCVxVdoqt7b/j9x1I/Ua8qfRqs1bArk/Wg4qRlBmqoZnZS6YmwHacTfNWzZ0
Van8wlpqEwM+y8SZPWWAZPNaiUfx87hcaAfmwRwPJ2l6lmOW/5XZoCdy56lnkCkroiyVhNpp8cW1
x5HiAdnyQM3LwjBjm/feqzK0uaSJMAn+CWlqXAReY8AaEGnWhLWcLfiEFtMhjMDbUczDKkSGR/9d
1RCLSQXQJUypj7OECj7tN8yk/1Yu9R0T6abEKNzYA4myxBuk+2JDeY22yrulxyiRFSwvkapQpez4
AXEVUTydB0nXUVVeSlDxBX2k3beQgu+PAcZpbO24SN2pd1rdrcqXDwRFyzeK2u1e4FuOMENbo3+O
aHViSvOTnXLa12tFbBCETPA/hix8LF6DXa858m0sVOxZJ1TYjXzmv3vizWX99eljTxKjXVOtgAGq
yhPyWjgubz/5bqrTwzc5ZZCSCKtsEcLf06O9BeMFMMmoV6IBsAn+81VkdoBOuFm38cnAC9T3IjwO
wxQG/2zGV0805iQQSdncpNFrEV3X8Xsmhi1j/hNSmo2nj/Z/GgSeremgfvdNT16i/2lW129ECSsH
1p/2daU/2xy3Jrai+upk2tIMaK3ibRwoQTcW2V6w53NdTdUnjIrmYSKTRCHZaoKn+qwlE2V29WI1
m0458TsMjsL9QTxaVmwG3mXYPG7ma9inv0V96Dh8VYLXmrPuojulo2FC6p+Zu3rYcSFI3MKHdbPW
s4O/Lc8Uv+83UQ1C3qUuHhMwQtORTKTL2dTZfK1E4Un21IkR+K2wswcCmnkUDZfkYMb8d55t+vWh
rOJ+kHGgCYmUaQXxposn3K0ekf2gY5ZqDWLq4Vtc0fyfY5d/c748Ywph7zr9+ZQGuteon0vW1n1E
SIcqhIOQUd/0nK226MqtwbtP7Xo9knYfSBWfnb53PszXtaEOIW3MZNGz2jtfEnC/N4mvh7i9eNLo
MPy7eLnuz0hFeMxYX21wo0sRbGqCWyfjc0vUYJPFL7fThwE+4phKqekKd2h+TLuRswPd0R/06sjy
EbFDHRkeurqvTRXBm9Af+DgFIY8t1ZN+Fn+72LrX4YGTxvN7QtIKhKdSpmvbtAgiOvQJ3KgYROE2
bfkWO1/sjjatjdH2fPMI3tKF9t7iqQ5zZVJTY9MdL0YICsGLu4lEcWZoPiSmt77LXH+mrquBMRkP
W58xJ2t3m/Kbwldt477UVFKxuBx1sA1AKFQ42mAs8HCNmktBC4Wdh5s1Or6CqH1qSjgxm0dcxrdr
BPpUTxG9TsBHnkd8cKhsWMGiGaVL4XpEG8ia/bw6tqMHdHqIUL1SU9eR/LDE5MtvB8jqSTGB7/HC
pX6Vvld939T7yENGHdOPXja/QX8SJi9gcVusZuR2G+vaMXOeHGW2sHne2DzmEuxRU0I1KfOZ/gGf
e5fTCbigFiKKkfxWRcIznyBenhDHs1adma9/uZz2RBiP/FbZJcV+ggwqGNKYthr+HUjdC8Lju0BP
JjjVgyMcXl4qzaMhMdPr4KXHeWxH9Yh7bmMrbXXBb/MvLoCBRQB1eZ1xje9zuiHMQavMosBSj8bQ
E/c2pCNq4I7MJQgh5Cbd1/ji3zcdbT+nZ4OnAdifpre7f5rDop8RvZpY9LwfAOZ/mZrQOqnIWKQ5
sfhbHsJQdMF2ijlXXYx6KAaebpxSGuFbBjjjtzH/TUecyVYKdHXCX+LRniaaCfnShr5MeiIs3n6R
iDgx8CmrugBbOZn72GM8YxdT2WHlCO476/kOFCjy9SXhTGkZ2fpwuX+iQZPJB8L5tEG83tQAw96Z
OHhHydkQfq3dNn3qRjyJ6TfiFyGmziZbisjqcB6RMt5LoHYH4RmV+6M0kyy3s+HkiXJDS9asglEZ
fY4xYWFCtsfyQqsle12Amcppg238KP+McQeq8D47nY3jZw9YE6mlwD4ffc9te39wGkCqvbXBgTD9
6VB2Mwe5vEJRya18Ndyq/zjNAzQsriG4mvFvYdSIXwW7mRXZ67Tne1jYX8GO/zwmgid3gtGTVNpz
IbBjiGIPzNlQ/HTl6zX+MMTS+IXKO64gNdIpuKkUCpDRiXC9rYWutzlpeYDSp9i9nmHrnlJ+lG8a
Mm6a5AXpAbpwGDSpCNlNmFvXg71JUru/CgjiRoxxxvnml+a6LWgAxXWlJlXQUN7HFJUtmJlw9IQd
O/CEs5V3Kpc9mkAbYjVk8PbpqqKaxsQR+qeywZGm81SvioFYoa54QyzzqLJPyco9ru7JLpq/QOwW
KMl2pCefEoP5F/EKda/hlyqNsydFniHupfRcH/iNV3RslqyQAzwyi2efb7S0il+UWDwx8ve/Fn5Z
UHXGQu5Un4a8VGX7HMSbqRZR/Fwk52M1R/kDfInxIpzuV9ks0xXOF26ajSTEaJPF7sx8eE+3a0nM
iLacPVanf+RWHX22rvaedZc/bRAtG6ixlPm3OJMnLbE79KVlslGsS5jWdVu74RnmTYj+sdTo96sy
AAem9u/f9kdUsXzfO7MiYWNATT/cD81P2zZtKm1z1S6yOAALZ0Hb78Aj5HIFUKMSnvBDf6cQjo3y
CmSugppcFH+ubcLgmwU1bn2oaVqDfuViwWmcBUSdBkf4No8rCbjJf2bGj1mCATTFIaXgGipO9oJJ
c+m0gSrqvGlFUz3YPMFPS1ScjXvvVzIpiBHr/UcRCDE6KPU2PWWUYUQetEabQFTKq/Tuc2AFwimp
gzLWi+qzFONYJldWzRtWdaMZ5fOY9qBABdGBMjtIt+1y92/aU4vQtGrXAsbAmXL4Atmoe0l9i5ui
o6HfW5ZAo2CuqegafoJDx1GMOVAAX62vvgHqaLOnQw9Z1fq8pgSGsWN0SgvwfR13IFQNp4v/UZJk
rQW7cSOeF693Ls1YQSXRQzi9JMiBrvz+tVqTO4HwlSekl9vO1dljDyKQ+eBKnTUvqKaO2XsSg8nv
dw3xtIXsSoLCJeEjqSimHTy4zmJsEM6gQCxVyn817YBjWICNv5ZH7VLMlh4lPuQXIYNq3Hsx6KSU
bNkQM6A+qEKd9otfpbekklfYxPT73lPntQX4a4Lg7VRCd6IK0s4Aabo1uP8zBVfcW3io+cuLt7FH
N5+CgiKtPhNRXR973VqRfkpvDgMNgeGvTNshhg8gQ5v6+mPP3Ri7TaPAfZKpLaV0jCo+I/596w4g
8OMWIuQMey6lPgaW4hLLTnMPv/lx4Hac3FQ5co8VjbsKEXVMm1gH9UQgprM5N6J7ErZF6dKPBqN2
E+Xx2cKvOB5VxvTUCYjsEBqBMNkb9pLqaDd0FnQ+vGG338wVEgre+auFeuyRsuW5pn/UF1n+43Qk
/6hl+WQke3yEXN2F/X+qxj+zJ9ZRkBVFOfkxwfPtSE+rQEkdHtzGveXq1TK7buYPnMoj3qDz5MGK
UK2CMtR5zWLehk0Pfp29BIl/HofQzxK2B+ZXJPNke5+4hbQpGtvPOgYFwCyQJPbUvAzqyF1HEnO8
yMz/stELDmab+MrQEg/tN471YNfdgF16GqXioyah8qf0JWwD4AklQSAlxm+hnWfkllaE8i4v5Uof
oJT7gvsX+Guoom3z45DWykRNNt2UPg4PHVEZ/GHZEbgIgcuGN1XUf1lv2cAaPKLg9GHHSlyFWhXF
EthC7mP/KuPbjrKBoW+lD6Th4XbthS6z0mR+JS+GCZ8wObzRFxD63bNYQc/j6ezkJFELG9LfJbRv
EOj/ggLvu+Sh3r7TNsXhMJ9e8Ha4ifKkHzeA5V+WQhCqOXcJsgI/i7PugvUlix03o8+BuZi4WF70
X7JLXboFqcErnr4ekik+krFfzc+otHeVDDQMTmVjcXH3Ti+8DfREXIux29Gmv6bHDPK0NErwBvhc
eTVehjb/mhYa1yuFLoIV/VifUk7iqIbtadRYgqlgUVX/iKiPGPDyM118Gs9nhzQKlRc2fVvZz8s0
1whfAsgE1br2HEEUi0JxgZEugG/S7Sh0c6Hd9uUPlDQ0SaG7UXaUoXGTIzVNtaKvmF3k8O0R02Y+
hhAcNhf7lpErGnxEg4ZJDpZmHQmW+MaRjQUzOK2MVPorJwiHClaXWJiOdGzF0NIHQVJnSzjA9Set
eLDhKtcIoC6FNN7tjbvJH+cRdzQJBH7GEx2WSMHlMxemyZ5fexTKWJXmYN6r/jyiJEQLc+r4MfDQ
a+Gdm+1xDtbjfQrY9GIGOwi1BRLB9MYUW0CWgM3/YCA2kkgeAN5fZh7KQ14IYQi2nWjvALNQ8t/r
/4AKuEPqYPdX3h3C33KpE9GCwV67PPMhSc2aRMmppZrrFV5QxnFZVQvFVCIYMqzvr30liTl1LawI
o1eeQ25F8n2HqJD7K5JT44oqzzEP3+etLiEn/zsUlFD+4q8npCazPysQs09//GI+Bd4QTD123yXU
TBSBsb9uTne1zQEw/dDcRi1JO1m1Sw6M8GZTzbPetL5Z1BMvLI805zBojGrdJX5P72Z+da1/mgnE
JkPKMxmhsKxSV7Q2bSDZkC58KWUvMqQIkIxm85JHmTA9Npx5tLdP2sCc2AhCQMgCzktO8Rz/I+Q/
7GYj3cE3Hj8bBaKwU/q70sMMQEfiIDAGY1GCE/fWr2mDB0pONkVky1Of+dXJ8mbRIq4SK2I78fUQ
5fZnSODM4qM65btjUqxhxNYcp0OL+3jsta0uxPIcBx8Di5gMO43ZXhHDgFL5v5dgQnaRzRcsMeYY
jcAh4rsV2cSA//ypUFoQs9nwJhVU3p7oC1vHBIuyGKQSZZiJYYI3wNI1qzwsu4GLJwR3pweNQ/KS
IVSzpzw4Xz+TuxO8SnItGNuEq+HYhFF6usz4NVBe3prrMEzfSwKH0pTQA1v2ZKDHhWeOdE//mBJB
AWJ+IOknbnqFyfJaTRQH/huEYl7jI61EYufst9L9jgn3fSD9KknfEHWbztyM8UWypu7rQV3Ggwlr
pK3vYB2lbLfiBSa3mopMsu20BZjGduPAF5M778p1P8VVNFZgxSZJfxS/1JP22NV8sLmovnSaoUjs
QscwH+OHe58DLFtb0e6RfXT/AgeQNZMWuCNNSZiJzIvs4XxS2MVHnfpEtsISJu7LB2YhDwqngZoI
f07r85Y5Bq5/dQGCssLWHzm7NlEdtUAxP9X1UnZYHO1tamvoyiWV+ckUVxYQYCKHjK3jHuKJVxBv
iAxkrx9sc5BuAUTgF4IXgLF/5zMV97hXSC8uDtSSqLNSxfMNAp8X/hJNKeQybnmKTD3XqMXbOs6Q
PEIlMTSL0gxpNSHZpLupQVij6QRmvPghymBajFc7Wnq+/PfIcVqhGC/xKJQb3w6ICKNaRZB6Rh66
ur0G2VZTNB0gLQ4c0iv3Np4fzhFEhHx+VzofFxTiMxF8jv7EvcQPoL7bEKijxNDSi5dRm0JjRN5z
bT6gHVXRiVIFPdjItSDhrWpEz2xV8Z0MRDuTvitAIR/JFQqZys5YKCzHN7q/lny9blqosUJ8Un1H
Bw2+M3hkD1ocqQC8tf2E//5ujkry/Qa7mWp6dwPmv08rnT3NGN7IUFgabPfE5qG09395dnGJZvpK
OlO1QosTtjldA9BSs7EFVAML0f4hcdGFfv1tDcGOCsGUA/yXiD8Jj0GzefWO4TiQK1ejvt5YO2ta
tD0fZV0cH6zkxn5VaF86aHQPkqGXhgdG++oYbrmsZ3yfiK923eB5R4N+uA+eiSofaj+FyZE9Qfz9
akKw2cFM07lI2fcEIl2GLejiBKiSqIrrarZCpaNQctpuNdcDoFG9KAXqCN6zTRWDmKzzAx1XlIre
405O3q80vbzY/VG+2KY3bLwJPD2iIso8nkALLLamiWEiVoNgn+Mdt47vQHXSMCvCXW/nbJXvCciV
hoa15wCkKZrFH+vVxJgljXqGlrPL8/dBZ/NwrdYl8N+fsYGhwfifhPKGvDTufRiacySnEmVF6Eie
0HW6czXoX62u6dz9WsZq6+MXkQ1iB7ztI60mzyMzfUzzo+w66RzWuML3eHAUerdPvd9WEvL4kAI7
E0egJP+6ZYv3yee937H2MDksH9KTXXcb5to0DlUtwjELCb46aFrOghRKWDKA9Qw4gQxU/7jeMgFC
YW9KeRTgU4BAMJ+i6HajXK9sK+MlfQjA+YzXI1S8dOTxqULiEiadl2NZ87nC49E6+unS/VFAIyW4
qh0qoqdw4CqEE3K4gN25RO9JuDynrAXlWzL2AjtEdWQ/JDgPoNsHUo0KW+zQIrRBetg7n5WQWXcm
kmzOVeleCZVvay7l3OmRdT3wN+7Dpxl4Z5A+F1am3w+k+zG26t06ISn1cVatzKw+W4BaT5kz1qLe
/ZCnFK8MKZ+cgF1V9uneS92GPG/x8pI16rq2JLFDx+lKJxzSNpoO4t7kaJnmiaiBK3i6yNLPC/lt
N4vpRZ2AoS6NgnRubx6lWUP1umm2pIB9BsRbXlbRTclzmVyzJp2x901VHp+cqUfy6M5zSIc68ltu
0OErDHiSolwHGWL4hbrC1qK4dQ/sSinvaYtTBu8/dVgd9aG1yKqA6kDDSQ8vG6CEZ8wAm+89at6P
kZbhqpm6OmwrZtNEsf9vxu9IGpB9IQRvK2g9vppF58pnJnoGqZlOdefRKOGnxYRqI1IypuhIBKb2
22PvHQN509OX/aXRZgzAJMlTZe0po8hBCWrcYqABctLFnk34SNz2mLoPnhpcm3WnTfU9A8tTMN2u
lGqESeCg5Ksg2WNF0Qn7NFuj7Dp/rj04UjWYVFNy5N19Ts7dQS5gZXL6mQvKliZsYni2ml7YsQQZ
DWAnZ6yxb/HeeuXWYpgsbIqoxNLakKyxd4kUD0tg2yWRhxs97hE9ZxFvyYv24utZZV8llkANqVTb
+GRq3NsfYc6xYBB9OLpBOQT2L5B1YX0YtIWKai1dKdLlST7fr9RataOUdmtMYOsfRwKPrhWyFsRq
PjYWGS9AVIWhwcb+XKMWFlELWQenz1eYg+si+v1UL42m1YstmjnsUPoU60Xt4kaq2Pq3+L11MfTa
hPhJ2H03s0+H/CHr1xnIniwSKBaz1DSghzBaEocZTCwOovbTF7PTZ3aYOvSRUbfZmK0WR41mXYaj
+AS/n+hdJQKmtExdELgRVQKrtVlpgjxEogZiSUGPJb+MOsrrTgELWNBbThRoU9Z0lZYKDmxTv83x
CBw+ETtorFeUNCLhG3q5QjlpsHuel1aVJ+TkNe5r2/TnYKP2u4//UYumMjHrrc3e1yvqXRA4sZRS
Fy9q1GrAU2B63VROb1kFBkaX68T6mIM0dYMjOJISlCgl/+PGrRWU6q292ma7qb/1rtIThU9k1Myb
8SDdDqji7e2U3sPnYHNILjpCJmgyUHPLU/RxOehdqEKbMG9HlYRp/SQoG//uci9sVLwSlvXNc2wH
pUd/U311B17cTO6bGO/4jjumfg/TuAqqzKxz6N2IvUkxYpQkDusFPaKfSVxHGSPTFOejEXek8ELB
Yexd8J9vmTFvvVNglTR87d5G23B2wL6bRA1kFv1JgHAfOBIkWTnk9Yg9/D8zByHxMVM0fMYJWTRR
IV5WJoCs1JSgcrRGoVCE8pXfr+ISNUSnLqbjvVs7X2XLjmzDo+ppBrOYnxhqBVpSsCS7Wfu3XKMq
45TpEk47guNrtQ4QSBgxYPlh7FyxhvqGXeB4/fMooCP5MPYnPQE8vWxpBUvlMa94Ml6x+UO6F4ri
CvC0fy0dYvW2F23FmbjHfMmJV/70f9HEV+Qpigc4KyeUhSYugWwV87jl003tIY8GXRWP9cXB9ip6
SdRYoCHQyg7qlMxiNesoSObSInsBxfXrVw5Io2Yxj5fdcWTDfLGOAzvHkEtfOpQgmZkWVbjNhqgD
KxbSfiGZR9u1oa0wNNHg5paObrGNQ3x/D7DWoIMKh84frjfJEW3Uip8+zrRgQfFgwXljD2QLawK+
iqhrWh2CFQV9nI60Fg7mCF3Us5z2O7BEELulZui4BiBeBXiVJUPgelxOtHdp80mqTCl/XNdpHZDP
W5p0f58Y/MrArvwni7pBbQdaQtcyFp0HVWvd9XCtzoHWiS0CYnZSt2LpMs26h7MgKtf1gzkzYFWF
+1dCpPrjDrnW6Vzdh8cng2fqr3yDn8dN5kfCa6cKyHkfO0wsUqLQJwoliSZKReLbjM4Utes8ZYzi
rH0QdyB4XGREshfT8G8iSqOdn9xhR52sXhBYbYKOyWISll8ZgtskLGcZTGY1TZwQiW46gjPjLCki
zDTVZGzOQ5ceCA38GnXtzo1ps2J7HbXdEEJGiTWa9JXHzRzvbTKZ1lQHlyiueC47/eSyLvQb0W8+
QFaajJy5yoxG1TR/VswgKK09FGpoVlD93siBKK3tnO6iy9KeOSlVB92DPhp85YTL1Ft5gsiL38GU
SxOsV+wbJRGC3vDDxx3ORcds942WQOxibOYgR1EyTWPcdDgcjsiDUvUcAY+gG8/kNFTFl0tgPuCw
rAIwjlI5ay0KXDoXgN91A9y2YJ7mOWDolSKyK+pQs/gMe+9SkPsIR3d/mSj4GtfyNqjWja9rjuaj
UCItG/ejIMZsjRPcQpPgS0kPr8iKyoCEspaQPBooTrSiARtvjc1yQ9tIpENfBnxe9TiwyhWel3PA
fA2yuZ+2K7XMHFu5zsJ6nGh13GJMVvPObGHksP0/CMR5Yul5zQSxfMWcw7FV9s3ZZabWffhP0cRU
l6Uh4IMSTlyf5bOFKRItg/4S8OJgG6U5vdgpnDYbKu6aLsiH9Ey6fxOdciuKBE5Q6BRTlmmEGSwG
T93xBn8+Y3ogAFVy3xJRZY6fEiM3eDlLgFEdAWht4VeX9X9MSA2bCWFiAzfzaCkqba5drYtm2owQ
6ncfQ1eHVu9uotetRTPAp3q4ZsEUBJdMnFTSo++rz/WLfzh1/5ye29UrjhSchq95JQ90gHrlENs0
fQJLRRWQL4XXNSvxgzvUAUlFGCqNJslvarZu50lduCgliIIG1fdNp1YA59p9mhKe0sq5XySjILda
Wqc98VAmwC5hK74Xcrk2mH4Tf/Fady8Pa4fsp8ii4s2SQEbZmSrWUywvKaZg4hjOyXvpjOwZo/BF
/cLZwhxQ5vTHf3fnr70gTna/m4wbaKZgNchQ8ROOsGe8RfyIguhluxNLEGI+sLXV3vI4jTjBP0rp
AqpaK/amMJJiG+M9+WjefQCKprCTsPJQ7LGQVXO6TEdgKhBJhx7f1gobUju6fCkpb0qYfWbw3EhT
uvNXM+La2L3tzNrPyzoWjN7feuH+ZBj9dYm4vSTJsip/5i4nk4MSTW0VUJEx5FENm47wTyESERTX
UJHKxObDdqSf8rGcj6+NIoMsDqeTglSgRoD7V3lI0l5Fn+p1QV7NvMHTdTc3iqpc7j1HZnneY4IG
A0X0FngxDZzNd/BCScaMV8CqHrbYC4IPl0jw9JymLOcmiHJTWB1X+A7QU4TTs74AOyL6x5Zw/6/4
xFb9iOJ5MjuVViSmuT7AAD3IkqxWdzAdzBtL7/8Xv7RVyRAz+PwUzEsVMtAtg/DDkaw4O/WRbKHy
JSYp6gaXr5LyKc2m+73sNecyDPs8zcOC57kpIIUWAMgOFMrHnDmWn/oL3B+eOKCSDFhLYk4RiTdq
DeXNhl2hpRtd7yG2JqDufkX6V1z7UN/UxMZJWnHsUslkkt0GIYDMIDOLWsaU67Xkca2SXz6BkbEc
x9AzVckxkJGLUKwhhtD3B1vuQfP3ncli4Pgc3W10JbT5gl04OAmDyiWRKCVB/ysTccGAS3XzqeNU
GKKv4ujdEgfMRTQpETT9gftGJBgAgJczaJkDLS5aRn4ktAeQLD47f039/iM3k5pple737jHL+Beu
vYnlPDScCex0+Uo/lzgnT094Om4hAPYP04D66Hw7rgEcee5zHsNr+KyfrVp2zCY7uV8Mn6ytdfoi
QStkuHsuS0uyhwRe8Uf9XKS9AN1PAVVc1kfhd/mno6rNOanK5yE/zGPfja/XFWZsSLF488C66Kj7
e6i+3gakZSMVHm7am7MKZquB+ezyk+jCuH+1ZQ7uoZmTvYsnv66RewYybWfYaoe3tKTI8i25HQge
NW5lVV8YbLpUsp0668ZcSGMUZ1iAZXE4VtAua38HhQCjvoligmWrAAwq6tYIIV4q3uoR/urLL6GM
AgAuAmC2MOSfABU+WquCiP6gPg1paKj67kSlCGfxrUO12jI7CD5wyixNuEVF37aWs7yJ08FPHwbP
LYUCkQiWwdzArL2IurQfO4VYWpmTqJh/jlCuE+9dh3lFnqpVU60bdXw4tEudgIUATg5RLW7Fgrhw
XVjqrlGk88uccIMomTNzJX1oRH7AYDWgwBFTMgnAl6dPgtDNeUF31FyyFMP0QEiS8wHWLXDvbqc8
nhllmFKU70Eb8lzrJ9IpQ2gzh/c+XhE5KLdKudDteHq/wUh+B7swDzVk37cyVIJ4+oS1Jn5ePGim
7fkWK2BchYP7LDGpvqsEF6oK6lo630sk92NostiW9jmxbaIuv6Yct6NpX8bQ9Piv64P2Pb63WUaB
rn4MSdTQ7g6Ga4J9s5DBGNPvQaf42m+Laa//F9z4FLV9/ZQPW7of3PzegSOfxfMaAlQ523aQWJy7
mH/peYdNRBv0g+vdC3Ma4euxAng7KWpsc7f+pQAktRYgPytfeoXN+RlCCD1TRvD/GT+O0BUNwpld
5sif3LsK+qNKJ/TD4yLKw1aQSifG8vwy22sB59Lav6duYV6iKv48renmr75mDYKm+ReklaTdwy/D
azc+xFH3pB4lHcOW7kFjW51B+ke6Fq8fUABUNg+YztYyJKO3r/4EzbMcBAsINkFZentxdF11q8x5
p1aW8i8JhbF0wIOoTBlVgvwhLVRVKpnQA12vKScjFNY2dl/NIoOXuqTFpggZqnbtcDrTX4N8gPNG
1H1GolLWKkf4WHsx8Bmzo5ZfUhaE/6mjt5qEPxgwCYMCMGASXDOukB6Y3qoPWZKnhM2VsKRjt03l
RuQ3rMxvfQMM/4SvIWE5kyOPHQKfGbmRgT6JIl/z/WSrZpMwm9pRfTLRbU/m6KSwSGqaOa6Ahail
Gsb3mVv64hkfinp+fsR2JY/KJ+NR+HtI+7ak48NDXlR4QrOnwuKjAIx10olLS3tn0dnkDZ5M7unV
uu5goQEQWUuOzr3QRbXLUdUtFI8bAUHludAX6qri0BvhbmRKPBsSHGE+MRMe3lyJPCsCj8sz1nLe
ylZiQALVjWpi038FPg0SJPiPk8OSt+1Uez3VEKGjODHiLFr/uN4aM7bcqS7y8PShMHVwa+5fmMTc
bGa5QmLD+l5S3KpM2p/S1uJZPfJw0cThlh1T9bV6ex5SpN6D1wtkeTss034Xy0fcXqBAcM+R53bB
kQZpEBbhpqXkV8DSdZwVGSsdDGbmMkebMotQWF02YLFbkBBbdIdoTe9OfIQrHJtO/YknmKIosfZV
OgKBM6yippfJWDvIg9jELeQ14Szp/+8npDqxx6/jzUDXbDIMZ62rrKXTgyea6ct+MbEJXH/IkYeG
qTTIVt2nHnr400wI1NW0+F6JBoER80scKwW6CRTPgkErOsKdONvOGXWpctdjljJU7pnLCrHwkLJQ
ZLIlDBI05C/IuKinZr89nYR1WZ/ZxH9/+86s86JSTpjM2Wmg2T+J2Q39G/jzbUiMqEM1yOLlgh+f
pg+ekpHgOmCooovcYnede0JXpEFR7Ez8PRt96yO7l5at02mCyesfPVV44VfKu9PLflOk/SCflwrA
TuskkCWAPraSwOB/vsl6aFYcvvCLfhxq/53h7x6dIK0rOXWUr6Pn5scmk4soh+3SKUhCAwJiBY9I
9mliArED8puNaRBsuT0mvVGrEif0NlnKHEpyR2+j6T8GHrvAb4uZ91opno6wsv1A+16ZpzT6cYK0
m79e5928LDZdKH+cGzPBevHdJnoTFDJpdlImBv3SOjLnYUPqSBM6L0GpbEdJb6JXlQ10gpieKkWh
oWIr+TlvmB7UyUhiEdbzzSerMVbOR0RZA6lrhW8ZHJ/rQavvtNfjt3hfgZUB/tiUV1lXN2on7d6v
VikR+7TNmvkGSjnXVdykMI+1h/2TBCWeyKLnRvKe37kskgTTyKmvyjua3mZOLfK+HcL33D28xgnp
9ePma0IM3NmASUWMIaAs4Re61MrwDx3IRQD94OoGLBvJM+oRXnKNU4LPnmjkvytpMnV024Pl84Le
os8Po4Q67XhtVaysMguixMff2kWzODx+95i8xrHML9gR1iVV9sfxZEMagtGbG4OeXfdJFNtNM44R
u7+HypQTRkf2HD7/ArNq6h2yvw+XMazxzGxpi6mcIUo1Bs0SCLbk4wogNGDIjS+Tn+kPyolDsmZU
n/aQHkHMAjAbHHjF6Q0ulBv65xvrUGep0qxgUEsxk4lhYnueaGeA2eSN3xsC98CRva0wNuRR4iFe
zaRH0kPfbRU18DU/JriLchX9uXEgPguPlVL+8paCaJicsQapPFl4KdIfScvKvXaAWJoYuDw0alcS
gZhbCuju5dHi0VafN8wdA416cywNtYuNxTfVa/xXvT5HB5nFWXP72xALjMLqg0eRLHvE1H85Jclz
Iq2tbvk7CU/iWBRkYt3DgcyMD+UXaxTs8nYJwKTeGXWTWZPzgUryxdpTAQM9mYzHBqOrCUHb4NHw
zGByuGFne7YnoZWGZS+417j1m8UwERAK3kmzXPU7xQFMC+ofRsgAutLpmjVgu/Q3asSRz9h4yab4
cbaA2JXJlrttvN1KyOmmiZSKpqZVlZRG/tv9jt0OOgOQ++KMhzPSfeqN6Y9sy3pYSesfDi7Sz8QH
6PxjfOJ9Pb1PCyI4UrKXL/8quCdXTzIGqRjIi1+/4jrU+/+8wDkE06YWWoDSlfOai0Yx+pfQ9bhz
6xTIf48OJlMsJ1pf/wNto44jrpZYC1OMZ4zCvtyfqfBsNoexosB8Kzj8dC8/yVruiIg4P6myb6lm
WuQuGtqmX5RWzvQlbelfQSI/TYQowmcR7RMgeGmBqwCl7cvy+LYzee9qWJ5Oy6iGIMad6PeXW+tX
/D0rUb2SqEavtOU2pPDua9filkOKthfWjURDJt6QAcFONRjvOtkCjHVPd5rySG6FLhFHKhKO8wP/
ZN5D0Lp1QckFYa9b5r12oPmrEZ6ICVkqlraMYSjy/nWprwhdeuo4pT8nUgTbMc5HlXwcyqrl2DM1
kc8xuozqwmimF3+YBq5Z4HfQVpbzYb7i4y19xTou4rpWsQQJn0BqSxSaWhyc03T0wvDAsMXHEOiN
lD9c+r4e9aOIUdidCJDWiu/suOIbjvFbPu7JtniTgCBTFwU+sLnUOQG48GX3WTn2wN2jH4mmiGHr
UJydUK2CISGGb8qf23iseXDobgdMNjL9nR8i66M8N57nOzZZJG8LvuM+51jJ/1RsbGSTuVXhadz3
hfc0hD8pgQqpthP+zYjsiOxbsUpjAWHylnAtdFBzxpHDDeIsiN5+7rSMMaicEZbbw1gfYy3iJJx/
f8WiLCA8MmS+pp7wUChVdI4qn4fMV+GMFmtdAqT7yVWV13MFJLO2ymOCCpW8Mt9Z/P5os2J7FaOH
t9ZWvj5RUS1jkJ3yjlBw0asxAovWvmg4B28MIEWiD3w3NnYDdASmq1zz4fLEX5vsmV5IdzfoWSiN
qlptjjkDb1Rhtp3xEGTlhhDGHzpNmpm0/Qxf2sNIRxYFhi5i3y2Cjm2uGhwYP3zlgmAEMOQQpQGj
Cieh+vXQY97ZR4CtOUoXiXoN4ImxQg7Aymn3Uc5TjF4HyFMCdWe/Hrj34Y8i5ZrxqQVOR1InwApP
DcKZ82ZR/V+T3YRPzweqPh287lO3cm3T0xGiUS0KCqiv4sXAuDEhYF2c0OXa+hA8wjxXZJ2cqymY
Iu9nfbrlDLCNjaHWAb0SStnQkrjVWVu+KsexEyUd5THvdfHHak8HsJ/5HKnO+rQqAH8et1RJzTmO
woLHEmXU8XFeftHxnWNd1QRYHr2sNVPDiE7e3B5d6z9dZihdkM9hU/V4RMy736xbn0yQbFoMlCrY
iMEzm2UH8Hooz0OSxyL37BTMKiHYbvTGwZ1fz3GFnmS6pmIHHgGkPDNSuiQxG+dLJWqYtI1x+dgN
dIaMp9+mnfAJJx0E340Ew4/VztmXGHN7PfK5l8VXpE91ufApPFCCTZ2OOSvrRgLzlgfiHJV+i60W
Dr6UKZ+vFuN1R2hQtvgHOWPu7DX7M2SSGHbbUAtIAiZQevGKfq75e1vcr2zlvZgFlv/8hI05NVG1
I6+sezEAIal/eyX7Xsov2h70l0xYYudfhINgY4S3HzLiROaflI64/ntAbtbTzUyABw41L4Wk7hJ/
UK1Oxr5h9nFYsL0qtcGdkAQc4JCh3vOk8NH1v0mylYp1idh6KrPOAmbFMq+P0cRMXTpNEVCj9GpL
8r0hvpBRdsb+MZjr15NCXqqJK/9i2TinoNM4KRS/BDe3GakMrFCjp5COkw9H33PJbcPeUvf09KPY
DiA8MJbPJw3lUn73tVBnD0ob0aceBCoVDZy9Muw1Rkt5gMJpJFWRSEPfu5TcSScaFbhrW8zagrbY
HIZ4K58g3NKu11ntWva2JRvpc50lIm/BHzqZaU7exUSNEhyU4aSiYBugczvkkv6kdWQrBXfHDQZN
g1H0Jcri89em5JKIiMy65CWWsSoAB2mI1B1Zl+KiMi4dVfPWnVWSwynsyOyD9aalysQZzkTz2pwW
HlVBBk5uBEsWewq1Dlg84TJLHZFKkl0MTS6yWFmcIUUUYkCe1X0GRXZOEpzgStBZSGq6G/VoYUFO
n7LaFisp2zIBF5Yf6D+sd135H+p18c/d9X6Y1BmFhtfZgc/LOQ6PxEI8IjkAUzNM8BjXb19s41WJ
FueZvlKt6ZqokF/Oz16wm/pPIXHu9/+FM/b6STUoQyitzHvfTv/Ljwit5fhs50UxWW3vecd895h5
011ALfAnhvjS1gUmPJ/bovhwqabHFoiGoGbN1DDfT3YJ0VZhS2/Yy1vgkpiDsYkf0IV51Dhu4tqu
8rwxNlhQaKmUJjto/GNzpBzDHPskHrPaLa+hYN+z2CkWkM1bJvmGxvSutmxJcXGkQcR2f7Ti9o7J
J+Zte1wJTFWvmRhZnzmOTlSKkWj0yovh/gCbtgbaC9ej430RhSU+xAuJQE2ATWP8/x4uArJHQHN3
7lbrw/xfXWgGgIzqQfM3zCuBUdGVdbk4CI6ajOw5dYiSWfKmp0sXJVmIC6X44iTzn6AcC2DABrXP
bCgiIBuNaXUJ9HrrEBn7u0hQ3HNzCacV6+k7U2BhveHS0P8xUmSKj/02HImIh2BynWm0aDl4+JeB
IPFP5jN96z1IAEfwBY4ZwY1ndv40D5IADPRM4U1uZx4hm0siz2uzTKoRku01YhxESLkNyGwarLZC
oaVKfJayc43htHyhY+Keo8IoulAQEI8Ct47W0DkY5vH6234AO7h/bN/+P44JuY64uyjZ6QRssC2q
T/NJk/Z57J/6OU+6tpQ7pU0n5+JmAUmYV/5dGeYk65ZpcQc/lnOlcD28RoS/6rRgiG7JSYs3UAPz
f1l/F17ru5jZ/6XOIAIKiLft49eOPJn5JJ9h4TyyyWKf/TG37aIwNAeuoijkzGohzpdPRmLRsSPu
mkGf+yBJR1hFcZGMkd/HmoXixGjbs3uUT84uuxR58DiwwOnwcBfj8rXeTJcctuSw3kfhUnsQWVuu
K+UXZUrVQL21oC4cdr9/uSgtVbuT2gBUQs3KTIbomcGg7O1IYSRvHlFXMPTV2bKNEdC3EjeXIxWv
gLOb20KneiacXFPR+ni35IrJrx1882ftfOLhRTldvR5/bhOSXtJ79R6BO5uYALYe+xURkcsFDjFO
LsyeyPKo5NB68lBF1IeLgASwq91ItA8NeOrxN20+B4a4atPGG0w0hvtodzUOAMaRMQS20jcy4tpj
bN5LzhIr0ZVS+XjcOvaCWYAJHR0a2FIX3gpO1bb1z9r5volkm3V4j3nKsYefK63QZLlEiOBP0M4h
Jp6o+ROpKtkrQjIZ2dN9CHVoiNv5aT6eY97CHQPqMZ33inPKXknCZ7Vny9KJZUhCevDa1j7y68vv
kXqgSp6Z2QIIWldY6z6JeEhsazbOESVhDsVCj2Qnef/9CicfWHHFvnuaustbtF/Q1uC2y/AR+zkN
4yi8pH0mMGFFK/FmAxbqLkKmNAwIbvb6WAhtBy9+wIDWzl1noUblHJkcxBvpeb6Z6eebRLXoG21z
/5ByES9WhbTMoyxXME0f57G7I7OnRNzBl9X/RYbPTDpln7X9kl3cJAa4e7Kc4VP11j9YWW0p3FF0
/QUhyYe+qdB91jjiv1mql3dhcj59AGSJx4i7pRkoPD43NgB/MBUAibBOX3kKBhhk7orUgi2KtDVh
SzAlwRHg6KtaNFLivWyjGqNKegcteuqbbMUc3naXWmQ7jC9+xifRkTrfp+Zc+A7gc7v9uO+VshyY
4+WShZyUXica5Z7MtVaM5Gt0U0J4vpcaJJk2MUhi5MvduLOMYKJdoE/vaa/OQQ5iLN0torvKRmCp
mRX2g9N+FndhryUxd5U91qWrUa7PDosRd9oM2dIhbZtKzrVjPOjFAIbg7JyZNm71wi869KGkDa4H
CKk0kUL+11IMJdifCM7Md0axeAV4joASpmt2THNuib9pzwut3iq9GQ/kMp8jLRs6aGZuJctHoknQ
6Nqwgch9uN6EIqWlenntctSRGqWvf538uqiZOEFC1oM54kc1PTKRRpOWj+nno/6yD1CwJLIuWqUt
JmKxv1rcheI4Z/RyjnjvCxaoLKS/WgagB9l4DkbGMJpWAiRXWUEpaoJizjhxFAJVzIoUOy9+7rkx
P6YovxlebYkQXpx4G/lTHnjuPheYwoMAjGkjAgrosEnSlimmFZhhlOjs+xNU8KvQEWil2ByzgZrR
Vb2iezWMsBR90f8yi2OZt/PW2t9Y7ZemIHEZ+RSBIluI+6bi1hBr5sPz0K5FuCHAkviYO+v7LyB6
kquiId40sGABcl9sybFNd9FONbgD+DDryjOdJgT7N1ntOZTXdILemdMw+3Al8rm6oMi4vUMTYXwV
lb8UsgLsGju42dyAq2VRKsN57RiJ6LrGjrBDNzOGUNT+InyT+jM0GUiKUf8uBQP07WTvEn/xX19L
HLO6c0piNgeV4b3z84XtokmsE7ln2vpUXfCGC536/wUMQF43ifrHqv80ym05izKKncnM99eunl3z
I+MTns2QIntTlGnOMuKvKyKfT6OFmpiBzloX104ITDHP9en8WMsXehH2F1rx6z2E8MuhBtPKOPzt
LH3bWyw+pCahr9rDbSa13i6WYP+UybtxhoPRglKkMVdcsByT9l0HCKF3czWSYLTNeYOyqi0A6piB
cLuTKtlidfKj7uCeKfjB96bDljxzCptaQ57Y5B6LxTxYB+K+HqRyvYFnA+0WMjTb3mp/QlVR4oo6
68ZBk5c7VoHWJx0Pq8H8bu7vQ22fHTMN1LcJNCnvaMzcLnjV5ao3AdSd3xCpT8uX2QngKpSSeB3p
YTff4myxgL4lwcslgd22mdJDNzvZvcIeuf9m9lYIzpDuyrFDxsIDBdv7OmOpwchXBVNPNjBEMvh+
4QdOr29dZ9C+P5N6HdEiedZb3Rwxy5x1JXPBHdqtOBOWDHoPjDrpkm+S8x2K5gudSfEV6b9t7gFi
s6argDhPE5fNuIFAgO/LVPQZs7NFNZYdn65yD1KATKTpDzYAUc/0OT61+rpE3x70psKuB6ozANvF
esWVXa26YU2JZhMc4SJeHIyt5BKK7z7BsvcI24z7knG+ulIAMbnr8fxO+EAaBF4VVgKzMRsL0b4f
vHCRrZgfPqwo2QZJOxmmDF6GSSFio/J0v5n0+zp5JAh2KqycXrWivReUzWQ157c8y/yncex7e83+
+v1Li+wMRg59wpVVSJXDi0gL3yezn9TmqDyF+SiB7Sxuhk/s2/8L1WpWfB2ZokEcGys0X2whX4fn
9XpHuvh60v603jA/lqmmHd6hAYmHkwUly9vlM9kK+xf9wBrBNqacvNcNLqp5mwRyL6Rd1W3DALUP
nlfTn9VFFvW4xAkbo/b3d7/huMZqPvrsOh2Sgv/ySnDQvy4R/y9W9/rMPO7MNtIlt1Rvo76ynPI+
biV6MXOgfk2Dmd8GtDIbG/SSvBoH0XQmVHCYkwnmdOTQ4z3eLAwxmfTqqrwvaa61eezkiTEDHY7r
pz3wRLbZTVWBMkmZFqP4sVHJZsfk0aywqw4ivPO/xiSaBWLNgV5pV4lUU106+a6tpvIQS32pmAEi
OMg1LeLqgghbYHv2XNkt4m+/QhOjSICrAhazRrnoTkqby5gzgmNlJ+WpARhVySg82mdcpJpX9MtY
Ge05bwWBZUXhen7CP9Y5KbXPRhKQzvGLjPZtk2ySrX+RLYcSsXCem1L6B3rIhTnsK1ryKLJlVJQI
ZyKaLsaulBU9XHvoKFZj4IvJmEdAuaD0VT5FVyrMvef/1tfaNQ3AeOoEBzM1sjK2SFP3bCBi6y4O
Z64v/A777uoldSm9yvPkDzZ1+UC+6xayOBECXC9wgrbVWNL8Awc+iYXN5MvO8ZMcPcVfCSkWtZPG
NLpo6tdUd2HDkNVtUjleVQZlwImwsrwS7OLraGunGeAAvO0RoHoTtoSsHxlwLTdPKKKbiJwfLvoH
njwuuHsWHi0SBAKLCvXymlDVGGL6NWAB3ddKR5M2kk4O4isbf5pYyHn9WGbZE4WDRgIb3+FV80xR
I2H3aqoaCp/c6q/FQmEjSPRJS2MBRUjOFh3qsIMXZ8H8yi84XXdgD+DX92TdLHsE37HI8HQeKI3U
SEbV6b5pZdJo1urYIZQemec5JNeMqxoZm8uL+f/J52iTG6NOwZ00QZFWYGFDrDBtc92+jUwwNASj
B2b4db/AgKEq6OoddL0NG70VxYra+TOHmLOdrWBOZFbQhXdAW9gVUvdgqaS02P+qw6d0V78ImeDy
K4mBHMsyKM7TAAgk/LBwW/YzdTp4cdpw2VUZ7K2eCfRO/MoDjXfXbcWdBuYoDgWnedLHsPPB6jrL
T3/xoNDmQ7plwGkUEzL5XgE3SA1tMkm+Xj/Wc1jsexrtr6139sKQbSSVxAuiROk3XcMbjBwfH89V
0ZARRK+30EwjU2jrCumfU8/gsH/mZ8jjnBJI1JQSfv+2fM5ZPM5SkVWUwaIlwt9wBW1duf4IYxnW
beWpNb88YaGIc4Qg2Eyy8MOlAmfX3wcmaAawjc040bH+q5D1IPDqb3/YR/2UEdkktgphQHOttXvM
fJKFTKPbtnWWqExMNv68++EYLQiAl7kMYAYSTiAYp5zGaVhYUluM7bAG2oevBLWnUDYFOS9bAuIG
ire+7bnDRlhaQudYmTuWgl50Golusirn1zOv7IjA8BT9q7M4cp8iShEGfx11DvKZpdX8gNZhbckF
fu1ZpMGb9jMAeilv0qDQTGlVc3EaBh8GOCGW0NcifMwu16eyMU9WYmFWf8oxw2ERRA6na5qpj9uD
JK/V7/KPDR2aS7EZcZgWahWZaM4vLb+bL5/asOITiYaAHmcC3ZDssuCdanru3Y5ZN0/M2nU7PDvY
PbI12K4v3XYFoIOyZ7uMT7nr2zyqUCsv+DfwUd6cjvxN2v1zU66wIprYLy1q0CbT+/c2wuib8JNg
cpSHLwWNChJ9Q1n9+vQezJV2T1bpdANDz2sOYz/5o7YhmOq7J7LN1VEnSyyOP/xaJn/Si8jNV9Ha
ocolHqScRUAojvR2L9uUpGr3rVrdRrudt1fm0+pRbSBQ4eFInMvxafFAqm8A0jSMZ0Lj0J+XJpvB
W53xw6awHUCx/k2nMn6v+W7g2JbKflie1vazR7vhc+eb8fkPXgFIx4bzTzQfGOAxs7GZnrgXL4h1
wqth1RFFa2uOFkcvlIrH2ZuFmtLF83+9/cONZWq9iS7wTyAQctM4f+mWuCMr4FhkrDlBHht7do0t
bku52YwaGyHuytxYOSvaopJ59PBPiosd5NVrcc6gMqKkKQVyneih/asQuZy51o1vxF/tCpuaRhky
JkHWPK4Xaj+DbIQsfq7UxOuuOIFkaXka1T8tkHkXhvdohjMbg5OJwoTVwoO2xmXqUvhFS1pt58LX
73wEw35fi+43FPhUACq4Mc6upx/nK16Nxp3nXr1wDr6C9q/1/rybX57yAmjTGx5q362Hn2sPxthz
xyzfspxddhzgMlvdJh3xU/ZeGR9P3sSK+g8zDYeHaqb6K3AfCk+N6OK9hFH6fUgxeIvorxm5EgDe
ZJOLEKKs1quBqsVGtrvO5wlg0eu5ZhXQVFXi6YVXkn1NAl84TgRWkIDA9b+AU4JV1xVXkcgWEoWk
WtO+BO6zNr1UUO2X1ZgZbgDYNIz/ljzEqzjHbE0aLVgXriaxoiLNOoE6b1ZumtxNFc0fr1ysEaOD
RzqLv6id4r38M2FeNQR+QnI82h4yWXWCKjVQmCgIAtcfSKPlMXEk598CFpOPvQjh5Ya/sUKWpsG8
PNgEOFxISh8uXiuEPwNfWeneCEY5Kngkc4GjxUkRDtoktZqOgUjjdU9H7sUJbpck6VxGWEKPKyWF
hPc5YwT1e9MZw01PZadnwrSkxIlysMQIjdJc9sjcuTVzQ5dxpBv2iY2QcIva7745c2jtOEZbiaRD
XlstJxc/xJmx0S71NHAP9iMxTDsSyYuTn/vwIMxes5dTGlATiYxdfQXObHXXlU54/3Z8c4A/S1qZ
utE9qlZUzqmR/0ElxLkJd2SiD6V1DZhjeqh7gdBiAAUmyc4gLcipUXenVSk9kz3VZCPAIGHaayOw
3eDUppHK+m3mMXPNf1T0XnnV2vdI8MUdd/IyEWTVT9HPhaIy3IGKsjyQvhVnllaBuKUiPRDgcti6
XokIDYLfDR1e8CDDhnvR7cvuBE7dH6XHBkpARdKzHCvT1C9IM90jn3g8yapkKZmGgBqgIL9AzQc7
NoWKyZd5o9/IUd32xwIPGacpNLJAcpM0e+1mWuSmBbDkuYjYWW7f3wZUC/bfRoXn2FRdjdgchUp2
LyM7xOlByMvYP4Zn4/clt0fS+gJXppMjl+DYU46l/g3CXd9+zTaveGrdkzxcTONZTmwHvnsCbTG3
YkSWTAkbWEt0sc0ciSbyMwnOJthMlHVLeIJKSDsLriPCVCBXhemw4kF8cV87yxSunqhF7uYdBEIM
UGbBV9Ku1gN3Bf7OXByb2gd+RGQrvhH4xkMjPoqDdLM8pLyDsVMkyh0wiH4niqiAq/q6Vm4yOBYp
Zh1SGcmLNPpxb7UKqhKK2dlYx+CMxv/oPAOmhwQRWgEV/8sgE0HPgSgeshNTcqX9Q2gFSbFirkiR
nO5l1nWWxqWJDznErFEOtd5tekQqhuNOMeqVlXE8pUf3keTg8k8BqvJGCMj5UiKjwJO8c7Z0xE6/
wcxLojyBdY8gJD0y2nvP0z4NrEwmNu+Rbo8Q4UgKmzZ6IoESLKEtmz3eQ95mGt4kq4FoBO6ks7WS
otqGjWHoodNy1NhaVc8geHZc+Ac1MKN4gNZKOaNbDdEEkPPKJ1BB+U96vefibzFYPCeyGQfLoS1x
I1gmRCKTwXegNr6GU/MephJoNgLvkBSQWhSbwVZIet4w3lDuyNNotQhp04TLjUai0kETT2I4YGIG
LT8Gh8weU4H6UHHGzG6M7dg+gVhwsqSqy3jWME4DTHsOBbfZ1Prsy7eAzuON02oXbWJwBbZqv1gl
sHdzMiLnBSnrrwVcXR7OxWMwiTruc1+f6mbbs2AuZL3y+X87MltiAdAEMnGwh38ffxieVuiPJj8J
kTCDfzLkNSN+kayRktAWK0kNBB6JtOsB0VFTK+v+qpB5nIvcyWnBqH6JMzcPR/UMCQKFvnMlyNY/
dWnFCFCjUYzDa6kPFh4n5/nmrw3IrmM5RnFxK+L8OpxDJOniB8adEw3URZt+6aPJdUlRdycA5EoX
G2aGiMposzxoiaS1o15fKSEa8QB5Qt2onI5ztGF3hSLAYSkGAs/BBYvB3MU+Hq+BqcSrGF+Ips2W
ksvy+1HeNWPswiV+HJ44aIFZileiUuA1ibNYXHVtn+xHmW2Pn89bJgfju3NR7HcUVouEH+64csl5
vPDkP4F2rikfBKUv0Pd+hCckYbghIo2yUmCmwfoROZaPQpgtjNP1puhvkDAKPpC9HsQG0+J8LWVb
4BphpGpQhMcAc8SQQ3VA9Ajy4AUlFORuusGtDeLSDrdI1jJEuj+gUB1lGyT7CAREQFSFmMepnoVQ
8I0N6KiiAdzBKcHSCbi95MBHpi2AOYW1QFiX032kGpI8qcJFGbmsUXmqtqCd0HZzRDLyE6+kICyF
EphUY4IfAlDEmN9UfheRh/w+uZf6E4TyK1quo5GPT+q37i/joVY79Is/akw63W7IZHLMDNE0f0t7
mrcIxQYhE3FlKWt1r1XDMIhiAaRvhdCyPB7tjUaQrdbmn1FM6FZfGM45jdNbzZG+MhgrgjLEw9fm
Nz8AbbZYWJ32/yjO6N0QPSPcbi1it1TwQhi0sKLQUwGVoaBgTKXMHA26W19UEUm9sMcIElo1AvbM
aVkY3wdSUaGX4J9MWdmi6EnLfi8zPIFU6VI44CbfTBPY5lkTAnNa2ERTaRbyOlvTKQ+93USjQM99
aOeEIV/1fSX8ku1Eyc2UOwWY8fxyjj1kUrlPveILqU1bmbfnbYg+mSYdSB7u3OKmqzrmfkBrQ5KF
FDWTlJX6+Dm6KNj/BmzugAJMjcuxlisT+8fBrjwx+mkG4rBAqtA91yB3B+Hqpi8H2bp6m3elOdU7
8llidG/xFhfIYrX0XbQXutkJjq57QULQCiseS7wOFa77dRxl/G7jvJLHY9c9uusZIL9hvF4x4Ltl
ZABMAKJEFG5Lj6Zo50cME3LYOYyPADYQUY8YggX4gvqtkT04Qn4KzOuf3cjmeBlVQwGjUdPtWNLy
1iZIpqVVx35rcwTWJ9vOFPJyfw57DJpN0MKkpigB/uXTQNvib5zHYyB2NsSHtSsK9BT1Cx2crWbE
rGW6YpTTrV2udewwkpLGBFiU34C/r29fkOHRWbkpIfVsd3V93D4tpLxyTcofRjqEoHWRrO/il7L9
d8CTpDWpjkufaKDwUWDZqlcv8J+jco7hscuzTC+OKlDKQnqrAjWjPeghdJPjsTX2KyIbMUdGsTu1
EVISM/kgQdq/cOL1+T/PUCwnczjfo3Df9KYmFsondvuq2TnMgievZTtkfSGfTm1VbqRnvYFzO4iZ
msHVwvDH7tnRGe4IjdzD6nzm9ppY5+7IZp8HztZZwiO+6/F2RAXrNHPzOPKdYmq+rc9YXCEXJpkJ
3XsycmNCkUEe9ijH61UIBkAo1RHv9bNqOxxI7wqf2OvZTR8/EC5NY8c+2VeGLKV7HCkCE/jgNKgQ
fhZu7T5V3PrZ+cg5lyWcU7qxVCZEeJkwRQTm08CI4UTVJHw1OzPPfjRLIRWE+1Ds09hleeFTl0v+
Eg49weR4siXUlgx6MIlfQunLyGudH8LiynkAmkko5hDXy3S801icfUscwF4wAFCYw1MMJfACDFf/
7PzpV/Njktbwhb4aGwytOUtLNWG3boeqy1c+i5rRZIzdlFK8iwq0n6AkYpMj/SNrBjLl+v/yqVlj
1RdrFOpubAeWDbCstc6qXQrEI+bKB3RtuVN0FCIOa0f5ewmX6wDyO/925R3pdCYRYtdy+Nj380rj
xd3fEUrBNEq2W4+nkLH7rh+OPpsVtWmYXcqcclFWH6rLYjFmOTKO2R1hzs1f98dKoBXFHxdJfcUr
zUdjt8PCW1TgI0UzMKYfJPSARsBBNzltAIltRaTAYj0F0cWcHDIMCEFP6AqVkbpYRsKXDaqQJwIv
PIeUJ6TrUUVH55nUkt6AS5vRoaFxjSmsQ5o0BZVb+oBC8aQMT0sRK9ZmaSAMaZmY0tjXjmVtbyq2
0D9HrlAq4jRDYFU0TY9smcfyadxFECUj0fS8lnaNLXrNjU/P1pMiq7qttOfBWtrKUZuE6du4dofK
Ykt+gGLrD4unbI70uUH8xCYF3D7pc8GKTjphbNan5DuPiZnE1eomxMAMyFkZX3c4WB+ejlLoC+1e
rDbOONNU+o9oJQ11A+XS388XOTdcYp/DyC0cwJWR06TDdT03kaJLzHG8WBnPils9jyCveRTU/Cxt
e839NueOkf9MknngX2+0tTRI1o0atMgyIc6L2iSJkVizpyzco1jm+hQB4giW2f4/uekpPr60QVcU
79mDsh+A5Dzwpyj+olu+NbIfbuSFQAxSVZp2q8I4DpDL4c+sCOIG9mUG0oQldbtgOKNcXBuvEFkv
2aFLJrbQHfXnKGqjPi3ND8ilfSiSzoX9CpX1BT1HxFjLZTFePXP3hw92QFG5u+RNS4umtyv1NVPt
sXXdSP3NE1DIY+dDEdBvVtvEdNuse9jhV0Xfr6OstfnAxWh4GZD4Z02NnqYEMeHEOqdoQH40XtsN
jJ5CY+L2qGczQQ8/ssocG9tP/mf33nqM2boeRuCxNBTqKqfG0aEI5LJwC2RGdQrCx8O+ZKefNfBQ
GIKmmM2iL7QCDpFZccMQmlS4JmDGep9Yg/UOw9SwpAqawxJzcvRb3d7BH4kp9hRVXtW68lT6Xgrk
UE3aVUpuTnOoFaFjn/XPKHoaRnxv8tipWDEmKkD8VM6KokH+vwootTzX17DDM0zRS4FnQur1cAz8
bGdKvdmNePW1vceyxY2OjQnUxpveetaDnt8bdg9fMTaE16V3YfIjhryM+fGTCb5jYOku86FQqZlF
4uouofQOBq3skLilRIKVCFHJiAHUUfdnwTeKUqmxpQHwB5OXwNz+s7Thwz8mtHlucEDnD4xooQPW
Bta9QmdLaMZs/bDyzoicbEkwgcnxDS5hivU5f3iIB4PyBwVnC8n0pHtm648EmoBa3/uyD0b3yTAb
9OaH12GyfXZhjdA+0NV2qsuiUgFc6KXJ5yx6dUwWNJa96OUw103GtfNJr3zsVCquhgVOlfC7cwRw
z6UCkBk5o9DPqnAGnSTmpeexUI1C6OiO4Q6bUY0NMUa9UlgTvdMAIfOIK+PFIvCZmEwfN4Hi65gd
D9L3C2peCBMZKzJ2vwU8ljEsEPdrGUrt31HSD2+/ZPgn3gu9T73blR+IP0V9UCMTx0rVUOHMZ3Ax
SUdiGNXMcpB2kcEedkTzOFivjvoJyojW96+CrZP59xPkPb7Ue03Wl/JEa3yuWuaa5hOeURjtfJkE
Qd0noiSFw7aVus9+qKjwnsZ0GnTi0OVXZWZdkf2p6jxoXTNXCCC6hfbJC8Mc5pjou5JoxsaOteSo
vRjCZtFS0IlFh3yQuqqB7fBTzn+9wkI0phrweP2E1Q7bdZm6AD45NjbMW6PcqZZ7hbW0kXbEoZTM
h5+ZqGWej3X98jXamkmtvBeYTVcO4ka3+HvPFX1NidcIiiT6b+6o/DVxob/BRu3LCVv1VVc+PBvv
ckYiWR78Hm1hqZiwOsN5bua3cyl8gsBq7iqU6Q6Uu1aalQ0IMThhbJR2Ew5Ny+cS8uwSmBcDLA6O
flyVqDgIrc7m+o6Edm3CHBa+JuinRMJ/MR09RwxJUpupgj5PzmZ+iGg14NcKpxNVA9Yjftz2RGoF
BqwuZy/DZtBjHzOk04H/EHWKL4mZqene5yxZcY2VOnl9Qmo0qi47pzxCJVzvYQwk8SwsSgfYkduZ
jNVVNJAbPGYWGYo6tNUJdFkf3BRC3xhjIkXHHmtF9ufLDwU2ypar9pU1LxB6gTvjnsSfWjDhr3g6
oqJmlqhlU10xbhOK480LYrp/jxcZu6YnE5GRsz2f6mYbvwN5IDT6ykcfK40QDY2VrgMZCg5cFgdN
Z9eW97RVPcWrzA3MYfQfeMtzXhgYc3ap/CWbMqTIrchRIz1agygysu5nBaMGO9KPYxZugi7G2C9h
VgV8ygHo5fa5fd2+eU563l/NE+FRSo4wmlYCWWfUJNah2Ep9p2mglM4uip7pkFqSgyyJWzgqlAbk
4LzgLAEVGvU2oexdjLiqxHrqGdAUUMsau3lxT9Fs6DW6qnmSFnNhiwll4Drm334PEfLOUgXZB/Lo
LPkYkJc31lxYHEe/GmXACgQxBWixE6sFsvLevuir4+JCP/GkDL75Le87n1gz422GLpiRbX6G8eiG
8HVUiisybBElCskd4MyCc90n9neR4co4lUjhKSquEltsGZ16nOls+pft7RTGLEr1RpZKnsc6EcAc
j38W7EdNvAoAXTAgvSMT67uv33m9OP/tqNlzPFD0yVj10rN2YmElIQipGdv2GB4u0RZt/uuWDCOi
g6uEse1vYkKTYu1ve5dTAJD7THhPO948ooEGOoEEJ8sAgvRQO4uaaXpc8y2ABOCkDJ2dO77f3Mrq
/AhgVxN3/8mFcfCygadNsMAvpZxwSvWndaBTQez+C8mgA3IYjhitVU0lm3KwOZ15EyoWAQLOqlvA
qAUW+SExabprF4kYanG9PkJOmEKt47cw0ARSDUbNUjwXkG1HAWDK1ZIx21lk5zZk9LWLuoERSLty
NhVrX0Nlo8f6ZFgBSn8c0BBrB/nc9NEM6AT1dImUYQDUPuz23iIoYx7aahlRxQ8zUabsf8XnmeZk
SCYDP4zlyyDjIEz7lMQdzlaIhz0n5waOd5P/uMHC45MJf2GmkbdLZZkGNs4XPqbG1JCcvnq78OKY
bfCeS326vf3aDFesvrmGuybEGPjtH0wgVp37iMZ0a8keLFEWBZcG1Svt00VlEx34oL8S7DEW5NuC
+sHK/g/win+7QDTUnTx3lSyb5gaOhPk/2pnIDg5zpKmlNos+sCQlQaMgwEDl65XeTe42JXhzTCrl
//r1HzKFjgYg8PwLSUa3hnLeRsbFKOumiQnD76MeqSjBSp/JsehM83+rBkoidemMXMqwtA2uJjSo
i0d/kiwtwVRZn+YNBHqXDifr8LVJ0GCh+nRGD0WKQErQOp0NS76gSRC5GyfzjVr4jWbFYQqu6Zo8
bHotYsgimuFB/77XRbzafAp4W8RPYO/KZbkqCgcFAdXl2RIbTMa0Ht0O83yXEAxhOoFbquBJbXH0
xktXlbjUm3gn0+doaIJim1KSgwCIRmkLn9eXQ+k4FYDFbU4TIHRAbkUO5spNfSeOxNDYmmTiNE8a
3AKZs8oxCdM2golYw0/Xjpgg2J7gPhX9jKqeguOkZNEcelFHYpaAEMXqB+zZIjOxEzKPFM7sjKxz
qASceyjrXbB5nL3tmVPl3+brGoB81JsGKEDISmlTm2dsHoXP/8wjEVNPQslEw37NoqJIyQw0b5Jd
BZJiMlbfxtEC/ysxVoIVrGyrlqQ6Qt0ibqOoRuZrNfk8WR1YviBw6v4MwYuZAAgRyQyG8fSMN4Fs
MbfS2EAwcln11nHXbuJzHnYfYILuBmb/hC+nbUnOIpbDnoqcd9rkP0eV1mcSYo/mYobkr3P6dxMx
tm/kojbrqkJ2Crpl1Ve35zJmZMscP0GNDNjTWRJpM4UI3k5mKrntMONvLpdchg+v0RzypOWv+F7p
yxI45V6rQvd9EJ8+NmKjaGKTNpDkmI/y1aJxgMzDaSUI1kIwd9YE1KVa1QWqI+DGgJxYzVSyjFGf
bMfLcs+CAtMtoxr0O6XfmPRvhBK07EMLV3huHmdQYMgclCyxYz9etb6nRcG8cUfsiNptALWJnwaH
BfFEUCALweEKogf6kxyQYIsOs14G9v6ep63ayewWx30nI5AuvAY1loODqgORTSuxAhu5CM98BvQ9
2gI24KMQNxaCuKDInce83y7zgBxLSThIU6Yt5D7OdoWS7pMMWWTwwM4xPe9BiR4SENrCPFjbesiK
6rRTe/FS4DPk24+WH4CjdoARohCSVWfcfw6QnGOzntyjIQivvwQ6W8DYqQcvpwEi1MxlNkFPdGKv
8kIWRMDBNaEABMWQh09T3afnwl1yrdB0EXrcW4HE/qfZqPqY+961D4qCMzEmnTi4smmw7Q4E2xM6
8tmGv/Z3pWlIH5ZGBcJWGyx2ak+cxPk8L7RXYjbdxPDeHhWOY/Ly1Ud6cwpTgN5XHurtq92xzAKo
LcfrCIu9HRxwhKv6UvwU99jrvE9In2JlZrLqwvRHA0Gif43SbNa8qCIyparH1xQcdgvZgSm/Hev0
QrzaQAD8MC5koN7+LjqI9/3vAPxxseh34qkPsScw3USDYVxV0KvO3im0t5IYsPHhzK9bUGB7FjA0
J5nfCing4OxxO/ZoI0cZHNSBkOv65K0VTpSoPrdpKtyEH3Hp1KzwP1fcWUxxfUkjVt7rztHjPG4M
3TWYjxfR03VW2gQ7HustN701xdxXoHzoM++T8/NWGx9JZqNctg+Ccj+50sst6EeWb/+VGwU+xo3g
2N8FMlOwEy2sf0GCySBEWB1BZe/ZH4X/gY+Pepbqy/fPtNrov0cXA+aJszS3Pq5B2l6xwB+eHrUB
mA3pA2lFtZIaHvOKOb6mk/+owCpCgobKAdai2E8K8yn3FDt4hwvjQsxmN0lLYdcOLgoeawa4+gqJ
o8ef4E7EjgKSXKG7rzdxPM+Elyvi+xO3ttPfXYJq9WSE2v1B3iMviALCdtDOO3VAi5/Nv5WAHr74
WD9+Okk4WbWgOXoe2/7Kdo0eTPeHZi/kXRHy1kTl+8DKCJbtEI47h7uwqvZtUXLj5iS9mZS6LMRj
rTzXZcgfbmABoY034W9Q/aEX93Emv/fAFtrGMvZfVyreRVrE1hpGIW7wHC/5sxtPLSe8lKT8oxjA
5BvZTODP5cCws3ugdJULmfOf/RzBsrAdm5Ey2qP2PnFRnfmsdVFXgbmdq3O1a19CnP83TCu6JYLA
nWT7sWkrRA7kZFD5+7100KuQljmx/bV0LbTfXI8K0F7YtwN9yFxW000Sdt58lbwlNrTsvnIcCWmm
1RzWkvF38xdujfdbX4d4YF8baSUwEmi9YeviDKCJd6zXHIk7mcvupcBXej6CYvh8yLy2WCbNiOzd
HBFXMX7C+q5bTlQrMdt9k3Zdyrs/EfBUrwAsoOajhgZdt4n2S75pv1T1GrojPtKgRe/ti5LKjMkQ
p9WpwLg0u9tyBkSEQNp1MrP7avHpqsC5No+fgnDJCIMnskojCPr6wcvxg82y8kLdsntjt6HJEFzq
8oJAQ09teTb/YU8zueKeNvVAabhptJayauKjdF2tP8RO5ai7GqVUoqO3CfhDtDwee+hIrCuSjN/N
amaO172AKPI2/ndrTt9XsfoKIJ2P04CXqse++dVT4adHAAqgV/xFdMr0tunmQq7u2zhm2ZZ3Izdv
71P5xQPjtFH1JL0nE8/nuCenLjuD6e4Xr1QMNlXp3648AWfMirGGarK7CUJdi3Ou+WQ/EMTbnv51
4Z8cMnoYWh4CHY/zJ5/3CPtd9HDKqN+F12V3uISZtbOr9yQLq0v3lqcdKRmcKpCFjPR7MqMXSeDy
holHH6mU236o7RvEwiSsStxrVA7tTwoH5hh3nnRrSrHyb38z0YczPv5yV59nrwvU9B2hFBUfQgsh
tio0W5+3hXAydQ8ctL2YDh9JBDptrxNgvVn24bN9Abo/I13GcX0+od85IXJejiUawU1vb5z25sfO
Lm0BT805DHZ3m15HquBF7Y2LIwtGBCdsR0HYiu92XfFtARMHYVVJCrfdaUXidFQ9eR1rwonDCRae
nR3f6IljO90C/B86yKuzP6oBjfBLKFD+DViP+Wa/OdYDsw1QAq1XulBQ9/duQPo3fTAje5aj7eXj
v1PwBqliu86G18CwjuMTWlpae/iS7geNI3zXqjcV9G/0PcZ/cSxW6fQciE+Urjpy0VLddZuJLdT5
Xif2lIe5Ddp+4WOTexvFkCf32r4Sck+4Zeg+PrTGPneBRZvOR6Lh9/KdzsI0MSY+wGBIUu95jhox
J1wicWgYqnwLjleIyBPjCQlROCdOGS+vf97hy5/sWmmszaqaSWl9QjuQxRkggVL9AYvrma5RrEM4
GajWcYRQBvyXbLh4LHvpf6UlUa5UWdu1ieW9zkMgtJwuGsoVXON2OBLdmOGF7vfUaaCkpbBYO+7j
egyTInjqrepjk9tnj2inNGNhpVO6EufvPgGpqogmhN6lkMuLbaiqYrpIdXpdL/gvmITbjcFmOng9
p6zRpYlq+wIr0nakGLJNWG9kSa+coqSU9QTTiOlTpIp21A+15rOvKrCTn7DaeEueEtvHiVm05Fd3
dfU83mY/TG4uiXyHxpo5C23tGuttEyzQm2dEVmOpK0ykY6DpBUwnEaa/eSTVdmCcVhbCltZvMVj7
/enUnm3NBaalLVm29iugqkLY7f5XLn9cCwnpY8XXBbhOB8oAciQAYFuIvWHSp+EgqZhzR0IsEEdt
Ib4BKqrRLVnOPfaNMkuuIluqrqTNuigZ8eO/ea86nlTelcbIYQDePdsebjFMIlcwhQYZok4p5bmi
uXkmE8CWaGSGJEVJVjZV0DGk9fj8SLnHbOUDSZt608SttRoS6T7dqGJFxsdGF1cZBRQOb5YDId5B
KurInIZFldXSjtRyxXyMRD42wTWnSlX47JzyZf0ukmhUUtrbAmFMOFzcazuh0EBW3WGQiUVtc12y
WFtmZzLmtiLzVSNB3fxiUTzAqoqWkQ5CDmA39ijHs7/WsJkqujrngBJyDwMQKY+7GrZEzg49igGb
WIIBWyg82QG5Cu80APnA1CbXMD6xfzA72O0doXLeZRlx0Hw2pzqU5BwzF2gNJIbh9MYfkzhri2vs
L/j8GPpjNdkXBoKvbZTwt3ckf1o0GATdNLoXL2uA1G+0Tl9sNNggW0PgDN3V0YGiI7HOuGIQBUZE
6KV+2AFPqTxeZ9s7KDnZyG5jr6K3eCIqOq4XJxMCXYJEs3ByoxSKh8DQgBH9LZpirCtA4FiFONqg
RyM+3RmPpRIWYVy5ArFwnvqbhxARhUeSLYDG3lLmvS8bMXzdNsgK1H8SKy1+qtzh9s1HXtLf+6hc
AcJZ1aW2VomquZIk+Nzizl96t1ka6rndrLO9KpSJdkC5XMtvqpWi7jGV0Sbq0D4BakQ6kWFENBIr
y9MxTVbm1yDfqPQl/RipW/EdsMngshTiT5SiukBPQj+FVXJmMImf9r0A1/WcEx2Fw9m3uSaBoU8x
Bz83MBVsUwk/GLXZh8qk33WjaCsT1pxfUuyQ96NN/3UivUo8WDt73uc89FeMLoGCOugvaPokfkrL
GIDnvJvGpeoiUC0TUcrwCpiNG24hFNsFQLUFHlBYBbJ51HsW4JSc9urzc6juVyCiJBZs/ml5ki3C
fXop5iebs0fbvKHtdqjST38xBFGEzMPkzjN5u2H+i2JGreg+/pJY1P6bTaUKqwh/Z8UVcPjFSav4
GqurXtKf9QXvO19fuMcOQTqZ2mdBDFuUDpmFoWHhWR91bb9hiPTmzCO5OoXGAZFuCSzuelNA6XmS
tyTQZ3OrowXYb+5Vjr+hGnVYbQeB8bv4xX72U/mfJglh5CYXJYAtl57uwHXNPEJJqyQFZ9ZN99IP
8ghiJa0LrIYdtN2g+yM1Fs9bGegmHXDgxYy2AfND3whpglsCM1zswgbvLOhBiXDk82RgLhzprLN2
Ngyp0ZEk2UYtnaFFr1QPEfwXNRwbbqlaCTY/i+tvzpp7jr6v0Jn2KiHmUFBKSxZyt41LN6DPlDiC
8bcqo0tdmpqFX0O5rrtqmWWMTDznXLf3IEQfuMQXcOoYCmTC+0sse34jE/NaBzgK4F7TH/HLvYoQ
SgVxSw5JfaV6x4eMpCB8Qn3oQ9SvgZODGXfy+fkDsuvsNC6wWkf6LEz/cgiIL1zBCb1rWdE2rAtC
8QKzIb+al3wEKVM+MiDgb0XOiQcm2LHUmAbdwixwS+keNeSbao9XaWBC9Onrywp7A5eDg2gOBVCX
8P7Zi7/L3MZf3eqLs00kH4Q4BjxA9We+rFrwfF+iFyJPsoCgQXCwvufyn1t9AF3l6NqpdjBtkPcn
OqXg9RTpSN8ttJjgf3j3WFwEBp6bG40XzN6e9WB4Zdstb1JcMkuhqoD5fsD1XhSC2hvvaj1TxoyJ
H/TKJIOK2pGeM9Rod8ix3lE532GDZlaT46vWqZ9muT1hY9viumW1rziJI+1rr4RePmM2wkWvZlhp
LlwuwTkHXWALYitZOOJjnBqz3zFud/Z8ukLuW0xpxiNR5i947eMLMDkcMnx3efYglwoTLRbGkvDD
cpuhpjtZsyL5oadV9huEDKQdqXVYwuu6ZKaF+P3t1AifYAGe72B6QbeH0Go32aKO9kdmWXBTd2s9
n3Aaw0VQdg1sM4fGgg+tZDRIYkDtY+W9fX8IHeiIpKDe8f2zQ25xE76InXxXKOdsxhjOYrZYl6Ce
KHYUlhAnoHxX7l8tB5ll5sNnRroit0/eACNNYucLR5g1xEbnVIQfWeNqPJlXMpm7jLavGLFxHmit
ZdiJpMF72QT/qBrsCh/NhGGrmmGUJVg3zkBcIMswu3n4uKYMlbZ8LTbloQ+MU8ygAr2Ne+IA4wn8
XSkMUzvtAyEKwSAVOe0LH5ymBAQ/dcxJbOkQpMfbSlcJt/I5eZf8SqKCOIIvmRgVKQOkdIvWcrtd
4cE5JmF4VBNPT6QDuTmWBMyQacWyePo8z8R5KW7fgrT1b4ySOb2WDeREuCCqYOpDvoGtPXqFdMXX
Ehp4i8os11fnE9FZCqRHgyz7KzriMhYv3IiibR5Ty3bvP+WTOBldEPT7rQNtNkGY/7nkeRJr7GeB
WU9YOkm2NZM3h1dykERLHynMU6lSUFsP6wdZNCEHyPDcXa9m8tg9xF1HCvbMzQYvwGKaK1VaqPg9
hj+g5eyuwNaMlBKmrDYR0TW7PN5Hls51IUGAxK2W8kl1fwiY+bCPi/CR2vkD75RaZCo/R0ius5wP
STzyjZpIbFVaIkDXPAN3/T6RKlpfBtVS/1YXfQ59phdgOS0rwV4csMXId5bHLun/5pSNEttHPeox
MBlS76WXHlChgPhoj6igl9q0EuNd1+f7Iydhh6A5jKjeU4zKsyxCXz2XgeUZ5AIVyKOl8D93U/OU
oX7VqY2vLmediuILhQ8MUEsryQGF9WpW9GlAWhf2Q3FZ65eW6/6EStq+9RSiMOVHjvwh4TXk3f16
ILwRoiUmtISTU2vUUgInULhRua7C4lb25wyetBQ6PT5zZ7TrJVUde2NQvQ7h9TbeXbv0jHnN/7wF
RKtqzAFiPl0aomEqJSo4TYsGX6QMQqr2ivAyMnVXkmsOq8tzP9oRQWHhPWeKue2LJmaXfjPpZ1sj
mCQuSX6pScWpw6pe6CTFu4tH5AmJaSKjz2g/EhDwN33YIpD99DCCi7ndFBartq30RJPR7ZmmBEnM
JexK+ytIMeFUH34N7LORDC8d9ADo2eBk86/uvBVU9DE4w7dRJTjLzNxzaOlFuBbTa7rmRDOdNZvL
G1zw3cZFhWtntD+7KjBozDSh2bKZgBAfKLOcV5lNm9t+VsIaXt1LB2szHcvw+bpnwUbskzvvyzgh
hUMSv4UKrHL7vkQHIt1emFmR6SXXqQZDPkspXIjboZaw75ryb5yotbuLCAhQdw08p/MEQjnFkgRU
144Y2xP5O/ZGBTtXK8UHD4SFT5g5LQ4losBHezYv/xFMdPUT4mIm809+V62CjE/85ZX9viv0fF84
DvMfpTQrHjjmsE/hE4QcMZBFIybVKu+zeMqIpw+U5FKACXtGATpe4Bot3orKxBkpF+rYfj3tgLUa
bHKYyTx9ZQ7LEKtEOmgEq4+j6xvi7ByvBftoDeY5rHjm5xQs2QmtwGDV3eauU0mHpB+lJYj+m39M
kHyCbtvOsK6LL1qt7gPVqByZhuYFOrh9PW+pctUIEAEMzvQSTZOKG3dIjTy4HBkK2heJf062SlDN
rktKe5EDfpWgOTavFmbGYG57kxyISNLRKqKp6WNZrWMzPvjGf04xQqluuhMjkt/KBbL518KeJfBo
Ha8SILpUr8426wIHrZbzvSzRvnjTRDTccWpRGMWnsw9Tp8wakdp7NBXuSj7J1szh9OmY0do2gQqz
kFV94Wsfw9CJSKEmM0p7oWBdrT3b6bPWeMixYzk3HGreuVBzWQOY29Vgf/qYWbznzzPyHaxl0sH1
HZ8d6I1tKNUtxWKYW3YVlphryqbjWhhx5Qstksjww4pQgbI/k69YvENMGenqjhSX8uRYQpX29Xip
d+ikjnNawihwtz1eG4mdT0BLHLjBNf1FEJnlYrq8Z7QfarWdAmaYx432fe+Ji65kXUmf/fkXSsRv
zzvaYOKqeZwlWW7sGfpa2cz3/f/HlvOKJT5dpPzJ488blDg/qwzuUGhiYV2GgAxPNJ1ugmE6fpDK
wc0djQznOysV/Y2Dc/PGtaDNfc5aKEctvbNLWTklf+bZJBNgQMAPFFsSujvIdr5CxrHXejtQThwo
bo3Ci14vMvbHAoSKSKYzq9zGIbY16T+xYkGdj7BgIvS6ZStjummIyep+CpgatoLnrVW7S2NCSJHG
rjtA6B1R8rJDKJxm8+kg0gl8t+Gbo1rh07zooXvO/i3cqDg8J4p8b7xcqnYthok9rT30+JCpZ2p7
v42lm9irDb6UnQKVUrAQS58MlvhnGWqpNlUGcM0sJftA1D6rlqCn6sVOHWjBBNEGiRLJpSw70mi4
DnKV3Oa5xuUMVBdFpyHloGBUN8sj4PBr/zPH9wbyF7XSSAQapEs62gda9i0eCS/ItQp5KIa6XGxg
e1mxbty40kjlt4nVpT1RPL7oYPmaK4wCepEkg5t7Cbl5K2xgYn1oIsAZchyLbnjuRT78cnwwuOHv
6o9t/+KcKlVrtC7nP2LUHi2L6jalbavdXoWeYTcR2aIwVnfnBeR/JCUHNGX6ovd8s+3iXXnSbhab
xk7BDoEYE62bjjBxrKf2uahCRtkHDgUDLA04Yj0lHziLnyKxpU3oN5cl1rOFx4E9ZJoBIOgw/92O
bHT+PGOhsNoEOikN+MhNVtYyUWD41Tglp2guR/zj3PdTFhPnvCs6R8n1ZE6mFxO60PWrgjLAf7ry
nkqaTew9JICwz5prcDGXH8T+K0Ok9NDkanFk/w5tI32gp8DM/t6Z0PCcHZU4yuslyYIyZG2OVONR
zg4IDUhxkfg/uRZRuKIQx+P8FFH8epW513BnNCYhfiF7owIUgyTu4VqSUG6MVNhtafR08A+ZWnEv
HA3Wg+qeswBKpR8yGbcvsw9MQLvH0dli6dddVALTDLgPxo6Iz7DplrcB3QuOqSXPol3Po8jfGNe4
6PGRUGxTf9kHld0Zt5Oaogk4flVKPewjez8JPc3bxc5XgfWVhV5yQXZrvxU25BjDKyn+kyguMUSk
WFOTXjlvRr1pPy4Z+CZuCHmA52Z4c2hkFLHmrFc7qkWeDKycxkYjXHn0NFsiqcuph8Bfcz2q+8XG
L+L43CTOes2DrMiKgnkmqZtbUX3Of2OcSxIhU/eyZtPGtJ89TRb5kaO3ToOxYMEApu3UdqM0iEUy
9uhB15qYOaUvLlNGSpyZy3hPG7s9G09brYGG1cv/cGyyDRYsNzL1AYunWR2Demfr+HYRZj4CA5pj
gk/0DqW4wnFLz91Es2euA1+Rko9qU99etPASen0PJ0IjfmBgm5vLMRi50l+QNY7QrMlK7MCFfTid
FW2glDXRG+3c5Xs0fL+l31co57a8r0aiH1oDzQDnStna2I+8oia2VtxINRjaCuzzN1I6fKap4h9M
VWmi3yZJOAe/dlwHsQEKg2Z3xN0aozFJLU7S2ei2EauZLkQG0i1nQGN038LQb4C6J9+QSeKIHi8/
GULjKI/u16RLaEZv1ssCpZN8XhsjzA+HdMW7/3V9fVzNYVeyb08nBw1QjLuKnoiEhmZO/PgXZ1+X
R3pRwwvK0sNSQozrwUpFa2n/tIgrPH8WMTeZLgn8zESGR+F6OLvGiBp7YsLcmbVlz55UKKIvGHkc
AOFMbcuX5+bELh6BFITOKW1Nb7Leu655tO7rAwTYVfa/XmIEnGhnzeBamtWD1CSnocmnNMvT8cPF
mwyX5MMjbKg79KCOCtUBZUmonxieEZWlJoI39GdcGf3IM8y0jS/uL8d1Zy5WmpTVUNs4aT+JiCXd
nUZtjRjrx1brzzr8X7CAk45OruXn36O+mPV3vdRdkoT+JrgkWO+bEBqB6ipxrjrEgjt+dNIzyd4b
1gkTjo6V4gTLesGwxRJ8HjAh3E843A+gG6kmY/ARdlHTaFykDSTdtHn9s0fE2VF5w98/Mdx91BaO
UumjU66Iso6y+V9MvHHU/rgbdeNtRQb8UcU9SP7B40akapu312dS3xAdHlVD+pePEueBZflCxvnn
EM+BrcMgG7C4z6JBahgcpJTZ8C65c7282H9+esxcoTajg3dtcrbaUvvKz0FYtgoUiOt9whBa98pL
B0imd1hYX+q7N+/6RQNFYgljqPNrxC6deT3K86G/81t2uy9PKElAraHIE89+A1chpAJtgiAx4eAY
YP0WjbuIO8kqwKZ1yZy6LPqIKtGfvhVudLZok+S9LQKPYZuKsJCJfGgApvMT7gpgwxWpW3KyuPjK
d+C7hqx00om8AKtZd8I2ctAy5hwYga0nvNQFD0k35GHwQMCiKG3GN+S+d+ZPzfSJ9OYXhH+gN15M
NDDXvx0Mhw8hxN1wLFlgYCb+BjdFHMxV/gh27KILUcAWLt66v0+/HGmy1bHf/TKKhYtUPLsCzkIq
aHm3lN6NAYeH1RQPfsSFuaFKC2ycr0OGYg6pjzPhR1WDROZPSiIMgIX8F8LltZK0HQgaMFo3UrTt
LtIbul6hQf8DSfA1kTSFsuWBtc2GUBU40HPFb+Qqbxcsv6V1Ne+wuW4gzCwBmaQqCUBDpmgKoBaP
6yUhhToUuRVnr8qvndJHl07SI7gqvDU6LpqTi1UED57ysOvTSdiSXuBYuqyYC6Bih2IDQaEuRVpd
jmn4kjdWZ4qqcmzKdSuX9sOin0+KNZ+r/94C8t+bz0Z+UycwdguR304vsXvM/IYO4aniLd3m+MBA
9Ir0LsAh9gDB6hY+VguuT+4YZZwOC7nvWWBFuk1XCUxg2NmAwIswCmJ9DQnPuj4OS+/Wd19vO2cT
3D9s7f20Fs7iDgPwaFsbZsu3M/YaMctK16FpyyP1Ln0btMLnngq+BSBhR/3P0GIVacB27ldW9Acd
T3j7TuG2g0bY1MP2WP221EDoRtqCxrGn0sZ7cOeWo0rGEBXoJ4C+nWGh+wBiDFXGhfV36piYCQ5Y
32PZPizQzCf9ZywrfWGMUzVUAf4O5v1Mi4a/zjHsA9UTJDWgjqh7qJXLqOEFNPz2gnpNc597eg1u
V7mGwXWlqwvHUrFsBEhDuZczMTrzKThWfo3ODqeLTYLFw+ik/V9BJ3N6Z1AMSJZxmXDyOknSEEMJ
H09nihykd2SSfmCrQt0HfP8e2S66nrLIax7/DlDc7mNhBz/56OAgvKZKq1RZRVb4cMw1MFKin/QW
y19Oos+WZ8T0Lb9LhYUJd8fmfgwy++EJ0KcVVjjDUuaNemmOQNdJCboRU2OBHNz7PPRKfWEdXx2h
lflpNsnDILJv73C/LtagQPmMki4VEL6C4Sd6VG2yavyjhmLaX9W6eb0VIAwZcY1118TN4Ve/EL/B
9ltIbkdyLqa1KDbK4i9EcSPvmHB/6b8BHpdgqlXi6l9UG/Fk0seOxxJQHjQEdY8xEXoyRb3jrFjR
ZkGOsfn0thDcQa6dMMWGN79OwXZRRBecJfNaCuuETq8oPH1B257mCrh/ezbQyLYbV3s0A6S7eKQj
HaizCu3BmZ8O+ThUI+iwNV5dxb6o38GRnPjGrh/17mH56oAncibj6qkFUEejq3b3hvjpwzeBSOKt
ELTox+do8EuDbQe+Whpi0q7ctkIeY4H8SP52B/ZNkuHXoUhEa1y6pYSz/QoDOjdLJKQPmh2EzOd+
diRj8UNsQGVITAP4U/mICuAKOxuonBu5Hs7ZjRukfP2rtk2L4SqjEAQ9HuldChKn4OUMeUl0Ql1s
O3fKTqC/OE6Mwfb3PmpB8xvcrZ3EGnEZvUOG3t41ndM4bQE+yBh+gGytZCjqjsgwDi78zN+LEwCZ
BPfmIC6Qrl+V+Fyf28RMOkm9173uj9ifdz86ygYm4b5KdvwsTLHgQt3guU9fDqR1+wGN2307Ixro
0s6tGeDhcmWDy3Qd6h7+6RubWmLYmvKozhK9My9ziMAoFrxuWxA6RBoQ+g6lSqhWjOSDVaHhjbAq
SC7dhipklB1V7gJLz6iQd2qRuE+6TEONhMyFdpurmnorH18NXF2mVJrWnvpdhkaPQn16DTKU3kv2
2Cn8zomZJZtxU5uI47815uEwsKWwZBCYuPAyMssn37sd70hj8t73wO9XQgY9PczPz3iaPzpsYpJi
szlbmAoKsq+M6/c9hxiEe9SG5zDo4J2DuPHDz7HBbo0HR9ctn46XApnDqXGJ+JajoS/RuOmaOkoe
G+pVq3vhfoTb1ygsg4CBYw/cmQS4O4iNZAis8/PcX2RPCcC9/YqEzzfg6p/mbN6IX6RV30QeFaK/
Q5zqJOXiv7GnS+6taDXw/6AByCZfndzhNMzDKVEWZagm1089WkfmrRAJqCm89HT3j/S2KYZ0YM5a
qIEFKlWBs+yicpAAryBsmOLL8skBRDKZbUkcql1+YXxlxNfh8/4kUSrnH3CDFfUX1FRhY0+hlcV7
EN5HYbWN6hss4sbHgjU+88ICls/ytIaYyDF6Sml6Xlxc/RDYUvmgEZFpXzTJzVMsyThzZhDrz8k1
gXisY4/zckAvNTRTOniIgYAlacV5F3olWdyMgipkh05qwcKSEbhGkT6raUbYRWp3cpgb544U7cqm
rmr85aWRGrVJPlpULTtFFLsdbjMCF0w2PeMqkAnXJhs2XnO4TutSkAt+HFN08/NaeVaFcICChSsF
n1/ZNkenfcKUlhz2PuW4kj24gDrUSo997GKMA6d2yG2AH8xlYaAlU9tL6YkSQ5Z4DhWBywXx9tgu
J4CteYayijmbiIc3U4K8s47JPSJcXAkoZUuXSf0tQ/jnmh0rfDxw0sJKHA2Nl5nOzK1duC391o2B
ryf4h5TuRsIyNhzfGA34uQwb49xeUZ30+hpLBtcIZkaMOZIRV5ossGi5I0/dUGEQNh2CYLWGzVnr
WZk9zChgK9xhaY3sF/Az0A5GzL9r1mgRds3avTHo3Rw8AyFMd34t8eZDD4bHRezDV+JHhn8WfIHZ
y4v35RbAFQqXKyDmlXTVRd0oeYmpgcIhJOCTEEFGWyIkaoPzhS1+KcBmt325nyUgs19Sjr/zSHBn
YFQmT04RPC7leNxmhr2kZ9Hc37tFI537GKkKC1YfzAIxbnmSVsr2ZL+nFczjjWN9/PGOKhRt9CnI
CeZ5XCh/nUGj/kzRPAEKrdlbPVngCB/AGrEbVf/bKcO252ZM2951aMszafG4r3sVAd3QnKV6ZSiN
OjAPdE+NeY/PVFOZsAV9/AzlTx5Mh+S9Gq1HpDzIx1HdlgtOqLWP22mBtwjg707OodXmy7fk65jn
WZCBzbB0SaPl2Kir5e7uoTpq2tc+Q0zN5he498pIkACzZrFJwqoG6vNYkPaZdMQAIaJbqVDv7ehy
7nLENeelCqbZ1tUN83PrSZlQOyQxNyja62lYAlFXdEPsvvrJZnKBC1FVk22degQv3fuvKfFMb4fL
C0KBF1dZG1imPqaUReW0XYhSCETBTbflaRvRO+2EidgvJjOFSjzZS5zN6Gzk7tOv5xfeVsx2i03q
235s3ead6VgReEG4kOWrFL88dHGXPL55piAbHlPJ5QZ0DEzVKNU/4JEcKW8W/AtO9bbvJAl2yQzq
Ppwurud8oeVtamwalR4VEp3AG0eYJ/IQ2dxFJMXYj3GIV7/JCGImHxdE1tjuryFCuejB4Iy9f0OW
jtdVsc/G0d8Q/arKPhyXk0H2VFqM6wVQgMwZbs0YAY5RMyWzlzqGb6uBainAzYTuIdy2ZbPtxmRX
r+BAraIL0edlz+1Dyo3PVULkCtBn/NAZMfPFEKqyT/H5CoZosSSms6XY12Vgvc3zlaFOBg0oiMvN
GryzCin4GXUApPelPWRq/NsqI4HADzLOKUIRponld3ZZn9kpupDOJ7r6hqq7r2rhVaAYkYy0sRPc
+zgsSzCcTLV/RNtodbHPIaxwfMyxoelWaICwlxzj/EUvAaBig1cMUtob1V+vb4CaTr5f3EqxFmG8
YRyHuZM9vvXDgbKKDV8Vbhzlix6rDp2zhxbRGoZ9sUjPDn81kKquRZEkwAoT+yjOuisVM0v7ALKt
2KEloU6YjUdPSiw4esWiNqoZ1HXyWSCNj4Dwd3exLflmr5NfUb6+fq4IUxTQSx+b9Nl67ysI5tq9
Ai4a3XbUeyb5NAKs1WA6wDinP/21MveI9rwf4sOPKDoEU9iG75DWkOijk2G0tQisxTfG/c5lkV4z
8+nshWD56fx5XrxW/XRWkUUxkFbY/rZsM4vlN1zZ4wWXQlgPmXiZIVI+4hRCK4PCtkj9TLucJfvX
uUbG8c5pTKZW38vfKLVZ5+zFcByl3IsTxux7JUWp4a9LlNILnZ8qkdhJlnIsWmkGksf6RzX2M4xv
2Cj7sp3Rm9ruUc7VnOLq/OTkRMprUvN//+7fo02o+UURWDJn8U+yC3zRnk7PZiroxyTjcaFAeKIj
LTppNTs34uX27Pn+N8bwnl7CeckH2ZyZaaXl0gIH3NqQIca/S6d+rmY4mFmQd9s2ZYjzUr1kb3ov
M5ot/oKlMoAqWbL+vKw6Eoa42yXwTOlBkAvX6t/ycRoAIlqJycZnZYPcGiu80rtUc5iGfVW2DqJt
mhoZyUf4gyoIPwY9+vvpcEcV6HmS/PsvtXwvkqzZ6Mgsh22tiu9C8YKGc6xf0gYd/IeoSYQodGcs
CrkQsmXsP6OlckWJuJ+SaZ/5pYLnQCkml1+9tv4mly+XRSMDKYcT+SzfUA+pdfbJybS1YanatJam
KjH33PHvg2QfDCfHGIbX7Dc3BGWLTWoR9p/fHy6RK66xl6qx9zHHwMixCdUPDeWgnrMDte/8wSeZ
lbV1f6FHD+LDb4oPsv0MtY1BGqdwf3jI9Vzh2apoqfLJGV7FzwZnK+xbFQi7eKMvRgy3S8UuxnHg
nyPJjJbw+oNnjk+ywVQ4rzaNDjYrxkMu29UdR7HLP3A2+egchlGXrGGpVIwAki+4b1OgQBa8Z1dy
N1o254LFz/96Iwfn4f69uAuSciEqRwARKuosgOwxoQpG+W6uJEtBZKj8uBKDeEX24tlMDR5fxzVI
ORWHrGFSq7dz+3snMTsexckQaGOwuSqNv4GM8t3V6OqbFnhzCFebHTseoBWq0Shpz4lmJMFKWPLm
WBkIngxhb0Qg8RgkJcr3jTaLaSFXLZJMg8qVJhAqU7ZFBqMJGscRF6GcjXMWVi4hembNXuCuMKAc
xP0D6dX0Bw7tChFj/N7q7YV9X+3tAcI73wUcpNMUOrddcqTwVJ8npT/GhXnyOz2U48LKra4r+l8N
gTTbxDYcGU3YU+DbM56fNFEw/uc7DEqbTdRZ0s5JNItg+8cY0xIPIHi1z+1bg7hkBGgGO1CTlqnY
jr2Cw+4uQKmjXeK+Vd5GLkQEUFLjzqXmVeGpYixUQnz/NKI6cGvxfwpv0Flve/QFHM+UvWwVtkv+
yEq0aNFCoinLEm0BeauVbbcliigUngSnvLGwAv4OwoZNW5gmfSqkS2D1ij3BS6HvnIHbiasayDGp
N3V1lRfXwFAYKPoH987Tlfc+WUMuYjMZ8qOHpYFYOVzoz+FyK5FSvdT7OVLx6LXGwEWsvreumtMp
Erb0EZ1RyD+Q+CE8MJpvdZiz0x3/maJbi6kBso4IrL3fPu3wyKhYUrrX+uabD2uScm39VGhbY8UV
XxnCymKwObDTSnFku2KWLMxLBxdMRdZTuwyZ41eWysH1v3OJrYt7M8JV/8t8fyoJvwIptmLOaniG
BjoVye44jC1aEnDKK5S4wSgK4YChrcX/Plnnq/aJc73ykKfRy2Corfg2YG2JT+Pst0Jm0nPV280p
eYMCwwje1NLvCj9UucSk2Zff2UKczBrwthX6T47bWfvUDpkC3ybgj+GTKztMFAsPiHHOafVJrCQv
mveepPqD0Lr3/26SW+9QNpeZoQ/7NicfU1GKT0nTZRB9b5Dkl2uJvPw2b1HNGR/IZWOSWbBAwQPQ
R6sxwVLUIb7sbO9d3tDXkHX6FRYWytey11CREwj3y3GIanHDR07gu8L/ycM1gefYqKnhglyxq8Xt
38E/K3DAmbu+TcYIu18DIQoCToJ9MWYXu859+9ergX3Hr7q+nqvTuDE9IpJkV4Y0Nmp4HTmiHlKT
EphVPzUhzg9yZVutP8QFw34kQxfbqaXPyhBtQdOCAFazWi8WuwByS0S+fGOiilKuMrkHPJkMGL8Q
y84ShUMZBAquI61+k4fc7hhIKw6zF/ydswMWa0tU01sH9aNc2iVPrErZZQe6fJmYAmXyHrSkaf6s
nsTXycci32kfDeAIomCansPAHjII8ioq1mQ3V+3ZZES1j3kbXEbG92wXAfB4rkPWI8p/5XrfTa35
fTu03DefWilpiuzhRx9s/mtQcsA+Gkc9kpILCvvyuJZ2LWcXYFPNAGOGv/epWamv90SPDbrMlblB
KKgW1+hQf3zlFYkM0/2HV6VjIw2ydwsOJd+LqBQrsNiOpaYTG5t1l5FYgcBXFKPmhawLIHPNZu44
iGtlOfDcdxAP6/eZbub8kcJKXK0Dztlik8yFAikcer1sP1iW27Q4n792K56moKzNLFJx9RAyAt2K
ECwE4+owGPcNE7m4GlxP4d8eyvMT8KmovTczjcP3eWQcUEVmY7zH5mL6/CMhkBLtqHAdKhgoeUzN
NbkUSM35yrXBsTRGLuVtm9UXh1kxbelos0zJEPQ0CAc5fjNYO7OxT3WtmiI/29rSz7ulFwek6cTZ
MgrBe6XfEw0YItk1+wfFrT9hwIZHBhnseb5TTcep365r2CXla0q7OqlO3GPN4RNPUr43PXugSbdM
SrN+6LOjlnS/Jl9muIvedsdgHND+DH5w9roO2UlzJQ8EvsJFl2JU34N50QjJeIHF4CR3dJuz/Xtc
bc4lgluV7c82aBmxse9Oxei1PDPVexf8aNuGfZoSgsaTnBUVIDkPYJJJsoRXMXoA8vXfZXlwBYS3
fqGsG2E/lW0xVxcz+a+3qV4fYLAj+TFD4ws8vURhJxk8AxMElJP2GirCNlykYNj5+lnMd9Q6stvJ
BOVGU124LuoHwsmXeljC46QbiTrCXULoUXhgzknRLeNtg35J8ub4yTDEc9+84tUknlO+z7AsBrds
cqVTJe7ET7b+Yf3c3AduPacy3FSIVQdM4mvwH4e5DjtXcKxtZ227oYA2HzAa+y07MO478tWhMvQg
g7ynL1wyFRHvU3KXsRZD7QyJKrWhQ6KZtAYnKyROCaFhM2UVN+YNHXrEFLbtQQLBTYm4sdNiX2oP
3q2H+U6C5zyEpWt7mZTCC8WVpYkjsaJDUJRUqUs0zGgDWoSwhW8GbCj43KzTB1PflPdhjKqo5/DC
YcfO+6oAwHazNeL+Q+yyHG4Dxs6w6TRSww4EuBuoNJXoqZoeAzoODXVHPym2IOLuKd3UJVJqSPI9
84AfGTfWDuAQ2L0axSUDb+p4pRyGpWRjDsWbj3pxZSs90FJ8YXuMp+HE/hQimnxC19iLkJip0E66
hhspyL9OrLGW1qyVxfsjY5ywCDxQTQn2talvjRF1vw9PUHpBb/esgk9d4BmHm6+jpRhxndKdjJdw
HcHwy//N11rekhU9b30W+BYelLKehH1QJ4ZQMUC9KjR/S6CSpMZeGBt2iX/HgXxuviwPirZlFcPr
J3QCnbZe5yai2N1SsL4poy0zUGIsgvxLwVQv/yNwZAv7QEqAVaT0/kxeMG4Etswhb877xKTpnGqu
HQerPqijvi6PSwZSN7VwT4zr/X6dw2z5hW1YdMsA3/mm0xed8FtMxBOVVyt4wiHIsqRjKnJC0lhp
fdxfCFBZ0zkRsSAUCNdtL76h2PDgVCyc6p3D0oYoy7QHDOKmsfP7PSQ/6cLz/q53u0RrUeiSBrkm
bgFprRW2P0kNj/Pl/haOxq73innlWsYhzkJopY+/ZLZNT4UDWd8L6mkuN9p3XvsqQKtUKQeW5rLg
HTpRXmSbcg2apT8rIWhcqu1fSVY7V12rQXHW0el+chO+q5uLrpN34vlKXaphrLtumyZipJ3bbmWw
t6LprMqs+fLh4ODIU2hpnVMrvHLTkP0CLf8xralFjGmcnJ79BdV/GA9L8gpDqH6EYBlA0su7TQPI
inOp1q1fCuDUtmAyAca+ZaW5haqMzvNq1NTQNG8cm2cy8H5YP1obtUTy8hUESMrBBuIJknVGe1My
fTfSwgk6JygjUiAt1LeqdcflmLHuu+wQf+BV82NIUrQb0AV4VvfpiuILpBqizJKulEMMjYRagSy8
MplDkKghFU+4KBwh1XEVC5MbLY+BpCVVXxShzqVCYAGKo+TS/IgrDVYR3Ecezp778kSkUlU1BDET
kf5d7qiNLdWntK/uP1JYBNrVa8k8ANrGlrBM2LitnPSkneexdSROiO+0VCD8ze79r6DPolnAPdKJ
dHbyeYNRszc0cdkbFofaqOKuh/fj41X5nTRTaQ6/FLPh6mSBXgoZrx4r54/Q8HBk5qslaC89Ao6X
mXRrtXi/ELJf9ywawM9gnnld4XKqez3N6Z+0T6W1wmljup6Oiz+izWmgb9X3gNoY/4oUivO3llGx
H8v18mmw6F7Di5LeaagNgNzB9/Sz6kCj6GRt072olkJQ9LC4jofSBWUaySEth+Rng8wDRlmPKFNA
7WattAQrF3lf8WoEolxhyO9FqrWyJJLUAtDIuY+sLczrKuzEpop9viqfQKQEEJNSXA/p/NCWg3Nb
j2Fcf5Uh69WzDezOyZ877zs1qcIxMhH8GVgDbuoXdNBGMv1tG7wuoR9oh6/fXEPTubYgzZnrY/CE
/GAV9erXmVSCPLqirjUUM38OGEC0DXQMwPzoVkfMawBfTQMkzvpS9erM8Q0LOCNmphxF0CxjFygP
ldmP+r5Gq6lR1U6sG5ZxFF7PzbKJmhNoVLRHzpPuK9rpNGN6O/53QJaKrRKObLDOpnKTelY1soip
fmRi5xzvr4Ao0USXZIz5sRsoPSHA/RVxfPkZD84jDo8ju6GqGEU1cUs4HihlJn2mkq7KitqGcyWv
r4OgwPVXHOH+hbTpuMLB7oIMlOB7icCi/OlxQNpleB15hHK0Q57iam8pr7fbN8CPL3WS35UmVv9+
glxEhsCJGQC9dVcy0927J15HuSSf2wJiR4h0omRyAabbcrxzmwfgCWnRrYfaWu/LaZkanz6bZr58
i0kPfceJkcBvwdbum6LV9LKmfHS81mrpgOlG6CAaml61A7uMt2FWQA6YVhfyPRzlbT89p0znyDNE
DPnXfgvrX4DAuXnR8kwUOZyNz6PQUAp2JuzzWz42sy4B94SmXiLIjbfdBPPyIwBqeX6aukW20nG+
Gy2eRtV3SXLh24BncB6/qXf/apOj9IsjHJtqRwrMKY+A5nkOIXSWcAZywKbJE7lgXZ7E7kgLu9GB
su2vOvIgRTjHdyzO+NYdabwLFS0TbO6ZfRIY6NnG5RFti+4u4iffGOuUBPE+ltK7vvxHf99I/e2M
uTVlJ2KMl+lBu0D+3PZuxhwZxPouZCmE+deAN2SroJCADUcKnmLQVkUPbIqDsXqi5nthVeq0MZYM
3gp0mIOzLd1GGyxgXh6oUl1AdAcCS6tVZldbru6yIV6AJ1jAQLPpVCMc71knqfN20hAxKIJrwybz
PNDQQs5HwJnMQsVwkab9N4+m7X7L2izSGTnRtUp++wBQvvHH1uan1lcQCIFSOXRrCxj8Vw7tfAIy
NtgYpiOKRe10xvrRZfSJYAKFXIHXR7U/odtXuGYWoxAzVGQ6izC+EMJxW4I2ySInSp3xDIneWq8V
7TbTXB3yLG43MwLoB4KZARgtsEBH97JraF7Zw9r7P4WFKpcrrzCjz7CAOdPZ2fXEQ5+tC8MbQkFt
vx11+HJh6S9J35SIiVFjvCtPVg5NeS+8VtdFaFtNh3yhbIaAHd5Ao8b5tddoJ3yX5g8FQf15cBl6
phzVM2jOO9w+QL5Awc2dbM/pXFhAu5e6KazGR7lVFrrEvfaR5pTBZGDoy1cqhNTgnklq4QCoEoPb
EqKILyYKSqOgJFkj0rOqKjmDYT6ccXp0f4psoP4SAC86CbW+2hKEHlxeLlV8ad1F0xRKtF/1EF51
O4jD5YXZ7GPPV/tHua4u9yVZVFpkND3AqIm/iVO3YeglPZlyCfdJYjGQvhfgUyc7c6fIeqQTEDlI
c97NI+qlsGvdtZJSpgoeM/lKP721Xu+bt+s9ulNaVg/iqZPfR95ot63ZTSIbzwtjv/shYqQhfWMv
0Z8QIMymXNbWUstcF81phKWFgHETqbnOW0DTq3GqLB3hATQ4x3VRac44dF2bjhV5Qu7SNjIQ42VN
vN5kcV8NQfrFOZ4UdJ16MIJB6nZrMNZPJh4aqCHR/L3zaE6W+MzR2XUFHl2Tn/3r8FfvMQAdqsRF
I4zhdpWU9YKohstDSfVeqlBWqU7V7wT1Deasmlbp5TgU0FP2aWmeBK7KO2U+V5mVlLCRXOQw5mxE
oFDbOH1eQOVNdBDUIqzW74on4yUSxj9g8Z17ckWAXTjH6MMn0y12mhzjEcZTkkBgpTd/b0cOg1Of
BqeqMjB0sslIHJGt3PCJePPg9bl77chW0+vBIRtzhkiy28i78Gy9UVarxDlfCnjhGF4wRIy8AfTN
q/dZltSZIXYqRvPgrt9lEoMoCB+w6slGT2uce1quSt4JQw1UGYzGdyE2zYv/opsfD6brclIJtI8t
lpxBeES/IbI0c7UBddG9C8ADjFOc5rsjazxA4DXlchvP/hV5TV+TynfZC2dGzJLkxq/WE/n93Dv9
/cBjjZoe60ExT7G0SYA5/x5IcInz/PO5V8/PMCrHoTiqzaMJeJzFocqm23R/8goN9xHnHWpugC9C
9qKO0DvdyAiHtxzdCGCmGfise01ypVm21lF+UjlrfiM6TvEs4w4dXkFyaXZg2OP4HV6ZQ53DZbVU
U1yK5/Ti684G6NYkZKeTshNZlf8znVuys2Jfu5m7orXpijB49/i+IWCmguBiwF2L7IFTu9VPyJ34
OQoCkRXNqX+9qV3aRKgcFtULf9yiGHOovOq02wy755r5pbltuCi+aek8Y/Fov7CMTtZMRFAUzCtm
QF5Kev2/K/uyr381uNaO4kODzBxcmm8qNmFVfhFF6aNZlzUSNojB++7/8AMSi2ry2A2lQwfpTHzK
u/xu63Y3oglLvU5/Q6IP/aAinFxn9DBzvinHCCOeNAEGUvKTSneISx8DwSyHUg0a/l370UkVdneN
Gx9mcClX4YPtpTiX0g5prTwSC40WptlDWt4e1+zMJe8423m30S3TV+X0VUL8ZOnNAcLc88OHyVI/
a3VvmBYaImDTuL2WacJL943C6RNt3yPHMZXag5SXoK+WYnIGyJG7Y4spdDH6Ud4J5Hj25RO7vCT0
Kux5s90mxuBcvZZdIff5cDmwoZN0GefjXIjAsrQ0L49pkT/bKork2kMCU7gtRzhDrtq25uTBj8cJ
ydoIakB8e3MdMFuxxSibXSxykEifgTWz5IdeVuMZkdnfGN2uhQeayW41e2XHSeaVKGdiEbmk8jR/
ATRfQzB0+YYIDWP4lwhfxZWVNU6KFG0VELOe/IuNbgHFIM4Jlpp4ukPAiQ+Av/5TfDk0VCp8XjH5
6gEnqcOQzeEh8Ukj3l8goNTa/DeyShU36bHr0is3UxdLNOL5bKGY0+G63r+3GoQMYJI5WSuO/JE3
lR72TND1VCu+D/+DYbVRdBnb/2Rp7Z/aP5fBG4kp7GYxNozDrmaw6sKOpROb0a9T5+9lb0m+XILR
I7RUpfpH3aaG/yWoxqEym0+fKaxyxvyB+W/hglJ1jBIz+V2kve9aV3uSWKik3wDs5UE6jkTvAsJB
yf+2D+AUSq7XYdXVujWVZmQKG/5ScIobHuE1QPdt2ofNnLZ0GRheG63tdzmtdfTvaOiARtYlQhkf
+U9lT6aKG+JywihyVh40usZ6yLVX9u3lz1WY1i0F+oFgyYAZCcmOTpIvO/fZoHb0jXqniAHZSVJP
X7vvoLIuVaJ8xVI2kCw2SEraEa1xtFScaXHPQXJsWccbjwsjYipylNQ5PyT5UsNfpMGQDZtv1ABz
xgA1B6FAc3v+3BsKFErWDUPm7F0Lkt9aMEykaUQNSqaFi8H2zvIg08keQsDl7iNGQ+qFdgKWplGL
KE7d9BwNQJhVRDm5E8SBZ7z8M3xpGl1H/eVx+fRV/O502Pdl35UsMTcHLkY3p7QANMNx3fbeii88
XZRFQYN57hqYH6bWORl5NJNZZiPeEX3X5diD7c+7mcPY81tWI5AKlVucpFbAHEVDuD4wHxin+Oim
PAYU1kz978k8SzYXuImt8laNNIswbEORWfb39uhIDXejBgyhVa1d0KfDx0D+ZahZwPqBIrq8WImX
h4n/ffh+0/8ukIC/4uX+unGmq3gB8xK9teP+qRddrPMfES+4+CABamaCKEJDyWbcgPTjFuTbf9Pq
7HRruOMsdAcDBeBLpDpVdfZa1CKuvYD5a/hlRMNHX8dH+5AVOlKyhCEO8Oj1n1uZ3pDDXSzAOP0E
inmjLO0GPtjovCNzGCqhWtxz/ggLeY6WfG3fZGflEMsYxRLR3Dz0l94tqQl81H4pCLk6EMot9Cy0
v5mwPJ9R6vhsaSW3CmHv7Rr7FLYu4eC6U6M6u3tLeB6nnil+i9E3scj9IwexIBVyPZt2xxqyN8cr
ATC603H2el7NkgCjwT/61fOAQkzIEMByKgt+z138nK7VDqBq5Aeqmvg5X9cuRx+KRWnwLyqDIXsZ
GUTvV36Ewb+A24vL2Xe7iXPdMNFvzW5GUDyRXt4/lIBHFFM3Ypaj2C/Ssh28/IhywfD+l6gcud+2
wQI1Hw75fyiWKzbsVYvpw/uKVkOwbaM6SwB43Tiuz6M2mWJ4vL/o5ulGppn8XLE6WOcHf+Z8wt6C
htXj1XTBFrjzmh7/nWpFl7DNY6U0X0IA5jhu9pcVbOX4264zL6gwDjBBNKDrd3nK2zd6Vq9zJfen
XI/i5SjATI3guy3imTJtaIj70btoemnheLyEFI8BhdIO6TfZ73LG2eQU7g5mzYL0R2pSOWi/hPSJ
I0Wwe/uvqpbdP2vKWnEN0maoFsxFcSpXHuBaiSG/pOmbheOj77gPHx2UEHH/f+a9MuAFJnsZUXF8
oJmyoDS1UQgRcQORL5DjI5mjvama4OVtnPMVv7USWAzCX1lb/VTStgQJlKSynTRSV8ayGvz0CYia
JVlJZ9KzgkFQsz0pw+I17I7UdsK1uqffx6uUqLAIihQDwaf+cRHaCSgbjBYcrNjfn1sgDpCfje0U
TJIZkr9DqoOBeV3yRuwMKZlzS9q6u0VQzPzQ+NbcXpj9QgzygwOI6jkVqbzvl4tU6gM/X9HiQesb
hRMSPh3jlIKrde/oDv2Lb57tl+oZZtpGxpaHTZhWsxHd2Behj9/wei29cyxz6ezzzq8+Zc19Eq1f
7bZ2aUNrFPutKCvNC8tigDWy5tVX4hm81WWSixvXRnI8U7CwhhGilGtaJuksOySp5xqZorJbH8zd
tbjyJ/Z2ztuI1gmuBrMPzq+tGKc04TIwQTbG5Lh6vsKoM38/g0YUIsGs7qW5HLmfgm+n2e7Y7HQ0
XrIca/4MId/Kecfw1XqFxzqmn6xaWkNisuYHIujntVSiuxC0aVb79ZKgOcS6ErmnDHlym0mkILpg
oILzbck/cfYy/FE2SAz+6+9chlft7VkUNwBxlUzcgR51wH585tgAkYpimtcHuI12GSIF1CTZDoqv
6xpBmVHia5rbJjJ/KJfJRbL3xXMH5+Me/Yonk8JwJgSDc9FKEQYRjqnywQZX3NOHYw+3y21ROTSB
Acw6HA/yRjZtlQQqCMHkGv7nHpfKCF0SeNUpatiV9VSpYEF4EndVqoIhfnzfR0a9hn0QCxVLG4B9
5sNXKIXNj6S9SnWxBr9w/spZW1gvDksVcxAH8o26cx4RB37WKUwPLZkk4Yz1yzi8oN5Qb82bp89D
056uRCZnZvHaX9CVoQCbknoWLhAebc3A3+kZZcbNvANrPWXK3cW1p5i/HCMksL4aSC+5GtFToubm
v7DPcFaV9gP40riyq+Jb1x8Zocp09eB9ZtbEA174mayvc5tC9R+lptGflfcKg71kO6SETv3nxoW2
wmX1Ol9X7iiGYAPhOLdaly0RDN7oklNRxXlqgfQUCmSKVZFVghUk7u/U9PCaRlHtFSmqlOCF0Wuv
ZN3kwss0p3Nz5PyeRdrlmKeeIR+SfNQTC7/fWtR22/DVk1t+pwF4MoqMdAw9ijgUvYlwkR8IzBO4
VvQU+qwDufEv2VH3laColsCQDd458lBf5ZSN8dmRkemzzmmrUwImvf4wyVcnHY7f8TiKc34cZwfo
6ix3PgNibw4onnpkLAY4YlhNRkbtQm1aRpTVnLBD2cu3Kx6CtQRkMx8EHEYqMhAZ7n/ngPPGRaP3
J/udMvhjFeIJEXovaoGU9HhZH9jVTKSfV1IaYHkoMjPHI4CfVWlJBxd8p5ppCCGZoN2jFXpihKS5
Hh0pqEwEQ418yIhsjW1OVSoaqci3bjlNdaA9YyYM3bDopWdEW9UC5hHxlu6HHWzaYMqvMvSxw1Xo
mtR2YTy7Jvcu8ePoOjDi548iTc32UMe2hoWi7dwGgEqR3XAB5NRTCd8FFjSpc2ZrZcx9XA+K2Hdr
hWcjJSJIgGjMfgeBsRWr6AkAJkE5RdzP0tsoF98HGhX600tGPV+JR19+N77VooRfiGAuqVG0fGsx
suUuqPAhBBL11Fi0VPs5Aoe4g8J1DYudprB1A92k56C64gXjXyN/BH4fZxlpeC1AvtOSBV+Ztvwx
bMK6uxRERhTx48BMvSPKBHvnmTcvVmQil927oHTd6x+XkGKrh0a+wcb2kLKU3O633wjbXhiKZDTs
VdhU1yWRXaJJ9m75nsYhDefa88xa/I/APD6tgPlLvJvpQjxsrYY6PUFlyaJXBzZ/bYETrWySAamP
SHeNSOBeRKkcDt9JjSMP50kqcSt+eXbsGCYktw7jpNb4ESWEqAOzfXGD4xn64czwl6BL7Ip5I2Qo
niWJ7EkjL034Tu9CEyQJshZwOJsw/lb852KXzBauYZvhMNWrPyss9NlU7xrKKkbAa3LLkunpTCbj
2k4OFyBbQ65My8xosGK91s/9Ac2/8ZVYzJm2BcEIR5OeMPmEvlcjCQ1muM9TtcR9GqtFPaAjNIV8
Spz1YRQEnLDwOaD9s8KhwcX5BjBbX3xdCkeA706okdmYvh26ghb7UgBbhc4UcWXVtWxn3KYL23wB
WUwrshukJVYlZvY5fN2suIMy3F+pAapAFdAvzeHrDfq7EVAYH9QImXqtLG4x6yUy+0ePIS6C4hnr
BjkdytP6jQEyA3fEaqmUxR7A5pU/XyygvzXVroQu6BpFidBVI0GhMUDBZ5Q3Dy41IFTDVAyTi4tp
H59YpDi8jjdJwXXGZWKLelRV8tp5FicEuaunn5Ymcy2T7UT5FKHxGBEtWybHpI8z7O18CiTPlmOt
HCrG9kcxBsvSNvZEhZnzzQzJoY8VvHjcC9cL2eRN6xPLorLTgEBkvHLgfacuwnZKJf0x8IodBWD5
0euFOeSFfEncstjVtXXHAVfQY32/6CcKpXJYvhYxEQcbyPnwqHUWYNy9XJprjTs7eezY+2XAVPcW
FDUdnpcfGw3INaz0Q5BQB1J/pXAYNbqAmEWGWRMFRubiEAzBq8PxTTdegRkYEHx1dqxW/hgm6L+8
zzIvxzc6hwqrhkaTqrQHXKqzo268K+dfLOFzamV2hiKKj+xN8Hc0jDbB8MYKrS9LyWCKtKCpbUd+
GaogO+5WBuQA0UJMxA8I49QIiN0EdHFWfZIDDrjX+D8e6Uw/L1q9OOZlrfJCCCrbxhRln0AArGqx
zOAtuKCvqDesF8d1y/XY6yaO1jZhQvarocM8BIiGIaL8yZRM8sVMK5/iYZCekuJgixvIjl0m0ZKm
O/DmGhLQGfbhm5kIHGo2wGyRnk7tZaMO4XKW0Hr0SAKH1ehJrLvn9XRqbb3WnteyHEqhDtAvNORh
7r3kIDgqFLjhTYnAm9PB2HOaqW1OHtZOOY+k/8D/qyHvbJQgqdOGwbQC3YTZXgylaJkpQMiRZGbX
0HQWNKGx86vqC22Yw21TKPhHcOP83WI+gbO7ljaLC3I8sCbhgYEf2xWpXKndfdyRHUc5mOvgZ036
DezS/Ls7nCF1Ef4PGEau6RB+KlQQ4SaJoijm8zyRom1SYTBvue6OrNMUid2ih5ivq7WHJcKgsIcH
mOHa2gVhM+e674l1f7DjRfw5sCylS/SinxqKswaq4bUlVwA4++BsycBmbttCHV8ViW4jtC7f1kwh
2kvE7zeXbqtJLjdi+SXkbFOAe6K9NEk0nzY3hMwRG1ywKKHlYfWKyg1GMjzrknBK0s7quZgsgmfm
DOE62ozXddltdg3/VkrDOMW55GR2rd4qDq760FycQ7VTJ0zCf6RVHBzfB19+myAtvcXbl9Y1JhRL
WPPWlo5YF9yqWFuQyMa8pNYa9kGf2venuilX0OmZNQgIXMs4qBmOQ2liTaR/41N1bbCpwDBfTED/
7kwJ4pLq8PBCkZp0DBDPu7bbMPcV4R4x6WXdhQ1Y7G2hpEkFJDipm/dM6PViUm2eH/NVZFD0DKMb
qDI51G9JaMyKetj8kB0J77KFn7Jzvv/7Dh56uruEa/1trcE0ujtrHTKGfqkPKw/FPrdWLl7t37ql
wIEMTv18EKTniwn1xH81tKrLZte13kuhuo2bLaF9Kn04eQbGbZC5PxEMan/6jrSpkQR2X5V3jDbc
QPg3QbHVYmTlq7nkowTd3b+OcXMhv6scv3v9pRqA+KOk594Dworpp9ZO+ryqpTbzWrvTy7qZxX0/
c5coVsQwHmry1c0cNMPCCcrpBduG6oz7H9YCndxlTu7v2sPyw1SfouBz1Wt3k30utmpqykkkHqGS
QjgMR9L6qEuNKj7/NYR2GKAObTxNKDw1cfD25pEAY7lzEV/BIB6ZYln4V79O0y3UiqMpBt+u++Yb
TfYrWq30NFc+JsnyGkaZ69a8APa/xhjgoyW11g8UJghcOOAQ2iTCt7onv4Vvb4RcRkRqOPMH/t1D
UB9NlB5UX25NbKJDU7k9irhaqz1cpebPztn5yfumIKlXaOtwLj0yV3EGSVCAgyEtIDOjsH63Tw4q
Hct4GbBTl/sbiI5M5/9sqjr3Mkrb9FnZNJOdbODHKoqCvg0GtHu+IJRFBJDRO8LVZe8BFQEVHMx7
s7MZ2gCKTWfAW5+exWxkq5OjM7JYvg1KmpmNPcO8J7IOPfP4Yvk3+jzyFa8JrDenezbSsXITrTfT
ZX8l+Afgo9qM9uOJnNiCxprnp85s/cycFUbLilsMu9OhQofYZsdtIvoV5B62ewCrNzCNKQNwsnCt
qTcX1h+dS0Ckm+HigK04HH3BiVoS9yTW7LPhIqIF+2RoIKaCC7N3p/eqPH1HqNgvjaWJQs+vSPIU
kl6PEXy/klLYGA3uHleUtmHG2RjSKLOHhn4vODW+kO7jSsz+vVR4DulvWPNVeTV/q890N4kpymU4
wbP7nTt82PpYJw+Npkt5CnmnMfp97SEz6FF+Hk5lOIEr4abPfVBWYFyKUZmENBHH6DbhNEKLTz4l
QoDDVCXtCP01GVwv4KpRnfSgEqnAumGrdKus5v3eVjzwHCVFTws/pa9nfC3ojVBv5079XZ0Ajc52
IdrJAYTmY2XHWgkHzXgAxcTn/KdvDaQ2gVxjQCpEIcEFW/p/5M9ssvcfjk5EwK74YODA05wgRU34
lRazfJZefWnOhqY+sL85RruSHByOLiDHR3mXwxhbtvtascBBl1ASZPYHfFMucgXx7ENBnv9XsIFn
auARdE7ocYvR8G67OLmRZ4iWNhhCUY2TUhjZZ1UyS5mVodAN9SYDTpgh8acFJnwPtygKcfjg/Fin
av2H3LROmMIQiuaI+q/bM8YusXpstq9RgHdMGOB9cBSPkT4KerywRJLfLtfA5jvlDonNOA0QXB73
VedyMAeOEEecY3g6tyDvxtIQapwRJ6cgoB3cJHLUObcPOxla/yO/0CQOwJfv5z/hz92U8TL5Eoqd
vL54v2oeo0qY9aeFJ3K5oG0Nr5VGbmAFjgQuRND9VnV1GkZpCFhaFFoShKUaTRo/PwJIQpXy4MlS
LPzArMy/VdDKuhCeR3tC+dvtyPCW0LbYa0AOCEdHBJY6GW1hbTQiMeTLjJlKoyVmcgbjx1Mj5W8Q
VKvIh2wRPZJMbLbYeMeJT2AzesfIjsBYLgyxVPYyytAOWpZ3af8YSM+PSP8SZAcUxxJCKw4ZO7nA
PKzCmFpnRiWdZOgCWZdey4dcUj6ZLtEYlOzk96WytGgHf5V66xObuRL1wlagW2IhXDA0xEwmW187
dxzsLd24Uz+ofGSo5h8XN1bvVBI6yXHRzB4w4AHpgxvUXsmly4wRlt5mN2lOcB8ocP5wPeOUT7YK
wl4EtVkV0fOiN0n1Gy/SEdME0X04nsW0n8SL8aaczqpOKxLyHMAwEpLPeHzTvOhaNPwjrzj4E8sY
UGae1JeJ0quv3v+uvVdOQrZQS2Leep2SUGQhQJ26xyyyaKi8GnExQ26lrVai64m04OsEX1gJQMMd
p+WwrGLJIfhUK7WWykq/OGTWDiV08YEhLQniEf6boSn6KnltdgLQG3OaT2dOpftgndHVwQ7/5qFx
WrtpsBCXJITl9XSRKxNUvdAmoO3V6Jw9rZo089xPKI2qj3hPIREHvL29PT0mDXP6yyfqiVsl6d/l
qnPzBNENHhT5Y6oOXBQPauQw6r1AAPzU3mIcI0DPgHCzGpfbnh/6RRtD+Tv5ke+9eXATHOy5bthL
uPj6tPwV9q+C2/6gN2DrYaN919DwcSpMvhqr9gbupKESmp0/KfcCoFKSNcblwn2AZZnb0C4vGnQR
G3vH7pjavvWHED0/M1GeUVYu/v4CJ9G/zvHcx2L4GoAeE2OGDQ9pEkKE9SHvQqpy4lbss3zGnJuV
IfgYLipdCYi5ES3oOIXC8t8LAXjy9o52bVyXFZ5ITajb5l4lsMTcjW7iKrpUnSviKWv1b8T7edPX
AkkeVVmuwgvBeffagqN68BtiA/epe0L4RFwo5x+UHB8ngp6N1pikrVn9fQ1wNzzvu+qzC01p3dus
Lt4EJTIkvzPu+jssVboRSWNCNYGw+huDLDu6qr5R7ZUWoXgt0oOg++JzXxQQJQeEjz12bWNT51U3
sClhafZdtvMJWDYmTwL0zVwzYv/LkwF8UtQiFBN+WoZ4uEHjLceIySJFMUz4bGB9aogFKY1AOEd7
+H93gVMjFGRmJ5EgXwv5sScVRMQOxjRKyHgAiNukqVxAHSAbcVr8t8szbEI4f9lDE5a4TXhNIbyR
h3SBfb0AWa/Rh2x6zWULZ1cqZWUcyNaAJbzRX0jzl3ezOgh/FvSbEt8vRUsJWJyHKVVeKsfOsMyU
sot4SR5mTaqHDn9cGAnFaDKkFNyUz8jpqrjuB7/yhMRNPgHG810m+t1jIVe0nVFrvo7iEpxfx5rI
cIcS0HYL/y+R+wksYeKLzo1jDpGpU7qYj9zThRphkJEZST+ykp71mABtSJR9W9YlGw93qLbzH04B
mn2bgxn46gviBaF1xd2K5QBiKFJh4hLQKGJJe8JrtFqn4n0oHYPC/iAqxyOL7Gtjn6neHoCmyto/
6PR23ClqonGLsHj67BrgdfF8Fie51EKebkwjkSNhObNcGC6kz6N9aShLv4I9WYB4PtxI1zBmXElo
8A2XVTm2jjgITZsFe0yJTJkBh8aN+ZsQ8zGwQaps1g2LS3ikzxZEhX9aJDTuPLhYZd0qCtXw9G3q
Jm3GTs8mV+1QgcjOuRle+EJKKtg7N1cNhfmdWf8Qo6GN+NGPwg4k90gF4tKQ//hDEbWbgdgG8whY
DnAXXfg9ngfz2yOEOjU8Jwnjor2uHbaeIlAeJ+coYBU+VhMukW7JjKuANU/y52A7k662minXSKnK
jQ9s6Z5ZdiStRxkvAYw57BjccSvKzCwGWg8FUtphO1rwxt/cGJvfp468hLbV2l0mPZ0UFHui6zX4
gA+1Hsck/LK2mx4DcFVvu1Xmq9tuadxHJIq78s5bMPAcHByWAGqNjVjNVtmVeiHfVGmR0ohXe3ck
VhV6UY0qSq8gPWMbxWRFFpxoY9FXqbbkRfZY6rBICdHlUgIXyvx2DGGOLlY7Behf2ivG9ZzSRwoh
mvwN1cuPmCd79mrrYwA+6b006YiOppsWgGtafuQwqPqZojG7gPiwjUzvsyfnxxXwPULsFNnUpMSv
PSS+iNEvUggRW6kR1A9obkglpglwzcewBx+vRjOgq2p2fdKZvdNoYyRllGuGIn3CxICFVLDUkG17
9I6n4hegbwq5BYalyxDDF8dSSX94E0YKidgT3+i0CDQ92tJvqgpCDyY4Sb0biC03qYzgzvAL8+Ki
ZeoyEL31p5oEXKIbgkjfJq2lkMypQjEfkUSozNvD0RoyxLXaaS9B77Oj9aUnSz9/6L+BXpHFYB+v
AxL5uPu/7ny4XAJfObQwo7P1lD1qEZ8t30ULoePCL/cbJtX+d86xOmCfL/Jq3M8La+RbDWmF0KIl
Jhy0n3SMcce8is7jW7MWVW+tbwI2Rh4IERiATls3NiqkLtRXkhUI1KFtoYVfSPGUlO/Mi2HPfm7y
ePCNAfFZsAd6Uh8C9Y92qiuAHe47llUTLOroht9e4ah8bbmw49nvT2adXfnFW0f0aYpBm35O/kgr
5Ws/p+WA631AC+ddQSPnIC28q4Efd9w2qmHypP+Q9IHelGS8bOKBfCDpo+P9eMRfEERlSgxUBG9z
cQZbETOeF2pRmBY0WotOSDH0G7lbYQnQU/hlGtDirx7oe3v2Ukli74xpX49BuqvZwo3LkiJWU14m
17rMegZoCrgVlW9pn9FjXXO7/OnEL3Mbpl6xUc/m3N2xHwYa7FlmQCWFt3ifbyquwmoiXH+bzRIz
L0wgXqToFfY21iZGMaoAqcXWw023LxA8SuMec33pNRnBye/pXVIJ2mX7Ktp0WVsJZxjsLBp1itJ2
GqHEkxHg1u4sDhJkj6i5sgJcjcAeotbWDRGy26/K6nc18h0ICfs95ZmYgP1Rffl7Yrj6DZIWn6Sp
Mpf/sAx7A2g8+RIbPPH5I9zXVKMSZOFf5pYtNC7hDXASBobZEZF0e/0vpRTL3moCUHKd6cfbaWss
sWsB5HXfufPoUbV5j7MKjWlhb0LTBBgZyxN5c0uZ2oGlj0NKTjG6z08nOWOmR1D5QqyCsLNpIG4I
ZAeLeIpdY0z7TEmR2N6f/mACxP5CkPVfBtNqaL/sHipH0s6WBIDXdSwDzrhzo0nACah8zAAPFzMx
oqhNCUKM2MU4orszzU4EcgYG7hvydYcFMTuFTOcyvbDOQIRbGCzUY92F1Tr2nBMS++l1k+O9ydHr
MqJzilG1HZPIl58j33JfRToz1cW5fewV+kkVO9nkDDgP+1Fr/lpxhBbOfdMjlBjCDKkLMQA/M7JH
P+S0+nQ4tkRumKR2w1O+adwPN/CzkHhEnejLi5RImdtieRFCO50hOTf7OlSQBrfVuGea6s6hkw+J
79vJAXSzqkXC8sWKBhmxwH9FNkHNOgRSek+DNvSB6/CuIXUnWMSwfDy05B/kJpx07WZBEyr5CSQj
8OSFKNt77cQHx9Lw7iiJ3jL1Ek3Pl3E+jtF3OcDV/3OoPo7TpA5vCpHtYJ0PjoyIxqnRdIsPctf5
ku4bXUYo5I4qoLA8pIQdiDs0jqTcWOtFhLjp7fRxk0tnrdajOiUqNXylZ6ukhJ3hod8CWqafB/HU
jDT+cak49ZZKzy3OYqJzBOtLN/ypraWOPLednw94Cx/mLW5tcEBswawTVMQNUxaAhtoHGzyVOU6+
VDSgXlBljLSR2S1Kd1lW8/RZInAv0YAVnMsbGM/uXqeWdchGGilCpIJ0bmTqEtY0wcxptpBf8i1B
a2JWl9ZHqIRAgcTXf/QeFRyFPmsSPeo9WqFnc7uKGby0UQhyjewLzHiSNy0K6/Y2aMRf+8bLYoW1
JSkP4udlZgP9biGUMaPb8fCmuFOON5g7eB8dXe+KTxX/LD+XZphJrfbbkgWnPrA/5gjBVsLNWfz+
TyJDz9aYGzxBodEudcTPhazOps9LeiFA3yU3RVdKChtjrAD2PhZQ9YNkzQZnFm8bFeBLUAJR+IV+
l/9ITe++JOLS2cm8QZpAX9So8pooERzqCGBThkIK6yJbheFP18E+5zWKqNz1OtvijcSW3VuvlNSg
VLMK9qbBD6rPX9YEJeYmUDoVuX6Of/HUbJDs9fW5ZioW9FmegKNGC6v+n2J7BVdrXphsGesLG+aF
Z+GHARu61eAVx8TtTBHl5Z+8F85Yqf2kex2YnCAJAA/SlZ9sBWmy5saHhPd//SpnXBKpFFFtRGak
3sHFoEtGEGNmmHvwOAbNn+64Xq/3pMXnpAgaZwO/N4qUhfXUpsiqBtsEiQeLq7Dcec7TI2soF4ri
gMMbgcaE3kNzvZ9vyBTHDflaMwpwuV2VbmRyDwA36LRnYViaWJCXIDV5H3ybQkf7jvsjWRq0hELF
KLZDyn1mxQR06uDRqJJf/hcB1m5emIHpuSSj0ExHR1N2erwCBvBI+lfK+zyVucws90SWQ+U5o4he
pcmEC5oOz53H8UqLbe4oDuhwHB0OEz4wglgQt+ZCJwAM5pZtXRQ7MdFG+KRB8rCQyhiGBeu16SEx
5rfgO8G8H1PpDUhW6iYkaJ4l1jiZaf5VqR8TkF4TyzPMoKnif+NWmcyIJfdTNp5+pQjwKquBzpVy
jzvalbIWe6X6W+NKAKPT3ohshTh4MH+jhbYQ75spCSuTO3n5LvqRIuRrKKLO1FF81hKwg8Hx4WuH
KbZQDKncc0rNzWXPFp0Uy0cqzRs77kaKoGy5yTFTE2Mzx2N0UKhLLDtC8w+Jdz+2DBwm/g4wdb26
4ry4y8qBRjDdMuFObnO/1B6H+sTCiAZZi5MbZNqMdnparhkHmhPfvgfTffwI8BbgdpHrL/NxCOBh
3kE2y1ntIQtgiXwaopvqLrBVFqtPjd0yaJpHF2VCSAWw6VUmdfmJMgfHXRrRdqBnoXFIGgzUDWIw
jCpJbwOJVuDtF6cc3SUpfoc/lNiRmAJjB3EFViLh3aZVU3M9HEZH/NA2z2p1fcmJWEolrCA728MI
nTCNbskEINZKcJ0W2Xw04pbq3uh0gbVW5Tr7IBZSdYcArU4TIxR62OEjXO75W3H07nyf2JLOkfsD
Vb8AhUUQP2cSTNiwylafjSWGWYhNYkkSiwampeZ1Ea+mgmHCpbdZ+UtNtAH/dGgp0xm/ZGTSiH52
mdja/1upoUl8wIGPzPNzrPNY42sV3wGE15Ly5wnhtlN0D33agegVVDFW9VWpHpzoP7LfghCKoNa8
4iazbQ2xyosV+HAi+JFgu2aih1nFUxS0xx1H29U+TLKKu7c47RPsZg/vklglktOybFfbA/BMBoJZ
bqFkmpPnzsynQ60QOH/B6Sq/3zrSK27Apa84Ir7kCttU5bRNjNDIYitdDe65Y7BABWfi+9fYXR1/
F72SibkAZ5PgjLUDG2fmsiGrFJVpKn2AEPBK1galQe1Bw2tjZLM/5Uwdj26JSefwwb3a+oEFG9dg
jWjqGCBF3qESNEzZl2JQvicgn6APcn4KW132dY1GzhYykbMtWUaV7TEza7FfekhGc9A90jnZqWkL
d9lRatcQemwrQeiEieheneRCaR4THsoC7/T+2WSif+KUb6FtcoacwRwMrb28NiBwrUhRS4H2WFlU
9chIA5xoKaeGkiJG6N9sXQ/AG9qtjTlYvS/YTPfLgVA6MA/6Ft7uzG8mX767lPUpNOVF5ZSh3NvQ
QaGE/8YSQp2wzFNafZzug40lW6aao/sAuA2MVI/9/+Bg3wdhLSHudToLsCmwDTuKPgVbJTU8BGre
36lUxre4ttW1jfywrvSDnhKtLxF0hMUGL2MwqhjYSDP7QKNyxoJ8w6Ivqt9gcnKUFp1qh1YLfaAc
DjM37opmKjraNk6yTxyXUh+hUWpn3QwTSuQyGsW6VGX6l4DSIGadonp+9xkyoFbv+2zfBotZcGbP
lSD5+Dbkzw7SjylDd4PvLjj7i+hRfOs57UfDCac7HXJIOf17NdSoxnMKPto2RC3QVClxmSkEBNji
V57udPD0BFjZpMn7hZ42goh6EW0nNcclD7cVZZ2lmNtcjFwtoC3wV4IvrHW8SY0raYRZJ3eBab+t
dz01r+7Dj5vEKa2KL3VPPC9ApsW619fXsm1d/9nLwYNBlXWBa6S1ZKD33q02VgLgXVQMvoZdfPaI
NryQcGsQWwkTS1sQ6iB2qWE+hFrjMfoWWPYcELVbA1cdH5kPQWK5zfjmDIinswE49lNr80LOK8ea
/0bt+VuFvysa36WRM9vzAxZ+IZXEJdup8Yxdy8SsLYy8uc4KCQxZ/ct0i7bxJNvK+3LdRca1VoaP
HWKz65el6Y+ykX3R+iXAJZ0PSnMqCl4Jg8IcVwpjbXyp/Hsht0DnoRV75vfGVOmQNDIfZIYd0/V9
+tF+V2/Nm5BTrPCUE9NnpoWG3GqVKU08QH7UuuVZDTLxeuvD8QVSDym7YLET1VxgmptOsLB65IbL
NRMiu1NqM69b4BpkNDPNJJouebyDehk5PEGnYARIbCgeaq2N1jlZ+ZtlY/cAEZwU5B1GS7PtapL3
OXm5/h/leSeaYlje1x6mOjuFmj9qB1Rz813x34BXAcUUbzZy92Nqd/uvS7IvvsUTmTk4q4yNCB1u
tETMjirbVwTgQS/mlkzS7AiobgGGHHpJ04NQyO+g8Al6Z5LX7CW+nu4AAAF7JvtoBVU0rCpOcTGa
dm8kpIISs1oga2204TdXltxJNBi2Mlm4eR9xYuyVVTa2xgmBpMIz9u8Wm5AObC7uSwGhWYFlknvk
/xQrpnBQZIcWI2C9McCKK+WhyumqGWfHWPP9GEN35cU9taG1X63w5xGInGNiCymKckMug1MHuExe
QPvCllg6oxMw6I2rQq5OWC/v+L6cGJjNa//qauWpsQir+mEQZQDGh+G77pMtehoA+a+sZTc4y7/u
vZw/0YleT+iaRjl+3FXeA4SIg4loj0t8qsazkWOiqJafTQho6u1Q0WR3kzp0g+gRiA+6T9hTfG6x
cge4/oWM/1ed17uMWYiZzyK3CtjEgkA1eqKjdw36vS9IXJKiceEjjSea7rxQR8NRhw2tkCC3qKUk
adNaJkIXBUhL3fNgSmb7byMDSl8TyFf0llH0K+tI8vQgwuZsOb+OToIYZZBF0DNIh0JztUxVzWjt
YLS6xH9VIqfwwEpY8lGgzRapCGlKGTEocsZejlQRnelqS4Hpeowd5UJ9e4fRc79+vOPdkkw4FAlj
7YxQIUSQwvcD1y7el3NHrQwdQ/hKn5mIhiYLak9lJbw9NaueDaqjtQxclGAHoGEOFTkKVmB9u8N3
fToXyXqtufhwrFHRhblHF8MHPy0+P7fM0bgI6g07yw7/2CGulPfnLCKbWjk+tzyJxuVJzLgYCRyE
+kIk1k1w6pWdiCfDWAOqONzrZrZ3mLXY59IeiDps3PJ3e3Qy/HUAHkZCLhpWtKx6jMjqnehtHVIG
ahOoQ4WcWXtWxbXrJwkAdZS+B52RvL2wyJPhmBm6JBcBnNrrdcZymDHnzcRnHReN78aFf+RsHidS
hGscL3dkI4LQCeMT7MezSW24sbKFM7e6/abW+RDRBpCusXHYM4V3qRNZI686PAHeujy7aLvUArmV
Ev3Ieum0ZixWxqUOgNEXTuMDOiehvXI0PSp/url8mjzaXftN9xRp9qOKDCIPEExB06vSyewr8Fck
BRfPkqd3TL6mHqpLTV3CL5/cW7GyM5AUxmLLfOZZdZeRRHWQj8eEY4bLlk+B0769RwoJPoBiMcQM
vbQV5sQRqB4pxWPx/0J9UZByFU8KxUMeAt0EPA/Ut7o90/5WAHDeb2kFruaxnPrWTiZUULsX0UhS
LetL7Xy8pG/VeerU/vmJPLYivKjTEZGNQ7styuJZP1kIGvgnQZfZBjbh19jKZ6jjM3xJzdFFurdp
P6LddH/96AiWxPaXEbUgio0GhnMg4Gnko9zuNxI+gQGYdaergOfv6n+0Lw4hKdcaUWGMHz2SAm6p
QpGbGw3ifj52jf9Luxk6zvNfp3P8Vj4viqwzCXaQ+ngrhGpBYiA2AVaP9Pee2AsjQPvpc5MZZ8fS
Z/v3DvARCoaG5/kbuu7yMQzmAL8F568JfP1NQBF6rmhKEDn8ljeM4BMiH00NXBDlHboshI/7vQnh
rV4WiMMKsCFj49QrZAkjLFfbTwN1UZmJnZyrHDtuV4Ih/bXx1u7I26537TSMEPLwakVdqfTkQ186
M2/5y5nKOVJV4RmUsujbP0GtvKUCk4Y9LM89/5ms6WfQHUkkM2Ti6gbrMhI6bLy9zDXKJnMPwmh/
BzSiGF91XQynittxv2IOnbtDjeDdKqF1UfXK3K7bPVjK9/g0IPOdAMOAFxddAS6Kk0sa125ROI1C
wu8y8pchqDRuHJCLes9qojXNHGFQegtD9QCa3l0Ekr7UMsMdF+xtU5vFCjSMjEfIoacWLny+RDS2
vcjdsTCMZGX+eclotglxQ3d7FGctk3G3g2jP+M9c3/9v6f1XWoD6qysFIw8xMye64vbB4k3nCifV
gRmmxad74I+vn7psYv6C73Y5j93bii0DqV++M1LZl6phiUxHRhgqKoUHeKQZDEOyJ5bq2WC387m3
vjda4su9wQN2RpYJ9D71QheB/9UWljlCJZtLXFk3VtH+O35K2pI5h2XBB9pA6dGxDMcrTpBGTTLe
OVO6b2OE+/j3uh1Jjg9wLwJC+rVNlVlKNoBaaqGC6acrNghcYgKGIhJEt8hUh4m1bEZRQAnX8khA
jx8g0FO2oZIZZcL4IxIl1mxhBgoL9+AAiNb/NptqUpUVeV0P39w8poLFkehpn6gxB2MKuaQ39Lj7
tGRnGESEvc35yndf1ylS3v+FNg5y3dGsfVyTYQ9Mcret0AU4WSp8HQ7dE1xIyi36+CXH3e7odF+b
NxwMvKLhZrTeVBXRhRHaT9TieomX98Q2qa7e48UG0C7ypWZI/FDJvZN+n02C+t8F85+23UREB+lf
t2/R+eVr5zZ/KQqRHIpZTuJ4JI1PTMB4etRfFGvCt6DO+6S8+hyKi7MEiTmu858DKyi8HiG4gc8D
rEASNipTx+ndjUau9L/o4dFm/bHDJjYEh7/Oj2zyb+M2IUy4wLKu7zkVfRpdDTqfA2x8iqpwmHvf
FWh7UN6ZzwbgJ86z3jMqithAb0axtUTpusuEWZBWNn/G6xorrgkge2tT/s4il32or5h/kFfoLJ39
4H7Jg+hEcu3cUg2hW2ZJwaTT0gzZEqbRrQUiIO2LQZfblhld4ayYXLBdnD7dZsbKFAjR/QhCdoY/
Lt/gGG+IgStcFiOT30uJtLPwBnZf6m1ZmoAzogOtgFLYEah6paggUtTCJG6Vmjk0OKdc65Z15bKo
wM7Uz2ymcFrKJ3tMEsgVCnvJtnQfgJ+JFC6AaH3RUCeQdU9URB46sDG9LzZf80sC9JDFEJg9FxR1
DvimLv6gNXUrbQcGPP9Yy3olqHDrm4FnxpzCaobYGFqleyAEsi9vwdsnkH4xXIbaoBVeP4xvDCO5
1bzGE3PknEck3eNMMJsmq6ngVvf8dgTPqHGwxKMus1FvX817BWicdj+3NFHIb56RIKSZOSnfq8+M
7olsMjCIuBtwM+o7OldXfHM05ZNzMl03Ffin3EYt9ETJF/3TTEQv1pl8uCtBHSleuAyzfVf70T/l
iQyqnOeQ+729BZkCxMvFHA9IEI6x9C4eIRHw+dZH+AYLQPT80yD48kUPXqf/n/Q6w6klps8Zz3Dj
IcGd8+8KDyS1O64M25AF851h2PvjRcAnVSHcjqQfRxUWXDsp6AVcaLqyn3pzkSvtQdtF7r9CBi8O
Zy0Yt2t801uOTS7g1r5wnaNbKA2vh5X7gGUvEcJfPfXZtqmxPu+5Fw1z4e5WucCqsf5Sxx+KRqWd
K0nr8EjAXy6uw1+IQGPD7CFmmw2ohih/ypGWnMVnYkY7iK+yeWJwxhegYgW3Ab5Ykkcq6C6leNBg
EH+1qIOf1e6LwD7Ws29QcROfyxjwkj3QivDuVZ09lD7ku98XVDah5xx83Y2fhuVH+2NKH5/uKsVf
d7yQ0yfAVSnuu/efFSnSEkaH615qm4ChI42K0Pwfm6knt1UVAlX4M3mQQ5uuoBCYS725V+zu0Qxh
glXdZLOINVfqr4qc2Gj4f5i7t/5A+9GuCCfkaqjaaYOsMDv8SIp1SMkrRtHGNlsVZ4XyLF0V7gxG
Rqn2nkjk/FDpVZxBXbo34D/QAuwA9JIU5nHe5rZ7pd70NsUaewRyLmj/7BlJ8xbwZT4XDrnhBN+b
I+UC+rH9mpaeYWVW/RZC1PUFrWnw4DDlY/o0LB8hXpgUPDGnNLa0X6/O3/XsQgsb504fOK1oVdFo
yVmbCvsXB8xPelJbzqqOHp+XmUy8Q/mxdN1F+J5nfBrFIJDHY/p+77a/m9kySL0I42JB1Qty2OHQ
9/5jB66sAyMbggpKBvauXJ3GFv9BCD+8ET234fT6Pe8zRxDLWquhgxipzhbdR+rTvmZpr6aI7EhH
QcLqrCUdUwnEABe9dsYdZbjPaqKs9xwDspgK+agc3AL0BpS7fbKQ1gUxjfzl9FadlsLyUlwL29A6
RgWCSrzNWD7IWAv499ZGS7nQCY0nsnvq/aoThxL2tbCDPr3ZPOgCUztpgjiQ7YVK3XHn7J+U7kO7
KET2cT3VTk0Ocq6QPlxViAbHA9xt0gwhQ6c/dtYfyR9Crh7qFmk1jgm5kVW9r8NmXQoNy2UHItOd
Q3TLchjSTmKsNUnXJB5Du87qX1Obgrk+g2VbVp9pcf8JVIBwE1nmyIHyR24TvPZgMBI2cgxhLuIn
Un+6b9l6kGsswf4+Bw4v5WAJhu2zr/1JS0v4Tg1XSfifqPeoJlHh9zVc94pUe5NSRUVTi+PVzoir
DdxSlaoHKTGiGpbJz85bTxt/VbHTG/0MxupuMRa8+ZWzFTcgZAXfoo3EmqX8YyZvmU88equW8POS
auZtF2MK4+UuP41WUOQjCCmGpkIMMCimEDos7791n28jVqlf5r8ozqSAcxIH8YDUOu4gj14nbQxV
yIlCb5yEL+kHiWQabaNBTzd4Q4ZCNYlNbX9DfK/O3zPuve6HzjLTBxMhTE0I1PXz5oFdufyxv8lN
zoHQWVLnPJQwh9+vrHF9iRT8VeTJAJjdUgPChrPv0k5pfGPBq3g2O8uJyptWQTO+WC++TH0HGYuV
mvHVh2xcWlNpVLniabVXttKlyOA1lWCR6QzoI5la/JQY283Npuw57uklzHzI1N1sxa4G/ew3SAwC
YDjZ7W1Goqv1eUpSn56kRReNXMYuJU4RVfLNEr1ZbPjmCw9opm9MyQSKDcbP73Ac1ZvorZ1Wibug
777y+FNlLb8ZDJfJ3fK1lx7WvL0BqjqKFn/uuStMCt27N8mn3F3Y+RHW3ysuO3X0UU4Jq4oSVrs4
hz8dBaMjK8hNA11ZAZuEBCthcHv2cAnsIROWBchGNqH+8/9FbJyF/DxWJXMgwSkay5Rs3xovru65
/JZOkjBNra5Ya5AYS4YfvDCjnLw706uzB9aNPfQP0/DO9k+I/tA3HNvT6yNc8CN0hc57b/591LGL
rLZdGWu54nnpabWIbN8E0JrB2/+n2vs0Sm4yJ4mGhwc4m31IYZ3C1qO32p76ZNvimZ8R6VY5RlZ/
6dn9H3NXZAGIBaM5A1v1dCm4fLcc3pDs28WSwx7htCfONfi+TeXOprsrR20isOXIt1dO2lJuioNn
hSUOggIvcNK+0evR2iMc3B10FSJiGtuenGWYUzhjCzirEf+uYCg4TN044omKbmPjZcBtUaNquIDT
a9FBzeIZm3J1ytw8sdUlEoyqDL1Bb9/xwSGUELH1CNel8NrHIsXzxA3tDdeigE0FCLqwTcx/VQ7G
hd7IoFP/7Cw0qFQEQ/OQa7Vlfr/aJMmW1mNsjX8mH7h4BOFui/1Kaw/OWxWVtKkF1+ZUnz5ECW/p
LjDl3RAZ9d8Rqu7JYIC9YnxuS+WlguvP9F+RhhBDUu+HeNwPkF2ZQ8aixAyxF3l2o/m9v9LTMEvw
SMKgIwgW5zq3X529CepvejEbIjNQ7JxMkP/t1AFw2hl6kY3rj3vW9m/38j8ws3tYef4kZhfVaPEl
2noO+QsjH1N3iUw8uyU3aEuel3QHvbkJEfjFzTWjJvTK/tXElo4CCFMu0f14ystMvwVN9s0uFihK
T3AG1igqvNcbkmbkYk9cZzaJgazhWITDBI5nKLxDHlgcxjwW/GJ+ucIHJgOrIqUT1KD2/PR02K+O
+9aawBWQgvJjEXWsEH2Dre0JItu4+RoaH0okLrNzYt/L5mIcT2MYWUE6C8ccxlDobtohsNd/9Gh3
kqXOIx9Zsm8+hPTWwlVIvbdzgNwlZRHrl/TKaZt5MrJJmHbWVA3hVEuA7U3ty+cjX0wflAoUSZPt
zVk7B2JLlASoWBxF8KryI/RdLVvrF6Bu+BgzSbItIAyqWvB4BS/sNIvShqJPpVYCLiYYMdapSIJu
rPU+8L7k7hZJ+FhMd0JE6kQM4jHfPmUecRMSUXy+SwWkn3gJrcHAQP4R39PGNaZQuwfAUVKOhaAJ
A8PN4gy2+yHN1pqZf3nFNhmk9lkRlu7e3En7E2pYErU2ng6uw9DtHj8j/iwYJa4AnJiX9MJIXU09
AgjQf9YOLj1Jk7jSqInXfOAh+WB7X/RZ1W0eLF1guAaLv9+3beHRPYmxVMdOWgXEpgmJ4A6tnt1K
Lo1ANGZkNgZgi0hqU3Y16+jNZgvmZSH5MrUzqr76MmVsR9EFMWR1pzSNFw7zojWkg7HoaQ/8lTQZ
oNPRng80e8AufsNKEdPpHechUzvaDlk6Qj1YBfNvgEaG9MbriICLSHOgjFTNwzDAzlC42ZVr2BgW
Yow9G6qUtwWlwoKpDyYPFqBDj880QULDTwfQVQzvF15C1O2O5mBfQWXLgfu+WiyyizCIc6cpNdvc
wbFe1Z2liDPQK7y7ZLM0CDOlbiNvIEi7Q/mPtstTdXMnFq2Hf+vYtmy7hftLyVOSwt6wRvWRFjVL
oipuNqvnWyQDFI83l/UeYr4ONX3ZwCj3NHXMhRpo6+AOmDGMLSQVll+qHnI6rx98Iz51HrORQEBB
FM5unVPrPUc6ZtTPuw1x87zYeZqhN3yqHO2ghfYMFc64ljUnVUdAgw97XKfk+Uqri4yzT9coa6v6
jX8fgQqm6fWgRq8e5a2+bXrUWtBsHTzYbs5LWjXFvDQ7bXsiW8j8if43YvRZ5z/GrGqMYQHXH0+M
oRO6CHEJiGussbInDnDjm12Bo4nhcOrkU/XenP2DYoVsMpGBrF6WogCLDwP4jEViZ2hpTLKm7H0x
JLEhUTpCGOK2enFySxSHEUcpu9QO8a5G38gWVQlzrZCpjPOhiCryd342mQK9Fr6mG1cLcTvUh7z4
55znhrJEH3Cdp48QWJl9wykUsDwU0Nh08eBQM0C7WCa8CQrjbl1cgvWQcgfLbIPOGGj6X5n8cheM
Rx4XlfO5kGzrhoXsJukMRWRxvgj1d5EZIzzt1kV+DPiZvx5K2hbzA96/82P9TLHml7/4WTj2MmCP
hOoB2L+ip2eaebPXb9X0t7Ly1Hn0EdnKDP7sCfm8PiJz+qQ03Qp5LixHs/sIjCzYpqPLmcgaP0XX
gysRiIjsJdM3TL4ITGL2kyQPdP2DXR+WABzht+6lUj2u8QDS1kWJdOS8ijsl+ubrCfSmFSc3W761
vDeP1LmvH7bjzv1XtfSMWbyNNshAMYRPUMJHX02jbf3V/6oqkO9lU6Eie8L9wRdA+wq5pm/1X9bk
BBIpueeFwKgknsz+YrcQh7e5nLrrDf1jETSvwkofpbmGTvOVbKqijeowrppdmLbZ3rIUzCs9ci3L
nZw49Clc7/whcUSHggC5a9ugTBH4drKSd/BirdoPaAvqzzkYjWTI9Q022TeSx8fSCFGcvhkw3qVW
qHO9zbNfqDNKhlG6fQlHmdWnVP0Km9kmSYM46EpLJQO/N9moJQ6mdmJKkQ1S6XDkRUPWk4GdAGBr
vFXdNOBS31xQ/DmGvb5onzQKjPEIsi9QQnMn463U1QGkHlw1FZe/eoMUTkRzjXp0xrKprPDysTzW
djkghZjGvQ33pLYFhaGrUtlemgLcunY/pI2l8ap5TilKMSwJOpHJUz0Q4wN/a4bQLCwQJhc+97RV
JuKiNvEjstFPDXZzMkSlvvP17La7kagvaRrnorGHl0wxFxfyDSgAXZNdL5s5hS6nbH94J6PQRcHs
oVRji5PNBonMGgYpl7/rndnBRsKYu3Fy1AuduiNX1FkdFX9a5XBXvhjkdrDHbh8McsMC0jxalUaU
og6Z9gyrXK1Dq3N1qQzjBzpwRz7LGKkfMIXd83lgc1DFIyXGTyhSXUlcWc7OvVmx9S4iGmBcBg8X
zd6U2x4IGVVtzh9ZLl+jOxm2pb7yq2niYm+seJtFIkxAIpVs3qPQFaVNOpT29KC/kWqJKlXFchBR
RyVaTmRHE6+S9ixHYQ/5XULgzlHdxA9eaGtdIOG++1JWql7gglWbwhXIpTVvCHnaXgIEBpprvwyB
Fcb/ic9C6a3FJCGG/WBdr08vjbZ0Z2oQxXvlcj6oP2+2TXr80OjYYtNEHPdRJXHU4zt1mloatkht
UaKZouHUOx9L6uU8NiZGXO3BrmnJPzLuOZU0WZ78/J9Vg7YGjGX0pzsFcqREx2F7uSEBjvbOKVmv
73MFiGJjC+SPj15MMcUawAoFvnhVYs0pVXVWJQqJB1ByZiR7/yOWQqtBmojh3JuTBuE/0Yo/hxHC
OM5iIb2IOwbKaQqbEOjLBYy5xGZs2PDc80WjRYBVkbTddyYXmOXk/INVihr1ZQncn8DyjedP6WSg
7mTXijvwmCkQLW5mMtbudulk16G5HNKtddHIbcuM2I+snm7JsP/rpADWUjUpuU7wFCU/KHKPNumT
E2lFW6IdrrjU70dLeknjzPdidWDDC9Nx4NwLbuAIinU/qEzOQxHfZewdaKHdl39rCibOK0kwdOWc
zExxo1vnwlKgwSvM6nsMRRr624oYC6+cUMVnfrlCLKCztFX985fC68XkOC0O2kpA0KdpS2Offxjr
XMAbXwt2PimHb/3YxXReAMB1JXWdVRlf2fhpKBHobJG19ODsUHWGNH3JjM6PQgPDjs1ybjEYhPhL
Ckq9b3NivS4sWSk/kmxybXKGe4+52B8OOfSeFfGa6Ksx6HjljfMTAPMiZbBzvgKu0t8dJP7+tn+Y
9ico7bYiZm5GSwN/dQB05F03xuZhT4y1cH4vuE1amKpCkExS25whAzqen2otJZkN4vFWbO8wKUbN
8LWlBykl42ooDhDs83MxlH4bRujHnu5tjSrQJTRCskM79iG4YFheK268SW4qeR2/MCW+dodkoV4G
lpU7nshE1jPGpjGiHVXt+6p4uhqKIoVbefHDT6eQYLOFgquIRMSR9lF7AJUeQuV6ayDN06+jfwgT
XCk9vpzmzeKkZkhaIRM4mQpdi4G4x05kVF1Gpqxc1jdFPCTgvW6fHJOl1B8wng4GXFLKVBDqhugc
214HV4Ps9pVkwdPravOVNUkIHORNfFXl0+zzpGq7u08F5BWB3Zf24OVBHmzaxfZeDU+eHnbkyulj
255rG8p3aAvOrdODM9C7Mapjn5OAk/RLRkDjP6OJQdxMWNqL0znL3JVaa/Q1I9h09v/h9Revd2JH
Fzx4uIV8G/TMiTiWnOOklJLvE9ssLN5sbVTM2Jk2T1V0EisbVrt8QZbG3B6VQRzlTi1+e/lJRvSK
wKGhgrWxkbXymSummXhGB3nu+wZixz0t1OJkqgkZdGC5dpNj6XQSFCfpiGTrzRynlBc6BXKvLVq0
AOLhnFQmCQTYF4lZTC/POYQZLoTj8x5HLZYjF+JOqJvtF8fabhNTh/pT/SDv04uW4pPnxYdoq+7v
5/ym8KrV1RNYoiATLkK8Y4/bKPjAJA0GJGN0w6sRo63bKSYPqOq6bZXKaF82+izzraitcCABHe9Q
DK7//nRexppyhONNoZVVytcE2C9ScqkaZihX2IwcpynrU/6zmsDyWQQvGJg/jkP1qzqn9pTZKsCz
0OAqu1f85XpEDvyQU0w61JnrefNaGTk1fMFjAGqpktF6SwSPMCPtBnZwalga4GTE6udyfCkujMi2
pS2YTwCVpUezQbPkg+nqz2GSu3qjza4oVrs1NeWBz8Q/C5/O/T61yOmz/S7EWFrzDDuZCpR3Zsvc
bO9xLULTrmj3+C4Dx9mhlOVUfW1rWSgdUaBuW3fa0EccR0wswwGSuMaUIavuknO0dHUx8GEAdbYj
uLuhperXI3noApG56+ocf6MaJ/ZsXJJ9Y7OhU6WvnUhJjukR3ZEHIvdOuRpOyM3ZQdaNdFmipfev
wLeTCpKkT3AB5PRsE7optI2/iiIPQQMxEjfvaaS2mxj52WOdgaM3weZBAK+Q17/KdBc5a5BTQqH8
0cCbT/tOWE2bjj4IcHMwWfSlB/uPNednmN/cQVRCC80WRqtgHCIrJDWkCemWsFAW3RFzc64G4EV7
zEexcdhNp6/NwSnWv8zF73i/dueeLm43//Z455PUnlKQKXb6aT8NCR5i9jE8D6nH4hhKSM0AQ/gA
lugLWkSbTZHERj+9rkgwgfmN6Ddb5EbAMW6c3uIr7Mef7ma6pWeK6PGEtl0Zt2+SUoIpXKZ0lx68
Gm5s/NHzFIUUI4r0z97emL+3p++phNBtLTqIYthKAfLGtssZLc1W+oLDYdczWvD4wEN3J593FVei
nAZrda2CUH2rBzv6QVdkfOl68mwZVZO3N8C6XYqrpkGGw2TNumPj4gydLuKwYSyuuz3rKc1pEcMG
x+v3fCwrmwaks0qXrsB0Y9F3qRgoW80EwvXyKBTsWRkmIx+Sw1hdOeO/20SUXbHOB6OunJbfhTKS
jGVv+YsoGydqSWnhv2wTfIEE/PLwU/JN8VRO1PbtiuCMFzqAEu7Yfk2tZpwlFyPbc9oZLEvTMhE4
/82fgC2AZnijiWxodRj/AwOOdpctS85aaQhzUJLno8uaqUY1wSzP0ZYOWuWE+/EHCOTtWncPU59W
dSHYrLqmiEb2PbH5xoSxslGawSqdGf6jobNoAOJEgMNRD7+qebc4XybgtPcX++Dzl3x5E9o/TUzi
H2KSLl0rFklx4Wrmn3CEDtBQS6fU+jSpQckGQkf1sXrnJngOpv2jibidtl4djB23XuBBd/pAXaa5
V+5yBA0KsydgXnLohKW+c+OlVWE55xuchg6I79Kls/zZ15tIGCiAb0stGcmKpQ1ueD/JC3oruzgp
LpdqgTBvTuetLR8hZrsVoP/lR6VKsu+TRXFyHPc9GmX6YDnFAB/5rqmDH5Ix8CyQbckUXlXJaWHm
rILFengaiWwGdMfQmxQAvU9uPtE6+Jyw209+4nr7fUkNUgKrfDRsM2yiyRZ8tJWQroRqIxTjq0Jb
b9YpMqOOcOJuNKOK7aGSqNPlT8CDD+GktNyDdJGkMQfrXL1hZJVGpTOMIjAPuWFqly1pv5qkoP2n
rB8A32Dkm8jHrhIj44KgFOQXR9s8oXmlBp69x4pAgX0338OEgenRQY2GfC2SKIfUGxfKL6DPZ7sp
xahS/R9apgzKGQU0LktyhhO0wWdAa89KC2cf2GKqfGWow9Bx1fDXby33R0nrSwcYkRFfGU+BLKBr
XHaxTiuhpfVXQrB67taQOVj6xfY2kq4iIllXkrKNlI/FSsBP0zbRYwv3/1CSOXiOmuPmRc2ZdnLk
IYl++HTY2eU0lBUu0yMU6aXnMx2wm42bK+JEpdzQVcdeIDfGPT4qGFlxv71DaWfqso56DQ1deDAs
HEUpFnt6ZVDb38y2Uesq+3xSyDUVym+DO3mqg1tPXDe78E/x2KMWE4JJGFqsWgAEI0Z9Eg1wXurA
7zCn/JgbK2kRW7fKUNApO/SjyGUwIaaRmUnn2NVKg+R3x/5lN9NPPnGPyUGxgqVWx43jYqc0KIDi
bScyouON/Hor72ML/cqgBDS5hoAOZsnQtRWIRhOvWZ38bOuP2aZ6ksh7uC5U7zUmFmw0C1O7ZQH7
qCodSxjezUYfUaG0VJJeCI3t4luFVybI3uUW5Pu7ea5qhK+EBJ4OabEXeLexJ88RipndPBZ6e112
Hec3MgquOlBEezy4rP2P4zxPcHK1/9YKqAdVNIdxNNoyUNOxWPIosYD1etfz01KDmKj900DzouTT
mAD5gYe/etGlqPzFOOyI3GdLb98F6HIE86Ypl5gHW2tdwSIaWLDAsWpigi9GxlDK3Olk0SM8HBxW
9KGxq/VZQHM1lYinQphITj5sR2oAUJ2x1FQ0YPv7Ck90rajnwtvGNYXJVsNDVoK9c0mH44qxPAuo
QVfjxsYMjJzAEULcTWarO5N1lzMde47gQ5/pMrhSjonZB2kPvO8OSTdmiApkaqMp/ZLpo62LkW4w
/3diu0S2qLlvD7qfwKUWWjo964JSeWKzqoojreMSDbPDW2Iv8O/6kviNE0dutzoLfls+8KDfxqAD
3iD6WXffODeiwIexX7lUNvg53Qu6ExhDaiyujMa+OtlYmyQfZOmLB8CS98F/Zl0HU8TnsCGppZXo
5iOlT+MyyQlr+QQav7s9QQCBHTqE+4w6OSppakPFJYSd5VDRhoDa44t9gly8YMQy7x9rKmVvPfsh
gFwGW2gYI6LPtYYZx6/jyvI53PJjQqH4cxs4q500Y+zO9Hp0QhVDYI0qzvbm1F0VV0+Bnp/y0sdf
J0Z9tWTUrveJoWEqFovqSBxybjX9JkxzCaHTEcLYwhCeSAOdzR2eQPi0CeKj1NgbgXNVjBBXyu/q
g1JRhntfw+y3WtG3O6zZk8ggshr42MOCKhsHDvcKMNg3BpQSQLipheloOzVtN/BIdgf1vPfGg9g5
bfIDVKa8i20AHMzEqgXUis7y3nNQ6gnIdmjFa2xQfbZaA3boiWG/OHBPfe7J6Y1DXgqJIRXzHN29
KtrHySwzWfuZG7QZrbx27X4krdEu4YO9eQ+Q+3j1nP8+5b9au/LqMlGJwaz71FHPk0SaXvgeNPNu
N9ZfPQyImknStImudvnQ4/F91qsZcniO2QLbUhLA3SnZ/vpWcnOCXCWoa1x0GbQvC+LHwgvYxcEy
ALkpfvVTkGacCFaESV783UcvRDYgnYZPmu/tyf3laAib7obX40heJ8EJqauJXY2S98K5qj/ty2XI
eM3FyVzhIBB3/xq7iyz0t3n8a74ElnZg+26om34sGHmFhynvy/bUFY2I92dpcwccyW/KehozJmhQ
CNnXTrnRwKF2ogGGjZvig/KKO3fhnqG8UfbqMw5knhBwrWrydvgw3SUkDD2wmFShu8qtxibH9aNf
+7u2iOmRQxKqn+CqlDgD+oXRxCJXQvC+9lwsttyoc9jKNqIMZ+2MhRiV5scEuRK8fi/iaeX0X78D
AVheD69bgTHc4dj26YOGu84sDIr/50Q1Lq9nYdPLi7rVRwgkE8Fd41CSjvlanHHGlCOEacDZvhP8
OWyvci4hoWKv6bpGWNie7aAghDoxiLjd6By8ofzCg2VpU8LbK2ruvDhfBXveqT0B6E8w99PfvX/Q
c/d1pHIP1DDiD7gY5EdMgXnirsS+g0/lAg/mysCMzwse7L3wNq1MPhypdjZyZ2iStQWKb6LK4a56
bm7UyeVQpTrpbe0++cpXeIm+E6Mdo1CPY5dkwKEwOU5e3akicflJ6NK6m2xRzrpL7seYe4LdtYRq
xDKEpJUbM80FjX6qmTJljgfn9Vt1PT4i/doEn6z7udGWncNH7zexYRCAe69rUTEOsNFg9/V5umZw
doHABzG6+/6BcB3VgrP0JCqpURpHoXiz2dttbfdT7JosH9NW6vtVgNlmNUFxd1JhVsG2y9hL2iIQ
MBBIQms47OJ18ik44GCCyE9c3aTDFZ7xArCbb9OUydu66vDIwzdqOaD4IT6/b76si5+lXNE8FaUU
Ts+gXOxti5cDAutgMdWeemEl2zChbBci2vnjyExuDCN9XT6GBLG38Hmbcg7jVZ4u39qVww81meAd
Cnhw+ezf0uDG581pnwOFapIi+RkELpdWjOHAkTNXGBetDXMIN7QfyQWPjxOkh40x/PS8k7fLynG/
zCcuDwysXkidRPxLbz+lYEf913DSdY+55mgMsi0+KeP9xIJTF9gzmXKOmL28gx0TkKon97FvI6NI
ZJbKQJKMprJsm1OOXWw7O+coXphNyNch4tf30o7PSBMiAqr1097InREo0h4BZ4+2FvYUe0zzPuAc
koDKxhk7T7b30501ngknkKUiJlacROmTuuRTUdeOII9ro7Bxd6g+guf67/BYXf6bn3bI2ryFx5n6
G375Be6P/OggcPAdc1u4krSndlDcBmlmL10l0O86vMwIePjTBT/IqUlc0rdyvhpdJahBDJ2BNZLM
+mrg5RnRsKs3fO7WUXpie9FuB+DwiluLpOqNrbEHyYazI5SYG6R7F0hGD8nFzyGd1ejwfZZheQme
gIlZd+rFTcHETWh67XyeArk/+4Zg2NeKA14+EnpssZDj44byKS+5OQFFrviA2xwGa3ICwJB2CVFh
JEAEiunt5BnyT++eO179vywJEesVYzk9h/ck1cz1HFXfmG3cDnWM8Y3GkfUdMWBPfFwRiXUdrV58
vFi39xi54oPeK90ZMVOP/dxx3qp/y4yOZ+Fx5UaS7iWCfNFnWKghErazfLLJIZssDa9f6wx0c5qj
fpYJwO1nXCugD9a5UE5FZLltn7Ygzh0HVQG1Q7FyAZd85QUs0Io/CmDm3xmPUfJ+ppThggPrhiyF
aoxpAh4dF/C0PuocRbF3/WQILta5PVvvckmgJeQQUewXoQijeq2MyU9GDf7KsBD5J/nJt9DirblF
d34MVyV48Ahd/AXxz6PXV1RWl/0ILdMpeonxuiNfu3P8zOmxWB7I6FSzjtqaWqk0WnFKrvK9bGhs
KbEc0jqUWu5TlJWwq8q8/EsZHAmkjThxvDizpsNHB9ppThvr7dnzOE1YNGzFr8iuFRK2m5EY7KWB
YiU8o8LQfIKThLHBIF8qj2bPPw0DIv4GVBsqr+7qE7no13E7C2C0QZVXgpQsUmXjfDk0WsOELzIF
oR/j2A0f8FTApNuFEY7oDYeeB3W1yQ0bs4+onoVf7buKMiczCiStA2ObEkAAJ7tFWL4wxtDohqV0
36G1ZYuiVFusz+rldfpU2ZHLFEsiOyvDnw6vXk7+z6l2WHwIs2+0jnaTWcBnEbt6nxtZEHxDBSB4
kXtcsaMj+G9lGjP6ZJb26JYHi1Wl9vORDRFzKDw/dTvPguH76lubSzOVM/9J8/5FZWEriE9CYJ+F
bSF9cuWz1rGWdjaHdECVjs2IS4eaD/pT7/gy2nYeRw1KLuZljeg1F71H/b5c4GMItuGonChUvWf/
lJLaXPpWbu/MgiEcTe5kFRdXtYmZqx4Z87vaG/jJ711pU9El5beuD5frfGg4e5qcRJGyFrs+KsAM
BS9PCPrWTItghBK1EWBlPPZz+VJvSHMDfHgu8LeIIag6z2kKu9eSEhOvlYzjUlUzkkrW8t45ddLp
3uVrFSdcqUb4bgqOEz4kwNvBNzgEsApNilCqhHtpzqOr/s8WhvoouDXHRlAlcd8Ctjf8rpgVm5G+
N4TBhbF3y9suCRRX4egNS22RpfhSnISBTDxWHAIGnetIayDgI6IZTtL4NFgTsSeDncPIb1iw3s9/
b23ZdOsEnxl+mPLkHXGG5xpkeLnn5jKBO9GyUuLCL8d1iRW3wME/aladArGbs1X9xMXGabctEZbg
wpwkrqXJl9hfmFn2FNRUrEcFE8oR/Qf2OxraJ5ZyDZheD9Vw+gZbFmcVvb7blGX8J6RxA2AQ4h3N
v+sVRXrarbpP3tfpxCw2z1h6QNy7JwuyphrkncZWtkWCqMjrIGlKp/OG3SVouCab/tPpAyODXTJj
4iEvPxMDLvyj+n9CKbGVvxyF160yCr1a7ns/4tSKdqzX05QEWKLp6iflvtRLZFJgm//oxS38JcHj
CGvY40o+Y0gODxB1fIEwV83N6R4xN0xawrD7bsWtwzNly7OEucqzDcnIPrEViXMUuVhdbZHpNHgu
uYmML1AFSG6Ydrh2mDF4AI93AAVFx2dbOEpiJGf7Lo9JWr8l2C0wR1Glgsm2BkQ2bRzBjd32+c+M
S9O/MELqytgFn1MejrH/YG9/SeOCHdv9fo3PdjKdUERaCmSfdsaiqccmbKhWssOYA2dX+0YRLTgm
5CJBS37MIC6yiA/GlbxNMcIJDneo4qnpt2l2iJjAisxyq3a7jBxBORuPTjGk5q4aQpuRV8oxXAjY
FKFBUGWhJjXC43nZEumXcUI3CGNM6RYDl4OcSl/yODhItbH6IiNwA6nYsPaOX084TNjbSw/H7A2Q
elBI0Eo4Q/YtodP5byh7rWfSWCy1mwRZU2pCvqGD+7io3wQ47Rgpp8Q6b2dKwMuNI21wpF5gnUfM
Utnputk76dHR25bTjM7X3WMGMvJz3XlZ9GP5PU2B+gCxf+f8PjeupiFh1/IpxeU3DFFxjxlr6OwJ
2P3TBF7PFIfVS818y3z5/MOj2w8PL866sF3pcgtFuq0jXaRDHowR9LOt9GjZNEGys3EhIe38XOl4
NZOxr5uVq1k2L8ex9LUKs1hta3x4QrwOOacGAHCPKTcSSYXkO11zMQtj8oy3Mf909a0Wn0KNMPTb
bvsBGW3PIMbDCnzp3G8I+28O2Ch7LGxpVVBWSY4ahgw+LzS0xR8zF5W6LPyDbjVLgYAKnHmJQggF
jexK0BPmHa9FY9IFNO1yDc3fJUxCSqifdKUHdhtL7mglcTGiGyJ3xAujpv13znpCaaWse6ck9hew
Mqw8zj7gucdAp3uOC+PaDL4PPVOjYRLXTOvvoL6Qga6oKb/N181becy2HqDkz3C0g0eZd1/ZGqnx
KwDH/f5np/5c4zMcs8FbzHYS0daUS1ujTyg3m6lpbUvyKaqE0LZyutJpSCB743NwNngYLnWWSBbh
mEJ3Z3hLV+wAQT2SDrutl6OftuAe51IGKREX/feyYwKGNCOeKI2n/Dv4cjCNs30qDMCr0CSZbgEF
bz2caMsATURbBfp6Dz+WfEt2oJ+t99QIS1Y3WG5mLqSeXI0LFt1dYgAKjJs5s2IbF8bS66UH9ah8
YBQKw85yGTimqeahxK67SaDVps4Me/e2V1K3ZJhbkJPrJiITwzGbBb0cg5OOfkNNjyZQU/KDVxDZ
Vp1jZLFDNzzZy3uSfHGR1MBGKvLCbVI4GTBCImVZQ98FTsgsQjVNs05KrCSSq+QTyCCJLTZhxi1i
tPM62hC7lMacl66p8vdVkIjgf/jYCgpyl3tvYCXV8ObZtzX2eYwpO7xo9kLbCAwkbL9hYG/mvMR5
G8IB1Dw513+5ZSWMtRrg0yNKLDNaB/jEUE3iHKYbAOBskBO8MMFeF1EP8ehwsQwcu+ebM7FbULHj
EfCE33IVUHSaoMeCRVSFxTI1yKB1A+59lbTXiUJAkLgb+XqLm0EjoPhd3Cko+diU46lRJoBrcpRI
QstBfronwMM5abNlNbgQMSAZCeZ5R9/gC3JjgGaGdpdhT5tPDSUtt2UCJ26gk2LdPLVsiKX1R1mN
JlWB4F7ogNIjIo0Ezd7L/uuk50OuMJ2urW8KLfM+5jJN1RU98FLkkHc71GoxJgm6WGRJuDmmTvpz
J8AfTmOY3ufOmglmEQcBQCl+R1Rd37u2+cYxZRPDis1d1jIEFPcfph5qwVjLWXtgeNJSTKSSJeB3
c/V+PJT4dMMwAX0bbsX4ou6wXCjxPk49uEfbZsZMOzvi3ABhAHjXTf/0d1sm7gJJbYG+egbBOXOj
5NVjUmjgiA/71O+AXALy88NxOQe5GL3fy1UHq5ZW+ml/SHB0kTmZFRIbFwUBcq0L/dBW0yUQKblm
r+Surs7G+zywUTOFn0Zbk1QVsyLMSVX5+kYPzff0gV2V3m+TRAq7mOH4fFBJnPpi2iEJRNHOAvoB
GhQOv609wPm+aHN3x1lXTFJCyKP3P3LcF0KNpxbdovp0dASgPJ1begMSbpSrgLG6sj9WHnSS7WcD
kaT5JwrnUZJP6PYP/HrSrehq58yquC4ysXGdVLqh2H4ilj4an02YNb2KhhmHtOMa65hi1dVxWTnq
Py9lkn35MKV5DAxpt486q99qubFV+p4YqcRmXVIhZZ4Qw73LjrRkFyxDWnRV/FTK7T1/5ah+82Xs
VG4zbsqVeuod08dS5zyqMDvufEV488w5zkxupckYZ0LwMaYAjJ3MQe1GLhk7v0iI6h5rnjsegIDp
PSUMIMUV+8LzpY0Mx5qwy9X0TnGwRudgQtU6w4hXQSkjR7umpuZ3uX9z2dZia4oFALmP2RqciWpK
v1F9sf2BBUet8cK4vjxSNmcxhw54jqR7OEvVVFZVYkQ0gem9jgSGiwDwcaDh+SzVjTih+2KKZwYl
XWyyaMSBVAq6FHt9jLDVYYcr46gIOsuQYMAaYzVI7mGH8BYIgXoeExWugAv6S29kjA36yH19vuG3
F4Mt8b6v0KvZTfWvCPqxPRuCeIjoRj7RpJ6CHFMQ4QasSj5O9VIkHhsf/6gRKtWArmAQdK+iy2Zo
oJFji/c9MeHlKdq/POajr+Oc/rsp5vH2GGxKpiWTTFkQQvrSDTCk0cD9i/EVRl+9L8CdkLiXXgiG
9JIHtLZGcGcwYLvgW+hM0hvhTw6iZMV76Udv4irc71hIbMvwhVzfy0YEyr/jX5C/C5HIT1S+q9kX
spEjXVNsMaWSjQv+mpCf7gF42SzyZtEhuLnnKbR6CiF/ZFR+VwLj/muAx5v5tSZodH3sMwvBP7hv
XS59xwUVwz9dENo9vhVDGKjeluIybt6BWN97sO10YpQucoTQJNjWUNJFc9MmtvmI6rYH5q+O/H9u
4umquSOqsodwbsn27/L5ldPEfLZvMfX3gfkmO2cgPHLfyeN3Y62dPSlY9XMOoOYgJfJ4NRyvTpq7
HbwQMaILrSGhNfu2fCbQOJFrve5tbGFHdhLm25YUtJg4rWT+Gu+5EkoL8jC2u1Wbx86UDz9fdPFt
LtqaV2ShGIQGqKRwnD3gBxvFD82KZsCLvbLgcRKfousSbRGAu+shHoq4FC62K1BvcvBQqFu35syP
Lo0WYg7X3VkJ12kWJBrLu8781+MPCwTwTXuhoVIseEmYGsYXAbHeR6Nz5eGjEDXPNE4WF1ESljOS
mTmBYy+egogWHe8OLggmGC/2XrhmdcTnzWbLf+yOQV/xx4AI73JXvn9BNzYj7nA0aqR0wjW7dAPj
DT56UpclPPHQrjI14tYNmrzO5gLFd7wtvzxaSDyNCRKBMpepNnTEg1/Kdb3nMXYgpY6TSt2GaFxF
0zSi24FdADYd5nPUfxrpOUHSfEArKsR5VWHDw/wsAWLpggIVXDpgoQxQrJP+GWT67j0zmGcR1Ku/
uf6I4kCBrg41XWqRPgfHD0VzbCwtfFtj5HkqSvR1g20Mh72/lg6EhX7iy62udFkc674mltge6q8T
qlIYxCoqF2H4t/MlA2EcaYBGmK0k4NeYhZw1hwKZMs3owLyuNW4atbKCIJ6lLCcOtWyYscBXfuD3
MXMmfHip1/Z5XtMlpr9f4h1c2R8hEqdNxzmatzbe7DWPXjennvWdp/sar7I5mRUdwaSTr+ywLhc5
sM6CwYj6r1dnEOQWM+VKxmzbET7G/1Eg8ZvFPFcv8DiWKI3g68qeCnvxv2co6arXEk6ZwooTvkaS
rr13p8bS+Supve/50KgT9hE0tMdpNVpLF8nnI9SZXj+OQmcxhOknZdwe9/+3LD5qIdWvOH5zou/K
8HEpOqno0kgnJ8wmbiCAajaxUglsmiGTe7pz27tvCpZrY1k6zT/iFXzXhKNoABDo8tG1HxZoHuMd
RHfVoxf00RHmF1ZOHu2C1mk49+MZ1b9nHkzVfXpgGxIdz69+pzWRTYREDN4VRujiZdkOe4HBgekk
/zZ3z7cn6lWnv+SmhWywQ3WI2MuS8E5MEjUyOT7h/v7KB0SVV5gf0U5zo+mMjmZRF4oHTv77jMsi
Dyl1yNuDs142kkTI3cI9UfuodCYcuUXxZhkrdlZYRwTj/63gpmvLmqbZaR79r3RLy0YX0HJHHFqr
Ll7Fs8vB7bfUfx8OXn6V/eZemNLASh0E7hfYWRqpsOb4aa60aPqc9l+ZEEdCXUpSaxegnyCNTBUQ
ontXgZsSnvy937Wpl5I7OoeMNgSEfiP31zUY0ELuXqlhgOWlGA/9gqt6x8EOLUFBCzjncMPk2caZ
xwFfRAt/ty2UOQTQBFCRA+9J8yyHCfQREgAKB/kAriQ3zS0EFdcE110/kcruHm9RFk9GZalGLO//
fVsNSSWYoLSxCnJkzaPZnKo4qqA8hLNXI4qazXvebnfHG44fM9kFsR5pV84sbRj44vNBH6Bt54CI
Iqp5CauKttpep1bjBAIwsK5NylNfAmeaSP86SYjDgT/bsX5ErrUi1mVxHdmCyn4g+ZcbCwMz1A4v
SQ6M1khGNhrbgBo0vNdsey4zwF+fs9tL2jTP7XALTLk+tMyRfLOzzZZPKJzR43hdhL6aFSHMXGot
AyjH5WckVXAI76hn85jWb/eMnVOF5kgc78quOkAZW/+s98gVQN4afc11JL+lBZOer+9ZOu5pKkwx
wW26D1MhIa6448I767IVN3tjurWSE8ji6Zn/fNHNKtkqOtz8OlXUX4MyLHwpmqyIJtW6Po5DuO7a
Bp+13rIoe6dP0iijl9rkiG1xnL43LVKd/CMf6pGspICebDXxr1jyroGLPJswbVSQ+Rg2Gwryp3bp
4zc/xq2pykETlASgYZDRJjYmEwJtB5AjIeK0JcDMt2VZFLYBpoou4ZNBRf+mA+uucblgNjB2c+9P
hdIrfgLMjM8uulQPL4RuR6nzHlbhoNol0UXaPUQLY8IKdfy+OVz0R+KeQT3TE2JNkS0RpQRnoR5v
qDeemDKOV03a3IRa3+a7y7oXeJNfaLfwnzkIxixbyxvZ7pNYgCuYq0xx3XUUaA88iZIMX69hUb7G
qQMEYO2FxaxHvqD8CxYXXirYKPf+tasZGVY5vIlPC0rCL4WfN7xXuk+teh9x9SkqAXnN93OeGAOp
b3l3AcwF/CB0ncHU6yoJoMeN1GC2wOrBPRFlECM2rXKnBE5S72QYivv+RNYQnGCAeLJiAvGKEt6U
2TG57ijexMCdpSlWqyzZ5gY9AcJYIVXkcitSlfNPMYp/o/BJfZJ16jwJcTRWGnN0aiCGrUj6pCMF
uSCi91d+Qfo+9wRxH9T6fPRY4E0IwjYJx7tqqExRASTESQ4OnnJlH3yK9g2KlU+qfOYgdCoJ/A3x
ygu8wNWexaqUbpHToYjQrgakCB12vPD2yHBA8ouMvcAsSWfUZJP8HCF83zu9F98H5+IQVZPQENQF
Jcndh1HYJ6hC1AG4pFFzBtYtVmYIt1yci7YMK7u/fEoOpLHs6OUUca/eYkAVQJaZpQdaTopy0F8f
oJQ2h3UHrZCFIMAorAyfg1Iz5DuaAj2UtXAHPUVUDUDfqGW5XzPX4KpekSTmJVVy6pXjEdzdjqau
6myb7o3UKpisHt2kpt9v/Be2lO1jmP4wse47BhgXUaKn511/t2bCjUCFIBSzKEtPpZRdtK4RRkf0
IEKp8mcpb1FLr3gX0eNefl42te6h1nm0OD1LNK4FjYzD+NzryTIPOXfnWszHzUZ9KGuazzz/ScmX
ax6MFKV2LesR9EIPN7ZP3CrMwvwj4GtV1ifYbY5PMvzR0ZcEM6XcBBkw7XpP3S13vRZyvyPDoXcq
oGB77FcsC8A2KbiiB3FNybPTQPuqajp+UJ0sAm6xRKuoXiup/y7p2fGVuG+h5NWrbMJ0K2SVU9fS
tI7RydvzMv2ROX5fak+b/WvNnlbyn/bzP9oSvbz5dSzI9GH/lwut83sQh59vVEvAfSTdTDG5fJRS
tKzOSVbGBUfOHIA3Vil11lyCdMqnZwP8jZZTn++biM1qId/p4DTvdAYRvS4qk+vBohqyghKm2qU6
RKIr2iOkgAUoXpp14gKFa1k5UsMbEQO8Hxl8V1/ZBOmJQbOkpMknxIAfQdRtuRxv+ZBrEzKbk9Me
C5yNV7tw6Ae1jFONiNxaqlShM3nHjOAKawXngxdEkL57XC3fYsUDrEb0cgEFECY/B0/eH36EUqR4
SlfunWcLAckXIiBJ+hdrBJRV8TecMuenh5xxWhSR+itifXKacrobn3ba3bRCgcW4KxWJolXAmv+d
/cDyAlAyqGhp87u2a75xUREpwgQW+fwwpuB5e4vcC5pGhPErhmCBKoM298dBmDUXdpV6jrmH/GKb
Nckat8u8eFA+IqbGSnV35i+LBBq8MHoiTrygcKCd2Lt7VdBa6C32AUU7t4v3KahJjTwZ2VgwX5Jv
h9dyWXvGG/x4XTohLEzawmdLVVRg2CzQ4KAsByMvJJurJWx5rt0HgwGcmAIScf+xmvlkiutfh7eh
1MW22U+UJ7tkEcCaeDH6xOqsAMv85VYmAnnUPn+jFEszGXekS/hiMnf1ARo7gqygcSdTsUr+UUEQ
Ff3gtYfTl8MQgFJbFvOOSxlMVWFu01WFvfDE7Bhz9P9MAM4ahahhHuLojEwehSyAisd0PnMxyged
cIa474ZRJlTzCeWI1euT+j2WE/RDaXFJt+aF2RmbOqJTTZFX5vZ7LAOcfq5pmgV5c22kYQMY6Si3
n9KRCwJBVM2GUUKrbXBvtgDfoABXciQ+Ps09p7tm4bL2SAQKv4qtRppj7gVrcolKjw8PMa+Xfyq2
rVJ2in/v7iLEFKR4ICn6MQTnE0oNW/FtLl5Of73X+42r8TtFVbltMRehU/tPOFXgXnzkKt547k7V
uM66NEoewkgutHAV98+PUpI92eGDch7420aR4YebN69piqd7JSQC5EWkViMo3ZZrG44sd9BHF5WR
OjzCazJINV/k9i+4aejF4kE729K12vpIswbMEQnPuUslnvU473ZJDeFQ8q73MMI7dr1Wcsg8mxS0
cQXxOFVqye7jmSNwjR2OzhXICmHAWJcmL9eUNP2yGHKvms7G7EdKmK3GAokr4BanWfO965IBSU+x
Gm7tOpgfnfzzS6njVGoLeC5Q6/K391XQNI8TbLV+DHjeF0QYvX54Fif7r9+X+MR4NRNHpTUY8hMN
nmpr1Xz/W49/nZu1tZiDVkYaRhaO918SUBCY4OUsPS/zPgo0QH9shdX06TtIHKR0UX0W3Uk9kkyt
Xozcblbwk3vN+U0OdPdkMYbOoZN5Uy9pC+IgeryuXWxU03f4NuID/tsndjf122Ub6fxIaKlmEthy
2I8PT+UZfDu3Tku82f+Aow/nGWPoSdKpwxfzaRF+WMH+B1GlUDH8lxoo/ArofwjVpGTjlenpjbSX
BOaaxKunDd4kHDL/v0raOaCjuN+Vvo2+Svx/7H5VQ/jxTr847Al3TUUQavCva29E+dF82gs88SBc
CXOWIZ2U+6ub81EcZ0uuj95EOY4HQOBElPYOm0n2onJM/9jhS/gWubcJljKnEaYRojLg0BmzQNEM
Q8eUcm4MimjlGHVTjt0dNVO9TbyxDoXPuWeu1cRLG6vhr0sDLtSzkn9vAkSL+5+s+fwgt7+8bwji
jVs/l2Or84T0z6AfwtpPt7XiM9vDIkUCSpyhy4YlJAE55/ye5X4PqTFaGuY9BHo5klLfaR/917mi
i04SJ/ZNRb87EE1pTUfZXFwXTovZBE2hV9uG5v53xsWgDAJdGyzv3FcO+52yYN6dGOeLi6xtJ6XD
TZv49oA6U8XA0OW+6OJOkzT7bpaZp9vopMLqjW/IKOQ/14W6wI+E4L41hPjxpElMnLvBUAKmaaHh
5VZxZUpCMi2+VARPoMEoEIs686NhRxdGtbtqKgMIcJzVQdvrVFQ09I81hiGK9YKIhQwH8robJzXK
O8J5Amh73jPsqCcD9L1+oVEIa8tGYRt77Czj01j4aCM4RCxwieVXTZbHcS4fTptWZpGR9mMa/aQX
+DUuUZKgDhJirJnqszBzb8DuqyBw6Yn7f/m1sU4Ut3bpN072qYmIGV6dbxUDP5SFj/kR6zTrhSF5
VSqajNgSsDrWMQToPA99Z5K6ZPfE04IZM7qWPQrIXEPf/nAnVWZi5AKhehHpLYi2cE5dk6rhASeY
7hQYKsb+aBHNCtGUGe0OWx2kItyEg6FvZuPuhJXOIvaIRJL+6dMuIhmacindoXZ0hLCcbxiSAcYV
isPgnosr0V1V9eoOtLkrcZ857qSIwGWoe3ClbF8OQSsty1+H1kgilbXGJqEiZsfYZlfBEFMrQdML
dgrIsuDcsOrPqdWifKvtuSAyZmXXpbxovpn1kakJYvdJDUl2hOdpoiITrluYtGesmIi6nh2ocnQe
rnCL1OyL8lwLOByTkHA30HX+go5BwBJs9CdB0uQlpaKS/V/tKIq5sQ6L25i38yE/1fNCjP/fSluF
f2eUk2h4oe7amqF8kKwJT2IGgD2DCEDus5rrFz0V7ZA9RM4G+CIIct5HYW0Eqgjc7BB56sGLzRXm
u9JfaJNr8cj+xn3MgGb4LyMG0LP0aKYvS1jUOh3mZjXxAEiPKO4Po+m2LwFGNm1hueF++SQCfVUw
9Z4eG4xYR7+x662Uz+K+tKrnz5g64wCeNJJXqS9CkINuQKmQ9XNE8qhDp2YY2//EsgDCL/8rzytM
6+7JUMF26hjeZnK0tWxyHuF39yQXrWuO3LxobtwcndKtymQj/G0Ui/5MXlN3tjM/kOS7O+Hl/xht
wu1eL98t+QrGDrATQGpFopPbLm6EISrxzKeRSKkTiU2Kw1LXFNuSzFTcY4iHWHZI6MgVhQr2+rta
HLNSnTbyVZCNJ/CBtUmgOXWXbUTUYLdSNP+bUzyH05To7tKBvfNaDZ48h7p5PnZFnhuyqoY9sErz
VEuaISXNUkkHebL5K8vWO7InNwejRulsJpVZQV6Dr8ssPBnJoJMVLwcZlRCJwdnsjRn09jUtmkOX
EDo1BjuB5s6JjMKDE0Uvj+DytmDJk4c5BQ2VMDR5OeFdU/nnCyvtN1gCV3oSm8u2xgrAgJp1Vd2Z
VVf/Uw9NGyFz9kxnAcdWELh7fPZqtbQ3UwNvattGWa+VnYwCIkIyE1/kXvxNhmiEsMId1MSPtxCq
KSza4NK9idREXPc9uW4Z44uhUb50Kzor0yknuDFaN65uBCXC6Ufs1Dru7/rO/XuPnBWRZ42/5gqf
jQ2mN/5fUy7Hmqrsl2jHOTK5+NP6s1o/EHKMFZH0DmMZAzNZ8fo0judU3oFwd9Iyb66ib5Dt9V7h
HsGaeOPBpc7HdJe7fs6/NbGZypNvMUKgN8oFSsXdytIaDwBdviLNo9G7H+yGyPF1e8PYaxQbNlO3
WTEce/w9PnBMvTG+n3CQ7unSW4q400KV7Lm+Kdj80dj1Jh86bqlhTiwEgGCAu9nlkb8aV4rxQlYE
ijA3I5XH5UkEf67JTbMLKQNL9ErfKUfH19NL6pQSXFkvkHWmxCP09BKrnk0SvuiEtMYPs3s8XSsa
ga5OiqIQgkXaUVyK1+q2aItpFGqgjm7mcyp3uaVfVSd0ON1o0Gs1bN/4jyA+QbYef71AxwoYHXth
mv1ctE6aTi52Zjxfnb/s6zbiH2NnIf+lEPcDZZleyjQ2jadgjMtX8GPQVKxj9Cb9/8HBZZ4FKBTz
Vq6ImZRzw/vJBE8pLk3mJtm8yuPCctsMPphjpme5eXY3p3bSPRNwR14ObXr5qRtOeUmQeitCrDQ4
bKmgqDsaYUZB5ylLn3TI128sSe4rTbqErESXI2upIx5U7D5xSiyUprf1Z6UYEk5W8757tfqNHsco
2qzTuH0ZpSrD2U2ZM3NRw1wUH9dYomgVp6JTcF2ED7Q3UM89NsmI0boCXZQe5bYEvFgM3WYe0oUV
bUWb4HNzgI7kvFIvrB8m2Xgz+JjFBf+p3UemWG0eFjl46SsTLPxeIOTvXXKc+JHKTGIoFDLoeqcK
QLKFqw4A2LlbVgvuhgWvCLwR2Hd40L2jwNb3WUYDvrH7TP5DPZsUstErSVGSPQh8mmDauJon+0dw
wrrEepPcpQl5R8wHH3TDWs0nvwI1mcZqADbfSoeArYpg6iGBw6Y20cKcF9DSokg/XvyTCnv18lhB
ZhuclUftygd6Rvhgs3ETukmXD9BkHzRRtC+/XtLkUdki2vEwcA4rzpk17PK5TxYOsLtsAaxeeuLp
+EMx66HJ7U9G/RZyYvQRYgC97vEcY03uv4qVcecvocTLe0BFnevE8u58ry/isPrv0fa3t+F6ZRXT
irYAN47SfehRmjhWPAn2AFTRO4tcuX0VUcaBTqgKxf8yVYa2xkbZSWQ7Ppks5Lk8Rq854anx+Gql
3sSGwBoLdjQeD/GdWqHe//vVeLjLKB/3IN+86592IbyQGie8cXRX89D5fUXgEHzaicIADynbe4YF
YHsa9z9pZPQSiF0JX9yPPRoVnEJuYU1Gzmz/CPefl0fuPOgHBXDHYeQ3NuWWOkEe7F6YW5VYN7mj
jyz0a2w6t+OhXtmp7GMflB+MfxVeeZOSIWnFI0NzxnNtmYL9FkH5yUZrdCyiDsCvcGpyhF8j6Ort
5yY355pzBfe7xyeHW/u5Ipt5/+gXbVYqurbdSiecMVKW0PATGcQ6vrh9+06uYIChe1S8eUAQa5WY
SEduHT48lpkhaMEkveN1hi0CJxJRM3qwm4mLgqfzUKQbZQbmxDl4xUyX0s4YGwAxz/z6zbaUZkmD
vZh3GrIFKrNhjA8ztEhiyUoUFTc508bQYon49bMJ87vuZqD8zG0xXG/AzupBMtPhnr2VBdxkOWAt
Zz+q8qbdzuReovXuyGOK8wO+UJft0MmpqYVrsa1AW+b5qPBwXs9Gh0Wvt8FbrxDShVOFFn7NdsNT
MPk8CrDtwZfOqJDixbvdqCGVtM3pgVvcfB1TOccnmRm0Oru8LXKTivIPQbbxYXdQRKgqaZKtdz+J
+ZU0Gv5CVodpvOB41wBhfPRmezishPGwJUUylHvKCCm2epwE5ZdljfZKxQHg3ZuBCVZcNImjQj90
vpCd0Da5mTLE/t6K6t/lEzOWIaOqJkpNFAyhj4nMNAmfJU/AdXGlaOiq2ma8ih4i5JJ43lbLvSxO
bC1O+zM6XR+77JzqnXJK7n16IWLlJOwA+9AX3bsyiShxmyYKDAtRtgCmGr9ylcV1HBRXiOgdnCip
5buDER1XcUzMPv3yBzDW3a5MKvlJNbRuVbBPixdN2g4HZnfHrZ38g/vy7LrEb9PgrnPjrS0V5vtR
xyVMaitZSjubq6MWTVclOUtwH4XHvv70566XobFaEv5nzXeZVZiA5lcs/w9xO6ihwj/cSgTcLLSK
ZXcK9EyiOruqf95OIDGN3P5VsdiJnRZvlKY1iapMW5t2DTRIHVwOu816nYDs6+acSWaBiEK/0rD8
HOEnBbOqFPhxWjgXweQ4/rKLE9h0I7nnfk0YTc1jsiPdpgeO+bQ1/nYBncEIXd7TFwswoilk01PQ
M0N6jJ6O++EsatF9I4SdlXmPB+pFBGxMMpFRmJ5p34v5u9UyO4p5W+PilOuXKIejMVgOOAyJWxqh
hOtKzaubESYDrLmdXy8pYpoKNuscb5y7yJSOVf5hsQzlfJplNvp8V/f28HzXni9K6JCqvgZw8QwU
CMr/byT4chGxPjnQuFMhCPNNLyqtKfbjFFstvwad+janYgz+PgMVtNHGJquE5cQD3/hNvk3UK4WF
5849N3J7B5j2cbCEj2tZDJR6pluDAqcfCUR6j1t5TPTXPmiH0XE998/XoCNVF7mvD0TGEVPYK9SU
Efo7eTtM9SSs9V+nputZBhO7z4w12DHp2y8iwhP78+roSqTHYYGu37MnIfKFQfqS4gjgtU15E5oT
4TtRWKsKSWdNAIwXKKusCSD3KhH5benM2Oxpge1sXsr4ySnI3k+PBDqWV7bC18je+lQW0ajx7ctf
nwsA/C4yY9BogvAbke/9nlL4dSulSs9cARJnh3gkqApMM3+mMAb9iXZHqDpoJFdsq2Ef5No8YgnE
kdep3iM8Amnji4qcT+OhgD/rE1wR0uMFWpLV7V65WgpMuwyyIdFDdT++ysBX5u8DJpZIQKyBDR6S
G3wTmSDJZm0knoCErGXQMNh24cyAd30jlRyy/zIXwDQ+C/2jtM3jVzYf2u8PPwGOpP3LqwurlvIY
ZXBw1HMJfF2y6GyoUs0jfpPCd1+vfLq4RRUnVxcAKszFpZe5eik4N2noWdeO5Lfhs084ISb9T+oZ
bTM1llkDKzMmGPFHZHSB8Jqm7bFGp4XTKpIkmVGRL1tDrf2KZXxKeTaLQq5mzHJ4jIF0QRLJUKCT
91vZcbTImg20MpWt/hT0tBnD7U/OhsXq4mKhNGyHLEbt+2czIHQ5ZTCJXwfaYOAnWj1ZQbzgLsq9
S6RQL0v0T+pIepJXdvkOyB0L5e93/0Cf+SGOweNi1A4bdAY9jwa9pztStKNuEwzM/S3l+z0s9wTk
zzUgloHy6SBqc3AgnaAF/QSsf2sQO9kAfE9ORoGU/6T4Dh6bJO0o0NNiFZPHfXQ244PW9m3t63ta
p2BKAx0UVeUyXQ86/Nb+lw3sBFD9eCxPb9ZetO1930Q0BEPotUPQr99KEbUy3nRUzV2yi5a9AT15
lX5zQlQG7UtY8j+IiOUfGYH+coqXhYUmtPpsuWNTVAVY6u2DNLeggKmb/4GGq6RqSl+AwXR550s4
5AUyrgORnsqr6souoESyXay0gb136xl7UjHdyazGQxXslj7O0KZ1CG1CEvRkt1PxU1AR0arrSKH3
J0zRtZQpWtPrq24jiCms3QloK5te95SUdV943jDeWacWopF8PCYSGAZMCpeLNJeW9YA43m7fs5oF
Aq9l/CzzYlX5I0CYHG/NTRQNQCb6+zWgVHwxPjGpkokdBo9OkcNgV/fQfAskXs3vkjwZkHsQ9zZj
hhoF8NKWKC4wzoHWOfXQNMHLrQ4hSl1gVmIBAtLq3GE14IwkNHxGSWd0ZYZi9qThepxv1qSAa5KR
9CkhcNbYmeAoN56KL/jvci4xqk/g0ivvks3jzEW91vpaGMLhIWzSV9P19yUBBOERYEmIfKQ6PG4i
KgD70MN+l+7e0wiDf0oJQYXdk2odfqiSwitXPe/JlqDyqVzjnqnrdG1XzQEb+L4FWCy8g5khovan
tLhJgEiFF0ZEk3zx1SXfPfc6bKJPdzqe5ALmdXG31MGdqEXkYwemrCjYZZX4ECFD3g04AfzMZFc1
+GTKQ5Mawqn1BlM9/K92VHzeDZ+GG8sgPWGXjO021GN8NpcbG3wnldfn89RhBDK7ZKGHp56gz4Z4
qBk0GwnLZLwG1WQDepdamLr7tuEMtk0InR5++PQ2hKWwyC1r/ltxrNtGeuyW2rREgpIS3N8X05r1
6TSvCsUmLshJAnPvt/zdfo7TQYyxOMusl7OaScbtt8CbIGm3C8Zrl0hU53sFNDHM9ZQjnes+52DD
0mJlKp9vOWpVcttMOuM48kzerQuhnF2evqMuln71wbK9nW9oj56Sj7tyPw0zjsFl4WWLstJ78R0j
hC/mbMzaKMyZKbRytXfdmiWg/Zjnsty/qZM/gI9kjFvUmh1RPmQKAlVtjgYi+4z1OGF6u2XV6gah
JTsh7WDhmyS6T5PkJ7XuNd2TMOE0dYY8W+sNsL2SUvjK8VqbgLSwR0iU/MlGjedbvl42mQY8pLRB
QY2GkcCAXdZrMc0ouFxf2k+cYXeJjsy6urqdsrWZL755PVh2ywf9/JZhcsoEzo9FLnJhyxdLy+QP
rR20h5gH81wHv/cm+OBPSAJKtd5mPEPz9CFNcI4kDUcHBFAD4aWNCEQIRQI9uYQQPZ3z6OkgjdGL
tTzL3azcPexP/q7Iz5+STg9vpPaU09ZTCqXVaTqVU3v7DTK4kLB+C5BjGpoRhxCVIe/HsSK2am4O
ysSgSH+gTYJwfQolmK1N5Kttf5PCYqEcQtsk0nm/xBRHvyZsazb6hU/bU1JXIo6TQZf8KYsAsdrj
grx5PeBzhdbXeE1bRhyQfSPcghV8BQCoAx98d0tsbRsBEPWFUGb9Z7xWBJij7527ALRcuJlA5E6p
709o4AtpGMsSp3iC4Xv/nat4pV7PiijGHhjSh9xk0EssifKuFBKweWatRaZ+BeaXFy6xfJ88krtB
PcQGorfqUsvLGi89aFBE7w2/wn+s7HlBBbqtf9FFGlfbHI7CGLPBGKqIZDvzjsnTUKlRF1RVh0Qu
Qc8IHs6w0nWVxF37uf9vUCw0u5AR+6hOnMxygUq18qSWLWbucd0HVp/x0cd/qiR4B67RJlv2xCaM
A1ueahcN3e9dgqeOzgWnwOYfQSvGdWA9fyfOH07BQ552DSDfFgDz0HNU1tnfCnewJesEnRngpJAR
m4KKAhOl/r3JJvaHEjSp29gQqZYCZ5OLdT5OE3aqR1qzKY0LJVNWMZyfNlUErTOxqUtRdZklFDBe
GdX5S7kIJErgaCwxGneHPTxdraiFNW87m0OSXthGsqEfUuue0n7m9q9UafffN6rRIbGcLm6o4rXy
JUWiDeTchFnFdW9g3otmQfRMKZUP4E/tNmuBxYkwh9YCf0w8rkNX7A9t0Tmj88XpAnMD4qBlrcQY
gY6xfF4r621JAgggrCCqbUhcX6UFi5BXO7jO5Ab4xCRfeadJGf7P12xn3JkcOW4EgLUopRmTtCs0
6xWICmWWhb560wzRaKKkWOo7Pr7KGLU12t5HqKp9x6maZyVCBTPxwkNSaQOc3llWqAmVlTy+rEx9
rS254dxAFiN7R/R0PR6k0LuEu8eIhcxXH/tzbPr2ySVGE7170zk9VprArUlyzogSnMHEXo30TXFK
k2QO8xX8bSbiMZOBjdwokfA216XBgzOO+/8wtmYE7f3BUl9hZPtPcEeqXYgyef63EmX9QKcKZqM2
wmN35gAc5eK+ppNHFePxxlRwwL3QBog+Vp4jgxMXQfNb53n1OcPhUG45MJRbqFR9alrFlBLlkUTs
0nvVoxTaSjiTbxEjUlX2fbBH44I4PZg8dEmwSn66G/VrX26uTAzRf0ecMNNnx6iE3M8+u7AyIril
kvlgibKShi0KpOpMQ9khRWBxtBfjjUDcqfyhvULnJQzUjkV+5sBsseCYO+TQSp91qSEK5C7MOTdu
tabkrxYFmN1k65x4iva5dtSdE5G4PeIs9liL7Ab15FZKtZLaF+bte9zsins0NH1lNUtg1jRsKD5h
9NvA2TKml9uApLJ2nyt35y7q4IysstfItdEVkNLE2+etox7klQL6RCMMNJsnBYADrFzgJBGMGYfv
jPB0CqZQz9b7bqC5kUaKZhQWFqXEKlYKr9udt4UKK59QeDurXuFpAnwr5iZH8LbRG75S0VhIfsYW
Jf86fljoPO5JrhfOOgY6zgD1p+Y9zMqVcULcU72e/UDJnf/KzXfO4gCM0bpJ/8L4dF+bFQzHb4Fg
lyLCPn5jfKQolDcx9cZbcqhYB2CPfHMucmuJwO2mBZetw7ig6ryDUJumWKx8MCOYyUO/kM1ldLTX
0/nF6J8ex1IsJv+AoplAzDQOa/LlIVcSlKv74I58X0UpGq2dqZudQ9/oEZ4OtPP6NA/CY4RGufI0
lhp4V1abEbK22DJ4yahWAgddq3CnAzVVcP/pWATSdv0JKhW2Q9Ath/JjtMUMGIiPF36FyHmg3aqv
0YJLA0AS44NT6874D64gEBsX+KBIMe2D9iQ9KsOKQ4Q29s3K0euRYYmLOG7y7myioCSV65XvP3Ml
FA+m6zRa3LfoV/uIwlMc1/L0caupZEVLjtfcIofErN1nr50FXP0xF4hJsdUV2Mfo1YvSB+09dZM9
8ZMT4zrNg9eLXDLqo5XMDAI5FVb13QtjL+dOYVNThUb8a8rH0Kj/6FTL3oeg5A2fALHqA52MjzgU
4lbrinc/ofx2kW2WGZTGbJF7Zgki944O7k/HsENxi75i8KeJcKskQpSc3+zQWTsUCN/3+F3bQ+OL
CducDmQDTovHeNIkCVqXedTMDxgFAuaaM+pvKbdQzmlFZR8jMkEe8zKcVaCawQHzs7WWAl1U6GJ9
Us2lA9dc5W5P8OhWJTH1SvZmoG8uDaMolP9WIjz6ld2n+rCZ2Sg1eEMhKgcUgdryFtAPe250kwQh
1tD+egwpb3xxTS82CUBPw83Q3MUlk0joT3+/j3CTozBK2wePvBUW5cJFJ1hHmwur6lildrAJ3ISq
8xLFR/f5F8uevQkOA/WTzE4VSVbvRVCvrHMkZs2tbhbdx568XxwC4Cd/DrqZZ18FVEMeqWBtKME1
dNn9jQgGkTVNtdlVNARdcpL4kulxFeYI7ozuSVJoFlXkbY8q91XaxfhTXXV6aNJqIbAeUBGKUIOV
9uoJiKgQj7pA6/aqavFbJTjkKJ+Wd3p4c9uwtUckkbknFLz8sC0L5tfjeFmS4SMK0vDalAjgJdto
4Xj9FIRrJenuD73xkK4p6qGv/O4Q38KfHrrr5XBDl/Lg62tWC4s5KDJLTC7c+eXKMEDB4DGi5kYm
wd4XIPCjQ85AikSRzxwuWzaBBTcRRPT/i7RRYOakD3a1ziudvq4fqxYpYV/CGbrwx8xrs84rFtGg
xZyZDKINJPlGRWRePhp3rZ2WBAnnevtkdbov4wb5+LZcG0GDZrYwNU6/ynUgDRKf0NfP1PvnEKf3
J/++BF7yo5f/ktijws7+4bi3XxyS2vSsSEYBg4mo8n7jP+Cxh91HBrMolmwLbToL7ESl20Iop7WE
05+ayN53tpGhRr5TN2S7BDxS8o3Hhu/nN2uehrbKlaNbPE1Y9zeTe7VuvWvhIomeWyhWvn174wnG
GF+IYPDvqt/zZU3mxaTilAR20CdAyMeyOq9idqBXTiIcMjMg7+pIyDJaBdrvAeqfkIqzYXHVWmMz
L51nSRH8Y3KkROv6ksT4mK9QJJ1vBmx3HQk0ddmhekSgUutQ83B09dXo6iQQbZwLWgXMYTg2xsRy
CuVYHdlmSuIK/Rh6HbNSa3KpuLHEsLmRm4SFwr4RnO1j8cFJEGNPxqENksi7lO6TdpHMCZ+s63Ly
oKTurxjGcLEtfIreu6eNDLBEhIntl4+hD2q7PeYZHgQQOclnaDAb7LAmpa/zePTwSrKXnnS/KGpD
5QxslfnV28qCtrayjlma4XD/BqCu4NlnXPWmJmYurfud+4LNHE09NOXFh+gKL+WLbiiluFy84Acp
kWMsHRci7IKTF3mp33lcmjNV3eJLSk22zeo1ZLp0JXt1z6wdceZKswN1s2IK5OJ1oNP2SGthJN7w
sCzGKhQJzv8j0XcUkdZEA5/Qw66BNCIpcwqFfvtnUtYUA/cf1xbpDBlqILjsIUTgNR8anL9J657F
d8yKQHTyDWxUNpcYm4Kt0iubx8DYcASmXAZfrtmX1Sul6OqCqnkvfWx46KhEJqbzj0jz8Eh2GaXV
j/uGzeLDOyvBqk0n4uUX+SVqscm5vrdYmJpG2wV3B+qfkUipPjvQXO19Z+qU/80lAlOWaDemhQh+
37HViHlzH9nkEoYxmE4AySyxvuQ9myZcmgzbTpWMJLtKCDppY0rPiUyVjmVCAh1N+KnCh6Ih6eTl
yjwpk5BrjlPhkwPbnMZLgmqoaulB+dJedyjSTinw/6FCXNU/Yy0MlusEwjvri3vQsBEPVdbpMqEk
YXXeN+h1WtJ+92aaWz+GTSpZe2tAo+yn/8Nsdw5XWlzyaEt4kjXHUX2+jaAgP2OM44mXH8OLC6Vo
X3P79uHEm00TlrZTrQamj8Y23dtrt+EuQKDH/HBqBtfecF2CwVa2KN7Q/z4cKIzX7s44i6LRkkph
ZEAuatzVZSqpCQUPbhQX95BSnABiRx9UuVdP1k3jeaukTboFSIS16AFMk0ZFpbpTiJUV2FJJqk02
wK9nxu1Hpjt9hUHCmp9CLw8Wh2d4O2UvP1cfl57LgQMTy1Lc8h2BjMS1DOc18XCx3dBRythRUF1l
2WBFbTthPqZJK/XGxJk6bc/SG4QixxTkYpi3jdVeTwDVEZqfQUjroBimh3aiX92u014jPmpRMGYS
G+eJA/Ar4LQVb+VbK1v7qgO3gtMkP70Jtafkub98fdalbXPg1rT1bScwgh46UU//5s3qJU7pVYLc
2cUeJc47NKbngulSvS51jhXilz1Q4xxI4TTMERvmXYhDYSvBqum0Z/0lo5Ka5sJ2QixVWqHOzWsw
olqq+5k7oydbecKzHVVD2aiqsXQnfK7y+cE94s3RWR9ckDnDH3GKfP7OrBv1v4FN+WneBjfo07Ij
eUV782TBSysbFZ4s1okE6DHc0SSE0d9kpxLUGjGuPQhm7XHA56d/ftJKkfaTOVPolRuwhnycnTsL
EQcixd6KP48q8zp5qO31yOu05UOrMAWdc7+HBoM11NTIPmLmVHhMHor+QBFilQ2M/WNaNdBTPfUi
QmAydf9URSHhlQde/tqkUlU/aAT4Wi8zFRo6eA3Mzp2Gd047up6UASs+wx/pi3nKl7Z0RcIqJfIA
OW4wOANOTDI9uV7sBdgQkAY7yf1TsLqBzu9TP4e4DASHLHLoTVYDytMG2DwLbP2Vm4i6LkQx5BNv
FN86F4wTpTyLasvw+pVN5etGx2Pz2WTcSRcl4Q3WGHlbsAhnveZM1/x0GiD8cLpu6VfxCwk5S0GG
EuYTb1IpFMRUBhRdOVyS2pQBIbtOejE2F/hSCektzkHvTshz78VkY4YS1zorwX2MmQFxl2lxdaBm
rMkZFzq5bVHjCpLJ1moNpjTxV//oZ06rtyREdcNh8/ftGMY+gnnQ0WR03bgdgp6pG/sRVW3dgLTL
g488H/mETcvX9C0GkAZCGiam74eFk+drOgUmB2SbJV9KwY1cAiZrpJW6wQSHh/MsbbcMZbWoXgvQ
6TgfgynE/cN4oQwJXIfYispnOz9AXiFWeQAsCZagnk1Kr6DZj+vEWAnbZUNiZvqaPkE9Mo19DU4Q
3pjfXHaxoHaK/H9nlDts1NygNYLmIzeZDT4sM8frEGPrX56Nb4cP/Pq6767QJwXktmuPpVPyTW9m
e15Nq+Qv1UOs8N3MHkmlzk5tEojfyPHqZ6EEPNlJjdvNURa21AcSII46ksWS/EtwGax/NGgLmVBE
/LPlJmSaTi7B9QCXxHs33bBM6cXk1gBB8yDNmPS8SBap3h4TLEO1D6GrLJSGavOImrsqWOuhhfqH
VM5AA083qCqlK7pndlTDEIUMbyreEVosnlRChdk1LtvacxCWpfFYqij6mk/45EB6yv7fIqg6RNsQ
amOiuJlYkkx9u9hWzVTv7cIDOtwb+F557G5jB7ywBUP7M37Wp7Rj2z786TqekJcc+KHIR9sGsJ4G
xSa+yOo5Rv8WzRWYqj7XcIR1r5D38JIL7OfzxcHCoa32lCUlYCdlcsX3pxvL/tvxOuMRGXpcNxtB
b5evYx063coj/l2xXcvb/j1vpjQo9CbG1iD5ZbMfxys1hRYhppPj0FuKoroUruXgzih1yW/3UcEP
87LyBogFbE/QMuFpkltujCxd7KQoRgzGV5uTq0eNsyu5l2gsOu07TTPWHSmb8eIK/4O8BsblFlqX
ps32I5HDnzbF82qqEAqqQYo4n2cOUl/IltBGpxa9huANqTa6opSOqmOE3nS4K2BEMK5aEYUQ41tm
bPco6vJzK7PEcGp5bom7Ni3y/kvOaKNinHFe99hGSSXxliV635BE6wDJAYCdI5xhXounVc//Upz7
OSQMTZBF/TJLkLPKzGfHkxzeLovem8z7qwlS7rDu1Qr8LoXoifArlIaNRg/SdZO1iyxazm1CT54N
F9CRL6rCGrD1BWOaFZpKXO6h0hsm7wYsWvISFwPPjUb6RoIGUmZvCXtZ0swb/O7zOC26233MaYoM
bieXkWJNU0S73rmDiSfcwC73wdJWRb3aanmqcdE0ewBZx/UFQJfw6sY4YWs1RIPNhvEtStrmeGXI
MdJRMCtw+Mbsxu7NmwTd09XgovFluos6PBD5AyGegYtpcOBbWqrnUXIV5guwK9ccMh6lwHiqn8T+
FMfsMwy/JC4cfdsb7R8pGLCw/aGgOV6zhsdedp9sMrvbrWg2hb4psLxPtyp/MbBkIw0LwrqUUsEv
EVN34ru3p8caHkxthR4GjenXSK4zVXgBtTCvsyM7dFNwfGctXCyiAI2g9TZamaQLYqO+5SmL5sSo
Qe9fHQh0XsHgXGW8AYEp0YbfpQIuKYwo4oRqdxfPK/ZS0imqjENSZb0CFlPlwe5pxXyz27gwLRG1
qw1LxgHu73yg1XLkL/BX8rc41hYFW5gPXg8OCXkmpMp13GuMRgcTCaPoRdVET8cde8Uc/tlULRJX
esn9XJVvGUqBQGlhGEE+5Ayt9KTX989oLATE2PZiFIhakzawZqda96vUkNTdTNWUqxX62RnxvQ+s
xDG2QqdKb2Dc3Gou1YqArv1/GwaT03J9LreQj4J3i/Eq6FXiRgCcViNsYhY7nRB4HzoD906mPLBW
Qyz9fsL1IA0Yspdyq5A8+hdoZ2kOrRNSh45RfIsd9rS0O7Fj9zeFdfwTEHjQIXQmddr+vXTj5txb
IwzdgRZdwHPkSgPubZcRUEWFVdRKDXY4nahdBBJUYWqXLeQCwPIcVPOaDkrk6tL0LK+everbjX1C
OuwaIL4nswzzGLHectlClTch+roJbvs10vsEz2Exg/aVJe27CelnSgvu4CPCX6piRLcl8OSDNJp1
De21pAQCIXRRW33jhqqYJdSKguh3TppS8pFnL+RrzWIXVIGhRacoRennbZPIXXhR99R5Qzjb0uYR
s1GibDWs1uxANqZLo9407ahd6cRBZeZJXFsLjuMXtwOJ1fN21/rh03s53iknPx3TZRZ0KpDKeVaH
spgFvepaLGThDlBO8O9FUbt0PiNKolloOkWQfnfsXSuEdqrxQbJhqeX+aqAHWnTRxmkRiQtLSCQB
ohu3dRZO9MUnHQqmf/1Jo/rRNP+tbNftxGESLiIUTUDjb42lbxmsq3lDDVm/dfHIKE6hKBw3hkoi
W3MmQ+Wvpq2N3zDqMoqFQP++OykKlauNs4Nu0yRoYHqV3Pm4Sot7/jACXNEwpvE57UGK0mIG9lLs
spd5XyqmJuvZKxl8bKKDxdRm7l9K+vz/21yYvgljNJ5ap/r2erKKJJ892TNdIhw0lG5uL3smZ28Y
/UrCSUIbtDu3eTlUxlMQd4tLujkZ7qZFd+GWXe6zrjrwGSjuFVx1tfRx4JNEqXN00jU4nM8hBIdD
j0wBMmgtrWl17jFQUbY/uWL/rixjquO5wjMDcw0JwKasREZz7wfPW3ig4ZI88UTnkJ4st718owuX
iUMQ+XrC8/kmALY+0/Ua9N2mrn0bkBrVeQ46f+qXHsi4Zjm0PhJFppJFQ8smYr5vPMOvSS0tJq0x
kmtkRhJ5k0sLmIzXhhP4juVq3CtmMSQVs01nX28ibjb6rzkb8zTYIHBCrpOwvjeRnJaGPsn74nqA
fkkz43d6vkef84MrTJKPbtVMgiFGcLPBAvzae+1UTzuYsSg6PU9ed5+lOSJpgsSxX19Ar6Xkdq5m
WeumO10N4LkZ3BqEF6WITPItqwrlpBRquMCCiS0IA/+BhekFn475qmJhVzucSmTgxzgnCCFVBKIS
KqAp3w9SMJaVgbeasr/37+5xOdbRAbOOSaaTVK4QO6hxmNBAOmuyDBGfjTspyq5VvobWq/ysVNpS
H5IZ2O3pOt38MKY1cxYsPZdX/iutQFtA8JTerLyfcIWCozdu4e/pAnHzrqlcuXQTfpwMketLje5A
nHFtlRnzEHSCVdpwh2EfVLpLYnupq6TJsVqW3Ga43v1H5YwprlXc/Ghbr/py7BK3bxieosbIRtjN
7KOdfS0ikWB3ayxVBrDBkyYKUMdy3Qcet3TlhBvS+UoATIKhRL+03VBxMuQktr+ceVS2kizU1Fm5
Bw8+YG08LVAusDSRCgBRwimbVX9+e6FdTzoNnbJXKmCEChxtVRhAmcdKIUkM1QIDifMXAAzUxxL/
F8JyRSA/to3d7NleEDWmmMrgbm1E71f55zAbQrGlki6Bnhui+ay+6DFgsP+x8v0QEvtHez759EsK
DphoiRLOUu3jQbDa+Kh3oZP2iCpaBw7V3bImOG4awfhdLX9Mrh1z76tz8J2A8owka7qAMojqZJzZ
cN7oMScVWLWJn7gUPaemnGwDozO29KFHKhE2n7UUoO4DK1nn27mss1wQi843YOhSm/vG/EM34QnG
gL4ajRrkMzY2Zx/t2EpZRpWAnLtmvWg+YEXGjfv7VuZo0LH79vQX57uk9I0nF6dniqz3JgcpJZbc
9tKMU4fd7Oe644az4GMCNUu9AmPHWGocgBY7oHWoEL4qkR3bqiNRHoETP8ekVkEffLFehFcQpxCB
hAnHGIELpIJ+4lYxDNLkqLTKjqI0OV3diHo+beG+iBfJksigBovSNUphv/Z/dkH3iO36L6bfvul7
8YTvSpAlzA5KpZV11iOHTbgXX0j32dTL7DRHN2kwbCDcqtBgOGVW7Jhsku3t2FiJEyCLRrTVQWoD
Ud06ZIPggHth8eLjzR2yemmxXHwUjshB+ltLSJ100VFmVOh91TNLn40Hrqe+Mb3GhMGRcsEEKLm0
UqgrGTzUO2/717aTB0bHJ5rbpGpoIAlOlVTzr+vTNz40sojRoWgf78T3RIO0Req6SMpRnKbzty63
HrtXkhR9WjEfGMY0Srva6R9+ksBSZDrpr+7GC1LlNwe9F/8OzcVPvf+gRXDm+H8S4iGO4pKXBYS8
rMsRINoMjoOlX16brNUaJuHgvNDC2Ztx8Dct9wXUWIYI4EKMiLd4Gzw0L5m2D20S4ihAyIvyTWjV
d9m+z0BZ4KiZQ2njrSHDlsVHEYod/tf9cyCDiLww4xpL25uQmXNtt66+8QiGjFvsJGY9nUuIGwOW
ig/2EojhF+Qk38NccxlygYUWo7pJ8XtwxbtOgB3hS93GiDR0IlBbR/mubHuUkR6K78e6dCj9M7GN
45y/yrBb0IX+UCrJjPh38jmxapubmCDheUgsxRTHlZa+kDc3HU8G9iGzg8OI/z/tSxBJG5/33Ttg
4w1KYtPsGgDH2Ykxht38nFe0Bq/1ptpievlQXMDK4iv6Bhm0Ibl/RcDlea+6eLjgmqeEG5Up79k4
CoZaArqw81TuBSFTS/leAaxo0wWFLv2UUBRJGWjMU7kBlXIMNefMgP0WP9hb9jHkLAwX5Vqz28F1
1xtN+ljHKEzjmoepxiSD2eKD0WqP7xhupSIeLup0I8fGhOMDsluYkLUzTRG6xl2W+ZOOCy6N9m0p
98o9O9K52S/bt6vWxzyxLlSGvd6ZazzV8f/ZIsSzXwsa8O0pADx7wu9P7IyzG7Yo4ivRK66DZh4N
iA8pcvm4SrIKA2cJc4Zeny3bt6li4Mcw5WffV7+uMRW3F1H7ctvRPniU23w00B1eo2qBhDaq2Hl6
I+CGeYFMhjTrotcMo7XoBaX9nGCnDfP6vNPReejtWstvzGR6y+iBU4c0DnjDZKnvzR6OZtSLcdgB
IBTvF4JCB40nE3YIGiKpeCsl/WeRjII5QJDlRtJLj4TuMtN1xfjZsAQ4YjDUHxRn67zi88MibrwW
VVMTmRPyBa+jt03lad19OjsL5LCpWzAu81fB0VfKu0m35UTFlwoy/5SNS48iHsAQcAUz0rTp4R2t
uTrOT6ea9hoaeAg/owBFlCrd3HItHz9rd+dcH6sMkjF3C1DZJc6TmBl24MYuvD644htLGGFAdR9B
c970nIM71w31v83IVk/6A4snor39wSpd8Qwoljgnw6MrVdmXkK1vR1k8/xoKsJFoG8MCjhyOoA4c
vXCMQC98a/HSQlZogc1Pz1W55D+ub9S8f0ELO6vxAwNIVw9HW3sUmTcKXwh/EdKUGs/gHFa0swN7
uxlEBKxmqm41ZfQc5ZMOCu3KHAeur/TeN6p4Auta1fxYd4ATkZawQIknfqfEK+8i7b3jTDS5AVl4
Nvn7WvzasPpQ7p/ukh3nhy7FHgr39lZeVbw2SMmVUTO/NZH2jL5XunrqIwAEbLgQ3KWMleGh/7kd
3/I4jLyVWUU5xEiFkoau2GCGDLE6IsojAL3bUvn89XzCFIgkLDKSa4tGNfXZPtx5ahCYfhDwj9E+
bdFjLK02cAb2t+DNYo7S/Ere31II/5JZsqLil/7WZHmB58ID50I8tfIlmJ/Xo8vAs4Y54D/MRXhG
nfoKFVRX92vpJ4N2UcOEzisOyxbU8d+ldq/K6LFGaoqjXpLtC2MkYNo8bGBQA4hye93AQKuaPgk0
mM31xsp+aRoO3RhSQX0qO7yFJe0WLWBcTtViac5dg/NaRRR4tBaoMqYlds7VQTnRJgBUMh3AiAOY
K8o1nFRSuuGLb0n2IYhpGjkqDeW+yj0i/qEqLyNZ6pk+GIcMd396Au7suzhP8ZH+JDbcvu2+PgQM
a75CtpOLZk/RGxJrpe6IO0v7jLinO8/zVs1/clhUjAIYH0WrZOjZRWWs9QuEceihMrCy+6rkWF39
uIuWvJv72N6BY83i+z3J667OdW9vfZJHZ+nzXPwRu/BTr09xpM4e6KJLlSYQjZAc2+TNs2im+Dyq
qcHOsa9LkfSAqj79rvX8Ns3FgpWdFWtRZ+WqKKSJtR4XrE/rvCc7uedMi058Nu7+WXRlGw0l8W54
w5dxLeUmckTcJ/9S/8thBpjexyJI7jM7XEcdjGcuTBUiw1elwiKuIMjyDb/m8rUxga5cZ+lNitQx
Qw2dwU3F+42ILwDnFJ0cxPiVO+08JgHlmtf842Xnenm6ObQsTMe6wvBXOPXWjB4NSQypF0GxBAXJ
ms8u928htHIViGA9HzNY4KFSVa1NOqVaWaj7fLUq++aL6RQGmBuuizUjMjapZabI6A4mVAgEXscw
8p2SWkWwVhmggYdM06gpmH6sFnF5eQPvJw8PD9jT1NJUAcDs6pbUbK1uMsiU0vuyrn9ChzVyJjB5
WJ9TqtGRzcYqv7Stds8b/YK34BuynOzYbK9Cjxqd4vB6TlI/zZcHJeUfPqml/HfR5JPOyieCIpoG
RyLxsM80Fb8qBgJW0CizC32fnhwcGfGqtH1g85ISu2E8h6gDg0Qu5nE1zI9fGBhk7S+w8cpgrizm
Urb8H3o0C6jkpiIBKK4pL1fuPM7JYRvcf7bGBvDV588aXHLwT/GoU8MrYJFsKNTt0Z+obuESa0/L
vcpGBBbKjZxmfJUAbXGUD5pWGlQ03zGqng9layZGRw6N3+UE3N6DWMTsS9RCThHG4Rl3cZYLcA+2
r9Jpia2icqJ2alNQVc0GBHKloYYeZ8sKDynhaNX5nI7K3/guqKrHqozEwXGJOfFLNxgmgrFnGcz9
oMfqzIEurd/9GY1JNRYnKZ+xxE9arqvFkA82nbgBBGfJ8Lb7uDCL6wkUe6Fy+akUq899flar2JLi
KqLuFRmWWHLk+Fqv5Fg4GhjqWxJOOFmOk7+oXB6kOUZB63EuvsEcSc9PwxU1lkkcx6qioCLT8LnT
0Unra/tDDU+ptaGOOzT3Snt9ruf8EnCDhTczcV47XV91f+CzTlMabedHyHcv9QGrcuJhjF0YMrEf
n7qkTpBTKYR1S+xPA87dCIQXt2psdqz9UooNi7hIwmfrQaNOZw1wxp1haOWIidoQ99o1WK+a3ph/
sXxYAeY3II76461sKFU9L6NiYJ5GZhvfWiABapzviRi+G3dVyAqVQYfT8+QtB+vXx8M27x7/qW1I
1AxkONzkUBfkmKJx+UV0di2CiGPz8z6QXDbaUEkChB4uUSL0GZwU2019DjumUi5kCI4YrQl0ysQg
zoFMMUKaef41iwbMjTUNHiD2KEV14OMw9omLjWh7M1AM1TP1YMCDtlqVNkpoitX4kGhPDzdYnFTB
b0VbQULS+BE1uZzVjkf+cI9+BwNGulSWwE8OeVuR7ihEvxk84Sxor9Qd+S8RMea/CxW7f1AHdjOW
sNvIOj22iku/TdP3W6EVOoaxgATfA+1WXy21RHE/ig7ELeyEu5IAmvToBxvfqMXUSte3IiZw6Nqp
OoworlN1MRfUr2yHkLrHGQ3qDuhXEWbMcrU/aaAtafdi5kLt0zmzasMnh+o3Wn7NdBgxMNNFxQ0g
5aARB3brp6acual8p12XqEF9Rz0g4t9Vg7+sYHWqnHdaHkVHz9B8igXXVj7BDh7v7TwN05hwQ0Ne
sYLZ0XTDJVsLCYGXw3kN2ABmWWKLH3hU+nAVpjHDwud5FtwwUdjh2xrmpnnLzWlrKwa5wUyIbmhV
CYrmWeggIg5gskGDmqdMYCnkJmpHlvFARDFThAqlkAFtkwfMyzbzktv9bqUBkfWftgkvzvwXalF4
+PEbiaIovHxQT8IpQYvnH5ytNxB+pkcmRXUk+WDlAaBcZmlpelZCLTgy/a66RKFPHDuazTFEos5n
51ligruigPWIv4ZnmGcW3k2fQODt+7R0S0hZEVOoLXacxwYlFZBGXtR5Y/d2ru5ry8tVdfl+rkAI
T3a69zdt5hZuRYZYSFDhIZ5vbxmwG/kimb5yZLyUyX4RndYpi8finXsLxGM2T/ZPs/aN3axg0p0Q
8Ct9yeo2+akLGEta6uGqxjWkJbzPm5+Ikui8tliGEZC7VnAKLfGgdPfput94dFNhmVuHhhfwFlj6
VJzuZCY9aP3ZVD0Yfg1SCOtcnFhsXAHfkE/kOK8kHnScewfzS5Hv7VjQ9a6gswhviQzR/H9ob840
xik3oFXEQGgyHKGf44SnZxBJi0nUiU75CLT5G/wFuOIrNq5tlqIn4kR38oJ+Hua824MhDjnd0ENT
bIX/ie6FmShbe0BsW4MjsOWmc5mvab4elNP+6MMkGuSqtwPNhmDj9kojWa6inK+CsFHtHYKJiaLw
W6wYjeh5H1bLiyOKvZOrMUZs+R33HYMPu/sczImiA1VgunKMIB05D/WbQcnky332niPYuNL6MFKu
HbAQ+WN708Lef6uPtte3LQO7o2mmo2teWuDpS8J1No/j8NME5lWW5cz8Ix8GZc8cNSp9/glmA6Wu
kYYprvnaPzc54NJbGHtJGFBa0ARNfto6wHxsWjWU0Xe5mxmH9hKmHPcw5a522Z31Cx+KIXj14cYo
oO/wWfqeY2ayEY6cz4WVGLLcsYnBLmjmcJmpL5XzLaVA92mshPVaY9uef6G8EQaziKFDDDuY4qmj
px1g1cnCdd609TeMcQmOujTwWjDfkDIp/JW11IBU6TdAmPXOFisnXeRjohMHPKkTl9COO6PUVNBq
YL7QBm6LU+jLWwg8YrN+BEVWjdmdhRg3/8uWVqpB5L/ShUKFk2lYF5m3F07HoX3YPnV8Piva7W6H
s121NR0PwCCNPv9I3cPyl92xwnXC1e7VybGAIIA/PXs8LHNGBwAhaj4qVKEVSCnDg9S8eHDB7MBS
Vse7dFURauzlFPcfJaFYSBFOv012XX9/v48ykfKWhlRlaVC9Y5kGk5vzQL/EbcvIjQxbaxNbex3z
BEbhm7nBFsdN3BneCz/0vunNWDCbOLsYRPttCgGq+6938Zq7alhxCdLH38IGzokAc/xxzswqw2ll
QAO2cVA9am1hDejDjL0FMcnm6zXvg1iLPn4tHA2vl8llOjY2XIdpdCBcfgZwJwbvaHtB8nD08OLW
n2f3IsCAcoMDk5aq8IjqN60WwPdAfb90CdUz44eenWQ45LAFp6FYj3bO5rhy0lsXWxwvDyZFbkgA
LujOz3lt2+CNUWuogjLAsaZIf4N+tFthqOwbV6XAe6uj9YdqKjyEF80wHbZQbR/YSwenHpM5/8XQ
KllvhOXkG+zsRHV6M4UGlRDRUsBuD6tvQbVNvTCxKekPOUR2tVHtcTd0m1XeDPrCqjpeQyotJqr0
zRoCrBhSXSA17NzE5JkNuwmxevPBwRhcTf3ZffxMxU0JQ2w8XF4Ixy+Toyjv9OZTQT+PGY61XYM9
nn0C654TkS2/vKa1QwfHm28SCQLXi0eAIqItJ4bXtC+J3PyW4l72xh12/85mgNT9JXeDB27ZDJYd
3+AbD3pk3wacfn6EtcWERx4ORoZ9OV8vLaj/ecrL6gdlzov584zx7ZaXj/QHTEPdex7tuSwOZaHe
4ipVFyArAtqzGCk0ZDNNR4RzfpRNy8Ou4s/k4WR0r0BFl4Yqz/0ne/PXAScQIWN0hrI3x+m/NhU6
SFmk5QbXIbbPVb3EQbuoOGgdkqNb7xTldQ+arGvYiJ1I7wpe/g1p87pqwCitWONdHEEtVJ/yHBpA
+sKS0Fvm4I9mXIWMDUA29zzy7jn/Cr4FSm1+H2m1epIMAP1onFc7aoAaSK1Viwk0577az+iA8P+T
Ze+zZBPVhCSdZ15VW/DPCfR0AaEY7dV/55tEzjuR3RLe2Pgic5S4nZ3c+B8iBgfZ1xGawNXW0SGe
nQ/B75ryM5KZIWrfj7gLtc0PkfuRmDu+bqwJolwQLnLqzRX910q2edhBJSGzquH8Y+4FrvHKdGOX
U+xG9aumkTuh3uaxczpAQ9gOngie1jLA22GNULhpH6DgOt1yCTjmzXntWrb1W4iQic6nSyNCcG7t
23ReI1+EkMT9V8Tsubb7SHWKHqfJ0jpNS642SRQypeatMYB+7nnYH6s+hXDKbmqmmWbLUu5Bkjt/
MCYRuniVzEevJCzGYW/5NbCu9W7uPW7Z2kEIiHRrfoVhCCdWGyJkviMHVwRrivlNswIzcoZSFOfh
0EDbx4Mnlo3YyhL4Xj/veDwk6GSrXsElpv9uJ+Ezf5wssQl3RwB0wz7rdUnRlAHocyr+7EoLhkNB
mJvHV9JQI02ncvuIbOlbsWMxm/xi0+qE7ZyASwsNMjMw4EVU+7kezy1vBwhjPEqo4HtnMWi00+W1
ZZSdgJ5i1plN/iFKXeCfxCFHNrfVIYsjNeqyWwcNd5LrmpqK2TGWBBiWq8s0oLOz3CWOpt2xcAbo
Fk3VFv8QF1YcJhuOebzlvUlyABZiqp4aeLOt/NPb7m0Yt6QqdBnPYQ0B9KXpecIThICACdETJb2u
4lN9ITB2Uvt/Cs8FpqchdBzjckL+V/FUPOnIwBlWliE6E9APoHvNM79/lmK9ZfMWzmZ2DVt2bcq7
3AjvZN6E7l1BfZ/nJnQhLN5wkcmIJlGHamCSlCSxfDh6MHVmKFjFO5CsW+40TcSZYNvjBJhO9jFz
mdqQVAxMAgzijklhh6GnRFm0JRQ8crrZmFfO95R38Fv1eC2MSdWeWoXulR+L9JokALH0iyUd9xfZ
AuDs6NWRyNjRDLaoV+AErQXlli4fAV9Vox/Y84dB0EC7dOfEKDyJQ1O9pvC3aDUnuBMCsEYUTjXT
kdsu0or+PgDeehPiuXL5gzqoe3ruWEF6GBptKbsxBrVQXCPc9rTlcBgMD1XbF8IsswWFXwF/Gthp
q5K79fstwqazapO5Rqt+wZDgSdQzzJDaaP4xp/y/Uf62wE2V3wAQ8FimNd82xAhB75/ytIPuXWCS
cvQGPVDknRAspqZ00kt2nj9BOiWUUihBFvFy9PRv2wuBYvnsLeMNxJUYBYZHGksCIwr6bbE6cuVr
KnAXG059uYopnXT0lReKQd5JwRI9FAbOyZ03olH6BEYqBd7xMN7LPp3VHY30qQ78l+yifjOzGPZz
OnDUYYXZVhQWv6Y6PtqrDS8ruikuQQvLM6KPfz/3bItFUxkouf8JCKAqlInh7wF73s15jGU8vgpB
B72bMrhxHt0YzANmTAUVs/qbbfcAn4C+2ANuVbD0AUtJFI3lc6qulY2BvUMYxVYP9J91KAEKuyP0
4Q0o0Vy7cQidMGFMo0r5y6UUMlJ5FL4niGcgoL8yvu19VcdwlMdwyWMYYQX5/JsmDvDuorxWTj55
/UM7O4Rn9TqWJspbRPDRqsrxzxfMUO0/wta741deFvqCk9ndQsVO9+4phIFuKvDYLcCNCMmrns1h
7oAtMc4z2u0UGy1jkd0nGRvXYxigwhH23VSk3hwe7qyTJbJ9B6Jrd3gxFzqw5wfvbsX9UrC+pKEP
Vge+g6KgEPgEujhBMVw7Pyu0jN8LNjwBi1CRbi42THlXyBmltcQ6/Dh2rMwVBKhVz1/9Y77wh8bv
UQtdnifm8mhpKhf+WyI6FtOXmV7+7sOxoTfwBMxKNXAjMl9X0elzveE57FXVPqBosWFn33S5IJ7H
1+CzCElbaRNPOVmUqoGApekBRXV0Yo5B+djidYnm4tgtfbBO1DSv2MhPLYvStM9Ai/pZTAJD+BSU
Lrxy99rFxmZLOHt5iRicCi6emXETcdJn47vV8cn7psmgH2UWXKCxhztsJU9AGIl9RVYX53Zo9rNo
q7fYcsZifIfJ/6+zivCt/CwdwgvmUmrNa/d4ZD9Gz4DSSLJ2IYaAPlLXcUuJAbDY6UgMNjClX2S+
QAnGczlelfZwJ6RuBZr40Ad8cR2D0G8g9/hjZuw571ZMLisF9DSJolNOAuBxkoxYu2M+uYPhq4et
dseVRAz0/AR5EvEo1h4qktfiFnYGO0aqiMBtFzUX8P6r4tzR3fl7abtDcEQ1ZKWcljJEg8s7ZfW9
PM8lWVsMI6Q8Sw/9kYHc1npg6j9V1sJHIy1cIPCScpyaq2qPJN60wnK35yrpPLbjBYF7zSR1xeVz
cVQUG0VRhXmCwrz9EJ/AcnHjuKOedJstMs3+XWHobYZWJneO8fx7rlzDitCZgpfSVBeVfqZUF+F2
Dw99d7YselUF4Je/A9JxWP6Gc//w3gjMKiCbWeZM1KbrS1P2n03mhyAX2Fbt7QO9xN4IMsKtPIyk
n9BR6qWRfFDPXZSHq1mydzhfHLZmu84dM424taWJzBZR+BqTACBLkMYzhl916zyClzjYnkK1EdX/
8Smy+wdmsvzEQ78SRRKc5p5YWbEkg9BiqfNTby7qolrb9iEtc3abG+TcTp+bCqjC3hpE1sMGgsGR
0I6CC2Nma3xFZrvFV1ZEufFGsL+9qMgw0bMfiQJ5IKqu+DgfBtnGt4SF04TwE7veOa11AP0uf1PG
KBTerZLqC0tpThMoygb07mL2O34RFKf+4nnWhTDDVJPUoPw68pbOMnx4QOkn74+EJqFynE9n1cQo
4t8Xm4pOh4+F3AC7hUxcUP+NuxWnj8JKjQOlrI6X7DP2IzBKdo/AGRaCmv1sAVBJFrdzJxMWWPuZ
nptkrKZGwfzlvmRfxV0z0pKDbemvdwwtRYB/FmvQXafhNgeYTObeiXBf+Jz6Tx6k3iCeJ/0Nk1HE
IgOuF44Lndj3IfGePmg2aXx3EqokDsO/7vpe7PNzd+YtYl0KPSxHGjWPquVk52mLdoe3zPlSlA65
MiDpKGoMQZDbXaj2XVlaIgj7rucubVtP4/iZM+x9t3E1Tr3vTo705LOyCImS30JrMm24zCvaLjLT
W6MIVhOcNbSYIhgSJcLidCj9YG+a+BiyyVosDt8zYHbEwQ854cZpK0OToGEhZ2ExvUYU5Z8sDJtF
y/Yc1dKzTPll1JPXO7SPMwIS6OHY+YL0gIOP6RMxi8k5F+r6MqVdOGdiircXIItat8AzdiBpuLy+
KAp3H7L9aZcJRBjfY+WkAXN4N4r+bKUbylin1yvlXZoAJLo0NE166+AEGPId4A/O+TB8VD1oQeaZ
oHCSqMrygycymmqXgCDUFvQTce56FLfqz1TW0B9TlNddQQanurf8t8E0wnzfP2M8zer6KijiqYn8
nDn6vScvOfjV/B2DS/FDrT7VNUBsVIYHbfcZW+5wPW+C7Bah/B+e/tHeekGdP6JJwbyzaR3+WVkX
q/E/1/mLE4Ucr3SdIY7NYmqDVlW3OsB34DtgBmkTpAMusQqvv/0iLkH/cZyKrZMHvQk5/CcefgXm
4W1DOLUw7ZBE5gdS8b0AUZhORWNEiHZJTIhlLalFpv0yFxiuDWkOkmkcaX79K4zrWU5Oif2mKrPu
W8NnEcFQsuv3y8zXOmloAkjxlUZnMBrKyuSkqN49suH29Y79MC1wA1gGIpEs+fg7FXwBz4foOb0s
11K2crOWQTt/h7aNtXbQLK2t0sSqquAnxecX8bhh6QDMoI5k6bkPf2PSYKHZDtuT3BVzwbTelMss
tsVepl4YFm9r2LUlal4ZryOo0E0+gDlXMFWteM8Nifp94xZ+f6q3XiOFb8MsKowBWX+Qw4j8+fqo
Rxu1Hfe3hGipEQbFe21dO1gSBS2uHLgaRg+mG7OrygU+CfJtpcmMcr2bMxeg2YdGhqETRHFNiEW3
rQJj9H2WL7hg9ivTXuRWAR5rgv46nV56AFIA1AsNnLyg8bZIhhfk9PP2/lS/WBZAPYaqI1wp4wtC
dBmMDebRGkWAJL9fa3gcg12Y25Z6ckTd8GYjmHRDXj7kAzXCJQlnc55ROIVoVp7XJszxChbalaXm
EvR6k5QhZQ8REqT03r3wo8G5bGZT433E3TO84wdm4d6NsmATtSBnNzyWN+aLzrI2mylwxt/rGZSS
yfy71XS5FHc6r5WUw5Ikv8jbruKG0bRhxBWJghLlG519i4N9ukGsSZ64fpq4y665UZImVFR5swQH
uA6wQinA4V3V8c/ZO+HdqBHTp6drTZnYZUHckbVbj4+TfPjqtoGT8A/PJXkcKhHLBqnnq5nQwFOG
SBrdLFdkySZO6T/qeQ/rWwl0UVrbyDcI2kCUGgam8ktyXFISasSn0+oNhIj8TQa/h+xZpE1UETyq
1BDdt0xut0ucEskaBpp/svRpbZ2EE6le/Tndlu/J5qrg27B+VgO3oiizcH9zRPwsrATorZ7XRbXm
4/yf3qcPpIXrH9o75u5WAWxcQCPKssCW3F/hATgz2KLo8Hxfp9yQDo4/sk294uxjBSNQNz/+/TYy
4AnCfO503/ZtOqXbq6oESdE2RwbGkOGgm9bovnp6EyHNlVguuVMJEOIbYykhqmUtnUscuXCYCtCL
fBi1cMgLpv7NPYMeuczi690tsoR7L1CtENN5UWQFLGQyjUpaVflDC0K4DOAB4Fdm2NtjtWPHr9JF
sqR3QIeH+UmNcXS79ar7r+gEUGu3YtbpFYW3CmdzBpKKpCVBRmJ1KpGr5LXokoX3H/295tA7zzfH
9JF0HM/vi/TQgsECCYbC2sg6qm5eGur64LUY+4lAC7HL6Uir/Lh/ElzpsPCYPjtM9BcDKsmBiDIo
S36Ihwj2jbtPNsUiClX64W9LdVclOoDwblyqLVTQvKJqJ8jFRwAJLLbdfdhAqHnjkx/QHPgyzTR7
1CPtZdwcVWOR21PZDvc84oo1gT5dInuHh1QL5MZrkrligHRoeXsalgesLKeVoodIf3Ix4OL8DIrH
yDSxBOr8twwgmqXRNa3LcKPcd4cI5WAOEWiQU2P43QTgXKmldeAwasf1m4f1HhWuZhkAJ9VzWV+9
zSneUY6GqqlVRKwJg2U1Rx1p+EGfX3lZLNMhnArRPiOmgGJ+d4ZHgMTdWenSLnD6J2B5e+SUNgT1
r5I2dcuTRATfV8O7HySsGpulcNBS/kydwb5NLJq4a0jAHy2RtBuY0zmjoSsMlCXeqCVN9m2X2ZQx
flqy7aunLlJWLgQiHy7ATdAhmcGfnIbPmch7tAjdNYzIaJNUItrpbKaTJvsxPMqwtqcR6BMerd4g
ZbSFx/ZHFgKj+rswQF7ASq9ierAS0aQm3yTy+yKRRSy7mVwmqJfmZ1Bv7riYuA8xQTdcqctX3vqp
8/8K4Hd4nW9/WH/UKh2+Spi8p/s22iihUkIvFfkCHLr5vEFcJhyEUHCC/HA5cSxbM8m5YtxafmTM
r98ESTMFG2eK2MPPbagYeVK07QaAL/OAYG4l8y5i9wxu7R4mo3JxWKeBuOuKbcEDIqiw87i0IlC9
S3IImkk8KjAGcGCluCThEjSpkM1MG6780bxqgWgtAWj79uyA2cSxDXCMz3UatZirNvdfW+fWKqtU
0NuM4/hDg+ZvH2bQS1totms1BpC5xOxPHNJVVOauZ9K9jLzs3EXLyyI1pECXtTP9XsHS0K3jXHXo
yJV2il3YL5XCKm/ZQddOAKAW53GkijxVKlvMpFijSOAywScv7GWTvIE/ALFpOwFEH8AmerU4aQFx
Skt7cVdsYpuu0+sFkVLkmOg6vrqfFGEVtTVeThJRXwCmju8fUd88HGu1s1uqhdtj1+dznDWOflhz
ZlscpaR8+Anr2hISjdb60uG0q+lDtX/5TsQYd/BsbqSWDoZQURgODktBboW5QTFbfZWex6GnIt9g
b4TuGDMbnupj5OD3p0N8qwEaqgVMOJ/QCUqvOAVeKNknDA5LXQzmdpTC0NMicZn7T1h/TwDJTzIM
mX3e7FCJ0NRc4SmbCJ9GstWfkKHg0wLtbfZh1QXkJjI5G3LL3L5DjhvB8OFJqBPiGpIJnfErenIN
e84XXuIpjpMJxREFT5Oor7TuExEO3UlE2n8c2rDzG9qTpZMyvUH83hT1RZX1xBivUkRUrTqW4We8
VlcR2Ta0gZn2o1HxVoKHBX2sVvJKq9lMYizhRjTLeZLVNF/itGDSe/ew4Meur16R9cadFG2IyevB
hACwZB8Lslc3eMnIlmWKkDf81z39TWLi9JVdu89n03T9TmWR1TmJraZOn8Xqlbpde54F1r8eQ1v5
ugmQAAaMTJ0Qja+W42PMVgPIgg7OlVFaLubE1HgcTmJlWCJImF7nXtF9QIHAUvQ9F82XCYUwCuG8
jBcp4tWl1CdCjgOwpu3oRKRnlcpXBjUpqDkjmsAQUTpGmU6a/4xK9ulW/UvIzvEm9xYZzzgs7eVe
Okv9kK/fxjS5Bz/dHx+chy+a90e++Tkg2/9pt+6k07p/SEEcdyB7HP8Q1zJJzJbSPUOit21HnJ/s
f4GoFRByW6MxQo3b4m3eBiLE2vs123PxuIAWDIwP5qvTaeaiKTnjRD7Ly4KLwZy7jqT1wPYJI4D8
Xeij4Gg/W+rrHv4bfmNokOc+RtYaBL0idsytXUuVlgcNchkEJIYlOXH5f5cK2sZl6w8oa6x4QSZI
iVbLqedWv6DhFv6qqkygXDDQispc4zC1eTBb93Zei6rj9FJUuaqI6sv8XjbueAipzDYVQrVT/N3o
mDyiBMsFEvJb+XqkHUQckS9yM5vuNdgEJLlR81jpDAOtzXwp1qre7NscEcFlRh10pjQm/B/wxbrJ
m7WOMigOArIAx0twpOmv5AopQjp8V4gCifgbKeKcMABXaLDaTAI6qdAVcquj+aOrLoCdmtaI1N6y
A8VTYzS2Ej46qUCIeYmuRzYb9JFyDi6a+oqccipmTMUhOozLKO84FTH1I2fBgb6FDDQzpXSDcM3y
pWwe/8CMXM5/dUNSnEosGBD5ZxC7ijwk+fkl+IBA9ra2VW57cIRl0rBobN6pEcy8SrORvPa2i8/7
dViYwhuFAegWpT9+UCJwAxJZy3/wncBmnw/MfHtwHRRhYAytkzRIlj8g0ZC7vEtEsLkYaAz2B8rT
4+xZNFv2AkG58Yh7q2LUDQrWqLPJ/6d0QZYqwC0YHgGPK5aLMcG0mUmEX6WMkxlGLe+ZNj8qa38t
37zsQs90U+nmDxapOXG9T07mvMZegXVJfV2d0F+U32ZcwckXXiUTVYTB6P2/brj2cI6XZQNaVfwe
60okhyjTWbiboMEJ9wWT4dWkDlbH9FcAJZrulYAdKjTWDzNlSygqtzvZzKlbDyZG6xlwtU2OKTIL
xLuyiB6PAc+wmeaIEY9rIgIw1f1rhd1P/8ON+O1spzvcTHeZIiPp5/duD1YNq4bzlpmrMn7LZdxS
vJHNTk0XESeMHJ7lVIGXveSs1RjFQbLRUOeC06y4qKLLS+EZDVQyjHIBjf0mLpj12EJURNRyHjp5
sE7xBGz/hIcgi13vAULe1afPq9ys0U6ndGBNoX81IGPM/Dupogye20AZm4IAYbQze+pIfxgggwPK
XV+6s7rxirDwCk5ia8dERNXR16nqEcfzQeLjYzx5DwxH/AFWDBcAyEhejM0RffIJclqixBmrtBEY
SXxbG5HCj5GS2NLDqDvMy22tWqLOeerUsgt0r1dEMRuk6PstxZcl1pWD72cJrorxA8j4x22U9+AU
l+pDEr59U5IDZO0ycfPO9iDHCltMaX+oJEy13WF/4O1yduVVdIeO2S0BaVQYCpHo3CV1cuSOmjzt
cAaguXV+qK2TBs19ZZcfYrrdzO0UNDS0fpdLqZeXGJMlZkIEVTyXKZqWWRgspJxJfCshs+9KXNOd
YUbUOmwR+g5mM/GF9XtjiWq94rOMRiihuZ91DdMZs7spVchZEfGO4GSlmXCING5EtGp2fLRtaHLP
+YCKaL6l6sjs6VaqAycglrQC3zyWwq4yp8ZKbd/yDW93vnjrQU7PM9Jx1a8RFeik/cXiqIRSYQvQ
xDD801EqWGewJ5qoEKUMykG/TFxrn6AtFft1zcuErzK/ajS4bCA4OnkPXfUJGJ48BojefqccWAEF
0cbfoCI+9tlU9BCYpKVd/ewX6Db3tSPdtV8UQpEH1lvplDw8ZP5yANxvwCSYjPMIIDi5Dzr1VotY
/EWlKeSRUQk+B4LFoy0wfTX/nRS97Rs1EB9lu8rBEDHxTNSjufHD8RQZ5/4q4u9rqF5rjuGvJ6dl
10eC8HZwiQsUgAnJuBiBmjc3uc/0WTwI6wyX9s/HXhhbB3UgeqJKxZslHpyd9x9Oz+GNpBeAaz31
zTcWuWRkTsj+zV5P9e7KemigHKrAQoR/kOYtXWjO6HX2Ox9DlHTeUNVEy20kDLer6KBXjSWtvBaW
Z8x7SW5RqhXiywI1qqc9+9XVtawloZgVmJSRFkDbOTz+27t9eS5sQhPUqbsZe+q47cKJ7ggELVuT
CG/3XPxDeCUrk+G7Y903NwfP+92gRheuoDvmLEAsp4rg+t8ROdorbF3xmbWiTMhzkWA3XSKzAvfG
BDTUg+c5hRKGt/3drnmkETMRCfrycM7BFR5m5yT3Xb6m1+yCY1K8ihUrJt9QZ2DQQ00KkVw9XA/z
I2xlemih54BnlqVQLWl1m94/Kzplz338wHJhAxFnOyWoAGcOQlvCeiaxieFsNoj5+jM/te5ATCSi
iIBu7HqwDOy9+Ebaq9QtGHBNC6GA7S3rqkTPWI0blOwvArUTrx2CnabwuI2SIuzH8aEjv0pJVVol
cGMf8OYOao1g9HyXTwtZB9BjLKCA7kUeQTXZP1A+E/8OumLYE4kXVgYij4Mr1ZD0KtNEn5O7u9xU
N+D1Imkw64C8L01JqSoWWFa1UjOcdA3ixhivg8ZUncF/fe8ZbGHyocQqkluMNmbUHzGziU59DN9L
7MRkPTI8D44LbAn4isKvzLTApWUBkN0MEmZQKHX/zumDYzlTuqbP+AjbZWi8zDHHEm4l26bxbp/O
9O4DDX4ZaUawaC5nyeR2YBz+RVCVjJcOSNNtLwAnqfMFy2astizBRaYYYF7mfAicmkmiriSHIzvS
/QP/iiimGWxxw9JFddLUvrYKCIGOY4VzdM3/xWDlc6eUwMzAX6QHHcY/NCIB0eA2UkZqNxNt0DS7
udjzRlQlRvQco5qHC4UUX5ExpPzMNR7h/MojDZdbgaUHH5s/Ri8humsvi8xYzpbKj434AP1d+zDq
C5i7H9a1G5j7dOv4mIOy2D39DrsLIYIyIKYv4Oxu34CjySPC3yLtaaEN2qBvAbZlGoYLbFYJazAk
oPLxYhzLXOPjCrS4RJY0LeSQQ9TRYrF3tsrBQIKD7BZWXa/kQYmD81O5xRIWILklE2UMX3qc8ZG9
lC2kNx0H3ES9hkudtn95kLOBI1RSng0pkrcaHzBV5N5GT5s38sR7LMXjqXD2p2Rs2yNgElUIYPrg
KzaR8d1PhXdvfmdSDroIPLr49sZpuvyoHpVhE93Jh4j3kg4yxjhNuWD07/Hd/x71Gdu/5gDLg1GX
vNQfL7r+asGBgTIc/IADIWk1XuHprb/VAd8/Og80QY//YxANAE3FAgnnO2RSF0q26n9WKpzZbaYl
r9xDcSAX/Jm+xBb90z5OTHJ9QEJUABYfJZUubO5C3qznu6j86Klid1DG7mKIt6D/ub2TSqqtIIzY
zj4poRicA7hhaNZdrZBfcss5MoQvFxlk5ncnZUKNm26vuJQdzYW3Iy5qhWwg6LFuhtoVrQm1O3qh
SJxyYn9RakfoqYlSly5+FK7YbOwxVBzEEkCRZmcFvy6HqWpm/ZPhf9fA7IVzWONdkt/y0OigxQ5y
mo4Sv+zIlxHyV0htNutuVvFaN1xP4Q3tvhKXpG1WSzQVVrcnkw5eFN9lKk4TsPDYYiQjPDxgF4PR
U6wuXZzIihWQoAEhJ45BpBvQj++jOfJC0gnkcWZYsrCyRnaxa1I7vrIjomkklGo6ky+ClM8qBNOK
WaSC+L4lECVnN2oRwy5519LLHrZ6WBNxrkp22YVbPf/8rBXw3ApRRJbXvnqHjzDu8LU2z0Q5mZsH
6+BtI4L0gK2ZLbnhBo7CuicfErCsRc/jgt7yY/mPGUizWZrI9aC8XPusTO57/baNg5oov2BybDJh
oBQ3jMhdO6fP2uvy1FY+Y3Vwv/e90R+RsWIkP/fxuSIT632isKw75sgSFddpzt+hm4AY+PLQJW7H
gqj+jOZTyJtqqlcdcK1MfkZDYgwnydWq0rMw1fR3Gm1pNmsGwAhZ0kuXyaEVFCZLWDDUANNG0uLu
kf3xxk+K78N4UNLe3dZ4jUeLwzAXwtBVEquKjauyiU4PnZN4uLMbtVT7BLjDdBsdV+f95XHqauMQ
1JfQy1N+7q2QgoWEC2X639I2isa2jmu50XSozOCpwYiX6ZATi1dktKHBpWWCdmvCJ8VAFTStoIWH
yD+N3mAk3ZVTxLv0DhpxsCeIugCwPiT66M5IkaJPP3IF10BfqfnKkAKUtUOn0a4XkPO30j7XHIXA
AfFvdVfh8kFTj7gAe6Pi0m8GMhAHaNqQhiVYfH5EB8vtaUh+fd1IZ+HYwiJ6R14OWsEZx2XTXrkr
+G7pgBsayqxT/1vF4dnHwedKZ2wEgi3pWWMljlAsM9GCUfuGhp4ivJuN3O3Mrkfl7IalK+9nI7XC
aE7IPG1piR/fb06Ff+D6Pahm25rwiuFRIcezQJIYCdZAwV1lRBlwI8TtF3f2PxSDlpCUC/U7YW60
93JtTf7MQbz9WD8EaWPFpEz2lKXtBwvH1XF8C9sm+PLgI89BxVv3BHVJYztDaFUarqJ6nlaOKQ20
MQ5oHPoaAuz1mEgyCpSxu5qcW36wNCMGlKsYqKGdwzIGQqK5dqQLdIb8bvIUARKkJvW0M3YVSdQc
UaDDkANF53MGo6dFnZGC1AmLo1njUpr+3P9Tilg6J2MQH+MAa7lk0T2pd2OPmmAUQVYeZS3Lxy4/
hVDwwt8cEAxxqPSj8INuAYvooIYRCCgeeVfhoqbTy/nOpQBJ+ZkRNhqvXZ3erCcXzvUmMWmRv9Qq
d3U1oisjqKIyQYnFhwcg0gCBinHoM6DBQM9HzXFeBibG8hcT+W4gO1wRGZ0EQFA83HvekeR5KWN9
X1UBxFK4OvivHZkaulaA/C/u1+vFwUQvuqR+Os9fnmAG28gsqVZyC10i/x9oi+EvYocrSbgANCv0
4W+Dg2DlUxzV+kQjIpduKVecmASWSCKP88WYTShkBHcw+XZv+kb3RNfoGayUpO14/QKxmdOJO7rc
pe0PM2MyljOioi0mhoW+L0IHiFTkfUAxkWYUd+x2TpKx/NKYVu6gF1o5UuXXPWVTy0TuYqnrF8fN
RD8oIjSf20ewJ24bLeewah5dCosZFZX6pcuVTbxw478bVKksZiUX2OFaQtHEWsdQZ/mOaQOJnOQ2
iAb8t5MVvI2WTSZZu9KkNRcbZhZ6yJin5vUCHQVWiKnBGDib3hM++lxlv/Rk89N2wss3RrBly4HB
+poQ3dmmfyNtOozM6oGfp76D8pdHnZrJHJjbdZKE5Y/mP/lsCp6wormDGsISP869TmGgVM6+pJT8
oijzU418zULDIUuumiWhjBxTGVgCpJrC/kME1gooIyE/KFUFZzOzQSwHInBRcSZLUSoQxGpGYNMf
Xe2KbCzmzcXPSL82XbRSKZ70a+D8Nk7pm8C0nJbMTewODmxpjskvbCv+cWVweB7Db3rBU93zO89q
RMo3o/HTJV9Y4bf4t8m5YTtu6z/smqYpFnHMyVuC32RYljTYLm/FMZ8ml/iMcJsCYcaUUEk81C7Q
Qo0jUpBPkViNqfU5K8OlCdI/FiKDynt7PiKqGSmC2hzsDN0z53kPj06zyraXBl9ZpwP9+Ahgc7h5
tGZKqbBTZ9kGW+zuG5DCpoM46luJsIJmaADVZgFlmuUOtcj2V114q2IfSOxE8im2aPFSTZv02U2c
jmjLCFSA9f/SZEtuchy8/C3df4AnIhtc73eHHMFArv8GUjuP+fMPMcTNQyEml9D6RBQYqT/5vA5w
Yz8m+oWZIuyWXuMma+XbUhtNapqwjiOQKgtHYJS2OoghT22YtthLsEF08F3VXG+5zlLk0l7O9X9G
tQxAtDK3aG2sai5ryplqvQMaW2QS/ycOQCy1S2XPJdiZGR1mDEHvSTe82DkMo8AYswqAEBIqswwh
7nhyP6a5cvTQGnockx+WdmyNG3bIWFbkdpZNpKPjYJb9E/Hmr9URlprNCl4ipug52RF1ftWPLe6+
IRYSNTH7RyBmTLcc3gJhKHEYeJ0+rGwrJGHjkq9NN7IClEO9CkbPHcNyoR2JsQhhJG61dvJu73dT
+VXsrBV5jLOobtdBJQBddgiZx7wjxu57U4D0Cy+4lAh9IMGqBl0++hYvkUkvFMznG2VZ6man31PR
EaRsI1zAQJpGn7ttrtFKiWobvADLgZRAcThlHU9s7GBtrKnDI/SP9UNuSBzy+JpqWAP4Zh+8KKDo
dt0Cq6TcfUoPf8odyypLBUvNfSmmfX71TrTNf4PAe2OMqlDDJB7DJB19tfGW2fkdUarZeVw4Nv/B
TBCkDy7nfUrLKuUXPiHaVRHlTpQWA9m/BxAMPWGr5KGwV+nPUOTJPmszuNSZVN4ZONgnnmyFpEre
gjjAVnRYna5VALnPb/3pDYLtGTmP6aClctdYeZXqkKFhskxwZ3cMBGlV3K22z5G7zK2G2Wpbf+ZQ
8TEDWbZu1ff2bTKqh7V0d5i4JaX9WnMLiKnsnGLX/Y870Ei5hSkpUd5Ft20YkrrvBRHRprgbqOQc
ahMA+8v5cv/4M1h8lD+x75lvfWSBtLc2Sq/EIYOJ+v1/6UPC3hFtZTRyqHL6bmUlReOjM6gX0E71
/En1XqYBbVso8kTW66lOD3Jyi/2wHxsFpCNX5OcmffwSqpeGR84+RW+VbxW7Jya12A7hfcwoMX1l
AJ0JGkiALBEiDHI8unfVdJL2Df+uPiBhhmrRN1lGmgU02a4O8LlUYTEP952q+6MjE0LnxBUw6Hof
5AJtTPH4Vf+IzKu32KgW8xrwUZ1DDMFP0xqZcYxPp8V3GiI5xcixkq0Qq0F8xZMby6MBdeHRQeBV
D1OUzPrnpwWngz6uaTmEpYnAoC7wG1N2GrGAQMKwCN/mPPvLhNzvTsQ6WxJG31xM01gNqcWk3GER
kQwjHC1y2PoUwyy8cL+2t1ZEN4DQ5SV2LyVNao+WkymMbqaruLsS3QlGwr9tw94a60x+hLqVoDFk
RVFbk/wMk8mI+70nuyV6reVWOE6gIAuXEUeNalWPrCSVAlDE6gIbBPJDfRWG7RlhpYjhgJP2PEww
QU2pQA52+TAGUgjnH8aRUyt11zfjj3KoFGraV1NUuROuDGVGDXFMgoIuAjnzkFD6NR3uiGbP/YYe
5NBVFy+EaB16vIcKru9E08ukk5YIM3TJL2mtwtm0inRXQVzUCfeZwNEq0bPVwE8JEWYrjfoqqFZK
cEmzK8iyGJagqC92wpAPWq042dOzMLhABuR+QX6fWxW8DhaB+NMJpLrJw2OdW9/iYNoltnXy++Tm
tBPXR4LHKlQnq3laioHWnfr/g3CUppR9CPmTWWH/7WCQWynD5840drPZBzoqfkMFToMuiAmlxZOd
pBx3SSwq/kt0cwGAzDkfuPaB7sQiA8+8xz97upC3kIryUEpcuUjOddQPHguElH7G5EpQrgwHJqwD
r/wSkM2B7Zd7dZkfTb1yIJymQ5IXL+rl6UnLvBMa1RHTXMlA8ETv8C4xx3lmd5bH3L0cTKq10nM6
Rm8A6RjTuRBk1iPj1wRYd2eGRsYOd6wcMSDFDdEdALE1QFVfstYc6pSWh9Ago2Nff789zTCk1Zdk
imzHcFMC9wqTchee0DoRhXTFVoE8ot/U5Es+znxv2dxjIPdlNu6AthItJ6jy6CfZGnqC6Puu5w9F
cOjF0o1uqTPzZB9Y8lRIRONaIJ7/3omDF5MtViRWYEO1+aMQnkola9Ybj3hrLQwdJJ5oZOt8aVb4
BcZ+LgBkoJa8YYETBlBz4MGf6+nbGu2tIWMPZJepk2Zr8Ld3Afo81J0wT/o1XPXyJ5DjHe6WmGeJ
PJ0pH8VAMtYfC8YSLlzQ0bAt/Uebpo0vcIIuR6cv5EemAzIOR8Q/oNXzM4EX8rdt3ARaORiG5ETx
xoBKhbOad8Xot+djCOskXNW8I+VbF8BfksAfTeCZkgPzSSKPfXeP27XV7RR9XW0wCtyBPvYKrs+0
YXLFwnNz79QlZ0q+GJXomZ7L2J7n1EIjnN31oA/jgYqEwmkt0a1uTScLMlkK19lL3y6TM0uKFLmV
Athg3jWAcBa993pAYZnWQYpu6LC6nGjdPSZH2nMWJVNZsp6out3aG04HlN4nxO9Ex9LzmcATXt+j
OmNRUVdCCbufsp8UvucD20CVpJ+eQONr96atQlbWRpowR8mq5nguzo0KRiGvBvDg2QZOUWDYXo/r
bGHa5YeitB0aE23bvScSrqUY1+scVcWVSbyJROOVni5M4NgG3IzzsVyhJg/0Az1LCRH5rMWyXvVJ
kOUQIqWHV/2TlWF1HttEBT/PrnJsUtRxEv7i7Ja4f8pelsfOF/iROhW7qmkWu3cXlCc0Zaxq1Dnq
+VwUSAiEOVYrutW8nJyMuONrymvAAE4J4GSCRYz3946Fu8A79bIsrXF8409XDGbcTXTNaJp5XMbf
wRReVFC0+whgX0AxH2eyCY4DOuXm9o8jHhAhqpCeusAgGYAvPQop/3B4nuEd8ou9SsP8XtssiD96
0klkgNcprJ9FGG9bdxszyEzh025Azq9WksCZ+XU7t0PXGrlmzBZcy+6YJORhWqqhMEi8swcNwwEM
6JCyWGa61sE5CpFH6c6Sqhfx5nSGybowsdTcUmHncSlz93/8Z7jdBzHd1OKKL4amVL1DT2cdNNm+
mcBM956FtLBmjjZb+JcxYAoREM2Uu6pNQQoIqS4RdyRx6mt3yvc2axz0E7sMERwOFdRrljqsBfEg
PHQP9HtapNkUKw5yBKaN72qSz4XUmevE2YA4DosZCzM8+T3mlWtaiuL+JL3bB5KPnNi08IadclTO
kZrB8opW4q8ayMd+mwmKQLUSHyzVJhHQX+UhuLXocaVrH2RzhULveF8/l66xGALVpDV2aIXdbGJD
GKJymid+MmjcpYP2DR5Uhrn6DMpY2SSlUUn2MsmVQenfkLYjVvIhGFIW4Jfc0GwDq/qQTYPIIkCQ
8+uDeASowPx5UYUo7BoKv821M7LssxJkfTIimEmIzlSybbVUmox8kRRKn5uzSvPhSGmwadw3Zxyt
i/H7f6HrCJ2H7/PLocGFLWnwwjaxsafVy8+hLRp6EWJJG5mhaHWZKrO25dzLGhtuL6ViAdhxFfu+
3IiYQmiMbXM+IAO/HArn2ne49itwzXnYpwNgitgpMdTgqG+jFwpRL1eU1Qpx52btrlq2W/XuHYIm
QCbaFDwiGG+U2M4UMJpZN3u0kcfbNTJY67JWXgrHpeyHzZP9RCCgzd3oYfzDhrqaD5rAu18MKM62
/TBJ39EVEVQQySAu6scqVoleNv7zqxPsH5ipvU5RfIhmVU5dKEIObL58wnAezIB3dBS9gEMzCB5I
mhMZXMlxu6xoKUW/f6aN/3S9reCN/EKAv54MgeRFg6mbje0Nn2WGeXaFb/x8ZCBck6xNPitYxat9
Dh3PL69Al54ePVtrHsJ642frLOWXTT8u2+Vo0NsQowd5+0p0H1BTAeUzGJT8iuzA6wKqSwJqCQLe
PhHe67yLwE+vZM7ThP7WT27d1Bu4ObYE/PwTaWf/mGVjuDFh8XRRn9FXsEp6iYu3864b2K13A6dc
1MdBiqsMvDLs8F6ACKddgEJIu0xF3uKIlI9QDozd9idOOG3VxSgdN4j3a8EMfjx5AUMvzdVa8M/V
d91EdDYKuadG5NE0u2m41gaTueBSiUmlR9Tp/L4y1ZCVfPYwWSX9zIenD1lyjoLKy0mMV7kSBJmH
38bGdiqKOBzTtmgjBL/8t+rUiiCTbROFztsGc0hOmDxDcn+Em4D1tX8u5oJPPXVXh/PCMvSeaNx0
DbYoNfYZQ+rFtB4z53BBx6YWhi4/w90agXaqyuY272G9zS2tiWMWiRm4WJFsq/PtN4+I3hqpOaXB
2iCVQqkjCnxQWJSdkJyM3UInzMWSZKSKnBSPLi9oXnfvHWN/7XSF3kR0P+Hx4zPZFyhO/mForMLT
iGbpPU94wCY/Ow7M1DQAf+9omFiLlY+Fqbu1gvjEB3uHkkgeRqH6YSXeQKPuExKbdPLZHdE4oNOD
lhCxB46kL6Tllim+Be69wsKaggiDiHQrKUlO7Zh8abHTHz9b4XR9qyBZaFFXomn58FzceCwddhdy
VA18Qhi58Q1ao5BluRHMXk7C8Lj4R8JkBoUJSx17Kn9gmK8TDTUQCzlN7aovKDY5gGh3k3rvjaMs
bFVm1fO4LIe2y9dGsCFU4KOc65ep5jlYh1QQId0F2zXP8cteSIxDjl5mBxPGZW+Id+eNn3VEehZ2
C+2taIP4MiNFRGsOBCqq9tFsQtgxQbDbI4kG9/xMOE0Q3ErWL/ZX6G+nqvnrxvK+NlPGw1Ehk1W2
U8eX4y/IOdYhjrtS4A2+MwkzSNbjiOZ7x0fy0zsheD/9Hm1QxjkVaq6R3IZ/e1X4x1ivae4YUoAA
V4+OCB11p6IPua1eis/G49xeJcOelwPL96o2TR171eJzcSh+Gml6ruIXFu1hWKhOoHx4LtMchbO+
qcN3qUFRgcm+qrnTHn7m1CcA+rUHDm/qO4QQxmtVTTTiaZ2r9KSOeemnOAU6MgjWbe7y4mlLhXQZ
fI7C8dqlxDSRzlLux6rfj6ZsR+DZ244Lg7QITJdhwgEYd3YFt9lWN+IpCmbuSbFLhfMKLWZfWO5A
/Tix67syCZk7p0QIDcwqZVTpif4tNjvpOehr6ITs/NEUe7k+XY8gk9MWz8HMiz4MsbuG+ZLe6yMo
oG3UizNt1IyyLK5znbcOJ1CI4KF5YcbpsStm/ZvppyZG32GkmkKQBfdixhc+wxb/GD8tQMlzw9mu
jmFT4xd91ptQnF8QGqoY0MrWmf9KZDnceRxEtPF/Ql7WUnL1D3Im0MGxpZ3+gTsh5bifhZmf9MPC
+MJWACUi6EgWUHAyUPlJS/GJjTxh4peF9Kag5Y4FSN5LJY9iPUgpRIb6yUOaMLQga5U5jlBPivKT
Z4B0flLcxzgaKNDcr0RRVMzANxkfDF+OkSbo7UOPGjOnZf1qJuw7mJfvREUFUjhEgsq4XoLCDWG0
ymeqqLLFW3GVZ5CBnfBSD91vv7XuO6LXK3oeZl1T7nEM7xska0abtocgzrtTpt1xugmSsIJC49zf
lf5NxKgojwwdQG+xbEncdulhaGUnBQKswFQ5NgW6rChvs0B9Js8SoajcBI3dxMMGdJ2lkXkMvd6/
RXQKLpyI8I96bnbLWnjUjbP+wacCC2XcEK48WBZGShE/CgH747OB+MNLOgOXF4+cmCYeEMOWPVwh
vsc6c3vFLlL77ZVpvCN803TUwU6c7Rwv/UlDPkFMYIyHyfyhr0dday98Kxf1eau0Zm9I8mwNQYoA
wiI9Qlajb6fXdxMvdO9kcGFdbsmkAS5CPeti74ce13vJ1B8LEIlflnig7aYi9QDEyoLsRUrc2JuE
eDI+KTZAYFLz0PsvTKD+5kmMKhF0x7gtSYBuPUKYAIAzhWV80Hv6j2eyYUXrqVufzq8jqqEMF24H
6RxRH+bwQ8svtpUWtaL887zgusRIthuQTBbcA2i2t02AWjEWfmYRuHpuLJp/IahVooU1afBJwlO1
iiFbgLP9oTEbFqojqhWrgf9TmiL45NrpF8dcL+XvUqI8NDkr+o1fdBE4rdQUbYkKzuY7NeslD9I/
UEnEgx87or4PPVLsHE9vGhiZYGOL0iHaSl5e+xiMvqaUClOmKXJJV+cOMh4Fbu3cWlKQYWtTOJbq
hmB/g+AhXv3+fDite0Jx3e6ntVqZ0JLMmH5ob8fLwv5TVkRcJmFdPv/kwjuG7xOEB6IKQF1/8pRG
vXAYPlG2dEJbl0uldJ84Ehx1MNNli/umusNz8qLOKVZXxKFAdAqir2TVp4hu6u01KgWlRbYJWL8e
pu9cHtFRluv6hY2THNsFC2zRz881XGcecrd9sMPLjrv9RHluXVDHhAiIpebB7+YSsPHweOOY6m8h
46+EijclVg2cpLxcheIdGNO2llPcFmSkAMtlXaClRAWqshVH0K4q1lqr0bcuIHBoux92AraTu5UB
qSjIHaYtaf4jXN/9Wqmt3H7GAvN3kJyFA5tKzp5qNf7k81MAR3zZ+AqXWHAa668bzOEz5R5vpn/9
5mqfN8IgsBUx+4UUbh0hZzmtHYdWUI2L+9zo8bE/E4PjJs+g999VJAtFbCg64Vv3GPip061ZoGZj
L/Umf4nEu3wiIpSLZOjAEWRfxBMDYMBrnpq8tiTVdRpJC/4RM7ssgA0CzoNHzMNDlGr/WeWYXtu5
LgDE1673kIIahoyDAXErp2tSZsyoddwRRS+StZa1wKQ4mudrMIvF2rKgCJy0mZSgEm1NwMOY+CfB
TubMmmZ3f6CRQXMN5YDZLDLiBPdT7gCkD9/5wOAY1YSxz2Sy2E7YZou7myYSl2c/EbDipT41qIOJ
84WBtWg3R/J4Qje2NZ6f6lH09xNL9eTQEZM1GoaNxTNP9sQYWlA1MFGs2uHDxnskBx+9US8nidTD
bTc87iNYlzmXn+YM1c2yuIco7w1fRvGGuyXiIta6XR4cR3M2UlrsbXs0IE/UMZbTsMjX+5d6nSDp
NiaV4UzlHHVOZbGTARoSuBHK0jxrutz8HqOH1cHzv8LIlscaAmKmCw8dhNG1k1d+0XPt9tJtn9/x
nB2Pd5iZhxPGzI3jq2zFfbh16rRExEdrtxDQZektxc8SfdEbihurpOfD640ZVAnjhwQfA1C5QyDm
bH/jrx90Q6U+lQ45MNQFlny5C63JlOVuJ6IlhPDZxIWnA1DQkeY9Cf61a/sL/AmzkywPhaC1bT1U
1ovLC2WrVG9JFI2qOuHD+q3XLiWPY1rXtlXwAiJJzl+nOpDW9q9bRLrFaT3QHSmPa1RKq9kY6TsC
MTs5KBjUJz5eNe34UO9JBe3xw+RiZtA7dEvoTzItckPGpLoSgXnzyfSB4Y/JaXuNZsioyKxFzWup
YREYnOEyzqasK2UyHjGSwQG16HvrfGVxYg2xxkEPXzmSk9WyVBD0Hzvi8hzrt2GaXk/T9IGMva+t
zC4b0eIfRSVt+FF0twB/J9NAtk0/DfkGE6KXcqHj9fCAjvnUXaVvvNZr75rGUPdSlrPyTg1XZTLy
ewCVbkgm4T+cysOeVHHHjTYWZVhLQxWp/iVeuvhvomlpFwObDV4NZ2oT2B0DucPZnwyxEOU29tEB
dT6wuE1XJtLYd8Axlpw2MgvfJs/ApkL3j5oT7HJHwzCmDDz54wuI6vS/r1KRg6wR/gxWVFF8jk06
RPESwN/gu9lUNA5PNuv+iJ3zAYZnW8YwPX1/mnlA2ZJ1A1hxbBKo1Nh8mM0jYBG3JZB8ptXHRYRI
TBiGQkfQA+AgTXO6PFj+86siEX7hW0TsL3Olktayp0KnjJNyeMhSeRa+RxyCxqXEQ8IPlQSHpM5G
rVPCwKVFn2oVjtzdPVUBE9v1XfW1qUAroPM5NZR6+PkZ7f9lOJa4scApsiQkxniO9LGk5U6Fs08u
wg5K7PkoadbfdV9GYbG+9gCP/hJvVxkkE5dST7MHZoWHkY39Qn7aQTHiICmIduVcgPc2IXKl6H2z
Odh1LTMXoBZuIEMxBqkXxH73M05phfVDRHv4lgW4UuCCGBAlTgC7O5hJBFlsW9tpm2RlyV0xB2x/
CHSj5p6UT/yGqUxvVTSQncoAwY7sS7pW1fznSvMHYYRCWhyu50Nd5uyNcVenJpI9dd+xDXWzLQ7v
7jK4wbyh6I/fbQuk6mqcuC+3KNwNirAksVNqkPbHwinegXs/H+AVGLzCvFWsckNN16ehfSvlZ2fs
X316wqZU8woIGxkIW1ozDHNB7ddYmtQ6oRh83p8PMe9dO55X3LolidHkiXdX5B3ESlPS27X8A+JI
Ez87UItKcPvoEMCHNPYzogHSDK7VW1zypt3n/zYFkwzYPcb/UjLF0LAlka5JviOS5BlEktE4Dpph
5nzczXA/RtwkChdCn8p2ul2tm6L97tdM4c39bE3ulU0aA8mMt2bXInKACL+/lhcj5AQ5YqwwJQPf
RmktyfOORynstuYUr2xbg1IDbm15zgjEsfznY/adA3HFXiaEtH9QEXSp+KuVPGhL9z8bM8+vhTGY
PKj3h7W4gywUROZzI98vZmOMu4KXSsxax807zYwzcv6S21IlQg5xXYZbAi80u1B8u6Mmbnumd2HW
3JNpOLKLvWJX6N95v1stjCr0G42cDhu89QbCDkp6J0szyvrl7uC0dMoUyoTvmASLuU2m5dUx4MwS
YUvVHdoUY1oSykUECo8eKS52/T+QRw7C4CVY+IS3Mx9rw5kCuooCjMdzyAp0SUwow9ZW0mLyUXqm
unFNWUVvQHS/vpTRCRaDar8vrUH1h6TNDYavdtZn8cxPGAhxOT3AiU1E5qqMS50tPCtZNE0C6U4d
K7FEuCJ+SJDsqjhsKA5DbjD3Ti17iWvhL3GGVuDmTox1sqn5dabGyiGPUa3DKNImxQ9KUl+OPGDe
78KiVcJk0F91LwEXOUNrfrUwHYepWi6/Fxen//xl2rzfOlwO1w7KOIqfMdiMYB2VXu/70CfwW7Ue
e6AoCoqgLc6Q54tKO7sAa2gvNmbSwRTr36Y9E0iD608bufsuPznIanhhHm3up1IqJSTEwajOBS7Z
q8u/+HBqlBc5xVSiH02LkHt9aWMX7cvGksbb2kXu5wFE01XDJoCSL1x6tYShnKXeytBsR6FsRrzY
aJiQZQHPjFaC2SWv7x2QgOSYKFVRJbdkghfqGcuT6WJvCAYMiIQjMgjd1YdJOzZhn2aqc3RnYoXO
LrO8DjgfEJseWiB8rvbriMc18nLQwFxwggPoRDdl4ssJfaO09WgbiYD3vVNOBlc/SLdSUWZ09a/r
NEJEGoEOybf7Mt02nJyskbnuiUO60iwRdbP2hS9DH1XZiqoHHrzHd0TmiU7vTqZnAV0GDabyen/8
2rcJe4zfschm49yeR8pLW/76ZB9PBUwkvphfR9jsp4iLK7mQI86EyVocRxvLrGUHiKBCCMT58cxt
/a4oc12LHjclrtlzhrjs4KNN6IfNZ8TPEKfn4fXXDCWeSQ6xiMxi3TXOnusAm9N5TbHrCU1mtTtk
6VG6a0TQ7v3pMFrjVhNNXDFELQaVI7lqbNk+aqcBnBi4jvS9Wf4hcInONK/9Tnbbofp52Sxnwj96
24CJz2ng423Qo6wD9X0c0NEx2kwLcZluyCg6yLnvLtBaVY/nmiWWx4ij+NWBiOCdcnGOTqQ9FpY/
tWuIFNLWocXD03bf+E/vbZt8Vyw9VJXEjFej44XrXKse8GUGziaQIC94vjJegHLPlYh4UwyXNhTJ
jBMDvoB5TzkfxxyJmacwlTCVQ1MCJ2g2SezkGP/vnHR5PSNtqDqUvfrzA8sdzpGwLAF1K8waignY
NgiRmtUWNHMbP6JfRs47Ijp54e1ZIDRVVaUD6weYP12KYlI0MkAeUnnNEfvgdTg4i53ERK1DpHQ4
SsUv1OLtt5eAn2OMzYX83pN7XZJh8Bn7Si7h7ZDD8bv1qARK2SJTLhD77WNbvwzmITFPwZC76an6
AnNTO0H8NmlSDF+tRXd1VVIe3tghWl/wjQUpwhhcr+iBICicab/OygvRmnIbLzOuXSnw73SxkIne
4hA+upaqrwrQHSj2rOEDBYVx1VCQTSXGbIY+m00gsyWFT9dvituf4eSLul9j/s8l9pMRXq9IUxTn
5YKdGZvBvT8BfNxik+SJKUGzuUr3L20X5O7gQkzF1L0FsDdF4hUL45iQgRO8n2bYyiH9w4wDWcNs
HA1rbN0E8raJA6oRANuItUGIdTdi6aTfFd7ZajKE4WMjhXcWEpjErXtkKIORi5UB7SZZer4SwghD
4SwjeQfxLknowoWfc0RDvlh6/4FLEz6kGLIy/QsRKp5FyCCgrVikq7t7jLJEFpi7g0f6V18Kt1nc
VAZVdavJY1bjXlk4xrgvwVTZKx0wTLzlefZiTFB4q+Lnz56uH9AfBwZqHBaWJoS6fy+le8JWyKw7
BPaP5Bfz9GOgJXBEfMtmEei26uCMFsO0JueWOECRgBRAAcRcnbot/Y70CTtjxWC1yVH167Sicvfe
cUMwRTGO3Y/6W7+SFmREdnWVUwer6q3g8x68rhnDkjpd0KAHcuoZUlqB+74lzJb5mAtEl4Uq9DT4
z2kSoDGpK6j/YVMjFtTe4L6ItekoIQer/nN3O7MB6ni2KPRRNyl7OXKCQMbfVNeOP3iLoz7Tisjs
XqW8lao0J70MCzB29rzz5CC5mvODaH2CXQmMPLU8Nbw95k2uBGx1laOZCD3E/OkjTiogeA0+49x5
Fonn6VL+zqvny1QN8N+Ur0wIaAmxNjL+J5qR8oIItdloNW0r/5GpNQWUNKwnYBcIBJJHvVbSyzVr
k4K27YUPwYQDD9XGCzTUdmHc7Nz/MdydzmA6fG8s6eONXRwUyfov/TgHxAJXANE48V0Yh38jkjTC
84S+THEZRs/6vzGfgD1WrXmiEab6B4YTSjQ/Ae/DfFWswgsR/dkDgljN5b+wQbFNEseFYhdkz3d7
LvxpXSr/EC49wGjDlQmCwTXc6ed6ypnPgkM1OI1mEq1SBjxoV99vpw4D1lYaZ9tKLVih7S0S26VQ
hmUQYY9P/lYKm0HFYLg8gnXf1FlKbYtxrVw2H4dJxbnNHj2lfxylBKIXfx+UsAiESorz1fKvEe3V
6xd0zSaAK3nEfFEFWNsDf6DMLCT8qohYGjpMOZ7SACS7iW0c1x7rQGqh8DWNS21aKDkWE/8V91Bt
+7iSsVRoBQ7ImR5wa9UWpeYP04cxEqS37L1gtqhGVXW0ahkGrBNzJnkdqb5gHAOqyQ/rFeT5wKv6
dxsN086uJ+5gXpu26dHXn6dGxsQxW0FGygJrALKqsMqn+P9MMa5aaA4SjEYDg5XXlB1H1LnhTCBg
pUOMrGUWutPbDJYtW7zzHYGt5sWlCpJ6ky9ExPLHJuxW4bphKXF5i79Urrmv9OoDrv13OxqYFFH/
GTAt60uH6N9f7fOs3NTdf0oGi4DQrjuxiqWePNIn6MwNp4BvPnqUeWV200MT1UO9w5tb9flT8u8+
QPMSd3UE9VfcYykQE48sgenVmQIWETyojhTEA8DmnbWwakjUPaEfz80DLakrycT0hjLZ0xFL3Qm/
vXLAJv7tT7PCeyrugVFXonXqkd5/4jc6FBuQDc10M4bMtAXakttzEDseCksuRXiZ+D2OzWfZKP6/
/A1f6PWa84FBFLGOnQYE1pcke6SSLE62Whc0jmp2DFV574BeULBmp8FAe5rNEyXEADc7BUqtSscV
KCE7TkENy9o5uHipmEdGNXKwaF6jQJUK2taQEJ8OZkPri9hq15T0pD9WSPuSTdghOjCOW5pWwQcN
6jxgp6ss5dMQM38oSOLm89uQCZhhh/g6/UYGiCzfJG+0lowokzu+8m8oQpgGjC9qtzcADaypE+z6
E1OxFBco8e5xxSqt2CE7k9NaEwSa3lW4LVe8cOz/1JltvE2188wVGr5RF0qrhbwQoEvCWlPO2dxa
dP5ZfQg92+meoR9ejI5EvrfkyBG3zFUEMsnFFY0vH52u8KeHUqpJIY2a2Gxnw2Pdo3aJa3KXQ9oT
tohGaLlaqb28+zLVmAtiUfM+jRFDJ6UPGFjdzCmqVCYikdIl7j5eq6WlHIZNWlknXHZcwLcNDdpw
kB/saHQmPPiRrvNHJa5p7x751O/ACGJUmq55ewvwL4wzT9OYoPVXqxo8jYm3GbFG2w1eYLWhwdgs
eCjINR6gIOmj+n0Mcmez0liqEgeg3Dp5KUmmD+cHm10LS3ycPRzgp1VsPVE9lFvqjXQUPWWFCLlV
OxqtK1vzg95GTaUoWcCPT8mX77icmlZzxwzBlo+urdhXSc1xvtVZd/N1Uwm841NcXke6+XkykIud
L5j+/maKVpa2NCjGATgZulqxB1vpVyJ/e6gWzBnD8B4VwQ3WHgq+ZfXL2Zb68lFA8eBNOVuZaYXd
6sPbJt8W0UCl3oHRzG7nRHoNpm8+dNlvmhEBx/o6Oy5+FzIKoyBUN15/V9tG4uSLJ+MIafmCeXFP
y29UsHsGiTAgKmH2RWV3NpDzHijjMiVF81Cmq6e6GyOBTtbExvHsYdP0+21lOoRcIsOUFOnaN3rD
WWX4zFGwYEKz8WFXnGs/p+s9Qt7DtzQ7ZY6NX8Uz2fkGbvJX4stf26lgfj0z8rpoB7G5HJPdncxv
a2FPV6yO8l7eIVEOmQYH/wkuYbnrirou8lcQx+MOFKv4nfQfO/5uSzjJcpw/aIpFxxUoM7nGGYDe
xeCuq8w/nJGjuVrmbIknsMFhQDEiEYFUWI7fvk/7I/T8aQFIrjeI4OxT2JToNrsYilkQF8bjpwwc
il0DJR3C7oQakBW3Oar2VR+SZ3jUOIj6QIt6vKtX9FSus/PjWWKmP1aKjtI5hiWKMdFNfyi3NCE2
Oob4UqAYsXsVPhpFkeW+3lfVQq29cirkzZu8goC59p8V16qMSZPfLQDghZCJg4rI+nYt8e2mJrvH
PkR9aPgaKWP/Zc9yzLb31VyF++LTOMb/tqwKQ7NcuraYexZWt4roLAoMwRUHMPlghm3dxZwCClq3
QqSOKoyLtDHQyfZ3jyxZQr1A04SNfQVlFcKGdW9fM0N3G9BkuH4Ol4hwoKZ0kljbDG2GPxOZ9ApP
wIDMUkhl2WU/GrkIBUotYWdbW1xzfeAsyNnBkmzcUOAPHXlBXohJsmTPDlU+ZtDRRXBQ7kOFAYcg
dxL0qrNywLIKMvocHgQoMfJ9o+HMuV9pmtSLS0OU/7PASiQrSC28aKnDsn+htO7v7O061gJFOG+/
5HA4r/gl3v5yA0he1VTQTJkGMsFxjz5rClvzT1tWUTFVwgJq5q/KkeZdQ9uRxNNt4dX+zDWjxiMe
m3BJf1KKk94XDASYuhLZH4F8xiqUTKucnPpi65I1YzqWpbMmc1QKKuNtcnEQRxsSjTx5LnzRhrFF
zuQWf2e/DcKL92a5bg3P2h5Wz6BKlMyNoohGonfnT6UUVYA10pi/1LxWTvkLyrcjELPGdrsjCxzr
4pgZz9d8k257dffVFBTCYrAcLmYcLJiluP23ucch34/1Cwrd9/RTE6fKMHWvyiZJKWyQWt6eqyt8
HDAZHEss9eadfLXgybgFeOBT7005LJxbOUMtRprsCrYWQOCxYDYHjtih50mxS8D6RVc5sy4eUyiX
547YIr4vqh4iSVXCeVdwyJQkWNdxRpdTYE7sfksfIdz/m9NWS4pDB+bDs3eCeFqpVQpXaWiWE7SN
x2DBY3UFl6xlqeEqLkL45DtymPK5ZaZMSZufv0E2sV8Yfi84wES4m7oTEdhBv2pC8oria9w7w4WC
y45UW7SKBqWkfDpJNxQ+r+1RV8mVLbfZr6IXEjomG+YWfQSBk6PbJb9WzwM1K2vuYoTrFy/YnYyo
hbqsMNUdTsHfCX86bXvLOPWUje0UMRzrhRq2khv31ZNumQogjril70yHYgxswvb8KF7rBCPLCf2s
zpm7kw52ZLJ946Ys2skmJwWNxmRmMqdkM+mhLcPDjdWqh4p/TRdnv7W6zqOtKW7csdWJqihJjug2
GRNK9qv2LbgVy8I2Nwdn3Edp2lIvhj4DkCUPZJHbhr+neqm2Ynp/1v95ktr4KkXqfHsch19ZjBDf
bg209cf2J+6CCvnc98oZ58V7lQqPYAbZmkzHwVy04ZxVNIFBjfSutjZx6JAnjkIl3cOBeBxT9wVI
c1Gqwt9ntzTZiOSfWHuslB+sk7n1botPzXUjyMtMwkkqtprCXQnTYSqKJkgwu3GYM0RGuVYyV7p8
dfPXTdeDAKHkCgCputM6h6hibwE0cZ9hbpGpqzgl+u90Gs/d3eRz+usjnor9DFustj0M77pxzsvb
37PkrsYKRvsll9J7lDomWl8aPqjwYSkBJ+BtKkJ1haqa8fuqXpiXKIY74DrgWo+gBOXsEdtA4y6j
5VXhRsaqfcTUYPCig+aG0Y2R8eMjP50Zm5VDgR1wZCmP3NXIoC9buLtNhy+fk3hfje1byNaWLCCH
a0LC/aWplp/kXyBu+YFKna0GzLnqUGFRtRW1+AA72qR83E765W2pRghj9ABtcqngzgnEXefMI+No
te9wuFfVsu4iF/Mmo8HRFjE9YobTEh0ccDdkiuEp8+6ttRwIwh9TxsDUPLX+TIZiL1uJfhW4CrLV
Thm/icw5CDLQ1CCuFNt9JQwVvWUmycf3j92RY6cUNDO3eEtEHDJgnH7KLcCFD/vkT8NqvU5+6gQU
VOdpUUKuZAg95/oYeCQqS9jySOIqRlwMVe1iAgKbkv8bG8DFcNDSrl6O0CSUMyRatlV74scfnS53
8YGkLOkEGdR6EYU7/F2KrF3qQFD78VWiIGnaYnwvaZDqWg9JKNeJ/wiJt/uPsR0fCSqR9fturNpP
5z0R37JleYTpJbj9UTinDTKyE6ifqKZAcXv7b1bROj6oAxgw1wQE6d8YQF2gq5ebXQyMFtNYxOJX
BbVBSylQXaPv2f/4eb/vxCXLpjOje0p6OD9hzGN2D5cAm3oy6qkKQw87Ru7qKayuLptRoG3zV3G7
xWs0aCHo+s9mFA+cKKu1tUj+CFK8xZlZuc6g3MYs3fokCt2WOl0FWAiVIo747VN4ZJRJteh3w6e1
y1IYNHxwvFCRoJICddsQFMGb9NZr6jovCyr0mJLJrJdoVLj6bNnfesgF0BcuryXfQP4z5egRsp79
O8EQmFcqk63iqVwoFzsv288Ev7XJAc0ggILhwh/5qsxeqG1OngxSHPsCbgZFAHUSlpWnWNLlEl5d
WvvOQNDC0c+Ygj0lW4bn8mRx7+hg8exfoBZFRl+BmtqCv2eUgC/ePOTluHDCamrvu+CVOGermlXd
13seG2sYEFyymT+rT4AKgvfVxEiYo8jfv7jnJg0VPZ2SsoP+gX50jPkiAt3zfwAloovBU6p6rkv+
GdBR4Y8cCDZ2pTcHIvQCHuHbDixl2uj5r0C3/WPqirwFeTSbFCph3OyJ8W4x5eAzn/4oJ8D6QyYm
YQ57SZU27ykcKkkzRVydc7spZOwVTlaD01lSufdnUaINGA/2GUnShEyT4LyAuE33Wl+V/aKMJTby
l8wrrbQrAXqDbqFEdD8HSzkN2UqWG/8GmEwNx6BLGG2oYLFe6ihNoLdnFmqz5lL317bVVC1PO/tI
xsdV1RxidblGKRS/iwhuon9jeT7L+KMso5SEvITEFT6R6N/+FPzhJlcOuqA2o5qKJdD5aaBJzbYL
Fi+U0HFkINzNN5sl39UQmSmQkD4y8JSQ+mKTpCNOFBs7KJYmQiadM8xn0/CevjNBWbG9EmCwN8ag
EgF4LgR8eHKJa5EnniMwpnglRaPvu4d8vzXC0+IXFEu+4JagiCdX+5MrA74yt5HYajFCPv6lou/x
x542vp3ba4p9nqJkyF5wccVYBkCWxuIvvJ0PP1pd1olZRCgUMLAnOjSZkD0IG8+cchOQhNk95694
AFbf0vt9ywD6RADs8fy+8ur91+nsNAAZffRmuVskmJD4N4ySQ0+qXDWFprYzd4mOw5zMEushH9wV
cCkhT0wDx4wAaz2w0DR9XQC+EtFxkTY2ELF/sfNX7zprNP9l5cXIQhQX1VzAnzbCMmRmHsCfRsqL
gz3Ivbn9pHoURl00kaWXB+utPuQt2RxH42hQTsJ9ABvW1WG/VggcVkuzJwjCoHD4Eus/ljgYITYn
X6wkrR0nAs/iYCxv7NiJBEUU3cBeFzGKaXhUJqCcLVymgxODMoe40LbcEqu9RiPRT/Ve/rQu0XhO
cWzPHb3e4KN48l0elAzIvney95WXfeYiLQXQ49MVtFHewWm1Jel/fNAAPU45EzqzMqestiqaWBaH
hcAEV6InCxeHQlXkRZ5Abi0yLTLxzAMb4jXM51KsrL6qD1JpsJK2cvcx0c4U1HeeZ7vII+rjuOa6
IdAdWYLwHq32j5Rnvaej+tIAsEPmRq43eXHgALz6/Xk4eMAXMPf/dK0AD0PViRCa3wQjlpc1iYhs
OotKvCbdrEXxZHvyQgSeniNCSbXXwUH3wTWgPuqGJ1mlNRMw+fB/EoxQPhiPTH2/VJPchXjcXd39
8sEtl5LZG7fp0JSVTtkdmtvOQpKNvFN2yF5qLscWbsdROzk0V8hJPyQoCWjl+kQuFW4nUcgqExFO
LozsKOheICL8FiKQytIFcRLbUEmI0zr2zcT0NjnKTYNrC6Wt5jXa8Di0ZUhap1GlPSzrCIElZvS6
8QuAjzss+7TpXOagddUhvFfB4uf3epWykyuNO58j9zs5+c8guxKGp/5xpbh4dFfyA3sdkKstfl8X
RJKpJPjBYhXtLwHyuneP4UvwD+hnjfEgelpP36SBO928EC+aDaXMUdAvYIaou6q6V7tqrdM1RWQe
zbvMD49hrW6nfT9cKToEr0hPCSAU6pzqrhzy/SuwSnqm1Ex9Yi5qJjzzMXbbViSM75MNTAPJBEpS
0LJGDaNPHp+8uD2OTN+/iW0iOGCKg7ps9+hTdTSC5sm0VRAEckJEKM4oHBi6jp7WW6VdtG/dM8KE
tzVDBxqjY7Iwx63aiJ2hZh+6Hwgz0RL6HiciycDW80zVxkF55kTasfwkslrOGjy9hu5Egmw8ZAgy
n8uMTaT8KJhw2W4Va74RWnFzH+QlbcVH76I0J13M/je/W4obkDbe9eFTCyXW5KjaOx+xXOQq7Egw
irzDPdKn9BekWqsbzQpPqDrhlp4v3W8oSe37utseQx59nwCbdVlm63/s32a6iA+ZnR9j2fFkWLks
4tEdYbXhc6dpxuoLQ0M6OmVPGxtFQB7M7/iEUFfTG2a2PWMqA9q80e5J1WfWgRn5XHNdNSZf2DQs
BgdD4Yk+6n8u7GDvxKQy16rI6Z7BJj0gDmi0DHcBpF9kgX5x8B6rmAXCdy7vnnisGrnrOdKQ72UE
8Sb2xmiRUyy1TRiDbHIpeALdcQ0KLm+rAdnEFuQH0clZuhGKFu0rOguABvJi4wEcuQLPV/avneL/
zloAlB3wudEuAAE9WD3Er2J9tP4C3+4PPwLuhOZ8dFRxLhzx+B1Sugt8Jr4x78/iw3uFrjVvMFXs
3nD0fq2+hPUZMMRZVtEkH2R+taNH80HtATtzCbLmd4t6m5p2rbVwVYnU8YvBNzidxZfov3ZxbZGS
uYU0XSRB81wNMMVOeJLl0aVOUbdFQ9Js/qYVEHtoQ8h/JflQN5CIiZqAiGHmWh+xqxaOJNd/Qee/
igPiZv53JzJgbx6z/EbBewFMcAaCDvT8o+7JfS1eKQ0fts0LXijzUnG87FKiQWZ0hDAc3aW24JKp
y4sSyKsZWmXZW5jMmI905CQQCrs8sLJl/ROH6jYGR/ql4Db8wDQoUnptEWNhtIPI7xiO5nn7wri0
6E853RbJYvh1zit3fuU6BJrRsNEjB7zjUTQRv6d7WDGQc77Zph+L06LlOX95Jdz+ih7IcbIkEvok
sDJomlw4LlTsZ9X3/6AWDLrMAbSQMGqeRUA8chXNpQG5PqFzFHHs8FQauq0dcskEBGl+yDz5ULOT
+F6FVR1bOGmS3jX4N9FccgT0FlRsMx8u/agyo3NWSarjh80is39UcuELnuKXJAEmN3yAmkAApJrX
2XNuMuW9U2twkAq9A7yzm9dct+ldyuxmO30mcYNHjDjVR52LSjGnz/284pEFRf8pDt0CrR6zCtu0
LD/bGK8i3tw5FNlLJ+YTaBj+NktlaHZ1Lq+WwmOuk2D9aKArg84Zu6OnmlPMvaF+mb8nZ+79y56g
zt1IiE6gJY173J/jKY4HSA7QZHBMkEfjeOHjZB08AxLY4LcdTLcxIipVUECRGoJgMzhohGBtZTwz
ul38sKv9wXjOOcmSuO8q1oRr0uVlSi9WY6QYqOrKQqUmlbJoNvWWZvmPtEYCRicC/lv7pWTwjZnb
V/3yFdaBr42K3w5wzBfZ8RRPThpW72uyltqc0jcTB1AVtB6y6mSrfoSyuCoGpVPpbaTlRbsbxY4Z
uGXPHPxZFp7lSnwdnTQtlThWN888z57Kcyxofuo1D0gQZHsWOXsuAmAeg/v8trltqCpgunRWcnMK
+FRkZnqa0JNSS3hx8SQ9Fy25HfqfXSllxtq0zCvxwK+s1PxWMla6XHCfVd5Av9JK9BUhSmS8T+IC
BUnVsFbeAoufmYBPuS+ErUsJPYoG3xWW49uE5F9Q0f8R29TGT/9U7xJZwAufFDQ+Jef6BymwnakK
/ZqLQUiYOASs5GwrLDfhE1NnzV8bDQJYq+0LPZwmLQ4kDBb0nurhCYURrLOUhxyuSWv4R4TDcZyu
XotntRBiXzdBHueeCPHY+Xy5oV1GbNGIS5yMbo7LN8z1Pd6QhadmxKGQr+6296MoMyk0GeLFNIpn
RXnfiNzDyywly/D5/a1q1Z2H2kuocpLNaUdCaiImyhlXOLs3kupXCv9IpAcj6tBab0kw18nCAkSz
7LJb7zcznc8HdVdCxervwzl4bKN23mem/NSxqz3ZhIfgCQzav6uYR+3MSuUz+8PizICAW1TmuXUI
sT9PznyRrQUYwaC5aJk7B5MqyjWouKlGGazv/mYryHyCz+qphABoB3tXq4A9hSpU3/HeOoh+7hGm
WeK+/lyswSjrnFWzfXPWB+h73TwJks6JjMRU5nhpKdwhP5omfyKzimWR09xmHgaUU34mGvj3ENyx
dmbG98fKtRe6XQgYglAH0n0xmVurEG7VchzzanUxFwym6VdIZ3qIuoBSTU5p5k4QXiXIXRhwQZeh
QZlRHQhkfourD01YpxSHjtjrjJHjL+uQuLzFdsFD1RRUc5m1jZBuICyAiQnaX58n8CP/NMt2eY4b
PbVOU6iPB/3WiuRF7fEo+5xUnDKGP4EJFqz8M1ZpjnP2xshOolx8DKwPtt6Feeu6gQ/K2FHpCNrY
fCeS1TBdD6PeMNcb8qDCS8tMF5Na6g2i7LbYU6VFAfJtEyTvnmB24aIeQ62/sDn/Nd9J+QzzZ1vE
0F7rpIrDoQt408jndEEc5kxeMUYiPOouv26jdQounBD0nZM25YFNiTDeHScgQSUroUDdHktoevyP
nFjQMiMzGwxERjLt6dfwpQLxrDLDA/EHy4OHyu8GGc7U/q4LPvFd3holN8aj92MdBX1eLSgyoCIF
ztpeMi5YcjdUZxrOf0K203BKHg6lLc0MiEMcXn4NQSRiv5JexN4AHNEYSE5sVpZXntP1lKJPQ+Xg
ifvvzMKvRdoDN8k6R9++QX3ENfGuRyZEzN13Lk9ijpDYhcB7PxgGzN/OBt5X4X1TuuvOdHT386bS
pRQDLL/zP48q/KTMpftuYLGSO6IY8NLpijFmZ9auZ++L1+pPaWTk6lBxd1Knin+MenfI93wNiTL3
d+QHIaIT34wlgkcvKuONnN/2hNQtAKoZJE4jF3BYbB9JUAcgDP2ryieP8q21UwIraRrUDhNpzQuZ
rdUd4ejifKP2eHnuGKS/4m7THLFXSBELoMURL9wcy5jaWCvI2gzTVGEeA67+0r+zpLuctw3AVuq3
vpjajKyjdR8Hw1Bv+X3FJfiiaqwtiBI42+YBIvA3Mx+58sSPWTCLokpHxK9fFTOsPyyLxeEtLWR1
/Mt8l8mEXq52qGeUcwJ+GVnIfCt1BUl6yeWL2+ubC/8itp++Rqz5C4QQS/U/V/26Jyo7GrSpukCf
h9wiz08ogQlFuRfePQJK8IxJwEOpINFVwuOzfrbXGTSn+ry3y99D+X1Udqr+9RqMk9P/+/xNB+tq
fxz5ZFiNBa+2xwSQG3h+Q47S0BRNmozcOyd+s35lXvHWqv8bVhDFcfwvwaxqvAqOfP1Odd3fD9Sh
EXMryv7XG51EVdZgJhIyUyRCEuspQFli8749/lC+QEN26b4dVIkTSPhaUbXKBoVkc+xZd9rzfdj1
3zF4G3+esBEIr1fFtlkLlmxusVreu6SC1cfUiexr+Rqg2czOrMt5lAXRyIaJdxTx+uNzSjdVCZ05
zhYYbCfkx2VyzEJlIAJsSELLYA8sh6QFcChSdMyhLZgW8KKO0VKDNbuL+FXV4M/UyPekyAlisAwM
Xh3earKGTZ8mOixvFSELdOzhrbK5vaU5fKuNZuFWD2SAnObGJ/OAoKhcARZUTBM6gk80Ko5R1Xlt
3PDjtae1pHkELnoARixMOYrHCIA2suLvpCxGMzu0ch2v1os6B/8ts4Lq4PsKnV+qJ0L9pZqBkFoj
MEfAKkyteXoVH6LEij/AU24FqkVH4s8WBvHIqkLQqkkBA/vNDBtEO1P4Dw29fzqOYU+zf1Jqb1vW
XPXcY9FOYwEic9TjH7ciogSUChTr2v3MYFY4DEWERVQpYCF5rzXRzfJmvCZAY4zQXePkinxIxZje
09wszOjPtvDCtMJ8Wq56UB0q2DUc4wVZa7Tmg+JK8ppzIWTf2f7ddrcK0cRdDZ3BjOPaQryWJL3r
SUQFfK++8TyX6reyarduzagquj6qR7yxl1rHPaxDoRZPUyYGsizo7YhGhy84TmHNck6XTJKRK3kA
74V+0488NVAia23NmzWD0jxi2WsxlReUfbwgI3eEAzyA52jeTswK6F9J8Kd8+U4J4ccHNqOeT/wa
jqppCHTsrVPQ7X/PMRUWxaMg67C74O/tWMgTdHFO6bGPvpgi99T8c7gAB93cuLdCOC+5VNM9gzWM
NcYFjgDmLeww1GvWotSHyf2cpHSuVMUv+GBygnmQvaO9UHzfw0v6mhMnAfZsChggIUJ9tSjLkR0d
P/JV47eF5Y0ol/G9od+K+XJIiDAEKZLDuZ3xqQwHV1q2XMD4yFhB3z1HHmd0/C3oG1YbdDCB0YGs
IaEfn5PT+wnrEABVMKc1ARfCmMyJzOBF6fM8HRkWln2AQ7iYH9AjPswDA2iWrCDTXqbHvEVsMTCo
wJkeCNMpKV7LqZgx7F/pBB6h2ZjywFYY0UXx8p1miS9/csdmxm4zvaq4PKQuiE6tSm/RXpPVWPJ+
xTDk1bRVUdWJ8hePsFdgG9LUMuUEmrp5uqM2iI5XPOaczP6dAtD4+OAlhv1Vhca8F3ebchexKJut
UfxqCcuMgXQahltXh2FwUyKA1pskChZDmSpW2Xmm6cqlDCA8V2+/29dfy0NmqokY6II/im3P2c3Q
/kqFhBqiGugM19pF2EMNABz/KTagKyqPeByTOYtX+iXHZiysmBGT14V3o58TPg4cSVlzWxyrVcQH
Jvil2tzTvZ3Gyrt+yBrAGLcTUhC8gIUSlVGc4dHzL1niAEgf7K11k26UTgS5AxGDh1NvBB380CAq
peEKTOFKI5kJv+Ze/MJ9Q2tLUQ2dBW+c4KhXHdWp3CglYj1o3n7LvPxVvhj1uIpV0UmjEm/vLk1I
Awp8bJBh5cXqFuIeToaRv/hBbBYaYbooIC4gG3OEf7q75yMX6yBMiQf0RIPtwlyu29rKWeZ5u81a
ZJh8aIdZmumRzNkhWqjZUuyRzes3XqJviWCSe5uCVtvMQFnNwNpVL5U46jmIewlDYOa+2P1zzvhk
wc+zUl4itpW3ewYrF37GTj+ANM5ls6dvpdhI3CilWGDjNWpIVH8tTWDb2ogRkbH/1HcKT2v+LjrI
RLApZ/dVNFaHMrZ/Yf7IB0b7hzID71ANj/3f7npoQmsjSjOZ3CfVCSU6W8EdUiHmfO6wmisp/mBT
MDMXEFOATxdyrqm7TLzQrjzzuCNGbmbZTKLRrGN3TNzA0jptH85WxgmuguuVl5qaEK3AVPV+NA/8
HdpguuGIo8bYgP+IbNkBeK7OshtQpq6NemHTnuMz/Df/PXKKe0p+/K9FdmgMue1sz2+H9MU/j0i8
bTdLYMUD5sQpKYdbcZ4uLUnfKBayIAxU4unTEDsNNsjAHTH9ktqYRHp4g82faYlv0znPCL7V1hAL
dNHQy2WS5kolhGJE1qv3NkgkM5mnjOTIFlqpNp2cXrenrRTX34nHqckk6lC9gfrUdFkQeBwHk3lg
ce58XUXpjvg7mrJzuH/UbGJ/yQ4oZPYxsz95PioXp5GtzYRPggTNYudp60QoDuuzFuNUF5VDc4P2
yDyUpunrbJQKGEMJ51wcnDEjaavtnu7T4RqA7ErslUA6TtxpPM9x0RsLsjNqNukl/PBBIlCzTxzs
ppvGEuvqFqY0g0B/d/rQ9XLixNezyQyKrzS6gcJPlBZA/N1GzNSIZw1fMf69HLm5/7svkXJdqS64
nfB5t/t02aEI+zStJ4a4gDa7wndI+ROvFwf076Lp8Vkm9QkndpUx5i0zCQGxQX96NQk9LGuIdYOw
6ktvT9icHdSIffsD6xmuKB3Nb3w8lDwUOu6BaxjyMb8OvBu/Nuwtkssp6VkUl0R1wT1+MA5HA7DQ
NAMKxWEyvVji/VsZ3houoaFnPwk/b7MP4mLjTBEGz0SrVaJ//nJYHMONYJB8yr1GV+f6xE+GmVO5
zD7/gcNFVLg3+Pzh2Hi0YXddsos17edJv/5/gTLN1WgLLnGjQIlhOrL3kaDfdgYsHz29ojXhhACX
kAJQk6HvEixSY29PHvnKhlWFSV9Og6EV1MXvHhcqg+HrUKW86arIwqSR1xVOfCIGM6QGDGK2hBvw
Owk2eYvcTFH0jyfwLv3+SvMxQ1+nWt0/Ff0zH1INxVTh06ltN8LGSJYwVng0ewSD6HKgh+qqlggw
vFmKZd6aIeyhc16au8PD8MHaxocTeOoZ/X2x7WNyIhJdANOUV1fLQ1OYS3g4v33NMtSiJ6zVxh81
bz10KCDrVQUpMEl3tf9WlyJXJxz68BbcZG8o31bmzER0FxzScYPIiJ3KQtz2bPM19n2vIM6F1JKs
nbc0n12SpUJ27W7iqpBN2mnaMPv+q+q6oDgHCXrrjtqzYqb8iTH2vk1aRTGFJL0evEzeInd4TfvU
ZCML1kNAvrNZIWMcRhjNDaYnuUiw3+nNHUGKg4asmzQOfYiOaZhSbK07bSRDd9K1e1RCydxItrSJ
J4KirV9kPbZ08Q8ONlUVRXieHWv2kKJ08mJneW8JSNgLQc09zZQjJaWF6KURH9z1C5Qz4BMlCB5l
Zu4TGDEGp2snXuTO5Mhxu12WoMX2RG7Ohmj3rzSx0ApNvi6ow+IoCEihlfT0zrWRKFVqf9ubGiDg
JgVwtBNQ+it2QQDpBbtdojL2JZF1CTHxBYm7fBvpDiesseFqMKinRqdn1DXrXgvMlBw+lDczy5zc
Kja4RXPfaRCFr4pDyhYtlWhbfXmJ/gw8gnx/bTNLBT605XhjOzTqzpJrHc7RaPco67Ul0FzHqVrr
JKm5GEiD9jWDyWl6hvOPQSVmszzTfsxAWX+FE11lp48+Gqj2Gpinqui0sEHsfnPtxhTOyipV3ehO
WBJ8UTMoV49TDvbJWovMWUODFWIKpFgH4FffCIJ82u2EJEfj3gWen3QYOI9YGMFgStS8RX+F6q2x
mk4EXQMEICoqBbd7UQivfRMHiCUm10UhavsanVECSzqbD1wxVaHsHZhvv/0bF8QSCY1WLGeVqqtw
eXVT0TZBvxrCDqq+yu2/LiUzbFXsaybbQk1ksp14cyRFYXtUW3k4PqStiC0FM8chOSUK1SWao+aG
x+78D6xLLdMKq3RGyCAFWRyI7vCuH/95EJ+oDfb31VHdR/B5zy3920swt2mmiXtCyaNOBy5qc2/9
zVqLoQHzF+R6MO7YYtX1QfSr7J7sn8s/yv/sSAFEE7xK7Y4r4Qg9N2unUZY+FwzXDgxUBpIYQKcd
bnjd+fz55PCB+UxTL9XpWk8w8KSzgzfJ9McNP1D4l+DOwsG/njE7MkkqcYe427MC5huXsnkwU0eW
qEpZY7aQQJYsn0Pwj+2l4GwHvfwv0lic1vK+H1bS2OYpPHfP597LfCj2/o/ufozB1oEHGt+C8B4T
+8uxzmZfZ1KSXsk4ceSXSnIcMTSrr4L6+4UzChoUtVTqMk5XxwjZTtTMaac6DxkmyZ9dy0GEPXQ+
uQCMKXbOjGf/gAHrdXqEG1XS1Zj1y2T0IZXvCtTCs7KdaIFurlgWWPF+K5KKbGl+vnsm+J5gen7f
Vgag+ZSpUKKWAymJCzPE8k+l6g3NsNxx7X8uXPD9SEEXMLAypQhGtbtBbNTO/msgrY46GwnbCPCX
Vmv38PnGwXZIR1+y31G5MRUuEe1MTBn+zZYsBp+AB5eR7CltM23AuV0Wp4gi70yusBTDU2uP8lFh
bklAqTKI+lSACRXZbsgUH7wytcWzMJ/Z13FmzQPg4mxr+n0XwiUD+jRGP4E6egKW8AsA5nluDqic
WWmKfpcDmjvfgSuaYfwwi8dEmQ4xiWwNVTiWROtGrugDpM/a6Fmt+XBhw9GWKUp9c97t+OoTZGn6
+uhUS4NyoJtRByZBX6uV4JVNgUfb/IPo+e5Q/DubGDRBp6qxKcA/BmPzZS/0KSeRfHb0qAlyccSo
nS+NdrwGHksB0EzTxS4MHAyd8SiGAXX34ulFEJIcA5YiNjIEDqt3rwNWiLacdCwFAjlqqrRPcmGP
9MS4jzZEcbWLsgenM/5O/vId3LJ1spsCtUzw8eeV4sWSoVT2CDwWBTNkZbeO0EAfDk1Hww5MsajQ
cQzeBv5KUBEYN/c9UL473uMzwTVNB0TNHUuhT3NWjnrAeR5ab4WavZkAVRdUHrd3E7Rcu9hWKsFG
/FeL0XVI6anf8D3OJbCos8dyylXhfD0MHd3SOvV9P3L4qu9+ORfXufIEYK1J57YDVpDJc260kzbD
CHvmW1H1nud5Yl1n30dsxmCqeojLe4dWyh+nUaBNY4+H5vG3IRb10F8hMe979WN8NnfMStsOT/0F
eXHYm2oymvwpPZI1oso1Frm4sGkA/O3zAvi0p4XGDTNpB0w+0z/d3VzXdQoCzjBljmIADBJrrEDo
6JI9JxYq8yKJqxqQ2eYjrdXI7UC0NT7cWOpb+ATuBiSIL8J/vHBmfTTJH0QHN2+P+cPT0oSOTRoB
Xhk75aRkaPCNexPdCnQdH6V6eo/ILXoMhkQX4veyISehh5vE1WRdizRTt51sY75jVqSKpRjFirJp
efHSHmam2AfantQM4ZSXeDT7LjClpSu/GKCwreJN3RLKJxyP44UvhuuabVcL0UEA5nH0Vaedt2gu
8LUR8W1vLbH8HiAbluD6Kp7EsL3Wtkgsyku/fymnpyYCeDzbyF2ionjMJrmbNQlUFgnKRT29Dt6q
eUVea5Hlf+SWiHNcoppArYVspMhic4V+Mxz1DrgKR6mrpqQcP5OT7gINeZ4pdQFdlyHB78JPjnfF
YnpdgpEkVRO536J+P7RIyceM2sWTYgthnv+VRj0ZbjFyum8w852Jwt7j8qgD8Ea7PtvHhUspOR3O
01Nq5IHL3R7Ye9M5/u1mrwu5nO9ogb6Wi4HLH+ueOoN5yoBq/qyAoJcOY5ktUgmGBYxuqRsUUwZN
PvHUwpNEVg2FsqX1RSoVZhS33mtr8S7JV2X7ts4BoZ6aiMvEOhNAgpixTi0gUISK/wJ9YY34QQdt
E+64OTMkKUN/+VV3UD5q+QOImpyEqBycOosEJ51hHaIYZsEzpkyrHzP2aTMUWWYu/QYjJOmYsHb6
85K8YIlh8jivLCOBGvn/J8VQHaF/S8t5HYf5lUtDjKsKsDGdWUVKkkEgU53bxcvpLBplOOJNTRqo
ulgJ8EWR4wM9srkA/out+4e8tTAvWbdb7W9Ypk7TEvpEXD4bnqg/h80f2tpp8grYnKhvZXq0Af4O
zUyXAmIG2ge5XY4oBo/s+/ZkPMtVnIFQbA9d+/LprQI/1O65DR1BwG3wEGekmOd5jQ+DEJIK+fbp
ARFCbyB8SE9Tapd2M8H52O3t7fnWDaD9hmU4n4X5fB6r/RhNu1f+P6Jyn7zoF7GQEEzLD0K8ldhL
c95BnQDBEN2NuQd9ooy68MS+1sp3igYbIYLwFOBVmAXoj1xBj7iiVpyGCZrf7bFi4Ic7LfnXKe+k
wfWmqpHfk+rrdogxfbmDH970WCVfL2JhXGp13BrAcTi2vqBECmSUu0L+nv8mCwdVml5RjT3LrfpD
brHo4nzTMhvy2ZZ51XT7BilhSUZ1mEFPRBP/C174425NfW+buxHBHEfKsAd67ZVA+L8r6uyo3HAg
SssGhjbaGQHwGczCRsfY2AEYgmdKzf8VqYRTgQ7BCimlO1CfXviRujxh0KssedvY2GPPlYXPkzIk
SELQudNCJaOCU81EHbaaMcieBeHDZK9UeXb5Oiel14z7sADHvOLwHzTnMeKOsLGB1V2V2Dlj6ALc
XAOcUooqbY9UPooNuJ+AFFYlQpUFtK1XeKwaXWS/Dn3CScXuDHlHwOqnfGeYljvwr+V1H/XVIn/W
oQCaFIxwMyfDJhimT974LR3AI0dqNhYpr/MivDdUCzffFWi9hjhCurHnvxKA7IM28j82fK4ss/8N
8pGHRfXq0w3JjPmyccyzCNdKdQUQEQ8QpMpBImYCkQhdnBucy8XrRbcNrQynDvsiPnqcXLEETLr4
cigeeHcOlsOCPNJuVaCi0tDArY9qGnZA8pXWXcBaDqAXAzU2hbhsxgu979LmZxW/ea1shpjXfqBK
7H7MDoLejC6EgJrtvQB7N41TfxxwYd5b6hKr21qup8yIoqoWWs0J7x3bOS6XVKL8e0EjsR1aSN2R
qdix9cqEY5/l/c0t0FiCadsGQfc4wCPPQAYeIU1QYUZwbHrZmk+IgOio4Kslp1AB4CJrpMkcniBv
+4CUzy3aWY8UWOuTMh+bhufVE84qTIglfbWp12/u2IT7G+fGdXROnm3uhKou+llPoaiykRJ3Pcld
LS0NZmMQUVeU/wo2hZEaVbwMT/NLlvs11RxNUoYnXX2NldfszWUpiXIAQCrOgZUA+Eqs+ZEQ86dJ
6PeA9CkiPKcXEUezgBIwdvLITtuA6BAl2RD4eP3s2JINPG1uq3uduQDLko/F888nD1qoz4eVKb8D
KAizF9RtvMIXkXF9oLfn77/MAv8jBOl8rB60rcBIfGnUvWdhl5kPRlj3klxFZYtuY45RKWLoZ3qt
d46ifimPe82kKaVaQ9xUUeeRWRDEWSOYO+bvHOFpYAQxIsuHFssHMMSs9bjW/s3QijukHhoMMust
BlhMh/2SI/09pF41o2IdEjiuVwG0cA+A5WmkqDzVuzwDjM9ts4Ykb5Y/7SiRKHiZnxMNIhgSLRPC
PqGcBwr3q/tAUU/HRE7lnGWfdRJK8PjJHvv14Zn+mwhB6SzEcXiwILIFozoUJit45451PwuDNlg/
5/W8tXKXLGGSiPQaQBRwrdCbWOkRDvlRZN3zZJF3pEX6tPQ0dvsqxiD0R28X3KkX1nZvIRbP4cL/
TXGo/DC5wD30EAnRuBW1CfJXA5wBqg/nJLfLOOmrpWUM5yKKNUd2GdVxWiRrU6wErTPcmQB7We9H
7OHFcWYykeJ2f3gkJ/3YquPJ+jIHjCBMfOAkNd2SCv7RaJ1A5+MclOh2LwBGWSz1fhdl7Qbw2X7m
c6QZEZ5CIOGVpDsFaiQXAt+U4hxZIchMp4AaLsOycZ8f/NTrlxwtEFR4bMHyrCq7xCNNtfhY9p1S
tGOPFxvsqBcpXps2pRNvHwMhWKl/d+YMm0OqPnCy+YTlVh3SZGEq9+yYzeoy94JFjAgScK0PIeg0
hdFdHRjYve6SUlqXbgrXYlFqPobXN/sK2aQkCbeY9sEYECfuWogCClp6kTy5Du406bvkHXl9lvXG
hTEDYg/2onjt+n0VkfzgK3O0rM27kPV4G2mpXyLhQlB2NCl2PVbjA2++LiAbn/RMZ0GyGS/BlKzX
GJw4arsxFzeOn5Mnu7/NxVpUKatcoeke9P1xjrmwK+/ZkMvP3jhh2CWOyaul38td2KfM2GYTgIVF
vagl0lBp8jVAOtZqRdZDZPzAo5KPutnp/tptthOZK+rs2CfFmPDF002mBKhj8uRcYi6FpwYEJh2V
jI/Js2CzvMCl20TgvZ+og8C28trVjxSHuPjnTTXK4BYuaUsmjNI2353NeyIog/WFNYUrXTjiQmxA
Tyk3lS2fEDVEIIxgnpmGAHvN4oujs+pPeQj3FRPAs+CwG3NSsdu2PVg9fORLwKKohqQir6q7nbCw
AfbtNJMTxR2T+t01XTyDCOcY0pMaQwgR7mRX2NhDLa13P7We+KFdHG5hTRlvsjO418JC03xi4gYK
IIVeX9p14hLSn8/PPmVgVce8S6QokPmmTFt3qwxlfF9A6svz7/fRF1TWNuR9mTnOkDadsQKwB8Vo
x0gHHDIJNpBkRvlR8v2Qw2ndxFFu39BkknQ4kBFxEocxQA22Fkc7vsgWMVjW5OvoA80hqspqp4Tc
wpbbWpEun+LmYwB36IijA09TewyiwLbWTCdq4M1K+LPejhJq5mi/XdDAG89iaHYrnjcNp6cAgArf
cNrp4jqCBvfCJCh3SY40jVwmA22TgYkrJsX6AjUbjl/FqkJD+1GytyrpkLajFEfXaBfP56nycP+U
2f4zppuAFV3n/nfHWsa7DwowL9HYjM9SjQCyp8L472PZsJ9yQo0AZw031nbgKBwNs43fyrPOl6LZ
8yHSg9JNnxFzkWKr3ZS3t5AtiuXDwv9snXNsLZwVRs4MeG6w400kw76a6u88b6X8/nO8SHfexTuB
moN9zFsjeFi9YrR/Co8I2EURvCwDzgDMgSz+VrYaIcwG8dyVr7o/aDeDmoNCVhWqbG8oqlri8W3R
ToPZCBEVXVAZuhjsZDGmUdmv99b4eJ8GYjJ4/QHE4XDcZ2gs+c0ah4tRdeN/X0EaALsiXj6rHi7W
zFLGbWiTFdW5A1fLaaESGjwT03SXwjJ1O6KXGk1ruJ8bzGQ3VrAgmIekSCZMC8KcwUcX11ci0NoJ
ImC/ZOowDfLIxwWh3xZHMtFaK4TbzD8O3xdgQ0+CxJ21yHCErVid93xkhsdSwepTwRMOivt/UGH+
PbOUtjzk1F5mwDoyZ9J00/XKarVbTqp+WfWv0bfOKCUWqTASG4b4LST/UL24gNt6pe/1sRkFSs2D
7aj3Rn+KBgE0iipQps4Mm0UURaPUqR1ihR8x/QttZK/cXvA0Oh+oy5pyyQuSD/myzfqqaA0stoqg
RDw3UOahcxDmHfoylUmLQirYLy/WsVrHyUGVuEKS4K5tnwKfalFwHMzr3BqHLBfZaX9tqVZF5Fu9
QTspfw/hJ4jXT179FHBbHJdWNeh5krGmfwYK97bmMi8ed5FPaPAJFXYxbQpWS+Gb5ejK7sYzdQml
Cjdn14SOcfmdV1PEyG5pUs8DEfItm99VlEZgVJty0uHOTryCBn8iEc1pQ5n1nX8Spxvd2K/elkNn
jKdrti+dqV6lAZAJMoIbQNOslVTWk8tX489XezB8H9tn2CcttkMIWbRBUMTCS78WRGMTU8div+oU
l/yPe7xAP2K8Mq2veWo59tuTEdEX4OZP8haqsxkBirdzpeXMqljc9PXpK7VAYiuShKOx/TVSjVxk
i73OYokklKCxv5U+CoH/GxrH8mq3dcwCMHFBYghQCHuKQPsygTBOsqc40/lmqKa15AgWwzXM/D36
wB96kUBSi3z8Dyk7uZBAXKV0lCBvNfKvE1HjpQEaaedzZogdoskJDuMXOY06LfzrlXH30EEw5Srp
SpNmaXIgirJZdES0GAAdYDLU793aTWEYRBVUbQo1FLF4Ye8PW5SknFgaHHPOIXkJsic9lZ6rpRmk
wECsG5/5zQ+QB408fscSbz6zEqlZ+51nZQ01fvSoxA8cfaQlJk9dDJ150E3iyS0Wx+4jxjDb4v9J
Zgsi3bYBazK38WArx9pYG7OWPjUXPTn+BB+dOaMYIgqdNUe+ov3tRTgz583i4bYTK0S7xDkQVIMv
dd5waV1REJ+sU/m4TmOtzgi9J0aszDuWpdxe/iRpzQcAU+i63UvcmDUpvVWFqgmPtQSJ2aTbjaaZ
fPo6ulYqkCeev6hPqIqjjE5m6Zyqvwn/6rFU3FK9EhRy2DNNo+LNPBVyRfi4gkV4rkF7sqxUEwrF
42KcRRzVK4k6mtDV+h9Mor6O0ZcUTaUahjlbgLs/vTNcMY6vw8trSti5xiXEcwg6RbpVdf47LkB+
kwOxgLf4pP/ii2uxlSZgl9RHUhVC1f5PwyGVdUga1eIxQzjZgh+XJVlpAMGdhKezaWkkqklBuZBy
gX9ZqrsorXKLGGKsijlIuC2bHwlr9iDOgSV9Ml6myOZ8IQaQYiH3r2zosxuVgbgE1taG5s76Gfjz
8RMdskHwirMK/nCtDWuoEZ9g/X/fjMP9MwyT9gvbFuphCiwUETpaNWOXNh/83eA4wovOBPcX4rlk
0quz4gbkH+lrHTckf+6MFUSJ49Jtxqwng5GpkFDbAEF2711wRT/ZfnXsI16UPmm8v8fz8aQj8+hD
N9Z6ZtvnbY+7Ew4+oULlAsv3xCNhBjdzXKxvc/yTwZKHqpNHJkQBSj+bl0bcmfY5sc0Qy2PYmgyu
7IHx+vgy8rHcNpYzwZ+HBOT2Yrd7Z2ykwqaTW1Y/ZNMHADhEtHHEITMEx8AIu8kNBRX3fbD5+X9i
4wRb+hfsNA4Gq4vAnIl8h/BiWUNXCruX5KIUq/HBomXozo1Ujelwz3DQAozhUB2y5xNjHmKX8KV3
49xEFWL/vohINjHLvqLjWszF7ClW0xHBDU0D+4xyEN7QYXy6ckt0C+xW8ZMVjnvEoES/537npHJ2
0kkaipyfkUN1JXlSE7Knq3+cYqXyFeXioEdAeZqwgEQsutgdMju0wgfLfbBLSjr0EEWXXtgdmpiw
8w1/q6yi1IGHVW86Q5OXgoGl08qTlQ6JY1sFbnw3eDGpgCBI4Gu3daqs9cVgZjV55mCGT/pORuUC
BdvXG9gnKU9FYBe1JAVjL9qJXoak0nYG6N7PNQYPDTjq7BGSX9j/76D/aXOeBX80C3e4nyoi7nod
JyFOwhLerKoNFJ6bsaQn/52FcefpUV7aT3s1iRjBr8/ujzk2MinFbFuqUjlfc2elMTV/Ni7GZGB/
asBEVzkZyed6Vk08Ae7MusoOYMUvK24RK1G2Ql1TW/kdAMjyS7AnNLhR/ZCjbEfcdbfrnbl5efhi
f8VMrR8QRnkVJ/du0zJxRiErxAVLY90AAgek8QFm7S67QvLu/WLNsXWaD9arF7M4DeE5+RTBvdx8
aNUIAlO8epj+lWLQwq7/Oc+CWl/xzC0eiAjtfx0odLkw/zfSSEmg8V8bP4i7A4PWCewkoPpIX8ak
EPJrW3UGMcBDSVM5v1zpoDBy8a98Y8OkMNsHC7qwQ9q6vB3L1ln/gNGKHhuhMEExMWacgdt1XdUT
eHDm1Zzii/c2ZSy5tEGtZeu9Dmb/nVKDtrYI7/3OIxy0sg3QtLcCLnPUBvmQzgg23WTiRbKWjNlq
OjsQ0wVXVLpwrOv4raR25I5ElCHalGd3O4eB/6OvW4vNJPH8sVFuo7LqSrqovJ3iWK1q3XiNCWfr
0H61hlwXftGp0FUHJH1zTpvhEfYe2J2ogfexf/s6qgJwLrJL/0ofgU6Z7QEjvPZ5biV8miQfh2k7
8IGI4nqlbxVBUz78N5qY1JWmw7LSb5UmawfdSISwrVaf+BEHRKZkIXZ4UGEH9XjVJq5BgQms4LvS
LxGYsNqjIgOCoNJEIf0TMVjB9apZ1uiuN+O9mx7Sdl+5SD9qqGwDNmhq1JiFd+CQw9fMFMY8vEGe
ko2Lk+cJPoUpxRXeZ41R8AlS6TE/CHRzgxw8LyD90N4Y+ZEOMiiZh5C3G5RSRYGpyfu4WKF1oT2h
aMkxgky8lhXc/I9rZ8ikucM4H8wDmNuDwyi4UKv0R305A7BJOJkofcD0HKMuMtv5LaOPbSHF8Cn6
VO+l1Vxp8stYdriOAqmw7ZGxUc2PyY9z9g6jKL2yLpzWj9MRAjmKyYMp0zqnR24KhBwydGgCG8aB
mS9cXUyRD2mQ5+2vqB4XEUT4WDXmEp4ynyyvspj5H5OwJ6AuHHvcvIgFSZF2QiX9T9CdIP2hmfaP
jcCXp5nh1x2Kt2TSoOMTImDekl5ENhUthHVwdUtPXmKcSMd2Q/KTyq90lbDVd+tKXyYhY5jAz73a
XcTeoFB1s5Sh5n0bk4oRxom9L7CUI1mVPEsz0ogMslaPrWSftfJ8mYDacS3DUg7IybbMDZoNtMPI
dc5elfewHp3InX9RXFSopOhcXi6iaU/ZjKPVPM4TFSLqvDvW3A8l0z/G9om+BhnoR8fDhv4MtVVl
oforBkFe4cGA5Cm5KuoamWB7452oJljtCBWNm4B6fxMWmEoKyuzJkToDaY+s+FwLQ73KacarcU/I
zt0lzsZJrT07r4wphDvDswZZohOpZO2T1LXDRRpY2mHcRyYQDMscQ+4J88evn+cfXXrYKfGmNMtT
cbc3t6RS9Ql8Jvsr8T5sTv9mZe0KEzrtXswyWTF//nRBrAzslY3vEPNbBCSoUjJeijojpmFI4r+K
C37/FOqKt14VcxbBiNMXm8ziBYfj9Uxx2Xd7nN3GdlWJIoRDT78/rOG7dMsm/ubdzdvcpPr+Wv/b
e3ZwdTvmCkwnMNfPIealX2qxYlNv2dtHUAg8HdTQFOE+0yLySD+FJVPDRCC1Pc9TEWsEXTfMcF6/
sjQEKzooO6k7BMcmsIWgNBKcjJDzgr+R0+XgCcsRo1sHT89hecOt6PXIOp7volChR9a0+6mVLIsI
bLT5A8NU4hda2R7usMRtMDgK9joeoi4H6VYQyFKY8uaBz0g7queZ953X+8qJH8Pmh9AXTr/5UJih
EDMqTOOslv4WtIl6WbiFJRip6zEfsmiCIfatJTUtBwZQe1f/LlhHtUWZBhyIXPf0Rcnvvc/MOAb4
Ew8g8SdDLlKCNwOiwx7n/OpDzHgPDkNbPdtEGzMR2F7ZRMFs1teY92+AACe8/we7ngvodQOu2xZe
IEa9oTFLqtzL14kmExGXvnBLa9wydYo2ad968XkpSS5/Qk8aLGMzn6iF//39tmCVUzKOL/CfjPpT
hTItaxB67nVxI7MG25HJVZFIsB6+LX2PmcV7OzfCJKtZl6quAyMFOl4KgZD3RtId5/nQDndYiiwg
LhJxa5JlmIIuLOmEszFpEkip5nK0OpVhsyoCQvmG6WVUfUAsqdhQ8lQXidowWX7oKruYvLzjE7mQ
UTwZehKv1SjkDsfSy63La+n0mU9c+Ed6Ur3axHHBZHjRDw73dJHsUhHj8SsS8C9VRdbKGvHmK0Pi
IwbG4+dUaJqpTLP/Wyj0qmDcTjJbfWQtoD0BEulAOHG15/x9Pa/alktl6GD7mSORhwFjVRR6nSRf
Nh3lH9bxQI31unsG0s9R/68EJy8OE1xY+S3fXSb1CGb9Z+VaICxDBiJOdfvE1+m6E21/0/mNXvJW
3nbDY6knXYYLLB7tTsu4Hgt+gPxPOXr4LFcmrKYL3Mhpp2UYjx2ZwKc+VvvGy2QilpOdmSp7ok5a
6VtIJSrAbXCPtUSl4mtKEwuXkwemERZNiOfDm+YpzW/PEaj2NpCzpClAc4agN25N6tJ+2F21ygkF
St6kjZpoijNfxSqqsiQ9eMwYc/bXyQizKHpkWvfAHL6DL2gxlqSqFbogkpx3UJpaKI6lkPIW4n7h
slzssAolTZTctSoZn30XC4qq9skZMwQx/pwHeTCzPsvy7qeVfqNuRZ/xkIPtMPTggQiLQFr6aV8s
FqhOQbpVEUJOmWvgGl8JLFKEJBMJVi5gNWWSvlN5gc+YLLhGutTMEnzBi89iirtZN6R8OEakOY6D
UvceP5SendihgbY3lKEPC1dTd5UK/AxypG9RXEJjf4waJi2t6biQaFI8pmACEt3jJPvZxXHXZ8up
GBvj5Xj6hzLB64hjlOJhHke8esLx1Y4K4ouNih+ON0dVnyKM1DzLWOi6ZFzUd1xdx4aBstGA1WV5
BTuVnY4LnzZSPIsT5futnjE/RpxSMyyXGRsgxS4YR+xxSv1INHqxh0lZ5uxWkFASicK9VbMqZjra
/PZuh+JnrFeKJfow3gvc53eY/KShY8GRAZxqpvfu+VMv4E1KTMZAg5wai0cjLsq1GolRRD54r+Lq
6/8oFSeXd8Oj0DL1eOE96X0PJWw0cQ1DYSuvDF+vLE/HhYtDtnb9L+U2bWnPxhJOAY3KEfYXyEFQ
iKyW0gXtq6cSWRLj3AzSaTvl9nSFhTMX4xikt6cIrirsxjrkz5BtJT676trUsPIfGQA452FHPbAj
WC4QKh25xx854y1CZ0r3qacDgHg7SBRKb1YrDFC2aYab3YBfaQNbkKcND1+kcWkG0lNE+W0SAYZq
GCFuSIHhfw5/8vaHJnByNen0aPr3HhQEwxW7/jsMxeqmKmWj25o5A966myEesvJXDm1BmRiR5MXN
7fRk7SXYFldQMDlAGIJ7JXXCeW4+OEmOKp5KkXRoyRmshyi5ajruK68kD06hrf6jF5OYx1sWQTX5
s8yXqXu2B+XWYDDajnKqL2f4YMk/n4DC2+73VKNJ7H/pyIomzWY0hkoizBhCXCfmEbFuEt/754Tr
HAwLv1mhxv8mcuwOdVzSMi37njAcaXqBWWZYu1tTVIH/QAd/8r9Q27nwcE6uyhg+OzjHZ45zSN1v
Tdpa/4zt+xo51uBjgZim178PVuNtkP3GgbJk79MUlXb6Fkhe+3o03ITqe4ApggtupofRSOu5CgMW
F7J51FK7fVy4kqUEryLu4OmaWxbfDYbYnzCg8+p3VGBit/gCpUU8vz3EuIsj8Uz4m5XbVu72BXLN
sVm35z+IypFwSRxJn5ROyngdTv5CsC97LQe7FiuwvjO/WgnBK2ayZmhyOl64bS6omTYD+H8ZX1Y3
KvcNsj73IidqVSLBTj9LODOEqEhfsGpNpfowaTU6pIqZzE/A8OXJDwHdwnvZbeqiPOn8g1Ez3I/1
0s1z6fUn+dsfmLYn0l1aF9xKGfLPAdTXdiT4xHWwOLbM7/bdK26VdM2qfCCMvOjEgAhpJ8Xp30Mp
RqFdsQY9QHhshRmKCRCOHNJxpBWrVBu8LHmO37C/vgpx77q5P7gLlttqBD3Q1A6fl1cTxL/UyltD
hCcYpBz94Upe0TRVnWH7x10TB3m1A8LHEFCKURHTdsHXagiJlKAjAlKBHBfVvsuzrR107V8RXnH4
GLaaLm0llNzOA9z4YA00J7GXhd/wsI9/m9H0+Xwul7BvnWO9WjUzAuhMKhgJKpgHnGerOkqaX2Li
XWhfhXIIEQ+Q2WiZW5G3ceUlLAdYpGV+2GglzmhQo9chmKWu3sea85RT+LDD+UoEFBDChArLtzI+
sEhzIK+klByEveiP0/eWLrfkI7m7rFi34Yfc9GpuMCwDKoPwuGXFj42uwJqlUqtJACN8g+CN9cU9
+OzG9+OMUgR83Ht5oluEU2C8OG/ZRoa3t+PxgRPGqgKF3vix86zigBILWyqhRDY6FXSHZgWJOZm7
5EtCQ3IRdxZqtoJep2JDdBumAkO38ZOCSDI9KTm6vSt/gRJRCocD2BUn1x73o+MagwIuMsdlIVGY
bRrNwcT5U9J918/bVhmbTREd/NB07CXMSyghzvdTUmbSukdfDMPXczh2re59dfaTCdFqd8pJR+Kb
bh4t7LDu6Fb6zet3lcCy3q7uW+x9Nsfvim9teg9OvlNPoosNdEpuxg4d/OUI29DChrbSCvb5wgsz
SEVRjrufxVwdubGxE3SEQaTqotC8ksvJI9KtOmIDQ3VbyA41l5zIGTzKx7RvLnVGls9IqZDDlcaJ
bQQZ8Covefy+oBM02dXqxg2QXpO6cZdxnq2n3U3yyNRrobJgSW8nESTn5QjD5Ta9WwFSVruYiWsL
yeSC8BVbb+V8amxHVa4pUduQypnote2+9MsU12JvF+5KPTcONLSZHavMl0njrL2Va/0dUFpNGxr9
bEk8CxWdbVumL7dyVJi3iuwtYPW101WvpJYPQgXyH4N0F7r+QZ7H0iJsBpS6YG4vQOkDePWPpS8T
40p+1PQFptkLmZXof9/6DGVjSKEEQEVqC1Ww5gj6XUxUN4DimDkZMtLcMD38okTWglaWQV8aRA0h
GYMJ+JFE3ejiBLebEXEuz/LAyP2lsXZMQ80rb9mo9RPsg0yg7fXvogR5jWc1/153iu63ut1glAP8
kjbHUDDeDBmWxsh+LWRJuLe9LtR1C51t4sdyFu4z9RV2iItfJ4fYSwWIGnEN3nb27ZLDdWEOkz8u
EgyPCLCGbFr7O8vz6192AfsQGpeKcS7P2Ac3M/nyWmbZ0TgEUIV9xUQWht6PueB7stfgyOFeLIJA
11jhnI2+obG7KuR04FyVrmkc+byGcTt0FHK33kqXcxToNbPcvfGEA+e9ByWO/i9h52NmqdWV0wZ4
qzjxFwpVXdGnNXmNyhi7CVT5g15dD112F4kWrrM72W4asxxe0H16F/AjMM1TQN/dHvZjg0UwUvG5
3GgsZoYRIl2ZblXl2ZfGem7VE15V9aDY+qElWCcaQBBHRJO9EUNCw0NFxdUChmTZWyquZGv2K8mX
uPEN35iQdLAC4Qon9lF1SJaU/wdEyLp+qBehDTaRQHy23lIRzdrVnPKP7b0UD29xvZ/8/t6rydCl
22UUvtGt+huVUoa8MfTdZQUJJXTRsPmv5G7RHNTJ0++AHF6s4iswdEhzEbAUMneSqlmjZ0vUrmuZ
QLbxiycrGBF3QQC/Px4JzugYiI/9lT9u/DRO8HGFbCUbxlU75rUdeMf/BPQlQareqLLHFoYJeUoW
4BTiiT0qnZtgv+zhi753wDRZbHSVss1fWEqfJ03vj4Ikc8BFElatq2HZmcD+2ZP79PeHLv05K+bb
Fn5lQoGpdMqjS1Q0sllLK/J7/44tpsrqmRZNAlFFFMxV8NjPaBPBfduD8wC2LO2JlneiCWKLRZh8
RJ4SR3RImkqU4OSDDqHJs8DTzYTudF+ryEsAkpVefe6lWdMuA6xHInOyZuyoYoRoO+LbMVUiJwoK
YijNSqhfA6cb4H1QhZY01092YG3yqFshKF6soomToqZBFHWEfLDcRmdu/TB7F2P7nUK8+3aDistV
HmRtppT84/6a99/1De8UFYzg60mRd+8OCZCDBLShMsyDvHstJAbogsXHIPFRw78Cv13ss3PJNauA
ThZMQdQQu+9koDwXI3Tq2gY0eRLrK0hmJwf7G4Fu5OXLlei3L2hJiwNADye9aO1FP0hkvI8DWkcf
0xTU010iMk1QklDwoTLLmzNauwUTkhPMDZ0bhrKQDA1kXqxHAN9UAyr6GfEVhSix0/kBFLA1qxGZ
3ND9pg345VfbQW5yMSPVm240iCb+7Pquq1SkRHRObrnuYnoJ39g84OJ3T31NCwbdEbvkvu/TY7v2
cjIdFUltWUUJyVSiwJgJ4qA/j7+STKTV5jl4iKGT+NOR74kbSc5RxIx2ZNl9W5iK9zFrth3QDqfp
KgsBMuTJKhtKdrDm4PE1soB6n5Q+RCa+SJTXkMD70PyC3BvJya90vKkpfB+Ha8fWQyKMhZ3NzZNo
GdOwnYrvjk9StheshefQ1wXQYZ0TZ8kJsYySKdUlu7HHha8ZKDNaEDrNMiNK9NMqPG+ZSTAIt/d0
InqqNTsgVcLQ9gmiinmj+Qm0U2ys+pNdZqzyv2YPd/SrU4S4PLl5wcaSCTpenJ8LRmkQ/nx8Kv0p
wIjeP9a5fWRPnJB0UKwrKuJ7F5pJwH0B/WwSRuRCMLcv7oXFyPAc2Edbfr4HLxAUL4d629hD90CD
coPxSDLZOlytV9W5BiYfYytS/VoTCS3MgNLQO7gKoxc61B94WKrHBc5ahZOiDN6zDvh93Ms88QZS
BpzNmEU4mlgCVFwULwBks5PFkK00FH/rZQHoLOQUGHX7AMrRY415JjNwx5riKXotmaNUz6MKCQdY
GqyzdAfKKxvLXu1imhWRAntmM1jNezpJfgPzsJm1rbU6KyhMCgS25YGVOkdsoXXP4bsTs0AtbtvM
NQWohnE1bbyG3FFYHWU0K+LecXuQzO2vbeOUsuijvIAmiBR/Nj1HBBQ3AAx9nub0507k0hMIOtrS
F/Xsn5gR/cHFd18/siq4/x7x7PtyGEwD2dgSkLJpXbLodd5fknmyT9o6uv94uxhpkFST+srEaHFz
e2u8LTACti4+JhA/6NUObYQt+7PEQPcz0vW5J0pdTspbtvGnkvJAixB8lxMKeKRseuspeq/Bdf8r
WMfcfmFqUS2dtUkDTSZIp340mzA7GnjdXT90gQffe7fHsxwxWZGlHXVCbh8MYaSwWwds+leSDGGf
cyMGeOeMjcDf134agcaEMco/fB/9IxS94wZwSFOnd3Zaac5/qXCEaNt1Ql3uzyMwvTaFSMEDFFXP
oRhA4NVSD+QQKltSel8pZ7nrznpb+vg/xW8r7Thoo4tzFM5A0YuoJ6AEeCEThGYg2s339OLCxka7
66YcBm2A/H2t1oU87sKNCAx/l7U0Hx6CIIgvUcM7n/gdd1E/v6NcejoKXeqibPQnVrwAjeymSeEQ
Ecl3l0Qh0ipIwQS36rxvjnWAb/EinAQ1PWakg29cnewUUcl5xFRVQEMATsXm+OXEAzXGqLxvVGoP
i8jtzaydnfVhYY0JRYy0extmMvmxlBYeSA5TPR1903xHYmoidjm8wMf/mpKYT9INmCjmzC6rMse7
qxAfYu+/m886nXVyVCSkt2l0Nh0nPry/XHI/2E8gGf+O2l+0BcCv9cLDXQ+jjypptyWNXxSqYpqM
/C7Xlsuadn+rbyR2cu+CzOCMWlIaDnmsxSC6P9A0NVMmYOOFhrMSODv5HefWWElopuHPnz3eUdv2
998J77DYaZZ/2Sd0SrHShXmmA0vXAlKgfLerQhJsSff8kAucahFSUrs2sa9yLMrxJFl5/wnATHL9
BqorWJyCF9tNmBTffxfh/K03wCEUKnZOMUm3/LbssgoOkALugmxWPPImIQI9x5K+liwjb86+GYaY
8CDJ5Vb+8X4YjK2p77+/oiZIC0BL7LCBKbEl5UTo59krgcQGrNa/YKMD3fIInQlK1IMIb/yO5fG9
Ad2mi4ZK67tdl48mxDg8Pl0fhkibbSt/4RhGQpjy23HhUVTD3pEuFQ2Wxhp85v0DeKuVMIK/jFN9
tof4mo+zthmPiRPp7Srrtn/yFR4ZYHW3T+iQK4qfoLZn6Ph8xk03oYQ3MLf2vqTmEg3eqGGgSC6+
EErnkgvq0db6tzHh31iFHw4Odg5jL4aa8Ux0y/bap3hN35SB3ElVo3TLZPsU+gGImMfjDDOlcpwx
zDDfqPxbzebw+BRGLzwblnDFK7rexku4OKz8Z8h/qOwfP4Lwe8ecwkIsEwSy9mDn3t4dY3wCyTVX
HKDVU/obfrnHNtJlZ/0jIVIs4NGRTjs8Wy8Sc/8iUonDRDvE2MNYUvpPn1QJMPy1DgrkDwC/kS+Z
mz4t+przu++krHLC6NGrH0r1dm++BVkga3IuHdkeecAVIkyVI4EE+tSAd+l5q5Yf0WcsWWJMvexq
ExhSmwj+MTtIvk7gckj8Zv1ZiQ5F3kItqnX3Sr7I1wo4xw2bjYDrRzK2491fJ7jegUpJNy68f4pZ
0ruSuue4C6I44a+h9poIl2AokpEHiK42Q87LqvRfxfOrRx5BsgcqnhTnN2ovqP1C7F+FuPW+QCH+
6LVvcBvKaB0O8cZ82S8oQltwRZPTI9JfAn0M3/e+kk/714+ZWBmdQYsSNm90MTzRvzdDWGcTwsY0
+tT+Uqyi8abtwfKa4Uhjhmish6cUZkwRAv33st9n7AC22/mpjgMvx5eDeQ5HFBhUSDgcJPEZt4U3
/bgON8vecgzZSu94wDcRmOawkOJXurWxgCSEBDILB1ZEAfDETgZbgch2XxaLeFzXJftznbPaQUNK
miThOthlCkXdb+5y7zXOOgsWgyVnr9GRpG8OoesZVOuFkR+NNFvOfTbwdqCWTrAMHFA4GOE/lT9K
D4GXml/nKTE1V2dQ14xb76d0EsmQLuI+65XGHg8pZejwGOO/0NGZVSq2zNmz3W5nj/cF7nvHf93r
dUDmQm3Gd970DQBFJ0q/iqglfXfjhScqgVk5cbJvlds1lIit9W/JcivqjVp2YLe8llESaEE1X7JE
AJyZkoXVin8yx3SO5Ng33x0ORhvGm1RaBCb4wo6zML0xWX4Ns+AajoRYC6d/o4SSNsMi3u3a4BzC
ZB6yGcHRC+NueetGzL5MQXK/Tr2ZWkj1bS6/2guY9hhY6nXWUdseBhjWGW8dIFctH1x8VJSkngS9
Pw/J9coyiIQCLW5vB3fgtuSNRVTUl/d70SrGneJOkUbut7rcRBF6TtT0hN9LJOTSKwFBor4CM0i0
Xy99nM9R50KeQyPw3QK56iL8Im6em0qCwY09kIPb/MZY7Q+tVHhCem3B+lN3h7rqIVIRWk0zNgcK
tkpnjPXBUnpB5M0CJuDBDoJGstA0eqLvnTGERWAiQZlALdhbQr1g8zLSFgpAKVLNWD8zmGpC4Ssw
yqJx6v31hlunxHnHU4NFHB92L4EGktHD1UdSd5kVh0inY3+HUYZRMJ72AFo3sLPtABTze8HpnLQK
Zoo8hmNFeYQdDES8W9VFgzh5DhesxQdVKPpmFeM8BLyJgoqkMxm4hSlOa6D9CjG9qS9MXGFqGfRW
Wv+EJFm6BpkXgxIric8gNIIH3Q8etQ1II6cVwCkW8amee2eqT0qmqvxUs8fIRwNGkH/x/y0yK0KQ
SGSjGjC2lxNoIFCTdCgod40o1L8wDRAxY2yG+O17vrMg13FQ94ZMfmwH4cbbLfn3mn49BMoL24yq
DI4ZUMC2X+30TANTOEbfh2Bise6dHyVU0e+HsEYjafvN4TSlUTLLWebvoiN94oYCsgodtA+heIXL
lace1rpSVgqQehioQNqiJw1AkexFFctLGv8o4rOtnuiz9ywwaPuQxpmR0yGzRoU8arL0NO0Nzwht
iLKpGdO8CPawZtzcsnt2h1AFZg0q0IrVdGnHgYVZyvM0SED2jdalkypaDsTPWucya+ZgjNKs42m6
C7Fv9gEVhMpUIpBI6JFnC9Cj5ZmSjpDKqwkR+IaugBQONvbz0a1zmqjY2Ag63IkdKbc+MXqDMfAA
e+9sMdSjv2IM85WJELihij4ld+kipD7wLlMn5r3AUU11AZYqtuLPNv6yL3lKp3ZmaAmCipdYphxP
Yi5+IQpoVeJsFVcYTwV/jxZ/QsNLuqO8LnGzKG+y0+Obr0qYVBr+DBuSVGJbIM4X36dsC6A7WicW
8eXgtsxo8EauCgN+qqGtBzSE61JNhnc9yAZ3ElBZ8C/XdA7kjlJpVyCet1arS4MOeoIA/oKCCDVn
W6OInsnBqXH6cJvB+L3cLMUgeE/0ibQr1M6KBlhsXXgbeeRyXpCo7v7U2PM4eHib+1D6+crIUb2S
x0jv9xNfvHqGTRvOw3/01YHK25c0Q7f7pijn7zWCt5AF/HF8k/0ZMzqQ3nXveJLZV/QSbk+TU3IR
z9/5W2LyjlhHODkcdzrxUaIT/fQEOVKypWVrLgOW8XUuJDYjU/84SVBeK1oeXqWKKssWuK+bGsVd
GjbQm1Rt+mDuo5FrYqexSHhZ+Oog122+7NYekpQ8ucaRS/1zgl5HPfVqG2YILKVFFdOCbP7Jr+NG
k1qKfiYQsJspwiuB317rs3bjDS2q729CKQp/nqSmDReyFxA2jXiNqEMTbb4SzDM6q1mRaS6Uhno8
5aGcxa6NoII7+5vmEXs5asYWFd/Hmyj2NEsB/RSMCUy3hT41daHLq9O5Hh7AZr4UijpW/avqjJQy
mfJUuzza1spjqf4OAwOopDS7FR6PoOBCZD+7yshqQv0YKRG63BJ9Do/981V6BPbxycXmjY2zLPvS
008JORTSe0Mb5L5CY1N8lFtCPkuxyT1oFRyTJB0maGg/OgwJStOAkjpNZz6WQWPR9fotyZ89A1aq
3+rEjSIczrfIMkKLqu62sX6qr+ERHlsrhtoRftd6ybMWHyreWXuYsk75ucL/PrrcXbqOXbUxTLCn
wDo3ZI2HusKAgNEXORkhD9voPzUcrXcKshgUxY9CfhYbYUHj3docmg26IvebXi9suyb5Y/9SV7IP
ucjfbNDsNAqMtGGRKebsUzjrssxM3N1wSvwmNQLTan/IfeZkLaxbcW6Pssfk/Nt/FJGrhB7bQVsY
8Dc/ltpDhJgODKf51oezjDCBNOzXTHnoGXMYV09OrJbp9nele/zuXd45ndngYTypoFf3863rOSYs
Jk5sTxbLMODthAzpEZnGtSHYE1Sg/3MaokTgxByHavrg6GQV/gwL2hCOKw3KR3N2cZJ2PWkklF96
PSjfspckoIFSxucAZygntHvc9LEuQdqnNcABuvh6jFrW4/rF2aYWiiQ6Wl9E9x/tApKb368EfRxz
VZe+q00lEMgkSjnsc3IxZU3610ztYGNeI7X041ANxJeJYOiV6v19TXLn2sZtkSOE1GxkvxaI7cj2
WqzY9DZzXQbjC4Q4b2P1aQdC9BRzAFK7imLhN4uDl4cdDGa1EDBHIhSkY0iD4aLAK0IeMuxzM1YW
sUuyLXBbci/5ZDlG9jmD2LDja4OL1xkSKkWVsFLJUBEjrBSbt9RgPrltPKLQUx5fO0QLKZ9OLl5H
QcNAkeC5J211u8iMWXlCt6HdxoGvR2D6DWJy6PRnaHbVfSqs7F3I29n/jr8r2grDxY8jxV0nD3AZ
zTN6sTKOP+NOnnaX1zX7N+2B964qKJErO7HdSbS1WAAG2HW6Recji0vUIl8HwA73R28qpoPZ06Cp
C4Hw/J2N6T8vuA/RP09YhWpbgDnTdErkzRea0auOZ3IVFvZgTv0lDJberUTPpa+lYsVrbQGmuLD3
ONQLa1MA9qbLq2hBSLZsDrbfyF35jSDZPa8i3fIenPxCbr/SXzl0mpEx6YS5a6YC7r4e26xf7rm7
izvyLEoQbeN4UQll5UACslDWuO/U5Ylx//qBMSqJzY29B9QuBP58VQr9je35XgXhXqeJh9U2bJSx
GKeC5swntu+tBb3IdH/4pPg16gt88cMRZs41p+z20XW/D/kxsEPdVmTws7tL2UEs1bzCyVm89rzN
YDd1Pt2Vd8eXIv9oPv6Ky/J4nps+siLbGBsqR6mNpSkyrLxR6CfBUxhRHOPTrK30DZfkZ6Yykkwr
SPKM0WLphNvFpMMh4O3n/hmLBP5hZfgdy3qui0aPZ4fny5Fs37rlT1jH76LPYCBxkwWAcB+orSgV
tBOxAyZZ/Fxjj35pNxO42yB06+e6/xaHJIE4+7sNA0CZ9GuEp1sWiSn6b6z9RNXn7OSi+qxjc3TT
sWiKiRB9/N57cSUoNyfEQrJ59yXtTxD0cXfq8qqvLuYHxcEA+NIck1XE7rzisyfE282gOlyG8eRn
78u6b8lbNdwGM2kIoYqJ48YELNyD06iler3b3QRgNKEDFdu7DScz/8t4quN6Ifa5DGsmPCUj7OY5
YpX1m2Oe32abqjyBn4uD920gmxWmEAcYZUWlMC7luDgC91KVPuGz9yhPEesm3bxt/69hh3L/zviI
wPa4DZFHC6WBqITvoCun/doWLX9jft003Ryp9vqnaANnnboK/vyE6mx0OVXRKxgQ/N1pbtsQdown
brxkAiRI4EpQQ61YfDoCW/2lkjZk+AWrs3p8VB2Wvse1GJ1+eochQmcKf4MPXZWBeuRwq6AGtU/8
Ie6LMZG3C6gSrwW9qcbrfK64YX+hU+fttpkrVdwg609zd+SrEFAwoQ/maWOQ0jHFOOylwn4QIqW9
GZ5C2MiWPRLlkYizKP5mJ/kg4k9E7Isgp3gLKS0LkSZwunUr8KRlSrZApk575jMIkmzz9+v2Pfsy
/zUFIj4alTrWn+ibzeYYQbwqt30ED5q24TtI8kCvTDtWb6HxOiBKzubVNBIfZIAWrp37ddZKcv4h
5510E7osoK2nGbbkMC9zs9sM9pnjand7poNR4VaobVRiJNW2UX70clgTuMg9RJxkeoDPrbrb76FR
WhXl/Gwvnc0nRWAsFF/OGf3qJGbJOZ38CXyhXfvzCaqy9qu6RQ9RI8K7Ki1UXE3Wct/rwAujrYvi
9Y5PiC1U64+rWsRrIObBtvIn4R/yymzOjstiAg09BlLzq7ZpthX2dCVFafKTXbBgj+7pPpqYUt+n
R9rEpMtqCiN878bIIHjHr2vkROPZewltIeUnHOWDVKytvLTVUp7nxfghpTt0WzEzqxDgVw3ZOIjk
E4hOu+Gcvct/DRvamJ/jqH3rJa45dITUgXhNpwvN5KPjBstLEe8Zke5hiNqGRBqcg8XfVeSsq4za
1TfJiqs+W8BRh77ANu1NJc1/bWVURNORJGHVPvp+lBjrGaGqLADHgUHIKOE4RbNXMFbUOuOJ5yb0
enhJerZXVTdoRmjwzFug/uIOFAkt1Y/JW776CJSckBfpiL/sx79m78fPO1eD284wkQhqnAOlPSHl
zmYGYtQlPhHxFw5Hipy4L4aW6MeJbETzPK42BAA1XZxJgr1a6X5DaIKaafbgS944UrxN1r+3brVB
oqtcbReh8vpr+jKX+daxgwOWW/PYP780l+r1w3AAcu61scEqmqbl8FEj6ntAVbCIDWQXeE79V/G8
SZseSey0JhH5qaBko//1XHkbKPyOBzRUXJQrIl+Bt+dDKBt4kbC8EDlyxfl4kPkdbUNYEj+FEY2e
Ehe0YKN4rD+fzn+uKWlaqkLGxhzbU2n4iIqDVwRlAWX4I0MkH6UIr7H0pXahbon9mB8tF5ezmfAS
Zjz57J0q8itEXaUR7fpUCcRZ1odeIQNkl7MechGrus9ek+dv/fDe7q5YWu+ysZLtLuJijRNYYRw1
SMhNtorxz2PNk4FWvMsoXAmzXkGlqG2h3C3s5vctmFc2rRJj4h1QjJhSgOaPc4FUHFq6Vs4vuFJ7
1Bbw/mYu2qtN+PlJUJSh5sT2Mi8OQ9cITuYJUTVN4mniGLDHE7zhWDcVfyznykubeNiEJ0d8p7tG
xd6po+k6PpMgofwGI5YaLvz75X42n3zHxsUMbS3uZUAvT3mdSo/8beut8zmwvlPNAnfDDnTVXH4/
1vlqHrPs38d+qEgFDeKuItqMI0yxcvIKAziawasFXLCwWzEBjeYcAzuPQgjyuBvj+vxlm3fPDuM9
ZIKskAOJWbOlCRhOKwGYe6HBDdv1+byExCA3edgcAgPKba1b0hY1UwUIKIrz1pDv+CV+M+PjJlFo
XMDCKCIXTWC2lr9hR2/9BNF6Kou9ug70g9uUsZ8Eid1KAjYh65tAvDjS4vLcK8qufM85Qb/TvmlK
fYLygu4NlXJa0m0GwxikH0p6AWqvklrb3u8hMWm/w9a2SFADQTgFaIi+X0wgrCZMlIwAwh08bev3
AV+GrA95V1t8j2DTkpJX0AittaU97Gb9s6/gYbviUtTSl/OXJAT0guZv1NnPSZwS4BvxeftuOwLR
sQjmNsKWTd2DXf8ibnBKRVtBW92RejsdZ4BVfCBvhA6h3B7kW/ZkKHsONkdHuhjsPGeLayGmLzAD
Ku8TvbxnrMYLEEVlzTOphcWTGyTQMTvS5fmVmdehDiIn+xZ2tM00YnAKYB3JjqdXbNSJKJl69yc5
dni3EjFzRmlz1Sap23bbKjrPOWFchdNNdedzh8pOkVGTIEcs/Hy05gsoMix4B8HACPuioHvYicmu
e+Ugz5KfYx5S+lKLtBYY8vgeYWMla63V3kYUMEi1cPCxFDvgiyI3zLBaUZ8dfY+MJ5T/XnjyH+fZ
JseaRCevby9Fi4A5ghaffzBOvtnbULG2AJYIevRQOPC6a6ePlAHTvZBSYtWKnDunZstN8mVOe1EE
ZdLiUVICFI+zYNwjsCZOnDXFeE4EkhCa4dShR4QIplyWeJb6mCZ0f+EqKJp6e4d34mfJv5sk4eAt
7+aFJOQleUTujbJZV0enKHYlIToMsy1SZfDJyHpa1bRUi8MdfjBDT+sRDDdEWGnB0glf6EmcnVu/
n8j8mKvqoyBHFe1RkNqZO6JOGmsbDNfwI19UuL9UDMG12LzGeqFtmnmb2VXLUVGfJSidyg4WInPS
KO8WRnKQMCPyBCZ3lk5eVaw47v0fMKFKNX/0+HtvucLm3WplY/nRDENl67xthuErHpGTsxZRhm6X
veYPTxf4qVW7uKTx5GkpbCoALvxyVkiuUxwcUWAkysidVNMDP7+JCbXj+H14YA++dHgFSj/sz5pN
AejdyxkGGHc52JUzUJ5wo8f8NeTz8R+fKQsKBqXSG8dCNS/R0RRRMHnC0yJd5kXzz4fXMck8ZsmS
1F9HFNCcxe6i5kchTswgUZ55fgeZlS9Y/pb4XJe0Q1ViixypZNLD+GDkQPN5w8vNFZypywBAQKoU
UJKCc1+qwiEhMaeXSOowEq54IaLGCOlIZA7agh1TC2YtuGo+P9CMmqFaLDYHBfO4jFSJSnpaNemx
BuuSykr/20Osd1Ydqpg2m/c5hBrl6l+NYwbf+seleT/pSwXth3tFdungt30lt40Wde3izGAPXkMh
0ubcMLPXBIDqDV3epEDKWMX3cuGgMzFhchcGqTXvxrhjL3P0IdcqvyQSkfW4O7yjiG136GHaFEpK
e2EZdT3IcU6Gm4ZKQv38YoUCYYGOO8NYl3A/iXicGZ5bxcRJOqrzjdwS+Ysh0pVD0Kr09J8a3hU5
KSSuMVjc1/tTmV7Sr9eGwwf2yJA5nKJTiFReMi3BgXaxLXqIYnVjduJEGuMdY7FSVNBsfPovHTwA
6AKmzo80Q7zEet95bor4hsDfsRD5Ooh3tGtn4/6yER86yPtbfSFsDcG0eh3vvnAk9izYn6LP374Q
9/8D9RNnWuFsI760G4r9aIuswLrrij4s+N0eqWu5u9OcCuU9L1af5GmxJuVrKi3PAo3idZJFJGla
i5O5st+PJ9Nlif3uiv3aZgU/jrV5cj1JXdMcymJIQeUoYcqCdEOFzNN1DTnxgVKVnNj3aO4N5G4q
wK7bxKvz106QL4q/pGVvIYnlAv2gnL0KPHwSOaaZYbRyR/ilAxvADa9RYmJtJ5rwcIUN69r0c6+n
Dbaj0IKuG/hoTjDqLvFpW2+cfP4G8eSdQtg6rAvIuXhLObBlSOeeLaHkk3saG1h9/kJWMXifgijb
olWdaHRf6Npa0QK8atEzLA1+bPjjl5TQz6LtAHTnz5a+YryNjiH5eXt9VHdpp+YYmpy/iCdWzBxS
9/eGSBX1D9TBLMa29YiekPXD+ZamQoAu85qeKAcuE6zMZzDSrzY58I+FC2hicOYl+Gonz6FQ4WA/
Cgy1Vc41nWF0c1pUuZ3NCnadE9YerWUHwtdL3w07vMQZqjhJZ9NOSwZZSx7FbyxuTIGOr7/wR/pa
e6FhfUCG/JDKUZP8NYcomKdxE8sqGGe7erEEL3FedoOcB6ayWycWcDIozKfrg1/rx1VDsvjd4wtW
W3AuToKPi6tU92/dYbZcWXANLHvrHNh/+tdhyZOeMLDwh7GbXbos2Wa5WOXuVoJOfVlETXplOLWg
5O429XqE/sNQuy3Vj9B1tZmk4m4x3nnQjBRVCZU66LenMfRToyncwPlTANFTrxH/peAuakN1o3qh
yKMsttZqAAlXe2l7jHP9bx+MCaHuzYGyBCJGGmx6jSPjERM01jg0hS5Y/lI9QEaVD2RW4g4oO60p
O3WINwnN4mvMvgJ3cTQmH7b7tHZ4nmd887ZJtC4a09n989DvMY5NQVAOG3X5DEuXo5MG3uuhORAy
mF7zQf/SjiIPT9Day3+SYg4a8NCSmXl0YoEC1D1/iyWfvtF1F+zSXkrZFxjPlinm+p4N5fEQcBW9
3smRu/fhlRfnmp3OQ5tgcKcQoRdSJ7IsWHFSDu+1qDEoAoit5VC141436OoBOk1YYZBVU6PXwNC2
s8eBTzae/yevRlOqsbuL1hWew8vfXQ6C7bAvRpEBl+YQMSJWVHoxsHt90cbxHWY6Wo0xT2P79o7Q
QlhgZIY5fnAbwiicdICNeUfwFs91lj4j0JQ0T1bXRNaC/Zt6rmq56MGqwz0WlQ4riLMg3PuuqOEW
dP+HsSJrhN38yhToE7qP6Bwd38RerLHkZ71Ud6+iHBj8V/BcQ9sGqpOl8TGDk8f97yx3nU8w2aDH
iJ1TVtNcyvYhYqY9+tTJbE/XhfeamjB0wp7EjtSTLMHv5zHLUOwQhnRlKq+grx8FH5i0qNZBaML7
2T2fTYSRdMzI/xwtKEeMki84JiqNaSsLS4iL+wLotEIiOlpLahr6lcppOUt8S69LJRXPzUDghtCi
2Q9dB9jrGi8wlqO2wC5lf4H0bWxRxpGJtPkGg8WF02dPm4kq/VLcrQmcyYz6q8gKFBHpLB/K5aZj
jWGQM6rwSPtHFu1qnGr5NlDYYDD8BqNp1VFwayTVpfEjrx+0I8d48Bgkxc2pCmE5GsUqFDjNBDY0
3tMi3mPZ5dunDig86jz2D+MewVddE0xAaPB4OU2SPaRDmwtsVLS0hcWsCf7kie9Z45hA/qjNAvTb
SRwr6U31tRVAMJfgjrx8NSBO+wVzEFT+Zlfsfu1Lc81b3sHMbDTgIXRI/sres7eUJXyIuW6o2DE6
mSUKTsA3Ud8zatKKY8Jx5Uo3yOAZdzCj5bWI8LJxs1v/FJ2uj8SORw/GZHY7flaKBk5fSUi6WOAP
u5DMED8qGeM7OlavvZR+3xdm7eA0sMDIs8cWRpjXICg3Rt4SM4PYVeWvXb/hxIeLY/50g/2Bnttk
sKAxg3I4u9SEiSxzQApRXplqUXpMKG+AdCYYOR24/l2JZuihyX7K15Z0K/iH/PJaF4nTtmN7H/ll
QFmzl6agYFG0C04q1BiMHLui1gqwe3X05xTQ6PIbVzEQKiedOatULx+ek+udpG+xGNXg3DM6JcpO
46/0G1afHv9ATm2b0SzUAL6gSeGVaoZBVk1L2v+lcK+AxvrpLBlAyvI9hj1AZpxOu92EAOo2jGCC
Ih2JV4jqgEmtmPChwIaXYCWUW1GiVcb66OOesGxoOsJ6l8tu3i7q5Sv9naUbROhHqkK78zczgIpJ
qnE05VMzlwY4jWx0TTnJ/mT+QgzXarTXs0tCkETVNvtqSN0S5bVJG9ZTeuUrTYmVLgjSm8gvUQHP
KiHEbnhdhzNuJ6Blre/3ueoLUpyp3R7P1ZoQ32fD+KoGtOmpxy9XWCT5ycCVj1RJ99X2x11oz1Xu
cSx6SHRWa/0YqGxGlKXG/2PF9yHuAj+z0V2lLLcsbK0kpcblzj335Oaejkev3JS4zi8ntviIsZQg
JRUenLpdqQNh3btkJLREen/noxvpjo9ZgWj8yHqyCSk2Iu6nmq0eXAUPWtgJDCEijHipi0Zv8UuU
iL52gB0sMKmdK132EbkKcZjW4fFQ24Fb88i2BaoEESJYjT0HxiyOdeZvxRIsNpuRheqqZV5M0+Vj
cud20kuxukjQEOv52YCVLwA8oaqtS2pOOusV+8YzCCkIq+dqrDO+e83055BL6Gqi4moODeZ08u01
HSAxH+QYjhqX2vn7y2fX6RbdVKSKIVE4uRk/+HRkG22TG2v+BiNTRafP6bek90vqXzZSnm/+nolL
0U8iyW9pGddMBnrvVA6ALa4xG4XBEODeXivMUifpYIcXEWJgUZ5Iq0q3EQHslx3M9a7EhWrBhMkS
D1SjXLa4FXyzmeSygxVya92sWQUK0DF2E8b1IbUqGYP8KKQsjIiWPiEZd5UuZ9ENLl//qyemYLMt
nfBCoXu34IkaHFXLRn/D23uURN1amKAzdi77lI/QSUZJr6xmMeC8UxBxorDlL/PKVH87W4QNwUs0
ala+CJVA3UU6YfIX0r5RfGVIbufSU6LJdeHQB7MVDE/vlJXsRULu3vcz33yeo7spJCdcpFmD5DSS
IodyPLIjWGlPkfK1kC/kB7lPhiAXtgOpU5uKYyMqCIYJxXu+xBA7N6sfjHh3tLjzY7uay1muFJuY
y4OqHFfnc1y9jwSm9/HJu2eIGW0J9S3CAi393PIxHglArq15wXqdA6GGMmFpmq30XpsKldShEMYD
EYf/VjWZXloppWrEAzLghquTlTZ2qX24kGZmpYjSxUFo/94ILH0WDQN1jIvos1zEV9Rgp+pL2piS
2zww/LwcNID9osNG2SNRHC0edBTlysNBiVux5ho9b8Bp4XGgwe63ZzZCzBqcrJpdNEC3nya1d2kf
BOPWSZhd/VZdxHgUdlznuTVxUceAzYMwFm/jgCck1/NK0NVwCTGnu3QnhwtoUIUHVoBj9XXvn6iJ
a0YGUYX1nAl0R+oujUjF3yx9CAEiKRLdRULcBu6skCb9/7KWWJ8AZoZAQ0Lv+gDJmxyG72uI/qzW
yNqMJ75k2egQVoxqRVP3fVVVWqpPDFed/qDwts/EbNvlQFUsXUTMpBhQ8yZouDcBv26+6QEDMHBg
L054QfJRESxybY4nEEswWwU7IV/SK6daCcYQ0YHW1uX7OoFfqHJMdkGssMrknrEmoWy/41jcYGjz
BAbfdQoYP3y4FsyI6+LJhqnYng3rXrE2ghvlqGidahNoo914Y4/YQxzVU+jiyX76bZ3ThhY9ZAci
35cUyLrfLs+uu4P7fV6eLYTHjDXC5yqTen7EcgmrYepTpQBJVlilCvc3rBnRx+cleJS0ohoZ89DT
meBIS6MbTOvGRniLrTnz36WpD2Ar46pjxcnwWFhPEk/3NM1Voo79eZcgDapz+5632ZHTW/aO0zxR
5xyudhR9uI1hnM6JNYK5+znV1Zm0r/zyxRJCiLTQCRN2JldfW+oPI7VHD+6ljh52W0wAobZtaOy/
JLkFnIBK9il9YZvc+Xu/NMjc/i+TyAmPC6VwboQdG7REv6mDG7EWHhrMiMYwgULAl6wwoZxEx7JP
wu4sx+yJhBa8wTMzBX56hRMfjPXgYY5lJw1cPddVxh1WMR4/0NrxeVJnuwHeKPWDEwvWGS395wQ/
vwytviwf0zBA6+9JeNgmBbshV8OS/o4Mj/RYSFG1QUFqFGcnaYYYhB1Yf3iUiLmFnxxiwKZCIphZ
ADg+nB086yQvsFppxyVP1RDzHxK6i+lDT/ox06aY5+OvI+r1XZH8ze6+GBtDUU9Oj8oN0+0bBPbf
Z+K6MuxLwqXkPFuhh6sY0l+U5y2J+IAgE2dZ9S2L8jeCK93SY0JbYJhxoX41JjEACnltfAfU0uS3
5QEouZfKf414O8zZfqMaZZ0xUJoLeHehTEM1M1G6sC2aZJpu2nsQx04LEoMYO1HOrRowvDuc1QX/
LWcRTp7auvqtimyr1qY7A/hI4oEhlTsuxCbUOW+bv5xS5d29iYsDvJsu3sOaGfhzHXovlvUK1bqO
mzzRipXmzxmxGAlb2gCiSu/nKSd3QvpCGoydfT7UqkLmRwbwvXAh5NHVO5UrBbHjz6Ehrd7mkiU8
aM6Rb//AI+a+9LoHURN0SFM7Au8+mUSyBdWTrZZOrSHXFq3Lybupz+O2OFrkh1DwFmqopoByE32M
5we/hP2dQPj/8RA0xbRIDhXLDgjImQ2RnFjQO8+tnQ16Xu2Dk41FMe5frqiSUZJ2I34iyneo1e0n
i+F7fIBRKAEa3feXAhrkkheXGrT1CKZsWHkm30TevUkT+v/88q+Oy1P5z7lzX8iOYbJcZakeDe+d
LAM85WMThX5G3B7v2VD6LtRovx7V/3e9XF48UUSajkVfnHgz/ztIXDONMGU8pZCARSgfw7IHTpmq
L3zLVfBBQ7wGEjAoDVAff0YOHPYkOqOnHX4CCuj7Qp+NTxuP13PXWG9KwqhmlvAfuOMzyhTaRs6J
cjpRHm0wWwt+HWYFOSkWRQ+i1PM9dKsKJcn3moOXa7XpCmsDH7AHIAXm+ihfnRdz8Q8oRqL6Mh5n
RJQ3m2rNzw5CLTxmK1HG7GgB87La234LaZe06VTGjsPrx/EWGy0otKIDzq5Mj/McEy0AHHh0z2nm
ri5O4ILvOfNgkOtyXSY2NSSrY8rov6IjDIexmjQoAL9iH9a2Ca6ueQbXOBv24VHvt1373Y6lnUfy
VzOCiB0KJirP4PIc3gOkO+C9ftT/Kpb3uDrn31hN4CV4LZs8ypRCS4k3JDaHo7ACfg8h4WyJZqIO
q3IupVhqAuuzIMuBxO6YekZczuBAdfDUnB2t05Yk1dtudTT6e4jLgBwcsr/iehXhT0HFhRJUsWRi
pfb4yTcaHNwBHS88j+zKcLAxv5+A+D/IDW/n4Kn5pdsC0M3J7sTQn7m2S+07QIFQgOPZkN79mYlu
ECEfUURDDSICzye7JM9AmEq77eKikRB/h2Ri5cLb99wGrH9MtaQLhEcbGFRxwOFg84p1oT4lzOLf
7WVy2eHrZ0SgmzhQn40ABf6/JvaXLZg8H4hIdPQc5/5V1QHMP2izFEPlYjoT89jif7aDr6dd3aVt
lPhPS+A63+1EI9KkrS5tu8lbtblfazYIODR+c98BQ4i9YqcC792ZWB+EuMBUoZZx29glgyGRWVRz
UW4nRzq/29OW1TWmuYGg1xy9kZeF2w9acCkJwSz4wWDV8bR2vOhaye0eh4IPYfZC6gEcU1UFy23F
UQPyUaJCYsu9PoKu57bePRVDAsR4QQNmTrra46aj+4fbilgeTpfPAL4pXi/kFrn5U27wJ+f01M28
HxAD9dsYNX5Amw3ctntCfaimLXP3QPBCpG8VgLNM0cFGZ6RuNZcUaTKpJdexncKfWElSv59Af+VW
e98nxY3Wh6B95TWQKnUo+Bo1HcAzc1s87iXls5or3trO5mZHhh+NmV+LC232harMILcch3TFVH57
QXLT1gTRM0P9hx9FligLkBA/BnkwyL1b14wuULyHVxHMVcAPDmq8dnwDY7lSkeOfVUzyV1rHofYW
zyD3lyLazTFEgFCJ3FGOHP8G1Mibh4oKrIcyANYY16D64rTFiBd7kgACJxv9Z5FW438ZIj6nhH0N
9v1QEuefzQL+ynz5+AkkCa2hs2Okxwym7ZhnOxZ1jNjBadrR7yePshhiBr+s959r2p7TtDUzU7xR
eMTMOfwhIl2RuY8pLLr6bRNHQx+vDxbJ6MpwiCzgznSaaFHeZTa6figuCzX0TXtjwj1kGa8xLcEa
2M4ewjAImV3L+w0sy/RxZrh7HkwesFn2dY18tMsThEnCDNgRcTxZ/uostvlLQjjXRGL41LqgRpjL
aJDH8ejeTBteoZRj9tYe8Pr01TMKrtjdLRO4Z557azUven7xVW85XWLFib7xC/hidZHvKQsa4fWK
1kVE+2XMe+plxoX++Hio1YilixyOGP2XNBp4AARYX7FU4yQwPdFNf2RlTElsqZhr0tvXVHmiPGQe
hFL+nIdYMkg0y9TSbzjFb1HYpg4Hy26jgpTrd64CVdDiZgyiv2OW1Hi978fNP/G9TYeQ4VeJdLDs
ti/Ru7zkAA1yR1+EZbQaLW1hXB4ZZ3+NO7l7Zsnv2MrzItZKQOqKI3y2p1rAL5ynDNHyLSOYteFB
BcntRmNb//c15pvD1dKvAduJmXIXAMK9dvpIB1hB5v8RVFrhdjEHuwcPeoZwP8jk5BCcueZHxfhP
GkP+IlD7HTzGheqeCJ45oESMvQzpBif+gHS2XwK0OYPwN5upYTSm0mJnteJkvP4AahSipBxm0pnq
2hdzrYMR1qrkv/aXKAQ3/GoNKkgiA2rdeV0bMlgMT/DHu7AHyYNZfNoJPgxBr8cwYS98GIwKk7it
aLnjlf/xV3IrzvAcq1lLraYgaxekNEf2oh9zgo612gb1o/MRZN4QmOgEcHJHJ259XQMql8I6xrre
EgCH3xW3Tn6ZGxGnLHpv8y7QJtlwWmu9hrGarcAO7zk5Oe1JZ5zEmfKPoQml7EroZxdnzW/aZKzJ
VKEct8YqGwTaTJRizuOqtK7C9P6Pe7b+InQ33BPm+g6zq9Fii3q6Qnrd9M51pYJjIa9ajxHi0RK3
h7NxCXosLfxDm4EU/meB7IsnwBAiPcw5NrIro442y+OwQoxQfMHVLB0BaeVnP2JDd4KsbKike2QP
O3iPfdEo8S+iPQ8O00OnrIMUZQwboSLAOYnCs8nVnp8PQd+82Jg/gEE9SzEN/4HdJeSbbvTV0SWw
IKGM47f9oDBF+5uDKF5XrtwCU+0ZMISY5uniUngf+pGOBOOFpihxxDQ6dLr7q7wE13gTCBTHjVq1
gnBZmmBej70Efw7Ou0vuUQ38CEhP4lxFP88tvPaovzrskkWZU7ojLAMjAXeJ8h003CMgBkUM9GHw
JwELLun6mCMH8xE2lT4IgovstYyBHTBSm5UuP8UNllpG7M+Ocmb40H63+MdLP81uXOtL2VYmyhL/
FGNlYCc+FU6r/fwZbW2kclLsnRmYmVd6G65hdbkNK8BA7UQ3c0buhAdlEAtv6ES81cXKC0KWTzT1
wC1P5TDOWJmO/DRxDkFXaIq8d/mKjdfIkfmz4vQkgUnReYM/Nn8B+/WXSJ1UmnmTtZeVNlfxu9eH
Fw2V+68Sc6GMVnGTDZrUi9etnSVIB9gwCFZJt6IPWNKqQPHX7DDLZvqh9T9qlkAdeQ8HKJDbsyLL
2dXIxS5PtIr5O/RFhb43oSENMpL9lgDOW6GElBp7SLYY0NRECbhuWLqXBFhGo6h3hzpnnCVOVNr4
PV/yj3pDdFmVK1O2glpT20tDauJ/px2LyY8O6DouYPsIYTD5flc23eIOCYPqXthvzXXVM28iTjOq
nRj56ihhYxSASOWbOYHqe+FHDiQiWjZjOsPKWdgYdd0UcMgou0IZvrB0jrYvvqRI4fWPpY1VGJmZ
+XkrppNjnWwxVbn+EiGGYJnHwOgYSI/1vkH8+nFUoSfyY5/VNHFvq6CA4L9oSIH03krFk/gU55hP
XzD3H212zutsCPiL8s9asj9GAd5DCWPsryko8ZJyk5rDKbpZTeLRdEQ2XoFLFnk/X2f6xyWRPAqR
SzA3x9hx0vANeJC1hBfwg23+7iWn56bTaSjDt/nBOqH8eDepy1YR8Qz9lEcqxVOoz85Hap/Hd8Pp
C2Dax/a6M5A5CVdFrcoruHa9Y7AN2h4/t9pTneSIFwOCVQvG3cYfINgJ9mvmoFScwaCtanGf76q7
yPoAy9Wmznz/4qu7XNPXr8ZcfP2Ovj15C2Fsfq+VDKXtziP62P52Zek3490g0zZsvOhI9tzBCiVy
pC2tBDoINidxj965AelgQJHrkiRPgAscKnGmOsHCOnmHn2nqWMl/R3dKYZ5VuqCAk7/R2ZgJgTsj
YT/f0dKPPZ0D6svUHsk8MgiXE4OdNvtbvuVPcfBqT6GDaCFVdRBtIFdRRJ7fPzj6Wk2ZOGa3TnpR
Qtzss/jTfRrYsIJWUuL6pwz223A4aAIwzL792wQOekHgAN6Wi4FYELrIurEZzEVlpeboVv7VjYUy
n6nqqJe592ykBkcF+ZpxCA7OA5EcGbpgZWqJ2XLNuvTx+tVrn6bAjCpe53Vi14RB+xCbLrNlPJ8n
9ov5qDtwpOF62LNrAj1a/o5dpPP54YW0dtuiTXe1Lh5/2bAeBpBjqGaNiRmoYG+32QKkRK2rzWFB
WIyoZld/rkSoh0+ABlNRJcEIMj3Os3tX4AXZ+PydJAE2b73jQRFaLhy05ogJgihXkI6+AqizFFNV
ulqjpk8p58I7ry949l53WymKch8BMRaoKEAYzgFVTAiHaE0wjCOqPjVjOJbiLuTSLoL5cBQDawkI
WTAwjn4VlmHtt1oyGbTY7crJXNmVOUFcnOVNBsiOYbvte61wHFO9hE9pPDjrqqVNjL4z4AG2KAVp
5KGaGbiHr6gVSki2WFGo8XuB0+QCNd0KNk8GopIfBZCq/UDPXVYcLkwwlSidV+hC8RTU6CrIJO//
s6nXfcZ2iWTC4UJlLU8aavWgWmpvrSJl6C9miV8Y9eaLdEsJmKpgAvchrHXNmj7WlxsAm9wuc00i
kP7K0bavuQEoUtmxkyfZbegULqJY9mN568LPCaR0+A8N+LgViWqfg/HUawlrH/cJiBOI3vgf6BO8
Gw3zqL6RTQvCOjMUgd6f46G1XVf+gvS5oWHhyOGMYQwh9jvXfj4k02Rf/Wxeo0a1x2h4ULHscxzX
ahNvwl0K2WCirv8f4jtKkgjzeMTvKQKhiED1/jMQ6xF+jLYK2fmVl7EVK+XMOv5q8XYyIQrxHkq2
yb5Rv7WFdeKBZ9+vQm0T3UIKC/LSO11HvddRYIWO2xJw7LW3FSeCd+jXNdnmBbu6X6T/j98Zo6l/
AyqKAoAenlXeFBSpCunqqN5Kd0CSO2O0XZtAGbgfHVloG3S8AbGu7ev7C777a/YDFvfqzwjoJ4bN
rW6L0jS8oYyK0XTnCp3k2Ngceb2HNTY3himokznf5pGE6g0FA1++FUUyli/pV4QW+pnB/cdxD80a
f6NKEKULZUnvyiYzOz0R1lYmdIovIS23hk9NzrmCoYGwtlke2uyZA13wifmKftn+LyAfewbxOgxa
NCrBVv4Qq82hJkH+NpV+Rk/TK7WwB/v84rU9Sj0FweGDrSVdlsnj0Jz2wdo+y5e9+NbvxToi8zdK
cCEM2ora0FOxmO7iB8DahJwefTeOmhRjaP1EAF6/4VRMXqpd4gIh4Wo7bSr2yxraiO+EBtgL+C7Q
N/+9kVowzPIImibuXrtnT3+Zp12O2fs5vFWtSkR6yNAKpOf2RXfYe9UI9wC5Y4+V6yJP06cbDa3u
ARdtjCfw4Naw3f1tYdsoyxLf8q8PKcP2xFDtRZd5uyjXKFaObET1URc/ZyP2iCOmEVV/WsOjg9ad
dp4y0Lvurup6tbcVkNif20ZjeL/x3fqXbwyU+/w9hzQyxgm2TJWpBfHjRYf5g4U4RCq4jQZVK19i
FD55gCVHjck5YxuSdwyAYwT8PVaXJSsu0mYxSuwXDBAlmiiN+jTiG8sXCbmUYxn5bK2nq1O0WOPn
XGZeupgQOvjEKd65zVhTyiQSy9Pan4ipn83RyhfSOq1hZ3Le/IqpqMGXCNM3TyBlYJ6LUi5XNJmR
46Zrya3j8/E2NqrGCa9q12vBQtX1qQ/U/7UQTj/5K8yxVy6/HtXn/P/PBjHW9G7yco0Xc4ubgifm
+AEg7B+cLNXchh+v12/114e2cTwGl+Whoq2i44vFBjMbnfSxBtsJiqDJCkpuxtgSB11J6jfskK0E
Uh3Yf6e3aaOMfIhd/fNnhc+aloR/qZdKIbZRlTXPIOOH4Zm5X0eFvruh3xQZ0oTvGO/s6VOLtsDO
8++XsvHDwiJkkG7pANItVaiWrfb0Lod4cA68EU7WtA9fLADpYJEFgx+/DX5g7Sr8hL4e79JQyQvE
BZjbb3ZfbEs+/Czbf5GEz0sWnvLMEmA0fRKONwsJ55lJSUpES1Xk/KHcavtF8QMqO4yQZK7od27x
vgeIRI/xMLH8Gxue9jMkGNALIpaTAewb5CB9XfyXL1dFnteLhuo13ez2AtZYGxBd5qPPpD7fCqdc
bAwuHOpvKanqr/+4BArR0FjWCPPDv3wld9zST6uPsx/5EF8rTq83FA/optRh68vI49oh7b2ktxA8
Z2Jzm5aYzy7hTuVLL6DbAebY9RFyaDPr1emAz0Fk9MprzdO3fuFC3w5sHIKVMjUK1n+Q4cheUUiL
r5o9DOe469zUg4neZZJPGoJwkgG1iTmD9xOecHQ1HTVHnYquRtdUvHTbhI4ZlAR6ULavkOewgrfP
4s4g+D5bch6jsaYv4MfiSTALzT0/mW5jaKlP0skHO/GY+xruEhRvm/2Yq0d/dprYirEkdtfXb7hc
TP7SE3Fmxlg8d4JBWKgeDHshwaM+icAQ5kBblK+S4/zZo6JQg0SHnYvsPevb5H3QGS+T/YDcMeTl
tEboaidGKBXTHPFI4CdDJcZvnxyGbFbXdS0Of9/dFqQyAMaZRomZHWgZEyyhR71wVxh99rdmZ+ts
C+aTb7CUKFbhDqNBt5pMpoTYN7sEG+Ocjx5e22XIYc3yxYuXQg4uazevS4XtW/vvgJBYevuhQTzC
1hwhVufu0n6yCLko46HRYEDVjcsNVR24bRHjI0D5Q9twEL4Jy4WvVcdtMXfQ2P/x3gu1K7Gf3+Z4
wjBjX/JZcsip//6TKc+VoEbk9DyE8hiEDUsQsduMQ8+9LlPl6tCvRSWuYVTpQCzNFj4vgPnXTa61
qDZLZwz4sHFUMoiUGT5F81ZAdBngO/e/WxjXfXM2V2BOF+YXrydDD/XLJhNTRUpXHEkKyrUiG6tT
3yVSQPUFvc8Jj+Bt3jTiqECZ6eIiPh0RIT/KAiQDzmbpWQQVSXl/F9JQ7MiFhREQBdZEZ1XJDD4v
K9gPujQoNUwTYKCrux+Wplgcb8v+cdlf2l6bVePVxlwWVVMkjAjrdwuPez0qgKWVEZedCMas7VWr
QvAxz62N2mMsWecZnWjDP1bMD1hjHgNwErFR/U6TldXVnBcTLjkF3jUSQlg8xo0aP3T81uSKenSs
SLmLkRVtiAO2iod0Kt5Ckwnep+0AUaspOiF4Y2W03WjE0jY5J0iaB45VCjNYti+x+b/eLvlmRXfI
H2qk7e/NJ8Wx+74MqyDcza+78afah67x1A9dzFOQgp7yesRnXrEi9wS3gZU1occXLW9BVMFJ6BaJ
6XNPrPox6xqyYOH1oZS/K8MtwRwIhMSwsvlTkBw4YG5XLVKGJkgIwLFhvqkqrxJunpAzJuHA3so/
rwewyRB2Zn+5bbAEkufDBAKwKoQAehfligGLzlRyMMWsbcSV0HZ6KBRR5nExpjNRTrrqQhl/A9ex
3qPpFSdV0ygUrybsIOGNMi+84/AXm6JmQk1zCzmObaxe/i/JTi+LUhkuzcImLWRLfEaqlg+GtnVx
B4j0BRLzUd4VZjeW0BAiNxk6z5Z/uTbWUizh7X7VXVkDn9FhOAQMnyjApr75njWr8SyJHagPcL1X
Gl2LdzjHxKfUYLU8AfQcYHfikHtK7l6fZCXYpxoAFh4/gXWd+z3lrY18Umec7O19yy1vEa8ca+CO
kQneB3CFAZVXWO4xFZb5xzFRoZ2pINmoWdiAW4Z7wm8cPW1rWP8+OOdsYv6DH4hyJrd3oT/1MM/1
71Rm2R87+uu6kuYskiv51tfx5fTBvUC1NvIAHkB3sk9XU5SZkcSGd6SqWByRclcFo6PykmDnJHO7
p/FNuESlDxmLY2HWu2vJGFSNgGRpyzhC9CxSkiEmhFNJ98C1CoA4E6JlWfMvYq2kI7ycd2nxABwk
yYOnXWt6Dl8ApSSjerF3TJzGYBuLkr2greNdkcPe8rrFrbOlAKO6ePwR0HXS68QsKSWH2IYXPMa/
kCJvf+J8r1s7GrsdmKpDA9CjugFtq9wc/7dSigO4TtUmfp7VNjPuB6YH/lUnc4tsICt7zCG/2udE
vFkMSI2jPQjJ3argZKqjMfFBEIM1kcZFWseTBvxwYn+J7uE7nEW3mrcilLFRghRylwIETZR8UxDS
1IProDwUtD7NVGeK3vaa3DLnNunu0VkVBlpqhyXDUAu9Ks1o9iFilTCYQnh+K1fJqTp44ybRrYyx
Ny48/u5mz2ROSWMqwZPVeTYG4y7EwHBcBLwOrj7OixzA3dne9hU/QuX54mFmOW0HztkVOPstpt8v
cyGpiih+6coZRlCSD2mLMbc8o1wFZdr1kZbTtBWA8xGYIrs8K523Hvh29h1Hvm1JHhr57w0OUF4O
WCWvfK0mtu2n7bNPJ2vW+THS1spbBCi+uZkHZbBypfjY0eczsM2PdpmMi70XOmdL0AGboSOOFNTy
gaX026icPqbRyauxJwAN/PVWRXrg0u9q7DrPJO33TImb4dR6AcfYyda+CYfOg2dP9HDC9ZyeFagW
caantwoK1v4cm0djKKPYgaoE3GfvXaqV+SBGBg5d73agPWKgrOTnzeFdXralIMS8oA2fd/C/qOSG
qsFeyzAKW0t7rWvPUD8R+A9ikGXnoOKCq+u1GZQzvXTYHiMuJhKPXmgnpEgcGqm7NXN30nNvFGMN
49zyiIKb346FErI4HYqfv32/UDNEA34cuDFbdnh+gw5QzIYCbOWDBShuEUFPAABdy0Dt1labcABY
b1t4+IoBDkReTM4o/QRiekzmJn3cCeMCRkbMt8SDoxdWRhl5kJ685A5i/egNQqTG0uNqkuQUCGBc
/C2MWyMCDbYBOy1bzsNt7/aEK18Eu7W5obqydGgtJMCn5kbVJQkzed36GQU/FLcs7pK/GlfuJZab
4S6soB5GpQXEfdybHctOIR8F3S4MV+zkw70o0OTVT3Kv9NJNWFAusPdDDgoMj4Kx/Ypa607+3Y1t
jYaztr7vyTVxroXPcNjbZZPP/0EDaQNcvoaSGSdMrhYASLxhmh6IZg+bWmc3XsrMzYNpzHsaIw2Y
a3vGEJBDZ06fudRS048Gxq7DegxtsLpBnDAjehkg1kbHh5LxPbtXI4OiGcW0t+/myGELcgFH2vfu
RMeYxBA/xwskBTLyqDvv1Ev+7TnuXBUCmS6KZfPAgE3qi4SgzUfJlUioNTGX1D9R09Vz2LW2tJuw
pReKzyNJsNZTxPoIiU9EnA6i2i7krHkQ/S0yMWVHzqj//P5yxyOAe4RdNEXPzSs4lFYrT8HLcoDD
vymjFwYx8RSkJXN75EjFWpcqZNBnnj78HD1hOkw+IgB4rvqkblu9VzNNoQo7YLEB0sjxjv4Fgwgo
v9lq68JR1oh/ckVKCjsPfTXfMlRGgrKFVZd8ZeuJsF/tZNnqgmQKrg3doN2rxbxrXVm7durxWE9j
zVn4unjFKY5n81skoWwfnOkoF+Qb5fA0BYwWaz2nLuUVBeIxyy2OomSBLUCGBJvwLv2wcWPx8LuJ
iETpaLCXG3HMHPp3fEoLWhmrWPhHXEO+A5UhOhuxIYdfylGPSRFLqk0QZ8gd4eZkpE6uvbmuCHA4
llztshpFrt1GV/uv+DUsAtjp5wyTyIw3027L39XYnCeKtgwiX+ls9MDfNDksy6BiC85ML2fFiCDZ
P3ka4rK/0mAekmKBAxkBw3bcB5L2wQRTJti/GcjoJqXwY9Dku3cs5MLSUSgX8j5i9lNF3/9ND6m4
dArPZtAczLOMkdfWyYBPSp+1FeJXBL6BRfuPJ+sM+rFHGZCFbXUAcPnRij2AaEtcoCp+5uURFyfY
tjvNbvrxd0wWnSuYRODj0/nMkzw2iz9KKxIj2BFdjCk4ALwC4bYgkRYD5p4HH3wFh4OoYqGwYr12
ip59WQLKg7GQX2+wj/UyeHfgo0BnSTXOEZ41GEtuMPvnUPNMKvo/BslmP/r1A8JkgJQLGxy/9v36
pJOb0kUrvSv5zFXGGGrb/g248Gz4J/MY553RhIE3X0RlWQAGZt/ySvH1Ch2jQ1/XQJj5y7pKLZEz
QLKtuayWTgm6BDEw19Ng9J03bPB7JQFMu1tHLrzpGSt5JknuqoEwnd1SeP/OaCRBfkj4ewEgqRaS
jgTY9z8zRYdUR/hfkyaV1M05b+yaQRRyR2iTg24XLdGdfLJxfA5Z6xv/S9+5PQ92m74vFuMm7UT2
P/FwFjMfgvSWEDbHNdej0v0xPgX1CKwtd6uexzMudLTdwJUWfxpJhiLTFWa2+n5mH/+gRS1QkLW+
RbUqSMmEG/BO9sx1rAk/0znQYIeVALy9H3M01avVtmykCoVuXg9Od7hZEJ3rkuEamA3xMBAaidrP
ZfgK7z+svPrWMC5TLyVkjVUsyvGFuDUi0zT8MZod5cRO9x2E1+kilkjAlBT94QJtF01iEpxC9OCr
ep0gDl8M5yIwzfp5AieJ7x5+sPO3BUKgXlAmhqBhyetMqFy2cozlHRyieqRoIKXmVpiG2iXqzAkf
b7LWRocHoSeF/QBVv6sDIKQiwCCG5nCa9iXtJUNIww1U1ESq1uVRtO+PNwYuyQsJlsXkRIpFG1+K
llSZRiFBidLqVDySK/nLZsjuPCb5L51RuFZwX8Hf4hszCzS/LDeBPgPzj7lSAQks9M1zmDGYz+Uf
tN/0PYAkob54r2cM+gBLRm7Stf6WGwT2qYM9HJjOy8woD7Yu9/pi40sW4MliSR/eOQ6yRCCueHvQ
X2ValrPWaI7fEra6KRwpwS/jzcDs4fEInSVQsfup32ysByg9voVS42FjMFSXh4M4FNTsIUPQ7VcR
4hIsyYPlcJP+4fBU8QJ1HhvA8vA1XC6y1KM1jnR2XlFJGaKIiTBMglv6FZX7W72FTDeVVuh5THU0
8JH8oaPyJXo+Ll8mpBlP3Lz4rQe/j+nPohcd/zvF3XuiMN1qJYT2stX8miErChLMfU3HQk82Ci4O
DZBndOe8rH5LIpBpoEn0nNRtRBk6rQJbmztOu90WlWIMSsAF8euxwiV8qhOtY+L/HWNnKvRJFCSG
gXNVsF9//U+GAgPFT3W37QmN4RNIzbk1xF+4RlzV2Blm7Ntu6Mde8rHOm6/OiH45yHvzn7Z5jXgX
h5OAXOilf+keyEi/BqSUiTK+LP8wGP8m6Xve548a9vMVzCkleJxYMtsZJxOU3DLfamahJk8Mj9Lk
TT51Cwll13gWZHD8RANbrHFR1IjPeuf9BTE8auVuij4Xn6JNl1EngqPvhrdO7KJTWGP76akONGSX
nZ74ZQNF56sfzRwHvhknON+hyWf2rZzevCLmQaqVWDNht6nqYhZJ29LtQB0Tt9p9calo7p22we1k
9OfUqR2yOew57fcGz72co1IhvotQBDUOeEf4H0cgqNaxIbgtTn/H2mviuX4fb0ug6efQdfVWZ33F
HwA5V5y5wTY6Nm+8Pl+HN/1ygsWVxWkMLT8TZmmibh8953/9YXXDTCivqlgdrXrZ4Hmapi3oBP6e
Wy6IjiydbDXrXKpj9GEnNBykY2Mw4ozchk7vuB5nJY2ypq6QSejoRGNigMfQ5OteWBvi8aqAWIn3
jCNsEt91LStYAMaTGwIB/W57iNEOH08eCrEzt2hfxmhe7wvkuH78uTJe1IoXEx6JsDxyQFco1tKK
Dc/pGWmfhY0VDa5tXyiYHZ3AiGHtAmHgVgll7XY+OFdOcOb4zqyOr9plMlsG3h7XFlf8ZYXBN7vu
LhfcUHxNsdspkjKuvTxYRvdaVRoJZn+1a7uMLmJMTd8b0nCnNRgXGVLYgko9pGv1MxIV6rXuouE6
wy5Heqe0FR4mxk9ua3vWBTqQEin9vXSB82TU/gxyFxlPoTt5qxuC9IZOVSDplIh9Rf062OG3tzcD
3s8d/7wS/vVtFhaDIHG7Z6aIByVSQMmH42oXChbha6SPavDJIw2E9pVFYZYxvLbtsgQc0dJDD3qf
ai9uCO35VpibBSbZMQNHYbuaJGaWXarH32/gKslp4PXACQ/YkkFzU+kC4xBaRIGrnRK45/omSsAP
CwRRfyzvgosB85KuyIxL/bd4xFSeDgFUoroFPWtTf2zHLeMcEh0p7MZufRvy9BxOCrKQySnDRSNG
Xx9m98XNvDrvfk4sMrMxlkZ1LdyPqN1qCrFUXSTSVKT9QMmIXfY7ttUzmw34IkpZxHmOMdsO2+5i
7LyQ4CurM+ljpFC1HU1QzspUV6UxgYHi1KT/wD4s/UtPcSAgSJIUDGstJHzqQW4ahCZJco0xq4dL
8E5ggAkGq3q31GDc5OPHSGQwgmA0k7ZT0KqnNs5VNaQvhRz7GEFtngh+6rdRSOG50IzmNkKXGvZo
vxovkb6dqzMjmZSmuGGO1MuMmSN+SlzVkZeqE9o2g6b27WeamR4rWcN3jEMr5rugx+Vuiy5vhZVF
yIMXTyrxjqBcXiCg+/O3QD4hIhsWjLCwIm5gXRdmp8FWAFGBDaoJnRVNFzTyHpjxX/ed4KEnq9mH
q1L/xKRodO9ToG0QvpZameuBoawPwKqeFR4P29bal6tn99ArsjUN3A5ittRqyoxEXNs2UspaP9D+
T8oob/QJ2F7Dmxgl9wgR40AmXgdUPWYBTMOO2SCaFrO9SjQyAe1F1ofBTc+g0ESxM8cxQOnoGVx4
TLKw7oC8ygIHu96I0RTCI4fky6qbLipS5FIcZyeEix0abNRhRkGd04LtMyHHr2PuA2/0hhfm8wRz
9lNjXMpZksF+ceUQlytQip6pH7D2W1mkt9WTdCfffTGjUCawrtfm9PhH1bGPDbH15yCz17dWwcHj
LYKkaAUrigfw5svGsfO/JrIz570H2ONo+U4+d+m8tg9CMDu1NaUdMUpUlLAJBg3ITEHO4WEzN0qG
SpzuYZ51K4zNBT9iCUdMBDD1JuZI4KNzEl3XW0jcy5NmLvDbWsUDPjCqzbnn0w4lj0WmK7pq11Xu
K7b5Xcws393c8AopkPbC6ORWiqXFcz6YYUlzzlGKpR3u5tOksu2hv1vyT51d2raKilzT6rMfY3JE
3K9KQ6lJe28/tvvD3GrZQRq6+goOtIU/c339C/Z4o0nIVDaMbTkijh7bo9bmjColRX+29KMKWUgd
NbcdK+GfyAR3swd5k2JItzSzuPvDJJeHX0IbKvJfs9mkpWoh3jgsIw/5EcXcNoh+C/WbBnVult1J
iWJmFzSc4SrYEkDpD4NVtgZJ8OnIqjvuhhQN2FDxOny8w2HUe3DhrfSHkMJuZAK9Cd//9oD3yUnj
Ot8rMeWoSlxcRgIa18jzDL4rNjkKATL/nLz9uuazMLhCx0Mj96Ubvjm4Gmw2VbrDyj5rUipE5p9s
V3Aixl9c9CRLc+Xm+BoHuLDQmk91YirICyKCDX//5VZvtWDlbSV6Ixue4wuhVmhnso5Gj8PHME5V
kC5UU7/3jJ5aKB25f2S6dJxFHZPIS6pa7XQ7ehNoiw16cE/MgjtKHOVRgAqGYzpCi9/nP26TSsJF
j3ceTa0RWBJcYnTHbLx0ReUQtHWq+oFENja2VMgpf6qirLdR+I9FhyCd7d8fy+zP/0VWUN/VSVzW
Gmp1O/lRnKfgVoBGzzbqecGo52Vi6TtIAXrDCDFf6qXaIN1LaRcbzdQV/MJYLtvMtgVqABRst0Iv
69p0vZq1oYLEcu+ZkefEIrgoiqDCAz5k6lmsIPlvMUHjjBvsujc3+X6iUaAopGe7lA4Gjuhtv7ke
oqJwzmorc7vJiDNueDYg+HmMVHdo5RQz8X5J3juAVoUu8H/rAXsJXf3RXopdqzA2KSvVnO2db8cf
PAFF2fg1kaNDya/09bDgAUphVF6lYCVNPl6wYXVKDRJsOf4X3qhWq1LlXNtY74uANmdsm3gxLHpe
qHOgws1aYA6SfWLXP42bakr827UrEdwYImdbVX/xXwptZdE+Ghuu8J19/5JZHy7ZLV35yRBSZdMi
Hdou6RcVuvYsjQNijPSVKXC0KQ818vh0DOliqlXbMdvffR6CZGoQSeQQLGKHVY0NYZpMHb+ZlRKm
kuC8CACie4RNLp94muZGYfhT5gPYsSHsLKlpkgtiW+3+Vlb378ejNrTVJYzAQbwDiHiydy/MqUQL
TyxMj1iryyzidW8DzB4v9aQqwx0tyKMlBKhAOOQfztSioP1aAXKxVIw7vBuE8wPllF+7tad02U5w
FJG6EjgK0fIvujAdPJeBkV8TF+K1XGve9d57QtVZKIp8e27CJko2gy6g94iu9yGufeUIfv2bbby5
g3bQurlGK5FSPlaYh4YagS3bACfnXob0OmBVATdD8Y8d+wkW1QWHUjvup+9NJFQsva5EoCnQ9h/l
t6mafvSIvduymAjJyQBP4sgQMTeYRVvrgAh4+bqTGuSlxU3crTMhSdceS7s95xOaSva5ad+5rno7
zQHuCys3ZopnnVilh7Q2rLZQYYoKHSBRMPumzXDzI0t4ZY6yfVXnzcli7/qCxvbWjN90ST+2Avl8
Utc5OZtn74eT5ApM8Q9BcrnbCSEBpYwVUR+ffSB455JuPL+EpquSB8kAHNrPgi4zYCnkTb7IW1U9
33WQB4Pf65ddDiTQ1VksLyXnZ7H8CgQlzamv5mR/AzvS0bKhtIxOd3w668TWKfTqW6JpPYkHZA3/
s93RwZ0Zx1D4KqxTzELaaekMRHwnnfRLaKzef4mGr/Ga94A17Zt+bD2ZxFPxoGbeSot147kotP4A
v3wKPphLhh2ro1aGpX+cYeeTax6Xy0FQ8X7eIR1tIVhdqyJg+djks+Y6qwuVkVTcUR2MQ2MPoBjY
YewQO3y0jGxybQ7b7wnIj8kpVhWTNJELabh2x9Av1TIvlaUdZw+8Iu2vHu/jhHauBGsTQJ8u2jbU
KrKjkOxGfFox1NhnfK52MxxXFJ26um7sd/WhvzkFQ3YwFs/diidA4W56/YDb2X1oGKmZcHNq3Pok
WJ1thyeduKM+anS2ehFC0ffFjPynks6ZbtPtCWFxCj36D/XMtTov2fZeOhLc7bV28bjnt0i0cCLU
jJm5FA+hXK2zaO8BHehsoC0QJ4JPMGnmqqOepvVRgOmEPiAOCpliI/2zGyD0heREzDlv9YoLwlib
4QhWXyH27lvCjsZ4uVw3Vb9HSVoa4PHx0W81CaqLj9UAimtq4/8/j7qkSL3pvIVLkHW6vnHq0Tfc
gBy7vh4hO4psZjR+4W5ocacbFC7qBaA0AqYRTWC9Sa7DiQvoun0XVKwlI/9fYZlqBTNPgOiXtbNx
yKKy/Ibg6xE9puqoEOWQXgdQoMftqv9SkHKfKpv/gcYzj47meFJxKvziI8q3/d2BtxoL3eqFjL5F
NDhun/kjPJzHwGvqErbbmlZXK3lh9Doaf3TpH9w2aymz9ha60u61/meBWUObBpcIz323uLx+EkVi
8PIs3HAsRmIoKZ/O3JJPxcotrp3jsjIG+tOfhQplSdpGie2xtK1+qnMJeyFcr3FBVdjVd5xnzwMh
D3XxKfqDORghmau+6DkLbzKvQCMH2SZ1GrmgBzSFRJJb9sOV8YoHjJbLcFRXOVDyQGzRuQRczN8N
i1pI4k/3Wof9r+5extLIgX1ghMoKt9KIFk+R7KiJPn6OpovhxBtRDpFbr+4OLzmGiv+uvF42URUv
qZM1H+pOycEpoReL3IIbTOzu5HhAm9gJBg0VZHScKRm3j5OM7gUWLQ5bhV1kJGmrGP5B5ALPeFdR
2vfb/5ofiD+3IIIGsFvwFg7GOb0ssmThit+73jGyoHGW2wst7wqBYajL0MFzKh6N87FhIMhKSXKo
AkrHg2yZXCHQdQ1Wp7ramYz+Ez0fFZ1s6uJj97uyMWbT5ycPprngym8kc2tqka2Xxb8iAZFToy0/
uS6fxCSePkYWn3Xx3b4TPfpQ7BzP0E6FCydXLpTVoAckNymMfTS48TmTO0ORH1sz1h8Z5BrQdil5
FWYxu4Dh7mfIETYLVhjgtXVPW71vs59Jgn08zdf0BmEEL0Y7/SxcpXHNqxVYy2x5BfshSAFoCOUU
xHXmb+f0a0c/fYxyBX9ZrEL/wqmWNrOGJrhxiJV2VzVkOXlYBETyPZxanfFhSTUJaNP0G2qS2nEC
UqaBWCddBxRcoRNglWM+5kRLHuxr+ZAvOmi9Ns4qiHpgiOtPGLiyJB9zXUTwNy8KaIzIEzfBXC34
yxLn4CcFptfk7tuNzaneJJMJUymherbe9XQVfb9xgsxC3RGQzEZBBTSaihltYZ1Aa7fimY/23pb6
rAVnA3ikS9vjjVh7UP0C/+nmbd3aFx/oq90KXhw+uJylpWimsQmT0inIrkvBfkaMb9gYFRja+sUi
tSW8pmXjcOCM08MY7Cb8zQ2N86l3QarZLGGc1TJF90oqdyPl3Wk9uGNrTXm5BS/OkDQgEE6LpXIN
+76NrtnJqIDO0Bs7fVFlhRWebR76FNY555J+ADTYcK4/FLhYh3Ie8aLoBuBGvZAfudeYV3LzkPVJ
u4phT47naTrsrWOP/VvgApr9w9Gkz5+ANWfwc2hCh9cO6YEb/GfOR7z6BOQGPmeElD0vqQ8szLvu
z00XE7rxkKOrjEwy/y9vkMbvYN9QM3wVcddmg3aRkJ1YVr9P4CMfl0nLyVpagkj3Q3RCtSn1havt
jpc7cyVxSgRYVgkcGuNDxks89oWUmgzrSBMci1UmYi/8WxKzfDWP7QIM2F4ibR2VR92d1QPhwxnE
iif2XC2C/xqT762b3lbMWRyskjjekljchRDz9PUqX54W0vzbZy9CuojD1Jz7yspr0Z7XLKITrKsZ
sQBUhaXPdJCVLf7DVSk2ylIJffkVtp1YyuwAPEaIF/5dj7vmd3TzVTYp7u0K43ak18jOEn6kRNoj
BZ6KXdHO7wJP0jKreomn8UT+HfS/GIiBLGaIf+/V0ksF3Ywyv42n+G83DIi0nwetgaOop3VrMT/V
pxXfa93N1rkV/rPFUnnrM8yGn9OIASAV1NFoVgndnRpx2JwekgdxtfQkvZovLROlLza269+TRKB4
58c95fTMXrqIP1mDqwjB2t04IJlPfPr8u8CDvKPZ2Cn81CcIG0glfe1Mvy9s3tNHlBm1IeLYAtnu
0L8jq/X6jgaPGx4qE14Tff/U1ols+ANALJMlSEWP3qeM61lrHU5Ji43cPrvsHyx+aegV5L4EvXZF
zpVkF4AHmoap9mFSopml2lRrlJtAyrczOvsYkaPCdoy5aKcPIFtXHtizEkZ1weUm13TunA3IymtL
E9hpoAMLhUegAqAc7/ASp2ppHmj/XJBufP9ENH0kFH+lbddYA6IQJ9zkTu7yJoVYm0Gd7qLoPngD
T3pn16g2eQch9cDUDmhw/MaAKcY4YDmmi8f72d9ti/TQG37fe3JDG5+/+S6qgYlb9ioNAxWZR0Mb
U8zXUFsGBMqvIqs0CvWaJ9ZlLSMkStwQahwi+0Oy5xkCuv2/BO7SiIYVxSD99BYvfozxEhwcR5SR
22kPEAktY8FZm5SgjksvIm4HQrj5THKxXt9Tm/dsruu8sZVPQ7rMeG4MNoJrRopHQAmpBBsHR4dI
pFF8SA7OHDRSVRp8XbY4bnHFh/hGnAKauvxAVngS5j/9hKA+TRoBpVvRq6H3cqhrBBZaERtLuk0p
dkEXY9GzpRrBuOXtJgBSS/RqT+N0aRVmdkkLuRnvUi+68kp61agZjYpbhXztu7iC73SDNbXFJbyt
6cLTIkTTjPikAZQRFFSNh8xo2U4aCTDqLEE/qCYRxheUGFjOYYdHwcSqL0ZNtaARL8h8jlSHbTqb
GZqEXXtNT6843QBBjviqOg1mhup54QGtgNVl/c8z+/Yo24Oh1CKWo3OCR6MuMP5k3BqB7SUE8uyn
/8G7bgNGdr3dRY1vs/v7kdVKEf2qOZmsZtem/YTR6jh99J+zakWqE0FRv4AdhMBb7nWd3/ieHipg
LMRkI1ziPPa0XBnxzD/qCVNeGTujsiN8Q4ON2+Br5ujq8uZydN1ciThkTS/TcxEKZxpHO1/wtmpR
Hn8I15MkzO3VAivU5Gn9oCUJB8iYi9199sIHoIDMjSrSAPuoKfLcesQ1uuX0ZB477Hv2pL4WxFAJ
dGSWz5a+vCV1svy+B7ozAX2DB80JDeGfG5OxPeT8a+Bx+DrFJFLwaiP6HcJ6QZlWc0sxxEq1NeoY
ySchHKPYUoGlFzPIbDFgl17dGXNTdqXA+hHYS9zxuIpOVQm+GkX0auAAci4S8gY6nao3fHPq8ZoX
hifOxvPGA5NBARDarouB+ARTr/TfH4S/QvbJg+lQrVrxKU+7V6ytDo19aQ6m4GDIQ+w89yPM4wx3
IAG3OCk8khrczjl3RRW5R5oQIPn2+0WSCqxZWfsgspVhVXtSm5LWjjZQFy6AaNS6ukaJbyLZeTGs
//WeLa1FvtCeJiNvoMg/BroCAyuDy2dFCqqBQqBmxdu0Of3a8vmytvlpyzm1mA2Eo3sy0HE0n3n1
NNz2MdnYmtnL15+DxgDun5+SgiACEFVxbYnte9TDMRD2fVfZQSfBeHDOKTVsvDvZA3HpnOMR3NJN
jBcci9e+I4ykddapV54rHPswLeH6gzLTuAfx1ZOTH9w98hvLVxLlP9gXQWVq60qgLvxcVXWDeMX6
q5uklw9huKYcGdxaudV/5zTHLt+EI6jOj5Hqo+9K3PPVusPtoIrfFPhZuGJX0I8a4Skuc2GtVusO
hE3hXpmikd/sw/wZ6hBWo+CcZqv9y445oZ3S/ihJogm8XNhpmWBcls80+Diac6N0joqZc2kewL8A
ED336GMchGHjblss8kfm/RugJTGtMnojGy6Cmy0cFIycdR0pbcP9xa6AEVlKAkHiVoJsZsS8H9zI
+9GQ/k87OsY+ZagxI5AlciUGG06xKXJoGXTdCGTPEhyDl8RzN0eWL31sojPQBlWzuvdFiJC3Z2Uj
dWOyVeWIWDmPh3VgBX1O8LWA3+hsDj4k4uFN8dlPdlJrWACHuFrf0rWLxpSV06F81qjZmVLZCGBo
1H+NQm3hHoZbW1qmMkqaS/yvX2Uk5EfdAh628MaHfLhFsvUMkhKC7b+5o5dTcus1QKnDl0DGn1Lu
3GQXT13X0bWhSMftLnAQl1yqo5qa7DjFLEJR+P07yFFe0PNcnCKU7kfN3HQBDmWkjj0ipIagFwLv
/bAuv2tyzth0uKXA8ofl4a5lgtvcORVtJwPuOfR8nGjKx+mvgmnWqTORLkwA6p5lvEEHZ3dbxvoZ
ud7NuCBkuE+0X1SleDDz0HOOEhUaY54LLL9M9+RWgiyK06KoQETfwLWV7jN3BkQYLqqxW40Wdp/V
1629tsnfd4YyQhaVVFpkoUUEqsdRywTb6l6vaSGKPdJhg1sZI3P7FeX6Tu174Ge4vWvNzBjdBG7I
cGJOmPiDUaVPy6y0uy6BPxc62IUOEzXUF1vhpQ1t1BJgrxaZYVbPNFFRUup088IDLd8/fEh7S+Hu
wSk9ywwgpAmS0ZkBMo27BnVkBKS1yihpMOs2TwSWMDhCFTlwvIZglW5+nrWRfeg1Z3sT9zf+QkXU
qSSqUS4lGsaCbxcbgQ2u3IO2W/HnOjsOTLJwpv83Qd1A3uh8NTPMTnG2zFwc0BIvbsw9ejIo/eYN
xDjjeWK3XrPvziBf95a7a73HFKlfxo558MaexOR2SWY04lSyz6qb8PFv9pccd7ZZy2rTrf2IxhWm
IzmafV8gL8kBQbdO1WLwbld3b9+a92NLhgvXP/rN1U+kakB8DZK+o+7E1kZz1vy0xxnXA8i5Uv2b
bb+0WuUTAtR3u8+6YfRNZ8qPTcDHnXk0Vk9qctdg6L8IBVlspOw+BwkhfCC89fpPYf2AXjYFHBEP
N5PYFdAFOeGniPzDPLneKo377MSTFMeV1rfo5XErINCS4L8WFxtj8Muji429NUOxrv3xDvWr/4Jm
IPv3OgHa1VOClvJrGN/mPd8QY2BaUaPHYx/Tx+HYSssd/spGPGJYxoYPHJh8cw8x5N3nhzJuD8Wf
Zv+JTWUhUSzFnGuQmzhJDazYCIOFu6812F7u+oRKAoAlPYhvAsXf/FH4ZZ6qipCWZj4Meu5JWiJ0
LVHQwYbfmosuIg+zHAl/Mx6nXiIzob1+Hbp1VyZCKX4q0BghEbmaR5LiAveJm9xnP7oqPHSn/MFr
YH8a7ThaoYqJT4l1QQMwjClpt+tK+AEoWyr/8FeCNqQ1fUiNNGUMNcGLl/jT/eqWPNhwoHlhrEbt
NGkYo/hF5xX90MehYGo26ybfsfK4wWPe4mFmqlmIWQfUtpugF+26t/qHoIf8HUeNi1RWapxRbSLx
Lcg0oob0tq/PyX7cwWSR/v56MFN8Ext+pkY9rKb/Xbhv2P85U+8VEuoZc8IKzcg3VUxgbxALXOeX
6s5vHmRUuHE9EEeB94YdXFiddXuykvk1IBezmnHbz8S/IMc2uXpKWG9lJv+rvlH34+ntwpMfuGKL
Eaa5LDFGaVkt/JM9gHbETWQpN0K2VA+J559YQAulVLEDdjVgF013xpArrkCkcbM4OgUrzcxXInKE
SIUT7qEGCd1xEO03oc7A4NOfUGH3Lhkbr9+F8rOtOfqyBDf5XwIhNiE1Ypatjwv3FG4ZxpS5GOQ2
oFnBUJVZ93lwnc5wYCcuUXGn+3by48o8lKCifXBKbTaHNaasRsvgzLWoHX3vV9CrjpIsuIvaUgbj
CAbHhqome/57/mU+PTerAnCVLC4tMAKoyLh6uq92TSZb/aX85Olok9tnnch/tsNtC+X6DEdO9nDv
BerSFKLvCTOh0lddtQugbL1yLa65h8B19IKEGJjsAAiLy61iUbuqg6D5UX0NqyiVKAl/7U9p4pmV
B9/TC47VFOxJEsajm9PiyX4fXVV5H0gkLNVSlYhNqXs8z+U2HFsGVadbCdrKr5e/WClCnyUZbG+E
TRjjw8mjbekKeN+i97eSEPUxaJrTifW95S+/FNOynaLoIUFwwKy46bNmpW9wObyW/EyanabS3QqV
V9iK61lMTxxHkS+CvF7UEEuiC3oQUS0sQJnO2bTGkDgg9CKfDzVyqdATCNCHandoURuxBAqbz8i+
ZQ2xoC/cFYVA9RdGFf8zK1rh/N8G/pGMXtpXT+eaJlqvywF4qjS4BdcEoc9LNTZ9hg1IXyDVubsH
Q5RoDwSIN4ef0Um9v8NUnsg1Fv1NeXbq4K4C+duesGoxdHzozQXeNq1DRGWeu94NU14FYcg+lwBW
FfPQUQIAVUNiPRoSPVcfq8l2PzS3P00FtOVvLgwGFV8wG6thH16ykUtIH+iaw8WWPC05+Zjr2YY5
h0ZRfY+Nusa7euDVYSoTlDvzkFC5XYje2zek8Oa0Hzp4JtRouOREyYk/Dv7W00ZOT/NXJVglUjrm
dAto8YuRQ1O773LotfhQYLg/ozLoBVcsuOnhbsILOcnywxaphLOz1p5MExmCHYSwdhG53dkXcxf7
mnweQsBIt1kb//8dwrTKdbFdVRHyvgCcW28Yqw/5PtWglr6elVEjVCAWNGrN2rQdnFsHG1Hkxcrq
jfcg+y/1x7KhlBWNy3mU1RQ5m0kT4ITePd/E7LCfxadLlVVHBmDBTMKriG3gZKWh371O3NPJupCT
yGhII9AvevdmOAo+i50Rb2/yzyWgLFzAE3kijz2e0jCr80aV2AV4aOWSI8BpGFpv9aHKQBINY9fE
XVclJ7TN65nN2gDGSLiAnrNa4mShVJ38SzOT1ysm3uQwSJFuwjiSCvK98a92hZS3c+YjRpT/Es7w
Vqbbr5FVj52RTp7dBhq1MUvzd1bMTrGSu35251Yeg/Z85aWvHICaQ/uXidJ3dUgpbotYTp91vlYm
ri8ELslB60zwomy2m5MC4+gbDaKACJIldfDitLjaHb6wwZhU6qCgvTgScS0qaa5UlzOS58cxIJeq
y7nvBivLfbrqiLvZPomI/rfxinERbTQK4C1lCJl+DBxh0EEE+2394+rmlqHS22SBUJouMWICBS81
c9e4rZuCalgAKz5Dbk9rNe5aP3SVBnzIsGZFcAMo192nOTaITCCYYQDYIO/9g8n0B09wl+MxjBf/
Rs/XDHKHL1BtIPyrAv9AddTOwI9VZowwQPGZzpKrIGvMWG1yHGG97u+YW1uM15MVWiKGOg/rh6M6
24UJI75SYW+h5atU7IaV/0HpdFy5tvKCpFgdWNaMIyOzTdfw4xRe7Qo+2gvVJufRBq2yVtvb+yqP
t/U2PWxG6HiPznkJBW7IwQtYAt3aydrMEHTy8vOyYydds6llzn6bZwIGtQzxYTnx6TKLc78b665w
umGkiBnZ1VuvFCKZbkG/poJOPjMV+AZXDD7iTzaRTealgispKifpE9tbrCgCTE6BhH7kKlK55+7x
ZgmGqlUHJKadchWRQYFLoZ9CleaWp9t95Vr6w+t34DGhkYYZMdYevTKRLnXPwgInxYx8yyyBEV+J
TMEvf+nnuCA7IiZppcGVAR5f8lrYUlyVt5TaKgYTCsJIr7ibGa6fFC256AukNvQTu63YRwZYRNsS
XoLF/M3uzhWsEul52RVBvecrWbOOo2j/XaC9IUV3RAoxnFm+H88dBLMZlVaHqrMHrFMPf284lprw
/9A4E7LIH9cuCJP2zx/34/FmmN9wKD87nq2Qr7cIoLBbrUex387D13vkpw9Gc4naDqxVbiIKOkUn
nRji/DPCFZa4XiYXL44lgi2JQZhamtZaX0HdbSE0A8SVrVv846C+rxEu0UJwus8epH5nc8P4QJQH
ju9SCT153FX4DxXsqtrpf7SAO8LYCvgriWch0xmzrHW0JMXd8EYB+UANtvSkeF1pFI0/yRP+ECFq
SAtHxgMuOTDwW0BvYdSFNL6UAxuH+8XZPCLl+PrCOfjAL3x+rBET/EkE+GseZS5Yd1EazGUDv+cx
1vkTEOzRc0y03N7l8JHHRZPlS//E12tByy5/nBKDhAyi7DvE5m5ccGxkAB7XmlCupZBhFUEQhUah
fKF7welJvYrDnwCJJQZLfARhDM83lGzr8Oq1hrFlTZJGAaUP4USG4wVNRggswzBuW0FfJbKvkTbk
ZvrVagv41vPs5ePXF5JSGjwk+kIqCtAozAmJMI85+sJeMWHYGltmwK+6HTEk6KE3tCWblwghS6x7
UpInLJc/FUGPgvZm58ihx0nGzJGVPp4+xNX3+Lcb7IySRWTlqP++S+EJxkPxc2UXKG8bn134WCAz
nI+IJjZk6O2qyORyV6QOx812mWvWf6CTCaGQg9hYUsmgxxccGo9mN9KoaZujHPvIG99zYfc08173
EFhRDacAYv89MtgwlObkljBRvHabCp+iNyqCb+q7+GsrU8+KWh33fGCh/Z1YitcUo9hjUU3hEhsX
0/bZWfppC8HtsvWFvl3OvmlZRWl9qpabhKfW7R841i5x9tiUA85WGB0fa4nN3wGGP33OA/eZFIey
dkdQ6hZwRYmcWDBpchDe1Uq4WT3auPIQSYfsnddRO1NUeLnrD25kSK+Af9Ovub9q2xlo3nmP+zYj
Ov5B9LnYjSvxAnfogJ1za4RDkIXOELb1t4I/bHdoy0phAFIXZrJh07+T0+fHuP6qIec+qcWd3do7
+BWosASNG4axxJqcCg5z35SRQ6nElhncWhZ8vije30majztlf9j3sphnJP6yJdfOBHSCupk/Axa1
zmqP4Mdozh+TWdnWU+qCLKZh4dvba2ALADOPi7Ppm0vcM/aNK197nt9750P2SqghVevtwN6sf0cO
LcCEjhIjXBkqbDFpfDdPGMPUE3pQDCN/NLtPfUfcZsN/JcE6BC7Qqb3jB6fh4SPwglemVWaEyH0U
XY0iSabZyPuk0vb8xwIal7HI8RTvWzb3KKT7S0CC9HzbP5K9PCaVeoRtvZwKkgYFSzQ7dsFOYIpr
LOxixB8EQDZ847sb3pznPHlj2oLb0RmK0x1xuGW4xMcP8ubOf6m5k67eK4M/tKEH0/djNvjmx13/
hACjynRbYT6L9FCrUltagFRqCBQucxSnqNR1eSGNFSvAfDSTsH9z+6RRhuajtiE+FSZsI1jNpvTc
tASuovFdHZ43lgpxmdYqrUg+K5rxu4Ep4yc2bVNQSUvxHZKNkunT++TQA3IbIRq4I+vgThuA8l2b
69jW9qXBYJOcbaEKWADPqvV4lYyuz/n2UEt1BPDK3lZ4If/1Klu7wKMqS68EzlNVLGSw+IjgiYSd
evmw2taRNgXCujU8EBv4Fk900E1B3ty9PnbUAF4OZq36SUIu+Lo/N1KTdYGucy5Z9J6HTQ/OrExA
LrrdGh9/KYyAo4sN85MdfC3Y6CK2wIeBr/5vHBVdftFabUGJ8Zm3nRTJwhJW02z62vY3itL5QmDR
tmlru0TH3nSpr5mtDvwB2FjuEf2GbmHF59z3Li6R864oYl/J93h1Rxdxi86uQO9Y4acGXx5U0DHz
dMDURgOgaGDsbomxmTS1+zcSwHVO4fDU3n16UEpK+r188oCgMSgZPjskDiR5fKyD7Q26ZCC5Aqk2
EdvSXW6jueV2Clqj/+iTIOdhccd6YQ6c9tBqJM1cwfjt8/mnaQxCh6kPRv5CHt3tw0alMjonlhfQ
em2yQajFLp9gVoBjQbyfnyfflBUE44Udv5N/oFRapP5XJexa4g4BY5Az2D7xWkhVqgPMvDxsgylx
sJSH6+0RHIZKfuBZJRXy1/SbRWrDq1jgVhCb+KegzqQUykHjIJTbYWKJqZWno7L+Ipc6I58U3+Kw
E5Yzl0j4ykXyzRTC1rl4ljpc7BoFbNy+VKsoQY8eh6bJWaU7UDkAmPvvMVZlC32hlSviBV6eworp
7AmmGiP/errk+qTzT3o7EeytEN+skpBylGhZF0B6M3MqzhN5MjIwrXPopypVvqnXE00KggdFGcVR
EsHJbQYI4+o1CDpuFlAhg9M/F2vij/mV+ASyBhH4Yb0MvPPUx2XFuxKLgbKt1ryqAnCsEEyQIS3P
/Mts4rdnu3P/ByLvCePFUjD28+EtuXMvqqOXiN5qCQQv3bbh4VqhLfqiJqet5cvIvZgPZbPsEACq
UhEtRxff/czn0C4rwHvzAzdlVh0DjkRQQdyzRwP75pviB595pfrhR9M9uhhcZ3gidFsp4lWf6Bqb
Demfx5Bbd9GbBKIkH+7XePXd3GKqzKGuLuQmEW9uREwmSt4kOr6IM8OAguPVRQy6V88yCYNqjelu
cPZ+5A+qDNzaYxrW1hnd9XO1kuL3gJaJjPzGUblVv4tZEVqqWp/EEcOpsTxtKvex+RwnK8yv+FDh
2ez+DqnJiJ8Z74uezP1LYbrhTv6PZyI/pioyBi7WMNEXWm+THPN4HC0Y/e8hERhMAdECS0WuEgd6
SsKradUv80GAJrbxOR/tDJ/xu/0fiJ5oidj5UXVXX+7zaCZVUDAxYftlCgtteYEAWjIeHDdcou9w
x6gDUQpdOxkK5MlftW0UqNWMx1LJMCXzx2hqKRGHQWx7Dn0e1ULwJwTkTpLpmFAraUjFNQiT87qh
sFg60m0i5jPrT0hCRuuu3G2quRtnTQUOxCEEE+524iR+0EW1tkGbl/6F4eBJdpyEowVxUqzAkWrL
W4kI9y2QG6UgXMY9N11549Isbhe3JSgOBlBC/NjcM2Dr8g+ESUqFz4hF1vNcFK+ujfWNx1T0pOiy
UdM9OBze649bG+1VQwoVNInQcG4ZDlTe3Kaxy0t1ukC8nwZaM5ZfjsQfRSyiktV89n0qcmXZLPDz
4Ow3WRBkMcn61fBY0pAIVIkI86aRDSig2SV0mz87f8AkyctIqaurwgnGigkvcZm6IJzPwA0czWrh
PN5QZwd73tx9+WpBsrNGNheIihtkXifenvn+U1NGKBlF2JeddIysVZMYle/3TUsTNy0k+KKmNzAU
b/qZSGFHnfTSxv3bOjpUTHNtKZeBI9lZ781DHEurtK9mK57yxwspZpGJbWX4XysKcs29dJvbCYI+
ohXjXJGd5e6+y12wGt4cK6Vi7sVdv7SRgU2+8/HZtkB9x69xsXGMDqu3L+2xBZw48fduh5Bh5T60
0SvAaiMweEaX5wswfFuH+OS37r7LZoF5uDJhfggqoTq71YaN/y6wWto2+elQjANp2fpJ7d1VcZPo
8xsTxDrRdlUd079zpDRyJ9I9YJEF9xiCcNeNGUYnd3WT0phu3MkqGrBC+EzhmHBLFl8fF7/JkJLf
rvrrluOAlNGL8385gY05xBcOUi0tSg8+cYxS8iVpBZxbWzG1QZIoQqKRbUS5zi6RpSqSYFB5XK0N
K7isKl628B9nlr4vl9E66Uhtcj3Z5+ZVN6nSGoXyrSs9vCbAtz1Srdm2UxL+rACDtBaHli7sIEW3
UAE3D9a31aN3WIPnKv56hs4NiQidU1whFtzKTzOPqGfLlNjP6l9qyrpvUg6J7r7UCiwEnK5rkLud
yqhyOf1tq3PsLJfM6b0EQDtl6rHYC0quUMWdycKZHsZaGwP0xjkc9rEPLX0mCyN7iFL20kNtw/9J
WVIDGLGNtLh8/hUCa2J+27+56aEmKz1M3tXmv+bhzdUnXwq9xjxb+aXofpre6TZiM52AULkLFCv0
umx4BENmhNciIQFIGQt3kRVdHypIC3UFhew31Ff3qpHVAIVsIOOy8+eCWfenNVRv4tolgR1lWBKx
1Fxb5vIhCXIrKDpWFsEPhJ9u1LjcsV/8x9VaWO1mDXXIAq9xsWAMEF5VLCfnR7MQoq9hZ1BTlXlJ
AMto+Pgqpow69bTJENBsOfUxhVCj0teGjTwzWudiiDnV5MPeFeHdbSQXVxrzT5o2tzISDqCkgfXq
AIhYBjSHnBb+NTERzPa6Lgl2YSwPgoioqNQ4wE9LENrVLrh0IdNRYmc07ErQvuvwgLu/Us5wZjlK
pSR4NnJg9s4Gu3qgy2VAG+svrVssGWM3tiNam5wclhWxzm0uqQWUroJAyn1vrox4q914gUeuPutI
FF5Uc9YPJs9pUJKWAtC4qXh+mHzeIsM48MGYadZQ9xJmkzHpfzmRIi2hsCGXEGewa/8miWsIHI4H
CBiYAb6zSV6Y4P13AFn/uzINhmWkq1GE4k6QLMh/oJHQlOn8m0ysZ/QTyvSR7Q8Opba3BG6W92xT
MHxJCu5qEEJCRc5Ghcs54V6bxKNEo80ZKPv1YQQWfUsYu9OEj/8jq30JokMLVsGBtXz50/D51Nsr
oReg/Nz90ImZFzhtrdXy2xSYn9V616qfGnvgnBQzTZeKxJNs8o4dy+h6SPHfhgeYEQzmqRdAiWui
KIb9Jocw1OU0H2Owje7PhO8tqp4EQTrXH47z3weKqBJDiBUGAt5ORaKyNM3MzTDnfxnLSzZjsOnk
6YdXuGwt/oy8UaFYmGdWSuwuA+3SXiZLa3KDINtWXbpiv94Ji6WJyz9jo0oZ44XPtGDzc8EELiuY
mFohJRLM9FmEG9xwOvAu4pqKzTSgddmn13VFFT7wc6vdEW3/dLFGXpmmW8FRvADe5uaNJst3zuim
ZrbQmOHnAlHDzlH7r8wzrKKnvCVJyW+AnyMVRU92WCUNdaTjM1xKI7ZZg3PsJ+RJJu9NHZsCFpU4
kvHafo6QMF2jaFbrW9IlgbAt7sfZVhM1mG6LGXCOoipflgrSt1i78+4EneluN5ViB8dB4N8gFKpr
ZPYbcPEzDqlkfBY2nFb5aeoEZp8jqiFNZRjg/wDpm1FnT24FTDfcF3uGcxp9HMo+3WF2AApVpU77
NuK7yNwXxodTdMmwnuAHixO2C4f5ka0zNbgava4+XvkTKiHqRfMvne7RQOfZcRYZTHtFtxIDGuWQ
wg6VK393EwcEYdU3oHBkCJ5/4k0duS+396/GzS19P0JzETCObB4vwktYARvduEvwiTAsiaCRRdgk
prAozh/32EpjCUGdJpqzEMC1jKJOKj6ECdiEQogMv35TmQoMpV3jJuZZG16Lznv7JOWdaB7jvMg8
k96T0lPltS38JjyYAlWNC6oGZBgCa5xTMn/4mksqZ4SvRAiXhG+mqAAdMuMUbR3JX6KxarlP07st
sJi32DxSaXVAHnmmlQwIQ/bxOMWwy6XyKbLlstLNbFo1Kq1/YHYiUmKsAQeACrsLZohnmw/S+gg2
p7H4EmIXwXSaVdAFPp4/DU1Oo9tEG1MQORI/2zW9k3Ksg/YBKypy+8hI33bXiK7crEAtcIk964Ew
ZCvGwLnmljGbJFWkYfOcdCi8ftvjo/zg8k2cTD0kaeqw9xNVyQyET/WIDf/KBUmkotFQESOLH2nA
MS63BySq4RxMpbYudjUt2pNFZ3Tdt47Qbv+f0C+nyvGTH34y1BgFfTHF8EXg7qJCFD93TCOBtJ6Q
d0RNj+fneJzaPGZWuRO3i9bRyq33NubYLlhmSG7TlZQ4jCom6bSxDy98TDdzZ3XTOpkoJrhabTqa
/3zwirrIi64fDOqKk0Cdrgjo7noYhP6Z9K5kpo7Ls552wWg9QZK6NpNy9WLKUuhaBDcHP/kWjhzM
20VgLrmONK5Jw1ziztGfstH3JJ5jXssXoPy1NKQAAiwbMZLjVugisXXpJSafzmUrrTY4uR/lz1tf
TvQwOoO1PhHOhrgITVsfxS7Pw/YmhJ25B5w4nZ+skLI2L+W3gaTWIrQRVyohFRZuG7R4yaHf0dbR
l7gNCUSwzWsRAWANWfuzd1tQQC+VDs9x5/KG75RipnoIc0W9MoP0c29WKIvcTFtMP2zpRm64wz7f
Flf20Kn/HjAo6WyiVY5ZqHYEES9LZL8/I5XR8ZX3PAMc3EJnTfshMjNTs6c+eeFfD8YX3KwO9Xb1
035qZIW0Ve903hjPviEG5Nrqabi1foHAgEWKcqaWNTUcopS1JWXRM8fheamCmU/G9lBkr1yHXp1M
wmjBmxkzRMCGl3jFhMcXkTkOOn28x8USP2SDSb9UmBRFGMy8T9H2JGByh8b7/3FyXrPmQcD4qylV
BCBNFDMlSM7dGMxBuOA8KP4ictjuPHnZYtDqhRBQ+n8wVYz0AY45M7OI6YMJf0vo8N54xac4Zgf2
net+IgpyKA5jOMiUE1dmjhz+JdCqcfkN5FlP/pQGq5jWt93dTtk5B4wDO7VhsQ5o/4u3Xg7v3E9j
Js0wlCwAL+FR8VEUphQajMqDvCRfNTpOBnY5LshvmdrfBg6whl5z7v2tT92lsxLs5n1wANH+9XEG
KFQ7TLtJWPxE/CfB/esnlSimuev2k3YjX8h460F6gVMtyDRCePQcGM3e/m3yvm8xX0+VpLXTC7AW
hXtM3SFBnnJyajtuaT5ewtMCgUX8Me+log02Fd0u6+5O0YOx1X3DTld0cOHYDfqUWOXZugJnCdft
mXGlOgiBdnOsEBnLQkIHMfk1QBhqYg9CDPOuAl0AWE1zF2EVSCnSDf0+TUMtQPz6Uk+gxAeu9FO7
YOmF2Y5eAtLj5w9XCK9eXwHOGUc/bZLdiZ3/5zoIsOxwXkrxz8VR7tTn5UQzFruaqWOn5IWpQxct
RdvMvSuiaurkRzRR5hwHN3fSJy0xYxpemDlU+vOlBRI0zHPqTSEeQrC34fPW4hd8u3I8etDtL082
nqg9tqoEi1vwjoq+6ntXpmtN0BSnQk/VWxwITs/N3/C5RUuabdOBv6wsO4dOTVPCvl+bpKziV0pM
ZM3j59Hgceael+HOm3YFBHhsx5KQdGlxw8tJkX+5AskfatEnj+Pr2CLWe29V1mkUU0dBkYOUx6d+
dROB7sDhj6Goaey4Vf5ZLtug6baL8tZhd1FYN1Wu4g61X/F0BoJLW/0cFVZjreKjWWT1UPpNgjs6
3b50arZQebKgO4uWxA5zqbCjPgo6eAzEKjNupQYcvB4/FNfkIx+715QN2q56LOqCkTaIKuFdswS9
xv3877sbhO6eg/HQH295ETcyD9jazv2zdz5vQu3DMQLPJ1KwL+fU9tO7FmtPRHO7R9inPPVe67yQ
Y28XTMHgGCHxgYHyLVXgmZgpd65XU9KG5g1OU5m26Ibskoztp1COriQ/h4aK/MbCbJJ2GzfiLWBe
mkeTQn/UJSnClGiqMM/0rOVGLXHPPQGc1y3DoI45KgOZvYJBm0fWaQrBs8eI8SaWJ8Bum2lXRaas
MVPvzcIcxtyiusYKnAQme1ZansvW9i8o2DP1OJquZlWU0R8p4cqwUa5ffF97VSWG93WspjyS0fot
Ia3ExwhDPa91+3/w6Q71nTHz34cqD/1wBklMCBwd8nkUNHyF+WosT0JPSK7SP1Pu0B9fpQ4JhY39
uULCtgbOI+KzwphAqAD+EIcq1et6TA1fTg+OB5lkJI8PrRJlBZSf+4UrR+EqhQx8Ua3dDszzKj9S
MiKFjJYnbr7EYADFjhZd0Q6tWRjQr5y2ngenO+6Trq4lSW10/8b7rOCYOWBYis1SqX6EkmdoihjT
wk0RssIzki59Kk+z6/iloYn7jllz6vYqxd1w5nqbiueNwkMAtfeNqt98gTu0nvzNfEpOSnby57QT
7nAKNAjLNRuT09PJL2/767YpL44IgcQEo5D1M8vV06jupiqAluwSuohdaWB13C0t1sWZ6d0cj1tD
P8vMP6ectC1f6nvrEW6U/W1PvpVYqqcuGn5XOuFK3M49MHKCcnXE3VivO5vM8IoQTGzTbO2kIG53
IlxepathjW6b2YP9msGdeaVuTtjLzrrLe33ciNDOkvTQ61rERGyZ3yY36cTbylEJgviWKGHroSKt
PLlMbMnuiqgN0eUgYASA/IfO6owPs6zmCagOPp3tDhDnRITJyKGbiwVvKQCqQUU4UIJ6a/izAYT2
y8Dp7qEtl52D9igWljNeskKKMvrcHNPuwuqo0p2anV+2NqWlyqrGm0ZQ423Ihelub27XmwDrWFuD
lbde9jC0J3Mmh7lEbhKvLOfJsFU0H7cotJ11ZiOI6R+hKPPoePOPki7qNe0m/bjgtyKPpr1RqVtN
7k2l6M1tmhK9EQBhcvLLaFG1KRU0IPLnVe+8S+MDBgS4bd2wrvI4FSKAMt50oOmk0NE6YB6hnIy0
DDh5MbG+nc6+FDu7RKbtx1ktTHFNICwIP8UOLGsC2bDIK5fcWUl3IoXBL3+oIwP5crXHMHKyQT6Q
KEvSnKxdaOiiYerJaEe8RnxpIVZqR8Upy3mmbSMm7QbS3HlizvJmr+rMHMerko5hPwuud0XYOs6K
00RgNo27PzHqsvPRPvtfDgPdpQwVLf/N8Z7/GykW+osLC/1AAC58g1B7HA8S+iKQ6GDZywVJMpaT
2HxpiZLB486x49Ayazk/Xd31wxEMU2pghZNftofBBeWrZAlxZFbt3VMzZKBRsH+571ts70IHSocP
foRsnS4mAakTryxxYgdR5f83YPfoSl7gugEGi2CVjwUtxQvaab6vwuyojvtGp/jQWDEB4+zkEmp0
Ja4SSVpkORDxhE6EJ2vhYetIDvrg3RYJzyrlITh8oy2GvyrOUqYIwo23LhLh/okpVTwX4W3pXOnu
8z60iRdu1b9E1tBuY16S1VTKDTp1iRmosbKAuw85kfX+yJrIwHSdpisbPnIA0co9apoloK29631s
bQT0fksflL3CTqGfgXr6ah3mKuqCxQS4s24M/bYLEh54PMOv1EEq9qwpwqzDRn7f+BjLt0JtQB//
y2aQGGxG+eRxyw5TAXX9ZpatpN+PVufhQTU013MfGLNp8cUNFXrbqLQKSdUL4FH7cSBnPY3nK2Ug
r6ErHE0G6ITxSlbyDWgm83tAV8/sZYZ40hISm9L49Hyy1+0mrkya4e0m38JG+xas1hlFKjJw5SJx
7im+XHyG59HXLImtPUAueLr27x3EcZ6/ku4GG9zbrnY7lLKnYMtxjljF0nkQOHOIbU2IVzJIrOqG
u38+TImDkjyS6wKSBsHGMIcOnJO5JT0oCIOfKzwmR8dJoODyq72AZdZ6SouaV8+lzPYLZi9hvEdQ
pn6sIRQnf3wCOrDfY26+lzylSnC9F0WzmZHKGtOn0gSKgDizhz9aAi5+dZrFG8iThm8j9jCRInV2
nuJ+DtBIkqvGeVtXvvV8uqiS4rMLrhJiG1gvUSGwGiAKRx5DNS1VX6jgMaGHMVlZSOyKvvxi3er0
Vtd7DVsTLaMeWnIG2joQK1yu4OJNAyIJwcMeeSyIUFNC0c9kFMonBbC8I9ZxvosTMCfZmG8jePWz
pXImMumRxakQKD9vCOHvSPNgx34mY2FmzoN/KN47n8QBE/XFa6t7+0ZIENuUTZ5VsBcLH1VzCfP/
wKHYMZjikkm81Ubc69ENUYyx/NHAulZu4sBoA2NuibwheVM5mdFqSdJ4GIgrwjozrEQEcvKwbrCH
Dr6uxA2iFvx70dV683tWuSvNOpYiYj/YNL4LY4LPTxBvwRjDwLlV6CuVHzXN3+BygyqiiHey/oQA
Z3Ew/Ubr2HkkE6qfXXbRTfC54vrkMSuaGwFTfy0k/IwuDvcj2XoY9ksT0jdtCCAbOnc/QpU04iup
z4Rj57DuD6tla7xb0ZuDgY+utLwwLEuNB8I+vA1MtyXq4jkSs4B6xnjCntyjSoTAb8IteL54xXws
yS3fZWzadqO2o1peapkEvgBBHN+l69rJoizogWnh4FSX3TtMAoSWFxSgyne1CAX6+ZRuDORTBSsM
Uu6NFar3JxZF96LcmHAzAMkWVLvcjdC6lSn6R5CB1oIdgOOz7t+2jgFREMRSFl7EXFbcN5Nr/R4s
uou2HibBIP+DIDbjbRyNZgM7o6Y+i4Ap9l7Dsts0VMKpY+5Gm16qyEIIvxWUR6D/3Ks4tLSni9Xc
1z6vBnNmEfKzWPtj7ka17tDQVpzQBXZnPrQvH7Z9cHnZaCDFLEzmNiigXefcjUbOWLbBgsEk7Rar
SH5koqQAC1b/gQOg4UxO9iG4xOjnpzNGR/GTbji2qQ0Vc/6O19hY03c6hSRTrR6NW+H8RtDqFj1h
+8K2P7TG3U4HfXROfbBKE18akma2LDradFt51WAwOOsbrfCRd5pNEQMt2+OjMLgViArEhtwOy9st
zuxbkspaC5w1HBxSsj2n375glNKAXkrSRFE2eszbLsoX6540iibBt37NKke6xIwN4lWZzPUQlfcd
4JZB+nQoub0FGGBQe8grPPsynoKUNOzNSHfTlsE/EHGqagrMlDtXUTiVtnUvnUbxnA8kyWhanppI
MVqdO+mO/dGgg/U0OGx6UxbwKBbmALSa6Ig4eqwaq7U8pOOMgCrnSI9m/SEHAUeSr2YSqk9z7qU7
N/dEkEHCrh4c9tsBQuiPyYHN8a8i5iymJkJBW1+k2zecNVyCkaB9uI7N0JE0zYiOpT4jcau2tfYm
3PBTaeexrEuaoCGMFhlEGgb+syAZQ1NjJGjeqd98hV3MzsDDVd8Ow87YHBsTRd7KNZ+86fxP/wBo
XVbGNz0RkmRAkQ4E/lK2RJ5sJgYxzVvQDGU5UorxDBy70Qv5VlmCZ2BE0Wry2ALhrXdVeAN3JQGC
VCBDnuktXHvlDENinySkZ/A1IYd9/zY3jiLdviFiIGCNcyn9Qa2ZCJeyGdeywrgA8SFDirnW6BIh
q3PC63uEdzT//6hTul/w52vMDzKylHziUe8eLz+9Sg+Rf4N8+KAkzCfeWROCx53i9O5dTOnTlrod
6trspczFsERxmyggF0mK9miAWkYkQ8rEkNhICypmGFED5bAtuvRJQmeDGKVt8Jwku+A9iyLxEFz3
qtxmPKow0vn563TRz6MZZuhbvLhpuNnk3jwdReSDPjwZs4B+FQp+MwHkLxUeqKQF65g4cl2czTvu
tItWqC6HUnQrUueMERHfc0GwW+vP71V8D4u7vBjkQB9NGNPDis2ZrDwanwobWprlSWSOeOArXVSK
PuHaA3foGQS83DxLmc7OU5iXLtd8D/nkhWCsd662XysmDRdXfBhu3THmxUbZuV0dv2m7I9QwzG/L
/47kgBE1HgmY5InwGgzuQsvE4RmsMauaxitCq5gRyptMoW1YyzDgh8TDJTFGfD3Koi4Me6VDqeUs
VJ2jFgw9HGpRKQa9Vimh2KqsoKw46ZR/7J+sPAc9B1VIDRD3LHMtuWPtEa7p17J77F53RngxNC8v
v31C3oCKXWNY1STIQX4kpWXFk/4i1E5sTXJNnNTYEBd+h2+VjIhzTL4kJAkbirZDjJnpGBJpMGRq
RMHGZ9rOAfs0wiMlLRI2sWZ3BDaytTIN3Tw3lOJQIP8ozedriBr4at3U3T6vEGyUIeObZMLE9Y2w
+VgTEtJ+bt3S6uyw0bky02C0nrRjTzPRxf5km5HRLF3ixScCUSuryvkPwg0WXtHG0RaXNZHz4TzN
k4StsZYtB0nA+zVSZYtZT6Lrz7vY0MPStMLls/kO1XlVU0kHDGyEAVeCDnJSH6qtgpTgTV1hctGF
nIZ7B/wvlhGDHN4hOLFmJpjjbASfW9x6miQdEtaIvg1tKSOY4DlmgyHS/wQn2T1czo68SOjO3cOe
+UDR7fZzL2+S9PeIpoEocd4G49KL3R7dA0ZZwQ9ngMJDZXaZbvsoJ4EMTD9sRt5FiZnzm5wOqeo5
ZAi1dmo/B6VUPZi1MbSzAAUzRVlu8o1zLxpzCTYGGUu6MwijqeW/kKwG1XC+vDi9RYK7rt6ZJ6eX
xC+grl40cJaLRmk1arVJU8hrIybQpwh/lyzEN703iB5K3V4NJO62MRlq8MZbrDONyLmiqRbxh3sK
YKfp+e2GIVpd208CD6bjew/tQxB70LgJ8WLugEj56s0ECP+u4LxfnZyeAZub/PnFIKexxgWm8aJt
CMYrLcB5deG9jwUaff/TD6arnhqM+naY7ihJ4do7rqhQNMo0p2NNFkAPCs3dc5JQ9DVNiUdMzhDS
H/M++orC/t28ECEPHPZsKbccsMOZVkaj8LtTQeFBEHlqZ21Bd7/WDA3oVuE5yhofpK8h3F/ud4BG
XsBfqHxlQPV1UnDV3spEQoj5ZhzGNUptW8pnwxQKPSRJZgDo65FDNEhITd65NSZ9nv7qybMX/aO4
yav1CdhcjGb/AUV3alBQ9trrnI8y8XWuTsRBKtRdAr57XSqhxiDXSRtr05mLxSrMZl2So6CKHCrE
t2hALo5WMopPZ4kNgCPBmvtDP9xSUhCCDyhs2ouOI183YecON2ofkf+JGwBCsLIu1zfZgdSrqQUO
juGPg+CYG6+7GDM7BKBf7aIi4GHSd0cOGeuK7ZmKbQnPHpk3qv24YKG6qzWdCEd9+JyGPzcJYk5Y
yIqfO0KGIUzTgLKk2Z/6UeQxh3BQh4NTz10ISKH5HxHV7YPepjmutNZUwtXrDgqpxs80/AffPgsD
8YGE5JbUt0QUQXa5QtblOz0sQxZqov//oUG/a5xTXV2neY7Sktbk5G0neSzEvyJSSglliWIfZ74n
AIWGlTrBzC3ezbtKyY885o5Es90uoPvkZfQTONU30VF7/fG4Jz1krqwBAONY3Y+Znu/DWQwT/qGD
2rWyBJn7G+Ib1JBa6dpDHYiW3GA+6D37aNXNPnTeOP6aqbjD+QMMr0cQepb6AxCNC2DqUCYBxSrq
vyhZn+N5z5Cq8TTPLV+HjL28meT5uQ0xtE/FYzpHjrc2OwJHTmoa9LiVz8NrX0SjWkg9rFGEAuEv
1h6xVRPog4hTJ0DB+qbS5V3j8+2MFOMT4Lzcd4mz4awHqG1eNjazdQZ+r726q+eigH7egDy2y+hg
bQ45Ik32tUZv/knkMp9ILAvTnZNKJTl9EkVG2cxTmlcmBtaCrlZJruSSUl80WtNFc5ZNqrERxQIS
3/Xd8In1o+RrvnH6E8VhO7eLzAx+Imf8o6JdI91WgU+/68ZkJj4nifg2rtg0FtE5BccrVFLRBul2
9JWegO+hzUtHdCrjrzkv9JrCwfKrUMfzpgmfka+Rb6riSffyvGdhL7+aB3yc9YFPft7e5fMpIJIf
1yWU/iY1rGfgEOjOKN0/7Gx0mhxJiGFLLNF0iTyrSOfJstJGMOGQFcR17hPuNl0CyS+R3KmoOurO
S9hvS6P36zDToo4QihTdBnyt1tfOV7rQKzikZKuNSgg1JYS2q505vRDoirbkO5KOqcvZt8KM99pW
lhdLPeoxyqSRnGYR3+kjL/RTK5EAKXV/IztDTYcwNzlodn+hgmLsjl8aPD48u7uiNz5b9OHkpw9x
wjstfmmRxnOuZiT/s9ti5mde4l9BNedygcKYPR5M6Fk/V5ZZ0cW59rGmk9iL6Ch9KhvkJRhKq7GK
mlzqnQ5UTkJCnYU3FCE4BMznINOGVR+xT6862MUSH4GJYG66wXv4tvSzm2C50FLaEHexkkWykKed
5l46fq6HHZkxWVDEA1sJA8k9wB91tUDqYUkwQaVSFoawIiwitOjRI/SXSGCRYEzryDavmnW9BaTO
rNhU0IVj1GhfhpyUWM55N1s4pIxI2+UjM6QbGFhEnrre4caDx5RxYsilR9RvaGV4rM2qFaME4FMl
75KARkp9Ag+Vqh77hFTOe/ewaOi0IgfuLbm+wYWzcMa+yuu6GCpL0olfcKcS8aPOs6xF+mYsiCA6
mWIZqbtcl56jijqYUWNVrBQ41L94hh8W+TT7GeNi4VvSPfT+mqqCgTZ3LFpMzzp4S7AwOyUgESKZ
sqMcwx2zUtWakibeYxDEhRdMTTRSFlLtMLOrIBGSr2TpgUJX7MdkTpLdmzICa+Ii3XhwU7ECXwik
4omE6vPrbewnz+fwVGPgiufiCLT5M3CK7zuJP8sBPLum9+eX8nkAQ4fhWXpgDkvrxPxXOE0dTeTZ
cIQ/rIg8NCT3LC8QnxhO6RL/pB0tIwUEjZ0mp74/3pZEeXzR7/M5Xl++QhENkefCYJMKpaeqdJ6H
+39IFrPshpfC14PBLsapPGOkiwq/hH1M0z2BPaM3RRdQwbA7aa6ELOtiq0wL0eoXUZx3w8fDqHxP
cUyeUnuYnrdVWwHxb3Zi/nslvnpb5b5I66eTVbtqIsjr9afnyGLxg4yoTobE7lO0hMzXBC/gG1iK
+AUoPyolBW2jOkdMsx9wMtKoUxKRwzlHe/8kjYPjWOu4qjDR/y0YAeXaDRZYhu7IO+VZzRu6zA4I
bAOsfo4Mb9zp9Bi7qX3bbge353x8DIXfswjEQq+gj+y70APR0xl2dTrjmQRyjDXf01NRovuYPKJ+
5tRNvDPbbi1YH9h0y3PhBvL5luDOzZ58l7bZsJauRYHwi6bwIpHPNRwx82vLalovg+X4t7tVNoxO
BhLZ/narjKudfhrItEwolo9ryheW3ssZJUXvNk1+W7nfLXNmIElcSA4aXu7QYKCK63/2JnBAKCkZ
xL6IMb2MCPayQhR/B4yLhy1PjdKXr+jMqHBQCkVYWk2hZdsJEuA5A1m4t1azpZDJ1b1cU1r2Qunw
W+LWiutPV/CZKU1X3+SQz69iSg0MzK2uiLEDzPPt1KuQGEbx+bCjfIfxzngTRHx/1bxgmXhbxvMy
EQW8DC+lGtv5j7lk1GUmcm15aB3+UkH5vfaFI7yO5FjPx6YXt+jTU32yVfcDcjvr129uleH3I49K
brAAaxaMqbm84EshSArLx56yZirZqbBL74Sl2u/RwsJ8IpPsd7g9prvhvmbswi3Ue1Dom9mf1DNr
xkXX0r3fLn23zSVj/5NENhWkSq7VqDTQP17Y9/wjHgq8fgr05LZPOGHmsaEycZzI9AktPkj/YOzK
Fdu4k0k3x4+BVQL6PziFf8V6PmppE1ttfPJEj2qXSQthsOsRR5Tu5Hs4K0Zgzdf73Bah9Bhx/rDa
d+PCxynL7H85bodV8Onf5thgVGkESIw78zhh4WaamTj4qzfJeKJRg9olGsfddVWAQWiPaJYQ+Ybk
vCbZ1Uv7eUxxqd8xhhV+axQ71thc6Lzpu4GCzfLnEPkCiEcdgxtrooP5K37VekzfsjlypnoYcnfB
rc36RzFmjbPNwpHdoTeayS9hQSqMdGiV72t8pWxobSFVZ9MkcK2m1WtLSjIdMiYLyeQ8QsjZvZhO
KaRGDlnWrSjCE35IJ55Wjn/0lVCahqtIM/AYugmDMxwRt17HzekrsYya+ysk5gjFOiBoDnhD9wcC
BSXzxtgiHtWiiFcJcrLQr3SziotZMGuVaOiWuwd9YCe8n30BNWG11RRJ9MH6s7qLZk1ujXrhTPVH
uG4ydaBECkzA7PaRtcB0IlWYsEJ4PVdGGGCb+czvHsgJzH3/Vilp8j0WPe+povm5JwB2beNbEciG
nft1NRhoCwUZsZedxOV3iLnbebD5LmkEzKb8Uzo0aPw0CxRrgmI56xvFyyIjrveQzqO1BAH02olY
hfLWWMRJo/uS93q9Rvc0oifmXdF2VZe6U7dA12vCmHBQc94Q6dOTN/F3k2lGQTEKSv5H5wX5sHtW
/qwfoOQckx0bmFcIVEJ/n6DBYca3Wcj4dAROfRflZr0PIZKcxeqS71RPfKldtOX/Ef6MyxawS9Js
Wh9ILTlokzygBfBJxx56L+mwEIxqUm2W0WePfJ35XNn9mCKsOq5PO8jwChrBQTqzGv9ZvoSL77TI
5Tu2IoXYl48vqCUqLni5J2GOyjKMnprb2YAYDxkL5z0Ze4iQ/NPfF+WTh2vNVbGqNCdn5d7szJ5R
mwCTfu59k4EC4deuJI10jFhG7GNo4kIuB4AwRbeuQqa92Cn+T3DRQ65RIWNM+j7d5Z9RRGu0lg7K
Q/Le0VAbDNSxMRauUmOHv8p1F1g+P9G9vKzcB8Wj0WHGPpxp9QE1GyuA+15ssHTgfn9D3uds7TIE
KosuHrhqVYqz7dvO/SBoahRbIP2xz76F2EThZdKd8ZL56J60XtVozgiIb0ktRNURiopOpFxFF3e6
Kf38JFigfhuda5WJoyqvE/cE6X/Bbt5IGLsU5Y0wafk1A+dcBMwn2yLhMJNBREHmJ7SY924BgaIz
kCFPvzm5tgHCUyH3iCkSN8okN4FaY/fJ9abwLaEaVMbaQj4zCxqG1Ho1iUpzCOpdyvN3Bpy6LmUv
qkq7OwrwRq8QH6OPKmJOAfFdHKkd6Lam1sgHatusjXSFZgBhwBAac3qIP5eefHyKo6IY8TjOcr0N
CjZco+Y/LuoCeqLVed8EpxBImgKkBt9+GF4huCRtJK51WJn3z3JEzf/LYrMWCf5HpmW+CfDYPPRP
Cl2/jBlKri4/Q9LGdpqoYtaDM6OeMlCgm4KFCCPBEPCyZ2P3RWyZDhLWZFhSqUYgl0PEjEIZRSSe
9dtfMaYSgmyHoTRfWn9AnFierg/rieHj3nL5K6vY7fyEAab1Wovs8sRT2as1F3keYUJ2KSn25jxH
HHJ9YyBAh2+wCm/JD898+GdcSLBFHpdAB+WgobHEtTDZC6qKGQde91Sgd77l73Dc9ZB0VVmrCj63
R0b7hJY9LqYQyann3dbqoOCHJ6q4Wp5Ziddb75fcyWmutTNh9pAu2fpNZXP4jTkcKtuKdxpADN0F
yDMfa2EfnC1lE1T9HqIDj0jKtDIIlaG2ZqhITN/xPF8+FQtbEM50sb//20RqK+rCm+lucHQV1tA6
jHXjZ59j8iOLU3pVvnLIulQ5lj7C8CXtnSHSuxUNYWq2laWR1u2zKowbKp0hX20nYRsXS80tENQW
7bX2Pt6lQZF40rHNwJy4m5kv0RffoKLNUJJy3NvoRDRu4NZxnY+nTQF7v9VuYkJj0mzxIBkaKno4
txBJB3goXKGgs8Bp4cOJbTxe4qMSh/piRuGMl/snxRSM/EgzXP7V2Bln4Mdc9tD5d2C4z8A4eejR
lPTw7XtONF8m5Jfc1LrDGHn6bSmXEbcpn8UsZgZImLJ/gJIQ4wVvgfqAJm8lReIFSYdL9dmgQ4tl
i1dIjAPcNDleFTp5xyog4r+9oyj/RUxEs7u+Zsen7NL2/1LaJKxWU9zPyAqpN5pD8BQYiooLcXyt
NKv58iriVAcXrnSZ37h4vvx5xxm6Xxeq6pV/b7V6a6q1URr92pn0LZVczNapGmb1PMF/1IQ62nmx
IYYDd17znf9eA2sAOwWnAreHjwrzammLvIc1HWtqX6Kb0vzIGZiBfUxu9FFbjzrfA9tGeqQ6GWTU
XW6M4Q5ViY1CbFJXz56gTRleh8Sx/VDhw/wBR3js5X8b5v44+2LECLV3xe9QAW7421tQhXqZ6bis
z9WBAb6s9+gCUjq8y12G1sIdeCXjo+hhmxFfoF9u0OnXvM9XcKFiNnJegOP8qWuuzNxLmT3JbAfq
HjsORcsKZFR4qCNb8n+KZk9f2AJMtJDwDBGQRn5NXZ2lm8FMpiSEOx0aPDGpfni+KkMqNOhV9yTy
zknExKRJJx+lfBVijIFeuQ/ReEhlb/OHulhAvKw/Kv0QpMd+Mv5OO6ygT40h+D8FThWo2i/Z2PDT
9VQfCo+vVvU9fSzTKQkt1VLNNaQw4PvoxYhUTucP9wC5U89BNUmEZewpuTKf10i59qs1kFS6fkFJ
iz47gGaeuR5dfK9+hrLIOrwaUwscy6Ps8zVWxO3tbdxtf+8QjUKtI70ATvlH3tZeQbnM6jYuA/kR
f6vzXuctCni6/Ws/2LtD+GRZkUDSADhXESsCeKUsuTeVV8Hf0RhUYnP5bZj7o6mr7H1Xk69LaKFy
8m6ysdMnICFSVfvbcudXxdHBiJZWN+2PJzVlVqaINa78z92rCu7zzw8BuL7qULpcLdIdfWzRrFpY
a+wruza4ZrVQ3IDeZUjEp5Jpq4GPgX056uvGUePMyLBnIqvNlo6/IKztfC2VR7bPWNxvILV4bbwB
TrfOVuRnKsbojCBmmjV3LkdHxWFgMxo3lyfvIJlhEVGDpE+tdfmAEA4TcykKQiW5KDfItFJpVoxJ
NAudVNyoPNcpPnd2I9asBI6YkLqSrwR9HHMdGXlIEs7uTHzWVxOCmbSYwx0WySaZWjSpRQ2ad+VG
y7yHQmQxGSWdVguaZBXpOooaHFaLWTBw8ofG5fWk5DaKBiQ1QT64zfKWTTuZvDED9NJ/aEtwTHGC
ZhEUsX7zaatdNwNrs3Xh7oWgEdskxiJvPcmcV5X6pjhmZTXMJIH/0PzllTO9tXCOqBa58DWZnnw+
xBvzkL2aGyUuctgmXphRxogJjjs+FM8n62Xfk+7w3XaeNC+oBkVYm+l1/QoOFhDN3wLJmD4oONFY
1Gz1ShJIZBVeBfAX3gYiHG1ZekoxXchrk3iUeu6BS/gjI4KI2pWx93XYeAdrlXynRQVfYy2Tpzut
G0rVZqrkSemxshSnWr9TvS/xST6ojSEHvfaoSvhfkPhM9qZWjLsduvBEot3IaiuAYlPk5GxfUuwK
HL/tWkHNmIe1S187Z3K06Q6DLf1ter7xAZWhgMMSnbdY99x2sYQtSTyEGdrjW0V+ILDBO0MwfUmT
0+CqzGIMWU2Xi4ii8AeI3dpL0rPIxFSzxD/i7i0vk6zetbwvbTiHWMBf0QPhs/q+ejgyVzJlUNpS
8CgliBdly6Cesjy5u7iXqKgOBhDISD2EZrsCWp/6k+G1PevFLh0dXVic7ebLlbKK7Z9od+Sd93Zr
MzefUm3b/3GUV9BfcZTahWMiDeyK3741fyG/QUj5mDmOWnM78EjLCGfQcBjAuL40dYjTvZVbcFrP
3Ne7NRxPwGtQs0PYoq1JMzFthxn5Fu6WgmkbmlgcNm6csHrK+MTmiHi6KfI83kDBIYYKj4xIK+Na
YCMJ0crJU2Iqvs/AAtlIt2hr45Ti62t3VlUBMzRkOA1os+cixDj0oldnA4F4+k7C7ET2OSqG6Bda
75oKLDSPIv83jXPqZkNJC7jHhMc/MpR/2IZjd11BbMc7UYZgqwnZ7CuRBWVVC3QZ8ORkb8vG09pY
TundUM6yDlFnqTS3Y0F5y6cfdBMPD8x8WcCdALNUcHDKl/i3/EDQtyO8tKkn7vb+hQY60hmIQsTj
0TwF7qGqctrUF499PTMZtw2q31wdvMl56HoTz+5YGL8lo0aY1NBKW3mgk1M5Kcqb9M02Hnz+EIwz
jQ+jMDaN5Y1lTnFuLWaYaRHQ11RdC74kK4TXN3oIRoTkHzJ/0qE13f8UXq5hLzHfx+kHMGoA1k8c
CmWpBw3NAUxtJ/bcO3ttlpbXhZOu+sCQCXYEYScd2pUo/oH9bWQxekLCoUPSbV9WlQ4nd4icCihP
lXmUVhVhDQDp1xZKeeTQfVfiNqTKdxNIB7X+aMQSSfuOUlyOeYqC+4LoO5f4kJmwqUWfmhPAFxdb
a6L1NUL2kQZfJlx70J+q9dQ4YQ4/HWeBaPChn4Py74uMzaup+rKd1b5xtzPmdejDF8VZHLashfE7
dkuBXUeSiZRztDhB6Q24LOlfit/FnZZuoH2MpfLb1g1n6NROfjjauLNPNRA8suYFEB++MQXklJ9z
UNSGg36DH6Lpyt2sNg8OEDiVQkW9lzqhVE0nsSqqCZUR5b5/LUEn8Jd22Zu1+g0nfi8YmnNM83IN
WjQscuZmh7isnlv5WBmHRan5xdiMoFqXPYC/z1gS1EIpit7X5TAn1DjaWASRqP9PtfYkR1yllBOH
dq7MYTtV/kDAv6wxqq3yLfjdzzH5hG3OtPrKnGoxX2WJOHK7VtLaqdBNqfJ1mDium205eygMqkF5
0hc+8OEA1e8zvalyJPCvhD9cm5Qb3JTHuNl7aBrVeikhCEMSd+ZM+F0raOpAO1+ucCA1MR4h8Z+T
YLj7W4hUbzKD3rBQ9Pc4IBcKgW32BTxGVuqeNHr/7x6InASFTzHmCjqsV2LMGNhHRteZHr3O/GFk
3PIFFf+2uCxLH/H0DOp4xtltNqMpMNifZkO1DF2QZgKVeUOJLZttYrWBYDjieuEoX84b696nwXce
gv/YsHfQGUGafVALuwCQ3Ga9dBda6eOzGlVWt55QkB2hNCQgzgwu1oO9uJvwlH3fEWL0Y6WsAlLB
lh0FOoVYAbK1UKO9juO4tc6EXzhGTbhW7EkLgVrH8S1neftxRiSBfGH8keH2LqJsWDZpxcAxAvin
pzfpUubzfep83ycRyN8g0CW/B7wH42P+25CvT9nwzrS5z1ri+Fy6UPm8eLUlYyBhLEbpKlZoQDoO
DH/D36BhQs69ucyicKI/9ELxuBdWECVv7Krd+qT8Jy9+f1zxX6hELkV0VjXtdhdk8euVEo8fRLSu
1eq8GDAJVKUYYULDWux+3yeWu8MxFU+zJQHb5sP5+ZgdwU2YEMakTz+rlas8QXb2wpHza5kZs1dP
b5BlmygpgoZlGqcTFEKaNrw14MaMPzLFVla/S3FXz2/3JAqaiV0xLsUNPNN1m0YXMVoeqKehmUhy
7uSEOwZPsm9Y8JBowKDeYyjXm3S4UirepP8EeRi0QBYRb18VBIULPKdHJlSAUctlsGD/iFk/VGtn
je9gqSJEtNM59ObragJGnRQd92sZUpZgvNrdQY68DFPdoFp66cJAjBHclXe3/utz6VJEpHb8hSi6
fML5MeBFHIEshPbcU24vn7v6X+s+3BETTlz5ArNydvy8A8vfo/8Ql5sgtI2WKP/h8+WhOL3A8dOO
FGC68dWLneo+ZyKrRKJHvAmg3W114DYorUk2SO8gpWzm3EzseYvHhtvxv2asnHvsQCbgDWBVDIwM
/DAToYcUQCKwAd8sDZar5Kck5ZVo0gYHYdzJXje8Fpin0Yy7IHjCGuMT9RZuS0wdgdbHfIsNnC/V
vnCwWogE+PG+gmRTbW+5SnuBVuW0MZAlW596fW2Oo72PefTP10e28otBuHRr4n33yL1QkLkL2+dk
GYD4NooX0osBdCEh37ObeJVapentT/otgi16O5vA+KSK5bWM3QOxdtn4iQRJMLqI/CksRAlLxIE1
RbgX82ol66BOrmFNuXSYOFYKHpTCIxx79ni+jIrydXweHpcYSCuMOiIimw+AIE+zgLYmm48hDoQC
rCz332xB2crgoX+x9MCg3Lua89xqVIct7zz3WavUZLUbwZPinba1iRcoKlyhuYTAgW2SdE6jd5dL
L2T16hXWPYLoAExKIRzYCP4Kjw9mrdC4dzS1yswtuDcHcaS9iwIFb0G9Y0xxt39opOYz8dxH5Mhc
xn5xAftdWgSSpmcbRr21B9QFG3B/u0wuBfwSvvz22K8y3cFru1WkHWVXK/ABA1DGpstd1Wg7SGjt
ZI4lx7WnChGtC+TZldXDi22Jwj3YcE07AeDRg4xLTxyfC+m2r76cPmUj1N2gKCFp1Ggi1A1e7cAk
ZG/w81GHFRlVFOx4GAa5db90Y/seWf/STPiCVs1aPq6zxsYOk+XW3BQafZ97aIGhl4ykCXnMqHpG
8nL0VBuMVXth/DtdTJJgZpjdA3ypGpYn9jCz4U2U8SaqjNltMvrCuEUe3J8e3Y7yN4yeQIaR7aYI
vYdmKVP10r097NqIbW0Bi70377dG85WLFhWKaOMhFj0UvQf2dO493Fm3VdcX0HheZZcnBOccKIfL
EAQjYg+K1ArVbyyUmMO75+v0gHdvvzU3d1DbY7600ZN1FCl5vFiLc0bE94rKGbQPisEOADBx1m/6
tp9DGTvd+yXDTAwD5K15lLVAn8IMYdyz7/MQiN7dmoRm7HWUchwbLQiJlUItmbYNySbuLFhixIw8
UtwqyB7x+vloByhRK8Q3+iA1K2h/2UhZL49kqW7m81NO+LRzHSXhsbadrPLKMxCyqquev0LlLH31
wtYZcjCcwSjopYdW36tmN6+8sk0tix0nnIM/Wj8qvbsMGauipmIzzLhc6d6JBLr+VoO+J1LZFKxA
FWd4swuQPdjFD8JXeaMWX2ROJYnPKFCGrl/Cd43KcMzwHvdQ960s/A1NAx9DF3sA5aZDykJ4xUj8
gJsLpSXmvkOgTb3IRdiYLNLoi6mslIXhFQxVp1Dj+Kw7TcSRpPzq4umKLDfD7prmaAmNjjln1AcF
V+enT0S8YrYEPOc37vpNeOTaG2uRSrkNyMQ3NkBz2JCZDDmuxpkV7/wXIN6taTb3pxQc9CF5no/0
vrfuzteMF/T1jJYjczBam9+whBNHqlB9FdvV8eI8kQn0ZVI/QH+ddB99ZANCMRs8tHyE4Y4Kigr4
6Srpr55fNn6TrLj7yTLldXAKd8xbQtKADavPHOX0Ktrgxkae5bapVV0CNlJjXfcZ/+at2Y9Fqe1k
P6y2i7tNVWwZ8mFcAKwXMdUvkusEBzRCFpxSWdGTp8SfhoDQOYGn9crlcAVkNmcse9d+8EM+gMz2
mWGs4SKPpixB7anwr6ygDIZDm/N4lBjO8+3A92xBDE3Vqh+nZe4vfHyAMPXBpPMacKfgcfCTORiJ
jiCzQP8Mi6+LWuKSJi7uhOq399+yngFXAwREtvt1VREANR8cBgEvyrzXGOIlUNLOI5F2N9UqWtFj
ydZxrGABnOcT3l2B5baSoTMo3unLcIOr4b8zSrmlvUU7z9bKIytO4mE5E3MNpNSAymj8GhumKjdl
vEMziFyBn3K//jEeV/kHShEbIv72qt8N6+7celfj6v4gWAr4sj7385ePPQXbf2t3Q0wRaJ654H8d
qtnbr2FLogHr1s5w961Q+NOGc47haHysY57PnzjxomCvNvy40RoTCwQkcddUZjOGmxpTeDiC21dY
VH/Vo9PHSjgyPvKTGCdsjh8oT44zqK4Q/BAHoZbIbTnKJqDzxaUf6LTQPvV9pZYcBujQdkQNHYN/
MYgsmiz24XkHUPQaD2kZ/LHrZVZLyHMRuXBpEIa+4B/3e1AZJaz3/aeNp5bnNIX8PjAknnVtxitx
NlFmWzHdzVr17vSxwFRIoEYPO/g8l3+2jWfVFkjmDjlmw6fV3dpphyzavyPEvhxz1XLhwIX8wy8m
oouhPrARl7TIBu/5P+SRLxlYgFGfUmQcC0EsvpBR+C9qTZroNow5a/UwU29UMCey4DV5Ch/PTchZ
W+GVhr53ACe5W9GeB+QF9Cn8YJiJ1Hpy7VRKbRuW7hk0SRpRXiMvLG1BZGT4R2OZUxOa8STYI5v8
AeiYv/z2yv6mY+untZt84a2Cckeeqkd8HY9iXC1fcTGeYFSoSW6dGqSDixphPDJZf52VhkS/eFVE
pT2NHZDv+bZQxGoq+XNvJVx2xWwZ13Z5SS7mVMCZ7CIMtO1UPT7Z/ETMAVPFfeRXyJm0+B5dcGrc
TsO+0v7RN4xZRq+PGmkJ9OiuV2YGfHTeOjHHxEVb1ZJwucDG9XlVdENySWcnU0Xoqfid4zY24474
mxRkg5IyuGvmStPv5lCLvDgpKJI3AO0ZBkp9dgJ+0aNV+BFDpTFN28I3VrQD0Hpx47BbZ/9UaypX
aQrcCpFi3V31X+Dq41Ahjc/qrlVIBfAytCgxnHCwujaqAEvhagzYrjFaUQNwWkQ1GuXI9kEBxph9
O0aWVNKzb4mivy96Sy6vWmpluYHrjGzbZ/Z2yWpvyfZR6WDtozmMNrvlHpraakmScnP9q6aQb7DR
dbJdWy4infiiknGzEs8iZnSxeAQ+mGiudXLmPWL36dcUF9q6+zZEZrhwInxialmikkAxIuDWT90d
OgOknbA0S+tp1BNWgRz1TctK+ith4ycrkEPwYTxr0OC5ECPt4mCUk3HqY9nPHzaMc9LIQzmf0O6B
SLuRjNUwPb1XizHVGLjiZmDZ34qqG/6DK3FelUSWe/HIwjgvCXCSYdbTHtwhM8nbaWk9a0hVPXIk
iXyWo702ppsyNrRW/17XokdpgNyNSuMYV7mXCYoZe7UOzXG9h7RGafB5jQFDdNKocEnMsEHPjysg
3VNZ/PA/UG2G6R1/MKdBRD5MY0oUY/26qQ+zovWSSvOz9/BnQp2ju+sPicw5dV+BMsdDBKU3yoYX
wtsKUC2TfmM7sVHFWlCApu8wvF5l70WgaDE9vfnZapW9kQylxDvkQsd7afRrHZHe8tRaixl5EzEn
5ACTV6/txGYNcHJT/uExHhiTDr8wUji1EVtJJgTIJRIDiEyouhq/Wd7dRX5pexrnPhnxf0qnqrlG
r60XRKUBkJOogYpn5UyIVPM0YhwRV+loSu2Ntl78pI/ZTaHIxvmH71Rc9mWz0kO5S4+EIdUikDEM
Hi82h/Fw1RxQDddtj2r4wB3b3kWWNDII2/4/5OKrikN0jTQNNesE8pdjq/nIZxImT9s5/MaMjZ6i
kZyfXDyI9ARD9V+HM96AKIaaNGXd0uAvN5UwnlVuqBYGZBdySQupvBMys2APriO9BAFktmqj7Yco
fHnqH76BBinZMDs89ffu5X9l3g6HatshEhuBoJk5skgR/8XwQgB6K2makjEUOq2xPKofnLCYHmtu
7bIcBXxCFxmemFvq0AT9QB/hHgTDEJwiOF77OsymZxCAK0bMUQNbFPWb4N2pvbBFuRZrEtEbOeGD
MLPe55hCfmYxnSYwvGxw4LJ1/ghyBcgjj9m5XUR/2dppA6Deo/sMv14lFnV4Dej6RM42dt0c/UKA
uqWFqlvUdp1+iLqeb23Ig2m7/sH5BRVE4O2e/NMPlbIfKiHTRagQMRPUgrjDqQRIl1FDNmzbfxwA
sSyADq6/jPWa77WIkp34vmri4ANLd8kdHaTsX/Rjw3beudv3KqWmFLmiVNjphWyX3rpCRG1/PnEa
1iA4A9DbNpuJ1amJKoZVnMuh3r+VpurBSZXKg5738r1whI0Hc2fBi4plvGTV7KcrmAa8ZMCkZBYO
tSU1v/p60Dhcrh7L362cTaHu3o7uFxDgQ8oRPYAWct5aVPpGUi9j89ZvjS0/9twIoidqzb+XE8a7
4aQPkSZvajCcaC13gthSUmPDILrfRLkbGxKWiRfLMPSJeb2hBe6MHiHnJFSZSLMnROAfl+NMhJ8P
EG9yI9EHz3/Hffoa8RMGqACScvfn1SpWjAy81nDvmiApL5hKQN6kkevgU06pQyXxe/QrJio6jAeU
Z7F1fbJoIx0e3EK9R+6afKbeNg58k5AqI5ijpZN2HXbJLmVcy5BpDz5FDZVdL1zRP9FYVSGBqnmh
oVbVm/f1rn7z9PJZxBu9AzSKN0Cc3Hn1IZztAcuvYOalosMlTjJxImTKSFCFxV22BQ5HLfallObf
jLiWJbU40U0XAJm2fHudUg51y2b/IZshvTWvVjSeID3oCWZ1Lx7Pu/HrmgqJ7LVd9aR3Ws0LlFEd
eLn5bh3wUboaS43DpWT1jSIKNROTZwtlSwg2BhBaMh8vRBkop7CNRQi5K5F5nQDy0zVF0jzKuSDi
WbWP1hWcqMqTDKexc49xTq8X+UXollN/p7Vtk73+dWwkcJvFK1yZkpHwHpKeMxWH5SyOJJ7ZIvpS
SJaKQCOZsiJF8ED3Tw9/9wfe9ErPoFaKPu1Pho4Pq3zDDFUAPIoKhixvKZeHmnK1jPeB07TIoJZ8
vkuRS7t4tU9zAz24NI/7UpJFGbtGGp4DxX5qc/GKjLGyKETE+ixyyCTq/TVbawu1DBCrZ2p12xuF
zB2Zo41P5XennVPYN3lQnDx4LvBGxYn62Vbp5vJtT93Wn+yBzmv73gqLCUO4jLcbVU/rq0U4RbW/
lBzDC4xbSanLPVT3xqNOh9wffLYxuVOT+z/Nal08jXXGtOzO7+ZRO1YZbz9vdwy20CbGufpGuRQN
dKBJyroxTi8jTADqndzia7rpPri0J05W/uifrLcs7MHJvoFkHbH5bTdE5IDFGy9ZTNcAyRbo1oJa
0syoebQzhHT8QnuhF3bxPYWSvmFexqzQmWqexZb3El8a3tAK12A0D/g7V17JJiqfgYewyTBYvHDD
CL2q3pCOgFbEg5GgMOYcD6TciImH2arulpS3DTyU+I8NUO1fP+ktVkpq5N5IP/0e0WHE4CW+56jS
q8RZdnyrlzPTYRPWgDF9mdKadduoqcFeqBHxUGbFuXpYwUwcVS4adYN/PJIay6OBuYZykq4QsQO/
P8gFxCp05cuIs5QW32ghM08xvYEgVBkyAcChP5gqV9uPi6mL7H4sg8Wi5XRp3Zlqd1LgT1tXxXp2
7yIC2/7Jjdvg7omFDMHxYKmULARi8uVskxZzXLpJEoEle4x5D5LwDt5uG329Hb3DNDEQbhK6Dj1T
hmNnlzvSGktutuEpbvZ1vbWNB4KL3Yykr7koiLw9kpAhArzuV8yQGVu5VdBedcn/lX+GK33yGRPj
PJMOnKdaPQQV3yJzFyyYWYO5OsmIasR4EuM9wiBC1VSSShN7YiA7FKYbL+vJetmkISAwbJ0VWtnD
AxHmX7CkAYBspiw4xp19WZ66pNa3eLGl/D+Srk6lHW9koJ01ZHz450+xoYRjyDbe1L9qWet6n39m
BZ7SQPdekwdtILWMK0By9bbHVWn2azwb+Oavt1ZxwrFKo2+KJF29Zkxhq3P0quAE9B0WBZl8FmXP
cYjsWCwsWzBqXEBq7ANoD2zQLjbu47zjQ/nD4bdUVADCbHDZ6xG/83JGL+BvSsGfdAAtGm0nlDOX
8RjwjUDjqT8cZRSShCULqsjca9J8xzCaPgl5u58x7x8qgEZDNQ5jSp5yNn1oBH94pEYnhLYRTNKv
4TZyoAHDqJ7VamDkariKumhUB4seaJM157hj/msCRThFTo8RmLXKYrQAWRG4QaD9p0MLSpYJ2dub
ziZh58R+4VIkcvXRRFDOxJP2atmcyeM54ZuxEFXJtaqc7CvJ5G/WKpk8RKSWWXfHtzWMHsVCoorm
ZA6BqHWmo+N0jABY3pj2L042snGz/An5JSc86C7JU3FLrOWQj0G929+2/Hac4m+bQkfmhwK14n3r
3xTdXuZhE/5mr1GsUU7gQSXBTB3i2E8ckwsXam9VPxPEelnHzYbl6UMbYovLcBv5y4l12A1E70Wy
Q/uXo91hmyJ7jQMSjHT35Z4fxJmqw9XtMtlvQPeY1I5UL795dd3/ehlx7QI8TZXQds4PAHVHcSdq
wH3yYtxcpKjwv51R9RdgysOK8j4nSyYkNugyp68ae3N3l1vIWnGeY/Nm2ErvQ/ZDxh+2z9TZ/mNM
7Y8rdVzUB0NfK4+u3irmTOQBPeBqED7LV5qiv38VXVGmz/h6aqmnEpVeIv7ZZrB33rCljzkCdhrX
dFZUCU3V2xYn5Pr1TbYxiveahQFbVAVQArMHPSa6OwSmGiOvUWW1W4hv57narVKopNKtHlAk+olW
BrmAvGLjKWRGid23k1hd7dDUcnrFW6TfyZhhutndMOD4hTH/h3onArTv5Lm4CSsr0yMUvKpi4Msg
VIQXz9ocOfzTQek22UWBuDcMGHz2vQ+afeW6zu+Xs5q6GHuuRHXxjxW15b0eusaKNX09ElWnEavw
UUWkKkckFAYFoy6LiKytIsTEZJ7QMFUHqD8LXPYItiBSd8CC9wr7OwQZZbkXElDecldz0ev6Q20f
ezMGARkA88v1g9pPZvUVdPPjYFdxaRR/oupk1ZvslH0sOgSpdL7JlwjTDv0I4b6z7STmQYKm0WnQ
hW3hjLBitHzp5H/jbUW05fBLbYquxBs0DiVXkldcNMtJcT5i6bJdlxv7PplbjNQB5OablvwAlbUo
1wXHk8PUAOz1Mp8skqkgSVS16xDJR8vZ17dfyPlI0F8Av7J7zNKu/Km6rh1LAfwOrLnL2rR+xjFP
EB5hfuhR6Dis4aVUh4axH40vE8dybtH4TTa0imqaNDakbclBgNslOEZEP1IrfoxYjTSZQfHorP4b
HuKm7cRj+jSoRNzt6qWGm6WR/11rV9uvSNrG6879K4fUZiJoIhkFQQZDCzCfv5L/J8YJ2rQyyZ31
ulJ7NotwQ7izsaSGeisiKl5rNdbhHgKSqpCgfFP76zq9hqTobDhCi53wDKp/XMRRlRXonagircai
66AtK5wFOn2aSEf/BLG7IMHVD6TSiWV3h8FORvuFXCQxmb8vaFiLc+HjB+Er76215r/Ph0xycJtj
feV/LvDvkfwUAv9cThsPk5ta+1uGCxOcaXHJeIJ+LCfYKwt9jP5fxR6Mb9FIzKkonv7tODasEyC7
GG/7vdXel0sKbUpb/5oevrbfpAJvzN8zPlt2LxOy72xQgvNfrwRWrNPFMHKqWWloxI3KkSP+Jq/B
+D2yQXbbTbkCcfjzEUHVi/AJTczfZOttD6s/tAAfXIljzmv/H23gQSxu1rCe8pOu6QhqD/vSKdO6
GH8BnaC7EuBJKCIwpFjJXwHu1bwpJ1H/sg1QEmVl9/NyC/w1Cj0zsxA4IhxjKcRK/U5842m5AOYH
+JIfxFixTrRzYIjBT6ooNSugc7cjkm+7IlB4DYQMswhPqMlEbQr14yAL2c9k8FTwe62Ak17wB9kx
61+THP9UVAqyHg6RkT7nNAI0dC8jOWxBKF0nHer2KsS4hSYnm8S1euvZQzhtKHKFviEVyn6V29i5
VpXbUCdp2HsOs8OvoMZhH3tQ5gX7cH2xesr+hczYg7kDDcuI+LIaWXeRettKbnVPEC4l5Nswha+9
N7wyaK4o+rVCZNWMpYvwXcQlgytW5RTEagIlggHXobbO/ftyVbq6swC4SvahHEO010T8Y5ds/hHH
XMpuCVK0fOx8ldAymV5ip6xiyoKJSAI94KoulzY2r8TR8XspqoD8Qj1p/aPUFhvnugSNnJ2/FMQc
6gxSJ18GAcndTYpThqUynOVi12Ox3fMF2eRAhIAnbpDfzmp3g6dl6HFH8RKv8yZuDoWY1oWKEqYC
MZHEDTB+4hV0KfmOC7rhy0BgYTZowejtEHBba6wlwJ1SHcEZUHo/rvSR83kRn6FvIbz4HXLCaVVt
5EGpSBACy3vQz1eDTFOsgFGmY0ejm2yd7/iR1R0jb7008n8h4j/alsDEGgk/7xGsoh5pnGnOmwc+
AsReNqsS9RPdeFfK1z604P0Wbop5qrBqrM/Aqr1HHNt3bPF7vBvlDXzSeh4ngnZqx4qu+jNiRpQf
bkNNseiPnVDS3wx8Uap4FdSrg2HQ3bOihvVxGfIJA9MYqPfj6LQy/vWejLy86fbrOGfiUJPO4V3I
O1OKJFdepS6NMiTbsf79rQVwJdNWJw/IHtL1h5J23gonQAkLrlf01xNcPK3OkxRlmoPRDO9Ue/Ow
r5RfKWqrkIGSeEVEdygVMe3NMNI6e3cNdeCo8r0NgqyUJqpyTXNFXxwPb3E2CC/Qafv5dKNmm+ZP
WZNkhY1vBF30IyKxB8YlEo9HtpDqbc7PKANqacaBlRAk9zmt5dcj/xvwko8X6a7F7fZ30m+JVsql
fEfdv+wxbGyIvUAP3mMqwsXBmEX8YYtRtNHx30XKHLyul3lWCDzILnc8n/Q5nM8/4QQx/hm+pbFY
IVmi/Mv1GKT2I/jIJ1ZGWZgE9/0t1gXg94106bZIaHKi7uQOBJJ9peekrt3gyx/odK+OFHLDEwi2
vod7n6PyXd5wx7ynBGuWfUtY3HNRPq7zNQ4VrCl0tnAcUskACs/KeXozXHu18Q5JtGzvsmE9OiAE
FhG+Kc06iEO23Lt49eYe0S6AmTMlZSlXwYBYGX57ANJXgZ4CVRpAoJIcpPaLzjKZl6SwBZKmxN5S
M1MO5w4XGWk73I5dbBGh1TnY8uKqjQ4mmPliiRvlp5KGvyQE5kpv6BkemBR5v+G77SiWHCxR/CTA
sRt9o5/GcXI0FCUtgqyfPE8PNdUtgafzvIA0ydX/t02dbW4p9qPRRcb8FpQJGEXqU1hE/gRpLwo5
Rfjkj75x9ZtDq+wvO5lul2kTq+NnIHdO+G2av52e0GcIIHO1f/CPa8QP5PMc293gmpznlJp88T93
LWYa+qqzQFMGoFqMCyiRw2iGH6AoedXw4VRzT/PiihkdplSay88pVddFuH1NoKqEi5BehwZmpWSv
yNp/aBw9JhUHwPYM8TuP88by2YOEa3UlFZczAq00EBonBAlQU8KfnBaTFVZSRtu9z4lXoNUGgiur
IGea1elwQOMDXzNXwX/vM2mKFXDXs/aqruyrLpJhxSyH0pQMkEEfktuGcn/xuk+b4RDO8oaMHIxI
dcbWRVRMjQLTGz+vpbMygQJD+xEZrtyIZmmUbXkjXhnOM/gXVCqgdnvvwqxg7BCbBjeB4WajYFxr
zjqQuUx4f5vWq8VZXyI68zqy11szrmtuv/Uzx9SPP3LpiqCo3fEyCxOUkbDwdjNRnY46Dm1YYg6J
HUiH5ix0Xm4hBZ6LgrbHdKvvVGpG1Y18qvgdi55O0j8kLcvgFo9lFjN2Q6Wgj42GZzrsvJ6L5N7U
jQbEwv8Tl0Lad6XFa4TwynvlzWo1PQ6+GaB2haIPV6Fpw32l/xYxhDHrYM83Zdf6UdaxCP7R+Or5
6cPTdH2EDQYUOgQfnQQLc6jItN6zRAof2UyvKT+VFmtQ9edHJcxDExBvsnmZosrvn5IcHjhBe039
fasl9lIyliaYMYpACH0SXUjd5aAkraEXwSDKRKr6D+ULkCVaagWvNTlX7z1Mf8qSYxwUT0EdsIK+
636TYsGozI6Mo6yhZg7A2cCmoeo7v/qoo/Vtb8a8J+3nKdPfT52WtFarh4NWd22qghqLrRY2LMay
jr8B7iUJjh7kdrESB0Y0OKiohoLYPuqskx56Siop2mcUo+l4iaMdarAdCtDoNennGBxx8GuSjbOb
AMYhOvCGdfIfTrxGN91jXG0E+DJLb4FOhQKq/QqOgJagMCHG1QZIo6o6m3XyfwBXC+Lh+q8XEoXB
kgkdR9dT+Sxmk2v96OWp0wvyxhNhGNil4PHDlhPbdLMhLTfB5roLSPE7vBA/cTWqKAn7fCXCUC05
Qbasb/d1Dk5hpbU/MUcjIUEgZ4C1dz0XBkokLD7eBxBLsWZvGr7Jfj2FXPX7Xvb/fWDXRBs4DSdX
6Y0kHlPiog/tWQG8/8CvPmjoEcyXGhQ3ei/Ipa+k6kflI0g9DhSCLrWjnbWv5Xg1QAAhWI/KTAGS
6AVLa6HqNoQVrNJLBvEr1nh/LkS+b74qMuOPxxylOUOgj2p1MIxioN0kzEJVTcEdV+NCDIWqDccd
PqkVKKDwmBS0uVG9kw8ZNIQgW5iacYc9Fo20BuUu0UIP6lW3QvQlJohkU5BYdGW31boO3ktxUivj
s8jJ3874sdIUMmMszduxoNjTjzQI3Bh904mhYRdL1c4G/56bejzmV/CvGT9IteiDVXLRwVhiMKeX
koAEG5G8xgni2eOfXa3ym6pyuQzw1//AyBZRuM2p4/9ygmo51YCyiRHLqQeNhT9hlefJ8pAfyH38
c98i6CQpfLBjnBk67N6/3hbsR113xqNvBk/WQYP91Jdx0EIfHhIy6P67XKPHgtXSTIErKdlcD/bR
DwxV4kcR8E5Uu52tNMi8fNuntd027Ks9S+N/WFsjdxt9LdpEirJ6N/n+mJg+9dtalYHP6a1ZDwwx
EE/JtewKQ5mRHWxnzV0wkIH5i8AU2Jvi66TlzTbdC/7DLSNK7ziiiQ3eq1g9S3vxA85gF/z5oIxu
SEas2uE0NlE8XTqXkATSxiMpxqjC/jfHysHlKsHTBc934Tu2NvJy95MWpF1PQsRe/f4Y9LTpGHQ5
PNn0SY8xjQ7nXUE2GJIJ1/K3KHz1WlQBaFFEw1cWO08eXFFFTZcmRHsXjZ8WIYvjEzXhQ/N/dys/
xJbgzvmQFN15kXuoNUYl1QgXlaOIQhQPYs37RuJ1o2JGC+n9VviH+SI+5fUtZBccQNgQjl1eJX4v
Sfhm5lSxxFdf49qiVHpvL+eLHmBraF8Y+e7wgvzv48ztG82HKNKE24TuNZ4KlYUKuXk8RFdQycIJ
ekmwDOtn1HWfPwFbl+t5LebWrRT94hITalCEQUp+2Pos5N+aEFndHgdN8gX4of36jOTtUf4W3ZKE
hBSxZAtDBIIGaUctHTwWudpJgpIQe9qxpp5j1Zz1Bvu3Nx0M6jCtnUSY2XdGUfTvALfKmEKBKFrB
Ndl5oAuNLB8Tyz3p/GRm03n6Iv1Ip1M8Vg2Cxb1J7ogxbpd+ic2qTVNBgVvxXCeZ1910kJb6iijP
+2wB6iUdmvZAJ5AI6kdNTTm51H9rieEsW8kzGMK2UR5gw8uqdmpbuMIL50MvYSDALOX3I27kR99J
GycOtwwrXmgA0z6D42DJtifkni2azyx2ycVY47FRjYmV//a28NUpOilZxBTkvLtpEdaelpZCBtzT
VnznkuVByX+zyTl92OsjasNa06ujEQPBPINzjRavP6rVgssymfU9p3QFfEeDW8y2AeNcVX6zni4+
eswN4VM1zVSQMox47is8zmOq6Okz1b1Eg+KQP5VVTGXng4iWEdNwCHummudyvU8gAF72xpzWY5V6
mSsWRdV8r7YqQlqXhXgD+za8iF+1sIX8XpzF3ECSo3ewAG796EwE0x2qEGbrjhIiuPBLnLJmBf/R
FKX9Q6SmT3YXxQJt1HnR+R31rDTPJ3RxEerbWA4Uhiv9zz34+8EuZ+zZw9p6xX35DdwRygc2LXZQ
lb/Q/dnRnCDlcJVFLNMlAasy5qoDAnVsl8k6LJwxhwQlEd22wGQ21G1O0cXtOmv8XZ4xu/66mLDG
F0vwLKMyzsCEMZiaSk0193pfYEvwE5IHnsI0ksdosIO/hyJrWP76wmZqjmMLXENFLYJiDpGHAmGS
thensQkSY8LC1QzSQ93DAYM2w5I5i+vRywBNzBwJ/hAYO18shvw1UxLH6tzr6nFpy2TByL5/utHz
/rYFgvjldHQa9dcGTsaBHDFocFmDCu75U0lW90qVIU3Hh1Q2oKmDrXuX4AOap+1nfBR85C3SCN3p
S/9bLAjVmEz5KPsktoPnX8lV7ukiaJKy8K9IzZsGQb1fmyUdndmNomdct8Eo/56vyL0QKklT2F92
82DOOeUoGzGLn9V1csINZb0X70tgo7FJfRcunuyTsOTDdLj75d8TzmhgHbb1JtgQqoC+b6NKeGE5
wzuAcl2w4ubOoNlhKTzTCEwQjKwTv7/DOtsscIn0ls6nSWcPElfxaoZPF0GlYDCH2qcYTayytWqa
NFowXoPzH8wO/8dOBbRs4xSyghsIyxrja/jxR8nezGMRSTVkNWVQVODWlKp/t+zALlY1TjpY96sR
wE8zwdaOKTrv0Qi8F+ruaiDMHm18hriAS+YknK5Sx+KgzpEI4NgA3TpIObyiMSGhBtJmKtiOEoJx
dtEfDhp/kx+mXqw0wsNvECapOOCGDKbk4yj7jM7ELFOrqYACYKqDhBZpSJugkMH6w03yIs22MWNN
m/s40jdV27XeftAGlXJ9z3Eluci4jcPtr3zWba1JPv47CxHAmvREd11msGPBdV88l/N/gJfJiFPQ
RqjSwzuHiiQFL+3wA08+vtxNLbIZaZqd40ET9qb9/Vartxv/0Kswprp978c1U3Ov8E5MKsFis65h
3EjQfqlY/36d1b1lbstGV3lrCWlsqzx3rCRlYR2JFzCU//B4ZAVeXtOSIWe/KSvVB9NJajl+Gqat
aLxNSYf5+S5gs5QHzTJVUEuSqmpdUOpidHPOr1MhsYHWxsakP5ITkS1Fmave85e/ULMPawrrEsP5
+SbCILlbZljrU81Ge7fCIHIXR6HTxwILHgFNl7MpJanMPkphGfHMStatBpOa5AA+4jYmdyawCqW3
2pJJ3hWurnzSStLWbfHBwgdejKdGn8f9N5e+p5+5UIOfy6mjbZiyA7kRlai93LNdZD1KaxhOb+TG
YX03r5e/2jmrY2yWceCXBGXUtcGx9KEiFzqwKqPwsz2FE64aEXZP7rQNZJnXepx/mjKGTTdV4Z9a
Uwu3cZa+6Wk9ORjo3VfFQlGgcCPz3021pkMEq16dnb7RK097Pdx7CW6cAiSoPKp47gOBPM0jXJ7A
Z453WZ+tMXFrRdzsVefM7l+GkXgbmb8+zirMoWTFnLKXt0wLbrOLhRL68OHPPDYhxXdP6oZ+bae6
dL7cFLUf9yDN/BvUyEj3PL5uFZKgZoo4L2vLgz6nYVMKyC/7/4Awo1SCrsEkxpWmLpVPWVX9FbRl
X3q9Hz8A2XxqMd7MS7aDRb1e/BMWSstPsqsTRbyEufi6IXfAW91hIAsCZnlfy32dajhBN9eu3q6/
0052uWC/cq+RW4pFahK/ldB6RxSKDHBFBuCHIHaFrMjfQ3yZeLf1R0yNL645THbiWASoQziChTRJ
MU8FCsAOF49dxxF2l1Us2yxmig5nYdHfbBusH6XqaWgxsOE/PN7qlIXWDr4kSo6BJOWCAaso2jWE
Zu8QdvmvVeuwjba0sqvnUkxzTsS7w+vv0/WsVNG3f8HxiX+eUNivf9b7QdOsB80fgBxZMFToJcJS
+Kkt1UTI+n6sXM5jRsOqknfRccmhy1BkfBVPtheU0yleyonbmgHXC/mWR1X/uQr8jWySWkXGLzKZ
JXYZWkeYzhvmErToadAeLsDqY6RzZ997KXbQuSLzHxNV4ntJBy1XmBy7aeawquvytaJAvKhjFdgU
qmvaGqHMsKIkLospTNN4yK0K22vGPSz8fCZ8EAdEGlFUU6+/WDP3kN35i5FBELbYIr5of9blaMQL
bAPC3ciKr/RtPUq7Bd9M5z7ZOx0XeJyMzpFYiGAoFvw2nILLcC6uMCLr5KZenIKvQ1NG+b3LYYNL
wuDEOnpbuy2H8C+CRusW/ptJ/Hqh+kWa39C7JrWwIepMgB0IZydf2bYx78I9i7aqEX7CJN7149Da
lOeciTfgmY3/wKwsjMNLMyEB3EYX25uKkaRac6cgvZOSWTqwBIfEbKmkmflxyZu2cOEqRXZ0lK72
dfJ7gjnrp/5zP5nB/XCqIa5FdfjEl1EEWioJjuFIJyRTJl94+XhpDYzgKR0UjcG15JbMDYx9oVQy
NotjayKu8K7F9yasqpdgDvLXnKb9wX/j2wDiqbeEKR5qK2ZdkomyV9fQbqb4QTJwavCwT2sLJLWk
3dqjkqFECn7pGIV3ZlW1jrFpHoJBAAqmr+/PHOWrQF9r6T0VAN5DjCV0LrERjZwaZZ+/o0n5YBd4
yIycfLETORtWpHUNI6CFmQ0ZK3PiZSIX+lmxNccDzFNmp0BeadqOVqN0A08H5tKAcc124cerPtRe
HKFMPfRwo3sLiVqb51zW4deJEUmg2jmLKqdJFYiqAQVSVEKvuMRXJlt9hgIB3r8jOkVmDfY+F2wD
rv5wMVa488Ecj0Dw0r5lVcaOD/s6sNuV3BgCqfIHJxoI885SCtS9tJgDr2r9BfVW+UD0XwYwOlDb
MVGVx+pRmK9bW+JLEEDMqrg3tSLUb++mtyvxaJfi1PDTvrJ5fGW8xDkkZBzOQl3xjpTDM+3DkU+2
voBDapUuWmQDt6L2lcbrpO531pzLTNzfgcAbL2u8oFUwEGEtE7en4pd5d0erSH4tth169Q9iI4qi
Dk6BZxaAF4/6whDwJxMgu5ZGMo7PJkEv8WY1KTGoq4FH3qOPnPbDAvJUHk7Eh+pQM5nUmBWfWFuV
u+dff5QSbOZGAn315Po33jmBTMc+MjKY5NEXqMW8sSqKjV96l/NwHRZ62Qju1/dCWuz5jj+OxM1O
f6BayTVkweBNpJbLU6ZI7+Ay0SVXdf28XTs1sz1Ta4lGdZzhPrcNiMhCx4cxH/N0nn4BDHUsLqe2
SYwoCmupoiRuggqKN6swt9LxJZUfeMB629cbKK0127czneqXNrmHa+A8ekqM4CuXnKuF80S3TIGl
h19y+iNQi9sUIFfSkG5AUAC9+VCVn2uxiu+y/kUQDtokLYKqycUYWdAn1/c6jpWj3KGhrYfHagNJ
YoLgGhWQqS/RfH2NgawRPuGVoCczkKJM6MPSkyQJaDKHeTRUTFAM/cs50EIZ9V8s7gsssujgHlTt
yXn4VIcKgNfmEBTvL7p059Mr2aMoANEtCpYq/ogf7CkevnDeK6Z4gG0NPcfZnDKeZDCqL5JnIZr6
DsocsXpW1aiy8NGKNI9mXdpSThc/dE0X27AsNRsPXjqfEpvrtSyl9z+G6IgLzZhdNZiq1UEhZZ3v
yQtowW++8bvgc/S8lAIZvb9SyMaQbhdJxzd9LZBGZ/bdpq3A1Y1jGQPnL9VNZrET4HifmT5e6xy2
lVu9+ZDmuoxKdEwkdW6535PwV4qCVJOHOC50AKg/lgZgd9OPIn6wKbl6pGvyp/O2BnulzPrU/vbl
d5RiiQO4gRAKr1ykMukZSusjlIp9ESu6h/7iBlTq2DyGQLN38J7FLKs2Y58Qg5KfbfnrSOAXaz05
YqNJTEucA6AzuouraOLUXqhCoQQOdpJJ2O+MkD4Lxx5FnLdLnklu80pxiAVGbkJgvto9ELFmAJ29
sxJEOF/PFnN23kkGRSYkW8EdjctcRcWP/SG1HXXCreE2vcrr2SSMvWVcIesQ5xJHW/wX4PCp+FFw
2t0gpOUecZ/6kMMXor/GreeSOOId6oekc/Kn2WSu54sIVWgVCC426ib0qrqZDJ7MFyrkApLgNaDq
kYiqr3pTZcPsCvCXPoy9P/xS7qhrfEL5tuhzHrF/e8+8BUMYak/qg6gijADfQxYxVRWZpR6OiDZl
EV4msW/91lRrKwiMLz8H+H9V6HsxF143oD2riXP6UzTbVCc/nR7xgTkVlvFsZ0E2Gfw+7/UMOock
WH2GANR/uV1nvT3hUtTWILYXHfERmPfkpqndEHjtI5e04QomxptmH7QNLrayrzOzWDFO96WKIKxS
7Q3ioGPqfgSOpiX4Uz8pyQfXJW2w5CP/BDa+HHU6+pEX0oftdOu18ENi95X8x2Wx0bku9wkPHv24
CwAieKY9tcbQZkRU7vF/gjkhAejg80BAg3CrNAWCBooHSvO7w0UcPmKom9uZJTTyduROs95Otod3
k8VqurU7kYoJgPe5NYpTL0Nbcm8Rt1UhxfH/8u/9Fhc+H3nWjoRE3LKSR0l8tzYdP+lqYZMB7XXt
IyIYmPel4gtLOrfzYekkKcx4g/qDrb+oOtyqFuj6FiDbkx0Fzla0/pOSR1j3LxM84dTAC9PHK0AS
HDAGkY6zdk3DFGoc7IGM9xfDSiF7BGICQEqP91AwurLJiof3Muk4ee56hyfGQzzcw1txxaSYZBa0
HHSgxgZeBVaqqizHOklW5YIGg12k6lNYtQoGDH1xB06pf9WkKoZfyZcI1/kFyO51ITjynUz+2Rbe
oFW/K/uoHFi2Jkz3ev6JVD+W85qUKwHl3HhmC1kQJRMgU1nQajiZ07njaG1IK+R/B9RvBSbYmEjY
tzQKfqJ9A5QKUK2TQIiWYhYHGDb0FGFBR4rdZ2rZMs/aJgVAKxDJx8arVdQFRLY2e7YFiJzg/I/S
i67QoMLqUC8xTm2qshTeVgnmlbAZoRtcsV1I86UCSL3UMJq0NqvdfyYD3ZJ4XZA1v2IndQym82Wa
gizW8lf68UJlsuIPrFz4LyimWWSsrUX8qYZRXKXaPVMakXwL5u7Rx4n2KPrhMRmp13hBuIG4ykE+
lNJUZ/N3hEeaOtP5KFRDjaS6v4tqCS7nyt8tCaAXt1AJiNCy/vicEBKnya9xvWeN9nfze7RnZE2z
/TNjdMz6cyd8ioeKE9ReNckTSS7QK/m/16HPlK7cvza6oN2G3HSTQ4yZJWmVmV0/tyQNyJVIu7rD
qxdVrzeFH0rhZiX/vopjJEkJTfVRBLqQ99+1bufLlfTtwE6D1sysDED3c4INMSt9qxjrHULrKIQ+
bwOIIwfdhPohHx05BEklWfSWjhomQfsZv32dexHGLG3Vb+AWezlKhQtULrs/bvnP/jzC0R+HpdOT
ezB7twclT7EeEkFWkFrOFYg6rzlCoB601LoZkUHNsQ60CO7bI9rkZ8dFfGwa8fHR5lEMldVVtHS3
BKNJ7dM9tFSU+003eTe5nJsWLlsc8zu+E7VYm1Gm4BZu+sH3cD8P+wu4iKGngvt4J367wxlrTH2g
AnFIjz4aURR5/yurYi3Dwk3TlhoWBfjJJG6tIDXURW3wTsYtL3DizPS/FQAFHl0pznkGx5tSZDRu
w978h+B1jaqhEF7DJZCOH8s9wpSU2iPwM3tyvGshSz1b8caylkwMfaxedtYzjuO1OX/ln3ujvcLD
JzjRXIJ0/J/L7WyEsecu80Ti268MR7p40FH+VQGrGR4QPo1AWF6wARP77Imy+8WzgZtRk5EQgNPS
3Ugz1VzyaQ2+OG8hfO7PsK3gGg9iCE+XA6DnTQVIlpJywznHhXVrpTuG+dV77nUVX4vCHho9Yl/N
DlvkaFUylTdNhMlpxNwMQKOFvCViNrrgFuNe+AOQTBIKd6yI+6zAKxJKQ4u0GeOo9RAFNkjfBc5h
9JRAStPvz3mVIKXyqNwnF/phpGPWochhIG1dQXGwr0Yb7ReXYzRGdnyknD3HE+dKGqV6x33IRcMl
wzGf31ipUVRmXnVY1p9boHFWWw+ZCwaxU+pyp0ST0xzJzW5iL4GlHthgjKnEJAy5oAGinOJNYh/G
lNO+SXYcZzp6CKj2k1i4RRut21EyXlSkjAGWVJ6ZAx7TxqWsqmUERqs9yL1t4wkqenfGEkHW/uAc
uGHa/3xWJ77FN8BY6WAuULzVwc83OA8W3e3sriw3tZNi86W+HE3XaAuyzSKjDMgdzf24nEvzq+Sq
wRl13OcftoAFfQsdrOGn7+8JcTPWsR/yZbX57UiVtmJ6mL9NHiq8P8G7kG7rUlaPb3A1FyZkLr+/
eYPjJCLkySywhglGi3NUqk0Gq6+poigT+D/oUAhFhKHQ0EBL+e1+DeUdwsdZyLm4ogIZzZZKzQdT
HNKao6hrWp2/wxXZ7CPMuzb+B5xIkK5axriOI6lJF3prV6phxQZSl4wcIhuUPvIxCW3bkp46sOwN
DaYjRVfOkckh+xZWHFVvxCI8UMjqExhYKP86mJlzXJ1cWcXWZd0wQytjRIxXCBb5KWitF3w59EzS
T1uXki7EZaOnB6tZdwMZERuwIGFB8YKrTp4Bdk/TIBOE+Fvz0La3zKFhe4yrzBHY4kax7CfddOiP
nB528y8TED39RG1MZAd2/NLyRCM/Q+J4daKd+MN5vbN2ggzTZVSIRcx3gKoHPI3wctI+LysTbS4V
vK4BptkXzn/ToMsWuc5SMfwT2HqqPujArxlK+6o7BgrjA1kL4McaEM+MmrEYka+H6SVmi1C3eNso
4AgSb72uj1nmVuwJRo/n8XQRJwlT/Ep/ulMXag7TMazE6+orCjcTsRg50mLC6yPdTTEeDU0fgVUQ
h1/nKFRdy15fVfxp+rX4e1/kNpG/otoNeiz8/m89kCPq+oc8rsLFd8jxpOjx+Qc/WsB0dN5pPwAZ
tTVk4yzcrBW5KoNZpK9X9vC5hPX75+hL0AG7+R3SlprmM34J67712JvS/La1uSwov+Bojx2ua8Cs
8+l8XMueG4gPo0Z+vNvFSgrZs2Weg3cpZimZbczW1aHma2r0Krh7wcBC2tQVIVUnGtoZOVUfOIsK
pobI8ZOQQfQIpYUT0B5xOeatWijYHISBLssWDXa7pYVqUYEJHNjdy+bDt3P2AQPZ52cXvhGglAxF
MRt1975Nn29sKAiM6X0hXUuQeddH/B84bKfaER6NrOUezVpn9iTtKNa7uiJVPXlM4/vS8EyHDhaV
L5FVftKYPI7GL8hl4LMatc0JlICz+9x0CGSNAhvsvykYwVXFiCljzOSct42iiau6iTE55OV05g3P
yZezJKaGcs5+nG66tT+ttvBmVlpHCIqRMFFTlUm8xaGLGE9Fl8ahMlNxscjQm0WkAcBjKdWv07NH
xm/+ETp2vS4QMGzrFSDXrd6dfDH5pCxc5BtWja6DPw5B8Vd7UNe6c7TVWVWmrs2Q3BbO8PEACQ+V
5f3kaVkH4kq3ss40UcztAWz/PIO1hlecjkfljLwKegtWZ/5cGWu82Li6qTcdVObTsDUrNHFG7Txv
FsOt3P5kEk4JBhu+Ojd2dnb1volPN9a3szgBAIpqv2kbjwZnUmluxnSASm2g9ciRVUt4OHhcbph8
pJAIzhG2Fx9TqBwiEkU/SkxNVBPPdG3MzbNL0uyeP7nMEzLEwRgi/zJ71UjzVJdHfO7Hz2cGasCb
h4xD/DUMwVbuF+J9HXORwB5aNYYetffkLJgokti3TRVAIP/BSTxxx7NUQXC3epsG7ZPt0ia0gcyQ
KfUX21TkcOWXq8mAvZR1vvk+AOAOyTMqfEvO4Q6sdHE7GKytggowF/iTy+EgIekht3hUdQbDYSfN
hzZBAU6fqLKlp/Gn1W8Jxj4kY6X2YEyBk7HXCXhFfisFdhdpKjhv9F1EnHETZIyjNWzeSBOLfhvh
5673u4i5f47eNHJ4G9N/IKpJqWxqMQqVBSbkRLIgiwrdEPVuG6cSVN/PL3x+SID2cDojaZWu7IJD
DSnsh94uZiSLou05kLen8EYWc2X8TuoPK2ZlXRu88vQuskZJRTA5xbK5amaad5p8QHTWPJJMZh1w
z8PpLYkLYEeif3WZXBy7yK7N5lHqq7NbKvOef12Tc/K3ULlhCXNLxpZkbdH3JeQy4/sA6BH1+L/H
j3weojt+tdbF0NzjeM4EYLFOZgpAeyrNGDv2EFi1R7JriVm4/kIyTOxCryl55yMBoR/saaE5RQH9
LmDwb8LUNYoVsJhVHmzkClEHJY2nPW0FftMwHrHUTQfzFIjEBGSaedxyeCS1RylI4kPIHHSNb9Yi
A0WsrzEyfzHa2WlPDDBqYITUKGwxfi0ot9SGk79DT7Y/S+bC143GEbHZAvPmcayyUFNwpOthwU9w
7nPrgrmEctDI3zEMyuAewsSd/yFAYMcZOXk0PQjuT8lzeWEyZnCvRH9teufvi5/QhymJ/L6RwwuB
+8LeCWoLuLq1NkM6mXc424wuuerdWHzXm+A2prEQYz/RTLqlCkt5rFhFApWgw5KKytojLxaGbqOW
hYNk+mbP8henytS9s2bCDwq7enFcYHDnkem1kgxA4/Xz0my4gbZgCCS01K214pRkC+My8BiMGoTh
acRu7ePuJ2yHY1UB4iw6rnBT0J0iKBw3b/aLBnnURuhT08S/r19INqmgnOVuGRrej+JAJ1dUl+DA
FnDz6us5wOraGaoWExUhcf+3Z+ry2av4I7lKcSq1iYS6SAlMo2quMVXBfmPc8gAq1h05kE/Tnt6N
hKCPCS8y9Xhxw9UiisVrEDKZTSj8SzOzWnt8UdBJgrY7CEzqjOlK5KF53c1D69ZBb2VG5F1FElTr
IZacqNWEomDvYQA/IWYhdyyEq6em7VKeGAqKw9KUrBURqc5GQb3vn4tGzvUpOv6zu0h7PGGwsPny
DcgMUrKkqgiKfPB+56V8x2Ma8FsDg4ViXw8rtX06KZNIabWIEuIYPtVo3ydIfR6p35pU0epXHOk2
mTbc9z7TnOyShz4Z0hsXJWsEUEBsLq2uPfp0e3WV4OMnaawHvdb/eOmqRZQ2dNWh7qYASY9c2t51
oSeMFHBOWLD/c70W+r1+PmaiG6b42RlvuEszl4znVVMSb+Xlq7YSMTn7c4ffKCsnUSgP8esfIflg
Ktzb60DZRSyL+ZNZCHX2VcAeGriGcvnmXKPN3KbVxB3A0D4dYaWrclZztjqkE/4W/dMz3s2meBp3
hiDmlEOBSbg3tqgVvhDEZVlMsh9obO4z4C9FoqRPmKbLKBJw039qiY6GH/6wlJUtfTa3cJc15smb
saOEcTV7Qwp6n/gILz6U+qiuH9bHk1+ge1vUmGtKcVMOdktbTMewV8zJSEd4XB5/9SROop4bjMrQ
BQi0rtw+4ygtEcoZZGGqjD6B9G9v8gDtd/KX7XsnUjy1Lw19aGERdZ5hEY4YlHMCCKzx54egic/B
KNHnZmEpurxwlVVOjfS1bVJ41ALjtS59T7iQTZvi8VE+qepk5aIJSSyFWsn4WBrqRAlXCRiA2SMF
dUFBEUF05izcbXG1JFtTqkblTRK5qXduDewVekXT3MZCfHnEFmmsPdegtL4zGE1elIiNXBEk0X0w
x2Sfg3MAyC3ZhbH6Dj4FS92wQW8nycBq+ckuH9c2PCnV4DksRCj4QZtRegojxzeMaEvv6Nax3eXz
Eq3+Mmxt8xuRT3HR8ULIlnhWIl4r1xrqblUeS6o0L2QuwKvVb1dNSym1+QNGURKfGkuVF4vnF6qJ
PTez23tk/yV0G1pdkMe1v0c+sv+AFWYRvFMiVZjtbCuD1qeXPp5Ss0lPPqKQ0SFd1SqttfGQDofK
a83PHyoDmp8G7ppgUxZUR0QIAw+yBD3B0s4N8z8rXJq5av218sbb+u3dAXWFSFHEnzGwXQds+XXv
ndcscGuq5V3w6fViMryEp6bVeiAYXzyiYNauLxN7pS5PH81ZX9YVhZHQgZo2Oxomfn5TVtgJzvmG
u8dXZO8g7pTXTf8mHl2gSVzyUp9K/3/cAPbQRM5kVQVozFVaZdUuRFjFSpp/kSzjJkTchUGkIp4j
EewZf9xz4nYtKzfop+ruCdw/gH9iflVxnbGX4bCCO6q5dHBrupizUNP2fuLFY9OInXCvL2sx/IJO
CaBc4rJtOR2IXx4QqxztssBmbsq1SmXC3BGAcTufdxY8Yzhmu6azVmSme4G99gICg4rwN+oPbmth
EKHTqdjTRcxxhY360XzsIT9lAWUex2tRLWZt6kizz0JCLvy8yVwvwY6xo3alw7uVkF9survwCKt6
njirlstq2Rpbp7QCS5+f6+6nB9uveRaxd/zQF8mKTLyVkq2cDaI3LRAL2pY05/PUnTCctw7AzVfV
3vYVBzI2zU+rDp6gUc7Xz2p4gsbiyIJLhM4xzpaHrM1uvbMv3BJ+LIKenZ1AnELRP00tShRZa0Bf
KPeNO97JaSu3oRMBGIYoUsPYFYCtiqSg2FipxiXXHOQSv3quD1ClgqRgQHAFN/y/65Z0LmUxPuIo
cZ6CDxH3jR1dhE0QdNwQ+YrmTB0QuNYQjfBTA2mn1vTGS4HQd2ow9DgdldCFHyqIkHbvnJxpTiq6
77ysQYHIF8Oyey8xPVWKcs97bWmQ0+nMxFxQf18pD3a94+3kL9pAaIF3neTWveLf3l/ZaRCCsNnC
MgXUE3pAm50JuyDv/hBRaKzH6SLqljh+Lazw/lmqr8n7sLf4UHxDrxEc4WS56h3d0cFqs1xtuG1/
ClgN+rJOmN9FhwUdvKdrRegXd/RjAErlGcUjywdTJF1bHW/dYpiitmeNm6zG+4ClxRUtfuMIpHr/
HUpRShDZEGJTwPCuImrpClPzXpekhEDrAbUqwbqpd5cw0XZsj6EEZzCwaX+l2zfIqESI06P8vMkE
tHCnRLZv57qjiuyucxrbwro76urMR79I92JQV1JjsZHckniANVsmdUOiwds9Cp8BaFL2j3uVunOk
bzxTzOoUNWlidy5AUqF8A+A/yPn7jIjIugo1b8zQqYtsLFgJGN5Wb+pTlfx77sAu2rXXRIcMsDF2
7pZADcz8wLPJ2xL+0yJidjxhHK0vI/LEWtl7eIdjsxVGj2V+SWrEWCfHXg19ICiEDG0uUq9LCysV
lo6PvGe+31LZFeHTPbBUUaJ+Gr+Gdlx5Uv4+tlzzxstWLZp7sHuPOcrmNPpzVpuoD/Bn09u7CSZt
kfwJt0WCfEBKh38W/W6g8OKK6D/9+xsJHGGjGfcW6YGXuOLeL/ZFzkxnRlWBRekxW/LzYZyZecjA
IFn9aOX+M3IvUB7QK/Nyc10wwR8WtloK6uBoyfd4POej+5/ahvvvTinTjeOcIGaFrJ7Xjwzpy2cY
UpksT76TcZWV7FAEW4dA1zTTSAu02NoksRdvLQNkAidoQxGyXcA2sCmxHJTV4DbJS7HvliR/tkam
MA4zoY3ebsbrgMlqhSiZxcReztP+1n2vt41/txvCfgbS0us3MnMwhI4KvPDslGvt7YFT1onqFz72
zQCvWqBBds6I6YirFVEBwRbsOc6XAfEkhyqVLWw+Zp3C8EGq1nZXp2YZbnQZsmuTnz1/9BIo6FPs
UkwjwggrEfzkgPuC9NvkHMiJt//C4fzHuwDjhv4SBxFh56bQC5zayLllJkdWUG4h7OqDK/Er519E
c/mjF3VFhIV7yMmNFwRnm089IYaxdDloXjE8RhrbGP2+BoXnlIglgS9fGq3FJsFpq+E/GtPMmymj
JpqyrYAyhw+9Z77mqo4d4rhcXShZ5obmKwIKtSj1inMokHvJdsXwLGHnHLKqbFs+nxs9d5uaAnnO
fGQ2L0rXAbMwdq6yHECS6GYDGKAhZyS6aslNvmCnbz36HbeyNCZoomLedDD7tnXqrLe0PlWjac8h
VHSn8366+i/fISU8z2BovH3ORON/JgXIF9PoI1058sJjfKmSuvWu6Wue7R49bic+NO5voPqsjajr
ZA8FSdWuphspGhKX7p1V6WE123Tk3AqDYNXpVGHrv+ARNt5wmtYCYetbt1USGoE6tfukpWkm8Dtz
zf6+WDjzvPIq+YterN10St9Nq1FYRO+AWI4QnD16X8p+qai7ojteuDa5LlFDc1o5FMSpq1TqzI/W
s8mkyLp3nBMs2P+3IizzFnpebljHkkeqzCS+ra8Ypsggn7HA27cY33kVIUY4pNvS04dt8Db6bAnl
dxgNtsK6rY2NAxF8KODRHbgP4hLd6z5JjxBu4E6iQvdoKf/A36x4NrGVpbukJmBQOr7+/MU0qM36
mrRlu7ryM1XN06+By9xmerzlO9SrtkG+acxdaUzdmDLjZYJVZXzl9EKo1YnWiqfMW6f8a2t8Uvhg
uhzd6shD+FU/Ophir/Nzzk5C5X9Q4s2i0r3s2o0/2SqlZvAVkaRtOUdUs6y41WwWunB7HQyqutL9
T4B+YaoEtt+dJJPD+5tXkOsG17Uk07FS8GsCzCVVFDaM999Z25D+/06ikkoLoi9bnVidl6SJkqSO
MgQ/cpZuv6oLqjuZcpELtUzz6dpxJXnJEGavqmpQ7fxsMk4MsnqJcSxTHOMAN7DLMt28buB1QS6E
qeiU58qqt52LYd0wsekSd/9asO9pa9UcmiFTFo7LBqVWsjmI5lRbmdecquV6uL8toRI1k3utvslR
jWL2JdOC6TVtcBpubjOG61qh3iIrLVXxAn+/DeGv451j1CmTkdiPaNccUNrVRxKqI+JKu9N4A3iG
TZSOMrteWx1PElpjWO5KnkfGLH/i3aG+zYB233aZ2w6HT8QntsMJU9n+cU5mT844zH6Yfiu6Gyuu
5PfiuhG4TcE3WR+eu0DXh3CfJT7OqjUkz+n11Uh1X871PdISTgNN+O/re1fW2HtjX+nJ/v6jVTiM
PNkVEQKcbSLY/YnJho0IbnArneguALqPUQ0rxx7xGfI035xVBCV666RW4DEg5pPFm7cjCePZtxwN
oOpiiQd75kPiHrN+mNqdvz5NQXr8NCALkBrDow49+5haq+wbxR4ew39T4ctEeaoP9/MBNr9u0kIc
UCp9FCRRK/Tvn9trsrEl38tjo5K4OG8xRevLGsIxouHEdABX3X9L4QAdQxgc4+3El7qx1T9P5aND
MVbTe1MUZnKuJLWmYq8oYWzA6djL03E8b/t1XKmeYUEQs7rAOLtNbu/XVF5M23WZvHU9VemIdOYe
F2TvxM5TaspUhUSoIn8AUmReaH0klhlIP4ZRsS6QG/zggQi90fu31FQm33bFScykB6tF+80qucZZ
mGe35ndMN6dIDV83MWtcG070o0Jg5djrZinKChE51yVgVra5B0A+kQv8F7kqnjT8Di8IpIugBaJO
6knLHapo1x+vfTnc3hUhYRBjG0P+KsouhKOScrNazIj4Kkw1Ld/fbbiB0RuDcDIUgRkWnYqMhxop
lzuskJBFN4K4WNnZNsgkroc4HtxYx0zQnmGPI7+iaRA+2z7CJnHdfajEsnsElNj0PPkZmybayCfh
mOp6URCDJuPpno6Uk4Zn/Pe37EYRoiAKi27sMS2FQxrsXJHHX+ri6ioLdz7lUYyqLS1x4YcRF/Ml
EdCssR8aLmwARDwR+S9btffGAxR3pYdh9hHuZPBz5r13+ZfFs8S9qwStb5/dJ8PqBHHa7GZhMEWT
KL0RgI2ZiLZMdRyxIeSmaY9ehRqIyNW0wRdpCk03VdImHkfQzkAhIhf67cx6Q6UZzoSuyjVjW3Os
KYzT7M3+dzuS6nXN0uXZxAaCPvy6SogftITc5XH7SNxE80yX1QOn/+vZgwGEBwP0Uvmt9Gv8s8rF
7E4FJcGlA/bAXFv1OeVwMNdkedWWK1rYAH1Em0or1GMDI9yEE+SR8NRorvLd56JrWyd3bLXkKINR
pHCG+RXFqjPGJFbIwQw6TZr+VfmadvMMs4QyoPSUKnqnLTCE7B0O8O1xSz8U77vLmQ0PH/WKPF6c
cG6JTngOqnxZV1Q9UpF3qEytjVYju1kl9hjdsZ3QBMea4VBGqwhhfW18JCaBC88qe+rw+IzhiFYR
8JtX2PtsBaYRz2y6re8bOWcaKBMLKaxkW/HXzRyDkQI7Bh5hl4ziZrsOtmuEKY87dRRcCnrWGKyy
b2yVJfLG5lm+XJMKC6hur0K5q2JKLk274nZOLqi66q7atN9P2lKAYlGz0r79IOR5/Ob1x1hqLqp/
qjUIgFcRtK4kokA0cUFy8DzR+xxKSDjkrVAixUs6slAHsEiSNxHvywQ3O3lOubGAHCo8WYAxioFp
ymYp/Mj+pXqzHajDX7pR8eHUJ8r3Ppk36vtEKAL7BqbM9SwNg+m4/D79Lh/kyADU26kQMOyH2Kqp
f5xuLQ00mmc1D7KuH0TgOvq0n0mL/d6W6wBBMgvL3alH9KdlN/FVAqZCQ2F/46Yn+LxunMo+pDij
J0IqDXzt6v7N0gBzxH7v6ntqKATkBLkW41oRZYA+7FE+Q6bKdhrsPfKhuInBRMy6G3KUD+4h4y70
tN/1dwB49BVByB3rb+2x8/rHjoa1PhCGlU6H6FNqGL/KpeAm8wYaycVApRbE8kyNhUg0tWJBJl8M
BGLMl1VI+0t/pMoN2zDxBJL94QAKrwEd7Hig1BI+lxVXHb7yTttVpTEmi9XRFqaSi3lobB/Fy5kW
vA4bTJm53FYuavZDX+f1wC85XHtGy0BlrY+DRQgs2Sw9D0+2csU90HWtxu2nsfJlOZZDOgutn5w8
n3Y3MEK4Y0xlCWX6hvzfwkfRWvbQiSK6mkR/vJTidIvKnGYo3vQa5cea03YdKL36quRVmRMiyFB2
d4seby/+QtDlFl6wPr+p06FfEeRAKg23AfXSw6cxL1l7nh8XNp2oR5U1MfvYG7X8IMtpvxQyk/uB
/38OmpY9+tMNh9g+2CWc4bzsteP2s32xD4D8OxqYfwa9Wj5o9qNcZh57BXMMDi+zHzrsFAy6A2hc
2P+4MYHXoMe+5qq9iluNcK2zI3FcxoKK3xsN9fd42WlO+HxrDZUDy+KSNQW7g8iV7KKSKUh4m7Xi
pFaX1hLpU+OSy0T2YPxmfHSX+3LCFjjsrVyjmT52yLFtbuRePOOsLGVm5tfdjOA73ZfInwFwM9ZE
R/HENm9au5gbUKqBhiGQjNyQAmaTVXjH63eNjYYTgB3XvUX4ggvkl/TUL+qquGIxKFsqrZuqz6AA
uAKQls6COYe9IiOEe3MdKp7gU3HkLi8ujdAIjAxMX7H906P7zriAdk5HXBrNpD8Q+32HEYHOnRsZ
/yqg3SqxfrCRelfOSR1I2p1XEvmPwBwOyXDPU0+mwwlhS/REVVBVa7lVGiduEmqkTiaUGZKLqpcI
ygP/0dJsveKqELaKp2sQ+Z51T4NrTTsMxnMx9jh2xi6ymhxW0CSIiO6Hu57K6BeFIzgkMGKXJJMU
7AisBRyWTXGPMV4a1V1WaAVfELiIgQXs5ICrjaMwHZZv9oNOAwOLZsz+TWLa/jSsQGTgXmYZqCbt
VR2aYKUYjG4EobPBnGDQ5/THGbe/8lN1O1LGm2bESgf7zFAalr6BhvTfuwWYwEmU9fq84v+d+C0d
4YIVV2kA+/zXAWUKcvBp53iq6TLf3xWhwA3FzySv04MhtiOCMjq3KYzvyevG28QpBwgoHV+YvdOl
X21RIv2GQG3Yic+Ae3CbBWOZ8sclSVKmdgMhMDSBhWrc3xvy+Y6675ypls+gOi3iaazttIY+INYv
ZUi7pSoeYMsxmL1ji/NWRa7J0UbHmzwjZQsWI3FSD5MnpX1aQtnxWki2NJctJG/WlF0BOQfwUE/h
1+/n/Um8DTM3z0YI4dIrZurIVxUPWnzrsqS59EM8khrfyviIuR9f/Q96THNr8K7O4Kp0/GnmESUs
xpwPpcSOTqhjZWJM32LWEtPXMh2iosrM6OaTZTdMjPqB4Iy6cPsHfpDe+M9RXnSdCQNF5tXrsOzG
DhmSdNajNSP2+gqzhMmYmfk+Jps5ll40A1/5jVjY263jDhJIU9rsWm7Jk6xQnFEBGtW6uTeIjbIR
GxYFQmrw9t51E5M1oG8svKZnTLFj9R8jrBOdZDjkobIOTMvy/yj/7El8ci6q6v3wnR7RElM88pho
9Xkj8UJ/0cKL9DZekjdczvy19GEJ6aFmFx6Qmad0JHm/gvDhwn0S+jTYC9376XQRGNEfir6OsEHh
6GxnVPZ4sekXBHLZygeYpoz1jCgoCgBb5mxUbU9ogXuooLkFyAUys3yJRMo0bdPrwptkOkKkewIq
t1RjpIWBgPQB/uQSAYKKdgnZ9+z8x/9BD7D8ot2OdOEkxOvdc6oMlt0Wl7bEQD0L7x1ncAli33UW
CCWHRJ9O70m9Sw0EAnW6+P8x+pWtfNg94leRlswJ9pUS5zWMhXZS1nXCBE98V8shCjjR0EXFLq+Z
rtN6Y2Fja4v+QEhAErXl6CLiRbWk+7Q+9QJOCS7daT693ywcaRLgnhUzngTcbE3+eUHW+O2wXNcH
4uRiHMC/YfeJNxF+mvn8ixM5ZGtUlov+PrsZtHdmNpqFt9Fc2T/AwuR2ZkpVE/NpelfPeoYFdSkh
C9khFCXymblSaCbJN0X4MuGsQMBuQ/MRyvcPmk+GR5QOQpD/0lONukfJX66WiGQghXRDnZHXLaUT
ks6RspWYVQ1vPitVAp3hwZygc10OvtGBP/9Z8ZQTJ2PHIYiMGh3OmTHRAbDQ/k52XdSvlLDTZepS
qd52QOSQ67ECcGjnvITbUMhhyuFccp3reNrhEIN8dMDZ7i1tC41tc8qOmEgr4uf06RU//r3glQnS
LJtEAzu/X+fGexbIP5oSvwug9oc+dl2DnGqMcioALzalHBSO+Ex+dxw+33nRkg4zVlia0xy0Vvlb
6vC4kTugB6o8DKxgTq8R48CCQURp6W6ibjLyauGx74o/NAfqKONMT9YxklyhiB0ZMHkk24HfqZGv
mFdLT9c5/aEAUhY72RHXcWGw2GrCjLg7GWPx0EV1bXccAXcLSjz182QISB5E1xD5JQrIsh0bMxg0
Da+E6pVXDVginqPKJSqY7Jw11GL46hQr56HWeRtVCn3FCBGlyGje9XPFw3ReP/H+c9F/SSCrY4bx
K7x8UFbQahMNklHDWq9WO+EIrg2DB+L3+k1E/0g9K7J6TRp5nKHZR9J58cDCP0DkA1T0IfgdRbTK
F375MPiaPtpmDED70rKgqZBk1aRZ8P23QIPOKDDsdxG99++R5KLjFth+scTi59bdeUkq64XV5N38
OCzY6GkJf+UXZBmrIWmQk9RfyVmyAu0KsR45t6qQte+E1w274/TVz7h7g3jVFm7fLTRENAlcJOxm
qMe11dOc6D6+ObbWqOztw61W2JS459fiEJSqc+vTvbEjoITmobT3YTJj8JEbSteV7nc0PZl3GOD5
ukOsDxhVEMIUZZqprQrTnVx8r7abz5ViwcTtPJRySD6FXd3s5ZyNWaQA1+sn7ev+LIzn9+mHfSUb
5YpECp9c1CqW73xYFU96ESl/gSQ3AU0TkbgMQzyNZEaUIMrnL38nEeqSu75f6nCeT9Sc+nJ6BOb5
9PZFakHRmsDS1ao+3fHWBmZ7XIS7QhuYl+8QHDWQRZcUHxEqQevShyc6RQ8WbKZQWWW8ykjICcqe
jgDHI3p74pttpt3YVVYWWS9xQ7CRis3rKOZAvPSeIqiNeoqXr/OaduT7BXqsyL76Q04ZNxOPEQA7
3te8BytwtTN6jaCn/VWHxuWxB8mV0zEjeH5qiLoJEiNHhk8wTFkbgQ86zbQ2T6Ae2m3ryC4AlHh9
smnYO7L1ZghnoH6eRsGL8Klq9O2+CGaLTQQ/9X+VpLrfLhRGBjD+6NyxreyI7PHqUUMkTKgIDuZp
UpM9E2vKvF7dT02URMgf4ZxzNnzcMSfqMZ7nMivYMv5leorRCFDb8jHrSG/WwiM6OPkNH6wTwjG2
/QIzNRILaVZkGaQH+saFkMVfF9Bkjt1ZtsLgk0CMUJDNMdze/Wn+9eKmroVXjqwK5A0s0q3GL60j
hAt+naNCC3JhG2Gii0mThT9fwumG0r6tY0iBfFPS88u+Pt9IbpQZ/Y93O4nFOxiE5jRpeT0eN1B7
v/bVb0eaiDq3TL9fxi2EwA5Yqzh635HAuTMIxoTmrEUokYpIr6/yXJ4ACWaNa8L5xaffUSYFfBN+
WwO2Z6TZHKllKpwXBEX3+GnTCnThzBYQv+LkNwU3MeyqZuiNAuN4IIe2vQoJY1RldTZZelbTYCkL
U+XBLi4N32dQyWEGo0tS6APH3zr9A7dKYmCPvD8L16XaD7sjo+WM/s9zD0SvxyVRaH0RFyAbDzuO
vTrTg+CoKoR5APCxV42HBjRug6z6DP9gkHTZTdylGbBNZuG1FEzr+A6GsBG0Mg+w0Bbe+N9n1ZDS
y3+o7tb9wOXRlcDHznTtAUCQ07Uv/U4cU6Q8+A9cchs9RNGuENsXMfE+kWDqzlERBPPqNriRYaVo
DLfDB7J6w49y5pz5Lh9WsVKUFBU3uF43Qtv2u6Mwi8c7oE7WJMuVoSHDsTeytVP6rNBJMdTjMZUG
Rn/jAcCj50j7dthFEPEuQAhvIy3bDl2qv6uXaLLznvUrTFm6NHSz0aZXp88znqFmE9NXoZJsyD5e
YzBGBscBy1z91XWLiCmMfwc6ae6IQDyVl0zrrrmsneFvz9yzuWN+I72Uq4P+5/spGQxpJWvIg5LK
DfhzRFdu+XNpfcBso7mhPIHNGJLTixIq+xi0a/kODS6zvC4lqzEw8lYZ/ZCRmAzEYRdPM8JkdWOj
IYCMdbfe3olmyhogW1hxkH7vpwCDgF8jvLDXBGNWGTz77qJcNoY1Yc/FXqKdsbHUnz08CR5TEgNB
1LHG1FXLP10HOMNDwiNPNR6jgLbtZpVXLfOZGL8jfvcg6SaroeAsuecWa57tDasg3jz4XcQZKKDE
4GaJw7P7OM8mf+VUbVFqd1u0CDbCx0MV0xfNRwGFV/wiJIrxfrrxGQ+/TT6NbLjmZG5Ew8ztqvIP
6PDTPlTwnoeXwovgJ0Jh0nxWR3cee6VRTfD1bwDiSIq0erZuChdZ6zcurIYcsqpPhinoFk+rTZfK
1aNsAiyeynxgVs5UD+CmM6L2mXFpuiDdsC39QZr9elvh/rNutrl31VASNYc36VA4de7gQhePUxj5
dlgiEKMHiBwepKWbM/iinrUpJzr5H2LHVd9ESHas9qU13EkOznjcx5KyCbjahUpiMoiGehrqqpH6
JoxsVsmdq7HYEMmdRbknCColPUwtCpihuZZwEKVHT3nUfCxqUeFDkHOvFN0MtMt2U4CeuXtbQwvt
JjrHsAzgBzC5rRxNcksljlyx6mxIt8y4lrxTcGTksP/porUeJU5d7ssG3ZtVtdLo7V3SirOwpi+8
XblqsYwNk41tCKg3K/ixo8q7Hpo4JumDGaE6naC1wsTOkcizl+8lTgXEdy9I+IbdBtfBGmkaGQMS
m1KfFC7dSgtaCiDQdkDU+JOMAIxbaed8kzgF1w8MUZQqe4W4i4fELR5uA7ypfLPDBj7MmfsQSgHx
fCLSMusDHbH9Kc0lvi3vF9XzDVw4SNsatHcwyERrp8pK1TK/gHa+h2npFVQxg26I/7YGCQ1BwkPg
1yLKlM93mILCxQeFRQIeBdpW4G8TLBNrBkUySzNUvPrfGksm1vgR9OPQbNEryTJCi8ITQwp5gy82
ERh7JLtPtMc7oKWBxvId9txBeRBBAanhBCvjy8Gz3jtAWKrWRey5CN8bs5eU5YsPQfJLQXkWwOML
xDDoB/oK0PrPOqeFUI68zM3mk+3+fVb7JP3aAYfPbQGky3L2vyo2t5vISHIP9y9/dYUR1HPUYFWx
pPB7XueYazChcXBMyr9jvK93iObNOUhdGuWbltpJWIOWVVl4KnGgaeF7V6G6FDbe4PKhqpgWS4N+
yIuuCZDhm5klxx3KzLHcyN4B2DYtcW1z0K8xANEgi9OoAy8DWkca0/sQs4x/msMNXEfgNIEMKivK
d80dgxq9wbT8+DzkpVcEH2j7Zcp9n7nXfa+H+siwtpjsGMHd78VOKFahiaIOT4x0ukZwT6TVOdiN
K3C6gNsRlS8wl3oSKHcTMmZaTVRuCRN3K4ToEb2EcfGmkYdazTmU8PYQ66UH8vmwK+stfUlLk0hG
FQO286yvT5q5qCextxtJHR9SJNt9AvQCjPQXvlrKu+6CgwwBkszE1BOiKxQ+ezO9fivaGGMsv/X+
GnsNvuvx24TpqOivD95dXUb8shOcqOaIs/7Ylcpby4FEzIn/y0kpcUVU3rnsq3qy5SMy+UylNGOZ
47S8MmHdS5H0MnprS41QNMd4Ks+NlE+X6Qvsy8ZAmww6dG+DpQcGIUQEc2vHQsHAySh49OllVidd
dd3dY348v0T56szgF5iiwNciDNO04cw7v+Ac9iRiGH5YfEjGrbC79ie3dg4DOaKdOWy8ls8U8vaB
q8Li1pG5KTlXpj6Q5jZYB5HyvevixTxksgBAMxl+bjDmfpLlm1Si7NZz3seOwphTs41UtRHQY4Va
oF45xu1zxdCD4+hDBgKpQfjeqLe/i+sUGtFpt5evPdv+4H1NDQcZ3Ulfs2rg0U9MI3a81m8/oyiZ
UCkQbQupARa2JEJU5eocR066EX6TI6aNAt4IHl40/HcJqLzFAHorPJkrZ4fRg+eKQUOiakm8kryT
dACpPOgaOYGIDZWfXxrqJJs16GkjeIcH4x2f965vrV0CCoqPSpwYhHIozSVarhm7Aet0x8UdUvSU
awqcTQ/Tog9ReXRAveroEOVKXTlEwxfSW+iF9ZxWKnKNzO9nzS+RKTWkYkGpkF2GRQuF+6Td3hJa
E/hT9PDjA+Gw15nLzf+VsvfysNyGxrItRe6rZoiZOvZX97NKfE+wGmeoO1A8nMs6xqd2+p/HRZbU
87pNxBWyqHQV6gF354ZUyiiOja/0+7QyOHrV7sOEsMzU0r+pPBRpn0s6v7fPSJ3trSJO8p58Qi11
RD0VSeY8hW2b5MYo1itXGa1Bf036FL6gBoWQ75i6wKWRRX1oKJ18baH4cwDbENFwdQMq9wbg0B5Y
7npxDyFGejwTCSXvsdjPnTEXoC+A7N27Z0vvD+WOMm6ki11upFC+hpHQOvm+c26sItLOrcrHt8Yd
DecnZXLAtiRWm9shZZQfp23Wr7Y9pL7bjIspUBio2zu/EloI3+zrQcMiGQNpuR2lDlNF9HcyPZD0
aKgrabZkWwfSarxGTyCznorUrpnVMb8RKjw3A6fIvJ2yHEWSdd7B72gNaQ/U20WLYXOIO5EZzESJ
tAQC+0QnK0hasj16FtgSEL50ZkGzO9NGUUIamjrEBan+MKeH/IM8Wa2ty48XL47acD7Pi+qGhzsN
bvvjCkW5bqLT8YaIepvad8DaeoSxIaT+MZHET2ZJwEiixU824nG34egD7SvNljogrhPWyoPAJ2ig
JeUzlyYXjQRztWCS31mut5nTowuMrF6YgA1KtHXSa2HoNPvw6cdgW2oREV9JraJnERwlwoJ1ZVGR
taegQBQF7KBNml5HXLE/BWoXFPWLWYWqQRnEulrUsnJ2LMcgRtlbfuShHRxqpb0JccTKLrUN4Z7C
9h6JExhJQiS6r5DPLVEQ+Jl65dBPUsLa8qXKpjv6OQqz/09xiY+z2EKOdYph0Rl3AndyX1pCgCsK
yEHktvVzWT95n+qqehrqN0DfFoCX/aaF+DZ2w4EKKr2tzP7TMkbbPAnzdXY33Sa8AW5Mdg6dm9Gr
xBf8NvzxjVUczgpVqm2uDQYZzca3l9OvadfG7NQ4mwD4/4BW6dDIOK5OtotxELh4bHnLxWY/SikU
F+BGDZV7iuPDWF7whr1NFVkBKVbjSz5Bpx1FBmcmzlDHn7RP04hyMCFnr/2k33RUOs02CO/CBCj1
jV0FdNiEUo2x3YPRKX+mJwj2AX0VSnD52qibfJ4h5cNiXnhFTE16NmzqzVXABPesrdgMp06yUMO9
s3z4i2jND9ZDVsAgENMjplzmHwhCZfLGFwZ2spNDuclmxsQhRulsBNYhoKepMSViOBlscocKVkE/
UZcud8UyLlkEtkYh5FDzDL/b0t4zwazGRRU0kr/73AGvWll3PwRrJdiS+UU3ztDNO1iEowOcepWF
Rj/9D09RYkSKnhyE37Ia09yaBm2ih9WCmOMADrVbvLnuaXooULbaccud5ZsplTCcESLHO+8iF0ze
dX636Tu3AyPOF4zoOc1itxSl+7iDq38GdVg9ZyKra1z/VkaeKLKw0On0d8HWIWlFErgWGl93ncc3
XFXp+vgk6bMaUZtS9uUxoyyCsTm9ev05zDam1Y1KdxjmA59VqOXQFvpBV1jHQ3Eoi5hDvq5Zjbo0
7Tf10c/AT9rki4yuVYdh6TN+OUyC5DwyTxKlY8V0cDwW94y8wuj+HommRlDYfjXk1kUQjBQfPUjQ
gZ7aeQFmT+5fPu3zeCkJ5q7jk4XmztPmEUmIrbK1zNQvR6OU3p1MC6YJuNTp0ul9do6pB8kKaL8c
jZOHM95SAoTDlejRnGLjgso6iK+MfPUwllf98DJi1C4m0AiPsmQtzsZFlxoCqZLvtz/+iD0pnhdQ
HKJlhJIFyF3dnXXIWt00CyAKu6lQhasQ0ZOOC3kjthe8aQD8xV4xVKd9+wwXMcdBddMdZPDbnYq6
2Tz7VA8JCP3vtl0klZBBeDktg3EO0z1Ilher6oBdu/YtzV8xEc2jGENoIg7cQd2YkJHEjlMTGL8p
scVgd9hLZQxxWfuRoqeklACgSStHguLBDoS0r+smNhnpRX+hdpxwk5nEvnYxt+uSm4GlJCUo0RxQ
VlgErd0TNNsaG7rgxoppNz1ISGzaW+aI/vU7eqEzKu1sLmRKugAthhTWOKBx4W15KY7r9PoNbKGb
Bh7xa8fYyPTp7iWawv7+eLInI5Y+kRVtlSo676Gznp7c+nK+EgOSIP9hGgIGzAsDF5AELbyOjmgH
QkKnsY+y1GkdyBOHTflCCQXDt3qH9WGZvuDizdNPQlt6MzXqvbMAibe5/+B7vjsSMF4SsJ2VUpUh
qCXBLSL6pZwwyIcSaoOfgxvo4aPFAy8IF3hQhzCt4s0TB3lsmVVIdopQhx4UFjSYghUg//H1nA5y
h7QO1JWIscDja1bb7UqKhuvaLxWu6TuXAEVjim/QR5K+EsunmOLQ3J25YxNYyeBP5gP4xQI7UGRV
G+lrn/Wy5JlHeuF6Mgm+wcW66RBOWZclAoY8jIubAMoSuAqG0DAnTYg4r4FPS8Gb0i0ZK2bmEMon
uBOhPvRPhDSwQnpAPT8kMHF5iSOA43TJ4fwmOFboyfyOVyJQYLXDS0uYAlaWIOFhFJgxbMMBnl6V
93N9cwA+Zwilv2HB6ofg1pm+ar2j+HsFFo+5jo+HnRFi8fRFS+gdfbUCG73yJJEd6zuYhUujRl/u
pxZF5uagKUkQ2x1t7L1JZ/00Np/Poyf7Bj7wU5rw4IL3oV2fPRmUH/BumhYlJshD9Xonf5UXI8eW
85T00IOeqyzeNkCvN0iBmsNjIMvuGYt2Xf7YdPObWkEYNQOhTXcVvs+s5Y8Swgwc0JqfnR5kyvcl
0th7rStoEfuuceCAj2+sWddI/lPY1EaooaPLhG5QEpSAROrYKx+3U2o4UMTH4/4GCqnv3go/+qyw
ec/ZzFANdNCcNUjPI3ycvO7alvfpX2HCcSgdr4dM1NTT1GmaE/BIMARYfLkJse7IUGgY5KmhnTT5
5i1JmT5uhgbedeijEQcnzhMC8hLfJ/6qb6YPtQrY87iKvGuJ+frfL+0vJLHLWcKy764l6gmsc3ox
S/mC9u+/APV19EyoqFdpYgJ05ZodFyfXvGgP4WTke64Cpdwg1kDep6AP0NAPeI8fhyHhsQYBks2U
AnTf96oJ63ez35dgZCPTjYCSG3S7krVAkVt+rui+4rYMR29Z7SCQXyDTqRg0/Dt0ztoZDlU6yHE6
I7BXnSKE7uepeTx0jz5vJN0m5i5vFbi7oQCDnyhmDN7n8fTVLNRq0pDMTcHzX0kJVT4fqTBrT8Xn
6v7VLcBux3jIqGlgQ6eqiKNy6LZ/AT4YZKVgKSb+pYo7EPVcrk81yWTOHDYQZCm82C1VrQOrwjLZ
d09U/Ex6Sx3/7Zzm+fZbVX1sgATuYPAim/fu5FccBGKxuJ7mxUFgNsQluFOj6GUnhUwI7ojT0RDW
6LAoJ0q5jDmN/VW81LM9MEYen6agYaEH434ZLVxojXFqINERkhA4+StADYX1dZ+BSAERWpiTlteP
NRJOaw1QcEErHKPGMjC2la43eo6v1Nz2tjLAZqY3hld4/EcInvt1kbnaXKhY6Qytijzvfl2KkpDN
nQL7uh8cq+IaK4By/ypDiQZbhUW1jUsI3t+dbbnFlcenz+iTLi/IhHKBRHjRmTKqprcw8rPc6/Bf
rWZhqV/mNPqMvXCuFcfqcMCXjv5Sgy1ijVoVYnh+lHnfQWd6MhpoKFBHSj7zHX3NA+xbJh3nsm8d
IaPx9JUUUU8ED9ZVhPlCU9ePtwdFJC5r+6gckuaRmKSUCUjH6ZHCDPouOkuYxxP/InuZ1rvncIpA
YspitMFDfDZdYYYIZJC85EXTPL1Q7Te9YCXr3Qmq+MnJ9NgvYCda32uJDFSzbq4BXkJUjR9EMRg3
D0rgObY/xFKpFFVbKx0nmwb2XiEJYAu+8uFy7BwXDOIHfYfPlwhEBYJd2InyfNCsqostDSRee6wu
9Il7OPe/Fs/7w6fz2ht7nZPZiPFFtEUSohAm2v2gx6Z3taLRBrG5mhrOkbIYN4Lf+m9eZXPzZjFj
5S/bO18IkqLbMks5iKIjpoDasBXcszgCQIWv6ZMjP3kUF4ocKnAWsrZLw6scy8DCIgv4HbI3mgWR
Vqq2SBn5pAH31fd84sUAjC6qUEOCpvGjtBe4U9GKc89MhRcACzGJ6/jQpOwqQFhNjysDaRqSqo1S
neUDH5cuiQrxZ1lJXiIZluflfy86AvX+7x3I3cTLT6PSi6YksEWIauyFHm/lAzWAlN3p1W6GQaR3
durMn3ta4vuaJL3W2izfOglD4ux9LaUQOtxRTHxFS2jbGiiIKgaG1Cek+fLzdV11LSQzwvldCwL9
KcJe2jMxE8k1XAhD6OcK/i0ncGgyvBP9GGp6UNRGUl5Q0JR0YgDwAFGfp7Rr7YY0lR7rNYXSmBm2
7l2bxjGhTbp89PvKyKKF97G1ya7WH9YuwkrapYDCGKgJyjea4ZbpJgWGFkA8LwRRWHRxsBvKTqdq
7CXNHCVpCDVmgijaDGq2LP6eAHkWTxWIQ7DDfELQ4P3h2T+cu3TsENR1NATa1i+WGwb5UkMA6ZhH
HOfRjxVkkvJ6pbzWd2e616h3Vn0s69AyzoyUKr0ZSg+CKTidWxqnT3IbIxcbiD2M4WAsmLsyT6WJ
erMxaLqdgK0NotS3jZGvpFwrCla9hqRVmcfMjzqv6XY+sTUtp3MLQZpN+bfXBYIWQTzHPiHogIZ9
X1SOjRaQeV04AA3rDDgDCy2sS2Z4uacPxHgdR/H2Wo/n9sPRn05D2XrQSWR8f0x6oaqL5CddhSwU
bX6WSEYsm6ShpHPIi6Y7ZdND/pgUZBaD7pJXBLeHnIn60VahEeebFMpVDDu4ssIPGnCP/yE4D/Wg
b7vRlqTFKPcnyRczLPhYYh7G6Tnnft7PJXjDQ0O9l5RHwF6Bapt1zLRa58vxvGCxgsklcF1V6cGX
eKQxufTF8+rUMZ7yAbulaNK5DilCzGwKhbSfE2+odUGi63uDqk3I/seFiIriIEZGpOsl7QvOjzfj
0dTKC/aTqzIRAZionwn8ufPiwQIqJllGiGWa6FDdrt1R4gdp9r5zhv128SDaBrwyXs6lrlUgu1YG
teTUMal5VGB8t1pLkSnGZkPWAYM/rHw+B4xOQs+zhac0EH3UbrNl6mTIN6o2HdIc9/Dh/P8DYOLK
rVCIH6jFcxkhohzey1w+J5mcv6T7PGbHGuc8gd8qzm9Y12Q3YY9KgCLW5IZIUX6lDn5+ymkiIyf7
0dAhx03Cui9UXQOZaonzPCCdZLJkQHmR5neimIrJTIGxOMhbSeEoPGJ7j68iXFsbk8tFPCimMksD
Cj9VxoZeLsb7bJ0+tkM9h6vdeGzDmJ0IVTszZjSo2dmsvRkr6nR5Ad+4wUcH4/nLlf4KwHuX43Pg
foE4/wsplU/uZmPUCvjd9dJUcCuuKDHh1WjCv2sd2rbIvz2EuzRQtNg0vPTTyTxIJGJBxufAzkZu
eW+fHsU6jTiyRyoT+Dn9av98L1IosOLCuGYDDhhwwOcMqWoge+kJMf0p0BOXnV6hahbxx9qeQaIM
4ghC6XhySNUDi2f+DVBK/VqIVm9s7jjmVeXC1rZYdB+8aEqf+PsuHT/rfJVm1PzcLX59cqMWCzmW
dAhGCkzraqCxbN4M0FkN18qqmxrHrgFQ8LhTpGzwt6Im5X5C2R404f7GWL3iNGWzAZ/pApF7A0OG
Kvdo6OHqSvJe/vJia6bHAUTTIXc1NjocT+iwLSZa/MbeIHYfcDHXe11fmJmEhhzOXDxaJ8IB+vY4
U0hMzTYxePVWbK0dQRxun/EoUtnmSROTqPGpmEFeImFVDRhLxPq15xt/dID9WuYbpoM5JJf+Ri4i
cURHEj3b1o4KZdJ63xrC2/lBA21QA1mDWYKzKyHMtDzWEeA2yoJsxW7agcjAuJZXL0MLpuXUedx9
5xtVq8aMu7y0Vo2L12S8Uv/QpcBQMZZ/wCgyTJeC1fOVjTCu7O5/tftZjvF0dBJituF/psH8z7mn
W1r9qF3izxrzpaiOhZD287ylSrMox7rGzaHa+O6dsbl08AXf5kbaI7csHie1+nZie1hqQKwMSkAY
nkPw9DJ36vdcLWidtIT9ujKHpsfSyEZRJ6EIDD3llqHCvdlLyCor/nZi+MsGO1w4PG//ETxpcSRU
7efnlud+X2OYPulH55yfpmbqbjyM64YYz7PSrj4AWCLstwv7tAn5Vwf3+51meRhA0tMQuCfQlRX1
FjT25vlUkryDPxfEZY+T3Wz3hkswhA2fK1Ld0/9JnsYcU2Vm2Jw514rRRAR2861jcDAPiFxUbvge
Jfbw0/4ffyJnyBGucbNPWInVYpo8fklwIkQdiitA8439/TdnfzjjAFZnrcA7y09BCGHLaRrnClm+
32Z0GYlhNcGAzHgfadyjjfNCS5lcGDEfpvsY24RRJ0/SSWeBobGl/iiw1WQK5cvVEgFrneDNNGp/
AbQvAQGtzzOBB9GF4WilhDNbwdqZdICqEXlntBpUE+Me9EdBDP/weNEQqgsb8oRlyBRpb7FKW+EQ
jynYiHbA/Mr8FqzfWeYb75kvTBHzeNeoR+JbztDLXZWVC2hJ6d3whNHb0JVYLTjqr6sLZvYi01yE
4z87GWIernp1z3bwMNeyrWu5lKWxji1aja4LdPdfZGOGKy+YOTT2JmC2sX3tE/9WFOBkpEP4cOBt
UQp85WT7cTGgREd837ueZX8S0cne7KrZUDrn+8mxTGVALxdukzbnBhjeaT27ThS2phPRB5o5pMJk
FHQS3OTPusglGMxj+1QYTC0NtbezbNDEb/qxzFSembxaySUr+8Ps6fyTqPUPaBnVhtc9cs08sCsr
3i1vUQH3oAbTO+twX+gsrwmB88UFXhUoqUjMfj7VuEZUNLtM3heAiXXTrIAUwlFS8Elg+omSUpqc
1cG5XkF0wHc766Ct6PB9pV3rptLHN48wu5xjLwNiHKl2MI4QF4CM577asO8FgR2zAiQkhsq+wr14
1rt+gHOgZ/YIY9eXHlQB1QsgBhjwWNoVdrTbIXYeiL6i/q/LanPjhyM9LKDG+aQZMPYPK9Wov0+j
aO4pKaQc6x2nPzZVv/vhOYFAArFXsIUoxHgXIcmEw3xh0mewSESqB76XQT7/jX0eUcypKVlWmg00
fsLtMHlZzxdtqzWWkKO/oO3431FVLYIYkwcfWLNii2cdNRvJdYfWTa5rhcFk03EJaOB0QzNnjVmz
nKHe5U2qk4k6Q6bZ3nwXFckAZlCPc16nnlLXbHJxCvCNOTGyUpwwS5HrReAIWQoSpXF3BC8mBRx2
B32OMIInpr81X+tl40RVte3MZR0PjShUkjb6GbpxXvee4xm+PiiMsttn/He4g+IZ6tUfXaEskWxk
aUK4n9018+jkzfe3Oh0XqSfKexlYEKhhwC85K0khlP7CSLzDrUtIw7B3+E7UPY5mig1W4RFeuoCI
Cqod1iKMiWDGx5JrPD5Ozi02XqIW6KUYB3icFwsIHVVFtBdmSbBhi+DEEbMIYfA1yRrkdEFF8HC2
/njuzxJqCi4OXwycVC6nmMA7PwnfsnJVWHF+JAVBNRVRDmJL7WroPzl2YMD6JAWB5aLrgwqbg3fs
QZiyKFhMg/18QmvJgUKWx55rH7mhIdmub/997CM0jg6PfPg0n3DpM0B0qzZnCkKjndhf1pdLmtNO
wWpxcbSdcMzqLJbg57OzdP2Vp9AwtP8j/VVUd0DJCrm+gMDDxMRcA0Vd9JjxmpuCrByHLeKCykMc
5BqOcljBjG0UgP1laudJsVqnR+f4em5jopeNEnlGkM7+YyYhelB6nDfmUnhBN9HbRizK01TPVQAj
iKnQypeOTm0AmTDzAD1dbzkzjrfe8s7zHzjGipNt1h2LUxkFEoHFAZe1GU/Et/x2G7gxpy7pIl9S
LNvFNN9BvAOeoG5nVMK8lYOlNPsJ7G2b6LK2A0DCzNbBOaSFmQZ4/EQRgfjAL5tFxgwNjeOELxSk
jDrByaXoamRdu/bLM5QUUM2YAiG/LhocibLaOil/eW0xsj+0Qtm4C50IyZzjZsTLPPEk9G91Gyz5
5w44A3lkk5RcCXmFTqxMeNEv8erU3SV8KRKx7plZCsLHGMR8E/bqvNj4VDDx4MtSE5ASlz5jyUAx
yMBcQ6mkEZpiOuOUl4kj1kJfntzrVH0Mk1M5EKCsMIzQTJU9HHpMR15SpdegyQZr0gqy2FBxKC/M
Re9EUbTh+Yy3aE7rhTE/YtKVAPadIKZeD9SD7AZzZAKQoKqWDchc8143iW0uR+y7ktjGsnx5+Z+Z
ScMJmeSIhlvC9AFBSLbXUAwmHWc9/nVBwMi4JA90ZWfRuIKhqr11sd5DJJdwQq+XPd92/b1SJdC0
kuX3NS6IRVgktBH/1sG3YsdvZ+1TOTtggG6QaVZw5WWDsAFu4nSHLAjI0EOQV3ePghwPVhkNBksE
UbjI02wTjm7I7XnGmlD8OxRF1CMaS/nUSPWqkjW22geivmQP0BrRSugMSsaUh5IjUR0YIVJGVSvx
BJVZ1IwRE4Jn/pdIgtwcR7gCU/7P7lR7pAujvX3NDDNw+Tq3ucrlWJpcGh9rQ02hjwUR5a7SGkJ2
brWXutePHosXolqYxvt3htnlF4s7hS/RJBjJfAzmG8TuN1lzDhxqOwyyNtwzNnU2yewn2GJ0LqkI
vX+iXFSamQkhT+dvagSdz3iF05AK6vzo+nDDxhhliMykZl31GBe6lU33xybnKsKC9Xo64ySisxyH
DgBFUJy+22KBtPxvNh2iCGt1+22TP3fDML+mcMAmSlSowTlZ60ClYsZ18P2Ild6p53wOAucK04TM
hxTEMwlBaPBCklaAq7tOrcJqieGp61kSipAK5pMPlp1snu2egVG7jfVNd+qtUCMb6eWoYJDL9XF4
QFOY0Cri/wNyMR4I18i36FInSjbTYSA81N8fZTuTZ/8OgbXCtTsqayZl74PsLVhKxzdHP5c552wM
a1cUdQ3fvvh2OZ+VRvfC/aBwBcxj1fxKrgUzCgjzLAdpclJfSvjxpw5mIh6pELsqKspdVoua5zlp
7i1b72EwqFsi7hdi3qh5x4NBSz9kp0wUrBhryhpcysa84JS6sL2227aK0nKDsYzAoI7KXObJ02oa
GaIUIsDBxr+mWAdaYWZtecco1OF5CqFe22nAnBS6y5eS1srnWlQBAGEAj4+dgtS6eMklkbFkoG3T
xdTj0qDSrHeS1Ma3uvaFfSzrXCxbr/yie1k1idViaq55FDC9hQ6cWrTEzlw06Sn6k0iqyJMA65k6
qp17Ja/yd0P7qZgUSDDaGX6SG1Zi4rYXYSgTrf+g3vAS+/Br2lvRWoNDVd41JRb9MhwKdeFj9KC2
9XcDv6kFaYkMABEm1Ta65pTXCyYggos11Odwu8riLd3bfOToxMb0yR8+Az1nvFG16J2BjIXxWdFN
NGKKMAk0WqwwjIetUB/21YepNYToI1IhYg1wUlhcZanYqlHvEk2ezjsTRA1Sjwjm463jNntQV/z6
C8kVTb+M+gIepP3yPhjqTYvdf3KbR8vgQ44BonfMWNVpEDj4Gvk5ljIw8A/U4cStsYkzahuE9e8G
rs7U1o/c4U7nvVMO1UWU9ZQWuB3EVzkWS1OaTQhmTclU4gnQrkqK9ejkrjl/wECSlTk/1BMSJJ6d
VTyQfQbEPtRhTX74OCiDloG65nmjMoG8n54zkn6CQVSZSoj1OT2WC3pHPCAgvf53OCHGFwwNz0TY
Ayj/5+DUPaTXpg3HUgUcsbUnIf1Z0dbYXqCZIlDjYPUJSBVItI6Xx3r4NpYfnquOkETgX5GofOoQ
YwoFU5vHL/TOhjXyIFDR469LGi/TaDBubUy5y3X1Bt4UH4chteUn2YZccHtS7Q3P7ytkylnSUjo0
5m6WOdQD601QCBoKXUTGWZZqNvdg4OxHuumoWNt4RHvYZr63+/4mp2IBxGh4kCqGHD8ZQSRXlM9b
CuB5a8pFHtRuyfNd451KGd1DpBJ7GTECUocjTttuF9V5+2B3kqdiKF7VgEWYliTQ0HBbp6PxaqTl
sjWep+LExKp2rO/TDb2rVktY9cpJ99dcnhiIu2q45Ho7YaZUWEN0P1xyhmBunmmbmk12LA0qrdtm
rFrgU+EMh4WA9bu+51hRRreVb5jR5gHbXWnK3MSoQ/4z22tOTOpV7LKNA5/gvaLMFpMhfcvIgak2
eH+8n60hUKaB+yRvMMujK11nqIi1YNbX3eLZuZJw4P1qfFJc1OScFWJ83DIMeOaShHeDy+C+YIMh
exi1dz4AMuvKbiWAsQlZ2iEGjWXsG09l1T/4402aQFmPdl6iqJD6hvhQOGQRrTbMKF+beg/6FzPV
gp9H18Dne8naq/7JQGM0HPf8lrYfWd/ziR4G061XTjIfKyqJEHej+PZIZh2nqU0JRkx7osWyDQmD
B28m9wscvEJAYC6wEEpubUymxT/OkTElqVo8Bfbb9wE92AQi29PE9CZCsPjRC2Mnib9xylWH0cvw
D+nzFxOVwdC3MX5Z8cewBaOmZUXIe3be2cyDaBkbm0eebGX79RNpEKajH9z1CxxNof+rGtwZDHvY
1LVM5jg3+2b2Qw2jKUow8kdLOXawTz1+GmPg1BBtxhd8y6ahIY6nkVOxwdWje1vuTbQn0NN7zxPZ
4XzPhr8u6KDxa1Old7il6k20pUV5gYw07XqY5EBjSlsRJfKXjmgKSYluoLXI3DFBv3ChX2/uJt+0
j6MpMzMxQ3+JYHNYnyV8VLN5nSXtiWN+X9U6lvr1+o+CRzNFOYFoOnZnV5SXmZr4n9KpGZUE0yZz
vyQIA1insN8886MyJaTyrAMNOhpr0AUUQ15jg4+pR30IV3PIX/43H/9Dl3uV2O+ciKGzMAHiSHvt
MzW3eo5iM7YeHRmR5DcR/3bN4Gz2cSkNY/2WvUlVjopnN3Wlf7hiHlqZmxDaHghoyNyKk9cAiBP9
lDnBUhGY37sGh4QIwRnaIf8iYAu69WJLiX38hmaFXKXI3kcPho8hoPcPty5DN4H+7aMHhs29VIk2
7hUlfYcSuCOUUv8EHYCD92fgudPvj7kRrNbkZPscX2kHFM8yTbqXuKt+206RkOuI8/Pb8SUK3UdZ
dVtmFFrBeAvdX4rYotImROGCxEfF1BVbIdj6RRSIVRMHFc/dWwb1LCq/D1SUOFrGspen0tMb7jYE
PRgIiNS/Gj8pFSUSPDTaGJz4nYl9wba/Ag0dB4EwwhaeJt+GoKRkC4ojeFLea61CsAviUGpSr49a
j89lj3EFL6V7aTt8R/eSCiF7CX6LPqinkVkpEU5npKv3qG25CmaRkTWYMuHVo33DWBEUvTqxtWGy
LKVZ+QY2tZXp99TPQC1piAnzPvahbRJOoUCOOh6cxTFMSEauSMo+CzWKH2w6Mo97LjqgZ/dMWVxA
FAtQvMIwOfQZ6KPKeEoxyYx1nNaCFMyI8839xv3m1YS8CQw7RqMzEMT+J+7U7u0vFq6lzvLrIXuw
/r5C1QO/B7NPe9fWa52dABWCuGBegPjRAW2tQjOjaHTxM2ylSTO4A3pCjQzg2ydRawwJamegN/aw
iGpmGvN2FzwuMJZpndrQw3DCyESYgcKT1IWI0pr1bJW2ZQHtXLReaT24BsgGLQm9smfAEYLCwju8
yPBYVnxPm3DscD+OK/Tq3QedHoXnSzdVpsdwi3iAOtz86pHOnXg2+klqzzg8st8N6yH5pmKcX1x6
uhygCxCy90VwIlJiHN31gKiAvX5sVK6KYHsNHaRl7xUaozm4lO+pykTxwMBF+FQhBB4w36YshQ0L
/4vrI4lIItqL1XgcrGxO+ivArxLYHaholB3zHzRtTVSkWaJ2hg6e1Gn592DjW90kmCv2PqQe5pLa
QLlNk3VD6CwzTqX73/JDyRPQimwzkt81hLfBM0X2Ia2HkFLS0KnMblbbjzTstbHVr/4l0YZ5Ylo7
izvqNZfDqQ9780/1QoyNyjyIgFxvjHCeioOnQecInUuskbUMnKGnJFghs7bteo0Yk8WWY7K0KZbV
VQUS+Tb/wg4/BK/JwzVOLfdzi1aPU0HTTBnVM9SAxrfHKNQxvLSIQTn23jB6aXCE1XrdfYSn+1T2
9q4oXOajITyVxrpgLn5LCoXGVDlEsgrLZqkeeyYN335nZBlG+26ohoeMcUCJ9MKqc2MDqNTbHkIn
u7msgdgdG9G4070YlwY+hyezx0nxFexdPtsVQog/ubgZfO6oWhw3/yZ0dQXNvQH0arZB1W9n9ImY
B7gENohBWQDM5H1S6j1U5kmhA42qTkaBU4phBko0ftSux2FDkAYN7z+cafmR1TzE91OS7IkECMNU
9Xi175kzEp9RxQh68nOLcthweErH22+Sb2+I3HOy2bfKkJx4fnk6F6IW0pfgK6WKSmNNsHv+UF1/
2vfI5Ee+BfPcRn//HySlQ4S3b8wMqs673PMdZZBOj5WNl2L/7/hB3iMv0ZSWwXWLXDF1Qdd4VcHs
WZeOQQq24AnwU4DqvLGaRLXHCZIJ86k0di99q/4lqNGVpoY4CDJMIH38gVWfPfIacCdnQwrXSNPU
t+9NAV1aWT6dcqQwH2ko/w3MKUOVg6HuMc+NIS+cVFrD3jFoWEvaQQxrswcEmG/MFL80HKbsaTG9
v5xk5/pqs/D3sHba7fcVmP3DVKzfZZhwNZwMvf8kwCx7FdH76ZMRsIe6uNuwmmuVmPRZjNzxiJ18
PDH9DNM5oq0YJaKAKTc6QsOZFj4UbQev9aMua9MntBksC3B0j0KK99CfcJy6xbt4VxchaWJjcYiT
A0H2gI36QPQ9aJY+2XrDqCh7mNbf7cmnc36Io7CJiyGawC5HVlns/POYJ7LBoC8DmeoMdJYbAxf4
OGdop5vmgzAlY6YndKDJ8drLsmZBamL6U5fINRJ2+BvgdbN3SwQDHZ+/Jjk6ghNo6rTltRtI0j3J
J41vBZi4Okr9yYYwoHOnTAe4NadFFF+hD6esXda1IBMBUw2vDdkL7jkhP2tIukEZ8nuEGL/eq7lr
fR+b5tlLr/YvgccFwKhK9n3FtLTNqc6fWipLOe2wE2r89WRh9YnrPHzyW5eZ2aIDhFelT/EZd2Wd
5q1y4jX7eU3cqSlelJSErSEFSDd+L8qmcH6D/6r8I1gGCFvrx9Sq9QgNVQauGwWFxQr2GfcYzIe0
hrD3fyXZikQzDh1mB3oW7IVnMrByXqdXb5eIKUg1VOykXOy8Lph0lwmd+sdB3G1HXhYupYt8GXr/
9m8BBpE2bA5zHBsyPEp9SgYXoWIcz4GEw0CRAQmNUPDNlU/6Bo8kXEZqTQOy2GfONGOWU5q29SI7
OelHHzt4jMx1Nah4s3kAHCj6BVtorJNm8iniPL3KX9lcXt8Dw4QyrJQTvC+UErSJFyIcAeVhy1qB
5WDBzJC0GzKfHrXZixnc3ASPS8+O5rjuAu7vmrFYo7I7HWmJ9HFLRVuaJRGofsfnYvVL9Wm/bL2r
LoqzNChh9eEiufOE+OyHjIeobKE0OClmB+ggwMBFLMYZMLgyveJBr49sMpNak6PfmUqZlegplBMc
MAZPBVkUSrUM+2ZXzX5umh3vzeq0wRqmHbZM7a285uj1oZX7GE7BTxtqfXwgvd6WiA3uA9UzUqgX
d0nzgkMKBDFZ7yNBN/RODPHYotRBUYWPQbtVrN1oSVp9l5+H5ofy7kK/+/pUUpYzVrEuHRFDIzCY
AQkIot6dZAb1YQPGUuLkoAPTx1xeVf7ju8CfikxI+W2dlxIX7hFiLDsv4zYzaut3bx3n5IRx7PxK
uGzR3gcfMyNOplsze0glTd6qnZ4RHG21whaOQxQRJxDB89KCHKGdHBkHVQu9lUIErkaWaiTC8KJg
XyeRmyfR0Ea2CYwFtPyts07OaxdhGLL5Rk1aHk/NJ4UO6Qr6NnlUnSu5MyruPPLD2Ka114SsC9G0
IpTPnig4vHZJwMxI7nqGvfLuCe+7z3J3qVInkjAJE7p/wdMb6RDEICOV7fWklWYZrJUKVaGkePV7
9tM2u1mVI2eG5OenezT4/GUfHjXRQ/Pvg4arVhOPG62ez/mDPbw0shB8Q9FBYG+gllt8GNoB3L7d
q64I0hHdN8KqP/ttxF3Ne4fP2Av22FiFdTfdEIiMRpeWTbRlfs/VcH0Ebj5mnadmnnYgVKRMHq9A
Dvjo5ku6zGzBoF70AZxlN+otPO10AhGY3MLYQmRB1zFlwIRcmtrTrg9Q31OnhpSie7ixrVv25akB
V8ksw0JhOEnAmeoMeZis5eKdFxgOGcybmKvcnr9ihKbn/EGSp1iWaGzN/nmO+PURPiX2tLRCsm9K
XbwzRZ7QLa3t4awU8T/SA7CkQ7jj9340cDrqxv8/5dxjlzktzV/YQRZOKqbi9/LO/FejSlw/LznJ
OBzaX5MHjwVCEAoyMO50HgTn1xf1cwfzDiBkMYxuuq/5aa0+kYGU9Y0f3OY10XLmqC53FvYAdjsP
E9gBRQ4pTJkSo8DCd5OqHkvtZREVd1bYOpeHnyDV0wN+3iC2dYmIXfrX5SMArPFtd2rIS/KROB0S
NrJemr32VnEwenWIDUmdvuFKEyggRPvBZVfCRTJ3rhx3Ew5mvTexYqTpktgYH2hezu+tBH7fYykY
SfnNDj88eDVc7vll/mioJE4fxd1wueI1NBskI0JKn+BbtmHEYCQ+nCtHuM6crSC7tegO2lgWlUhT
CCYl0hzEQn51XyIVKAD8vQtlKQTamxqSCbS9lswdHx/EGM7yM1fxVzFxoOgCYz8GY2i8tDazmDBw
EzpSQEOS5BvisoC6N+q7mXtElloRVmcGPIgElHv/A094PL+kLzW66B1FTsrOT6+PAFqraoQyWWC3
NzxkMfysiwu0xINYEa58sXTPB7pB3lFJj8COJiSvzCNRrUSzTfdJggdiDty0VssFqI2oxkPqo3l7
xrwSaPEzs/gnTR6EdJ+bh9i8Bb0oBBYBPgxS7IHUgV6mYbGshAF+KTvuPskIJMx4SW5eTrrwkYBP
bnaoXSsluoEvDsiHFvmb0WI7qohulLNQxEZfjowSR6azqA4yXEge1Z7iyqgKm6W3kroFPuktQmd9
IjHW1xCQJYwFQ8Ol5xDSCF6PP361Y+/zaSFm9nQ31J7TWa3326a3IVCr5BBf7vfYE1aCWDXmtcxs
kdeBlZWOCbWp2fv6pGKtxNTikErs2Pg/lj95qFfBE/Z1IIoMzHoHgCKrtZiXLUCj2IrRbZ3Vkd0N
ffl1D0/HOCRbjjaoyIsmfBT20sp6Wv2ZbqZGTIsETT0KIlOhO7AK5aqzLTpeGF6pbncN74xlHDEK
HtU31nzS2wH02TWlRXBfcwovtj0/b6q057bwwdWVq6T+3WrIC/Ut+L8ZTV1VD+Q4aT3QLbTS9zM2
qYgZwW+SsK3QrgMB8w45QRbqslZbahCSOpzb3jSSkgVGmtmbceDe0QQK4hkoxbrmxjookbj0A5lr
VLjBrO5KUkqzkveGllQpJk6ae3pTz25XUjo13VI+fSFQh1DfaDqtLUwsD/2vjlNV1vdKzPHjPKqM
rgosgNdPWJkaZvDaO7m8oyIPgYYZDpkqTIcvE0OCfQ3jLHmGS8JKyvsk3TDS+WmcMZHoOEq0yZez
sZJBnW3s7zS4uBSAngxnnJkniSjxiHi2bq/O2rMnh4YjZBDZf1+lOW9G/z4JSUf9Hh8ANrGf5dxq
w/KcUp/bXr8PhI+ZO5+F9GzWvnCzuwmMbkGSt9NkOA7MvTSAylcoh0YIOdFYBIq0zB/T0q6PD84/
e0BW/AK4jr683k/LYhWpPnOFXrXvW6GKpOE+f98sLLQ9XbjQouCpPCiXKX/5eMrj4DXcGxAbz2Z9
/yW/WS6/3oP+8wfTtDxDf0M8uXeAChdgK+Dgt6TjlvrPEYAup4n7svDlu59tdQn26JsKxf6KtI71
gfXGC+XA3HFJIowodyRIprCZh3ajaiC+lgoUJvuPp0sCRoxZJJLM9M3LKgmbL6IioJcejmPLlIAO
i7/NejY5MqV6rdXqNUuzL8imgpAAa5SK0DaWP5DH4T4N55s9dD9U5w6odrMRJyHEXwDwOfPdwbY+
r17thTJLsjscBW43frw2jERlR4M0y6q13dnWa9rCoaQeQIHqAPmel80ex7a9jNXCTIhxRKfanJzU
x8Kk93Jzs7Eo1xLqL+2qanZk4NC8xzpUXl+hp4lcTASkwVxdJ9/X7iqT/9hm1R+q8M+C0k8THXfR
pMeUkvPpt6im0QegLMMKTSJic7NanlMOt/8c1lKk1o/ueXB06PaojXVwY2G91wtYU+5P18cu/v6o
ApC3ct1C6JrMEGuTNSEsD1yCzkXxMzQE81cjpQS7yJwkPum0UBED3o3XzcUnm8E+dsp4Hsq0i7PH
MD9HCcH6aCWnl21aFfjCj30GccSiKkqvH7hsVIj/3pRSvR2DC04S4L9cl8ocI+H25oGoGEkEU+8D
AGttsjEcF8565GhTo2pQPyyFfQlfp5vDtkgkRoLDchWv7/iH4g4dzyTPKb1c3Rbtlhn52ToYttp0
xLcnCRAnovLYGtTlbeNBNfHyhLIHbeGthhC3F9Zx6b3n6Bdphd2zjSI6kiVF6tMDdutzIvCOLRnj
cVbtuhZJII+o5+HgeQ31frs5CgpRYuJJQbp+6E8pGNNVPgFiFZIulYuINMIqL2NpS+c1A1IdK+dt
8K2FxscdXCbJEYZy0mn1fDSUWF27SF069kMu4F4F2TO4nAFeTCZi1iH56xBgrTCR2+E8XH3pVpO5
b6DPEMBH+gcoSRaZZGn9rq4QBAj90aRT3u7inWvaYraocP9BaNnNVPQmS2Dje2jdliDKmw1v9CL0
xBDvDhCoiNG+HlI0O+8g02OmpZ2SALUGAe0KaICVPellxinCZ3SqtYODOgi17VnMHq7+ffdD5Z7P
2Ep6vJc1yFAJlipiIuqBsC36BHlgDgEG63ZPb1+UUFOEkQq1sEbyWy32PlcskgCjFwDxApeg9Qrp
gMcMyRFIvVloKMKgvyZFvCoTliBiuanfZZj7qMIONRF5CFEbf9yfqEQi1EoyUN5X9JRc4RykDOhV
k/nRQnNuQpzxrsiHuS20qTItbTGu9eeqnpCAtRKB7eooMshZGJhT4mpfF5WbzFg9wgM2ydTim1ex
+y3HaT79lL8eaPU80bfenCg5g14pdxQxP3swBvzZSWucxJfJoIcAb29nr9EPBw5cz3eKJXtpHvvo
3AKG2345oaJP2HTC6t94vE8aay03OUSjulm3kPWzNrb0SAdr7HAhg5I35CW2HQcGktT3K1pO0K7X
LQ/WqE4tnmvtFlG99LpSQP97Ll/lrA4QKLkc3R1ePp2RIird5xNku6upmLKxaR2dsSK7BxAhMIYx
59uR6qPCzxetStrwsgHvCXiAPmaHyjBZrKsw01LSABwAhiOsKacq6LnD8N5IJsDUF6GBkt60QD/x
fRk32XIrNi5RPvkIQ9HihqqoE9oSc6vEl5Rvw57WqCnkPilggUrPsip5O1syLg1XtjxU0P/jEYeF
+3DDsYagjQPRMuBsi6lxhMtT/X/COKkjSZZ/mk+ubIluI6g4rW+Z/jo1aY3HVpxe8lf6DbWACDT0
byi+ftdT57qBna7uEk+nJn2D74Hac4ahQAzJU2oQYdZMSFy/yw89lMoKBL+rYqS8a+r2BMkUV03c
qzOQSokoLMKXDn7/gF6OXPzhkOzu9+LN6RwTin/CKyI3a94wFOTDbY2RvMOvlTC8NRc+n7qgQ1TP
lKrALvhBOh0qgwhEnMR78o1uEUp3xvXQQh1nEvAneDF26bQbSvdPIyFs7YiIa+ehLeZ5ydiAgv7W
0Sjur/m7r8ye3/e/uHnisfCiSRwndviWxRjCVhjIJW6tij+j/CP2tANhD1FNOl7aNlxkHgDMqgTl
gV3NlG9MAg596HxCeIZccZ6kwNPk6qUbJ8i+8msYCbH5EGQ3UXX4GSbJeknOrJSnthLNU9HLp/Da
A2Qv7tyjnu3/jBjrihPhLcVvIjwVdit6fzrktAWAmZJwhoLTRSBjOdOEvNcFX3p5jLT1Amd7Z9Za
02b7cWBO5p8TOxL6aDYEgmMFlCgSFs5Nji4w890G6noYvp3u6jueTq8fjAnnnba+X3eLgI3li3cw
kPA0wWb4c3K35X+nK+7WI30unud0N3VusG+lNfMFUKiu9onikVULpLYDE6mIAmZQrj4t3NHFlONv
k39wq/nfg+7R0Sar0sa4TIgKm5cYdKsmst06yfsuF+/f/GlrJqWOqvQdOu5rBPtNPPgxMUJQevx1
9ZBx+U0kE1aCrZ4a3gJDZ1LW/eKgHHJmbo5oweU9nG3S0f6fh4zGPnJ1JeNNzPd/38xQOWE5OySB
H4R7d0bR8D9MtY3SkgoSJ+hcahKnItZP0n5R8B9bcIn+crZIrWtHQs00E/2AY7+pTjoh/3w2CWpR
9OxVrdw/dNU8eOKl1zLShc2GSpeBGNVXQ0cwIEgaxSOHgVgyP+3c5WbORyZqZW9GjjTAkNdEvbC9
MKkh3ajQ9SkT1rB4K0azCiyDAqaR9asAGEpFyy+ZT4fAt1/CzTxP59SO0J4DqroVdSlj7wbBtfp8
fV/aXqF/gb9eD9ir7oXQnSH4yUFs6EA+nDahxcIf2/1glrwOiDIZ+Pwwgvhu/5/hHVW/hPRoSHtN
foSvPr6weELhy/ugAv2Guzvz34uDjOrPyVm7fcZ0aMVA7mdTg8rvFsj2ey+VUqM1opveNDVKW9V5
oTob6+86MH9ZnFzW9q9ZAUkzcMdzVvkyKIw/IwFFie6TPz6G8x8Zgi/oj+VOgQJhJiYPpLxNLBnJ
hzkabC+2BpG6ER+ZWp1Z/ql3U1ICqgT3i5pKIjjdvNTJmNgTUrU0A+ZFmX7naCtac5eZxDgIWOtR
ik2AwfcTovn5BjjJawuQKICZA1qN0UuAzQTHpLWEpLe5a72xrITd+KzvN0oh/hLvIj8uvGiLoEvZ
FIA+DCsZ2VG8vnw5F98PUmq7MFZuQE0lAt1gtt/oj/76E7qGnxdvDYuz9w6oBhpKoMZK2o5ROIVS
MJfkvkSSZriQ3ceYr/wzyvpTP+G/NHLV9oEJ3az89NFT+e/g6lof2jNhH+21GNRpWs19NSTP8KON
VKKUrXYodvcXMPhH9ZuU7F1uvc5oQ87yNB1Ze8pZC5tqvl5vtj99asRykhHYfmFrCpr9zWji48Yy
aWMNyGjX7GBo8ZL6TsVSnJm0dzzE4+6C6wZ5JWZ/0p3/zwmj8uy+oVDlcv0pxYfoK4qnKQQHcALF
tuMh5UrUfKgYT4ClqogPZLLhXng5287o/LSExEwi8H8IwMULKSmjqN1OqfkW9HSDQ4GJAVPt5K2J
KYou8E9lOC6vJvpU4Fo19eMYjWxhXN3cgFZTdDo62wbErLdYcPZYnARuOhrlIlykzqlE846xFKSd
VVlPRJwvXBm4pp3bCIFgy+FrPsGqYIM2h3cAEKHrlWYa+jzMSO08gPV/AJLjkOBlu8ZPwnH2uLsP
tsE/OBXivXJqyQ4d6CC4O5BSIrphcPVubO6VKnc5yGKcQqgInT3s9Q4ghI8Z2CJv5F9Mh87uSAUD
BIMaJ7F7M4OMgKROJkzxX91ywSE8Lku2+/F7QBEbGDrqKANNTr3HOJLqs0EBg1x7Kh/a5rngrJhA
QihLVvvOib/UhpjB+ebs703PE0oWp0IsKHp1RIY76t52oVuQzI4pxcG4EDnVy9a8ILV+9lEa2S0I
8N/HbAWoaIYeQfR7AKmDQOQLam8Gq9jpBbMGWz9HBqAqhfPuAYJpreHisLXLptLGzd0PKoMG2/bb
AReXqu07IKfkCeK6rnbBiNybEm5iGKQKoehMBmGunfP883lauKA5FHm7UpapBjzHX67mTRq1+azm
ARNnlUgmil2lBM9/YU+HXDPT6Rytem5jXQvY312uym3otUtg4RZAz0vVzMR6yBHmVG2R0pGpbCJk
t8P1EDDM+GRXFl1ScBtd+zp7YkV5x4EviN2cqcaYHn24pciT2772rXxJpa18vhhoxDl1IfyJBkyR
ISvTCOcYR+UzKV4TD3C0mQtp4pA6lqORQaNRhedCQcL+N30Mvj8FHC1CtKNAKwbUWjVhCxKsidaH
h2d4mHVA/yQKlH2jUH1pbhCHgL+r6Rr0fhpexUjcZVj+doVjl8vLdEAXfCUyH1Qtdin44ZCDrLha
hSyernBJSdyxdpFk4VGbF/+kNyPjvmuVSJwhWW3ibfsgx1/SblM0AwJ6tI8yq+5auM+QDZDNLYiW
Ghc4IRTb8UppOpzVneQQ7/qi4NEdecR9n/dp1zQ2C19b0BxL80WPnjzb6QWArlU11sNGAtdhCsAB
6NcYszKtY955o0QLiVpwvVIXb9f+tacoumlVqckBytDZTaQzWoUXtbsHaz3Jh4oX72E0GkzaWl8P
wUWFFRcdDp7CuKslyvQflMkZ0QTJVVBXQCELJrKBsGSwbemnDBKPq61bxT9qQSOT5/cmebmkhv9/
qyvulIJmJ6YNAsd+qhFQpSJU/ZonRv2DTnXaShE/3TurrzJPVB+JwVrmu0/ggJnLRNiwqJJwqXDt
iceIIypIqosECnQ44h696OD2SM9A9/OUTYyCHdvKN+BmVQx1Ji2IW8I4kCWe+btgq7iLfhAxTnOW
6YN9i6zksj7o4DP7FGtd2P5TexnA5nuIcLCIm36D4xdQTc3+kv1H2YjciD6C1E6bi/a7lVKF7wuP
wyt6Ajzn7JA9ZQDdf/LibjMCa16pzoF4i+HgbsIp5gJoafF6PxQF0/idq1W3FopBCuMENF0UZDC0
S/xO2CVT+Wvn8jA4JAAq8ezLi6zlKYMYyQP02Wzx0i8o0iSeEAs70rzSEITP6RXRKy/f7wGYSW8A
fi+1SWNoD8Y0YRGdsEH4VnvpjIOBfKh55nQrQ4MiFU5e9GS6HTOGjD9ZlUSLViwTqkNkL7lPi9Wf
HR9Fq+WSllEZJZC0vi0jcdVTOczc4a1oGebeReKbSr5eipojk+C2Jekq0MJgrMns7yadrmrEvtaW
UdT7vLXfKD/SVIwtxclbS6v6Od60ihfNKEX3M/shUv2RIdlo6Eh3uZ0a7DEr51Wc+pcPNhlCWmxa
fPjbVA1sTL0HHZYTpqAfzZVMkdMY1JYZYaLGE9UKjxx3CGelioL/QWSuYisS+Tbr62chjbIoeWvj
ctMg8NEynyV0J6SO71wtS2NfWqjTmGG+VRVk+zLkbRVgDoBpAY5H7NjY1A/fS1G27uLhgcNr5CCy
573EplFl+jX+BhH6xr0CLBaJaSZM7noFtTUkFInI8LYvgW3FV89yYyqoB8f6iAE21NpF949Uphbt
ySKp9d/n717JD/0ZyjnCWoHSXgsd78adrc4r0T2WoV7iKhdY40QITcdNz68hZMq4TFZLST96FcBD
Ug30DqhDNxs9RvMDDCRTQg55wEtchojihizSTUuBrSvEk+qZ0xy1A55wTV10E+PjlXj30BINlNZ2
utX3HV3H65QngF/c8XI+jhJb9facYTavTD9eJu3W24xjHPni3NV6jb4TxtLaYNCBUQzp4Q5Gn9fE
gfpB5Glt7xoMhkvXMPX/EgWCGo12B2xV6q9tEiZDoo3DGrlgm6jcHgrCeGHggdwICT3R4k3PINKh
07ybhmTuv0y48VhvteXh4G6NsziEMR+W3QbUDNa5S9vwYgIoPmiWHfzERXJx+fcC1qZNkRfK3Rcc
ymdIKg2WEqC0XLIl2opVfAKDrspkEhBn/PO77GUqiFnLgO6mfovaRexCenjH6cp0nX+jYs6+Aytl
8Cf/wnmphkfpmLpkjvU/O7ywg1ykZa8Fj4vcKIRvdh6HP+KZTGDeuzglowU8TrLGq8ffrJWEChdx
gpXSNfHT2qzZZjWkNoGkDy0Lf6bRED0hlc6tBJLt5cAJkMbF/MfcJKQ2ivin0YdFWylcSVMizaRk
ofMXP5h501GxBllz50SU0dR1GMLKHaJkd2o2PBaeYiqmBPvlrzoSyzq6Q046Wml9rehXOFjNugfO
Yg90FFxjL9e1lu8hN4m9ZtuwIbndeHNGUGFI6hP36XbB8Pl/rK48bd8I3jHkZoSFAIRYuErojWml
/MOAH9WxFuZ5y+BoX87nVOabW/6VKc//KoeVsru0y/UNrXLSIE4AAYnT/weIle7LlRuZqtbG5U8k
Cp7EsOZ2c6iJdI/u+ICaJa4ut2BfwU0xqi0ALMCV+EBYAUz/OOcEW5/61rzZSQK17fN8zXc0akJU
PDmzgCxkeC5SCrWAZzJlmSawzq1axiKpuCOLe1U6I1ZlJ4zXDNcOTuDzznb2UyDvgmSIp35yVLWV
Pa9UNtXYmDHueUj8/vE8UyEj8IdFkU5IKvKUK+Ev0chp2NtDcFq+b6/RGTAXLG+/SjCTOqXfKjd9
21EoJRfvepBpo+Pq1J5mn77DkVV3LxYr2EQh1xtoVwWbJzVeNf7CP2CLGISPf00kCESFZ6yrfHKy
+yO74KATnaDfUSF/x4JnwV6EG+MSagfK4VdPnrl9oazLXUxvc4fae71airurX7OonzUj3EuoZAfr
CuPyHeXQU8WTJIhXwVlaFP/xgcEGpjsAT6WEi/I4jOhGPXv3UaoBghbFzKx0dgfgZhAv4L7ekPiv
VeH7kzr3wH8xLmngX7SSiEUKEs8HR2jytgR5g9C+NOdcKmqvN2ZT81gJCV9692JbOIT4XLsy3Eov
6Z1bUlqfVTNc4Uy+bO3ZwJhqauxWCZdKzFVFUY28p8lsrGkGfH9MAh+WMKC1sA5OwFXVUbQndRWJ
T9AoAjgWgxiLgGGW4YJmth7ZczbZpausmMoW0As1KPoZqVfTeZE+uqAZ/iI8eP5Z5hMlqqnCXu49
HgsRG6LY8DQuy4diDnw2w4QM1W/cpoDpuPGchpxjRYzrkHbpMmIBKGXK3a1DsIN3tFb+9pXBRYbx
3G6zKzj5cuY+FwlkvSRtzE4/oVdE7X9O+WpVemIqjhb7S4kPtH3twqP/dCrPR7BtGGj3hZ+fkAQ9
JAeJaw0pfXp0Sxy1KBb0v5Y+PfuigUeSGcQtbN4lkHIA+v3tiL9LdPOH0vvLC73uYIRXWsjwRoht
YL0JGgddDIclz7wIePmbFP/bKOBA7Uh1W/X40afMa+3yrtaZWgUpk0463f1oIZkuUsclLh/RnqGS
roQZSTw2s2jyjHEgHkS7qfzG8TCWVjKa3um5JcE6+UzwF9hRkhm9S4Q+/AeIQAoHUTbI7WL5n+yc
gFPE2DSPYZZtJb3EzFkhpTiE60GLA7h/zvPoBxeehAMnHCmgVPLA12idGqnufBf+PMgfOLPPLrVI
sc2LUtr8jGwOwHPHYfp3kChrOOMxYQj5dgcmmgYvGW+Tb31BZW8Os51COivPXRcsHlAEbwwoVbmS
4iswqmqMa2nUzapujVVHdd3LFSsuoDeKPFxy6YFDFM6BYOWO5XqTdqDDD/xCXfT1zIzM+F8WZ00C
7KtLk94IIBUPES8dXus85zzwssHyl2z0qNZLnNSD1VE0ogQZaxXK/mBbGf31CFeXjDQMGr299AP6
x9jH0nqNQlXi4IECg3ozGiSjVsO5qd6Ma0E975VB8taFhcUJPiuHPjwXQhRf8gULy56ff99hcsv0
2+/49SVU4TeBFJIOIiBbnveAtAFRvemSmXazdzSvdY9sjWmTBPbaRoNGlz1Y9UFln6CPoMdujexX
Hjp6dxA8MWxnaSyf5jmZzfflv82CGT2bWivc//UxXJZ8MhA0xNiFtd0gPwH+PTM7LYQfIm3L269t
WkDyv4vsYpXIcsNIgtYjRSl1mUmZvfEcS5AG+wUGDxQ1eGzQXJRXEAm7pbjmOKS2FUTkeOn0kG4o
SSYgLQBgGdl2r/+2kJoijzRfRlqV0sv9RNQrNsH92WUMIIUH7533wbQczu2QdqO9Gyoe223Izub1
CYX0VP3u7blLQGusMHIrYfQnMJhr489exjWhsTRKadk46utGOH+d+owdpZCaxGLTaMEEsq/V+pZP
13sH+uN6/RHkVIraUjT+bpigCBf0ghN8QAjvtXqpErLU0Q7vsRHl0y7tUgxexXlwMCVpbvgqK3S8
Of+oeGegfC6gweX6ezptqDGhnBR7s6qQQcAvgTW+8eyq1AmsJJiE3MfMqWUjW5Ksjp073wmBSAe4
z6vdHjLGvBJDV8zlPmXfvo4EyAegpMCLdK1yrLYgG3zB8dJc5KgQ7cJM8DMUV2HvQjNrSgPFMMxM
72idqYO14uUl5ISuVtA5+t6z1wuBCNtqSi643Q2AT8SRX0yK0MWQjcSa/kZykCoeTC3S8Q2vKSRs
b7voD7HDNTyGtjmu5S5vzCL6t32zexBmTVpw98CSJBt6iEamQL3Rp7FGxISfGf3lbuK+9NpdwccY
CUr1lGdTNZKgU3kMrEyT5PFvP02koXxxnHAvb8nunAc1uONkcySysSTvSGFd1VnG6NyIiBe2K1X2
8OnzwTFKCUfa5fYllbuFFME/BNp4c0ekAbxe/TUOruEAm3VYsU4uf1wvdET8j46qX4aw0ti1SmRy
CL/KlZeWujlivllhr/gDt7One+Wv8C4kb9Or5Wuwj3bYlT45FOxmHIJYkvRiRCefj4Pno8M4qo0a
Mg1AyylCIf0Br04zlsmJPK+t+j2udyApb8+UtyTf0pEKtCBG/EX9jG8OezEKkaQDzECsObWtnFTC
IGV0ZV4DzAsvUtsmsjBJnLdMu18eLzn+nsLBzYfCK+Pnh29MD8QiiTiyDVOqGBH7qnUhpDMBPlrx
CKfYSliy5S3fosl4PgXx8n20464YNnfezRqY0oSusL7fKDTr9rQ4bKWKSKHAAzK1plQaI19zy33Z
GgNbHy7LGpRHV/4hQgm+NgFDNOil2FMNcu/N6knutBm0PhPNldyZe99yni3lVXtWnXlWfMbzst0l
eXT97MMuDHEpUVyoKb3mdEZwrercDHuhfCHcDx1RlD9fsO2tExbKAn7uIm5doSUAN47upqkqJDDJ
yhEFW2lCHfOBHvMj68S3kbTc9caBVmHmBZ2waVVVj8oKlyemqXg5SfTayQIb0mciZqr08nwIQoIZ
UvJolpXQ69q5LGCs3ZUqh9dmJm9hexsQjTj5Yfa99KtAg3U6OYSq0JWgSPUrir1EBQeppP1Tqtvu
6McEcRSntRgUyqFCLRCztvQE9+vO2FCwaNxdwBrR4/YyBHOvpiDu3+JZg8FIfV8sotxOtcGLlhcl
fAJoQ49sVuTksbVYKEGrh45O0vRwRZ2wnI3FolGY+sjp/9wrUE9yZBEg5LjxhqCqWZNVkvd1ai+t
cJPo6J0zA+3RABmRPof1Kmd4/wf+BdN1smxmVe+BoCvFcAurYJohX0OZTFqJNiYPGH5Y3jn6QhSo
ocHJ5tr4obSjvvKWerF6ReauIULGRUJgxkoZrrg6h7H1eILOHZSA5qwpOZ4miRPSgLjwLRIaDBTi
ZUqUZnb4FBLJdq6cKpgAenDR1I1Xy/otgOp8fPvpMsgHbg5H8wgQitYCp5Qd4EjE0Bpx5hK7C1iT
GKm92BeFOT7iw9hzwVI8BIgFUA8VHbAeiVE0oYqRLpGkVVdnzEXe3sCpFqe7x8OX00OcFkc/5OHj
YNPjrO6dTCHAnflkmu37z8gC1xMRi+B7kaZTpOIlT5pMy4kikNZkVsROtyFpMAt97KfgTupyOhwv
gGG/3wXKZdjk4eqUFGIKzJAdUtt+0ynRUfojFwaqt4AwdS5OEH8Wa8Mpc9Rm7nYkTyGeaeCM+OXH
l9oeRikFTTt2Mka6AMeTlT0mQlF1E7GWO+iO97A+F7JicaFbqTEq+GbBQvD8FFXut8GtGkF0/pG+
9AAHJvq3DhUCHtpSXIjlQwICZmjMF0dl5IFp9otDvY41I4IAvuxcjngAzggLNvnDW7DvQf01WSxC
h++mBw4VNcU5rZRFWhbW2PgTFwIBPxFl7RbuU89cHkVoAzJBgRqmpAQ4UxMksUheVfB4iNJkDoMh
+0m9BFNDj6iyNBboCseNN3bhAoLyrLE1ZJE3sE774hoTpoW1luhCaCMDnal371jLTe3b8C1nYjO4
Xp6qs0t27XyYXy4LGQWinwRj1NJt6lwGYwzvwy6hnE2GdQmIKPTLTwvthSLS7PJsvEl72tlYE8FE
6Nw7H6/54Ijn8RJue/esVGVi/qFdjiteBTR3EwOvsynQVU1JfXnTCFxbkNdnIdHmpZ1nXbj2uUXa
9YuPBEdtyJD4kBPpHGPCTIJA8B5P9WmWmE2A99YC6sOBrlgpqTXRZf0fNkMokQn56o5y0TUw6aqQ
XyCq7yFkykShIA1fwT6batTYvPMDgQw/3cdPnm4gC4Ydvi+Yi+8w8ZxbZYxbCkazU62BdqtnK4lq
g3wiE33x93XTKiBNzr1O0yFzfd3VcE+hBAuIEdFr+iP0zVuJfrEaJTXmMGsM1gemblxhxbgIpM7i
ZHAAZ67OYnvyJ6577yMer/ACj67TzftWFcIS8bmh3HJSa0hrS6cSSYC9SEtYVaPMOA4RFEp2V4GF
4qYQ+I7+GX5wD+77VfggxOq8Lo+ejnW34BhIcG6Xv3PaKAoUKy6SS3D2OERnxAFYi9Ul+hfrhjgy
3r/Yb0kP48yvnt+VYhQhlqv+GWzvJPDNGaONCq//ql84dTYzCjhEkn2MEe7Omx8jbwie4aGUfzQ2
SRlz9ZLXpTUOsb64rJOPt9p42yu0f9sFKnHh6BfRsjGRhfmt+K5mkEcGnTzAWt04bxv/OCqg0fRu
LDqiftt/ZNRA5v4Ck/899SXDBkaMmh4Sqf+9x/69KB9xJM1IMc4f8T8OyMn9Ql1fndvVxigUdlh8
uX5/1V+GEw1dg4zyWIXA8TD7Tdi1hseg9IIzaaVncILXo3VH0kcGnkY/G+Aoz9C8WlYs9LbMTg9E
5WNZ8IRqfNZUx89LiT4Sx0tY9PgfDOcW8iYqZBF7IJtiHtOhbIgyKnmY3jGKLTvpB1CGSwx22aHw
gAkzWvULTeh8cSc+ccFceAmyENorcTFUo6imYg0slpKw92cio0u3Blq7W9f3Vsrs+J8xcpBJxKhk
6WiHJM+7ByJJDmWVQ/YAYwzcjw8dYOovGxTufA7BYjF7zVYaixtHBHG2pBDi4FlDLJckTidk1+sK
AFyQdLLWyisKf82jPVxoPw/oiD9xlCOze5D5DWZKFRTiELIdLlgRkkBarc62lDVrMOKSed4AWFXW
aLyrFzCUWUnAsqbHHnhwi//dA0H1RbbT0wqN0jcQE7N1x/E8TuDEp/HW+OCYeU+QYVD1Q73W14j3
ez836991jLuxrrX8amFCCVkhkal1IAJvrCgsEvifKkd8/ZW9R2BMJL8DVjtfiee/jywoKZazMpTM
mDU5N6QAhaZ33exWQyAsC8dV1a4RSAnpDcAU7viB3bmozXTx9nzolxyxJ70+rwLKvSyZofXALvYN
WYr95hNAToLFKj6RwiIRgzI3SSl4HyZl6xnsimoIG8sC+sBdxrlKXQO1Y1njIIjAn4tOJgoOxRvQ
EZLd+pE+UaDwdczapWqwbHfjX8Xy7BkoGh4PtrSCzLQWBjstA6kHqZFn9ADkMBTV+QNpzUBmJV77
BUecGvc9DMXYZYiB7oTyo1ImmHARioQvRGQoCHiH7dTN0PTwuaeJAuNhLf9NOecNOYkbGCYYk+TH
4vZaMIBNEjTGKUsYpfpTAH+G+yaPz4vCScSYKSY4EN2RCO7SLLY/mDBrWYL+ZskCAlmRe0ha+Goj
QXVrr00xSionY5IDeXtkv+nekkSJGNTLab+Mck55+PuH0zkwk1TFp+r+TIy4BW7eI5Q7RmzP9g50
L4FIuUsxS5noYfqANGuSqYBhtpyjPKaMc8Yn1V+yt9uLtCmXrAQ4nRmZiegl3CQfuAe3AoPqfmhh
8t/u0TD4L/cdsrKXInhEWiojKcheVrUNKti/Jxr50wvqX5MRH0Z1dxnEOJkOPV+wDarH18jBFW4y
PiuuWOxXV05kKzjiXK2mlK6sgtA9zUhKxQZqxSeie7AQwllwkvuiOvPOIhjw+WguxkGeNtVxRaPO
+uYGjA88tMut9YLI05Xgf5lJpZwLhndVf4J1dwDazGI04608CdBhqYRGXz6alVsMU5/kxhf8CaZs
7Bg7bFGusZwCQPVomMuuKQWP6ASkjG71ExAFptm6xZZfJTf0OUO4F+mZUPLIDhVxrCkyB8losIvW
RzowyUi6qdFK0YH1Gv6EAvz8qT79NweJ/5uhstk/TPmArUQ4mOUi8PPgReo9QvQDaJG093ylqUot
rOQE0JBS3YhBOs5yPVJwNW6FN9y8+SO4QKaapyZlHhXkHXr5VI6epnoeOqM+a2sKOs3Tt59P2Goq
DU0wNhpubsjLYFkFB3onZSag+r/v1NTjI0Ys85St0bWcbeH3jnmG27mtNrBMD76CpD/n8TREHF5V
bZMX3lRevzsUSx9jCM8fRazBApH05/j5RwsWtbed6eRpucr3eWByAjvQGVE5a+ySihBurBqpDlGv
pEDxQ1E3LzFu1D3YsSvRietWc/igsehauKy8hIRtcI9gDp+Qs32FNupyCYhKJ1deb2SdwbpmAzCO
mrOa6Bj/99y3p0OvEMWfljP6iB0gSNUONYzz1sbd7HJrW45vTF/gz4lDoEcP4+rtHLs7oO5b5ode
S77BBWuLUv9pTwMNCNZ6OdGjd7Nb39meDA9QP9eFNZcXUezuQT4nh+/UBU9nIL+o6xJg2cjIclrQ
551UbgfSzjzUFs2dgESdpbz4HSE0gI7cCeWjRQG45+R/FnlKETzcjNRAdljMh4kGrK+DZIUY9vO3
o9n5ueYstMqkH5gyEr3iwwp4ZxkdrU8D5ZUL7qp/m8R1P+iv0zcVuRjGCcw4nCLtE1eC06wU8iUi
TYJqrjmnpGqibjONX3NDcJl5DdZx1xt/OdGymmMAdXtFgO/+WN36oUXbtlWcaeZVv+4Gzgiwd7kW
Kqhynsn8UQ883pcODE0bDevgb/1KsUzvPHQp8l/VvxInVGqIFHAHNJTZdVNb42FtIx3vrblApr2O
urCO6R13AvO6oC+3q+b6z3zEQEu3wLPkS5jJLYGhV49973Gn2DLmjTpJSJ/7Cm1Gn28WjNLqg2ms
69JiuTaGF2eeUdLZxuQVD9UWFNav2cEgl4BXHJfRLSTq/HXKPvSfTFKRqgELrtPo35KTLoMv9kqr
nxJnhz5iu1BxWbnpRpgR24QksQ32GpDjiQi2tC5KhwTnIkNXPiwS8hhkrZPQETDFoRDxOTlaQ5yp
pdrPG4HkCXgjF/dNZ5kxTfMYZvDGEnapCcfw0T0LU08jClV61Zt+rbYETS7iepl/OnZs8GBrju7j
Sw8u7tsmU9sfSK1mPHJnOnayLCI0SB38HWPNX0VKQdWfS+AzjGqAbMv+rm0M7QNycK9RVqnXKfK3
MKcW6pynruDG8gw2AUB/wG/dkwNnGq0R48an5bZLI+RN+ERO978nEZq62s2rcIqfgWtBYy+a3f5m
8o8vHsGXcQix6GBOqc2xN2TSA2UTl06MFvMqjuqkTNsXpf+fuqVWeBW0g3Dr3XkCzs8XGR2yXGPm
b91qjx6IjuHbjazAxREj08gUUCeDtMaZj2sAqnTdmF0v16Dd+89J2iM1Cgh95kLqmdG2muKWEjV8
+vlq+8cx48Xm7oRgOqIkdFSRZF2HuhcOMl2hH3u6YvW6MP4Ux4afYCY6YMGVQSrl+x8C+rGrEErE
8y7Jx3UPVhluq1wyWSGmQXdI8d4Xt5ybXnICAb7+bkg6JZF449UvyOiSPTRF0aaVaWn+swPEehgC
+XOUfRajS++xm/b1NUoB/VkWcut95utOMOYBM2nUku8G2mGe/ra+QdBq/dVPalFTHwUyxnxSaJq1
JTX1Tt0IaFpuqfwjgD2XX0B/NbmAleD/SlmbrwGRsi9Dk09h6ypLm9ITnAOwB0bgOQFMjxi0cy5Y
69SOlaAxansGSXFUaQp/3J3dQwEP0h239WBtkuRB2+diUJCNTitKpu7QDPaH0BJV7cPmJaAxzcVT
m3rrTpYDte5DoZYE6F5smjGIMP4jB9VsgcJ1DCvCOJT4hFafFA2g3UIebSmTRuq7djfRXLPdD8Wj
fQbi6sPAC/pPWy1pJ2oTIWybjaF7PUlBrfJUUpL5WBfR7JPQnoaCdD5g7jTN7tafGIg05eM3Exz0
YC4CCdEyUWp3GjdAXIDYMvjTdqVhXl+AK5TcldjMWAUZ0D0gbCyq+P6VhdLeHPqSEc8sAd5wp1cB
HsORHqyRh59a5FqCWfE8xbZcIGyXo5VN4L1+qUEdktBiF6ktWIeB2FxFU6Ehw/aefnCj6R3KC2cj
AFJLl3rqMqd3I7LjdtSj5nHH4CQk+vqqGE9cF2UeF27cS/LoUho1LES7hBP8t48zY3FoSsK1ObQa
z5z8UO76dGVWgoQu/J5lrvjakZri0pI/oxBWLfAzbcaldJBg+Mxu6VGeClEzQs2LgjiDhG0vbOHh
e+aq3Y1MYq34Bwp/jVujtchU9ZQ5wdMgs2yD1/0w2LA+F3DGulES3NtgrwOwgwBgiLRHK39zw5ZE
Di4OrS3ntj6098UoWPATIdzuFZC4SgKZ1Z9tEBIIpV/7rhX9D2uy7qnTKZCpePlplU9r9krO+NRl
cN/txj4hWYUauqUB7SXUl8DO2C/bUruUBpIpu+S5yx1MNaTK2TnqXjxJYY92nnnvKxIZREJoGN+8
b0a9Rd6eYydv38YhJRO4OBShFLGn4nlvBfYR1uIDtRKDrWZ5pjIFJ3+UPly2to0tpUV3kVZc4nhp
a6NtlvCASOXJxApqJxmM3uLeAf/0ifpfHIm2kQj250aNJn+0ZmbFUF5Ll9NPWpSNmpww+/roHc41
ft/MZ7rwSOs5ZoFPnx2ZvkW1B7IcYOvdPoLn4xNkS2Jo9X4QnuATkXwN1Jrrb9S9+ZyiT3HTF8Po
WRW04UYZbHdi7KOwImrBHh8Z9HmwRUvuh1QrHpJ+6jteUU9eKvO5ecm2p/jNtG/d0ktkqy7TN/fv
t2e/DodzMAquLKeYVqdCipNVtM17uBZ2BaoXMyIlLtMXyrxgU7BzSe1YfFu4Fjf2ylZf7XNwYeEX
UW6fJhvJm0xmoBI3Gir7a4jAOvS63itF+qVqiUldcE50let5tOYm+Qmukcduifsfixrv3h+KYHon
m0k1tkCytHyinznyfF84NubCbh7qXdAgmtjcpuvyBGOA4sDXMnwGFZ4kFUlbQUhMQxzr0lpxMgAK
gSG6FS1yklS/FuDI92ru7GMJFA0SIs9V6bw7CXR+m24CyMyRODHge/XlBXMYzTluZKkBWYX8yQx/
xtYYwGVbLeNm1T4Kmp2kXgGIHC65A1qKCbWn+qbJtLtgUIbkhladoRACr1/65ksdeEuY9toBOrdS
HN4s79haJUFGghxqXFYTzEWdqlQR7odo5gKGTEgFfLRsg9Je3a2v6vUwIZPSzhQ81jfcAENs8v4L
PmpECPc4RVTje4bBHAzZNVB3NVnHQr4BVbXITILZ+iDD8yXrNFYhkKs5b+nTrr3SbLZpWIowJPOo
tdN+R/kxwn/yJR7IMy3/TZxURUpx8TEFUmRbhOpaxnqbEE+/cvvd/OgavhSzytpN3pCDWvZqvbSf
RfMB0nCYoZKO+QH/JMy659extYep8yM4xBogATq6GWGKTLs/u7mnSahN0SfU7xQr/d9Nrz/tZi1H
Mg/aaOw3YqZ73yz30cFHj2fchc87OQV+txkIR/HuxAhcyXDr6S4i6iFT6H6e8DX8X8K4Qbj7US8g
y0VxL5SACNqHvhCkROuIXObUPAQCXlu3rt+KjQ+ApfSzXO9HLS6ks6NPrmbE0sGs6A4CnBkXyMZZ
MBdSpaXe839hwrmvb390d3hfMpmb78j7sf+qxp+X3r65wVBVYzLxlb/AMbVrlmnV5WgCzPbFrX0X
EvfcnF18IRtb8INKNoPAmUaJYIv2dsHFCKqqNA43dr7n/EKMgQIqxlm1hi1uJhrXo5lr8V8PzK1L
s5Octt+xbLQFwM1nVrLK0VXjl+yi/mAC4KCoNSwfbRgYeQylFHX5hEhTqj+ilcb/27zGHsWfOcTk
ryNKA1Kx7osGFtVwUcO0JEyRgMWjbIJKDknz4C2DCLuDILVoqt2E3i1Po8f3BMsqE3u1ldlw6im2
nl1CdU9nv+eUNU6gPGIYYWCzgReEmSYCCZY1IV7nsNBpW0BmKLWKKr2CPmRNJ5s5Q4LJnCKjOM/o
pnmhLLkFgKJAdVPzgCCXPOhK0vPpaV2nuTfCj31rdowGW+flE9NeBWpzZLB77Oe9dhnumIFyNYWX
U4sSdl9cd1VgCLVKtkQvy6xYp+ujzxTzN3Pz8O9a6nK3qDZdz2hBimcCf4KcWuFGcf2rfUFrd6/h
Lyfd0yR+yawweGQECTmITh1GlLU0BQHlHXdp9hjgEqGGXL/j3xqziB9RDmTBM+CmF2PDCA+GhSZp
WAisOhejgY0wT2waq6e4zhzR1I4tsq+0fGNn3vmcIcjV+2bQ6XfwUXwjuA9tOjdiHkFS+oZZnWfH
/3SKLpd7T2sjI8wM/fJmyxvVHfvBPRuE/TP4me7+kMCXCVcTypW6rxb1N+1pjX5Ogprf3CZh/vCl
RbFyOy/3la/4Q9fF8RTq97AHiE+puso1pSh3cYJhlGPtMEvr4Vj2JbM+0Zp2uMVeEVIw+wlmTp7f
bmgWJw+DrtSaCPnHz0EwEESr4vu9SU0vMNPtOWblZVuJy6gyFIZP5MaVU+i2o9KMpb0d4BXqhQ+k
mQJAZTbvN6N6ECj/SJe09KgTBik0beUO2yFUS1luJg7WjRF3ejmoc+zR0WD1vtxyrmCpRIrCLNOd
Zyu2pZsDm/wSI8dpceXqN4uYpprpQIaMTkCoKb9NmbBW6Edl/YHj3/T24cbNhT0fCHoyinJFMHG2
rfWXfR8ttQWuH3GIGgxvo+Yle3XpGSCJh4TylstO6xQ4cEFZPqjWMfap2KH8IYVLpmp83b1430Aw
AxD906GGmLdpLyD11IKYkov2NRuKBfLis1RB5fka3lOc0xXhYOm4eFsyZEhKqpYJogFYdkw3Iu38
XKGms4Cgnz7S8rPZYDz9jJ/blgI3nJQvvb2D4FD0p7ApV2RGDnUpmgrekUxY2dV8md2humkcirfK
/StzFQq+uEroNwvzBKC5xzkKVCamiKDy4zihBbA46D6fGEryPaw+2Bz6GBty0s+61wJVe1vVzZF6
QHPxHToqbAmylinoqNinGAsN1WHquhOVc0El+jKIpFbr38wrmH57nYzvxwyk+BhqI5XZT4R50nO3
CkNiL3uWjkFcSor+7N7wJo6fEQjoAB6MWFqGpWw46nsnXiGdXw7VLqZZzZlKrqyG2E2u8ZPQbwss
Io7r1DJg39UERe3trNtdWugNQ/7LzpzBz4kNMYHwTFVP6HxnQt9Xsf6TQAGIxuryB2NGgeTyPJcU
+5HElSXH3pzLegsb61SoN+cldOi7daPjc2URBYQA93uQhosZhxaFLoIYCShE+yb5oK1GawW+Nm6E
9ws7i3aqZU/T1Aa50QD9JmCRscnnm+kzlC0X3ieLstrd3Fp8IeT/BWMVwp6ZqG4mFzLUp9HKYHEK
LOhm6FC/6HQqG9Fw27y3A0BszA3in8NzTRWfmctVQd4VIO6UJcUghQPkl9dvgn0hEFX4WQnQ+xLL
dZXjHh+pmZwitWU0bf9zXyha4rD7U2LErIMOs9DvnCJ99Yif2kDGtPlRjBFLGzBMrfkopvKbYN/s
o8MQLIZJpCszbjVZ5Zrmgz7e/K66/RjPZrvDnDFCp2EK3LIgR4eCJ8fy8ynp7QZ+QJwpThtYLca+
/iMz6+MGhLT5ETYUotmHWXINovjFPMdmjKKdbJ0do0C7BRn9WRKmxcyfFgekQaRo7TNIl8WxWM1u
83W912X5YYL096SqLD387iNEvWMFFP8e9eiRu8f2f1H0tgCVrmA4SO8Br08+e9/pE55jgklJJkGi
VZdpGw3RedbqwASJfkfuBgU3QYM70ACAlwhSZTVdCpS0+sB1R2l/XX8V06E2NTwRvoRI4SLsvYKP
6EvZW+3S6uWftvySm4ZNStFvpWV3RtkWFPJM/tIqfINQhadk/CqyETpE+4Gmb4UpB5rPA16PEVkD
8euUdK6ynvYdXeteJ8cYqf6LMjqbGphIfga46tzpTb6X198uHRKtVAEX1antqp0z0zg51Ot2HVXi
jNQ7hGOti/YQsn7iiGwhys5un6jvJsGYRh+qTAtH3xEcIwpH9FoIf1BKlPdNop6eYwS5Ffo8fkBO
o0pdT6CveWhfcTEzQu6BhmtUi8QJqyfWAvzT+NCT4cRa9c3Yvrb8s27NHLJxoBEUOGOpHRyuFwSk
MZouG1rBUQ260qjb6IfEvVRQfT+gQxAHbeIiIFtmoHfOC+SBbv6iSist43HOASE8xaTzf6fzWT5n
JjhIqJrA1EpviM5XSDZJH1alGU263v0Hdmn2o1v8wy1xQDHGMEPUEP9r1I5KybVouEeNwkNlEOKU
oIdY9UwSOGaa+nKCbQ3tqvuV8X4nm33kWmRY0BATqrhQL7scbTA8c+/d1tmG5pLyKbZQVJxfVSkc
RKyEoEeX07/NjUPVvb14oux48XQWnq+Zk9ZGObZB2XCwjN9zYsE6HFrDt3Qwkf7BxOhxvZjNfKUY
KN4+ZE81Tx/nE+CMxx0GNs1zKqWuRQZ0OP/NOQyt/d+AIuxwlTISP4D4p1bMjxxcyl/tY5cjNa2W
YOI3fhFYCBcFJWam+DAdOnJ+d2zIJAn26CPfbZeYTlFtYsZThbo2gYBB9mSxhfhGiY+0EtE6zJ8T
RBAu4d3C+i6yas02r5FhvxB269+IumdC0T4KmsL7r1bXnuUuDZCCOy6qqmhl+iP4fWL5/0SbT4/t
YR5/P2/8OLacz0SYeO+zNeEJAs4XI/Dc0EQnFzaYXFnh+lMWWlnAlTs40Qyju8kVTQSEAXQvOV5n
yrcM8G4BYzPmHf8GpWxnE1morWyeVUphZ6E5/4JfVwTboY/NSAwIXB6k1Ty98i3AOS4906OoP+Cw
OOABJPdmAVfLmarVNkHRCteoR2Y8nujU0ZLLdPBi+QZ/ArvmQMo0D11ZWbo75wle0OAB9H0NjF/E
U7NmsHmMdPaTOuz4Yf3VbRhYmgM3bDg66SPk7rCQt7o+o2Hldwv84ivoG4Q5F+wRtbk3eyhAnoEA
6esB1P4bOUVVtBnKkIxm+7JNJ+EHxB+fv4KGsw50HEFqjKdNlCwGsbgsonzs1x8N3mdoSmiR3IQU
t1OoNIwLBV8GbKIZSJMWf59aeyFJLiH+oO0bep6Ovj47119ombXRIDPewFwrpj9EKVCKiTT1fVQp
vsaVqmI97kxDpAvrdWANz01uIVKpcsWLtlp8eoPswVz2aHtUtybF9+tTD4sUyTK4uUWQabCBjeiO
mz48PHKeiuJPcGc5sNIYcBJshIFxsc6clC2XDk/w17ASMQ9D3hHLdMBm7iyYB7IVa95lSlaJqBlu
vr++55QpATPqyLHwflNcAz3Gixv5gmi2G1gqm+/+DGycsISeFEI9opldPCDgw0smZZZx4tvVVsjr
7oI1h+6Z06mc+k9GBVtXc7wrq6em23Kf4BEizIuHGeKZaM1SUkVVpKoSphwMSPKghXm3KtLJJ3TW
Mefwfv5bqmQF/AGcO4iMIq8J/y6T0zDsjA57rPcjZ4WLdUvp6x9W5IZhqtpYCyPwOEVHGIyDTHPR
2PRjwFPdAU4Vh7FLQG7HEk50pRzbYR/j2TOwI2pQGTp4lp2Z2SQh4jrC4xPK1nnQ47WR/D1YW4qz
4XRRmbuqJA4dNIhwLeINss8C/U8w1IW1dbemb2hd3uvzr6cGlYkMF95LJMDkF8Oc1Nj0RYzA2xtC
GJD8qU8o8QcgWsSwEwdDzjpPdoX3pg3V4qgYrLS7LObjvJyCQeNW5CBjX03iS5yJkOpgKBC3ioqE
kSPB56tQz7NagtKVCnDxe5Z4bhAKZOcy0QIyAHTJ3lp7u876h5hBA6OttVn/50OG8qnmEW40vzW2
gOKSkHf0BEqO+4FJvGZQItv8agNjLw42rE7RkcTMxvp66XRYz9aPq5j/SeYy0+hnzLxaKsJMl/do
VlwClFGksxYtm8gSGnl1YJTxOx4IY6AD2V1n2N2qgExZWPQeHqBySPHrMjuGF2FzoGBMifHCLLF4
XGMCksIF0FBh7klwFfOiM7z6KPQKM/p44P6YD8CM1AI55DEJZvm64vObqkiGjdBI2KrkJB8JdvgJ
3y89B28CYX4Wv7FZqRFOfMx5vyymmXqbAH9VZoIXdDy/kWVG0fTOD4hqfMxUKQ7AiHgEryulllUY
+Vj43KS7yNi2ajxwDR4pJtDL4fuqggR6RuZiu1BBoX+a7DE/zxjX8ipy6WqWvDmO9wvZKgVA5AwH
RpEMPhrKavWO+dYZL1iX43r/Qy4l2jSS8PL3OAmB2YhmgTX5nQjqNl5cozbmGdTFKQdw61dJ+tuG
4ge9ymeFREyFqIkNecfymLb0+mwuEmkAi3wm0zUjAwVR37BfMdF7OV8ggxuFVC2A6mW45HfL7HG8
RFUzMnCb75oXgJSdNRp5O0Dr4snyUk8OomDJSdxktRrDFznDFNx36bUvjIN4ScUeT88CSDEPJFRd
5PE/60IWagxK+4bvEGxvsnRPwoR/sS1DimiJTbe69kEP4MM+MP62sPQwJ3HV78RiotsXaywer2L9
uTtsXi98xWNRUhZPdEYWNNv49SiJOJxzK6M6wIAlva0uyjinsoH7U/xIBr9coMPbNQk4mWwkD4Gy
zbypKDwfifZTRO5SzhVHW/uq6BEPHOrmhgSOKEQSH+hOk+sfwzvC+QOCehSEZotkFyaCD+90SKNk
eKxnwN1UYDFIduBg32JKbXJ+HJi5g0ChJEWpaCafpDUFhFvPA82zm+0ZBzhsuOh0ckfJAKSSVZfs
KDc+OoSEMCAUV1lmCZZbSQmCo2wbQvLTVUwpuzXgWNDmCnTEYat9WHiisuxolfHEvzYNngk18uBL
QOK0QDwj/C0ItkazrxvAr5nzFQR23cc0iCQpNk5mwrJOj8sH6a+nqtmUymfeEl1RkZ6Fz36ROObu
19BpZtKJR2pywiUm+dohjpIB60hlNuJYAfHDHJfCw0IC8QoPW7sa1TcUQ7kspQPsGlvk/AivxLWu
xoUZZU/33amD5CskpjaH7PaaGrG2RAf9NpMot0mg/WrlYQMMfWQJav4SeMz6ylvByY/OamxDnAMu
PhjV6HK04Fc4g835lEoH8ZNlsSVuzkVBbbv4EoNIUdiLNwqjr5iNpqkjJeqx+dABJA6XCTTFkTc2
EgCxF8Ft4gtAx7oFV1fJQse8mnSMFY6kDpK0bdCNuv75PLJndv64x+ixExk5q61N0aovUaHZNrcn
ijD7+QHt87qiBqfRofFhOK19g8G8b6BPJaHT0WH+IkDN+x5Q5BlkeLQ+61UzbKqVNWk3avbh0nRh
ns0kV+LeSVN0BGcF5GH/QpkG7Fc4mM9iLblhEIWijtSfzR5doXNxNKDYw7Yh/qZHrMOInOSsG334
WIzQjUCxXmL2xz7ohdYKQT6I10ECqbuArk2e8g0tpuvIgbpe8QuRyDcWIYj+zfYbuiCZBkpx843c
WvemKXUeQ473VVtRe/Hx9nE6d0+BvIRe1l/2hLySfTWg+GbRZeIqq2b+26qwnPc91QWeu+ZftSlK
huGMKWNbeiZwXnFAwu6IasNZGn5xClo4zNC2dgER2L04SwiDGlJvtfUt3pio7wcfHIboHrHS2q5A
9X0hxWlyqiRqfiGv3UKOaD0MO+f1omUK7NP03S82DtSgmPiHKsYBaWEegrknHEDZVpsJW+Ak7aNO
04uElliaAcy8QlRc6JbVDVyYDEjHBS9Besr8V3TiTf+c7akDI8g/wNMeIFUHMsfpxqD62ZNELPKV
xwP6zApwLjJzv2P5Xi5d7X/EZQtfxXTGwvX4KADTaPFHW2JMqCMxnFhS80PeXWgO9Ha6b/Sfjhzd
h8OeMmAHza9CKoUOrNn7HaYFPnzTrmxqGOLDL9lz1eXtlpp0JwT5B9jClSu+XXZuyq5/7XaaI44I
jR1E3Er7lhevjwTMGkX0GhsDOzfZkZzfkUaLicnh89/PSxW+hfgZ4eDIYHZcupgP93lxg2jld2xu
eKqdCr1v98EMQB2k1IKB9PBEaU3YhafwU7nW9tHmu9ntiXIYTgWKsJ5A8AKFgfy6XX6lE5VmrFU5
9kiSx3I5B0qNS9ctPdJ753y+2PEvPtjZpZq+Dhu+TAs2Yx1ZeNhLwHWk57TAAKRT4DrbeZMEhNgB
tcbPO5WrnEyDRPok0a0ehQMp6M1y4kNtfFnds/CMqErTD/qg90X6bxXU/KIqQTfzIcgBz2SJGcUS
53ilAtusLyPPQ8mJmn7ax0hhWTFWdChUt3RqrYncUNeORyfpSuFrm8oQFdy5uL1yIYbU+8qEQX+O
hxbI2hQiwRjtGH8KYU7gOtUAHa901mdIBw6L5J15FGMLLoPlspaSvg+KG1v7OlasXKTuLsB2s5uS
R4H8ZRjO/9Onw2eQRSs9CfgryZmYNWgAB//EezYVjAv8/iIkIUfWP87TZmPpYtL9W0G719yzn6Ji
MkmXPIyqZ+jFgKs1pyxodpn1MkAc633qRRVgkiFddg8kHrFuCA5yl+HpJM1gTt3PhpIwqH+zBDkG
5ufuTV+7ITcgSgd1LO/0ClBrZ75GGr2MFomJGi/WtQ8loKqNNMn5XYg8D3KrPvyiKsDCg7U/gvJZ
YxMw+gWpna9BSKhIKqrPYh0bwYqr9gO0etHIF9lCR6OxMz3lkm8WXCypIWZn4yAtB9WrqhrLneeQ
aDCfuz/x0OZOZk77J9/Iut+XNBF3xrYL04jLe9VK8BbfqSblJkaJbDUDj4VsO9aXDnn/fAaUL0yZ
1AD3FFNWFpJCfCPI8YpWOLcE4/Vq9l9stkLp3hqBtGWBzBNeyfR8Tt2FlI/xRdF5JU8wV3k3FL8I
QNEXFYM+S+q4s6GIly61+mg8/NZxTDUfu2+3e70PHPLJtA9I4xGO74wms9zyOAwApTa4NhbviKpQ
2gZIM5Ny4xSSSB+WGL5hp2wZPHvNcW9kt4cdXf0nUb2iM6gWmHtEjEodFvoC/gnjVaH9scvq+Rid
MUv6xjZg2lHaT0Ll4E3NAAZzh4c0CX4GhWNsMdLmXsEoAZHJSlkRfq6/TsBLytc8l5eKeLQ9SVwG
/Vd0Wtc0ghFnayX2vlkzj+VdLjcroPCe42WQd6gluVdNFT1t/IgMwIAIkKRUOUH7qK8TzHksTila
83ezsk/zsZS1Ha2aJ9EuIEK7xhr2yGvt/DJLdSVgT967zHQUlFyqpYovvkAQ/V1PDzKiWqDURHyG
zpE8E8Wf9D6raG/FEKZAHQap3cji3S8X/Y7YiHI1iwv21rSUR4pE434r3AtP4kS+YIR7qKR8pf3w
K8RLS/P67FlIK715rHUWNUCdMc5PykSHTJsekC9NKkJJBzU+55DCQKhlZYK1su1t5t2YxFMD7ABc
yWxcY5JS5BgmRHOAlU72p3fNnZuBYvsHAblUfL8AnoNRUhWGQwdMVdXlSiVsjINo0eZ75BmDDzzl
5rFZZ2S1l1YOKB2wDZa9fMH996D2l1TosJ1uge4ppf/aTZ9rMnga4gnZuXuMgr6FlgK/WvpJgfYf
9QJlga6N1XlURTYP7y7ifvOqptDknhMzuVWNx7BTBipyVvisgSMWk+2cx8IdeTSrpGeLiO89OpdC
zPVu6Wl484U9mL5oJK7G0v8pGHN+YvrlQLRsKGeRG8sTRRUQm6OcGaf5BTt+lyDKqvR6OexfMald
1D8dELIprJDSB29EyWpuvpaEPcBELpkl8UzpMbViv8P25MS8XN4XceZKYpZpm/gh3lheC3+izE6F
aZLgcbyPJjxSJO/GTyUAux/Gmtcc52V983LmqAIvgJItd5zqRER/eszQ0a5zvz32IMXcclHv14NO
JrA+zhxr6WZ1H+qm+e7lbLP26BFv5gBh45B4slxjRF/yJqPK8ifGf9ifWcr3pfV5wsTIOCoV2p+U
5xK5mSwOwWrefZOmmm7VbXXwhpDyK/PIpt4eM+bYBxV38VJmcEQ4bskDkMwX2woHQ2y0Sm4NHj/B
mOyR/kFn3jvdzs8VKlbk0OrXYn5ri2h3hJvaTyzOS3kN7nk050lg7/eO8Uu3j/wx2wEl5vG2eItV
IVxelx86J9MRtqQQGjK7S5m5s5vXIyoPQfM809JWT+E3Pr6Oobh6DOKjADci7NZXSAKtRJ1rx3fM
Ei/+LSdL94gtODRWC2zkMT9kzzTPOQlqDvIS9Wr1e9QRtZV/FH5abfVXRK5IT0SA/nsYNozzjBBQ
Dd5g42uIemooS7cNajxHOZaRc31+A8AqYQuuUsgqwZK6kdCe4DNWRDAoJ/h+vintfq8/wALUT9Nr
8skQxwcNjOXFJJ886XjtwxniSwh72Oiam4SJZfk9ujXp9Mph9uhucLIudGnSrmRsRvARlxYHhHPq
peJvGaSmyOfnZYmatwEYjrbSA3hmRl4PG5u/uWT58owtgXte/h7UH2Y0mNGdgynGc3R9y6KH6/sf
r3BrKVgomaO88WfIxZLHyIT7uZgqhWiXI5tMyGuqdVK5905YRIkpwsrysEDCdH8RbEHH1gHBSNbg
BAaEI7Xzq9UtSAdxntlNWDV0lhjd0CCW8gZTkciWkwxWxB6zCk2UKWqE8thJ1xVYznfgAVDQkPsT
fOoJK1NSV/nVk3rjTwp83FNXFLwHf73oPDEYIq4knUNZCzFtVdQvl7kw7KstOtL8jhRxuB9hfnIl
mpY8frKgIWiKZgJyNvyKKBPgdquDNTk1ThQ/iEk0tjC9x+zm+WqioGs+zNojJeaR44j2Lv2+rMPl
JRzOFhYiO39hFpnRUxTHqXaLIuUs1L7JcpJXSjhjdOhe2FmEo5P2ZRQ0ecW6yZ2phdXyIHpdWfEi
NxWCjrSF1UL9qW0BeegiaT2YZWhC20pH8ba7GUKa6Z5xOSzrspKm4ag+gAYvcaQfZnfbOyghPkeR
Ln3GLpVpNrTfyiCYSIIPCoWergb+QzY4hYPUVNwiZtYrweCPKjjDjHgwddThfD8karde9uf9m5vJ
lnPSyxXzv2Gd0WnBxuCDrduV2WGOZNiiZ7AjvQBZhSmSDmHNoWi4w8SafLQkyIQGZvBih4R0YrEC
FxewKf4fKSSgCX2vii+kHH4+KdCx6mDMx5g52cLW7dK/mwhsO+F+SlrXVzwERF8zBy6Bv4xtOhBw
qkIiQRtWznDPYzEK/s94t4NYd6E2jBFR/wSi3KZGGF/nUCr95QDRlcOm95ZzaSAsqd+Trk9RSpj5
ePCyd4BCknlTmfn9pEqh4dU730sIDwL6yuvCPZ06gMejJAI/2WFjMwqeE3iHL8s9s/Bn2tMKLYGh
Frac244RLkM2FwS3vi8kW3BeIToVIXLBRM4NAP2OeSTcT/pjR4bYMNfHuMtSpYDeK2B/TULicDK/
pp9M/pihk9H5fFsUZ8jZ8nAB/9ay0nNKjKv7/TMwCCGPLwkXH3v+7LPkp3WFPDPFcp6nuB0Zudp1
1jZmZ0lBpW3R8yoC0UkWSITrgDrHQiP1F5US+HqgCAYY1MNk2YtN0AWFDlmAQCE/zQz2vnuFX0kY
IVt+h44VuV+jiVY+IAsclppR4hV1NSLy9C2jnk8kJm29DK5iznEve4w+4TuzKJU3ErIyI+44uRqb
3fw3iZhZTvpytotnjdqfKIxipIBous9cSRswqG/clkOISiRyNDKJ0gGYq8QVKHNAuE/CnpyaF0KK
xUOSFm7BzXUV+VKGu7NZM34s+mtTu7SWqUVvEfbkUUvaevT649GujN32uiy4bohDlN48DaZsQlBL
6i940Y0wFxT0ek5L1QLoAot0203DuLYL9aVuVVvSgpVrI66Rn7EwcuVrmbZvEvzUAz+avn3a3RJu
UfrRcfR+ns1KxgbUtiERY5HTLw9odsn7ISAZjKBparL13cWrN21wg2wGglVuTquq9Go1qjYyvthb
ZwK6DO1QDCbv2k/ACpSj/h1uASVlfCdMDS9jgcNBmybc0CJhYtdK5MNYEanvnp6qUdT1Xzn1tNDV
5xVrXVLD/CK/IssGGeVvRaFznEUZIsOWtj4Rby2JVi5JXqUtQ/AU4iAqpOhsdjLoeszyv/FqKp09
qAubuAaebt23drM5KewElcnyMSYIU0ZZsWk6vmaSbgcnQe9fCWvucSuzW2bMquJ9uylFCmBjHQkl
rHHYXjP7QPBbRHz395GVkIlvgFBxGxZ0y3EPTwG4mlIfR9pSGNFOSwP+lDWXEHpKL74XSBSfySZ4
GrTXujBmLXdd9U/GcFKZMCBCRdFstNY2lD4rOWQ6gwGffJNVp6wiL9hvDLWpxC8+BRYWfZJENrW/
KhZIOzOLr6453cdMSe7bGLAxrxZzJbyvUK5PJe34teZEHQMW8o1jELNUU1LeRHe5n6sadR8o8aRp
qUDxfitfTlC6tn7H5qHZoBZ1vDM+0kBYYUG+qmdIZxq4ykOqZCgipQEDegcYQOX7I+vPT/eINnXr
mngiVuJCF5GIhiueJrNzrsP3m0hxV+TN5nNdg2IA8BvCcgAFuM47l+mU5VWrphLM/GEJY/ONfNmx
/1t1Sjg52doN0dKo+pY2cwgV/X8pqMdCmGl7pqWwk00ZpAiPc0OBLTqkaw8ay4fCuT249mmkPe8v
L8hryGnbLVQj6cRPAqqAeT6N6hfiIcfzKInwO92l8fuXYBdLcbtVy+q8kraY2T6JbqBxyWjlw+Bk
w8jplFkRI4bSIUOw/9pWgOc/HDnh/XryUDffEXoggp9qyyRtZXIu1JzNxqdQtmGJpMgvFv7g6dLI
Yta/ZyyyriMT5kIFbHgPJRJlubJPR1ih/UguhYnKLubSg/pqs+2IZnWucHgrzpBt6+Gp0HTBB5Av
V5c7V6ydoxbCcn4RuDa20c5dLxy98EIQLLQZXqiyqM8vJHZtHm/tgC/ud/cUXFiDm2GFzMMHqfPy
6snmemHM+6V7v1aHLIXcBGPWgJIcN8Ppivt3sKo4Xyq6VpJPCLEEpBtwp1tXu9fBMwEq+l/+HYKr
cAHqKDFo6EZV7sLM/UuVdcKoZoIJduKu6jQgv+Kko2d4mpafKI+bEp3nwF/IR2nTbLd36H9nboh1
94Kb4Q3sS6KoARLFpm2eMCOrt+2TGd9T5Oj3VR5Hulpv1IGzTstGalCLs9PBlagacU1wvQyfinOq
pWRG5ZMhsqdGdAvYxzw4wI+jzr15Prej/Euu7KaZmdDuIneCmx3gU50OoaOD9oZv9pbucalhPnWz
hBDsfR2MM5ODTLy8ptOkLCOXeOxRMZuN3AEcv01G6aouGvutDxd+NHAleSRassoajwAoD4GuBv2/
lwfTXmEbM4NA5EVjisPV/nNPHwBoJtjAkjkjfrGrY10gmXYY5j5PU94r2lWowILibRxSnhL7u73k
uKY1/8PgaladKTmF8j0r4d1vhSuDOSQrHBykhpF8IYYABbxfLO85UH/9OaXV6HCHv7a6co9w+sRH
h2ukFWNBITARlx9dMoKHbyZeAY6KASfPUZ6HlAmCVr3jGZsy3O1koIYkTWb+LV2DtSTobpc0Lvc+
0tOU7mxiFEGx6ziADJSe15g7p3EkN9HAWI9o/QjNHXWNY1cTXsYA3nqP49ot3aDd/QnVQWRk60ir
dYViB1Ts+Y+hXiNjlXPqem6i/zJjP0buWxq/+8Z+gU/B8EuGt9wRrS8Q8VPEvz4NgONpCZZ315qc
Qq/FPNJY+WR+4glcTMmIho+0Q3gUHlq4ZVGRfc0NY9XuM8DQXWwE1aPXK8f289G4+0sfk9yfMete
pXNR2iofG/iAHjMawt2jr7/PrqacRPu6jtvdF67mYvKo/oTbypq//BqUDylRHv0gSEaeP1/Sred8
f4VM/fJdrIj/B/1G51Bf3NT6jrGEoOjPrt8tsS/g+C6E5s3gyyf0ysJBMMCoCvps+btaXCzYK5CE
MrfoQFGhvixtR9itOpKRW+ZUSf8ZatMHLHdQyHBzNCL2SKd1f3VpmUcom59ElnJ9jC4R8zZeZHUs
VEl8Vqz+pHJ734k2aBT9yURS0RSWEeAHXLSMlkl8lAKKJOSmRIVzbAEoFEezev0+bfXDOajFLfdy
MvSDHu5zqXeoUn+g7RyJ8V82CetselVZE5w8uhgcfAM3YRArVuW63pH+Nb8/3Vy1ucccKl6t2ONn
ddIiiGimAV04JEWJrjzRTcsh9SpXfKKZIT5YpBmGAk6PWYmvvz4PsEVlcG905lxHbp9ZRG/ZhfMv
adFkHc0hslg66EuG9tBGkKKafVvjh0JDN2TSU/hzJEEYC/Zth9nK8eMs4LMWENlw/vyZ78LN1NW5
Ml5JY7fBzSGaxlmdVyD6PQCLWHKZ48W/R2PYyj6fWXXAnfprqKkECBKni5K8LSmJjgNU7MCW4Uhp
nNJGjXYpqZomINNtoQxTCsYfw5eDSPGYcyGrbnX7B9ZKSNiim+Hpa0Bp+XR6nra8I5fRqjzbfDHc
sWVXs5vyS94rrUQa4z13fiD1srAMPgNeJ7So2UI3Ppzc3m79CLiS+RSQk09qk0q8ab62WzuJG7Uq
0j/mJ2rOrou/NSBkJDDP3qIgGzYklezZ1ucpi6CG321leRyhx6AT/sOi947fn741Yg8KEHeHCzAD
5xyA4eJd4gq2FaedV1h4r4nRCwmhWrmUtTfXOY8xOSnf2rcrYJd1+I//llMTHyHiUlGeIQd4UfB6
oTcXYlKanRC1V7BFugVCMTpHTtoRueerF6Eq+Jd15IU7y2MULr4qRHWcuuIR1LoueYOCsNa7u2q2
e8thBHY4rMYNg2U8l5zGJqXgV/mFmKocOSqwU2Jfj7i0IjTy+H7VnKR32sC6jQEyYjwrEt6x1bRe
Viyu6crg32tDEd0Z3568afeG9qekjdfc+3sMI0UPkY5xHEfJdpN0QnDOaGPQWyqyyxw+51LSFQc0
9SQc0VWiXmfzSqaMuwn1z8HhuP3MNxcc6ifgD2KkdDXQJmFgzKWEu+QLTLnlNy6EXA4zrKmkd6xy
SM6ZTI/kE3GLzCdh2QHroIQSLughrjHukMxvWEaGs6bQP8bwyAVW00gS3ex1tLMldtccSt6ifnqN
oJuNmPMh9f6eKg3a30VL6uVUeIXsrXmfbpU5InhbKzgnfdh6Pdo+Ip6RgvSLJqKQhV7KOPjGKwE8
ZxmAqzgvNXePnCKtPTJ8uSm8OsuWQbd8ra0iIrF3pw9lI1JQA9XDBlLVKyxTHaj31Ah2caK0Y+hH
aM7jP3G65017lf2oX79qxRVpdl5RPUr8VoSlC5EYqOSD4IEN7YxJquIB+/lQfA7YWMqyF4P6OSf2
/lUB/Bh9mvlAMusV/3GgBoLsVF1T7oKx5b1trB3HPISNPNtvGXmqGWhuUoJYaQAom+qu36dyW4cI
ZKU2brpqMzMpF7xxV4Px8An6azjJuzYFr+EFnu3zmxJlwc4wFOpKwNXaWwdnRNW/GTZeNMEzpceG
sZ1Ni3ecB4AVNB3xdSg1kaHYERuNGRNZvev7bZC9q180aYqT9K80TGVB1ykV8zKIT8O9pJpS+cim
XPlSd6SMiSTM0bVHaPOswTnwvGErKA5Jl0EcrmbqZ69MXRwVpZUbF53SnDgOzAK32eHbroZXlqhM
cQglRPIJpMFBXFiFv/e36ztokSL7K2q7TftM3U8dogmV3ml2QSXRWwvh5RFt3YlaKqSQO4RE/6oY
IMmmAhp48WxBQtOgZQHXK6aKGFpkODspgC3W1LDo03SvJ8AfWYgFjiEM2ODGxJO/Ylek/iVZv3jo
aqCO0REvVpLVmJQtQzqeZtZu37AH3C8to6gCIi7OPUK9UUgnY61AjnmpJa5CMinrFhwF2ATBms6K
9l1NTOFWV/6OOrcQscRMgN84yFqa8ETPB4cMNWlS9v9aHlbrpUZnpfFAxSMhM5j/rkjHRlpM77Mb
aFkEWyNLjE3D4GEGXr1Ovk3HDPrVdgTui9D8XR8vcr0JZJ0hBGkY7n67aU/KgMH//19KyPkB8J2b
b9EP6/QDzur0dWvXp8ojyfB0FWkPuGY9J1S0HpuHfVFv1ACLv/wZbH9OfVPK7MsZjDac8tvEpZSN
fVqRHfFlOkt2KASncb73nugDijxPa57z7DyDgq8Fj9pdC4IWgM7Vjx4bX9FIpsv7/xisgmklXCsp
G1BJXMR4XHcmPcVM3Vufi97D3htiZC/fVV/LG3BOVT7CjlXOratYLwNU1gN5wunVQvxhJ+yYNlfc
GAbuJF2R8j8QYlBDobOStz8tlEr0G/kO//kWXSJkoiTj+UcixRU4NtnIq+btOAwy+gkmkd/u9F4t
3/SuYSb7aYENYX12qJ7UFm2QjVvkuECjyhT+5pLCuE6dUbJtydinTGkagkDykMkVA8j57Dow0cqf
h62hjFfJZ0bxuYWVrztFlMjBqYZg4HgjeIMZPBA/gQ0ClAPyo3BeqlfPmBDmmh/JOaRItwDvM7kv
NERLRWYL65gfZrdO77jLysmlYoiKuXNQECtAhuGWHUK/LyOCoxEWQuxb2SpdX1bZzdnmr/Kwf4e2
FTAnGeXXO/l+ra1zAz+VfiZJWJux2bF7Q5srlYNU+RjCmhbKPFo+sMIOrFD+1CAz1sHgDeC3Id5E
Wi1EpsNbQTh4qtv6JoyJVhDFk1OqWILuk025a1VnXd1C+7MGmVsv1Dte9AumLZgEWEcWYnM9KsMA
JvZhjPxNEGyXIuEZYaAq9KT+Qp+fMlJHvMsj+pj9U+0qhTWP+zZ0+3hveeSslXb4KEoxNgZWZDt2
+WQMWtJIQUP2gsUjl80VD0Gc/Oxhnr0vQ9rPH57SOpuHAz1NRJdKoKSGvabKjdcGt7gqQssJ6pAQ
KPrxaNiaaFPYIOH1zappSLriBgcgQUdII9yiJCyvZVrFqwYom6P8vcmpe8JZjv/gO713S6BCVYJE
hJ62K/1vrT0AnYaiG5+yYt1HLYtJD86K3fPe0Mw8UjJ6kD5c/O+Ty0TeV43kmZpAcVbfwoeAQi2R
2QHV3Gl2unqOPBA38MfgJeRfuv4fja5JjHiuA9I3HCzQbz9TS8RaNfAFW2D/xD73SBkV08scOBCt
d8CDP0o6dZM3h8Q0D24LPhHMvQegPhPBpdVTQ/Ex16v7CVoad6HY0sTLMkN1tpBJo9kr76c9Kft9
UUExbQR7Tp71QGZOZtrLmAezI62UTjHn2I32zBuP+2IK9TEII6c3dRJIxym/slc+Kv/qUwJp6lOD
PWaDurwZFI1yYUgFV012vJgnh0WPs9Zjw+5gmCOyRSOyqqGBvKnrP8lguawmN3xgs4JvWSOmm+cu
bwfnkZNQcZPdFz04DIriS4vDFOAuR9nDGgvkWl2lsxbN7IllMpSvDxbIXzjgFnHdPcLKAP4t8OxM
uDfPGYWgJwq6rvKRBjeh5fjFvDACJ8PBzrdXbHVYBZVKHEjVkKJpg+CzZc/iXvYHEW+pdYgBmrmP
02Fk5K2aGwR2GBLpw3zqxIZJDDZ33bIQBREB0RNma3JaiqqtXtiEswrl4a5buVN+gqggbCH9Jusn
4eFooIsuxI+pX/mJC69LGe9hNQ98RdklBRSbgE0+bBNMhSzYsHnYXKuc9y+sX/Iu0sed26K7R0d/
jvJ5tHzjLie2qfwIyEq+i9cHILeV0OakAcP2jgux3i400PqU2xyaN+Lz15LLYBiE3tNv76XTadiq
Xdh7RPNpOm0WbYQThX22Qz8RMTMIvGvHzfldzsjYzYnjTwQ//dha+VNXbD2FrUkUIbF+uMUyMy8Y
p63e1T6oN3RR0nc5heXDYV08HO1AfExFd3CjMG1AvhFIs/TEi+pjALWiqaMokSUVaTKqzPVtE9si
gC8ZmEWd7XQGlbD5GIgpbXcIjRwA1Q2e/+rsqS/8s/7djP1gJrwYx08sTCRK8Ktk1VNpgSzJaj08
qkraRzrjmvtSY0X7+vjawDeWJOL/Z4Ui+OoiS2PxfTtDp39N16YO2invO6qCFZacNkIdrFOkL+zL
wp0yNQd7NPbHqx493phlDNHn3DOotvBUL5S627cUOZ+EeEwkQIoUPdZygwfeDWXPFKvKZAyPPIJu
qb/6VUVtZAEWaajN9UC4lJFLtMCety30KLDv9vo9X1JtTesvzo+oakZHYglWuX1OXJAeiFk5B4cZ
3JDVTYWRpNOAjb9ZBxnoKwkRnKZSBkJOqts+SayDanRQaG2Q5mFtAKtKfoI3pyE25xNbQ/xKwfuj
VyzR5+3aqb768VT5yb1/5oPN9+M0/dQG4/tKJ46XoPqj0kGuWIGhSb2Uxc4ou2rgg2EG4tfAbwaI
9vIm+v99OUR686uvfaULJRigZOjqD/7HFyMSB6Ml7ZUmVfOUKcwPlqjjQC1JAGCRPgSYOHJDH6ty
SjupTZ+kCMuL6p7Uq3ycJ2Baudwk5MPGzltjKkhNThBlxx7KtoT8aIdGK5gqkdDfPGjvgbD2YRGs
sUZyLmpBOGzDUNrHhDqc8zATignz9jkYSWo6DCCgEl/GrwzkMhJgjDaabhgJsVDLds1vxaOTp+oQ
/t9dZse4q+M0+QQNZ+cgOGk7UQWz8xTBk/bYz0rkFbbrun060Wsmg0WRoLNm6cUO65eboQMkUzHU
qxqni+qpHZ8Cn3hR/ohO13XnsujdjDDLgVjYkcyOeXPp+UL8569Uljn01xoBykXNQNf4rxHqfG+X
PU4SKY4KnTXw8jYYiyJnM+AyyJd38nLMIUaYaQYMNxCs0rPLCWyrEaO5A0vCznEQ1P2WGZ6XOXv0
nEostuLJ5WvlxUYaT5X3bkVPIU3RaJXCXie69VevVUP5N6K5y0uOiUToJd7+aSD7scC+ClLfd1f9
RMeOO2EqkmYI74v30Z7q0YwbvMXjibQXnxykehbGTn5AB0h1iyjsMMtHktdI+D5oMmds4yomoRTF
pIvMJg+ae27q/SMy0MEhObT5vYSP0jjBvQ9lbqcO2jQNLPIk2VAkdp9u7wAWxJR/tzurpygiWmkh
x4DgSCLaCVuMqfJIgLY7SJViQbmo3YRgXpfnWSDOLirX7FwGysl36L1KScMZN2M8S2ZW1xHlBqws
C2nJOM7HAr0leLcWN39MAW3+CYIw7DpiW+YKTlkVppSq3EB74AcAVgRKjs44ZK3xC0vyDe65xAea
Vtlb71KY3cjA16dXadAyI7wGBSbgZzyrnSm6w/NKzT1gGr/itBKEQZfPjfuq97SRPeglxeSmOhmu
P+XaiEoU6sXvWOWeWgm5rjsQwqzBSZz0na9p6t5w29QIpFnVCtoIxpG4TeX22PtvXJXBZ7HY8LKU
cnZH2LMlIL7lDaZq38qGc7EBnFlBX/Q8c2eZaHwXyEr3yqUAKcVm5934Ssnc41sp2WOj+6Hsimba
nI/tu0WQiD329emdoVaUjzYEK5KZFpknZclmhuIoMgi6cL33aNsZo2iCAbXWf34+Jfr2244XMpvm
bJL6iHmH0l5va/NPpKS14l1u5rXftAwQMCKZJwPDSvDUhgtSNV2ukpH31YCzLWwf4XI6CryJXJ2G
pp/ZWivcYrzZl/v1ia75fnZaO3YtMKUjO8NRyGrZBYgW30xFXq2VDELOxLIOW2+p7QObFBqxR5bA
0D3LQ6vQDSxE5n1I7zgywM/TX8NUP5pvpwBvjgua8UdCfCg9H4XzXW5je81WeulrnWfAJhjDZpsR
Y0TETtIXpnhRujAOzqIiCOzeqiJwlqgFRvkWCqK6/AvqD/VU8OtjSQbk4WZ6cvawvTFuYth2bTAK
AhRFIY4p8o/SCOQz0kPn53VIf0cqG0iu8a/vptKG0hZvqQ7cuA714rEbtDx+xFq47d9qo4OMoCXm
5fXCNTb/siuK10ph1QDF6mNycxbtPEugb4Qbg3AoHJIkKaqyhJU4H2sFTGAXw0T+zSSuVMWrj6yx
zzLoJv15BPnnEI5Zm5WadP6npRP0hiOh5Lb7xMwBNzVOjANNzC7w7TjnLRIa2K4plgnhVw+PS6l8
13kU3TXqG/sD9rDaX8LAyyzl9ZdB46M+xOLpTIhKs3qnE4tUjnC4qDT5DMNI8A4/HouMBk1T1V4P
KNFD2SAUTaTt1vT/DCAfUAKPx/S/4CMrN4dWAVlttPY7mj1Ldok4bQXLyzkd3NeobT+s+yxa4M8D
7A+jN5X8MBJFno7CLhH/2jWH+oEbHUsf7PjLA7VYA6CuC2A6jlQhNS8VvEoQchWsQN6mIp+1odN1
YAHl+F6+k7r2tnCmWmWmoQmP8Z1xjpTUXOfkbJjns1S5QN/veuoprDhae7fP2TrGiP9dnEMv6uP3
1XGLFsB3cHXKZrkvQ2R6p2wAC8aGBPbRNKDlM//56zl3Xm5FO+QfktKRdI7SCDUoERyNQQFhDHaw
qf2uW+oGWgsAwp5N5ERKl2SrZzaqZfxi2ggm20gOvoIzz3b05IYHraV2D6A9aR9DDpD5IenRHLOX
wnWY2Hi5XS2u1KATTQPcHICqPmVa98AvC0hRceIwg2OyAeYY/VvZj1AfpGHtmAuoaAfNksHbGz2j
tfT0FZ5xjLjf9P2rmCd5KJQsohGXJ3vWPiJxb/BIDzdYv8V++appR9haTZKcSOzvaoKtKs+BUwG2
dgcVBNzCG9kCBFF32F3ozbKWFN/GATiHLt+kCMw393/Rrd1E1MxBeYWnMDWQiOrdBfaLlBJcfwiB
Kyc33r9jLCSVainHBf4ZXcDuVjd+9l+b5IHfyx+uMYSEea93SyaGFB3WKhM/URMPs0Egi9kQy0fh
TkWPDUDAAxM14eMnD56fCC51H6eybgXguAoY6yTL7MRQnaBSv6zduIK6v+lsrU+MFZ1LXTbe/Fjr
OW72eXPaLI6mt7WCFXim9zX1i+reJ62KgARVnSZWwyll8awvx5zznVXOYA1bPC9omHI0r7VOPT9u
3IY6YLb4Pm5tiqCjCZHfq5fwh7F4p2Xve2uyN/h+iTjlC/8bfDzkngHmZeWA3BDZFpbVHV89tu0l
C7dDxQqWR3OcHPhVEF3HKxd+XW7xZQUIcjp5Gby7CZkM/E9HZxn4/b0uH1bgD7Fq6uLyYsxJBgjG
uO/siRvK+1gi5isQdyQtxbl8We9Mos2hDyg3HI9pF5tsKi9PC6hOUDfowfV/2b6cxrDfdMY6Yt34
450If6/KDjBudlQRlk48+oxq3Vz50JFkCdLKpCgYUaQqcFlTXnmp6exTK/zpUKz4yA/NjdAnqhJF
PFwRgy+HlNQj+IGL9dO1x2AGmfw6cXGPc5M4zWHsgk729c9VwobuGt0MpvLWYd8SJl8wq7GVHEJc
ckyiXiIAJDuRV5S8gREN+cw+LCxOsfIZ2z36rx0hWpjXhXbG5RV2ujQoqWyEM1QJVTt+eJUwIYZQ
6g3UIzOUQKyvdzWtFWTCsu572Rj4PF2oVHOSw6IsVSfqX9tlcxyjMMCBXJDIlT6sEcE1wARyrPzD
Y2mx5yH6jWsAjVB7A0dSr8zxFyAhEalk/K7JzApQfhADwDSktacMvXHFkRnA2hkzS+W01UjR4/FV
CILBTvJMAa34RNa+ysyq6xBQH9yQc8qk9oBh760qC4apboZmFaPtkyfkCnO7sDnTtjaNHE8YtU33
7Cnzn9WUTNCkZETjtw+BsuJklhJeHZnPoTkEvOYoEL5Pct/Bei7mK8LEbjXAB9QkpEjtWJ9ekqA0
2Jt8KuiXHY2Kei58neC/qy+ZGPatPKKfp0kqjjqX2MneHfxmxZ0bbK1NMTcP1RnJVA4emYU9WIY/
aVAzvxVC1Je8BLNJUo2z6Md3+PoxJmaCldRKop1R6S/esWfUus4/JAT09lnhbOnKNHjn5Cdzi+ZR
ApHdHhLoKu9GVWBBBp/4Bvr68LZdTHxE6pjlM0rLPhKR+2wrxDsbM/BFcY6+LU4aepqkXP6IM2lL
ZCd//P31H9PYol5kKEtBzevmmgE7K865B1ZkTiOp58t1o79UWz8kZN4DGSU/gc8NThLDhgI861km
S88DRqw+uUSrupZkF3eDc2JeqO9Xy9hXObvrVJujKCjvPVMgbbBIuvymrxy+Gw3D5mxO53ryWKFV
4rDj2+Fmua1nQI8/iqiQ3Gyood6xSc9mtt6zkc97G+QcSewPcOaTF9Z2gcjDlanB2OODT1Z0bFta
0gJLIgk75ls+rZLF7Up2F8mniws7QnVDjGlPbvUs3bR3PwgR/6Aw9Zmes1KTeaYwKMll7mq2JTsT
4HbgOf/zSZLp/AqDxhu4k5aiuZcgLeiz/i8U//ShCyENjiYERbDVGv5mLCOh34uoOJUqKqNzIBUz
EcI2kf7nKC3ynLLTsoTSpYAvsXZWWIL8oLMnP/s6LEPo+O4Rr76ceitBF4rRT5+eSdpvHdKhxWvM
UxMPauXKUCgv1XKxyHwSX5G0SUw1hOkK/o/39M7Xf2L+/H1Yp/6t7CX7hc08M/1CCv40CcWt4Ufu
G3Pia4lNBtvhpuCztsfXj8XvDWusTiS6kNf5SWRlU/TNvGx61tYUUvSIY3kXm7abXVioHK9eRwTF
jJFmYNDXXe0ZTFVmAH+MIvi1xZBW0Av1+RNhGfZgstSUmuC2rWxKfJudWbPwHk8XjloctL/02zxR
HkIQf05k1qJqGrPcxOHKWUSnuxDoBVgG6eyaOJCfRvEgZRvziOE0136mLj+lXFYo8sRbhmQjofTP
8TNHzdLpoN4pB0eqYymEb0F63E2WfItNivpziquOfTF39pVkTE+RGfHz7R8Xc1rEIZ88BWkgbwfQ
tNkJ2MN/RCSkzSi3ze2Oixs0eJFLiGVtaW3J1Mfqs7Tpbw5qZOiIEscnuC8jIzwbaJ6lNAMUtDcY
ccx3GGAeXCk4HrVjWcplSp+XsntF9Dr5CVWkcNW0DQolAVF3Ax6RbyZdHyLWB52itlTkwpOVibs0
IZrPFrZlqVX0p1pkasDgrE/wZjs8OcAQodJHnQVU1qI5R5OXocvliuOOPocYGnBITk2s1z3L6rab
GPCLPGQOZfdspU/a35jBzqGoCtbbnJX5buTxezZXX4Ku5e3fQVDaGQDB/Vw7LVftiYQ0oWFM1vn4
bNAA467QVaUl3drGY2wpAxPJTo7iePXwGpB0fEIWwJgamTA8jJqQ9/RI1B3c/NMd7RSrCEmM9SXL
ypteCucBiUbRZgmuH4nWeejFcJLWSxf7EK2cqjhZzvelSD9lmr95a/RRMatusAefkbzzfjUPoKXE
lUuCBsDqeRn/p5nVVGRKUBQoonu13c0tw/hOzusq7e0XG01YBfhP/z20LwHxkc+40yF7/IA2rIcM
zQccn6fXe6meqvVcQK2LnDjoK4KQZTZXPVOZC+9a5cxnnXfxzP8ArLbJcQgtP0OcR5fCpR59h8LW
gN3Vh3Brxv623cRl6DwOyEHHRHpOKozGNdqu6iPpL6KRoKwGL3jUVuXIS05AsuBgZxgH84B6Otb2
KS0RP0eatdukjetLAxGqRVqZHzQJQspulV3lqQiqBlTek13IhpZqzQmDO9itgVml6PLYTd41oVcu
+PJ7t9aSBxPhbvBrTcMIYmviW3llwcFel+M5CEfBa5XIpkOxoT9Kd042/zq5b5nycOWPQht/YOKW
LpJ2hTxj0xzFxt0q35FheU1jcy620oZDootRGSXjDFUtb8Q36jyJZvfoEj5qIxkoFXNq93kXbODC
q8mbKR6CKqtmugrleRdpBALUmBESVrDemVCfAIP4wQT8BlL4CV8YWQ8mZUsd3iuBh3e9fmPPo2Ks
UFYoX8ghrq6Wis9vofKgJenxMgaDfJiP4OeKi+2meesjDal8VR2XLt0VKJrGphlJImVlpJfv/Nlx
OU4mGK0v4R9sHIX8LUfHhssSp6UE9HdPuJIV6KUMcbjAnpMHn+JBmCxjqHkkIJyvTSK6uiRkGFcq
xzWWHAnRcXZYFFzDvZ/DMOlaxlpRVcYpVm7n2RDqO4tMoff0d9L4JY/sp7hN5LmWBIqx4ylB6Vbk
RwrKD3oNFsAOVy3M6E/sRP0db7SgVjfUOjFlPTSJWJqLvAYXN1CkR47Nvt7Ju5A9Hjn/xWoKXkrT
zEx/b2+5Qa4zPrubkDdeSzEXj/vtqacJPADqS9oOLlI4S3eiOoC24duOAFIGj1uzSoGurNuENt7L
rlWPcskqRp6lJGvxAccONudB5nRXU+cNQLicJ8Wfcjs8wwItyghasU/haJsB06bwWJBa+4GNby2o
UwosCA0hNIRdB+2327MS/j2KMiKZ7zGYAdseLoJfxJKvBTRFcFxXU3YpwsiNdZ8GmulTEu7xf+xH
FKxUFFWTDAdw//MP1G2V47CLII9FEjoba0RGQwQMRNVZMWsDtEF7W1U8xj3vxn67Y5r9K1ekRO2h
CM8K/JhHADoMqWWxMwr9CbXmgem6I+bhw3q1iSXSDoV+e0x+ucHWmqm0NFkBOvS35M8Q7iMESsIP
Q+v3o4eX3AjofXb/liAurDpp7kothwkkDEmj4rijzya8g9NHXO5R8Ew8JPVIGOkoW18vM6TQU3Rq
Ji8HxJWYpCdxYz/79ruP/JzbQHRD+UgY9xbyoxQPYDG+yVZhwiJ4U3nHvwWZH9V+cYfKy84JyRNW
Z1VdHCSmU5rCy5uZOOWFrz02x7EK8Jb6mkWeKo49fmvMbtaPQVHO44NVAwDZ8IhE0xoERWQVbmy/
juB2tRHuIvilgfb/PcTwU4WdpmyGO0m3jsS3tAaInkgGabSIZ5+M/bvFv3jeH+nJP/172hyTGpmC
biDA/nRSp39g2VsSWeVbbmpi6T5KA9zfyM5TrV3X0Vfg4oqgfj5ev1lJO4GXIaO3ttBzOpLyN4Bx
ZdULy74pFziXhM5SLSyXSieOdOvb38lPORCer5PToktbj7aDiGkIXJQszWSyMtKOXx1w326H5RtM
rvDTnMS8i6RzB89QLaNPV7SMJCN74kCUZHse4cZrzvuRj4D7P7zMqdfMxFc7ZU8DJNomvqhxJEtZ
nwbXYsgkt0PBsAOEp8Q77+yRznN6Xzp7CA+pUmcXcA4Ben7uFyllH+cmP5+PRuYH80ykFYcGQCra
/hVTZ7/tssX9Ygn/A3L6HMBGs/AFNiaoLPK5I+N/KQ337XaBpZR0ChXDHNvklmcLRGXHT37pdbr9
FYVne6xxDQAAE2d3lfqQkXue8pYXmtmWyYDToC5DwOza4Skmmg0o4NvbjkY5KNmZb5W7cwqPw0zW
1CpHZd5eMkipLwy05H9mpsg04kdrh7c2iDOXXW72FGrypa2WtLlrPJfs6s9TK/ZY3DB/Pe0IP0Ud
ZmL3BeVvdtxSIYLKHqlUZvZE7fr738/BECCLJ9cwaQnNOqk5jTmgDyviNCYMwmrBlRsj4Vtw5Goq
X6cptX/Thwd+19auHpZ+ImnlouDraRHe6BzWaTuxmG2i2zvIrdke98QRV26bj8O7z+j2la8uYSxh
bSF0Lm2dhznOMTgVm+aFPn5J/fcaGLoV7wDdnlORP939z5z24c7OFYLrR4L1xYE8haK7pzIbkyMd
5wPZZdN4M89nEF/BwORuh5yE9Id7bXVXoqb/FegxA5JGxMl/leQ8rlk0kdZceubW5ebMVWqZDwvJ
JLt29KZN9iMUOYSvsNN757nNu2N53FJlbEi+p9CI/E4VHGBtJ3j6daPFgUaIMUk1iTCLMSnHITO2
SN1WDzZ+MWGq4rZzM4Eb/lYrZtSCpGHhuAQoysB4IcBFFe74aIaGc1PpewvlCmGAWQg1aOQ0dsVk
kaiDp90tVIn9taXUnWWHQILeGHhJqlMzKrR0Lf7EPIHNmqhET4d7CrTwlX8seqF7xwvdwrNTsq+u
QNht4sJTOeWjPhDjP9ggyuj6eenFTX4PkcOMHfVag2vLpkUzcaqlyfple+tamjCtxwko5j7+CYrk
4YYgeE6qdqaKkWridLpYkVWKqSzk5RWFXo0hUt7drrZThXUBZGy/Ln2a+WuzxoZYQJQliMF3w+L5
/MuvFd7rteVw6wBhNJZmi7tUyIEBiRsg+gvdCjI5AsBQdJe2EXv4Hbx/f+fhEdtFNt4NB5gjhUbj
42MaHVywiYbZa0gWeOCZ5trnH7g1diLLMTmCyZ/6lU8zlR9wMiyhb4F2G9cHvZOCCkQzn0yF2sMZ
RX7VY4AN4pRzXkcst3xhHeYg4OoepaO3I3tQg0k9FMHxJXBy+f7WOMmnPzlSBzNUbTvlP9JybUD8
n44+OL+Mo/PzuIXugHfVOoHA7QrnDzGCZ+dBhWbhfVbAZdfl7IC0Y6CwK5HKGv4i4qm6QUzklaW0
6XhmPTRUlIfu6Gz4fVrZ8ZnVm+HwJddmNH1dLt++rtJy6J8L5wd6bYAe4+f/I4CktNVpJtXhcfqn
/TxbA7JiSD1bKGNabYPxLGWKATnx7ackvlTebBhOuTHHierQAcZomM6LG48kyqK/9pvWUu9+R4ex
02W9lfkKunOkMoE48LP+2xqy6Mp4wd/P2+qvNk13SSFYBEM1U8Zz/635+8WZsOs/xy035Pi+3fZE
Ud0zBeq/0DoXuXq+gRd8VQF5fRevbv37wNxF2Tn1yPGGbxUVt7yhdP6yJEv5baykCHijiUHD48cr
WCKHL/yAOqmXFnB77rBQsPjOll4QBbmiVX54EefaNOx5OnCzUIFD6wtBSIjNbivEOgLy8L2nrBgw
/S8uDO5UtPzW/psxU0pBiymCB41btmrusuxWTLxjzq1VQLq1qfj9PZWi55Qkgs8DwVTaLPTiJnFm
93a9fBsGnWBaFVbjTtXhxiodO7eS1NY41+xQzbixMGXsgPSTvgzshs/iIWFoecKGpNpDVoWlYZdY
T7BIzoUdg3+khG9GoQ94QKkGc1WN3ZHQQOYnngaiEfSLOKEgRrP8kfWjx+mTvX9ORwUyisuZkjHg
H4bQVA4jiPBoin8eP/Y6i0qshiI88nHuPNTxGLTT9lz6e8jX4Xu8hQCKatmf5719Inz+LIwkjV3N
Hz37PiEk4CuqP84fOeDoLb+2Zf6rdiedo6hFp7ldUXgRKwxb/k5dZvw1gHcb8eCPN8kQe9Cq/KfC
27sfrXFgdiuZzvlrxZXbIlorgMB9VH7YCJQ5f4beJNT972zuz2fCFg4LoTJdTuwyrqMJKndyYQaF
xmJTRmADpvLLaE3aE1LWlBgzRG64DRdZqWE1U24fJfO0O2D7JE5Cc4IgI1gz9XggUeI/ZWj4TLT4
C9pjFAWlTkdr/RNSRfKSPJRKJ0h0iM/1YFWkzZsRK4KFfvG/PtVlbdd6QFaVpe0Y3uaxY7DvYCTS
myqVALYmSdQy4Flf4YljJgTKGqSgOxU0VU07RCCoYEmeLQGRukQ2UzIinmwqsro23wAlbHW5KdbI
mlzRSaKA6ciPHlFLzwaoNXDkRYy5YtELkHWeh96wZaVWJKFbBRukrN8g+7jOH2OcqZbAnR5ffdA4
BoCeUmR4BdUtf7/phQh/bBdSiqiUrpulrRRW5Tndh528+TAqChE0CV3/OFvq05O7nHv/gcheyMTc
j6gBV2LU4te2lnDEmbtPNOjljzlkf9JVH+7IGvK4bEUT1nDegIYhrAZMD/q1qCsotJYUBdEKnlx6
Fxo7WpMhLZ63Ff68Rv+A4hG37VTZpUYCPVRXVzifJTsv1KcknBYHOfrzE7TH0NroonGWye8gUK8W
ZRkXuMufXQE3eBHD6gZ16nDe+YgG7aahH8vyLNs4rfHj7ErzeM0x0Bpay2hXo/HkXrKjrxPxfWA0
oRFNCCjG9XzB8kmuwV9Y/bbHAiiQxAVPzjrEq/zw33T0Z7f7IhqNvem4jO45RFdF71w3twbpQ/BP
EJKDb8sYbI4pnuVWz4eN04h+wp+8DxanXunbhZgkq21lkOtq0QPXgApDRjWuYOe+s+y+r7newCOC
eOeqMpqqxG40CCijYj2lAb/3Yoceymb2ZwXkKfZf6xJHOZ8ffCKdXNAP82ojzsYacPKjdXJZ8vh/
TiXLFIOqyMlRLrz0M+YFYJwHy75tSD6eyuVdNFIBvq/QMVDl+R+4iw7hYKTZqFaj2+/8gDCbpd4G
MF1ZdlwRKSmYx2PxmT5UNYlwBBvkXqZKfkpfZIJQKASt0A0Fui2QxZrIacBuDranWbEELCrP2Fxo
7lnb1032/2TVX7/HrC60y2az5Q3CM/pY3vhhoCoUburgCXXfYNM9B5ejrDuwzTpZ/YF+euo8J1PI
XZA5MX1/H4LiM9CxuvLM7KGe6WSXsWsS22vfdtbYTEIQ9+lTQcTmOP5xmPCk/c9K5PXhHZRBjgW8
LMTJPwivJqNfORXp5rSu7ABWjwV+1WW2omctf9/QRL6McRdG0uLJPDP3q1nQLeaaERxjS2YfPqB1
enyQC2GJCe4ZwcCwq81NTDlGxZESgnFpe22lzkLRa76WkkJ5SNOBTzcUzw6kAd5YLSn8/J5x9pIQ
Uq7o0sGxMwSunF6x3rgkbdFmX4W6PIfCJ3beEceM9t/t77WbifxS+cUF9GOXEIkMeguBnuodbEXW
ypxiYYUTG2fDEFiEh8+S4KJPSs/1ONM16zI+ONlZTgWyOxU4mV8EI+OsDYhgQNqgca1XB+WVeXu3
Ts7UOBRxALyCF0gLDrjVtOhdG5ekDDFgxdZgViGTBLbI4rT+kEQDBb+5A9xu7srSfOJE5a048WZb
HDemkFFlSl8vI3dRBeOKCTox4GD3adDgBF4miBCi9hNH18/yMcWRC12LACMlqkeTtFS4vh/Hrbom
Yf69AAxMoqM8mRQpJ1+JqsjcdqueFicuLU45ElFEtnyp8+rWp9cXkV9YEOQxFpJdjUcPIuwuRZm1
NLpSV0x4+ltJGf+c1PXS+Kf0QpJJer31m2C8P5vclwNW/xaYeqq2qq/6ohhzEz2zz3H7L1QXDjO1
MnNlreUhqDQ9dfX6+GkjukCvXcsmrr5nmH9fjqc3BzFoK5VXHdvIEw0BAXmTop4a004m331ZoauS
HPvYpEGVwJ8EKt1ZNXbYUrDz8x8CNT5TfdiXPpLXejzou8qb3YsA3TuRCsP4vuJgDA8oeHq/ANdk
6+O1CZu+6LSSfsY0ShPRNKZVJW4sTYQ1eSAKRzEmHU6p2RBilysKMIPySEY5iG2+/CqRbdygLfEm
YAr//kMcazoMiR7GjOD/YSiadHmRfFastX+SUVTosJxcEE41hW2nXkW8q1JffXQcVPJ5s42lIcuQ
i+hm4Ta/RaOMCcZUTh37qy7Osa3UBZQD0Cuftq2ZE+fAJfWi/xKLBTd1FfbbZfs+dVuYcbVEqqVd
nwyZ9g7oLA5PY9QvEDOX4E6l4zy/y0n4iBpwVUzIB3l5GrGUXu9NS4m7kVaT4gyLSt8G4euKypEz
iHBQnQM9RwZnyLwgUxQcDgnNfFQIUBb8ciXQEQXAjmznSL9TFSiqx0umOGBXVmUv6NVlvR47znpl
dxXGK8UluDgo+lGgp2lyH9VvhUmFcIwrmj4b5Qpseb8DxTaPGGI4hG1dz0FvIeDfTRFdOCTkoLYz
QWZuwhzQweuTE81vjVP4oTE+9ye/lZSQdNKPbc/noJoTWC5qbx3YHBkD6BMvBQXiAaR9CNilqhtc
44AXVe5MIt5w0B9AxIOFfBlcqaZfH4No3nHeFeL4Hqm/YWPyTgKdPevCtWMebI+d4R3VVqx6M375
NXKUwC+XGWCS+KHsh9PHbXs7jAHBO+BElCO6S0UiQ70rzDTOy3GkyYKdvzagHavpAqUyv1lHWKxv
FkWUTcggbDIEshzOpksqcLxBpefd/XC/OYjshLcJ8Ly7N2Mg4DyW4Q0yIeoZ7jqdH6GDm3t/PRG7
tlg381dc8meKnjR+eemzN/GzeERf3TktgdrvhrNmwcIX9DZ5sgmy3/EnTnHwfAP+MlvzTxV7gQCc
yJNxs3ONMGBRiI7zNOMKsqRXhkjA/zBrSoT70uUTReDCnjQCacF0yLMJFIKL6IZQgxY56ggDe3Sm
q7HDSAmZPtmwelu+nZmADnrmF4Qc9hMYFByPIseZRI81ojNiS3Tp+kpqiy0sEFck99g6y5eV38Po
BEKDR0xFHzJdh3Ls9TTNn5n3uEbTY3i/+04wOD0lce+iBJasKfSHpGiBQ5QqH/wL4Cx/pTGRdvcV
nf8qTQHfuHifdWNyBMaBF3lUc/Wab/qteh2fmSccBB0KWEdtupCoPmJD+BNy5kWKm7jfowQg3geP
e1LP8rLITzG+s9WDNk//PyT9cYNFWsFmkLojh6gkpkhVY4tAOuUvNtr6S9jDeANoibdXfDwLOk2P
KgSGlUtHnWOSTBKU1+q/Eqt7oJwH4JEyYNQrcXCH6rCZdZHBi4aDQHpsSv3p6JniYyeFPSe827B+
6pml8pZEhn1hw7YfXlDqsjmx+H6B9iOmoOiuurHwuODELqmFYcxKsrMaLJLtK+1R9bW50/tv/yEC
V6fVLdlTNUw/3PxShWegfSnSC2OpBfvQDfeKRZOl32OPejUo2j4O7ZLyV+B1SkWrQKnG3fK76Ma4
Xh+KTvZFH+A2S2vzGeNdVQJyi3/DOlHFl8ayEdtotLqHh7zgSwictMwYxX2l6JJbSQ0TBBcZteS7
Jx4XlWPswAoT6KEgS/zqPhmDrYZKbLm+8oEnvqrrTXHuyxIfsJmEWyLrUXIbATimFK2RsB182wDj
VpvcefxVqQV468e4kQF1HWftkcziT1BaTGYsy+txfKTHISseAs2dtyiNcGvkyIU0nPnrr2iZ7iCV
EhB4jhZI+ZpGxF2s5HweWJcP18X1vDTDaVZ/pMS3/K9Iz86SPcAuZ2WRMO+2GRtRjql0kgO0ynNh
pGwkWy8rVVv2ouWWSV/kv/gAaXgkC7BFortvqgm6FoA1Ny76PaNyjHb0nMnUyZ1764sB3L5R9cav
fqo7hurD11ek/776Uv6gCcN9OVcRR51jZ8MxyG/JkGMLrh2xRq6ROE3KNmHTUqSWZXlJqxYFVmdj
CkHLoBz72GoSTS/py1ADR61JloqXcclUcKoc3fptPbQaF0eTzfsfEza772crsavKT627KHvT1yId
qjM1ZOcu8zJSfav5S8q4HBK/VjDOMHG48NekHexWtoecAow8osu0TtCAAJ8jwlX3/1/GkadnGgzD
PMaUoYpLpjGjwMPJ7uZNeOyqmPmFN5G1G4h2AAvJK739yALMkwXgZnX1rnGk44TloIq1ZwLCb+Hd
4ePBugID0yjnpBpaEKva4UL6nxXgI6DtaXEZqpGFh0tGmKX3QHAuf3Boc0s5eF/XERxJJApMTSwq
X1iweIViHMZbem9xbQc41uYz35Xjg7mIhtDVG8YlBzIAJyD6gi9wp5B0NwuYXicXSrqws3Y2AXVb
TvU5Iutvk71KYQnZvbLw+8FTRPs1+uST+/csz9QzRI9UKeSU771GvDCwzE3JTlApaEKY+k2Guz4s
4gsOtq+eywoGFXvOh4awIhM3ZJwGgOpEQlF1aUOCnujnOJgUyDPZzU39/x8ulRwun0xffu7JWfiZ
6ccMf5v2Ub+MpMpjdlXHe7GDRtn99y37PvHn4aSaGVIug4z2WAkAeFPOKBwUUZNytbtFof1A7GvE
RH6RckJnPTbyxLPr5KfHhkCVNtJirHGPdfJ2wT1sDvurVYMDUmJXlVpyE84rWCDz3Mqgbd7Bn6ep
t/O+pb3cilCWqL1tHnugSkkHv1xWt6Y01i+pRCR459BoS2Q1cq0FMfaD/O8L3hejk+uyCZBWwnXh
bAQD4VnD+9MhG2njY6Qjpva9wOTNjan26Gt5kZASWHJC/JEFxKj/gsi1O0ObheDQFCm+FgTKFiyr
Kro4gg7/UIlPwy0PWL4nYsweu89cfJxOD48virDyb1X+mIwjhL1xdlC4Lgl0K3OkC+53IcdRMcSW
MPxOQxryHHHPxFvtOOy86FEbJaWtnoXoLmA5+zxVbkQAwKTLD7JoGWhSxqJOJa1Mrd7DiVYyuRHK
zM3BEXDaNJWvdzGBYXvgdGte1nmmUALLCR9R6VUWCbDVBA+1SNvc/TumgYuTE7GjlVmZTHzKIMg/
c2yILc1Hooxo2AsQ42Yq2PD/gkPeHf5/DtTSWI3vK99OYIhICC0IE6rgOHn5H4v8dwjhUp0xnm9k
mwUvdywXp/yE8Ftvuq8HZsnSz9R6DphEUj4baA+1zdhWKp5HYbd/P5OjcwgAcVSS9J4VMx/biRuk
rgoQ3vHUuVjB0nEKN+qM83PWwQOTZqIPHUcUgvNGiSx1uIC8h5t0qUouBADZz6ytG/PzJoQRimXa
L6yu71NtH2PpDQRj+lVI57ZW04nafxVxgsXEJoD30uzh0ekPyoTwDxEx/4wn/I+GcBdVxeOXhUi6
4pI2gcG0hWUV+vE3B/DkNufyOMnxxR6889AFI6z9SZZ09YxRHpvh+Ebw4e/UQUK/K33HnqNUtA+C
t9ls+GeIop6uAdN4trN0YrOelIJ/mH6yQ6DmLhEpDlRcE0+jPddAhiG7QYC0Dm08SC09oI3iqplH
/wwlIz+2Ja1PCkqRnPnOJK42KDYkmJa5a1MApVZcGrWW2xUC5eg9jl/P4bECbV0hlWLceElnQWAc
PhfMnEn7TCxfDAfW+QrqxbtII8QojDMcLSvmtzR70Apx0Fotgmmal6y+LwLYQpdCZSLsG+RkPE3w
i2f1fwuY+W9Qx1IWxPm75lVRtWSnXri2ZJjTjUV6mzEzvLrDzncgJXHE6rWjBCQVYmOKCR+0COtA
DXd89utudffBvdOL9/RMfyyHJMCNwlloK4qehTZMnk0/n70Ed8MTJ5Z2DFdefo7W4Z5S9PCG3LMR
pwcFOeqDzodaE7oWVMNFPqL4NcKxqKJIBpODbmgyYmMyB906E9ytI6zkko5IfLJJPFzYR2bd/J5y
slCBTKqfZ3gRFKAKxw3nOLSMckl1mF0TLuVQWm0+MuafjIqY+BgxGr11P0vD2zEugvwY6ydpTrzJ
AlTWilLPyTkCcrWb7eRtMD2d5ctytGrudEhQbcVaFlP+ue4RZFItzE0kNcTxd08NsV1w1xselU9E
rG09xArzIdLQSRnJUoFDdVKUQqwuepWL87dypf8yuBLi2+e8OWsSzuGxPIsJ67Dvk7R3Ycve91pg
5rc7n2/2jW+oSe+GesOiWzynUM5gHEUWK9i9/OgO5MdJVkZtrTBuIGW8kHZz8jkQfRvDRH+rrMeY
/e30Cscz6rGNMqlmlneEGFe4XVOFlP7J1hg33DpEhVC180XFHXF5LxIA2M1SjXxnCXP8pfeJNTjI
5H9JqlZ066wDk+xObA+5O+LPWF/sdYSTaC7SdtkvT/3czUB7TECGGWIVlW26B+F58AMiKSU7JKNg
3QpzdgYCZnFnMlRAQGT4Vr8L0wqMAmENyxsjx+Sd3kIPgN1TTXOqqCCn9gf0bLoomZ6aOZtqxsDc
qpcYGr+DnxVv+wcENDoez9Csfu9q1H4/d3NmmYBYnGkR43GbvrNZU32jw6pI0O8bbmrAKkgVelVS
SJaTpXIVZpWwIdWG/AeDS7nK8y/lUnEgji9PBOSPzDI5ORIB5QW7Ub4NN7P02XI1TB8xEOyssDFX
UqcL/9p8ZR8bxE78ACAtXL5YN8QTr1nQYGl4cepgD6CngFSsaSdN4Ci1kau1kAereiEDPlyhflBi
0RVrVOg1OYAHwVAsmCsv9y3Jf66vqZ/Vqa46t0Sc177EQBItELy6Lipbf/SeIqU5kVUNC25fxL3V
2G2jE/7JpicaTZt6n9gJ8fju9Hxr6FVvaacoUFDK/qJYLMdBDS7+mVNIOI1mVzbfaTTZjVfoK2ZY
NB+NzOnc/SU6kaurdjMaBMrYbx1VbjCdb14mvRSA00BSTJlWuKQQsATrV97yeTIXR/ONUyDTqqrR
eQiwFlmCXZg4pWbArdgaTxfRCvasO26FQe+/p8apPFkOXy/Owz43gyP+KqAxbaRy4rVnWjOWOMMF
DpG9GNaFmzi0b3mrq8bONgtjMh8x7fkJOMF7Arjdh4VaPIgD+R9DwcW2HkMn5KabzWJmjxb0Qcpe
c9IRytzVhBWys56N95Nj/zMgaO1iRXqs69QZe1SFQiESzbGodIFsM0WjecXkM8jVCpBjDN0E0+DH
IpR0Pt4icUWsbm3iSroQBhXXpP3LYZZqxry1K7CNprOi+6bqdAb00Mt5IARC3Hs4gIRAYxvTifxP
CxI59QZ58hRDpJiRKO6GQG+vbvkaEs+4Sj6l7JnGX4i8rgO+bF6y8GbkF+njquAGdF/a5MZ6Z292
ce35zg4p0CVGu3fbDj0QXm4aUa710Zrj5kdkWFdsZWSafkVi4gKXn32desL6kPDHWdfos/E8YEV2
JrfRkru2eDUgfDuf8zadP8GcYO2G3G0EBQkl0mlEnf0lzy7urvhqU/ZyE/59rPlvBO8CQmAU00Y7
nwJG7G++hP4ZpO/6Xrb7ov6Aw1rPyZqvc8LfTnZ64B+dQf1cNAhRt/4EEOeVWZFDg1hDWIQdeuFf
UpvpRxPxY5SoOrpeqRz7qb6uFskRB5iAqkD24I+URTXSMy2CWrQiLPj6Ge8C0y/xVBYZx0AHq1e8
6S+21Ls/5lYE6wIRH2Te2g5WCVc7wOE91O13+rlGqjkKTsGg08VJiJKtdctr1wmHX0obVWeHLEfc
5FLFsGJ5YYLK+xgJKKNNJEvOcFjeN+D0Blogc+uO9Wr00212L864hJ30UYgaglcld3vZ0Xc9uo7w
U429jO6f50bZ87miFx5jouuOMAOYwjnBkpjp4xVhwjGeexMKu5LB94CVOYc56H08xCGjt3WPNnuV
0AgW+Jq8Lvx0wpErT7a8Fb61VAZWnNhUa22Oiio1DbjRMruq2EM7EzMhwx5yDm3i6OACUDYsPB+D
02cHTO2JyS66FMmrqPQJzNPweDGg2VQQPI7OGqzt6q0d8yhKUI+iGKAWNB5Ew6hI4xKjET/53ANi
lOprDgvsVWx8Pt7Lf4HeJNLLZnVgmpvpN6RAyhOe7YZbHitKes31OubPDfsMpUNiTWBliB90URIi
qQpa5W7fuo98j5VZOn+oFkcZSDRNJisCKGmxPCWavOop7P9hE8Od88PpHnVUetfZdQNdYWBCaoGZ
2dhLO1NDAnLZllpchQkTUm+08kaGUrUuXHEjZZ07sLuDi6GIzZCjLoWp8Pcob65j4ubQU/RKmPwK
RrvBd+pRCB9dnXEfSZrxZVpSaJmhV2B1kfIXaq22nqPiwdE3+RguPHDqqjNST2x347zt67JQ0dZ4
qLpM7JrBybeb50+NgQztWj/WV4cCojJXVb9ykj9BoZr81YjBmmkw1dl4aq6x30hlBbKCNcgfJMA3
YeqZhTZurbmNfbx6DAaRzIAx3lW9SyMxKNvGZHuKtUytpYkASrzOOMOqN7cfIiaO1NnT2N7R7cPl
rI0zK1p5hoOPGCOPdt/U1JnccDhcs2FduFzYrDBOdwQ5c7yZpjKLD/S+7qJj2u5MfGNbgkYtVEXP
Mh+8137aGjDn4dM2IRYO3/+oUCQsvZe9sgNoIWdgEUW4sLCgOHYhhSCpkXuMlM6U7hpqCB733e6j
04d8UYXvMTZ2hxlfzAm21cSTsmY5lij9+l0y0lAGNG5osNCMWk/eo/UTtkQJQas+f+UUMy8hWn1g
hRAaIanIKuSKoOYjzBiCtov5hdmdaWIx9xsD/Zvu59UC7XtYGtGgFvfF6Zf7rhOr3QYLTStoLliQ
tjTtL9zlw0Ieoq0/PPW6oG0/ftJweGkpJLhpuanEN7nUvU6r5zmUhKnWcvwl/8dleL+8yKhY2SiN
D0q2sf3UIXScoif9wpjw3a4i6U5tD78WgXBAaGgwuHz59pLrkCo5TxuYHp9q7XAr5Lzm7+a5iQqX
EsMzf6bi0MNo/6MHuqciATtca+9NPtC5Kv70rm3sUbJ6Sa3l9zeeh7IJuT/ns9QTztyKZQhumuOq
dGTlKUcDDRs2kLw8LLjit68UbohaNYy+WZUktqsQ6pO3kMJqHiZ1qMZfi1/Q2wHyN7Ac69VAtzOg
Qi4FmH2I/I5FSvtFZdNB3YN8Lta/I7PFwVJIaKM4w8buzuU8ruSaDRp2fmeVPrr+V2NKMhshhltJ
MHNHd8zGLNFFsSYWcOifBBlTZhTOwTaD056Q6qRDIFQv2uo6oLM4Me7HkwC1dCWnKUzHjx03/bQC
2KA/XeicP3NaarkQrnnBsCJ3hzFybZE7krthdjGC31UD18KN0IBPIDzhroKeSsVh7GX8aBWwnczh
Ikt6ApFKS7sAecAFAOzh43vyQtFmxJJA/Yi5C1UtOsIwwbFJvs23mlKPvvtSHERxPEmq/G/gKCDV
KuwJglOGyoRl5MN7YoIXWxErdmpYxYasL2koOGlWnSMEeean/paxcb6OkAbaIFX8e4MYgx8w9tE2
wJ0uEjys0Ag77pCZyJH6c1M6AOwkStlXooUSOur45aRYZAZulX5fjp/WqReAXMQkjJnlIC5j5i6F
1rZhPE0r5YrnEu++ecX5gmBKeqq3ugCx1ksjQETP8Gm6Ipd0JnMMz9tMudLSDXsz76s7B53lbFG3
HxYnznVCUp/MhguRMi6hPmVHWdK/DYWN8e/F8e3PdCoIX+xYx8U4J6u4vq79iephXBASTRslQtHq
SyoBzCFA+PCA8sZJO4IXkMREuMOM7wixTVnjbo+jlYTH1Rx0As7GKYWiHA/uPTaEJcOa+XBtP13I
6svcGfTmPwHiULuVPt0K4uhIQ5tfC8G9CxX14EB83swaT3SGZ5CSwoLZJLaRCQNK93NSPEanWAl9
Ho11om1o4C33vbY8Rovjwm9LRsQZFF5BXU9NQuyVLjX6RTuyg1E0vmb+vFHHgbHsx5vUif0cuBW9
cE34O46QA9HiAUYlzhBMi1WYSckk2VrcZipQKzpENkdF6oFvmXT3BLv+rwx/Y7doVYbd4qa7cU3y
yIF4+zmWpWIClBzrzv2OO3vBTNT9omY+aMmYvtNAuSFhi4oI3uJ0JavN0Lrf/yIv36W2hu2x6bFJ
OLmEKpqqP4WoJjTpS2ANiO47To37A5uGkJkJbtF3FvekMDIqglpCL6xem0dR17HG6wn/J5lO6aU+
LRZb3NZ53dSqMDxI1zjvvDHNyCNXodMboFNXLtL2TXoPkKB8NPLkud+KEjfCrB+v+/fpLWsY9B52
HHS3r4rnqUdCLDvx3HE+PaPE3fPAMAyk5VaF33SRHXBS+jDzMLpaRv3Z+8exkyxjqwIwplHKtHSG
wKLYyd5Qd6zxgnjaCAQLR6QyfwYZdxAdp3LUVJheAs+uJu2et8FX+KzmxO3TcAGO0IUFy39mXgsv
p27qXjcgjxZH7qFF98gYqrUtzzcRz+oA3CJG9zHV0ATN/JI6Uvk1WNo7WJiORpHGZWz0XBpHBtsj
aAATYI2vkcl/PWD01IeQps26ROi8xsGVNHQ5J7BrRYGqrokJvvIqIkzE6St40nTroAPRwPbFZmJ+
tTvjvX4zNmWjSSKZ/lU6z9ocs1wAR1qu7NowukV4p1GFiaxTXHnuDbj7a0tfQFtQdxnpy5ZwhJHQ
cPq7cD4QI0DAnyHb8aJ+qd3yPugt2SPZHcz2rMTHMgMrivOpoctDmSdQm1hVR0hXXzbarTUq8QcK
35Msyqk+JAHuKi5Jp3YgpSUhjz7NzWA/oqimxUXTqeLByOvJsDhy6ySUIe/ZgfX5xZQ5jDI7ofp0
bjajg0s0Sv/jpj3vwVqdfJ8aejQE4JS1+JMeXMnTijJOaasFGjExMjmGE/xdhB1v5fy/uT3o/k7N
oL/Z7elk7x3ZeXY1erBHjaSilLTlUeBD+lfkMy+DBm6uHrCmi+un+eb8wjPiOaaX8Cf1CtGaldm+
nyMmQNDEuYdWKroABt51N/WzeZ5wtJhr9yyirox7hQA/AgjVeErn3RdIh6LlyzP9AZtxYt95PNN9
Mm+4elmExYjPAmTcQlMYQq/IjZDoR+UgJAwiYDWueSc4yDteJnAxEpgL9mbeMtp6CcM2G6dxZPS+
7SmrjAHifc6a7y2k66AGyqJ9cjXxcHFK0ajDmkZOeFA/E1fRjs0rqHQ0VdR5EA8kx4SfNX5w0Zg1
SyNMN1lVgH9AiTYWZ5VGcP7YBhlw7IlbrBKYel5jk/+kWsGaMP1tdTNBYDyEzXLm7pXf9kEnxBlM
4q5bzTWCt0jIa5e8kFAS5pBpo+FsOUfkeM9YZ/wB3IdO8C/Xgs1F3nhFunepppnTF8w3wwrdIScP
Tj690qHc6TAlIUEXHqe+b8u8V1c5UkGl3IS+bLQYWRdeeIENhmgdop/dytnw+Fqb8bGzs86k+CXd
1l6Zfq5smMpLaHWjoNUQnOYM3bQrdC8/h1zY63T9E9w6AJfWebkFWbVCESoXNZAhOaUXl5LQ8AKw
VFiSAhQ8PAKGwYCfSZIN+G2x6xeWPbZfnWUDL5YDALVrNU9dosoMBSzIwfIV/u429dBHAig1ABmT
x9xfJuSL2AVYYDMZk/rZvPxcvgyZQ3hCD4OSVHsBxP5XhBaMpKZmgQJS97TNS5ulKozpZRrTajL9
I2IlrsbNFlyLlzjQ9y3XQJqV77O3iy3VjFGqgA7Mbes/+QhzIXMsWNnLBhXaFa7kNtuMbR45QYCT
WYTLCvUV+zS7CrBrSOzOii+Y8WTdpDkydSYUYHTpJbIwtnwGV9bHK5n2fym6oXD7tlKFBCo3WGjx
4dq+MfRmkUbkdvkNfkP1iNlZvAYsIfWXZgUFQ5AxsNFftgsXX9ZVtHyxhDAmUppuzIJ1pLSweqFE
6lATqbIpwbrAoXUIEVWxuA20TxxU8aJ/lrb8Wm97g/+FS8cQpOyhSUTIF+4zsKeu2FK2FFZXgA2o
dKFp7mQUR2gVHqohCFK4/MO38i55ordtKsozadjwxw4zQ+/HkhSP6PLnJ4dTUf5XuBiPC/W38Udq
9yRAkBwXgMOHCtsVJBThZB4LJpmxeMtmx+A7vAR2SCoHCBk+Gl1vFKAG8ChPIq6i8zDLO0+1LgW2
9Pvy2WxkYtWS3JaWX//JMmDhCrXcpmxUrDn3Rbjeufvwc2rWUYXWGjomrRfunsKt/n1nTtxZzCb+
TkoG5sWcxAzynZWu5zjaleGRGAFKjxM+zK3vbl5K3pFi+GTUG3BO4yy8VLlol9IlMCACEGmuUtIR
GWQx3Nq/zxwwJJAsshAJIZNTYFqbhUgpJGwH/q4/Xm3uBJemxvTP/6jONvDTxLmsOpenW8e80PPo
ZmvT4RxI5mTlwjWMCVq94LX0UNFCxCmhnxxPRg1jkVrLRlYPBTKGg6/Nhoc3SE6aoS5x+mm53DwH
wT6792wfV/O/3FzsTRI9zGdc/V6YBtPJgLFMXIYrbDFAxazXMp0PRlf999b2W1+1E74QQ6X70oQI
RI4/CgySXHSDRS5tFutIMiDVmoVZ2eOwlOIsQ1rIm6biQzSRtwClu2W//YWFTZZClhJysR9JaKN7
QzV4Cm1Qj5GQ16PlG3HhMK7dW13Kf93o0jZybWKs3LGmxkYlxbnFGgGf2eqiAinD5eRUSxTzCuhA
xLatDF3qaWni45KBGHNI3tjyU4d+QYcOl+KWg6fn95J3irJblXALbi+/CRuozx6DcBv/kiC7IxEI
cQrLTfK7en0IQKVMzqFnq/hLL91EpelNoVfit+XnqNC2uM4+jumNt4YVwCWshBFPIcHzgaf/B/Px
xFHiIXenSCPe1mlVQLqW6YcsIAScbczRz4ovt0TuiaRHRIWBfLx0xxC1OLtT7KerjHcMSSzrQFmZ
TLn0nRyvDe4YJpFW6jkuy67ceBvg9Bt5b3r3GjyaXdmxA46i13s0ynR5BNNEyfBNSkv8tTRLu3Xg
UHUuQwIx+Ks4WEmS1J/W8MFy7mzckjr6PY9VmxSKy17y682+gIMXkZtCtUZ+5HPm2sBbeE9L2QQ0
j4A20rkp+ES2UDeDTM5rnYTBZIe3XRVtTqUXbViv35v1wGW7TBWQJ6h26ks/YaAARL8muV8kOB3h
pJSXyi+L6kX3naxrEejnbSgY9a31EumJBLMPYfsuJ53ub4HZMGW+hfonqtn2JulNnluOBfW3WpGP
xVd174elIwD8Q4MVPjiee3xOiS7AGN48egq/yW7sBXeZCSd/fUpDnrG9m2ejpdexNSsynEWqghFn
KyxmByvyBhA4DQX/AtOJXG8DFNZcG3mpcFLt24Rfq8jZ7SpJRahsQK32SFp11Y+idrQPLPDEEH+y
wkSPLNZtffmZULlYqNaznY0EPXBdrr0N2GJsvfDkw1PeuR3uV4bavoHWdzyeoJY16uxbrr2VMi10
BhbJm9O0ijTeoeENKTxAEI13yTjiJlxi8ChOC8Tk6+52O1VDPlDp5ziW8UM6KpojsNhC8Ks0Pg+p
1RK6BgWVIpCAQ57EWBkUDfVZ7P+f+D0F4doTz8G9ussIRZTSpK9h7NHxy8eaqHgQd6j+h5VtZAJh
sfkvO9iV281eKrz5k8QIvbDtAiQ9zAPTf6oy2Old9zZ+uRFl9RX/l0macodfZF6yHuJ8pfhrPwom
jEIlMdec9B3Igjkr7FiUiNTXsalA2qE1u5Orw9DB0+5e/WVgN62c/GCGNtiicMJtcXWFcLTo4Ca6
GZ2SO0MWIHU6my4mIJuhllvDmBCDPGkDzzWAEWYtWjuPIzrabqVCO6pctqQIJ7vfcoyyZ+m++UZd
/cdIHr+Cgg/2gye+0ApviLJ18MONL6fiUFcXFVyp6vJ6dWW5cFTEu+kD43l7GdJQyEDfTR4qWa/Y
OzYhcuA3+t7RTHgTsCWklRE2c5X+TKiXihkrJA6FQhAASF8VWJDGKMbNJTb0fnV7blKi/uwRu7tB
JDPZ5NMeZNn7MBpZQX83KK3NBc4S5Z80cLStWggu0Jo88RQNczphIMe9szH9SyzJIqiEHuisiStU
RUJyC2sgW3Lw50PxW40MlvTHP4EOySVecBk2wt8zmCZhWLIX/9giT2UyOF7PdX8noUMGWSLjPKJZ
QA+kBMwuw2SF7WGD24yUweqZBCncBzH8rnZC6drCzG3EIiRYkdMuWbYRJt67FF1M8jr/N6Jk+oN2
dXv/S/i337YhVPO61TpIKVEid0ZsoCkbQT5XDX1++FrDbhrNl/a9Q/PEnlmoglvyU7V4+pNbcCQm
xuZprbZyMgGdOStb0AI1g8N1iESLpNOs/zQsQUq+C7zvrIXZx9ujNoERoZg3aEdgby9WhRW2vWXQ
ikw6PSmZzFPrC853/FHaJ+BE8S+8g4vVFYkx+PECKRehQlhbWGPbxXiLLYaY3HaHNccBfcXu+Rqy
cRd2qb3h0+EoTL1T0QUPZs6FbNi11wk6XKvhX/pOKxXlgGlHP2C38bDGCvCNdRWPiA3iFebdqkF/
tEOl3VlOnLSz7H5WzID8m1C9BN9+GH1Yr3TrrbRWhqQs5uV+N6yyZgmn6JCDZ5ljXy+bDrcRCyUC
VAk+Q/JqeoR/imZLgufGGIiacjDfZEr/ZhKU8tgFBcCo2hu2vbsSgoDwRjhXfK0DbTyhSG42RuaX
LjXeMDQfZj4UEzjZUIR3pYjaPdP+Wua+bLG1FuiPdBbmfeixLG3baADlxHdtmNrfzsu5FphDxi6s
2vaf22jjKMjJFbk0+zZeQLaIdp+A90bVW2asJ3XSY8ZT9RmM6vis+GMKu/uQJ/g+lyE+I2S8O8el
ETn3DnVY0TnwUoxgwfOQNu8WQ4hWNyZOnYzb5tJWU6p1Ss31RwiKYyMxgE6bNw/pxeteY5v5CeUl
VjtFOZtON3Jv344D+7xElZZaGeqWuBMCjXHVt9AJK2DY0iHyDMg8ZaorgkaEsCncQhwI5ePcC+8/
M5Y5BBq875jM0yma0MbYuupSoPR42eLCyTMbXYfoZ9id/aL7KlPPX76wLZJzSM/pbHHfGAFcX7Z1
9TVw3iYf1/waKZsxNIf+bseVk7dO8jmSa46qqaAA84bXM4FmNeEVVVYr6Fl8dLI/uE3gF1HgOECA
Wrf71QMjLAzCHJCmMhzAQigft4pMukOR60H8gUsltUqSfWfkLlAT6b0WHgyV+47Rv+7l62+zeE9C
aVPolEo2NZju8/uT75IVcXbcrukgk4rdsJZkQU5lWloZtCaQe0GVBlCYpJofxp5tW+arryq+y1ki
acc5hAJUt7H2slsYuwHPVaVoZbH12Cu4akm5teqIUUN70hKQWDDS9kjFfcPmKpPO6kaBuHzcduAT
oYOIPENmA9H6RLlGAferUkSt3DYeGC9HUike3yLnYgCzdR/9wIFlG8HFupU9P7deTx1KrgI83vwz
lG+528jRd2akU+iI/sE5OYhOD/REs9TcjL25GYo7kD67nlmOD0jItzO1QZFCHE0RYw7wBor66fo2
98Yu6Ugom7gLqEG/DdQMX1uMhSTMCN8iFKkZzzILp1jnej+ZP88E/oPFr2drTTDSWmOHi7EZhUUm
PLsGpMLQ53iUJH/sR7w9Fqrvll8ykzphMzLp9gOWaQQUB6Ht3MwaxFa6YdFIIeHNFYBYOVoKITKx
y8psXtaeXKvzJbutH9QoI0SN+UEmjgSAfx1mSS2doiTY2hzKaN1liFMhx12S7g+fuTVmqVKRrAHJ
VH6LL6qZ7m4F41TXhNTQf55Ij2mGBuUBdX2JEfpLm+waklSeAEqbMa9SfGokPYDUoR7Y2PU0uvP0
WaXcNiFJJy1GBRWiLkAZyiYTgX10JhPT96MR+MCe2b17UTe4PfQ9p2kaodo+KKrRitv83lKs4lU+
172JvlLXq995u+SObeKBal43uedDaLl8hpJkKZKdzmEeEax3GIHvpNdCBQTWtN9RgLo1n+7rr1+C
VfSTMVoAWxTis0tZfcIw4jgnjowJU1TPePfLYl88db/Tta/0nf0j1t/RjmKyOyVF9euXziv7CwCy
asCsYoT1NUrmufY6/jDfWKTlg+aVQ/4MIeZPqnIa1HTNcKJd507eFte0H12LooE4S4SGdRAIKwQR
guofpHTdT1HXXN7zPWLZQUMgvwCFgkgka00Op9A+luF3Rw3d6DFUi3KrPA9+ilebRDcF2ANg9xRp
JlXxckzX2/yV17JvpYxW+KW2okKttQva7unwzulSABtpIBU3CRLZkIg+lmib8TRAD6CYI60xva6l
5Qqu+TdC5aUeFqcAAx3t0BQRKPKspgWXGerOe6AKr+Jm/BbSKQrL7IS9vuweMH5pbAImdizIVtfZ
HRSlXWUEFg3IX/DcDRLxLNnlONI0hJKXbu11jZVSqYlb1P2AhCS5NiYwA6/EAWmf9gSVrpFjwJj1
HoMqW4/bCjLaqG8TVB/KKoE4IpIFgbPgAI9y2n3BJ/lpq9BkdwrSYl/yWynPDAW3gE9/xiyeiXET
UfNt41yq/sOBcOiY8qk3HUbCFs/BMnvIkKVm9Z0TNf7av7lqlHO8N1ZNbIXZ6HtoVgVeuGIbftwz
6GTZvrcbOu8kgMCUUephVyBFuaPvWmqRcJlhw3tn+ZRp7TARIHj7ly2+/YDCOQTOHLZfwQ/2r6sU
Jaa608WZaPUuz7dWhzvi9bE7YKH3aLyU/MJkPpbU1dXY7zzqMAxpI3jfKCzBq9xdyq1DCa2HiJ6V
Vjh2T2khDq9zr6801N0b4mQOJUagkjsqoJvL6m5Ag9RRSYhxv0KKKrHBnrZ7EeCpQVNi9x19oUgf
a44AqFG5ZSr7c4HSlk3aFVQP/RYww1q3V8xNH1RVx9Sp3LcKVGuNiu1DM0iQJwhrRgGhK+AIeqJi
k47ihCf99x0LVSxE1FA8z/Z59IM1vI7kAmLEQ4UWrEgv89LF/njmHzGs5MiihI7J1srOPEQ+t2f8
KWe6BUE4W+Y6dr9PiIOO05Theh8DfaaOwLVD5xGUE2WKdu2+XJfVUja8+vg9VB6H1rQ1Oz1A2/jE
WGfc9i4uelvezvnRst37EQ9VxFL08eqm9IKHY0VCC8LN4uH389aepiYED+daeILs6CVn84XNwT++
R/Jps88uxXBGRGpV5DGRHngyITqiDWEwwm5jd1rUz05iGIRPwc8Vtuo+JlgdPYqiLw1x8ZTvohUw
wWXWTlGCdnpf7vytOuvF3Ul/ohHnZqBqhiaUs/8NlOFOoca1/VpuH0mj3vI5yxWLcfGnJemTYXlx
aduIBYztJF+e9i5doM4E4U926nwILMIxQisdV6AYpnx54JRjRMvF2BpXjRBYDdmd7yT8VZi2p9yj
ZfUbxOJqvIJUIbrwD52ukjglFQSZ97Irm3AqcH8uN8DErstswWYGQhlU/Aq7p1pgrmMTS1auz/Su
9kxmD2I3KA/t0FVdGCItbZAaTeS+XXt2JiB3UUG0+u4OaDh8tb24TSWNpI8tSl0s/QgtHM2fKVOb
yXGG5eNubAhpijQRO4HCltICJZ/AYjjW2WGKWiYYR4A1fwvmmZtqErpMwcyfhZ31dyGlKg2goYxg
UcOQoju7C8jTldDJc2f5gKwGWbKscIIkTaPCuKsw0JTm3v28JfA/8x8UC7b9TYE/e9hHGCl58mhb
lKoJJzMV+iqOR57jFc0ahPk1EPxkcuiZ5rnj2P2r+47kyM5FfxxZAG7mY3fgGOIWvhOmP8/Cfvji
HS04XqjemiWxFCFaYQRUNI+dCqnqKYCzGwiorTmUvPUFDn/8LIV1VuxHxYQmkuXMqMai93oGpZa9
fYECDTbp9/ouHsisi0JhmoQUv+W0tbYBhpkprTQ91mic26x/feS5hJ8JAiX2HZl8Sixe6wxz9CXS
XoxzTznywCglqFn+c9zK2ZLzvnISZSwPXntfr3iSha3ldi2WAZauPFbZ1UbIOn8bDzIDovAbtjuV
JcanLjdslp2Xc46h3OY3xhKk2/ONLk9YnF99snSvs9+A0Ayz7JxZXt3u8GIdgmL9uxfFAIkuMmpt
hfQEh3I6ksygvUbq7lljgpFAZQ5BIJkil9kSChN0GeuK5NHvi+9PRSUyvvRhSK4aQfsUZM6hZKgU
n+MIyAsUJ7UzhhO6Y+5pW5A/GlbANEE6WlPsqLCXSwdWUlHRXIMTSthv+UlqndZZ6cep6Hp7EisY
pXUY80UYud1cLH6aeAGUyWnBCwOQwV2/LxFLN0IcNlZZEXGTeXaf1ySoYatljBvEMK/gTeGEAFoE
ls9Nvd9zGgh0D+wEcLKt7YgFm8ZHZgm7+xz0cUom08I4ObozZRKWwp1+NbcTDrA9tZFO23etJnDi
xgPlmXJhvw91EGLP0FXBpdxKAxKdqY+eOGrGs4+aX1LyEXPeWlYEYkiG2xdwkeTAh64cplQazYDi
fPfbzkKkF+WHvprpQkqI/1e1Mhu6uLz44kyV8tDmuTAPWYu6Dnk6kfV5jb520y19jGtDobl8ro1r
GOjxsM3Plx2Vy+dcwkcJh1F6fErGkcgOum8/ph2/z30kp6YXW/8bfu02BRNAMK3sE20KPh0K9jjU
jLvS6E5MJGejnOd7KJeaazliOJ+Z3mC9GmFTCm1y1ogp2C/Q35+U+4saEKK0IhX+as98LUea6VqU
3EclTfwvugPet2T77tsvmcPMpPn4TXLX+Mt4BPD1tqNr3Yw36lU/sfz5P3UCt547GplNIq/JQoVc
XMyfKluMES6tWQOcxe9c595eidOSJgybYn9hzZAuWApw44y+dRvL2g2yhU1he9IqJkyfabxUtHgF
ZG6jzza29IwWh95W7LM1JcIPQI19CfcVsIlupFzHdSy7Vtk9SQMTIUDxhh7A8Nk6ba0TEUf8RdVi
9obpobVBiMT//85gYkL6Nm1UwV8GojG+MTS1bS+JqK1Wy3yx4cMW7seMW5/uqPHfYxMGu2qLzHZX
MsB6CqJL0v7j6XIE55sW/rQozCq5CxojxERiQ0mWsb9MH4/j3rHHT4MiQ0JA8kMVfq+NIYWYZbNy
cGhJz0D8Lr2HAMbI/sf4oPtwc1rq5FYHlwEiBkQL7Gy4BGGAMS0QRUd/oafAYWlrUgnAfgVeAhO6
4sxbJ79xuZEnZegBMG9WO8NTuIMts0EkmNmVMFVqs8zoe6CM0sy7K+d/riC/QJhRnoteT+lFOUI0
hDhz+Wll+kJPQsF/WZgSvuF3RZkqYQI80vOxLzWn9gsphb/1cahqCRIMwgFoNc3wnISFMgLSPt6O
4L3fcRFtRSGAmpHoEnqs1uHK1fp+4+mU2LEZ3mt8PxX2LM2TV8Cid9LIZFGM66CoCO/lc7uow4jm
6PrM0Fp5nODAW/uPSrOwCA+bJLGG0bOpay2O4w/Kms0uCgpOOYEb/9zk+YrZ/rsbYqjczafYCX0U
a53PrcScqr6VGN3qEDp/hLCpvJXf3cP/ucaOqMMxOwQ6wiO5zgWJ+5vDbfQZYc5apSLq8/oZVMmd
C652xVWjEke7vXE6GS+c719nCasUy0f4EChkgS470+g1tRpyaol8Mlketu+7hUKnMUEz6ZGmZTq5
KSRqeNIOy0NWu0WhfwKW+D2KvwF9EqJUNausgyq49h5FP+fT0ivGd4vbnrHBsrAIojL4xd4KEIgQ
EEvuUv1mckkDW4C6/wjPs9UZXh3oNU9m6j4X+bPbZyIwBd5wbExSxaG3vtYxnSIjHxvT7M4FvNmQ
CmY3wmiaNW3peMLo0duQ35YelHEOABMfH08LLNPlDnKrtH7Szhb7199OsE34TPX+xTzshs34HAH/
idDNqz37cClbWv7ZFVGDl6wCOWHdNS1qxq9hjyvyP7PuiXrdAaUIyorDxdiXWHDQddmyBJyjsAOr
tqUj7lu8G8RL/tBvG88KUpsyXMjGIqZVXvByPHssp0T4E2xYzaMgYmaFg4L0ImiQnwynwfpRAv7i
VJeXpUscrfV8PXS05iC0mX5BjbfA0oLgAbuMOCQEefNj0PaMnnlF9TEMIFmHUc6SXhlMpIzHAMUh
3t9VZwersgRhI7FRCSSS8hhIa8MhtiJMDBdx5IF5CxXe08oTxegdBLbokbquJjG3MLvKe3ZUDoyN
4nYpZ+sSGRbYX4pw1LJUTwbeufOzKC88pmcWdBwUNsuJsMrR09+zN1iE+biOLz7yHB0QeMLoiNIO
Pxfoh5jvoa90lgUXRBeAmJyzpH2xqlJjWtVaNRI1TbMfioNV2AGpznfq+A2Am4MOv3ClzlJWlNR2
JaF+1CrVp6vdVxAnbEaRz+Vl0RrHBJyofeGMw4fU2//LkipGSn1IjCnV2cj3ehAxHviE9L38EQzr
O54LqFKiXgn0MsPJ0MNup9/vyfm68z4NWuFGoYc8cOxv37kYfcUKZmxmWDV1UuL+CG5JI5X3qvHY
aUfosdF1MD8cc97dm45i3d+NGd6hTo5aPbEl8Na2D8YY9pNCHLjllv7QCgapyMNfVFCtIHMzxtdK
z7UXBB4CNMm3lzAJ4qZAXIdA2GLkS+fU8rDbjefNamjp1BYsYpIc7QERLrvaa9OgC0dn5xmtOx5p
uYj0w2/1jhrm6VJzxBhRzTSp2TCMpSNHtsT9f0PqB6v7mmkImlyP6IQILfJI4F+/xWoYpKYBmFjk
1TioOMfaQgg2sE8ttspGs/gtu5rjtSt/zX5hmJSFx/f0+YZt3TQ5c4ZxCfbhXQCuwwaT+K5vQkD6
V01CLdKVsWh+iz629ixORIJkZzvy31K9p4T2L2m0cISAV2GDCrkT8TPnhDoHstvc+zLMLavOs2xy
kT3Nu3o6Y7Dz4yv1+Y+jdJl3rEkN8lDr3aE1PBDCfEfPmReKRRLy3mNj1yfBApjqkDVoou0YAhg7
Pxc/2JJp25mHsMsT8HGy7R/DAayR9DsJOR5iycrIlbFVB8jgRKEHLY1lU+bwIqKryE6VTkcWc62m
v8udtI+frhBMBDADFGz8asIb99AFwW5Di5f1VKzgVwiXfzppI1HHR+qv5G3C6Tz4NQYUNq7Hi07X
FPCLw7+9nupDXQwWNM/Th3dn38tC4USicSfZ64UZVz9e3ZDSK1Y+yRWXnOoHmbc8kva0q1/CsUtF
XDdUdE86YaPVS+8O4qsolV7mm86lE6mZW4KIPzRW+SL0bdaR3Twz+AzjmiPp2c5WPx5gJJIBZLlF
Bgb5akyRrcNONBn9Hzob2WMnOktW5TWKP2p3Qf0D24F0OWDaAOX2AJ76tdrQ36M2gVyTCAd1C+Fg
nV4tcTdD8tU0s0am0unQXAsAeGmzsK5eWsfZjwlwiQOsXPPgVlplXA7uY8AP6g0n1k55I4sNO+AM
36GmF88BEWJybVNGe3ZrM3fdnxLejqBBa2N84GNrxfakMcayXrLxy6KgPhXeMUMsR9oBdPWX8PLV
zf/LeWNKdIu8QK8Ncy+VqHA34Y3kTUepqYbCLC/9PIj9j5Y4yOrN8U1qaU8kQ1PzUrQE6XQtz06P
wyXnBLmTUWS4Z1pU657JC1uO4HQvuE8Ecn4YQDUbCNqbgCUGNxhZSxo/ALMMX5rJQyi7PuHW1PGg
B9yqE03J+awV5QPQ/gpurBZQ6dJSJXXSrViiHHMbKg/JrPiM0EC+gNAB2sW8BgEPQBx2A/1b0JoE
gWL3SYWrsXrZiblsVHTEW0lMdCPhC9j2ep10Puw0NU7WP49EAOm7dABLNFQ4wMcSgD6v/1mChQj3
kxvXJ+Dsk0vppion0d+cBSJgc5VLZlA3GQCFWq0ZGdomgQbl8kz3nbDXD5uERq+kkalu6de/NbY2
PMPrBv8kbUvjZEc3YZZbaoJCPG0AnP46yQe2Y9ulQ7sOk8FnkF1EIU8nCk10+Al8VjUKMu5SFE/r
TNRLaXKNZWag8DpUHk0q4VYBxQCKDGnG8WfORlo2r+TVOilOYjpm5EWHuhYMWIPjkJtLVR11gNR6
if1aQFUN6RGvtwIH81S3FD9ByHPWB1Iv53BW6W3dkyetiC0YhyfPMpCTJSL274vzyQb7YcUqeaRz
AX1MhtZGbx0s+YYUgM4F2tDieHkOjhrbSkIMslP6Caps4ATrKW0n+evKUWIiuMFCcIe3CcHIZe2p
FZBUN6e5UxwFO07uN3cWeb2P/7lbnIsudYp05U62TgfG9id9VRkLWMYr3h1c84VRtmCBCjKEkQH+
RdyOpBvtCB9Mw8bjyWbdJejKAL2jP5Be8MYfAzj2ruzBv/k7LFbrVXWTbGDnHbyE5sWFzZSid2g4
d2uFRCgmu5EsaL+gE/SG7xxUPsSkec7GK2nS7Q7TF5mKEJidADPtysF8ilL7BSJbWlUUVYf0rmT5
up5OYYUW7gNSoqNCtbimE560MGtIteojGF3peFjjdgADHaUEleAPBeCZIjHpcv1XODsdKXmOJRUb
DKZANI3ZR5E0EWsdpeL8HKRPLeZoONS2ByIfxcZ1MyHWnv0aasJQham+3FwXIfX/X40SaQcxoHuc
wF0O2KsR/YFXZOHL/WcH2Czt0YZ3Cy//BdipDRz6KYZnrfqe2txPDntYYf9xeirPdIOB/y/1I1nh
V7Aq5NPcAXfG3Mc7wjSdUFE3bw9sYdmF/TBmPOO9s0yZjSPK7PseezL3tCHPklJ1mkKWZr4PLCcH
KvvrnhxpOeWIwUUAFsCTxgz+TmkvzAF/6HvLTb5ZVhConnog+NpeW+UlN8G8DtZo7pxQu21zRyIu
k5PoDRwfvxul5imk6NpMSxyXMcG063eCQ32spLxRaKfUCzX1PqUpi5zu/6NMuD0EAMbao22b1/+A
n0EfgkoxDj+f1a3LzliJ1Y5Ko0v7e97OdBP4kHnBfDnh1G5TRvgBRzrPYflQ0tuLZRTuVDkU3mDd
0aJleDZA6Vvv60ov+9feknbPtVMdKfSB4QKAhFL7TFtKn+bP8iOIM7ZQhMymIUVAvyYieMXU+fep
1ilG5AHovg7dW9QSFpMDcUJt9uOralJw9wliFi05JiFGHb93cke4f8oScmUzas/xJz3Dwf0gpnWo
O53srnkXWG4/Z1qIz6hLujndkEuRAIxO+DK0v76tTdh6IDm5JwHvHOmjE4NHZZaL4fi+TkraKiJt
zJnUXioSqElRIuFDDq57lt6XI1t798aSCd6q6J/zCRrzAHu6Od+0Fesis0s48EflEIngYLJ4pMxt
gIWx4/MmDJm+xwaCXiVK6OaQp7eieuLPZ7x56UD/LyYvKKJgSoD2/asIsfolLpYeR2sHeJaiGEn7
Fr2VTfdc5Dh4sZCnjxsAYuI0XKdQiuA7G9iUFGr6clBa35AYFTZx8DbtlE/QmH2Y2i4MNUeDcfIq
ZvT4U5yUuw5L4ckZ3DzHALYyLm5CWXPCJs2+hhYYHPvQ1pJwRxTI2oxczlK7s2Dvh5ohr6LdLDlw
wNPykzlgc2B7UwsBnJEwUYcY4XV9K7NfE4LcacVbBFssuYsSVY2iSLlh+DEj1fmmc6279RsvobJg
jS0yXrrvY1z38Zv5Xk+Q/KPvRkip7rT337vQMFyWJ7pnsH57FTYzTHXOolKBS9PqFlm2nKxpmPrF
Go2eHIpTmyXnrD03qgcKzbjQjHDQgHyVgjICZZeUxkoN3qHhbCb4VPl5EL4ouqeAGNP/bFOfCNxT
Zpb/VWHh7L0c4WXPEtiio9OFHlwarACAoxJYIZdeYuKPTQHvdjbmUh9rqxoUTq/vBRTmmuhTPAVL
lB8XFJgsP0cXyqiC3oz7nZoHYrYQ5P4i9OKok8WEt4OMTi7bN35meBASJxCwQsnRM9ItfIzCFSz9
AZfA3V4hLPpZwqpOGtyx359eKGfN+yVMjZqlgCtAUGCjZRoUpqzVS6WtpnYf0FvTpnFECbx5j+lp
NoLOwjaHy/9GMl77O+pqnltjXWHppeKD2UuYD+VIa5psuXPrb2r/nnvMJEPqwIyLYEi78woW/Vgq
FbPnapNdsDhMC3KAnrr2AkLDIBkjrJrYNlaJwwkVmejYrUNWb5rZrijumWpYpf7Aw8YBU1FG82df
EPCcmq2Gbxh3/v6ZqIpnBoITG3yiBSa0uwP84ZJjOAWOOuTyVge+eioHe7E8WTEqo0qtndghzA4r
vKOgeftO32nVPzLn2DOC9g+HUZObkQdJ1XcXIWTwFyWMF8hPFNzn2+OcaqJGiTIHPUOG9n5ftOye
7cE57lfSQi1G9wVOGIgilFdtVL5PHJJy808/88w7Zx7qErdv9q8eT0t6n45OYLZ891Zao+QiM+fX
G9Hq9dPRwzwRjNJYNbB4U0VziAR+UaAW7a6i0g9B9tVR8Z6a6GFZUxhf7CExhsPtRK+CGYA1CKL0
MBJFjnoII/9e9pDhhT2zHpK83Dujul9oO9/H8DAfSIvljySxRtRUwcfLeTmaw7FsQl3PjGKRsNfw
K8gRy06dofYU8GBTN5F11yydDi2iHUZLP+RJTdCJstsyDPffT7ALaeliZIlJhw0Va/3qGKZR97Yp
ie8bkmt477xA+hOeddz+rxkdzNQ6WvHD7tysvhPRfF/nX84mANeSFYasELTszH4AmiesU9fQ0xDb
frto7fylQa2gHCV6/nuSVwlmnnTpYufcs/HubYD2zsECY5dkzwNBeNRMcYEkv1WVXj+Xtwf7NbgN
GHYDUtYx2idlRs41I7qvaCyjjc2NW5TgAbFuoXUgDkkQyg1GBfK//6x0WtCR94LaCbuQoBElBmKI
+zNlFtP36rbMXGGxhBHoenTaT2A1m54svVFVj8AYzRzt8h0mV+Sbvi3Uypb5WUofFwkhI2nak928
grhvZNeKpdVFCln4FUlVoXMdrHbncfveh0PYTRHQ7v/lUzYtNBDzv1S0ue6Ggv91HkscRERUh1hn
HQEfGGkdndXAp8rZe6JchzSPNP0NqYJ4YzOePnurnwZ2c5hCuKCX7R/YttpRoSot06SHyP7mr+sK
5EfcNQIhVgNTnV+QxSuKWLyqXun2HFyvk/OEDOqCk7WW0VUkcg8tG2pQ6DpeP4VaH9QsVHy5qJXd
cY3t/gi/Go3UjD2xb4d9gykkGQ/ZR/DZlcMU+qeTy908EBQeG863X6mKOrthMRQwk+LVbp/x5LoW
egrYXif856O8EkEYfvjezVr01SWiP7EabT2Q0zCWzgyP2cgCuIRBnhVHcl9ynSbqI8HctF5sHdCi
sCe0jwELZYNHrT6gElWAcEWMkA8g0G9IwKIbhF4e/ww2jPJYN9a3AQ2LKWxIoZg/rCQ75bZ+v8/j
UvBrqHy3yyP8M740ojVe4V1MbmEJ+jJ9WHpeHbmoopoCiXLjpbdaKjEBo8oXsuuV1lUvjn5bk7rC
zDUv7pUb8TyOcX3l3rwquXefWIwpAV5DdUdNCGU4Nq/TIxNHOXEQH0ny3UPKqE0otGYMyxDC/c90
XCvsCncRwrg2LcrApbotR9dHvBlG2rh0llKNBFODwhlOAj12xFH+AGyLg09cadRmOWDnbZKUovOT
SqSVQYH4YIOtMqkW8ERoCAfMm6aJqIzqhU9ZIXqX7wnqrwPv3vV/JmbzsDIlrDvFXLTsiLhW5dbR
QqlhVV7w1LbMPOCBBYTSQU5zbFEDJ8kIe+eM5/wUWV8J0JjbZ6RrUye7R5WSTCeRrXT66+q7C2o5
3TwYRG2Q8rwKvAgQAMj8cRIVwUn3JdgYl9oN63wRO1ie7IIcd1Sw1PAV8jTBEWcG0AjiIemAUUtZ
JcszsE2xt8I/cpUN41Qu1jWEF22tGJYbgWwof2HmZ/m0bIKwY14Lbxth/Cyazrh4c9/ZLElhiVmj
PJQyv8pPWqBNaom2KhWK6GaaCDBm/f8imhAUNvMHrRJ4kjFtZTBS5ikP6jsygfDSKKvkLueLn/Qg
6bTfObikUmCQa9ap8QFM3bALivmWP5h/vtweR2HhW86xom1Sovyg3cThxQh87cFGwJ9wgvpDXeTm
suWz2GhSGbRznRo5yVPWKKD3h3xGS7KHJZE1OvJqI7lij6H2eANSxYQ+Ao765vGTjMtoxI01Fg5C
ESNwOIFK0iGQ6ruHQtc+ju8CotYnoVg3RyUKfE9WdjTzU1AAbj7GZR6scItQ6/7BZ22qL1fXX7fB
pnFcxO573Ggu58Cos6Dq6ZPxcSzbdUdX+GNS2lXbhgAXjPgaJBQhBihijr57lwFaJPHsQaQE/Ycx
HGdx10HrKaBJmm4PC4nSD0AqOJFKp4GmSB1w4xssagCTZitoYbXeorrbe3SsI9zfRnPvHKS17mrC
p94dq7D7Y3j174Z75FRwBLPwjZKCPUhq0dlsOc5+uMXUJlO1fUEvb1Z2aBWxtR+2UDy7KP15NOok
seHfCRA9r53hubZwZM6/bsFEb4UpM6Z9DZtk01aXGvAsS1Bjmm4c8CRY77tG5WQn3EZ3EAdcLic7
MmHAXa0tvZST79USrBfizuQrF1tjxP57fMR+ODovvf/SEsSq2frxYD5SPNCV5PYzXyM7f/CRVD4K
HhpEbqmUanGa43sjR24EnFK9K72V3H/1GS21E2BHO5eGAbMZFjwTHM3+9ADz7axS720eMscSsWxu
JjmsrH2pij71fnd5EdpgqZ1snl7eLiG52I02GtTVvDCQpek7FbBtFzh6kKjA3oTi8NQtTBTgDEiZ
yMmOYLd3fdxayfqDsenJADoiXqyzf/4XRWlm3OxAZVEn9bNiMAoK9+LVgih5gvsNcofMgNSj8KxF
YihIrxKiC5ZFehKkv1kvfQpus41TsYqXKnqof+UYUPnOqUp5a7X7N7ogNGsoIveG92wK2Rwxn31S
5TTPllIquNWvcAwHsaAiR1aHqQjp/dpg7rCPtPGkrPP9+pPPVKHs7nZjC+WLauRqDe8njA9JyRR4
aBw0jxwaXbhiyb6iEg95h0W0d2YPslxx8PZszvr8jsvxBMqzDhC/X2E/p0t7vtmNxWhCRXyLPfc6
7iQVXq78VoqLJoK9xA4jbrcPa+IoYG2ReeTmSC0cITa07qcO/uffaif+SMoCDUqqywRvlLKB7jIn
CU1VcleROomU6K2KwIk4phevTGXud3T+ZMuUsc2Nbf81Bk5yK1Z1DAYVuEenWeVWrDexnuVBdVL7
ExQ+QICfjcz366Ep90q/8twGph7EJnq8GN9Xs3ouFyCveI0sNjnaf5TCohZhgKVpvE9PHqwL/3xl
zLMrodIccsbVkkiuRDxhfkvPvHacqOFiiY/KY+Z+9x81k082ML1IZ5vd4i8jP2dgzZTcXGoGA3jK
d4SBvkdU/58DSf5RqT8sW6SGzaMmey8rPBNaJfS/K2ULncudh8Sbeu0JjIV8G5njbIDq+VVwKqau
XfW4M3mk1ggJW2KQKNz4D4l6GSGhg9HgwtBor4LsEmAOzJ+lVS8IV+V00CV2lnZZOO5KjtoOiQLi
G7O1xwMWngj24d+LPsZZ85ysnu9M3Gmc44zBAYOze3YCovrMuksFq7RCJrYIxnkNGSaPSoafdMfW
rjZZvoEZq2jWPpjzREWvHpC05uh/iJjywN489DpNq7fLb/ECJMPvZgg1GpT/sVVpuaGJDKKJ6+mN
G2c+3slBznHbOl1i/UpOJjLTa8MpmD5VFEfqHuLEuEWhaEFuFE922kqTGHcwlxqJhOOIspn4aaf3
BUWgOfUeawh90qkIHwo1xRXTlS1hPOP6f8Ce+SMNkLd4+Shi2UG7cwu2Mv6l2WtY06OCNyw+7s+O
DFliHOYyUZ3PaLVk/3KBqh0Ac5zdI4qkxCJLIvL330uRYFo5j+QvjukHm7Nu0RgPQwr6PfA7m2Pv
jFeHDbql4ZhMFDdpnFSBpYmQpAfWzwbSeaLUo6239tWRcQ8j1FcR22ouKROPIM9v+YnNDdRBht64
Q/L+TqPJKaP+PpBqB7T8u5MLKE+hWqeayd5l2Ay9UJ4x3CYvsLpxDUSLzj3w0VDKtWWF1rSqzLcu
M316X0MOLi4nS1siagZTQu9bkCQEozhdrG0MUyTr+KNzKEXeuRm/SQxmrT8G0p1W8/dh4BLoCXtl
o7O1puaVr1RF2UtaCNvs6w7+n1bL1A4aYPrMTnpN2SxRaV10Dv61r2URS8jzC/Wu6de6D4VtJFIE
xJyOXjzOIyAGd7fQTnnT9K8brXFbdhvrKoKE4ppfqwYRUSWBx+63STxunBxEaPmSjvgFhBkABSEk
7CWAzno6TPnVBW/p3bhvC5EjZdz+dLSPtzBG4AO1mPNhiZVWH+J1SPzJbrqG9JkJuXQofKTI5zD1
I1Q5amkoa+Ku3tH1UlMPCy+THMZV7pYnEc2JNJzBwlG4G8DfzNAfvXAOqxMS6XJveSCupHIeLSv+
gPy3GO9kpfWAIYvhyGinyLxFNvnqQGhIqWIyyMFbIbub2OlWjEi6YrbegQd5WDb/rZurZYSrT8qT
Esuc1X5V6dnCiRoBTJ/bAMHdMafH5PpJXd/LJBQeiSmDsOCmtnwfp2xUGdH8o6OuV02mlRyNs+Ae
CPgLFagbrk7giN96Z2DQ+Va9kylifDR46ppksz+RBR33vnFtaPokCo47UsoRe+IG50G/nj3or31x
lYnMdQTRVNBf7jBe/Ut7wJRNrMTkJGehhbYdOXx19LoTWf60WL2qlpiGpo19k3y/RtKFwpgFw20a
vS9Pkk3oa5J2Z3R737Jf/akTtdQeRmI3+zu0U/T9pqdg2oxEW1EeiBKa3ZzvVIf6mAh+NXCqKNgH
Vb0u20/mTZpIFNTsxgafM1AAfzA/R2WgfxNOeFqRn/mCHyVXaOUKdNu4PoZ/SGakIuv6Ea8JfK6N
ERpIl8MqOmf/U1FwA4vnMZLvAIFpnVR+C17BL+uuPr4kROEl6XDNYaMVg33azIHjqi/OMUrR40t7
ciho3gFUuNp9a33BUgwCtF+kQMOsJQOIz0nkcAUtVcaCXK7JHH8eEPN1BAbagQztGqvdvVWTUwI+
SAa2lv00lxdufS7KaZWOo59bXyAhcI3mUcd2Ze8615ZEIIDU5TtsmCIV6ebpPm2RA6RDEwLGzRYB
uSKZS2DMlbr1jO5DqVgDc3vqyTnuMxhTwzDnA5D++fkGyfBw+eB/zXZDXigItlX+Cs/+PSROKBYE
OOl9ooWP9+IQPqKU8Fj2jqaRYcWSda/fDl7xwC3a8+csB2Cn1M8YkouNiMQofJw/PZKyVzxGsFJu
bfPoN3fnQD7HjzYVBQ5RT4fJHOjSVip3wfNKxe9JGjFLmHGLfsvdC3HesaQPXYaInYVbB4UsHH49
XvEsWbTV2Qx5rHqqqMRs2Q5+Jz8Wn49AQe95oId7RNfbiqsBuD32S3l+uN7TEMl/ph8qEwh2xiU3
4BH6XvbTlKL+Gvnkxxup73fRH1NwcJ72Akch84Hx7ZvldeOPr/9NBCTbwRTUOJuTQmmaZYPoOBnR
BBf/DQqbQvxzPCmMCZU8v4b3c54OfmVfSUw0yFvrWGbnmw8NCK8VJvYf34kPk2beshqrCC05caAp
Mfb+j2xIyucYbG7kNEQGGzX1mf6R0C1YAv+d53tkw5ms8f2mwvdvz2OOlfSyDcl9wIbmHBIuxCs3
Mi1aTmFvXGZW7EvtpYGw87mzL0RBEVC1kIwJz7QEyJy9zQaXZ99r7Ywo8Ycpl4Cxpcp9od3EnQs2
sjLkWjfyxvi8yqJnlb9gEI/6fEsbDTpRQwhK/dQWfGvFVQWaey0fh3jwC8QUAJMcppefj8r4Wtsn
jyUt2lXHPBCqjn0DSygfABC/ZUToK0YIRAfhpbQ5y3e9T9IGzRVjEPeltok3tFbEDfRcjFq7GUXX
5c+FE+qBELbBbw5OQKufpzZrUn1vL+G6L9/K8+qMj5kRtD/8J/+1C4nm7lrz422fSP2RPcAqMcd1
g/bqhbc9hz0dA+we3iF/mwIqTEMZgjKzvm09FuIYqW4LcJfBt1Q0tIVU4DEZ8eiy+WYR1ogUKOs+
uYCqtfjAielXAPjFKsnxg6zOJW4Jd7B/BzJJyrFiI2ST8EyGJ1v6ZkcrF6/j8kE+LiqIyzjpmrsU
5wEWENxv8MPbu3gERXzrEjwOBAXzWS6OwFudN609ChmSTnVJUZNNPyEh8uV508N2u7dFRTxjJbRi
oZTWcvlwUciYuiDvlI11wbepaM4SY0eLnOqkcQrsIPXHwnWsgolXYAJ0jQQTHPq3hKLzUKbA39Jz
Q5lbXL81NvyYbgZcHeeUPpNWjAoPUyjpMZJOX38o9YALkeSWdC05RsRwQpghgPl7FfbaYapC0KPF
dskNKLQX508LN7TtukgC8SAxlOxVgf7vuCG1DcxDCXsWgizXbWPZilXaeMT6U5+I75GeL47IzuBd
AifOlSP4ADvNX4aQ7YKn6H2EWwwP03rC8Ft40ctK10ADd5F83wgYB5ZmrAwKz2stW6gehpoIbu0F
QBC5ihuz2WkOyDwqYThLgDSLUCL+r4zrqpfDp1eqvqpZTKf5nCz0NY5dzTe3w4Z2KRDJAUgBDPvM
/5YmuENPyX4uP8/nOoxcxUyKpJjmlu2JlVwWoNTHkozFD8ThD9XjTvN2RTBkWxV/6K13zm9yJ6Ac
00uDX7JTz3lHW3X4ef2l2tg2bI3i4OM2B2wWDR/JoXZ8Eq8LwBXFlOhJlsn6z1AwmEzYYOC3MVnv
v9oPMZSnOePQJk9nNkGDB3Vz7skHwb86UYxEJhm80jXziqkn60KX1Ia9Ue/FnwpkgexHTUG9EI3O
dUzQ1Lec1zt29tjq/nJsHi9pFh2Pq1aq5FN6KIa9r+w0udcH0CXh4JZ6hwuBrL4bRHZuPQWxkDHD
o0G1YnLw7TPqtVeEk502sON2gwaVuiqBWtAwtnZ6ZZ3ZQ98bdJKcwZeeJWbGTkow8kbVqj1UNDNQ
dWL8+Ckq0eRZ/VlEEhgavVr6sLSBYPM5HSfTUQZQhIfaU+fEyMlduBxS7v69xr+Ckz1J1+tpIzoL
cbgDNpeCuMtgK4VGiR/AltH9pPBYFxlfLHimKEshjFl8sXc8TEI9ftYxJbyUPl92CckxgAMWgeXM
USbNRUkYjv/2Ja7d7uslOqyaDKx0yPnUJrAUZkm3HCa5JoHTdXH7oOc8hmX2nAMcdZsTqdEbG24+
d6OJftGUlUXeM/zyD9PfO/p7BrLBgVTuFdg08QcdUdQCiaGW3xqSJzaElxP9Ghbmt70LQgmnzb/n
XB3ui8wm/UjbLhXle6KiZjSupNOYNoSAShuWFr8O1paxipLEMl4A5EZx9bL2ERHHwIr1HTSynydi
GiEZso+Aia2m/oBDRjvGStAlcfWMTAOCRHTlgc1Ek+CPJUOnzpioHyYz4LVV3E2EB1ZMjTx+2dLe
k9oHQ3mkzfT+Yn5hRO5xgO5KjPPiM2eEKr/K4zpW12d6ZxyRj6NL55YIIjasXe4KV3a7ENti0AXR
iXfJCeqQbJAIsaMKAOOM/JTlsui1AzOdAqeCV18ommIW4/A7NEmT6McDafMDjY+QxohHS8aVQtt2
u68AuhMM+Me5Plct71CwiijKfvBuTcXnGQLJ2cSyhYV+VWFrhOglt7PrZKNkSv2I24VR6W90jDmP
eAjRTCsDcv6bC8NxJa7Q5W+ddKvQm5oZzA0jv22X3PDTNikrvgwN+fsX0uwxRusYBzlwwpBSn3Tk
yMx60n+criD1u5/VVst1vhvKMlKK4b226LT9vJv0hePtjM1nBBzKVCIum5jC+G/HqgS3xknPWtCh
FNj4P2vE37l3mq/NwH7qj06+UM/k23pmUzEtuE9PH3fs8kdkA12Pasf0d2MkcecZ48oiJluW9nWx
16tF10kKVpW6bJyL5ZwzRpS1GyDycCNqPoBpGaomMKkCuAmUh6elD5L2je3CzCEW75KkX8MAy0A7
FFitV8M7CTfL6iLYBTXQ2032pVld+E0eoEn1EqZ3RVYrmJXfctWvJkattzQTfnjFeybNCEQiW6QF
vtc66tU+SVfpLi+kCxWaTTBaba0IUIajWRg5SDRWjIn7yJCQBhUCUxoiJG1QH8LU55/Njmoq8i2q
OD239vzIx+JhXKC0F0l9TKmxtwb395OZxmqHvDbyk6sXKdFQRyA3KZLTDUAXfBvgKVIuLgR8Ra2q
hEIJ96Eb7+45Px0Ea2rhKTXCwdd/XjKike9iDPtpYtHrkn7pM4wDR/6SsaUL0kNXPxjmN6sRc77i
0z7DUOnX3vOwDqD8Xy5vEKW9PRJrpAygIHS5GWUiBnjbNgJZUSKymMqbV6htnDOHxTGroetIoIsd
6VHzAsROKetv/IssbHlxkhntTsy0g/+NYi240yh2jr9fq78+itxod8IkMGzuUbY1i6rB6XS6H2W9
LFv7KEKC0Hd82sKv7LPXSCRwW+nbFcVwJ57f/VWkbcFCNk7bS+tPWhSn2NzfGPhsP4apwYt9qNNS
zxzijgYDfdYYa04s9WkpqTA4hwmyF/T83sthNK+RF9sXsaM9cYXRb71/zanLO3YW3fEJ6GEHUde1
dyazyPkh+9kWJTkeDY/YHRPbtYf60MItWWt7nmlGIS4GKN/eRVKP+Vz1gHu0jnSRF43gQ1EDOywe
rwo8EITDZEVblIwVqK3nX9ho+VXAj4ZPkUmepphBld22rYq74tYuxeikkZU34aEI6DlcjIZnIIvV
wT8tB9oBbgNGJF0J7Zuqn4dtuB+Rf3AlrTsRE3f7FgKSm4DAn/9/cdqKP43w9qznuoffOv+hW/za
aW2kI16ZCQ33VYGo6Y2qFGySoC/EXwCEzuCrgJUuw5bg+yHsUWzglDQf5Q5V4mxLnUaLcYv20ypd
XmTLFASZ6eD466+q6cd9fRuT8aMZdxLRdP0nmJIjxP1l1diAo1syTj+SjxzpDs2c2aAe/MVIdnte
fG5e773olOpYDIYZbKf1UAYQXH6gguHJxXiIbCu4etSf+tYDSfzys2lK9ITb4UxiA4eoHYN0zPSE
o33jHTH372Qly664zQCCT7nVwL9i70BRcb+uyWuKluoQdOi8+55aOSRaOKKnYEyalBCJC/ovILvg
47yGj93K3l0jKFU7zkOW0CFEghR8ZNzckoqTMXz7a2ETMuFMtDYTvZdVDTN6EBmbL0lpWTzqFy1f
2CIa/Lm5Tu5A7SDbNNHiyDY/JFwKwm4s6K4vTiSM42webZKpopoS1UXyfQn3HzVnGKyqL89hfUHh
3G4gCVMf/mVeyNacKU1mQrvKXHhag9qGFPMWBq3NvpVRhh0cjKEQvHHb21pA9TxXkmFB8WrbTKkn
tTRenU+nfgy/q7n6hGppq6L4BJMWBIryEUx9yM3s6l4o+rxYn0tcqZ+ODrh8CA8MRRrRQfv7OR/2
YpHNHj852pF4O7VK8eeuIPTmJQNQ9PlBtxxDPYgZawkaumNC7rQ90Mq3KTf9br9WbvjOu6wtUBbI
alUZOcnp/YHY999dFA/zYBAR+eebfWKHhxjxA+VFTHCQqo/8KUp/phkydSS+0sfgN89p6tLCz3sP
9pHGaf9oT2MxJw68SaB/RX3KpfUGXXs6GviomKbKLkq7JYp1G+qm1vFAHWU282HASrQSOuvURdqq
vjIOjy8cLeLNFPeL7w46FLDW8cmYCaCzkj4HyhcglpBTPY/Y82c23HKB+4oiTxKhKU7ztHWgg+DQ
ajsVQFbO+gLKHAOMs9Fd+SYfkAVbs09dji2ylufGMmG3bVMx3W/6vxF2IZ5F5JmePnWazexkAN+n
2fNB3nqxC2JXhmhqmmafXHWCkj7BlKBtJeOQ4kvUYyVBUb75lqjpQXqapOi0O2VmA0iTF4sI0Qu/
O/4taF3Xmlip+O/zP42lFLQnKgidEaSW0+MTIo2zkb5VarVz9WYhmsRvv32ODSc9o3RMuS+RYEDu
HzKCBSVrIHx0X/1OkN90+3YJrIYtTIOFM0T+LsmO/CF7RxYojU3EjiP2zpImDipII/AQuODHjw6b
N+GMKRX13G+zLZUOk5YeTi6WYmHtyCQNhuh1Ou1m66etjYgeRXNU1HtYeNms8BbgHRCPYMpxxymb
/DGXYGSUQ9bt9i1maqAP6+tC2ZfSjko4peb4HbBWVUQ6oKbFYDXDmUIoJff2bM3uq0ULRpilZvpA
WgAxlMFCfwlAHGlIZPXZbZdWCcndvpASBlv8OG972TIQOqO7/C+tmW5EHxSYk+95tuCOzIJHMY7r
H0lP4hirk0MEIgn6oHWkSOLzXGSDo7H3X/f5rggaOrHLEsjICwaPde/S+UvIju9vl4GwRodLwtOz
Uz1EO754A2PihDVhZLjuPzdYG0i1WG8IxYuscgHH4RRUBlg+TeSlH4PZf94DJsmLoMZB8HvqbVnw
aNJoOzoU2dhP25a5Tm1xPs6/l0MQlaSRTLjGhmdQJtOAyhsNG6xWp3MOxQIO8Gb5rfWqGnsIlx+W
o+HJKjhQ8PE5V/jCxdeOJ55J3vd88rFXJZSACd/DrOcUTukakG0OiDZ/4hg2kNw2x5KqZfcY7A8j
gvnuNOtnEv45gB5FcBi77spDvicTjdNgC32Fxx345RTORLRVsZ6Oo5pwkmb0H3H3q/Mc8gOnnCZb
Znh4doYshfkp3nm3UPaSHbtqbldYK645dWHf7y185j+10x1edxW9qPQQMZ7yDY5rufL149UYR594
3A+Wu1ubgkRRHlF/j+sCn4c5kiO5DWLb/x2rFwCBUCdcoe6RkGwbdOEOlUZiakxKvTi5ArHQypq8
TUEOdpCaw2Zpl9keo7ctcW3PZsX+IUwOxQSHhysOrm/t4Xjb4JoWc7BB/j0DA+2+WsRwcs/ck/cH
ytVlaldxrqkC8wwcrC6GiT2UVb6pge1kAraS42lVMKLiJeG9LBI1VH4d3QWhfVSQXmhyJpvU3ZUx
rm1MkcCPLuvLqkdBY43JUDI305GLq5C/xCo4UQaX4MGI4SG2phpj42sTtePe11WQqLsZ6XLQ/7Qi
IESym3UJ+9+3IXuSgCtWK1QPirYgD7C/MrieQ+Nd9EJpDfsU34yzE2oPhNc5tHZIvPfKNXCnxKMW
JMdestKXUgF2TLlLfokfNKc5LRx84qaD/UKtUqIP9w7hdszHsX/IA3wrth27aLFT4qxxwslgS5lz
bLRMcfBwpEx/+iuksg3YggCA0re6oDTpFWWAniKzIFbMQHnMaOVTO5No2unInWh9TCbtY/e/Uwo3
SO++gKmpb9QJpomBQ5Fl0qzNoQZaLkgjIeXCgI9swwrp8AwQ+2B+PkDzLmcRKZeXPlSaUZBkOXtv
mJuFtmRebDlCHBlaZt38VYXvR1pwr90H40QDjMrBzPQ1YC7YuYbUZj5Gu+fMPurRgcHN8a726BJQ
p5uNtVKhTKIxQOA6EPWjJRTw1LhspZDQ2JEcqsUBNyEogIMLxI+xYVdW0j+rzxualuan4DKtToew
gGsK9NXotxhbfd8S4Pj3/MKvqpJXnUkS993QbxZEbKaHc1Mn1Y1W9dT2DDOvtENtXwskWUWLX1kH
4m+17kF69LQrrYYoT8K8sbkKsQfaNPshFY/2YRfDvCmdHuO4Bll47RJSz3X5NJmVfph4rMr+LuBG
z0uA4eyV8BXLNOwoOhZOvDoC+vfYq6YIBAZOdtHRPLl+aYbxWoUmHsW1QmeD3UIHb/BAC5SCEBEB
NrlJf2Ni+LjzdPGQBhNOxRZqzk1xogjGYlaq1hQy5ba+3dwAxa0c7o3owVSMVhtFsY51R3QnFQuE
/vsdS+yH4kWX8W3ecJpoD24HY0GR2qtuW7mHQXGlTTAFLi1r//7vgWUm1IgDQPUwuAm5HlsC1rYJ
WfKnc81VTP1gcMar5S+Bg3f4FBXEsI1EQMpZUdoy80ghYmf3WBeamTYGcJKQZZ8xJ/w0HpB41Oke
P0tFJ+kAEEzxbhITwxBgkW4OD7hZsLVjMsL3B+8hj3eFAm9DXUx48uxpf4+1CymS+IIuvPryT5Le
4Ty1MdODhhj5I1Xp2hSNJtGSEvDlPf5FZivJTM5CEQNNKgDnmZ0/eAL4+hERY5Bg/pMN2yn1MQOY
GXTeOSyPSamWIcs3vxYavTAZhS5wFLtDAkinAbRODsRItLMf+b1J84bkQgSRjj3vZjt+QkS/tg+9
+PxAjge3n80aQYk8MMkGsoC9g22lDAHXkKH8gI6YNZ+odu/CjNFStbe+gq0TieGcDuekrqBFXfg7
Lmep1qjjnXEEkwt5GlrTGqUR1PQTlk+oW94eB+fa3f2nmzqC+m2xiB2h50H0//9BmiHrobKg1dBz
ktfThiaqmxp7Zve7LRulG9JdA3axmpoRbvz4nPEcvB29S6KfdqYH34UypNdXefpXTBX9Aemmc0It
GI6mS7e13WmH9tUbFQzkxj1Laf7/w5+HAYSZ5MgZHM25LNpJAiH0a+fBhVBetCbG3tPM6nTZyH0E
CsvVb4JTVNs7RypLKJiHrwSmZxtvPCZw5sA9lK8c4YYnT8OC8vPiOFxI9rIKC2ZzMb8ia6a+SkcX
59MBvQgcOCho9Zr+axJpEreTrGwx561RvFjBsGJquNcfox10X/kuHgKHE4dK8wWAT4QY2y70l5T8
8Ed1TwDnpc8YYGR7VSRqIAplNyvAlsT481z6gr4SFKupA/s7Zsd4Ihej2EQ1CPHi+vKiAOP9iqzO
5+leosltzybJwvg7gGSLI4rw242DWB6U0DBEyNaDbJe1aEL8ckZcMMAsm+422eih3QOHRdgGKbHg
zlg5wEeaiOCBXRZ2I9/3lO+f6du+3cxlpqXktV4MuKztvQRo957jnPEhfQSKbsuLA1u06u2cBUxs
uA+/j/O5hsYDXzud4JIxVyAONRBxyY7pVqKrdszLl00PA58iMGIrQZf+LNNdJW/X0zF++rLnGX4M
jdtma0xDpWCfXjt5zROup5bRuvb/lnTy53mRZ/b+0EKD4qbqt0al5vuaKDdlYotSJINDeD8vPX6u
y4HRrmWIsoP7+iykl9iApg0wJp8VIioTCWvYXVReiQrgoDdUqTqbX7IcO18VTDwTYAlD1x5H0iF9
5YdpVNrwVvzP21BsgkdAMEQfISow3Z97AZDixyhN7G54yhzPj1tphjUBprj1iMBFwpSfxxy/H4r0
HibmEdyoJ5hcncPbPHhcGjb2FOEOA6OEC15kTEk+21WzjiWBnSMfGaFkwoXlshtCUqZzHb+FO7y4
YpwVZaw4dbCMoH3R1kEiirRQrhQfJEDgC8c03ODZtkHbZ+0yAIyZGg31CoTi6r90QphqgU2miXwG
44CJz2VSlXI+j1wMQ/biRGGj72HFqRaRSIxMKAKoswHU8QqrQE1UsOTMVHChj9RosyRAXRBwAgdT
wUMEJjZOfQwd21jMdjFEgA0AyAwE4pRlkU/H0Ho6IfEdzn55Zm7LVqkoV2CVOGkOkNf1+f2MgAF0
79Lit/rLqhPSgiqMzjRxw9yn7AsUuvCHm1Y3mQNHeNzFdMTr2m9eAE//jrdcQRY+ssuTV18Qw60e
V5x4XGjf3gVsbgORB/PwMeDAzQ7lWveO/aHHbQuXl+/ny1xCTl+dt13tko0WChvM1o3iCAsPgzKx
enz0MLV33xGO311HTrB0ryL/e3X127HwH6jTn+7DYGOrr9HLHcocwKJfLiqgNzQTbD5Ro66yyYIl
pwfzu+GCbveaS8EarRlWzywyKO1E1BbFQfQ9H9m5ysU1Dov3sTMCKiZBCtdMzJmnGfABLHE1KXkB
Kfh1gVmVM/IuGyE9hNdyRKYYgKIOiyexcVWJ3AJfud2OobWgjxiWiBmS29/hmLA99BGwTyeTdJ2S
8vXD2G9qjncJXnjWZl4hdbbPFnv+C7rHtjgS1/B4K/SQ5ZhUKvbn7wv74SGyoz76dxsk7jFU30HG
wbiwQJsunYn8ppLHxp/GsTCe4KNuI+0/sbWwpxLRi4AVF5Vrl1x0r5SnYEiboPRr8UFj53dQCGWg
Eu1Zq6ks7GsNZIvkM+qpV3PJ8byXuifKOWnMunIaD2M55oY9MiP9fvAxhSx0RCfAkXXxLPGfn9R5
s4bNUMhSSNHY9l+0MfWqDDnPMQf1ILVVjxZHQpAQwO/7yQZJoHg0R7sUM80Uuk4vQ14hRW0vkMgw
R9gqZ/cltrCqNliULutFh2WyTM3DTO8ykOOIsHzYdSh5yQbDt8OrC2600HHOTrM+mS1myUmNSays
m0NLrMn/Mbo1Ne0BCiIFJxqN0PS1wc0INHzHp7992sFzL/o8LrUKx8UOZV/nakg2emAd3hoAPI39
raBpFfY6JVf9mg+LeWqtHfrQ+CCx6bxtgk4AN7LKP3+auF64Bw4PTqQqlQYe08F4uVoAh8wQTSht
BP5xzxU6aIjRtyawL4RRq/Xi30r2xb7o5w9DwpuywAdiOCrnEdQi4M/AmRNVNtV43s5dEqkxvDh6
t4tSdRzXH1SysrMJTsqe6YvXfVcOkIxHQYPDdkZRJu2gBF8/789em/6WLVQOyKzQ2F7KnYZU/Jl/
p48doia0loFiNyLL3pN8zZPNDZJP1vbN3dppzJfGEw3Lt+2NnkA8KuQ/5Tz8qfCOmZA3puzh/pjG
5/lCxFGFsREgiQMbkJzRQzM/vYm2MWlEEI6sLNEXL5SKR9dw9wsQEown47PJjCm59wquGsZFL2AB
uAFrbl2CjtS+UEnBKmMVaQDLNWpL0qTePzV8rwaS7Q9C7B8Lc/vBTMn8s+4fMjB6cS1vaRS1xzD+
sh89QmdndAeQ/MLV4BUMJ30reyrOSYXAnxNTBj+Qhe8AX0aHRZF78KA+t86s5T+ESQf1ixclT9+6
VHyl27DxnXcO+pcF1wUl0thosBLyMEBI+Vf8gEtaqz90gAqV6fOYhuW7f7tPW7oK5B6BMurVScnw
Luxww2sJGM+M+5kd/UPbXvbZHnGN4P6TyOBu5gRJXhYPCYXxM5bnjy95VJMf1aeV9aH5fTPUlVI+
Q1KM0cIpOP4krdNIcAA0rCRKDMx3qti79stkPRmQ7RK7BIrOtXoYZO7JtLvMpz4X1v9G6tc99WM+
nsRTrTbt48KEg/PTgcKPR3TETJIIxVUWHC9ObRI/7CX4AykHl2J0DgljsCCnyydeucd0TWsj0ix1
hPW4XaecrOFMVhci2K1fB0CVNp5FiFXCY/uyvVmHRDiSYTOys9+rWn/zTU0ZIfyugY09kAqYXpbf
ZDl63fBOTiwc1MR4e5FvAd9HVHLTvyYGD6pJtBYQDr6alVQjiKNTHKB2cgLrsELLPLMfW94eW3Fn
8vqMm6xHmCmjPP/H/K8qA92r0ZGPnhhUlMAT0VlmP0Y4iXWHt5sdiqGq6Zd/U7PvA2vYIHeRS7Fv
tIdI9j1WaRhPxyyekuQ6CFFRHBM0To+EEnmtfbSksAZ4E+Pjy1ioerKg4hbFu+NqrmxpBjztoFVp
2tRiHpcIX8IpkZFz+aB837xmrNExbrr72in2eQhjRqs7+maSUOUhAMtW4c3nFh18CIcg/LogrHAp
JH8KpJd0by+l0zonFdBbjf5WDdIFMDQE8jXhcioX1j7YoebHshgpRShlXhwCXScRDUXRiuQCG9Xy
nD29GC9RuFQM8h0KcA/FoVZvxGWtucXmbVVP0SuIn60gK3ilQzbiWkFPKYLKzFURcHquOhNea9mS
9xnJgearjYNeRtha5YjWww50sh5YRbbddsDdmCoced1reeFbR5gQGbW1s/8UIUw8kGj4j1ANFoXH
WWOzoaaFtl55XvoscJnGkEIcoD78D+dUzi7mtNPwkOAvWMfltgq8SE61CtHZMZpzKRQ15mIRMa/O
DBNx+5jCiLv8jRDZv77feEy9vdsSfCutV/Xy8MpD6vlY+4bE/8sAOaQLHmld1DQ+QgOwRqPsAH9z
Cw9q/aH5HIPNiN/0s84itAOSn1RTU7qG/fJSOlJowTT1m76KB3zOJ9+SfyMAI7ElNA+Vfc4PWMRd
08N0ruCU9/KZNdEcY5cXjte4UJ4QXbEU62UJlrAOoFQQwXmtE7ZL1BK8q/MZObKmPwuqqo1XxbYA
PYPTRhHxM2XIEvnlcFEE6nMjrLQq4iTDr7x9pi27K7am2MkEHPlBY00mDoABn42Fs0GE3ZMdRv8z
Ss3V65Mu/AydNyHLxuVRSb8AmNRWEBkwrMCBc0j+9OzB+yHetpjMEzG3faoME9U7ENa5tJhK0ZPZ
YsWZ9koiYjHMC11G+L4TPS0qPQyavQinFMuw+PMTIZfWfuPwZ2FlyaUQiKg8k9zdxC54wwmC7ndk
aQC/6SOxxMH6TBOJUNnNQTsk2+Kn092/amgH47PaC5R4HN704v7XPXkoRrHZqj4fhrUW031KyLAC
I7W2TTZ4dKP2/kWWxgwsstEbocaE3yGa9LzrlAMzGkvbV05cll9fAFNIxssJvhUmTbhzPTWuCZo9
1ROdJDVqpOUz0ctBz6Ha1hv9wqJquMdiL72ynIa175UtNnNlku5JNgvqBvRLJNCGFmngopomxe3p
Y7eSKW6wkPDJzrJxmhmNPFlzIYI5Q9kxJ+mwMrPO5ZadpT20YhEl/aKQlgngh+QPfPe0S0CpKrQ1
K/bxqhdRKT4ow7/f0/szEABpRI/VjjTWVzW5nZyp6atPofEiQeAXzuO+ujWk/HBqKpWY3nqjb9FX
GZWwGVUFaHBm0SjFua3n8U9iITS0sv2t1Ve0FvmHi9Oi3nFhQyr+AQsj2SNYhMhmwOAyIySZ0j+d
65BpXOchcFa8d84+/dB9JwCI9gK3wXYFp1mPBaIsRtgiDxOPOjqWW5VVcV1ftqPSdBuRPm51ZBQR
zT7/Njhb7VnA+nUHiPmEqqZbW/NSzajhThZ8tzFNeF8cH6DBngiUdDU9zymLyHpGjKjacXWzV+cq
welRFUemgOKmrZvGBMIndR0fVNFyjA3+T4pnmvNXoCeo/RrTrZgKKe1jToxASu3QpNVcE9RTAEHd
HPsYnTqpWjtRm+ldqmihW0WnOmp0bbesMpAs72SQJmaYUVYEMGVgV3GkU4GQ8U42XBFjRfTkP0mK
JZrQ/VClxMfFRp7QIY+LsUdqLs9VAMDUux0LI9ID5rw0F82YLN+uYXXG7LwKgV7+OJjfENsafblO
GXYdQO9914pkAihCG9jJIpAI9LxFlO/mzKEY0D2HpEugYhiifBcJXpscmEKN4m2bnuFT/Hf8Pccv
Kn2NxVgJC85dqUOKaA0xMI5bohQMQaqIX42gSv/L4adZlNlyZHKwAIZDDJWlaS0D/qyohh5KaF6G
JMmnzqy73pA55WGtgr8eELnPxO1lmwnfVFHZGtb+grwVdiCQiMXMo46aYGfePSvHtYmXw++dCrod
CDkZM6ln5z1vgsPEjkUy9RZtWAynbbBqNAPlhGwYsDcIFeMM2xQZ5GfjlGjdtmsdKedh61z2l8Pq
AREiedKXvPWCWtEafjwb3FG6PpctzKEgzdPP3oU6HaJ0PW84xqybx/Yh9orRoGtBA4eaQ/ZFYBtP
lW2bcsF1StA9JZk5WscpkMCERfrTZZ8m5wTFTM4xAYk9W8MaYmt9OvYPxZUA24wzYevI1v7/Cylk
ZkSE7MloeMzqxiOWrLybiqxxOkrrSThUtoF8+YpOmFOOYFcMSoUYeRk7wGF7izGHJMk3XfjsJR7h
5W5PeUOQhZdXrfqzSNOjgSr+Pn5UcBsq9VnY6S+iSK2Lf4Hrt51mihBx/8FaPyajezE3ltlquMcN
6HScCerObHdZOcHJsDB0A+v2LyJWliS5yJvVhoRnEWjkM3348Cf3Z2WhO6hqdVmvdarg4JR/eLlI
uvmdBCvKpKbAjXc+A9TOWvRCQUOxPJ6uu32pxdfwJ6F67IABO1nzwJyizUsgvVDBiir12eJJyK0K
0/kiUDLq0r7zVJ+EXc5SHgxWq8X+Y8HslHlZxEOfj42pueaxeTssqXZHURXOFV7t+3z842O9GWss
3RpJhhXu/vQ/HgjFTvp7AyXQJQweCoZ7Vmc9XSmai2Rn+DNWK4ysNyM6qsI/S5PzXuyIgExaHXu1
eyNsUHKmF3PGTynHW1mAKGTLaeEQlhpO0/URmARxrpfTht0DAgnR7HOm2czSKgu1XiUSxlIhtAzz
dnvj11AYoQrzWONyQcKNaAl8Z4ok9/pAY5r/riUR5CHTuE/EjXBDFZ3Y9Qt818ZLrvXkvU5FP2vj
81h/0dN7qHb9WHnubfVysdgC/2gUhEW9mNZzMcZNOUEyEwmrOVJMVGuqGz52OQWHxYw4YsC54V3j
LNFJyF+MR/WgLhTtppbVRrPxMBqF6u9NvRMkHptpxHNb1kNBUbAs5nUZieM0wW2xkg05Gqw/b4dJ
vStc/ftR9e34JC1TfxHI9UEyHqvHMYLVmrO5yRqnHKfW6MmE4k3dJecuBn41fKi5O5C473/9lpxs
tcV77+PNT9dVw0RU16OoSiuR3uvG/227uNrBcXzIaQbYOsrpAteOe+syxMuom8QlY1M8kLu5kBZv
860PWwaB9GbQ6b9m/c/zIO/12rz8DaMjnHwL4F0EO6Vg3C86juMrpo5p3bvFuguXRuTd/Nm8CU7M
BS96z+nGf3Ndi6tfoks16aOmRcdNIMTF6Ue6YdPjabetYjGs+WQl0FJDgFcqFMPFh3KDtB05w/yT
VDeRfKSrnBTADb9KUsc5X3szdstEDCR85gEdHoxkOSIwp32nrU4OzyNW1HsI5rbi0jmsSqCJTRcT
gTEv3W30+/9vvhKv+dsU/PjYMLcWvp5tOFypG3Pgj0RqPc8M1iyHkfIX8IxbSDnidrrwMidlAkbM
w55Zw2eEm+QbPLoAHL0LQPnL84TDxJmX6p5DRPV9ZDjB69x1DntkFe6x+a/hxaga6nY7vR7H5sNw
Kg+8NqSvzqunCRB4dX/ytFjgzheRLxBBPz2J2yy2yzhtS7u4314d9JDl3NFIgAvrhp2HqeYvKHVs
6zo84UlQ+Ujknvh/pVOllZRASCMuPFfRp9iZwxsqGcxHNf4XqwV1c0m2+h2qJ+WINsoY5vIxsRE7
zNlDpcZNdTuufmD8/tciUvBSgt6/SiJRzXLtXpyixND4lNs585ZTh/BwD8N5ezk3R5aQwkrrsBgK
UXKi68OjZcfSfkLWJIfdIzD+uTn6LotWPFZDMAsTmXbs9QKYGGt4qqaGqQKlt+tYWGRLDVNiQAz7
s71cU1HVfh2nXTD99uq2mdrnHBPnjvd9Y0Ij4ykeSKhjeXS/ruORKOQlSBGtcVcBTpqJ8VyBINZy
91Qgy7hAoXJyDoucJyZ0ICZYiQsofuvlDJaB++bn6X44iG7g7ElxRu+VHkzqsks3vk20OGPN+zPC
XqZ9U5YfMhYWpy2BnpyX6D/43LujdawtDb7BKz5M6B22w3pRtJ5aQOX+PVxSITpf0ylGFwmSAFgm
JAwvEkNuAOAo/x5WNhQUzEAhjycIFqapMvPj2Bi9CWF77p2+7dycHY0gnIrWQ9X3SuKBtWQX/7RD
KEtdHmY0TXhP+4EsiBjRevC+LJDJuf76HyfnYrgWSL+1EBwyjkrtmXrw2Rb/eVZXKaaTTV6Z0llz
ff8yNdHEsFrBt4dJJGs66rdDGTgw8q3iotYELFbazVKj9INj3sJ9B+fWtxEcEN2djUzA6zBa0gHT
azCQlwsu9YIGSsIfICNRk+D2XimCg57H0m9WpxLiqOpKhqrh/D/+t8XLhC7KtawOsctRLi3jqq7Z
bnWOw6oat7Q7pVgsbW+sFmBzABmPljvTrm3ktEEnXwTytg+WbKaS4zYXmeg8/L/eR7LLPlsFGORm
uskq2mzC8ZDm3XAjAl+zlYMrzc7bMwfCcajFq+wRjOmChY/EfmC1MmfQ8CQINwJF4QvXBspA0a+G
5h25UNSttDgJ4AHJoSbMCzJnGAXaSYMRv57qikFTD9HQQqdx0R1dklaibH4tZNY18dO2AM8cFKkg
w0xlRaJqsxN2yJsODT+HTWca5dtD+cfexxMwyPaT1Rqb+Zlm32VbnfvNS0SCAT1euVy0iotmVmRe
8YrkR+KU6HTTVJEd+YY38uiXSCSzZ1PCqQKhjf4fvzAjMVaFQf3xU0rBTYgTxt1kOq0KY23wgdQe
Mm+Uc9AHGJriYo/sG6xVU84z34aP8P6ewnjlYrmtyQMRIzFFW0rhWroqJW8Kimx95ibNEK85f7Vr
tME5iedTPjvVKlpHeEJjeu6w7AAXOrvdRWyBeRWlKMIrFqTpSUpRT7h/MBlLntTIuWu5ynZUNvwC
Z6g8f+UJlTiQL1TXAQ8H1wNzKNOOvJjjf722u3jv/nMGOw7oa3lsr/VqCo60Unec+HXtViCBRexN
U5gXV19n0vNnD386w25fcY6wdssKK/yaf2vYYLNgEhv34sutBaQ4MunHvGjfCXd8Tyj3aEr27bHi
Y3Dsmyz0nLnQyKPdg5SITGrNkJSt1CuOkJir+4Q4uz6whYHQthACk3BroCt154M4x3XnRpZZfWdZ
sQdvaMROWkmc+SsIaTH8n5OxhHPwAFnEYy6BRFAjUmc36yDONQ8KHqc+HyhsrJuRrlCp3dTKmfNT
oO9RmPras/a77NyUw+3aAyqx5g2xYNOAhK68PSTWTaa3DLWDRl+yh2vuExCAi+G02yEZGime1rQK
od28Fkii3YjeaJWOHCnY3e3UUGcypRnxDGZWNBHJ6OQNZwxY3g8Kzt/KTdi4n9yOwT49GOSMnzBg
BRCQ+isRNbDNSrgtNeWb1e2AKhPZEgb7hXtzuZ6ypLviy+oSMg80IrSGpEO5ExLwIjG0/dTPAeGd
XulrVJgBXD3wGWpedAMt7bLAiprlesq48w5orYKBx/RAvOIESKmzSpEJB9qo+oLmC0wPqIvyLTVJ
mPMnqo3A59okVzLITI8JTa1lVlNEkHzbokqmFN/lRX/cesX5LgEahA/9Gx4igUgK5NojUHkGUUCx
G5KPbZGtBCj1iULlddaVko3FTQZ4G3iT5h6bYcki7yJtRfSfZf+XRnXX16Xe0CnZYWwFC7b7unFi
atv7q0TG/wYcmGDI7MtvfwM+RQB+hpQ1evl3RnDeorSwSHphm5iX34tbHg5mcHkCrVf2Lpbdsxc7
gnRu28eXxSb0rTt1+43LBnuhVmDbQ6PPawbk1z4tPIlMjvLGJUBDPw5KjBK3Yu9Ws3wCE+/8zevl
Unf8jIFVJxaW9g2Yf/LzqekA2e5+QDgutWj6g+5JBop4tEwAR1LqIuT7dEsvoF/h4lK63n5RdoBT
yMBVhTrF6ryTA9EsIJdLjBtRIf3QghWVVHmIuMNq5ERGyd1g3erKFUAlUhIV3jHbKHzvCEG0coIE
iJ+XPQOHYYkvarkMIIDzmstpDRCXjXWo1d9jjjW2C02nD3z32GPpA1ymtELQJpqGa19mdegFzhAU
uhP3TnfApb30a1pbw57HbVRHwAzModPyIYIww+71PZlCc2UV8CT+QVn5hbD33oRpYrxG11Nm0pZU
VH5jVCws5ssocaom62yXuC+OxwB5YVkeDlbnifpuElJz+mpVBu0ssyVKORKtO7xCcoW17udXc2eV
OY2XlPLet/zIhpWMRzSlJtuuZXP9vvBVsbRU/PtzKl9f2b/7Nq9S/7qE41Bsqjq/KM6k4wRffeb0
BZfTSjUmRS8qA5/cesJANfWQnGXUviWF1wNRjzcl0zasyrPf8Ep9bco1VtmSeHgbrg3gs1veU9Cx
v+lHMveo189sD5q5/vvWC9EECKLelFdIgl6onpSqb1oxKd5q89A0nqPFXL+92RV4RP+NucT3bFVw
n/3S3Wp69bSdsyXSsjJUlh9mh2wYoaGwkPt3E2A7f7HX2dWo6qwDe7PzQZUc/7JwUYWFn0K5XEzh
UEd4cLWcAtfpzVcTgkaYYYxvWWdAdrQ7WXbTy+VxFnYSe8VhNYiQXbXQ65xD7u1XyzM/nqd/AnWF
qm4Yh7HWUSqsYtThi8F4KrfvmDS3ae4HZHs66MWKGz6NasUSZuGCJ+sXDvSEkxzKqsYQ9Fy4GgNa
7sRUEUN5tVM0/ABS2IcY37J01qq4MJ5CCI/+DCyhSibQhmxZv6W8+yG28zz1S2+ULiDMyG5LmPqO
nC7D5roiSoOMFZ9zvtMEqsm9R5jKah+wBAHp0cKfB4U98/O58a5vdHNYki6XL4TSgraBBdn1UcoR
N2pZsTtG13GGmjOqNI0NUhLXekNhqRK6HKryvB6l16jCBAmR3whLFRa8KhkoYg1z6n5qKuAfizV2
CxWX5Exef4BXlWHD3AV+mriWcEpsVVzgFcznR46OZjcev9ZVR/qaeeHFdMNtuJZUyUXpdtYKqHKj
lHlkELHKztL5nRSfj7QdkYxAhpHTrR6iFEyRr9evY2ai4arX6xv4an0cYuFarBHzAExCnMaHmgfp
2x0PKpb9NFXRBn29a0S9ifNeup9OP7QartuTwbvbO9+6oH9BX8pEwfugcVLvtmG6EAGaHQ0vRXmr
yLM7IKQyBJmkMBGCv+7GvpLRscJmAa0alpsKDDNenJXae/MUo/APLlgWq2eV+6FLCUjSGGFLbPjm
1h7Kjl7pWA8KtJBubsFl3pAaoQzgXKc5O6OyR9qGGGJWEVLU1fibIY/6KHGYFo0Hp6eWWs8OlFAW
2TeSIOTGmV8ClVp2mnhIvl74dSV1m7fQh/jWxbTNfrFdKOkQJL+QB6nSy6N29n1qyUhX0/L1jMfY
92pFb3AL7sOFRpAN7tv9FLMPtnKLglBqAmtV0uvZuQb8rkyDdT0yt+YNHwkmGd+Dfin6bdfzGVyt
Hkii5o6rVC0hUZNtobI+q46N3FG5NbjkkC1I+vjyjxF9XiHGpwG9PrSZCt6q4eQdvlDm5FF7MPll
LydR2ouONrMz2Zjlegm82QTnRfOZ9qMGFoAYDlu+8eV0yFuTygxJDdJcV1qmKpIXrVveLCq4lWHA
QkQu8eIt7v3IJ4z8i0dhHBqDyVmTa6BufBMPznsoDl+mJhkdBuj+yfFQNerdG9H0MDcM/BXMGLO2
Ern8Ltl11X/gTRq25G+Ifkbv5kD9e6ZEaYfKDwXxUTykyUk8bE9FE9fa2B4PLr1SCBK4a3JgLneg
aBZESwaDmx20L2G2Oy3pRvReu14gum10com+c+JLICh3IYkrJV0vgdHpIPk6CqqPK5mJwyrbWQru
nnKU9XWKT5JcNGqIcvHZhBJpqwrWvReeszWZM7rVfQ0bvftxgf9k3Fu3WwpfxMIKpXQs6CnDzWst
ltKloyp4JSQs/n2xhY/bl4BXb8ZAHDZqxOWLTqjFOCDzrZyvWmjBzi/yT5PWvaYh4Y05/TCEONwm
/oYIfegI+fA7Owqh6usHDjnzsvYzNHELPn3yVa8WLlFWQ4+5EATIIojQCoGfZsf+i9WjHp/pmXbz
5DfyyEgW2EF+7YPWBpsnbspxZj3WW5tGNkSdIDqH3yCriHgX6OlKAkK8aD/q+UUt5SUY3VkL4Bg5
DsKt2Li7n5RfIF5iZFxddr5tRD1vGVm4DgUVV8rtcCaZdarOV1uKAk4taqms/pnx17QV5TMP152s
zkJmoU9JlQVC3CssSxRyiYcgk7bbwakMtmFZbD1KKn7NcRd8zo/7YHyT47mBK9MoqJKH3uRwXjUa
ismTLvbGWQ38o8SnuQKrFokeQd64UmrHtY645trZl47V3Y0KUGr5ZhHJHpDf8yGT02bo/Pj39BhL
eYBOO0JOWM0TP0qP8p4aCcdkNTlqYUpGbGoQ7MBCJlvwe6m6+GXx7XFT/CByn3eUvKEn4mW03gCo
+bwGCUdXxBxba4eeuKSyQwVLSlkPhsxNQ70TegpycEK5GMU/ataz26i+D19//o+hr29xmFvzmZJo
BM+9LaNojK1uyAXjBSucM2l6Zy5p4YU4Ex/v1exdItY3lpD4FtRASRDo+o7iayrqZxJW/OFtl5ca
7aVkQDGs9bnaNk5BVIiC5UWp7ObgVWKlaHf9EMV57VjftfNA28sWB3ANbuojSQP64oS02oNqlqsg
He2LCCUN6M/ZYmzIao1jNXk8iMe2ql8SUGtyeKDT/sbyD3nbNTXIGLJ5TiGDXFbHhKINz9TJYeL+
hMF8PfPRAhTYAbaYDiZXL6j8hAq7ZNPvyERT8tNwwZJ63jfuVI1oGtEc+FxXlgUKW6jJlDyOry6c
YSPQl8F28hHenXUF0VLo/3UXHB/IB3rOObP5hGVkvfqFWdsSXBEWCzMs+Queyqijq8e5JXV7/3tA
+y7Fx4j4WvHslKpOAv2DvernYJ5dMVBM4oK8A44DHYDA69/Bdw1cv8nimgDIUbBIcTgbiXdSSxtN
UVVo4+t00FMlB5uJAl5lVqeUqM8PgjWwHhiehm2jg30f0fPLEatXwxiSg9Hy2Xo1MYU1GtwlMxjo
/eiZGWfQ13O0Axju+v9G8tZaJZzS/dGvQ2j5SCGGiqiSqHVET3w+k82aGK1fRnhSTQTCHMtVUdCP
t7xSjDBhkYV5ouTGMZnOzvi+1SHp6Jda6jX8mtXtqyAdod8L/bAicGPIfFLjizUy2LdV8c4zAA80
ZhO30euqIBHUaaoTA0HoK0/1ypVhTkW95BGRwEl92YVKmZVNKPLhpYYTDT7qOCu+jIrgegQ+sdwW
07kxZMu5xCmafS6MPNmXhFmEckPGTHBSszC1egTCk4d2tbhH+SNLmpPq3IGUbUcX7Xya3tIzcgFC
j/u6eWVDO6Eqk6p/SxwaU1/QcPqVh7xo7TFXYITFmXVvX3nFMO4tKx4Q6RiC0y5vEryXe6MrUhGm
nb0TwEOWXI6BeSQhSwPYPF++afDCyJXKJ+1QgM+9q9gaRhZgO7mwFheCwS/wJquonUni9TGHbHhv
qwRgMANOBKo4/FgfOAywx40q6yoxxBMGDXNEzBVm0oo0sPs8DM7TMq0Wu9o8aCUl4i0k7iWJL6Np
ZSHgtCtUw6rTL0NigtjWlVZYb8gCgiptNW8L2lojXQcawHPwWQgr7VsuR22zPzO71pMJvjwMsfiA
aBDPOccDZ1iqHoDrr5QDUynHiuDK5oMf5JfrLcmIyZN7pK/wP6C67iKqiXj30jA9jUWRfaWg+dFD
BkPGhj3ttUoYy+5uDDBSPQBmpYCi6Ma8VpL2fbR/FkMtRIKpRjzcfucOSjQ2hs9WLCwZeJjkk+cn
8uzrnPnfUS679gv75IY4T076mjoC/lw+adM42yE1/2i4tPtYmzKc3+JzlBVgByv8vkHBeSLasw6V
4bto0VxtZTUXQ8I0ipHGwJGDRsADaFF6jK6DCau7R1CbZak/CkAYkidjTSG1mi6yXOxDhNCx3vkN
E6goh371MGgAL+OgehJS5ktjiDOhOjSRYtJQKGyiPkARw9bBmUUiGSAlOZZWUMPjlrj8gTKMDnRS
tgAW5LijGoRqyElQLNbiWQ/nXvYq794LJFb5KrBjMh8tvqBl39t/ribW7Raz8TIJwJEWiNmzD181
2hLxIH8vD7BUpoh3KLK8GO3Bd4gnQ0uOtsIDiRmkggnjMo5MSVrPpSjhs68mTGcogMiJWJxGM6HJ
chb74Rx52yfZ0hASxsTG0gpbtrBSsh2GCfzPqZgw2NIkKKsl1mqaTDUAxAp47LSeQl9fYtsQw2Qg
dpWG/NZDOzom8L+kNe71fWSitmhDWvce7XlDLF1X1agF7l2fkErneuwZvJJlzaKsRqTzUjhyi8jP
SdgGnZ9TTvp8f3GM0nxteJcD+s3mLgIH/seZqsICeZnTYeMuS65u/+KqD0Y74qzmikuyjYDN+jAH
TQecW+2r4vqX+Otqt7RE1LZFovdg8vzJxlt1/zA+VsL576nKtUw30mgyIBZc4lBFJ19R+QQGfLEy
mf8fZ93qdfTKxiEsLg+gZnC1jvi1wmACgSWzcdSIcQhuS/rJWNC0xfIXkCuWTXZGGZSm2zUcGSvB
b3es1W6j7B8ebISl/rKWx+ym2EDrVp5jUhX7PR6gyzjOwaNenKr2zhqLJQBrW9pag2inVse+5CxB
Ne8v6/YiC+XyHhjBbvNWFRSp3FvLSv+joQLnmciX8K7JJFOAUQj5/+Fw1l8jC3x0LdlG2neUb6kx
SRKG/Ux5TBK3/kVzyztyYn2yHKLjvVi+8BbKzw65lem9TJlywB2M97oOCAJVDeIyp4X6hWttsSYu
5R6algi+sgz9mjQmvRQbE/XRcuW0aTfneMQ88z/t1IQZ3PVmDmevyk0AonK5DpSlhz/t8HPzOHYQ
p38mbKEjCUly+hCAu0LiUlJHDDVW+MgmDyp+e20/S4rXspK9wy/4g0Rck3ztQ6rSLqrKYYPsQq1B
FeTYf85l7vudWq3FzC1BKm2UGv7XLxNbdVRw4IsxZM+tEvsqRWiQDWtvGWD/QA9qiiqz5Vm0INxA
aU9lrJQJ1uC389yO7D3aMqXtVDMg8OCqiDmFzmC6He2RkGddacNCGXkh5AQMNfURIwvFQ61bUJmV
J0iCnS6yBJmlAJVt+d3Kl3iOwEKKdCV1yBXtas2Zy+Wd+uvEIet9APkSCjSC0Ot7Jo1Fxrtub8p+
ha9jzB9Z0EdWAAbZmZs27+d8seL2v9O9SGzD4DAgdqTfFfHH1eSCmqhFKem4ou7AiygftK/9jJir
cQI+zpKD/raDp06HKVb3VkeSYczYyH27bOUu5VBaNJ4H7SRF7lSe5Z7NVKyYRrxl3KMHPoFxR4E1
7+GieTMRY0fXJNAWgtF2vjyG9LsdZIs4RxMQK7qNX2P7ZzDx1v9ggodf7zWDAbkVdCWQwNSETrUF
03xEc/Y6abyPojw3KtQ4Ip5VLxDay6HSgLBCIoR3TLk2t917ytXSbpy+wtydXbaALgrH3yqnKDFt
YcQWL2Vfwx+xbfKG/LjkcqRj3tlIf6ihL+k51OHvwRgan0RWN8CM/ud84SE2wyEsGUyydP93G8MV
rui0/C9alqLqvEXJolNQVQ6JHy6UHPBSWz0GZoWBRX19Wo+9bAbma4Oj3hVhOzkisxTyGZ+RJKBk
jHDVePHhUJw9UahFNbnU8CBxFZFSztm+jXFQP54f8HJXxLp6t0iigSilTOVumS+zgCF9O6w/oztl
qnMPllotEY6I9xLCApo9dvBYcTqvVFeg0IMMzEVG4tJolKpzlgCbOJg34Uma20FIjy9tz2Q7xdZQ
x+J0PijnVXb+2ZmuSg23HLhRCz6kNeuPH0h9H+2BwfNtVvhd/Bbg1CopzpUZjKhuhpSJ0EJPK6OY
YKhr/B/YKrgKyCcxQCNfqLOEBLBPvkhWp6BT5JNgPnhybEuJJRCrytNDfDnONzbx3Yi2wcJxlE6N
srcT1y2wNcHF7OxC1zX8FGjMlu8Vc4g4kXXhwMPhPQMrlE4Ej0EdgRZVF7ieK4DIkL2gkrao7fRH
cXtm06h4shshWkbKxGo+NkgiSg+Awg5RgFlfYw5Bv7BquXXk26WOHYP4CNHo/VOGH1tdiPpHnhKE
5JTU9d4PuwEygR+DnZDDmnIZ+nA8ThmcMrP15J0bauCy0u/Jl+cLhtDiHmn/1NegkLp4eQBUnTom
ARi8WETA3li7YcHTbRmRwo0Fg6pfHEx+j5dWO2dytVnGd8VqYeKr3yP6IK+D0qCO+8JzA+nXCnFJ
KUsl+nsK3a4YUZrMNAgiys9ULWWyOEvX3pMMnvfm+9KJgfGFh9LSGz1r5pLkzZSIMt3/8bNqxqpw
APNyw9oOybPqDqK1QE3FC8mamqvANK0j+kUfxFuggo+eDxNXw+pCMQm0ep1YpoLbpEZWm5PRYEzu
a3t0Y+FkUVweKrKYL1VxmvZPduxjvcnj0eRgidjzzyj3FhysIxT0PPacYyxZcm6+eFKVsmez2cNk
kUonEHbUFgkheNy1fNtd5OmBJ8cEqo6jZ9fnNvV4J0O/DBNawoZuJDxyeqnAcdfXoRC+s0sp7stU
aQkx+2mZsg3JIDuJAfe+KHu/V2ve5XMfxbZk6b0BgaTQkASnDx9qfgk8tOHv+Jhgmvzhf+xnjUZa
f9XCy5R5SYvLKZ17WmRTJlUtyvrV7jEO7W22ChwBlQTxu8O4gxtpcvLPp2ovx9gA2GA4J5tqD24O
du+vGAnq2zwjUehyyId9nyh02ghPAuyEmOJEopwndoO8HfprR5ukJKF3dsTrwSA2fQ/mWVdBjgki
uNNiwiVvKus35TZCyiA1SM1NCPNcrjwRwvth6KTpxzpJRRoBNaLD+yZNddgBXGcmapKelqqzmlxM
EGQcSXy3/brJsWLopxA0GujrILiawzbd2EgIc5PXYMAXDnEZ0iiOvyKg6zaA8MMd9JJ+zjH1IRdP
icAEqHSEoGygcTUi7OW1VegMe5EzjglsgUfA8+67Nkoexocn/CRwnvsZu2+t+3rDYZehfTg5AX6p
9ZODqixhneGglqKamv7paA/OqMXecs84SD2+nevjjEYkzEzULqPNl1pKrg0LMSNzEHqiZlGkLL1C
qP9StTF3/EaMdLxeQmqTlje9okxHYhWx8HhfHdroDlhijQU31P5xsT1rpUyTyFRt+IrL5mo4OLtJ
/mnAxAVEcjPRRRpOt+gaRhUi7ooa5cZ+ffJLNe3ShAQGEq75mlgPyJGDxP9G3o0uzcshRjZISCfi
bq/R00Y5ZhgeNjPKFT6mud4szAUTZFxvh2nAopNSnzKQTb6SCX7QAukv74avgbDJLSY3ZQJY2Tz4
9RLwYfNTgNzkGVfO9CM2IaNgZl/kl2oTEEGlro6eQwjoI/MNlfcndSSKeuOllIXnoFIH6rkS/Lts
D4lIhEp2VuS5PGNh7rLdvi9qq01CCUviyMn3rcMgzBBzr9NZf2PT2huQ+9GteFuNQ7xgiuu/+gjB
kitA6nkhp+zl5DerNy8fw+9SlilIIOJLqqOQey9ZBJjnEefQQ4o30jeGJj7L1Ts/HZKVfn9N25OP
sGfIX4GNVq+SSqh4qk37TgpGvBaimsNY2FHIWfirdWG5NioOsCmlapdR2U8+3Djh2QID5+2Nb86M
IjDV/4AHUkPIbkX/MAbE1A6TaLjGkPEAG0G1HqMYnDltUME1sElC7xDEEG9jsyVCVVG/XnQroTaL
6V14syclHbRQK4iTmNJNplHySMW6HDaoTTDX5EIkmZcmRW7bQBvPX6JRB3MkRYUN3VSaWO8kZ0kE
Co1dm9e4oXwMe3Vqx+TRGp+e09lfmKVCN1BMpJY/aW0z7ErExAeRC3cMw/3zRQB/pAAP7+zYIHXG
+bne7yoBSsE+e+h43eXd2oPdXaDK5zrXcaqZnJI0EZe9iVB480GpjETJNp0uoPxRd8pZNaFVGdIN
q2kKMBFKR+fM+bHzGvq6VtmmiJSXslKguvPVo2SH8zaqrXpOSXrEyXhPpLEf/2p8e1nO0ctd5Ndj
hQ1U7wDpg+7d6LxLujLKPlaXD5rBhYo/ElF+A2tumk3ikOoF3pZF2c78XOAjwkWRrw0jedgAHVmn
eAyZ7wopZjC5+mQu4UdtAqct+zb1pXE+DaVOMyqPjt2uQ/tnHU/aCJ04RfYMes70jOpDoSfSS0W0
AYZAwKB+sly6p7ZiiyGPD6sQtRide9P9f3SUkEe+QI54ZgS5bHGZfMwJWWN4mmp7LdOjEeLw+N5q
NGo3ae0y6/0R3HrTAWu/JJaaqYuPCwOJqeoeNWirhsvUB3rvNl/W6eJA+EvzqRKteG6btaA81w9d
HILgvDjBXhWzPGy1/s5ZRlHMLa3jQfjFh6XoluJbqdFJVLVz/dMX1r/aXhwE4u2q+V5doT1LgG/r
81tLqixXJV2nk3lkAuwerauGQ6dX9yhFAxmdHJ+ffBD8fk2lTdCioXL2phgpjPYNiHtUxNgFMus/
LP2uC2Qvq1LOtiItM29oSCuM2/LJLCtE56Ti1kwLKIDL+SPkHJ4NIUc5cPB18Merp6tsz0IOFvyu
V9QJkpzjt+0IbKyKJzSofwexZ6QWtX/37fok130i1Nb0Z2sKbppERMXSFcgoD6CL1AFKnw1yAqT1
B3DO5bbOKqzEqshj4QyRxMi1E6SqEMYm2jRZkW4SKzpWyCM1B7M4HtVM4Hhlu7qo4D7BBJXaBW5R
GebvXn57wtG37YoKP+AQ3cHvsOjnq0/TjuPk2WBSTllfdm1/bpY4obv8SDSa4Q5+r8ZYIKY2e9+I
PJ3o1dGtt9Qtbt2Cgd4zadVGATa5sC80liHtmhR5fgjbUEPwImkBXXCqKwMYfb+VXSk7xgPIjlN2
1O5UjXOdb0VH1bENbaj96CfxJOvoZANYOlehjozUQ0YgIQdpliBFrx7U0d1Bg4tE/ecyFR9c2Yao
YVELLpJuf3Wpm0FBPBBwi/gsZwGvlTq9Kmb8ryDBJATngl9dxA7fQqYeR0ZRT2+pU94sEdCww+Rh
wbDdsDmkRNf2k9AQUwwhJvNiqwiKxH37cxv0cHM3P4BKhHNSruOjpwouhofqC6SuPq2CXcRowflN
rwGvuYxQFnhSkXETHq6oNXh/IPYD1r/XU4m1oC0SeJfTqDfXDngk+efR34P1Ht5HPlD49AxDhqPI
vciq6IJ7NLuGr68XW2m7lFcsMfgA2b6/K14ykpYbfpMAh3SE9r7NhZpYhVHUqnqKWGMNgFci/Ec4
Yfsx6T6phHgKwZy3fNWTIj55oXxqoiUmb1Er8aK2MlkT3CgneSzbTiu65Wcv0iKETTdq7sSxtae1
fbsyl3fKwdfQtahX9NBEGHzgAFhqgcai6rqhXBGz/xMgSyrfsxk/omJUhhzXfvwgxbHWt8/VXfkT
nJ/L8+Wrhjz45DtR0oe7dG7hOVGteOLECOlhF4/qIg3lwqtJCNlIkMRW9CQmcn05ShOQ2SVIVRIu
W37v9DgX1MqN1Mhpoix0iIBpHSex0J96nHEPVk47icj4dqtSjHahdbxxdgluc2fWBCckfP0l7gUT
rrRx79ZYv6V7onxuwgqfCiJRKxs2c8Xgmd3YBcdG0eirL4NpYZg6IvvMGS4maBAjb/ZqeylN4Rw3
GLWGwbHSw4EbEMxOofSCJEKGk5kAc9bayvOerHarR6l5rtOc4Wjpp/CaHt7I4YZk4p9X4wv6rKbp
1Wh+gDxkuwzomLKUdCY7dyIADiZqu5B4jMRqUYNhZOzEbBBOjScuZqvI1ChbjOB23z6+KT1z47yp
PxFEG4TIrvXvx2jOJg/yyxyEF6m04hcOw7Nu4/5fzC6xZEHdFONRVEQM7ldk5a34MV623wi16CWw
VBYmqfDjiNoHvSk82DHwW2hxMXBzaa1PI8t+FabWq21tF1LkbNJN2aW/CLxhe3LLV1u9iQ49RNtf
Ppkun/lXvI4N59a6JpWkqxkQihmeq5vl9wQeOIsHIZaDTZkWiY+3Xtdo6oNWPVQm2qm51ByHW//h
TT0hAO7pNeL5etKRy70e7PCnRzm373++jMhI/JgVSVa23c4HcsBon/4xyTbdzHORRy8Ye7jfYKjl
Xhyl5/ey2KF0PBMhffJeW2sjGzChWYaBz6GDWsYGHpsdYvg6C+yqMPa3KZp03m9cvbweqhlk4c5m
IwdkH/VkBj5YzzX4Y4yuC+9S1SM3YNjZzVYNQLG2Z75RVLllWmY9BN7XBt8Jki9CGT319mhJHYYQ
ZlTrTK7Gxu0/ubTl1Shs2fKPIF3yTCkW+2VOc0ffAJXNFsmtUEY1ShX9DRcBrBjYiY9noYX73blr
9jHOQTD15zrgT7nJZ0jen8IkFbz0rHzWsPcBBEjD73llopzRPnRhWbV1HcpYyytE9ar9ihQvdOKH
AaJoEH5Lbw2OxPNOwyLV5mviB4Mq1bM53B6kyEI8ISPy/2pe80FgPRZmwZ+U5Mua1ipQer8MuEXw
kWvyIPcCPBJ1OLwOkUcJpOUzgZjZ+JtIZ4kpGxiQpFRDcaHinwHE/iLvnTDAVIguLGcVZoitHmKw
n4MD6hWc56HJgPxoDzJLocAhr4pJ2BzabbvJksaD0xyuXRBDnppQvzpkw/dTc6DLeyEytpgj7kji
gqh09OG+IhS6Ww4lRl6od23gwWKvOxaqcQKjfTWwKuMooxQZGXgMexGD/YUJYKWEzfsmDfUfPdYK
nHRcaiF1wZb08NofbRh1hHo1sSZCYq5AuZrVT6eIkOl0cNKMu8ldvHlrV/26DpQg3PqVncVXDah/
DkfKM4+F11iok4TaufFXMt0QQhZ+HkddCpzkY6LdqCTqBmc4UJGoGuGzDvkAsoRkv5sxhBaWQUoX
v30ivLRVHaye1U5az6nTE3eLOsQHoQz7N+Sb6J2wAPo0FUKHtV8tuI7t+lrOkljSQTrQkk2i6Y+i
Jw7GvIAao1DrrB7q0zvHb/R+hlu+UWKt4y3nHX0Dtuzmd3FMyO7efrv18k0LGhHU+9yJCTrdmAtP
8ZiNaAIeICBLNnqxYRAO/hiGLT5DJztGESaKzBhnFL8T880Og43FdWjBZJQ4RpPm6azAYYWyWhJ1
49iWn0HRJJmFbHfoIKaZ/zEVOAJbl6UaIzH0+T4NYRFCe2VFsxzyuw8wx80bWSgATGyTCxMxnPRo
JMDITBWsLHElNaqaMk1kzIeMZIo5ERpkwg3lBdseQKesynuGKkri9GxIC1B0NiYPN+eh1cuo/B0v
CgTCdn4DKjXNKyISj1txFo3Jn0EuygF1SnaZBRBs99TXrKvngUtHb2uEq9GGFd2q54lzJuczVoRC
0VujWfmMn1AfXljY3ZCBHJLsQkN0xK7HOiXzhpTB5nB88fRtARzVa6PTUz7VI7vLf8DOavzD1qGx
zhPqghHKWvhy2+H3GFfm9NV+ro/XMNEdfJF+SMdzgbJifQoQ4SM/+VloQnKfKZHhIOzzRo77k2O5
DqniHnfT/DTFVwgrMd6yTzcIH4w5B8fHFP8uMqkOC70kovnyB+2lZucSY1FVFg9Q0r0X/ojW2wXz
Y5/DhPriL4DI5fcSW1Gpd5lCsbYgd/wT+K8iUgY+QLFHZEswTN0p2LyBy4ur4K4qizIorp51lAcD
eLZQL8vARrvhbp/+m+s8DuaxvG9+15RY4/1otu98to8gqgyP0suT1huqtkxNVHPmL+J+wJVpBpaD
n6WeMuBDccA5fuVX3gYtfOfGVgV6TbCQC+ORmhEyy9DEktMH9m4rKHyIcSvuvWu3RR0JnPDb5whl
hmZDNOylh3oXLW0KcqCIXGIQTQ1YPtU3NSQ+2NuCmJdxf0i/GC6bsWpcOEfD6bFswnBqjCQ5p8ea
UKZIYioiZbFB+FZxIYm+MdENpzWcPVtWSdqwwVJnOrhcAtq9cSXiSepUMSPf2dGJVIoPyksVru0G
YIxSOlHz+23BiI1MWeaiiH7G5C97z9BQTHLYcYZcPIrgyTgeJRFUzYPAeZMt1klwUjLkVAb3ojIc
tjZNVr7reVQyJIlrtIjbVV3PaB//QLo25oyYF2F7yA2U0W4oKvmhbUu/wldCyGVKUdo9buDFMbJV
xhQej6a+dZ0PTBXIoVNLjURHgdCHdTmO5xirMepu9jmHh3E/CqUL4riISQDg94m0XeC7v9qfd9mF
AQkJIiJCSqjf/KXQ6vtVMnJaMdJlcMtWjQFhffpnng7FeC5XbUXSnDB/VAiR710HAI594Zh/9f6B
kHtHKmVmyyNzJonpsRhOgYsKYHtTGQTQrEWIyYQZkdAgVRWxots35SYREaEA1oeFa5lmoZFVTWZH
ur8WndTI1c1RnA92J/tV4fe0XEBzjoxE83Ekm6AySeGIREeOz/IjNb+cBnhp5/dy5OhD0fraoEqj
fjwrcyQafrQn/UAhREy31RQa0U4F+KM5yS5/Cbj7wKYR0axjrdqY3F3sGoktE1mXUZSzOVbdF7Cu
1hgFKtJvClHrONHl3aN/fnBgi0ZiJirX4XeAxVfyC0YtOUZWlXwaqsWw0BSO8kn4zP6dAp4wIKKy
kcDuQ6lmuNw2izImA1rPivKY7cpcZAiFcb0SFjeqM4RhHUtmOILuzZLmKBg3e8lLexVLTb4ugaRm
nRxjhd94peP8vA9hhjgItvLNwlRDUIpOm3ND97foNqzJOZde3gT8EBlmjq8LEPadAA6ARpRiCXY2
s2ia22lph5BdR4RzGNP+5KXsEFugS2vygVOx8kJbj/xhJJ1NX/er0YVP64Q9f2YwBTSZc7RMfniY
GC84kh32d6JcE0612IYLld/uCz/UD1I1HNCKPor8F2t8ax1NtLf6q7GDGzmfORhjlN7Zs5/FEhAQ
t4vCFJ1VtFvp37a920WxOY7YV67YYHqBadsDnwPS6dDibe+TeGRAr3ChZ1Ds5Ih/Vb4oxaeURVY9
UfCw/MX4Mxb/WFiHcmA5c8+WmYyw4yKeqVeGHgq/dhd91GWMRw66To0Sxkwxs9DoWX6qLQUD2MF9
/v/nJdm11RDI2NB9A1v9G5UoOv1j2I5SRtldgMKvBBK2OLWb9HlTgRkCkiw3uK173CA97a3q9b4W
AK6A/dPV21gu1/w6WTvBJvZ10v6doSnJYFOvenKQQIJetNA/+2aKm0CniUHV/M142e5v9hAhxbPO
FUsJw0DI6Ipg6pCfjJdsFwjnYgMjVilr2WFBMjgKvdO7njnKZYe0+cXNWghM1qEOPdbXFOvJrovl
O0b/pzOGQUuIjMvpJ+xzkSyXpSExiwWWhUo5Gc3kSJa88Xqda6QloQaicdhOMfbZmlbH2lJBBegR
Y5mAoOwiUGVlSkfUEyM7JWDgBrzVOhGWKnARfaDOA1LgTTxtAQFQlM3WNL3GQ9qwLV8PR4FWSWRK
5Qo0ur32eGYwDD6GW4t7zQCKFVa5YPRkCOYTgBddmQCYoO2dFzWFO9LWLp9dUcXOmn+sY2YLjLuP
j1hDmPzQZzA4YAqOIYweNG+QZo+VKY6M3p4VxT3yZY+Oohx7NdGj1gfC3oCbtOUk9A/GwB6hJxxc
gd/wdaj/RSXc/R3+UM0BGdgY16qo5RpVIzuYs/ArUwbkOZU1o5LJAjrGm7bUgrkXVJgS5jdv9Qan
B0PJB830U/J3N3rRWyEpUuL4iHUY0GPWg+ftyZC4bticC3gdpr56eoi8QKBZmNftw1voI5ouAvju
H5XM4wpox5oEoBEqUEPaWfTV62jOair4rQWF3SkuTQb9bRFAcc3yLifh/mGGVLtGFgQHezuD7URl
D8Yzg9QHIzEkUShT0/nhB7zxckSMr/KXpN7kGbfeOvbkgAuLr8LoWfKkqvUNJCNcwhgWZEJkQSj9
JvU9uWIdZTN695XcrMcEmQiovAZ3QdFDnIeg7YUrd0bJYfzvFkr206Z8R1jlo46GBPN7hNNW7McY
L95fjDs9VEgTJAwxoQvpfr2DCINwwd9DUaZKQ0hpeuu33LlZ05Y9MHJIM+HumLvGH+fF9iu1j9JQ
GKfDc/+HFY4TRq7y2icp52e5VAx8cO1y0IpMW28ed/Y4JjqlAMfA1BqO6mSLE/wDLpERO7JM/aey
KVV3BLhZkkmNFHwGsSEC5JB0Cg3Ye+eSRTNlDPNShwO3quhjiI2JJCYm71yFf36MTrSnS6hh2mpn
YQaqIIBi8rXP35ocijNVYc5elKOVSUv3kB/SpXZnF+kcaHaMEG8uSU0MtF0gOpb8gRCs3UKoBdvP
LGIiwcyf1Wi1wNAWMvJksg7osCQP2FYRJlJ4AqQmKByT8Ps4IXYp7Vi5PQCFyPrKE9lLltonZoKv
Z7UP0vxGvgrLnxGaEbtRdVsMybYAfMGERK0xPLp0ZM6kozpQb/CDEsVQZwGEhSfYk16dRpaDHVL/
Ey5rGlS02WhufRrErW5XI9AlkSKnGEOGf8BOLuiqChSXUl0ndsCwafDyHXP0OqKZ0C8h9SJirjKW
SgIRYG7d7bc16NleX3loSMnZtkeQBBmhLUtz0ec/UHQmV1qDxZq8sJawAvIkMgg88QkBAYGb526r
OvS+R/iZrpvJM88D02G59YMVrrTRfB7iDQ9Y8CeKw7T5En+2Uj6JXl0onf7qOXWFjm1JwnAnjyeU
FXtCm2eXORRzOGLy6LqxQ3t+wkeXe7dJ3JZzS72MwbFoVUYB/+6m7Y6r8ClnNf8Dr6/tY6+uTRT7
vGymVSpmsnGfN/IXBm90DG1i646hixx3BES2j+WkdEl75y02NhYZY6UUTTj8k7uHa8Cfug/sAY4D
6JLMfmCyW5h/d6RoeS3Qy40Q/CHXlAWQgc+PsPeGTLHfbKrPZx9ppTh6SQ3b9rptEObM+QWis1Vb
H5oCXug5lM+tNk7ym3ybaJ7khgDhIxmGwR1SyXgCY/5v9ZhqapUBXkm8Rwneihec7bza2Q/m2CjA
4rp+2j/mm3M+YhC0+X5mS77DmXaxcmMxVHoOnwsyDOu8534Y8zbO0y94cxOX9RCwtGfKVoDARDzq
LR4aWxWWo+yas3sESSBJgYIczGMtQE8aKao3lkNokNM+kIXx6N0XX+iamCNnshYztxGlgsKFmq5j
xNUyGj4WsuiPrEeUyfp2jtD1M7hTw4BWTBc1VuxYVR0T6G+0B7zQIRCDfVzsnfoQAzd7lo9BmfH0
+RYIBPO/cjmMV70H8T10AhH0BjKJ8U5KVci8Yzx2+555x/mRmZnRjvSfA8t9Q6n/8uS+P54AMTLe
viJiIyMMa/OdZxf0xmAa63s4gsFQaengg/ui1RACIEowGZ/5SaeuFlCwa+9kBcWyWz5gkOxNxD4I
HIoXuKejVHeLiWkF4stxikmMKKkGHcA6ttlVe3P26/DQHud+aWLxUQNsNRwZrLhjrKaxgpFidm3A
aOodUJ4TUNOkAI6Ry2+ZOcGrgwqvvIIR35QoSXDF8yP6TBuBkhtlXf8rFfDmU8ZAsfzB+bzGMR/3
yqvwCu4Yt6FL1QlsyAKfCHJA5lT5TOgfcY5C0rzdA83tmLwk0ADbgID+W0pPaHsPFZaOBxNPLJ2S
aAreIy5cyYpoykzLY1tbfG4RkIXcF8TItCAxtCNb+dAaW7wNa8qcO22exciI4KvWVh6RDI7jD+3W
pZme/sazmrEGUMJzBXfbLkPNtXZvCh+bJjiFXHdsEHdHSZ44zs81GLPes9iPBpxLmRIvRVVbml/l
+nkGKD7s9WAJfYneM8dqZ4Fl3OwPuiIT/n+nRwSTMLpt65YdyzVoEhiFTVniTewjmTr2HTZ5w3Gz
i71v3go9tqQoAdrhfE0XbzjraAOpXeac8Sxjha1hIoxa1n82aCS9Y5M69LWoIaLVZN0zL7loDh/E
iPFbs25RRGd4NwYjP26esGsC0k4u0LaYg6AFjo7i8OHIHuk51aMlIDNz8cf+MCjMxjF4Lskcclel
F8MAfVOk4Ce5/bqYM5Dr/lEA4jAXXzgspAHsyjM19m5I4xpOz5XT5r3sry7Shp/XY7OWsBq7Lofd
uVD8b5Af2SC6CFAq67HsFteKwzANzAyMy/tL2Xs01pBcmqGTnnoseYilh1CxxGIi88xCz/wK+CUu
uMmZvuWtvuDIqkwitYl206RdmS5PZO8ZVG6nZ5CCB927G6FsFxgCAA5UspNNwudOR8GkDSEJvbw5
qmwOez68V6BPVnNbesHE8Xt3oiAHo6K44QfKIT1BTlt6QQSgLY80xvIPFmdRGxo3uXWST4DKSOD9
jj/lEtS/RqQCM65QNGLTkuTr0dqGDAkFIG33FjLp086ubE1U0sbNj2I97DpfippJx53CUeQ7E98o
6/wD9bbn1yXuBpfADEFWhsp0fZfYOUclt2E6015TPpV6a2yO4Ka1RLVhFe7tSe+gGmuKqeQQS+Q2
vnxI7+7zd0w5FGpCKNlGhHhHbGSHIvpvovy/jcc9mSLMTXaf7NfvNandwtXn7S7KX499TdmUvbYe
3awT8zkfxhLAoAjniQ5IzudI++bKMkJ312iL9669qU58L7/2pKzkClYHEfpzVIUazV4VnYnvoAMk
TiJiEVU5EzROhEQoklzM7q/rlJInywgwNOuhFEZKKr3JyrqZyMYVdDyChVupH80l9HMMbaXBMRHn
MQFlHzuFVRWs0eZ0R7l3SBXAq4y9F4jjfCeTZh96dBOcSmNrFZt9OOspvoBIVmMJjP2om6nyVNU6
0wukLx2IzJyE5LymPD0nM/rE1cIC7gk3ZKcJaB3jCSuAKr5ul1aDLDgULFe0d//L+ggKoYEh0dl+
djlZ17OjISwbOq8M4a2qDGOXS1Ph9ycYmu7SU8oEAxJMkIG/JtvmAHHdHeF0G6f2dFmlsTqa3BFH
nZfhIiV61VXbBndtdAuAMGC/xR2DDMPBRcG1krG1L3YED68po22htmw51YLduJPrrQpbvzkrKwP3
BuqrKEvpseWoEKFP/3PB+N6DQVhTooEVX9DeIRft0654jzIO0zgayaHGK1LZy7nTQj5tU8NB0mbR
l8EQuvDnQuHl8GxF1C6WSvWoywWF495eRNG3mZWebSuGM6laW8VzrnACpR/KfOe8J4Wkw3GI4mWm
GHZfN2/2w9PI028px2tu8vLhkFegpynBXJpvPm5IdDJH4w7T5u3lozH1T+hk+mAfjGH0fx1hwNcA
ln3xPdrduI095dFiX7HKCFbCxuxiXTtenwVSkvaEGwrcwflgdOlsc0/Pa2RGwDki/hlxDqRljns2
4aLQmnTkIWf8PVH4G92NqXDeT2BnDnWRkuQ9GI7IwlZZQ8odDv933aJrszHPV+S/7zlws5COqZcz
Son1tOt7Bk+kL3EneeWLvvuqnSnO6v18a9VQUXDw4l68uNUIi+Px2PaepOJym/y4y44UU3uRW7Ke
X9KvFXdhdo9JPKhFy0Dei7/l3Yw4Gef2vpSVnoM3UzzrJ2ab36PM7+Ho8z5cY+gjogowQ3Mple4B
h5O2mxNfcCeH43wlwoPVzu8xqbIh5QgdRAgNfFFckMEhEtBNHY3vPJRboCSa10MDCZeOK6glqE+j
7ZCOcRSIw2MtQFVADwJA/lByPtAIp+4Y86ThziMn0UCTXVjvfUE6LoZJ9BZCM9Gr+So1KcXr3HlS
pj0ZuOGGQ37oDKq6yqECw1fSQuajyUpCP/UnkrMlhR9VcnIUNJsSAbESY3hoijMN6WwnJrVLWukA
FyeyVb03Zztn7rJOyDgrr4og4YUQF3mhYtTD5MyrDxO2+1u1ztOY4dAS3tiFtJ7gCGkNxJvNAVnG
X9Z3ClOE8ZbGgqhIYuB6NL4QYKU4cp5vd6SM4C533adFMQ22GbjNueBhffeihM/oVMYcPPIXUIJj
mDIpKZtPQv5t0YCLtqCfW8z5OUcUnFsyg6d9Q9WxL4V1moMfADKvBx1JnmirBa9lTac5ONl0sdQS
Qj5RTE+1sdqTjogCg3h2bHQBAfizdWlxmZFd1lTHoi75EI2At+1OgvFl0mXyo9Bl2+9t1nWVW18I
LlSLLpLtx2v6dzRbUmJ9z/84k37WMhQ7ntathbRWOB9M0r2u6lWRqijJ7IUS9oMVyjLVk0xbCCs2
FCsV+95Ay+ethTEW4sN4JG6KxX5hOd7F76wf6lM/kFNT9owv4f2Z5M6TgwWaK/v8NUD2B1AozdUx
rWkWpkLUOgs+SoVsWyjjaZIgzjc+0yceCoJko16bsCcg3Rp9EWt49gXR+43LMj7ZZ9YndFagweaW
jrwKwv+Z0d4Zgp4LyLjZFiVkKgnEkF5vniPd2ahvze/PdNKgtfIXc/kvvAA6nWrRI6mrYnoQKECU
lVfA2HkDTxutsesV9aWark29wR/JDt4PQ1x+JY8QyUnA3eBNrY2mODTas2Uq0ehQsjMyrwCdMta6
iVUo6ELBO8R167BT8bpmCarKKuUwlq/hl7euYkifpKdVFgNMP/RQBV603HHBf78gN52jzEXgxaqL
BMt+KdJQMdm2QxzbMqf+A5bf0Qy236tiv5GXui04WMeK2gF3Z7gMC/kwZ00gGxgFgvxinFpKjyhE
U486+tgMHBoT9ew/fq9GOo0wWMmLijt7nFnYOtZUAEaIgsy+JP2reH7dCgz/gz/doK6RZ6aaYAWb
wWPMNs6JftuyHwMp0Y5WHUUuFYmC4QlLReTbBy40fYLqgAvIKLPHPdDGWhvdeAl0k8uiKU02l+oW
WqfUVRbRHgNwrjXX1jqEXYGZgBv9vnBZGl52HtZCW7pMzLUaD2+src620oplMrE4fmpapwR9swT2
6GlElWzU41snAXGCjvh1g8wlYO9fAiLfNkbANka73Zi3y1qV1bZ5DUzpvPkCCVW2qzwaWMsDWXM1
cFwkxbHDkCaC93DkltH2mOD3NWLDNRMyV6k38lznINIFybq7cUWPudcGsQub1M99xbbAav1zKQ2a
OZqnd3ljwhuBCPs7wf20Ao2fkKQVdc+e1JNOQTLZjrdBK7ArVSfeRoePvdoIYy/ozgCs3I6PXABQ
EaErO7jmy+aQOPNv05eFwjy64G416o0AWdJwk/49YdxDdu1ALwvmwYjTD8Br8eNMmHxy9lY8YXL8
0AqqTVrwJIdN+di7xYSbU0m2M/sO4zoyT7lKJJA+lz7RshXb77kH+NG8tzdpmQ18IpE6zQCJi/LG
VYtIIdA1n1VDOw1W7S2UwP9hNzth4ECL0xxRRzXT+uwCmDXivdL9JSy63ANg5C0uxapIowCJptmh
2kxFgYfVULyfL4ujXPwtD6rmWyvOejPjv6YNYrqCeVeuA8+ZotoO4dI7K9FUpWFhOH7ZLKuB/fnk
+VJBeZhHYR1xY/CFHHxWBrAL9cVAf9IhTvhtBsEHESKcDtUDwOI38niJ0B7/2HKsOl8GkwF1JRRG
KojRmXtodPD1g3OA2vIIlOB5FR2AmzPDKauQGSzlSRfR9+yP+IcM8RFMwcx5AEmCOyA985IF1P+Z
ASGeEmfZbgEdwgjQLMbRGQiyAIOvVdxsC1Gi/ckyo+y/vQqekXGryU8dcVwB+2YKWcp/obvfC3r6
p8e9kl3FFKJJKPhN8cKnKdwJcVRelekNoj+dheygfA7axHjkJ6iBWex2lK2xRJJqdMSuXYYZuHfX
6RuJ+0XVn7pZwLp1ApsQifvTZC8s4wga72ac6YjifdlH6BlYA39GvSGhZ0IxLKSkgLIUD0dVEvpL
3Xa9/tEvK7idfsJKuAq+YKcZYXUppL+5V5o8tlC78eOUpoWmw+u+tYkruPIeydQrsbPIAJd8IMJf
p+iEuqjA+JLdeeN4dfTjpwsyHAGHXk8f0r9tAxcqocDVcEDhQ1N0LbclDV6PoqnvOVNVyQt5lwVa
p1HMuEhK7g1kr2mbJXKww1EO5qPCYuTxZzgQPMQz0+AFV1u1iESeTO9TkBOus2Qd5bIZ9aQxgEW3
8UHKU0DpaTZUnfiBfy46wxpI9RKYBu/4GzLairsZRydYfMqf/aea+tkLtdhqmkMYTEXMqNJWXbos
uccKLAsC1C05fZPMoK3aJhcuK6lq6bql1QnWcpKvBe7QBIlhXn3iGtjJLPaevnjrHCeSi6XVgr5k
7sLffly3Y2baW097j9Mikn6wv2q83dmdNaH0mRy5Pw6iEEWh/0j6vc190UDEBsIQPic4lt4LRzIE
yXyJp80K82LSf1wAQ7Ld3C/4gf4B5/oH9slodVLgvuJDyxg9NwLGBDupp1le1cLzIj8ZI7R3pk7L
GqXzM+tAGDeSIi7ye9/S9ojWBxUnBVBrxKGZ9RX8PK4inMZQOWohEoaF89OPqwzG/RDnQHZO8G6T
PBD3E/5UimQX1KFX4xHg5i/tHoXh0Gh5RD4ywyIm37xavrg4osN9fqUt7lpQoMM4UzAuEuQ201VC
OYiZMkAgmO35j3Ue/PirlGhkycWFm/1UFNVbN3tVp18rmem3lWwGHqrDmEOPeSJpWOgQebVV3xe8
QPuKQk1MFvi9c5yBmgNxU0Gz99pRhl7dU4Jyu5wx/DfE4KwEKrqDjy1raGQjjw9yfQt3tOGh2JuZ
enJghG19G7FPenH4HF7DkiuC0vWAQ1idN+txEHSqBAxP4W8ec+t+OBcQToWU0Q+1CqL4aBQBZQC/
yMXCirAbpSPonlN6UfD7cXFysGUDLKjl4aa34gFHVUDg3bPG6KMvLTsYS2MZV156ybxbRaycSiMq
50baZLrz6JEMv+baslyhzCUdx6XZAPnoZ32/JXZp67YzK2Yvx+GCi2epwxtUHjnbQByQqu4/cEUQ
9ojqZyjqDyNoivgQmy8dUqqYaVFwO+XOKGmsdBuz5XUj/ShSwsP0odYrj80zItlNtT61z2fq62pn
DOgF5uVuz2Bu4igs80WnXDIVTuj87O6VWJ2b7GCGv5tmQzEO81tNneZ+cNQZVOi2KSnCDVyBOSQa
3HAR99vMHfNctVix8HBBf/s1LF3H2pPrwK6FWyiUD2pAR7BOXcXTAo7jj4XjJskM608z5V34zU4i
xTk2IRVtXn99TAz+F8Dj35OYI/u7ZCmULXSLK1kgDN2/FqV8JB3jutPfajr2bf6OgBh26HlT34yJ
TYL5rTXIYNGV2nINB3KBpffOeLWOpW9GqsTjQaOcboRT9keHRrUkpHET4xeANkqATom6OkqNBTVS
wyZuQ1A43Pcof9EbzqacSLh/ZzTigFR20LQHpTkD96mR4THmoSm/z1aX8tASCljhd3zQj/CW7aqv
6pRqnMAUbXmh1GP75ZLekG36Xp10DAuht7/tDU5J52tB5Ye5aQEpbrzhHsDl2oYVH7k3MmXOKgVS
q9Yb9tIgHptqlcGjzmcRrydtsBzq/49TekO2XA7V1wbYPy1Ixn0rKBehn92ilXBLG2jhtst6Z9IL
1RPY9N+qmWtlJcHLyFYipi2lQnvHOMNVospIqtEjFNbIT0e85Z9LkVfcfZrz7j0t8Ceb1Es9BRXn
s2lupLhN7ZBP36g6GY3TBvp5DaOaGOVnMOUSiLcb4Sop2I2tkt8pANTYePXhqK/toAKGdtaBWnVa
dPP3YmCgRDrV8OFX/Q1qgz/JMomObAHbKSF/dmlWo1geVA5qU6NeB37SU27oUmBovPSJSi5KkcM0
BgXWEezEEhLTgCvtpED2G/XWhH1JKDPd9d/bYTJxGW/kUUmCMUXxDOtQi0+s3dQ7cVzboRYSV4r7
I5WlsEwCD8xCeQ8XfD5thosS6bFOJpeb+bJldlZpu4ALmLJxO8kpI4KvWceG5V1yKtKtumBWIXDe
7YqNqxWKJiJ/+YR7SZ6fE73b4niEURwaoBLo1XtDKsHDx/XwIpBWCb11sUZKdwSG7G9o5AFw4rx7
qPE+Cls32K8vb0XLgZeuVEqv0ilRmHUcjk4VEqWNlYsfejYkVZgovp1/vf4M7hq7VzH/m9ITsoeK
lb4mxNNBWVuewHhh3ekYAxPeWVbZlgjROABJkXbTrUdpwGZmtlJUX5vRpWcMtUi+Iir3vh4yO5M9
kD4wbjCUMzZnzxQBhAC1yIemDbwhvgm3E3s13Kbgh3whGyXzLBJmdBHb0dW/M8WkktOXaQUYMxzu
Ye9M4JJkmHVlU5vejtc3Ez4geQaaVUPcMVIU4AoMH7li10RLZscAvrfTs2rMXVdM5s1JOMlJERt9
0NxuKYxh7hhhfyGH7XYkJYcOgmIu3+/h289LoTBRW7RWmTD9go5TGl0qcxyFZqB0wSPRfh2pS3oX
qBLVDGEnu9P+9ER92EA/KJC8Y6kJ1KqwRUgLgE/VL1dJcO5S0j3NpEQlADukHu+lleE3k3oKDaSh
ZRozqp6lwGrjHlb5ui/5958cBfafnvse1Qp8P44MEYnk5RDQhFuQR13u/EBxLtr6Gz07IdaJzdyY
5olv9qGLx/gw3n4Kk6vZWTSblXZHU+TAoal/L8HKdFTs3IMxTlszOSsQ+8QE5MXY4z5NTn+JVk58
b2M2ADCovv+iXP7NzjgHSHG/1rKHxQh3aj9rFBe3TWhVoJZETP7ZOUY6XTeB0HAjEmeJUnAsFajf
1TXI6uxJQtlduoPexPJVMTq4RrXA26G9huoIZqMptnhcuK+NdEM6ojavbID4Kg1X5ASLsaQx/BBF
G49lJa4QnJG62IO6s4nuhYPUBurEpZKjWU2VWG1gWXcKhKct4XsEYOBXKe8kZb7YzS/VA2WFX6k3
4VsZ8mocAqykaaYYh2JFrOLEoOGOSQHiCHU8K9nnoAoaodzi2Z8u59XnK/Pj6cEKbjiPzHlSh0Un
V1Gat6ms/1pbQXY3MTWDn5FVWlH5Pb09RxmsCXt7U99ORU9w0TqUM2O+ttlWs+NG8X3j19h+l09B
6T9XAGGWPk6csEiPpAgNBEsywTQFZXeCktyvyEuyrWq2kHTr5XkT7bnX3y0WclVPmc/Ne3LIGTK0
Xe1megV8OY66WgtqhSIjekY///VbaBEwcZUbXe6GJ9BrGCKDmLFiL0e1WWl4LgS9VZJhd1GeHb6m
QdnDzDYZYYXfOgOatoIB88ZwVHDWASwTO5lpvfKE5QVM5IoybjPH39TJuggU9hNl7kGVGohCLi91
w15jKi2yEcKDBVe+lGE8uoG7O9oD+F+JXYiLxn+Piykoep6Uvuu9UPMI2nULGNKEo0a83ag4BxuO
9XuACMsD32m3ZOGhhS8cDbrXVAB9D8bG204ijq2/98ch7fUvE2tNTX45vuyzUKodJH/eQd4HAAXL
62TRqsMHH4z+dR8pBSYcxBd6gaDtEZTGc/a8DN+Yo7qNSapv58THnvTbjIUb/J/OL5M89BsRg4oi
nWUSug6xxb+CPzt9Ja6J6buetsf+MO2pz47RIkJqCGYtVHOsigqdHKIZ6QyEnXvI4Tshd82dDhaR
yxbCY1WPPH8Nj0bxLxlc5R1TcuhFQ6hTpzsqwu/wOoBQxigYyhWy2gwmlLP6hscMyToVTbvpwk5C
qRm0D+TR+TQa49W6YJpKHLLwP/bAVvjlp26EEe8BwWyyunCR2+enjsYCkEBfkmLnzS2sx9hzkF+n
3rVM+Gy2AU8sevyLNRyXgR3/VntnnmD3azrm7nWPjbc60BwvprMbgFI6mZ1MiW1S6pVFcf8VUXZt
4eKqrEhuYQugxytRps0DNKLYQojKXq8pCfU9pe+TiYRv2W2ZoUeSVMhAMwiprlzARr7nW3doL4qD
UCS9Ak0itEAxrzhMBDGWXut6vtE6OP62cuYATT7ySkd0GjpanSGf6uNoVLx5iXKWbMWNmmCxLJVB
9/CYNbxU0mQ/mJ+MpqSF35OScfHhsJQcf1t+Fs+bBrk1vSKApzFThX7f7MIJJrVnPR++fzOjG5Y5
xmSkNau7Y5XVm2yO4/gCyb/JS1RjbZpMSvit8EuBgQEqREri9ULhrWsldA7XivyWlEsK3RUZL7aQ
OkEmQC5zUk8+y45F4F6/2M7sALFmeRQuwr5GQKTGFikaM6dp6NIevswdSQCVAJhCFPM3tBUXwEJx
+e20uubpQ0Dxx/GY/rgCEjI5wU/fop45QoMceBqq9aDGR62azTA6JYZTRAlw1ADlZZlEDP9J42Cd
f9gDAfC8JAqzoLI2a8I7eN+aJ9bKahYAdFG9sL+JIHfiJmGWhR+/SEggQJGGpyCEUvjA8XmRgmJG
2PCkG2a/kBimm9l87wV0/GodESoZzTpCDyAeW+25f2dEJMoy/b4quuQUbdgD4tpIxZsTaQN0lopg
EO3Mv1lZ162TMt2F1NbIaB4IcVSKK5libILF1ng0DnjbYtko3XmywoteTqe6tBWgOrypw9XACrSs
nVA8waAMpmaZ1QQsEjWu0JlLiRKsNyLt0djQDRQsztg2EozEIo8WQKy6+/naV8RMeJz3PY8NAlcC
h32y7+CWwec524gWTvqblXfirytiAdIl0533SeSuBAvlLKRWuUygJxkVcyCeR7BwMsv/wHuoppHb
x/H3j3weQWMMRVQHkEiZ1SzbkPUFTGCOasrkvPsVMjJ/xFvtUVLlBD6Fo9dpaaY5bPlXxkkjRpDp
AcU0zOm5ZjaXyhzzbS/IWGJMs85XdKcJ5gz7bdxBgelE6lEIo5zMWBSjSNEY3bNd+Rbe9m4q6Oxo
Za7zKIijbjdE0lyGdbmki2lXsyYtFu7Krkw23pjYZOQL+OYApZfan6Z5BxvZGwOkqL17yD/2Z/eY
hcs+adyeuvMbVo7jnTZRevzU83+S7Yr6gZwFgSTi3Yn/zALSkCAJ0HZfOw/42gIR8r2RaKyXocp/
DAM44yUSEQ6KxTa+NMENsCOzevNK/aUFimmVzJpTCDvX8WvPirSnEHakE03qw7nXLFCuWZ2qCWIc
eMmRlJfxLZePFSKKOdrcayNg5zIPZtn3Y/Q2wTvD4599AgLX85s2i4BDhZuparaC6TT9Tcx3Ry7p
R2DZeeuvHbysrUcEH3nvLRvIkwmETZoSnDyn5PBRU4L28jzT/OgU3VgFQ2jcfwA2sj5tFlnHwn7m
27xCX3fyK9QKbbhjNwtipfQEwC63wR9xsE3aytyntX+IpcKwlTjipxJehfGHMPy8iW031gsByHcD
0fEsEAAU+G/hXFYT/7AngRtbeUIzwvEmWeMnSYOZbuCJLbiCxr2QIHiIW5LWOtqV4Rp3uP+e4DFG
TRhN3ML1HSh6e1eZv6XzHK3OByLtIPyq5Q2aQSyf8w+pPuNrXl356BphOQvM7XdiNAkBx1dvBoc7
J4S4lJ5q9VMxTkKilc+tkRjn2htFCV5WbjZs66mnow641dMfwW4xJxuFd9VqzichBdYlBeJriFe6
J1WAWrB83d6qoLN3w5kMHwmv3aKNXyxQ9g2+SsPQiPLVo8q1wktIeVGHl1zLurR3qepOjg8uR1Jx
HJty/tKGZX063d5pKkjxk01CkL4ptihc6OHzBhJ4wbNqQJC0c/vnl6+KohUew/jT5FoZ6X6Ozn2h
9UcLglgC404DPNkiKEhaLDiSNiQ+20dh26h8RjXIkH8XiVxwIaC6kMVZiW+T5NQuszYYR7IhUE8L
L42ws/k5ILtfItKk8OAr99S0Z340JRBxhJ3Y6rwnDnwZ7R8Ad8bExdRB8cPWLw+tTP0fSVOkeOcp
bUu9oky50RKJOe24/lWL+05dl1aHGRTELyszfsJz5RvtY5JGgoJxta+hP6XoMlT5HDnrdlwS9ntC
IQICRHN8YAUX9ehSEYG1+kkxNgRiXyDziCeto6UEMwKLDiBx6w2ZNO2h7MTNTl9mCV2pXNnh8oDl
GNgtzg8Cv9/NHst/1ReAIwezPBjQkzceZBRT6aV9V5QV1HliICRLyiayfDEY59oiluZabRF63YbO
mdmdnN8I1o7IBtJOQ30vdPrVPcNO2SnlFr98EPVG4ULDGbNxDmXTrsR77n+KBnQvCV3kH5jtP11K
FAOCtFM3kNvnGdVsm4U7L9uLxnqOqixv0UXRn4Ki+/BOgPXdhhRYx62NQbSo1HbKopW/NVxD6beW
6W5qgJdQ54WWZnro4U1XfxQ3VZTDQeG4xcDDVQqSbjIj+Jdm5UcVHRXHrTtDMldUDjBx1qtKz2m5
pZsIM56hJ27GPTJrEWAv6rQc+OTu3UtVRA5MrOxvdGxLfnHj9o25bj+8vQf36bM1AcHGm51+CXUq
NSxRS2epkw6LI9uP5z9conWP/oxRRpwZQhKilX2wA/vxVbW06mKaIc0KgXsgwCmtjxiTz7JtdcqE
XoTSt79ueDcqHY2In0goZ63A/7rgFDs15T1JxfUQ1K5c4+24o3Nl8ScF8WZBU+A1B4sBNjCG9qK0
9YxIvuu6cDUxGyOLm+K3TlfvuUGD6x6LaLFDh1/b9Xd9XHEQILb9rd09rVVcmPMxo7sVPBdpeb7x
EtAStzDIncAWFYHmN5pfKNhAHXzFf1V6M2gWL923HsxI/yCNvOKvkW3D39E1+2GQKhjVeGr3uqJV
f9ZJRnkzMSkwK3iehnCnYuXecRiJQgyQ04yW0Y3WwL8oJZUXnjlABVt8vsVjkkY61ia9Fn7peKMe
ZsiSbvj91D/+K2doFHBf9KE0OCVQnuLhdsKhNk2x2ciFuhEjCjKlMgBZb0fqa2GGCpXhzKGNTYte
imsaAYBORMxSXuSwSEXcwBKqhZrt+nqB/06giWC6Dn3X0NcZqwEGFZ5waZGlzQqv42DVuxnPS9Ac
vkgSDoe1ZDPl/dfGKEUyCn1IXUL4zRqOhrqFFBQFPq1u0/rWiletxaSrDB65PYZ1qt9UKHvBZm5H
M6rAslcvHjQ3TEqMO7BnnGCjrJ7V/pSQO6zk1lLHEMshtoX0r0zY9MuepK8RKSUsDXzdwufc5sO2
OfKLqb46A3iehj0r3XrBi/E7XRzeE3OT1PN5fgI476CCz53Q0b5ffyoS8fnrn8nCmm+S6UY1S92y
9uOpBeqKr7ej0NrQAVeZ9XZyPfgV4jWMjJAuJfdjiAdhyINEijdK60VrGS9auW39KEPsT0hDEKCy
mUqVCjMbyNMVqlF4dqeU9sP3r+26ecLAcyfaRjlAt/aW6Jvq/wvsN23ZPJ0DNSsaemPo1ABlDU5+
KKzhJOrLWcSOWDJ98IwQCSrTyDsThQD8zjKS0L3hhhsz/v53ZkquuZ9MiHIi7ckUlIoRGsG7lY9D
czfvXuSL1UFf64G4/7CbusLbc3g3ql+5PVqvIE2tOxOWJqZnmpjt60/v9651gelomFe0Pnr3/16l
EQzgjI4ao7mu0xho3uyjJZ54Ra70IypVo9e7M7hmh604eGiSyV+GYBmJlZffT0Yr3Q8QYpjZ0MQF
SLmrtOuLWB2G3UAENVx+EBEkYU7Yyez4oQ0RaVBse3z/hjGrxP8qJQGhWOzJ14b0yCTJNwOtwg5A
lFEegU9S0td7zWCC61/VHSFQZUpH1YwIm5Ix0Roe5NFohpW1LH/pGiPW0o3Vx5bUENkEbBRkUs+B
FYV89hrf6CJFtrdVeZX6Z9lwAXmhT6b0rzugC1VMO+n2gwWdffEiJ0UyjkHaIbmeUtPxFCVCaMuP
LxMxKYVGgxwEiJV2B9+f9HeSSGcv3x6lfVh/jCuxSRfKMvtUcV2NxQ5Z+ZFgrUhNdPSfi91OAZLy
4gbHOviFpjfvYN8i3KtuELTXr5yfedTjXvOEbQsouRjdl0d9ty5dAePLN6qeaoDWWJpv2rLBsYXT
GMzzbFhjd+4dZ6bKOJ1/L3jD+8HiRA6lG4VGy8pSDHkLRWt3FgAdBKv/VR8ev8Fy8B72juoaH437
0i2PB7EkqTwBk2yKXA9l4FLFIVp5LA/rkzE+sDTSN4aDpzr5AFLsd8Uv8E+8gWDb/Pom1UGTpEka
LCEgqWCUhBFi4Q4CaVN8bNaofQr/rdya7/6REq6guLq0CmzGoIW2xLhgjoBHzKzPB5OoDfW/AxaG
rJffa+WGSNfXkMnLzg3VDlMG8D8ByjBMcOdCCr4CEB6L9fXHK5qfKlgabBpUDtURtaDRqsBeJEZm
b6+tdsHDQn6mkEb9Lvf8jXF2ZXvl/g9nhEcnsMcRNfv7+pA1WYXjuHG66uFJYrjnllOqF2bHh4tB
3/Vx5O0nNa/aKvl7tt9pLq/BA4t1etuQn+jdfse+7p3CgKAKmHqKTJcWGuRtgsX5zxe4vyjQFKBq
DcjiXI6a5Bs0pWyIr0KxuPtY/+/lweNjepPdVdYbfMs8TMheLDNdN8mGNgDfFauPXXSM0hdNnqKW
TUfT9TlFE9bMxQtqpyaifK0cyV/jS/OxAqa6d3p1FSMLLAjcqrZfFQfIgUMquh1nRvPt/7LxjAhC
eCLw3NUhB0objEawT2ivByo+Hflt+TM70Ya0Z2sCjoGPABKNqPLtBP1L1dIQvTfaYlJB6zS/DRjq
F50oDmGpvE/jMLeJdwQ34bh7kQ6z1PrrV5uwsx4cwwE+lcvJnrQ2yXwvLgj5hhC46bi/dWE7zHsq
QjeamkhP/pEfuOZIZ00Z5demYYpz5F+FV21uejkidYborxNE6lG+vtFnPm119ZSSTJ6iUD9XiO23
997tbTD1d0y6xwcuK4lQlElIzXnT7qtTQj8xgDO2aM3hYoM1lpK1qKGSjQytWbfY8LpjcqijY5FO
QURVyA9lxmNBsrkJGJOQvFrjJEdchQK+SFG6Y0b9j5MyqdMyjbR1w2pPMn96hoiWTZxcJZbrOh3V
4d34FcQ9sYxtPZvaAG1u3tO6mOYKNUJqib5ZcGmFBRTZjrvp/+4UknjiiFk78xJ7jrhcTsIpEJa2
nBWUpUMHCVz0AC6UAW102VHyYNVCSLpA/MpMbH22UEAFGgHU+VWucWa/b0SXCdnlw8bFnUZ1aJIE
sGWc+R8i1N8nQQ92KF+Hoc215snzIhakStPl35+nEVKCj8WDf7eGLKwG+fMoQCJ1+4sE7616L3sK
I38h42PBvb3i6xcUN67hII64L4hb6joKqYArt3Lvng06T4WcIe4TVrRJ9146tiS524v/vkiFaLPS
SxdAA0IMqPdPXuDB8LkrIft3ZXxV5aPbtVKVKOSt21ydqNsx/INzRz4IWSUbQzkn+OxQ7zdm0Z8y
7JtCbF3i0PXShbLKMdkgPAiulP9msleE7o/zdylZQX9jfi2wVvEW/tZBEAM6MQeLP25KTPsdZ0eK
1SzW1L16NQzlr0PFF64U6fKpioffh8gQjtkRkq89nQKA1PMw6JXjVzlr4EAv4nFjnwa8GIMfcFuX
gHJsFMptTbJVMZopuKbg8pkGwHZa3aHok4nwqWgZfd8PxhLuY9QWqd6CK3XJcVapZU10aBs50xrS
ObkswJOjr8QtorIQPechcvxxuenW/5tWHrWJUhZfeYDJkoUlFBt8oVfq3qsxEz7GM3RPsOMnR4E3
NwB0PNMt3vdwaqD3+7Ppa3QxvC7yuic3zshmsgzL0HPHABM6yUgeeekFFXddvBEQHHSNVZ28Z+lq
fO1OGDJNeKfRmgQLbjI/Q6L+ZUjGiqj+qx9uBZWIvSoqmB0KkdqeNZFY42ik9ARxc2QYRi63cgMW
MmkPm2/DbBgCW7duFdCuDgGSjq8IH7L+MQswugNdiSZkkIGRAZloW71GII0bGRPhfRsk60OplSuc
1Ne1/PVEpcDuHxKcaRaOYn1Ey/awG+J1mO4sPA8qWk3ROkJPN8jrzun2IpD9LH/JhQW12zkQFf4x
2l20ZvhCOgXVJREtrxs1XTQ/6gYMP3OmESRvJ4zIRIsYD2VI4XCC17cKxsYjRbJdQwd02pFeFgid
NxQpi0+RadAvoEt8A1D6iOOX0Hrh/uHu6Yn5WpTBPMudZ9VHjo25hic7Vo4KgvrtUEaCJMd+3SNw
xQOo0mOBueZVzWFYQ/PFCyDNkocD0yXD0FCo++Goi2bm0ksj5xw2De9PiPX7/lenzZZPfZMKJB7c
GVAGEmLG4PCXSDXt7OQT+hamv120t616kYQjfs4o2yWJW8MIJJcWfhGWRUz1DBkMPLwIr0JqdufL
eoT6Y4eqCG6lXKzzNoGXVLt9mNdEMy+2tb5BjiFHE6W6iq110SQpfUfaeerJIkywkRbh+w237LcA
NJTqDFIZmAPohnmCaLM+dWvQGYFScLWrEw1QIEdFRs7BBvKysTbad8Ml4N83u5w+3f71Dkj6SFFo
OFzlYsWuIvGE0uqWU/5aqeNykX891Rdz7oIGZV5fAhUr7rBb2zNrTIG677ebnhj4Z55NlLCweJg8
sFQY1fVa+zJ3pDrLx0R8NGFxQLlh2Yn42trfdMSd3e4PhqKnf5k1Jmfoc4u07VGlRbsFONDlVmU2
QFMFnV0VEvDkGhxlEpPVislvUOZcGCf2sg5+vCCncsnOTY64bbuO4Jdt3NPcX8hyYik9WLrHkq0z
Dh2WbDh0vG/qpaPTPgpBhtaKW7WIuJk5ny77aXs9ZdQeNwjI4ZBvq7DWVxj1MAlFYDK5Rjez7Zkz
ojY90KCJ2aae1j6qNohvs5cVUgHDWtvbKX+zJz87mvAQikDvcPMeulccNj90Rlays/l9XDqW4Q/l
pS3co6U8GwYOpeue8YLVSkHFX3CrUeLqGyFNWpO4WnnpqWR7QeJXxZSoiw2ChiQ8fic5JfC2UJet
Lgp49kVqw5g2PEBTSELDxAmAVnwTRPoJSM1cOVC+asWoGMrg07ddYPG8JFnazka9xrxJMsSyd1i3
ZVXpqoUDCjkMRSp8uRLzVfCWKRJ/Vgtvlw+ZG5MmDBiFq+zKux9NS5k87GFQGRXdNU19HGEhC2PQ
BtJuCjSS5e3KQMPYNKmNTCjL/Gz+nLxqF/yJlKhbNfLU+YCVoCLAugGHumo+g/5FgLtSjIf111z6
DO9zOP9uSEaxBo5M6wJmR9aRb2i532w5LIqBTedb0TJD66YDEB9nuWUt2zhMyKOD9JAp4AYEPLLW
gH34YPTbDOHUiiet4gMCefzNRCPwyOSHT0RuaZZownESZsOg/3AbERbJbwqLsi9jeqPflpMPC6e5
Vw0LPPQNa+ovQiYCibtsyXi8zFQJDLKeNEX5THEYUUiYnzaBDmvX2Hbo9Y1a0uba6tvzuXCOgXmK
Y13IQmLQ17elWmuX0MMtLwjh/7mFPTRDPBZDZ8QrwhuFLXL/ph1m2tbJWBrN4GXoR8utJWQ0cVps
fFgK5KNAPoOkL4zRk6KML6o+uT5epm23NpYN2pMtV1WPSJGjPXvnFmuzwfqZGxZBbGjG1biwG9lh
kmseeBpG0VcoBmLcDdvHc1FR00rStVhr9d5zOxu6pvCeOPc1CN5wPP1PxOZPLfjeRqQjmoRlGbWG
CY/IsBsWdHmLhI/Z6b8JHmc1YwWul+2BASJoihl1idLFx9lBRMLgUd2CxpBHulX7MDhPMcqby79Z
o2cGoRITEv8iYs1J0O7m7i3+INN0zw0kjYgxERvqnuUz40vCvv9oISe40W3ZiT6sITScW2fiV8no
BapKk7fom5R+d7MHQC+fHb7hYXQogSmky8PZKd+KEnctMuI0YpZv2/BWymkcVqBwmbdme/zZzXRI
/w0RozTxqEALzgU7pWjyQuIiQg8gpGUZZlP9vp+YRUoMWylL5ARNxvx+xS9YRl/FD14HAPj5cmau
70ezqpQEpRdP/2SCzccsC3xTg7hQ+MlXCW/TnJjb7DzBZC91zKbZQ7c4OZBkba0GcdimgKuSLFcP
5uxz1auBh//S58xo4KFLaFJT41q2+FnF65C0RmoMsVbYlvqvsEzHQhy4lVyzI39oAS4zJQbWGSl6
hGCpv/4tEg/C/Sy1HAOysfhYbayAXsEwfreMUI8xLdYRcsIeaDuGjCN38VHuBQyQjAwnQvnabcL+
GqvvvHbZr42J/1V4KsKHnf7x5H67ZIxhPKn9jQcob48i+Cn8BLPEld3Ios0TNWqwZrY3zqFlNRGa
TfleFkbI5IuCq6eKGKCbgFvuR//jVAdJZetCFuVJCR7AEFIynSOCSl7Gx0GU6TD5jMHEPkS7uLSo
BaltdzvgOKzXPMm8y3sY11xk4mkrs5SPRQlnPDA1hZmOF4CFU23F5usg4l0Bn01BxMfP8grcGPkt
y+Bs1QUz8fS4G1nHy+YMtFP2Vlp53sw235AHaPcC2EHcbk3Zmv7JOWdquj8pjQlwxue52l4/Rgcc
gkPlo0LCE3bkMTt9+6gtbTP7jzJ1k9EVG7ctCQIUGspYpx8KnrB4fuL15I7CDx6uc1uM6aRAifW3
IMIIDgMzQ5xB6XTsQn4RWIlKw/tYQVZuv2Ym16S7vq5esSPhPxcvzS40IioKDREWgvS83jJb7JKp
ysZSgqAYdYqsVxw5zMxuP3lz5/2WxRrevCOvi2PXiVGWxV4Bk5c+c9kR1RvwvNqNVWACiDoIq24C
y/5ZBfl0zmLjR8O+A06i9+C221k+toezhwFqRYBI2Q+GA54PzW/wy/JnX0ZwnC3b/wiLOEdBWa/r
pVdBQeExwnKmK9YG5C+ucyHC3DMcjgOwdcoYBnSYzfv7W6EWZ6VR5zV/Bd2sVh71wx9N193CO1R1
y2pu2+1cLzs7oOe6UIy3CQjs37aQiL1xSd3+LC5OhXu5fxtQt4rTLvgB39ISHgUH1crZIy4X8FbC
a+jkyYo3HtemB5KOfCp5xYpgK8oRXKXLXOS7rbnjnZehMLvWt4XOmuZ1yFhhqaX0mBt7NQTSN2E2
PN1ayxLNh1olA0a+PqtHp+7SZ/PdQsDDHgYdBaSjuoMLOlFNIE9EHXAlYY0HnWBdsBWE2RVpuQYJ
lChhN6CYjdph2cbge7R/RcHdowj5+Q+1jlatCpniqqz8RyS8Hkl84z9ENhWhyAxZZSK++aOmqe9K
4L+p139OS49BNRTPPXF0fb8kuKTixCPfN9rgQ+we/koYSZaB5W6EuaqBVkQQM82/LC5Z+VpStYCS
bsNGobYCR6qRXXtiKK9RHOUhzSaUtepifkJzvrSQdTCFPN5ghO6axNloigrAYumAwNrxFx9guxld
X4CEZ+NscVFl5K9Jb6nE/SmFpwub2Ncz0cJScyzDYl0iDy4/BKPFBN2znq71ELBJYSQgFvAPdE0s
vgHSMbarDoKd1aU+E9iv31QoJlL/hQpSiNF7mn8WqoTFtQqZWmopmAri6DDzZbipR/0PpjwG08PA
x4MQqlZd8IbWXzrgaccFHU5ZbqYGmlCPQQm2MKvxnZhxZdKAnoVZAyX0ICKIVZom6rJp5uFkM6zA
tu8pZXgilXg/ZLAc5LRfYaoR9dBDTd25DrMYA7ZNAANn4y+MrEzvysWmQ5j/UqY9cgvv0CNoU+WV
6SBUch/qc0kr3YKCCPg0TGF3XjDOlnw74XG03H10jOhnyMLVgBvvgZyMLHrcLQ+50Gb5H8NU10Q9
t1dxSs/0Lwt3a4bAYHLMIP7vDsYCCHH5o3m4pW+7zVdPZUnrPuE0jEGtKeBhAFXnqIJR4TFRl8vc
KZ5NfKU1238gtcvMObHfADGQYfDKmBO9eaAwm/kDOhKD1OshMH2kr8/3ssz5DniVYbZBOlo3h8hg
TR6E+xfkJrH2Sfeu4ecAnyVfwxmWG9mbuErck1PIXUTck0AxBEMBVEHEb+9LyxPjW5FiveX7hedA
tQiQ0pQCQE+rH8hi1TSvhaI033lGWbfejAfE4STQqT4DDsMUl2kLfDVcgauxGlo3MyNqUICU7AqJ
dYPCioKtnBZ/vhJJX1q3WS1EZZflkQzEF/l4GK/V3QaNLY0bC9LNqBDuUA+6WoOs4r1c1wREacQC
ZERg030ZkXzyvxLh8XN/dAX+IfR9lc0dhqcUj1AlqbLISLiwayA98FrOhqxxzQnu7a43BzTqCty6
wP8dQ+jggpkMSvX4N80gLCXEc4wGZ9RoX11ZvP7mTRlXKVTAbEMpJb7+lY97FupKPoOjULCYsFGr
WW3dzRqgHSgpQa4k/XXTop4+k93zY0chtoinR8qRpd2Hqv7tiw0O8q8qT+ASXFWLso6eCmQZditY
eMulPGR/ggHIAWker14AXNScqKfSYkonVX3VWZZtpUEpL5kiVcqhCvc0I2ZaRvEGpgCawSmVV/Ut
eJ7UzcMNy/St71xxAKMD/5Dp8UesQdVrJKMNQiTNlD7PeOq8D33kliJcNflUKFgNZiWIwAmn7zN6
KWs7ps3R0MSaasgYnDaL5oiwpcfmNy/UM/3fmVbOk8VQBV8OsBgukHVdiP1IY56c2QNg5ppR2gm0
6/YtUAjIQhT0ojNBofKNz3s1rbZUI9l9S0d7Pmp7xhYv/0RQtDz3WmVt2SsPVV6wmuILa6j7Cyii
BCOm1k5ZhKTzDq1U+4m0jF9JsrSeqfg3DQ8sFlPABBYWrxZBKClnqzPxhCTrunH20W0+8xipZ2AG
b8+0CslYeoM/3zidUYKhEfF0ADoz7zZjb8EQRv8m6uCQns8lbkeNUQ3QSLSf1gI6xJK1PEtdPeBZ
ADMhnrsWx0ArdbSt/7yh8NGdN/vnyv9HBbjfgOWVWDBgk5CVunZF9VTzVkuX03DXvNrOaXLadmxi
cUTVnEDbbeWbW1bt/urVrixd5pIX5ODdvZwqzJbgGwUB8H/0/2/haH9KrqSuBs8E0ADg3ASUUhxH
1IJtYj4I4lV1dmvrTej9kMH6rG1IWcBOUc6mQZX2OcxpGn9KuYKi+IqQz1znHTH6n7EWR37LqGcW
yrA0ofowVeUJP1AkaJKGeoxK7sXlfOwzb+l1sEIjMUWM/B24bJeeH6kw4YgvMfUxRinhw3ltMaPx
3V/cvurVqhPT/sxJNDjNfdgznY7vbxLPyYiNov/IwVVinJtPF/Qr+a3hCcmclcB9lBfQhYKOpUe+
IzfuDnkIpausGdJxG00wBsLnGeW40z17oSXJtBbRP1kvky6ru4Yb8egslsufXW5Zxurzv0AcFO4b
EP0KScEyTwQv1fRXSIJ8eAYjsYwt1QIadx9zOyTd+Cg4U+7Md5CQj6NrVNdtgmABIL+qbPFOF3p8
g6RVqZ1HPHe9Y3F2gmV2PBiFsIpgrNdPbO/6QfWPikMAfMtqJ8wVyM+ezdCuY2KYyvh7aieh3sqA
zehoEidJNmBndIy3W+L9rSM9UWkbOL6gnKr620/M0pUAOESPeoz4CeqV2OPGoq1XL74KrxR1Xurn
DEY22dCMvbx8VDrz/ELj9TD9ZOKsyzQMgYHhcyDIGjxMuXnNQOcE+l2V80fwmPup3DHVVAQ6pi//
1WGkjRP3GAUbEKiGKwGM6DFkvhQFUYkkOVVTJEdpA7HQywLpYcKemoZL7bBfolX2YvPu053vLZ0y
EJ2g+Pi5UnmxXVdnnwCirF7H+Idqj+xY8gbitGnUFGSqwOemiS/WEH1e2JWwFB86DXi52d+VL60Q
jXnPHL0QwvGfR1J5kwCXEgPImaDerFAo9zbEOtB/u6safFyGDUTHIHJulrq3T6fBDR+/O/L25TWH
cj+xc/yoyXihTy0oD1mqSSf+ONIb1F2IfBRFXb0Vg1lRUqoIhbfn0+4JYjwBNXpoJ11cUeiJKJkb
9nBJG3HRcXuXMliJxTHkfnvE33R87DDvfjU01aAjReiMbm0w5ZFJq+4Y7aqIS4KoNZ88UV3oO/HV
O1OM0ao6QeO5QDWRPw2e+9iBtLkXoBYhJeq9rHc0vXfjBhyAaE3FjP5uVVsNhHqcPRJbJ6kjMs4f
UfZP4nrSBI3PkbWw8Mm7jdXTOSh7bIsVSCZNmAm1IFlLzahf39ZwfS2Tn7HndCbO6NNpaljc68zA
fHQ9HpujF31jDx39bB6pwiMjouiaAXDdxTVt3Tzkjw3S+qaZJUqL2+NTqFxObP/ktT2rm09QH/Ge
G75G4FVH3sKxmsamXR/2NWZ7gHudOkm3QabqZ7ptrHZjhpR5ntEbbaZSY79y+cIheJVG7d7tpK99
LDU1N4Zcq9TLz4Qh82eAGHAEacd2D4Nbt2kB6aIDP6ROw05r2XJUV2x0oCxlX1YdJGKQnX3t6j63
sJ8tZcJDOtqvlT2FqLQz9QWAE3I4t3e6lRsjgecre7hgi/W7aEQ/BmfCAkcj1NqC02sochMCphqx
QUBc5RBjl245t7KVmE7v6uYfkPqmkLbGItNaZeqtp9I885HKjZ/9otrupf6bvKxi2q/Z18MF25gP
KDsEn1GH+uJMQObJ3jt7BJBOzMq4gFmA1VI3Y1n/VGbGk9goEHA8XJNFPJTT4IvHMGfTUfkuxR3k
ITLmguDJJdje68AjVWa+gTG3S8E4FFce0v9cz8NOaiDgxXo00Ahbq7KMHbBKvr16XR7EI/Oh7WVi
rpGCCdQhvzvdZ5RDO8mJM3PBQUBY1KstouG5uT86GinwXLuRV0AUtAwks9hpIeVcDB8lVCu0OmTT
YB5zunZFvPc7vVz3hBnGQo1iZvstCzAFyO5qMsLND7Drq9JPocT5HNnPOUOzflZAjvEOSixFGJgn
Vgch5gS8/3PRhjKVO3jbFZYZOGJ0kQfcrBayqn0rnz2jHKNeY9ytcK0vALC2fZfMSN+dlNXjBSkP
R+DA8sS6eXK8Qdy6DnHSRy8G9jIn2kH6rDimdYpW3xHk5gltxj3AwpNzWGvSXzPkhBnsPD0t18kQ
B404zR7JTy/gTyajBTa10RvMXaaP/EYKWMBK+dbHcZjuuhO/ZX86tSWmg2J5ZYG3O5ZfKWxHyY85
ie/UhiUQYi5azpM5cXTOzPSLVKKdYyRfUMdXNR2ZROzwmG0FY6eUiJlpOIOjD4Lt57bE7WjM7cLI
4yO33CPpLFrhTuoWzBAi3EJfgXhKESixA1QVNgi5WjVAYtZjs4F2NcO0+CS+gBAF8VUVZ6eLS6mA
75h8T6NquZ/4+CwLZTTNktBY8sgP5rx8xHdSaPu1dIKqeQJi15zWXynxUWuzBrBVYNeBxnH/Z8QV
Tsrc8ZS95MalvND+oq3knikMA/zjKjU5f38fY/rw3Y8Fac+bvUoQu1ByfDBRBTeliia9NUyp4ngW
4tKPKupfjpWxHWolRCAYy++ldAQDDGGHrZ+Sgvno5K9fQtR/+6skzY/MurYsJO71tpu1TwYD7f4+
1hx2LvSMADNG3riA/lVInljmscCaKejjXk7TaUkT172cSyEB+YS9Tfh6cTgSNZ3DHHIE7suKQ++U
frimBIDrOi9LMm1tg20gSc+F2DH/0tYPXrXIK72kBBl+xKIuyak9HXjpzKiHo3OXnO5ldEFvbl/p
YeE2mpJZh1s7eyk5OW+ASGAyKojZ2qsM+VvwLqWzWwU83fBiJwAUoM3mG61cwRNgn5BzieM9Sr0G
2lL/ebBGcTJyQqcJ/8GLRQ0Jpen0CB4V/egJ9Y98PMV/VRVcE/adTDu/frY7ZxwM665yohSyEAcH
HtWKquFMzk2/hA053hFI6CLQLyrGfRP43H1lilFT85YRkaPWcI8ZBY5mGKy8tRlRilJpAh5rSRJz
CYyoJ5GFpt+J/5szVRL6xJ+xzpoJhw0GGEEspYhcaYEfsQl1rQQM028G5VREbK7sNNh9h4XGtuom
MSzqPhhhJhpBq/FKlWh6o+OFCHaE1YfUumHWqaXI+djEci2BzZuV23r0xJHITgztdLmh3L59OsHY
okXviyBe36aooZRuvNgYipgdr0n7PpxQQzLc4K6CT0kaRelgvR5YcsKtiC5wogNsve4n5MLyLr6B
dHGJnQDA7K33T3nzDl30wPWVvehSyfFf6BVu8zvdapDaa7ae2pu0u0dnCw5TKgjY42dfyBarJqP2
FoD0uACAMVROCp52sceKyQy7yEaLvpzQcaZxCrv+twxMDQspatejvawOApNmpf/H6kl8BR7CF01j
zbteZWyXQmcY12ypQZlwKGcW6f0YBjyYrPwJPjg3bJkZhAyHwK/E1/D8d05towT3svWxyutQM0jS
2eHIWM5uBBo0+hrwmYL0alkFtmZyUHkpvR6NS9nXORlUQ6dTRNwn1bnkPmoKPLqSbCTtZppx+R/w
eWAdF9UXrEs5ive5Kvdco7f6wAGFfAP+z8zn+p4fI89vax9FeiEspJEk/tL8FXK2XBWXbeqzY2wm
iui22wocFy91qAWw3a/s4FG8ylBgK9tvQu91sejBhXfFPjuYF4+zMAWUL/iMV3cKNpAdwIahMt+q
gWxEA22dh5GuM9eDSKRsIW4g+iw7DRKIzIJ9w9uzqElBcxBQ7VhlTlc+Y13pQrCOqGZNHP4eCO+2
ERu7NWOlrjVzwHVLA/IfBEJPrvmbfVSxn33XA5YIX8KQIbXAwTzJn7LlD5cxZ5VgZPv9zkUomCFN
/GViMvvI7MR+v1PELEvOPc2nEfS26snFIoeM/46Lgq+AmXtzeH8vSI4akF6ZcwPX7dtqDm0fT7HQ
RVhhlsN/5f6FSFZGoajMxW0rQh75HifjdAyLVaKewcEKsBSt/QGvIqFG/OPIJUYOGhAtxUaAH7ZK
ygFLeuias1ERiIZTNAAQQYzE9Ez27lPtBjcRWKCicTe3TzEPQ49NinBPMPRjyB1BHuJmJ5MOsokb
21r5oScDV+nw5ZnWoRsJutALszNgzNCMCz9x8nD65wUht+8yToqDdxtE5Zrh95ipDjqZL9huWrX9
c6lPoorob+vTTjZDnocADocbZ+HMLNnTv/rWeZVVG5BurVqhblvPlLrCT4IUMJCiFWnOjQcys5R8
lUleu8cuUXAIqqOMfIpU2mJUD3rwqTnNuW6rUzIE4btc3sAQWYSpY9W5oKfn8lbAjG6sqpjl9M0n
O8/gJOWedLcyWpmiL3gwU9dJ7oqoEG/1ZuvdrgmNAvxL+WPEEsb8ZrxJeoJPMFjWUqzie/meDBk9
X4jXuSA/cnaQuUNxni1mBv89yjys54Ei7gYd57bYVvBCUX56EMab6zstWG66G772qw9Bk9uyiDsF
HJdKW/0IVGR6swNWUW4hIsWC9q/TPm7g4q4Pd0sKYSWvivG9nnsZbt89+sT3gXm/gW1NVofu/HB1
V+rIbn2jcG42ZpsRFRJ9Hv3+Xaee07rDv03NnGvSMil0zXxM00sUR9n6hHqtw+o+P+CSGbf08+8p
BFT9xaK84xZif5QZr2UdDT8X56zZh9M3v9ag77D04YqKCJgdYfxcinDdADr2Z8DrLw57DwcFSmHP
7prM9Co0n15Ij8JAUwLvyiGzVmz08jcl53v5rh6rs+a+PWzyUWRXUIPsr4fm95vlh0VNq1PDR0EH
3oYzMmsFZ+8wsuR+pFtetzDcVTc4GKb5MaK6E8DGMWT86YUNHZd4vvqbcMN02GdJ8cONiz4N2d/e
aBZRROncvvjSGYiIVjclns2BOk+KO4Jpc3h+r0ajt+bq7fV2iDHH2GqWz/cvrXjA12bybKukl2r+
qBD0i/2pfnDUYaGFHie+UnDqIe5fai2Og1ekT5QyB7o99PRAgH5RonfqBtI5yeWG0NvkP7TAecOy
jUMNi7Kd6e6pejz+Fu1VmY4Fdq1FbQmOt1f1vQ5nRLZ5fOdfLSMbJz1Lgbv+ywM5j6TdywTiQJ7N
1fFWxTYRRr5prTS1rqNHYB+PoA9k0883OXV/yAxFiodNgACNnvm/vjkF6FCQGR89WcKVX0inyWuB
zeiSGH8JLP0AdhniFoo1lRSc/lAa6kurWVHHAnaJhGVWMjg8TPcmdl/Yp0lk4VQMBhnI4SeyRKYw
/+hOmhBbbiYCTbFMGbZJl7FuQVwXWRyq+V0A8PCConojDTlSHYHQjCpPpsMpndb752gKDRSd/0//
OHB7lJ63TjpTvCBcSFxuEaXwUtm3DndhB6BPvykW/1eAuw1gWqIx0yoHdjDgRzPYlLIbG6Vsc8s7
QTnRWYD8vwavl/R9l1eamwnzxlOYRySzbEIFjo0yVLO8iNJR8DZMhKm2CJ9Vu4Xf++VfEYbtOYhf
qg/0zI+ZYUIEBaqDRvWoEiPG3FzHMj8bZ2H3soSe/j46d4yTTbXhtnKqQ6YTh4MM5sD0FxBWNSR+
YqnMgsK9o+tBgfotRKqA+JFiLBp3fSdX6eJOP/Hkrz1YJtbygFtZseJb7NdHEGOHPIFOsjJWN88Y
fPAsdtgXZrq386St0Pnik+B34Wtzd1vl3gdwAjX/ei1ZRP91CrqNg/jIvLlqNvCSFPJ17/rMY1Kb
YIycy9xZ5MfXg0D2ph6Pxi+zzW8Zowugw1VYxTl11qkA3C8P3pLeda6BGUe7TRJgJsuD8MbDV3YT
o+Ix1qPdP56OMqkgiO0h7/7Bdo6x0LR99AGnZh5vgVN91nOSmR2rWqkNsSFTfRESP5USUOYO7akh
ixKGe+ET7EQBkeY9docNIGcLStkRTVp8LmyyeWYE4QyRyVN4qYI0EFKN1ddZ5+IA6wnmKJM3DfSb
WL6chusiqtW9TfomPAj9g6pDK1viiKdX6ZlED9msX5yDGCcaINBHJo4mOtBHuqr4wpczKKVWxnMd
SkcbOzdg2bLhpErGJ3qu5BIcYBc9N/qN+QYTPeCB4VUwL/6lsLe5/jj1cLnzMRBBEXxZgQ7If3fc
3idOxPCwzdktH5KlDG6worL+P/ZwpS+/LklNsTR6lpnKXqpMtcH/bV2kStnLC9Sz+M1/WxLQIZih
Nkzk7aU7vhctdqbxzr8FY+K3IRLBZQDl1p5UXqV3mZU7fITsO/n1X0WPK7GMmq3d6jl3lUIq9dKN
LXgR27O1wNxwq6ccrJgmSV/D84rx6kcXm8Y+pBHPSo5IGyELOx7PldG2ZOIbDyZbsdCyQVCY05QN
m56r5RhH6LNCGFnfUjHi8Hiz5ucT12dZQWyXKaBEmRwMOawJZj9Q3nhn8wHnyNCM+4beQLjRIlKx
9Dyrrv+Rp6Qq0yGumBrF8EPyx8sfHq8XsJmRT98Tw7lM7il12bv4R3OsTZLbLo1iKFinMfOsPSOE
Dl6cX2VZo6VKIzdzTmFMS7XCtqG408ejVcASCuupERBNIjPOqZE7YTeJuYquK2HFHULqyXZgc/65
3SyQjvqyTtSoS1/DC4o9Ch705KtV7Mtiu43CR2Cl9P9UwbcDwWplQoA7X32TKIIsnPq/c3tzrwnW
USPhNURztdDbSLUZLFp9Rd+Nja1Wud4o3ubBXF0jVu6YsBAPYFtRQbuASI0ajD16sIq9/tZPR2vF
4PU76h59zNtcyLj1mxsQjhohtPtUmokxxV9XQNuqCBveDcn0p5HB/BB49LuMfwqV5KmPEcMXR9uh
BQ3tlQo+xdcMZL2FNs5qv927NNaYA8SD71gqVsUiClJDt+chMaG1q9HncHSUXJC5ftvTdOd7VmpA
P7UHuLApkRd4Onfk3AOt5VXbGFW2ApvH1+M3/qPi1V3JKwKmMV9+LkwoKKN2xYpMTYMlSQxcuBBI
259U8XRfFsH3iuWZlDpjPWU+dGQnA5EkkpH8NqI5mELjGRUcYb9vVL93Q9wnUMKhJgWkPVcayj2V
YJIOg3PgqvFh5Cei9K1jnzTmJgnyQz+2SoduYGH1u+iI/NGOoK1PTYUM+0YGfEVFypoTHaSYMPp1
Xmp8V0YmQ+T22ndvnMCOeHFFG0HvzPWE/MnrqD4yfxE3II40dA0zl9J4iw2pH4ICvUTg3ODnl2Zp
AV5g5yTuk4C17miUttqGRgDxvpyMTAzbLz3xhkXa5FHa+cToMM5JS1LfsuaUhpbE69cqRkFpFhOS
ro3p/E+L9Kwm9PFQvJfvvLIVlE1OUWXPedCFWZZLZotYtMKPFqDky0Ohux7fad3A1pL05hYxrniv
Zmc3nl60omDcWNQH9UhTz2NMhisItkx6rLjRklMo/1nvuwv0Lel0gcKHEBxW49WHbw+BGnMX28QO
BHG5FGXkWCRRSAH0D4tBL/E+f9TM95mhvzVZg7Z+wtMMrJaBbwyzZzZHfyr207jXsEX1DGsNES8U
ewK2GyzO36DAVgO6Ya5eEKsz0l7lRrnWPlTYYWEwwjweDu1S029Way79rqVz6mkYLiQ6IESJJ8E6
rdrQyziRiB386dQYQVW4kKHduNz0LyeqCYdPhyB0VMZ5e9+Zptid6hr1Kzf91Rf70LfGanedNLk6
+nDb1LTbwmkxC8hvVr/kl205gFIGnr8MihEPKWlRuOctm/qHxktrl8UMLErgBi9CgWkh6opW21cd
fByzLP82508O4SWPB5HyqsSMxB6VVLKf7Gs0BejIt+RdBrVblA/cARYWHZEy/0srobnfLINKSru3
+c96SYySVnWVr7xNBAcqkDOKhZfAAarfqLMWeadsrGWsziPpJ0jdphcQ6aX1jmRd9/s+2QQnyo4y
sbIMINSlIiBKYqUH4uwtZeqEQIWccuMgDVHStiP9jW7i2Ifu36iLDXey4tP1IjGwZ7JvgS8lbF6r
v/G49kXlAt55WuKIgWkv7YpzmC+5o4+PNbK38xUaTmyEjnUP0j42rI45ytBUygkfrOqg4bOLBmju
6+ZVtddcCYISDSLqIrtgflGi2om3xt0dtRZnBTssr1NDbkK08wJcANvl57mexrrN8LK9uNJ9rQRP
7lZEz777sueVD3bTwXB0JFYuqHrw7yBy8gv191LY0fXj2FJSqqxakH3ejOzCcdS7LjGH0Rsgfzv5
aOqEZqbUXlefkl4EkerMBD4vMLjkNNRvxwsEvR6ZvXr5S1DQ9lce/1vOp5KDb6mFxTYhqWQq1y4Q
a77ybvNKm6EZUyokpcN+hccpIRHqbVeu7xlHqp/xEV/i7x3bpl+dkGRZxhibP9xicse4Kn7iyN+7
BVoUMuKjA2beS/672Y8yWLCa4bUByCTm0pjtaqQuzoaPpUzJat0xRq27Hlfnz5VLdLhs6RMuyWPI
a/k1N+r3oBWuV7qz6h+4Kf1s1Avw8/tZ2TgXj6N1+7UEudxsA0DqjTcG+8KUDyYOGRCwcKK2A0Vg
vjK2Ld3Hlxjy0uq9Ty/hY1ZfCjNatvhFJqzRoetB9n00sMzrUgy6ceeBBQlgoXfkhUFVXsZ7gZta
+ZjqzHchLx1FtWC1MvNlVANXpRUjpkYoOd8bl4xialGyQKKGUtUceV3PLZKy1bJlmtUWVVzgh+D4
oofC5RKCnCH53y8AT13T4hSqySqtZk3zSkdVzmuYCbxGsh/FevkYQtOXH8Bri8Tu8O8eKt9mFCeC
mIreGEMFsS4Xk7dTiOyGcBRJ54LBxfOaOkyyHBswJ5PqFEgWOXpT3ZYldwu2YlIl5G//vVAvVI0a
CnGZW8m2Bl9c6gNODRLcwOZa+2GCLYLlYR5LinNa8WNDCfX5Xuixh2z9+H2+wqOwZitASczBDpre
LQfSmBbNmXOkw7qfMliX/4fjAWGfSxpDVagvRF+XndRF4R7WHUOJ9iUYiic762d740PLlquGy5Sx
Nm8mEJhcnreOSSVHHly/ESaMqjiUYWwRcFFlRKNMtQdmxS5xCuqomXu3gx1xajKclt0IQ1pCSxQo
VCalrHbwmqw6kn43v07gjS6VhYe92W5LuS+XMrMeQSIITZRhkxodPZtlfEBOVLlj8abKi3BWBKMN
y1YXNFG1b6d3Z3+lrO7RV+O3u/GvuB+0zLKUcVf0cs6IK5mfBx4Qxj8fJSJE6pnRz+2RW5kDXrQY
tviOWQiJ3N7Kq+JLxxm2RnapXwMWZ2PC8ZV1U8dDhzXkLovaY5sdFnhH4hlR8GfITLuZJ0GNrTdB
Q6vdcb3wr9oVrCzm+o5Lf2YQlGKkRIqczWDUJIB9obVqRLjUyGQBgfbaav4QM0lMtxIBdpw+q2xu
jSIGX/IkQP278tRrGEZ5ylInn0bbmrcQr4MiRvdAwqG67zo9k7x31/cF+ZxoNxr84XAO7Twrn/1Y
HvdUAGsqFZeHHTQ9MthAuJY2k9aswNoTo6Ag1u+YhqBllJHycXwTEjT73Exp2RJsx+Ud8Jd9b8Mo
HhRwHXps82FS9w1UY4LQnoR4Ma5F1DK++LaJKJt4ljy/kp0azJ9CgBOb8GdMJO13nA/r207DSh2Z
Wk510PH/Y3aNTIgw16oO6WkUB9PRhhdbH4SwE4L2fpwH07xixiMSK2pu6oIBOGCgX1Cxujwx8XTk
w1KG2h4dfRfW5XsoyRMExD8TSekRrGAVkeJ3j1mw4CeCIhKOW9N+rl65ohAWH+sLSg+BXfcQScUk
Hr0jqTUiu4ADRGYhcSVaiq8qD57V01mERRGNHN5fjhavYz4X/IuG26mfvdm2yqzJuAbtgas3OALo
2liEllTyPVXp0nsut2PD/3enzflwngfv44Vj4vRRf/2mviUqQBzWUK77V42MIGV7e1SWVZmyKYnx
xdJKEosJ83+irvXjcegijcI7ZLOyMgm+vHAly0sYP+I7ztx5hI7lfImkZI121ETpHruRSszVlW+Q
Xyu260x4wtKsGna/evjFDYgkubm8q5Xx/XI3yUwqN/GmoBfFFObbgz5tvhSUkzEZEADTXL4EDyya
SGLQCSjY9EYbhwrmm2CROH5SzHV0EQQoPlzSDM2dEJ+V5bnM3fQNEkyUWIMNzSyKlEQGAlwxHemx
AI3w/PN+r7yzZDHx6WkIVM8ItYVkuLmIXiqBOf6rx6LjP66DJ/8jdcIv0SyTrSo+xmkqVVzZ1y2N
xNcyu/KCTHMppxYOubZJACvV09zogjdXY/S/kuPN1w+TlHjZkzhoHWSR7vzoJY0mhTGSXQmwWi3H
3Qx/VSKvI/TToIAlAih8kJ6jyLStyFd0HLLo7KC5IrZM2e/ddcHPortnoi2F7g2qDVeB7pzTqpA3
R0S8EDvnZETlDRCslkFguMw/cGNVjKWXx3IPkjM5UTC4HzkRdn3AS8N+5FEwMM3cBLuTDJ577Dn9
1suw//CrvwqTIl9OAJeZyPPScU7C3dnHDRIWeisj5cNWtu5JaT5DGpWb6Ct+T9GkZXfcO8Fus9CY
1FHL5Iqn9xeKC4JGHi8sE99uhARIYW9+SiJsPMFtv0nAKSQzg9/oIOHKn0+YzmuRnrclGo3RTMA0
SrhNdVFsy7QAB1Utay7xWulLEVkWZtJFGcEg75b5djeC/DkdDUkEL8TYec509KQup0me1VuGuveS
uWxreNFJrqgQGu+Otdi2aCwxvHdfz6DpaaBeQGEzyDrI9DX0ZNoMxyeMtVPSLXQWtzfQl+3jm22w
f4/FjURNc7fNSJwxr/zCUOQNRqYWrj9a3CWYto5AQ80eT1hsboEDcGCYOxP4vuVVqnKnMsiEMmUZ
wenXMKxvdwnWtPl9Vs+SmVg1BJswkZP5Q2iuwnRRRsRi/lmVo3aIU3g3ZB/shht7wOCj17q4c88l
9JoQhBso08eUqjtxYxhsh3osC3dKAHLlIkOU98GADZBc/IH+t+kHY7Cu5uM7vpOdQNzdcLzkypnT
tseK3wDPb2DMKpBk8IEZ3XVioOlJCHG3j6WOtVcraYBTcf+RDKDtcspMgUkIVJI8Y/lz5An4ccsn
WLiGQUDPuMJYsLlXpAY5VsFcw2iHlmcricnDQOZC4OjI4BlSQs9KAy5LlArSkHSb9YI8zKivbj90
H8jdJFbBpIfcK+yxj3WCv4I3i1yHmynNhzksfE/S9M+pBs+H0iNYQPMhiJFPzKkdvpTrAfAfXD/9
Jin+Zz8tKQjEOLYirqtAescaJ5PcZlGMYYEz8Rtbyq6+KsA6Olu4UxKfZG4nojFjfzHfjpBvr4wF
DhBpa5hxo5sL0PWtfUMA9gtpXJ6HUDOyG7V7xvsIAEivW3s/axVYEEWHP6SGvQwW4MYYJ0hO2Isx
/m8kzLMIKrhUdK4ac4MlapA7WXNDdOmJtqm3ldM5B2pba9YVQInCe3CnLr0YSdLU3RVA9KFRpSFW
9YmSLpxPfB/QpWR14ktRHdAELIzQT/Fg1m8RKrUEQt0t/pMyqne5V0mzb5CN5xWybcQv6Y50a++p
JAZt4tiaXW/635AbUrLvhIn8rpJP+qMNl0tM54FMyt78zLBhlNH2UB8Q3kqhbSZUVGGkCJfZPcK5
rs1fY1lBUV7/Ewvmf5zuQLscRltk9G3uBdDgve3MKWoynnwK5qSRCdWc8Vq1Iya+6mVmtofJtnc+
dD+Iei9lqqLblzCBW6jpyYJv131m1F4A6H57GdW6VIhuEmVNcl2AkLjBWUC7M0ZaZvZRBfcHNCR5
FRfeoJ25dzAOZfe+/zggOmOb4bE75JSE8XW33LnRQeEde5qklywd8So920/GsufW/xmrpZCB2+Eo
+oXmomlfLB2cydbezEjxrg6j5BNL92CC6A1GFSOYS8vUQ0ot1DaCX9bedDKnp+dQKYVV0CoSJdRg
dea1qMmNN8x493Q21vk3ozmImRDFde7SpERsNU0UYmu86DOR883v9QCMcDoLg94qP4Ehb2eGdOKX
d94rvWKskboX2rdSWfDxdqsldu/LVnucqUsKPwcUyeJX+ZT7fb2xbMerxLV5FhgAQEch7W7H/eFW
mNclBvRG/p2KASTBgkuAniX8k3YUvO3OyztJTk5e+dqDidOAgrucN+nTZnxlXlz5lIEm464BZ9OM
QeRM32UXpZ4MYFelmjiCbDXRolVgbIB2dnVDg091Dpy1fpPAqCuvGZhltDUuhSwuJ5HDYQE7Hn7W
BxETkxBWylKalUwzuJLOCni1B5AdQAuxMcgOc+daO4/89GAMxE3IY6dOdQFtULUuCryuB2ZOA6a8
Fe8O3cHXjwYf5aLWtOdy06Y0gKyojZJwCl6PwyR3IgWgivINM21b9bF4C5xTk2H5zooBMUHmv6+Y
uhnSj4Uhgbx7I9Qby9GavbQ/j7LFC9VKF+DAyS6yKUzushpL627K9XiuBBGacb60/6qSpdwfHyRs
qSlcvZ48Kuh7t/Mk7GBYzKqHAtFFxx/+PqDUhWisehaVbXudxe385r2rli7huH1EymDLtNl0jnJJ
jsk+06WQg4YnJ7tUCw+d5ocI1xJGDUDdiGwEaxSpn6Lo84JeDk7yP6hfDQZf9+sgB5UEqrneISqB
cA2W0oDifMW6WsLLmcjX5HQoBt2sAatEbAEOFGe8yTyVgZD7w0jQc3m9qbYNIquRwZn8LUnXh0LI
sjPn2PQW2a/9m6YhARzPC3rKtr6QKdq7eIKj+mowCnvDUJT5f4o23FcX2zAAfGA8iBz2lhbSbrI0
texkyYCZiFVtfOSQriU+Y7G3yje54yVIbgGGmrBIVI7AJlTUP48m0l/mdxViDcN50yDjphdrNtyP
QNUxSd7N/PCDaqbEVcN9B3Y2sIrO+L+9tlNUTZ90wGN4wBXhGF5BY48XUpFRB8rCjcrQ1nFgNnXi
gZWhRmBuIqIGELmStROStE86mdSfRkCSykH7O6ZBBCAQinwYC/8YKVGuqGR1OlELKmMp8q19IyjE
UqrNdlqE+BCDFdC5WdDjScCuHuppdJ+BIIbgyJt2FJbTPO344zXEJpjAksVAsW9vAy1jNznHSuTA
29BTe8jOWEJ+T2fY6NfBMv8L5som/zHYRFRRB71Ug+ZEVJ8fgwrkdWHezcN7r621el8p1Ih6CZ2B
EVIJTlczT30ueT8D9naT4t72uCtNQQn/qRK7ZSlSukVPBH/acraXMbKs0Sd/lnTLUq3P87TQViAX
bZPCYuASaU2Qdz4PTkb0tX9J+vppETj/6ZKf3q0XSspQsRVsNq8WaXOk13D8QRYVz0MeIA4HRkWY
xikXR7IeurLZYKyLlMtiqbsfOZsxyfbEJuEECvlxoHsJ1OSe4RGFaFTpZARPewFLRsEISBVh6r9C
6VqECH8uUJb72yjmKBvmQeGaMZ0bVKKfh6wpKgCSiofvyd+iF3JnUFW9KtRFUidjPcbkDQWu+fqW
kPinn3YbAOkm1NRurhfOOtM2GZGnxFK0YyVwmDinQAQdS21uqLWrtzTZKo6q65VvcEPr8Ywlnt3w
A/M95Nc5TZFFuNZymurNPh/DfUc2Wcq++xrnT8bziMrahMJmhSAD2EiSxjBjlvtceFIDpK2MVExF
7eXil4+CTaIg/YqPK8zVOt/uk1EzXBk2DPvJpBSiPK5TjXuU5AI2tSmlalyEjprUUVOWPAd0ZwGg
ONcmkM0AWQOrwWT9ySCEPAn/WSWBahTNXYyVFYqTso9Xy+VcVj/FIdIYLRc91To3JKDx50vP6gf4
/muWxC9BcEFcUm+4OutLaR/a4TEw2oQyOjCiyH43ix2NoFh0s2TJ2odRUwHudBdypZHy1x26vi19
6vdXvWY7N1DZauM54Rr857LXKqRtL60SJbugaRbs/kraOLZdHGCW1/kNYi11RE3xv+xRxm1baK76
av7BwB/cxXjb8zcHEoPCkLuM2W+GKxC6lUEEJPgcGsRL45tUivSGd3ktetbyL5YMJtbxELk3tYm4
gsY3F6/Knl++Pej35mbUK+Tf4a00CYvfhtqYeBlROdi/2KkJi31N26cKdCkRtG7LU/szuHyZP/Is
zXrDtyCjkmNam54tYn1yu5q4W9442O/iy6NGUdCMIyzF8nO7mTJIxAUszSI0F/XzRgv2ZTYGb6bh
OuNn5/Lzq6ti3VunfDhyhzYMhlpMoFiFjlSfZe+TuM5v9ITgKJ4rbc66Jvsd3mSCP+x47Z2W35MU
Rtqt6TdmlbbIiSp46/XGnP2igf643I6D5Kaq4lc+pPAQ7ctAjjVkftAmXgJB9vLTCvo3Pu7RJoMj
zCYMIlbTpryqm0EtxTYCOO4wTZS6mjgGocvoUkFOS5n4Slf+FGw4ss/OPNvs/4jqq3y+3fxlgvQm
eEvgRjdx7xGpTzphRyu8o6ZuujKUDaahhew8Xl9CSouRLZrN0F/KZql1hCeiNRgntzbQhX8lwy7O
VoTEhTPAKK8rzUSBalSf96IVDu/r1gtfUFB5lmWROmkm/SmMUWjtp5hXn77EwxumX4T84vAVOiwo
TENd/f+BwonZpXZjVdfTWTp1GNYmfippka0QR8GxHflhAQ4BPMgz9n4o8ps1B5acwlbNMkX1k6P7
m4YxRBo2a3SBZxk4eSPB29v4XCC6u4gvl1zqMAMHpeNGqIAqQWWSw/1x7u9OGAvfKfjHIiLFDBO4
PvnJMEgd1hR4SfW70mDR9LafhCN2nBxPKS+NJ1O/WOBi4e2lwJzRDLtpQUI2OdKm6dsbgFlk5vCb
XVyvzOASZP4M+GyKi4ZKFbnxR20KqabF/ppeXfPBt8i2KF3OJ72S3uFhDnB9o46qf/4Efc/71Iua
OqbG8PzsI2vSITO1px8P75YtMGohEU30zJANcnlAfpx4sMhmYu/IDygs1IUc7hJ+IBcZVWA3jURL
vNE9kIXjcTP5DoV9mokG41s9UNWpfG70ym3PN2k17cTOfy/B6+qQa1ZWnvqKtGl69IwhMHBoT0sK
w6RamlGpFnY2DvxVfV9hIsuJcVAe0Y+87aEwONwiZQp/tZtUdewRdANXI5Hviv5yA8JsxL6mNa2w
VXztquVt3pbNM13H+WB1z2LQpF13JeQnNG6/bD8Xlis+HDzi2Jl8aaiW/3DmRhod19HbwRIADuoD
fJ4oe1FjAkfnukUycazM3csuxgvcw7BIc8EK0Het1Efvwox7D7Jn7bi3lu6QZCc6PFxan3uzq6Jt
ZFpLr7hwk9Tu5XPe4I+7MJSn8mjguBcUPpNy2R2guyevPHpCnmva/bYndIrn2iposR3AzTvAX1qa
nBOgn8poTRzdoI6Pu+WEZrXGxz0d9GWMA2/una0XAWsMGc9ZjugXb0rTWUZtZd/1G6qFQgwC/D14
eaD86lJk5vUVqxtcaI+KYeu3QefjEwbSA5xSqrXDhgwUVUjXAHMWgAKsvQui/XQG10HS4+FHcV+B
XdRxVqE3J/xj0zx33Roxvun0DtGrxzP3N6m9ZfHI4TFNM72JUE+FFcFhA8bHV6XLOMgKWFXVgT+L
7ji9qWm/Zpx9WCm+8T/TNWKKgFV832cAyI2E0tE5SlUb9ZvYk33xZjEwSTpKKXhPXpEdwDAvQlPt
asN8avJ8DM0z5JrXv95sesc158eWJZS7Bm7naH2n/LAwSj3pEjK0BhI8wGmWZxM1dQzIlxchXtw3
wogjBnBx61CkTBWCtNexjyeSbRx23/SPcfNXwF6SwAdSJTGuLacosqWfq+hTIwpLrijX73u9fyBB
P+FzH2ciRPMwdCrTL/YKh9uEwVQO/mAkZ61/NC+QRM2Ty0a6gf3rDA/DpqVCTGQYyy9/zQ7Q5Un0
AMRnjfwd8UzzNPckNDjo+Dp8/9LEsJs0YylrXfF1n4efFT3O0pK/f1U3VdPaIp8PmIgNca/sbwwN
XcNOcnYh0i4AieAhX5yo6WMeEsdlaCmtjmEwRQQJAdOi20NZsf0E/3iLhTdH7NyvTapiA4wenuS/
WggReVQi3DFeZhtMu19W+WdVmTkocggutzANRwDIURAXYSLijSNqO9VPViSlSh1Na27z4mqB8x7C
CnRViPaZguAJ4aqsJSxd5s2eR91eRYM/FQ7jzMVXxqAawxypSwU25Kg0GXdQAAvcvbVLGq5xFRwo
VT0mvVs81Jc6hzWCjX25eXj0Kq1WKllxhsLmm7DGyEke4jHXc3cv6acbPLxoT8mEAu9HAplgp8iB
xpCDzenS6bOOcCRBG8mJ+eMJ+mN1Tx65crb5PC/OyM+oLMj/PksvVxCr+eCk/qbGpZxih0Q0s2ac
af1pw4P9gw5JlYkV9xkqpJPNx8si4NCzNEYwzQkGDeQqcqa0+mNY5ZwFep0pNJpSZXUAiT4avfok
JthpnstY8vr757WRleW/45fWIEoSS+RPBYMP3JZa8hl1Cp9uHtHOUArwZ11E6C47ee4tnxkUXXkG
W/uFkRtcYDGm5mNpIK/gzrwA/Z2XzE7RqyLz0OJqorGqJZMv67W4XJbSO/aEbxYa+st95ESYC+C5
fzQ45jo210kIxpqXIf1nJTptLE4GOxw25uUvYFYeKo/09GN50Lp3hH2wbLFfu8TPO8L6+pEFcDxp
qEZ5iwsPDfnJG6q5C6JBeqKKpOnzpVSJz4392LpT73f6M9fApsz8v7XHvuqeHxQS6kj0QKJepTtZ
5nd9/aKm1PUjnHJSz4xAsTWNrHg47avvppn+IoGp5hfL92GZhRLbbT1rV+bJbSOI5MJ4U6N5S7zm
mnvtdCifn0rfWvWvcllRcl32BcjQZkXAYKjpj42+JC9Xg3Fgp9ccN39i8znSLliTOpYxYFOuuuKI
RvavhpjHGno0tSkxCDDKSekzvhmBsXdK8UShk6tx4PAE3nixM1gFYWeSYWJmb3BUF/Cnrc+J9sMc
Xdg+cA43rgEWV82y6YGxfvSelWRKjbBo/CwzVQNkGpSjhu9zakKLKnTYiYPaj4WCpqK/1bNwlCiT
qlgEx5AOOODLVh+MADthgbxJD9TLVnf4wgRLFRg5kN/kFbQIez5jQUOUe+m9WEPnciRMZpG41FE1
GDNpZdsABZnxWZ8FFGs501Gpu53+WD6BFh8HjrI7pgwECQtQOJx8ICbQTBBSAQ+R9/MT29H8Y9Wl
JomhQ3/SqMrph1futVYQI1D5X0gECbulUmD0AEip5yoGgu7/MI+qflizUzaM1NsTbOkqB7f0OIWe
3X1miBbnqcqO36lsCy4QxlAV/zpYwtejKSCEmyETQIeSDAXofwuyZWu4OSx7QtM0e4hSBwFp3WXH
N3UT9ilQYkJofM+Vlwl80Wzg/UnMsaJC4T74nu70mQRcFXtt14eUmuo/1y6K3VP5BQdcQxW5djlQ
xH89lHbPcCEpQvEo0jN9tcWVZtKLPEdHJhkdq0fSixiBwT5pS5IQzSWQ5XMTTC+l5em3KE2InWgy
aRQegnFx/uRknGdtnmJiHwag3JZ4Nzz114+L0+uUcVlXM7H96KTD540qs5inTHvYPbPIiBdA+j5E
Q/DZ/GiARNd1CjL/UW7DClXapMTWLRw2M7uibUkxCdp20oiVHJniJ441nutZcTRlFGp0i+QQK/ZN
nmRiyW6Drp6Kpc/f/GCfSBe1yIxWL1NBo1bLu+TOFpcbVwigylfhKBlkrEr2zkp8iAo7q2/tiNCZ
SVWWUcFocKTj10Yo2h3qk8WoEuEkwtaCsLpeGS2fUKhTpYEOvvM57fmKhfeigmCspRbVclMxGJlG
zykGrxzwCS82k+uXv3d1ibEezFxcIAhs4IMfEYuri2WgrimNnZLhxKiRhATcZHZT1p1yz/cEFTLJ
Ns2iLecmC5foN9usZ3eI53EhQJ/Yfwrb+Ox7OjG75w70Lak4lHLPAgac2QNJ4VxMhNp9DuDIfjiW
4k9OYzUtR7HntOO+6p4UBA2iugwCiBGK3v3pBpCrILNYF/4DGpfy9TPNstoDv/G8C4AsCkZK5WjH
mKice37y15bQSV4UDmXkE1CzdAm3uTHUa3gbhYLbaXs9/BxfHuOJ9oh++OTF/jGixW+t4pCCpQ8F
eBD0U7cV/TNht7UHcjX0m/JUkc4+sXI5PFqodiJt6xlDePbEcL2KYRlybvC5NFROEXcAdctD+o0o
SL9nGXFA+oe4lGKcIP20TByIT2XcU4U4H80m9nUsgiu5QbXQdMaXUvSHEYbfFhuv+UaPkQW1qoMZ
Fxz93pCYZjOqpxpu0QP/b4D6hcWnhgYdPp6WxlRKQtFRhYNDaCmsehg+Ec5JjZKHccMM0ROpQ9+6
IeQt5UdGbq26SlU+3RtlB4nqgzYbjWVoCM2UNMIK6pPyRajRLfKuHfWmshDNfqRWBIGoGXgZybhW
/cClBADZxgIuoXGkmwVTYiaEPV8g1PJiPq4g2hniEpbvtdbKcRBmHMUHy+l4+VX/RjG/JgO4BLhf
DJ/pAgcnO+yNgy8x/6b3/gi/EiuxL86Ii3GWkHU6FruM1fPsxrwEOqWVcSrMiZxnuHU3ONx2i+0i
swCXEaYwc1c9frXbVN9NL+Ukyi/UMzESCXWDDvtJRjIzciUgC1MaK6d8BB4/Cvv7fKVjyic8L8Kd
PFO0x7+x2iywVhLgW3kRb1WhCXbE44s8yEwRbl4UO6ce7GHv0c2EQ6hCjEaTE0nS9o74a4j12/uX
VpDyQrX25VmcNJ4M/hR+g7a617lTfTNuB/itiYLL7JXiLeA9RJky+cB21j6nzFe3Q6wFQLrhASwG
reTaqX1Y0DMJlJllRRWzdWKcyrqLfHVWAgQcic1Ga2jJCEqboHA8VuGwOYSuBOFyxIbfvEvSZTaY
VZm9KY1ykBKDcDq4m8n5LZ7D68EJR1/v/vGgAqTvOLZisbHYl5MMuJa6bc31PtSfsp3aAGZSgDUZ
al5AmvXrJ6E8daBP9OKXZ5XPTz1EdMoycis9fxZHDboHGBJXVkaCqzJHoscNQNnCQ4YvDMbKYAOT
y/tasAXEegaCNp/H0zwdhWXJHNiSWmF8lDZ50BN8bYUM533+cnRVBmQzjCb6nCpWdj427eqcacAb
TMzNAL9NXzKjJIlV8LPm+wK2dnt1BdoY3wNZADi7fBFj8vK30mPGAg6zumuO/hxKdhd4Xf/RIsXu
djWekAqGnvGgpBHKHI+uWwhp+q0LXlHqzX8eSKJJPmbvNIF9uYttW9EvD2otsZTTfeE/dRThMkf5
51MfUWcEge6fFBoibFuqLcKQcDUgp2GVhsNyJRrsYpxE4uOtXFfn5G2zqqgUi4mGcSD9Vm8Op0uh
n8b6ZbZ21t2yC5qoskbocp8fipI/YZvoCZzM2rwIgcC5JylnN8AQyEtxes8U+fBJ5SM63ETm0SHx
g9Kl0cDzd2IBfUkOfDpd/7/F1hmeHPVfvCpm1c/S8LeCJXFMp1UdU5WJTWiWZyu5+FQWrGzOhvTf
X72RNnFYwi+c/bIoW4mmzJt0QFVgaEBkkgDle02PaHpgWvvpJ0P6l6fv0kA3Kdc01si8leP2au22
XVVizOUfPIUTi+gwymOheWEK66u31IObcA1RhI9DNQDL6E2T82bG8EnwAjUl/7g9Uon7k5gXCsH9
HVl0pfgSRiUqeIp5gSv7uzmXXkgJUxqZqr2gf7kfzYd+6xhOqbu5+eC+Th8y3s1sCWcyZnt3u4wh
DOeqIHdKvatDdmUezZV8VH1XlpsYXcSS5mLWnSo7oY+uZvirMZDDiCe4VUmWcpF/SMcAumE8id05
qhmu/WMJZY8EOgdq6Cv1Vc/4oFnI83Y1XX+wPTbZJg8lukBG1dIfUTj8h+H1TLHCq6pK9Wl4xQbb
GIBuM4FgYmL5B7g2tXSsdPDIMAjCNHrDNwu0SsaQJybmnn0ASNb/ErgfzRLFeB2Q14QJZfh949+2
MBLG5pn0VgqVZkDb5t62cFehInIhhdIk2oaydd3hvtoLKe1OU8R942YXJjisYnQFHjSpPN88mKhh
Q4E5jbiIx+1ounH0KfmIwyCIAcLx6CiqV9dwllTDED8lFoKxKne2IqrpvOvZcv7mwolVndW172a3
uNQK0UHBoBVTDQTLTZBpXAtDSBfLRn23Z4yuOoOtnHCr6YIfAlfBGoEjRoqMaM8N3AOAFG6DC3sc
tWsGBvxwa2857ARtb06FeIDIVaSd3Wy0B6PM8shPbr9mAQUPpWA5xTvXL/WXHEA7WDQEGC5CaEQq
8GPPqOmdLc5BfZdj2YXRluEpDLZpD25tOkSk+c1uahyCeTRdoZA1uJNE53x1/Q7YGmqUWe5NFg9K
U28H4Ge99pa4uQov9U7lXQOa9RKFRVr4n3eSdTgXnvdaFqFmm/cGZkq/eA+0MpUyIV6B+57nQMYZ
e3aiZbnOvH3EqdpAD10IZHHESubBmbJkDSlS8dHgXfxNLA5QuQPu+jGtmUMUN6AApj0hWN5wrEsV
21MuFCKOWIeDyAbGhrnz4r2i9aTVipPhBrD5zaLPb+gy+bLuM0XascTn6Od2By5AewDIlSJ0MUOd
XVYGPg9VrSP6qEahzbWpZWGj5oqugZ+nAfTf//Gd8yvDmy5VIaYMlxS2uMTktXC3QN9L6LRnD9EP
TH3rvJqg7GHMV4m1pno+gz42AhwR8TalKDGvwWI6YrzmpR4ZqFA+Ap7DXbGwYsvkiCMdJMUfNHE/
dci7QlRr4kL5hRoi9JtotSu4FdVHtsszBLCiNEDOoaPq1uRbun00A6xgAgaq7nr8en/4HwEAUPGG
SBe5PrqgUHje5scGpMfqMwXKb98Wq+TDwnqGYyd4FVHavtxjyzf9+Aejhl5EYbgyubnbs9q4V+3f
HmTcCE/kaW2W3bkbo7waQusOrvrrDo7dSKkLxWOC/H7PZx4kn4aA5OdAi1ci3F+k474m3QFjqdvI
LLD7WG6ai+63y+urgmnKhgWx2Z93UFNtY2EGBJExX8L+gzW4viBPyU+8B2qUtDF4gB0lb76gpYap
bjwyy6w8ZGBwO7O5Gjf9MnIl53ouUhICLAW9rykL293XZ6q8PR/XA4tf+xDgAuHKXzXp/M8UCiOl
dO2DdYxJBmWfYzKYcfA1PzvrdBYGRJr9cejQf9Tguim6rB3VM9w2bLkW+3B6ziQKQz+3DJaM8SkU
TADadJvnYWIo/azLXlYrzwUPG36XzUtksIlrBC5oPSZ5syrF1PwNJDHGlcvKflPzNuedAB5vPEhi
RoANoKMBL59eWn4edluAnlZS1ZXchVMrKIwZxV788wJqn6hiMzSokCdixUjOxwEkWfv63mJ5nYTp
XurmIjVMB87dLKu2syosV0zvKsXxgLQHIpoPh87oOxamDx8kYEjvVOzTbNYrwyC25bzKsoadeRsP
cxIUYVx+30CjtsVEcFU7BME/K8W3Jj8XTRhInyhJlkWIdlYaDSSSx06qFiLdgHaH7oQY4JQ/Mw8/
gkLyueCgcdt91TtQcVRX9RxnYzBKdVWrX6rVzOCm3tDOfyUyET3K9//G4SfYSkYlM6UIS2t6j2/W
eYIL4781hVJaJrYfE1Tl22Uape0FqUP07zqmWsa2XSs00ZcRbR7oQMB6rFc/d1ZaAQ7IMLTsZ9ww
f1AS8yB9Kcce47UhNxmMZZrBkcxfxAYDD7JYhPo5gUQPNYSkXoBoDmQNPt9JDfpg0Ihp+a6FEXhj
XTZXhmhtWA60bGM6yIyAlBhdqVa5AFLO7I5Jeq4yZELF2HQkeCYocCVT/cm62oX2eF5Ll+HnJOq/
NZYD17eV6R2/ujQAc4jiOA9R4KH90KIsG8dE8/gvqtlo+SWXSn09yOpwWT7eYKa8eqZJGzdmIqqw
1I3WhygzuKaBBYf/Pbta73bKxPVl72/pnB0d0ZPzqgNWPcdexl21Z1y1XYN0aUQ0XGlbFOJfI4ik
OKo2Bb1uvRtM7OXPnIUPON94zGWfvOdLiyx7L2uJB9COeJAifT8MnBKH+W4ZbC9J6fm51vlZkmxZ
9pqDoMaRBCA3bCjpEj+XwrJ409TCTr2aAVtoggCBAKt7PVHTcfNAh9ly1ynLUPGBHu9Uw48A8XDR
+ZAO6EnUD81eOcrKK2cidsqVCT2pNrE2iMsyfKSul+WgKjnbEfEgSy6j6ZbdN0pOTVR3XDxK16CB
D5kTJTuIZDxx4lEXxbWmFV8lUObMl7Gn405U0AIjqpp+LbdLgykpp+3+eaKFepQZsBGgtxgf3CzG
ywceswbEpWnURwEen9wk7PYYCLgfAadnlCt1SuWlAJ4n405IiR3/z+4JtgNZ2ts66id1TGBI7ORL
1poHkgM3EjBT7loH7EGRwh/6FbTSMCSDsbuP00K6slU+xXisWX0nwzSQwUdFP7oWlAeGDSDSYmMk
E1Fsb8lJeCLZ92NWYvEku23uWiEAvjjSO7CScpuO3XbJHQBGDENcJ5b1/fY8Jqf27ga3wyUalzTC
Yn8CtvTr1C5J/ZO718W3+3mLkUGwxqj0p7iYL8Y90l8VN9uEHmT+AtvKSNoLKWGUsuxOyKf742au
S0Krui/+dU2x0ITi486t0VKssTDzOsds4gH0NaU67zwN/04mFa3tI+UdvjG0iIClFBS761G9o+zm
Z32g+iRig2ToMJhc7HhnVwmpOB/fEZlbCCcB7RU2ItyQa4UjliqVoo8wLidV5W1WDm94xsKmafvM
5qivGLpmZZpoJPR2HN3Gfkk3O7urhpu8JGEile22G7Y2EqPVcOL2ZVwechDLHYgSRLoNTRDSyt6x
yEO3wlXm0E16dRoR/hImUxbNTzV2+dTvgOuMP9PZ1093BLOwQ/Wsxpt3U64AmJTQGtBHh2gnjZaY
V0pzQNnd+S5OQlL9GVOVrdhRIW37X1auKcE7lSDmQc2cdtAUWgvqfaketV61HBVbOznNKg+Qf8CM
hui+RPQ4xaOQcfqD3n/Wjb7dF+X5NpXy4zF/j3UMoiBDXFNMKouwqlSK6iEQFwCFYj/EYZHRyCvL
ZZuekx+bXg91QpSbVSR1MWLlqGjfwt+V809CNSonx7RHKKhUY1SFzvzArhjMR+aXT4WC0Q8ClZIU
ZvHSGJsTOVYomoWJWsZskvFixat2NiulSyuJoN4/vHoR5t5Zx0TjfRyfPep1jHgTxQ5V62ACzvRR
ST4J0JIPBtq2GpmMhvwa7xLQjXt8rkv6CgDymy/ibuLxlhRefhaU6Ecidnm7kIqPLTW2Sje60gWm
DYUOxUbkOAqPOLyv2hO0c/6Xl1VQLr3y69MTGftj+fTOGgVQ47ILx7BcD+XPFJ+2O9UcutPccOt4
pExzzydRh/0cjHmcMd2Y0F+YgkRblB8beiYqUcMtHakpLlS3FF1MALMHRnm3wEfg8UCHeHExKVMv
jhOjJZmJTmUDLqwx+mofdUwh/8Qnt9sZAaDlH9QrKzVMVNrYJLHZkEMc0hEKIJaZH1FEdzoJBDxi
Plif0PIjwxLiDctmhEvI83f3H5Encs5gPNxSIR55rYlSEpKZUc/jpaXFY7pG2hEGzw8jjgmy6Qxn
qAnVTLA5w65YsVbg7CBTkeAx2t3cdYkSQTOduNrlHmwUW/5i4EyK6Qls0asxGmJt9IAwZBjzcFz3
jjSRhjEL7oYcFa70I/ejvll+y6OcEU0fl6XXoOQAK9m+0LO7fah+r8HnOh1PmtPbX3NTMjJj7bx0
LKNVM43bov0Cc09Jq5yvOemeuYMHxS+qWhkmRDV1XHHf6hUFR/EdMyoTdERNbVlZRl5zYlOWi3RI
sgG8HlYPQWlnqQ4EEz3SRqsnGIvpkhboNPzAoCmlV7gkGksiagBQmbGyJfaqNNWSlPHR9WdQZ8U/
TNd0polGcx5XA01Lg+lvifpipe8Cm39Yc8DigLVWS5x5CP/Us9uok19VkDUzOKQIbC/99G5h/PgO
SO8F3WZUQsGecweqKEMlbbCu7biu5B+/t/2tKRYfkZt2Jvi1hYF+g46emrbgKrxRxceMMlLXJQbE
xHkNcDlHf+AOqd6/8pvARWqLiDY6vNVJv6Z5QDj9lCpmJnvWNazG4Y7uzBSltnkjNDunH8Sn9rHF
uu0002dDnE0ASG15qSrtILfXGyb0+4SkxIzQu1dUtyoIIMTzbOUteWn1a/KVwuMB2QSNLEa6jYcB
Ha6l/qLWxBx96woM5adCG7JHPq1Gso5EN+O80hWsHlRRtw6WeDPP8MNvgSCzUVyvPrkRWy0lY/Dt
/9thIIo+uGN7QFRI69hHiSMdsygyIy+Wd7vFRKmX8b+tJiDX/iYgU8wFD4lWSkTIa75Z48YKtKIA
vrp9wkHx9VEAwuORjyJFJYYnSIuSetr1pQh99YFFxFQbtzPtIgiLxVAiQr9Zhd3x1LXtqJ2/v/N7
smiUG3XP/9SxBn5k2NvoSzMgjdz6Kktur9vOYq4XqVjbonSwjoQuGOpoFhA1PL+JpdneW5hjMG3H
L9hbkLyqIykJcLfIy4/GfyZcu2IrXAourtLcIfCMJqxtMdjmsgG2OM+7ahieWl/kL5AImeEFUPVQ
sXhqFiyNYeh9gsia1NZICrrvtjyks8PciGEanp9QMjkfEnXb3XfE8qhlQ1HQ7q3HyKW620gcca9c
ZP7EAZAVHIuMdgRtuYVI5kEwLp1W8fcRanf3ZEQwf9S7x5JGVlGjBO2oqrfFzXmvAYUTNLEsIYi+
pWZzy97B1HVtWiUniFMNQLECgvGZSbkvrDCJJaS5X6WFK0hJFE6R8eIB7aI7E35FnL3k8Sv+puKi
DegN3mvSCVsXiCH7V2Td7HpFl+t2tyOaxO98zoNGNYZRlm6hKnRx9UXTiJSArEzqsCJ6TBUTeuGU
Ig8qraWzm5DwWq+0vtB6enWuO7H2UCMKlIZQcdJC5vox7pnH3Aa7oqLgKEdvaWmNp83lswqQoqzl
LtGp18CGJ8AEWh1cq6RHTs2U/Tiug0s9WWcuhGsruYWTaXMaWPfhNB0GO++6jZ2YkY84/N+MD/M2
wnVWdKPFO9iL6Ysksow5iZlO3LWzKeFcrfnQ9aTanWzexqPQTJ6oarBuU2xtvZuAkxEJtHUr2xsJ
Qmeo8TpGnxFbhm+F6q2N0xLuVz2wVdqAyNyAxjdGOqYXtAzlG9IafPQnVIK8uUWgEUze6mZjwqRe
07Uvy16Ht5JVqFIj25jPfv3gTcPX67aMGRvrA7DLaQS12feGLU49geHKrsi2Km0FSz9RwScVsaSw
VQ0eBpgbqbkA/Fxw7UNdyYWlFFmDjRRRJuczENaxYggYF8G5T6CpvhCy/aQbYb7UvyEjTgHwqYup
VzMDLAM90nFWjNW9gT6Op1up363rBRx9djq7T5NSh98FF6jIcBt3ou5PFCJdQxDNCc7uZ47mTIoh
sKY9sBQq6uTDKpn1P1ohKQnBh+HnbBtzf8gpb5aq4vf6VKR4sZp56d67AhZ3mTg7zrI5InwjKxMa
3BV2uZ3BuAxbpD3IzAETw0zz4MxQW0T6c9l3vzaMMYpQ3rzly7hXdCCWGklYn+66U6218pR0vnHS
h2/HhRsuO4CqHGAT1kIJqhd1M6koFN72WYV07jaZ4YK2cnDh7AObblhcKuw0DxPkNU14Zv5/9llW
+ktNULdr0YqPR1mZOgzxysA61YZaBcYWsrJ6ChQ7pb/wAdldaIsbxqt0wMn8xozdKHuHqVBnHqUw
Yu2o6nnV3wPWhNoKIc2xDPquHR5otTaZdKIJbkK8TANd3qeAtdRnlUIoVY/srykt3yE5XLlQZkQa
0OT9MWsDvWIO6IfJNkvsdoGLABhXM1cKJThmzLTkGo0ozxP5/ZHwjZ4Cr4PmlH5Hec9ujCwx16cG
Lf2W1hkoWtG8Ao58ivvP8ihGnABEyTqvAIMuZULVi44ccLUnevZcc1h/hbTThhF5ZOCNb8w1u9it
F7GfZJStsAku1w/WTqw6ypSNOw+W4mvJREIl/zmfjaq3fPHy75hzavhnQhZGczjSB2Q7qZsGUtSU
Tq/zaIQT0pZCx9+qvSBqgwRK2Q3DqdlpsVYfIydlav+jt+2jA6DUUoUD96GVtKk1DiWYG7JWHZuI
Z/SoDfJxndzTDcv1QQAxGuGTTwdo9ixqUSdFdjgu9m6nOBmHxXGp89oJqroVdk/iAzBC1qLpIa7o
9HQRgqOLjzp4GdIggb0SYFei+pilr8eIti8Pr3hFJ7TEJWXo8hE2phhwAMpmwbwUQ+BeeiTRjPmZ
vu8LID8WvcfjvIHww7IyIeMEihis2/vfSn8PZdBCcEwqkM2XNNNAyYtdu8YC3OQ95ynT4P3Lmg2n
PEOZFZehoEVgDwHQhxrazADgvDSW2E61ouki36H5MIAZHZzG2VHPzZb3Te9/R6C7SgHvCDU/8ViP
ldIptfwpw3dEMKyfL8pHIAc/SdY/BkNord9rzdpT5x6d9Euy3vIHvSnLavHgntB/LVNkKlZKh7H2
i3AeeGV5tOMkPRODFZ+6L8WGh+naP8tu9MJ3uvWeP5HHdhrTGj7tF1odYOJCdK5wsethirdSMKYQ
iLcRFnf77TMssyxSzft/zAoK2+flHnX8zVCL4XPCNDOWuANMCFfu4X99nlfg8AN2yQ89egthtNX9
XVwPCQYv0V/683O00DEcu8W9xeUtmTw4/2uw9KSiyMWjoIfTyOrkP6Zgirf2+nADLlT1L9Pbm/wy
6Yrz7j8NrtUgObnLo+8tkIvxUdsi5+pbUQXDVy1lLxpoDB5kEmYO3ul4CldF8KgW7NxPvtym1YoD
aLuRgwVoEguwIHkeN5Lv35sGaLRAwISUx7sd3Sdpq2rFTk5dpYwOImJFsnalgK5ny4JKBAUwdlOl
ee1Tifu+wR9gZEY2gbQ/scuyKkyn2X8rvP//1nGBfk6ov8Un2pf3MJ5Au5yOEQxn+bLPT6fIIPcj
ohSrAMV6JJrvuNcc0ZqzFlq8QNsTDQ5x1tGwMx17RwWgO6PIQiffjZkVH3Na6OMKc0ZXUew+nS93
CrtArfBiUAyd1ys7tT4rn0OcNteWcY6aeNu6h79oKJ2sGb10g3ADsBJHTZpcvNADkgWwNsUgpdt2
dgi3ctucruSIU+Ak6LA7kQ2MFGqMNblDQV+nLXhMnYUs/UggN41CdP6aEPDDSu7JCXcFTjchs43V
zS7wCsenn94SQXAt61bqU45Hz4AKjxi7SvEVB77l+iJLETfPSeAINDpxFch6DYduSt2uURWW15Fv
PuDTMKLBFnWuhEMvmKIgjRVnGFzlPIipdhIqGtwAbGmBpWj8IjAwvrYBARQOfQEpECgCa4Wpg+EH
AED4woAo0SvSvvyeUjkhEgwSQU+fwvQ3pNI0QR7vWF3TLy7MmOtSkdVJKFljurLBNH6FsG5TLM6U
/Y76ezUkTqhX7uiWmFxaJB/XsTpRB4sv/z3Uf1BOHrw1CBPppezfMgdf9Pz2uoeDtbAqvnYkBEcH
d8q+b8G3az4+zUiPBH1q6P3k5HNv9TjpQx7RAoQ6X82rCW3TkchdGaEylyLBTy6cFWu/Dwfb8DTF
LGzqLfhQGI3uS47s8SAy42rPCu4aSUORvo0KjtX8xvosISbYi4vNF9k7xhm1zzzRwYtMoAIz84hO
oz+ATrYv1J0l7fOJv1dTzVFhE+ZykXkd+lZf0HMxHylfFohy91LlfRTI5ShgPA/t00trMSKMBV6c
nrVg82Lekn1KL6tmfS6hliDrvVtLw0FMwamgWYohQfWt+eD3I37CYuluG3uz1qiis7OlIAaPCXus
EZ4G+7UunAYMYxg//x7U01SPbMg2fn8t+uV9Vjl6Jwg38y0GXFSSWtcK3M8HHc8qMemhyIKLKEGQ
hyeTFKzK3cI+O3zmqJqAJ5G43dcNncEskcPckL71JuDI3QzZtRpn7H1I+QQNSCxoYvCbi9/ZxL9x
aFiug4zrrUbZrMlzMBUp8Fn7pEBsnYdNbZyv0uof9EAbWOD+fHMeu494Tztm0rUv1NkpODVBTnOZ
KPV1B3/MEM5yqvmq5+JNwNE0is6d43YzPTmH2fdlrgWV6Jvh1uF7MgtcnBalvRJOs87juL2PKwk+
EJw6ZrSIXurKhdSyyM4SEFJNCQmCxa3KlCroSMfEzMN96hpg67LHP3SPReW81StTTuROdFIPo/If
CPsXjJVSdGk9kWA7yuoo134cKcDoM7AH0y9ZcQI2g+2e4fQM78ZC57W5rFVpkejniJ/w+/nUOlIL
q6w9bKRRcLz/Ewvc3/2wyJLlpKdTDPItFFgfUmS6p08V3ZWNN84IaqxR7fiHQa2dZ5tC4mKQv2tU
X9YJWFQHRzsBIOU4H9TmXbaopduw2zYqbARONQHFM7wSzRZC/seH3TMr1LXzO2n1jGEwSVMJ4qzj
koaasNE94nuXJSCoaZXr98Fqt7TN0TMkqPX/tubnb40T/OI1lG+e8taV4CDJvBD+vlwIdaOuyr46
lYWzZgivLNg0t3uKbE8gaNxfwSqqDx6gRM12i1MMfOXbs42ELsbvE0IBc+r7+INN3kw/WPVRnVm4
PVzH4collldBTJyW974Xx2y76jLGCqVeGbcGiscnkqR8Y/h86itrP18jLHIhCj5yaY/dhoRS0VCj
49+9AjYVlvbqk9EqvMyIqO72PH80DXlVc+f3Mq7SpJfzlrpuNuafcVZzpWw0D9X8Q2ewALsH5Bvz
zpGFnEUtdcx1WxW8T0ch3bVsc+Qe3hs3vJ1e9N7yoETuKmdTX21MNevqDJcg38ITuc9guFj4S9FR
lrpuo/O5DyXx9aVUNaAcfLRKVJM2aTUtr/ox9o8rfLnFHlNir+DtlSNEPebUORG0goN/45AyE+zz
JkczpP8MxU4yI+H8dz+XG5KLrQLQKvlwiFtq/9vlapojAl842lr6lygEJvCr4vII3nR3JWgcQmSJ
1p6C8wJwx5ie89AGqDhnbcGvUZXhV/7mxNs6sCWpicdq/p4FI1AlxmYw7h38sYGHuBatslRz6alD
qArFXv/yLNB4d1CIctl8BsCrFhWn2Nn1rz/tH7B+iY1TyYsk47gcbfDoyhtH7yK59L0IWfZC9Pu0
th+zpSkYlNwfoqlrpYD59aVK/Pu3QHHnKpf386DXlwuGqbNBJCyShDIV/4zescHLLUPYUqmNyCRs
I5CuYvr01Kd0qaf+y2eHYHi+V3BndsTVFUZt5l3iLlNFaTeBeggwLRQSrDj+RNK/hKqHv2vbtg/2
wIa+hSpfNgSk0rygzsxIKvN6QnawuvXRUe3AedOIVZoZrtUNC8djJ992h67vuNQYreSNXTe7Qsay
5x/HhU9MIdXblIrevi2hKGdJa6WGzWDpLdV/wiKaEXtGdrtUchgGJ3s8xgq7/soZyr8KuWZu7Obz
Y3yz6BnUpa3WFWHaTCnbGPWejhqEUf8mCOtF37MrTJboXS/qQP/mnVgNEGbdrmneTXIQqJIp7/Op
FmACcHBdBD1xEv01a33CupXSIEp4HwtXzhTWQz+QFDsP0IoUs8fcOonOfN6a5YPNS7Uv2UwFtWOC
6u5xpFx4YOH22nlSKVkrLswAxdmEYMmzlmDgLH+LJB0IufszZRsbBP8Gj1swGLoarDC3SXq2QbgK
pZsPXV9WdvXsxf0j6ICMct4GWEDeXAg7Vs+FN55t0grRhVHbP8pT64EX/ej1XPNOrfE1fGKdn8h0
xNjHUAYEMaWmwFhj3bMTBqoWVM/hWxkT57pEhQ5VkCbNTBiCii1Wyj5FYq3HOue5HQLcTawjM3Y4
XPYFEvCyRhEZqlf7gbSNL63uiSL0/XyR3vYIYV2JsoU3PcPZwys+WGAAX/5vybbkJD0BiRDfS/IY
7ZtyyLvyHc7ustHXeX8RHcV140e4QG7uGBew0iia0WXP5cgyJ+lyqaL84eRCWE21uXpWeiV1VxmW
HsSqdTmVhpKVCXLqXposbAHSPW/8Ws/OFC+8C6IJsPrIKYxE/aD3hhDrf06+xgxZKvcPmYdSnet/
DCVLWk8bFSp1V8m3IAHC/K9ZEAz51tNdPgmr3Zgx+4+OZmcVYw/2FJ3Z0rwjB61nWXR4muoUZPXo
45fPUVc/UGpgK/f4AlpO4lfIg1gc2GJKVbxQBrPgW6Z/d5FfGZkIF53sA+0tF+L8d5U9ds4UUDEC
PTQJFqdITJF1DasQsVKPRQ47rp1e8WToSOHNwKoTAyifkbxoIlp0wwgwvNiDk0HLGSKFAxFmxFnw
oj68eac7M6l3mQQ2FUdqIePSR+oBlX54Xjw/S9IQynLDAK2FjffD0iuH5xsd2bN4aF8v9ZexLmnx
35rblvIzjU5SR1WAmJM6+b70q4qIQwQAJCBwJ1lGwIqX0XxmIQMeCaVQqBhuF/I+E0g+y+nRXGbS
MMqDoNY1b/JuF1vjvwfFF6ht7rL3A5zvGh5vJX3UswSx0zTVwSM4bo/5z3bpJGiiK8FkF3Hh7fYq
SUnqrPJQOYvAzw1jKwkPkdk9pkAYf8dbQpFPQg27VmJlS+Zcl86kfA7sgKj/Kl/AlIN0GyHBl7pS
GXS2w/yEk+y0XvFnfVTlZnwN1QkypV+2bmycKaTexRfR4G1ftYjTpYyHMw33qNFNOlpvkDOoiNz/
H6E3BefNrE97xoJ2t+l+a6iMesrIrLS0S7W4AgR52sGaW0Zz1kJ0AQgag7i4N2CMtQrP7vqIW8kT
FzP6HqdTyfSsqFFaGUJuHCGsdHmUripEdweLOXE59RIW09QiMfiRjOUkbC8HzO7N0DP6UU/vNEjj
s0/HEyrKf+3sBMLopDR/nUBRoNV58D7Q1/ststHivWKzS2oxuQQ27mQwnRCdC4cObtxGtI0uJDUv
Lb8eu7+Ei9ioDHCq6niBSJdTrSerqZR7k2GBYKP2yIOnsd5YMyIzDCpx2XSw/odQpJX+hIjIGkYB
uoCrbwrPZNLWxNrY5879PzFTd1OVob470ipW+S7lPXdt8Hv872qBPNK/1pGufZt6OOeZ0/CgeAPp
3vh6zfkyt0IIUJmRuREb4mn9jbXkz2pj/QaguOV4dMS8wPQ7vXPD9ZXtlTvSnpbA1vkBFqmbjy9p
/hJFaLEOokqpFKJ9uw/vcNXeVTizegcHEfzEAKSmrDDmMzMq6MG9WhfZsQbT2CDdm6/YEBDzxbpp
HxCZerUxvam+Zi1E18ohED7qXmCdI6adiJVZzgQbRnYh2vtTdSNymqWKBZHl7vRessk1LL+U069G
7Q/tO7Lv1fGnfXxab3Mt77pA9ISGbg9G1bAFz2BR1NRNE1MiWN78TeOwFXAz4SE+EbrkutYtCEyb
UYgXxlD3KV4s9XXripyxUfpLYBPihUvs2bJBFgYuL1VgLt1hHEKX13YBr+5Vq6PG4CHgZd8m45Cu
fCD8+zE11HXHXdxtCnoW9DAkQ63jXocPHjuKnzgb0nztQj9nC23yA2NgmlkIT2JxhL40bywNofhU
hocdwrjfNDn8PPoy2FmfEDv+Zx/btvsq15gWIQ0vLo5/o1kNnbyujuWkiOzCjxhZxT+CUcOnhk8+
r3OulqzgOPTx0v1Rcsso/pvswhktdVNY8icOWK6GGA9XspZ/Yec2Ffxg0c7qelfVmupuXyZPd5Ct
lZYcIO3dEiY96CFG85A1Ia/Q49F3BEjD/5HZgbpdl85XgajSX7BhRe+7UfbN2CGwBf5u+v1RQjHN
iWpmqfXoTGS2UgVwiOIvYMz7XBG6weVZ00Yue2cQMaW8SsKut3nNRV8VPDBkrmExZ6nGTiszZOle
/tI5FYbHDQoBbFstRhWjC/bApb1RQyJbDNXwV6lBtwaq0eeZQYvLmd+sA8oBZCcU/R3S7gKBXRYN
Ggfg8D0u49c8kWIOBJSSmcN1/MXf/4xk9ZN8fHiKkX2+pjdUbQX8KQOfvtZBP7kpPZR8QF0V29Q8
FHSxiQVIdcIgoLnZKeR+ixKPV8f/ynX7vJ3JenCjO1gg5pRxSfiXMUz8IkcqT/GKcOzBVVEq0uKM
PxiXD+aGy62zDUwGcOow4TMzi+rEFubDNlaWniW1qHxt4y9Nom13imm5KuIwmhmlPVFCWBLlVZEu
YqGiaH/2qa2Oak4Lnpwjr7WGwEfCAiJ5l/OW9whM/TXWEgOCer8cMpvB8rE7DD6YuI1HJSKHcpnH
mZtrFU4+eUlWuA6mylD5RAZDN1slkx6KHwewCRg/eusCCGRjZ3qzDA14ndPD64epbTgKbyPyoHem
i4SYtag8sBFN6D/n8RfCPT1hb9SDL9IrV8YrXZUKvFKktZ2AzL89rhSpIB7eczI8yl8w1HjIrlJf
DZCXlxyx6RIEFrKPQtLy6ZvAXRWQZogbJkWGX0nAUW0esdukv9700lMwAzz7GuFSae3bPdwMDbG2
cDV3FhJzS/M+k9XCJyhj1znj60NRznj8dsbEBT8jIZNjFlQ5W5MrSnW/bgHs3v3OC1EyEvobthJb
I776/ZDcU+sDUI9ZHXc3CPjgbZb3PJfv/9lf0p50XSRUudnUttSGAZHjYrzvKBbKE7qG5WqOckiL
rMvANwCn8kb/52M0Co+x1SBhBIxzLSfej5ZUaKmzcNC9/QcWuvEDDivSBPbiGfZac786TdoZyRH3
f/48tSywWqwiflPcj94+eRCvntb0g9cmBH+F4h2egC556lHHI6jL58Z6BLQlJMi28eVPgz3BpU0B
mu3mPR1AmCLR+CMhfb5rQdLRkfyNqD2T79Pc42OlM82w2c7GmhYjwzTLdurD/BFgpfVwbRbE6V84
PtMIygdq2JFxAJ92jmkzbSdMy5elbQ3NPf9FMI0HDbJpjb5snqOYI6qyx48/aMYJbSXhni6Gehl8
hcNksIuxDjRrFaBnEjcBjQw7UeW+EyQz5v+TvvZdYlUmGdPNrf7/GUSXjc/s+KUXskBcL8SJtHnL
Tb1L470fKuCV/AgG3e8XmzHH+QzLsn/oVG4sHJfXXevoevHlsZR8LoHM44LbHKbGbvzVpbeQhCg+
JgRItLdKXlQIP5hbD9JjHIzS4aE9V3sUM1nPKTfaQwCP3stYtP4PBrf5jxi1D0FURXtv5sfTfRcx
6FfbDiJ1HuFDGJb8vNswqtuonqp8uTqclBYqHyhncS2jhaOSdZNpILadH8eZFeypVybWA9evd6VC
OGZa7ZnbYt6L50JaxHTFwwUVIDKmPZMxy3LP6tBm4nTGpa0Z8+HsNivt4M7JTwesxb9Dfr4pvIdd
1mKD2kGD5fZYpk0tZJ6XgyQTPTOibPZ6Kis/6mciaBHpzRHsuJdLbMTln+oIRKNBTEQo/3kTVe25
PJG0oljg9BDmp6TwjtVKZi6Qa0NokfegSJKEI+1nNUEGonTE959Vfs6hS3obZVls6/Cb3X172aPE
WB/9qmCsDzKVitlAGYRVVuks3z6kNhpWlB9cHrKlCLoEjYgzQLcWTqA7IZElgke5ujvVA7wsk7nR
NAFdTdbWsTPKW7KvIIeS9y4AobAe5YG6YTp9ozpWC5UxSiUGbmFAnp15BV1oY11AHlKTxwkO84rd
HTnoK0rtGlHf3WAflY0alDwzkaycVsuKML3oYtAlvNOd3cPnNFgKi5SajriHdyTcGKxfmwfnT7FZ
RCL/23hokNxI80xO6I4tnhWqXd80q+/yDPzMoRvHlsGXyVsKlqpAsQ9EqMUuVh8qkwnhYUZkGAui
nVCMsLySk/xX8Zp1mz2b1szsSrnLSG2zBfyLH6pPHLueyHoJyrOCj+X7DrpbScDCEeovwPviF1V/
scEbAIruWti446IreEV2XWpX5nek81+iQlWsuNZaL0rJUzn/eKn44oXGZM3Shz19+90ARaP3wifR
oDykY7H6aamjXY/kmDJGUzkXmi+nGFxwN9w3lyRnaOmTOL7qtZp3rP67obWfVx0mD9eSKQ3B6d2G
PAgyXn1ywW/V3DsvhewWX65+LQRkOwjIhHM756ySHo6WXHYk3MMc9lsL1WfGtcqdsrE4DuYg7Yvy
w4AlZ+bK1I+cEnH3zBp7xmOfzLHZ+52qdE45/tXAPuOV8rSlj1SG04NwhYMOYEOHxjD1LMnMBVoB
wTHt1bT7KUc2vCYPq4QJKNwDLvoA6L8kkQJBQ5cpOxFxFBUTRAxYIoiIzS9J2UM2P1DszrG/hkKF
lSCexNDgfF8HKmIaEEyEDNRBeAMT7Kesyti0iIV0Lo/Bcvml5I/KTAQHfUqeLBndcNBjKcL/a9g4
5rc2VlGcIyDfd4G8ZiXBbMPuTkANRQCd9gpLbWM9iAXmmzyNffXp1/jNEUTZjbmx5Ygq5aPX60dO
/FJxwCHiU8vy6X5MKW24o4AL+aMTK4SAsigqdCDjS6i+Xi/RAHSU7Xea/IW9LssYxb0QVsMZB3nw
+MMXPfTknP4y6xlwtG/F1AuE5zfv337DyEjfU5BQa3kFQNEPFENq/gUY3hvTziFv+YfX0mrhzMGj
JiOQB+xhyAOcBrf1RCLDTGpDO5QwWRtlhrNb4/nWbN89GJWehFVxrlFkyPzH6IscQjjqyqwcdstE
G4IMcucj3x8522wF/ToNofJWjytlH+GSIDwaz/feh48fMgGvk9Lv4ntpfqInQoMgQsE2R82Uvac6
wdMRRW293yniNwXlIK4Lp9aexD917e1L3+PGIj2z7c6JmPYx4lexa2aAwkbHYaVkROV2J+Hzm6OH
+RsJ2h8vWgktm2tkmd0hU/9fGcVbzF5zf9CM6RHNDe05s1aVorb31+LrCMoWjZvgWjkX+ngdUdqt
YajezVDMCISJG2B+qoEhkzjPbSm9zI6OA5IGm11fyW2DxoZ9Av6qQuKv1VHpIa1UXWURb1S27B9a
cN46Apd4wFsTomqdNjPZpXg3xVE0FFHf1DT60xvKqzV38AzT5bo98rZrMdQvQjYZPaJsEryVQ/7t
2oIKaFNHLYc6by9BjTI4h5PyCIjrV3CMWC+mXzaS0h5EYKucFKYXd5L/RGQaB620alMROTLLT2Al
4gVeTduZ1KbckuwGi5KxRSX/tUeKvAcAqavcf9o11coKdD4oMPAwsJh9zP15k6akNDaB62n3K5jQ
ZkMdCXKfE2LASxy3Wt8QQwXImt25YC17q8sY0eLuzb2SVPTq+C4ZDrCI16mwt2i1ksOLOrDDvpC8
/7qYQBHskFQFwxQkmDCuuqteVG2xU00fgK3lwbbPpNeik6N27ZA9SSeZz2UlgOuGHfgsIqB5qh4G
ao0x82TEmGLmRD33Vrt+R1jF8blHgSeMxvGDUl+ongeSKHFRPkDw6ZMbIjM7zjr3vc0h3e5pfs1+
VxSW9k6m26HOXpvq/uemw8V3UANJwWGMfrcPYBRpyJEyQT8EA0TSLCiIUXccjUz/P5nNJOYTN7OB
/Q74oJ8Ptt9yGiTxAjZWdgWIxFpmEqJb1HAaZpsmKa7Sl0blVFQu4i81kg+roW+9RqBPxKGns17Y
WeNvYxJ4oSBiZU+/JPe05ztvEJuIf1VZkWqdU3ttHpCUbjEpymGwXIolVZymew/KZrM84N3SFXfc
0bluxVcBI4DMcLsGQrId6G02CbCFUtB1/74VHXFgkXpSKhh2gyKFAkBXvjx1co4mk+F38UFpzAt5
abEqdmla6yjlBWGLLHGYazbh6fe+sOwbC3yju36fa9poF2NBRsBHrwrFy75cUpUiUrb9Bny9ejwW
4t18TdMMEWaYxe5Y6UNhiCr1r+DdDaQrK0i0TwDVVyUyx+MJNHQB+H/cyUua1gjLdJqhS/89sSkV
CBOen4kbe6/5aKD/jaTdcSD9SaozZoqgF66Z9i1YDvuz6J5jOM/Cyb7zwYxuyC3zfZWdZ9TdvMwX
V9CcQ97P2vCPG3RrVyWxz0iHVEp51sYWdtiMgrXIaW/tcvswes61hke0JfW1zz2VgL0tpkQFk5V6
xdCt32P7ObjiRTevoLsdRNjk1TcZ121lS3W6h4zzcath9n8BVczzsdc8Z/Hdk7RoirXhp9KmeSrn
MW4BOFSiD5HiKtapkTw0z0atzkEyv5debnJYVrgqg2F0rkrPb5rnamUSeltJ2LTYxZFMlzP7w9+H
+bFNF1SgtzUHbQqObpNzSmb7XeqEJnYgVU86XERi1o2AtpXOO/17qmurhIIhT7ABX4mm6mh2PmKN
FIlzZSPMTQJyrWQZFuXvHot0FNGHPl/dz9g9GBdo/2PUEYstAgVhrMohNu+I29GXOJMMTtvW/+bJ
kWQZK8sY/+mhaby0a1jGlCVG0ugEBSqxlFdJ5Qvm9CR0HwN14kXXAtnCTjJpA09Un3dyUKXhKdHK
o77T7yGO7rAsokz8tBhuPenk8ywWzweDbbxJgp0TaI27jwrsqldNmzATrP6IfIYXW5jqFiNWRCMT
MfOSuwVHFFtiB6Fn66RIwcQk/oj91UTjC0YZ0NR/8c443g0pQHzat2vCLSaMiOM6r7MPlHDKP++h
VlCf5Ri0Nuv2X50G4x3suAotz33Rb4TyKNDu2bAHt2AsQwOfQulz61sI3B5l3/ga9XutFDJFBMtg
g7GbaLNXw0FDlsTitYyH9+24SUediHAOeox4kaCH3Cy5ckcN62NGBo8uq0dyGVJ90t5bAD1xNguN
w1GzJiW873vSamJuvsf8ArxtQqaWt891gPN9IKSXztfvcy6pl9OrijYLcugh7VrexcvMtNs3EoHJ
bhZK9/DlRYbMuZgDDVAa0r/lRw+b6Djxp42loJpMRQ1esi1HSNwy6OKooOP2fhnBElxdLlu9hVsh
HJrIF/bCqzbhHZ/XFBZNvXXg4UJITPiCGg9f8I54ztmtxuAA5qfXm5d617qqgPlo+UkBbbGZ5c6A
wO051XMmOpAZoCX1UIoDwUiJMo2TfRSr7V9EJnLB/q9zNuqyWDajkvsEKhP7oEh9bfCyptJbLxbW
UlggJFwfuZ6YO0/yxesyMivMJcYxIHBktoJQON24MXKPuoHTSN+fv5IG4VLekoB60IxsxKBU2EgC
a4VjuoY5Zyp2GnGBo/S8FrpIq+RSD5Zs/wC9fi4C2eWkYutUWXR9sCHnVQAd8IiLA6rJNNLKMAkt
GjqXndhpc4t41fRH9P2YqxjL9VEGpWDO5uDP90g3QzWkbIA54ruq1NtVdC//adK+I6IJ0GZ2c9RK
nC2jI8QEG7nXakrlDPlV+oix+uGR7Idv14JNTo+Jx7OHOw/pgwFT+FHaSioFAUq5Yzypkh6Tgd6f
HnO55Gx2pu0TEksPcO61IpBYxhXkO/eZyWbywneGaN5iSfDBOmuDLxPk1TxWzsaIakmLoqx6TuUb
jV0OPsFkcBFYIP2+MDTMC7aj4pt+SSdpUWUfs/qluJ/wRJ9JbC2EgsYc2vWV9L5eyn9wNu6LJlfj
vAe2tRHzWttqDzpvyxrWh18hVPPqw0T1uHj5pYK7mJ+qsgIVOzVVV5LAf3VKpfUga9LFA/qaERyJ
3e1wrucCE1QWQqA0/s5kL856CTzegRYGBFfCLgDFl7vFHznHwWUzeuNYNcfSWvr5T0Gn20jrSOdR
cznD9fcF8CPDa/ptKpYmD55L/IGEA+XLTM4hD/728HDw8zIzFRd9YANTSB8Ra+TXw+AxUMDzMt1O
qQT+2PCCwsf+Ct3hlZ5sVAM5n7Z+BN4f6F2GGR5/iM2yio/GqM3Pyb4HJDV/w+uJ4WaRWqReGjHY
+XuaKXEFpO/xNHouKxvDVQLcZuO2QYYghNGAC5qdQfvglusS5HiCfWyLuVfqoZoXJNCSQkDsYMpo
VGx52MIniukyCkI952iO1eXWCB9t2tbQ7EErZ/FsYgOuW2AkFLRp5ibe2hF9K0AQAYGkNOjj5lqh
8OkagJPgzFQYnFVtH6EEoRe3mxs6aW/tzkGhehcszjrtWOGGAd/NNMr07wLBdxiyEj2xUboFVTRR
Z44mReNoBi6Iw37eR4b+JUTF1dW1nSPdMYB3TkkkHJCW7kMd2JUHHdnnaFmdjZqb9N3xYyYmP5dM
7swAnaQ064ydok6Js2w2pnJsNkS4hCUqp0cSCeT5Bt4/fsZdrfqFuBhVa9graz5/428AlRJTU+f1
z0ZMBoUuA2q6LymRncSJ147aswZY75s9S42ez+MPrbeTdss8lJWbtTnQ3Oi3+n9+Ju2Wm0imcbuA
W1EROF07QgwIQFvHcn10PhfH4hhJLb3xO66AsNnVIJtnD3sT36/9nL+JxyNXeZ1Bs76ZTc+jtBO1
Vrjbuw5qkgpSWAVIjcy0V9/Rk8lISCSHBJc1nd/Vw3YQUPB5e6JECW0176crQBYANQYOzmAOsr8E
LgL3zVZP5nIoNbP3X/PtGGWRYv4H+jYtH8Fcz5JMtlTzldnT32O9bcVCmfCrSWn0QBvrDAUctxi4
boU12qy63luax2LuiLDvzZ92BeXJuyqsexQsO3zafhtJX7I/lwUVRuRdWn3dxBQfbAb4hN8C+uwh
Ir/UCVJFn+4pRy53E5XcjXicoyiSE7XvUOwSNl+zIiuF1Uo4UTIxfi6jj7G3gGu2H8bIXoPolU+3
y6wvW0glYIHYxxkg3NGth5wWIeGl7vAWaJf0Cc7+joVGKZegboJMfKbOvO7tIqSWTdJoPhRcdkgR
houhYLVsnpnikD8YU+/EP8OeMLOnNL8mXQjAoAN+mTVfJRvhhKEfuZtTcCWwM6UBPn7Difh7CbKj
Trx7jVD7uPDf1r8f+OdUXeuHQqU1W6+MC/Vypoea1E+AUH7oEE+o+btnrRr9oA3fHbbHBD6LRi6F
bq3Ji055VgjUZqR3Ycy0hsjwa0jHo+8PReG0CLfuR74QD1kznmrICMgJiPpMl0vrMupZJErB/EEz
FkctPwRyGyUS84Js9ALx1me5ruAt/xmbVI8mjRwAjHgaG0oCcrJt7LLvCAWKgBGJU6SlUETZZu8T
t1pfxhBfSbdq2viDSoicoiI/bBIVz5DJWipiqlnjdBbdZ55EY4dL3W0UfL59UiwkRR9zsP7KHzUS
9NYk5nhh44+IvYAgLf86lMlG1qN42epsjhGO2owj0znmOEZxKyoQewgCK4zAphOtbJ/LhJNcekSe
7p7WfvnQ+SZiUBhPzNN5vN7Ols4Yyr/Z+QTfo78SELQXWbsquTlAGaHe9bqyHkdc6CivNAR0lVk5
pMfvnkEjMN7V/0oa/KAr5/GAhg/2Rc4x+tGoU3rqAe58wlMYf9gVrAZrRXTDiBBdXQmOrL27Rr5L
HbFwDB6T1rseJTkK+zPxJaA0WJmPfPKjiWyjMhy+9n5VbWbfCeHqblnemn0wnJeFsij4zhDSUp4l
es5oAAU/LlbsklpVHYgzEf+hPB+WYeOsWMb+c7F0TcqpuofvaJUClveQCB8WwUDRboesOSAE63Rw
t38p/ZpCHKmd90mojZU577BE4+5jCoyMKAceHf5dYcLO5FxnXhNo9uyNf0K7UHtieLFAOTGhh4Wi
DPOoFSfOnXc3cNRwWD0Rb+qNjkQ/dYhSb7RUiKltSbGC3N60I/xhCsIOhFX3+CWO6JgDSS4A8ZES
aOcd6gvtzuR7o/Vj4XY/QaPkYftOMag7bYE6QCdcdYJjYWwFWg4K0bFs6J8tK6XjBlqYVDRvK3he
GB1M8/F5cVKp5kJdHDQ3FqhUCBWRX3Rv7CKUZs3cBngITLe1CPQQbz8cEElncfv8Gl/Cgmdda7+n
LHRKv59KyHU1SGNbXxWuALuwrUCWBDgAvpIlYYYKv6AecijsZVQJrHGsZujfvP/HLOrXufnVhnIk
YcMH3SfGrAdspGk7I/c0cSittss0oKzum+PokELbyCtb+RbL4smP4Y5VsGcWacVEtRUSByesix/F
Q/rPGY/QvQvPSCsGe8gv0zmZgMsvrWxCFhUcLb4+YF66hIrsDg+N5cP6rWAo6i38O6oJbK0ytI4K
U0wjLpU6/BFxbBJnW2OON/q7tLxzWBx6Hj1KPxD9ATX/FtC9rYtd2ylNvSKxCDJC0/6HnWksRCjm
6toI17UQTBzItuVFRiBKRgJd3tE5r925+w3gDMJ5hIHpwDa4xSHNRZWv0Y6MUDjQxCD4BMzo5Wd2
Z24TcYzGG5Ln+7VwOuL08bKvb/kBGy3ueqZNq1DlG+PjYLn0zmSNTvEqinGpFBDROBht9Ym8BwRl
RWZyVoO9cW2l7H7RTFcdYrOicQX73JLvYrqeBiZWBzu2APIUD1pr2ahVRBaugAWDdz7FUi6K4H85
nfueK7j+Xdua4uxPMirozC8HY66612GbXU6rrhezuDa4j9G5lWFiXqyLPrg5n8BlDPHmd0XCAALF
Pym7u1LklZU8v6MFFp92BKrzNIoU72Lryc5widmuuFOAfnaBzhUy0cm3aEs73tMPJZN1rBdCbalD
6bgPR4Wmce9SXPYNmuw3xYBewqq1UUrm0nbUINU56TXVEQoMHhm96wlV1XMwA35TOZgzcw3EEGf3
lCgevMWEZG4seXQgRs7uhMqlEYpnYCjDgtcvDarIgknyJEef9zd4XIOYkCxkJ03cSixmpO2qI/l/
d3L7qV6o4CowTXilsl/d3ojpjLhKlM+YC1in/lnPFT6ApVPGHysO79uDamAO8DQvclmfvtlJUy1d
XR3d6evTPXJW5CqrvSjwyVAIZfb/L3AsSWY9f+kn1fpHHMpT/EaibaX9vYJ7biY9pe3lWAOoxzZ/
sscis2YheAQPUf3iGspg5Q3ls3v04vxWESK1I59UxgmzN+yXBHiK5L/UlnU6IBPp9xqEZIx9hGIe
saD/2ge5TdJ35aymZ1Bm9vRT0gfyBVbtsjnhtW+p3SltVsumhgkvPgw767pM3W9W0E6FJ2yKourC
pHGzOvT1pmpPIrUXDIuyTvQmIkSRCGpF4ZSn9UQmbZXgrf7D3Sdy8LlvbFEbILxJ+aJCbgJ91OIa
viYeC+PfqcUjRCIqPrVmPJdqRhPg9giSWEsd135c0jJSgW7ImOEazQKx8THjJwpo5FRZAGT54BKl
vHECwcMpK0Kh3e+gzGwRlFq/kuk8d8Y/r9R+kd9xLcYLmWwdsrOwXQp4CbCy54+U91v55gF4cM3O
/vxPVeuym+7qHkKzi4TvzsRo++tWcQJ6ZKs74PTJmBVSCoTwa79NGe74Zv05mwiz8TmB5UMQe8Dn
JOJaKvIcS4LT5uv909QY6Kfm+ry2fVb9ImczDSZFEybj4ZaRDcZgIoaO5GuIdUhQRShT2mqRkuRP
MaF1vg2yGY0JJn/m5ivIpJpMHX+zepMOKciUJcVdVMb2zakTPTKsGEz8ZNRiZBPcHK502C4QcZQc
TtzNy+wlLc5bt5WPv0Tknfls/DQMSy7VusuMxx2N5uHlxZC0W+SVWSFaoJKwNv2VZqV0zy9xXdNe
LizAaUWg7YIwwCg6h6303mXgmYAEMfsWG8EIdII2T7dGHRkvft7e7tapjRPL0UQORue0exgtvXiD
bKylPeNF7LCKLPmOJ8KUquHl4lTCdWSfR1Y0r874pFkWrCBgf5v9EBueihTcSbVe1+n9vnpj9gNj
nr///xO+kS+iyvAUivdxtv5DBRevscrUPXHV5GB48f//VbYweOpKDJJIuOcsNOg2wMYySDlcGhBC
KwsBiW0YVG8MIKM/tnHpi2AlstaGu9krcb6VVS3Nah+0O2Xa0CjbR63bsbsXjznTvdTpe49/KqMe
8CG6ImedZczOuWr9JbfpSU2ppYp+ayG9081ej9RRdZw54ucRC3rgmbfqMwXA7QOPrLEy2X4L+v+w
UpoOMcy34Ml7NMveVrH1W+ThdrEqdwDEPkE3y8rLRm2LP1LTmDa5kiTimf0G5Yb6Vswu2BTcNPlf
x0I8CjGEqLAB8trSPayYpmTczAHSNkXgK9zZ4t2H1kTQ0DsgrvjzpAA/97sishr6D2sJ7BCzbpY5
IgTCcJvBvBXYv4GZCqo2J69s2Fz4ULaL+sHsm2iVjhaHt0lVr8JXFquHs2qaeyRMotPkIQO1LDXT
WBFkmdlz/jqOa1Eipj9zq9BrEB7hNiKzvSMLpYRNeQ0U8fIhCItRWlQDaX+eBuIR+F7NJZpHtjep
jPEARat1iMg/416R2frmA+geGWkgBgTO18c4wHYNjgFjU3LNFd6kGUDQ0QtR9s3n3bagwi556NDk
HSB4OP/k92ChLOttMP7XTR5azxvcWTVoHxqpnGyqjzMEpo3gmf6cZtufGXNfnUoaH/0YDXDZJId+
Vf4PHnWj6ZaFPh9E4e6BF/yAuKwY7ZskwrJQdzXAxL4RwTGFVCHKjKdxcIVDkbue2FabRiLmVFbc
wLKSuYVSmDVSKqDgu5bUKtNTnA3y6y0kvNAzuM00yCWt2EIY6xT7ei1YyW70be4DW4BZ7dz1+sUV
2oa8D6dxGOqW/HNp7s0fmaNABEyGjtFSDUWq/2mM7CKopqN5BE8KuituOrh2srF0fy16THTaGRND
i2f//MnOKRhHjalFbvnwDPf3TJvwuqwkhusTJHXIBhsq7/Qf7CHuwuaW6edXAKFHj7wadtg3byZe
Lrd5A9ENZWL2wuUMLlUtBBi1/GIrIxDFjFAC6kkV4wvM12MDMkU7Ahi8twHD++Hz/ggDSVNE7CK+
YZ//EjEPsezEFdj740HG1kzf4t6DifzKO2uPmiOkOqD8Jfw5FOAll8fQ8/I16swaqa1uns/ram7w
OHoB/DUZXKlfElISikbcpHbV5NLARfgFJ0+jctdb8E07pKejzurfhstg9affSA1dDuQ0C7SI6T9U
q1ZHb/MDs0PjMYtwiCeEOz6YQ15l9CoevCK8ENnexKZgg5oxLZrSL4WXUADYGAUSo/vGsSI2+I2P
Skc6iy8ewZZbr4mkLvleKvsdrGjVCdNYMByndEtUTj7gjetMQMMfYGbFZdPt1rL2V3twaAXDoEKG
21P/Q6tyRB+s6k8ln4qNLHucNdsjiBpZ7zNpTiiZl+77VChzQb6u39ad8mHjzWXDeX2iUIoEdgBo
2JCvT5HXt4i4SpDjUyFN4GG9j1qylnnsNhpBcqMKJtS8srs13RRG+dLa9kArlWnaejPxQSyPNbil
1tfgMQnLGjGarTWMKh0YVz+eAEUzCI/OzCM9c2PXrAmXp5KP7UFdvk3C0tAo0ztSVruSk+Ai9XKf
DhxJbhaeK6ObeAfIdkCDhsAq4FR2e1O4fc5gCX0Jr/svG9twopIp2ARR/ckaUOoye6ppP1SPQyDp
NYNNj8XNjxhRzIikWJLwLx+ReddUS1J2ibgDNOubYpfGkJwuxWZBIAxaYNXnORf+dFZmNxlr+LgZ
Ap3S2RQUzuitTJSbbhXj2r8hVa4SGrIOeL/oqwG1rYczamVdsSa7gi0afMvsKXebGKnVSP136m1r
w3bXL9K25kYUTpx60o4Om+yv0l+hy5x0rvD8sNgwvN0Frvw1f3vELNoa6F84TutLa9T/11WiSkGg
PhpsggLaiTEfcKPjGBYvN7iUdN3gGYPpZ3UqmXkzF7PYCoSTcxt28qA+x4qoeMjJmSxVx+3i6v34
tn7uQtazOwqz7J28qEJltI9hHijABT5BZsj/IzWdLThtC9pVQNwFqCuhUb2aWiMZLlJH3fF3Y2Fv
X6JDJTIEzq/5cdvebu1qDRWXBaLnFyrgKHNN3ymbkNuRgLnPc40wRNaDf7L9AouPRM6Qvti+Qbfz
NIRsfEQmmMfSFDfpVC/kFJJR+yquWnm6zd31z5l2AC1vE8p/pYya5X9DSZtBRKI2T4g/CZmWxe9M
ZttZQY3tXYfcNww5eSz4y8DoztrIhbHBiaQKW2dQI4IylAVgawKulfSXzP4PVZELv/knbcDWYovg
QYdZntmIw6XrayaZUk/YB/7TqjZr11DM+8PSR41l69y1P4qKN9sCtvSDnnakqt2EkWiCpqH4jsKK
eUpsd4FxT61RWWaH2/bmU3/L+g7xIoIaQ/oVM9FsmsHqWmSo+9LL+GYN49JS1y/P1uqVrurSJFRV
VisBJLmmWLmL1bqYf0jqBS0ZUM7JEWuXyCyQT609ZUKumwS6h02WbqmHS6Wpy16a9lUla35OSlla
UAa1vFJRQtRyb3akvvvm1XVh98ubPWRDYMqEtOunduEMI7UYM2NiWSenOvbYNwMt9kcrNTamdJEo
1RoMMM1HXwRxlHxG+Jg5wA5Xk1AG/moahuM6QNssqXVqUUFfDMssrja8qCoFMXqNtraHLQrBqUyg
KRdUoN8vQBDP2+Qjig9hjak8BXcy6zmbaWc42oP9YrHA3c7YO3BfSRQAGSEadw7Y562nIWlH1h9L
w4HWFXyuwHICNpOYhQHT3k0wFz5qy+zt7VzGs/eKfBXyQ6VKcvEvBt9IgL2lBW30MNclV68VvXaR
/yuaNO7MqFaKOy7GtHuT6Xud3fbTZWvKvh1dZSLKcpNfJcrfQOT81s6GaTx7E4qF+He8Sg23qFBx
kqNPkMpYDR5sI2JjkPV7xyjJyKwdZTDDNXotwXci81A6IZewAydRAopAAcMu4siLHyYsQb9xmxNS
kxMPkTCqBxcfu+42l6a2TWRK6O+fFBmbqCgT/IytNUVZNrYmg1/RJhx4K+CJ+3uXODnwFszRAKK/
PC5EmpWHPMUiBmPGb4HOhYZoxeAmuEfWlaFGln3/1AvL4mdCM5LcMOQq/QF+U2T69jsFj0PV/fCG
1Rjr25+b+dz4cqXe7KYnocRFAR8aV+WpoScTpx9S6+McTJ0YEUpuXlLLbJV6gD9Ba9AzAN/Sm1zE
c2C5Fjedb/42Y+C/Dtjz3tEayOdT/jycKf6o2O7zwT9gtbfhmI+BF6bleOqAsQQi0tM2tcnvJc6i
tMeKKRI6RubN3xczfCTqWjVKMzSBB0iQeM/8nvqJDycmBXGcP5phz7evya90OdPOdlx7QNF/J1fg
8JT9pQh58feB/WMlZwDI4VEJ0Secb6YQhFbv/ull/mA2KIU02MmWkk+WaehyB8CNNgb6e199zU9P
iIvqrEgjKXWi9574TjdkswQMx6GA4m8CnFH2iKVgC2gHPJ5D3ydPYuwmTQHhMF2eP8SF8PWUWjIT
AOR1dmDlEt8OeNKajMw0zRAwqu0mHdc5T1ZHMzqH62h+W+Me+kYTdwq/voXAE+l8ecQqqNYkhmt7
Z5c1qAM0/kNkoyWMGpikMdiNaUgjm5CRpzIHMhmuH44TUe6mBMZVS1uCNooHK+97VzLiq8YQNTzr
f8cJb0T9EMCu7b/kWSgB/MopuR1XPIy5zs434gx1s+DhDJbvQxaiSiWpONZFLG4u2vwKDV+nRfUu
4i9ClIl+2LoBwQvEWqrn0RG6mNG6E6FygNjTuCEekVLbRvuXY/Hsx02rik9hJfLVxaqzYh6LYfwu
xq+F+4Yo2sBWc99I1fypWyX6ivRC1FT9D4bcjmKJgZyWbMYkq6HZqS9WrOM06OrS7KiaQzc4lYuO
HfzXMnTkEbn9Un5jY/+rPE4Wz2egWIl9V5IA7mP7FHxPaPfGBxFSfYlw43+6+clyRV/Uri9fXYah
zV1EBFXGzPOU9qPinNWlxLIU9n4OcWRTkSrUMINceS+mvPoXTPAhP7VNaFEk8v4ogVsN4dJEPVgL
JfWd3yNH2T4UIJ0HNUXYOuRB5NtOxJA1H1naLANtjv0PWoTxY+gunv0WRJZkXYPxAaCfXYGrZp6t
Dv4Adr1KSPHS4BzrPvtP+AgR3M5iq7JwFpFOziEyyuB8hQMvri3NJkM8pyhIC0ukqIJ6rIeut0EX
EBGU4ip8O5KGBfZd0TXVI93VbKPwnb3DdLsljjX6UPQQ3YiRs6aNTWIm2pK8FcxJ4WPtFXQZ2q7w
Y79t1kKteuF2rxqexoJc1IRTMvQhy5+FohN2yO1guWwbaRzA787nQ6HOfTimFy1SRrRBJgA13DXu
fCpUYbVHgD0gwq+LlziqaH5RdHTY2gkfen5g/MjOM6nUecqMyEC6u+5JHVloMd3V/6FzleHz7kYb
nZzvyb4tFtFJPBrsE9GpFHTnqZ4w+Xqay7OkTZyNNqHs9GK3u/hcQunHVcPufBrqGuZbR8+B5L4Z
VVHm/1OcvfAzylqk7KCw0O92BQFmTjqJdhuneQR8qAA9D3OmSUBT3/Cmy4C2c4n5BrZniwGIW0o9
TAabr+HNMSrrneRZZO6iw4OCa+JJjtQ7mdSECIGxNgyFZNJvonskfUPb+YnBmfeYv2Rqm4PnlbIc
3qckJ6dug1ngbLCHXvAJ9Tri9tVT/R8MwfxZ4OTHp2rwBNIDXkH3oj0QpkT8MCzASLL8TvkERybs
Pz85CbxfhrwbxO7Ey2zI0UkocDfmL1W+4dxRfWe5ETYgc3clDARUvfB/8/ETicB+g4puz/bBksRO
AW1LRNJ1VM9Bt1leF61taKFvVksVeZQgAMkubFko5GQGQBcmuITVP8Xr54f5mDAplta6Du7tZfrv
WhOVKf02fNFDEk3Yu3vfQMUG10c9iM21zWCAHvhNEKTo6d+BYtb4/O1Kx67EMGpPrW1ZTcHivjnA
rk4PPISwxwZePX7r1unF6i1d1c3Qulp/pH+78Cksh73d9FRgxpAXX6EiX2K+Al9S4iFDV9O5hqQ9
2qWUNdLrFbHgmgAw3KGNqaUbSQy3Htpe/mp80bE8MeHYOPA3v6zY06eWbILPTy0GsQd+ubx+OZnj
2qggcyqQVxmPFJZfcun8SPJZnX/fQi/ibm8M1IRaMp+sMpUpkeyOMRcA2m30E9Nx0joLpDBnYtZ8
o7RiClrkkWtZ9hUJbwL6vPhY6fsPaSpUlWnmJrp0MrYU41SlvGplmbtX6DOIeAfvku4G4/aHOTts
4hYJGjsYseNvI3xzEjlWxnPdQym1GD9gN51beK82SdzBdvYwtTULzhyHFCCryYFfZdfi6Ya651Wh
DRKLfzaqjYjoQ2uQmkMcmKTp9KV75Ukp8XxsCUmCXmZTteUkeAnfnnaxBSiEzHIq2dV80mMVbJyz
gxb3SnVjgIncSp0DEggzxK+87EC6RkoKZtNJKBRmaLk1jSoBI4pwdNxswiIr7km6T2+7yAI5Uk1l
uf1Qcb6BgswOUJUY6HtWUj/hU4vSczeAsyTq69TFSTdAAHcRrfhmiJB5vPZWgk2+nXB12cSgUlZQ
OAL1rz8m4vkH/GbjiCn3rRM2LOpgSNbd2bPQ3uPpCo7h0gQ3NJm044d8NPt1zRhR/3iZtGaOd1LY
V4ajyoiiiQg4gWIC8LVpuIBH09fuJwlhfkDLx7zLDpvWM5P30fHM7wwNsU+Td8S4XjFjckLYj2mI
exK5KsNJsrwXGpw3pSwx3vlu7Yjsw+WcPav580RUc9PEVhLBmA4uEEkl+fFLi4YSh0B/CBDuW59Z
MuwUMonEAJXyGB1DtHxpRMEVkMwOgpumC8fvtOsWrqr14u1beHSwycuPZgL+lFlECdUiiJw7VZ8s
VS81R7HALsQdcLe+pgwKRZIpXbi6JS24foudEMlDvV0WJ74qrjxaHP7xKCaTuJ/EKTt5sbvhlk1b
EMVJSqX+mgmUeYO8ZhfVVvYVIvnp+jw47N14U7ek9HLDlyA8IU+fPyt764YozKgh3EpOcXpmr4a0
V4XHNr37r1/kyjfTjYrhN1jp3gN8PEOT7Sxz8ay+5ky+2i+UXGSE7+7TZccJmnzNjwryU2QrPhXT
kLd9Cvm776+hj/nTeJ7r0Q7STxWqgUkegzAi8sNy/asGY3LWXw07dQCIKklw6IExfroNYhczIpQG
IXa2yYzqd3hQ3ypiAVqEfp0ljj9Ob9jxvixlU0OJgJn93aJL6DVydMR1aFCgBmWb7Dpl/VekFgjb
H7AJek5rkfakEPtpIK0jYVAqrdDaCXo7QyXHM3D3styPvf+KP+1aybsqB/9wUZfVJ3xQtAZeyBcI
W764Jk/Ri9ACWcZaLDe552Lq6kZkTOzPwOVsYRPq17/m5JBccvnGt6hWIiVJ0pLK4ru7uhmnQtKO
dBmtZ0y6QFsHD2xGLVcncvznVKXm53wCk0ycnJuszlJO9njSarQjhjqAqz+0JVQSy4GlPkd8gIj5
JJD2kHG9kgEWQwT4En/5/5PsKFrFfwl1Rlg8jLEp05S4w2H6nASFb7jpAmiHnuO2jTTM/p6/+f7Q
VnJs5ZWfk8SPH9v1P94Eyh1VCOYuuvyGthwyMmnvEJE/+//WQ3dVBw6LZzmGvo+4aXjC89a4EsQf
nGwxBz+sKEooSgieh/JysHYlLnxaeHcOn52N0kDYWZeNYXcm1VjdcxgxDHwKqbwAdzmXtSVBdLI4
6QFOKOAv7FP+FgB8ZxGT5YQAjWhie/3PREkM0R7oOC5Rv8WAYNt6KmJVuq0ypITJd8QCEZZxoD7b
0CaCa/vD+Zczf0em66dzJDbx7hyUM74kkZ0sHb6cdq9a2VYm/vON2nf9zbjTB8atkH8SnOu2WaMN
GFY46KHYM9YSGt4VtvhFy1tWLhXJu58IZaXaJRNquFDKkQICA6KYqO5zUS2N1H+6RhLMdb1ohfSP
NnE/erAccQG3/rmieWCsCNx5BPlMOuPapI/62/RKDysHcm+Gc10sUWlkY8okUw3VVdtjIgRH+bIM
7EW0n91Nv1GAuPX7RuPSU103rznye+wB5XqqjtgtskSisl4jf83CrwI8+J8D3T+C1mS8mBseD1vj
Hmv/F7UGH0gT5bHDyHL5lPCYWMufTTTF7atuJJIec1ivpG2D3xOwZZBF0iBHq3TKkobM446yWcrg
l8lDs6ql3ntrE5cLIgSklKNT8v/uuUX6kJqni0Y55IMC0GIfSrgyDz1NP1nHqMV0YGlYkBn/4h3T
N7rNmXwvOvWHCZiIMhB7subLQfZQoc0CS6F7ulz5zEdqM7rKTBqcdKA2F6ckB4PtiRzWJzJV4H+A
712bRBt8DMBmxPNH++U0DBlCgIVj0WDBxTXpPRupkK8C3d7+87OYIAnNxx5MltFc0IgIt2dpnpIj
g1rCOlO6Y17q8aN8ofE7UXTFf3gGaZzSMqq/RJe5LMTWUJBi3DJ/OnuB1Oa4XbPeeU8NDZRBO0Mp
3COQ+JZZu0gKd+pCH7dO/NvWusLiQjxejFHNFRxM5E3mAfrgk6w+HykOHTu/bnr4XpiQfwa/QW9/
nwQKslDCILuy/wWoBDpbphEtu4K8VpMbN+oZlB5Atj+dn7aa5dDgzl13pMw+m5aaYeZb2MTc3GfK
k4HckVoJPsJm9HCDLv2jPHzm6yUE3TjNKuRQGTPxLlBeghgH/kWMQAU8CC8Da4h6v+fINsUdTV5P
1JypPXrh3X0/kKhrPl2hDxhj8hUHkwPiy6lQ9HgCx0tC56WZC90rknJVhMtORfjpdv3RkmANOqvL
I8LM7cwtfkg01ENnyvEhkWGRNvBcIfOrnNYCdedhJVfmzvcg9OHce4VKmoHp6xyjEewfFF/gRQqY
YoMCT53BcAl4hbZ0dR1j7Xb2FmD6I84IZqoO5VAKx2KdyGK/5u9+4Ecxnhoxf1W3HMg9HmjM/mQ+
BuEhBb6p74Tmkmqb8IzIhmqr9TP7Xe+6NrrQpr68WDEZpdIbSyYYjYC7PPnImAVAJWpNfCfuaRcG
y8Wpl3+V7cQnXoUXDQ7a/CHvHXSlTxRBy/mH9OWpzSA1AMDUJo4Uu6c++AXDjJlvj44PswcKoWfv
MzOF35bLeMcshX4hX+6OrNpBS+YGJ1oHOey8M7Wocie+35TsqCrsFg7cVAkMEtwaYrLAbcpM8V6l
cSSH7yCm9i5uEF8LBLeaiq1uDkGvS4ic0DUzgLli4smPtu2gyKHlGYklWbthpPjXdwbllINMK7G4
jewDHuwl4Fa6IasMCb3A3ecI0DE9JXiyWrmx1tr9zHux5xp7zIKZ531YG1q5RveUPLnoI+mrJnvx
29PJk01fSDF7cJd+lpF+zR4j0jL28sNca4TWDj20FtX3oktGSei10dzIa/7m/SVqk75yQHcerxEE
StXfvmAkcOxqrZsUwugBYh1Dmf8ZyoEz3/zDKxTq+FpB1i+jNO5vz0sozY62lcUF5IfQ7YreEtL3
iB6JAHSMGsclp1utoIijzzNAi+5pU2l9GIDEMr5Ti+jCLNDSTkTkPuXDrXj7AfQMvH/+3FBsmJv1
T1eT/gShsvdz2MuxZ+jXWYbB0fVeZ2FEIF50h2ZrCjrDLoYKmI/L7wXNustJCD7gReVb0NPY4ZwJ
GyzntMSJ/NZ3PQSxFXOR38+RNvA/kL5GbWlfAT2oaA3knVmm7d+5FMQekXgVYzOAZmaDq/PWxDEj
p8ZCjksGncQSXnHfxjttXLmXBFecUPFxwHKQ4KA2TvOIsJpvjA3G939Et40sfi4rFCRYSVl7CyNT
FuRJErT1s8Jje21cY8OrqdGGOZiJQMjy2/dsPpTX/ooSpthwdorjk/7qdVL26leAKssYPdccjEzb
HmfOZUghgLTOa23ex1gxjlOZYyuMD3IgXgIxKcYzfqx2ShuAPLXzrLb5hUTvwAy0kfkXuodKNODV
/zMH0JihBSnb3bGniiboOZzSVERoQ4k9jl8OFUxLuoXApA/kRIoWke67p9Byse7WhFrZvpXbPByI
X3aRlJ6iUtWiKqP1FhxVCgSR4fAY0RgzCiNxTic8rqjSDkd4PIab4juaehRi0KhAYTTLoXTi0AZB
xMtRQHXgxXgFUhljgHtGuPq3zH4udSCT4lSCzTnFcj+VkgEP8pHc0a29vBfRzw6K3fmHSoEf8+3X
2NNzPCkFmnIB/GSUsCUnhFxfAGwEl8X+OEqZIIGjBivB66Geyc9n/T9fuEsfkyzCJtmmQDbz6VOY
hOvYdS5PlLWJtGE28p+4zTwezcC0n9xloXldbrzpiw1Sa5MroYz9/cEM7m8r+DrHPSs/IdvLlLsj
//0V9Jh/NpssMc7VR3ijuMAK9SFsu0ImKchi7UPpgYSWJsIkjVqHsO+oXH0H5pRw1a9aypaTBL8B
F108sLDD3IfDZJKcjSsODhv1UibGuJCLV/VUvLUAd4xvchduJoGvHLj6yToT/Tb2zwU+PtqAQBnV
7FlHjIZt4+OYYqxW0yL2T8ntP/vwU+6F7XcskORyIpYDzY1OFsOHzfcezSZ5DP8AdkTfGv/r2ZLe
3wGfj+c7VksSDllnjH432TCrTrNByWT0JB226TTKv861bDfITPMc7ZakSg3LNE+5jKi6wE16EQJy
9RWfqPa1ew/7zgcj9+k2gHMMyRI3eutoIVJI/Rd/tvJ3m1h89/n4+SnA4NxpXmDrdk1I6TQ90wyR
hfupZ8E1aCvR1/rwpSojxy/subbWSbJ0bT5sYLwKh/I6pBIfhqO6uac8FRTgA663Yq+Bu38viGlQ
pzQ49mdM9vE34iM9iNsFkqu8qaj0CyiiV0QCU8XGfJEcpb0CPrw9yYCmAnvDztsXbRh+n2qEwmgh
pHCK/KaGnxHi0VGRQaU6G4Gs8TGVV0kBxTJ7+ufY0FJ0yC0vhEpmKiQIjN2wS2nt6TsZWAEtgWSu
vkDIKJ3VBqrzcpANCXJiitQKc98ElI8SwS7LYxpO/6hWU7oOiH+9C9j5JDOQ1YuUNjXF2PwURCHO
tJW0ix5O8MQOY8n12pBuXMoIaGnAUrCEGHJ6Off1n6HuyYBFLFfjEr5FLVGMXO9vt7epG/KRRW4m
KnZyXVYFp+6QJhoRKbCCFAcZsedOtVH/B+X0HAW5V65V0CVnG7Z/u6n6OS5zajaPVFgiwQV5RzXF
L0JxoEmUP+eCAD3WqVimUkIIJ/Erl34ff6Le8uk3f5i8yiEzj4fTamdp2REzg0N/zDwN/O/QY9cF
GLqP1sTR1ti+GVe22eUsVljoRg5ojLYZ0YhsNGwuTZP8GTBS/cjrnKinwkqOUZKSiZ+PTzWiFm9c
rsBkFI38JNiwU0/y7oF3eCOq2MrlmMhGl2bS8uyFBtNHgx0LsnGcytdrxR+cGniwh799tBwDg54I
8SGvPy13MPM04RPtmITTIHQKysKvzTB5mBfSvx5iwHAA/1fWU9l+1utYPCbzp4qJCq9bAis7uF1R
CnvVldYqqje78rTT4juvlZitQe9qM3k1fNMfMd3sCAvqPNUXGT7S2WO1tsP9qXr+75hELViMxFxT
Hzsh4OFnK/CM67bk/DxWZwisDpknbR+snpO9hbIIvV4hsuoidSA3kOzCJNOefZgoJTaSI3rIst8A
R9o6rOlbQBHp/RnYlRKv5qpmIlXkmmWs49hVdHH3T5HR0jmuue3vU6nlvOD5ktNJeceNShJS6oIv
kBKd6vBODZXmso+3fmCHtHB7fH5aIDUrYhtYGdok8Xuw1qq6DhQMrsLc/9RI02m3tYeait8vcTCA
IeWS0GNo70hTrzvS1kQb8TxuelmD131cBNk8F5NfKGu3uuPN21IBDt021pL93T+zwJjVJuCiGS+I
94TlRTI7zkRf6gKz75juWeA8O2XrFBlNcqznoJq4ha2w09rFWfaDyUznEr7zqV0n6UInaMMAM8vh
JYg96+stsoh+mbtprtp3BByDW4gOJHa8rO8k8Bc6yvQegSM1GCZNGXuhsew9MHiWfEA9VkG3FpSd
UB9EVW2Q8n10wnJ14TsnRpZ0J4Svs5hUyacn4CflOB4sGMDfd9ZJzJd4f1J8GgkJ45QmTDBQjlGO
tO7cy2laTMoyLCpLGgVOcWkgMQWZo//upjFrrcoE+yerW6x/Bim3fEzKOXum8/L9jMGrAQjwOu/L
nlAXIWv4vNBLNtqEJV9+xfp94u/NFhYakrcpUBRy4RTA3VneAlb9RtdYcD3X1hgjnY2VWzqzzzlK
v/tXu9XK3Fexnbbpi8H2WklPpBL6xrXmblyouogH8vim8voT4e5z++QQ82yiY7bmCwFWE0yWpIUD
MJNQwcx2r7+VQK/X1ceKXMlXicNUMuI3jQ3SsfSLLdVFHWB/qm5GQhyYP7kfZJgWy7pv/GEZ4MD2
BrVKyX8AHH0pM+DDbDHzC5dyr9Wid3tw+iJbp9gwzqLEdlhfgxM5CLJHd2E8tTiDhtuEZaYRhTtj
5LKoB7Di42NudCJZXtDgcF7+ETFzH0F8MYnM2h/otqEurqJEOZ1s+ryBwZhWJf3avT1vIGXZ/093
xcFt5Qrg6heJFP6t5Anfww0GhrFa/LG99vWXLBfaspLHeEhVxQhVzrnZti9a03jAxtLXcTM9Cecn
BlJBd1z5scqT6Cd0OBC5cXMAYFU3bp25Pr2MGnvDyvBPVWzOlBIm2HexKVluIZag+92A8kjFFyM3
4YuU/3fQuU0wDsZJ4fMGpKzY9WhK/+Y1RYyj2MDQqq3eqYK8DiKRptBmS64s+OWAD1pbmQLhxZB8
Du/ZegKMSLHTBB2RQykhnDSEibytFl1Iq9LFQvPc65o3HS4pexkUnHm4ytFxP5qevZpQRG5DvHr/
rwvSdGEg5yL0A6wv4orEujsO9JXR6X/WIqN9Ibx9xaAVmSxwvowuPPUVfwE66B1pQNvn2qmwxBED
+3DY4VXNYEJ2dtLNUsQS0PLfDCeEevgGr7EOTd0OFux5I3Icjp8XX/oBzcDuDz3CChmHn+4YfoW1
1cDtCyz29KpZtNUsCxm9WN+/C+/GYCeGno3H/bvTLGckgEJ+9Yvn9/kcYb5B+i2ThLDZ323OuZb+
swSpA/E2zgRM3ke3MOPNjYfOIiOqYtIS0tMHlqhjR/8PM8p5aojA+b6DnHBNRMxDishqvcK23TCA
Si5g2/WiVmxIg1LBfJj2CXO3kX4DF0kMdSuChNwle9iPypv4v//l9W3IlxeTW0owdVQw7C91VA39
a6IlXTupkq1yinCjwrZFg7/IQsbdw8+CNdDPMZT+r4t4vQi2m5zfU0tElRz/Ft4PAjGPusw2/StT
DFTGLmpTsuOL/lP4finX4EncIys12BVM9THjmGz17nAWpK44GIuWLI/ljmEhNc6edsGSHbXM4kYJ
Ibxp2hX4s1Yw0Nryz66P0+yUEBipvUdUj2li2XccXQNLF+XH0U5abdvu6ybh6KOcTqaoCgslCtu2
4rU+uCgVP5GhtuJ/GAS57LuEYtt/4Zgnhy2hj2mXONhFhwJ8QTSIL9w4Z6RdQyHGIXNXeGajpNd7
XzbBhadFoSCAwcDm0sBaH+pK8r0Kj5YJZ4Yj58rplh7EumnFVEs4yM21lsOoeWnR/TkbHD+DPcva
kxCrdJF6tbtG3Ta87xnWPzYezHxH3AlC0D8K6NTTmZq1KC4LagWegvo3i4irZrNsDyfz8qfqnEMF
mAF7g/tdgVZokCU/JMoLikG/Y9Js37gNrLamRbk6uqcGWfrmezbMdj41jT6wmymS8GDM9FlmxJbH
U5HRZpLEp4XOrcqUv1QPWenG7AqDuw4iKIaPMRyVkNrY3ECGlGlHnEGmmZruHzfSOtySFZRfMuo+
kHonCcmhTr3Jt2HOonX2n2jxFdPnRkUBoB3s5YiyTJSTq6BNskusCDM3xoInITMq2qxcrDHEto3Z
jiKG1gz+P9Gw+X1DPMVkp7XnsptOq4VQMaEj7RoG1xluR7ifgsC0Uj18Rj49Zr47qLqpTHEbrN81
S5036pg1tWmYQENWmzHhVpnHbkqrXbYqn/bYQbSKpt6In3YJCs/UJTdJ9PR0WtLoX43qShatj35m
4atlrpdlirchY5ojPHKmR+81e3C58icxK0B+LVjZTaimFhAbmJMWnj5BOIxqRyOPQqK2YoWi7fF7
Zk4D/NgjyVo8kC7ljmLDvflW2L4gRVDddJiWltuQEBYV+bK99G77mmN8Olhxxy+0rldCULkj3q5/
mjczOLF3D897HTrlpNPXBoevqXzkbfzTzO9v8oIvFIRoJaygbJtHB0HELFnuVQkgImAWnJEliHjD
WmB8NWDMIaJ65rBJ8w+q5OPiCNW+NS+bX6wKyyt5oIsgS2MQlwWmZR/QAVN1a9mewWN0pwCnhO84
94KLBBPTJBn3ZU66TgUn0ghXsRXyZg84Fv0xrC7Bd0RZRc+4f34IWfk+ZumuKElWdddPLKAv07GL
gpH0zBMVn6CpuyVPoUqzEAjWn7gqe//mfnNBrJQKoGBZ7yrCv3XWHnlwRiHCA2jFP7w45WMiEZlj
jrPM6sQMAdqH/luOJX6bxiwOnzYhQdY24BxFs76llVMMCTCz7Zk5FUk8h0zrj4dXNM4pkKqNzc8H
RaTC9VX1lBw/1Q7jc3XTdTS2e7UFI66MJpx2bHJFA1U1d+KVxbRT978+raaa9ZgosCElUb+JatR8
ej3tuwKxvco61dUvqNsX17V4dp4zvrT/OB6zutZNDd83RS4gj9mS1PJNM22rnONPV2/ePcDf92VA
YiweGo+uheMgkmmr2ZQhK4wRMvOpYxE1DMt2WitOrImgIxBUKIkF3Jl7uEEsbw8sd2mUNZGppa5Z
j9MVuNRsiRI707BOk9VXNW9wfF43uP//k0Lgryp9I1qJySic7P0EEe9pu+pU1SpP8weJpscXAof+
PCaKl3OisgMBhS0AvpehQWwsjpLrZwJIl0bsy5Y7nF/exIWsn7KgqlJlUgo0cCFXUjux4nqK04t1
waKL6LD4zGKVy5YTmQf/bNunWQMyLozEWWcrEjkgxGAGg92EbI1Y2VjkXPk/LDoMa95k6+Xn8xh7
VItPyMfgpRQVN8MwxJfrdfoOZi2N9xzhcRfKsFlBNHarso/8x20ym+dMt8vhBhQ0ZYr9SYtI+Yyq
2CH/YBjGIdBPPXvl1XIx1953FfnwtN5SLU7h2VOilp90RsZBHA1Wrnk8CHEF8mmPFLfQisrKeaFt
eaxR5JBCR8FmCH4h4H/hPpVq5qZvpv+vj6Bisq05NC+o1DVYyZWeKa0S7V6qKf+i+q5pLX+A0y/T
25nMWKP2zFKuSa0jXlmcMilIKRZX6Sm63QhxM30v+fALsbYndY1OfYJqiAALuuFpvtsbGaxzRB4s
NB9WO7XfRPyvTMoJh6EROGdtHvLcLUnZS3on2fF7vxyXGDjK4Zp/u2dKeeSOTPKorCqvTF+4EmwN
Y/BZtv/0JeQa7UObupADZKSjefrXcGzIJrtPjbvpUtnjiFPrnT+ewsyphA/2FAklQPX8OAjNoe5e
dyK7BOh3hcWz7TIExenatEJP08SYFhouQMRU0m05a11kAqooDtgjvHEQ+rnJpkcHoUAHkkrP5igl
iTwxd++jKQM6pw7ee6d00W/JzqxLPz/YKJbdo+n5JL6tlAZqxxFMUya/he2w/SHRQzVdyGLpu/G9
eqJkrZeOJ85m1M4f+LHF57mftktbDbE/NkaaA0hHM/TwhJlh0E16Sgnk9ucPHXSnPC6gFrW0hLH7
4+dj3NYlnjsGij+amiGgbyvOb+4NfsvfzY0TfHZuV9BWq1TQEmxo0UhvWE0TKt3Na+UQTz8exDDB
qqvzAPlKFgSSLs+l+ShkWaoBSzKNuNQwfJSfaENqZ1pR1j/rW3yByM9TLGOWJ2tmz+kCDp+7ukuE
h3mSRxLLLF31APYU0iW2Hrx/OHIqIuVTVYSl6e0SrXXSglzrYC8Blq/Lxsh+oMnG8EnRRLmr7YJD
MP49mk7Ar4A4J6q9t3zXh1UnjZwPfzlDNSUskJEn5UyT8TqllIW0t1t6WVUV93ChgiJgadndYefX
yStKqrgp47YdOttrYgmWMozPKqCD1Bq+jiT38HIXixkUYVSksAsVurm/x9o6VI5qHfdZfxY9kYna
u73csXLC3AEpWBUdhoUi2wzSuQe2OQ8wXM7eaMDK3uzBknZX5cR/b2XHb6Sato0OEpC1+POzoxBR
ZBFuY8ZiO03A1Hw8OYwZsNHBOFS6lCcgYJGb7HxJpT2nhmI0uhhsfVzkJd4bo2B5TYzPgOtIQAxI
/8Gwer/KFgX3sF2HFTLgwUgqgrv0B5neenRs+M13uaPIcyeDdex3px9FcGPgFd9iGfbDZtSD6KQn
iD/ZNPaRNGysS7g8iyaDRQui/lhtueOgNIUmlh2v6Ks057+ZYfwyK9mgLIbj5JM35/BLAIFvsZFJ
wzYbE2OIedis7mThmcl/WKjPLizDDrPvzMxeD7aWXXz4Pa0n/Q3KBtvZyGMZzt2EW8+ozug27iko
II+hYuK45La+sGg2ycsC1xnAsY+52vphk+5L5lhSowySomiHzA0NaIf9uXQuKWGo5qpO6hgRqwDM
Uf6aWZids0Qv+wsoKlW5ntIjgZoNyypmJDd0Ckck+h0Qu3mzvNz1kHiM/22UYSimVy0domu6vavS
K5S7k4SxOu1scw++PkSqBzCsPqJRxx4dqlDU8FZz6keDP4TNztPeQ2zgL1j1bgHD5BOp1iSfs/uQ
3clwxJYUqr8vC2mkGBghueVERqS40u6zIMNxm24vAUqXQv9zUIH30dVz+QF0MJwMaWSb/06jeIzG
JVLkWUTMKYNRd1M+aY7V2LLVbzv9KmXsV91lRuctWgaGPKI+l+outmyMCRKaiPfFm7DQcK+LwXLh
d/jR1F6YRc00kLqW+uXfs/VxHYt/NcfnecHFPoM+Hlo3S1mYNscjeEALsGfg65talaY/J7XwP+iF
OsMQx35Xus8gEVlmC6cXbezHH1NKFG3QmnKpDkVqyAC6D6CN7CeMdHafXhCb/x7VMC95jJk5IwmF
bgXjiynLo/L8MGinLuGztPdk4gJgmYLau1FXntX0FwIRffYstwDV4KLNmvXdTgquBUXYQOz2lrsp
JoJ1vsz1unQqhzr12K6e8hXo/cMxWF539SV7prrpLHwvvjWTWyI3WDtMNKxi8DGg7iigrA7pRSjA
CauLDzJdPghRWvCGKJBE5SU4U+FCV5cZnRPRfuc0nTqKYXuMzVkhR7qUpZQXY/0nPstEdQHNnUIj
a0OmG7A184ctQrEZYj3jBAknQI/HwQPtjqjV62Thh2J/uLbLhxwcv1teTP/GjIajtRIaDcqzX7eC
D5L4U/HTASTGxHNSLPRFJW/9mUkucJ4iTnZ8NLH7hPZ9pM9IiOKYhNPZATuWXFTzkc8aKlgooxDk
H3CG30ADp6kWlRHfJpwPafAvyYIMwnEYSn6IDOCy+zPXgWLERqhTb6ZXohYvQKF4nxC2lRlRZ7PM
UfHLxx6Y/h993g7wczsZKubxEITQWakdof2IeD9mOfpC4P5Xx2+ZweBqhlYS1yGqLKQ96KOEPzqg
SuMFeInVaDT7snbgzS5ADA6Ip8hKI7KuTfEyod9zWxHjYItZKr0njUIj24or0LrICQltHI2JKgB7
jiLf2nS6DLdAq4QvNO4wuFEt1Y+SGp4gW2O42RGlxfJjWkudnHm03AoQn28Bw2HE0lJea76bwXDa
BEpEvxdARagkIgucbrHZa23jEOy3dnuOYuu7DVS+c30feGgioGU/AwIgkgYQqSn8vdzet61uvCdN
cz+vQ4vW9z9MYrIivzx9lmpmDPZR8MWDdq0yCSRg6817HfLD7gTjejLDBxKpdyKDGMS9ybjn/Um7
Cq5rv+DtefiuDOgtNlvPMJrFgKSw0+bLL6pqGn7bgRW9yzxxwxL6xLBVDXV3K3C83kh9PXidD01c
0uCckS+D4cu8Hi6E6RvF1nUrIUbNoDVUYf9O7iJaTgqSufcsIsjHZpPYxJMLKCy1IhSK4NPoQfX7
WtO6eMeAL0xHV94giGM3jQKohD6oyVnUxazujMJ1W2DO27YeeUc+g6XFwDBoxk9awfC6v6Sy47N0
mAiOVqN06ndfZRRKMMTKZPWm0LtKff6XYe+a66ZqctW247utZOmJKKAUz6AL23Zt/5qWjeXrGPmQ
pdQprE6Xxc2G1Q/jWVAfofwRsjIa/mydG+orh+7CpgaWQ7bjD4GVzwGLzy43EQfRrso24Y7RKedY
rtF5R+2lmz1zKVJU7GUSlP1n+P8TYlOD+sIVzFa6mK/t/zj4YRw3zLWHZPv5otI2P4tgFQ27R3jc
XZRxNtJAK7HcHXF3+LJDOEeSF997XoHONGyuwlB9gh5q6tL8O4ZtynoowuSkTx/iEhzReNpbnqaI
II/ciuANk6W4mucAyqFmQcUL3k2YW69Tre1Ij/lo57IW5RoARBjJxMj9f1zj61/yJfRVSQFeugFU
fRWkF7JfLtp7V/zWQHPml2mna3BSCU/YZztyqdnbp4Aey9GZJI+wOuYX4LsfXrx6pQHPJPFPDYKN
uohqyUbeMMU68hEnAUKgZ7USlEuNiZ410KDh7+q78Y0D5onzNbUN1cfVm33i8SOJB09hPS0KQncE
HxAoZFSRlby36U4tF/CJ9LaI7TTb8eYAqA7MzivdqX2P2uoTyvuNe/KJQtQIoKM2Fzm/Ye1oaYkD
8VoS7espiOB4E3fEA/R68hL7DElCsmTcYXrsoT6aNST83r0bMs1EghGngP7dG2tZrGcTYaJKtA0T
phDRxh1DGBJusfSHdmv8FEqr0bRDEiz+/ufUF0as6yzXOo8QZf7WQfe65UmZ9d/sevfzMbfucyNR
Zjt1YxIlrks7MQ11CAI1mG6gmX7qqlk2T78V6fKkGWxnr76MND/lGQ/cXzy5PrJ0Iet8lHyoXpA2
IEV5tn9eOu6H6kduksFs+g/9STPKmkSIxxmGFel9JJTK7Oi/maZMNXvfCrEFD6+lYgbu6P9hC/Ci
oNU3RRdd7BXpaYTihkBq4PJ9LmMfpgAeBDMd/3Dzov4FiSuXecG+SX/SRrev6JKjjTDjq+By4wOA
AWETMCRcufIm0Vv0MkyOr5Zb1JQ3ih7Ujl5rCMVXLB6MLIteM/pHE2PZh5wLyg6GdKDyOUhlMf5Y
yaop/uHstJiwF2Fdp/M8454WMZAgPkafE29gUwPmSfF/RFOkGMgT/117dU6+dTrrKjcSFnhtiScw
cd8Ud+viH+Wtzu165g63wiR6I+XzvpBEV5jcIZ+MbescWeDkOIHlC5qir7zbGCpt6eLjf8W4VwsJ
eKjJj1aZtIoWz0lssXGbGBfj/X8IbEC25mTIN9xFp+RTTURvSX6R537+J7x7tCegxnIBlU5gQudm
DfNDzEwYFE8/L8mMFhbQK3OUZmvxii+tEVYBOednDoE9QpN47v7fq6o0N9k5TWsHXRKDSbIYD1DL
TIeacV5qIg0DD8AF83gbbfaB6jDXSJEx5Vu9vKOLJbXlx6AFF2+MRDo1+VYG8wbrWfrbdG2WzEXc
X27WNj9Cbp1fl2n6G/SxEZACdZzgjQZHTLB/eE8RO/FBqqANH71MdWgZ0k7hvRo09QVt4HLSDk1u
qwD69Tnwa2FD+9RVzJT3KbcY4z4ra0E/IYVJg9kAhSeJI3XUaurX9KIwKeVAVNZhSKsdZpvP+K9C
dB7eGO+dPbKH66+DPdsrRodm/Mc/zuti+uoNRDomcp48uoubzsfT4zqz7h2GbM3lJgY0x4SMzW7S
FJivtljQ65bPxg7KzdnbMZ2bQFfelZpmbO1I1O3gpQsU/oTkuMf9vSihK3fHQaNcjOlCfagBWCaU
hsBkhqM8mbXb/zRTd2BUbv33EtJcvEIoutKKteuq92H8nYhhSjqpVaG6fRTCrdQWOWDheVcPYRA0
WRxEw12lbbZb0VPuBUHTX6rPaTtdzRYDiPdu+N1YKusmyy83s31AZjjJ6D2I2McgYCttJqRqhwth
EdtkNLjEOdHvsifeJ027EHCmYL4bih53ra51tpox9gkO4bgRUtVCq7FPBrJwGlR+u6upWbYQ45HQ
fxdfM0wHdRUtra+H0/Wz4epWAN6fcyno+vDMsC97W7CXPzt2teSj/UrpMV02zgaqrwyf+UMuvDYc
BL2HM0y+Y/d8RZphtf7Wm+cXSXGBRVTo4AMOOu5qDNps3NHwGDOuyfENrC8jNL2xPeKJvyBRrkMQ
RSj8BKIs6TjUMy94Q3S7WDO1vXNID3ffKnFzlE3OmDF43ITAY5jRDnole7L+PD10TUoWTWft2dKd
jxSWymu5iqz7lxsinXrhLxA1gPEAw+kVb77QD0yOikHOUF95xNqp3MAYlkxG7p2V6LOdR3RqP810
ir7WCOC962dsfSMkpWS6iDSmJzMm1AlXKqegaolCeUk+Ztacc2jv+QDEseK8F54ubtMGeLLjgiZQ
xUptJo84SVsN9Kl2u0BXgE8kxZHn0MkgUbFFFGzYp70KUqOlHlYeFLJ0Z6yw0ikoOyLZYP3h1KzE
V+aqDQxyT0wZg7aW+jmXkrRyQoie30Qg6rk8Tn+xU9YcZUL4RxBCsWnDixP2deAqIjuFq/l9s/mg
4qlCzjqIVrryWL23gqQ2si1cTHUVCLOTKyyfSsJKMDWzfX78oEbCFC8EzZMB184tyVJoV2NHO8k1
We84We2eR9vZzqlNqmANmE9K5hvY9W/KEEKyoqjM8DZ4wQlGt58n82j3t2jpKg0WL2fD/YFmHkAD
tH3xw1jtjUybiF4CQMe/SL3GSwwfVcOA46GxX405nOEjGPtHTlO/MZb+GWDYIT+SuD6iuL2j2JmM
T5E4Qtn+HSXcI3TboG8F+nIBgbU6YVOKfFFG3pfvAmxiWSLr9AW+heC+E7Aiivt0yla6b8FEQuWB
SUY6HLZzQk+ahHADwGxhKjZ+EvLmbxOQpsvy33B3BGtlBXVUHssA/JZsc1mtndFxb92TUH3JYnUM
0DEs6HZXqng0hIDYJuwvkd4vyvT0ZpVhCW4/6Svy2LEh8VP/05/BYEtiX17IKF1dwhQSWWWxEDvs
k3t6J/x1g5rpTCN6gvuyvH4tYNJF7rn0SFf0RJNjRyz5SfN+xbVbhdYvsZySaefGiJfxd2ssVKZk
g3v9JhVRx/uELLs5Ask0dnA9i8+y/w4EmYhO0nnC8IukooOILNysGcZcHpsT7Yoqb1KiP22XLQtX
4ZABtAgqbpeEKRIAI0OnZkdw4x2v5onjuSY6ixZK9Q+U/hpH2KbJYj8CMc0tlFvpWjABrvOn5+7O
IpxfYKSVNlB2Le1goobwXLm4RhsaecuJAbeLtFfZSPNAMCKpTS5fPdH97h45PeR9lIK/s7/6O2bA
p/ImfgsAXnQp+zk1IYCbGxPk8XuicHbDn/2+69yNOaeu5CkQFUeq2r3SZglu/AHYyWjylYt9hrn5
NUYvJqWtzh/uQxA0drmRmBIO57PBdOTNyg+TLKsFHaAh6iZK3xuPWUihUpaM23LqUmSYuIPuIZ3C
1NPHgGhYUAP2wDDJvNWiqB0XZT3cCJPS5ZjD3EqBlFYGFPPI1CaxiP3xdT1KsYBgAPW+w07D/rse
XFHoTy1tvJ5ij0vpqFMJQbFVxeAo9m1N1oRF0CupIOrvylmtlbA6aL6j9ziU3aHD4VzD8zkoJbJC
P/3PWVj4umDgarSu4Yt0Tda37a4PTaIOHVFCY1qGJGNSed/TjyuGI7r9JG0sgwGddoxIgFZYfBrf
aAsIeiSoZYGDa1CzAmWJrzdmBjbLDS7ZN7HQE3/ThARoFYDxeCkWn1REABbIO010asIIb+Z0FwA3
RmU6MCfs3aLsEfDAfoSXoRhkKdW37FnUzzJiTmnbP4pwXKj/OwsholICTN8ZLLOUITW91eziFLEz
oZiwKwd17x+k1ejOonf2CsHJ2BCyyhJHZtlF/Zj+nyKC/7ZJED4JmfP/4CDSgdZ+9kTG0gmpWvGZ
nLv+L4y2Mlf+VqFz3IHQdaIHCPC9RtvnEo/0hObopQso12Vjx2B5osKMlIiagK0D0fIWds7XdM0u
X7//VplknaxVsWxTA0UoClxMyXym46MrNyrFDgFHCMffdEhPurTvp/UaxvgVD/SPg1N4PnF4pv48
NtXnyTptP/8oKQ4HF+6m1iL20Fu/e+eZBzqSLTWvUjypkgKs19Yw9UhrivryIfDZsRPwe7x0pRom
Ui0YwAXKY00Th85UHA6hwq2Y/Y1aMm6+N00CYk1+dJc7KdEty5Gk+wHAyYaM4I8lXtV27Nzg/p9q
nuagmV2rabgpVF8sVapCA1paaH0ianWvhpczd2ppKMZISKzvnLu5Q1GR+/73GTwBno/HF6F0PLDu
5dBOM6uzyC4/Z3MEoRX0+LNSUcHGW6FGRhbJcSZ+I2NAMDnAZ1pIDyzSdns9VS3ZTFxPLftfCJMc
0jd5mRBUoP2Oqe/lAr5SU44TCwrId8gifiCB+50MSZkPl29rhZOciLw6MjpyH6SIeuPBoRNZeAJr
f/cKhdo57w1iV7KeZFeKQT1DYetfvLDXS/glfuO/jdkyE390HaixFn1KZ2v/UGV7YJEusdJ3pV/L
B9tqK1/mkNaRQxDInSO+DN6yXoWdVKL3cXptFIUj/swWgvvJ+gqhNTkB07swtIxqngHGRkUS7OU2
/k7ZYF5Lss4kpSF7XtKTTK4SPWWo7FnhkSAXuWpof0hMErR3QnyLC57mEnThtjLzCCpGi01inHGs
pO3t5hyxKA4huYdINH/HqfdUIYcZd6h8lvCvzQ45kpzgZD5lr9pOmYV3PG92UNsuGAojRLvF8/bW
U21xBrOKTIFYf4O3gdR9NIgDRIcMNpSAW0Qawo0lA+kBCH+lnSuk32rissa2QDob3AtSCvYv8aB+
HVqLGV8r7EsIEOW27gc1pfGJk88czzhL6ntBuAZnXViv9xA5/Ky5fS6bjkDoB7Fk7jOb9UTqu6C1
Ns4/G9Jp6f5mLIIHXo8hwOKBzqN6nQM2XM9vfJNJRyNGT0YVx0ZbNXE7iGgBBekJm14Y2mveutxB
o7xfkiVXYlJx/SrUx6f0qJcai5YwVCPPS9Jtc4jkN3WICkaRvD3YVan7A3/0RIVucSy5TVsvw3Bg
e21RdpDXSJcPrulBYYVMQuFcMul9fdA/r+gxmcQO+vnWseW+k5VrJN56bcVg5Unhl9VzRczziLYc
Om6y1UFRU9xxiWXGD6zGadLUxqYJALntgqzH4QbcbrLdlNqyv3V6swbqJQRL3Rq15T0LGtY9W69a
LdcOWX4OhcP4gudFGkszgC+PSdYuuR8innJsuxWIrA4HIwZE2bqp3R/kePscU5mnCYi7vLp3QiR3
ofSRajD1iWN7JcOfznakjVPPb1vtiqvjXqF0KQwwBEwqnXWJzIJPvqXGVh4rcKezCXn8fFBYlA6q
FT2txEApluy08XFzO95LCamYKkbjTOIVJ8zEN893aLOGfhCMGG718TMnd4seKn2uAC5FA1r8JvtJ
1xuEKQbA49O7kWojDwpY97qnz9nLGekA48BokHYC7ZmiILeC9jnKGjkgr1I0ByphNdTUmI/2MaFf
QXgEhUI9kkUDMMIKVzAvtWBQ2vKN4C0RYKmJUXhmRq6XzeN21Nz4JOlbhwXsvwsTiHnRDnGVPGcT
WtUSjcP0zWV0HvZKF8diWdIEFwfH85BUhEiANYUNBH7rvlUk1GAl6HAgtJv+kn/riufPXO5vEIdX
ekwjFq/fAdGeUy5MbtlLmYtzIsqkE9x/9jRrb7nOrSOsFCGQ+XnpRs9JEyNbe/RhGuSs/T1yFq9M
QYtZIURtuua5fQmE9qwqB3tjzyoKAQoYRaxLdapkdDGU55+qC8jxIlgYfMBoXH/tnbvj92S9NMjf
XzE4cCBskorhsnx49BYKNNFLvBeEXjVoDygT2Yt2GKZPSna1aj9OycdbJ0m5DG72gBDTVtx/uxHq
c30ivmCLhZ2I2u1u8eSvrWtcUtbXezW4O1HqXDZUAPJJoTIjNQBq+CA7SFA0jpLeA5qi0hPmTqhW
yoXHZ2cYxGf3tQLUSIHR15PJ7kVWKkMhbE+99d89V6GpuNMgG76GSNhKlEHjycVXChHOvhfVv4mD
hHUtdTRO9nX1EIpboruue91onXPKBsIaoVWEALOrqM0CUpMvxAuyK6KMed5+7AsulXSnUoq9voA4
TA+4gQCHg0jrCNVllXbJFLv/OiTif6r35o3LQ8ocidL4T2e01HZjErYQwBHT/DyeMgEdfCHAfIrU
hXz25vs+qqx65hNXWSEnwPKTAivqPaC4keSArJWbHPoArupOShR3BXZgnQOtDvuVoeR2BpjcSumc
N2vMrcmE6eOgizVtDb4jqRtMDP5ww+9yAdghz04A1FfFwN3J/bqRfeQKNkQOOLW/YWJkrN/mbVg1
0Otvp3FWqrFMj8eHoRDkgcp/UT9K7lbxOXtZpzXbpqSXr6obIO8k064hz4RLX7eDlB7m8OWe0C6o
YPz8KgFviyw+e8jRmYTIXkwGRvyreMadRJI1PRMDBaKXo7e/YAfX5sw2eEZ66ygStCtYqjE/QvcU
ws8/AkxjIHrXG7O1ftWClGntoSUhxXB429ahRz88lKARzH6oi0kriEBtneCiSUxqIgGVbjhxAovj
vVbHzfF31757L8iCu0LZfnD6c6Fdx+P73y9EpTcEChVdqk8Bj99BWLyOiVg+usaLRufz7Bzh5m6j
VsWVcrxmGDfPgDm8yIi2YygOfIczEQf23CQQz5vNjEe5P2AmEmGjLnjuyA2a2bWy0YYU2BU61Es8
yFSmNlLt7QMeRXBHgD8UIt5sj0ZwSreZnyyTq1cxgN4SejUpAQLegv+y8SgVIo/Ew/KcNGhE+PAa
6ZK4wjkbbUwy3+5zViolE89BNmMSzGHSyNoGxPztWyCg0l3ygqe0JajhiZZajdxgAaxAPasoEylw
YlvYAHTkuaNeLOSRJ//oEXEnVEm2huK4W/OSOqzMUt4dvVUTU3dlNErphOKCjBu/ppr9BV/OQ6s8
OwaDPfkFeE2mNwkoiQ3vUH+VlO6LoSaCmUNX36A+Sj5kHgioQFv0i0fi0BR7NK/gw7Sc5MWC+e4h
rAgc8WjriS2Eq0Hp63hIWQZCdv1nU/WJt/Je2QfVSGiZZ7pC+HizmHjW514OH7TphJgubtkY+Njc
2vyNLYr3loDtjjjVWHP3lS/+dxf9gvddzK/v9pvYOD8fY8y62DpYZYFARxWPOBR6GcFIJCx6X8T5
XTvqHINoEdxHkP45szOjNNLtF5LjoRVwFnAAevEUhLQ9y3rn86XIG6Osf6o9JzQ1vzxCNi6F2Bkx
JrosVyCORRWsRqk2tl45ot96yCjCjiBNDN4hnpXahKQGqiadcIg+k+9SZaCDsrUmapI79ZCRHl5l
me+EpAM3tgSOEtnJKmJtf2bXHKZHjksAwMJVsQ2rXP4pcv3Z5EWFo7gV7xwP9gdk6ffCPs+SUoHm
8rV/MuJh22XRBbrIsIIPUV0g8Pq5AcU6AOvJmFU7K++6Pr7JhhLY7UjxUgSXeQskHAE9bFkkUz9b
Quzcu1H24g3qXIJ11Pd7IwmU4ZL58ohMqQ47WOXuMvEmJEaTNZThn6+i9PH/Z6k8ZSNLSAvaeyuG
xrEqWyLFk/kcgtYjrSsWzCxBDHhPn8Ana2oBBd+oB3lsqjTwUM7lqjY/l7A0MwcLXh99vsigpsgB
wHWzWrZiMyMzvI3ceNTJNPH0QAeEU9Psi3UnPuGnp4/DaUW0czjune8XIgolvof6CauHjWQrzZGT
IorUir1361rqyuCYGbdB86Jk60OtX9oA9W7YVqAbGfLgc2T/C6EXHYePNoMe24GqzMqvAnlLZLgK
5uyxHScON4T+xi//nQ6rXhSBEQpkUgXXe49zGm4R1YIYzScO0lxTkwal6kXmucojWiV5T3DuFP8J
+6KlXpPV0IPXrWst/1AQ0ReE47Io0vsnw9uwQGGgpxAAeBMqLp0D0xXSa/AhzMwu0Yclyq9sdH1K
o3KYkf+2VVRo2uqVSFLbEDKnmFpp6ocjPYh1VHdztyADb7DgHMCrekIQHWU5zSvMPxoEgyL6AwPe
jiMFJ6ZsWlbRM9vxQSjKMNzP9pnz72Xd57ky00eHQCdIMkDg6rGv0V1138NZiy8zeegq0MnUYM+F
yecoRHPkxhUHL/q/0gXVtidSLt0TkmAZ43XBT8yEtyhI8PLzSPNK2NG0eJqDz86rOVw3kBrdCIgL
PYaW77EqpSIkwOo8Ydrl1iL6jrcsNP8KdX/rnwnn6y6330Ip/WyDxgesSmtKq68bwCNT+5DfVoss
YYANNe3UVqdMdMLXb7cF5u8axYANk6eddpZ2Cxb393Pq22DnC2rDShvvvJ2VsXiiJJyRm33D1bpF
IGeBvGNWDL8EC9lyfhpEXW6EApMIqR7mMwV34v4zZjAURq8jDsZyXKxzQY8+GYvt8HkUR/Psvlct
xde23diVpheI6sWNrJw6Ns44c22/kCkoe9up4rr+BTAu5UbiGNszfR1qpY3zAa4BnFkOqS85GKG9
TqqdUwYxF/iALYAXjBMLRQZpyfRq3e3zgTFzAE4qt03oKFSaW5xK354zfDCmbQU54YIKrxjbXd6q
kb2hOEU+N9SiWKjFx/DZkp/6a0SRpUasxqeE2eSlpNm45z40hDUD/0MwWbEVxf1hVdMNoxXumgYF
bbIl/0u4fFjTKyKdE4ONqQ5AeIFxEhhuGqn5GTrpMx4+iD9tjrt5PIJPq6CVURkqryZz9lSFXnig
py3LnPbG2CtT/YKNK+/kbnwbDhgHBPK+j2O7dJmQqTJ2senufe0fgC3FZoBtCf6ibH/4jN9HXmrz
ReAtJVw7m1c2V6hbfQvKzJQWdn9ohi0tWp0LY1q4fgUqtNXGP3EUqYL/uM/fYFoLCJpVP9dOE8XM
a25ieYDPaOs00uMGvu4Z28IaaVl3ex0+gk2cOZHSEZbsQE5Rm0oUuB/rmWOAW4ag7jS3y/nG4ldn
fxWHFoaEhQPPkp9DRmcbLNskqWAf4b+HaGTn8tRgMxhB4fKLYoTu0BzKY2gaA4gHAQuBkRYbix40
XeRC5hvHURgudS8QYkMdS5NbWwIFtdVGf/pL3KStzlSpF96+qJxzM+6aT+kn9Qkh3trdzi4zan81
xkgRXy8qGfTBkr0+1xwmju/k4/2d5kHsgXMg7PAMdCKpzxXWAG1zWu9XEQRvrvVAJPJj8SjpmhF2
JptVwtm++QaaW7kqBRBPcw7bTLkbqRnMODu6a1/+u0JlUNjXGutlrwZ0GziJnmQhCDby3rOoPgOd
GFpdTm3PMx9u3Cv3LYEfIYjAYV6QMWkEG7vBeMPI482kC9qS0tSg3JNLe70vYhGE0nr5PSJCkwS1
X9uIrBo1CY8xqGYjpNM/ezmD8ED5pR4XpZq0e0EtrNpF4mMk9FwGsOrKjW3dZXNB5Y0kRXWgjEw1
EGJBtx/C/4zst5lve7Yq14IAYk4AGEObkQqv6AqZzXGjLXOgkuyYoICnRs3zazQwGp3LmWGa9nxk
LWAYAWA/VRyWjzujYqDCYGK6fGmeM2Zd8fI5mBGVJk1poztxM0x7t7X7/xjmPvLO17DLDZeG+1kL
f40aU2g0l3ZucYaU05wpQqWtQ5u2He3CNaziviaC3H/XEJEk1JB/s15ZVW4fJsGJv9Rj1JinhlF4
k8h54qatEsuh88MdNX/cDHbjHOnrI/DfQqFOiauCCql5xPYKyskODo3Gtq9yYAnhHmxhfKZ7m+uH
sNossJF6P7iQku9wA8IRjxhpM9JSR/84lQiPbgQ/FsKsz8ytUp/TUc2Bnnv0NRIjDOkQFzDDCes+
hvFwSNsDXzakMnswHoyuntmL9ygCa7IAvxs53siuFjo04+sGNZCKmo5l2H2AlQP5K9yi+0WWTTYK
7v9joAgtj+TP/fTLsowMwyJO7j6y0uHGFcuuG0IMx0j8ROiIoXjNVBOVpeB2fsYbw3UhLBn2S7d1
oaPEPvatcv0icGhsib9vmyUZufryG6WlntCXGsfA+GgPX34THurulWEpPCHb+0TdewLcZVDNyAZJ
DB2l07kuah3VnnGPPYAGc6sOqqj/oRxfRNAXooR5q4h7HIVSauuIFkJp1U+EnS8W2B257pdzhPN8
7NE0acWA855D6L2y+r+gia49fLlby1g8H+iFityLPpDXVwXVnM5TBN/Cyy1ctVlkPl1XFEUqVZ2t
jVgKdARPsrR54IpZlvgKX0YFthfeKDWkEExARZl3h8o+kMP1rJDAzjZrzZmn3PhB1sZtcDkaHW+/
hoygq+l5YpEgM+MfdHQTkGVGmib5d0BgHeqgBrhGI8oHLpqM7ilUyxJqxIrUgd1NACPg4+a5QnXe
KhEl3umIK0ZUfq7m0jMTbNtduSAEOKU6fTDExyjmAjnl4cxKRvA5zrYmESakRmejNBx+wnbN/fWm
jGs4xRsPxRq9IdxeSRb/tXncx7NSDHe8DlNV6xRv4161s3m6dRdCNXrJD3UTAL+qwR25WgKpn5tW
dCkoIgFHEV9FAkmN4knSyPQKjIMNPcrR6yyaZeQRcGWeexCaNIjJ2hbDFSm64DxMAphqxbzQP6+L
OkrSquzpQRV794S93D5qUEQpK9VWxLYeZDa/QLyZvqxsTnVOFfvqLAYV+ry7sIkSm26KgreBesj3
NEJ05GTFi8JFl1GcJfx0zOSNzX0r3Ni3KNXEkCPBeLDL9qIrDEuBD5NjkqxMbE8j8Wsi8xor97oU
7WYLX6KLBdAQ1ZHfCmaGqgfTKXr0+VJd6kdXVbi9vFI7pQSIvgYr9B4wOPwRWeal3eEdSz3UQ2Pq
KKUcu3fF1+bEG901dJmY4iy1u0VtCyoIelUsFSRHfzut35i9hu4mDtHYhksBLLguNjtWtKsZU94E
MqHNBRDo7zJui4Y6gLENY6kfmNeNt8+6JSHTdU0oqOCnLsQMfAj02ehsBM0GkHhTH6xDmbi+64jE
kHLtHkZErO+MJnMzyawjAVq5eOHlb/QlXjc0Ndt+E+izXudkUdoPVKSbGMUyu7ae0yB17/uO0whP
Qp2mj5o+oMOVbMl9v/lwr6dSZpJOjzeZCqVEHitiIIEnuyxLV+WpYy2auJleruMoINCu4d9W5YYe
MqYEFTYfrVv3EcO4GXH/vbAIPKRTFdqMrcfHEcNS+6A0LmpTHBp9wdfcJvK84eLTlbEhgud0GRdx
buUgwRDXPgCTEcGM+j9nHpN90z9kkXvFDzTgCWArANsmWCXh6I+vDVDxAIGBDF2a1AGlOZoBvnkX
MI+lfb0Dqsf1CIXTY5Y7hH6ATibocRX7WKC/LKcNMplRD9NRQAr0MtBgZPQ5GHQINRNouAFdsS73
bxDXB/rf79Wf20g1K4Bh0VPr4k3BsbTqp+PMpKPWBbrC6X6CbRr8xSWrOC+eRZPNBi9890aEgedo
QwbhYXU82xHdPRM+YINDEznQWS+DZ50H/TeIic0itB67WQO1hSKOpXEVovYKKeU8e90QUJ/+SOGO
MyKRYJWrpWQCPPjFMBwsuNuaU5QVtvTNsMb9c3U62cbB0YMkY52RoB31bxAZBVfnRWkey34k6X0w
Sn70by86uFUygB0/yxqjhzpVvaHVOwm/7PpqI5jMlgJaPAn2c7fpv1FdprtKeu1bXNBP2X9xJZBt
SzIKIV4xMcGK8Q7Z5L1T9m4ksoZaCi6ToMM9/nEm8kPmEBGnkKGrlMHS6am9n+3QnZH+vYFx5xqQ
BrVWz9BqxBdIHucp6sfUMuBp6T6n5YF1iEzK9OxjfRD0Ndy51emq0GUTB3nbsMOGOuKIPqkgejW0
NIUa7iIrkpSN277hifXATJ7X8RTtv6VP4WWc8E4UsrrvZZHYw2IKFcHOQ/TyEmuRFrKj1g9kBgxy
qNYHOGgJpvC/0QYGrWnKANHOaoZV6cMp5QPvAaBpx+HEDMu5iy24FvDrbHnBOdtKpwIKBUKohQLk
cc/jMhqhvZ5ZYZtKaivjH31bMFYU4ct3XE0J9Ost9cU14szTUdmwKX+THD55toEapu4e2rBeX/KH
82yipMw8zIjZdrxnJwPNSeZK4vpJNbZvLtCm4er0/lK+BZ7If5OAX/Mlq5KpEnhS4THzIk1frse7
uYsnIfIc7O9Bm4S+6oRUguCEIo50Rkwlmju45hAfD57kahb0s8/JgGMKOcFzan+rbV7uawzzrZTZ
HmSL2mM8fi4kSDNFGo2WR8Em4KRyTNdVzjjoO/Jxmi8Mby8vQPDJeQWd3roaEdRpV3aqzrWAnPA3
G+UcEk1l1t6JqFKyubVdCmj2MJSNQKbcJCma7VuFHprXxbSXOujuJtT/aYdRJwP0ji4iSXSvRV3S
2vljvWARxope0BNUMEA07Scjw3kMdOvDXAv+QlS7PSsLD6kRheVSe0FwVimy+BDyHa2+7V5Hk1LY
05Cp6YPvk7bqLRjffikEH+6QIAaUosifqFsDIf10clCnzjKcCFkIqMvpOJ/NNs5/a6WHDFfc16ah
4XLyHue0Jc/lBOPHZaWC5i+k+BRWQ7jIJtOSnZmQiaDF7PpXcVb98QpqT3hu7CIUdDXFArYApQ73
vmuUX7gpGNP/rAaRT0uUeJ9H4ChCjqdWQOHM2MELRJjaL9BSDnUisOr3esfhgY/S5/J+8zPVXhMo
SVxESegUBB9XiQvm+ZC97qnnf6A92uSnfT5okRK44Hid1484+ehAixEy6mvTgfG7cGYHAcgYbPlR
kRzLMGoXHtjDbrKhqXJnJ5gC65xRbeUdbZSg+/ZG73IT1DxtqTl+yrrEyP1ObGZQBEmUt4VAhbtv
fTpvPXgvLkuhnU7qTYh/ZF3GkSXzomuGj+hmKOZzTS1ECNc8IX0qtoClyDR5NqNdJDEfiwZDXrxU
8hy686D4bKeLPJDJZDw2mwak2qtRUayuYIuk5jt/JoEY1E/oIuW9j3s3gGwzxzMMagLLclAHcV+h
LYm88+DbTpEZmXYskUbYK8Rqu+ttJT/A+QdxuvntmUZ1mLdLg0igkE1wWH2vFQu9fjhOj0Io+fNn
YgCtLv/VMNt5R/wrCyzHQiNgiYcRIbmG9kwA7Hdbcuiceg/Ve9nwDJvBUdK1+2eyCrmu+bPNQdQr
VpyyRmXbcBzomiYGUuplXFvHUCoUN3AQUiqHWxTETjDOysWOao8q87uCpxMRzp08B5Md3Gfyc6oD
5SVYMYWNNWNsm3qgZx4LvHHVlPIdPiYB0GSKVunx3XmeT6nY/YwBRLT0WyazcLTiOZghFhbZTDMY
7NKSbSrgJD39DzGspeekehxMIk5Zh/iAb02o6yULh72paz2LC0wPA9rX9umC/6Ynr7Zq+j4mFbQZ
sh+qFwFqjfJYXgOSOuvQ7pYCrtKsVRZ2UpMZXszcGN566/DY16ffEU5x1E/ySUBzEF9pCqXx7W2B
zZzMmmZPlWOsP4NK6kR64iYe825aidtLK0cUMJfhmXbTyN1/UDJsRLuT8Gr3QiL8aMw1vo/sjO4b
bbzME0BlvTMI6gIagtCO9PMcz3ySlytMVMrVcBd7+Y7IfllP/Q/SX4SnazfM+JgKFmRNAaBwO0Wa
i/PI0O5lscYGl5UUSwzDpKRDUF55fLBiV9zEi4b23wCMXLnQtwDhlK6Qdg8Mj+g/Dqqo5Qm0H7mI
ElNkf+fZ+BmMBUaxDcF8rNquyje7bMRmrpVYP4DeLSPdxqPA7FuWibfJ0RnvafYuVyzdIO5PT7fF
lyykGKJFZH0iKEwkxhOrPJrZJp1ikvCTRaQPJ+5rkNFJunns9+9pKP5ailV80GUIXY5JlZR8A2Nw
foHWvg+Y+EKlxXorFX9rEo+MJaD0L+jKhdyO0zjvuq+TlYOtxNcYTgfFG0X9y6QS2o37JfohX/ER
cJhdX0D/2dlyt7gNU4I0ggPIZuhNxyAY/sYzwy2WkKipiSu4PuMUhU/uLQJi8qr09eNleoh3XfMb
QE87MN7URKakaOGUEA563EddFWT5093gbGO3kZojWWTeUlX5kUBmnLuun2dEptuXgLTGAtX0MzYl
+P8HwbpOYC+TQtHQnd78X7Dbkxk/urwKqgDQ0kfrm/EZa8AUxJo8waJ5i4+aW4GGX8vTUVLU+pfz
IzHcR9cmKiUbzdzCG6PX15IimFyxefftxIK0WCuOYVgsR4UpQA5OLFGy7qTtJCrxm8hGcAapxBCH
5Xw6yu+7zglKhglnMLY8qphzEcEvu05Y7zSQS+Lnu/Oaiay+mkbYiblTGtAO3wz6BtzcWHqAIVF8
GpXYv6KvIa863rBZAjlSMCoMR6oU2UFVRlCUmNj72Xckb5w+v2S48ivxltUF4R2dD33Ka5PmKU8F
FpA4E2S5qAXsK4ZAIiqCAvVJTNNXIQz/7+ZTb1p+Ut5QF0aePTVc3w/LiK9U6DDPqoxifVMVwHwT
5LXjD7lIR9SFQ1Y24tKp54O2h2kg/vkp0gCgr6kSOwC2aBkls06eSbqg2JcU3Zkqsys+1Al5bruf
2rky+oQa9Iudke2BMs8Zka8rKZLoks854CODLfyrbJEzgBNw2TLLQJ+8lsf1MWicaJPTE7l5Ty6L
//rulr1ylseR2t5+A276q8PSqmLFL8n51X4rMVX4XBbDV3FNyvFbWAnrRTBuddEX4TKlYItXa7iw
32C7gIF9Y+KM0Axh6rZC1mFYD4OldXV3VXZxZwwREdnObUM0CEKR5Ercdm3MfCQimsqR8kGXt48H
LxP1e9VPaKbGQ90uySvIcToiTLw+rygLfLwujPAwrXwzRrRuUF8Up0m/ILqwb/BSLAgaRFhLKZ6c
hE67a9kDZlOFNP/XJcLc29dXG2AvJW4RqtsACBBDdqecRaDhxR9t/HUKghwljttZ4ettVuR04oA3
TWLhxfZmo+6ttWNHY3r8ONuZIHPJdJeczHSlEsM+vJVYzqBwBRhIzkoO/NxDgjXY2USpLFsmarfi
KFNdb594UTp5tS1c+wAoJRr/ngh41EvTHbI8dIhs/wq/DeilrO19X0xIuwkB9OZWwET9lgVp/awn
OiIV/OiWxr/l5SyIayIjxZD1IEJ/o4MzLsNO6Dals1LB8E5VGf0Uz5ae8Uqlsuwxx1BQPlPiIvy4
KUH5oWeNK0MbxptSpFp+ntjpdVFjFmSyyVuwh7WwW6DAsdH9gME/xROfu3b9gWjZPyuf5PgPNPgY
8zmsNumFYDgVnzwNW6+otNq01KRA+sSNUcdz6tuSY6lOLdmu5NmmSFTDFdgCuMkBhTfuvbBr5rsM
Pt20bn/PB49K6l1pJjyTV7FUDUISLegbodLRyyECLbtxyAf0oalIsJd99d5SVg522yLYjjig+Xv2
huvyEB8vrIvO1VRw2Go/NBjcVdznyRCdvyfUqQzmcGSmidK3iPQFBC3UCGFXJqNfDn3AP/Cd5yVB
cMRgr1z91SeXaH8j8M4lS+/+s9qPGY5rm8kM7sLsNAiUMAFu1gemN/LtXw4ZhUdmRD1abKD65Tfs
R060JxquDkRAOXku+/XW6duKqEjqTGiHj2K7t9N7I6ry3X7dZkgW6EdF9MpZmLX3BSkY5kiOuZAV
BUtOXZKWTnALwxeaiYyEs2e675D1czF6H+ePONC6KSjtYZHk8pcdd3A1ClJAXBccenqghmqKktu8
vM0PkNnqXpypbGCDCsGdpSEZurKZWvoNQwvn3EJKwUJjwQ/KrJrNMDO+VPuGD8upA3tS9xgY1VJ4
XHWBoSjl2WVjQ2JIgZXQgVGYuqbCYc6qA7qj70N8aEaaIZ/936FUBqtG/Q7s5HiYvDOhOnf9nyYA
QyO+KGaLeiObgIFxppcLvucTQ4T3mzgsHsLa7HyBoifPFHGsocLvLZ+Z7UC+3liT4jMjRJAEH0/A
0Rtt7tPYGYniEE9JdwcIVKMNqs12wmwyKvdKQ0djh8But4+VgipwyA8gpJGWIgOeAsF4hHd9l7oY
3dR+gjdNQKKId/iFC8Mt2B/zSHxqdD96MVcbML23GZ9uTz9D3qDqripEoQxC4vC/RTgOKiSFx+o3
roz9dpvqK6SJwwfbLoGOpQkpqf/qHVaVet+yUkoikHFoXOUV2z1GjEyITQZdl+QgxuIbfvbuEdTm
2CR8n0jv77sUgnuGuQY8lUC6mPoSoXZRU4cPU5lEItNAV26VFx0MupU9eQWT0gzZbiNu9qmAnkrs
8litjMmg/tqVyyeELGGpQ7alJiwfmhgVwue/v1gxsmgEhW4lrI9jAwKNArScTqSgKCbgQxuAfa5e
h4i0821/2dqXn5y2rpkLLzdcl2PoHSLSQZc/Kb9BqZLJ3at4BWkxK/748v9rPdjVaT3Vcqi1QRhl
TCSao/qjCDK4IP9v55eqESrfwx39ZNnAfQaMQQ1ng3+juK9laE6bpwNfrtMTJFeoABo0W45HSx1R
xy5LZccyZ+LQ6ZANmd7oeLBMgDJU05KRRfqunX0Gg8K21EnO1u7kWagtifHLiLIiHgx+a6Z9G4FG
9sMm8yubMDoBODoVk0Jdtimeq8gBg6hvHtbMU1x2kSRCwd2RWCcYKhtqSlnq/Lx/Jfar9Vo3EYs3
7RHwBnsvf5kvj1e+hxKviV2io1pcQGUvqT+8VOfY9qo5tWIXzEeLSxHXvkLjLerkcrla2+SJqguE
E27FkRyHrNS6qSqLCKzjiaCP16xg3gaQtr4fvLqChK2SA/QS4+B9VQ29wkW+ftOgidXn4cuM8lc0
ix7flzJhXgMHzr71PJarX09lSh3m/Jk/HsA2BcjqixaG6539hRta2BZc1zoodDHRNeCb1jiv5UUi
ic3mqTGfbnqc6KzwouypkWXR1yWgbyww2omyk/opfym4W4QuwNLGZoMlsfBFECMvEioIX7rlpXsK
xEGmCoG3pyzizwM5pXpe20eNlkNLt/OEX7N3LGDiTHiL6zvkrRhf/xb+ucIHlBN7I1ZlK/X13vDJ
oeqF701LoeaSdZ80iOPtkEQLUnDticiKtvsydwIpLIzalpN6KkHsKvVHatVZUWTMyrM5IAV0cMRd
wScc0jY2uFvJhYd0mCA7ZXc2X/TY5kXQJ92/VFGxzn/HJeLw5SjD79h7tjpytOErneGTPhSXGSxP
Y4FcJEHJCiLAo9auYqigcNCF4KbeLM+1vwGpUHbNFW0zicAw3mPrUHkvYRXI1wQ3FC2oN0L1ybVr
oaI6xRqBZ6rZ6ToFNjBckHo0os6yLKr1pVC8QVOCcAFqLOByg9C2Uw1nV0ne6L7xCQCV4GsofNEw
REI73pv+ou1/7goWjGXOdXh+ASnmqW5tLn4bKoaUu6u3mZt/A/4BZgBUxJ+ymfPr5dXO5wxloQD6
4SgdnLOqdUGWP7rvuOIm25Z+dbrVjI5Z7D06BIQCMwLyc/Gop002xPIs7PCMt8Sw2Tr9wWwvQ34b
Y3BWgsjEmgJcZW6yhQEi661M7WsdjAh3pPJ1eCr6nlAR3wZ7v4Y75UzLe0rNOTniUeo+X+oJgVLa
mLY4HFikK7CpYnJLb4oq8v3N/KHA0oWHqdVKuwpO/EbWNVumG8KdEKXOidvNP6qq8rB7Pp2M6keU
viqWQprsimeDN58d/icLNEbkDQwZhB51ul3nosVyvzcuBtaVaPqxxcVA+D5m2GUUHq9sNAysRaGt
fgQwnsrHz1o+Eghm4xTHfgga0k3UkqPAV04yGj6WOYU+FXAqPCMHZFg3Y0ptxqnB4+kM8MPzVxhi
1FegXd2HFZpr5lsOxF1vlCZLb5pcP6IS8+zrorLwxeGLLOzYysMr1+rY56791iV0tJ7zhRvCCsnL
a8BBb4YQVdF0Sk4TXuYIqAegGtDa3XLaKJhxHqQstyHJRElG++bUX2k22p4ehegFDsTmW2zMnskX
dEjsnDFthPPdyk2pj6r6aFxUJi6SgYdtScrSJXCOJocyAb1HF+NkRBNMc8gOOixVwCuQ+qcn4cJn
AXbuMGu9KgU0r/0GI9i21KI+UjeHB67SjpCi3n0FbvuktMdeATw3xK+haVH7e5p64F7fy2s1AknZ
/jc3/vQb4v/leD4hxmhNc9w8cQjLCWKA50IaFxM23F+ilutsJvYNZS1XacWfDMQp1KO3jX7ejlSR
lr9MF5eyphkkqMlPI0nzwW626a6+GIa0wMaJXEfYd/2iqIiQD8Sd2m0EzZNeip1VxPZbA7yz9rDb
km0cQHlj/WFbSaRmPY4F+zDNixDYsVZ0iqchfaSsEpUViF9slQ1llRjtxuMryOUWmBZcTzKWGpNX
VmCZT2vG4iM6nOpijZzZUY1nxbf1W47j7Vl+7wTcAluolftF3iOc6Ni1Gz7Gkvj6f83UdPKJq5KD
QCheHOWrBNVgXMfv/UpQhHdfpwWDm2t/pj9dPDln0KEzSrnAsKb5jCpJ8/v1dZXmoUfNr0ppsQE6
GSYtaI1vn6o3l9tO3o4MWiJlgnNlaaz6ic0P04eXmlOetYO+Jn9gVSZ8qDI2TBJOM7aG3V+FnS/4
bPHcW7pxmcOqycPBTba8KdxiCvlAwPbIx7rKUz9vwmz1rmLgswbhf3YFSzlWnFhZmt2jrNlixDGW
8eBohLTELt1ZxO0jekyuMY+IRJLal9qKHgc6dK2XPuqA3MxfDp6bOiKNYyYZmqLhKAuCqaBZhzw8
sF1mCIvvgGxp4qmUqqrk7uqS7DoxIctELUXkXs9sPBoDxOdo3wReq9xE/GZgZBwR/XV6c5sL+jN2
mfCg7TLvkBT+lsX1MedMDoLX56Q9gEIu+RWID7fj7mGVoVPTp8FAC7J1C82ngXPNfk4XZU0cIpxD
VT31IvFWHLP0cWZKZBQ3GcNnLzAM83UA3fic81mMOUWMJo9FamY6jZPYLrUfeuYVh3b2MFY6sIeX
B8zFZ+znDarlKpGQzkN7GuFkoyHvca3V/Q3pSWRtnCAmHdXk2RpXTkYF3D+NeX6IY1gHjVfHMNAU
XrH4oLDUGgqD1dYQO1ZgpewjBLx68jsunKJ4H2pFrcfd8xcuPTuZae7Y4Pddk+5esUZZ9zhFsjkR
Jnfo00c/3adS397N1gW3Le2heLe5yWjMl7qE1yLDJJBeUigQm5AoD+tO40u0vmO+bWwDXsitEGvZ
yyySgG4wkMHO3O8RMdv+m5VVm7oPD35uL81a0qO14qn6rdcpDkx9jokBy/LZZxP4BV4c7Xi+bMjW
iEzNPwEOIuX6Aj7j56Jq3ptwWTT5USPKJ9c3YWTz3O/kAYcWSxTbqllT6/rMT33SPFms9SWB8bqh
vDQ86ZUXpjx/skijgOCkik32jvze/E8DlGcTGgtMnDh2XJ7D4DrKYKp/+CIuEhpGiFcxO4/tTcEf
Q6Pe40BCBuChltu5svA2GdGYE+gmnEwdsPeXMk5YtjqX5qXKfq4ie973iU8z/8PqvwZBghNKMzs7
70jkkCCWptDpKUG2QAqZcQlUDDUc1uL2EReCnmsPCaumZzBWe97B/1nIowxtgImB0wIbJi94hfit
VefevEisdhpElP8mUF+fe6UI3f43NlzV7a/OttdME0A7neuFfMhoEeh2Kfuj6ZrUDgnIVhOV0Vqp
JhAwhxVnN1KLa0q8jVz9Sf5xwwuFIm4Yvnr5+MOA6nHpaGBMeStRseDpzYulItmPKNq9ZsDwui75
7ilUAunbugUGG4213UdaVLqWENPBuEAktB1u3/n1TIyOuDso1hU0j+7jNq/dvgCUOfFMIo9Cwnxi
WwDzz9/3iFNTT2LBaebrHrEuYTeCVqm6MoS5QxH8pMuVYOtPUaZFPmKbIXM/3tUYJL2EyM+l3VNE
6TXFbGAsL+DvE9vRuOBngbFUQEqWe22TFz6AD/ewN2wRO6jUdhGwnCGgmdKAaBkwmox4H40nGjuT
zM767llw/1I1B0C94JCA+nhbiVLjb4aeQalQy3qXHH9w9i7DLw52m89v+y7wROztBDSLCK13GaDx
CVfuNfY2UNM/5Hvsgj4cCreFrIJ5zfnFUtKENI1u0WosSKFBD+obW2HO9L3ExVRfrvgHjRj2FHYF
kRauLPJNJ/0Q0MoPKD+WzP0uIjD51rZzB/QR2jdX1Swu2qCHiz9DSsA0RuMf2O/Vo3theIlreaHS
IIpJiqu/SvUe50lFG2lBW6fvir7opic1k5b53gUmFWUvwAuN7tsb5uSvleEcDHJmZxr/pyMOmIeI
jFmn607a4Lx0GILI07wVuFyyZn1oReB3F6x9ikSTkYSN8HRORl+MuX60BXzsd9zdmJrYuC15WBtA
ABL8bComZnL1pW/olzkqh+HkHdOoGl6rvXg4BHcAjFCZhr4RrkoZ0IwBUGgejmDrNHumgaQNcp9L
2EH6zT+OO4LQAkmF7FmJAMkn5+DYYuxB3PT2n/dfVumVJOSAOn5BVkGmQbwKXgwb+fF5B18h1qHq
5MHuOieTI4KMDM5KRtadAKVTpeEUlLOF/ylL1aA73+aEtgjifdG2ulAcyLun55Ns4bZuk3erVK/Q
S13/7Fy9Lk8NbFf01NTWvpCBNhcrFSRXU3Dmwr9fNTDUDxKfC1cYR/6GX+iUNERTRewM3zcNCmvt
/c2srtt4Rz3G2u2HkFtikg0iI9gKHgWG0wILCan8hxAL+BXHcdELWqxtIhW2e3TwQFuvjzFgpsk4
qbUad953sCDNSLOzogNPxkpliYb3FEbrDdKNkXiCHJFJSPzb3T4eM+BtZJbLruV1dtvXVw0kd1mK
QJeTFk6U1rDfK4Xrpn7mC68pl3AP9z/Iu6kyzcdGc74YUdtbviSBhVOKeayy2aVpuGG52iaeiNxq
rXUYSq54yp0KghU60f4iogasSRI6v7FrkKBH3IG5nII3nlhp2/jtETdYrQgT5OmJ5k4OCOsNqx75
1uZhWy/cmprkrcIgaTKDTaBmqphfHvL7NNk/ObAUHYkA5+W7KsgHi5u0z2v9bvRyTx9AxH6ihY9n
Lg2Sf609kxsny3jnRD7lybMy+nciS/yQ+opR74vndpEAWifZQGaG2clnGVmJtl8ESzgAkfazOmdA
bcbWC9vXhKZG+UIAePOkNSub5DXsxwmfMnl5O72fxZucW6h3QBCErJO2aOOqrxeVMEpaXaioxmYk
efhp/aWqCeHG9B4Mmku2N7SynogNB6/Yu2rCK2aw9Uy2Aha7WStNjmvChfDwjkekaYU2/L5YoB/u
M0dJYw4rbHBQHOFhzuIr4Dd3RxbSBgyTuL2IO0iNmUBfFNHBodPNvxveP5E5G6eYy2uSCW3Mg5Xi
o3Yzn8hqcsqps1v+dzCecfhIGS0w8AJeL9coCZRrD7wri6WhaxP/mCLLXISaj+qGaJhZHZjdApBz
SfgskcbGAUogUKboKAI6yNPdI+oBIGJli9+VWT58jkSwE6z3BgXb7VCKrLIblzyZrSL9/DbNaM99
g+nPGxn/uAGmLu6PswNdKAa8okb3WDtCh590NvGwHL261ppj2kGRb1ThNi29wQKTgPIl25z11/mG
PXpkqO3TDbDx5gU61Y5nl2WhrDLAwLtEa7ill6byIFJW7tZJci1HO4xEskTlYf6CCs3jd8ZUC57q
/3qOsYqVu42T8wtgkA5W1aate2qDEcTw2AggMPIh1qGeP2flD3FCJ/6Rnf60j8kHnbpACf9/3hGt
Y20ieUETtBgfPgSvqG2F0ESG245hHtsDzdXTg/7U5z4ZtnsOYYVyKoUVG8C7LGAmG8SRpgFRoQ01
+30KImXiOVn7AQht1pkN2u7aD0Lbk1PNo9k4D22eKOu+OlV9iEIK8d+LzvHHR0YNc1akPaVSzpqp
vvTNjAMGtrwyi2XObIykNrx1pubMfVpYeh3wJ5m2DTS34P5vHajX8RaJ75wFcdLT5nF6lPnzHlvS
XxmFJOti1GR6ma+uxaTnFdglj7Qi8fW3VbAgvd6uW7QuwzbsUAGxFUTxoMWFcA+UjGL1tmZVv/cf
V2rAwiNEmQHGZFv1XACt4NJE7XytjYysOg8OGq0Z3QSdIWQux0qqJgVLZLmeSeCdd4uQMABIB8dq
swMtxeCXuRS6mMge10Gq5F4dl5+6sArsn/1nkpegm3nidEZfVVrS2siSOBkBsiZjUqD7uZVP/V/t
DeTlqL4gyvti6VR5ZUiQ2XblgW82tNgc9UTrYsUsW7gkPo+iBGhTfsR584b5fumN1JpoL//i7KjC
QDFspiMs7vK5DBHIqATo6kiGWvSO06p0qk1lvBcJ6IYfokZraHdFvwJLjgR4jsVQ1YuED1Q492/U
7jy/snitmX0HLfluP9gOYbaCq79U9oeyqbvdumMcTkuYuXwqhkCV93+E/+ayNk3p8fjoqERrciPN
NolWSJg9hfe2GjWhflObkIv+KBhhpk2Dqvz0QBXsOgRSYNn1MJaOXg/0AkjFDiLkFmLhDE9JomPk
8rRHw6rRyyLGJoI0jnMR+T4bqiOcv4IDU5cnp9Mwo6Tq/13vfeElosqrUYjAVZFAVpumL4dkWuCW
nuRuKxdITMwETyQOp4lH/H1nDGnKrVMpvSLFHCuB+019luOu3uaBzkmQbumIBThmmhJFVXudLX7l
8YUXO+1AtqikM0+ygYheX98jfFhwEHzJJVs6nviQzcV4qNYNYu+EQzJpq1Nz9eAGYC7omVJhnnbw
36YBp9yesrgODtHv/THs+xNaRUQ9JTFEt8ybNHt+FlpEZ43176zOnHw+xG+UHaO0AZVDlKSu6L7Q
G8WKsId5VCc4cV3zMMrK2X3mg9cUlwKkwZmLyolDaEEpznKGmr3Gtqrqp6EcyPC2FW1Gdvx4Hm+2
B/mVu+LlPxU0o4R9KAWqNWwh56ypeA0q/3yLtZ1fF3R5qtFVMVIUhhyzLAqb2BK6xq9YdJyLnNZi
2X3FpHtKkWkEhny2+zvi3zUXGxuw7fBzsk8Uj6qD38WJ2qh0Bz1TF9bYFMUgaKAt2M6lt3ktbIkJ
+8joI3kwTFQ0i2+cmYdQCNajSvVWqvI34PA5cCr0ypTRn3uHqhLoqNtyBsNIR85g3vQH5O4bTtTP
4Hg3sJXyao4cEFwTW3SZ1DY2BkAE0jb9ZaNGIpdi6R8OXTDJu3Hh8QTO6iV/lSTTk0MX25MU8Ms/
oSnEhVzFtH/EnAmuP4kjQ/MVk3YP/8vxclWYOh95JDGSQIvDEQq7m15eozU+6rxkVUxTYObkR/ec
Nd2Q0fdnPQVBrdDHSf6OwwstekjsD69xVro2jGfpuQDXmlHAFBp+SW0hQWvkt9GaGyxieABbsQO3
LsP9IaBSBcYEaFyH6cjK0ETl0H8wqRndYCy/C+nssvomWuxrOo06UTdjwIA5UAPYDnRUAxLIzIiH
xcPrEKvK8sLC1dtoxChWLZqvLYrPFqYNwIDY0qVUDmu69OJF3WlxaZ9sl+icR+TdZxqUiUsvpoNd
a8sF2cVku54ohaUvOXECEFz3nqxUIfy5cWHCB+dKC980cJvh+dUb8QoCWRSMFjUe+rxbGXjcPoTr
9CW6U6cQnp/854ZoPJ3iyAcpvRatJxX4EkYFX+8V65K9sAUC3Px6ikIdCIynAayOOawIp9qS4v9h
7SgrcY2GYzYazWw5MKBoe+vdVVOFmcMl9zBzOhCQT/bdBvjWYgzY7MQQCuZvpJDK/xIlwqQVC/sG
IcY7isvHgxFUyLlzWxKG+daI0Tkcq6ElbZ6rOaE/NAUvLDvm6thLks7GtJ5K0PwS22C+pdaOd4Gy
bnldFHjIjjLKzRFA+R5DVEWLeJXbfEre/xzH20w4NqdQZnvoQEQBiETGJQTNpfGwWXyUxMA6Xjza
ptrYoopR5g2v6/HaYH7GFtXKzqCuwjmRtgeQ0FSdfY7U3obYvLIgNs6lKspgzswSA0w/ipfSNoOo
2T2uaA//QydAtyw2kuspeAFDgr3uNVSHodEpHUDsZ7s/phrvKviPOvScXBnpwtuGDbw20KSKbvYb
lMKrzdf9EtAaXuYDlbHdffmt9zMXN5eiHKbz0D97Sj4uB9AI3muQi88hIZZCuc8XAA5T9IKgeZE5
o8kpcONGke/HlF9YFuwfFtMWxII9t/rczratJW7GQceirj7usBl0QEP2TQk2/p3Z0RrTSimBC33z
qhd2iyvoSnV4TXit+rlMp2briSkGLfkC/GssC3SCnNKtV8di/Zp50o00QPqnAHKM2gzwsurdNlop
6DyVgXOg3CvWjUEx9WEAYYTlRzxLkw/Ll5cFqDeNokdfAN39t80dWvpHqFB+I/GNaDYwVcqNBNwm
A/bLz1lIyuAz2GjugH0jtc4G8sOnlKUK+PQM6vd/nBaQtXkF9LBbRWYvt9CRrj6nllaO04TMJ7By
f6OS26iEvu8GOco2MI2FozTeEf9NNH1vo3Ir4d/exbPJgiDR5p78eBFjunKkfTUZqTpC6bNkOtTL
dCTnEsigk0WZVsHyVvMVsZYtnQsMLrl8R+v7La6s4Rt/efIPwlZ3sulzPqwRlLwQ+bLjOZ4SEKpP
AkpdrKjpqByjTuMBA5/xDnGrE04ANv4kIUempSt5lXPdoQwlgW+0lc77Fk8Gcr20BEajHdduFR6/
6E9ccrnAAVyHBjXIHMjKOtuWyD9zEg9HK5Kqv9nKFfA0KagBi53FauPsgU5JFqvGAc/PlD7y/MgA
GIaKXKOzJWKmTWTaY4Dz/cpT9HWLkVewen/ajaP/hYINRpux9INKxXX336gbdlDcUIUklJw61m4X
aHQnY16TIceVNO5bQ7FE4JHQ7+8sS14Siq51Y511H/DT2n9FkIu6IpwfbHNFXRP+57BHvEHhiJHU
oA4mayGAULgCC9BwZIzpuOZF7bsubqJkotwD7fp1l5yzA/9pOC8TSIVNYH+H/TeInth9JudT41K0
lVqaGVF8DUC3PIxtRdQZpp6jKVnHorYIElBqaEJ3eHO1HaJjwoe4aFWhjWriC2WPWV9BMCnFeF8s
IkO+nG7AO3lxjX2oAQqODc/FJHVfoD4+em6eSHuYZ68PYvSYWimVhrTJxnzoASeta9ipidgz7EGV
uDQB46ZOSplkUkbKtXzuObLUoK++aqZ6lZdTeDEwRe+q3KdoYQ29TnSXQPjWGhV7Vd110xU7TA61
h0aHmXAfOwYzxCC4VCDoTtRW3/WkFMzIMrCNG9jCFCUDBDayA3arS39QkgskWQoINIFRSgTfy8Qu
LgDufx1ySVAExZ+xZpqUOQnPSMalSWUg5rVhholQ5wp2irzGvsJKLTOILBpOpTXMUEldALAiRoIp
YuaXC8G79P1JRLDQyxkRHOBjOZNv/8PoTXe0ZzO7Mxc7JXw5C5+SCcwyKLM1MCHddj9fV59nFW4H
hcguQYE2up6HykqUmaUEND3gNyddVhGlB/4uoQ/NyLhfoootiqjQsKhCc3HZKFncNOlSvTInFSM8
nY1YJfGWQk9LBCrS/tIMfFnG5BMBT0flR/H2ALdYssrCGey8GJ1G2pGUBoTTFm37e5QXlppjXCe5
vURx9L+QiWjYsBsetSWe9CZtFr9tPgOBBMxwxLDad9RSRdI1z8UVKCqzeHVP2elwr8TsDM37+8ZW
QJbxEitkymNTsyVjX3yd54dq253tVOQBSsR3Oupxrz11OoZbccxmGHd3HHqc3mWPMn8vNV8fuOSn
kFCm5VRkO9pk4hDFFpITMLQUyyVYzJXfCmvA5qbZQKoSIvz4w/bMX5uk2IQ6/OAvFZQZfZh5MT3R
OPbHvkgqV0HdjOjCo73WtCvmHTL4IAmadbmcRg5EHINh2p6lCWnyrSHEbPakh+7BkG5Gh9nAzX7W
x09+ofCwxROhO6P3JxDFWwD5aN6wnOW88tyVXrBhbOFKqUqvbi9jWvnfnwr/gklZabMEZAi4/lgE
EpfFKHGaEC0xi/TtI13eBwfySj2wGsW6a5g+XU2QyDx92tIo/fBLS9C/BPre+PJLg8qTETnttpsK
wZrtPYjKcTJbJIQKWPfi60DXXyGpXMWk/CoUrC/1h/q2OqdPJ9xx3zVd9g67tWAfsvP5S0ywq+QD
jugmF7RLB+idjbM/KosnNRg4OpeMmpAz4K28DLC7/HsUu6ABVgmk1PE21bdleDTnMaB0MRA/AD/7
9vBPRchPQw9/37UFDcdIVF0pMGxr7RgQKApRIhuqw/GbIzHWjfbkDL28/cbg2qX2wqz0/NSVtder
oxC8Kabebq5AaFA7XkjNrNYvKFtXSVz8mmneOcxcifD/u5Jy8O+4IGegnND+sQgE6N8LDYsEATwT
JxwRLkThZiMvN+o7NJQHFATCKzLIYLlhFiBGh1aPrmh7Vw54KKnv9I5egcWIs42sI9ltT6MaP1+W
2JOLekr/utu1jjGLCOJ+q1JfZya5774rBUqChPyvbQwxrGYQ/Gi870+HQFU4JPPcEy1T9+nmxRo6
8+DfPeEZPgPZzUvP09fUk0RdTq5KJSHXivhHBSG4XbeFpA8T+6G+y9JuyG9LUNV/ttoU2pLGv7O7
ZE7mfvokefeSVvERLaDvJ2wTgGw1V3qgRmMKBsPO6D3XcwCJI3Bu0h5Sx0VYABtlIY4ESMXSZf3U
H1MSXBRwsgEicwicM4F9fD96doIhZIOcPb5LupuBxAc7O76F5cm8WIB+EIHh9NL9dc3Ld5c0kyfh
NtAITQuHYxbk/pMhPKi78ZHcDaw56LYpDJLZHLVT/EDbmPq+SlF+L5+7U1HeCrMg/Bu7rC7VX+8h
/CEOpJIPwo61q3VpuQupnojlEEQ/++k6DbzExNM3WFkVwagOCFioPb3GIQDf5oeJktuPXjdu/Dfm
YpF2yhHJAT8n8fnX765rhjfthp4R+ejz7WaJ4m9qcoy/w/DKcF8nqgjHVjLIS+E2Rz+7IIONUUBS
2jSVTpd81f0ubGo9BBtJg9UUybzl4R2uL9hOkLZb1tBT1y9oTgK6ndsNkQ8bnFnn3eO2r8ltvHAd
0rJv90jnoyisaWKb44llhEkJgzaKPAoMdvkHg/2SfpCJ7CBAMKlqXRCBwfN7+ezM/7mIA2oRws5x
pit4UrvegFRl554bCYcOKdEp10Ir3cnVOJnD1vgxGoDTZX+Rd3zzJM9RXs6bj8b8bwiEqqEkuPYE
SINF95njfzB+kJATy9TnwtZDKBNXw9GH4X0aQqQfPLQZXi8g9KV5wQDmn0Bxp7H2Tihsmiv54uga
ftaRynxdW6wCpPoZj7VniezR8anoUmee3jWWzsokQZmKV9zDZCXuj/Gm9Pcmma6mSQhm/RjxNZKV
SpNhZfB5dr8RisjPIn4QWDAbSarJDbtSdopccMGUFfVfaCo2Mdt3rKEd238yUkanaf7pIV1EcI6a
l+Z5MaBlj+dLzpc0fUgjOsMI6e5naLSUaxFsPX1X2CnyHRjoXsj29BrDODD+K6yK8alPxWO1KEs1
MJjGwouTyAhyRHX319qEXtrOuHyofiQk9rXCsLg1TayyS+U3AjHQsBiYoXDIeiMb8qADfaIvLYVf
9AkvDfnJtMtTH4HSsKo6rxb18jisIbVsgX2gQF5bG+yUfIGBknO5XwwoMihdnwC4R4Y+WjNcVpgD
2y7gA9drHFjZEOmxJMj8nQmTdCIEjhymbF+KGBHgaMxKacTMxI6or7Cz1OG1FgSSFLNmjaFLO+p/
F1MFM/qp7iln1/3+QWy7oOO3AaWMYrsLZrbbJajODiBuESUIxUAoBsAEXVoneOIs658lLYc+LBVL
Pu/p5Tf9cajaCBidOOXPm9GjZ/WpZ9Mo7Ka1QvFg/JYcm3ryqdLzZgqFfvjw5xBdBvboeAgzfiL1
PNanPPYKzkm7M1Oy+796yb45XcBE1pBeJ1b44S+NAro08u3EYPmcJUmdY0a1LTkjKSGzwYOOM1ZM
DOXVeKSVCm5GMxNymg9xLYH22k6PKhnza+ipzfu9WdRysiE687pbky2y+ns1I1SQjQcWQacPaJ84
nzv+QQCI1XTIQToFHjZI2sid8y3I34PNWW+5Hd+X08oL7+y8UCMqAhlwmMSWzZZIUVyB9DVhQ62T
PdYodpqloiv+OjVqmn4i4+SD+5OjaZ2Y/4th1WPUtZ7atYy2VLpjoTRAnQVcBoSEEhKZHf3YPiDT
I6TCfEUbikYkwX6NFvu0jFr5C7V2rm3UQyBuoTxyIofbQibXjdIBXniG8W0JFd6qUYCH9Y/YVkqv
rgr2sfSE2w0HOfIcsFMBwS2EbgEVXs8/Ini2iPrwa46SHecAOPE46lm5UkAlbhtlE5PEc1KnYCT5
VUfqMNFrNOk+vDrrDGlvvtpsXbYh/kRgR7Tw/YOn81EfleECF5CpHisvu3KMcIt8bfb2Y0Gr2S64
UnllrAkf85/0PYrzjwkDb38t6HOICRuXrj37t4kLvLfrZRZqSKaWAE2oCA1k6AbIZCLr6HWKKA8d
thFcXVuJ/MFBTiaNm/MG3cfUrNn09CQPvcWuK4mVxVwYuenyfMyUkeBy2NZLX+v1K94PSEoBGIGQ
B+bLeb1oaHO7GNr0DKrHFL0o2v73Yio917CrhnKfu6nPoaBhXperG+tQ4Gm7s3ooBS5zoDrx3VkI
qmxulX3zvEQO0eVgdj7AuVVsQIJKnJ9+hnq8F6dqlXcsxWUEErPk9e6VW2Hyii6J8noGzq0zvwuB
Ev259LlU3OqJimxfosS49ht/oyVbgblCT3jnCd94VfBcRxrr2NRGW+WkF7w/xxRDylsITjUqrjBw
5H4g+YMFE/jISz2keZXEhY6/w+nbFWyg/ELwodkxlhOJHwlHP2XYxLgg+HAo2RJyXmUewHrMo6Sr
Ut0gfu02Qe+B4vQY1HOZYqNXGzF9V3Y/KYg11CFx5dNCjmeR9SFrBY0ATP5VfnK4Fhp5e0dUrM9l
n0J0JvTRMFWHl9vW25y6z+8Kb09LbWFJBbch5HGlFwAxvW31hxmRFSaaNLxdxoSwrT6g10UpQKiv
jK3cMdttFE/cpycUuHYKnoNilrtiSS0Cl7xwOGm2d0GybJDBsP+NIG3vVfPAWIbhP6adaGTV2EfH
0/3gMiDVfANQ3iB50kphMkBVAR10TtoJmRLwZf6mh8tQBRB2EtKmKgzIuRNybIGJCno+aWikmm0J
R2cbeCZ4RsfqKF3KFQ5YbzLdwW/M+/p/g3Ao7CfuTYWaNElO1TJyHuIY+fVT15Xtks1P/6GQ5L5L
RpVF1JWilvRwxSXIpHzwTzAWSquVO4JwG0qLs3nsQFhCoWCY4tVavccBldW7SJdsgSJwnuEwg1UB
SatLDHLVtBnc7Lg/03DJ/C/4+TsChK0/ZKrZ9mbT6mHJVjpz9Wz5QlbmiWsm3Td2yPc24IbPbJGl
D+HMby9KRNWdJSfMalFkMaw8bASxLMIW4Ce1sJaqg11OnLtXxM7YzpENmjbHZEMSrpraOtDgdix1
d7mm/2v51+Cgg12SoCt7Vpe7El3WwA6NB6nwz+yl+6jhNyPh7q4upGG+qHPerkki9+CYRHnUuUTg
Upw8k8QuXVymo73gitbBA6TVzzydmYP3W89puXS/FmL1TG/HDCeXWeCDuxWpEdHgLVY8xzD+iTzc
4/qZXo7v2ChaGfnUsIzmZdB/svADSCg8OE5hYg5DFqMQvHIus3M3Jup+ZTHiRnShfp+wy6/Xj6XX
J3nThIYzhknYXGH3rBMiBjQAmGthbwO+5NBZDphBH2cBb5flLX7D2aL/biqmelPqkERDjk/Uulnc
bHIsuVmW7ApB7Xq0sZzRrDyPo6KFBU5z6DfAG1b8lprbMJqIMvODbN+NWMOp5ygCZJetQyYezQiB
GmA9rVLoOK/Dmc2SEZmLLABGNwMp2n8CyhSytkKcQAmYBfrco9CT4Y2Dz7DEANeAf6YfaTDIR+cT
hef2NVPM3T1CdMEfkhHLjLzTPHsePJmDzAbKEAr3GdtdsZlV+zJTWBRBFKNoLBH/2YvlOvaDxbHQ
9V2gdgcyGrWW8W92KNwa+rx6XKaLoMtc19RT6/vQwHfQLssAfnbl7k1thgiLsza1hvcbbXQQ2LYb
GTph3Ki2d5wFAV/2hMHD8rpMkHK0TS7wM99C8cOq9qMv46qqKQn0h424hYpklZuzXbysypiANKmh
ORZf/L9FaBueUyqMQCT/pwBITg40Im5cEfzFA5WZwpEl2n3u0kVwdVXagTZVL7YkeX7YCzaxiuht
8DGSv7rn5Uqr09elOBYt1JanBZLIOtZ1OdQi2nHL4GBjVhxs1865P/Tzzv32uoooPyrKOAdS+/oQ
SG6XWyu+6kTYXzT7sCOQ+IUG7AmqwOwK5mJmnNjX3HOlurJGiSeLv771+R36/seNBRBjROtUV2uW
NrcJaWf7zIAY3aplCStQ773B50cqjlfjze1JS47wtozDAyBvMaUjtjCpM/CIqJxUNLQCMbV45jhM
54mo4RRWKIoZ+DP2hk1KqNSmjoogoQgI1BhT9s8TtBgs/fKUiWOzTt2joAOqbEPZS0WaeInxQ1zB
zTxcnaSEfWBzfOJ/+7NcRp1zwwBNT/pwD2Uig7bXh6UQq9YCtDSfR2IviS2bsGNp5o3E3UJ4NH8P
9eJLK4yJG20aYnh3tMzXs16WcgXMy3cDqnE03a1x32zQs8ziCRZZrnFpX8klCPTH7EN89VDxugGv
sAU/lYuSgZJPKxGsk2M0i/6ey2wpstHqPIqVNZDP3O6EwQYjPyw4eWA584ZnkjhwUT/yt6nFIMfQ
WFrL/CsSKBNX6Th7zQNMHjqivz+tPinQ/odEYDxYRrreyDpQJ0qBgSbSWi2RT5bvJbJxnoHJAfK7
muXwbOqHVaQ9VaoYoXT6JU++0I2LdWEE27sWoKiJK5HlvF8wKb0+VzabY8bAhQ4zfCqf5E6Up2A0
g2bL3gC3K2L9j8a3+2pjr/NvQSuTUXSew5ikHL5L/zfcFR57ra0qdphpFSpHm/XuvpUyspy03GoD
sTVIv4CZKL9phKHQ8rRl2nC0bIlteI3C9MJF1+bqh/ILoayXs2o2opB6QJxUrfzwuJiy3fkAHRm5
qRDnexTBntDB2jgyKcVc908yQovcCfyglV1bUQTSYfCxvHIhnr+qw7ybJlwyEjxFJKZfW93AZUWZ
B25Fh7SYN8PlcUiMttOwL2nvIwS3GdiCi/LPK1B/FXBFwFkFabVD0TppMuL3c4TsxjHRIWhbLpCZ
eQSKEwd600jeghiGPVW5irjozrCOqiSXq5TDvzKyGYJMPbOI+/K9XsHKG3H4Cno/tNtVDowiySjR
KJ+7LyIkjwuA17XPNdzRDOR8yCrz4sgST6MW6EsMPAwl+Jbbcj8f7IpvYE0hcGi+E/+6HIrHxqIK
bfkjU2UbqkbuabdYWOn35X4p2rH/nsqXT8dQLpfjm5jICEiT9oKmkLpPfpTIc3M5UQT4gN+RuYKS
9fkp3o9Kq+zVauheb1E7o8IwwzO8SjQrR4fNYBNMK61SP5wfV9qfi2MytDy97gk8qiLU3hTsCOrA
EkgqFfAjWHjoKSJEkznZbmeZO7geX6GxfkWqFTOtOoAnQZLMn/3hqxJNsjzxsXx9N8QKMR8v0uyC
6UCJu51lpqPZcHRhhv28s9zgibOHiPygWZP9S4K5tWro7Km9tnH2W4TrW6e4InXG7UkwsMko+LSc
p/Ep6+DunC7XTIEnEvk4jpdFgKXnm89Bl936GZ0ces08anW7pyrHVdLYU26sKDYfuNskFFNLzCc2
hSz09UNtamsrhbgO84IdGj4fkIzGSwnVEeFtlufqkGeSPjIlVe09a1Ycfzc0Izs3TU6Q1KkAVZar
WlaX18uTidrjeORP9iTya0KE2T4/8KCZ+aq7iJ/ySfedEKUZM0dSYhiWUUvvuJpGlkrl+jxybQEh
1GNI/FsPeqvmPb/mridtV11J56S3zJ7yV3sxvoa6W9F3XPAQr1Y6IWLj3Mbad9NsWAz2MDWToY2T
K2bcqmtinYMt9sO0aCNpqDzW5Rrrr4LJyBp+yYxzbKNswl+KnqCanxPo+/RKdsY/vuhpXwr0YmKQ
AGB4rkYnAvL1pLXFct4alsdOv/oN4VmhCs8Z0NeBI2k2iFO0Fx2vdBkbmIlVy+dTTdXjWz/ObBm4
8RB4Hk5XcGBOzpgdlHji3oYoqfa+Qp+2pqVEoH8MjnZRvB/CWRI9ucelWhGT5w41SEri0oPMFH1M
gg5dZoAWUMcD5AlSfyhv7nCq/cc03bSWQ40RJwd7kDmE6sg0YDufF4wvYya6yOhYoenmq+B+mWDt
mgRyaqhT9y6Bg9LOCFvkD2TOUMgFa7Xzh9Jwm/mUwxhKsmx3tIwaQrVQGXjxko4QbIk1qOpNxVj+
1N7uLIHV8vXsoLx4jp+KN20yZre3m/8rjBQwOZWTTLSheWqtFk1w52teBaw3hjs6eNhwndn2WZ+A
bfnER6hZn+ylYSuKBXAOSvWshBANGu/mGtcVuUYQzJU9FLufJavs5Vt7Ob41DWFE0TYkswZeW8BH
qSr8uTpUVjpogb/qg3nm5A68KwLliLeuqvEDeYaRmHGZI76A3vAqDQyZCLgKb0lBtOxaTTZyKiis
TTq0J6mNuB5UNvu0Jr8jje916iyrfkbi2VjW2puRQCTh0OriTYhzhRu/ywexE796vQDHJizBFyAM
F1Jfrep1lfdsPkOsEUGomt8imhUIZiCEAQArEWwpSRvfhZskqsOeo+hSeFk45hwuwsbqmFCoPnk5
rGfKm90ahigF2kL9Z0CQ2lx2xKiw7Y+1TPSI2BAhWNsAZW5bxQ3wIrhjw2O+JOf2EyfVUzSSUWmu
VSXkZ5FAkocfGhtPEaBeBrDMmqBiKvFfaF0FR+XFW1uOza3u/td1jXyk8ASns9/fv+XfY3SzqIvm
U2lOO54YCd4NVV7hfKBLlM3PbjFBAPR5+eIgjOTALqXnM3qoVCDOlkG1e2bgIlOrJBvADkd4QWqf
zDgBCx4KecsJBShFKOH9jOm2CsyJkOwVflD1f4tJwRTPbOnZYMWdm6T7pezKucSLRE4qbZbmJtPL
Mon7HGk7utx4lvC02vCoKjXaQjuPLe98MfCtdjo4lNyNIp49w51pcEuA3EkxEyVWW9y1tttGczKR
EL7DvQQQZVFCSG9B0j6wNiJugkZ6h/3RFcbHgbpn222lE/3leQWoycCoRePQzjglb+TASPo+3BlJ
slwzXKvJyjv9RhhSqfKRddQY4+GgdjalxQhvJf8PfEQl3J8ikiMNzjqVmU+GIYrsq2xEl7Rkuh3l
/swpZFUcN9H6YXB2mVrW2If0OTaW5yrnUNBhJVgte08YaTPs+mb9LcVJnXcMLWHO+YfRQ/kcRl/v
XpE3xOVXuZB/PtiMr5dawQH8idACk+xOpbtI1de6YP2qzQXjD/0d+krxC/ODZRsPxOUQVIHrGm9V
PZAPWOPksAKkHAQpC/wy5OvQ78CyViEwRmiC5GpqwodU79FZH86W6ZI1xjGCysxRd3uoYN2g5o66
0TryzUUkJgO08/OyHtpCds9lYqzrHoJQk+/GJOTnJ6BlemjCY79V9BEO7P1EkDjomRQyCg4d8fXY
0YrE70G5XKqdQBRe+kZRIpD8A3FpIfcJuqeL7TlBLJMjIJxRzrIKN0c/qOvkLwRWMM4B4aBrL0kh
Kd+Gz+Tt02De+7TdwaAelcPK8jIz/OiMfAmz7gSHadQZgfVYNAR2Mj57o+3EXvC1haMgy7O23f9X
eE7WOElC//gZ0hmyKLV1RY7NWVe31Y0H9XdumOnJ8ZrDIsam6JypXOVgS+EQeviPQYhImC9HZpdU
9JP9ZkFjjilGpkzEFvKL7P5q6uIh83/mCD1DfqvFmPJE7BmUZgdMXrwpNfGx+flAFjpn394x36te
lLgh9KMtMTXjfSMlDD8Z1yg+msjP7jR5YPg5SifNILArQ35/z68hzClKg63GbRRxpU60EVl9OmjM
gR9fCfSli25zVU2ND4evWAgN8hQJHQb3ig6W+vdBjODENC8mOwJttSA2ByAA9KUjPRoTqE5RB224
ZjX3Uo6qSJVHPoabjnj6ax0aVH4uZsOqFbE01hKfARUAFKHVi/Xf9swxofccfaE/7q+v5nws1xjx
iEtUVcM6V+l/1YqehONURBaBHK0KOQ9P+B8Uy9VWYqbsqtSx6L5Ft3+fkd28E6NliO6O8VItpYmj
f23h6gzIR7s6TjrogGHbclOh3KkptnKBl4tQZ3BuC1EUTHcUU3IKC+8pGGeMd4hyLFDHSOEVvKDw
jz9k18QTum3TTAyq92x2cjY0+lbzcffxV9WFspvUsy9pHnw7wy+ghGcV+jVDvJ+kD8cDCjTKEbEZ
/gpU++bvptlxQmeKYbjrSnhl8LRdnTRLSKCLRBxqJGxRTN4GBjnJz6abW5iS9Fi2E1ohv/oZbzBe
5qg3FAyyaXoVj0EELgCUeQlk5g7tSzzPZoA8zpKfH6CKjFJ4QHU+O5EWhLYFx08Z9mJOqrNCsMQc
Odq5hGJAa3NX5CcoeNDwNi7ljKH9uSygh8vK6EbRrqFGZyW/DQU8SfYH7+idx+cuNbag21FQ8525
TixTil6vW1DX2tG783qNagzK7rMBfkKTB8MbXsCH19i7YGIgcl//jukcHZx+GBo1nAcP8VgCTgjp
qhg/K13vFVWfXxZzlZ9Nsf9kkqpdrOydw8YH6ulmyZ9sKBhdwmwBSgZXLZoOADvDTcUuzdwkz+VD
QKFRCp57CeIorNqkkDXRzHXLEkTkcpvygEmEVtOnPhB01ICkgAp9kLpisTiPlnE6vkedEEz+U6MO
jRNUcjS3qLJ+9cZeKvJIUQvfPhqTROt7FPWLpVM+IKhZ4BbF2hnyge06ZwOUAjJHpF1VhSonAPrx
6osy4DMstCDL+0YlaRnXay32ALHUVBKPmjSnco9PQOKxUzMrNShZUkIWRZTVpgRzS+ZeV5F7VQgG
u1fUYWIB29P47fc/hapxUcjV3W145Ql8/FdPNnX+/eoDBbSEEpYh9wy8v3Ej/OKX2PDQpuBlcAB3
KrQHRweuuUgmbWFo60LW+z5Daqw17R9HCv5ccHcTTQhdCJstIGeFVopQ97/dMi45bojEESE3mBNl
MQFIgzEjsJEbBxLsmoBK6TIOFJcwsLgWBBU+dCZf0niPS2lg5TAmyACj6yCmEqU1EtsLJEGIP5Uk
a2TscLCluOvEpkK2eKq/htKMf98mJ+sVlows3usCB6gHIT9b8y0ycQU+z6UJkkJqjqWB1WSe1AFA
L9LfZN1SDvBYwE5RJHKr/jpOcwVRwEDX0UYwtikWAEClGyxcY8nKdw1PFlnBM6g1+o02ADAW2O5o
Ndp1ghASWeLqS6M+DLxwInmg6r4EArt88ZKweXbl2CqxZ5Mr3nQCFiJhYiK4y44K8r8Gj95RZluq
PGyTGGzZsgticQXS963yMikb1PYyKWLy9H8SWDAv16LpHhVBAi0yHlYpjuq2AXMKZEfnJySipREs
bYURSgTG+l7TiYUAJ2nO4Q/sMzx9XbrpF0m2PLr9atiM5tfUo1Gvkg9vw4WYxlrJ6bfHpglmWVD4
WYjHQ2fzXyRC5BSQlYiljdm/EL3AWRbUpzWpt+VL2OUh6sf7VlNoGoPyyXLEWl08QlsgfVCHSJnS
L8Au/1mfFuuAHoOwm/mSkCqV4Zi/o7dwJqhZtDU8ZdokpkWHOH7OvzehPUdywjjJ1MMidst+t0Yo
EbNEYuxbsYUYIK0udzsIA99VPh5RFeCARq2kEx9gLwk+t7iKTJS9HU06i/M0YMMhFo43v97BdlVH
dIA4OUZpWYQkPGIvGFmso4SoUY61E5HcQChGd142BDYtCB1zRm/WwdvI2gNpt7zbVSP/Qhwz3AMv
CSz2aGkXQDHw1MThQieIzKWR120CEOjv+r5iWQDVhaC8zqT5q2ojaqfiV3TlNm6w5WPr7WuMIOEm
+ORREzxAr2lu6Vx8bzmUB+N9zgCH0f4QkyaELmCPx1qaNHm8CV2SIJ6dE2mYOIrOhsDGhJUxfnOw
7zckWnve559v0RNBAnQ/XRz/bF8u67p91XwqHViniaXwpOZm8QeQnF3jISg6GQK1CdKoVMW0av59
xRmfHafGiLNi6AU59T+fzPpn9dpalKsER6keTOK0/Nhn2+CSyC2nA2nqQqfTWWWVeb/4Q7en/2N9
FEwDbpQRt0PEPHvKStk4j6BKoRToZKGmeliA98wXO1dSljs7uaLML0EPbqxsTeKvq6zBNme8ipF8
CmPpyYk5jurdGjQqRWh7K1968HlyjA4FmX9aJciAcG1y7K7zSj0uGdDElW0hnBg+993S+pAiTIfo
XLmny2VdX+idA7z6vrUOamheqtTLFI/8cYMxdS8DLMgxL5g64eh5mToZliFazYjTlBGcFNiZkXbr
XDxMneZgFn0pQH6LuGLlFiTOwn4N6zGI9wXq+gmkhCAmITCnTNDoexnvsGyPUrUO0H96s06o/DUr
J6QvlYh1G+Sq6Ej8MFaRjJLg0V7mROvZzwgLP6JAHZgF4/Vbo7ugS5Izb0k8z+8utS4RYOlLAVLx
32Pm4o/3+ApGTXqGIW3bMir2PoP4z7cyvUw0SMefMoeIZYkRsIZqE777g4UC/RsWhc6l7DVHvJQn
vbFLJwXTsAKlf/kWUbA03kXTLXwDgP8YFIEifIydDH7Bw9PoL3YksJ0CyvVYeovDgx82Z6BtJ9CB
HZs2lIE1LjZSZY+/UjDiQRxbYbQeObTd7BSXB6cTYcSAY/gZIAyMLhGVvfHg2TAjUlhg7gnYngEZ
hajfsoVzztPAMLAeIWLEACgNSx13jIRKg7lEZCiA//1h6XpbLjNF9AkZXh5yGQ92Pd8RV5DTGfVr
VZqU36dBEiacdZFg3dFYNX0W6ubNbfJvIbBWn/Sqiqsy2PPZqyfSAsw39uKA3D1lESAID1AQSY0/
bj9LfcjCHYU+zl9K+o+MJVWkCWzPvEUlXGC4nf5R2hNke/rkQEOteA9P0SlRAQ7QEnxJelNpgm+/
IDU3pKvafEDu3Ey00cljCuH8loN1T1tuwumaVNEFvOptzZ8t4wrovdwhj7jdwFuNUf7vCnpDNFau
IOY6ZGEsmh1N5MbHm5sZWMO0pT3hmLb1ChUsiCkQL/LHMPth5iwPgqcxPVVR0VzBMnwlvCFeAYuR
aR+8fZh+5NUOF2vhcJXE+oiLZ9GbkCk5K7NaotTIkSmEOygBn3sPODqjQXnD5bb66any892lxj4/
Y3gzdYBydYP0Zi56rLyVcTsIgTy8SpgU8QnYilf1twEacJ0lavOcIxlv27E7wuqluBcoYahd1ddq
dSQ9cZJDA3DJ+wtAoqCjWVpr6SWccVRbHD4XIdsencmVSJkT4kQIb9JaeCXdr8kCx3dRO39ADmTm
j2s7OO6ovVfibuzTXAs+KAGTDEaRtCtIngrfeI12aEATrB8hC9TW8Cvwjiv8LvRmBwXzbTw5eFd2
UVmuro/gzUje5AYHLH73TprYdnkl55nip1+D/NWJeZrtY0JAbuqQ3C8cCNB8ifd8Z6xNrssnDCZk
X0i+Xhr6tgGJRoEVGfc1WAbw/Nc4r3g53IBKpYZqIx3Jae/t6boBS/ekMoFpzarnzaapfQN1ojtJ
vyWlkF5600oRPWTH7GoFR8ES8mR07nxSnvKD9ECNyWmbNAKXRs1pVXBMffMLVrnMkV4yWrK52Fri
03JuAT/DBwRNAiYI6emg+xW8wwtnoA7lWu6kyDyZ+ky66cNPDQV/NizQBALtsUmTn/IN7S+2JrOL
XNG5R42/PWpDkymCmX8SNefATPdohjOoErCI04Ejij/0ovPuDyhyATHakd5Z3lNVSOhzH5eqU/yE
2mt/8G4mKApYCQq6FywfDru6UqiIsc0yS2ANPaeUcvlhMFiRNsp+AiZaiLqDrMaNwMmFySJpmiom
rBBvOkYZJlNBzoC3kYz5kUY2YugHQpDMrqpzjDrLvgIld/I+9BDIVsWHBJHMLK/Dr+mN5C0KDor/
3LXw3FJqG+yM2Y6DoK6oCZC9D9RK3NHzJgmJsRYePfcOVUos6DBLdjl2USHpV5jQRgdnaxcYZMLd
olU3Gl2xKZWaCKVMO9ddfCwRjPwMmo9UZ67ttb5+WH+nSaFPf3Pi1ynykdtxVfhcmIQ0gf3JsKEq
r/CFWpN1GrfqWbLSbe/le2Hst42y9jnP2PGr01rNV7gUugJkgBiDzEas3iVD8HDi4IKFI9F9Gi9e
GhzGzUvvqTs6/vmDJ+SJURowPx7VGUBTEu4vQA/VBvHQvcapJyt8fGACW5vEwZqNMvhOzr1N/m9Q
eX70knSbl5bn1sru4DoOYKx1fjXaSQEl0xvA5dFnQmf5yCoWE9ru7wWwy01YU5FV9UV/LUz8RSR1
KMJyLSVg5ABbQcmjcEyb3o1s6yRcNKgZ6OAGHJIingvlgdnwMyLTfhfxDYgSDwM3mPYcgVrtE5qY
36IGKLzgL8UPpkVWJmPccMnm4U2G4UR2Wgxn7hpXnKpZf1UqN59UDUxPDp424E40D8Jwya5X8bIw
iZzWckdEg2evFeXdhSKQ0EGGPewSfXQRbe6PfFzyKrBYlAWuv6MRwxoEkgUDex0wgxaOZFd9Qp8B
48RhsVpD/UwWqwZAN9CSdkIM3EJlZ8dNTt50uEfOYe7gK/JSDp1wZoKtsAxajYRqGmXRv2FrGg4E
Sc1gkH1deVlJFzDLplvwP0hsRssNvYA+df8ijsQANP0jlAM0GUndez1RnDB+J/miKE0DxrtzfCWV
KNv8phkkdvS7jmufGbr+PZbtmowCp2c06Zwfx/SkQdIg5j0pc3CIWO7uUT52HV+YKSP+l0nvrcdZ
q8a53oCq2wJu0uC3e+EJ9EA9g0d4M1L5YjvvTjRFA69VEC74lEQBuwhgqRK1oBfA2Us1BA3Ikqsl
iQcEV88gwYNWjyT/ym/rjhZFheFXxFN74JYJLdbnc8d0m5wA1vxNQPXhlGal3MBSKx+LWMFdSdqC
KR+5CcEWMgQe4MiyeUZhb9BLj6f5c2M82yut0IBM5X53pxFqXoGtGNfubdhxLHVf74ibUDe9Kk+0
w0ma5bWmiHPVuA3Gjvy3/uklZIU5/2K3hU+rViijEaJ3obKksBYMOP2l6sCCix8+6GvGNVGf9B+y
VWINPky1Wji8sEXSTxosdgHsECA193y2wVGgqw4JhUD44JrWNnQAH/MF1vrTGEaAyDjw2j0Nf5x9
Akb9sV93hE0T8vyKqHNDpSjdXs/TUfXBGbwLfl/IP4VzOlpNDm4afVv/SbJzgCqT5c93fO1zn612
i6oI+kXSG+FbPsB1xvLCpCidnTFze7GyqSvwZQ8vrfgI2/dueMgS272Sw6pYmyRQ9VeFJxdC4PPv
0b4tdrfB44hktVInqSKecKrAJdbXVjYDEBNAN5G+Q1Hk69BVfMtfWnuaaDflb9f64GY8cYDzUfzK
LnYG60vOmmE2wV62zIhXQEjeh4k/VPc7ZBIDGhx0Tstdn8L6p9fvKF03yvKa+/jhpTefGO/Jr5oW
0utIvm+KWCgg4GitZsQZK+wgZXe7htcQxo7uPtia8HK914tJJqb+Mt2CVhTDlh5H3jvcrqM4hqCs
BhLk3oWY/QXgOEmz4RxciWXq6HLR3ryUjK/Rdf8x070DMuc3e8OpDZ41bl403Bf48Gh7jFLR5/SR
DDeEybKkx98ItFht2SJkcPrxr3Z/V96I7Tl20x/4bxNdXckb58cC5EMWIjHy8DKDutlosHQE8AQ9
ntwJTlx1xYH82H7dg4hAGrDFqcZtnaz/drF5eshbOPsYWde1NDKLOi7EQb0d/5FlqiWXsCSnaNoY
SRu05u6iu7O3jD19GT2ikCwz7x9JRU05I8mk0wIVPAfQgmYPXKrbC/Ig33DSlwCfOaI44h8HN0zS
2ps4Wx1PIVjXzypsVrImgCFeCq6YdpdjXNZH4Wh20MrLdLZtNHUN5z0hX0qFK0xJFsyM6Apwxyl6
Nt1Y3jrqikDk6VK9U+mPIvH31DJQ9qa7liQaxAPqZ8n73Ih3vyHn6Z/5PNU6aD+MeaciVW2HlrsY
azK8fZT5rVo0/H8GiHgj1JjHn6VSPWeDmSP+4bL1wJmIh328RcCWubo4/RzzlrJaMYqYncJmaUpU
wQmI9rIf8xpiOzJVXjt9yBv3F67zQ/rvlkSaeWJQZnXbgf5qhp5EAjMllDHGOcFstObWkweUkdth
Lj0EAgW5uapPjhU6ifzEbVjYQa4qf3OVOrmn1coDuwXO0tSLMUKg6PfDDWeuMKgDquBYnzWnSfTs
Tbu9o3idstFS7YcSF555UoUu9GM9VrhqvtOglvzXehQPOXiEWHlIz3UeAPzmBg5pIUIgeHtLIoLr
KJtHLkzhrRmXy6qhIHYswifPDm9KUmt6Cd0uWmLX95CL+whFOd0ViOIDMLpZ+6TmwVTj784aXudy
ndGDi9cfsknu+Sildhq6i647Di3X7DdDTxveuiJDPydFNtzIhtfNSw528KMcpc9ddo8XSS8ZLuqj
AubnWzpQzvY0Ozxtn50JHq9xtK2JM5QV2juZnlahRB7cCxJoCxUxVAtDWWrfZ/CrGSEs1bz4obfg
ERWzuYC4AxppQkH0G98CP3Q9nMgBO9TMrt2a5mZPt0RKC5WodIWNPcD9SkM99N6iLdiBGoITc53i
TLvf/vg7HZvrztaThH7gyFurHlm2CBZWQdgvgynez/cDrM3SFl6CnzLykg9/FvAWjFbuZSlUIXoJ
Urzn4eBhsWPhQjoABqPasEF7D6NwevmZivMtG0P3pvrvpTRq+d4B9oh7YRIfat2z/4vKZFkT5qV9
fOzxIMoYVJBySAmiSERzkmbnWSZ9gD1Ef6+KaCEb+OR/GerPVfYVAZ6WGN5pgsNLCf3woBDGiGSz
KQS5kfcB0nNcelkBiU6V4xT4puiEHMNacAzbCNnEZQQfd3bkthMRVpRwLf537vqIp9zt2pMbVHHK
kGZoPKjK76LPJdsfMVbNG9TrkVXqvc9dUONSuZl6CSeazj/aL92pUgP5nuREtg1lqY7WUF62c8gp
m3W5u9739d3vNQVuIJsJq5JS3URF8LzHTjgGcQBkvFHl7JOFJzWLdm+9JuBguqAtFGMFkeSn7wBs
ltk1vrypiIzwmevYWnkMQdNMbiUTZ898Pj2afLG0lEF9NzxIe29sHrzH7cD6cgytsHmbRlKwhe/E
vtJQVs7It+edMpBHZ4Dwf4e+u8odDyVqyCGTOoCSNyjO7OrHrAsE1kCVb4y6sR+pj7r+pXaVNywI
VjQpjaq4xN8wBjgvKp5K3O11CJfOrNIhLQmTtNkT+SU+9Xa7BUZgLMKdDlfmvEsbXQg0OKiwRW+e
4wFcoMPw1dAUOzAc0aXFsY5sx3EuumORV3N3E4Sc5Ji/EC20Pi6tdrusyMHaoPowRPU2A6k+NqRQ
HGJUbFAh+tQ7/dnzFzhBbZZOR4IUNSv5ebbfWuOOzDakqtEKb6SuVCxWYZFzdAhsjUqUQZyKag57
dm3sPJrp1OFi0kYg5vi4h5sKZqVkSyumDR9dgdn5KUXS5wgY6Q52gubJpwBuf0cvQwsTCJ3As6Ol
FGibHUvdgoojB9xX3t9aimtkcewJGycKl1re31gVlixRZ4vP68yEhoMmaYbOd2UDcITrfq5b3QkR
SuAh3QJfHstj885V8mLlAC7O5A1trFMaEC1/rq891uljXeVhrfX1RZJKTN7Wb0ixDk7+vsSLc1Dm
MQOz8mE9XNVOv1Oqhb/7RcLh/gQANMFoZbWeNZuhqXZs3ZcelKbM0MUHw20YMseE9wTvd2kOqHf0
kBFe62BV6BYdBE7fMAOASK9rQRg6ZC/XrkZN9SqP94kApUZK9ajtYO3vfDczYvI2begu3cD5Y/0y
pb6C8KaYhkMwPSdRCD2tUdXAfpVhOVs+ltBZxTz1hyudXqlTK6hnctHzaQEQUmxaK1tsxWMRFq1g
3/yzGTc8TxLIu3REm5nk7FkKfJCa2lMESV2Zjup+g6so6kibn4gHxrYUoWJwHu5DzpeDgr8l2k/E
Q1bYlF7XJTqsal+N6zq3KPNSmoiMsy/BeaXqNeIpBrFVPW7Z1HNb+Kqi5/+GF4bv9tWtfa0JgZGP
J5qDoKRmJxzPq1PgBuxcfJfugmRpumEaYwZfosn7h7Z7tHcxaMGE2geIUsE/bE4mUCH9Im5pV1jE
RINbDMwOOagt7MFQXIHWa6oJ8VdmqdsfoshP8oiuhHwYt2KH48EFbur6nIjU3IKGPb8u6YAvnJAy
KEMyEx+gPPJkYy3HfSXavzRk5mUrxbXXx70Qwn7twGAypHpIiywm6OqFDr4ulm52Xx9RPdgdq9rH
w5Aldm3R4Wc1+H8PnTsIDGZsHv5VYAKLoNRFGT5M9Mu7ozdrOaqYvRvef2JNpGvjltGcY60OIOJK
P0so9EHGfEFPUTF3xys899pWjKywJdYx1YyfNc4bBsBIjfLkstRBnFEjV5Ivm042Uf0+CMx9+HaK
xxiJQeTL28EYLiByl9g8TowpnJ4z20SSOBj+xl5OImxTzOnVeh6P+ABYKIap0sgdE8jmTWfpcz3D
dtaBMr56BRPuv07O+EiF1Lf0g4SD2bXvqlHRx7ilOQe3IcMGvR69oTQdrW1OI9PBPeEq1YmsY0an
lLlROMcTAwzwLP9aTB0Cf+w53ROP5fKHUAXdnGDTb+3Om+uW2T0IxnjQuO+sFhVuEx6ERQIThmLG
ObzIzRtorfgMDT84clL+kyhy+NjoPnraduP0IbWbRv8vnwzKMeY6xrbRJ6hKLLHYWhQYsWh5ak6v
JafbeRHVSbdWacI2QIlx3N2bWbcBPataQDvxaaYytM2gMP13k9BKF5196bGT7NpjjYzZTjeJtjwB
6eC9qCy9MBnMtrHFQzI9PZfQ1NHZtNXBcUXliHCChSQFmsUumkUN99eV+SxHjJEpe9Y7xZUiea2g
zpDv2IdaDEMKer2ngSJql2C163VDdfyatY41tFlKyc2dlyWRk4BigFEvuRZTY2C+Cfp4OcpmtEXS
S6xl9gvc29gwGZuF+iI2mv6kgTjlkrrgWIEuZf8u9mHqG799fbwI8XfZ0jpPRhwqK23WjNEDtPoD
2o5FCMa7A4G2bD8JrsOCLy3Kz31Ppso0O2K/x6mdo9nT0g4SC/Sbk1c1D4PFRtQ1N3GwEDiSHKOo
JIohwKFtZ0cV+dcWs5M7BpUxsO+qUWwaq3n6JO3chZ2pY5I2MuipM+f7SvfGaGMxNz0a6OjDnF8Z
PaiTq/W1D4RCMvAn/O9YXQm0VeDWiPYeFqrPXwzvSSUKAZPZ+j26Yww14sVqWVa0URZKRNlkICV9
szLCMoajytAO6uwF4PPq+45FcywcvWJCKnBxyUGhys8+pdqDFbsOdXc8qIu+OpY3OrTCg1LtcEAx
9TrIg4rh/1Cn1VKec9you+VrAvGX/+Rhzx3XWOl40ppuQiSfsKqu9k8n00HmoOQXAkpKllvRHJpn
pdksV/XkoWzhdHHALUuj4BZHPzYLc+ON8ZrL5YsQYBeG8W+/sTFPrz04IloOx9nmgXu70Q2XZYJM
vR784Pt5A3bEYiYfnz9a2FnPThEVrvcP2wQFQjsuPFP4umMboZdQnxuwTc8cFz1T9WFBVUswJiab
H7jA971NoVK8AHFCtpI3JhXYpCCQOXn79IojPSFE55hrxLHgJqFAJlr6+dXPvW2MlnjoEN3ILo04
Sv4/6l/4CJfdF4S6M+Jz6DLuyE7Y83cXOc1IN6+ktYK8LgZyMNuH/VZh37RbCBTCR6PKXQth8Q48
g33tTxLGnTLWKIIiab2Sdng4jyEXI+sm9Ofpo1PEohLBg0uRA6eGtX5Iz77c2aF9Lt5b5amR6rlO
fSkcCkEjMuKxo85gyH0V0c3UuqwutciVfM35qofKdm79OWn8WKjqRWABgbUekIzp3BnL9aj9CJwx
1I2c4NaOqczRUGW+NHDz1xjk42p1oEzH2hhZCPuXJW59bBnvBXIqfiGLeBuG4U4wFYRZOFciTB+W
uy+ZIKrQhYA3nblhVwnNkmjOXARhK58k3r0uZ4H/Ufb7OViTevNG4pqst37Ysrhp4m1uTgMRjJgM
5AUEHiY2qKrPXgbWlhatxIX3rommHbhRK/RfsEq8nAmFxpuHLdMVd1rD7DoOYFYcGtGPadUj/Eti
ZY8YcyxWf9sLmXPJVF1Fo4wYcx+JkN1IgPSWCnTlkKzszfJGtsAwsMt6XESxDTUbP1kjzFoiZowS
lfo7npbSSyg155X0oxbF8PTWz87iZ0TpTXXg4Q/dE1e9cZFgV2p8DBFKVwGn+T8Xkb0Hk51Rg8no
RSHZBN+29KKv+Q0gi48/ux7+OJFg+i1dPyOyBAYFGBfvyGxb3MDRT9fT/f6JHAEJ2UonmDRgNtEU
HVecA6Px1S9+n11K9uAykRCSsGibNqeOe4YpVpoZLdo4FHu7tItfQOQClEbhYcXP6OKuQxWPLZz8
aTkycZ9CYtovMpcfd3ZR21pPoU47+0EAHx8L6ZMSnAfUQGN0wAPQVT+edsPABFpNC34WSvMKF7ik
rtRAlCPM7tgI1TO+yypnKx3IArhAWxoLI9IG0al+PXz+WY+pEzKwVk4tDlHHaygDWk6QAZJ6yeE9
tdiMsEl7DQvyW26n79FP2KYB+m5SGgt6UGadw9mMXog5dMOQApY7VbaAgbIOmr05nwCx0aX225Ts
owU+nBqPztsQXLBuOr1JYTv4rPRL8hS7bIMVAduAUmy6PNllcG9rLfaJjEx/Y9BcgcKz25yZneNg
HiLZ/N45B/rqss9yMtnOthCyy7fTUM0mMNmSMrjTbfAmWNXxeKvk3rgAxB6sOO/aa3CrQTvNxbAv
251WxvCQeusknyBMHAUZVRshVoYHTEPXY59ToQEUTZ2Rl01G2ARtwnENAGmYU01ALrwapdN/KMRI
ThusN9KZqd1+hzKl0FoI+lmKzyTVErdU1qxx9VLc6Cnv/Yb1jmPGTxfpN3x8HhiSdt+CNgOneYBn
FpYiaSv28hcGvCJazHblNo2zdnhWmdQxCcbuAHEh5UuWIkavqHWfsYPl7BF9AOxyG8sPvit5y9U/
wVXRoK0GVQbVof/aPhFHgXcaCHDHbj/7xebC+gUmDUDGW3QOS3+dBy9os/8/t99/lgK+TI+uImHl
GTaBEY3V2NWOUe4cCFJSqaUU8fCFQr3hkQ9tmbZB/wv49QZ+wtm0eWi7u7ioki7PP0TUicXs0MAs
r9F5fXes+7VRvYnsDW0EivyGYRqg7fH1Jj8DyJ2fafFpl6baA0Z/F/6NsJBgPJy3DqJ4pIvIB5Pw
nSstcwu3BADBjwErFpiTkMV4Zgt0y/e+TyYQs2cBRFzk2IWcNNHilQIeKqYBlzhaDh3qa+giLWEP
8e+ace8K7888uAhYKWP6TzqFxCZWAFtybJMMM+ESNeVEV+RqrCVixOIsI6M1nw2DC4FNq+zcKOsD
hBXQjKxKTPxDywFkEri4LppP4hyyQm5wKpwKriHZY05i/hhIit4JHqO1R+MtV0ZJMM2AmUfgIReY
f+arhNIJO0igkBoGur5Y1wNGHntXk9MCdNs1tey9LKy29ZyiNGnLfwnEF3p+Z31BBjXhQ3SzSFzo
Lcfe2fcp9P4vm4grYLLzgqG2qTb6GLz91JyURFrU5rlpMc6XavVgvVpITyhBWFSqAWrxPztpz9t3
Vf4f44/4J9BAsMW+rR6/4S0Isz/2CqhAL8EIrr2dt+aJtFzVUlmJDYZxYB8CoBV+k6zFpPZBiJgd
G54iN2/94L3B9J/nCIOc9x8WjJUIVSdR1bTiT+e0qb276p0jJ8SUDxMKDQvV/b/qVQIScQSnzy90
y42pxZ29fMYhp7n92ZfJSQuko05hrundFU8WTkrnuzZwNr7jTa8QEfkDl56TLbiMgyz/Cn6z+owG
vPSkmBKgNTkPhjD9eiFelF07JN1GHLOBOJ1hDFWzInE98tU/3w7aeBQTYH93kvDR/w/nS9QyVSpx
/0qZKT+6RqKPWyD5DioJB4cH4xgK+MYQbRFP/dd/2oorutzIOg8qTDAU/AyDiS2yFzJdccNoQlTl
UU1kY9P5kDTDKAPuswYN7cFzDWvcdB+RWtNOvghgvfYhrOZkT3Bc9JHAXj8xdWeRSn0Yqa1D0hja
RffntGSz5dxKCeDIXt2wZRbl48h+ndIFISFddae9xw/I6apavjQYKOQqqLWbeOlEzP6jwy6kZoUL
OmTI3q7OHzIpge57oaSpFnJ480FMk9SXBPmlRs1FA745oeA7qEudmxq2Rz1iSOVzYnjtycQHd3tZ
ebTNNr4CcAk8cuzodbcaS4TbeuhjDhYUGipumIGYTuReZ76fi9vjQDa7nozrcFinF/Pp3MU3qs0M
Yrn9pctpYXitLjLzaIb3kuT3HZ+/85hm4wMAbL9NZYghrcGzzrCLkWR41sykUerSJxyWvqp9T4g7
MT0pMrJsYg0NA0Z7T2fVk6PhiVYcv4CAMv0LEW7/qV2GchvhsPI4P9TBEyr4VrING8H14Qc4UplR
PgFeqKz+hX45jABtVmLlWkRU0vCTz4kLv9yDmRDvFks37eIvvduOYzDs1JSGiItR3M4gG7tLrNjp
tgv5HWF7lnElX7Qd+a1qvZ1JnExgFnjTls2thx3tYLnHTpfsRg73ccqcQio+itXEnSwxUJNYQxzU
PwVOsMBAt1XrS7/Nkh4Hn3sl5KhII88R2b2Joo++7UU5jUeyiZZHoFquj9KUuCIGiwRkpH7EPycu
5kvw82mdE2WlCoC3s5A6Q+XSj7++RblaWSKHSeuQ1TmaWwdACrN9DuGHTppb5628MtYUsNjEbw3x
b4sqszk+fmAZqRbQFKiDZDIsBNvG/lwRME1d0qQnR6TWmTH37Cpk0EFMPkKJmbSChvFTEFJT8eBN
YTlefLg7XxnavzOB9utIz27Z/xiRAL6zitAcopZSVxJYkdyLHHGRQmY44xtM3sIiiztfz635X0nU
FwQuSbXYTKkfTEcXAaor6GEJOMiZbK+pCwOtTN/h7OL48g4E7O66FabJW2NAN525iuM13Oa6Vu9Y
YKXXZy6E40bK2rLmISOVYwYHLGvlgU9tVxskqS0VnNcfLOxThi7WkV3nt6GU/PqglmNnhStrB4qY
Tx4DRmSKqW2uB6n7nyjtE+TBf+F4Xk6O7wkI2fLL0PQWTTOf6NrjunsEOC0wtTfMWxmcv9geMuBM
LXoJqco07HVH9HTbmVYYGTjYQgGrMWyc0og4wvj9VjKsQ7kypfCgxLcI/a3xuV3JVU+ZgxIx0vkP
YrfLPwufQIbZ/rXoOFqh8zGpjvah6G7rKf12NOGGUFTV5jbhBDF+NCj0YsfNfsBry0VUGuh2DoCY
eTkWHhI7cRocEo4CgvxPaF4wNNY102i/Jiij1f7QGKd6wZ4/N1ZjMN1eU089VNVrQchi4ijgRDXs
5cNVLa0UAsxdDXHVaUqmTeymPGZCYocpdVt0liFJ0h9eDBGmT3b4wXcJ3bCLWIbwTWnYfhouXDV4
m57kv3nIJjzy+EwLgf9JSPMyWyjBUoWIrt348NnnCcAWE8AxZgS2vfzLKz5S0VmX89I+6yHYP0wH
IBwIQFMmkRtwQDhscEh1Ixip4mGOnM271Q4foKEIFjTp9u7fd6ruOjodbogMtgikgtr6OQX3wK8E
YVx1JDW4pw7lZa5+6NDW1J0XsKSdpLfdsAPRKie46Z1qDFiJ4Yj7ztF5C1Cnzlwx49vA+2qY7qje
sGgngKjcqtUQoF9+uVK5kadgQs3JVKjcXr/OkDFv+0TfsOkfONbawqc4LhplFFeLk4Wf4L5+79ks
daLAjTsyRdebl+BoXS7ik7bQIaUUbFoqvOuF1iBKguMzHMw1AJ+wdeROb9RrrC3GlshHLqR1OE/1
suZKxBs001hPSx4SYMZ1oE8vmKTBBt2NcO7+bON61m7i+H7JuTdXCodM30WClQUCzFA0beEFmddV
LJYkPqUijOqHHXKuNg0F/8L5aE9davFPrkiKSMFcqP2Xw5YOuUfKBHOC+fsiHavHKoLa7EMutZQm
thAE6H/Jo/GQoFh/vpIR7YsvBku3F5EmOkLKoetJsLS0wCRK3u9sXlSbVuzN5ZEX2HIGNZaY5Cp2
SjWI0uCP4Z9VJToz3V/EpVFgiomkTrPAIKZ6svxcCMB+IsAmQp8rooNZTSZAdYMgtXgo4Z4Ks3Rw
h3ES7Iopd5HMHoARbi6tyJGHVnRAdjlFI5bPuOXRwPHZFifUGW6YvIT/+GHQjJnysw8g7fY2vDgd
Jnb5MeOY/UMBek9IbgwqnVsibIXUas5tX1vTFhus6x+iUyZX+IMAdolu2dY9D4UV5+xY5rAmz18I
OWxiHJvxrib8A//IkXfolHZ5kckas7H97qpI3vKC7luLKYu9eR9kPSIXEkN7oVhSjVm1UrOKMcuD
TYLaz6pJfuI9I44PIYy3b+Ie5WHyJfwhI/MbBEGDgP9BHO1QmsuwO+UIj2xxGCYugCW3fm0GOkEU
fBEnrAHj+wz3pZkYPf2QrmAL6vgGeNgAX5dbWyNZ6qQ6RpKMn9FQ352MiAdw7g09IlYs8kETaNtc
X4mOm1sxXNi84XHSZ6lvArat87uhRiAbbnM+VKivfBYUJNp3HlDu7ef59CYyV974BAkdDYNEHU67
Ce+OSVPGWdcvzdESN+eyLpEV5NWmqShrEh1O7te8uVufVE2xbpYy5DcdM3O1AyBT/J/SS4X414EJ
uzw5Gx4H3RLYzM29qfoUnmEZ66mUd2bBYMwwps0DLmH9F20HX8xiIbtKJT/ckRmdCh/R25Q8bG17
dCQMcRSl6/PE8LuFj0emCxjlJedJwroboeFJBPMcigDzqgZoNeL2adw6TaqrypQPZaeRUhtYb92I
TM4mge0WY9oDtUHqFjK6dfWOK55c+x4umYE4ou3f5AyJqToL3HjEGp2RQHyAvbcwfy264bdfm51j
k0Dxy6Jnk5pHSUQufXZA1hQngTKGWplZyWtnwuX1ho4EOjI9lL151nl8ROPen4lT2DOVdrxk0RCt
S3m8BQRWFRGn02KJ1kFqXSZVGBnIB0H1sTE8tDm4m7+pasuUginMcB6KZpMEoTeK70yRUgucHCoC
/5Vc5BukB0vj0RDHjypOFbz/m1Vx2H1sKFA+oOd8inhg2BCdwfq+iRkOmQDNI1USMUbgyTZakLgm
VHOW5EBliNdmB/3snPnFgaEq5INQhRnFmmTjENPXDqy08cdrI1nCsr30th/75+VQQcLeErN/PQ/v
RejaprQNLSULW9gBIf3cYWOmMp2hRF/Y4TfTxO6SoGIwmYpikgh23csxzKJbE9xw5I8VafSXty8b
juNmeE3jmUXq7HQwlG2Vf74+HKoWk3XJvFM5Q8u/BSYsjDq8fwuhn4qZiprF3fpJoz38SPczMDJh
YYLFutMcLaVPq46zrQzca0SsCd744GIw4DQjpeeZGuL942ck6geY5y6IfjQCN4U/mtyAf4C7lDHx
pw2NEZ3VD1LXbXjCUoZ+3CgZJUSFrhSVAVOMcWMUpYLvTy+YWPWZiCFOQ6/zXKKSWBY/nUQl2Qv+
cMMQeUczhLjSV/ujEpeA0elm7W9fW9856W7YZDRGGBDyT8RcIo12+iQcp63pxfOcqfu6OpjbjLQJ
gcZ8opVD7TotMCsjdUkn9pPF0CdUnCWUrNZbINKg0otleW1aN7Gw+i50A6ZqipkSBRZYQ7EVbD/u
NfvW8XLPySXKDjkPiSc3oaALoJF1vGvbgOJDTGsmOSTi+DXf8L7h1VkYRzMs2HI+p4eKoXP3TByA
qtiEwm/AO3UqMx+6ab17REgBHJgAq+dc+ILUZc8Qa837iPBhgYMFhZj+BFWlFOdAfNSsDlTvOvHH
s7pHQ2FQd6ki9CHtW0Qft7k0isUCMrt/XB6PsPriZuqc+YjiPtnsyqLKMmS3Qieyc0JzZs1LQ12p
LC6Z3Q8LTFQ1tOgrWtA8mC6+E5KEzPDGFbvNI512tiJU0A7QkctNlY9sIcMb1b8Dr5IJPckkQbsx
WPE3N1KeDZ3O+7ShicLXh4C5DHI1l7h9ai0Zjote6GBPJ4hIEaOtYS1l+Z2ZQcdrY4ijINKuo1lw
iuvfY/5HpbIXTHvoxs3cn9kd8o9wvMLEShcyFsUii0QVxb6xDTBTfxWXDXd533Svy/LEpkuJhTE5
Kk0lELoBAVXg7yCtFYM0BBqLQOTkb+F4L23W81FFPmpY41XBmd7V0120FNW3oNrnM+dX7pGOMPWi
uB9URjhL61S75cgRCVHDNRJip5SqhEOJmLnKKj1l2Nt7oeBVMRzPN2r4xK1idzc8AM3k2P/JNYIE
QvagflpQOYC0y21meCPRb4F3X4pJs25s2l5FfJB/1R6GXy7I6PSovrqmL9svzBQI6Jx10y1ysZOS
msLJN/C8sxCVL44gfTH+L+ZD2Nx+WNsPNJ1ojTRNf3W5yCWoodULh/gkTaaJEziErCqCqIsXTtRL
hm1l8RP+6DhlodX+FHA4bvV5dP6yp3Mit/5BhGy6y7nXHPmkTAdTiyeuLAKyaxCJe8AhlAstvV39
Xj0ZNEjXG5sePv7KFmmJUp5YsZ6ieVJkyhEB6CLk8h+QY190AzYN8u5wPwr9a3jHkJrOAGlbejI0
qMcLdaL06fgcEz9r2qxBS8XoDBBLGNCokgsEHaNpghddQaVcxMuT7698wL+KoYoSkrDHeIXnWr65
rKKpIuGs/ttwlrUQp5+KDqUxrQiLa5vxFUKCwOquBXtLxyTHTvp/XRXS0Zfs41H+TzFpi0WA4buV
qV0yYeAamTvlTCxWi5XpWmbvs8FSnZIXSqWYVG3UqmJYRqLXntCh07yW4o/E6G1NqmdbCOj21/Wo
1oRiNk7Vrf5ZUhwPRPGGz/zp9zCHw1bvuKEKq/SurG6sTmeN7RC4WFsEWxMJiez8uzwfke4ho0xz
wrfqz8h67Pvoh3VysYBJC8AtHtb5aocOY9yAH2UuTMrKSxVILC/H34IR8ZIndNLmuxn9rPplqxqk
uMfQfyPZN6J59QV5UtpFqSaijtLlrJhyweHwNTpudTeLqpyJ+a7ydPfz3MI8zx8VcwYYWZXfU25f
KSyh6uWgVbjZfI9i4ZP2ECBo/n4MNdJdl08hPoRy9+msux0OMZ8FKD/3x7Yi/DZKzX0FBGgJpJKT
c8o0MtQ7COG6mvddT4ZKaRKmV6b0EfJ4JU5cAqVwQtqW2xnkyKwyK+tgiQZCMRg0JlA43/i5ol2C
ZQbkQd65CPLQ7eKi4nRmNezIhFrfzXHpDWsnun3xLxWpEbrf6DKBKvbbq4XfQhLq2r+z0Mvvm3pK
sWM0v+TUE6HW3nJv8j6TXZF8pLXzGFigjczuwMmIuUZGZ5iYrTZze2rjOp1xjV/V/pB9l+BO2bkK
YifpGVr3A4dPHBvPh4+NpDfa7f9zhT5I3OvFE9NHO43P52ZrphW7/JeZeAMPy54XI+DD79goHT1x
YwhwIffsJ0u2nyEj2TBF405txVf3zQF8OSflsFQnTxnjz8rhkF5iCYKLyrM0cS+LD+JO6Xl06xoQ
rCY0c4ptMKPdc8LJ1DqOB8WkdWpGxvzVedBqUA1OdqguZAbM6Q9bZQJsb9XfO+cIKXOJoBCexS8F
17TjpPMH5wNVpnEeoL9QqwaUiK8IH8NDGf60TiKa1pr7rMleMIGjx6F86fm4HdMePnseG+QIQk1l
u6noNINl3ItAcFoHrdaOKRQYTLIR8RB29bJKsjyNChSLwhUk7XKZyj99bcH6fcztuKcAsTJvX4jI
yoQc5dlCaxAkNe8W6f1wjfwulqNsggh6fyUSGgHFf7kjKG0C8R0pdb0Qoj1RiAiAO1hnXXQkikQE
vbwtZ6ijHdRvA6Rcs2K2N2PvBayOdMt6sZkW+iZhZxLJ+XO3IkZSocTAeD4WMw4VGlSsHD+Ccvzk
zxa8NzgZ7IjT0Srng153lyb01Mq4tLzIBk9OQ/J2hC9M6H0p+hIArF5yNfOgi0R8lUcmIwTH0b8u
f8VLky95wGR4z9V8/FsBDcGtgQNWfAO7ueCFG3CavZ8E1FstAHQM1QG0nVMhWMPqfQQ0rmdN3u2t
iv8Pf2HJVqyOCVRFre/d+RBi8jDvrXcYbk1mYOPh9SYcG2FYy5sXzBO5H8rgDn1n83JWDofSluOi
U31ydiEvXka440gNSir0+R3Phs11enToG1e89VwswSHCkxmEzyN8NH/TU6Jqsx5S6UA86ypyH8KJ
12pTwKYmvgsBejECzkdu3Tz+p9tDvNQAzCGKOzzZfyglQ7sua3IE40i//km1PfXc62dino9JWYhT
mICmL6xMKlNhy3dIR4jAV3bYxYyyIUrlZMiE+dIpuaL/uRjbicgDMQJA0LBxV3tLY8IlGdxD/+J8
hndAmQcUCuBS/AU4ThNOs+SLoAgNBmgRvdx4OU1jwhJavrE+kIXHFc1Ongdh/FDJC0Ewp2V3uMAh
L/k18jEYchSEEIMUVmw6LyjLDd4JsXI8pVeEBRWHYo+gKeCoYNFYL8hSrcCNjyudcboc8unYU/66
pwjlO1PEVubtTmqhuxJ5ALv5USGaAGDZQ9k2LAL+ZH6pxoo4RjXiThTXKfRm6589ajzE5wusS8XV
UOLFzuBy9OaCe0s/VC4Asmn8WqLPnJzU5FybSNwgsgHnNCXMUy4+GNsdQUfVqwO9EAjwvMewcwRp
rGKr1Rg4sfHfqeJZF5WYTqrjN7Gtk3ypNy6WAXny9DAeyeQo2pcI5tOpqzOqqgGQ1SZYizES1pom
/Y5HiQmKb7RvkG3BvzueWy7MVglU2NSAlQ/xvEkeQlB06FdylUJYyr6Z90czDYlnuhcM2dKRkAJX
XjeOkSwbCfHCtHautszsMXCblVPOUNffPsLlnsf8GAqsKQFSvg229oQhCf7zdflgXGQrGbCfPkNH
R8dPxJComQDTzsW9RKJMbVPzS9cb+jH5KQFeBEfrvht0FrEkg1l5jKJhjAZleXTgbJkWwkdao2RF
MmwLiKSTnsczq8dYIvceC39tbz/8kSVP1BUBG1vkpW8uEmLkoe8uFcjqlAZ11VaGtPGJkUZ5cQZi
fnbYoQZYBM9W/EO62feTW9TSO3FCEEXaNmuPlcokJ14lvkTJD/mot17cedatY2lzXrOI8671tf/y
JP6SsxP6+EscnHW+0H7WSDyAg6sNgJT1Z/HBLsk32yhzZ5Qsc9991kRH2EShPu2OEqcIYj2d/mxU
/4n+UFfdCnQn0Vthz4yl0Ui8hg9VdKWK2u22ikmBYhuzQAZrOTuKDMajJ0R8ud9IdjvWeE4OiWFu
gHOg+H58rE1NLFX0Y8EEhTpQDFQbtoiEApmpVbeit8TkSWvR1K4efzYmubFxyJO0phE363ewLE9h
HoH/7Av54cG2dowfd+lyQ0pkkyLw41Ku260bgbDbVZaxh5MkvcnZNT7nppLa62BhVdzaCG0ldlvl
rAjkfeZt96cG8/ZKKRRcSXFAaib+K5hJ0TZeijFUDFGXD0fTEB+nA/Mcq0R7d+dhvsuAQnKQ+lD4
CR9pa6m/G71laVXe9ApVZ2fq35q0xCLCpTH7ITqWYugDrSpRJbuvjrcBT/2mh/3Odb7I52Ffl+JJ
Jlergj4TYC9/lezqN8IPsx1sqPT5UMBv8U2TV05Aj1xfIEitoUKACLdSbGbYunvE1ZLo0mLl2Na2
otk6HZU74/yZPCNn+2PIlibLS0LY+/oKzT0bwV8N2bJwFSDKpzNU9upzew6HFXC3e4QbVIdHrwto
sPTP+W0BIk+VD8radOJwt7VALcpRexUu2UNA3hkCarPcr0px2a8z1HqoNq94VTMMJ5MaAW8E94u9
ALx3iZzIGqH0cwuVIU6AySn74qpiU2gso7D6ydOQ7LCCMtdQhfHZJjLmYmWJtVXSRcqxnv4zYKhd
IW6Lio8oFa/MUA3hU+2l1XYWl0EkjezTzWLbAjaaiYpBgSCl4DsTXdpd3lTzrtKWuGGMcdOHKhiB
UlTIGPYC3Aga+Vo7bDe6MuMUsH513fmoxUmUSVOm1LAIAG6k7HLxVYH7YQygxK5mKcyta7jYguBG
Xv0KQUevugH6pruvHErBHOWIFUXY9RgH6NZHTkzZ1x9lH0V1LUW2JvTJ7zrmy2443XUMgAb+nj5v
H66AYU7Y50PCaZfwAjQJthsRCRT+UTUmnvFYYFRVC8P+AV2XVtJtGd/gQpOXRwLEBPnshkZ3z81Y
PuDWUg6Spf5TNkJDFBhHYqgqcHXyCfJ/ulssAOXzAtbcIFi2C/glbCA68e1IfZq6bD1L2ilyQd7v
J1Q2q/4mkU/CzRrCawpKWbBGvGAjfYLroc2zsQjigmjZ2QkYihpQFGHuKvjoi+Xp0IiAbkasss3m
47CrxbbGf+ldxWHWFP1noZzipxsPnvu4GpUbR3stuoTa34B5020mXsdkkA5sA8jLgcgN8GBFm01x
D54in9+mvbLvsY6rw5UA5r3L1y+XXdjpa679iZK5ZdttPea+zWERutlkNGK44WSfCwQBa0fd2s+F
kjqxDbOvyXxVNfHz4hZycKeLuDXyij99DUpKts4mGIlA7uZnp7NA+Y/KXzR4gl154feXzvbWY+fr
666hE2Te1tUnUvJWg1WXmMvPHXpCFlLzlsh4hkmHhzOiIF4m0iNLFjRQjSEjdk00T5kNA54I1OZE
Iryy30nSaGjMJaNLrVz3+eu7p39dP2xAjb2Mm9tKASVlOjg4DyUJyu2BNjGX/tDiBl4IV/mANCNB
/6WIDnBIJ3CGasEK+uTQr36f77MatQ9OLUFDhh7gP1dJt8gyQpIn92y4Sx7/KB5u/MA90zw9N7eO
epx52qlXhK6YEqFL83ZJsf5XQp0cl5rG9HSwAXduBE9TkTRoxbLiNRjeWWHTId+qEMWBGRXv6Y59
HzFh62lBRInEcdUXnWJflDYdW3wQJllGhbLHEw+JUFROjnyT0Cv07gEkxIojQo1CQQjeFwDwwnHo
QHAVM7+/xcVBzOiydKpF8+vOWFTDVBCAn53e9NC2vqzyOLgiCSxoGYYGfgwmVPGnB0g9hdVm6Hlf
oWw8nU0Y1dwx+BYpemBjsVdppP4+zYBLHsxTaCnYcoFX9VTexKojKeGqW5W228KCKDL2WhN/48qQ
mXRYuS6jvaIaX5CTsPnvXkYHME6zav01YwRm3ewkP68T4CrFhZAd4sa7wQa+0aw9mym06SQ0fDNN
OIDBsyTVlOfiYxbaWIQLwpKXCxNHWrEkweRgHTqb7ylRaUp2VlD/FrJ2J+4QemjNzNaPGJV2ygZh
CngTjg8pRk+5A4JwCA+yF2MCBKCtBPhRnxdyaB+0e85LMQ8GqbHj/4GZcdQTfLmPVPe5XIT4Y2HK
69jrtxifYYNm7h1Be5QDAFuD3vjHPFaQObtRn2ayKUpgqjzW1dyVd/z3hSjohexOC0Xdoj7yQBdW
V+X73Cq0H4Boi8R68xqFBFstX1iwAsLSnUIOn6z6JftwnyHYwuAMo8I0FG5BTFi0v5TnV6dB/19s
YhoL1y4exa/cmG+jY5jn4CroHGAlmLRzNTYQutRAo2Ve+7zyBHClsQfpX9HG9nM4uJcwR7qL/JiF
X4dX5JZW2KpUirVzR1wuJhXA1tB47FVfV3EdSMg4iiuw68p4aOFIVGgN5BhmnchFLfZkNZgvMbGb
hTIQhLQjfswyW+/LXhurTkrF43zXCJmlL84KIo6mGCsP6urQYECGjwJy+6wOzzrePotLeKWNXP1h
dxToFaw8T5YMuEoBjK0Et4rhBvZL62ZunjyGIk3+eI209rcEw2XNhCYtMkdAtyZIZeFb9vG9NAEo
AdRU/XFxSM2iBkM6b6a57f/VD23vylI1YjoFEvSSk2zmcygFSOfphaKLIijAd12HVe8lQGqrTsVl
Po0q9IPnMZjVut9KThrpXuRgESHEAekaMhJ9bPbn5ep0C2mvhWx+n+ZrrdBsKU4QKR+LZ9by/kwd
500yekhbERPYDb/6MW3vwVbg7nPYQZNfF6kJ24T3yhfo4qLZSzgBWWQt/e4fTTL7VoXE+PuXa2ZP
MQsGksL3JWgL/oMnbOoaV8Z4cy15DEAm5hUdGHC5UTpPgFkSi4xJGc8bcv4R68AvwVahN4vxMsaC
7vAxVfP0WndoPnJqk2KRBdslGJdigf8xe7Ktr3Ly7GiC7MRWKJ1dbwgFfmfeLLKMMCQlpnXhS48t
sRIRywtSmcuhsX1CKPNgG6R0Sh6/yCrwQJBNRM1P4am6NbDzWGw7/QECWTJZMGoE0xWO/91DK5rD
1rdJMM93r+v2ae/iKAiJpiSgt+cq3rXPHluX0F3dFfIOP0knVTqG2HBpvR7Oj+VAN3hPsATZH939
SNU+6TTTaikvNUCJO/9EreLrHB6c1G7H/1eYxK5rAj3SPL//wO7vUjor8ZNC/dYzAQW75PGjCzz7
gmpxRxvFyt1I+6sCbEzzl1McN6eqyKbaLssONmCPKl1wp0wg64NLcsFpkoBSMkHEvU1mI9YrFDiG
fyJvuPhMFxgDxwppV6oGRMO9M0WMn44MDG88weAZCge/4GzboQItXDNh52EYrwzKVhlTfN3RPZPW
ZK01/QDCBNSndlk6yRF9/fF9mQO91guQPnmgiBUnafoypgbwCT8AEvcfiI46vgx95sv28pn99clX
QiLfClGsnAXT3PQQPDto17PKJy8YFxxxJCViy92N3nE4ixszxBzhUOZND3gYMHaKTe55WgzjIykR
MAM6sqUzstOXNlPd9B0cTP7J2iIgFr+i6jMtyNgvkaJEnAV9NQ0y0Tb4Sb//D5lOnjY2y8IjoMeX
odkQTOWVbjLtRD8v4M/t4uzesFexq1oticPH+bET3La2bvoSVpgQHxYLBot7+lRCzqZasr3r2vzL
ul3RQlM7ANiyX1jDuLgQh2KPwz1LVrvD9t9hA0dLG79xIJ6FWZE4vHsjSYoH8wFJHtIyMPpo464r
rWz6MwHNVGlNuOar3xutfSSf3WePI7yV21/SSO0lEJA+Skz+x4v+WdDbE1AdnXFNynygY5ySKFJP
nNf1zxOOSOro1Dy8KiIXVuIEoU3QXs9x8PRrysPnAMQVMqwRsq9I/QCRZwCvo83PIMls6T5BLgQX
mw9GeJmx3Xm2Ea61L+sO+YsTTzw16QuxkNusXJkovRJr+dCUrOCV4pZnmRmb71z/9o7WKHAOgXvb
qmsvn08ABZVmzehN0km6oioWjYWZiZ0jW4tr2tdWkLSyx2AhY/LnwBsCPX2xoy0bGY/678mNM9Yi
fo0CLd0cEF9GZa8Q5O2F7Z52VIgLjRd2ok4a9oCXZYCe/2eIEtA/p2hSJpmJbztHf0RAJA2NiQXC
FlZJNsWL6xQs1Vdn7IQTkzASSIfsmtRe8MtOriaCTa2l/Og0Ly8vLL6GJCxVweETyd1nFF/TAxHv
GZrthyQHm55wfQH7jh8mwJgi0ZRD/PdSQG2v0viJscrUyEkEUVoyHWUORPFjZJgh+5e+FUJn9EK6
pehrpLlbanVyZKHm3g5FyYLSqOD4tZth53gg3NrQTAnphLPwlk2fyPbiT5Nw6fGsJiCiqv/uFx5d
wkUbTTFUcTEZ2Xlvptk2rRCgPj1fxkReXxsC/+gMOQfO9tu55Jp81H0w8TOD/e6xfTdxRPm0/mlp
Ym5DxHg7d0YbEUsXqCHCDemDmp5Qbd1hmEUfra8siYkqenwVJbD3w/qLV+d3Z7obwR9HHRNHMSLP
Z5+ajjwyzbMBOAJuPDmrrcPtOg6f3Q0VoY4+owGVheUGZFQT4AmparDsX6dVDVuNXYJIZXMwvTXT
Ts9My3iB1L+T88HIQ61zMYGeq+er2ztpnMPZylo5PKhg2jANDGSM2v6EXzGhm9k9ANWJdRLewj4M
iktlDTkyPMR8qvaLfamPxRz1pp+vHZumy9EU6PAxP7fgmiggxYTp4t4RusxXXolyHgBvosghlJGU
NuEfY9+bv/kObqCdbk5+oicJYqLJPx495XHk/tuKtdFXZQhE04sxEzJuRtTSx1WMPGVCTFh7g1iq
9UIXORn9BRwEhMJA+1G0kogGDAwoSgmMyiZ++CsIIH/wn19KgR30/gvEInWu0Fp7kpQa4A+y+sD9
uJC60fBgZy+ttcCdzWQy8oUj0LMAjml3G+OlPS0vH4ReNKC2/bZe1yZ3GyWFN3ev+0PPWsm3Iib3
3cBAwnpMizq7WrIGHiQ+tdIyf3hcjynNgUHw1oWpuHOxtBC/uuegqYsHvT+t5fcKSKinl4H/VxOr
CbSJh+eMwQHc8RyWPBnrDXeLI232iAsjUEWtP4H6tqqw5SF0Lcf9ghEHcpzbeI2Pm+bwC954Azix
oFeEnADI3eetiqIfk5JQwy4Z1J2rWSnxhpva77N1/OctW/HeALZ8BVXK1TA8t6yCEtdMT+i4AU1v
tm7jxI8PMIT0gadE1THDGFabp6Ktteyh4yrgYPRtgDrrg7i3mFlzJlL9D7qPefKlajAeFBN4+l/b
gKVzjW5QSsVIx1+7tUsxRqABkRM0Ujw9UvaXhgE+nflNAilRtXC+gRelqMf4zXpX16BOq9QLET1F
MOCVBZOLUT7vAPK64tFOa+ajG1BdxEe9KaQTHGFRUF8C9jwhxrqZLtGQsa+L46SPyD4AC0SdgNJY
alKqtqCoNAsgRVtw/MvHjWHR5uD0ohB59V4vso2sTCtSiBwC9IVypPRvX4DHdaLgYZCkGdq68kw+
lEPG0aprm0N3baMjjWIaHLmZ+iv+O/WqZDhFI1GdMnWnWbsEZ5VwW+d8EY2a4fMjFncGwkVDBeqw
CWKM6NMLo3+WkX6vdH7bEmRGt7Wz2ypiXMF9fJKHazJgfSmUBrS908aDFH+auNMzFW09z62rvRQl
ZqfQF2wt8H2YXMqhbE8HVJQWsgntTB5TjSVOpU+7SndI3ccWSyiKWMY7YSL5JZGIS6AJx4WNW0aU
rfKerjd3GU9B5hiAEfunxlC0eMO/uD5hNFW1Zk8+XMQrKFHA91YG4Y6Nx576pSFpm2LbVrKafvat
qyjaAvBMz3CBRLWatlHd7SRcU/lkccqVjK5GipTHzX4oRU+4V+Hj8UnpqOJA0ZQltyeCFyrc+rk9
TrzfnIFi5Ud+MB1yyYP2zFksZLalfeWojWic0UA6xAOTB3WBghhvC+VugJeVPZtrFxOvF7QTsU3T
tylRJw1sTpK7P0BvGvClFkDQDfbjwkwbz7FKbImyu76WW18ZUrWJLWD48gC+iKifUd0T7GysvuHM
KwUhctEcgTMVC6N25A1a796GJ7VYpZIcTSWv0cKl7bCZD12AgDqhxCALOCtKi7oe3qjvew/BRoP2
4BxIdjKlabIZJw/VE1x9ifEoPvRS1b+IvsEVkBdxnJtmOvaEaxs+iWm92/fmQKnKLz8EBJAWEsSY
FFc1XxAWmkGVUpwpB6sFZ4yenJirEzulC0R/gUi7GyLFjfVAZ2ZUxYSlXlFDF6o+qlC/ZleMoKWm
P2CAHVda4JJIAvvbS1H0SuV0S3CUPWLA/+OjL1rUUMLCwEI69VwpRM+QlHnLsiCd/c2s+nVHmDK4
LX78K4ZxIUIGKwWWCffUy8/peKeK9xw+qAs1ekUFl6S80ausvittZ02PX2E+3x94COb63StLTNsE
bm3W+mEz4e/1gK9mODUxQVlcaiR1LSK0EtH6Ef76zQw8irnn+DB83DeBUCerm3pCyzRbVz6cYGkS
jeJ4Wh5YOGPpqEM2QYPgSR6vRtFa7TzpHs/WUzEOX5tTh/uWQKOawl003N9bcydL6MIwJ14mJlAK
LH0rwynjehQekEPXSHo1n3E4nEMwYR98DYL66kGQNDZl6StIOiZS7y72gtCgpjEzSSs4tjUYlnHL
4Df/zYn8J5uCwelhX4lAy0w1AY9lyV0C8UlXO6FBU6Py0MpsAnNa7oywSf/1lxurZKV1+NjBjCeQ
7uth7Zl9E7ZL25pFslJNd76V3tfs1qA/fY+Q/QTlZ3E0lCIzr4Ab0dXDjvk2sYCWbRpJmS5gE5MZ
Eodnds9P9bk0zQYI5Y+1lqL7O9zigFChmma8mqJikg67SyBsK6CLT+xt8RnzMTY3QSH2mDRVJWps
lKVIzF5x7ZiH2s6shvNfhzAtsUSOgB3D/faB9UaKqBVtkrc8NEYQnGVCtjgLQIAu0nn1ktF/NT8v
4V7UXxyeVsN2vhpb76Us8GH5QFb3YS/RuNUTbXkPjw9j9wNiT97Qe7yVwP+/GW61Sm+T9L6NAbhI
TDCe4CgQcC1PEQnwq+ITlfkWC1oF+dI71Z/xTi7iHmTBko3qcftizHwyodllkM6J8XKulHXqDJmh
kW/T74TdLMt0z2SUpJY+6KqZyQvjc3C96JfqX/e/9bVTHG/VsvRrmGrJUfHNo1MMOAmz2Eug1Ev/
ri5567mMP27ZjYfeRSRpd0lPOakpIExXaVaPQ4hQwBAfmWbp7eQxA5eU3xHdT3+WDfpO2jUo8ZRn
zyPmJ2VO9v/e6nHbldaEE/pL9HojY7J3UYxI3xrf3Nr+3vFnRTwoReMEjDBKSMEvv67XPzQoTOkJ
minOzI0Tphf4iQqhQ990Bw+OnEqdBNer6nzENaeRONElkl+7LzR96nIEaDNrfqeIdlKuP9gjYUvc
tyIxJX6Z7X6c8n84udO4cH9vVpVm8+jsYlGch8y3Vu9YoLe8C2+nq4yqfW50WBlja5g9E1zUAeGC
hjg5Xj0hptchG7CBRvcewJOZieb+08Yf1tmv+LoAaZM4wklGrJSRQx0DSSLMg2zeL4+a5opjH/VU
7ARHWsJb/eWMuM/oB+TLii6nVaEoBEUQnEVwjF8SzKhXhX2aBi34zsTfYEEQXt0aqSn4mOl+aQ4A
nae7xK+jlsrp/hGJO2TTv3qIMXA7Aph4+i/Jv3o3llI8yClCQuOrBf8EPaoE+mxJBWlrHbe83oO0
15yk/F95FAoJ1d0T+S5qbkZHOPm+BLBmhDqCdrxUsF8GFb6kLoLrcL4oKWUKdRc9XR+1J9+Cf9wV
75HWyrxZ18lAGp/xHfDjvsm9TnlnKaW6DcTP7QNWVaVuJMVvfgqMH5AS/raA2Nb4JhagMlXkY4NP
hCwKUgC6w4MUtSpj9Mjy++EYMi0uB2MGqIgzzkkI4UiYZu0UJSoGb810NXxNgP4D1ODIWHmSYTiS
ejYsrx3oudIz65Bs0gtyobVvlhRYyFvYOY3yxNfm6u0Xv2lZS60+kdeSxNHTZ89b7LHaSfoG+3Wg
SHn9+cA5JYvkiol0eXKExU6EI1vUNK5Z4gsEoYPXZJwUF9M264aY2Cwrax0jm01CTlYocvWKei7v
mDgRFN920ZVQdnbB/9XHL+M8c811bJ9yJkRjHRlNz+wny1o3jLLzp3NXHRb9sOoHDFWdSGFk8V7o
S2AqIEGKcM7FdEAu4QGV27HKr0DwkJdKFzu5kPxR5sS8CpGJZwgobSLpsy3WUcPb7uB9vErvKWdy
YcNqCi3HQ29GPTG/a/VCtPBHdsbhLe15Ldc1wOOBh+sNBmU2efzEpElFxUCoXQ9GK5G+EbfBRPzv
PPwKL/7WVOgMI7r/wkc9z/2j2vyivbcXETf1diJ11XFOmXC2g4ZSYb11uzGfo3EuY1z1GVxFVrmn
REI9/V8own+XI7whL4FDEPvZF5+dfmFN7Oiu2M0L8KyrcMCHB6ToYL6qX9ii2Ov3MLbs2pO4YgUH
auxckcMT4cvpjvLfJkE8N9bvaKJOxTFaD75g0mNjWH/JtRABQu3wmaBPrEBzHZPevkZxeXk9LD65
vQQgBu7pFuZPnJXfX0+F8slFe2eUuvwlrR/9vxRUemLUHJnsVaAaWGAeIXiBAZzk/L/RDqMYOdEy
XtMvc/sbFMl7YDWZOZ54PtIN4XO8MH6XZa5HL+3mjWRW+s9G9uXrPv3jkRBslZPmV2tXJZGphDsN
bcf9pwefMpZN0x/sMNXbl1PAaRTtCaG9Plm6ih7s/u0LvMQVw4MUdu4xWOBdY0xuPV0dn4N8nhmH
HuA2CDR2oo3M/T2BToJPYJxXXGNt/qngIw8H+A68RFr4KK16eHBBGP1KyY5XqHi5QUo4+0PB1+kJ
ZjGX8kuSFY98Xh5ilp/GpSVhWkshPgeGWbAM+xSpfsIjhHLV3W8n/yW+clcOM9745FcoTViXuCj8
Cda1UFvnDVDLcxe/otXrvu+yLb4LPa1QRyV07l9wCXsB9LLECCNkY02PTlYUBRrgpFDCS5pLRsjy
NLiH6HFbvlRIWPmbvA3/MgPu1Ub34TStemtXqC97iEvgQHux0CNJMZKjvfaHk1fgtnvTSHlc/vDF
NLArTMSNWRYnhZTd+qWl001/cJHrw/ZvjMoT0q/bo1zfnUxlfHivptCycCGh5aiZtVBrESw0TbNN
qJ+dkXsF3TeW3l9pkCdNjUZmEvwPDBO05fT0zmyyGkGOXPoOT9XdA1IB8ErDNWolZYop0fwwlMHi
dooAr90R3iVHx7U9Qq2evVVz/4/mxeGd+6bWCmEu2YVzvxF9XdbPZ1fYOGqt4ApT7as6K7kRIAIC
z+X4pDojNNrJaeDptaA/5rYw4zg+iPTCQBw9QkgwzirvdNJEmMugV+QW4Ba5BzxF7m3uWsB1tKrA
73ebBy8mzVf6ptLmcUFk/PrEbuVzuWzbwsXvYEa2Wz2DUZP7uedWNHo92UP99rgOnvBcwjvI7k2I
f/LPCYDm6l2rQ8LKsKmCmaVA3ZoOJKqyayD1HBNE/Xl7OZEHY5Uky2DCXo5D8jZoi8ZsOkrMeBes
SMYnUNUKFFYdryPFulZqhydvOenCYSiNrk9/7gdh+BfWYqSNEua1RhiRqiNGjkJrU5fg9VGr4l+x
6pNQ2/RdRwpAZEmQE+IW+FwdXFakap1GhBKhosSZv9/M+Vw91yf0AzQiKP6nFwNkZsrGAruYEJzM
ws1j93k4w8Gby1rDIb1ECwQ+fjTbB70PjQ9M+NWAyYe9II8VN3JITUziuxXIeNFZx7rvfZG222dl
Tq7SysOP/RkSQyRf6eBeeaHZiUhG9nhNzEEjSFdqf+ug52iPFde9bnYZ3w0CAkxiZSQg6i08z10M
FgjGI05XPBtsFH7sgtfk6Vd5mxaFwGyuMylOOJsjmtnLEti3O7f/HOwk9LNoUuse6sdxAV2desTf
JEw7NDA9I+4q7TNwilrzIaQfJCW6VQLDo06+R0D8SEI7tzO1APxALAeNHZ89XzV4/Hvf0B8sDACt
axJyv+VGQjkm65fn3E7D6JdSXWoOS4UDxa/fIaz9ihrrvEcdsBqmdcCT7zMQ1Wdkg7urCHh51IbQ
theJotOkqFJ7AkAOAYQB+des39MXgVj2vU1oiqlI0e37LlTnXof4bMP0hbrj6/ETJWTi35Qc7Owl
mxSFo773brhUQBiaJ+YJ1gKuo6wEL7z8qQ1/Lbaj+G7AQlGNTiMtI6/KUs9Sb6EjHC+6JHWqrKrx
XjIipUR10u+W1Lrb/+qZyVYHU2J3MER0ojcM0K6m8jvKT2uakBJnspIeTwaCPfwIGdSiQ2Tw/d7W
sXgWNoeJ3JXCn5e0AHfrf+e/xRbm1FiISB0LoqDbLbOhGUw5ZvLiOHZgPSo8NaBJQjK0nJEtkiG6
hjuKlDG1II2AdFQdkWG0qMx2u+X9feKl+7b65J5ioFwxy08WD3oXZ8sdmmKXKJ5R6wDXhMufeA7R
gwahmz7c6nl5RKmOAWlCCylMRAFOa6K0UzCBHhcHfD68gQO+LZ+Oim/UDJLrPh2AT/OYqLDblkAF
SDAPcLMnJAjsCW73q1UpcU9MbUfxDSb9O0WahH/1wDrsHshj31EYZkgRKLyDJP+gPC0/bc4ZGksj
hAdC10qIbIRmgJkWh3WDx5C+2c+WAY7ggKBX16LP+GYItsthuNoEwDgmZQwFCQciuhQHM62Ozevu
P87nxQ+vBr0NtBHijIR1RBIjvG7fctdIm/spR/x1jS3r4MYqOYWz0CqOG7D1V+DuPUamRVQ5iGVo
94LjV91tl5fWGAsUt7rgTEgVOw4S434qbQM91T7wZE9PyQFI1gtHephV5xky5PTcN5mhEJHJHd33
WIhzfwQEQkNrVwztk/218vQUh08bhDVPUMc6Tg7JGxgjFVneHo9qG1gdkDYuwmH+LAfSYPGdkCwb
3rTk1UDiSUWHiJsrJZHMxZiqfJusviPjP2vVWvDi0TCRouQnZrl25DObZYjqcc5tNDK+e3Db5a5v
jTb2ucxg5kOefRlZLWBOw3QeGwaM//u8/Dj2nbgOIsUsHudeMHROrMtmaLpvalBcobmhxav0hYau
P9GKSS4+dh9Ck8aTHh/rGgNGdfah7xFHLR0AJovCEDFTEkMEaiGnOuwsJz5J9aN0GBakiVOrBkWe
N+ohMsRaY+CH8rIzIt+q4sdJXLLaqOIxrS0R3ISw7rrJenjmLrmO3i7AKevhM37X2xuyWOCFDB6R
KYKONSKw3iKtA1r4jqaZNj8LEYcFw20RahqbX3sbqHfhuCXaMLOgEKsIKGawwZO+eG6VtSdsW899
8vIiFAHYsYHH+gaw4xeygnJueD99jDEYDvjucm/YuJBM/ZXx8WDYTnutkC5wdH5pyoxC8sAfNOJP
cY5B7ftYdgSMO9KriEFgnKQBVnbAmHPOFl2f3svt862Zxmh8Uuw6hOwtDgckXlHq9GhMaptoZEnb
abqO3lGkoIEwC6xOWqjbyblTm9oDfc0losgS0nctfwQa5OLi5jzhyEaK1QV3EhF3TLTYCa7m4Tm+
QVWZBG/ijBqRpPVpd88HUlSNuDZQbGdcOnr98ZobNaElc9ELDXnFlX4xgn1ilpN7xr4DUTBhtjrn
WzTgmFzY7qlbHRUQJJVkYCFuG6P3moDI46vfTIKgoppxD9irRoT35i62NY8KVfgzYz1fKP7BdS3/
lYrvZGb+aGJejlMJcv2NuRPRmZyxPwzqUamv5SSc8zICH6o5sok5MOTDGdthjqoOunrQewT1Ivci
WGnBgCBsx3sLcRiJSkCbxKlKp36Fr/9jIgGrqFxt4allyNQWggc6f4RVQmnEAyLLBPgn9/WX7zAr
j5HhI/DSasf2nGp5GOomEenIGzTTMuNMHScmLm14WOYDyJ40FVjSNvYWBrFW8Nxlxm2JMDnxt/3O
/7WTpy0SpQXJvdHIGLUCqrIKlvKLEsxNDE6lyMwA4a0yATisx6b8un4bjSyLGbE3zFsNx9PJDjzc
l24Rlsl+M50J7XZUj+cDefHkehP0yNecbfB0fPLDxF/kaMvNza+dgZRIK2YIE1IuJnaLdviEMxg2
Hp0f6wEbaqpNeCm0RJcgCGYeOvZyz8aOorZgu70hBbVQtiu1bgTjwBLVnO0qxRDpU0bUxeXiXkQL
Qp0n0iSV7b3ZnA4/79lBcYaXdBC84YjmSu48JPCytonfW369sYEkxshlQ0zTpboT6dMOe3RS9FYL
zyJcF5MiE8E0Fpcz7+JTC5Bs18kumQuAhqpFUmq0DNP/+xDKK1P0+8MPZvSjrdWybCx9wd7/S7p7
5N2rEbybw6i9B08B1GoQeO8iZ6r5kBJpgEHZgvaJ7P/H+PV8B7CKj2iWQTLZHtM9SrfnwKcjm6G8
9TuDIe6hzpGzBW9qUzTBEBKaWsEwnJeYlBG0k12UQXcanNTUwy0Unv6+6+H30TCPlqOYyzOUtj2V
fxuhBXJXk2Q+6Fr66io/0ZNK4aWi/2QyAwlxbuYc2O58Mv3r5ifcKmwMkdgk5+xDZn7Ny0CEANX/
AL0tCAEw7bh4WYmv+6DiK5FAgQNTHNjVwyIuHwug2EPoAl5VGve4XmzP9PMTbcfmsdbWXOZwtnS7
KINkqVRVhMKBAUHc8v2gbziVq03Lo4DTdayjdbC4cm3hhM2EyrEs/kVlLPToqErvbuJK0jHcCaDo
SIOOaGQ45U48nTMUJJu3JVMaay9cm4r+RpzJ9bcL4xTkhAdenu2wMPtP/BtkGO965gLxD9KXxcc4
2gtD7BSORtY3N+RtysyAbGcK55mu5W9RY/syzxcktDhygfH7q3gJGWdC4iRVlo4wrcOvrGUAOsJ3
HifD1onfTMW642PsUbLsXathvhJbWimK0EoaQFGBl2yiI/+1RZwsbrq2CNT2dh74I6mCnK8lqC24
ueWMN5to4hJK1RpbJeqPiV6e9eBVib9cgZ7fRl5ez56L7fDcbiBwALvaoTe2S+wE6IRRhGVFLwvb
ObQZ+p+o0auktpBd0xHKyalAseuzYMoxFWt4T7ElgY2Ldc6mHJEHx+FZCykjuDLA+kJNhluPsvTH
Vf1tJiB8vSwjpDxvA/PDDKlVp7dTdxisslvtPjESeWt/FnACRqUuJ9Uo3GSww1vKFSGPL/hjlf2X
CrzNoEln1aI8rZCGi5ew59Cyz0zZiWNjMURS6iAgigIt4cFrXk1ONz7KCaHFuYwEAfG2o894Laid
1mfrQAWM6oGDy6EbBlDIaRgED17D+ezXOSG2VwhVG0568mfb2d8S0xjMc+KuQvl/xhFquvRiqBno
yLrKCf7hR+t9MSO67syWmZffO/VtEsY4/IQHk3L/IUFBAPup1TomxsKzybLZY4EeGoHcPqUJFBFv
g77DjcPSwdkCQowkX96dnihOPoT6zZaEfuA8+x8HUB7vKSdnf8A/jaC6fAF7xXLZKumdFdksZM8g
gUazD1jN043joTA/fd+1ezdpxxoRysUZtn1uvi5t7lzEVP2YcrWsiEQ5YOvEgBqnkp0ToYFscERx
VSGcbO2kmdipmbC889hx/9bFdVl5S7p2Ew6bXk3iPVFKRt0l3EiRiORE3c1jJO+PYZ1M4KVUwjzH
6rpDHDHTUXJaxgo2H4ifdyaaIm1kIfclaDk6dqAWX1vHCPH9OrEsCmK2MzhU3uugNC4pGuD/BxKf
YAESmIKtyJUDtgoKpjk9wcuue7XBDw10YdIinmKDkCkITsR6YuB8yuBPGZN18JAlWB4P9BgjSaEl
ic4bVl0RCnvGaozmvRFTtajrrgfdI0Oqn0U2g5SHQgEVN5LYgx1qoVMQeG4s856+HzjDEZtnT9du
opCL3UctJN4ArrQZ7h+wVUBNWZuktWz4OEX0XLd270duPJhx0MzWt0lXo9tgi4QajnR4PNOrExyp
in9DcKSD0rsoIgvK33dy7R7JyS33TwSqYwR+tZhbON326cigyRobG5RD9WIuzfmj/8hF9G7ipHjS
UFkwVAwEk2UBtyiISngSGiIA48H3aVGWPeeljnynHrjoWwzHjwGAGq88Ss3EGJm263KyFJ24WODi
2H+XEExbc1KzKsIpe747sBk3dbuSPDhx7oAScj6FqIO2QfxTHQdeda2bhGdqSqyVEb113er+7vuo
RV/EY9prCtJTQbeD4Bf/W8lxYQwY0OMR853Vv3GBJsSqbZOJ7MOgNLVVDWpbIESixQsU/lHOD60T
GFcF+12rWGQSygV/4uS8xQHV/HKdXT5KxHYfsnmBeibWCuRoivUAkARsv1W0gfyWeG+PhxpF9tVq
KF/MRgt+lnbHinLCkNaWvOtpuq5NmXszBQkvm4sjODi/CjleMUhpd4W5w6+6YFbtmnNCAfmNUJnM
MbfbrIw9p0u1zLMXUmdiaHZ5r0dktpIXpeKbxuC4eMl0y45RaMGKXWvj0+wiL4q3YatnvjjwKin4
47K8KjVoU98kObOe7OJqXhz5dAP+u7pMxnDKHq89M7PUVo1+0ILL+S2adzWLADl6GQdBlt6TVgKs
WIO+oMxs7A6YFnvhQor8g4CDe9YXmfe1puSidMq1nCgU+D9x0mpGxYZ/X//H+GvFpSlLz+l42sDU
N1S0X1NFxl3WlhZB06TTXjnU+2KeKSGihP/r57EMyj7Xi6r7hhHEE/br9CNY/lNJvjo1CCea9+YD
xWkU4NN128EeFDbO78ZtOyFvt5wekGBv/YUMCLfIHZaI3bmwnwE+Q0lE102zuQg+fVDSChGaK5jA
K3LiOUeCtW52iFFJjWtH0rU6UUWsEPoOMdkiTMrHts3HW0QEbpm+OtbxNnXql33u35BZ+Wr+Ws7A
22YKxTlxLhtcaeGxYMixiF7w4REXBJRgW48ZyTcmcivvv5rzYUvnFgxC9n0pjX55ShZfn3mmP70u
Q8U2OfNccFODbmNNj65RkqxBkueYWvtcvkRA/GFj4poE/69abNb4iYyesvhuQHG2daGc6ymliZHS
ucICeQU9H5P8sKIlHPNPUd1Dx1q/RAaC3lz2kv68Gqa8HfdRInwfiJO16ZPkJjmzc9u5Sb6kLT3R
Oqw1iw3wgCvTofxJlLMcGDn1G7E2XQ0WVTrOmqvA/BRzSUFxrxxcXzGmx243IbuowfGMUBusyasV
Kmge8BtdTlkfWhOiLH15AEYIhikIzl4JDea0m2YFTR3yrRYLrleaaXM9fFH0dBOlNtR0t2Lq3sA3
L4/Anv3dn/JCNz8PBGe4wFvy+35NAfP4JSCeqsPTGED5LcyopzGiCc9YA/qxUQf01bCvnA+ar8Fm
xLN9XkHaQhIVAlQNY6kDCzwazK1cMxScu6oeq5vNtFXxRRw/Y9wqARaLV5Q73XA2TsdOBhorxKPE
OsCEzyy0lD1uJc/iSytH+uHQJZAxuA0wtB3axEWS9EQJpoytuOxMx2Zr6wS72diJq92ba/PLzkiU
GgMuD2K6HhU0l0eW0tcBupl0A8JcZQZxRo6rdGa+IjzRyA/dgZ+ncwIWIt1BXXNOP9UCqt4lCAax
nSLIUrQJcuqGMe5eJsiy423VGQfgyvYltxV5xXcZwa4MBdR+YLKtILl9NPUtdud3VT57WITLXJ2z
vMf/Jl59sDbLxJC8gWWBLXMWLs393baDzY8hkEVbP6l1E5RtrDZkADUAZcroqQVV6Vr1ehHSEfOv
fWxQWXDmZdlxIo/bR7RNnxs9RpN5GIlX2l04evCEZdGM5aurIleFhJVZY0lMDPFpfO3I4/uTZ5HC
HIfOVq1at230tSIoZChsuLSt+oaOSp2PC0MbUL6zt/QLPprOC6ac5So1RbzFlVLGZj+fk2nJQFDe
W7BwGGsnA1xNt4WRcW2R3Es+yMV026Yb03yhvAX326Of8aHtqDIe8likjzPLzMbTaZecL+LCnlaT
uAHv6eSP/JVaQCDInZSIBc2GgN2OvgHWPDCXVmVAwgsG9niyfAC+sVjXSDhVqXaWL83/b/qJZz2/
SL7SxDtL3WHn4BtO8KXylO+dVbrSz0elpkfSuraPXCrawTgrZJM+puzQoq6jGxDc5VhxVPPu/Mkq
Rfkbgs6ksgYy5NkDfdt97BYGrRvMan0apqO0F5bn8IXXP+FfogRwgRWJrN/noiW89KA/GYavGe3j
mmv4P46+ZCuXxQOS4cjmAHIwVTXWdkIoOXqhL1uWebTWNqcJZ8bNomqZg7Sr8P/1kTNetVsp35ad
EAEj0Bya3JwRYOOuxuadBnIWbIiahZfPU169GSNZcMsB3Kt4ue4wxq0zJJGxNg/+uZPb36nR4fwz
tSzHkfOGlXZYtk7yUDooiyBqXhT3G5LQJEGIvH6c5IbVFEL8WK1TM6mLPKTLLxX5aYrhaqPEBiCO
ExgpmdbQekptTkKtja8z0OJuSz7xbLYQj9CDOi/D8INSzNwqzES709hNnZfVCK7dkQ6t98OgoLEt
vceR9338j5ToE8KUNjXSf3VuBWIu1UmBxfpi+T0JTmJYEqrOjJqROfHyrmpR7guPn/75/HlvXsWO
BgHhm4HoyEsaPYEqarwjlmxggQmw6a1i7ZWSWprFk+xmRt3glL0wnBBk4/6wPGWiDY1XH5aufLfc
RFnz5+sOeE+vrp6Ww10I2R6XsklxWCpfxaTY1Fs8NAi08YGd/UWMZpZDAoaF6Dul1GvKw+/T47HW
fj2RRubeqaywFIEtk/XqLrkjM+QOI6C/ACE4Lzu1PTGAPDg0pEZl1Ri1U+fhDkZfidd2ZICCqYpL
87SjmgJ5SyTdKaG/nNlfxzg7RGi6Ewvlomup23o8hiekAn+I4NmxyRi9nhibQxqNWTrZKW52f4jO
gVF214IItAOoWXMwabm0y+G8Zu9ZT68DwMTaqHRY8ciL7O7d8LW9HF7cJrPXTknAmKbDaG44BS/c
ZIrAEJHjbiFAoD+BfkBlRNq3H9Qeal8QWs3vmZmWgs0VPZCnJ1SsGYvS4tMB3nFIa3Qpmntxcjbw
nuS+mk0Nv6uA6XuyEcFO3M4mA50ZzJ+Xj4TfFEk4OJnecXl0LKmZpjg8Z713FYzAfD58BCvWEFAn
AMClZWifM7L7omQx2rFTXM7BmdujvU2TzjLFTuJWXQ66EVnDKAzBTWyjvJkdzkB5RQ2SQtsKMcL8
4NSRuiEHA9zVXpAapKXuWfL6AD0ri5rND9ZyUBVbPyE8uo9AHZK4ZJ0QZy40aINPJtBOBbZN/RXD
0AivYxNCrhib9kpr0ohDYrjiZRgn7k4OzMpIraq9D7KFuOu/6zZcsHh5BsJ5y8l6RX0dLAJZI5ZY
DagtZDXLHOC+5N20vxWWB80XCsIHmqE2Gnn5HrLGnOqavMUTwWo+Q/w+lQvi/n5UOJDlRwkmas/Q
Z/wIuT5zqC/LEREgRepMHj/NpjuvoWZ+dr/A9DS0pTOALhQZnvaR3/q9NC/trPhWzQH/rH+Nd23g
uPnDBzTF9sd3Jk6hiPZRZziot9+ecP9CmL5TctsaABz0/bFxI5LCe7Fbva6M0Y6Gjl1XngZJ8FuV
VCD63KVn4GOcuF7tstUIH9J9UP2aoZjlT9VUFM5FYh20WezEdMEGcDlBx4vbh1ajDIWqVrhLTTPH
wXgfH3My2X6RP0cstw6o847rK2tAoHwGRTj+5WR22ifBzkoKwIYbdbm/goO1nFQiedBAUBI/rhot
HYw/QGtpoRt2xIHjn7/CcwnsycSV86jds0bjWkpN64VZIsKTXPscR14IhgTQeNyoKPKVlOYCamDi
lyXNKQ4AdA8C0Uhps+FUmjbReowgoLQlxMDSXam8SbeKMW15cRHskLsIOCJFOLbfw578V+YJ6/LN
dbqkieUEQiIjpn/nKLpKRfm46QyrUZlm8lvgo77CZoegRKbDpRwSSno1gywLPTSaLmEg85yE4T21
df92BKw0gVw7TQ5IB8oN65VBDJsnEo7wDlAc6dMQUp+rCICjahSLMNH/22QcjagHkcdO7H8IGDIe
uZd7H1vzcYnamAkdAhUZMv0SV0EI4PyLmMibU5IrlSMlZiWNjvtRQs1b9+kvZ7tEh8afFeWCSIAK
O50dD7x2JQUjNkeLKCT1UfJ7RX/AxP+HOSZahLCHwty5FOYzlzriy8bnk4B5baxkKmEChURmwJ0S
D38rw1bxxf8UJhcUod3hXYEyhK0Jk84kxd/p9VYBBKKcQY3BlhI7o2ugcAqhHWlysjhZWJAEU/tj
8NNGKTu7B0GA33BV2S4qEOHSTdf1QnIX7y/vSp5m4iJWOFterIMsNuaw8zwS9F0Q0c8pVy692LMl
vRZtQbfFBJ22s2kVBT8a6b/8CrGyk2FwG3yhLru/C0Q6nZKBHDSZyttG3mHMat2IoixWpBnIrAyW
Lv7rI4KKo/P46zagfMw6c52FxiCkXtZuySneMITaFrPznyhyz1NOKxcfqxPIqal+bAgmkxbsBPMO
9FsYpzTAW1cM9pbGShUd/ceXz/N0FKjnrfrY5dJ8p7OXimGs7rnFEwPgM7QDCmRt8N+uOopLm0y3
ZJyoC7OPcVmjRiLuKHwsjKE8PbqeCigBNJQDi1ng3WDg0eVbOEHPHB7jBu2hhSQtOSEfJ3jkG7p/
QS6dYyiwCMV39W9EyfkxVLqb1wa/+fube+5UgdRK7yaCWlCwzRkDRkVngk0iB3oEN19lshYFwD3r
Sus1nusSrWBd3SLyoh2QU9fGzqbLS7fcO+IbAdcs6HAxTEYyLVSBFelzpI217dQ2Z8gOCqElYGFG
JMQpGToZweo3qlixJ8eg9P3kwUv721XdjyvKWvj1UseV1Xl064UWWnchj92k0Q4sW3bJSxeeEPtj
/cSg9QhCvCUtJspPM0k8rnDdMf3V9S4VU6Drv1U4VDeIuTHbonNcLvAtvM6NzBUsRGN+Fjs8L4Ma
497cca9orD0ZlLs+vImJmX2tIvB3gPBEG3Jvzs5Jybqr/hW+5/BYiP8zBFGiIoYyWOKB+YTuPg17
UHKM1AQeph3vmLt+xKieBd0LQE9Fn1AcPKLFE9oNJCqP8+ATBhWSChLV0MXJSNxvQWP7oqnHrYsI
kjat77t1wTF9GrPcVHxy1+OVm5mjshVBOU8y4HnO0h/oOR4sEd0wc/VSqTWstWFNTbP1590JS1mF
Di0M3sotXg7L/3Jo3NNG2337kvmPbqDHqVm8d51cwvkNbJIZOMQws7nCH9g2XVVWR+pYL91V4TWA
lw4JJmrx/9C3HST4J1KxBejHqsstpYwq2+Lv/GisUKTy0L3YCnzP6ecLue+N0YExpIKVwMnIhAYW
lKvH/C6cUxCJU/FwmzIPEpGJ7gaUVcdaUS9qlSQ8H+uea7GUK5sT/SyaXyQk4DqBgGSYHwS66dxU
NsVDgo1eX9JEc74OeOTAFMyex2NnG94VreIIYFdijmU/BoM3FRHaoq9AfLiBXqupWjdGhz+xhp2i
ULShQvv4rLYhBLwjVgn1HrRGK7bGUfT7ZvplT3CUkXVCeVDdvEFitMVhYUboTZIeMfxGKJujSXst
ZvGFphZLP5KJjvtoOXon+RSMmMATROngWcEM4kHiovGZV3MDTaK1H1IHqXNqXvcuURb++IeucTx9
qYQ3+VY30WbLCcggVGLgZCNN/nLxsKZJUgeYJEbfpeMbb9RlNzEm0fTp0faNNV0zsKtZS7FW/1ZQ
woi7QaY52vupoQGEKkyBAYZqrceHXp2YL8FMvrASOWg00n5zsc1WHItTfp9n735kZkreHqu25B44
b2rlh5DKTgYMHYqnlVLpomTkCb08QUAMNSu/sm0YrYtfY4aHw7hBzBdoxx9MGHgBPFQ2V45hvhUS
qEA1chaVcCMqVZwaZYPrUe7+VH8TliEwK1d3myT0kF/Zg5kHmnM47KKrOFF/gKtB/BZZRdMF9rAd
AKSpecz9STiI1vYcXq2MALzJ+wKDy+GrdR8m9pkJRPUa3IaBv4LpFVDdHHYRDHhMmXBMkqgMdbD9
VflzajWGICK8MUdS18GhmI4IHY7yCNA4xBxmUmHjqTBKqDGS7aWBE4qC9/8uTfxU2q7C3fvgoglJ
9D8tWL5S2eYSHOmxFDCUdiK+6bExGK+n/LWSAWGP00rDVk6b6VXxJI0No09JTBgUQYCQP7DyKYiU
LynuWV3fRYr2+EDfvZWEU4jxMA0B6wAZQXIPuoRjjQ7sUd9eZpD3PAg9h2OPFcy87zGwym4HTtkq
UAJY4lRn0MQutFU9WCVl2sE5ohroLYF5vokJGn+IPlukKCRX9veg5l/ZIYNiQq6wIUDBfRPhyqRo
F/jqfsuZy1KXruYe52tw1+81ZQmFo0/9iaaYfSTherV0bfrv5t7h8NxA4nNbS1x0yd5xirpYiU4f
cpXe3CtqhmaptYdpWBOmCgFjp42X6nzAdSgLVwgOIN0IHklK1aSSSZtwxS+CT+SzuPhr4VGxRvlS
6t4llymw++FrVhCh4Z66w5yXMaxJjeC+/E5qTcx4+EwnSweb5ft1wOe+RcjWh7RBEQvnDcAWhzaa
EDzWsSdXlIQRPDJb/AZOhIq8tI7fZOagOIF4CACE9U56KDzZk2axriFIl2dBZRIDFR0RCYaGWPZL
dRLeOBLjjx7QzjkdcqqTY+vTiH9R4kqv1MEdGDEBb8rc5zWV5UBv84UQaO4PXcoBEem5ULKtcwvj
JUIP90zrk5vLJkrOR8Gz3fiiKwOJsWinVLJ4EfOZhN6YucyuqNthD6wP84LzpKTUL0SfI9KaB95+
jzjCssovzV4iH2dZfosm4VyCrSVMOk433Ujje0X8ddqRFRRfxepnQT3ogkz3gwuk2DdbH8Y05QOQ
MuYIWEMypffzOf/xgdbIwSQ+Wu6gvz5grEsWBVHWTrtvUQ0omP/baoouwh5bo97yQ3seKrdeUiiF
E8nhdZf64NdmD+qK/A7G48KqzWLXclXWv+QLfBNSaTmOMC9cWElDBVkNSsDhYqm2frl9k9Et8GoD
JCsKaLDQnzK2K4P/XfGWAnBDpFlqtdwrQvjywsSPpkb9WT4ziOA5UcymoUxtM0hxX3KeFWhhiTaq
gzMVrKYAuy/8O+lFi/pawwePSkWyAKTA4g0loYHErMWizTw4WWzcJWleZ1nehl/RNL+9vcL99X8z
WQGWyLuFM4nSLdkTlx9zvune1oDIByfnlDSpV9E7/+uoBfvAV5xOmuBXJt5v5La7H3agaQH7VBPh
e8MhDli/zAr5LVy73PANRINuU8CAUGciV4SXwRRU1//MHyuU1J9AYPMxgs8Wg10RE1FgED3rsEzr
GSYTaMeMwMiRwQC4PQn2t3b5nhtRy6j5g2BGX0l8gCurWtfI2j3qg9FPRrgBWBlkSBio1CXgZSFd
TNPLuFtoc8/OkG/QQ8cziCpwSuoqaEPqB/HjkshW5yeMy8FOyWOCuficY8YgxxgFxz1k6/71xNwr
QTjC56ImlgCjc1Pqaa8U6B+IggnKI7x7Av945bcG5BMdSouZ4T+r3AjXnC7z4b4DiY7OZcDCCfn1
CpLNPf89wG/mhVpE7AsE5LPSlu4XrNS9ACrtmVV8/lWGqZz14fArcRPNKQ037gfhoGBu0YXQmdnP
bHtmvQWEzMyjgxYgGygC8JafuM2WMiaxryGroYILSO1c9UEC1wo/DQcu+ON4QVPQay4zEI+iB5vG
3ZQXWBgMcG2MmckbnNkVWqvvnIrmK4EOIOyCNQiLVhs0nHRBOxS4zaiNgZx7xyFmPCnkTyZaxlhx
B0kZhgBmNf0DoQX6UC3ZNyES0SxxhMeEtmHgX2mB3CNnqIR8KanDEjwuFnVN+JbU3BklkC/s/nO5
SuN31O4EUOG3307vARukVMTIp5BJuJopSFUh3jNVpC9qn6OEx8YTbeqDdOc2i94HIxrjogEraDCl
U2Gk9IVi1898TsKtj4yn1tXnZs6+H0ag5Q0RaP0xZKabixftfXdwB0urEOtIcTdcYpZXzY58xqmy
rjKZutJH1TSD8mqabO7HOkcGoz9BY6JQkVEeUSlNGGK5ROOiRubM69PAC0gQ920ywWO74vp03tXJ
ZA8NYzrmnL0u6hc4Eioo9VEBar6M2sqZOACzO4ndeCTPgKWrUJ3jQ+7jW/LaclOts0CpiEzq1BxX
xJjAfAO+wU8nQRz3Eg1jmbb/opHbnBjkBe8pfOxU4ZqxdGNMgTsYW/VnloVl1dN30+8dIil0xQqg
LvV2nyZ+e8lR4dMhR+r8ZpL8MC+vWSjY33+9Ss9ynTSG5DeE2ycaBSVukeV11WBHnCbQ36F+iMZ3
E3yvO8q0weIj7DfudJPuHLcBAYp0tgc+pxpx727nrOhrFijIdbPWS1QV4qtxOMj3p5KYG1NlOuKf
bguKo1NXRM730kp3j7HZjXQm0yOh39LCn2dCD/KSvvSR7qB6cgfXubNINecBEMjA+YjflM+q67b0
hS10wYZ44N3AxfdTToK3XxNMmjLmVLF7GxfQr+CVY+RJPWxfNbIhoQj9iFgkLayzZ9m2Q8iMmvwn
wQcr1DGsvSXWwqA6o3SiLpcPUAMPDMS0SBTusjZJABLq4IPjiKQEX5GoigkyyeEUiqk/gj46GCTk
SeRPAJwtgzg3IRa7/FHbk9cdsMvNuklJL0FH1MAMC+QbQuIsftjlMQx+Pqenqz0Bpz6XsbtbSYcU
y0pKvUGPlEsSPCb0BMdWVb7+j+87ziPqUxXJsjXUCOoDZaYu6cDYVTkGiLocXRpYcu2pZ9YwKs5m
k1+BhdMPJEjb/bYznY7g7lKvyrQRZFZtzodfkSiyQcDYVolFZk+r6PDbC2UNI2UxOlw2UiI57NyM
5vwOJH8IkiibO7vxntd1yJoGbopJJ7RA730HSZsdd6LafxlWv1LRWDK4ox2fWh4dCY1c/LXxp865
7q2FeavPyii1Q7tdP2tOwFbAu8J11zPot18iEeZckNOaXsk8tZE5DUFomnzx3rZD3+BK1rPy8025
ZEbPIgVVpfxCj1PBC7sq6oMx4wjtCwQL0N0r40XDX9LYtzLf7He4EJadKSEKRcpWNjhlcqZs+Xiv
TXh3g6v5Yn+IlABDBJkXdmL42UMuAq1t/lZMS8CEZuy2MahcjI6ysizuAIonTvoAOrpD/w0obih1
ACUemQj9uTa6oda2QvWv9R/rlPQIzubQHX0f5ocWvyXA+UXyaeggbhlt8gybpURQFYZy30iJt5Zv
Asw7G9V2NQll+BWWRvNNnf3exWJLP6YieN3eXy2sxyVoXg/kX0+f4c/ICPcgv0w7MJ0SvJSmv8Ue
JO2muGKhMXPkC2N1xri6uho2nt7Jh8xzH3hiqUE0OZKKfJWLCuphiRDwCfsMo36HN77XTu099Fz+
atDOyDzo5BHLNmH0VQRBWUyawAZqoPFdslEAx/PuGj1Kv/mH8MgDHvoMmeJy/cmrWQvtHxoNGRsB
ihHaOl5u7PnIYHMRNhH2SK16sF56b7Vr1HMM8eFvHLbK3gZ6T+M2dPyyoV9s0AjnoPIdMj+pLppv
oOnbkgIWem8xW1ClieLI+b7mt3gh2dQwpxDvqScmVwu4FnRCWlsGR9nbMpAZeAJiqNET04XTqFzJ
794wkzZ2sAofgrjjZNTTS46MGDdGDgQyXmwyReGZdFIIm6wYhnrWGf++INdW/3+uWyRzXZOFGY8N
4pHlHzDa4j7FkcxfQRtbKxtWITOHmKkyla/6hveuz8yaXTgsGfLyJld73BijAJDwf4/Sumq7M9OE
gcHMdZz/cWs0RuDKzABrwyIzh/oyDrpCufHVilyhV0t45kOsxUT4nEOKNZZyWklVrtlf3wusRWu1
QTtTsIjk4awFYU9lTyGDo2XU/3D+miayAlT6J7JbYiGV6i3Todl62Xj5+7QsEk7BGVD1YcVKU5p5
HObKjwfebxZuivc/0UeasIrTyz9XeLC4ziI5e0jRjM+GaRVlcIpPMR7t1z2uYRy7BueCYqSblPic
Ot9u4aGGdO7WH8xQL1GETejuiDB90RbMY/JXTFWvsFz8yZ3+AuxUhkakFuxJhU+gqN6vtI9m+11K
aAETxNb5YF+8IP6XJhxY30wqM93OSUUyC2OCUqgp8s/BNLc+4wOPR2zGQQlqVFPZpSHkxOJPnjLY
BsyGyU6sGqxhzGyeXStqXwIhYGdi9xBy1te6a731fs0EiNygQgxkmrQTHF+VzionVqNAqsL0zPGt
RbSHjQnVoumCVbQO2Fbs0Iv0NC6JC9ikfUiej+GKzdBbk3Rc51x31HxTtp+BMvWzIiQy4MH7ATO3
uTrUL2Q9R6bXnWWdPymqiL921hJRIq+y1kLdPOViaVUIDtptqCRitEsZWfIfGZlmWqLm9Y5Wu2jk
2JwrozWTcAFyiobj6DaXLWGAQDUjwKVP1qrqzmA+6OR59leb2hsKmyv2EGriCg6VdX7YjaoAnZqZ
hRCH/VHRH/EkYz4cHnj0RsRdgOmR/EZm0PWttCAi8ll2UPPpYWZPQMPLAGazBNk4z65xHZDSPMQH
E4nvRg83I6gR2lm5WkfrTq1fQeeoHH8M57DKDXnL921SHKewlBDZTLiuwy4jZ87bmAAlAWhL+Iml
zgj9h5on/Cz7/RmfYa3GUDiUmNEBFAvzpvBPeXJfXcPzxNxXY9/nNW99JTvrOgPPe0x9OTSJfxcd
t0e3wYVK3+siV5W3z3KqwI800Lg9kvQ86+W1HtRC7JuiVtCSWWKuiHsIQlMHFJ4/4md+H1xS1KfM
vch5un+FqmlohPAT4ZvnH/N0yFEZyhBiWev1YzT6XCXs5vtGZwf5LVpRwmJQ1nFn3PjrUqe1AaYM
kOv0aEvL/0fQWecjep5FsbHZdp22aljbGw+mS4yp+HkTi1y2/YHnaOpfBnrMtWSqPlapI7w4XP8C
oL5oMZ0d8UqxS6pchSKy6q9PpD2oylCg9Xz10rMgesHX/49SbC5WBDv1+5wuuLR12olVBprr4RSL
oLM8APqyFECJLh08ohK6zE4glFMSuuiiRHvjV+mSYmHYSLnu4vvW7JzDGthLrLDPTRfTFXIEXN+0
MuEPZs1k3PUSrYrRYK1qYYyaDzpk3UCc0f2HoAMY1iDx603KTjMTHqGOZJ8osMcQGVeE8dPZ6kLw
XxXsAjUB2/dP882tNAha1xtkd+66xFPpEvdeTBDpisVXneGUSdLQfEqT8ftq65CEUOHKDCg+pO7d
A73ktWOebahDO9OPXLMLizSONKvy6vsqJl7Dw9x5F7ttbHtOx2IURcBbvyvRgMYXqZc1F+ko7g+b
1q4bL4saT1bo31yIV/THIwSCkf+wSbwcRPqKiKOY8Zyu1DwnX1lVVCAlUcEQTujB5Kobk6QE9G9G
QRYq7JG+4q1o2QQgYARUsMWJ8VlLMxubkLuQa8QoE1at7++BDF7UiflaOUe8ASnHgqeE7VskPw4Z
muqhybGPMdHbWNj/nTKbEiv6X8BpytnXK+7VBrgvKiCMxBdHTfX+7DNRvqjlzZ+XfRyvcPKWollq
R47fwvmkLiSE22xZiu9sO1PNKneTbuDWNADMm2YanoY9sJXExCZts47BXE8Pgq+boUe9XywU1Bof
YeJyrQM0hhswd9QIPtdounp93uMU1qFp0jjMzSIyoDAYn2lpqMq22u0YftVkJKaLuTm69VqpgcNo
NMYYV4LFdLbh3xIVv04Th6uz2YF8+EJYSjOJ6+gVDfWxIo11VmUoh4pi32tkM7pePaahAjW+U0/5
82xKxbOAsUFywn2px+V0Kl4pyFk5VQgY2a3HeOqhTSXmZxBZugz7sBlpxbjpb8+TOdImIG2UjLmU
zxbZT6wYLIsRyyxjIt/OF3JeE4CCPwyTQ+Jc+EUqmN3Eo0j0ksMQuhDxfZqekykrKEr6r0XCaFkR
eiM/IAy7qsHWlzHOis7gFbQrUlTZ5Y9VXAf0bKtK2Xw++rO61XswO9yqvnVNlrz3tIGVwSyAtKkm
0y2B6CzkeSqNApu14x1B+kaY5lvr65SJtxK9FyLVC9uPvifqlMRmjfr1bbfyzfN/Kb5Sq4Ru0W8K
0i99SzmRfqHWyyZrDo2sdVNdJjQiGdjcv2sGmFhezufQ4/RdLDrex3F4cliqq0CkMoyFoJKc6zC9
GS9NPjseZu1j9h/duXRvFdragcGIfbcZlnQWif49XCyUBUpmtPsuH6F+481XXrx70ZZ0fcjtO1xa
VS3l1FAVZtoT3VeKgPxmwydwIy/aHS/jbhAKeLSeJSPpE5QdEG7mXeUqSWjaveS6xwwo0PqQhmRX
P6iTPArjGLSBDUYrMNmwK6IUuzXYUA35GuPaAVWBvQz2apwZeHeAa3QOzjTyJXOR5Q2NJ1Jlw2sJ
Evl1bZrJ4X7vpisDPqzY5dr7rXJ5QHchmRcI4Yo+7vb/ZiAwvdXqwfn+UHtc1xOM0Q0Qy3uVhyJb
8rUKVujhXpPE3ymYiq4SU5+L1Hw1/Mp3Sb2nq5dUJTkpUGUDPV10NOTu6uQeJbjlUwN4LYY2Dkhv
NUOZ/N+bAEtNfkabRfBtS+YLeP2ORnWhaUvW4uwH3yjZlrVTd4LA8n+TIGO3pJhw/TYSGg6uDCPT
MjNCwTwrSFVsljXfDztKNVxnM4sLf+f7+yhvqBSaBAjxK36HUD2EbLc80fH7Yp5BwRjnSNM92B1a
DXIiBvd12faUt23SkpKHt+mE6OVVJN7veSywtFAi918hqjDsAWG5ilBN6rlX3SK+kwemh/wOn5OT
7AkRjbUrjHNEIG9t/YdpTLJ7xxD64XVSLC0UTwHA4pd3t6wgyREcnpAcqQfZ1gTddShRh3nde/H6
BRJC96LLkxBmjZAT4rTybi+6nA1+O4Iz37JrPv24MORCR3KXPw5lBcbQKlRfaiYgr9xab3MAkoFc
XhHApCttG2uemGSxk8Thyd7DKSipfnbtbhY4Xi3am0Fi84sESCzPRatj20FsCIZoDj8258nI75q0
f8iXypDikBrrk0PKA4bHBnQEdycvCa1D+awrlmbYU9lDjI5V9aP/A2nPa7oh84Ss1FdzBAfKAbFi
elCVRmdcVamV3yDko1ocMxmGFNt4pFSBHNyToXH/JXpHqMNJG2dUyFcUsIOrfjLPiKA7CEnvV7jd
NWGTDebNZ+XXcgc+XQ6QnP2qR0IVd5A0l6b9V0KGp+ZQKuXXiifmisivSzp2ag3lsYGsExT0X0F6
Dt4uxBOzUxBrzJYbVa2hqYbgzoC9qUdRo9PyiKvt8kdCEzRNRME3j0NfaqfEtcpGWe+UYvfA9zcu
4NajTqZwwrb5eLvOEW505vmRoqsatm0Sa/Ru0fLfYbmPVXGhyxEkO0C/Ow65ZqhIAdykHYN8hOfU
4/HjGaUAsw1wJK8Vm92C4Q/zmhy/ChCkjknFaYOl8KTJjLT9Fe8Gdu2mBfdl0TO+GzskatdrlboY
IFVbzo+hD/cJzgA5+5xIHOpzQw0cSUM5JVwRgPq1ZnDbJYs55oZ5Z5GI64QTft4Y8m2LIlZgLNcG
CsMNWiS7sRdgxHPY66U8fDG73RyqAJJI/fY2pPGx2aB1qt+FV7xFrWsZTcl6FQP+yoLm45HvLF6P
lLL95a28p2RwfvCKZC+qAvG/4rL/2eD39vHuJdJuGVv0WEpnvNq8veVnoApdYvZO6jppm5jM+uB5
cWJcOF0omCMwa0QCs3W6900Y46hFPyYyDia+SbbJY9ZwnJQSian1eB+ScomVv8ENOfgGQqPEo8Tx
oXauOCyLB5kba5FD3FKCMi236VMy8jVOfscIB2pLxG1kLooTNXig8GtFx5y5zgfUVo7KC9i2Yrav
BlaTed5JoWIf9ZdrgUE60WJ55aaGwB+sLhyVQhi27lBsuKV8sXw8HAGu4UWhIgBoctvl7HTPhW0X
HA/dxyUn1GFi8oXO2jAk/9a8/5XqnC4rqblmJeVTLXaD0/cIxdcAryDf9vDn9pkYME4TLJ2qyxHn
13Jr+TmgkzY3iEEj5E/wwsaynMC7cSfWf5nNP7wCqg9+uG59ecAuEYI0EYL8Q5pD2Z1ppPy8rIYS
2jK3HIMDLJy2V3AlmyZHsq6dc56mWKdZmmM8CjZYIbsordAOL2unii5lpti33lBFIfB6VR1Ridop
65u+VIhX5qpX7h5KFPpvjmJbr1bN2jvDGjAUQ4MHStkW50crWmzVqUBH9iTnF1ZT751L/3CdcbsE
szBCI0ipB13LSx6kZa+jEt8Fgj4l5rtZ6uanMrdYUF0pF2xF4TlERBLqj28Un44D5qOXICYHH+FM
u6dqpwF+uWOAS4qAKXeFeJ56KFCC4qNV9moVcCPxs41kcOKM8eWnQ/gzLuxxU1J+Ht5ixiC8HgA3
tWJEjtiLxYRBCl6b0MYtJlm2BaH5Hl5WaKxQSqtwMkMy8o0iJXyMmJUc114oW1iBC/SnkAVZ/FBI
L2y/PQTQlp4CfcdrYLuvkGgbuxUsUmVoDpuxN9NKNzE3lGmc8XQCnFBiGs79IXzzw3jxAqeQdJqe
M57KQIGFKUFRV4t+W4IwQIspTN/aSluouZd+ZtGDk+Z+zUPMNS3gv6ErHxjHzSyvuBp0JeED36ms
4CzHfApdDOC69CUesJtAF4RnAc1L8v742Wkp7cWJXzJ6aE39jXf7YstdTMl6rtAunu89ugHteCxa
k0C6sVjmECkfEJwM+2axR0ZEs/u7fTbCGMq2bEGXSro810fh8439zXkggrshb+FbtUDHdufoPidF
lka7tQ0iMX9/vIVXm46/ugQBRE4Pr/nOT+f9RBKJMECJtte7JkSYwqvAczpiUGZqBWEZUkVRIYWx
ts4y5NBsoP9ZhFcwPlwpr2yzlXIAwB5UCWtyUMYW4BvV1CGOw+ejJ53a6jzVNJW0A8X00XuxeToo
mP5xDS5AUPXBiIsu6LvJSMKB1yR8LwXax+SnOUPwNKqdSJtnspyiknmAz3BoxL8vLW+/CTBV2ggV
CjeF5rAVOMjwR0Z3vn4uI6xEMoilmZOHG543hwo1b+IH9cuJ7nr2Gp3/iYTZUO3gAx4dDfCNKyIs
QvzRaRjmqFBsWewi9lja64KzinuqJTW/pg4Cx+2GeiKhVGHCkXIdrhoMMj6tFZfbcQ8WJFmdFXOg
CTdtb/ZKbPZOP5DDAkHx4HrAM39e/AQ1upY7Vln/4u47yoRVaqp/pH5aCP41mi6ZJMS9XREGaQMC
nkcs0raVR1w3x6mj7KrF/MNjMu7q/ufCNQF27PkTw5RxYgCLhLpnkdYuxKFaJvwrvHf7joOFlimZ
D+TQuLNrI+wavcrUYFaHL/Xwupp0tYEAhEPZcYBGj0NIFNsNrImjd/3eD2lXjTx5PUsbW/OBGZ7A
s8368IOYlpflYGW8wsBv/W21jperx5nhKAdsHZgLkdPNIjYwgUkU08RLTr743nxkqp/HDqPtdw9G
xx3G1k+Mm3XE9jQkQImh3KQvVUSkvxJAN0W0sbo3/8FFnmMKgEA02+3r7aydt6tLtIG3sNBr2QYW
jErosdhVnaAkqPhqeqv2Yqr6jyVaAvdoSmb+bQhhlpzUMrfNdEXtPt+lPocfWy6qhG61h8pZEZUr
6BptLrgGPaBwOHUnCOOtm0K0+Yz/tLgSe6+BfWuVv40bIXOHgy8RuJO3SBguQOMrncdAUlWN8xX8
jGQR73ZEzHn71kMlPZgJ31niXdMGlkEfO4fcJCqSDCq7D7UMA27fBbU3qaLNjf/HPU1xm74OnHfT
AsgNFf8C8EtlDxAqw353S8og3LpXokQtyn25uLPEqXoVoBK3euwmNrtVKTilTzetFZPDSPihMf/j
oWuZvq2hynEFbwRtDwBpscy4zV1dfdapbrjFs4i2AHacANDrsQr1CUnYCkvwW1ZH6p/IHSlAPnqA
sntzbqdlbarQEB8w7sT545rA91lsIa9ilG9ooViyZf6RzNgli3vWHJt7ZH8mMBAovoXSLSXyYBOW
Wc1/kWCEhxdhT9QtfHxWrxezXMAXNSkuj2V3nkWVn4hDbmua/wFj8AA7ocJF+DRM0u1GahK22iYp
GVuz3D+2+ggaWmZscOLdCvwA4WYBcwPFrUwiYN619MBfjsojH8q6uAys4Mk642JHq/RPCv9yvcWx
Ona+WYodhWSWw1IVe8yTDkWyt3WD+MudAUpiALxvpVdfx/5ngkj9XolOdRGXdoYoDbFobeE6TIWD
wgjbyc13g5dIixfMA1yQ/Xy6qgKB0bBeiz7lVujIi/apfL8J+j616GEQY6/Bo6wSOU7AU4SmCm6X
oqW3tlcNsmHVkPJMRV6qR3wdVel32Kxz9R95JQo33OBk/Z0eA4PClU6xbm30JdP1ghOjrrrmB82u
x61tsRbn5t99DN/H6PlEa4veHOb+AVNxfk5BQAh0qjuQCeoNIvVeLM/E003dfVA3dG1bXXB1QxL/
z3Yu2bjXRVGU31j1ZZL2cBsQbpzNpDcjBFIW/ukfjzvSGFy76gOo7ZxC6aRKIVj3HZ/5InZTU9xb
lETsaZGjicUZhesi0y4iKG84wUYJc4Ujs+rCKkDSYOHb2jh+QWIej7alGNkDZEC2D7LnAYGHFUGu
rKm82r2DLodVtaF7ZAT78SIQC8ikPUtLD2I3x1+eOyxw6RRIcgiycpUzr9p2Vsqn13/9Fqfq/LLN
K4IgSR8DmHo4bLfOk5ukRb30ErwhwZ/mdjddHcJ/qqk1J/EFq0V6RYAJNp6xALAFq2VovWOvVKk0
nx7MBo20TaknMiG+oGXGBxnIveu1J7w3SW4v3KSvCHk0KjhDF0pNnF9oALHhb0NEvoP1cyzX2pZt
TR6A7a3qlw7nUKyji3W6JX8KuU1SR6MPm3c09ntjUmYkb+LzEIpTY/YeVFBVTbE6zZumJqZmsOVw
53z8mHqjp8iyi40qO3R+BjpGUrEaijkOam2w1vTyhhQkes51fyrT7ru0Gcw+AOca9I06L7Ao0G/9
/QJnrBT3lf48+wQI80baeTdMb45Rzxenq/Ige9Hp26ujaq6EFluYPhsNiNvsxvh03RNFlxyQFzEu
BfRI6twwl4/BWxCnWZzGnglQq2qpJ+WJESw3ijg7N7fMl5n9pJ4/a1Rc7qASnxhC7kOt7eRRUqBu
QN/Sum3OZ9zWyCIJw466rBdFGLDdYfpmwvAXkzjy4PsEmrteUK4mzn5uY28AUnOnp46Bq3fPmK7N
znTnmSS1H1EMldQaef3ewKgPbEByVgD9mSfk3PUfWr3Dg83GTZ9AKQFQvAqFXsFN6gU+r4pCXrO5
xAjw47SwNYTtWtRlEVkPabegGGn+OWvKlX05jtXIsAAhhIdzR3C4SWy9DkKPB+F+eRTj1jSfJesv
6idEl80abOqqlH0i0EbWRGn6piCt9vTCW7iwP1H620IqfzcHHIfZVHCstHew1PjawpChMshnEAMb
KAqXEdmGA8kxYDgA44U4csVgixqNsk8NySM2/osqTgAS834rKczpnkB+JQhLwhUePjOjlPcMaPbT
gOsXh5HU55S0A0VT1pe3Huyoo268oybsvMM72Gku/PSzWgIWaqLxa5bdVkWdp33EoG3n23VtwcKK
EzzbSsYb0ppz1glC79CEmzyWN1nfznMSwh/VLlH3Ff6PeFyFedwUOsMLuPkZLm9C95b2pf0RC4sC
Lw3Vm7UvUpCXy+9yaRr9iINxe0HtiLOp9fIlEIxkxQhXcQK5MEGhy17SnncP7XFqZGu5EaSfnyBg
xKG7StGkph6kgD8le/9069csyUP8GdZsTuLAj5NsOpDoQvRbsBm8tSADk2NMfHp6nS5szJaDFzeD
h1Xyg4J6he/UAAdCx0ANJ5dsgnmW7+EW6KFzm4JDFv+MEBtKnbmGOCypzcdiSMEIA3nbCB+zoKkO
OpWiAfTRumh+TM7rTEEOaOcC+J9K0d1FRrFUHmD0EU+bDcC5+qx1PhbEGi261C4KjzWVQ58iIWTE
B+79CKW1gMhTWsKxJ1r5xJ4QFfuXNgMKsuCFqFTP7rYFH0y3SKAJNzCPQSkgbWE5QJJ1ZemL+epu
2Y+HfwR++TujkO8c/qjR/JnPOUmTrhaE0ZkhYup65L9f2CMgXgCO/h/cGH1i8Q/F3S6o2fwrr9NS
fplEytc9uyKZUi3qnsMuF6+0hx9+h5mBmWuvXLRIGAz+2+fgrmVClr3le2+8LTzEpfeYxM2tguSs
YNgXylg3jPE+7W7BcFx0jo6L+38q5yNM9bMOTvA3w6M/l/3oAGSINBlk+YtEVYaQBPCuNCpAzMVL
v1a3ljhp4rDrX4s3RTT9xYGqernNRYY2RMghyvRbHCaFiWvSsMN09rzniqRFY+ADlr0vW6kh5DYJ
HkWEWTW9Zf8fvZ0XOxDGiLG+sdavj5+mfHQnVPnnhUIKIU3J+AJUbPaxEV3qNgKyiBfU+REgUaal
N7JJ7T29fc7JsYQTXC65zgeaAKQjH4ep1Ff9dyOaU1+EB6QjR4HkGYdJfhKRLcOJqKJYyA13t6H1
89l3dGw422krqveNwr2YqMTIGhHeOr1fS0e555rvoshWK0DNYB5wXrb4CPPYhU2xkdhizZ1EwbWs
WI5g4g7xdOLtc/BPiztodJJoAGOQhe5Gt03ysnPNXvraU+Gr4hx8TxANZdHPkcZTkTszPPSIRRUK
GVHk1mxTIlZzSeDuqn9yqeHU/bTVq0FmQwpOdzmHhurEiv0V/AjblHgWZ2vf97TkzMNqS0YOcMVC
qMbEo6/DibrKhe3HRfjM8oHxGS38NjZXVB+J47ZO1OnJhvjbwATjPjb6vC3DOBEGdSlxhuq1hSkx
r/7fxbFtMCt9DtKviWT2iMsSj7JbNdh5AIn+nPj9aPUU+ZR0x2rX+N6XZGCmW0MqVzpz8Pntvfxb
E+IlPLKkMKww1f3r1dZfRxMS9eQiEbPbtpnE6Lejgiwjb6qhbVfeK49jK9bBZrb0tVrzFTOLqL/Q
FisnInZ0fzBulfxgfhnO6H5XXuEWe2ttHI9y+PxsCNK/13IIPPuJw1ZJ63YgxYYVZqibUFpgFVli
nCDi7Ai7ZSe9T1k9vQucj6/EyzaFl+wjJWdl/ghRsZGEhmOhznx2j6//Mersr3nZl3Nr5RTCeDxv
f7goUgTzyIBPj0BmsLh1hVcPmQbJuTVcHO8qa7FfLfef4I/33dpLFZ0BpaLx5i5Vzu1T4EPj8wg0
RTKOVqIwckmrV++gRe7Iq5jXKZrdgyIVOaUKBzbHGyYuyEMAicnBq4/wuRm0ZHvE2S1RXazwlxj9
7MeyN/xVXNBhDk5LGYsS+dZ4jIlZ6DnfiSRAcKmI5181tEWoLcsZmlvxzXzdsQIzFjUEY3sxtHXq
BhriiU6Jx+sO7Ux3GJyuDX7vevVxn6zGAfGOlaZ7F8On9X3GLZP1zbAeUfj9pvrGxA9NdZT6otX0
sTwoohH7B8dBOKPPJ9uYAigf92KjCIlTLQeeTlkjhyTPoFRRcIlczXJEMfgQ8b/xbkNCRrn8SJE3
DbvuaZU+qJyx/8hBqMK0K5vvj5knQy3hE+vf7X95uYg6PZgG5iZKmzE/N2RTt0Ziu8gXiX4vDAzQ
lFVFWP2oDrV9MEcvBNHoJ4RRkn3sffoTW9xkij/Rpkh7kLtO/O0Sefsp92gTflPvxmbg/CHJrkjs
FpVyvRLVqdR0+fGYXrKAcVi8lHB9Oe2QPm2UzG4AvoTVkKeONlLgz0NZ8fDnammeNV2Ajf1v0e0+
+RPqZbjCDMVEPu9F6LezV4c0Nvi5Vq0lLAkBRfOsWtfVfc1V6MqNZ+yNSTqxjremiwoxiEC8BReT
4DXKevo4uTDDIrVsYQ91BWtf2Ol/FzAdjwtCGpkpgzIeibjK/04dhKGRVe6M0wFvrbIpkOrQ4DLk
g+zTePKYsj35brr1h4sGUS2PAnRxHH6sxfcgyo7wjpqM+07JzoNtNJmqVgsmBAeuuCZpCQtJQ3uU
2zEaZGWnD97hrjOAfc+S9mahbsVRokaWCu+Ak+KDRt/ZCHxIXdIiZHck/OXW+F7NF712gl+s8LIy
ksomh22zQCUICtaJVwMGNAD5wwqCn5aLt0+RfAVlFuLFTLna+1JzG9bDCJCpHFwm82MimnA/fEhi
1fFYaxVZqY87uyjoeRkPrSdktWRYeB7pC1nK/BT0ceDJk+nSI5GUurPAKmF8gWIise43PQ7Cz3tA
nAOR+HxdXoHO3r2U+37frNsZY4+ythzevp5NTTYOi3pdSYxyYjkBXR3rjX/DRBLeyytr+w31X8kC
AeWr3opiV132dnzPLUpbUODXY0/g31AnxViA2NrP/W4GwryZmrehRS/c52yDGAnaZuwS3pkTMS5E
ThDzbqALJGfXDNxDKWKfLCYDO8R4QnleJwEYR+OQtynB+y8g7bk0ioJ2edA/m29A5LVIcPKQzFtz
AJ2zN9o286LeXI72n094mwNwPdeMtRHT7GtwUy/k486LDVjDdnHATPoAWlIQhFSs3tmr7E42FpgY
wTOvXg9LvbiudPN1wU8eKs9varo2ii4KhukyBcffUHRRnMD5smquU2jZlIJ0go5qZF/fGOZlzlRh
N2lCXrBVHMhfjLAW9TSD2Gk6hBG+XKo1hReZ+L7EFlz7ON8KTqrUFwEM+MUzAIskLDIlRdVun3sn
7OPuN4Zo7JflKbZ4NqY7/bgFEc4C9ArHAsKt85QyXz5L9n0RIJM8FRtcgrGrY4amaEBjFP3GhM6Y
ir0sfKMZNGo1GOH520UXUNCNE+Z/I4CPYNsdzPuBcBBtn/MuxcDOmQlPtu9GgkaBs3k327uz4H5z
1+Cdm6evT6Qutrknu/i66tqa4XjsTfbVaF+jxo99LnzeadP4fVnpoLDy80PEJF4nsrfz94I5SXul
54M1DHzw/++if6DhHfpq/szcHEOv7fJvlRKMiHp7otqnZu2RV1Dj3COmiqVxnb1ubDx7xIxpBz+5
tNO6i2Uok8l00q5069/bGpjV9wEaaLpYtFHyKhhUJnxftIba9mEk/Y1r4FDxjtJ5ZDuL8Byfadfx
FHG8dPLvvCinxVHVtWRlIa1K3FDsuTnYqZS9xf10T9t+n86dRXHUI+/L1JYcli5VrwaTX57SoNcl
4Wc12w3KwbfQxeG+NOYhcXO4SwC/5eVj1POug3DM/yoEDBRqZwUudYqucEqRbwITIyAM38jgV2qx
xZJMaXiX35Vz9sEzywgqvgos8EwI+U19KFNwy3buqW121eGMSw9MaJXIGzngPvcPS9Exe1MqsORR
DDSkDFUf7/po6psbw2Y7DFGQUyUZm3lSA+05Cr/6iCQbkXr6DC7fJnqTtlRhXeIQKNSVT2ShvjA9
BB+y+/9qPNF8as+6FjUHOwJosAJjWYtnsS2LUXA0F7eY4fUn3G8Qyu/EuvlOSwOrizJsXHMlkp4E
VHn8+lEYByHVyYtoVG+64h77HLJUACyREGByyRFrh1bgeZvN3NJKZs5bxI2J1jxxbSz5y7xxLl4+
GNYQqm5vHUDBIX/6XSd4mgJS9FSAeuvkXuz1mJT/qRqQmI7uH+TO636O7AnLJb0O6tukfgVTcqZC
oolT5ioPnyorMXRiFUxn3Y70ktUPv20Q0BJOcQ+QUmy8/TivRBlgDouHXcEi/pIOp0CVyTSeVZqP
hMDvs+XLN92tGJQ/ImrJebkF2vbIS2K0KdKL6FhqQqCOhd2Xu91lFePaLLgmCESpdyJWkG4WYBy9
3OlWv0Jc+PpHrc6ygU2NttwpkVKWxoOpzXL10ebuHOo37LigyRBnWSXZOheerhu8wExESYq8kN8F
nAFIPWmzJPiEySoJmCzNjZSItWWXsuyIVRKash2Zwd5lpiU4LeS5F6xLAosZEStbmyUhSbinywZX
vBibSox33/icjJDQF5M3TSaFDP8mqtetuc68cNBIiN+LHgiWFgHA5THWK91PGZ5pERBNaRR8acIK
5TIWE4fdPrnNG5Iz1mro6CTyyQ5e8mggFKdGn/rQqycQRwt+LNTQ1yZrkWcDv/xJm7Os6ThHQExn
F60M+la4XAIpQgbIQsKBrZMSFmG24aXLRCqY7ejWHVlz2lYdC8xeHotLIrbL3g3OxHRpAAAs0/Pr
FQzygNLvh7qapTNfG+wSCzE57waJQlWlk9Js+YHoEaDlvcKiVPIQMAZzeS27nrvUkeCfIyNmVVZe
tyc3M59p7GH84r2AaGIDV4X1hsRMnnjrlSzZ64AQegqBPMukz7N1kFqVazdZw53BlQfRAuBfFDMC
Y/20QgYjegdu3yP+Z3lzgF0Gn8mIhqtneSQxEkFAAomMODPxWsvH9eiCZ2PYqNrKGOBt6Eg4p7Sm
mUGQ1/c9N9D2zEuI9V4nbKRpfIuBmZ1L6nLOsqhOczSqupbgTzQmWtHIxRVnRX0ZlgTvgTijQx8s
Yl8eXej0GV8bd6MkUiHyU6BZB4MEWtJ2Ie80lVov0IRc3LiigBw3mM0YzNgVrxWaQje0+9HoTxPN
JWWxGmXFQ0smAgIZg8aE9Ft5KqVgir3qqOIZl2I6C31hpUMR1TYcq40NURRwh0d4h8bo7XvXZYPW
7ZYLVmpE5IvD0A2u++cQXESMvhsDMCF8XprDsrnFltKHH7Sz7FPuAoLviB+MkAecRWAsFTWLumS0
s8W7sPIHc9cUsw/4YR2Qf88GaLiYe3Y99SwrFyjgvLuq1ZBYc5E9UneGphK4xIrVKb0NxH4LdnUz
+XNYDDYrXn3gS7323pifNFCl5jss67IfZk3YZqMhJn9TwVGMR50uvYtoXYSRSa/VVq9VsIcjNU2j
Jv+9jbPDP379KSY7o2C0xeuP8XAWVeE5PFcDIXAeXVv+UYjd/Jo1Zy23T8yICeSq/F2RDZ2HH4z8
F/t0SY2tmfSFjRqCau9diwwwxBnQvJLQBEBCFy/I8hAclzQJozAq7wGLfpaNKS3Diro7bRSQLP0r
R8VfXjreGK8vH0iUkDvzXZt/w2A6x9FZKWJ+PGpvSfgmym8T+R/xAEK6WJFj5MNdzAU6rx/FDy/3
LqJCE4V1pZUeS8KzH1ehxzyVhG53qdx0oj77fx9f/wG7A3mBN2SjiSeWGlD/Q1TJR0t+SIHuRU50
5ExUJLjnt/sBiMBSmdqxZX793jENuV+sCUy8JaF3PbxW7zarknrEvd+rZMlg3k5NVCN1gNsKVvHR
YZI4flODTL90fRDHYLoFopOiormiBxmzrbs2qE64ZWzvG4kE+oITN6BiT4Cr0ZKqbS+rQ0/jHLQc
gLj6q8tuowXGNidJf2TS0MVQeWs1k0MUlFrwpJDisKBJCwwYYouN8TlCLPbqIVMYmcsvb7qrmhgt
+e8qVMO+zI862i572ctClmYGR7U/w+5urVCPOINeKEG9Cn5ejhgvIknZgUA41U5lrcou/DeeQfNi
g+QnrKSsZWRVKvhXT6apc/mCe585laiMndVDXb0i/td6geoZPudUy6of8KWDm8v8U9V+9BM0fM6K
Z+v9QNZ0Ta8qA73H8U8Zbi371uTb73P85uE775gPs/Jfga065BMQz0krG+M2olGOxqng68jc6zux
pIImY6jw4U9/46dogzsYZ/e4HoBZQJLqlqxU3Cupz6SZbooMnuEBMkdWz8a6+3uPBQhn5cSx6oLb
hTXdEyUT9mFftHjbAy91DzGql9NAVS+MuDdmBUD9zDsylb6TvgwXub6Ae7+c5Ft1gIoZEYHjcXSi
uhKITxHd5IR2W2ZMe7LHsuYtZGF61mFxK7i0Xclt3/g8KoMm19FTeRI1rGlJtOEhvEMplyHfmL3N
dgq0umekWdP6Xi5TzTMavreJAxLuaRf7354b8eumxHy2zM8eMyNe0hsucT+5PpNhxCxEBTv6ggfz
Dekwi/I3Ar6LNYauRCqAf3G3yGKUxV8yH4uF+0aMZZuTOfKCLFkjb9Yo0zPhcbIFLGZvU2+BGfTa
eDOJSMGzIld3hwLBgnpuh19X/U2s2e1am4sVFHmYBFoPZ0noY3U0JNgpYBicE2bqJzdlkXohDMZa
jr6P+NYC1gwPtJwkXs0chMCt94cmOxG87NOY6EM+voiqmUTX5y2Vg+fNucN7qhnYu07sXtjjupJP
lHwHZX6B/JveZkrIdlOhfOrWgOafJ90d+t2fXwXIkp3JRKD4iDH3CX6PFLdwb4uTDV28l8/XkKTo
b+p14fWoq5S4Xb2CWgg3DMQQwNjN19CNjsz5KGZOcQnnlo7oyK7MN+CM4Oa+iYHPfWfVB3vji64W
Hab7aKkcdO6Vnx/TtgRxWeyBDgjP6FrlyVSb4KTAF8OXKNH6Lqml3oyx+ZKb8XNP6H37rjgTrMbN
cXilXW0UssLkp+4PkdOrRCbEkVlmDZs2RKq71OnanX+0x7iPbqOzSdm7Zp73ufTRckN082UO9c/A
V0ZV2Aa9iTQg8PUSLM98yYXPyD4IgqVoVExnPPRzlCiQwpoYAp0/AXRDb44z8BpGxp881Ooch2AP
BKVTNRbYjcHqOoIropjpSHMTONYit2PqaOt5WTsFOxtAU+CAS/xdjUSJ88TVo+vtNGKHx6vIr+U+
XP7Q1wOPSYndPGR2B1hu0h8M7WFk0/zYRE6+EHH7nZzUSDLTq7YWduxoFpq/zmP9Pomu/qhZma6O
lzdKXeH/CTFYob1UidiOFKea48FracPUcmIBHcWCYpFVdY9wbCZVRMu+hFvQHRJ/KBMAjSKsMRqA
Q2Ob9CU/PKfhltlFS9pZrgp10SjBZbFp7eS8jd8lqhGGKMrwCvfIFUXadidNvLSHQiMQEQeccFjZ
92Tc7G4ovsAZh3plpL3/Eaw0C3nZUmxhR92ENgZ7Aw2Vwe+RTymdlUo8VewjXLkYPjWltg5+GDaJ
gWUnxGquI65L9CtRguZCW4d2vG8YSQumMeLzxpNP/grouBYyqCmFCWlBG9oxeNrxjgEKsmWUVU2s
UvQPKefPr8T00QC92cHq3AREJXFq9hXm6t+LLN1CO0cT0MVdJ0dMde7+QyubREeg07dnuXfgEIpM
hY7wa8/s107GgvmoZ2cjgRtS3fz+iysgVnrKdNG3CE4WXindR9MwJlXcabYLtI4MiNbujEYHkJmS
Aj97ZVkFwUc5sIHkRIjCKPq/X02g9fPKrc/A8HX18xDhjs6nrT6SKzsCE5rAd2t6YEUeQVvHlPV+
EMW8DccOY4VAn1NieEz2ARTYkdiXnYKSNErRgBAgKCIy5q2Po4gdB+99XfHBDYyVA8Gih7w69B+4
SmzvHUaR9Ifqa2WhrO0essAER4cSOe5WIqD3FqTWWMM6PR3GUgvX4cr3PjfO183kXOG229bbRGUb
Duy+gbjYCRm+aLXf2hyJ95vE82Crh6TwxEfdoNsToO56aGAmKqABNCOHgopQ/PSIpyt9ssH/6dbU
6qLZ3+/VxQtl1hDK9tRkRSZSOjj+9sRe0qCoZfHrRzo0WXLWUJb7nqyYvYrYyU+zt7XoovjFvtW3
rT8NkjC5tH1C2hWUQQGecCDXXTNWaN5VIWiLKnGGZN6i7FXYqTpq29CxMxLOaZdDgoWJn3ThcmrB
yrvmAt24V0oa8Z7lXRaiCc+VTATqZHrafF7aUbGdAkmAXXMbibRvzB7nt4L+cc83no7U8hps1hiJ
WqhQMWM0GD1O1Vpa4jWQcxk+IfYCkqb33+sDSBm8MPqYHEucnDEZqjWWHcrvlMGH9fDAbTUfC6dO
jBbfcprN+PlkGFVdkaRA/7GCyFo2RLcjl/HGFwNPNc10DDzYsiFZDzo0trd2kex1jERk9eQ321Fs
GI9LsjlMZUMguWEe/UR+FYhLhX2olJ5DUCRStgNw0CUxPzoj/uNYtX557utr40e7C7cl+WBX+N7R
ew4+hSfGqEEgIRc2VX2lhJ57YDgYr3clgGAlJbhPtqlYjjbS7OK28RqJR6/ZnVuAEijm24QZRM2y
HK/X3aMw8w51oC/0ihcaaducBiMl06EPxDKVW3grrc8S+zV/BA9hLrJV/0RG6gl0tSaO3uMFT0he
IsqdTk1zlsiXytABZ5B0jF+LFldyxhECjixog+JpCEMWrMOfMQp/TSgeVrfhLMqFCwuSsqPmF3Lu
toHt2KBeRHRJ16+V/JRxFw5gkxhsLJoKpIqDA2uBEKNyw7DuX8Wl5z+HUlTC/1+XQYpuPAuKAb6v
QvFhOVD30/4KwXpOsSSsVVZMoqY8adhQxxCWGcorzQzZkSahMp0l81jhVQO2d3/+tWIYhw93GA+S
J2bJVfU4L7w+L/wADPLKINnxanep4UrZdMGGuObg6Gp0/bp5bCFMViLKwX53N3DljWOUOBom2PH1
LVev29Er/ixn54EwJYeivvVkFD+MZTlOtOfdD7AG3WYYbaHCHHi95L+qqzlZn1AOUKGWb0SgFwgE
oAGiLVTZ7xJxNEy8hxyN3IR6W+zK5NaaAO0wQCdFpc19Cs0BNGuxXPodC+ccliHHxU9LTi8JLejn
6mJB/IQ+aRB9qVr+XAtldVfKva+rkc1Cxnl2ZwXFoqdkyHglxcbpnPuNL+tAjpQZFabLQT/BF+WV
0Xi4cDSLW3OIgNgfXb62C2K7fYefDRW8uH6rPpZpGcisKNQFdS3ZpK+GZWIcwXuDrvLJiwmR3bQs
xkhCIUpsGOjjDlUvj7xNV7fiALZXCLE/WuOas8OZg52eQTNQPFS1pd+pN/XTEb3GoDA8cIuHqjnZ
+I4nirmvwRhGPtFe8xeb96mIciOYntn8p+89ajWLRXWVXQT1BoH3lDJ6UYB7Dsx0HzkpC3MoTyB8
cQch8Qc4/ndX4Z667onxEn4lrTPOvE83HxQUkHNXBU+PzHHuvwec66mcOjtLp5eIUOA5BtjbAx6a
I8THw8SaMOqO2fIhf8B5GGPTmiSI332b7HLBv+oUzQMOZ/CoZtADOqXaG8nxWjknGzxzGD2HmcLC
MnDQskP2nJ7OmF0vY36e3O8Ml/8N3x0TJqQryrm0E6DjAmj6YlXvpmtBdoruGPjYjhNwl5tEmeGJ
XkVdIXh4/8YKT/X7SfTTRP9CxT6bxYfq0V1Crq0Eqs1GJeQ6IYbu78lSNUUnFLxMUevUdrGcb/hB
H71i0VVNg7/n3mShOLIsjWPzISCITv4a8IXEMEjhrY2UJarkylBfuCmybUDE7GttS9JZE6xBmz5i
UprWufuOMS+jyuSH5JeEqfqkmnN2BnmraRapA6jJIaRMvWZ6AwJ3PZWA9LC4peFJh1HadJdtcTN2
rkQVcGkb0uV2CkR2mZcMqT/usnp7m+C4KyPqkmHKgF9QuLi7uOloup+TObbeqUOoqEhSb+UujP4/
lyR2Zn8rQRC2lIJUnmavRCmmolpNHiUljhQoeOnHyI2YqMAHPoaxcPnR4qAkah2vDbBRSCXy4jBi
7QiY9FZYW7c/h77FLSYRXCmuFVuMGuLyVEG4wzBNxcLZq9vWH6dExQghsv+jKzz0gnpP583yaTAF
MNz22xGcjIJGfsP4wF72D6kdA6NdZQnkJDqXZygAcx8np+sZRxpg9/2u9b27PBgynejScarhK5uH
Nu9tmIJ4k7lmN7SPPmc+LFD7qe1IZhN7WfgJelcksCySGI9dc9tXnB7oupeq7JS/tLSsGVg+0cPY
P2BQJJbBGcQxJ9/HeAXAFr6WSEvrphFifYEVyzLwY271S0c4DjKaXgi0SAqV2Rs4sPIOzxKTKvAq
ZkfiRXVswLbf7vbFEoqKCzMaC8ohEN3+SR5OwvvF11K/85J9a5Bd9hemtrVtu1LEegFriGYuaonE
eN2AtnMpy4kELgsIXYc5ebVki6/2jb+DDBzWNbKswdRO/Cozn4nIjPDuHyNDRtkc21q7Co6UYlQY
v01l0+OPdv8lcnaCQiIDIX4sJOxb42ZQP4zhg0g4RXapZvtLauG8FlyV/zcAw3WqP4CNYLxra/nd
JCvChiY+HaGf+gxaomKcUIUAgfWPL/zmiOTEWI0imwwGwhGpeiZWjARJX2NUELr1x9VcfekU3Dmd
z3M81YNhh5DPw+lsTKNOa6GTDLYzwMoELoWDK96I+UTkFLYc3DUlAPjT7ARwS2ntBtn7I3Pj58dS
9rgqk+BPuw93yVHf+mUVhck9CMPdOkDlqsntCrvNqoLWO89f0wq7WggYMVvTSfspwIMoDv4DQ7BM
GOqx7slhq2KEZtuWkOUwT1H3fENzLW/aNgQ0bu8LFlukSBeZj9AXFANIlAaC3vuL/SdB5Q2vGNUC
14iA8BhPfcEoSGTuKs77joTJkxPksvXI7fpzHCJHZ3rnLbGAnDzC2eyh9MNZRsvmbPVhXTxLVY0U
R/2dC9OD8Uux7uLJ8Vlhx3eeIsEwkMtiqMLVgkr+/ULDsDEeinWVfZ3zKZTk9opkVZBRMbw2zyJi
EVTGiRDzP9XMb6iC/iciC+CoDFr3LWvDGXa09nycDQVLLCobHaBb/9AH4C5CUncra2kcfipJu7/R
EkMbNZf9AMkgpFDwGd0Y6hN8i3IG91X69/1QHB29uEUNKPnEuDuq1uIh6oVHdEpX01cQFICw0nz5
4CvRdCk6ZQANeewyiQEty9zl+2/j0rFNukS1tp1dPX9kiz7AUvZiC5/Q50XXj5R9HHi7qZ0qebJL
EAhfSmOu8u7LtzaMLxHPmCsUACOkBBwagjpOuyH/i7JoHpRAkFTdVWeM4vIuuoYr+d6z/LRJDGzq
Bp30jPemAyyNafxkVRj/VyHuGCBVB4ydXKW+9P9IbjrIwU5yayhr/MMZ7abNh+DfEGwIymnGAHa2
zzTMS5bIN8Le9Wb7hYYOnR8L/LHT7JXRD0f7bgGO3G8OYo4fUrQ781RJurumK1bz8hL8GunJ9Geo
DtWWk9OXqren+0gN56Jg0Un6t8jkP4+sTb/HVtmkMQLrgVh3HVKkEMdlVrvvSXE+hMkO7aNtalHr
i+h3NPpdKhVZ9t+ChFoaPgE1hs2NxLL9dkgwv1A+hbAuOSED4goMCx5sPdp4IPeFonXjdQrw3JhO
h2xHGT5aEYqwewL/4i1ImVE/lXwYkBjNpTn7/T/Cp1W56mM7nPJLyXyucpGOkoqp+oHUBw5V0P0Z
/mazSr+1qnVHeZypbyUoLHDBqA+flvysdebC9t5kMeBxLdbF6XRqizzvfa2mOK2CjfZBBG9rmEkC
qGcsjTppHCKZwRWqlrG/vGr+Pmipd/LRfWT6SNBjicOarWyH5WWBoGvSFa5avot9K8CsicyhMXtn
WqHKnkKox0zniqRIpm7L8t5U/O9ZGpLQ/LFyFTOxnSlYb4mWLlOzZh+4V2wkRzC6lZ6s1FFruhAK
mHw5fMLUE2j5JkUlMIfzdJ7ePB/X20u1XF/OPKRm+89sO0mlRWjdM36X2TFstdSke82/O4cyId6v
H4LFMemEtbf6qqqyr7fAN3ZM+NUTNSTtzt6ktXfMI/nf/UmrXd8SG+BQcNEdO7ma1JQEMlu642Vp
IvFtn/pmZoD6PUr1gRHlthyBu9bWIhf57mR18YYR+8unrrWaR+ODWE9HYqa3iq5QXbZjgECpJBAS
yewFVUnHN6gqk/giUl7canrqf1xx72u+TtTlo4+S0ePDsZM2gZQY6CMaqAw0SSL2fuOQt7TTFDP/
JZ9YcLLBghpaJ3Nn+7ed3IEIAjVsFxLUsG6cTzb43cirQjjWqaSMbGOwKkB1LPQIZBBGzH7dXYLY
sqzXQNhXqaBJjEPME7zD0L3ozu/vL6qGBOC4x5qvIPmOK9I7pNdmRiiwC6nMQIZHk+C6Lm+3kWoP
nEQmiDNLPwFE0+gm+y/n6Xd6ObTweC6OctCMbtfvVz0bwhV1hLdeEP6A0lLgtdfMO4yTuelXXltC
6I5zPTUKN6bQ/horR6KeamLYlQzCIMdO2MyTmrw6SI7bthJaDzKYBRdqVTZ6kWLpDQgimJtAQAcR
yA+xd5Ee00cV6O8QUbmGW6/JgUEqKjmnh/sgkqCUHU6BluuSSw/+OoetTpixYoyG5Y9TFsKJqAyG
juVxukqAZaE4/CBWg0ItKm8YAh0XcIBug4SZSilK3euYnJDH+a2OBtxqZASRh6sb71OPv5M7Wq/q
v4dKCTE3+gGNFCeHiJISAdb3xLJPuqNyPnmtzS1kh11kwe9d+o1c+QPgmfCNSxgCDyhyxADaXnNl
pPJFjGmYgISSnl8FWYx/wCuW08puua4pm/3jTOoqA7pYiE+g4Gj1+zsJbqLNk27zvbxFMtH2A8c6
omwhoQ7/2lvuKsIkB1F4AbBIyzYLNRVb+aqEypue9j8PsejNGNRY6UcsX5aZRmz8xtC/h0YazFo/
T6iv93Nlzi3WvQyBDWTdWfNHnW0xAFdFs4mape7HAGSlW0AvGjPZAe3QHSLYwQcviPrWwNuEwtxQ
HD3UPvY95ZjA3qKjAKab60SGdLTtX+us6x+vINAv6CydH5FgHu5BdIi2O841mKB4XTYvN2U42amz
miY42GlgrEVfcKgOQMCuLkyOgmKjczzMyNSYI5oWEHnK6nk6s2DxrZDCoVXpWDcUP2DnOWud6Phy
eJ+rsYutVvSvONVZA4e+AzMncQdYGOgdsdwhQl/qfws2rCY5vUY1ZSlH/6RMs5oq/PQsbTQCq58W
am7JKUyx1HzPm4HQKlC6ZREVuaBy9Qstz6wkVKEjx8Il/C6UtLZtz6pPLH6/uyoPzLA9aHMJORUG
g+kF0avk16FgxC21tXGP7sRlv2O1yWal4OdkSXd1cqET0KUCtCQ0uBotWkpwoSORNfC+s3ehPrWf
/PXhbLI/w+aksx52nOqHoFl0YsxghKHe2VkuUnsA4/i/13CfYOjcSs0cuOF3gZVVOXMDUO4yarzh
stJKaD3V7UAUzKr4fJXVB1b+xMjDvBfxUAxgltOeRaRsn5eQVkReBINJdJa2qPjvFZdJwEZrZ5us
umBQ4Pi5OZLQ3/jf/D6ziOU9zvVFAlwokd/+eiCEuupOVwZyBOmqFqdhQgyjV9y1j4WSfri2Tx/q
CS9VsydNKMZqIBTVePZZ5fYS+Wsfk0LmVVelM1Z2xFX5t1t+sYDKR+3kppc7/9eY+8Nkn2vmYMxF
BWNUJRZl67672WA6rH2949QglmszOKfGLo6ED73yjqxCgOQuZ10457CdAqOAbCt0aQ//ywWLUjoy
1ReHbwtgOA1c5RdBVWPiiYmxK1XSXQL0pLODS15RbKrPf02qJqZ8smTNQUb8nQCu2vcPdMqdt0h4
2b63NuvzDPZKS+BVnuSXN3iK8cWNf5RrSDlVIctoUufNbMo4qq8syiADlC4iLXl5MrNAjbj0z05C
5EY4NucJLVOY1r1mDBsXIKsO5WeHT6ap/pmBhYm/TuzUHHoMuhG2TZ4rEjFGF8zxOQiOuESsnDYw
+YznQ+Ln+zTS+VLp8qyItaEzqxiDi03azqPRvGUHkTFcZvQxL8Q+qAQ58vEw8sN6pj+kMMQaBPGK
sHsk2VSS9BjImlAnep31Prhbukrbzc+HFusc5Uu8eNXEb6HcvllZWS/qzq+jdv08o4wIrwwi4zNZ
bPOa3erA21Ifu570IGo68tybwmLQAk31NBkhbQftdP1wDcBnGvdnIOwnhqN6T8aewdNk/HU/z581
M/CC8Zvl72NGHeJuq2MUKzjYsRfFjYAdgscefqQ1IGblKYmUIStQ1kI3cWaN8Y0dH4QwB4ocYTKE
vHlfWU1VLDjw7QY2KUJEx8fGMjmqRumCcHd+3VLBxslbjlQ/pC13f/B9fslI27eCg1Vhe+iandzG
Ffk9hij5uI3Fe93cCs4qxl8GsTErszFqlZVQOJsueoGdRdAQjpUhDKw8zaha0y5oUbDZs2vsYr0p
anyWWcptUqSi+JCtwvL6BORqMXumtKK4ZkekZH8Gtgl+CG9BIrOM4G6rWRqRWoD6EyoH5Fx5Q1mE
xgb+PYUdE+5OyTsR64w3Xu6mdX06qCc4BG+tguIjdBIZ2ZxaN5d7D3doYx3mJ4kcSdKQvzhugvc/
N02TCvzIa7MHYb/+9nHKtIHih/c5MQ6YWV0L+w1/3jE2/QZgJRUcGqI7lyQkI5U0jJzy4CBpJUHT
XdhQfTfv3NKQCzbNtU2J5n7DgTPMIXpaRec3yNGp9FLPgAnrbYBd7+Empc3O6s3y7Cc9kGaUGYac
l2HaCG3pEIKCTbRZ6EZwuPVji5h5D8nGLS3k2U2ctm4KhnUFrjjEN7hi4rF2O4iJAH6lXM3d9BU2
n1m50P+hDJAcq4wIWZOPEfeElfAah2mCNBg2Xl8AWasKHzhfrIxjZJ56mswsEfwHVMidQzi36ybK
ocnDOpmCH0gjoyFsTkJVE8o/EqeYA+rwakeq8S3EmoeOnBj9biX5MrWCiWZaFB0AivF3GpNoXZMY
pk5LosAcz0mkm6G91XjaMsL+ks2eiO2GzB9WUh8WFMOhpwd7UKtxRGbRD5EFaeqKcOZ1uy6aQz8L
2IomyvIBsU/t6xs+XNE5tu8dljigdQme+jQIMKfmsvVxvIRWpq8hT6ps4V8lWsn0Fbn8tCNM0/2z
YyxDlsbrdpKzqz1XFFk0wMuFcbdUU1p9ikqsKfC3/GWwsJAjAhRpguEa3cNH7AjNRzPwISFauVNH
LaIz/mrZ07hxJCcnwSZm8irWJ4FfDGVIx3lbMdBInOLQEbiQSmC9hJYN3128FnIKlV/1uWFsEpty
pvTw/jpO1WIxoKifqDiES9ISNw53xFQpePsI6pkOOl5a9sZeF8+LZAuQVnib4rtH93IBq/ltuN9x
BCkorqMt2A2GHFLkoEwFlZMzE4xK/6PNiAIW232gW+PPhWlL8RnANTTXbmWLG27JW/RoI9+t6qoL
JVINVqoOhKxxDocdanHwatrix1iagRKDOFe/GnaIJgwIZmGpHubzuUmfjOGwpzEIQx5ikbip1yTD
Soe7v5wt9E/X5uPk5XjRk5cpKgxUbjW/wzVK2uc3Nf6mRHdsb6fpvMwFiOI/pIFoeuu8TOpbiLK5
SqqwRxfaE7N+JQSMe2bEnd5XpgyKFkojhqOo1Rzmalsac0zFiThzmWht7LYsjVz+eaAzfZsWa0OW
us8RfEMwafXv59VTgluPBk0aIp9oPNw4e7eyXNclyBPBEfTIl3Sx4UpEL0hfI3jPsPUfIenoXfeK
RRY3/iOTly8pptWcBztPTUPHkxGsngmUFe07nZ9F7MVeDv2nv94M/6Y3/br38xI2Sp8BDsJ67Lrn
D8ObAIEkc9Wxs/wZAoJD4DBYm9bXGEOTBN0AjgvPI9BCsjC5rt8MSkrij5DhWA0CZekCz6R5yCTK
k0hdQ66AtWShjQhLUzGjUGROITPTBvJojQcZrc5NK01EF3pvQuyG5k8EKns32z+CwAmgJkZ2Oisw
dKcAo7eKg8Xdd9vgihqRfT0Gg1kijAW8rkpKO/D9aO3sOO4urc1UwwW9stZrYFdcgi2bkWNEKOmS
FJU540cCLzO1QjLVPEv6ViKY2GTVW+dHYDnbTOhAQH9pBHvMMLdjTiUuzJkS3w8kbLgB12ClH+Cq
TgcR9WXadYbWPZJgI8hl78lJBIq3Y1jsII9+YTtsypOPLgAPO9oBOQWFBedQ+HCy24iuHIOwZ51q
godQJLHmQ05H+2Jcvlc5MHSFe60FCms0o3GPvqWJDHA8GNd5ZQFmV0JFOPHlzLzN2TjcTzW17WsQ
5YDyJs9YJnR0ULZfM07Ef1PE9wFTFksm0K2FcnDVaNMHpVOlUchR6Y0MDN2uA83JdfcR8eGgpKXx
BMhZQ0RS+Q3f6WxsyTA7Y5dk83X8YGIzjgK1ZxgHAZa2hcediCrYOmsbwWN87IFV2L7hhyX2ejD2
r72bShnDyy/AeiXymKBbVU/OkTkwF9VTtvRkC56KB7qsAU+GxNSLNSpw/euJKCULpGH3vumsk+9T
4XrxRkgIg6HfL5ubEWEV6RkACaxwxpbthMRseryrGCsP5FB/64RMHPkEW2DgWqYTXDRvSn8zV4Qz
FVLftNdDSf3pJjqH6Ij9k7tyPmuFeNj7MrGm/2kQ3CC2Zb6bsO3YEBOhqhxNCf+X0139uyw46IcW
tmVKCFcYPDFnn7jrxXLGQRp/HuTYh22BJP6x3+TcCw4nqLvPIOxNN2eMx+kascjYxWj+oALGbk2T
2gnVIqDvnC8BkiecRpelgsTcU2Ur2gN+Hdcv5A5l1A/zYVKpi5jF/VFWCCvh6FOQxglNhof99nX2
2FT+56pTHBnHjkYbN9X2HvLkJGeraLe0WGptV/kfavwG/e7XmBdaKFWCoT6wH791A1UvYLKSCmrn
xuTU3fTIWnLUcO9JtZv3CaiwzWQvU5zgJQSdM1vWl3DW5tq7b7iG5IXE69GH8ShMg8r4eF0JDlWN
AzHpo9dcZAdzj1Wp8rluheo9eVGYV7eVdPsSRS76ZZo3uzdgvgHG1zV3KXsRJWAnpVjAey6OBuYa
+ZQd7VbuQDJEQiG11zyRtyFejQkwhVh5xRBPIqlcHCi1W5Iekah2ytM59wHyisUfLG57sSLPtGLk
0dzJl5l/9S7/uIg8zQvg1xSv6ATynU0uJm5xCHahVDVOtUN8OnxK6/UOR3OYEdMnf6fdc9Z5PmLO
LNW/VoVQ7lscCRm0FhANKITu0C8u0KuLaSJs0ru3T9hYPymcT1VMt0F7v6uBrGGc8hKi248NanT3
niOW/QVr/oeEiGj3onx4p8oBOBKidPotnImQoVWZZFQGviUe100cevwwmF21SY2wyR1tu6nnhKkc
wkxVHp3gDpAtS1CczjCUMo0KTP79tNtFHM1vsLZbPEcyrWq++n9U/S9UkBGWX7S5lfOLMu5SJmTP
X3GMvfa/SJuFiXHzTnIHQJisUm4vDnABqdMFhAJ1RgyDmflZ3tJXURKMQyzNXmCRqhEPUMWMof4l
40I1y+whDWtGrIdalrd9M30SL/bf8Y7flfu2pDh1q8dG2ySR/MdeU83cn986VPdcHOjm+NcA3nBA
JUiz/ytV3gFqkj9BPUT8XivrN3udkDt9kMofnxJ7g/9AXNAxN7yQv0oDnXTm6gOVpwthp/6UO6Ss
2FAkOw4uteFTIdCnv2Sau7xNbTdRXsbuMtWbqwvBLZM/wQuJRUGtIrAaPVKCBGMU8jxfMHP2l1p1
pEaxgHwBXgseOUTdUjU0kiqV2iuLQliv1biVNn+ZsUroF6BSb/iFA1Rq4yJzzD75giVdwx2frEMf
4bEgV0P6Xq/4AcJBqBIOYivV35KM6vtcSFQval4De4AGK7YSxzpws0qQDzdbx1FbPKvVXNU6VKqG
i0FdLjy0PTdP3jXY7gMEaarexgWbWZtCgGe6ID2UMX4nXKkmpUXsZVwHpfc/vT4p5pCLh+FyYMOi
9x0hIJdfVH02ZxIE0HxV6/OjzvkzY9PCAtFiY8N6QXd3RGF1DbQCiriGwn865/9REFNM3jvtuVSu
4bCynHuL65o0jz85gJLsP7Y8a+4gPp/bAEN42904wHLPX2SJj+Yg7U2O4oAtVi8uu2J8Qzlr3BFb
mGlTbULUdTY1Z3qH25P27NH0YADarMu3d5JPeo/OB+FPhZnyd+1cBzoo/sMciMbFofB9myvjgF8X
wdCy8lZgpxltyftSgBmDz/2rK6fejbovKbwL3aP/jobN0XntcJj/ueKkfdluBlW9mV0lmmpb+shy
PyVMnsIkbDdsCV/6r8S9rsSnX3Cp4tmtJae970KuDCLNR4sPP53RXhi+RuxIYG25UD/NOMWaE/Rm
QoP0H41vJOUAl9ZEAJ4+K4PZJPuqM3xh3gj1Ra9jBEp50k946Vw3YHgWmDd/U5LmC8/bdD40Ous5
4NUxrlklegNOMaP+TcD3CaLZtLVO5WM/QjD1Wk10V94YLKjB8YwElOC8GyCDAf0hYPWpsBqjPZMR
0EhQE0SucO6ke2K0nOiWTX7KN8rUKFu/31UiXLXSSYUQxNaDnILkpzl3a1HP51o5AtpIqSXiszbm
SDVvsbH50uX2usIr7rkfyIBeD9Dl+9Isw9PeigOn7GBVCXhVQFrcPHef4nMIiTpDHdqGbfx6zCVH
MHYRckVNVkOyvcZ2bBGWGSNSQg6bCLeyzc57/L/UBSGnVCfkwe07qB62jjvoXL+I5zEZwHWOZ63Q
RU4GseXx1lV/EZeIhNB5toFKcUD3jmhGcUv9nrEODSVZCPsk03BtfLt32g8OqqBQypIlSPrfGuDU
CBjQLPDhUGjUEwgLvXl0dxgae/4u46z48TEg0hocIul1TtizjgZBH5wbb+FKaVAnbm9VUSIrFX9M
JP1tA7PZYUiKxqFYiI2dqcnJs6KtlU47Grech/lsumPN4QeCxXipAsuKRNJOJDExIdy6cRH5zIcf
EqeA15ippAfTEy890j1YJe6xIV2YdDZ4ywWjyBSMoqnYZreW0kB6cGyCXv1oJvXtCCvJFBVV4umZ
eaHfmh43sxurW8IgdRrCtv5BVk/9TgPJWsu7bub4WpmNaGGqconJs0fH7LD5KyvO5p+OiWiY8Ggu
hfTo/vj6PiZh0Pou5EiBrJPtR6bsFLByFzqDln0GHn7rQJXfJWj9ANDBtEAVJqaIarqn+4QMgRRM
cYiNvRfqKEKHXgKkoDDOt+wpYOnhziN8ljfdoRkX2dtwCHwH59Qpx38+d0ZdDQnBK9WtAQS5+AdZ
qoaCf11ib8ARroDKyWkFRudpdGqU5ajIVyrMDxYsCSeHARr9rZIjHfO/fGBSYmEEQQeWZI/WhM51
f3eVtecmYbNcCfbMBXcRMY3dGRsR2NG9U6OHSPCVJBobdBL/2Yb+Y/QI9vBdfmxcb8J9MU055DNe
02hZ2cUTkuP3NK28BOWZ5ob29ln93gh9LWBOpriyZ2D4pUzclt+gLDY5tjLdX5Pu/q1hM3JUSvfr
qhOgoYzpA+k8KQtCYKXo2XOCudoYGPGFzVdwQlAJBiTA6g/uhhUgm8q0UdidyRPPxXyzaEzISfgi
986OiDBamfEd27aqd7/c+EVW7CTl3OgXekVBfrcgMKEdwvGHxQiJWvxzkpQ1G7jFbWBuR5t8Bsgx
3yxL1cih2Y2vw2x3GjyvweYZnkOmsKYyXq3tUYoFEWywiXGq3WTLdYshtZC5wnTYluB8PggOT5Ox
2MHKDulttoqH+eqqDSnb+MTeF9zEoz8mtg4+56MaTkDCfRMxULtbJW0ARbj1TUWdZ/Aq8QVpMMxJ
A9VCylH3bWP/P1I/ZfwfpZpF+DVaFnB1wsgYc5UzJPm88hkMdKl5N5UtQgmS+CGU4YBDS28t/uB0
xvuGjswxthHNlAggC+7OvSvkPV+nLILn3vB0vtWcdAXzqIROX0kcyFaQ9NL3u1dBkCFkGvsQ4ua7
ZWrl0QRB5Qa6YZ3EO9JCYKpEB5IZHAh6InOl5A0kkKnDmaLkVz1IFQwhPm2Sz1TkM2xkC0muEz6i
cv6l8CvkaXefO+j2ERiD0L2NF2UUHxiuMPKnuW3DBC6tn8cxJ6Mh6cw2fGaDSVbI6SQ6eRxRQ7qm
gjbBJPhPMfoUVU/Car5BXweHbic85HAUr2ON5QUyHSZYkObTBkpFUo+kAWEML9RQ1SNAcgNIAtMg
V2fT31nbI34jI0FzlKjPFw7luO5UlANNHxesXL5SwF8UGhPAPkt+WjO+HkWxHRbwo7BI2a9L7wqm
YZ/XMoCwojCcdlGABvYajEOJOMZNDuY/KXLoiNT7XwYaWbwxBsW38pNuWnt3tdWkJ0JRlAyN5hzq
7O+EthqJsGrm961EYrToyLkwd9RY6L9W9GHp9t5CBhDvmBwqE9w675MZGVdFqLNUjSh2QwgweFq3
Fs4qmjrNuT7ruqYn34pNR+JwbaRQyKFd2IBtuhqptLQa6LMl/njMpvnOsaS1I2VgXBjQcHqAfyNi
PFrf7mExWHXisYyoeP1AB76DVLcQz15Hf5BDFsNqGMMYapaCCs0hOkZPtrU5bHz29+gkelAK9Cfo
huv/9IXa3a9Ssov3YOF+mpovtj2nZjNUacDbR99dmtxWvOiTFmQ2DXqHlfxNJv/yqpPP4bTx8RL6
+GEpZK+9TH6Q3G6+ptd9KZrAuvWeJgpkbyBK9C96LhpsFFLa8zG1j2jo0xUgeqywHPOYMN6p8V7N
E2TCTkeQM+r8WVfb+RpTxIu463lkdhNRD8I7v18PKWfrazsqZLrYXmkWCzLKnZxGK37vRbiNlQdo
0QPw0niWkzpinyfD3dVvxgXZNLidGbpkK8Nn/VFTSszRhJOW8vL8Z8VW9Tww+8qJQjQD48m3kz5w
iD7eW/TrF5/RE8UWb/NqAMaDvVKu+Q1KZ4ym1Z2ACi2QVx1X+WUVRydjdLrJyLLCSNPyujbNDPWd
N1E5e5FalE/OWwdWrrmTcaJ4tPLoiWWtzhpJDeof3iH2Fgcd5xvWZvMl7ik27nFfpEvH89v7hXXg
EaEOd/GYdhoxLWMMeTICfZWdT4g0soTKpGr2t8XORhqD2r79KEHDv6394qO+ygHaZVwXuFWvqwik
wS9COeY5LJeYDTDNLedHiSNcylXtrcZiCGQZuyWAHaN8FWd6q9MtDqxhaoK/VbMerRWkhFj6zLb+
VIW0Hc20rwUSB61vO5P937DVcfSqtSZL1Jnbss2wi9Yx6egvBR+p+I30UZcaj4k7t7y/iUCkCG4J
kTSO/JmYdL7EKWbqcN6XNQadEHCUm+jlM0IZlu8DmQgUcO9MyBiEMSB1JeWPB+6yDvQwOoKXq1s9
U5fufTqWm0vp7kQlvWWJK/sMSLOu5dURROspRSgt4ZOXbQBODjV7TeJ5iHYQvLcRgOj8XbNSdsGV
k6fmuaTTXkTbj8+bgsJ1oEQYe/NQp/Khk8mkWPOHN/gbryucYTI9zONPZ9ikOaLYuyDb+TVhjwA+
LsgnRCwz6gbAPnOKx8sYNnFZqqIId7g8X9fK+N7dwXrK57Z7+5tufybWdUculUDL4UX5QuwdHsWa
dA0/T1yz5aXYU7CHxCyF/Yhl4z8xpBYPrCp/clLu8QlneCflSHAzQ0u8NSwwb2m+fW22XsCYqcVy
n0zXfYukdvJk4eMpRAinmoLpLzD+7rWTpp52D3U8eimXmsJVUUQ/xmRFYbN2ckNBVEPtgU0q7q1J
B23Zn23DND4rVo2QJqOi5z89/bg4LWAAnzEtEEQhc/RulysjDbCOxI2TAdEjewTTaiYV/CbdzjRc
+v6WyGznHy0Oty45iWS6rUFpdLGPS+V6TsCHuc+/CgzfnkpDvNxB+NdM5WOsmtcflutWd+E5zwDq
RhFTUhLDer8C9qROfTzf+yHGK+GiLuvQfI72EkrJfSjvXLKcl87ChElp5mSdlQMDU9znq6tfce9Y
TBCOdfpcPMmgBIiCRVhIJEFDLtN/QVYfCfl8l9VUBdwcHCETDOYAiPuYjdltISRRT1xYJUS0pbip
ChXbEfwCM77tOlEtdOreei/zNKjvqKsDSLqVUctLLThVLtpKOujqlnhquaQ2Vvzk/5v6DW0Ydsjf
9XY9spqisIWWV3GlJHm5dp6Q8Tykz2bYxzpxNi7CXMMvSXH6aj+RibaJ9kdtSJtb4hDv6md7NGTC
pETNUVW6O1qznEOxIAgD4h9gh/yWFWjxFZOMSWXu7luWh4u732eM6dt3LY/XN6sHkM86ZE+PbngA
lAPdC7yqK1IrS15PaWYERB4bR/RJ2jE6R3DGdQ9gpW1PR47O4pKANVVtam+oQ3JBcWSZyACLoU1y
l9HU/fiQ2Bu2Vz6+Gpal0/NM8pemE+lFt5LrdL2dzFwV6BBv8wwUgHilTOmeyd5U9PCHBbhoSYHB
6aUq0TVRbyz91U7zh+ARK5T4bxzIRAk0GD/QFg88hI5irMA+yl+dL892/wdt6yyGtU6mtChyEdhE
uUymi4Rf1zl08N+CZWlZlDE/PZXSAXcjBXE5kHaIkf2F2dqZWElArnPad75Bh7TADcM2EhFVQSNs
5Czw2nkWmSwj1tyWs4B6yLBwYKaczO/xpFppE37myn3WWsLih0zOO/BrgX/UQzFelKvWQ11fpzjX
9/QtmEFF2fEfQZeeLVYqML0uc0CCRKDtP99o0eeNyZjkNJfjAd+b9gEt3UypWeUi9ufVhJhye8WG
lvBdcvFI7o4a0xpH2LJHWPgFa8Bif+6HBBIp9ETkbc/AuoS19vGkkU3o63YO3qQll8rBHEoneea7
NKsVwWSutqIxeRoZbL6qSd/kOSzj7nBU1lNBCECFrZp2xGbC9M6W0V9qtWg6inZZHKCm7QBrpIhu
hZGPgJ6shHkG02TOw8M1xEiMQ3LwZbHSKN6njebYMY7sV9wZWG4Jf7Cp7P2C0iBfJOiSNRKUX7Il
DSnvHP2RRY6FTVwAkLMwelEUvOdbcQRO/KpLCTABCllXfq9aPRiZAL/yJ1SlQzSn/HgPWCszu8XR
H/vUEeox4bv16KSJqgtp3r2FChsJXxyNEizCsUDjKGCgmgfYXOLGtn7gsveivGv54WXYzo4jAlZ2
JiSlWnSDy9AfOww5K67Nl88I0frV846k5NHAnzoA/w9WPInB/dBYSLVIcTuQKyaEFwmIWu/bAeJQ
F4t5aa2zay9FN2t5QG2RF69XSHuCkbEzMvv8yyT3vsZuFdNL8zvbJI90LzSxExFLHr38RyOMnqLv
lAtQS7DaCKoQpboCgdaY7xWPZlbP7MxLpz/rRUwMfpIO7AHZ1KD8X99u/m0KRL8gQFzUjhBbKDDM
UcPel11B5IUhUm8ZDfXwOwWUeNigfTATa1+37LgKDMo0GW6nJyLyJNMvkd2yJF3+YtPlGF4Y2vZE
FwXBpqWjU4rokfRQ56A3SEFY//cfa4Z/JT6/leFhH9LUptvwN4O58/Z3h+TlTPFIneU27uVSTFME
hPRVI4vyBuxuQT+og7OToRODGX8HLE2uv+EONHeO5zGsC4MwoUG1h/r2b9d4I5SU9LWQ6Bqfh6kC
plNQ49t5Fq9I7TETxgDhQlM9L6pE0bbWZfHc+qeeBbDcv3n7FZBMsy9vFXR+qxbxe7kuYerupWRT
gvclBZNOn7FPlb4MucMRfdFkG9vmwzWALuyZIsMDej+faAmSkDFHBtuuZX7qt2/UEKflx3QSPFOR
B8zN4VwbobQXzHB+pRNJb+8etaCq56oSO5ZGU8ez6WbVr3uCympShg9soCS1Y1ow4AlLZV9rD+Sd
TPSk1fu/BbvjgwN2xDNL0AMPVW/PALIJHC0orZSj1NDbzlR/Lz8xcIiAWqNQHi30v6vyaDfh0f1E
K34UB9moXVwdXYLW/OfdAmFp/rkZpARhlG2dFnLHOLL8VI6MMbsRiKPpN432uvB+/+AFPI8mJm3R
JLetrs3mpQ5eaz3QVXitmhP+FIqv5UXGi0ldnfWSc0pWuymm5Zubs+7gTxOykSi5pZHVq9FqXTtk
b18HdeKy0S2syuMaCeohDDf0OJdrYsuK0rUlIP4jH688gTnvHaWGzIwDHboMfA0kg9lGAx7hBDma
2/NCMwT0GpMl8uWb51WxhZ8JJaUhyhlo86YKpOhs+PMzVdsTjv2d2eVHArbSmoSvZXQoiHjWaXyD
/zs7QyA3uIZFQuQnrBDG1Teaqk6bn/eZcOZZ78Y/TayDb7QQ3Q/xzk4gq2a28Fjvvn3zIKetbFyv
yFrMvSGj0viy/2B8tua4LMn00cX5d5kfLNSU3N8i6aIrbDfORxoQKPHl40tROb9QAL4rAp4NAjJT
QTIScmgv8IQ/pzRr9WjclQLwxGTXB/HUY8+CTsLUXdxIchoq28lspbwe8LA8mOxPDRt/gHK+BizA
sycb/oED1GSunKFQaO6B7WHCZKd1s6ulJUmczDtRzYX8skBWoWmj8mDkNQMlmXoTAvo5+jSgEH+9
o52XCTbkz/xTi+vu6/gplWvyOJD5KRiPALqDGUy9At+VzH7pLQtNEoT3ui+GbVKZjviOnx0zL+oB
y6Y9cgyfKztg5ngv0Lh4/DEDh/iAm96nEQj491EGx/wyVk0s7qEqyjEmm0uJoLbax0//URF5HjM/
A8dZPdqLsdnCvwLhpu4iLoS/ARTQHjuGIBi/FxQ79wZ+F2aKSDK7+UF9yqdk1hh/4yOX6q0eBkqM
zYVfaPrBW8C9XcRdIuFwHjDsiRwWhPQsPtiqrmgMiAllWR0BDdCz59xZETlIio8S3T8yEkgH0gLh
Ya0syn2VRLNg16XsxIaFYcIA3USDbg6Rjup1v26hTqU5lmgK4ud9xIwgImIhLxozdElTwTsUxR4U
RiyEdfdSGUHtCI9s03BI+jiyio8sUZUH/HyXuPthfXFrgQR8rO5nSNUBywOh3MRmjW1IpPhldICw
WIMlLbAPdZ2byQH+kfhfDr/zNLafgITkvBcLCz3/ky4UHsxvieci17DxwZAjPylAEAsJfvs3XuKa
K+17Sv+rWukyc6yCPK0Jr2uqvgBPiD8ZrfHeT1UeuVKuJeUrNn3OPfAjlHQibjvEGdo/7Bhb8uuR
60uzLFGYpMNpUAosDd1uKFRvsgCWcehpAjCV0RKSPwbzHKT6/c3MiEUG16wGJbnQGgB0za/hXobX
OUXcYMsEw7m9fknZ4MDdZCwMTXbkSdZCKDZw5ALjPJS7NbGTEGwTX+kFYOJ0aqsM6YP/R7ZEzoa8
HY2eZk8H3fXKtzBWcSzCfprSJLL+RTthFax14tk6Z3rz/bZrOsHLE7QiWEHCUVXMgQXRaRU/OifW
Ezbohzo5N17QWCGp6Joj8MNfjFz4ZmHaw9YupHbNu9YDzRL513HvRdvUrt2RqByCE3uUHb/2xiDk
u2Lb1J1H0q49Id9fDd3g9n2TxyY9IHRrJFTLzJeztXy0JxpDEp5iGJJAnYVDS/Dvvk7ZXDrpQpU9
/ojF5RfniOUVUpiw5kNC9IajG97ISZXQb5C1yU7UcraO6k6tEADyWUOBQOQPwn8z1zPszNMfrzmw
R0i1cn2ZycslpVruqrBSkpZcPQto8hxi5qdZ9tF0iFFHbKj1xiorRIDtgK8HSKulWExDGW6hYdWv
F2i3bUhiEQsT/XZU64mNJxmnBA5r5SOtrv4ej0eppsrfnV/0ESDNeYFzkZxcpW6LPpmYOHeFwKeA
bA+1fO3wzJWks2gagSkL8yoHNHWtgNNqa/tDHAqmtLaAwxqM3mICkniKtmxElb6bzSccyvtBQV9b
1UsPL+OWfzLsmVaYul2pXk4Y3TWOwXDGO8ggc3uUhT4n6k7cQh6SfCt4N8L0P2pDu+tuc+cULaEe
hzCsdcMG3aLOOTfPqfmyRxn9V28QhWSWFeUWmjbduD0RCikyo+0lhuEh8NIwV/FQUofq1OjVObgU
f992yNdt6994JikSSNrO9y63sBtyJHUaBB0u+JoFJ5fotMBf11wwiAG2hZlSertPAod5KZj1hgiR
rhSPK8xmDG3oxJAd+mLW18ZY6cGs7D4l3Iy1lGXGUR55Q2lgEDwUPdfEOkkDErDInIkY6DQwPpco
VGHhMUCzt8Qq3dbz5fOQkvIB0By1msmPA1cwH7E8VjHiIecjweZFyxsIy2wiZ9b6YWkvjRfZZ3EV
7PN2M0hnMINqu9VrmZm2QP3dezrpXKFgzPlRBlvOPm0cBi/JqMLOffisriip6jRfItOli/oc+IT4
2jpHHKeiN/aNRDPk+aSfbqinq0Z7Zsqpm+6y61wqdVWHCoa3eQ2acXgFiFS3HzreaXV/gIrmxDIt
2Ymfq6pIdYHfw49pfJpR0CHu72072uAX2kpKJMVr3tI+2U074HPYTlZk+HWjf+Cr/sT7G1qXPY/A
AoblRmvYftFuDnneLL64oQMqZyhqPbVZK5jp0y5N5gWCDpORENFfkY1BWtneUTHwXcuO9W0tl+gY
WwRU9LvW8zoT5fu6waHR46NtIE27SigM9FWoOMseDPPBWyqF/KvYhP96VzFBu1m1Shg2lfiIojZK
W2WB7TI4vZgMOii4GiKQOCNuNfUDUZ1p5Tq6nffd1KXZCRzsgyqWitZV94d22sRZBVqLJO8W6ojy
6wKVKImM70CAN2VcHS24SYe6VGuTn1vpf9YIx2MCsQI/MNTBXgstG7rgo5B28UwcPugJUkrDO0y3
kiRVUI+SUmsCDDGRH9ozEP8QsjaRCry9bnNsDMYPVljOCieYaBSYczX5fj/yaQFP6rs25QxxCl5K
Du8AB7E47rDpevzo/g6gEs7TB44Da5GJjaaPw49bci0+6q7sWbi5aCYHyoZ1tb147UZNTb73SRXV
/KRGh/HbjMfgHKkQMBijYm061OsvDFyaSqgJcjVA4j8CMSjmPVTUp4YgqFTiG6vLmsbdSFhvJIwX
mNI5wnBQQZnB0NV+ccE+NlPmPtvopX9TtsN9GERXzI2jBHLFKdScx5VGuorsgA/FoTCT5XJTa59Y
DlzZyA+w9PHrwivvT1FD67KOW9mGLYtI8fUGx3ceVww7mQVFYGdqnH4j/CI57SoAcRcYYP0qDRPD
NuxHhCp2giHRmYwod2cHu179GGVL98WdiBGVs3UivDIjY8BPqNpiSr16wXdBQqjI8hqU5eWjvGNf
mwbauD6jafCtdS8MCfOYYhwD+zqsTBgphZQWNfz364c39t7RcEnG8YkMuT6BHmTzh19q8ZOEyxNC
o2wkZWQ98Z+JiCt5ZGvjYMV0a0nARjMa073i0tIq0Br5JW05Bd3LH26Yxp/L8g3tnP68jrAMpTny
UngJhGUOni1NIf+FwwsgfZy3KIpgt7olRjyMh2n33fJWCgn7XW1m3hI4XE/D/d2h4qHn+Os0rNuh
yehLLjw9NRNoGSCZv1AwwJFi4mcSGyvScpNJ8f8iS6pPHtsHy10lueluGslvWyRux1tVPhghRd0Y
tTnOQKsgXXU+FlS8EtN1AgaTNtVL408F3Akz+LVJT86rQ9KdrNkp9LfLFO9r7VnwYNNef+1dJ9WU
Jj/+6MpCpJOe8esmkMn+8tWTq3whV3dcD58tpLGVqNT8VyQ4AiV/H6Dmwh93bulQaT+fFbHiFlAu
L00S7sEBJTBuVmQpL3Bh+WRCYPp9BUPMmYk8kxA7GsAB/Q5tXDH4/xknp8xPQK0eGE+bYTWXXgtq
Ja2JT34JGzfAp5x4J9DRQfeNe6R58751rZIscHiKT2AdnOin2L7APGQX642AnfZLtLV+1BqflOX4
uJmhrRpBRIKhgKFeZ7mghkzNdBdxww+BGMNoe8RJUFg+oKz1gXGpnRp1rz71LlrvbdIaCSE8NvtO
/kxmu46C1KumPL31nXRYF94dMc8KXuxFeOIL8STiarjGR+++zSqc93SdVcSqRViTv56cIl+5gqSW
w97ZVwNYVp0yIhpKIhmH6eKrjfmtCSL4krLPTrJirO0bXfc71EKRPN996+2KDrDI+amST/BNzZ85
OE8ktmYJExjKrfk1wJnQhbDp9PiKt9Jcuc265pLE7Vcv0wDzaWXPLEpE154mCUA14LOPVNMMnCEP
6fyS5d7hLsu/YwwAp4txsQs8KdD39tOrvu/F877T5PkCmLG8SzTAVsnuMZxNdLc+SxOzlFo2M1up
m7EVUmy86iqv/IN8/JflBvENbcG7cJFzxDSD8vG5cTgNEcEoBMuyhxXSiagOxGKc0qb2H8cr4Rhn
Li7vkQJ+fVOT3cpb/LFK4Bzdl2rgdCutfPdV+6+snc2aYEVRMtiMuywlWEBfiYLhfDhmEpdazGA1
xFbx47iGGrXfllgGgOQPg4c2Nsj67zD1cuyBwmMAA8366eOrI7n53ixHXxEMu01Z/q29peU2+7GH
3fymgZjPfH0Bn8trTbEmDeHW4Q6zBDTATFep3AABQyXsIcndUMj4ovrb2dvw/qMY54FxuDeVsJME
7rKRXYLBZsCBQGFAI1BCgFoUQwAJpIei4/fSLrLzhcMyjcLNTR+UD3WyGbD0Hb/uulrVGnsW50bh
91+YuVvwsu9zUyg3tYFUgNw3R54KnDvlnPExRTt+iUM7Gl/wKrJUUjuKcRDWvzOr/Zx1nOPLSg1N
D63d3v4VCEFB2wlfJC4VYfsw1uut0QWDyRU/myitwfsblgvfDKlQqk54zKlfuvYWrCXUoG3gXRjv
Ubv32O3VjCNo2smB4fYtRFLJShh8eAxrpNYlJyNaCsSNZi/epdqGNUbOlNDmi3J5B34A3wONotHy
+Bmvjl/OcSSpOjLnTUjHYLz0XVZCQgoqigVxi0yYDL+dRq9+5c0L6jWBwfItZiuKq/tIAdWYkF7K
n9nkFGgY03zzHYv9vki6aR3y3Qd9UL3Z842uO0xSTHCYGxFiWmHdjusOYtrSgELOoLuWWUW9EWF/
mUHObYq7uphicoVMLeJZnm5yWwdj5s1XEfbcQn9UJdm1o6oLqE4tKUlA7ioGaKo1FNo6zXR8f840
pBFunMnOSyNyv+u2fLKMyEzJJCOAafnu1hvWzwuMR7GAJPR7YNWIGJ+FZThvqfmrTt9bwK8VwP/z
4rk3BtCgTqXQXhIyP9P7oPFWuYYf88019GJRvBH6xafEhAU0iubSflS7Npz6SZ6CtAy0E4RvACi2
a6uWMbfZTwKi41FwBA38CkOqZWFtuEKNZAY9pbXyHr2LCSQmRR3YCkyEbwZuLxNyfMeSHp7qM18W
fn6RKt7GFDBrfSLBabHnwCNMgSZlDJBNpbrR31BzrwIbJpjjswIy/TRFY7xCFsqUscjQc6FiDr/r
6YnHxScrwdzekPP4kCosJQUiDRQgczoN22hxLOz3vaLq9RN9N8GuCugpeD/fbI0rgdzK8XnkffF8
yF0x0WM6+JzkS1TlVBebNDYIgqne9lI946eKlr66g7A/Y3jb8JilHL+Hga0GObjx3RFIsIqwWSG2
+VIOOCJyB875JG54n/4c1aetELbC0uC1FZSeCaA7NzIoKT0Q7PAMIfqFJ+BU20xuh6OzWSqSKr44
v1JGsxUF8nT2L+LUn8wLKN9vWVRlx+3I88BTK//pFK+EDkk90IXq9wWUcLxpn22M67+cd84KoNvd
GYMwa/KN++ugffMiGIg6xEqHuUg7ZnpkTdSUH5u6Fxzat/O1jXxk1wELeYzL5Sa/7mpe0YDuWoLZ
AtJkNwOHr8r/wEU7b3yUjZwOCMyqtz4yIEtPREA5kYyE7xtGhJRdt1BPkGP1RlSW1VLUg/+S8K3t
dovXEElt+HZkrOLU1BNEnumWEqst/Ui04Uwk1qK4yKwxj99ESp+uxGsGdZkCFeePGC2gd+Gt6Z8T
40bz7YRWAoA8MNPwjA1znjgWWkyd/wfZ4oIrjzYgdH03rylJV2IYY7QvrNC5KA1rYuf/dBV56dPA
zX0re8aUysy6QhizEzHSmM21COSbiPFQ2eEbxAL+4YaV1bSvSerwObXFO9Pbm+APz8tZCk3HNWNg
sZY5clyZi+PRQqu0zOHSPla8BydAEVWvzY99LxlrsFoGfryGocyuv1yiVX7dpwXAnv4D8JUeW3CS
s6sQ/8iqebu4oZvpG32YB+xLvPAlj5cl8jgf6MiMwV3i3aEyCnJn3jPobDy7RKS8gXNyXCMTKtzQ
oaY/hMbZCNtjB6NR01H7GeTPTym91Kljzzt1u1Gm0s8ncsBpVHZsuuVhuRoXJjfpi55d1mE9d3Gw
kXItJFi8LL6FX7V/oBmhqKIcyrcTmK13u1b4VyqAWqKATZjshClCZSUQ/6vao7cTJzIpQVi6RZYJ
jOT9svV0/e5KE9a1hZzuUK/p5jdC1ibljb3DRoj+S5m4uWLNLZDtyY4HOyxLv2RcOCzoh8ZXyNqw
dQKsh2PVNLEvTdU4J2/7emz6eBxr1R2huZsSvz+x/d6XU1933klg4Wa8NJnNRRXu5/a7voY8EqRA
DUtTUBGVoqlhFDA0OHa8Ys+3Q37m04ESz0ngTd1PMt8Qh84wDDJxnU5eiqGTc4aeANyelDLMvGXm
VOHX1c7STUM95zBV1AsI8HjwVksRrTG1cOZ5cWrZ0NNQ13FXQb4ZUgEHgp4ab2K9ziXroOvLPR3J
jwSOiyN95Cn7l1TEpJYVtcbIcEVMrMqNqgltspv09mxGO0SBzMJ2JAscUyhVXjG+/0m73i4agzyF
nkVNAfR1b2NYV4tXWh4e6NhazAoRm/2lmcF+vkWUHZG5Fw6xHP5cc62wCuw03D9rqZ6j9OQE3vuJ
JZkwF18ypxvsWiTKyUx4ESlw100PxVKvIjA+0+uK0V1aO92Zxj6dY5xzasggpR9MDqRSx+H4mpzE
BWRfOIS22ZedihaOLliqfgJQz0sfRlRk2UlVUjEEgpx0OKq08aoLzWbGtQ8SHbUfyvAgnOVc23n/
lWTZVV53QO9n3Njq3D1U3yRD9PzIWhyI5WAP4HXc8mzlivyp8KUDqmzbta4C1VqijVt6Ae/z3yi4
no32fooRpItqmDZK+bRhefkWczfuJXrw26lsaiC2cYdZLfDB+VxsPNOenrCKZ4IrO1iH6GoAnf4e
0wElHxBgbVku/5jhmYCJHSwLHfNNYBaDdDSUZxvCmJCYAQhBDpcy5/JEE6zG/XOGGBtsHd+4vKq5
Lgounh4rWnVTxvSCByItyIbxEUe4+tjuS+VFPzqX8DcV9rP/n4zDLEOn/BO3ZY8GcBya8wZoLe29
voM58q0Z5s5l6aYTON1/169zDDuKijrPDXZKGxVUuMH3zvrwU4IUDTGtWEUqQnhRiCjXECySCmYJ
yxxsskDTOkfQidZwQdcdX4cw+qw+yP/P+Z+EDaFVouJvaeyOOu3/L2rqzkADKrTVGc/qzWeDIY6b
zHLTgjYG+k7GLWfnpF3x/5o+hfSSiu4WmL75jkMXG7IYJFHXSpBDPWY42/4ilU7VK5jgGlHWZUPs
EZ4ec/CFil2I3lY/9pONjX2VnFSSuOSsLhZXqX3s8DLvrpof1D0hzoTGT17oqQosCDaAibrLvY/M
agPJAmlJwL8bKgkz1ODgrc0KTkm0/tpMxo8suJDDdlfbzkDF+eG2n0qmUJrpJ69s8BhyyPqRyp6h
UUIkCuKL6kBsEyfDt0nfKr4Z0CLagDXVRbXmgvsTLeEMKKJga9ak7waCQOuNlaS/vyhspISWGeqE
OCLfH2tySBOASlumIvEPb4DpRd/TKMek+QAApfzAfjQf11kK67C8Tr2pZX2zzmfWpHoSP2QiIEEF
hoKleFdCvXMi2KqV2aJe/UoWYMWRhmiNxS2k/lbe0Lh1MZsnUMon272kr/gD7WrCyAxPVNpHx3sv
hoI0EPodU/GyoH4vBLb6jgYLi1D480HgphEP2RsQqlT2gHefUmSbzTnUi2oxCXEi2w2XSME0Zo4Q
mSwgs+BZqibxByGU/oJzX0mbPaobUm/i5VS/4vQol31f8bn0C0oWMeiE2+Q/vs1Qk3K/k9faJdA3
GBVDXlkDPmQIqqWmgQ+HgiLbW69iOHX9bw/1gi6SX58NPXLWs08lU/SAm4lZ2+4zUM3zvvkwLIeW
k+ORlOV2uZaJl50Yg0w8MwwDvCPDHbyDvqyLMysoXhbJQVtjIvywxz9ZQirLGXqC9bNsWQhsNpfx
R/M8a9ZUbangCEdOGNkaX2skVNHTAj80c+D6o1aUbBvnbZLA5nB8gkaqxLdDK2cK0bVkWnMFFM/U
sbqAnuGCqniqQyg10RGiuVqabV7D36e1ZRpma7EislMPrYiRBCv175TGg77o71xsjvm8pOKSE9RI
0d1tRc/lS+w4fDhRiHYBV36WGcnmuq4U8oGGTKTU4/aPJ/tItcqrYO8AbpnHDoUonPlszvyXUsiZ
zutxqZct3WqPUJyigrnwTAeV32Vb15LTpCAulOwTxuolv3PbIH58g5okeyqhDjzpsV9GTJ0ryZyk
FR1xhZGU81QxxzWiAy3V0+TDCMUZOMM6GoY1LazcW61h9LtGEWPYiu/NC5QUjkKeolf1XHPR+8qA
mDNyPkcX870Psy8Fw91kutjSQbG5NnyQKW25QXyLSzNDVdB/x38VFGKpFoJWbqo7w1Kb3BfT1cbu
CTi5O3xv8iw0O5iMqvObjTdQ9lG2/mYuznJh8l8tbGpFVKtfL5p3UH80d0Z74NeKS1ULI8USF0Lg
DkYxrnwetC23m2jn5q7MeHcaZ6/iFUrPyXJdIDHun7ux9HxPwNHaHjVvFa7xoiV9qoNhoEvFwlVl
G0nonzVxq2+llQXVn6GJcUEdX2JEvbIqqSkuzauGDfHODAUsCMuWYGQ+JaAAJpYx2RDVnat/DyES
zn8vo1Od7b0yTYNcd1muMG0ctObpTpY5MQp5fcw9od6zWrpCfmorPNOjqhQPJmGuJQvYfIHsnNLg
Yj8dfVcd2lu3pBvOvKB/zXqbOgI3yg0CicYNMxsLPsuQz51jFPfx7x7uD2OQoeF8M9C4xBqJ0V4v
xpn+086kR7TdcGQNQm11zPYiBZbiPCjofFy/J2nN8BKC5pdwyTpu6W8z2N0S0BSB6DZZDZ5FgFum
mPfcRV420mB2e859wocSW6txHcmMbf0bMRUMlK+yeePN4aNt0OEwQbxF/ccPTx7A6YaJLlRji5z6
uv/083PPQox5qjaGYD2bslDZ9E+lM6PEBVmAVhnsJCaIa0Tbfc8fXG/sHIx/qi6OrpmyUML31ROW
6h+2ELhOGFbH/K3vhEchDBW8yKzLaM1qfsPThYggdGbey0hQQv2aTpDJnVhpU6tHo4Z9deLAZPvr
FomB2Lwu2pB8FJEze7DMZtcse8B9VTkBWqdXhjN5MukrpbPx5i6puniMw/hu5ZBlKOBL1XoIf2v0
nW2bMkfPWgrnKp9Hp+asofwoI56SgHY46nKRCkeo+KcyUZ6jAVTwW8NiV+DeEwMm2LE+9a8GHBIr
OFdMPxDuoLO3kYysIuMxfTHJSCTk45ZZui3rT2KlGI4ihI/bxYuZtpKpbVu0u6uI7E7Eu3J5+I2u
oFSH3WiNKDJkWKh406ZIEKbJ8V9Da8vEFZIKn4BrdFanncC6CU03QVQFET9aVtWxYKYCAmJPtNCB
NXq8iMBzsTdJ1e7eycAWrptQUIQBkrXVvhUB0HxX0VjZOF+GhH/CNHEZxPaIkinaS+X8nXqajeyx
OUVi/jrPAV6Gk8/cCyBtYZBuj9LyOV4Jn4KFTU9AstqVBNzc0FAb3TvTRqS4OWdDc2TcpA62YNTZ
Cpemnph9pxH4o3BJEgPF5++VLzXIBocuns+um1dXNSQj9OINNoZ1JvuYq0Hvz67NjOnSYJz9StSe
8/mvAtNkXpdmNxpl1B8v4e/36L+EguzdR5ipWpEiWA0d7XacYmN+tQUKctGKAYMcwubfh3wdHcpF
TayLHK3CqeC4MEpeEIVVInWyG83tzpXdjck8Nf7X/7i/Sw4fByLdO8nyox3caVBAzlDYruRkytVf
Sx0npg8jYKLF8pNv0GASD7Ftp2pvihs5g87YmyHaDg48DQDEiEVi8odSbvuiDHucMesNDSRkCE9l
Na77owQ/zHBog3WW5erCF3WYo0sdwMFypH0ZXBB52CkARzbXaRgHgvBKJ8whF5VuDBY6SacDQrys
iszXjye6sTJ3YcI6/IS7/gfvP5yKDNC0Wfyu7efSnVlfZ04m8NsvCgD0romDftSHgs1oGDpnU1og
rZz3XFPFc5EQaYW+rqHzxn/g8OWaSmxiTWVxjA2Fd1N4psB67gA72Ph5jtH8gcM6mDjGX22iZ6iF
6PhsU4EWjCXCVpbDK48dvbgD+JBLdGBWPdM0+31Ao9jZ4gMbQa+PhTQ728tH3kdz3gDBvjUBnz35
hYdzrUzoLrsu49kbIYFZ0e0dyHm8AOJE/cR11xoIITmYpbUxPmDOPOHsuVdb4SQ1pPZ1uHmof5eE
uKelZjOmQB7BD1as05VPFi9m+E0H1UIhkXrVj6jRovHzMO8SBes3vo91Ri+xMUYYGVGFs/5ZlGZ1
dQzTgpWbY1kWYXGKBtQqK2DRscqRxXVdiScGdczIG5qCikHXHHGVg1/YraVZ5sBJn2jUkJIJtp6n
IQ44XOhItkG3NndhEa1t3wiixWJkxJmB5Sj2bsgjlOf/m6fzr+6z9p10QblZhZkh+Wq2PNnU1Snr
54rFO9vi4kD+em+4XHqUrW5BzHmqkJzXt1FQfBhXdoadDStaephG88xE4ycBwMtwGU70ZnePGwR6
L9MjdeXMV6q0wo54f2iu0GBUA4GsKGTHA2uoul4wQqKJo+bKM1MSz1Zq3gNppyfh2YybY8XCBwFd
v6t6Rq98o+xLsPNFWA0XJRpTyyhX/EBou9Qr43MAvmmDl6TPJGqT/wexilHvhZKX2NigA1GvjgZ3
xoFhsaHKwROnDaFSx1X2Ayvt7GGYbitRLm4o92A54qSOrQjVlZFLnARJ3Ur1T+4j7XIo7wmW200T
uQVpnHK+YTJPt4QexjHyshabFrb+ZppAgkGDFidjHJfzdyjRphe69WUo2nioGHf/qVxjoJD3D1Qs
P3tBtSonhLsml4QCAXu+Tly9eWnMEN8YfujKgpjofjmhzBKvrspda4Nohgqfw/0P22LZqjeuCtU+
IDxS/LZRn4wS+EQdDWdZIkURN9YrS+V2m48MVEdqimkCJvrRQ23Bl95Hh22WuEFnK+qRHBaU0+LJ
A3ANZ69Ldk19HqfIhKjMHeDqbWSM5hRC5N9ikfqjiKLpJ4+g5ywHeik3/9f7dpbzdtVgPhm9wj4h
t9X+M0tBKshZgfamoYdnYlbcu1/eWHkCDtejbzCNOCSf06gjt2VpArDcsM/RnYii0yvNWQ2cO5bZ
5aSSUdvzSCJCNYbqhGVUXgNmDGWR7f7CC7/yevykv7oojL1ELwSO4zATGb4u7m+nMZnRHD99Vzqy
RafuI+b5iJ6fdxRtizq6G6a6RAAJzGEOn6zcIS5+o5Sq50cBPJIOwTPsli4jRcaUHFS7RuwqJVZI
BPWcMKmgdyLNgSMXEbfmpAPgdyIaj9T2plVOh/ScSXXKzEhgkkwfcOE6Klfhjg8klzY0Xnjaz97X
vdYq/tuq7iSoqyw7zm4z0s+WJxWL1nZInJ2OCPMkM84uM6DU7YZcuMeqtnITKkloQeviTDl/6caA
iGteEdmfNc2BFSiRMx+3VVvk8GAXJlYt1ikwD5YyuSjpoJBbWRZ1L/4l1hnOUwEZFRwHmLXy+h7v
ZthvlTf42J/8GTlp5Ou5Hnshv8mOJo0P5go5ECOJUsRASuFtJ02I+7dC45ObuJYbMJpQTiBZpx1W
bHjA7RcEby7vDJqWspL2RGT3fetuJCrCot5q3AjdBcDYEeSt/9vGlUqxE5JHw9yeAH1gTSt+57pT
X8WupvE3UyX0lEUaDqP8tO3rV1rajmZzNPe5lEVb/4EFjvk4ryHJVNnbBDGqWOUTiZCFtcZlORdC
AzAwuLu4ZaTPIdKTv7y6SEyhaLilbMoRmVJVYyctjp/34ArEelocWBgOAlTa9Y72rw56cCpGjQzV
o3xxITX2MEr08UK8QoNikpsRRjHV5YIVPfe/4QdbcYY9A1R1k2GSJc8fn6po4RGU1YsaGTNsRmlB
fkVz5OrdKlbKTe/1v3nn7qmBOiweRibbMZlljC7++3lay2hKe1GW2gk+8d7FzzLHatXklOU+Qu4w
UlxQYY+sMiZ8JCqrp0cYO4fzsVgFmDky2MCI/v5DVfwCqWx34Wg6Vi/qJx91/A4F2JMn5rcCVeDx
Qe4iTvHOju/qlAwgDqbj7pOPNBNpbzaqKnXygdxvxlcoNPTASAlQLRIkgMA8lRu9DEX9Su6zp64f
x+KobwO64LC7ylt7OhMwi/2nasiYMZW2GkxkB5a2foTCWr3kVgpwIQGSf3TXvDaiwnT4wTR5RDIE
4RXkbdSWHAeFxru/ZL2rQYHR+jLNcMklVbl8A+2ifxihjgzb8hnVrGV9rMWVE0OE/ZQEUId2zbzD
5rJdDz2fa/I7qAyetZU0cT372OTNaqURHNhdYd6F5zzgZeM6Ms1EQIjjkooOqCZpB1eh7tKCgCPo
J34v35WKthUynjXjaI0we9sLp2SvVPNOCn78+ymAzvg+pY0SPIDYCzRgPkd/aqS1kDsSxj8aOPZA
rXAliWGH3dBdhfM0GZ2EmnSeaXfzdlduq+72O1LFOZOO7skXKWqiMgTTIFYZH7ISiqSkZH983Z3m
oFQN2LudhPVs3X66a71d5EWS0t2VCwsYy1tRHw/NCV9/ZhywBj4HK2Ny4Hk2aOrJuTd62JzyAUXx
wdaUVlqMdCTL0zODPB444/Hxb34P1UHSYa1LMuKY/1+Kcy+9yO1RSImNAe3/vHoPgnribcNEQoa1
KUEz4+CbXTIwAdVNeuJOFPYaDdDqhEiv3b2+F3w3N1s4F0hCGyyFojFkZhoE6qfvPBKQqasBXGnf
W0yHPYcrH6iW76/MRGY40+f45jAeOuj8LOYOshf5oXxfgJb6EXxmfQgW11+t48Q0Nuayr9wvBM80
zCyonq32SDCqMMZ+bldgpE3oUu0t3mQ7hvV8tdf+GragxSnqguLvnDBpWeV0WmSaVJomCKe9+1+Z
YO/zZDLEg1ZHiQsdCf7eGZvW9sC7xYrKmk+O4kfGbRiN5StUzcBrzSUNwwUhb7QXrPYpUGmecpme
JrYhP6iV4xCpIQUXeoMcHAvn2hVMV5NhndBoiAQb8polYy9mSb18NuVWDsM9xe+W0GB/t+EuZeXp
3jyVm8WkMMQtq40hnuFlEqXVQ9dp3lq/V9JH+u1CcZ2EZiDKoO32//iYbpEUnGT2zDsfMCQQyLSl
5+beYEDLFpGutWCAT3OQx8BUrXo3MMQEQ0xwFPVwG3k39op+NWsp1sa3/TS+r8sV9jSooPH/LlLE
fHWWO/inerc+NwoeBDcCT/DVDWHpA2IXwKk0i7m8QvdpDC++5M952ERD6RTx67Hvjds5EyPd7h1n
jddXkGoo1npVJh+kxCia/cxPeIg8v5iDIWkGF607hcLERaGvkqyYeEN0k1z65Ym5otwifhFd/0d2
+3sZb38ti5sGJU1xN6xSa5DFp6MSAQ0BkHuW6Rxldk5l00eioiqXZ6C9+fcXkqoQRLCGtPNt2kP5
yFtM9fLVEFlz5DS2Oxw67nLKHRbgH3fP2+I+Gm2YOvtxWn28lXAe3IXjhvvOphRcNyqenUeGXNWu
/eGXrrJK3lbP5I+vPSNkl5YmiJyCqARogWV2EhSkTDvbn+x/D58+Wpn/p6Z9ehpZvbS/Yexl5jw2
KwbYQ/IGGIoq+HG+rr+UJ+UhyhvSEx1QxvIofmfpDqLfclSGFLBzNi3A08BRrP1Ca8q3GLLp1qUy
7jtpHqbA6uCQnhMsz0j8S8GLDAv+WeDFju0Khnv//NF/8BO04+s3Mdm1LXX/3/nl2Dkw9O9AzcHw
qzitNR8hoHHXqu2rD9k/9800W14USOaQ3gsN2d+4dqjUuJd/rIldcbGBZhXz+/Aa1JlvutSYL82X
TZ+UllbZnayqlMGkBi0fPIJMlChnsR0NyhOVoBA3X97jIkHG3qQE9Gat59yElwbSP0squTvtB59f
XyLH4UpKtfZGZZi9qIXi406gXyZQlKz4l/4iHCxz1GbYZ5tXeBFHNDTN5oYaPZG5H1rGLRS4FczB
lR3Ryx5kZIy12+DBq5GPTJxdNjnQuH7ZCbhSd9aB0c4cQKTQ0qfb+7Fef9odrHCe3ICIce912cWO
U2jLD8BWHdkSgdM/TDPPVjcF8LvBsXMsb71akyX+RG40s3e0ZzXs5WALY/3mZveFEzs42C6sCPqj
9CkCjuapFAwAA5kLBRfqB9qnf0OnHfagiDO780oUmy93JHW9DFZ6XkpfDVXZgkqeOWviRh1XmDJa
onnfVo3BAkQQkuf5pu3aso/xPRhortd3pexHsW+N6zpry0u1jTXKgV0/E9XeA++NXw5C9wqpUTUD
r0KhnpLcug/HY2W937+SPAMGUbeAnbJsZfFkwGT9AQnhW6ImNwWVOfzBwPUyKsS9zt5vpwuib6M7
lDidPO2+uEBnY+LV28SAd4MYi+SyB6YJLzuiSta0lEeL6797XE2sV005lWdT//ReRRFBY5QEpPxt
Wy1xiXSlub4OvjNPbUZLdu2JvHIOafw+hnKSwKxK+NKaaqUazxC8/cUy9Nr7GXG4DG+4LXIvF0gj
3CZGdr1HA5y0sCfoXrYGmxGsfwyqJcvXEfDgyTIE/EKm/z1T6ZLdPIikJriS4SxFM3kVDB2KUV/q
KccSj2Ovla0jEFVfcbOR30XzVeWbTQWap1NHNYY9Htenhxm1yqCu5X8cfjfxegOXZWoNVpabrqST
n0zTavewo2KFb+8fOI9H3DRJTsSyFjUlq8zSInWThtW7BC/yJRtL4uK0msrwDKbIq/gz03uO5lLc
1zwsYD0OxtoWDngV5Tp5N0+Bt+fmmXvhEmPpXly48Om8y2S7XlCw9PcZj2odBjpMfMGt0z6Zs09W
eaoH7p1n9uqi/NcHbUoTRcjOboZc0IkJn4LS+/Eyk1T3qN36rH7qO4BxWmwMGrD21521nFjkQNlp
YIx2h7w3bEw6CPYfVkMlwai5boTj4xw3XzZrmSze4j86fUb2bKhxCt/tAR6BbMRNpyp2u+IzDGaB
7Qwp5/zejSCE7MDjNE691hPZcgu46hpEe2nlEGobVd9T8R+9+dA9nCagBJda1eIt09/3EPrCHuC0
t0fsbr5B0fjlr3/fe97TFyyeKEhzSe/rFW7iHsGxdrVGBQCJInVUEEGSTRNgMmIE/SN3o8NNi8rv
Wynq/9JWvhMurf+UYKpLs5TroUDzR58vrDBGtGIZPGMWx2rKZZE7AXEShutDQyVKpG9ILMJg1nht
H7YLuN9Y/FCGfgdNpOUxdKFlVV19yjncsBGtlPct6n0Rg4ot11vDzBDSYfN5Wm5CG3EgbMkSCGbE
tpFcRs+G371rMjIoTYEYJRky1tKmU0QEdQcwQyjdEN7CHULkN2FlVtLzmssQnuQWuW11pTbXqEWd
q8K1CLktg+8DR0EootkGkTbdnz8eF5uwgw/QmN7z3yZY47WXxAP1wN6wvnytXyxq9TIPJiOWP2Xc
1jX+W2PiqtFgKAiUMdgJLXonZrdYlKyKs41aov9C7km17EAbrYZfLoGc+1c6Cy3KKeyQSnjKnFK8
QDqZoe6sbKGZl8rOR56Add+ReL4hsc2RktbcEOoezkG8FWLnuOpQCRTYd23y+Of/EP0wzuRFlqdX
A7sNdCI0sXlAj270sng3/smVBNElhS7jbk8lHAyTwpvlJ37DM8X+FqcRsPDyVn/aJTIDGK2cHUbY
jVnd5IFwkatPUBhJ/P/fiR2qGL8JjLndypW1KLZCYtlR7ApHDOX+eBLxAIfoXnyGMdO/wcGHthAZ
e9hLr2cp7yut89Z5wc04sbWJvWCneQQMZRzTl4Ll3Qz7jXC3iraj+9GyMNR3144HFPhQm4dPev2i
MkNb+RO+Aeb/z8I1GcTXv4pw3hOWpwT/4F196SyDo14MkvUJUR5AH2AJSJIyzx6Qb+H7DwtxnN7l
qIqmlC9I/Z6Ql5TZyEKkCs2Jn42KX1aEVJq6P18AZvV1HRuGmm5ZG6V5qi/GxpFh6C+wLUUeldNy
0QDNBjNjTGsygYO87qYTK7TwxPUcA1D58Ob2+R8xoy2rm489bTIk7xrVBkjLWU4e3nG7q51xF+2t
jYebnOvSgsCK7cvGRoXDSyYETJb2tglZKP1HKGdn9v4I5eMfL5RSqXwi5ezZMBpBs+X3PnnUpEXu
p9I4hrV8fn3OkPaLUK8ekIJsoBUBSBlMyXL7fxhQDtePtNbMXviN5qsjejZiWR/l77/Fhzr1Z1Sj
VaeAcXT+7xTz12t3p+6dzmAkPpaD7MVv9915Y9sXuPIlikNYBBktFixsYqzJYevAOA4//lfJT03S
cvS9YecafW9LVklxKjKID2R8z7nKK8O5R0ITxat573qBNi2hTWcc50i38o5tY42ql3qmFltnluvt
LTLycDNjd6zU4Ii3BoLxryye2WJt/9+QJGyDjkvHqbh9cmxlA1lxmxw59Sztn10wG039O4Nf1w4V
+HBni3qY//l41tybkeW150jPlOFp31r89Rz+HndMNyqM5T/rpJUzWI6zk5hi/dVPflgtc/TAwWte
rf+3L1y+NQ/qP+KRP9S4YiP2HMmCNnr22rRloo1kk3e3X8FIlovzmZXbH8zeXePBAXXc/MQtP3Hu
ZqQvGCnegcmKl4iWd+UTDkqhTye2fXOQ77XOVvkrmPYFHfQo6FmL8pAZnLq7gZYO6KbnuU9Zf6Pb
2qNN5R1DM2vxmKRqFAN7pfn7pqVUApkgOtGRQk5+U977KnvMEXhkbpXXcbtySbITCaSBwjzZ0rl8
YiQ1LwqSvBLOHrljbEChw7d70cVO5zvFYoL6JqU4TEp1MIwCOkCGWI25kl1K0IFhukU75DOxiWWq
SwnFpdHjbjmlbhEnEDu9tS0xNNVxU3i6Kr//XWpa/JYXEThsN01SPYIr2AUJfTLB19f+Ss2zAPtG
CqmQr9NCMZgAghl8CzmvhjXWfPOcJox9TSeymw17GiLGd0ySi8Bw65SrEATDPr/oDrLWoaQTBG95
BUcgVYbgWfmCLNd9+7FfWWa4whrqjBmaSWkuvGmxzdPXtw6OT/pWJ0+KNoQB2D6/blgywga0U+ky
rTUVMLAgL12TIDct7II/yFxAnZlgdT009DL1gE6YmO2xys2CSVa/8wkrBbAL1iMdjLgfN4VwAYsA
5Q4X+DkJI9MtFPOUvztf9vZGDOYeCi4ktpD1XmdfjMY1avbkRkGvJoT6FeiDCB3hytKIhAzusmwb
2UrdGYeOWjiUQNqtpvcJ5xzj5mCzV3S3KpUziupKzXl3zqvBWNL9jQBQBDJof/gVWOqg6w1LICnA
yhYt2Ald/TcKggLgl45mCeg39QidHcrCECb/GVXdTg7NLHKKuzP/uzg6tkm7IRgU5yJ1CJM8aGY8
DFXreDhFmfstqxL8WuwLpmngzcg6LgG3tUA46GP9t7+wGNdGb53MwG7T51jHWh5GXKdkXtaCZCe3
ABlnABg2IW1WaGN9Wow0DPy6D43//vED7aTP8oq+HuTBE5YSAWz5MWf9hwnPrpaDrLF/nZEASk+n
IWCznqBtrUr12w40S6+mDk/fHRuFPoQzlQjjwoGKrb0qbCDcVeICsv1csCVYb3Wku4A4ZvQcZVyy
5P6ItyYdLMfufZwZFFgCVXrvmsh6FpOEltetBuN/DNV90C4kzQkhrHosCg1kAhQXLk7h2dHRfCA7
LpW4INLKdSB3No2fJN6pX2kQhedpAHSXldaAhLLxlRgmR71c6BPz3WQg0N/1cdHwwnJBmeEJ3LNa
uxMvObifA9w9nBDwT/K6DaODmxzB2JB0AHZiFxwc39MYyw0i6DMTzdHJcHfxkeqbe8yhSZ8gJ8aN
yhU5+xLFYw9/VlynecorbS0gYa8H4IFSRrITctZX8ovQnFKLVZHg/UNk+6ZemO2TryYDaPxFcJsC
OD8yHYTHgfw+m2aMhsdLa4Bk585ami9a027MIGWac+R4VhJU9lcjje9cbE/RqZJQFbQ+C+mI7603
04w+WehP1cPKVDVSnuoP+ZAZ74jbGiWWz3cnidbG63N6WpFjyGTeVNSeqEGBXwg0edHXVA1lyUq9
YC0o7VkRuz5N45CD2o3LiFC36KTKmaHapcRHksPudY1ofEQXTjstb7WvySbc+by6ID5AhP7+8TaM
JZZgweSjYTrCCEXUKewBECdJ8SZqMLKZbl/ESWXorRSGGAHbyLyUL7NePAPcxJ1rDF3of1IH5fuB
c7wBuw0quhQQ8uuAWePB/ZnU6p2Fpp7DP8LeJIbCIpwJ0dwM7N5S/pY3gGJJ8IvNeIvR3WY88ipd
/e1cJZrAYPETuCr0Fk3Q8sRoXLpV04hKBCvPDQBW3wnmtSLrJ9rNxenknGZ+92zesQ0lAVI9tram
QjE0Wc2Smi4/JtadLXVbWZHXPdRqMvtNGo+iuzX10AsLiQchOadmp1UC4gwkFRiDD9JSZscdFZfh
QplcvnFCEpef5BtmEEaaESHP8lybdWJ06ylEBY58XokB9YzOzyqv416okEvd08m3c1bL8Lh805Id
DuXS+Mjt69tRYzLed5z+wsoKLupezGOyYv2MO9Ql0NZrnZIvG0km1Fo+zdHKJ7UkO7HpH8h3E5TV
ogU5G9juAszNThKRvwaxahESzb9cXVUCR6mysRK7t3afAQMFbCHoNFylZ/zc8CDQX8i/DYNCoekS
YpHD2wkltDadLgMds3ZOtXo5h8Fkb7YysdvFTt11E8HFaWXCkulxG9RIoAA6Z9LNLJ9FLwE+HuC8
nzJoZAAA2kKQHj5ETawJYUbk6XHJqnzSm55+5MnC0JwDpedbUnUq9w61yNZEwhj/Pz0cL6lcVcPG
Ho7wKM364mzmmJlbAxfuHmC7DJ5DUeDNdPwxO51ibNdngshWXJo+4q4iWCvzAtOA/YiLR3HGSUrK
tSNPzX7TaXyPR+z0nbDIbZLGRiHz5UOPuPawp93iDS0szhRFI1BQ6srtdyiDkEX480NvqjSBIZ32
QNaJa8NSHEsFrlSX6vPzmESUWsxYACYirO38+SFScS6HEAaAcNfRD0qpdJGkyCJEiWOtqUxmpFA3
esazSNe7X9ILK3uZwJEfEVHVyTQZNZOUgz9cCQtzdEmhhP00HDKzHaNz1rcqAL6plhb+W4gcSzBM
uexgoPVe06eYT09GMsN6jEMybSMCcPsk4NqFduQ32JVNWr119Y+EcSPLwFHYzc4T0iVq2w1Boxzw
TkmBvtBUayyXPKwzputvQT1WKoBGvYYRGaPpKp5sHbcQvkvLSPevni89TDcjPDkgEijguwLaY+iu
t+MXVyXAz9xlTaJz0ddHPHyqZVXPx74CfWj2I5x9ZbGl4DfCyne8u6lVwRjXzoLlCcClVV7r+kpZ
2oBspHnDWrnPwrOzcSOZIQKqD379iVVDfX2UfsxeCRh7lz7mj+s0nTCzwJngc+DrgKdllRm/KoNN
cNpBRc/j8o0mreEzf3dy+ser8b0Dibme4G2kYEx4ficpcCAu04OolPHQVQ6jzcVq8TR8BBAbkVmn
UEVNPBdgzcOpyuEAuua5uE6Buvepj3J1GAy52AmK4T64J9TXsaxygIZAXO6yJYD2rl691kEst0vt
EQvNjeqEIHHhcAO2B3VL1RmiL0kdKLJXZ/kRbuWkI60nu9oLNVkpSP/8bdtMK+Qdj3eo/gqYD3ya
KzKl2VP+VcjNCcALFC//hO+UDmj1cUdxTMbKyGyuejA2STFtD1cDOYedMDNo0euYTlrTpaX5x+VG
g9uKbsTpubb5RhQrFLpdimR1JVcY43FW1j5wWyPkF7mKQYIR/ea7EGvXQN8fiBeQTIcKoxQiVGrN
mup2DViXCAbPQuIvpmWoSMDnAuTCuLkcfqCIFgmy11AVYrxDH73HTPWMq/3IgNK9IpiltKmOeFwg
+WcLsp7BcOi67O0ZxnUxEzQ6eGkbIpNEb+C1Jxv+ddDVbYd8CANFCtxwx4JLhMp42IcgL+DjQGO+
MKx3bnCJ/AhzXUMYGC+2b0o7mBcpS70WSqPa2fv8xCug/bAYhney3pPqxEjQQYIF/Y4wv+h1BtpG
McYXkcujhhPpE3FkjfXl97hbhN+dcR58s3ew5Q/jHYkG5tK1gpKjOUEVyeDjzMlLez138xb4LOv6
SkWRbCSTXJ27dKLxpEjwx3PNKwOYAPm5KxzTjK5A2p2PRhjCBGFryDbMt6iCwctwwyelm58NOyWX
TXMdLO7Xui9Rnzngu2BaFzPbkcEKiR75JqMzh+X/XrL+vaKArYoMNfxdLU8f6iyUwD117SWFAXh+
y5VKrf7l1dGoo1r2C62+H8w/DeucctDxSqmNEBmQjSbotjB3YxP6ZYwhkz7JvxRmSDJawdtmN1pI
Al6Ujl92vP9DerUSFv3DYYZOMjZvTIMlTVmX6sr3Ge2D58zVKGfVEsxGl4UrIruSf1Wa4Qy3Wd/z
5xBs4TyzWrdrZW0cHJNnO+YBF8SvYckSdTjvzTkDaCw6F6GdESmaUfM0Vml/3qM3r5v6tQnYk7zA
A+32an4Cqu8/rbJeToSPgYNgXYF8mFfoyolJnthsDlp7JhCapptp95dG3qzZWz3tQecp1XX71+n/
cGyEEfpbmnjC+rjgIjCVJorWnsYhPMTNvEot8LWiZ1txGt05HfmkN/vt2zjguWfHXDhT3LyyqOFm
le0V83IHb/DahedjP9Uu6wgTYBTR1J/dpVc3YLosWb2b9w/kkAQ016csnBkGHUe8GppHQQi+8Pgr
sVPN3vcYgiZGutG+O34fd8iBCc003/Fm4LTI55myc1xtTyGqs00JdIHqjrhSbl0Fr2x/gp8OutSo
trLapZbPC0W8CJItPG/dNJToFh823soOvtwaqj/6zaiKu5rls2/AMTkbMw0ae9oAMmvVQHAI3RwD
v1hRwRlZoknGr+u6d4bJcOrhdNSouKEmjCh/JOnoHJMGC/rdBie18hDm1r9AfVpKTVYMxdM3jo90
qBWlc/S7CkSjWw6NlCTV2/Rvp5O7WhxyNuyan9B2SaetSDRWY5lx2O6GUdSpbblia199EidFtQRc
jJXiDQ4H4ELE+YDkTgtIMAqPLeCLPnEHYQ6kER41J8yMPF1GhyPT2f0/tbu0oZ1jzqe6WOwVC6g3
Esuw56A7B8tqixAvtwbcq0OYRa07ybznDV6by40VWBHQ7kSjz3Mnla0Q1lZS4qGpJeF6AIo6Fvum
sGI2ca9C8HPjpZSsTM3FvVKhOZbHWs8bDdiRMZNzQ1jzLNJjiXbNBwHU7qAlu0iB+vTVSx+/0vIm
DDTEDx411uz2cBtYGehfB7321ACjRdw5cNsEsOdQCFr842za/GF2aClEYEojlRpW2KADjVFL2Mli
Zm3QRANrYyJcxASeglpbepk8x7s9Ru6megUkvPb2jnLcaxOKVQD2U7mlHncZaUrDOUaEYDezmMOK
i7iKyi9aDXvLpZsKjComFNm/A9FD6Fjx65se5HBwDDQEM7hrMofDTNK+p8oQyCfq10YzaYi/uD2M
1ZarR8Ii5JPF6Gl9OMDA6NEVaFnM/IZoHv1DK9JaHLMpKp0RPKbeMMrtnMgZFRGz/B2HrI6Z/QBP
+7oip5VEpePsoK58/KBqXbR9U2ypKwsDMAI19ggwP+kwCEouB50HvvRaX91ruCv54pqMovHtIA1t
EZ/TJqrQ9gdaOtMIHxoVX4KFd0kuveQ+L9SpOUcOCOVyhaOkPZ33zC+FlPY5NuCuqVHh2durdF/q
ODtbQva61+hKUajBOcb6tLnXineyl219prjrVfrQ0mQPFImuTK/kidMdRDOEpvClJuXhJO2xS8fz
Rz/QMOoLKDzvkiXmiczrMV2DnBfpQ1mPVc1vUsLOTDBt+ttxA5viZSaqd46vigqX0evjOVr8iEMA
1mioo+nM+M+Tc70PAggSZO0DKHQUn1ttRPvSmV24LHMa1MJUG3H8yLNreEzz5XUZJPDBN43sEUb+
Mbh7X7HOUWR4zfZ7B4jVxuYufOMcaTGF+rrzVOvy/ESchWXMp86imHnr3UDJYoDlZ1G4ZT/J9iUs
fOxYGqpV7vQDy8ckfUgnEjdTzmlWeY8zfJdTM0i9wELHc7hstTAfQ75DXFu8e5e+ykpaP4Yk0v4D
1IEwDOTqysbG07whtPnLmYChutzoGbdhKsFRKqj+jvt/ZkMrLqdgZIRiJSRDfMduKtZZDiQV3OHA
MzgHhtUemV7dW5Nr18in0kq7/1phbqQUcV1yOBGYiEkojXMBTtvfVHXDuYQZWHrcTanAB4axCjSA
8BMBq7Wljlk/Txd7r+l/aqiiSkS0ltQ9I8Eu12Os2eF6NZSQCrP+0UgnE6JVNexy3ggqoKULU6bv
M6LmMkd+Nw/ZWqhLz93rt9tOq9ln1x8qwCKYkKXLhsCDrPulM3NDKlc7n6PdosQkapIiMX+/YfSX
3oUtBVExlmaJJBtin7L2f5zxwWmPDcYLFCUTA/c0yu0wFmcCXN0K1Z9+q+cDuRg6J23SxJCB2vxf
HAVSEPFVniLSq59P8OT/AWF3rqJr7Ld9OiRicX+o85ET6gQ902dkIYfG+hqxvF+THwr/W/cry9m3
KMZCCU0tCPOxXio5kTQnhyPes/ZMVfqGcyjv9Km4rbxSxBCo/jZiC8MRAxX/ZzkMf5fBPDDOOCiG
vHBvKTh2DtJHBOsw+ekfKqBudo0o2oWvNOisQwGYADNh5Rl77MQFxC1OPev+B/IVVh9d+1d8BbUH
mGoFj4LJiSgaZo7bIQAQWVpDgRK5sKohVTdUjOv1kzxLAEQUcYZvAuYSDk6BOudslJI8PaSfW1Rl
NCq7kvbYHKCtAMKx3hWpVmdpPYBM2s2J64EbsBVRBvbUrCQm4wat6m3LQPNoY2yWhzn8DvyoBBOz
HfQ3Huwit2VWggaogN5hmjWvKusr4GL0J8yZSHUora1pBKfY3oyzTi0qf39E0Pxn0h5VEzinzyOe
SL5nir0rvK+VzGedJ/e9MXcRSx1yU9/EtuFyzrTyjXVsnlrR0e7jJTuslP7w0UGvHMlSoROp0Zeu
ulMixErTo0MRKdrq+koP/E2GHAfd+VEB0UIEAI3es0HM0RJ22utmaxWxaEs5OmRfAGuN2PkZOigc
2GXaxikfkKOqjiAtbdtGVunVpfaL8tLc5eXtNOiMX2PGdR55qhJTwAbKZ59hNjKOxBAwNFSsHwxm
ViUVJOiQnzlM+54dkskAw7CxZAtD3B4r/MGfbIpa9oBvxMBJuvf305O07DR2+NkQZeK8w3Bg+3z4
xh03TnfBav0tyP2s9QSPnj8MdBaABaOqY0xFxdufaGxE6WZm6H/FeW4rwb5gfiN0w1KuDSsL0HTT
PTxCnf0UekGsNaLjaksZ04iF2T/Hg+/1VnABMTJIo09CIzoCqWuy/t1QuoQCilkmx5UyiKuAnLuN
BwtGQgB/IWl5wnpXY+/LwyuUZVVwG/5bQIeWZ+FPTGh3BIVdsk7BaRbxWdJjYGoA5jkyJvlzpFGU
GJuH+ytfunlZi31oBj0Y9T/82MOzOOWR4jc/5i3zvUS4ei8wb/679fv8nyU+YSkt+NImkMR7Qgb4
A27vkkAWB0EM/erRZnCK73cFghUg7NtZanPv5LIjH2Gh+HFzVWyK4l6hQZy3X4SvMpva/7UenBDc
uM0ENOfslOtCeNDPCBJG1YOzNGUbws2CFUdbOi5js6MeE0AhzifDbMljvSr2t5OKcBCuYRTarqnU
254Uj0I89Jbz3L6wlt/SILJ3qbSzv8Cqof31Ce48K7YRAiqKmbfGEBRycD7hfuAyjq8fBDEQG18s
o79mLid19gSiADpkMzW6mHCSDzNem9S8e07FMa0lKPNs7bQY91U30cXwMXkYfBDi+FKvDUCE4NG2
LY15WuKtxxX7IpH+2EhO6iWPXzH6Dmm5mFCFvRnsJP6mNUi4S5rIgGrRh0e+nr9VEQpAaJ/oallD
7naOxwPcHDuHnM1wdh6hs30yOOUQMyJOOX/xur+iCCqSxzmvam3DWYQ8cp7ibCOxmwc7d3R1ZV5J
pD3yzKVo45yGqVhGG6IEpDWBdb6vZUbwBlnh6a0R9x2QxJrxloZSp7BxNO5b8IdeRTrKWsXIOt4H
/wd58j9NIKyI613AMsYDtb7LZqL/mCG35DnfbtwzxKiALDjKYyxYUT5xGC+YwwKbGUWQw3b5vKIM
+qNyoT0vssE3kWIehac2S0Qx2Cq+gaQD51RELMCqPwwyt9BIgvvHArj9VdW1zmXvZv2BI1vZfcAC
kHfPrx/Ci2BrguSuFjSOfeCqIBiFDEmJxl6PUS+rHe9oek2WJqXVVcnoYzx1sPrD14gGFPLlPY4m
8cKE3NwOf3TKBrcW7Txmc1fvVfRx80WgvVFK1N6jmCYr9Af7pFDuKFp6IeozcKSuFXKNYw1jW/oJ
/U0m1qNI1R+c8IlrlbmkFVSFYBupdk0u48omkBlnPULmegMd/G5WJs8b/XqEi1Lfjye10axHDLQJ
qFO4jCn1lV5hOzoALJN2k6TrO8zX/e+AXS0OV+Zi0GNumsELiWx1/0TkQ17IVc5u4T5cK0k7mbl3
o8pKMxIyjZyBiW2QI8Fx8Qnmsg4zzWPTcnOtUv02PN62P7bWdTYCn5mYnHdBvhtnfdXjKGDqnkLm
RsP/l3GKziim8p+P7Iv8mUir7vmnC+/QtesROdy6KIXJq9rIbbVDHIqspRETqagTvSSQ88aB6ebX
/SRjNPge+iTqaqaWh3lI21PRZrzl1vvj5E0oXuTkaG8b/8LhGMNOoBvKyt0KUvf/Pv7qGJ3rKfGo
7fSNfHMZ2v0TFEIqAiJt9WV+4ttnY2/+gPrBOfc+rYQ18ksufRlKo+9FfiS0FwXXMx4YTqvT4Uan
H00piQY+E3/nIs95LVUhrDCiHNszPO7yM+Ms1x9tdCCzSxEFsnChIUOSFPt1hGAgqCXMwUJF+qUc
Y4WlsIviOELX5GKpnpvTjZir1mOZW3nKXG2aSTmJUWqtRTdsTMNLM5V1q+qbPB28AmMrwNcV2Qvk
3s9JsZAU2Gbz1qxS0AOFr3mL/T3+QqcJofCu7kchURcab8pox3/KKn24y9QLPZ8v9GraP8o9fC6z
za0FpOesMWPoIZo1ixwOIuyMDLkpP20a9o/y5hBiXa08X5AlrNHnnXP60FoVL9dayC4WskLbkzeB
ctIxGl1ARSVo4yL7YsOdyF/LIIs7QP7cHSPz2uAgH0H4FQCm5BQmS/UE71b+3KaklQdPyowX8ieb
hJtE3ZG6gyGKobL3Y+35Cdnu55/gjcBge/v2+95StjhIN2Z0Rpi5JgPByIjjj6f9zm4ZOb5PfwZg
vCjj5wLMJrWf7asGQH37xVDTeONmcImJJnXQ7Cw/yQLhchFXPYjhXw1j5LcKta8KtFkNhVDGM0W7
7lJs6p28x5qogORs7bIKqrrLHOAhwUAP/w3D8JK3NkUDwG9aqKk7LjkZ2zjhYEexbuw69NeXChj4
6RKJwN/iPebRXIs5IdBn9EL1zfMqu8o0yGEN9xRoET3Pm9mIqyzycGwx0dlwneGz+Aal4SdnJQEs
P/8zTP7xO/E49ifArrXmJkbBtJfC/Ftsz3yxDmHdeyceGSIGBM9l+knALRvMEdxPOXuZpOLUuYxX
QurxKCylKn/qrUN+SxK6yX27droB9uOSUfAlIApp87nKf8oQzCfMiTlvpn6SRTanJIgDM5JEAV6r
U46LBzOrZNwU/JMAtDb8JyMzawF8ZmCy6ByDAuvSjaToHdGSuAgQez6ZCxn+JJurrW/yyYNSotQi
eO1L4puguz9M60bxm6vJpoGHb+gtRGqu+pY0xIuOONIOpSQFGyWGXuqfYzeXyCulA5xTYxZzJdsL
dpC0riNQ058iO1pFB6N8stapP4+eMHSiGXJzYq/cUhCjFVQ09POfxHnpQxplRkSNzMvzKpL4NyH5
d1iYrWIK07g6zWtoJNeqQ7A4e19F0OvAhcASSK5l4xp6G1nlZxuTzAC1JHldzDvnZtu4Y7/ilcLE
5dzDnYvVAKceTjpfB2JgiG+Ls4RT3xf8/NhDepQvsD1LgIXHtEyymhshYjpdyVR22leJFLfUZh/A
m3taTbKvvZOfXzlwHukEsxAdZ/a9d+l25/ZE0dwbJY+/u9WO5icWv19/UbiWYDWRRfxQGEqsYEKT
+lR+IB2pYhRaZBTNzLfxVmYqyHoCl2GMLAtHosbErPt5VL7Ezilo1nMHJnZXQLGzZQH18pMV0MCi
wduu1onSg14G8n94zOoKB70iOOC7bhOGbUoiL4DmQ81+7/JBt5i1cWHelkChXf6iIufFJ825Qa08
LDu06YYXxx5nXR4hACWrZY0FFI4Mrf0Ws7hwM/VzA4tZD1F2TjPSLKMrnDni0ll2naRv+5x2Utcl
9WOthdblu/SIOLGErWauFWkXpOXCTwhE40eTVz1Azzxo8BLFslHGBU34yREhNgxW4L2E4V2o3RJN
9R23t9Xbu2KreEHPicTXoOXwdkpS/NqUjm4RgU2vhUKyuQ15s7Vyt9Yg5D9l9u41WO25OZIdXsSG
HfHyM4yZJHHfoTLqctgxj9qOzGoRuCz1yUtlBGmToUd91ICz1AFG4KkddymMggpavle2ZARQPkhL
qwuz193rzcM1iCEwPPy71bI3YyOmRrUaTtzptdg97B9el1RW0GEyNMwzIkZ14sc4SBimHuoOe7SG
XgxBTG5Ieprgb04R3QYBWS1Q7WnBnOW+XUkUiJXJMtEcBepHSZwyN/kqLjOnjpuPKD5CB4eSLapc
4w0I7KqogtZeiT+je3MapnYocfDErZDPLyGY81xGf1UPQH6BzLsGUSRmLjfI9GEtdM/gaOKcorOn
kdQcRsfULGotSbBWL6hCIAN2QflbcHMOC2a54hQ/J+rmgIjYjy46LSks27cfxtBrOjjHHDYmTKO/
+jgQQzTDQtp6VHKAPuh4/BJaeuyReXy/c0n8UYROSAzXPLOLlW6itR64fXmIg0jVHnPNRLSeXsHW
JRnsKwI5Sf6RewctGCA1sU/JdNV4vls+o/NJiECbTy1LZshOLak2tllGvEPf/Lg/rak0E/1gN+2A
laA8MS5sagEljQZaeCpx4hOm+hCKD9dGInbgfPEe4hXy8CTo8vOQdTyGungGk4R6GyymN/E88MYK
lWoK+DS/Foyy2pcv4n82QvAZPRsycZl4jZW87IppnwgYIBgSIEDv23+THdHqIFa7IJLvahhFO3uN
CWj2Hva9/2Px6AQ//Zg+ewXr6yq2Q8MY7UKvCj+7DZgghAK2ag52Q35xMFDG4She5hS2kcEeZFRn
h5HQw5d3t1j3gNvtjWhf+ngLXyCA8kXdzYtWI3F+APe1U92CvLZAFj835FSZ31DZ7GnK3OkqIWvG
oSmp8g7TfxMkMgjYBq3HKGvr2nfgUZCABrYLHTqdlJ+brg1YxYOdQvFnDxTzCA/03SCpUuX18D9J
O+89LVv6BGXTYfy4pUTjFvypbrcMFCj4Z33tz12t5ziprkWkYyhrV69t7fmviSjl+rgZBP3666Rw
TmO5kMj/cxdkLcmDEazw8TIWme+XHw0hbY4vhV9BPsQm8UvM/h7zjgdXnC6fU8aREkt8aIRGCUVQ
Kz1DltnBRUTz/zx5W9m5dfIavy9+LJD/M4mj7n7RbSHbJLZefUxZl0kWLVCzk5Tj460L21I5VmQM
7gcc97lABFrMPfc14MUYFZ68vrI2qXE6F4W3b9zo8aoEv1RBPSpxHoh7stJ5tupqW+BZmi0ngGYU
Knf+sm/L76OWMa4sw657adABZrvYJ2Nw4c3Rqz0e2Bgq4CcSw6OOb4vohLb6QMra5SaX1H9AbiBM
sQ8sQkPKb213lBDAAftX3UpMKfWBfDAsPUkYQXq5QNG14vIcqhDECbBSA4kGDkw9bFxwfNRBQW4E
oWuqsN9sDK0jkhcBsiZhTC9HiXtVXhnMXIB8IXOPkdxqqOwFtgHl5BBs85Lh7pQCTNdOLYMOjicM
/wEHkUQZI42ydU2j1oQ5oWGwF1k08YsRSCXVkwR+K7EhYTYHfJZBKgVApVqADtW//pB7L5FjQKvb
HUhSqPz7Pwk7HetXMIANqTvIMduTtepzpMgMR4Iyayt3G5/5INWfISPvC8ONJkNbiKLx4ejfyrxI
WSJQaqmsdMMV4WiwI+Af7cKN7+E5EJMxuqzSTYN9cZFDXvCyCaJW/DS8uT4sAkeiebVRXEDdQm8t
cIAf8A8+8wF7Fo4gWkSdDVcyrlQz02wFpNW2QrhQ0j4vy5fNQ1mBioZlfBFiDGLMH7Mzmb4Pqhct
awZk3VZ+Rin6oUE86HiEc48vt5JLD/s2sGC7YWGkT62aVheo9MG3WR/Ui17SdGcvw6Nma8NsRx+c
1DEEwzLPWTFMX/cr6c7NGc9Md+zk98fwdXHfHOJKlSnvuL953iEctk/1lgP8plyggSSwIokAdaDo
vxCL0H235D2PU8MrACgJErB3f9hzrbH46giovfRmMvQX4f0yiywmD46oBSwckQleszfbF+ee4NFS
InE553HrSsiYoRcep5/kw066HzX/Q4M+hC5pkHfgnfIKdAuwD5a7jKfnZskBln9M5cRUJn0EJoiZ
n3RHuOXh5X2jxru1Vj/wD5K6KteglBrdQFqJ3nK6pJ3aSVXaSK//rur2fdQrS8R69yoO/0eT6jKG
wdZkO9FAf3ESHb1NkTqL5yD4cWCO2luH1223Bf7G4dp3Pz9mZ1dM1J/6KY4DluiDpol80GGy9hdT
rWuvF+PBAz+m6OadjnNxVOE2e2ulRxb/kuVAj23IWXbiE8fGc8zn2pDb6eEIV7czuTtX3wey5s29
E3TyhF2ltHoyum/T+mRctdTXiojwh3cWzxi1XPfeHcRWPIv/KRr3hCpVtsJ8ieFx5VzB/WiE9d5G
GDhR4qztAQpHfOsfRrbiOQJSw2Y0DyMv9yzjeFzeHhL93IwpqN4SAjnl3m/W86MqnO/7mL1jx+Z4
C7u36rx2nsydtkO5H3LLRdLy6l/a8S/Lt6B7dbJEarQSGTQUds6BHCGyCAYsVO4fhy9Qu8KlQ3Yi
GrFvhL4meBqIYgQmqvms2tWk7BN7dywo4tTncSiBpS8trGhH0JVqC956JjbK2OxQnObur+c0IWRf
qmm7cudNfYWEAFmZyWSL6sZ1grgRwr7gXtTms7Frwq1OgHWV6QMHg/W87PJc10hoSNHHjsI1kLwP
WxUsCLQ59VLXVW7RPb7a6XnMgspgY+NApcugiXNycohQVKTiVbaaplGC+ItQhSR4VY8Oao3wCCx5
ELcW1Zi9Ep6LJm3TnM9Np+llm9KXlZ++zPZAmTM6I/3z26S1BkqOyVybCcK/ufx+WEz/YbG4bCvl
dhP7MqkzOZFHc0hjz4Kn51G58bNcA+iTkLKeEukWbOlr6nDaILvlZ4Qo4wsuJiiXJA3Nz4yKAWMB
RcqT4ZvDJaxosiL0W3II3QbyBo9NsDCixoXRyFwCV6wmuWiKL6QnCHqrOrQOGUO6qyiraMksLcL8
JwaAaDcfFCFADHcanKCQpI4vMkGXYWL5uy8QGtnVo8yeNqFnnLDyiO5wZRDrUaTr49AMV8/KUOuD
/1iV6NrsYt2/iVRG/HbwEwK/J7CdhfiYDIX5W9zG/ZG1LzNeygSiuPCD21NhK2A7x5Se0wlRUl8S
4sM+A9F5Dw1VnJEo+yCucq2Bcc1thtKo4YpUQpPc4yJDUkWnWfrVlkg3DAaTNVdQANOceJd2sR6R
YT0QqLa715OA//DftrdO9zGohzo/osqVAnzs2UnzB+Mk2fzaAHImEpfq6RwIa/QjN6rsiRqmc7q3
i1798YnAR+5OA5/sXV6C7CmUVrQtUpbApjYeGEam6dXubMAqM2Jys0Vq20Gm6KeYf4kqBwMRlnQD
PpVvcpoHajO/b9ZFcwyQxSgv/vrZSEHEDqEFC/bZWMchMeZxg/hJHqdtjSASQBPxmHwmk87zV82q
U5i87A8UXXno7SeOXvA2Sh6owfovfya/xH5muid1vXE6BmaY7mmp/1cBvVDXGIqUnO+EraG5VgUG
ERjcJ7W6XYMPGWmVacX6THIPqmm8CL/0gUeJhNF9IB4l0ABKdcMC6PFr45aJuWzmBFibssfWKYmL
f43jv5AWee6EzlYSGDSMTilQ6r3D9gNFnOpUjMvr/CYTIF0a7XVhv4t1g9z2cMWoQWdog1sDES6c
3oTAGNCWHEa5tplE4jQsrm0F5uJoLRLPKa7fk2MoEFFMOJpacv0RltCqulqtS0DI0t56sPZNzb/q
uctjH9s8ZEOoDDlChJRNZBnOeVoyMoD4FiQMHmUS1afTG86WlEstkWtp/XozkFugMRrVDMgpywvX
IVdqOZ53Em7ZPnisUWjp1vL2PawD9MhF8ya1WuVx+WZm7o9zyBmrR3EiRbLGmChmQ830I5kE1n0+
p9omn2QuTWnDo7G67KLOxLQPnjWPwxj9C0TJzM4kfJ9u8SFHhE1YQbnEtFaHoxgndWyaae26Oxh4
DW6QjhprJZwpEZ3w8nHnxLktvkzqoegXlwLqyPUBVDznT/PmvOBUy3vgCAgcXkwUf6hdbw3F0tLA
ZjCahN9rQvfj4j4cxN5OCusMxnM4+t2AF2+zMTyoBAdR6VSqt6ESNalwgq/SZqUostYSCK9G+Kig
N+f0+kjHBXhiZBTYxgfkJGNm7hB6RxOgpXaVRcUHOtmfvj2DIECydsRAvsYJPQA5atIOuFJ1R4K+
+opOH6cpFDIyQuvYtZ9ttkskXsoOxuaUegYaaKETHp5EI7BnxBL+M4LECNzZXJoTxYd18Sg3vTsp
0kKhNWkjVbfcgyXTjRFo/H1SabE3MkAg6ChNnzKXyuDGrI0HjE1sc7VbSzoB0dLeLLczSbQWlvAW
XZTNTH6EDOwzPq5hos/St8bBRJFt8wwmkhveJUGpaE5OFoarIJovoQwImRLLmoW5zZI9eYQBOvca
VRdbFw5j5xi6PMkgsPLGgyxhfht4pMAtS/DwbuXy1w9w5GIIm+r6/R9xFk2yIKIJdTaMMrw40set
NNI+njcB1adPOlOFjvcMgksh2cmI5WtKE5Uhc12tWj30tFfBH0OptMkJhsJDgctkFgdP2u+O88kR
HoPihfkJW5xZRecoxAVPQhRLk4Q53FA3NBfnPfF1KLm7RQJzj9a6OeNol796I3num9n6GgA+k2mQ
fsXO7nP5q/W+4+AzVVHYU6oYg+kS+5P7C3SkLljdJzvfnUcVePySAyRjIOrLud2EOK0wkr+VnC0j
GODkfso6xpVOBWTdavPfQ13GwkJjhRBuq7tMef8XnEjVhzsUDtkcY+1OlG4hOa2NdSt4veCZ8Ku7
WsAUblwpP8oA1SH0sNPWxi8i8UBCtQRYWqW4HH0NC+ISvWeYzfMAdv1IJlc4nYyApKCvR1CJq6qF
ZXgsCChTKbgzgaGNY6oBkvT7r+gi2wFVO2wtc2AtFZ4LOUxBH6nrgrqqX4mpP3ZSw9BoNarsYuWw
qmrkoM2ETScxr7/oBU1IpOD2nY0/+5v01y4nmhseYIowtDFQyK38ppvekR1ySYg/3hrIZTEBhsAz
HA6R0sutEBWu8AULIRWeuHqp6DGRGWyWmwam4dVlcTmTm7vDjwr0F43f9G6HpwQak/MwINPTSp6E
vJi2bwR3UYQPoX1oVMvDhqDwg/iWmD2FWKLDnvPsh90rRNFvVoJPH+lKPX1vjyDhWqAK3RPg+wAH
5hnyx0MJGT8UZpUepNRRaeNkY91Spn23GD2sl+mBAxVKjmpjGPPEMQZk1fEgOMZBQq5OLfmp5bCv
cowNp4qPiC1xPVViGeYtTCf+JPd9RddXY5IA7cEVJrEcl5mREjeebaNxoQ/c5FIwu3LmNrjvfI8X
ZY4OGlG5mDvOnlVpjinYwUtWGJk1OW9yXKN7T2AuPynRqckvt6WX+f4QMaEG9fSLoR7MrrmvzhWy
EExri+x8KHsBJBgYj1a4GLpF+VLAKZRAjE9J8m4RuI3aLCS8n5v9rHKGHgk4hj/wz0OQXJEu/GcU
eO7ajoRL7YPw7tSEmfXe/gnIH89kUUDXcfWTAWIUP5qvRc7e8PdAdgm6WjgYaOdgchrFr959ehks
EGWZSDV4TYKDAOP5xVWoQnSlSCGxslb9gY3mGjM2FeHAZf/nhZY6dO1lPJSJERFmfNbaEe7pIfGU
J4xKiK25KDuNQ9It5zf92pI5WtAU/nwibAS0QzQoWVrJc0uHl8lCPGUiNhnUKBopgxa5RlREmcO0
ZWvYvaWj3xBfuAkAE5ftXBLtikx/7VMeBnnEHSKRq6uavMpk9d1z1hkY/BKJaISP4YI/l2tujVsK
Gtem8q9rBHTv0jpSBNvIOW6LwJqy1S7YBLxysgu6xRvsQ1kd9Y3bJ0cmQ7FoBJ2Roz/Uh+qFguKT
914Qw77yj/hUQhr+/RaVzWLtBDGNHXM0YbyECS/lYIvZaL2c2tsZHdIz7Qhob21LUWuaUalHWs0A
ULhAhnoq5Les/O2ejq0VGNjZtH8bSvi260NTZ0dfX/J4qsZGIm12n/x4gzAokI95LG3V6lRzyE5u
heSYPXF8siuLUaoO5RN1cyWWlFrbD+oRHq525NDrVkSnXMI+vD8AqytSE/NiXIcMrQuD9Pv2dsD/
gcovNtjiEL+6xidZPArBRMEg9QhIlS8WKU8XsLLPH0dY7V+1vf/ojRSBChICA/sUX7h19sjk7lPt
9HALPzzEpj8gVFuxHN3o0j2yFZZei38WLDZQYOKwfXSZXAb1ZVhAez/kVh6IsyKfGvykiImg7KBK
q7arc/ZeIuhi6wh1m2IAQvo/wqUDh1VQEkN3Yx8blcq0VT/ifvd3LNUTn9D3dEZZh0GgTj83iw1+
CMjnwSpY6XdDSTe+3xefB2vojKZG+iOFU7dUKkmcbTarvemJk5NScoy/sMprPqHWY6d/8VoSfsez
yx6neZWCR3KHiAXXM2TMPWC1fZoPc76BEGSQmyWTmq097Fp33DXZdxVe1vqDSut091Ncj8v6QtjO
NdNyVBoNt5ZzYmbZIbp6dSX8UWYM0Pgmm5ahrCHvyew/qcKtqAazP/wXFQlYVyTk+1mlSXYJ0diA
RAqYiFod8ZGaQTOhE0EZG8+oZ+MeUnDbNDbLmI++Q/Dj8Qp9moSNhdi59pfIXzlFKIT9r3aQeN7X
cEYtTSoHyjIP87rGDcoslp1mzl/55R3v9q+7QEk0pWx6fjJVclTK0dygur1oU85Gete7Uh4ccnVa
Uv2A0JuGcXW3Lxgz2ZBRNbx4xkyEr8X7jt9XKUFYs8dNx0qHrensOaLa8l7zGcvIDDOnO6544/JM
bCjwGpKQn0K9BdCcF5QVuWsBPBk8FO0ts8tIrH+GTJKW84hGLr5B275d0w6lfu+MOF2ip6ojdUJo
sy2INCR/+WmRT9C+i+HR4v1NQax74hUhWQgpmGil3oZkEZF1SgFdjIsPPsn8XDLQY9yd7RUddFlr
h71ZcEpyog7uusGAeXiEbp25qMROMYGG7fWo/JqcKjMBzh6NqVOindGBfrWSUzaTs6Jzl+scu3SM
koD9+D7da4lT+LgedI5gr2LviSC8KAd75AHckVbFqXsunGnmXhrj7ofhJbCduC79qC+CkcQSnY9r
CCVIy7f87OoR0mR5qef6c+er2wvvD42HdYJ6p9pEKQNqu412L67FKFQe8+XovknjLbE7iUvXtUNC
v6J36B7n36TdojvMVCVkBTpsFlECcHUHVSVKkbQPWu7VEfc72mCSW2dsO1qdgbXIRtsRBnd5kRsL
edNL9eyTCIqlDZI0BpnPfHz21aDGdGrrkwZnPPhYlYsLZJAtW0sumDPdfFODRmqLPmmfxhtalyhD
5u0SMzG7txsIX8R/zbCEDcoiiwvqzJElJbnY/LuktfzntRjLSb3K62eT4D55g7EphkpN9Px1Qt+2
qeSmKdT9qXqmWaE0Mi4nNHepatOmonFjdJA9PLX2ViJckqm0NTIK7gxFPomw41jY6VDw+8250Z/z
GZnzVftTLzEjoiVLCjp0i+m6WZPKGVepj7AK9v29ZOUIUDK/AA1FcmR2+S5MjC2hkosz8cqsOqdw
eZm2PNUFAS0VBWdmqSmYvERj2VJseY43ofaecWQaLa+rNKRQbTGfQf/Ij7DjNai+bjrJGho4P/Rs
9rmKvu0LYcor8TeTIi20iK39s4FFZgz2aQ90K2fCygXsnvrMMsqNZBVl2znrqBKzDiwIjoRfTyEL
9x7L1qiBn9+KZ8K3w1T+z6OC4F1yRo/6uXlIQjta9v2h/XaRkEXaLIVK58uQ3kRceRoCiFmYgWyk
3VVAW8oGd75gKDRje5MlJnskb01bcQZfJSbtc3diWLvqd5l8c1SM7EiU/MLQofKdvzytVhNEDOpm
3hjm6huewIPeJ9UbbDpOXo4qEi9D3MtCFwiHidGJjlLYRdjznx2q7JIF3c1GSRghJF37g46qKmts
5TxTSfEZ3MkGSMq6w3oFQi5odmDW2zpImCDU/+/MPzSKWNTecw+TQmd6IEIVZcKYw2nHRU0uy1hF
SqvDtLdL+1GUDKvFlBDaHyw4WdalMWyHyyW8biFA34wzRzUnYPUyCGJBEKTydstOmSwbEtS//7oQ
3bMmNhl7esDaON7Wk12wBK0Wh+HctKkAGKQP8SquPApxt+88Smi4dC80eSwZ931QRycZBhbgEYGt
wQnmySZkObbx45iYubg3qtF2GP3SMdK2BaOL7bGJur7p8N3YziLgYG6md2DpV+/coTsK1SVqYLHL
VuPJWzq35j1MfQaaOUIVWneDMM64pYGCSp6SyWFRTmtD5vS1l0x/RDK6V18m1n6yNsMD+mz9IHJc
nOfCvlmrlMr0IAOgV92IG0fQvcZxIZ+K0i9rVSOeYzneJZgNnrIIUBbzrCRJ/k2nZDNhNoQcsNl0
pD86AG1GLEDs7ZGMXYkDbLfHaeZAZUBURkLtwjdODfAYKtPp+g0T6a5PaKwhZkE6RC6TMtKpxHa0
QhEvvASgCZ7nO8VtooN+TF+Fuyh8PllOPUvg3fCFQu1DxaDR+J/fHVrUcQgf9N2oPIqdDu8TEOsh
b/wJvGXLRDJXC9uZ2SpmhrYLdBD/SNHhY64az/ot0df13L7GNUzq/KSTTmzxhN7tMGlIk9XMcr0o
SevzjtDJanA3GZ1365TlJtSq7d2jmKD7snvfqOVCALkCy9+OFKXtKjPCAJWfHXlvxj+GJi4WkLfo
3fXStlwPHlKKUlpHd8LKMQP1vpUxOkhef6/jq1KvXy+QSRr8SzOdK+qlrLAA5AOlXKRo/bWY2+UZ
oi2mlAhs/0T8QFy5Vpd7AMFYBX+EgjMUPMraTZnhq6bOm+0lBb551sJinbcwf/1K6e/Oc8jhYbpJ
ly1UxaZa3wirddlN3ylJ9vsMOGGi8pyuzUvuUvJ1p0NFm3g7U5X1QtOoJeLO896AJwnOwsBBzrEK
Taq9amf/Kx4GX+haDUARNUHBIrdskxhO0taEi6y62fo0ap34XqLS7LwCGm5vUUz6tA2Tl2eOwhuu
843xOubKb1jzcsvvBvsFAFDS3Ru48JwbNvzuD3Uy8Qv9f+dYQXOVtxdfkmDqcd/tS0ffv0yvOrjb
dMRI3l1V8O1FJJH8eVuuedWrbJU0TpGxmPsdBwiuIRvEGqJapWcC/oSumHxcAAp78wf/toT1PbN3
GvjD5b7/V1BVT+xygVDa3bHZPP6gqLNaSfDlEsct10LhRuRPP9hNpJXAaiZqCp5aLLXD5oC1SsMq
TpcuO2jUL/UVjDHAaMJhFlCtNhZR8C3uz0UE6M9G2SUZk0KCoimFuKwQyl3DIwWVv83v/PU4UXPx
D89JUBDbWdrIKNdUUtHQNCL1Yo0sXV/Sel1po61Qo1WfDfF31JgcaQPvzzna+zmbRZPEFtxjO3R8
F2e9H4SLMAxGNu8h9OHP0+ndb3kQLOjZ1g+qKVct13Lj4ap+fcSWYcs0tQkn4pzk0vMbaWXGQ3MQ
3POrrzTtCN4Q5xLC7aEDWygxAbOIojzitcnD1MYdAfp/zDszbT4eLBN42T6EqMCmxsp/Yh0Gy2ky
AivLNKC1T42VCbN35sGTpdrs6KkQ7zQuNIQ9K5lSL8h6CZzqM/588tD/GhH4c4KYKPCDHK9fIsOs
30HQJQ4kCyL40fkowGwnT/t4RRAbfcYMAotaiUc6g4gP2bAq87nKIuLbapQoyZuVDVWmQnXlSr0x
VIvD/xSaAL6MZi1dPxMWOUVFOGmQwL/CBMUg6d0G8CRfZLk4EP8vs1QfU4X9TuxmPQLy7yZFbg48
ka7+M14evqcnTZHltHfQH25AmhqFb0VnQyb0/DmI23cjUyhN9sq6eVmJssPl+Snx5B06QnVPOnME
0lgh0beHb34RBFZ007yYAP96XUR4xsU3+FqvJ+Ju80y0gJ4wPhzgBLYb9q5lcKm0DLFK5eAfCJzE
aj23NiTgow5vOl5A/5iWf7mrkZI9lFBeJjunwHzNUPO2N9IVog3ROGq1tz40AZuBvNqeuEgR7Ssm
f/MW5tVfL/7K5w0r2up3uJ3eddacOzlwCTuxX8dt6TCbN9GLXW0XS6boqK/QtbCclVooc61k17Qq
vr3q1pNhjHRZypX54Xh5XSBRp5ZMprWoq28uJ0ylbWPylg87Iygy+a3Z8NM9UckoBTxBcRMZ8lB/
YW1jG/ChaWWsgnMT1JkWzV0a9dn2KPwna970NSUGrOIRJat6Adm5vgI+pdUQf2H2zor2Mzuba/ST
tyGmmfurj4mifRdmA8jui5Pg4Woj92P3Za5/h9+5LABPwylo5v6rjG3pV2JEGfpB7yPWTK3X3bAC
l13mu/dghnGh/wSNUc+MTNAUn5Z5jjN3YD/ijRnR8eU5SW63E7p72lEBa1/VTyO+0B3zJK5Zm0op
R0a3PIhQQj6otaML3+UvpLpG3hUjA2NGRiAA0iLtUZkOJVVV1/kd7JinMqOzT/IwLXr3PFJvsWYI
pXUCZGfmZNF8rhDhgI7ioQJ5XgVZq28ROrzlnTsmbmvnc5Wh/tWoVILsEfZVm3ZRLx0NlzFOjEVM
aVo1K0BVV1hq6O3u2vJFwGBiV6tXaUuHpRfeOr+ovwieRiTdzexqsqP+xE1y+JWzuNmDfa71zndw
H9H8OAyvP8eGiPYNTWdXCx1+TKOlG9sYzqCUM+Nlgfme5yggrrwGtp2GSxmaK8z5Y/lqwCP05rka
1GIDYvLkwAT7icoRSXAUjcBZbDhm04FDc5SPVyV1BQnb+DPSFuklrB6scvhexHWJR0rfcQJ9GyYj
KTqHvF1L5VTcmp/CZxaElvCpfud0wFTHQsJjSrEteKLGMj2sHMXDCsSFMGNGQvY7yH9QiElopUpi
LsfPzPTZBRFFSU8tfzjseOcuFghWMsvAwoygKyq2tVNCETED44VzTA9SWKyPviJUvKc8CDF4B6yO
8GlX7NtgnjsDaz1EVP4ZwquEaI3Xe9W13voveFAKr4nq46eg2U7D9/oHVzD+7K46WPy96sPMLlOd
eii+czNERXRPTs/I4uoPli1UTraCooptrnn36judC1FnVeUsdzeRdQrm2kOFVe0OxXOpSoGvft9M
3gDGmFOL1uNrjyXXyhAUzXgw8eaUkShC0CFpow9OaYr1YjoDyCHlr3+eaq7NxA11NGCu7rdFOOBL
r5oWp90lreKowCRaIBYzTC5xRDv/BUb4JPWiYtjswtSJjVrl6k1KdtGtO93WdUMBTkEnYpFQghjy
ymWAdTR+PdxjIQ0eEdhr/MyPyfF4f6UNv/V6CQTJCPXtFYV1WkxyC9NgEHORlJS8fH+ZuXb4E2fU
seFU9L4vXqoEarNftOZELZ1PhZDgoDbz1vD1a1m07oBc8a30/xKaV4g+zuirYPc4wsAenjLdsNtN
55lbRpUfQ4HI4Tz2S5fWJuNXY/sw2ilUIzIymecckFiPqZN5MrtGJGJBG622da20Ow26pqUhgZmT
/wHdmbfNmJAoh4imw5xiUENFKBeGQUi914BoFdXurvcAefB6nofTJNJJjUWtPEf4Q5/7gBTnDaOj
LWI1iPF6hEeImNschZsFO7tLxnkuD3YbPoGBCKUYwi4LwLJS2vRmRvCNEr77z1jd1azzy2MOpTBW
ebRFd/kVFqZYHvZkVSKZPkv7DrcOVN1kbRg0I3J7AlXjl4+G/6LEWecKkaZccs1r6jRrHnGavkP0
dbusMRyIBxO8O8IIsyVViVI4bvL1Cokfq2vK/KbmaLOXJwu/W09rp+pusa/ZOnh/2QX/AUnkkBbO
QYfFMA4zRVLt8LG0lvx24onFM1jb0OKQQ3BtKRb1U5hQC+a/VOKP8npehLQK8Wg4sma/Evl1bl4O
CePuJkaNH2J7AO3OqithaSKkIePbHvhBeHTAUhXLsv4cyD6Yo0HE3JNX4/l7UbblkJyoti4damgJ
RBO47hEr7/FYJM5/pFT3hG5kaNjv7d8DEvsrlMxSEVNuz0JK3AvHozEv8DM2xPePjF3oS8jL8PSM
0rdeC14O7/R8EqaO/bToVeXZG7rVxhQ18QB0SbisluS7AgMiwzHZSLWvRY/BtDFcvsyMAWda9JNS
gz2fJzNYQCRU15taR/ncbu2A2VF5/VdXX+QcAH8UYShKDCVJ5KS2KfC0YdoJb4nnubs/y8MD6r91
CKI/vUXtLIgL+sJtIBWx6BHOKNLO5gnJ6CNG/RtBdT7U3ri1n5ZN9CrZs9GO3aDToLNeL5sMlgtQ
V+QtD54G5oGfcmCuZOLplPO03OJpYvP57zwYiDvsiLEwoguN/jReDxu4hkaHwYZoJmC1BQX1xfCG
Q3yr9xpCaTEIt20N/rtTrDCgkIXpday/t2vRnamcdZo7OaXpdhzYTGll6QGsi7f7GPooGzMUD3UV
Axf0F+SVQi4dB1lHDPNcG3m5q69fcavXiMM/PE2bIVtEObVyoMDYGJYfnY2hJBubEBIfPXTzQkWL
MZsIeNnlcSy/s4g4kGPTRllld/yrAVImfJkU/rn/XFffHGgQaMtW6nOp/fai3T5RTxVunj3tfFW2
QqXgLo5+pZzlfasbjk/FMbkzY6E9uiUaMSgAnT0oR11f+bxE1q5E92EZs979EMC2GqaDAf58SUjO
HhG6nL/SfS/CMr/+mxuBrg+GPLWlYK8wIGU8gX4m0icCz71xMyfnqVUj2unlwMFPIBYtqYlEIOY6
+mz3+N8Kdj/pYK8pn6rAyZl82PIHVv2Vjg4LB9HKVzdL5AO1CCrFyzLN9KLI/KVSppA6TDE0pcI+
G649PU3FghN1cQTvx2dYQJAl/a1kPtghU45PIQXokZDPQ0UlSHpZoCPozUAJuWGRlkb7MTO6NPMf
xc/1IdmX8DRCzjTxBNbWdn2DrFGI1hlMp9xUNLzapcmPdLR6tzLfHDmr3kUIWZvoqm9jT2VToNOT
BtPZRLlDXFEIt5p+OT7wLMU5+gcWofjCPNTGpwtVdeJjtXJxVzLSKvB33iPJQ2a+F0CfnokDo31k
+YQ6pb0YNaJ+c/ZxmStVLbXE/2k5QtXWZwP6RgVVPlCbVZEWCvKrkYxYhaV9cG+IPmzdKkoR4IUG
k5OQnEd0r4gYU96RJ7+Xbz9gjGzguwe+dFHBz7al7Yk1RXNIvCP2hs1NjajGeu2AnzjqfEOA6Vlb
k7R3GWlGt9mQy7UVlAoa2jR2G6NipTMVucQkqNtXIyzO3AwJ3/WvN+HJud3CTD8fH1zedaAHawxU
UFsIguU370X046mYwmUjWCue5XpI/DxutjFmB1eNuK+yDTD6AMeExUSwwfMW1rrY62kB3ZFcMGPZ
27nuC8RELPxPC4ASKprD9uX0D1s7cKXljneNHq8+6dOvQII5zd6obI3OdmVL/Qf324XPnt95CnN2
QKnTeoi3tkQMCvPLClEEIXOjnaAZqKGHtcSzG9XHv91TAOH4Vx1yuXttNqOJBoz/0kkDDoEtcR+j
6YjUQZ1VUfyj1sMYJvSGuVKb3Ln71kbwOlcpZ8/jQyshbuf4ihc5zlLzUYntPZxzHSSLYJ1/YupF
dtsNnPLgFLbrsztKAjtsE+o0un1k1tWXJzjs0xvy3BuEiaYXWkAiHTPSc5Ysn2gENZdxvWRE9OBr
PnnVidGkFEdU7gaCpCv7gPa03eD6xh0WuBl5nnO5slbm0jQIi7dX8nRIcb3gjzKLnAgTdKFhvLac
8ogRUBeBDxVg3+mJFtglov5Q1HG3ocWfEsDW5BbAWCtSuz3yRVtK+ElfLOewk5Tb9kHoqs9x/3RH
mwRK1YAlqzsiSMf/beAHISH8Wnqi2+HFRpp94IKbkntH8tIX59u6UL1YVSqtoT7jgEGuGV8FAmsT
SziOrx5t8ixt45awZGkfKpsUoAtTcxhAwIwefXYbnByF3H8U2qEdnrgY2EwrCus5Ixq7suTWaqv1
sIohw92jANCcMd1pRAzMhirl/S3cRfETzDzt1sBfI5zw2V/phIS2vm0IaswR63gtv4QsBuM0PGoJ
JhuUXedWJpDvZBSzNBl4F/zLbxeDMIxsvc/IqoWiz9dv+Z679x7xT4iDe1ZOzl6Jq8VumUjwOcF3
OiAcZgk+3QE5/ToklPSoacNUHUzKX4BxxqBdLETHCLM0zS2hE/DzvBvVL1uPOrUfcleVqgD2h6qo
VyK9WZaKq8nk4qTe2Kq+BVAwKjS+mz9q/jUzsatTs10rZtgaBGtWb7LMY2gkWY9TxukgBAH5BVfk
GKJkdcgt22/xFIIqJK12SGOEZeWsGbaN2P1AX1rVgIEgeNhYxmWsOxwcW94ePj24pxRKlcu/ATVn
jqBiQWwANGmtD4Hf5ILcZr3Q1VG/fTnv0FlXY2YyjYFB91MTfQoL86D64ozFokGQuaCjcN67ITZY
6IFI6FuCm3XEdbO75R03juQArkD7MvnF1/5o5Aed9I40Zj9v6tmKa/zGZ4SxdejznY13A2dDF3ds
dEMloXyT8zn+DpmPOSb0FTmsOaFJ7rxEt3yoLl9ajkg06hQI0kJdvHsjU7Spaj9Bqp19pX/NMloK
Y6cFXzVdc1VCTrYT9884tGnORhPcJFa4UTLm/zsg30Xhtlln3AIkc80xh70mVRWgWKKmquhx0rZU
0giY8mCXTVbcsiwsxZIITwWgykIyhExU9LMOviYNBDx/4TVx1tbQMLJ3H11014+4dYVTqzuU6p1g
W9fDFWZNWwHXMEM+ZwHC2DZdL1LXSMIyJCf3q2VUem/kexoDWeI4ErrbV0hx6JaWJKFVprNL+GKv
PssAICSdhhxcCErnxUPBqBrKysHCOktxGJF5uMFgIKdmerIYTWofen2wTk0WofAPHgtzwSOnHeYE
0vf8ZowTuoAJI9BrYuSsF/oAeDaqxfCenyl/kmXqo+LSUlTtNKIv9gmR1+/gEz9fyjdA/CTe4SI9
hFHPooKagjt9xmzWIgPaLBP+++sZxGIHcBgT9VmGaFeA8pcDFhEkBUU/IayPKR++O8zgDXwuTmI5
/M3g/W0DcxPQ5wAdKR7HWWwA9dkdhLcUl+gy5mC9etaQk53SDJD0O82p4enofDfH3Z3z2NEHcHqn
9gekZSqogTXNdaPsx+AshTGCMhN1Zkx+JNfwVBgB3WNQeeG56lxvm9ZCaN8nIyMP9md/aP16KNsD
38xJ1HvNxgRRpFNJ6Kq3BpyvtlHLkEAZW1w0Smmuw+noA8+BWyU2UssoFeD9ul7ccbucy2nynIsJ
lHYzfretG+RqMjFe5lGMkSAIOt88R/UbQn01FKcE46t16e1X+P0wUHsYkYgnMy3Jpi5ijfD6rcIs
OI/f2uL5hoCwY3evzHdNs2dNcUgZJs6ye9F1Mi1Bs5ZJEtI0P7Nw9TYUezzlsAJo4IfzQ7+cGt89
mw7757Q8qsEE9ZMLVqX8lzxSxSJVI1LOLb+NXeTQrULYRyCJwYImiaq80b87hYqlIiw3df5/ZF5V
SKzr+xZQms7Ir/HyFnCggc6rqM8VYBpnSwGBvPzQHPA6Iw74xD89DUQFPesA+4cAqUjXKFLHg0Gl
mXjutvOJ1D6wDwT7jO+CvG4oRFHcE///fg5Z+InZaxccagcrUSt9VxGO3CwokWHCZWcTETofcDtG
qhKExmOp7KmBhQi2avRLgITjRpHK96l89FD9yTNxbDIiGp3BFIva5j4xaVplp35ODGf5l2HnT2/m
2Ma5FmYnmt+982uhekHRWLJXUeU7kg+N2Krp2BTNuCoiwdEtnGW5JzBMCIfzZlM0yc674+aKHufi
RMWM3gx4oePtbDLU8r8tL8BtHYxiQUb+TWldDnUVd62gVtn8QecZKX7clZQ2Jdj58qXz1a6UPB93
C5ilpOJBFw/L5+8YFDwF9Ua6pDsbukEs8Ki4maTeJTG4Wcqj8RzDoc7yOwSzOYP0v0lrqf6b4MM5
gTxoetN+cjBoLQt2R9wyqN5GCHlJ5+oJUSDLgWaL/zX+onSZ2dsjaj7IWQD241YJthl6l1Ag5O8s
/NnRPwxoq0MqxFeaw0CXePUjghGzKcHbBrjz8G6F6te8+r2o4cTP6ny3WUrxqHNgiDVPpjqe7dnQ
dZ/sJMJbSCCnBsOYW/KREGXO2cCso0nEsRjK8awqPxvm3oKeAjCTr+SuEP6wzK9Em5IYOTtOTP02
MpwObieDT4cnfy7KozPqaqYXaIOcMLhsHZro8a/QU0FBvffPC+ODvSCJS4fMPuqC5Dz83I71qhOl
1+SnKWlWsJ1Z3iqO9n+3uCwYCjZ6F8UUgnWtEQdV/8QCsvojC/K0wnj+r0Cyzl8BLxFK5KA/Fcq6
DukQK/JCrzbaGG3iAJbPdCGP2H8EWUZij5NFUQFlqL5GbyWkJVNNU9tCIpeWMdiFWvuMwOp+Du1v
KJAr8zzNbKqVLd/DdFcAAYheE3JptaEuAIsa6mbo/SDuSkI56F/iUbUuKh7tRIWJ0yaHpgZnHnpE
erXW/ykg2AKC09Q/vlpBUi2+ZozpGpCNrUUWbFvOI8uQPhKW5s0oodJr4lXBxdlrLvnraojGix4J
lzCEXoSdXQisavKpGVJn36JLVGitHQGKWvTL5wdVJeLTQltvxSL0YywnCQtnlfA8hRWeBe4czf+j
7we4rgvJVBixEcTYEacENFcwBDHQ1VtdgEW9QIrsIqZPIL6VfSKzzPA871IdH54MSeWeURXvEY+C
uSTUexye2rGxPwOb38WmJXnaRyxODBH2kREG/O2NgIyIDuPSijVYrEccjsQBBY9M7S7FpVDK/Z1M
YadBt1IR7kZBMjfE2Nj2c1lYDx7utDZ7iq4qS3GNrYAm1dbyAB5gZKNavegAWtgfOSZNE0aWJ0gJ
U12N7P2H9OcT/Dq6pJHTHNxAH76eF3fJJnCcHr4F5SQQiYT28aVBGkuBuV6RqwAyNRH63kW1ohUa
4q9r9jG1Q+VP//vmRsakIYXdCEIqVglhvfkddUSIIDYJmhRpCRQDnbX79LWejE3mgGpnm7N9NxEc
d8S0iAm26nP/hWHl2Gkxn+CDsySZOpBlsmpjY4OqaqIwjoiTQB/zFstgVaRZvYlI0zIqWaGHBCfW
+NgecM236cjmL5K8gLS+GluGSD0WcsEb1DU27ktbgxbwCUKTvaobcUZNP84/A8fqb0Nwl6bPnnAW
WFkyfAcjW/VKMBfeYw9+hYOKFsOCGndqM8nCTccDAWbI1F1e4DhrLkSVLLf4kA+8WRE7Q7aw6yTA
Wx1Dmf/JY/XDoKZWOYrm9jQsw0I6hvkaAjpeAy89TOUbYvBiSOk84fWj6nc47KodWW+/oEs0vV7I
7i3Rw0BKfYKJ152QMjbumKug1AqBP4Ckw1YU/vycKTmFPnRYQ3snN56tRx0cg0IlblwpAgJcNfeE
so1KGM1SBKGir6211TAZzXadcuo3eLIa3aI+TTVl5nHgOsXf1/yMHImFGDXsyZ91cpMsvQRWupO+
2zKY2VM3iUagVJ0z4aEiHUiqyFzqB39+Dh1zStACXG1rzB6XJdvCCruomRu2wWTf136lJ3KYxzF4
6IAMsL4zsYMk4rBZ4YExX0imbH/RdC/N7SCoHrdlqPLiLmTHaSEo38tYuT/KN1SUa32be2wgGaJd
oUFMsdRHZsxTNxVr7a34HggvP/KcTC9p7v8qUJ3wZ8o6UaiR1oWYogcCPmOi0k9olpjnf2NCEgWd
I+QTvOVVEO8MRxBf6CIXx79DMdCtIvrQF42dvLo566/VS3W0KP0u7UTChc0ZG7thNnCyKSuaInqJ
COkG2pBYgKe575RdvZT037exGHBh5IRdhyyAfzjHanKaZ2H00dtTpuMNICX/NF3P9aklehRbRygA
+kEeo6y4M3dBTtew8BGdvwGCHgWgGlm9fSU8utd5B/ZdnrwZTATrTXDG3N2bD9xLUcU/WL2JJUs9
2sx9jz/VgDOZEtbLp7Eq7x82zjQyS9TAhbFAfaif0EZAvlYApw0qjqGk6x9x4ZJkQySz709VnPmP
I52wmsGV2CQvmsdU1bHihvkx/CbCoqgnmzFnBLGt3mqVezscyr3lAvo73xj6U9tlITWrxWWMUlEP
U+877BMeRiAQ9mjJ87Xqp7qf67kgwpiIoLIFqMz5T20sx0ENIDe26ihp1wONyYA8uTcmShVRNGQo
PlqfTdTj5wNAi4TKML9oThz2G4wcXvao6jqp2/rKC5sgpcdPCxn/hbwbccnCT30PUfPFCoyZvCyk
GEPaRN+MmYWQeOl5CW8dZE9zvUosc0LbA7i/lnJD4IF/nuRdY+CVqAVVfijbEiA3ONki6OG3HO3I
VzE1mG883sPmuhCEqn7uaMO8G7Z4yQ+XkwJpuiDzehdtt97adpEEMIChvdDL2NeTMGLQ4eQ2sI95
QhfwWvcJO3cuA8b0RP/3uy4REurnUwhJEGG59H3YtQw8jFeDXty23cwF6m0LNlmR1XiNJHF29zzT
rm5hS2YUSUlhmCSiZlLwW8IXoSrp7ldyvy8ERAeHmOTX6cQrk+0mE+gl1JesTLIYLIdiHSkPn2YZ
yWkWITtOgfww7RNpSsgzaXUe9amhaIlUWYkdcVGe2KqOPbrjH+jC1XdXPFEU+yNXV04RkjLA/QUi
rOSTJ7KGqx240039wpGqVZS4DhG5RHzffrJJrkJ82+8zsNWqCiO1pvuXYt6cpWaBQSK2XUUbdtv4
JyvVVr0AsTwzaIP4mq6TjdlmfpFMQr8zPYaMvVkVUyDQW2hv0qOeR3Ywvz1rmAHa9s13MOuRidE4
pbCrgsCwmI7pivVJmoCKDyntBwAuBne+Cq7gluPstSI9Q63Cyfy+NHEClN4Pg/ZB/Fj51dOti3lx
mT2OBeMOG8CV2Hs+DwC7mFalI88IowwG4+/sPTJZ8DV7ljHuorKEgGG9PQoQj43GYsxTJNBfG39u
QW7vkcRRMLzkv/dPWYLSggWTjq3sksLEvgNNPZidjFJWf7hw3+YWCzbPGmd1OdhZjb4OB1ejS5Z6
F+jMihxopeS5lyBaySeLW0W8UZHVg8LScTcuoryjNUUAi1g1ceX1QS4B6AmK913l1eL6plMeN1fZ
3k1ZJSUO2RDhuPAuVabbTbCf+zAIN/Ao0/Ji4OLJ/Q4VYR0JrxkfZczUoNeLNXl3UT70AAuXhfU/
4hqWb6CPYxIudpz44loNGy2MBfzNnSzB7UP41vtVf40ve8cyhczdaN02gcz00+3E+TeZqziTUY6p
+DdK3Q40EYPKeEEPpuVMQpnCJY5KvHHXmh2i+hAh/bLNC740E6bnFc+tyFipOkx9XFvf3ZVGjqx3
VoGqbxEhSwKohrIbMlOwCSR3w2t6WdGUC9FZgBx3K8eg41VsTkZYYoyUTlbedompJDtkg/nhxpIn
fVL6GhM5Z/JmTYnW5VARpnSGweLj8kpGe6jvOueoIneOIXxYQFicwodQoVbIU7B/IJrYr7a1UVw9
mKkj16kgxLOKmBUZIUBJcv0xhlVjurmAwLlkBaG9evfgB3/yEJ+O7B9TTCeuLndW62kg+LEGMGUg
R9mcsmINtaMNhVFmAGGI0wFAsxOepqO0scoy97zy7HMsq3SFLxD9BlbG7FOPTvMxBunaIWwxpgMA
FcChm8JYWJaV8PnvXLKEw1q0BSavLZEQMBEg9KE4WPUSxpRU0BbV+IiTeiwxCJ9Vq5+AEDUlHZ9U
Z9n0TBiZFUG1GDOj/LS7tJAT7MQX+0b/wQR9njLDPCMCygSUHIL323Da3mtyWGoSmduNHvf576Xp
2FH+NF2822RbCYoqDWzlyG9lO/y+HoM0QPKxXAoM/vmk++rZivBNzQLTOmrEaq/ABu2RgGykBEK5
tUB8iQLzAJ1W5NyNIhzR28GQBBgIdBg0fUtwUZvUgdKN94FJerhj53svKnVOPh261yxM7xWK5L/m
Ygq2B7CiT3K5riDTuHeLbJOabacUl8je0ErU8bVso75EPUfFS0B7FrGDU32ABJ3wPeOCmsDsd8Dv
6hQuF/aJHu/umE2OwGfetOxHsUy24bY4O/UPiTTOypiZ4ELQqPr0GtFCBIQqoUygb06Ym1z5sjJT
Oa3FrUPq/eQ/jg867Q970y/FYPNgd1/7Rkau5D5e7sxV4JlSXRL1jeYXlZEforJKoT6oxpSivqmm
vgEKmsdehML5OC9NeQRMyrevCw2ywOMWeeJxu23dWgblDoZ6hfVhL0+YbJGQZrKrnshR6wgfEbZ3
rDNfLZHy90fPWHRLD7Sn6w+iREALDO1eS0fg0AuEyaLbmFj3KQJoIGyuamY2iymSmfkghqKBiPVP
sQyZSfizBTilYM6vPxxBhvkTTdnhdi06pLXesC4LgGQ0IEoUDgKvFDtOQ/RS9vidgRWynD69vjRr
u8Z9A1yo39MMMfH3vlrITJyzbMUDMzuCarv5MaBSkjCmrBXq3m0vmLM/CDQJmHP56jiIyzOWtiIa
cjQlwbDOWsJrJArbN3uT8BpbyMHiwg4vY183glU55QRQ5jEzsqzyzW0/iwF3hb8fNaH2HcALWH6J
zu2rL9VtoGP35uA5Y/2M37VYJdLguhmAL4cQ1WiybOuIP0CqoP5SPEv1HHOIYYg4FWPyqF8OgJY4
4v47x3gqVIg/KE0v//xJ3p1RSosCBzgXXjwB2qydIIwaVrMWB24V4A+3y2EbDwkkme8ol9dtw2Ir
hzLdR7spNO+iiXb7AQAV9eqzissoAkVP+u+i4H0sjvteaTwI1gEPgKbOLPZc30e3LB4tpsG/i6Oz
mdninoh2EDhOHWHQjj8Z7ArfHdyVvO0OZv2jn523zT7TgVs7X6NbUPyIyb+RysWQ/jFjKZM2iTmE
RobVraFoJqSSIOW59IYKw+ChyovOv1AmdafTBmL27qrwhrgh0X5Xm3nj1nK5gDIER6ffnfRZytIL
fZmdpBlHuTNVQ2ujeMGxoQ1tmggMRzO0qPbx4g/IUO0lYLX6b9yBJ2udD/JJ2oOQlzJynuona2/P
lY9otOXQO7LAEbOZIjlHJq0N+N1xc5cKUgUdtfqqPEyzZo+mmSQrQC4dDg5fYU0vhj9gjCRkHYOZ
7p+vR30HlHzKMsMSHhF6+xsUs5J5kOf/KbocO7k68QC69ANYt9F7LWOyDFdwWKagDig4ZmOcmn3o
BN/9pD3SKrJ8hpUuRSVzfykUAf4ObtWzDf+KqR85QA3Erwy6wYcfhTbkteft5FXWFMYjrQt7BWC3
uMZ27zH9ijfm6AvFXEO3SjUCxNqTMGeB5pDGkUNpO1lKGyAEFgDZvfqnL2o6TuFeop3E6EiS9bri
BSYjH4rmzNNUuoQ88gZzyPkh1BNWkfmk+gEwezpt1xZ4HagDPwe5Ji4PC6/36xiNzGkLV/IGzw0A
DFHL+OYYt8Lxb8iK4NazfsnVVEonXWhrpeZ+bVqlOwY6qy9767YVtbBnG4+18UGB0hvf1G6W003W
oreQMun57UwSwV/xfMlETS8Hk+kO4E9FToAJpRMfb3LEyCKZCvxXWBQRuIb1jZ1IYStdvHLAGpvl
7yk+V03vjDwSv4UXtrXKc0HEbhOLG9HIYhWPLwmPeZI25EdzGTKxjRNChC1Vl62ZSVQRLXfGU9WG
ve/IK0dOhkJFM6YlQkKzToMXHT5y9uh6plMdFVPmuiSbtQw5s0+K6NxvU7t0i83km2t4Sf64GAX3
EN24Vc3F/zYP/nRjHaB2t6ZOJ59bd1R9VJPAex4lu0HCKbfbpAp7+OZbtj7SeAA98zkele8rBlYR
IUAXsMyqdokU0tuFce2Ih12Aq9G+sLEsJauGX1dCkqSU1A7UMfNVpvVdQWPotkh9jON1o1OMLaBw
Vd289KXI0ciDng70iJOwLA/GzQeJSWO0SpwjS4bvbIlQcZNqxzgJpUEDSjnGIANWUIyuBYEGVyhF
MTaTPcxF3bNhINwQhwUvNVJmdDM1optBNj4zJ7NbRPNiwKIs0CgLwKxFCZReMtfY9oIMAV7aoGK7
INln7HSETZjnWGAlwVjY/TnVPPLwC0z48GUdIhos1F71/f5tplKQZo4Baso3is53w7Eo1Wno4Byg
bF287gpHkzFrzr+M0O50VnnYuN8QVr+lmg3rEbgDmssrayhcnzlod7g+jIfLYuEp417A5QJA6+3C
YBYy18pfRkGntBB3uevs3n+zU35b5W+dxrB4HyjPXh7ZkNkwuagQEghF7Xpx8kgftLBfdFxMrdn2
DKyI8SrqlE2q/U/rB9qdsHEfPR9j8s3acFt3GsH1eHiWMYWkyXKvFsoKfLyte9MJnseF1RoC/TL8
0b6EBUl8icsxaE/W6TV1b6hup/6NZU7xiAplA+mgCnyyfZKOHMo6zPm+k2nNBDYH9gKA8zMmBXZ+
2R35v/yR7RZApEuPM0t8ULNBdIU/+sgaU2DBCtJaCjo3YQ1nvJvA2OQRE2zhmVjTv66Ssh4Tg/2d
TjC7JbfQJyJMiVdWrVGKiME/5ltYOC85dEyANVRADH2Ku0EORGm53VYTKB6d69o4+IVMMhHkHl2Q
WivdAQSve7ifQ8KYUVMXc+ecB8e+xqh229CG17Vf0NRCHUOZ1GHOWY4JDxpUcWCIBq/o29s/4Q0+
JO+J5JHbcBVhVaUK+TKdYLdw/ObUOJhreqbw3MOw7qdQRCCyA1/YmT4HrkoVZ7Q8kOij3WxuWPpi
DKvUhTbTYhR/dLofnW/+4pLRuAWOMKDOH2WzY/5gZGStsQFq76gcueJf8P3SE9LrUEcmPgD9XkMz
iI/VBDSKXbL7fY8qbruWXJpi985/zoTtqov7PWN4u4avzEcMZuXE60mO8HH2X5gy479Upf0Ocz0o
3AMDe8PiNtbm1TdqxL+weyCoAZEh33Weorlx9IlECMHjNpJ4VECbfq7KbEIYeXDPtpE92DpyHgmc
n8lZ1TyqvHQP4STN8ppoOToakA4TannXDhSsJh5Sa6iDgL+r2uFwtgvNMZG8tsEjKFDJnSaj991V
79z3MxyybWT4BYD+AwVnAryLXaHuIFNPFEh9sQL3ljH/g8ATDClfe8oepHaPwSyGiNvxKbGzPpvW
zCtd/ofd3AdHH2JMSkDZb3gFn25wZA8wXSHwIT/2pb5Imrpt7d6xk0MfyrCpeqZ7fYi2mr+gIaQx
o6kHEWrxij6OuRUpT0h02V+zNCKv4GLDPeuXcV7lmrezGiWnGQmF6qsR8OccggdZV6x3ZFdtQ41S
3UbnJ9cvVj4pqx+k/3awO5NTAeyjlWlmBOQzvadjDRoF6dA1b5bLrpg0aU0tJRJoUE+nFAtYFgg6
006qYLhEECtma0l6hh5GFf3bX0sD23PF0pcuGphA6ZTK0Q+mNdMRebCuZF9vFVEuj3uWyPWl5rQL
aFcw+DITR6/1/FAJEvT0WsFiQ1DScDYebnrEaAOXVn7YD8UOVWRrTKCH1io7k4Isjr/BltQ0aeY/
ADdscy4ESVEHGbPXYbBRIEHVoj9BdzayPEniTHZNdJBZUBy+f1qsnnItkSkgT+UdT7Xt/w7sZX66
SvSACN/jnjPcILeewx4jIGksDEYLZJ0vSyPooeXUeRk43Pw5chwtUHhEF7eGp+nZ0fSPaLNRuZS1
u5nK6j/9XLWbnglSCxx6NBppKc9U2ZXOagPL2aZYPdOVblWAkgMlQLNJcbZMSUknzVf447xDgwh1
dzGAUdg6BWgr/IB+hNvBLohNswzJaxTPAahf8Riktpw/8vVBsDMgEHrMZ4fVba946Z7RVdyZfriL
Rxi51INPIAd6SJYUH2ckSt0nWRrRbLRL8dpTqJ/Ch8MdS98VU0cizodhVQvtBcl3YPo3jht1lFPw
qdaOXLebkZrHNHsQsD9KChnn+56gGcRHfojrCAnrdz8kvugKA5ba8UBHn257H7Kw/YEwEtBP7NDZ
sAReZSmRP/7zHQ9PkuwNTeiStqfiQQNBz8JIs5u6hP5beXvEvlX93Z8FDpkUER0HAFGp8nR7T+5N
Oh1mjbW6jjfjmSvOxBlMaGiXe6jlVqh8Be+N6LWl5Oz9hXYqBZ9yx9imLZI/seS1qgr419QjAY28
Zl0eQg9TY0TaOXAuNIDP5ua4Yh7qBHVzc+f7vuJhpXPZZg3jH/4oWF54wuZBpvWltJ2MyOntB5Bb
Ihv4EQL1XsbMeh5jtYpgX488u8FiYge1YglEfCe/O6RwzVzqXeyF6WTZ/GhyYxyb2U1y/FhZdHSk
oF059qri+Td5e+g0/JOXqJheli1AswO3HYvfG9dDcZHe22FxPX55VYRA66nTLGUfb8HwMdwU+uhH
fZu2jo5H88og+4l4OVOQUiwpTvCVz2F+ekAHctjcxEHUxYSe4ymbdRUPJlly5a/rSqRPKdaae210
CWaoUsOgQh6LXhkUaGOp+b/UNxf3wPw5aB1vyvn7YpskFxQo80wTP0o8v4Fdebq4SEZ4IwglRuCZ
1i1+V6BfKGVS/llB1pT1n2HG/TeSa5jnerTq1WU4aliwwCyn7UqrFOsKIcYsjSrFvcq9B1r83Keb
Z+7S3G3EEuU6sjOFh95U/qGlqQJUkS1t8WxlWF2aGdxB6WKP/la0QBsQR/7jaUK3Z9rm509b7Laq
/8fhwb11MxWh49ENk6QUlcBL/nkBkUts9Bte53PHC02nAkYyOpWd6YB+dzLTVnh4Nf9AnjYdorkA
Q65HOhHfESlRZ3+2xtw9CZ1j+XIjBgoxw/F92F+7zs1SXWekfiFyCCXefv4eG2k7gkIZ0hXMwEAR
rBziyR/cqEp41HlRQiPrALjwarzAXu7i2zWARkUk+i2QQQWw3LOpCsLp0cGMMmfmwLmSCQYWUy3G
77S1bwOAd1jmZ6KnPRQOCka6iyOayG1tP45h7PbjyPNUzV+Zvv60SCWzAi4FfqKLAeEi4MatSJ9c
fu42MFwjLx+jDX0AKM8VHweAbHqwUewduitFucSsKqpjxbyOFxKJUUIG5Qaz2cgThnL1KPLcaOyc
OE8CsxGSWm1vliZggWEyNPyILy1xpbZm2QpGAPNjdqEhd1plSzLJTubceOS4bsQiICodkqk/TBik
SbdIFwa5c2xZnDKNylzPTiP9LL5qeXo6o4ONx4LuFzMx/qAgOih41PCgnM+2TDtDz04PPaYBrMf6
ew6EvaVE5F2u6L/TjlVDyLYxDJaxkkalVxSnrty2bhWTg3oJDqjpNhiSlBhPJuCajEv3pfwRGna0
zLNtfgWy4Uf8Dtn4vm2so4tOg62wUBMMx3OP2biwyfEvGIAtODdNHOoeI4SRTdXfkBDjz4v7Cvio
vONrk7NcTrRjgJ1XhYnAwwyXwN6mskxgTO87cJmKRkAwzpS6+EYkp/7tBRh2dc0cIH15StVNYEDS
oxAW3pkeb31nQsCEQoX6TAtvvEjc8GogRgnapk/AG0G/KflIlBIOiyr+H0gH7iWhTxKAULY6Xwl4
sGNBFYmdBmj3KzgTzhiYy170g4ryDX+LXSjtcVbBM2w3myW3qSgFFtaIKR9JZgep/3t7ROJEqL7H
gwQ/o0bPE2vmTPmHIY1SJmt6AFpEH8j7N6A5V2djx3lbUnXPLNmkq0cRar8Exr0hMyTdhlb7n6bo
jsVKW5qN0BG6VgztjyI2WV1xvAFk/wOcAauqn447s7imdRNiLVy+owxv3FP6c4GBjxYGbzdzPq/C
PUMkKUHo5YHSzoITZFDCqkLWDMRMjAIDc8kCk3T0fD4nDj5enaMhbdCuUzl3sAbWlyQ3s/+BiUAG
PmWsHot6qjKJaC/Gx2USjEZBQpxY8R8GTLgBmV6/apIHH5OboKgRGXqkYl+TTLzVrbYVHn89hXhe
HP0SPDTQE1SCXdg164YQKsOaZVMOphcm8RdcaP6rxddaaWCy/GWFgWjlAvJYI+6rVsu5jnlJ5f3m
imTc/7bWryItYnlSV0YIfOnaSk0QHL6HQW/7w9hEBrgpUva01lSkGARnyIaWHk1r85zt+8yIP2JX
hNLO0dRY4PDSp7P+ghKAjU61gM3RlVsZtjJ+ip+Yc5vxs0FSRiu23mMll7RmqbyYVmN1zlKkQ1Qa
VQEPXgEL94VJlM6i2N1YYwaXOvaeSnTyaGSEAF9rOH9uQMx9gVWKKBSSUFQUbYHjx4Yh7/oJGKcD
XywCoG3PM7GUej4kXBgWrUXv1Obqwas0k8IYnkbPC3/+9FCHfRFaRdwdfl5RhSlAA3N3mDSe3tKg
S05DxENOyS9qTEkjNRQfVCkzSucYm+RWTrRz21h5oyBeyZR2xKjfnijO/FenstpiU3FSFlCRbw9b
qipLkouRx0pIWT/ReVwY2ruIQNrImbA9XfYusOCzhUyDCrJ92Z0ev+Dx60ALTLxpCHwHnG4T+rdi
HDKojmpNBuxNccXz2G4sHqGmuP6Hb143Z3M7cAhMjxxH9R1d0Mfpegk3gQ4zqNXiudmCqU44sw1D
2u29fyj9TKHTzFsNyRoKBuK3ZIjkLg2Wv0QdJRPEnrGYk+0AwcsrTd1CuAiE3gXpl4kikolakJAs
1J+iRdgH3IeDAEg+EI3c5pJEI9Yn4CPkfKRfjN02Nq+Rp2HjUUAsnOOktxbtQxUx1LtmjZzgl90G
/q6gHAq6O+Ochd6O8dZIQk3NwlmPI4bcl7UdoPdqLrUxnMI0MsBUdOeJRg35Cm36o0uEQRX3bDLv
aqDedAyDQ0qywSQgWC33V/sC+9xL7Yb3liKeAy7GPlMa2K7HuYREd8RAdwq9keVuM93KJ3LQJf/9
Syb1peNm+DRzSef0y2THZk71Svy4RepijGSm71DYRpjjPoIdrEh8w4H5Xzet9sBdr8S9F0RF1dFS
MibOYzjtjAmZyo53IK2n8XCqSY6IeBAwLMQ+du+JFStGXMkmBuRC9GcYBs/OJr8E6Ef9dCoAA/1w
8lOtEoSLMJI7ZRNpvu7ZozTLlIlBu6L2iy2vGwzErMUwJ7wrdT1AJFF/D6jW3nZjM8aIquklH3xI
rmQWdugWwb8xHHa49slO4jx21O6iTjV8Gb4MPZ+cbSHpp4rjVB2WpmQzvknk3cDzho+1y39RXkah
8LK/067eFMluTzAwtn389vKhyyRqEeovKKFo5wlDWPihhOuG767ATswqwym341XGIkXUkjMbLRKc
Ri874x2J+ugUVdiQSuzIuco677SB0ntIRft1Dt69gTWGqbkvLeimlycORIsMCQ9MMOUGr7KyOrnr
TeYsuWLtyN6+xmgNn+BaM1rx2SrRQzpzj8zcN/nws6jTYh8uBuQXhHKRRKBAlnpAIrMZrCEzDsco
/o0OQNnipeDgX1tJoDqaIFEHCrEIEcAypo5u8QmthBguHH1QmoDG0JoXQkicelsqbAysxQn60pR9
npZPkKhTtq9cFoKiJmPnk64mN2B8HC6PEwREd0tGxqBD2mHJVOoDjhb/BNLi15OEK4t/F2H3721E
71Jet/ZA0rpi68heRNhLNoBhmF2K9tMHjcwm+IBy/70xcs1oYMwn8LA215jVKIc7zn8ZZ1L6NKpj
I0avRT7i4n3oTIIlH2yVWEl+M0oLhAEafyjUXUmLqcz8v4Kii33bBthG6cF1GSXvvJUHIsUjuuep
d5T8Ft2Ix8giBCeCZ8Ko/yqnW8+3NJnVt4RGZNe/HCDutkGb7lTnmleTe6TRTb6Xqh5mSBzZG3Ii
mC+RyakDwDc/+1qL7FxG3nuK1hHUV1qYmpbOgtMGAZ1t6htYSyGtsBGY7dw0Tca7GvJBT5bkJJeP
LHmfWAZs/iJhZ5XdV9I1oXzD+AOUVmJCpmjUi7+GTGRWhjCvG3xUl3SOMmv5ks58/ztLuyOh2jbJ
31voshoc5guFCpbM2WXjWIHIOthuo5z2mOZTvZUkMQNavQlSV5HsjGoNt1g3S9tfZObSRwQzIT0k
NyUjzyRPUSyT4aYG9Cpef2LNy/4yd7Dxzq+jD7l3LSgbUngsgcv+L/C2wCZGugKIdg2ZCs6d+I3R
U3wrhi1l/XuU5rZp0yGFBYLcjErZBRsyH9U5urdKDl4UWfV4tZjUIERiqIttFpIHTjj5ct6QSqfg
QgOj7Zt/C42dQYqCDJX1mOy4DlMACghzIWoTs5tL/nfXB9z+nMHgLDkGFONWIbvaOQfeHhV/asHV
pdUrkQ6mndG7vOzWXvH/OkmLLCJh8ikCe291ljBv/Q/hWvaUDxfMBln0q1e6EKtlA3S3LSwYM9lb
MzSPkMPn+QtrwGpIqKHB4VBJhavD0sNXlwbyH+plK3pZJwTb5KtzZcYh0c2Il5zK83L7fqXo6UiT
9+7zQLXNXRHG7rzgY3kMQ7fFRSqGkTYGSxtKsimajPvH8ivNJmJHimIf41pAomlyS4dfc87iwsNS
hF9ad2VDNcx77+XMCLmteEYV0XLuVr78OzuVeedCf8T5hRTSnb/cWiG5jH6lzYENF+4qArnxw04M
I3HYtyQ5Yajm2RbIzniMU660Jce3a2zWc7pa6A/td6CyuWV3g9e3OUEb7YI35aOP+U2T3doE16FW
xQnOVcWgi9TG8coxHHwL5nkAmPhRKRQMu5tOsFY/VTKdc3arZ3Idztaeb6w+dzWdjKuXAcO7zgjG
rij29xh+CWkM6UE3m55KL/B52+h/rRfD0xeYUPyGUv1ojboF0Uu8JYd9T0m+z7C9KUAltRhJfmv0
CbNdB1sPiDEMYZgw+nNDIMP2w8JCE8NA3OVFG8Lk3dsQYhIxQbCcXLzI8b1STBOWs6kjGFP2iyXW
q63CIx3BsA/MAOw5X3svaKiYp3Bwy6OHLLLfoNikLfH20fbDkYGEEWIy2bkmn2V9A/SPkOlX3XM1
y2sUpcALJ9U+DAVvNEpewEgED0r0YsN7T8cWbnyvE/K7o1NSfGyM6ZqSlVnJutIIpBJqtYfUl/94
p1f4pxUKEDnZ/AQRVhtkZ0BisNCTA2wkzjCVK0zl2j46bwZkyVugFruTB/fHe+LoO15+rVRHbR9t
1dDOamWdFISYELdVlsawK1T9EDUl7RylDdWmun7i3sG96B6ENsjeuf+2XMYLOxABMuqX0/LlnNzz
CK2nXXnP9IyKwqJSJ1Z+U/c8yX8Gb3Lq2ZBKtajUkV3knDzNJwX3QRw6PjSMvZm9pUBOW+HOUkGA
TVv3+lucBlVPXcUO8xU/19hXYq0NiO8ev9ulViqzhb+8SFUmYAafhI0Pj45qSpi57NfX6Fqiw+c8
JyIvxpIq1LuJRpaxmGDAWA4jiP/FGmxP1CIbEws7X1L1798GY9C+6JpBnLM0D/EddhC8td0Yur4W
cikoCB0wQBsfb5RMoBhUrcZzAJe/KDuKcS0CgO8HSaH1wC5hITG7zdIK/vHkei2U9XBfoKObgFff
ULtiNqwK+fQKNSVqA0nUPnYax63zGVU77GVUGwZUVj52st2+SJqogA6ta/2wUBJyKeQeyQBFqPCP
YO1azTOCwpY97yHBoUN1288qGr1sIYnsmMe3jlQFCvMVUhc4Hidup+EyGo9aYzVoBQ7AiChcDF4W
Wfhee6AXdFRPdQRk69M8HiO0lBzXNkfYjyERrEi2SJ0OXaj669kcSdjmcIKpvsDfzdUPkhRtfdKb
M//jWln9IAvdapXle9C9XbJ4IOfTstcxzFM+VR0KSoN+PTSKThbovcIIlxdyqS2MZaohAN53IWHQ
5irrJNkJyGThtH4gA13zz9ZGvjmHm8lBsgtZcDMcnv6dLSP14rbWWyNCqJMlWuZQBY2CKqi40OqY
6sIad9UPt295spb6gKLW7w8DrVthXDEbAf0a5NWQmiFzEDHvga554i5j6Pa31NNlsY8j2NmV6FpK
0SslPGd0IlbO/XT3MZ2nVbdVHJylJUVgJbAJ2grh4eIFEjU45sdaIGWB5FLIdso/BkEn1CfjiJ0D
ZalzrKCDxe3I1ZNg49nA98f7PyXkdzgZTsswyziw+RD+JEhfbHyLrIyyaaMQaG3+Tfvh0PTwwxhs
fm7Rk2GYDQ4Mk4RGthgevr1y+8SJv17N3nXq1Hx2f92IapbL6qQ3kF+/iIHS0/vwRtUZn5hHwf5h
nnYBQwpW1cdnFyoCuK7+AV4+0v8TfVJxsre+usZxu9N2RLOrSTtLpnfrT0DnLuzaIcJQ91h/n/Zn
c6DtMpTZZWpnoQMyTEPh9NrKzNxnt04IdPpYBMANv+6gDZ3Q4Nagb9Rc3zR/lUpWotyuA6FjfmBF
lxM0rcKA1SUVrTUUQYrSfSPMEg2r5i5ebN9Zo5RLq+On21ceOdX+/H/mVvxtkJyDIBCwNZxO+NuW
yd5Rl5dV9mJCQDsdJ2RTD3U0zZ5klEZb4YyCYA9XxQEwQ6y//PlSTeLzw5DzOpK25JaeuhppHXgL
t6H4l2z8JNwJw/Hirv1kadG2837WC26kLTj/UUA9fvDqmyNO7lF5s9H6dqKMrG8Ck1UBMTP8Vhn4
1Dzoka4SaBAzbwrJYaF3kbXo9516/wtAOSCtjB+SYSHpfa6Yb1Yo3ZEOpkzEPewpfeu6dbMPFY4t
fijlRsA1Kkf2/r9zaIkFUXPehg1q7e5ayl6CmayqCLQeZyDmiPAx2CYQuDD/0FQQv8YU7YGv2ApS
u28ZgMeK6EutIQzWjqrV7b2S3F1xLpDoPX92xcW7FJOD0Bu2pd9OK4617nxa+YzFQqHNSAGbewZ4
zeRs+cSuFsOnO6DU6hEdZrKZk0zPHLMicp7HZse8ugnSACcnEiB/6CCEXoChsHJ0nMwV4LnPkX9Q
UoGMfGLDIuPMnXKNSSY9ELVq30AxrzH2GpxScQhWlOtQ1svzkTgXV33+7asYxzc9OH0Vh3ia9yUA
w5smIUVNPNpb35B23eF1uUaOy+CzcoMnqz6XF01Tv0Z6l50slyWLHsgs6A5HNp1mPYbl43brSiuP
rSRCzhxtutCpNsaFLrD7FnHu80vesHkNNv8GGSW2GAS6uxFXdbfSWHOADXZwFRKquK0bFUZBuPEz
DR83xO6Ovk/9mA5KP31jyRGDvNoHGXnLImLTdHZYbgCViWAbtL3JgEvzuDlpEGfzqWKXsN/TxFrD
2e1RmL9z9dJBG9CIsfyKIGFx2X2XOIsIh9vw16OAuIEnzyFud1DTmSMLmiomu8DlMbmqHvQXrajR
mqwmPEGMTbRJytOQ1+evyjUkWzCjT/fWbp62CylqBglmwNhD4yOoz0gsD81gKRjOmMQ09Msipglk
0Jw6TWqvYi31JYopJnwDq+j55xhPdGxnpWiABUAmpw4Rq38kZ4nVBuH3pdTcbitVd0sDhAnFibEu
6gsKiGYHTscQnAaHVr65hrNN6EkAPP3GZ9nrxdat8lr2rvIHbqHfW02yBDYrvOH/C+9yIDbV3Q6z
4Ma7jX8RuG/JzcwCshrxM71W3pE7rN/SzeTZF+HUqO7XPqTInkpUcqVAAt9q6XThpL2aqtvW6wFU
Kl3/AyhV2AQHUZ7/hTkBnrVMg8IhCe1CUzhP9pilMt0JvE5Rl//FPDdw6Qm/whJ79xhQsj1ZhHvB
GbM6Vld0xtDvCy02HxR0Bo/LOuZ+xFQurjWacynYMW6sM3Fkfk84fjuiay7A3oDee7PyXqszImim
rrNZI9cyKCgTS4oNO+LRq8fezYRG45/YAjUONJewH2qJEff198sFDZxUY3IYEaf1Kx/AV7DwAtdq
doQa4EyXShCgAiijZu7umQtn39nWgZboAcLib95+qBKvPCrv8FiFny9bY33nEfCavkVFFJfFkS3w
jmzBKlqJvKkUfPmcFHcX2nSYvOTFlcGtZzuQUSYnQwUhkJYjNl9agYxOfS0tHWRWccEZrXe+1f4n
F+OLpT4AYPMknJGnOM2qBs3qXTgCcJd5BQUOXJzHMspyE6I/4jORHmuDUR6W+hkN7z+cKOaHYx6p
zffoBKqTE3veqTOxqfCqPG0iHcDoBacbymQRiZkQ4j2NNyA3v2ESq3NtH/Hqqg/+QwwHZjUmOF+i
nUia8jxY1CmVum1cwDhWFSDkYc8szPqO+lTvKqEyTgQc9OMFdLZ/jdzx03r6euUb8HY+NhsP2UNT
3ev4wz8sdaSVVO7rrpqHf7PCWfAhd9FkVKiv6NF23Vbas8SNcY1YyEXT0J3hOOfhfEHCskrOWPHQ
2bgEvIlAyfuPLsYnq11O2d0JDAY7lCitm1SCkAMDC/Jkn5PxiWTaWgzhzn7v03WWT707Fl+x2aNv
LcVyiKaoiUj2NP6sASE3/pZGmIwtArp/N41cWTe92ulf45t4JIeN6TKD23ArJ9Hgiqb3s4eHWTpU
YDCMdSpecbMXK+gqozFDpCsy9ki1/XxCiiNg/YsNUpR6p3Qdm4JLy1McdgqVQcXW8+Is9ARxqqgJ
hsHJi1P/h8JIRdTQVfkg5n60Gjof9hOhXBV8Yvbpr1J1fF+Qxms7WUoLM5ABUn8GxCQ6uJBunPU/
piGoyvJamJKQril9LPFLUexijqPG3Hw+xdFoNEQj5L4o6+Cp9j0geIrve9wMTOWrT9dtco1mb94u
jNlziVwv6PoSh8w+OXy2OwDiR6vYQ+TE1l9gmSyk6INlkJk5cfeaJSBd7Mp69Tpsa52Oj5vpYLyQ
20nk6qJ6L85iHQCHzWwgon6XZeJo2ophVNwjvSjy0yIE9SWPGLptMrbNEjOjW+PVoo53iy4rzuvM
MWq7Mwrjvqi0tKwCnClV/A6G/dxcRFcgc27Rco2IWWlyxlf/nC5wo9o/P61IZ2IRXxcFfOsvQKbX
twGqhrXwMuFWcuDYeSHSGDXaupg9QLTN2P259R9tp4jQ9ZEvH6R2dmtyxI/sfl6vX8KK3sE0g6ql
BKwh9OB9vMdJkYYYsy9xxyHMozm0ToVx95KOyw2gugs2RTQ/1iOmQF5r5h3tci2Zyi95Y4Q4mJN1
5eutNspcH8TvqSE/Rp3RlPPh7eGGvQMAp5UEOGLUekfGwVoe2AiPg/OugR1xhjKXMT2zRzPbJwu/
oqb1ZMHBOoaC9xbIDpbzw9TA1yTUhiirxX1TLHuY9rElVuJJPGJPD6E+6oSQWapid72CgTIIL8vi
UTfZbKrAMjZpOae24vTPyqGnhwIkym392lxWbHN+uRdWSApKQbDMH7if09+ZpSKH8ncxq6PMqTpG
jpYPrD59WAT4Xg2YLqAV7sfGQh2YJMPLZfmEwE3iN98Dt+0Rn5HXxtSRsRJyvu+EK4FCAxTQqJbT
8LqgOOlqD1VSzBE5Ufb080p8tIl5EJwvTxMJ/65ntAG8b1jJFLW7seU2oGfeE4nFhfCd5TtzZLFf
cxciQCWb9TXjx1SpV/hz0gZqoiMpIQvr8kO3VnmanEwaxd0++kIzWWJPsGuQQBlfZx97Et0zyQkt
+sLAd3fyl+LDvgzUskZFZesuEv9WhxCCOQ04x27CMJSXv4MLC8KaEABMaORQhzxiUN89e4SMLgY5
LtBZ4j+Uywh3o92nF+apBaEDjt5AD3Y2gHzX9+4Iwb1w8gcAuW36L+qwCygOKyvoi7qFSHQyAry3
o7Yv9nhEqqrCghX8wFN9OaKQzPpjdGnn9eRNk63cfcmcibdTvCszid+ia/KxscjPZvEKhNqsyY08
mUfYa4NFuWNPFXhG0zIRdrtuehjZVlwYkedR5LZs37yfJWHsXafN4kyES3iv6OrHlaNzIRAvQTOT
VwiWCrsVrrVJDu087Xr4yRGQTHcxcY0DiY5uKHI5IiNEKpOR6b2uM8gC17093hFZ+7Bes1vrmuI3
NJT1r9bxnhkqAIu7Ydg6yDh4XM6/mPSldvt1lHOjxSiC5m9+VqM8Q7fLzOrUGcwWPY3Hk1xwtGEK
yvIVvNLD8LRLDIyajdchLqscPYvo4Mvwp3QZj5EGLrCLy29P8PA/ZczTqOf35EkAvkjeQVajZ9V6
wzjuV4Bahco+/hLXGfVsdLkELryPP8Fe1hlahfb4SQEq+VPs1eOoLrrRaEyg47wm0o9YAmmqXsly
1FR7VuUWCSla6BL7p8AAZabRhRPjWMbkNomCKfmCdeZj2cy7+dhStxbCwwkCdgtP770Ob0WdjanQ
inxMh9QMO0V6viCbc48pG2rXLGPp+73Eh91mh3rn+D971ndcM1d+cvaxYKEqKV9pxVI2GSnw7flA
TO/lJvcELNn6dG8hBpQGr1l/uJ5sRrDVe2wDMeAuWX9RY7uDngavqE3AhTQiw62AvOcaDLc/2/5D
/WDBBY35DQu9gKJnG9J+U5+2wcOhgHqnctyyMYxb5ibZuLwkx41OkwoU+DZXJfikSvZCaS6Ul6xW
LtteBBGlSK9ZRHXPAaBSxp0bFFy8kYjWWLDbAMjQbVnCaGT7D2hvqaX0Lbl+cyEhSEzzSPNfX82U
lgJds0efznAB+yKd1EWsLqAFG+xKZ3IbO/Ky0Q7mpmG/20jccaYvXEE19sIIScYjhlrZLim75zcR
vsdSGb3f7WcLvossiWno7BrxfxH+2nWPQBjNG32YXfC/W5IyU5xSFT3S8oWzB1MIwu6K0Nlyxp93
k1LLnfsl8LA2nNh5IFW2Vv73oqZlID0STymOGRwtIQgQa4BSz77KrA5kes6TCdmUAAqi2twLF/CO
wfYYW3RG//4genmzhJHhbIom82PJvfIiqTXAta6gMejqm/7vdrzOtlbxiLYJ0YCBTCsl9Y7uwKZS
kOZuZ2ft7o95N6AQjM1i1irv7ywMUP07+cuLulm/LI5+m1Zn/l3xd4n6tGzGib8tscmx7R4GYXv4
FNiEylpjQNKZsn1/0Ir20mJdfVRVLtdBd8Q/D9gypjedT+ryWnHcCnmT0t9iH5rNUyCi3iVSIjz5
1xaPwtlIehYPwiQo6G55mmmLm0CVIpXqByWxp0sm/aXtDXcr8IWO0hZht+tOlA72QYFCDeSiUaXt
9bjI88NnkahMotT/q11mKz66XAuDJe/4jJMjlZVhCj4U2xT1GS8fTCCF/0Rwk+wYHuSMP/t8rP5k
HnED88VYz7PxyA0QJIqFrp3FWedE/hs22h6A8A9M5pcORc0GEBZep1I84PAB6uvcRyK9Y8gXBJXJ
M5UGY/SjTZ3fxH4eTyim79xynYCf83VtZJ1h0+w+Iqv/0U6+nUzqldwN6R9KK6vTZ6vjBXoRwBqG
9/owqnaOunaLEJdlig2BPFcHe49m8xFyhQfC/D6aMTQt+NM76xLIiF+GZfQBoQKvkfl4nlkE08jE
0ErvFhLqmsj9iufNXSCiNIUc9makvlaVWxjVeamIt2s+sJ3ussP8IcYnDoUK/iXDOcEC/bhoT/2d
NwC5W4QCoyQlwOMMnyxMDE8DL76XCbtmRVW2ObTcOqQWMXqc2wNL9tipeK8ot6LgqPOs3EbnSnXK
Rmt/MLqbjC+iGuKAbjSVZDugGhEGdkuhEYHlyOIP99XTg6P6lfZgB3A89hvKkAM/UglSgAYzIyl5
dqBNz8H+PM6YF1p6O8ELoekhBpC0XONKKnboa2t1ouDPQmpPgH7Qznun5zOUR/22fBzXHrSZpSmE
fVhNZf7P+SonRHq7iepW5YKt3j8NE547+LsIIof2o1tIerPAxAHibrFizkn+5F3WlsarAh6xVSRY
WBNztinu2ijQpDw375G4oJOp0D0Hcf0boNhvxIYgjpj5z67rhaoWF0+ZvM8qcg8ccu5VXcXCZATY
ckg34O7LLzEHu0pRTHaPwrhXlV+m9aQniRVFRevB85/fHN75Xa2SKBDhAut3vrH3NexlnQlMdF9G
qZITkjyDWSXhzf+792XVePOnB6FXUGDba1yrQhXg64rsDWlufswIrpMf86TqNBRWRRVxv9CwwZby
FmVQt+xPfxihkTRJNK/c8OaeYhTkW/Bo55ZPVnJdWsewDiUDTgZDUtQjORrOW3bO9HU52QbCL62z
0fq2auV3ApLjXA72n0BSgmssQ0TaI+teLIsoI74UqY4IHYfbB8ufXjgm94K++oEUEX2OyhwqUhXu
nJ9dZ6JLQYgDD6AgNGGvXWhZw6b0Q2Nqzwje74W+GTtV6mjX4DFsb5y8wuyc51G8WxLipHGZONKV
BdNmxIYtwm3gAZF16cZK00h3D7vQhmgx+xK47VX5CL+2aAwC1t7rUQDynnDGGzcMXyq7xj87c15M
YHT17TQBR6yEtg7hSpyDMppDynXWMH1WDWDln/XZ714XY4+D2KnNN0bN6ii9yJxJobvZbCHb9Tn6
DeBeSddlBRe3W5UPHbVm8iG6Xhktt1qvG+2W3L/5AD85aCopeCVoVHjrdeRfC4hWxmOj5ezUf/X2
oGClLk/AGYLkkkHpfXbDRxVHDXlNZ7B2QgD4cw5hbRnbw+LuWSJkYoRGz83Bw0HXO7X5TIqKeuYo
wfKdlDUWbwtjOtcUKq9A7HV9EBJN8078jDmfXNysXJg2tNaj+IsuJw38oZR2NqPF0GK/+nQtLEZH
Hw/0eVd3RSKB7EV3D9f99QLR248eVEx4htgPM7nt5W01uugwpI5/PKEjWyLQ5M8L/xNNUAZZ4r4j
+xnKsCCuNnFjsOS3B4Q12Z6rEK11sulzS36J4ihwGSIzbPnTMu6yMZMbrKxvx8mbsTPcxjRXKFNA
P9gOSnnOg6avlCLWSSmOf2rhLvKalszUbBfwWUPNn6QGj6ZiSOwLTP0JhBSoVff4ga8C687wicYJ
tEiI9D86E71M2PNq3SkH8T4qHc/5e5FaNUeTTbtKYInV4ne2Xp3YsayPxt3lSH35+6oELfr5d6Rb
znbS+cM3s5Dzx/G+yayOH5auKqsjoT6yHMtQpdYpECIeqiiOh8KMICgdba2MIBFjAhp5fWppuDQf
199OUQpiZAjQUn3neDlTZGm5L2r2dU1moAB7u3Y68Ee90Qe7e60SeiecSvHjdX6WRWnME0s6IU/+
bS93oc/s43HEhjZ7+UVopBckyy6bpsC6FoDbkMME97EXlYJ0MFZIyW4kUfNqF3GShdapfY2MWPPc
HLAJtg/trloTbI/FPC/YrTDKzOPhV7D1ISlcq6foug0vm9ezIvTsbD+aOPNIPLFs/SeUtrljt08L
hymkSWe9HRY4qTGIZgeOJFHOztfDUodQnPZ0ej1h7Vy52TjITwPin7Ygr3YQIQrAiNS+wBF2cgzi
QDAC8yKoVdPkiqY0gPzqt0i1xFTzXkBgGK9MN09W93HlxqOzGUHNUbpgH5k7o2PZYYq8icBwfO1I
iDJHVbNTogZ2ddwdU4nN2KasYBN/2cB9Y6i6Sd5Oylxa1UNc+O/G8QdPkwZ1ICrIY16MKqg6MPMw
raLTH5DHIcGF85noSki7O+SwvbIHSBDxhwGX1yXrP2Ke7qhhu+KDBhJh0Jb8aAd9Mxxfb0yFkXzO
N4SRrDQSMKQfaRmAc0TJ9AxtuT+cl+XMGS6GHrUGo1JmRQXcYFey/JS8n4h8xZRRVmxpyIvEX+vx
/GLhrFRBLyb/RhXefNzrElbLRydO6Ovuxmu0lfN95yioTXeTkBb+wT2QNQ5CtzhiIx7DwBwwjaPV
LHF4Q/IfTerD7lYqaBdIEYPGMjrhZzG4KzKfXjLK0Vk7Zh70HM2V+mCdu4SJVv5xkdmy6SSHw9SQ
edbM9J7bAkEQicB8sEZ4WSYVIdjFegrmAlhnOJ0wwMogET7btUlUtGrLhFDasRu44CKNr+ce9sCf
0xsSf3YBpihGMs9wdh9CjExIJV4mnssAB8s+vsVnkYmp0pMxaLSoDh4m2jGoJyvuqYU85orIu4bE
J6HAQ8FB7O6vw33cMusTPdmFR1GtRM/lXcZwslYc3miTD3tuj4JBSafNoejgMuZQXR8aBaoPv9Vw
or2EktKzMeQ4v4ht3B05VqPKPAMCTvlbIUcQ8A7nHFyDY/VWKS4DKaFspJ3QaGAHdNuodDcFRmpm
HrahaGRfgdqmAixJH76o45e/Ouzo/dWxXUorFk/jFRqY6wED5bz+rDVr7Lm4z8IPJovoKQotfy8l
feJgT8I0YIWmiPgAPXsR0QdJfBg+6sTGZodtEydlNbznZfHSK37XiMLQcQucxz6GhmMhwY79rSAz
sxpAno2qOJuIBiSJgc9aNYnTIv5CCNftdpKQovXyzWaLWB5lU3k0YVdsFQIPiJoDs8x1qVqhqgLM
mjoDV9xxEdnWC8l3RNnETfAk2MJPHImoxGbSF+Ohk+M06wV6aaM1Csa9Cml86wVk6f2toWc/E6oN
PyrtxgAua32JzykIiQJnfOYVc4cHMIJwm5WZSlAX4khXwh8e5CvyKIXi3PxJe3IDaGUCldqcki4U
hn4hlQLEQv7DvwuAF8eqsx9OuwXqeBCbeYLtJhrk//AbxjhXzJ3VxXnaC8Hi/28mGNcR+l9VsPoB
TyTGaXHlv7H+C69y/XkDOH3U8iNZQnw2f2D4ppQqZHCu10YYA1iDrNNoSIyTNd+oJ7roslPCRpd6
R6GlLhfMMTr0+D/B/q0fU77WP2bJzF2vVgXSIdxdVv+GPnv6XqKdXqVU+y8X+AmXsOAS+Sul5sxg
SxiEVjKnBq2ur6+JNPo/roOUAtWca3K6CvukCAPmOluDba+Xa7JgHj8PXi3uFa7vnBmMq33Et4M2
G6dBs/XSBvzlAku1oGYkitD7WQGRtXaMXATR/VRstXS6fM4NjdZBKZV3qeExp4RP9swjwvZYS5++
/wQ+4rtt2rnxCxmyVj5AjkNBDs6iqkDsAD/Jl/s1st8jOXZaRQ4tehXsTfoQJI7RuGrvs4nE00EQ
9B3Z2zGW4ax0fO3qX/Uzg/b02sVr5h5nU0u9ygBegzkRiNqC9qg23k0plf56XUCR3vemS5y1ObqU
jFVXmFF/yAayiW4LzXYFEQ4J1BQU4jWaBk17TnjP1gijqGiLxg2MJ62pFEPx97oT9mIkHIppK/FG
xFtDGIDI6jCbeFuz0YFRwwId7ymMgQowoKtmbEfnr2/pHJGJdHn4cq8+LUJ4vscBOg5h+yY9D3Ta
4VD++3OPK3eCzwFt5HCyGaS2GwEuagEhCWbDmuJ1FjpR/A1gU7cR1ear3v8MW7U33hj2LGQ0Onej
zRmUIYfuBUs3lmAwytTSRVB3sFlQabF+dxc3evuhvq4QnZPlMBzlBEo0bkRMNdf5O4DS2csfo5O7
iAK7V8RTb1zLoDyCsUAXjq1R17pQJhFjwYFIo9a17EnkAOA557Wju6btu84EhzGkactDisp09wIn
1AapY3DICyCqHdWyt02GxZnZWoyKyexPI4qvxnJUgMtVzEv04IvtYf53IipRSNJnKKXoR3vXVwfq
LH9GAM/ZqiMz39stheVu8bAvsviJfnB18HOrAak3TDrXHFk3ysSL1OI4ujyfrMAz5fxtvzHjaAAg
ZtQ6RiSoK2KI9NcgqqOuWxr11Uly+1h2cvFBs1p2in8z3/ucuytLcpLCjSohtBBakPhzuubon9zA
BYnA0Vt/+xmoAFQCKZ1b1vUEXtIUC/uIpfbHRbvaC+k9YgkRvKSlU3tPONGU8p1nDDXh5t99KF+i
+rq2vaICgx6iUI6/wI8mnPMsReWBPFhsf/qa9PFnsR267RyJxX9YABC9z2jfWkIF4viZo5cpsF/d
e6saEEArjgl3SJr3Z+oivKvwgqQQfyqKFtfEpt6OlYGsX1y73ebsF9nAzjUzkvLtnRMUFn0kfHuY
NRrtZ0uG7O+6i+Gr6KH9pqvUyC6q/FPoEQb4u8IgKupshnykFLaLJC0VLWquaABIS52i/XS0W8Vw
3zCiJRsmh0YQ+5vmdpLJk2apcK0/ASY1Idcn+PmTNIaxzVA317VQmh/McSKG1Qh7qG4baZiYgPDf
2iGcce7vnhPHLXbwXPbYH//Oxr25qaENk3PV3eciD0hQKMbQC1/dq3FN5YXgnfg0RI4P40d8WOJT
+cnqbNVVL8aQZTsrXjPbKL09vXyLbl6HfRkSRmdj5mR1xAtZR4U2J0glxUZ1Te63w5Y04gpTVbqk
km6eS+zOpYnxGYF+z7zaCSAi8/VwBz2Rz5f/ILzhZlpcuGf4YTZm1w142reTgxrx9zlM4mACCWNw
tuBoNdFg8kH302PrC7DXrygiGO30JCbucybIhWn2yTw5dYO5Al/ytI8qec3eHLVSbwaGqoFFGLHo
MynxTQS5Z14PuAQsp+Fkfkazg0SdCDXKOYaORlJz+DTurF8VNVREP3d0ethecci5EO6CqxGc8xHo
VBSuW0NWR/MZiRf4gpu19CagDLKd6eE5C8w4IClj8uZ9jO9vqwAn8MYRCBgOs6synevTZjo6Sm6N
n2ueT73mBYg+evfLmkNT93CyjOmAcKbw5waMG+55UIZb7z5W9UXsUumaNY+WTfMwxDyBHxIYgRjy
hfmnXWAYVjtc4M807DQ28EuxgfvBZzX+ZFFzw4DjdUtbhTd7z76a+qt9bHzNah7UwLn5c/XA+lvB
dNZSLrNGjKVbQ3g7JKiQH+MOKUjbPhw3MFEVh7U/Na1mc0QGUBI9e7gcngFPdBsZ/TGPazH4n4BM
autPr0RNQc/WqlGnysaIP19F3vXB0A8K2+4nmyORRdwNtjeIxrNoW0GCkOPgpEc7Js46msRM2egS
TrFxZfRt56R8B3fZntDsWRqsPRlkqDP/ZkVyoK0sJvYExuEZa0l4Qtb8bnRKNOY4lWykysJ1+LAy
mJ7Be+AA2HbXVk0xa5vfqs0XUWoxifbt0Gsrc1furJOlxig+z203HOQPX9bIoZT58oCGap2zc+kU
C8Muz9gEFv4kgUTUrIpOkLNRm5SpM+9r4j1U9yPiTMwHUet94oyJxWPj5ciyi2OsnprC/GfvCTlV
E79YUfORlbOdcfDZAS0cxclqOFrgbJcBPVtou0IqI/kgvUJrMvXXndhiIpJN3tfprY4qUEwUoQi0
mHL8KKCvsWv05xuyUCBppMAPb7OpQabGItm/jtA1AMbq8Z1fgtjcg0Ev37448ro6oTAbcyPFBnp7
XKQqjfFmbFmFnLFAO329Ter/f8wQdqdHqzubBtM+9MY+cMdCJAivCy9q2nVSVmSk6SqnpU4jIWXj
1fpWwwCgM1UPBgziA28mz1jzEY/jUcPg24FPfsmhJNSB2GOKNrB2fl1xusmbY5DDnuuBm4VUODNS
o4zz4/+DVimvsMovHMqPNuyEfHh0RhL4a0XuCw+bMI0wGqv9TY4qfX2HMX327YVGUkhIPI5zlFnl
Abbrw5VeLuOytHxNUQq7IxFrWUh5XjL22FNaO7SY0xyGc0C+aw82vo8SekSGc27lufWYc201c+ar
UrgQeqf+6ZKqffX6k6IFcmLhegeG+t9ADTFdg37pKiC3frJc7t2U5vPbtGWbVS6UFAngPe+cUgkX
a2KadD0JH++qaPsJCFRoA9wKKdiHdmLzSqs8qpjPhA9isdPaRNJ+XeSIlyykx04wZvsIyRiYP9wA
sEx6i5swNRLu4j1j+YdU/9sOYtWHTVtU3DXqdF9OT5YpVKLk4OA+yQAI4hs8JtD+jIJYRdfd+/oI
puo0B/zsV84b1fx96XPkOGLLOciVSdCFWLtu9WrB3GZm5FxFgABIWfOXn1SZxR3YTX+rcwHgRqVC
HlH+dJCcLUjvENGRujiEJvAxiEnJIwvOvIE1n/XqDstGZB55HYBWdI/RZWsiSiDPZcyHnebHvyq3
/AmyFreNDM6/PTT7JZ4E0+ToaFehgTSvWEIQ5yPnpxiPkLbpC5JrRTCiU9raxkVZIe8znHOkxjxh
ZW7mYzNcOzJwkCUh47pynnDec4qDhzQpmBHMSU+XrF4MKCGd+8PHrEkZk7/p5Z/H2wISiDZDfVAi
vVWkfZKZtIfEw/Zo8lmvbhfXP+uyBoUY06+izcarkcJVEgvweGhTvhyt6M1fe1gIWdQ2j+gnx7u4
8wy5RcCT/79Gvu3StI/mugO2eF7XwOfPs0OwqFtL8zVIj7jJyZMy6KqAau0fryYpx9KYYSQsqCza
rGmw+PTTYAuBYSS0RGlxhdJISzqQ+JGXip1PeEpvx5lt9E+GU4BOgiw7NLcYJmyntY3//oGDIsM4
K2kj2HrHgoqUGJgz3DKnUjVKd1S9ZHqalV7+GAv2Bx8c4fI+/JNU+vZgQj8v58BwK7cIUt1cpOgB
CGH5qJrNxCPzaxSqKr1N6Lqyz9DoDtYzuo38M4c2Bq8js2OMZZ72H1ucNj/zALHCGXOgKmkyFctY
d+JJz+LN0HccpZOJOyoNTbLeoIP0lbt51DhsthWIkLBm3v07Q8kyNziT495Pzwn2QUlvCbyFnEp6
qmSAlW0V2VWcSsOqEwtIIYXSvaqipiGsqgYPgeiCusV0tSGJzmUaoC80Ak0wVdN+MC13Ccq7Qdb5
64ftsmLfn/NN/kII072eTyTORbUI4Zf9yxlUAs4BSvBbTDjAbDXeit3wcO073r8TmQqiWBHJFFsj
LdZg+Dq8wz0uOWJMamryAn7RuNaOr0FPuscCEo21V/dC2+G534Y53CvoL/Kkqmumx3IOShbVS6L4
fwtDkzQ5eEqWvYSAv81qS9lTjaZL5puyAxnUCAOyC+vLtxqAIKMNsMLgHP1YLZGhLGofl49hGD6U
v2+IxArf9pEAmTfzixK78YUbkfxKtEx8ZBaDDI0oeeLJQzTShZDNY+JxVBNeChoLOcN609GTPKqz
dSu96huOjJnGxg7nSNP5OYy7HfA7BNvIIH+VmFDNUE1wbeg/LLXi4F6g2miExyMKHYAM6zk49DSH
lLPmVKNEsCH67NvEtWcfXuwacCkKCBYL60M4GPEQiWfNFwynHC4dPtSdqRpURhz5BmwlfU/bpNw4
iSmmaG9p6epRM/yFq3TevOB7mVL+egYZMreu42LW4mSFazyw9IzQ2BP66jogKu5SFIWcpdGKxCMl
fM11eeJZ/eDAWpmSl/xgiLRVULnkN4fyYZj46WcU0OdWThbV9JKyroHHVKg4KYm7sTJEg4YSN8F1
vbevhsIIQfPEFJZBbXcvvbR5/d/+1rQ33QuYESSj037+lAn4A9UBrxM30RzVbr4ZJfj1nXxbe4i6
GezQZMSppaSU8qd9bSaxXDAAN/Um9rID/dUWkKq3lA0FkYuOxwyXW+U0BiihTRpnaJWCOIUWaU/W
p+52h9l940v30HicWL4MCBY25zeEP0gE7ywJ57wPqUaOLWIWbLQ+AwdtyaxFp9EcNNVdI9qga62r
0FuFqDUCgYrUGJNuAImjJEEnUYQv8u4cNFt7KuIScejYhi1wrM0sh4Xa6mjkoays3aZwt9TWOZF0
/2CkB6HGvltUchtkisR0NOPWsvcYh/HUllEgHoiYXsf/sgg68q6RLd8yRsMXI6m/iAfm2LCBc99x
nmkHE3cmarjiBkhQcc0Usfh1LaSeHTGM3roYRCu0X7/t8COZqUcf9Ag4aJbwZiQHBTRWs6ctgVJN
0NVH+PEj2Syc8bd1fjru/AwGf3DHEE1M2ntpL5xf4ja++RBNewfrqLyQoceh66iBz3i3gqFI7oI3
PqdpNdXpmc63UBO4dq21p7oqUXiPiPveMPs8kDVuWnZ6Q1ezqljJZLyK1KFXaONJRWq+tFlCdFj2
AXmqTfOrMyVcaH4bjXSaQtMenTEAi7/DdHMl6fbjT2MvXQP8nFcQIJdk+ssjcJAXRpknEt3B9LpN
CH5X1Ktw8Blsc3+X2V94sqjvr1RPfmIG//mcq90euttBegFAxEbT6w7lsl2BS0Pv/U7HnR5yRBeY
WAT+I/uk1/7JdtsPdTiJG3LviGCQOCDCImbrDxV0bvEPr4MR+LwCKmzXv2NwxJlmpnSSaAy9j+x4
pM/NuOQbAjOCI4FgrW6XKVS+NS3PCjkynA6DeFWl4xNAIlfmUnTqvlgcGGOqv6YqjbATCcmDHD0F
NtmRLEtWSL6nTa8AHTOV9BE03TtLVWlvxiZlT5kIEiG9/kwqbhnAjuPqM1lwm9uLUc0uoGmdKGgC
HWzhpkjNmOJJH338xmLIYOyw2uCldbagsTSjOPVI2u2LNDatFypanv2tkp2e7tUFss27kkW4bO4n
3TWNml6kvdmDQArSRRrhtmG5pHU3tMjL2JXAF/RxWHfs8CSowEviOhmGEZhusf4X+qa157JRYlK/
5xxh/s8WNYr08ct6o7SGXtiJ78WnlZLtrDnvD5JtLkuAhBOrOdidlJb74EoKHG8Qu9HJ7G9OZycV
s1r3Ud8cjZvsDI63Kv9I4EJsAgNom6DAhmefQ8QYUPP+eKmUN/E7RS+XTiUyxWXO1USYaUCVYyq+
3SUspzqW/t9ktWFJqF4oJcd3PD1r7V2qCzppF91ZxOj2GAwO0oaxSaE/S6xHKYVDyVHBFkUq5P1q
UiJ9tMajxVEIZHKrSDT/MKHeljeZHCiINPsgBIgI8N1o1sjB61d30PKKUmNAgJ1HTUTVNo7M8lz1
tPNbaBUytWjmmD2UubHsOl02bZHS5N01BxO0UhaabnNfqC8v7JorLyZd0+Qit8n1X5LgJQBFo+TX
yqns7H0lREAuVfpX4+CBQNLrweDxB4OUpUrsG0VF1xXVnWZ3aJgPS0+5ExYtcoumtSUXSODrMtQ2
gY4WHnSgDZf1eVH9E5a7kcFo6EDX/QACrJ+fuUi37HhcFyXIsFfiaZwnD+KMmYW9VphU2oewYVor
i/6Ima8cCykd6wKFVR1utrbm5zzViyuAUYxQtEYiFR4bTfzStuLvAypGEl4p4kxmoHeJRNIS0EAN
UjT6BN4fGK2y4d9moJbWeTlF0qZZ721aSvO/9Gv7S90Me/hJSsY01D9yQaUyNYfA+xZbaRfbjUEf
vOsZ5QA6UY/GK6YhX6W2d5S94wtQhB73wwRBTVeLTZwQaafHWBW1GJ63+iW8XWZk/7GqbFKcOgI+
Gf+ELCorgoSKGQCYUzq/hwgahAY+Dz9LbCvFAPyymcwt8QBhs/bT4sJyb26GpRNrFh0P+sNeq0Mq
jybeg3qsYlKqkgRy366sPM6IQSb6ixCPdYwgKmgjxIj6hpSx74587PCGr/tAbufkpkuiDQOsoqjZ
saCJTIqNIc1F3S1Em3xZqrY5Wsptk4ypohVDPR1xYOXiOV8e31/hLLpXLeByvcBU9arQWypaFhNX
/VHOYFRlbCmgQNCIa5tHj8/OmjwV6urJ/1vrWBw+8ZfWEu3KVubKsn6QgQ88j97VvS77/fE/8Kwq
zEaQ7KIHJvlkKcrY2Dq0fcw7cHpYCFzelOAA2j8IPBaMl9ejQU8WYuWnjEvN/V/OKxX4vyyPuTtd
0p3894f5r9m1sk54RByxKkreATQ/4VJE2dmK+lP4lVLvEBlxNogv0/62GLgIoCg68T+58r82JQ3l
GT9kNQQGNsgnVXzWqbqskKSZCASSkNXF/e5BS3l1UgpKjS5dWRe6O+bY8iK+bfpYFwB61a6xRBUi
UnPhaPA8Ki994CbbK83RyJ4HHtnQoO84XCvzF/UPvVJ1T13hlHqkrJG4H1CHmNKMs5UpFx5Fo7+j
nE3kTrqbwPtmkK7sTxHtmrhFVUm/ziKlEdNAMdsWHriOddDCS/8Zel2IPpX2K+ev11iiwEzYRwgo
mSLSDF++T7jv37ydwi84+epqs7LbHqsxL6hmqEOmEwfzkL3gwN710w02eMUapZ0XqwJaFUAn3YQy
KMN3BUooZynQ+KnWjCkXplkriT8D0M6DcaanADKDrD/lczTRPvUef6kMNpXT3Qbv56UjhqnUOZqx
MC8BTPdaqFdOQQvHRPE1KyniiAav4yw8JUf+u6P3/YycuLjzSYGZWFFDgPBQz5WNCzSMSYfthUm5
n1mll57Tzc7L291MwEVcP2p64UdurRVM9Dxkqo3Zezwc7K0n2ibqUd8y4sGaUO8qTg3Expk2aN/g
YSF9SzasCMdmhAFPOq+XqMTFuo7uQjijwQxNX33XZUmwE+41Ts59oFyl75xE7ohfemUjAk6KKsis
Wmo99Vk8Juuy/3LKk301bwcX2uaMKl+EKTXUCKM8suIRSuA7+4PUuvTFp02j218feUN9lrVWpU+n
Bk/yQ1tGbtwnHZUue0BUUgtn6pagBCW8YkBaoDVtzu485SAcIhruBev8mTjimNAy6lKQ4QB3nxJg
HaQQ0AsrbenY3kpkUwpBncBSOAGFg8U98GJ6rtb+GQ0s4Mpm9c7+wJGaq06I4H2z2ItVY5xJdc6w
3i8b4pSGmo/BuNq9+/VdLjRhUSU5TXdC0EuQ4ECf/Q2in5Ve7ss7ef/TMxl8HPeEipVAAJwuxV7o
mnxdAMnGz2bke9jGQv56k/NEgqsJvKhipM+nJqW2rjdDgNyRMCL8gp62tqWXBbi1vK/J24KWhY8q
wCqtHfko36m3IPca8RyM84+cysxJU9Z/1v090Zy+sCsxTu/+ntln8STZl2+COm9xkV8HbXMZPX/W
qAJZby0BTqf1YyefV8AOhtS16e5VKGvExM5x82M0uF+TC0rnfDKibM/QLAVIi55SecAJqQrX4PSU
UNG1HYFLw8RpA8tHveIle8BncNnhqc5z6SmD8H2TQlWkYBWlEXbVhrIVVipbQirqtRQwKqZT9D3v
Chl6n4bTCWZ1viPxdPIIOnSmo+oqr3ptPiJOA8bp6UiVq3zLtatEChwY3CMGAI67kWMvdG0D4Neo
OUDlQ0D+4hKaD0f71vC3QmIWbrsU9q133FsqnRsfCZmwX0H08dbC5VkN9o/snB70oVcJl7Dno2vQ
RaLKJo3s4tkP4tnv5eGA79cQC3nMUApBoVtuLAjP85IaO+NC6l/EMSPf9gVn+uGNiCaAQlcNGy/q
sa1AtMkJG52CyBn6bghHiSwwBcTHv+xlOrGEjGWYdPpMiybnMyGsJ46sC5Kg2xUhvOTP5VBsCqpa
o/RmQ3WIl2jf0PWUHYlnJwKPjVpFKEcP3KFkS9pMTm+06PgPljVaRYzXzlLf9m5pq/BOJ9d64ysY
w27Ay3O+2jiH/vsIUwknuGbG4dyzxyhpPPWRRHrILcRT9gBkPdj+yyHLUJLhBvC7YmxwwCh2ZVDL
Z5qnQ4gdOmxRDQtC/j4xr05WMl7TpxIUkwwUSWGAB0lEIJaZpkMqWPBe6Od4MHrqR1yX/g/QzzTV
AtgP68pEn1ofkbuTMDcEHooGRtnHyhE9Q678LTUCYy7LYXwYxH6B4O+4BGrVVyy4Fa5baaEOuZdG
FAuZN77JZVm32288WxDI1PNDTKLd+UttDq1H/1/CLPLMeGBb10eLzxYtCgzI4KiiTNoLVPcrMtkB
fnMxeUsw9m9oxpV8/DWl+rVN3p4RzgJaBwnuderSpC9GWZfFhU8KkmUys94Un4+UpkBWzxpfqgBQ
1yerQhp6/7j8fB+TETtOzh04zS0n60pNCqCqs9xLdEr3YJXcQWh2PDPhqxTimsrcYu6B7XCXUsJw
oqVg/7ygrmvxasRpW3M8Cx+mx4SxYOXMtCpHgOQXR0n9oQOz5Ej3G099jZdNDeILr3ApLlvPbYZa
7k9oi9uanU4uUjlYf54HE1rSQpN6gW3irdTZU50+g9s0635hizDeHTirHs2KNLGKCGF8Ht8imOJh
TLEqCxRTTTBZH1iuJEwa9XB9G1KbNemGurBVvuiiusqtl/+LTjc6VCe5Mke04Yp+rY1MmKWF7ZbA
Ut83VvoDO/W7tBpSh1cv+r+JGLa8mrSZMD0wzRvsZogJueQc6sULjuC9VZ0eD0JFmZDlNzIFo2Fb
cM7frNA4SWUu/CpZgJqa3MwYdclRlq6hSNqpbJMfiSQciJg+Jw/Dyr4oM4fTR2sOFPp1Mn/ENgfi
6sVWxFml7KaDnoP3Cl2t+4jRPmbo/PFuSMl6YlvvCc+bxXC/7zM/VZnMZITt+APeywwHoCnkKRJs
n7WRFAzu4IDxUXJ/UsPtsBqU6fpQJ2cPqJsqdt/7+Dg/77FdEEpr9rkqYVFn4hLvccOJlik3sQT5
oQf692q0cU7zossek8sNH32F2Tw456LTMuZccAfJM1wLCzTW0MZcVtsCw2Q9Soq4qhTbXMNZjvM8
3O/ZSDss2+FNRIYn7m4H0hIQ1VQvhTYAbpBeJP3axuUbA6CrmuFkO7caD9YIhoR5hBRN2zJku82O
zeG32dpssbSu/6raP0THadjSyi5ngC8W/GTCyWjKyDFVALK7l+rVsjSlWboFFI43iqXG7tciTQeC
2AtIKZhXuvmix/DBUmhBEOIoN2GHYJFKaqa3Z5V76alcuuMXA93A+Jvv7cCSUU8evtkJthZdzqsX
Ng+FwOYZqPLgfBDZ7Vf2tIApCjYQxHdRcs4HAKrRkTUx8V1s/w3o5k7hOuZ7dwgzrpOtIJPbtmOX
vljc/o9Xh92nrxOkO8PnzKTcQR1hr3dKi5VxvYJSkKYk0739bmfSvWNGl51Lp6e8t9DcKbgnHPM7
1jEtzXC80Eb+qi0E/28CkVw+jdGoI/ht700KvOV9CEPyWMDqQmtlqUsG9KWQUk+AoYw4ROU6q/0J
dmK66mciukSsEdAaXsxn+FwcgOzMbsBuxH/FMku+mwYXMmzESAsX32wlCk7W2d0jxXnrjQ8iic63
iINvzLYJcr6y0na6nwdWVXKL+yNL5TZ50ckj2qEM+MPTQqaE8bET3kr6YY0u3zch4R3tyA74nT0l
kfR7TJBapM/RAUuiKxy61KWd73pZv1h1bFLqAMdLB4BB1G76iwS2UvSUBqpDogKlMLLhAM6PSZ8E
9u3RZoM41W8YXK7CtcgochsndiNZQU3xK2peft3GOOgl4Pq0FtHUZGyYBXRk71xgDDmDZ7muGQnj
ZI9Ls5RzwLJILKx/pqXzH2784YXS+/iye+xirXTZxPg/e2rO2g1gB33NSMjHIb0YdFRd0HKaTUiD
14ePb1yT4JU/EyO4Uxi8d40fhgvmmHd5UZWyDHLTmuBXbYKGSecHM4xcqKKlS399uUPN7Py9iyGA
hOhVxESKAfEb034EQtFZvz2eEum1wvfUrhx72Rf5Lx4z4MKR6mTWq2wyUn2Q9DBF6JVehB9KfIN+
S4KW7/Dvx2EqpYLSFa6HS5o9j0OSMi7Ay7jzFkXdheHXUnERGrEbEaE+eWsYmHDXjbaxiA2s/ZSE
m2gUfHXuPhkFP0Z08pCtUa1zK4pwv3pBV4bUL4OVESUJVOk4NDqlxluXoSSZnJprmQdpwE5rDGKU
MzyITyh2PEWnFFFYtv/+/J+cSTcnaxDA68VQqgt4jOidaAPRsvu0R5NXiW2657y5wBqTNv8Bzq/R
6MgDMWghsCjQtbYDEP/ufXzPubiyhauNekHNnrmXYMPCFdPJXZR4qSkiGYSfqcZWFtxJ8yb67URd
vZcXl1sLXNNYNE/eMw4PCjn9kBewC6roGiRymZP02ic1OPpCk3HhafPUxhkpp9kjUqwobqgDEYwP
4RBMg7HXKx5RYZDi+P/+QRSfqHWzhYLqZsgwayTZwJfPLL77ff6SgmtghYmkh7/cFkRoZ0LkGID6
TQPDbt3BGgJ5StlwayAX/78q0COhf6HZkOhMGJTQV+H75Wg0hmaX+bfD9HsMaEnv19OGeYFsTFgv
0WySI/Zi6Niu/ebgAgEaRY77ecE8mcq6YEo1y7aoVPHfwIxJwJwCqGaMrKL1yR4tBgtM1aNsHPQE
AOSUpbx8qMO1foz/7eSvteRq/z4AAzk0FHf9trW+J1/uOkZvgmZtTv3lcMByz825mDnWdJdnXnue
h2oEibLRI7bKuZgyjkwFJb+5ugOsInm0UOSiEXWfZZnVOpM1wHR5RYcWgLJY70mDzg3Og312jrE7
1Nwhox5m27InqEyNetPDvPkAAGGr9PGlha6xBPNkdRp44cDe2U9OtDBmNw7daCSNUYv0wcaIoDa6
jk5Jz4mcMQOOGjxLky/TZyU/G2Qa3enwdkZO8n4lSw+hp73D8OAyzAVG/LJJ2KFZVhf60v+DWjRo
wEJJswqZiJaj3fMxWmXF9ge5hE7FfjU7qO3cO5gSbXp5J0XyISko1Q+GDQRTHsb+r1GBQQ3efi7T
6yELzz0rDlHkXM2HlLUfzI00Zrdemyt0BnVd+1t4nORXtB/N25jKhgClM9S0+9Ec3lNfDGSaxshS
ashdKn2A+Hf7uWrf3LSna+C33+4eYo17+iUake1t5PkD8AhojRwLsQdebtSXtrXor2B6ns51e7UI
A9nZkA1x2tsaP3nAI7L2/J/0OpZLbWtIrMCm1hlaltudF6MkfxLkSNgnM9emw9ANe+7H8sMvFGvr
bZHej5ZkmE1PgK10W8ToMed+9FY2h/VORSqpS3q/YpCqYZFm18Hu2u3NUY660ljKL3BPclvJMery
1rmm0txqC9m7zDjz8aes1mljgAxuACp0Wvu+4/G/3AGMhOokLdznK35Shi2BOZpZtlqXx7Iuiegx
tTBXPwCoyPPBgNT0hq3dk9PE48piOff31+AoRp7DEP1RL7R+ZJJFCSYMchO0mHPJTsgoPmdNugh5
BAotU7Nsh7xjZS3puydd/6NYd0VCMCYkmG/ItkVyrAI9m6WCGrg8D08exItyL8jZzFBo3UX9fYZJ
LKFSMc0pVyh0gs/yUqZSP/GiF6O2dVpLpIdrhTJOxW/sV/23tjk+X2MOcmbnATEFsO15BtJ5vN2a
ErorsY05n1+367hPYUZMoEVvSgT+Cry1xfv8VuBaauh8MqPXhil6herkLoqoyXXmUIErfUq/37fk
4m4MD8wDNIApg8ZMGXk9L44Pjye0yGTFnaPBdb7znufQZMdAbtqk9Bt8pY5eWaQ1SucJfRo6clku
DKVKDzxS8VDFuEgYwBNO9CY0lsHFfKzrcbtV7Kyt8YJopdU8k5eJFIT7uRhAVS/PGMDy8TvXDlnk
JNwlsvBvavns3HhQfxOuJU3uEpWlpd7jLNHEu7H8vs4kzrIHFrPPdRZFx+3VhO/Deafq2jVoKiN3
HnSo637Zj8kJ/Gb9eovHmMDYANou38F0lOKN/lCdVn1oxxyVXMMvQBObUA7zrNXToPdIz/15mG/G
MCvDXU8HZv2waK/rqBv7hRJn9LRIMDVpOI8A16fA3Iuc/hzYINQaxFl1Ww5mRlisQIfWwzJkHvMY
86DfEDS6eZetNEn2tbGfsDpMAzxvhLXvWSl4Op74h6l4WyEB2qIjD2rCCVNqZJqFORpCh/eJntlu
pG2saSvDMziGXshywmA/Pk1xeIOmwulnz3KGkLPbiLV0WqQRJDPG3mVe6zZst9KO+vya5h3u8fk+
3Q2LCCPE6y2kzAei1M/CXvTHP8ga6iSPtqEOrMnXMHd29a7B18uOH3kxN+8sLyxYyqRFQ4x23/Dc
KYoAo5/r/Vjo6l3tr+UzBaob2t0T+9ci7rP79aJqVtpu2CQDrGW2VEWC6J6/QI3ENGuNMWpCeI0E
UxEQ1U8z/MqLhU4kxZWOAJuWb4/AtR6frQGC/h7iKtuSg87jRgL5ahScLtvFxAjZs2ZGmIccZflo
y6Wa0Fzv5fSUcmkgaM8ZSCuV7XT1dUotbFJI1+HGvL/+q3ym6qxNqe0NXNtWfG+EGZgsB6VNn6Ih
Z5iyhTXCjkWxDdy8b/EG/iyLnxucqy5NyfCyiwIi1+5IVu/CE4IfJ2ivCmXQkgd8up16kVYEyDG/
P5qZNwZqgBL9P40YnQH84uC6x+a8tVjJnj9rDYHtYSloAzeaZWnZN+CSTvDibmn1hiOj0XhSZ2ns
fasglUP+g5eXhJGKNWojdQ5sxgLbhOd4J/GLK3Cz8QmJUlh/yxSFUjMa9OW+SB1XFb1G1PdOajJd
AvH57aozNq+lKk7zt64mFa6CAgmlZbRlzZAjHl/P7eq7/RyBWLKpIb15iUywPLHIQTR/MjtQImOe
PDMBULpT9t2R8HUTLhpmnIEj5TGnrDrs/vCnA/03tr147ovI//wlbYzjrHrvVVsyvRXxSe0ehGOa
9gh0jGrED03A8dgYIymwYSdzHeGMEzrJ14C1P5aotJIHkk1KLCuuQGfHF++0WP8jOz5L9IcAn//F
4jS6xswsL23yCZs4Sob9GdWnAv01TkDeCSNT3VKAnOlUUOSm9nnWfDXnD6HvUfz29CyIwoRbSZ2W
Gy/0Wy0086ItFR8EOqbAGi69s6aJGmQl9Zvhe/LRGl0PYyUv6bIbobp4sLkDPl2qHe9w249GY4Qo
vCIaZyNi21jJMeJRbeReg9CkLskKBQAmDOEW/1HIBnrJ94V5yEaZFvm7SYIyytAP9hLFy/de8Np0
vw8dJrYnVGHgfvCt7Gsflc7f/KS0L5/Dar9ltkZNEYMtIDIVZ+JJTWQgwaheWPpmuXPZAB//x22v
tKcv8XvZaf1zvhQct9hWGk+APRYamPdtF8CRHMCvz5CRpaGjhP5+/j6UotbZC0JPooJapcJ/zlgm
+f3JopWDvfW6xuGH/MTCEbqhyNKMEtKLAW0G/dj0EScAUx/p9v8WbFcIKdqnypMFTvPlQTPvOBYD
fUIQjhQ23TozwuyFOSVTiLm0udRMEQPMgNOSQD1nY4MRC4/aakgV16gl2T1VM2RY5hJ4co/HdYEn
kJ2mbFvDzQSV9xTsRAucmkPaAYM/oCWyE8EbIEunzmcSGL43hMNZkIg6bX+jVWPVpZDYXOJnqtwv
75Iephr3JiLvmPjjq/TIhbW/0xdqES8YObnSNnAth7S4FubPoBOosUK7yIyHafucNR8QmT9mAzXV
XRGVlHMI4kzSVPQej16ehK0PQ4g3aL00r4Jt+HxPYBOFUVJtValZNZrdU3BFL7cNAB7ajEElxVbh
81Nt9Rx32m2wekP1TtiGLh8K9jXbnnZSZRubwoUbfEJnxo7Ren5vS0oUPUYgPEHCj8S1ZOTlfYB6
rngWuEF493jSO11Q0RD10luTw9wzGPNWk1Ho9MlieLFwEC/srUW7HPjBjpyrfltjkB5pemuYoDdi
oUCsUpszL6XqXQ2TvrF1EOwspjlGT26OsZ+wnWXSwa0T7OG/L6aZnqhIswAinYOruboapmrlSVK7
Jdcj8COzGRMSiERjbNF0DFOPXVe6iSiS6UjnlkXTDOaZp/cSTPNSUekf6Kn9iOMnOFs82QKEMtfx
/vp5gDucDJ5luVurMVS4rk5kYlbFBQI85H4+t5CYUXlhFBUQKhi5B3k/oNyZ1uMDSrhPuzh4HKlu
VlhP+h45CC9zKVBMn1o/SF/Psetwn9K7KmrogUans1ixZqbLed238Cj95jU2UtbQyTo2oOBoBztR
pVwVAWGIMgZzf9fM8dztBgrPn5jDiAQ+5234zKTPxqWlXkAapA2NDg+8hJtPWySOAgOMNSPizwrq
yqS0cRQLqmqwqClgsvQYqMgzvC79Phb0l8dYk1JsB8sH3fLvOqA63ArmoscDJwPkxpEvEQ0lime/
MKNC356CA8vo0TVoIFGu+kaMouKYgHG/Pa/9RADTVOnRx3B6Ik6j8XBK2+am1ttZpv3CdpZG33rk
YzmeAAi/i1+SK15bLn0bEQBXUxFw4Wu4gUmkCIlo/a1QznV+LPK0Bvj1IBMBGCtCmtUPOmHZtRh0
jfkseEnw7pJDnNnjGJ3aJTjI3muCj2Op9x99juiuMXbJzoZPZ4olaJSlCTl5DM7+yYnjpzQ8p/nQ
gm+60J2yToIu9CFNpCFYRlkaJ0oqQoNfsWtbj5Uf0DGJvj8HNQNWPpqhX083suX7T7mHgRtepdMN
x59En2m4nVbysqio6O7tb6tPFTalACSWjd8+KPqv5HneofvKKT3nx1vsBUYwY4arAEktFXbOjLBs
M/CN73H5UeQPczjjJyClaPG9oyEgpc0xo4Kcpk/Q4QikRoU7PMxS5dSt+oIwJx5a/lEkPJhG8/Q1
peHejLeQ4UqxPc++lDmgnunO0Y+DhmlekcC56VY4ZP968XDBKEhzHmO4xbtlO6pCcnSVpmxURTp8
NObcHWg1z2VSoA6/CrYR49PjEAmPgVrzYwmNfxrBCYm8aQIZoNHzuz5tIvucJJZ878gDJypg4k34
3D3Ecek4Y2QDz6ULFNYTcVay3YyiTIUtjHJaaOy09kQNP1SSqWzLKduQ2j1MVrYLEOt/BhvC4k2Z
MgC2VEgqKNJy7aYTnGd3lr1ve1FK7KDSRBN8X+Xc+sN/NlR2enuya9Uy7KSgAE9rxztaWB16jgAG
SCCa+nwqrHOSZBqZ2yao2fudUCwxt+oFwTjR5pxYqbhW40L3BFUyouZEushJn//TDnl1VlJpqurg
+6i6BDvlq/Ah0xRKivil6Lmc3NhxCatnfVYWaORboQSaedeyQlQuNwZRrdH55wqoPRc2Yvre4cIw
i/Czz/T8ugQ2a9m9G+MuBIcSE9R/cEShf4VNEyDapZgRe4uKoqmbu3tN4do2wdDDJdDFONV/1rqZ
E8PyyfvkZDDpYh9E8tbtApX8pKRLzysOjDIVDGw44wooQe/P588gPQOFknV3Z+OxsBcrx8KkR+ku
FT8h6czcIetJaW0+thpuFaFekj4YWEjzAD1XeojXjYri07TkvCi0hXMRJRCatfOCtUhqzN80SoYo
ug4RSK/gccFj1dbv89J3xljXv77dYjOxsRhxgjc46EexhnhiRNLq+mHCfIIq7WUI7dMftMWtTpH6
cG35sPn6TnDiJacEGKXzwvurTd5jKIHsFRLxv4HYGxlSxMgpk/oc7Iia7wGU+EWK+AdM+1AvES7O
LTU7zoheZSHgchzj60Y2GwcvHvcRBZfRg47AqbUncjgb9w9uch8SV1fWi8V9PsWHD5BRRjVz06NW
1+dfxi5VJNHLn5Xm4AHkb5shsCeb+B9ZnCSW/h53UyAk68X9Nf1jZbjEVDk1Xl37KM2jHIO1om6i
74ZFnla2/7J4PVWwJFNmkBx7k3BG2+4rvOFUisemDrlNtu55untM0FsLUd1JUqhrAGlWIqvUaLnN
3IzL5WlVRDzD3BJvYKoYblaIAnl7RmRneEXBbMqlgVhOm/Em0/t8rrnSBuZohaUgvvUcNrWNB//d
ShydIbX/NgKXG+YZC5vM1Wjw5PpvUE3JzS7g+kRjqm//xCVjlf4QwrTsILUMJg3pghMVAUvmrKHA
lcVXijYa/kDBCxPUgEi+1i4c1g4llnIBKsbNE9NQqRd1P2gnLCZKggflduRxyAiRCH23VL9aIJwC
/cfWqHUn2a0suTIVV4szYdSAYCnVcS1nBel7+J0gwNsrRh1ePgnDGdHk1Cw3zbW4fO165Cvg/iUf
46/pxoHiKzLEgdBeJnpW+LWdmRRGxz3Z6j0Bgk7ugT0a14uA+JJN7Zhl1jrSlxUJANMjd4v5lUuv
wDdNa+fe6xjY2LM/5V1UMYjAq07ll5qN3CtHbNRW6citNyz8HsOB1sIry5PB7Qu9X1GUBrvAkt/H
6Qu1edyPYBERDCwAS3mKo4rgUUo1HzTJ1g+znPiJKU9QuMEfWaKiRcMoejaxFTFurnMvh+w2Qdj7
VkI7WODU1ffVy0h5Gb0vstteXWaNPbiOSkcwqMQEOd8sGcrJ4rcyyBdKQb9PLIaJMCPWots864Mo
nRnpjxHyHjJyp7iFWZU9Q1TKVvIf5arZjZaascWTClpyBMM3ahyGXoK0/c4I8IeS+Yz47YZFzwuT
1JQB1J8W49oatC/1lWFkYDVtGmn6aWF9CxGg0alsTz365njhUm+f+Yxi3eNx6HdQnRSvzQtjS/eN
GcUZE4JUSK3BKDdu3vAdVVtSGPXrBnfx3jA8HDYdNX/oQkkTKwC6qmQqOVPAC1pbOEnmxpD7nyZR
bkkdIyNJJeFqkmGiDLoADdRPE421gH+sG11aRjPE6idYbFsBeIaM5ypInk0POBNP7ll7uPc9G/RI
daq7xPSdVY1ujwM1wx5takp7atGk8FHSh9T7CQwsBXJ5VimCVzR320BxU+LbXvFLFiPDaCzW15SI
achmK+lUfIA8Ok6PC/JOKxz97HGDbW3jTgK8DV8Vx1cnY19AIy/fgaMLKz01DJD1o2w2Ck4LI7iz
Sd/ukyjl5m7wVSj7q6voCOn2EiAD0EfneuCKT8Czby25yin0J5r4B1swC5q2EYvgPbui+tmp4/AX
ebL9QgPMhBlnFzNmvKHUZYe4mSwUZoXST2IIvH5n8H6czhTf0SVjs+eq9fcXpe8Qjc+xhbuMTfMm
5DGZ0bUzqq2IE6YAGt43ud5yxv9OlDSFG12JZAstUZNiWOoNXHpBVapa9+ci1gitb47m+i/QFU0n
9+EURkwlcYqxJ9mI2uXjDdF8j9YQ+8LP/vBXF5DcCxS7BP+4BGHgplNPIq4BdZZToeDmrQBEzIH1
cIj0+CpI4rGcj/HQZje7nTpe+K3VtTNkIvUhmaPW8ti4Z9Ju5iGtQOu84qhURY1O9eN3VW/w0EVr
7Gith2vrTvRFhj1+0KFRA/l2aaUTLfHpFmqgN6ipmgRSmSwfOKi+nmCicjHmTVxruINbQnKY/cS8
gEQQdbSLkthslVPCBoFqMn+hTELeoIFet2L9vv7g5WVjkEBGiqEqDE8QD7BIF6zBfh9Sj9iqo0RN
ErfNP8akNzuyXVAzE7ujhoElgK0RvXkeutyppCPhEV+Rp0/q6trsM4nqbU7xSxcLzgxs6OhCmIrx
B2SJI0fxz5erovgRRXmaaFCmAXJ/cD9onZGGpfbyTMMqF0o2uNGFziuWl28P73DR/NLYV7tzpOlY
kqfOR9WxZoPFrIG/psU/LXuMT569ZMV1rIOyR8eEr+wvLhg7ObDImyJeyFVRRlXI3Nm6un0PM+Qp
kWwS9CCgEECgE/XHQZkWWDwCWp5KmiLc9QREMDS+D9lI3PNjZVzRYb872If0zIMy0yJGzJFYsU6l
5qLj/upjUf3T25tUuZajb6GVONKt0mbaV8RxcwtuG+/nwy9qj+jTE35mcHB+1k8qZmC8SgIzd05d
wBgzqA1+wgQNSQiu2HVymlU52HMiWruIIWjqgqUw5+HKKXrzk7pl1kNd4UMqxs2nAS5ZV34I4Ww8
8pK1EUWTV514dFJZftmI/a4H5N5dOZjBx6VgD7u7pnlHDrs3KRP3RaTmjIxM59NvjsANfDP8F5aK
IByaHtgqT2yW2cZu+Kqlke2u0v7yyuQ6tC89nlB3xj/hWIBW40vj+cIMiHrKaaPEMtGHvSeZRV6b
rH0oizBhhuiI7hZfLx7HdjMUdw8bu1SP4VzL1W+nv41sSbMEG198ivHJx1Wub+peoosJFjXLaR/S
TW6G1jEBO/dxR4FBNKDnZ0DkKhfhYLc0b/zwgBMpPbRIRH5cLUZi8T88MmAikeK5y+TePCuYUWbR
uWxKhge1s8lJ5jCv01sQfifqN8JdumL2Bio5WBH8gU7Ygtv80fZHEwRyBOpJWLKhqBTj3zcYnilR
DQsg5VP8pigMwbHiJoO9ffFoEiOLtQ4LCuiJmmrdS25jsDKVWTgXdlzFifLpzTj9mpiifwjAVgAz
cM+Q9SCS60g1yE8kCfQ+oy81n95KriyJ63eEW8oPd4bq1nQJZYoSsWaO3S2h/X+6LqHL9t2AW2L3
Jzqf/+IlDpofvveL6TrTHeagOVPOHp6opQCt1wxBPskWP/KGYHv/9hppLadUP8BCbxy7Qm9CI4ZR
D/54ZVpTSytIwlmWWhnc/cvoREn5IzEYdl5YzG0+l101lvDVb1tofTztwe+qjMCp/dPVqtgjDrPm
SMJjhXJ1RIU1DxCvqLN3JwrpREqvjilDi9dWdEbC25EkgFTNvmXsK4nAa0lSoGUv/WJZAHVSicf/
/pp1AL4c3DvbMATZB069txjH6QVEOf2RK8PcAcS7tUxIkkJ+JpDtb3swN5LV4SpzrWKrkSZXpL1d
bNNGl6zbnBsCn9G5FdT8e1hJMSSkM7dLy4yRVPzkSJYNpi0eMwalc7SbFG6finzJKNWKv+6+qUxd
3QFkEYdjqWF4Pw06fx+0fjC4hwj6wCuNdq+FKlazlNIfplkCQ9EKdz1akRLpxRdludKfPWoIvpyO
ds7RIQEWnTsOL6SIscCGMZgFhfcGb5nGuXxvLOfnauc08bfVO897XYYh7DGr2alzTiC91woa3/Fa
wpBocG2A9urgM5Vme463bKsXV7UfmOP1E1gr7FtaVi7zzDc9q0FGSGX5ouXUGMWCuXxE5BIid/63
I7MejdM3lACRhMzrBcKKFP4CqBzbgL9PumwZ3MkZf7/S/8JuMGLjCoqIL+p8OgS7ObMLY8zL3hi7
Kgz1NeZxJRHrfjFPuwcsQduH+PV9NuLWUDZuDaPVSmUo4jHhyVEH0iYkxFVhaFAjHzx1wpO4K6gc
PVXFz9guMRAwDATPBPlIFSXIhzSewHlQ0To5csSlmHiQK/UCykPreTJ/FPQodQLN7vqwToyBQrBP
JV2I+rrUuX9/fc3jHD1t6tUCF4KL7OLYCtmBSjGlSGDcLXkERzAowcOrpAB/Lnw81tAceI87esWu
zjpC1ycrU96/Yincs5BBGTV8Y1AjY4j+merBjiBVicv4+Ms4ja4EsUudRjRHFfHEQVS9XvQXx9ow
ichn7GXi96ioyMwtF1ZtNCVa16FptjI01Pil9/5ZslhrxWkC4IL7yBRCpvCfwpE0GxfAWUrkZBmg
sUrQuCFSE3/D52PDqXlniBgqKj2c4JrwRYgeV4IMPckco6Wil3t2ZPCHlqvKuvgNDV+nhQsVeC1G
l9vLWEfeQGqnVEgj1aFk8kBDKbKtjHLt+670PZewdAw8zMKg2Q1RAbX8uQNqKt+fZaynrQ8hOmpW
dcwoejwxmr84IjgztcKPHXfpmxoElPFXfMETug4RCtpDsdtbNrujQ1iVquwN3E3uRco4/M3w2Nxa
U0RDYBbCenpwRJKbDs4hAtnHBvK1Puuoj3rkUzAkKucNWCJo/gwYciebtWJ4I2S+rkQuoT4c89M1
Yyb+P9BghrFYaRQeU8ZrISBkdV+Pkyqcubkyy9IYcPrUzG8bI4hVKSagnn36lRC+zHH53CnsxMoz
lJ3IEVJ0VVSLs0UZoMHMhMK/dURlAH9qQZzdtYtvJ3MqTot24Jx24ssGkMcM4Y6kq2vTpFdAeiCx
1Ho7Cp3eGxY0bcSZZs7vTUuz9mM/H3gDWn15VadSn6S5GdST0BJPPro5haBDBxHxjTyBKEIp9Ssc
hjBJvOk2MKScaKwXMwCl0Swe3hiL1BfIcuEI05PJU9jL3ZHOJMSw7AIGn7EdMQHgHbQ4awC16ZFw
dDMVUfahPklSfQ2o3xSkCHh61CQQ9mJ7gDplf78KZLc758AGBKL6XmdEBuXhEv+SWltOAFhZo6Kj
GU5Pl/tz+HZ48Xw/yzc0H45ZmAlgM3M6FOzDT6NvMhBEZeu6mI3kxVSoiclcTuxMD81/KZF6xVm5
26/yZFkwUlH9BZK+5goQXc5ICgX14BdDbk3vPu0YO+UwO5CGLQcPGT5VvYkHxVnrVjvVr9QckOxk
ouhG+VNdBJ/Uz9W8hiJe8KiON6s/N+tyv3ET0ylFLJ//ccgE+YaYVdP7TVeELdHUwhyB6swyfDqi
w1WGzXweMNrELQUOkc1Xg+SkcY1v8SfbxHgaAkc3eyIbpTXfpNd9LyehfClvS+seFfFRRbhHQAIr
ss6b9E7msVfoCmePpZ9w0Y1ApJxK9mSVP2b8DyWqH2Z8FLd8Oj58MSY+O2GHYMUYcqgqmpGgC7+I
mvgloNcls8VLnghbbgJI0mxq5tpkQZ91K2mRGszNk/A169BJCQYfzm/VkAlxOnX2ZLPOrVIoffBM
Fujp2/39JCOvkhi19c+8vSKzUY4ZC3w7HsfqzpoIG+TNzbvirpeW5jcX22o0MHRuMwBhb8gTwh/t
y592ycPP3N842j5XMCjWA12roksf5678Os0olMRYzn+xKyd9VtnOVs5gaE3feDN4crJXa1QPHNEy
GNZr57hwUaM5fy28DPGP/trsSvvPeUcse9pHN6j49pWdV/RJC2w+SI5as+0WuMLMJZYVF68jPQGg
HlDrkOCVih5GS7cjX2+o6FyLM09oq0UevImBJAMoAWoowv9uqD/uSFK3BMjTvt4W5u20RVap7Efn
dmQJhdccWzTa75eTczA7c0XeFKOIk+Gzs5A+rrbI1n7lAeVgpo4yWaJIXYUcSNXTVJSeXmDK7Q97
y+IwSqpd1kO9KKY1E0niYQiQlSKx/P82x2J1HWPfH5EpJ4kvd8C9SC07yrINXWcGtkUc/MOTDTLq
1zhYcad2UBCx2+Wp3eqm+mDvEKGypDBJjajhXz40TY6EVQ870Q1KR0RIyFKl38rXfVHCr/Owto3/
MhZ6A+cGl99kEoBFXpQVu8HJKpHNf78kSZNr36n8t/9JPfceJnO2270Tl+749AX2y77W5gr8pLwd
DzQA3M1/Q7Y+ifph62SJaM0tYNAv/4C+ncNGhHjGkgQ0NgqzcJArMwWGqC82zjyzOK97JS1Dk5kW
LB4MxMitfU4qttGzpx2qn51xSV6YqceA8KcmF0kAWrVcMMHyY1dHx3yxeWSD8VErp2JbJcUnrWWA
TKzDfPCxn2quzVeZnZWtq0zfHxboUycaRl5RUWMFtGHgn9DIHJjSN9Sww1PN0pWFyYceDthl/M4/
s/zfwx2YReH2XgnM+0aFAqzQqwKl8C+yhB06xIoaKljDbsM+cS+Cs8gZBJIg3Y11NIvgeVqgFUE9
1Mye+GTWv7QacQ9E19bzgi0eEak9oilUVRZ9MJP32iijv5qoApPYFRu8PznJ3G/FHPKlf9jPg3SD
TwVvAuif6SdoTwqnA0Ajj5Gxft2nzpdtRy4vrdT8ikhsr4hlvnLtdmbQ5VlCMWsaewjAoNkPrIS1
HNuuIx9i+X/kqisW5LYp4Aw3xDFQDcOscjuywu3I0JyXNHa4j3JvCj9j2IB/x9CDqaaEGmKaOteM
oQm81YIwDr4x4+Urz9BWtkRtySh0m0ZYIKOUL0FyM8rHHbuUVKWd5RLFS+3zw6zNXDCCkvaBrGpe
4IpKInlHUwGyvlbXiH5s1yiLlNJ5wp59nevp/+AiBrr0+v1pas7XpxkzHC7ZtcHaFM21r8bvKzix
jG0FJb8a2Wh6kw3sLDNrTxUUYzBhY82A/9eH1iTs9uVNurmgoX6IH+wR8pAWKUKfRsp0VBfmu0vE
JSHjoIW7DmSUFydGgW7Drel5bsKoNhSLwXcIxLOnaAJ4oA2UmAYwX5te/ZJqwKWtk43NdoJ0ihRn
AQv/TwbblOMXOminXe+RxGuB498lN6rB5pDaOv1JzQvrPgm2QFEc2R4hcTpnuv9TMg/Adv3suaZb
XXQhTGfXcGI+ZifyACtV2Z74IP+yiZJFNy+bbgI9rIg4ggei0wIh61VFlUWaFJ/hAgNricvLgDSN
aUFB4h3NmvLxY6bUZPx+qkr6FHto7f+0fveO6mlaTg67iiP1s2p1xpYmMVZWo3IAQ4p/bkiPdMxb
Q+SRf9somDsjxeL8mLPtmalPJng7xy/gZp0224uYohP7BbwNrlMb4l9C8FMEyc8cqH2SQVF2mHD3
kovpUulxoNWAvpVqa71qOGuyIYHdD6orl794kg6Df6wX8+kIO3gfY+kEnC2R3ol6bL7LO/jpCRkz
zKln/UPxsfS55KBWS7K1Dwj361ZQwsaA+18XjuiR6Jx4YVTaY+C3TQHT1m4iZFxfrYGrwrtAfNQ/
GFgO2rLyoss5c8i7V9wbF4VHTgtSPtHfiwD3v61smqZCs9Wb38FgpKSj3NhGgdGbe61vYYKWpqs+
3Nhubcb4GTOK8jKYOFGZYkt7SnHy3Tg3PSUQacR5C3F2QXI+IW58WFcuTSYFmq5CxE0dz1uydR0y
YhSdqS2NBU4Soja+YkHhnwzt9bczxPGjBjC8QFGoT6HhRrJkZugj73MfpQIokitM/93jIlZ6paLp
hVUnnag/BmCPOY+Yufockw7100hmoB3kGclICW+tTa95vK6xYFNkublUvLL5e1mMgjtrdkoPbYUk
4jaJi9k6FFIt9R5p/00RSaFockoaSxs2TZOcfp4cVdZuu67pmk9UMA7AHS1QtSE2L+hLyHUG8gis
RYRhpkkCmydtv0jkGBRUXY1lL3YNF6f2Djdb5hsuwIdsivohRIw5HLZoHaoFyPASuH06i0xR9wqC
P35ooKBOcjKeCCtANOuMXZv6Z7CSTQTgmdhClLz4OCKVCzA0S+heHfEMXBz/yxKyrkDdV99Ly3AA
k6XseUkrqB2G/BEEuDwyHfCbD7pBbi+OZjZbo7WVYXv6HXj9v+hIG8iRNG1QLzI+zX91HecqT6Wt
o1ZZdLR7OIuB2TYvU8ijwyd9kVOhYLuUccwW5/9tnRCQutuTCGHiKMaVKs/v8CfMTVtGzWO3hZfp
l2JLmoGSVTIj6xUuFDqToKmhWryMhdyqi5hxdtqq9/gnicOSmNsmjdyXAGlxJK/iFuuaWbUf4h25
uL8b7S9yC0dUxYnFlianiW8p4OH5n/p+71hlBYN5Coiac9vyqiUJZVpII8otWfP1ld5cLLlqKyzg
tMg2TIIka1HCvil3Bcm2tZKimlf0RtqKwJeyiquT57I/OJtANTUQb8UfRUmP/D/F2c539s5GDDtr
4sfcK2AoXGJdVEKsrtFZoGYJ7enN2dCtg8EyLZ7NfYH3QDNFPkb0KvwEL/GFv/KMDcQ1QBLqxGMx
UO7Ahkpxg9ZxGLCjHcVTQYrKIicc4t2fzwyiFGT76N1D96D2QN96O3gGNCXUJOu8QEQmeE64ZN0z
YTQpNeTk3HeQI5txnlMVUDsihOBmRrzCkx0LAwT3UN87wN49FkWMY0eTZ/QwS1fSQC4AaS74Tg6k
bGu1opVwnUUTCzBHBntnW3tshUpFd9HQahDJTXH9w9O7LzxqHmU6VGdSMVLnUs7N+zlNMoEwElbi
VzQV3mframvu49mqItgmgNr0vVmz5kS+12Eswyq8FqXEsFTcgio5KrfsD78ucdMvkS7UbDKqBwQa
IX9feD+L0CgvoYUiFgeMSnAj7wWTaV2VbxrR9ZxIvWaBv1OSTgRbRNvmpMVMFQ4eVzE/1wSTlDJe
fp8h+sPSENZLCIgC76UA9h9nqNY7HLTTCwAOaCobrwaavuzF+1h2OM2fPSbUZTrcn5XOHDd0nR8+
gnVDn7piwy2Qhapwzeo/cvoDF75owVnj/t7Jd2vCzHUKBgNOyEgQDSQCpaSgjEUpFXe9lt06zY/9
yzkvxtl5Fnvs6OAAK7VuupwX6+JssWcr3e8yRw6d2DVzk3d8Ua7ZxF4O8iReBB/p+10Iz0yPkV/O
NRHdlUpuCogb85e87fFQM0Njxc3jxpMhvyPpKD3zM/BmYAb6HrX4pOv8bQmKIM51XrvSbCsqVT+N
qFxeV1Nn5JgMrEiAXsn32l200h5bR1KGxjm2VVWvpTa2bhEviWi70eUvQd93+KVY+M66jKURIa32
6w3ApX45z9Y18V8hcXEWf59yP8PvWLJTj+g0JQ1vAKVPIriXkqW3B/mlfgXUf1Ds0Z/2PQHWMQZl
y+gxTDGckwQUxxODVl44ihCzCAjd7uptohqoqFCgjL88QLUPSYpWt8nO0j4mTrLXRF2ApTK3KtIn
R504lS7uZXXQq/6ABGFEMovhqdy3vYpeRw7B3UwXETxuIdFc86MbBjfdoLLLu2E5v7zPbQOeUiMc
nR9X9vPNIw22G9AE+fAVzQyK5ngUqahHq8dE74Dlp+DTSGp7SkvJZUJgErQn5aOB4ZpRAyXS3h7Z
4NWBCXKVP8NG2P8bLGvk4IDptOBHWT4FbqkVt2DAv+mBmpVqstrak33b5cooTnMnc2bpGaR4uBIZ
BZ1GoVP1H0szWWMQhZ5lazTqjVbIeMIS+uO8gckXCFTt3qp0modozVXsCHcXBNZC77XFMDQY8PDX
b5PuaR/u+CSKXDNm2LWASULBIPDnz247oHfEWsIJ11CDjcMOtKFZiNjq8hdWO5YDUfHhHp/IR//C
r7jKg9uGLMbdI6mLslJQlkVbppVeVcYuoQLEwMzIiwr7imBwOkx276x9ZDotz8hhx0UOOLXmiEeD
vYVz4l17tF13aPr6WzGK3539rAv6CvAJ9sDu8MbjzYS8LdDtb52OabZHjeAzMbKaXgqMEvCiXjMd
V6WsNXEVSm8P6jVaPJ3ZpTF3GiiTt9PlY5Lr0TONgN56lOByfOBbchxonrnYtKgHlVdbqPXTK0jr
SpwQkkE+WnAfekQHcCScNijlLhXyOpvlvc96osovzJxkl8S0CiOnnLaExX51aLDeJ/KOj7fBbjdG
g+tzGYngeMsmiJOlLZY0CXNdeiuqYO3MvgvXdX3BLe1d2MEMDk7ibdMzo6gfbVnhagxmx9zjCa3Q
tR/IFH3/XpNWJ0O8/2MshLmT17Zb0JfRvnjiQJdNEJl7EHWX78JLDfiyPx4GoNzNgJ8jHPCBHl4w
qMkAkqG9Bk+VcfRIUikybBSLSojopJ9M3YnS/r+Hyx4t94b9q0BKZQpu9j8W/NOnc1heiv+M2adi
BleE87ulrV2gICWLD8HA6gs6ATZcoyxEH47Gi2UTItbgBUmX2b5/tjT8MlJ0IciXDMJo+skowbh1
nX0EVPN13BNnMtneVf+ZWKBxph9KO/G0tbJDqklGHgVPDXbRwL/JiMFQhCx1s/G9tAaIAGp3Z9WV
ImFpE76A4TBsmLGBFO/uTEYXK2UoLiD1sXQ+3Fl93VqKkwj0WrPbZJ/4/CJoRHyfwKDMYoJhrx9d
zOUoqjyI/ay+zcy+y9WJqB0IVS7b6fy51pKI5LKFOzsjNsaws1UmuYlRWtiTjgw1x7sS5lH7J4F9
GNfU/+MXUASVo1+cdjzleaSMKYkamDxdtJjrQPpLq5QgDN9slGZaP9Htbf/EXroMA4PI2QPltWFm
Uja5/Rv1qTOpSwdt19Rf30A2hgu20r20+iWru707hnOBKj4KoktlJE3yq7OwXiJfr9N/wcFKzHbB
Us+NiVv3nD7A+cvZ4Ci1859PDBL7HA==
`protect end_protected

