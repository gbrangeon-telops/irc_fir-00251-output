

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
jtXjITQ50a0ecf2Im0hc5gDMz+eLQYg/zzqRdEOtUonTsMauUR2I/zDZca/cFZRkz2Bn/e1TcNfn
wKr/p3+6Ew==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ANnTEQ5JJem4BDOpiZXGW1BGnlByArgufttfMLkwemXR407wjOM5c7+DduQ2B6Rws3h4VtvHo6rO
wrBVcL7VsvPq1+tV939t3BGzv7HmeOgz+bF6BolXyM301AxlRkWo/0oJhXt9sAWYr7zYDeoXtQZb
l76HOHad93vrCilEPkc=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
XmwNj23lI8XFGQYG7vF9oV5Kxca20ebqjV8UOZJpCCCr+xVAS7ag+llpfkHEOHuw9tSDfsd4Eagb
WTNoLsXhoBdOAYPEcNzU+W9qGu9/wjx0qrsJ9f6NyxsR8o/IzcMAojV3xWACKEn/35hhcf9UXdPw
jFtFMZBq82H3pspBY7rQB54QzJyh7kwXdtgWfJuR8vKgpz2Bgw+sWz2/D2DHqFf2M9nR9Jj5wsYi
jA2guHzbYFRqb3Hyb8w16e2ODRs1Chv6CQa8J/8jZZjpfNE9JYFfYFbj02jB3GIgpxkUh95YsKVS
nyG+AAIy66AvGO8wjxEaZssb0O8bFU7NUeHAaw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
jhiEXYtW8X8urAKsC5DlhfR1BlhyMUwpr7b+LLkcXXJrwnqMhkaTCeeV/MLdD2fZlxbKcfLK7F9V
JGPVeMHqW/OgkDKoPYInFHgV4dQ8+vVlaEgOkFd21VNxhDMogpMeEu/OUw7EcrJ+uVFRL9Y4CZQe
7QVrICfnVX7/1Uf6PJs=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
fOUx+hBZ6Yu+THnpJi++K5FNQDW/3h2F0eesEGevzvwYAUzmUKIlynhcf5gdgPU7azk/daFeo+yk
Krq/01NBV0vQpvK8q0FHFH+ghuL05juk1koa24QZKqKLJESEoqe8+SMhcjfeA/1/cXTmsbZU0sOR
598davhiRIPeODK4SAJwb2vC+fldvr29ZQPfn7IqVQ1mWsnCoHzWBSYPyy4Xw+6asrFDW88G8kf8
wyRSd13FqmDW+hKwsLgtlOhvBagW21tHVBbEEW2kPEAMrlmNhaLMf5utkD/lTPuEPBItEC5xgDps
hn/cW4ZYOpIgB7hTnFioHxnAEnyoEZ+mfU5gPg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 23952)
`protect data_block
fgJAJNFU8n3pyvgjJRjmQGAy/zQw2BNtlaWEzwiuMl3ElumHzz4s78YysF1Hp0QdPnkM/wTBDMLC
8IT0ITScJPh5Yj7/ujr1hnAYvgF2TYWqLUldT83+tXiRuaBWYlN4u9w/A/NDSiJLY3O2wCo4ZSVB
t60TNQMzoM4p/NqVFCKR7jGYHIXOmIMyZ61/un7DqmbG6Q6aqseiC+k20zXYGX2TxkL9cQjLpm6i
36jVbsEMcHsAe0qabtzS3Ueor1z1e0R3U6MI6wBwDQTFwweFoBHZbz4AZjmIjbw1JSx9BGjYM44r
eLEX2O7A8k89U26cfVVzpRzdag9bqae9FBnKcuDbE2B1HpIBF/GbW/XZ8VOmOMgbuImS3DzDY8TH
nd5T5k20NZJQtBipw1xHb3x3uK1A6KCHdKPg1wlo5hQiL2jNhabOjhb/6JOlPbN06Ad1Om+QWjX8
sTPI1ngTux7sff9OU+CiYmdM+JXzKVTQNQCqe4PJjU29c28oEGaucg5mvNuFIV98jQRvgXvBqcdu
HDq7MV2XuwjKk1nJqGCE7u3skFGna16LJUv0vIXUOn4c1TD8Mufhj375PG3HxnRn3B2JKJ01Vyf3
edJrFfE+FK8/A7vOwAJfKL9igBYn3ls8tQcd0QowwbYiWek6a2GDCkJ/3mTTyV+NWwVC8759V2rz
fY2Oer7lFAwBpwXdVP5WbJxDLVC/FOnZrPId8lClKnt5qc85Mxpk7cV29DbYaDrr2kEmt96MzDmU
Fuywsgk9NGuH9I7eE54akQpP1xy252ClH4wxTvqkl6Tn9qNxD2wYZp3hq1GfIthS4fpkd+HuOWEi
54tIDZgeew0nFyRiBPh8e+77fEspZUx5BuSzKHfhq0Zonm6ja1yIPNAecIzNKZsbGaDxu9t3Wu1p
fzFRZptfFxqCEb4cp+zd61qNouNxby+w+AtjNlVjGJQF6HyupGBMzdcYi4fyF73HO2KggK5aXogi
rg1hYT3kzy8ZtT1yUOdtBvP/6esQjwQaoUPz8+s3/mod4Cu6XacTL1/r5lo6A1bPPZDkED2OEwc8
SarDs9N5GzuEAMaXBR7HTbhi2Bn+YUwF9gFJnnBy8ZXXEgQFrVh/LulB5Mo6h33f5MU521s1GMfx
B31bBM3Rz7OMn51N/Od37jpLScCQWrkFDixrhokv7X5bjoDeteb9oR5/RXsBvf4NXkZryXindVxn
SK6q/452Chu9hZ4HUG1RGEd4BAe2FJmlV4o2gmRZmyIg+1rzNxxBlLhjwKzcpVCue8MMCeI/yZ3Y
RUT+RL3bC9d9etpkerlWWqP9kodjTha1b87qHJb/mKHUN8Wri9tDJLRFKulH/CT0h//fGUYJx2kW
sMbdhu8OPiU/kHcb4+TZ7JQYmDO0hLIU+wSoFlWvxlwm5SGm5lYOusXANxvHCH2sRjXS4QXYxv3Y
+pQ4eCHQ3kx4ld1ttWQBU1CXni5XgtSn+U01DfDch+vme5bKQiOxTFm1OtEDHb/i6jghHy+mCymo
9MyS6ftEw7TrUXyBykbS2X27W6m53AspsFumEXb+uTlyL1tdgWczFVhsgDkdbJ6KfANckG8iRI/K
es12FpOvCldQ4vx17m0n1inlU9APlcwvbtPQ0Wgp04PnG3iBC6Ywtc77nPFTQfS1XdNJFpthYWSh
jjZBbChTzNV+klm0TDOsyUAvlr6huldzdBhZxL2A8Fcra0DJtCjx2Pj92PKFaxScYuvX4mODGQRK
GXRw5qAlDQtP5DfE8wYmCH0Tv3fSf+GxsOIyrUuPdbHGHZPPJeQKJwebfuGHiHqZoX4/Rg9INiXz
B3LCKZ3Pg2koJnChqNlGTo4d+CELPyc/jS+u0kwdpclgalyR04kjbRp+X504cpsy4pOm4pdOCWa9
ADE+Z/XSEL0RDW84X7ECyXBDr88+6RWO5ds7iiWq7IgxRDCcRhEDgOjbXkgGWwUC77P/5blov9/C
l5SCZTGZDsQSBUgROieBl1Vixv1Fs4xyLx7Wocx7nJKBEci4FOz5kJEiuBFI5zOLOrihu62AwUJ5
uHhYbWtgq2T47Az98E1Gkpsmf+huFmxg0QmHjflsYfuzjCXbj4fJ5fCh5vjBcw0GgLe8iACjtQWG
DF97nC38yVQdJxZJoZvEltkaXgShdtVY5VN5owgoNewwRXxyfeXDFxtHlmXoXINgZdd3XV/UraNZ
F4XDTcjDCX8ZxiD0DGyemtTYaKunEN8Qt2/D1gyVp1Tb3gVyK9sC8UU8MZXPMRs7QGc3URD4QN1P
PPJxuyZusnadFB8tNWrkoEVfaNlo3fknLLF3X9W0ibghU0kKLW230GTWEJmrjkDa1ajvWAW8uzcN
lr9bguK1eyxnADpoch4uDaYWMrr7y2ly/pGTjMK3qSbXAjO2Lsth6oAWLa1a7yIujBYoqDoV8QMK
8HMnypbEAi35TsETE+9x6HvZM0/vEjusevWRGVgtq/8AmIZHZGrjXFaJ1g3v7tHkZyv8w0QfmhYC
OA73j8yHxfUeUhaX0MGcgUAoCWGFf8yLU/DJKUhVg+izI3X0p/dkTgZX+SdyLN5Su3jmaJ67/t7Q
PKa8Mvj8pBLupF8Kx9VszG9A2kTwUKY8Z+BymxNlUmr1J0yXCqb72J9LPsrwboIA5nPcYJhFvl4n
ocYIpAb5XB5LFvtBligt/UT5o7CJxybtOBUVlqaDHp/DNAguB7jJjnw5GnHSyyd/NrLz/p7utaza
mayRkUxBeC720Bwc7dLNVrZEQ9k5KlVzcef3Q15Zehx1Bs5hAOtE46COSGjHkO8gNzJ4VBdp4ZTU
TUURdVwEcH3OdnesizBhEhbBenbWq66pzPbJRlVMD/curbpcsOyU5F7iIHLcWXdaVjkH8FzlwVV2
Asyi91KxGh16s+CMOCCR2Pk5IJolAD5L7wv/ww9A8x1jj7EpuQn68wiFU1Hbzq6MEJDxA25scuO/
T2J+nb9XLXu9zm9gBp96ODHbWGfSVggEmfB9KyDIGxSAFusOpH0Myo+OHDaoxEhuot1M/Oa0SlRH
h5EeSzQpFDRd3y0poh/VmNqXlK9hPOY8EfOQgaH14el0iSXOVADr1ymnzwBufEqs7chvgwp7seRt
K+CWA7V2t1VZt4U2fbh1RgZ36z8fpzXktLt2/nlbQTv2MSjqLUL+BTQ+zqb/WoO6js7dTlhah8nf
VO6P+UJm81cJ+7/JAoSaqQjAd3E9/nQeGIhgsP729O6HoCz2Vtwj0toIYBxYpD0Sb8MHf9T8dRvd
yzKKkONM8Q2Fezinj60o8CJBMtnRRhDGJHA6EIrEJ4phqZyhbuniu+7FqhLoN6yCpq3ieqBbciI9
Q2+2+LBjDVwfBKSoqr3lKNTnHIOPQb8CZEiSQxPA8qyS3oacsyAuIty9NI0kJNF92U9TZrsoi9wN
1Vxys9IbBrqXB+1nPcDcwdkq1xPwz79ljKTnWMg0JpXfsBHK7Y2nbkNmnM2Yj5wCFhN4jWzKmsnK
07gznNQZmN2g5ElITh/WCGx2d6UWvE74wJPsEhtqDREPhFRmxrWAEq+huZgXk9TKM5L/8cik/Zaz
Bg3Bwh3l7ySnYci4YkljZ3KN4MpiRZnT/x6fsZjExYAvY8rILSY8GyyuxCjT0cH1lnBS2fc/gong
fpaDAlo4yqB4eu40811AQWcRXlTezkSuRYPv3CcOpxQTIJlGkZPmrs+sHquUq25icpQSnL8TtpJt
zQbsocmX9aSHNKyjfsZN1WljrD9om+1KnQrP37yTa8Pv8ebRXrW7Xaaq3phD5LkzKMQeDpLEBqy2
6ZvLvFNGCcdKQBW4iR/l8lFobR3VV7X79gI4NU8nHMt+JdIr6fzNLQ9K1vD04Y1mxMaCoo7QVHgd
WzAMLQoRODmr41782Dwb2Bjicfo9GCIHYbaotvKk7HRjs11RN0vFcfpFsVDjwlyQSwwFhS7yWYij
4/0yNmTkt1a48NoXUMRYKD+QCTxv6h8MCMk1skf3YNpmyqfAqoBa9wGjHwKVIcP/Rwpv7+gp+6IQ
VKsYKem2VLFjcU42N4fbks33EdgEieJdXG0dehH06jTYCQOaM+pJsO22gi9rUdlz5pJosaFPUQOP
lyKmi/42BSWVTlLMG57gAGBYw5psK//jqvbyOmOiitWRGlKJeLdDH0ehyFSe2utDgEUa0WFxFZAe
BUnhTY3jZj3Y56A/R5trc71nBuVFZ7mX2kE+MBAD8Mkg1+tG2gcyHq8jR3qaDDagB9izikldV63Q
cjp0A/SSWMv36vDY2YXM7Q6uvYq9r0q8ibVcpAANWWwHd743V4RjrwMPO8OHPUfywIMwD/DkOg4W
wxnY1vP1c7QbvRRkcCESX7DGPXetrzcqC5kzR5jHBnriIf3JN9NfxFLsfQXn7TPkSqkuVI/IQgeH
kaJIndyLAsIfT2tNZjsx8Fz4tf5dKUbMx+ypYccFqq4h7g28SWN0O//AiiK+KwRYnUcZYk84jpGg
WoYiOPJCNv+lL/4P+sbRfTfmbz6Tm29w1YxnSZifD0XcfWFLoIeU20olAMnDIWucxgmC90smM+N3
yvMKv6Ng5R4sIoYXIow04vN3HsAwmLkLCUcJ8jTjUpgSHWgTrFJlbxpmvk1U8IGT24eTR56rje19
EQfq5kw35v49a8mYcqEGMrC8/FHyLj0Nny6ou3Hp6Og28waxDJAhviiv4pmZ4TJxfbU/VoNH8al/
cOvAqPhB9BD55qv+jodpPQaVCvM705ksdINyB+991qUWVLjnuV2w4uEOrS95pm5u/c+VauUCnmSI
wbD6sSej+MvXu+ROB8xOdZwdTdbrEs9cMq04sodB0LpkFK1sn5Yvqf6rFxq8VpFbNZlXYL37eQAF
mlD+PV13MCmTeRyuwFWJhde3O7X8F4ulSUTrLLctGz3/v3NeDO95s568nL497uu7Pasz8TortxnO
h13PPS6mmFOJfFGqRh/jgh0xtceCpltSodYXEc2dXbA9zcfHdSmUxeNy8zymdpb1UkZ6QR7ovks9
gEAW3YGN4hBKGaj/qSjzhPvvXvuqwStr8dneD5JEy7+2tH21ZwvI3XXLJBERdSCalAusDc5uTMYw
oGtIplznfhPYp5w2yq+Y0GDlq4rP1w3G63DB70tW9IJ91ziO3HC8ge4rI/iXorm/4/vyzOpCmnJE
VvnW8QD3h1tnwm1gd7uShALve7jT6RNOu8Ryj4aX1kjQDWF+g+6Zp679842h/lFL+zaHJM5pmc1W
17EfU59llJ5UjYQJclpWhl8UH6n2ujb9TSuMZIKC50GunmI9cYHNK1z7xU+EJdya/nbSGdcqvvep
nVqXG4RtVTblMHNF4RyBwyB+cMjtxYRMzNfttYbAFYqx95mkdUOdtcAGi9N5Or0fOVqycCxrFBAZ
CxLI95qHq+EekdpLSClA4M5Kzhe+p7eMrSkz3VnKpS4uaegeI+PVi/gE/7zhtNAoHqrTw8hGDe9V
EDkjfylIZkrpkZiQvGKLQYM2vF/gNllScmmEK+nYNq9NfZRH3eZwvArjXBgI7IScRVXLe+a9xtr2
P8GXwx1CdRQ6e3FuoV8ToLotbx9BC1c63uDR8S6eKGjWPs3I/JwKwxm/4DrZ0FZl8YbvOkysdCDF
n/S/gju9YrR1DIVwYLfOCt9nnKeFVygr6FS/1bkKNt8bWdM9BCMUtcnyNjyRi6pkTYawhG0IP9qL
wmrCLADKm2ASBjwONfVaiPsIV+YHq5r2vFnqkUgYd5S8UvIZ5107izx37V7EmLQxHp8zC74g3pE1
wk8+39Yw33WOTlOHkhc3Lt09Zj+dJVwr5SkXJMKba4N5rDTPgRRMDM8u7k+TlciDnBeba8OOJSlm
P3M0I/Fjr7l2x2oD/W6M1Xxxm2l7EBUGAbuMmiCn/tfyCbkTohoF8Wqi18PvOGhRaHEN+S5nJkW7
soOaKEtphek1ZN22padPfeL3YChzfStjiXEOp8T6CtHfe/lppAbtxZEViypc9WrCAHS0cSkqSRyz
uvTqLZWqe0GzZj6+8sE2A0YAKyIlhYzjhfy0Sstr2xZx6fu95L+0aqv6qTFiSo90XCkn8DToMB5a
cxDuMeb1AsmBYal8FrSQWIA86SqxXEc1vPjlAXx8NPup4nKR+a8j9Xv+k0B0fIF1qShV+yWZONFD
hYOd1nTAbdYgCA2c2RqbOQjuffj73eReflKSh/MDrV227VIzKzeZeM8hoVQ86b9RRJgxeL/UDuUx
65L7OEYcSwHlFhwOMQw9Dc0WPnSDph8wJH2XyryOLOqjc9dB9JhAbs1JdCXSEW8L6I76b+bxFMu1
zRAYewc5wgOP242adZzSuNTayyFbh+n9FjPPVpca50oLNT1aR56YL2/6t5htYp59emGqAj3dIJx7
h1dvdk8hBF89aON9DsnxzGSDQOdyzRZZo7y3olKUYKXyLcBbKCBQ4AFyf9U98rHjHUB8CV00kuei
9R6+0jNTSOOrHeA60rzbus52AL7ZRDn2LcHU5D4B6crgj1Xholn0fZRiECGYZpUOTUZgeXi/0G0w
9MFGTSgbrzBZCeCfg6k4IFhPxllzrJ3pNVupHZkQugZhKNeLGkEcMTZwX/NuVadeB2BgSbvOb3+o
j6BkOnrXsLmwyHVY5wHVL6l9c21VkBClp0ia5N405gebCJmS11tijNa3fmVxj0ZMoelawM4zW4OF
a7aliImWlRWmgm1tDlo+hpFlB16rheSI0Ek04jl0hNBvBhrV5Q6OFnWNlGWCONATgcjQNEt16SaZ
VVgTn7HMtVOklypzZwQuECnZXqFhcOwx323ufJ8DadwrQDsTnJdTFHdFu4XLh32qkOBkp2EQk8GM
Z4JDR0zohDQoVHoDusYxN4USPdB23uJEmEx+DmhdGnWOzIKgHPZa42LSR4x/+77mbo1oSg+NBAcr
OenrCjXXSp2DMkVob+thwu8ekuP9KePG92I5i5Hx+qquIJUlDdBiqXwBiTi3AaLLi+VzYX2H64yi
3ITMaRUBJtSbT4H2K3Ofd2yW+YOhODig64VZJfE9wWHVAG9pg6iVahHJSakDEBUtCXSaU0h1/Cex
plZcvYrWtqehOYJoS9nddRS+A6PvSd3gRocx8mucIC3H2DigHHFmgGfm3yQg2CY6iOwIQK1AeB6D
UAOtL/me6hukt0VOyri8tFg2Ao1iIoXwcRTh2g88NylBxjO2RMyivhsa2DArLixpxv5mn3npV9V7
hA/LYyqNiIeZtVHeckURCXOfBU9ARA8Vn4qCUT+WaMdBrgux3mmuT+/El43UxBeEIvrRWJ3t58vD
+dyVyH/XRs8HlteH3NAxuvrD7+y/C9kQGHCHRm/M54vF/PfXbft12bAt9iLFhpde4sl71vz7WNVZ
iBpWN6qtkuY56L8pvCqH6tGS3cUy5sErMc+2aGIIVotkm+g5voB2GYATYE2DGFz4c890j8UePk8k
oaKKjdr2+mcSEF3bltOasIm6sw0EsRxohu1LGlSrp+Idm7H9Bvbab9fu39GEBJvWjjyBPOfa97uA
e3yWOTq4kD9lJW17ryMuswwLSC2O+uOlZDkwJmzq5olxANUlpdPfMYAZTB+Jg30iMnZfAPx4gAp+
tjydVse3TUtTEkh4qiU0wZvwzDnL8KudB7wwgJrt7nkjSd4ArUdyugvcL5kf7HWe+L+HPiMMYO/F
HLotvUyA/CF53FdSRyvZ5/Usjqc7Afy3GxjW/8gy2N3mjN86/8rjPVJYbrClqtf9/DRQTxYJUiGY
vp+opZ8wwbVfLaZYdTZXGgdSX3BdRpR55geUWB/mAGCOZRZ2PJcpZl+93uGQwLotQoIdvDCsWMGu
pLPj4y9eyQBkpatWQ+sKCaT1PNHSY9UHQChcp8w79am/+HZ0dxYZnsT6x5IqikgN2jPyUcHAlRXW
nGsuyQIqP6L6qq38fyjhdRBgwsH2lVrKpmTmnntqMG/rICy53ql6pSjqiEKIhlVI/LnyRdWtvh2v
e1wfaBuk/vwFplaOzQTECVR016+o878PiAbgYoj5iyRzxnf2hdVHve52VY9b6fIxGyXtUzbmFKAN
+DYo2HV/ewJXtsDJ/BaI4ppv/CrBEweON53RIxY64uz47O44mKo25UzJgxOnoA3ciJxqWcuihUNY
O1Stbe4CtVq/ycfgCJugMLRbmjb4HxLWW6UnvASDr03WDZaHaUFAcEgbxj3HbEvJpdpf5RHF3XJs
yzhft+l0bxXbT0RCdmakkTuj27b+Sc9G3PWsSd1mUyE9kRucZtHye94AKe896d0xhIOPlpcQp2bw
Wa3qKSUNFNOLj3R5Vs5rMKfwPRXWqcX8f1A0HDoCJTYUYoUlDjmlWg7elZFx1AGDYeqjWa80m+hJ
whsa2PMNCnTdHWpW3PSOpGRCKIZ6OyOxNipCX8jAih5iOITAmdvYmUsCzj84mzufXr354Wj4p7Li
af4LZFDc49kYFL+GaN71phB16xA0ZZ8fKvRLt3teCg5IDAiFwcMbuhQGq9e4KK7OiNwW3NJDeIIg
zVfoNNH+BWSnKxMqLxEtxe4cQfPeUDuu0jIvsu7TIJQpbP6oC4qdfoQ5NXx0alvUy4eNmghOM88o
V70BBNz53iNkTngu4lrDvCg1MWrpQSFuSoyA71MdWg9D05rTNPx6aWbm5tZgiFMSXLMPUgNgrKsc
0TbD87HD5Bm5PQxLlRVGqTvrnWueDyDfbJnZ2Ru3KRYH9jWorT80QH5LmkCHAmonqCR11OIhDZcR
JZI+sPaBhnwkwYmwNXcBH1VMrUNapLeAxr61wZq/tOGCSSREHFyqCOfwhue6r2spznn1NC9pRcry
/UcUMIQo/8Rfv4K6SnpIL8ZPZKZ9zNAKUH38DlMM/gbPvaXay+x2HZde1r0G5slImp1WKZM+ogOc
T0aIvga1Io7PHp0Nunp/Y49/1cSVrzTALObGQm1JM3RFl5feAacql9dSVoRhtzzuISELmZWJJukT
XPvLIYGFLfVTidhws+GQiE2uyobfR0sYAmz4Cr+oYoCbVGInL+fhdDHUlxwk8hu5bCh3Q+3Hixsw
kN0WXSmlRC7Rxq1ZtBF6zoAUcl2uT/A8kWEXOOxvDTpQ8+VTwLns1x1W+osY9Jb65mkAQSYg5UBf
EGVjJc0ojSVmaCiMh8jzGI/QKdy4FBLFGDQQsF4xzeUyeRPIkcPULsf3N0OVEPydMMOtrGhOGAh/
+tOmD+A1NCFiUKkdmhBMyB2Pv2mkkRXQJFD1C354dI+W7Isd5NOut6wdMgw3UndlwePSeXsK5cYt
kQFjIviegGS1+DbzyqnpkxExeQkAD5q8ICGfyF5belof+MwfPIeOXSgVnv0IbFcPL2U4CQaIUJSm
jf8hjZE/nivSr/NjOgazVKjRPNCSGf8iciRj7BbmZAcZL/087fI5+g1ZPtZ9Nuxd7DgoxQyEOOcT
hTLhFI5LHbsZK1+gCtSPTpxSN5bNkT+M+/aXrlxar/OhDIaEeMyYFhcEO36++vPu1PtrqOuBd7WO
BT0EacGMECF5T4rnwnOd68xb9hIsV5+XirXN52h1t4JbRMSc34YhTtFdAST70XNqeyITuxmzTUMU
T/c/icMecYSz1/DcYexrEVFWpnRMCOjOcUD8NiuDHaXxP/ifsyDWRFY70HB3EViiuQcbSv3WRTwf
Ed9d318n+NEf72+5hUcn5FtIpUKOROoo65xg/4F7e82wLlldbK6O8uSxvWCeygdRWt6JL+TXVrAZ
56X/3BEQIfHK8pXdlmeHXgJZ7mz51BPu844+lQRcJLiQ/jrseDXdDDFwTlq67Qzc6uclb4JLTD8D
2rAteBkgOfXU5FYy+Z2OJz/wcd+0PAbgsZ7uYZZ1jHmM6hP7Ed1cYnaXHLpqlqOFK5FQuSqe9m3r
e0dElf6Aoe5+a+vBjHUQ10IPnTUC/tmY2zkx70wjcyiwTkmOT/sO6Uy+oUFw2XAx7vseYXR0jv8+
kJKz9tcs6+zvuuvx3Y/LmOUcX1RsONAZJ+v3xiSE6MQsAaXw42EqkPYLBKajSV/tesA4NPXZEtmY
LFV+DrGuTd5BwYxU2IYDsDsAHOgssKt63ttrCBxJxNTycfEf+CaSmjbH4IrP4pk/kkwuup0jnnem
oQYufDR65QJ4k/MpWKuvtHanr1edYoYGgd4G8LsiRm4H84Z9nC3siy4Zg7w4L6CqcIIJZThtRz0W
H7FMCRRgdD7Hazh1/nDgJsdD1ZWIA08r6IqX8KAO/IeIhGzFNF/ttk3r5TUnuQzgRj4EyUX+GWst
+1rTd6MJ12UDxUs9ILy6EqwwGBpTBtGjaVVk9C0e1FpQRrTduRZzHP1KZqRK12ABOK1CmjiBFFWu
5aDr+SoV/kRREMMAuL7jbuc4uYOoVO3GJyFwd68+iVmOvvXXYVi0knCHH6p3f7uVuMrss8nmLlU1
MOEXz5JkhcU0j3BJFfJIop14rIyKfgkdgFjbzFjgDwnglUzdMgIC7Pkc1ZNlcODbd0O6oMTS7qCW
1M+MJy+kMGph7O+/8cf9dKYz1J2FddhPN7IQ0c6hyYWsOOlkVeOQhk3kH/IQPKOYtLHQpBbBOP1t
hN7MXcT0i9xXAKAGIzXJ2Pkbh5l+qmE9aWSNoEWdGg0QJ6s7hLzuVGCaJej+0NF1mJUd+VVgzshR
P4J0DOvCy6LcVefh/pQr/ig8jmBg4+OFysH39qu6Kz2m76odRxcg5lorqMolwBvNjZiUpRQl4Vef
gERkodQv0zNCmvolpxNrKIibh4MMKHO6l9SpoZagXxSxPNrcM6nC8oL7dFpr5VcWvYOCb6zcuFJH
UrrnTFBDLqpOtIcTAcBsJo/zdti+zPHhO5oZ1vML85XYd1RIqCCt/UL7zVcy4BUAvy/Tkc9Dy+3p
dt5ik+6B8E56NUPiH4voI+tS8+SLr4sremMN1hUkgIYDLcGsEPEPZU7pLrJRmWxbhB6vOXwNmTuG
H8F+u+myhI6bkjliZurrCwLblRhMQnhtviJsLDtoBxHaS60i1ZoOZpyZR64nRUWlb8yYNJ9i1TCe
GZ87m2hsmI/c9/D4SFlWwzHvgUtmZQ+C4DSDey+Xw68eoBZ/XWgIrZLmGla7Bod2RUC6/k1A75kx
U5eGSHBtbjWZfNwzp24C7rd0lSL31KQfsnpFRYXJNojejU4EwH0FXLIC5uSMhYjCbWPrxpfmNE2f
UwF+FOGsZbxoKtntes3STMVC5iWobQup+D/B86DLHtqMF8Vyto+aAXdLlUuBcYHmjW9L6mQlr02u
6M8AzhGu129Ky/jLIkC42ZU/Csjmom/gXWN5vCQ7xh7zHu1owIw1qyC7/awAvUvd9wGCvGYf7MsH
HLWsORgL20P+Uofmd9Ruw+m6R0trFgGmOL264T9l1wnDL/pQ8xGeOqw9lWSG6cEDhHVeKSBUMZ5C
V3cZYATSL0gzx9jpCUV+B9jSjJ5DgywfeFGOpknIcusLuvlDYt+MQV8YRKmZvvSfm2QHGKA+2E3N
4LfyvS3EBVim3GHjxgTqryWmQYrYVDj5VNNjMORIbs2FSVP85u66XuxFNQMsbtNs5fQMCQTt4chZ
ztj7YCoNSZHQk023OzgHrZG0WGRQPmV7s7/OFxVXmAmDUiVONzKRXxoFB/L2wDm/tgC32O9ptAzX
EjaYW91dORb10CCpC1gFtlcD2yeMj2glDFVJlUgRzHThSOPQh12hNZuwj5aP3FUkO43TQ2D6d3Im
+gevq6oUYmoB0L/HvySgS0+jQbi+klK0wz/yiIVQHkwje40zxRQEGzR3y7gKHs8Qa/1RhDf/D17Q
CJ1osYoCpuLW2uoogJVykyskMVE7E30SqwihjzwvIK0TR6dVEmBUOL6msostjvSIeAlpJSjbPjVi
N4DHm5sSm9qSeoWzrVJVrgviBnLCaHtMDGQfZuMcLOs53RFgqFPwSCfmqmWOTVZXYorhfPg9hCY9
3NvNyp5dZTOnae3wN5oBWKZwJ+2DsgDeKSOHOoZhFKbm2Jo1AcmJzOyyIPU9+XsATt3xVGa5Ru7J
7sZxAaMB6CXSFom8F6/9Q8r1CZdaBs0xc4r68XYYCgzrzmsEd6bzxoS6tBt5YCKMBE67KhONBEie
kfzaPWCN36u2lPqdJtx9qBG6saaeyCxZz8AsbqdgZV7+/EhyiJQg2ksZDn25O4FBOiUzb0aEUJ/o
uMIMt0zQHkX6Ihlbkn2Y6qM4VBPzDNakvv5QBtvUsAplIXlxCG5FV7+Qo/1RWfkiEKSOk31hG3m7
kciRo5QLKw1Y/StmqXn1P3HddwY4D2C52cERQXpQBuepK/mCeZ+i6UzMa+RTfge229oKq+wmZoSG
Av/NaWarIciFfcJhWNl8Qc4DCoOHBuGDzCm6pj9dN5Kc/rVmKmZQNUllO+41k2EidXk51Fru+E7J
wVX7saKSofle1nFpn7ALNtcDEwqqNOyu1m8bTr0jWZi+BPcN7j9xLgJOUFZMcQCrSEcC1lflGvhU
HI0YtOYCkGp9NvJTBgqtoYqkzndXRA7w8BmlxjeV+xYN8aK/G3Vl3Pu3kLmxbNy2p6Pzdz+DrSzc
f8B5H28t1LZ4FXCgeuHYZ+MSXrWs4gF3QP199lx/bgoyu28WKrFaNaAEynp56kmcmhW8/+5B0Ngp
BpmboIJRYVG0witRUedS4/SZraxPPcztgbkVmeBZp1AVxvTlu81iOhzQxFuPRDjs7exGTkDsSwPY
mgzidS2HGT+m1N9rccP0bY+BxRnPJwDv589RpCbi67EaAZbtGMVnsOV2zwiXeWhdU6q5Lsak/JmO
QTikkAhCYdWeiXSk4n+8AJc4U53EnAlHXolpqxv59icJLJ8Twd3UR50tQwOxNh1s+BtfOTTlgXdU
n1zscwepAHamXAhN/WxyqqxwMxL4VOep3Yg16Lw1X8BSm16RBR3WKVzHUdZvSt3XbTs9uoba3XCG
6fDYbGIA0S5ZRqj0lTq335WqERCAAt3+W6D9m+M6M1HVbj41MoXKQ82lFLddA3JtrOQeFAoJ18od
yINo5aGrX5YfRj/cFGlCVhxJsOx4pEzB9WHRIafacaB/Ai5P36g536eVMGqNl5hqpr8vrriGzX96
3oRqCftkufFOG5stdZGiVOPefrodWV5dQTmeooK+foGCsyjESXioiC6+b80JaNwc664Dh8REGfDp
bRsP/QgyiRyqMw3e9MdKCAPkqjLUrs3UB6azUYGcXVs2j73UYgamHxj93zosN+YQfvoTe7+X0XzD
aj7qmq+BmeU6+Ltxi1tdtsaHPSAA3AeQlGrrAMGuUGvpvIi1ODf9dNscvWO6wkSJMKjpveUTxAr2
r+ulDeb5lRW+/scF39Rube3x6vSJwZFtsY3nxBQXGnU7SgShNSCt2BJjx25AR1rxNZqwmWVOrNGq
/GEIWo4AYFGPcd2gLM/TrZilKNhkWvsNV5ojkcrmYWR5G5LouL2c94jGIKudzK3ZZ7cjry25N4Fm
G0XmF+1z/PJTXD04TYMvzzQ41MsUmuzPbLvSHvHI/Rq+dpR//vP3nCbF61d6yu0AHhLuKmDjRfEt
bBUQiWGzz9b8VL7f75OfkBu/U/Tp6r7M9wwJmDMeM0GR2nqLZMo+AL1WAeWA5EHc2dbm9+5vvsRW
mG6S8e6HDveD+ZwKk1EE++qSrayaM+QdbdCu92iQ0dbWjgt6Jd+KIM9/9Y+Fo17TTH5N6WOPVT53
dMsgb20RzD8SPTKJqEHtQpVcEXrVH5mMZeFdnXwjm7XkKhCxV51Wxs+HhJgCcXVa6lDjJwN6xGTT
wLzBFF6X86ZuY/rVTvrlmWvQMYsNrTJ846IfGlmVN/ktsLpgCwVoGYSuVGIb+iJodi3k/iK02neo
fdOgnplIk7kW3TvtFOIrc9z9jsECoZIyHVj90cRRjnKh5aJpluQ2O4vYCrcAf9Cpep01qzdNA2V5
O5N8chvB94ub/i6D+xaDXWvns+AY84igB++PJA698px2WkHncF4JAlDNFUGvaqVrJfHoHwxqaQjx
AOOim3OjW3/hzNPKd4TWyIpv5xCk9oRGhSkcYMfN4oAIoOZAO1J6Cc3aTA3BYBM0ocnKZMfBhDqQ
5IJTLjOV+kZ57p8INO56O7/657376lADNCjEvx94l8pkV65gg4eI7dVvaQS2zcQSKHcnuCISDdyE
q3Ortg0smL1+q9Hh9UBfQzGTaT9dgVvC+40astRX2yuNP9LF8KCn2CUTQHUiHysw7VXuLHJIleEV
pmRdYOaMSgheRb+BqT5MUA8LG7xHhkRTIJTF5SCp5k/C6eWKxCTI5PgYKQoPs38Ucx4LHwYRfNto
pNcxpBVJDkHQfP0vpnQzUkurMpJpIkHbpYDXexeMsJvgICncRi4SvOyAIbz9LkLfSaic29u4PhlP
o/ltVEUJqtLao4vXDqxTVEzoQssrmQ9Z1Jirs5/bBSJyUIqw8NGd7RghAMs4Mz1WzRmormsW/HzE
C4GlIidtQog3EpccqhRZ9DNVcigys2Qyy0GHeBo2qrrjikqdq4U6GPCuladZ0FLoo7Qk8s1WAgfH
d/tnWA8HExAA2TqX/iGXmYXVmPWJGxIrBQdjAsdW/EjhxmnNjYbLwhfblx4iBnQQahM+UPoySip0
zuwIyrOzXhdOWcu7eBGdFkv1zubU6/AensPXEvPYZKKTlbVBVbCHscU1hxxyXlI6VlnTCSIHya8v
s1InBuszQsQcvxqpNbv33R/AFgsfNzgSAXOhsNAFrUA9IfvRy+e7YJ9Irkqtz4+A3F16gI5pja9L
NZ97JjQRED020ZpehRASpjM3MD48GfpY+/7EET3wxDa+5A5uDfqTJ7aWVB7CCWofsAl/IwvF8jKd
uNe4PbDlmVkfW90obuxZ06VoZjMVt9K3TuXPRNRN5nxw90k2QCGWgNfwd37AQRXvTw3IiHIP5fIl
lJrEJvjPze7OrDjUAgOo5iH6+vWrhaRSUgH/qq19MpNkQxzeNQNLasygq2TULMtdmgfP9kpJIbAS
N0IF9qYZA3OurP5tEEuDvjz+243QiS9oSmJohRW76AChZ1Efr6mzspyh1zdWewRDTnctx1yqRZAi
EIcx/6yfLrF+o/CCQt382L3oFH5ztB0mfFSFa9WEEnjcvdPOpoh/+odRvgjFnE8RfcjNIfQpopFy
kR6k9iopCpwN6mgsOe18dsQePhLMhv6CdIbKewSB6bHI5S+E8ay+gOzu6u/LoZIMFGzzmcPGlFph
ddFxbOaaVxtHGLN8wKZqmrW0WoPPSP0DTXfApqiIDy4SKI0PG/YgzoZqi5MMaO9Urf1EHL/IyH00
yUALIpoSgj0bm/i18etXHlHYiZv+jcJ8KLiHfDiMlQX007aH3Br1qv3JVXn8x7XhY6YuXhbA/RCl
eRK25TwI0bpf49IszalXJQuQ8w0P36haMBgRRbIP12FhcFb1AZ6OF3mRMJ+MchKfjJsBDT8WCyvY
Ho/V/a/5UfqmKS+tlp231641SguSU3ilzBvjyvQM1ENsDwHkRHitSO6VIKnNkB6o24UnHWns63I5
6GhEbB7K9r7lq6gt7udfUZRT4paKpZoSM3vAv1nul2lakzepe6F1pN0qtUbDyjZlp/G2NAhAmSho
RkKfJViUdVk7UtL9J+WABio67DqoxcClyACoyFMKOxKRYLsONPIWcIo+U4UFQ2ZYoCMxWl+onAI+
slYezK6mX3G3vXGQLJAxxsfWBnDgYMTk12Qge7s9coKxVDvgj+/l7VauPOF/AuglI3e5t5iIUj6f
x+5i/t2LlDOZLhJycGSyExlNzqBHjEG4hPXplH+BrwZ+iWf2zyxcDAXfRTDSAzvJ2oZOi6+bkMNc
OA69s7kafRC6+2HJ6i2jrfBZ84aFTDIJSn9OglCmmGoqC91hvqFl2Ga6nRnbdXVnE5Njdzbhze66
cPvrAY5Gu+4z4aexnsJ7idnByMWh9MG1UgROgYSNrttF6nVHZ5u7ZqHj87iJBdkrlv56cQG15rOl
r7J5BjjQlmWytuks8mv4F0EEKsXUubr3kAMBfdn2gepmuWdcOnFzwXqZxbzXocOntnYur9DoqtE4
ZfxDlwBsh11ulwpX4AknIn4535Ts+drtEicRWZP5XSKWCNzcX8UzVebq4Lttl5i893jFL79E1leE
K1JXfxxwqEkRkxppoKne1NwGK0sGaqoSpGiErx+jxEnhlR1hD33uZvoPphOjRrHWq6jJdqFfJoMV
qsM8Y8XHbLzruyqPTqJgPF5KRRqZ6tH9Txq4rJJKytARwKWW/A0eeB22Dy1YU0j3wzKvI+7NW8Mq
Ot03SUi+zF4z2Wj7KnwJmarmtYXIWAFpLUIjhR9R9rfxpLC6xX+V8mfuGpAXnz60hdOajdYD8hWM
zIs8pwPkjLljaTIMoyXPU6BGeeZ13MBYdlgMZuNbunaL3EWHOI1WIc7bjzOSQ0fMyBvJI92M6Ntn
/Kv0p8JJMpWT3nkZzq+me+b1ff09kmhjD8vzcs7O+UB+RB/35J8MbFxv6ux5R3qF2peqXu14SKlM
VlcbFUR0L6r5hpAvL6L1XM+xwroFnbKKVIEw8rwNQlbboeM4EC3HtA+dN1jJOLUndDgKyYTzZAq/
agjD99Vd9rPdrqvcKYUVX9yhaTPR+Tzkim+9ZPwIXkqcj/hRh6ZrlKLwLeHXbZeGhaPQXXfhkaLY
/07cVxkZElMSaRf/aOrqBnwJenGqk7hTlzZY9eiu9bVNvBRXhOp/GPtQZAqKuqUDugV2qZx7ZWq/
H/OOpPWjLGhwzQ2H9udlP4kaJ92XkkNki64Iif45ZCnnRq78efDIMv4mgBOnm+RjDU04wzEF9esz
rJHm3A8uxscv8XDuXVu21tCgOPtC2LgyVc2ZrWu87b+4hRqorz6l7cMY95EorpuAU8MAoUkWr1u5
On2wCHr7vMZeK3060g7LuanTK0g68rGz9NGQ+qTLHK3CKTu7FuNyWghIWa6fN+bu713tCxYOoumI
j/kEPk81Gx5W9I6MH7FDSdxZUrVK9vYEybO0e0VBEZjN0hNiGFx0Y1AfimMVjhzzq/wGD4QvW9Hw
YxOeMZSzUfI0SP9BtBu4A7YHpfURLLjvp9LPy/nzPFHi3cF2FeVEYnVLvi/otgJnp+9iN/3PLdgh
ZXCBDg6mwpngSc7QQymbp8Cp80hyRPUncPPy8kbr5C3fHIx5aQavqJXWK1BT2jtSVxr7cws+Ez44
mfwVBXNTaI9wAwtGiusObVLa2pnju1fqce0fIxSdXyYDV/QpS41boFsYLcgE9mok2YjNvg6/i/Ol
fXmLXoVi6aUc93DeIEaQz973qvz7+VOCjVBy6K9TGEGo6S6266KhG+a5n/OPiMvJKd8Kc8TmgNLj
IKCKZ2XiJ0pkNibGYPVxjS/vw9ZBMDrL/UYs9wzJ3wMz9ZQGz1DPDtZYaotV3t5NbxKkPmAw4X2B
MJW6fGwLwi1aKyJceNjqSgfC8vlPnk3TG+86WZ4Fsyl/PYKvSRskTOZDDnsExGjyD/7bW8HL4Hy0
ub+SC7EZf3XpVyefdFC37epVwY5jkHrANujyNhtkzbHuRzNUohV8wjav7cBMx5RN2nofBpW+tvnA
XPkORWIgmHnL42NNp6u7C3PmsAVDYkv1KeSni/MFjR5z8/wh5y3JreE/KuXCqo1U0aPofHt/Ifb1
uKjGc+Ry4pvLzO6iT4CJSGTWA42rPJJr/Vy/Cc3FpBxfM9u6IfFvCjcLk+RMgZBxAtD5l8HK7cja
/kcUjEIJU9j8CzxpNUX0ZXdsk+AzxRu+gfIJ1Blmri/FqzP0SJWiQ6HV4OZZFtmyf1LhnhWneEtn
jz4HjmimdVwGZTxHeJWyv+KqU4dbXgGDqoEqSw95crsGHNhkjzcB7CMSxKLopx+rKCt2q7gfxLW9
0jKg8SgOEqHfOgFNcczgJa2W37mIdsH7yU856vM+UbUKUoJSYutGhmJ3CPc+CwxQI7CxlpBVb+g7
Th2ZLbBHR+DtJeC3T6UK1ZDSE90ntwww4XQgZf3Ou5O+aN8lLaEuCYywUvg2qgTJzs0qwb5Gqw0P
YmSq0mcDPGz6ArDY80rbadB0UIGZtDD+lmvNGFBCWVtdUtXdDtO4y8jvTNbrSaLK0OK/P6/oMB0b
dW2THg891XR+euB7edlm11c/1dY9CYWM+1pYoGXsheEOjQjklsuGGIrBlBVbGeIGPoby31DlxOTl
DZDnjA7aU7Xo94/Vl5g0uxXES1tXkozkc6hU0KiW5JDR5DZ9raaZ4Jcxs+3dCehXczZs6HhkTWxQ
vGSdgXmA8w1GTRP2U29j0ZyNeEKKDj21zdG6Cdrn9aBcj0TItOJWO4PF/XBWdNIK/hEYn4LzGceE
DoLk4baf50fb29gzOUsX/EdGdqsPS2eo5MeKWh17e9f5Qy5IhCUGaqM+YlZ9vOmH0uuIR8/k3VOg
+fHY9ZhbkIjRVRDGjgFa4FfF86RL3dfXPUx1TTwG8eN4ErXM5wsRMCU0ZeGdZOQDZE0UQLOTSjMl
kqcl0JTa4rG67Tje1/0YULpuY6+/5nAAZyHlsxjR8s4cxds2Usm3Kg6U0JtiwZTVIkWYDMj12oFS
Hs3h4EbjQCgJyLwKr04c4EuwL9CNA2cTJBB5EyifayV5ZNGWXd7oQPrdszudBtpDOcrFQ1T134TU
3L+0uKizuzXbetRlSHHThUYTw6yHv0KpTRkCWLcCeAHEopsWQrRLbOr8N60ujnCml/AATuuDFYnH
x7PSXKjqM6Eot4Q0lIf5tJTKQIBcU6ILUGfAqrDNYdXZA6JQWaPuLUkbL7kLMmqq404/5qhpcunu
ZSdsvcyxXb0xWemft4zsLnYdQG54fH7QqH7C8XeAx75p2RzcDPCK6fv/uhclfJL3shIpa10gKASQ
6LCSYve9HoCI44BBvleXWo5PQly4m0sDyX5b/4oE5dVAktdPz2QXNQbT0q0QH3oS4xY23l+a8W9f
NHKnzCCA2/4iAUgj3gVlBPho5HZb1JHzjrf7ewMIiQrgpakpIUr/snQQW2/K6uMIrT+LQqUTI4dz
keKixDAoCO8fbGKZp3PwQ9dXkiQB7lRgdLRmCvQvAS5JhrIekEl8naB6yxV46f1K+49DxP8fMp2D
GdLUqhje9o8Wtr6U83YjFk6+GFbBl+CxL0Pa48PGw5t/hbqNAGoh3RS8Q7tfb4Ly+V/E7vPkastf
1DUScabOpfUd+KXXv9XvIzpc8ffEmJtmN8CQr60PRFre/y1H38K4mrMUxaZFn+xVz5MxDF3e5TY7
fpM7lJnCJAHIbQTQIr15Ce2wPOKtgSl/9+h/QD+aUbyQycaWcglLiZDgtoiFgTbLoGAcBV6bxlvY
8X3kUyqgCkf4PkEQ7ujqHXDAAw7X+g7z7UNhxcH5dKnDzSeCI5Cfs9a3f9sZolfCtDZXS8rGeedO
uaImpWXISWIt5gS13Z03kxez7cyTsrA4pvuFYVxAn1aL27t6hmrUgcxE2MmAoeHKCujVFToZZKxV
W8ZY8UXBw/HAXTkhQnZ1g53KlDRkIdovkfQMH829PwsoQ+gHsuknP3Y4qihKExqnjPrfI5PvhXEb
C0FUaSCirwa1lV7AD7UnQ/DBTP5/Xopcirs7/T3yIWcQE+FFEQeHDLfVS/tyXM/WfyCeFA8QMHvP
R5eosAkRiEcml4fbE2iUaFhE7Yf4mbjf13/750ueH1bDSn8XQaIx9zDQTX14XKrjXawZgkzsKR3V
XyxYtAeCLf2wQiGOAssmVCgrUMCPArhJyUPCcxRoVgMrYz+GOLUrpg36O7BBqrkzj/A1S012YIhh
j+o4ZF5NcoSabfqaiYIjdAvA18RpZQHKwj1F/06HZRFCx4N8n4g0r/XDEj0LCgXAlL1ElXoEgJxU
ic4Lt//CKGaU5e0XBj1UpuKpwcvyKxW3mEdC9OMuwXaJAvKUX68Tu/ZjSbUIEsGhErkSG0Z42FoT
j3+MED/EUnQDUjUEk34HnXZhOH+x2ozpXfJxae/sp10hw7OqMtHGRcmKd6Xkwh+znbk/E3ns3/OT
JGY3mUBcD86b1EL0DtbIRAO/lfXf8vRHSN6wcbF+rmUV8gnOWPxbctxg5Hepzyt7poJ1/KWhw5G8
cu+TaG8/AjZwsiV2QX098dhfWBU/zkB0khEnZ+s2QgNHdYCUBRNDpC/YG+zkj1S0YOrF8O1ISMzO
jXoYr9uJMAagP8QXzyX+iXP/XMc6U6Bi59c1gIdP0XCd2FkqZwnXPikiQJKoPztqk26HPQu6y/n5
QhvPG9dMgPpVPctRHouox64nlWznxQIwitIOwRKpcJhpbr2P99qHDtBcVAh4ffN9LSVsKshJ7IcB
1FBh5PYLDszqi3s7vLbkm2TmMKtQL/T6ijxbfQoWWlCYr80Lea0VwNX0ilDyDWtXl8KfuqfUtcyh
lzQxBfDAV7JypRIr09HGtQvXEIml97rgobNxXbUPetAgzCJYBXxQWmoYl3VLOM0GIU8L1q5ldXJ4
+oVrBk5VvajqtCx1L/tTprytRC2dgDDG8Mir1Pbb+2d08Xs73eyUN+SrdWO2otut/UwQmoLogO1/
bOpfFtsZ2eKQVQYiWOY75C7+sIJkVQPuLQLLTqyMwYAVMPXgWzkwS1SEzYAgmLlfioFFLok7vwa+
NOKl6MHCQlL4E+yuVc0LMAvXXJij56PubtsSWCJprlLpqHxiRfmcNrd2f6nJf1Hf2Ep12G7vGMfq
HlUBGCgJmt56unxx+fCW1bPT33fzfkkB1G+jDhbzWVz8HkOgzSOv/lvGfTzYQSaGigCP1z/gxXAr
eHBq3fx5rkmVqLu9lufAxzLYeu2JcZUAEoAz4auMJ1gzTmuPiHK35aDwvjIHIUYPtC8t69LDlSbP
McrdiIDX1uIY2YrHatLHGQ3ynuOUcvTbXqdCMxq/Y3QGGw0dlpW7z9h4lsMn14RJpEev1iUHCibr
zxXk88nCCOkfHikQHMtBHwYJcKS1nQnFpEZY498McxnypJr3UADJMC3gncNBSSEFOkCJhcWnE8g1
ir+K2EaG9oFvK8KTWUhziM0xP+H8UKQv0tVOyO1s2M1v9teVlYDNoCeUDpST6+llu6zwoiRG1YsU
b6/OZPNUoIrNCn90DyuR9EO94MpN8drrOd0Y4uYAjLki1eswybv9/Kt4Ru8YslErG+62uRoFLTIi
jlUbHHxLOVBWH7jfsc2BZYIeE5AWjjMQqGD7TDJNP9X3kwBua5+ZFa9aos7CHSKL62pMw2H9UyOh
8XdYWUVKZcgMvqrLnPFa/ycqe9yaUzCk64Ha8OIoFP8J87tY5lpmiuLu++68YGSxjdhq3rZZs4QM
QRj3c7dCgwhpYTOd8FoVLzo+g7hEaGsfQD0uMg6Ul6xNj4R4Lbl5sepuEOgutStCvHlMWGNX+q2B
NkdTvvjRQiLLM3LCKaOt9KKcrmLB9LNBgybzyv0Uf2mFgR8gH2SWCCr1h58yRnn6ScJB3aR3eXmc
88IRfZw6zXeO3EFf1/fqRPGCrm2yP/WHuYCx+9SNTlO//LaTtypSF+plcEmIHoLA6o1m66yaJv0t
mq19MqH2EabDkoz4b0/scQnupbGo1qWpkybol+BBYT5SNnzj0Fl/nRIvnIwcAfYR2a1rLUFHjAPv
Nz9PUYHuLhZ5CrY2JY4NNW4rtpG+oQErdRdDQPKvm957jwgdDBPlvcY5zy6sLMzqdSe377t8BicJ
0Ar1TAtdcGiBMlodA0R2BlnrlqnRUvpuJO4wS4Bs8AfSUkRwBH+XEIeJIwK/0i0GJujGydaabZcX
8pQW6K2krhGRqhI4Kl38chVlXYc3mPp0hbT8nOFaecmKquEoe7DS+NtN39Ljm5ylpm/YNodrTMBW
UhT6hDzila2BSetMT3lmWxOucqk+2BDqEUt0FWHpL6HnHGSVGZWyMEY8hEos/qffUVASTK5P1j6o
N6eVyCUHX2y8xWSUPwR/vU0khDA+BhAacSvHBkOnhuOMczc8fJYFP1K+vz5AvEJatsM1biV03nwT
scOkLwN0B59Fx8CzlcuTqPU+uw19s+0fNv1cWiaPJnvaqI56AvtjqJfFeGVtQCQxu7Ex8LtNeOdj
U9mOYRTULurHJe/HPBtIR7ovwfAYXqifX46Kh19K8mbPhu1PcPNSFIlUuVWiffZj1f4v6WbimVtt
YPppewL3hKSztAYO6SjamRlnRFtzaQf9FxHokBnbaAoNeoXxyAZhy01VJ+cFPuoETafxBG+3NUVc
arlF7WECfOUf+e3hdEjfjBnobrwYXVYI4N99GtGm/6tUAI1bhr3c98f40jVsUjuIUlZzcFEPmhju
BvC2xYSA5+lnPGpESA956Q+dF1H2Ezpr5vppo5GGjCcJZY0NJhNSEuG9W+YyM8ub2mMlsq+kujAq
iGL+OU2l1mT1+EIUDIxkzC3tGVqU1q+2H7VkV0a3uU8+hQ2zWvO1GyrD7ojdTDDH0MeROtPuXSiC
DiZvpJ93w6bbM7yR5ffJXRpYqdi7a7czTqd4vIverIR/K38jH2JWvSL2Wosn/v1nWBa24IpCxcUe
bstS3w14r4zgkZzrGv90wIm1+EV8yNd6FRvu7MEmqP9OYLxOk+vUHxh09Jxk8eTMbXDNVEDyyReO
BJGyZ/GtfQXg9iS0lFd0GM/RX88V7g8jyyjKPsH+UpSBOqc0L/8vw9yTSxeErSYlcyjcjncjFgNe
aYjK24BLiAMl4Bkwt7B4z7XAGh7WAEkgctsXT2PUw6KJHttRQVvkSBPsEcuZHCajw8JRUmxKNT3f
T8BmQIRe6Mii9zFMAQuF3YQ7yKF92byUcXrKE8dPYuED98UIDgbMKhkiuEfAi40ePuskyuDsOV0J
pvnyuYbDptHBPmTAHWGCXngCPtL1EdQENiDSkzzVjngLWvByO4bos1xBKqvrnmpBIEwKizzsEryc
W/kZnGLzPD4tVNSznaN8fNdhk6xLoXvsfTgEFXWbe90yb2U8lRj48ALrvn+xEyBjq/UUoNp8+5O7
k9HE32rhfjpa8u/xC3XJT7r+iotahAfAysiGzL2o9r94DEEyOyUPGdFdFKE+q6n4PdN1zkVNRi75
oenJrUuqOjpPfTolnBBLnyJSOltRR7Uf0taJK/4O0Py0M1ofy+NXn9b6bU+UFoW0jdrvM2s22rQP
2MtO+ojUAFTbLv5uiehbL1NY9EQ3ntxIRDATuI93hHMC/hcsswho0/Xac/WiX3tT22WXg4xdN/9I
GtGfdfpjSB/b8vtCLgSDssyX1fp9PxI1JAZBW63M7Ldi8S2UPWnWdf35PlVxVniG/LO3ZKbfUnLu
a2+LNpcxFHP330uWJEP3f73AHrFQv3bruLle5FAkFsJ3NO+koJ9kSjITtOe95gHpqvLOX7soKSzD
X8GdTsPM+r6ffnlBQdnhZJ1pXhfw+qBqOSjUW18qJQ/HwR1DZsio3nZ3OvMyqLwfxdZ5Ou9L4cVQ
d70bE3YMwF1qhdakW5lso5TCCpzUPcBjBPliqRPtN3ZLpBpgJYHYuWEzWNOF/8IboFR7QKABvCVy
UVQDqtgXg5mC3PeYdACkU2MW5p2c35xIBl5Ql5iyTBWGl/7z4Y0JWPYPn0kTQoZF4jXTB7dwPQSH
qGfm/cLRsGs3lwZLgFLQtLE67M3ylvWun7YPY47stAM9fQNi8qc4UJwnUyeLeWXzkXwQ7KeZPfxj
ziZbAt1NjQSThXdIeGRzIsiIQB4zLmbXkFJvV8PWDjL7WMOa7xvlb0lNmw8ZcmVN+WJC7kuXCito
t2W/nsU8fF4tUZ42fkEFlHzY5EoE+Ut/q0nIkmB5pBsY79pCUJ93v9R24pBCD6coVO+wYfzBMCfp
9p6OrqxKssQP0bj6kGzR3ID322m/FDbKdTXf2RWqyk7DaV/rbqdorCRlGMYLpdiQ8EWBY2Po5WjD
1UWB7o1pP0PrJ3P4BHjdMGN1UHDzop2Ud6vlFDYSJfLWf4hvsqI0NPkjk2/aWtIPYh5ATMIsSUBU
jqWJGonIBM4O/nH2NkjB646J4DZdceP08m3Dj9p7xXQHZwU2UZGBNZc0o3PYjh7r+9RR5nIYk5P2
ySDGosunLpwRbAGyLZr/JOqWL85bj4sYwcIUaHYV5DuynMI5WofqPbpOeIx8OJLvbfeKqeiwtKNf
i+rfgn439Kj0UExm+22CY+3cjuszbf1KiM+DFbgYL9Anbcl2t9uNRNjAJsq5sU9u8YNdH3lDTqii
HB0IJpGqSYoa/2KEVUUGJGAT6JSv6bE4G8+y85dKrVwX318DpymUE4+K6ghjodk4S8HDPo05CN/p
CQbujtfpB6MmNzKMf0QlfNYt8M7CDgvJjfxRjoQG94V6+lSowtZ+KtZIAcfckBx7mOXLlIvQb7Et
lblzfM3GxGDC+37pV6UbSm6mEAIObzCN2ExHYjxYRIJNicB1NNI265e2sF3fQDOpYofvo56+iU4j
07YEkb/DMA5sg0Pjf+UDX961qjSGMw4L+lGFprv0beWDGmkDxMWcKOil0F+HZqYQiLvFJFyUPiUb
4LbytAm89vmh/rfMPjy8BsDwDuyYvspy66whOH3/pD+hVzz/WmbbmaunNm9UI9c5AeZ8aHytvy/u
5hCRX12C70KfT+BZoiudzo3g9/+mxKxaa2RbzpLnSTi3hCu7DoSxW98ayAolQ35NOFOET1fBjr+X
ACWDi3foJONH3O3pOYfIiqJAA44MTst20wtKtr9hUsHbYntTuhrCbxAbhsrctv+52P7Hf7d4f45F
0Ar0yTAVdUsisI78LSD1AYVX49NpfRGhitb8YqWd6acCAAu12t22nzACE4NsEvnwhRgC0cbJ/iAL
nZtlOCzdcZbwJL9SvvltGSwjaQlM6LLuJW/L8m2qDWbMq+6j5HNVRfNTUkgZKJYsWJnHXImGs2IB
8kKQ7stGCdlnNrCfjR4cq8t59rhwjd6MitvPzzDlCi33ELcal5kxfRyUtlNmbMt9EH1xhOGV3UHb
MEvGaRK04y/BoeyrM0iBAenHNrCRRFBpbc9ef6ME/h+Co7Ox2tvnB88oK2cAxPkJewE5fNqBUwKp
eUw7W6cSqsDV7GH2uwOebIo6W8A+KxFajwgy45Fev6QneZKFj+yssk9deG2KeS4OqluaCKke1K5G
3kPKH8vHcjr0pPhB2jrMnlvawIhi+jFhuYJBX/jh15dQ1nU2+g9m8BiQ9i3F4lKFQZWEeHlrZfEl
9SIk8pKCrtEV+xxhcJoJR2+gEryEZ5GDDVD26EdZVQkMVtqXj8oX9OSaraKapdnrr/s0JyPe2JSp
NhjEM6zV1ziOyMJcGdS0shtaFHTZM8Hy6T5fsysL5dPOoj8yagRZSGSE9hTZS+ELbiTC3aPa+Wum
16p2h2sjNkIMu1PUc4wBu+kZB6OFYLWZIICgMl3Sxc9ZTwQ67A6Su3puZlDDjs9clSJ7PrXrgxvU
S51LHNotFvp1emwpV1K0MxvJzjWBYSywhq9k6clNyg8yzTyXhWwwAcb2ttkP9mZJgV/fZjTpy4ic
alxaFvrKBz7Ko4fXul4yxRjUwGVTHPwwRyWPAWYZwosFWq8XxXTYc3WTsFMIu+irjFVzCW3Pp5FB
jguJp00McPd8Y1RdJOnrT+xjCTt0d5tmWpYXQEMXHaF+D0rQ37WgRojkgACJeugjkzwzsC3rnguV
k+vmkumUXPiKBhBesL69//kduNqKkpSFjU1KxhpDITYWr3GP4rTauxbZp090D6N0jEhi9WQJkAHG
/aR4xQ0yzUvIk+oda/5Z/6J4V66m8xsyRo+55aYAOlKWs74MDje+779afU+ydS8rLSRY5DT1Q30J
RmHQuiyYHFHl85vVtZ3QR3z7onyOIROyb5AaUEHmqFF+poByksQAlEyyiUT2TaQIkl1dm1BE/yoV
ADMgpgsq6LyynoJXcVERanwrsuGihWN7yGtkJvOGm0Z7V9ADSdXzzDnq++ydUv3RxC5jV78SITjB
h4faV4TVf/qjwZL+oK5fLkqUMP4wmxA+aZ2A/ZIgwEfCR/Aw01A27Y6HplYTM08/EgbxQanSGXcs
Lw2HCXM4AKuXYGVKurlZWGwwXjV/88oKzWimPfLdGQlkesSXvP5hn55MRlxyL6fpitxnbiCkLbk+
u+0kH92lvG1CgxqQ0jxqtx/rfu3HD/bzBHLsPVkKRAumr/xx5vfj55fjgSRP+/2ZutkGPHXujdNG
P/I0nke2H/o6kyXvqwnd09f8LkI7juc6ebHLHRZ5CKgt3f9p0CMUetwFSEWF+LW4rA/T1tN5Tfbs
b+oaeb8N+enMyFJCaIsJewaCvyeBstgSuDIcUy8WLdMnMeq1iAWEKQoqNX+q4QEinNpCc89inkne
gdJT6Dcp2cEPdfSYVqoaOzUXXv4v24EmgS/AD897/pldwtMejQu8v7OuJIxWZ+AEA/0EiIcOh+G3
pySt6Io7QWTBK6PeNtIaI/1R2eeMn+Rv5wx79XVs+TqvBwUyUYYU9jwRf9eTXkAdlaf5V+oQPiZ6
Pa1qXu9Zae3UZilAjePm4oYJV5R66HPK2hURnY4TUwwULR+E9KPH34+EhCYe2B8fE9zuCLpiLCnL
OTNEzKeneL8B/cGz2pcw1Ww3Of1Hi0nY8aaq4XqipkpdCl8I2hl9jpBvyQ04mdBmiiFta6SdDjZ8
57Um95vQb2MuhFAlL26cs7hGoFiwq8eCuO+F69TrHHGS0MLOxPPbOk20xN9CyNJlJt1R20xSmWb3
XFV7KBnA+ykfl5hIJuVPgDUm4iQ34Kb90xp68dlpuuYQEmYRGNBw63P0DpKUrVUi3/jTvmkxxWfr
C0DuB0SgmcdQCeWQBsokVBkTkF3HPnbuAU7/ddn5d8RuE6OZjE1OQCJlQh7HgWqWw/i95NrG5dUK
WyoKKDoURRG2Be6AxOa2/T4ClWLsuzbaixZlY7S7ikyxHpxHnD3eTFGNgWSES6Evr2mpL3iBm3RZ
EslO8xQKfxAAPp4uO4x0+tf+Lg1U9xVpfRtmQpNFQZrFJKO7OvQY8SDD4rq18HVPqHb+Q54DZ00N
nTTvPRj3KlVWb9vj2Q7QxmcMie/ENpIV+uSNjgt6GK90/SSoczos8x2qGeUmpZAZJ8i+jAfPeIsk
so3/S4WdnFibsKSTA+nVDgKZ4dB1CzGPgHtYe9oucbPry1VDeaJkI1UUaji0UYWWDFBRPekw9dPr
55PTlgJ9ef4afBaosbqcSYtoLTiA6pfG80mQlGnOEztFTOM5uJLXiYDYUAoARGddlm4Bxba23//j
NvW5szE2JpeVaKRqO5+LhUZG0zqTfzcjVpeKlL54DMA4LApTHSlfcpC4oWGt5dGPxcFRSOd1lUZO
1VDZ6siJcCoItS8wSGLrQv1Lr17exgMpp53gjUjd372kPMcdzgpJy/ymL0INnDoH3FsCqzu9AoJk
ZddUdki0j3vbukRSpfoLfeEcsIVRSQBPkj3mMMRoLW5XjbJnsVlLHSBk77bsnvk5vKnk5ytk3oQB
qy1vEZgHo+ExwAZkEbB0R5HNDyVvQ/nheiMdV3PYEQ2ZkoWs9r6sbLy/iyJAEet6NQyIn3td2vsn
TRtO/bx4LlpefjQvFgcu7N8LWwDzOx9TgO5XSGGVdBlBtVBAIGPJvdDidVmELS5lSLujopdjbJ0a
4EUjTCT3Z4nRhmM8y4aKS9J4vsJGmYhGwq036Cu89y8rlPBOERt/ByPtSzo4Ghd8e6CgwfvUVLMm
NiDsRNZDOjd2hw2a3E3KlbPwDlO4s9N7/EVCTY8q/w3LRb2DWEjzMn1ami3iaej1oPZXuuVAPLxN
s0xMpRiTFZvfruXrAhSWpe/NfvYDqBRvGNk7KPIpfFsEjtx6UeUweJkk8ZeDrTiwne0rtamyzirW
oaqZ7RKcLx2jlHgYhxy/OSnF+mVTwbN0+J76Qi1pbbb86xXbjgQjmYnsfbH9E/3jSqo2m53+fuSa
Rxm+zndwzcIXGe+b7VORXyriUzceXJxDHKN7+nna9jkIA/s1F04N/SwE865woX3g/EIFYckXik2k
uNi8JTQHzsKvE6HG5vyF4OVQC7UbsqGe0kJTrOld5005F5UMWkgdfNgZ3NbvN1TrOTXhHh6UYZkR
6X0865WR54IQgBQxnKVicM/aFG5QKvyH4X4/L36cKK3pmmAGF4bEdNfL3gKuSIvJ3Iug2JxyK3L2
ml/AJb/xZOaaJp5JpladsnwdMJ2KeDqRRbIClGDHnrcF/SAbKx1uBMB6JKS+RdWDTRFMDTAQOa2l
fQ6XyEJUZPeFDhjEULmZCNJjAz+Fm3elYdfvMU24gybsrofq74GSlXF+BDLpjsn/993EdTYa2uiQ
yqcFZMIdQtjLpl0A6YU6yBlrLY6UwRToKEWUJbztRGKnTDk5hPzBaR42KkrA6YnqNBtmHWq0I8ou
o4zhfjYNaaQBONp3r9w/ZJTeRy6r5folK9YdW2k/VlNLJf+S+2OV6Hkrk/04qgVNC5LqF4ONCT/E
15oDfTZCXCEsMG3f9Eero+9mQOL2Nh6UniQw7N+SVXDWFHoJLO15lBYygin3GXCYWA06ID1+vywl
e+ZauhhgNaMMLFRXpVZVfnVXTJiU82kaB7laYg5J8oo2Ek0ShD6eFBxHDOoSyJpymp2mYPM0J8pq
vcOiJU9z317Rsn1GVPkbwOPWwSOR3GGbfu5GdLcQjfUXzhAZNIg9GYKZFe09E9hpOYJoIWWr38Em
S2fz028YG0ZSEcpJnAs37HrQB5vdB4WCKCP3QScQmDV4NrFWY/ASYjbT8WfdewqQZKdytt/eLu8g
VCqitw9UHcCoHgVho/Jq/TQ5G8ISjD8AlRMMfdWkvHyKd4BkbFjgv/OYrvjpv3b7oBQsHNjaBmPn
4ecL++lQoqzwji3eqPLPu1xRkF1mhUh76I5FwV94+zSVdLnDOCgv1WeKKcEFBkopEmtHGG5y8zMd
Oks5CSBOiYEOiR551h5YMY6kTL/mbIHTGqVpNBYQocGcQuZDijqWTROputwMLd8/sRAf0E79gTvY
GJ5Z6TRmZyT9KBydw6Ei4z+Rzu+gqgrWjJq35z9lyplKMZipd7fce55gMR2S5B7NTdTphdrITsl9
+E1zlLD3BtZARd2HF5+k50JGOX2k/wKg/r5H2lccrBc238syHj+mEL16S5nBwEyEgLrTVvHMwySC
+R1hsHjN06Tryiyrq3E12o3Ogt9UglCeYXRVcAbnr/b6VLx7Kdx0fDa/O4qYD+KF53DrGIwP8iiG
aLERTHf8cDY4vfseQkm5NnuYs8uYu4o1fssLBlWmqFRPq98btr66kjXktVGFml+g3ceAF302PYPM
3NeYR8aIyYLNf+NFL1WKfYqAtoLAeaDEMqYJvhTRy+aImanHoMd8QIEnGPIQio76/WBqfYvpesCV
U/woaDlmqpBo7tWFvcrU5hC8KRBMsCrwHeU+pjT+v5bUSMEqtIrVgTEikYntlR2U52s1LhcknheA
CRjOQ28WEMaoVvz3WCZ+SUsUZwBRLt1kKzsnEmRgcq6SIMPvnZjgWpzL2h1CKYXMGwvN9VYWT6un
vbfI9I5zkz5abV9TwXcdVphL7Y8rF+gD6AVbaDsFUy5ozkqI3RVASgbEdg0nCCNVcqiFfT3UJXzg
aIzFOo7+jthasd5z881OvUIwG/EQx3L3p83Rine2gg43aRaysp/zLWn66HkUAMacjdOSFXDwPH5S
r8ufVGgc9zjeOenOkRU5LpbIxS/oJCIG2JBkKeT/jP1Bz6hiYtaUX/FDsZuszCRtZ2C9yq4hVxj2
ZhXnLV3b15nd20HcYC7rIDcLt6Txkps93ysf+/MBEgbWuimkND85Ij2D8MhgL69n7ihwrYpKuGFV
7cYBd8lKf2XqoRWQxnsQ2fWD0QBHV8+vQTpyH1j1qSGGD94yPODKCju9c0WGBaALHf1lVZzfvsfS
YOBd5UYyb0rcek7kiRLWvO6dbYvESuGaKIDF8A/gn0bsQf3BwXKGuk9imjaOgJtjXL2+xjQjLM/E
qu7YMZ497b98BqgvrPTPfUKNOc9uB1Ls1ykkbQIlBjgCRurhuTNtR750bt6Bo2hbVvtIAcnML7LW
ZU5qP+YKnbpHtncJE7q2SgtwVQBBFCK6OuzehRmSbqumKFkRP2Xiy9LhEN/7Tzk3+GtUOhrfadQx
npkqTKCeZytSTewr6Pd0O/sgBcuoIMVpJ++rxAhCL+aPrrR4UAOqNugwn/a1IYb3U3uiH6MhLbBz
E33jvNvkLoomYFkQlx4NcGnKzip97CMGEP9fZ6OaYb0I+Rxm9aVhz3Q+pJX72Jfz2er3YGYMIeLN
p7Y+3FO4UhpRgqSIUu+xOUZYe9POA6XD3EmHGqC5UpKRdas87kNZZ9PblRUr/Kr/sVrgLmBx7hj4
tpIUzwr/ivvp1JTXfFtGHhy08L9iyjzdmocViqB3p5V6je40dmp6ASyOBmmhP9Bh1ONkGj3hlAb4
dP5W7JSig9+phFMOwU8LQkwqHRaO7fYngton8IoZldWZ4H54xB0lw2uTTATu+9VfqVs7eB5SEkbC
qljRPSxxqQGbU/hrvn2ZP2SGZ1MBUpVcnlsgh9QplVG4QWI+ZfTtxluHxwe2FPV6w+bezA37NCFa
j0lYjYtK2+PIsf/nNJKehIh+MtVif9Agzs3mtVOKY0X0Sfe7X5MqCltyl5FsOq7WW0XbvjqhIJWK
RYwKsild4U1+sBF5Nujk5FdkrpIzkL3rLu50OxtIhEbRw8LAyZi36z6KEzJy/0zhTfd0+B9WIZtp
4lmG7H/If4LBQQcOc72J+4vAv5O/veRKRIoMDUB0rtX/5QcozWGU0wlvz09pbdW21YoXyBbwBS0G
+/DWQj50NtJfUGu+w8sqzwXZ5Y1bNYjswDLyn9HO1y1X19AHF5zlE3H5/DQy5JChSz0kMW79Tz0i
UYDQJwToEq/Mnd3QanYoKMcS8LMpIwqft84sBA14Yqu2A3U19L0IkZ7JC0YZ02XuG2N0DFc18myo
fFAWpcWYRPRRDTHD5eP2sf0q6xbyNmpbq23pI9lkoAq0TcaN03mQLUOGeXyURfgU6eB+RwW3G0/j
9xfrPkF6mQrQgtQlLgRvUC7NJjbjz6M71VGS+aY1FcA3mWVgBa7jNZeAS+pJiB2SALyWvtrbg+5h
7Bij44PXSULM+wsFwj5Px8I6IOLa/Ee/cToB6Lvf7ve/xQXCOQfZ3MsW9KTWPp1KqFHe0fH4jLxA
12k8/DOBPbTQ1J0m++p/5+6ribj+gIQbttPKVPuRj0pMpClcqpbByWy4tXBd7ZPdySZhbx1i++S/
FwFvWJDL/3NizCEclwTecRDKZsxvbzoKalLEnOifhPLb02SNyQQ2Q6TdlcYyBUbn425D2soCf65s
0wwWc5p3o+yNWAZsivqWlSJK4d+j5zV5NDXAbTwdNN6A6xcPqah/mdDnyfLVy7h84IOOaa1dzkmI
okJSYTKHFAov1KXL//l4pzqDNl/l6fsw3hPkpBmBtxx9eyif135jlibElPr/f1ihndnWpa94ke5a
QFP0u62Mvh2JupISBrV9zFG3e6HIiEaajDXYvFBtjVpvg2pFULXUE4WIfrhMwL+11C1XQIwBiCKl
qP5p9oVyzKKvynIX2Qv0dE3jTBMvKS3b5w5zcKAz2vnFhEsZYbnTyIlhav2Hyfdkap7eWxyvGPNN
rNVMYDVlf4sqiEiB+BXfWJ1LZXtIgiL3jSP0XGvJUNBb7/afbZY3aV4e93odwBE5GrADmgxBWR/Y
0AADhBeGU3Lz89cJbM/eHRz9fcLZprSD0MA9FLgNTmfr+PMmhC36WDntaoIdQGB5d3fF3gtFtLP7
ItNBtBiX0oQkhKsQfPr57KikGe8xOPijnopiMau4ds50lueomDCr6Ia//JzW9zaFP3rWkK+R0uTn
VfwW9XOisPTHNdg3bfBw+RoZbDbvkTee6dyQEgDUQWi6/j7rl9Cnr9lSrtrnbHKk1/eERNcQefjy
rXX8Xjrfzyey+Xiu
`protect end_protected

