

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
pTeL3lbzyXpg3zBlG8xXBsi5mPcSaOx7zOxONTRBSW321/dGdDH2TpaC43BqFdYZqpUNj4ng67vZ
qArBG995Sg==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
I0+MKhxg9FScVNavGFQn2xkzaE4/JyCe16C1b5v3ObJwo9nXDzI72pLgwgIfWMASSmFXtaAAw0ml
3uLnAPMYr1dgB/uJGeAtmT326qa5BMsAV4vQ1Yunxch6eAaFBVMMeEWawv99YiJK9jkH7yDAOpb6
smI54SxBdohXuGVE7bs=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
bDMpPv/P03hJ26zOMeRntjG40FHNolyY3dG2sIAWSb+A/C9vMJYUZduiM8NsMGgn92oqltQI8itf
kfh0mxfLeub+eu7+DutH/IonvZFuvU5PDOu5gXDe5IZcX7PKYSeWlg23QrTg/K5l+bblhZE0trh8
gSCxX9Y5M/tKkk3Ah7QmsxFm+D2iD3pm82WCrtLPh7JqPCGwGw7ZkIH+rqgZe/fQHahkffxj0VdF
wp7Pe3wFKtUoiMTg7uNHWsoKi6g7a0GVmS4unE3L9HQtqDdu8p186XHZQqxkv2iNX9KutOONjQNy
x1JPQknSlGZ+dd8WmzTlL9rwhQHGdMhFcdrMGQ==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
CqlfcKpSPaBiicqGT47t9PnrRSQ8njMbqaZWYqvnT67KXQ7fxmLQJl9EXGvFoMEq5tU8J3rLbBm4
9pWLf80+KgxXgS9WPEn1zRTKt1wiye9VOUHfewp3QYM+B5lPR0EENtCdssVC8DxPUBy9Aythtbty
2YxNBkGFMjMRSnj+A14=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
jiVIVHHI1er6oSZsM5uji5FpVlbZFUX1C20PfTXKPYBzpAjDWZhROWc8xFgszwvy5guzSmUMWOgw
XoJ7z9N2ElsO0s1NH9ojznzy4rNB66tyJa27TZfjI9UYZ/9rfTzXHnlr6WpUX3IChRrS6x5LI1mY
orERQz81jyLKT8cB3O8KkjO3g1Ks65ZIeY+E+7T5cJHzOHJQcoiTTtwLajrQktJS0RpyUJr3VZHu
CSADq9QNuiNkf73BoFHvperz6rZhWbdV5MnpWKfmllMNlSqFwzZuWbMdZs7ZNbssXYmUZlJVjM52
JpTXdo1N5lXyKjXVvDlv7kCHkBmnfQZM3rMXlw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 17184)
`protect data_block
2POBc4apgKhD+IK3RrfwXU921X81fl8cmSahna84jk5O6qclFHItQBq8gMsNjQ5yUQK8tNhXxVR7
xwPLwIipbbMzOjnRHxLUjJfQl2pD3jzuxQkcsQ2Qte2SZksZnwkwuOBNswYMdG9JwrAkCGgGthAh
TYMb2EtppHgTzjbLTpOG8kVDChEFAUA7l9K9F9D1RiMNqEZTn6DMg8e5C9iRrtCGH/Z40hneGJ5o
qtSh5FBY3TDj59/iG77E7m5/SAk/MVdXZGGGf/a5l037yaPGQvFPpZdkFGfazeZidt+AlXXekWrr
V8jfB55I8XVdJovWOx7amwB/TB1vKSqFs7iOqYRd10WM4eviBEeK5sfzcTxt/oFQNOiiksazz7Lw
VY2eH3WAM0cTZ0kxaLBxgywf36BGZNJoTbvC2WeFEHoVXGTp6wyENwH6WsCYOMAsuKnqFNIIhQjo
jwonM33mTevSKxgmhojgk/uRouCpDFW0CCIWqwem78zYnsR/jxs8o393E+L4ffQaUZI57MwEXrB6
rGkam5iTYQhixbwVEbIcwkecooSLaID6zpCp6xz2xieQvXd1VWrhJ2Fe5Y/0xIqH+xqOsvPfgkem
SKhFLRfjz2afuWyzAxqziN431RsclFwQKfP79syOuF7leI7gEu9TxNLuNQnMlr68lf9oUl+Iinir
FudGAiIVdipARS+etLoTcBep/w6ODOHAFHHZfrkOiXhnaVFy/H804EDZ16g+o+7qT2SZlSrmMVJw
Lgtn3ETNfZZN2BSIZNLuwSyfYg/EZCcL8Djv+k0nCuMYClthLyJ0bZtbSraFZ2tFvnx/hL7m5yXh
n3gE45/QMcPMmN53ehYelUUchGhIZk2KX3uRE9iWpVLfh6GfHC4qXerW4XaFD3exgOFLtY552JE5
rYqifv83p3+DCC1R5nCNHrSEZFZ/e9q92HvDj2P7RKGxqdKWSTjYuxCU3XWbOsNmyCmIngttJ1Cq
pSy3rg3rKeimHnSMmThxKWZp/WW/+d7vJk3uZ94cxfB+SGPPsJyv1+ic8mTXvN5Z10DYzfZGfuKt
1csyKCM4RihB84uL6chC0JNw4G+ArU+fWlZzTVkpK6JVfuJoLG4yFyUrwoLvVSfg7BJc9gY8EVRI
iYOdOjp1L3XeGgVxqnMKfws7U7w95xrAs35AcOhheMBW2UPia9zQtg+HhSY3HuvWVk17okSMslD7
RIQlkZabwpB8C8REM7Bq8BfvuvlIRKykn9WXZ6x1/m5PtdvJ/pW3FEkl7Lv2JG3IagUBlI6c7YYi
Jk1g/O6px4/RPorCeqQNCrrcLgMFrAk73H/smKsRskF7O3RCBSwBzIz+BTyQYvIllRQvMWFbKa5C
NyBJl2CQFg4nBT3rXjmZaUp+9GmSYTSdGy4HHA+p4E8DgAF+cLsaXBozwrtO+ns+caTqDGGi6Z0K
RHAy9sGo5Obk8ULudWaUP6D0RE4gHLXJeNrsYIhqUV7yvLTpJyXQkWpDWg4iEGEaYgASV79aKnuS
q0IjFm9YehB1wCrrEFQbc6YAqpxngItCikUMiBFliEgrZWD52+kWKuPEWDWqDnXXS3QMDZzzhWPB
7WAzX75nucm5gyi2UQ6jPQKlklhOHoWwNoQux9TJ+JbpDax1j2t/9AEMWDwRflOxcttD4CkIUuCF
jwDK0i58jTb5Q9+PoMawSxACRw7OZ0da8v1v1ZSS2io5ZggURTCeETFOCxkNrNLLXPalCX7XxYND
00JR+zAJHLB/lv2EBXwUEQ+CAQfjp5eNUwv4W6LtKnQpxW7UuUun6Ootw3fZJNU8YMLrjFIOCaKC
vpFetTdLsoc2uKzKLR9HDNZ9PNFqzDKtodX4lb8Bugjw/M2OlcB0YcOMCsbQQSbJEoyr92kHIYP3
2Y0QHkYHVoQWzlmwdKYAZT46Pm0vjnAcMyC0uCm9lanisRoesgXfn3TaE6rVsiRsttXjeD/K9xkd
tG4gYh+0lgTAWO2VRTX5pqB66/NX44TjSHSfh0/wT9iMr3NQeczJjKcfZjCwKn8xmfjAiaoxynAV
ZxqZcBUbDz6zlRaMQjNJWCKPbTYBIh6RXBDU4N1YiAVwHC7KxTPdiZVCNdrHLEFPTBmlua+1Bp2y
FcFyLo7b8Y6imKnyFkHfmYCJZIpp+ZiOc2FRCIqY1/vrIoHHjqbUBuLpzvrjQrVQPmXGs3RD5aoi
msX+K7SrMHEzlj+fvkuRM+kDyq0fYDoV3ZS42TSTiFZbXTGipKz7EcWBhqDQiEhV+Vs8rnZ9OAID
Lant85rpvmNIaWelBs9eBLxbscVaX7c/e/w9eDG+D+BD9RCc6bnHzGaBcwqWG4iyrh2buZYc04IC
LL0Pl82UV9MhAEGVTlMdwIl25sussy84ksTq8Frsh+kVDsA5wCz7dU6WHmFccUkd1vX93wo43q9x
fuY7381AiZ/SpOOFJu/iAZu+5RRXVx9HtYQjPe0AUULl5BoZnkAh9DHDtjJdm9n8WEWcu9yHaB6r
AAOF2X+9DuQL/eitI7cdmP0WkNWfOEwRa2EprRDhyWZG6BJ3N49fXw9of+/mRLQAaZCi1cmnt7SY
MB4gxivRJfztAwSCzyLY4FfyOIiW/bywKj3hHs1Iw/8FtcHrAXYi3AjtHblekCphj0stthgmJHzi
P3YGp0xK/1u0D6T9CEesNrER2g0BUqu5IB/1D3DXgm1wg213AIqPgeVOGmqDJnUSjCdtb4GCOaHt
7zhEaouPcG9YMyvfj+WNp+x+vb8/63BrJz0ntEqqgtXfklWit3frQ/wlB4wzkaP7eis9H5IG7PwZ
8KHn/ZOit5aTBnxB0JIio4EsrZPwrygfICI31DBNrU4VbdALhrQaCFSpT2quXKf9Wnhj83rIkMcb
JDNwS3t+wwZTZGLt9kkCA+sFA0/8BWDVZ/8Q2gKrmDeAi+YJdeXypjWPZpCe5QGhs2a/csq0qtvD
9ZXq3WTwolGTFJ433ChNhrKSu5r5K18FWa48/dZzBPpExJ2juXD57GfUJoEMK0fQ0DCd2j2U2zOM
BwF6hs2PkWRJg0rkd7GLYfRQ0Z5li4ylDLOFba2Q5qQ8o+tHFdQgTKl9lVjdvCJZXoRYVnry4cw+
vFNLGVE8co+SDXqc/HUWUMlLqHXi7dhoEE6H8omwY6FlyPixIxaBhO107BkuJFEQUYaiWKaBFsXy
Kn40w2HkjCHBQgtmZ9ZyrQAPTllVLMeeqZrVC2fUp0KAMIvIdz4GpbIPBynimucnFRknKmELj5du
N351BZapAALkNJJivmPz3A2WiOLd3JpJ0EYtMIKj5jjFTqTzDKrV44wYBXgpvBMzQCKSk767+GaZ
4+4hXOv9YJXHJdWNkChqZvGHKO08vsqtsjYp85gdRa45bAn/kEKnIgFgG+Bj/OVIQ+eSOcFCYj8Z
MP77qgn+8U1zfK1KD600ZovJjEYAzfB1gaFpj5E5JUPMNEnPGWXiKj4v82l14OnVI6VaC884qe+d
UrIbatkjYjgZp1fWuPngIe5mva3JcBCw4R7OEWh2uhQ9TncsSKh8cy6PxADzKk40ZJL458bW7BL3
4x1GkdD0YEKeNmxIhVz1IZfRNnyArhS2pHpK2lZ5x/NMQU9j5yOLg7yBSJQiFWuEiSGwrBorUGNP
Jn45MT9WNExHIEjxL35YTQi9GjrpLI4TwnFG/FK7+HQPF8Q3yFOmgu/h7BuSx43mgf9V0ytor07S
l78NEYuSxx/MAzf7WB2tpeUKGRNoN+VDe3UOGRuy4v6hsKpkytMvlLl9ZTARdJjupwsxhFOzVqcy
IHSkL0zKOL/pDHQTcff5dMigBLwqDXoaxR4t9sxemK7IX4xy8JUPi1kcNblevjX1d0LdynIP7KxT
UrEorCC8HAQZ28+6wyXPvGud6vb2YWN/HhXLYM7EZLiVS7TwIcCK00feokCZYuZxubtx0bC0wOgz
ayMJt72VjqZoUVGt+0Hj/96t6vKBVUdzogoi13XCcbd86wcwNAw0DmR1UQ026IDimwNVlidxC2ZZ
NTXoQf63TI3GVlXIYTgU+bo5tZmSp3fIevCg6+04Qf5wELcQbtwao3eyJQGk5MpMET0QkdS7aXNN
cLHj6KsauNeU0ed3gV5GmZrh9nikDWJXBE4mctCmBGzyb0/HgjMGsNSQdqXbBwDyZHftg+GG3g1g
dMmrb9a/pcvlrDxK9dpddMsZaikAkIP3vChinZCeq7i4Ir6JsFpPRWZf9A603PCCcZNLzGQ4LhcC
8AhjHNqyKOJhzePGm4Uqdh+a0DUGEvHOJUB35o2g46vM7c89r/uisOS2EbEEHY6HR2X2InC9qI2H
KKfHcxU2E1TGZcWSKoUCWhUIRyJ9wvnYmOJeVU4dENDzhsEiHyF6RpQvd9UiEyOH7AXL0vpbtAxt
uL2oL6G7VJRdYjEY/CGAtAIz19Nku+MkipiwUT7EidOK+iBOQHDaEqVPdwHEquQjy6BooHscr2TI
jLhYfXPr725IvI+9RTCNgfl7x849iGoeWZxiOcakp8E+pd+gbymkFpAUrwFO4aMJpD+hVL1w9Xfb
lMmNZqJ3oKRqCoczIjEV7dTfN2sOEZiAo2v2Tn6NcKCXElpagA84kXADsR7R4R9Hlhjh5T/vcRAs
fTW5MLHG9L5K+HHw6aldCVbPVsnNKnLzjNp/bVpnnIBqStnIjaLmknr6GEQb+Dtc9HWZIXRid90T
SjGayauHG0CVVb1i1w+JQkuLbzuo+eHqLhiHx7zbZT3e8rBoWqY3OGCRmQJCmRoFcSeyZRbRhpG0
2V12vSmzB7X+kwNtspyRLWmfsVk5gd5ENZiCkvjnjffexz/6eMPBSQ5F6SS1MFDl2CpV3Huy5Fg5
280bLbZGMXMF7tn2Jw0lqGaPICa4fxfrGCfDIQOmH7esWFXxtavoDYgUMh9woRxVs0TlHtnEcrOc
pt9bOEHNZP59UQZCOqkWjjjidr1+kOblt3h0M13T06UYTVXOcgrOOzTy/HqmkmuUl9rOWYId3bUn
yt8DpEAY+fzqbUf2mTSxVkGlDHzBh0oGyaulMJN09o+YBmmsB6uLMKX5cviE82zfe/tu4icrkIoP
cNImpg5mAtFb2WZiq0jqyZ8FJ3iv13QQURkenl2/MEvNUXS0QkHGewNYSfoLHatwks4YMSvrtHky
L1v0LY6XG1/Vq/MhncNj90PUJedxQLw/nK/V2kTz9CwmVmvFTwK86q4TbbdU8BWqWhO8hlsohJCc
NZ1MlV+hrKAXKOgIo0foUHjxdYAzEjM1BPblPDp0iYSywOpcYg7tHPHO4zeekyzFaBRlu6Wd8ByX
Q+kbnMzRvJXYu6KbJRUQlRsDN0WwogtIhF95YYpRye2z85gPJ9khFUwuqbv0OdmX7lmYw/3KJCzF
NW/j63GR/oLn2SRD+FZi4vzPy/7+4NOR6O1xl07RJYAl50nFTOue8ap8/+ft4GN/PP1OnBO2ofSO
0i7qQu+kIA0IL93BRCUCIXXDbi63rfBhoXazGFDioaOlUpNq/zT+adI7e9GJiDJR2KlchoYbK2v2
OvE6NPrlCdU7GrbKLR5EgPWKD2R4DZWUqBp0oOqwcYPZqCyj8cvVHdKLp74t4cqMvr75lliBGEto
qFuF696DVFqpwHEvp5usrjAi/7TKXg0vqIkEG8yDiXd28ggtnXhywWP6wh49i8MsJeFEWr5HbRWl
MvPUKKGIO5BIHAFRtnbUAr+EKBylu2JnWiusbBvbbo80CA3kBryHpc+5AHli5PJUzadbD6QwmMMM
k0yjAgN6feD24GsApmURb2gYT3M3ggiSPJG6x4z+HhW/GjucSh+/LdNmmVxu6Afur3MPYNqLITtP
XEUgsNtWPvX997t47loZ1QRgtS2Zjn9xaqSAnNfLtNMSLKWSHpwin+3zQYbZiM/rPBykpk+Ym4qu
f2tcaVAUd7NtSagpLC8TanMuf76f6+EbLY8Iqg0jGAvQyhwxq3TeM++XUMmIzIG+2uWFC66RFLnb
KMHSaNPtSVFKuSuWU7jqGgnRyfL75jnoN4TSIv2xrVRifCJxDm8n9FQneMPFzDWe+NiA/0KNe++h
6oWQz1Mmh1te3A5ggfgjMAK88vth/caRH+b2D9BlWneuQno8zQfF2XGI+PKshbEMhAvaGqEPh8H4
V6LpOIN7BWGi34U9jQx2AgVtP14UOyoAuPvkKyYoIiLU3W25bcCGoYl4ww21QfBUChYBxcK04A2E
1jf79gNwrzQyIF1Zh43yVBqvsbhYquto9Z36UPwAPUj28/HKKPrk9iDcamAV8Ucmpv4KGJTHUpAw
Y844vWLsr2AJ3+HKs602TNchNBCsBPppXdBtu0+0YjzL8X616WfOjen5QLdmHx0dgh0oqpQhalVw
5h+A6uhlTDR2JbfcvAuHP+BxPTYzGdRnyJ4se07XSaPR2WcYpSm3BW8dJzobLJE/BnqicmHLXHp0
lpaeE6tK+prThKXmTEkPQMZCXETue5hlLNKFCfkzLjubRGtRwcSrRF8gZnL6sCszKLNlwxOpSNAK
gWLXZE8tKwhMuIhCuKx+d4/4kG2QMD2QOlIib1Lzz7s0kN92yPdPSFeexrbO5QlP6uVaKfBbhkRr
JxvSSIAgceKrg8lC8+F+H2gXuyOi4JhyNc0oxs9YrtyXQRygyuqdBOzQMVLcnrNe3EcroEUvEfsb
4fpU1LdzZiuVkxmtONI8M3ula/lItCOcqp0SbHtD2bSChs4qpq2DAAVcMmCVwRga+66QADy7fQqk
Ec2sUqfHqam1B70RkMWITuI0TORqTq2sSl9+qc5TRX4k2JWabkbHerWIh8Bv8llZgJ+v2B7LuBJW
MBfqGeFzQ4IldulS4K0hwQs10fZmHyS51IRD8WlSZ/DtpjVlTCvtP/as0hoVRU7Z6mU/lK8LPKlS
+UDH84fvV8/UvMCL6ZWKrqQUM8zstAhEOToMuRj01J8iWYg3VEcdnDh+zv5r8HDnkRic8JXPejSl
zXXcbo/Z4wkazbInIrdrE8TRigLyBMaDRYZGrqBeT74FziK/X8N76es10X7pmoOuZEvKH1ts1n2i
YiMTj5bWAucpwLbYP/zcy6gz6qon4OHwl8PbOry6pe4qq/34tqknrBC15qm8X8TMurwRmQ9xMvTJ
1sMlJ9lVs2rX8FokjrNLkiJrM/08wTl/Jx/BeKBkGYete1Hcp4ryyB2yEqti//IUIe4emwCnT/lY
3UBv3pPGA0bzClJBLWk/GdyirV9UJfJxzVPVbxvOCfWYSKe+TF4KiaKU8bBjaLta4k8361/Mge16
FC+oCv23HvcK1dIE4Bq6iVfORZXss2OYSgB3nFi4r0SqmsIjjxTerD948jMRszVM9BTIsSL229Iv
Mc65fatf2wqJ5Vbi+VElQXxydrXb8ioA4kExPA0Kok7C2GhkQvhzesgPSkpn9S6gzRUmrItqtZBT
FWp56813XFeNx61TD+clAlKbJaajsNbo7WUiBxFtvs2I1zaEzdxQCy2NjPsaXqWFvjnvUGyeCuTZ
prSZUrojtmgfcqxrFdp/PgV8HBaNV+ufAtuwyxTG0vZdoqv+4t9iFisKj3sVLPMvU1+H71gzCFYU
IW0XklmfoyWArq3UXZxYMxszHRwMHGqq7n382M6cf6h1QqOddWTnEt3TXzpoQXglyYgrTabaUsDn
03+BK0Rq/j1sgnqKQlLPQNbmvt9r8+/r+dqn0WAPHQlYFHzkRYPk0ugmDec6fPCIOl7WhFRC6CQL
jLIYTJeyeQRwtpCeXr4XTNXqo0hMs7nANhwNnWhjQON/4/DtPWlpqJT+Pu/vOB/BeylMD/qKSL8t
6gXGutmIdH7DB9Z4McQcTrItGDS1zGEpiAQNNawjS7GZrnWuvjRI3lAtg46IGFVsBn3Ad1knOHq/
EwKJZmO8PMEtQTjX3UhC5KGmAxvZeR2NomPCD0vMPK6r9tAztxivC4IHfxVdEaw9Mm9BDsHAixUe
t2iJIkh9MqNKKNp54gGJtaP4aOQr7vQFh6M4tKky7u8gL8Tvnh3RnmCIhEqIc6/0eYC+x30oBNky
b2REubj39KQHR9k7BVv4yFCOlh9Aw/LYwtSgEA+Bbe0JsPr/jC6agsHFuQLmvneP5Jg5W8S/pITp
3QORO2ilDGvKI3SqPbZGNEP1SuvxKrKFVXe6OtDXflpVnS7ZPdRLCcdbHGUzkX1x/BHqBXQGmEVf
wdukCoUmwhmKC9ocQ9uF4Uf8V9Mh9352aP9MSrEzZD3JQGPHy0G7MmE3Dmr6savvL+YSrUYbdphG
9hqCo1LotfS7lUL0vfKlS5cvk8pMAMVR7UzCxjsCd3YXEIFOklwH9A+lXx+gbqUBt73H5C15TIXl
CPwtYSRRazme/vyuWwWXdMTvlgYNVEMZaV6FWo0Hecetv+aumN5V5EpSXDSFh3NeIjdHII4GzgEL
L1IEWjgW9uzDOZIsuoEc2jIZ9NLZH8NBPJ2YeQWAXXdDRpQUQEMD5ikay+BeXWyqs53z8qu0GYv9
17lKq8txbyYiBtl2dwroxdJYu1yhbLrg7Bmz+rwbzMlFGpZD1VONP1LW5gZXtGX8yyC44GzoMtVF
NtiDilO4dCG7UGRB8hBCoqUNLxiTHRRiJ8WJISkyoqTHgxKmIBtoFIN8MDamAWbwau8gkFnVjx5z
jCfHUlPG06onzA3dJ2u0RDdeaqX2qlHzcgYf7rfHjkOUpS+vEryZmAlMKhD+TuCXwPTGOWsoSMgW
j1meOeNxBlZF/YcKZ2CUTuQ8bqwatQER/0OJAi8b/vWxU7IlEOvCStyIBXriNOHDrfxQJW/FSe/D
y9hay7AhDQDgZjISjZTzaJ36qGSHMusTHvZDc7akpBGXAZoQWfZMpEMiDDBv529iV7ykdZfTUToN
2w+2Xn5mUV0cba6829gnmJGHnv2eI2/t4FU/bKB68+AfTuypJn+KYj7NahLRUT+AXckCsEBU8ZvC
4ve+U6ulrcmNO89lPtCVf81MV4HPFKJ5QSMw8q7zl7/HQtxX4k1PplPVnxH0RfDW3/klDgpZWkWd
1HB5nRfgPVCa/f2lsqTUPlCWFoDE7izwjmEk/zU3M9z8/B9k6EOXR8V8GFVlk4tsmyNyaJ0LWwFf
DGwU6pisyhFsey8NjgkIdwVVupwaWQ1MtMqzgklUrV7bADhAOdnyN8ZpByLpmITSJ5REdCaMZ8MQ
wtEdeOVwVDVOoNu3VciQcySfqgZYg48hd+b6rdxxGtYXDDJhw5PLlNxL/AxwTK7prVMcw1UBMA6S
yQd5qvfvojIfhOIpI1BdTLIiu/yNc4fAa/m5KD32qBMggQ1zVkODpYYtDCG8BlF1PByw6nRFIQAW
bseQmm/dA4mHlwhYPPsyuV5O3BP/x1BlvroSewfq0clLEamqFF0x2BOSvTv6BYkm12uLHYTS54J3
iGdxK1YxOTbzM12wuZ0YrWrV9Xr3vvVUmwQj85JzSc06FGN18EBPM4if4wNGNrQaLRO9HDhPHgcP
2zOSEshTPxzwM8xPw2pp39MjQfD9KB6kTi6ok46EADbVx1Klnj2Xf+5ib7K64sNIfBmq7WiIBWFJ
Gx7zP5Mw7icnTEJaTL90ej9F09Cjgy6BeFq/mBssI5QTh3EHr04OWVDzI2n+N6r32A1nxx9TfFzs
3sFOgrTUSs8E2PVLu+LnFsPKONJHo4zF3HsKosKgApHL6BN0W13Vh++C1oYTT0ht2jsyKjgsscij
cDR2A/T3BJA+Y6kqhifhIxkhS0h0DvzUcbEVmL4KVXwgE5rRHHWFQWrwuLTv3Ypb9cJoVGqALAxe
2EYSusKBHPO5c8ut0wQnXkvC37tTlmKgULEklSMvXxPW7HGdCDIdTRbDrgg6lk08tCmtDoOKxmtS
4rcnINlIIODHJCP3wHoE7fSgRSVwZ4g++EsrlS3iX0VhCjaAwjHX93kwK5NwY/qvdurv2oFmXxQQ
TCtTtpX0Nil6TparVHFsVBfVESm22JBcYS3Hw8AFG3EP+1Eobx6zb6C7C0syF7l0XfGo/DBvo9xa
h/wrOOTfgqPdVioOBhRIVyQ+8Yx5JGcvSI+EE7te66yXiGmaLBV8erguZKXOX5JEqCsboREy+44w
aTLwpshLZC9kyc0k05nx2vWBv6SszD0mtm+iLT1zSPXLL3JJluekP9S+g8uPxafFxtydqE+2Liye
EhFKRxxSjhPm9i8trV/+W1e+QZf67VZ45GW2ro0cZP2EuABpkDAyhj310DdJ1ErPK2mThbYaSLIo
lo2JkMole2igE6BmtbU36dDoyPBNl2dSvLU5Wt1JjyUwpEMlhmvxoC2acH/+ELLvhIwtGsHQTdbn
C5lMB8Lzhe12EOTw8OQkifJPGCYzqNza68SlMVoXI2oloDyaZUZPVFngokGWJFakUmfZWv7ir4Ji
Lik6pK8e6cf38IhnuBZHsCMbxcG0/aDCVDb9+ZsIVqk2/auved3LVaqpQKlN7cmU44wCxsa/Iqjx
dI7V6TWPR6OVh6igtCW47lZvCCliX4pRPEJST6QsFqqRZg0mTjnUQubnZnU92oX2OWmOhDIewKfe
OpOkbZS53OTSzOqhsnMZ3CAxDKOHBezpZtCQLGjUG34f9fsJD8379liLknp19s/a8f4YDanHW6I5
zSAudqjKRiMDUQtCm2lGqL8vWZsd7fEvTJuHxggNpfvX9E7Bhg8fLlwr2ILkuwdymy3zUyZgJ1xi
N2k/dNY3p1Qf5xHm9UKkbbk6OPU2VjvyZxqJkJozYEgZ+Fk4oi99Mt/KcUmdOd+3A7wD3k7IWFSn
moZhNfg0dL79KrbTuUzOKNyJN2nvIZHvdsjvCM2GpcHJa1dnsd/W99s2084VgpsAlpOo6EbkHxlk
9Ug2FdC/Hy24CkT0PDoODqzQATx+rSgeUY/Jqs6/ipZatFrGfUuvHbWcWMEVLAZIQQFXmj03JboT
Yf8GYcJNYvVsowzw0Z/xwu8SFwehBqo51fhWnZIvEZv3UYQA63Fw1ROykcHLDOcpf/FGqDK6h7WF
p9NnglWb8x9cSoJOvPnSyJYHD3R5YKsrANb3LsghH4KIQ2Xj0r/e1/woA7LFCK6BZ8/wXToXg2db
kUCXoiisBIH1NFEiowW0DFvoe1oF/LBMYE7rkI9j45JbYqzMrgvyKyiCha+dVVVdLKf/dyo+JN0Z
YcF71oYCbRXS+Pa5Tbi9wTypHupmNNrfAidZmIPWp8ifn+bLFmlFVnlK+PDueib9Bb3JXq5mGNdp
cU1DbtK1dQofBUlgF/Ku1i7Oi2cKweRfIRHu7w0vBChTysPDkzJIR/i2UznaeyAiePVmyGIHZFMo
JHWy5GuYpovAUGJXZ3BoCbpeuztdw5OVZVZLgp//4M2NsSzuE3PS9V2hx0aSsTrrUF4HsmfCTN9d
adGlsV7oaTNrH584ytuUckOuBH/hgOiOs8I0EwscIaSXTE098oD2CdfxVdW9TYVEVv5NeEehbX7Y
UCvPN4u2U2Wh6s+1KJv9yvspzeIj5dZhoPC2cpJWtsYugwgjMOs8TMRagmshfRSpMZLr7aRS72di
dRehLGUDQPcXdtNOkImZNi5g1s/vce/zA9znOsGQml36b7CHwKXKQW3Gnv8H1rapXUyfvLnKKlf9
mRBcijFEimo+A8NGtdkd4XTMukSKS3nU85BQXhW6E4OnLGumYtHqNcK4o9YQudVOlf+/7YhSZ1Kj
DvgcSIdigL0veBABXRLr8nnBBdfz76A5z5VKqg1gE8JpQsVQBrEZ+Lslvjz5OG2jzQKlsKC+Rvnn
q0/PrWaO1kbPA6GpSthBNjH3mr5D+CHJj2RU7zLqZH2afpN5bmKlgSDhE3HHQRu5R0dMIBcWxSpR
qUgPRSokcp8lYLxplZuTlmgD89E1/jzZocLWCkzlGwKHhTur5/RomfF2RlFmR8kDmbySG8lnMmvb
EUMs2bU84lCMA7cfHnC4hTTghd+5sZ//ezs/TZLbu3tjE9QfeqUoISFiDYLANfIUnvnkNYhmvqe5
GooSQqZlrG97l7wBPiCbiEg5biHEnQWpeb7wVXQITG4lA9EnjHbuBdz1kbi+c1T6MmRkUs+EGLBW
syISlrzkuvj+fPu17rVaMKhx8dPdnctjuWe7nkQlMjh8VHjyDPSJ2F0FAaA7CATM4GoxjI5Dg179
kEcW1cYGvNYQSM53SyDBQro8fOgd+HHaJWjsYiGJe4I2JZaEks8EXlRNvJOhFpeJ8Rg90f1678Qf
3Cj9MsNS1ZEfICCurOQY73arlUhrqRTyO5JrbODtXuEx14b9QtKFQ/Xsng36zRbB/uAxoVDFEP1E
xRYqdUaOMTNIoItnIfCkL7axWqekD7Y2azejQUFqpvtor50Evlk8Qik20XjUn2h/S/Be5f8Krz/d
TSu6Y2zN6adkF3J+pbSKLaMCBJTcm5RE5K5EBAnpKEfATjwA58KVZ3nJSVvidmA68FpzieEJyBPV
OmOTPwwfCP3NLtl5YQDNh4ac3+MShrTt6l2bg2vAPfQTWiuxwNpf71o9qS3T2TevGOvvHKIrUWQK
PG2C3TEbRznjPgzNn5ZGs7ma/zlQmorz86vi3x2H7EHIv38mtuEVo/8ptsfInQD5qyF1DOgZbGmP
m7UH0yafkF9CvJmjUTJ/L16wCqeBJZY5O66dZz2BzFAoxZeJ/rnZFien9iGPbfeiVac9/fkvrfyh
PPaKlpOMDElRWfU/52kzqqfkeV0rbH+m6IKjq2iqr8ZBxu5ezzxadxnGnSvqFF5c/dlj640ICXHV
hIv06xJ/w7Ut0gukSriH1FpEmeIBDPh4xkRryYdyNMgPpXeGLiMbSMqXVUANWfOoaJwmZ71+NEQb
L0J/5RH+Wb+89MQlDbumrxImJRHKSuqm7ZLLWxK6/fZkMztYrp0Vvi+cl/E11PyFGogsEBWFfjb+
gViv6a4SXtTLJrD6S/dH88LGsS2yHwD8mt4+PcPP49EdaGiNsDxy6rKdrf9QtpauFxjMzTWPzYx0
Qv1tLLBDP5GcW3YMpjrGvwTKWZIRpwMMlxhN8DE+43U8a3C6SYSHPv6Oz9aEooN/sHA62OaiezVn
oLHAN+uRPJtJqgihB8OPDdSx04UersyFHjGlzEZEOU0PhegoOIotm3wUvJklKGCjXDbhvaiZF422
yHe9npYwcKQOYd7jGMdU/jPj68+47qk7uQecSmDN/6jtyy4EE7aEJJqzzoIFaxFQMx7sbHCwOcRf
I1CC6sj4ulnkfL4K94FLrU1493TJTM6WHgfSbwCYbz/PLLSSm23uFHAhqW406Q7XZ9dn/6F0QTRB
3Aw9u22pQxZj/1S1o+urDXa6pCZwXRaK+iwEqeDkDwJrh5rQWLSGYGq4ehOBiygClv5v7bW7GbwL
Ff5wUdIGyIz8M7oQ2tK+vzVRIFTBImo3akbJbGWkwdTMXRNjdyej/r/DeCmtMt+6x28+SZvAetKb
tM5eTQti0XHVSwV/RTJQm6RDoCNkPu3L3unPt/LXdbPBWZpCe7neJ3xmxzyJFeI7QfkiGisPYF2k
938j2jYeGBhYNaeDBWeFzqhwkReFNVx2q1HSIj2jt422ahWm/A8il9w6v3I+l4+WkqE5tO+jgTr1
EM3z/L/YuJu8BDdxlTTLVWgWq4JfBSBr42D/WkHRb/J9oVONx0QY0RJrCxbL+2j0PjX0yyAIdG28
TdtScqwf/l5u5ASRxyh4AIlwsPkEWsXOsB5WodhTpCcRqWk0rB0J5jAYWcseG7d8eB8CB1VAJhgl
WQtJkLioWmRaH3028Zhg3jgwervMJBwFroV9tSwTV55/lc9/likkwc1eG3i4xWkN0IRpwT5Cx5sZ
RDJIfyavt8CaIb8n0QIywwtP90gPnJSI2rE5tLlTbyivPPs1eTpjKkdP1To4aL2/L3ktH6jrrEDy
GHt1dZ2Byb5/MWcHuOG+j+I1PAkQX6W2JjCMMnI6S9LU2wf6Q3K0aO/RECz9p227Dny63fg9K3uQ
EgS8lmIokOzX0pujP3RyrEb+ZdfqhMSkzo7Yd3i0yL4Q/WYIq948m09nShcw/788XcsoO6v/0Phu
AGoTTl9FGdx3mT2D7YL/ztCxaeWo8eQipg0Cl2/Hak73lu1ANaLnauhSqtEFOBgDFK14PSA1E5iC
pbvtuwqAQK4VlK31TC+OAbe7Jgr9y36Qjuj0pMcnYSi1yQ6iPc8sy+m95ZHMw9drhwGSzCoz50fV
PWh8uA+xkcn1RwTEDRXmFUrc8gsxiNDQERELOtNpUxKl1C8/DCcy9oLcBVsuYcc7cnO+eYstcYkZ
fu7aY4oGrdKX2jWeIl3qem5Nb652Tb6MbkPqv25F5yf55q/gQ9FzRcNV1EBZ1Rzo+PaQquR6di3x
QjZcD32F2FZ3tKyH3unbKQI5ajEmzeMgU03bZz9VuQohqJImnfaCOG8UACerTGg9N+aqT0UiZPRF
dIZKypL4GKKoMjQ4aCPAEhwF3N41g0d0MbAW/iBxk0vmvGzaeVP6tPxaIU+mpI1uQJgIYAlXxY3H
GD0YJgOvzGQlnyoaQijZgJjXxhyj+Qzks+01Ffla/gsnUgBVbW5zBqMh5ngoZ17u7JWRz6opjxH9
6bCHUw/hgdPevAl0VIue4HHOZBiGgj/7dQ37cW38mbkFfyDSko7tYwWHM4k4EQScU4C+Hi/emZvl
/9IZBStA+0inxqE5XqGEL59dtfWqB/AWujGdhFTcqVOWGbSn/0mcOo90I+jqOEGg2y70FaQwqku1
k3olkUICQgo85VT9KyKNI/pTRlRBKFxoVxoibGsrXqYI5jSxDpBdtQyeT4rQg1aDDW2FGwQ/ZL21
Ihkwn/LoJslg5gw/+eD6peWPzYzw7UGQ4Q/4Vf7jUrDG2ygQ5NMA1rKjjrEJpf+cf1OOvYVRAOhd
DWxMNtXwfM7aaXwzhBAJtFMditxepHZYOSHxobBq9FHMl4aR9D/aHm9WBs2puFAcNGmVyb55/f7h
FWYyV26XCqju94Lbdoq86ptHZd7klHsQ+YJLmZfCuIa8fYobviMe/ytmQBpeOS6ZwnEgYhPyPJ5+
Au8a/KTazWQK120r5TlAA3Oxc2RAgTyloWUPKzKFz4ZqtDZ6CLtwKWb/p9j8CqH0wF4lGEbO7Ot1
zxuHiLF9WiroOC37PzVLv8XLOYl+x9EJF6HERj6yEYs1N0j3lb0tEJpwa3EpJEudWMUNCcS7+tZB
88iiUIw5Up3jJR7wfD8rPlWNJaIJIP25au+MnijJyeSYVlNatk9sSYKJmTFJ1kfWnvAK7zDuSY5a
AcumuNRkm6m89NGL8/o7/zKkm04xETwt3CfmRTqmTCKQZRuhJOkGNHgGaji7BIe+YY4ybwRi5WDq
KeIS2aDsN7w7YfkyfzenqqAFC10IGdhPXAhr3wBvyvmlWKnmIbDW0fVlfs+uTa7XXVegAMbh0WUm
F34VTUPdIapWdroMNTRxO36K4wQDq7qHTQ2TdcGySVzR2d1yDFsPoeeJs8IEfsfedjr/okH0xsFu
/A86yBRYfGEmS8YcBETOIV3O5Zu+bJ3iFFFfQlcshZjMDOMiTkbm+LxR++Hivu7RfQJq8WwOmnUM
TlBV3oGsFZXgFZRuFcdYm/4eTDKeuPbgetwj7Ahbs+AMRyylDZqNBSk0bffHLano1ynFu9H+Ehzh
MH09M0VituYy0qv3yabgFKwJJYCDCcX74A0t6DhOZjMqDned5IldwLlJyra2NMC065lZqnRPoK49
03E5FuSY1XePyYBwDsGQR7Q28PkipK2Z8omfyzVQ3UUZUnpZxkQRAgkJHgmli0Ik6FJKiO2JrzOo
19PQHO4t9IY+3OE7pHIEkQf9vrcHWyj2oWgNF75eORtmK14RunNkahHZYgkRiKZr7vF2yslGDEUg
HAGmynVUmtLEhMxw2o5TyamFZaTTVqvxn7bmsD0lOPZVnz75enUo8IJaljGFB8R6RXBFcLVfceI8
WKrX/rzoGdSyRcNIoEVt4UuviNOP54agMZlIJQm7rtlO4Q5kVHD7i344AjtsY4810X/B4qjZuRKf
7QZxUt9VxvFp/X+oyXewW//gDSz6G7Bz6094N7F87JT+LPsWWD3PtOLAVsi9oftaRvgrSJbdNQw4
hZ2hpDm16pvgvEMRVCCN0/sg9+WF2EFW1FHte9G+PCNeUh7ZMCGRhHf4kQRBe5nUm/gEbZF/W8M/
1eXt114sIwRlnItB+JDsbMpERqzDW9rXvOdqR3G9i1iveKIdD4YFMxlaoNgw3uL6dond4Bb7MTe2
Uy/La0LjYuccMlcwWYWskNrE0CcRqWYWDZnff8+FjcnQ+gI8tDlXJhXTMbAEgOjSnJEwcz2udHF1
FBFB3t/G/NLyjiLuD8XxQ54u+mII059f2AN4j3PIsjY2l+w0n3RqmEFS86guumXrBdsv+WkaSNg/
IsWskcf5xfD/mPEljjMzjF/MespSLPwckGXadqnDcP8J4KXXChaUUeL/TuGaWpcQ1HO/DhdY8Vpx
9/xPiQGPoAAw3My1twNRxaFh3r8Qz9qMKfP12E2qvBVlsx9g0XzVoJDQKqnS0Jj0Tpt1gFacaxvA
q5BxppvYx4ywB0tFKc6peDbELIp1e45lb/ZndjACDMxnJqQ0HPbY6EnfDI9+o96RC5wh8aiWFvEP
0hQ4LDlFZTfolimIl8IiOXEKWDArOBf+bkXeSO5StibWx0e4e6wfp4z1SlhLdsLEje85/bnyGsN/
TXeS1FIHnU+excbdoqPb/46yb1rsnn8UfgK/cogn5SF9j+URqr1fct332NVEDSisZc9c2Inrzbb8
dxGekxk9lfbrN4nmk9AHuE39vph4sPgZFVgzq2QxpCY6F12PaCxHZVANF9YXo3aC2T1Ult4O4Ee4
NIF4wusS1Z8nS1mLLI28pHd77r5SlsY7959MxwJSBn/YzdbQNjlWNa1y14nRCXquixSm4vIA/lDI
lcoyyVZXcz6VS7VOTon11x6X6Uo5KIYGO844EbEFB3IlLbsXgkOKhGEVOCD3tr/NszLV9NbLVVI6
D4U81IL83m3t5bmPnkyemyH0SJDT5v4Lol+5PSGYSf1YqPvHqnNtNPwNNqAEISJzhG4cV1t+1U6L
NjFzi/KCg2XjhIfioy1lVTahULaBVqPQvTmCw3zRyevJokIiwsOX+ivBBEO5J1cDgpSih7UrDvXQ
h5Ru5kq8Tvwdo3fWRmH1wcRbUMET1d6H7u5gPp0gpul1Hw+dKOwETG9GTHPWQn8KGDn75X0iaBT7
hsjRMqjpsOSMAwzQqop6yOIIBA0LEcI04geQ2y0gvIzT7Wxb/TQaKZHU71C16UncfEITDK4YioiZ
AnhnliUhc4/pi/PRcMBGrqFJmyoPN1W8CzQ5B50u4IfhJfLnoUy1Civ7pcJ1R8uhAELrYo0cS+ag
FrxkSx0hliC2rjTRWYat1YWqycp9YK+ekX/aGLu4+6tX9GwnypEAqqw0srO3VsgyxrHsf9AWjkwN
WCDkiZyuPWfzuv/utqLWR6nSidwUXxm6CbDCrFYHI/93QPsWmOB9vcty2SWOu1Y/BX47e79T8azZ
WOfvLQei+qNbRyBfmQmkDDps7v5u/1GjgNQr700xaIOjAudk1xx8heD0V3L8qsaPlBrSnjITl7h1
vB6K7SYJP1Uhu8YodoMOXDsPKVllw/IjYOgpIN3Detqtowpl/FlSHF3OVgTAxIXxfhyvLSg2AES6
04CXmmuVHmwJh98FGI+zqh6s4Em95Mf2B3z7Obz0hjtd2FMbZFUjndZMfsgw7vcx4NytZreDa/5r
RWZQub8PvxP5169dSyPM6o+Y1OfpaafNLwkGRVw0Lmgrt6zHXaYi5zYyX4Mc+tZ/tqNa5S4za2Yf
4yIlxu9Z3lDYyfOSe5mkHYoVMc+qqj45w6yAfIYVVTqinPjXmx93Z5uXkVuukfIQ8FxWnpZrZu1T
9hX6HEjcpcwC2oE8QtlBW/V5k03BDUfK/Jn33us1DN6ISe9Bfcy/88WHS9wXKlucN1aiRH/I1Qy3
co1YIqpKVXN7hG7C/PY3/17rM8TThwQ29fFToGEITnGSc1J6O+pXMWYkAN1LQIDm2mnR841zRzzL
QPqeOdrUK55svG+wpTNZxErPH3tPeYQMJgqAPbYOMssgpcDY+X1/2BN1btqxtUzP4hU/Gg8bkfek
F9sxwBAW7qIW0LN1m5RWsv+Ov7tigcMLoGNYKFxHVvcpubbl4DNaqY4JoHun+IiJ1KHNaINA6z4F
a1YJJNgPWi0nw5il+Q236LPS2OnSiGunVYN2Wl5Qn0d8YtZAPFeEcxDagu3FI9EoUGZP8CKKf/Lw
ZWoBGqo2qquHk9CJfApI5XS3+/DSCoCJb/4vUCCdD0uwhVE9WQQZOKnezBlXHrMKwCv79E+8cDMs
XTVCwwmjIMzKQnRnQtGncqlqrFPVJ0VFHxSyqqKJtS4hUH/7VHhkV7PMxLwbQc5sJhnjXSE/ccRk
XX5uOhkPPM9z68aB2A+ztZ7xnErz1YRqnZBj7byTYItLy4hfkX4ml3mJ7NcS/CEZOhhvJ90SU7TF
MrHcFlKzxFFbJuqyhAGv0AIUpE5zgZFWsx/+SsYhfZlT6s0G26xT+x8CgAp6ZjHsbydexK75/IA2
L6k7rNA+8/YGmtKpSqTzrKuDxn9lZPDPfJCE3r8g9E9605JBLdhn5iDeYmQaWLZ8EMsiMOmmPZ0+
9YWxpnWI3vtO49UtzBTfrmx8qtPjLuQs/pwqb4PK8GRVVrEnRmU+R2Z/0yQ0qFtgBXCmyapAR0xn
bytR3MaXwSWoIPN+ZkAy+XFpeZf60W+KjHyx9Be/1DNV6V4dlVKX6uzCKWRnbUi3FNvuRK5fR734
NZoB7ZqkBB4JE4AwLG3gqqUnhEoM5eS963N8otLFSs/3fHKEDTHfWE6bWwkeWAIiQ1FzpEGWwWJj
OWGX+MTmlGyDJPq7xIAq1uCsevwn4czvoZZzD7weGOfrTHrjoS6qVzovJEeegyjyz4mIYAZ8FVUp
jIkva2/NY7cdsjvKudteGimAIwFiU6Kg9Ni0Hs4i5BzR4KTSE6kBHuHS2gp0X7RIjRfv66nO499p
dDPMUawlh3o04Cchr2LKdnNnxxiULP+EYWL5bltEp+r36ibEe2V7Usd8tOp3OsZ0lupzL2ucA7a+
PKgcyKtKnMekgHoKKAcqAlk2yKUg14/81enxVtZFV/lilgb81dn38cRBm2xyxFMC0Ip2hljrUnsL
HKRcvj9VmrqkHGVFYTSq800gGxXmWpoJ83TfpWTTE7VBIUr/U+734FIBXQNTfbCVDNbMb0rkrcyQ
TQi3Miy/QGvf7/KkQ2zNMgGHFTS4VI2QrdIOx+yGKNdeiV4pxAbCBSacSqsWML6hvW6uONLQlTYQ
ZKrxauCeS6DOpshrufAKx0be4feJOLI2tyFTh7HXQVS5Be3d6KF4jfgtrPKkt9CYE8a2DDVTk/j6
Y3EKJY2qj291ckDLR0ts+mXfTV8uuqoQKd0/rgZdZCBDaPtL6gnXYfQ4aR3Gvr8ogsXYUZ3drMzb
cDcmreu7W9GTSEr3ixCycbwc1lm7Y/Qto9eFu/l9y57ueXVTYTy2RINxDmtaq3Dzy8DtfDHizU8+
OAq0ZMbneRaxovPQyGNhlXAztfVjrFzAefJI2rFxPLGqpwfPaaj+YupiC8dXPhWeaYIzJG1I2qa9
TzmIozpwPpsjx8x623xlfco5+mEvEXwmkE0rRRp68t3+upO3mOJVscvmf8B9LU1LwwbW0Lkt19AB
hun+dIHgQLTBQURNGgiGlxJ1LAeKTuVZVOJccAkOraBH8vbcXmSxnpsTx3Pra9BWLScB76VPMuqU
Jk5YJED2C5+zGGiwWH/QUVQOD9/IlNKTFzjDGT54rNbECYYwjkMpu1UKwnf7EV3A0veIA7fgetA0
mdNMFvB4seI/4Ik2OVqxxhs3jPOsd97ks7385op8FvDrLPvJ2f1zE3/MW81h6H8NC8+nefWxgRXy
+TAl2utji/20MI/avWomkwKHe87GxE3ouUx+fD49Ilrd4x+eyHOfnA48qfYHl4wZ59/pmya/knSe
0Cv2fTFAsejaMYk1DwOuAbSA4qh4IfdsG0FOt2hv2FdgqCQ0Wjau+aXzLASiwEAWCzhAOSemZtGV
IzYNkwdZMV7gmB8V6zRfGGOlEDP2BjBwde7QLIEh5XCm8ZFh9gKmebkY5XZSYfUrXXy2p1UwZBhQ
fZWeBdSj75dsZ/CgZ6pfk/3Upj+K6r5P67bZcq1iaBAaucTOMWhYmWu5RvV+nWRgzqC76OsQDPLx
z2szCzKEcOh26cYogTR5JcSnTqqGonyRsaaAQpszIE/BdERMMjaqR3BIipqMHE1dvhtXcH8HfXla
7ykn9fNO4H8XX1L8QB2eplPhbI9FgbxZcwLKigpaooQvNNDelGfFrJu9R4elhYHCmpq+Q9DXG3Er
4I785iTv5Y7SyNQiJZdDdjmDIMa/xuj8ahOj4/Tp/bFegwkcn1ZNbBLpw51HZMDUH9SDFbOf0MNV
EZ2kBnWd9kFfW5BvNfTYm9RWIeimdEv0pInRoS5JKqAczuJH5LT5DGiQB3AiZbc+4XLZcCub6hBp
yDTfc9viZGixiHiBvbF7/r4vAnSq/wfwoWj6oKwa0VCpuPeQxF9Wxis9rqjdFaOPMB/tbtOI2bQm
+4gGZiGSA3KIJlFab32/SJFfmY1zPcunybRaDzaD8iuUds4wWguAdCKcFjwWCJNLNAmjUd9uKQKv
FWh8BZWVLAG/rbo58eoTxXzaAfPdijcBw251R4k0KfaA5bJMjvmZeYNsrfX1HfrEElTJ5j1gbG1a
tRH9g8sEEbvbuhXreQo7u+8NWBwXeLtFJPJGNg8lUEUtFzMK8XypF9YsWdbgwU+scMuNI0jSuerY
aq2VlBFFUBoqI2L4aSml+DhVBDw4UZ/RMPlxNXigFqCFfmarPogb0guZ2ZuRzTiSVp1i1GoBBrN5
7mTf9x1Y+N81/C2+jNw485O8lI5nPZN1FXAj7JK+k/l49tzg0ASTVpc0EAVvbKGCsmnW0vOgDNzk
kTvDDYNTdft1e9Mre2J8xA++pqbIUHjS1gVLKxfjqAxa7n61v3TfcQO2oqY3sERUbAgNVZSuKWap
Ci+XABQnjs3j0NI9mBE8HNKYMAL0M1HR6Nc2nbV8+1qB3fQDH499tQc1T1HueqvsH/teIPEkRzLG
Q0CUf09a9j2fsoWYWwm2DeU6KAk8MDvpy2rbxldaQhhZJGpD6Gy48XX6ccmoP+c0NfzdJ1Sxeudp
ZJVgXiJpABfigb8kn1LQI8pIDmMfOU46ChBFERHjTWESFpSz+7sFt9wnu67M8IbxGa9lpw/ITyKz
8W3wyBT/FAQLWaohWarnIc4gwrWk/uGonC6sFtVC/VOSTcG+BVXA4UCRwsFjZhdVPzSyzObPgtWc
KYPsK3bvcU6CBpBdsRujaAa/l9TkMDhpE8keBxcDPVr8Jo4QQsXKSRDIbXHCaALj1JAER1h3E99s
IhX9QlIh0Pyb28659T/vL8WSrjNEuRU/ViaYcMS9IpNGEgqtLI8Y0yto/1yVitip0QESp67o3RZi
mA0Zqymk0joQ4s2bLuy/EFS72gHAPBMLHR7bA8++Z6Dt6EA9hJ+j8qN9e8mureom0zb3wxpMrpl+
1NOgBDh+jL8Rsooui0HGeCb9mcDzL+dsWkIqu1H6kLckDqn5n4EW5a+/HsFSG2ELLJTJqa/wPP9M
Dbtq/1KJYHcQgOxd4DqHkE1cArQddzBVWvIgGxEex4VfEbLmEM5zlhzOuw7uluV/iouh//qOtkBw
BEHHxVR+/0PpSWc7+y8mc9+yrXrCpsi9saaMWdlQ8FLbvuPFnPxfVVcvDUKGr+zAq6yp15jqMrDs
qFB0/w2gC5cyCOK4tbU0xqYGhgRdUCUts1Wkv8PP1GwPM5D4O1lwu4wA2Y3+KT/LbVCfP1Xfx9q6
lpKee8mt+nJZnkn1ojeOqhFL6hgVAsMg8gb7b2UhiBP04W/JqiYHjrt0I790LLO7NFBW9DG3325H
SrcJIPRI4j8KePClPt4OmyuoYD4LNjO/kCedEUq6fn9LcGj4Tg5Pj869KKlj7KX5j7VRaO1oitaB
rdvsoRMh5csuyWhxFrDKfG+Wdh9aVvCgyzCb5fQ8vDk9X6dWS+w22xhhzBRpBKHhvzjhXZHnP0RZ
W7jNFPUI9Xtm1RjBiL3WKke0XvjwNURv6K4qGWBQ1f3Ty9bH17OGsd6DiI7wQeWbfxP+nktviGQQ
dnVT7tK3Ui2CZ7VrxBAKtAaALclhkXVIlq/n8gCZbZ0a8ZvJTexOVKQ0vJ7XBqEm63FaimISn5jI
dkcs/JCeQkTbOsnJUO0ld2eXk/tTrTuWxo1hW3dR3Fu9gZDlAl+TLH7Guyow7ttQZkLgBvEdfDkw
wD1VbofHz4hoMZJtKP7SzQpB+KWoVry0U9yLU3gha/6IMMC/X7ZLv8Uqueb4Ydvbu/gJM/6PN8MP
MAkcQNRaedX6HkHtRmqkX7ntnzenjxWs8YT8aKY2fQEAVOZqUIHo6RlwR8/LNYDD9aTP4f7KwGYn
g2vzG6+w9OFHnnTJSyaah3Jvh2/dg99eX8u5aQ/4BykC75k7JVLJz35Jhz9QFC348qMTEXYvxjWl
N2d6xDm2jok899mMykqClBdtMMA8yUyblSfcTIkjpHAXrIZWhEm4vNkC43Sbn9P0lITh5s8TA0IU
PcETokosNR7YpTAWCxH2fFiCPcbRons11yPCCsVNO6S6jnShqDVd7vOGPkbp/90VVObLws+f8ZeZ
E2jgjW3w/3Zq7J5sJZ8nl3gvgAA49gGjeDTA6KA115KZ37gfrwkhJq7v9ZOHcH2aKsC2w5/6byI4
+E2/tFQ1ccp+l3507XknyJ5CyZYQ957lSwCt
`protect end_protected

