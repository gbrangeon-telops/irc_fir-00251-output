

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Zt+Kvzwu2Ua/vrjhNueC6ZHFBDEZvqw7CYHtLwQCcRpSvR8qcFedNcWPERpPju3eJt3nf1a3JFkv
PrBPNZe2dg==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
BgYona2Iv/0k72I3J2JPeYuzuEtaXjhj+ZWCoU9nVssKXxrxRKdrDHt5tFvberHeN9tDv53k+E0+
zSJEc8s7HUTXqNlaEROAMDRbOb7ChasXXdVxfl3WOvXTlUGfsx+NSKJ4/HfkR4Zaiz3A3zH3MCLl
LSzFeWSNT1Mt1+XG8HU=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
FzDw40mQxR9kpm1uxLfUoItwH6249dxMvWlSzzE19zJKjsyLJvf8oLgoShFkGPrtSiP79qKNxcUe
hzH0hyrZBcM+hC6bI6Mi60dC4BhdqclOgz1qMMvUNpZqrzZ5JB+kSMGHVFW8GUXvnFCCxYuu5mP/
ywkJGUeSDVEZY2th7ObJJlKEA7icdJ5tzO8g4W6w2f+MHJPOeHFy+SupHzB+1djuSlirLlm4nhaI
hraNZ0zRKoeVe6z0EIEqhB9JNsFNiC91BziwCnpzBdkOsKtsrb3RxMWbRRWbmc0XLssKg5Ki5yKr
zZaZTZk48RIng0NJRYTCGlINVIuaWueM3WuBUQ==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
gVm/uXv2qQX1H4bUmXuUswxUb0GUskWeA1MPfdTQVCi9Xt+VdX6mOhlgO6EFKXSas+dhLpimNzTK
aBHFEULIiJVFga1QEdJchUQ/rBMO2ShyfVm62wP8vvP25+deZ0Ac63uVlMRNhE68fori8KTc3x2X
Z6Nr7gpu2y0w16PhA7E=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
UyIHMrvI7wZyM6hLJ4gE4jKiSWW2iEuHADz2BcA+kHWTu+vXmBlODWfGdNNdgy52INFMV1nxlqnJ
XDvv73yssq80S34n064XoTXJBVIQ+OApIu1S7Z1OlLjdyiOtUW3Rq9q1U3A+hwbuiZ1x4LA5dZoj
5xr1PfS7YeIFNi86pALVL/xngSOmrya7h0pb27Yqn1ZWp+ZFU4zxAnMBdh6smb7IVFLN7MVgfSOU
BFsRwVHyMW6sC4c5q5LyBHJsVE7Cty+4Vqow0WWDEITa8OtbnNcM2JZrP1+VHJVzH4AYNHP/h5/v
rWvTg/dH3ZrlceYDFRqzQnHfQLNZHJkGerETEw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 42448)
`protect data_block
T36NOtummwygMYmXeLvh0BwJfoinYGC+imtONpx8khvs9dFAH2WsqP8oJ+C7YCdDmlOn1DEAsOfL
WSTJQyItQgppyX3W2Ujq45HOs+/+IJ1OzmLf9VWzK9FCKAnYHHCvRxUNHRbn+fGtDteLcU5P2JvB
8F9A3zZGWsgtUJjw+fCfKQOjT+mm/RlUxLOk00p0aP2nmt9l0J04Fk7N8pahUXNfupK4g7L0D3jy
WFFRkRXKSMZjPkp5CGe2JhxVGmBBkoDZQaCTcV5gfWMFI2YhVmiqwY5it3Rre8uGH0zpIHcQejH0
hJFmB/LgmVGVy8MeCgBExtwk5NtqztcPZQkYHr1Ep2r68Ucz6tUU0rf8bj6vHB+JOIXmBUmLDWtU
mm6gCsO4mmCisOYpEEs9cRuiywvfkv6pB55UYQvYCCLvnTR+LmVpYh6AJ2tg598FtE5EXAZcyHE+
+DwpibS7oszPGKQVamHYKLnjbxfJAmDDJVlZJwmVNxwFQ0i1eWNG8s0hCiTSlcx+He3qQzYwkWsK
ZY4YCsZXchJTcDUu0Uwf70HeHxygyroCdabD/H/qA8IcxHumB6ztum47ZAZ/OTlAZm2kmox+7EL1
0D5apSmkC5lYi8e2zdx8WKxMb82oDlS3JYIjhAlUwR2QkV3SLhDbUrPtspyQMYRl+lvhPwtVU1uh
6NLm1/LrId3LqF+phuth0zMsbN+TfZDruVl2AyvyRn1QWjsFCazgtaabTIl6g2HPjMQH0+CLfcEL
nYmcb2dwOuzg63zksgclCODsCmia/fNosccrt+nNUgqp1tG4QtlFrufNm2P192McVW9GdnfHxLyt
nDMWeI0dCDiSFjeRs4Pcas+RhyG+JmfmptmueQKp4nZlmaP7RwRiS4Dx6LzsyZlTlzQDtyFZTt+P
XKhQwUIKQ7v9Np0wu8dB7XTgAeZ1tpfEzfaEt4ihBVssxgYsPl1FdpuLfGyb/jGHoTDpxLyN8aQD
krMFaihLrT6hGvEeCyNfxmYrSS1ZCT0RRTt5TLO0RA6Ou1sjPTrRtyvjrwdgqprScuRV4EuzcP78
o6ZhHG2s88yNT1BQC+Z2xaqBqwBjJl61yw3Sw+KJ2naGdPorGsF5Tm3tSgxwMt6TShfI3i6nrNVN
mg0Fr2I7teKn4tihrh/CrdVYe63bwB+zDaZY0yqjBMSxojc3ORMblsUkjBFhR5tC9HJ4rmfXf9E8
BhK+YYiac4PQY+sSDkrqhKswwRjmv8ce1CjeXc484tMgaD2xNaLYOafqi1EKoze7wEyRCSBnymXK
bzh5tMVSOOUbhaTmIgabLUJoSxu2uORDJnm8GjOPR/x7F78PSNt2t9Vw1Ed7U0GBljVIw61K3sYZ
BqxcZJ/u/+j7m2Aaessnrxi4qZIrRlnGJX0XFsAs54RGjaCkf+RczpTxnH9RJEwIQj8zvE2neUDg
0ycnVaCNmvqLMxXj9qCwc8DQgx7o0b4Iqk69iRl6G8VzgAE14xhJNqhNw95uVH0WPZoNPb6FL3DY
B3VIedcGGiHyErE77eFuw+5OXXk6HYjDnLz+XzhjeErYDQqBgUpDHyy3FKy2YmfCDn6xt4GjS2x0
ZrVMN0D2k8Fnm0tqY1P37SPTGrD1VlN7gncxN7hfNksa1JJ3gSMk4tbn+5wqZ8zZqeXkF+hFf6l5
B4RJxQDkOmd4XWtAVlE/jdmJ5BNX0NaDy6a5jix/OfLcAhA+j6dC9Kl6A4GluIeM965Bb/VRizSV
vgZdhx1czCW6C6IYA95tINqCdU3t3G4IOKwuL+1NQ/M+zkF7aGZvqOkUlLj4zz7XTt1b4zzR0ySn
4IO6sa+EswTRtpZPGoqkzgn6oSiOqWl9rUQROQU/W6IU1Hegh4lN7Xf4UX4SG5jdejjKcs6aBAn4
SB8+75H083y35mEB7GuWe1PRkPNWd2bYSaAKHnT1MFUyC7qjiifAnGXru/rPOF5xuVIXcwVKjsBc
ZasjVWOrkzz6q9EjyO7S4m2kuzajbTP0p5RPyQ7P/hwZnWlRr3sY69r/EDRLrnRbeJH6vOUTWsru
dYqIm0DVyMxfyMrJqHhHphWfSTBRRcg/naRZnEPh/brDY4RgAssLo1+lxZlYX3UO2Vw+11d22bFh
l5+lftvJGcFFTOY3K83aGWu0RyiiC4rg8T/v/SedZytJUUlgyIVeDXWvARUrqyI13rxOOFzw+xUa
WSTseliUjP/f2Gf3D70kOxjJPCWVcXf7xectk26Nwy0Tre6sYoCRr8yCoVpWt06plI6kOJfrBrar
nW1zHxN/+mGqwt2L3SVYo8BD7pZ1OzMB1P5oczVXFoTie3e/ILCjkIyo8QYh35ft130nQe8Qsa7r
oql69+4JVFFBGNEXn9dJ3ZD6sUKWtsSdRaeDfpyARrsMcbCnP1x8QvwTlW+PUgLr+SVW3R2gg/3B
CDOel9vbud4eG5CZILgR4Jjrb1/JCJKWbexGmIMVG+QUKfeChe4fgj7ohDsWh0QhcpCMCvoWy/CS
2oaHZNsBtLYmsT0+DtY+SvUJ6YpaLtp949hWFwJ+F99ZTOpTtYQlpeifHcc1itddYdsBAlUQy+iW
DkuHr9zcDfV7TabBxZ48zptmAIyTBGGTMd1HkDyjkBN487V+tzbSsTJJVbQIbkWga5hcM1FieioU
wUSTJrluPFAPjR+u26dugpFRxHbvRu0yWaya/Iyixb3M44t15t4BelAckZx+Pye2KP7gVPu4sb/u
3jQC7wwBdW6PenQVYd0PHJ+xKBe+XargROsDGMLny4bT2l5q7BwRpSHxJ3ZNF81ZwMg1jMr/qI4Q
phaWt7BCL0Ex5vyCps1EyiSCF9noA1yZtMXcXUl/c+Aqovo40vuLiMHcf3oLSFG6Q6Mpq6udJmBl
736rVofsF/PRTU7yiPYVd8ILgJD8F1/uzdffJJd3wNKyJlfFFbZfdNGhCPD5qiD6lpg/n/tZ3Hi8
lMl6oQsrbU4QzvGE2c+rm9qTgv3CxtXjaOP9kCdyzSSef3FsRLaoPrzOvf46T0h9R+azQQpU9TP/
CnsCQIPB5Ah8AzvlrIe1KNvbI87RAqgfnGaao5FWOQrYgbSt2qA2kRVs00QgvEnYsa35hQZw07E1
dgJmDm/iPAmbRCsG12Rr/FOKagSzvecoeuOfB1OelBI4i1/GV7jquUx14R78nBPJuSSq4Uz/l1w6
XOjHZUVPG5XAPo3Eb+3y2SpOaa2zZBzaAlsbNvfin/hn2NQVaf7di/twl4DF1vE1JXinMWYVq+Ra
+Rdrj3VhJjtGcfKMchgDGGlEKB9EuFgt7lh8ag98x7+H64ewCGXLsFDkIGQdWt2JdXPMWZ+/HLb1
JfLn1VQejV0QmV3fq1E7mEch8MW6FBCcdf7SAY5kMqk0n80t+KlqhVDRJ+pwyJUdJVosJ5B6cXrW
GscPkFVSxnRk6GVqv/l8isaOshYfjvwcm9JjPGrRib8QyCw4eLsYqGg+bzsKy8Fl/t2KYKL8jbFZ
jOeX2lCGCArS4cXvOZdKrBmoLq7G8/ZwSzT2PZCXqbsjftVHdw3wbx52mgKOaNMcKFBsnsmTzlS4
blXnAzmym9xW+h9YkbeWmYC7Pdj29pfCpDKLh58peG9qYTJZb6tYyPbojg3kITZKVhEOhOL2AQp6
PsvSFupVpRWqOKUE1rHx9AViOJi/g5kXta7fxClz4VFsi7efF2t5jXe/S2HHhMmJXgTeXySLT68l
b+NDI6OFOLnvTa3YucUN2O/fuTtWukCMMSzv02zzwDjn6wzLHYDDdL3nfFBHlqfhbF/TBPrAUyth
TdoFDGHL68QjeE5tUdk2zElV8fBvIGHkd4i/po3GRwSmz7AVE5+tdSJc7ejoMuB+W77l+Q67wVEc
m9LhH0MkKpP9hZ6PCqjJmvFih6mX9u8NPtPtYfOav+pyiLnZWOLAyiedsTPoevd8WZL9MW8QfFVI
t9UlAHeB7qrX/qa/THzcP8+vFawi4SYcuMbfd6toNN4wt9mhP6zkbWBbP/A50z9c6rZdioa2rPOP
BoIBZd/GDHHGxYYzMzk8Vj8tQu1QlLyf8eJ4s+4hbABKm85DhJrHRFtBfUXoK7IzVrZpMVXxTNRg
o5DWeBHn9A9WkWxtyrbrMgvoXg6qm3GkLY7wbZNUXY7I5KvzzJ52XtSjniDC9ff4RS5IyxmXes2J
/pv4s+fmmgOSeq/IO1Gv0eSjyuOm7zA6rBBn1cE+NL3nFsn+u7+TSZmmKA78qNLS0KB7elPIp0nu
ic3Xg2VsP1ss4GxTU7DfJbqNSJi/TVktTr3BtAdd/sQvCIG9vylWi0gagV98uMgHrBqIIn5NFW4G
2KO5rLuXhsWFj23s6LQtwdN1U9VVrVURfGdBHrs5qOAWXZIJN7POfiZV1zYoSeyUsBE7H053oO8F
/MAdmP1DesLVpfMojIe7IQvP5CulqPFmbDH/MFF64JijF4FHJRDzmKRawVX2gWklBTzsdcjc1ItG
wB7HZYMpZo4Xh+X+Ihe3p3AvFLqlreQcKGnnDR4QfHSRBMaTgpjRikjQtaRDVkQaidJxNXNfJVyp
M4XXbAVM4HTsjfJdSWDhw+tBuAa7/EwAtYATrD330t61GhnLJEgR3unhwo7aLh15rlEwGRIpaHge
ktv1PAwKb40YVFj3iInN80OwapqqkHZRqWWuoZUajyvL7f2fl0KTnNCESwuOSmiPX/4CcdqOegpT
zba+4t5wn/3pxzWIlONljUvH9lFbWDUp8MuKHJl7hNSUzjuqYanTYHJ53EcMwC4BWBHNbPHoyhyJ
Wxw0A8tslh+M5VZGrGpw4UOZJ22B6l8BDP5S8BctmLWFtb7/gGiqijehkHt4OJfue4W/LJoQKeQJ
Z6oRKaFHKV79E1f4JbcAZ2P73giE10IDcWcOCEOOppdzChTisoyvRYuZmiAnsh/eFm8jCEdtenfw
04Ys4q7zEk3FzgPyjyuKygtWiNBrRDHhRYJN/OxNX4lO2xNUNEGsWTQNVly6Pxn8OILBlGo0Ny3S
KY3DLy4MCds/hR9EPceStkeWFIq1JEUveTu3igMX3VoJucvjzCDtpQCtJEwFTBb4RWOA59tdwVXz
OoTH6BEX4hRYiTH09yoswzoI6KB+Ji1fa++7YbHZnt7BHLbHnLRCkJfGUa13keb8HMOU0kSawRJy
IVy2aJxKQn+X2Lcq1ZQ+DjKXikRpCS5NGTRomzRGGfHL1sNMRzQIYuzQelRNR1J9xV4TXxaN4bNO
hqG8rlluCYJUHwZ4mwqPrfJ99ylQhJe2U4bh4at0Igy+k3Di9n9A5aNtcXjSYINjugyk0tZ2mLCY
CENAnnridbZRwgTlmjFqJ3XKN+DNCsTzH+79Jxy86VMHbBIGKcG8wKWEGhKnhF8H6KIqptJOKQde
WkIQ3Cdpz6RA5EHXpHyucrrPrqtviPOeef15o8JGgMU3ofeM8lSyonaPmJ4KdmY3pp+HZg9fU5d+
lDCdvinTqHkSiCleCzfUzm/J3+eLK6GLzvRhAgmi1d3mheI+Xr+HF5un/zKEBo+YHt5SvNpmWyiS
7pNe2VSD66Q8+K4HXyEUs5Lvzb/FdlEvxmSQU4n0OJUOzs8l3AwZSsI+rs3U0iGawP3x0evZpaoK
RmKAsCKj3R59MqXyICwsIspcg33ML8XBCAclB3UWRkl+Z3QDmelBFM0+rHbrbdl9YmEqEIfJF0UG
eyCt4fVxMImAsBeHi7xc7ePWvBetUKNZij3+dUBjK1y1/19yrRt7sGMJ/jL+EJ0iwY6PdAxx0mdd
Q8ONhtgBH+VWxaOsi5Cu5RexumPt5tow9CEuYxo0H8cbDrsoJ+XY9ZzY+GbGlvDr2zIKJmvhYriD
+acu24vOaNwG3wbGdcZ4dR88eUe7JoWsQoMfTeo6EC9cM3dgAQIM98rC+HG9oxYm59IrGtKBa8qT
dRkgQiae/zZJZZSvpSINn7mYH/ebC7lOOce4v+ueJMGUDkob3BxY7VTW7cfqV4RBRoudmCwDJ27c
t5XuaC8gRRSUG6gMQxbHUEsyq2QQdjuLQ+/oJRZMjLbXePER3MRGriseHAJRBloPu76GtQod5h+f
Be/ilQR9WtRKAryqEPp3iqgYdXqyAzX8WnAA61pmvTk3Dpi/Hs4MMRYwbApf5nFob3TYyUdIvzk9
ITUgc3Bq1zACJbD6dKmm6uGWpIOcG/HbvoiYAvQ599jRaXriLXPxzK/YUZdR0rkAZ/U4KtTUe9aC
WPw7vnoe4IiF1NHn+hX9LI1B87G+sqVTu0C5TlNDBoCk39bEp2QbiskETGVCY9v9HUF9BVEFbQOC
nMGC2AZYJ5NKLaze87hkrnULSxpXs0YVD20YURXR48CT7He+g7a9hdA8sC/yhtaGKAPPzZnscxjn
jAQPg2ZCDWNRW9oAb29hh8G9Qy3V0Mk1n7vq63envB40LGNE9XcDdv0Z7tAUkYOp39NaNgxbUJ3j
snEVTE+22Z/T2mxE5pkADFL7x5j4TkLbg6FgoUilm+1HUOtt357ZKr7femGfLAotWFwunNVmM+mj
d/V5pN4GUucmJ2YT6YMaY5pRWA9XQNJ4Ym9xTvL/yKhGzRf22t5FwGskED8QLofoPgTabQccZk8S
Nys3fRkLr0dvwLwEdCrRA/4wbCsvbGI+rJYjMktzs+UUn0RSvxQktv+FRTX4uY4MgoXYS2ZCDpam
ZrfyExApeHUn2rvZnKGrOTiR+7D7accXINZ69jsfNuIQ4JpEQjXgl0DRdJ/pGJ6JB3U8JrwePZEI
XCP9vIQbPwmgeWv/YXA6sEdHNWKBiuoAPKv+2PmCl7Qt/p1p/YCVukzv/w32OJzvrc+sHC36qXO3
zL1o94eFYHH+f//9OUW/Y+xn42rM9D93q+Fw1cPhn/Me13lKPhkG0uRzdc1snloTG7547p9o7We2
BvyvvUEHx2hR7qN2fhKulmYEkVZf2zzvK4eteZDEcsTSUgAOyWi/29VgoXd9JtJVd1BL1t7P7XfV
VapyRJkV/+YirQsdo9Ps67O7e0gjhYDQQFQ/insKuAGBB+pUxG4cthrgDMDFhoZo6q7bzOy+PCn9
ECwU/OpE4smW/l2UDzm1ofCkUwz2ZUYeaawsU4fXAm+ZeZzPNGTzApvDs9oGNrf1yfspwoZJ5BhF
LccwMm4Ce2X5tBOOB9BnLpt5ClceTE/Bn6FLdbETqP3uV2Ec0gkSyvAmua6chYEvlfc8ZlYYaAuy
ObLY8rkkA2AMMoMf4ElmiXtE0g1wFq8hy6sP5Z39oYkmvEQsxeSKWHkx7TBFXRVOChpCbLVFOcbK
vl0j3tWD+Qh1NNvlC/cBOwl7bBMp27EGODPVpE4WkDQSpftWH5y9RmiWDlIjlhxlhwyOUaI4EdxK
6A/ipdqfsGJa+ni6eLt2szPI5tqDST7b+vQcWgfc19ciTznN0Rc5/vbT1CaVQ/v+qaSBrzevDSAQ
/OIyK6x4E8mE3tzzjgMgJc6Ocv179PsOoAUPij25O5099ZeXJ6BrVsEB9IdvpWYqxHUrPLOmQqfw
DOfJcOTq1TXnm2ticLpdqm6eRZJHeab7b4fi0lprv6Y06s5MHew+gT6d0/a9CF9vt71ngYJQOL3n
ZUI/vsjMLE1LhTCJAvhm+no3M9VK6eqJyJh+9zyN2+Y3EktXgzNpx48l3f3XV7AZsB7CtX4XlXix
W3MZ5HM2q9pbuiizXQqE8dwyVLmIQ+siL8LiqFLsrqvyyePdqwDgbUqQ1aDVbmZf0htNcrso0kZS
4Mgg7NJRgaYoE4C+FOSbEZr2ZAct138G9SeQtuTdQ8uaz4KpQOyi3WQw0TZLfG8+r+eBPq5MEX0x
dz4U2WZt26KR6e/DOvaZbs2UNCkQ6zv+Vf7CbdD8jxhuYYpX2kWwkHy676R6L2uisD8TXvO/83k/
jY26D7odVTc1qYQnbaZ/1CH8DQeiZ69IsWwq6TKW71XLBwjuoV+yMoQgmAtcskRhdITZ2F1MnNKb
WE4OR+msRG47kZtMzbm/6kCXDeBHb50XLbnDSje8Oz8Cd9CpMztkYFagY1mm6/9WHA6EVedqz7cN
NSpxIgztoF91IsZ/axM0VjxhBH6CYFuvva3f18hdjaxaEvZ6OQAVfsGisjr2En4mLTLcm/nt8xtv
3g/Kb0aomewVFFNsiZjpl/5FWrO58Q9l1+AwhZegJCYdLFOCb98iWsa4nAmECkQtrfFgK1JAYnVd
cdtLZHxnwyJxuE1p+e9BmFfoxHjYfS6inousSBNrIdzfEBM2Yhpwlp6c0dCiYkp8jZDQHcAdD6sh
3MbFFYkBDZu0CxYl8pHEAhXzgst/zk50m3+iGUDCiNmwuxoA5LyESEKN14gvKM/cgWXqmfq+XfVs
/l8F31NQ69BqIv1VHJwIKggkvUcxg0XYBSb7IkHUI2nCiBIp80OGwtcDH7xh69B4L9FbXkcNNQNY
5YZIy1SFCHaE4ofdhVnzWiE0JoAMfMX7HII4gDfF1ffSofmxeUn+ojk4X+1SAiCQ8xzUe1/eYVI3
ALEAHrz2ZxGb2PFXJBMD8b83pGPlSNs3YwR6GTRGiZdgZUuRmE6iD/llPseOglAxTS2OKvypN9wx
8OFhNJ72tTavrIGtfnE5ASr+iMR4LxeF3X6CM0mZxMEpHkfu2SVn9S4MeyxjFLXseWuIpLJ1AdDd
69jvfWZTDUcVyj91x42a6sPY1a1kBJPEYNsaSDLRv+xwqptRSbaSFzrURuzh5YRcSU8V38MB09N9
6Fs6zirtWe17fSt3qkdAr1ibccZoCNYzfW+pbshV0th77sAX12GVzLfkEolfIKSY9DKiyh6OKOFm
WTTg+4MeAhBHNkB9w4cf5V4Rday73gTqvgdzKz8YEcMiCo746IvRXbnCGO8LlJ5aVibzRlH8abmA
OB5np+6ywrx1mILYDnAkihsFzeMiCydYazYfr8hwdQMhofX4KmJLuPb7SqiN0BHVIsOt/xKtPuI/
jXfYDaugQK/LzNnAmQIfC/qlhzeW+CiT7/hNXvtpcB5H2rTLYaqZPMx2HvjniID7PzxUfVX1yLdc
QFJ6YoMB/+XducNnkQ/AGK4RIJZvCVTUAOxF9YuohBqxThJXAEJSlC5jvYxkXKLRc/NHKFNrAKTT
S1gwzCGhkIc302+W/Ca/mlnwT5ZW5mxGnurhDjBQNZIpdoYRPtgWGa/wtY/egAPX6gQwCVQK6Q9W
tYqc0eHYikaKLAQSF3S+fV9hh6Bc9+LsouBfPu7ec21MAKdZTOqIKX9APQooGE8st0I/AfEwybA2
d9RPDlgMUJ8rRVpfK4s+ITWnd99cNC7rrmml1T7f1L50D/QZCZYMQJ/M0Y9iQkK1w7q2OraRgpTP
b9RwN0wFx0affDSSajSRxO9Fv20e1aC136nMkK0FGsNymlL/c4BTHZgAf9cKjtwZkQKoNJvuiF0B
U6fRGyQ0VvGBJ8Mhhq7uvJH10h+AfQZi1nYTdcm8ng9unFa2wuZoL7DTFfGMwHc9W0nVbMjwC2HO
gZlY6mYvijJ4NC12/YO4hl/JZL/wvgZD/Srq/rm6oqcRvTs92tUS379Qn8OV0/F4+eQWb+7dKwPG
iRAxEu/veIfpnJmlUB0TdEAdFmb0DYr7QAPfsatB3pvTBhYizn02Ri36jcdCGKs+i3IhyTHP6Lhe
HAByWsFSZhGYXuBF8jgNw6TOCiSzm/zUkB8stLCOoIIpSNbT7q+s3hvtqRXvR/noZ1pF5kcqmcqY
WA7p96mEcvqdLgNDstLmPvzJUs7Y/BXohrdj1izQeqWE/7GgCFfdf5CLHW6odrRa+ifI1SNAn9nH
odk3oouroriwnIRL+Y5R/CrfpAMrye7GnHlgiCTFf92o016zlprhQOO9NczTtVY1f+0nIsuhrPDE
bINxqbJMr+ST3ArE2SgbVmrtIX3wXSpOwQdoNHgsFRYWyZr17PLgr6SwcKvx6sUJMtQVxFwzL07I
GNKCiWotfaWz/dvBL6r0PcVgw9z9sG0jDQ/iokIMJHukyDx1TSt9y8rmdvimNqN7jBoVrFNzqqIA
daEiGpHYge4gkOEY3vdsXjH2tJkT8SfCv1kTeETeuSGatwh3aZBbSW1r8h98VkuU52fYwyZsNaM8
LCHo/rcOv6qjQua928X7yJtdS186tYyYBWAsnUNB+6LQNBvQmrKuxlTVftMgpbFD2YoMg4tMR1iq
QBYLgJ2G6qhZrXopQLZMkcNRfL+yAxK1hWHGjAf+N3D8B9RyMQpOULVFFpTZYLpvs9IMJ2pOJ8+Y
zkblIJ6Et9OBAqDAs8xo3bpqAd2NaGU18mciGELHdAVZkQ4qOu+RxbyCzgP8zAm86ZPvBHMS5sER
qu5IlaR4Gq8eMnxfvS3zaaOFvAPfK01VkgrU/4IYRUka0jh7ZlyHRmDrwsAnspOQ25mc5eZy1PA7
gvm4ZqJC3rXJvbgUGezsmgsJ/kVTH1+kd4XG1gI2p6rV9vpidVDLEpBEHNx+BwSscyD9vcROjvlU
4zkxmGYtJIBmugb1EU0VmoXQmMiOHnjvS9qxnb/f7kUdX/SYXjmtvi+rqBdpC3ZiOpIHrWyMFSvi
XMhEjmQZV8FlL54eduUMutOdk+VvioGBsdfNDPlIoasP3fP/u2MHDBkuhcihCLEXmMT/DDdAuu8Y
DOsL/DLz3kmB+NWg+OjTSoGSeg4tmGFRRJtSEzeAVf/W+7P0xCyRVcVVuLPuxHfR2lT67TF8R6sw
o+Dk85f35Hw8ffDOBfeQgSOQtpwm4y7QvMpK4IUDoLDjZJnbXj7j+8nDFqeA3cFUUFUuVQzzU932
d4hPVLfhtn9R8ap6kj6/arcu/nfBCbeExzdZjvJXvUDloQ0yCS7CgZ8tF2L+bOA/zS8jpBehyrZ1
5l8R5Ohhqpmw6RqftQGzAQGbmRNa/D4pDfOgBHChb1+ggMJursjOUQuJ6a/C8Tx5Ffcut072qO46
WEfBMHlEdfzvw6zfnA6qBqkgwtw4PYrQkNr7ZK4VuobnwcbtEAVRSoBEUh6dp3FzFm50c3Q7pxko
z511C29qHQ9AabWSvuxoAwb94BnBytqtcns3yUBt/LUlZmdCtjeRaYAwiaMXS2FOcwNYPWBhRuH8
ZWQLuk/3uREwefOAQ13qC/8x4LrNAXtHFS3wqdCMIA42jmmq9+NXIwaYDPg3NujMcN3yyMDPJtvI
0NZyxnlvBQ9dlT4OUqwbwUPA5dSoSWMyYSD6YXAuKoKCZbf7Q3z+gA32/MGipbNtlRLmt0dXEAc9
cQwq7zA/HMSSlgrU6uRqwCpM3lnXbiO70ZToTEh23mSEVRa6xfAEnYwFV8OWFkc5SZxF+e4bz1OJ
6bxvZhYV4o8wzLME17Tegv/KnsG7gQzGsnj+naxnuC8XoS10D8Jd8bSeJFPk8hQzAsOFwUM+a0HY
lKRlosE28FimyQQoBt4ghuOiwESyglsDjCfHaJz9P5LMlKMfFfIUI+KVU4hyQ0ECV+d5mLva6e7R
2qflEal1++u4UEOCmYtUyFmecs6oTLPvLP95OXmQ3FAoKL/UopN+HhzS9tLR2wkvOW3wg9MC6G0t
+EHrl6z0Qoeqex2r6KqP4FR7lhFd5tK7xrSqQis67oxpS32Hg9bFWUCZ/VZOBK1xwKnSwGltxDvb
RgGVVXed1KsAL4uxn4ArvDyoGapr/QgMjFb2/xvGT/g6gUzAF3/ISc4WSWClgYggbZvHQC2gTm1V
wTexB8XM2ZFAkb9Ulk5IRq/0LjgqX3CsckBWXz4CBNGrwRGn/nbnygj9PvRyxIa8pWWIDL2sS+6C
Ze/BknzSYj8VVLOTrkjOrELPzKM1o4kYZ5829WbxO8/84tBvz6LqDR9DvElVxZ6d3iZYY+8wi1zq
l7RTZwaxYB2tTFw3OwYe6SYZVqvDUP6y99zsy5jCS91EUezL+xWnLvUgnwXurx1n5SnlfnCjfQBj
Ujz06rBVQaG6hjgwaSBdNyXJB13T4CziZ0ioy+bFqrUNVwkiWQXyW8FOZd9KiIjKg+W+DjBAvyuH
9HV8RUyeX5jWAawloIR0d9uw+zvx8KIGCJMhYwdKfupNcKqVMw1gg/Qcdyjw2cHPQs4LN5I77VYz
xMGlYpAKp1cAvIrEngB+4iUZrKirAWbO/S/wh0FxxBZKx6MOOeHLcxef8wuALcjwb804y1iJeCBZ
C6K1IFdwUTIQ9VnNnU1dGksdueAREXR5oiTcbwzvNEnPYuD0gSnrNFa2Y5rJdlOSvGcKFh1ntlfn
awXM3sTF8mcNWBT8+ckvsN3Qc97CTkg5rQyauKjAnbQTHbF2yLoBRNeAH6TJ39fWvWvX7ZzPwPVP
b5TYgjrSgbJ88XGB7GEEZHWdnORBelqg8AtTF27s1oMMbNXXKUW32PpMOXVEAOh5eHDZMwfA10LW
QXd068vLvxtBa/ei2ceiPL6Tg87hDpZ1tO+z8OnilT9D07XtoTMKuR4dYXh2ij7VwADmz3Bad42l
jZbz33BLGRCX6ik5rVHyqCUTR0rJ1aLTHwrJs/w+eIzqL+hja5cJGUEp82pS3r3PVRsBrPSgI4Uh
C/a48fOAnK7giYUH1LqxWShXFqiUhwDjfFlR+qX7RtRoiVkMMzWNVGLkbstkjl5PsXOyP2OTp2cH
lXKeAQ9ee8th8VOzVcWPQ/3Gj7/cmO7gB9Dcek4nLaghXPo4zQ7NnfxOAac+6Iy+qlkOc6Lw+uE3
TlU+EQze677kilNXBeUoFu6YeZjnAcWgsxbUMqFZxU2ZZCl1BBALk/qANbQpvog4UV7imewZz1Ip
a1p0vJfGnEJql4/2gwk3NWCOJ8SWyyK3wW1hjx0RcIZKLk0XGQXwgxoEuzmZabHlJ7RINdGy9QSF
w0srSC/m6Qc1pNOOmDRJbX+nOKVXzJB453khEz8UHDL/A81PTn9AgRrikOzW7KJGKwfpHyVHN33a
R2mFJmzX+9+hwRPwpMON45w4dVtmf5PAoCUsZ+SzUPs53KHrxjsuP8dnn32eZdVUxifDiFhUAvTA
UzqvpKdVTWoz4Qz57ojA7wPvw+3kFA2k4lvWjUilrNfwWh+NnhIPbeOsB6TiHa2dInD5iXJvFUCc
vOWZYRCcRgObrJ065uYNMbsm/+H7zZsHDVgTe7KLeL52w758sNYdihIKd+Pl5QA4CV1Iji4mf6Ca
jBIEzIqTqY7519CVuXfa/wMxBgNwVUj7MoBED0LZEfkS8wUSrKb95+JmFqomI3F262RUh8diyvHF
kb78JgCs9ruChp423XcABJ5B0aY0SZtXKqulzG38pkIFTWzfp0Y8RpDYQ5YyCDX81UvwZp6rbDjS
vDEXQDJuFnn9IEzHli6QdVJFt6U8S2EMgBxwKYR6rfhOw1dNOdoSHY/J6HCWFo/T0vMK5j67Ahkx
urBQ4Z9uoRzB6NGAD3hC26ttdPHiYTdNpzVwTiaElMxBr0Z6jcnOODhVOxKsKGDo8VZRxvH37RyR
wF6MyFhmWlndzQo9iMcVydKD3fo8QLqIVxyB2mgsaR0WBEqXMFkWxqwKl6sXXjGCUdYrHlFQk812
cBJ6ZASK5ikGjz3Wz+PhnjdG178XaPe16O99fuMA47088kjuQ4NfK7NO+eTwP1BPJkSOLdPIpA2L
+gLm0J5TGMinrYzyFmD6hyhhneb7PVK/L7fmM62qiMRFRDHhj8IHw0c1mlufpsSCJ8fwCmB6qSVM
yZR8jkRPnpvc+m4oCTizZahdx83fnCt9jEZgBD5uY5pNT+mpmq1tFV9O3nhlkE/7/s42+eVcEvD8
Rh8SWX5wgf0n4rbbIwWNfWiE8Z+dw5NoNdB7ZF5yi8kF06tUJsZn5ds3X+GKRFTa1iBjhiHAy30N
/k+hegzbwqXOz6PGJX82J2XNNAnXAJvnrhs7Ceso5L35BsYLqkqVUAwWW+c9xfZq4TOEAPjwmF/D
FR56lx6lKxadOYNXQ50tIQnYip7UFfWS/2bunaZpy023oKThtXJGqkoDES5qDVkNUXSsdyxRWoyd
zy0ikPiBEY5BvCl5adrm6lfp5LpenoyThLcHRURItkn6g0BpluaT69vRM4luLmlqk58IYil505Ij
NLDetKOvHxfMvVTexY1mnjhKM0ug/RCiGJlqw7v7rShXjAY6Yhixw9xk933cDGGU8Wp6kB4qmp27
y80nsFwFiyQ9ACGZgJcK7aV/ekT4H8PFfsm/lZvIuquPZGqn3ttHUV4sN+KH7GygXvr7u/qea8Ic
8ddpjex49nMUPJ+rHCz+4BlbVnFLOM4lL0q6uDqXf+6jg0j7zy290oY4BF0II09XG29C1sGDlwP6
PZDUL3f63KmU7RG99MSiT7g5jzqw88KaW3KzsjRYTKEtmXtLomNRbL1Cqz9/vKpOPRxlkDWgW4yh
umObIpsojM2TE+dK2xAlgxHSs6VJ1+3MjUl00c/TGcuq4RHLHr/sRUtgI5on20UY8ubey93Abarz
ntQcJhJUulLaa8+c8mhwggyd02GfRHSde6FvuJtaM8LQ9VKLkURez4wQ8XIhidQrRD9OlsSXVKh4
1qbIQ8azhbUW2VdToVURaINi8uRb9ZM3pdqNRqO49Qwpnm58hmkHLdFhGszCVf+FC0eOJOdM1Y7F
7sa90dedMjLReY+4AQrPUO9bjoJNBrZrwZMWteqzx26DMB3uGjSaxVUXd7hiWIrS6UmL1NQtAZvS
wbOayV4/1rFhUns/QdckIqJBtBMxFfMIFTl3NGac/lEfxaYOfMJWHliIiF12j0oQDDUT4qCKOhQ0
IZZzR6VysVfTSZ6vS/A8KyJn7cSYZ3T2T8hXBaGg6uPACsYKOftHU34aJWIvHlA8kCmqxqIeNNZs
Wkbtf0n0mBaz9H3pmpPNIOqryhlUhvTBbjwuW5MFIj9Pum/KYFvqhuLhsQ3fI93RNYvKLJjwnzPv
6mkyW7eCJ8jJ/bQmTRrXhTDQKHUSiNmkenj0NYUEn7hTLock2NjOCAXarvksk8btWpZ829IvmiEa
cKOxcBh7NCpDUge7dyEESDEHXy3Evaknnk4bH9KqFCwJSEvJm5mGXyng2Jq9d9gPhdBpzrU+0fDW
qmFnPdY+rpHaPsU5OECM9GTHt2bDkWyxhstdLypXfh87VpdhU+6JwAP2Bs29PXuMXkMMxh2I4cMA
612m8Sx/8ikC9cp2FXX18K4ugunpqrpiHrMlpmZi7kxK/2Tw8ThWl+ZoNjXmLyFmGmeqS/YY+biS
+hBhTidPmklK77A6yeTPWH8h+D879b1xbdgO1mgSR9FvwAhvoE/6euZaY5ZiWStRYb3Ck2yd1bnC
iboqqV4zZ1/Cq0isysU4M0PN4sZ0lNuUYYh0OoQZWZsz9Z92/pOnrhet0CJJJIJRH45MuGwMrpKK
L1At/x/cK6m5eWjaph7e4GJSvv2gu99cx+DQhn4DaQChwTyDVRPeVNRxPnDpWtoQEs2HGW3VpwIR
1O3+rnmuquxr5PX+a7yV9GtS1fOiVVNAeNdE39UrSJLjMdgotCEojOZJCQdpJiSBBW2nK4tLjrGw
8CoGxbTt2/E3FcCBwEM4M3zPrIhBEdpKdegqucuJKJ6tw7bUAj2SzDBzlvh4hz/5DJKgi24N6L22
mcGTbbOpClRIKkPnDCAQYqkG1zQmWox1fK0VIP/LBA+Ffd7COo4x75OnmQx3WoClsvyfhWXP0tT5
rbrGRiljtkyl16IO8CVsSlvV2ErCUesZCCpJEi0WPV1sNwGUsMY4A41/wCFZJb1/8v106hIiuLpA
t54l/xEDBvEQnngFucwT/1A6sb81FioU+aDcTl+JofPLi26MBfYMEK0wYZQwKFTOgwMLKSyMn022
Bv1P4E84tkkLyei4R6SpAv0qU1NhpZ4NVxQK8CqSAN9K8FTKUhf6pXF8WJooHIif0IaIGV03VxGv
nGmezShftBEB3QHVkZqlA9gSO3lyO16V0lYy8k/9NnXiRXFe23Mt4wF9HBfEvWrd7LSrPQ+JkQRN
HEE0winNnx5pOd9NHpUKVh13w1Wusn8abND9e23OC/qq1YuwgRPA9vtlWvCNsGPpt0Td8t9VBSaB
ThKlgD3fZL9mXXLWT0pGRVLS2OXHBgLJeGO0qOeIEzb6IapqtH3V4zJ6MkFpISqclb4xJYjzdK3G
DZE97zTCDwcq5Fdm5UpnA+PLbPdBjS+w1l67Hu6dCDAwHDp6dfIC5EcTFifTjtTJpJuluHnwl68/
lcn8Qv/DqlRMGX1ZXOteG8PlrOu1Y1snCjBca7+Gw/JyqoH2vh1baW70fvFJKOxfMZnqvfXWgwRD
qhuf6FtcnUGgOr0vXIr3XkwTs4B3ib/sk0NysGvv0VL/1howVE4pAMUdqLCQ4JW8CsQ0H6swS9A9
hbs3Lm/V18NzXBf7WpX+IIxDWQbbySIyXGZLsaToblV2wnh9F0DfuG4bDXWwmYqWCTNxHzsmed5/
LmVFfV3HbM1w6Dltjx55Yy5LCjiAULK/iwjO7o/Wid+gC0ofHh2N+Zjb3asibKH+L8cg0xqbF4iE
uw+W6kfoIG1WqvTaO0poFb7OcbpGrQE+HnYP3vU6AYvldvCSaEN8GGxKhQCVXcjyzrAqm9as4her
T8OcaAM/WgNWfJVp1+1v7Z55gio70WWUX3hF2vbVcn+WC7McZx8usX2il9eYkp/5lEzLnVb3T2Ja
nDRkAwWI261l4cKpvVr+tDCjWP6Nnh+m/wUt7MVoGlytcxnB7NbNmoPVGOenB9D2aOy4LYDVLfNi
vIo9JhSkIeCjNWsNHpv7AImg0KFdOEuXfMTKMCSxYbrj5nNuIoavDw0TUEJAJinBsCW9OpODdoIT
n6dq7Iz6kSN9TmnSgH+GuI6i55vGrhzUSXHGialD2IgxD64VXk/DxKi0zNm0lbpY09JLq6K6vJnK
TXAlAQtXEXE73DP9n/15OSQtv8Bilg5K/FVNFxohPmm7Emi56Yop+f5aJnunC6HS4b/ZlF4cAl8+
/eyvWeY7dfO51l+Ckcp+Libopx6TE3VWebG76LVkp4QrPpr4GFJdXpWpDHRBxMggZKEuQqKt9NGp
MxTthKyQOw6voGH0EPwa1pOooj1sPbtJ77mxUU/IhtKWM+tuMCZkZxsV74G6M7ti5CvKUgNiB2kf
SVTegVd075wCrLDR5QAKUT7W2/b0osAAOmrMGSwQJ7aMYSGXbfPMjEyEcgwG+aV+c8egEk90q3vH
Le5wYYUYFU6WMEEGmpttLmDCbOWH6LP1ITdivfYO1vtYnH7H0aRSbDUwM4zYtOFuAZyuvaUeWhuf
eF7rGwlq3iR3exFJPYm2tGZ/tM3Cc46X+X10BGXXCdhNmBtMY9BxsTBYq9yaFph6bZXOFMZ5rvhe
5+VXb7JfSnc31UIfwy+9EQgApQ979kT70b0EQEjJb/3qfZesinVD3yttj4AnVD6AnGvzhMjwz7Uv
ycdHNxfDTI4ythhGDY+T76ZrLqVkHLb9hEIe7iLsABWnoKwisGwLwsnw6sZ6HgYgxj5xpfshyrMd
nmEpPhvuKpW0BHS+60Z7JGYPoRqnS/zTdCmY733gxA7/ER7VLVkgwMW2wdwDVozwBy518IAcZr/5
j4tHeDuk+vWmk5hDXSbVHO5f1moeSBtPH8cr7BRoGwUFYiDPF41xNT1wVXd9Su5GwXv5+0EGcj0h
XBEdNQY/FzxuWmL5r+vt0G7bscc48kjvGbeLnbIJ+EN8xwc6pZBEmx11dK8jrCgYEo7H6+ReFG72
UruQ0cQ+bmPXqPdiIILwvB+d9rY80UeUVTpzJr+kKlods47jI3/4GcIOkWs/M0OkS3LAJtCo4V4f
eYfmRi1RNrBae3S2PfrDRZKyX/CNkJ/vBv4J7nwOksnL7kohyy7LCXO/0aWAUhTuXHJ4pnPP2glZ
EbCMgL3P8Y8bep7oS8cOIGos74S64571R87GqoNwNUtp0mNTbZAXWjWVcVOOLlA3rO48QOlotND2
udA8dTiieaMRim8696X0D3BE/WihQtb32a5ZR56BMySYUxWkzAeusDB4uLWTd/dzJJM8XZ4d8r0J
IGxSaQqTy8+LdtLda0CJysFBC6E6+wntBGj9A2acOoKvE4k/QVgZmpB5WPnqajkJeGUpMgn6+RMQ
vPMXrUZUnq7U5cmCKUBDPYVMDm0mfM5c8kmxXcp8gmCSCi03vDtJ8yjynurTe2hoBA1P0T+jXHHq
s46cnqJf47TU3rCNu9Wx4XLecyWBzsDHKcP192U4VoEsE1jiDgvFsUH+5QH72LF1NvOIFa2jl3a5
pne5RMkmWEmDCt3ybVAnshC+4eO9qX1ukMYhI3kSy6cDw7GTYvEOQ33DQ5CQrpNdCT8kr0nQz26h
U3ZUzsmBafD2GW4TnnJNsNE7+RQSRs0ht/dseYFklJYxjyZ1MpaB7JcanTgZt7jPEsrCpFxPnx7B
tA1O0fgnsi9/BNBK0X0oIxBq7vxEHNlLm9b0on0tTwyktAAl9nvuvATR9rs0u0ARIPIAvOTuqGYS
WmlBRidnGb5cu1FflrFFDwPVRXdwbRmrg1irY4k20Q/yFP8w4FUqXLzcJRcn2hFJAXUOng5P0KsT
DaV7BXo5o+ULGcIHGUXiqIbvNPjV1txsaEsvum0Xo6lfex25m1UryEq5S2sFrhuWqzHys4EL4Vbp
gqqzONFzmNgtOKTK9eH9gzRq9FuRz/5F9xpqJl9aK3z4Wv6rleotAmzNm1w/TNGLRKRXppK4IMRX
kUwfrQV2iGh4A6ROmLV973BEQGhf1fwNiQzRw31oUJN1u/KLubrEeoZsZJUVpUgLlpNbY/qL94Pt
01iYj8N4KQlqmRO0xPJYyluUoyvzJAUW1WFSxJaCftgYJBtTYoeB1NEc4hpFy7WPowH9qzAuso2X
DRa0jPgBl3qr89cy0wUsEjd725EZrkwDmxejqA1DkXM3GadwdipsmNHFpL4GIDuSeI0Y2D4Z8eNh
XrhWwOiq9brDVovhekN2ZhwvQY2UB+ImyBcWUYyCVPxh9two/2MP7r7lRIOFG/Y3ZphQk5UUlxOg
j70y0qcNwQuowECaLWfe+Q1cIspOP9Mad3aKqd+LzI3cSW9jHX7RrIUDhaJcPs3GP2ykF6zgtmek
sHgLd+wMd0BWrU3FDgCbv1naX7gsCxDg2uSt9q6NSpBwR+wbyXK2TfdQBLV6pptHnyYd4DnOgaWo
z3B5Z3cqz6DTPOueWNhVuJYB7UsazNiVwC1JuQBXrl7s3I2UWeL3MlJbAhHk/2jj8UCNEzy3YKk9
TOqsZcXj2eS+25jOyEAgLGgcO30jJPSPu+56b1v3PQ5fjoqQAPi4oV6gWRZudvd1wJmtQEGtcIZZ
zFxpkPGtrTbZ8svE+99QZg6N5TVKBwt/Y84QRxLyirJcymakz3wN1K24t+TuTavN4dwmWu/F4SEd
HVED6nbnuRt56rz4JW+WXUxyRAW7dSnLIm4BUB1SmnXuVULMLk7Ctur6KByN49jolHPm/vsCb+xb
VII3OQp5EdAF0JzmBpyZOEfvvK+IQWH3bECk1nEBgQfjjBE4Ac2VIjLzKz7paIzb1o3ZdEbAi17O
WVSmE+TAf8HaBxGsLzHy4GbMnb/Awd/oiMA+msBZQNdL7+vNl7pbweGVEILXkk252rVZ9y11mqYS
t9FycsgeFGUJXrtWO72SmK52WL/HfYl3TpOHlDwWf6oJaQfIg2ZTgMuCa2Dwirp9tR59RAd+px+j
865PvLj5UorntiCBSlWDztmnCdpTlKzXxirFFJrs7MjtSOd1kgD0ih2AQxlHuMcdd8+LBmgVYFa9
N5nrY0Bd6Zx5I47BBB+xMVmNG5ZQlMykbL/YvLwBg1X2gYPgTVzmmPVSUS66Z8jduIe7gq8dUyoY
H8UgVWu0tjjrOWLj0rS1+k5bw0XobKmq5SCBBGGQh5/RwzO3aSBw6Wr8d/fHrRtMHPCYYtVAufVu
CDP8rhhYD0e8GKboKjquE/QE71NyYSo3YPWhUF6Uezn58wiLO4P2TNgYZN8LTMAOhNzuNau2gm0B
KBzkCCkd1xIuPSyGvw6cilzzNDs/d/vC8oIFVd8R05DBWGPweVqoUJpwOEbs5bqzsnkwexVbzaB8
9Q8irKd7MMgwkZ8SUxOEIEiGIUMt9q520jg9qqS2em6M+Gkas/SXePSbMBQQwsQQ8f0LsrBOSc48
7SP7y0iZ+qVLSHkCUVjJzvHymfD8AvJXG4bwXsGP4jZKE5i43p1pZRp5BDZV4lLbuUtqUZW0VXEd
ET18tVG91JT1cvPVnwl4n7mRlixNWf71neEKt00J+52vuT6VannVtFGgH0CGABSl/s36B+pJhglI
8vfGeOltMaFi/ABBGyBCSoElE+PPcrjO07m4SX3XIcQOnganDRIVTJNaGOL3OZ5BvUZ0VwfzeSmH
pLgkrs9W684HY9TYVBiPJw2rX0ZtDuIPlGo4W8bmiMb+ME3+C/WQwKouI8U++ISRJlEO9sNwYod8
VIA4Qjt8gE07vydFWwDj6MZ7PKv6vmuEm7yJZnKJxGBeZclZAgnfj5Q2EQmYwAzlPDUBTULdYuHc
QFk9Sk3z0zhDl1/G/xf9a1ezHNCUZVepRyB6AMcZfKElNVgLTkzXg2U806ZrU+ZfyxgWROuUxkWR
1wVanPahajj05J4EeM70pnzne62OfwwlWwCOqc4SWw+1zAiEAfTSpgny5JxmaOILz5q5Cd0CrlG2
nUE3StcE8P76w7SLeT5UuDvFbyjZBjCt8DngkukO14zGnxyKtXt6ndVM5/dUHm6ntZX77GBAExHw
elyRYHH2IS+zYiwM0AWmrmbGRcEWrYNyNJMMP5JbL53Fzpjl3NqmPhl9ggkkvuDO/INfcSr0m0ca
K3kuqDPWTq07V26vDIO+qpZB54xUVlt8UadYRVQU5oj82xXDJR8A3IFZZjHg+0PbBgLtte+MzRvN
4kGLq1g9OfKCSYSGpxn4lBppYW8z9j4D4bSxaQXQ6dJZ7ehNtVewsgAFsYMe8IleHZHg70v4KxiQ
TEwdOj8bZJ12JIdHB00I/3uiSCv1onPWFdJE8pIgWWeNZ8YzlLT0Q1FeNILyjdD+rdIfnANvYEQu
t/gQrTmaNGxlpOER3h6uNSEi+wzzdLpTf9jLogt9+FdMBYlA8vNAs/faiKTZ4YX35yAKKboPzkVv
A5J234c8vEWV/nrKk8Q4aBUZqtJPqFqetLy0rdSnzVxji47CdDUGsebl1uQQIrAWnP+I2rVYJssl
AYddMf8LlTD7CTYiEwkDR4wLeIjOQ8SCIfTcPnwKEgbLWZQ96gXSBqrDf44bkM0j1J9zoUw3s2fi
MuGFdIkvEwgB9hWcnqNZ6JG6Ww5NboDjRA0PC2DqAn06owbjohjwjY9d88LYN8ytR9qfR5ZTN8Bn
dV4izokfQARKUtt9MgAKWh1JNvJP9cSq4vU6hnclDeYYR9gi5qMXSKjw6Ka+pl9q0sM1NR64jVY9
N/qwhSps3HyMH6gwnhsThAlzjpaZfyFKHbH0DDbXvhRY1lYM5F8nrEvLxNWRLv55mrvKmx2klHI1
APglkcKPbdhLFFQRJQ5Z1eNAqM/M4HS0lyGk/CghQxtNb0pbaTTY928OODJozBnCn+aA023KSP6V
6SO4LkjhLMYoq8h4aFBJLhyxKSzH8QX9ioxtFcW53FXdhOvWXjguD4Rpeg3BHzNMhEEHC8LrCJtZ
Dp0X+Vkixa9UUxhSQpqGY6/LTH/cG3DTl3/o+Kev7Vs2wH9b1zD4mN7I31oJB6xJ1zrJJFXwZpPY
mQDGD0rawaKwOC7AqDbv5uYIvCimxm10aJiOzn5KoHgipIQJEqMZL3HDj0/smriVw3Gx8hN++IV8
Cz3HkmLxSszKnKOeDMyPkuwk+9DciM9X49c64JLaCclynCnL4M70+/UisAU6bu7gY0rj2TMmebXK
nT0wmMUE3u4y3TDwmE0qFDf/UzgGATIFqYR6MSQi+ecIipbjyDAGVuLeKUYQ5tdeNJQyvrESvT1s
+AD0+Bzq8X5guj1U6C01PPZwsy3dCGFbpxXFzOH1FBgWdGx4Bp/C/yIx6ryt9YdjiIbjhpV6eqS+
ZM7rGOhsiaznfgyJfW2Naay7AM8mcNDcmhczDDO2t2ob6uzc3XrJlvt20gnQaIQQnRRzeu0HVTbS
gag6GfVZuqkZblN0qrAc9E4PQSuz5OVorXMmYf7UaugKGwjqrQz4+hEpS0lEilP2l04x95Av31FX
7ztALxtJytIX9SyxP2/Alm6EPKoWyoOF8wjyvcXS266IlDjq5ryeCE8opkwH/EphGXFOPgLzxiqi
MCmFCFHsD9E2qNwz6DpWKF4tSYWNcTFG46/JRAYU/QVKXeCVHOcQ8qoKaNtdcrLN28HszLmUGYV6
Enk1C716No3lFb6DmgIdkeihHH0QXzWqeNHuELJnzEmyePBVHk10SN0YZ2tTUJcK433wR7AjC1yJ
u+L3Q22HraAfsr+L2DwH3ZRfFkMzmdZXmNNot9h9NG3a5W3rvDbGOWF6C8fR1oR7cN1CyhsRQag8
S5+r+CnlGQFP86hNGoLjVT1BnMF32WYm8US2wedPPUENdOyGJbpy8GOcMV+W4KibWxHt+oxlq7Lh
UImjefMNLE7BGkfQ54r785LHDFdGM4xbDicBYwDarVSiicBwX3aV5RfyPPEig5LclfKBzVRU7mou
5FbSWGReVqyfYtOOqtRhPYPft5VPimUelQ+MdCPLYCCQbcGBoNnZdV3ZWvBxTZqECIfglRSCVzfb
rSIIzZRTUa/3U3UFJRKtagAjH9MOt7dORU/NiazRbPJ9S4i7xKleRuXCJ5/VOBDbdRUB9jwamhxl
9A+gYk0MygTv2m/Famrn/2F0n4R2RpZPCxEtpKp6BthHYJh5rDZz391qeMP/se8CUjlfMA7E4kg4
6t3OdfBG6zCJZLSmeD+HE/L/dnBxHpX+tdRi6o/GbWc/C+jhC0v2hHHYQ65AWgCap+T64uCVFcpp
gcxCym4qpS7lhSDAQt5Dl+rRDt0sWt237FLk+jSBc65nOhIuD4G70nAk84Z+6a2ypJgd0M6cajNa
lqvfvObtntvuuIQ4HlluGM9s3eWcuTNaZitbpgQXbiazvd7ghPv8pJmQ/O3ChFBsqWyFDybvvwyA
YwhwcE1b0uH/+djSYowiH70Z795UExARvPpoTnRhzSxHeIUfcnBRVXAQ+NFisgzpVKnOISfokvLi
qOqP/shFZp5b81G+KQm6hPwlvq+cMC8m0ZP9NvQiJzaJZxvVnyj5YcIaImSisUbx5YoPGKndw24z
G0GmKxYFoUU3xnH6FSoLRZemJTsURNIr37MTQOSvCwvhnwX1a/8slbu8Wjm2z40QXACTLN7+MgiV
0rNAKR+JeBk0DC3QWOnXTsgcBoMFB3GMIHfPnpSB8Pl0TrzheEyjqbvYVFkWmPgYkuNwTTtqlKKU
m1Y6zGD0bM7a+fxnzjM9tPOJTOsRlbhP7aRj+mn5KnFBgO8Rbu5y+OttXaJJEQpJ3CWGu+otdnaI
FFJtrf4Q86SqynM4bkkLwCU8dUNlPNgU1+Vgm5RxBh4TIVI/Du0iWN27i8FApz7hrAfmdSiq+BUi
bLSvlpsHc0UuY6Suxv2FrQUJUHir24uIxq22X0DF0ARZnVI45nuxUtA5SICKJblaov6w0/w8CPb6
SD39rSwvGr1l9Rp59ahK38YW0IkTO9xnkU2VPPNhldWN9sqmvLWeYwJNsQXGQggMtiWREgYkO8yY
a2Zz8qWce0trnF5cwMIcNeRc4P0R8LbH2K2D2oNTLDbznDDhnmGHl0AnUwBN675CxPzyJLK0x0ot
M10ChwYr8ASX9JDbudhgs2EWkeumWeaic+uaH+L6iPis2/4VHmAj1Gnxpb5Ag+iWtiYWPovelCQf
3QMmx+QqZHpv1q7QaU88KEzE8OFWoPshXjH3GDtHxEYORsb5B7borTV2J1DDHPXwrj54gJXT+4sY
UUhEj4bB/UUZBNtfY+AD9X7t+V9OJdctugcgSeCiAsrE0DnxrJqwyDfC81JRKnIq5XbBeffLRDMN
42wG0FtMsqDpbZuT6FdN0cr8eCCAVN9EygFTG63taiAMC+5HqZnCyjHVaICCvilvmETM/3EEf+xI
jWeyH/bYY9vxsjsHaHkrXRu/nZ3wyGfkEe6O/ypDN9VGj69qdGC3hI6BxZ6XT4WGkFQJnBn2xZYy
73n0uea893VtpYQFy2vZVVYK2s9ch3nYEEU9e2qVlHFMwlYDvynsQ+LWTEm7dEpGRRVe3fif0qMR
VkY1C4a+uthoLpLEHjoSer5SDZrxOxTFF1bhkWd5JyAx9ZrMH/AHFek/O0QKOZMSC5A8H9BvCA+p
PR1x0a5eTBrygnZPReuY3cRDi3JjrlRJYUFEbtzIcUZNVS7z9cJLn904hLOLu/pWPH/qncs5Du4p
d5lwNfSNRyVQ/ol/3fAnqJbNzB/3wugJCdElXRSSBpyZn6WXFQJCyVxZyY15iNd54/Gfz3WjMedx
s2Y9sZnKT1pAtSM2FRU0NCWPU5rdsQrXuzeGdl+OrctPVTej83r2oUQ42TUt7pqUCcJC1w6r8yYE
qdHawTlY76ilvfMYkn+u7YSEsgX60uFHV/SoS2pCz8QeMI7r7Q8d8gcqaH9T2gYPJrYEtVNQT6un
j1gxBWYtUc//Yp1HFO/r/hDX8RAukFM+xMCKIcIeIIn35FuyEb8Mt36fQ7cjSAyKrlPTiGAqfn5M
c312X9GDJE24gT69fIY7ZZmoexROu0HYCbBlrzlHbBGTXAcdUpyJ5gmE3jcjRGmdwYKm5JqmyFsR
81Rj5LRAJC9nRcJHAsazvl1/+XtsHDB9r8WKYclpWKT/EmW86YfxSiOdxtp2HMTkKRU68wmiPzR8
+4U+L2b/ROsW54+DxmIpKZxzOsJvXjuAVvkXlKrcYMse3TGx/T8tcjIxLwBUTUV6WiSKmWka39ez
uQaZtLd42s7N3mmAvc4D9F8TQGJcVK9FoMXCcov0DJomnuXiS8cZnggP7pQrjzRgkDaibLL60dtP
r5WfPY6YG5/lTamKRfavov3T33UL6XhEhJSmH8xRGMaHL8tyPZ0amPm2t5ZrLSjgym71LU5NqJwh
k81YWyqVMczDD9vZtlhAdS6uHAU0nwQggB5QQ1UFuMd041J47F74hK6c0I6B0jzKl9WqbPGI3O4W
sjE7+dCN1nCLCqkUCR6xgxnm90OBrgTbRcfexGtu/cMTNz0xiIOXIcLNGnOlz8DcdAhJ0K1d0zqm
d/vnWAi1pimOu/IVSqqzwKhogEZvEJoOCHllHPDuTB4JHCel3CQAMPfDuxvFFsxFlR8Wlrrb5UZq
y1hn0+T1Fab3lT1RxfzH1xP4QfJ/vVweh3Ma68LCFwCkHx+uSyPiVW7Q72F5xUbxcpph+GhwWE2y
g4sK+CufVjh2ZLENYpfamklfNNUJnaHRQ/H9GDdfWrYs7TYFlxIGldfUSrXZPtIZKyHrfAwhOPyK
PxMUixAsASX89p+0SEiUgwr++enRUKurk/djHIYKuLzxmwc+Ff+KHk4ROoTc5zVuUbTxAlafV63s
LmNyrOGv5tC3v3X6GoIVFtwoPXbGwZ7bm7tkDNmRcfUQOteJmplmD6LVLTnrGJJUADu5ETBSpefH
b/UxytowZqVi5slvG06hOPs/2LWZZZSjd3cOcJh2A+QfoPun2UxwNdFDRdK7iIUHCghrSEyQCwuF
tCGD8SYQxwFsxTpVpQYEeQfyXxSk7sLro+mYplexhw1UL5l3DVyfKLuE1A68eCLRNm07ibSefOq9
5cNHGjd62GMoNijcXwiCCiTI9LiJAh5gdZrJ2/6S9AO0RF6/JUyFInYKm2iQGGF86mAYttW54yU8
5stsnjbUCxRY0HU5uWe1YdNzs2PpRetMkRFhqk2lqB9MwMRE9mmIsCdtj41L1DF4QeEOgbPzlMdN
Y5wGU50OVWQJF6kiiLL5NXmWkc7wy7QxXCcHWK9Fya6sRWzE2u6Nq7DX3VwsI4xOtJHiGbjcj4qt
IUDRCgjBYkOLDXvMoeEKWFXbkPB1owADc9E5g7H+QXiYsFL+D6FctoPt86KaN9iqsjrpKpo3KKtC
4H2sIce/2Y+IaN+7d/CUvv+ybHv6bY+Wp560Wah1KONKpOEC9MZ5DroCLze98umgHY3du5YJFYQy
bUoSW4PmN764Sqg8je7YIzOgNak2T/hOwVdyb1IlldlsNrrJ134uwzLRCTk7Em4AdZHRuaettLhw
1gq7xsD0vih8j4wwUlq8wr7/ONGV8gvZ0SQea4rgk3BxjK7iaPFF0YWQfNqSxw2iS8PVJW43vlH/
s+VhnfVVT3xdAWxqWY/u2bboUbELoGz2NY13o9fl6U3XWVrAYhY6FltyQoiD3Ea7fXYGmK8MTp0T
tc9pT6AcNQ8JtEmkXTPYakW/j4+ey5lPeRPsoNHy7PZDxJ5iJze0DKa7PtT67IpCKpLH2anfCZbm
fkzSzvbwifrNLBT2j4NTGVqbFAgOBLmwRGi+mXMgYCW1/Grztfey2vpNbnx0qd+vDIWcNa9letVJ
JyPee2n/Bq1wAwQ+PHhSOPXAl9ykNS4/JmsLzqU2GNa016wS7oc54uoKZC8t5A3RiZ6/VkQqRucc
M5L2O+Oqc84K8N9oMqQJ0yXWLNjpURHlZMfhLLH2UXQ4ONeolEHY6PpN2E1MTeNGjLJj/T2W/4fg
wcQF1enhNfFQFsPOqxKZsc46TPc9SJ+yfZsiOjaTVv9YTTbQ5ise/La6q6G+2MsiLJGLv/NbDaa7
mtM00ewwcfs4q3aighm7TdwmwhEq59leFLEN6vB4rMHyIqC6m7zP3jHXQ2MR7szqiPfJniGUk+Fg
PxE04FMggV2Kh6/EIShmH9TgaE0T69BH67TZITO2+SZhnvbo8FoFWzlJMp5Bbw1JAPUruouLwd/p
hm30GZ9skGNQwWimm5JqBSbXJiNBhtnM30eXzzXvxwooblaCCy7jwOz4RQ2PvGEyZMbyUVg13jFx
BvFs7FHUSmOdjdt9t91FbShapNSpt8g/xj6B1Up6PM6+V4l9fC+e+kiCwPTIOywBpMoC2k1WG4T8
CcWRdHxhdwNrXto0Psxvf2LNAvt6deBguD65951qszaKo86Q2QXnDumpqTChJwkiAy+8PDxKff3C
kogjWjtOwC67923w11X+LQWIGnV57s1+SHBVj5jDQLg9VLbftTGJFi23nKrcuUHSO0fGaUflw42D
pX1APdkTBu2qM4W2DM0KnlSWlJrOSfRkFAo1PhlkPvedVLexrFRO8K8NE6c7LEx0jEllISmaQbPo
/Hrgl/1m20sX4dqtzZCviK4wcUnG5pI++u5NoW4JYMISjQ8rhbq+lFz5ON88IlCBTp2VSVDAapRR
UMxGqvcM7BvSRNKOkVKba0quKqkYpwojNxz3ZQhSxz4cmdnaKBuNA4QeCFpQ7dIGMWQiGXnlAZBt
vIe8HymASZ2H1uWnZq8gCmNtFf+LpkdYkzHIx+gvTHTuwzkvs94Tv0JzGYX6hzcIYhXPD4Mzlp3U
f+Y+GcknpiCtPQErTSEff8JfShZaVg7YG5FRj8XXZel9jx7IZovOz+8OXT9dWrCNfq1d534jRCUP
MNVdzE58QDY5zmW1qhhQv+Qnq0cr2YB0iRxuBTk5fsL9a77wEedugnPcop7atXaLbeuMeaW2T6rK
6KMlmcIUCVYZVVThgKyVGy2/dwC0BVrSq7C3LSlhYBkpWWFpWyfa7az9U6OiiNaoHuOHuUZpADEH
5S3VUWml5hVeHazgm+1Zqf8fcIHHO0MQnmYhGjVPhROC6kJjPIcGqkBlHGMgAuygILcqb3OfX/i0
AnfD+m0L5/KC9B0NJQmGylT8iefqlw38r8cL4V9v1/s5jJGCsb9fgescW6NFikoLE2bs6qa9kXtv
BDU1Y7adMk/9H5YVlE1hO3R9qtFRln6Xv8A06rYgCkgeKyt4OmULPRnIL5mlCWaEaCud2i09h6lW
gWAfWxOcxE7qID5f+YYhZYXK1hNtM1FuFPK/nEE3f2wff9d8knV1mMs16t0fcTIZlfDMwhUnIae0
GeHQ0AR6OQBwYjFxlqikM3XsRPyJmHKpYYDizqjuXAfs2WFF375GdtDLPmAprzwVmNefZBNgwiU7
TveqDy/+iVSkeNIZBmtAHxniznzPJi/acPPN6JGHUPGmRNgOQCIKhCqCWxLxGH1Gj3cP+nvezWmW
o/lauNPA8n5xnyrOBCT1HgGLZUJZ9PMiI/CdmH27hVkCgdMm4M81dkK11KjvszFm/DExuokGlGpL
Guv+0kJnLLQG52Eej+rJtadyiW//5NIFHHcyCHEu6FACm3Ie1lhpQ/9C+U+NoWQQYUjygAjOz/1B
8F4eZUXcB8/H/80mZQScF8pkxnkbKJRro/JZgFXb7do6Lf265qLoQibt3PuF2lNKY/xbz830Lodq
T5O8hziOra+lgZFTmY87BHAZsogQ2k87Ms08S/8W9lyME6EdjMChaXtVGN1GIkkLoyI4ez8702Jg
5IwdDQFlcSu/JHx/s6/4PoTC/i/e99PgC0Zc8xNiETpLrCQiXSpa2VZQC5i3V+1DUl1AcrikFr8U
b3sjffs1/o8fYRLQoGHD5Zu5CP2G2w46kYy9bw4OsDHFAcVgz3zjRrjQEcQqnnP6QK/CH4b0qQaz
7tv1EJ2I/iMB/VOyOIzeO6JAYdh4kZ3eFoq5Q0tMiBSsyNiEPQ+9UlwrZ4gV9r9Qpt6hOHHxrGz4
ptLGwJaI/AI0pamXoEQjdJCcS3LVbRdKkNeXErFX4NFzMH2rP0GV885JazCQjHShrojzwswAY+9Q
BCB9LOq8WsFZg2l57IpSFkz+K498QMg2Zt+5bpKwajcIlxSj/l0mX3u5SiCb3K/3mUUvOHDPYafO
hK+r1hMXRJGUwgwc0hTXQxMTATjDvD2dXqsbB9jMPL8PA6LIIP5rYDsqrQRmx25bt8H8PefnXVC6
dm+s+vZP1I8oxFudL9T5rEGK+1a2alGgc9Shvbo+GETt6wav7KLT0wde1YfFBqMHGmvhRTsjHe+A
2bn88AbjLTuC3uUxWca6NesmKQrdpF2UMgTPIXB+2rAHe/ffExGGI+8ruXDfatYwHm3apfAUSIuf
BIR+CxiAvQoIbnLFyfdOBXCrZNK48E85gEdNf9hva8CGRL4O4BOJ+XE2rlJWVDSUPfFEkIlCsttl
q13TTkNa8ehAujvSur8F10wnlfPOHCJcEyb95ghP0osqStZdONMnQnjR4cxqlFLVrfwV3csN//IA
+/dLRhHLhpgz3ZsyMDZV5jdxQ72eD7K2UlBDJ8D+oFeIp7gg/kO1iYXtJYsLCqHU5RXjlAUNdKrf
swY7axXcvC00Z1i2mCG2Zbp6C+iVKVRVA0M1xvkCpLdCsVNQB0WukeLFeZtr14Y+UZhfmjvF9XXV
1hwxREeQrxLySDcFVDU4bJjZ0Y4dmRm0CP5GVwjzkOidOG039dlazvlpdIhB7TsFBz+MCWBCW1Jw
57h0xOFU+eJ2Jhp68Fe5uy6NkKPORg0ZEGRZWPMbCJ+aBQHEc4bPJZ/HjZWNjXrNJk+NmDp7crBc
S7WRcisOesvVxrj2soNhU5V5LPzANA2ynBwiHsAjPirO37d4ra2t5aT3B0Ozx33OnBMt6OxG9Mv8
kQOu+nL1boGqINNusOlZcobjREEysBrqmm+aHDgkOISd7zpZ1AGplhyPKkEqNyUx7gP+cd6lbv7x
aO0GVH/hSHg/LCmTt2/DKIqf/YzAp1sJNOEqFK/y5p43AI9snSpmtb89R+2k4GA2H4bTe1aO67es
YH5rHwA9Awuz3oju5nh0vkPlUMZQANz4IfxapoxS05tHexpxVvEeE2TpeIU7Yl8i6o9aXo7KBf6G
zacdx9QsWd/3rmOs7D2xurGLKKtjhOOWAbEsegbIpKXqtz9efgJsgnU+7M/Azf7CYBl4g8v5vg47
jZgd5dqQGl0nHvZJqInUaXa0HvEYeFtxisA6nRynHgt1XZCP1twB66jCc3yRhdL3XTrznCXu/HiP
lHWJffSaeXIIQGugmC16n1eArNLj8v29gzO70Ygdsvd2nDC08Sp0c21RFfiSxJ9M71AcSt2TMuv0
WmyUr2wBg264jnX5w0942zP9a32ro5j7goFlDf3aymUWWc2ZCuOz24mqk2YsQo7yGrOxwhm9Bc65
H8cxb93+dQuZ3GhKbEfDn2pIrUm2KlG33BY843JYySjkIfdhmgORaOmQHmPNIOoMY9fp9ZTlFcYL
RveOmVBoWmapg3VEQ++NYjE57OAN7JI1ANrFYovWQex0patPqSP6xN2mZc3GtrUCUjJE+zWcVyAS
rdd0BtJGhyzuKRyxrSFIEL79HI3WLHrYzhSD3K6yz4au69m19I3nFAShf7gT6ehYyeg7E4oEjo36
mHlkZ9grHFqYrj9cEJ6OLok0y02+fYyyRM+/sQB236wtbwA8wnZ7X51cV/jQ2uM6U3JQjxvjVV5G
bw9js6KNG26WFygSvFRcaKKYkPNgxcRu9XLkRS5xNyXwd4P9wNuISipx2UNk0i/qiK7cviwG8Y+m
96s98Xko73PnY0G8rJ47+/kpiCVNAOcqWY79OPZ59GfHY0MlQYSwBllTYEgp+pEM5a3FJEiHr66q
I+qwQs2sXVUUQjgKx9BXsOBD0Y20iWVSD2zoy5HbIixBrj4FUNq53UZdDwBRaFGUsykFH7co8m0D
lyO6TAu60zMCoNdH0pfnX9FivYDUTBHJPqWOSvgKvTy9t/Ew3QCrhZawk/E7eja8XKqe0Gnhj79z
fTxTtCTyx0bMD+OykJW9KlvQ9A11stI/26nNygWF2CXpz8tSczUfbk6QM/3wyME7Vfeh0C6FnT1H
Timy1v/pLgeNp1se796hjcblWNp3ve8e5BucohH4WXpPo05NXiF9xHkNZYdMEN2rgrJR/2/YbgJ/
iPf0uJ0rmocc1YMSlyT7MIi2lQjV2ftTGt1vIHnzGJkiWnSaKJ6gKVc/P1wlMLX+EI0idUYR1pFJ
K93wZuBfs80+SBZlLNMT/Re3lVG0td14ks0Vq5LUOgVjCgwhCZpF0nMUfYQSzrfoY03orzLF5Q7Q
eOGL6dQTEZr6h/C+EDwx01rEMrJ0m9dR36hJK7wIKVAybi+9r+GafRWAD2AIQe5hrNEUoKUfQpKh
hBcbuvQFOt685FlI/o9KisdoLAjwPWMGn0oUbvVv51Su8oPpsvSE5Im3eXjbVARSvXq6X2TcyAEy
CsggT0tsk6gQdIYFCi2TJyGjIw7OJ5yRRS3YbpPvZ58ZRfaTRKfeqic6RillAxGF0/52n/TVT3r1
WhsFjXC94O/Xu9hAH7uq9GJEopLjvQQ4oxIx3SXI97yhNs9Z70jR/voS0wnV3UixTWKA3SmVa7Xk
5qIfu6s834HGrv78Ow3wujOL5KZZEEigxEx5JRAbkt91gU05oeoekvj5vlIOeVoM9IVLrwfHeRdi
yDsoPt+ALtbLtxH2jR7FtPYpbHWSCGU2GM1Cpnu4MpUTArHrnjKqZyBDxWGriPOMLCvGlGSKVqTE
4/Ybk26scBVJt/KGdKD23FGNbo+iiiiihojsDPH3XgtnyKnz0Szxb88j65Q/Wr3N/7aByf97FN3x
eyJborQ13ktdr+YiE9PXFQgm/5dc7WyiaW7Ayb1x+/hdX8tZYlO5wNjC36jRKbPAKscccVslQDvI
sLetWX2qQX04c0EXfibPrlW3kWaL4OVvGdjxZhr9rzglwDLZgIi60ptg/eFxJwhjCdvXBiDggDfk
imRJwamBszw0cUR69HdbkcQlelVxitfZclfaon0vlTfU4UNMVKFL7+CD+s2vqNONQHMP9pV7nuXg
aQ/857eRY3dZkmeHfR6rKbOfvjLf0xkqRIx+LU+RJcl2LC6ud2gUipW5zKr0314aJRm5mQbPEo+x
EvBqq/Rs8gbNiPz4NNS/LDS8IjfBXSpXjzZDxAAn1mntC0/02x6KEZWqkljWBv4IU5VHideNC+rj
vvsxsfNkQOxvq9sbeOzS0wnkVQEr/at+WpJYY6FhsZzASlH4vXrdPzK0bElWVXb3pqozW8ABNQ6S
aqGiG23/K+WmC0VSKeIIftyAgqWJDeEjTXoEDjMpO9QktNpU4Recz16EF7TzQccr95CKn/lBWSH2
EuToFrA92sS4UxZiNy20p7mcU+LE5i0h85G8RyswjDT1rWTNg2m9UxsLcRuF6kZpH4TSbNJyYsaX
LDb+99xF3DrQ7Str3fLnat20HKLODFybP9kDMCve8Uev9OYd+9Dm6ytkEPZo0P49KoGfIhbjuo+O
5HPgm1Pgh9d7rRQfuUj9bgQFHAVgH3tKNZ3qIh8IJzL7midbmfiUCega890hzcgCBS+75A5jAXGi
t92XHFB+3e/A4b2/k8QsOXjRsX+a6RI1UYc1rNS4RqoM2neh8zLNhTxBhpvPCLLw2VG+rXc/8klB
tzjGk1KXOHj28Wo/TfBEeimk++Sg7X38sYEZ1NVRShJ0fHVnBks24JOm3MYBky4RqTU/6/DLyTdL
57Vz10V7N2eg6s/1RAq4g+rfPOfSqcw+29ngXRT7vB7k9XTRrfDEkRl076BKJdLexTO6LOAA74Md
qL2KNbb+AMm4XYryO0mxnZIwpKihfg8VrUPTmbJASFqq+dHTp2/7GiH5Yp8FqR+RNiMEJ5z/iTpB
t1zWCUmEzrLkLp9Fy9z23QFdc68X6TNgbQsRs/QZBN0kMQuzMHERtPPsjakKHav9LwUJ71bkcgWb
eBZ84agehU9Me+KXjEf/lrXD+92pz1Bkr7WtwC+M6Pmr/Kj7cg4gPQKz8DyiCkLdP1nnrigf0cWc
7+ZQ1U7np+nz+4l9yaPVQM6cO+sury5Zz2cpJ+8tfCghju1ndAgoTsqCWLS6mOKR1K/nj1grG94K
i5K4PGi/nFtlAxPrYJP+zK55/Re50poXzOd3zUTlrZq8JQygelqmcOKneSFB1TZD7jLfPuxcvwC0
LLwJzx3JvQhnPynp4Awje1Amgx8qpNZwMDrBRsFn1QoxJBGTZF1noYlCi+Kc2YyZiitkifYEZnBi
ySgad9szFL07/Z5nAacYcTfU3Adj7myMU/R/GQ10IRtt3M4q7RL9lG0vlydUI5B6ppnYOthQ+mmB
R11WCBxZZUm2j71ztRyo068y3kBqAF3RNo9l+DJgujhyjRjIcVW/beg411eql2qsztyNAlEs9EsM
6KVOzmfk66gvb0hwyVawvCgYibHWYjnICzz4qP6KSivRFmLYtTwocglqlsj/K1ZzYvO+67CccN0L
MGrXXKYCdEyyPVaFOJj3/HGUz3FBS57eFXkLCypZUsGI1TqmDbKwJAkgq7M6f4XiY0EwYwFd6Wrf
84Yhnp4MkFB2Yu3xwTlyST6FVMxG3F25J+TP4E+GJ+qnpXyYy9nD71a8NlQhMHLY+qxWTfYcP6PT
pBYSBOSFKhK1/v+s03I6nX6WRow5e9om76I9+KtmrXyVAiCLK5dM2dCZhbT9/FWvbGCzMrl/JeYd
1IxV/UaWmThkQ8s2PD4csNSL5Yj5u+vuhwQiuIbZWWeZxOYQz7Gi068Ftjh5X3hvzj6U/dK5AaJB
hK0NM4nurTlSlHGk4zlGt/de+I7nfB4uL1EAwpWxQwV7uyMId/rmc7pmb+N2Gaun1vtxGu4vg6kE
el/FVrGcDJnCHbCRyCg35aFxhY6H8x9kKyHJL2WIHdx04PXJbNBtlhm1NRFIVGmT/9GvhJrj517H
9yCwDDIMs79j3sY7WsHMfQScuHjQ2bl/QgtwU134gtBxid6phsaLb3AGi46rl5ObV4TSJGwqj5Uz
7L7mHmN65OMPk1p4/YFTlW2IiCW9TPliUQ81xG9PXaFnitY+l2fYDVv7kbo77CMl+RPFTvhbDPUQ
1TF5OLnIDmxrMtk5vuXreJDLc+JLI5GXPvBRlEH2edb32xblK7P9Erf6o2rKpoErVx/ZHJ7JO9vn
/bAik5fZnMhXkO3u6KxlLJlcIsSxqeMFeNsIr5eRA5aW8T51x9hK0qGJbUh2Awx8dUIFqPWT8wZa
bSoG+ePMQFZJeXzSNXM99tV3iUYMzgK6HCk//p8Y24gtHDlZlBhuYxNVe5+ssn3jqXtkUuMiVVXA
L+tvS/16e57NCaLv3H+g5FitJp5eoB5DF9ANnWGIUFKl+JcLceLov4Yr7fERn2oOyTHLt8v6D3CQ
cUMC++EXs+Ej9k/ZqMfTYX7znSprHmPYVq7Cj41ZIPGtoC3/fTPhR2QGASYpDssMqsdL0LJv9Igl
+loG6DPqDXURdRt8O6nmdmKgbvnvYJdkoXO68Jkuc2utt/4L9C39L8Z7sne6035ldcotuAHG4V7R
/3DNRaKIATQYa001ehoA5w/8Uk3u9tZgpqSJZ8c7VFJjJZoz85PeUBZZE43F+U8T2QMaAVL4iLx2
9eVBf0RO0Bvh+y9fkeGWiE0B+CEOLB4tG6JN9hXrdHOT9u7UU8gmYNr3KSwstkig1qtJAz5hfPzv
eDqQDyckaYCTevsFmauMKfB0A/Y6X08XhsX2wZPrfr2bmYlwmR23pahECrma69DLmdEZzeklwklp
anqFKGkeeUOdCiR0mHCKENOA8SDkmR/oZD35/eBbtPgmCc3OngKb5RxL6jPqkT7p94WRv1gIYYIx
rX6g3Ysy5qMF+2to24OARfsBZMooBilQbPefGkNjduAjqwIdYRNF4CZ00Cd+0KbboCLwqEhO3sBK
jsx7GVZQWK8+itCSpLh/zsVPrHXw4K3+vXXV/i+Pq7stpjynLTQf5J98Vw/WRz2LKLSvzvn24NM7
ptZglUM9yomN7ON1ZmcYC269DIDSfuIwxUJIJIElPbKss9PoGuFwHRJQvN0lel69rm851/1ctr0q
44FlqzGOOnOn+eHWaFV8bXpgch2bF90ThJCTO1aevM6ruFTh63cOSyQgB3UGnsnbkJl8XjitxRKD
SYvZoIgWTfvVUxORhXlkE0fEXELAfhkMvO5F2yuIH5Qjh1wUEsYK2QHdKGguOR1DXlaIUM+AsEPt
zoXjqeGGKJRWMBVwW+zHHuHZuoBw2hHlaUMDd5muBu5ocT3KiQiZfNB/9NaMR+AA0dvQl7MMXPwG
zedG9BAhOg/DtRQrHw13xHP2mpPKCIdqntWv+kDLOa83t5mElx5iGTM3Cff5q99LF9UcIr3sXB34
kQr5qxYxq14plKY/UrX7HIRd98gcX4rQdNiCB6eYxtXknas3KzmW1EZrrnGVOcHdv1Q5CLicCw48
EDd/QZ2NSZO2JPnKrKOVQZP/T3c6krCCxeALnuApKPLH7gKp+BCBu7QQWfkjURINw4C1v6PYG5tH
uzTHYxoggfLl3TqvFtvmIlqzff0D0Qeo1ipcZLELOn0LGKYwOP7gc4yB7p4NigPyKq6M0Ype+lBu
1mHCdn/PkSYTXZIBWlSHi/3rl0yiicvQo0/mtIf2K3WSmMZBNZGseRelFWLwac01X74Lx3R6fE9F
qat8byIaDt6/d28zZTiCzn1Yk7IHZNNKbFS38MDAwK/im4TY0idCBNrmiwntm2gazX9l68ELfSw4
exCMVj1zvuk6bSto+65bzjpZh+FTDx8vO5Wx3nnf+pCnJCtfIF94fpzaAaA/AnAcIzr5jU67GvOn
r0ROu3DaLOVatuzT026m+RCT2vQTGMMelkArvcf6xk13LdnluBZYdG1WaMzrJnT9M6gfs+rq6jjp
agE4ZLLOtHMMzrKjXnrHj/3e95EHxRLgsPmI/vAOlijReJH8ilU4aS9YE4khQ1xRhtkvJKMJgRIZ
EumN8KFOihq82GKefiTm6hX2LJRtFcCVN+R4RvZDC0ywb1jg5++53NhP1wbttPnXCejvWTF5Y5ZI
8EmhbnGSFLSWyiUvTDfb5wFxxvGY//Y8mDN8L5DaNQ51bZg48XCLRK6BqoeWz3yJPCbXcNRGgEgn
jvObNjwbDHnwEdJpilEfLFLJANlWtBKwkB0gy1m8tFYArkzkMvYxiJ+rTSgIUmSGaNuQMpXb30AX
ePoKBPTNIGubDofhWdmakaRyPjpTD/syc62cgVNrOpfODsHgsMJZm/5CNMwiWNvZxE7knrqoFeVJ
QGeX3N06c/qS6VCxmuTUeZ043/ZWMWq/9WKfYWrd1inzdOgP+MkgWTGHcQLhEAUXY7pS0K0Rnicp
Or04xv/gQ99fmpMey2uEF92fqTZ8ComjqGLGCYcfEYYSxUR3tlVIUZq8/F99gO1xLp+tcd018tWZ
4dDnwv1MqMHlcS5YICVw+GEgWgxNTrC22vk60I02eJ659GtFwTo6z6x2JnSKk7HMnh6+KUX+pnx5
EwPeokfK1B0VmNE3lRMdxgfAm9Z/Tk/+AR2DVc+7Xa6GCM8hhrovofIVSy9jDzdpz6EG2gv0aZqF
LKYMJa5aFe7v718d+rGl5BylolqIyFPluHtnbakHgqKprCY69FVQ9zIj68mKbEIoFeQ7Nf4uZ4lm
8oBrncWy3VTfh6Nh4h6SKhnjERFTnInfVyQswGQ4mBrTxGxpqYpX6s+gIlFZiZmQIwAqAT6C4SzH
Ef32xByPx13oQF9DD0I9YfBzBmcZeRjMMhvTAPo1DeMct4FVGBfk+1oPsrsTnSSWmacrn8vQZAyr
CjTDvw1IEZFwuo3r1ICI0k9J+SFwh43HhwXoEsOX+p/uvVKE4T21BT+DznYQkoffq8L7N80ZxUho
5K9PjvnM3KjthFTxqmK0bVg3W8a55Q4i6AjOTLQ3wXQabX6t3oXnsiJdKAPAnWpOGdgB+8cbsiyu
bnR72iXMJeqVl6v+a7B2FJHvPF20e5tkbN6xzJzCqJIsgoT/hdH0mjQzUpgO1fC/9y/18InEDPsL
bDXVJZGAgIGfatqYhvULGuW1RgK2GaiB3MXM4EV2mVg/iDjmRSxoITrDj3824TtNh/7pRgWAxuLx
Eh33jdgUC5XfT6JrjMsBhmjkkYfKuuFeFFgJ/dI35uXG5Z9T6ta2KrVbNSBQM1Ub98CrolF80GVn
3594fen+FeexNCRxtOtBL2h/dKtYLZGF+BudT1o8IwTDEZj6xSMfREVHYC6QJmGQzWlJ/k0Sfjyb
QUJ12rQIyD6yecCLqOxGDJJDHuAuE8wtwHcgJvK5hb9kRZSSvERhV/Peb+wciTcP/Chl1sS+ygBP
LvbcQs5Qy5OtshTieow0nDG5koWW7fbhYvr9e8xqq6eFEQWT65L8Dgvsw/JDBbFD0ei5gIDrFeWl
sPiMamoKWP0LunIjC2S71fitUMEBvlmMM7asVs9w895DH0T8nh3rXfGaiad9ZKEX6A/tsPk02ay8
cJzyWzFyjaWzzAmBu6RLtH7KO4jyXHiR6IIgCagzXjxKvAas79kkWbd9Ibo1QXmflbs9cFhIYjCB
vCN54Dbt14xDQycnhT9CnxKWUO8o8Q/1zlDe0u0JkNj7VJibOSyqlhEDfCi90W3x2j41PbzQLfiG
YfAJigrINxR604aOZq4k08JoPoQ/Y77hgQGMrWCafN3nWhSdPkBiqFS6iD6KMEe7hf7nNFDJQaXk
upLhiMP5z78l45FuElddNUzI8ohC+60SVQvQ2RVumouRJaEAeWKzwvyys8ybHjmfsKBmYPoTjrkh
iYjXKrbdf528HBtKW8wDthwXMA3WDpUP7aCMyqvMtF9d+l2SugcQNuqGCmm+4An/eHnTwNNQwX9r
KOM8iq1NTkDQDemiQi6tXdl2by2EFA5PaPCOE7/9BVqS92ZfHqZEgJjF7lKnBtX/wfnL9Cy9M2rW
L7O+5K/ANwRZ69izOF+ysSFwK8qv4QMLMXvpfON2ZRgUUfodnkFejvSHaMG9Fx3KC3Ejbud1B8lm
szld5WCzzRrh1J50Qxn5vsO6k2wkbJ8l1zUIvZ+4zg8fmXWGu+vMGlUJCw9fkkOyUPecqh9mgqP5
ebbFRhKrzypnvQmtkgzw8jQEH1pw5wgkVbxYuKUPv2pnCRdrUtoJ8QCzlN8QVloVk+jRVi/rn0w9
fhVR/L/gd7tRLVnlM+X497bXiimphN4+u4WmgrS/ckjtuC1ONHVwScHPLW2JL3ntawsUF/QbkIVL
zMjtiMxOtWt5+lopohn66ue2OOd5z+LLfeo2RcFLlCbuGyiTjmdfApZmVKsgpimkoIYvBBZ8T29u
hUsc9Ce0J5Pe0S3arEPdtdPedJtiJPVHa5r+9etk+5pH4hl7AdHSSQrKL+PsPIVXJUj3zhoRP0Tq
iT5uX9NUZZ5+pDEtlsNeWQUMoKIZWkvGgrgrDli3pVboxsfRYrkcKKmrKTruum0XkKaeJ6A4d8AB
uGd3IBKXpjo8LuMgvU+RQZ/XfWOxHUQtgk+B1ETkYX5U8GThhPskMiMa/Jdr1bus7NQ9riYaTxTr
W5v98umIX9QWNowS/wwocJbTcqFclKhqftbacFx6HnlhqKnEQQtPFIGSxa/mgkngoZAMLXI6niFr
QrGoSLI4SMDhJrYhxARFKBf0HRqkgzORhtPnDjEogQ9Kplr1ZeZv+stIRuDtYbfUkbgwd+6e+yLR
hGUGGie9Y80qC8GFo0kqHj7UnNZ2x1F5iCWbnKj0sKSA0sFQB6nCW6pfOdMux4dWKNpFLV+2T9em
9iNGDIdRUA4zBjPD5tuMbxT3mkWYteRyId1oXDxvHpFlTnnZC44Z7tuOc2sm/d3rHBmAED+YQ5oN
IxT7H9trQcgpnIvYBsWqLwb29dv0dk9q4D260Egsjt9cmuwDiEXBf1jSFEAVVgGMfHxvbBiAJUaT
F+cbkg5Tvuc/EBGiY+x0WqDF5mpbHOow7EYWyfK2Gzm00ht6B9Sw+pV0zASjDoTOUfjHQ9JIwBCy
5aELB+CTpQaHvPq/JnSiocVwKAj9627xHcr91GSmVb/xJ5A7bAS9S4YE94BgJR7iUIQIqJoHhDQj
Lly7BJ2NUgAwG21KXcyViGJ79XIFgesDbJDpEst4ZWHFoTDFUsmjl0dZ9FuZ0BQk4vW7uTSbqg+0
/7cN8v/yxHCAeO0EIcT+rFUs+UsgOA9WB39R0C6S1EgUBq8E/VnqYk79+TxefRDf3GKY1pN0yWRv
UoUD5gl7ACMJr5fJJCzSkyPcaYRwQt7PT7aFJYw6JUXtGr4+drVrElBirpvgEMvbuTpQEveBUANP
bJqKOBPOqmG8+Ps1OATsIcUKSbNMJcx9MZo0imFAm1as0ieLXYURyKOaCxQvUiIZVq17agSwhGU0
isDkEofFYd93/cdRq9Cd2tWVAgAdsKd6Xc6dO1U3/h0geaIc9Q5dJx6TZGk7wwKjWmvyd0Z/3M9x
ZOsY1Z5WfvluRJSaC2s2fv0FuKXcvBWlAGG/I5A7Ie7RLRVVqmsxsXuPRK/AwUkSF+J80sZazox5
vYW5mt4mXqY0YSW+D8/d2qkDx1m7FvhXjb3jhhD2FSJ9mAjyZnSKTi+UaSyCyqDnK78S6/toHq3i
l4WEKNOg3ti3JMl8EJlWjoFKVsI3gqW4mo60fOFt4Jp3weAoRwqYace2peken8sun5C9uDm0ECJb
BmD+ZuHOKaJ5RMykwMDenk4MA5u3AAM7Ys7ZDDpx1GX+Zs8SF6eVU6qMG8A4bhb+73oxmLr/D+MW
dPkurdYdg02uPjn+SEFPxhk5/yLejZUfIrr5s2qENUab66QhhLS5GVG2lwR+ILmyBZZ/BHwbqzpI
g9D0yKAoKA9EYKVs1gD3a9alAd5MXLbycCZHvX5AJ49sTGILgp6kAc1rS+Mkdbz8ci7a9f6jfqX7
/b16ZXKnSLL4GovypQUCM3qxnF7mL8TPGa9hTKVZnaMdDMra3Orc4wYZVJd6rGHHIUBArz4WuFAl
3w5XxmwpiNZ7loCdUEEcG1oItnelpuYUYK1YyUCMFDE2tqV6DkAkI4y1fhbQ5EBnfYGU+MDlXxje
pBXdQbQKS3tQKsM8eoZV8Q7nCOZAoh0anjrUO+Yz6VwlVfUgt1b83TlSPO4ChwwDzn1lAnpdD0bO
fUXXKfaBNUqwgXYEE0Gs5H8S0x687U5sX5GeaV9z/iAV1G2BdG8XfK4t8T94ZlPdVrBnXUoCnrIp
uLAOr17d22LxNDIpn7ImdzrMP/JnGxrulTFXGJsWLI7VeQCKXS7Q/YkMFRGrSNVVoOKXbFRsgxbc
C94MieBL2GhZXNnUb9zRLX4otw124oMwGSYK24X28lKW6DhItLFPtAKFNlmdcvcDOJ5T6bNXdREO
aPOAs6akFjPDFggemGanXaR770FgJKHmXDPO/PRhHHcQPUMcC2tcIF71Xw/FvrVvNd+K2apMWTz9
8RUsLt8yEH8h3DjKwnGGMum9GK8QmU+APPPSktUYkRa6rqHbefTqnyQRJ1cZxf+M4OvdxN7f/gB+
522e42brRBuXFFmmBhmFTq+rroD6boc7iYkCr3FXHzYXjYRNy101QxADjGvLUpDARG57LsYVKObq
RmhrR8gs7rVUGnw8fgLG5UtdwHvKDEWzQheuHCtB32KAPObyQ/JcZ/o35lfu4xkPRKluute8YYEB
8AE2leJ9Vfwle10D2VwYxs5jlDlVNRHjGjCo72v1SHxqR+uo6JbRoiQDABhRPB2v4rn5ldpHUG7M
xn0KBH/CDCbGeYA6d0zyuhEe03zCmxRcKC26D/kj72SXv+p7bhjkU6AG3NyozJ/M9qomcFz5wmVd
c1BVk+x1SdXpHzvVpEdzGrhmvmT2JQO5b/rWG9vNAqvJOM8Jy8O7qyO5VcYSyjoskYcF2yfRPUAA
G+jxJ8DYqmz02a1oEP+m94YDlE/gMM1ULSXY0J5ts2M2MqEQBSDQm+HuUiblKUL233c48wCphkHZ
narakbMR77AX99MwFdc4LqSet1a7olovzGRYCBANbMxJNFb+INnUsVSNaKYu0rsObdeMatOuc+qu
AwnP8DSP7Pn+bxiLcQmyTronKlBj9fHiggGuxx3J41eGIrKnjTE1cSA4F2Qm8S+2+2AkXPvZw60e
QKaDuenSVyM2z1yZb3fQBzC23RaqSWzfD61KVIFgFTUX49RxaHqbRiwCpnEa1+axq2QfPetfC7I+
wV4xXvLgJQYbcC+fSu9rlrzyBUhVe9JxCWdD5khM25HNI0dxkeuVNjDADgV87dNFny0Vdw1Hzkum
1kTRSk6eouQH8AWEQEl2RDXhm+mOBnbjBZ7YGIVCTJHeXb0muDbVq4Th7TG2NT0vLyxSLRMmMmi2
L4f3hhh6UfpijUKJczlABiyaFC/ik8mp01QPPUopUHalf8nOBXyGAr+sYFRWLWKScsNYPyTKmdZh
jtLJ4JyrwW7uM4f4ukwGEYL+SjrkZXLkV5ZC5q0oqB66PQPkopVt8tNQI1UTL8UiPNo25olZuEVi
yWkcdK569MSjUoy3VhwiL22X+oV57mcNVvG/wJ2wSMfADal2o3kXKl7INgkm4NOX7xpFQpKIkCOw
owURGB/dyh/3YmGAUojDayKF6vR9KUfm0rcwwHNp9cRVlQBMWMuvL75Mxvdcrmh7WVosQLJbCKw4
S5Uqc5nFEN52K8NfGb4n9cg+raLBs3S2ppwt/AnKFz0E9HM5GG3CQnbC3ZubwqDTYo5VDShSTYv4
8EceLu59QEJfObPGX8WPkinhm6LpbZHU8iaRHeo7i7ln1dnflNpMYyxvNbQSIAibe9kCqN90mWG1
mRj30G8g6xK0nqs2dZG0I5Yh+lsoowAZ3KcUxMZwVKoLWMv1VrPaYuwlKu/6TmfLy4hlRM04VaPl
CXwC77DcSL4esR9wJ6Jn+23g08q4jtcSK6s8E0pgazAY90bRlhRHRrvfqzIRxjVaIuMQxl1Id+Ql
7tcNbIsotLasZOK564juMuSplY/zLCRHvrz5Z0Ob2g6R0S0thXQM22bPOWRoqVccrNWhaQfwmEhv
O+Rd5mOyffFYqHaOxbf04jdPUKBzVP9+LBdJVhMfqhj+qH7cKd0OMzuSsmeO1Xn/L0lpeNZDVv/K
xI/oOlKtBicqFrUCqmdCrQrglXXZ5gBgg4+cxbdr4G8IUjLWQIzJAwxQDweXJ7KGbsGeXfzExT/V
mDQ0butPiG7ZZlea4vVkKSH/gbgwPAFF6ouVzz1tNEclxYFHPQgL4Hvq1X9JjrgWt4DxrRKiNFqz
LyjScvTx9/PDxMi7r6bL4meZm53kUouaOlVreezdxmJOxT9IVKK6Jk8q+K6nv6aNbcLDIugImA8D
5hrhI9Ialqye64HZD4rQVgbdF7r4mN+4qmrrnHpaUO+jhtFKoyo4HMHH0+K29gRaIFjG2QIY2HKm
I4O2U8H+8dHNhF1HkENa0gpfRYF4lByvHuRRA7/tnWh7Fom6tfjiyE6LBqaiOh42WyXYDg7DUZFb
paVPKa+gB3JdeG5qwlBszjlxv91RmtXNAihSuoNtNAjnHSy5oyug1wux6dD8rsTzA4ywn6lyN2m4
AC4U+MZDa8HU0xs7SbSYEWtGiaplGPF3CvpGwNzkcQRlobj/dnhUmEtw/A6LqpbYlHi/+eAt6lZg
sVCN8mxNqajDM2iCXvXNGIdlFZlAA4pJC7mxdXafifhJ2PEFzcQwOJkGXo4AGVE7QJXrP4uAF7b8
OVOpazyJvfJm3nDXzgASHI71zMk8D53q4UgMn5LUXjMot1pqYEMTX82Zl/UjQa4VNwaZX6ZMwkZm
VOLDpQfnP1CJXSDJB40B52ylF+HWCyZKASiFR6seJ9DVxZBhLZk5znh8zXYjm4+xVPfa9Ss4wdUV
J0Csq6v1l9BvfCIjXwGqSyNV+HL0SpIMazcBtsj26WYOwZ1URqFuhh+LvlGV9OF94xxGxHt2NcXe
EX6xyBSSZ5xUjxoDDekChKKY4CdZNbotB8zl5Qbu2YIQInNDc7zoUC20ob7CoUkJTcPR69WSWAOh
4/46G1m3Oci27oFB6G94wWg0MrJXu31tihd/WOXLQ4SfDR43CWWq+UpeAJwGzPVLPvB2mWXnV1VY
6nMphXgJCD54rVsBjRIkaTIAoh9bPgKM62cixaRuFHUZbwXfs9xx5qeQsGppsQEnYrJndcGqdcpQ
5Q06Uw7zElvtw8ixfd1mZRDwB1gdOKBWUv3HEZcSMOHzgrUsUzsFZXT3EuU6NjgNwDWCs9dIW6VA
boMl2NMrUyIu6v+3QoJB60ozJVBu8SFYl/T2k9t5fWKb203L3WwfIw0RyZz07QcCZkv+ZEW0eijK
TA7NRz6ypl4Iy0YfvrIyLukdPuNVhJ1IVGUMN5livTpIXLOU35BwI8WcsYRyK/bwMzCbwKrRHmdl
ZSNVa4aRJLT7XQ57JOQBuCH0exWVF6nWUsJDNhgXSJ5vZzl9CKmE3Dtc73gPcE7LKO5hmnbj2TfW
o/cXOgiey+9MqFLqALmHWbXTKUzO5x+rXWpdsRd3EdHSL7irIWJJrNkO3E1ajs6wgTN++Dduns3d
oPMcjd0PXVyZ+1bi27AULZhOYoAKxGy8IkLBWmXjCYZbW7IHBQCRR9hRcoH0ExwUJ0P3o1epvISF
AKCHgczhEIzOFOO4CiZ8RJb6t/W7mGl3kiumYsU9TM96ZBj/xDY/ZahQ43d3tHiDwPZ2gqmamRF7
0qC2UHZDwEdOBywFKZOq/7cwWARREAwoYtS3TBQptHm49/wu1BOtsvEfZHmiD2BdOzMScRn7XLQL
Bwpw+Euft9GbPh89Fo7vUJ7F5M0AMDnRwIGlzuqbmFMlHzbBw3EgpnhOiInLcPbemfdxNhWxSxRi
LAxIJJsSC2EKvmHTfO/uhJYUdcP0xvFk4VNZrOp/lgjEEBJyveaV02giJV98qM2oG1MsR0HkOPhM
bJjXlGkcQ3O1+T09a3c+jhmCRmG1TRj5z6B+jxBIemvx7asRwuZpYe0HpaeEZl2L/HQfQt+tkhLC
JsXAq3UJkVJsnrH2mv/UNkiILiU+FK98LvOnsW1s1TmGpHoR5vUD5rYQq+oorDVm0K3m5K+cPcQv
B/rpgb0qgyLZofZoaJLsAAYTuw+9+t+PyXjiwbtpKNdfHxEjJ6R0OiiSD+4psNRFNfzEU+OoyOAE
iLGHKVnPZihg18Q3ZvWGiVAmuIM8zjXZsd+K5XqLeX27Ol7cFMKzNAssW/w4eQ6X07moVgyoN1MN
mdqcg/UH9M05OB5/XWF3kpcVgikzI+7HqQZFUOVel9sNSbUB6I7eRLBu8oN26JwT5c+s5BrI6RJo
Jy0/DUQ9M/Lnl/7pe/khCdi33/7BtrrnrOsJ3rMLhFAtDsf5xBZ2pDIhipysEGWfXT6lyXEc/66p
loY9Kd75FJ3pyLPV25vxeWJ4s7ewj7chhsFBy2MKg6QTQf/c30B3l8kIdy/AW7jr8MwfgSTZhyUI
PMi/i3Q9CLKWBMYnjoiSJDX+lmMfW0S589KKnf9/ryt6xbVAJe11OuC/2lfw7LOT/31k+jbVCL5c
W4dokXJZHZHTgdLLn8bxEulYPcNzQ88NpG/aCNZn+f0nP0Y/rEmzt7yk9IOR4ZizCONlvmRJWZdM
N0HzdorJFLr7eGK15lTi+Wt6e6/xIxFpXx6UiG8nuovQeIW0S2X9z1y0CRgm/zvFq1HjM7GM8gU1
bayBVCpDsn8U6Dis9NSY1/VcoVSdMMrwqb3sGsnHDgYAeHymBGKPv/ltr5ps8yRNlEwAWkHDyQ9b
dhLrfOE7qK8dldvbw5jmgCH5IOzjFOwMa2ZmsLFxyNKn4j25oe2rxNltNH3qX2jy3uTMthIflAK5
vbqBhFB/hw2mmQ3thmv2WwVK7tH+5EEHH1uQhSAS3J7h+ZUZ39hrv9cycAUlrD2Xqs26v73R55ok
Vb7+YwSmtIcDjpaRSJHIfcqWXz4Gg7Vx5uc2LiHUZwvjjF6cwXKyCtgDISeZ3Sq8m5W9zj8hNo/Y
wxkBq7pmdX0STpjQZZS9wDXuLXzNqzR9UHLZUlxnqV7eLndXZoDKDNt6MIeK7M4gj3ojyiHRc1o6
uUt5wnpCj9CFIyyDMK91zPRJ5lFE6YJIqS0VwCDlZCam5zyJnzZ78dcazUhiCfKdN2uoFdqtNwJb
rZCfbZm1vxHXyCKbhs06XDEnkhlsyVn6QoZ4X7OqcawHqFcdraDYU2e5V2WPfKG//NKV6qGMF6r2
jCpGctDTpZzxUgOHE+AXAuZ0liMv2wMNIYT2fCwyd2HqbFLNhHWpSBFCTASrj5ugu8GXk5KyH3Nu
D9H4UFs2Q64FaeBke4/DqHn6ye91om2LXFgJ2siJ1zLHDsL2jqfIevAPczsw1BV/DtKmhr4It4Wz
LqKBB1JiKmelC3jey0UVf/ABV3aL+QYCgSfdlQUL7KF2aFvncxiA6zMKJv1nU1VSfQ+a2LvN0gRL
5CFkImfXWgIaKyy52RnS952L/qOKw2unCx7FRYBXzEhZxgkMwX8K8FOx4jvWTXxTtyRgUvF8lgVG
ejLndg0Nu8A6XlLHPL//8+G6Y5UsjJ+er1FrgNGgeViXKCiiVsUA20UW0AobxmXTSurTdUWOu6Um
l6fpemR95hl4GH2iFjjtHeMijoiZ4gPhzVk1UUj4s/+mWkZ4XQM12usBPC7ohWcsx8lrtFThOyqQ
JvuS2Xl0R3/3txwFsgPjMyKPkQpGyMXOa5pwxZj3undzPpG1bVXWNd4D6asAlBSDYnKmqnkJHNls
50JJQ/Yo3jpf4UKQ1PHUIJJPWgIbGkLCzMtNHaizMv2rCIsc0xiD8SG/+HbBJctUCWK+dN+1c2xb
yddFfUqZJyfJaHE8psTqpO2980Gys6eGSuzhpXRapjeG9mcFp4kkFi5KJPsaxSKGgBeEO5zXHzVV
2sDarcoSlwc1/pgtVTFzDgStDDNptnJsfvYS385KGtJeR/R/mhYqK1tXF+8KyreqLmFHWcrVZZ8B
sx3xrZ+e064jWcyAcaYr4bf2dEeViLqQFBd0GfYnz5OcjJt5MkeRV7esdHLSAcBFsKn5KVQ9IWQo
kMklbVGPdNa8NwsJq1x1KoUDKbM1y6l5ZeJoySfxu4IsYxI/J2w9DlygA4U+wyLMVEZbNDEqJ2Fb
FLumdvq74CqW/bZkeeOJ9QHNHzX8rygHM2BdmQX9U89ZuKzCcVuROXy9l/CSx+lUsQpVPWr027oi
plnuoklKH75OriIthC35A2+G3t7SOR9jD5gycvW5gpj/9YfTsi6whZYnE0UpledFIzwkBearPPmF
guHWQrEJupVbZ5ZqQ9XuHSFAms2IwdTmOCQNVOJZ86ovVMLGxjRC2qCtgafS1yePgJ6KkBvahCBx
78zAEesvbVAgs6R+XHWjaQVj+GE02HZn7nGbgn2LQd/Pi5TDxa2Jq2SexZP2QRSdspiJdkvRcy6I
MW0apP0TXyl9fXSyTHNotXbpY3COT46jzRBar/JKq1h/e4kNHNGJATOXIOEYhhXHS1hdsBzE/fJa
be+LBcdsb1AMaZkjrfIQ9UstSqCMaOcCN/Ho/MpgnX0WgNBbi8YLV4ORiaj/BV8Sh2lNo1kOcTYb
qbof8YZDxRgzI3oxufyOAgLN7j2J5mTmorLTA7Rsk7YFkcwgSx+IhY33OHkMI/S1Tj5QnZ5W01Um
AHi/tv/fhvXkFBEGSVfgOuZ/FuZeQMIdt6rlchOPUZzkbMVJentcjmUMJozlpmNanDPXotL9zvRE
rVeXHR5ddKBpwqVQJ4a8KptI9+bQ4FiSddNZkJufMCmLoVJb7eXQnMAGfr8VXiXIvK6onN5RdCVY
ZOS8rMrnaPHTnWTWddHJ5MpEIYBaUQNiVLuyCiG2AfqOb4zgn0f382YaOrN133pMPc6i6xAih+ls
xBR2/uAqRE8m4HrC0RqFhA+A+ZI/X3root8QC2jW3KiBHiYNhTxe7l2th2MwomLQJXqGguA1mC9r
OsUIXWtPSacm9VgPzaPne2lENsJG0GmrEmyHNNGE833gcVu4l9QnimJ25PWq3HYgdsu1f3FIeeFn
mMQDsWULAu76bHyPzG3aqn9TTOoGJlPVJk40aEbX5R6RjBI1T4bPn2FHucZyeJGX84fGMzSdh56o
KZTPNiEqJd8MeG4ARozgiXzSE7PT0sN82WyLCViAqesp2eAAt18/zVleYz8pZY5QgAo5CtwzRdkI
Ud51OemzoKb5on/8dvmhQRa33cRSCjd1owKEccHCKGgMg2+B6Y/3vnOaPJFQtx89CfEVvyhnb6ZS
hDJgpK149yEJ6gp+7u3Qf1cYfeG0KOT7AZDIBNVCcngMz++Rbtd+eum9KaWhzpNTqnl+pHjS28Eq
ctIQMNR+6TzSrSbdmh0Sy7ezYcNchVUOEBjmuDkqz0jZeV94MYO8wztpxyX48tp2TTFCaM02835P
rWPI3WmESHVK+JCKf6Cniy2Df3L8qC6XvjylK5xAN2iYnxZMBgb3a+STw3kj1ZlTdaMC4MubHeGG
K+pgU8fh4EIeXNLOyrk5g/1IyAeWvc/z4WKYi7wlGaODyrKVjSPJYD2bmWcc8Y1IVWYGCZPRqKb+
YVVRoWHhdBBoLz0Ek61RXJpvlLEcbo9qEZFHgokRdij3fADeLOGST1DQfuOsTDF0b7dLIOpznTF3
9ftbMYVguKTIIGq44OhlXGkqdTkEgHPiMRG3Ew2HqXUvU3GO3UItmAl4ZcA7J1RWorVKgB2qwhxn
/gdjXONLNka4O5sZKYrKBsZJTIOPFetca7ri4D/5BcDDRoXht94y7VTp4LEHJhEGV+vQm98sh2iI
eSy9szKBDNPlHtlKQO0dCUgd/nhgdbmboDEkRXdfr39w14weESAsaZB3opEecoVCy2MlQnkXyU2t
ArQxT6Rca5LjKsTdhaIXVw/OW7F/nk+MC6LPJHKzJYa4tpEx2juAsu1TnIKAk78PR9XsuLnotJYP
a+mGbkoMwYXAcWUXIMmln/dhri+jJnuRgN91O4kK7iknXZNIVZch2A8DLvYCYyDM0jHb8g5tMxs0
V4i6HjYJDGUpRmGFQ8bwzx3KjyjdiBywoC3OSeb1y5FLVDcP7mha+2S50awHXzrYqVUPRGH+YBLB
/gkto6uhddIJVx/2SAVF0YkdhP13ozrNX3JpzewIgVUFEMV7oDgzKv3DK9eXNnebpqHUhslSnLgW
wRd6qPrhjQvb7Xga4q9cDwyvpzhIk/+OK7FU4SSA5AsnGynhhkDDk3bOXw6v234nNs7KQPwdsPlh
twFUZ3/k4zcUnQfc2ZN3ozDx8v9RqxE0ABCBllBIcA4cXRmNZDeMOKCQYCNJ0ObXswJKbLFj8pD/
I94OHI8i3QyrGvHEAtVBrvxYbGzCzJaYfPXfM26ReG/pjy1S8yftjoqAVl/ynw7eyrQ5y+xcSAKz
QDPSFCScZGYK16JaHBFVjHa6T2JOx5nWW/GJwNQX62Pizq6l9Au1J296tNBOfeS4BTQEdAPGw0PX
gyJRSasYcknpnJ9qJ53MLHOq80dyx8RxYs6vjhQnmUs/uy+7MoubA5YltJdeBMZJNbJztMZwfRhv
VrtK81GGy7ogkB/9aMe69OaJiP+JvkHEuEeCHfxt3lX9laJWabZaw27Lg0lo22T+1RSoEqQTyrtf
Rrpop9qoJ7VGzLpzbjIO+4GQEJWCcrj8FNBCBH6g5AfTJmw9NjUM20sP1sFrXP8znL0g7BcCHwy4
HfuFqbYK4h9XwAMKYzaixbg8mOjTLUQhCdcr6M4xgI/XqeXUpAg0dw/Sbe6vcGaMoIEjeB0xfg4I
zCoQ1QGULVfTDl/c21jhaJ45wg+OAoQpUdSH2AwxUbGquzrpQliHgSG5gkTufhTo3JSHLP6DY17P
zDX76gzCq3gnnge9EJXQJ5HaL0a8ud/reX7KRi+DHupxosgRu74G+i1uKtuyvW/abQB883bTDRrV
8CLyioRhrrsl/orfkdXbj8wboasH9ayGlXnqslXh2NApu7JQE0ueanye+LVybRObsH2YIajeZJua
NfFBHiI9/fg+XrvvtXQI1GHDL/rEVnL4L8ytFDXqFeqmVn2Tf/NyHieRjGx4kmP+j/cE7sfRpeMg
KI19JjetxJeWOyze3IL2RAwDWS+rbPVwpvdvTDU5URHwIpE98kh3LVrjKK1+gLARhDrdjkxn6TR6
Yq6Pq++cC/NhgHfEhdWTPG5YBcFW1eOZ0KfSM4qJdApZFbWIBQ3j6X7y7A2vk3KKtJeA2tcO10im
4sV8kIOYMorlJGvec0pr5kJpBfGt0fuzDTYt0nPRJsJ5KQyjeX6Hdi8Si2Wolyr42igW8LrhzUvk
8DQA9hcAlLqEtfZdHEQzFgzHd432fjZlHlF2zhy/kZEVeQn9Wv1ODH/dI1D9HW0VNYNNNE29TDsZ
JOzwvFZrpTnGbBO24c1uwAWITzLm+5TmxVMQBlQxvef0/8ZZjPzSCpXW9g3BkkzMxbzIy4KnBTAT
5xQ0M1km44w86DrDTEfHIyE9KI16KLl1oRO6tjRuJjUmA6g6iNOExtXG6puhPDW6cg+sSLBYqxJT
l8vCvP3ElADcUWtTSFL1kICqii+ZODPCu8ungr4RUkXOak0RD7MLltQpCbXo/QXzusnMSyxrmdNx
nleGFcHdRd+8XcvS0C1liQyVfHL5NlFgnoWnI7sLqfslWv1emr5HD/1K1iPCyKCLzwBZqvNqzO+J
EFOYX2aTlp4SS2Io79f72TjbxlMsUmbubU19wbbrMuRat+ZVuLmLYEkq9/5dHqXp00YOTkhpAOKN
Ia33DGnLJBya/i9LQGDM/AEQ/MBjPexWayDVV6W9fU0DGZh9c1IpIssGD8oj1lYWBInrdyW1tZ93
UiIA9LEYa6IEfHGrfq8ypgvfhxtL65mtd5zvbKH992ei1fr3Ga4KIK1giyrKfm6JxHsfhUFWG2Es
xRD/mMdF4NWhcaFzdad3tPXbhWgOopArBxCd3K55PXQCQFX/ypQcqDSR6qlqf8gWmpyvPfVg5qRq
cZ+NC05LW8lEWpsHZu4/rjFeAnPnNUqUje6z6P+iDjtg3AvHbl2yQ1DjNjmi7zkuE8nkDRndbrFV
s6WjH0areg/A61W9nReNkqirmEX0ighILB9O353crqZn59gPJ46OlhSAD49qwc2R3+JEvKDuM1d8
Z+djaOvwx+peSwUDePnEWi3iOKYzosIb3IHEil57Wdp60D4ADOUnAyT0aFP5rEgxiHUR5DT/IA8K
2uttnbxuecjXMvi/xTzlZxr+QHFvmkp3jJQULweRFM7PKbEuELjp5IoycAaWeWVLHg/PvDjxY0KQ
zwrGfKpx2lg+8qrT7QGlFWfWS9Ram5pzoJqfKYN1VUt8Jobj3O5EUHfIRRHKR3Op2M74zqqx4/R2
PRzFjdeTS4iIVu5yoA7ZNu8o0/fVnx+b2wmK3UGDcj8cRmeFHUTmVg4DjX7hSw6lmw9tWT+CJLMG
lF6pIXwIxN2aZ6lYywRrR/zJR4nDCbhkiICBiFCYRSRbzzfp6k7wEW6jk2GknZ3CnRM2HhDVsLNX
NJe1SgttaqKlz8VJCN8JLePd/M29eQUwdKZiyWLHG49UdOWW32U+LUMPiZ6Ggkw2nMwOMvy1BNSA
ptUTBPOUR1lj/rege8gi/nuD9UVluD5+u7N6m9M02V/GrjTl/XZ8E3b0dLnXQ6Cvr7VVQJahRKv1
8Te3R3CJGs94X3n9dXe5EB8pYzrkg2EBs3ypTtJdbwaQj9F/B7MMcczTWjQu088pjaIwb5sW5Fgk
IgyzRjrg+uJ7swfj/pcjyOkd81KvVTumyMfxeI8w9gAK73hlXrYDlgJdJMTBqbmBj4Jtez9HEqxF
247RL2dyzbmk23EF2mpqMJH5TwJh5MOTnq9Kby7q3OZlMNsNkCuEhRJkU6X6yQaE0yd/+GcmOO+E
4FgrKbiO9s1cmtbtYPkuscUuIh221AaAFgHNWl2vGHtgmA4WcOE/KUY17eTcgbBNrg40wzwPVd5n
RlaNW7W7AykkrvI813bHEXODcf6oBQvfN2aZCajzb4DWcxA6p58uYMHupmmixW3FxiZ2sSVVf9Tw
QjwD/VpxZJ+h9n39tkLcELkuoYvQ//lIT1snUXK2vhEsmAnigkz7ivQQj5944wn4DDmS9oov1EUb
ZgvaT29Iy9Ld3i+oYjJKsrsIYBJCNePIt2NShyAdgablY14L2rpFB9/xaIDB+bdQ931qBmLTzwff
aACxYZFhlT45ayyrWFXokQhgNKa750nnsmNbRlbzktfqyOg4LTzTfRTcefSHmaU2uEPDx/7iiD9A
oYe8KtqUAWF6QzG6sni+OzZ5hVxthGCRKedZuxfvmnMSm1P4W0ETQfJSaV+ZAwhyeLYB9ehWgisW
lukH2TTPg0vOuWwRdMiMS5lO51xJxeLt8+nOJoMoiCR/Bnou88q3PHxqaeouJtPB3dVuZ/7vW8l/
vXHLDDLe9Me0C5zD0RalTAyrkgmY35sfzkbW6lRPdsFvgwHKOgmueYUs2KD207f8RtErM1ZNQpwJ
R5puvTbl3iAlV43m4svHUOye5ZbnJLMPbxxiOSSXUK6iThrDUnOWgf+VfXBXwylutCbMxYZVgCNe
OqVIOj9ZhugLV/nMoHsj6Mts5fPw+DLdzIore3Rn6h1cPitwYsGHLt5So/Fz/76PfGYfNn7UElzT
aAO++LClNutySiR26Rh3dP8hmc5w8YBF2Iv7xEcyzx2QgyyMYRIpBhSSC0JjTuNFNCALhja4ZDGM
2q5EaCy3TzaKwoSZvbo8YT8f6ATjMMwcbxBCqusjzk8/5EhuY30XcZnTj45/FvetjCHT3WuhXCXB
NHPHCp5K80+Y5QrkoPu+BwCpTN1F0mlSTav6ujUbPVRG7mVgzvwQz8c7tWwSUzWntK1nsiCKEoB6
ILnJuelEj5hMvXCJRi98dhA4XePR92jotmbdExEifANsaoqzGsRmwi6OsH1waY9wlBzzd6SbvwU5
QO12zwhnFPLvznw0SZZmQtAB6Wqdl6QxjEbqVdSp5pL/IV3zM4tdqShL+6Sq2pcQCJrRLf3OhGbu
q9RQJSTaTZU/bbYZJOuo7JvJSYghBim8xmuAuTWO34Ny8ezV2TTBCNekY3fYI2n2CQr8YKzTT+BS
mQeAZratvOM6eONSrFBbZynikpIeb+wJuGIQXaW4c7Csom8vJS5b1PSE+udSNUSfMWqsV6UO/mRS
JaZ1hrV+a4PS4cyYuDqkZhDV7nwRadNYGmoUYp1S7YbSBcLWguEgX9EezsKj9cSp5N95zFx+YsRX
xlaxlQI4jGxEY97bz+isrdkJ+Y+1BorxeDPkfTCv9zR8+uGq7kpSX7R8pdzoqNrUIdnuv1krC6cG
kfjLXsYi14t7ZBQBhTFxK1DwHFYpwLvBo3t2PeriRPTSi0g8ubif7+f/1hPCrojhSxZSHrIlLwCP
TC+4KkXDWJH1Pnx3lKKoLyxsZxdtuSBSEJFByxzaQN153LCKwu57tBcdw+SDe4GvUWuVZ5JzdsRd
JQXlBAflTZdNG1tLehtx7o1bbBjAm61YMazxTGY2saTpjhB9RkzB9ivjxaYJbn9GYaMEyuOlCgxk
viwltq9o62FO/cRYBEVxUDsCwVKiSs44fbI3tNmGyhcjklj9EBdWI2/XY1iFhkjIytjTDvGw3V71
hlSRNaknQsr73NLlu/L4A80l+e5b169ErHrUun3SvnKdAb+qOYwnrQzN3KgnfM4Z+P/RbsjeIvZC
RkHfcKlXABcOuaDKjhaOwQCQKQbCW0Yc/A2Ve48XLUk9N7GKDmSngscw+BnjmryJJ5jdbj9x14kr
IBLsufvi3EZ72lGLvwTPP+z8IbLMwOFofL/XNoWvnn0xTeuBeH+BzOO0LhhGtpx5Y7e3SL00Y1EL
T7xF8jLSEMQYCVVwv/c1hRqB7MkAz0z5+n6dok3lN7nWOCLHYyAGe8KDmWUb606+W0YrHCN1foVv
6Wqsd6J/nPs4+uZwWs+HpLIuKH7VRo+Q3ch3LCaXEOveoRsg64gziRwol7B+KHB5OUImHIru8ASo
S+dDNMvdRDlpl7arHeDpJXjRUrtkSRWBV+JmnbI4rxvwrfFMBp51gmMWgG6UdJoh/KU8RPxATdKn
s5Bl88sP9UukxJvZJtGl5ro+KLyx34qNO+lVKdGlVxaLLTrUIPLdvm9zIbOEyKgx9fWVN1rfDHzT
s7d0ZPaA0rJnatwtLbAlGpl+PrSzjLk2sbNzpsdrszWWT6VJhNugqJX6yG6aSaQLke3GBKhdbDjw
RNrvbMLAGikEuPfjutrSLKOp3mXVjqoSErQq2P0JtZzF0Vjr7A62zLYTEL2+t9ltz8jnhGBFxa/6
/NalpQFEazNf8J1LFOBi8QeKlhgMTE+UhISFaHQJEq5GfkArrWU9Z2N+/N0rwZK9mJ61PQyxvD2B
ob0AThV6ZgDZRy2M3KreoGRURMnSSyKJRFT61jz4co6ZdlKmTyCJqZFQ74EgzC3OeeGdIAKfqAzW
GHgjpPRMozktm0ktnPwxIOO0LEtF+9hOgXnC0VhSyns4ER1JZ3GHja56Lu7cXmtmpN6Dffc+8Src
IGjc5t09cu0ft6mHqYe+NF13GpURKM03rZjev3KX57AHo0p1JPYHS4XK3vqJoepJ7vnFfHUBmYl9
Mql3eOgvXbLjewvSZKumia4DpHlkBUNvmuX2sKNLJgOq2dl50E/yWOfrGpPRLzRvTMAu1azekPN8
QY7D2E1iGTOZoUTaLpk9lW+3ZXZnmM0WpLtehgnAcKAd0bph8j8in2ex3kfkLuwPnWPJHoh6dXH3
v00Y8w2GzMvtfEMtb4d6sfFqOjfuNw85q0s4gFPHVFOj1Lvx32UtfddGYRkb+te5T45k5L5DRhT/
MKPYvDHGytxQqcC3pyBsN1JC7lSBG4Jk1b6JslhO3Nh8bQKvGcyHxqFJENHzB0mBQclNahkVhmt8
wQQMkM1vlq7qPTWRvksT+/wtfzX9H1SWfnQKgTc1GA5anERrAbOcwMpUWHBd1Kiww96sRNKviiGD
FBnUG98Z7PRy/gg3jj2AFturzYiSFQ17l+45f3yq+Cy9eMEtDpo3NrS/xdH4oUaTCGABEbA1yHso
Sk/413HG8sb+keL42cPvOAU2a04s+OaHG6CB59S/IR9BgGP+6OKzQGTXb8LfnSjuj9xApagRqMlh
HN9zXOmaR8QtoU1G7XWJ3CL0nkW+QcqjCOQCB4FoI0R6zZOsUYHmtSSe83lUSnkWUi6DuhF+vMDA
dDOStwBa3/g+ga+xyU9sph1aK9OtojxxHJwVWOlUInheHT6VgRUO9LTRkzLD++ndRYxsYVMjOEv3
xlguXyYIZPCtP6EqwARxlq2va2tv58cxCFKpMa8+obnQG3z5D0YAvR++jT6gy6fEc3sKZ2yki3n/
DFY1coyOQQALYLzCdi6xo9UUlcTWKf7Xp6rjvXnEQoqm5V3GkASz2/JaZeUH9WKQF7SnGKdNVYIg
n9muNS1Ngx3Yi64dxn7qQO+dfj78FTgtoD+fk5ocQAa8EtfIw1kVOjrJzu6aXU+8k0tThr1kADzU
tSWfK1xugXUbWuIusDvgA2U1Rr+B/G0TIyDbrfKK6xWZtXAUrJIcwhoxluKNQOUjmXr+aW9HRzwk
I4XxVQgdI+PzT0fkAnvHG85hU0L1UYXTxWjGb9qXy0IxS4rtR742ARvlOCBxOc/42xO4mqLcCF0C
tYb+34E03kYfnz9Cv5A0uP3tIyQIsn3VJxxAF/zUAdmX6W7r3HR/mr4WB3TmlngHF/VfPPtn+bV4
CIMpq8ytjLwJsUURN3BDZ7nAg73fHWuq48+6XV306YqtED19K7UOYFz/tk3MFZafmEn5H/K0AWSa
8Oejm9SEXx1X0/wCcEE2buO2nGIuj7X39+DDn4OzWFkkwxbW28Z5n+ktPgC8krBfD5U9wftpXxnX
W34QDaj+dBoG6PQ8Z89Bc+V7XMWhSjyEH6RcgAYKZ4thg+eTjBkiXbWiY4ZXNl0abstZVMC1CxZD
H/LuE7O2Bj2eBvZLIuArI+fvoXoyorVcSWAR92SfTx+8xjwDeCfatrMrBS1XfiPlKkdAvsPk0Qke
hb0p0g2Dm0UsbR/fvoG9iLk2dcFMl7nur5Mqd3yP6q/bQB5dTe8SCNwbOreOxbNXI4IsD+Ca1UDh
YpAi8CR8cWzZU9YEqnxa+nTxwn0Y2Y8mub7OoRBikrirWx2/UtEsAR2nvAKHPHuvY7goENxSf4iy
zNQ3zt0x6274c5/TEtTFBfd3a+mhq4rRoJ6+wi/FbGG3ZzKNV5m9unfzvX6vMGpeHr0gYLf1rG6R
3tyT9j8LHGlCHLvD+mnw5BBWOy/ehbjxgpZeRiyZlGt+82fb3esbVQsAoaXjh9ANi4mwNe1vB1Jz
Shg0lw2reD4uqye8CUTCdhkzorwFLv4X4AQqAvAPJ5n4DkKUKG8VCybBVcqCbhFqL/s8V/aokE9V
RtFFjd8Oi2oA9ov8wf/aKS0V+r9+tHN8JcmQrRR9bIuy5T95ECwgYGReNL7O8Mir9VmI0cHn7+3D
5H65O8BoiFr+4qHlESgsx2tnAP+UDwYJMc5LKQa4v6GVP5xpWnBFPRVm9oUm/kK2seVtfojmV5wU
6QwDQGA5RwLNzmqzH5V7IQRz/MZ7mnLO95oGDvgd2znLIlpx6ZrZDQjvOIQcz7dRJASE15WrKzea
VdJB+4wxu5QmKQShwLntC1CG7XBLDGukQau1Rw2OzHUl/QAMtE3OOTWcfj9Bo2Uh2rIyScNcBoPx
8ZEp5XvM9V6jIKNipomJ9hpxgstl5C+2Rrf9ebc6ZetEtzGAR3QOgbdsTsTtbEcxf7q8Gaw62ILF
UXxVSHHmNndyCa05UWl3cbq1+JcfmegYfs7RRiQ5CpvtdaQqESfXWrQUIr+lia/ogbdOiwcyMNk9
pJ4O7DjMzP7p9cUECrofZM+TlipFN4et3Ve5lhS4rKqduRx29Goem9/JneqPI5OoKsgRDhDnzXz2
9Rr71DbT7LkSLcVGB1oNYYm3+xy91GIhSgq1lqORAvag4VOrdq50wL4kthHNp7Tk8fkXPBh1NtW6
3PljXfKKLrxDGWo4sY9CMM7LRNzpRUIg5ckYjHjdn2suHv+96r5xTgLaL/RRI+dTTch80MB8pivZ
dYx40+v6QqbxeEsovt/D9UiBPF3qJy6TDY11MMouBrWO5QhCFWOJSO0yVBNtibguqFXDGrRDwzC5
m17A9Vm8UU6EAuJ4uh9Ks6Bmmue2MSr2SAZXA0XywBG2TycI51BnrEGaK3JZ6xPrWeD5kA7UZ02c
6QRgRMzaVRKU9+/c/sQWTfzzsvom+KOec+PHCq+KDX79hVD0VVb25hbhLBcdkZ+sNy+YeqBFisiu
mByEmJtz+URgN74e8mQMsgWDxnluHjxu9WRxmQ6KttFNhag8jQQw5Zg7ywMob7pfYGhXb6DjByzv
QYjUMjLZgIbH9bh1mnqI4E+zc/J0loMumMU0SHocfRHW/76EyU1mX5I1hPxjzDpiAVY+M1Kk0tGT
AE+8bBW2oX6FolIscXM8BheRlErZwCXY36CGpf1yJiO/gP05Dai3+Cl9CjlyMsJb70NzGqlaQqJU
Vags8KjUzCjkRmvrNxi5aT+dhClQlbRC9chIb0GPJKpRbmolL29C3GR7qU+wpHAHsaa1Iqakyr+m
IEQ//yFrXkeimbAjZzIu+DwpkJWn7c5WHiCkJbxT7maDSJv92RQilA==
`protect end_protected

