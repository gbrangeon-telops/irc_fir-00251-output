

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
GuWEw077quLd3kfu8DABFf0P+6oHLq5R3U5znEygNXmkCks1DFRW7Mt6/jd95Z4sdDaR5vCLL2M6
FB/Ff+rNvA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
jFvcfNCzhBWpeT533DDm5MsDXv4GiB5r4Bmmnk5Von/5jho0+BIo5IwIRMf+AlV4xqtSYYHC3I2k
BVrljYddp4kTGUJvHCrm4WaY6cktxQlEnZCt6LbtmRJq5bQ0+BhbjRb+yhnUtxVO+mqZJ8X5carS
6TiI+a3eiQyqjafsIxQ=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
3uk2ioXVXgv772p2rHBKB55nN0zepBz6/NR5erkVu2PDHMiL0sh4KhStRZxPeDNzjzcvfXxTocKd
hKd8wwyqbvI0xJMti7Zm3ArPWxG9sxsPGJWi/HV3nwjRdbl8Q5i42ko8FFW76K8gPbQTkcXqEX+f
TMDFgnzTvHtLMrE1Xm+zXTsDfz2iY7i6oQ9oV094lrdSLAt80D9E8ysTFrLsOAY7rvOt1c8o26ui
lfC5xFONM+l+w+GytYmCYLC1g3/Ymlqj+CUT7JBGrc9OLEVB2jBY9OOPdBfOl49VdH6n2k4l06g4
tPQ+CDbASlaP1IKOpWeipcMMiP2EcvQEvzBqvw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ODN1qSeI0EeO28pILhOMZHx9bb2qYpmwvyQXvKPrPhpTBylybxluT1/v8KSBCRH/tKp0Ke1TAM0D
rxIBcEp/+xGCTqhzkt5p1fRCsGDy/1Kk5L4fYaTlJRk43uSfOTxn6cMlcuTzjFQ5x+FkobtNDSvc
hzmRwInNRUY241xhR0o=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
dC/Y1fV+mqTG5rOr6IWyGTQ8KnFRPeLZShUWaAXrkw+Ng+xoimVrmPwEeCnURpwc/T0yNbEjCDB4
bGeW47AlClSVksRroIGKMbG4EdH+85GyM7JEd8UxBfmIEn2qUdv8H40fYW6ndPlPBbIsiprcQqu1
BO1TrP+zbizezYEZNLdme7klmciNF64y46dVM3KfXIDNKQvoLTlpJYClTv0K9dc9pDZOVD/5ly4k
Nh9OSLv/jIhCDn0y3M3rX1DyQgZeJYBkDd4IBP3NH/wojvEFQZAcMKJEqADK3qsWu81U6IIzKfXC
PUyRFWat+MUxb64pAuTyWw3derZjtBnOfD89TQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 54432)
`protect data_block
m7H7/hfsy4qFfuqncGcuU8P9arCUg2eBH9ulPvfQ5OOUg/AsNz1uf+wthyUKu4hj9cpTnxX9bi4e
11Cq21Xx9ro82LKLcgYT0KXTEUOuLEgAH6lrAWbW+SmBAha/4X2au4JJskpKg7LeYhhD8Utaw4GV
Vx66CEQmDrLK0mGSBuWzMK9kAJ6hRgUVZqeusXW5INRDVNrMyPMExOP/T1RBginr9QZasR/BYAOj
vUF0wECkBrvN/Hq78BHjq0ik/YLjhNLT5wnhsvtzslrqWHS4/ADlD4rwKP14xcv5JH7a4heb7r5D
U6NMWFTM/RuE6vQ1CWjTZ3s409UDuQwsFY1xub2way1OuUwsepXfQ+AN8sBpdb7mf5gOxzozgWS+
AwQKW0SR0hsB+XN9Cql2gBhztqsrEuPkVeJSGU87z6s3prvVvV/pX0npal+ePGRNpq/ZXGCGJRvX
Yslko9mByGJX4SDDGNHSv56KktlAkFGZJ56rnlq7IeZHcgoftnk7jNB2ak7orfSDP4eL6bG7WBN6
z9pHnucM8cViOqpAcRdfYSSu9ViJ/cbri4m6SQNjk5vqYlqvNVWeCsIaUO8j+AtYmXnFlIPNuTuU
+WIPjaUt73Vymev3zCTmVPtK0rW3El3kfT0jXFiCYCCpGOqDfoGxNeRG2h2k9bEc1FA8eLwZbfc1
cS5Zj6FNjNin9avQl1EW3EpyRH2cqI8Q0KSkVuvJzjnE+Yg4wkxSzjUZb3x+EoFoCEAo5Z9fjwB+
rbcmwDdAuB5ckcuMOs4VfM6PWKYEop333PIx7oKaBziQwNas7Xy4a6qAtOMngmJLK1A8kwphpWa8
UfQ/tuV9M3ODG0yvMQOJ3TSYD0ybDXXiYtr82oY0J49KpXZEhZgo7tK+mQVCTP+jvU2wA+AgkiW+
wmD67rvgpR+QIRbsxEaJ17bIY7Jp/FEy1OQo8sYfDbpAuqjwNiNGG7pS6STTsan7uI886siB3KGM
2z9XJ2AT0l+pRtk4RtTCgK4ABZh9Qv6T/FeomFdvAqCfSxxgMnuSJABdkdgWYSFJ9nTZwtAj04tC
x5OkM/g8rRJMLoPbEnBwUJro+J+S+CG/eB4GjhFEVprNYgdEeigRjR6XyYykBnCE6v5+M8zsamRb
3xfVXDP9goN6NO/TJPZnqGGrKl1zsrB3I/wJmOsbob32N9kOfpsjEQMSQMrVPyBaMhsQWdfjNfAi
vvsGwkIajYQX11NLmawxt/sWgns9BiV8cLk5xaMVFTU3T2zYAPGuc5Wg82+2HtKBx542s8sPY0I2
eFNO/u025WMXwh69VPZEo27aQnSR2/76qDrUXi+JWUl9d6Zc/80b5lzYfEgjrT7wp/wIHE+ou6Vl
lxSX9iMHYxxToxj3P7Re7V0rEYaEVN/zol5YB1J5FSuSd9ODZGZg/RkHkrJLACpsmJc2dqwISRoi
AuOk25Nyw5ra8LSCXgQMXHc0GICAkHiYLNXpllFUA55JXdCxQRXsFvz+wB3X8MFqvzJMcsjpL+SU
HNe7SJ2Et3KBIjeTf+chCrtZrKjOldhsnLYVJYJPBWZNmnYZPyqHIDMbcUxAkxUjSoPSMi0SmeIm
zBPI0e0abARhuDcAiPmuM2nP3xOz9m9ToMXeN1j0ujzgJomzKuHxtuwbrQOGQcwwt0rVlXfBmY8l
xUYFUHx2iqLdavrxBKkljLxq8ramLWfhxYc3OZv9ht1FJfe2qxa0cp5Hu8dWZjNMoUCA5Y1wwlMw
U8J6eGowDJFNoe2fRoF8bGjSoPhJ2is+u7q8LYeDbH/X3Hoysr8p+B90wK51HDA0FicCEmXzAxqq
kn5hJqJYJfXPMDC3czRlSaEAkWGMvko1xrfln42kndP7tMH2D2j1e2Vg06B64qLfJEj52gsyMhKa
tNy/IbFkBFLtTjqGnQJH4L/SrFeOjly92bWvEtLH/ablMWQYKgg5jcqa6TamEqLDPEurKShdGSNv
xnxin8bsh87+RCjVtgEB/IJuGRCeSSxEWep6ThYO8QzuDEGjVSKvMmr8woY6busYve6SjdI3K9eu
lPtgllQBjoAz9saBWMJgzELTmywzvvD1j5j7tDzX4bMjUNCE5SCYymuKLq5SBJ+DPz2/E1zTmMNq
vTsHvVRejHDTG6rOqXQ3QwJeHVRJdRmkSnVENi5RD3bhZrq3KtJtozbjHamyqc2044ana6JqnkKy
hMn/nV8SrT4pYKJ9/jH3gxg4eixMxswx02LJxJ5S7SJIVGhVMdIdC1L/aH8Ydiht+TUejs1nPsUO
kdYjrHUBwZmrr3rYAjothapExlDyZNEaCq7NIi1Zu1kDkG8A8AqcCO/RrQ6HKKIzc1L95xpibezl
6O3eCB17fD1BsOevoxGX6aIJFEpDhNIZOOrn4e9wCgFJLL33SRGeOZfW43EVsGs+TqjVNvZyiWe4
9yohERITFWqlJAAjTx35Taczc6N7BGzuD4cIdMY2dsB1bW/jkb9MrHDk92E9dlMxNE9z+jjrkz1+
p9vo4DBqcZ4SVCV6h8os+QS3rTD6RlOpKj+tnVFg6RizU7YmS5DJYhcim+AN/u1sYUuu1evz4suZ
rfBf0HZr9w2XAfjmVPe4vh1lyI53pv0pmMg0etuIvRfYEWQv/JgAfGazbmuDKuCSFWNJn1cnHAKb
1NEQ15RpKaIR7mjPlQVpx1uSBq0DS0Le4WcMMraZeMpZlhlREsK6rtQjibVAlf09Kk7Cy7xCWUYD
BTWn4wl3+UwJOBvm5RQ/5U2i2PZP8wjGoTJ4pw3re8GxaoLrldRKEnk173alLBU0VUg2/5fxDngl
R3SX9Zm5vNTqSF0gw+5DL8dM66YeykD9obAWhQcTOtow9hBUtKk71nXnSk7GK8DjsXr3+Nvnd/YF
fV153QIxxxQ1Z0mYCu1sXwHEWOpl680V0CSD02665/M6MpOFaFnpw++ErTtCZYPEhYimI5Aw0UIJ
RFkMGaWAcONP8ipiidQXOeJSIilBVAQ12ojknr1LnKVCfD1FAntD3rPflg9RnkcTDq2z9VfqMYaR
1kBDuBvozkvPq/6LzU0SJgSVAPuuAsSfWVMHw65fcGqgwehd8CGgY77U9aimWhNJatVObnPC/iAf
YSH3WcrTynUloIbGmHbGXbTOSpJPVr3/IlN8SdHbnx8r5NQvCDeM3R1HaR+j1yF4WOkM3xhFYzPH
MD6uZyiu5tUYdSDGGmXBWMPvn15paObmVLovTYzizJSHmcc5tMDKe0c9CMjLNRvT6QE7AHD8JN+x
kg51Lg4ZcLpImHfTMi8AeVv/71OwhyaDqPXprTFzrWga8j4yUKgF5ZaxKkxlJxsHrhSEp8ABzyH6
DQPesa1XvdWBPRjPRgYA9D7BmrUKtj4pc81KsKiQCN5QHGTUI7HZYvHC7nchdC4XPWuxNqyDKq8a
wkj7hztd0i3s4ftRRt8vgkVp8Le7XuynrjYiMzT5csq3bv4iL6BFkN4nfmpzPlaUGPnWB9om0stb
QHuLSGRIf/2uT7W3kwnYMOduLIBddg05CrO4+IcvPdf3iaOwUMoH2YVI4w8mCwjYkKKmNixNmXL3
di2o0GGUXQ/u6Umg1VZtNvFuEjX8pbeOY1qOz7h7JlkJ3OQNW2ZTZcgHX1px7bYJ0TcTAzrwVnq2
T9XQcnLtTxDWwHZh1/iKorezu0ZEsALEU6mr6lrBxmLj7dKd7U2G6RUeN19uxsFFxhUtoLdaI8QO
8oDuyR6DlH+bDWYXVRST6wCfYQjezQFC9yKnrD6G8f4t/0C3Jdt46rBkUGXDMTKHEgyi878Y9rvF
r5uU6pmM5p+799j0sZvxFj0X/EEF7EWOlBKyXh7I2FKThN+CiWQpBITNMNQAqdx4nMiNfcQUjK94
4qTiaTXbAP5f8/G1NQZ6OS0F7dNwY5MyDvYsKM3kDFbTX4PUN4YspHjJbpUElsI9bGoJ8WrA4weU
c0fhs+B2Axq/Rwh2PWeQcbZ/7RzBno9yju/TEMshxTIrDpC4wSS6UIjPW9Xq3G7u3ROnRnQfv/q/
fF2wcfw6FaVT/puXlwGer5H9b1KRipMR4nRVTmFmBXgFCynfWyiEYpSZTf929kUyzKmOScFdUGjD
yLX7jkBzRqnsWWpuPrQTdd3oxjoMCDgOtD8lJfDer4Ecb7lSMC9zEWbVeWN1oBShI/CFF3p1Txvm
waMNSKUjqT5PV2K4pEGZuI5HI0AmnyDdXUSyrs7L8USFE7uiExXMCG+H4jcqNh/4OUj2bBhFb8kD
zxiEsWwrYCSSHcacd2e5iYHsCxHZkfH3rl/UjNix7ft+rCI2jHK452bJeEGgC8mOPpMTGReWysNx
vK34zkcrNtNcCx9B5QG/bM2yXX0WibFKgoZnEVQ8cNrAXoSBsPM31EliUJTFgZwft3GViHG6D0cj
fiaxGquLSgwcYzcuNqJjmXm/55d77uUkMIA85Z69VB64cLzPEVhuuNx2mUwjG8DN1/FdiLcX4o5x
ZwfcwJXIiqL0yoXFc9b4hYPAGjQ7IoUJ+rc27r5qA2lX85etTPkMHcwMNlCPfBaydvuC18iG1lYX
xMAezepiu0n3wkZfHqM44CHvriuJTHYz/rzQgS84itaw6FPOpTf4VJfSWHv/7hYQZFQD9e2Di57r
YI6471ZBiDIFhSxPAUKO6JKUFqwUXJD2R7jUxoboGE44nXv0sLrJu/rsgUC8MS8DstOo2XGaJJ5Z
spOO41TrqQxGEzGU2OaPkCome8+y62SyXAvKKi9eXn8Gmd/6u+SDh2VYJEMxj+CE3MHCuqxbhlXt
PgrJGC1soxvqhEy1W3Fpw3u+ogRAo9lxOJk8uk6Ny45OqypyYBWsPleX3JYxHeM9zCsmzMVpng1W
lv5b/OSw0LVHAA/tBBC2+wb4rgO0leIh6LakH2kYBOnucaWAydlt1++XhTwDQhLC7xSuarSKan+3
btpUs1PBuROSSSgHwmkgfN2w4Iub7IBVEstkV1Q48EuzMaXah020J4OU5greCEmKXgcQmsBxVyGv
fwx4s2bSCK0Oh3m+a+5x3abbXLVzocRQEn/xUAma65IP96AIvfOTo3wUBaAk3ZCM89bMOYSZlYPs
svPmmkCAe49xDhHp/B6YDTD7vi8d3jJPF9T2aVs/zec/Ai2C6DQ9u0Wc9tFINbQSmEWAx8FrbaeR
KiwsKGeKZ35Kl64XcSDSvQtoErVoG1nOXuKtLxBLU5gahqNsftdwu/OFoy0cctcgseNDHjyCdt64
2lo1zMjrQvNz5HG8x8ftAVz2+2CJBcR3KOqPKpklbz1g/W7a/oVys0OxKTcfRpCFqsI/Na2L5Nqz
aXc6uxcOo9PpTaVMwrEUMjNpbQFfIYpdOr5YL+TVABZ0AYJyBdD4Sf4m8gJwMxN9jynsKos774Ha
s+JPPK7MZ0XESIVpNHU7hFhDrIgt5udx75HhlhbBs/E9Xh3AN1R//xSnquMn5NIZoYFdV9FgorqH
BVH/BHD7IgVad/uxkHwA2l5IhaPT5LbHdGFo/CWIQPKo3y6U/RtHvmyufaUlnhxm50WHNEP5IsDA
SROJHNGRSf7ihFgzJAP3usVfFUuGzFmkMtN5mRX0hde4bIQ2lBsNlwW2rvqmVbiJjLvvAJ4cKxKQ
/s72zf/6qac7nox+qLYO5FScnkMy8fOHo94ziMGTnNlnH6j7KsjXY+abJ0ZukG3YiwWRiTzcNU5b
VT/Y8QxFfzaCh6K4zpdT6MLmxs433xvUlGkritbuuGynL2whN0aHJwajZ4Ar9lgGwwNBHoCTl6FB
Uzp8zKMC6anY29EYJo2+vN2P2l/bGPopCMc3dWg6xDnd8On37+lHBujRrTrknJhwx1HcvpVzQdu7
XbL3YOY0LiKtR3en+fYFTPSZSc5TFdeu1cPAgWhwV/+rorkR8id8P56a9DpJo0yePmFu7eThsVzL
ZYrENK2afPVE7Yk0d2NvVRlt6G7wVMaR2ZfePEzMklN+gXhga6hiM+vjh94fF6BllvL0gOeKjtFi
bgWXmgKZhLifkXaNefJ0thf6SupRMgib3R0qEZp4prXNtW1rnLnfFfI7esLNa2reDn/GE7aCuIMK
teIeJV/HiLAR2ESJ5woCDFPnuriVoGrSZe7g8O//5a7zlNC7zSFGuFZrkxR8Wa6M3pwJMEY0OtJh
aWRfy96kM50ozJb4WWVoNmjpY2EGMunlsj5xwXPUyMfMq/bt0cAtfvItEURjarzZJgJAKbIUaiqG
VYpXyP7G7t1mFhtgAamO1NKZfXpQmfgJ/G211lsc9k4974uXLuZr+mRHzl3O09m+nvq2goZx5Hdn
ruHS0X5jbjGYAvuHXLqxE2h9IA56z3tipU+PT4DjusBbenDkNpuYXqLmdkAHlMQQZ/dRDwtzL2gu
Olb6RZdhkDp33WmGeoV+Sn6DQ1mkn3DVeGNIDGsNkKjWTA5+hU+PuVFHUbK4lkUtjXezJCZTOBIk
SUf/siB9gz35zNzaUtgUdUpKPaq+faoMlKTvbRtn8jbqqt35MEr38iL7i2GyJty9Z7UNfvbOfNaS
VMuoZh17DYR38BXqUII7r0g3qZYQgQeYszegBwMeOkunfE+lmmRw1VkNqC83u9pEuC5VDiog+PQF
7lfaga09kLJQnVs2MVvOQbOvtC5D2+qx6pr49jfzSN7oDaPDgxb/PneMVKjM1AyOsWvxaKNnHT/m
jXtPo78tED9RWsDzDBk3nEowyRs9ezpO0BTUGXsBuzUanTF2aDfgwq7NfT86+JDnDziaD1eMK9tX
n3KF73B6kxtoyXcgQyAdoSu0E+qpgDLTII1W6dydkootIdXF+mNKlEueJpurTChdH1IFbEBP7LkJ
yoGlc+j08JitDz2Posv+yS/U/lH+MoPheTVDlE+uRW0fW84l37uV/efLjnxnRFwzKUeHCosSMiN9
E6xIvkbS9YK/k9nHNdpauAODVNdv7krCSbyrNU0GEPjCCUfijWTjQ+QChN1VLCrWZRuAUrVm9Sch
iD2ltam5MQqt1P/CDbNr1cmYurXYX/GyTuhE30xFAwDDTz1iBtYU+PsnmIFmv10o8yhqbTXtkt12
BI/7mIMYHp96om4AUd3dGnEoZyjpASSuiNBr4AXsfPjwlED19rI9ZfLtM+PZivDDyqMUr/VwpB2z
oIHnqYuO9LLA1EFTdwcyhkimqf1R8SOOegbVIk6jfhAhjjdnS8kVqwvFTNDeUI0aFDgPdRwgclYF
eFWMsrPoy8YGUo7YMIboYGlY/a8ELjdrBz79YifgBBYvDwXc5XB7QlKyNplz6ulqgqQkAB1xk67p
9/bAUV2odt+S3RX/LeEs5P5HhsjDAHsKM6IaKQYe4QiZ5Jo5Jxl4HR2IDUWfSQj/nzePTjGyjXAO
lqPhOogShrFMOyFIAWcBHlF3LpeM3a7A2pw5RaiOGoGqzigBNZPaIq88t0rVZS7WiF//wJwQchXK
oSXFgy6cHE1SY5PeacZD2oQsNIEqvewvZbWhQPgpSlS3tXxY9k+09LxW37gPfFmwA8wJkR/C4Ame
ZX0jurQfuVYXj1UVSSNtQJoOPRyOAN8ST+0QW3abjjP4L6EdgWebZzBeTYdte5OY5cDjAG2MD6xY
1SILYKLwXMODzC5TRWdz1nqHouve+agkYpUxPe0jzPSfu//z2e5CqDXMFPsNzGImG1dCkkwp/kNa
keQ2jBv1QEDY2UFSBahj1XzINH4kU/Kr05M3M6Dhy/fjwHHjVT4Y2zGhaXa1f8J4TO/OGmBkBUj1
ZVH/JWaldV29SlXodUVzeCPU9im/x/w4VxW+jJfUvqHOD4WlqGhrQ5GPbzKkhQMig8UIty143uXQ
5hVelWideWSWtNh2TbgG/xmqO3uwnDndhhGLW+Mmy22+X58r2+rd4CVNGhTMUIPuY89Ano/f+KUK
Xqv4vMv6PFuAlPPpyIuBrSlBy8vO1xfFBG42F/ni1SclF3/XUfugtqPBCN+2x0H7fqc69vxc1qDY
oqKrY354ZLExmHm42TuM9ohkDWPMPmZpSKiohdIiBwm52tysW96OdpfWI9cmmUj3IKcopXgVPHBN
YOxw0ovx+JTEHSD7ucmoaFCdgBxH47dxWFaL9GaXLh7qxkcKP0KdgbcQLwwz6CPA4P9D5wN+J1ft
2mqXmWwQelk5eOvezjBQZymPmzcDMaRRRIAEy5tRXPpj+64f4aTF6y+hz3CGVZEdqJfUGmtfnEIY
ntoGj4QL8S41LGNq7SyDNsuaVWQSD/UYYXBbDL+EG5Gn0KylW6wXFWTlAF22lYU3CPxWeFyoVwvs
jmX7ytB7PrIn1Z4wmnOxLj/VtrrvM3l4szq0y/rok/+UFib1tyb9ecq+R0j+65xb5pOcex+e4Aro
Vepv6KGFegxmOvwbdITTz5tV34ODHSc2WzXqLprFGAAxToLBfqDRI358lSfis5YvsOvbdbXn/Zyj
mb8oE2uJfz+MO598ogW4XlCxkXqwOauR2SwXW8Ox7hEhE6H5I80M0JVVHmO4CgwlA2hs9mpiaJpT
U8cCsGbs8LkD9GLoCBaCI8PiOZEYIR1vuroO/u6cg3lm60WOH/3XEXuudqTLKpuqJ2IFvwKdD8QS
/2DF7aEplmcesuqtmjCT+jYJN+nLZWyMMxnc2GhELVzXoBZcyF5nIcmg8qlxqQAuQPtBTCte3P2B
gFu6/YZzb4bH858LWrMUs3DAS63bT5D1ACQaaDfdmMbVv28q3/PHWkHbEyldjluKaSiHxQym5gK3
VHc3mL9A1xs2ewVFv3fx4eRY+EllpNmcQBVtTZqm1KOBjKAA5w6JcmUDmpQvcMIKOoZX8t398Odk
6Wq2aR0YaAiGv9n9gf2LCVzaklfW0m7adpOdPM1TY7I6SCyS4kGHF/yoeI1lsxlkeOhlKOUY7ZRb
kNuALR1A321RzG2HQhzkAR36tbZWhkxUSPUT61jhanjeZY8JLbv3dp/ybBbKQ6REp5aYfvvfK4pl
LvTPYcLg7syY6S5uNbz6fevsrVG21AoXDP9b5BC3s9Lx+7CyPpQnuwdRVGlhsug0UgUJHw2nvYcT
RSJaxp+bKQVa5WqO8Fy2h7EWWtRSbmynBTjgyu0ZaIqqOZvF1ZRBHFlSKOnDnJLhRHRRY+vauBow
rXCyL8Uz1VFy5DWlM68qjRCQvanUIJPSKAD+QdFA0a2JWqfKqS8FC/NSdMZizFR9V0YTzVxb5ocD
yw5W3OmL3Hx2LZVanbZ5gr26Xnb+OZJyavB11dNM2TiL9upnYzhclPU3MzleRChUa/iTO5Ucsh7H
3XCdjBj4/REprQ6Hvw0zDkqNvGmK7+l4UFQ7K9EdmjL+PPUxzZdXGslk7CB/r38RIT5KrycTsxBI
Nwa4jzJyG6JFVPIOSVntWnW1j/nHCFw14oQ7Iv1HTT65bk2U8Y6KA01oHalMklPq2bGi4S4OpjWM
PmNdasSIdF6uHGW73Ug/7t8g175dxPc2a6YMMhZEU30jFQztbvCWGWwtm5QLJoSick4UnfAKGl5C
St3+k+KxoXkDN2Knq/+GE4CwKfwNkOx1+xTAsoacVnYB5HhjA29rIMC94HqqKL17CHoOAilfyWYB
xi9AgvvyjbhvxBg6+6X1Sbjo0HoJglyAX+V8A4alh7jxXBuRQSpFZjRDieZ9weDEc6wBps9JggwC
ru+ICKy6lML5XpHJNJJ3HAQw7RjrOEouAxYhjTuFm3cjHYLSZSg+5nTcXM/rs0YDZnMqTbThGXln
nRV3xKxiWQ88W784mKuv5fnfjNvXjn/oXLMFDSSBQ6lM5dt7GTi+sAQX0zNcjmuwaf3w5s4slyBk
iDHpN+S1oJbw+nr4FqfSpMfIlsmbBWsBczgV39Xy4jQeyMFtlKys3bCqLnitdGGGCer86AN4CONM
6jd+MnwiX0dtOHc5csc9fhaNE/ocJ+vOh4FDcUoxzi14d5nNqL8bA3iAyUe3WoXyNm1oleYOcmbQ
JE9F/PTKPTFLG5T5f8t99d2o9P0dRWK39Ym9v6o89XFiHAoyIgCJaSIcCTznzfgINAX0gFbAU03R
X7o1vndpdTzvp/9T8fdzssde4sF/A9mCAdRyM2bOZaCqAgqwEjMOkqVdqAJRVGCoLpB7ARIW0/21
IR5l5Pn26PjYXcpp5G6/EOBroGKIUsmA6QK6WPi8UZs4wb7yAvkynHxbT1ZkPNK8PPjUiuJiS9TH
6eJ2mQcYYOH5z5z4e5L8/iB6fTpWG6x0RO+4WfvW+bfMJ/1qIfcCu+8iGFmdRkKLz32S15BW6egW
/TJ0aA8sK8KwYhQGpi2jxpIZXF4ZRGTOgGdtGwsGY/C8GnfptAnjbVSltbPoo27fAcaTE9zSE3Ja
HPySg9NDHpSSc8JTu8e2q+TecjL3njksmZh7985kEd0WgfaoEKjgf1ua284rbS7HsqzWnzpa+phr
L0p7EZJHn17PD6u22Cqob5owJa1Lv8D3xSjV2WROQDJRCNp4DgVtVw31ZtB2XxEA5WCwfGSBAGoD
GMrP1QmdB6Kocwq66gbGsmKhpB4ohwprzlAUtjo0Zp0EjyVT4AAsDki5FPWE4kR4qk0KWId4eMRq
0bp2g6arD3h049ci6sn6ic/Xg29NQumro1oScKybq0nqPiw30NYKm4c6zJEYv8PFHA7CAG2sW3NY
v1KpTXQY9eV3/tzrn+R9RNlYBOvXTuq0ksDK/6ikAyklwmVGexW0QOhBxRzN34pvAUa6ftVWXiA7
2E8nYQ6xBYm4qXie8Z7GnfEsE/FwPv1kHCyNuA3HECOvPCHZJAu4QxXot41rUb0hdZG86CPg8UeH
rzXc6eLUm+8vc1fuVHjqrizRtWe+4URHP5X9Fgz6I3sSzHJg0iDOtze1snkX+aZq9t5iEPr46ghZ
pSWA4xKqEQU0YeMoTCVVujKlKpy/RLpUN635SH6sH1OJU1uFEwlGzOxGlaxzfTfqXth0WN5tvjCc
1hjFCGo4zxhsic+/8lwD2UR6ZXOynm2R5msaT2aPJYVyHkoUpfwn8WfjpJh+snhH52IwZ43RsQT+
uV0yAK7BJsWpARMw3uJF8IBf18UkrkpTkpj9iXzyvgauxSt0uiM3AFM51GR1/K2cmatg3VfF9ps/
aIU6bqxg7UQpn6HdkQ45FgTbgLfIRb+dQezz6wKdwbXQLQBmLv0THnFNjgo02VvyBGasWLlKT5ra
bKnfjKXNLexaMruhtstH6Ih4y4AhNkhIBUxYluikWiCcFCp69xNUlTjLkMaMjcAQI0gwK0y0WnlU
IQBszcAL+zxpztweyRoSKtZLC/oay8MPQu0WVglYeBxaUYGtR4wkmDbhHgPNor29iF32r/AVY5+5
rCpVgxOMbo/OPkOrokF23CEH0aJFURHsSuL3fmecegxyxsz5ut75M3MgWpQjBaDav+ZGC7HpmwQT
73AyQ1HDmS/s8A2uide0Exo3wRDRJ33OqT+/XYM4DmnQPumQlskdXELCk1rd8c0sjC3qNUFLgm+G
5ifEplAVe1hXeKBV+AHtnXhJF0S10/02hPYzqL4cnJ3BuDLn8UBDHRYZcnCuMMc4Q7VxhqSj37bV
xG+wI6UK7tNMmuda9EmKm51SWi0o/5yiI2DhNqEZvf88OOynCYi2HjJyuPkmJL0zydvPKt5o26JC
XZXX22KpriV+Zms32ku6cYsgKg7vg+tgqVGSlp4SqgBVv6tzP08kipSIvutRY3nq4xIPKxVCnZ0o
y7iFSnDTC7PQXhmH8NZWmwi65cHNLgOhNZ729YkrvlentLiRFsSYDR/N1E0aDrWmpwGaUcPy2x1b
k63mPzyJE2OYo5TGoS9bj2912gZLZL3xsApP3FpriAB4TiPuanHe58mZmhy5qVaNg+dkUN1sRN5J
3QDklve27n1luqGAXWmTwvfVLlTUL+dbCfuK7uXvLsOqm9FCgOyihYr7WPMRQbArq/d830rHaDEa
9v0UGSacURE4Cns858H3ND3JkTFrHYtboUrJQ8V+1vhGM2XEs5UwasXvfcZhrk6PeapvH2GoRGph
wyn5AVK/6OQnA7Myy6n/LVJIaiNvimUzzuhmnJ4rODb1N0gtCTe6GknthBSU5TxqaPh5BSJroBji
oO/M/QUa7tPPL+fHLt7lcpdk1RLemX8NBOPIkV+m0dG1S5dhRhnj8eV5vubqYo5Ehikjbzo5V9Px
dbFwv9CHyM/87kUcimnVTyQgOw+PYnJuzSKzLZdYSJ9LlYmTdYfQBp12PsFPM/MNvT2L91UZ0r9r
M106YpOHpAfL76HNiudIgshOiMd2zTwtaUx8YVXer6vi4tn7PQf94cNICZrmRRGcGaClNfvneg3X
7Ec6iGA0cGbYO5mjZMTRx2TjCOY+BtIjOygTeevc+H5riH/Qa9u5KPfLsMKQ2IJBxhwAF/Wb9bwm
yjJKWSV428RrgXuSgaKc8rN2Jv8Q+Rcq8Mlzwd4FRIVKBqGmolbuyCjb7LqKiM938AUl1dUU7OMH
tg0OVwQ2IA3s7nWLdWx36+mJTLDr5FAz/chI+DJ6mO8M0hznpn+0wdBQ6QLLJX7bgiHFOJR6kFs+
zu8goupNTaln19qhQR6niBnhQ1mDeeih1y2VwpYl2QjDPnRqAsxVv0v5xXLo7VJZbNbuOZIJ5Xcc
XZuz5v7LzM8pED/kBPpzF5qIBYYVhavsz63BULWuhr5AaIVLSi7zlaXxPNLtNrq4cGuibvLEkJXF
FVIhXMuqfrjzSiHmKdGHIOsUg8a5VUHBL9t/UauE56sCWG+NimzN7XOt0WaTkw58iAIfp4USm0FO
e0OfWEjo1olrO7vITXul9ZObbZi8I6JUNh6xStigK8C2Wpq5l3+jsdf7I5d+w/f683UooPWy7ylB
O284/pthnTdjO4ULc+VXst8y/9icroEpzzwPJQluBTrvcdGMy3ExsAbZtyBAlXCRd8xRa/lAgNWC
MynOfiiRW1CFzSdFRR8FXIQyzu1dg4w3lWCvVqj9QmIscZNG5fAM0OSpo6M4qds13RlsIBVF11Lv
iN/CMO+etkSP4bN0uPiv8AUZ7cBagEbib9QQnY/qO7SjC1JkKBdZ3J6Jf92K6oaOyh1tBj9QEI94
IiTEgnWnib+HRJQHbH4XxceJJ41iWuBxZBCx5JQ/U0YwS4oA9TTARlAe6wYLU/wMN2zDgolwPaZQ
hUGQKk0/k0GyUxrBJqLFNbYr9VFtMxtNG46jhclgmREdFYjw8OW4kC5oLv0iwVK3gVYHFHRDzwUZ
4dRigLkr2c1+ak1VgyjfLrswksIUKJ4OpFuDO9sQUqtJdTzgxIeouxZLwyJ9Pgjwh5AzmbCSB3KR
6kgLWQVZ6tZjdGhkd+Vr+xVTVdzBZCd3p+vIT8lZMZXvpyOqXX0dQTJdlpMNPuk4GGjHYSaZ7/ls
UKUWzgv+6JdeufhUlui5AJHXBeAcQMbrBN7Cn/UNeecNqL6Q/zx877X919Z1fXJ6va4gAineosw8
wrUOKIjWU5X789f5rAjMt7hZzq1bsPnF9l8oZ/OtBOkcZ/cnLsFqqj1JqGk36tg9UiDY3NsP8+NF
NxxSH81mVBxfwEoYBEnPadh6FzA4Tsw/+Gupo+ufc53tDtg+zjXgH5GDS+CAGxRbxTMRDBR8oeAr
EUPBiBG2YigYSfhYjtQy91YZqZUQ5GsvauqD5dkYqs5hBA46osFIYBbq0I32yYnq3DUhPi/3ktXm
LbIT7TPMyX5uFHF7BTDt1V8u8FE3+FEHIY8OV2yfm6F5/3Km2MRjZ+YmhSX2zwv3rGkM8jqJVAI+
nC9d3qrOFFihVV0ZU4A2G49w8wWElrYm/e2+v26NwPpsEW0trXrybdJCDRUTgpiy3hCr2BlbM+t2
+qsGTsbzIfxR9Ve6nZt9NXK9rZWaLaQ8AzkRZ04H/SSriVeh4hIUfeh/9xzomuibwAStJTLqmi8C
I4scmXud22nNBTQUDabb9tUEA//bIB2oBKIzRvGgJjBckDnVQ5s7WBI3RhOiYd4c8KFM6VRZ9JgH
TGyE5ZliWw4o0sL2E9vmmf2FPk6OsF4jMl6UWVLYRS3CHhvmshTH1qwNzU4pmvHNqQUldxSlUGGj
hrCzFlOw/rdYhZqK/o+Afv1BdkoNAAwX+SxhFkGtdt71cyIZHNCMY2s+m5RIICuwfn9/QBRWg8oR
BEtUcnBjf6UPBN2JTBtYg3vE2VSNhuV4V8tfIh1WgFmilFoR2yvufPg4PiyqC0RkkJ7er4GBtf7w
Km2elS1FEnzKgh5lEfcG8m1qrQaZG7A1W5yo/cIX7xxNLBsppsUv3FH3aqRAJQhHwTRAm8HaKwYV
q4CYKhItRv7mF/YRp4IAeu0wFuEC+wktRvjmxdM/qokbLgJCogPxeGb8Z3DoKe/YGbXB4Fl4fdTM
iwG8mFD6hVRe2d3f2bVyluA63hJ4NqPBhqTaNOlXqPHMEY9kr54cM0iyiVcr75/QfaeM3G6w1SLm
AzPR6bdtgMvNuXPTYiugr1yes3UpWJAMJroVShrrO9nS+GiVdUq2Cnhqv3qqj8o6W+3uUkgXeTXO
syyLUjCm6Rg+OLhQCWMQR9ausrAPC1pmXdr5wF/vkLzuwbahMhk1ENKIaA6SsgjXYukgzY/KrW61
/yRBT7NKWQRjamTK6tZlTtVaJUH2Wvrdr6R8ikwdU28MLBSojbhYu9HbNIZeXhrUwG3KWomD0DjE
na+X3oJ8R6VbXxHJxRu655BklKPTElaELUxVOmW1btVqzLNtfD1f43MHn3vCmEGp431BU8Gxahh+
mQjElIpZAyHeRITTAtjUTYMOFkH6xQ8zacVBWLeSiyvkLVYpO2LWgMa4ipTOFXr4znb6dxlgbO1e
f2/Pkcaw6BjR0LX6pQGmoxpjs2ykv1DBSjCTJlV2flm44J28h77Kzoftnk4XiyTWsnwqEqQutfID
MolbzH31oHk6UIt2MeK6NJB8p4uXw6TIgBugUeraBn0f0adEzDzZfqb6uYwM1C1mWZ30fLxCBT/v
uQjd0it+ia/caWTIao0JGKfRFW9+mMIHn8cmEDw8Uq3rtA1Lti0pqKULnRQ9EksgMn1PEz+GlOJW
yD5sUXBvplFhPdtLWNUH1DtPU43AUnvbn9cXq3d5srEVkDS1HNv9iReMPJejWEZ0EiLoJhvXBmjP
Lbl9xvzrVf4GR4X0ujEbp71VkimVPfrpnW07xBY7iAfLRQCNtugLzYF2eiLqE4OvegKvBRMGgAm6
HZtLJn0Fyb4ESdCfAkXOzB6cbpH6cbX3au87C+k6/owLS6sLMWWDPzH8fe+o6q+F7OLFqX5TBGtG
SY2xFWV0BdcfGsfpCOr3IJJGpo87z5Kicncs5ApNtmI30Nlx1yHL4DGRIR4uAccgg+wFYW4ym14H
btTGWoKJ8NkLz5jJTgcrw9F2TrzLMZEBYg5op4BD/RiD75eRzawwdFArAYg3FQerlJHgp4wEFkpz
kGr8dbk5UJBF5KJ96QjSXOM49veVfRNKLvp7KPaunjdJYb0MM4bH4thmdocXqVGPaushKgmK8gnf
XoU4+jT4+xDQSMWhTpIWR+AqukLPeXp8p00sPZOTshnuoPbh2pa9LKSQ367IQZGBf/N/aPrDRzaj
SYJdlgEHrlv3FVhAcYd0ISNXvHZEf/EgwyZHKg7dMMoRFf4jQ9q6MiXdiK1hstDEkCNC7nMmchuc
L88/xyiPY5MiF99vcE4OO2NaRj77ibXNQiGBabr6RB/L/c6JqclXULgZRcSu4epZL4l4BR4WN1xv
VaBbKqY5jsCD3X0K0fP/DPiLRAporuCXzNmgHgF7E59tjEUX3leWRjZY9UlmbrcDsHrMrl1Qp1Q1
MgMDFJNXLmOxkav/QNQLTSXOO2NY+BKc7ZQz/Ey0HYRKVmoItbpUSvv4OVxM2E3lf4vGbeYtEaNp
2oduA1/tdwTXbK3Aaz6stNVX9Qw/np0fx8sJKdDNsy543zmRiPCGokRTDTR8cmZ1NW8YMQji2Gly
7NHdlyejIADyUhVry7pj41WI61WezszBUQzZS/fhbNK3udUE1ILF2XAsmwQsxy7EG8/5PrXakj6s
S8XoWsuN1PZS21XI0663AW5ak1swcnNLtf4A7lmjDDJvGBbcJsFFNk0i8wPEcZIlsiU37ZQ/6OhZ
x/ilJGhAqcmZ4jSrcDMKIvBcVVZLFOMjhko7YMJ/ovgMQasVarbfDqQTJfxhe3rVp1ZgBZbdmPlq
z6rXm3TgFKY+9nzyW0Afi5eeVb8mm8dS7e5Z+OU05DmsFPFQWQR7lMewg5ge7lRhNL2T2Kosal8X
KVyG8AcKuxPtpWQ7+Qgi2Sh1/+bxBUNvcKB9C1GCk5RYYSmzcJE4znCxUkWGIg2vdswR7A0J3Tzl
a9ocOWgknBTL27FbFYhcKkAFBZUZDwNi76KkYillqIeS7JI6eN3uEkwjRiX4ct5YM8LGSoS8wfQ9
7fzQ/SYVOXgRoht925Ngs1+nPq2v8d4xX2uVd6PSN2RqbW+APmPOr+P5gndCu7SDEESmWepTfgi+
fphBQ3mC7W5hZWeB7nNIZQ4LctpEJ9c11S8k+Qd56RkUcd/Y8T8QZ+nYcrWFPWV1THia6Bnwlm37
pO0Q8wmnYbvmIWrZxzxqMVTCSyJkgCC7+Vsyw++gLZ4JJlFdBqhSv6YsJZ0xPaU898KDMzjGFB1k
Jmb8SQ2FotgaNVDqOUIWxNTc0cwPhlkgr/lUigZmGO2IwsJIaI991hxeO3VZn/1RYW4uziSXvI7z
qIxtuBRIb4dRuQcHKBrLCJ+zmTGIzL9HyqItz2WPzJTWJ/P0hVOzDhQCs7QN8e9IF1Wd+xkH+ifd
ZbHRh+V1b85qKJhlXuL1ml0tOsq82u7Rt696egkx5MOEAAWQnN7NuaT5iKkOfTaMDt7vuyu36sk7
Ipitq4LEtMOV+SalyZpY45q80jDVNz7jCTAnvHE8JcB1M//gspRpCpbY5UR01+F4fAiplrw7mxpj
BP4OVd6Qx0ic2G3E4zyRhF8QvFmTNLTBIdEkIHkNTu3k/onRIqBYoIOfZpnGLC0fMbTAilekiXg3
rpT3tgjk651Z1GVTwZDR4kJKcNKMvygkytLyKb/XlnYSRdqibDup/HsA1lNi+VrPu5u8rhgdEZ9N
OdSYZimrZPJp1zE8t+U0RXDpRGx+9kMWk64XqjK+GEo750CaXZKmXjX44kf1qlb0oOyXcQaS2LXL
ysTKm3LXGu2RdbzYh7YMPJRV2qcYZnUdFg9WH31R2RK8C1CFrqpqDUw9cXRVTl45ikN9Eob4k8Pg
MCQBAzDnWW/1X1xTXwHR6BRA5d4+zXA4GL5vxQlgY/rJ2aNMfyz0MtAGkSPftBphwUwaaQdUwL6m
W8n1DNOCRyMDzHgyVQY/zS2KKiVRjRlK+TU9Mip5bRiRUzsmj1kxJ+6Qo60N9386OF2LkOURdjBh
RM1/2SR3MObVCiqxSKp/pfX8p5ncTtBAF7ZSE0S+jz25efCUqjTbO2hjljO+XTV26bDeQSkKfgLT
HVrf3amW5roa+8rNIiu8PgerFSxh7f3vLj59v0wY8ZiL4mfyxS4rzcxCatm+vOdJM15ws/WgAZsf
OMCl/3HO0PVsIlQfXybsMR2PKgJzkcx4GPzTL6648vHlWDJq1Uby3FPhVc0+Bizx71r3Jhe+6vJQ
BAOgZVB4c/NgWahL06qj30xDAOQb2JSNsCJeWcQez4mxW4XsRowJg0YHoOjW10tyQuoqBkDpamjL
sFwU8McK+LGoDj2mamgXycUYEf4RfjaFBOLp7q2TQ+9YAbSTfMWIS24Jyj6TuOtA82v5Lb/l04UJ
9YbKdReip3mClky/4g1jPPNBJiWLqQ5XQlxTsTzd5c7rEdm2TtzFcrZOz7A0oVmWSMyEh+s5okKl
/SsD8qCGXTR1nwvzbj637isfwHfPxFLNy+hQkkprJbkTaTnnu6tCFyUlRaV8fm91wMPVddnsjWGZ
eHNUMvSn5uyoZtuGJ+T1Vq8gEN//HkambjGMcW12CzSGv7O7BWei16g/B+tn50iGDRsJs1Wbwgof
pDGmi1jC5OobWq0Yk6PQj6b6fJVvTrV9rh8bLy5a5j2OvJZqaLRL2RofmsuHoeb425Uzn8lo4zhj
X1uVrW3hDP3mEmGludOdtmI86CMn2HNPW9r5pNmZi0dZJfPAp8pRXRGMQEzAcDcPzbZZMhlcAhQa
zqywonsjQ9KxljhB5dul5Q89SIxprYvlTqx2CFHXpowjGYftoN4ObS9A+OGFKFUDHeGdEOyH0FdU
GBp4jo4WusWOnDxsyZtwyCys+rn1imSL/qAV74GPJE0pAPIhJ+5zazoCYgxhaPgbEGVV8pS95Q0t
4qa84V901m6wSVvitK4EFnGQR3VVpi7PurDP1u8AzQ3SllUKIdevoeDXvT7oV36g+VJ7W6FM2LkF
q7jFgQ/AgX1d/JXeb5MPq6INm3M/awhTxeR1q2gbf0+NyYAnyyaq4IpJLC0JpRMHhQ37Ne1K758Y
I3XHkZR/1bTzXe6mSHJedLygx+Kr50UuqdIZP42eitj+Ts1nOhY73IZQFuzsVH64uZG1wTVDGXvn
x72lFxVhBGKcc/mmbVvHJi030pFLPsm5zni71JGVptDUzspS7qsylyK1uKseAfQUi/dDa7YLbZ62
+6oWtmnKHPQMsKadryubwlQOvAmkJLCIP3ronAWIduqibODoXz7GN2BUaJoE5KinqgryQf7P5rpd
uvmvZdz0blNUXn+2xKUCOBTwPMl4D7VLwH0B76HvbBOO2g3jI9EYpMyHGXdENyD8GV9w1M8l3rST
5ucbUiuD8DUUHla4X6pQxtFJmXON8oc9aN4H4Tj82wk7nGPc7AIzM2glgIhIHy1FNQRb8ZWAyj3g
/xuX/Q4KmVPTA/9wUssY8/oh3wHXWV6gIi66KR/9Grsi/UcSH/Deeh8BPWdowRrqjm48Ssu9+L8L
7s5MRHmmk7ET4+dIuE8m9e1I0OQiHfWwa8c29G0bOC+O0I6zwv/ETXTZWeAH8PYG85zIgzXcV6a5
tVpW8MdRt+mHxoYPg1Pz1DshH6vYlinuhbTFALdohfKQSfscQAWPpvcnVokhcF2aBzYmaan3sYD5
FBYiJUFu89bkDkras2AT3NGDEFLrZFOt8kDa7VsV5fV9XyGZDImIu7PGtVt9j+rSbgRvX2E2eg77
rakouXPaQdqkUVdfkiyy6XQXbU7g+qMkoRJNrL6+2j0S7qmWHj0l+ag9g+nduio3SFdkuoTLBhMD
LSEBiItfncAp3tS/v9TW8nITYtbbvfdeeA7n2h9jSGR8d9Rh8NM325+QQMONW879/l+mkazhPEKL
NqGDebF6Og/t5aisxKfDIZk2dX8pe8+sYwwj3s06rCMUwi3lOwhreQcT8akM9GFHmdbB0SgVwPbC
/gYG36/FKNnFW8brxRg32QwiLqw0zLp01D90DsRJSoWY3ziku9+HmC9Yh/b55dyvAlH5runphsZc
uztLwGV9UmVCx646b7KJT8xfTfdo1iTbdJU54ItnIkw5DD5du1TaUsQ4+xtd5zb7+wz7CBuaD5ij
pyGZuDCBJ41oomSNrX4F+qSOtkAaG5olySMaDL8jyqP+fkWvts2zedJgtGL+yd/5Yz9l7wPu2uxA
PfzogM2HdYCTKxEoDeh/6zhZxKOMwy68a3qbeoznIcWJnvMDHdGqhD5arZTMiZLgqLbw8ErsB8FQ
YHdSlKx8ojL5AVVBEVbtzPKO6NK6tAryR3gHA70XbdT9zcGV9tCohGEZXBYIMRCXV4LbCYy9AwOq
bskVYRUF6L4TjeJ59Gin8dc51uzksAF0n2NE2a1cp2vSUjF1dlJC4w90l+JvPyDQYUGscHjKMa4O
86Qq2J0HSIZcmEOamw3b9xfVO9p+5Mh132Xc4odzWOVpjeaTXwcmB+7+aSY5FHUzOCk3u/uMvtdm
CIfmQt5ITqNPl5qI+pKy1KrAOGCu6YhpjpAtodd0s6Lau14UJROP6dyyFbNcilY2+hexc8P9gC95
89BwkOCFL1+x/CFxRBTHXhZEeTqnW6TFhN54/u8QEYgpaCai19HnZtsrZzVTEs9RClilDcW7M3eN
/qhHSilTXJKSFCJlMYZduf1UliXvq+S6g/4BNSPVEI27Skd0JIa3dvMDff6WxIh8fCJaSi4lDZMf
fMIW8jotSEZ6SzJgxfwMmcLUgn52fnpwSD7830DtiysXEu187dRyO7vKEJPryD9/Z4pPzhi8/WWm
kGGW4LMk3lDUzuji3TAEuBk7zosb9FEYUtEYbfWDTllBbLLZryupK93G216p76sGGLAbPKBCVQxe
uk3lVhfkbyQ6mfGJzGPZTuf702w2pqy8paAimVlMTF2o9g1h6Zqi0BMZCASGT9943U4Qn/Xndrjn
nhWnzG0z8gU+dt4QIaCuMKhJyw5CtUTLFa2rT5EU+bEad6mFK+g7qIvT/+ANVb6uoBrhsBwho5EY
L3his5RYUhYa8mfftn6haH8xZSiy2kJc7+S0UzuMfLS3HNKVRuaHEMqLne9NE6MrjeJp4G1IOrUN
RJ7fpPgfo+Yr8Kp3tMnqNqd+HnRz4oSPGdN50MpKCA/+SCH7KbI8FMbRUOSGha/Vt/R/ndl/+lVp
EocbNW62Gr8dkt4qoVllNmiSDbmQF9ZRMFTavSShMly738110l6lRuSHyFvKcEDycBC1SYCyKzCJ
s01mnrGzcLzY/+AopcM/q0z9Z/aQRAdBoKCu4pi21b5PjMTuY6QEvk0nCBYuAkRlKKUbm1FvymV/
1Oo03NNpawF0HhX1n1OG9w1i31tnCKMcvE/pHjvOFtTMZssEjWnA1BOjbhpTriIjFfx9vYpnnmFk
5u/E0FlmD9Ryu17fIL193UsjUj0URTFlQxRx7E4Y3gDiprVt9j3grbOY7CI+PRx28ZeSMhl2iIa7
yirkKYo15OQnuj0Dt1GPag2F7DBeYGQVfoi6bOBZcBO+RJvq0ahlTWyX0KYWBKnnMqx42mE99o28
2KRyhLNaFNXlxwFNYL8lX/S4jeo5VpaD5P87axNRUnfL3xqUD2EwNFnUo2jELvXbKgqMs/cGYttk
eVEKTU3rKHvSYfCcgbbSS9xcI9c1r7+O4oqh4Dh5K2Yr+7b17KSRvtBlTDGSUk3BobVjk/cfNqL4
Rn2lXFFG+q4UfyT2HnXeoQXovtn5g78HwgaA1F8p3iXGxAD4MDbPJqNeWE/pvuZPZF0j/56WvTaz
JlhFV2usgUTDBDRPA+2snADIu0QjWStccQwtrIjh+AXubNi9ZdfV1kmdIoapy5uoQch1Kw0nDLUr
6beSXLBv5YysGvXCkSSSfbgZ6XSHQHIUeenWkgFYeWR2vfBoWbpyhSMJHK/GDu4A5msF6IrD4opa
uPF+ZGT7Eytvx+vISh3XzUqPT+eCs5RP0qK26vhDYRlqx/NZTX86TQY73FCesejXRkS7ZHRoKdn7
SjsMYwwBtgyk2mOywEm4T2kQot0VTzLQNRx97Kkb7tOIkraA4Eh9SajV47bSOwlEpRFw9eZUf+js
CliAFU9umIBgZNEJHQrN6+o0KU+CGT8cFdGYdga8CQjPsCsElSykWBibH8IHbjotF1n2pyujaoKi
drWNVso0iPqUNk1xbnzqoPw5ZBsfyrqQNSOEnXC4EUuOOoWLz9i6VkDh74vcMsHmTJqPznMQzG+b
HXrEJUghK/kR1N5xRDBT8WIJr8S9kCFYIDqUkocsA2TLpJYAyivqGrG3mwuTsIjOZoV8uD6EYjWd
7B0fePcrANCF0dB8UJKQtXVUkSpMqGpwRPblsihacYnGWSNBGuwiCOdDNOkFs/RcssKpbCjJbIsc
LvxHQ5Lk9LgtyUEwhzvRWMSGgOe0PDVNfbRASSvDJmBmM9yLs/Z2JxWUH7GsI/cZ8axIlDZioGs1
oc0mlr1GaL+cEHebT2DdyfSOm0T/5bsuhpb1v3gSb+Py1B6JKA0LSmRkR2AA7WLlmIRxYHWo2AdE
TTHH12/0T06rt4SOSecF920luXHXbbcJMAS3EVslV5ZUcdNe3kzzaz/tDswOffEEtzWdSuM5rl3L
4PS0QOyJPFvdTndqpVSYk+BnMg56HIf1xi86VPDmTwpkrh8f5+PHW8g/zJSdug84zn+UBqx6p3ps
uAXFrQVx69HecmaAH1G+RFfSKinswhVj0ivkT3snFYC3EEUHMCA/KnSBigp1MjjsIJbbfGS/L/rC
nvYv9RuzgO1Tn/IatX/9GR0xVJE96TJPklzKkVSb5mOAbMc+HZ3rlDilL6tREF5m/XQ59toHevAV
D5plfGqO+3W2L37jEjee542fZzOfLBJYFmskBAou5Tq8jIg4Rk4VDOqtMfnlWFBRpmj0Ep38tjv6
ZD3TecdpWrrG3YmgdVYcRKC3GL7DtJZ8be7QHazWyDUbRqM3LGgWah2zBFzEGEqKHvBP7OTi/Hw5
YxnVKzB09rGhZji9tFQA0BKhoO61x2YsGYA67P7OAYjl99bFXzf/IaaGuR7dgQEudCcQgdK7fMyI
yesedNJDPHInZnuLRbWsWvuAx9mdY3TbgxlRJQZLX9PAbjH06Jr6McNwBQ7C2ceDLgy772MAV+z/
GA7yNWEowwj8qxrxwPsIeRYFmhKTKNKgnTHcAyEO/gibNZXShsQ+lEwQmisg6RAF9CyF8BWiyB2F
rdwlmb74BAmEAK0ULvDseVd78pcJcg30ip9LREIeu2wgaJccjB2l8vuy5Lr8lxFLIVce2IIg9TSa
gTCc3DWApFccT/E7DLSXR3kSg6Te9M1QaAfJA+hqfga96LWbeMS4nKeN4ObD14qCXom3hy9x3XLz
VRYfwLHInWGU/Y1RvEeqB5QPCes2n35+SfsuFJ2sERGHfsYj4sa2e6rx8taxz0kiqPESxxKwiHzC
rrVG9fw+2JSztNLG86rxuWxyphotBp+3ETCi12mjmIaVdvobvvJ/k5k435H9wfcd4lh304hIVicA
ly5jfntQmX0Xhlg1PdLx4GEEbeZIpU8U/Q/Xu6S2yfGEiPma74VC+Z7jW5ZjKTpBbroD86jM5TmA
KvQcekutrxAgQ0Q3EVUByesk7OFE55P9D7q8cTR7Xh104P7GycPOuyyD+AmGeqvdhdhbst9pphlY
FKu+zO7INVx8N5hefGqrgaopADb7T8m+T0+/tAtWU/6kpESkn5Wd7bWAnSdnKB2llx1D2PaTHISO
F5fpQ3mPnrD5/E4JRQ9JMnPUa/MJIWyLOP9ke91gM7X9mw9TfLksjEaJTyB/uYr9brCGmaPolRr2
+bJtYOKo/xXycOU8LsCH1bM+rydj97z7wUEyGd8vpxYS3I6/AWpNwiU0622PlHbAiaTNEhyKZkgy
HPSyHtXTepjkWaGXsV9xabndbL1tJY+AhT+OU7TRXlU9tNwqrOncaj4c24ukiBSu94RpLS9WdZkG
Td0HuQyx+NTAsXwai17dMZMR0nJlrp0Hf2y9B21y3CWpAW4mxzrh4nPgnqB/WaLAPX8qDDfnBdnO
SSEL4IzF3jtSuwVMhsmGLq4MiqdoKutsvxfgnrv53Mgtj53bwbt00FYw+FiptuJfGuzQm8X5kR03
dyJwPzgTzTINTIPKbZYEe/49afQN7063qVVCWDjESFUuhSgyztxzQppbb5J15VeQHSJtuHzS7Kpz
kME0+h3PBieBeutrWQD8DtGk6ekDL6kqVMQ5xOppxQUS2kjSWf0aJckaDRFKz2+flOJraYUUQg9D
pj0Mc84UmAHljg6jMusFaPtfFP2bfZpwJjWz2wUC3xRE9wyOyf4DAzbc10QWdhd+28dQOXdCnFL1
yxVDIQYMGo6iYyIdRJNnuBSOFbc2ZQJm8ZGrUZSzCpCXZ8RxsgFz3oGJ4w1V/pq10jIYeVXbW1NG
0Z6OZvZfkfrOoM3K8xs7qHVx7cOJe/kd1RXhFSHJe5Rb1mcYg6tMU66pNJmNGiKPXSMlEsRGfes4
o4Ywa12zZUdA8y7dYLHJ/egF1tT/pXDVAHJEQEANLcKSXZZvxDr7xLi09vGnKs++FDnPvGFpZBEP
4nGCqmoc8XQob8oVgas8syUF99ow8YpYwYzP3qsMNsPWhvpS1cTjOlUzcNFu6cp7o8u1XHmZtE0E
1WMpKsWo4vGeYtprLMuiDGwSuJsiM/rw78mtS/B0r6YGU3NzBKT+g0No1HH6BO+CX6RJ0gCRQ0AG
LEN/0nlD8WQhgp5mhbtLb8Xy8Uc4Wou3hSY1XgRuuXaNbwxe5xziMVvpNHfgCqBtrXVF04axg+tq
l/xu/qXjFCkLgJRu4ExrwlLTlf9ECsZgqLnjovScReDDQi+0fMfAgqENlSlRlWP2GAKTUwlMTwIB
MIGIpbPuNgJoHlkOQE5F/sGjTwhIVSFFhaXkjggfCd/3elUSdgm8tUPG7HAAZE9I36iPcBV8k5Hx
AY7Xkr88wsJQFlsrspaULnJgbJw6FIgMNx0/QF6QdLDWGXHZZ9kUYlJhRr9f7k03kBoWxrJeVzsk
q+EObQ8vVnMUlZhVSNHX01jiMp1bkNTCtscsZduDr9t6HXPLLzIgOzO95b745uce/wz0xSwEEuSN
L6kFiv6V7jLDx47ju9UsepqWmEnMD8ltoFbQAxuqJuNJTxrgWXYXh3oWdxvIEXIAa6/yxrYYXHnE
nryGGZ6/2Xse7Ui0r1n/MtHDkf3U3d154s8FXw6AcncBr7sRh3+IN8SOhSiVpjYuKxKDILtkJ28B
flFAvrUomOk5M66seOjQ/HyGEt9DF83wBSce4FBvgOX9e3YzxbuR6L1Eb6xFSqgb0/K32oIBwwA6
cfj88oE8Bict1nhEvS7TX8TmlhU+SW29HhGbxgeSYvqrSw7Z5bff/MDJdKuL/wh0fASfCpcfUnGc
uXWQpM6DXX+ZoCbh7EXHwWHtFDwJEDvA7cfIzpAreHtl8gGqP7d1iP3nOAMEDkRIinLofUjhwBsP
xb72GYnQPqyRCExBY0v6a5m+60lSCW/P4fJ3IoHE4ryB6xteGX5XoZWYy/f+kd60KYoTwBNOdYVc
UujZyGrBxJ8pCcWl0csedrDuCfYLd464n3fZm/PhqbE+kODWMx+qU/8eei0OJ3KiJpvzjqoJHSLy
FPuhOuMLTG4t7eKAmtpGNXdmHrAGP1RHVu/vIC4XViHDZsL/53EohztZDDwvkFuLl5vFHU8rqCfg
9BqTIGO0U19JBkNYwtBpW9DEi711NUO5YEpo09fB8ELqj6NHvBBoQnVqDMM8ud+dUnxi+WE5imTK
IglI4+qwEkvzx2kCMeDJLD1ha6aSsmgtytz3fhqUhpIt+SLvsJM62qkRSCh4Ea1KPtSs7n+G/MQJ
ZIteBTwOCYM8OkJHkGsZ8aRmsktxWOefHPm+D3YymcCWIEFc+SvqzGRkzWdxMzT2ym11CZYtow6X
QooGrXlONbIZ34DQlaV+Ur1OijMCuCsct5aHiPqMB9+3i3Cq9JGWWLCS6i5cJAuNJW8EewL+Z19H
ljUugq8hurnsxpIhZcTsLZyvgxR7UCbKxZbf4frGdLVfAln648pBIUSSI+UAgJPED5eqpZECUoBj
UHm1KjGhGINk34jZdFFPgxg3Q1JXSYq6mwQoL4kjU3kTNED9MiDcLjCkZJ798dmqD9jfX4f0gUda
eYzf99VUDrU/2wBvUztXYXq/i+pdGR5QkFrZvRuw9K+KdsACitP19bB3CwoP4JUo5siYPygEdI4w
RDP6XIefnsFaG7ElMPb8yfJn+ypA9dp+S5vWpVr0rCgfSqdIESc0oM2EmPuDWa4tUI+eIEc8ImBi
j26NpmNMlM/QL64VDGEfDr19EjRCTMOA4MqUH+/jSQJamN0bNIkGZL2AfaQgATf3vKBRlfzOP9R3
QMm9HPs8CTXi5ueZ01TFwCuUAX4vG1yAsWuSgeyK1Dfzv/Bj8bi6iCeEs961lJUFeqRqG66j6BHM
8WR7EwEuuNrgKEqgV1D10PrXvkSzW9AzDpQxQZdrOR411aK4Wm8VBF5N9LIZNzW7UdksIEuB20zJ
gaLUd75UGStHV6ws0kJk334JzxqEanaej+t9ejYzJiZEtZonmSIwiO6eiMSwx2trz9tr/0miHwnP
ueF21KQiDZ9zVf/lqP1ibSZ7yKLirwN5McCKcV/fKiAnnGFUQlxxIOIWzDau5yFngZ85d+b32ocC
k8r2E8Xk/+Gi7EsX665539v8m/Yxvu69E7ykhNmQDMterKpBMr4WqiM9/mlxzpJB3mMIY2w9zU//
wgPWI4T3H997C3KElqh8NWGvdGK6YXoZ0cdtqP9uLmbn2zN6pcjUMzOb0kzxW7btdZuAwILy2TSR
6l3AfCG0c3ESuyWIRvgcol2xCW9jpn7/P+Rz54FK0mleRHCKQ0ipnI22dw9n2gwztcXGbtwUxiyt
PCwZEhHd45ADhYc+E26DaG0/LMvMJBccegz2McQijcco5pHsX7UhHdxxvRuFWiYZfGfiXVRJbiw5
Xw3A9cAkSFjePtwahChyNBUXofE553uZZoBwRlSPFVl4VgwFFxfoWlzPMHJ0Ui0TqbYPesoLmk5t
GDReLi/RBrJuVEK2y+Q0wvFlh5DtIA8r0q4O6NmRFaICBD5Pvt45mdBjHyll5JOFFvvcXrgFnbqq
4F0w8j4NKEfnDW0Dp/IpNVMkL/Lhz2aBAqFBS7Vlb434IaACheHVi+I2AurYj6mg0oBVJi2AMNT/
yeyzfXPNtj7uR0qO9ymzYrUqasWDUtG+grlbrzcWl3xFJveYSmrijUqn29dalaoIOo/Rhn7vwn5B
7ugb+390fg0nP38DBUlGB6sF91M7gsEmBfjxJKXm3WrqQRHUw+LDP9DDRYlrfyJQNDrcKTEo+prg
W9kzHnIr2BLCdtSJ7yhvPQZz71swFg3r7zC2PnfEBGmmfx/CtNR+EkROKVKTtW46Jp0fBzhvf+fl
s4SMElPDZOunLxlR1ysbuHBfroH0Unsu+vfBOAE8VYRMPRCVE76bTilEIlBUWGaR+Feauvv/iF8g
vAypg30efGC5Aq5/8Tl5Lf5mOaJgnL5vkENiYRXEG5wX78NhMgz4cZMNlZFClcteW5aoNfFD0jgX
P1Zw4fV/z0GDd6DH5euw60UsjLBLIN4JJ7f0IH71qE2PTqCx5Tub+eWw9SZIN6GqNo3lZBrRHsGv
7vx4uPSnGdHenoYfyfrodmLhJATcLIPnV9gMJSbGafcA4PQtbCWbrF0Fb+M1K6nCUBdR26orhoHI
dwDl3+bL16boNKodRMjlLMwXZraIJomya5B/XpDguWDQXAxQCFbp2/yggeBBLJxl5nyoOHDmZoKV
/uFb+k0rK+hIDKk9Im9HdAusmZivTrvzensA+8Vdy4NlpzPOxbi34MdWzrzxoSzSCb8u8nlBDOz0
NpB8mM+X9M0+CRvi6wEdiFEGEnHv1g6jNc+FXlQy81o/muU4bBL1V/VPSG5R0Xno0KJj6/Z1e1Hb
dBhKfcTF/u5xCDOVBorgdH/ZbzrUA2PvoJY/DxG4J0sqWUMDr3WSuEb1iLbT4fpuZk+sXUcQsBHb
t5bHPdpvCWlGyR92RmXlScEv4BPZcgm+MFFgM2XI02kZKj23VF4MoT6OW0Z0dLdkdcykOFJy6aix
d+RXfHEzaSynRxcIeX0Kzg5x1TLfVM7S4qZtP74+xPHm6sbCfoxEVwNMkNbZZXJMRt4+PGopsSax
7hkSdhRuVsFDny+FvI1wxfTripkaGUTfgXweYnGdtS5MDvddDjb9uMIZHUxjoTO80ca8Vyhyh0Et
6WpzFBS3TlEzzaICjSo/x614FpAIlWFh52L+YwdAOKJ8dGjHk7jCM4ANs6Qa/yIY8jQjaeOEAb+1
j2IZvDkF2de3gpvGBqcEtuVewakIWKR6AO13c2CcW33hqFLex/buAPP/1tPhgAzk/8AxK+nXz4fs
Ar0xiE1upxHnmqwux8S8xmk3sQ31pkIKOtVuFZEpYRDdfIes5DTesXEiPUeZFtHaxn4drpe81oQt
c4/1Tvu8O63bX72YpiwJ+RyLbghhXWUEqZDL6HOM5KAn761e+yIMtoDHyJl6/rqP7r6h8hBScyoB
CaT5VrDfDfKMSlmqhoKIZiTC7bqCyxQyfWMTChwlHmjHTPDW2VHkbon08wLtSRUmD0ZJsGZFpdKq
CJe9H0P6tnpX7tWdI01ie8mkODCJhVkpGkamlOFyWrZLe1LGOC7UvvNBZj0z8TQtvsEGYvXXjB24
LjW+eNZUzzVk0eOytkpjmF+3+8NyYHTAyW0uXrNY/r1fU1binJQVVwbysMNKOhJq2DVRBaGKuSNW
+9MzCakmaKQ5Qtyay0tYu16DGixQABZ9ueOD3Nc8JJ4Zmmr0U3pcxa7SPwvulAzTy6ipM8mJ2uBT
rEcodhOOxcOgN0JGd4w7jfIbMUgsf8OhcSIhlwVGLeQyamNUUZx8b3rdcq2FrkPWaneQqS/yI19H
Ja7EDuN8G6+08yRLJ1wdiETnYz6KNjrCg2kqNYwT/Vz/FSXmtEFPsdh60LWxL5g6yD11rHViqgAx
dhzOrPC3sjGIu3pf/tjRQ7zHDIZEpnM/aURg3YNrsggDAodhRfvgmLePHR4OGTyoig4QUwlBKbgR
Xncxq1TXu0Vw7Ld9sGrb+pf78bdLl+CFOE+nNdD9Dw+qbZVSvpTe7pQdELgErm3zJGDYWsDtAWI7
AHhoPTBtnSt/d8PX7bZjGSjipW4x6DAgBM3Xq2FmYwkKkoA6dTdlLsRlr16bLM73NK7qcM8SaD31
8YzUcn28W1MUdUCByD6hjs16HhBl+KZ6G3dF6X+8fxUGgL5Js/EMMSrYLgNLtCk1FPVOOEYu9ijj
oyu7zM8UnWqYxegJrdxa82tgw7XFmvs/0Btv8pRbPBsXdUzgeT3+yn7/on3TUoV2rAMWOGJMjJf3
fZkuIR7Kr4DY2UfOSVpeuCD3y9xRJussN15lU+R2jAv6TTumMyaf9flDPAUU8Ha9W+yeDFbmY7fl
rYx6RJ0anVOgFG2jrys09dF5hDnXpuaHDWHZz6Mo+HIU7SnrrYFF0PjkevWPpfCITQw4zX5FF4Lu
EjIuPYP/tVHkr+tgTP4FamkZbMRMFfGGVCxaPeMQr2ETQLBbTgyhZiIIXiNE4y6SeMUYXO6UfEyS
p4LO1pAElOsHluDqDf5+bdg9z+nRef5J8Trs++0tx7py6fW9C4bEpZNkCN9itUw+m3V7mrpCTu83
z+nTyUbTyYWRgQzHjHpUO7mkqFw54+QF3W7vaVJKQPvwIXWAIi++hziVHnvdRLJEb6yI7QU0yf3R
bxEDiqmV9aHHdX4Fp03VK4upvY/O2sd7ca1A264V+OPfYa/CQZ9GO6BwvejvNuro6Nxpd1aBDBu5
WjPvvBC9eWOaoTJM8OOK+7B84yVmcKRLSPb7xo66hpqQioPfCgi90MLPjuK54P8qoNHPoRRlof/1
w5zDFkLs4Zw+54AT/5uecU4UDuBuwj7jkBHwOSbji5poj6TQ8TfhYH8UHUlBxPxkRowqmicdpI9c
pHSh8mq923Kt7WA2aWL+UD368wG/SZa+Z0bNVEhdKvHgunapfXpGslU5Wvv/x0C87nGGiuSzPmbj
CZDSTuBha4uV8J59AL9hnkggPCf10rd2mQ9H6qa5LupcZU2oI6CwEumOP19uV56q/+agBAm81zDW
+YhPG4te8dgj4bsA959LGmmBahCMeaKJ+48Wk00xgkJ1upgjll4MKBpwaQUav3rh5zSRJugqAWZ2
qwknJSSobMrunITCfFC6+qtTO8oc0ygUgd1P/oL73LzgHdOdaBHL3/t64NGwWJZp108H347GcHeq
kC08JjwEjN11AVLiL79p0Ffh6SG1k3fBUCbbRdLZBBsCLFBdPj6zyvjL94GN7W+qujLJYDxTYjbU
hPVfS96xsfy+h0rEfR88PsgYLyFBpQNJDV4XTGU5DepFQ4nU5WxpCL9PTETQcHKh6EV8HhcCABUI
B/bePEtv+islwholCTcBl2pnni7s8lJDqtCddY0mC10SuAxPkJ4fMj3IKO6SVWGld7W7BWPpgVtC
g9I1HLRTnZvXB6OSx453R5Nl+sY4AsVU4NPOqk71BqY35Nqqp4w6L3yy5r5FfGVIXLJLJueM4spK
fLfsDkjsfBLhoAVCVAKd65HMqF4jVfXi0e0zb/PXaPm4m75bLIdJhjPd5UvuShY2yfsW0hjXlbpU
CwxSBka3txQR6KfdHdI9OB2173zL3WV4U0ZPpk4eZ+YAxM0Wl3KC+WacFWGe8WZjbgKoTPEgbrs4
bZRsXOG/v0R1aAFeNi4836DFlDOD+s0RdeRUyXv/8XJNWc1mXqegZoOnYTFLNxFd0/nfHva1doqM
9w/cWat0Il4hUKF0213ZpHLgFc22P5vc5x7t1i0Nsi4n5iTp8vjtA7xSpBdn0AZmTyZZSOPYBsVn
cuVc7f0TrfZqdAAWjquYRZg9kM21tGmr9qHJUTKbhmU28EFEDGixYn5I06OrG3sBrCSYj4kp8Zb4
PRbTn776I8op460u2BZElmKk92p41RFSXDnZOzaxQpb/ZUSylHvVxeuF5oHLvtgInxKOpPrEgDwL
HKYw3f+ApXIbv3H4eQhgh1NmcfUXQGO4aF26jSirqAtOB8+IpZQa2U8bfAedYWqPMeRe6pmMr1rl
3GNt6jkD8bejC0E4DMhExG6Batgl+tb4jhrPWZvSi6ZgePb4zGLj3JbgeN4i7iErDB04Dm6trXXs
Gf3KYVaBEiMkMZt5OtKQP40BiEuCoqWd+sBAqYfrpId0I6JR6AyzoCTaUsWzCLMeqCyVJD8VUEED
yAoibE6WvX/uI4IhPFXo+UH7xa1fGwoX9rn7Zj0/49QEKNoUxiqDKNgyPpdojioSz1t9ql9iei4U
7uN0RpQphD4xtR2lRUUtXUUdP9DaavVkVieLzp7pZ0A7SgEM7oYkoQ45oCeys7V7BtC2MEZOgazn
pUzlOppa9zJ1E9zEoP76HzNy7vaV1IOynbUXH7POwyhnDJ/+sjTuWy/TZrFn2GruezN8vBwrariR
Z3EIr3KYey8n1KWfmVqRMkwflDdeJSE5fjGBOZeq+Cg7k7ezmvd+wy+ldnLlN8mW+GPvqFcfe1YX
VQcYiN7jbZuhj+0Pql++z4QR0v9216nWABVPgiulzIA+p0B/fpQbjnprr+6MYrqADHHfL8a2aI96
hifXbE5Nffe2ye38fISyO1wub9X2C/WCOddIh0T3gj8oG/tVCu7PYuznrKbkL4SwFwk7epBWKazR
/4sEJS0kt6r/eImTUZziX42sE1MdqZ174Q4pfxyd5r8y/x2q2BlMcwQXYG0SuHiNaLn0A+D1XHGg
dPOHR9fXKae4zb24mv/0eDfMdesahxTxyO+jtjtkE8eTXDF6ulfZiAOyJUCrcWwCX++k/+BKzGRg
/aOiHsyloG49N7whR7X0D5Okofsam9Rcc2mxjOzrRXZptwORWlsV4T3NZjyZfPr7kvI0obmuZnTF
owCk+6W3htv0Z+YE+blkZCZLFO9L32GIquyBDKhQ7B+EUs7fHfCweyTwEZKKmtCa2LXHnJHSNdkV
6jAKjcIM6XzVO4jk0K2xZO92cF24yrrWV+dbHlNZO8rdaczLl+X4ZRQaAdW/cpMjykfufsP2JJJt
R4r9Z2PdOE6ym1jUXsmvjY8+um3MY1KJb9dWRtQ0GUDs0rRzDx3pwX139vq4cuVNPaGqndgstkkI
LdlLTVjpndhkyPXO19n/kWi6ke2qvRP/gLjgG9OWV2OiaYDIhgwmAbPEy7YbKnYndjc5vM2H3IPf
Jv4U9mxIM2n/xYtKOTVZG95Ghoeqb0SDF9kM5wFVQevChQPjP3l1RmAhkXgzffzbkRClSE5i2DVU
0/QStArZLkv3XpfoOrfoZCmzICqmPjzSkx2a14/U1hIOz4PdUmccq9y2btjJvE2nUuzmfBX1H62Z
U/af4REr4N5pRJPhS6kXCejrsrhLoQx0A6e0FLjIOEgviN4YUY88p6tvVR3PKH0wDIPdcB9CCETa
Zn137a4TWzlrWLnQJNlvVahJCLKc2i+a5AcwnKNONczgRuGvVo41AgFDlxDQfREVZUvSn0S5g4nr
kvGkJHMYz7/xFdrMi20AQlBkA57hPsm5lvigOMqLhpWSRkEg5MzCVE0YpU/zf6j2kJNZJEkkSXcW
sDuUEmog7NhPi+NQiUfE/BKAXJudFoEJsKRE0/n2o9xYX/v6/lBiXfQgU5pymOy4qat+bgshIDJu
FPXZ/+xKJVRYiFBN9mECbMDrpWXipwRICLJgnvFs6AIEoCzHmY5Myp0Ts5CbgEJBYu70bwDT+aG6
wZZk0NTDci6FVrb8ULqXhoDYs9tXnel7ACvw5gAZPoPuoU1WGAZZId0VcGyU8M5wMtfctUmazk0J
U/5AePUwe6/T0wnzGwAFv+JKIsP7EWacBPtE1nqQAvcHO6M1JJIwNB35h1hLmqVu3s7c34RPFmdr
1z6ZRfCkH++143WDe3JVPMGbTXlCgS9kTNyvWax6+lRl0yrxvBbbBSQYpt1RoTW7SMkDNONz1WgI
2/L3JypHlQfaVO9yJCQRlHJD5XEjkYftAlBufNvnYnCp+lKdOFuS23neSoEoXN5Rjge8vCEH/jo8
SJtN8Zc+sfx/P3+l9f3JCuCpam6b5LSfk6rQkk9pyp0tSIc+YqSKpm2Sm5NE9GBfPNGKcp6M2Tt5
YEk+BJaCVLaK1/C1SXOi3bD4fTvwF8dB1tRhykyLiS2bE/SD5hP4agFVirVZdWIsuyXSkDRNmGtZ
Wc2zMnTuSydPKcnh+FGMA9yFwTYb17eyk9vNfobQXohPcTJOgLgVp/G9w8GEfdveQbpG+AqFB5jk
Jd0TTfJFxqWd3lbWuAQsKxQqXVawU1aseyK3ZZFDqq8hUh/vArvMAz4fzNau0Pr1W9qComitOfGw
MCmP1EC1aCx8QRnYSwt0WMEbG9slh6HIyHin7NuJ17HyAlq2FZFgHrqTV8HkIJm+dHXZDCQob6fZ
i3nJaYkQvV6e/oJY04bNK791KZjCU1VAb57zwCg01K/c+zor5v1ceKA0rhcAvewmksnDDAeSjaB+
R1TSpeeLfYwSuYZLClSj8WxmVUVCpyz0zr4NrWcnlGKUyqf670bTHUSzwpPEO3SRVUVRX0fkCCNc
zcN9Msqjk8PYktFP42bFokd0dhQF4snIuPJISLexmjjzb8vo8AsDL19qpv3nRHfDE+bPyQNnSxbN
EI/UiUZvCl105URGbG7KeTAOlk4qD4eKJ0MhqPxxhhSEHO4Nqhw5RL9TQmQpISTshCJ6kPPj2bTj
2Yrz8RUv55buK13mXFRQS8pz2DpF5i0chDVd3bZB43XTxXnRGZBPyqmGIh+IwxUqyCCk6AICNWZV
EUu1s/e9SA8Qpbwgy2w2ixmCUbBeoDiX4tCcSYL1coPdqP9ZddKDWJbllgynOiZHJ8VrwWf2JN6z
wmH8LyCPYBUqlDiEHwDzoTKbcSJ9zN9fkHxgXWjJtAC+la/1jtQ/cQ15T3wmvpZlactsBRNCrLL/
WRaMU3kfaGmtzCI9V4BIEuljxa7NYNCJeaRnZvP86EBzwCNkFuA4r3gwhZcbKnSiTWEHfIVUXzpR
ji6m2bY2Wb862BnT+v71pwDEQN1TH+zfpO9WD17rEKHS9vAjo9FTwxM8La5w9Dt+WblJJry99fd8
BfoqHfwCN5ZyKhgoAV0P1iVVl9/oJYOOd7PH7vl5jASMBuZGHDYAgrPjCO+K8UR3bLDl+VMej15w
Onc6h4zHMxAdLfmcp6ofUQCvaqzkMICl2ASSjaO4vJY38Bk9yQoAZz6QSx7JQBmopq/OR8oKArCa
RXHhM9WpkPfK4vMRBZho8eeFx+9M0JrsjqTEv9BkzRS8YvtUQ1GBKela757PcWjlqatU8YcO/nPv
NNleMxshte+9ovCh0ZsSy/i33EsPFlYB/akOHvwBa/t/QjD0zOn+brhn2NMiluVHiVAMSpipP4ze
KEoLz2NLnuAiQ2NE32Jjgc/hADLFbYWM4iSc7qU0mhDthhiYlEHY+muHHtcZPa7AG/AXV9DbI562
zZbXRepMS9GyvYXx16xtehB9plNWsDGyscfMMqTFls2rwBucqjiIke/6pvrgKLFC7jKfAhi1J+/p
i5Yge47KnwoG6covv5v5AJpBUEp+oJA2r3J/0rnwpmzwGt2IDsbWrrdxRkuD2rsSrxQrjKr0u9MS
Hm5Hb2qCH78fbD0/GsxDvDMSXrp70yHM8xj4hG3vkJkyZk/svni5f7VGgFmfzU+lw3ayDsTvjE2q
GGg1wwjFXaWsjXNC+obPybB/gpYxDRV03FtJ8ax4Y4ksPWNLszEXgzbymclU1be71TzjJb5SugaG
W/UyDkX3Vym2cM3mB8ivt/AfvnbE3jYN8aUkJaXNK8B9v32doSihCHpHmODln6Qx78Dm05pW6lhs
bg/RpkZnbPNEEdmUbX6f7ayeH6LZl/2FH/tW07OUfNhh8Y8QBLt2wmSBqu2rf26Mk4I75CH4+VW5
rZ+86sc2OMhhw3MV4xS+WBeXjOk9BI1gJiZF0NWW9moZhg45l40GUGA1fOjdbaTP5G2KEDrQngxY
jFwUr3ay2m5R48GgF7+B7N+4mmqyP8PFy0o+FfORamI0QjSEgWEiftXOBXHWVFIffyyxos+jNooT
t9F0g41xhZxqoMDMYbnlltKplR/hpZ9tGGHcHsD0J6D4+GMe9E6tIbfg/j1WasX71lcPnzJQU2ww
lsgHOmZs3ShwKa+Wqnf3s6TCr1ER5EjbQCcWw76/QLTXAX+TFJHqGJ81k0GSZZOefmf3FmDID0SK
tWTiIQU+1r4oDG9UDvIP0lYX+wJQQP58uT60dol9z9T7nc6/AUwF86d5SvsKjPj61elwznjw26Vh
vS846udGLLuGHaBQl7ie+z1wVNrRuiiWVjCCBmsuGrrwJfIyN94EBq434ZEufs9bI31/q8ESdP8U
98zlG2ekQtGtHXHP948LpBUjUtiBQ3ahYRjmpp7YaDk7WtRfseLPKHv4QqOjYPcrAWM5YHN5cM/Q
VBM2dHCt3c0pcmW9OvKBvrUQjpC3BJZ2O2OuFsR98ocucHsnsIoysSk1aL8enr2aP2hsefBBpv1g
4hmmTnWiG6zsdFshEfBoh8ep1mPB0tbeBy9havscyLNYpPKwc1GpcXVCzkxXR9D8iZ+XiEI0kWap
YhtUv/tW69YC9ed0v6iFFjZm51fqANpz/WiYieh+OvlPoqWGCQLxSP+N1qUY/HMmUtKII6Fa2bPz
a5mvz4WsJMgkq+t5ae33pAxPjB1Wb1XU2me5X67Eg4AsT0bOH6EF3ztipaNG7OOKDZqt6i62Ppt0
bVWwdmB1sutjOXsXKdqMnsJYEqx1D7ipfnZsjVOON25t6eoo/Wj7O9AjLSXDsTw16DJiBVSA5Zxu
POsQXvUFc5sRuuYVnVg1XEwwUZydnTnCRtLoHG9mc6QJtSCNDCxbUbZjCoUQcAZpn6rKKYvlDbQC
SjFUcQncX5l9ULazjFE5fAU5TJLfzFmxNPDhqKQ7qlxi+jqqsj887IfaA/rwtpLuzAnCbRhsSo72
ShK5I2TSviA9sk8pVaPWJb2pkfxMTZC8C9cyu1LA0vQR+sNBwfcwPkFCaw0mohyPFcc8WdwfulcK
SXXxJJi6lk1GqjK/d1FkgSflzO36ri2kioXasShO681EQZ5tUdgWrRH2nCeqU3qQ/rr4pNWzBxQX
pt/tIsivyTrQpSGwqK4QARE4VaqpgnSnqE+MPnQEm/CuSD4OwotLu2AHfh0q5aY6eLdwVpJdCtzr
NNxsEQqAZp6bhceqBAmL5lzYIDFMkeT73svSOz9gAIzEeySFpV+zZHK/O0gEB5cSI+w0WoD6Xvc+
unvM9+nK1oEGefL+9zrKEtfojtpfBeSj1rV54gxZeDz6rMULz1ehhrXMpcgVWbtPC2HPdj4i6yEk
u4/I2lFeXax1qaBhPtTx6brNo7in6j528gQ4jKqD28iJmhfz8TxlFLdlKlZVf/2jEtZ/Hp5Ad8Mu
tzBq7fBqOJceN3Auu1kabeOAN94C5dAua36cjV8aoQAP/Bx17lhqE+KXWvSpYiESOa8wGxohfo7p
YAJrOqrTINgHFBj4VVM5nQqbF0GNJ7CfJIkTpqVhZXeGWRG5nnm2CHLsPYk/5rIjg0DGKMo25bAB
T2TtHjMoKHu6ftnn2KjJ+fBMfp2kAB1qgHZT03sKEIxCAnRE+p5ZZxtyFFh1h6i/OIuTd9YL0OwM
Jv0Gl+iAmU7rkHtWnfvfE0IRvBozTbMjjH8lke3DL904MyeKoRRhCCiRNFdbI1/OxMxs4ZBI4/NW
QSbjsSaNki9vPMUsIK4JWAZhaJcJbQZCRucWvOdjsMB0SYRDU+EaNRDOgo4HxAm2E6IaRD+/3JIr
HwojT8leJwhqL5LJuMtB3o7zB395piFCma+dYp/+04ou3CcSVos9uOgkoFRNKTkRUuPlrvjcTAEE
aP/z9Ly/b/iRCNEdrMHa+nCaOWldfvJY5Lmo05cA3pgelXTIfjBkckqd706NrGvdW3IkIik6DQ0/
ULvrud5QuRyto/9hmfC3yU9oIDpwCQ5gcY3J2PfQbYzGtE7beXngCrpqXGejYrg5zTq22YYE34BR
QMioiynuDwBRsgxOjETM4YpHsS8BqzDba8G+YHMlyJYONp1QXLHIJNn20B+0+kWW9tga8vimnzS7
3p6FA9nG7UdL/FMxAAw3lx9ShcameeuOCEy6SHWPPwT7In/RShIeHqmvZCA35G7yDM6+hpUFqCS9
u8BnWzh0DbXRszOQropYW3fEYZtdrqYl3VgHMULezrBpxzjRnCGO9sybPwvO3dL6V8D+P8YTLyKo
PHeeeDt+XUejnfH4PwcgM3KR/tQVbEtjtqgvNbPqsKjsn5kyi5UdPFKCzwuQR7DtlE9x2UPnQ+Zb
pHoJRTmFWVfLWiZZ9IQUM8WdA5Ve5MoTD+m8G0s/JO/7V640WjkdSLGbYTUmJKdgsdcF8cYbKzaG
/f/fJ5iLL0cSsoyo8PAeA6+jnugmbep2NAJgwszbu8FZMON2lkxaDl6HIj1x3ORb5fszDJdyf0TH
ksxxrqRYPW9k81iYUTfRwRULOCQLQwIO0ZoRRbc+JoM219rboQKN4tjsF0uHISAG+xamTZCy6qeJ
Ufoc5xW/IDLDwkAQnOFdBO1JSAtbWJCLEpdIjWZdR0954vwmysaXgY5OtXPNYsM+Ndpi5xRO7x2O
6cALgWbFXQDZDWmJZtYQjTHu4KQS5Mgo6ltlLViTuhFdSzS4oYGDWUhQuSLrUZkUIR0xeuH92+bv
NjxTXKbjVFahXpV/7q6FHecMc0C/i8hSh6P7xDfzoXH3Z5DFUoIWJ28rizoEEf7p/81/JVlBMtbH
ccUzzHi6tvGKfxJCx28PRH/rV3gBxLthH88yuEiVYJp1tejBMew/LAcZd9/6apE6xL7s/nTF9lli
DpftiPUcbQBpV+Em6Pndks5vknFT4PnGVCyFqqMTGGplBP96BJ/Y84Dzg5EhGy6GxAaayXzvABoQ
Fh/Hhk5il8szMvC5itH430Ssi/6ZJu9GGLyrG+aQcFbLOfWyJkLYAQMBHkHJMYPMOE1+K01juV8G
CFi412+9FQg6fEUwpSoqtpHYxqPi8oyTOEnXRn6iOdfIP9Jo9IEWquFL8N3Nm6qrZmgp8Bcr1ZsS
AaiXejAA2LHDn/gSuemMrmxv6kzLKoOJf10hELZqrK92nd55lyRB0C9hfWwScVPcVsiMeqMF4T5H
61pRhtgW31eOTy5YRzosVFjqpMBPOBexIej5ppNiAgkRebFPkfzSl901rlwj3wg8ASSj/mKYLC2b
m1KwyggOpQOvr7yeQ2/Nz/lnoSjetEyUopdvGrD2JGhCG6Qe0jzoA0fnqrjijYKDf8dwRHdwAF9f
AG08YRieKhsH2/Lzf44YyfJ6shvtoBFBolPAs0RHsFVQSmtijMbDLoI9JZFyqWlBQ6B1r2f3Uziu
XDqh08ihmW54plpqzriwxahnnXyzZUwY2xq8jdm2sQ2lH7VbNrv2JiClkm1MYhnDbj87FG6RDft/
VGTqb2lisfKdU8PNIANeeBN9RF8ImtUz4HbvG7PZW8lL42UHViQxU622vE/7c6B3PHbObHtsH7gC
SDx46dNdnP3GRGQLOfRtLt1nqebF6yZmI2Mqwa3WOOYzbCPS3ZM7djANdENAPFaIF3RZ4skFm91A
dwHqb2eN7ORQ1ucLqL4xlSZTKTtKni6TVzxEJ7eRpcvkdHScR8J8xAMcgT9ngo60caXsftrzRDHz
8gRlnGSlzBTsjTxrHR8ev2TLyZEPMHr7TjvFINtea2Sh2FoI1/7baK7Aeb9lVjD9inO3ecms1i0c
gcg1AyXT+s5AlZ+s4ctevXcsC0H5mQY6OfktyZRSaK24mwVIKsGwddOClks/UAliqxuIaz52tucF
za291jkDydjfCQ+LS0GhAto5S7sfTOpCXtUyaZNaYzp2Mt7Lace218aqkYKuAAxgRyjYuEjA6w7H
zb30DtgkldK9mAqu1yyqLbMacUHGOv60noFx2DjXyWlAJWZBfbAkrA7bzDoGCHTs+RvRk/eJkHwl
T1Bfpq/GXt21i7xxa2Z9kgA4v87AMBDzJmd0tkd27zlWfEGHOAPJLvhOOQzTotfRNPVYl023oyNo
MzYu33khAMYJ2JgzNDbWxNpW/k4QFYvaeZwgnM1NlgmNLHOU4FYwRBaky8HzHKUxGdRslPZIXAQc
EcNJCeHQft7GC1hUMkDuNMkM9yauIlyHPUjkz2deOUttiWcZFYb1jhUbCqvzOz9+2QZMmiCeT84+
/kFC3VdqVcGxCDKXvGBSe8Od3bDGlRma+xUUXdaMvUTpW1ajhf/dMEAdtMLoOMECYbbogIOpnSPd
EQAe1CzrjsEterfpM5o/3G4Too5ukSS+452/73A/8T3PX1qawmmTV+qtOgdDYct6FGGYTdoIRLhF
U2wL5jyOAonKwZ3hO3l5JloLpGJlJ3ARlUXv892zxml1cE0+0/KWKpAzoSY6ChU1tFvOA6UBB6Tt
BUFDyzy4EIG36JKvBlLFoUdyLQUpc0yC24CH4ZacOmnZ179TYq17yzTYA0aouZnki4SJmTEmWjw7
4j9xTa4NZkeevE3/t5kSf4tLgyg1I+l0rubaRdo8ZLlj16CxXPAqbBk96mG39wwJ0v/dkHS5OCkU
JpHr9KSjmjwXjgPFPp6OplK45mY07Eu4vIsCu19qudqXEJEjylVpPac2bcFIyaregv9TkTAMzSIj
UToJPwWgvCgCwwgjYlcW8Wo49MkIfmIbDMn2s625dohhPQexIT6dfqxXWWg759YwBKJtaHFyrQBS
QC+CrHsoz6nMI26623RRoeu0HRgxHFOVJ1lY8WMauVZTYijZJ0pWN0Yafn/sDzVMhC0jV/+V6xyp
sL8hZYgiKKqSwNU5EBgLH2R9HV98O0yC+RbvQ+IEQe8sAV6eeZwXiIsqegh3B22yjIFXSVKNMrRd
RHM/BFCQTSs5FW/NmrvW/gVDsic8S/Q3RudVg/64e9OJ/cnYVayKv6obkayISyH3+C4YxeyjKa8O
dOzIAQvZADGygb7LyB5n6s567WJBb4gAPQS48o8O9XjZgRCwUU2AQ2rCBcvWSmdX3HKCudyx82Km
T7S5dWmFImofnvhOfnhcopKI/19pwN7p+NNf1W8EGRsqpKfHwGbJSJUMjH7nIXqpbejiOv26JlNP
QtcD/RFe9BbK6ipYg4JjSfrELu8wJiprxpP9BFqv22Way3G9w+tlnlZpFs2c8vQNHh5M9VJCDuA7
T77kQZ0mTto3cHb1p0gcdVI57Fns9b70d6tTXE3W8oSx1ydS8FDd5xjRFHdDGColAh2JGk5K7qPC
VuMbSWDRcJq5ADYZ5RI8zmcs7P/VndKSa04WAyHQswqR3IZ3BJ+qOWlYsyI0DsNEgSND1786Ldkb
d67faEN7MyQ9b8/07ZIbjXel7Jj/SLPNnzmOUyD+5WHd6+zyGDhrD+DOq9eUdbHlVZIs3WnSXPZR
PckBCkXaPFWhF5j3tgFGGRcOjHJl1n8/wUMmewvEJdc5njm9NLtxA51gpJlrqvNQZ+l+30RQWJwU
bNaQYZ2psDGZWxEtmfqwdm13ai4BSd1lqr7GoU1tqlby61lPglJ2z77hNboxZOKnLENz8txeO1oa
NG2IFWXhuhV454KfZBPJneDpjC7bn/ClI03hapXF18hA37ZV0htErn88deCzl0ajGPHk+37futvY
6QR7o7hJ5O/mdqZgCtJ64rk9TJEidBgsbBdybMPViFp6DJOyYmo2trIWY4o39VoKsKQ60yEAttEO
yRwwHJ6fjj4o5DSJsewvPE1vX+iGhccsQEllRxO33b2blKFN/zatGnRgKv1FkTfLmr/shvPu//Ec
6BVhChvLudZKJQuecD460xc4ydMzDqcljXswEcIQuck3QSNwRDDtQsoZZ0xYqwWqNtWWQETOZfMJ
V38Oaj9QzAnQPU8VPlhOpFqb/QcY2bNhhuxuKrW16egWb/2r6CQPLgby9bUosOidyBBkz6/CzBh4
vqVtDKHzE8cU/1WkCAXbnZQy7ySTCoTp3ldpg5smBoGIYiv9ms/DJjHaTYmczelFRo8wMA50bp8+
gbAOfXRZxdtMOdteWQyFY2gJ8FfcfLpWVCx7U3q1FqIabqIM0kQJhfjdgpueRvg9Uq4ngtQdEpS6
e8XdvBo4o7oH+AiLazc7JGRl8V+CKTITUS64XjOC5SyQdO9DdsrELft/HPqPqrgVgiV6cxE2mBgo
+aBHFkKQWwir7sc3pmH08ej0JwFrETVzIzojFW9l23lCbrWrMtVYPvqCS3+CHItKamVOoYwb0cnI
95Ymu2KiDCSSbPsDqH5S6pVnO/CVKGGYCD8NEXh0imRXM6WZ3U1mByeMz42PM3LLsBKp6LPeena/
txRoPNSNeZJcyUvl5qFf6KKTKMUUJtDZG62pr2UkXzWOSmaBVm7TINdijhqdMTvO2J/bka1LfO8J
EeZouk9bjOkmkONznlp/CnvayZ3sVpUtd/gE1jfybrK6YpnTMj5gGk6P9FQM+ZmZTWUES2P2sde2
jZenFhSVUJgMnXRz2U+kf56hyS0KdC7AdxC/knOikE5lkuhYUzaWnt/nt8AlRD3eGGTwY6ngzn/y
sUaxAuEo0FDB+OW+hQpIabIneDsiP82LM3fiGG59lic5iowifXqkKRRHr/+C3KcFlXXXNR8eYeVJ
TS2qqt0eKtyr9Isw0W9uuHuRsa2/OdBUN4mbtZPlGrBkoGKFB47kPcstDAajE42NumdU+9Xtx/dg
2/cAclk6vjKWWKl3NISc6dXHpHIQviIdhj7iWI+/nZpFxCbTkFqINXzjaEIlBjqDwkEVXq0wrdtC
dGsqUbfTFJrxM3UYgunuJXBuLjJsB2xyWvwAl/2VRYI95gL9syWsbSmcLJklPKs6evAQNw6dzhtV
RZ7lQqUZofYHekfKWLy5ZFE5Aq6RoRjU7E4BFfAmLhBBkdFUhNbAhmwwZV0vGerV77tNI1aEarOS
TgvknkYXjih/tR1dR12LeUJ0uHfm9CGipK8+fUBgcFbQkNOud0iqV8YepWOoPtP1aVYckVqBHTZj
qZhPZ4BKGGwZ+gviGCUs7CGEkaRIoaYX2zpV2n9AdGRankcvQZ3ssU0XiAd5Q+K415kYK3QQdCzq
726GdnuhkxzS70mt7pb3CCp7ySfnJym1arvrML7hsG7gG4nTqrs2iPz+Dr8gniMgwC/86W014d+s
3CYMBDJOQCZR4RNDVYTzmXuBRMFx/vTSiHMsT8SK0TT3H80rX405OGnRj9dvevoSwvtVmSMlNBw5
rvzjHp46gAQU21dpFLPJV5T7GOophVCkEaAu8Y00oZKsypIlMM0r7RdOHS2+bbpANFeWYvj7qJxi
XIgBVPr06SUAd9oLINy4Gtno727/MJoO4DMDmIpdHAauZ7FzzrNMxwN4PUg4ZhhX0Q0X8ahPax2c
rXjsyQsu4b2gTV/JJ7oEodDrttWAWQPI9WqQd8dQghmB/OdH8ufxtWpmUpdULnfpIlnvjKyhT1DY
7L9VEHP5FWkR4xPZEHYTDKDSe7VtJUu2JCANM7lp14eRU9zsd6lkvLvLoE3WT4hST/dBoiEkaIp+
TeoSHgk8sUwHCkg8WMug3isxDbHNTwHQJ7ZxbfMYseN81INs4Rf382TW/nRfy7K5yoSTpSZYSLN7
7vpXn2luWWi7UgOb0/vGi6fOnvyff37YeAU0ffxMmSRvnpGvYfLqE/y7JnMA1PAhSzbfD6ey35Py
dtRhKwEwVV3TUSMWoVxTCxl1PAR11cvqUm3Jg9MA/qsBjY45VT48KXoTWes6zYNBkZDfCq2qfIe5
b5MDqR10qxa0olNDTBVFlkyLJ9CUujKkVwkwNGbIPasDD8fPShMoDQBW5wLws+LJgf6YvX9vPxVB
t8C69c7idtOk6eBtWYva4JbgBS1E5RdK+ZyWBL889OeZQcICqo/5aqHV+GUrJpmG2JozcpkUbHBz
hh+KIaTvOdu1ToiawI103c2XWET+GtKJRLnE7hwwetYohgWJVjP/MHSAtIpe5Y5r/E3ZVWmxdYF+
Hx68uNnXzGeEbmXH25RbKzLqmdK7Umt6TgZo+2ijRlH+FLGK/T29N2nZFPqemIJKAiuqUU0nMJ+I
2WA7QwNXVxgrrLED3vq4OEFL5cS+OZgIibs4J+5eY3dEuzQLGf8G1Y9TV4AHj3aOiOW2Mnyma2zP
ezc4wP9HpvmYCYwt0ZvE2UVTPI1qsqahQla09C1y6EtBwZuUQZk4pOugXhyQRHUQ3La3YKw319tL
9am32lDpRsvv7lNeb+aijU9aSXK84UeX64xbCQXx6qi6JxK+acO5nXuvFrxgfG4S0M8VuBxUZmXu
/XxvqcnCFRtFSGBqkozyhw5y0nTloCJ3+bVmfbAYFHrs+mURsJCBharFkK48s8m5KiChfGHga0rv
mhhIJWlZsdNxh/nd35KqklGMOupVd4j6rUva6iswHN2IxV+C9UYaykrpfzajyahU62YOEqKR+FZW
+NAGWAjaRE/HkpHFGGBtL9Tb4U+X2Xv442tAU/fDM85EJvco2Pfpn4QwBSdlG4Ax09TrjQ0MyGN6
3nLOhVnG4R4OmgOLfXqW167eP9F7EbNPrSoH1faFsjUI+UmBHu4LNfK27W8c+0vQ0c0OszvOEatn
j593Vhp8+g3LUH60bfbiqM/7cSXijh8dbTsKGqeJjZb1r7xcpbMqz1/Y+EiskAGwbJP/Owx9u0tK
B0jqKzPkY+j8ohzmI5OitSR8W85g6ZswgKPe/v4bxgsq1lmU0v7VeRE2RIIxk1jXIVWehDX61l32
of202pa1RFNFOGHJpIpCQk4NyYTkulZbbrx/k7xSUWp8ery4vjkP7ZusBwTHU9O0I9tiEUgyhQgc
VldjSGWB/9lyTgrbYOiDms/MoU9TZaoZ+gZ8I729yPOjotSktSnOI+BsZWFPyGb8jTwYini7pNhN
iUUfHzgIm1bphAaDezVfXNRw6MAYGAaTiyDn81Tty0dgN+Eyc4O4NZNRBUG5QxWEo6EkDShkTiZh
HD+L5ozhCyS6W5vjSNzpNHXJwXrYOf5mvvS/vJRmhNjl6VJoOCFuFEVsfYoVeEdVGaalTCRoq/00
o/WYcblyySKH48SxCzt6dqKuefGeQ8Vs6QSYmV4Oy+UkqjhRfyDUVh1Q6pmARieP2Kh7JpIwmIOL
/XchN1Z5+cMNUiC5f+P4OOEP119eM0VnxldF8EsStY9ow2R9FKojaOYY4xvXfQOmxVtT0OUjqyEu
oD6zdyrVwOb6lU+J20rnODrjESr/UKZKQNvuYHIFMIluSV9fSVTCrslIYjrrtPtmUqil7AAvxebn
Ml8SCqT/CWbNJkZ7bSadr0Yx/guVzzbv7Ik4EkVYzuODW2NXhtmOGXVq7B0D9Upimxar43AuJhQq
wAiw1xPI0HxuOzfvXZUV9gES+PEBodo5ojgX5vtG/jR8SnT0zN6VBs8tuk0XqhDSIXxAt+YtJHL+
eOMSER0bBydTEJVwzH61MGTqFoo4cKvLn4QMpBS0slHbwa+g1FaedWKftEe6QkkBhbyIukRj1GRY
oullj0euBJPBmMM3BtYZOhilYPS6wNaXIpQJWuReP8GIgGGP93kikdvQmZ9LQhkRGy9byqWl3ayy
plqMys6JQztAd0fk/ddgQ9od67nSq75G4cJDtoJTarz4a7+4c79sRiNorkEBoHJy5gFv6qkplgYW
u9SWiPtwFgfgGup16DOxtcLX9/7eOITpa2K9fCZEILCCjp+ysZjWgEQgqfHkewFIuy3GqpOvIS0f
bLWdDlABy++7UgcHNU5EpkuAKZv3uF+8TndqnVxRj/Lsx8N84ZMueqSCh010g4tt58tsSVIp3KEB
FpU97Ddf9XQpv8cD0uosW8TOHHy/rr2E9Ee1OnDl3JaAL3UobYrUoAFKt8KjLtlihYSm4CpHgrbi
hI6M/s8n8/RO7pDWJSIhT35L39G8/nOKH2yrNrjfqT1nRzd+XPjqFNU7C5Wc7tdESB13YnnMQwNu
45T2wBl5aQE9piXKCP621ii5OpBkMmzonmn01Cn7E1t2Qf0Q5sUP+HR1Bw6F9e1Thb7PyoRJDZxE
T+SUCVzz8ugWi6gZZVPeA0O8ahRpE3SKAuAZnBnYo2TZeVDmRa/46MmXvUa33u0cimvw7BbOjBDG
/t0dhGVjpapiPJMLxEkOsgT+vBJ1ABjsPS5aEntac74hARH4haDt/CnLjWe7wWCUyJtag5Ly5zlE
WrqHjS/Y2QfI+dB4/hOAv1Rx2qQq3azjiSNdhqitscGavBqF2KuxMMJFsv+Hq2vT2DnNBBysbgFf
hOTVkFvsXifH8J8OkqjyiMlf0Oazozxu7Carg4eFn9SIgZVveYp9jOa9EKiNdb8gGnxTPQGPAZkR
x6aildoL5Oorxs+BcB3YXVik/dEp9qYA09DYCmAn+pttUqS1XOyJbv1bXDUBThxYDWVGNlf2FZgS
FjtnvNNQuUQTYZYNUffMEjYLBu8AmXqHY9aDv24OV8sWNJW64qzMZVAI9mmQOR7jH4Uc9XB0zton
Jfw5purF0CR8hi1OBvaBnp5Rg+kkN7pog0MzKRJE9h+cidEQ2cdoymXP2cHHdzvwY3IblH87D7Af
xbODcy6ri8x+LIziIemw1sj+dZkfURJwfNHVXhgDdihD6Uf9+Pb8oeJyioizzWYsJuhfXWmEsmFm
aw0Ak69d/OaVMEJa2l3FaHnrwS6ajlEnHfN97IQmPDNB+s8bX/1ft+OQ0N9V1QvML0nUQOzlR3nE
2L6SRqpX9aALH5WE0ETjGUZPwyX5DMdXwylST6VR2MvMzI533a8tgdb/WSdIxgJPHSYE0qlYpPrF
XfUSADN/k/Bd40z/VqFI9v+E7XlwZsEFc31ei1dA65AKnRv8C75bp4FPwI1JazxlTqiasLfN6lqm
mwMtCHSPk/g41J2XvkXM9c3usT0ZZvY9FYoDQYppBTnR7+hy2rDetNvbbvuiguK8h1sU9JGu64oL
3FO+tiZuNXLDzbUq1HGBDLvJUJslgmRVnZIewkUsv9Gy3OPPmLEEP22c+3deJvp6INI/qpUks1Eh
DSAVLgkFM/o5h3vxsFss2FQLtgG9kEpZxJHJJneyWey+OqphQJws/UnaZrQiKGqLPMCUKM2zkMdy
wWSA86hQfYej9Kxm3e/AMV/fb2EIanc1fD+VbdN9nIiIfCuzmEbvMTxNy70qWYeR4iGbI21kT4Ax
V3C66nzhs80hOlFBkZQncnBuLVJOYSERcRRIkde26EZmOkw3owDoWvN0DjbljA/lsHnBnHgqbrrJ
vJRXmnbpFWH6QOc6nZsJiAY5bAbdXEtE9LTm8MuRLYpEJ2yzHcAk6mY0h/kgL4TFtcHKeueabLDa
7cEHrXMaTGPke8Kq53M9QxIMuiXh1tFpZbwVZAuUeGTRKVqU6pCWMmy5I8p4/XQmTZStbO9jy6q7
rsyeFgWm2VJpTcba4lnGu1GVfjfwn/TRs+fLIiueqx/j76PjAsYDzRWIJHKLD2sNb7qBpd3mhyNh
WkwrQ7GyxEQnyhjzxM/yUB3w+QwQK362nCJ90+1bAbFR41wYQiEnFwAQslgg1H7O5utLv+8U51SJ
YVsNRGrXNfgVgPGaLt/R/h9AF6C4ExL37vtGa4EqcBl89yiPC7UHDipu4iNVnMt9IGwVcOP5pbg3
LRkQDT+XtTBlfoM19Z1qp+nnn6uuxwvq/XaHuIU0UWjHh6ESlurrcinB3WIetvh8xJ0wbKWkX91A
FKQ6ujohAbwCYIOcMH3h3jvoNf7io4b91PKlicCMFMKAn+5z2zmNcqOcQ13R74XxEPfYVtrZ/YuM
3wtNulRoWmoQQpgODUa8VfMdUJ3kq/1Bvxybg8vqv5Pn5mTwZzEvIW9yZQKa++Za4l9sWakc08+I
r8j4wd83eCEEFkHOt/xaSbN5lcESByUEDjYBv+hMDxbmgZ5VseghfR7cgdiJ1zUnZZ0yaNYryUB/
Nkt4eTdobiTvEgajIdRfNaKuHknb0VRhjwQioWChsqZKYruEAOlzMw2zP/CM68gZdupjgEgqP69N
A2nyqXO0YbAmQX/1Rp3STiSgN6QbaaKfwXCllFWm3RqRQ4sJIe1543odUgvYW/Ti75qWstemgn/a
qRD3aKRaftI5hrh+YOiuLwCGY/qve7O+8S1IFwVhF87qntS2h251hEUzpKypDKS3Vmjc1jbZ2Mfw
iHDjgNHlW8izshO1fVuH3X2g1BaQVBODQq3pxC6H01V0pXQgz87HPXcdcum6jVd+1VvBy/XA/QgF
VocuIu7Ba9uBDuOa5PIgtEHVKFyVnz5ACDZEDSjZDuaZF+izOUHkQ15bTqub+fCG0yHKTqdFNrE2
MUiQJjY225PVYJf+L5QY3h44a8BMLz2UQqlLceGWc6ROhQJfq8nCLjkcSomHZHCeyi1gt6EWzdln
70X6vQ4dhT0R3SJqEOwAjBPHdvxgPzp464WoQ3Zfv0jOBKkdNwCUpcNvgX14feMGrpAZHeeO5aX8
RlWm3e3aprnQFsqJkr/OHfdHeHDsZu4+RoyTjcnpVM8VRytXVu2xm13cfRduodp8mcAlffiHa59f
q/LS/v96uIYCZUktT+hdYDiBWPVAXK+DKnrvwsOIjt/Itu/YOD1dH5QJrWsqca7iDf/FaQEB0tTf
mx3DL9cpfLP/CEi6KkvGeeZpZkpde/XFjFj8UCkzMOmUUIim3uC5ZQjJZ/WyXfGTIv6hvYEGFZp8
jeLmQMCRPGlQ8AWDbOlvzSZM1+ZApAzC0uSTglwFOk+krDt5x4M+4Qpc+t97950T/crHXw1cPxpM
/wBsz6CXxlu+CfRmQG/u5BWz1kJG4wCz/fVDteQ38fsVkxi0FT5FGK/Gl2LgyavqpaojHWu2p+r+
wQQ8khEQCc1Vocpi07BvYKkzPH+reealbwTzLjVb6GK8hrl9S1mgsVPa7fkXSWdCVA6mcJ4Mu6rY
4PMlAYdXJJali6LV3xWW7lG/+h0u3z9nb5d8kYiGbz4zpQs5CfUQWYro2AuH2cj0S48liQA/Mn45
SMcPQ61nQSH3DThZih5fJnd+wTIWax8sQxVpVqmwRK3DcYE/hk98oXMT08z9X8RUm54Q7HUNYkcr
r53Nj/R5kP3uZweIxILEzwGwVI3+lFMZcdEH6cKkyOCdZ9pXmqIPU8BzZUsEy8kHhrWrZoth/pEX
2djLeiJGHvACQKlIbLLYvYrpphrEshbf+QUfegY1zb55t2PipDeHwV0R1Hmb3r+0VQgkLrfrOmHJ
Tqv4J9KNLrPfiwfbbXLsayoYtKZC7OTzfuGE+07Fgdlr0ju91DWsbSFtmP4MDIn7T9PhD10A1CSq
wbf4jec6UDr2fahA7qCPwwn4P5b9y3lfi0YR/bBoGveGenGPza0RFQOZ4KurSAVzl/U9qlVqlfFR
W6Sn0idD6Z5fLbGVmpPHab9ZNEFnFFxZzlNR+q4wsTdtbgeyjQ8p3pdYTcnJpPiNu+EynhBREdnG
URMW15XtehfqtrRflaYdWYy877wwfC+aLBJY7X1AIgqwk2apaPZGvyONiSOk70ZPPv4niCV/qBQZ
ypLKX5dhcG2mSosNtN7ftoAwchOFdvdJlJQt2q/Ay6i/gG9EVcAZYhp1RE15m12p4EPUf/rbPWZt
taD2oGgIE+3QXgvqdWjn93yHUb4mLIBnMSH44MdQorjqirvRvcM4nnvJYE6fEq96KvrUG9dlgZpR
NGDe0dkL0MSwH4kA6xLiff2s38XjZVY64aaRz9NBPt/Y8l5kmoJ1JJKKmhN+3iLoeH05ILNwa41B
uuSxQrD9uKnYXNLAejmaG/4MJ+RHq2rvvnDmyhS9mMHFtAT0RSRnNv2APmxXOp68wjOLEGJYsbNz
2LzGsjZGVCBxVcaXa21DdcUElnIRjlXE+VwblOq/DjZsp0zlGJO8ydfbHrzPVoiVVJkuDzP3C+E7
4FcQOESWRYzAiLrAFbVPsy95ewTOPuFKuqiQZsG6JPKIMgCwhrwAuCr2sIS+G4jJ1YvaVosywA16
05xoaRdKrnI5CrLRk5J23UxbfQS/yyqvlP0K8CndPeti/gaUtChQZBrsebzpsYVLEk1caJVj1BTH
yq9pP69thpsZTgqC+dyGukE/z4nd7TkPcWnaBUin4C1pW+eEteWXRkqkZAPeg2dSaO3X+eYX0PiN
oVmybzgPGKAd6s4f1UlmTmSczDcjw8Dw6neBvObT/Id5f3LoxcYNtGNvi8quV5gXM+UJ+YUFZfwZ
V3TAW5sfwxekIGrD5xaYq6Q3W0GLE5e9XEyaqLTfWGwv98mQmVKxn0T1aXSdkQcsqu6kAi2crwkL
Jo4Ujrw6o/ayWZlzj00x0jdUt3WqDDCTC6doQ/kKRe/13Kp825tLGygaSsEweyctxNYsK2EHAV7C
nMOiWUOdBDccz8HlkViRXBEphDpHAkAq5qzfbfWakSK10G3kyxSdvNwOQyIlaIertm/egZNDwO5r
ttz+LplP2IPu1dWxKZWvY4F2auXGK6oFDT64PxwdAK2WNzw/m1gahAIN6sQIhGJi6yjFTtbQS95N
3ggepJHlcqf35jBPHzV1kXA8ILgNjeY9hWkdkkUMD9RpYnb5A4BYpboNxbR4aZqbxotX/Mj5EPic
DGdYxE0PRnw3YnVRmKJ3U6XmOI1xtS7yVBDLhfsuK/0ISUwbfI9LeSASC1eORM+CX5CykcgyIRx+
3eET/IB+2o41auBgBFavp/nupp0rmrr+PSLPEjWn4DEdX+vSp5U1Entwr/lIEz+crZ1sMnJwXQzL
HMw0dHUnXnawCkLBNmFxUslRlv7L34npP8r85V/k+9RTGe6VkeadE+9AcfF930CWImjsZkOyF4gV
MIss4N1OVmuA8asTNSMCUKiIHztXw7VdReCHWFLN7+9EtYtCTzYNyifVa1pl/DpeHuFL0TMI1Qa8
z9nsf9n7mPaejlWC2mAqRTCEMjOLejpdDBVLqGedz4vzCFurlNz4JNFh46HbJ55TtjHzb5bcFgXP
zpRZIEkhny5Y6DV98Lk7r5sCEeGwmzppDk2zYg/0LWiqE/5axmQ15fcaHaVvHCwnS7pvKtDLexZ1
lCjTDvF61g4cKtiGH6Lskjahx3Rmov4fBz2GBGvfT6oz+rC2a/8sNmnvAh0NcaICXbjKr1+J/46D
txusPbSRu3ToyQdMGcb5C23gC2/hYmv1jGvKGVRnc6c98RkaikiSjp0KHc0e+Qow5OWi6kcRxR8+
E+S4vV/fgkfSSnIrDAYE8NdtPLJhV2uxT9JOp3zj5mlAuV78aZ2/wxxcY3oU4cu2vF2pA+7iy7dH
y+zs+/VoJUNO8BJtJS/HKuBvpU6U0oZ+lMx6ORVOOFNkL+XPKeRg6xJNI8RIGFvEVwao7qxw7CGs
62zQ9A9xwmrB4iLKK5eJhte1IYq+wllq6en5ur50rxVzQ9vPJnryd17yuHHFWRywMlC9NSnn0rs7
Wml8YL+SYcoKjTsJYRpEb2BELyPegwQs6OAcdRW22LFxEX2VBclcu6QHesF7sXA0tkw+cQwwBOcv
TS9kaeK5XHR4u7omMaxsvBytsZICCl+9BGIGwAmE8E43sCp/N+mvngugwIOWnlqIwaQQNR26r5v3
Ytk5/kRXmLOBBmD5O++YLQmGetWoJr2GSXdQmcBsF9Z50H+edQaZYKAgIBOnqmTKpiHIdbWzHnv1
xpoP1FITFWrM4DZE03dNkT/w55ce+Uj0yjq5ekFNVRrMP3r5WDbmnQ6mKeQgZ5nH+AUliunTnbKW
oWWHTJ36ZETXnPWiBllTUxpdO65vFP4w66vdUPl1gbjeCeF94lk0AQsMzK9ibansSH+z3G3T++1w
utQoau6XKSyyZXvldfBiSKejfWQafDuRGy2f92UU4GkIJmf7beL6GGkjp0Ru//3Eb/gjDHLb5lZA
W2sFV5/IagtPUVeCswXR7+3U8ZnqaFipInGKTNpYYYANe0IumHFVgdpH1CySXfwCOg6xi3QdDikI
b/3gn0NClTPo8wQMn15xDhHhu0aoTyU4K0ZNrVO/Mqyf427E3taKVosyXFngQRBj4oMP6vo5AxaZ
zP6hJ5N1fdWGR6T+BqFTsmxS0WtEXhJVC/OkZmQsxgRVp7hcCvlLJBdTdZATtzWBNU4tR4Dj6MEB
YSrvW/0iMytEiejN0/47c66h6/QZ9bykjQfVapc4pEkcEToDVMD+ig9+bWHH6qAVARNcQKDbSv8l
Svp1z9WRS0caUpFwgYXDT3yf2vbYdzCCKZjmFhZAU5zOgR4cCVYsNcO0CLw28bgqzELfYa6tvv7H
NZ1Oh8sw2nlWKQ46Qiu4PcDXaD08RL8TOEGWUp8xZUn8P12OrGiARRb9eiev4Yf7g/wK8eL+a8Th
aDCZqypT+jQygUunyIr/U9BLiH8njszmLy2I+TUBuLHm1mKbVltbTDPF/I/t/n2IPJ8cRco8cS04
5sKXoWn6H8WreRlTjlJexjkqzVYnv9qFT99GVnUkYnDyb+a0N89aW4LIvkT0RytM2ee6Nv9OErjo
T2WGixnatQRTtg4wnliCzjQO1ez0hRuCiwbJrb+J8EoiB1humnTl69u2KlksOqbOYz1Tz0OY5ezb
Nf9WD3bn2C1Ea1f11AbYpT2cictAeJAMPfI0mezn1XvcnWfmjazJrM9qmwg0vX79Vov30x1tpC3p
3hrt+HHIJaS+u2vzZxbjLj34Nfe0k6ZCmalttz5v7Ju6Jj83XXEerVC6xeC7zJfbKh5SY4mEpdIz
8q0BbyIpwBFa8kkARd2ANNXKU4yh8Zh3kLL5Ng7yEr5RdXHEk40W2LCLi3WgNzyBJrzw54LH6r7i
YkG7MKOloNsv3ua1IW1BgCOyw1NMi/lKEooV3vC628dFyDebb2z1OQRybOI4uo/5EWNccUVmRdMI
IBpqFyyDKueW9+tCcz92psWfASTYa7eLdSbcq5ggfC6ND63na+gkg5DRuakkH3C/9ocVRpid7aeZ
agYATNCHYVqxepZDuc6S5ZxLOag189Wo2ZZvHostuYLArq6ocrRQCCg3Sq5Uej3RiOq5UiMhOekh
iDcn768yJTGyruuFNOvudn5quTy0U0yZKGOklAVIiUBHDD2y8RmAPfQ8Mi5yOCWbHhHoy8nGzlVT
RCaj8TMgTk3C69q4g9uDj3P0P081zQRHOJvK6VM6Y+r7R7h2yNAAcLcyHwRTwL591DE2VP89l9D6
pP4fh5wmxYN5Ge74POQUoj7/qqsWjtb4FCNB6ZdZh+MV5wSiiRYZPCPIaRpieSoSshRVWTOqHKqW
wh3Ym+XVSmBsSQHH08bV6yoy2l+aAKb7wStElMN5pTv7PTcJfvAG8pko3PtqIi8qSnCSoJUpRo1u
wHSob+SPBIdch6teQJjawgqauGMb2Q4rDtF2pxml02BydrlrZtq+v8ZWCl39CCfFrUTSSwGaMm+q
jbuO/qk41pEih3UyT9jRtG7UOKex2ewSHGhUPjppSfb0JoQjXJGbu30JkG0UnFJkiObhZVcjG6RV
mxH+JyFD4Wr8vheeTbF3t4XKdJR7jYiNCvCmGwT/csUvSMz6qdhAvlVCdEgFZSdDoyhF3fbBIBlm
UVbLaSHeuRno7M2WJ6vDPMMbVmdbNPTySZDOlrFR+fboJSOy0CfEPfC9FOa1E1lXhX7V5maVASNb
unhnQyL7MTcyrbzh6mY2i/MiFfI6PH1hc6T7hDa3GT4Ip8ZJaTkduYI06JrfDk8CpbTAfuFTtChY
4eiLjzTcMjL2AIKKFpvYWJuW+wm37FCi8nGSNglRbxgzX2/D2tK+nFAbyA+U71QPlsMtvifRO124
Wa00v4iOYgyk3En2efLYkxv3JWXDqlIhYPGkRNyqp9XMOeOyssW20naAzKn4Z7mTNFuOsY8GJozY
g2J+u+vWhqezfssZ4PKRtbE+zHDe85jkhhoCvQOCULWNyGXZwYU4J5h66zBrOiBKNaAo6OvcLRHB
YO1PERgnigSfq9XoFhGiUt4IYMPDecf2TeSAWkhzZy2pWct2XSjQqoI0byJv2Fnj89qqhkZ50R5M
Zmvn6dKpWKJj8vC9qioAoj8pwm43gGnDq/f7hOibekIfYPMhWxB+ZhuZerAn8FJFFeJB3yif8KU+
NDtuieCO5V+xQqbArGetaOcROydDwr4C1bG00JRyCtuzX1PZYuEXzzOkoeYnj69iqwAlAbnzm2UZ
cVz4dbw5hFJSMFd3ige+5Sfc96BqIqeOm/5Bv5/X2/lBtPrttoDD7J9oskEI44e8LW4/YINy6mO3
8uJDAJfdmGBBQUi1XyqQuD/+luLH/0YjmG64MWGLLoZMacd3l4oZ62vZwblq5TDiopx+U8aQdOrW
OpOov9NnaZuOfx0r5Z9PdSQjdoIlxF6ux8yRo/Ym9wywXZ83YT/HkookD+sDRIS7xaIs/7da+GVf
U7M9L9/FG9Vf4zfszCHhSqzZTByUnSHFC/EVp+NwtRYc5NqTDLeguJk60B3MSue154fj/S4WMS7c
nhrMd99418zvAKc/XChtSIqTjhd8q6j33RNFYWZka77Z8SjxhjJB9VtsM2YhjmwUrIr8CswMSCnM
mx9FV9xLVmJRoGqkkuuKAm8NjuGKxn/fpife4DMhO1L2qi5n0I9aetNJ4IgVzg2udOpB86K0O3+u
QJZkUWDk0iLLncB7Xte4vkHBeJ5GoFUIw1GMAAkYWA3QfFZ44Lq+kEOWrD1kSevjAH9zCoarL4UV
dDgif9IW24md7kyPaA3Own+xLxQQaPJglOWcdxJHGyqNIsmpKt0JYjczHKPP4a6+dvly70mvJTHD
t9D3KUC+VFAWXKCsra5KlYShfKoatJ6IdWrw7AK+MtdKNw7/kvxxZLOKRa+0sSrhvPiGUrhsVI/x
7xCGp4JhYCVPOjQepKuVCbOhr3IDaP0J3X3D/QVdlVL0yPCYxBnGUGu7Yp+AULKA56CcVLkm0Fdy
1y2lbPNTGyrlII4zOgOJJN7Lh1KQQtKnfbhskhY1KU+KxfS2NixivSDkp7rATc9aEIm6sPVIs8IR
IqXnLMxrIiFXrtOZDmgpabBeVus73GEhsZmFPoDosiDkh1PdfgZ/k5kjS04jreEiFlEw9oYnzyUh
7pKxJwF7qhSXvU595sIyEbBAKx+fBpo6VntNhCvBjfFJlIItylpnr9fq1sJgo8wrDcO+Nv9mVunl
pw3LjMM9HUIjL+RjPJtKM5bg71qn+9bUCh4OjOxeaSduCp1rses/lJwitm+75he3S67mlK+EKCSd
b1GVddejUD6vGAO3R9tB8ka2rV27oxPuvUPG/m5LsYnMnYaoVH86FOpz6CIygL6IyHt7BkWDio80
eAciUNBmrPrbMEJwx2eKgHnnDxgl9LR9/1uThMZJySYaPA4aDAFU5V6BbwPsZtR0OMEly6lXKEWJ
1Z7JpBV3z3wlQs+lPeoYB865LL4Zl8umCBxoTBKY1JEBGxvP84S+GZV98hmdNLNm85xYG3rB+5MV
zvOzzFUuuUzrNzcKaghZkKRLsnKA+YUPFOXMy6ZPjrGoHr7dYIlBYgeyA8opPW8tZrwTQn/82T0x
nIlwbIVnFdUK+e/uaklNNWATgPV4kPlw7KEhO8PDDChyRCLlZk4Atr9kCGoQHAbO0WIsgWnSxSKb
FTNYuhgTR5M5YjhVuIAr7SY7MfRqvXxSIVW8nvd/sGYj44T8OhxuDSFPNOG72Brp4Wmf98tNUW+l
ilVT7Qayp52b+ZrrY4FtCeaSB9Rxdh6ytNTLr4jc0zVD0vAp13L3f3FGJOtxvorylfueHRJS6PCI
CqlQmWfyyGeIUv7/mDs8I8ea/GaeG85M1FY6ZtcbVUiXkfCTr4V+A0yrBJvWNIIB/kHCXia4Fcrw
t4aDFgWD8+pDG7ZZXiRzIHfUdiQksT72x5gmXxNJBxXSOhLdWNtq/NGXwiLvFU1r5ag6QDQ99ccz
HXVuXAeU8voe5n19XyR6fwYhZUSHF/Q54PzmXFH3QUHUcfFg4NHPTYu43ch4VVkzUPLqGxOPgmUC
qdvTq7kIYpxZPFVPoKgQcwKKRzslQwxqDuZFz4SQLrnX1V9iswL3Q5NiCHUP+/fHsypIHEi+ET19
MvSA3sMVd1leKm8a5jg4Lr5IME8f11LPkGXrww0LLUcztxloEirRdaXJXNzA1bmeGesirbh+Nau/
FECagc7/PuPdayeAXlcpBtQzXk0N45WNRwHcCcit7Y36Szpj+XCyGp0v7lCR8BTzUmKo8Qe8YfMD
7OErd2DDreNEYpnsnf0btPYWCUoonSL99imPWxANNmK1IlrQqyjHvmlF9LoK/8mE8JvphfJR2w/q
hqAe83U6hzPiAhFhUKPza5xThd1cbBIuTKgbx8vvP3E80JavQ4GMwDnVei87GvcmIx8KN5bYXgfW
Rs6RmJEcb0Yq96jw4ei5QH06nu3N6WIU8tTM+X3umWcoiR9ZptMn6RC2ydGX08fd7tXI7w0syI+U
sBNAygYC2yGBA7hdo7wMlWRF3mK1QFWUqC0nvGwC76M6E1xYO0qvp6FeHzUTMZpqVQ5qgfDXKBQX
IRTVBHa38GUOE51PlQVSrlj2ge2/3Cp5psrbhoecEFN2Bmp9JMMCX7AA3woFe1Rmnr0qkUaxJif2
GvWJPo2GXpIURFvQfguhtv9Cw8db8ACti4l9tbm92FtxrNYRvWRJX77OQVlTS5f0YH6itawa1xP/
MjJ1akrrCDwPCsDwQ9JJAuzBAs9VP4tOIcvrH7ozZQFXbC/cEUFzXmddEOdDJ5HCQEquzT/Wa3lQ
IuCw1eamVrDCVIJn81c4omnuhqWDX92zRc4d6Ei2IpOK1m4YUMGk4wavlwSjd+uSBxgAfvNIi3MU
bN2Jahos+X6UAIZsW25IrdU+MLakS8IfD/HXUeFCwmSysn6JYW5yEpoFjYqlMX9KAwk0A1Y9zTdB
PyAtYqkrAKFAn28HtEdzP3OoA5cA0wnoFttfdpUly8N0CLrk07l92DYMsdvbuvRIOZT9VG9QIZPo
IjRAj5FG0ix6LpGboxa7qL3UQSc99Or2+PECiC+UtuL6ix42NaigGEfWdNyM86HnwFD9uslCUEah
BjSqFitVLrTcwJ1GU72lBlVHVhfSpSbUuJUnClliGFgxyBaf06FPh3ww/O9kWT7AI7qBlcj2rkU3
JKRMUF7oDr6hBsqjqu8Ma6Sox95CXkAQSRhnwMYB4bGHN6uC6lg5+W2ncIN/wfbHvExs+0Up/9YY
X0e+OlxJXIcoAf1v+GTdP05c+Gx10CxkXFml2DkKa28LINp+/1gc2EetKA4sXeCRGpSoNlg/s3Ki
d0gq8Wda0swrjrB9oCj7zWn3NQ2fKXin9pu5skVNo4ulQbTZ+c06QAsPOeONPfa2NtFI/bKRvHbV
iocSGQ16oFLnbo7eLEZXHVBcsyi9t4XpToP7VBjGsCR4vULnNZZMZpBbKM5fICAL92AQ2oikp8r7
sWEX6huoveit6RRqOqaeQe0rcP8rg+JuHwLBLZMLd9KuRnvS0ZaZ4aX244rprjiAXT7HCuksG0mz
e6yG9qvNZEc/e4kpP5TGGnaalA+FA/Mb1PHbaoLeURiFmjMYhDF35xSQQWxeAIaFe6Rm9Nsd1q7d
RrGPbutbbgHEsGHqEW0iXg92Hd5YXTNWs+/8RUfe2pgHTA2Qclqoy0HiV0F+Vr3L1OLhbCYruX/I
Kj/1M+96hgx2W3bodyV2JOMMz5kugLfM6tKySEHk6hdUBpGMDMqbTzp+V660CE94FXLZCXamQu1v
z0G3RLOPXmf32fZ7SavtIHuXyAXyuibUf4mAuR5GzaZYoR9pzIH3rma6CrkstsrKo/fWToCPUhgS
tn34d7PXdkGMiz3fQXHCOFmK+O5pyU2NUDvUMouHuXVrl4nHmg+J81LpNy+uGh9s2iTtWNjhrnPp
Ss0XcPg2/YkNntkFUBBwp7H3s33bpQ3+h7vGQMM+zbTRONOOLsgPvvpGaJsMtibAZP+FuWKt+AQr
YIRcA61NjXjbNXL1X+n4hdx2GDtBnorm27FlJg+Np+AnxYZ6p7J1pl2f3PWx735IVsBCbLTg6wH3
5NSloRTAryn3dDc5iAeIIz0CSkHig3oEaeMQjzimiDS/2ao22NIgskKGMgbaKEwQQOhXONYJofug
Ss4KNXylvLi5dSbnlqdpjeLSQH0jqQixyB6gm4ortx62KmUlziSVO71FzPLtNWGUDYjly0W+gGCk
slk1xW46UBRBMhrdTlJIVJkjZFK+suoqu2RwO12GKXVX9z95hj7uZ2vGIkRBjQqnEcPRMpr2NCWN
vYHwfCo/+LKbmUivBBMHbl/4s2tEJ3bCUb4rENpK6hAR1eadPXeUoeC5Kf56TbqZry72IumrwSe+
LGytcocO89E7lfzYb5pcJm5LHqT46460Z8kFQ1Ex+5vQJOPjNhXD/ibWj6I4cd+OmVlFnyRhsOk4
NUyY5/OmVFpoulXqw/+AczuQeAFfPtG3z0H8WztR2cxhYidsPZi8HVdGc4eJKBvBrEQvpgsM6Vlx
gUV4w6pzqYl+voi3ZZoP9jeB6wgNjZtNvPEBTiArVcBdA4RXy9sFpaKTx/ZQ62DhjjVehZO53FXS
zeZ2FY7GUUqoE/SQ9hS5aHG+MRLh35O6iGGSERnzlArAdAdD99EDPWIZs9dMicQMWoEITb5l6mQf
oUzzmbWDoCdUtBorvGA6lrrrpFPJw9zzfNvfa+5TEOeduDwfbqAwfeaaJeu7lH8CjxyBJpAy2Eo4
sG1qt8ii58MoO6OBbmu2YKqZTsVHWyfwrrWRs0tD3JOE/ktgyPZlVoqeSXg2dNekaonqHNitb8WR
iZ7nOhjNdNs9CFSYzB6fWBjKHfd4XQib22/dS2mhkhyzELvaGuY0Vd9mf893AgK93v/m0i8clwjk
dJ+nsNgKreikjQUR9BJmaQxmc2DQx2jaDsAz0xOxjljsZedtV/ZDB961EcSCIkJV54+OosX5FGgc
f8S8eZ4M09k1tPsxnhcFxat1KwbJ+H4CHNkRncpcV4dB2hCBd3YlQG8iE8imuZ9ukJgSw1NCYcpS
+2xof+1rHR8oAAXwQO7ct6Qpj/H7BpFILD8/XbZiSH4HyvrC1kFqDgRDXF0qxyqMBIfaDutPEVgd
Z6MNeUMMyusnTuzyPIt8v6PYs8dRHzP9H+ptkUs0Z16Ki02cRfBn5MdWOrN2oR15HpbSsvm5uv0z
94L2DG7CcAlAScoO/ti8gXugT7f5C+mwICi6JWrHBb2AwTiCPrsjaiCCimPmAG7/0q+nSQEmJyjx
EeXGsm/QNPOktMY+/TzxVdId4y7siPRzMiaW5MHwSBxfk9Sgdre+g8+JIBk5vLUmzd/Vcf+s1XZn
Pnc0EhQ8jtID1Ji5C3EE8Zk0AhJhLZXTqYPuj1xD9tz6jaYbpKd2bUxRerDiNDRK3dkc3JJUr/jj
CzCLdV4smaIFQ39y2BMB1yE5u3pSL/AshT/EoK/sf054czngvO3Ed0HiDccPY80QC6JnpJkLbqDN
8od+ZJ+c1NpmySQd+SB7zqfwA/t5uhnHd88TZcFGx9vMa5avGvmaf+UFQoX6l6qFctxm5Cs2Q/rb
i6zeaJvXb0fF8KJSXnhHy7U8TZQydRBKCHNEXHXkdI9KkZJ3V3kHbkZS4FquoVwruoZds9JqNM0+
q1Lt6of/0iiNgz8wVNiIHR8bUzrsOss/V4z+OXCD7kIRAI97OGXiVC0D3SSLZS8mGW655uXQnQAc
Z26006BsaYM68OJVaD4xa/QahASB6np6yDKTr9yCVGUizFog/Ru9TulSGIMoEpo0qFrZDaJ8amo6
RqpeSbKWIy6urMHmNyteufkakLFjXO8trU0MqWMva19KNWupAcxSjwad3A0yk7fI/0ywj+o6D7v9
CZ4z2/Khf18Fr7rg3u03uRr104rgfBCtI2Tueuepx6noYD3Bu6jXbjEgtf/qXCKIaCB8qxqZRy5I
LvxXAz2UzBrOWm069EtYR1PfMB/jWH+yzI1w0b4iVUBrMtg9+8WDT0rabEKryyTSxu6D1834KNTP
Axq8z1rWB+RSWk8B/kVP/k1Vy5/T2OxUlcnS8qEISm7gU+lQuVeK3AjAxm3zUdjfIem3LAEqicGy
bIQgQcm0M4xy56vVD4Fx+tueU+4oQj3uGGJhsgnYDKf/oMAi/Z3/fIj+4QK/rxrxEbSWO3wvCkWO
fH0FpdUdLTeaZ4ONTCEEpO9qEyDCRnemhlEtFI5dr0Eyjn4pOHVS8Tye0AqDuUhqHml8HYSlBnVT
w+34/dPtG6g56Geaiz99QbDXl5gnaeo3pA6M/5n1Wsl+rY/rDoKShZXfV9w4+k/msVm2Kp6kznj+
gtGxpXwkPeU+kzdWrjnOKuDFrGttNDWdUtAE5KYu1Y6aGpFb6OBMJ8tRBpyeLAkkHNi5eim88ZqO
nbsZShugithBY+xta2BKD/2NA+1Qbax63LAgXRdVBBFcnv0hfRgTYyxcDmiIaAODgAucZhNCL7eI
8uy+PA1gM/AXLX5HnTFBAwgIOCjKTyRV29Nn+DMllOfW+Apg/vTJbrrg8U01mckPkyESTXU8l7oK
BFZC8fRU/VhN/Z1jLvo5MBqe8DmpmUpyFrSx5I5jGvMnI29UGR65mAmbYMVuqz/ZPEllIovbnmXK
uBS7SZ3dbpN+YuYsEfs4YgXNdmfT/Aktnu8/MwtS/HQwgB6s5jO+2YfdRB8wQBy8IzBfCt8PjyLZ
eiddOhf8IpUdH+i1ixY74Uy30eeTgL3SedCr0wP4x+l40dc3s34Z1U5kMhdecOHqHy/ayraSVlm+
1AHMVwa1yGV/BqVMAuNV+4GKVNP8QTdpL/zofnWj0Z5i8h7Pqm45CUUVF8zF5Mg0jWIk+0KP87Df
FdKvlOLtXFjsjvJxNqWgXZgA+If9/7OQMoEyg6Emb/p7EoNZzivjrNF2tDFe1ho/W9PJWKWH6aDT
hHm8+Ndj803CiFfr8gF8oUin4VCf7w+JDKZsKqLw3bp3ORgHyQtS/JwYIOuUFPrEIDNDCwIpZeWd
Q4yr5UJ2esArmDFPiBPZM7Fn3z2DSTQEuFv/GICJg73+eN7W2AAlyycvNpmeVvlogtXVIXLagUvw
ISg+UzB6QqQcQlGKmYSd4RqQ3AUtmUePZrvzWvuR3t2qHY2+1biil00Al5hmf4swzQwzJKkJ6HeK
Ir+6ROC9YW8cZYX+sBsnZGJy893HXSTt4Uj1KgGtAHCjl6OIPL1Uo8wpIs6wnS9wJm3RkzC1+E1X
MKTVHVjRRet0Ggv+1b76TAEIYPcNNY14XcVQSH3w58E5xhYr/sUTARnvjYcgun95MgWzN4CZpL9X
U+K4gvX5VBTrbU63XdwN8ZbxMawLUy2T6Yl0rdNI8u7wOoLg7SOfs+ZNJpAZkuCgFKYpDoSs7YMc
8fPd4MrNtRLBcV9QNgT5alvEKWmNpo+Q5XqAGBN+evoFD6ABWizWW5Ci+0Gdv9I+fdcLfAYuispC
vyZdR/PVqIleTEcRt1OUBR7oJ83cObxF0AS5IxRnuoBR2MYTpeE8nYLuvkxuk/2ny3gGEbKCcMIv
523wO4jPVZruoVN6j0WuAeb/tZnwhhnyn5hK2AkahTB7GwQg2cPS9TwcOVHQM+sPt+JWoLWfmTUC
8ttFiGJkhGYn0l7LeoIRBQKOVbDStghqPA27zYIRpwEUONDY8szamBHhbzJpQCQSUr2uOnMNR8tK
tD9qesCbH54fcUrfi+ETPGWYXJ/8n4eFODf0P16aYFYBC2qy6LdpllbOAh15HTbEygbx3Lb905qe
2QgMbRrN3RW+sbFIM7F34uyqClMOXLzUUt36ZHDVogyupFpKD3OloKVxyXhVp3LPnhXfWmDWV3yc
+URT8AKSIiX3j+Ld+9aLHMRqLzfw287LPFcxJEOTUArKTo4vmev8Fcr24rKqYgD6UHCbVMKvMK5D
z1aar56vlCnufTbvm9nLoEJx5/njXycj8+n3qFq67v9A+TfbPp+LIBQaVvcEazet7CNWkr1gFYwV
FM9ZCE/uQW9XZSUUyRTqNQEalWl2sOG6HQhol+bIS8yyt8r1afSJSiAhC28dZ3HvXQ48O1BoNUl7
rtxxPYcTwZyMqyNtHfa7YVFvl2d7IZbMDwah11t4VX25ISF+kO/n8oz7cYNNeVbKSZBv+f/KUVee
Byp8bsypDbhhnlqvDKzLII19fhLerAJD5oPbj1fclnx+7uMlwuOeJJipjwSHmbOZodAYJg5HQEg1
HhA19JVP4DKMW19Rs/Mcqi8aUslhvvFZMMFdriToCovq8lXXQ0DVrbA4clNJEFCAI8PXZbBeEdMv
+OMozxInnnRVMmQO8sTQgjfvN8Us4aFyisnuc7moyu6lWyEKJRVbtEVHK2H182vIqS8acwcqBfQk
0koD5mUbXKPADWCDDgCGtDeP94BrnMjpQN217lF0nfcm37kLxHPKUDrKByolwc/POX3qjzWJX5d7
pjK5MxoYc9lRGgj1xA/yNaLVn1/p7P+66cPt3VtSWitV94SaH334cW8BHdNk+R1gqx9p9IlQfvid
gLSemhqio1KOYtR3mEkVq7IrzYpDawhOyF66GbYhbqmi5U4ANiJfat1FE0VEgE5dEOR6AtWgBgJJ
VRKIf6sPm/wJCc3Hf99R20ECyjOW4mrFbOVVXqCugBOV5Wg67YR/Cfz4zHAlQc+arqsw5o1bcHJZ
F1M/+p2q5rrOq8OgiuIRrnK/zobQddpONYVFB5bHJJWM0/kLNuiwHrGVHWd/M/quYECT+Lt81Eji
4YcJDX3GbA2WubrEhO8/JZQj9ipy3uE/lxd/eUYySm6nAMSvC1a2+4bUI/ZXKrHNl8BqtSFX1uL7
x4fa0CXxWB4QPwTAQs/tGNj4l0tO12Sp8TCf6hns5RFSx+LbKz74BoXi9da5amhxU61Zta8gAvYw
NFzkvGFhN6aUSJj7WfEROIR6Kpl2vNnqk2J+RqbU7YZyknmrVdRah6NM9tTyc2jUaMniA5iSC5sn
Ud2O4Cqe+HhkJhobe27cp3FqHBnwsuyA0E+pWBAeDTuUOy335sMHx1Ow3Tj0/1Rx+pXF6te0jdsn
hmWtj2Z3Dv/mEwZtUFuVneM0JGCBD0WpAEbYADzyJYHeRYzekja+t0quMwkLw4DHgnEkWz2yGId+
LAwAmmy9QAesCkCO4x240ykHB9EOu7yk9sPfs7heKP91ousLtWVhQRSHckJTlIJgP18ggz0/dsH1
9JqUUyz3n5Q704jA/QS11b6H1cmEDTL7Ry7ZcJ8IFg31+oxBZFuhskTCmm5yBihovJ9ekK+oOWAm
Bil9iiLWoYieINzdopEJ8CUn83C/PaTn2csbUgsR1tIWpDxyGhpeGvO+4gwq0mnzyoDRHxg4lq8U
xdwLQNIuvjxtRwxim0x0239CXTz+Vt107kNWwhSeB+xd/kHYkYB/G6NWqibpYxRVqBOz75ae/olF
EWy+qbE5jPVuaMdp2TLHKKYDQ+ruKgep9zZ5+NLZJ1Fgwh0CZqYjydVx57BpP0GdxZb0ww9ZntbL
qohL/L3WUANlDSEc4XLkaSQL7HVoEfQ2Om/CRFQv9nRFEaw9ZYeL4G/Mhoq9LH1Y8PJxUkoN/Bdn
G/QDLz+uDyKhKjmNLPhjE5H8y++4Eat9zKjpJtdbRsAW4O6qyIZgaKJMGWlHAOh9vsWiIMtglEBN
lmBQ/rV8e9MFw1S2kLiGDi5ZrQXZfcG4kKaHIHJO32R7x8ySlzPkMm+nM44MTTwU8zT4EtpHlfym
cf60m9CCNXnNE1R8jjtVvv91d0sysiWbp44VZEVmCSMAMXaP4d0i7xT1mzH2Fa8o50+bq/PsjcOb
ajhcZ1MRm/ao+o8cpX06PxkNLV2oC5Vop8SNgBhXoXO5LIsWf3jUclDwoTNIGDKBje3e1nfnwPCr
zMBWzTsX/wCt25e3CZEen7IpH+x/6ogHfRdYMHbuD98rC4sxqPp1ic2wATm/syrGoUos1NEf7FSb
lOyUyj7znbmABqKruRyRcS5VKauaX2loGBdJFJYTK/AswT6dg6ntrDXh3QYDjWPFTE6xhQYKiG7r
7XsLjtRi1aVvwa25mHcXBn3vZ9KQFqLa9QvfogUWkMhstzU76qz6gj5W3IAIEzXnudP+YC+es0AE
RTnGZSRTv08ShDG2NJicakntPUYBMAhddsRfmKQHsUodpGTpMD8cquL+XjGXouEIIPqDVzfY6RQH
O1IXpX6pVzaoGZ2PSOyHEIzCSQUstubE7F3lXs5u1Vq8U3j8FTcc0LGfD9uYIF8PjPMqvRurBAQe
kooy2weu2ECQ5V7gK/3A/bUmKj1KO+DsR9RnPQpxPBXgPnyzrMDIwjWfT2GHCn+vI0vwsB/EmgF8
KrqHlpdGKRHitDNIa5ctZXuwzcxCJzru2+CVDzgln3WGT1dbEYOfacu0+l+OgciWrFR7uKU/Ka2c
2S27A/J2DPGtMJWc4CDJhfsOsVon+zybMc9upIaWwW5SMFF/ziDibci04QlAX/Dkxgbr42fps8qS
aezYcqPwNx517/PBlZ11Lb+vMYjh1euPTRYwPvn1QuVjAaaX8BYlF4MJgv25HpomSAyQx3L0YYv5
F2UisxJdBIG4DkT6dF3yYJad/XVt14Q5pPs37hmRDoCqIdVmrZJEJHCmxzve850K+5f9Ad6jJx0F
KcA2L2K/vwoQxGogYlyOneUjrll667ZPUfyCY7qWdi5Z/2ZOhxyH9c48C4+jU/ikH/VEWg7vog0b
tnRcQYsPlpJ3SxOyd60QK3XTP1u/FMFP0qR2x7dKV/D4va//atyi0i2BJwM1tMeVUqrV9qQbgsB3
2wYGnKy/FvXLnrcN0FAPZoY8qNxinEwqV12pmLxvOsK5vgpvLdchT5NUoEyNPv913fR+xRDV1mB9
Ae0yPJTQ9kMY6ZoH6Dv/07msFqVIw1yfUDPGxwWWU6+OPzse5/eURyypiaNZ0b24wtHQkoEIhPoL
rFIk8GrrHz2NeHLjIHFza+9c2yuiwIURFEM61ax8FGDpW7YTGs5rhXfM3nUXrrzcvNTgOV8/2PLw
wTGVKTvQxqTkr4RZSOl4bL3m6le/WWIgFMP7eZh0tEZ5qLl33X0hHrfHHXRac8XzyonayCEGMpae
c+W8yEe1IodAkw9nMVdvu9fRdEvJsXFIFByn4Ub7DldZ1b2FwjCIqFBtQmJaKcmakYCtMeM3xFC5
mlPzFoxDl3HWV2yRWqdiEZ0zmJWqb95rQmHlBWLuhQe1Vz0GKkQlzJwS4suCtuhAzTwbyf3c52Id
9nqMx8ZKZpsjlc0isMRdhd8Cn+Gy2v1Ey/2cF/otTlhnJpCbszTMGlmRP+YiZd5/WwnAoi+vI39b
6pWLSp2p28JHpECsete76AjL4jiXGp+Ga3Ad4yk5x9NPL/Hf9Htv0pWPrssW3vsJWkEz8+0sYo3Z
TK3OC42PH2ncSEi59JJG7knz7CZI5lMgToOaqBPMP6/gV4djtsEdpF1SfHlntqoq9+fsHNF+j3oT
SEfMIf1+owx/skJmHIC9CQMHjvsFSX+WG4OAQaKJHuZXBKRI8jyoNGJWPw5mOijQXGrEjAr7JUmb
kLsmdgavWMN63n+VLEsp6ByXMwrZjoTIpviH56NnaP+4kpTY6W7LGseDWryrTg/xh23QmL/dcFzs
xUFGpY9loJUUD8mw9CUyqQ6nPRfKf4BHUHZGpQ8ox1Q+QnE2Krsm5DShd1cDkCzoJmGxWpx3a1R/
pnaXSwuh0CRBfSRDch84FHkf6fNAls5CirreLb+sztLl2ELPno/XrjQbPMYkQd2ZsnT799hD9rLv
S1qxzii6h/Zv9D0i+icRfGPy3PuZdqh54JT7L0DgAv598AjFQ2VxZJt1RIIeh2Zh7v6JFy3kIwBC
phZm9SvfWcwqB+W0xji4lHexbNSh487QSjyQus2jhtI/43kqTaz8YkUh/LgcwXNbiTJRZ7mtFmQq
m6a1u7BNV9Ii/mt0fZm2sxsDAv8pJZl48HEBez5OCEGJ68Uc6XZyCem8QW9v3h64vOmHFSQQ2LW3
/e2Zh7ZTdulk4Ph4If6eS6obxgBSTf82KdKD+MnttFq4ypGWo6fpsM3hDjqItbIQqIJbRLoUoB6S
0/BJRvbyfIKkfAGSCYdqmDaSu74TtivIhzpBtzPl1NqWbfjuEy76b+Sz7zM8A357Buds/j8T9Bjj
YKVtQFUgJVHnF1L4d0ZByRSBq+kCdNgUvTHMfZD0kolgX6kKflk9QbuZi+tswZXOcDwS1aP83uQ1
U6VtnFE7/WEsz8jFjLs/110tQlFSwz8+Rx0YjEO3uhwiu1TAQAIwc237E1qyDOlrlLeTQnvkh3zy
0ULjIq3TJtGZ/Bb+JrT5jeid8BaiwOnu1JQ4UxenFjc8a1DKDuGNLzYr+DOh/TGkqW+lUq29BGbn
jbAGu0WXPSCVSjkbUk00QytByM35NDEwZvxKk/B11I0YoFHKEw/4fTaIqiGmWS+T9+UakSAU7tqj
FItLW96gAyNU3CoLuHGcV0lnt972RPmiVg1mXmN1Q7FExLtmQughwLgjT0SzAN0u2qtJV51dUOnL
nhUFexud/EQVXHLNuZ9jhnNsO2QLfBnEJiWBpa2jGQaI4jqBcIAfz7JRxOIOtar5PeoViICX/ack
NvN3tjgbeTzByMxJmHI98UAbQlJ2NKdVIStykY83GaTeTjbAcOXp3H7t+E4FO2QNOxPS/pMy8Gyw
Gy6DJlFwivnfVbza9XaZZH7MM8s+XzRAI5tRlVDpDjE8Xyetwi+MfLDJYCmwspCBXXLhDT8DsZxe
aNRU4KZBNvH1C3WtP6g5YOPx3AlRc3t6+3jN9kAh5mdV1tsLz+vGkhE9f4FIejOUauPiUYSjZ7qv
GTko+HSEH8WcgfZQJXzJOF0BM6td5xVp6rTLJ8iIn/SKJuBrfalE8aPGPmYNEoeSHhHDFLCyqAo5
kZ/x1LizYMibrvZobupuv9/HvRbPUWJjwCmUJCOW5aJJLdelpYTxfOYPHraaPILa0rlrDeE6YkB0
qi7AEWU3Bb5EUiJjwcjQh5dG1bl6MpXTLkHtklvkJLY+06wJ7oy8P7HvQFxzTtVEEEyCh+QPuyWh
ITMJKEcManJqJpUd5Ge1EHMa+Mkq1dbHIS75WIkA8n/OF9nwkCz3OUs4r4mtJTIpZ8wGHUEvlAYF
MX/iUoyFgjPw2b+CgaJTDyX+bOP2R/md1BqSjSPkphr8FsEEP7vcS4/7JKQI8BOamDsickI/Qdjv
cleYHV41QCqAcC/w1GvghIaDMYjsuQgY3B1x1HbRc5D8pSbfbhuYv2WkH9sfmZUgJsnJg5sH/BcW
jJaxDPpzgTb4J6b0EtaS72cza/Bok5IK/rnGvtp/T8ZAJh9wBYsG8DdDW6ZMWqzzKY4F8hdSeeUT
W9CBizJmxb98o3lNYFI/aiUis09xbCiuPYZAXBAIfv4uDNtj8/NIg6+M3eyRMTiRU3eAVAyj+TYq
MZfNG+jYdFan7Cu7Qkg4f8P4MYjKATEoowWmfpRAgojM4KnCTAtednolZUIoWFNMqCWVm3y90jlC
Nbt0SrzJGaC6RLv6/5DvZTvQkikiqQYtRpa3wvp+0voFDsxhBL/2suSZm0s8W2//modwGEMmm4Mm
iP3v6ufJ8hiFKMbHGu4drGctgk73ODWwYxrlccKvnKWeyqCOdLk2wIHNXF4SSAqQY7qPTbLSrpqy
eMS9T8Gfv+dBMeXP8bbrw/Ff8zIvBp2A7F+9T3lH8tF+Rbn1WcY5o1VKClvKcTZpdtFFPAatoA3i
VZvFp0jX0W4tTlWcv93THsGtqI9KjLVd/oaMW8qMwBBwG1EOXX9T2Aq6+QvkzJD6LJ2OQj7upXBe
0PYsVQ1NahAaUA678XfikcrDrXaJpZrNA3XTA8sDw8HmWDi0aUqfGq6NrPBTpQE5sZ2WO2pJxO44
FGaye8YvR1pglH0UCeYY5CZXszp6hbG2JDewtRG4pgH6n3H+iebsO+7sv9hlGSwcq8O7Gr4rf2ky
6HuXCXmEuzM6Stg1MkR6Pa1UE4vfXMDdbVCL0fZm+DrRqOB03qRF1U+29Ev6J49ztTpVCNX1kDxs
5AYTblTrhtPLD+Bp2o297YF+7L6vSiXIcrk/VWwE9aSD+prkrwpySDlB+5LbYIXHwx7bkCFU5m58
jIRBZ8rR3nQ4b5oTz1RmH4SRwHLPwvlXgRDdZX3wNVN7D5dmnojzi7YYxaTttd05ibfPFMAPIKtW
bJOR1EFwWfV7HzIEjLkRbrn8Sry49Ei09qKsgpBEfVtQfFtTy2chxMP6qCgJKDCw7g1NtvGd8SHC
VraATLXAPpB6CZrEPhTEb4f1hkzUtG45MGslvdWEEAOYSN4Q9LZWAEgDHprQcIsH+uMFCkKb1olN
vajbfwyDFqLt30MCF1y/q4j8BroDmZG1K6/XW7SD+l3AHshww7bSpca1nNo7Q+/PKnn14l6ZR79O
GhqJxBCVQ7FjtDJQgJplY4ZpoLEUM4UAUEv2e5kTAXaa26XHI0zdDD9FHWEJOSqoELdOtwE14msf
UDvyVRaEqaLDZuAMmEY0hVK5yXWEN05+pGYT3oRPTcIVclB6TK7vTYmd7MBCZgKhnpkXsGoaDne8
VpVcUMJZkCaEiz69uJ3hdIVTL+VpuKCSqzQiHYFbCpNj0HuyYEHWycx/+YBqEhMHkK/WozZMuXF1
5BBKiygRZmiMqfz5295tN0NtdoN9ZZG9HrQFff+b7cg785kc3LGGqWyeCi/Ck2wmS54lX+520KqA
PMZKva5KAnHzixqyXhPDJK8+bmglFD+ws/CCsyoCsv3lMe0r/QCeQDJMozbA7H42Q4YrYIxhP4tE
Uc86af0CtYumnfQXiWBFb4/zUJsIN7SlUiGlDlpSjviFZMfrwjtIxRG0gOjnjkWZ+N70IZ4hvU4N
xYjCQxFw9gmJ5NgGyS+o83VNp+vFJbOj3Hl7ihjisIKG4nz5ZGOMkIr39FptIA1fbtvfPBm9YEEe
azX+JcMCICTJzAOJS8jnfuCnrBJlTMeWbkAGasuKJjyviRMPtBJfzLlQYOiiieoA7femA4YIFFnr
3INFp+CYLBqdL5jQ+Ry4NjTb4yfEyLqDVnWTzu/7h2gVn8hPmdV51wcBrP0/mI26pG8vUCj/miXa
fqxAoWMLnvXI1OXMCToNOdFXBzJDgmZJK4c97TCD9I6pgSm5diqAze4pUuFQseeyXixNfzngwN79
QS1xfsoNoqPRY7go3oJOaud50Of2fDikLEsIQ3hWCBxuapzeqhRLa3mKqH2d5tvLw3xOlutFSnIc
xlDWItjWWfR6XPerL9lbDNXSZdjcSTJ7HBO7aHw+PvhX2gdmD6rqQbH+4drDKw/aW1rk5GpA7Kew
GDmCjzESSelvyK7nefVZdTPL7UZ1GiKD23LbMYHRohO3xjtagmDCtMBp5nmyO1Wq9oAg3LLVxyIz
w2kjIWvzc27cFJVq25W5oZTkH0TBvRRxvkzhaKI4s35Y24olYTBTmUWjLvznhKmeZXhf/jHch4De
LAHs22TA0l9xPvPCvchMYwvasgNS0m7QtOf1wKMelK4rZT0mGnMWF0Ci/63wzMzU3R77nLUKeQe+
yq67FLCQ+TbUpolU1y8vp7AiZjMp2/YRZUsX2WxAUJAaugW+Y6WgqmZCUGLu6jlm0GGAz+jVTgWp
mk4hGSX+K0tqz7SeTL2zeA0xlzLxf+6+tY/kdgNmE2b1+eqO0Gk+NU/UZpRJ8RGJlBc0mwLRVbP0
kzprOLwyJHzbnr752nipaKTx18pdObtarTxWAmnSw/4qhKItYXr98bwzGqOk/z+o+DxjHhYp3oY0
+IJZdrd6TxOWAswsIMRNnHdBWSR27hRpRpjICT0aEHCR8kwDeB5e+mfFD+kDWOGUh/CCQ1MaW8FH
gsu6Nck61WqEHCglvLCky3HT+55M79YBVXAKaXHrPdOSqja5K42FvPEu6940LZ9FfWW6fwMjHVHa
LOPdD1TqdDu/nrHjmPE2J5wiL+LjSJpSCB0/sg/tr++cT2+rrEfDIFB+DMmqy5QMZ9JtJH6idrSf
UbOxJeEHul8R1yaDoXL9pK2YNXptFVKR3HX2vAzL8e5p6WdpGCRuTrJdNE9xgH5d5oFsNI3TOhfO
s4j+cwD5pdilev6GIBi0pugT/I7pRYV84KuYX2YfRwhHB8rakC20wimf0PReV3kG4UExEk7Il+No
p5SZT4wOQLIFQ+GwBvY/ZK+hvIZD3vPaShNBGjwAqxnZbx/hPLrYDhBMA8Xr9DC4NF/myjcHoJ0n
rb0/eyQzUB5fidBXcbvgWM+X12uuWBk4a3BpzFQd4qcvpXcAQpG2Z0P222+jxrZyFjy9V+P6HrHN
2wwaalMljujoBVhBtt1BXY/8wicpJD0dixFy7+ueJM3BRAKSMlwpBm7jm4F3JKX7oh9jpgn4Lph/
0j5ti0yLI1lUL7dmBQXQiITQ/6E8qPJ7R+7TRuW7eqkhKS7WR1ZeW7y8Xi9ntiYpmshMe6eZBIpn
tuZDzJlTCDdJMVCPW+9QEUm8ayGVQJtDuASGwLgIQEomnlZR5rEnqfAkh2TkpK+qeX4f9io+SuWm
Nl89syhM+fzYTDB6K0mBEdfQKpRsEG/FgOVth0lxTUIWBGU9wySjp7drWsvMEyB+IQgNfLrmsfaC
uQOLEucb1aKvr0nw8yUZgfvAAskuVPYbcxEAdeQ+RORgi50I2jXDGBmUeMQsF9tQSlMAC3ED7BPR
3Fy4N8SBEDAL2Lisp6TTHbvbsweRVESMMbVPXpEn4k3fxNwjOTzT5lOaJvfuVEiJTiOXk1OCsYPf
UQKS9kGjwidh2FyzVpvpFvk9u8JAv/QevcJU2hHeRjIewzkvnE6ZcNxejj0E2YPgBKcqpN0aNW4j
/20CWT8E60B8hLS5kC+tyCojeQ5/TLs9+kQ6/cB9fDTKRzukzB5D3Z4AN4vRdSDSs4ZkNXVSZxvh
c1OdEMlN3a2Ht3syZUFRLYkL74x82WYxPV4eb3+7ObG9hfyB4PJ4Bofw2s2zlVstRMih+XcOo9Jw
5aFvcYYtWurk86C9zENBttMP+Z3A70WR0LY/oBFStCf12NButi2vMV5so4m6kbZ5Mbh+JkKBErDH
nzN2Se2p3DoiImZMtD4FInJHHFUYPc+vLlkZBW4yiMi+K5H1gI5R01DYaiPX60bqwI3Fj1KpoSUo
lw5lB2SOkCvvUPenBMrJUOITi2LmTzKQa1iBzjgGASZ4YL02EkT0yyGvv1k0vyW6lrqFjynonSG+
BMYaBYsvSQoR0GIMVXNHEmFytSRYIaYWqAegCFq5kQeoVR7Os/XkGCqc4orGyV3QYGbA3IKG6199
649uP58kKnv4XxLG9/UWltQi9KGwj01pwyVBJXhg/MfY0L+l+mIRM6Y4Uj5mJ0mHC+xtcTQW/6qC
LIIJbNSGOFvHyyYPgq7gkHckVkBtw9VYQ+bawuMD7S5RJP66+MCJzo2FTYE0cbNSgvjpg4LZeWby
pmh5d6jQpQcyHT3FaIs2js9iJKBWRN2L81qTeRkwmdk1ycQ/scSU0CUkhcwl3UgaEgZfwj1nuRjL
8I7KBsDGq3L8h9SJU9c3kW5JSQSJ0MeLzFaJ+Sugv5ZdByHKoAS0tgA5bMT1SYFTGFnjQlT1X1sB
tXkvAYwaCTDmMNcU+bn/c+MTZLex+lVbSQl7JCJ0q18giCCzEAiJPn6GWcZyxhP8Qs3cIbcz0EG4
SSzv3OGQIUDmzoDuM5LrfdGpFIzqvCaM9GPmmvWHCA7MH6H39II4l5OpPbJdLoX3W4QWF/UEyyAU
Dcp0R0ddYOtVheQmZcuD67D0IYyBcY6IJu4sCczr0C7gGx2VTcW7FQRjWb+fxb6pnL4fLs87rMki
7h5IFk2gpL26lNeVTSsCH8+sAH68/ia2wB2zrCrHDjbx3vz8dR7S7rcNGhYHR/tdSq+kAgBbfdCQ
GibTewHt082xFsGWM3lLYvtwh/P948wcMo2O3JCconnnKP2FwrUpuqdhZnxERB18bsxbPMghRP0P
J8JPJcwJRpQzeEW0RUBERgIQdt9HTO5C9U7Xlb4VqS0IRJS+gN0zhtg7JyhaPtYakzrKoXHgXZdw
9VSxQFYChu9bE5kTyoghTpgKgspO/b/i1uVOiVHJWHaIFmDNCKlDQRK/rBRfaqVg2wUPbmGXFDFe
NbIbTuMYs1TcayBroq8vz9g4Jp/5cRrbRyopyKiaASKrW1nGszPZ/4SxVmYCENTti2cyt/SICFLP
zbzZEAtPheroLU+fEMcWU/k731Ib7DWznHe7B6EIC6s7TWkc63XB+IcloL6ZXTH38vSxblhkgjL/
Z32T/q+toXoibCMKgml1c27XUuU6hUO8yCaSzbv8QQ5iY6q4uHXJW89FoII6nafcA8tHBBCJMBuI
KnrjnaF/RbDWGdOftslYpAKz/9fuoJY6BaVqtEtDenESWQKINTo6Mi6gMqo0mlg4u5QbE1uFUKCn
EV08bCg8guAwDm7rF6m5g8SDPdVjPzUsmmtzP32J7nLV7qpHc6uM1CfbezTm1yHmmfg8xqAGb1Ak
++8uhVYlcmMF+TJf5C+tR+TNZJqIMOhflZK1OexO1uc6KEz/5gYzZZSntjEO9WCxD50heJn2POlp
Qa36aE9YjNsNsW1+sS5nJuonCToSGv3Hp8fxynwjPjZffsnsFwmZP63oZ1/b+spdnS1uT6KYKr3X
lBUZDhrb51s6Y6qwifat1G4oqe3gDqF+38KEZPApVwntD2GaYKUYsZtSg4TSihyjy2C6iISJPCw6
9xUXBslcCFnd+EVTGSQE9EAs63WXELDmmu5S60ON1x7ya5xY6SdGZTS50JEqvVmqVTVs0Iyb5/Hx
rHzKck5/oJEgvQ6SLOBdRromXgUx/M9Rf9WkDrxaAH4d1dzqJ0oIe2XVKXMfHMC5qMBhazd7fIwy
KhNi6KGyFS3VDuKb0EG0i8VKBcj776P6cVO4EvbqUTEG2LtSsEqDeu2WQ/JmSBgUVEt+fAz4plc9
07LVNWjw/15gnSmwe12d8bM1GKjgWKMuozJEbEs1caiuaL1svNfErimHIjZOjLn96iF8E9ALYrkn
lBAakXK4jIR0UZ1wq4+JZ7YErc91zWNnCoYlEe0VKU0cUTK6wvdZJCV5OVLvkitQS0FEriK7KE0R
u7guqWmPIrLvzuZJFHEo4hjzPKFT56qwvvqWKDNJlEeV9nFOXquj2A7Na3SIIxXATfPO0jD2QRmc
VsgLXM1XD7fsoMmXAO5C/+2QfLXRoqaEIguWDikTjmE0txqHFldQa8N/ewt26nucPzj7fFZccFhg
uwjct4qbVkLxfkWJriZ6mIFeMfMFJHQYbrNTYGlySg+FmKfzgTTQjp6W+OGx2WHdVYE9WdoseFTv
xGJ21NNS/DJn2VAzaL9L2YJfFsmMhZ3sM9yrFfyHcC5rdgATJjmcCFSM62k6WuuA6/HLLMq++1nS
V1M7Uzl7LhZMscQgY7aIAJPhRE/L2RyjXk6BO5aKZ9w2INjaqpUhLheXkwbYLvGgdXj9eKSjA86i
qy65++Z+tna8/vBN/nFR7ZQTjQ7WMfCJQCnUAjlm234b1TBco1vPCc0DXB186ak93NOUyFOvv4XB
nb1N4PU73/iQjTgaD/aq1AoTX0eY0WPNzD/fOE2NkG4ujXnfZ7fgPYFYjgSaTdEeiO+kPftTSz8M
4X0ZDXXB5baBEoWKJ9tcmP82mZNWVF4Ia+H7PqK90Pfg7q7xijrqF7HDGcEVzuJaysZWAnxRMgE8
vsiUcZnYoy8Zda+om57qAKrqZx8wjWMoXQCkFobK+GycmYGmk6dZSSV3MtgA+owGhc/RFgMvGeo1
FO3rbddkmMmJxnLtXyA5QuW9im8I6c0Mm4zGFpmpxq6Sfa2APddrN3gXuKEQSXzjwrgGGgm6
`protect end_protected

