

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
mwxNacl66MFUVIMc1Encct2aHZOcb2pREujQa4vWHOpoY4Ryx1q0qOlrkehqJnJB6VdIGpRZ75ar
fafQO/Fcyg==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
WTY81lfpic8wiNg2xUTFY/9pIQI3CKsiY3j1Z19a6adif1iCy2STS25TLTe/dZhZiWj1W1FKdbVN
mTJAkstRD1IiixRw4XPUhHS0kg8DebELiBmCxBLwbMicqplV5b6X9QbZ+d65v5AnURtcySKvK9fO
g9n8up28DiiTZN5JTCs=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
wSJmxWNG9Vaz0hV3ma6xxbW6Q/tt4VebLF5ALUnEWrb0oMwD9MOvKTVg9bgiL2D83XqOs88TpeXX
Ifg7m/wa0qnVENMQDpzrbdsY0X541kchr6nHO22IjxAZU0y34IzPOD4wlt/LkBIeRhuE2oOUmiUB
mj42HGuDYM+OLJ75MJFObfMegkawW+dQ5MXJZAvaZb3Gdq+Nc//x1D0rUYdDzCYkIE6Z7scW8Wik
/MJTbyzmOPOK9ZoDJMjaYzyR5QyLAdSzLEdKbGH7TxDHRl54Q3XCa50pfJuN0PstSuaixGzvKQtH
Tl8qJKpy3o7KeFGSzvILj3NDt+zm7na/fYnOyg==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
TWs0qYIcIilONYk/cz99Kwd1RIRPFnNZwYyu+ici+iMJ2JCkq8jieFKJjspKJpdZ8Nc8B4CnG4qj
aN9KKPyGY83yGWxxRkXLLk1fDABMFcSV/QWTMe6VkTZV7rSzb+eWC79VK61VEPbjbvhhwl9UlHat
EKGcZET/5AsZpsdS5rY=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
J9Mi5TzDBer7RNgnQmNNaMr/oObsCpVjypskaWXDXbsUL9Tz8WTWA1k8rjWfCv9Dmq2LFoNWohyz
5PixLjvzdMk+0EAtGJRSdyjvZnuW2bmu6ekaURxk6HvWMfHmukxtVO9c/su/PcWlhTBaWmQfDEOk
MXt2eXdYnsY9DHX2xUQnYdQty3UwLIiL21L3I3SO1yyv2PefA4p4KfovFGDUvBPco1deVqNYRLx4
GphEA4vKS+OANoIaExoVeJSpvDGH50O+wbHahIOE11SE2zucQ8cWichU4yUJXYALRvrOZArC8ClG
ouWj0ts+fBWmUc+Q65XK9XqQ174/nPdN3w6Fsg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 38784)
`protect data_block
P1tJ15FufyyyvU+FvKE+xwrnnbfrGMhx2B41sKFSSlIdXz4Y+3TS/+l0EWX2jsaxRlY4f3i9bYm/
MMZTnTmY99Oe2oA4Xsw8kDAxSpXp9qMinl6aXVB5gNBUastN/PhYpzF8FI/RfC1NehH/M3OuzI54
TKtJg+Fhlj7PJiPdQ+iT4OD+UqUmZiloUTeq76M7ISaaJq9oEInGX0aR/Hi1L8Kmv00lHZlk5ud9
EdZOQKu/o+znqnbMnV4tr+IAJceZHYJ1owJXzXZvRcabeFstmChP91Z1hiSBY9VVC2cKKpGGO080
r4u29j1j0oC2Cpc9bvk3hqM5y2/mAiwoBaJX9h/pao+ZBzzIVfSzw+vc4nxplX+ZAdOifuapEHxk
r2U1+ymgAzfEHbQBatbELD8gRlltTE6gRxOw9OjuyCwtdR9GK4FewwqKAEvsDlkeZTRWhJxKmOzo
OkMVBbxCQeowj/YhFCh4OW6U2y0n415mPgJKflM4zIEBPPPg/tc6S6e4hSas8z3dFDA/nIJ4gQNr
tf3Rkeh87EKA8GjNyPLbtlJAzs32CmR0TJckNiWgnUH37PBhHdkHs0q4ORRh93HZI2f7EhB4vCrp
v/NQxPXIFVnOnpUK5W4GzjN/HiKmXKLK50tiKiR+WHoeLM2PDFibjuMcBZs/F/Iy3TT+/It6iiV8
xn3XbP0/z05mJZDXL5p6cV15Pz8tDsKK+2MxM90UQJfb8Jl0aO2P60jTTTnc6TFBYdwVs1L8iYoG
gvSlsjaIkpTplqdGbOKuIhDgb87peiksYDguG5ZWg3r72qtDHNHAJZYKKFB8z2qAfyALy+aqNw4a
Tg7aAOxRUs9ssFhqrN2T83g6m6IwUqXREO1Qn43VooppZGltWZ7YrnT4Yd3qY8hoXwtSq4fxW/NL
/gRjgHOPz0vf/GgVucmVoKWiIpmqgNYyFNy5ffoNQiEc95QPabdz+EzljGpsmjW5SVeDTGjW8Kd1
51ImHQAFuHbctMylSp63XRvFW6M17wzq3i3Agrk1e4b9eDfBkHmh72XBGf7ZbehKfO3AmE4MmaCd
NzyIwnOKyEH0BGdNkDPPvWvnO+bpraHTFo2nh2D8YIOT+3QhQ/5O+0gAI6qXnDfBJw5AqqwZSxSr
1LSkk08kixsS9afv8aXIQvEP1PZ/BGzaz3OG85b5kq8LlQAQjOfMO/zUfpxh0NHCQNd9b9Fsmds2
UhoHym+1E9KaKdSNGbL0E8GKSa3uTwxtf9tSK8nIWp00rJPXvak5dqAHhlG02mjtpSxFIu1BHnt9
WoZ3BAjZZhQDNp0ci+clbBNbsd1dVI+A69766/ki0gyqi06coyhvHhb4IXE7IsXIwP05tsZAv4lH
vLMJjIeUNq5XqqoZfJ7efKJUr7BnvuSjityZgLnHnF9yJKKuNx/BSSnM5jX6O9unFzJGKg/LExeX
gXS1mllb7aqOgxXvrJkfb5i9lq3KGi5M7LPn1edTccEEVCwfYQJfFX+DBxyGgkGEEDayO+Yc4REK
6YzPXOGXe3Z4D9OvsaDA8yTEoIN3s8OMJeGAzh48QuiEX9HoSJ2x1y48YqkVE7T4JnNbBsRw9Jja
mJvItKoZxcylfcIU0pUt50q9Qb3FjAEeDr34NacZZ1N0GKtzvlxxSGjrGlLaCinRhMp1Nkkzfcvj
yjenbEkRKiYM+Y1ff7Na4BP5Vm5At0cBndybKWUumTXNQWCMsX+gfbSAOU43SuAjRZ66D9Ji6qhI
llRP4LtUnv7oGMNnIRM9xqn31SVE/lSFwfAn2HVnl2v2iyrMH28t0VC5Zt0rvSPLrmnVS5uDUzRS
IuwcU8l23uB/1mONgeqMt7rvNp0VDkWV1w+JHKZ3RX/a9mTaFElHr0wIMGrXAEFjzaoiknrnO3um
WSFiQCIA5w5I1NBuqMVQdoWj0mUEDTkEa+1RS+JfRpP6rQAcc1m9Swd90ko0DiccbwTGG14pANa7
4BgZG8eF3YL8W6MmAZ8TBvcfvYqlt0yfxC0yP9IOTv++QPikx/hmLTPcLZUCKuuuGsQIFDoCTMfy
qLL/uDjjKqGvgiVR3icBj3TGWPjFwJojgJXV7Ba30y96FXbnnqByF8zKAFabo7f3iGtpx4tEXxOS
uDyEG2lap5sNfvkyvFt7UT7jqzoWJRP5AYnRXV9ZaJpGQt5vZUcsN+Od30nyxTkgLJlno9X4MJs4
do1/k6eCrrYqQaP9Gp/B45iMJyz/0bMkJM+zwMuhoQDFbn2KXJS86s8QVmLxfdvpbdLhw2CYD0ih
pOfzast8WQxFvKCTRipU9xlFzvjRrpz/J/7n/N0nc2o6oFT4uxsnkQ5wDboRuGxhnLdzV3LLQnSl
70ID65/LJSY3t1zgJ0Hh2xeziJHh2JEQybYqWTPiWp7jmA3u8++9fXB2cO8n+mTkHMpXRGZQmyi4
1Hn5AqORqYCN2eSqMykFoc9XVGqhSldriQgfCKpbj62aQ4f3WC5CX39ogrT24OL1Ft0g2FTLLewi
BhmkBnA/wXe4M0zo8KkVd8ZXugHAWPhV/31I1lff9yB1lcrW3G0ZQdIAyl3iz9wxqnN0Sb5HUAKm
9lPd6U2Ykhk5lzkFlFNd01g49KO1mr3/alPuCerjR1Ke0UDVceRbUTnzGcq5NOw2YDk4nfbzqh1B
8edyo0thMvEHyQV1EIFb7i7r1WeFLtbo0Ex4n9RNFuXtJ7Gt8TcLHnvVSpv0TxcwwGLQfapU0TNV
tibmy2W2W9i4R6PBuLF3utzHkpBEkI+CBffDrCrknvCqaGurnTS9fpEa+ED9qpKQeaXaJRDXlDHY
eenx3hKoPAWULhnQpuxxbeR5C64yv+Ny7j3su6f9BlS9X+cATq3nq1DuxW+rwyoDEOfDLRKYTv8w
WtaNlRDujbV5B6BEoKBKVVkZnOtYqMV7YGg4XZsnMmr3p6NLV8raYz/QGbsA2jLbxRSEqWUEKpQc
+4IF6R1I6BFQHbEmO6eRoBJp/gi6aF8F0O5YafT+nxbTaXMgNP2PpTz//Hc8TaFSUf7OlOS6uMGj
551icvcgSj5kL8vzpk/lCGNVfOZSND7iPnotuESOeiSXGv8H615r8RXbo0viqZdChM1SFfT4QTWF
66uNHQv2gr2b2Pm+mt8MHT2+kISydHpWjqWxONrgACq9eYQlGJDOFwIh17smttP8RTlR6cLXFdFG
ePzzNhZh7rTObk1bCQBLV/QTf2Sb5K84eO11/ckl+bH5IjUCkLpmeNl+hlMnIqrAVop2o6xo8AYS
xXRmpK2vJeJJ+actb54nFGxqQ40dagDMq+M6NQsvhPJUZtL74WNcVhaR2VAebuZDN2BaPl9PFW5s
XX2Zgh+oGZ67fPxwfA1a2v0fC5o0756lLsrLPyuSXWeRu1JnoVMrPFoSfha0YNm1aCiQ5+giru7p
YEhx2Az/GicxHi2VGMMTD2bkEt6sAgtkFjWP2VuU9PO7/c4cdunIDm65o/UZYVVxeJAPHskU819H
XBG7i8kPS9MfDE0gE8nlzxUbxYqsngiCGka4JJYPbd91SWUqr1gSfZFeOoC2G+kvMKhjuV4bjlQD
jTL6fgrOWFUY42DfgwDTvLFm+LgMZ3f1yrskSWhVBKpOgBYv1p7psUnZvlXv1h6oSS8laxpYs5aC
MNjcZgLhpTH5Tq2676IJ5tguzCV0HKKGcGJoUSQrR/aG9kVwUUM1VtxZdLMpVpobbjfLjWrDn9RI
EdlX5jBhVuobbv1Fvxrelro/2vnNYJzGTAAA96MV6HehHXjH4EYhBKtwSU8GCbhATrBS55osV3nT
dzUOQvQ02xTBKL14ITTXiaINz+YpJPASOjJzNGDjMscAPA0u7/mtsCj4AqORGVNXYSOQKjdzt7Co
oroE0NHy9u5vVJT5Nyf4rw1pOlBbwqaO037lTlKHHNL2oH4OfG/uUFyWCGsJCFRd2FRjSwoim5wL
Prk4pDMa4vw99tX6VuD64hcq1oiZAyNbOVp4ULr11K3pv6Mcg6Bgx/ZcxRQCai2Ol2BC17bp06kJ
uwH92J/FrmIHfj6xe/SDtnpFQ/f3/qKnknhV3bpemq1P6vO+shYLwuHMxxb/nusHalmzYgx/8lsp
Ug0QBvDAP1bn8YfFyNgdR6+8OfAIhAknmSIeiNUREOcAV8Ft3RPLfySG+hYdtAZMNZ/EwtRwroby
eHEu+Wh5ng21TycEjrtDdAWzrrQgxFAdd6YQLNEntasXcomt5n1U5tKUSEWu97ogOOBvCZXnFV+V
t8mhczyZf9oaLGYuBYKuQROS+JnXFlCiIZM3LlP8eULZZKdOpeosukvJXJM9UE8422B1AdQvRxzs
hut/Tq7b6JNrR40mgNBQ4SDWCmuFwr3g6Tlm2tA6YZz+Ewh/ZVxxG4l9P2k7ON4bGVtqu3sqKwqJ
9MWmnU7/CpxFL4DZupgmfVWqSJuhmlhqb5mKuPXzlJDuM8nkPk7vMkXOhmZYKwqrWey1E9IXVsIy
My7Wv/7Ns6Hxd70+rPQrSPRE6Ro1qzRb2cZksKZYOYP3Q1o9Axk0cKvXpAE/zmF/19kKK0Pax+tK
NaSRhZQgGsSZRODZjyoYU9qecx3tCfGX1W0CotNJAc/SGQ6LThGW2/mxQGv67wWTChjsFDBnZwUO
mGcPyrsN5JhKhn0Q3lKGQs5vfVwsLaSHDTSkf1K8PVihFf3eQbjIQZ1QTvvoBiEa7BBrAsKQOt24
OE32o6WvtGca8ENRmlNEvCfLVNpMJHXK98i7zrqiLfxVjwTIwfCiYrrbBZRhOigBGqvSZiiKHbvt
4B39cKCcc84D0EAYQy/MkrEG6sDuw0XrTh4t9eZ9z5qaoJVWmOAB+lQcQbIolyTEeHpTDry71jPm
YNdh7rVnGy2x/TFmn6veyPsd70dZP1axBUd4f2ynV5k+0BoYp5oN36lljrVd7Ii+ovtt4IyOsTEF
cv+//AW0cfBrmikNsiRekC21AdnPAJxJSCBF257fhVov71UQG6MrBe/MNTbJxYe7m+W4fDYZASX5
oPmr+6DLGtCYsMNonSqQazsG2sSoRBD2MbjGMAnYanQoRTXpmQRNpVqpEsoJ8Z84r52PlZ5gJwRf
JIJTmLFSHVd869iDgFs5yBVu+dU2hb61zLDVkI8bsue1TYT1ya5bt1DA1WvnokGz7KuIzJ9Lfy/4
wAmPyAv3Q0yYq7Tno+xjPhBKp0RFehuzQDZza4oxr+VOksNPu84Or9YXDuSslGXLPEP1D1F8nfU6
IApVvV8CyTDMfsXPnsTPkFEYy+YJRD00E7NL2iU4M223C8FDyqe2Dn9/7oANwg3YM7rx1l/78Prb
yyaf+vP9cqGd1RqeuPYtLzwjZxBlvJN2K+3LMOamt3PQr4Gxr7pFwmLMbgG7QdJPa7ulEACzYVS/
Te/CJAj0QIN+E6R4TqfhDLx3nhbFLsLExtCRl/lt/PrISBaPZWLCYoehI+9ayv/uJjm3fGvGuxDh
AvdX851QX80HIqSgqvM5aqdAeW73OnAHqxVP+/DOo9Z7bzw4mdrx2W8n2Nwc9AoPFNw380HgmJAP
YDGXbwVU2LEXhVRab6dOSDG3oNbnw/puPaRbbjbq+Oey1JTGDOrngP2hnWUjXYphBUZO7RQVBMtL
vtr6HEVAF6ueGFJDYaqccl8spjnVVobeA5F8zCkL9ehiUG+7ZK0MEVJU6bRFQA6iLt8oMcOuSUxR
5RUai3tSQUvI5zXmaCMA0IhZqOSKIQD02/YHLhskXmJdZP+M40GbBGeA3fqdPEjaOPDrshDIdtjm
TXIvmdwuwmzJOAg+/aVi9RKlR+KUbqtPWU3mT201ZCe0tFFEuhTSidrsdOGDfX+aYgY9luiF1TMN
ezWt27rbJvorpDN/MiGeEu8K9Az5rxu7NuSas4UO/+ZRVDlRQkbSNTRHyEM9P/gU7oVQsgC1Goo9
Fuk+ycSY7LJWMKIkGATMJAaBg1XmQp21J22ID8Knovd5OGjOhxx5+opB3Fg5KrxiFLjSTm1P0yqp
fyRU104jUvsnRfzjRnjp7UvIbkwmWbLPBelHVHo1pSI56dU9WlapmTfB4E9HI2QY1ZHqO8Q9uAwH
QrGU4TAp1rgepFeP3UwvSp+FCAHsmsQDTMRxPYtob5PZVsHuVUEp3/m3x/rUvw4PgCZs0+Opnh63
qXofSwOD0cCLg5RznZ3mPHh9vH/Vq4fsY/IEsEqNHTi8nmyQDb0KzOC7Dyuhh5u974BaBuMze3LE
o/VNROvPRBI05Rvh+KSJh7aSwm1PwStXWytSlEN1xiGfK+cch2JlZ9+X6Shc+3ZUZBaD6iG0n9z0
ATjsJcAjdeEoUasSfrNyAK00P6jqKRjEAHPNdGYtVn80sCWWIIKL8KqxI2na1K/171AARf0WduOy
OMbJn2dt+zscvLLauGPY98BL43gYy6s3OsSPPb6WDIcZgxxAUGyUjuY4kJGF4BNawbi+0MQx1bjh
ERL842LsZ1UTJUX/IcynCu2qWU7hx6Hj0jwhYV8DtvA9nfp0+7+GuCXUOXZxJtSj6G9CBcK6QTDT
HHt3KGcRAQXcHXPHyj1IzcK1cBJk3n+F+UhaponHzw/k9vXouHUTtx4SDUJ9B0ZjKcX+p/GDWRWn
Uw131n2Wg76UfE2dYroTQi4Us6cBQdOhOm9seXhwyk5jlWDPzOR901XoWBMqL2DBy7ym0Hl1X1jH
MAnXxmnBPYCHToQ/KudMZb6DFvrhuqIAc5QZn+El0V57dLbZzTmaLrK6hZQ/X1EaQTCCroTBuhZI
ogZ4eLMrdR54hbaex3w+IQNTfipg5jAJFpUCjs8SITbP/reuinz2QNrDCD9/eYUKXYLozXr05fzx
A1iR5luf7DvzhTDZ0alXfxs3/ZhZMUSdWoU6IfRg9h53DPuYc1l6fxe/Mc/vzsGQaxrIr+wmTSBh
mJlAMyd3P6VO5D/0f4uk0rx130Z2IEb9GTzvfuupNxFLvkm3eV9GA3pOHv66AeilHFBX1vVrR7rZ
WXQYy2BOBl0Y2eM746fFvV54UVzhWNO+OvG5EI5yL6c478piS3dsA6VFMfFD47GLfB37gDHtB5Pv
w5iF1zJcZyOKJH49jrSygacFQ8mSVVs8XwkNAc0jnlwZ7/uW2ucBQiOqr5BkWyNRduf32D/2t8IG
gCnI4vG2NhY+4yRTXrD+IssowlNnICWGScpXs605hA1aLAaMpFZTLaSaW1w/JAsdXTgG9UCQ9xDk
N4Wuw5faN7ZCcer5uf9p80HWdbsSU7eGFULC+24y47g6xbMUne+G1gHOXKmWIBWaPTIiH6NiF5LA
rsqv900Pj8/nz/csChxwGFpbtMAbOWFde0cV1oZCPxKlyF8Cv8eRE9TMmzTLWr1sNwHT6FK5YCx6
UwTI1+FVnFni4zl7wS0VySabi826g2yj4+5hsTfHx3252gnLWgVEz0R3nf4eO4H2q4AhXoniOZFB
zrPXIyxXfx7TDU0zTDIEsqqZQRPcweO/BB+ho1HQ/v9M55ryvaxckeWQCm7ixQ7rtIKpdzvKG852
i8vlUdA+t+dMJTYOEUMlDFcnItOt71dXkgJ1t3s4HO287w0UHcAAuB78h4m6Rse6c9n6wWCTYw7A
iasdIFJRwyva4vlKnRDMpoDPbKnB/3aN88qUGTnVy64h16dqa1FrWmzNLxxJtlLNSIuon9lsOG20
J386JqGfRG1N6t7jKlqFt8eyQz6BaFm4uM0u9Wtu7jhQNYaI95EolLLMyPBZ28skldTMLxNUn4gw
s9DESz5DUQMl90QCaqpAJMBwzGLOyOm6P6Vx602W5lWjPt/cTFJ1mzZnAyCyHm/B03vpY2wWadeM
JXKqOZWSalQ1rmPzvev3z+nvL1olbCdO7kgvDY1JmTWVe6pesjoYLiZTtNSS3dPBeqxxDTv9bx5N
5yclcVYo0k2HJrHNp2yTQipG5ctuAVtek7hqMljqhgPFVoxM6WWMdJYsau/xU5wt4fMgxZK9BIcR
QSqMfdUFt8DuzmFcEGyewqR9dZFQxjXLlfOY37De0PgBD4fB/x6mieLoFaaj/AuISby41SC0HTG/
buDZSPGZFELjv3ZvauqL0VFfLfs0y9aWxnr3+hQwFxogBKFbWx7Ntoe1dexSCtsN4QksNa1sKl8a
tHg47USoI9gg+/T+JdRcvjeXYXBVv9ewSEelgG2MB98lAaEWPYyLrak678uT4pC1QuqKYgBIUUTM
hHw9IIs4ca1qxJHtJ5bNKqZxF0RUYVh0/fr337bh7yqPgtaWu6FffBJfiYg7C5lKTDz8okvyxXRD
a6TULZAxjvlIdmApUp6kQwhuRgmJES4AStoZQ1UrOsEIMaYsY9p/eMfCLaw0F+abXTT6AQJrZyiF
EfAgjXsM9vI0WlgNQsf2xDZMIn2a4uKea814Gx0K190H1AJnNzVExrRSmHxwBgU/OKoU922BfIGs
aQBiPQWfZrzi6WhoduQs/gZm9eUnlweuXcWPOQMJ1ZOTIOouVjOdKDsaPZIt0xwwot8Iv6PvQK7e
2gDTBITyuEHc/kXMK65RJ6sD5le+9Pa+iTearfhH2CFsFrPp0JZnx0J/kTRepr1UvtBZ7YT1Z6aV
QYcnLJko6vXziN/Cc13mwPrFkA13qWDwVpq+UQGasu5DkXr06dBa24R6tRTjzXXS4Aq30vGX34OV
ZGyYyKVMzRZjQPA3tQ+vTkxU6l+za5Si4D6sJUqDzbb+csRk77EqAFvBYwXlF46doC67z2gfvAB2
h0pppDBzBP0GDLh8HZvI/Z7hshs9yojHZCVO1V892O9e3YjK9HBDPDL9lwN1fs0ygCJFZ2zASn9c
q/LSYLQZVgwWt76IbRarOKYnbtm7zcRZYZMk0bN7RrMcT03Y6tG+0HmGQABCTiB0SuLLtEEgQbos
UWe7vZ3WiozYZ1kAU4+UHZ0PoPCkKGWE8G56lK7uzdX9zdOgLatkdq8UiYDPT0e5qNmRICgVUZgj
F84e0Ne68Ax2y5NcF3bvzEUNiZeaZY4ykOyoZ69Y5bNWXx45oU2Lg4l4K5/WCumG5xet9vGH3kln
3Eh/io2nrESYrliBgXVlI5j4/yoJ9UoU6cINDR3pBcYTZEjTmOwHtJ6fRTj1mFYmmlfuTG2a3nVs
0pyBwCbdH18PHKybvrRpEtLeI8bbJy2pAjzd8ysoI9He1OSQ6Xfkh+0vqBxaxJOQ1SVfTFnB/RLC
O6PrLEgIoxhpLCa+wlCX+kkhVI0aVi/DFCzR6qDiu8zf4xDhA4nbKApPDxBDnN1h8VnZPehvTVmU
/GIjC3Jx2uiJMrNXw0RltPdPWNjs+wJ3t5qFS/q2dneTGcNEL/mpDgSQF9sgsx6nvyuf8Pn1fpw4
N8POoyYJgIJ/BO+sU5PG8KdhpXWGaRl51wcAWMAo/GQFGgX/LFkfPNs+eB335Qc0qhOEJAGXRT44
q0G2VUQ1ei9X6BEZjqmpyj8i7y6F66fDsw6IvADAtneQ6Iuiq/wlOncjojM112ldlKsdHpyR7NeL
mK3TsqvZ+wt23IiZHdLfWBBSd2jgZuOrK0KoFmrKCBPJR+8AsCo/bKrMHs5VPTpLui1globOhNSt
45Sft8+pgKmqqpLPc/7FkQcVGPdRUBo1dWUSxEj0NnsWTRcoQ2d82TD8vy5Qo53kdTZg7HtdEJ72
4QKSq7vHuNJIk/CZO2K1ar6Tgk9qg321l9UwflmAGWD8IUcVF8BYqBF4HwbUK5xHeJcmX/YpmC39
zqJsQv7fsPVFxEuWFpln+2kpItgRw8zvfx/53+kkslUjtWMApXQzkNk37X+nsrhV2iv9FpHepGnb
bgRJPFkvXM/fi5fly83SLIM9aCQAvTuK5ZADbDFqYZbDkgB8k/9XmZYevAn0LpzaIQycMAqCQfny
FyTiGkiITOImoT6A9w/+sDyFyumbU6OARmkFnYPdqowYvgMAtB3XhPQScvPPJwHbV1siL7lStRO2
4XZcOIjk/X9B61M8FmYujskO6cGN+STKIsl1CAaiEfxMijHLhcGGskKtHqRY/CopBO9DjF64qsd9
vsshameR7ij90ODr4n7QBWZ0ZMRq7aj6L0UBwkjN9S511O8pmoyHf+GyR+5gVorO5clj2zhMzLZe
AnUqVZu0JWDqaJBP5kPbyS5z1ZPMNAPHibjx8bz1KmgM6invcVyX/6UM1Ipjjc1eEnvUqJBlH4xT
8sEDjweA2dAK7AOclTBsMo1g3Q9yT9gUmGd5V6DHvTh3kMrcq8/rxBhIQp9tGvrJrE9yPax1t+Tt
rjjU0bj1ndjAkB5WooOp02+/tgVd2M2bBIK5uwhTfaMIjJgqxw06tjF6zyCT3CP1uoZLY9upyOjI
/m2+w2u1bielbfFxkHqtzx1Y8WLvMOGUppRT9KjZ8FzSeluHT9c4CdxkiLpbtPN23EmVNikIZo3T
fb3mAfKZBMOmayPxCKpbBvMo6++i8TlnJTT6FxhboOAaXV4v7c9QVAyOHdj2LY6HGT+4h9GxK6Hx
7orzCGMjOuxI/ceZJqNxtwPWLby/5esAZyTPxN6Rg00iX5H+X55NhrXsMjlyS9FzayqQuwzCy4yg
fBWY3ANeXPIDyjOHFlWvLt6H79loYC8guX3BvxwphTu0aYDZMBrdakhvqyvGf2yUTW6AwOuUXeWs
VYDqziiScuDw7Pn+QXFBxQTWJKolT9iaayMawHM4CIPLeSzxHA8OLY6R2Lcq43kk+EswptO0H+9N
b85MFNIf6t7HXmF+3mqnh6KC50ZtdiCboBuUKX+ONsJ+HT0i1WJKMCjm0/IzhHq0C6fuojKiGd9F
iJDViTRmkMZqn6nxeZDRWVLRGl5qkgaaaYdzaXwIejRPqDBwUHa6kRVO0A89/zHaZeggu6Lrqca9
aGWfi+nXj/zPBtdPrt2+eqU/M2GilvL2NCMEMtI27g/l4z7xOBClE6OgMxTt2tgghziImpqfjPqW
M43+2mZVzSfk+rlMaBZmH1lzx+c6hhBLkn4wBDajExk9GaMneJGrNurF43S4+J7OYOdjP463lJdn
T+e+6Zfkol+qW2HkuwtOZsK2lvg+Pt7xAnrpAv7km7z3sNTjrMNimdXkU144ww+ygs4bcnP2Q7e+
0fEoAOHnG/eMHFxYAsAvGttrh4CiRnbWX1ppKQomZ57biL7zZFFm4sfxN9rz51se9zx2DYY7kWE+
cU4hv4lAjqAdz3u2HNa/Wx9ACO3IrwoiKny+RUoaezDSOgCzeWFu5BJCWAFHa3jAKJ6kYftfIajB
RISS+7dYsCVBivZmCDhgC02Tl7fSSBv87Q3n7sNHlBstuBtOxnml2El9qF6H+12V33y0J+maBgq7
msxecUtPjgelbGZ8YuFtGiuAR41AYAF05Zl14LsJjkYCenaTY9NyRbO6RvWJkWoyj7vdYk3p3E6K
6VUWFYMfWiRKP/zn01WN8HRIAM1Iu9CQYBuu9BKka/xSz35vcH88ZzhTU67T0/E6CkZ7owcvoWDG
doZmAH7q539ZZ+FAQ7qqjcRnxWruWmpUE+zkwRrmzFjtlrll1hMZaAvAX1UYECSPsekIPnhoZkEY
pQcQmREpKZKQ+9i1luUtRkRtvFEAyy33ly3eWQHDu/y/Uc9RBKOKLueg91Zxy6MbPaSZ6ORHtI5P
mh7hQi8dxrre6BV4GdjbVBVLYR7kcGyMVNAaaAOHOjmLDKgqvTABFlY9yBoQ9K7SQPOEmDeM3bEW
pxEs7oTdJZ9xllUNBNDUAI8jzS6w6Ce1ITkerC7r3WQttDBKo0WXERSXFTnSfk7BV6muIQbk3XmB
S4DZdSbz36ewewNddcitd1dg0isULnkKeKS0RjShchAyO8I6GbSgsU7gN4Tva+X7PjxIKKPH1NxE
BIj0VuqOcDLYPDRF3XHY8zxOq5caZ8XH7bFUJ6onlXGFmMjNWrloYtCz8haFYD2CJMPsYTGcHtnO
SB2YEiVZ2GoVpl7LyDA9/ThnNTLZH/qTaIYA4x7ovvd/l4WRa+JoOVeEQ6olc6Okvb14ZyQTAScG
6hETQe9oYaKAFozP/BqO/CqBfTEQYf773Wev8DPYYZYAB1Fj2bpiqG5fbMYu8n27JHu4UWskcR/8
eexmyfPJDreu9EXiRh0X6GQgMs0t+INhtkKbrmUqKPa1aFOzsD93HSZWiH19ElPP85ruW/D4XTmC
UxR9ljzwSXZUUzU1Wevvx3YS+KtJPJm671L+zJnx7JhlabYpqqBg5+bQEyJRDLJljGyzI6dCUIHz
J5ktqi/H6fdGEPvSk3oWQhRMooKC05AFH3tUbFzXghrANJUE/AUvy12RJilKIDqaEog1EYLXRhEZ
ipIRL3PTb7XkJ7jeF/IT2/Ni5LMRfwE7TBmFaR35zjYZMP1CUXwnvAaZAdgDuLPscmkdxQVwLqqU
G0a9kvRyIZp9WXRZbnCixov21NZK4azi0r+ZqLzxrYBHUNV/46fRrBbp1XVJFnkUdIOzLJ6k1tBQ
4jl7dpwkQ5NUghTilm8Au0kYROZGS03RIohYx8aO46Vpx2pKmO+TQMnQE5IELt+r4Rd8vcQAoU2e
9utWMqK+B/f79P3MtGZlkXwc5Cg9b+BqF7+W0jNoLR0WCloX1Tik8WeXE+DdiHap539tYD3z1Y7i
pifBlJOCmmkEFBaKMoyQbhe5i1rPHoFFMq+7RtJJ57/9t/eHOc2EdkEDoktp9l1fSfOwybhsuaVo
SfEN0sIcOhsSD6NAoURZE70Fwh4Y9n7NTg4dcH6NSfk9XXKjZvdbenzjgkTSFAUva/laA6QRT84c
MCcX/1lpqPAex7Of9DGz94taOrJ6yo5SBBRm254RgHFooRMhOZSZ4/9+l4NpKhqgJqep5ssRP/Yq
4bedleB4GkLUbJDea/5Cc6AWxhz7T+8jLHRrdrqEE0b1Fh0zhAVv6bsx5rzU+2vAjhhknVKGGeYZ
nkcQsPcfISKVrPceAr88Ok3+BYMlNokK9N+ek5Og0Ue2Vs2+05Eq6vJmOznKl0vyUO6VcPuZtrZt
bIcym4676jkRwpm3gc39NZeoLTPLTMx9ICugVHdfuG3Pkr3Cr0sYiuIlDo+WXK9RRTqzD+6LIeSY
KpCuE8Lgts8pv31/oIF0kc1uGAJnhn5qTZEtC8or2bhNoCpge4SmVyg0Pq0TUSPDTWBZYryKu+Eb
e48uomJz3esAEfn1ke5tFToKFATjzLPUTD9lmjUQb/HrBSOURv+Wt2TklnqcWjstbFu0xfC68Teu
85j9hDLS2slIFvQ8ZvNEwTp0CF7RW2GH/aKsOrZ79f844F6bk0Uid2HjdOdsKz1jpKgkFzSX0UMW
Evhul6oQPW0/H+7PltB06s0YEivAWV6vW8nS98CcRzw4GbohjjoGEBNQZ53X9v4LOYNviOSNeG88
nohvLhH2lN4p/8JtD9Px7Fiw6OmRN88phDiTSW+DezrUO6vl5dGkc0U2dRCySSdd7NPdTC0IQWE1
QI9KqMcG5Z+sfN/8DfcCA4OtFAtCwX8a+fwtjeDVLut4miV9HOaX5H3sIW3uyv1ArjIOhNwLw8lv
tjRD7+rJuxDGgzbzFHxM97svnD9kOXZNCMS48wSHfghas1WBKEiyL1ZQvx4VsJheJsGuOZ5FZF/w
GlI9rpvuFdwJT4uxDpazs2JhThu0UeJl5S4Y2wPWaYohWMhnqzL35MP1H6wMfa26JxE7YEqiDUoB
AEhAz7fBefLvCIwjAsQohUkp60CouKqKU4m4OkSMOl2MTUDTX7VUbCYwtY5A4njtUWgZJNMG2NRi
c/LJGvkqDDBVTZff5gfgLUaEuGdIqqMBBHu33+nBzgbx2hoI469UcQ+UcWYVmZicOr+RazfcjeNL
+g6VV6qALgbPhUiyegaQO8kMU+i1tM874QQOlqQTlh5wzSi2q/s5jgBADSspUtgyQnJZgfEOaD7j
nERtMvxTQ6ABfGglFls/tk3cLO0sUYRFaUwQc9g7gG98qxnifizAVLZ8xIuMOKpSbFQgtdfJ4ogB
ExXZ3AJP3TY3Wca32CxLZBSK5Hm7j/LyqyfyIlCt4amFowKwP/96EDPEjMMe1XE3IBpFjKV97qm5
WMf3YcUDx4PaOmsKFlXuAnRHijXGT5vvZegybSlzIaW53FT8gEfNxSw2xNPBzJUSMbrRHzH+WVGV
1UxfWQ2Oz2MX7XTppjFeQMZY82gjKzUIG4ux0uAEYG+IJkNWh1YCchVtwF/YvsQKqdR8ZKq+mngj
xUXEeqlKS+ZGjzP30nFFsDL6j8jsZSgwKKAzPp57EafewPYhUM4XsO/KJmBCSIjOxokXU2r0zEo0
A1mvZnJhMEvNsq80wLJxoMYjIyPUu7cL/3pLUUpAjXxgTfZf3QH7ABp0pgn23hQlZy0DRtmH338c
iV/Wc0zugbdMzBQVThOTNtwEYtuHR3ejCRtArQrqst8PNos9XTh80lPBCSfnEJkckcnJGgdMedy7
iHrIWAg7K72WDquyQ8yoPfbtVq7dZbDLNwA48rfjv71VFfkZzv8Ur3UHDGldONetkXrSuqtF/cx5
GewshsgshaJKguzrYXI12Vt6KRnhWAkE3tXzkg1qU5/JCzlw+2//CsZKWs/IedoUXNHuA//xrpDJ
UNt5cAbv2mXzDPi67/eDOJ0dVzhVpuXtp5B6Q99H0P46OlbNMHLzV8puK9JfJvJtnrY4PcKL5TKm
12fpTz+WbJ6DNB40iZcpoP5XAgiFOFYVECUy2GStdOGjCGgoxwqLl3nsjM65/yMWXN1hU1mIqVdh
TK5KaCMR7SDMZ/KH9MYp6bIs68ZBwuVehfsaoa2PO1wBejaC4GBLv7IlnYchSi66Y6eOz1WmOEmN
4H2J7uug+D0MsJPDeIsJ1m0sJSJLkICJ65RyhGEI64uGMQlahba9VzSv7DgPFzKmfIG2eSP5K7tP
I8/5vGaJEn6LH+pEr0L4/28XkFp1O+6/kf2sUQzCSP/QxjHIi6LDt9BSLIYx1EfaImgeSZ1muDBd
i0OS5bA6AVN/u3eex+RIPVdYfriRnt7In02CIgnmC99SHQcnEzUDdmyXAMhjoNbAa6nc4fDsBsGL
6E1ZyWj9A5ir9MWsSiwDItgfLcgIeMERhsZZgbjJ61N4ohoAyBk6sarrt7G6nGej41KcauRhEjJh
WQX16v58NBHV3bCOb10eQfOOoJ9nZKbJAMFRYDxb/EZVM+QAJ1CAOoy3rDC4qdh7DArWcUqcEFx8
YwvHcc3lEIx3fvHek+tRe9f92aZRXOA5/zaRiSg6G41Dq9l1w+N9T0oXpA/UviRL2rBdInPF4L74
yh0QY4jWsFStlgCaJay6EBfr2Ul7Z1LFCcI7hCgkCmVnPnQykbuQzEq4vPaCq559vKSeSudbfzyC
jnonit6Zb43OEJi3qJxzUERcmDEtSArq1vnLiDUpisTx/w1E5LSLZa6iEkvj01xltP6GhER/c71I
iGZhIPAShKZmQNyAGR9I1MOtK4a4BrkkJq+2g/SivFDFzIg2OZmAsaa3TnhL5S7mJUN3FAHJ1Lux
5nJVaSn/rv4NkGvAJ4lSrNBMzcim2hi/e7rCr4iLIODVt0UQxOkrmWtJ8E8Cq3bAAjLSsoTygQYc
H4bd1kVBFsdC9aio4O6odc91oynuo+XizGJg27IoVijCl3ZqJtGII2r35aY6MQfGgxI2SmpIFPCg
ZsG9LsYaNKR0dv6q+522nuowC/xYjhIjRJCS4yTUySwFsgFFeD6hXqaQpoUGRaMi+RTnyGA8Yn0E
BF1kQYW0OZ86b1rLN/8PsPVrN9LZ1mHTzhjTLBUkW4TlzIDQXjSucpO7clXlOW6zq3mJiQJM6Xy1
C3am+qOwx4MzYisEAUhFs18aYl5nEI1Uw9zej2K5/Zjb3E0dtbRWesclsunAoMNbdtrIeRemxluZ
CDI2jpmsmjv9bT6FI4gMY+YyQasxH0XGZj1F/XqAJvYFqRLp4SvzF6MRwhaYxhhZs5v9WrCXxqir
aPa455WUFO35Qsv6k/gfPnjq5JO9cicm2ytgYMKfTbwCDEI3wL953y+Sdk0JxX1GuRM2ihDw+mMd
sOcIylUbA4iMLotVoK6hfI8XA+lEMu5adpht0XzjQzvM4XMZLTSAw3EtfWIzNkNkIeJfSbwD5+L4
bx83+b2nKZHyEbqVp83cFCDdaGAHB3y+HxUmNrBIhAcpg2EwogOfIsweXDerWecd8ziiAL/rsiee
r+4DclSC8vgbwJKDR6oNWWthswtD0Aw1jlf2agO20sU4jzOXK5goiYyWLEA3irdrQiy1xCBrRR8E
P9zrpfj+XiteHGblc+jlnd4Qr23n2iAbhYFpuBHhUYqlYoqiod7hPhw1ycDCCZKomEc/p3jT7H5n
/1tFgPBX0amUPqo3zFfzGWtYxwhQomieXDP4zghXOLSoPZtQLmT8iIYprOS0Hbr1OKKdDicTLhH3
ReGYjF7FIdVy0pzoXY0bUac1TcwN0rwPiaWb32kxzUredUtJNT1qKgM8bFms7Mj1yOn+gwh2q+7R
yEItPKFWrEYrzhTqpKf8hXk+vUY5GMukCTBrlaTRM3+OLHbjDiq2DQeYX3F8Kk3FYyu9D0haEtHA
JsXNMGKAmVOFyYF1fnYG/w+xHGsm9mM4IzbKs+l4H3eLTse+SNNQEAFihcnwVqn5GGX9cg8l1LAK
pHFtKojQrjVJDtzwMHbWl8+SqIa6MHGJykc0HyiPaW19yUJg2t4neDD9DFjtEli8Pm8HNk+NNUfr
aPsC2V73DHsrgGgnCpdrbcUn8xUcxWshD7DXeoa9cYljzUFn1qEX/kOzGaxGygoXVr4luMljtngK
Ki3hHAMTHl591CaVF2XQSyhazii9m2nemnlh6Fz7jb5FsEzGJFNdnBwzgHDE0hzNy9yWKx3NxnYh
U0ca8RNX0L+MSyx9AI/uomDzTazBDrmuK1XWuNncypi8TCsKZeLeEOMb6UkFpDFY+hvyvc+bMjxC
3CSKWCrRh8IyTVdeE9F6PYAOb37cu/hbbhEZz5d62VHpM99ATVU41ButplyYxFy12k92bB01iafG
5CMWgClxrTKx44XWuDmHG/R+iiCQNAWzvupx0aFZN0sWO0DUpDeuRya/dIGGPyna5WYs8kP8xeJA
Y+dt76CqHzV2WwU7T2jUHY8t5A8UkZei5ilZULdSvoQwwtnO/etX3Rc+GQHVgrHsaxlX8h+jvWKs
naNwF2HimWzGgJMuBqpU3Bm+tDQJC4nOlqkUBfLlhBiOnICuWdmWSAMV0z5O7Xjh8jD4T/3Ctezl
GLNoVTAJiK8jqfjcQ+mxTrQkH7Heiknpfla5T/upq/lyT4sXeYnz1G92RJL+ZsE2s77zEUCLo22W
t34kc/OO38bYsVGK68xvUXXlYwcPVymM1rsfuebhG30YagRuX/0D2/J4oBONf0cLIfVmOw3KcsCb
8TMBKix3FfLYE4W6GYRIU/UWNAJchGN2qbT3hdr4a5XaXzKL4V9vR9zRSXb6tj3QM0JjBv1FUXQ5
/Sq84EAzZAIF6bBTvgEcMxcxfjU00w2ujBanyxgOnFP6eWjqZd6ALYY1NwfSUgavj54Yuzgv6JOl
kWGwv79hPw0ZWOyzYbTAVCBmfdNsejqvihlKJwQK7G/dn3iym7Jet9cdS2NsYP0kD6iq+rhxbz5o
yNnQ6BdvVOcki/WVJzqZfDAp/Ti6AecNU/15GywDmtl8rGl+lzGRJQkEtUmgTw3sOsPE5Afw/ej0
1+bs/sL7XGyC1qw0hc2tbJdTTFu8oCIWEk5R/MXfUw1XjmJHqGSma1Cs3ob6ImRB3j6uQgusCzAx
q6xDFpo6xs3ckjREsaKIggC5xsz4VkLx6ZQT2WkeqhLAMPuYbDWoTxP3VbTgzd1tGlXdJlQQBWMJ
xen/35xPPB+u7yz7xscarEmVBXLiZBGeD3L2jkwCNhZXPJQEtexyo6PiTLx/NxF4cSp63WiHWqTR
IssCskNYs6GbW/mx/ZTk5xJyYhRpRig4OxwHDvwruO6QJR9K3Pnp0uA5JnNMu/lt/1P7s7Fc5hzn
3zC9fzoNhZibZFUncZrfnqz0C9Z6Jzqlp7kker3T1nW1QdovG6fryApDESmtETL1pFf0QRirwyn6
VkG0wC9REBYlKIo1DWij7cfXJnh15al4+cpyeVXgMTCGgXjw6tey3vZwaxAyKME/Wusp3po0AAkm
qCZCCKbbK7LDbQbCaq1OYG40d902ZAvJIZn28NmgGmKmEQ5ia9kQ9WxSJx/Pubu/Py8lMLDwiWCt
yxQUKFd5kTcC30Xt59u2XBlt5IwxzgERNi7LC5rSEt3sFS/eGFtIpZTVFi/5CKtE8l4w/VLFl1/w
8VumEpG6+Z0EAN3TxG0v4VqVhZnHWMOXluajecviMKQcXloKzuakT6Bc/d9GFcFpcoQpvDQpy8Mm
9fa2Pz2RrV8EuBAlQivlK5NRxrMVjYuNVlCKXEYRsC+gIz+zx4JfIrIxngZpEze0pG2aMrADbI/S
nP5Zytps+Tu7JpgusryQMtQScVk5zpyPr+d+wlf8LNhRBbSE0p3cdIJ3oC1NhPkdMhh595mqMF21
E8jPNRstS2i6X6X65SFBUKzVp1nNzucMfFWeZLKognQUnRZS3FmdgGUbzObb6yWdkFzL30vpATMd
9Bl/YGUSY9TKkSxLRC5sdlY5wNAi30f/ytgIHKue+6RvTQmQhI/L7BmTCRguVekgfDVSpS/5AY99
JlDZoe6EbPHd7o4D/R7t+jt9NooUbtl078xcW/JWK7TlJNFYCF8VlZskPeeGkBS2OaCShy/8B2oC
NIGOdEu4NBJfEb7jClCAMkmcrLALmLoqsi1HrjhugEFBByqErt0i9FtRB3jQ/WspP0LjCgGajpCF
qh4lIN++EIf2crlqYCtKWUILRFTeyDcdW6DGEDONPTJUGE0M5kUtaJUpwIazqDTfca+ABLiczpHT
6zqpJDBXlOmeLU3+/felrxaVTbp4O34MCvQabhy8qLC1N1uYh50TANjZOLGYZiC53NOd+YDsZ6Ip
ZNgsGMuk4RQyV1zzyEUJxN/iboWNqxJcJgNnoD/7SpqB7E768c76DKzY7Jg2akqvMqsaZSx3VbEN
bClp1KQhPQogwohKrWaGPzzZ6YRkY6y/HyRplU6hDTzSfBajrjs247o2Dx9bxmV6/juX3XO5VYpc
uUJwmI5/dsgiivZ2ruXFGhXLOqPe5lKgXVYsmJSEgMVhGvSWt7ZXyVkpDhSKYBPA17fS8qg+DqML
5P83vojQnp/fOzcqTpSpHkMTbZi1+uX9iNWTnSCeV9F3uAFf0GLLXN4RIKCIShp/qB6HfpB54934
iM/uyCmR29ojya0lZYTqJN/plcnV7iBP8nQzZUs/ZNACrOGnk01Pxc1nQs77pWsrfr9b3IileRA0
Vbg7t51BbBpX4WfW8TSZl0qm40Ckn/pft2qL7k6SxaCJEg3DKP8evKDilqE0aKbdJCV3SyjfYKNB
+CwY/lNBBef+P8kXeuDkpB1WcvUcJIICnHsq+Thznoi/FYjs5ZZ98Wsc785kBGlb4lVGD5XjP0Vf
tmaEmdMWK3szcbTOKpLM4DSTO/tb4+1LsRTrz6xMt915oaCakz+pesP3dj/ZhxZqluPcPMFddJaj
ZCpLIfSS9DaprVyUGnQFtZi7wv9SDymxz9aGks5Qwf34KEcWut801HrTU+MCkLWCIZnUDnHKvSw0
bsyK05FhhwpWbLWFyWbOwLBPTxNyEK91Y4eb3Wo/5OT+j+KnitYMNqQR95W7ZzhZq4JVYG3zbRIR
U+mZ9k94gpW06TffFsjvbKTAGqq7MN2PNfH7s0cYJNyk6BaijZSl+FkBmTKihT8jBzzG8IahI9gC
whN+jNTO8uzMk0gUXPKzAqHq3l6DT6Jg2U2Ti37EuWi/4H97rsGwygrCw9WHZHP/xIGojWvBapfs
MC0fvSOgoe6aOp1+OCuoAW+HEcIBg+i7hPyn15h08jatNZgu2ysiFoCSvhk/sJsuR4fFmd4J7+87
HGqmSxq5E79XJTK3RKr8fxh3OEOrSKRSS6kxVe5cAYEZDIZ2iL4W1qVop8fRLhv9jtlJlMs/+cBR
sOE8R1BkgSe70dgBNk9yMk0GRxYrJZ/JIPLawuBHGcLI2jkG3It9sNZAOyDyKz5Qomf4JVyVhdho
Nnl1Bvvycf+zV97er5hZn6oCGTY3z74PkphAqD7pBBSTIBcCATQpe6Z+tOS7t27Set8KZ4blzWEH
qom/wir7BM0PeYoL2goNCQTBDHxX+l51TuxOf2aZQ2q0rKfBzagUbsLBRKITCt0murovEeCI0TGP
9ecOiv1K3qpnJDfeCTi1uwjaJ8IzveSV7rtDfwobhivgy87Nyk+LVEuL//YEROi9pLAn2/tzBvId
/K+m0XTdUmciDMYtXaq99XohHizWA1gdM4W8oNb8RHgIgoSMt0ANTTA5cJpvYFnuEUe9NRl1a1e6
vsLIbr6Np7RsDvM8A1ouka+Gk0tPbYwfKNjSWIzTbeJ2Pt3S7wCnJ90xsvAUWWzYPewV8yjYRqd2
uxAkSuR8fYmsl55W4OMvKx6YFbyttJGn6O9/k6EpjlimNTpu9e1cHjvTnVg8s/yt6b3ll4C3z0ec
g0ka0KrK9pslqDt2AvMNfTisg7baqSe60pfTqef8UPuJtJ8s7U+Kyp3Z+xh6sBS3FAcx8aZ4GSQ9
Xu0iQR8myKFS7mc7wpTKeSFauuJRpRG94CCjzlb745k4xGv3nvvlKx5mtrtBLqG73zhv4pESxgI7
LeMv2ATxvz3ScG7yINaaKeeiyJKim0PnGjqeFNLgIUz0qpBamivnV3TJ0paz4KzqDlLZXHc4os5Q
lknrd2IdmL7vq2a2Cfh64bwSKO2X8OTF80RLObdr/shP0MVJNPCQnDsJsdTsEBzQbj8vep0aJVP4
gckpPlAXxEwJtaZn7qMoHz7aiy9T4Ffyc1zELlwmV/JtoYTKFSpikQpQF4gA4WWglIqM+Vwm4UYC
d6grEYXTYHsDiic/ytIAFziMPbMipaj/HDEryPCiOmko41i4OVr/Ohfvfccvb4DuJosAVfUj+36J
97mZk/MUOpOiwvxnWpJyx7hFYhsZfALvyF4xDg1zDe9gu7k4Q/Wux2mT5mWmvdVe5qMGd3QBJbMh
efRXqEbxih1kwGPfu5DbqNLJMiSeNxhcdK37Yxca1ydUh3wXNU2cGbGWJ2A0Qxu4CcW+uTA+12Be
Zcr64FUgIjU4SiPxn18z5nYOVPgRTdQgfFOJHL+qVlUuuCNt1lSy260gvu4EasvRryus6DK5KV2G
CO79cwp6TdzkUQa1nPTsg5805Mkw4b7Dmy8rSbybxSM+Iwg3G0Lc6PrpGprY6sAgV2cDzHVigIxd
LgNGImy2ERnQyhEGEkAO1x7QEXBAidsGJhAFgTxyN+hKecaNXZDJSuWzmPwzJ3pVaemQC/8aVlY8
44qW8I7y23WAR/LYPsL0g4jRyRqeBlxp5w4esrm7eXzle3sIHe9dC63Zt3OsBXkgPcikcY/35MNo
ELZd9oB12EgabUpDtdfG3z/A7oPDpLdJNQEopRKQRMN/2rbJsQJNjWo/EMZM4W3RhdakcqwqLecF
FxXlPRjlbLsRY5Lv8WjVqxrXkShoBG4hN8klNlMkrKp1+oL192Lwt8IQD/TWoxsjCYqzaY7cQUjo
Jf5DqJGsbiL49utQRoe8cXj1Ar9wlrz+GS++JrXmXdDqKNKOPY1CRXJP+XN5b/cVzlJk6AsMh9Jr
IAuHyOtHP0bgiPf1xUUw77BFRS6b3LXXP+4NCQLTkjdsc0tT2QIv5ABZqggzdVYdvFMVwqYwP9+K
7UC13lv3ESsyZf7U3m3Fj0lWWpEWaCqroZcr8CjFwK/Uk7/ugW6FA0cNAwvH1eY6nDqNy36LS3zg
4Y4A0/YBlrVAaiE6NQ/twaPgBdGkWHmh1DNN/y0eerLUwoGuInc661udmlNrl8p05yc4CNCsYMtu
qeL8P4GfIylnZYEeStYGJph/5HNsurFq5JtRFu+oMHn72vY5kPiX95wev6814Ae/WsDHkBI6LLdk
k3dkV4sRL+l9WEoTZRAE2ROn55Lxdmhywa94dLTyRwpuPMdc9YZ2vsL9VS0xeGoc7psgMqBC24JM
VdAaY5fEQ5tYVI8S9Flnkg4ajls/f/Jtq+CDkGmF1hNxAI9xE7pOi2JaCi7YgrFCOPCLEF1880TW
AIuTmrgEfsalxSW3pG3iudC5nfBcApiK1T00mxAYS5R6rRaY6Y6Ox9lqi4jT4fSAdwk6ohnnVbPd
+y6FVdWqFDxC/LJ5gWuJ28Sq6c1TWyw+7UWnX7yEucfERlXlpcBUoRmf34mCJl7+JGR/L/YWI0Nn
+FoKmAPV7KZxv6bioIfg1gsMHR9uS+z5cSDEfM3v56mqEZRE3hqtA0FBRpNihhwcI1cvh5fGzetR
KEVlZ69LwRePUHuuIwP1zMvTWZRRuLAOtSGsXFj/zRLuSp9+OjeUNVrXzyPrROTs1y7k8dgOcZEx
dRlgvcO5fqG1QB+DRQXJFitOLcJZ6QZSTSDr+6BIKzqKgPDCCcRnLOVgEqdJgnF0pIkv6ihFB+gF
RMNFPNAOiXif3jlBTxCADT8lpICTvGB3EUwlRMhqK3hSMHh08r7LV7qwTkS0x0QxDExgxSNhr5x1
aUjMg94vulWt2RkXp3bCcDKxFECIV2IVHbFJH83altRssqDK6AQ/KeC53d1UwKv2YRN8EP6AWVsP
/u/6KPPMn5q/rqBsrZg85DJoBi27A11MkTuTY+16tRzhKsBUWM6ALI66Z6jyZkiKxel4IsGWfTsH
H73XhM6RMjQoIh/c8Iqmrt7CQk0Ifxssb5YfKoVhX2l24zqScecRyOy3ug23+xEWYMuO5CtmVA5V
fyCI0HcQyI6IEEUlP5yw6knSE4almFBh89mT2pf7+38yF+R8djyRQPhrddMr7oz0SF9IWeNKQ6L8
D8f7wr9OfoiwzAzylAyZrfcHB8uflbJ1UympHHSS/UVC02TNznNY2aSwrUQvS9kmdeOn6BT+8u28
m7CvQl84/u7HSTebYo+fJ8BMLhrRdNZEwk+0Ps/ckCuD20WnCYBUL4YyD9IQJDrCm0d5E0GbQaJZ
TwhoqvLjhcN5PO5Hv7H7H1RG1zHyHL38MECdk8PN4sZ1+rG5E/rttoNvKc9cWeKRP5N4KFx0T2bN
RnjWF/djjVTPFAF6YMkZoOYDzuE+oTw2b5adjTy7v+T2fLpddMWpV0qa/Uh5UlIJnnNRaaa0lmtc
l0chvY820BFnLRE19aFTjQhDPHEATPspuqW/4GcNZ8Zy3U2qclaqmZvC2Bd2NpCqQAcC5OEPUzLG
tjhS0oGqRn02VAf8O8x6dgAU6RluLrHXqTtkhG5PfFwhKon8aCW3pMix8PgKtD/ZaYap/nnQ5aRw
Tufl3Cv9DJMpUTUDMoV4hOsGadzAPTupjXO9OqaozSe0MqIvHu1NIi8/x/wJDZFQKsS5s9z4OJXd
Kmc3D1MRSTbyBKom6vQZLQLjQvuDaTDwT5cclrEHthGQS2v+6Czi3MDtl8n11G9G9lMRlk3FpNud
w6R7IarcKNBZrv2OmqeRj51xikXKBRp5Gy/r2VWH9b7OfcNZH32ZwARkDU+wX1S1cTX9wY17IGSm
gpQODDBkWPE7b0bZE4Eh8YgRSj8kwLe72M/zi062ItjA4CFkRu1sn/yBZPHGuNaWdLiVPUzl8XJA
qI2+gXBuVXGqLrMM7mol9fNwRhv7ItOIazKmWha8r7Vi6rsvZB7ScIel+eJ/7t5C9j5CoaXmcIVM
g6dfcLL1fU36Y//GDoRvUp+QvPz0vXErfuNi5L683UqeAhAQp32FF4XM0+N0usleithxQtgga0ty
wTPjvhaeyjSCw6Ekz9A7XyELDpYpTbPA9DnmF41C82E/KKGvillxb4FDpJmEU0SJtCYpu7tcUh62
Y8okNQb9w9Uoq6UIfGDxXtl/CXs/VOV8LB1w7d/R+wXDOVrWh/gUQtqA/CcbYO5ZK38f30x1CqRW
/TVDSv2mwzzkxdSWy/BMo4SS7hsMZXLz1o4NFUABWIWXB0l636gXxcQQa9YFa37PJByRWbIPFUAw
nnd826DtjIQgXEW4hQb/zfI1A2cCr1K0SvdZkZVcSqftQcmjZANg6QIMEDB71SfADyUbsHerJQWw
e1x/d1I7QWppH7DR+xQFb342GS+xvmLhd+StxetlQpS0bDwgrZsx9WmAS+4fP/A2fdH6sYNTEAU4
NQuC9zMJOfAz1spqZrqqeT6qndshj8Ojrn1+3jKnjXaYHL8UPfZymUrsMQzoSUKeyNACBbs6lYZ2
AE0JQWDIkWsOIUilUuARpbsfeQX5NbbdrHoyopcfpiJGgwg9xXbY0a9cuQfz2BDSJ8wlzRosPejb
mPiHsBKuSXFXYyr3wSL2/F2AQWHCJe3C+JxGoInynvcsjIrWad4AVeEMTXMfTMOkEdnJQvCWcodc
5B6YLjT5ua3l5ibbGjbWU/O76oI0vir2kmzLUkUIgF/GKNR6OxlWEu/xfB4AUu8rnuQn7hhcTsXu
8hg4/qSiAwTQ6pMfNQtvLbphvNR2CTYHMAXMh8vWHZaFYxpZbgAJQq/inS54HphqWtDdfpeGh17o
l1hvrzvSS64idzVpvCUgciz1rhFDCGLIVYm1QFyV3CFeo9tbetpACFpXS+KyNcrEL8902Pcfai8J
3ywdEpt4KWoKCnbYvXytwlXzlyg8Iv1QnTUdZdVM1V8F8tVb9ns2waLXcA9y66KnLRtx5VcJL80H
ZNjfFG5RDj/cZlnSFph6g+z7IllaJkQRZaKoSjX5AA0VsUIt7d/JhkoMoKms6RcsI7vVNwj3zHBL
cGEQMhIuEIXXmvejJGm708KIyZjd52pP0EBYGpmeW4D71b8PPS/OETcjOt5dq9ebRWh3IoHFtBKs
AlrDQUlbmNDg3n+qP+d4qQqVD4f9d6f1qeTy7mn8LNHnO7T8cxHkr6AlVT38w1FiUDw6AxFzN1vb
xyHLUpHA/ZppSifggESU09re7XV1H1GM1R/sNdmsTbSLcNCU+YY3rM9RB8wWlA6BDDnAHQP84RPe
5MvZuTCy1A2yUD6gZ1U3EkziVcs53o+Z8GppLTCXC3fYR33Ge5mfi73k+VSYgBi9mXLwiIu9EwHE
rqNCq4nK5HiF3myM59qRtie/K2ZrCmhEw0cGqhcip9VZi57JqGjzEEE7QsJPArSrCTu590LvHv/l
mTLtrwoKZN3hM2KyvU3KqtLdLPgow0G8h03ORGbzJbwA0STjfhSLzi2DZT9/xXEorARSFQ8+ZGk1
5TsWI8IYasmaIEAz6oZU6pVKnPhgHBQKqvjL0hIMtE/E9dlllnbEY3cVu4K23Kn/siPr9DZru4TU
+KatYGc4LrQxpuyU5dnk5Ou4NqqtqRKMF75Q3gziE7zv4bS4xWClvVt66dI7vTvo0HDJucDLnZ8E
n0bD/7V8quBLF4PswHkJ7/7ziu86S5UYxBkzifk+mjLgHFvB3OZOgyZjy66BLKnCPalTptFfdBpo
VUzBou27Z30u6S6/bZvd8uDefmfvwQg6Zps9xxTLEczMk6Qy3pcbsQFdYGbgchFxdui8+nw//vxW
V7uAaocMcWzKRs7I4OX5EtzI3QMrI60+tovZLKXMJq5aX2yl6VKwjtxbCP12JTkuJQbhy1aBIpYX
cI5Ny+fsagYGilmYzkSTaluGLzBwWRPEsJSC0qP6utsSZR06vNMiqAvQs6TGbQeBPjwAZeiqUjkS
h3eOolcjxutok9c7kR5sWL1B/Oacisaxdt1tM6smGifmPSRLTILvHDG8K9J91mUf/PK08MuXw23C
DajYgycFRqvi8UMATr6sz+wO9KC7rQSvF4WyFgRRFGixUJiLm3gitkI6Qc60msvfHZH6PmIlfjKm
eo/5VMdPQ0Vhb8rds+bwU0lJxCnQ5iTTSGRQqsetBSSU2HLZo40NTtQdnNAuzlAAl4ihCEUQdy45
6s6PkvvVEWQ+6mFDEtC7RpdBm+2ZbaNsnN7ZRePDHVQ7UtRiCOIYn8I+K03RQX3e6rejFHf6p4FS
igxvsz9FRt5vW2YlL0ineYRjC2P+T2nvy/gzoU0Ozb603+iacjzY/ABblGs/V2IL2RZBQdFTmdL1
2YXqZ//rEmRjIyJwZr6p6Kg6THWREoqwdqtGNx4ItRIFtq5m9lI8oSNGjdpDPtLxkgzg7lJ5yqse
JBYtAbjBYxeSeQIT3VVKv8I6pot3VwU2ctMIT1yw/XXigoRLwQvhDige5dfVCI08XAHwmvqwI2MJ
JqHEQYH+zV/1x0SucPPqULt8J9WMS2/sS9mZZzYcqG1oQZ4BM+l2m5bnf7hdtS/gwU8SJTGuFVje
wbvQ8tkvBFlr/aob7/VP6TYAV6HHgrIl5/o6zYYs3Ryn4U20KzhbsCdZMpp2toeoQwOFOufHk309
86ZGcSBPtP5wF4YaNu3NcS+UIARRCeKrA15WkoRBiCwQ4k8UBpaoJleMaDF5bb3SlkAe6+F78ce2
/KC1HxC79O/N5XnogBc23NzWSHNjlcDeIYsIuK8+NhfNxz6o0sdQtSKJxALDC2L1AWZPhjCGrGCy
xT1h0Flg89HzPu26BjXHvT72bH6/pxsVBcCRCU9cSmKX2tg2L6g2Kk3K7j3uzrPipRhYCpBFrVvY
qAxJq4WeBVZbqRTLczNw+xCsZ3KqSe0E6Bf8tsEWUO4bq49na/FC1zlDHrOQx6F4XA940G775+Ye
hya48VSZmdVD6U/prEM9YDa6Sy1kKQNcKKBI4UvwtPNwFJiii7qalwrXWp+t+x8anyTBX/TKqua6
J/HAKRRVV3Zbt37mUK1x98OZqTyRcpdiyBZHMag7VepeDa5+p5LTC3sMhTcl21rEhKSi/Go6KBTD
9t+R/gjSBM8h0eguGN9uJj9ozKFR3v8HkGk4D1dASpDxQeCCI3bQwsruGydXw2tRynPOlvBmYgo+
sYkd9IeM0oPRFyYKrmvcHwAbfCJ/bIjGEDo/XWQY/red3wd0P5laWlNDXZWTSAYvzqB7pCb7dzSL
SMPgRNkci295uIejmRahUN69q4ZrKBxrSnNbu5OhB7impNyW0BcGE/h0+3Rgi/NpvCtlkpiGmx6L
Guuk67ldSbWmCS5H4GeydJMuuKKGSKFn9fHSmsSCLq5JZFw9NRLBIlmXf44mdW1Hv4V/cSaaIyJt
s2H+1qeJGSXWXNrviqsx6+r76bN2GLuYCb8zYGtKVozONzRFgpJIvhl5p9uzq5bREKNlCulRTZhx
SPlnke1NziX2IvCNEfaDQ25+JmO09BIOOPzU1Hg6G7qaCmGGwCsSjOzpwHgjpZtbUf8Heg56SVP5
XEpXaNcrkOpU107ntpihayoEIrHcwWwqpwTqRNoe50bqXxSNT5SYAMGZgw0THN8yR33yeRmtOpqj
XYu86PVUTjNQtn/BVCCY++M+hEdsIKMRgeeWcFLSrHKr87HhH7Y+pPhCOMfSEsSnyFNe4UddKmBl
32L/CvEqsq8qg0+Z4Z8rUm8ZGXpKs5mpDbEQv+AGrKz2hfm9NpD6o8z5G5vyGRKf/VLT8qPYfj8m
NaaPpHAy8cCqi1mohNbvbmliOsSTzHBE1pKNXZoKn2jCqZ2a8lO1XpCuMvx1SSX0+QPmsIhQR5eU
qIw/GVne1R8Y/H5JgHmNdDm2QXzrTI14NWNo/Zg7XxeqmDd+iHvaDgJCj0kw5no1UK76mrwd9uEU
Kw8+KN1/GCZ5+yt34Q6Zvt4Qsq7nhfHn05q5zCQk0AY6H/GpWLn2GMvmA/3nWQXeug/oFCHiRKXm
TZYjV2RsrGgfs0spGQiLneFYhjoawr7RfQIFhWYwyxV7JjqKHS7B/iRChMcS1IIm6LIx0079vglJ
96R4T2gEfcEnhzQ4b//ND1USm53+emAqpRAltlwvfYAPlgEFGm4lpZstohwTtaFMxHG5Hw/auFWz
CXfdBPXptLXZcezxOjMeoYS0lxvA0pecYgsufVZhd8yedhzCaIjOHc1wWzdUbECTNRiH2szTK+8o
3LZmgZwwpryoKLIN6bM4TX3qG+c1gSNrN24QI6yxIqyNmAZn+99lZakCmGB7+XAseSvY8N9GPVde
80vQfid8NgWvitkHwOm8j/UGLroCumd0OIJM3WGgwnAastsc4qnIB5ATnJ8WQeO3zpdKwExeI/rP
rewcoGFRpsAHka6HNHNmW1D2nsKSL7WDrIIc8FcTVccMuER6G0fSooMmQ2K/JizwcQxPj4F+WtN5
bd0jeEsp/bqHuzylhk+pGCp7IcMdLhG/5QEF/WZ6Uiqng0pCsxVOYGLnusTMnjgaIOpBhd8k0Hri
BnGytt6ZtZbidFf9aOvPFxtef0rj8KlrAKCyUi7DrWIaZ6PQ3BX0ymQFYjfGQVQReNIsifAeubTi
ftAaXyyMvi8ajM5sfoutI/t1o88wptIW+KrMbeEAjDAcUkbs8bYXacqe211inEJ3ciSVBzFpXLbn
GmjSJ4U0v2Bo/rnLRbC4ESMJpWWwtzXguGaZiV+asXtjdA2Iw4q/wpB8LP8mjeEKPCs160Tg1x5J
fNIa94VW5WJ9yr0lqELc2bQLvCvamnn+uEKYSmCUPqmpWQaMKFMYG+eErAo6fWnITK3MxtBXBI8Z
wl9mmmxEKSH1g97gilzmIbQ2F2+2/qy3Lr3zRIBloZmizM8Y1r74DAAGhQJ/aCDPJGrI6h4ozp4J
EIWZe0u/y+Dwdu6XQDAatVunswFQMuAqRPCEy6ifwmiY5FwNMT4g23qk5Xz0zcduQ3NaUEOzJo9c
ELKuk5InHRvPiZ9axTa2M7IdNyvoSW9LlehezLWh2ipmlsqG7dYa66uPygDaw+q/6s4JlxA1Tb3r
cpzPjeT8M7Ku89gWXXMssQwHr07MvGb3a6U2HENOxhBn2+nCSfH9kK1vcFM6g9TRehKAHCHZ/3q6
Ii5RGCWJo7YnxCHLjmcwZB9R1P6mW5cTCf4AMtInD24x/6Z82u76fgpsryeZnIRvBE0ezbHma8Ue
S5fb5/AkfayHrLf2PvAnvQusOq0S3CNTHER0HdRzv2EPdCAfQlleNm6sZ61pn0Aa29U03nqtohNr
C6k12PvGk42iTA6U4c+kYI7mglgi303HaHC2zkIrIImPPxpcTV1cJLOIuuQ/K9pdM/5j3KGIkvQ/
GL0EHKTdq23ejLun1vLictCqv6yCcCHPKPFr8xBv1ZCOxpVmdfZ6/4RCObT2uKy7z1kzzKT/MUTV
LUizRlp8vnA/lKok2kwOU7ublrNtFdcR/SLn9lFZJKwgnpnSxx0kO4wjGYDMuTkctUNw6GGKqVDN
FgOmWD7j7U+Op4Y9W+Kw1S2u3NlCedyUSBn+nXpJBSy6SoVxx2CVA4Uqnj1AWlmyjLVXur6cYXN+
+yU1qwPk8Y1dN/UeIUmtmrMRAxmnPYtV2NHZBLKEJuHJBz8WN2LJ2T9cB57G+zscdgG41tQX1q6X
jyHGy47+nMiQWAhxj7ZCa1F9boSPIN/w1/+Ipkrd3IuOWXkyAsYli3rLyvD3gFUNHO7ENik2Ypho
IP+Cbpjb74snyMRwW2JGTK54veURc/mfZ3UcOMkB/CqczSsRdQu2LYR9a8J1u54D/XcUp7m3XG0T
qrPh0tdxRtohIL7H2lepNgDJutI3bILV4QUvkv+H9yl7mNtdZU8NqR1zOLBY/iw0EEuTrfi9pekI
dhEPYJK050C0eARClNi1bA8iu7dRutRepla77iSQZPNNDemdDQMHVUt+X6v/xj0rVUcmZCstKhxL
/be5Rxo2P2OOllri2znCT6UsEPMskBl5wkGSaHCw43tzQoP3y84HlHV/eYKscO6kmCipNiHP3fha
D3aYed18TgPlP6gbmjPn708yt/ZmOE0VYvVSDfFRjTdlxMau7uzLZs2yal1h/LyFDHFaohxFvLla
R5731/mL09IsOjaI1+n8sYj+uNLtk5V8r1z2F7Yg8uB/eWiRku1PToRfKZaxdxJ+cYPh9v0dFz8B
YjSdQufKJSLti+HUDj1Rh87gB1+YRJYSSkiXq7ppCblManEHmBu9iDzqikJRgQDzsDcBmPYuc3qP
uJ/6S2+oBKDtRahOsMp67jUX8LxDE3NoAGbsfby3yEr8u1aDitMlAKidwXN22iw31QooDlL4uqQ3
T5fa0tYfvt+NOLrMOzmbg5MLUaFDXURtEv1DERRbM3QJzRCEHVE4CdId2lmrkc+AOcnmKt4YXQfX
spl52EYmvM0ff1u00N1JN+3TQZ2dEjS9anROjXz0hO4FehmNhYK2gY+kNlCKdNCqeLPVpunXmg6m
uuC+MdKyeTO8CgEhG++wwmiclfcU6Lj6KRuID1n74YEfwIiv06egCyfMY280uvkBPLX/7y/x75Vg
tC6EfW7xgtNT3HfmQzZEwvNrIHkVon2eQxl5UqofpRmNpmbMlpaVuohpU4ycoop/0f1qbIza37DH
ND/K7sMkfel7mZGmm3XpMW5zH9RyYjkWrnP5m0X8wX47jOw5ihJrfYbRaOT4VcCJYv1QIDCTKV1D
5S/H/7gUJCGSt1pv4xkPC8ElLcBv6fkV1w9cD7ZoQn6ZL+kQwXYuest0Hp8+LT//rhit2L3vr71W
KwVO8d1Q+k6HT+dd24Td0eE5jkOCwYzhY8dLSeyxEs43X2uy5u94ktmICLsn7TaMSc+IYNpP1r/y
0ZdYNBKJu2bhcgRaDD3oG1zxRJUMNmcUzezEw3QaOXlD8q58fjgVhjms3qHTUZ7GxLEk3NjIcOsu
JWPI+55XIPlhJSzPxQPw8FMYf4U5ipgJTtyPgm/tuSMJ1Uw3LJ48hteYCUugEpOcrZImZtRR9+uG
c3UovqvI8iHlo/RVhXWya1YyBka/LxmDGq+nNtTWFQNPWYmq7NigKa6OhajFJCOA5ASIcnWt2t9W
PmxUdF5Dk1Qx56WO63agMRwQsfrovCflVeptI9UBtPCh9rHWTuQJcu5YTABI/dVrApZoBGCwm2AF
u8aN6Pj8x4BetVrTIvXqgdVGUdV9tkdpK0ZlSO6mU/DSyBIQZihl6PnBERajjy0weL0LM3oqEhgH
50WDkzUKFKH6DVCBxwMGi/91/sOHOe6gAObGlluwGyhpp2P2XzzztxdZ88ClFEhdHNA4OuKm+/WN
7chVIgmbTjeR8k/9TxtWS9rPAE7kjp2fJHhS1CG59ibg1XsiXt1th8LCS5lS48XLkKFEJFVCy3v7
C1hjNouPD7JrWNbBx6n/2sKH+JNZ7AO8sqy2kqpnNXExK859XfWBRDMiaXeNhzt/7pAGdpcW1Rgv
6jDkhVqlvcEa9A2Bfeu79Kb7DaALccmx85GM5N/zZXRoEoSOsRCXDx+FA5GGzidWbRAQRa8e2RMm
NZ326b/rQ06/fkJ22DzOuHlowialnrjkPC8HWnpzecRmSF9rvTlsJcjVvlGVPX1cjkxdpi8oFHag
VXIW1IRnmghale4Ef4cgw4asOly/c6DE7Dyt+jXgpb6bd9BaofxOcrU5ROVd9/1QnHbl6hruHve4
M9QDuchMm/nk5rzozERMpYL8d/DN32W/GSiwcgka6tbEzQzfJQ7KkVDcesPhf0TRSSGpCWeCgXGO
ay3XA2BNSgzQ3jRiYpX9oJLUgVOmfsSi2jDoNtpZKxFwHyBWI0x/wNmDrD1A28YhJmTfW0V0Y7JT
L/v4VTw5An6ougfDNtMccIurD/UXeqDz0u5xoJqBT4Rjb7j0emP9/Hhw8EOpFjRLzS4baOx6KLHF
QQZlpznjZPUBdw/A4gY0YlUGAkrv1GDA13RBVTNo4/vkbwLmDVmZ9YkJeJ+9Z4jYtKIKzVP3wAkc
8bompkzmILQCTHzT75Li6Y1XTZ+PxffjI0Uy1cepFYjJa0j0Zh082VsBslHfGAFiduQGY5pjtSnr
7jj40Wr0mvVjjVFTUbXZ+uJZpF706VdWrroOrF0SoycXcP75qpaZdLydikXi1anTUr7S5Jk4z4Vg
rBIzSh7HRScGWXrXXlwrqtIblKMRxDFV2/MhPCsZ2BdhD7hj9xIIdyTnvOCuuJ/C73hk007rUwKt
byq82zpiFViqOyc0COXuzUu1R1xbDys7lLyVKnyCSG/Ke0rOrW8lSjYlyT9n2ZmwUDSX/n5tNO04
qwzQzT5Q+ehx86HFYn/vm6LReKuU7v1eOVuS3atN78ixY6EmbA9eeAxDebLD2lAcvqj4xcMzTZXr
Wi813hsJRg1fBw1S51OYnM3Zh1n8/5eT5sJrG56Yy8emgRBMNs9YdOGo5qxvqRpTqCP+1yMJlyw4
ndjl3XyVxbB08w80J9xx5TItiD22gPu5I8zLob6E3tAxG0HV5RIxBOHDTM8x4TQg0uh61t40QdWc
hAG9516KPcinPqBS6pPoojMJSxLOsKsguc82miLu08IHPK05pTsdHZOR7m++rJw1T9SJ3VMvHgss
afpcOy6DHOjuF4SwF9vORLwISucHYVtV0t1yguHZPsihM765LjgwyaDi405L+TLYkIrLy3ITxoeA
Pp+Htcu9edFe51XEvZHhD5ThFfJat50faAwrwrx2aaSX/BP8INjBk8o1h8WnBq8gs6FxymjSP3rJ
chXr1PIwirdlRWizI21M8Yp6SQ3trAveE8nnNT7n45UQY7+KbI5tnpQh1Bh1VcN2Qh9HwJ9dZKS9
c6sTJCv05Oei5WL6e6ZLFZzlA2++nYin8vCshfFLlkM6AJ+PhQSkXex3LQF4v0X6W15/fxSnBuRk
Q/sIO12QH38a6tkdRKa4y9gloWg5YK1ZXMrOo8yEoVeIufUecEvzOvrIjkfEL50L7oX4uqArQhVr
xvMvT0/iwrvFtZ8SVKzwV7wL+fzUKf7xkJRglEWDcPiFaTkG37ZbHvW67UjiDenJVXc0VgCjLlta
2zrbjCedrMlG+vdQPRku+aG5ymsxbSVLOIyuiCJcuvxBMP/+4Ak5FezJbALUNHl8xi0csuHJBXz+
eLNyI4v/W/8zi/arc0Z4Kbz1i0Zm3Yapfv9GWw4KBa+czGGHQ0fPY3wVlLpPolb/y4q/4V6ZzOl/
iPVpT8kEU+KSCnHO/WgPLLiGRYZfJzdrJEmgrFmTcDf7qmjnQoEbJ773EwKc5RANcE/A+2gQ4SMM
nIe2lEVFNBB71W3POzyfOW2CFH3iyQRbHBrgF5IntbApRhPWcMRDItTwoLlDeLMKwnZgTu08s+fN
EsPobxy+75xHTY6hA2EjsKrVIluTyZ/10zyw02zmuzuYYCBBfVPGHFE/MAPomX9U0R196Z0C4qKE
mk6campXKvJUHxyvQzivd7ySsfWx2l9NN1D4SK/2QKEQXpu6GwAyIqjOLmmith7ULgQb/jTd0vJH
N0eiU/RBI75Ai/V0rwrvc7LmTc9sLqH81H7bKTnrNVTNqRSFGKCsOlv+vGMe2IOPtWR5MuoaC3rf
XXDs3lc3a9CGIEkaJHsRFOx//Q6Uie2vP8Z3p32K1163H6AcTy2suPDUID+pFbhhXZjes9bXfWzq
0zsYJLGx6qDRvVx6gJh6inxlTxEJPxVKdP3hEoNg8jSl3ilpqTHlhSGr0YauTef6GUOiDcCWEz4y
Czq+vwA6IrDd6qEl0pMTF1KBWYo3Chx4SOZlvdw4wLzNRqXnvC5RGQTS9k7IqiHx91K6VtD1W5Sh
JZ0rb61IiYRYANeyK3L4mH3DHP2wbarimWb936+QoV/Oci84m0UiabWNLi/KFw4F67iEoCLHNVUo
l6eRm04eMDpFJgkg04630nhA1xAj5yM5UHID4945kA59h2QCG9rfqBypdGX1yGG9C3+ShSx4mQ6g
vTmYlal+VtMOi4ZptYTAdMzJ1RyDtJRJJKhIqH3eARGLe2HI1Si9ilMOns18xi+gQOCrzps0BHUE
VteQzz9NE14sfFC1oSHs/yYINu4CnsKkMsBBS0jdjM9K8SzDu6mMQNriKfEv2mCJIbJ6BdqAVVNU
fCJHxsUeIDAaVnIfDNWbKVwcKEQqx4S2XdZMP/DS33AUMms8u7lZz5lpy2gI5xOwkyRwqsaCjlYE
rw84ZoAj0sfIqKWATegwczIkhyGejsj528G6FusTiMXFmZUFRmAeSyMjXy25Gh7UEZX+BAwUyLdX
8DJaeOBrBywn2Bn4/VkBp/M1gEJfYUbhK12TO5rdUSRHOFvUr7LLu9bwCKAqyCSVGdccFgt7GymQ
hh6rT4KsZQvf4jRN5p/aImEyYHYj1BnLpGXKHJWQObdYV0MdzMIRzi80zi2aCB6YOmocwQTdlOY1
am3/8l9ob9w9eYv9O7fzlCYXT5JdnHZlek8T3FiqHPaFsO+UQ8PqBFko3jAurHWna03xIuaDhZKo
bSjRXNvkqFcn1bMxmfj5xPUK1ZrZjrlY/Y8bd2zYSnLu6ElAacT9Lt/y+OVRwnPsivoDDgcpxNDH
9msjC2s6U5VT2ybWbWQWadFgE69gYwNpCU5y4jZRQE19F2BHX+3L4N/mF6tcuxVPyM7F3XbA5rWq
Q/+BpPPiOBDBzaHp20HqT5hn++U6HLR4D9yMjtLseCnh23TQiRpO0eEShcQ5/aGwU75KORKEyb7Z
bf34RF6sP8T3+fwTIzJvYaa/csE+QHh8RtyNKeJJ2gooynBw3XFqggt8x7ZuRM16PBPYP8mwjsjk
SQtm0qv2L69s+BdHtcAVd74YQtQ9PwqvyQjtY/DpRLRQlxyUECtG7oiDluYGJ2mrwY5YIwZDEYlf
3xSPPgGYunGpzPlaVamks7jsazG6VkgCqjFH5zYF2u7qPFBZ/zJDh/fjuexEnsK+1i+F5W5G5WgG
WZlmvkv8eH/oD9UCTDBFgBbpNzmvZTdaChAqk1cTUM7eKD5eMcfluBm6yrMxrsZsCTH/b3/btWAD
8jelhcrRnLlntC8X4tqYLr5anZTVRCepp6atauCyP7Anfr1olLgVO1rAPqNYdgzLZGNwc3oETaTH
2R9LSEUNvxDbGbHlvnQb6pAj/AG1fAHwaO2t1Yk7AqwzaoeQ5q3AbPO1MGWNTP0/objWgH4nT35Q
9hClT6CIpy/9A13p0KSCWoEMysvSKy2zfj+l6s45GvzdcVH+5F7MA4868QZU6tmRuEyN4IZeAk2E
ndhQGGse8PJUiRoyQmRt3hoAgAvW7Cz1BEIqxNqKGiDdYVqOVnPPXnB0KTS1oFElKYEBWyl6KX6u
NKDp4NRLpit3Bs+UUTnhkEAKW3bPjjn8qM2YuR8e/peA/oG5hu7gIyLWo4GTJTXDJpQCBJo+sTOh
hX0BJhdsEMA4kxH5wP3s+fCfPLsdBY9pY9mVpjitVcR5sjBMFi2WTBxvycRTM4A2qrqeouwe7LFT
iINh3xfJLpEunr1nRPYYJJUlK7io0lSxt94jK8F7Eh9RBlNrUAKUKtpKQmYuCe/o51/h40n7BKFe
6IQLIJcxQV4pSHyHE+bGhLp/SNF8M4CRQZ8pJNQk4CYJ5p63I3Ql7ZYIzpiJMefQK0LJiwwJgnk6
QziE8PjGxMPxu6hmAdj1jMWo4ObnTf0ktGSzL+7GdieWaMaIp0hqGUavlL+ZA6D+5yuquhol2AiN
XmHr8JeJWqj/n70Z1DplAI33UHE7I21mYz7Gu22BDa9eMwdA2hv+GbP2I66OH/UGg+H7e+V45Qi7
uYcUFiUsKjeQj4LdMEsHMcEfqmE7fTo8LOuvaMqsbpQGLquQxNyCu+dtTMa10CH5uXbY/yZIHFWG
F08jgT3fQbItmrsHU5B6YQvKhiCBQFEgEkF5S4cxv09RAptB6nqqBY53hqFipWO3VrPGEB40Srhc
YITY2t3i07c0Il6/8SegNSfbwPJnYMK0CwL0r21edG7S9iSCs/xspfqwcZtyIRWY63Em41xQaAO4
OF8QB3Qdzncd41AErSRHST4huojwJ0gS4B67n+D97gUxICn78+OaYz9TKdye46Yn/UBsNc/4kRip
34kOl4ath+GxtQp2nP3NdWusxXCwOe4EjAJq19F1GoIwgkUgvhlFuUrSm74qEKcFYSiC4l28R6BL
JYwqtWvy7VbdHBeoGLirAOI7KqO2xJ5D65bpUxdF3OzURzbRzYGkC9c8LeiPoio7keiItzUUpLg0
4S9BMfroFvqoeIAAcy0ronnGuj4VE4Lh3JJUQX1FmRwUBCAtMPW/M4b/MDo6ZKK3lhk0zeGPyguD
+7q8/6sUUzLIUu3gXkYATg3W+8b98Ys4LV5NMKxNZxTui9lESx1LKQckG5HLiXg72//QrGAc5kCw
lDl9O054oJJWCUkBT+fqXjiJb+339xCmFsqevehlGZ9czAFCOP/loHf6jBRACEZHLgaazPf8viUg
V3ZZaXZXTGiRU8YyWPEJjd0ltbQf5Tyc+fNhbT66nTNbp8dSGBpLS4Qlrf4nZmwFbkHVcjlrrdD4
+HEG5+WX5RpEvXUVGuGeEzIXEPmu9vh3QAX5xXrFMnj3b+qjGABxTE8OZS7AL1iIugb9gY3y/RGd
eFma+v9GY/2Rw+opfyk7L9iYScarZ7dSGM6xlIUerR0Wj5KBh4xqERfU1/fVeZvKnhhadFImbxl5
RzMtmS5+3Bd8sflCfm+DGKnrp6xbnr8jSu9iqnkIFhUn8h/zOBZZV+C435FeGoFJFj9UmZCKYUsk
yrOhCdGqSkKKfPPAI1t6Z1N0/tgLhX+jc4WRhODGKzj8U6U8HG4jlBrteO7XYXTR/KBGWGiVdBMz
q5gCmtYZRBbsMMQBUfEus3DOOw7qSs5GTyOaKRblj3jw8c5xKy/uvPKOLecCd/nO01shfcXCAejb
4Ra7cSjI2tLXVziU1uNtA90NeXe1Wj2NcjPkw+npN4ZgF6LKjXtLr84659PXdWDqXDpv2kdEzIpL
y9paJvo8ALJRSYL8WEGMZ3QqJrifV6AhCuRvSQLCVRZnD4cgtTbdiHqQIP0yhfZ+ZWrc6QmkENWr
fuWQNS2WJMJWRnST/BYzlz+3JndV6aGoSAyNT4rksnvRpNeDajUt3DVBZqs6mvJaYWS8EL1XT/Q/
cmErY1i+4OGGSMXb6oTrZdo2Q7Uz3yOWYtJBxf1vatdHWP3ARpMdNj88LGPI16KvvcvlYJnI7mVb
ce+P/sZFhm4Zqm/2sMFrZrYny9fYlMuRnUr/08EQgeeptedIvTG8kyJcW/3c9lDcr46Fu05pn/Xd
3KhreYDuowoDGPKQqK6Z/Q5e3Lnl7IwhqTqr9WNTt7f9Y4zxGFjrVYiz86/6Iu+/04pa3K9WcXTb
x5tudBRB86PWn19gkaH1HMfIBKKO2GXPLAAHDTR/yIAsugM6NQTaUvFAnF9bZzGYPNSt+Kh4VanV
8f0lpQGgsGK6P8JjCbK3ZeQKduUiLJYozV2+VSxr8N4m9/t6KnRIlt1yV3leuvAlx00VluxUoqEY
2t+e3aRGasyX5Wt3zxYnyXA1recWkaxn2zpKwA4AhapDDCoJoGmtY2pdgtVGHx95cDZTraBiy61Y
ypHwKWFh/9NHPI8muBCuZ+1H9qlqo/Y7ihT667udMRZwnJX3g0On4oY62Y9t6nnljSRNxYRVCcwZ
fS2aYg20qzrEcabw9nKfv2x216qNFhi3Ojab3pXpi/aFAY6ts59MliRMq/6shPIp0o4v/wJPQ4Pc
UYzxRLcvN0wcDhzrJgagmyt3N7KEZcn/jCMbUt1h60Q2PKEhei/RSch/NZtSLkOvVbS7TDHxFs2b
LWSSSLxQCDrRpTs/FWyLsm/nDQMlT58vCWib8eQshF3Qhm1lmkwrn3BS48tp6XkE0tzMd84sR6z9
8HpiuN6EXeWzsHmtTBOi4fHH3/xQOWZXC109n//2+mGpMWm81yr5MzLn6P254d2NzkupbKnfo74p
1YcIwzlvr3qBA9sBBxQ3Ne2owUMBnSCdwMq8B1qWPT6Ue2p0rhRGFcsJraESjaChMY329Nrq6+Aa
6JgFr8ANLbOQx/rcY5XPkcBysZ9K9/yrnC4uVg+knMX2hGeKQ8V+0kwJ84pVRjjt9kKcXmf+NqgA
gL5rf7crptaShhEC3kqLgWcIrzoAEQrjqbR+gK0DztjHQch8BqfZRujAj9ILcMSA6JjmfPwxMWiQ
Mz8uDrgoy2G+tlkZ6tZmJ3Xwe3tfdepKuJ7hC0wTOqBFv18mUt8YwZ/XXoCV7dssTpgyM5YVePU5
yYjjClhNIr0xieXqBC6jaEOfc26aUG6brQcam+7jA+gdkIoPUXq2EmIXtxxT7v47hVkO4HCgpz0j
T4S/x7Nb/Ej398r3q9AoD5q+RVCm2JMpFrasNnUdd+Arvxk5o++u9paUePOzyDCMhiAmpNguB4fU
dc89jIiCJlNeSFnUtju+ZzEG+yvT06q7YQLh1gFNp1z1D3KfdLcUI4Zn1WlJNs8uuuM42fgyVR5N
ls1ahtRGFriQa2fs3RU0nQ1AJn0a6lRwRr0pUc3CiaPY3tPd5DNhpzGQrhC1r2Su1cFhMUUIU18p
d9vNcK4cA5Vv9GekW8WJNU5KhYgV4DY5+ejgKzEjsjVhBcx/JITzHFwGo+E7TTLrOeeoZuwhY/OL
BT3sCE7x7FkUlIrwJDV2b4OQ25gVA1P7TBMW3pu+gENrToy8udXkx8h4gg41qbiqBNKtHSdLjrc2
f7fBnnwBNMzi9tOCBptugspqbwPv/USUPr8ZhbT7L/2bByX//k/HN8T+rRlEPqYi0Q66+5wO19l2
AOjnFtfz4VIhaxJZnrzdhLmzfZiHLRFQCPevtPnV1p4gvk6fhg5ht4clTwLsRbdIrGDY5Zv1JmHw
udoTGCATZi4k395iZEgIZHW09fnJq9QbTgfluT4nUSI2YfsZKgxrcrnJJ5gagjOvpQFRqnojuBv8
jQgtse7NlfkyewuZO0kebkquBUXx3fGWvJoy4HbWPB/RJwSShvjpFome9z1xiBL0KHzjzwuoAyPs
QKiKLUT5gpawJnofwNVlwrj1hgBw3wnVCSDE7KVYtDkbeoR5VIJdWANqBoTqzSdUCxztoKeAZE8J
ad/lbmJ/Ggt4DSfJG+vNh5VXancMqeM8+8q1LFRI55CS7NMzXV6lkJR1xbWpP3BML1TYwdWrdxuz
1kBuBX4kBI8nZIoYPM4FlwFqf3CqDR+vpiST3WSI9Bg6hmiP1F2CF0hUj67R4vcK/DjLyhqfJduN
HAXXR36K7GBSOJ0hb7elVsTLs0BK0yx6jAnXnJ9UJOUsRwh+Vb7PHYbj2a3xsyeFuldq8VBri3SG
oeY3lwLa88J9KkkxRswl527AO7bXVQMgFSsdJkOE1FINbGlgpgXiIKSnqoObSlmgiwzJtgbdONRu
eHGRJUlXoLkfr8XVXd2J2D3Ikj1aaqhWDuTd1Dw0HjQCYlyFzLqwQEp+NGSg2UoX3UiYJpudfWBi
Ht2xkJ1RAuXwzjh/apNRDnOxwM+vFX6G7BFpdG94pJz02sI55PFEFLMll7mkoG1C1iMPcAT9ZTh7
6FGNHUk0VA38xM34ElkZK5oFcyU2EFLvmA3kY9WkqMt67rpPqVYHLdxqunI5DRyYjHO7foKgYtwE
VSbFWmFUa198Aq3aNR1Hjbmdbi7K/UActntitADbLlTwe8Bz97+TnJnjzrcNzI9GHUssxbMiesDE
CI8GYgk2JBXxboVUI50arWKu8gBFa3qJF4iPGumeEXWpA5Ft8FqxP1x1udzw+gqyDZU6gR4ssHin
4KTfefitdIK9StMx7anf62HN84E/UwCnVkndxPcD1rhjzDD2u06hxs8kXClDaQ1fBJz6s74ODvzo
qa4USEe0f8Y0hEvo9Bl+LhMJismosuGBDa5W0XC0Axp6GI8qW1kvrcXNlMwv8xaUnLVAvPLQNGkT
Ycygl25kLWJy9KNREF4zWqzyfl67Akd731urTI2xYTUbnMrR1CzX7RcDzII55bCexDQRpiwdbxPR
DPJFFFVm1QzEyYrZUe2Cs24K6sXL2IwewnZIRgrGboGMLGUx9fWcp7wE3v4M/K1oeRLN/C8E+4CS
KfOUxHzbk+0vkY2BO04+bynHnoLMRDukzXjsSfSW4OoSc3x+pwIlbXjhcwkT2fFiJqB+1VC++suL
HemTLbD0vKUNjIKiBZ6aBNOiwLAs4gxS2GzJxSKgm+48w4MZyG5AlVF5Yc3n4VKJlHv2j8SOTZZW
yM2tZsurHlvN63XACyjGLOot2qFIahxeBdm+I09FuwMuyq2gPfa79VlSPlSQvpORwSCdvcZrHRq7
/KhgLpx8nM8p8Gv7yI3rhHefSlWYlS/B/bb9pmzOXxgIVrJfVZrJk67DX6uQNR42S6VI9FHl92C3
NcoUmEPhc/GdF5C+T8gnV7SkTqVTCa+p4DFO2L3r0kWyo8oZiSIfvZjwG9h4bTW7nqQkHFPUufq9
+/TLNcX2xlq93bZLnWUeQ9XktyXR2qh2rnEoAuTtSbR1NZf7n6zQ+HirHp0iXVUtOqrBp1+4Xa/E
8KatHJ0Ss+VQE5cNl2dowRZdY2PVfk2hqYlGWX8ZrQ4eRhoIX8QmAKCm5hZTEWC3BR7Fx3nJtHwo
TrQGnyyReRO8uqtY95LLNB6JPas/ZmZaiAcsVpiBEzEEXebCuamdPonqdVZiCErfbIRXFrKsoj3g
lMrHa35qJQENT4GoLXOZ3eZR0Dr+uKs1j946bPEqSvcoLreUgR0RFEzQlwwDSJfvB/CC4RrgK+dQ
L6dI61Gn8CilI7aE3jLV3gkwvrtaJDymCgyD0E9d21UXMAHEcyJRElh6WiRN6tUK8MvylCsmx+8U
xHowINbtzVUIDPFrTOplG+bobBwsQltxb/RYtJcyVKtrVLVElOypENxcOPQJ9u/2U0GscbjR84H7
RlkO4ujIkFBi0/vfrNvMBJnFFVgTHEqHlmeM6XV1IRzrZKBLEFwMn+Gea4lez8++sI8IGmusGNys
P1NzyXOoZ0WqIxl1e8zL370tL6HaOP49/+LH6ENaoooJex8fN7ACHtYDL2L+oe9WNkm6Mr7uUSby
zUaaWFlnyf+1B7q/4XRwf2sQyzOv1D28miPhhxL8bnci4i4LcyoNblRR/VGKvHqVpkAPBOdLs93e
LBnolQ6JJi/Ep/tHNwokCDM5LxXBInaqz4kGSvCGDQGZxAV5YYl5yOYQAhxox5agd6HIAmS2v0cp
njdRI2+Kr/BHFTbcJr5IpST4lO+mRs4U9wsZoHiTbTtGcWqG2NNFBnu9ASQXjp3fA50skwwbOsj6
3ZNzC6XpO3VwTIJejuSAOBdHORkgUFYPgICYiS6zBLyXFGfEIx57bOQ6mrqDB42omtfcc807qICI
hbmzKyhyX8NjQ0mglZB2EnOXK/vEjjYzwit50otQxGdKkD2Eqq6KFXxl6vaD4tjxXw3KcBGnRVHi
dDFrokQTzpdhEFDQTSPFTy4Nw9JcZlNBbCseljFD7h4wOSqI8oOzhE36GAXjXaqrQRW6x3D2VauA
SH16ScY3n9lN1mzMahKvfsIC4SzKJo0flQh7JXHgWE45PpW2NN35CU/uNtCK034jMP+wH2L1BNLy
tn9D+7yKAushoBJkz4o+77SlctL80cSA2pSPqmslmPxKP6EPKCFTkK0DOfZ66LdT+UVKicd2mojF
vQ1so60iY4VSSdI746wPiavjiioKRpPv5aGWBRjIyepbaOwzEhUvcLmuRAApf8Xv+Ij5+x3Z8gPV
8eTGfI4X/NXTx/GKMJATWlo2uHBpMoUJF8tRXl6rBwq4WB7O52N1r1OxRuoYY+Bb3DrCKrp+UqhW
0mnlgY5NU+6zX6nMrOH6jEsAOXSE2TxKePeT4B3Qj5v4Ny8WyxSPJfQ3gL7v/pjy4nMYsuJOsUUu
NN0vqRcJ6TS6mH1JrEmnfcABbp1KUwMQZmmS86kwdn4ZoeTfGAznTKSB4Gh4XJsEUmXWeqiE4YGh
6gmVhTdkNSeN9P4DHmI8l9+0bU55dO+StguKfb6k6wNfYX0uyzRm4/aJ55LXfKaAZD1yVLDCQIsH
VAccUCgBYr45Di++QwFEVolIANgsltTEVI2VVFCVwyDXOJ8t8B2oIOxy0JgWlVeYUktg01GY9xSZ
BUcx9e+aBKCeOXHIh2ohJDu60nd6TgDTBRi+iliGvYXJmPDZdin6YKgSwrBrzIyNUc+TY8DdP216
tfNpGWeVSFSoDxnGnErnBcnZZYldzu9QtuTIkhVgVRUGS1BfQJvgF/Y43G0p3Gw5mWQNE5/xbq4t
isGS2IZ8CyWgEsyTeNJCf1jgWr78STB3/bxAADn6G3FeucmGdSPvdOfyWoko+mCI10/BIj5xL696
xJOZHSj8vCnlHkFBvRag5zy8YI8KD7445N2QhAqCTVPgHBD4cMWtv4G8Ho7zPCHWGxxw5qMm3fnF
elEFJSjSbRwJhpZkgcHz7SllTid8OWcqUiSaRtQlOEYS/E+w/8iEBKoRyRDrRN/KQuV00FVffg7I
y8ZNPh/56/ZooREujl9oDkVsl1OS4Xrs/4xR+zVQaVyn974yAL2fQ4GsRs08N35Neh/O73Utu7nt
LuT7UmUpGz9UU1OKx4KQbkes/jWpyO08MpFjEywnqJ7EqES4pzTYvAeHzi5WyVPRNBKwdbGVQtWt
bqytwUR107U3YgRDy05GQkCWJJKkuSefQp9ESNZbghEKoxhHBJbqFjEfydg41LEwnw+Z+O0Nj/wd
uX5vm1XbL9rA2eE8FjMQdP9zDlJ1vB2QhzN/Pq2RMfsXwlCTYrjpdzgeiBdulK2UKUFFC/mKzTUK
Dk9iinXDHmWV4NRe1bV7XNDBZRY24nq/SrfXmzZ9UzCxk9fhOd1rE3MMC6m7gEaTEZ7a50aOkCxq
myxm0mGdE6f+8s22KVVHS7ge60sRZiCTe/TyjNqKezSfeDRmSa47jMIzai7iTxFGmaIxq4WaEo/C
MzT87iEoSt4zb8WlF+keybGGsJS7dy/DeCCZA5aEcOjBeih9G29P3xY2JVBMgSEHvRrbSmOoeAh1
tU0wsV50+RIBovjKWdeB+v4plGGlGdVCRitKLMSupNuN475aoLI0xq0v0VYqojfFnn0ZZyORRfeI
Z9EQWkdHrBiH1spF0idRORLb54ACaJYfVl9VTDjz+QsmwWk4nQER1M1xEj9zETG+Weg9ar/+55j3
CjZiZNKDzvc4l890hVG+bnOnEMGBHBQCS99s+xkPTdR3WHCd4vMkPPkU1K2b4u380TxNhG/QuFrz
43tjWOn3zAzdqLcKn3VqcBRmlrf5rBPh3sO3pomuWvOGgNeMYPkW7JOXbsyeHTv9I6JKMYrkmj4h
QFzXlXkC+NzuuvDvZtQwebX3oiFmSMGp4FqIBZTbtp3gq6386/jItvKMnrTaqTDcxLpqXjincf8E
2DSg9E3ssS0iAv1ILmCo03MUwkDnqgSH5Vx2NFEpCBi46WyzYF5Te2AQIhl1urmRAdKmJ9g+fxkw
4t6JwE3VQXstpHyWkErca706rzLnwJBONEZqiKLBD4riWC1WEAjsZYI98n+/i6BxleQcJXT7u28E
555gZ7mL2y1WDishbnIXANeeK7uXZT5GA53T3c1ounqR1hULgLK446VGPBHQeZRpSXQa1aNkaIuH
uXgrD4v7bK0WcWh2ilZOOzMcQ7cBeNtdl6zSUF9m7MnhOi+N14hiUy+yQPUFs7XwqbrqldPXIQWK
xXEEIOeo40vXpBnbFjaVkxzO0G3juqF8pq4SulsJOgskqav8XjFuygT6gpjtj53QfdxcitGTMkKu
LqDbebSL+kzHVCxQDUZraN2nv96r/6ZMM8x/Rp1ZJaXm+BFLe/aLj/IzXqkKt+njRWOVd5Yoa9+3
7z/NrSCkLL9Hvn0jtdDZyqk8hf5LT7/2OUOM0lSrWnRcMvekUZJWGdQTBo27WTpVv6HpChO9DPVb
nGtDPS2GbX+nXLFOMd62c4PSRTFqwLqXJlwuylmYy1vE7TgLdzihLBSoBnqSUUXOnh23frjCqvlb
Q9b7w4K9oeWjgwTAvZSJ7TnhmGbKYAa6vNySBXgQA38Ug6+31/aBiq2sO9STcB6AL+S/jyhFm0G5
yRAd5ZFuplMb9xX9KMmCtwPbR0ZJOT7eY6rwrA9yery9jCmr/o0hoYRDQ0jTyhdwui8E9ACKN4Iz
iqvyQGYaDhs9GNEPOP+HECGaGBRZSqc5XlkGsY8ikiX3ewF3yv72ItN4XMMUlBRJTuelbf/GKqAu
W6FJJuLTGn/q6ceMYGsQY+Q7ZW/+0X4H9oqPPArF3RY3KjNSOO+vUyBhpJTMrB4sYmvcQwZ3cZHU
XhI8rnaVNifq0cuY26EXDnSdJbhrWJsvU8IO7UfwqLPP6fCyDabXd7LkgAGSbsmC/b9mc2DR2Sb/
FFJWI8I0p9k3wKLoUJ4R9CX/HHTMn/7hTyvJrk0iVxSq4cjfDkN+5C6RUSJWhk2uPZM/wR6CzPgJ
MsM9I2L4AK4wr0BV/4fLJzM9M29Myb7JnJnnUUJa9cg4XvXa+UDdIJDv/geHQn/jrUR4nw0QlotS
sBLYNRQ9Svg9ZVyKRh7GT/pRgjc6R7H3W+55+PjlzNoHuPGGpNNNOHXTEoZEMJhDqdmCTGvEzAMX
k0kjdbou6n2+BSesUI9F3aRSW7TZ5xpfLXDzSHVm9lFvRolGPY8cXZXz9t6aN3f1rEy4H5Lxhuzo
KSiHAGt0+1J7HW9ic0oNG3J6P1Tpwn128CljVmyzbz/fagzK9zMupDQCtFjbuW0Y+p2nEAGcZ3d7
wcH9qqtage9SAJ9gXm0m/6Une3uP1YZMZAcVK2OI+w+o8UWb2vt5h0ABo3e3TCD26NZ5NGvjentI
CgNu8qIz8qAckysnwrGmJks8eDxIpZHnW4A5UrtlyI921UEoXhZ/mtTc3DU0hWCqKKEjyNPnsRBw
8d+dbJ9xN6yVtHvvNXDH6yoGScpYZzSzw5W28BeK/610OuJomsyLckxY/9wVlXPzeCptZH+MPrV3
NhPzxGxLo/pUaTdi/PX5nhOr4lDklL9kUIZPyn5XEv6KgMO2j40NGJ0Y0A+fvr/LDDW/8D41cvTK
bdBehjPtArZhyB9D1VEUj7qazVxDX9EYgbKhUCqyMYrZYpJsY/jciGpGH4cmw8EzfTv3k/ol8RIS
GCBAi/LWBCerTI+GBYyKdUXPfctvW4/B8T9ZOwOHHH4sFBMsHLfSNSZMpEsH77UxUCFAHN+Jo7vV
thrAJZyNa/340980aIKhuYs/rc+7t2kqeLQDyyf6R3T3ys0LA7MZVtTFm+Ost1f03yPGOhx2ogQk
dyg75rwCuI3LzalXKR6Mo6mMDd3vS+NAO9YfFoLLaPixsUadk5zphF5q/wYli4dHRWhHICH5NC/f
o3ZJckhJ+k7c/C06i9DBCQQkp6Pl1p1gJV9n2LL1E+0jZsSQyD5lU28FC+HBO1cURcD94aqZWA4X
VdyU4UuCeIKc+WfSHy3LKITo7qOOvHLU3pIFhIZxywqFqZ0861RN3w/V6J/CPggiJGE3VNsx4S8v
NOZEKoyuyjEKSnJTmIP26M0IbmOvwhhrworrhi2jwNlPs5UmFSaxLT4+QDY3RBc6Tn8KfigoEjly
noG4XSTVV5SRaW6r6cMWtspv5zEsWT06evRdfRHZAntUOCJJyXyBvjiCEFpGZnFakSH5NoJdU+Jb
zFZtjzUE3pu0pzvEoaNFNcvJPuLk9SVvPmN1MZvDdkZMsr8z28cPAaFJMy6EzKzvMO6KOOoFXxRt
TzyIUePdbaKMW21b/yy9zEzx9o6sRQLmkTt+fVlmYksIB9nfmVJmRsG7bFWE2m9Mpg1txijqZqcX
loePCMO+/bfeUjHpSzvbp3glWgG/dFph6csrn+1T10/G4+J9jqqhU7Qns27g4WrIvKOBevn2z3CW
+kFE4tk5jOWMYumGNa5dKNIu3h2W0x50fZP85OV3ab+3Jmi+jI2DmrZ//lUa3icYZ9EPsKcUMhZn
RyTTSpBFGYAVFNRnzi/LtfaEf3IXhT4YI0ehklvXbYv/qgZn+ipgR/nSuUvNgrxsSC5m9Cs4/mZH
/8ebyr/6XwPh7jA4kCG0fFSAOzNK8nE3ZxOXlIqe0XPREvZl6IqRU/h6Bt4G6sbvGa1mm82n0qLj
7Y0TU++CN9mMNVI4fh9Po2vtJ47ofhD4Zsz8n4ryarvLx5pRV7o4BPDVI+E/MZOOg3JHazauJupR
gQu8IETzgNXAOPZmm6+h8IgTG2FWNWo3HbTk15SYOCHAqfaNJon7SbxrLDls5AaQ5ciRA8MRvUkG
4LugHtXs+gJ6863g7vRPvOJ8vXP+AK0EGIIT/wdBOdUiL7zY8hLnde08kBDhj+v7k4bmn8AuGUDt
Hm1TMLhRnYw0oLUQMAOE6fTl0sNyIpFbrOkVcQLr3VC07qa2q+QJCwjB5i2SLq81B9r1JwYkx4Bg
RUdzKGZXXJtRXgBsvTPr45GLPWY/iTtkz71V/xLYe0FSsgMyvQ9u2/uqqhzUqcSv1FREXNTHJEI0
s2Y3itGLZ16mn+ISQzG5qXF8cAhdPC0gfpI7Z14+HXSm2sgjy2oCNGfYvbAB5e9l9jW1LNdKLYjW
7leJcJA+hxai8W4Eh/1dTaQI9HHyDqsQaT9u15eRbLeAXyYj4IR2HMpCSw3qAl0txrjdomkLWKZJ
Tys6fNF1S0cbUuI8UcLLrwmPLdBvGIb2YD51T6AZKEGWXkRoLH97WA5jR2AdU6kKUcwW9W1YRVy8
pil69VkNvC/lgIpzhXMNzCg0+Qh81XpB304lmLGnUitEYpKSgMVE3GKjnzQFfdCrVGpWR5AaEj1k
q28ZSWa1XGTPo8RKgg4K3S1q5WHk0i5edkIPUJice8vrfqStT/7cQmT3IJ9qvYglDYveyF2wvZ9A
OnuAyPd6fXoPjPLlhyl4sRoF1hkDgZYaPJcGbryGI49dZQoL0C0uUrue6U5nRODxrTg9jNeWi10A
KnJsuTQKauAk/qsGQ8MMP8ZBQcvEKXs9/gjO/uM16670sPc37k82TguCE97SLru0FMALMm5k1kl2
AnvVxyWH9NU1d7xKn5Wu2SHRgWLaGdG9kezfHQinflEFE1Drpwus/tUGrKh4KqUltdjnziys9KIw
t4lUo28ehlwQj8HUpTwaj4VOHwTdIss7FUu1wN0DBUg/O1TAXccY3nAJy7gl+gkA22fors6lW2WK
IeOGfwDP6DwsQFfTePR8Mg1tpH3VCdRx9QjMsPDjPOR6YHbaEYO9KgOiOVBo80DkL6GQuerbu0BL
FrkNYICTubq/LbfYGDpLeteLj0TflipehW3yZMBgUbv4YcqOtb/kE6Q4K0+1N6dC8xb9tVxd312z
pyigHh14fw3s+OnrE9PGDk4bF7WgkRuKBTBimdsFyTs2E3yIvUuM/v8SLXivsg/UYVf75Y3918RC
/U4TEu2Tp02NVGNGWyYTTuSjVbFa+s+quVITH9ufg7paC0+5TZyAtuMfBDELctsKLP1VERcKsL1l
nyWhQE3yaCBraemR7Yr6ILBLXSipqVKYFMGSTilfbWt5b0TJzx5gkRjnbvryjYWnxKGj5MiKb3Dy
Jmy/s5QhI3SnGZChjkPQEW0nD2w8fIGDM7jpBM4J3hgiFu/E8KFR28XjZ1TzdBHme5OJRm2PmZeU
BdmBGplg308t6CdF25ewzF4smcmu+O6MShVaBfEHgFnqMIO1Diy/DLj/V/dfMGolsEdwyrtTtjow
+v3GquJeSD3bsvpUiKYOQT+XwKmudig7ylBtZON7+vT31RxFWJ1SD8X1d6poAlHMYxtGjr84Wduw
VNNf1oz7ipgDE/7w58oCn3hslkHcx4/SbfubKaTW6rrQItPH+bazIRsRrt4k+cmhHJ/vMU1wrT9J
nPOKLpwbm8tsowyo/yqYsPvxYVRliwMjj9uUz5PHTTGxEa0cyMtzDqSLA4qFYVMWyhq9DPTU3L0o
ZQCNEtcYUyYO5alzBmPW/ZUwVd9GhoVI239CT7wdHg9A33q3EQ0qoSiW3NDnXsqmifDAoCF4l95M
kPlO1qJ3prpmq1ENzEe3XFSMr7Nnc2hHfXbqC7Lg+IKCrkaQUyEbS6ol1GSZCMdLb23adPKfH7qT
Xa0urWSYbqIOrYcEAYKrbIiwThrnLwHtrvvQz1MY8vVxRE67769ozEJ0jPwRCrejYKX/EAp9y3gR
iNw6+7/2RKexuoaXy+7G6XI7POHp006jEWaTrVeYVY/HQdLfOyQR8H2QUl41ZrDZzAfAPOampzlL
und4O4il7GUlqbhbWqm9Sp3ZtcYRcc2Dsh8NMLeZqdKRK49hmlMRaRYk25mNSqGdV/CoALG9WkkA
svMC7SR3Snj/4hDeRERUL5qI5WANJBWJWWr55alU9/R66MGC2Kw+C5T/z37mCbXSJdsxEpjCfPdv
eE7Vrd1/oxJtJ7Lv66YaHlqGKwZ2z822OD7XJd3F9e6/AK2UhknQMWX8uQIjXSa5Gvo8iecavhZp
2v5xXAD4y9CaJ6NJQT2pk8bvHmyPKzNlyH0HU3WcUREfq4NXJfPFQEnLLGl83JexgKSoDq2H75vL
YDGwptjAaILnicYtPb3THva8aK8tab6Lm5cPtd/ieoJl4ghtvlW7jwNR3AB9Lx9x9VsOxAY2qmrx
UpiP/mLplvn4pQBeDA2oJgwx3Y3MNvXM2hm6D8x5QAF7qNjscdwmW8ibVwq5CHqaZEbnlRCB89PB
62V9jDath0QF1TqseUTf2kcUOuZ5clu7XjrzGPPXG0yfuAYLRB1YToDsdsnyjh+a5XS58vmTpfrc
kg76FqL9+mlrW50zbdFGZ15LgvPG9x7cikyCpXX7K+26yqG0uagq/e+cNEHAyZL+5scgzCzBCBaF
hzSWnoLCItlV9L/XX9j+fk8fDhkZJtpAc/4txpNnzdUNOh9wQnp83wU+llU0UssPo6qiNHiIFXT0
RkASKN8SU/Ya2MktINfrIGQOFgAY6e3+S9UcXVKfHab62oXDGio4qeq4HL3ufdNfAZ8IpCIqPFId
jiMRWJGUFrqodI7VbIYySGYwGCBMjCx5zHyyXFIWDew9bjQAFrwCRIYyrW/xrA2UK0yf4Qhvf1PP
trWNmryGYlRl05PjGLiKcf+sQo6d+eujkZW6s0xZRgX3KMhOUIW2PpUVbKXoBPaRgCW3XAbod/KM
5DZ+zhIBJ2eeSiy0XQlvOAI4JyVj7UJLA8znzh0d22eXF/f3XglmQxozWrhxDhKHPFwAzeEwfmfn
0mu4bgFDuhbD8y0kBsB/NBWwEF9ZYsmgSDcI1U6F0DeLcKuFC3hlejE3V9QG2aNQa5iwD/PB3d8v
5IrxGgD5wM4MAYiVfUEsleILrDWy3XcOeILoEZC90m5NpfUsNAoTEcZw0GlzlMNMt9tTPkeV1+sR
HsU+F0uDFKSFHkibretXZd4R9TBSDezwczk3zfTu9Ogb8ib8rQopBRHupA9t1IMXOS/Wxmmf5534
GXy1EJausBT3erqJPPU8225DwCRsFvYoI444jQqeGHm2GZyiWflNtyV3SVtM0zKJAgfP85pP0W4A
FEF7SxLuXlUjdUO7CSO6wPMMmbRGu2YZcAaJDcs98CgKlNK+BI+BETRBgxGylrd30k/GyzBVbiXy
kI7VMVOaiGW/na77sbQqRgCQ68eT6ohT0lWE5UMfvW3qQZNrEPGnhceri6ypd7Dw4eHBbk71khAP
tg9hKvzdfyUwj15xIt9/lp3h0goQJlI84DEefpblEFK8TwbZoYAAbiajFpJ75IaMpIXTCnrp7k6M
bZjDyvGkhpyTspNVCUMKGqJdgR5asth7X0nzJIChuAmxM7wFztvEK7SkMe7KxLuL8nmtILllC6lP
ecKnGqS1npoRwSswgsNb+9h1baLLeBON4Mmp5rd9MtgZPzKEmR6zAFcctojHWsJ3fJS71YjavMwG
CU/ReC/Kh/lTpvBwbgAi0tqctcnTz0dO3f52tChwsxyXDTvuM51RNVtEhboJdFQ9C6sCxr6XuM02
7qZKUmUVnIDQAgU6QAK+dHcelAR1/DJqaoyGZIABdnteVhe3dNBsjmqgCUV6yhfV/YyEkUQ4sM9u
AMcqbGRKqtD/HVLUb4tvQmYd7AZi5fL0gJZWpKLb5BuKv9oAlyr/vZUSLQIDG5uKnYfXL5CU9/hh
7ccCv/Qiv5k+fNwdDF2kKKmPTATO14AYy48pJJO0+gP0pMPVikK2cAL0ioiidg7nWLzloYOx0sWt
swTbu+avx2O/ddomWunnZN8X0WMQxyH/NwzJXMNTC4qBZtd2fGuD5KFFesiNeGWcnoJZAR600yt4
Y8drvDdmXRaiEpurZ2HqhEaFhj/vfXc3SvY5Q+jw5N/0eY931WpH7I8/6meKNaukVHxuieZjwPL1
zy8XjBLs2LAuanWguD89fVm4fgEu5+eT7Ux14zIyMIOPpze/vKb7s8gjhI0H1qmGcRabzlOLvw5s
7mayULfqpeqzbNR3hRxxIbDV9AsV6B0eYuxsFtaHX2SynuMqVnfpp4NWMhEnbEWECkvewPnZUXVe
zMjyHtN2I/RrKznUF8xOBhWHcFYzAc6SKGpfEA/Nu06S4Se0qy8Wr3PDnRX5aFqVuMPwEWrHCOJH
H1fYBJQoVSRKtzerFjBZlIVY1KUvX6H+yMX+PUTqmpTYzpjtgPCVnL+6ahi5fWSh1F/W780O2Tjc
+G5zbM2mYt0Jl5OBZc26/hSRqahXGKApN+v3ZiKa8XK/NrLOGOAB09mvmJmdjduUzKr2QLhJSx+N
I2MlKK0ziWE/EDHTX/nVV4+GGF5zVJvCqgEE7KzIP/ukFkyfZ25I9myvZX5L7QIsXsbjdTohRxcf
vp6nzTqWEregWOOs8To+KNOTQt+URrFOy4Qc3X7dujwWKmZ04IAuCrC3K1D9upgFMiNqPjCJWL95
6dWtwd0uCht6qlNoujqDA/yQym6CUIwz8Hm/2YJjz0dYN66euyeo7R9H0SLEtkjHYEnak+J9mi0J
vr0wCMQZ6JSSGKfHAsIXReyZ0EMOx1w/epAtSYxi99i2iTfh8WfifmS2Z5ifEZfFiFkCJUJfhe81
gIUu6+lMPXHcLzvUoi/iPvrUo1Einsk0j9m2ExK1vIf4/izg8oOhUZlsWffS9BM7fjCrpD8oLAdU
TbhXrkTPlYkE7Erzp47ngqHbkUuwKkQJKYXfsCY2msOjACAJv0DPU80KgvFB8zqZ6bnFdUYZYKND
k0BnyXtzqS4msmdg19+ouBv1TuJgCi9fx9GgCAW0LLWeHofl27h2743q/TePPfG0zpOGEzr9SxvX
G0A92Sdw4GNAGjcn8gD3qpSsmWB7RPXSbbwv/EV0xKK93P2KPelO7/OkODzd4VGThrqWzhOPY/Wn
zbYNAfkUgaP6hAxtah4kZRZEKkviWTTMrchp/9t1RiUvROEL5RBvQNyjkpyAbMz1Kqk+4MK93w18
+9PBbuiw6KljNuJWeFcwB8nYOvtGijHcmlTQ6+IyPd61kKS7Akoxt4OMfqtkyxHGiD+NfSQ21H8u
0TN7sLGjBQvLPv4ccu39K9/wKTBGBsM3X4vDdtS/wFbJz5ornq9vftb1Kh+dVGu7HYWn3CQbrbaP
nxMZktubFmtKyZ8E5OqWulRB0FSfi3TYk74nL9snU1nyHGu2nAq7hGsnZpyzrDWsbHQwtd9uPgHF
iUtNaGXC7ij6UqJ/lGaOLwIR9XhKAe2mCqpVoCvA8XWMbGeEN4Uv1fcEhNM/3PwWY3DY8+GanI+0
ckn3nN1JGx9w6bA60lj1LHCm9jx9LhRk
`protect end_protected

