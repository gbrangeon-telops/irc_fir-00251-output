

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
lHZAv/MVAAt3F19GG6CyO2D9ozHTHXUyHUqVqPhHJ9Up8V3v4BMtL2rZCdPHvvrLl9m3lxdPLeMd
yZjuwpNKug==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
V11pDh2GdTX922gInHRdE4PGQC5LocLJP7s9hbeXjPbTiX/dPLHGusbEN2B0toY0K8U4vuWNSniM
1aH2SNR2JV5BnhJYTc5D8l2e07TnA0V6ktY1z+NOBfbsIHPai5FO4rlYQdX0gfNxjRiE4WpTGufJ
+8B9yaPmasK5qJ0hmyc=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
0akrUk3wQb4EqzKkib7F59nSOOeoy+q3qc0fQDYykXO49Ll/FgY0ewL69TWySlFx1Cac/+BCy6vf
iumuPLpTjOS55mFm1JTMxYzM9NsagXEQHLi1lEkcr65/dw7cjFH/RPICXrv18S5beJM408VyZvsr
NCAeZ9gbVAaeGzkHq6VNPIh/P5GGGWEK3241GOn4p1v1t2GkteaDbOSjGK7wX7a4kTfRzrAH+xYH
86BcPdOp3oyEseFdQgL0BZboHxt4zJr0bXL7Ln+oOm7kGCKk4PXPdudDDSsXKQUPtDHqr2MHJwZk
LDVjKe6pX7e2DnCF/lojAxyhWqtc4aJmRRvYWw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
P2FMFi4MUNbCcmQEmOw8kkGKpCf5liEfyrVflbrNDPfCQyQhrfO1z3elwJF/eYuRk4Q8ng49IhJM
QbJUTOajY+rTGsCSJpmNj13e1oNpCtCwEA2TBzHdzEyAxDwQ0hUh3ZqnFSNQ0MMnavo9wEIKRylK
MAHL5TjDsmLJG1Zi4ZQ=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
GFuz3jjDcNus13vZfabnTsKTQz9Q9tOYpUUTv0v99miJHiWg9X4Bm37tDSsBPgge2ZWYV/fIZNhM
o9RFowO2ZPIK8CdMOp5y1r9QlxbgxiEVYj1tH56LRgvbv2A1ghGFDDY3Qvyz5G2dmEuSZ/58uAtK
A8Mm1zy2Ln16qChURWHrjkDuCcIOuGQ1GysEn2sqg3E/XWxojTbAmy+LaQrAOqIwoDTGFZ/Ek5fe
49U6fyDbugt8sjMOq32EEkOAQwWmc5uVOZWv3KIDCD6tRxPMIg8J9cwcCTEoanlasaaRs9KqN5go
7g24OWiCSjQz8Pf4KXR9USnCWt9Xh2mPsrZAPg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 20576)
`protect data_block
7EaIDnenVwpPzXaOgVt5FAxijIe2We3jr2MtQIUdZ8uc19Of8N24eSBaA06AGU0wFEZe0MLXSLOA
FWzVwKudI2dafiAP7CTJV5n72fPSewApCsuM9uENVw5WCjMorXxgcMaQsQ4oBxq6UIS5iQ3AuljU
r2ZwNVZDnF5rLRjfIfI062j+um4HCk57T7Q2PZfv8JMzoyzP0OYtXSX1RsiDpKzRcoxTWOrFGRu0
rn3MOsWoRZVLgRLcneEMGbiRVOyqK1WvK9+raFpMzdHJDPyBAlrk/D9ZFkCdL9DSS7a9XWqvnaMQ
/50KMqMHCh5XfL12zOF8osXQbfBD7li3bWne05VCoOLtaVKUSGFWMPt2zUoD5GBVDcjtxPh8MBEq
Zy+uCYhvevX26dqYm3iA5NImbvqk5EllQTtw/EQN6MiPjQRgnm/7kmOaNVfAqNjE93oANx7AIGC9
OHLDkG6tjBh8AM36DNuc1u7oR/cLpUb0zh51uNeD9PpV1lNZHN3QXUj+D7K1iWBZQSB8FSMl3nnC
pviX4k3b2SlyIEBIP5CaNxX8F1xSxpVflScJ5Z27/oH10EIl484BCpejWGX5WH6gqzi8scNc4lFu
ChkKKGoxoysf2obZwI1vH94xCxCSPp+jFTW1Rfr+lUNQKmM+V8kpKY47cB0tAt/0o2Uxcn1RKjPx
JqcMd26ZmwBagx1DzQzsZV7jo9NnBbZOLqO52eKpdNn28pEkMhLHMiUMBPniNfN74ke+3NSUpdb6
5lDxfaOtuf2WyR5o6nAUbQckCIngxKRw6DkzEQzubAUj3qNN1nE9g2/zRbdaZCfKuet7U+X7dsY1
J7Z72CKLhiueEllrlo5u0ehC9XByjsbeQyLxJrtDHyEH9ru2tpOgWp2KuATJIm9dTfLhyAHQdEVA
Hmeu9oUBxl61vbhSeeSu8lCvLYhiKl1cNXPf+2OawH/ESWF0tQyJbVoPfF69ZRuyfdcnbY8tkx1G
4l3sB4lPLvkYFoXW4wM6Skemub4+L1x2RVzpYnQZGCJggTOrRQjZpkMt4P99WWVf+bFB6D0bSasK
LTey+OkqtxCBEbj0tNgqpMUzPpNmGimNZLNlHmYMAoom8m1nKk4d/Qd3Mcgmv/w5EI+LKwJqUbBw
o4L7b9yPpt8fhJRsHr0Bdz8v7NRkabd8toLoqpj2H6JsnLPtjHsU3UUCm7v1roUelQ8fnMrEXY01
9VQlTqKUEkP01FKIb5ifkIxmXNY19nvyAg7Z6tFLtfa6MgmkwrpdeMBJhFYWx/psUSOw2SHvZ+nO
b3zhYbpMsx0qHRXphWs2hGj1xKwQQw647N2Nn1VdkNdItuc6vdu0/nE/oHEW0iS6ZHTZ1f2MW8Fs
Qg8aoDrN5So46cQ3KpuRfbmkkQOfxabmmTfW2+NTG12b+Qy/bwY1I2XYAzBg0HawmZUzQZ26HeU7
hgJ5RCR/rIY8YRm2dFgH5DP74tFtnwG0QwW64CTD+4V+1iXwVMiqeS5g0IoAtEtrLtc6n6b1frGE
r8Ilv7vWXCS9KSqzIrbrVp3SKDrFeA386ZYOjLNCxl7EId6uOrru537slhVtNHnrtuAqnbDO7bxE
9W4KIWU03vCy626X7VYnMIGpcNVYYJyMfh5ghRaQdH++0efjknJszgxBAwQi2lpC2fA8qCtqCygs
fLmO6d/W5zrchK55ywPZTYNs+RF8GDKtzNcsswPYiyEnZ3B0IO9tUETm/KtRRDr5PfFCuM1Ddfbp
KvYnRw4Grh+dF9eM9xhJvl3wfQNuqGfKYdlM74CtqUIZUdgQSLluIo5gQQ4OSa0qYLkYMNJXXkxB
I/guYKxpoQQsZKCEPqEaGY/UMBJy5dPIsTMLYFZAPNrTn5zprPChKYtGGVS7EEP4Y16kUXS3gf9v
/8lYiFGzEi1nc0gFhO/YsJjDW5loXSc2/P8/znWakG4ZTvdSW3XtMgt76YHBkidBfGgOztvRf6si
NFvqYI3vYgrLUNAMO++fXEYXf0JD5SRhCt2g+I2yfr4LohOHkrlLNOuF5/P5Ce0DF1IQtSI5x9NK
9k4Uuy7UeibtCrkmo5CA2XZW90fE+B+Ug6nrM/+datCGFF9SR9CK/6xrhrLF75oOd9gx0EHt78qD
PGJHtmQyUp5214O+yX4cZOvxYQWSpN2Zcaff6uBrQsQmEIQtHiiSFWGEndo3bUQJpT5MbH/LPMjS
ihmIUJ3nuyxl5hZgf83rvR1kOYRglzeLbaLawuhOf6cjVqyqeu+4qFEhUhIxwvkcxB+Q7lKj3QNu
EhrmPx0wv4ipyTI1EiaoWotkGk+LM04wiwfh6PNUitj7mjcmywGQVuG4x9Ip/Aexf3uj5aEG373R
S3Utl08IiC25ybw50ILXiQNyEm0w0QFjU2ejzJX7KSdqBTYGI18xNwAa9LRxuXDUvfa5SqiFi575
UrlvSsE7KY3pV0/GYrkNtkw3/cP1uAGnT/Gx5yAjLIeZiK63IQGnBNlr6TjrOwZLNQ8+amRQyCdQ
IjY9sBfw8cwzO380G/JUSVet5Fd4kk4kjBYpOu33BXKMZGB5EDVkLGPWQMOTg7DRvN/gBoaSHPS+
JNJRQwklm1kwXfLLsTcuoqQEpUWKTBfMiGMzdLNstVil/CTAuRQ7AKd8tXexpIgOaQL+FC/AgEmD
06TIBuk1QTuKRhtIEYun0A/asAsPwWFWHc3Nqcr10dMjpWrDFPilhJWlTQuTBSyOAr1vlqflQyEn
WxL+awz8P2byiUIyJJdOy2FtsHwxP0+3Zx4cLMCefKkzdm+we0XnLRNfxiSJ8LCUwn9l+4dj9feH
fksR3kjaZj9MQ4tiNqIgyBohMG+ithh3282sBHbsFi5YuYK1uzSGiNhQF98wMsIOYJH/6cC6IfFH
/XtVWfnf5Zz7P0RqQdD0L9uNrxAtE1FybAgQ3VpJmRebJDoF9V/DIG5pY7HJvzjtP93/bzJroUTW
tGdqNeAJKNltPlJXewZubx2qBYLgXXnbDrHkWeXttTLr5fyzPowWiuYm4hh7UmBI9r3J7ObKIu0P
yyh2+nTQ/SR0slQQLrZwTfuy+4TZMvqEJfjjbfiE2xyGRHHg+TQy205ar3EV69QuCx5bNrNCHQA8
eZR8DLCmG+kjWrLYTmrZY94f0Nh3cbZBfJhgvhNMPHJnlsFUGSqyXqsWmY4RBL0TiJ55YX4cAcW9
DaW3N1q5Vm+9b00mgHp+qcvX/Ut2If/dtUDDx/yUIgOZQy13N0oF/W4ezDvzfAqM0fVj0J7goLlb
2+d1bQ9kXfCS/zkLt6orAr+MyjID3elINLYF51QX+BF3JBOsO+sVdCx7HvMII9yQxrgIsr8KHKsH
YPunb5nT+1xgX1Rzt+KIRqe+E7+mJEpvVskG5T7AYchbXfVApcbwdUvNQ3r4CzReyRWgyia4gC0L
hKqDrs/MJElZPLO8UKkmQ23+Tpnvqg7jOEtkhGYN2cyy93dnOHff+gvqf2mAzdSpamoLCkVsqkkE
p+/qIvCrz1ZoQenYo9FB0zGLHfa3tkvKLw/sdSeK/3ttTaSiQUQ51tDQBc3DrxaKuS2oFCcj+5Vp
b8QWJF9Eot6uuv9QzRWUCeAFhTpqIZI7350yi1ETgLAQI2BaTssFF9jpIKrNan1AvqhY3+2bZP7h
eiVOxXAV8vFc8qdPtK0sQf7+E3ovMMT0gNOrqNFPk+FjvwwSE9SPxbKA3poYpCH49LyaRsnfm9Ru
2mLjfqo39ZrVyfB8IUspyhr7onQ6UccismXhDj5KRMteLD32d5z70rTWaaKouHBXKgdDEWP5p2Ru
CvxHynUK9HpDc1TLTrPNQlBrwJKtiYkD78tz0AvCiev8bC7hoe3RB+wpVgHAw2QapUjEOwDF7mXS
fac6rVokEXNuUXBKnVkGvxPlHfN6HYkSG2hPFIWogPcknoImpBQT3ovHDCsnRnai9BueMRB9PmBw
PtWjLzbHQoaNH24E0HuDr92HtEYqjwwn/kXjPooeQelKxRD/valxbmxmUScN6O8ONre+i8to4s1A
Cv0YifRzFAs+eXY/7zY/FJkCdnGqAA3UIewGzQXR0TY1IB7Kx1TYQJGFhjHCgM/1utWeSXa6GJzJ
FzxK6A8LrCJR6lKY5L2tKB2lCmCQK004mHtmQ0oWvE6pWD4zz5IKzPACf4tOmEiyfyumooXQ/QMp
UB/CrBtXIl4cMO2J0vbLWP7JDg2xDey0sIkl5c6PWgMOCuyYygfMxDOpdGC2CRdcRC35Hdl5TjPy
skUs6/ZcEH4BI2U022zTYFyeSlsRp09XlAMTZesy0XW9AvA7jko6wNX91KCVXT7sh3xnDXNkFOST
dE04b+IYfUpg0dF05J//o5xsS842geRcSe66CXKr89qMzblJ/WcbxDLUHHxDRXvIBqqJw02Av7Xc
qQnQ7KsbLB+rcRLhGiwiF6l/nJ1XSM3ZcDV9jibZY7asyt6eeyfhNghZSZMCe/LEGhTfeOkNbtK3
l3+Ljzl7hP5+iRdejJz1GGaC4ew9jBjDrhEVt0d3JUXruZby1GZAIOsqN2Zpo/PXBe9D0628ws/7
wbcojBOxMR5SADUbIWF/YhCJS9kO40LtiTrwtY7dznYdCHKe0iKX5wSvuMPMgacaxbz8rxUL89/S
k4cFw7HTJbwzsJdPY/qtRxFJE1AEH/wb8wHH7dr2r9a4d9afFudisFj1Ce7NVZEmAtUVP+Pgx/V4
yeEkOdvmhraSiXDC+FxT/1kOFEb80YwUFHsHDtFiqHTDppgaitMqOjOu06jiJVwVf8ovux00aFl9
qybA/Ka27eVsiHGciI4QASU3Cl8oUf+LRc+tMwFvZ12lmuxOHHKIsge90sqbRc8vlGRQQ3Y99amP
fdFPBwr7n0fW3W4epEygLFKTjLxYstUMA77BdtqBWfnOQb37AlRWfmXWL3zv//jMgMSJgGbl/HsG
ni86knOqdD3HeejdGuxRGKFhB9UicrJcWxygav1Cs51FsX6NduGD8nF2Eebgb4/TexZXxcp2N9Et
Jk3h1rYCLuTGlb75G4WPSQyY7obWPpPQxYpVAnTJM9Nw0Kr7i3dFqWJU+XBFcTWFFQwAMFC1Hjf5
i6kua8QijPJCvON/63gl8ngl0pvSRE3iYitvP5J2v4quZtSOvpMKyQmuaeCmyndeJSP1rUSGVqhf
LAmBr7qe1jul459REKaTYPmKTnKLUN65adHRfNs9/IzrHxky1VbfAjziepKTBgk44GRbDgrqMLr0
MxQUckVxO1NZeSLDF5ST7VjByardTDAF9HcwXg5dyH5a8rG4LhYfkqoVfICmz87IZ/AGXrGJ+KEd
ZDEasrfonWyMM0BTn4Pb3FDDnmllOV9uwqUJAPAWRpkuo2aKblwLFkbU+UnZQ1fw6whrPeESNNG0
inzafcN0CkzugeiiGUrJmxnDXWmeP5QmO9x57YgHj+TFVdT3bzhWj/+qNA3MVTM1oeFH0P1THb0g
eilOTuuKL33ZbDQeHVUqY0wUHGAlLwpySiRcj3lmWLkQAgr7uG/YD8OafzoiTKgs2hMv6RzBrvVr
4LUdxbdn+fQX/R9A/WnVDV9RtWkkFbIe0MIZow4ZEJg/8Pf1ayq5ec2r3KXkJZiQ9FwN1/tvkm3b
BsAK8aGArFL/G7Bo6YHMksLFMu0qR8rHdRAuV8aUcIz70brk8CuNDgkRih7G3IzQbdsyIWb2cICA
TZl/lpkV789rbisvHz8sMf7j8miS1T+S32JfSsZpymRttbn8Na7hU7gkXiHHMmmqpv/HWDlkcr9v
ma3Ep7PJ4Yt2/l0aPqn6oWX3GnyiyTA6T5ljkauevga86sUOv4oSikmBHk9lawynVBAh61OBHXQJ
OUuKtoc/zdfOvx8sI4MaC3axZ5xz/69bFJ3KQ/z+vxMpREKIbRlHMVXIZU0QrudJuRntc0AWyM14
Kxxeu1kfOLrdtmGpu2bS8bnQRtL26nMdr5f0MFTxdjxXD51rxfpQOlDLEJYoq1XOJiR/VBTA4L0f
uaXsJMnI79hHzFME95OYNHlsoZpYbmw2Q3Gx1iB+WoYfQJ44ezYbTf6KpoBvcED4E8QzPbV5FpQx
IWk0p0tMNMLoUBZ+HMF5qizOgloVU18ilsPOpfhV2XKRK6fV93wlYfWt96Tyi5NmgZFbS35x7N0J
KBTjf968uqEaqYxqptSsms7dZXWmBSCdPwxw796j9mpwDjPE+i1DXY+VzDsMAYyLBwwGorhF3G95
GOBWPo3lDdqZOyD7XeZXnWVt6OB6NCQ5xcW2IPUQYVIgKXQMdnWxbKMZe6yX+4G7F2o9AthyuTlq
fyk2nki7dS+u6eB13SFrY7dkK8beEdeEY6VC3sTevV4JmCtIxeO9k4dK2o9QwcLJiI/DEv6u9Tdp
gJP+SX9g2qHHKiXJdm2ychHNFNmfD/wxz/pbH5bBvozij4UUyeDALvASspmyFPkY9h/ubupY/OCQ
0SRV6raB1zQetgcN6N7ujTg9G9LMNgAi5JxQ1AwU2CiepzEtiCkmA05bqLDQGpHCrcadQeSDZcog
NWVtXuLgWGxBDacESWXC9CCxzkgqMoHphuRVm4/L0vPTEY0kP0UjXfkElNUBVGbkcQ/O7qRBxcXw
cPBA6J7gHrUAplujQBw6SjWlg6Xa7oz2r2IMGr9nWDMvEWqExRo/T0JzX0PYFI/1MTQksmrqHS3m
C561OFSzSbj3LcbBnS4c/00s8WdkX+Nv3xxopui6VHrAOiHnfSqWgcUk6IQ3hrjwwAZx1nz0ekFa
vv67Z7uQJzHTOSiHZM07DlwaEWti9AQu2pPtns6MTTYKemw8rXnolLWAvClsiA7/CWQLUmp5JRck
UISlGUWpnGKEQThdoKffw6VgPSIX9v2gils2F9Z4dvMR2+uKtEnQwlYbnJH9EkAGC+o+ptnYInCB
o38P2Bsfoej5Bh/UA1zbpqrhV0Ptfh6zPT+Ef353JMovbPptJEOPMICoq6XAZDtQMEXRb/Dgqr6t
lZupORekcy54WC19c1YC0fmw+11M6dlCcovoqp7lwl1EMIPLs3KMEJjWCJlk30j5jdJ+lzzyEIJp
74IXaySYYxsMp1jhRiEKMOIOJfSMsUoGCHbOsOMoBLB6eK2JgAv0EV3a8JtwNVLy5CfbgWrjm+xo
k0giFoxJJHKSaOtCiQFmryqJ4P2IuxHB3zas0tWTZH5+hqD/iHtYD+yOPGs6L95tXxiSoFMoSu/T
XW39dFqTI3dAxyV3z+uu0OGl4kTc8+5x//zvxZ+oJHTy9M08EqDQXThQqW91DDTrY8x/XLCc+wIa
bB/VaG+Zx3NiHwe2USSHioclGBA76hHM+A8mm46y1QEHQIPTSeHnHCTl27M/bEmdHtAQy0YCRFwJ
/NftqWNQ+gjXV/fwl7cU50FXWCQKOHq9D3rIokRt3FsNReBYgW5oFSn4tQ/n1ZzxD/sttNV2sx96
NFaZHJAywUn/v+WYyHd52+D35f+nNTxFISGE4/hnW4V3dr86aJHBau5GaEmlkQdss/tBbLEBHNnk
As5hE6ge5QCdDB2+jO2COfI8Mn6OAxQCXEZLlMg6JaG+5PJy5Qgmh0o0C3vyxlfir2TtFBsL8Ny9
Gn9fPS6Ol8UmVpE4JDCn0skhkjSgXC3s4ylBDoSZDKM9zhCXerz5Emft1oDoOkBvdSViP4Let6tx
YbeysXmVCAjjjLRVMvlTs/cXFPBVMp/IapJS6z700RT0sSC46enGqYUgIX7zB/3nHIv9ToigdTk/
WIVwVj0mup7uEiaroMrXOu69hnj7X9novcPqYsAxf88vqej3QpiSl3aWAa9KJSIQFr2nnfTNu/DD
VNfUnzC01+fvs0PSyp4qookhl6mrcDHIL6XcQYvwnis6qTwuN8YNqgFqdvZ3vW0B8I7WzfsQKRa/
gSiPqyuqshGEBKPoOEZi7oimsJtRshCS0PxOQTSxt5+U5r+hfcdypN2IYKcfHniXj83aQnumLBUp
GyhCc32IEO+ixUwDkE1mEQJq/GVMxW1ySRJSw6kUUhdA+jCC4gHNm/Z0QvbwXNgCsK4PYEJ7T/Pz
xlEZnxHcXkL1hJqZwPrZ1Q3ml4kgSwrtqTrePTbDnvvryaEmRBp27p8PglK0gTum7cqGYAmfSVAX
PTqvnF02Yc2AAxPR+MW1/AGv0hhA7IVmExC/ZiBwkVUkQrFDdvMThfKf3aAcXWjby9tgxlRVbmaS
ImC/u3hvr6GFiAmjhQESRRM3AUnM9JDKk1FN36JvFXnm2saYUSTBzcsA+pPo4ggym9qfdofKXkvS
JN/uxZuwH5y4LmJqkSNFEgazBVi/GUq5zMXM9Y32dL9FWWSh978OcURk30J0lP38QaD7ZoVOVw9f
emzy/5OtNbmidTDfaHXXDzpY1//wlsUmEaDNcqGqnyIxvzd7SxTUIF/+ff8Btgx183bdJD9EebId
zR2fjsGjKFYlpQxGnVF3xW1SdI3MgVlXhEF5VLPsSOpKbauwZ+ezxXh5Xgum2CMpyQfUU0XzRgZg
JEeh9dOhDo7DK5LjXTrENmVe1KIdVdC82p12uShyS2QgOWN9ScFFg2AySpb9pTLK6VdAJ/r//n2X
YPN09z2n+/tpSOcMNXcj3xBGXA4plnO7k0DYf1crgzhLUFuIX3wAy/G2L/CfxD8XBsifanq2ddoW
/iEvnaKXWYykhi4flhhnWiH22hPGTDv/6LC3wC7AsMREIYtAQMosNTND4R+gf5nuglO+HzQGc0nv
ECI0IWwYIVSSSRfUvDpIanOa58pwogynPHIXLuZ+kfPuTCZ6qLUQilfhAngNck6ksAP6sVO9TB6o
d4qeUZ7nn5/iViiMVWD4muE3W1YZDFKjcA75EK8cHccIbRQbj/bC99omk8iWZ8SkSW5QPHWeku1T
ijhfhpCnS8rFnTpcERpjVYgu3oLoBCPOWQWSAwgG8q7bn7xDpqTr95dYzAaNJ9ahMqqJsjWm9aKm
XC4176231d2PTH9XLnMOw0r/MJp0qEtDVtpS4b0IUQMBuQqvdCIh7Dcbgm/8UV8VF1fZoyi2m28Q
jICc3+SfTnQJFOZ0VF3SpnEP4j9SwCMKvDHbMCUl02lIxPsZU3RSW1V5D7K0CN5NxoFQMcMDw/Ls
TQM5ZClz6w7R+zJopYgl9FOWGNi5NCIJbT4c3vT9tX4RTElLGTxeylxH9Q9l6su9BLsa3e5CKQkc
QS1r+/QCMwHEpAwUGV0waHXL3QfohWn8jF1Jj2cPMKrhJPkFou6RUd5zo2SR5msKIemHn70WYNyJ
v8xKVpnBH2gUKNbfvhFy90CbumReDT/0JW4W/ka8lDsD+2enC6StbNvPm/2bgXyjCK2GkyOy6+OI
Urx4QOzVBMTYQ5XPS4y+vW/yCcgMo4AGq3KhbHEt+KH+6F1M4ce66CzrFNjQ+B16PkKDqrnhmWb/
XvDXbfQ7sWu2qlIl4/SKym/47OIvkF2sizduXZQDjuuKDNQh3L2vKj1LuMNZo4g1plyG2yurqf/x
Q2xs2IuSQFwdQSnXomWZ5JAeZvsY7cwEDo5dsa0qnwnTLpzRIugUfm2jF0xotARxJLNUtuyiRacu
+qIjoRrsW13e/kATRAFiOA2y0SL0JxABsMcgHDWA1ul3XFzZx5YloPTB7WeOc9sqRUJaIUmLSeSA
jfkiRzSvoYQnTo6v5F7ENupA/yGQNDGwrHue5BYfraab8GtWOOtb3eGtrHZsm3mYcXeqYRqCDTzL
frVPwJMTS6a8GmOd+HZ4UxIpEPT28j/toMqRr2s39R2fxHzrVeAwwRVmzIH+wvBaHPPitk6PiGfy
hr7PjeYqNUP7HpvmsysvKWlDvEW6dPewkHNGX4FZ8E5ACcXxCPFUu3Jg3fgLkO5JYoC3M3382YhP
SDrPvRnZcxkrrl8O6RafuT9rg+oGuns91sqpkZzitvb8H1FeLAuko17TQv+xFpaDdyLCxLYI5Qho
8FjdtMl5CZUXgNZ7b/qgYB5o5X3f25i3VnYZCmz6LsaI+r4NL1CumSPS6vT9SUGxVu0MiS+SJDZX
ni99cC93Feaj3HA/k02/Gwh0FnM7u9L6/VtdrUdGteZGI+3pZsYkLTVz/5hdoMwhU0S+lJJe8abi
2Z9YAmRMjYBtXcPWPFQ2WAD6VbYLuNYnAnLcBIyTSEF2qxFr4bZkfHinVHgkOdYzm1pFS1lowDdf
7DefZVL1fZN3PtPkUZnj1rqEnTudXKtP59DSVc+VonySuoV2D87EaKdfBW19gI/Ld17mBFPs/leM
K1/xtzLSrqGZab9ORSD3pC7S1HaIjtG0hU2ZUyAW19coUqTofk2YZ6hlktr+QfK4sc9Ca/q+TJO+
0FhkeYKxDLtLxlKZbHBY6EgYr9ZoGayheewNhGTPQVmh0Jt3SJSC75ZWblBJCzqU8ep/jkh/scqE
HiFrG54SRQUDJOHQohg+0joERouEk5FGTKfyIv3XI7lOq44L1yJzfNkzG4JFVYlrWZyXmf0eQ+Ja
6UAyu7Yq5m7GvStLMYZ3Iv1QAjf00tgDepC332tmLWz6ORKrCpBMfPmFYcYXgq06nMtFCrRoOqbD
XY68DQPcW5/dIklFUXmemq/9iFQALr9OCDIvDW2hdzTsUqUoQYFlmLWx7ptFsYSZemPIJ6Z9Kgw/
EUZWSgIFG4vM0sB2CaPEhUlrIC1mOf0qS7KW7uN/fz6sSaIOX2DwRECCUO/Ik8PQzUnlMAPkXhb/
tpHTY20gSpz4owIxsLs3hPXOh8nibcOJODCkc9miBWFhMkBfreESbwPVYP1VyWafwcs1VGD/83WG
KPZJle9MNnKigZHVaq7cscV+6zoHXFNDKJjFx0/wqBAutW0HEt11lB6MKcAPShed7dJY7YT2hM5s
kdBLG7ibbkH9twqe4Nmxicky6bk9PF5UCumqlce+NG1W2zKMb91A5JrXZwplfpDR+06CoRJHOOT4
LiP7iWeoeCBAfvDTd6ZaNxvsqLLb4YK4uQs+q+XkOF7GUh7b0qe5L+jR7lCJ7mzpGdTINVNbnGP/
CjAtlfNFdWFjWSJbr/6ZBcS3jhkmEEWoL4Dj9hQPMM3gX2LytOi4bfBPqyhIeJ2NZ78Q+/gUs3Uq
YufvM68g13FomE7JYtYCNmUBSq2CBYrcUmcYA/8xtlHGl5lqV+1mxEvxC9BMNDsCyCMQvBcW8jpG
9EwlMrlSfcY7JIUPd7JtxBdu7SFWVBVCA8rQLNyXpdFgCW1yv2NmtQuL62C5fHojG3dhlggo+QRQ
tWxizWPcH7CZoDQVaL9UY/1YE5GWRvqYS1vFxxTD0xsE6UhtpuXaUZNyysaVFGu3jFfoEXrFIW+6
75Cd3F4N38pA2Slb/nW+GepxFyV7MtG9ToLxi8dfkEvwbgcFGL/f/ipz/TPSnuBKfdZxdxMkpM3i
IkRYKDwnGmz02CkHkfh7q0v13OMxPvXgUH7Rl1gG8lgnhKslKGx77+WGaEVASIdzG5PXkv3Kwjfm
sts1rOeBnD8lcTkbaXZf5ed4XM3s+J0GM3jJBJAB0xPXZFZkVUH9q0LXJ0QDiSFEwU8JZl9A94zz
PKCWuMJ6Hv1O30g/xyWIAoOaodYalL4viedwK8ASDe9YEaAOnTJvtSUTIo+a42SHiVdQyneL+O41
btix4x7NtgTWVSkm/bdwuTUc431FMAYx82jiOkCqoBGn/XPM13EizbkasAVcpW4d6O4Lj4pU/pvb
o/iiJw1z6SF7E8+5Y9qqh771qozqHFKemRB9VNDowgUTunJdYyaCiR7FxN9Po9W0GA7QHRHTtWqB
FR9nvGjni0WG5CK23QlFYcOf6kQGAuaDJ5Dw8GH/8xRLrOYHTmxMep+NLhCPe6W/xPxggaD8PBV4
p+NNO2GF3TIdGnaoq2C4CX8F8cTFeXWPitO37CnCd3Mc5rVofOuT+fqLHtpz+BX43HJyfjua4zwe
DzqLk2fPWSXM5FPMM7CXb+VKjnBXyjdXFvMyck+yqo3GXTsA6syQIYzw6VMhTAJFcAIonTuqqFg+
DssJTOY9maUCfv8HuT9r1KbinOhRXcmfg9iiKc5o6wCCZ4H0moKnozjF1R31YFuozFy711TPNisz
lxxPITFItNR1JcnqfBjPqtii6QeYmkiJTolXH8hfbJNJT1xQX6+YZmnvlBE0dmqTBURPwyBIgIK0
fgqZyunUV62kxxIitWWEJh/PR9021rA9YocOAktHYAVaqfLgfo7vV+1fNF4b+aCldAfCci5Nnqrn
4jh24fq1BaX68Aq2Ew4yfuv0fjFR1JmuZjmNKw8ShYcWp0c8wkw1k0up7JmqnEj75P0/tjaE7duf
jvliShzPDS3+joyga9tDTNXZEJtq9zoKC1UKOCH+/A0GwHat0sFc9bFW4l92Z1Tvt4Za68iQC/oV
ipxp40EHcmHZI713U4Z+psr/GfYOfEOVs/uQ80TXz4oUevMoSDs5s/KFjaBaFVCd2XwTdROIloR/
LA/ircvixEKB7Df5yruTBA+8Z5u0b1+RiJbqP8tBgHD6ZcfsQKUThXlt75G+uFIsDneGnaaWfmEC
OTV5Iq7bEuI2D97BbDv3mNY8vZfNo/KQzeB3TtGqHj8v0xL+oFYkIG0TcDxbueFXmT79+ZR9ToFx
Rf+jQC//llVdzoIsXySInsu2TRol6aJvao2Tmcg5mvMkQ+Q1oW1MKhJnuNH4SsF61wWKcWQZ9LvK
EV9CynDSg+EjERWfGxDGtMiNamk6IuI+rqeMrR5dAxhMWG+TXFbz4mD5lQKTqIV/YhfjoTabSQ8J
NeaO9E16yTbwopd/2Q71K81w26C+UfeNSzYuQR3bqW65iGNpRccNiP6kht7mW5K80GMryVOpMNsZ
ou87aou0JPPHEM39dQfdgEjgFEX6132b7jrc/cQixk18ZJ1xTUq/ZEzjU47jQRBDBlmbBpqdh40+
QXKw7W7FPIsK8ocQ2tr7LKhTI1araMXHMAsUhZ77eeXQ1LdkMXunk+R2CI59T2sf7We/bj6DL/MO
Psbl1v1sdvFN2GT/sHzSq/2njAV6a4hlRTC/8ByS+aj2QlCMaVWVyAdNa8hy3AYJI2iJubSIeKgi
GsEZJ9yTcAgttzs+EGvwl6undCsZo6AC9RXDN0YG1W0VR+7Fj4tnPYRbw15gVBKWKwqUOhK2kLP9
Mp6TDt+xkyofs6qQYkT/Z1AnwAK3A/Cz9IUafNuM+z0LvYRrpHxxcoSXzZqs0wBkMXKMSDmTlkFr
tiLsNNcAqVeEjRYUZWerwSk7cEiQZs0vUSJ0ottjKKb99Id5bZRU4/vnVnAxsTOCBc4z0tYWzY0R
8r3auR0AC3gEgbuJA1Ed3DomITECsCNeY9gT5zZV/Ehg/QckmjqLdwYzN9lk3oeGpXMbaGzhldmb
3lFcEI1c7LuZiD2ttNNSRVQkZKkmdwc9wP/ulyGghrneUGGOCXKaMRugFK+DAM74FnsHKsPmgffT
+xKPbVPjxw41inMX39bGGIWGysMkeqOaSh8DIzzI30vVOQsiazuXZ4vkzenYZ98qBIFfA13F+BIR
lTC020Vj0847onQsWyiOAEnne9+r5QqDot8mej9kzjahGLWeC/4IeowO2QeWPgXxBVM0fi556/wZ
DBNmH2Wt1X0Tn+ZGnwU3Sfg6wVkvmO7ocFz93E5f/bSzt9qIN32kA/FKWmRcq8da7AsJaaA3BOAP
oGx6NghaOMRu8ML3JckELTV7gxgmY1dySFAMqMYcsoPtsXEM7oX0jIhXfmRSc1AllDgxUkoBL1fw
LiQQFC4WfJXDzohb8BAWJirYMrpJxlcBimlCc+UpuI5fnBy038eYMS7U1m4TcL2VgBxCOTF9gDeg
5c471VDifRxGJ9pMQajkEA5+2WFI98HS3P8qTreCvlbzlcWda/72ppQlS4VMLHM1bdO+cB1UhZEy
NJj9Ert6rvs44qIMiIVimEoRGdNEyQlcF87X8NKt8mBYLjb70vvzs1JeVxfhQoQGvTjXWtBn8it2
KVAIKxVUvQCsptsPJJmMFwmS+ANGMllT6gZKyoCv6vZocgY0uUnZLctD47Y4vTmaoFbnzILtwUjZ
jFz3bAAUY9jmcYb2iRc27eA2tFMjtJlvU/3ShoMU9hushfozXE+Yhr2fuJQztCzDgwlbVBAamYA4
zlF4cLIVGnl3E36YE8xyRDIow2Kiey4XNW2aAV2IN7gVQ672t5pgE2mGr/Qtzx0QXoaKKfqjrJU1
7jrKXY4zfSs+LYopqPSclcOcc9+Ub4kyWncvT0pXiGgFZd6JklL7tRPDPFIS0hLAk1nznnddZCLg
p81O90NVKNQRf530/FDiFyBE4mVlp4VCfQ56KIzBRXff7UzTAblyz1K5IFBlWBU/OnGWFdEBaOd4
JF3jAFhMOZOmly/q1NdWHhzqRL0Qn7ahcXeHRbJMqw1Mrf043MyjuYndkaZA9HOOJ3jn2oPC2WcQ
21UbIdy26dCFlgfaSp/n7yxt856N3nj9EGi+2uFe1/e5M1DNfmkC0tdReENZFyd5VJAOC02HlMWh
3sUZj3325kCrExdmpJvusDlbmw9GlSOmIQEB5nM4sqYy4MUFpikL/EAMtxIRcCgu3p9r7rx5Zxlw
JtI2shfqhkNjui2k/Q8Tzl82lGfQuRyI8MeUvdp51kN4SVuK2qYQj2Ehf3u99/AfNVF2b8roi60N
4d0q+8DXInAmIc6PaN8tPow2rNoOH2G8YRqvRmw9JX2AmZ9EGPkbod3FlD3XODvWWlEeNUpCp+yx
j2vQaPxRDpffk4PIQB6owDjHOSLa8nKv78Z5P8pQsn/9p9p5V6kVTOEwkieUbToPqz5u24cEeCYB
cycQAwXuXWw3lR//iWtBxfGTivVA5FsacGcvOopcHPtl077a0DxFx0hbiL+rVYo8NNeNny1VwtBX
F3h9w618Fz78ErX4Ws7iJLsWoFgv3tVZ5ytwdWX5A323RaNMb0aVcaO2GsRy2Mk7mKXpdUsQryru
PxMDZ2jx0FPlJWDAUC2lPp11s4Fm7euFu7hStY2kRJO37QxtlN4Kzf7NL03cQzhFBIvR07fDmiQn
of1ef3CzLB70NevtFWKlUCToigYn+UEnUUPUsthuJoULoAuE57SW5oCZGNjG3odILm2mOxMzk7Zu
Am3n/IuLgy+E1/UHU+75StJKwx9wue/oW6ZYUYirQppVMhWe1w/WG4YPUip1UvWTIdps+HJfbH5o
84ahzH+oe32C7V92XdtY6IoF1XMSqup4oA+gNouhkuTlJG2al93TkVsxAjri970E5FkoOd7iORnr
3yhOag3lhsT/3pTX/MMNTeiiXKC2KlQIbtoDw0S34ESJcICcfsH8KxvqPcw/sCkd9ftE/rpXpHnf
dzeANGUSuaQwOwsl57RO3sqhlMj0PGyPnSEzRTN9B4kNRdMVw88bijxFdGpPNrf82Fl1fGGT29oo
DYIWbUnLwD09Hocfa0A4rgv6C5gnZ1fhsQT56Qw6xnZNAIItfXf/+HUJwE3pBxAARXyX8jwY8KtK
hGpLqZhm6xT48DtnfuBy7Dv95GS/5d3LfaW1hU/3l+w9wAd9QA8Y1J45GJeYpXSa+MVOfNyLGYeh
SsvDRzdghZvBaCMCX+k+cKIWs4uEYq5Yb38AS3H8llKaCaAU5LV2jLaML32Osho4ww/ASvQSq/Te
x1b3bO31030Q7IxyCo1JSq/rPQjFyLechgjEGuGOqY2m/KT6f00IuWnJk7gRfyMK2gZeO9zQ7g4L
5rKJZf3HRHSms2/NJUH2k/6zjiw88/ZG1+UTc8Cb/3KPXZNcEdDIvjGQ3ocVh3IfJglq5c5YeoVc
+Ujm6UE6S8e+LbI2qwEgh+BgxWr1lfH3jcFINFU0g3RixtYogO1JpwDgzd4jHeaOSGf8vsuNYAdk
PkzzgC+QIcX3xcqlGFbWt2Z3aKwAsK0+6l7lbRHi63xuwmsafk2+o/JBmOcu9bOJLFJ6OcvnW+K1
6HNIhPs+Ty7ItpUmB2x6qo/CkGCyAXtG2PdDPuCHGFw5y1levoooZf09wVbn7iqJzSqxU/Ipu39x
XTOJQq62RI30drK08wZn5a4pa1vUOEmuJ1XIw8CR2emiUxL1ZDF2R7WgBVF0OupM9rzHABvFzfCX
l5hq/kKzcfUgfZArRrGqUJQZ/nivyekDOw9VP9CNb4tlqCwedVQwaxwmEDx92Fb0PG9Qcy+TMLc4
aL8D0QImT6RtR2fxizOgqmLVK3HYsE/E/m754F1x6YJQxDj/p3ZOf416bQo6phlpLzRgDx/kusS4
/r1pAfc+G0jyosNKrxjVXZF571FXaFSdVHToaeJwNYiqIfpq2GRol7+NMymsnHFwic1wTKfyBsCe
p77YzCfIuqwslxC3Ot+DX1R0OizS3DxsSjpuyJVfPk5mcXuKr+iEdevQdAh1ZLlzCfnO2ijgbdst
xGjm7r0QI8kr8TimG+4VwBChlL5KCWqyxixjM1KzM737I9k2GyoCbwFD/UIle+hsawmS6+/0UBh+
U2Cs3BYgEXsmbq/2Rz+hhbqEpygMro102WMxfLSglHVM7QxgXwgvBsU7AAmUuRYF8w7fWLjrOspE
8tRHLGvnWe1xnd0g+mo0VSl0/jkiE0cygvye3u7z32mwynaYEd8hHA1+177hNDy8LomNmNLKfoxk
c2lwtNxTHuXeMFmkUm7SPAJoYF31sdZYOEuWMsIdtlGdp1P16mZTuXPNFNjKf6MYO+C7oieePJdz
of/JaNPEqdPQ9apFTXiy55+xSRqSWlx8o2NvPu05D79PEQGaor/pOm8WGParVHlSW7SPX+gzDQhp
dB4qm1AqiG/pJRLhUAsW5nIqaVw3yyW/ngIvQo+cYcKuoxYJeex/tMp1LxTjkMbwTd2kWgNndxfn
xKYq5ADmU+dEgP2OfKWhMOxXff+KudbVW3eGyVZQAAHE4mqK2k3YksuJMrswyxUX4MtNwMS+1LpT
JGfXvVhZiMRJCFg/ESAajdaQ4JmdyiXa8qDoX1cJz4ZXC165qDTm8XJoBYmvYu17JheMy+QKmYtx
Tr3faOXXr+I02NOH4SVx4HIDOhyYIGdKlYq9AnhG56ClmDSZ4AxB+qTPfDkbkHKxZPWUPb/XoHR0
NY+sfq2PwKcirwxdIXe1rIsi96QSlXZhVNRLPr9lUkY4l5zKUbkaFDCbQSun6nPu9dwrdyYa/slp
EJKYe3/R51vgJNIt9rnD1mjywmHdVB41qAPcOgeQezqkdXN9HnEjmHlZjyjUOXyMO6Mxjx4zdqho
TlggJro6Lo8daGqQEqo8zsXBlzXwtnZwcnk4MpxHPkxZzphw3oiFdDZKd2/cGxmYab0svwPb6p+N
HpSeCxl/ZRZUDmib/hPeuwG0AiLaLePXQWyccA7ojwj5+IZv/Ow3gz3Li4oYhm6QUDsb5ilDXIdV
b0gnXDhrNIujljcP+XRRfj+5YO66iPrfYWpiUATMdjEZYaVQsawoD/MPrJqLqNj3qKIBi4GyySYU
ObDBn3TMbEgbYfsawgGqgWnOjnsnphP3wE6i2i3zMMOVtJD0Q9MLBSU3OMRXr6ywrEs7jCodavjF
av0gSU3qd3JAzQeSCVysSsCqdDwqxQ+EsSWoykNo3qM7L+zCWj2af9Vx4mXD98qvIgBtiWgf7eCV
XSqjcy7Nx1HGHbZwNKSeyety7UOjeoUVsIimqHnmlzZoIj6GTfzRZGRMqwXHyQZVdufM0LkBhcwC
YMCRziaHfHekgaX0MlxFCJv63uxTHmLuCCFN6Kcm8vkslTrrrt4wGOjpkM1j2MEnQrvwRuJQjmT3
Wonl6vXLdLvk0IPhLLT5+PUKTXaBWIdhTEsCONIgw0ddLNR34TuawVHjBLPv46KRLPNCSqr9FK09
c4vcMa7wIE131Db6IcG27semy5BbaZb7UQLBYFpj+hGSLjB6GDDkt6l7quIiK8D9D8t+619+AwpR
F3/PWJuGFgrFntQ14iVG4Ei9BipgU2aPer2GLlwEYOtbA8w+oPAOWzQYvUT4ukG7axtYq12HPi8j
2GHjmNCK8A0xHRoOZo2U4csDytXWZi4hUQ2DMCoBih0gM+YLc/VxbwFEna4PZwYQ5XR6VbVuzUSD
162XtNJ8yK2Qnl0B/9pMFlrSpJEdkgI+Mj/D4VaK6I3oNJxtfEROb57/ZF2G6+7i2cpt5aaGUSnB
NoC/khOMeXc3WQGYFURgnDL2Ga5tsX73u9VXq+nI58QrIR+Iwq7QMNnG/Q4UTL2iBCylFgAiqIbV
hpYq8gyWPZq2mWIevijbg2AXucY15xjHAW4be9ZiL3y56LkbF7V7dkXKb5EDp/ELzZUFYU++CutI
wYXwxV+vs2xjL8pYUyt4iVTEwfh7Q6wrvy1Oao9cmFXR6TxrOnChuI51klMRO2ZH2tOX4zOqMfQJ
1FL35fCm5+6Bb54EVhzvGe6m0A9dtchdd207sNV7qIWDzLWTkfqELlVdQrsXgglXgu0nFVToa2f6
YDVOuZy/pOBhhTCi7J7KIFGO0fd6jpRe8KARDddmvQbjUa156cP0DFF/5/YL2FjfM+X3o6CCpvZS
b1xNi5K1RUHfR44KqiJj/uUnpWD9jLAGwrQMUBl+hEEPpG9Ac9fTM8y8wDHfZLjWxSYadMvPnuLm
1rEHhm+hZObM3+W0TD+4f9xUkC4Z+DFn7xgdvxD+j6nirO7audeF3CDdfwySHAFX8d0A8QnSbD09
I6sQ2dsCxqGlRDVnaoNWpI5J9XuaaiQhCt+4SZoQVNUf3qlBKtGMRe4oTHdQYaKkzH1vp49sqab4
IP0xNDAZzsUx/LauA9OWlftpVD4vtEqfCSGccCEq/SEPhjvocpexdit1bb/KH07bfd49Q+I+OaY4
MwlbjpZeasEnYt0gm8uOGO7V8PvnvkC23s72/PVj1HQbAsebcOl1JeWsg0nL5RlhoHRw28T8LHg9
wjbADzKmDn8SfeVbGH0kuL8FvxS/YWNoSA7CnGh6ZFqWKi5NYfPJvK+jubKctS7BEDkzWbBep7kV
xwYvBAtJ9Qlmy/Jv74dja2BF5Ke4wTNOXX+7FqP0FUeV75gmbPlYOURJwFbUFkAhaqo6UzmevGGV
G4JnRdNmn3l+yb1gYaxb3blCRmnbdtvffVVxq6nzEGs6phWts73NCVCTMCPARCkZ3i50fN/rELHE
qZRPrYmkyg1ztBo7DNOl+yNGXlxRq364FfjB5xnV8UOWgC//TN2iNw2aNyT0ZGDzHUdSvxlMUusc
sPIPEjORKgo2urLcYTOZa1+4FkTA7xM+NK5kLFfHRgRCGzVb+tffbB6FpC/LrceHTTtjCc3guFI/
SdRQb1bF/kQFjnUW544z2vkioxPOKOkIbRjKcH0Yr8zfahlkz6A3Ak2Hm9wNR7SMMhsiVg6etpp5
oiCDKVzyCH44ZF0/mkf5f5LkkLRE17q1FIo2VKVP1u84puHah/J3o+YjzW5QS/3n9mn0ZOQpYYGE
o9yzsaIArHPFZ/jM+0Ugnek4/1hiF4i60i3ygQFLiHMTdtsfzPt8sHOm6G82o0hdOo9fSh/g+Qqd
zq7adAmx8wvAX6XxyLyNiSVJCMQgkFQ1b76XTyEol6087bsKTTORh5mJEk+d8VjpurNmmH5OLmYp
vBIzG1Sr2rmYYkqsaXMiuVsePNjIDMJfHgfmf9jmR2kLTme9l8R8KyUnu0NtUYwzVFapVamVke5r
KiYiH5H5JcSZ1Prm+0OjbZ5X5BerxwV3mz42fJn9PTc77q4RSP6sKiJjByy5kcmB3w8tJfUqe7Wk
cIWPz55JdZHvLmv+8iqOGvNBoYg38/IIXzdgLAa7TaJ8QyTqzD7GpqRw8hs93SLuGRlPqqUcu4k0
YWw4WxKx1eIIFHGXM1eaYIBRhUWXXyAxFoAmy6ePxtlylzEsRgRJR/CG9bgMVz0dx+Jtw3d6i/sz
op7D2bmgxQPfaFmJMHb110kzDp3zk6Xm+igipVyOZD4l2esCZFCGUQqrFy1byE2bItsmAK4xtRoF
w/mL7MOw8HOFyeKmym24aaRaQpCawa813doQ8CYnm0BC59tDyWiLSgrp591+vFP9f6sX6IMUvMF3
MsdlmNdSWS0cJQlCrVCxXmtmglKi7obcyLJnvYYUBXibbJzVsh0c8TpvdvWWQed6RkSNuysfMUN+
M92NIcHHtBFh2+Pkw7kCOMs1BzV+ZvCsNxy52JgwNQorB2IxUgR6Kwv3tLon4tO/nDorHa+FtAbQ
fByv8LlZWF75Fyrdu4mHxwH8lm319rQcmyeRzmVXvZax57o6SOrvdHpi9pB9WZAuN/iWehtZiIWX
Cnllndl5oZimigHxFZifxxVpBlBSrjwSgEAOwMhyyYKOSU4uy+tJN8uhF8YHc/YNL1NMgFDBWF3m
fSgteAVIOsuZ23nfIOo+j09ymHG9nJ/TKLzopOhIN7PFhWa2icIHW6v+D0xEm9FafdI/A1YZc+gs
UiQtOY7mVPsAKEuh9fORGu77UXkh7CUKn7tx98OJQPNyEZwf9l0sNU6mqvw7k9z2xQK0gcQQphXU
Q9UsA072QV+QOrr5LONmZ2Dbkrp8Zi8jJsjEEaC1TvpMALjQglo26qdYk1+GnAkB/a5meKKuRBvD
PX0OeZRO9GHqAAM15ah2L6u+IAyPStjs/DBlV5JmACmkVfTrZDhiArws301DdVXY0Lk/+1UCdigz
TSfGXpHuXvxqagFWfJtR2rXmLSoAJ+gBoiwhZ83hGhKTkl5mSMM9eEqNicB+todqW7+L2iUWku7p
7e3wmJuVRneGDBh2v6TyliE7N3fmeiXPVsU6DFxKNeo23FwTtVtxgPikZZwj/u2Bb575Bv0pJ/9I
ZSLcGNTUBKK6srJxjMMEe39FUXg/pC9pQpYM64OKljpBj6OdlvLoj1r9p32NmruP3KYG/OFV5jeC
iIl2kPM/1a46AEbCsk1Ap/m75X0oCXVLQh8kg7kTd8iPX22zSD1vw3uW7xU5AypFCZb/+Kjskle7
QdXk6eayvyd7qnlq1iibW4st65fSAGN5DcDjvMOG7fiO8Kp9kGj5/cH/p2PuBMuIA0c/g+1DmKuc
67EKE4exhjAC2RrF4pT1lhrLAtNRwaEXsB2esjgbSs6Ab3rmGLYFqin4ar46NOoW49nQWJ+wio2Y
R9ZrDyT73ri/zJtbtJ0w/Fpvn509+HczCQIC8qEB095AiD3tz0repm2E/FwYa9qv9w1hyTv4Rowk
buoSfx64QohCKBz+3VQv7lrFz1KPu+KnhGSGuER92BjBgGwaWiG9qhehum3GJ2Xr6I+Iuy2ftNfZ
7HRPJuvI/tnov8WKz3LZLr7NPt4Z4/0SnIhCS9xL6qUAgvg142AKQEXCVCbTp22DtGU2yD0WQjnb
qM+yeuLNyzw4JjhSCV//0TZ9AiRirqRoHG1vMxmHt/y69g7SQOb9sEKzUfFx+hrSPUmB/JFu+CN5
N2AI4gcUYmqQom5wm+9nsJbrrHqJJ68orqkJsw+Myuy7kt0ebWR09CFl7MZST4xKknQcLP5WyH0a
p0mKDmBR1QBH+iOQspoHHw1NJE8AJAHVB96yAWbzj1/pIQwLwZjqXQIh9JRJIigUlUd+fHeqA184
NqCbbq0BAyHKqO4mmz0uknkyhvVrlcGkJZrCaw4oGQWew+OJDHY4oSaSMX4bEohvslnzNwJmyQ90
9yt26VIQnz5ZHHUfjx5nQ1FWuKar1cvXH6Xih45aMt5qQWxzspOTYVjwiFwkRboI0FJ592QOiPqg
yqUY+EXQuQ3ONayPJnuhF0cPkyIdp3fve+UvK318O3BjKrNFhI+t490yedrgcxKk3aTiLEAK7zUg
2D1ahsQhZVJzGO/XNBEgAKR2dlxshxanLKDj4nnTR9A7Hwqbmvbh3h7AhNCInCuxtjAHvZxUP9p/
UFh3le+xvyA7cNh9LoLMImc7E81687vB+FOeU0bUL4DGfXnO+h+87AD1n7L3SddWoYF6OTyWLzTQ
9o2RQB+c86mp/rA7N8vB7/biX34KtX0gJ5VodznTFHrldSnoacuvysmlKZa3Apd2XebhnjfNOv5B
yHW5QzfDyCyo0LJjmu42oKUo5dPq4Ed1qqyXImmnX6DUGYxWSnPbGfgrLm74d15NAW9lKutICufu
Pw1EcSRVoMCkEFZ6rVDZsfrjU7z+9Lf2IxF0mYw0JELUL+tFUcXlGZu8dqj9koLHWU+vjAOoyyP1
eKyUB9H6fHJP1E2jqLhVCT0eedbOzASXpIyJkqGtdWUduUzlGgPh1cRMEYkaD87749cVQin8kia3
BJjPlAuIxxUk2DMf0rCH0VrxPIOBG3Xe473HW3bTWdWyy9swSISFFTaZzi7uk/k5B3hM8EBVz+cl
AgiIYKvaICd6e9HD4a936jZqN6eaSSHYKXMvtN91tgsbzDGjUpUhOGBlM9RL5tCdp9x4mgyk7AEc
kJEuTjsVoU2ETMlh2ST0zVOF6M/iqdblTU+/OVrHXVqcP2GtbkE+b3aurD2OJxpevP/xcGJ8vMe0
uN3tn9O5YrmGtCcbBtaCQQDfkFMASBLsK+5GKWjJr1yWvHSMfFQlz0d6xejZViOvMgWUoUgDhqkU
Wy7oDCjnckJAENCl3DReaHoZ2ornIjPF7O/qOLkbPkilKn8EA4HVpzLZszeTKy0QypgdfPK0UJVR
2M5sDMVCCueXN1iG5GljOuaRD0RDoHv3oM1UB3u/XS746ofZRGXXCki7t1uk4/7qcXxKOjmS9MJZ
udTJ/8WPsNRznxSdGkCf4uu+Gxx9HlLz++mdwLqN4OvCctoTQ6PdfpAJvD1F3OaBkatUsKX5ZjfK
5EqHp+Thp1cW7h2d6uxwmaBB8UFD2bwp3NgqjjQpu46c7pP15N+2G2jlvJCoUGFS5D93qoz3wI6Y
fUQ4s2MrElKGunAYO/f9eSrwPnOr7xUgoC2zMyB0WFaSHAmJ5T+5bj8elP3ByxnNIe9c3SFV/2qO
2Ps9Pl4wiYFe5h8XwHTgLqo1iDoaPtvuItWUzHiyFe2jnkRpEIr7UXDILzDYuD3OxFPePaensKRr
3L3iNYGQKOgnZeM821fXfbby/tSmZFxlRr0b5RuTUDY7inhnwhnEH8uWf/vcUx3NThxNg9ck2V9k
s+u4HdbUfPQPRogfsMglSYZEWqYaTdE0mou3eO7zJuNpkYre91C/eUuHG4QzauYwlaBvb/+T3Vw0
+qk7FZcb8/7RIBd3ZDvMbPDPXdrOHOXN8/Nsz5ze0k8AXf/etm5FJDRpytykfiyJDUujeTn4pNH6
s0K0MsKXXoP/NFHpPhkAsrnEd/zk81pyJQ+mlPnX9puJrYz+qkc54928Dbq02hgcqG+9AVZgew8W
m+f01KbIDE/68GeNraRCYCZotLaDyPcCGIFhemfHeYPUVIZRBI/ioEyEt4GXeDws4PI+wg2qcPVx
mNnLyn8osGx00/KQfOHSZn523tNW4AJJqTWloZpFAW1XYmx8N9CnhgmAdRsLKsSNtUDzq1d0Dnr+
nQ504qzvlGZZqll/K99QxI+qvCViMXhthdGKehbksnokW3BlRmTMUMM8xCDAneIWmMqEkVWU67wy
uecbhiBBIAUYGOzDAxei25gXsgq58s4Gu5wbbnn3KUFRIu1XT6jOyMnCTLZXcVAcV91b/utFfuQT
VFQOQWDOHrCvjcoaYncsZyYxDAZ03YAvZdoet876mGlobqbYjhBICqClbhpdn6jEdwlUtOZM+nte
s89id8f3ZKED3pNCWbHt/8jrbYwWjmMrOx2zLdxtgTLk8XN++lhiuePl726ysiy991GfnD/BprlS
cmelmWVFuIL278JHX/E2w3nSabn777sSFJMfCsTVYOKJ0pux+YSfDq3htGUjIZreqD8qOVJAKwJx
CjaGtz5rQU6hFjKzinsExXS1t3GFtpk3n5KrLwvAUPvogkKOf5XRJlBvV6sizcoIPNEXk5cROEys
npMNxebPhwkP8Tj4dT67BIzdepOLtKXIUr0feTjfMVZEbMsCnrAqVpDFMDOzbViDqg0VRzyjnvxX
TUzmsTlkbleR7OoNkBq1JOSaQj7VOPJxQd0BoYWAC4Lrp+tk+CzG3lq7V9IVjSD0UUSBQSR0LM9G
gA+a0H5tjNTfDv9AhUPRts9Tl1iauaLNHPLxTPljw9xYEWZB2+gKXSks/ruHZ9OjgkVgV577aOnu
4YttwrPxUJrgZ7qwqqcfysoceMce913J6vRcYNpFpWUcbz5S/E82n9HHpoZqcR0k0anZQds/7z5t
59kl1pz02DKgIEeZPEHRNyHtnPYheoXp/qcIlf8E6qXH4iVKSyTlv/gcjrgXa+//PtSqlXFQqw61
sCsbwmvMr+FNuDh4fgJ3vtMR4XJIbcauj1TYTHkCYbt7hWw2d+C6BbaWMWXgyuI9wFWBCVntpccZ
65xy58jJXMvVowpStkQbNZvpcKUkr1RDQ38SEEvQfDkkgoynVCcPZpR3rW5NycjJdhjNdij/wDU9
cKlRwL/2gcoGd9qcASaVC5+OWRiDQBWfU4/TowzVqSHkKVBgrXyIoFRlurKqJMPTH9R/8/xyRuVL
pIgK6/vt3b7Z3fTxiXFD5CNaeuMxO2bO04iQBQEcX5uk05nBCcpGxW4pUlOkhdUGRtH1oevvfzDm
flduthgU4CoQhm5XreesdCtDjcUfwsrzBO53pCLGqmOcIJmrg7DSfS6QmaV/rIDoaabc5Y/3Q9Xg
Ayom60JHscmnHFuNQD6vQ1RiTQxAd/E6ervNZ5QJFe721tG+F8FZKbQFaGc74LVOv1JRM72RkRAO
/w7sdhN9Fad4cqFrCLSF5OOufm5Nz45C9SqgWx2i8x+2c82DMi9ixjAzkmOQvOuJg/O40JHcE/Fj
GIcQhW//tmwKuQ8h/dZeFd6jBSAL2zkf6QkQg91IdlQjsA62h9F4Cxz8BXycpTuJ9LzW4SwBnC1D
6sZl49KvR7WEfqiumgOu687Slk0y8IPZtiGjPR7gknUOgc1datH1RdIsQumJPFYr1/Qby+OV4lmT
BHFJ4TUbmGLq9qH9aSQepZqSfjQy7BsHf7WvGoDiTJFh0fJrlu81iKKpYbLLPFo3So0uot4B+9Z4
2f6vdWUnlyTVb+2izySPYODOOKf0gYuiJZIAEf2RYKJzIbKux/k5vxeWHK8aPlYHEzqhEfxBX+D+
70TEwV3zpZUoTHDVo53JefRMOhyOMs8klIsZXii/tFW9tmzOcSitM3Hu12E78+kqrblMct+0gtyA
DTQmSsOXUBQJSkpt6Se0IDjxBVvJSGCTxaA1rUVgAYm0hCQiAyFKGz8LOcqLYJNqs/k8Du+vJIaA
vUndFySbWyQkCFAlIK2jHGmyI76WKQ4su/enZ5YIAwKIlEjUn5hdazNhdX0NkSPgR/ir6oDIeULm
HdKwLTId9HELEFrCs5Kf1bEMsJOWmjoUaz0dLJybu1RGs/ZMToaClnhaCGG1W7V4sj9XaHu4IpS+
senDB4gTbsVAJdAMm1d3OHYqGEqqw+f47//LQpMUAPX0kIQdwkJkwpwqBmJ+pnsTodHjTnETK3y6
HSaQfJ9sH2FtIawGSOzww4M1tDudvKt8Nfq/hyquBjy2hHXRUF+cNhXeawHiJWdJZM65Mmgb7A0k
vQtFHeztSa6EW9m/GEDW4JBxjeiCgV2zPuqELj/05FVRKmgNrAuoMGoDZ9MOZN/KVwcpnbArwyRm
Ah0Yrn48a3Igt0V+hHdlii78eb/x8/LXbnwBrC5domVNZEqR6ab/ja4oPbbRsC4D53VSfEMWLh21
NNsp/rA+L+4aqRwaL0ibmnFtzgy6f7pdmPTmPtgoD469momB/87ABlI4rxH4m8ZSDh4FbttkP6Ag
1ozsn2RKxCQDaUrVzR1+AuqrSYtwW10OIpyKHNjxI0t+fFiu95nWOS6+gh8hZ7yLEozohQf9QO65
zbvcncwZhG/TL0m/gt9o0ye9IcpPtQ3io+LDIneeMgb1VUFGCvMiCRgY+/t33JT+oV8ann5isww+
DqWuZH9Xb2hiw0UDXJyc1r/paCSXHSlggaIfSWhcZfhnGX2pL31haLLY6ANBU090ioeUGvZwai0f
GFcoCCKY7wS+qjqvdcwupBJ/aiXlmqOO5GnWyNWR4vdV3uBhKnUbjEHEzzBA1pUYMwYyKuVW1zal
GEzDbqT9EGjzmVKZFhLwz++/kt8v4kv9165siV6bPBQnDQdQF+y8XQE6OBL7nqcuo3yUOhUdvUPM
6yctbIVbBQ1i6ly1tHqAI/2s3bREAdIuv3LweaHqIePQAM4nIJ1irKAnkTM6Nr1ZLnWcTabgALZm
9Mcjh4vtIMFeJfirKtfXDWqg6XLgN+4iF+nf370l2L7CY+Ltfhz28z1fNZkh1mptsYJz20IoqLJ2
7XMuTEpAMAgHtzjws48i731h7uxtCN3qfJAIpOPdiarWCHTWJAM5PWQSxu6rxd3kfy9yuegFc099
sP94S3V65tcs7Kool/KsQEzbnugq/v4sdOfemCs8iOHBXnltBPFX5sd6DnM6hhQqw6y8mGYJkzvg
T0AvfRCggxS3jbtPDPMIH8cTJMb+Z+Vu7CLlsViJ67faSw/5qGAfs2jK2SFw8fAX8prFWlFOmNRN
bjn6KOvPO1xPQQ/oREz6pbIlHxHtnjToDCIIengBJN/Dh8B3zTx3LOvXoxE7cFLnJSHMbg4k58aL
uQ82y5yB5zGpF8a6ITHuvJ90P/JCxZXoRm7zHMHvNk28cVpRrAEU2/tpsF9b+ubj9261SJIotQwD
fYV1tTYaekbqrRFkxSI4Wx0J+bgIaj3TnT3T+jvglft+oil3JpCo8F0Df5Q6E4d88f5EkbEjWx6C
Y/gazjrqXn/OcuBHsWAcuefCTTjg6VHEMEscXrsP6VAoPDZG3VsPzUrG4AnQRVkLdlGAMjaqeu1i
En3t+3kSK9Ww75hG7vfWiw1yyix5Q6Lvt/ez0JMGZN/SppkVjkp7NrB16Hl1N6vifmNWDEelvkVU
mVjje6A4fBEv/MzYllPM/H9Szir4cxJrweqtXGqUYY1OPFu5Gj8a0ULMwPvwEj3YdXTXVZrGGVLF
g2Q1YmqFVyJzmxlTdV3YYkEW/gP5vfIqqqGDlp7ioLRZz4799OSUlFu+mlG0AE3krF48SZ+eWLN1
HHVuzQ8Bv8UuYtVsLQG03QuMH66OzjlR9T/EaYzxqUxaH/MvTeGKXPsEzmbF5WnFhYZzaj3WQJaj
/SySBbHGEb+LH5ah5JCQTwGqmKYIfgLBTbItWUHo8kETO7ZE4bLMMnrgnI1vXzO/OMpBB41hsS15
j13q1DEBVX7CgzPxuUBhP0iEVVmdCxMwJB7qEphXjCch0tfw/ztk0L5JuJBEo5tmxmRRz7gy/Gxc
oIhOdF8aGvEG/Uu/BQs929aq5Aj131xE6jl+q3O+OmCDwWMCVXGmwNhcGaMQ/e/nBIG1li3ipTM=
`protect end_protected

