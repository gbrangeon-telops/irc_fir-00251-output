

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
JoMCOWeb5WJCBfHoFXpAeueDDgvCDiGp3AckCc481MQYfkwqbKzf91lDJ35VGRkR+lnFDdba8hVh
ebdPAvk8sQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
bZP6jV/nU5x88OLSeX17wUzGVM/1H7fFl1OvjJVlfPM0WRyEzOpDDBDAUuNgnxFvzLOKKYEuQdGX
W9Azus4jUwU+zlgsaiCb1S5W3YMjUJKtbRQ/PvNNulBlTlfZaMHLAox9gfCqP4OK4hzymuRCwSK9
PA7SK6I+FbKAacX9y/g=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
38Ya3DupjVbpSJ4i6CmxC3OEuL9qNwdAvGt4GnhSmvDhP9C+krqPc261IqfCwYzwzxzaeMibTDWx
/h5fHzYF2I5fsXilkoEoRxiVUecJo1YSbQfTJW8OEBtN5aYD4EfWNZxg7GXemsfNXYAT3IQ9OGaZ
Z3OnlMzYiNTbG4DNtpaaHWOF6C1ZcpZaMxg6JA0ZIcSPls5SVALLcDt5FUbDAqBNYpV4JoWo+qsc
FnhESB/fKp4TYpfMu8ZebNdGwLZE/v7NBBWsur4E5vgpE96o2V2PrhB/yUkeOaYd/sqFfOVAPPYH
mOxmomWznEckwZ7yWdfaca/+EES9Dh2xe5bnww==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
D5raxCdsBjNBeucgp+JNk0QydQuZbfT0hk9FPoXi6WfKMKGXanrHw+M0M2EvNOZMUencxzfv6CtL
nCmVqYCrBCTP3KURzHM5DqNYzQyp0kj6XGMA+Q1QHtCCtnTEsuFMkRdychCBXeOcnfn0sPqhPAb+
dDkLPxvSvOkSf8WjYwI=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
KE84+0MQOal9OYCn+WiAXywM19zQ4xYNV40iodnIlowR+vSp+kbADs/ClNTsY+01AbPMnO8ZTgZN
CGRjsRjKcpFcdHcCbRqcEDPJE7OK/v9PEqPDH9NFgGw1pSJUkP9IpUNC9/uKTepjTRYkaMQQIcwb
MA905J1RyQ1JTo8+T7ZjypavwIpWqfh9+/OtTNQBqe8xPN3IUu4u+7M4P7P5w0QOtT0XGFUOVu4C
5WyMVCFrGwdZoGJ0XcMR+keGC+lH3zgKGf7XDuZwC5nPj50Jr/CWT4G590JXwyjmGrh+LuEInmJ7
dRdHoyo/UrKvxi9s4oal4X1UmgumWAW7Jj7wfA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5824)
`protect data_block
SCcgaOjTh7G77hRCf6HOotiQFoKh3hRDNFz58CRebe6WUrFQ3cPEFdS+FfUukJ70OP/miAMzPsas
lbbzNa2Apboleq5RXuqIygmZ6pTNf+jctJ0HG9Tj1o6dDFk7YpwmEjFJEiJD5AFLSSmJX+gO6vL3
gWaTZwV2PxfQsKfR+zibj+dFifAkPYAslt6FfJXlOcQG0bKVxE18tjSevuvy7khs/d9rkC9L1cH5
CqpTPiLAIbBatitUpduFhjagIHYHLSSjqyUyGvM9Kr8YvmYJYfLUiM8+HwNh8Tjr1ADEwgnWcmXe
0XhDs7gvQI4dAEXRFveq1YvSljn8V8gUV+iLvZfz5uD0nE+r3ezLI4SKAYSoJtWMNt09pxOjZWr4
YYMmeAFgf+AbvFSUIExOLmLcg7Kabbqu70cj4CHKzvD4wn/qF6FwfHk88W6Y7sVbhTJWj82iRxVw
SZtAIniyQm1YbZsBX2HODPAebkW/u5aRPKzgHwBuFdmrZSsVc+REWzMbfcD8fU/r3nrKIdKm+Hq8
bODQvJ43CKh/s9nIg8XVBTYTYZOF04Fm26IVBvkgjdc7V2FJug56QWvX45ASvvBVxrNdnSFaUfFe
cSApZRPoru4RKvCO0hQwFcJcivdjzOovGDJOerI56sip9aIIBEoIoWa5euJyXRUj+bpepiW95RZH
0+FOXIHAgrrTqkLquMgq/UobcJIi9fkF4uxkx9vQQu+IujYmzsRIDa9TWdsE5RiSqIapQF0nTck0
kS47+tcPISfLYVMz7wQACk/e7M6Cu1KSRk521RvX1nvDXSp7NENykh9ormlnz0eWIOwgcIY77V5k
r83+W0KGxKZSsjuQW0/cW+2cNwH8AMl9QMi14nO5WvTb/rdEq7I/31CKu4XxctfyDKB6SeGO7Sx3
7vFk762Y3rjGmHgm12e06NKd7FDA8ZJTG6mesMBvE/XNFcNddgRE9yNUQEz5wE2u9uEmW/xxyJGV
Vtjwm/6zrai2DcBLtrUKVys3x4Y6J6RRd28cOH5WoBI6pMfcBVu9W+wIk54irfeW3PqhLOlj9Eba
xOx//fPtRV7WDN1nZSlKZ3Cy05u4OZFaYe5STQm0QHTIZGZWxwyIlbImk9KQxh+MhNwi4U23bOJa
aJDYm+uYbcnOlCLA42MpAxI7SnWEMyKW9Zca8OisnoqW7VSjiUZtpseEORVaL/+73cj8wRvFdmpz
towuzv4ORmDubypZaakPprFG421C+wfiJa1FTyOaNdnO6+vXPPNhaMG8mbobet6k2SmPJIfTSO4L
1sqq0mNr5ZsMGf/3Fzm8xPpaL/jcybnH1G3NHma6v6oHrHXcoR6vkwBwynxGtxv1VnizqXJ76CBh
AgPoGxeZ4xN/wAWEndgwzcx6AIzIU/FABtg3hf1/hsLWddLJAqKILzvH9RdaBLvfsaueBPbgtjrg
mrX9laIGkYHqN2IR6BaDRGAi70kYjtZS2kVlzkqPQNvnjAcm8Rnci/dzI3ROIe9txQZX9wtiWyX3
xqx4yoQPtrdUaz7UOsBr4ARsNLKc7Gyx13rENj3laNTerBPxX37bkxCZ/xgyUU+PXc+rjiYReGMo
+xzdA5JGFCe8nN4TyKLddUUU/S2FQrmaP33xuY5Sly146JOAPUJw3nCVy+PsLdUhl0WlYZCPND40
4AznfoAPeK2xgTxY2gjxJkgoY4nwMryvIIo9+5Qbsi704xI5AiBepCxXtHZv8i/SJ3HP03G8y65o
pngXGjy9YKUzR6llA1QMJT3d7ZsMrz+knQK4KtnNqtCd19lzsm/VlizbUlOQYb39TgK3dcCHdryn
p5GSgrSG9p9LbSagxcvKdr2XrpEaRvc/WSrOtjvSXfT0n7PU8Iaaf6zA39B3LJjzC603xoFPd0Le
GH5PCqzcwYaTuw3bf1Yq/goO3K76HFn/+YdcKwGM3oPEyuUiaE6BuiJtqlam5hFbOhdujL5P7IaJ
wBGkasaYNsW2Ag42Vj64kSVXNB3Fq2ejElzOkYwLFmpbdMtmTs2gckj4r1PC7hPZIN62Xz9g9ezx
sTU+VaZNlHv1ZnDVm3YIahGRjGoXJqLb+WS7PTuNg9jp3d5zUFR2BhlSZut0gwVhzWSRgsjVjCIN
KYFqVqnA9WTghbn/WTuLznQ6Vn9dK8mhlndxdDCaZDoNGs73u3TaCPaQMTh23WMYiUweyep3lxQY
+Aj5D2gl9wawRp7C5wbY6zD4oQiZdSPFldrbS1jvh1YlCGbF0gHZdDyZ88rXNCrheKrcPTrsSvhe
K/yNN7T8NE/jOtQRbFtWDM1461jHm3wyP+0QeF3YaSQLkSQdUFKUJXEG3qfvPxJtc/+0BmUY7/YA
IcgGfVF0Xl8+a9seZRTfxWHHMZMo2Ndmu9/lRPKWm3fyVjZ2MevTMKEBvENPFQ/irDKPwLnkL/aj
DNSS2I2NZhOXVHUCC0jNA4WrVSq7djGYBUI/H9MVW8P8x96LTsU65gFUXciBi3eki+v+1NR7ZFTw
v4DuCCqt+E0BRRELZYp0k2cpQmuoPTL8sQtlFYF9P35fS/9JCgVQXqpvrIVf+yW81GsOEC2VI/R0
ND3v2lCjkpnNG+5aNMBYqPlAVZTQarIcmwZ9VpmUxIioeABMl71yoN2VJnkyr4d/oHcZS85gOLjJ
0f9Mokh0OnXEy/9Uf8Cl9nQGy0k9OCTf/6X54PZsSI+jArGqvfUR/umdenPkk2GlsvAP1fSLNfm+
tXxW4Mq72R0uRDR4uIeSKOPs4sXGr7XvFM0HnTlyECp+pX9IRrsNUR7l1b8BnqvqUH4ZX13FCJFZ
iNbkR22s+Fbu6pwPyedTf4lMnUKTYV3QhdBJZVdB1gsBQTxlV/MvbfstxgComEnynKg/cP+MwHIi
XAgwHlJ0NJRjm4uhqo0/ydAhs5ggKEXBlss80W0y5T98LqFClt/cdtp1xSp6aONuO4HE/dt8GwjW
dojKxTnCG0zKNjBmNHwJwtR1ZF1VE8Bp7faQsuI1B//HBmqghylNWCfnpLFWAurIBjpNPa0Cgzje
R3WbCiQen80zRL0x64DDD8Q0FO4+CFYHkGpBSPYkbkV+qWJx4g3hwmIsZhwX0fH/OpAm2zARI97A
Mm5lzAWqRzzdJ3NRGLmm+SHZO8Mj1mzXRjWJWRH7miQkSfHBPjBPK09mW1IgCr5vQcXaZbzYG90Z
oMlNZvVmrsTipL1/DgeVhHx57dNmmjc3fouUlzlL1mlt1a/mPTYVvsIx3zoJ8MfgBB85PSiLUl1K
o3VhOwtgjJ5wuS3xuLj3Ss4ipxKzfYiT5BIqHZqJa6mS178Z7O9mTx2JCr1YMpXj7eqzKOvjASvE
X7M3H/IZaTl8UoPdY/ESHHC1tt9JouGIoXoYz3KA7YokGFleKXuZaJYHHskIcGRDMZBB2KHanmpw
2yrq8pBch24Ord+SDazkmAYlpTFkr6XvbLooh31ft/gpl6O+DVPBpaQJSAkJZ4wl+Z9FUviAqOgh
G5uxhAxyPPGEolRbNdCq5CyIZr1/UOx/+wCqP1Wfy8dQv2LN+iNl4u8QAQDp5gJOeyd0LmZdWBEc
vGyIegVHTEq8GpgbRLZ0WseCMFXjq7sI7EjgFA/qjvyKHRn9YH+oXIn2cj2ATc98txsPwdUC7sXh
0KEpOsEWDedpdYTtFr1Lf7LnqTYeKK3A4MdfHwyI0uuMlkdl1qO7+HOZ4mJet8dWf/mYCbgpKAEv
zN4SlxoHOEHq9k6w+D6HF6QicEkujQ00ftru1Iden1KsnEMAAEX+5nRsvzg4A2YjX2d7O1rIIl7a
C2v5V7Y0/eek5Xtnoz2hhG/30Md7b7UqXvjJZb6nYNM+ToVxNzOZ6EmhokrBu4GN7/f+Kz/BiM9L
ZunknPzHPIdJOxBfd1qHO7qVQYenN+uYcjyWcFeO9NxELOIfB28NB8L8dt5yCi9vh9J2pHfNjrij
fe7ZM9mSYV1JtjVe7ia4xAr9oT3TXESRbVikOwFhiMghawEmFM1h89Xh/v2ROd3cNUa/mM8GYzsS
m51Gstsdu3unBrOOt97uvjoCHtYLNJkeWMOHVDzeigyXphM4Fi9g42ZQewkBeXGmuhdAM2kwDCv1
yfO2YHuSDV1/B/MG33ZLZA1mESsG7duakN4PrmsqTNbA43HaK3IFSoMrmlVtLwNMNg7ciQzcm9o7
TbXpxuRUTxGdWh8Hrsf3VphN3AqBukwTQoQsuikclkl+viQiITDvP8OZq/bH8YeyBZAOysazG5FM
zhSeHbBNgN+Xr/9cmlbj8El4r6Uc+3WKgQuCipQo0lRecQPcu8P8xhZ1VQs2DNbMd3+HojGHlxhM
5yXNNOkDK+citUx/q8I95o67zXga1b+phjwQOUw7KBNznXtLCmxzFVAbTE6ds2zd4k6SKMCrqoc/
CnIJRyt5V82YNB2tgbXG+/rv6bs6glWAgvcDm+XDhSvu2DVEj/OQRkL8+Dm2p6zy2AfaN15wc4Aj
9Fjk43L8PhCiZhA7HyQrkRfpZOONi1JeaQaay9UZsFYw6vC2vX9KEN0/SCPnMDOwynPOk8XmJM7U
qAI931ZjTTeRidwQpkbbKNVG6CA89uroc+9atrfoPvKdGTKqy/wzhhi9jvwM4O7F7y+XGJXMOFEh
itm+v5RYT2MAf5ZwopK4FEntwJ5zXpj92DZdWJ9o7H3XVFDJMXlm88BKgEdN5LhO9EWW1fjIkXmr
oP1KrES+sE4eOmmSB+cm0++2fYyj29VPRf3t668A2m0E6KunV1x5RQ9iEmx8KmNCtQu9f9c1XS9O
iBWkyzzvNrEMUXGT5ExeGjhhUUz1x+ffaZxm4GTpTI0W65tnohPr6ckBSMmcsJ38RZdek73Wpwie
Yv5grNsL4gvzQVMGunkPo05OUDdqmMHpjeynwvbz7Ci0EeuSBdvL+IgbMMuzTlTy3r90owCG8g3Y
bsi3XcHK1q7B7e9UlP3nMujCvlWee9c893v6dkxahkB7fd9P4783fpEcOMQhh6U5E2W5tCnxkITx
mj0pplBhm0nN8PmH0izDJ7qgwsW5q6gWScC+8E4vK8khPF1SHkuhpT+YdhH2thhmGG30irkALdRY
9/7LHrGfwtxhAuBmj/3npgCson2cwA0ev+rVw/906dgEAvqJxKfalWWBZupqfzzw5/aUOtSkS2lR
Svh8uGuADOi0C6LZBRW91eOvwpzR86WLppfPYJdwiAUeIw3O1arbItm6bxKrDqHx/uwd7AAMoDBk
FQRsImfhDC6PUj0plfavoNxu7XfUwp3AiimiLLLH053QZTCB7JVwg0S9CKzfzA/0JNbNBrWrjrsg
zCh+mpjweQXg33MNzo0zB90yRZicXj6EoVgZurW/Y55MxHiBek2v6psUwc0l+T2ODsYa2EX65zfA
umsH68N9tVzCuVScS5VEQLECf/wJ8Mu2NQ7jjTy33b5w28wh+wfkUTWianIgN2T7Wkm9Jl3jDMHJ
/tKYTSe1ii16+SNuCrpQhzYwhUKzYU+/v7IRPK7LCiXrP2VEi+v7nc4YgGXiE+0tza9+2GYjGm9e
Qki622FFVixNY9tWxMdOt3Cmo/6+JCzz5xgtWt1vc6OalYGjDfNFOeTzWKPe1DmQSI62b/EFhRIs
ELtBObFg9Iov/uIFrikSCoCC/wkjfel0H1DcNawycnf/TRtzgGPsLWOieYfpfkY8VwgkXr9ZVVcx
f6Aw1hCk4s2GII7O2JupxROmqPiQe0WHBACuRB0vJ1GIKHiS/jOqZjFm7rx5V88dpN0bPE/9UrQR
ZifoLydrQ+ZeiBbnG+ULbpEsfzOhQvfr3MEnGyU8H6LgbOw9TGfyykCcLf3bUfA66ttKwRyNmZoZ
XqhjhRQDOEVsU7GneL+chgPuAkmU3+8mvg08gOMeJ61jjIArRsBK/sK7gpRcaXHjz60jxpybFPx3
ssJAIJtJMElivn/uzLAk8Ps6SbJcFpSXj6Nug+eHYx656M8X3LNBqqhrydCjb43dRNMqsmxvxTIM
I6insbB3Z5NIU7nTSiXNGr83fdzwzZykLAN8YwIsb4tQpLcQoVnoOZBq8g+9IIz33H1C/LGm99nr
4BlQ4amz7FlN85z6mQq5lopO6zGBqnU6D8+J3h9EeWDE9fT+0SN+Es+QsveAQwZVB3t5CtPia+0u
Hf7Zpf0VeQey3M0fDStBg95JMjow3aRDlYuGV8T2sf0NnesI7pNJU9Z19jWTShrxtAuXxuKwz7ml
cg35Xhtejhv5B9WG1FgsksXcdbZsRHmpaH7p3bGxb2SJ/WCQ/xo8FXF7Kr3yRrZ4bYvWs5ahm+MU
iA3MUghKCRaNIO+592Qp1T3gGkzMs8Kws/5x1a3L0yEd9+XN4Y6z0QUbTOG7rqVZ23eIIPx2nwAO
0NzArwo0jNvroSKOe6sqHrKVJZ/6BKiMMxS5bujrPgbtJR0OOTelB29cXF8gQZoTR50nvoBu5WZM
6ptzrnPbfyEEJXS4LIHWY74v9JbsjEOLqu/xvBNh/Vi3j/OcHfAKekGRwMWaqRRGbkXB6cIkhjHT
GQNH3glCiiO26ejEiEOkMe8sVYNNPK4VkPpj1JTn0r6z0ESm7Ydltb7Es1ym6vfuacV7hg5uYhld
jvEdi7rgBXjLRJDCY8tJRvhIjEvY5+WSsMgS4JyXk9FeizU2A4YEqNyG3Tx0AlDqHTPsJc6PJmEf
04+kP8q13YRJN15sE1KhE/PmKcqqdmGQYPgUII/enNni2fSdH5qzkYy2dctbH0l3gglpC/w1lE+e
ypXKtzacMn2/Ly1kLjnvU1rnrhukrwS2NMtALS9Y7Z/0vUYsY1y8HyjK3NcM/F/DtwIcznNGgT6k
kQutIzOqGCKDibelvzzdnj5ge6q9wIXuyCJxuvAyXk8zOS135c/dQ4y25luIJtSKX9CpaJ1aXrg+
D3a+TILCV92qBcU6ZgZ05gYY30r+z2KFxsJrsaTxYJg9B0t1p8vCUhOFez7sI6+dQaAfqEpOAJiI
YIEbnnw+wGWT8WcDHzOn5iYpmngacxwuZF0UDkHnNR8CAbbroSg/crU1zqcWFjdN3J3oPXtoX0wt
38e7+iyJXdZJCGTYNwk/FOcIHxFlln+F2ASBSY462eA6jD5M0gKOonpoBz/au9ekvXkoE7UJ9EzT
aoGPKdWmrHcOTKXJXT39H3D0m+85R4GFjHWE9DZPr/zGzI/eN1rak0FHNWF8F2FLI1dv1jLzauUZ
V/cG3ptJeH5y628I4uDu5QcrHMb8EQ72imQJiCJIPgGK5ArwudxP1k/3WY6/+9c1dQtlRYJP783t
K/V6//p66P4ebGVhj54nsLsbkKdg6AvyHw1JZOOTOjIZnW7l7+X5wrxGVDyNsl5YRfqb4dGGajS4
xxvDupQwjxHnJ9wBkfMwJsyLry13/qjBfCfU9I+/DZARfYY+3iwOf2+78W2AqvC7izO2QrH8TDly
weetmX7wbrrspohax0kDbz+0jW75cY1Ak0XIcDT4BJM5kyCWbBDCSgBmeqHV9utAQuAWyGZh7X4P
SjHRb1IOPHSD5pbiY7/Nu6BL9QgvyA6nXCEci0KC7ReRfmb1IY4Z6kNaTbDhAA0iQhWDTesAvsC7
HK7jupPcscTnyWcKGfIgCukKK9ZGGEjvV/EjLSdudq5aWHkDeZ4hi9R2Um3eHhd2tmOrpRv2jD9B
aTiQp0mp6qA1Hjakq7S3/5aDBaD0R9zxTqNDPPXl0etljZgSRq0+Q05uLimmJF4hJ4rYD6Qti83n
TYf4Am8HVM6a6w==
`protect end_protected

