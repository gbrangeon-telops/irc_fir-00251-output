

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
q/LTCQu22IewzFL2xoALv0V8R0cS+n3ZGOXTlz6zO0tHpf0bhYU3nG7YhbNw5H8bMFnHmKPTo6eG
UeGsZXmzfA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
RYLOlBm3BPRhwpOnNgJH4Vt0qZdXkt6+qKeUVOFaD4rlCQUegbI8dSeedwyfmRhRBYYfcasAbBQY
SHt4NDprJvJn/h7vAd6X1UjRiIi8OF1s+lR2yqR+Y5n/Ai+CRx+BajVy1wGHxdjiCnM87Cq2Hq6s
UytlPbN46pRkluJe6NI=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
5Onxh89dWZfdY8AMW/MOzaZUaP+doVdup9B0riUkkwljU4WHOna1/K734H9kkMqSDTQ9ivkZIsmH
DErXjPeoJcAWqHloB9UX56vG6J+JtHhxXpnFa4rDUsDzFadXGZZrXqt/NJt/7/nP2AP1p1qeKRkq
ksYRHunueBYG/B5LuPR00cTpoZaaCYuJroh/pzkerIy/CPNX1RAKt047HCKtvFBXH7wuqo/yaUyk
Xkrxw2AQ0ggYgz1hK0KOdWT2JckcbGgVwPsik+mchcvmPUBKx8qFAnef+ZSGsUTy+3gjDznrQOsF
sJM7rKdsAjU5OLq3k8BWR36ur9hbMdk+lvFEHA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
fe81XuZ9RrG7wwwI46b8GZQ5C9RFsRlLr0EzhGvkV3ZMeUUoQPwYfJl6GHoj+GDA9GnY0KeJe84A
xt/fhvb4h1DNhpVnvsOo41gu13r2msE3kvHyK8en6IodL/Mdh8CmalY/a7ZhDb0W+KP7rEAgisED
MHKHkmm4OWbTY9lIJCQ=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
JHuY2RJ1GBIZ6g9aWOE7BqrGN8uQypqLnY0uHGFvCX6msmuceGWWswz4xbJBwz2/gb4ZfVDTzfAB
RXiuZlDm1B8txxWQYaxO0lZYlxtzCU/lUn47fRBxEhyn9Yc5lQx2oW3B/G9c81S8zCONQlmapnrX
y4OR/jDZXLz2wxMs0tkWUSXHisAbuRctLOTsTUfqMDUsJS1g+TDQCDpUDXL43sWg1LCRd7wDn0um
3q29OwHxtysopGOz0DxmTcK07ZEEnSJS89piniLxLQC53j2zOhAk7sCb4iRKccCVkkeasTjlcMTi
rJCab5WZRXi1gu1yWZ5s8tCfrKbGVSZTS8p+pg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 57216)
`protect data_block
GUMHeZ1V7ePa/OieCwqMo3AAN7YA+4X7oTigVWDt6aDsEyeCR5VdnjpczSTVE0toni2pU/tDxzPN
mk0gNvLOej+zPEJk1py7BhuUINi8BI3O9xoNZLWtySczOlHeHA5pgK/zyE+CztTuhtJz7qcemAf6
+7tqfyHi89uP1CEtxuJYBiSGpsTvYiJijCxPhadZN/GW5Fe1mshKFPky/Ekntsu+s5hiyc0HnFSX
89+Aeb/Xmy1GsTQTOeIy6NuZrVavD9gcsaYJNW2NGF8YZbIGTK+1TfeBdM83gn1e5qYG8iyCaflO
iQ8FDuwTYknr3ObhIFSb6Kaf4upSxAzgb9zKOkGAGOyyi9FF5b2t4tMeIDKPtTky9TQ0aRbzeaCg
UwJpixCkTAnaADUhLkEXEBMFpIJAMAqMsAEhlyE2TWftc4xRl4HVn/KeNXdwGWDyljuR7dhiy0eA
6noomxzQwRetSuD7k2twfrrRAt3mqMLvGo30JfpScAcp/0UhJj+hc1N8oa/t6/KVYWnlaevSYH5w
+EqTB/8DYwPpiMaeh/ponUU123ra7hqaumpm4Xlwf+GaspTWdCKAAkQ0mI1iJCMNk7YgM1AQeT/N
Ipo+twfqdJQ1tJn5/M0fjFfjAnyXbv065yqV9I57SOOnQAhzzJNR+/5qC5X3TfwkhZ8I42TvQn+Q
mgG8/D0r8brHGeq0kPQGDpf9tXbz1fUeHp/p2DW2XT2YDYm5nwX7xI56GdPebSMHTuVUTlSSLMkT
5qfOBkXrTtc/0lBEV0hjfG5tS/gBle/xFjxSM3wry+BdSh/LNqiYJlAMc+wYf52uQNTwWR6LkS4g
JAZJY+dnnzziXv727mMBGth2uKZb3uuqWGqN+Y5f+OGXwp7o4zCjHHIVAQq2jnAJIbZMm7aCMmrv
hxfCfuSSPI5pzLlDttHuTNGc2tfRwghKm0aEwJlhK04bvt4sgeBKWqrBNl3rFea7RBEBYpfahJ+2
dNg4XomUtXc/ZxbJEQymcndDTpV4ZktuWi2o4Us0V4GtnIe7Ju2vH1oM1TLkeWghuBG/hPE4n4xa
f/ntWjPit8KmbZGOjDuZeSEuZuNXikFc1vjmy1VlAza7Zu1LtmrvDphUrB5iAexmS4Db2lDDJb8N
E1wjIudtO8D29wzr6ZnWrC5njC/Dc1Mj5wujo5F6GsQulkuF5v8d9i2ghp+YpodDgp28Ctvo/lVN
7b+AOVLI0l4aPg+W4bNjQVTAOYnBhY4GkK8YDFN8pfXEm8gTKSRDTMH3XaZbyHOHgA+cv2YzB0r/
95UM6wjcRY79nSpIlSf+DuqrZStUQfCnKfKDpcRY6etn21g1K+RX1bvULjj252ZbUv66lsP3r+Vd
W86116yv+t5Gn6dYlWmZTZUMZ5Nis0PPyW1W8FQXyssxxV+3Fqjkt50kIKXwsiJUfulIMJqjBUEI
naw/LnMbFHctj1uo0PJar58ZaSCk/pBSnUNMXG0OL8/DyAtLwA77MVvMiURcj3t15za9gevGH8NC
Pv1KYXbC8x0YByTn6fl7AhM7T6u61WcNdssZZlqDj0gWjVc1xT4d+tTAMeo11tR0ZzzSWqqPmu+P
E0AZI4GPLPzcxfEYM5ZmvRZY18ewCIUvyPxiyNnecEuzvcDG++shJW82TDzCxIkxjiAVyMhsJcuC
9VNVOWdZJhSTMB9l8vRFcKmR+geRDVKXEp8sf5lj0bnafmjEpE+zBgPvCYsHpUVBJ286cZhj7ZfG
8DJ+VWtrgrldQofoZM6Dk5tfQNIQyG1gTEVs/h1lZUZrMGE3r1Qk13z2XOZopJzrWoSollATWbVT
egEWxuu9ltVcVmh8RuUPSupAuH0Tn5XzOHQFHB7/PLs3f5uvpdW+x3QQ1ryfWpNM84SvQyev+Y7/
UmC6aFLmDWq4ujifJBTjYUKbm4lMFU2IIGNRrDj7xfHk4twzAy2JQBKzYzpo2ei++Va3h4COHhwQ
Q9DxOxlSq1pVEfk3oFkzdFpPRV/0swV+1b5ekBTtSKZ9IZWhFY5fYDk5ltpEb24s7RH8I+9yJiPm
FdHC3bkeyxTRYkS+XCgads+gXEZQP5YmmypG1lncF1vGaCSqb50pSOnJjkkJgrJaF9h9QMlwq28w
/lgu2IBRB0qGQOQmsj8VWEQUADrXfY4s/ZN3D5rvtdXRG0SM8fJCYVSZks5ZdCx4/YmnD8dGCBTd
wu2xC4WRiDRSG84hVaec2mhGizvg5sOu+ztt28zhejP03KP8CuTDxDTbUeVZnuFyq7w+f7GiXWKv
Es+nE90dzm8z3XdnQLPxMGYJbsuU94db1Wtbm7TZRhcr6aMx4/V5FAFeYeX0AYU6c870lPbNbJ55
NdlrKD1XKpXry8qBJLpOsATX9UNSExWh646RnDkwiHM5JkkcZ6EoiUUiAM6H8PyZEna/VI3TaMRA
lU8gRS6B5v3OaEvtY2vib6WooFnxJJyGioeImxWVD7dbbURScTr7t2JTZe0CuGLDxCey+4C5FOdn
wW+Go+rZSys6jPaGBMtW5CglPYxuB+louXXSXCQqNYmSEAsDdVtEXDkSsBjN5yXjAqygJsx2nrC1
7BSmX7SPM5ZLbORoKHE57kjf7TwU16Xs9a4+f7IejbAqbuzIsUBv6X1CrM4eQtl5+xbLs1KWMP1v
yL/2oz4mJwLLjM6nO9nmOfpc+mMpgc7CFKG0A+/2TK9vXaMeam20zfd0HUWAQxGfwYMj32ukUMRq
FsgYoR+VBUGa7l1KutF85+Rn2VKmFlidokRb/RwoDMcz7SHBYnqjNPzbet2632q8JuOdowg+w05+
erRRNd0y0zS6lUlv+J4Tq5EeQxtp72mWV+8dHkmT1ThBTZ+k9OUgMcQJhWV1/EezHLjTWtg2+oA2
NbV5A0I3ZeOUvx2sdr3TjsF/WkDl4CJTGEsBrIHC4eJpAYRFj7GQg04ff9zH9FSPLMQa0J902IA+
W6qGy9SYj7ZdXpNFEaGXpZag+W0UoL9x/Ad5GBLIF3bRXxMOkvQd/BrS3s3bRS4BNsQEyEa8dwFn
rco4qWJ/ov1CScD8lLy8oYIt8BWhzfntQPzJG2P30Sv8guIkb/uV+N474SEZ4sV1DJquV0gxJQ8r
7E71ra2iVU8MM/BPacfJ7SGeFdop+ym4YVPWBNnXk7DrLEuYjiM/wKF1G6RPWiHpG7wdPZzAIYyL
cvQsRZszbJV+6JDDtGwpxZdI+tIBjZBsK1+pMtrYhkk9xkp9P8O7lmVMhzHsEPDnzih/0RzlIxWl
xaR3vsLDGccS5APW1msTJQn9cMiISNrZnzJ9x5uamkhTEHrFXQZ91ydmRICSi1b2pKRWVQ8sILub
4vuwaSsvjionj3U2VjxJsxXdTyI8USiGQl9D1X9HE7lZE8kh6tfV8K1RmEyt0wHDMaEMCKLXBwj8
xIHktAOjahOTrnXFk0b4W2ojvMUPcTquOj+yn9vBDTX86CkmF0kjoPYxTljJBNVEnjtQXIMvVCJE
UeI83earuM479IoEMyYi0w0J88Yo4Gsn01QLDNo1TJkOiTSYQK+1gseguAamshmy/sq4xgBDKV2y
I1oZTy79/K/0MumXXpBJ2wUwRrFafTl3a5EGh6y++vMfKA1CGoFRoq57qn9cpf5lB57fAWn9k1l9
XCTsg9CZR01MXVtiOleUk3JTnBNDBSRABcI0eWvTxbscdwqDBhE1q5GtmdjaiLpgbhlPv+5KnyTd
/gBqDzkAhr589WrP7VQJiJrIzoqiIOt4IBh+SxBHU/KKZK6glod8fQ4OLwgWNQP2D8G9An64WPq6
XDa9pFTmMbVDrJ4UHBWb9l9umrndLvEbx2pR0t2uw92FPDuGRtUypT1SrQ6XAmo9V9eHnhPyEEid
lY7K7p/4nh2dVfVdhSzsx5AsVrJWt8NF95cEIbgqI01vfRkBJGYGQHR9cru/lfQzbnWDJWigPyLM
FDF9JTr0QXtaY7g7UENm+lw7dPym9198Jw+MylYv7DzS2Zi+FG326Lzi6pPjH2YWBP6aeSBj7T8i
Z5pWDWV3jdJjgZRBuqZPNyigvD+3FwLHIcFbuzK8+x/NuuOMjhDJ3R6PswIdncxI3a+aXVtGOe7G
Cpt9ieKVk+A2m7Sc0gi1DRWR6HFqngBO5v9YX57tT5Ok5cDFsEKk0AmBwl9ZvB7WQjZecfsNQ7Sr
SNRUyB27qCNzwB93P+mivR9pFVcGjo/GnO2sDEhHDQbIXRN2K8Mp6mTkiy6Sq5k+P8XcPctZ+unA
nLuFvaheWUzIhfPSgg7v8gXELpiJVKxdrGCXtLvLNXjcYefvNKXXPYUnQih0cfgDOQmPqvrtTA1W
jNuAu3JZAuHiKOEuqV/S50PmAnir6OLQRQJzrWMdoLjT/L/8rXhKYA4tClsul6FBIGWPqFRojGJq
BqpUahj15zx9+Mh2J7/ah6QanRASeSA+Ln+QJSksDCrDCN7FXriGSTJbEK+qoGvRIi2r94hzvMcC
7KxAk96Ld0Gaq+yplzgaZ5p3aBINGzEncHfTQUWXZSwGG0l6IpTNwvPoMH1lb4ykjfNt0aI9anps
mLulFhCyMsD8EMpa/76B+InWnHApvlRneCMjMin/5u8vX91eBVDM3q+UbHNhJ0JFOOVbbKtSWr+j
nflsWiU+qjUhdlYxPEMCjNX4l61GUWyIR5Sq37OQJMCPLi+uTnFJ9waKeWanj4cUu/9ZCTV+LecX
DhSO2hLXaMsrMnNUWLLQsKgrLZ9kAg6ldjMGjRkFPxpDb3QQXCgOwSV/elR9UFCJbAEezfNe+dMH
E5fJl+axjqc1CqNvWvgDvVDVdqkWWre5c381E8foVYeh73EM/t3Y7i3FBT3DCjkFO1AwZw9FU+st
AP0s+9e76SQl4qrFJg25h/MLKM4Y4P6atc2YBb2M1ba8AZT2UL9mG7dHxDZ2LaUmg4Phsdxd94wL
VtoFvJsYsUevoOYs9tSRvGg1pbeXySnAz8BCKAZ9EKEsO83UdqmYSyxEaJ5Iy0tGy+oTZHLu8QC5
eZHCDUzs3snEtVfzb3opkPHGSWF/Ly5oJSbZzydoKLsQRJ+h9u8hqMsXG6l66jdJ3gToaxQcljR8
oFLgUsaJO20Hx/u88zZeOTx6wjSIRZb15LXMGlGdvFZWPbD1Dt9iCQZ88Yhqx0k96CLauAH5t1P0
EfYRe8D541/7StJla7dGEfB5fwiktS9iFL+fnMQjJh3aF9qAIICziNsZ/Jcaj+F03esRlUj4Nzwt
lKBATxFICGdcnzv+mi0ZyyyuGN2Jj+DlPt8FgE9xJ59x78ioH2yAjsnTZVFI/QHxpv1Ih+ZZFJzH
vaWRWayM/laCzb72e8I86TpYdWGvn9pOlud3VNII7eSexeEDpOMCr/a8qZjTJOGflTK0qtnkv+FX
h4YaD2gGZAbXw1WpB9dwNT6PMOnldEZ57XSVsCODGnEqLxbaRtLTfuFkviYvr8swYU2Zx0LIefw3
p6FDSFJBPIT31/4RLCB11Xt4L3ED3VFTfZzRCHW5PhMx1JzIJEv+qJQPz8+WwuNBLWpkCzzCr7BH
iYIGzMO5nZhdZIVrNP3MddgMMim36Spj4FWIkPkNHP052g/8leSjTA2AbomxJIfcmf0+4AWuq89G
0qPiftJG8hMIblWiKhnoaR2fJ5sWJy+7ZYe6cxhk+ms8lz+tOrqTDR6+Jg/NvTZqaZKV9ENYkATN
tffwx/D+byi3w7JQak612OvGyx2yLGBWH3SCwCypouJO8QXe9LZ0AXR3OJvqoi0DmiYEqx68Gi6z
2rdKPcc4RV6+P6HOix4czqcFG91gAS601aiC8JUjpucsAGshLLdEuMlEM5lnXYEDwj9aZvtmI+ip
XawH7cRO5zjKnL5Q/o+s80gRhcFf1XD3oDppeambWZAz3fgSstgWReEtC5hizVsi/H7xYPxfVOyb
xNR1wdnWPvXjatBuW2rDKluQlp6Omo0YPUqErxHbHboRttKMDtv0ZR4aRNGkCdryWaOEVQCXu510
9V8OYCEgVqfqklnK4ES6POw0sNWm0abIP0JQtm4ic7FeVyQFAxD8htr5mP5cCyjBwKpDzQOJylmO
+AaxdoYdWSVufzDYOP7dWQUaNA70LjqnKHjdEfDUAZToBS2y+7E8zks4vPFi/oJdKfvuSVN7mPvS
Ert/1W9pkPOoGSRzYq6Deqg2+X/QM9Olg2odQ9uzUEuI3+8jxZxo8YgTe/xJBFppFfzL93TSgY+O
B6epIzDGmjzfPdM3cMRhmESWGXch5JrHgvRXdgULfxtYbw4YXTX3uXWpoVGGt0fD3TB95JhfPIZ3
V7fg+9WixdJ71hglgTNJUCr2arsny44uUicPo8MfW4imBmcQUoJ4w+OSsp81c8X8CyiBzY9MnNtz
eHGoa9ZhnP3PVzgyBdFPV0VIYdfsGT9HeABxjsmWazfHuDZfXKBKhBUPNVJz3sNCEHJ5+npmvYlX
f1cbUgd6sNQPOTT71bPvnwIeP5oTJh6sKxMr8c/ZS5kByiedoRAcLTzTJX/6DAOYW3uBzUBoOrJD
Uj89ntSAxhBm3/YLD2WzTjBgFBNSlryEyCxFGUxH8JlaVfH3wVCeGERLMwbg5gV57oxYtN80gIow
94x5XdwosoQnI0HfWRI8Xo1IPZP6/Jd42y5jsLnJiiI5KspKikJuVOpyTYWZuoc+8GPFDNiAdle7
MeHZS4kVZZnx17oTKWViEWv+xWN9La+GL3rv2SnXQR2jzIshG1TkwNA5ZDNy7CuFqPQJUOrnBOj7
XOl9elzZuzHZI1XhoP0hK4NW+u2/jYuy/DU+iknpxY6fBc7hG/lTbVACrbsfjS6ZxK2cWFwMY7DJ
InmeMtMDAeG01NhPxymkvo1PORJFEdRy5HsT6bpz9T49BB4RMOobX9VBaHAAZEAOmGz4auvqjtzs
JsiFLLnMlVDci/KTk1eHfcWm9uFjg1TnLWA91HsTB+SmNVutSgCdjR/lhp4S8PaQ66quAlB1sxZC
umIxBTjr3Og7xFKuLqW7Z04u724GakQh+h5RoX+biQIxaeXb1bwDVj8dIJfgBDbPL8vgHS2K3ENB
pB+XOQIZhOMdwhm2x12XZg3Vm+rjbvu0MzJT/CDz1H58BEJo89XXZZ8yWOluqA/+ajQkcsQihOJb
vCCOvZF6nLlcjYuqbcjNK5LDNyF9w6w3kyfZbkSk05eXv3uEi4vX9YcJ4HQiWw0J5C+F5NIARp/d
twgVbbFl8c0VVZCpJvLTuMtevAzs5fb5pYYCK6gHZm41vWRj6zrsqCDHmGEjDWOHIJkF+r/yJDXh
/QXY0XXbm+WJKPW3ouNrgxpknhaMw2fEKXHd4RZB7zlrA6m/GJR+c6lRhNV4B4SWqJ6J3h+6QXD/
nrsWRz0mpRMACmdd/PZsq3L3IzbM9/2RvAxg0rPS3zej+R5K2DuxcPx+FClhpRBUwg7C8kmwT6Bc
PT8Hm0Vk4/RzFby5A2ZVn/VGzkpsqKie03gn/kST71xZSoECB82jMVOVlzaeWMyc7gIFEFsUyEJu
SEHVwBHKmmJTRPzZ5qlhZEz2ghGqngIJnrXUOQOPS9e5Ym6QrSBqM5OBfmHnYivxLJh+IDAD+I4/
f3Cje4yGn4kIVvzo+cFnPygtaTnEP6XMnpcEmLPFkoM6E+nFTWyf0DjxB6WW+0digdKIvPCSE3qo
uCQKNXq/oTPjKqyyj6cfBrsGjngb2F8MXo90oIRZP9TbG27IwIOlOm9F+GWDnlXEAh7tAbZDt+Wq
u2B6TpYQyZKSnlkONh+IKA26jRx4CRC+RlOd+KB/3PMbNCpJLR83VR1/OynM4tl8004Eg3DZDWfA
q/0QdCvSMcSvY4om6kK10gOa1xUWcQ5jfOFPOcJknaMx3D24d2hBYdkinkHSW8a5CLbnTbmjorwB
x4vFFeiau2LPPX+bgwROUrfGpzgvO6ikfi/lo7tKxE9KAYiz+96uuIpd7Hu9oHpz/sx29BlGZE3j
k9Mt8KFAO94Wnj7QuDdVCjbTg6xiaQTGdvL3kkwkgBVkUnvM2qlxM/tjgHOiW9Lo91gbAvS9bag6
itVUVV9zuOsSkBcQ4VV5XaVLQQfWWei6MllkvCerVb3UdpqVHjocKarRnRbaWjeaBIM4Ve8Sca9p
fiMF6lbz3WVWtGJKXuOc2g1MotRAbVdwPR6GYV2Otem8v76Pfh2wzgvI2sRCeeqd+ByFuo5faK0e
Jy9MyxsA+L7Vhs+fLr0EnAx9+zZt9mhFF/XM1MPjEYyHGE7dU0W+IYTt6dzLSkro8Wj+9e/tbJDu
zzOpmEN+oI2F0m20Wm/Vj7DqhiBzZFxjyfJV3uOGO+LMvJl+27MzFDXjC82JWhS+3KmqQYi47DHe
xuQ+nuc1a4GK/LyKWvQ+WG75iR5E1Ua3h+t478L7jFWqcsrqzHS2nhfPURTpOpUjyHzgNEQkwsh2
dOMIzfnGY9y0SkAGup30Uu4t9UQcOGrMackr4kOcJLz42EuCpDn08UQ6JQXvMl4pfxAkIGzbPnT4
lNSxSDznkT+dnuLpIheYzFgTLYJW/LrLzQhRwumoz1ZE0VuWwF530M5b0P5TwW1gIza6MbpOlCEy
3AiJqvKuQTzHkH4R8UntGac7d9St6E7/CezeV2wi9AfLDHEslI0il0CYRBmv1XpD1O6Dg4Xze4/Z
upk+G9SALGkAOgRad3nR9skzCSsh9DObdP7MEoKxvu74QpD5vnSZ4QzDcHHvFOFUC4/6T6EOadyo
zDJn5aKyosqUcxAQntt41LFRqUXQkMBjN1GNnG3C5rC3MzhNo786s28/8RH+4YUu1S4cUY5JSV1H
5A7/kDlH/SUSUH2GYYAOAJZFz4VZnQCS6lTBHN2pnXopWAqy8Nu8UT7g5Se4lMCrEjqLn0HVt8NT
HSqzj+OA1D6RdaKExCgrQvx3MtOuogVWzxMpmwgKGCyYWIRGwOAHptsN6ig/rKs7XRB7HfOafSrZ
OHyjv7pVtqdzhLXUlYj09SIeYKMr2QNDRnyn8m7viVqp65c8gPGXENjZ/HAD5iSPz4PMv+2sfxbC
DzPjYwTOlgvaPDbv+yW7N0gjzxsGrX0/NygD6tFnHi7fKan8L2Zyhx0KEaKn9z9/hYHpcqQZRhOA
+6tjDsOHx0J2aFmTB5Ot32rkYPybm4HpBfq6msEcsftjJ5FurVmw+lp+QWDSULBmC3zb/9LIvooK
I9Ai/VnB90p//rEVlaZXQ/7qUOZff3z0Jk4yYFuEzhopI65JoUUM2ZWO+xYoytGwCcV4Z21G1zNW
5F8nujhj9+J10uAvlZ0S4BD3LUasAJURUfFnCOVklDp12OTuqq27+pQakH/i3W56s7in+G0c2/sw
cTjg3qo26S0QEPhLaHA64CPn9RZljuZYnHD5ouRI/+TEE4A+UQnzdooBaJUiFCA+0gkoQT0T6Ezd
NsUd+PK37lrCkfPSPUkDfzRIBJPVpVUkqlyDxDyilBDE5OJFQMIdRLZ0ONyWdRofRDoL1OVwxqpi
QY+rO5dEnXMjjILcMc2xp5cEtu0U9nL8x3J+FTc0LhK9XQwBeza/KXDO6uZZ0aZSoBcz9tlmZU8z
XwtJ22lT3XXTMMtJcYC8kYxaRQmSIgronsDQtcLWxXU0rwYYWincOHwhelmTb4ok4kC6Bigc/Ltz
OCVLGvMnpgiJ4odoj9YOhdGiljWTCMCr1uOv3ltpgDvToUPuYoDNamzpz6mcaeGHRFHI6ebzVYne
WY2331ICTO20relC+Eyef+KyeWAw+WZTdBQHI97AQqbVtA/K5awhfqEVNYm6tQ7NKJsQhDJn9GHH
Sl6MUtdsbb0wvtTaUm+njb5Nppg5cHeWyv5x1sd5FgR24e3cA+QNnW408tBvqKb+63NQ0LCWZGB7
h/9XXchBsiZq7yIoR2pJDwVv7s10smMEQ91Fy5beH4fbMCJfH36xlshz9WTsxSKLwNHAIQ8qpcT+
X6TKldvB21YBEU/qMzCFEjOkasaD16N5gmbrUmilw+kgL08jNJj+tal+0gQ+WQX4kyMfBH9/PRNP
43twMS20HNUTrnr5rPeQF58j8/RtN3bJx9KqXk6f6NQdvkXWkCKejCLNZIUj5PrvjoHDuHv48CAy
RKxPfEzDgv4tPoudrtQ5LpEU3UxJGADKm6+WVO++A0H8sc0ARs+uFq10cDYVyyVG/Ou6fnJC2Rsd
Tb4rJZGpBjih5bLATc6Q4pYL1m7AkU48K5dTXtxOF2jM4mhenTGhgmG1IFUHTM309LB0aKB/ARpw
VxvSMbEVphOj6rp6SffZiddGV2HTRvQF5/69ticNgohbPPB3bIj0+LbSCcF+VtKOLqzG7fRsK559
8id5wkZQyQOVYXbC+dcSgHdTrzGvnaG3gf31L1hAD1CAHiEl2y98a+O84xv+UTcwLEtjzSMf24mt
tbT7MKzy5akogR7M4wZeq72q/cXoMzd6YxHvK5je+HaEZ9kt2h9uXEa9cQgLCel9rpZdMADo39bv
4K3C8XZcZ19UeV22h4uHYHk95wcIlS0mv5oKCMHy8cgzQp1aMYXTyhY0RCQpym1Pyzfubc8KlZJn
Hj5VmIB4WYR5XzTjsjqryQ9+7NLXUWqaJt14gNFq+qu64d910Kf9WbiJTHb+33dTteWnbcEg1mM1
hi8Ivdgz/aF1cluc4J4h/BwG90sq5xWda405+Ht2a0QMK8LRQafuECjdQFDsjsUtXLsKkCSemZ3P
rwehzOsIbKVMxMe5OUA5ZihZBlVx8tkdq5TdeGFWhmkW0b0+l1Y0YazbAs9Pvr56VfW+dgNA7+KJ
NFROfYuxM7WVKunekRm7U2Ob8e4jvyNlYN2IvCUxGaBfTf1YBy/hwOfdNoIvPs9E5oYkA6bbFPPH
iECoX1k+UlwfDM/lfIJb+5oLQr1UkEgdkyvoLD8tJpEZmhyCwTzoAwKvuDpwwK+jNFVQMZ5wo5HF
F1Uwsmjwme9Le6y+vRaYFYC6npbDmT5u/CgoQ7D0A9wiAfMBFZ72z5guY9FBdekDXyt3R3E6ewji
ogtm8POURZ+ZrpLewTP+UARDAYaDASbOH9orll63W3c96x1GUkEGdvnAtFx0jeOyIkP5ZFPJZKJ/
LnqmHSA0bmXBDwqc4Eo5OdDMz1JkSYAPMBDV5EgWdsu1uZKUXHIRHPCrt2OCrVp5RbCuKcC8YbJf
1ufCtSAdbhxtqQG7UUAwvwTrEpPz+nMb4+dvW0OxWm3d337d/hhaUti6zuZK2ltPt+kspPcPFXUZ
doKWLS3bVsPZpce0H1eNNoYw/T/PGx147bU+vpkXoUnFhziURh4Efyybb5+QGynYAylObaDWYQBT
58dJAQNYO9s/+BH0EBNQQlZ0Cu7OVmF/MbLMcQaot8pcwQpeJ+yrMKMGp4Woms77SHemwuhcsWZ0
qJT3R+XwT3r9pMjoZL4Gmwq4D36wMWQ31wO3ENAtt7K5dg4V1QUoPup8XTMPrSVgjJkt0MTRmrne
DZU3n+XLvWEqKhRPzo9Ja9aIxhYMFVHj38LoxWHsYIHvyrYH0ibJBUd2aenWEI9U+7Cfa6zXZtVH
xD9ep/ORiG9TyR+bLiIuJ+OaIu1XUdH4IW7UMU67pBPyqS6v+SFBaTSZEnmLxj7wTwNblMW8EUIf
76BLy+Mk/y7bziBtCO1XHHu1yBm+ULNPSAnKo7Ym4uqC2RWIY//sNCROIAoSoW1YJT/n6F/6g8/g
ehVGFnLuB4MB3s1NCfJqmlbPSJEhwfspKhXzUbLs75WL01DGwQYSYMPQtc89Y8gv9GOw4MJHNzxW
M6a//uH2vMa6b768RT/szWbwrTRhwdTGhIHCSO9yW+32tkrfLYK9MXCxI1c2yIEfokBKoMKytiPS
MU81A4NBUmF1ITc++SVCkOaLbiUmRl4lFoYfPFkyZ6mAguyepnk0IN/8QchZKofo87igpgzHbzvQ
yOKQalkDJwna5mCAmhRby3mw1OL0mbwxoXUf1jlYgEH7IgzlCt9OBPyIyq6PoBJS3zshbaS70k7O
XW0Q5kx8drQxVv9p3hH/5VDHrkEx2dg1no4oL63NaVfywZtrxqDSS0Icwj1DHPlOC+A2Ul+rF5m9
KExg4j1/P5BnzgEiPJLi4uGlSFsbXvXgIiQGSpiQPI25qgbxRvnouYyNpAJ+/S5M+0TV82ZyEIhl
HC2uL67DUOxWXSgWav+5C2BjXVRCQ450Wq33S1Zm445qbezCcq9tSnSoMzZKHtoVGO0LSR8YF3ns
bGQ6acUIBAc3ul70Qx3eiVGDx3vgRU5S8VTJpe73vBtM/5/HBYyYgR2YKR5hZ7Mcp3EInT2GozGO
7bxpNKT1pWuO1sw7lWkLqp6/1b2z/hVx5kpT9sXhVw7tjtOd7AGKpfCNArLYFdpIgSaR+Skijob+
kVgrShOQEZ0+0VjZfWQjb/4Fz2kaadfNfCFHxGsAVhTSNEAbPMHZOe3vH0yqruOP8fYmqnlW6A80
t2PvqLuG/0wbBEqF0ByueaMOYWOpA8R7iuyd9pvDyssUyDZCoViKffcZtLOafoXXeDg316AE5f/Q
HFQBwrxsua4uwHOuKoL/MR3sjmFJ16gusl9Qss9tqTddxcKWvhGtTbLcM3DOGA1ZBWRgEI1VnrpQ
r3BbWfuBG1CQC2KJ0th9Trm3wAjdnj4HpOeGKrTqDtpiZ93/TK73uomNGaoKi52OABdX5+QESKGY
gwJjiUTVK+gnN5oDJGRXcyFLjbuPiARJ9h7CyKMXvCpc57pelIE/Fq2Ty9zPrafIJMniOM8uK4H0
XuP/JYJEDr1GZTdPMUCQSnAjgjCcAmpdaVCUvWkHRfAsG1qJ21L2pGjNVG95yM8iDKIPkCRMn9PG
p/OtrAWsL51CrrzGtjipvywco+ozLcS0tftb0ycP6OztjL6PLuxG8l6b5t2bSfzXs+jvr+8T04Hv
tBZslvfmvQlmLM34jsKgV3mEPEO+6VVcSsze+jPgOoKNsF+QNYeuhBJE4zRYd2yxCjgw+0X+Umsg
SBAeI2oGceeK/0oaaNacez1HOlGtahtRfj7pSuD74PNdS7FQMzqxiSG2FUzquVo9JMsB57GLcU6M
7YXN5IA6gzvTzJbibbBMSCT0EZV3ca9BmbrVVMCyi1flyX4nGDDfpz2L8E47UFokHa+8pwzrApCY
2yjn4yc91S6JM9otX3iZ6/Z/bNUYZqAfHtjiLVW5PLg420DIU+79uFkxygZUj3rbH/xdcKebcdGh
Dcr15pdDGTEGqjSeNN0TNRDcG5jvb+BX00L/IZqpdA7aMPVxE1G45IKRH+ZtO1MCoPMCNzhwrXJf
uzEQnlagqSjYNbv4KLN7KOIZ7hrRFwiCuqn9TSlkAHXokqOlVG7CJ2gGX9qJjGENDFzcYs7yH9FI
c8oCn7wvJiu2RICaFH+mHqZCOyTtzOWSBOFT3vG7QHkkofXMbzu20FcWMyUm/WK59j9uS2k47FRl
6/FRicnWfQczyYsIr1y9/kD3c0AYCKaQGqTC9IDjG7XdAt4HPAtczryWTIJeK+q0gN5ZW3DOXAuq
3kVRKpHXFv5YckyyywC+4cG20TnoUeDSGlL3Xubn7vryOKQ/1EPbVF3uuGDj5aArBeWZSPadU1vw
EcrjylzB62ljtLoKI/hHvecYENLMHpdeFIjM3nfDYD0vXElY222e+oQDKpDyj7/NQJdPM0lzZO4e
xSuiMPf2moq2Wu928KoSkhTXQ2c4gnbZJJRA5+/xTXoqfq/9DGAkkrwkD8stxsu8ZiZRh+rVvkNQ
UltEpFGF8ETN3wxNn6QZqxTFZxkTQPcVUB6LvMxv/8Ft9jTrdLABc7yy1ATHE4VDW8eRXXLsl1mk
gM5T033zvGypVKRq7nvV0aBYulhjATe+AmwjjpXocagCHU4nft8p9yIOs6p6iBElQYw3K/A1oids
eI/vnJ5az43d2583RTbwjKRoIf4CjXCaLhNLAlV/Ff94B89aTzvr96q0bh/4BKqZJRYsefhKpEQz
EOPN4dDqVOothstxd/MPDXG+R6Ms+5+AcjLtpD77oihueYjL/cknvffj3FOQqzQ3rTbIGN1xmBE+
zGCeLu07UfiUiOx989KuB0vQh/Kp6pa5vv9dtwtzgzSXYxtqyhFJXIrT/r1ngPwBXcGqyTormF7b
ytokGWP3saLrBjZ9YN6N46hNwCY4cfcT++GCNZnq14+fPWR2W37qHsZ/OZ1S6C7s0+5hCtnJXexh
S4+3GFKtI7CkGc26WKuJnLF9c3sMMPl8uhCUBFbcbTtcMCPgh3U4RqATvYlbkkpwLCvzFkLm/sr8
TTtZg2bhQU/I60YpxH4MZe+qMvVbA1QciixGVYy33LioDihTd7bxHXGO/WvDrzOBRKXDllKUxebH
rzKOcC55beBhUSUCSBr8IjsqDkafePIIiGui52yzQk22t0L8D6mfR9n+ofGXr1IUC9T34O6bxfIc
Jg89hen1AhzRBhtVCvE9KiL2ASRbvFHgza/Sv9T7A68SUIaT4lW1pJoGRKIoTsx+yLmD/DYThbQe
vo/tNJ9+04fvyl85hPZPbWee5mn5gKzgy7d3QfacJ7LJF2yI1AWVcKvZWEmDf3ambf3xLzysHyb8
SqSEQM7W78XjfnuejCJ+Nw/rs9Da+UFWza7NpCwR1O8VP5X93f1lZZgJcLzX07EMXbTwkUnAa5bI
Jnvq3/qckKd0ZpRA/M78wnoEDxyMnJgK6jSE/CFmBABIYJVaRwc+gpp6RnU8eV+sp2/DxnvvSphF
U4C30HRW9B/OYAuhQvw38ExjP+3Zg8/AByY/pEAw7FAyAHmlwGn+zRVj71YJ/YtQLj50Zhc82Bd9
uXD5oiNxRmc95Y18mcu3X6dahR3dMKM9Bb7xiMlKtE4x92e0SQqq7qMBoWTBHWlqrHE7WEAqjGqB
lu7xs2d22Gco1XC63J/i6QHPIEbCkejYbCUlcVNAnk+uiDMuq+X/UClhkPIm6PViWq4GWpaHRbJI
/frx8bZnyUBUhhq5PEdnJbiOWZdWl/uJC2UVLPa5JCaDTb/gd2IJMPJrwCr49amhZl+1CEljm8ME
Bd7YLH/4kvMSMWlLTtqrKEWuYlGj19E/or5GYVFhO0FuxIjzRLABHwHDp8QiJWQ+VvIFU9MTqaxD
zbdILqMiqr5ZHG1BvYCEywJpwGXap89bXhecAqeesDSU7h1sxzMRKihPGcQlPmwaE16JHXz43f9/
cP6phGMv5gWFMdvC7RnBlddFtDtNpiSyjlWQ3UGijJoyndjJoloWBzeAqoT0lHcrpa1/hohrXwmm
TXy3iZZjNrmiTBe785oPraweWq2H0UFmMR8Ls5akzAQrs8NZO4tzZzWE2BI1K+8VeSOQkNJTaR2O
GtaCpqHC6s7NepWXEEKVSHySdpNolrE1yrtdBgVie9jFXK/ejIRyBNlf1G9XJ8FW27yzKYMm0ASU
hX++XyA1jBTpM7PM4SBOyOagbPdjv4xtH3wIwCuXhBVucflMnwFMruXC+uo5WL5M/DU0fsYPRfNr
Twzswq8Q+pnayc+JIaI2GPCmvCbjm0x0s5Mh/Jtu+WoN6Z0anR321IpjRZJLhsuQ44xzSu/6uO3b
k+NtyjiedjbTIGLSg+MDsSO9//a1h04ANuvORJvb2LQ/iFT6ajYYlFpStQ/qs/jE58XGFGk3J1hk
4EgFQsd+jzEBArQkquVumk39XZYvFgukZTVXXT7uqrVsqNMH0aCd4q7yW2ocT+cDgDVI+WZDgGCc
jdx3+BUI/kld4S+IoGSuwm45AzVJWlmZW4rRiBjCAgLW7QmJTl8A4w5HTMScBCAY3m9/p2ckgKLr
iSbo/tSp0G+dXGvnRqpRa3JJQLT5BqVv98VRyBcg2bGyKonlhcAWz9Ihcz/cMcMCV7GSAxn6SQ3A
cejJX/38I0hNH6uH/xwMko8QqRx21PcRhgXpHVZ/9E1qOLxV5PVUC+dXnPNdieJpWBFROEd3+3QC
1C4xJpUAu0jdfpKoBLEVHWVgK4FU/4J7xYqzDQsEOGYsoujFqI/4KLz6r8sIqjpQgNeZD0O2KtBt
NkdROvZZJDTJyfk0bLkFiGAqUjlmanCr71BdCgTrDYujfookjWzACrLQdAxPcpE+6w6KO2vadSbY
s6TgOQ//Rk1hZK9jiNwLK9SGNAvpOyniI/y87fuV07xhhDT3DbBkA35vQ4PiAfVlCxyvLlkn2Rpl
CuK4Id1KnjeblhbUMvj4Y0BzuZgdsBjhJSonMMY4TY7nHQgx4dz04B9sMxVYg2Ywlkj+msS2OzLp
rg7MJrGUzA+QdUlAn3skjZ+AkPst4To/Kxk6/R4ymrQfrSqm083rXGVTbFusuCqs6Q40voFzsReU
Kyy4XLIkEHKRpck6dHzFiFCGGrgAmMbncV/DGvypQKJSxUtGJPFpDbAmmEB5PBdBTC5VFDUs68nW
MBQTFlCoCEJs7SLTeEv3kBPAXc6xLzrH8deoxBDV2UAC8c35obcNMr7tCJcPtPGXdWtWHbpr8gpd
duhjSH5ewDSR03BAi8De33D0TC13L2rvY0AWzov+3S9B3sf0ThdXrrh0KKUsEZ/4T1jcuQjqTwmD
v2yx9rY9sX3QCXRTpyCiED3pJHUIbGtOULK7sMBm51joXr+/SWR+UozW1UfgMBQBBMq93p3WdZOb
pVGrmxyAGCmwC0OgCRclAODzEmrfEAXpcQKLHFfvlll3+25YwAowrsPFY7dVbCt+MrG+wEe6d4U1
4fnw3SWfsOs0umCARU/WLgxke9JRTxs06W9H8VVRriNU1xqQuJtYWmnAn9hKrrWurj+CFlXd4Rxs
z5HZ+LvYe8Rul2BjyAHXBuBxPeR+U4YKcBVlJbrTGZLWHR0efcbUkzd6dQLEYHlKqKoJxHe4/VCP
Yl66A7TydYZ8p8WZOdO0/FMM0AMm3IWKlX5AZLamFNl2oh/7i3UB9om4+6aAqXvPR3u8aVhE9U/G
YwUvEz+FQD7CbSsCyiBZUrYbCZX0RkcKMseSSSctzC1LeNcinwlfSWUnDWjbpFhgy5FX4Si9iuNf
wMXDijSjJMzSziEMocgFFy0pGWv1xcy0o0ZpENQqmvIBIt391iwKLoIBsZyOKG8eTbbYpWcjGn4h
5Dt3aw8bBTOsyP+sWtIZT1ecVBjX288Sb5KDufa68COZoo6EX4d7d3RWlhFVsr4UGGV8r8j/401X
JRVBHAVn32SSXuhJlBYeTKvxCXygnhkiBSrj4ruHlyAMa6RYya8Pem0OvrdYjm0Pm0r+AR2/78XC
S1htQn+QKwPm9nHXlsY2iXa5tqTlrfKQxViBbUPptv76VsGCMiTCibmZ5PI4obrxjs6yC2z2/kzV
jx07xPGCFW+axnBgM9xOLMjdCJsKGIC/H+A8HIyc2sthGVboStwh86uAnvZIUlspEW5R0h5uUSUa
WzBOn2C4QACOmTaTTA7TfWjKNYJw/os3S7dPjVU8Pnv7uxrilvJG/oJbpOhOcfL5TfstIx1qRd80
SywZmotoZ7tkdArBhFJ6c/w4OHwig7PvXHMNe5ShOe3VIdbQiXWWKS/U7VuXL6W7uZqZlTX+ipUZ
XTsTDo93IoTcRgeByZLjlTYVYcJfONoMgiessz/eucaw/PkkIKLaGH0v4fqcOpHu3FUZ+is0G1ui
3gBXKP52aHo+68Cfo3LAunLBD896qaUJ94vwaGZDaZPdFLlsG6xN8cCxaivqjLdVlJIYITLLaFzq
wh9lh8kuxbxShBdpsEoBBodvtN40Jj8ow8D+BVMtPLH/gB5MENMh7g8FogWHZNZlBDRIgww9KbBk
ZwoVZxvaPDDEC7wod/rnlUsO+lQWsYlqq5nJfi+2MsgEPuO6k8QRv4reh9hWyuCzSB0h0SsUXtMU
5AEIGCESyRij9YMpVvYemZcaQraXnLoLnC0CbiSIXqX8aca9sLTojN8riYDPVID0ZRlLC9RC8g+5
RvVJUZK9pOf4HLFcwwmTdoOa6GOcPN24ijlWK7CveQ+WdE2/6Ic2wWRACXxlQEH4Zoj3wMdCWQNb
hTZE6KBxYXRYHnaJZh6L6hvVsoX6S9f3RzNTW+11KeIkdA4N0qRb8byx2w6Cl2ypMsErTfPTlaWB
NuksJFGShXojZ3ZD5LVtR3DF2+9rIpjaHHMLHcNHKZRhX/bQx9qldFsUCqPnY9xDEqUEneOO5Abs
7n0/S8kJJ97OHS0LoJQPxiwmaZ4sevPZ9H+Cub1XVExTyLmKB0iRpw08P9wNT9i7pXTDD0FsRf4u
OZDCei0ISTU7pzLVJ1lZb54b/M4/Bjt6lHN359fH4rAbEmlc9gSpWAzBs7uRLmQ0vo3hr0oHizeC
oQpSyqnesR7bieJbVNJOjj0MfjuqDMCJUUPXaebOmXgt0UZYZOAfxtINHhfCEVPvuRihh7aBtlE7
CEz+UGIsc1a5jipK15aWPilGeFKBE3ll2pWHEqbiecnmMF/OBQDRDimhJFplPmrobfMdcaSbhH1P
3XswbKyJxrrDULrTcnDdxUfei9Kwpe3qpuWi11X56UVlEs/MoMrY0H4EqpRIgjiA1uE3Gqwep4l/
BWTKGm0Kc8GtKg6cZrFqOKCdFDHk9QvCCdT0GI9+3ooFndN7H9dFOYF4SH/72IiB18XNwTHBmmR+
fNrjwft+71zb1xabeqZ1KrMZdlyF5V25wJN0oAyMBywSeb50bdjhDY9bUll0DyoK9tM7F0DhWbMC
kooeMCX5JMfX8uG3yfUBlxC4vf5U3+RkRxfHTF+J96VGQGEmOBBOTazXwIC3f+MXMdVPzE6vDE4+
NCCb06cpmznAK5fINjFYW+AbIGQOZ0gUAfvEoNWTRbvT6pBaS9qTVwfwH14m98hxpTYuqfawow8d
Ue0RCGFyRtlyazaR2BI927Bi8t6VFAtIUJUXv6k7+A1YJB82/tz5uBHGsbOHO3suKbjgaI7RLbrB
5+cOsOsTynx1lbCiZNvX3tH77fPk9VVIeVO8ikQo5WYMfwOZITE9bwGO5/fqDYtSLQOf74L2NGuJ
793jNi8JDuOZ5Vm8nT+SXSGTa3vT6aGG4LIwNL9A3BoTiVUdCL0ICrAAOR7J6dugRwBtFgwkmCUT
z89Kwu94zcEQUTBqJlAY0vMfotrq1u6N/3ZYSS6RftIHj7t6yMfexUgw5ZaWMliSlVdDi5nflC/O
XBdEIRI3aIv6rnH8pTzBgfcLxs+vj0t8/kfPhMFlMv1pfBErIZZIkk0d8rsb1X8HXhF/vPjStwl2
SEke9XIsMfALbrZmo3uVBaRe74nApNIF20JAwrxQX8dj3oIUKvpzYZiuvP/j07lUVzA1ZYAdoqfs
fHHY5837BHRoTjwCAVyUnMOENud5PuOwc+5sQHCRjixrP+kUpxw6p6bCvpQseiV7+HkFogR/duO0
B1X4oDpHow0963CUb/CWbnp25ZEzH3+eT+Cpa9fd85BsfBTzrP5hSbm4aObP/GLFDx3jG/uSf8cB
mi/g59tt/kvCH46hmEBAfeyvLYCr7BeaeBs8oBqI3k4M48tl4ss/3LXsX2DikigDB3JGIgsDJuXn
hXnTCkJq5w22dj6mrrhBB3k+mHV30oBHaPwGdGuEV+EvzhnmZpU5+1wT73rqec8wFZ9tlKRHJDwP
ILBmrOkydswcJ6VmZcbSlhwyfK+shdLEYEp0s84qimfyVH0WPMUZIPIhZ7hWh7jGrC/7HsQ8P1a0
h310W55txEQUS3k5gZUqjYVinbaxTrSWpWw0vtlsMySVyfzsg5apx99Vdk5rVizkZmRsvo1RKNTY
ymIRWe8FLHmIfDKYbY8PbyROXKAvSY1Gx3Zcm9sLwDpbVEZPwUkqv1sb8pE2ZW0AaUv1HltY6SeH
wADDtvpeE+KG8FWk+/NE2yCAPOokAvNbkEEPzrMpwjzd2BJfl/iwsBrigt8+to6mj8cNSsWNL+9h
PEtVp2I4mF1pYI/drleCJafeY9pf5C+2ReA51mOdUHs3OBkymlo6pud4S1APBBBoU05LMHFdEakY
8a1Cd/nBi1dFYiR7lXERYUpxFgYDGIxcl/j7gu9hX88YNnZrcRqNFbxmPAUN2VI0RDF8ZyvyDzB5
TpG1nS3P7eUXJUz5MdWje1zxFn+HZJRouC/Ou6J6oH3I09BYh7tAqQw1h5qkil83T7TooFH9jWCR
4Rmx8twWS/bJ2G19I4YbAH4OI+9u1GjLN/9w9NCPdsZWqBhds307UclvpfFWevKGFjUgJZaZGaGE
tcdKpS44zHbSzFcAOv7qDs7EjSh7qtfE1ahtpgbP1Gie0z69N9uVK8uIt7n45KL44DD7n6/wnzFv
6UopEPBmp7xFLdGwNyNp9n7F57iI+MRw6osQeBtTj07DRKBlIG59KnLudKg3t0Z5xr7RCO0Texqo
gALygJjuVX/Ar/8VREbl8etqzl/pRBlRQJq1R+uBoLVbSYQWMzSI+99WnbFZqWD0Ys7WBW7NGRz8
iqzqZ0mI0ImFJ3JFYa2u0/f6BDNjdF4sb3eKu1ihGM7/SFzaZpd503u8KXDac+Dv9toU10uGoJP1
8oaYHNs0dNpRJTuz2CqBeniv21ZD4VDeIAQ53yEKK/sVlPyr/v5BeS5juSJJ/r3TU9AHb/iw3Mwa
880tqqdPAmP7MlwiRbHGBLFpw+I/PLuQVQyFf8zVoqFK2EXzChue7RKSObeGtWh7wLi/84AjJau5
G3yFQ+q2Cw8qA3rkyjIYV4VFT5NyawgQUaSIpjgQyAzRmho+t+F3bxw9R8+qMdisaK+CiACLN3AN
2/NgkdhGg+zLmijjQC98ECvH7eiWEc4RCO/D2bmYlBzscvhSRg2QEFaUCaxSxgaM+fEWLnuOks3z
J3D6isYDc6+TFhW9mnqj7DKb7ZJbp0+dogAtY+Y6btYRTIxvOBdW9IJf1sBLSl8HcNx64kPknkMS
vhSdJ6ja9hTQ5wu2OHLd5BogI5RGUnAAjKnVDU5ceHk3uAGBVAc43DMvsgCPzzrp3mw659tlcwuD
5RIWfgwR/UwD5C6DGeNQgzTNcfiwUPnEUuctTlz7x+mpLNg6ErH5m5KQAtZwJ3PxDyXKy96kmht/
FK6S0uz3+8ddAlpuXcAExX98b3uSgXIcqUWk1GUyRWzckALzpoL7Cw4q/UbFLVThztpOjC+SzB+d
N3bs06IAfaaJcDtBsFMro7r5P3q50kBQcQPiiEvVU0E95LbWmEVmn28AvIXudSUbVTAAtGmGzqDX
4HoWeqMDvGq8DDHjRonZKw5xklJzJYBVhIpeB7JZNe01m7RhGMpJ+4D7TzGf7pGeVJ5QlY4KvWQO
/m+C+xJYm1mWWMwXAjppd3mwdKolx7G7i7wcamgvRT1pLlQYGth1Nc06zkLxY8zDkcABEvn+mpqv
rEwjpO421vo9x7NiPOzRWCn3GUXZS0xro/OO8OOImoJBug2AG07tF5Zl2ev861XQ3npB8l/prk6g
yAJ6Mwqr6gjIWgw5jz7eG+90QGJwwwNPLsW02wRbxA30beo04xnH3021xku2yy7C+M/5k8RirLQu
c70TBPNi1wr4HQJ15IVViXeDIcGlbY3pNJ22T/b5DODP2xGQKD3WxgOq8cwPgBu8INzgtwh6VhSa
DB6ATOyzl6La8mkZoFlD/c3rePAqkwdHRy1bUL7rq31w/07QkCCSTSrd6fi03muLRXo7yRaqffVu
aeVt8zZngA4L5bZxSdVqrrZeg9j1Tm9G3XeGFRRsCunAcV4qBN7dGqtOlJ3iYlyHvyYaG5U4Q27x
TsxQZ1EM/VuxoVc+3ET+aQtLiUgk5qlnzx77DFDeegZ97Q6qjGYRvta/8auG+RJxysn9rk+eQC86
4gCMLW8vDTwOmAbYi2z8NfZmGZS2Vz29ximVOzEbCWPa6Bib29v2caApBMndudP5T4Kt88uA7lhp
yLAQOT1uDGXWDV92Oke2sLUkfreYZyT+B59S2DUevoB9MeC0z9df1ZlEFQFOttcOPw4hLv2mFhRX
f2j2csBeFr2cr60osK2OUXbIa8xN0QT7tIB/tDh8KogXYeOg7lpR08/2rDmjWrIJc+4438BP1Pu3
ZqKyV78zN5koK43XRrGMxKKB2NkgG8HbBM3k+1vNzy6z6KNhYarxV2m6i7z/wTbxN5tK5W+WO3Xb
Qkqo/X9FFSEt2UOqEuFhtyB8ejSG0ZxIC2NnEK/cs9IZ3iBKQmfiEJF6Zy5FWM0Xe759XYUbbZkF
J7GA3e5bVdRfJiqcFycIbsA5DAgN6kCxN35+9tDLKFlYrwI3X7QaByWgg18Bz83mOIV3tVOyn+Py
dIwu6pv8JS0T1uTrLvKzuVCca11rvpADqG2netdi5BlUjbpo37WaIcITCwg4t94TRfos8p4LOkBD
De604Sj3xqdFYVY47eOIGmIIQ1TQ4jMzSrfYer+CVs2sBn9AmsT4RZaIsCyMNMNzkbKDbfoC2rB/
rFsqDUkG5hQBYhS0FK07yiU8bxxvvZvNeeUhaI5UhUcg+VyvdgD6d97Qtx5u9/D6GFzaeg5UMSLU
G1KteV2WkB4lf7muYXHiLAy2tISy2rBhCkkeUxTSSBtfJOUy2Gny4Oga+d7UVXrak0GVeYoQ9DbW
1jHvpTDJTIJ1OeTi+ZA8ltGagiYoUZr30KAC0ls14tUsI3C3yiMxKHCXIwV2PyK2sreuaIn1Ywel
Xc930kAfzHUAnZrP8r3vVkFH4yqPWuMJRt23MpbUkplMvR6mtlpi4ly5YRLNE+DkFC2jL9vfBrmc
NNq/CxyA9qoqXUjUgAcorICZnykwYApgj175IVppBEKiXv3WR7ouhB/iILSOYuRaQhXjvkhZgelP
op+MCpdBk+n6d5Ibz7M12NTAV7SL2dWR220vlmmnUeho5kTL/Jf28GjG6OGZiOQntc6BjAnscQ1U
HmZ8UMRMEOk7qJPCgeJCA5Hd9Iar0+LuJwYJQ4qAsXVsmgvP4viKoQ6hiD3+BM26Sku8EcKrSU4y
csXChB1pGogQ7Sw8TBUiZclVNKmHMa6lYjENald1D0uu43aJAUr28zESrSaAqs/X2g//pn+0x4kP
ZmMHAvyUQoKCAvFDOrpsQWdTSGO7USbSPOPckOGIA3xW+ogCG7SUrIXoaRw8gYMrTVhczfpXFhDe
zfCTZUYt+G5LaXLGn0khd2KrvflnhA8JKjuMCCX2pALRiEXeTq1tW4pX33Ai+uzX6GXwZffmsN4n
r3XbnU0Xq+wYpTMeXDMU9hKgkVuP8nAOBYj8dU5a5pGpmqGsBB2eF3BuYPWuXmLuL2K2v1/tMrEA
a5NJfqGXlrwlfJkky0gWLg07OSASoZv1xKxfhmu+vtqevC1iZyBjzuvFMi4v8KTue3Mj8WPzlkgI
Tg8cZM8ofrymFB4jyQLMkc8+WSyi9/oAXyqd6O8hdekaGMOFqvFcF+yK3eUHzJqoASRKvMM5boOG
QHMfP7PcHqRYIQhGGNTxMcPVYkKLtCT1Y/NFNOXZs6+NQsIEQTOzQ98mTUTRE62XrAzM6Loa1PCt
gK60CftugK3gjG0JTAoo4nkGhyjdfa0QOLtorICMrshBl4ZDWyzZ0ExVvXZ8iEmEWj/kRb667DZ8
luYb8EMBkhKe/Tp87IvRc0jDBohCYzbCj00N5uwZ85bX5RNa1EfJRUeP7pLmHhoNO/SAs2QnEYhx
BqN5OJ1P8uT0PGrzBNZSJ9mZG9okJLKzfLQToZY84Yo6A+zDzwQWxT0ql1+x9c8O2nFpoUIjJcI4
0tsQc2ETRrVaovQOEYB4nEfEzHOjwFf+cZhGU+OJS3e+JTDrOKDhPI8Zg6kayj3HdbCnaalK2ucN
DdE1578T7TjC2nOJpXFUJhRAj63hR1CoT2sYZYjFx5fiWnBeR0wlC6Df56Z4xpUs1P+bSf1+cLJe
D+q0hNOfc9AQVX7qX+MhgR96aQEgDbRU/UKamNC1q+kIuBcDF/uRFylI52z6eABCeXyPu2FJbdom
AMsfFOLXmQ/9IH6izq5jTlXCT/MiHUpE5hZXsqFo2z/q1KnWhlqcaYLgeVWmhK/zryT1PIRMIVvp
diuGJCzLo75jLRrzMZSKb/PrAOPGYmuCGL+Q2ybucb53CWk9ILPnvniuUGA//GO8HZO+91Y7rjlR
8tSCJ18Mqbc2KnGOsbmKt/1faeHvce+eUjkK2CpuyU+rz6YP940FyTi073y70Mk8iVPDieBg9Bpq
6RQKGwXF0Gcxj1wpos2tmSXmRfy+DJGpwEFFU8PxTcAsm18aCkQYw07ctj/dvaCLMoiwB1jjA3qZ
9Pdjr0KobF+/dkUs+iMJmCKIRacPPBrmZ/hc/omBrQMAdfdtmB+tsTSCCYOkQ6aJj5XLNMuUh/jD
wW8CQe5avDxmdW1g7dzQ/wNNvcG7Y6XWafpLxbO4LYSJOC74X+mK3D2TpSLlOswkMzsQvdP4DSxB
5w6schQ+C66qBuQakXZvVrXdm33fqTfWL7GzSHepxa0pLxTebj13T0NRdwSyouQrpRo9JhQgE7Oi
RP8jvK9Cg3SUlt1VPtb/5AzQclKwigyvWcTqehNLeHrl6KQBTp1JPXF/wnIUOBtz5e2gYa3l2UFB
G821JaTUGa1WzCGjSK/QSNlBXw1U/cM03xRBsCLLjGq6dNN9F3GO6YAKiZEczjnSPucA+A3tXClP
NTVUh8U8xBCuTLscawWDaqCrwLqVgvUJm5aZwg5k+J5mjLXkpPKVZr4GgavRfJBQ0aEr8vs0bJdL
l0/Ne8PlUZyhxHlIXWdJ6h/8Yx/6oeCzBpyz+wonqrNvV/cz2KX1JhkdhOmSSTyBQky3va3iiIDP
frPn8S9lMcE8COw43rgpFUqA3KlG6z/cDrWWkSnvIKpQSs3hRhK5IosJ2aTWR8JxBtnVJzEKC8yl
7REoHNjCWFfBkQPmutY2BvzmKsPVNwPY4Lyo/d01uWVOP5NJ7IOZdAQ5a0AVhirJRTiyZquLBXaE
kf096bBh7HXXRqmVyn8lPYTMY3aFmOY+pcObfHm0FY6KCjNhSaKZo9N5JyMd97+rCel2EyQwmb+n
UbJ4lOwwb05er38CVCK/cKjSs5mPvxmipd8fZTP+sD0sRL91bpnItj/+kyWG8sxu53byDI+Htmar
cJkGamsSv/W/7jryE/mItGDF9pAP8Vt5hjOvhc4WX3rauVmpPANJu00Tyfume0Bcfbo1geZWLZ0X
AYEm+2EEVCrjB7eGp8dO7x7Y+EiTQEDuJ6zzT0XURCE2v1z7c60c+mpSQiFGQMCKZhAq2a9t0O7z
5T7o7z0SxzeUiSEhxFyKGN+M9a6mxaqBzZdkGnGIND1VXC4qTfrp3jcZs1Gt7qByB6U/s68+3qQB
3cFItNCoKRK60wLpeo+yeportXIyzOA7j4ZY7qTGXJlIu0KUH/yDLBzAb3Xugf9XBz1mFIAQgc3k
VsUL5YLbhImRgVLdlurggLI3Ad6NPh4Si0rt+98puSZ8qu0qRkRRgKgxehX+VZJ8vMaUofYRZy/3
jNX/8J1ZZERNhpMQVLr9nm4UoPKgGK623yZhDGfu2cpDZimXmr7qHrwxzeA0W7Go4cmvGLN7PMPb
ghKfRM0t83Hz6nQVpKaTZqBiaGjJRdTzIQnW3Q+ZAq2K9qyXrzIEa+Dwgh9Fp3Ge2ARa2y3sNPm4
80ANWN18C1iaf2l92Iq35rbku9yInmjVzb0tHeTZIMaTeL8OHA7VFigT1oqilxihXL5HXoMXgZqi
mQhMO/PzjPUp6UP9Q1QZr7q83dHmIuqaNdelpBuzdX2gqPqlbF9AYxRFMV7jK/pi9ZSa9Kejvaom
5MYieUZqps92QVinaNeUM+f36HS3+mD130yxYfYq90pmtpoU1b2XKDX/CxaGmqv+GpDwq7GgrpD8
cFpAQy+8Rxl0ynsqvkjJcpS2GQHpSIocl98GIqBGdKFGmxMXmGyUnIXkA6EwyqSxq+aAcoPDZOiu
9M9DK/50zxH1DP68r/KrSGWwk23GQioPLRGtU7N4fwKdIThuyerw1ngI57CPRYFQ6HZvVXG0AwNU
oQqWdjOF9osCTL0L6rikV33oFSYBAKNKUPAtSa0ThUGhCT3qW+W4bVz9vt2M+cA7VV/pzn9adEDU
osWWM3m8D8GvICNcSEvRG2yJmHDXJy55DeoB/vE4qiAQCAbopBjGppZgnugsOOsCkJHgoL7z4jUQ
uYrDixWdcb6mTqhx/Vexbdj50Cog1/Qd2N8Z64FpHkXL1yv8mcRp6DegSaW4l6IJCkcGq4iX+1r0
J2I2kvLUxol6ufs3aQQ0kPn16BsRBin2ZfH6QkjWtt6q+pz+GiMQ5Bcf/bHKZ9NpVt1IXv95p0o9
FMpu5W8kwygiU1bawmloVGwrjvicp2Isu8X0G0FNJDebVk6xK/zELHrhNg7p+EEPL9xRk6+y/LZk
YsBTi9iFPOMmHzWe3eehpb7tXj+zBk9F4Zo0+vA2XLOXkuZ4DK7ASND4LZpuowVkJ6ahmNaBdCoe
b6+X1sJULmQr6Dq7qZ1oPzq62JEFu/PMoW7YQ904xu5xXd6dRMwXr7X7EP/CrasfU7ImHcY+Lsqn
EZeGOsGU4+HhAV0dmHrStE1rAw0HpB5c9d67Rpp1tYxURhdqikDyvfZzOoRxce3b8Hge44hSyE3Z
fh990OJ/VCg0hJRGD+NF0+WG8KUTwtbA4sVqztm4m94iZ8v6ujIeUSU/yFAc5QUR7qzfO5JALyy4
ZS2PtKzh3Iw2j2WH9mj4HJ5kU6BsDO9F68Z4FbMuz82nV1fZ7u28W13LrGwT1Ot4GTRfkzBOcwy4
gHi2qtqpfg2sby25wbUE8Y/YZvsbfeOsQDP0MC1Mp59Y2AXgQueZaHNvyRHspn9ApVozNbcp7TYw
ohETlzSqUlqDnr7+Z3niGwuXfdetUn6Wp1SVilRydLNU1N92grD1tX7BDtZalAo4vl6EYtbyV2iT
oZ2JfeymIfFyvrbn1wsu+E0utrojVs9cYHi14m9LhyqjTBVMKsDpDpxCbaYqQQNTyLZHviiWnAZi
t81lz+2aFiwU2al3pDDKeTeAhBWXsY6/u0xKrHOPtsis44N5VWg6L9xBvgzmjSkkOGAQCccReHwo
YPhzDEyahSkMVob9MswTWwxoAI+/98D3tjDkwdNkrOVUaiMf14re2PaxrNnyNlpXXstoNNQA0asv
FTE8RI5Jay9ITrvJjC8T48DvLHKySN9ExpeBEK+uZtanQEsi0616r43WgW1NOrzj2KJ28fAjFO1B
VD5sMdVNUE5SvVvrLWfqxtIcjiT3JnJGlKvnjHxdHG4At3zT1jl+0PZssJxYKetw5yeEWeLoLOaF
II1wh5C260kLX6dud9Tp2kPlhPAoI677A7PUHg3X+4MZNZExfgUkaisTivo6EZxgfTyGewnzyyeJ
DkhwKsAO4iuhUQy2NgHIVO2pgdqJrjrIJM+9p19mruv+pVph6H3gknhPphWaecXCetWaiphdl4ID
Z7Vb4zAPQl3KaR43320s1MZ1cDllZ6AmQ000dOq0H2d/6SOy4xw+xx4GEUdCXwRFWaxT5BqtDt8s
BZpNoiYElwsEfruH+MhH+MTsR+ZOoN2qCUveol3PpsijgwYubuAgH8xod9lIMEdvDUOmEIssYaov
RrBaqu2cVI3u8PWzmG81x5caOCOxJieCx7MlVf0MnCxUeAhdzev+qnjZiSroPI8l/aJsa/dcdoUW
6s4qNobA+AMgNffz5veJrCo9alDeNLJgM5mYCGO70571x9K8nxCmakDU4eXboNtuzYlL2aCplpwP
UsLp9bot6H9O+iV7wO1G77lJGOgMLsy1e/imIaqWCA2cAOjTHsptaAm0Da/5GEl8b/tR13yk1uR7
TvKbagaXd4L6uQW4c2snkSPGRLGe/7EmcaK0FhlqfI+Je2Oip7D8n8aoFcQXD67XxC1V3PvCT0Xk
WAjuN48akjDUt40yG3aLV7TTYHAXmkwGthFU1xIzfZVnkib5ha/16+Z3g8Gl6lJD5zGc6MFnrVAR
7/n7mTo0v+fDSa6zRBugihpU15sUrku5BB56rposNZmzoR8BlnwdhMDWsxBTxKijmz5tbznW7Ye6
YqxjSAer/TK26EnjpyAw1v2+TSXW00L+gKVPIINyvXvPzgo+IRwz1TmiRh47avnUcuWlHbjIdd7/
ALdzACXLQNhlmMxdb8yN+SJyUF5hSxue3FE+yZNj5vRT642NabtEZMdTIBcH9ATHnmYwATYiG/V+
p2diYDjE1XM/FKGcXLUaXcRZizKIG1zH1o9c32fbVYes/kDki3Qvat9I57TLWjxfzSM1CLefWXyq
obZQB3/IrbijwjHFHHk+hQOYIkPaRsIfNUN9zpdKvRwpWeMTq88KhBzzPd/Kc0RFygvooI0fOBn0
ctlngdSEnZjcuZZvxmo76vsON82WvM/LHviFg36eENqnMPhfz0TVx18qskQ4yQrkG018wGq+srLG
dsdXkMazJDceL2abwKSnt1qwVqD5VZOcA/m1aVoA5Z0C/+DkmrPXlkjWueeOUMapQLHLmg93WN02
Qqct4+SvgpBlmpgFoWo+VOnhmUNnIIulwuQXqFUf2eCH/geWfNrgtVSHWfQNAVSGd8pjAW6hGlot
c1XABoYC1iYaBu/fmaRu/P9LICFaELGWP+NLv22qgbAEcJCM7RNl2lKODzql600ptt5zB8qjmY6j
EmEFBwJGu0GBlSqjjGEAnf7bjMPPJCfwiUdutdpNY9mNXzgff3ELg3EsYktAsJgmP/Qa4vM87OXz
GZ2/kHfZuivmVo/V1Md1eGgWlFTf4R4Dx6yK+xsE7pHlbaRYsyfO2lSp6zJX56QojKoPPponBtZW
TGvcIM7kvbRdUOecOK8cTHKtr4m3wDKdomgshD6B8Dkxy+GWq2JCxYfE0eTY1Tcn2ZVO9UZjD9bH
G/sNi826Zv+yAzplwYyJXqCsleQvP8i7pbyQZWFcEcMz33vurpyOjnLhOULnjLxJ1/ffPPrvrwsc
wge2+XTM+qnP1n2sZm046Bj2U3+g8diZnsOgbdjDtsXbtPrKCDHZw/GQInv7u+eKYwQXpOhKaWGu
v5xQW8NEtyLje9rvyqZ4C9m8p8ut4hfyT6VeJ9g/1lRRYWiQEpRHB07rOiBYNaY+jjXYLuZQGZJy
MHudYU/x1tkOt+ehilWzkIAdXEVgj/0JLwGvU9nd6NRr+66UYQzn4XiMlxVDg2pfvaFkOBX6aVPM
iB9jLd2N9oYm+C/fLaWnbhb+9WPKLK+K5tBKrroQP457jyuSILSHQA22GG3NP7W1MuUq4yCtm6Vj
VxIFF4gKohMfEJwz9IYrIby6I3z5KLJZpdKxprTPsPOf6YS0PWBK+7sCCrK5M9GWyOWrJ1Qa2Z3D
Xo8P0IzjOLvjEXlxRiPmQL82yk3K0UDwjamlfcW8asunxYjwQ3SKVyMhPhO8yOW4szliPVW3/dIX
W/2PxSik1U9aarthqXZc4rj9U5ZUredrbs+kwGvhOvAXbICtVjDY1c/4IvfhE9UdBB6Pu20dqNyl
LabG07dF4ITXvf9e/Dfov1Nn2HXR/Fqn8YBuJJxC9+o9I6UbTXUsso4Ksn4PgG5fjyB3xlqdq4Of
CfImIMHOkmQvy1o049JRTho+QdBSAUyDPkX9g1ew69z6PUt7IVk+1qwtGKONBu0Q5Fcbzqi4GdxA
qpUMSbPmq78kR9d9ukN9QTBpu8Q0+vjSjdrmVHdy0+6zFOzmlyyLDHrbA1WWRyb1YnZSdVWOGG4E
a/DPLe6wpbO8VVO3h7MCd+pPHJXnHQoLM5RtSETtXD2W+bJJilx+8ulg3PlSJMYM6yr8RD1md9gX
1QZrMK8pilXT4WlSw8eO4y5nm6w8BCWARKlKVhVuwxXuD4WC5b85BYykKcye9muqKyiIAGhZEK0w
JK3GQGd4DPrqSTtugdjaHaSoar8JfS6HWzSKFjwS+QW6unEBzO/TdsVoyxMlN/iibX406Veq1aLu
AagRRHiBj2SK23LFUwsIKkOSf+NVWBAe/q4D/rtM5d6xonQeWorWLFF+Oufcwq+MNtm4dPmSz+tz
O8q63w/R4A8JgTAO/+DX6jAE/12rsC/tC5hWrzfpZYq11xOL1yKxz221ngg0HHbBphgYlFQk5O5d
X5Mz/WwxpYq6HPpzAuxBxcUszvkyLn1/Sn2Sr5EiDrqUdYA/pJw1Wc3mZzxMcTBTCsSMqSADq+sT
vPqt5vDX27oDeTH3q3PuJCoYqEheUz0v1EJS/1Kn/M7BMSyFeJY2mVP97sGNddm5r5P2eLI92o53
n4VPlQEvVpxppW1vsJORbzxID8senI/h3OroAcbIXZNArDsKbjTrlxgCOWD8hREVayDqIt6wpRqI
1UXjpQDCOicFMdxmyFTb49VuxOZoH9gOh1Qcy+MSa9KI84vkPjx8eqWohm9AhgW/HrMZRt71oBdj
RINFYWlEcpE9ov0cWt0ckTecYu+ZfGpi3c/J5GK/iUbKaxZhIfZj1b1fPwdcfnq42L86QtSIR7/H
Hdp6z4k8v1bmm14l+Jgmfzb55t8hhXc2GPditvRQUv+2Ngri4koB3BtGdtp+q6Qs0NOx36wzV12E
eK3EbMB6o3vE8PYIpemIkdVZjFryrkXtlZGaQGFZIbip+gzI7ZmJWFm672ovHIN3Cgn4ppllx7c0
V330bnFgAXBuwzJCyME9AZsDrAA+70AnlyR8KKMQ/y9N3L5qyK1QoiYoK6ANTI23JeNKiabFGdyT
nYZFxty/0BfWkSSkmEe7yOjO5iI/rsyKCUmxj5ep47HKYYJ4ESk4ctN/B2wbYFJzSLa773F72pbm
9HyWOjeIlcljesZy7coHTeVu+nhp2G0yQlUOygbDy3k+Ea/Ka4R+eHorOWJTYwKE7uZ514kzj/b3
7Ky2nptlMcy5qhs3jxW4DhgGl1e2aaoeI8y0DFbERO8zHLyUCdYQRmDd2NSYyQQ2dwjaHhrvVr7m
MH8ptt5iPbxClUBJRAZcYWFUdOzGsLSX2iX01vSskoH5/HoMRPuKC9R5cetUvWnPonBxb1FYzVCi
yjVcRFlrXxyg4GcQtl+G0iYQIe1Q211f0I9Hmq6JatOhyGZjKvDlMzTVpR5+rR1ow1oT4+k7ux7D
u7sbmx1/nFr0DSVLhfOHyW5LrvdGA+YIdFAVx6TnWT0EEzPHPRaVtd/9BkMi3mpkTSnZ/E/T/JIV
ObaA/fUjZd0pYfsy4BnGqNKnB/UiIyKAaMPpG6IcnVAexD2okdOEDxxXbex/D/1IillZ3l8u06dZ
7t3kyQcvVZ6YE5f9opXhEJPYBVLr0xtyx4Tgq+IfaAdgVYHUy2UeTNRXdGKSnNoaFCOkDXQ5pyBT
qr1OOaphyVc5b9M0QWoYx+aDVcOUmO2rtklES+HrMxRLmTOsrKItPI6DlAOjvNrPa2n4WtpW4fS+
F9ExPrcxU+TDSRSytT/BAzSBnz+WZAVI0g+2RWPRCuYJFuYyNwL2em0V5Rxbyh585q1fQ9UBCm1h
H3fLavAcb2FG+YhIYVytU74ngeOYaiQPdU8zibvsWr2GH57ElPbLqhif49SKViPD+kQMBiweTK8h
X8BocLIQKMte85P8CfPXqdoTiw3lms39yQCE0BtKizgZlHjYGi+0qJqSn+StiM6uS/RnJKQfkjYv
xH3GHMLY9eWEovvsqOIirjLZpPhFnKfQ4WQpYx3HYfuLbpwcuBq+08WNaz5IOMO5Zcdg6R5GLtWh
rmHq141OiqT6Ioc6/PFf88t7hZLDzXpal9BDHYN4sBCr5iH94hKzD+23hFKK1yveUexgfljhOGHD
oYM3y3ghdDfknzQum7GiS36GBxfHqYj00e9bG0Lb0lxRiYwtjSm651koRq5Q4KzHG5yFSnCZrdmq
0mzhh5wVpxf0bNnM2Jgssm2vBMkCsjlFBwd/dlkFOC2rumIe/qYk5XpjjkqGzwpK2HQhNXfUejSD
i+kt7ekQLh3ejEYa8Ip0aPRaZHPDRd8d4UR1oTLAIcIb57A0cmrFoefvVOdDE21pJ2XGyGPA696E
tNGHd02XlyzCCOVF35YzRVM3a/qPSUKYbkCs+5SlmcDdxYf3i1qQQNQRhiXgQrJp+0PEcOFNxaen
3buBsNFAD3dLspkLBxepSiFDzftvAsDAOqVO7I9foGUvpip0ZruGBpBhRtCXEy+HRT7eE69D5c5G
J0WiC2c4FUAx8lgdPtWS2UL4sYs8YxP3ckTn5pt+L++/x0dtzgvETJVeLEf9bgYZZJndUfeBPyvP
ZFJ5dKIbrQmbeKivqQkvvpw4XeSWBBugiMZgKcUZ/KglbRh2xWtzrQr+ljn+s6z6vHmCXkWBCO6d
e5Ah3sRAjGNtqTYntSO2++23Kg/1bgdMFn0pezJOJy8OKWTk0ECXmTXw8WTp8qSsd9PWbN/SrffW
XOnE0xXlQKJYTc6QMcPuHCIHE1GS7jcn0ggEeSdwQow9JAP3f/yYOi1cgVIgTx1jYP2Jd81G0ASs
L+JSDET3zjL7il/SVgtMCzI944zIT1ge1EnAFIGfh0LA78uCw90sFZBk4+U4DUU86P3DRQBwvftr
1AaBe7PHyUPulvf25vZ/ac41EZxaq9CSoUA4JuSPT4Sqk7BOrL+iohRJuoj7N1kxOm8b2eYiX46u
uTdws+U+rpZ5+C+km8roQrK8oX/EAV0ymmB2C9ZZewGSSOwkRQFGmp0x902AEQI9OeBV19wRSSze
bcdJDvG4a2152BPabBb2PpP7xJk5dnNsKX/Ileqnh6nkpGqc5479X51lZpsdD29AfdTa290qJPMH
MT9gYb2nViNFoHIfrPfeTtqK2liJxR3K3Wnw9XWDb6tEDiCOWS78ZgSJaBOcX35nYF2zrjUgUjsK
y3ctD9tjKFaME7fBla/AtRIpv9DCVF0MTJFPCkiR2uvMjvqCnO3H1qBqaoQSyjnx3x6YKGwUmvR6
FmJf4Rkatmnt/ND+9ntvGkKi7VqP5EYp++6zFl1aOk+R4WubgZUimio3eYszCnTz82IfNByoP2nY
M6wshbiqwRcgZRnvZrtmpcENpyN75pj3vSxAP3QwzVPVrLeCp/ObShoe8F7Zw8odwC1vl5nyqPVy
tJTmXo1qEKPdY4P5IPNcP/Fxa8M4cKasDPHXp4dNcA6ZuoDVAuTOie8M1T+GqiCqMVcUUF3LRF7H
v0B7yFIMqJTZdJGDIx9iYPzPeqZHdl+qqgIgpvoAULoPmc80dieOQFqY1M7JEiWbtEr9DVP74Iw2
/wl9rkIqra0tA+wNJ3ykpLEtqBo2GtnyYFbo0iGc20yhCSTjpK/1GSgtb3qnCICO7d2uKJAdTOQ1
EmppZKqhCIxuS7tpqVSBsn8XizvQ2+ehPy1cil80WmVfr8/rCqtBnmL/8uL9v50rgDu/7mcZi4ZL
vDVRLw7t98JConmi5DqQpRUonuflA+ZdyIm2VijOLdHoS2cy8/dBReyF4vm14sp+FvYtlK0ZJET0
tiWM1WXAvyNJ3mMpvboeelip6LJ4HXRSfLiIGT1GZc9EW6V8Ox/c7k4pn3naNcsnMsipZkhLnonC
EiCPe3ViHHLi8TR59GI5CsO8bUy7FzFF7M1nkKAJoxeSrb/yTVdusa+HtJwfIF6CY+2nOMLYT8TI
MErr/jkA8gQBWCCIE14ktwSRgxFuEfhs0lH0rvYUEO2MG4blpXdPKnz2dbZvCiHQrkF7gozyNWQ/
8eXtZ0VayGBkqE7Hm6VoihIeAgiv6sJZvxqtV3LWFzY2YVWWPRa7aLe7LMK+hSG9R+j/bj+shXnC
EStOvPVX4WC4TkixVEM7Rb87pQIu4BkThFyDL1XSqC9rqAuwhUo1uCS9RwqWFudnlhJkJsSD7ZLz
Vjrok+6aAuJ00gVsQpj/vnzfuA2v7bc1PiLMHPlMq5Ok8AYITGMdSM2dYkBLMCD9JrP3zqsueSAz
JO8FMeTqGJxOBb+ASvvAUv7d/eFSuBirlU09HWHXHbzCpSmEXWriQHlL7TfqVx3Z+ZgOoxiTBfcR
4ChIu2ZbuH1Nf6YVJ/v2TAyop4vRyU19rC9Kf9mdLkryPW+E9gfpvYAnU32kxYdPPI42T1DLc5QY
fow/IJTZNIjE2vlNYYiiOeIdTXd7K9+tniJhgTzIIO1hbnEAaYDcuFRXbI6bU+b4d/7psTO8/X2t
M3vBVvb8OBSDib7e+xfFvtPueuAGyz4F60Pe6YT17Gp5Qa0Vn7qd6/aRr781Q0EtDptgJb/NvXzF
e+dfHtQLYtsUM0lkSX5EUP2MbS4V6OyyXvkguA7Ko2wpEIMs676ALjmwwINqxPqQDLWE6IpgQkJe
EuJ+pEtPQQBdm+O82JCL8nJc5t8pR16iPfcXWQEArQZHD20GjrhWZO02nxKNuzsiBY+Z3ldKGLsy
LmVt6VhAc55/cVwazAT095GzVKbIbLfRPB/FNKkdNfQiTXA4q9tMurPe+u3sP466jo0010YBsk5m
eL5mLBklUjV1CjPAKbdHyyzFdJzJKXxAZAS3fiYEx3Y4vdOs0WAN6JfJSvpULGCAGvuBENraahDH
7PMcRLXPRQts6WJeuCslRkfoI07Kd8ZLrcIFkN8PcjVHNbPODLPWS9e0UCwM25ofZG20OK39Gqlw
jePWOvM/Ip7FLUivD2uBxgIEy1ueUtF+ZZyP6xrH5Lw+Mcfa+fQDcMTJtFvoeEmVn225cZz44b9M
m6iXQqdNGlcVgJT5AP8/mjiqS+6AEoqajNm5ycgULvfx69dGm7B1egLwpw0Ni78+PlaTiCbwkip0
MAPiLCtNZ48h/z5gy1edr+UsZlJj77xps5Dehs6JhzbFFE4uqY0C3ypW7yzUL8TWxoqqDRRcooc8
r1PXs9LijfyUSrjVj5/ngu1SOb03PKFclKePLYgYjTlMdOSgf4jTlYgPXr2UnQhYj9FCExaP18ih
nEKHphTtUnum7VZOgWw95H4ivToTrnI/0zQyYv+PJFX6PsuL+kou68AURvUe5CcdEhPyuHpdcS7c
9LlL8wFFyq3tyIjPobb4VGf3bhfpbDKN1tlcrN9gEA7EQoVyaNjJsQcb+r4E3VgQ98B8YwR+B1Q8
8kcaYqQr5uTp+zwHLtTu0Ou3P7ZasQExwFokkDbX91FQtfsf95qdia5h9dsV9VBfu2dmR+8v+cbq
kSbb5lNau/9LweGH/95aaDy0lc11CuPAlMRrReNUVF6z2Taa3R/oKDFiJt8tOZLk8bVaJAcqBZ/h
wahtfXMBU9/TkfdSlJvXLJLNWbOXMOZeWVSQp8a/lb311VMHg4JK8mkF7dwQdBlPuFSqWJ9KyY3Y
tY7fHJpNnmdIIvPh4nkC+tUpWuDLVxr6LIny2tsFKg8MTJtG/NR2dKjwd8jZ4dCc2rf5jqHYwBNU
GTJfoQI1IK2jcxEJV4ROXhkyA3Q2bF/QRubr3vkMn5ut8PxBVPt57pSPPZyaf9vHLgiht76bw+cD
U53IhYeFpj1+JNZ9tj9/V7aZrwK85CzdXuwL6eVBX+0COfB88695fzVcxVIcZ6WcnFUtDpJu/9ge
vRnKV9dpx7HQZ4nbkRnWoEEn+YZD0/qWYI/qQM2t4ZPHIZ6etEqmonobddKFvB8TwyEErN/+muVs
DnhhEmphcrGvywNWxkilEQ5LXN4t58xfwkWLXZpa3AhmkQmFjZORCeTrOeT6bbGXBARhuC+7200t
t1kYUHXpohpenNy/bl+wMOoRmHl2rF/9fxcIDE+OTpmrHw2Pa0jKKDaWMjJ1If05dG6fcO7Bubmo
IJN+0LjJwFLaxN/jzDHbxv9FQvXcIK3l/Qg6MFj0qthJyesXQWRGApzoqEh6TrwYo3shwRCg5Wr+
srzh9M+onzr4gXnHu0tkV4ifxV3HxpYHFfkQit4af4Kk2yj2NNzG61Nn9bPI1JEISp+2oijZBZT/
lOwbXXL9EzSJfbBeDu1JHgcNL6PkUr46u8yHs8b96yjpmMKs559OIyXCmuQMGFqjvSKl0Qt5pEj3
wxLc1R5uCwXB0wYnHeHrxEX0wxB4hOvPxroBRlvAVeBQsbY39rzUWWeJcLneOleyS/feOXF4SRF8
MZ+olVmO9c+wMw1Z33itOyFepuMR4sJjAVjKx0FjxMEGnsDLVh5k/B4PxqhfggGMKq9jWrWugso5
LS1jkfoEXe0Ml1ltOANuk173SrXjNHkkgQlrVdTwCk5VJl8E20CqooOyZv54H0izBE/HRjWaKEoy
WPQ6moOueOI1amF4jsizgz6i7Tauo4WPdwxjBzdFQSHphE9fPXCkoK/6qhkVUkNw1J5akb26Qhod
oA6JEFBLIQ2kxhKK9AnJ2AVIpaTEVwua4pR3qH9UoX+mF2KwiM5zbllGLbjejywue8rjR4fk3tZt
uSxXRo/USeP9Y9Aq0UqgSDfGnG58+TnYoUeiJ0N50qZOn66w4tV6YfqNJ9+h4adQFm2MWvhbsrkT
BdKMIB0wpmZw7cl6E9Cc5guqPXumKB4OC1ReS2vO9uN6uzMUWtC4ce3ixZMFWG1vX4TcDYYp1KBN
/Tc2SG+lnyjqaZA0yZdOpL9BngUIX949364IY4OqzepmjP9s1su3OPMhtfsRFIb3MWcyRrA0PBWg
s3g3P1/xAjXaRrcyt1YNlWKGbf5vRR8WuP4dUJPGerI6wMBJyugLtUPWqDWFGxXxlLqla6OI6Lf2
gYnnPRmGWSfrYIApHh9d8davHYX0IQxaimJLfQYZn8aIVwpG41wVaNQ6dYeTg8PLboWzV0VV1TZL
3TIP5UQDCNj4wTjQW/qwAvfqwHTBUdnd24BOnhwnSd50ukQGYhcXBSJHSqK/2OJH5hiaj6b5UjNJ
aCtjzKyC8v0uqsnkvJfj50D1ygfhZd3P5puyPXTwi4v7L7hbCRUdYI3dRbbIyaIBcqH0GtlmniyS
unA38YelmZJESf/42847rqRcBltX7ybkxPAM6D7tDumChse45mp74YkbPsUGY05xoXWaIZiJQ8Vn
DqL++WSbMWqMhf22dsBddBCd63PH3HRTzrFoej7z0E9FM8ZvSnkfZ3rBY/4aHmvf6eRSgqPrcoqi
KdAV5eMiZ5m9L1N634KnmXvbB7Ca1+D1lCl6j9tIM9NayajAGuda6tjmMytAIep2TRynwbdKPbnj
uK233BGAEhPvW3nX/Gehb0en2XTTlBCrbj4WNSA89mU424vElfwpC9cg4ZItFtNfUDhVjVcUJSEg
BDGYwZLG53AL44R7/T38J+Yz9+feNg/DwUKCu7K8g1u2+5DqtTsti2Wcs3vWFv7cysIiUoXbt8nj
Asn3nyaKZMa5PGUbo5w0R7yZPOJxGkKIe+PHW30BFvpPwt1K8VjMGf0WCoobokkhYUU91TFJaPMC
UIDYGFTQ7BSDEtfywSNeJATACzRXxhclaNkyzKwFrrEZjYPYLx17PhXdVMg/pNI/bfueJ75/J4IZ
Y1kHqajpCErJW0xQA8gjZyC7b03HfLFDz21ikWub0na8xhMnCaYT+ichbz3aMrpT70W7ycbrfAoi
Ylof5ToAtognt1DSvjh7PKGRIrbRzKxwhJH2o4fc0vU/loo3HiOsh7lqPFULvJDXcr1VAsBWOUkp
5M37ISw9URIYMOa2ooH38UCwFwFN2jI5PNoBJU5TTJbLV4Ko/7/87mDGkFeUExI9TJUwDkd80JBh
G/sdgEzWGvrbTVFjslo0wH8YVjQQd6wg/PDXE5qnwXR6JS45lZnQe0/vvBVaDVHYvWfGlsk3kk9A
CDmuElJ7mbCf99rHIZa6FE3Jry3QWKIFsryWCGb7ieJy/h+4ZIrJMbab/ZMNxm2UCokNmCtqkHw8
HoWMvZfmJYsSjAP3MZCyjQfLHZFNScVpe/9MOSGQON6SNcB81EtWqulVy673JDiZJt4Aabxf4kRJ
6eP+hwLYp1+NjA/HNZCShAmcUWj5F9Nw8tHGq0UVkdlpQMrBj1b8g0f2jQAcylOCH7D7xuJVVDm1
x2NbyUBqflnP5MdsyWs662MMI4zlPrttA1tFboHXBbinHS1yj4nja+0zh/qxIUtWaH8o79ikmUIu
w5l5MkSvkt1Y63ISBOEaBa+tWoV/C8Hn44qLh/KpLSH2b4RO5UKE8ikYnfs+WfhRqBQuTOOjzddT
EIh16zU/Dg3gdd83b/ffhEClfLYkPQbBQvYL2lYAVPQALE4WlDpntPJ1WB8MQdV/wHBt+vuveLPB
3Bt98B2abblrQM8CekM4y39BYbdngoCAya+FhWDrkAbeKzDEpeDihI0Hq0xNTm/ijVDJ+Gi5N9Tm
wEMtUge3LeHT+17j4ByHOiyT480GL+Ne1jVL3srCrEw7Asl1j49TZJTGLj5gdVvcFZjWkkvnAZsd
8kOpOYeoLb9rLJAx7rQIHw2mOZC7PT3+uXddVBsOPw1LQ9LK2D5Yzmel8FO4WII5Vexy97uYhd1r
UMzoHyUvWg2jC5poEpsjM3LAljeEmZDtsZVl1ExHzz11lcQ3JGWm8EVSeI0Xo/Eh2FznNekTrXbu
v9hAG3gMsBgHjU5cCGKZctSz+4C2oO9tazsvKSBzOS1uD16CHUCEKRUQBOvT+7AASQnd4U57loZ/
YXSVt4wieohJalZOwFlEbFQLyMbUs9JIXqYpKR/YCTyy91IGToSCH/xwjNKSWQly8DLxP3Vc2xzw
uiYdYcRzxFwzFeSDzlqTAOMo9aSAzRFoW4hEDXmz1VOb+IVopRLDDFJHKE19QrRvyHwVMnTZTFSW
GSsp3ouRxwRySHImS7+3HsxfQv3XYJ90FuMnbAbweliKC9TQH65i8NpYBsMs0U4WSpo1/veNhAPG
uroyzt16ImrkP/tJ/msWCQhf382e6cK/YeQ4TH2PgxYoWQg0x3wL0cykPi10xgj0jFoxLalcfF2Y
oLTxiT3tWpOvOBI2BWpWIGyUJxSmTOGx/hdGFYvm4WqS08DoF4Ud2wmQeCrU2fOLY3/UVnGNN8eM
W+1K+qi4QgscPL96DXlQyxHzn2ObRPKGK/kutYBI3nuuRVuzxrd8fYe2j4J5eEtFCjW3qwJHPmYm
Shq1jVrN+/5JqNSLAt9HsMQzTSYRtoNxF8SXLfpZwm+L2AnS0OSgSgr1+2V8MldCaZopiJTkxS78
JyzFQUPDoRigUR7AJV2zatOK3vsUApcyO9C528ZEXCRrnxF3hkt/ZkSA0FCQwsTvP6cy+iOp47hr
Bnq2CSiLq9uCyQJQ7/4IOAKK5rjIvl8cRn1zxvClwcZlMEBfTgJwGf0jDVESd3zotICczyHTkBuD
b3m9wWg7/ibKzr7FSs+pVl6nc4ohpEY3kJmj4lPqFV8jzNwRNXouMj3QTOPaoNSreqlOySihg47L
2zhjQH5XDcn899QEOUFgWHsOXhMXP3Cw1Lac4RL3VQqSL2Kz30bX3CHvrm93zzWi/a/D29W3smRk
bt4Z1SY6ruLTLnRZIUUgF6iWzI7hbLgUB5ID22q7b9FQl4+ZAGfcHpQBN3vv9o6kvs3/vEOtenGn
6+s0RDOAfL0tWcIcvQc6yo3PqAxuECglCV79ZkM+/hc//oaW2/XYFGLVeo2+Zhe649MVuBiwzZhq
4sTBCVZ2T0snmxDVnJaO7sCKFX03aAQXrByqyLmRWp7ageboSZETKS3UkwhfZZ0FnR5FcdgASZdt
RCh7LJFQLXx55K1dwZm494YXfkDy7bLFawTXD1nAQ6/1I2eiRyvOH1oV4CcQhDYWCXcjcx3DG0Bz
PM5rDchD+j5ftLu9571ISBJtdPimoYe6zoEbamJYlghUCuZZVTolNo4VkTR3dYU7q0psQYeiEpss
b5jIcauP3HPTAAEIXo7aPh4kzECZCrMcbKwG3EXQU6V+RXixkZwL4xKYjdRf6kw3zUuq6kWtM33l
DADH0XnN/pbmfceTBzdw2/hXi+Y7IRnpWEko4atEGvmiqv0DK3z5AbUizWSSFyB+yC/0gTv7t2Fy
/AJR0xW2mh/lJoO1BeZt5Ukivpsz35Y8djqbutxKnYWHT8T4I4lsXj1IdLszI1rw5h5V/YNMxkQH
8lJPkgiX2vVh2UEn1QmIthCaOeEiu1ovHvmncHkB1aYWOBibwCLtbiKNVbgh6Vr0tqlFG3Ywadq6
sg0AkZELnMDEkMUumXkKeq/5V5Ka96O6JQirOYdLaZDTFyzTZGnFUZm6AEqNlqb8FUa8LrVlsw9F
3zyCCfvwedIb5zCsHGvcyHc+nT8yh/qM+k2I/xs11D8AgijzhnhN998SHrnvXeSmhR7HoIxt+ghf
Ph+BoePDdL+ayrcICVif0MdWlpXdY8WRzNIJ+374hwc5MJjQleFl0J7yMJYSyjmq+drCdZlFDCRA
EfBEaXLq6lpP4fMTRT7RXkn2Z5i0u+EFmOr7tFKmtiywaN38qJ8n1qez4cuC5NV72fezrc7w71OG
PJK7MSBehF7tXUqpOVLjE9iGEvLrsdmPk2xeZYRAwq87SV1TyWfhjpdaEf0uo0lBddpfso+mqbC9
VZT+0V4wFT+Luyps+jbLDRESsittz+/8pAsnqif1dX/r9Yv3qJdIUXEPCS3xCf7onz4E/pprgIZ1
ZP3bSN0asaFrsFMEVsPR0hBnYOPveurapBOON41wdy35y60nzmAb5Db7AyO40AOwFjTEMSYH8V2V
0b01NfRGI2o8qWaf4HebAzKRNeYxHQXakHCLIYj/Kn0EbpR6ksQmJ6rtPtbAgoWZ7Iq4YDulj0Z7
UzpjhhhC1ImzRkMzlYmk1dMDPoDpNyEVuGK/cWd3DIl89PXH4kp6xEf9G4MIVtGefqRiUfWyrTLa
7dTpC9Zl7+QpCPh85rat8vBCNTis0fsRC/RJgGacb78e6wxBJ1JEkeJ5opwsh7EcmpggYG97ngx2
AdbgHdDrDKFWN/NfzRji/qx0z35OFPyJMV9AUvixAVFYZMw26jRYsz8iI7HSbZkh4LJrBn2/r7IY
6TzJO2AvZpEjHIo5HMpd9qPf37wJYILBg9EHUzevwQuwlZP/7p5e1w+f7JxLzPaOa9nsm69Jnk5W
W7IPHNIw/PnBTmHPO11dXgjdtM62oBI7t+lRH/EGxrhNRXitDl6CuqjI8S5WiSAo4/PiJtKvMmvR
2c3lnfvpR4N0dn53jwOiMnRAg/NlQBvEJqaE9YaA91p1JOfTyFNKbPXnrrVana9kj3nCbCKW8qzg
tSIsGLaaqGA++J8DG2J8J9uaHTo/i7KfAJIawgv6po47qy0mdQzRxcYd+fSfE4Lf8neGfpg9munY
/vIgSj/b2AyAN8tafjmaUNjs1b/Pu/jfJE2w36Zm9+Gljcyl/EDGhWkfkgPuqQ2CRIPF6AP+knDQ
1xMGINGfH8GmW5t1SK9ObDxX+NWKB2T1SpeGp3UohC6uKyX9t28FFKuH22noiagz+MyGB9bG2ByT
PfdCfPFVF5Typ5oH9/8qGuQFMj0MNLmiUyZlSYN/EGkFRy9C3wytyeUpQsnNh1Kf3RvrjH9BqVur
rbijWOpS8rUwyn1En4g9qPOHjSRUZko+GIdRaGMxduUFJIR7+KQ8UiyqVodDuOm/Kw8/Se2AaU4Z
otMv/XXPWwihasIMQOz4yK4N/ePQhXlT38FcxahuWQCuDnLB66XNPxZxI3p/Z5eS/eviKSqlPeMj
/DXiaWQhj9fKIjZ10XzclcqLpdttsT1pjcCwWiV8p/S5HGtUPYNPCg0iMtrtrWj4wT0udN9P4qjZ
oKaJhDlEI0vyAVTWgugvdjw7w9EIeOe4d/ZHoiJ1gM+1iRA+z2pJnQS4bVHqUfhHfdIhxvljeBhC
z7jX7DCcuq/WuLxuHQWf7MsFfiSnCM3ojR/dSxruoKv5B2B4FNGezBVOSHbibH5bFryShf5SKA1V
mE5fb0udDQmRmwlQEsrdIUoQm1nN49jWcbY6am1i4wENDeS3m4Ikp3RFm3vw8TbbeDFwxW9eQ626
Mcwiaiiq4B7uQJU8qAkvz2+ErN6La+11ynOcHvuKP1+dRs2gNwnD9ch0nY2biEaiy6D7KFHD6l0V
nZohrpglXkmIQLnI27oXLxLafk4scc7gOD8Eg3syrnUvLSvi4k2zoh8zDvlHbpGSpKYVBQFlGKpl
viNn8hcw4j2wa5YLNM5g9H3pDsLhHF+GioIFHsK5zZMxfmkFeubtU8lz0YjGRHs5X9iBD/WEQ5xs
pliH8FQfl0omSJITFtByd8V9LoX8fMd2h+b0X6oGh6JodaAWAAco1WWJpcoYmzyTjq1Cjlm4v/an
C0s/WmDlc1934kqJOZ+yruddtoXTWa8C4zkRsuWkM25jO9ygkb1GH3lkQl0H5auM9hi0Gd42p7Qk
mJkzAPE+tsd07u2chV8/yRZlhapkKTFAWGEC5rLme/r0oHPbWzr53A1VouYjn2piwUBrP9jKtNj+
PLoYr6ZpaRm5v8TJ2MVIDE+6myDkp6koUqnUYZCkF705lUG18BsbE4i8mrW2CDri9ZC7kzKqeBJg
6iMzSIBp+AC1N5AN4wFqWi6/SshI/zR3nHvjrHef9EuLggaOmlu+J73yBUOqcOoecrj0Jcs4CkoG
ocdjpkBQqlefaly9S/hgPrAeT5sjXQlNBk28f3nbPugGrTC16eixWabyx0Ci2aHT619LyEvI98LF
Mdf/NLBZ2MyUSB+d65kA6lT9eNT/YUVUam9br/ZkQ2wbYW5hoAavJV4BbNqdiJ/4KNNDTmOm96L9
J2s2PSAF5a3yMXgTsCKFuL+NJuDjn9SSlmRSp9ylpvZO5UuL3iY/atIumnr41zqOsB94zJWI0Q9F
6/zct/8a5gqO+4gvaVX5R7AdbfAmH8s2ZeX9NcZdHZ9rC11Ril2UVKqKRUibR4gFeLGTou3DId3o
jn4DASxcixz3z5nQTRLXHCd8QteLgsNfvpc9LIwhPzKsfiMyiFp5jOkh8ydEC9rhNQfeReOeLD6t
t6WwTnswME2raf/wUsNXSqA7yuqHqI8sZHR/e83dKV6Ny+Y1yDrdCFHj8MpHHsX8Sn7mXsWRD4HV
+gB7S079bnpwuIFkXl0XelvwjsGS8F/uT2GHajg+XvmLZqJBG0kftBnT/E2FkLC41OPVwxfqRSQm
yyXQlhw9z9KDsF5xWkJKRDnLWMMM+DGunuTWqp49DJ65JwcRDDW8Qwe/IQW+ZHsu13zFIlSwHcmV
XtUipR9cPTQUUpDfB80MeIfWR6x07MIK0HGezKqLSr4/eTOCBJ0tBGNxBqt50o1cfDBC3UabJQm0
jCLkmRYG6Q/oGuEOdW6/qHUjxPtQyJwRVDR7HiRfKLNM401I4A+2urowDPsnpBBVXJNqI8l1Z+Ji
augBLEg/8EChpqx3wjSBrdUhpNiBXit5YPb4sNI/XRL76Ewu+etK54goDwWgrbNWR9a29R/d/6je
d59Th/2mF/JXgJyywCKGNwPj4cxabSBcoB9Uttitrr9F0tz9bQnO5HnWSipuZc9Hf0Qfv/cbzMI4
HSCu/MK1/E8qrS8INIXaujrwMmvDvOuxU6hoakbsceAO5q6z+KhjNApzuyjMYtQtJpABa3N5jedq
pZxPHyXXYCYjxUYWgW1sgnND+adqzUAqOlneiJd0NvuVfpzKwU74FhWnOkNxCDC304OA+pM9iHS0
Mkl9KhfzYfwfd7Zb07YloYXiP9yWxYNEGeiUcBG9BqFJOnqRk5hUB5Dqj9yHhzITeo4nOaDlkyra
RpkYl8QZ2+arSvnFrIZ4fmYL3CEAUxap+VQqly5sIoWAham12zVaem34HhnnDRXXaMCM9VQehqIB
XtMKyr1C6f577yXhaa1GsTYdFVBE9uC11vrR7scIy62UYbzdtdSj5B7RnBuWETvfpfjaGjPCgfb5
PD1j+9KAhrAKtm3LkY528vneUSWuTsqQauzFmZewYUyKRLK9Me3PJif3xHpKTLdJdacM4PwHgWXr
7QAksuZKHvzldN09x2G2p39P0lgWDK4bYsGimh0ePiqb7TXZfO6ixniyGB4fyFnAk6GZ27/xcQgI
asYrcHb6oxgnA28p9Aq/MEJqfJuxMFpz9Cc/NajJCXbGWqw35U+Ob7San6eFoXToJ0XcnJ2aKFtg
/vw2+HuNF5hDFQv9ZsuXLAI1aidgLImkHoOsR2EOP5WMyBnaa9ybsAuctvZjI+RN42oMTK6ra9W5
J1OhsJH+HJEh9CxtB/LlOtKcdrJ7dhFMLlifV+jUXWsCMP+FSFFOLNW8x54ciB//cBilgROmkv8Z
LhWohdHErueWperVnUpqnjy6VmscDVMGXqCGlP80iB5pVKD71mzb/AQAnG8qqZH8/6Gwu6F9bI7k
1PeJIh3hlKNSLIYXpGfAE/KYhy4DsMwJrGL1SjyGdn78YKkgNO1zBWs8OB9NPsEyQXF2OPpaBRE0
ll323qwuPf8kj8JSF23Ydx1O1JEU9n5cbp697GvKng1YywdJ9tzz8AHPzNBL3Q7x+pQUajUVaz/p
z6oUjgyMsxRwvDQfTjYrMHYIuoq30EeqaUCDt7Lp6sWIrWwKcqqS2EDq1r8iKG+2n5hFh8/JYIxk
V5SCDt2vfYJM2RX1pOB4b9Z86RsKEXIw2JphvgrpuiQN77dQstby4rF63KTPGnLtYgXE2Xd3kceR
IKAUWOhkfMGKfkZXqlV1xNWn7sGAh7W2TPplg2fndZglaZbyhohKIFWqUhMWkdkeBKrC5VpMeQUx
usx0L7k7HME+CbJlv89tmnVHMtTbslH5T/W1L7Z5/wmcg8pn/Z2GZEYjppVenO8ggdyLQATPE4QA
GJEuJ9Ie15yFhpy/ycMlEHEFmMWNhvuBq+iNs/EN0LVeQJo2VM2L3dIAfXkNv5zNj98FS4S51cSz
FttnsCtzNLeDxx9ckd9vLeCCnoEIr0F96hUncDy0V6bn1ixlS8gIpNAMcJrJa00guQEdg1sz7xKC
kIawT33n097Fta3EqEjtwvIVQhaeKArZX61SPQ43UOanU/leQIBPporEd3DlrHjANDMucJ84d9OB
nWkRKXmfjaoIRyG1jjjXv743kymYdsugM29Fy4/3JYvbSefyJoK2Z1E6ZxPQldlEjHeXzVcQCVTz
xqO8hXW4qMYHMrfb85UyWJH/7VrWcZw70kAjSsvSbqW341ExLkTS91WSzNoIUG3gCarOTs4Gjvwr
8URXEtfrkRjpIgJPDWt0qXzX/fPoMvZB+J8ajO+ykZqfSSYOkOZ+knSQPu7uvYchtyOSuvRVkNb9
fqnqi1uhX5Csm09E5l1/DIqQ8w80fIclM8zAo3nu8yVz6LhDIi3CHgSEGDKD4dc22kAYz2VBAhr5
xTgA+7Y9EbI6TVBV7Wt0hBjwl6EuZZTZuSjFEU6fyfL7NMV7c+i64U4ws61yLBdq5GY50J4q/00K
1G6flm1imzrHfFHWf5He8aeco8EfyU/126tLgRVCKDpTJaN6HBEfD4cvatHs+oojbGLCnBQyztbQ
2xGwv+b8KwJ2Q3P855h037ADg+pJdSZ/pTH7NKPWRebAoo/OtOe9eBlWnZ7Scg34eqZhpdIRyOk1
HCWr0yvnIwVOy4t2NDbnLZMnkyIjjuogWAZYbem4tWWH2SIf4fa7eKQBv/PWAwrkC+JiM57rjuY0
nCDLocaEUzCOXwQF/UxKzCs8wYr0pr0nvcmGpbDtVFWwACPkjrhbVNeVmCSLSb1EV2OHetbPdtsy
ebYxrlyCgmcwwV5TIq5vZOmZbIvI9wf4yPJxnxdAlZXC+0bGihUEgGr4g0kx9Fwr/RIqd0Vu3NEY
EUKlzb8qypwYoHvOg5ZiCHBC0IfSD0hSPd9y/V0boF4QE+KhiSHasx5n4n/GoNOQeUzalnAnePQE
E81fq6rEQ96B1Vh/FNkapNeybbYzOtKG19olDTuuDrqLzs9arAtSuATFvJtuRq89Ns7xAXd388DD
D/Puln6CNe/3IJSAeBxVe5OKhukkubvpOSJeB7NL/3CPmU9k9QLSDWbXFhxIbO7tKRpYLokm1A+G
wxen2NM2+raiJ9wE6nBMzwob+/aGvl5i1hoKniY/rjKsIIoeHDllSrJ/MegvKVUWwJGhU23tTxWp
+J7koBjZythDJ5rFxFkc4dqY9K2w7ytKP5Fd5Uz0lD08RVvwS6FQ1W0n8BAe2JF88jGQAxVBiiff
dUxGnNK5Y7PsCZJ/pSLKpwcLmlsH8Zjl1X22HZ6ExcizsPI7pFLgAfwLokzw3SFj1lDLQXhsfW3P
OF2fMqzOeYHJKrONaS0Q72D5ndGHpoL7Bi0ZjkbX/yE1PuLm+lhGcIy9wv/62zd8LCd6yU0CbzCE
U+dOUsYiD0IFNi93TnokdJKsOIM88s/2tj8S9Tp1pw58FTy7ZWcC2kXYhiJl+wIUidaWwPSfpH41
AiUTFSCXdg/7BAkZZawzSa65q+RnNvXpp+0CnIvwPgOzjtFu4f1VeD5bEsDkZSY3DaTu62C3A0w/
+7nNzGH9GlwT/1LAss6JW/64afefQPfvLiuX7hFzdzDP2qc4jfq6KkxXkPBALOoPwwfeL9gktVym
YPm3tfHaH0tNi2uIlYnMbCYt3VjCc9ovbS8ukagRn5LFLfMMt+rsbZ8TaBbld//lCIuoiAQ2+4bM
B2kF43Sd6b7dVSFZexTPul0lmddsVsHftx/Z2WR4Z5j/3Xe2AUki3p3yIBkwqAiI0wJrYpGpsGCp
kzl2ZLeN/nwV5PX7NJP1wdjD5rYhTBkTNzbbvrMpiYRyToqxS2/yHy7tm6g8GwWPTj6Syvt1lcDl
ZVKkDFqlZ1ZeASwj+1CXQKP5DhfCuDHmCu4OkrvjjPSquk6zM2bj/QzjXUqBaSDnX88UFce29m1f
nBL11e1sy56cQjKxkeQP8gLlKPKrd3SAEz1ElSxEeLurtozH6u/q6b7C9nyhbWTkOWj8O1+kj9vH
670ydiIKFKxRliHIlBjMnw0UnEPmjL6awCCLcXfVPnzdo5AzDKE3nGxB5h7NhQCNg98M9x2LZ3Ma
m7pDwv879ekqlcYnpyCnb3V0lmE3+wO8wjb9fbRicOpJ24TaLsRIVv1YUHuEqWlJ7Vul5YHmxVvY
xzzCLM43O+x3H4oRy1Nk4UcSHXewyH+uynpjIs7ZzC9fTADuU2fX1lfQN5PnpARX8MnOSojC4Mzg
0LTZwmlJHcyFfS1itpSOD4Bj3pY9czioLc6SHFRSTv25Lp7YkjmnC7feOVXI3BeRnkOIMk00Y3tA
VOAMQepqGVHL+l2/AnaeqVBtlyBy6twAmhNt6cYEQf1ZB0uePEWfmON3dftxigx0Tea3BEIFxJcX
/dAnQX+UIJQmaiXAw0cHqbcHcZ7tEkb/LPUWFIZ0nZjQIjkk92bzPsTRvfJkup/BbU79amyug4no
ehdnD+9i2m6H2wdcAX+HRCzD8VL9psbiqQvrtQa7esQg9xbYE/NjZkBoEicQfbRSPQwdkoBsI+ky
20jTi+ilBZx/uu85ppimGQ5bix+RZSP0pNv0VbfJ0+SQag/UBnAYeNclI4XrCSD0yWUytxs9u1Cf
Fy8cxTuVpNXcLlCxsX+DzJDycpgPXn1O/AbHF7txBTBnYBEl6U+xRibNTY9XsTmXLIQOS68Epr24
U6JjRg/ZG2J91a6OIJjFBsDpdp8glrs5p239CBYLJoSOVljUtWN/Ewv6PtN1fYBVG932j71E3yap
/UQBx6I6poYoKO/C0S11r1afDUwQKHY0in6V8ZTCBqzf6mLs5yyJEWKiWDk00ysWcJymKqz73INZ
FaVw267K+VueUmuRwxPqybtZhrgwhTGT3jrI72Z0Dnx4KI4ykYN3t8Dp4l/mrETzin9TTdiFvexH
ts69t+YGEXOdXyPpnlp9/t4Tvg3B47x0EoSotCcAb0AtHIEozSmjg8echq65Km7VtovyTVzj+UjC
QfbPsVQg2OwCwAhDEG8VdSATZZgbLDfZo6bLluzJrs8kML7No+J+KaawZZHSyswGdQzTQ0PkbtCa
rnCS0VL2zH/n+RzjPbYW3APe8IirpxLiYkrGDlNgAiob9A67h3tqFEsPfXUT/GFAVWgacKr5t7Cl
QahvIvZxYrNuFosz2dy0qCLc2n0GRjASzIkpLuaEfQ+rFxGH1Hwm9mcHHsAI9Bm14J3IosuLfEbX
NPkRKJZyjsf4jExiC+jzjQsnbxoNkbPcuOGPuIDYJCV9fweVY5z0Wgh2FPyFFRYlyA2z1pR08QWl
lmbEu8AN99c5qlHioJNuSrQAIxWYdw8/OmSocgK+08Q/4zOSOgOBEs6UZN1TIpw0lZ3xiVW473kZ
E2dZzY6o0I50uEd2UTxpXwON0aqki9hOaI3zrm4ok+jRrjhR2l5IrPMc4ziNahMk31fcFjDqTfrj
8Fkx+2eiEOBjIBzpPxUnl2oEj1lZh9KVg+pyCWoceIbTvNaHTAJM+zvdQp+BiemEakssld6upQ1d
1bZSj/0Uz9pENxKBNxIi1HoWkL9yDWTYqrAYSNbHFkoa7EWn4O1vGukSGv2te1uYBbGVbKJdtS5+
A4nj45uGnISJOUEnjh5QYSwKPGgbOcnWTqs2mOwl9+5PvKTZYs6uAtPxvrOWVFdyMDifdTIMj+Qb
B7mYkHVbdnmVykCcfuJxy2n626XwmwDjdReZHHPbzIEkYbzxl06CGn38dvrr7w8Wfv3VGjk+C/dO
qmV9teQiL8/aXMpvKwZBF/0RJ0/VrmqCpCjc/7ixlFGd30SyCTNLKBOmz7+emOsrQo0KLry6KuC+
ZdAr2LFPvVAqtZgwcHxqzF2pbqc+UuawNCPVwODZCtwPc4Rda9udYlHWudkta3rdUxNRDbIzESvG
mRL9IRzCwUTPulCrY+OVnT1TIPfYeXefIHxp60JmVj0sjyt8h14A+2kuEZIJHUckyxT8D/FCAzM+
BgGhUmpyBIMidaCsW99MTlV5K7RR2O59XXa3G7ycK1K+X//fdxlyraDc1p7jw06RvamI7i8dGjw/
XLqi8UFFUbrKnzTrJ0End3qTohWTDPtxChSWzkWYb5iTmMvH2et0fJJaO8ZvzlBuGDMhqJez8T4s
1RjZD3xTuno5a7unyOvRJBQunuDTmkbxKGmGzD6ahwNFyHzsE0v69NcYgCZ6UIfUBz3WSCxdO2Bp
VT/WNA7yz5pJot8986hGN+7MpcMIg/5TYzs8Xr1eafEGRt3Cbqe60pmqio489/8sXlWl3R9TDGRI
HVDM7KPDk9oSvv8vBdsskTzosCi0CtMx8TVWkxKcmYPPFw0xGxvEZbvKMa/leOOKk2p3GveHAGjH
ajqnilK1rfqo4dIL+j4nEjdQhnK84Z8vG70WDyizwgaxN3PjCVF6f1logi05A64mCtGp0HxwlDNc
RWzHPFsXVy15zblSjvHu8dX8oevlLfmDNqdaMuJJybvkRD4veFtkjer17nS8jFldQuQm1h+gsrv3
Ja1sxzEOgX3BNaDWc7ulKFwQ6ySajkx38UHWVxZ0hZrLtMa/zpnItc2McwgEKCAO9YGtQd3B32Hr
pkzvkuFVzhE6pgWi5z0G88QVlXQqL6tSa0y56BDdeFe62jgfbhnyI93SL4T4hjWQj+yYHEZTDdNs
92RAURBIBBskFdy6OJi5GMWvcuhFwSe5FhxA1sYw1duBQulhR8LyC/huWep8vY+kNijMg+Fabltb
Mcwhy+wuONd7PvvxDvyn0c/oBGAwh44GgtlbhoSQZHhpIKgJ2fKBQn+QYWKhdM9sc4dwTF2BOT6S
bKtIhOKHRiBbs7l7ADOp+IaMES+cMD+o8MFnjswHH+haCMJ/+s+kMb2k8Ay43h/ICgxY4pUPB/k3
f9bkWY0Gjg4YVt6j0t7lb2L4w04HH0KLYgzdC7VZ3dtBr85tGL0kp/OngE3HWJq945owKPXbv6GO
hO0Wxboty6GGhxkwbVropJVqx4FSJBXDloBvJb1RBLi9ochY7C7D1CrMDOiMlIgR1St+lU5iUgQd
aeKcf778YHpNKjgg4FOe4/I4dLIfjVh541iPKkVQzsvgeFQhQw0TqyFGWJgmknGXGUdKVcbUv+Tp
4RoSd+yDCrpKRo+dooS/LB3gyG5ArIBTDxScKsnpQqNuB/Tu+RJirtiMOut9pRlz0yvFGcacP5gC
EzEseY3PhdBc8qPilaaZbGib4Bz4fjG3lfjzY6wuQrlrFxhCrOcmm/mXweS6oIFpz3Qx7otSbI1M
mQTYPsqXOX1nhYHq+1sWn42HSWSYiowvwhh8uUyZneD1rWHzIOnBseCLatLk6EzVnqMerh1Wmw7K
WJT6cj7E141b3HNf934SF2mdZ4tI7ryWJcFLHhknDYPcPrfqCLpuTyUdvVn4RXnosZQXCc3SrYW+
ONgjv+G4+GDfIEjJQdmFFYxpNdAlBb1f6pwGLVonXLsqvm3LtWuvAsq4karhaYjnhwQs8xjLTzt+
geeKuwDdQ0jC1+ce+NVYtY/DYwAJhGN7txXqeWRKXnZVgkkPpCaXAvFFew9KzEioOPZUFmskS7NQ
ZtqxGFdD62EqiPpoNdMRT4mDilsY/JhLxguvw59KunK9ZXMnzX5yC+pcBjfh7MyUPceCp/gg3uAw
sAZc9DNOXGq7K4bR7TN9axZxVNZl+a5oEZKgI4JFSIx9iqh+Gq8AsE0I1MrfjS+wUASn4jkN1iFO
0MTt1yS322tKRVM3cGIj+E7DxiKoKOoDR/GCgPPq1yMKH7g7Lvv6OXHCQWdjLwV6x3IeCfc7fMhh
lsSc2VPyFuSx5QMKNTWwS/L+TYwRBszjyg4UtxM/cQjtHpTE1g/qnLYKSkpZu7mBFw9773rqdPI5
r51xFzxxehwf2NiMPzb0BuPJWqzZv5IjqB53GYzW2KwqlPBbRhOH6j1sXx5yZjel8O1Jm9u9tXNk
lsVb84A6a74kgR8TxamKxCcJeID3wJDIgqK6NbnMPjdtv1FW+ZfNfhxDioyFM6Y2nPesj8VYIJak
cyQ2XmarTRi0oqOa9jJd9UW/LvWZ2TV6aVK8g24e9DsCv5wcSBRP5QB32MYC6x/ZgEgwC4Ly/kY6
F/7ZIQBXIKh5jdE1dYd+X+NmjV/5+8A21zyFHEfCItLDj6AElNG4zgf+e/i8u4IxpidmUbT5mg1d
0nFPmSa2VU3HeaoldOVcW3QFGwxi8PL+/9GJPggcOMf01t0xcmX4AlICGuzrdQK6MKmlq4i6prsH
KW3z/XbIw9QTOejqbuoPEY4Uz4Uj5iOWxflimFG68HPPX8h4LT/Ht7Awg5bNLTea0QGio+dQvMsW
hTRxcU144nj0F6mA0gsST06mjAbd9KU2ZbRDKRfA7uL7r2kZIGpQz38s412gfWqdFkHVYzsZfeE3
fV6c+6iqUe/6s0qMA5sFg2wnDbGGVpBllHFhyxpnzs7eLiyPA/SgzNYBKtCKmBTW9DT2ciKiKg8i
so5BMOwu2PlFrzRqOjUGbw3l7jSLVdL4Y7BFF/L/0bjKm83TOfExVZDcjGhiEouXD8yBYPwhKVAL
ue/LuBWqdCfJHf0+KJpN6KnyqxJiOp6eNwyhgMuN7c/lrZNTsfm1LZWEDvjGqdEt/n4i9S/oxdUL
xQHMWyu2aM2T5FoES4zL/arXvsSEhaeQ1fVisx4G+cwuNGv8XaQuwuLAqkdA/t+XIJqdYGXLoBbx
mf0i7TMjkYQZgUBG4QSLYSd4ipqmWFlTvL5ik1mBKsGlvJ6CVT7JlXdYBHconTI+vdF09joJl6pJ
xcZrXqKQHr0cJ4us39XX07bZLBiQ8qja7huTk6aX3xmf8xpB8Lm9JqvvAOddh9GUZs1Eh0XVpvW2
V1OfN1cNOvHZrILV1LeRfJT6r9A33jKkT42Y30+RkYE5ITrr+jcP/NhlushVoHXicZ8X9V9qx4aJ
Xr0SCvahhS2pKj9RN1fHI0Is2qxeCJmUzC//ed50HdxmT4kHwf6xNkyGCLAmkF/J5caiadwm7Zrm
OAC4NzQgwGMEn2m/4Z9D+XepQRyexRI5yKcZ/TA0wvHPbmUN73s11i3tjRBNMRaPA9oyu0rgAlH3
BtaqHoPffnummpfnzwPFNaMnsY3WnZSJ3pTvHMxkH0d7Z44v/CDOGGMvGMWbv4/rZQmI5jb3+FUF
K385+vuKxINAEV5WTziZkYdmI5Eagz3/lmmSqOFJafpGmPJU0OXYu5tBdH0ckOMQJEf/GapYyzJf
WFwSLKhcxQNfAxrOKkfVaVQmHN/Dmv7mL5Vr8FbJZjC+QHqYw25I6tiAyyaqqTP4KYfpqBIRoY/D
b5vW4kl+gGUAlpEerfq4nyyzDnLGBOKCvGgoJQzPDT4x59o0FbOpFF9jCEqz8Dnnu28rYLaEsLND
d6P63WxKSv2k3UFvrQlZutKdk1nhsBnF6wWxfdXjgY7lohiOR3jXCzEVJlZkWiCm65HtvPJK04ER
dy5FSwCuP07p8ofo6lYafaBrJ13BrhV9CrnjpVedCSk07AA03muewlrjP1LKnl4n0/AtF8iJTOPY
BAM2gx1s7cjuKlLWL7vRU7jVK0h/zaNl8MU8iLeyD/0gNfTDOKiBvK2Z9H79zPWQuX2VyTjZQO8f
Wzxu4uRnOR9m1SBCU5nm2/n3pC0dTbDANiDchGbNJS7I6qidVhFKTuMqQlb+Cu/JZAKOws7W9Wni
qfijpTa90OTXB/k3/U4ca10DDnVN2I4xL9vShZVRxNLfkKimJftjWkWdveaPbWFBnVUNS7ktFaJc
UytALIdRCxlTiLHRQkPOPjWZGKZMkPwERLp8NbP2TEIIjdSQ1TSHKFpZwhQ1prn6wJLl8iFxVDjf
1s1vIFkvOM3mdBJgv5CvrApRXaFnp10HhMo6/FczGtK1L8iKC4iNNd75OkzAFPKiXw/MeGd+UR4g
kKHFr5VNo8xzygldsow47BdCOqglLPCzI6kBD+1eyJ4FiQ0Neo7OQ6400hKln1CFNQME9sCojWXO
TuVffW1w+szZVtDyJ8aO6+lIcDla9lsjwtDg8XQbVlnC5dEGRZAdi8GTCflLLF9hFeEL2u8T0Id1
g5ixreklLG9rQcEu+s/FWZFVJCzuB0ttZpBDvkSW943bus94TrJ+u1e2YEFwVKksjGmOGHEEJ5+w
GNbERvDoSQH5z+FoYNapFgdaLAg79NhefAUUMbjplHPpaRDuCsBF+DGiPtUnvY2rIS/JRCyuwQfX
mtt21YYNIblu4XeyNObHsGa0SIQ8GW3g7kFRUbHzX8Ao8uhtjuOfI0Q2zA8RtVJrr/mqzay/+qml
BmMdkpkCy1ReqNi8UtVAC3FKZf1YiJUDNZMZ+kyKbQKjwtejLAuC74VGyjv345+Nix3B4GuJKsLX
OHjVZvzFgMcN9bpYHE46nbV63zB5M0j7f0RQbFPECCUzHQ3X/q9eaMfOW5HH4GgyHtY6gryN3RWt
wPj40+3YTgqcMQOW9LN0kgvEMMzlcGWhhXiA/HurL+bQ6c+OFxSuqzDv6aPteY4rpa/BJXFphuwL
Zd89Rl7Zje9V7BmSU1wx5EL7/r057H4P9Lfm7SdIIOy2axcN/hUlj1bI2XTL7XdNdAvNSgYVF//H
cfAeMwSzZYBjafCFOjLxBiulLlxgszyZnsaXa6whxdt5Z7YNPTW8CcO66jkPcBH/Cju89BarE9TH
PLO/SCH2ogW9ZUkQuxK38TvaHTwmgAXj2/l1GtjrHc29j2Fl3a4OdMv4+ZVwDvYLA+Q9ruMxphSV
zCtn9lbGzpRX7Heei5Xmz0ZMIu6y9dFKQfhrDEFPM96bTQyvZCnzDqrIRGKsz4qTwthbiuJT8qc/
BkBvtWYQxGSOmhx1YcorHG4WRKNYZD5vialrKOe3v7c7J8XuWMaB+k276aSFsmoEUKLrnCmr66nO
NAhHtbERnuSRIi27Qacc8Np4cOQsF190Gb2DKo2DLmp4lZ4wM+TDi4b6oRogORc9f38cvIZHEktC
PQQ2Dwd1v8OOm7NNR7QQcF2p9ODZaAYLiXoVUHK4/cuFPcSyM+Q9/oJ6JQd5Obpnls1mcSxhR3eE
oOG+0fioAUtuELbxrpXMc2+4SBXzQSBpPgZX8ac2cveNc2UOKMj96CdlwEV3HmakXcF+5Fh8hWlz
1bp6mWFKmsgLtaoKBGnUdEYMrzdtJEFOXkoEbPhHpsqsawhPb/TiaXJLnMEzh1lUKvstuV1t5lHY
2cuHjMUuyL4vK0/VDrt+LnUP/auKYae7Jz9kE0OyanDJcv8dgDICIs1UL3QPA2IKH+2rOkcCRPkU
cbJvAIEDUID5VIfDfwOEFPY4cqZ6r+SqV9hG9XtCrjbQFy5NrPWM9od4PYho9TeMM5n9a+pkwn7M
IQCZO5e07T/NX7iwBZgbo86oll1/NV1VX+wHGTEFxMooSGDqK5oMfiRo/YY9wRXTlH1aWkByay+Q
K5C/TEeddBIg4M1UkedE82xctSPy2tiXDYduAVDbduy8UND/lqAksK3XjPfAfXOe9JSv28UiWhQu
MglmETKlT+fRK5kGXybHV/x94nCUlHhm2LSGFy18vjiYSCh62C9Z7eJ0Q7yykpT0eKJiSqJ3gQTK
Nxp6ZEYh5WMQ+pnbFy0NRb21SQtMkkrmRVeqhERTsPhTkuZs8PatrBmDVLrlVTZ5AfdSbc6/aTQr
ev7nDe6Ppashy6mdvMst6h3Zva6yVl/eVrOAyGuNxlTLy5azFnjc+rysixvWdlEaKkvcj4fI8Jfx
W4luY/VrOV/gi00tkCvTmIp17SM4JeeJZnlZrbXKD9NXZWsfncf5el9+s0OH07dkr9sKFBw+e2RI
a5J7IpkO8/KCipOzrn66JLcrMhmuOItL1xnLB9CW5cu37AueTd4UvHX3kvkhAcnW4XF7MichFZmk
bzAkf9BW1ycj+/YDae998VVy/BdOlAlW91glvJIM/HsX+/ym4N4TrFn+tpXvcSlui1f837EVlEuc
QpRAwSc42s0T9zupyEAYTdFLpT/+tBtL8o+aFOv9x2iFlaxN5vw+ke3v4Zbm+r4Coiz99QUo7y6Y
Rpd5Shameuqulx9cl5oN3wntLOc5CWfjxNEAdx3cyClmH0jCwNDFwTRx5cZ1VA0YSklw0e6XpWzK
ON96P2/LE1gBRD5L4yAGn3RhpJc8OwF2x8akZVMiD6eurF3FEuJap8JMJASO/pfGLk4mcLNhrA54
7lM9LGUaGeAZbMkf6caGafJXi+bhDinVOJX0cDOD8RDbW88rL8uYissEtSFsn/5RDWnZriRGlgCw
TU6FC3Y4UawDrZw9v546OWnr6jSVRAOARMas4q3N2p4xTkGThFjXoH/LHfFmZ0vwh2jcH60l2DHE
FGTPlvslOYSTVzcWsJzJPzwtWoh0cnsKF8f0Ojjd1mMOnPAwivOfkHSInEwOSeaLZniWETNUfKo4
zEn/aF79Az8YY0/chXeap4+cHhqAU7l8DV7/U5MFjNA6x3ogf9tOIj/fSahcQ6X7o+FgekCKHUqK
tvXaJTowebaD4Rxb62o0cD10bpJrGE9Ak+rw2G9zw8x4+waWz3r3enJ/+S0D6ZujjCtAeDk/lZI2
zigEJ8Agrb7afbYaPS1cR0elYuiNXGR31m8JdbQ9qHIe5qVi4+nSowkVKvDhBPJgpP/Z6L6NxOf2
fAHdTWmrLwIAtBdqEczHA362gcVgwyeKZWZ59i8VKzKD5/vOxDZUJ64kzg7chkAHI7BHx+YyNhZm
l6NlpICiMOEaiuRWwtmJ+BvWgviYqVq9dzIEAGOfdarXpaAdNA4SZQymk52IGbcclPkVr9FjeWVs
d/jnLo4S1oj7XaMmbkVBJLNeqUvQWtWeRuKXq4YcBrtY4BNic4wak0+t644HtHv6agJbqg7Ctswo
03kAoA4T0iQ64CaUeeWHYEyY6RMXJB107Rfwn1E584WFWQL9AIenI0JC5kWLtXKXsAnJiL2bQPWh
IUB/SkqKWxir2luK4VTGp7dRdvhYBgqVRCYoAO4a070fFm6ezJUSWxE7xDT88gY4nz2o8F5vldUY
5qe2e3sHHHnTNGsCtQbZIXLKY2d3U2J++cfozzIt349b5FDzYaevpKnlUmVt05T5VjmT0B+08FPJ
tk+KNm5W78Ue9VljR3kngV+WNToKTjepmLpy/2/4bvJNRHHZDA30WDiQ/1i2QnVesnrlHEWCq9KW
0OvgryDwKtpRzpPXhvSgc4QV1p+H8mFKKccroA3AraShZd55PV2a6r4/Y9ZqG5G3g1J9G1TY+N5c
vdwOWUuZqlIDRmNJ1e0yFMiq+IffF0MUKbUdTn8r0WPQDFvKUdWbuS2emHu3xfgIo6TNyGmwWfqF
BV0jKf9NPMERwUuvTHAnypUp5hqobIjZvUokwM7qoH4M5QeMmiKUStwczapKz3eLggcpXEJ9WhRc
mJrp+rEPsj1VqVCwIP83kPKyxZba3cyUhtP7Kim9gdI+Qp2A9YNvLABFTnpVz/SH+d/uQ6sd2uuV
4plzEbC7mAJEqtI0gXp0mrJfs1MZ4w2uwg1qlDuFg21RvcMI+nad2K5pxDzL/cnvoocaFk6kUvCK
mqp16P4MQl0AP8JZUT1Jh+eJUaIC7ARrFmQlWRqzqfHyLaLdTIWyzzRvA8AMKSxmzCaX3u5IRx50
nx27I4fLxLaESBY3fpc3NflbCwq2eN2iznuBzIKPspIFQcivgIr+F7wk03bOO4W4xkizpFxIJ/Jc
Ro5e3+5j3+Pfajw/9/Wq0Quag0eT/vXwS4wozFMa+kYEtwRvzE9babgv2aFaucCkgMQv/U/ONuU+
i9+QxB3q8VCdR4RRqgnzK3GyMWRAX6X2uqYhsIEE5yPV5iAEq7brqZ97WmBqGgWJpwh5mc07msGB
eXB+vdHCH0SxF5eeeTPMDch/dc7uhRhBvKY6ioFslQGkmDkdT/MzRl9lyBuLgQ3yM/Nc69J4J0sB
ClD7x/M5JQuZ5qa8+gLAo4GUrAsD2Ryh78GebfVFucUA6lzm20KQquQmDdjg2pr9z53Uz22vCzao
qVKJt4OWMuDmXMZCOoqwbEKF7LcSHD8T2N1/AmwWJtnaTPDK1GlXZ7F0x+GCNfyu0HpMJz77YLSc
URa7C6JMYWIVuGCbS/r776h8MxPkS/nh5pYrPCDK9ExqPqVcaFkMUy6Pdhgi4Fu3VV5kRb4RccGn
owi3T1+IvY0/XnagwaeUIhYsy9pzFW8Gw7/11kHB6ZaVzgRRBIgXGl9o3KiOwwe0WgQpoOsu/Z1R
YSM4xDkTWV8iIZVeaKILIyTpHfI8koe22to6nFOZxUUZHwuuB46aBuXN7XrBU2b+EdhTjM5tZ8SZ
513Dv5NFfKAJfyyAZmjcxLeA4LoO0mYorlYjvEqH03hGnYJoHXcZnO2Xsan5mxOm+P6TsVWFIxkd
7BoXa3Phcdbyz28+CsR/rw7W0f+fZ3hh+5y1wyvf0LzJJ65TQNRR3aU1pWtqPbb6UFnPMAuLMfc1
SqFQ2H07B5C7g/dFNw8gyFTSA4yF2j8plw9KvWtwb++G+3zxj2MsaFHzY3aSMGyU63t7ZJoQwqFz
e0DWuCIfJKuY8qcvfMqmuicW3IpHbdpx3Uj5LLbc67Mo1fXlq1T3h7jGnjunoV6PoxSkDeBG+RHH
6YhUQ358EmqHBqPCX12A+2pDzXpyk4v1hppg6femY0fvqOp2zdwZlbwuP+6L9LM7nCE8Yj6x5G05
+E6o1WZnUwZRignPqNiZw4pbWg4BsfgV9HMp++OUFVV3D96GoALUTdyn0LenE85fTSvknKOT5ukY
rbs7MT5uS6aWPG35BC0XyLxGB/u+i8GqV2/BZOMiXLCfcE1eW63AZKtbmWzfYZYpnzPEsCw/J6Hv
/avMaztFNFYIsGy2Yvy5Y8TYAvdD1DaOY//hcYpbFc0hRXRgu2jOQ1MAGSL0+nHSbgpYF94j+TFt
f8Q64I6ge5H2LRK6JjMmqukZLCBCidLJ8FVbo/KmW/UGkTnGmoqEwMni/2+VB3z8Dd5CKn4/rqXO
YHt3L4Ylc1Yg2OZkMymPtd05+DNu1tD0saLh7XGI+32Os+S4NNyb7PEedodT7lBjyl5796eRYhmy
kbw8Mcn1IijqfqEAuaxNt42v5nPTXlpKpv7/3cj713+S3Exm1fTuDOH5UsSfIOwqQhP4/zj4JchN
NMh+4u0A0ZkSxJ/XXWypPb+F2U/sBWosNy8sYGL1BNXS3k0tbclyDOULo029KyOQ0ub/b9EMqzi1
W/KrTG0CVQO1229uMtWkZ3+wh3DEbDiRXvye3QzQRBgQhfZ1+0LcQ9+aaPHuuALr/FI+TEPGniau
EYARJB/oOyzjj6EdfKgGu2IptufxDjr66Q0qhWJ4YTTQ0g/I7CLa01dQ+aMtSp/LCg3FN2pQUNOB
jaMNk7EZPSyAzBsbk6JwjxSVEz3wYmX2Qrf+WUsFwld+gkQACzJC/FXTR5MclH7CEE4olM2IDn7L
LoTkfL/oDxPkHDplrMUTHEQ+mvm/ErEh9ea6Go8bUFYA8TPeQAHpqphSJs4sD7PaxgoaDA20T0v5
7lJwg1qcrCFCBCReeyuLKSgbOKNIgVheT1Qjw8+ptUL+Gw6LIp/As7MY6hheWGaGXPGH/mVv4oII
ID/x8FaDPTo55C66dAS2Bps5f+xk4eAt9tL76bBSlH+gZcbEZ2NL7isYwlH0vS1TMUlt/IIC9yBm
QOmrIjkMEnRp0wwf5wHvR8/GKw569cEAULmsryGlEfpT2CyWVOoxus7pHU3xeTgYKhTKFnSRLC79
hNriOIEr+xYxPdHMOUiILpm73q8l7P42NUChxWGLqTesC2nhYMKZpbmczao2T4Pn4sWa2F2RVH4M
wTFVDMVBtnn8v6Xa6viFL9VkmdY1qs9zVwKeCSbDabHIOCJRo9/z2GhBq0VC3bgluOA2ja8aqslQ
QFPN0hrQgV9A4GyQ4isYUr80twzWsymz3ec8/4iz2aStQs8Eu+D6TW9KDdPfmIYx4euclOYyBYap
17A1WYJ2PeT8NYEIkKPVSIuJqjaq+MQ9Q/CvmIHdHj1nh3rdQN+AfsFM2aZj1aQnK05cRIs79JWK
x3FyB5fwSr3kGOY9Ajiw6yqjOCrRf4M5kLPFq2ZC7T1YNWp70++o3KqiQA4KpyJHxxCO9f7UfY8k
tWHB4nlvdV4F424ykzGqcyIppjgcSEM0Jz2HvKrWDWZ+Q7bsBIHqPSlBPfivRtSX5HUbm8ojoBRY
l7lnEH8Wnwhh2Ff25BCOl/JBYKpE/ijr8WertDdZOmzP1QpQr1Xygl8tkvDRTAArergPsIB6h0lC
f5TUiC2nSzm4XCbE1bsWnmRyjtWff9SvZFs6+JhH1j5aV9XrlnxLBAd9iQZaDJ8//i7U0QVRYoxF
MiVzLH2eSJX3RjtS2hgfFVvaIct/tjk5nbCeByrcYjOFa5NPrd+9nPSVKNL8nSaW3EE9bQfoBKzA
sUloOshanLbiYFBwSPQqG6ioP30c3krBQP2Bfi0QV5oNw7e3rLBYe31Hqi29GvAauseTBdmb70BH
IcYv67ZxwkA6uZxCtuTYzNbR5F9eDDeEnnXzvHyqwy1n+c3UdfQhVXwA70Q85/rSQSRTJxhFDC/h
QUTglsVyGL4rOc9op82yvsUth5Fv0PFPnFQbJwtuQeJJPU08M2lQ7gh1yVhvaHuLo63s8qtDLVoH
vi9NaWPZrU8T4FPVaq0RI2XFKcdNhfmGTNlkcqk0JBcxCru4pQ9yw5Wbq/jpe4Wdf7kwjVeV+xG4
ZK7BUsNSjcfoi4TOnbrVrCJL5W5H3NoXGLOWF9brDCLmZ/2mzKr+VsAXu0hJRqd9cpSBXOtXBGki
2PEXWwCsvFr+iYja8gbqyV5uBswNlg0igYYYPCXvZFbojDpiu9w51gBvc/qeGwx8rb4qbBbY90Mo
ih0vpfohfkTZnX60VDyWhSst7xW8hCP+YEYg431ZYCSSvZZHbvvv+r/ZnnexLOGULyhPrbXNGiLv
vdQyWylqMTwJLNRF1aj6xDtsaetqXj9nVsNP4ZocoFcyMasM21xAOALzxOBHhGyy2H5+9nNzaq4Y
2ym/Dljp7qU4mXaSpzPM91m81y1YwVXvtvi2KojY1JQE5Ju1s9Oa9UrG1uJmX6U8s7XudYm1Z0cG
S0UYylb7u5IJFq1wK5hoEaWjOO7I0bFJ7mp7E5yMREYUhbuxLB+r9XtZncQXR5en5hok1tnoN6Il
jRMKeev1EyQuzqzURK4Jf/7EMMo4Obn9SYMj680J9cNk3QbLu9HdmabCwBcBV6zC37nNDvtNSkcg
dbdqd5RLGofgsqI61KpaIg5uzeKRNFmhrUJxqi6ye0c3DTuqbufXoUzZXWHk1Mlw+IGUydA+RZNk
z8uLCQbRkHSnghQfm4gylHmnr1rjXZi+XcWHn4BA1tFhYKHn6mjI8aBbM0Y//h+FUSoVdHFCl8R5
OqTMECGo9/haRIBc6CjjqHTMfItVz+4vq+p2Gw2094a+WqEs/A4jZgcE1NctNyohu4exOytop+6Y
SQvmNjg6KFZqABr4nZZStfLejIQktjNKXZFyYSocYn+//mXgzNTKi3dYgTIe2PGhko3jLGfKUg1o
v04ZhG7i7m2Lyky8iPgc97yu6c76axxlQVEgl4A6P2lEaLuXBchr7CEcqkpx/3MUaq6gwAXdp1Ul
MQbYdaINnzDtBt9hcEdarDHqWGU9B/VCBpxD6DQEEtSrGxNt41JpDZyVEmpmpadAo56EZtuE8TYL
x92pJ0Xgu+TxqgfBBmca5D/jD1edDnTUJn31OmFzYiZHVDhFYcYnwZN/11E+Gm35CVNzbOEY2kcD
GPRlx0KLdk7BGL6d04CutVsmqSnnTePevd9Gvt6rOCLAOwQSA3fpPoEGa4d1NCERbtpp6Qv+7rox
hEldsc+4rwkj6PZDoeJc6x03BqApHQSaAqPljKf2+XXQrATdKva3eEL9oKwSAkZ+20JeUInU6hpn
n5B/cc0SH820iVAWkSAV9tRK1iFKg1W1+P7ll3s3qJIa5wUvQK6O5NVDgYxD6PvUUlG35y/wMvOp
BcEDbN+BdissYAhe0YQvqgdgS6lP5zZEqJF8t2bz6waHFXP9z/Sp9dxSlS2Sh0va+Ehl8SpyNdeH
OyxwRHZ2UAK41OBcYMlkPVe6l5QOrVyN66+I+H1CnBJvVS6R97B0kfP/G0t3W8YoPGa/R/0VoNit
Saisdry+kNzzGzT0LfZBQTOFPMV/71cx36XngDkzZkfLwNeAXtrI7bWxHOkg6cZDEmaF/R5G5FPR
9buPr5P2XnCHfloLdA8+SNgwDtKVCQWWYBULyU61Te9egrIsGcHQcgnSD0szInmQ5O7ua5Fn8yU+
1k+Pb7JUJy7J1AZbayU2h/M5qNNU9iZO0k03oiaD6lGik+xUPmCMkfYML3fCb34HsAWdOU9/2AVJ
/KUyA2XSE1jKINX9mzBsjWuZENjTAd0t/B42Pg+qd6wAnvvvVf6E0Hmf+dcSBCAL5BPlTIYhcxht
64jhs7102bCGswWJaAsrXag3fFZy7CA2fafsBwLbWw+wAZTe5M5DTgrfLExWo6mO/ifBJEXG3aWU
tkm9FXCcCwbtlLXC74oRKTxB4a5faWtYfoGUAPhru+kErtX/FddQwmzsa2igcpO+HDHOyyPiqdtU
vUCyb0iI0ogQ/jpn9rMDWnlO7obB6V08DrKtyuzGWaj3tq/5N355L9NWINpi9FgK0nsLd3EUPmWY
gNHVVBGB9On1hi4B0L+gzc9G4Gwf1qBRAr8/7kJABuuQMAC7c3R8VNAlVcuf/XLESP9ykZsiDtaa
T3AmVN+M3EVp+iViUqVgHtcXoggLdD6EVHdAAHOxMtgJ/xgI1jGt+i+DpdlRQoQKDCCgRjVG9TpO
Nxq3FDaBAbXl5S4ei5c9TFn6X04boD2WLEnrxSF12kpN6puru7tglibT3ZNg4AGF2Xj9KhPPZybe
Yw8BAjZOo9Q5pBI+gVHaJjxroFVzWHg2YKOvlRoDY47En3Uyir5poagRFlpNQiegb3kDe8t/8MoL
HgJxb9tuNLTq8Ap6JClwrFxY1uPNPih8U4onxHH3IBc9ZxiudFbqkM+TwtcQGnITj3aBLl8hAaQE
SYR9RGUj3NWoTZ/EnF4Y9GeTUhaPofPXF930Ukp8QiH4bwUtc3jzlDWcA3YHwcU2a/3khMR2ocLh
QKh5FmTiuFwgEIS5Fm4AosK9L+UnoWgUAprwFK88Yph6ZDmOOYAtFmu2//AUd0mggiFvChzK+zew
PCt/IWtfzCILByOmLZ/H4RBWt4creMQYSwPKhjvAJoB7b828R7XjFXspklqm01/KBn+kbWHRyvWd
eo4zIAA6yCZ1chwPCp7nGTlN3HKarYM0U+wmpDfTpkiRzkz6it3ELv7ijp1We2iWErjUeojO+K2z
5WBMV+OGOb20ek96I5Tn8+VK2SSNmohG9K1j3vSbW5ghuMv5xVw8NbPbEGD5M7Tr6CteqE0kP09k
2qjyZ07eH0Q6g4+c0zrh0pnJTny8N/eAhCtPq9d0q6FYS+79WpV5jEarEID/c/mlOWYaWFIQWiCe
6trDlDOSvQykZgXghLTyhkLWGd9rBTQ9d7z/W5Fv4BPcGtSiiJ1mB34byk2vAiEbGlLcKv6J7FuW
P2pptQQIyMXziO2oRmI9Yzb7gu2l4LVBuMgoR6PPAr+gLecx+4KCZNempTuCSmJvebMou/t7Nr5a
Zan4yzbudetVt8aW3mQfXVhT3ZiqhGVxcEiX/OHKS/fg3svX13suCCP+AcuEdICbPaWQa8OETucy
5s1DOggHjj6tLaKC+0+s40+IqNsoMT1M+0qw6sNlPd8u0vRHGmHdgoJi+Sb0+mCIkncHx7dvEVEO
Tte9mnBwXf5BXRcfpCJc3TbrLqIjvx0KNL5lX1rHjA1hBpT3qmpItkeWt4XyRa3jGDauo3A9a0hf
bkYEo35ELo821fJydHQAZhXJodrTEgcDap6JeQ0CUMLLR6cDq21uSMwyvFfrw9u7WNBU+eH6OROF
8nZY/V5HJxicNeOkctxV+2mplm0yxmgeFLYJTcWfgCPG7AuP6CuhQlQxb6QXHWqfgedDCBBYmkvq
qLDnyrgpmFwaKEh1+7KkZZ3jK2/TLrAHWTNagq6VpJj0YE5aJxja6oUIrf1sJheCmSw7Davn4wcg
el6el1iL2bGZ+EfA3HozUPQAeupfcn48CuK4SWZhV+ClSFOKEzJqvU1SiK/kZwniPScp8g0YlXZr
qQRjcapkH680ItU76om67HyTEAw/psskTuO8DCRT+5BHz6VpbruAduG9r8TLuk8M/z92/uNq/S+r
sa/8rqEjp7kk0Idx++cxYWly9H8y0eezt6+vH8+Y2XgHs9+50L6CRLh38kx1BtSTbVbYxQ+MLexR
9meoENHa+BNgG0W8u98rSFMXNZIqRHdaJJ1sQcDY+Kan/d2+8gMadV3ktTZ1S7fFUWlVo3/DHw0j
43cYG3sPAgKzFNGdMZm8v70pLM5XxbRc6QoNnu+wRchQiokqox4tv3C5QW6WAif7bOL1Rf2WnCp6
f3jCEHR4tzwZrcTs3AYFYJwZzbjnPhOskNOVr54VsrNhasqEjhFKCx2vQcz40oW3U/c6VROKi+dr
u5t5xkKzInsqe809HRr99nIgCFqFosRf9G1zpC24vEVyLaLeflCxdpF2G8C2Qgy7XTEYNxRJdLfu
Bq8o2MSlzucjuH2YBv4SWupwBeEd4m+OtUk/OD+rhg/FNkX3RS9Or4w60s0/bnwsq5+mny5Qf2zz
7UeMMV6o67U/LfBCzkc7/mmHiKqY4nq2yh3DNeA4wP7Kq2L5YQnDz40LAe4H8G0saRJYAXiYaHG8
waKKowiriKgEtoD77ULk+Q/VeYRsoPGsy08sVmoOr093Qb1XbUo6+06BjI5EGxExNFy4LHt7AGBT
GwOylPoPngIHiFUgcxg8yC7KPXCczvKB40mrvJIkVo0fXSz5XygUrbC+e8sISlev9/h0w8JXYjvt
1rLDACgEYQje1+7N6nqjEaza5UJSlODbRyGEmxvZWp9ddJu2DL1imIMAghZ9pJhRqBs4cCz31nmA
ujQcqStLP9/RPLlTQ/4L49+cAQoWVUcIlV758O3cjR3C0hj2BuhcgmOyRTzbPQKAB4xxuM+LyRUk
JoKea9CaHVGCVwTuJBERm6RBWombpWqru9L2Ulq81kMALQXoBOKvPZZkod04VHsah0VKLNF/7Gfk
0sKJGFPScwQsHNpB7iEJ1CDRU/qbxFXTw33lklArBG/vs6MOLezA8m7zTYUx81SGG4odfC9ieviJ
HhJu+tc9NRQ/S6vLKM0xE2VtduJ+uD/mCBhLoznC1PYzzvrB382V8ZoDvVrrI/hRNDCFWIulE+wG
Gm6aXY0X+Z29L8lPAOYYmE993+qVNp/xMAC+qs3xOG1HjB/GCD0UVtt+i2KVBGnIXIfwV2Ea17O5
mlqGPM4FNorjbm5y9Yx9LwX+51qpvOgc/Xv0iUbky3UPTJJ8fV//Is3U0ZaytLc3zHt6f70aP+qM
et/7OxOipVr3H+aU68Xbv2qHBVkGStbmaAbNoznefI6UtJYvf5CY6aj+epMosNDkG6GIX6keg4yZ
kSu4Iv4mVrzkwP3D5Qm+WpFZHA7r5x7f0RHVhdxYGI8o4fbZ5zuWSD++MRtQ2uVuUsbzsGnL0njE
cgKIiu7W8TEa+xYwp3zvl+jdSQ7C9VRssNMwqNpbhW9aeH0Dj7FYlvTEPX/WRXAhl2fBR3aOfv5q
hHiVYWCKZs1A+PsSadXR4fAKrVe8Xi+inO9lnU2do8qbnZb3VgP/yJ6/+6vu+Q6c3HDCcEqJbt4X
4+IYtKnG+MdJO/cisVEAYRpDM4GWgJREOrWVb/s5Z+rDGZfIJI5SmlC/EQRqJFF8CEndi7aobA9T
5Z17LO4CodAi4I1+h7ahAXP4aubOlKQ3hxWdarVz+1PIh4qSvp3s10DHu0cGqUFoopvwaZnqEdIM
f+HVzY3jNKM72HjG0hBFQWD2XH8PxZPPZrfjt503ccptCl5abOrtHys+4fXGr8vN4dCy37dayNLh
BJNfCwkjpbv2D4aaPHaFAanXYvFyKt0huqaoldAj5Lekh/fIS9sPrbtLe8Bzi1Ioc3QB0Yof66Rf
fctNmY7Se+dS492EIlO/1u7/CL+ONihUk4bm5KKcb3zKzhvhDEBKzUNIhCy8DYNHrj+qonu0DKFA
arWLHQkyCHCHO1oh78V8V0EHMDon1lgW1YF9qI9KqnW8UAHW+pcuRtn0G73RUgMx3Ba+Af1EmdeG
sxCzHTdPsjm4qUHm3oXloaMa4PwlS0uD81ZMhYOl+SXgBF16lM3vOfB1RjNSl7PB70PDNA48hl1l
xI57Um87nGU0EY3vzGn7G8pORDFnRzw0oMOfcQXYEH3bSAHOKdDW0wTcEe8mM8rsRfIC72pXJcVx
b97I63V/j/q4b5oIN4ZfKWgGPhT5cjdzh5pZ36vFj4DT+PDlTNL6zLBG2CgJBhLpCPVWdK0ujlFk
DMJTC7LWVNz/mKV4LJzb80Usnm1sel1ezVlWxir7tSt5L31AbMdR7X/gRo6GhTML3xbxjZBE/PAD
i1eCdZFeBvIt4erVZ6lH4JY68nc4N4yvfWk8i1ceVy3p4KTrQyto6ublJ+tEIH3J36E/QiW0RMBi
z/sRP0925BPntoIJk8+y42op9zBp1UGN2pqAgEFq9ZrfhZo6tDedH2ejhGzE/9r8n0d+5ye9QhxV
2Lau8wiCRRs8Y1PfpAX9R4iiXzrNt80pGMztfwlFoZK5YeQ7/EEAswHjnb7mF9Gwe997HDHSsx0m
REjRfaxHFF+LwdW0X3WUA4zsdcqzLJYw0aSGwgThbHkeFo4d4sT+rbytxd9qnZ5+4wWovda1jkG6
dM5V9eElbdQOi2xz4qz8Ii5qal3987z9Hg4DmOsN4/kAYwf1R4jq7cgj5twFCJBqDw9aEgo9mlev
NUv/OXnfFD5rX45Wj0lpBe/Zzxpsd7IC3NaWykm6j9oapNOMWuE16U4gHsx4H3OGv3k9RRN9t6ku
CC46h0xLPDYwid3B+bP2xlXuwa7IQ2Q6HN4nabtYDNKH2loIwnMd2whEtI3L4a6JchRCDBr8KsPi
Lalsje04z1Y0YiLeOCyc9qVBRGo/cS5U3ldYBpuHsCa1jEBkr7ELVGFJrpqm0AsK/6Js1703Z3sh
f4qq3NKyXchdnAnM6RS8rBMAOb6Z9GlN6O1E2K+IgeJ2ajb4M1skaX3V4l9NoBkyITiMEcDycVRN
Fxo61yGtKYhj9mh09E4B0+UqihBdVppfSzR4NUj2eykbvDpFDT4LGeTMqnh0SKz4ZtE59TxNg6aJ
NUUcmv0Bie25grnEHm714bmbB1W275xO9Z8JFWdlRShe54tZGK0Ii/NFNKy6hDaWDHrKxiHRnSTV
iQrGqseTWYNgQv9Q6KkwpNjIPvYfHnnUu8IxKE3BYICqEXY8C1kA+D7moPBvsigqMTHvLZ7SKPNh
9z/U0C3F1rFIcuYfz60g9GbYMD/k8m91stb3XDXAY4T9TxPQ77r+qo5b2jlBjPhJanMO6CV7y7Mj
xAz23angtM0KeIBkjjDijqt49vR2X/Q2mDzgP2ybfe6kH/B2D0zuGXkFOkZNHLupF+/YYITi8hX7
XKBfz6/EWxEPPGJLQk0wPv3zeb0rUfSzDotkE7c7Xkuh9j+sSukZ7YYTfGsHnsytkFyxFO5e9s1J
rkND+im8XIVUXiqov52iT78tKIFWmbAf5efdI8kOOimVsF1RrlgSPFPZPVnqiV5NGmW1M/6JZbpI
IKn/J5LVV2BotS0kj/z2oxHNQ8gz5bnyPnfzOKBov30WcMxPUrZktAMcHjOFvQBIjOxkU+HUWsQB
XMaxq5jywLRSZsRCEBfsLyZ+n48l5moCf8gxP/HMMVivN2YMHU1KaIKxLqevynoF4szJDiw1Z8h1
B8BkFc1fUYerefk7iJBvgU/iE2Rye8cyI8jdph5ifzCfpQobAtipnBzYe516lFUMzG57K44wlCUd
wHjIJ2UYO+ERwwHga7o3VFvawEEtO6u9YeXm4I61pOj3vWeEr1P2AR1KyGPoJD/xg7LExJWS8xMh
LYhqXxbw9lmAODtmudyh5NFHdHCdqexTdflIo+vWMVLzlou55fzh98wDSnKQv3JuKuuDewJGwS0q
5Gzp414ffPF99BWjvrFFr52TAb8rTiMSQSRsdQqOuk53nK9rg0+YD+R91PYfKPzofYnSCMGDG8pG
o/JHbNuTJZ8tFfIV+YCmMkZOXsAz/fXMVw7MKBtHTlTXAMeJMDtJRRkkicywPtSRnSUTmB0fkUpV
BWcMk/5LJHduhf1BE3y9r+P+r0VlPkvYskM3twS9M9sfSn1PDmz8Gd5FEqfO2F16Yhwv2iLsEbtR
YQuMZchDE30/jrGuC/dHVsV/N+JIJQ/wHB+B7Cvu21QS9ZhyuDq5mN6V8k+L8122DA7yunYiv7QD
zylVWvqv30YhMqzTtyv9buEMakuhf3dXHz6qX0kj+WUvYogb+KhaqCoq9X1EvrV5haYDrEWYR5Tm
5ZEZd1O+gHio95V/xcHiTh5SGK4iRUxvha6PKtidI8CaJXebVT5gV2dbIc22M/72Jxa1RvS7uY2D
A2fIQXPkZyBrpyY2NAxygvSBQ3wlQdaGn88Nd4Q7Zjt66jeOI+ZmNp/hO39O8u2/bt9dz/DbffwN
T29/kosAkitPJgT3KNBOSicsXSXqku+SFBceTrvV9gL/0rjSQTD0GkcehKNEpOcX3TWP4bErjftS
jnWtnohUXvAvBjMYvEbGv5vubypVtSTYj4kP5MN6SusxISgZgZRdRY9ukQzrSMCaJN5af9L0CamG
ZxN4JCQ50KiEcCQjzxWzWONaGGrXkVVyYNbWNRWKolg2PGFUc/7zWvD5ZldBwFnLpSYkenujg1ut
Wo2LcnKVCHI2RZNB2bVh0KB1mLAf2yl6F3f/vsBvgdy6IO/PJtwOwxpG5nyBN2TLN7Py4w4PBw5K
QR3Hfz9YUsUuPagpL0igQHS89lWFTqBv2cP2NoZglpLYNzmSm9CwthhFtl0mDiNUVQPUtQlpI4sL
jCP71Gcf0w15QMBaFEvGM8+IpVQKJ4jrJ3OTrInuCDC1IlKif7EuQR45nWn2bFkb42e+8FUH5KGu
3dCIHU2e+K3ESlxINmtw97F2Hi0SH/xSme2cBomdUnZJr0TQERZ6jMZ4S+X+YKcBp+jvts9gJKw9
KHVL9f6SFbLg+UxGSibXLCqCQqb0g2Gq7u7wcB/lzoiinNFmxOK0HbRTMCNVbNsK8emYqJCVi+FK
ARKavKBWDMU/SlvpPrrTA/9WItkQfjTp1LfS0q6wIArHtG1QKqO/Z3qJ+FZhwP0R+TPTNXBQXLUO
mrHz6GCMT9RhW1FBst85+/DGrWxsouHEBHDjDzOCBCjKPMy9zNEX2VNUKe/NVX8+TI8NkaSAlxsv
i+UVaorraIrzu9UaajK4sVaUmZETxhnsio8IsfagFRNQcT9DZY+d329jyLGs8tCxpwoNMylSF2gO
zQd17dR3QX56xEHf9FUPUCJ1AYNVxNJuLMDIwfxq2W2NVsuL/BGCD1a+WetNU4PWEFtmgobD2X7a
w9Qs5ugPzbGQTc4quMV9eyyqIV3R/93dLqv88ice6PkHCA+IaFd/sdo6JNy9NV8UbMVLTstQ0kZA
dJ/1Iv7uit6hBlOTamnExpzzg1lhsHLjrndripVP6qVuN7j9qhdx4HTIqLIQqGQDxZt6mOqDhSJx
JSqbGqgTQvGZBDoiTHe/EBdyI6uW0AWpghnVMG8aN/ir7v7xC8x4Ci1jYzlMDclnGHdu0TsHZYV0
3xc2zvsvfqCKu8ZlkahH+2yILZZusdnthODfpODqCidD3gPxcPGjjrXFFbaQXu8D3tXYJPY1Ez8c
Ec2S/p4DQzfPWqkAfIxLvITv+HhhAjdKraA2z8CQi/1npcLB/qKOxekQuC5T0nb98rAaDbQgcpOZ
advy6bMOaZCzdmQNlUval2WE1iSniPQ/WGZlxEmZTnFWCmtsUZeT6+kfrOTUYRIp1RuR7LilzW6u
vNdg4lLmwlsETDJH0LlRntaEFTieXH2psdNX/FCe6x0HDnZ4Yx+dpsUFCOOYzh/iRpEGLSrpQbAK
kLFk20CN6FVhKcyb5fLoJ90IZQcEH3TF/Dn2EAEuEdxsEP/ka3cjUC7VmYAWmXJEAicfXqoYkRpt
IBVkjL4AuAJd115UJRPFpZlnsjKyJTgH78Lo408HC5Vitel8G8K6ntZ32rLMy7eDGeWTrZKFZQy8
KtULOPbEA0BLDGDQZO9dL8Zgb9DrhTOC307QTAN8knUE/ug87xNQxyNTUX7Xal+x54+3P1JXff5I
gGWrf4EgCFivpK21grcRuwq3+8GjmIRrr7FarYdEvm1eELhmJzUNKnYPYYEQlyvtZ8/xu8AZ8jam
EluLx5tWoSkLVswZgrojexSjkNKlaTJKmcTs09XExKblBwvy8jIWoX//kDFLrzmZ9mGOhSgKYDQD
ixKMrFpTYHnlyju667fHjtvUzabV/xeDYque1ijftk6qq05kaQ8Sq1HO6Y0F5Yx8bixCZP9M0GuV
Tx2yFqTBBSY6sCGkWc2GqnpoKfqnt9b7B3WmgbZxI7N2NJtrpuck6xPBnjvvRTUeyX7ygUc+InvU
hI0sBaCHYRpAcTYrQZ2w3xTyhWcTir6WWGHavRBrl1PTfFoj7zygWW3ElogstOxz31fkHSMMn2tq
GX0iqBpQ2wNshZUOuxFDCifOA5do9dhZNlTWSatCiZqrcdRuTi/xaWcfvGItKK1NgbZUapFLstl4
eFvOOXThat78cmO0Bp1xiNAbQtGl7qwOllvzJdsM+L9AFyeL41g2VeEaAhh8MTq/tP8ChD1YJcBH
tgsQ3OrAvXrYtn0l2T8JUvRtmeUggXINDqVcGTuPY3Ft6GxyxyJyycgniANrTHG7dC7RybZgZ7CL
4pnf3KZ5EF4NRMjqKe7L9YlNJdycxROVCE4q5W8SAH4fs5Ob0fmf4hu9Rc0uaEinA6qH/GukO2Ui
x/K3xToCGTq5gFv3NoaZ+zSgfnD4Xh37JPWEpnCWluNNXfgycomF/YADXTSDz4OEcBovh9tHNEb6
1BlQyH3Aj+OcqeqHEFCilt5H0bqrY+YL+l1BqFqXjsCs53DoyggoTUtmcFYK/AYpH8jJHTs2v7JH
W3OMbeJggaO8Kq4LRFfcrn/DowkzvSg/7H/3BLdrNHAoWyf8Kdpm3Ea4TkVsQtOMrhCi8615rhgw
7qunUftvgV55QsFgmfO5UwjhVbDaTjOb7DJkHEHYgbmycjcbBSBBHeAWTFjd1Jwsoc8l+8FiCiNH
g3E2g5a8DqwmgYlzYa583J/2IJ59qfvHW7ikfzeNi5m+WMaHuGhhMwlGX6ftwlXzWuE06PCYNRQL
9k/HqRwfMLNxQuR89Up3IPH8j7KnNPa1fVGOdKR28AjnKewTjctTI2/vrHKB0mttRebReIyy6+DA
qJW4nCWQxNOk3W8DrFBq1VCHtcqLwefUHojveULUF+jYvyQogTeTGzsRMLU0Ua8OjkeDI2JoNotL
kG3U5q6yeqMNiZItpbM7S+r3JMSdCauNSZWJIbPbCDOo9XnRx2fmHzPg8IlE5aJiF3NpSOLhKMjJ
ahGa+83bO8sOm+KkO8DGGqn+L0plTtxBPAeKwD8ari2dXXjCZKPLBqKAVretb4Zse0ywD4kWAjBp
iL42hBxmo3FhLpyUcx/K856wSrRXSf17cF2AfBLBO+cBS9Ze2VEPwDgG6gqiKr8BOe3maRwi5yMr
0mi2d7SdFMEdrpS9HpOkAhkGlvz/4FINy5BQjNXH2DAS8jzu9n4TRfFm8Z5n4rpo8v1x7t82ac49
lpS9xIdKccE7RXJw0dTkBrvVGtbOTRfg2/r+RsASmlhQw6DDn2FBVdwcVYdhfChWr9WSMdwIJztH
hb2Jm3t051AtsVcNYj7Ro5psKEobZx1HLc9CF4XhTR5J0CYeLA8PSEhBhfTb4gvHok23XqnZfZQ6
zUOCnO5rX4Qk4Flk8QitL8CJPcD7IZahm0pcxBVIqFADnZu4X2Dc9IgjLWqr5DKNiSXufW75KO5S
NltVt35paTyt3zQ9dkF4CaYDa1CFi5NMyuvIcdqVW8CjZdtuKe2UoPd5Cj+7BpA9fCIzBryx3gCg
XI4MHRIq+RATgsUE8pgcuf8MXr825tpy+IqluKfCmVAvWPLX7c3gKI9MK2Gks7rDaHk8X2zEcm1J
gcsnaCZYuDN8NZOXFehwf41a7nZ/5stcrcEsXeJpE8DxT74e625p1esp17lDQ1jP3+lhz0WMesNg
zVQUAX+l1PeA7aCZLeWK8DkGabYjSI+4pWNGd+PrIGXS0qoLLc1FX3APYiMUaINfEMLb/wEMH8Hd
EPB5bVpLy2s3ynRrMaqSma7Pi89ZRXHjk6TozhJWWMGA0faoKpcCc9MLhtffn9+XFLC8X7dV3ojg
osxSWT/Vi/sbstO/Hn94hohIP70s5e8O3y8ErFrm9FzDnyOU9p0MoHqj30g4Zn36RsAwDKGnZ3/T
P4ViO4LEamYmBOt9rBuY21phWXDBPWNNiKxytb7EfgZenwYs1vR6AQ5F+y1sfKzpg3qKtfoCU5G1
u0QDoz3DNHUL4w9naPfozSudGwuv8S0xUiALTK+OBTNklY863VKwryKAocGexWkJ7Z4PRVvibR39
YmFwENHd/yYjMFDhFASUwjUKsDHElOHU4lrSskVZngYzcebrGMArb5ZdEnoDK/0QLf19Ttl9f6YG
WV8UndW7St3zi3pCnPNC6vd6H5zRGapLjO9qUnSktdObn9BVE+lOtCHZruodrEDBpbdR/R19XsMz
Guf8TrbUcTn5YKyePd/A0SN5NaEd4VWcyfGrZRhOeX18aocFgfcF8+VOcoR+zKqsKJpWgTEYIKOE
zpecgZhLPaR3+7hEWdKHL8jtLVsuf9zlIAQNX0wN9WpcF6qknsWdPKU9x3GnaB8vrHjBWCW9dpZJ
uS8qmFaL8VNGBgPlAlO68P4Ya2BfHE+r2kYMq/8iSD88TJWi8z7IniAfv3CEXS8P3vFFX2jeSk1l
ih8PYDeEcgdnRnb4WBZ4noePbRlrLPiEsOL6pxbroSQq6bVX7e44pNCe7iKF0GZJ01TwvtqXhIQB
Wj8PNuteKKwJKd4ct2Kfsqq6PFRUBvN02pmlbiy4ewPO43oVIinVu/lv/tCKbXGQYLaHDSY/5e4P
CgX757uvsrvGYaMHK/K/KQUHJMAt7sFH3mOEVKlFKeRx6jy/Lcc1DPTNiFuCgvFqFe1zrkhkQZsK
DSYKnFHYit3LGGT6zp4S+2GWyLrvmVDEulyrgdb0lRV0LUKW4vMuhRvXaHhxzIDk06eD87CJdXjT
WUXdvtCpCc9eFc5visX2NYOwP83wDitxbrhPQ6/1LQ4GhJQHYEbzw+S2Czl8M9Fh5KaUfF4nPdN5
b5ZPRkJDYBuYyIgJ7FDZjrmyqvKiyD8VSSGGssarIgsLp9FVdoPEZULw1REq/U46gJmB6JxahlVT
zY9dkqURbsb/8mq7EpPfxJuAg8byKbxq8iysQ3IsntoqXrkNHgeOLhl29lq45B7uI3xjTgP1+da3
kNhEUQ5JPIRhQIOLlGSUFtzR05HnNsfgnlGUBW/Uq8bT471/7zsyXz2d4j5+c94Yle/3fExauQMv
FObpd4AeCyHV4m4oSO17wt9yhCgTF1zVa2+LHFsWwKuzaT8MDpErc3KTB05QmFi91qTgkh5Cid/c
0SMLvOaL5tLrV15Bq1U4ovzLD8glY0CNcOUS+QfReiIDbGNHNjQkGNKuBYdbsUNAQVg9Ve0h/u9t
cDFvsAHoK2fNtAu68RRiWFLYjHKM0iXY75kjA77K+60sS0HH+JpEN8GnnJrcJq4Gt9Yu9NC4XwU0
5Z/ZrWePc1X4p/XjFoO4NiK5wd/vlP2xQsQMWMSWQmse3W98SXoEwGbldMXbD6b2E0GmoO5MGGAt
IBBQbgN3TYSFQgDj9XLUtEOZX5fIcEq0czTt1sPb1F16LmWAABe6b4N4qskVUSZBj5QmzCph8Wev
Ll0v1ssQx/OlRdll9jVgYML8d4syvt9l5gvg89aWzhD+U6MN54QruhJBCK4h+XeRpBMQ0c09/MMO
wNzi/YX7LjuyaWAyDbgC0A9koRnILXZAvQ0xp4BFzu+3+xxJF53Vf7CmimFVdsmhphNVzzUy8XPv
PqJVAD+DrIy1IZZpLmZH7eNlOOfDtM9QnjpJ/t+qAjM53IDGcSNh8k39tqI++ZrlRa/9uRIhM7S4
UcOoejsUI72V/waO81JZVqxeHmr8gYAfmDSkEIRSjXgFyOUs87t7PEU9NJeP9K0u+Yn/f1Il5ocp
nFQyL0bPkK5lDrpXo83+IWC/pg3/sCbcphbIlY8CUD1138zndjBaiFCH3Yd6iMJztKvxcZWWP71E
BssRtl9gCSrjMux99X6dfPSO2PhSYGxh0jacEc3xHZDpRIaEStU3GSyw047YLQkKYMAAH0C8Qu5n
Itqa49xAYd02VeXgKmDnFS2Jv6yIjp6GavSJzF0uCGYmSzLOrG+YT8xnHNcLiXiTGrMw3rRZ/mIT
LEiCKv7in8t8amUbnq+m9S9nRN5rkWJa5FCTMfxYZA2E9oH1KYsOd8lYN9VeszgPwt9hb5XewnO6
xayYAk6296xeCOezIEOmekIsY5/grpnBgkKm5G/UzmKWaGDPM2m4VX5N09YRpx/OAQ8poQcyY+4+
j1Rx1GJ7OXd6LJoXuIs1YDxEltnTQ1DeCDcGHIt5Pkly7qgXqDijZQ9uGM7SdxxfB9ha8RfQecBP
E3kZpflhKBMG/g5Tk54waNpgITj7KEtZ4R3HbVSBewDDUOImDTyRLuCfFSbt/8sOjbkP29eYwBvc
VES8sTlfx43ZtHfytrWN4lv3c2HvuMhr5nCscP/IuANUM+VpgFXhlJvV7j4CKGR2hsYldndpLW7t
45c2wpMHnt65aPQKJ5v5pdKP252Ag5loBUhv4DAcR1Td0v0YxfPgFbe9WRlHSD2YeOlPYejVt8D8
RC8byLbYFpSHOyK0P/ix+KnAnM+1RKlmmqhiXA8JJ9833nwEUOXu1kv2Sv9q4bUBfIUD4kVJdVEZ
GgM1/duxgb5fjMeIklTfir1TF5X9T3Ej3rTFDuodFQ8RgCHSlPp+Qp9a7A8fAeZhshjMcHCmVBLk
BJmszZLgj81rGH78QmSKGAhE9ugixl99YNqds3sas2Azolh9elFWWIIfznrx8bxlcZLh4+oLUHiA
S/ME8kSPP34gPHKiAy0Oku/DSC8slHChWSxoxLe+1zhDBFFOd1hUJTplLMyVl+SlR3wEfQQJCs3a
hRxnQyKu1ZAqPJZaRE7EJUEcmiBnEtJcNDnBEeFKfcraggdsUgjpaOZtgSNwQH9mP+yI7dOmUhTV
m2oLGO7L+jQv4MNineuVuR0eGwedcQGux9ZFlOif8PcF0nrjQYSAsp/UZplxjl/jPTT73IedJ7HA
mZKxAt8Qx/OpnhBJzYtWOK4rU6CePNWCveO1qNNNqYmQEX6BbeIbQw2/ew0eTx3FuDv9J9I5FowJ
keQ6jBrR/4rjmtrwpI5QDaCu3CdIX1hsVatN5dT5qOSo2lKCRE3m3aMyqtRpHJsyCtmLMwnIUAFn
mBLiifvajonHEv3lfrWej3qdl6tNgGzD/gRHr7e/afmiFao4eOEJswcSo28t3YH5JQotZPscWICH
EnqysP88YZJwc1eo9qStL90WLHRkvloJ0dKxtAoy+IROnNti/UCqUvwxWOkyb412/egVsGtmejyJ
uKj4X3ayOTPY8r3/l7YmfwbG38LM/lfudAMb+cY94pskQpOIOWnmGtx81RdWnak1xRcHaZ2OdUU+
MNxul5qBHrYFnaSSQQog9ez2EBg7qPD/1Cmdpn4y14pODn/ZpL/K2uh/WMTF4Pi5SYUFhJ8V8O5l
4jlPdrdduxux3/VG9CFBzagQD+aKkPRtMGEAvoz6dNcIthfgdxLDnGjy4qR+6C8Q6j/KF7arV+mr
Ny5dCm8xopn61aUJ9MH89f13/d8/Yo0EV0pc3lmJD3pLulN5gVlDVm+SLBllDQ1wBzvVI59mdzCq
UrqJH+jjPzqJXpkL0QnlugBJ3XQn5DZpbkxfmIjZTY5XUHIG3DyYPdP+BMf2rdPAUBKXP6ongKeH
DAvep3DKgCRzLOMWt/YltaH1F0EhKIgrv/EYAqnkY/nUvyCKDsvZZ1Te82r4VhN5VXJmrfMwEvYm
gTmgPDgtmPlrV5m/64D4+HQoGbgC8BdLIA0VRRO9SU485m4hcSNJPpC42i5tz9QPvdUkoVAUzALy
Nv1yCdJW95GHk0RzSPiJqt2vCyM4cGRfgJCxJwLlk8WYlt8a1sirr1LDfCJPKNz1WO4F0nWlQ4m1
oNGnTr/MWwsc9dbqH37ye8gIJgiX93KXmvNacfQvpAYTxZ4XjEoxkP71HvtmQYZhrLGjSiC8Q3Ht
zocWhbhwJ6WAgTAfFhd4h3f6qCMtSCBmOJFzkrAhL+lFOu6WW/XNMhAPelXioZ8k3CqlM5iIeq1U
9BatmzUBQBirX9nA9Byy48bBslPzttgNr7jYg+J5MRlBI5XIMolHqsykqk9zQrR9YQuG4nhqbKGT
iY26Qe/IiI5zxAPl2leiyiicpocF5erYye8Dom8IC+QjuNrEAKa5QBl9S9Ci/Ka5NvlwyBv0ouRh
0LEObyWNI+ReowDsyVKfHZWwM2/aaEgih8cLUY92Xo5yDxhhAlHw1YhgQYfHvdYEOvk2hxunIeYi
z77cS5bVyjsI2jrgomTI7sP3dRRNMAmIeC1X7Dmg5IcDybkp8GCxcAUHDKqtbYbEyaqcW0UAqYou
aYrJWPTg95PrDbI58fG5d2bx/iTquQPBO9BbGDee0zq5+CAQQ0PcwG9PmYyNVFq3jB9Ca7Cf9i1p
RXzusF1gpeqWBXjJA3v0G3mdb9Pzja0mCiukI6lWBvLD/KBJp7vn12AdpMO23l/2koMDwYj7b+0i
LsTqfRfnLHdj7/4ooNPk6JIqvYzhZ4IRvvARf/wgf+Hpr41dzqSw7nAH0iY4ldfLF/YF822bd/9I
42eAZRcPSQFbstb8gYj8IHovzb7dtSL0N+2co8YTNUrMWncJtDInvaOVw4Gxj51o6owlm+GaIIqN
QG7R6d928IRCtm0nd1Y/IZEGQZt0yLU6aNf/nWWhol8VtEkOx+vOrHj0xFy+4nw9oon7iSvj4l6w
eL2hSQ/Rmg3u3u3GYN8QoP4mZBEFhALZ5j1M334jslbi5Ip+eDCmUaGluLdxfH96m7x5DuDo5mrq
3KTBL58ob72KPCbnmJqk2db8BYYXV9mo2gg7kAewOfdE8wQA8srLybKTEZoY
`protect end_protected

