

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
VHfaMJ2jDU0R2eAkOntfC5B4/6MobpZ0NSnc7trviKzQU5KHakm896MNUQ/U/XUDUOQl1Ix9hEug
uFcdFGHOlA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
jZ28dq+cqatvP/oWT0j+kbhevax+rcvgcOVET6FHORIxsClPAe5EiSXk6mDgtoieHOJgnr3iO4zI
pViSw9QXhHwC7nkjQzCL5GNnIAYREubhi50JKwxrsTofbyKzT/U5b+jDP0girnK+nPIjwrQv3vvD
PHropUlOeQU1eg5rEJo=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
wyTaR+5BBK3PMm+GuCvq0Bco7y5f/oiFqNMyoEJ+yA7qA21Rc24sV0Xv3v9W4doHSIdeeP0oUNh7
9I5Dbu7bsdY24p4a6rVQlpW5VOJjg7abnoTszev3jaBtBOpAM+FQDIkOj6hl9ZK+eUTOGH08ap1P
3rtu9S06fVXB15p5GUL4qJ+pbX9as7bXZJVw8JMDVFn1WsdJ/zMn5PNvL5qC5jZb/F7Sf9m7DkwY
x8I3vpZz7RsD6/RmMhT4lv1FkcH4MpJegB1J0hL5KoGG72FOKCqONCLsZdmnqz5BmJzgYmphlYZC
jJckdSX4yOLEg+jbosSObzMclIjrm9gORAOhKg==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
qekQcsRlt2+SE3/eW9XQwKmx/wWWvcG3c3jSLvuGiy4GIetXM6PaXqKAuGTMI8b+mux4A6dEdodI
mIX5ojnf5ZA1jyISA9q0jKtn/LDbiV/JtKzm0pK23fPqh9/IUaTz+oirXN82WQzZFKQ5TKpwrFn6
ZmImSJcOKVgUcM/iG2U=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
tlEZl/v6lEdJp5aVMLYyANJmLh8DNrpNnDhyEkIUHbeTfiozIDqQ3eefGpJHd1yUjxDr+M7d69UI
c7u5loKJo9CP6qAEjMhB9NE50dWkO/cRVvdlBQSlpGD8Asrd28oTNAHTTge+6t1TRCmYfvMKOt+b
zBqmGPTyIDG3LI8DiLXNfUjWjl16n5IRikeD/e8FsFJjAF/a0Kjal/N8CzCmRiQPdsZhdMiruSdi
vpIRkNPRNpCK4J6asTfuTemt2JkEkG10IvEYhZ/qTCco9PECc5G9y0loOf9owc6R54o3iALi9D4Q
T0iTW1tROVF1jLbRTIe753z7r02QD4PyC+02yQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 24176)
`protect data_block
K+EmP8xpURQwFnIn4VV2qIQ6j2PiN12d7IwIgEKnqSqHz9Daf6T9ovzfaDgImeF2Cv7/Qu/67bXO
Eo1gaINIzo3AyHtb3N+UaOXQCPLi53V1Li8pnRowGcXOw7LnI9w09/c/a1Le3ynd9qnhD/o0IcKx
qXuyK2wnb611uMbqYKeXgdLNf0MvVI4r/qb069IhqQUillUZ4IugPZwBlI9iUF9TJvPDVo+Haw9A
T2u2Uumbd9inLYHyHknbuz+K29HwGobh6/7klpb7RCDd9nvOBfhnxK+oNK910q2MC7xHWlBJpybE
k7/qw9KaQK42gSLZ7w+29odKR89S5WQe01fxgKIPdmLLs8fPYSjyRPOXWOuL2pAkmOFZbxXnDmkg
qNNFUjyRBBbmBvdDPj21KZykEmZt4px16GA34lwEUU01AZStYk+zj6LpIPd55FweKIn1scjEtIcS
+5Z6yaZ/XHfGOuhFk68Ekt1fp/A/T4yZCcI0bfP09ptJcJQIW4zoaFBng6wEwRVOo/rBdntV0neg
dA+mttlPxxZQI1XIjt9zjZNnapUbmKIO07O8WOal71Crixw6D1H8JE9jEWVxw53BgaaUQFpop62G
C2lzJ4k2nip3pekydoBzsND6lHAD2twe8KY1ucPWtDYl8wteDIwQ0OXhhXbRXsgDH17uUr9NoIrU
iK45FLAi5JRBoVC6Jk1+1YvLLQTQXCTbXFdVuJPKiK4OY6evb5yLAhiwr1W4krmf0lEFWXmDGEok
Kz99v8d/KCa9HzKmm3XzDKZy1o02DJibyNRLGcRW1L6ySWSTSHOhJaEbWipjYnjxJUchr79ksv3f
1yvKlor/tUfuwLdM9yxI0czdpsjKxtRFwZC3dcBgLHyN98Y2uzwlSQtfSYPyPX1G7afPJaDFa/RO
6QCnMTTdw02hMGQF5nbomQL+yZnM5V2tFHx+RLLYsp2rX37t+6yNEvCgLEoEmsK2bcS1GypAprqc
xNEaMrCaOS0bt9nm9blmHKwCubOavrKqX+dYm+q/V8lsl7k+BTB4ht0oFqMY69anD/EfoCmtPFp1
Y5wkejBwZmR7IPbqxIZ3ZGIzeWZwuWbyC068IC+K7myRJXt3apq/1YXG13BLOlozlKL8+BpP/Z3P
B31U5s8Ffvh7nT2nba5XJkUJ0bPrYk/FrGVRI90BktpxHIoLMqwixe3YrbHDZgxTOF2o0U/k4YSB
Q+5mHt9TOb148jdXN+BP0tXyqwcZM9GtSZ4Tku6yDUSbrHWM4+Po2ebS7BhULkkrsWFe3qUpPaFT
2gIFXBR0l2lzm0XXL4zr4k8S8fIfCeSQUi+mRnfyG4Cfm4olQvjG91X6ZGOB/o6WWdOD762tVEej
+PP+cr/LC1Cwjkb9Q5Utk439jj1X/wD0l/qYNAKCMWTbAr6gN4+TOdAHX/lUuKJ1Ih9K5V7FkBor
eHMf4mtbc4T7HGbB0FiT3LrGfG6dTcMFpWk7zIFjc/COY96vJ2JfPmBOwxsJiFBLCI9OY1DNUrfQ
3Ph6nsFoRTm3JXiZYqxzsuaHOV2jmbFeZCzhvC2EV4ya0izdXTpOMkLfdh8d+OVHkoaRrBqzuYms
4oZtvujHeXuO01K+BS1KrxRAxTHBvtoqcg9Rg+fhJWTzo+9omramAsSHJfX/KYzxlS1pvzmmcaEC
F2uwCWxtvpSvJeeFoSXKGclNhoCPyAf6VvELqsdV1jrbEt0U4ta0Vfwv38WBzZm11P7bPsARoc+A
7ruJ1Hpn9cfF4KRgBNtuLthIvgMFlqR+dEW+GpE2cLeFvvVShMfqRF9+FT7Ny3ONdJXxKSknvSgW
rMVFba+1GsQ8UqG3dCc+QwsGp+NimhFL1Zsw2s/zZ0AJIngqcDjFNw0R0pzFED99nlTP4yM2Jj1g
UAmsDHHlPqlFB/lrltqXfObJ99MThPOxGsmtGEdf5nqcS9CpRoh2VxxDQvDuQRU2Z02Op2N5J5Y3
SGkr1oVL3O97qN1UPSXDWUsi1Dk74q9tfPB89IQDvoLOorUkYQcxe7PLA7u1kT6alPuNRtZ4zQj0
lUXTYXvEozQfRcLHmz1AFd1cQDbfMAJVT5u5GA49rclr7R4lBCRF3TsqcmPVMgUTVj/tqLREL94I
bW/CZ7R9h/YPq9UIWNI42nO22MDdo2PuV1xjry1YXzovAnlbZd8tBQIYraOkUcs+ItVZSlklgOUX
IqP5lccgrhAJOolHgVXlsUtfhMS31x5ts5Dzc9mf5Szq0ns2pgFW0m6KgSZ+TjdQVy4benkjLMMJ
xxfFJgVA8rDs4zRy9TpiVA84rZgm040WQVbrryaMRHp7WHF+l663BAfTdcBEmvdZ1dlYTyBgwFHQ
YYcH5/PRPQQ8QJ2XB2EsPOEwo8VUI1J/pUKAlwHD18ckSwGMEDxMY0hJZEUqhn2BPq9iiKQRWfpi
IQSoeDbF0bWKv7s1t+175lK0uDYXGtzAra5sNruvvRSupw9MC2sb42SzxG7ao2LrVR/KxIFpd742
qpYPYJIGHvCacja0CGtpUirgc6eTVf7m6f0JAzSJ7UUdGIxm7bIregpmSKBDZPNK1AvdMZ3dIxot
EevGsp40n1MdfEK+IPkqwRCfQ/T5bLHvD74e7j9G/kt9qYvGNDm19+VT+qYE9QU6GYSsCV8ypgih
8v8aX2zRgr+yFZs/gA2I5RYNxFF93oVbDfuFmhO3eJdn66oLpNVdXZxSLFwBNGH0Yp4EDCc9uRq4
R2qhHhcmFG8p9xE0JPpgz2+IBmOWeGUDSbxRROsmJIOfubbYSJLOOTiX1lDmZ2umFUm8wzEmAeWD
kYE2HUKauxN+bQUVjX9TSNrq01PKLv3iDmcmJKaSBd8XD8bFjglPE++8ItanvalKjc/BhdOJ3foF
j1/D3/zn/ELo2VWtkIAKGmgH789sfQyCFbJNjlQy1zn6nfviqWfdnleqK+F3fMAv0tazexHJl+H4
cMqo9O+cjSFQVvGw5jxMbxdNPvvj3699rVv+U/Xe4lb+B4PlsgHmIpVowj+zQCpSvBv46ZhYA62l
4JlVA+c7B8hFfAQ16Mzyb3eZalCytkqnCzy3vr5j6zFeYOvhejxVexuvfUaCVaZSl8D3evebz/Yh
QFXpgNVQXu+6aAkqlUdxJZxjt88sdBvufLCKn+Jz5qMABTU3qmfw/xzQRaXHYSb3kAOm8mwll2mP
BvXg/b8dSams6dXYHO7n6NZy2xL3MA2x2NvIQf8OfgB4gSocUNBBdyoOikZ9XCUZpEhIDAT/Hx3H
R+7uq1GZmi7+q0sv2TiaVPZ4JcMdpLzt6WZ8uTmHZaXd4JYvxPZfxccXFoiJjobcjcKXbpboWorl
PwIfqL3H2WtVqtZ9jfavu/ieozrInfyG9J409Et2xJ8NSqm/YWPd7kd1O95fxIu/bDBd5F7BPD/9
OT8bhq1F6HnfFJW0MM293r0P9oouSymmlApMuZGbrR5ZHAISFvPNdCRr2/ld8iAUIiLZx0o6zQyF
GKqbP2e1X1hDHclVUFyqoX5aSB6QWFEuCHFmWXjZGSAkbyJyT9zGiyoxXkrEmaYGCMwurbRDGxRx
Qiz86lNHSBS4kgOklJ0d5BQ7gzYPy8NDNN2RrbSqn0R4cXF0ztxV85Fl0H7/o5TZiBmLS7NaW6Ph
HccCA8P8qVznpHLT1jkpdW7aUBgYPHwb2ZEhqQStN9A4GqIA1uxUTG/W+SSdbNh66DDVwM9oRT/V
vEUzxsG4JfoYmv9pZASlrIhie6CYmdKPdEAORQ2CJ4Ch73o1Q8y69cXju4ElKOi8Y/O0wt+2+kJG
HX8zStl5oP1mIbEtgPp2vI68NtIJmLmyr994ddUdQsvIwtlavWt/+VCFCIzraKbEH980Nh3jM1Rt
gZ8UDXJeYSMcbuXixvxJhDrKY91+Q6YzA+6hH/Lqsd5LqAsefVPDk6skvbPU4Dp5PL/1nbvwZd4v
0FJcdWCBMf1RawDg1trd5msxo1vju9J5npRwZV6ff6in8cdMLcw9co73YYfi0rwbnXE5VKKzJOeb
fSYD6/42wN12PFhFheYNbgUfp1ojwDiZIKvhGQc4vr4pp4/hckdVmwVcTMViyjhK4B8yPh+yOaAk
HIbOqKGHRZOSiST8G8Lbm7NAisC+TZGD1jBhsIXGbZNtTx53y+P2wTPcN+4pwXkH9390OCa7QsGm
V6VJbRneIXLhsuOPulmi+UHS80ioYTfLZfdIVydG1lGnq+1uyQQMb2EbrAz7FDgs1I510MbH/lcA
g3n2vhVDiNI0r53TWqbxFQSqt5RyGzHO25tQEMYyRIxKSjlIhBxXNwD7ygX+p5CvgFKQpJgM60pr
hnb3KwR1SnJKHY+bI/J4RyDQm+dRwJfpM0V7oVtiqFOAQJroDb5QB53FOHFj1+ew9QCaH96nNdXc
g65dAT28oDDZZ7+4M44FzyGEiVHI2H8AQEsQ2lA68KK8750Bo+kW5nqz8p6w6yJMSZmMM3oWsWv+
KmhxCwj5jE2Vr98uUc77QxZDgIn6ieQlR/s6G+VJGWGFKI633JP51C0JxRQUPzWSkKl4ACGE9fM3
/s7c43qwXJEvG0BAtulaLz4LTiempX7Al6URqJQowSc6ZZUgCXuUURJu5ROfaF0YqNzevuOtoyqi
thMHApA1rMYjZUwx+mApNyyltCKgfqFEUWHVOImWz8rhFdxziqcEbRkhg2E8V8Plb0cfVxuXI01K
12gYtLUD6gc1SQy6vOxDBguJKaoO/fKJqik4z85nxurud0SL9vKbofU/r91czfhmrFby2f1knL/Q
EzyZazvSZLbypKkisNLerihVkh8XeEWOnMNtrYA0rvW2tqSW93jEUAGi8C1/j7k2E8CKkqZqqg45
MAiEadi31TTuMKQz86faO7vR202QAJ0TX2EGw/TDRFF8ac+CzDGX8QJgM0qVubs7C9AageKA33yz
ul2PzKiWbDfPwYRvgwGdAqjTE7j2BgXc/8MYoMAJXWTWK5w0UEhAoilzh7ONKx4rtjKev64C34DD
wjOThs65kRqV+mwdKV0WnXjLihSLW8i3wZ1bo2voGrTpx67TBenXi357pXkutnfaSQ+NuSwqlRJC
UBu6oJ6Q1mh4nBouuv2XrjqcJEwscs/WQ5IziWJnTrYx9wt10s165M+jyMPiuTzWcsD7pb1DgrwQ
bSTkQ7TpPAPpvsaY1EVMOfWQu2/i2Qdvo+/HLhLMv06iTRaTJbOoU6PbtSWrPZYcMraBp3Iy9/uN
J27wLImraLdPHYH/njpp+0AEwGxJDIO27FarYox2vxyHhygM3YDfBmPX5eAdsVyMZoqfRHv7bfeL
lQ+zUMVcY8keCumrUqVcGcTOxAWzjS9I2p6nlNbopH3tmJIwEeTgJmi9vTamdPfOl6P1HVI4grT4
KVcrBefxY5s6lhePFjSQna1fuNOL3sWEAmJUCht9GhFlzZ5HWXRaZg0WNK94u+DscGWn4Nn/3R2Z
uXfReqrGuq6m1tHBpuTE3HKCsqePntckfNnVi2QOlOss5w/CVuRFWKBcsmltSBFjOT6axv2Mfkag
3ZVinWWHUi9NgOXTQOWYG2v+MX4nJ92Easo4WXH+/nGVQu9FAJPjpyQI4we9f4HDuve2AY24zQQK
awN7xmOYIyttgCc107uM3hI6ggob1sRLj7nAVYJEKEQHU0JcWamfo8jxu50qOfG3dexiOCMBpict
G5NBUeptijPlmDQwO/S+wE4YDrveoF1iOjQddh/TJ3mkhR/kQK/2cMBtBU/1m8TQ++uJiz+1nu7v
lJsTCFgfqsE2gI81Czn70U6VKHH6wtkKh5oyrpQXWzdpZEySy8EitZ33BZHNMeoI7+mjhZWVS5el
8/c5J2PqceMzT1KIX1frQc46fcbvS62pyvOegLv+a5lIBzUTEBO6j0/NgPg7aV+Sy0fxU8wkbuPv
J38Ws4NJSTLZP2aB8FiPsoyaFdGG5mHt0SCwxVxMQ5Q74Qsg89p9gpMT52b2WMH6yBDbJ/j164A1
61MDeFnri0l0OpwAc2uOy1A2Q3rh6QYD0s+gkZB89h0wi5L+Qbv5mV4BEThg/wrL/MckpKiBX+WF
AFOOEQCKHXsSOMpXU9U4/CmtpYjjHocBQZ0UxkBWLJRxj+pWwrdeD9oAkcAtgACjyMzaiHK+KYvz
uVcLc36oc+Ym9icTB4gRX/V71pFIxkO9YYkncak+NsdCuoJpk2yLCx/hsQd1yaLVAyHEgCpILOTS
y4rD/UNKWc9iGeEXIWy6PDytNJOqBhDBoi2ZKUKUlyaQsM9faeEzxbKONEmCJ14lGSM9u/IGsUQ5
Lf3pnp4HSLeG3nCyCnexOqAEc/UEtlOuwPuzLmqs0+cFI6mek9SEqGh6HrF7ixd9QHcUEj3P5LQ9
8STKUcf8OhtLu4dJ4BKyrShuMdyY+Bhzk7XC617fjzHKa22aj52tkfT7dYCWD6gfUER6RZql5ye8
9dzK2RXC3lSL1CWBRWl9Yba805me8J3gGREJyF+vTWbG2q9ratWIE85MGMI+YG7LSC7iRhYcPy9C
93I9dkf6FqOTyqxHhJlHXFRi8o96fw2jkixX2Ew8sMKIv3/zghKAC/D/ybbOgOW4KwheKyjMlsiv
V5YGzl5nb6kNqYD3wFVvmVjdFGSZIBrhTtLkNAF3PslUi5JdVQ4mGDwIpfTC+hj/29vGKAsM5pKd
ed5cJUJMY6BiMXaaDO0HIy/HGydesTJX6tf5hwqbs7avQCEccLtCdcHpX05muKPeDeLWxm2dAMZt
SWzfWF+97qBXbiNXcM9kYwITMGTJ14HEMwW1EXHAwIf1ccOZ/HoYbPE63f03rxiSbrDfX9jVVMaY
Oevaux0c6V+UHkAtUtuM34YK7/eFtcbWvj7356eEYDQSgntvz1THTH/J6FzOaUS+kgl7l06cvgvl
GLgayxtNUDSeJaySTi8FGN81uveclcuVKbSNns9XqDZUY+qEeC0L44r5XnWsoATj10WVlkjx16jB
XuKUgfH3CxeVniVkLRBhRYJ5AWc2zAAcEN3Z5nSFNR8t2DL3+q/gtOtTY6ZEVxJLgzaB7knTdAXr
PzTnw03SmeLUbFQhm9PJsmtnn0RnRSpOp7udNQz5bybrHpYnOgzlRZ2dhSnBnq2XK5BMiZpeGI+s
YSS6B2nCs1T0LsxknFJIqXnV9+5aGC9wi9ug1hC/B2W9Eg4+4C2e1wDwE6idRTwvYeRjZ2y0VR81
1a/H8KjAhzBOd9oB7vFBYDpDCQjEcsy/TG6oXBmi7xNWtj1Bn8SMLm7tgP7olL0vatUIC8uzXKkO
ZutnD0XwkSrS5UlnVRBdhFe3tCifg1oxnb1iJpsj/cHT4ZvaJ1LhWoA4QP/AP8g3gd5+cq3XAuNB
I/8OvwnaidAFH+SrlRj1GnJnqvTAvrr+SPlv/vr9YVt9c1B24DbW+63gprtUn935g77svDIG0zPB
MXTk4nmksywTMufParll5edP+9J+CX70pff7CWRA5h/iJLXYMa02upHO9ZQh2MgMKdub9yyEM+1+
nxjspksn7jS2UE13u/qAJC38h/XdLsXYRQqkOgudH0Jt1i3xtyqQIT+Ipi9eM/VQa7T0s8x924Lc
TFqIgOGbS0KNtfnJ6cK9tkJ6zsEGMC+kwYuOztcXuK4Eer/NXTbBFy64cM0soDMaXgHI5CRccjJC
bwlmV+ccY2hRybupKD4PRrnr3XvE5ALajK6k1z8yG4N/OJN21hhDIliVoghbV8+MIsuIB2c2LOgM
Y0r8UhX7W24GNMI3PGe+SUeoDQKxzc0DfvDHX5ErSgmBivON2q03EkU7UjNqLK52brKuukk6hAo9
gdp0mz6haeC07DsL19EAmh07Vl44G3aJ2Z7A8Uc+xJz8GEZ12jpznIatTK+oyLYCJ0fTpCotAxVX
6IWcNpSPGL8+Xa/lbqqEmLF3z/Hxsd1L4s2qLj3+hzR+qFf7+LCBzvjKnmV3WvAVLNKXP2mp9pd4
ws2Fykp2dGUjEoJej+WQHEaoeTYVSEIbwl0gtwknrIaJbSy1HJz7FoqppbQLEnR+i6wm87kpJ4Ox
5QBO3ini7uQYbRoGXSEikP2eMWd1fvIkM9PiiQqRqymwhjNttjbTGpxo0v9Z1lGJdHJIB7VZvs2J
0c+9ZlOxbR95ZU2EpgzYMSPNPgL/hLrF9Rtfb0/dq/FdYji+FA3F5OBexWnTAeDhdg/g5z8IgWxS
HQSylD4UepiXEdXuRMmUF1JCn+ifS6yJcowhBugBhXWvth6kNQn02n015OvNtGWZ+kJs6ZBHI8qn
3i98BQkk6ZI6CN/OnHEF9W0advxe/XAW7Q1klIbN8mkIFd8yH9uAILRcGwEzts2b5Y07f7BMPp1+
3bpIotaHSg+gmAkU9ff37aDFXwMjpQ29Tnd7dNfVjSpcXP+n2paOpucZmQlT5VIZ2hZHYOWtcKEx
dat7bHIBeyY86xEcZKq8HJYgHcIMGu9zsxelFrpYTohWBv0vabGg7kcv8J6LSc0WfBtOa/sUCQCG
mjaRnlMhVyNrnC2qKbHrNzH9KoL93gMFYrxw3Fm3SM3UihIZ5HRkoou1Gdy/l0dxfcFLjbbHFE/p
o5UZ1m7YTEpr/9KbTqXnJLpdE4KHVjPREMFvVUn+JILD1O9XebVmNkQnKInsVFOqRUeEQJOa3TVu
kh/66ee+5ldRFugA8bD6LEsCYFSaMKqC+r/gZYwwzdNNDsRNaSeQK6U6zkn1AAfKfnZbr5ZwfI2y
a+Di7t/2jnMD5WOcii7k9EfpmAOQZXcE0jUwpMznIly4DOFp9MqfZcDDJhlpK+msYRwK/paifu+2
1stjPZakiVWHjc8tjEaarvERmOsXrl181Y9NXEB0RBleRqH5UkQMzYRIF7k99H73esJaApwqWygT
6fVohml0gxKHIcq7+7/gB0h1IdaK3XxhbV0TcRj3p7eiMSsc1gSyqk+w3niMoMKBsA7dpf63fVse
vDQVtYmhsxmNclEDcl/RiXunaair96vIudsBv+9vEyuglMrmzJ7IuiTAG0d+DDG8ZywMPwvvv9la
JqDBSjrOGAH6EgqiEcOUfl1rAquq9jO7aPZcfNU1WC0E/zIhq8wacFluFNXps26U0Ud+LuBT2kzr
FJeAiuAbcJBcKpQkr4C6ZNbwqJqu/MWWAayQ5vSbCZeiBUKN8XN4AAJBgOFBqZ4Cldt6JJ0Ciomn
afymF5Pp7GQwcgDZw/MUtrEzTOIAZe0K+3w25nR/TfjxQqS4cK4QtxaNYbpm5q+ZBn83CyXbMqYC
xHjqX47bQ47PzVNCWzmrftWmN4zwGT/6EqYEO3vmQxqIacuZOgUAvIq8zHqrEUCYxygNmh8FKhF/
7kG8fvpmWYjbdtTIQYPtURMeZ+RVy1rJ9X+fpZHe8s7zJAwNxX9DuUCmPb23hM0Y29YZtbUA4Jmr
MWySOk1+uKiUx4IWwvg90M8CxdmkVgHLQLnb1KDv0WQFMgQZEQVOKpEmZ2Uk2R0mDQIdtWFrxqIN
zlkHgIzK8DfHfpJm8QHzDvy2fuCIlmz0wYbSFZopbS9jS1XEPKTyhTYYwu5uK8mrla9E+R55Q29B
dC9epWcBCb5ZGefwBZUu7AmZtVjm+Q7K0yo6ZogtYROiSBfSXuYgyqctO2mjmr4zDDiQEzpa8W3T
MD5q4y8BolrhKtHxBuh/MKxEi/PhU18Idxp5H4s5Yk9l7GC1bAwdE2JmFoVjerkmXHdgQGHmdHkp
KLSfZriv57RIdTZ4MTU6xRTSOTIx11Iz44dze9+wrnvE3/hspaGlGtQ8CO5wJjzE8O22bw8rkO8A
YP4bWyLEwPFRZAWogwVgiPRzDBOuhkqWDXVnFeScKu1pTavBkYDu5guQD1RDlVw6DH91+i+u2C2F
cNuFmSYLvssrfog8lPtjhLYNxcXrdPhvm4ZzU84U0JrIARR+coySRSQ0VsLLeJrDvQzK3PqaMss5
mIL1lUS/CusBlRQy86WDmBnlaaj41KyJK786DVWKyxCGvivuym95fp7grTSpd51SMAvdI1hrM2tP
NSc3EFv9d1SrHyCyrb9FhzN2C96TNiDUy88y4mwGSkf1R6KneZ3nbFgrV8Fdw8t94LgCQ4Ys6AwW
LUxVdlYyTdUtJ7qt1OHuVr/sfvl/6eVpgVTsjW0WjtBjh8FUYdrd8D5vm4dUWbrTuLSew0jKG86B
IuDF1vCkeNDsYq3KBz0c59Zm8vpKls7PPcv2pMrNa4NpsmTIo6GQvyxB9HtHuMs2iOPBYqxDUK7w
l+gpn2h3fAFP3hyAPqQ1m/FQw/RHkcLLZ1grWtYRro5i5v3i6rAn+JD7LMHURonEMjazUndJ0y14
CsbziHYkZhjsqZY2tvx29FqIIw5dThTcceD1j9gj9is45xqyIRk/9NYaSQklrOrfKDDakpFgw8ba
3h6Cgh/dYyxjRA0PjxGlAq3t6CimpuKwUrWQF0s+76+y8V5ax2D4EFOdbai3km0jksp0bHd6xh3t
QXqwpVEj9w30F6DacOhJtHy1XM/q+2M6WqepvXxc5IOpJTcSxhLvfouMxCSxNi8Ug+CNbiOoP6VQ
SPq6g/Fb7fzf2f1VqOieJkcxxnRXrL5ChiqgmCHeqmhZQ0HtUUvm4GtAliyCqFI3vHmKjccmACyv
ST3f45D/iFMY3QXd8wXzQrxVr+mG4BEzhaGKH1z6I5kFGk6Nj+39/Abd4SZ3MaNIWb/XIPjZ/+Ng
4CUpgelv9ir5YUeGOUQCDtXBsCvLqjg7vgB14CSbIEjqZdYxJfWGfccMnhXEPJXliXG1OIa/nfg9
meiWjs1UvykmbS0aTxEqm3lflNWTVbz88+2x4x8g3HkdhqNU419VeSBgF2MLHCPK4WUHZm/ExleJ
08KU32/f/ubEIjPyElMQ5kra9MIrblgXEJmQsKKnR9cBFqu1Mc3VDvr8upxSzM7gKlGENFO3UBWn
wYh8e8ZTpcB4AgMqO5odHQpzJsMQcFbplJQcKk+yqZrYwNzTjz1KvNQreS1AVk7bzwfob59TLl3v
Qt1nbw8Kxu5j3mbMZSV10UCcVy/R0ZAn3HksBOStU7L7M3C+KhF7W1YDGuRJvWen18nq3tyYaHso
ekf7eq69u1VERBG0QSNceZGoXaZfZf7MrB6KK4t+Hd14seyUgMuA+LRnGk626/+lhRsoItDllQa0
sD+VjtgHxPV+j04UBS07Kvi5BORkcHKfq083HHIUJq0C0p3vrXjq4/eCuZ9/DovhAdwdjpj2lWri
JGnE+gPWJdxaQzK3XG9v1ax2tXxRZ6tr5eUqdNODTjPcjrRjX42ghuKvBAEonlex2lz5HznH5LXx
F669Bz/nwShy4wkXBJPeB0A9Sk56ph70EHZ4b7WsznpsSX0XOrhOfWaALcmmgWVViDoHomdBRQ+x
nnFtNbFlRd64Bhmdcl5orbdQMkYjm/Unm1W60iEUJkErAhX16amQiTofQvTyEkir0InLM7rEU1r5
D5KVJedd5PoW1B1KP4BoEdbpCkIw6trgVCVuA0T0c2YP7IhZbsAPgxmRHVBqOgipCkydEdX6s5j2
kvJ/SCj7Gob/sr8smstptUBD428k9kLFM3mh9LiksULHpTCR9iLsoQYQZUr8nhJD+sC63xL8zeQI
9YfubfhhA8lf9XQIfVFJTv1B+8eCX47Gpu63WdqPtB0faRQHZCOUSeNUwXjGbq/vexVmstH0UkXD
BojJCz8a8YbxSpZwVuHbGKuUWUiHM16kqTcesRueqvBkBOOJDADzq2bxTkARDXt2xg3f2aCd+MYg
zpQLbdjEEdnW9kxz09sExVIWaEcxMs2QbIMkldZf0/LNxcBpO1MhxSkbNViDQ9SbhHgjgN+ExUFt
71ORWGwJrzTMcidQVmXq52sXvEVZuV8dgkhOB4T62M7svcBYtvPD0zuM4wrefqf0/IfHnyLCT75A
WA0vivz51XuUC5ycBVt7KrU84utgJhXOfMZJv/lDD5N35+e+P+Vbc9Icq7kbQt7IH9HaD4W1ydve
bOz8JMVZ1fgSHw0hcVjv9v1zdS6GW8ti4j/j78CP3jEGSb9o4nYfmjrUS7IXNq7pIS50Vh7U28rQ
veK/ciEoOiIxV+VruN3QAu2dkr1VAhHfX4m1ISgPh/Yfii39n+b46yx0tXSw7gIDItm3LpvuVn6b
6GDXwI+Qo8ey1U87X0h54AwYYOO6h0WrfDt2iIXmzRRTpWs+VGcXjupmgAY6GSB9865PuJ6s/33f
OEHuV0qN8WI7bBjvxrkpJUIbuUpbyI35jVBjE25X+SxGG1uI+A4V4V069OL8zPRsK5jXbHM7dO21
g2Rb1TKy/dI/v7rkNOCjaw+IQpbves57oxLMMtWkboPNILZ4gtpWjjCFNrqXS6vjQcYpzLJb3S1s
vZRH9Hw76ReL5NTvs/BWxxGZnaNsDZbzAGXpGKrx10cVDfnu9qk8epnpx9jssyMYJ1iiTQlAuAkZ
28M2ztJl/keDm5isVoFUlUOe69SZq1HIv98m9973XsJHcvRinsvth0go+LCRqguH4X/3npvhaSqO
5Qty5Q2Z3q7GVFgUP3PTD3Cu6Hp+94c/tqLns30FZgzhW3+C9qeM3p5+IHmOcsJrwRaZoqWRk0Jl
9uQ5hBiY5JPMEsXszfZuyRwQ2xDFmucXrUBaF9Ejf2yvxpJswsC5U4HM0ktb1baj2F3hknUijKIE
fsUwqS8j7Y2+zStu1/gRoEtD/CgePQJbhB1d8ADinsAdtCBmiUsPtE6WFOak51USxM/CzdWK2sbE
7rhiHrkfeoykqvx6zZChBBZp3sQ26xZgIahpqz/knSRVqO+J+/WWlWQNlVK/taNkYAIyinxjva6l
TmXsJ01jZ0DfqgNm47A2bAQz7ReUQ1/3yqblFli0QTDMYHnjvfxwp0HU7iaNfZcpy0VGjabv1ZhZ
X+WhoE8scF4ZAPvKADEP4iSC0u9clr8IUO8ovbBEPIl7iKz7HQS0vORasRshK4qi3rj+hI99QkPx
ohjTC6d2XD4qeETgbHCCTUslmeyQCy7XhusjJtep4zYR6JW0JJWXYtvbKnGj3jmzb8QBcwkVeBJ3
F1k4ejwKH1QZhWOkZmGGqa7oPkg4XzTifvfwAVvMRdX3/GfMvwdTUOICD3jwKEhGjrxPSWIgEjcM
a7pFX4Vn7V4XB2oj98yccYUrpzbjrUU/NT4mZHSoxQUsIMvOKwUyiFPL1vEV+AH3wxUr4tE+wDJV
I7jZXqZvEDrPTzTxGU7rAoNdv4YJd6kc/s3MyUkkR5oZmb6Bs6Olcj6SG+awuDbxsVBYAo1AKxkH
7bfm+P9WflB4S8K8r0mfK5SGUSLghVj+RkIrA/M/2EtD/CC9cd03oWfiuJtliHZG17NrFzUc8xND
u18aeAOIrRXDO1aKTvNdFbF28zFvLy/XHRPWBF3NqvPWjVaUHeylhB4cruaR/jT2k2inVfZMMocg
xNzaqbWCwafdNaieP9x0ODs0CDXbwGqpKHA6oEG31x8jkhMe/Xwf3ci0Z5qUuo18j80w59FbUuUx
chGwVmVm+SGFo6dd9ev4Sk+q5LfiN/yIkm/iOeWUdYFPD4Vb2C3TQ2ZM1NtBE4SKJIRwU4oLiI8m
7dagXD7phJF9ZlEftQgfhL3vIJ9MXIqeeoMjp0YKD3MOrJtXWyJp3gSx2Ke0lN/rLw0Xi3pFxzld
mYxGaIKhg5KNHqQ58kKzRNrpcp9k8Z71NAXZO9GOaQ/8uoAij5//RRDDqlr8i4HGwLz5MDS+4shG
HLsCFB7uYcGQT3EA91D3bKx+4sTHp2Uv3V/rRZT6rZ/6w4HXC9ROJYmfnSAE9o9MhTngiDPUlKTH
9jh9T7vGAuuxSWeVVsBJLgpu2Ra3D6jbUUGQcpOkIK+hCrNQs5tEoVjnFbptB4DMFi5+PZXjOgkj
GHM0Qz2G9w2SD96T+FtULkArFFQUDFxM2BHyP+rg2We7tcBd4keqFfE41Ziq/eedG3Vc65SmUEBB
5kHy3SBnh0ZEK6+sjK5X8185CAFJDektqhneL3rb8VOogclIOmJQEI0/2AMfdZX8seGMFjH92nAh
6a81FyuuBP7S6jla4kxYjlTD1snjS7fuLV4SpHvJlY+eBLe+hKfZs1abvYY9rt1kcgnSyDekaUg/
Xrsyz6SR5IeZNDCAJoVkLpiZDBNgQpW3OPG/D75CReFpxTtjqw/X6BHklPG5QwVf86YbgAsWKsSv
tZGodcK75+Zc+NZiX2jcPsHKXvHfFZfCoPdLlWp8v8aeW134LtcLP8WmitnSz/iQxSPbruUnjQyb
os2XUo3gkTry5PYk1y94X1YBJ+M90Nd7Cs86iNUUu/ESL7TDIppxb6VbqTh5LNErK5ixqp+wXWAU
rSkDdI+Tr766X1RQ+TvcEKa1l1P/M2AAm8T3FYDMlBh3586hvlQ9H50uW2CMU5voB5AyjOJZs/7N
fAEM9yuWdzKH2ZehVECpGLfVQYXnV0YtoobjiHfcVmoxys4+XnC4+Pq6kyJbfxAAI/39pKrNNMsc
frOLZ8r+lkJ8XNH8ADNQlB54vEsBICaP1YuukJ5/G5FCj6dVC2mFT7GvJ+t60WAaoq6zxQNx2H7o
Pjk62NxRWjQzamCsV4EELy3KplndoJ/Xahu5qHXYvkc4HzhHFjv7gcphNoay8l5ExvqEVKKF9JlF
7jg4F6FLCfY64FJS62xYaYp7Wkcj9Gw79nmDmwPvOYT6u/NP34rZqBkeFwjyL9qY0SZpShNHI3EB
0Hjhaae2LI39bsO9ut6Vq6ur3MBM26dvP8nHChpd3+XlvLGC4N1AE7YSo1r+penUhZEaxxut9vji
pcHoD7ZeTCi3FteNFPEa23XegHQIMQKdaJhkFmuHHXfAHPjToVgdZkjiOPJHfm57xbGxUc8VU4+U
lJazmldA4ZYryx4+0//xfwj5OX4Nm/u3FSu8y0T0ulttPIPIvadVSTDDf49lqMavjgwT7vXwLHCl
BxzE4Fl5Bpu+Y7DxyB4qvaIQtqL3iBGtDqp+seTg1oyGk3QSgEj1j0PXUJtaX+22/pp5POs2daPF
wxiHgN3PlJpx1p8CNaNSGAre6IKOMrb4/bjCIqisfCCXhumsEkwHxnVj6eBG4ipOk30DSJfHWGts
hL6WxJkl1EF0iA3H0s11oE64CFzDIkIeyrzEn6mcxd3aEEEk4Pz3as3snjrVnIC5vQ8ZzSKnr9Ec
9ta6Jy+JeWh9O0HFfDVdQ9mbYC3nUfic4C+tcPaEEpUf3Xxeg//VnEVaxgyG9+DRlO8Q8kFzJPgz
ltU65CrCVqnGGZ5gMETYm3kWw9CTEctvAXkytIn0viBn3M7t0im4wsb4eKQMSfZ61SsV+4y9j5Eg
hagM8NfRSCB9g5lu+Gq8AjVevtuQcyRvH2xLQLpUOJaIwr6tsx6JdS77J8I2eZoX3LZ6NNKMZWgE
TYBds9dSKeJmpyGgt69H5uO7fRVJtkWM71VLeKWKaDJpuNwlzKVSpy1/qa3i5stRioBkxkIy/tsx
ctwqIe8i45aJbdiOjGgBdITJOUqKEg2XyXYpdgCIwnMS727fgtLRYMLH3eIYrbvEQBMCJFi+OwYP
l26haHpwJWX4uEXbKLv5uaEsrVhbTr8ZDSUw0U3oAnJMHU3TbcED+vneefkRuA6I7sQKkx5QI1Wo
BfsPzldLKMNPmnA5euoSwzxGOgQSmQ5x5fK0yN5eYTcRtVx8RYAJUwLfDWSxxy+ZMOzbzH+SoVIq
zhx0D3C/eyuo6KoH8xmxyUCCXTYTIZ6Vu7F9DPB1xdO8oksxkdms1cJ4O0egwSZxtG7uZmL6QYQN
J8OLxHQ/Aw65lHSztcQ9dv0FiR4diPw2FoX+POrCSE3UCoOiyLGbuNK30rIz1ih4BBUgSpAOd/Wt
02FSsRdpg8pT7P17z+BA/SqUXuBHhYCsHuDQbZzzxz7PzRmGCoHSJOv28jPA+9o7r8G54Uf5ul8h
5fhEk+RyOj3aiglvoxH9WpT7CDV6yAK6FxH1O68mSBaARNJIbVsYuql8ndsjer+SN7PSKfY7CxE3
wvfLnBfp9fSwj4GLm1CfWxV+FRBT/MfHjLDVLBUSEqgavY9APQcS45xBOAgaQRKktfRfVAbB/lJj
/MMQvcJhryffR44OT/b/f42oTKoAbdyPpBRBXVDz7AsN31HQq3ldEBabRBX3ib6fcIwIGgZRn3JI
KXsolnjvGkLVZAvm7OkS8axWsYMsgE+GTRk67yFCqCj6xhsAcinlzJEJqv3b+zATzpHlFv+/CPQE
ulnwZPFsZvO9Am57mta+L915/5Tf1WsaGdXW41X9+gVGlCccr+l6zvLazqkpIxleca5y13Cdi00B
O1ZDac1pTkrj3g1yP+kM48bhHQr09TYoebM7F8B/3MDC0Dcn1biYnrc4p/RUN/EfbQqxHDyj4Uun
VbdLnVugdHAqDXtSuFp5wiLQd+BPW9+4eIhzBrI+lLf8rc0hiJJWjqe//loldNs0G61k3rrl1rcK
WbxcD7vsVXQYpLJkvKBqda8mTq79W+J0YwRKh1CBFkRGgvTjYozThhxSiApnzUBvOSqBItd4wv7a
u98tP4lAMqWoByjjdSZp7OPT7v0Wb7n1a+ThhwxoCHaCScpeZSqxNU4w0j3JqOIU0j1j0emHNI+3
759cPf9CmpMAjwB9jV+t4eMIECSsi0JP8LsIikFZHzRyr+deySUQoMs7FJmeSyej7e8YVvLn6pUl
C+Hs8Ag1Z7cPn2ZqV22RP9eeYPiA/ilkRv3+gtFfLtKsDObb7tO0q2NPnCZxRLk0vjRbyWWOGUWm
GJNsQpYalxyH3kI9Sz0ySIAkwN0NUj6kGuC76/gJ2Aya3d46tuzsLaVdzi3QUY116eDBUWsYmmjp
04AOtkTf8nmh0LwO2qoBqX2iodA05bugTCzbYbRL/kSaQmAtbnvNmHAiE6fNscyflu6ecDrqoq57
5ALUBDYBEpY6gpmcqFnLbpGySL555un6wUa2euJRodC1hCpQAeDR/vTl/1PbcA7FLeQ9c3izGIMC
ZZWmVKHDRVmzObcQzDUo1vHJCq9/Fp8soPFlgGgKRxkVUL5g6HomH1pr3kagUkaCECWqeyhIorpm
960DhliJzQEck9IDkz5g1+uhlIC47H6Y7ep7He67SiGIEd5z9JNhG53k01c9g4Dc7+CHM8kSAa/I
9tyIjavf44M8pwVJVihfa5yq4XezPKdlqE4STgHuF0vM/mWVcPvVarkoyyL0vciI0vkiwaNwwnjI
a4akEVbPPSc+rLrhX3FhiiFYaJE3gDRnDuMIMawAkwlezLxFKRCgbflR9f7mF+h2DLEOOEuoYHcu
sn8c/x6dy8XNqnhcRsmotFgIZ3thVaKUaphBHO+iffPSsRMhgUyG3C9yPXbHnM8WCR3HYar4UuWX
kJNndDRfOWsI2gGSIyEPj6OHLchZtAWiotA49btu3qnTUuqjv8XY0SgeDJI4UCzWZug3m9lX0qBz
ezDHfIsgCj72yl6OeTIEhl1cknf1ey8QfLDF9F2DnJDqYh9GYs92Y/Qnf4Sei/q86iJPUPEgYINw
00gRpXPOK3VHmJJZU32ydvX+wQkXEbBE544r8sKSzhY5Up3IpHtf4aTU7HhoC23+zUyoWHIfoTCM
2vuqy0AObyY663VxDpKas6jYGxAtadartZkmG4A/BxXI7hf5+EkLZ+ratiH6tBDb+RjX6QUZRlNr
qELYdYRfCG603DpD9o9mhuUM38xqPqOGyuRAUdtGjyhqCm6XjsDTLkwyH3gSXL92+MEXI9i6PmL9
H8jLiPE9vJmfJNXcpbVLyLLRqBT1813JMUerFZC2Ab51WgxBsiHaUTEEL3vkKXM569ZUz/g0OdT6
XaWkuh/lRcCMkfAfb6S9oLjFSFAyJ0+zd3EsVNN31DsF0EuSq5iM+W5k25IaOzfP+Zih2Tv9e6na
TPimtY2BtJw9lX0RRLC4501r1AtosrNFU0DoQR1t3vn/OU3U3904ppfeR/w2+UVVuXXiXJ5gxNS/
uo5kiqgii7Mq8nyC7n8FGqSgVBmTVtIJaxjWkVdHQmQY02uLuTakcwc/TPAn5PNfCANycIqECuQY
8WPj3CAr0wfpQ7LEJl+GdfvXYI+W24Y1kt8IiIe8hsfVr1dDH7JGm41RbZAaoj14safTBCFjXI5T
7oO3xV0VCBN4JyUlHNwKZdPXnH8NUrEoceXC51SNpv+MacR4PIw4CLtl1LCgVeJUwwVhWPXbC6rJ
p0kd0iPK4l7CUtrEi03i7GDV0sGL1M8MUskbUwh0KjBRX23ifg/D5qxiTDpGVhtqUIg78A8LDCTs
ixpHreDaXVD8RLbCc47voDHtnuCSb/WyPjdj+Fl7hN5AI3DmYzUhbZp9ZXYeqPL+/Gb1OCSKE1Jf
6Nz+YOF3OSjLJvEnehPVUQfM7Yn6/cZKu1kt6rKSFxUPjqPiEyMJMvvhrMpGAiD42iy3eNg/TVRA
/1k5j/vLfa85MOzopHcEQULeB+mZZyx8LNFuTqSs0GOy9yMGFX6O2XKO0/BTqy4GqWUMBbMiGA0j
l1eJXvsUg3X/iYviz/At+tAWYNB0241KrxBeP1Q9DvS4O/McUByMk3CQRUBwGu+E0Ssc6k5q/ZMh
2ZiB8dyWwOgaZj3K0I8S8PrBTge7ZfzNR30/dMPQNor0emn/WIZ4LsKSgVyKtTDPZv7sYemCjvwI
Hfj6sqX9OpBoq5+lzMjb5sZup3KdLVYU1DannBWMUNUnS4AzdcyNrh3CprCf/jBuo8mTxadlqsP0
jg6wpjDbvQd0LRlqYnRfXcBc+WSZ64+dHU6oTxiZD8b1tUBgo/z60wOYeZTjbwKXFQPg4lwVFZEP
otx6fw6jSVSICEaf068BoV8tOegDPcSeuyGzd33el2JGNT33986pqnFyxfXhLhonxvP4HOZjSDGy
LVB8rL/jl9YW4VksQ1NhI6KJ1v4WZecmAFi9NFOl/T55L/g3+CUFMHY1oJClzeBiY8xF1JFiRHjH
C5oOezGad09vm3HKmZ3wAQZF2r41PbjTVXBIjBhiBLGgQ/LEILp42mGavhJ+eplYiSiKaAzFU8VY
uy65KYCFtI/ZcJCQMFC9NYsVVG1YrzU4tTqQ6oJ+HGcKXuDQrTkjYQ2PwIZpzSFXbqdwMdRtfMra
6w91ZgglW7S4l42ghvRRGBz4DyFgdtxZSQmrpWhx2q6IdYSNFeJWan3EhOLCN00tsmaXA6bEF0ha
7s5agkQxM7PNbWfxQazuZ4SfpRXpfmNkNSlO1FH5y9UNlWH1VAmgiJljJlDok66yDL8A8QjXj0FD
+05J5egBL4mOhVkXwLfkr9/I1x2NmHjBtW20HnRAbXQSSYxS6BzNq0sWnZ7ETylYVSztfr9wzmN2
/vbW6PRjeCgen5A1HtDaobXRhU6Wz7+50DQF6hCPwoz+kIasc2jBYmQK2NPt7Y0Lfk5ATEJmmodT
s1SSoxdRQ0CtBbdItjSFaA57lJiTyEDd9Jt7bcPGZ5nZhFrKOfsZ8G/bscrLtRxu5+wT7zqqvbMV
exUo7GEEMtdEvt7HtlqijCHQB4aG7cgoKFjEt60pNMeW4ecmOrTYLJQOkgxKB4yukd9hF5WeEG4e
HJ3Mw4Fd36PC2wTYDpoHI0o1pr1WlWbBLJaTYSgoSm766XHJ4JQejctqwQXv8Y/+kAuKe/9iOGDj
iigqLHtoNgsnjgavTFYW0IA+RGIgIop2fGg4C1cUNFzxIugrRK3AQB1EO3kJgHfAg2g70ZRh52XK
3AKRxoXmF/PTA2uXObjTWGfJPC+5+B1QVseY7oEizqQxbQVy6aecn4b6NZ9WZjuR8TzjcjfpR1pD
9rW3SeO+rxC0ZR3pQeVCt99B79SDGh+tNFg6Hd+uGu6PG1y/0iPN2C39qvkWjBukDHz7Zhrjlp90
xlptittO95fty3Uby8gTdJBL2tmMZiROWNXhlmgX1j7EjCv/lxnIx/xiA0sLz7Gt125Q8sNcbd+v
4M0lB4Dbyyjet0A5w0WA8nAAcYiSp+nXAXzu6knpSK6bS6Z1cnTHYPTxmjaPKiTKCnoh8bMKosXs
8xWFWXWutLJuR7j1PoydVhnmESMVusOtvoytWijIkfX8QS1c9kijBtFjaDXUAxywju6c124QAgpy
nWOA9nbn9vleFz/3mjwGJmiNHGijpJ5P5BTkjLUwf9eMcBZ2v0Mgmi5OPAWYVLVumwriam/h1PWH
MdCS70ZGTKfgGwBVzML7wczRv4Pbz4q9vLHGGJZRPhe5PdaKBWMgp3Gr89qSaftJ9/6oAMHv4f+y
n1MNszx2790dT0EuqMMICY9p5bABzX3hunOK30nOsyo2zxiwOk1Me3rzxj1tzfPye+vMNHheaYDP
M86J2u8oZqZvs9joWtmtqvcRaeIM30yDyGYg2Y28bROFssVmI26rn8mhULg9kT0qhxFSnnzU/crr
xoTSj4l9wns59W6rAEuCxZ1UU1X2WO12mr8XczqZcqW4JNd14KrZ2FfQ97L18JpW0pwQ6U13cOC4
5jlfBPnR3dtJguM0T8iS7x7eKoe291sPi7couml9ir4Lnu8sQj6hYnb6aVx6lut/x/BfYIgcsNCA
Ou+jyOYAIZ7qvv3ur4Eg8Cgv6BcI47aoeTLfk8Cx98/2eBG3jDG9WOCCTxQ6iuCaU7ertDL0XF2g
8K6I4fFjUHPltxXX8MG1GRgmQbmoj0fWzLruxuRW6G7RG0WJ5XQ8N/mD0/tclbCdJxCs6uXSIE0u
E9nVyPKdTaSADlhnYu/hycC5emDFBinkzZJJjeWckJPzyQ5o02DmIqWmVKnjJ1A1tdyy9inWPKgU
lmjiN3oHCDVEpW+XgKtyE4TcmZMFwGcreyCPQrMMwh1Oby4PUtY9MIfl8lhMYngHe1mdoeNtun/a
m0zxENsgnGqh7/cRtr8bzzYO+s6s1mqJXM5nOGcE3IuAszkdIBUzI4weYHOlLz1tE5JDkkdJdSd2
lNuZCO1b5evkjsk78wuEpqBJGNInSoHvjT+Dddv5PzLPAjSUy9RBw4MylTycobxAV5HqHNAKq4GZ
YNse0EYq99XSp90YbNp11xWZTYTuqGr/3CtAg7pRbXG3JIErPU4GSyJga8Utq2s2/v2x6eE3Plt7
XYKl9dPcKS5T+pv5u+7Dq/VIFoU95fEqFzofriyCQyWWlY8P29rFBuGq6kNAOGJvLiNerylVPXRU
0S3FbRW2nGuKpGmj+klWGQ/LOPUxIuRR2Q0aOA7P0c4ChgOXOyL01/6JteyMgH7utbKazp4Wv1HO
5LF1lAh2A+QdUNYWUG7/ONCtYxkH83ep9s8TkEhJD30CtqioTtj7sGketau+Vnf0zMTMKSLNzaeb
720Hhtd3Z8Tgn5Oqh2jHGBMnBdiGZ9M0zrTkJJbMuTixeYEA2RQC0LcfpXOxHOvxHO1oDCGfvx2Z
0/z03me5DBji23mbLOGBv2+fPXmtTWKIla/yknULAjSYhmbNqtRQcfLlhwBW7ArCIvjyoVpjzQW6
wGXDEpVXaZ1VRAvDWuzR72ouduec3KHLfStJIqEyE1r2bhkL89QsNe8iWEz+FnFAcxDVv2qHOy0O
81OjZbGmTsuQ8aIJE/npUSoOmCsdags1U67OlNy0uEMapxoOBnsA6JFLYaV4TOYJI5KIA3jufdOj
xQgBovOz9j7oOomwD1x8AKYIUlGehu0V07LUO43e5GMvPeWaNna5ovefnoREUmD7oDblUX1f5iHj
lve1XCZeeXcf4NqnXsLEBLMP4u3lhVn8a0RJ+vSyMD5WNN9nQkqPplnndU1bG49Lyww8ZpOYlVRF
Pj0+WuuTJY5/hvsV26qScPkPNjazfhSGdiapgvIIOlVzdbSg7Mqfcw+5Na0RPrES38/PBrUs1DTW
w7rBgOP2+SrtHrZdEaeMt0hhtWD+6AzxsozgpWXwzMKPw3rfsqWl4weFQsNGUrgIVfTGfcbBdiF4
5ssZpYswQwiLQxPCWK2iqxj1f6TjDVmL7JROxjpFQSWpzyUCcv1T8NSKsufpnbC1tk1dvoELgPoO
/0kIFYLBTz2Ui7JV9NmvRxtRB2nDEOLrr0nxznW5nnrkLOeCWDZnv773Pk8JczWHwLPQYv1031sZ
DZeY/dLqn25fPnUSvBMYnhP3mpw/e33X3Er2Xv2DpdxO90yzDspc2ZAh8noEcoLU+Dt11HOxBgHd
tFJY9OS83WiPlmuOERGwJknC7H2xzGD7ulKZdj5Zg/90rl3xa4YEdWpy/CucGuNM4xvxWLYdaxo8
2L5tmwBHHpar3FYGH7NqJj16KpsCdQ8Rvk8PpthdBgFsZgo2k7Td5p4eh7QyStu9brWfmhzE7dzH
3/V3y17Q4VpnTpkeOCFJI42LsWJ/s62H6w9P12wJXCms+HT0HgIY27kEN168pDpjwF+zlHX/+RoZ
69h8j0nP8F3SsSYuMmhwsQfEJnuBs7UIbbdJdwlitTb1/XG4B2BtvkWPAF9cEvDyn9Jy9U/BWxjA
I8/zSBWGT4bDjOW7pC6PFJYZLfqtK+v20ffflwL2TD6tzP3Klxa25NqUhnnOeqdHSTUPsI/5JKO0
kz6NpUNfR8ILrXn1ZF/oMb06JAQiY2rrmb60fRngmfieQJogE/ylkz7R/YdYnDmTgydbznHIJ/zA
UXj+10KkwvexNNXf5AC5WQNHd5gEi0T2eq7Xs9BMuGNkJ62pwyDTNo1Ra+kYctevcctP9cR1Rl7d
QnXqii6btKhjIFl3ZLwZFYCbDqyBbgp3b0pbrEslcWTeUR+3w3dqA3rYBJ+hw+uyyG7OePMIeTvf
XaX+NtTX4CHOFc5wTfJTQcxW0FOuSQLBaSXD6dwgVhQOrALKDMe9WydEdomDOshVN40Go27U3/QD
vYvhaLFVOaEBCs3ly700MzZxZ+6J9kFS4G7s0TI8gQ61SEsn8k9OL8Bgn9dQAmm/q8QLcZhRZ/iN
VU20HEOwiLdNDHAyAx9kiwRmq0tmuEfHikf4Hz/13FKUJcXgsZGUf9lYkLYDKYPCA8ZLbuOrrRyJ
RHD3oMVa9/ncAeRhTRtVKEMLFQ5W10K/w0ViWtPK9qHkcxndtklUoyBczzE/4p2k9j8YJgMyAjuI
L/YSkXg+Aa0P4fEc1LKdBELnIHtk3o+wEONFqpfRnMNIJucZo1rWOlgxY/RiJWy0wWL1CZWET9t6
Ayfbein5Dpbj84JqJf9VH3fAs/SKPtEoeZwgkc2+QBLCxbt9t7u2hMaNZThfkz50FJn5uuZCejAw
6k64N5fmmQ4WQTUKYKin2htcSvjtQkeKudajYtZF+7c07WWh8LZ0GBaHQ8T9XT+OP4eMI3smDmXD
aTrrtsmeA8etC8nWlZGe19ptd+A21ZCBd7zYByeYsga39I9erIyxtVfCdkl0bxKjBtXSIQgJo/6r
2+jDiTe6D1RXl0xf3LDasx673zZnUo18MY+ZJn5tKUFWPtD4UGSsZ03nwKwEIhZbzbgNzQgqbdXd
oIbDvBrG6VtSYHOtelvZlJCZiPxRlaNfsMGaSUVkJi7kwAJsyLK3AXBH76lzXAqMKC0vfov33aci
QDFwXtLfTLVvwkoJsLX6kqrEF2MJUUpUtE84APuUqgtT+jdEFWWouce8TC3WNijQpdWNfKZuE5rO
FfdbFGapGZSiOVnmS8DmVDZ34tiTAipztfT03F51xF63eIWii0Xl6Em7AFNue9DbNKpVvpfY+ez6
nMK2a9MkcVAh/VpKq/Si6hmoajaZEwAMJJBETaZ+FFjyEaQk71LnA5DOZj0rJSBjHsufaOS+amMF
KhbDIerJ5lI1b9y5m9ycjkdzh+6iNiizADXZ3TBwBd5etrc2PRT3Oa9gBAdJueiRlOKnewe0CGto
zkW8QmW8r++HC5cft0Ydbj1i1564reVnvJj7sK+h/excej/wfxYTOn/++PZ3wayopjHluw6ix7hR
WpN3sMBTuSNvPMovNXpxa7SrTfe3BXl3gRFAPfN1SNJbhJuIzGlrzJTgi/12qqQQjf6dHOSuealC
C8CgHKbn7Mypv+auduYJ69BnQ7JS6zCT9BzUDZGB3AYd05pegXQxz1EBhzRCYWcfDgBqtAUEo1S5
rqDzxNcEZZ11GatZHq+zmxpWDCr9tr3ii7+CfjfEPLJh4hDqROfCnIdrO3HYeH4sE2jONddignML
O5sTiidvkbZ/S85dLoc5DxcMWo5wLH6PMu70YRMiSZzIVvlrAjJTFW8FwVY7I7uvWRcicbfSA5BE
a1OIbzLxwXGBkaxLiJXRAz8ECvcTIbK71YrIjvCnnUkafY5YMm4+kIwbT/P4mvjK8dN/oeeEAzar
CZSJHAip/24G4wHhEkuCZisuzKV1yNrd7NT8eXD9IgwA1XAblZCYOLDg8j2PgV0X2Q+uLW75qbZb
cuM+N2iDMAT+95FG8zIKye2rh3qVrBQT1MGk9XjBOpIVNcaUzZ59ciWpN528wvEOoZ6o+oNlnqVx
+71Hbwr0Yo/Tg3+VkHswyfFXwHtVrEjDzenLqL4i6238aYAyCY7/KCM9nK2qBC16lflY7OywZMkC
zorrfUyz5j+vNp9tPjIvzec7OQEipHFwPE1ViSvuuNJvOusBQ7qfiDHHL/BYi20v1lq7Pfs3HQNU
tRGYz5wiquautTK/FrpbN96p4BxtTVQ0X6NYe9BdmmXVfRjz3XoZdqFPlSfU93x6kqoGlCSDtEnv
EtUHiualOI+LLOB8i/X1t65VR/ti6sZkDxXtY3GZR32fP7RY3oi08xrhR0zN88mYdwc/i6a30lmh
+s4VosEc99C73D9DYuBgzzAkKuSG+qqNuhCc/QOv0XYV+YT/nfe3FWVl58E/2SSOPSZ8q1xvfjlR
BfGr+Y+G98USAiTrvOd2kn5UenReV3SAhlChxS/RLeH462WhnuhVp5yTGpSGQVWEIkKUphnSmslG
fOqK7sakslcSzlxCxwULwftgXmTCbldMMsGrF1FfGJxF5wnmkRbcVpFzlTkpUouRXnwPZbD2K+5e
Y9+six6UWbeJIMNj2W4urxkPhySELQWnnhtWT45S8wpkqcIX4xCzMRv6wGIasTnagI3VI/7BKlO2
aRVWdWX0sgxzKVrtSZ5uUw8JFqUVCgKQdD5pqFAtkbWRu0DANbefAw1Fo7VrYeMEKvlhmu6CwNdt
74f1VgtXvEYJeGCf5mbIApXKet4QrpbI1AXoeDirxjDkiNrnszOxH8hCgCG/IxqB0z2XtFD2XjVz
YtR//bsRmzTVsag907PSvh8ecdeSs+vYs3GTglk7TBavSEEJPLBsc1esFVeNdPkRmXo+NauvUzbO
8qrlj8qxOyx+8ZGt0+qG2nt/cu82ssLYRbDSPNmMTx6BhRWh/PLwpvBFmDk29DLj0DqWKP1/GDdl
94yWBehnBGpPx0ET0NeEbLWR1d6jwGiIQ5I5j2MuyPALoY3M16DqOdH+WI41RdFhUvAELbhcPNJL
FAsOV+KH8gDE6hlXchhZ7MVztJbgprrXVYEZLSkYGq9RQ1fMYSGPSXEh5m2oudwXTFqhwakFbEPx
gC6vvKTU23oktREB0LVIfPWcgF4DWYumsikgdKGha/5znnY9YOU83eMMj4R5e8gd3g+6m7YAC2sl
ejE17oxbJExwr41Xunx0C+m8TcFycAgu3xdHoINeuL9HMhIQMIYtKiGA9a4b09nOQ7o/7f2/EC3/
NyMcDJxpDRqW0W3j/HuaUPJawYQ+O1hIssjrdgl/g+zFkIk2lv8+OOe/Cdwq3ikEO818Gp6yY8Je
LhR3Vcb8Fli7cO7dsHou5QkvYyKnFQjCFUSddZ8gXV8QuP9MEMlj3d72dFDkvbfvODbqtzX0A8NH
a3cGTv5s6HbFZaU01lSwynZYnq34z1CG9gcY4GQo1fPKCAZzNHOnfH1nptxnEnQXksbrMcvjnujU
gfKHx//Cvv/RCs0X0fYakmIbZjAdS/fbEaQaB7IC91+sJ5FW405GTZbOXFUHF22VC0U6qWNWd8I9
SyQr0YpJH+pv24tl2VzF7pyHQqeola3xpXvvwMdtreAw8AKVROCC0VQQlUIOjJTIiMzbSakIFyck
Kg1DOh3fGFc23ti33/gZZ2aDQMltw0m4gFBEcPZ7KDcFqQUKtUdyy6tnIqohFwQMllp4cHit/OQe
uVu/6k65bthIr1nFa1OwXchmGjvKeN/EJWoK/t9J0XChCvcJ2g48r8wB/D/WB2qOPxRdGeg2GEdm
EolcxqYp0lwAtYJDblIlkPpHbr1hDItVoC9E8SMNscl6fYWzU/36WkZxtO+b2uZHRQZ/8vkLLaDr
kvMgej6tXIzoJcaKbr4dHAfSH7EnzUBb9o6zjZ0GYM9tsztyeucv7TPT3urG6YIq6n6FL/2nisub
z2nEK4lRl/bd3kL4++POHss9ifjBEZIx8I4YagwLBZIonRD8bQOwOXRnyPN79gmgJi+tA+gvWkMl
X9ClhHc04xd9cyoPS88cbSQjiQ1WLfWxgUzlA2EGHWjTxMdWiVRZmQNGNyDu2VR+cBrNEKzEejHf
CPZYHLkmvNrwnCdmMkQlR3i9gOAMXeGrcvnN6mkAdTW4xN39/A11ZgLwXw/FEO9uZVyi190g36gg
ctY1phgDoQh4zHNDhFOz5TW13yP5QWkRy/5hgij9sh35NRLHgJimgZ5HkNy0pkX1DjDaY8Esh2gN
1aXWynhg4LOgpkMIxc+Q7trgpIepCerv61MzdLYr0wEkEKoQU1OaSFCQhQkxDX8j85xDQdyqOHz+
eDSJgaNQuh7DiMvb4OFFZOqC9ckMTZactFn89qCTgHcvC0n644FDJR+5GtOYQlBjcqOG7dh7fhQe
rZv5fu/Pyjhtk9QvTUSZeBddaK7/UzPTqaGnBQaqX9GfFMLMqJ6g6CT/tjl+XoOYbiY6VbbUUIWD
1SGOcKBHiRe4aP1VtjIqLD4CbLbsS3PicjpuCdWq+aurJNKPy1Pa2ZOYhDh3C0pb1Xr7uMlk1gb2
wo0C1+pKHobHkXycx3aZxnkLSP2rfNaaHVHlzube0ah1WwMdMuYTAI4K/ER4fa2EtOI1d705PwnX
6VS0l8G1HKr+IAA7lxwGdLwMVpMixXQR2cet+ku8BnPlOWbwTgl8WJNpu/hxujR2TksvbgfLbqHk
fIp4iZNtljVfSLKSn7b9EKpPNv6jExjPCexsG9m/xrBjmVqL9FHc/9UX3lVRQfXG943pjGJ0Pdl+
vJmcm03ejoO6tGwpQCGYOY7vPVBXJ298Joh8CPJEhEobPgJQSV/pzZ734GKrGz2cAbtfosYJMqpK
b53uoPKhu0rabXTrISnhaWHfbyvHsFWZxiTpa13NOpB6ZzZd6TGSLuPacu1B95PiCAVw37jP2otO
vHmPPNsnG/aJ23szw8WBQvTvA5c3dQms2CWjU5mriQXeWulmrRTga/DoS0q1MlgIudCRkOFi6uJC
SHi6pMV/WG5fuzCh4QFy9qagy1oGIcgX/RVPINeNGIVDL+IQo1ZRqqUKODEfjBChGxl9Q5o80nXW
405ermpIOg+LupSIFJKLEiuG4q84i3iACi4u4dglF2JAIlu2yYtHsMwg/cV0yousUcFKPk6wpAh2
edRhQ9cYWKI/xh/Te4E5oU6qhoJjHpuVAvnJKCWx1sFwwolHmwajsff2pF1c9t38Cb+alrUloAOy
+lnK2wicyQOCRo1NBQKNA0cJ9QtMo9v4Btd3G/tFzZ6o+FFbM+nWlO0h06kEVpjZJsYXYveEVHW/
P3xtUh2scF+7bVpaZcdWGSwadr9vMkYqlrzjqj1Bv+2LWHQP/fiMEoZUiCUy7mNBUNSE2FEUGvM6
Jw1jsBKN0r/0fGxIwvgzlini70HjfBnOepZovfEayq51Esqcp49cPlimwGLUrMO7WD9tecrgWlBf
x1sficvw/bxS+2O2pEBJYP0yqWyWFbeSnd/VPmvep0DVVswllZrDX9xjpF9VhhGX2x/EFEivqdwA
r2RkSqtmcPSRiAGlzDacl195SPvUrVnmlMTdDRJSIX7FMIQUOvILXVZvoGOYRiWBBFyGVd7YN8/0
uX/s3D9jlVrkpjt3G4PXCF+hO3YxhnDYwwsIY9wvqdYeCkWYjIVfV/Tspi5oHtGLb2GIlALgdP4b
Cx8LJZW330ulol84nhsyjApq53BPJG/iLS1nfjq7/uQo3FeyVGfpCKYH/u/S2KbxEeMuF0e4Jkyo
pQ99qgFqJq80ft3OAZyVB8mTfzTLCgRolb4EBcNa1noVZr3Gm5RyeWrnJwirxa2NO5JJLWFt3Afd
q1IMexrer4jquFpWAh3p3KoDy6ZCeZfo1dB3KWMr+U9b1OyDASZ1BqFfztWlZRZAMHfusltipGeb
StLKUWC/Ij3YurevBuaPVnE3PGaUEcfXdOcW5vuJr8MBRUnYqhuWPa3veViK4t41eEFaHBpgagfx
R0laL+MvbI2bSs5b0xCSn5K0jKXFa8NkS9EEQLNBWCj1t8Xoy7QCXJIiRTUqIwS3Z+iUHIWuU32S
AYzDDln3pokSpoqvi7wM21OU+kin2yvvFMnnkyIFTITaeuMlW+RwV1hgQJJbmicq72g/H0q7HAaW
wJRHym9gvaedqpWrQ4B1RWspLck6gA2g/C0uif4oLXudCuif4+jSaUC/3jTEkmxb3WIHl8Nirazq
px3NoDbu2VMwOzuj708SF7wDT7HxvXsnYaUdVwS/nE1/JVpgBiyD1inIIsfeV0W9d2J4X4cT1JpE
uZyR+4MNnrpRUFURRYyCOaad0y0oBpgeE3HmEu5sMy3uQkUp2hLK3+ZkKHqtVrj7IUDaPCRhgNvb
OxL9klE5/PS6cftCNfexvjWV3fUsUA7U7HuUv9z7xTYSnEtD6P49FicQBQqhBM+VBc1BGzQKHap/
XGLRDWlhqDZjNgEghrzekEGtoMFSGMgAMzn24+urh82dvaSYT9Hl0ga6OJpOo1rnh5LqoTcylOOq
ppuRKhRmGMr/bKno4kIBTK03/KitlKEZ5wqf35fxCOWfR3qbEtPI9UvJNAurJ0Q7lh2nviGIvkWH
Wrxx9sGoLK+/sl54LaULUlEgBo1K/8VxQDE1sXxcfPA/J7UsZKzcOZsHQ7zsHKgSeZuzE1LfdTqv
nsjhmJ7B4gTQ08P3HNibSX4CsE/4J+vFNirvIse+u8M8OI5M4D6dkOLhBVyjH+E8/0X3pXeiOyUw
KWGVvTeHi6HI2IPGYod+Dejc+Ta83cmuqgz2CrpNPWqDUmBI+jM4SZentYGui4v/XdhXwIOQ2vk5
MBwEC/MV42dO0b3cDKkrC7SbwfwzMXja9xWhWdj+4G5LwjyXpQ4NoqDRXokQJsUsYC+rTAr1dttF
LNmZozbr8dnFkoP/Moa5OznijY4mVGpCUv0EJyDtZdhKKEtsqkKdnCUzYTojI3GaB9MrdIMAd684
4Uw8JsrUoT+6WX2b4J2FwOJujm6nLMtBQBu3f/rNVO+m22tDrCtSqY23OacU26kXFW5CDWHgXBSb
j9FrdBp0sWwdpJ/nNV3M9JPbiOxxID9FKhvA6c/GLoGAsAiu/6ZtVq7DXbO7TBe52SIt49G4081j
shTvf0sU148gGWtdVuyreYJUJ9oOTLanERicbQdL3C1Ima4O6kDBdOhHGAL3dLK3MY6sc8Ga/RRn
zdLE9Kw5M/Z+1cVk/C42tJCG4PySpaRwgwsdXa9I5BYi3IqsLQEfPkh5I++jBsb+6DLW3ZLMo7iI
kfCoQ2qKjrXeLQ3Qb+KG7O6e7InBgCuyqERTqrot/cdGyWkQOJ9FaW9+5Z6grXeUJRWAfvCnyljn
Z4pXGsc2XOi/fNVBtw28dnaxLiQtiYyhVBiVX8fWDbp2Yq5aMKekWvxM148nZk6Ax+Fn8luNA0rB
WtSre6v6DDUCcZcZbo1lmpt69Yx0JtRd3nj0VziDttK7cZzB/SV0Zo8Xv/vO0UaoiVoQmYuQUVFu
wEYDtwxBDfRUI5ksCJaJV4JoUjaAa8yVpYB74maFDj3CtFNLW03XsDzSS4oStyD09eWXQCHfiGJP
b3fI2rARMGJ5HHwylJw/JR+pu4jvn31nvqA5w+G4Ikf5KXs0B6HKZErV54AMX0ugjVdlKB786Li4
nG4iDY6qo2J0EFoMH6OxSWfp2SxGalbTA1q3aYSBMS+SV9AZktvsNGTuTrSNwVYNHinTdSZZAfT5
zCFT+VFK/GOxKMyQ8fW6iPqrc3Uy4UKozLAWYjcjoOMTg1TeGp8SP1wKEXt0i9WQcpso1/VfUFMr
bM0vDHC2LCLHOoKagUkxd4BvmIcNddYtzcis3QO3XdXuEMI0iN5ua7nIgoCiSw/XoPNuwAmsjoej
baagVxhJqsDkMeO3g4D70MOl6egoVNwtJTz+GPE4496ZsSOXyiciamyzFlTfnf7C6jrCmimciVuN
kLavEvzMOVjGlz8RK/WUDamPBorh7QeqnPu7xjEx8+HMETBEtq7IHIlVdb9nPm9dcvQOYHUTGLAI
nLtBtViftRbFiyJaR04xe1JB5OFg7QGQRXLnWKZL1d9jL4AQGmppQJb4a4R1JZb5yraqB4WwKbBW
hPd8mI5Wso4itPqRGex00sb0LgytW4e3rVLa15SbmGR/RKiZXWB3ZP8/T2KdWiC2FHSt8cw0X4/K
NUD1bBYnheqCQ/FLh+mZxrZMhyfx1ikohqFVtKDqAvRD+QMVfQDPNPrmxRVSM0LGBvsVOYerlIxl
9BAPTNufwx423t9cpJQ3pj1sOIX0NC5NEtH5E/b4nrACZ5btoWR083zLZFUnZ4Efejws04zBnKLz
fvlrERWKhW0yPhmOqjNo9mPX9+wMARSLnuuwKz0PUgkK8HoW5H9zYr4hPeDs2DBQTPlwxumcyks/
BWcsRN557M9wcy01XU+TPdDnBWeEt+OWtPo11/J/KiDwTEIFj5CGAjkSd8k3rFJdGXDtYb2MVoqu
CMTrXqJfNGpH1rgeWfl7T5g+X4GDfaGPeI9a8dIGpGJYTOq9RR/jBu1xif8AOvy2r8CTVgBTHKIc
Nv315gSUlTDRtb4D3Af6EmorfRgUAxwSgC7/0sLtYeFcLP3H9ULr06VgQbA2WpRXqAA0pX0ro02a
h/T0xZ9aPzxrPne+tDv00B5zYrLL+AS51d8EGaKcqk6dQPYu2KJmohfBjJV9Ws16RJtigQTYnk++
LRwkT0YeWMItQdKSo0x9IEoA7pFTf69OWSUHtcqXax8lidKTqm8QoFpEuVVUDN7OfJsD8IPadvhW
MGt9OYfL5NWsjnLQpw4iEQtbio4PdEWR8Gvl6Xk6LZTpxghrda5YTkFNqRHWKMFbjhHS2uaOWlUW
Ym9KQbxQXM4n/K4EB6ryc91RcHEF7/rVy7H9jgfckzlUEp3n/b+7YA0m+pOz0VF52hBnYNXeUXN+
L0aQ46Ck8B7W5nzIpkGP36X2stXTxmAM26bOKDzw3GJwra8jC/W2N8NKn1j6h8V3NMkcqW8yvPXe
hE1I9ZrgFyt8gZc3P2sF32Y0dB2IgUmsroFmrIevsjf3NX4+IN8bsEu1Z4aj3nr6NBy8UbN1WB1x
Oznmt6L1Hjoa59cAM96DNB6Tq8hWjCe7EFi8UaMue8/bX3kJItIDCGUfuRczBR3hPYTcfUxYmT3W
+EqXUD3zvhuUL42/OXFrPH/SWo2HKj8Y0Z11tqMFVqLTyeWEZz6wQzBQocd0RXT+vNp+WaZ07w3N
jqH3AC7UhmGeQJCEz0jvWNTpvrDKgZtvjQ2FJvW+WfijJDCYb1iARzPuUlZ5VeOFbTPpRTJ1nJN1
6PcWlhboffqa9E1pv7vaqSX8AmmMYcis+XQUHMP4YOjhzlgTeuWp+wXirjZJXx2vaEwVi8403Q/4
DBwBBEGU5r7FDa34qJee6fZrg9FHFu2I0lmpd4KQJdzWAURWb9tfUzVoSQ1QgWd2gqvLiddx0rXb
P+U5oAXrVK0O/806OLKStkOOZag8EZXN3lEEp9qQdNoXN9OIpBL3040dwe5VgA40zbjuiYdu1W7n
VEyd9Lvs5dQ6jgJgidjfJyh0vdTYUNhkeg1i1D4z1o6YJs9cV82KYbQ/8Jey0Ka/2kjC4w6LdzoM
kznMX9Z5wxIyYaMNFC5h0MPggW4XHPrloEgqcpN935UsTP5s5niP+dysKKmJSnrHVjmxxt9z7uhu
PIoJkO+qPMwgV4Q54dM66FuJmv9XomiFtp8gfnmteXXwDUX/cyyBs14IGd2I2a28VNJMqDL9l6Su
Mi/lq9HCpSM=
`protect end_protected

