

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
MpZqUX7RHqqBov6r9sp19cCgAmwWMQKz/kilwg6KfQHVNd7thNhiMjNr9jWB5lhCnXS2Dmq96KWe
V2+V1FG8hw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
eHZEt9aF2k9bUkzJgCuA+q4yfEhMdqCEDNKyWFDaQseZ/ofqbFQAQc2uVVXTRkEXQs+GrviVm+j7
2wxr0JrS1Xw60RqMKKhLpfqRVe2BmFAKgU2BRL0PnA5WtTOSGCOmSJGfPa08juK1otVgwc2Gzis9
06D0/bVknfjjRpJI8Po=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
s0TU3tsqHiK9WgquIx4poaAXQ17I+2l5Vqn12DnbEwMyPpn0YeINJkDaKFxRf41aPK1Wkun6v9Z/
YYZDqYBgVO9Z0NMkbD4LC5C9cZSBdk4ezqdUWACnMS4IR+6qI0nvPM6pNZernzgmYtMGFsG0h7AO
2CLMNIzANr+bYhHkAqpdx/KPtV7Deh8xOAkQeNSD+8rjhU0z6Gg+2FjdPjkTgWwsP8xrTSENuxiw
xPh+QM3dvd2tDQbC1sSMu3CzeLQh9mMzJ/R1uFQDv4VC1TFFFPI7VMPMlrl3y0ondyZNERO3SeHy
Mn6aVbKjlR68QJuFwdsz80LSh3ZTJ+foTk16ug==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
uIfIqnJL93Nk48nDUNvQ46MGSw+0jZe8QEp6D5vC3ytHCm6yvGspxOPTR0O/6R1kGtbYGX5AVD6b
KvoAJRDP7Wr2E6PTOWfFxWtEHCKiApDz7UksHM1gqF0d7SCMfsYR0KKn9LnLJiQxmEJD5y64ve5y
9s0qEeMi9k4HxMVPc9k=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
XH+fS8ngHwfDFxF50DT7MdOHeXbY/uKmg7Eva1j7eQ+2X+a34Rn17d34wKLf1Z56AIT4ksXzo17E
WT5KT9rKAQNao71yUm+YQAunOwqKEPRyxOz3bb+3Zvx3y9p+F7xTeZFLan3KtqwByX5rGkNJtGjN
oI8H+T5FEpTIirQ9oxghooMSVVhKX8RsayssyrgajR3SSX0Q0ggoCOy3XtjsFKfrcDNlt7iEsMAt
+8vV+volJUxGGSYbt9ATDx7fk+pYKVnFR1jV5fEpxyqiZQoGjkjsnbN29jqgiZBfhyEe2uAb7sF2
RnfrEGY96pFoR0k3gse3XEc9radVftI75N7ROg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5808)
`protect data_block
HXZGXO4sbfKIaujBmXbj1prb9v4Z19I0MnoTx+Fud8IRWSlYHVIeqBGMco18CvuMOTR066iGSOYd
fawCuo3UC7SG8SM11LaI5ApD3HzkWmhmc5SWuQpLzP2ieSghmkSdE5PZXjznMLfViUWYjl5o1FAR
LzU2NOhVy/CM5xicSFcWGT03mb7qOg5dOKVXNmjYJXS4e04EJg8c8+FqdZ3LcQbF6ZJOJfEt4fHp
Uxm0xgZptfwi4nVZZUoylEURZb9aZGhMjcqPCm5TotqmtNQ6A3WIYnelqlaxairSkEGG9PTyDfxP
Vb5CBtG2lYD3p3GNqV58BBwROwaj72TKNek4kotBFvfTrw97ou2WEmZpDXIRF4RjLHFML8wiH+e2
b75GTsWlRK0VKeC+y2eL1r1xYRacexaTozpYk2fyPK048NmQvShTglUvXVo1lI64ibAgEzjol4E3
/aucTGtYeeIMWwD+GGgteVC1+WAoYcYogUgwfbGdNmYbl224tmoNHFkg94KiIprxsiV/GUxfHXYU
G8Tnqwv966pkHigKb1DXHjb0OvzTjcGGLqFr+YAFM3f16+f5XgYnURQ0GOfLyjlnhYppMuEtBVFd
eOLx9x5JgS1tSVnZL97c11tHXxOLZH5QDJN9ucGgoRGl7Td0gJJxA2cgCUMgH4ZCweLWi+6QGDR+
ciKXjKif7e6cdswiMF8vjrBd4ot9wNgUlT4U1VaHmnO3rQ5gUs3iADuc/TqDlYV+rSTpqhqY4iBT
rnqlru4jMOILpiftnNVQ3ZMpylFC44viqiHB8BkKsE1pHSABM2zpC5CD6j6SF+c+v8JemFRE1DDL
768vZ977UV7srxGcQAZNkmHnDkBYq5EZ+6Tdt7jZ9FHLG4GIinl5+9yJA3AM4uu6rx8DmvCaX4Z0
54aYTDB5TUIJIXriRkw9Tw8HTx5y3rlpvn+iUnCPtom6DH3BDdXo7dwskpLE4Dffe8IKL0kHMNMA
6ZRfl/HZRrpZujYA3+BoYI7XMuprnRUOumPBu7l4tiROO55v9o5dZPx39Pxy3SNdZ3oLxR1zH0x9
lGrPfCfZRPnSUU+JJWF1EAbtDWn1aDMAPNoV1CtCH4ZdZiX51PCntsabzqDCQVSQ1zuRQjfBsm8p
rJgpmRRnc17+cQj2jgO+g6uOUtRkEVQnwMbr3+1RRY2maGAQDJIUSYJg8i/u7XthSDNnxXHcg0+5
V4l4cNZIPhdm+vz7vW9mAAL4Y+xB5Oag4zPx1DtVZgi/xSiUUV3ODsoddOKj6wiHaXweYf69xnOm
KPBfCXx/0aovP+WJO1XFNSu24OrGSl1Z0bxHsRpJQcj8cyet5BTjUdJxgoSazxaaNswnwoYGg8x9
oidXTaVR8Rmi3+i/BQzL0xkn4dSrG9Orv5g/5M3NyrjCw58sgfROKUE8uwsmnPRzdv5iMbAflVot
foRPHzGaBSQUqtmDNsFfldjP12NFI/4JVJtBr3NlNvOltQqS1M2NHMm8Ck+sSVPwrnGtAS6Wvzei
7vL56bg3N8CJwW73X9R76PvOepem2bT2mcBQedqIR+sEsp6BPE8OLbFfObCvmyyd2+1jsos2y8yP
WOn/HxFHAGIhPYXy/zGq+S9l/nSKzgpRhlSVaCYFsRmxAnB/ekVfF1qRsMYwgZzk1A98xV+i+Ie7
3wEPS/0GUt/6iN0lhRDPIv8yj0E/5d/rgbhvJjX4hNK2eLv6gK2V/kxniXAIwhoFPEv+VGjYdNSc
QHrqItNjz9IMH+5C2xBqG+/+hSufEsf3uTXXWp//GI6qNI/H6vel+boe/XF4T1InI4xoFy7XbIAL
0CHhxCIjx+b6qBeu6lVla7VbIEvz7EFPF9hzbYeb8AjXog3GZf8clu5Ze828aJIi6TNAlYQaBgZ2
EH4S4f6djf72PRLgfHYgC+uVoOHsXVbGdmZXWJ4oMDwVpKRkFcexQ6vjvBtrK5ABmwEG5+fLx0mM
rjNEyr4X3muJZSbzzM3rAW6akagL8LQu9PSvUVzyJORHtZ7plOBp0aA4jqemWyrJyXIE/PEV0For
VROy7dB55XSk4KVRPLQ5z1b4w4anM9oVTM0pfD42MHNtHjTknmGCE2FKLFpWniRPi6Drds1zaTKR
VSFYAwX2YoGNuv5cR+OVzI9a7+lpBfw9bQSZpCm3CbUdA+h8+RoxajBpX74uBhnb18bWoFZl4AFe
F7k2jpABoYPW6oPq1+w7noEUrOVsTpEP5AppVStQ2fqdOw1KssDs/f9zJmWk1Oo2QDjnhkAIRk/p
Mw1Yv7JazBCg1AiwixrxWAH0X1dzt8k5MhG7+nUJ4bUthcsfgh3qb8dq8/SKkirlY0KZsPoBR18J
Eo4s2IFUgSU7hLT1864HLJDkU12FTuOxC71DMkX9qoEh5hNumBIurUiWQDWmSgjdautF0L0cI9qJ
OwrvjukMLUPxmeTSnc+T/lcbfwbDRU35Q8W8E+gbDML9nWmdxSq8h/q9VuKe1+FexGsZFIk5Bz/O
L9qeB0g5iB7vfzuQsHor4wfA/AnIwzgWD3ZL1rcUygUCVQfQD/GfRpuyY6S9NSyYYHlEhiFkio4/
4IHKaa5aJ3NPzmx9PUeYkOJaKgRFp4xSCDakF96JHrEE/ZH6WJO1vz455+Yj0sFx8EdegMSZNKSH
fu3ouuEyyS08AjgmsIg+WBKe+qTAfP9b4vCgWp8Q4a/TK4g3KBbMkU1Z0aXGQW3Ui99pmXpxH6xi
HXZIHeTfPHqpsuMtxWe5KX7gZmPn46arx/dJrSLZ64rWfbh6os3MHPJcbinAEbt0y7x654R2raEH
NwKKTXXvMf5kl9UPmbNtO1b+BopJtsksRMKdkyYu1bJJWKyO08ULOyZUF80WGdbaBsw0FBIqovHn
83IaOVgKkslvucc05a/IljfjlaLPLr5H7AVgiStlmndn11aXiFvxQVn2mI1EsVhW525Un1/tSoYR
nOVydJusuEkXcyzd6qaJ6UC9gLVQXV+Yk25N3wB44kpAzXjBEoEpIL8Dw7o5kuWeXo1UBLT8JLfv
39op9/bz5foA4iP4zhqANOQAsOxOvLUp2exUpx6wZaYw/R4U0+3MQFXOfKzUUOh32q9vLbfppPCK
dfXenXkTDC8CvV3N9Qkx8BE+GvhMyW19IYgBb3qsylVygCCXk1EctR/qHUamFBSg3UuywSsCC4Gq
7ZFoGn7L8T3DWiEJFHLJwJmVj23yHUEpqsAv9N5LJI3zNS/oCrA4t1gZ60H6/sBETMDoA199XYKW
yR9TnIu2GIoLwr8LSKnX3n6iA5XfDOKSohfAT09bVf02IVUjQWbgahRHPQLtBlR8LVl4kxqwSZuv
kiJ3yxYGuZllCNh8AJMRrEvtTEfxg7o13IDY4eN6+dz65JAOou6Ud3toj+OHiB9zMRkhGUNQJKNR
+E9COpOBKUTi7sMkp7YGmEH5ZbUk0ZyWY+668z5DKwoCRx9AZVG8xdKJEzrhuJR1l+OAkG/SIn4T
lYp3PFYwQJBlxXGHcfeGOuf52Gx2WbXzAunM+UygYEUps2MloA6H5KQAVIKmw2+DQuXLS3kkOQfH
/l68WJI08hHEiBdV/DIZH6dmU+1lT670cJEewzkVqSI/SQ2fWagHB11oY1HZDyPHBOQedDQoDzeq
WIju3re+CrvuOXmE5CxG4bXsUkvZSHSy1LXEwYNSG8IwxnJFbjhrk30ybTPVvUUeBacJ47SH7kpr
gZj6QYgarCfogrtl1TdC1g7CHH8Gt3az0z8OyQM9IIi1NsX8AWxQNFofskCt8XDQ2tI/u7uNUKEm
mvKA/qCA6hz4HF2zPJhx72iHn8oXCeaPpSMgk/Zwrf8ZFy/xVnfY5AapGlWZlXJ7zdYCYHzDqrpc
4WltM4WghyIwFovCy1c/lpDEOn2TMzjpCe0Y6GhY2X1i/BurRr+fpccAzMCaNlhbM7HOa2Z+/B1B
TaeV0AmdAgwulB4V0LNzmx+XcST0jVX7eY0nzq11c4o89cQ1fWljgWJn5VWUL6GLDhQCQHVa/3+k
jdZLkqZ7wBs+mQvQaNbqCILA90UmVH1c5x7IMDqz44h+0+xfv0IxtqLseoTkU0LR48hhWFuSda+7
djxLVHGqaGsuibkR6z5jlR7f3jo/vVPzB0lg70cjlweEpUGCWym9lGjYcPycD34EhFwix8bBFZqs
GObGM+efPzOZM7U0gKvSdyU4KQku/A93NgvhavxVN7O4eqI4a6296SjSuaV6fPXi4ZbIJqosCJvb
tn61ySNcK01VkJBIIZiFkm55iH111MOHzt4uCleK/Y5JD9sP0QjUzxgRryU5ZCkva9z+NO1sll0H
PNaSVPdC2Bj9rYgbOVAlLi1bLOgq/QOCEcw/crEn2wzQw0yzt3n0yIAiruoCbXyb12ONHWrL2POX
m6ggJFLu2cr6v48mGBKHrnijR96xgDu2+6wlRIMdTORIQLUWTRhSOOJWfi0h31OYrvTAHlG/Orhx
fB8Hz8dFd5ihTUB1AKJGOeGQ5Tdi+PpJs1nJTl0L4v9pgAj0MRljzQ2U7ADzrEmP/t7JdT/r2YZE
Z4Z0qQLQDIQX6AnF5cXM8znYyoI0VefXnXd+0tXj3zENhLWZ1yQLjOK/FQED5iQGR2MCbqKBbMPO
HQpZp3lhPAX5hwFpTT0lXqDnrWykN1DYqRxFlrRzovcqzlfUsH7okY65n5aYYDSqNKTDt8hpODn6
B/vzMT2jMFaJbVHngkLyMSgojY8qnk2P6Ej1+gfv95JEg8HLpaDndITvH1+tG0jIZDxjMKYqEKej
U1c+dShYHknc0e2sfcu0U2IodAzOKuQ0jknoeoF98c2+BIiQ4KvAjf4urpKcEuhc9doaHTBGoICt
yhiHgIUwbaY1P9k0P5HYJrxoVSVZCGKOk0RRlAiwdPdHSc6QAs1PyH2hZUTse896RCyXcQGgC35W
4HiTXYucsUTQNMKGn4D4dFMQ5AbnOuv/DdoVZcUGAWTW4oOAsP88BypQE/ZQSM0XpyxM5UGhBRHM
5B5R4MrF7oNbqbex+jlb6JO7k8kpt0mCIKkZlFcgbK0kcpt4FDDtiUk3JnEyEc//c63iMRyrTvKy
ZzbI8dKTbpOJnGJXcl+0MlmbwzNAtzB4Uu6fHTuk2oiMB2Bl+CIU7X3g82o9cXy21XqsozC46Bsa
O7dx0B0ORuyVDKW5xQUz3J38+GhvUnVWptIy3RNGjNpgX62vbEP1Il/AnUd5KBSHWLH2amU++Z9G
fJ4p14ocz8pO2DzRidu8GszaXrYPosFnypI8R6zt3B0ClGSouXW8OmMgdiRZ5Hy2KC4ag+Dr/gUx
OHFKGtyC05qQnbpFF/bhHmc6VWiPSfACDrWTw4E4yAXn1/VMBfAPOp+4JYXmTeqvO5JTGGidlrtB
tZJfY49z9LBlJ31SWcteEJc7yffbUQFdaxDvRDjKgMRoTJPG1JcgmZqmDBM1hdqIgm6f39LvNvgE
1VYjgv5+dYLob4Ib3nm6JnlndlzOE4EexpIYXvMc+PNQNo8+SOvh33cv80Izl0INMPqz0qMwLvR0
xfIB4CEgUD+wzJoDK98b1BHOP2QAnwpX8Xd/v3QiA6CqMLKatzbSmSPRzfT5KJ/0wGot4HeO4FgE
Lkcd+tD1moLkvlOei7kJwXKTbU75LnaOG86biWBqi26IUyXhoBmOB4TPx3k0Eue5WJ7gKXXAA3fK
0PRnXGs4YZ08GjYw2h1fjlu5DSsv8WZgwB7TyMi0BBwbqI6HDRcrrCxUGx6+g0uihih5J3UXZI5h
/6bUBMpX9H+afJe9U+j+Zxpj93YHVN3Qnib5rnb7ezAnHkFJB9MpN45Rez1ko+4qJ0fPx9LvUwTS
dcYSoJv+Kh2TQ5tzfn6fKS9EG3nmNqgt8uV5uGRFbR46wSZ4VI7X9evsqIhMmiJujb0/vNwK9zhl
5ujaFtxh+aXbLNVcQYAcBnv2E8W1fnou3IMqSwpttigrlo4RoT7E6hsUK+/YsbIqro/9959Dz937
RNrApC9zp3mFP6QGK/tTNnQaQ7G1yfNVPSxlmhO052zg9QWnm5p4ComJv/NBZONARqL8P6xeXPos
9X3IjG0t2hJRUp1p5zTde0/p2sGT6rnYi5S4NjPkyLAj0aAX6HZO2er4bMkqXB8Hv0yfda/Cfoo3
cfaI0D8WC32RbT2QEXdyEuFsLxNqo6fvomF/VpeVTgJjHJOSurh1NjOIJvWq+8JioPYCmz12JSxO
vAWW3gOW0RA+yG9TytDfpaGf2rpM3KPRzc6IV1I/ZCPb4/peOR2NzUnL0pSakIx+aRMnEMyAq5ry
JdccN7jA2qJj4JGvgAnxXLGj6Hv833EkThF9h5bsCj7E6XlJ2C2ydoGLgx0MRbVQD/9D0Iwbl0dW
m224fffDbYd8Rg/Uvx8LYg9nvBS6+a4C9sQ2ZMk4hdOQx512YbKU8N8lXxEfK1jeXoKqE4DeWOAS
CFbNDUgITTaoZhxM5OZBIHq9zas22khGJoxwT8VduwKi2EfaxrSMvLywvphGmgkwUgiY+si2Qf93
z2MOyLC/7gmwskTY/TGDINN2wdKW6rxD+3QqRD7MxzmjehS8HQqVeWZ73UV7IEISjkmtLdi9U55h
HU4Io8xP5DrxoROVd1aEO2M3Aw5ECfQEJu6NEKjDZe7pYrGvcn6lNuDWb3krKxR0pxpTusCvBTSS
yeCjdVl/Runsk6bH+JGDi9j/xt07ZgzkNsoULPF2ybLelroBAmLveeNQhyfL+1WfUILVmkj/EiwS
4iNx/XlHKbVy7/3KGIDRGeA/uFcrzg9Uv6sa7tdSKyeTgX32dqyx6Vi+B4OTC3+KNzP+am7uSPyK
ezHEp8cDmJ8x39RBxV5VSZfGT6MBdMkjvL/RwzPA16ECWQoUTf4rlyr+IUOnUfEvQwuzUVWWrdYJ
nxfifdQgcaOSGFqomoqkH2MDbtWMqmf/6cPsjnt8pUdqwNa0EW0HKJg83hnUrTtx3QEkjjsSiQ0b
fV+OJR0gHztyY/IYFVdwMG1HxfeVVHK4XZ6lbMa0QQU6kNFMOzRYbdNSOs7XCYSuSvkb9HYVi5/D
Dt2AeUvtRSgLVoLODzk0Mt23hMasJgCK7seEpaZRG+y/Njj2j2j1/U70uIb5gf3RF+lNAjHKSyeh
yxN1QYpgXFdO3etdBUEsB8M1ZCUpvHwin+6eRbhBUM3s1m6+rTmiW4BU/uM0q3R14BDqyrGyW2rO
prCQJexMGW/LXANMVjqLhpy41g1wRoFZ71X1/0wb7k9vnWcR/DndbcgSSNRGr/bdO24Bs/eAsXeM
mhncomjHBfMiNWnjcfoG2jpTGJj1VBVN9w2CBVF11NVXKd5/TPIMO71WMZycpIa8f2s3bsGOl5fi
kj06Eopty/7bx/3IVzcn3spJo8JA82kDBOoA4vd2SsiHqe23EKo7QT7r82Kzb6tX0T6pj/lJ5lrs
YkKOrPMvlxsYGUAxE3TgU3l3nnK3rKTM3KFrNRDE1FCnEkafvebwalo9qUspchqovE+QjCdmHC9R
vv5D/FLLiLzkrZSlXjMUI5qr8PemK+dSLoLvIUO0b1F1ezZxfo6wlLCvuIqh4Y5D1pT2ce8BU2y7
/RDtIg4Z1Tbf1vnlG352lkHC4MlwLFFXXA9Rysnd+ywnq6v5xh7AAw12Jd7gvdTQYdeJxHsm7PZy
on/8uPXjQ5in4yG4ghdJMj+z3w5qc4B4cWlJLqQpNgzmRE4aVhs/I9XVe+m+vXEJPrAh
`protect end_protected

