

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
IkKQ7UnyfG/i0Gz2KESfn5rIa2XG6JjMuNzaLweotYfssoXFPRW5MF9/SJXIBGc5jwrrtn7ZIvXw
ZMKFyJ3FzA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
A7z8fuAKplZhDCneI9mNA3lof0N+J7iQN1H5R3Mj6yF0lZ6gCWQLLnnmsEoxkSX05NXSzlh4gcEg
7rRfO6LtEEhf+XGNB65vpBYpfhGyoq59NAHhGVo4SvBM+mv7uMxOGdpTeOCZ4JbHV0AkjL28mjov
93MegfTkvdkm8J0Lvdk=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
xuMQUwo0GDzI3cOEq+tu/2nUcDmn/7fhQTHPWWNseJwSS2v3l/iZo4evCcnhY45ESTueA+ZpjAko
WVoSIubelzbNSlntY2uMGs5oczMZtiztniKkMtgrjy3EW9dfGbHhtmNrOHGIHH4IdMr3kAy4Vh74
ZigAJ9A6+7kI6MsJi8v3mT1ARZHCR6MWsQMcVGsi2drnsGRWoYryCO5xQR7B/cwBGzMymTal23NM
pQKOm5sZ3P6n60ZuBiOsJmbRp0+LVYxKNhFdxlNXd0mwyAZQT/UOuOuVbjlNnKY3+syFmjH1X2jU
BRKqD7PfkYIVMVQ6XvOwQSNLyki/t/1FG9LntQ==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
2lTj0FQ90PRwxkOhP58Pis/0pnBIhVIOGqxXo4lWUDsJI5sRS1Q5L+Q6i9o+BNlX2LRPYus/9Dnq
5ATglZxA4PDv34H6B5xWMxj6PrHSWzf271mNIoMFrjsSBdzp3H4BqkwksoU2N0BujU4mvFktBj6s
VuYwP8rZjGtZ8cTr2i8=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
WKc7lQN7TOvrS4DJ7NNUxP98rrzfIQuz4DIZ8eAY+GKFx6NuoyinV7kCt4N2qBg8IRnkz00LUdTl
h4FZuBrLJJyfOOGbqIiZNIhgdqVi7fXcxV2ef2SWPHLvr6kIV0N1TmRIBZht7FPZCej+/BNW8QYG
B1Rd/mmsAB7hXx6GfVQ5u7NRsVDyxlcEghLjiM7GAdTaOWl/F6pDM3aRwjjOmid8Gt7xmiYfPT0B
Gzk510O+OqDJRqmdMvwBmv3K/y+M1RxYsLOpwIle5lGrJoXR6zj5dZS3g0EOtylaiuYJczAHSe89
8ncn00hUVfz/5JZCkfgcxZH1LxGTI+Ly2xY+5w==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 8544)
`protect data_block
558TeFkw58K0+DfX25tfPGjF/TyCGjJdDI/QAeqcx2rHy5O2mfEjB5gYKlP9sy1R/BjaLSEPKZ46
34OZG1vsDs8UHcyl0UGrG6TtuwLUCgsKmUNYF2QZHBRaZcIzDN7k4JLV3j/krzXjAQtcr7hNv8cq
F6LVMpJO6dqg2fK31oR7mY16+Yom/XgEne0vmiFiW2UsxVfllOsFerWh9oVOHURLbfXLIEPUQVf5
8y8C1bvQnZBYakRpWrFxg/xzFOT9MrMVLSSEdhzIxfzXYk4uuQX69GhzavLssTSfI7fxZ2w/6WdN
OsoOfMfwOCxamYwl/TYG5yPxW6UkzjItJeApZLuPFQDYG1HlbeRtPiNU6zVmDToUQO4kjfU3GqNC
9lcZJO8OpwHcBTeuq+gmUY/dzJJA2kx6aWh/ByuGzrYV8Ol8zx0jPr0HG45ZTBudJIsYvzEUM597
/A3b9oCv72e1vUd3PYIZ66bb/esvFASSYctwdgxt+mXS1R7LzLabTAa+qo3Gy/zQXpFwA2nZclo5
wuKLV1/H+M5F6qc3xj1GKa9BH0hYGhiU2w0EsRt0q1ZWYcAtqjukRvO37RfrNo22MZWjKsCscaXR
P3UmnJSRMfMMrOY7x57s2d3NDKbCDpv/tHBXvYmA9gevT2BDNlV3OSgzA3IVtzbd2+By/qk5dSYc
pvuI6bki8v5Ecis/oG53pK8YJ6Qds4QQhhcXbh5ijNVRV8UNjAsEo57CTUExdfNZTR3J0/vAMKZf
lnTxMpAjIaJ8+IxuPJT1j+1IGgU+sxdDUCOOajNEt5dbOCq7TEZ2h0l7qLj4LF+eJ0H06cVcHgJd
8OaTlNx+8htki3l8qCm6SeERmjNhyAhQz+P8jBIlrehklalqXgj/97/jnEQRCsnvWuiD1ZKcYW3V
oLcUmej+e2PgNbf3wCaK/OVqL7O3GNSGy6N1BzR/WfmAGq9zcLf1E8yAutvQcHbk5s0beJR1Dk14
kea13ktVrqkdxWwhvaw1VhjnJD+WjzN7Udo5Q0p7WO3NKYFuG4cIyB0nlv+NZet0D+WUaqut90a1
8fLl3hBmiwIUaWvWPKMXoZIIy3Drc1PNUaibQN98vUjYme5bCdBEFTqj1DAJMmBpu8Zg+/WniSPp
1ipuucmeUf22kU+vjLZTQKj/lMpL54u/V6DRB1D4DYPyJn+HrKPAyqrzwuWltdmEHNcAh9xvAhrE
yJxFcYnMfvzge0N5Paf+kDF81t7KjfL4AbpFbKchBY4PE+abcg6oOpFCyIwcs9iKONctojPBgCZA
gZ3iBcEac45sdJeaNrV7M3kz4sJbvccJ5FsCpMEqv6DpDzoNw6BzRHcXwhVmP/IBQrmg7RzCN3gY
C2j3SBaouDrF/8Nq+nJv/L1Irjd1HmQUzglrvfX2fsrye6ms2o2QbDwVbd+4hUChrfK9JRiir1WJ
+N95jkwkxywOjrJyHn7bvWYRAiSK3ufqWKJb9ZJgrSTi6c9ygCkJ8wUlV7Pf2rSAj0ZUFPRub+H4
Rw/BGPN5SXG51tNN6/OISI7alFW79Gis+Dor+pwZRTfcQtnKqzPLGPrpQ+jhgLzCd1hCTJDQmM4B
90mCt8zyYlMACTc1x0WV/KTKHALRzk+gmLQUiT+hiCQBslHY08xUBkFDnBIGpxnJwcqE0iRpjPVi
6AER4NhoVf3oiQQE91ypjM5QStqP2stfObMbyBvMBIbfiIlrauCCXRsxpX9+hkmEPV0SlamdhcIu
laiopsmi2mESeXQ411SmLCoyrnOet1oGwD9PTRxVvIcfRQ5M8rguarNr2yla09JS2eaDqyJ8k0O/
aGBl9FH0B9R10aDNLeNBGZJe50kL/EWGl3qLDttV08KpFA0LhblAjKZpqCOvYifjGTDZqs4Af4l1
gbF24pDxV36U6zQts3xxOhEaKcXmgg8AeU7dV472sg+3e/UrTrMdK2GbRBucC+gZUjYAdSrTPHk9
tnTXpJ3VTpr+hkhRWkUIPO9rDPufhojdMlaTHBmg9sugdLPexRoqvqZNp1XG9/jtw+RBY13wcGrL
J9vsBy/qTSa4qW7iDdF0bT823mJoJyyO/IBxdlRXF3HS3C8Gg6STbCal/VkSO/xF7EFjcLwBWFuU
Jawf1H9qpHPAOPP0aCbDclvCf7o3SFyFPGRsNRjH6SfoHXl51aHC/yxTZg/sWNpL5oTCl3eHuwYv
Sy8VgaGNK3cvjdVWk7mDBgA7ciIoNl+66SYQYcsOBDJC9y5nIE/Dlam/t1qs9XLvN0mc5CXqRlXP
o9mPnT3u6DxAhmZMLFwSz6WagQURvT6cu4zF0iXD1ZqVcIcjlPy8RULSx+CB8Vw2ibLtGk35vcOE
kWkXfer1yI0w/4BEVeLfpQhkcn0bHHxt+jV+80/1adBG7QmY9pFNRf5LbP8k3LrT+EfL2W0GsK2+
nDuvQSvBy+uRP28SKdIqVAyA6+U9pgnuYO8BU0ayoxudYvSAFIzQDHulh+5a9nkg0pP+tNolgVME
OgiijSe+B/M5laixsnCx8wH67TOf++N0BSoe/j3HvWGzvscaspNk5BOtaSZZNZRmFCZd2KKp15zz
d2KP8MVzpfSi2LbcKPPtOb30YwA59P/G6ZXFdrvbEVA+enC/40i6xfR2yttdmWRyVw7SSkvBL84z
6vC5rxzka1TraBEh+/MS99Bk/m53xv0v3mQm8btQxbg6fFKcE0G2vNhjhKRMkHM/bp26p91NE0fO
Hw4P4tTp9SzYRRe1GPJEM1V1Uh06qumVZDBUoEgXKVSwp6S5r6z1XOHuyWF7l5GgPzAnWEUsc/Rt
HQwGq6NoiV4f7vH3AeDAogD2A2iSqCD6WLh5Al2gDrEtohKGlCygVKrbe7a7Ut2TPUo8faFi99D2
sip8NWGfGXeA59UjPS+v6RPSw9FsFwIGUf7dBuFpM1TKaz/hpC+aCofKz4RePCQE+WJ+Q1hlZGwR
9BNwXycjjMyMiSmWhMX0lkpYZbno61Sp0nWkzR8186olWuSSJfbVsIoIcfbR+T1VoFbIjyttgXlB
bChFJqDNCb1OrUdVR3Var710QDViEmrx/ESZnDh7wRzPr1jyw5lBiJn10IFCLliePpgB3fpB4Pdz
1pT/2eozpR1bPGl6P5JJ5D+rMUrZDklM2iecTCTpKwqKxmMae+4WVfc/vUNuQeIGMZNhaj62fzMu
xaAV5XuhEBAQghBpNKEOuLwWc0LrpuVGQoanyyAlc2JrbQVKxeHngtg25fBIC0f/K1UW+98weUEN
Z62mAEXUwEFBhw4S86iXtVam7pb3dQJa5nTiqekGDgf9v4Ve6Tx9QFr8VpSzY94ULx5pOQLeJJ8A
24NOOs7YOAX+FjCZfTuc/ZcHHz5bxNuVqw5TeLnBd+Rfu7QKwAGtbbQpqu3HzclKulehK9FY0sS9
5kQA9xDvp5UsqyTDEYKjOXZFGsGcvWicQRB6dp85HWA7xLQ+NFvDJ1vg0fq4mqgPpUe5Pj5/D1Dz
xb0o8YGBwoG2vkTB8A0kkf8AsvfWj+H61Niq0gOM5UOW0hKKIcwKkO3/IlbygwQ5qfkzpbQlA+Fb
B7vI/cLidQ/CqAtG9ze/1onRYkHT+oHr5k48DJxuycQn0v90udNgdOey4CpcgaEollAPTPPBpYh7
79j4uDLdTALeqNnclKkwGFqMHpjn77etJflMZQRzXASKVDT1ZhjbUwPYY5N+ERGkg7szlOlxItfY
F/Zs6yLMR5AdWASy7S5RoviMl8WVhKRP6MZZ1kBuBwvDpM+WxX7PwRqtVsvoO/ufvym7rFoI6VIZ
CbQhKBWbO7fsACwsBkGVxuF7i0+K+bDmn5qySiGd+5EEbGLugg0DgLb8G/n6Tc7wRR2lnwvthMql
cES+j+UpecRG48UkqkqlYs2Dcw00YA/hs76gT7Yq1hJFfUWG3A01Ho7poi0+NQBtEjmGLE1N0afM
fdLc6+j66s+5CTRdMcIxRTQPjYAcAepPLZDgWWnBiyYhhMvwAEM2gp7wyKryxby4+L5b3jx8SSuI
77VL4Dtzc+eQODjpY172uR5aDB4T144G+eXsLrd4YfIeE1oZTl56Bmh3MnaYOZUV/no37abz6oi6
RLOQ7hTAr2Vr2Cn9WPjpL9vwjmLIoTAgo2QHhEx/I2LgEatdWBxL30U5LZ7Dip3C3py20xF33vfe
Fdl35J5/PzFk3cUqic94Suf7haApBjtrUhP2CyPDH3p10GZUk30rxeMV872OhpuN8Bz3qrJ9O9Mm
XkW2HG9LCwEDoojFsvZ2xCk9niVssbxrL6Q2UDgTY10flrKgKVXB2yWXH9aU1fNiudmB44oOdszk
cwQZDtnQ3b7XcwEF/EJNUr/lZMxCobIKp8L76NBjdOgG0IPf70486KT5unGsEKW8c5bHOlqlB+aZ
aenihjldjHJc9hrzLhAkJo+DhZYSst/NVN1WstJ2zW6XvHM/bAmFaBSu53teyESiq1NSFAOiRf98
qlMZZElK5Q/jN6Rk0zOshX4D2ujaVLoPKPKuVd8tcEh6aipJ7rbWOJvCePTtILs4z8FdX4RwPjQr
Llge5bYRwN0pkqoqzDn709iP+HRieJKJVw1Cr5kjGUwg/Gpbn9Yv8/pxD2iPOc9DDM/jfZryr8Q0
RzxlC30CH7YdBEzL2W1Z75VS0xKzvi52XvTheb6dilwybFiAIDaX65K+4uc3dytxTgCxf6Hjg7Qj
iuh7tMJmoOt/YsLY9WnZRRvktQBve7FUwWWXm1ZBG8E9KIHvu5i5NfkRTkaOhbcOj2+fBMcyWVE2
Pxr2puvCYOLM+0xxH0mHM7L+3GR9f9tjvHcyLrBGGI2fv6fLSh3vo9OHF4vm+fTSXd8ZPWf4ItG4
wi2dDg1s7Se88pPUw+sCXURk8BdgF4mKhUvbwkxd7iBE3qazbdB6VCxMZFqtlhI0sG5i4fde8pfm
T3qJjugeWxJQn3HBQNJLdV6wXvbDnjQJRdjhfdo0uPqSBswZrwEiKGIUBMbACB3rs26vIAY80A6L
FIK0/eGDaCjtB3LYaVqPcSYFLS8BwSqXKr8t3/rlRvoB7Vjb+Vd7AWenA6rWt+RuJW9gN4vcZ/Kf
B26wUHeH0QjfL11GyvNd/gTAW3R4iOiz0AAr9DtdFF+8iZSbEmSgjlORitIAx4b1pDuESJVlxDwN
bjQqppRfPrw0cqvT2lILgxyBsWHGuT5bl0jc49f+QUSdpPqT3Cn/iDATAaKtsnhDubBwYYgKu2Zt
k29G5NQkEkMUXfl4jvt177HxHrxoABWdvz+bky/puLANh+2h9DZNGQOqQZKWJ8Z3Hry1Pme2b2TE
5QBqKX/6dFYaYBmKMSU5el0nvhIsrqUUbGREHhhhF2alJZVEcb7nhyxJgim5LGSPNps0rpubBCbX
Fyj+Y+Y27WH6/Z+DsfwAMldAlg1Bci2OIAXQPsoOj4wCpntutAYY1M7l3ofSVFb/GkBxgR8n9/0T
lSmI+/YTC0MdJ0mlG5VmBMzI7hfI+rBwHPAjaUcxJt/BXLGf834chTdUbYwK3bCHlYyVptvsYJaQ
ox16xj51cMKK5V9IEHniIm/g/NYdBzAlLn49116NF0CZRpAg3YXX8behk9hOum509jN02Z8X9wBy
zOf3gSs/8VWJVksLzAKrsplp/AG/G/+zHk3/Sc4JtDO2WbACESkDfxiXhiUFm6L6RMFNCI5g/L6g
xDK80Yx5aC/F5OoQxlepnmOH4bXb/POaNpsfMtCWpy66T/dMrVpGSxEQXHcekrZhCSY0arayJGfq
RPOjGkzCXeDf1a5zWkFAioW3ubYAyby0iwwz9kL7XEqNld+ES2ee3bKk0pmDlJPos4bDI7dL2u9E
f4BKc0KOWmtlCXKMCQk3fiB3SwAAYOJ06/Oj0aatYDj53jqmG+Xetat7pOkEMKeFKoG9MIUfHQWq
UEV3AL2xoI7vRmb7Tk8vFiDpp2ldD0RtTjlIV/TAcoAZZG3QEmiJZbG32WALJsGcGNngkdUIrAHL
jbQMJvm3DJTO0PIkyw1owb4WzxPMrNrQKdEiOGLPcJfdlWXevq27dMAvEsuVhXnlinndO24tAaSW
KEBEDqgxGKl1I/cKCDufkMD44wGN2+iZ0Q352tY4EyfDSIeePZbpnauua+17gh+yAGZj3vv0hBVE
89WZh8MiSoiELFf6X2J3E3dTRIgMLx1SYaIQKJEt3XB/YQ2+gOvVMkwKBtNcLm72E0zMtVLmTqVX
14cVvckUb60yqdVf54vPG4P528IUEB7/XnAkn/OOw8K/u7jIr2kJwL3GPkxBrOWu/JLYMjNHcCzR
gfAGr+mxpTe5AHdgm1ZvMPbtWpxMZ14R6vQBbZlaewK76jz7Iz8Um/zEuH5J+3xinLhS9goUfzhP
XVg3hAanjqRIq1yGH45fGfaxeg/duyCeJP6Y3CAwbbrWNr7QJwM08/fbJyr1ewH7dH6KWWQUVtbG
YoaS4NGMkwW3JOv/8Qe1KLdVF0UNMr7+gcXjB9Qen8cISu5uHdazRpKSqEhCq7sHlLmxqb/jqs57
i7nNRuRA/HKm+DoWQc6dBH20fXayC3OqXqkoKVdzMUNP+BH8QkZS8QFqb4LM0L4bZS2zf9RBhjyO
f0S22V/n3Zc8RCDsJ49I/LH/45iJFd1Tu7JP1l6T/GU5RVD273H/Dd7wwKcD7K4ylZzEt2LSEjL6
sqkU1afSFEqmCrsWN+MVJgmQ3nRo/fpdlbr+TmDiBy4PUcttTzTrjltGjTB2Z9tubeTnW6ITjtwx
GfVHxjdkFv2MfaBqcFixxV8QAhVH4wbIg2a4ElJ+tBR+IvPiem3prlj33Dh9IA87M/gY623SQrRT
gNsU/t7FmgOwZ1UtQDYr/ZvM4MVTqjDBL7i8mudEI8p8BgIlSoHu7r7IvVEST5r3eTR0q9zqBNqt
CUXIkXAzcfYRF1wTbXZUwozk/4KXJCiZD3Qz+onhaHVnRHrND4mlwlldnuFCRUtN5prlTBrbjQHu
6eaYSRQlTbct+LkNzoxVqxC3P1GmHPDm8Clwl+VYedkduSUL8ykt0xFwfCS5DGiiub4lODwZS1fb
qkbJrewb6uYV6oQfL+yYFF5ZUqQGpzTIqXhPABbV+4Jdd4FHnT9vjdCOqSRp9BSqjoqmx0Pw4yvj
7zk5lp9F7eFi+ETdb0fMsCjrNNqYtC7ypDXvDEoeL4Z4JjcCMycP5dgWVjh+XEyhSxi6XSjjqNnW
ZWBgpYP8/RdrOPqIg58NKmx6ziKZvQVPuAnEYqY+KEw6iiARe+krv5EokIGRMw9hqJid251wl4FW
35taaAoiUp8XGxbdEAn4e6H52O3YISwbDaBPIcK+WB/tmuwVBNdVtWttC/Pt++ByBEp+T0exCyS3
GjFiQTWMs9OjF72OXkyyWnESQCPDleZIhU5n2fHBuHspRnH4W+Bwk+CtqjSYAlWGq3XvTVQpsL/Z
7ZJ9LD53nMrdXuvBphoO+baTU2gr3iEt0DiShW+JVIaIibvvfRdKcaTzlTppIkzOqUqm0Ao4wtjO
qtfapL7fwHF80v1Z1wGyZ1W3YUfSh4cwm6YJdZqVpgG+qS0vjAaFPnyEzAXxOqbVZ1yC3wxBTxeo
tgJtbcWNTraiJcBoakTSl7fMKxvjAQyNTZZvfNlyXmTBpV/3e8yZCJokUjZIxM/yF/hpaq9CmnY+
Tkc7PYX79GvkPSIi9nU7kpkRvsV54wZK6s9fyfjXn9dLVq0MBnNrMhb4osMBn4qPzwIPIQD9Z54p
eizPrXmCL6CFYh0OgVPRVfbCo/Ndl5jJ0VF3jysfi+Ho6KJ1WHrKAh6ftR0f4Q5YCLkQ9Ap/jIqX
Xs2TWrt1j+NDzsXxG21ByFbcKvMNlHBd7c8CL9z+q4jig+LXjXWzNsSOufFS/mmmsclMPpdLMmWb
tV7Quk+w8LmHZAKxwsbtXMA87bImHlQ8d4SFc5cNdLzrTE5UeqpGcAl1/7ZtKXZWAHNvDLaKZjgo
cz8jwFlHXPy2XNbD9GT7piKI6GQpGuw6jAkqo2qZdNKcRZ4SaCKp049nWriJ/FRfp6inhMcYwS01
O2rOxZDSSfJNs/87G8f6+cMWi1JZYAQMJNwhw6rNxUvfyUNFkC9tBe1rt/NH3U4NMhxj4N1GAcpt
Yr4d7UOHu2LOt8ud7hg2orVz04+7nbXfCWLe+a7Dy+qNpT1errTQA9+hybRZ3Kgqm2l1NgFjFIV9
GPXNTFikqLlquBtN+l0xsxAEzluzl3RoJjG89DmALU+tLYSdzCQK7kb8ECppdq8FRF3vUxH3NILm
mRhqSi5Lehcmq8yFXWbpH7wR3RTrMqyRa/kfw8XSpgFi0RxBBpHV/+8gLgkhRpopIKtbXw2yblkQ
GeTWzhOy/CIIx0WdUXGXzeQjVdqWf1ynwRWA5Iug2ea5eUz6lSfrJ7Sk4Sf4kuh4uw9Q/CdpfiOv
FEd4GELk6E1gROO3v0gcwTSfmAnld4uiNyWrKX6GDO69uGrsxv6IjBxBPAgrb+GIegS6uMElsx1X
09i33uyZoE/FDoM684am6IGtkxYOCBf/9WNPHLPdMPcAPzxG0uCBfubK8OvgIwXD15q0Mm8DbRRI
BND0z5b8ksnzHoYsJyfGcD3TL+H/Up1xe+zQlzgzXrlKsvyyIc6vun/490ktBlEcqx3IF1gAhJui
y3IeIzOqWz7/L4tc8uBRw+7CJVQIYLrJAZ2qJ+ll3lI/6XYBlBDlSQZpsqJi7wMFxiFlzIayF1VH
sHxyoQg2EorpVsVt/PxK7QmkwMMVRilECkPkvXQwvsqn2lwMagX86AJmI2toLA84k71koSOmH294
te048HjMltOaOc2wQFIgB2XA3hAd2wiycAros9VFhqlZN0yxeDyJrXe5lpOEQIPfRMJJfzd35v9/
v21l07QrFTKTqVAdIJ3cRGvu1vNjcO3QpKUBf1wixaYYrmQ8JP6EtlTXTXj/A3uxErIgVyLWDbS4
r5ZghilRs0gbCaxI91XNcYn/6WWC0KD7dcCQzCaOD5ZVwwM0DQyCw+F8T4r0FFUA05asQunc96s1
aP9UWWG89byESs3lT2oEtDil4Jrnguy3X8GCUNi3KwLUwxiSrpsoW/Cc4uGnKpOKVbiIu0wU3jTR
sq6ZBIPqD/59CuLUd8H2ny3qavx1Kj+p/R7jitPXyZLuwsRu1BywVoQ6FvJ5TraOIyN26z6NGWtV
jofDfUcxHvFAp5mVYF9oypP6HxamAnkXNMKMltGS1tO1Y5Krqkqs9xd8BaUAaNL22T6A0ZXXy1xJ
CW4Zr/+oBJejzyE0vgPXOj7IP1ZVsGAztJYZ2sNXqLCm1JOXjToqZCDTclu6SiYeCAVsjIfDOGen
Uz69YcOKAef6Dwa4GhzdaBlsICqQrwF5N6aV++AP3R5XkruXlSaz6bwDKdZBfDo0TjaHidZfjTiL
EeBclatXhSyEuKD5n5Pa0K8EzIHAiFr3yzjh3qYHL8RL025CAAv2bMlwPCyJheb6i1f6GRu5vN/b
AXpSrL5+a/VYzTe9pJk6V9iQuPtwE500RbFpaayz1QIKJO3lzY+0ympeaE9+tOotTQ8D3KaTfzJ3
+KoJoswVM31HegT9GruPHI7ybqu8KIwRJ8l1Z1AD5cU/duZgOpAPZYHEzHwUpFPPidr+TeFs2BUz
0CTFhX7cY5eYTAVIsklFtQkC881OkTGtYTKKgqXhaIwjgtKWygEixeuGrvhMcu6Z8KgRbLNw+9B3
D3bf8vTS/9zuPIssFaHM1SZCfV8MYCmIelZx2wllQG/zSOX1y8amqVw6lJc4wltgEoIUI2kmKjaS
6k96UjF0YkcRnQNibPVw60DW/TXB0A4Jws+FycmIGxZiVpPKTxvEteXKHZ3SIAQNDn9J3Y5iLUhO
tybGVqfJrRczYrh0xpRy/UR1nxnFEGedaOnxBP+PqaGFdpvHaxAyLXJjP5NZkGMyF0sku5+MJLYj
ZvYaFI5t14FO8dANMFo88oGhCFld7vJv0Jdgbkeabf+vI8/A+8FcZnbX2wbMlTZudf/PAjF3vINI
McGqZjc6e8nm1ZYYszMyIHsM+1dNGHsWq1MqqNGiQzjzdvuVykf+wsv/4atFuSV40btOD/SyZ528
ZiyRTpjeaCIWv3tOAR8X7yun095w17Pe60l9nNPjF3VaHuNU8hK4rop50Q4nZx79y5IOnpexfAn+
7JPr80V0+ymBM0uFue8xj0K0WygnsJG6/iu82Sct/JGk2QGCDA5la4ueJ6qBxV84caodPHnfG3QK
lvtrEYMMAXfZu7CBfWQ5VyzPhvjjFKojIObgk2jJ5SB+Jt1rK9NdMdFHXRS28qk5gaKARtMzfExy
vzpZaLKuFt0TbLQNUQ7m20yPqYdyrl5Hacxe9lCN96iRf4mxHAT290VjoR5HTO+HPn7nxybN9nv9
w7gfAJPenVagx+j9pGDERkISAqDhbKcDqUZAaRgWZ101qflKBMKAuTur5jmtdXuTkJTrPibbBDYl
Lg/NvdujI8UnfahOLK7mlOM1t128hUIU43LYhqQnRp4HtsTtPC5J71rDtgbgCOZDXzBOC8po/ZmW
NU/VXITTkX3s261n1+0O18tybylfe+WKEOcAyb4Czrx3HLN0HmDa2IwEAxBHFvI268PTG/61t3wH
Elvz14xRlfNQ/8gz8SBSyWTBjvOlp5DqZurGCQaGwKbal0JRahL4xSkD6h1np/fup4VqD+OhRtjP
28zi6TdApqJ+QaCdG4K0sLW1HYfKaATh3pcr0Dc84KR+AoBxsSA+rNyw8mQk21cP4J1XiKpSrsw1
Ynv+h+KSnH3aT4GdQCxXdICxS5PDGaAFbDqrB+ULVepMWd8XcOhAO+bmOirKKwkbe7mIIKB4rzXp
Svu2Q4mJB7NHtnYGRSKSTv28t5wga8u2Rum7FrspGXVhYQzlsvyx/dgn2uOwtsSf3QbXlwJMdDZ6
QOeKTjg00IWo3Rtnwnut1l2R4VQHNKhShgke/8uoycKwvB4RQtUD8Rh73lr0tVG4lxkit1VWCOg6
/FseSXYKUK4f0w0z/u6fkOE/yzr00QY4DQjh4PuSPuDdLJLWLP/A5uplETb4aEKo575sx3sISpKe
3eyqDVU+26haMKxrjyp0YVxqB7THh18y6EqTyu/edElKcIS3JCt/0RtH0qKt/d3VR/RvCM9A0gWI
TVEhc3c5xlKGWamHl3ppbVXGCMV3XDkmRimemCAHRB8MzZdfhyXlyoPV5b9sq0gOpGrFzh85ubTg
muCI/hq2D2u9HHX3dnb24hmFmGXRcULDUH2ZnlStyLUJGDEYFzHovf/Tmz4Ov04m5zTaAF7e4Bwf
j5k3rMLTmvk6IAY0xmh1UCBgJD1OLFFZEoEEp/LBGcTxP1YAuchh2MQX4mCqvBUw+NnH
`protect end_protected

