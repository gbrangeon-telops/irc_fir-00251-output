

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
nqqBtmqfflVo0LfdOWD2OeylbTCJPLX6XaSqFQpCXkHX4TF1QAXZspyiDVaQlwRkat06cPZ5E411
bTzbr9/qZQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Q/X3qbnpTyRXgHhmurX8chlDRL2XjwnbHjo5m2aoqrTNSVAUPYEYGIGJVoJhRP1Bd27KZbGI0BFX
fZKfju5H4nz84jXPUC/rcsp76WTu945qoXwdo30XI0Qhi1w21P6EhLXccz1l4c9zfTwlHtVuYV2c
xkxHRh0F8KrrR61HDHc=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
jBFh6UBl2pQmyl/KNdwY4r9ld/Frb+RgwTVitzK9Y6Fp+6xDwrsib4d9Z9Trd2PuW5z5/ot40n86
vR7VZpJnONM8UmDjWgdiB8rXNXaI1rBfme4TQ3jj6RaF803c2cAi4cdZ4qM3X7V29W2B5HXbYsfA
+fn+v+caVjEUXZHZm4HMyIR7TNVnvmCWeeLj52d+u3MrD7UjjkqtqnRWdy0ckM9p4TE27eiu/nsz
awiAJoiVLZNTMmdaTdZ6vB/sS67SAe0JjX1nTwssfK86UYU1+n0NLZ+SLB4lkqxmhepGPNojfE8p
9hJaPKOTV3d/umJbTV97L90iPloNPMXpGK/m+A==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
cwUUX8orCEMoCaO4wbzIkA5h1G/QOLlup3/J46IxMYEEhFnVuE82RZ46tcCa958uxg+L9/l1SnQ1
1Qa6GFDzaEz3zEcSDS+t0jFMPNI7VUppaIgcalGdkOXBIX9fihrhASeWjqmTDrUSlTt7Vzyo+3TY
n3HFHRbTrCchXcVswqs=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Z1XHzIMnint6AvJuhSJyN/+kraiZwIT5ZFNyZxcRS4ee586ZcCrsBlqjvo3awgeNWb2yZNQKbtJY
UBJT2Ww9PtMdwpg4MPuZFMCTECdiBOLjqX7gX0K3iBdA+35RXRVkpnaon7ABi2dY8SU6a03iv3ph
ed9P79UVGmdGucbzSQNo8vkiW9pS6ZJElXKmEibSc0C9Vw6VmCNdLosnrss+vUEVkPDu65r8MqDO
9/2zcjIio0kfnpSLOaIDXqGefGNR89nRv/NxKymzLnDjvK13FSfKq6qNfA+cXOtnv8oRuf0tdkh7
e8F12j/LQajA5bXDfmPQ3bNX4Qv06vuQ9+MAAw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 89616)
`protect data_block
gLP4cAsKthx5uLMMy950XiX/WLDbKygZeVPjONk8I+vi0MD1dGQnA8DlpjEca32z9LLfs/2+APog
4Upn2KN/V15qaXQH9p8HhHhQ2oa4XGd1PNyQcd3ufFe7cYKvbY0WXrK25+EXPeUQv/GRZO72w8UC
tSjAyUv5KiDrPLgk0/H2vgprc4D9RFaSql1P59OAbbcCPzwfdIUg4UYmEYloRKXeLUKF6WWQ5tnK
yzeKVtnItICVeaa9N5ZZfLpfgMk4swPnifIIw6H+vPZGz39LC9DHkeSta9ICgEGjq8igzyG612hQ
6J7ZTT1pOz8d3QbUxwJOduzDiN1h/fpP5zL4kKcZCe0Ks2I9oY+iLh7aJp5GFyiW82s4jLont7jd
+ibtnHI9G01DH8y821hCfuYvyVl5DalYz5zB/dQtrsen9Ra/sx6QxuLs2AhITlF14vLI8zQ7MkMh
bf6IZAKb7NnZp9KxA+HPoM5Bl5o2GYiT72Bg7eiqFDfUDXxgMVkvRcArSz4MKgoCPBJUtdokibwi
wpdFSH2O0myf/oq0lWmn4j7CiYs2hQN2b/G+xTPFDx0F7b6C6akgzJtrH94F5F+n3JgOW2aDIvJa
Cr26oWpUK2tAVgH38xZOwm3xHHnhRAdpFad/vHohQ80383fHBXcFPAu3Mdxh8yZxLBULVC4IBStM
YrKJANCM6XBjz+jPgRrIlM7ErTRifIpJZWhY45U6h8gTz3bb53tHpmUBXD5LVU5zSAAfBroD04vS
/jHxnmY7ADny0PkEbZmj+voSqzSWKqFDY5WKuvCP+vllzY0vd5x6P6X0UUDXeklUehiOuCH+ibfp
Tp+mIZ3F/bdDCUUhATDxzX7hF3+08HaBczPBIgxAO5wPDBrIkROyVK4nQkmdUTwjgpsBJ99bIUMS
vXV8+H6Icxm2UZPhbHNd1NtWpTRCnbQ2lsbDiAVDpBMubGiYbAAsRe+/w1elZTlTSrbWeOsReF1c
YuIg5zrzhAgOIj0wBoPRBtg7ihRDprTKpOoAjswEtRuVzVcBGjX8/gnG20pyfX6Q2eJR9j9BaZod
+i1twu5rFDAPCrOUnCMeFlzhkrW6vleAFYCGT8ZOZIlCC26IfCnoOW6EgYywBNJaaRPYJ9oacu7k
taI82EouRWFlxJchGaOjUfSGQfmklsG9iYey92inOlQZnZltxulc0Q7oKsl/5Ric0L2aDPWWs669
iZr75CtYzvmVoTwKOq1vNFwwfya8ImBYDfh281JhytYNHM/alFCvRg5sdCL5af4VPoTRLeyhgZVN
53RBk96qt7GHNC7zfHVFVwIcargZD8pbKkNAgKBRDRMPqaAZ767KGP1icojm1XzHcUiTX816UrVd
VrdwbozgMmesOY4adoxlvrXF4zecEcPI77a2baBKXg9BhBHYIwwvFejUgPXvC+WoSoF67Fsse7cH
JARKOhZ3Inm+BwHx4aP5S0yR8ShG2LhEjhBZD404m5aavVRvqlOgeIYQcsyQetSiGHZ6MFZgSa4j
Dhi0atyYDSix+Ht5Mxfo5rQOD/QQvDjvj46/WBknM+mHOHgFod/DGNEzY1vxTaGeyg2sMX+5HoRK
7vVLsXBSD8OJ22Etro4KIsbXX4NARQWYzx/DnfwKRUxP48hb3oRh1EP1e0TUPbdSo++9I0UOcBxC
jMsGJwkYF615IWN+PcJz6QNLFW3GR7vOd/xLZKpOyTB3QBEG26u6QpU32UXIz9qeBD936hw1vT6d
rl3AfMR9iJg11kqWVPlRGRRcEpTZGg/wyrJr/t6GnbGgvGavFuJjySTq2im3Gn7aH4BNTpRMm/6u
I6JIdnGyeZ6niTDO2RXXze0Yx3MFrii0wnQCFGxT3iLWorFpfDYMs9zRpPvxVYrDHAUME+rKdNze
VZ3aEnrp9bHDoExlwyf2LYK7w+TDF/5nSEM+/45KXsKySD+Vt+gg0kYp0LWdfnuQqJz9Z/DsFnSW
XKUoSpL23NDyLfl//C/TgBGs6O+kEfsNEt3zMiIQ5MQUv8evOG2R0Rs2C0I2aUbKdgYAlAiQM3yh
+XOj8rz5jGjav9hQ5hRGTwXOCL5vb1tqMlCoHguu1daiWTwab/RQbT37nCw5mYqaT+RSUELwTiUT
C9TvtE4CK2MkcCEgNKuL5cjtcfqpx/VLT2WPBcoD6f8bliFHMZUoXJJ4tTSQFfl8hGV0YQmWL8uV
+ilyfLoLLu7OnYtmuXYERmY1jl+bfRN8IT7WfCJCnLUljyc2RNy33ZZcGrGfk9EBEmqxpt+sUgit
zHUOb9RHvI1XxikElrRD0OZwSbL23AFZhT5uDFmsi6BSlDd9jbqwJLX/H07h6qHXfW9Wdc8ZBpvC
67HMyOmYzJa3SpMQnhxgdxEu0x+idMX5U7kyvhU1nGxrwRofT+AhmL2AAPJ8h5JTOdh0iqJYZDSb
UksUHmzU8ALMHckD72CCUFocqYcqg+UmJ8VyMWrbKWhaOcCVUsKoaywN4cAizE1VIe3bk/1xaNh2
rKQZGOde6bwBxiCVr6FFaLZRpa9N4jflPkFHPS7Y8OP+qY5d6Tqf55gcqI1GWB8T0cd+rG5rUoBn
hiycfBTJrFNAaVc/DhsAsb4g4m0ynCqlHImGwpzx9WmJO9wbuQG5iL/H/LqgJghn0MeRK4PVsyiW
n3nCI8dQBHwJtkuYdd+S36xBfdRqBH6wd6QBrZQkneuNts70dQ1iY0E80+GQ7FWvE4qrNLi383r6
avsp1XW+b3B1x74rQKGbOiOFS4yqleoF3BekJ/WKUp91wwactIPW8DTsQe6/YKpXcpnU9TYeOF/H
kHZPHSdWIE2+MhFCB2TP0q3PiM//mgCEsVELsJ6O26S9L6JL1Wwhdav1M0mnu/dCFZZNjE9ataHz
gDx15+NoCJCYsIHGQ8ZDW2wgUDW7XEalaAKM9tvFrCqWKqrgH+oZic4gd0k0Te0ITO+WA1Bb6BwL
crkyCAdQAGNqLSPeDXj04z0yXzgy4ymOc3t0fAcXlsLyVor7D2B2wJNXSHLR7qnLfibvG+S7osWy
6L3uVqYPw/XCEhJ7C7s7ZwVgQ3ggxZf2dbUl/hFF+VnFY79Dfrspytfuy5Mjq4HoZOXppPGJ3Sqy
6Kp0Ku3zfMThyMLfcmh36z+LRwuW9z7IJeUBlAnlIEn8Cscgiu5hFHqi4Uu/OQ1GmoCz+uBdG3JG
DpkM/9M6GhEJQpVeP3KEoVdbnRSh1h8yY9KvmRHPGbFa0RP3fVdVOvDalMYr2abldurns8Zq8J6v
5zSuHT9F9VjwRsxrYH4NxNeI3/Io6+xUyeLkl3n3ycKW6WyYu3Wt7G42BW2cBaZA7vItbtBXosH4
i9Fd4e5bWwz0gX1iuzLyXldMXXqgC6r8SznF/Cnrg6BihhwwzYLzeI1Xx/B4iSp01LyxLzWzuBaa
I2kNbBQqTH0nxKpkS+5ofDG0dEQ6q9MhkeUjDCK7in1MyUBYBqanM71uy0PZho2Gp1maWOlQj9go
0YYp6Cb4yc8xHc5uVFN83l/Ph2o/5GMYOmvxh9jl9Ajz0+B9eW4Chsd0H79Net/AR7Y8aamCPhHr
ODUJNGnXBfFYOfWjgUqp174E0yFliAqe/KetM5Pu7tcgGRy9Y+bQKmXsLNHAJH57LnqLrta37DW0
NXRsODc63rKz7k0L3Hzr00twbe3EIoHMpHucDSPt/oY/QBFvtEF4uaouIgYxeJljIf37QBTsdnGA
vVl/fMi6U7I1XA1lWhf0kKJPQlmdFneBanM4hTSrbJbpgf3TMP1nJLhNlcviwgqxBXNdVtGyhvu6
SarGwrzQCOelUiAeQ5ZihAkJ/MfzYAAsyBDt3oNIFzsYG32GlwEcfI9PlmqvuvdpR+V/Hmtmy2zV
17yV+XQ9CDPJZPTU4Vm8xbdKFiK8sI/pP69haiCxIk+e9UZAxiRe6PzgJHKGjrCo0j+gr69HRjTV
+syudxMEdMzP4XxWSdEYsVtCUgfBcmfKY/hP9spuqwKvTzzIRfrBvSIYki8z4HfSkDLClqQvSY+z
KX8g4/FGjkM/KeZUkYgnIvovTW/KbRhHEg75GzoOwNTeKNGeCRp9fUmWAuyZoWL+iinSDxlU86cX
nfC6oCsRUzT24WAGMu/YHBzCqP0cXBjSo/ZpvEJZvdv2wqN7Uc0AeV0sX1w6mZfcea3y15RxCmpT
M9R4jQpg0HeauUiYqvstRry/CcmERO423olCErvzLzT8mrrf+mHq8MoZHi9jtU5QWwx+Jtxu/bIF
7Tli7wS/rloT3o1aB5DBQw0ngo5Xa4K16tc7vUmWRxKlVvQuyqKeYtCrj4r7GA3JNzt1epxM2JSZ
ag6zzZespzFBGH+50vbM0prZFtfpheJrDHhbEUbNlEvekL1chKF05rwrAbgxcLl4AM4lZp75bV9m
p3/LLY5096XQfs4HDeH7Og9AKu19/2+fcHAndVArKKgW5qgocTjmx8Y2p1KMVN+KUuWkgnNWH+tI
EnXRglfCYFF5XQHd7D6fYFfy7CLOvb62hA63z8mT/nINlDg3bLzc69cZJaObZDiBjx5olwrCxToG
+2+sXxwOMaQL2VuVDa7J7j0OqJKyrXwQG9K6q868+gZ3TuQk1KKbQpmEDY3Mih57DKoaPp6fthZc
85o0oqPt6uv6C1TKjXOSi0/7AsbYob/GpkXgFe1qOXSZFfRSvOG6XQ4ooj2qgDq/R53REpR2WUgp
3il82ptWmcyeMyh1Li8+Pi5/CqWqz6317DYOl7VSOP8TKtnWQGS389PoqsgHpnESi/e1ZXFWNOfZ
Dv7h2NMBDsIOr/hWFiZZhQiieiulG9ERHUC8nCxt9vmrDOzQ9KhIZ7PSChwnCjkGJ6DSqZpbW204
hwdMpTBLpdBypONqLwxZVDfUYlX+8eFGRpAdm+ACsr734tV+F1qjcb3gclIlYuILaDMHPr9cl173
vwey8UjHXL//2lp+TWBU22DX7kTfIejVR8TCC3kgQYVvVH+pomDIxQXk7uQGvYXJsFk+jg22WeUj
SlBSLcnc42NUAM29Tcd+dzj7nMC1/NVHk3vdrSxfg++SHQWiwZLpMqLPyxCWbwQH4uNlPTeQF6kP
PjE57JKvvn4MZfUfFnKtuXmL7x6U5adSGcsEs8xDYT2AcuXsJ9/zDI6KXglwD2fGq7IR4joQjCHW
v/t1TnPeZDqrei2Fo8FeizivGHbHEwA/GuTLxFSQMyn7S4gu62xcNRCZS93DjUQZ3GFV2GQlucMO
T9zLJ5PkaoOwzp4n+3xJ49E/dtFJpKjeWVMMG571UmzM9AS/dCRZhW5ONIS5IbIPuYzZRItDG6lz
nVAlIP21kPndSOovrsi+NHpgW+4oyXSJbcv9ZIS57cWm3WBlkKqUvVK9W63R93VpQ54bvSVsbqub
Skcp3xhTaXk1rP7RcCXntnnVlDZefiZw2hXyNTnn+pRHGK6hHm173aHNDrS0kglyYzis14qC2Z8F
Jlfqt88aI2eJdNAExlX4TjtzAVcChDPeakw73BlTw3QIcnfzKPmYe5dUJPsgEq0XSp9q6VHOfmto
FbItBS29SUqeXAphcrgwRaANLsxBtNSnfFjhPjqDJwDfgOyMbgmDEiPHLpQBmLa2CHYju9j4zDSb
WaEwkuoEOmVOOQ7p1utQ6++EzhsXP9d/nzJQBSvGJkTR5ZD5VYDaBnqJ3j7kUYQ4e8JSm2FMgw5S
W+uolsswxNMubawtQJFNybi73HGlbADmDVlZHgmt/D4HS6jfxZbUcecSImedJXDm3U4YYzhLlQZT
JKYc3PlpJ3wBrGQEuybEHdy7eOdEwcQ2OjugSPOgYNzR2HOAbbGK6oL5veVUasVmj2iqgYON3Bdp
z2ZtlgAEKnNaTe639DrOrv8mdoNy0dHJgS4HkDO6jLocHeZzP79ZV0Rs0oZN6zOg0BlbpU3rw1/g
3/yWW5fo8G+IKqXpXe6/kj+tU76mTM52F87ewfyAWid7ADYnLax9w2KFouROKcW1WaUMOknhxlMF
5eaoR0zCdS2zg8romoObd41m5j7Va3rtRCiSc3Zr8aRhtSk2S7kdmMraF4AIORPFOZSzt+ZAEbdQ
0bAOy6ae3/5FRiXX2rI7oEdRvCSXxKoNrqJgSPuh2aZgmVX0wjtme5kjvYcrgZYEbKWBGdE96Cj6
TjZHHmU4t5aO4cDwaVJ7+QbwOyVvvxFD45MKoGFCsNBzZKwtdb07inXZOa0972dYXaZWieI6BpuE
Xa/N40of80Sp+3We6FLlf9363g6BknzY7tD8vzP3NjBTN4ZN6fYAM1f1WkMXYKdHf402JJPJ+hc0
C0uE6ZsZ0/8pQXx9i3k9Ln6ln9RYlEquNUr8NZSDlAy7x0nwMfH7gYWYx42nsXETsQufx5b4DyIR
9g1T31HtxFHT8IekUmIGSaLJJjiDjMjIL/jIKJhmyzytCxpFLmP7S3PZ1x0g1rwyTpA9x5+vNvZl
40ebd1ElAZ2GjkhNk3UeAjcMtmCGuUxaNlU13wQ3CQIrgammTRxmpveZd6YfFo+Vi7aw1L2WIixf
EohAZ2LK5yFwprZRIrBGcvHKMN6/Gee7QMAuy76kU4VXaSINYSj5WwkEEoeRv0md5fgLb6Nenvly
3DSb5ddYe/mnr8Z8g46YSSE0ikeqIkw8Bcj9QwLxF1IWLchLQ3c5WnlkheN8Nkn72RE8S5vSxQFf
p8z92xLnkrVkpRuUZE3XLfe8avsO2buX12bXVKKVF8yJS8OMpMY4yKctxnhd3ZHW5e1qlR5woTnd
w7Q3s6SAeP9S8slABro6RT9fsN5Gn49WPWTjii4WvfKSg3tRwzPkV7SAeoEqwMhU3dd9pJHmt0en
6VqNAix/trYRX1ikgzet5ktPgtf7xZaTjjZYDTy4f/k4FtMCi9nm0IyevEvvN77TZ70VnhdbOsHh
T4kG+5OvJFYxsN7xkuczWVrWdj1ew3ttvNbgI9RviJ+rWjEJe8Ywos2AMGDHuDyAy1cFOTUvAv8d
JzLGZayrbfHqL0KS8Y4AC/5/wmj8Yo0H8K1woFvJsyU+mdzJm2PnPyx0Q3VFK4WKP5yTXN5sPl8J
xdHOKcA3hpV7CuPJQl3B9nyJ/eTOyGyE2tk32nlLiesui++YjEYRwiRVlgpJtkoFIF31DlNOcivl
3znrwUdA8YIA2gCDE01TZOZR2ThGKtIwUP/A0HsUp8uycW4GvMy2Fl8JR3pKAKseEG2eOWBdWiUs
ZEpMFbODdoWGC5w9X4bKPOQARpler5e6u/Qv+6JR3UKbSgxF1I2UbT9EIkPSD7yt6pbWydnIVcqq
gTFrk1fyQQmBenxnGzEzZ2+nMSVIJaL68FKA8dKvbjg0O6YWqoBhafG1dpLD6KHrULWpsbfYlE+e
13pG7P9qTBNl8dbVoITqAs+NL7HcTqXlfWb3gOqQbvtEb//SfE9KBqVLoTbf9ax6sHnM/bOKg8Bg
8McVm7VFwwRYerAeUlD8CXDn3e0Fwao/XMzks6bKdMsR9iKS+d2aeN1R1DRx868FXT4ht234ZHqT
K1SvTy3DgM7eRIH5ZX5j9hzmRNVWxtj1WopxGtS+QdVTfIQNIHx8GZlg+1hX8tzaGTXOVa4C0KIu
aSNul5xBxK5E3a+gvtCaqKhNE+uiwuNQ1+rTKz7Q2UTzx2P/VxQEW5D8aALLnerq34ACWPl3YA+Q
1PS8GW0avY363Efbajjcu3lLnN4OD4Xdw1DCrvuKOMH+NJOAfxGBNt05S4BFsEmcIGBxdAEAG0kY
BUyxs+YGZt2MQkEgQNnBZNcVVGs30hQn1YbWpssONFmm+gFOuPSlAt7/0Aojvwz/QSqMslcKuVBU
+TVE3HXWCh1YQbdwkDrl8LYpB/BIgn8JU1Y1l2QZKqlA/2xwB+BAJsKAcFzzHg1xTUZo5f8gqWLO
Mf6X9of1PPuTEH6TCTokrymTI7epOP7iY2UgUihm7oHvVMqZL9ziEeIbgZWV4Kgw/WdLVauOwnnd
HWfT10FunatiIdWvmXVSFPTW9UjvmLkofvvM15r706zYWp6Usk4FFm2Mji5PCF4PPNvro0Sn858e
sOwGAOOD9Ons/ja/uoI0ykQTsXahOjWsJUG/DChrv+c7PsSff8YkDw49D98m0PGD0sBEUwMQSZny
cAi6/Zh3pSMGPdv5jAkuUZ7BLofvW4YD3CbBwKm0t5Q0lWFLYu7kI1qlJSWIrdvZfsVx8MGwUFMV
4SMwkPCwiPWy01wrS4dpwMeVV2PVGJrlj3SD4neKe8tweRST3OgHrOxLx1fvKoRlY/+qdt1IwMKh
nnCDn9IchxHXFwUPhW9GoNhI73L0dTYSxg/vAOK49qVqvt66i9cCjHx78HPqkKFb7jy3V7seVtnu
/pQMFueqqL9ADVUAbY+njFyLZesoxoZ6ATYdfeet4h13wztPGq6cSHbUDgbXvvnLep7KlnqYVlMQ
0RNFYEh2V5CzXV4h0zYNQdlEGanf7XY5w3hBqSr/w7wvchUX0q0qZPte3SKwqC3XkDrwRiEZF0HI
GG2BAlq+tANb2Uj7YlRx/PPcIsp24eIEY/UhlqWCwqqISyvH5rmZzpKmQdBKqZrNrCzdANfyig8w
r84qCU9JqjQx52Pqrut3ELFM7kKYlutm0Pc/FFvo2VQFO8iAsoNJcWL7p/nKnw1Pc3YhcOONlFhp
lJcmWNoTMMmsk8rOvAst4PCfomAuXvD40BtWShVQLQpsm7MZgQvEEGxyaVWT6RcbZgKggiyGB+VW
CdXoAtCbPd6Ffm3rnDUe1gB4bO+q9LI9yZ6TkB9aHLyeXBNwf/O0FdsKvlUfV++tglUjomkF0ehA
HlGPWGGRLuDTh2t/KqB2wZ64Ge2GmUpLBF7KimfprHkPPsuAgc3ks9PlfUZm7+f2VuOPCB4No2X6
GPmUNuHvBrzv6SRNRytuZ5CzKTlb1YfNlbFfqLyn9RDvExMhgjSC/AhSYdLDyscr6TYVnyAs8pat
ZJ8jTG/TRBwWjcE8KJV95ifnwmbsit7DjrFhCHQEb9+av8fa5RhGiHM3Drq6xNyFDQ/rpCWUTSWM
uw5uPLGz7hoiLNYLf5YHGXHPSFpwyatPzghBP5WToqTSeUz2QKOkVOMtedqoTu+Z9TemvyKM2/pp
bT1Vw+4KIHSAq+3MngGyEqDMDFAZSYFtiZNcOKIQkjVkrLg9MIe7KKTHDorVfMmXEESf+izOqMFl
+sKnUbTYjoOshTkMH0A+lVeKK7hZK3/FMOzvoFqllLtueSktFm+x47Y5MqP0p1dvU+qjw9ClCMm2
4gfP7F1Led5IYN60MUOl6ZO351xWZP+sRp+w5Tz9ebxFEX+Qt+eujQbYwSrlme++YSHqWh9vBdiO
+37j9Mwg9sF4vF7d1xqcNNGHAQV0GK/9+oJzlsQAM3lsAoMy7WpiEYhOf7WtWmRJP5xIqS5P7LY1
XJKq8NPFx674HLI+I6teegHlF/OQVnWEl6LEzTgDh/Wh4VaLumRSbq/iF8owiDZ+y6b+YN0GOsb8
GRuIkjouZsTnc3HEjjJmTy3aaTZ5UcPGkoIgmCi67wvHVzeBi7ZwAGqyiiMhR1tpzmOIuEqnFpYL
dS8vU89TaR3llmLAq/wF8V6Ll6Y0huNM6jSsyRjtBss9mvjpKEDGBCW9/f1w7gdNNLApjj5WzpG8
ymxgOiNJELTlZpy4/LTdstR9OH9DUsk4W2FRMBSo0wCuLz2MuuZh/JPr9XEHNloGpmKpvzQxDShA
W5Ktg/DGtbPDcjg0L0NuDe0mAuqHWbJlHeL96hKPw/xkVYaG9ViNAlXHhe0Zs1eC7VKhe2SwOUUh
t8bR8JGhLHujP+xSxwu1yRyvay00b441GtXIPoVWJCx8gdBXfoTHdALxbJyJiI+esEK6vUUB4SzR
BahwL/ZB2j7gZDHPqPuxvisAtbAQMuVPbHW87Bbz5F9yxabCiL3gdCZyjeguwHCeozpkeWoFRLzH
8AmAl50M98IkCTeR1dYZY7+z5EDRywu8gR3cupbNwjPBfnj/pCKYayT25HIOfsuwU/XHFPhT+d7X
5VSgsQtPdrTswCCH+CQHgJQWOuo6hslibWoBob7JUgOX2iQ6fpP5f2z739BXGrcS1znDJ4TTT5ry
VNkhdYmDxWAcjWkQAIMyEe+7DmlBlXwZgoPhVDLsMOXBKfPUQwgc3urcir5M6OqHHkqVdBh78K4d
EPZGXYkaY2xNEDb/yILFmcuWdU8IznlT4fVLybsx7pftOgpx8a3t+08fmAwcPvfe09qLgTA9hniG
ooZ9wwR9XIRCE8uB+usg44Om0WKKPzFX6RJPOjc/kXEwcqY6tRJMrHMhGeYdzgg2XqsivNDw8UfQ
o/Cu6r8hoj44a4J7WIWQpdMsGFWBIDirubMWGH1csURHsbQh5MwsyQjUNzgZGJDTH2NE04ADE3gJ
DkDSuhfxf21qN9ZbIcVtTQfvOIN9T1Zi3SJwPqoxDthWbBaFvsEIfTiJYLt2wIrr55by/mow+DfI
gcOWoxciRcZScH3h/xoTdDnO5QMD+OCEakrEu2GqEs4Poy0O/4NBmCmUd2Wr4Juayf/JALXyhXSO
mWfBotTBNUvQPZNi6+TMSmgfiHMY+dsRpRRFBGO4DYVOqiZ0Pk+s8kpHFK4QiJPpYHf794/UIslo
tlumSaifSH4U2wdMD8QXMD7GFQo4AkNbgaPao6JXVS/3FxvPGEdIJDlnwTQIKWsCMCmSrpNMN4YU
vCvf1NW2nF6gYzZNZg322iiclLqkHxNyJZ5glFi27IgGzUV9O1588f+coExcs3KQdYuZqhOoZu28
/Me7TTZNbAHXH51B49xDU45IHgT8R/4Y4wS9VFigeYVBoWSL4IKOwlX4mfJGjNfIya+9Tkfg99bK
MP1mBUx8tp2+fQc7M+pfb22uEkIWWAnPBx3Xgr1dC9KYTtXvRPTERwcTjDSPqerOL8oFAyxQLyEG
J8Limeha+IxDPQosnUfUvg9jtDZAwhKoc+Jr8HfHVibvDCYERf3FM+YMW/fupvPThv5TyhQgoegW
Itxh45pLekVvFr5BvHFYOIrw/q/08J69ngfH2x1NKOfsmYFNAUOqDhTlUjGHKbgOp/Od/msKrMGw
9Rt6CYwalYwwO6h9iNqA3qfhPk7X8SL0Rl8kWYr1holRcH/IOkD9tFAptcGil1Ic8TyuBEbRODaq
Xd2UNg7Lhl7jdd1haW9ZyMzWVuyjAW2A8IyRW8T9zc8Sqb2uVfym4T+nqjngYWmIvO/Skowuj6Ka
AAmnNyDVYYHqSWe98KaeNdul2Wb/tlnjiE5+xHij8F5AEBZzfjerhxBOT3oMORIDfPH7PtB2vnQG
MOQfbUR8NZmmJq0Bm88LUCTN2B0TwPY+TYkCLHx4A0UCpPRGuFb7I5T4qE1AYDbbq2BHvAXJAumg
yz8tpS51vSw2kDiGQOCnI7yU8ZV3Y3Cjp1lFdEaQAjodW/Ty8KSReGY3Dzu0d4+MkRznUH6WwRN/
u/bv4CKSpgWCYWL90h9RcCUOxzI8ReyyG0FuGo6F881Rs0Th16azIM+xobCO5F74Fnycn19ZTUmL
63Y1G48oYrdEX+nQHxNd5FXRhNbXtvv9jB7e4xKJ4Dafr9g80F0x3BC31UQjTdgvHarNo9wgock8
kIf9CbN1nhU+5hchmcWBVZ/bVtcq9wi7frBNULYqlGCA2JkaHealKqB2xX/hZXsrkhpQcpYGyRN8
YvD+LavVW46uCIr8IqZx8UNGNPCGu3ZGr0ERq3yBOXasSPG/HUI65nAnnuup3QdQx2P+PvMdfZX6
Jr+9G+zLtULNvI5C6b8yA8+PDtaOKA2+283NucS/v1K7tK0yWTeJzlk3K7mtVU0nUGiBh1Y6ez+5
daru8DlNutgR7GeyjU++9bKPmVhaxpS7HuwR6Cy2p++Ns6yRZ60m6c8ODu/iknuk1kglp/iW1SLV
oqrWBslquol9d9QVHZk/IVEt5fkDibHpFHtUaDUCc6SPQQ9/s6hjBoe6gvUGVcsO0wFECJ4Ppjxn
sjzcPzt5HWXUra/DQ+F6EvL2oLZEazwKvjHUn2xJG0eOrJRB40RQs5DhpWnbD1AatwhTj3FPWiWg
MMi7pDJCAH7etHBpo+lI1Uj0KL0eb6lmZQgbb9OF1JJ5rwyFXA2pP+VAnOnGj6AG0iNcZ8SSi9Za
NVEFV3e2md6t1xt1kcbw4ohpef9gmj788bSVEea6n6uzmKEOTeD4+J9j6hBk2ImwaLOh3mP1Q2yB
jRN8ptFMhlyhv4Cc0I6C8Ybbx6cIOFgk3LRNzI5SzGfZ/D/IY+6bVNlJkzhT+zgl+R6G8pw9W6zc
TLEH/Z7lHZZgG8mAvQmiTfCgVxfhqmq2TryIfWQALda8bQeXbuaXBIp+JkqGcpe4ZoljHBmSSuec
bGio8M9PTsceKUWxBYKtJBcsnJWPpGgY75kUNxGBrR6/ztyRg1Y6mF4qYMLOz/TMix9p+MFVBUG0
JWp/EL2v94SyIcYXB/81h2z+RtLEb18BZlHmE/JpzVzo778oRMHHy1z3gwSK6RLea+31tfZK8aPB
PuJmgvdWKSdjKe82okxyllH/lu4wqxZz5XWn4wqU++qdb659yhkKla9GrDitcKHPfEk6D5gh34UV
x/cNxIU5957koWKLoDxf4bNsLZX8P8weRHc2vZHU70k2H034HSx4BYjccMaGU1m+6UeYMiChEFZ9
CUHM8dZwL4B/F4Uvm+d6UatlBQUmaCsut6qaEZr/MwbhKwGYoR2AT35th4dXKtLQngI24V+XUl+r
UhnYa8Ry8zCSrbLHONMEjmkdZhEuaz1cORoRWVFpuV/oig68vpv1ui6rO2/z3LaGljC3qO8iyyVF
vFOGLiKqjyvs5oFPSa/XfV9rF0XjH7BflgenbleeAycFZcy3huVqFg8rYpUsaffjK7pD8PlFMVRM
GQ/ohsgXqiHrbx90Ern/5uUOWJyaKL05Gt9877c1Qqexl3LAyPaBj0PvGOPf9K9e+luD1GkhwDUu
xmSjG6yEa3GMhXQnNNekXxEmyR6+xGCVaM5dCQpc0I/cnve0AwDZGH9biFC+jS6icwVUzc/YBR2K
/vsYPER92HeMSP5miWM+LeJ9nt5oFXDkGtalJgUYyj03smWCGpfq214+PnagYJwl8/hD1L4vIaYA
wrzHv10z+vZAeIdd36qlhqcFXK0w6BzDzlz3BoDoFaLDBeN/1uUoNX1XZZWKumBPdlLdAMbCbNE/
gnM+u9jQbd/B8jiBdEfofUlNvBtrWv+RV0efRZNzhDTOlgtksThia6HyB+OQ64B9Nt9YDc8WNvI7
SYV/xfTFotr0RUd3gtjmo0U73Jbn9eoQNpleJRxbgCW9B2fRNI+RIKlXAdy1eMgB8U3Rw7A5/Y4w
hmrfk5HxfVXW6ZmkDBpOh/oIfGiMX2+dsajazXhWEbOC7yrxlRAgZyxg21HYmjIPh8Nt61lhao43
0eUmE/bvh4c5xtu4f1dHMmCQgnZYCQIFxC1OMv1FDZCIHxX/FOhziE218aiMgBOfaCP7rxx8MFvE
S7H46bJeV7F25AmW/IiAoF5U+/dBWS4MW+XSBn7rYmrs+JQr0LiNZgJYiEbrKC/fVUchlZHLDQK6
wXV2jFXqSZpUNHhwmUnVS1iOmlaGQ34tr5V53KVIkoro7ZRPjfvvrONq5STZS3SsJka7NyVxujxU
p1NTb5HCinTF0lnUG6PxZwXInYq2eM+nuCPrn+QhEEG6VX3DvXckuzAexCaFXWQ0mhjoGXilOZa3
51PDKQN6seJqBcgEzPByuo+71A0R8QpSnOa6MQtyVHnH80cDvhMMvKm7hiuMu7OD5eMxKCt9UA0W
HwpCiCf1KhzTW6iie0tLAQoE1YHjyVjSDSycv5kLZJ8/awXX7o1ZKePGO6rOES3b8XGeByPtnqW8
gRGSZAgCUdgx/NhMYYymgN7Z3tO35a5bKCn0I6UYk2H1wmVn6NQoFJKZoyIA7KF0auBE/5e9CSOl
gKsFbbXy05DirgV8f7dH/ZK+3A8aPwYzTMJk3Ikch4rJn+cmazGmH6YzLpcMKm0Tp9yJnNCSBEdE
mk5GcXPOW0o/W+DIf2qBhqfTnE7geMczhFV5RJdQ8doXR/jWnESISz/p5JAPVPsF894G9vxWQNe2
jogHGDGftpA7zH2ma5/ps2wrCqi8OMHyd6vMaykKf1ln/ImgqDgqLM8y6bpCOCDRQjqbUEhPKsce
AyrnBJSTe1h77Ct6PZ8bEOcKNt5TM719nNZuyTooh1ADQOynflQoCnASoIKKc9tvLeliIo/GOxOq
E5XJ5mnIxW609wAEcMxTdKa1YRvw4gkVWG5wRJq+TyNmXcVnIU13bVCBJpmEudQgjR9L1xCrMiGS
jTWFmppt97UrA3q7BNSNODYbHbrpg3AKzBNeXK4tg0sFgzrTnKUcYWvFeNphffrGOUZQqFH6cKEO
XvfVwGSAwjtu6vkPy5f0giDweg1xBmYVb2JE1z7IzhDy4UonpYK3IqZWZUxlkfkl1YyGS/4qL45o
u1bagG69rZHHbXVXRrXfOhiJZUkVkhpWZ3rD81x88uSS0HYqJ4ZBFngZgn6q1YHyHh5GiShzsLCJ
Q4rOn/NG33LOrzDsNc7IrHdfFs8qjnCZRLSPMjLd49MrDgk+JMg1wkNhNma1hDWFnvAUwzIr07wS
28D9AFEW09owLEd5K0a7uRyLQiwqEDeuREMkAcp0wN4Z9Yt0/3jlrZV+ac4ozY0ypwcDthbobmwh
QBfjN2AfnGFE5wX8SGgoovLS/xdnjkb5IFpie+d2E+Qc/vTKAkKSi9elkpI740ps5B2sOSNzrevH
ya3gU5INF0E3sBgnuIy8e5CsRCfySNWRv02chF9s3Cvj3ASLWIFM1oRXC/lc5hvH40dmEgecGYHX
BqDGbnx50abwXg5Q8eSxFoetqBqS0D5G29rYIZo+AeF1LAHgei1+Mdn4FMD374X50vyXiT2PxIVB
yTpHXYamXTq6bFhPilnlmURjvJ/B1BN/MyA8usNOu4ldcSZzooZk5DjgsFP/1p/7ECzoSkLZ8BlM
lEhf+FIhk+2r4mgKKuA0wrx5qe3cy8EUW/W/tjCgrXyWxJ7icjUIhTDUpiUHedhSu3OtZYBh0mQ0
oRpNqnrFN1bryHIm47qZtuR/I/U/ZX5yDh9Lm0vXYnjYg1Nxhv3FFskgRa9Wm2KEbO9r10QbpSWQ
fPQ5OUGZXfjCxbsGeE7WFgzeWmBMTcvksaCqAWGI89a783Q6/OuD+Nzv93gSzasMX1D7mFKa3/CJ
+X40gJFyspukfvIzAJ7xCGqg9/ypAKNoyhHvIHfaYynBnMNsxV36tgvO2FlMM1kddpRdxFz0GhUR
YFgljRRlzWrDQJe4Zzmtc+KBzR5NK2q7h36ZH5+3nwU8Z/ZZW+meLc3KyWShz+4tl5Dzw/VmEvfL
2hAYqm2sFcx4Bi5ecfkcpLwpkD2vAZW+j+zyT5am/0zn1nY0hx9HSEOPheXX9VVBccluKxyZ26Wr
fzYeXSlPDZp8vzJLXbcA8ymIwXAPhUnIBfV7w+6fz09aulq9Vik/FVZa7I6L+hM1kO3sBBE7AfID
DFeZqSXxoa1hrSZX0iU/A4Dp38GDRNE4BDJIRJJrNbLeYRjzycAXGkUcyrzwN3WVTTLxFtre24Lw
/FWUm+m5NT3DRBRBIpqA+ygf/6i4EahieAojzi7Hm1ZaCHDJLDleeLZ3CTesDZLb4ri8cgNy5U9C
/u6qhjVFCMf5kqyJ1g+DQ+iBjtJSm+tvrixXttXlnKVtRCFMxn9Gaohz3rsi8ExIHUFU1QA0XCXB
OZvI/vY8QEYm7WjaqRtYkizGDY5F805qZByETwPUI5cRhtDfTUZJjHE1YVCUSvghjWfXt1Ge93a7
el0+xTd0GQDBHoEhg83Vlug91FpCvX9Tkb0qgJRE2kKBMZ8S9+NWrPOKyoBkN0C6on1KK4UXtuXT
zqhsEkOIwrmn5uTPGpkCfCH2m5aEaqRwtkf1cUmfoj1SHE2PIXPrMzkqda6E/6JK85upln/52I9s
JbEbgf0KTGhxKLRczB66Mxk69WxmSdHmIe8RIgoKmxSpgnO3SfGcwpl5Z/Mk3q9MhxshKZslMkyZ
gvOgzUdqNbUJ8bwhWrerd1a4o5fa71fAGnGnUzg1q2zVfbrLmzzoEkOHWgSDADotRlgb9Cp58+L8
Der+xdvSQzy+IEyvfoTk4Y0WBCXJUb9Z4tifQRaspvX9yME5PzkSFkWUO6YwfCqr7KGunBkkQpbb
GBAu05v511R9nLquXwJklLzB1YFiQAgQPbeQRG+l3+PiUaKSWqakpHJvvVUs3e4F1nld/OlMyLD0
F7R9+THzXk+2VON2a8C8+vXM8zaint/V5ffQ5PJ3Af6h51vaBYlKOuvWfKVnHeoe4qvU4L7GlV8E
NywJnXQz2cxf50hU/aK1wdyIXJnPaBsbsmljfWn8QNzt120mQa1qaURY7+95RDvAlweYPoRnO0MD
z6gHX+LV23d2tyKxsOovr9fxGW81HprF6iB1QmCXOyGdOTodhg+TwP7E12+zpy0FXjMN8795whcd
/rwI/MxmGmGGSBLD2Jb8chKBTLzuie8j95YLlPusEeitpBfwgxOUazjSHiQi17B9iZk6Il1rqwn5
eiNJ73nDIyEDdipH0upAvnBBPAhVP9+Hym0wAH89xzFVmP64ogsG1HioGVpE//+cGbW3WEYa4S7k
MWK8hwibzNmirv3dz6dXlWDpRpqWSLOb+eZT7TfIKxIRwqeozDOMApMbUdm0eqH8Ee0lbnSaIRcq
uB+ryIudZKWyg30d5jDMJn05paum95HcQ+0JwrK5+zmMtgD4wJnjdVohEZJsO689cLJx/n/3Tl9D
YKQuWn/J6D5mYpMIN3ZdLU8HMswkPZMEagsVwO5NckSpy+vcrO2nnK0dyRRju9rC59PNGaz5F2uR
rM+1upLI40uyJ0PQ1LOjqUIJc5hUW/odDL+8LKZXVN4EmSzCF0zprF0HGl/yLc8/rr2CgfBQRvvX
v3Zb6CaQMAlGXj2nEyNrUlizpiOMWf5PTB3EO+kYZYUgzJc0AWlxZSxgJB0/5f6ocijciDcVJ0He
4sqMgh6BwBDdnUP+kCRWAP484cNyfe1EyjcSXJLnX2pzCoGa/XCZpcZg5tlnBvhh0obJ3NqFiZ6y
vRgrP/eshzdBKYBRogN769knVebHjRWl0WP3+GU16NdY9JxBaxQjDdvx8rRi2WWbjrbqSbHXpjs9
VPZ4Vny0O8f+oYhRO05t9xzRNk27+q8OtuA+/DZUm2HI5bbHD+z/hxnYtc4vU7apEhD3Ytr5PI9S
4bkgVWccUD18pUIuAmFxxx3IPZZ+EPC6XUJX11st9A5KSyHGnvycujVaKOcqzMggpYLAXIqBIIUE
raLzYdqg9jiONB+DbdjQ2MjBaEJ6rjF7afMK0MtkC0ifxCyzmJf2S6rGCOcBD7ABpfqcgbk9fJcb
kLLgo+XoZ7vnFpn33WhuwRV5g5/AWMlJ51bII+Wkf/YZHrys6D0NHmGpvDBdRW+gKZy2OnRtce8+
nYgZJ+Q+Dr8OJ7qz/ALHoN92+x+o6D2v8U14Mxv+RXGR1BKKegpHRB53tFFAzCIpwTLTr/1vloKw
FZA7nJ7fhgzDRrOXOOkqJXUZBdnoxuV9mQlgflfJLQY1RPw/lBb3im2Odve33ycEYFbBmbyIDMl4
oTvVi2LOVXpjLDEi4f9FvZnFiHrGDhbJ72VfT3K03M2ZZxjyfRlZOpjfcv+l1uiOEZ31S7LLa8ih
y6Jsl3u7pGDkoZlYqbTX59NMWC48u2e0ybknax/kkdbYyO9h53ZmouLxcdcA1PZyuDKME36zmlwk
W71xsHIYi+fl103Pater18wEFrlDF6yQcHFVBV//AuQ+Ee3p4DX+RSYhgPpdlrSPxkqaLWo/YoMc
VsLYPW2zO9Lbo9H+JS8zgrRZWobAqt7Bmd7UBx77TtyZD0v/EsS9T4EazSyyr50OfaTTOwZQbXY8
d0QuNO4zx4Ygn5X4qQ3YiCXnLb4Xhbos2ZIOdY/Ap/uqv7Sv7nqFYoeWusRymkVLlfMrRscv2+hu
BOO/Lzd/cRN2+/QmtiYRTYci1UegEmJR3qJN92XWmiphMebil59X1HE92S4R0E01KuMyzHrCSIAT
mBQVQZ8Nc5lPKChPvK/vR3GWgZNtOltnory/jtn7U6XjZab6MGIzm269Tip9ydFjyqd/3CQgnA2O
UHiy0FxMKOvVvWyH19S/VVxI0tPA9dI2veakrjIQGOETT/9/4rXvOR5AQSM4yaMENolOTTwsd1a7
ZUQIr0/KsBYoCL/B3aXac/pJkfvHVuNCDEigdx6CH85ZNxaf9Wphn83g6HQyQ99TLbZIQcdKVut2
loX/Q8cWZKQACJw03B4NAXeqSYhga+oWOtXCbhmbDIQOqvv9N3gLIUKf+xUVF42HOcxs371GImsS
2oLu7M1+7LCnyKLTt7A6IDCZk/ojFR2/XCDoHCbrUF4huSpe+x3qSEO89aZcjTIlyhuKkf0dP4hJ
rvsz7y6xAbM+SPjSsysVUGO7MzuUWyHmJkP1/rNnf8AbPS43Z6gkP7n5HsMIzwhgdGePht75/EFE
uqDrgwAVH6MNhKcmEF2TYGGBI+Fu/tDGgXv41Qr+XLAWjaQuCp/xf6XfjuM6HsjVDgF9m/u57ejv
wxjNU82QWLYhehQGPORqpdKefzW76uEPMD0LZZQSWHBAZViEX+xmDOhBkmncbRnEbFD6ZBVCMHiT
5gbkH5UIjj3nWbJR4iJiQtS12EZ109PFZvrj5zzDZli3IL0AbAqtTrISoKkkLB93Ooi8rvsPtZN/
6WSc/LH8uwA5uWWmparfQ2pd7G96YK40wnn1fu3nSS78xyTltZUsk+r9q0NOxjxBJuQciKVnCrjM
ZKJd++ONTXSMG8ZAwwKsa2xu8G9a285UHYfgLWvrxEi8nXotvPI3McakVIhsOyiiAUleFhVgOX8c
lJ2WuNzkhlF0PdD3G9TwviK032cm6Ep33QHzFdUW11iROxLli8g7VCN2RKd7O1VCKEmWrHW5IZ47
cohhys1jmZJUSSlk0ninGDmnD+iTTRxq6HXtkFzhuvD4I3SjffnBjoxr71O2ve4xunIAwmS5Nv8Y
k9s26dUdRyTo7pWeZUjyObvG4yHO0iTflkbyeghiTu8zr/jy7njSerNyoLx3cdNKHUUxBrPUhBJi
JF2brzd+16xpMXcpjfOe/ZmtCzW+tPoqUGWm43yH9Nx5a9StJ9SwTy0hvMV3TlLIKhR+Ywf9iS1Z
yF4LmhH4NuhIy3DVUiJgiYaeVJLkmmP/lE+Nb5WKg7xXSeOTTkstWYlOkaZ3VyY1Oru239xSLhD6
V7qnDalnqmL+8hzCfLqDNP9XNukSuM8kiaPxlN6RUeiw343ntTekcNfEUwXdbhaChRGEClP5Gn6Z
ZBr4EBxZPvGfqoaaLb7PrnjeQfsS7sop5RMbFketOW8Ont1G8tTJSc3LIfd66x0c7bFHjV89DARh
sV2pWsV3u3NtWAP69+LJr8xfpqABlESLuuRIz88DFyxCge13rf8wOnJHRhqTYf48Gip00llrnc+i
9Z9ONkZkZlaG9WmSbod4nzM4R68ZjfvkgW2Riq6VI7o0gMPL5giShQR86rzMWWa1d8HAkeP6g5ff
/oRy/4GHm48XARm4f9Kakx0ZXmLTG1+lVio3A5tfFt345nayzB9M4yL3IGVmhQJfGU5FwZwH/HMr
zF8JL5yUt+ql26bPTl0/VepCBf0q6eMAHYk/aOI04pOMjDO9apY6XlG7b2ttaddwnUfXmXJVAykY
jMOkyJ6gbXy6bPVvXkK4SthCHpv92bMY+PlW3bKGpAiaPQzA1rpMf+jqD+Exv8FTsrQymy8/BLfx
M5Rl4glZkDs5XySHHKEiuugFPXfghC3BkJ5hWrlVOMf8m1ALM5bPLWCcP9fymdXMzlsSgf7KBwMI
QDY+N3VIGjOffXcdNS1p9xLG5ELbQX3bzBDqkquc847ZutVIRcQyectMTuc5wTMtgZ8LpYrDp0NB
Wb1kxH91vbQu3/HoboKTYVjKc2iz4/Ug3oaTmkhjsa/hrZ00cdW8byp2woM0yHSDwFpbdh6S2UXq
+D4Exa90fHmBRSjKZMMLSeFiiT8rPbww2AgjmWvbjmLK35qz1NCa6UE69yYh8QPnDjvmH9HfUGSs
6pqP9ST58eUn0anJ1e1Rec9pcrn6I4YxXQV8+bA6rIFccAGbA7WSOhiopoY2ELuWNGVWvzff/6N8
VIazTkRlfk9dAetCc6k2mNekdytfKxfJyVOTyukQr/C5UOMMs6D2Mq99E832q2fut6ziXnlgYnYF
iK0edTqbdF0Sff3m8NFvVRt8MtaSlYcZjlp3LsaMFT0VCT+naN8mTVJg6SHYY6A1ESqADbcZlbBE
tjsje09gDGiNrUxD2Cz05iw/yU9dEwL+t7RlISGkg75jrBVOteUu3tXsVvWP7YSEyuur23satdC0
AiXsRT/buY9xvhG5ui7VWAXZgCr670VoTnZ+/zR5PCIeXeAM8eEf7Ih1iaFZN0SpMf5mpz2YLDGP
4I8dJG0dv6mza1r7xIods+U+5DRq+yDRyhkAoD+qE6DomKcA7JxVzuoeliSQ4w3aXnC83J+dXRy7
bB/sytOFTyiCQ0Z7zJD6nNebJDcgYlxBnVZkA4w1rHUTRqOzdnYhW3THtXpbpPY7xUHAv+VoSgHS
D2GaIBVA3CXWSoNXGQacsF0LkqlESnzKBh1LB+kmxtR06okNkhtDOZpvzhFMFRgiygGz8ubcYKQV
lF+DBzqy2dMDr+PYZWvIUqK3+ejT4qCXZmecNsEWmHbo8BMHRO8VDCM//3nyyhpxUBHZpyIpnPP2
DPMbi/W5vTy3ImdpEyCpB3U8d8ESUqFK7gBrL6xKBj2nKdhKCIXRIBFK8aUj5/gPfIXKWhyOdsnY
6m+wC/TK/ARZdgMuonfVzC4MFl/yWE5AfN/c+VT9oeQe/MX1/Ytz7IWwqn/YUTw7tkWuM9n/ASKO
l7anAgpAlI0A7MNRxcCf9TeB7LwiIc4RxdBBgI4llEkwvaI3cdLfdC0pvyNYXS4MEDp+0f1H3inr
oeq98qrJMe7F/6yhIjkf2YjTL4V9W67+AaqjOMwMnfiQnSW0HlOFnTgasqwt1c+iYp/lgzae7Qia
pd8ZSswjAHBNLeafzwxvJGQC7VBCZShh2uvoSvieb21Z+5GZjcvjhrObBcwi2CF/cyn4Eychd+cE
v9DLhx5GqBvWCRe8jQdyjw/DREaqlR/fcW+Jit+qUdNM2ZHoLuPb1kKAdntjR15SWCyGTob0dkfc
zyM1x1aaJQaaA1AKKFLRwnrAP/9cKnpC6h5QHjh3D6QYMm3GKkZBmOVnL8b+pb0RtZepK4BaJkTR
HxU/sznyuvoWKBtEPEDA5Jx84EbaxmOib0FXQwZdBxZ4ldQRdrz/F6iI+C3GLZNqyO9VUhQ3DsIU
oBLLxn9jNKVPcWyElHOh4EjvjBQdO/KkrBSfe5xnnl5ST5no1hDi7oPbMJt7txNrJ6md88Nt/vl8
WX52/8/Oi5c2ZMe3/sq+naQk2B7TvXgG+jU0pouHekbepMH/30zfIvUcqylJBTK5m0+T/Axv9EwX
HuOl2ViEqu8Jtn3VwZJj0pP23NcSZi3MI+7pI7jkX2j6s/N8jqAmhyTsiwu2TXWP0eM7KeHPnMCy
+aqjiwVoRa17sN0BblHAi6NfQ2fl9IWUBuhs5QfVhCKJwWJqh2cLgqRD6+UXO8eikRy8F84B2NDH
1zXuz/Tgndg4Vw0kmtQ13srDrIvzRaHZxB30ifVNEiUg5v2quZfZsvQt/brjoSJpGi4mA3sweq48
IdVHsz1x4LgyOxIMYuv+g0Js3gBjdfIkq50ygzNGWWSd22k9tYhmsBPG7Cbyjt+HX/vJr2NJBsCj
ymH0O+rewvkFX8Gq6dg+RatVT+oYkY1RrPSqHhVeiaI9eBM1/A9MMKNh8ogmscku8fT5X8PyKP83
UyAeIV6IpGwabDB5EfC6NiOFeiTtLnVNxqdjp+2ANpQ+jxG2C9g9fG46GJoZCjR9yPb28u2sutYD
m6x0Des1yy/7zAlJgv10pDn4bwUVCf1DHmYmn6bieTiTW9rwgnQlYUjgOYClYPkYf/08AnAr2bvk
97gMN7US3FuhlK57gK/cwgj0W4Q7NKouvKxqoJ0sNrA58oNgJ1y+Q0RI06IrPNK5D7IEpE4ZF/TN
o2j1oMwXJqr6NejUmbD9WrxP4Uci7J6CITYtwTvCXoLPbFqBnYAol7hmUeSmolBgg2BoUVHd0Bpu
hlLqUi+ji3stCokOHgdVUUvmIleU41sjOY3Rf/rullc8Lk3G098jtDut1QfslhAdLiM72KvgyqVj
KkdJL17nhaGxET0r888PBFdISShmyhqTB3RL1G4onMPYWzkcbJD/zL0x7TjnHR2YbAZzmOzs/Oe6
pBAvUp9InSGtUiglMkDAoqn4ymJsGysaMZkdNfiwSN5uZ9xgTWO17vBMAkAp5yZ2uqO9iEYMCgL+
FGzs6818zT8nzlpl+y2FUDYs4+x/EYFd8uLmhCpbkX/6CM+ttTeq3Q3qA3R4XFZpcot5caSddr3l
Rl/IeK9YlKaZofWJmzox2EqJ1C/aK8em7n9U+VRoDapSIFxNDM1mWrYztvcnoBGz6t3CX6lEBlVS
3hJzeo7870qdw0ezMnDhz7EcjC2UO5js+NFfGJ8vbrbIWgEJW4jBeJtFCkYlMzaaKfuTYpASxfsO
6iD6vY/39Lc84xQlN8izp/+h7XSRxtHB4FicTurycFv+GC2arStaqyB61cDkO+BkYMVemqr6d5p0
upPxcQlvUHryaOwR9m8FP8mj/9pmlA43OhRGGdphThQgwPlHpsMt92YgE53Y0+Kzt2oTq0MQIwnr
1BTWvbi4oFmL2b+78j5E77DHoAyxjZU2xno5LTHTaFk6fg8xPilq1s/+ftyabvjwF4SveOU3nxEr
mb+Xsu+uuDb6a3xC5igZWHGyRMUM34yOexFgRctt3sX+Q2xrC+QGsaC48qH+TEFEJNruct9Op5SG
LLOLl7phqEcghTcawLFeQ5w1aUJbOTYOBca2RgMRI4d1/Akq+G9Y3I/3MK0zx+V23PeIszmZlcEv
IENf9s98m5S3Cr+Wk9RaPJ/dAdNtDjkDk1cC9nwIf4oMy3U163O5GDOAuLllcdAWU8iWWPLhp0Am
42GmpaDJ0B0R4y6d1bRPwNbPepgKAbz46BxuU36LhQd0pmWUOlmYq1BSQEv1LAR2kD2SNsh48iAl
d/zAl4e2uuFC2Kw15mUK16WWxyQWfJpbeDD+TUyxwihHrlkEs/OITgvSeCu7S2MqmTej77sEFS3T
UaYvlRZ8MX1iRQjyBGLITBskEq0heplyo2pMUGjc3dmdYm7axbEXpkoCuwzAKInNp1Bbo7aSgiyf
98YCt9ETTU6n3w7zbeqhEzq71/zC5bn4Nw7Xm6eyiK+DsFYHtX3gUdunAEovk3cElVoNyI6k1qiF
z/T7P1NhZH9v2VvOScswrc1SS5UsLb06hTCwHiC6XsfHaRMWdLtJGzRr3HqrWTsuj+B0/FyHTMk6
POYjx7u9u84ITWG2kuBWuPJUIVqTuF6rzYAxVu+Wxz77WuCJtHKqbtVHcXrcaHhY4YntSZTrAAkv
UcxnG9aAQ7+TVxGaO0Uk5GlvpT/tE5PquQQD0AF4Bx4Ax7QZddymOH6fzeIUqrPAaqEHbHcNEFjV
0H8XyDGfIZ8B/aYEUJyGtIizrJhfscBitXeTNurPylPMkcu3nGx8/kg9WlV0Sg6V1nH3W8Hfx6My
qVv1ainbKpflQ5Bik+/TEp/reP+sPKCllrYhTRh4UjohXtD72JKio6s4WBjj+tuQtBIFxksp7pnk
dlmkCc9w8n5/fBITFwHuXRSpu3A68bjI/9V/SQvNsUEf3u3BMMkJjoNbWETHIhc6BHbOCJmRflla
ShTc5AroQepdb/K+1DR5T72zGwKu0lFoFctXub9OEloA8MEy0Sz40oksZr8+olRIDfqlggUJrwXR
3A1YWMt0LNPkgY9Rf2EvIdl+9apIRXL2mJdREZomVn9nZVL9+hEoBKt99CwhPBMtGYL9ZsqzGegI
pIKOO7zTa/5xca3/ASOW9ul6l8V6AD86mWufldtqI0Eh2Mz2KjQDtb3/Rf05kPT4IYCtTkhLlQOf
WcwLPts9+6w1wijVZ/PwfBCrrNRlBN1A6ZW/dbWHl39iFOlpJ7Sq+WzLQ6DhrKT7QYV6qDDdPMH7
rphqWiTSfuPYUAi2wmGwf9yrpT2hL5ZecbDO5htMqZCSdjWANsze1+AGJibu5o5K5imrAPoRtzDx
1jjSwc8ruYMYF9KcEPGWe3HNLbAyNnh+u04aTzMmexxvTQXUVvDv9CFJvLQ7qQEIF8zKCnD5oIs1
vPyHjRgIwUOQP2IY7UtEdCqaTvrNZ0VV55hhMdAAJfkrPZzV6jj/4P9vtHMmHIVJXwEnPiMnkfDm
z75oOyzBlnWYsv7YdPNuLMi+lfzBSq/P3rtTCYwQqK91ksgmxJH+eVqR1cvXpj9rTZ3zi4VdGQ3v
ivEpTAYsXHALpznIQjKdyZVJeJpP6VfB2EPhO0AYBxottla8wZqvC05TFfJvG9Nsqn8oKbYYaWT3
DtSUpyMGQ1rmlLbPxLg6sD0oCAjfupCmQGvJGNmFkPFcKEglZSP4HNF9WSBANcCiuEO1KVNueg8M
hlpFyFJgLPY6viLneNWX/j4L39j5nYe7wW+pdRf/cLNthvPFF12AJ8vxxJah5CXXEjklLNPtoBo8
oGSrfrJsugkpuXsHgLgnvNmYpb/SbS3xC+P/zmg5aYdFvNHNewqh2bcN2xMnqNRYuNmhoikO9V0K
nqDF3jRm02bEAF3GfOUuJ96Hwn0I7uYEoLntLDFKkCxgATaiDjc28lO7ZKW79+jBmlANTFMETBtH
r2mJr1UTdRoYv477b2crW4ETigjcT5MDMDYl4vRKDw6MPJoXUX0zunugfWC99Yct6oi93yAQfyqU
JhCmo8GfBWnWcZWAolsgZ5PKgKqeBXxE9tzGxkqwkctyPVXbg8A8X4tXhkOUbwVHKHAbNb9EEi/6
o9ITO9ebJ2KGCeJ5X9XgB12L8jDTSko1IMlccYYmYmWmjfvc8y38V5PW3HBn1P9MHmcNeNtUhrmA
o2L+OsVKlBRA1ve+yyEu9GMs8FoMvWdheuK1UhYEwZ410wWT7s3jy9OTiSSVdMFIRgLorpbSmAvF
zj8FMXsDTNdOGrJ+9G/2ujmMvCnzm0AhfRahqbzD2h13z2vQiM0DcBIIWoNDzlgqwsYoT3Vr89O6
EfPgcGlbm8p11qQ0p6CBAgHfOqrcIEvVVJJ9sS9F/dWNvCsF0UfSYH0qFBste8p5NeKwe/70G1h6
7NtTaestInb6l0K1ac8eUQhr0/eTGAKrywiuDCrCF4EqWGiNl4KoZrS8Skd35cZeschxEHn6P7zX
FnqPseWZ1njMiN9izPebfKWIfc7ZFaEC87o/rUj8P5u6SaVsBlJd69DdrHu/9mWYXoFTUCOcOmCH
Qfjb7nITG5tMBlZNjpZJQhmUqUW92igyvCiprmw3dvFDrSZbjK/1MXh0Np1LNH/hZnntV8Mhd3By
IkjNmV2QSEp+G+PVHeRIRXO0oijIVvbHXWaQ2LGB+4Ekp9axxJ8mQ3CaDoHc4pbYjV5fmOBQ1Qfk
qE8y141gX3l/xGx6R4xBDFaZ3qS7RtaFCF6YV817YzAAlSc76APTi68qFF/YhPbxc3VFM4UrSd/K
eXulLxOod/DoaIABPFwMv0HW5JyoQFAbtqiKa3vQ3dk4xEE7HkcVri9fyDVJdB7kNrZ1YVruXnpY
YUSHVH9aoEpK4Va/E5LmRtGDfYnMTc+zkltxmZ+xhkNIiZaVFmV4XT+KhdaDcsc7IhtT7DsleHAI
EKWaIPe0ixryaguuxeTikuE3KGUCL8C7b3YBeuCmbO5agll9RFmzfAjjQ2pNGjPipXgq1m7hLmXv
1WtQfgA68/f1x3jr0cog6EyjvMj3YuOn1aXtjuWfmQGOc5d15PGQWe6W2Ee9M4VpByTffooRoGNe
mlTDc2ydL7haovY8ZhukTiCjTc4BPuNsPf9vINrJW9qBgMwynZr8kkzdqcN09AGm/LbEn5Jg73ii
Wm4UK/4Y03of4y0gI6eSWEFZ0t9tJlb6/1HImWPD0T8SHtP9RjZuDcIxJ03/OjiG5Kfuxn5DJBfU
NcKFprR1wMJrNjEQkGmWWf4gC9S8fMoJbmxCdUNWAa2SvSoS1naBnBMqZQC/Hg84MoZBG2QwcERi
/WtvbySAIPv4YQYuSJbo+fX0EUACxPncHVvpC0/8qn4OzC6HwB2qIzCKL6ds/aWkC465qgQzz+ii
VATumORo/Ivi8sJwyqCphWdTBKRtk4lcX2r9/C0goAydJw30nIymFmqKP1ZuZ1uslzNG9zXQUVA5
ogUlKscM6nzeeail+xNDOFw8WF3d1VaaTmiaMOi0LEw836mrV07GGf4FK0b6bdoDWp742T6G75iW
DpXeDIQYHtV4RPX5O/hwd0ZMe4DTNE1drZYblWUzCrT5iQa8X8x1ktmOoLPpGUhlfIYPdqqpAsO7
+Pu5ATmr9yGkv26+aUShCSr2imq2MjM1Bhi5X/1JIFBd8dzpYe4ATtmYn+RLOx44Q+MpsqKsFJZQ
cIlbcxzH6V0i3QNAktOacUj5ZDBhTDU1gdIH/7Xg9+tuel0JEQXnjFRRtUYT0MTHSI+aEYTyGndD
BNzMMbwX0Rktt+z5mm8ebKP2Ai8fkImeAKKGb3Kx2P80dhaFTCqZ3y/I1tPGSU+T1qsXaJYqtVfz
d4eogOxtfUNRpCBPRfxdc3NO8QRqp/UqCLk3/pnvJtyA5RvUBnGulIaxPlRpVk2xuTbxSSuGwL0m
E/31VzGOfH3d9aK1CMu0O0e+sZaqqIcj/UZw0UbSKC03QOFDVuJAUVGlntuKWEzHx+a1j91ZNODW
PYpPl7FKqHhIUYxrUsQzcxs3AKUb0tmhMWy3y2yDW6rMm5v39WjJ8RjLV7+L0RQrSwhBp0mH7hzq
mYXm7rLBH5WGJkOJXfR7tQzv0lwXdMSEtQXvntRTJquRYfiR/ZPGMymYP3v9RpuuGxNY22RNIRi/
XJvh1tDlh8bVnjAt4YjbDpVjLRkUcc1hP9vf6+kKnRoT7EI+ZmUks3PjEKIfUbLZHtxLxEmtQDVA
BRbmsOlRAyQReD3t/xNEz5EMRZ8MHOzoOkoQaRsMeInZNTg774jAQQ3tUMxHn4FvbCpIh6mFZ9TZ
c5G7Eak95zNIL8gba+jvoIL1spXcnWiAQlRx0fV724cSosvVY3CwAQ4WgJ1L55wx9w0ILscUKusO
AgqR95gtQqYiLg7vBx8eABLcIvy18LfAy+/pVD4dgG6JoeBtc3dUy9hN/y2vS2zhr/urm6XUgbuN
RnX54h5PGX9Vuc1GjqOrTO4gb4nUuD2j/HMM+aIVG4yvlHTRCxK/XB09gl9kqdIClNQMo1rKJ6vX
Lb/BpicOf4a643LUOkwtsDdwlvWnf5CGDERB9+Wo4G27gRQxqWgeuDisp8qwxS3roUclqU84dc2U
R+wX6BJWRFzqRmAQ2x1bX2ugrqJ0N+LrO9n6UnMMBPXR0CPPMRf3GtNw72s5DaLWbDHdBUJiPzE0
QZdICiXgdY0VQ9oGLIG2AbPgBXjFcEY2N7AqR4XSnPaM0A1mIineWXy6g7vJTX7mJn7pOvahFx+x
LUqF0C6nurWPcrbuFQDNjQplgwZrbSXvJvhOhOZVDIknS7xDWEkyIIatnHnVVFO1ZVXp9T/ILVwt
kAnWKtbjMYd/xlx1HVF1P+lGGy3EUYpqAccTBWfVcQqWzTEc22Y+/XsiETomusuZDCw3vOV9wgUF
f2JWjJFbTyAaHa/0baJjtN876LGiOfbrzD6YJfyZUy88e7kWL5qYw5JbONNTjf07Mf4FJsw1fFe+
jMM0QOPbo64r4tOCAhQ1FELWurCe1WYNLhsL72lTLTcWHBllUUpmYGJluAxkuugaS8l2Q9LCxhIe
Trnmh013EVAZerCxQ60V80r8XIP/fYTc4k9u9Ek92b6BYEv3H/7KZYb4I80DgmtdSrEVnHN4RyTg
SsCUxKIx4JfB7Mz/m3r/D6pzerrcPTJcpRSb7U68Gy5ZSCssNAcRIPK5DUyoRbM8pZ+WrQhAfpW9
R2WAOQirxbwo8JaRGgbPgXQrSKz1meccJrBBhA9TQ0QPHsXdGs5mpcmen/gzvQmCyvFQ5iEE3v02
acKoVAK8SCKft5u3W0rHbiysO7XLZqeI72Gp+xusTGXWUoDlJb+UxBoGWS5uxZyAi2Rld/ZA62lB
BaB2uC4HRqgZ8KRAOyoN9E855+auwhUNNIrIr/zE99irKaQs1dNPCy0wb9Oa8QNuVqS+GgT0dkTh
Rbk1NItaWI24NyFCFerTyNnXK2tKUBi94v1cZ2IfOiHnEWXt9/BQm6+xbMOIpxs+tHWxZEbCe5BD
16v6GS9tj0Q3IV7M2FfxrP2PjrJhwcfmeRQInHn3nR9Li8Ni6bC9UPPjqB4tQrYwsDVuThOr/CfR
ge0ZieRiTJDO35Bcb8H6TkO7ZWkj6+1qR7VP0vmMWdLHy3OjGJSyjYS/P1JVUpietGW2/BJvKJ06
AY8NuQcQYrRGxV49JN6dZJWR+2nGhpd3NzQkziXiDdNmyaIhjz8lG6tA6H205grYoPerx0QJP1da
UC118ydheMWlFc5vAE+6bkV/A+/QTY/Ma0r78tqt1Q4icpYpFvL+TzNawVFLCRei0EgmDFYAjOEa
t+xVNNgTSA6DdesCT/61uaZgqGLanREfK9S0Ief0GpDKx868GEt1xyyzft5KBseoxUQxe2LlDVYw
4OUrwSTSQgFhBlzCCMSUVG7S3yBe+IIuPrOkQhdb5N3rbiwVBdueUMRZZDKllG/3Gd7lseKFAmRy
ZIJ19+++HOYKaVWlpVCeR6tCUbmvCkvOV/wyfnkDqLVkRfCk77EZ/P32HdY+NCRrecohHzwTcQvU
O5aIXddUQkeaYwsItW4wjrSLgJ6zBGmOiU6JzT5AVhKLenJnGonVZSD5DLW8ORJo6Z6Uzy789q5w
MIuR2YNH9IEmfeI88f4fMoXojIG7GqTTLP/vP7TJE5iruhVmsyF8Qda6PBkEMv6XhWfvyXimdveb
fgQ5ViXUU/UZ03oyZ3aHMPKF38OdRz/5js75J9vr10pkz8Z2ttd2e4JgYsUhSRdNfDTIFh/oCNjU
fbB23mN/b+V/eyBBWxKot1SepAGN8VfxwSe8M02rfz9YSbYA3nTXAdGWiatjurvoILbbpJ7llTLc
taBPfOnhNtFO2GuB0WZFWzxjk15KdGaFjF6lpf+eS7yS6byrNAsv927yc9Yo9fknEf6pzS0OTmn5
+cV68Sn8ph/g3n0BGUR4XUps+OrkDL7XcLftgvqdBlD/jlJTcGQwkloBGDOVPYqPFMoHbaFkfMDm
zJcfm0e0Z12Km4XabEqLGwCVAHasJ3vanEI1gp9noO8LzGf64iGDC0sb11o4rYSBdgKpZeXhmPj9
LTQemOxHKMS9SMJ35/VMqzFyQOSiyFyQqsGZxm0bvek8y6cEiS0BVL1nqPgoUHQ2LBOPwc7Lgybq
5zVrzp5ILW7JAaTlwb8NuZmng9d3DEUTXGn2oNoBLF00X09Mpab1N6uU3WBRAZaOXjVZ13judMt4
Wr3NQ9d63hR+Nf6aDVwcz/HTdW1TQK+0YGfjSS5OhX5CXm74TD0Ou7ayiDkuknUK8/1YqKRl8KDp
hHLijg+iyvYAtfySLA9kQNCMX5QQenE/4dTyRUJF1krrwwHNMBpzbrp1IrQPuu/Wt0F0JnxBjyXu
IzFAMyw9vTn7ua7VM8g6mRaxHsDH7Tf+0XNrW2Xl3oCWWXbPmpP+IKBlGC1M84loXRN0rUZ++u5S
Z1q8Vn7OBtPR0jnPk7GNyOBMLrDRmF1AOg8DtNhAlLDKUKNGuBR5ytKMiRARpzv8BcwSJKqNj0X0
gmg/VZX7SsR4SbmfEWqxHu2WpMx2A9z3mqk1Rv0qMbFPh/sfkLE2vfmA1BqWkYUxFNHS9RBwsWEy
hW+HPvFBomgANxfKVfpzamYfKMHPiH2JNgeYpszZWKXaC+NTzdKXVtU1ozTp2sH4XTfEDB0CIxCu
wP3KKAbwq/2GxQ4W4qZM5MtHR2AT9B2XH+2eX2YbqrHR2zKzP4Z3U4GcEe2bQo7H4JMy2of9MEN6
0kNvQEY7271GbYuckoKhzFuqJtC5JE/Unl/QWxzQeaFCR+ZMKsOyL13yeGQO4Fu2QII9dk3DuqXK
YYyVA69BsAGeDBdnGKKcWkva7M0UpHKkJn+XpmRo8GQTJpW+sJ4F5Br9dx+u2vpxN2PYSWbbXgnV
lVT6ZmzqaV2yxN0lsM43r1GYBjjw/a52Z4ggul/2iNZzdGiU9AE4gRFcZmgpaEGzYn7IM3dOIEUD
UAufclZKWSB0MutACtCdqGhd9tAajyh8+/yVhBeBgKeUAlZFvS74ItTUIbPIzf5Do3MrGjgkNbGE
A3W3+AJtaE+GPG9QpYeePbaxYUbEUrLjPOBCwIcHYrWvUZpG40C0tqrEGe0We3YMWKZAAM2HJel4
ZD8A4hnOMF1LMhuqfep/UZbTuuFlaNz0OKD2FjRa6IYObWLHyQ7Qwov+sdctGtWKKCD48y6rDG/2
Z7i3VWlREzzYJjQtaRsqHG+RG7+y/pArlzWbNZ/Cc6MEbKv1n3Neybs5r9vjTl//+vBLU4KSQh71
Lo5eR9m0rp1rm73OmQmixP8sH/Ks8BrNUdVHW7fVps4B5v3p9hZwvW+Yo0xza3OLSJA+7LwjLwAC
BAjtcJ251uSGrBkVMEbDzIdxN39HOqitnLguSgtFvcRfvUtV6OVoVEGVmqoGmtCfHWf1NBvfU8a9
k5dKcHUZNopuVOa16jCJ9GzBkgRVUGsUAP3dO1k73OZog/+FeJJbeYQa7z4dhyMzwbfvXfyehq3R
joz4vOp9FiDW9Xa0rkSGo3Uum+w91ED569qPSCLl4M7j4KwEz49ttlwPKpyRK4qPzzHphxmw0toU
I3wbW8Pgd9VCmULnshz63LbJVN6eCelA+Pe7LYGSBGGeOinpIvrFQ54kMi/06sDfNvQ3iNbacoks
fLz2Kg+TtgET/nMbwQSLtO9zRSBc0T2Wk9aKhMpkJnmnTzBnsJed54Kk6vkAFbpI7BkOSml0tRMV
jDaaY/HvO1+1Ah/WGzO+ChWSR16la28esMsKRCJt6GxM4BJ3fypPSeQpaB9OyPF2azWy7O+d9CJn
vAKSGzBN8NUx/bfGcZeMHZQ3hbf+mX6Dw6SX883FS2FvNffWMXa9EwgAoe2oxg4B5Vj/v8A1Drr8
b+L6nyVAqhvUTNzXC8VAwrgRebd7Nyjcl/kuZHvdytIJg1l88rbiVTznUFdLTGBjxhtCJlpjCEux
ol7IyoBeUnafIdiemmBurtKrQKwTgV6lkpgsBxXP2271qiYjqwyjSHi+tlMd8/Cx70xvFD2XlsgI
ZMNw2ipVPjmmxfx49wIfTrywowmupRaipS0g5bqxPiGCmE72lfJ/3GTufKANX5gnn1w4sZzVfFhp
XkUqgeMVks2N+gZKSSSppNInRomVDDxk+yH6UtYxgRGphbkEZdkzXR9r9r0wTEVXU4JvaVs/A66G
LsnGMxYNkHn+n05NWbUbqiNS/SNqZvxdiwecKfOxS0f1ITnzeJc9uvMv/Yollaxa0kBYJgdG0XcM
b9KJeEMosJEIq37wpv8WRaCrqZfbvIU4XLxURBztEbYqNhJz08bjN9cqu9jNLiVXra4U2jCP1Buu
9PjDmZdWHQbaH+CDax+5HdrpkDg6x6fHTP44TD/y8981dNpRLndq02tYOz/Ph/dWCKPgtba3IHPo
Wy2OxTYDbSAy9mhZ5toml5T9XnBJLhkYivESJO6QLmMn9/VpBHVu2yj/HsE2Go3oyVbIVk+/KAbf
QK6hTiClrxYdKQf8efyL1C+nV6MtdWlRHjy/W4l/yMzBR/YOQf9fHQpz80GYka98m05DxBcrG6pa
qYHXpY9Z8I0EEtxcqvksoseZzTok5VzKgrgr0xmPYHCoE8pxOATn/QVnYdk3hSBxwNz4F+owPnxE
2yILYipg4wG17wAtbJkHGu+hfepgKZqlxH7Yi0s+Or7zlVNcnT7Mf1ln4I+r4WjP/tCYDGlcObGg
JgLB1jWdHu0ByQWnXdnMVQCp4v3uWf6TWeIWBhZ/QI7MgsGTYx/plOdEzvL7cXglHb63trZvlnpH
jXvBNJfO0ElVHLO4d3eSkzxYBTGDFRyJcXQYfI1RXxxPnIQ1zI95Wvkh2rdK1XHzqD0fLhHONy3H
I50ILpO9O0CbHVeusmdvnPzq6Lk1cqtB2bCAARSfduEcu5WI54JXWr9sl084Tl+mSBTws+W7L9Jo
Dn6JyBLRjfSasS9N8dfDiYLI7ntaoNq04Pz6anTHboPFSFofwakUdokNgAMC5rUhUnWACaAZydi6
/pDfR+8lcRnCHFJLvpoMO8+MdQ+FNVjl7FHmzNzqD6UbPuOcVG6PrPgDG+HxAUnvNf1cC0Ev/AHk
bNwBfo75r71FyTCFZBrA1Ep0v9CXrO33lUAU1FC3DsV4pnyL3/Vyx07Jnxh+vrQr6LNLjfrw0bF7
94wvnRPLlaYHEWVQ3guWqQEoBkBf6ARlYL+5/17plFNYjIbZwRLOpkt6c+ZFNEr8+Ar1dDg4s7GP
Zbbwwo2Jl3hyQAz96zGahyMbYvZT3PZ65FdVc8XT6AzRoKNGHU9B740kk+mXJGA2Gjr+F35/Kz12
vnUJGyfSQq5ctdKQfCP/mN+WzZDuHxCfPAnIEpQmaFCHogBDQuJ6IzpWw/Rcj96Z/4ObjFm8pXJk
uu+iBA3iUtobpabMhREtTfDURnlk2KFguxc8Q9cqeZglA8/aNJpKnM9Ddb8d/PDgpfyBpfo2wFGE
f4JjHxB+BCxLCbvM6sCoRhTaxbjKz5Uud0CSw+TChL6OLHBDpaUw4wllBHjKx840rBlKoyqyw67R
E4eVouDu4ZeGtAaquDLz+kZqUzsboPplhNEum4w1AGrhpkn5+Xbag+zgLrQ3aKK20lL9PPRNGY9S
xCFfQGQhrqwSo8usGKzsi1okOlYz15aGbhbz5geOIa7p5I920rX97VgHFER48kq+A0qvQB5dEjnQ
yoFU7dAdowFZw4Cb9iWE6ZIwOFgquoxJxionujUN7HC5VYUoR6ZJFikB+OM0PZOcICeAEy4p67rm
0gmbaPf1eyXpn8zJH7y0Z2ubbcZreGA62Sk6KCILs4Q94DLzRwMzCTRU40GY+5mdx6htizJ2PTXs
yTMchc7ifmPbrkeJws3E+m9H+A3R93asI9Z8h92zOTSPfrm7dBWS3dr5EGdxXLecNQs78udbXhe6
P1NSlQ6jSXFnRP4A+q1x4DLsokSvl4dDu7Q9KR678AzcYZf1tI96wf2Y3LbL9IMbEfY181Go6pgi
ofY+p1y4gmmH265cOAV+6F2dCH8MhDRzfQP81V9++g3Gwph8T5Nu077A49ghDvHmexXp52z+ZBx+
cHPp1Rz206/WiP2WMisgk5BSX2wx2taoaBkDs5UXexn1yIhCRAKwWwdsDGTwUWi7kouPtHdPKKbM
NskVnkjRP6Tmuvo3IAw1B2GL4z0FCj8SlN3JipirBQ1AQe2hfHUloMwTtMbLE5ccnyYQ94S82+rT
sSWAjQ3koJJPv6wthamUIaCuB7ZHOjjJh5woJ3rJmN7KPBfrpNXpxORBBzktvGBZ8WMFPx28NJHH
lgHXB+FRZtK0nFZmFWdjLJ09G3auIwEIC0ZnpkA0hIxieSAeAQK+T/JU/P08MyhurstE97KfMz+n
3cbfLOOJxvlT28C1LM83sjow+Sgvnu65OvriM6Ofwb0uviDjAs6pgEoav9Z25hXCSgeYLv2Lqp/b
qTTH0MksMAOPmWD0q6Yp1+bb2PjL3YqxYKTwfLBsJeEiNY+6+IMnVa811g/Wzv1wfPbTGpbm9nxu
Hc+IuSEy3sVdvjpWDt+Z77KFMBurcfXF3uVbCCffvgLkGDXk3V+7jfW/+Vx3MShZMCgyBpfwUnyr
OZCMxRXuvjgalIv0s+80+W5OSnqtliFzeECfL5TgGw1N0ey1dYDyeiCgZ9tSVMf0AVv+HRnpsia7
lhB1pWnzNEJH9LwjyQ0tZ+ZcKFjsTWmu/1rwSGL6+4ztsUfzVps+R9ejPfcfg3NKiofW1ZlViDTK
v6tQfGjQeRzE/6HLwNdPwUQjitjWYKsoLK8br/frKWtKP5fTByeNt8kymcET2dTCk7+xESqjqLmR
sGK3zRXk5zZf5C364loGcfftxGpzvmZHqE1Um3ZJLBqMg7FbYPGA7xaiMJCVYBAEksjdguYVqS5f
TsA3ppxLKBqMoMJvOx0pK2T7ggIwTZqcKhyvaxbODHmH//vDP360Fo9yG/kSfhPHF6vEKx+3h+wg
3vdo2Ipab3I7odGjScsai3sTWmn/E1iGwuLMXKg7wmwYDmuG1UyHSE3HXQapKvDQ6w0NAfEP071Z
1HFGMBdWQU2sMYq1klGLLNRsN6kwJdULleGGwh5oqZafARgEamaaAQKazsfjz5Tj/1EcLVJA+xxf
TTK3A5xvneR3SxchC3ZvHTrSDkCxImxm8+ekFbLjes9zfrFKa7KN1tDoAfbOhojoKP1lL0OW3Srj
vGG1bs+b9AnT7bInDlmw+6RRkNkUDQ1Tnew7w+3gHJbjE1t4gCb6iu67RPs2/cgqOw4gMNsxFc2e
mLmKE2UQpH+2sdAPDk+ELgTFkE7CuHFAqLGB/cPmEdnGTsB/7Mn+pXfD7rNpuMBzL2z8H8qbRdQD
ZGxUkhyVkruMlSMHufd7IOyWC01NGdrCLr8fLKdI9ynqtvqNpKZxhUPisP+WVgPYYZERVSuC5E1o
KiLMH0xKSfbfWjDizUQXfBo36HBSa0MWpIVlouxVAsOWYkwT4y3vhrjvj3RfXMow/aAXg4YVywpj
YpeDjIXk2UL9JBrPS8Tri16GMxf2YPSiB/XRkG3nIaqq0K58ezb37CqfJq0hG+kbWAiY2h473r7b
PoSUlp2WPomHB5PHK8kgTEAIDLzp0y4kwdKFTBIwS49Hb8B4ddXwIztHUWpAMbV7A+HTj3hEB6m3
+MuXo16YU5EumGW5oFVFUigesDzOFH4RcBkHbMJU8OtBLDLX2gHEvJqg5DUAFK2/whr17rVeayGD
bdV4xQlQDu+Ey8D3La2RgHWZKg34rFB4Rzx/Rj/IikbDo+cB9d61oZjQJLkDSKcFmqeNgReC13qZ
ADgrfX882HFiHw7VAG//ZbFKmS3OskA8fRNoG2O8gf6s24/hcAqmssewkaazDnXfqJvNzHYP52z9
OgoaZJJh9PHNf+yCUprGL23oFuU7EpCxRmTY+/C7zHeAYnE7ICilXeEtT5xWVJveKAi2EDXR+uxk
zoXJBWE7fR5J/oirdXyj0l/TmFWkBynSlgZ0/3Y8KH50kk0UXMtBIYxqZGpJjsUyekFDJnokRt1B
BtAWEC1U3UuQB/D3kuNojojMyisAkZB1NhGL/VqWtf3bFblZlgmRQ0EfEI+mW48OCtOresor1Xu2
cEhdqriDYnTirr9Hyg8zmQFMWaY5fZ7Zz0JH7qyu23ozo11B77c12VcsNVtsj1n6ka9YTGLqP1tP
Lkpn6sdxHy/Dv5AoUzhqgkNgzKU6CTuygMMDpIhiOaj5Iz7jWXuCmjUsdnCHqbWSvHBbld/QUqP0
TWFUZ1EzN+bBrh1+4fZT46/FmlXl+xHLE4Wz9rh++Ob4cB1Puhycg9v/2a/GqdrXZUbWpaJqHljh
dBX2xpeFjQcyA10oXMtIiW9l9s3HzlvtAcndmVqKVWatYpFcYLxaKpMlJOhMVROqQieMPN9NkyCZ
bX+ygqfLPKrsmutOdzp0XD6ch0chvoiMPSVtTWSBDqjyJUCIRk7pKTOYbOlKg7irfFnamvFQrf3H
aQ+aPflQACq+FPYsJ8cahVs79CVLplQICHjHVi6OPrQ1KII2P45U4FNH0o/ewo9TrisUdMn2pEAg
xDaPnVpiGHImXLzhNAmndgilDOryoMySini3RiNM6M3OugkZ4cRF/TYvuyQ26OFbAd/axZOrcZ+H
kGkmZloJBghzDW3+6L9EPmupVuRdK/5ET7ruQr6jFXVeAGLJt0oMp8Uc9HIikeXVbZY5XZTG4OsP
VFQK/PRyhuhMqsQ1HSw1+9ebHEaVxW4/ti7pBKpEaVH0qMdJDV+t3shH2LmqIBjDPleMq8AONkNJ
IgAWpih0RPZyZLAGUyTRfqr5jxofiRqBGwMrFud4GoBKgzzHQqGhutloPrg1P4eKbllv4HNv1Utx
+r39AwemCfwWK0PEG+HMFUdl/rDfA4ObN0F1xajB42a+nAaoaGvEr1+Oct8OEk2THqDHZiVZ1UeK
zKAlWj7uXJDoku4wINQFILPQ3UB1ctxWERtxQACp/pu9B1HUewsEe7xX2UD2Bj+Cz+0ckpqMjnWD
RHkE+2UKpwNIPTYYmuda1/vd9puVzLRg9hPE89c7Pg0IWCcWEjmrzd+URt7pxk2rT/xBo8bJx71c
W4Q4Hv5N/DJnkebNLIpONg7+QCa7WifqCxcuZV0N/geu1VcSqriKj4wFDR/fpJMfbXOaNafmjUEs
WTpAftOEEikX73EcZKLPWuLRN39ysI/YFgM876PnyevWPdTYZxYYP+XE7AFhgQhu2MU5LHExpl1m
KEBRyiMTVBx01tYIErnXzY5IQPBO9ViYLUNUQt83/blpDQVrbYtlyuDQLjdkrqAkhvlzxv92/24K
GKFwb4cYd3biJ2JshP5sXkpoPeATP868DwHBgYd0jrSM2CNLq26KN4L37bUsrBCmgEZwKF+8loxE
uTHt50FHuGJvM5y/9rQZiaH8DzR1PqvgDzulqnIW/Xbaq0dxPwrmBqjnrPvXqo9kH8+OdFIx98xa
S7o70/PTHY9HXkdvdqcuWkZd40c18w/E6rn55lzttBCUyxah7iPJ9Hsn/m8UvudwC2oF+reHbF0+
Jii18UlsOzcIe8Wu1NIg7TbMXnTM8H27wURFK7/OXHPwhB0cqMxesKT71NP381IXqvYw7IITQQi1
y5/hciB2o1tTNVBBtGDx8M3izPlLk4T+QdzUNEtVdrkh2peOBgvY12doXe4cStb1jKf3IvmJBGsT
+Ww2l1wBknoLdsu98sBWlEO39Ni3y8YV/BAxL1evKVUtbsl1/BRdcASwh7xebwQX64p/XLi0cYxv
mR5/30cDdyaTzOD0iRI+tl1IkvPRAOXk/ZWW0svX0DmiJCUKxDfc+RQ1TpBqyV0aJFd3dAxyfH4N
imEWK3o29vgpzn0RDoiZMTqWi369AlsJ8bVu2ZiTz6JFo5mtqdNF9FV/nVLT6I3+hkqsr/KLf2fH
WEpKo3TRuI6vFeCrlqC9BkrNIj7WfU3jQWOmMxyRoHe2SKloGIHf/aLZ0PURCTLRxsk2lYD+MJne
zMh09aT6PDBgmx8gccXCqJ/B155jKTSYa7VLDoc7kZUZRe1UStH4jhLZqe/jPrJcZBCgG7Z1yLsY
4m3KDGTNmiqOG0AmtIK+gR04QPPgZ27yffsGmdsku5Yav+mZsBipcN4W/8Q/kSUgH+57QJpPYyEG
27WSsS/fQGu+DFTj+DIOKPOu9NHUdLVVxXNzG2oSBaF6+XWRPWrG7Be515Qfgm0LoiNdGBWgbD7S
UpIsw0cqTEcRhjPDcWXzXyTPxtBJ5Li+LvqdfexFZGWHZZuW7ILx3ZwyQVQ0VMU42Fmc3LQoVtG5
eXzsezp95+AzuRblhC2VLKoSS8ASCoyWbBAq4Bsw9+U30MEaEKWlZRGDTEzPatnfXggxYslEAm7d
RydM/SSsuaDM4bx2tFeghLwRSa69aeQogckN18mW9oasuyD0wonvZvz+O1Hf7Ax/CWgLfoSfRcJ0
xVxzpYHlOEa15auRa587Lkr7WGpay4dQ05vQF8WSXALTOyMrYgCc5qHPESRmbvPYfzbwSAQs60XX
Sz9ZkHJLp+VBxj5hlaqzELgaEaj7uG+FNwwCt/U/lTCNJA8eZyMxiGFEDAYjCQsilkZ+u2YJGfrw
nj+Q6Ezu6VUHk74n/jy6xOo465jj8yLHo20JYqqWQHQq/ftVjimZrlod2bUISJ8X5VHXSQWNY11q
WL1LxXwkho7R9NL+/Pj9Ruhlwt4oKdZF8T8kr8gOVG42kXye5dx5fzrNz6E5VFYW2qBYIBEpAehS
M3KyFUBpjPPD+es9fj/WwV7WV2LPqfMKh+1Y5hwgH1I6yC4GupD7NVYBrWQPCcgSPqqMxvvBfsQI
yMVQlv/MtSdnXhRKURJMF003QX4OTOddoQ+UslkGQSgAqrsBn1674rcu6KDOdc/bo5UIXQhyD8zd
KEk3NKtELeNo1m6/Btc/rpaewd9/EctR3kuyL+AJCLnarsIGrfMUqdsQrkAgNbR6pHiwODfLJfPw
B+0ZZ9HQs0/tV9DW99rilOEg2EurKagn9YEQB0VO5Bdycm2SieTpoDDa8I93ot52ZZRw2rqKzK7Y
USysQfyh4wzifXku8gBmhVdC4KuBfeoYHOZpm1Z76YymCjPVj5lGfzUNjcr6qvV735TGlauDU1c1
CRTM868AFbevAqexeZGuFD+U7O6224kYvNsKuhXhpHmIP1PPnCHMIarlkd76XsbL3KePjVmQJw4w
NS4MQsIGQPnjg2+QIY1c7Ss5ieh60IzbJTJBgRKPmFlNcVOfv0oFKWafLVJAFGR3f2pZrZYfIMPo
K/zWcFuIbeiSIzYNSD6aDW1i5CjGFTETwJH17ciKy+2cBn+i56QVBAx8yhJiSeLrXAe07r/BKWW1
4c027rPbHYGAGwmFebq/+OUiPXZYg+KV+PeubxAbYpt7Xptfa056ePyrY13a3kZzlgarSqgTJZsS
wXiYIa5tj3QS+8GMT2uvixXE83Q62A7Aq8sss7fdU3Ne3FPqxinq3W2MnC/HyoV2V0szafq2xfuh
GpTgPABMtIlwhpnLwnDYZh+cus5lPWOfOYKJtxc/kNI9dPO2yc5FfWBNc7lU/hbmFctmtTXThVl7
tNq3hfXqG1fLJ68iXPL8fpIeBgT1jJ4v0OMcmT5wclN0teWO3NlTW43FvN+dW7qmcO5eyRbUhLJH
zRFN2TfNQExsiYEJ/ZHzW09zXzqHMkYL36ZtvCum/KK8YK81KVfP9l/J2o1CTpojPKYN++Z62TGi
9csW0UtOATe8kxHWQoeQpRVrv2ZFR4X0XiIyYH+r9XTHQBD+pomSABZmFO2p5XHcUNXMiG/jMpnl
/Hb0B8yDQLybdU/Y95swW5lM03ED7FN4yGnnrmiInLxgaocrS7H+DgCNdn2ZuSZdtjkcd09sL/TW
UUKvm2qRfEdD/4gyDU+dv9rt3cM3q4kKmY38x10IBp4R1rXP7VC2idpQPkCbgTtzdkBIsOMFhiCs
QOjI14KPtMTgkZYwXlV4HrnPIpYeE/cHwUaluqkk0857wN2KFDSa/gHOoQlpERCF7EboAKLocpdx
S21OItVGex1Kj/TPCU8a5jAubNp5V3IrOZkMZozbaXD9Tx+KeQLvq6Gm/AXFO7BcQwLgRRBnlt2x
aN5iG1ZpoP8fTdy9ok9O5XL/E6NsK7QHSQwntMLLDLiaYFjR5P0rdZO8akva2NEn4davjlbyw7El
iJVcT9FL3OL7MT64TDYEZWyz/4i+YGJKYw8qRnTpUUrgevvJC1Z7myExmPyfSger3Uj+ve+S6ohE
zVUzkuPxPpAaJHw+lCuL87QPMoixBFtc6pzHV+cxGsuO5xXB1WqnhRr1HQHi1slxGx/hJ5pv1s+0
gahLq21tOdDtPn4BAAza9lGxmVoy9ocwYBeTba3+WO79DRqBRLsWz6PYZ+2CIDRCmWF0ct1ONbFm
gsKLt8qGjtlAyyyYLM1lCk+zc0wMRnrDYSFBmWMjpIyLINVB725CKG1QV5pUEXAnGTq5LV5yEkPz
/79fitqR1GEHfYtfPYdeGyzMq8SsCg2r70Q1OOkprEXuvp7Dh4GBA+xUZEAJPDKGvZi+oMyX4MkR
6bZP57bVY/bKN4XiSTDlpaZFoAd3TZckkMBA7rFt7b4AVy/2cXCNyAAMd9h8y/diOYyWS3rjWiB/
KtSQGjQNj4SuoIqcgk4sxDNAS7TiTBOa32ByrhnE8hUGI/cgdkQ+Lu8K6WcP4WB0focT7k5ctqWv
/Y6uUbh1dfT4oC7TV3/IL37pXfE9x0eZSJBM8A1FrRBPDW1ENY8yOAO+WUoa/bRX+ygKkCiGo2Ya
ULCjuu6xC3l7krEFGb1ukfA1xdb7mpFkZIA8z7cyAmbF4KltFMbbDQO1nZuV/0Xgogkf5iPz/m5o
myIQnhUEgSzYQ1IK8p1zuaUZrqDhSZgPg8VaCx6bxwtFErQKOK6YtSSEcNkpNrKrtcAF2yE2v484
TEbtbmnjnju1cnW3WgXPma3r4fCUWBawBpuMm9iAe786VyhoV18NOJuWqCtMDQWNWLH3vBGlQw6o
62jy7QNGLKjdWq1W+bq56JFDTwi5M8GMhU4Eo3HQoFGRW9SZPXVBxTkrmsW791IojL1dgQOa42AV
KdZrwAJZcq6eq2ze1o+971NcbSCpZWygRdkPnvqWKX95tkP54S1/8IlTs4Lpe/VtZr4yPvKcguKS
xXYz2Dx4hFv0RDzCpNYHUolilIlQ5Z7kjNOdiXqauQ2HHiDASYRHxlI7jekO9H9Xqtqi9cPllB63
VRpICqYMmGz9Vs32yBD975wgcruSVa+uY5EvmQqsEv6JhuJukRX/v+isiYWtU0YcBrpO00AWPv6p
R5a9ID1J7I3n4xoYktLJo/ROc/TEpoAZWy7KwmN0uxi9Ed74HQ1el/9OpquGiQILmHwy7yEctNv/
WXyvdNp15czWzJxivnrCMACSXxYi9UqjrhwG9QpPcV5Bfk0Nt7z6k05U7F3tWvzLwy+JlgYEquko
2VdOGjWpPfaHjejHtDj+V9GZrrr6X/o4/WQvFeTC2zM/hlGdi1PlMAG0jjMvYieuI7PqhWFnT4rk
N2JxJteE8dQ/R2pEw1zyLRLn3Bq9EbJRhDRhw+9Q3htzK/oHLHGbrbl/h7jjCWqyICcKgTZ2i40x
GmLr3reSsbE2osKEjvzAswITuQgiPa6JZ/+rXPbVitZ3fcqSo/nhmTlSwS1Akwyknrl3ORmYCEeY
xb7qTxkglMBZJhHD/8I5kUZIjVuE9OM5+v6wg3S4oLMbrm2W74aRpuNuKoIIL/Xcztz+WJqUtnV2
p2au4+Ljk072Hcw4pCFK/lsyWhs3Jgsl7yBVGFuFNuh0e5Mp6dcDHohiGac4rRp304CXO9b4uA8Z
3Moatdr5niBNXGc1cH05md/1CdKtDtu5wnur+Ku8tRpMBCIfudFawraX4DZkyJak0YoZtI6Rmllk
n9eVbjUWGg82emuFf7cw+bJ2pjF2bG67+6Ryqgv/im776bXku81Hd4+DwbQ4lVYx1mGalUoloFfb
m+50nT9gBE9/YGVi+/PWhmhS1fzbiNKiItKcXM1gxtu2niO1HvI32+hIOIcgeMMJjTaT6gVq/BkC
HQvEmamFiEeCCvMdyBMEc2ztC/XVxt/Qt4/9htaVOtwmlIVvt4xlDTg/p15ZrC4zoRcdBC9DNRJx
UuVhznV9Zp/8wJi8yaPh5rfnV1n9ImdSz9sTEtRZvdap0drVqA/Duf91SM5q3RTv9Kz01ysPxFV1
P/DMMtAFi/8rczoH9K7JfpSKfEgSU5i3jmaBPXwbVh4P0LqrLNn1cVd3R7cD/xUB8rzLALiESxt3
AtWqms472Uk/Oqxfn3L/fzwpXovUmcNwNjygLUj5i54C4aE9TB9+OcWbIDK7VV4BvFkSDFEqhHJc
h8heWSmJHgboqwfT2cTDprJigVjXT002Q8T1sr8+XFxwadgtBabwpTYk4TBYROSKYoeownG1PR3t
xzvMWtZ2SHWX6Y4D0QWGCGBHypU8Z5vBbwqXtdSMiZuR6kD0ZYFeGAoDHPewtpMPL+NSKBDC1+gc
CFVCY9GCTt7SRH3W2FQcgRaXhLaECCyLH3f/kAIoleRArC6O91UM4fQFScvzw7lWhjpXsjw3mBFd
sCqGfsJf1tMK/S9/NNNmfzVKICIAuKcyQfZchXXfIbbV56Vv2PESghgt232rP4w/yfLTeEber/Ql
rWRlJd2zbErtiEdOBgTg2UuECLnSXy6nwbsZvy8+MwnP37ypXCg+nbBPl4k1hn6KvqnZTkVPCqxA
B2AE0KaTeTFuw2bYn5Tt7qXoLaUAh2vQ+Sio7qurf2pA+3acXHmvKbA7TQmL0C8H0fSFNVJxW79R
d2tDAjsiaq21DTlmdjtin0KylB1/zWoz5UUyM4FohnWu2CRdS1v1z0ZoXXlGgk9m/tNDFOGK7hMy
CJ8r48DpWn0jLOb7BZgIK6SjdJ3BSmfHPurhWCtmmgQV3pr1en95bOaGdPjnVDFNsN/j0hLkzIr5
ytdFFZQ6kS3N8GxRiAszue75N25hU7cOatmVGJVHSAmIXNscgr5BxKCC1GD/YJmYMBGbunsyly9Z
Olsh0wFMX3zth61FcwISc9dynY/cg1KfMPhWjgMc+cnay/HOOTmfzZkf1sJCGk6blV5POmR2Z5cA
ukwxUxnU1lNW3CR4MuLD3FtQkDAOBUWB1o5uzVH5WwN58W/ROgjsiNfvW2Yu5Z4OJJxnzgrdjN2E
6lG1Z2XhWVPmHh0UWR/Rs38SCYqm6hyF5F5OKSXUdFN66xAHjOLQt03VlYfAI3e1stWEDokeahWT
2GFou2mtztSa9yP7FPPHyLSKRUWsmbFGJtnx+DZNiJTFtTjS37/1gqSlELnlhDwrpMEb2aR7DBu9
dZnNFOlLE55R2kswq2Vm7xXn3aR6ib+Q2jV5EqE//8iAwdQSuSMJKCCE+Jh+Xch9fuDMzDXsFvy2
LekDVyxaMJ17PubA/nvIAKjxrbWH0oSgwIi5zne2ABaqCoqiEjavhOcA1awZjVYiu+c1yELT84/f
8WtAM36yGL7AI2G/RwiSFTrDEYtO2Po3FNUQ5zo1bt/94CJqA4ySgmaEEgvUMMDcbG+ZDPLObG2e
dcOqePIxQiPMO7y+j9S4jvM3fHNAiDeA75YkK5J8bqBzKQXufvUaCTxyiiM8AgmJDnCVzvwL/Aoq
sb19DoEWM10EPebvRflPzNBNxXCxu/kqW7tdaxN2sdkF2qHEQbc42usewUiepIIa1TZsuVmwoLHr
1gqOnAfJEAaFGOXtFJIkEge7/90/oeE3Rb+eR/xOXfqyiHE4uWnBzsc4f876xINQyKiLvx2ZFOCj
Pmv/wabd7iYDsNQdEHKCf76GwgIM0lQX4Bo2R+yiRxV00ImC4dleFGu709SLfG0LYzQTzIRNwvZn
uWfK0lpDlNXKdMg4+nY538y6jyXlG28HkCgyl+5gAEByTnDq6iBIsY7P/xQtHxRSvGfLrm/IL/mH
6785Ltf4+9RJ87BvttjMVCDnU/yO+8vUsOjB11eKGjGPWphcf/T1jHvLSjeiWf4qiddcodjUznk6
/2jqWxoWuQFboaQgr9qKy5/F6DdgSZVyR9L9+Rpq4iMeQ3cPHPyPrbl53ZQdAVtymF/TgjDNpgOO
WS/2vgQ82x3zeq1+gNADMNCu0nngkLVVdwZEKARlp/FsY2R5sPX/K38J92/AJeUOK+ViFQvCJoEQ
Qlxh7jnfR2WIDbCOCdOQCOfV28E3QXCYfmTX3Mh8JGoo014klrcFVzstPC19tFofruIZqX/b3b6L
y9nxq7XoGoppmlc9A+Aoq+9qeaIe4XQY0byLvuXFZSKC8J0FXEm38xb3zdDQAViWZRKW5EQXMQpH
Qze6srnMIDDJzD7mFWV9Dk2SL/35Z6DBng2WcGejOBX2PPdLReKQquH1irtpNBoDW0rJI7L7EyZM
EcmaSJy9+zMsZu/CB0xPeBmjrVGBthObJeFplhP/QqSMbPsdLLtLQGoU9sSz446vBejzRlgUOYpk
BpUtubLbAo9N75QSI0P/+uddQflqoPJdj523vcjPIoBS/ez8QvDBST7L0+Ksi40jqN5b2jG3mk0w
FzX5xsyJfOLjZeCA01x04RYRNIhDFkZxIABCaO+QMlEOSRHMXagP1ZkZNGO7ku3cm+nIMGJS9em+
/0hcX1OWFhZO0L36SLcUuDToD8QRV2FMpPwYK+psVIp6njtWwaJoKgYSlLj5Bj/nzm14J3ySenIA
KXJyoaYj9pF1eh8PTHlER7ZQ5zLJiTO4eb4ZgoNds837Ki7RM/HAjjPgPwWFu/XPD7R+Id1ZeoEb
KCK/i3q7pawRJ9GNuK3p+plDqav2NDoYaSXv4XVCaPdq3yUSuThFhQWKuhljxG4qN3MGVbOl2U0u
SjUCAtQMA+97OD10CWTtH7ekEKehyEaEZV4boqNXWQz5waQsK1Bngel9icpvU+CELHjUA3b56Fo1
tJGvHXXtPYTLZ/I7NGZ9GuVV0YHwhzgR5E/snp3n26l0yOgD+S5C4GIUwgvAakdx56zIVg0XG7v7
xrrvQpnnYz2BmFdaA2fRePu2xaR/gx0ymuTuzyy/VRIfekli0sPBGQwBELEvh5KwUawAjS1E3HPW
1GcVqgMkg43YpRLt7F7pQo7QHgG3qKsJbf8RsxEc8kstpdpqYKMUjrZTNTIbif6L+TtHKG0ULD3q
Sfztz65mx4zuW99ZcaatxnJN2VtjyB5f0tKlvkytaADWRCB/oX62gc49TsF5g+EHxdfzrgEEQtvr
dUqTf5xtNaDz0HkRhASMTaDad8+bJA5Tme5bVbUQMI8hErrAOl1wssjqpZrDC36tLHfNS6K3g/qo
GNoueNekCtzoBcbjcafZLVuHLk4sq7XkvSuLpqvD4BsPgsiqaI4Kfrq6J2kw6G7jRrQoozb6+yTd
MB0NsasNULGizrZWtxJZs0pl1kts8uXgXinnQaAbL7KOCI6sIxSFTwkaB/H/79h6p56ugUaXZCLu
Sx9V9BgVRnNT/G92JaRoeEdGj90L1KV3scIi42oGot4sE1L+dYdtsH4ALcQlp/AAnUqU5VFTrgxp
L1kVO/eh3SI7vwFrMsnhNOg7IJzXunt5FZN3/gs5d+HxF4Bxe7W7pkruQpyb0qvsm6KyGIfWkzsQ
0VR3pgbe2jL5kfRjpiRG8IRrILd2zifDyRn9qGIADgP+dnYDuH/OjR2atSf8LmICuWOhtDG+UNXT
e2CwRqB52lDm5v2Vda+zr5cnaxLP9O+38ZhUd3o7lOV+CKovQ/H1itaK4Qm6KFBZZs8zwZU0d5B5
jxTAmjBaxe0AmCa+ySloD/tICRI/XDPSJwiHbfENLaHUkV/apA3xGj6sGGo1mNui7jkFUzsiUSaH
F9eWwZV87McEK/bdxXORE9tWJqvvp33rR7EQjEoGnBQcHCnUwr+3LybSi70QUpPtBscAbSmC1ezh
hlnav4BBPv/PIvturqH1DK4/LzwNBGwKTyyhUGRBETpASeIxT5xj9WKR7xQ1AvIxyiwBD5a/m+Cr
gsK5CebnwHtrkpl63/ihO+nEc5sz2txhGGnQE2GeA6t+NERjcRLBki9KULYo6do9YW3Bg0DnoRTO
CEiRa0Fg123ZNfQba80B4izwmMRyA0AXBA4l2YQr/dl3EkvqOsojrT8OYLHhhZd9TmR5lByNAJpr
843ON/voNCyoxcQ6j+rKNuszeVxT3V8jsatLgw6ySpQn3dgPYrzNFEvd2E7IG2g6908GqwWXUwpJ
z2+h7U6QsVkkoDwzWX7gS8Dhj8KhaVMQ9CjeqU4OxV+feVvnQgoKOh7Cf5MzfYmOc/chv7fDhWvk
AV2qCHJHKTVCylEg+/qqjAyxyy7KFx6/rcvsG2GJkSsEFEF8qumUTMK7LSP8qzgYGR/LqaqhqeFY
Q1WqLuDt2V1t6OhzMmP+vON3WY6EoIb6B7w44NZhysWu8nZzGXoWsGq/SZPgFHXNb/UA3O6irNRC
hOhx2E6ehoLQYk2V41WalWEZZrl7x/OeeXNsbqGHPrZfbYWzZANoCvSLpQv+L/GHrzyYFgmW7WD0
cgeahKRd/TvebH7qLCOhBFFKgWrBZ4X+GPvjXhLR/1F72I35DAR5qO8JFVrvV+4ZCdEgHwmky9t1
f2/jcOoq0nknkUcKc2lA2j7IVCE9tbxr5+gozQJcfILTyKQoNBmS2I5WsAAYfrEaBnlTy2dhWEh8
X2cib+Zl0AKz8Ud57CasfKjXMSfGhswGaqg+fGKbFVOilC31LcMjKhVMNRNNNB/PJYmP7BsrsbFB
b6gd6cAUGOwwi25e9h0RgbZUOJXqa2Rds4vFVUp5jbmq1dvxNWlNIAq/Zjsr6otLZ9LHBf19dy/M
dHkgJdA7d+7AAXBlsPBXguxBo+zj0C/dVrmezLFHMpqE0aCZELITNASy+LrUumw1z1J1J+RflIIG
b1ZgyeZUxgz4CChmhx8Bhq/xCS/qK0h8ujfgw5KRYPeJCx+4I9C9ad6fYv6PmBDwkzkjB+UDYlSC
i+3/2F4EG2XUZ/3eXdBmSKFOWAyl51Yqe7IjGvXZPwBOabqpCXaDRtFW0zC7PgQEt5sThy6dX+Le
IALgyVdNCZudGmHL9/la0eXZnFN1xSosTLV09Au3jJes8WkSeNDDc9DWtClb6rjLwIUX7K4hMmHv
PtIqLFHDOkYjX2HPfrEA/rtZHB50u+a07VhbRXRvh41/WU+nW76jNGlF2UwI0ityyDOONiOe+U5Y
A/3Au8br1CErZIvJVxK+ksU3nyc1tT1k87aOsuWAucZO2E7An3xVYOapUhUOMeLUMAsScguIpPd6
i8G9YOuW6b3ibGU0+jl97JuPH9oNahrhvnOUXjgs1GDv48Xtj9qp34mB2ZViEA9JDdjVw8VqG+iM
JCo+6OgmAPQyB/4hogoaXNZ+tDWgxSvHaNAv+8yRfIVr7j6P5g6RomgNChDEwm6f4Oft7PhsVNj1
n+ZyhBasIfB7LWjx2AH6Iy/mggiFB/FSAb4A86wfrc0N440y6VVo+hHPFqDCNz3rnB5KjiFGjnEr
tsNKVo9k4BgUjBDr/pfi8jcfruYNuKj3vfUxNC951OHMXSKvJzrVYP+rbQICzeZVPND9BcoFGm4X
9J4tdgblFLGAcjcoWHQeo2Alfm+5onI8rJgxEqffIxDzQ7tsJwGeo8Cc1z/RkMJjuQsqOuIX8Iw6
O/1S1/4+cnouTvIeTMtG2QzCd0c7bkFZsQfS8L/Wodii8tYYfX8LjLawtBZTEUYstjIQ+hkj3SoO
A2W/HfB0K+lo4mKkbBQvsesqFYQ7lOaz7MCPy9IykKf657dXIR5WffMc+meXWWkwSvzGdNLLq291
ZkqIhuqom7eGsU1SvZV1s+BNYkAvhs7uSDfAV6xOYXrK7ixEehpWdvvwEvCrfHigLqVbuZKUjA1I
k8iMrQO0tH0BFKcrQLPni7TSjj2iVp5OtLAkZR8vwabZXhZy/9ewpyPh2gPl8CB6UWv6tOt7mwxn
wmRiQQWcj9TO0Zlvdt8iKmV4/YEsk0+7mD4vJH0atFdrugG9BMhxcqFMXymhZ75kSiX/bl1pm7Ei
I6e8EJ0aYhOg/pwjZPFWKeJ6OSxbMq4uzIJUZlLSFx6YeUEZ6yXMLViUN+wmGUBGLppTj/e0HLvL
E8cFYqv9XeUoXdZhmUogbY/zo28NTw+JGa9GVPDOSigxR4yAivR2nVET5YpW1mqZv0iIVrvwCnRr
s7GaxTNyB0sKRi7Jx0ajE6RzC8o0GzY2Ruj6uIwqOfz7Zbs5Slb87TYfoYTrbAEFMotIKtrDDBU3
IR7NJ7pl4W/YoaQ8eeriA8vbBPPL2BtbxudyxDME+RaRVwZ3/V2tS6j+fLtOZElAFIi/UId1AVnL
2l20RCLA9InwHGJvehet7j4lGzKAUBCKaT0r3rOqTtE1diwDOAQf3hdNA/Xsg14A7euuggwJUXb/
a/GMIYqTds9xqjw0RQsfQNVs7R0QQJpCLP/zANOA8XSBDms702usVLQBxBmOSSnlIYd6BQZadKQe
zSOv6ivjKUV/NI10aD4A6OdSqLurB41H24Ge0lfwQ1ou/t9h6lpV77mgHBDJTXVR6DOjO6OiR+Nd
vevhmAdP1TtkhOzYmKV2kT2u5PKbKFM8XiR7DrZLYjfVrs+JPYL88Kp9LX/KBBv0S6PkBzFo4zFq
OxVIVAN2nsJlp/ptWxEoyBISK6IFRArBUH7pfcDa1NBv+x5W4/0O7iEyhz4q++T13dohvCXoyAuC
wLzYfD9KdfYPw/0R0JbYMrZsRTSHcZpErb29Jn4yGYHMbb6v0OsTqOUdrQyKsDkYqSS+9xKQd4V/
KOiROq7rz+1F+gkvcdoIkk5h90jOm93V0mujemoPBsjFwTIn4o1AACnlWWxROOUEX3XwGUcuWSzw
6HVjfalcw6FO/cdpxyqcgKv4XKzq7+nCquNqaSrYhROHv5utD79jEGOUuBf+2aVgYUPH/cl1NSPy
5118WPMQSs0/n7sOmkm/3r7A3rYYJAzqUWipUh9HrmsZgHWrIM6J7n4o8oebantDJTHvWhlq5rno
niKrUPFqw+qwAk7XsMmyHZlw0btZbJreq1Idt8FXP1kACsHWgLsoDylU7rSloPoOJdVXmg7/tiff
OzfBdJlZ358sNDUphzluKbPYHQn/V9zpzif0shjqUmImlnnvlK3CQImIMDcaBC3XpREMJaQaALPb
A5EZ7NVN2bVGsk7stAusrdwfnGi9YFM/5ISpNk1yvsUvYe+5Ht/j8nNMhdjV5m04jUHzEtl1oed3
MK3sUuCwTivWDSVzbf9tcY/bADAjoLJ9z8UhOU9CElTwr9CIOeXG/nXdgSeOMVqQQ8lUJWllxdJo
H4nNPBSJ7CLEHGIX/m4RWmdlPlA4YFrbilwrgqcX2h6tpQ54Nvv6K0yxgSyWgizzC4fESkKAeFqC
ZtzvwUN7PJQ2Dt7zHXFKIzyRtcMe2ZriBYP/07NmX6DCj99fEO4NDTA0CP8t4DowCv6RsXzb4RJb
pOjABujErITPeaSjiiTRhe8tr+iwOb0mP2isviWXoa/ONLTRtOZiO8SZx/4WwsN4Cu7V6qFrxlP2
p7PdSz3eHTPyR9akI0fRSy8KHDCaFnkmx4hUZuLr0SV0/IvGEFjgkwefqmG53THk1uW676fYNTiW
Z2eeBhzXTrbyn97JMCXaa1ECuzaqjlgdcZ/e0fBVL6nwlexyXLMAk9e2UypY5elXmwNHkWvOClWc
sUsA4wo6vvXn61i3rO5zUS15trXXw6+erHEc4Du2dgn9gy8GH9560a1YSbobSD6MlwlNkkslRyuy
x/ht5CkMkPTG/7VoJMZn7O1Jm+KnL0N7/e0fIg2jrtc8sUgwNxAxg3HZ0alUvRwwZgNmoND/yW9v
Eg743LDOQNyMxUhh3GVnkh9RCrLIkJxMj1LlD3TUKgrjpmD2Zh7gebu+6fp8O/GB7jHmijoqg/dE
bYT/xcubkk3C6nRJHNqLqxW249Je7B0igPr3lhgTvtuUIp3w88xE9/LRZIrZrYJHTHktv7JWoMrQ
xg7al51u2s67bAEu1M+y2/2X8lOxF/rK56LwOrwTuzje3XXcxMy6BGhBUaa8VWW+tFfbb2agDrAJ
EgQJErqMJkKwlDg1ienF9TCEY8y8Q9p0Eu0lwtwW/tpXV25CamYZYvu42VC9TravjF3+6bvwiDNG
IBAJkxGlo1KEmM3IhwDKGVOWGBDn078Q6X4E8w1mCF5ZvvByi6by5KLCZir6+aDJvbmm/Y6EPj5A
s/t8uAUmpEE0rMCCKYCWzeuiFU2fM1cPxiktb64Pv+qRYLqqBmX0cqRyIOxT8i/c3GPmR1291Ih8
RvXg1DTgKqBoHLu3MhXnYfyfUiIqM5rtCALKkrvjXtt0jwA5sgOxbi9+jDhL0Y/I6aF2OBj8L4pb
L6suWPl5cGaZuUWSb0ex5eT2M3Mxe0spYOeyh8G88LDLJlOu6chZObaE4NMdaymTl58YtvMgTtH0
74NxRBNXIzaJ0V3bk6dX96JEO1LNnYhfDSLhqlek5uVZ9w/n6f5cDdPXWxQ0adJbS82e7loT9L0h
RCFC4qjgUuCcvSorAKKKj+4BxNupx0yTB9KZYoHCmRupgBngYW1v7AOBV00H2y9cwJqI8rt6SDeE
5hcVrl2F3Jy0uek3oLXTEwpRUnpr9Q0pinYWvATmla1Py6QtxFbmIOmhJmw4ciCCMYwf9jgjUjyN
I0aRTFpvNf3YJVl8MOAHHazXdUp33lL6E+kCalBVQg3Lz2VzItwhjnZ9obdTK3PVkByNL8vZWIc6
K55xl/geyvj+GIKIMWDDOAwKQrwmmMh7qTaTVPvZc4tGAI46S+YyHQCf5615MhKBdC4081k3rEIP
vr89h2JOm7CEXdnrBs9G0/akVSrMi3im6EHAZUNDaHu22O2t1Ua6uTAWMjwLt7AGa0MBkciyGRcG
KYLh3sJ4EoC8MWAplU7Ia4uuzrzYUNqY4kOwSVGrjNzzSkNgQWxNyysqtauyfmmmcYA2gAUsLXXm
cYubab4QK8QEmucTZkhH21vUHtyNBN/SscfkMiKYoQk8j3LqMoYBrzlto5JsQ86yAJaB9DsgkRfD
V7lEYzuoGaZfqDxbLGyMe0Yr+31GX4njZPvpZbYkyz+rRgZLR7R+VhqbK2EKmQE3r3ymfQ4ZBIFD
qifQPJvIBvBWvy3WyNLLD8uwZg/oBY+NaxhJKOD2DAKR5ItU5HaUBof76XcWhyN/4rLjmNbf7vYI
sePIoHGvBtM7iU9BgCrQCTH5FEjrFg59EGGBAImNVjfsv0iJqrJSqn9uOqZ//Oup3+JBFd+7fetN
uX6MrkE+1SVCLfBfn4TYk96uMK/4S8tY1O08pumqoP3nwsnkEucBP9M/gZP7i0ZjkdL4sLTMkN8X
CgRXcWquudrnlgAguOsmojLl6qvpi5PRFwXFaLoYLgFaw9a8do05iQ1Khj6EiJf/Edu2UpSoSeEZ
daxoEafy1Me2lKO6VRXEsSQa6SmM3F+ZGVa7PjYxE3rCJCuM/yOvwoUIEKJUxiIgYMA2eGqkUaVG
OuO65HL3w0/zd8cRmq8AJSwotxfCaINXrZDXSLJpdL8lU3GPmxW/IfoM7gEQe+0YdHXgtrGlJMBR
geSaZznOeq/JyWGHUTugkcqMHPW0i3BS4eZqwIIjCZ7ce+oksX8eC14acgTHFCzN+mciuv18smUk
2Cg6Il5/aVOe5vgjy/ySqUiXNTLlV6br+0P9VegkIvNWzYQasf5/RvbzMftaNWOVuFthg0VbPZaO
Ao8ajOIdZESevt8aJcqsBN4nYmDV3i3ncngyz6rWaTJCmjRnRr56Xi3ElzGCcAWgqre9++HkwYB4
o1hBTNob9iOAl72yemQ+krY6CaGxZNyoTAKgquFoYiqllGNlLkP3D7CCNwhpiDR4FnFJZDX//Gdr
bIF0kr6Sr8SLtkzyyhJ97QuykWS7ZTzIPg0NfL4dnYbd5y7moi2rJY3DJJy+94B9b19/rORnM64p
Vd8zyNcn0QhlKxxfMwZGKvlwOCPTLKcWKverJfFI1tLs5FyLJBc677sTmYtse6wPr/NgefYoL6y9
HXzgj8kcd3dlTK5D39jyeABz2Tei8ANkPxD0is4BNerlanHKmcfR/odcan7C6dbhK1aR6OREUlLc
73g+NAwEPLcEYteP3dq+XGqHywH5XmarjSl0DRLtS6CpkAd/HFQLYHzaQDSuGj+mPZpCrsBS2Z0q
1BgJnGQqnL6Oo5pixrrR4Ew3XYN1mLEaiWThORfOO1IycRgi4yH18Na2wxU059mzPkKqeQVyBESR
NSXJaMMJTRDvGAu1k2Ul+ln9KtpMhqhNebcaKgszAjT0dtyr0W4jiKu+EwLv1mvH7yNqjeF+vYGu
TpQn+v2C9SnKoFXGo3oFCyjnkxigqVGBhKJkq09ZZVarF1gHAemtQ3CoW0ty6N5usWSe9R/V+/cK
X/cDm4agEvslneBI7P9t3DZDGnozscMf80djakJB8dbCKDgf3q4p1X9HMCM2kTCy3j8usvU3m3gg
2gPQCxODVJtTLvWwPxGOTHc9+/RogcmWdubW2jUDCPg5uoaQqHhbBEOw4KSD8gR6Z9lVk7NELWNX
3oD70SygRvccTu9iEqcprA/I6+7061cG1pvBfQn4Vzx1w8xFVPpscFjq/rUaRhjd81kqROOKwTJC
QZVpwCrNBZwAk8WG8E9K582et+akJhSqm9dYnQweiJ6Hg+66ay5EUFepJaHmKm6RVUz8bE6TL34I
OocwRZb8eu63xQa1TBRItfZENtpwZ7DbAgSw8Rgevx/6AP1OkaO/hZ81219vEM4DyULLgXbiGWv+
H85Be+oQSxn81mbGnvap2z3qRW8f+ogBO33lDRh/5RiT7lzkhlCsfNIzi/9vM+rdiqtLcywvnqi1
4NjZqjz5/QtjsIDemGr9FTrU/KP0t5iyIIV3wpNUkXa5is+9Sgv9/XG7iIAOtg4b4v2GC8+EI2i8
eaMFQ/oceLtKCG06hKfZvKRebpf9zzHZ0TjUNawYYlrVL6ResmTEPOFeHEL3sXVlX2mbUhHu67Ot
Tbi428TSy9S4r2wj5gLGanXAYtemcUiNCmWDOte2QunTUJmI2uFCH9494PA1/gz9IfcVucbHx4eG
bl2iZpQrWVrXhEZPoqk+OjLfHWDOaIw+tzpBY/wbGD3YpwYU86cosIvaTMu4oEeuxaSQ35iB0N4O
hzS8LQPcB8xeOf/KVkdBqbEF/3E7H3QpRCCtgM7OBgQVNncwPQQ2tsaWlowyiHeLa7YY62D97C7O
2MF6788JvjDs8eyRAG/udEevPTfGasArQIOJnUpcbcIkYBw1Kt8s/7IxcQOrE+lN+uO0HQJxh9ou
bZoQXYKmACc4Ji5Tng8rCAGVFqMibuWo8jTBMGjK2EbRagfOuExWyPWy0TD/S6dOCnUIAGkmPdI6
nzX04GmQrNnTrYl0uEuDymyP5KftyT8v7nlfLkYaky3o5MMYtx8TTuFHrm8wyZkCzSs60WLEqpGz
jEMB32F3NfoPcgXAEQunqZfqPwQro3wsFCJzsV/zk7lucttBbIYg4wNVmyjJM4pgZtxWw6frSq4j
UmmzL4xtXRRh9u+yK9l8OyraaKS/ff0sgZ3flNSwDwiqCH4Oc8UkpqADs13mlh1TRZZGY6cCdKDY
3s6pO8G3uhaq4yC78QCKirpfr/FkquNf1R1mNhDuJ5IYHpckjVOlWd8fw3P1ZTvIloU0HSoN7ofC
XLXSDjW2fgqrVYPy0IBXIYn7QNbIrSqn7cOoA7F4FXUIeAUEvxQ18rcaQeu7WiEJ5Cfy0M28o8hG
1T3qPFPSooAa2T8WX/xTH5rfGrXvESAhE1BqvwhPMrmciZWqgUXtG/YVeDokkSMpnO6o8mKrkA0q
LUwQEDajIJu1clGhK9lv+JGkfrdqZyA+rBbsi9T5SbVA+LUN4KqcK0nXsicA5O9rOlQpYUmC9pwt
X0KH3VNiQ/XwEUZddHcOZXYFnVsgXkV0GjiXT4acvkvieSFTQWV2skTAF17CJdY581G1guS5LOwJ
e9Ak9suLNJbyggc4t2AKAH0Uzcjwk2ER6/+w4YapEXbTEx1X1OdgVuVfnXGsLCO8dpnHY6oo5bv7
jki7pQkDYq9F+VIHq97HR64BGPhB68HMUVSYtcuE6hXCwMeUkw54kIdWJBKESxUgmwOPnukXzYpH
5/Uz2KncjI4jg52BUAY2ztWcFNnUshehaF1dem+RORUYo5Z/L4CCFVQIvj2lIfP5PKRQKfaL98sx
S/95/fAIypwS3Mqb62wwiAZ/AMpGW+B2+zKGVN7Avs9jljpkQblMAsev3bvUmJkK5a1YhyHpiyRw
XRPXRqv5cu4EHUZRnau2dZQp66o+4Ti0oWN4JKab2dA4jdQCUe/kNvRe8HfKmownYgNkKT1n6Ih4
XcwZC6VcmfgW0uFNguOAUqTuP4McHrJPAI8ipqT4PP6RyeWgdMx35pvUu/Dbc6BEa+fZze094bem
Lix9lFo1VpJmVscna2qEaM2UuvJpUXeCpqTkRq4T9dwXcBURnj5Obq30Lg3FAok7EHqRkk97wJJW
0MQhrIC7cuqn2xwOzoGrAgWyS24aIeqgetKwvQWM428jchk7AuOJpyLFqbWO874IJqjI1bx2pV23
d6+pzGwiOd9GoDGecApum3KdvCAnzLgRmzQKVAzMVM9Rz/PUaiRgH6nByu+EPaRIF4Y/hWAmubvW
sMGPj1aD6b1620Oetq8katd0RTDu4f+dYwOMT40Ft+Yw6EtHRMY0oo3aptlzQkmAkYIdnhrmdCgJ
rkqGoBhcHDguQ4KzaVf4OxYoHrOmrCWx5ACVBFYmRztbfDa4Say1O2NOE4m1F5c1fvRH0D641nGx
2eU8yYSklACUsqtW2Gw+f2etSon3Sj1m5aLWlWlfOrWRRevYiBfohQqIz81o71l+bZIXwPdqBlbs
GrXv6qezSplCriVJX3Rq1oFZMG7rgdrzYcdxIHJlydJ3oqKxU4rSRecGhlCEufNuqHQjeoj3ZO77
xvtKeFlvhD4xalu0aw4xTBmtLq8Z82T2BJNGDVdDfEy8GXnZdhdc5OpGpbpafIiuBQ2srUEIrjLw
CBicE75keCO1MzzuvD4141Upa9PtKhxRxzJRrlBcSYWzLCURq6CpTiWsRdFtDPli91O7xIh9wqU5
0rTfJbfVG5JYAbquUIJPgPYEId4xFQpgJu1ZYuL9zchcjuv7Un794mvILnrPHPGtPrY1ffaa4zRP
gqnWePjCFwNNXOWgsp2vg8i6g7wOD0Dq+yAiB4UzRkNh9femN9buILqzKpdsf0roEqxD5Ygnm2WT
VB0qpMwUH+auFfDcSITWebHvd5/HdDF4XEMcyAdcUzx34c0EIb7PDXPvzfVuWcHjPAliUJr8rUQZ
zFgY2OJZC4ph/hQD8OPs/sRT0oWX17STaAFHTYIM2/lNw3xtJE1mzybOSkF/5t5cCmr46WAnq+1d
siTwKdpwx4wl12o5ryn0xwGR0EI2yr4NbKkPiA+8Qo26akpfI+TiwZvc+R6uRZnDrCHnOonOOgTV
0PWfiXbbSnuhEvKitYUlpapIrqS6Ic479Fuwg+bV2cMmlhylZs1uuYjnGWUCp4PyZ9TCoaUbU2c2
vTP2Zo8JPA8gYcFoNKc100W4dTFwAOa8QD02phQWNphOCzSA2z+ayDzwYp5n3LvujFDt7X5tBHeG
mXQMa2Q8WrQyJBcfiEp2ZJ2wbCntyC2DjJzebRtImRMZCe9IVAJnnxn8/xiDwGlxxhw5zfr8XuSK
uqKG0+XBXXXqXAXWz9wYO86CmLlwwQniXOCVyQmWGW0YbtGTPE4hiIH3vXS2MUom8wbTuljJGHYB
koTlm+nafqFY5kekhROKVAqeFKBbJIOurBWja/kByYbeM7B4vCA3zhfHZhBwHVMfjeC3j9sdXZVl
aKGM2eiqKQtb4somRM2Ogm2nlN3g4tX5uMazHhCXJSXCGkiI35eAONo/ELh4OeX8w3iJcQly2aj8
LywHgCLYqvihWhPDmFCwEQk8jQ0g7s0GkvF1M7tRtMGoLWOwRYLW0hKV/h+n5kx+KqlxkYS+m2WF
LkZ2nyoIKM75a1IEXwDket9yDL35y63SrftvngPPm+Fb/bUlWIjA2TV2Xvu8fEK0xNs4aXdUz4X+
wcqqCTJ7XmuSH5AtldMn6znvHh8apBIetBU0G98Ge2NAz0iwqY43jFGEl/4+hcmoI+NAnFByE9o2
64ZLvZ7cUf0U/meb+WLWtMks0ctBzyG4Q62nYJF+eI1HpuRA1k6nZDXJ1DLdytjWgBuC2uoiRQyF
4cL8kMFRGxJPPubYAKffO3y3sKqM7LXr88/ArS/CNBVTDeLUA5n4t89fVzn1nL0+t+EM9+kGQpks
D/5VTx0UdFmuarwXvz/Ve/L5ziAohU6cAZIfjsGdN+8H5OX8jTmToXaH5HdTj62sQ8IG/im+b8gU
3dmvflIluzPgmayIlBTqazL+jIsy30UKCJPM4cldu9/xUferOYE5CuKRULWj8L45pm75O27tDIZz
kD5IGSyB/RWrrsm1ci8cVusqhOfieEg9GAInCTKvR50l4IZiU6+pJYBjsLRx4BmlezfHQwc60me4
ZHrCLgZj5caDaCm5X2hjenU7L1+xAN7smhHDxYvpTwyLpz/ZP8R01zwkF8NxNWgyGF3zIQq5Ile6
Vr376SDtrxPysi4uMHJHLnIv3pWXU7/1V9KJ780L4k540Ca4K3fR3xvBFKjGXojuJ2Zv6eFI9xIR
vozN7kAVNfDeXmMqf+uNkmg2qgYXyiqFW9rnpuT0x7bztdFpuEIgp4nyV61MIUROuAlxREsXF1dw
Fc3JeUkBq1EBM+d5EtKnFn9i5VVQY5WgNRGazdNLcUXN1UJA7fwuTbZPNJ6EZgndyfZeRtuFGKEx
OitT1KlM8UnRIgRDcRdPRQNZDdCbG6SwiDz3lxqh0VjzDolI1rxrO2etjDsCy+lBd6DJESs+7Yha
h2jURywZyaOg+6ac5xm+Ie8LLsqsy4BKqC3fU2XlbGQDUNaIpVA+kJx7MhFyi5hzW9UnftHu1bRl
TsLDMWACj+XZj+yX5jBizwTii0hpzjEvGKXKr9q6GiPcBfwqzH7/rqmkiF0Fgtsh1lbfxNFjHs4t
BzGoHeVNROoFDUtcRNA5aUVeNSVv07a+ABbXj5JU7036w47NnfQNU1bgmmeejfZdK2Z3XwChffCW
au6n1+wxrgBUUUM9ULOmXLl768QVAdifttIqG5lvL8IbEL0xmAFMrhS5g6gJ898B9NdeKloGlryQ
TUcLxAXhV3sofSaFDFDw14da3A4Bagyb7wtjwwXs4bkzev+DvycJk0IjGTtOewOjY7ebqyvcQdKN
NVhc7Ll7kOEjyytMm0Lxya5uW7/R/Kj39et+oCNqDVGLnOyhX+oDzv/5uNPt2/YuZiw8Oue98wKI
JjSWsdIdAaoMaMYDtW0lDoNG/Ps5KE5y5b4RdRzmtmMJKuYjjt1cAeKFhb1j2TOtFYfk6nFtW4Gf
/jy3S69VkmNCO8avS1oxk8BvQRnv76Z49zsiQ1qkbYdqPhaPHJ2zeERGupqJ3+MILuKFFRDXymqy
0vBPCcE41zr8SKGR3XIa7xKS+Jt4ds5PmaBQUJCImFoVLJQzKWmZ/NyfqlcIyLcOKxCtwRjdMM0q
ft+fO7miqE63CLCXVI2fsfqO7Wa7iz5j/ir9tAx8MLRyW67CQl3kTHBmGUIwLRVB7N+H7MiQFPqf
qh5K6xOmUkDWizUMd50O+A+EUJmnUebg4WagDx6V7dLUzglZkwbQ35gdHO1zWWXgemmoGq/5Ihs/
ZDxRtVJhuSld2N7cMCoENt1f/MwkkcZem0s2uLop5MgUXC0+1tZiPDyf0FcTXXBvSlznnnK/Rnxd
luEMUcX540JLjYTolwBaUlOadpeHdasKxWZMhlzcIoza3mc83gsy4FP72i07BhI7xHFhHo5xYBdS
tdElBkheSHDYC3x+Bm6E+nUU6YhfawOA+IprHXJJQs6cbeqbzTNpC8Y0ugELdw/n3/BSlelK9NuT
YkOxltdV9oYm/q63MUsYIZOATApGXjob4VyFH2Eb0Waoc2fiE6hBFnDmOjJVJG9FVebBW02s6VB0
vvL/21NeQH8ziQCq1OVIi3SMxqxCXE3gOe3fFGXIAzNRh9bxC0TDJ3wnoW8csXxrqNY4ClLsgXk0
dQvjHFNN0ZzMZFFEv57zKpDzmIsxkgEAuQoQS8uI8F43lIylY39ktngxBlHlWuC/4WVS8DNZKCb4
O8WRSK8pXsIZMmMmduUE1y8816+7teXX1PXq9RwM2RnFzghaLm5G7OUIuKa6pDvKTsOlA46izaX2
wwkdqSp8ffQbOfBnOJsfQwPeAEW2/7+yiRDzbN8tqetx9k6SIa6DUzXTIGod+qxQtA5MqWRQYz3o
7HowekL6NgzPyD8Eadz16rdGacp9tjOYuXBeetp7lHTbj8rpQUPkgubXaRK8c05YmjILKhRc1ozR
SRjNZviiJSkSadULpPO6lBjNYfxvcbU9admGOPZ4jDPgro/wNMIYYyxqzUk9iD/AQYnYeqxSyNrT
ZNTfY210buC2n7kN9z0kKGVG248UnzucCPPG+hJeaalPjbM4RGVInhNxewFtC7LImnlufsnJ6VUw
ihjzAvw3nbhUYI5XXJK7yOW9SjpkjZRpTRNvwfePv9RnHkxKBsLeO+U3Xsopmso+2wI67ujd77bc
KnUp0Rh/l7gYRKGBchkyjAWaA/i331HCBEDQyv+S8RHeVIVjORxW8Ny8RRdbe4CL82cb7/AJ+S3G
creLMtp5c5q+hYqb+1Q571AyOvKD3fED6uNkQasACnoyLdlZUlJUtaLKUIO9/DK302r/opBpNEc9
lwCDeCXA/euGhQUSdKZM9qSpZs6RyxOMId+cLZ6ru0+0P70QM3hiT7mp4IP8PGFVjsUI0CVTyc4Y
lLVdGMGgSPRWjR4SuGqIHQ8qUm1paFldR8Yzqt8R20yt6kXKSPPqmlMt1jubeqvV7WLqClAa1TBV
nuQvXojZT62NNdV9rMUt3bR4AklBkm/ahVidUl1ixSpzzxUHjtwvKSkJvX3+bmHFwfKXMbt1j5tO
IPoB6dssHXckafon8mcd13RdOwcST+gjGaT8xXNNJofKgwdx6Kfh0abH3w7PBNjGaDckBnD8NKkj
VyzyZNfRnXXnjv62N9I6Tzgk3oLLbBCdQqLYRo+aNUo0OX/8DI7bgwmC3e5yKQElSOZqCqQDk4Q7
ZuTIB/dszGmLg75FOSLPEeHz2RzboVzlfmI2a9UVyJ0XBcpanbFch9irDov4xPBzOjfeV87XOVps
421Br8xdLXiKsHPuh4naE5WFV7iFpzU+CYMbw7vSKCByspAG51jyUoxUDUfRIxU8OqNKzeP7lkUK
G3isjrgA9nJD+7/5N/YSejIJjzQdtHN4gS6ECjpEvYQk5B5hc7zxj+B3NUdcsBNW+L27Px9YhYDE
ziRopjE1NDaHTcyPV1f8kM8NE6kTKHVk4Aadz/954u8Qkd0z+fcQknGkXjg2GGzWBr26fduNyBrn
HZ+6CO1y2q7mPPTUoFOOjFr3gF7gvB+Se59329zPiKXcf0I6g4MalfDozQpGVir1/UJ3cBCK6eeV
6LQK0RncYulX2qp0yB8Kx49Xjg+Z5GB8BFr0k/1ujVp6arxI34RXxPaqtHk/WDz9gdoUedy/5f2+
xqxdLF0XXRjtnw7hbA58gAiCWezt48gH8TNW9c+xt8cubSTENMvIiJ0NCGAM/d/i2Jtb7rsUnkYu
6KvkeK5gIeia0QhayC0vZgcy73xXLoAqvN5juQKo9pV3P75xPzxxcLOp3RxKqa+ty22mjY+IC+Qi
OXIaVR9wfCTxwhEMJyrPqWno/UJImA6upiRC59IVSLrYbggVknLE86daSH9pwBpbQ+dEt7cseVRI
YEazV8TzZIOsnzQg39K7PdKaXUJ+jUqiECChOUj6t5eMSqJ+O7IaACjxnV04p7/ZHO+3fEExUoty
RgOBheykFj2DHAcnW6kIKadMg8I1fY6ryqXhZTSqVidQY/Hpt886e7E0RYK5IFcSg3rVHvbi6bZT
IhVIDM4WhWMadYIi4eiNJt8EYp5EHikLDvAJ61ReaSsmCoCiSPZLOinLYEqDi6cF6KTSylWygU5c
eXOQc1xC3Uo4HEgPfyLJWFVjurVjJcZe4A5RWq3p7F6IFJNV7r1MbmRF+cHWle/YvmTGyC8G0Tig
i/EduM4bF0e4oAqRAQDiMuLCXiS2lH4Aw7+XXoUaDZw55lMYHGsUsePfcCrGedrGm86Jz1YhzjsQ
MMPAcfhV06rw4l7cJhcu2GgPvlXDTg1ghdQ2NBxFpcVn3TXDHllXhKx+j4A89n1+kA6HMffV+DvO
Asy387o2oHkuBLPxISwgW/7Di+TG0jyXbnnPiKeIbFxzT8Kbaq5mTqgtC1H1HAihzFLbtIsHDAuo
835h1SddYuWKuuI//MLQ1Wqrl0wH7nbzXOg6IIgYbPgS8S2qvFFei7msDSORIxD8XATbVKHUPI0V
u4PS0Lq4TPT/+dXJtysB1G7McRN3tVIWoL5VrikZGBXjKwK27ZGIklohTyb13u94k4/oXl59/SF6
grdJRRxk08QBkxSby38X3mt3ozIfT3Kiotf5fWyHt773JheQrf/1vQMMzWcSCs3qoZyYVBOia5Pj
sOGkmgaYVMrqn5k/WccLbjPDsleMpC/gvI/6uFzZrAqauO1vipQIu4zSdAEZyFB/bR/fdgeNKMCu
H/aCdBfdn+C5pTCD0qPvCpbdI2/7SisW3UFX/kcU13sjFSHglYkGeiyMo0z7GzsKv9Bl6yJSWHfl
s+h8qtk4kRv3jouHFgA7HrrmhnxWXYvXZT0qn8qpeRsLrmrRV7vJt0kAyFka/UyhIMWyoTjGn1Gd
F3O1YbmOq+IBKhRVGtNFfizeivALHRrhklmN5IX/OBj8Gs74Q3vDYCyTTo69jNXsdWJ0umu5DYVj
wvdzGFTVAs5njLpf/ghlK6HCJ5MnCI+ZCvwbB6Z+eU4HlnGOSwMoLTXwnWPYEGgZYlo/f3mFN2ps
uFd/8OX8oVcgOvMG9qO7ECqlXJVolH/4F//kKy1x6hqGpm8ZtOZrHnP6vJwOJQrNAeCm25QPwOaq
NbQ/Pe4QcFBx4rTMdRRWXkCG3wbRTBCbIMi6L9dVPEw56DMbbxGTSFOlwfFg3rJZtd2i72OSt2ux
xrfGmiIFZprChFlnMXbdgZcQTNOZpRFZf/iWWxgc9by7f9wdGquVoHkqTszx2W8HV5dq5bSuVVpR
y/aCsyHACZEMWcmp6lAiDZSiLcs/jVp++G4Qi9r1J57Vfb/nSgFkR9++zJ/UpEUccPqquLoM515c
WfMRZnuYKDSp5Vrtyop/a9sm6R4wAD4wNe2W35Mz0+lYdqQQbQCw6R2k8O437s5CTiRl/docYdv6
Ea2FSxwspAo8Wo3I4uratm2dhkSN8LJ52X8HajebV1QcT1NgY1m0qjJMbZVlr7p2Wbo+g/5t0Af9
KCL0X+Oxb+MG2+0tbhOqiAuyMACtHatKpV1VAPmw4f4wZwcKIOewZ+SvjBdnuoo63VSvdAoUokN7
vrWN6MfQiVctMXEbU5GhTK9egzL+JKeaU2SYbrXo1hdo7jMQS5dg0GjJP5pG44ssSSgQe2rM3jLX
a7GPl3XM7haiHfXRM2ZNoyXNiWzqI4JDkuXhn61YJ4CCo+w1XkntIuZhmkTQAEsHtuifbbZKkBU0
xieBCgqviBUDWc08fjW2aEXmovCay+5YOoez0rLRCJjVXIAxsVC8QgGRxw+m0+N9rdP440ptoYm9
/SctAM3PR0bn7Dx81Gh8pq0N7ZSbxZK4A+KSY9iOxyCtDCIUhTfMR4DWU51DG19QsYNhGgjNA3y1
eyP14gIOgHwRBjQDQajtHtBvzaYYFWY3eyQAW9pVuUchMlaiJRliqAHoOEg/4TFuYAzfWCzI4VXJ
fUKxKdvUZH8gFnbjA2AUd7Bfg2FHaQQjPV+oA7p+CgVfwqykCBnn61zg7BTmGXXAktzoFHNCk4ma
aYyFQOUp8ifzjhRJm/aYgj2HNVa6NGOnEsCIzXG+iWeGkCK0GZEGcdkvxOGVRX+n9wXV8jtJbP4A
q0JKMPMmQxI47ZxtWHnQ1YpUsQTkU2KMdnWFCdSu10QDI1DfZ3D8cZcWWYKYHJp43mglcfa4nejD
HA5SX1di4nt2vnDCHwTfDEfPv89wrif24DPwXFvVsvZ3fVO6db2R8vPir5VQchq/Ui3xCR216BLr
HHI/5YBIiUManhN4f3eHExGjQAgny5WitgHt3ANQUzZpku7gyAfuQCxlFeCKI8UlGxG8hxcskwhg
6q3BGNU7zWIBigStadOmc8NFTn9EniwYtJvP9XyuU9+zeOe4O5kvs2mEflzAZ7vyoT8EWDDP2+0Q
Q2QSDpxhiXNOp+AC5QPcP47ckBiyWRbYgUVfUPoRsM3NVasee1NqajYmJhwSgeaMuhb/EEbkFLgC
jooa3sqTb+PbxYqoZ39A72Z2rX82s4VMktvkQPTvGY+OJZOOaECXXWFcWomh+2MtJEeXIPNsyGFq
/0nsFo/oBKbrAdI8is61bmmOj5pj3+8WJS5GsNDbTXnIGoNt5cVU4dQ2DCpitBMPeiHgZQ0rDAD4
OypjM3pHw3/rU5OIcPemEbiul6sg72NSUc1p2Mu01B843r06cVDbmQ/PDM9B8Hi3am5tqBoG4MjC
792tR+x0IE6Eg5DAGimF9Ri4dEHK6kD1afQUA6xozqU/ZW/y4RStGmJ+9pBFAbg90dCbFIi6Zd8U
QJ4Gxb4+abFNJYcu6fYUB5YlNZF1R2I+7SmPz46BrFXg9P+QsgUK+TJX9Z7+wh6rPK3bxOzlCiom
cOt7ja/jaOMwDkgiB/HhNP9TeTNCPfmSFpAC/Idy+luVuydUK4dVfkS5A4FNF7hCWZJzRCRfpWO1
+l758RkqX46W1Vot2QoikoyaRyZhKD924WaxpzCnWYaBNrV28QSMBBqFRisOqKjZQqdhMthwmXYA
+6jmVF/7Mh+LGR73+78oz5r5SduEm9uQ5KSxZaUXHdTzJbl1Z/dSvvJKZUe9o6HZ3I4+kchDo3fG
iMNgGtXlnPwowY/pj/+Vb25AkeNTomu8PrWuNm/mDtUvCqb+uImCSeJAZrzPBnxJaBuAx8IM/bGs
z8yP+jPcVfWJlvbsHQrabE5tRGNEPDPjzDsjpQynbwO9WjeNrlz/Dpi1lIMuEllHFFQELcS3d/lp
Nh9Zaj6UUUALnzAA7lmqyyq9pxRBWm1alxEQ1Ur2lrWqG7C1SmaRbqn3+SYbUbU8h4d8ymjyDf5k
Kz8Hz8GQoT3JeH9mxKZnQnSM5ar8rG1bJpSNuGEYLvnxcAgX1sKS0Nf+VX2nFheCd84lD8Nv1Y/K
5WkUHpsY/rRJO/SLEne2xiFoxOhndvZYcbPsR4K5+gQH84I1EZmeDmHR8fUsa+CchfGkcy7t09Aa
jIhQ5ulXDAUbGzxEdT4RzCjyb40pJ0uZkXiVTFkO9yi5K6y4TFrdkL1mg1jZVmU9w5wLzvSDDk03
iWuqFVM5MAoV2DSCj0U8xSYOkxwl+Ny9ru7NlVh3EEUDQa2taqootWEsXchcLmqpBAwWdRusocnW
xv9/EkTSJ4qBPxvFunITx6JDJKDUx7o/gr+gs7/k6otSIJUznyUNVpUchxWIj1jzCZJYPqwTauIB
kYkRrBFIcMLfj5edINuyBx4qEO75t7mXlfCs4bHomTNE6tQn6pingRFz08KXkxqrou4Hap4kFr/z
hu+wZ5tRUg/GShrCvZBD4pTq0Y4QcWLkKLecoDLE4Cxt2Bgu8VKVURF/AQQw+wD3Ib+4m/wNg+hP
xHbSyoXPbjIJ0Y9nd2cQS9Nlg7HVBRFHJp6AhhPcgDl0s8GO5qCLryIBzkVW5eqVBEfOY17r7ArI
e47j7cZ5fN0jhgfpTb83F1xSeauNvsc8wpLFcpBGcJq0nziP41qS9IfiEQqXrqNS2y8zta3R+r53
1+baU6ElbG6choreeOUWMAaLxfz/2PMHxX3PDL/zZjbF/sFh24fEuWqX6IKfQ4RapmYd+2mjZZh1
4z9ohPpTkr7dON9kM48P2qMGqxvW5+hEE14/Ogt9ejeip8D9E0AasHT5e4hBcjBv0UPmnDsrkzNV
73YIJjd5eT/FNlY1Zn3OgNYW3O8m721VwhZVIhXxvd2etpzfN+62heT3A60oQ/57CETmeyVvhgUQ
vGCQMaXfLOKHJ/1xfRDA5A0f/t7DBO34bVRYu18Oq2DUPAzw90l0tl9HHQOtfa05S+b2XSGi8mY1
06MXFyQTkhuymsg9zjzv7MEF3pEyVpYmnaCIojtr/91Ug+x8GSE+F3xFX1yf2DVMIT6Xe4+SY9Zx
8QVvwm0n7iI7ykhQPUlPkh0fKnaTXnAgW2v/b9Vh5wsDBY7/2xtmmA/upjDZMgigF9iRM8qAGRnA
DD9JQz2MVmzfnCya3mwF/wWhJmZqTKh7Fu3Q+dgPpdPAfKUv75RE1N+GESefpZvbWZY1IelycWRQ
ilTcH6lqVieVWNA/yXrdsqbqEfYCRI3IqIXHXL0iYcGx6tUK37HqJvx2JFg5GN52qsYaHXvV/Sxh
Brp+PD5YVO56GePIWU3XLRIhs/lCHdgmdmq1UnAqPYLLM5ObS8PE5pRc6IWXssw/YMdUbe8n5/o7
pSOIMAbSwyotFuEabBORrrNRuThvyK+AvjCfOR4HX5qD9aVGdQx9fjO0F4j+qSa3ZM16of1RTZIn
sIYrom+halSTIfV2dDQoQYB1hN9IWyTY904YTfURjW/VQ2Gfdl/bi/7fhepCSFWmsRuhURriTlBc
AjTWfDRV4g9MFVV6Zc4xFnUsEPDUUSERBFpdv5grjvzCYLZBKs42hWxy0CesgoQRB2uESoMrOzpN
9yGUpjP55dc7oY6pMWHSiBRUCSdAknP8nIo7n8I2wbmx/VLBF3jEJTop/3mPMHHP8BreLrzqmf+m
eDUf7z7nGwyY5HB/Reya66lvR0V05SRsdln0MX7H7HCxCbRapAgtqd5fA96wmnejJFsrZd4aJ1Y9
9CwHEB7mFQAlrw6NS6K0DaIcdPF0AFncCgw6PO+tCt8XrQD33c3WJcCvRaYLuxfgPCbK2tDuC0rF
JiLdBNmC0w5f2271paoztWR6PtLMm6Fg2bVM7G3Z9rFDzI/99RXBUSJ/KVixQ/osQNdhgvO0z4MV
FYZvtY6eV4/n0GBML0o0rkuDdQBKA3KvwALk0Hw6fUwo0AH1D2yeO6vAAL1z2QdXcaiCbxC602ns
glj2yH5e06ftCDGLT2iyIvbTTP7GUi8lFXkcJpsrArnVLv93K11vQJzM5kvJnDMYNQQCuU4gYtgY
YSWatg86KvbGrbwvTZv48DVSo3A/MoRItU/v54lOMZxCsYPLiDDJABUXPRdDFZZndB6SchbPsgwo
E459T/3/2PlSm3htqoGNI1Ap84Hiv7Lx2p+VtaI4UgSWVwub0i1/7ZiKzchPhUNH6QJBQuF9GPvH
xXpHSzBeHGiUUEP5XmX93FfYlVT57GdMX57Lw1Fz0wM0HUAyBIH6BXcJhBDK3hTrA6BS39GiDzuE
/wDdOsMGQPfbxGumZ2eKbj4s0C4kgk6gWYdB7C/I32Xqyn7faC9/eFfLZpd2Om1/sB5CP10+3Owa
C88tWpl4Qs3Mj4WB3sNOyOtzf6HPMF+voY3riL2sP8tKhPvKHDEvm6sd/m4IyxSHlaA+sQKtP/sP
Ht062McpLRzA3dPlVKt1tfwnQnQmQ7beiibApRc7iWMgWdc8YgD8etbWJTvqWcQg2iU/sVk8nF1v
sDcHKAOLWKXXbd4l7Xzi7zH5x3C4pmBt1vAxF2P7xQR/E4mtKXt+7SAok9wOT1pKWoDWSuu0xPUl
neFqH1N27iRLQUlylNeZCZ4LEXZDK9xRxUouRo1XgH44NEEKihlr2By3RfHD1rdSrdairOcYHBDN
tNyqpabvTvIKkCIxiMHGhJFFqGv51Enz0+XO2O+dyeTaXm0TZN/8rBB3e6ru1lS5lYfC3s4sINfR
OHQ2lfnEHU7WwVq0Vx21UpOYccAnc9SBalG16DE+Am32HE5/dvPF90LPyWhOTHTQfHVEEkChzDFz
pYUyImIT8j/EvCV+/O7acZtTSzl7H6MkrTl7Sld69LqGxmEXoMeGdBfmo/BznWG03wGiZ2lc7DkS
y2z+ZvMuU8dnzmSSd6SgIi5p0fooqg5+iL1kqSmbdoYu0+JUGz4Cv5T38CfCnrhuzn/idXzxMNBr
D/4M3IBhLv32xSiDmdc5dzdp0KkO0qHEqC0iYxT1T/GY+TFW3vcDti1lv8/1HswrVoqm7Lx2LE3l
7xCdKY7KaZ49KGw5Kq569CNUIcc2Rj6FWjfg5TbXYw0tXGft/tavRVzvMjlJniqBUKStV3Ny5Db5
SDA8y9FgW6MGSO8IcBJidans3F2Jh3O8lPCLgLMJoTcTNJKzpI1wTyIhPhb4P+8xBpbbHV+3t/Ia
iuOBBAMmkVnBi8CN7QUF1/35LJnOB/UVEdYG4S2GUO9TT8Wn/kjI3dgGYKi5YxWOm/9HNB0FHRmz
rnldDGcPwPBcRIwhN/fNaX718B/WuTnb+EanoR2/y4MwLsT2WkDUnoYcUk+Diu35FpkLxspwx7mn
HxHTPP5oonBi4nzCjnXxnQfyTHTKSGYN8wxOu66uPXRxf7CoLdI5kIU8NdTyWz4kFJKLKD1cupv/
L0XAMRuVcxmSXTLr1NCwu1kZX5Ic4LkW956IuHverjYhtp2LIPy+tXtyO4VXy4qw9Yr0+OdpQwq6
T++ZDfvNM1NDJv7Pjaa0DTVd9iMRiso2srsjpF5Yfpzpg3KlTs+aqL4kns9vHpYOgLpe+YYX52OQ
XvZX+ouIzfY0byQBT8ORaDZSJZ+877NP3Em5scy272w+Cm6eWoYxYFN9X7jDuUUOvV0s4DjyLSwW
mwYDljkN7Nwftsqx5jSYvYpWORnl4bDt6tLfvRu0w8FAon+UjcEkivEcYNl7P4xMuYnu6Plgef2+
wuStJ57ppur6I6jyebNk78eUkSGbyP9TqXNdkje3Allzh+5WdHtAK2t89msYNj/yJHFOnvwwmSF3
VtJfQyuO/kkat3yzq5VtDzFBfXUY1DvTMlws1iNImHn/BnWIJa6W3l487IUQyAC04lH3r8OPKbKq
m3h8LyHvYft3BwJZBmuGzrHIL/fMOGGqzKitFvx+to14xeZnYYA1Toa0cmLfx/VLrOhgnzNM9qug
wIo+CjJc0RxE8W44EiFVkbyIe1vmB4bt2LK+uOg9HWgvGXbgcaOEjC5A5g45EVShCcwU5eQGLlZz
gqE3qJO87qV8YYraGQstvHam9ygegUIwhPZ7De89G31uFgfOnWjjNonZDd07JDZLrQSsVT/wh0ff
jM7gOukZbSxys4WMPeWGm0eS71c5ZnX12c28/1ctGPAKEJD73c5AR8asOQyNvCrpeqDJj8lQ4mCY
4GTbITogB4JusY2TAmGcpYpNY3S0fDaTnbYlmpWCVMX/T6xkdkcpv4yK6qEB3AppH12HFFE4P1Ok
enID68xp41Q+4Z3ugN0TaW06l3cbp8pGhu85bPiz769YAQAkN7BhPooC4qO8lKCuubt5WuiCnzNk
521m1Bwf2lcXoKpgCujYsp+WZ/xpqUIfXwdCcfjel6XWXLRdk2crSuy3Kt4pFHmjF285AEBOLO9j
OSsRnpS2WvQjnF8sehCirHlGELduKtFdcRLbDFCu83pnKImQX21DCjTJnHdpXib+XpXJN5U7xy+4
3VqkEZ4edALoSSs7DPm+/NUzaJepTJrlpHDU7RSmePmPjRhUzi7WsgKe35IJNK/SfG66ne8Sqs/t
x+BESiN/15SyNZmucLeaV6vFAAIB4JPJCSWWg14XF2AMYHH07TDP0jI3t8GotLDVTzFsnu1WNIGQ
itH3CXKlxkBEwiKqIfsOksjA4SXTpilc9RJC9HLLfgaXBzWcAdaep7xqH8UHVY0VXWLX0zjt6amu
+B/7VrbqP/AmG52R6iTQor+KycHl/qos79Sctw+bLxbxQZmrs6wyqbc3BU3zcCILsIxOD8MPwbUP
fzvuSpQyHvezBV32nb3eM/yDK8oOId4Qy85lrG/pruJeZhqCqNPeclS8hUkXdu/nRjj0lJ2nTo4l
RiNON/26NCo8w8A0yvk5ZmBwkEfhaaskThL9STeWOLnEYRL4K4gJ/Gx5l/gTHeFmqG98rZXfJOo7
xMEC76ThQ1FqgVOg518qvQYC+xh3I64jp4jF5Pa7+M6ocGHN7ItF7wB14YgoDwjhlsAQNEXTbL+i
DQ18R99k59zFkVjAcBViEx0AgtUBqw0CHqsfynwjswL80N4bv+68yGRZ1z/7EIvgSTt77pEmC5/d
f4BIJu4gP846CxTYyH0o5XdMf+GsfA4HFTkkcTGxtbVcNZXQJ9WM9LH+kmYgQ8T8Mpng8M2e5uyk
/2AHSrJLmwUje8ZKJm5PhrrRcM29WFIbc95FCzzTy6dBx2C4VPOYkcXO3pmZDqHT9uem511LoCW8
4eZO5VBmPM06JDyCddnqsSOL3o8sgxoYJNGEgrJpYqH1b+ZLgrSbxhGdqxoXMF6ut1uFroz8Pa3Q
Cn54pS3QeaZQ4hX8QBlIeQN4bTGqVWqFkg7GLKcoD47oocDq8sFKoJBBHe68OfPgzFulyNnjgcmq
qA0anxhP65TXOZWO5YR8z1EKoCeucaMmBozPZm/YtxsfWZozP/W/trsJupiWfwnqOEt6VvXLtmL/
UxBL5p0qduL8q1OOUfnxRKzSqsN7n4uR4ES05sXa026wHIcuSIU/ZM2cM2tz/UZkMcEu+oKmVwZW
nmk9foYDzHU1OoWuwAoQiECk9sgMxFIacb2nBrmiG3k2lkHrHMKhAcUUOGukHvMtYTQJLZVwGJmj
0nSR2cvj3nI5JhpWDTqrGO+it/YLegBBGomJse5zjVFbhVlZ1OmZoNh3ujJoMUquT1SpyMuIkiQV
6DuDhAbsUtqAL3yNJr2hvS9iEnRGO2UgCh8O7FKVnClsZ1LuEyQBb57s2x8COvTvF+3+/H+Zibh6
HZM5jVAQJOcur/QdvFuAhW/1/iJtCHRXpQXeH9uiVjXS+5YHP9bMCp6gxIrB8TG3We4oVbp/OUYl
j+ZvDaGs8K6izNzQO1krJ3WZoiTT9JOjDEOsnzo0SZpRP6pP9p1qKQ3h+BNaqTFc9WJm/e01TJ6k
brgeFzt5E4QAFgMj02hWN8U5Fp2MVjrYFBRr6T7IHqdRnIDbgKQIj9dkLSiykbgVm3paATynmHRq
HBoiUIXviinveajKCZ6VutHAkizkP6nag2meITCMhcNLal0YZgp3yZsao9MW7oAO5uF+F78LZn25
mCd/ntDbVlUZcLZNP0qqNQHXdQcGpJTnQkqW3FNRc9JQKWN6d9tQA8UbazdaeuflP8ntN8PmTEdU
H3flqmMzGoYqhWz8TNahoX9BPaUvPOeHuRJl9bYVGBejn+5EyDsYVKVR1FGE598ZScepsDfDASU5
Rg7mojNzPPYIBYML7wnAo4pI3SeESd8muS+YCuG4cSYGtH1lJkTyK3PXe3IxBuJG1yXP9a9kKto1
LCTf4FoDCJb4kKPXYcSPEov4qmEA0FlQnwFB8XbzCzTPsBjcqT5vfgnA9kNk+wDKeBxbzicJ/KDb
F8zqfrqRrLp0jkNGmfHbX6L9jH1ESlP1v914JIO26xchPdzgQgfbQBnxgObFh+cm1E2jRrcB5f3k
BOfYbzDCm4BDZfWIR4EQ5cdh+wAbr91vtiVvtnJNMBsz+6P9ZEsBrjUpbA+7Z0HVoy8yrGMH4uM8
Y/qFuc3pQY8hIjYbBtHGiGRMnGnSaQumVgc0dk8YX9JWBuW286SGg3geMbGpnBSPTkeOXy5tkY1z
zUYQWe0pmDgICvnRs8+60MQ8Sll7QgC6xEE+ll6wNczhb7Wpg79hhIKYgKOapxEytnnMqSjqvCBu
HBjKD8+pLTENF9meNJWpgGPMRzsKjnMJQHz4oZgn1SmOfXnXyRdIcTq+6XMo9etkmQp8WQQnIPAq
BJvA0VNH0akbf7DtuV1W+1i99VEDNjtv8nfPjyNxdCwBERI/nHPUviZI2fHfKiGYDUHFbHKXniet
mqlgrUzgbp5porzXaLLxQnF6XcZhcj3cm9k5y/P8EltD3kZ0u/cVZzBDv4UtAEh3ed3caxgW3iOT
zW7HB6hCu2O3xSL+4YaM2dk/SWrnJxq6+hBBFQKsGY5ClNvhxjIJW5yBzrLbTVnR2zQpSLI2Vq2D
AgZE9JADqd4qS3P4csrgIJA443Vb8xgZ9hrzyxYW4hZwfaE5BXH2Miu/YNpVfHZACnzVbZCHOM/8
A1kE80lKkTuCXz/vN4g+fm6hFLCkaNjbxp4cWpp1M9y3Kh+6q0EG98A1953THJ2qz6hv8qRFEMlA
1JOdj5pbxz5CT7VJcGaeA+teOBnnkhKCmNbUdSIYfsnCnQB16IYspCeeSCR4LJAsC9A/AjFehEd7
spLTytgQA+vUFu2/GlN0AADTVP/JqhQx6SQ+e+1ujlG5JFI5NeGNawbcpGNSUoBhg8wIfar1Upfj
vJif5DeuT845nKUcNj/oIGVpS2caqDubAfbP7zrwklT0zNGd2TSRYk0VHApSxUNlyBtZAZb+TDyX
vU2VmpCxu/23rwkb/t+aUNSqYG6siit83zxHPtTs0L1VyB3x9PH59/qumlNP1IL0AiPVz0+Z5yTi
rILk9QFpK07VXXghvheCfReMaBlAOK553oTjdj2CSQJf4VNc6B8f7fEWwCl7WvToet1ih5tOM09K
tNg1Dpr0w3XyRxhwRD32pApYsqp+X7RspiYHH6Nnw5P3iYEqRlo6ql8yGnaD/mV1HL/RZAHWp8cS
9Z98bA8lUnydf4syiYSWoQSPPGcRqPRdmCMGgTlHELEcg7YnH0EKWWZfhGPWh8XTLRSkh9AQguvx
WLggbhD1sVISR+O7+lWgb5XvC2USR5eyQt899k5Txu2BLb6ra5JJlmkHhGG0PhhAxlvp8ECXR0av
PcEJKmILtbD7t/IKyDa+2lnTCF74zVkeK7T/FyS2BsIrQoY6UHcfXqmcTz1Uk33KGrM37XioxOt6
aXsjMJExokeYWIP7kHXOx+VpV9uG4go48vlk3Hc5U0mcVBW8sMDqaJR4a1JReiMObQlhGvLhExOh
ldyFvuEbOlAJzHyfeuRP3Jaw1mwe6A5pPcSSeVdtYIcOIBCpx7q703AaRAVgGs6M4SDv+nf+woAW
GTQyESENaZ1/dNT2uZrp3JXTGHYCJr1N8Bo7zKP+DI01c75aYsEte+ULtHj2fHBIexicUfle6u5y
B9mkCXyK6xyGDjzX+VfaD9DxPbFgExKUnLFLixO7W8x0HmfgED6d0CcjBOrBSq+yL2yyTnPqlErP
6bGRUfRIY/7Cr6Q9szHt4MyA2VW6I+wXFRQL4HX+a0SgP9DvpIv/Ggbfx4bKaTB/XcIeyIb2kPaT
Sd+FDPEEPUw14yIGuyo0i4bVFDuJuq1gT97fhYEpyac9IDtE4bReTZ38Ufw4qAonmZNfyfpVYC45
PdZjKO0AblmiN7e9ZAeSnPcn3w+u23rJdt3/vBOMBn944pRZoDS/Lm/Ka0aP7cDqZzBv/ZHMdB/G
leJkFmdQGsX0U1HiNjDgS8JeWcgxS0wWLWfe4Uws9/oLQ1kBHfKrl8QsP/vJ50q6u03GYcgdSkpB
Nq5//zikO1V4cuRm8vR1bmqx/inNA/gWeiOpzBKQqfTgTbJpOsIMT0kZK+w1yt4FbUD0PU8HAx4Q
VvMKkEe6aLrTlg0E1fbDyfyTCgWye7qchtWUfYmYL+pI0BJwRj4OyC7dl71aJl6I7Wr3VnCQb5Xl
9GwSa0rhfgJ/n6RaNTSR/1vb0ig1iiuxQFemgBUviIeMr1H4zWWo23JiqUyfnobAYA0eDptPNJMF
bCTMISpRVt4EZ3+MVidm6aTNvYqs0UbhfXe8HVm9vjvSrRABFJDRYIaEzvp0WDYhn207qFgQWTc2
hTq3S99eljIxrMZzg3dYKU5tzRZY8ATqdHQS4iPVKKuLkpwzhNidqhbFChSV418qxtiCbym8cqH2
bSFdJuxfeOeMzjwz+NkZ5GheW+WFpJKZWuk9atj1GuuJBbQC5wKEDl/O9CEFkY1xZi0hhqcr6/E3
uTdP4ZL9VcouCHDUgF/WUdQ2KqIcdF2X4eqoIZWRa+Ww34FOzxaGY4Kbqb5LVIVTnsN3o4CIf7Z+
60uszuf++dKVChjSa658dpu5fgO/aW/txe/4jyoEiYIqu9EW4C2vvTN6VzFD+V5PHqhKbWTUpAGu
FZnBGThYgTrCd0Qlt4uu65mpNQ8qAWdtprotI7KbMbCevn5IkLByecK6vJXQLOTSow5s6b38A55V
k6VLESULBcycYLXJ6DthBrw59AR+c1fcHS7ebY9HhSelwyvYVo/qrh5eRLzyyVAK0CpXRExfEar+
RFysOWdXwO2bz0YpdIwlAZBvntO1a5NmkeZB5qwNka265rdCvEupsrVswKyzfn3JfAftIT1EgJPC
fWLMD6k6qd+Zm0HaxcwQe5RwvOwdicEzWiUggcXgMDuJ6Jzqr+DvbjxCVXP1pRb511SNeICb+pOt
tu6d6OsHYxmZKOntQSD3bSYWjOgkrFrZh7AGzY4NoYAeO1CMpq8RgfWLHpfNYgJzQjPaB75mDGXW
82qZObtDAj17bU6oFGZc9K2+9nZIRQNwuy9tHm9B7svpaKpIflNUaIPyietV4bZZatgAyeKs3SH7
pWX8FQJkY1cwkA2BE9jSCMVaIjRDYruGeWekEcR+gGEPu6Zxh+8cbx6+C15hI9PWqkGUGNbXQ5l6
04M9KvQADd5y726XHhvu0ZPfd9VM3psekk9+hU6kgerInpBskdnnzM3Dd9s9R6i7AP49bScxOVEv
nZZzwz9rfTgARodoOJW2pHhrLK3YMfRzU0mepUQ81VJlQgyrJhaozk/S0iQT540zAVb6MNbghWI0
+e3q39rWb9ecPNxmJkC9P6pWgC+WhQZyAwDq8o5bVvAoAQK8UUS2QfW51yr7JQFlGfjPuWM8Jfz3
ATIeeJqbVLub4qUooasp2CbcmCKHO1bAf8MgPf6lPUzdcJ+ag+QswQv1um9e1nG4frTKfJZlJmzs
XxsPs4s9xXEUQx2kyJRbwZaSmJB90wGXtPwhzqLO7vJctv7K+jEItztSWjsQAPSB0CbUUmcrNwnQ
bBqA1650Wp1m9o5JCcKztTRyh7jQ4CP4mbumjFKiDwrigMCYxd961QxXk4yYUx9XpZB+xTAG3YeT
HUylNQAhaErQVeuS7Ax+qeOzO6yNnv8wmDn0MkHx+a9yCI1ZJGYA4jwd8XHkNKRiL7PENYiyIHlJ
fr8hU8Ph9AWnS+fbvdUBbDi1pF2nTwQqv0gkjTNj7lXlcTYmrF9iPsgXV8Jg9E4IzPZ4qGpqsOYg
5p5Bd7aEfcEcpFF66Bm7TV0oVPy1u6uGjs0tAJFbIxamzov0o6dxxJ46za+7zNgp9KTiToM/FP2A
m68kpZ9C9cGaOMAxTBvYqV3SAWUWGrqjss3+0BMLH4XDbkz/ToE962V724JU0nSRLbbYV3p0/nRJ
u02vsAUgAubqaGwCxX0BZzXlJReotb42BWVwLGUCTIeJh4r0zGwaxmDHgaRV5DY0WAAaY7BreHQ/
IQrENQWxX1ZIYBPBSmr7l34Pfngb1/nO4aqEKd37XoS5FmGCVcZ2xGxB1P0hUHUeTjfs20Rd+n7R
Xvz1zRlLLrrVMZkL68wMo0iMqFFcu28/M2zWsy/6qpgBPkbutF9yMRrH3/QMoAFhP6YV3o4S/6Fi
ekjr6ss5GwDs5c9OpmE0Zz019S42lGFgA7C02WNMbaFtWDO7MW4BawOLNMuGZxcIxY/7FsJ29vgG
lDrGyAs9NO9+x8iEA5jxP3FxWtFTLK14k0xmgfHh+9aBzOgDXBbaZVRWauTU9ozuSQzPMuRUiDV0
fK2ldUQJ2flm9LxO376+yrfgVnJHYe6+z0d/NVkHaq/C1qE+4x/rn5WQhiOD3gfNRjAyVq3x49Oe
jadTwmQ3QlelTQINSvB8l1Sd/cPnfQvAoItDNUmJ0FnCStvJ8EVxVYsdf6H3EEgDN6dbAjTjGHPy
Pc13spisyFqtJk5E7tUJtYc+B4MCKHZUBqAA2ttfZyDDYPEU5ReqvdO+PZA+N+qrda8vivfiX7ZO
zZTC1X/Ob3GLPhRm+ORZJTGL5y/GmNFBvYo0KfC05R4DoBfbLG6qbYoFQ0cX7E3FpvXp+GCr9Xav
8Old+AVw9A9NIvhpRLknss2y74ZRpTPvXuO68hclGrfoONaY2cucHTx0V5iKJ6/zpiiolfnXlwFB
lGtl7bIE0ogrm6AbUJQe9dRPxB00KtbAqIRYEwwklNuRXnnblxiOs8JYINHaWe5Onk/oXq5cVegD
ywSvGAM6F3dodRC5ZGkUai6HsXyHNZ/p/adXMeC07KqgRUY6+XibHylHCoK2JCtmG+Bw8VQdewqc
Re1C/XTfhBNjNbVnqXpD9KdljA5IWlsEgAyxW96uKkeE0buFqacvgWBFs3U+zl2w0lBjA4TSKchm
0PEWK+AYrFVkKQh9tC40sZS+ioI9Xcd8HjFxWMp2lpZwQP4gd1Sjvqycsp3qU5xud6rkgrz6eEmu
tK17416Uy7ocrRXKqcE+29KpYIm0FgF7U2vYMncaSMVwGEUrGootkiZzuIXc/EKRKAnPhZr5N8AE
wRMEP1jKpI1C8czok93T3UBEhlFm3DeqYkPyGonEyFZGssV77dPWziZQ69/HKbIBsVuT75OmwO7I
MJfSyipNOZ+RzSXyw3PJBSucQT74j5CJmGBXbU2id03hd7tUX6sk6WjIWlurKJyI1UYUQz72HOkQ
fwgOC3LIR8RhPdVb2tVwnkvQDwkZsTN1dA8dj5/yJ7EL8zGkyf1ljLO4Npr9IVkHXBcVCj0GNqDL
B/FKXVSi/55Y1dMhkmbYsJEkAyXipEKWxUWhrpittyEWPzwnWtZwOTt7gS2LiyPjmTpFHiLe1l4B
WHF6/sh4bzHscwpsMy2cXDYxTKRWqK/U7zDD1WNXB7HoPJIxQ5+X2yXahmfWP4BV1fTmI4TfEmWK
pC7Kfs1fhXC24ZDNyaTqHXWaiIfrraAiSETPhtscEyzw9mRVJUxXpWDi7cD4dMUQmNoDsztqhllq
JrLpglG+efsZAqYWgX83AhAKbjB4DNnia6SE03XoRSIBk2K4P2CWXpQ351LVNGdRU9rsFtYawLxD
DrzFzmzdpvJDeb5wkkxp4rNugU0ru0snd257/2HZer0/rIX10kzLxUP6asI3BihQsn2lFaKbHVUo
DZkr0EPGbO81uGCwvWQzotqrKW84Wi3jy22Y3oMWcI/Ie57i3Jjuu+G+CJ5R+dSa72aktYLxPOqn
ead+WMbgzjsIZfmmUhpZFf3BVombNNCTXCt+6QXwcoWOkfP5JmPEVDR2BJyW0Ch+2mIZ9ynm1g9F
RB2viIdWoYtiJVmPlKQc1M+MtsW1Z8N+bCmTGrTE7Abr2ebp9b89WLPs2uI3GO8zknYLrMf9PYYu
EpC70JoAIaoJ+8VFSLhZo7gTDZVfgmsISD4zSYK+JZqE67WJC5FW4F5sHRmoC4S/npJ5TPVFA6VC
f//YvX9vlyQDAPrysnMs4V2qvVrpLV+FRMDrx+EcqciYcR8OTTIqeCT43Bf9OGttbq1IroCjsNTu
gSrUf81MXeaZrAPUmWVJSv+WgAzTbLYTVpz9Y/sogzEtJPZvM53tZdrlxZRSF9YkIm8IB9S6RiJD
vWO8UimoCNGEe0z6ZbWDD+YldSUY2glR0Pr9OZmKddaRMNTUIyvh6lKQx2tNiHDNAx7dTmDgukPP
ZiSBHld6shs/Fh9afHCM2o+tP7GaMo3LHTqqe6e5VR8aKVJZZr1johDQJBUrAlF7OvQsiLUMuq7r
0LFD5aTg26BuZRwjJ5HJY1QRwu+ptI6GL7PFQlkNiVw6A/ERPBQu7j2zzemznd8MOJPdQ1byOjyf
2g348PUBuM8vOuZynDopWmeLe6X/VdNtEDOi6EcevG00Fg8cZsaCN4/wGt4GEMS0SLeZtfdk3VwI
ksUaoSm/Gw56FalRVdQgBZHaGh1YoiRJVEVpO/9E/V+e1gUqNJgtxHZ2S+0FzL+lZs9hoFvQlJ1o
iVf6xSYJ3CtfIgtarmdR7hgVmHV8fAQvJBZTMY30yFGtGh0kxhUatlJsQNISx4dU7k+9tTWCVX7a
oDHYakcbKg2xT/+Awy+q0sh5OC62+nzL9oSIbRhLvjIwbO0ZjHWvvYERZ9d7N7PKZ5+AIdtbTxZr
vENsBKafJ4fLf/RcdXFwkl6ulJVpFqZ3u/nEo8SH5LBSir90Y+1erk2JC9O+YTS5SEA8cOg/PfM6
tqStVLHtaWravoQLfG12bp1CR4zQVNIsCY1Iu22S0HmBGJHg2DazPgRWhIISva6dsn6O68LFoBfh
7wHB8mLVShffbmbcbQQZqXZxNj6ZCe+8QYSrsLcrrZzqbm2897UIlt5NzCneN9edkgxnXdOvA9RH
xee6zmnB6sTJKh8ABhujLYkMMp54U8g1PyKo9y3zjD2yvNCSlbjue5/fXFEyEIhsyJe7ajOmEemE
9MVUYDZJpSx4wJImUKaL9dXDGcHE56lz3EKiJkSvm4tWQib731c1M/mXyEqFdAKdyRJApc6+eNPK
h2wSUo1PkaWEEoYa27PFwnvhz48hnrOMiiV0FDi7FTPni8TK4de5Qi7dCPGf27srisNY9y72QaUO
JiOeGHfKHto5289BrgbTG1RkuUvWomKCQP+xewDUFn8Ch90vhc2NCrdujgHNImamtKooke/EqOr5
B8vfMfWdOWrE5BsY0vNW/50E+0FNH2c3IwTZWC0rCPWbNqb3nHfhvk7TSbkFHGFyDkQQn3Im3rm6
qfWna2rRZ+Q3jw8et+NWK1vs/FNG8G4G8zrFxnBbQNB4CNo/0GblGzsS+pVlI1RqPiWI3F7dOrou
Lzw83tdXS9RGEBV5ZyaLMVGl4JNaxyL7caijIXZRJPku7gvCZ0KEm+myXaf6YVndTxnPKG2TiiCv
V332R5acqOqfkO12a0DW5McrcgteLPp+s62dXXAdgHzKD8Wr17XoKY4xfZKQrt03FFJRqcAJpWcN
RP7CRia5R47BYvy2tw6xxqVOjpgP+U8ArfIiycuUpvOgwjXEn/PDDrLptn0v1BHN7/4RQrzVK9N+
cfNkTh5DPE5qESLhm72pUrVjgavcq5P1eJA2S/mGmSuydnl/zHlMiXvHNi+WZ0Vjhwl0U3c0cbPL
Y+NoPRsiWABgshR5nABolaPXka3D1UQq/JOhui3EaM3KO299BUzJni1DXOQ9Vul/0TS4U51jDmz0
3SKXcicpZXYE9m6NlIpsM3uECmqv7ny+59eNyb2+X4kfob93SLvv2kc8xooMfuFcSGo1N1qbnmGK
GmEZ9dm8yI7Uhpck0HQMz7NSSXKSSZftW1EKACQPWahEK8K6YMKVLvFPn8u/cNraS6TZyu0+vygx
NucpVZ1zxplVeFFqVxIaqcDMYxrVZDfAv6qvOD1lWzraE7uhoCDG0I9hDMjuBukplyb777Uh80HN
uGGuP9Yb3seXmRaHyo3MPX5Ti0Lum93eR6ZWEN3E75DMAp+8n3pEMeG5SuX69jfqhezoHO7R9pNK
Bm0wl2E1uaIvgbTT28FoaH8tAdLI9gm8HUkKrIEYyeDeBFLe+44/NPloM2+aKcY/a5dcIOPcyOPg
uCAHjwVZ0S9Tlz88ZxtnUbVJc6hm0tNMZqANJx4bRMf1edrwqsTYHjfvle49OnKnElJqxSyGxK9m
ArZWZpIoUvu4eKzudKopV8OM2Ihfwzk46CaulxbDHBbSMB+wAzU/iG7GOVma6j7l2S3Pm/OrTU52
35vLUkvDtBrYP1M84b6h+TCCPMdFnxvAC6dSsya0TkJK0TUSsdCfY34U8aMwavlTzkWueMj5LhsT
m7IhXs7PxTm09AAC5p0+R6HUOdfjPR5RVwmBfDBq6ESIsojeO19p5HjUFYwxwfNesBbD0J9JJ10F
0f6u8eXhhQn5IYgXkGNBcEZf+chQOcsMFHx60df8dIdlTqco9XYk3fqy9rvswDQPkFYTKpz96ikH
cy71OK+NraBff4H9rbO0YzCrVPGjdg19qbxxjqtnJMV4PyOAjNRyvPJop+4PmUCTkatOFhJoufDf
7Yf2svBcM3j1xuMYyCEoSHN87coSBnQOtluWj1uysbMlZbJzBo4GeUSVBfrlmKamT2qho+pwTRdZ
w5wI8/aiwl69s4FkDNKqobHeQrLJg8KN4NGn62Kzhu7bWPE+47oxHNg/mH4q5tdSfrju9twsSc6g
9Ei384Z40/dClSI7uXASPLIPDB+i3Ane8MnoPsDT5z3oG1cu5gsuJlZTfI5KyZSEc9dKv+IskhiG
I6aBN21pkElBZgHRxCh4jyTkbs76yVzlWWvP+uLcEao7Ac6wJKhtzDlu5fLpVPzqu4GUKUpVAmj1
rYTR1JG0iJEyhpiojqz9RdVB+n4xu2HuEQ7qnrh7bZ4gyIfBs87Zn0YWHdf7/AakIR/FWYslLIvy
CcI+RdKD8NGIxHE/OF1S8eyguNZAztqBQe9Z+VtdfVromdrTJO1mPJCSKzHpJacqLtvK3Vzaxaak
rL/4LZ3nEa1bdgoowQi3kDSg2E8Xt+JGoxJvZt1dEWP9U3hz5IYCpFEpQEG0NAYjik1yt3FrfQXE
7hEv7yno1lW20/8w9doxwo18+y82GuazREPZocDTih9nOhXdq6WLsMuMiAbCso39HtbZlgZenGIB
o/cNLpPI3M789rsZRmfS9Yd1+pHPXZrm+2hv8rFzW1mrPPG+1Wz52lLNe+PBrCmh8M2eZj1lIx03
YJkAsiZA42tkYUMe0u6H6meq4pGy9a7BM/HIKIEY1IWNCbK9F9mWUzUELa6/RpwSknhiVJkVW9Qd
t2d0hOT+CZ2giJKIt6ZRBEqfWLez60G2smLe68yH7vm76x0i0GKOa8DXe7BHJsJxWG/0UoalPmg2
Qu6G+AXiOzo+mUtCINgdMw2ccq0EJ0ObOQimcG1DApwDwwTVkjXmc8IfA+tO9YJTLHr57RtqP6R7
jl1LHWK3wMTuzryHVg8GlbDR6OcHscUfFZNNlmywgPR74ykV87p+nrVM7ZcPBf8aUe0znJ3kJTxj
K7eLQD7jfcZio3w8AGKan6NE0X/wy5TY8pX06OsYWZcOYuCXRg5Nl669ep4eXosj5wKt7pwRNsey
CrAwSg9taxaCsX2Hh0Ud9KfZfJwpq0G+OLfengogyyCt0F6tRpfPMhM4WK6omt21yD8o74SfNfwh
rCtCUIK9eQB5xpHfmrso8p+ipESxoS3lEOLr5OB0NQIvlyC/wWWHh61Yp4Z1PxDr6ICX8D0BzdQ8
ycrWoLfuOQ4usOMGEls5svhBa4i9WQs+DHeFe03xKOsqxrAMScxygdMCpyCZllo3fQD8aFxYk53T
qpfvpgxDg4JiqWPSppaYyQzFlRKujXHLmxXF3OZBVppTx9SsBzxIXJX6vOiop7Gh4nUrybVtwe81
ufZ2tOg/IRq+UPPcrZKACaLLH0QkC4475+ThYRxS3xR1uj4/fvly7ovaTurgtaQvdmfEXSQv7nXl
OMSqbULAcyzHtTxR9Txzv18NxF+3Wjqwer5SNknGBD3VbEE7IV9MNUuJlrGjUALuS8v94Yq2cLkN
LNRIUtfsxDMkjTk3YaiFtStIYuYMty7453DPYFha3ti5lLZ6F8psqbv20bbJTWhv3szz6RHTzySl
uopKVfvLazJz5L1PthkNCdBF9SQzMeA1OfiCe7taG9Y4KC17rnnzZbHpcJFICPqYQttIFJz/3SsS
qpRx3wtIPDKPY+BzHZiMl7j1biJYQIFH7tg5uNJpD1LuLAYq5V0zRJVyBlxanEAKAApkvKF1UBVC
2vPaVTMsX9WCf272FGyyEg6Ae+8qjbGA+Y9WT2u7Qgtny6S8Dn4TayvTe4OnBIyHW9DKPmAkxKxl
4+U9lHDtCRNEn+KAD9IdTFZfOFuhShCYoQ1U5BWhEuDE8VdY+EuV9ZsPl2SVvXSN57hqjB+Tc9Kp
ud6MslK5OWJV1OV3Rc5tz9gb96lt6/6a6wtZwBkryGdwxM5jbge4x2GTZ8ewPgcIgskdwZD/5e3E
FIAqmSJkUnpoj3ZJnYSplkQE+OdjkjuygYGkGW4Bhor0OJnHnUetxgIIzIMysq7lAywbiKDsKEnD
wgT5zDXb+nqBUPyMc2e03hOIgwbyPtY2tuI9nWue2cK8ekfG1tR6T5qtdbxP+lIhp/At4NYD6lq+
dfGY7U3lDwmoMxCP3CAKXOmAXkdwkUYTqtxAU14gXZ52TKxxk0yXQPhclrnjHnH2fN+uV/b4KYBQ
k6SkSm+kqTqj08udrybr3liAvoF4yofw8SEOOFZYStbNIj8hzNQZSrpFYw1UpwlnYM1BV4eKIsBG
zyJX9rDjJ5ZzVFWwTHkx44glZhADK4D1gSXQkvzbTjSm4IV8TYfrqjf7HRMrDfnHVs8blhNnCK9W
ILdNJsPH965HRgGcBpTu2sX0K+OS/iVgQckRvQGvSyOKGnZUiJo1t0r9s6LyVN69r8hP0oXxzAh3
WOPhCSrnUfHeB+9DdDeE5wA7DzHrAueGpk7W6Xd88Op5HC/QhdrFubyImyKS3NOJGQ9l8DKhq2tl
WmOL1BfraAO7OcgxWJu+OE4QXmZPk8Yn+vyHODO+j8Hy7BdjBclV/2HvH6mswx4kwhgw/hAY7KnW
dIDb9KogKvMzwV+aca6yWgCBTxqxFTyiaTiH6MPYrqQDwRo30K/pm1Ny2uIYIu+B1HfypzcgGht/
woH5Liwu7qapP6vOY1kqnNTCDBZbwUyGlQUGsErAB3NzIGiyc6E6ALwjX+b8rj2KdO1EAz153Fa5
A4YgRLzoGpRbBDUAo5vl0F0ENCfZAkUP+T8qCxhEN4xT11/+ZChgRdR9m2+lRv8LB0c5aHwK7fSY
WJQdJHon+aZPaoTXox12Y3nvAam49qFUqH2RcnWo4+8yNRg7fi9Nu0I/TJRGn9R3xS2tIHFYzJcC
GqRSMg9czhh4/2Z0/ufOVtEYmA6f/0Im9NvhxPyZiGf1fbUEcpJW+hdpNjfv7Y6M0MZ2YeIXA9o9
kBW0wY8AHU8xBie1V59S/1IITuVhXriq+RVoSe4B6tBJBSMT0rZYq+ojYolI2NmuYxXhzdIunMfe
whzNs2Qndur44n1V5wHNpnJGbeDl6eR+eKWbKeEwn7wzJTb8SEpEPe6IlxgpwcBz6Drod1cLh6kr
8KV8+9rKm+pKcMd3c7nyHeseDAK4IZG1JNbHzfOiNHU9tQ+/5Ydy7Q6ICopxEB3aeuihqRLtXZsD
9JI0R0DsJ+Cvz1NMsXyqYzdbrMHTiw882cG8fnNlRxNJ/1fRwA+LUbS6r3xLfQ+dbGQUSoxbYt2o
+IU042nIKde+o82QBSNDav+igyK5R7y2uMiBHxjFTV1eqPMrvuwb3pk+W28+LlnrbUlng/5V9+Ia
jXNQgIdcagLesY0kZX2nq544KMaYghFhfrn0MPAZswF/bbLkKjCeMTc/Om4rZmG/ydVOqExYfZsh
96yMXIpwq0E44xVjqbYdBXC4RRmFtY+SYNDp5eQQJYTB6JI7AtWsc5qnOT1rI7cI3ewmY8UOODNB
z/86GlDsjdbmH4/CeB8AsJ8amATDKQi/+KNBW2AkGrQVuH7EpTrhbUkOoOScQ4IFbeoe3suoM/NA
wy+FL6xIQA3q2OyQarBmIlPq09pz8/UcHeaTy/mqVRlkxasXWQmkPpbZmLtcqPcNk+Yl/xDxznUU
X/cxdfJRhmclu7AtPORVX21pD2eJOyl80OJmnUCnFL+0tPK9nL/EeGfV6+TyAduJS/G0VAX8dsl2
nbBBve5SpndziPdc2CXANoE+V1fcptHuq4LTJd11IXFQq8WbBLrLlHpkj9+Bv0/VRzNd6ioudCT8
nZ5xlW2BbWj2K8XNx1FpXRM/ih8uh7f3/aWtg2MwgRMBBUXxGjdSl5pMVpwc8nKRkn2mYW7zliUW
7NRfjj/fhASny273n4KEfEPKMpkqZrmsdN9cXiJEhJV/LngRQxbXaozC8qe3jKQQzmCjz95vovo+
eN7CmrI6qSoRPxIxWUv9d2pePlXUhrvq965r1IuJ8HVxvjBeCmGtzk/JhCIFWAlueIkUH4RZDpAw
0PoidvBv+29cj2MeaR6sCDivskGeYE2AL2HnIpKzKZWNJoko/9V8yjyaLMgRepjEyah+y1lnnDX4
o26Lc5c8FDyKzjbVzeYf8O+Fe2/JcuOcWVgDtTB89hglZy3UICX49Xwvn4bAJm72/H1/0RWUzlwa
U+3JLjzgxxxXZYPVzrcnpEIzoplVhWS8mtuT5Qw83yI+S0KfFKsrGRJxC+RpKLRzXIoHL6SszWMU
lKbz/l1k9E+2KjG83la29+Zfe/uak6fkEXYsH4mw5Ede+MSY23m/cI4TDdAVNGgVVbIBEi8GaI0r
4CBgltn8JBHIijt8SFiaoXFb1gyLjzzx8+oK9zt14+STJZpetVOS5ERx4MawVulHLwdV43/ZZx4i
wX2jWngDQYQqclA39jzoR3q3nMm/CCQnBS3y3ybOqxl01cZjh5zx/JZFIvwnFSDwtbd2Vuswb4JX
AZ+eyBM9YejCHDoDY4yGS3sQ4sp+tvxZxeaqstZUBJ19JO13N1UZuFkFrDFUQ3mld2Zs3qd+0Yx6
BApsqJXT3a0K8rHp5eM7piSw5w77HwqsSKWrPTALBQrbka9blESDfrN9yyEjqACtFDf7nfLpjqLA
p8peQ3WAmhqDyccJeqNwwqf8MVOMcWTwrfhsWXo9bjS2p1F6KvhxFD7QYvH6oOBLAmoZprTROYUa
VIECwBJ+NbHXfj7DbHyQ0wkfPI/T2rel1Hf52JPIaYCqbCOYgcIWk4+BPrevN/WuTEKjhkYRklof
xXGgHvOy/UKkwUrmqEiHwy8YfywZVY0/i1UEOMmUAWL2Vz4F0FvBZbgMcteJZ/9VdCYN3L7oBHwv
BI3kqQNkuily8huIfR3vVyj59g4+5wVs1dkhzrU4RR+NjNfYy2SuUv1T+dtK9+Wh+0dfAKNDRSJ3
gCb4loMJs5XYpW5/W0sP2wxLzsHlE0PW4OJ/oJdmfc63zZqJRnrQzCMqKhrBSkMOGWtUMeEbytYk
Syoo9Lb6o/EXH0iDUcObrgS75uhhVVHhqFuYpzDE9KD+aHuywQwn+s2Oa00OevhHMZE1kiB3Pp7x
RbFX2X/R1CupbSDTAGBA9nTE+h1e6nteITGPz/UCNcHPXVcqlQxL3vP7XppwIN+eroKAEioRb4UV
oAi3TaN85N6eqneBHzj0tdnbPw0QXHlY/xO9TsMQQRJ7FbkgmoZTnWaYSQ6Y17t3WWtvSGoZUtan
Bfpr0GCVdeoV083FIRJtrUj6Y/lpsymLmA0P3b9rIJzPYqH0sU+21tfVJH8yy/vVXIFVZ4C+7AK+
Z/MR8G8gaqVbFVgMFdxip3r+lBfzcMgjZn95zu7plpZr9d22RiQByTor8i/9pYWX+i8J592IZHXT
AaymgDnDKLRczKhtqyZuRGz/Zl9D9JeaylMviRqU8MTwfV2Ffkl5Wbs6qJomVVetr/SpnhU62E3F
hom0SvDoo/fEwsy/DY2lo+IACe6AcvM71QwDdepuz85JfVhkDk+Jf20XdZR6OoWFlBOfFT0rerPZ
ge4OLC083tzCPftJ95EMF3AfpKEZpJvXvpVF9SJwcpjmTFOP4MD8U6NukZtITVQZ6JFJFsgSpFBo
jHbku5BR5dFuZJt1N0EiX48MaNrD1hLPhyYtXam/EpzMbwXJw9H46T5yea5fXNaqSjoSNEB0WptG
us1NzsuGA+o74a9QggVUg7LG+JIcWU5tSwltI/kogsy7bMrg5SiqFEokYZ2a/vxHJXG7HGwUBe9L
0KL+Bmpjw5w8JPsL6WzO7omryZWYordUqxZQl7Q9Q2xQkDdDYXRJP2KKvTWZP497sQBMDg3iba6u
Nj3Cot9pKSc9W+YCyS5Y1uHiPFjVs2J9fY+YoJT5p25Z+iEqNKgdRuRKiTezrqlQBP1g3zr4Fgzc
1P+Lc5LVl6KmTVePhWM8z1bvwqkocxGVhoLRSjaM02RBv+1Mslw0454Pz8MZp1nxniqKcUcUGFmO
eKHhqXfC+VlGMkZVAv7C4rVyg+7vA7ckfV3fNjcOT/SfEsiazW/SZBJ8TGpzkD2AEfjd/jXjr46h
Z9lYMlolIZQv95XxslXMxHiMdW4ELOsQwvrDqaXggayxcaajijKODhbS4Rjqx6lZmW0dNIPJwQw9
73Hxy74mQtiEWh8/e/0Cd/MklMDHMK+0KIv9ux3aOiU0Sk//r5axan1MzSSx4wcCGXF61SDYq733
6pojzhP2xO+nviOFDOKqpUOOEmXzIK6vtqFf7mb54u5H4OsJZVEZvFquztcQ11LpcCShLDT/VGlC
KM8TDBdrNWeZjnTBzUW73CWbHV4CWzp8m0cum3Q5Wx1yJqdmsQQnOZta1fc0Jad8zgmMP1bXBGzo
l9NGYT8DF+robR0pGGYiwfxrLPu1L3DnzRULH+KxU93dcPj+GfNb7Hkidcc6vOXvWTHw+GQu8r4Y
0h0AbSqoL6dy5BfcIoOBmTpY5ne1IjdX0+z1NvycMq2HjYHcP6Ty6sR1YkUYd/tDN2X0bKeKB6au
i7rYxm7SXquB086A9nHr4aT59sYifsXQf/TBt0p49bY30ovktrV1oj5THijsBkel8sJQ0XQ5UzYS
yM18rMze22lCXTuJHW2W2yGFJIv7OoQzq3zz/zfvqfpjV40MvB6Uke4GoXAg1OJpFIad3h0EgpCN
zt7dmbvApVZ2GBxiYvUo43KQ2W2X8D2Kwrf0vfCFFvOCtE3IAymBZ/lMm0quqcqTrXtRdXXZg0XD
ta+aif0cdL2pkNkbznhJtHFPuxVJMrfOE5I4Oqh28J/XX16MN2jDifMYTQk8LGlI1ZzVcn2KwQk1
jLNax3B/r5pWRpgoe12FuTapsKx0obpxrX/9GR53ObqL267aFF4GPjrTs1JkUkR0CtKkj9PQjSeh
j/ilfZeTckh1WHcUnng5g0mnLFw5Q4i7cbY53uCDAJpfbjaxNqwGeGnK/YuLLPmgOSRF9QT13pRf
XNlV1G+IgBWysuyN4pCOth8bpe7F5tmOA8dCs30hMJ8tcuZgshK6jyvuYqTw5KgdM2JODl4LLTkF
wETu6nIMZz4S602ph2H37bT9icXtQnkbTsPQ5VPJ/MmDdi4Ikj9Q/fAKhNCxuy1VfKTNyQ50i2QD
eJpD/KLsrGwhEYuutkSp2G4CWRwAMw20l31CHT73QLg7CDkBF5ndMk5CDNIX2iuTm7Wyr7Asm921
C5nVKlQf7LJ/VbP6O4ysJdycf8ac4pb+Ae/e6A5bCgBu8K3RQoqX4+HwBhF9drNMwXj6XC03eHgE
QQElmUAI6sy9T7EnCFp7Tktlr+U6a3xGE34F29ZocfyH58PzjHCEXUTmAdY9aN7SygY/Hy5WgeXS
OPKj8qN/ve3xYkR3CsKRF4jvWfhjDhR4ICTs2VA5BDLI1GfW/kE5OwpEsIccP6M2JcxPOeiKjuCm
zJ4F8yBrYMsUtsPymdUtVc6nxO1kv4wC0JiJBOebcRrpj9GkOzbktfWo5FbgBXO4QFENCWx34NqE
8QEgA8yhIYryxtvv/MAOW39utlRxptEgG5hAuSy9XINxaNWVgaweOI3gCsdDalK0vRxOpDcBX8pd
9KyBcftsiE+zEhp8nmjZ0j6bB5Kny0SDKyYvu1N9Y9tStFLC1YSkLdz9mVck/nNIGyOVsOQGTfMX
zwqTm6uGOCB7wSYNpXKLykamDcVUQM2olx1qUu+zT+7SOhIosrjUYsq+nGYEOknga17gIG18Nxtt
Z42zxdP/U8aaqFEOZcNN07GBsstl/U7K/AZAQzNxOs7EdTcTVcsO4fy/JI0oNW0hlHvWgdmT6wzA
gWNL3vMJcuFGRhVPi5K5kwo+uX9qx2kYEkJoXMtpnAcw4FP6pt3P+W5PeRHLfmtf1VvYMvfrE3LX
aQoyKchS5sgGm7D4qD1/zggeKqSZgK4Qe5RM+9WdZgKh4Y4CVLpZ/a42elwCPcIZIDT1SztyAOUU
P2z4uj/10z1fjqmftrGKs/BuBA1bX8oi7KYf1zH2X2MzaxUAb5rR61f2WIdAAma84uIxJ6zmMVjq
H2ctMKeeTW4VurnGWZC1acrXMAMiGtwAikfhAsEzQ4Pud/XJAD8H6yLjpIOjOVk8tI9+0E7jOqpi
tWrowywLA6HA1snfSO66KuEZZqcDPjqdhL9lf+tsHKqeboWD1t/ZBdYcDGPwN/5SfDpkrWLMqDeM
NPZ5zLQ8zpW7/B6+7cxGlRTUbPXBLlAXw37Bukhrd2yzze7rpd8YRgK2+DCN/8q3vjsxkRT9AsQH
HtNFnwdUiVb17qX9OvkB1n8BhK/CKoF+jyZITjZQXkuonZGICGZfRC60NAHvIuUb3DNosEW06fiU
aIr6sY8UzsuHQd3H8HXB9E9cNY+OnOflNeVE/o78CpJEA+5nnDVrHzJQNlFSfLeyo2ZfEdY8BKBm
NUH27Wk2oWb88KDb8MHUSF3gcH+H+3UzWaf/90Bko/sYbgtIcwv/yPs1ps5DmzX1CVIN+85BfY2W
KFBEBXBX+PACO2rKj2YoudSL2yFbdMzbXA9pTXjSWjPwwCNEk10P4WV/YCByaVfG4S5otTtEEwHd
dfBz1/9SP9QLZndM5ndd4LXg9EE7J7lbF/Trth0EPaQyBv9Xm6FG9qLDfRDZ9p+lbB66aVaWUgzH
ANrTmSDub8bOd812Df0lY49aJ6HbFSBtujOfiMSElGHUeufuWyQ8GvE4dDpaevocZTtEh+TSKrER
64ohfKj+9m4vaL88RTOupt3K7tcl3Mw1bDN3XoPtGXkjqnsfD60W6dmLdA7QRzzPMwuk2B0FFRH/
qPXX0R3r192dCC68hviQQesH5bnxmLUQJzDCi2a2WiusxfgKjNPlJ6fPKgua3J/r/BUALVqdUAFf
2xS7HLO8E3f5HdwphArqgMrn0XuERbUIGkL+DFdSZupL2c/auIY6L7FW0ScO/lAoX3N+93bZFLeu
XNCSMHx+cPrpUlUOs5/LOXeidlrqjfUxTc0Qyz7t2LWMFX66h3+WxJhFAvYHtBfdxs81v9bV1rSX
K0Z5ni3Pg+o/S1KbDLHul3Lhz2kMB/AercHsNSEnIdCHfdSntUG2AiQPuSuQwsnv9KQSc6tKFhd5
HMTx6T/5TX5pTp0h6j3spgcRAALeGq9qXyffMYfaWVZ1o3HKJwpiXO8qEPUdCW6yH1/6keoT1waT
1b66QhwB5P83sOXcJaxTM9MdVT0R0XGjvjcWU1NW8yzSPkc9vPHcSDD35HKjoTSAQMydrtDpcZJv
jgmDb5370P5rNhQaK4/faYbgl2Inaqht/YUr4UGBDadWrVMkYsOyZjUdmw/seD+8OX+uCTrWhR8E
rLd/tfVfTAJ0ofXvmr1DgfDdl5fTyJCTR+CgvvxaOXITo58eTFivGVpcENJQyG4HRr+c2zVY6q6O
GMEB1sfvYVMPl0tXfwurOuMS2gsd2vqNCwihKwClZJjG9Mb4nYDQ9t3I4PuEw98KMSHMCrAhR1Xl
xLdxbk90IhN2+Po+chFXbXlJvADHm8iS7gluuYg0c58ahL6u23s4RhZHUs50UPg/9SkbHjx/njhE
4Yzbpnla3C4UV9hoj8+WKa+pS+2BgPXoDLLZPZyyuXG5rTUxmPOlWhb+NTZ5zCcT0lGpy8bO1jBM
h27jKj7EkonmfuaZbDNYpwNY/oA19DL3HYSqdsBUC7L+fcgEsvMjsh2gjJ5YCfAyBP45u45KeJX0
YJyBVFguMEskNvDmw7bOLhPDtWfdtxgtwhNQKV97CRGyXdxNyTJZySGLdbVbSf3ImgxYAWXOuR3E
GqxOIA9aGgijb7Zu1Xw+KYHMhxtVozkxbuIuZb2PJZFzIa6yzv96Xis1nclpb2OO/jwlxEK7cFLE
CQLK9Mj7ZzXM5Tr42eFz9kpn3ln2KkraXVPqJqoS+dqpp33ZSktXUEQ2rGhDuvlLVFQYelkRBtkP
4Ycs8mwy8lzlZrpBheLZOBqERqkHW8zzYCqaxv9a2c/iow3f5ryFghUnxiSBflwEEQ0egeQWggpf
a8cUqPSkEhyzmqyYrgHvLK5Tst+KwcJVUD6eZtrYLjmsGnzAe8nWc01KtQGpWbcEN4b9JwwWjS20
ay0YA/aY4U5PxmqySMglHJda1hG46ltp3OBJ4LM6Bs2QT9RG+zFJp6iLmC8XQv3jsOK1LXV1myQ3
5AD9yJXvnDXzc2XUNi0oXxb2x9GIWYUalgIzO5PbR4jpm/w/63lbUHF/YBiw+/VHp22Sh5Sx309d
vhICG1/EwgNppoa7uRbAPLtHv03soKefd2ER3VJ5Lw1sgXxpCD4XY2vt1jZPDsKWnYztBAYoCiW9
9O/7UPVmh3V1JBZouYnElixI54JaBCbUrvAlTGiojO9uAmj3FV2enFoL3qehnAL86EcMd7ewDrgY
YjBYzPmLo3I1H9lqcUL5FwaJQKrol2oajwd7uFIK/PMqb+sC/BaEpFNHijU0qsAu/3lseeUF60ki
j/B4FbjjhkiAU4sVO+2EMPEIXunIQ8tHUI/AZbLcMF9qMdKz/DjB2skgZ//pZr5DpXtefaN93Np3
qyQeCegRdeWtIV92/fb4H3wBvxoo8JIIEw3inHzXv5mzQUWtm7KlvL71DPBaZVsdkcx62bCB9XIx
4piFiyHS248jNfC+s06Wos4Oy65xM2vxl8klIjDTC2VnrC2775mhFzfFxmJcT2oDomUvIJOb9fk6
5uGFkbRz3myghkvacPapibtZ8wMjrWyHb7mCOrlD4F5CKC75nyX3O1QlNwzuVaNXrCR/zcqRB6mP
2YpuMcouEsiE2IOHwEmN+zBVm5Q7JRZLEGfkfNnhvYaxKpKFUpzn3nRJaI9abTT2p0xHjzQnPakp
PvJNTQcshrtPG3qydkuEYccSIGXULl04miU/xoFtpxBajLdAXpfCera7qQrhVW37MAn+VhEFDIF9
unXIAU02LBebzT9wd1iPTOzgN9WoKmeTD7AhMyk586T/f9Qc04Y7d8zUwibMpYWjihBZPSktTDxA
VORqwCSG2eGFytJWkiiE+5wkM4W0i54ERwcOZHhP0L8BS4FzejF+ZERL1qQulu0pzkjKtNuoa2nj
vqkikX33c2Q3hAIW40vfDy4sNxXnw9tdESR0MRMU99GDCVJKBwIvxZMEHTKPJ0qHF9esLc64lBvH
fF6dWxXU687n6r/S9fZPCyCYVMe4DlDZbylz+QLL4HXst3LqCb3JPoZLVIN1ddBVAVtaaAwCZI2V
PZAcI28KhccJs/Ckd1KnkAbXLlDL4fqZjv138Emg5Q+19W0bBasXjXNWhnxwDygq1sTSGjuEeRS+
WeB1F3Yb0pKj0zSVW/UTvQpGKZtsFO3lsiLMwiswp4zxAJgU5LQ3zFAuG1SADkgmlyYFU45DyC06
zWiOJ5sLefDca1UzMljSPMDQ4RSJvD2U52NOPtWlymFvSUF9SczYX5MAbruAeCEu7HbBL04VvkPL
ch2uoL7wZM/cwUuxnr31ouvWfQChhk+U1MKAhxWe8WmhenAHp8bFkjbrVSUQeFc0hStLLTIJvFjN
0inc0p4pmkMCK0TfN44Mq8o6+uvT5VtVPU0mAiKkU3mwlYsxjbvvN5aQTH3X0t8a4rWmVFNXWn04
mwyvNvXZqgpPgjXKhsfmHk6Ad+2kWfr5fFxmFGpwXJ5PKKzKrYDs7Z6bxV+mC0MS4rSqAWiGybb4
n5Xz+GA0R629slWTiJqoPzqcNIIOPCnSS36eErH23KP6B4Ux1TMl+9EqmW/o7rBkFPO3mCdDVAV+
+WmAAZeYBKRg8iUHn9nzNFGlvNfstajTIIjCfD2H2ej4gS9kEdvxviG0K930AHWC+r+qgdi+RerZ
mUPW049fEcwtCuJ6iET2wZNUji8eEHSBYPmh0msn4OSEidrvJlxBDbgmuqSkZ2pdLSIus5CxMtK1
LHUWLLKvK+Agv5vG8fZLOmuBDGcNvMkQW6cWnFWXa4go64RfUK0JLVuazDcjMEOy8VPoNNYSFuBz
iWsCIfAB1BwWsp8OjNM8GtByDzB0S0TEtHqDimEXrBO427AlDUh+leTCUiDmDVyOhr6yBFPTl45T
ZsGu4ZAr+QCduSAzdmYuR1sSxf8g0rdkgh9bsrLWcNWKIQo+vyxrkAPm0n2OwqgeHPyJmEQIFSlZ
rJGFj2vaZGxWs3v9b3jnTy9oRgkVvCDhO/mXLJY7KKx7FI0fHrlk2b6nNhYdKV4vL9BP2aMGrO+q
iYzqD0Lb0nIKYnTCpeuXcuTNRzzhUwK1Um6sOB7vDs0tZB8Y104GQApfLy4gwzkAltjurLQ03Ym5
NpJmPEEaj1HCeDNwtzGXfJO65vpvxHWf14Ln+0aQvk/EOQrIB1l6DhBemFOK5rNTizh0rT7CWRId
Tit9AeYEPQaN8EEeYvHZZbfE3dAn71/HrTDt9rjy3Vds36veA+wX2xUzrmJeEoldhrHGsXfiPObF
9xpW8FK1jj2MFzxcHDTsYIc9sbFFgNWW025N8za9K8xMrKs9NUmdzmK3GbZjJvTBIXtAT0QSHatV
ByINPwBco/OCgffLtYPLHOh7JwphKiWl6Wiuh4oAMxK1KufourQnxcLvfbGK2sPenEOrtuN8pWuv
68yoRjIguIs0aPBCV5WAn1xnBo+sGEA8HVa2/+/GtYn+jkgB0AlKVjPozx4gzrYfIrr3CG3i2mxz
/8zllCeNHhtn9WBzRH5VJE8dz9BU8SSWcDjFPUVX6QEDgPfGONQ2npotmfHn3BDhexOWO7cd4InY
0BEQDqmRp04N3MH5gSFc/wL9ryqNyWmBivjOXWl1O8LYmUS/ZXyCdt/hvnUf1oLDtDecI7e+eHNd
uNOiDgF9ZfiYYyk+J1LNvPki/GGJpYmWDXlafW1/2MEiFWjIjHxcp1EyXpIrdlZvtL1cHqAgGGt/
BVZXea7x8v14JN+YGT0aj5BG6t71o9gqq8Nhc77JLJQGxNm646M87zU8+B0moko1BR9S7cgWabp7
vAn1H1aIXgeHpmWwVWIxE+W+uF4ZYrOkqDAXR7pDmXhyLv1MDYNWuXetbGGDny9ICq8NrshI+8No
kdLM4trX8PWm9wG9pCL0BSPZA2imoCLgXoTjk4pNvPCHpud7Blz69iwYxSQsV+tDzrfDxpR64b2P
4owBa8EP1GfnOP3oWLaFx9MyyjWwfp4lCv/V+MeVD4QJvcbHILdWctRN4ZFSSNV4PY8Td6YshfAH
WQzaBxMc6CM62O+ZnMvUdEK3+As8EXPPM/Z75VhuyaXdqvT6TJzanmrDD5W6WRhS6Uvn2oJVCHid
R3WRad5afDRHoRc2/pi0Xlp0pYAKDXUWogKx3UMDxChLQbzus2THKYRk8IqzhHhm+KXCRIXMEGNj
2KztMndDKPXrvfNsY/+vuo7gwAohnz9NNMcXuftrd2iCK3H/DwDA5/IKphtXFxYvTsXFxOQD0oo2
MoocH8Ms2bDFmCfEL1BwUNzzY3JXjhdIkGx4kD28rm9cgh9B9+uc+l+3HWt6SUAQY9swZeLRXEA2
GcY1iiNqgbJjaZj4KMlYljiuSnAj/lZKl6TBtl9FvqPjzXqlQd92CcNzO7M19fm1Pz7kpjM/fVUl
YAax7NnASnOUT+p6ubiyVeXxCxqmwSa45iZ5kim68xPjqIKCg3qkkKRdX0c0T3Fr2FKoWXk1GDSh
8YFUmkOcSGAobUN1ZBvKGaXP6yeJfFpMz2N6WIyfmNfqSOBlW4mnXEilb6pmtXf0EuXiYpe4fX3Y
96/KxCQlbLe8t6oqQ+JgqM5ZECUZMwYuQm20zpl3rIgFSsymkLf6+2GvQ0EHWejMOPgb6MREOl2Z
xKKzO7Gs2u2yjDIYPH8Q7KcHUaKciTC/+n0oPm/8CZZMvz9YapRodWNe8xmUJDeyFzqmZd5esfnE
Ocp/KRW5nAsTy40tdIv7FxkzEdO+XXiuHzfkzBeptOktMKSgLQ0Hw0tITiRiwivXJXr8c9JOUefs
IWaq+E0XXZCnpaOqkRp1xybaDi/wtti18yt56Q6/7uq372wrm68FKlkxYti8XXGMWBan1YAYNb8O
YExxOER3oX3viRpHD1qIbvY8b1boz1JmDQEiRk2QSx0V+rkBjyTcq84htDQg+8Zb1JIaRKni7thJ
9UEUpZn797L6sNYwe1X3l10HuAaItWGZd3Q7+IC7I77WA7YYPEFfCcwWOsZJzUES/eOTegFEUS91
53zGP2Ofz5uhfEyunQ3IYHJihm2fHTqKbNrL5HS7d3g024CefD+Jg6n2XFdO2ZHyXR5GvBFY+svS
updHqQSBaBNVehXq6Vu5Fp/UMnrAoIzm4nhxpwMqOITymz9GORTpkQ5IEJDafB3J2wRh03Qp6Ao8
57iCdPY+ytwZZx6gH+sHDtP+LrGEKXyFq/2m3bYId2KwNPkYzJI+7YrEr2STC2HQxgHgBBxHxTOP
X24FlzFZpyDVvtx0YDMNVuKUy7Rg/jtG7EqB0Dd921tR6ANwYNyG2TdCS3DBtF8JOclr/uantknV
VbKxSIf+2I0UKDMGb5yqXX9w9tf+obI4wHPRK0bM+QJQuocGQRWhPkoqbTb1xRHyb/b5ds/T+Azh
nLJ87GfSLKNHmJGIb+hyUWT2zH4HYtK9zlayspra0mIb8Zp4WvTX1r/2ilyDdnq5jvsLEPSND/oR
w/j0LzB9toiEfcJgACMMmuh1oqcaQ9MJ5qT5Wc0KhyuLDY5iY2hcFBJyZfIGMBCrofGl2Hp+a5ww
UYulirH0R8VfiMqJn6vTGSSfHF7Z5I9cDe5wh20M2W/aZTSq/NP2lG/qunrU7fhQjvIPHLAzDUxA
oFaXbRuDAk+BjRypIumfUmx123yUoAqHpUrZu4b15Ac9puBFnPzP7B3bk1kcvsNciP7o9q6983VP
pDeK/qWqLfHeQ1hGOqG2u0th+Y3YLtOKRYTqBr2ofcKRyjVMtxbBDfK6A9uJASnD+YrJEujTE9f1
xTgs7UVe+FcDYrnPScyIbsxHm/zERAjDoGyIdCMkzK4uCgwmqPFKmjBZrRni8uupIbmMUWTarC+5
FGpIHH+weWHNyLNM1RlFOCKiW/BY0OG7n3wDQzfW54rBewt6oFxFHEKHQGa1b1wjVIa9lGmnw667
RS/GoWugWgHibXvkfCFXrACMmn5p7caevZO7xcdsBPOfI87AATxId9BVjq6vKnUJDmM08v+YUVdO
G0Ib9l2UqQuxytV31fg8fDPIczy87qTnjjJoiFmRz/mJYo1iIiq3nBUTk8w/IhDjOrovHBLkc6O+
v+QqePzTRSDVzSTnFPqDOxQG4O0+Ozfup5F636Y4KhfwZoDTf2c9iYbVJlNKO2SBmfbiR9XzhJLY
thqUqkMlBcKhAKTKCOksllK/A0qb6ho/X7Gb8KmgjWmKM3ZdyB4PovfW4BxINWA4tCPs/7qne6eZ
l2K3NweEBMHrPAghti1vr9JdWRiLJrweKN4X9SetR175Tu0b56r2h27FiH7CWkfCs9LEK11Vdo70
u87ucKUxao+KaTNf23dfOM9CCniF2oxQW5RXS8YjjznIM7z3Y4ZptKhxqGgBr0P6MKzf20Veev32
UTToO1FTuXTrGE7x5KR4N5de3j5uDxT0nNdRVkejmoNnijDSCRmwufQZvUfqksRm2UNjc+U3wNI1
zOX1Si6EhXhNAAfHaCruOTJ+R7GMfoyqC10/v/yQM2SNa0oDDHQl+evcNkOSVsSgQDpetlyLysNs
2RvBw/DXxbBvuGaqqZk1eHqDXbdP25r8wW0vikjAw0gohdPqZiy7Gh0dB7jAYqyIYZcbX/o3LHxe
eGAtxiDePQeu2axXWGrhBizmHOrBVqwD3RR29DvPqPpM9OlTngg80oOFG1WBo1gxFY1RS44NodKB
XcqxrXe6ER8h1QtgE4k1jmke6FyHj4pdMVBGBgOYRVYN5T/MjbO7ZIDUM0GYLQSIsUjZMUhSQtGt
maLdwdA37VLoCQFMEHnSk70UlclcWju27VTFrzz3vAM2REzi4oe/5/w05m6hqyRLPFgUXpv1N+Ew
9BALKM+ixaVzD30RqBSKU4h30VUUDj22HGZHqdzYoVaAd7rG7bCZrzIs8kNRhDqGhZliGxs1IYge
WM9R8fYo6bZ3T61ucT+WDeY7u+lLjEe87VJymQ5GAJ/4wtXUNQ7s0HLBl0OVV7yuGX3lsy8kBCNX
gJ4A7qFYE1KMxiF2oA9HChV2KQPAE+4bUX0IFGCvQ8mrHQYug+ZOV/W/UrgyvVuxdpY1RrExN4Rb
2JAxwnUJMlUelYiXfP8hYCvz8ZJvrnv++W0rT3COsm4GmfgyYKL+N/Btsx656kLQhXC5y8ebl7L5
W6FfrtmW5YMvZ5uRK64GoMzQghBf9zAT4mbiW6xIv9imlFXAUJkhgSnpGaSB+9FWlaT3VsKSsR4f
FMM6WuFDxhBpSxxSprAVhtkZ+g53NwS1SmUe4PUTRZuKfSsvEXqB/0ImGWFEBRA0NkfJwUd0blLl
gXAvjXn9jigeBv/mPv2pHs2eZQtWa62m5h3le6nY8zKTSsKryZ6aoS8n1KXNOMvKTb+n51qlOEKP
B9E0QUJVobf6lDSfLhSSBUPUWFt/DB4lqDkt7uvy+OKy+GFBoXtxVR01jOln+5u39mDRoxomlBDq
67iSYzn6AIVTS3+Z9ICXq+JR01THe0Bcpxa5w/GSipZbGKGyIvWn6P/aW90uaiyYJDT7z0oQH6JL
qfQzaKVJQRU6UJXHkDQBmzzjwlIHp4OogNPxegrxnJLA1wBS+Xbey6C0s1kn8WAKddfn1Pbxj9t9
d+Y38n+RfisLLf1E5TtpTP4lRsLooYGof7GSD/XGBU2tJBwX5YmTJkwO7h9ukty/wR6j4NK0MZV1
mDbuyEmJsCTSemBGlsnH0mluc0n5pqs4MQNGS3SC7zI+Y9OyoS6c0sJWH2GMRiALXkanxPxut3WZ
3m7OsjgZs59ZZ+xyPwTj2zTSrZFmdQWY7EIzwEwc6uNFtVO3XBWjqf7cO6dfKed8tlPMCZnb6CHV
OxR4oTrnrcWx5JS2rI3N7BmWtzDZZain/HMLAmjG4THcdsKv/oEPEdPLRDPSgnXtbXbG5aSGWyBG
FRZDZox2OTfYgSD/o7PZlP9GVZZetC0kJ4HlNgEgPR3DuLNZeliWV3NHJ6c0KgUiv6aoycDyGjsz
YgiEE6kXq1hRsOSvm61gfYGM96GA6GEo8XG3zEhJZ5DoYcUyTkHecvcH2fYJd7pEWtWmQAMNpw4F
BVbk/Wbu38vt9MjAybKMbeHRpYIJ7yD/NImjree1HISoucTCnL+wrPwEe32tWNdfrCQNLnHaX47U
FvwuTYl+l+pvFMMtOGwB3lvs6B7n2N4BYWRgpTZCrXD/B6kj90G6/T5xQmHmK6H+KdCqGKkd+1Pc
NigmGYJWdW+jaIyBIurFDuoC/vXXvwlnNKRKcPxByFP1NTU/JnPUvCP8Nhn8nZ+k28ValGjxa+bd
LkrcpilacG8Ce5rKx2YvLSlq8WkltbbLMu6hsdqtv4PU5BiZl+B2kghxRF/waEDBOhajihtUgOl5
CcLRAylKf+tIpd9t5ZNmaX2R5eVo+japIf0g2cw+HDhOfH4HY5zozff6ybre2Vz8/2HTO9VRmjWY
x5c/GEKMs8iuw5JMA4AjAGP6q2dF50JK3RRGch+fndI07XKUjTpoKDdgtAO/J/6gAmieMxW7QAVP
bFT8dQQ4gHLC557MNPRiWBWmLfAa4cB2Pz+8R0VxezpzmNd0pY2OSdJUCguOWTIexDGu6+MgWSL8
38x1AQqqFpVDeJhi5dUtj9F2/bHF3R8KLY67ib6/yGyjJx/aSwfNij2Hb0U0DRSsbls4j1JT58KG
sEUes4Gnvwae1YBfZlEp82yQOTOdHuZf4zT1p+HD0l770OYzXMJj+/omU86d8sLCyFCyFTC1VzLB
XAClxQ9KZn6pmRbsvmbww5zn/4HlZZUfcejvVPOVledaY68xzx9EgM6pARzNDYMpkklYwOrwGRhf
Ys/oDvxMg6mp6sKEIDk2vcfRCfscLbUz7KpaAYklFoHlzsub0YPby0aZxlrYLeigxkhVomYdIauI
Dg7wEJKtb/hGNrYPkEsH3uU5mWAOgmrEKVSsLYcObeU4uBbAcfDKk41JsWsUBXxVLPgroaCHoCBP
C+bkXAA3V06qgC1PwbKeXuO2EL5yah0BWVtxXsIJEucshuXT57FUaieCiSPDLNEpIHBd6TZuSSiE
NyFqpxzgDYUR0QZueR8t8Bc1LhOHlIUbZA/RjBIn3AbLVFHxZBRU9I4oOb9shWxOmkg2F4dxvd5Q
ufOUgV3YkDVf6zL/6b2poNJPrbQ7SYaG8fPf8krjZiG34iDsL1B75JNinVTJQwkgDniBnAY4ImoL
SlIyqxw5G0pJYlnyJDrHDyWA0rN9ngciVYonY/YC+bROQl6fORn4SHRzJxXNx6S7ALsrDA/bWfxa
qxQ/7nJ3IxyOaatL2GRvaNJ76LFSEH2UONalYHmPK3ETjdITVit18lNsWA0fFiKbkZWK3fmssOH4
ThOY6MObYIVnw9qh0On84f/dIemULHxIILwS2CqinVUec38fsdjNv4dbH0LgIK1dgh9EhuGQEj09
fgoY1G1evT6oS6Q//eIznuwHVRDKA3VHM/Oegd/NiSRiT8eS4Y3D+AuWqoUkHXVFod4cDauE5HRG
4/1jmwxcawFi5tr+uBaOfUNJDAANTALYLKYQUn4Txn8Jb0ptRboEPWgU0rAkBk7Lkl+aNaNjzUXG
LRHvNCqOJu9WHc5ClBxw74g9/6qEO5LsNXdcmhoZl1KIgylwcZRBvYnGfuwW5VkXvtHJ+Scwe6Wu
MarpYGaleA09xj3vaLOBOLAFFKFjbbLrkzj/R2DmtjGgmQYDkUTT1lnEB60cViC9OEjJ3RH3bdfk
cHQ+cV3563WcDGmFX7cOKYrSqQrSS6Z4hoICDlisW0WzyIGElZsd+HHRoly0q9gzj3bytmh1er5s
S83NaexeriZeLLG8I79l+uLZVB4HKLxTZgBbKQJMkoa5loVuQL/inJvv5pJLZ3D0xcmdH81B/ZZa
k0riyF57zgocRZGchBhzl1G7F69SUiFART85e6R+rJ0FYQNA3Lfy07tzyIEVgqoB/bm6OU2KzQvI
YT5VHNJ15eW6WoGk0tiSnik62WO/tdbUoh/uQ8XzQfLRo6emjXaGcBsDJjCWa+eQksqSj1ISJScv
2SMRWSho2CMgCw1KU8K24YXrEQ80Glcve/eTWnOzxeD7jdniDT5SGhKz3chjihtNzNAS97y5V2Ba
jPDjT1NhbC3SbxI1ahquljv9EKr9ukRgZDaJHHeseWetGuqUSdSIFXakhEso0dcvi6Ue1qRTGoXA
Ya7llcsS0K2E2EbIq0NiuKn9RwPsnrxMXEV/ruG+zmqXdM19AcwAcpTC5ZFcaa80V8QKbTX3rSX7
Q04XbEge68YgQzajMX20u2tX5C0KXCu4yRJW9hZMJIQT+YwLbRskRGflpInYx3pHALjIwqo3hot1
zXjTWpi9gaDb3FILWMsWCJx3l/9iZwmhKWDUqvTSZZNBNaz6LDJhC48zc8srp882w7pjXV0hafSd
zcNuv8RCyD61zrNVg4RpfpMTXHd1LS+5Vnx5xUutQJlRcBNLNRBxbRoHGAK3SPZt7ewCY1He9FUi
axKr3DzZ2P3e4aOlt9kuG1RU796AwVnT8tFJtvGBYwV8q2TR3sOhMPX98HcT6rAag3naoNm11fjD
ZwY9sBofl0ywMEjCAMOhor3F2Cf9m71/+NQr+ua2tyxEUw1uGX5CfRbPtUfH95+oqa17X7vEPbbh
TomLZgPNJ6YHITNiLQ0o0jk9k+M/tGjA3jFRE7Wfb8CEiYG3oEbLcehaaX0tWVFU2FGbGV/5Kqwm
n+t+WGDbLhfMpqwqLj9RLhuJYNlAiZ/HeplURvi6TdbMs3I7B5sgOfEuGbfDTkMDzpYo4dq3vL12
xmprlKBRsz2KnTiXniwM1xHmCw3aupzKsdzWgGVBVwOhGt+0BnZ9O9qzZFGy79eCx5T3lv9QsIBw
RXfcLxjA04g2GVOszxzjpstIrzYpJtfj5x0CYd6EXjiKrNgk9bZ0APGl8w+wXNBwri7vbhYiYlKz
QbohyJwxks0pGk0UWiNc83ocdyXWCXwS2SK5hQhTRtsXyTq21UyDGzXphq4wXWrUueiglOsORzME
lR+U/hnDiPzJvpAbcaCZtLuTsP8XpBB16Gv1Wt+zRWQIQLa2n0yNwPJc0C3urUjUiipe/XgDVO6j
Zuq3IEaBTK1WI8C2M0GnGIwnq/rgWKfa3Yw3mJLKC8AULTYvmXj3+e/vTyRW/7ASwlYuhT4jstW7
CxtnKFDfh60/p52AltXacvg/s+KI1CoNPmTPJvgl1rdvDJwrtI0j0AgjoEH1cxLEP2aj0tjpckoL
G6N5yCKpjaxqPeHuSJhw5dF6g+AhRVzHe76F0ORfKKgjAhdANNVaQRK+3hdUyNaqmEOC/1M3PjTN
4S/ucasmIzynB59Z7vz5RVXZx436YKnHgpSL8hV5w9XZoh5/N4GyzmLe9eI3ijh3I0XpDhXhbmm4
NVN++EYd8V+OaY0xUyFZDZRxA0W/l5jdeYF4lo1ICWaH3aGN9kjQ9Z2a1n3/atrQSP0Wro+Cdzyn
GgQzD2VfHV3pKrv2oEEPUO3DeCGb214mBTjF17R1X8s2u5YRj7w0n2L5TwWCUY5HF8pPv9EMMQej
Sd/DK4TaqgqMr1y7lQhAlanihwWN8apkUPwS2WNCH8qC14/a+0QAnZxRbqIgWqf3N+7xLKvv5+U7
FEdSlsi0kdb1PuGJkCQZSMB1OPjZmQWqC+tivwtQmPfkwnie52lwDUADpDRmjT7YU1ZbtKKf6LCI
/pxsCgH+fIQlh9UBQ3Mn+Xjw3ZHOVTLpbbazXzoLk+TNyhENwknajYiAR3CvC4oSTusah5fm9PDD
1jZuCcgkcTcfQrkjIsV5wYqywmN4Ts8yVUBQO63TDmOI1uEmo5Mgi1MC8ifN78bZisK/LS8zAvdW
kDX+xzC9/gsrLWpm/X5DPOiFcwF8N6cg94srWFCw4txALF94ZiBUY+uHH0UGj4/wnmBS+HW/sbY6
DH8zvHgUAlokf1kpbRvhtkntcXBxUB6+MJKRqjPGupQ4jULOYGifj3jxbm0uvWY1U+jsaALy1c1/
V5fXbqBfXB27oPM7segoTraQDLmv9dD8cV6YwOCvNeJfjT48AfwWLmQr4dQ8ZQY5zpVAWZeKU9VJ
mCKBh8oDphH8AVFn1X8HnniBG+kv1kJTy8Xvuy0RMrgjFCZP84AdNW1MU2j65bpLPITJtM3J0z14
k1UTZZu3t7OXSO5oaeoL7IETz314rudmek0KI06Lp9eVpZKcYhN0KnmExxFKtNVNkUbH0oW6AqHR
RFsQHzY0d5DeNSRDjt6mwvclOrvp63hSxG/UMPuJK+7e9iXRiW9rXMRLJsO4s1GyQphX4fl703f9
bXdGzVNizXGjEo8XoISoDmYzTb8q/0/pLXvB6Q320GZC1efAGVdhqlhtCz7XdCzV4JTTPU/xzRNm
Tu1ue0B42j+wBQk9PH9VwDgcNtSPmlxN+SON1HIvJtfOfFr9CIdHZQa3ISOiwlZDF7CDwxCs1eMW
RpUAp8qmfj8nM5Hx4ela7flr7fxMM7zgBF46TUzl/3TZxVC30g7zyzqDvQcuSqkYx39kPGj/3LBN
uXNuhZr8laSTML7IDHVLlY30K2shCKhPJXkekKk6iCf7hMXQmtrRaDAeDbx7Xv+C8H7oxDFmygG9
cKXk77ExRJxjzQvFd9QU7CjgjS3UMKrR2riOiBGTn9rR0uL5qqeWumHkk8wCfg69vmkEgRyaXSWl
uD3VTIf77VviFojwM5jSRXUzAOUtUNMwBQTiguO2LdvErx22FrdaxYOZPdKbSO2i25paimdPvseu
XgzRqNoVvSat9aYYVIG0SwJfCWswfTaomXpp/SuzLMZKHgHZc8f9C7s0ylyRZj9hsby+IIWFs0eu
wApg8E0AFl3KpUS1FgueavfAsZt1Z1cG1YAOCuYv9nE/dFSS0gu+xoEUhYLoYLpD8JisVbA1VhSA
RUmGguiN4ZY86Vv3H/MNPohG8eG6NWxN5gP3wrNG9Ma9aqrqWbaFJ/bwpSzTjMySIY/ej62J5XDy
PkHbYYcJ6lgnDamIRMR34CZe7YpW1caA5cSGEDMAO1i5ItjKX/dzRMqOyWCJm6gPYYmJ4L/IFVXo
ADOwHbEM17DfTTWf1yTEQXtQQm3mswyHn0kizpCHCzIrnHtGrOtCo8e+vAXzfmhMRa40c51l0rNt
S4FE6Ig+LshwMUwVJAQJC04soV5Q2AvfWlegKrBjFLHiaI7QOQlXU+FVEJD2X4z0rliTaBerW1FL
RunN9xX2dJIlryFWzxea4EJGp5R+gbiZjkGkwz1EPUK7tBSoGhUmHOX6q8buHQnOJ6148+vzjluF
lafM4c2mTpML96rxxzgv57s9NddcZNhq7BkmDTGYZXTWCrppM3BaMbVzxB/7eNBy5Y/FPW4Z6sYl
ygYxshCcXk0aCtojacV6V7QRo5QSyc2CdnGbIyx4qZmfa5O/N8Jp4NIByqGZFDtQeq30XS+WRc8f
FhsihymgYfk4KKEn8eRJ4gwCfOjh9pdZzSw6Rhwp6pLeFFk5mjTKky9lk0ts0S1kMPodwEWi6byD
mqaQSKsIptApRp9UE8D/IclKSbAjvyzEP1zGurkW/GI1CHatz9avGaN85xP9McxljvZg0kfvmRh0
CCVxuf7myaNlrnQsGsMi7l1W1b0lbAgUyK7GG3485Uev+ezVCDTKOpIHmBStdA07jw/5yb+qb8cb
Nh1sPHzyH5c9oKdQ97DtV17T02LI8Rg7VvVq5NGFX8RHd7Rv0RGxCFP4u4AauNYOmI8tJo+KTmKo
OfGSP1021tGsNvLxAYiwf6U1oTAbV5dDwJEmwCJU4WqdYVw+S+lxf7OQ/nCaCfXziy41PJKvQ9UL
/NiQih7cCJFnh3AiPtj/DYxqAXWfVBz0suJ2hyUIznCkRZ86Me7+h6qmZ8AHmvZdjuSWFrfk6rjt
bzQG+tIrMVop8+Snp4+JwRyPlYutLFIS7aPGZlA6iHFUp424CfwiDQp587aTN0PVGTK/zxin05nt
BmRxxWXu1QB3tlOH6yMNFh3PJIv3Hb0fCecCDq2nZa15NFfh2Eb0eVp6LOz6nqfqwzcpbGve3rYn
17kWVANO7T867+xxmjB+MtCX1yIv4EZran8cuVc23bClsWEpCwMo+2KF1My+DkaQIuZ3xRJL4HAF
1QfcwZu/+r5Ga+jqJkxLR5va4M/xanRUl/l+ndy2cZ0B7Ahrh2xZqAePTkQHZYobDrykj4eLiBQC
gZNtbngA0zz6Q7iRLs260sYPhUc3N6Wis5ZsHB2lH9sLk6Jwcex2hk7TwmngkVUfcJHE9DrIG9Vh
82ZgMlYghw4M0DrUly0wxkw86ak1WnItNF8H7xUPq7L83Cwj8Vw86VPLZ/ru0dQ8MrTbIg5ZFgQX
3xceEXrtKRYdhU8koGGdK0WAXmQL/CxcMpgsRjmfz9y7ytiOJlb7Ma8prkR4lnzF3VgBWmAGCUGW
r8b8f1QoKQJpkptKesC1kKH7rhl8F6Xff3Me/ZDNJJ3fj9G1BlF57oVibaD1yEwYuU18Mss24ozm
LFTZn3MkD5qnrlMLTAidlgaNR+hXcGpXSOwhRDr6qSi2o3w8xK/5Iqk80r6+o1829fA+BVS/jn7d
STskCpj8rXVnJQUZSZeffkQaAgc0u4VZFWGR0J/iM124ZWH3sYI1Ewz0dJ9l6VBazUW4hhUikj9d
N1borrCxKLznj+yLbfz+5d2ZbwNccIj4L9skPdgNBF2MCuXH9PG9PXhtG3OjXFm+i5O+dwq7mI1J
2diVd3HwiTZkXyN5VSuxA0KqRdQa8jZel8VqxGVjAq+/y+CI8NI7ugCNLzY37g7b+XoLQ0M62K1Y
Q3lirNLcFVZW9+3Z29D64e9YzOXpDZf3+g0ttToC8Q8MDGxMPk9Go3Pr4tS5MfiFjx+PAcJPD6Hd
pGLedACUbuHiAcbPP5jys90anIcGF3HX6aJnI1X8IHxFzcmUxahYytz+8jZc6ZSVMokNop1WMprk
F+lHehyjbtU9XG4+fJfOBt6oPByhkfFtWf+e34ZyfpByaqr+t9UX/UuqB3xy9eNSUeBCSHjIev7r
NM8ZAf1oyTEJqvqQFKVCrApVaTREkA+/gfbOkO7iHOPik+/SRNqZcO7uMgS/gZlJ4BSV1Ru0uBcw
naAARLKRqwBHpeL2H5dCrnLv6nllv857DgN31+IX/oATJfmB6SQxvUkLSA9nKTlEgjh91vfRIGWt
/Jkpx981jokWDkTDO+ya2FYxJb9pvE7p4iMsmxyBbOty95f6Gip5YD7UD5lbuFQvRjQASO/hIsd8
YNt+er0ojL6H9pv+tbYogEriJ4ZU2RhyDeV7HC/grXmS7h5oIa4ImH6OQ15XuFKWIPdm15dLc3Lz
VmyfjMsa/P7OJVk1ktSXitDXvdopfHhMVutiqN0/WvqvdXFmZEpJspWrX3nEx1vWeTZqbqBq+oup
G87n+iAbwCsUvmErnbeZYhE12f7NN9pJMZ7MbRazP5ofolL5VBfi57OVAauRqOkLCzSyoWbD5Hjt
+86n2ywxk+7WDiCzcsQBYkedfTHKb9b5KQKWqgc04sAi63/QYDfzx7ZJyiUWUhnVRUgL+TF3PEX1
HJupycAH32HdRLTAX3K5AHXFBBFRPQwMIW40TKFpzxQNf6ITw/CP+58n7Ww4GT/YT1Tv3OB3gxG/
RXBUc/TjAQkxcIIVKhoLiggxjVYcnhRQI6Z+A8G7VJ37TYPlnMu3EJdxgUCUqEZxEGEN+Y0ONmSE
CDm0OgrQwVlYe4m0b+RBFLpwlsARJxi9ops5Yv8kdReFCDAy5L+tyqej92mdnRU24KOjuc/NCZBw
r5n4JPpcP4rMB1QqN6KkR9IqBlaXEGPWOGdqYJ2BxS6xWJ4Upk1mP1ZOijxTj3IoAFbCpCTjyVdG
BU7iM73W0LKAsX2mv3M6lti4JC4LZUbPYJe+SnKqkwBpSS3ciNb8i3Ou3zkWNv2Bf2Wrw0/UXh8e
yDZ92Ypko2FQd9F9ML8/PnBJFvSW4bz9YHFVnOU/faMiuHMzltrfEFM9mUcwNbGnXsEFtUdJ3VYz
lH6tVlu/aOuwvTOpR+t3GkttcVl9hVXo6ZLQ3OJ09ne2u2H+3D5Gfn4feYE3VZFDy0W2PEP17NAC
SgHlh0Zxpde4RkPtHz21D08XuEQ26S8Z+z5s2Sjb+QObfxbt91FcAoOjC1qoGpAR7EiZ6+HSaluK
14VvNv3gf1cqUETmf6l6V1w24l16XLFO7bQMhEFiSGdCq4Sg840Q4DsGPkeQgwdpVIAmwcN37czc
PG2+hR4ZSOS307/yHkOH/9YspXPszxTZXWO4HMaFJSIh3dLSTJkaVCkMRtecg5x5KfW49GrdQARJ
0aHw96brQQdvcedgsbqLoyyuLao4ONs/d74t15hVB63uK4+L2UPngOF66JA9d12CRQ5uf74Sp6gt
ncSvqKP3odwjs5muf786n5ET1+QqDPZJl+7/Yoayz3EDS4+TJFkx5/6Qlbb99+r+z9+nJCURV1mH
c8TIYfLGgw3w7I/eOpjvpb9rIdeRHshIDBJGAnW5QnNVHoHYNKUaPCL2epI9zUf+7iApWFQFspAw
rrgf7sOgBJnhrMzPD8kuizjCcm68NkbYRtno0Vhe30AJsEXuKMDrgVl4+81btwkCJKe7PLN31MlF
kLJE0UeANory+ke539yfbzm9/Hn1r49GcmxaI6Oik8dF2IjlB+nmx6c7zk2vKdvSXnMfjzRJLQsN
QDh8OZadMvSCKDPM5kOOVj/DZrlXXWHFWC9xE0XCPUbPGffaJ2eOIGTHgjVge/LQ7f6JW7ZolmXI
QP5YUlUm5lfF77qH8KCEj0wbbh3UcKBqbH+CJl5A/JxKo9Cwhuqz8fpTsAlrSnVgosOKKLw6KSB+
NR+p6sd5kVvI7HS39rltXemj3hZpSiVqkuSVJjbjBj5BptqlCs7pQHtrPQWGc0o4P4J8hFMEVBoX
8jKCxAKzsyZt8EAOuNBn17HFXbVYhiIECalTPaVKAJOVcgTBRxv+vly3PzrXZ1rSOtEr67BRG6q2
yn+JuRh6oMmTAUXPl/GUWqRJMmVF4OKmwZptLrIlOEN+DgLzM+n3S1q1cafmtiXHDlY6efnAufml
kz0ROcI0cT1PpVSTwxeFaTaUR4T9MdCGCldOFMfQD3WGRsyNL8ZHSATDPk/iXVUGbH6H9886LZ2q
B0SaE6ZJaAraALxOtX8Co+9c8YoiENs+LQ9VW5lOUk/+RsAYgF2zQfg1htAoIdfSbqkS+mXbnyal
9m6yP2ZAS+dXJK88O76lTQmyUlYnIxue6Cn+VYQXpZ2lsllSt060fJdzzccTv6umVcB9cxf3jxcH
yBFa+xNZ/wgbf4iEYzMVk2ecwavmD7LV+wS7TxIiHXMn6kt3XTPzExU8UdBs87FIj5+j6suxt/D1
T5GCFzHCIIH92Rt2PXer5QUsV88tL9wgkaTGiScyuvf8x8Ge2M76LVtiGTgmP9hpyAdQeKNYAKzH
M9F1SBjGS3dhDkpHr/yRD4r1Cy84RkWvtLH//q25/e+VylA+Fs8mYCHoFu1dR0LO4360GZP9F5mn
rBY0wNFo2OxfyAPqfdi9fii9/obm2u4W+8EmtH4j/8VOeqSd9un5HAhIWyVppvJ+5JNYqCQKdagE
9EyttfmfnkVsBLjN0QhXxkU04LWsjD72Z1Xhzy/UR2G51LCnX3As5x6yhoEiBPqyMK0eT6oMCYq4
yMSYOXY7OeFTr6yP/KFiHvGGPg9osgSrXB7oOGMOEow/Kk0u4kriLKPgxus4thkCXNGa0buqUO55
Zq6QX9b+fnhH3uGhW/tyQ2CNlGzDxA/lDF6jcTftli3+v3WvUOyRpLeYTJoZ119vjrZb+aImNVep
GM8d8u/0cTjJN9WKzLqcHujmnPJxxMmkrclPSGvRH5LO088kL3kxgEbmj5Zx+GiDDO9b0raXVC9m
YCQU70GyBqrM0AREj8zsbbEPsGB3JhVaXX5MpubhoryfNJR81igFteFgmJrUEObEQ1uyUgx5Qybj
O0iICKxweqmXAlf+qdd7PLzyQZdgLvoz85ATohhgRrPXKwcSbxaY8tGo9gIcBQ13taJpxV6zGbz7
YlTUBTfKn6fJCNuAl+ZcXLLSfE+9ttMovRyNbmu59/K57NYneQS7lC6P/qP6q307yUW5E4gXBHzW
FeVr51TfMF0vT+U9sp7pJaVgtCj6+qEw6/2GsgFkn8fMvvyhXztcFXXbElOn9Pck6K24dgs/Sk5e
SEUYXGCQCgvtP7xjjauWVI5J9m5f/GIhleYrp96bAnRx/RtUEv5XmjEB8bjKW7mo5YMnmdeESlZg
e+aYl0NpF3x/ugvcEdRnf5P+fz8rz4VaRXSMIa9es0swNBkk9RAG71rbfdumL77os57RGkmVNGJ5
m5VAAxiX09C+qWYqcAqsi93+2NzhX9aCVfMaa8IxcxkVdkgPhrbk/7px4ty0bqQEvtVpH4exKHtO
eh5x1N+Wtbauu+oXhvS8cldWbJBBZJWTHJj0vyD+gh2DO/mUFg2OIe6FvhXxonMza9XBvXJ3uIVD
aKolMSOP/Or9HI+fxmsSXiubdcI1ggNm38jRa37vCCC04PIMU3TQoSI8CDiqiYkZLLjlIYyJe9X7
TkxldsFsEG4h5NISosVYufzR6V9B/uUNXw8FbOcyV/deQeZtih6vxKogv6zrbey+zpvPY8vd/tja
wIfkw8Z7Jptm7PB0l9B8n91SF/BDkGgEpMSBFKIjOxC+o9ZTDqz13CmDqA2fSLngi+ROqMsouuTI
t10PVnc3w+GrXlO7l6wg93pYF5dYb+KrlGsjeo3dCnDQcBnWhF4HlVZgFUccVmHD0b/KI3MByrIj
mzCKxsASZal0dleZpK5k+eAjA/xBZ6l+xkitS4vGEyJuk8UyrYTd4XKkGTVa9jdp5lOcr5c502aA
kYZy2EBEndOs7tbcklYFyUDCWR0/i+EjKIKfyWFnZ/K95UH4BTboJrd4OXq/0MmbVNdK11WDhRsy
8/tW9HuHhOSDMEHgd/rvOAPZCa0OPzpvMvWeKMWXye8nVUnkWOeIiMBD2i/aNCWI4jhhADotTzQ9
lxK6mYA/xbF88HeQDVjlU3NPGKEvUsmAAaXg52TmYMRBXkh6ikgjopCWEVAWZCz8PGHsESw6JY1p
pCgMSCPmrc6n1dXvhfNPSuHXHgxu92AB8a7QovM9sARC0RciFAxPLYhuqMunyuclHQ7O1XY9g3MX
PKZnD0KzAN1XOVsS/Oe5VFZXMxrCoYKfPgfxuLdh8D35CZi8JlJ7YtbrAoRXgbjmU2cP7GfWS7Wl
o7k6qxcVF1b0LJk5rwclipNq7O9QDZF0r+Ej6cyY1X4b22U2Aorqp5HW52t9SerTFJItbQz4w7zs
5HTSd40c/Jit94+gLZkMhXhp9bmN30PYfZ30ABlChZ1QJ6RT5D3jdy5y+2yjjLMhCeGqxPm6V0r4
/ASbyxm96WH4OgbP5AICECqArR4UWn73aN4o91IuWyNsoNCnLoz7yCQUneqxgWvDI835iX/b0mgD
cHWkDFcjtfyTgw/PAxreGWmJStrq4I+e6JxMxj2IIhhiy0CmteWV7dMbab3NIvkTQR/E12zFgmdw
DnDKNzi3fj6dWYFdt+GSG4fywemoxb6DGGQavnfoVQXn6WulgzV2+TWrNohKxKM0W3zOBTQzAnjd
tOqcyK2Z6/a8OQhfzk2Osjm9D779okLVHAIx/TbS1qkmiT08HNmiW2vrQPMjIH6NzhgcVfDaP/pT
ma3w9ht3BIET0hcjlo00ndm68h0eBUxUTRkedsPr26RMjim1K9Y3ew6b3LvHhI3G4KP8pwdFzRew
Orlz+u77/jCDTxMKZAMQf/zbW4aCFLE+UUqdH2Oi4ET+3Bfb/haEe9N/Kd4ysfjzl/5Gl/GALvIr
p7DuqONwxoEhcmW/dDTowq06qTqsAKUgA4TxE215Gg/b9KKTQWdrd3M1lAbOP7i6st3EuwRRfPHk
rHILQxnHxI7yVFMXdXE4bB6KybqffDKsTgq5S3QvmdbuTOlG7xCcn+/T7IkoOHTnixJogVsxzY9Y
QcezE6XLgose7tTMU4dheYHff+TBH3/buoizs4Gcxd+drE1dAeQejZkjx1TYTt9ggP4VXG8zQ2Bb
SNky7Q7eymIa2bihMdcCRwF/6CLKjn5FM0zn8j2mqRJ5F2BMeu7Uuv3qgQF+VGJ4eAFev91FpEiB
wEiWEBdiQfI4cy4tU40Orcth3NBhXlIOty8Y5opgpU4hYmnBacQ2Ay/EsmZ+RVkvD8OpkPY6bhsw
pJMUoOqF+rynk4qqbaDdlZHkNlZjoRZQyxc6KxHkOdOpMgNtVYOIwoOF/goNLejuBORr5up6BZKq
9YRN3WeKCLsxjETI7SxfIITkxR+DxV+0nvziqer17EUW9wrhB7ZoJd5FIzQ7UEBPZvV6Ge0bKKcX
MtBpKr0Zr65G/t0i7N0YeZ0cwIXFbvmUOelDp41yIWzaAMa2K3r+OZsS5Ku+MPmjag5a6a5mldFr
mSKHXlaORes20hUM0ob2gwuEGGx6Ir1OGnGhrGnwXcJ5E4172G/nKZOtEae53bu1Lf8UYfX123cM
4BollqOTnfUtq4hCWRoe96Da5F9AZ1mloBc/vlonm/skT7MvfFxVtYHgbcBdoAAdRjw1PLoWPSCI
ho7TJ6osEo/+1wYhzkEv91sNtDpe+vwH5z7aBu/1qwf25rKgRCO0ukvIncIQoXbzZWjMqliSYJpY
O6tmkWjmA3O+N72ZO6r4UQF7q3XJVUy+got6S6UqbspM/QKdEmqhBjN7a8SpuMBlcrRIYzsxC14y
3A9gJR/lVKqkJjdkXjScwfxUBbwgB5130uYCh/K9ajkcSvkNk/wPLZJz2RWIdgJrFspk0Pwh0e5/
Zd0fR0YoBpPwp+xdCOdzh1WRHRscAhsENhagA44VKJcKB8ZNhSfnKJuiVbwyAPTzGUSHOfU2xvn3
w3xEAbtVSiJZMa3BSCpIP++bRvFJj/YxV3q+xBZxp9QdUmGXy1DNmy03S6P4ewwaAiVrAzM+cxyI
/wAsbW8teLHqAGU2zHMqZaqZMGXXs4ptk3kSotyb+2FKr+0T8pFTFqp/V3T4GHVhR5JmCjwcc7wJ
K0qEJlycdVqd6oC/M4l5h1b63H3uY3m7aYT14X0NZHjNiG/KFtTQXIdwQPMVtUyMr99Dl2yQRJUv
znR95Q8PvoDP9ohqHatjVW5MxxkSyIIfBcWi824zg5JKdkw5FLwf2UvwLZYgG1v3WyiACWmk4DON
0GKMC/TUp69Dud6BtMT2VMxEWRc0fFnqX4Y3Sz0IoszOUZYtlOVAe0my1SKDqdCssO3yycgDxdUD
Sg6FDhduRLipZOtvE2d9tbhMKs4m8ho+oKUfC3b4Cj/7/6qdXDycizWvTAj5+75ZYgJFk27ygQC+
HXPOvsWAWi+u6E5wrfjJ1rFlPkL3aOiDGE/27wh0LUg2Ik4I2MALsIlwyR5j8KBoJjU55VPfkllv
MqvWqQVmX4xaexBfU8RYIqyJrDdFq5MPP50jKrHEft60MkzmevDqpJl7CzuOK/14yrEP93KryAnD
ZuiHK292ilEOlf2YQ0BMQ3wr1mCXHYw1n3XKXuN0oERJ2Po9UgWT72H/C8hKCMr0bwW7nkljh4wx
NTUuC8h3Kh8tXP80OnK/WbWvVsLN577PycY3i3gJRODX8RFm/AIibhhusajN6fdDqLebFd4PQAV8
+eSD5ImYQj1jRYsAbbUGfleQKtXt528jsNRGo0Q8rvBEk/3TLiAocSVoFSzc+lR/oH5KSYHjQ49j
M7F7MXtApBsr2Y+Ean8cSQOZ5pEVpIvNyqwxsm/7epiMDNf9EXDanPDfEHz8coEuxxRWIq408SwK
vLHhnQpaufpw6hNnUrxYuO+aIPHTWknMEY/ixuTPOXFO8YE3l6G9RMZGdn8ufdMZwR8r3i6qhIxQ
RWmqz1s0SwY/JDKOCGtDYwQXNroEi3nNDKyIGruAASMzQzUc78tKjRu+MObQnZLoHic3xXPImnKC
6WMlhd62gzWDuIp8IpwGYT38b24UT+3mF/yOygUijfCObwTACg8YUo2jijXbYEogM3NGi1fhTDHp
8lp3q3RCq7hlUiaq5A9gtlt6/fn0LBzOScOhKcI2uzerfxH/leA2cQuUeZuAwkJaXZpP+uxNaffQ
EYAfUu8fJ3svw+oTpQKB6A3P2quCu/5ysiEqIhN374CXSUZqwkgUMLr+iEj1sCNz+Y3eBxZCaVK0
m5GJs8Yh1we1r39QX+K89AjLAeVEtBFLj9XNpwGktd97SPXMGvTEVqXZRyMjTSFKjnhZhUWOhzRP
6yAt9AlZMDBtfwES6mLlL2cQjkkR48MpnT6aOfG0lZ1snk0QNFniwAM2Heu9EZj4ptV9qwUat9KD
SsaaMvV9n660XsESz+gST0ovyV2v5v4rv/PU3x2Zj75rVrwD5y3KhaNaAEWhH1v4La2eNSeZZkYc
e0GW7vaKzpDC9AWsncRFbDKNs+uvB0vlQyRbTKM+R4O5YyrC53whN21k/7thJeaaRt5l2of68DfP
kvBJmb/e2sblqOs2uZgnPyorurFPqM/OuV0moLb4zIHzdiNqHP3g/hJl7z71AL70UGgl8yJDx0Uh
Nnq7bMVA4rfAeVjjNsXwrNB85NNluRRKfE7s6Jrzd9YoNafsfADgLA8j+79DFkqsXg0tif6mtsnc
tPhKdlSnANWZz9CudJGrXwzDJdTvMn8tCP6pFMQvS+Zlu+Ip6So9Fv3nmP8gyf5bA5lbjyU8OqBN
clYdmkagP+slQi/eRaq32fernvjvEVX3P5s9wAP9OPR/x8DofqUMMD1WIymfoBFYck6hROYih97l
OK482PeSMZd3v7wX4YGPSNxG/tu6k6MER2/VQxCF7ioKD+zT2M3hL+M+ThApfZKBlbnAFQLDHC1c
XA2eYYACRiviKK0j6WCwm9WKtaaw+YUpzDAONZOFKpOTqsYLFoDV1toltU61cnCRQL5Q6XjFu+TP
xEcklkXe0lmLi77QtpkvTxsm+QqA4pXHyWCBCtbfvu/ZbL/cmlevqNYHGT4hiC5qCNspHHwJV3LL
CuyMdRn2euQ7gOXA4t75GraBdDMQUvFehvphBRblhtzEr1MAin8GaEJQhjpCYRB0vw3DgPJnxLzZ
a1MTn17LdaR9TKEhkqYHb8u8A+ucBcpLOKM6EU9bv3GEy3ivK4VshyhxgDqVG/uMc9kjYIiH32Qx
7EdVEGWIIEOuIRoiGRzi4VBPMWs4BUQuN1CE5yI0VvrncdrpXX1Mw1JsH96uaCbSKX+ee1I/n0Jo
dtOxZt+8k9UKcZ7iZLHTyufqy3XXtHkpYOWybFEmBe2eHokOIfowWwJMfQhE/KQM+TnTPaf4nMYP
MJav5x6g5tJlcjbypcZdTltGORKkF5IXRvqiTzAyeGwfDKDcqNFzvGVfyMjWhk7bCkVDnKU9b573
buHRWRM2L2swSZ2Svjc7yKRKYVGHPyJyFnLZnFavTKeHcBH0Mg0gM13/lEfD4n+hrNJIM9vOwtgf
cJmy+Hkzi0vgzOZjd3/A4Uc4raLD8tdlH82yq8tKfzFty5t2SfmjRbaE5f7q4Y+boY/cIVDZ/vra
IyMWzbuu740qrVbpTV2eqDv/8oh0oRKJ6/5Z/o86FEc1L9dqrxQcKc4s/HM3SCdFgh6OVDYsmSuS
HtR7mJ9Q54F2o8vJ7FSKPXULRsNHhQca2G8UCfHrzhzlZD5VrY4yT53RCLmG9awIsiupuliCPpLc
NOGdYAVjv8e8Rdfx6JXbZnIlDYePAkAH3x5yHCrqCNVyzrm17JHBua1BWc2K+E8db9sessBXeJ9t
M8giwIuCutocFm9bHDtiGaXjcNSe7BnaKz0M74ybCCZbD8yW+bUH857TWlIvCqlAFBJL8Vwnf4M/
MWcBIp7dRIMWwOzt1NXUWY7LGVzahNwnshwkbt4bdNAuxK14obQ128tOGfFK4iTjGIX25DZp+25v
9tGTJFmKnbbVvrfK4+lPJD3pv8GGByp9WiFaN+4sgHUnThkt44NG94yPWqDKwUFrhBwW89AQr3vR
GdsNdxHplPkYRfV1Fev4Eiwsxv2oVdnA73JhJf2r6CVSPQFa8OgLLt5jfCv38Rw5I6AGlXQX5seR
Rx4EEhNFHAIxppfQVjIs6d85Lsr9jvye4TYMUwutPhOLQnKu4Mnnxj2id7eD4BamJa7/mETTCoMN
NF+B/JT9wQtnnEvU0vI+gk5niiPl4X7HpnMtZVcVzf2rK8/Kflp+PeAq7ALgKvb4gjh+kqFJRe0a
P3DkVPzLGMfyLDi7dWsSrIhJJRnb5uoi6XSR4W3eW4rUpu5SzOd7Gh/t21Q1pZtw8RlgOnWDEUQS
FBEOij4CSkX4LCiAa37WSdvaeRus9ByybIeqxFw3UJctgt6rjYOg+ClOJZCktSPOOrJnaNv5ZMRt
Mh1i2UadW+3tDBclRmDC4FfC/ed989FCzIWBkj25hO4TsBGxjcwKpeG4o4E/cxUWeAHGl71kwpez
7dT5KSwQA4XrscZ4JTO82xxRnB0JQ+CMjkeen/M9kIj9J1JX/AehPS5eH1TrfBFQwQ8B0X42q8/r
o/cLh2vyJ99L7hbkZlx3k4AAmvO+KQ8RbdQV8eJ9jBWyL6BoEHN/zwfv3uMWXq5lt+3/rnDJuage
Xciq1Y6wU494f3NpANrseo+aXm/D1z0xm8caSdOV0wz4rZLHwhpz2OEnUMQrzDbNHIsDhBMmUpwJ
PxiqrrNjJYBLjMVj+d/xYYXmFM5oDtD52MlwEn3pQx3z6mXbfHjEe6v94JG8cI3rAcTZpbzqSxYM
8NKV4/SbKLb5Yw3mnyv8fcJ6nkUDG0yiNIgNsbb/Kd6ehVejHg5QYWcKdLryN+4ANg/43BWhAGnl
qUaVexszN66yPYUst6jBN6LNO4yJiEuTJlppqwkzYJ/K7voxHH7AaGn4C6S0ferh4p+4YfelmBHl
0d5CzuPHYpJEJgHPvd+kgsCYPlxkTeCM5sb2FU1Y4rHI2wRf9DVfCmaSu+kP6o28D8R9D9CuZ5Gf
JF4pFB5FuA/4AIublntwXKaTjO0ma5ewJtz0xlXC++MvDYzCW2LCWKmRVysAmQii7rOLA82L7/MQ
rSlt3EO3xtwExVgZ74sI9cMDXkbgALl5Aa6wFcLysfr623grQyWmKt9MBtrooa4s01w5c2DjVJdQ
LFCunNB8GD/tjaWAZzRItJ2yBACG2wsYlwt+DtH9JGU9Mw3S4Vow6J77h226WkhEfY4zWNe2pUoi
pQXx/BNStmv2elIkmynd4DS+Wt/2jFYMVx2462kodytFdcRXzD1fJ+sMu4hgNPreA8QXz0Spvt8S
Pmf7Fk5UqMRTNk8oSlWbBeJadmwaGAwN3RX3B53CiROnH84bcidp7vDJj6Sg0IWo8B/OQJyW438N
tFxHyn7SpeMDdfiYE7ccgGCkSBjRAuEwWyGFVnYtJIEkiI/F5UaHs1Wkzg+bQPrDPZp9o+hb1KRt
yRTk5sCHJTS0Qe1M25XDGVhXEglh6S8BT1y+NjOehWi+NC7rBSCKVv93bGMQCJKkH4ieG+TUNNbb
WEldJmogaSQGZ2XexQkVGICfV0BqA4gJkXroJQtajRHhv+oZE022mDN/VpE27HzlQPttro9GxCVT
3bQlG53rZYtbtk6i1ceKQbgxNZMVQZ+uWX7976w1AC9QqzdrLFK2THF8Hr8rKXAZyOc0VZm0FCoD
xoh1TUE3V0OOgtN48VjsHQ+fHPYP4X9W0+WWOTSqjY2iMFvy2LUmXfBJPsw2Vi5RM2ckxuAATBOl
f5HI6uQgkUiQmHC0k/UNG+1VRiA8prvhzmeFfB68mgp3dpDxEvSf0CobW1UhUniiPb94wQ+S6xEN
hEJ3ebkkSDBVsWAxyYuiabEuNnSD8YobCqFkJvnTyDTnamPKFMeL/27uYDlovae9+s8AFYRzEhjG
pb2Usu3pSn5M1TfH8PvYb5DfR1jkek7cq7FqH+a8tfejupDKVoqBjbrr02qKsWG0u3la9tSlxTGk
WFfI+vKhRWKyfG2Q9mU0QysaN0qAqd2ptw7Zf7k3eEKwFIeTaWttUQUJmnUlCmIZFzlyOLvuO27d
gsp0jWemS6zFzFqz0pkwIIYDRYzttTKkuEy2QrTIuX7F/vO7rKvCYRyFX/7xTwB7GndvpD4jmrWu
mbL2FBy4hKVNv/u7bWZyOGNWkujoMqrIQACSFeR58x9N++cg9ELRS4cxJJILyx31NyxPC/rbTjsC
HviKPF4mifF3y2nN0xhE60oyPu1A1sBOlRmFv3OMqMJoBOkhBjt5O5ku+HnfNe5qA5UPc2kjSljV
hHg9xRhKaVSbX0l0gP4I+EUUkRaVLzw747xfGImuYbdRJQBxVvrR4T1vCzMU4eNwQ/xUynHw3EUG
IbxjNEKZbxbfb8HDxxPrLg8ADGiByYrbkbpWfjSZdasl+p+ai9Sjz9NVqhPEf4t57p9CqM/+HGU3
yX+XtLWvDXhzNFOg4N9lxBhEYh0pBL6WxnqzP/2czNxio7A+Oe77PYoz6keb2dLqt9DwpEMAdtxx
9SNuEPQS8jeiFTECKIY4lK1JOCYR6YUQ1PoNSxE2p3BbVXyFyJsZGL9iL8UJpOCrhA4Dsyb84Gz/
lJ+EzOaihUhVRcLqtUrj+zuP2DvTs8tS81wHz5jmAR/09+n7cfL0WEkPvsdnrkJ7eSXkJYH6KA4a
IxJ43todF4y/tnngrlJVPVtfXPVQ0a1Jh9WHrYe9uvwaw13yUlM4GN8e805ogpvVd1BofMpqqH9b
B06ZpAWhyibWFfb/ayDaP7kGM1kJuoTK0AYxi3mFQ3zwiJQBXggoKhoKUZrYHjJtdBhs3iS7vkiZ
k8lA0vRwGZGTm65U+RhVXnccG9KeVoAO9aIPF3goqoomAGdKt7qvSZqsDCE3Gzh6AsIIjBc7VTl9
YN0yqrLT2F/l5n8ebSKtWp46oBLQV3mb+2GHDRadSj0tTU+NbxAJFCHGAbu+dR92T58upbPUih1C
tPP5NSkCatn4iDQ7hEbk1LXFlZw+ESnLeOw6PSAGzW+ok4KN7Hw7kR7AJerNbXZOQJ0l/KrTX8bG
Modw8O1d4Rf34GaTYmbPpkbeIDTnDEfvJjY/+rgyvPy0nNPEcL7/ggsC14oHbsdmRXgBQ5Sv+xWt
be1nU76aWs7dD5hrcBvJsMMEjEBpZX6YjjictDBF3YbFAjeXVToKQEZQQk0KJgxBmmI1ZMOIWpwo
wKNrrXJ3ZyK6q55gmIz8JPDTm1Xl0dbcffgiPjVzUh2qgGhwbfoBcgxJyb4vLWlbhj5bQWD4Xaa3
s+BR8ruoMwXvFsFn3d72CURKNcluqz/COVypxeQ2n25AWEKQzD4O0KzPuBj07tpaC+ac4x/8LoWv
ccHSiFfV6+zzVVvT2iP3XB9/XtZRRKr6I+5KmqFHPh4i1Xvr2X5vqSRDTDhZO1U8NLaeXQEopPcK
BihVMgxMdijw1JT51zxHulnsnFo2BUR60I+g79S9XQ7ZFQLSDD4flHdkLzKVh29AyJoUrPcaDtKP
lhBHJFgN2XrUs9LOBXsj9OTEU0ohrIWW+jPDXTSe6ju5sgKNfvNV08No9W77qR46YixGrmKy6a44
4z7kuNcyIzA36uzmrN7yZXEnGLUcb72xBdB0Srs0r8oSriZF9jKZsarQJa7AVPL7VAisrHo6T3p2
7khjH6SH35UTJoeGlZF3bTgqX09idnzjPN/K0x9WHbVNYRPS0YaguhecE9tBEwzg5OTM0uUcd1KI
Ex1xYKkzEVrffL8rY4fihsKAV9O2LyWtsAyb4ZzbbygtRhxFKLBjrAo84gtnZz6gVJbzJnEGjQ6a
n026PgULIQsiAVTd4UuMXk4faz2cIDICn13X4cW/MlcZs5eyc6exUNw9yWaxgf6TqFFJP98t2qJA
dnKynRIyBqPWzN4zszTQlUQ8K29WV/p6RS6zWF8F3RTgM16/Mens71/50FTfDIRmiUjC1dUYyggU
qTF5g6qEKpbR+s6t/FtCJ7RMcO9omr9Pv/TRa1St9RctuY4EvpnPzA3JqIiJJ2PWM0XiXcc4lf5E
1NiFdxfGn3OAbzXHJ4wArKS4Tov1S4kVOCKOJJP7zvT8ZlayowFRR9yxo5cpJVBFZRBcwViwe/ef
A7VtDDOABRlwM6hUgF52jSePXEJ18MkpNdeB/yix0BaCpUZKha21UbMEN6kJW7EVMEwUGvvVuuzN
Hqx9JXfiPhaqdmzVwkST2WqEuZL5Wvtd3DfG9518Kv+sfYQwNb+B+175w1QVX3QbqoHa/zyVnVy1
HCZDQe4mfsLAfunT+yT95/sgjcogPwCrXesJxtE8xugFBtpzx3ZrqDr1kC9JcczYexrwSaFZ9EI5
RAiOBtmQXVuj7KZJtvO5+jgbNb+GkIn0JL2RHIo/TLvwbocHn2rTGedCbAzrSqu/ggcYABeD4glh
hS3w1KUlc7uAFCGEOI5qv1JwW49iUyUPlzOB7ggWbMOV2+GAonJ7KL6sgc32lNeKw8B/iEjOn4S1
roK8uQjxRjYCx6E7YiCCdex1DszB0M6D24Sg9wQc8a82AOkH6HaKI1KYVVK/gew9yuLpB/KGVO+I
mC5tCj0sISz03xbja4CuwDWX+UbNnu23KTOWG5U/Lz4ssQGqF1yMMHitvdAA4ZEgtCUgd3ZYXFZy
i+0YXLoLRtL+KAipzdU13LCb90BUtjgGfLofJ1G/QdX2DpXRWid4/JT5Yw0ThAa9SWgTzGmjIsrE
n+x+6BsrbfdZ8CsGGolVAMRZ4a70TCeL3nX9BWPMvBf1OIsczFmU5jPg3aTM5xK4RDK5EMo/IBx1
dFIb8GpIpH1+6xFRwp+tuYC42HYcFtgCL2W0AZqdKGr6bSNxtQnmqUlanAtzTGM+W/PxFpLGKXxm
Y18Xja8jB13XvaAjUsJNLk5jSuX7Yk3iomG12WsOuRShPiM21e2yFfzwwtx5SpOQArhXhsQCGzHq
1gRpbgyF692R+7r4S2VbwlfiiS+0dPr/qt9DExRSOm8uemjJOPmnw1OI1wfWZfJsg6/c8r0OlvZX
CLF+HvGKsTkD0j70Dm7DXqLlrWtth56wRvHtVsadr8+Ylkvh/m6LWGKxD8a0jcjx7bSurzoSnUIb
mD5c1LZhxUEwAy6xFC4EwnW6jBlb23rUZDVHcrJ+Q2SgEh+M77tt82IwFahCUH4XakBlbl6RT/Sf
aFwwidzXI64rMD8ojTMbP7DwShNEfUiBG6YXRFxiTsT8MwzjahtJLBD1sRt0o3vcpBTF/hm8lItn
7irqf/wbdNcuz/+W9yImefiI3J2WZpU91wf/YanraKbIqwf0mYjp8fAel/j29KUbCgQ2QAfFv4iP
XveKdjM5NhfMmQWxIxUkd1RDY1XDw3aOtcz6Ar0ioWB5XZWY1Si1jPKHb/7+9PV2S/AsSQc+sTeZ
fKQ4xZY7m/ryTXmU+S6Wp0NzAkmDCiuK991zqE9AYGDn6safHqUl3IRtTcI9FEBhjn3TdlTtZFnt
6jHKbhpgB68Fr5TKoisFgbAbC/QE1rxTcK9bpUHS/7lTomcmdipiwa2f+HELNj72Ce1w0RFMJmNj
8lsAkZZtOhlSLQOvqoEyb94sw9z72cO2RmX38PCh9mQ3KRmPZ+q0oydxkm0u10sLCV3NeWjNUDs+
neb5F54G+KgI/Q5aC2Ud+zCUCiMBqGwelLT/98Te2NTwIGPGA3B9ezmQzIPSAyw+QXw7D3+xQTAA
XkYXjOXXSAIcsSgOLibY6vAe+2VAwofBW7sNJMxrY5NbKgSjtYCFVtL+UMPGOfjcdf7elE7xx7SM
+5MFsBKybSc++DZMzs9/4tJmi0RvCjBH3hSMeHzTOTecYYuNOnyOXId0rwo4a5ViTY7oR3nv2pSc
yKXJ0ArG5hkshxyVgtkfjnum3QyTBqgHv0bdRt4MEn9UndX4SGtWvZ93j3VNBaSO51RPku4tBSDM
JTZVIVt30IZNy/woF1PzEOU9+oJAn9Yp0ktCEgJLsPnzHBaZeCHZCN2UaKmKj39EjIiipFQdJNtb
1yUScrSPUlG3F0oTKpaa5z2zOPioP7FpiqzbClnQQh6mf3qhPZUY0Rv+M4tS1FmBHRnA3p+2VF60
HdcB73oHt0JXahDIH//OP2dHdns4iY8lqnAaAWHR1ONICwOJKCtmqNBLIbaVJbj7T8LowOcFWf95
eXb/rv65LLRT1wCodXENfXNQ2FYaTK3C22RH/Hv0LL+ApGX459iGkc8JHNopLwaZ6Ke9Yj+aXfkL
eOmbyuQc1CuaUf+CFZyRqZtx5KgplMwy1AueDP35q893IhhgbTc88lmBzSuUQjlkQUp7mO3v8HW5
W75yD/3601jlUcV+M32L5gmf6nVwCaxNn9cjxMa28qfuWyBSDwtJH+JXqpEXXSqReAGI8wJiJBeM
NWQYzAHe25iiTFVnsGcswSX48mOeTUwvW3E/9papRjA45klVMoRZEfvCLCYLLqf0CuzwYiCWKqjj
gTNgEruaOs8xug3BydQfdi7WIUafWu0K4Np0ZwfwNT+W0x+X2XOgSAvFEDcqlWo6KUmhr2lepU6v
kwnCLixdh1YE/1MzOkH1MWa5mwjm26i5m6F0UreOM4bc9cLlZfP/5Y0jqQWUbmfMMXt4EWbN2ziJ
0PapzOI0dReJKZwDwOYIMcdiNrSeSjIfVyOuGAosi6Es4DuwxQMkaT4rXCpkiMzAi6UcB//1qIve
fvuL2pbmQgaMSCXJEyXArEDWZl0qVbmW4JmAs3PNhaEn2ap8MOdVeaUs9NA8NMg6HslVnXQJaOQB
fyxf1h6yWpchzLZlgjo0FudX9+VEXn15YtcndrKAcGE70zE5E7fbQ3YRcdMGfBmnOqoJ/pteMbnO
UDtT4OO2yzA/Tknh7ebfhbp8tjIdH/ydjPJHaG+Fv9DYFqqlkzj9jUjZ2dK7s4RzEGxqYAd8jSzN
ZUTZQKobb5oQTYF582+37yMinqPEi+Ts0LOIpURYCMy8L0L42uCW44g2RKPDJ+QK2KBjLtOEqycT
ohjO54ZjE8LVZqSD5QGBoYM8zI8gxl8PXmoGhc9QGriU3mHH8Sn6XNcOp0aL/5Lmyvyur4HO/81f
l0QBd2iymvJ9pJ6ASejdYoQOFA1BROyb99s+8YZT0dCGKD1NDn3DTyKuB3wkUHQ4hI31wPabGaSz
jlylzjtll/O92fXXNeP92idP4R+D16zd3B5W1NuDAJjGkj3qXFp7/L6f2m4N9GxIDupr1g96DmoP
MqO44mMv4XY/bXF4YMjvmQXpgRBq2/svsL+DPeaTH9pGz/EoJ47Qg6c3jcSbF1fa0ndIGDMDq5l2
RABUD5hqdTbd1aiS4h6emR8Jv6w0PZCiPH+gy1+IC4pBn89RjYsM3YzUcuAsrlwZT59nAd9dB1Jh
9LRWBGHe49RkobIrAIyqJXB5GsluR2Cs0vc1sGF/AOhagSVs8sK0xlmzGHyrCWBqVOnieJ3zqCG6
8nSkTp4ySI5Ve211673fwaBLJ2rYR+fPBl4dbiDLe2RuxI38bb96djhWTn3Lrc3ROAnin0Wzz3z8
ZTGj0mpiQQM/VtqvO1ScH2uwrWpDxb5Kv+h/ajygFPtFQBT1r5U4hwyszQSPZ3+BdbWu7UP7G0f0
z8hlDdcYbtQqYZmcQqvYg6iZw1cPkReOwSQR6/8tmrTMvvSiALQXC8QJ2o5nxymxbTsSveAIoSFO
bbPBDAGw1/E56NM5hgJc10jV6sc/NFGhVjz7p42xWQ9LLzQ/+6qRFUQFeNxYC52fnpO97wDl608D
zaQuL8MN1DavSieLiudDxffEPu49ObwPTTePuZs+WNUtkb8yT6nXCDx2xTOKjpRgkq7bNG1jTA/O
qaBeFq09h0goLarohIZbKfZLB881vDHAX22mu9EeAbhDa+/7najJtJin5D91yR+9fyszuO/V7FLD
wcw9qs6eOUg5neue55b77hiegdkox1aDDe1XpomLdqWkuTbc0eZ725XnPDTjXiO48sp7h8DlRAdA
891F4ZbCGTHud8DBi8l1OLlBHAHMqHVIQxeh1cRJ0O3Zr2xg7PSjmFSE5+Oal9E2nhDACgtFjonu
KTi0B5GCfWJ/R25caUx/itRWnmmeueoSZ9PDollIV7oWS1GKHZ2vmHlF9qw7IwZf6yd7msPgPYy0
7tRlevTURdnanEbG
`protect end_protected

