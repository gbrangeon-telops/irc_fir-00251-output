

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
PT1CWY3UnkDDUklMeaNBhV6BliNbBJfbhqNG4kOV7Gat9/z6WihgIxC6lRE+3ldfsLvMpYhy8uJ+
25GNPlskPg==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
UvJJPlyuv70VHT4mYaiqDRKTOeGm/bTLqTJOIy8dhI7h8MQzd+YE6IQThFVGwKNg1149OMGabrJO
oYkVzjNGF4B9Aleco2wvOpKfvWGZDwt0GGcY0bPwCYhgwzblbjwmCgPjWkv54osNVTW8DzqpXiHT
yqTtBlllC+UP6StZLKk=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
IvSnqjuvUH0Q1DG87naNrsoN4LstR88Fpjj6aMMwh+f6Fho6xAvTtV8qJudD702FeycqdNzlt1ai
QXhCNPnT2uuSCS75+mdCpNaXrbRjxmX/iWoxCnzawaHjNORHnFYbE5ycb12Je0b7xDgqmfK+x/mm
Rr1i9nWC3k0y2ultNBrqag9B7JWz2UiAxNLz9gIhkdjfo9uuq7n44on8tD92VMcRgnjXzhfwsV/R
WQcm7g2SVj3bLFjNpwKO0qkV9egUmW/eEov7KDZj0D4B6HRqmpo2DevGwrEmNSVhbBsv+hYHPySs
vJezY6TBoybQdPcPOmulaKi4zQJv0qMBHUSRhA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
N4Lf2o4qQIsZJ5JVKzqV74g/C10RJITmHA7UkLNDA0jMmd38lQ4sUVhO++1w0lqqkNK7gbVbdw+5
aHqNf15gjyNPjYW1ZhVXHrYiWWCWKhn1CmdTyUXz9OVBdu2lqmPJnjbOZQNbhaspal62bK34xeW5
H7uey4lH4qjMdyRPWyo=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
WmWXhlbOXU4TrFQt6FbjizC0tiQugH2eLLLRZI3zQRGusS+51Hgzx4mz/p2wkOrjF/inwb9EGctX
9EIb301sFgIc2+iI7RGNXRFy/HDMZa7bViPHFvPX6IIbSblSMhaUsZnDGZ9ShEIypX3t04pywLmp
oC8cxeW8KJ9jku9s++a0XQ670LJrlDd/u67e8zo+xwxrAToVkNJSGwQcgXMc9YDwrXqUemdrJGhD
qf93Ms52+vFz6ikE9Bpwux97WA69cn9Tx5Hhj95T7V3DeqQDYaa0G162sFOeOncPAYjRFsxSNp5b
cwcMCxbjJE/oLyWzhKmrRPek289fPpANZ4f0zQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 45744)
`protect data_block
ZEnbEpjS9XKH4DVoAMBAg0aLTlKESiZ1h29c43Zt9ptJZ3p3qkBBSaLhGZwwUv+UyvNHHaaojRpP
5EWPk8AzYMlWr1yWAOUE9szxeFD/wtZ1Zegc7scNHZrqJ89OqDhSxM3UB7qLGx5wq6nmHMlXzV4x
hg+g3pjsOm0QukIKUyY7Y3Gr8+93XUNLYjFSuDfK9Rz8FZJ2QflX5SnCtJI/xOUy+Nx+vPsZ2BwA
pyAE5vniVNrn2R4qPn/xVejJXl74bJthUUbX3/r0V8rJXawk5r+3BJLwtqF12eGglaEk1DtG+p/j
D2/UDTtAuZPGNfSei/7bregrH+W159SpBr/rX18pL/QI7P55xlXX51vZJRnQWXehGnRTxpi8kkp3
G3NTHWFG4ZmgnlYZmSNWuvoZ5/FHb0WZ4A8qUaQ+Bybwl2PBO1WGW/bhhCx2enNlHUeG8dfzDdEC
u6GysrusUPc3H7/Oa3BmSSjxGieb4Dd+2XY+MxQdRkr+p/QhgTQaZZRxpCwwPCx+KWdVe2txGnmn
tpB+AeJc9XbG73mDGpBW9HVxDFkA9NZSMjPxw4xapHy66b2V2fyVC5pGJDbCWe4rhXtZ8fY1MLKY
cayEh4OKbvG45aKLM0l3a1nrHMyzkX2UkZndb5w+VmsauT8XLfrEK8YcwXtqyIjBOelT7/mI8teV
dLWJHsVbZIlcu2jv0bfxTK/gTwAayV6aGUsB8TyP2r+ax5wraLX0SJdQyd/7z6Qf5Dw2nBpufFXO
YCDTF+HHgYxiw7b2AxsyOj3D+r3C6X6MzsPqSaji4Wg11l4mwLjryeaSsKsUCjMWILkeleBLlfbt
A8l+XHVumf2AW+dvUyeZWf47quAEgkNtL1UsL7wqc737hD9+b9nI9Rwm3ScbfvVsY0cL418ghyeR
sk4w9WWhat6nH912RdXMj/EAKbiAT2xq0tU+MCz8NEEqqccB5hEv2eTORWI9SrmLirVTxnIKDPpV
m7/3NJzzZgVKmMG6/DyArW7E0kgtcouXRRkGtWO0zQ3x7/pReH829tSatGaxTSUvbplX512KTSYL
T8z48NelDC8oqi4I0OPeLHssZqFg6TT32RfAKPQg04oWpS6w8/lwc/3/TdJjiAgzzOUCS23l/Sdx
7nu0NKtWybfkeWaO3YAezPIpEnQ7aQVmT+eVUrUoVGodfhk3ETwFXTmXBxWqQJw+zB4L1fi4JLlB
cSZU7hbghdWLqFylYxaxjB+6Zrc6CtKoIBSwc2cvXCzPI4v+SXzUJFBc5bnBLyoT4olUP+kp2Nwq
OmsI9cd+/c8jMPb1tTNHj1PvNfjRAZSIroGuAPIVJWf58QAzsS2QJESxqrFrNo4Lw2pL9EjTmhay
kMs8sf2OnE2rlE1gmVSW7tb2YgLf2Tq9KfFCgWfkwCisNLTyLWgGShsnsXPm+G/zxAfBYHrBpZZ3
wuXbTTiTZkulGnIdIixEpL+e81/1WmFnau5VB1cmTaCEgfp6sMCadnMOEbQ3qUwnMAEG2iGO5mkw
friEVaIGTSURIGWFp+Cr2EKs4fljTUjvYQUcX4yf8WvX0G4asa8YPwA6gtylMYdxDiTEv2iCTX2L
htmj1bAh/RK7CEZDm6Un0EebQEs8zRN0q0JuDNd5YmwA2O4qKXpSPobN5EiPau23FpB8d3SJA0PP
vtgiWcMpVjUdnxQJ1lhkbPAdey6Hr1Bj5CnMOsBDrG6tkTa8tIfLZna/XPW0EwE7LW+kgqAfHvYm
s+ob5eun1j8ybP8POaCeOf1bpJVDSLq05dtoI+tfJni6Mjs/hYIU50UjJg+KazY4dQ9shaX9e+wp
DYBixUGybp8Oj6rDdLcuKmLpgQQRd8Wuil5ga094zgvGUEHpVBeAwtKZ5FjvItyO//cwDriaCYpG
UONz3ljOJDALe7+hX00gzSxfL3c2cvWSA3VyeF6Vx5UeNaaqmeESL1JlZ4DV9L8JdXWDC8tPE7S4
PVPNksGx3UJoa/JDcs71/kjbHz8xmAXGN5M61QF8WTj/rwsgioR2/1bxnhgqLI/vhq7hrjp3X892
rv9J83+miK3fPdM5qblNcT7V4mlEnhIfpbtShZPRLulrQA0dAicbcrrOBc8WRf003iNcjCxNfRRv
MJdmAo44kacGl4IAy7a5cutZ4kri7FoHI9csiBYaRGBAPFgWsH9G4BIw7UBzBRN+G5w8JhE7GAZA
PW9zN1Qy1WrOuow7sEiAu8CIoKHqkjizC9MPwvj5a0qYIavPfdBdcS48R1TKPnGXUfTWx0ON0iHZ
213uMjcVXTJi8unpn8188fWvmvTUjdFenh2Et0nQFEej2jOOJ7MxCbua0uyeQd8jXBZ7/Mz/SBFw
OD3EFdCWDrSJHPcfwnQRi+qpbAXCbKrU7QqeuQHdkwfN80NvpWYS+rzX5vkGEZHnhBcc/eTAG1Lg
WrZLtqsDmhzQb2xoqv7B4NkZeOoVU2P6B5/PNjnWQqipQB9pAq1Mk3uWlP+lA+qyp6eY7OPf6Ryu
VrfamsCFXH33HmmY9suRfvfAg2rkJzp09Ku6BG19Sq0OnfjavaDRNYD8iFqTUxRX09v7Ux8I8Xdx
h0+wpB6Fhy9dJrmCE0dsEGxSHpEwRzfVeQGUV5bNt6gMPvPaTUXyLWXBRXHRvnGDay24fQN9Bzif
QkAE+DetpDLWPSVMXml1VQ1+1L+bsES7vuTTGmVfiFTPfBPlY2adT3AvtDhkbCI0MLha0ZDxQofr
0NVfIJXGDRUyfn7BE5S/b7ElBBCGhB9JqqOeloNqovjSLudwb0zkYIqt6js9QKQl8rv0w+gtI9cD
iv898vdxoO7zmfxfWWrh1xkCyoXG6fbPI3E/bIHnjOTviLinj2NUs7fVyuEBg9vkQoQRamb/arqR
OKeJMX6zqSc8n8HNzuy4aARaIEwCufxqQktiJWNveMiXjqewUIMR/e40MpDDHX6J8YNECHul1miW
d5XrYzInORsiz57/SxVaa3FPXGDySAQojM3/uE+QCGizatvA6G/Ij164WwztR3pVWzfjjQq29Evm
AV+ZcSeuvsh5S5f0aQtEY03oJ6M/YZ2QMAMHWwJ2AMGFk+bxTcXyYnBzVWVDY8txes5AsHBwPpv+
qX1Y+KYbXOHrFLFH77/Z7/4WOkNvsrN4zmrGVkn3uPcT0EFL0hFDMcZx/wSDjrWHuhnY/tR2MC5r
Ngyn1osjWWX8tupbTkHN3U44kuvzxqlEb7CFkFnwD+vdQAv5ojaKrmqvo2oAKFUP9ohGlaRANKci
wpaudjNSFtggw9p9nvg7yxiPQBd33Vr7ZkvkpkVYDgxHz59J+bHW5a4VpuExwq3EevXvRfDKDOnk
LLnVaimVyhjJXXi+cqyodRrm9Tr2KlgW7GLSWB3qcFGSS4i/932oIqnL2WKxLnjjEAdlR7ObGjwn
aPqS7ArPTOwMpoRc8DrRUxk/em1WR97Ra+Y1NAlW3ezOFeIKCVvMokMgWl/k/RfVxrEhzOCccCAm
mlRoz7A5n/5BCfrWAtJaXWy7nsX7wftZYxrCcxtS5FujHNhG8oF2j1g/uVuM0+GbhPzNADY9DccM
lW8YxlmKTXc7GXA3/EgZbhBH5lrJah1pqDCYS4RiCpljsSRIVwjvKc9G2blTvFSF96DpRyoM/H2v
zX5L7Y0DOLQESA6eCopuYqEmLinxzY/bc6rb8U6Yr+Q0amfK9488GgqEtIRpRCjtCstpy+rXk1mU
53T8bNmYwmBGQWEYYz//rmyCsZCh8PjNRvLX2LGyp/huslXjUM6uhdi783ooBNJhvP1ZLtT6RP9/
kbj1il2Ny3c6YO1BlciwXMqeUNpLkxFW8uQrwQUN2IWXXPM0di4AIlcwZleQy06ro8ik8Rdsno7t
Ud2biheuLm2QgqzSJdKo0f6EwN9HE9RlajK1Nt+zzYRp6261b9S3xI6QRjYsHDHH+yw3qjGRN+XU
ECVdpE7DZ+Or3S7YePMcO+3+SwLzx57iSBbIulDDMr4zSwWrrPkDJTvlTb8BmjTLp2C+NrcaIx/c
MiQiI0hd05+w/Vr6mgv3JFEGaulixfU4tuLi8nu+doE0G8/gGHdsC/6IPD0icf84KTgPaD/QPF7d
AyYH1Z6uvv0izcnsovjjvt/u2drcjMLk3j3b5YWo9MF17jTX6bDEP7r50XYGa3RxxkK9ZQFWO1WU
PfFscjJVtERgmbu0g4BHo30F6dFY69L3AC8/ZjduhuzlH+Svj6ooHmhNSpeHgZqI+Eb+kJfftnMB
HnqBqM6vJv/wsd1PfLEBO5D6FPhk5er/ej9cHHA4ZUHqGRJoInitML3X8S2jLmeQ6cpWYgOUYfMf
0v0OWqkRCKIs+HsnTW10fYZjxxlOaGgVWMMcXsyGkPBLuRRUizD71QbLYDfWERRFdy/TsgwCZv1T
IjJKej6PUtVjzMVOHACWyAbrDB53yzLoH4PDLevjhP02pHqk2g2XYQXoiTUkGpua3la1fKMvu+1q
ZYCBw3RJgFZrSHnRpSWP1Tdz7VMEt8YheDw6Z5Rl2XQML6Q8PL4Iaxs+nlovD/3QUBPWUCMp6r41
sb+I7yMd3jhI6T1qgiWgXF7MW/7hR0rhHV9v+7v9+fGZHbEin/+clEBE99YGgpbCCH7YPYeRzRH4
LOKcUPWm011TUEHIpOJdK24NELMVG0V1gsr7/xJoYaEisqvMd5qa3kU0YixvNanTKZtGeYlI2tXT
6sjghNgv9CuoptOb39rkLbFYWUxivpB7g3TXjTYUZ7A6miM/W7MPUe8YdifKy6J5tCVwfOcilZPh
aQKyh7fQUvh4wAsdVYvxSPdOfk7fE/6Iw+sPOza27Q0cMzoxDQ1dXrWwTirAJh5b74oFc4jiHcXU
HyiBQ+BMBkXp7rbJLFnSQL3BMd7HRPnCHbcRZGA5erEv5OhRhJIid3bR0aq4LzXRwNePEP3qNk+v
xbEdnnfg6K3J9FyTqD/uDaOY3kN2LxPsz4yDkOFvqNyNfWwmVZqI3K1KHbKxf6FMyoHdDxiDuOO+
bdq8jtbycS1m87Z1hV6wlHDKqrZ6XqE0/xXAjcxRpW3HQRYmxH+TDz5ijaEfx6xT+JMlEVaJ/B+v
AaZbYSis5aG2WctczZt90otaalVoYrzZBadclVIHOiMLqpnvUa3BR4m+16m3G0dYC1EChQxOX95C
vH3K9ij8hulF6pF+/owS+GqFD5/F78esb0zjJaqw0VDMlifJqteosaVt6Mfdc3OJFYsqePFZU8v5
AS2xOS423XPXanGq86YQoTJX4IjckEqBMO58MgjPICa6joR2Yo8BWCwc20xiP+JXB3LeRP3CLA1E
NJASsBfHV4aWiZfJcC4MrK4mxc67qFdwxywoqfh8d+Kkn5+2vKe2gNYHHZliUpxlPosdq9vgLdoa
w+nwWgxNTtbsfRp1zBU47pda4aO6loRTZQtJYTmarLlWtQ1omzpe9p/oQZizHcMBl+lUeJMkxWKt
vCuf58CZRdzWzyY9WAf/3lCCUowaDihJp3WW/s7ZCAGQ2QkG9cqjCspSEkgUnlPolPd+07Ro+vyf
ebpaHqz2mDS7EB/AwA355X3EPvewlYakxj4lk20jvULBDscMkgEW8wsZlCnDdFXBfRO2WOHPclA+
qcjfhFogsRq9FXujx2qC0+w9658A9xxSCaVmuVgNS+8r6am2hjfqq73HcF3dKRBUHFmsvUFL1Tbx
RqA6VkyA6KkdqyhxV9vMsMmdJ1SzzUrwrolHNWyAIdIoRmRkhgQiS4ENqMzKBFxelKFCkBbb1JJq
g7SPqD1aV3tNDGLfpngaHETZK3XgTgIhr9DC5ZV2RFZLkVU4NfyyxRZUrZ7bB5/mupJsdn1V39Vm
zsykJcFnDSkMouxMgLg852y02qZ/nnaTJq6XjqQGA5fEdLmGz2mDBMHnNrG2iVkhiQxtMLnJxYfs
d+LdiPpmokLbPLiMs9VdtajcNs838dMemD7j5z2X+vdlLPvVpGT39qyrhgfhcU/0g+PT0ch27dOe
qDnyV/pcWaNUEnXb6RWLpLkqIqcg3YqnU8yeBwGyTZCgK9HMTC4lYN+cvbuPnacgxiWRDCOyRq1b
s6autJIibXqlsAIOGYpPQtgns7gAw1Px2cCmXRzPIwFYyoljerFm9Lju0n3yB1ZAghWvikgP+HLS
y5flYsfQ7kwmVCQPjfsAlVuIoNyXjOhZbC0TC+x0s5ZnvQniuxMfL3Bsr+q9m996jMXuL2HHLlod
DOZTOHTFIyQC7PQPxoBoPOtojJ0yeHVANvCuJbjrjus/7phv/U64R4aUhwjZpuVD09x7Wsh3wTgK
tw2D27PIm/HlaqESJfzopUQOGsgmMLq1bkbKhs6qy1q95S0XQvZ16kvwwakD9afqEQxNLZeFpS8q
FYghg3KFuqkHL6oDGBfCRRLNXbws8bSAFtrhHixjBevAahLTRWkeb20FQTdQUki4rftUA47ra7yN
1y7yKvVUqLUHO5kCrEei1TfHx69/BLNP/3RiuoRJK8qqHlwqaSD2ylXK11ri9XxP0i+elqSdR8ro
SnFNcL3ikddPedB41OEGqlA4aEjHtOdmpaQ/N7focwq2ld1Th06yUiagPhFFB9XLNxIiGK32/tyQ
nmPpJOd5B1JaTKxSddI120nYwbwaVCH6mJs4vPF0SOuVXpt5pwuZNQO0Rf2ioRxOiLrWeBXNchxe
lhtTH695ceijO/ZIxEFS91QTFucLt6Racn+7bBxJq3G/DfZooIp7jNT0cQCysS9gcMVkYdXQOS9O
xZ3jeocB8Ul4IQq3PDbXlhqESzpcIIR0+x3xO4QGhwaRAg6JnMGg/dO2d1ZxwTOoFW1RhWqDzgg4
kcZ7hRYxRcnbsBZ03m+onwAhzPVeBE9q6MUtzQ5BwV6YLYHiCEJZSR7Zw7NVD3uSa0jugE5Ax2Ee
GHQ+gwP0s1fvcB3MWKjft9zeCDSp3ADX6WZjb7AYiHHYzPZBpmh3/4JVkHdn1D8kb0t+qdx8/TGK
HpA5gochkL6WrAo7OXjc/OE+3r6QQIbDg9tyXrGz4i/ySSb2PWUi80Bn9Vqb/2TqzqkM83/y5ieM
DI13StOz1QfsKJePwKV9gHqjdrbLYHQPgHydeBEUs/d6CFuyiSXJHjYxtn/i02DwSdMebbW9k2RZ
2X1KPWIPJNJPoHyDMD/BNPbNRCpptrvjAR+uI3HItjKTNvqHIUMQhPzZ36OCRdkLFA3S7tV5rL8b
DZ7aJz1VDa+nf61Fl2FzjxOJhUPlusAFSEM6l8WVIFsULnVZahWZzDqzVhr+wEXimUHO54yzzCPR
7JUNz0vpWWTgZ6fEDc3GRBHfKilWA4N/Ltym0E/vcA7IMcjutH1HDCKHqEDaN90UI6v4ozsj9G6M
NM+Nm3PwEhszr0sr7QomA5ViUBGNLt40x2wmGADlq3/2Y29uwuZzourPZpXR18I2XpJnJhiRpcq1
hSaRcH5DGAjL65Kt/p4SkKhheIwBehGapa8IGQapoWHjJy5XW6mF0XsxfcBRlE4G4Cmyj7vODuGl
BxjKFz573/aEpr7ZM+Mm17zFdFA+aV2WpEBJDgUS7BQ7Akjy2jfw0t4pwZeRZYNdfOFlHdy+ahD0
cvhaJ6pzSWOT32KRRxGtpLoWPiBuWdvQRJH9JJdYp3wMSo+DhvNJBwkZpYjFVrwCTB1G/5L1fE3h
hAv9EgYtPJaTCodQEj0bGQQ5fAur9NJqpIbQIT/RIt1lu/uftwkMCosEcCnMv+eaXqxCp0MpRUbS
Uvt6BOtNsXT1xChcl16+t0nCv2KyLyEuDZ+d7608AQ9BrjdfD0/YeZjCAd2iQvUWphFfLgnVEEbW
GTsgxNAu2qA/0cx+l8MM4zQJE66A6AXMcyK7Dz9d8MLKHkWPOKlM7A7ESeQCFtFJUFoqzFRvVa7H
9erOs5VeS8ElZl6YLLfWASyJE3pA6WnHps1MEvVNSr9gw1xw3Mdjjiax9Xr6nBdHT+KJi83dnrto
Wb5G2F4LT2rJ6r2iAMHY0n2jU6+hz6j4AerwJoN4Ks+HdPomunLyqeHzbz0b37T2rGSt8FMmEl9z
qZkzhjVrogRcaUosVlatK0V+TnzGyxl9YSBcfcK1YG5jab1Y6L2mca3oM13XO2SsKADA4CSXkmvL
1BpEDFcGTncP53kbE1A+gVb/G5LNtJq1nEyO+4ZFtOUGnL/h0zhjY1Ry+dAx50vGlsH15AB5/HOX
a5jN9aBUeKiyBbAtdsc44thH+jdl+ZdDUa3CE8eAaAn9aiYYeiuezIQrWXF6g4c0U2A+26BP8j3R
igmAWvCGVBARCJkm6KaSc3SpHi/9GZSHU/DVRTt0LGgGqxoJ1V0UqTzrKtvz1wXvYjZ4vpy7CYAw
qVu/lcV9yvEL5anPBSpUWHPitW27wBf/FYSfPwt6pIrnd73d1pD/SGQmW9yMm290EQ6M/0+ruT+b
+CdTyHu1UHTKRbAAo4B4nFC0Kpgr+WWC2fluqiGu1sLE4YPLhdsFKnEzzqukDNoSA8NWP/7R+fzd
BTT6BHzmJf+O8E2NfaiW8+n/JCalE9DZPGiyzeCDM7r7QuaFKuLZLt7D4Xn76ZaVa5+36wq6bDUu
0s645ZL4l+eXW2Tvee2o0KowIKP8BGF9t2oQdfI6WrsKMpRykrYg3CEV7py9hANC+0zRKQT3+Wfp
7YABrzvb5z9W1liRx0aqBONKkQczKmTh9SLIlGuAmcByRxu6LD8uohIHBOT2h7vuas374g+MnD7q
Sx5TCiAEor+x3OO3YS7OGhlRPiRV6FawYD4pclfZuWRLFj8/3joN9ibL9oiJw/H+cERcZmfBcX6U
G2tcCP5GOSWtslItwfvOkQlmKyCOAC7Itv+KCXx0os8Xp4ipflRS2aGX/6v8TDVf09B3jDzQEVtd
TfHghItooI/pGNFEf4GcPqgWTNxnyZ6k73RgSuZawkUxWa+F7vd3ItirG+Tx6S1WI0lE++/KUxWL
U1xU7HzehCWg6oByFs3D9u8Vi18wrplN0PWUad9JwWRIxG6iVLvE1nlNeEADFH0Z2um4/DnCxNub
uj6LhneEP0iPGMSdZkxuDsK3KtNGgU6G+HZngx4GY6RvwkYYEeK5ciRP1fCJt+S49er98vowN7KY
xiok/mzg+LEWraQlnlbrY/YdWA5ogFMjNCosf+Xz09HjJdXxZGIYt4ATNnBn30uc3TKVqwHVI8JW
nbuAMWpm7gEFPV+5Rpg4EEL7dfWLM9i1TL4iZZhNd9I3krZxQSCkF8ouiSfCNrg5FWcTy9n8F7GR
GnkiTi5+sWPTR4FnxDALF7t3AnBRSkcbXiR3kG39Edz2aTyZFZ+1eyTbAgytU7XcDihc8z5o0z6O
V5nVVDpflSPGZ1WgliGGjQUYiX18ZrMaCIZLVEwr18TQueO8I+WgahJeVsnobXMt7imODRIl5axb
hOAsvQ8dwxvb6rByMStmSfh7BSPG6i2VFFHnMwH32t7QTRITo4S8qz+okTwIafd/JrGpQ/VZuJZm
C9e6Sink4waBolRDkIerxVbOO+dviYO1dcsJ6esO0hLHZMs1u0h16Vgk8nkM/Kk2+Y8yZ3fyZxv9
v62gnw+Unqg1VBSgQLvt5pTx5ZGtSnW4PMn21mhjxDSeEqBOh+g9dCx+vKOt6suPCI1UXRozZSOh
QwqrBoQkMNrMvorG4FifMBEJ0DL8DNv5n+HC3HclHWjEg7Fwi9MmQzpOlyTziO2nwMxOBarGcl+B
1iJMBHSk8U/Jr7XnpaN41K1fYHCvsLtqBlzxYt6koBSjhd/HLil4mFMIxLow/9kpynM0qt5v33o8
Gb0HvTTl4XWiToUdCJAg+HB5dEvGL56cw0v9Tp28Ou0NDyKeuQsAMJkYQ2o/H2cwPSl+zHui2wZN
dUG/xEdKSV/9wJUDBQ+lwz/Pb5oOQm2OYQ0sRY2TbKBbZ66N3Ier6JtXTv79W+ji4ARXKM15Qfk0
iWGExLxAqEtVhgdOd2A78n2/7+YRrqVxbtLc2Hawg/H2YO/UEpEvQ+bhSvuA8cYqOp5Vcpt6SDj+
pCqIc72cUvKM8K0ANsrPgbWwjpFifSRTxyApfiThsGiT7WTkSw2DMBBuacctr40SiExMZZvri9Mf
nDgXYeAgzSYDnCmFIrz1/uS4l3YPGm1R647YJjR2H5eFr8PShSw1b+R8jxLIQnNcy+YB2uoW0PIl
xjchj3yLw1hDPeylnoSmNwmb6zbVzUtP2qax8/IG2FVAdNsGCQQE2coXF52u/w2BPwmGncakqVt6
PyCUBXev8XUvLNwlHhoca0hWtKLn6aVgzLDYw7sJAPh2pwieaji7tmkFwigzU6XB3SdwfxFl4Kb2
a4aNfArptPN4muNQO1+pDpF+2otXuh2cx37sK1c76GR88m2Y6/M85yZ9iR9G2tHuWKcyUYEt1Bqn
tzTgWRnXWs046leigdCYz5Zf0alZmZ+fDdSbFneIGhHcfmEnPYbrFmT9uSBoj6t5BRz3BLepJQba
83rWzZB9l0V7zUY/UoByxXm/f/AaVNewJ5XBaE07bNwboErG4vFwJkGnh3Sb6+HEumgY8R1rE/37
JuwtL/F2ZF747hSUnotuoqH3QcNFH+MrUVH0D2bGpbP0FlyoLbvH61GDOq/uQkvpcKgt8wFEXhxY
GzMzTR8GJOwVdXgYWsnwhrap2AJWy19pnWrWdIBCPiaWM0PZd1yTZsVida0teSRZLc9yQAAHU7B6
d/rbO2I7b8kAYB5WM6XNvWhy54HMuMlxNmpDwugwVbsBNeVhdobvppILcybyBUFi2AVQPV/jOtRW
mngU/evc96D6XPlcDyA3qbc1TEq9FtrxjEXEOryWit+s6DSIs+N9cBMhk7qvGSbdIuIp2q/wEsXz
wvtiM3Q0AKe3ESzAEf8OI86E7DviYyZBbQpiLGM0CUHQVv4XPwK7wazwoLA0+xFePN585PhLm1ro
dI0ELqnurE9Akzm+CNHA6EtAnHrx8Wj8cQ/VaEHSVLq+7n+q/2cYtk/4vwFEe2rDXQj2AgVS8uJe
NYo9aCcSwCKd7h1GNP687V+6L9Tg4ewK4Fqwsw+q3MOhLu+2eFnmnTzjEwpJFTYnITi4F0kuKi8f
5KQcRm0YrqYIeX9O9wLRvoD7GRSKz55z0NvECUBTVB2ooaRuKYNiZw8qBMWzEcQn9Hy6Kv8uC8JO
HxauCgRot0XI6Vz+bz3kckdJ7Ht4UnaS1uVtNR4iNLgg1KLo8uZ8kW9l80vEUtdYiQpYLLgIyzrO
yxWGbxJawpmamF3xB/bCU/mx4/3fJZJnZhKlMBy2sr8dffOeRtGPgK0OPzheTBcP5/+jrGS67j2l
udKF69WL+XaG1fNSHxoyfe47U5WiyslSDsxiHjr132/u0ok8Mt/VO0SqM25N178HrpejFzoPFthq
Inc+Bss3GK+J40A+wXO2nFQbYXqn9QiWBFBsKHk1cmmY/pDR48mVXOT0hwp76qPce4U5oyw0EQHG
1uKTvu1e+4kaXP3hvW8OU8YvPuvBHIA+4Oq9zwbyRVL7zkcjKDxeW3nx14L9YPNOSnwumJQs7KHQ
kqpOIXak5RJXG/UhYtUaJ+F3ku38nE0ZX8JY3XrFZ2JYzWcz7/UD8iIyRCUEFTBQTkl/9u0JIwoU
wMOGAT/otO+8k0r0CmMd8n5PLl8Sw5Up34qFrtAVCs5Hh60nKIF+dprmiYMOeZx3CKjNRl1iEmOI
i1siwKUzgmk6X39ynpd6PYVNm72YQixjvYPSbsIte/6JjFKYGfoP6Mt+7dDxbxJzrhwMRJzXCjHL
8ifkxcrKSMRFnvkQATd+gfPCqf4U8o6pxkeQ/k34HEjwJm8JTVopYepBn4rRUmJa6lNIxfo/g3qV
y6J1knTN+umn8gC0/wg0m/7r7ml2zEuQxME2bTnOvzo4RQAVmMnFJFzWGtoDqMB+orz9m/9kBPQT
v6fFY4qQ/UTqIXlgeQGXjmxfq/0pxdBvbUcjE78v43BD64FueSu5BHSNBkOA3fcNdRDN9L73Hpys
tcheB6BZu9kxAuNVW6aiOyU7GM4uc16F95F02jFFHo3bQC1CkAODC3QpLanUA/58UffSfEB08rsg
JxzQiTvYmyNSO72/l5Pf/mnpQYF4/Tt6DCRLE3ndcabKgqYOnkW73uTgMuwEoAvco9QJpJa/pgz8
Tk1x+xF5g2VOjyb52yrAXIlro68Ao65lAAktWdJGm5zRQ9BrY3vbu8StGlfSQyDi854A8XwyBNEk
GCy5YwSRwdiKQPM4wP7KBYc5kXtSmLdLVUNm//Lk9UnIwRrv3PCSVL7Gyk4WPCwx+/pGW3cLzS8F
015LUcQ9QhnT2RoV7+oZeU4caFLfzPJyz3+C7eJAZVlkKuKfvmp+BbgMRzSvvxExP3KRqHN0webW
2X7gJGSz6OMsRkYyVw/qPUYWCWYkzSV06An1gbf7E0krMKn/Z+qGL9vhS3cbBG+88kJNm7DoLqc4
aI+kioOIu5BPHlrwz08j5n0sgTiRUcjWk/+bffVnrLWevq1KsBopFPhHs6Y1BefW8BbD6GxxetRX
pvou1U84Q4ykinkiy8ZfpVTdreu90JW1Y5+Vuut8DWZNKtetXLYNsUdYnwgTU4r6D98xx7298hlF
0KHrv/K9D+psoDVjTzoMaGLXQL8xpz4ztDfEtRw5h/w+KZ9jHlU4FWY1jUuVihE4eeUtf31XoF5N
kVudWQe+FwiGFPgqRdCxbNKOj5lrNc79IMuwZz/iW49n275WMuo36nJJq8wwWSTvNmzBpH0xM9U0
sfF+jxBKkGblUOjfTJzKgFuFSN85Fi+MIArj4rcgejYJfBQUlZDKvE4YYVqHQXvvlbTy2HFwvYYn
Xp4fkPK+1dmxvqSrTSqxCzu/Vh4t0Dn7mrnmuOJLgUZN4P1Ape7M4RS5pX83GgS08z1Ab3cKMfaf
iTt3UkD0Vtx2mTqqiJPE4VMiYL5ZE6QrJKaYF76FsNOst6GKkQiLK57Ravd6/7o2kszJd+xAQvP1
cxyLJlJiFP7XCUa/gTG1FrmYoSBITGU2dAmiHN1f8wEokooFw1eib7XAVe1i92mdJZldPKektu6U
uyPJWslVtsuG+SH1vRsCKFE9xZpb2MbbzZngAQDhDOaW6X7iMtqHGSQxiXFHJp6NSWkAZ97FwZcq
13L42p7vCEkzeSF+2asFdnIOZOfUsi4C1eEkchpAaeyJbsEkPcD8c056dFJmABeMZAr/bNJC4+gX
W8CeUAsE3OYKK7lGT6ccf576gLlhJY/Ha0uTA64VR+9Ia8Vi04xIP0UFJMGESMFrW3+BCtNrduQ6
NbPitj42YaZpgEEvM9TNVKhwLqSK/IDTf7SUdVhQwzN8t79T4XvFEmMWM9t3ulIPfsDXLrFOmPv/
AcqmIl3COMhlBt1RncnuBVmZvLhgsZAWyrWLOQpC1pwrr+h2JxizwlCiA1YiyRczw5DH31gsPWGk
nCHaxNEv+XHJ5XwLbijToazzx7LiMCFrleL8+3aAm5UD3Ruofi0OviTCGTiAqIAIo4+mBqna1mgS
jUYl2NPKG0tKrXpGStoFBk6JM4vbHOWPKHuaEMDgLZo8LJp8b1W41wpsU0TwdS6kbPvn7rnGck14
yh5ii7wusVefc1/UwoDJWvPlzL0VDY81jWs3M7fFsrZg5AMiO2NbnV7nX7B8O/Jh8Em9w5l//IHI
HTjGMJNPjD59Ccw6rE/PdvG91ksJuP2QXt0/x9Bx4RKOKJ06yzo4F1omKDXwHnALgk4yaRK6sEQM
niu/aof8ol7yXrQPbiDCHNMPK7WiaIJx2lWkC1L5LbOVK2tSn+qq07rzO7lvHCpHvUxYmivs8iOP
bPHf6r5CXJHh9/d082IHTixMOjwdZvzghEA0rYWqH2NdzH3rq6xRkxSddZmCwk27kNz0/zjbo3Fm
gfRpHnHMXeKQuCRaBq37AZifzhF/n7HxM28Dg/nlQWx3dE6KUG1vVxc4A6HXifDmgiATCPWLZ6NV
dZgdC+uEbdqrCWA6sGHYUUfFWUO3AY0DruXglj0L2ntvF49KO6wuV4bFiPqSAPf+zlIc1GNM9kwM
VgXJ5psD7GX/6F0lQqxyU6yVAZSRhgoBv3eJlrrUwO9rJhga8MS0Jn3b3u+ixc/Z8P8bxvFZ/A/h
ZCvnO0fBT+yRJFW7jc6EItm9nJkno+VeyOCPIvTlv/dbfZzesTWxsfD2TdczAft0yk8aZ88V8D/G
rLIc4McsGcXIAOg9B835n7z1SmikAqTFUMNbOumqMhEHfHOBnI90VgFU+jc4qtW5spLIIQNS+1Oz
H0i17omidLrOr0MlnqsBaceKMQjxrlzRnzrzfeEOLHhMFXvkGRYVf08qXhcCoAwbWiwA3jytp17W
p1hAha5sQ6uFMmUwDcGNgnCmfLXdTaFIBkkBSWa6fElEUDHF+9n01ySkq7PkP3OHOxXMuah9r+Nk
pFd6qy4AAFfK5Krc1Zglz3qznXmNMFC+XVfJjKYu3Y7gLlwzSF6O4l8IbXeLRTovcWT35eHp29DU
CGmx/f8vDIZ3RrRKJ6SYS2E3SNntNL9pxuHnbWTfsaXqI3t8GFUL8YcKxmke/9fnh3zZR3tBsLzq
0PwqX6ZVMg4VpEcZlReJgFg8JjZTo9NU9JQ/mZQ/a26aBZStUzIeCwb9Wft5kXkW8A6pkJY4PJ6O
4O7mUrsoI1NwYTL4YHczFbMATz51GPP+Jelj5TurFqEJru0Rq+FqgMYwJCWcbn9PVLZ1I3cWfoDz
Xlwz5TvnG08QCAM52LIkz/0VPDNTUCPKX1lLHgfUH5nECbPCeP+9KVRXBc7IILYEFSh0I+pdfC44
lvrEhjLfg9iKkxk1wtCjcrOx0XF+gX9YU+hZp6/rSEWYsAupR92H2AJPuCxH45YU9If83YeIy9hD
ajeanx9HdqGlh3ja1qwSFAx1fGmVbMNeBNiFAp3eOQTLhnVF9GgELg/gMoTh4gxfYKg+PPZ0ca/V
ZYNTvqYu2sB66WL57Fta1JHgDaKjE4e8VB/MWhDyhxvQNkiXUcCyNrfUx5Mipy4pHpIonQWbIyuk
5XPIrncSYWwi/ckoOlo0P0Q2mPv8iu21tgTJ9HxJ1e7JHGToDtX3MqOJJh3VboHwN4JxxKmZbzHg
w39TeKqIuMo8drRMfLkAcG6FTM9j3/YSJkR03O2fEqWNby3Vdk8QB/1QWoQZQyd0DiEjdb/+mHm6
nmXbqY8WV3GqRj9nlruudKIhrjeMZ8qWoaT7ixzPCnJfYyW2XxyOqpdOkivxZxck+UTNbk6OUvSV
POXoWwP82E+04XZpe0L+3jyYlm6Emn4/JXpceivLZPGG1hR2r/gTFJ7VHh/4kRvaNJrYJRrqN8Vi
HzPA+NBdqyIYSyKmm5hNKH0Kw8K63tMLDVawbJitxGPh9Gh89RyiOODv0bBIUrE/ia16RsYtOWbi
4pDHjhS0sJ8sEI7Oc3JzlD4xMDDI6wT0XbYzfHaE8vLC+CtT5oWyH5FqCv67cnt7W2cLd47Yl3dQ
RthMjKtdLpMuXvQmyjWf4mjRPZe7IeUeCVrbSt0iDIwIS0c60BCCpRQDDvM8MLZj2oj5Vn6I2L6o
/+urZ3FRgSRHDxXhqpvu4etq8uk5UPBYRLpuZ3D6TSzy3e1rGtlj3zu2eAXMxCI4Dqa0xAkRIk8Z
fb3kPFd8DVRII/Rayh9G4jdCaWHKxY+KbikEGziZ1SXa+ckYEZH2P0iuEhJmr2RM+fj+CMytFAiZ
DipISRJC76hWDS5gU/Mrq6yQgXSAVtFP7Hy89q6Qqew4Tin0XKOTY2zkvK9daiDpLh/K5XdIH0Yj
R8uSwQt5FXPIoymjzBmvYItuZ6laXcDusi5SI4i0/Hhw4w3ccF47xfC12LR1J7L5tLAY7MJef3Iu
7p4IDWRRWf6aXZbgKlV/rs8OnnfO/xqKTXNhhLYqfJ208qFnu/2E86a4oVMluGfP/HoU4UHrMna8
FSUZbKHNmf6fCkx18jygesNvyIHnIUgGLu+J1C5AVYPIs1TC0G9uhIEqYk6J+n7so9TDb6OrPFHo
b7YIhNkveVCJrbuACxoTlqqoIQuehCpnkDf//AHQdaeSRdkHROjZQKe15WnWHBIJF8e+AQp5aaWE
7P7sZh3S4MvH/8RXBHJ0eOEr0oaJVEuidqhP/wnpbtRgzLBBsMTqATcA/hMFcq4qOob54KT5HoCk
Mlkt6s8pW/3TS5F+9z2x7Jr36545ll6KJfDoPAlcDnUTGAQilemuK2oMZ7FGyL3wvfiouLaOxAML
OdlEXguECrznUd/qquV/6s7u/R71etBuhtDkbE4TjhvC1T+OKv/RQhcVf2WCytRnR7Yh6YwGtqrA
vEzt+IqIecwCbIt0nFcVhGjmbsx06DockjTtJXkkYbhBLdYqhkMhbG3IErPQOr+nGgRBQcf7b95w
z8HUmDHhPABYwmeBIUZFKJ2I/rWiIKuEqp/l8B8lDKz9pLVIaLQaZVp7VyaUcIcrnfmuzeSfAam+
jx9rO5crqvb0CA9a24RyslSXqE9dxNGwQCY9PdbGT27xi/rGCCKMAPS8ae7Zgb3nJh05niXrA305
gpleOXOcVcakSEjww0NBqcVpHMd7UHPToivnGEr4vNk7kduj7qQAVRYH47iYG8TK9vW+RSnzYH17
yfaolAD6OUy2BrRXpwN4lcmkDy4X9z+zKNCk8ytutKjM4+Qy8z/BooLgDuI7Hg9hWmBwHcjfbx89
lscaU8UQWwxye8Pcafr2O4CTVSVvW5+HxY5GakqP90iGFpF4WhsuARJvpc2iP0JkTXi1yiihIMSv
/XOckGO/bq3Kr7upUpRbBxRj7rJ7qOaefhTQPBqOatyOGy1fIRW8XC+joq96uo8JLdAAH7R194x0
tKdhGyLHmLel4aMAQ4Azr8bFtYK2gn5X84iQ9ukddgsz4fbQ9E5BeuKbIrtmNTI5IiJDMERPLPli
vZq7daKMYXGtZx9nMZ/++T/t0V0IAK7F9/tm1jfkmxhnHuK76ejeJv+oKu8nZcUQPBttytutzVqJ
/igKL1jLxH4e5vynamVrBOmbUbaFZTje1Q2L1Rhi4Gib3CJc/L4xOUGQOkMhGlMplOXs6oLU4YqI
AzvjTG/5YzkY9InH4DjNExY20DRMbOD+XKNtTgf+s7P7e7a1Yl86Jef05AdvMN2ngCwGTLIdI9oA
Opsst1KhNVCti8HxrczqRdueRxyVjBhz8/KPFlm214pNeC2ZDAArJR5mRfq2gGxAsmPDIRtA2RzL
NgydFFqk49b2gRhmbscS2zD21SH+5xVVvhZe84v0GMWLYHnYUxxrkK1/2vOdYit0U27SBZ2Kedqk
ioRqrcLaQM6iTO2YNiY3ybbNJU+YIZSdAfkLSChAPHelvoC1dRR8SC8xAqGUsbEatOHlDXjaWBDq
HpzbAdY5/SDTBcz0jznwrURrBlmNi/JFsSx6aaxxGmuCEXB58FqzUhcrYlX9Xy6IaNzowDJdU7u6
TgVqz/Qr8/BPjLM7pY5dnEztze6m6K25i0uBI2es8yP2R2hC2ip08bJ9xH65lR7HlMGfheKuMTbx
JRayMG/fRLFr9wadXNcNi77GxJ7ebwRj8Mu7ID5SYCQLNyVadDPzaisYc4NOt+lCbCYQnE4f5gjy
KKcorFMskTIl7Kk1fzUU826lF7XBllDz/JsAaT2L6cekg0Sg0DDFB3dpXI1iI0my2BdSKokQsALZ
5ThWs1RJ1/h9QqGxo1CfhKSyg/7qebZnfYqwe2OsKQmkkh+FL3HM3odYnxUNFk1iHcio3asur9X0
JhekfpF9XDuH7/3HptXfiYy4n9gu+5RxleDd4Moh/Jz55We/g51+d3OoqL+g4ilVLw2VvXJRbfXm
PG4h3uJJV3XqfWcqP3SI3bKMvKPzJVkgWNT2BT8HURR9IwZJPtKLvIHP7Ap9CMblH7uR1sS5Pt67
Xayf5l2lfDMNExmkrtUvcHWYJsYDZPRl6wTufitmgVK6ncDVJutNe8sy5B2T+ECNjMbO7N1P9JxZ
ZY8Eq4RDl4/G5cWAolRAJM++5pmcjOHlGJ0ijrB1l0UgEUcrlhjhQ0n3X7kn1IHfbKZAbli6ZysG
BdHrPoCXdY687nZ09XCqmbw3lCmQ4kk0HX7IhmgfcbSsp0vZcHXdXwzW+MgUTdiNruqbe62XHeZu
UHejYpfXYg3cU8fDzTTqqhH9FIgAgZjQ8QeoE18jU0zti3g8uVVykxI8rh4TIKX8wK0YQaiFREbr
BHzXQ1r+2fE8uC/8Jj4VHjffR7vL4lw2VESC/0Xfm/qQTaqDN9mbg8tos4xvOAmWR/GPWLens0fU
LY1aPGQ3AEp/8KQLnOlE1KLX3K8uFE6oZehFCcLtoneiMoO4sg3q/RGoOQPbH3D3HYSozPCGV4aF
eDFkk8ecAtQfz4W/ZoXIGhHgh6OmmgR690OqePF5vaISWDihor1nRNg8Lvbkb05Xgu2gjAnsOCM2
D4DTlo131BUE/JshGzn78sX+gMtwQp8OduBncv/+mQJDiieLav/fluQwDLwL6cJXPfHF1/RZZGdz
y/359pfZyArIRTAq2/p8S4mi9ZrMgtByRz2q5AIENYq5IpMSOWGF9OLf0ykXNpU7bqBBdKiF6sO2
ZbotTfOaXQpqhcB+iwlpkkqfbsgDcAewcNIFBdtuJLTp9wMeS8mWlLEyuj5OdW0NMiaHLlHGeNR8
vrWWxqKANmZ8GouIjUW0ulJ3AIho4oMl0sbXqTMlWcDLZ7DqUObZziRiST0Z6Bwvbv7iYYIWS4CG
TQL5WavrMmEQiBnSm5zS4anCd9/dTCCpdZv+rzmKzJRPJvr2rvkQHNSku2gxtLvtiGaCZdhlp1Dl
lx4vSCNLHZaDPuAYxF+MSnDHIdshIdHRlEzGtcGrXPZufUZGfTIQsawB2jOMFwvKT7OA3uCtKgF0
KQx7+b3ppiEIZjBVJ5nmg9+XxC7te/CuEofxsNZCvMyAs7SY0joq5Sa4HLklGGQ9TIeqbFSIIdnv
swQ6B8w0pTG2TtPGNBoDhDWLKbQeTngBQFbaDnFLPrIXMklYR0Frb9jiuCanfi/ZrMVMZVxZyX0j
7lmGDZsEYaMomLA+WK/a+zk4V6yd/hG+wemaiOppfb+N3eicA8ZP434A/5opaqeiWeOQ5KbLeUW7
bpwUFnrEnNVuvt47ncdQlI/sY2rZ88BM+rh9+Zfx1g91PVxyxfrQQ/NQju+ypyZtfyofmrv4yYzr
UYJkqfyosX9yFm6oWDLC6VY03ZMc7WJNkqPppelTnZEo4CIrG3lq3vxg8lGdujwISqfqVs7V3NrP
WIzHKC/1BpWXf404DFy4QkZn1HZS5vnn/6Rqgm2INXjZRdEzEXw7kMvdNQJgpSdXw2swxoqw6B1K
pqlDj1VQ6PfjB61/hWZzwjseGmXt0uTmLt6BLOh1zgCoccEHqD+QRGD10POyEQQ2xvPa4GyYV+ff
Q+ofnMj4UvK9pQdc69AtD6jfVLgX6VH4HHqZCfE1KYWqx+ZNBB5YucDs7sXPQGz2WL2PSaF6MGWl
qn20ygu9H+KPxfH4yVJMFuNDkYm3d7f+nwg3k6Q3YifRTg30ffRu3bfaNRc9hevEfvR21ghypv9v
+HCzEmWGRe1ct0V/kXeDFqrHTA7MZ28WJk+embAggGVoJUWmWrG3IIUgAvW4ix3jrmmLQ+zAm+Oo
PqXfj+dH4LS4aZiTtjlIp5cBhc6wVBN5OlxkPqcL6g5EUMI045+sax5W33fEuUoKy5YAG/eKILTC
CTNFEwqbmKTUTHOuFfGDkOgpRiWl/RcCeVjlT1EHUZytvVWhtPaE0FNjR+f2RD1zEQS1U9gbJ49I
kHQOx+HZbO+ttxVOYykP5ZWOtILZb+0Cd2IDoEvzzLSA7Fu5jR5iQcw9IJvVmOU4z3SgTgVbkdI/
zB8uvl1UIFgSf7IRcWQPczgJQhtpe6RfzP4EdbtLwU9HwwsWnj+12KzvQKysdk6cA9fZV5e3V5/x
p3gQ/vLFhWvAtmRHqpujnaGDNhzefw4R95OIgVh3zVnm/29wR+b3SeAt8W2I6ASz1W9QAARwPK5G
0nqcEaXogn1ouDCaG/W/XjWHPrcXrggdXQD9R/VPGWWogUQNP6Kw7yTLbImJV7gDrlNnjILaMSBp
aMXC++NwHBMsARNO0+/Pj+MPqmYVKh2Vw+ySf166OBUmnigoWPAhXLhE924bj+be9oLaYjYL/+HJ
l5bbvYESy/A+sguAZnOyM6kG+LPOBdmVKGwQUTAwlNsOCtP7eo8meDGp3EaRuuNBp+SgE+LKpUZY
DpwEJoU5+xseccGjFQe5H+BERGM61/qYgZo4g0bOX/qrJXrI9BffpxjJhi23RcTqR3a2f8NRchy/
hIglVZvGZfwJ78FbxsRRJwVVHwWcZzxJmrJrLCnFmNlXPb9ELTDbSVklv9/7JuOYauV1DPLdSSSy
Ebbu6gvkryaMvD8X77JgY2Ot0ZUE9xPQGQ8UjP+kkKviJ6LHYMc8BXTItVk2jMyM86yH/i8xnm7O
cTnHXzwtrLgQ3GeW3Jwf6dWrU9Azt0jgp6k6HDVatQtiM3IenzyvZXpi2yZTNHPc8gZsuFgU8rdN
1aTSJ7U03JCVpEkIK2nwdQn/oUM2Ek9Cdq/CBbh4V9jREvNo3jEzfA8KUPusEdSwEKt7vcMKL86/
6qz+igVMxZ/Io5vEDHCocY79LcL8o5/9IXqugwiwMjfWxu8gm7WVGHvmloThjwjyxw8otg+GyHkv
7p5IkgUnLUJYJE75XuqfWH5lG9NbGQiGB4oz3HwnskX9GGp0p+0sG+Kl14hZ2M5gOc17c4J4NEWW
CcNvkJ8A1oMzmxMuqbY1ij2zgyzbrW/EBnUxZc50IAPzyK7WxXXmRz7hWcRZZNH6waCDsgFyuWZN
YpyGj6T7JBc38yROO2e0v/AJGW1MlTRgve6ci32uvycZKqwy5lVADOlHqD1uIaRFA0AzaTWu8Auh
jnPGvm7W9l/D0GLg2xqNBCwonlZ5nktlLqxW830jzPQl9f5TciQMUfSVsfFdxQjlOSM1o1Yntt0l
L0FMtLP9iiEZe3F9faMDDanAQc8KYQ57dNSSScQVX8QxwPlSkdpeFlOXmJT/VEGezKB39N6v2ob9
4776uMtuKsqT2pCGYruob9rvl4W71YY0yw3KJ4dWyzrucnJdHbL9ZPN/c4MlWH/DBR78WzglySkW
/Fz+TQ/K5PZtAMbO6PDEsZCIiENqXZxgmDnVTLuhVxExiVexK9IqsGKgAZDijJx9b504ji59clrC
o84bJrMlEjO0fkxlrqDS4IPHBPP+yBgVU6Ww6LGT/1f1Kgh8kucKCSONqjbNAMM4YMPN8cpHXEqY
BQI8FQ4zvqA5DvofmBH9EWuu8EBsPm4vN7AaqCITUYExEujXA1QTaovduWUNfsqTYND2W34uCscs
8AZyxQFRLQCNHvyP6Ptt+cMEp39G5Fepko116d0NMOLfv86jZZryL+BeQODEYWSN+sjrmMMjVAyr
SzM52MCrOlujaIaOWIr4htNJhAfEZd1ZRVURFoSRp/jfCSRD85ct7t+RGvjmwW2T79TlLPIxmtwn
TC5XQx0PGjNdSqS9a8TK5lV3HNjmvNtpMQ2CZHNHeIapXnJVMnD0wVLsoAcPAavk7zNO6T74n37r
rEuocML+2dGM+QwopCrYXIM5yp0CMZHxZIhzoUqzu4DBHA1bNzRnjAiLt7EHHV9SvsC3vxzwolu5
vlc+8NL5Dw7YO7KAgRqLILZwof/NPjXIEeDshB5SrGV4U1khK8aT1DF/irqdwxB+nk35UYRTLloW
3VWNzRHBHXvon4F4FyKAx7pSTyYZ0ajQdbqYxAYOOU0TsiuEdW4xMyl03+efzJFFTBbXjgNrGgd7
ckMTtET3Kqz4NLdE+6QOrmP3hShy/DyLEBpDAnJ2E4cNJuv5Uno9//wLaQ7x1sTdv1Koho815W26
nDY9mqWOqujVKClP/6mOA0jMul+Jc3mtgWiRUGCPhKm33BgT3XfiINzq6TnpTS4sEfuSH46oO0X3
JfXszJcXNATs3SHVoANiK8pDg1dA9rzzTgFXjc++2KX0oqFm7vNzznDT5KchnGEJ+l76IFwvp0jR
kHPI4/n2t4Z7FBTPm9hJqEW4ToTIJlh64EccmGV0TO/ZQtvpeBg5UvN766lhIVcLHjMFSJ3t15/L
63XYf/2HUkatGMWO9K7feRIoFa78daR2S0DR6oXOr+X4lfjHFPtdAqXDZMTX3pWZ/KDdrL4eFlxV
r9sQY564kolZCqqPyPJ+3yzSuDIt/ysSbzjp61TByg97enZXXAHjaIicihvbsiXci0Gkd6wkUbcY
yy3BK38AK5H4NCa0isPMftN15Xfkfs+vIxuaIxQrgwksyJPDoGrXgJ5pvPsFfvD2E5hvn9ZxQqpj
vAw2/7TWy2RRxqVIf7JgbGyiciNCY54GYpLVxVSh3E7HX4y4oGmvN/UogHsNh91wtJKoiiDnn8M0
4IB06zAO1MLgQBXhFWegs57czzDq6UR77r4zKUnNmdWTkBXtrTuGEVt3OeI5BOgR1SgY5YUNi/h8
WVZhACh5v6fKkRN146qKzpuylVAhzWxiTiRkHMjjX9RjSrhTIQbO66VYf5GXXrzCQgukRI387D6g
16nHMAnXBWl+iOd284JjQyDa/z8GE5ehv+wjeJn/dIGt+SHhBQpA31YkvRjXUrAoP+ZJsNNgcDhV
nMOSZ5nIFaersd5o2/UFG+4GtMpzfLwyWFUPOwRiRyfJHJQvTeDEU1oiUBrPM+RUQ+WXCvhAOseV
bQBwZHzyRQl0g0asclOSsWWVJ78OccJHEo3RIqSRQq4ddRGbbcbqsNJ4t9RZP3dDNYzfVXs3HQPj
Olat5ojQjFVZOmtUB8S2Xf5JRlMZ2+LR8MMDK8fcm+EszAvDkewtkwTdNdhuhX0GArt4O28ZYiX9
RdIRveCVZF02lnbz823zRjZhwNI5qoUwicIhTkZ5r/cGehyOGJ9xBqYlgZIOPcQj+Vj2nR6SbqP6
GFYAYyvzhh8JmDHxQcY+awNCbCcTR/Of8psv+Rj4NadtUZzRGmfyRVKVl0/BdS3oXOev1mR6KKgB
oDT9f7t84B+vzlwnso4ueB4wME+p4us0PuYbUDgsTs17vn7N8CnC/OIseb4K9cRJo/rWBRsVVt7l
+CaAP3RdLn/qrmOecErEBcphMSotE1GVrq382SSvK3fWmQMColWcCJUJmHHgZpRYMEgG5ohQdpFd
92C1tZl3ZYu2b0XCLVvcLrjaLliNu2/T9wWTTO1Qc2FrIxJ/0mzQ/siLvHwfCZqNTjkiO7erLXir
99/ypn3zmQgCtjUKEAgPa8x6PjCyKJF1OwsvF5IisXLWWs8tWJZiSGalQvOH8Y4MculPCM6bSVe9
2QLbTHg2Ubi0IWsyHOt0BRCHo6Og7eCTAmyZeWVRJ/+zQo88CASdQHmUpKSBGtdZrPTdkhQ9Zchg
mJhOrfllBb/l75hQhHAOVPck1uBuB8OoR5jWtoPQ8yvJwARQQDBXp+R03oHte+8hD96bB5yMya8n
JcxcsLFza5I4Kn++2izMP9ss5+xl+sq48LSM0bKFZ3wmbA6bynldCiDCQO/d+AIdgcmkCgtPpUaI
qrn9PtVkg8M4tPsZMb4VBdDUiaqqC/LopxahixRtuJdYopYvz4o9xfvQG6STxYYjdh3hC7FGn989
F1mPU7VQ5XJwGqAJgkkKprXN+ngzn/aCaMd+biOnsZNpDxu0JlswTFSCPKXedFd87PHAORATtPiy
FdJdvAc409YfdMmwf94i37Wva+z8Qrv8PZgDPFo+0Wvcok9C70dgNo4IkOGJoHXDaYkhkn8ncA47
voR6B451a+YJx13cfP1R007l64R7EYNikHAdt4cI8Rxt76fTyhnQqwN+2IIVGGaFVQ83V3XIbjyn
v/T65whdByOTTar73f69113Gk7F7Szjdvjl+d3Io8FnOXYgBiC/YF4j/dHYhX0e6TeUTSG2TSYaX
OW4BlBBZ1WLsFqon9T5Rm/U2tWgMKLsmpAxY21dUZ0PTrPUKzgZFfrSfNlMrzroUCyjra/FyBt1N
qVgx4GnJu5h26EsYaN+TelTNZJ30Fopx8Wa0vZDxDw//azu7oLIJyk0+vjh2G4WLkTy7tK+ET+gW
nhtA5swYH1byniRt73Om5Xlg/5+ibtJv5Zp1QARTOZF9VM2e0UYDjhd9LOq7qPd7pUqSHQTqrtJ5
QO9TwktXILFDnLwA7LrMLg/Ow2Zr//i0reb9O+iKbg45CuLFMc/ZjmIquvm0pvLYo14HMnZOLrdR
/y7SnoT84a3LAgdzwAxsQdAIm+8d3bT8svRg8C9DGSSU/ApLuxsq6gA3aA1aDjdLtPxhlB2aW39p
7JZtvb2y3i9nw51iybvOpNaMhZ0OjjHY+1kxg2oWip7Z/iVFRAkc9h8yOp5sqFlf8KuAlR0Uqr1f
MyENUTQjJ94Doi5bpz8LXAghZVuR+naL1MH149iMyGTaPPw1kHZVxd5TuNCizsZ3vOBHJ89wp6I4
tlO3LczYHa8rludXPg1sA4wNC2V6rC4Med6aaOHvFxKbQNFSpz8ADEACUJTQl4EvnBnD5CbTlJ/M
TS33el6L3XYzcqgrV9w5m28QJL3y78o/QWcBdlYct9GGR9weqP8LPFyjtCY97/Sqv5rl/OenxeL0
1c8NT2nMvPQW/5MUaSogq0ejL7jBPspbRJ8n6+96PUIYQW6cISX12ERPCE3wkel1xUCU1gCEWqiE
JUkaiWgyEb+PfY7IhPortdnrgGi5AaaS+a7K/WFubyCMWxgjOPrO1VFlj2mThIYTJ/BA42Tr4s8Z
22/Ov8oWXJraLh8e37SY+VamQOqrbIhMpQkgdN+sb9w+uAVS4I5z17TAwNrOCoCYrrne5MomICpm
Pk8cSV/7k6a2zz++B3YLOOe1TKonEkCDaBx+xgHT5c5tE/2pSI2W4xGIJtRbq3RLBXszhKi/4+F+
epJr6L1KVDjF/BXUpasCrSwwQ1TrylhUQvzGWkWai0S9OE4pVku8/N05eK/aKcoTp5zJnSHweOln
AHBIHBti1YNwax+K7jWCgZ9YWmcKTp/WmwF3eHWvXetaKPZa19QbH9w1yLkBfBEfps+W8hmR8/Bx
hbDMm1PdwM2G/+llRnFs1Zv6KTY3B4j5ljjNs4CuGmgjtogJ/xORGWn+16aK6H0TDpkrzAY0Tkj6
poFO0efuynMw0Z5aDElxy9hxI8hmClF9RG/8r5TdcanQeAFIg6CPCe9SBvD2EfH82tWGCobfBFPo
2ayK1RPnzNDPo1+0GNcQ0cckdofVw8/EuGdI9d2bM4f52PaPelGhIxoO30YY+oMiS9gZ3yd5LasL
j/33S7SMTPhnkKoGpGMgoj8qHtsQNjZuda/OyIYVaEDfg18BIpNT3ns/uQpu77YKvir57fe9L4xK
Qki0evJq/osz0vBkDDeYmg/A7fgv4c/vAZFc/W8S0K7kgUSbE3qSBgvSDnS1w2Rsss9wBkWt1jTr
eFu93pRXZ5QPjy71/nLuM5kjZBmf9xhYl+m2/CBzhPi568C0L9vc2Pvwj3u1BsPhFHYBm4l3emKF
tq1fP62JsRpLbhBXdTJaUnnegjyNG16UUeQKOtQwNswNk/7Un5YKVwlc0xtmXu160fPi4QapeTY0
9z7pBsMCYgMLhgmJ5t2cj7K7llZrF0SlAyv2RYu9CMWV6J3K6usDdKBJt/4DcWpFDThTFlFG4S5s
qS9v4h7yp1kx8KORLHv3lTT4zJpdDp20e5v01JlpAXzALZKmOa3Ryxbm7m9p3L6xChyIW/PIdbvk
FD6xb7Wow+flFPm0Rez1mNP0Pf6zD7MAGPBVMZNCCYG8LccQi3xxnp7nbTrqeF5CA1X7LTf6/9H3
KmKIOXuQkPyULykHFeMwYIQovmBbUOoyMRqYfijnB2EynH1acv0XEdWbhUOPHU0chpQEnq3uOK8E
vLyBfD7JGFID5ZnxzuBPKWhdtnGpEvYzHtdXcnip1FZFFu/0TqHbOR+ZU4FxzpXstacfvcivuNe4
6go+BKnbG07YnbsBMcZioJTBvDKlsND09fjjQ8hYAY/ZWHws3wPdBVpCcjYaI0iLRjcnqIvIfqdK
F2ftFvdJ2pt8eoAMQQGf+lAqpX8u8wyBKpw6+MrA9tepJ9tStufE10XVTbReK9llqckSNnIYYg6u
kGqbL7LQycS/SFBRi1WTabbDUCCYWQuABd42O9vovmEH8YjkKb5fa+ma/SU8yR9q5O/goAc9Aqq7
u5Rr3+MENoGlD8nTCDY6lF7B6uOyhNz4nzwxYrkryDpT8eSqoMJh1UG45UOpFG07MaWndiEDbdmF
iN48RaquOMLocIUyiqws23vytEOFwUDcJlfV+PRShO3y60mjfvnh5K7DdaVIubmas8ll/2YvFXSs
X249aTuDICrDm6sW+3i7Z7Oq9vkZUCcHQdTEEdYu0/UBsomtKJF59LK5psOIRPVFisisO0v/iLxo
E+xuaoAnzE47ANyLelk3h7uNIqTeTqzkmwgs4at9qp1QdbyzQwVLP+sE7zMAzli4zH5VrsjYr/zH
qf92IzatuUAg02q5GKlwVPZDILPY6SS8GFlWgDXtLFuk/57ehxvvsEGuL4n5FQWP4iDrVQiDyFRX
WQ+GE5tVe6N7bsRWOcRM3U8mYyWFVscOnJXAdYNjA4NX/u60Z6znVuB+e9PBZZAm9VrJUToffH5p
PTFej+6M4YM76GMPoHOf/mWrAw8GUO3PJh0d1S0G8HzWHzx17O0PS0RjRhiNVwl2FiMrp0R/l4JH
Bp5/NUZ3tmWU8h+u0Hh3FMCIAqAJ3wIhM7Ys66Dj/Um+xF757SlJlmedCzW57Ts5PIqypwA7oI3N
n87UDe6VhK+PTMjSb+DZz8tv7Svs6RG2WeqFKYxOS5jG8PcTYqJ8gepf2S9qLAT01uwpdioqVy29
+lsEvXGu/SwaAYWtA8EdEx6FqwhTr27XiXDTZ2xQ2LDXkZSMGcO7DxUC0IuGF0L5hOf5Y1hxP52m
5n1EHyndGUzyAopDVx9wM+8Iy6RmXoAKuGa3DIWNpv0/V9uW8fa7kCM6NQ7HXhC55KoUxsvNegHB
4omymom4MYV0dTmjWC3xKriFaC0wrAWo70MTNjsaNnmgTXTjmI8ykmlg+G1h6de+R+4daU+yPB8k
FFX1RZiaQLAkiWSI1F1ukVLCHEUodQAZ8o0JnXhNMv8bZDoAH/rhgN82K8k/emFu7JOuKeSk9W6Q
EOiy2m9bJ6XYCVg9m9jGDtDhnmX3K5yvUB9nC1QYzlb+k0uVxyCUMBHZE3wtLdXLxF7bzMfXzOAS
g8QehKczn4cYvaU4p3iEFYABwyUNu8e2dAqi+Zr7G6zLeTXkp8XOKM30t9SvmyddsGMKtYdXj2TP
B/pjuVXsxvZ1RPvZo2DCK5hy5bva01rcqilF2ZQdMWmUD6EEAmhvFlRanmXm5rxrMmjrmaz849lT
GymQgAHppHm6dfUykg25F28iajEyz2ZQ1B+NM3THsgTTLVdsEak8frlY3187oSg/ZhJnhmzcwNpc
Ze3jDaiFsolqn2kxCIPsB2/JFz1p2KyaNFzZAgs6J9W2Zdpl4mgeaP10qaBHmdjJyF5SITtwfYBS
aoQjQHuwNOBij0xfc5lbTXX0MDOnsmHa6wdb+xszjh8P3gdPsRpjVoV97sSVRdGQKDd34iTmK0Fg
jw8sLSicPl0BQT4tS5LYLZcuYCel7oF2FFiQVCQgL8m/easAJRI+mWxeTLR1PhY/bg0OSmQm5087
p6Eho/r6lrLrUMJWO9q00Wsl1jUyOedYVmkj+TDCbulIubT+QudLs2dieMz3hXqurSErVmay6gQ5
ssy0WSaqwS8wzS22tPWpokymhrZ26m4MM8r7Jdj3zz5i4+X5fr7V6+7mNp2AffP2B1/4oiYDXZbK
J7hZAmSQ9d+YlfcaD5Z73YrHI8c3hFryESW8/3TxXy0PcdcWGL745hn4rddL+AWJnjrHqppRgURF
hzmzn2Zp7Oi4zZUPpLQ/pum/SeKAqzLhr7Y4/NW+Y5snPEye8q1dmcTD/QCEoOj6SVzsBk2hb2le
BtU5wE0xmWktxVqZU17Ibc+naVAcQb3ThYPoTxZ4zquSD8/eichSkae9lza3lBTuW8xd2h02lcbE
W1HcyrZFXoHVXTS3F1qVQyW+V6VgcBHRzBv+7MEygutcwCjPl/Ooco94jVodmQABK35QyjWluYg4
gASUou+h0CohKMlgrF4fSnjox/0v8DXfIlPfqLD1k1VglXquumpWI+Sxb3S/fDaMfKudIcjrTBi0
MMStNmTeJk6rCenJ597Ao3HOFfzgQ2jIC/30RxKi7UH3vdSSjD7G+zIJ1Cp6Cmb3c+lbpkYET2PG
q7UH5OH7Q4m1qSptMNLlmH2pNl5NRROt7a0pW/fiO26x9BMGos3MKq1tjWbVGsJASjPOFmDOT6SY
DA75nw07oWTspKAc5u90EJX1/Na7Xo0T90z0sCv1mAOGK80HH4GLkTbh7vQyI5PSOQTtDD9QjsN9
NKjIM7w6xI68ZmN6o2XY+CmZt7TyuvQUFz9S4w7u85gfrGhSRlY3cZYZGm34UaGtouCJnB8WP7dz
NNSJwyoMlnV31Tny7LZKJoqFOWRzX2NZ+VlzrN3/+TjybLE53pOp/iDRXQVJerfgkDrlJCHT6EHq
DYkJdc9oj2vGX2mJh+JVr/Zphfy8js80pOHYHq47qr4CA18J0VQhGyU7hLL7H1X5rQzcjRG9vYZD
I54H0WiBf+JW5VYj2LtkgKWEOI0EvakYUQ4nmhmc1rpYpBD7Zk0Ifcni62jtCbV0kFIx3ST1RHwb
ucAW9ZvXW0VlYJr3eV2i+HttSOlSQsZyAEWTP73IA633MemnWW9mPWgA+A7YuAEJk3RNG5Yp8TU2
VrV9kRB8Swb1IfrV1OEOEhqryTWWQKXERHrR2KhI8ubUcuOX6tsir6PH/1iYkshqFCQOVImamYsX
rtzfsQMqbAwndwPyNWgHlslPxE9JFCgrIGHYzZUDxcWNd2jwg47ND1xe83RkJz/kaQYcqud/URqn
ktHIj6MmL4QPKLC36NsBLwkIMyNsk8N+NqwoFX8GYUmz/WKnUcdTb1y/Br0q8VdtIpiG3nUYgzHz
fWBAK2RODRmn5Q5zyyluboSe2t5BPs44iu7lpPpmScwV1qKQujzuQtJvB9rDse6tl1MnNVY6Neit
pLy53k3Ixm8eh5YTx2/LOQo95S6rqQ0SMU6adtMvoeXo4o8qbNU3urvgItX+KKTiOuMC/TGVVs1K
ITAgbMhzgSQjSpZ2OeZKy0zM9fqQnSdykY0xKwQc+b2zMX/aQjBVfc1iPsTkkcTxsKIkRwwEnu+k
wDlWDFc7CnToQ1aQ71gQDPMlEKZLDLi0W1lDtjI0dz8Dtw5qKdPtAq7IKJNJabtp7xv8vSskaZdW
Psz+OpUu6koYUjbT/dp1v9EH4Da1l+SaDNRyPpdINfeNfUY3PqXOEC6CWsXA+I2VXK+NRWGo3+vE
eXuIH5kPcH8vi7HjN9sgJiuBm+m0Jo5UBTDOddNxKsEyfBGy0GfUJI6A2MuWMmJhVPQ9yQitG+QH
kLDlc7m+mnGbBxhS8MVgVU18rpkZ5RsMDW5+RISsIRKoaij4vC+56mkYOClsqg2qh8iMiljQkGU/
n2xbez/2ePNLZ2FHwF3gwZeSKup++XMm8TqQDMnlhT0j/Q9/uNz+RGA/TQi4E5LOfoJ3OAIk0hbV
kF0/DtI9Ro7Mo/8aLvQvRyv86PC/C/gDAYeiuSxBs2vbl1MwBxGbrjOcpafgbUFo90HcESdqsCZB
aBN9F40kleRhYVAknSXN/NE3pb7KWfzjO8+bnLmd0KzpBcrBLb0wW/QC/EEuiFsK1QyKc5l8phqh
G33TJepFc4DbS9jBkufYvzlCYfMs2O3fFhcqCgn0eQweUb3iMBTCnHCykqTRL7wxEQtxNyQdyX7D
M3O7aylGXYS+ytLKUbczBWguQ/wjO4wEKr/40+4WsAK3YSkmXwDqYfWkv+nntnHvCIJ9LSt2k/o4
chiUfubkiYVpH0NKj/hAV8kA9ZGHgxdEtmUL6OeAPZbK7jOEcwxJPAwQ8KulKxMNW3lGLLMNamv8
TOfB0x+5o2CGa2x4ogmKjE1d5ORhiK8kIyBXfLxbcEQQdM9VEyFTH0DEZ70lryKB/IJA7oIBo0iH
lEi34lU2gaw6LB9F/zg+zxyl4WXr9wqhgIkSEWAT8VC7d2x9SM0bbvPWS0msyz6CGQzzXqj0t9Wt
Ei6hxRbiWrR9YqLif3AacRwcwjXCHsgzzFqu4NjPhbZ5DLT+rtjoA/HGLBPYvOFdnai3arB/UUKX
RkWq8o0gQ4plS2ifKDfxW4L0h0BGg3vBVK5gez9OcSxwzvZqN7nFOtE9TI1MHfTjK5ov6Su7UicG
AAQLMCWEc5RMqUjVRHQvmNAMC6sVL1meo+v3UrN0rX1xSYTVEZVUi85sj+2Ob9+4HRY26jCEdia1
yRb3ntnstr0ASeweXApMygCRZJxKSrenfhgE8EltqAQhkPFBKZ3ABcodjigqqxYgKXpZ3v1RTZIo
mfDze2IBwYTN5e35kVIiyntxdub9atEqIXJFOTSrihlCKdI2s++KRw+FwhZFWsbGB0WrHuUJMoFU
2ab+8AA6HhXwpE4XNBdwSMLkkhmzK7HTmhn2t1y13SxkJBdHq7DjRoLgA0+bqcYvthpD1IjX/zta
KQBhL5ODH8g85Zq9+XrZf/g9yQpMk2QitK+xW8+P9uIVzvCxTnRz3f7WOSftbA9p4Lzi37OplZNC
jr/SNpfCwaPL/XGzTsjDgibeHHddHg3aI7Z1cpvYdCh+5P23V324zVxRrGqw1XvrHAHO0DFTSddp
Y4zabQ4IvYgot2OlHgqKqkGDWkJMatchXDpCBiI/YYDaGo5dLzitYR+g4ymUFjGtfN4AyesCaqxb
HdmwqrzY8wjT2o759dNYqJH9uvSDmgYSCcv5T8BQpxkkCRsI88cAx24QS+zc+13bP83sr0L+Ztr+
b3UvXDinwqPbE1SrKKte1qBib+YnHnCJ32Lp+qcyRYdfCbpzpkHtmrXnlfDH82vTWVTGozllB/I5
3eafvkT2iKexLcD5qQjTctHKrkuqXgBUXA+plJ8eueEGwE85l3BD5X5k5Rw8nyjG2wV7/hsursDN
8vWeHSYqOeiptfIuluWd1lR4iWwtnYJgkGoYEW2WU+L1+1kmjsi9xew/uFscEOi+eUzVUabGM742
FH7/8ep4ygyrm+OJ0gI/7iH+vAJL9rBz1xLPQzGXY7pGeqP1MMPWK+sL/wTFNDzm4Ub7puS6AvBG
2CwfiJ9vbXKc79KunaChPusoTg8XuKE6pXps/SoePCXcMuKeUGM+NPanlyXu/32J6SfCipcMZzBR
Ep945r+509uM9c7asQk9j2QXJQnAQIe8QsSrzs2PoSJcOV+QT0caCnojzKsiUHZmGm1pNQiQTrU9
YbXbqDg4VB1LZoZ53Un5Orj9/pIgfPIm/4qa7uJKWuhoiysBuhbu+p8WO39NxAWZq/ZaRdTMC5Ta
Wq4safMU9+VRYvgs3Qioymw5CGClE4sP0tqIvYTCkRhiMkkrxZl7Uso2nX9HS5SIbSDvZQRJiqgA
GCr/ZATlscXgxJUGAejnAJNerfMK92F2DHuJ301q2LOtg6enrsRdf0wIgZc4W7/Hnhbzs033H3Bm
MNwNvkoplVUym6IA9C+60DscBVDHcKyAMphXLBAMOQ+Lv+8VZhsCyppKLMgg0vFvAgKDIs2bNIIn
sD2CqEQyZH6lyptiFbuNPyDecLY5G4P7eUiZug1xGt8qOJ2Q/POYJnXpGRlb6E8ByIG7YnFxYclu
wVmk0nRHW8ge4rNbmx/pdA/yq69UcCbGQQuUDdI/aT1sKUn9eyjzNPl7Yuk7eDBry318tSeAOOCj
Ov2xJ9sbsQSahDVkMpxielt/noMhpGFnWY648xdxCVbVeY32jWOMSskCefFYuwj7ycjqK2AF2NGo
EsBtjr+ElIPftlXMQmwF/MyhhE/DalDcBvWd1nwvtlpTPpkqPEwlEaqwZz0JQZInbVJ54ny0HaHj
CVSxvwj8H/PSBiu1Md82BxXVF4MTyTHeRBFS/xetQGpK9mz5i/CajudJ9NilQdsB8MEaXQtxC3RS
08UtC3FueiXWphyPkWxBsp9qjcxcFqTMdGEj6UQ96LHua2dxotsW/3HCmMYtsEQJuARZW+NF4Ob/
yxyvlOce/C596IKd5Dp2JvB4eGU86s6dU9uC0Si9mbty49VOS/dYXAKTlcABWbh1cm+J+o3CFUos
Re+sl6RF1z4eZORnzEJnIQ2bJBNDtCwqeGjH0vJTi/qgWz7sR613DWzaOrqE/gzxFSkYfTW3Ej0R
ylmdtFIacAfqoNhTdY9lAhYe98un+bxeip/+swnzTWAO4vYUeak/R8kQ8CrQ8RlV2sicGHT5N9SB
cn35ZaRwD3WykjfYauVa0Jc83lhFRmrnN3/KqZYI5YeXNbXOnY3XzyvzRrEYzR92TWeBVQnGPY2E
UUcvXyBFFNlO8Y9O47fsu82mxhFT07kbEhX1rImewt5XWi9U8vEM6P9L0pfc7EZpwPwPGRhUut1m
FKPd1hYGc3bX3xA631VTHPtHXG6r8N7IMpK0AvKUeJauEWPORO7CiZAWza9oordZeMAfnSps0r6l
4FXuZpdWzL/IvajYTa4kWEFfAOiFLAc8tF8RfI3LXegV/TczkEi5E83cQV78T6AeisXWKWrpkggO
WIhuVdkNgXfbdXvHgYDQjCD3rNpwBlw+Hp+tPnLgT0wl1BZOIX4arGs1FWUIOyAuPJs0zrF31MKH
hN4QqlF/g732IxcVS89fb7D3NZbnKJkX7gDVrRL9rHu36l9/ALe3SfFB1aZ+LDhBMXi7i09KAWHr
SekHyqLL+mlj3IluvWKKSQOZ3sZYfxpcB9hvC/vkb6ZbaEcAfzidWJT1QRvrNyYSU+uPIyMKrQ6L
YuLj4Cqo2hK3cJ4YZH7d2r6MWox2WOIrE49d2+VDz6X/iBHDxq+SK7PS6DOoD+86FDI/OdsMio8p
2GIXq98QAjkrsjBWVJ7njI2+Y/vSgJ3KTB+TXQlM0YLgx3LffZ8nFx182Ykn0TOq/mDvERsjYYs1
XnCYcwAwwUSk9WSmWg1AnrCZ1+ezUQ/gwu/+WHe066r9IX4WHBWUlxwRwocj3X9xlwq74llXGLIK
SQiu+FPhyFMPrcGZvbUA+z+B0RLwYWtoZcwsFc/AoqDmOWfXRWtK8qlZsVWS0jnYxWBnwd71Gfwo
Vs2LsmqAMvDFeVs4+b5nJ3htGem7yPNibWuNNM+uGnOuKnq0N+tqHHJtS5lHSKntIZWARwGk3EO4
ynCEfDPTwc6N7xfCVGhOsxbSgfBJfSigDL8puKGJsUre6yerj7y/A1tK1BgasMA6Qks9ghcu+Wlg
6HJOvVwOWU5GzsHq1ZwH5GBTOBpFu19NErSnTLS6AE+C7q/7obM+73FQXHbTOkNZ3gDSIFyoV59v
QsRRe3lFPecwJMdHsd8kc2x6AArKM6EN0XPDTcwxCbfpDQ7CTg5U2SW8ZUjWJnT1PZrPbILWFrkl
Tn6irowq29BLIkoKpOu6BP92OeTI0yvUvgpFb6Uaw/8QwfdRZO7F/0tAGyiykNQIACqnc0PiCVJI
0EjeXxyEDcHF063/sc1pI0+WFYIaY0FvSGBFEngEdKVlBVyMC/IzMJQ9W7joz+XC3dkO7LT+TBul
eFy+UeOeILdmDJN30zrDzlGaJiGVwVLX/byGZKyu4/P3vgr9muhloNYI0s9vZswtz+0T6u1Xnqvb
Iw/kgB8cpHyA7SuUuII8xQjhnC+Q0tS5mqyJrfkuANcQJU6KcueP/S7qofE55QGjdJGv9vMsebk0
RcVDeAzeA6QpC7ZpHvzLiNUCc7RzRTW1aKjMgTFuQNKGfkaQbFqVXMSDTtIPSI6qziCiKiZNvsJc
CeQGQJVnY/QuHmRXUeO9WzgM80pu4Z7/wEDjQJaG02Q9fYPMNBNUoHxCjcLKmMXcSQJxM7sgFEyv
S/6FEBTI7kjcAa0YSh1n3rtNej6D9S7UEn2PiHz3Atg2bTAV63mjnhhWX8ezRcaCdX1drgE5OQYn
xJ+CLUHAXiQrSXU0ZQ0q51qeNC6qzdohBIex7YIuvJhgUWpm26V6Tr8yysLlPE9irPgLILn/WuOl
8NE/wMECUrUxsDmx9EP3+Qdt8UY+62auY40JRUQZOqnZGxEVo/Ud4lmWTYgSTHli/KbPJQ+tEM1k
5TOKCIQGtm6Fx20OASUhw7yJwBg26SDONkvFyv34a8pgdUUWvYgWEfzVG1xZTFES93mQZWXgu4cO
I8HwIoT+s67bYw5OzoOWI/mfmfBIIlS4+8PHI5o2Q1gCMESFqo5HgckuEtVgy3OoDNz9LmnBb3+7
H8HBR6aedqtxG3oo4xWtR+rg45hJ2EWECejt7ktYRhtCz9urTMKy3bxBFaDhwy/7hRh8KLNhlZgn
VjkxLUND2vgRYN/8QIMNPi1/fr9l50XCpNrygPC5B2rcwAZ6ZAA4jsJLc8SYj9rfd2WnpRhDzITd
Yn42gsbtHlsUScn2lJmhUlC6J3xu5z6+/KtI7Yn3tm5+oxSBkzIN2RydsjQLxpltuAi69oU82vGy
Lty9NvgM0LB5587RVnoIvQQXvu1ClU5DDjJhaOhzET2+4Diz0/yUPqghKdJXj38AeAbSjSDVeAY5
iouwlM5ieFbnsYGLRwHhYCfgwh5Y+Zi18yEJUYUdtAOovV7+ihJZZP+tfkDAI/qBvZOTSx7uwN8F
EOQVvuHMvYH1kf0VZ6iQMbNllGdgjC1lEBFls+ihgdTz69DhzLvWbkQDr58Zd3sHIub8wTDtPaWY
1vpli+17LO2mqkhI2RByYawobx9EAPI1EnSfe4XwriYPFbYJeZDd7UW2AupKeMUAvNhBQHlswtCY
KS3kHJ7obOG0hoza10A+i7vMuo5Oh8oaJJsnlJ1DnWMgQRM66AgUfXzE5LMl7xJmeVqSNl6qjfJ/
UeExriu4oS3p0RY3Vrjlqbjt3SI+mCSFPzhVyMUUql4LFhEP38LebejRg0Bp+7tqRaQSQJROuGJa
6YKG4KoJtnmYbje2Prw8Yq4d68lY2JFSm5W2s84ED2xcj2AWX4oH99/wKy6qWpTPFQ9k6yQVEf86
b2H/gPgWsQYrpRryEkCmZKP+PM0Ahu51IrolXGVhlbjPLAhma7i3BHY9jmBrOUcFIVRBdPE10c5c
gQizmlm39kNoN4FP8nOaW2jUrrpG6f8Np6EZ7+bsKMZQkLH7SWvKqL9vHexDlucQboQrnQKj6F6V
0zOeCYTL9DSofG8bMIWsCuTEUfh7jNR9Nh1B2t0cgAdeXtx3qM3N+8E371Yi1NU1bEyHMjGuwkb/
uBV/rh2XgvXhEGSHW4wjXdJdK9FAMHWMThMO4urzNNh+ACqoKkVIVJkTFQYvF5qt0Ye41j72boAa
gHpe6v6Esw19s+hBkC7MwUFG3UuvMQewVjQIKJjD2wB64w0iqBRl5QxM4H5GRcHT2+/y7CqjHEY3
46xWFkpT4SxPm6xmYc7oIkBHr/1CitrppjAJdxlVtWNoqjfHLrMF9q96x+u9/wudmQ8Vf3btUgHB
few3OtF5FjPrnPTVDkFORh0QIe5BrMpjMmKh3kmpoGUYYtxFWhONulu7uiuBZxcaD81lhai5Zp8a
p459ZvIzCUIkcw0/u9zKqmNIy5Bax1D7AGYTjTS16AbFx+VnzsXmBWabwy9ohGKLfkP3NQmazK9o
ZoHhJZT9tfZdvI1yfkUvWT8qi2vbn9TyQs1OoK3nT+Dj727cu25+4b0iUiH6GRaPTJk0Vdp/tXd0
vQ0XyvzzSVeahpb5/ELyUrn8EHGYVyoyMrl3FwCRIt2DaOMK9F9sYnlDPErFuyOT9eBdEMk3cJnL
Jv03L1X2I/T8Gk9RZXqDFW9SNhDtWLOXL3+iHUupztnghYrqYOs/Ei/f8ewcKpUBVVYN0ZAvCJsH
gbHrkZ69cv33zlNYNFruV6+pub9sSuMEREG6zua9R3epYGlyjIUljXtgsypMx4QYZ2V5WprNm4df
JGfNc06T07L7p7IB50yNrLCvoFE512dI5aXT8eKgWCGWYDgqFi7U5mZY5z8001/9qXbc6Vawr34C
Kh/y4krccidawmCD/9tC7XAJ+3bYIwp8v+HeJNQrcOl+jZZWc/AxcPlVEOSVA+o3sjjGNMr9XyfS
2Yo9HarVhyMzATW/eiwj0efDVDA89IG+U1mxV6YjDVw2MTg3q1XGlTJsMd37NXa2haX+v9NUi3F9
A5MOXDWzUyNIrt9Uc3yCR6YfVUooHBykQWPl58gNVj9WuPf8nj77xlTYE5qCPbMy6aUSXX0TkbzW
P57S757kusWxs/vFHGKdjLcNkTvikrwbHLvlMRts+PZ1tbtZK68iQeKlm3cWfNAMzQHq7ChiC9s2
exV6RjmxncJEzkAriceGSugYL9PH/IqASXKQILWI9nC/00g7xFt3uzfa0ohsHTprYbLg2/rdJ+kM
Zer9+Y1JaCp5klcjs733XX/MEoHxSkoEY3ej8LgJPJ5h1kTqLAzV/XnxLbmedznwbv9gmS9D7lFH
KmEkicQmxz6SxNFpFZfnbdwN9PgeVATBf/IxPrEbJMbDAQwPNpo1alH2LKFLhaneoMPm6LBOFXDQ
emgwH6Ljv2F5szFrU79mY+EPNCUQNRs+S/YN+Hh69y66SYcJFCTmWNTeqqMbkCOt0dQHimZzkcXY
UJ9bsGe66F+n3hoK3RKUeqi+5nZ8dXc30zmkM0uGb/dkqJMwkHqq9k2KZiY05phcy70yDc1yFWs5
fXN+XNHD9KhR+ejhBWOFbMOOgQke62pwt98P0DqmzaAoI3YAu/EWpyV4zxT2rCWzGw0UPAcC5ctY
Z1kN8TeycHI/ITKrR4iQwbVQKUrSjELMmZOATH9InaNNFznzfowG1oWaeYUfBGbhJxrQh2S+ZE4+
Ff5kkmYOBXtI7Z7zTI6akkQcF66zCZeLavvXW2ky3pcfuFxCUWOvMDZDigrvqfeccUeOJ0lMMfo9
AoVsrsZak5LyWuRVXCEmhJwsq1VPdb7r19dtUvLmZh1GAWB+4FoBPmjp/k7D89oSySialOiphLTG
ITxDr6+/wTkhW+4ZG0BgMEqnv7ZaYx9bBtoyjYOegrkCMk7Gfa8Dyy2o78Wq9uDy2MpgQXk5418r
RMDePTh9q+UG7pbQT7ZWGD6ASM1ex1vA3Bj9Fx8N7VHBvxcsZUKeOnOgZeCQHZPFnILQ+7xyFFAi
4wzLQWclY20nUh5+b3X7x1RPIAf5Y/hg438qek+HdZIOUs+/KaT0kRQPY4IvFnYBI+aiYik/VmFt
CTIY8BqP1ixT8yklrhmG0Vme1aSffh2+WxLxHen/wirG5H0nIIFSeEYMAguG5OQyZo/RTMNBL3f3
ggU9RhYLyYELZ2evS1zm/rTMVX8AwrFdDPRwX1+6pk3nm7mii2fUVWV4A6YfYWpUbhWCehV5ZemB
/KHHeryL6l/MC2cjz6IwUWt/6M3YcXxmgl+eHhDTfa4w4x3lN78487LnaPCJCJ41IBxGpK6Jgq/J
3IW9UpLKAvy2rrfqYcnSYoS9vjlYfs04uRP52btDnVpRWUJ7lwiTU+cNS82jUUEccCs5M+yjcgMF
4qWvt+hvYfcjK97brhcePp4d8U3xBsiMl3Qxh9xy+1byI2TPB7rw78MvoKUpdobkOoLEFNNsId5u
2a/zd4R0ZnEqXrST3Bxo1bUE4CLjPqHlLBAhQcpYcj3M8bb+WieLcASmhpJuqmYvFdj3mBUxVr66
UqHMEjtPd+FfTdvaFe3X/LS+XFyW8T6C1AfFieJP48uqmRo2GMLTO8PRJeikRiiFBE0iVnWyRmLb
9dHXL6/fVoSmYAOkh0RYMmRGSzOQrrf2jYxaH6aOKYi00AOvTBAYoGzcR+jIdt14dC0tmuxj821q
P4KiEZUAcyTb6LUjAdpBNroecZMlPv7CS7YUcyHWSlz78TiNC8D7y+Pt+CLaL0LVCYQ2jvIgLpFv
IsWqPCm9qdelnpiMAPneaCqdNC1k9dq3XQNwZ+hP39S0wJxIMcID/oN7bSMRCNt7H0J/ObzO6dqs
GZZ2+/PMsteYPmB9PTN6ZOxCuR652asZcSTeCZFlmKlSAtTA/572k9TxPzCJDkk+m1Pk6OHDHzYm
nifhZQEX6EbrxwivKXefNu6h7Zq4XmRcOjkws0WUpaCstTn/coLBGyfKjkB9oTZXoHqmq6YhBEyB
BndcxvqLXVkmbyhPV0VPwsj8TQE0QWVPyyQ8MORyqZFbJ1Gk6NLbBMAzvdwHU4YdShifitGuIdG6
SJVGn5DfaQ+hphOWELVt93OlLnkpS4wczejiDMUFFR8gmCTcHyeDIWyeEqI3wAOfRHfDnME0Hfhz
k037hPL6cBUPnc3YJulrLkg8K0JevXGYgofPeC8K+sq6iaBUFO879h8EJvqu+MdsNbS6u0l4Flda
x+3ug9KQ6xOXiGOfBijoUJDUr0ECKX44UHJJkp4Eb3UiwRjRDAJs2UKsxmSoeuJ7WoZxoKGMAuPg
NThmxyryYAAsUN292vEwXLLMgEqEww3o0NojDgE68NXpStZ3cmj++fAn3zwqi/YCCtIvGlIux7RR
WzF3pNX0aq2tyeVaKKSLjuAI8WWpvVNSSRWs+wAeH96INGA28J/RfK4/sBxhZxkfpHliWtNiiWx4
O1MTK2HfZfMh8Q6WJ5frf0viJVcHQyBDq9BJFo2Qb+HjX4zq9uejhqxqp5u1KrinOVyMJR5Ux+cj
B+R72I5TMAph4elRvcG7+QkvxPaCH161/ySh1kP/95Y9OS5GnXGi2ofwf3KGvO+LxbbnrAK7blJp
ksn/AfgmykOIvyt6DUYLVQlGU78VNgZz5JmUw+q4mu+VrIjnTCsaVkC12Jt7o0hZ51QfADcKywYD
bwSlW9pTM9074fwKuQaN13Wm/c8LkBEyas3HRzuU1w7i86iv7tj1edwKe/38OaWZLQitqcjELze1
6kHj0hfklxaW2fhdI+cXQ4eBoqzgWcfDr5JdIOFHDzDLiziCjY2WiU/xh52DU4AHWV8KdmFXJc/4
IsOH/8SKSN6MyafG+V/1N0gyTEUMqsm9Xp+v6LumU/INMJkh5qKMP2XcKYt48jymhYI6E/FHK5V+
uIN+AXeRER8UI2G/W4K+/9F3SxGIC/BE4JNHt0ORVJBt+BcJZjgVtTzk/UEFRpF6I4a5unwjedqj
NFbWMhupijTZuAzabaCgdkYfEv6Zy6cysR7vc5xQcYZrS7fmdvl7YL1gjn/PSBcuh6VWClX/ziPh
PabVc3XEpuCQq7v+GUsimxf57TK3d7+dicIMEtWRG9gR+0YPJIlXowZs2t1OV7psZ6C8j5kbO+gx
WolYFqMjOWEYZu+wqlu2IykUJNpoOEhV7ccjgRDjgwJoYT/W8kg8WFxnnxfNqL0sYWRFmc7WqyJH
IwT6TUj10OOUc1D/gRVL/pJHW79s7u5TAGQo/VSDM2vh3wXyAf9pzws6lJvREn1OzPRYhk/AWxd6
PVd6aScvJMiIRQnCXvDGXTDMohhCFo3QAhhgGpqiz7dY5N97pvcu5AXFIdsMtAguKw+2pUV96wqa
lvxiM+KVwgHle+A48mjb6V6YLEqMflK0lthmMm6Lt9vdt+UMsCsFpRs7gPjQG189Tlr71XSnZdJV
UKr6vXn24GeEeeqb27JkJU/8o4XIVbSaYK0mkKpfJCMOI89OgcKOIB2GUxLFNKR+509iJ5Ne+VCT
FM/4wyzL2za6gYPOPK4FG9H7kjEhuNElHO3zXIj9vwvtaxbF9UGgYp78NA2/KGb1h5dhxCxbm5Mz
yeCrHRwhcK5VAuwWmL6exlk7ldb0rj1/53iajmjDWAMdv6RCIpYvGNo8HBTWOJfq0LODbWX/FyfW
AibYl3ErB+77yfqUnWBPFg4MlAWTrIuYKwrobn+49QAzB6YrpwNPXKaHgxsmwUy/YIIMqHMPyxWC
dW+MzLb/dnru12edjVgFTvegfkwjum7UPcU6bH2DIZbUslaLOqUm7FqWGZ85Ze4/IYMVvjGo0SCc
J73ps3rgqxkzmZzcZ7Xswdp8FXYv2dt5KE3K0cTBxSsIYwHuN7B+4tpKsDdNo+FYEp43Fn8kbzJB
+C2Hd6V9vg1z0/h839t6OiYq+J0DiQlyO4VGTm3NOtAu2I2A8EOHztNwk/wsr2Wuu39Aiq4a8D6Z
CjDjLCe+/4OMRVucYNbMgIcygLEYOpVD7we2wpol5sb4li8n5es1Xleahk4A9h2ldarKDc7ETtbJ
04cBc2NpKMTO63sJajrhWS9qmveJrgIiOXRvPXPvIaQJKcggsdMq7FM6AmqnAY9UWuqL7KWY8hMO
OeZTR2pV7J4wpNv459auiqDHVpXLKOWMMVOvKRKwprD76sZkd2Qj9+eFZfw4twjj9/ESNbyd0oRU
sEvul0IbkhwOnpyY0Y+fSyK7c8c6fZdaiWaRly3UdrLFXJDfLhGvZ/AA3gm/0KDmfAAGB9ximeSM
bC2iZSXChD8YruSmJo5wEm96OldFDHXCyPLhoWf/jFt4rgZafXcdfm1qORAMZn9dOrv2KqHp6lh7
zxI91tWo9TU/VvegerojVrVXy+XRn3cYE4yvbZVxAOX21LAqgw5y6bUNp+N/ugejwd5K3bwwDvvd
ySL2tI/dRS3PvRN1fXdwYIdTsqoOy+ENElwVknWagzjnv17oMTLeNZMGu2UNuLGlT/gRzRbHzUBA
zjJKLfVp3Nt8tcnDTanMH/S8Dta9PRFzBi+SvivLi6J8erwrozvhXXhP7bKGIJKUsSVqIIrxhD+H
+vMntkKw/Ak9JbmOFYBp5VLVHHKxJRhjmYtq6mXsUyRBPcF5K8PKirV6IXPBqneYrZGlpUE/tBTb
wleM4piviwTvX+FvTJVYlV5Li/zxPxQDEtktooFa5CobYkx/6Ciz1Yjww41WolFCf3CuzZ77jqss
sFLYPOxLNJyxeLs+/SmGQeYirjoV27E9141SprSbdgCEX5iQjL7SXAb357ORtEXrUbRbqrc75GD5
LHT9KV+fgJOh5c6i6H7msbArAKWe01GUjzClyTiVhr9RAdU4PxLCX7I0O23oRG5Kqos9ylQZ+/EC
vQuHGsTnK/Jd6/+HRVCeQqfPlRJNmqKgE05+aqKIwPXUizSOJEUyxI9Qlqgfe/6CTOzM3CbybuAi
8w7wfnK2nSa3Hw48FSzLj1ahCHnHmX5DA4Ac9Kes4cYNYRCRVRnIRLFWoU0hfqBJaIj1Pfo2pIi7
GzHn13BGd9A1N3awOGFUAmnSiLlI+2Pm9Wb4lwxU0qZ4V8yQ2sZ/PV3HMM83/qhBS+B2GRJT5JOd
7S7MkvcWECREkC7SC0Q2GnUySk4L7pXU4MqJpufjHI2HHgDgoMteXba3yIgTvdnlwmdlyE7873BD
6iU/AT4nAJG7qsq2fWYgo/8l6uwb3vu7nyKckTffyzSuUYfpsRVWo8EASF49BTmh+wdCCWM2r+Le
OzjLeyVJRnSEqMNsnMQ2l8Rg8jAtmYP5UCkQIkx5vJ+gTAnhNDv6C9O49DIfSRkOHLkGPPZgLCk+
FL8Kg4D5gfrJN5X4EpZqqR+iJ/q+BjTER7lXg2ecn+kvZ4WCFkv/UE3zbau+xk/srA6S3x1O9okL
gMFzTrDZgd5v/c0rxUR+sGFNYx8pSD3+O5ILfshjYPlXV4vCNlkZ11VVUTixR3IUwUM1IPMK7zkv
ejH5D0NyQZ0AA+uRj43wEBcMKI0JoFH9KekmmLBqoKKXz+GOme7JbGiy3F3GiPoK/d8VHFpZ7c84
HKHQ/1F79pSajmseFT1ESHNN/bCAVlcD/6b92a7T6FUOYZynnuwVwROIy5ZruMQFk6gDgtnnTVF3
5BmS9S2zFWNvWEDG0iXCYqbulJoImZPhH1nAjbQ8rf1BUZx7FeVKSHs6HCIi/3cmilmi+HlsnzOr
XxkbjlgtuHC4X5LVj8lypnhwM9OuqGQZDdRp2smi9tPe6N3Ux1vPRPWyg2+aqXXVE/gadXNv2Fgi
4ZIm9IYQfmYo1pkVnWXQwF69qWrXAGulXk7BHarNN3pdfSAlQfj1EDimhvw++30hM9ICJSlTlN3o
Y8UsJbzxcdAio4Pfc7pyWSycax/rlQK/skdar8B4/6PaBsj2kkn0qKLFDfSj7WfHTigRc+AjSB6B
aonAfbR3AZV5/UEXttuDj68rAcskw4QM8WIWJIEEoT6y+xL9RTAZrB6Nk+uMv2W/Xp0cGvx2qb6p
ZKPy4R11F4wpmsQXJ5a+9YNbPp02K8WJNGOGV/3X2V0GJkx3j4leVixsJlPNL+fEQgMZtf02pS10
Wb3091ohORhH48/G43k036ypMfJ0Jqu/bJ4t425RTkTrfFUPn+CpkjkHQCr/wSWatPjpG+gu9r4A
IXk1svd6v0szu25vqKVS+infykaO6/4iTcCzx54Wz9sF+J3WPupy+3mg18mqtp2alC6Ms8Vl3EO8
yVBNh5II4yc/BPYrq9ao3H9xPOikO6jIqUR69/w3B63GcBkXVpHMxWDulriyU2LMe4w8saKAJp6l
bZhShEWaidfibm3w/bOPFFFZwov8InS6Oitj4d/sCKYaBcA+K7PS23XW5Frkm7FX32Y9uGUB8gPk
gtqW9VlAScfGKHMfpDP5ByDLU5feDk+0+ZLwnOeI4hgA058ZXX9paFJxyTU7SJzqnfpb+eRdToYC
lr0ax0dTiq6DyWp0VJ8cHdtucq2iIZ08o0s3nVd0ABDO5atBDfrxUK+mwZpKn+V0ysiFqQ3FDcGR
AjXZwn3hDoU8icwRaWVS3B3f4p1XEpFLqXEUK7vGC1lj5oivb+tRfvGbikG7xHqoH6tFXdvCh6li
O0t8XRKl5BJOlYmjrnMyYi7qgy+feHdAYeGD0mTpuVgykTgpUA/VWGtSle+Y6ORKgx8Jgk1dDd0O
es+3RPi5h5cAu4dlmlVhVanQ/yXDv5/R2yjGimebHEMAWweiwRVHk20b7BHI22yB8SM68wjY5BsI
pNbK/yU3ZfVh3uyY8ZetMMF9udOOq+BuPIJdD74lvce3yqylF5HpqhynNDO/Z+pjcYNJK40E5lvk
HztECUlpu2JYF3G8nl9JQH7hAloWXTYwfZlEspvOzgqfWf1ACLcGgxtLbI9p/eyuEkEraznfqlGO
c3W1nfuWxshWZDWHExTT2aIqYUfojpDejE7EaBA1g79LqIS5J3rkL39ERmUoBhmbYTRtblEK3UyV
gXQTMt66oX+mjhyIFfZ2uKwhoDTHSAs17llZEOUfxKRBybvw4K4PZTQM4xSOK/rrFQj3RLZM1z93
I7Wjpm5qblL8xKAVcTby0wft65tFdKPW+5EZgIfGy9o3T/k5UZocSNUc4lembFksY5I1av5S5wlW
bc5e+hez7YGWqeBW6AH/qRo5XTBcsEcoR4hxpLcXFM2BWql0iQnK+Ho92XWtd0HF+OKudopFbBmc
FfGyne4Mk3k+XkQDDrIXTqI5zr1EAULzW59u4yPG3KGsV+HBK0gFLal68QBOW8TP2hiBOPDq3+S1
GSpb9P32hqVjvGqTUCugfi0QFRNwGmfMijKDpl2Nj96zuZeHRzQbO3RKTqTTNanOZNJ7D2n0S5Z6
ZnXuL3K8WKcSnmLYftRhXV30FHLCFaHg1k7dR1euxioA2Kskl/2IA5GLL3hXXnmejtqQLZvZWe3/
S/UKC801kwIu47MS9jMWOzSoSaFgsULWa4meBhr+6zRZ6nmT7pphVSG1OkSuOyKNruwDuYaccjY5
wZ3U+QczCC6Vvo/Oyj3Gs1JnzqRBX/nb1f6oUzZcgQAQafWbrJRBiidwFh9oe6rxQ11edWC1VNiW
0qxbuwlRKZftkaxCuaX64+4NHTMf37di9vr2AXm5uziQTjlRz2NhyIFeCe4SzyZwspU+Ck6Nwgic
hVja5bMFPtTNBv6PqYZEd+xZKWgR+KbgCM/Wb+Bzecx0MkV45QcHrpYp1xEVYwjShrbW0oWgdJ0K
gCbKFSKej6AFDdALJ2D+V4JD4NBf6mtWKTni0VpPVKcAGacQmUDQyw7Nxhx6T39mC5YhDxViGASE
ghorBk8Q2YApcD/uBgdwsA1bUxZ+YmMAHJ2HZF/H351vsNF9udGmiznwEIJl2s8q6aulGIMnjgQb
410ArjuauS4fUNNJL0epx3yluksd3tapqmVpTkNvYAa5nrsVeH89P06g/YM2YmmwSEdKfbdGKxCm
QUqp/iL86gvGA5NEjf/UAnljS1b0IwanwcFiI4/roAadAVPrXqqC7RJEbmA0STyTDGvwTf82PllL
4D522wBvuAFP2mQN+8/aumQXyiehwqQfbuzp/xZ6URLMAoHREdGoebmSu5E8mAGUpRrWKuCIVTqM
v9VPoUk3Pp1BcAqZ9c89A4IqLzWxF16CtCMuQFrFvfFKOVkg9MLl6LyNYOKm7Flcwqk/HMLAU4YF
TlAfv7V/uNDItg0CJBIrqINhkXzB2nwtiETFDb1/e3vXD6tN/S23PE+jHc2YG22sE0AZv3ee8gwp
cT/qlP+Di0o5ikCl966mcBCN9yH1f2JlURQTPFr9ujBZvCkBJ0c0DUYSmNpv3iedRbcaIQwLL/KN
Fo8uU+dHqTjKrpM7oexX30L0hXseV/lkquO47NQ2QP1F7/9eQ+O0utS2AhxMNHSqN3PidhR1eofh
B9rHrgt+VW9LtGjuuYBI20k1hhzznDbyCTNzDkpd6Fnqdc5RHFXEisHgf6VAtm3YDLlP5UwJT/ir
poxyXvnEnV2MPjIsz1ym7B9SeGnvtmnW7jfaUY6oQeH17mHd66klSs063qpfF74dqMx8sQAiQGaH
KMxR4SzxWNLN/eMQUjSMkRWMKpoHUEDskZewFIS96poj6xT8v1RBByXtGndzy/JNh1/l6ZwGPnp7
QCsOBwFiFVjWjoQInK/06UAgpdvaxu51ZQq5fwKc+6T/636BwPy0y5A+H0olrvmY7YI50n3ckyOh
JwrbMnoMvcpM3Dizz6kQktAI/NKpBtLjqcUvADx2WC5/S8pNKHH82WCZYaOokGPC/6tQmOJwAkcL
/BeVPidp+exLXfLuAUYsXsl9VoKGOgD2p/31B/v6MwZG94WFhHNWouw0/kC0RsZfugQO42VKIvZm
nCPuCLoxPJ98qxztvvobmGPYo9AlOdaeAxqH6pvxX0F9Zoq2DqWOa6vyiGfj3JqaD7qPFZzP7d6a
whA/VWsTCkZQ5VYmZeO76RfEIR9Hvrb3l1zS3/BPuM/MVzFiI/JvTpE3n1m62N+rm2Nqj08qV8jH
oBhXPcxi+eIroOqvtuJG+lU5c3w6RJN1REn0xjD81P38CLGEV1Ssb+jPs+pwhmt4X62hnOSTBrnL
E8olJRHdzcREv+wPGuoLR4Fi7REX7o6QVJMnlWUWqJLEwgMQ1mzhotSYQC8E4TIP2AnTL89stTwC
aCMLbovn1sWCj9VpcI9jm6UhGaRVQ+O5QvSsCkudHGkw39tlHaJ6LJSmSOsl6EklaXDwXf1cxqZM
LQft5VIb1c3hUpK+wP7WRJsxYSNOxbfZ7BnxINRsdohyMXM96nlVty315Bdc7kvct6Nbvv5GrdwW
UIPqaVlTwaGcr+LLNSIgFxPolnaZMGcyNaC+iXmoG9KhZE1hN3jMSZ829XmFBN4ZjtpmPhQQvAy8
Jp8+VKCkEtoV3TOc67kGa+pYW9pIwsjRuzdT437Ifm6WwuOjO2XVDB+QWBPugAIW8I1j4EqjAJLc
U7aloniEz0ZafBFrYlfaAZ9TG1vNuiTAq0mr0CtwsonLAHl3O4WVuVj6iOowfOGWKYWmidm8b2qY
J0PlqRxZstwHmKmhleX7nu2+RDHG8mEULcpek8HIvPIm718eXkNMVnwmyNOFQjypowMjAaPqJMHa
a1tAFXfJVcS2JtV3+4kVQY18ulUA1ZOaznp2SNOtiubCuzfIU6seRiegcCIFQWAhM9zBR0gmEaCy
1sdk94FFptaOEBWHL4dw6dCgAjgUw/+4tZrPUvug+ks0fAsTqSfroT8yhrbT1LSyqMwtcqj10zhY
UazuVs9el75u5nHIn/0GHQcXPuZAfwu7uYEtOPK8ZBoSZh6MP73hW5W92RKtURnEArDHfdPOWjji
FwuppDVvEJQmr5ae19bT3DbmSeHWELjLCCLPuKN0rUIJ/Hia4760QaSRQdPmSMDZgCC1vI+kvEAq
hqEET6XNibJQXRQW2NAXknL0jAUyZeaBYJ0B2wLRrwkPgBcR9Qv1tdh60vRn9gxie7EPCAfGpEl2
ZTqJJRq8Te0F2N3+EsCCTGTFyVjnv35DlmKdZ/MRj3WM/vNr/j/DV3ddLZ3SOi3nlMnw5E832Gmo
5YMwPBgw1DWEMdE3RhTtQvz+kK20ZsCK13m3rZ3+EDEbTUbhhc9fdXaOguD5KVT1YqLRfYd+49nA
4ve6aYFhds3DYzoz7fQb+xHgPzy9q1Eoti9jNQ0rPkb6oHyaIWNlGIicfLEXm427cjByzuA0ws4U
AXd40u7FE05OqPbSiNYkUl9Q+mj2BCPg9NqOAvCa40GRUL7kCKYcZFDVtSNfcjebiTwnEg5178ht
mXPBQC9jVLOPQepvxYrfG1yhwpg1/5EbKSVs+7O/xy22SaQRxpNZrh9nZwD9RwHmT7Lz0WoLsAJX
Y4gzn/YHrjiWXDOMjGWImlGxnvb09FGetN3nyzAnJu9F1kma4yXWA8yz7QdGIA60pl2zRDvdDXLY
Lj8j360og3+UOTSom7XaVFBOF28cYISoLkjKN5bL6atMNjhzSBFnSXcylMstxek9dfWeFW92+LVn
itpBid5eCN2WXCp/InQSWpoRy3NyOL+3PZDSk78YsITqEG/4wDb6ee4l8QEHHT09N10h9892WMJ8
ZNI40jnYzgLoVyScloFgG7YyCAGcVP2LbOWTcnxwlR7sdzXmC/pz5fQc59sJ5V6eHjcLpAdJSfMK
xu+kRoT9zDgAWGrjjar6bm89ldCh2IvOfVbIWrRjLv/Zbx/5fTGt2CtpVexayyeosX3Ta7TnrArU
aIvAMc0cwouEoF/L4tSgLyWFmvygQoZNALROpRuMdrX9gs6ln6eplnLF7Of5B6JLqhNjN8ng/t1i
3aUDEr5qOObwyxUBG4iRJ/Cq+94gQop9kuEeQK7pfEGRpZUbXOwbPX4+VejCicuOX0lK4CsWvj+J
gjAhhsKWknP/1iBiuD3nwVzuqAjXnIYQbUPwKX264J/eHIVmNYNuw7qCxTQqfCrPgJCoL2l4fK1M
T/Cvn886gFa9wAd/IDlIzY+D2bR1tHsuCCYz9m8SuHO12U2a7EWmRozLyO5TPrMjMxwKawxig8kG
j64JmQC96Zxu6gYmZeOHvGokeG/RqzNLFPcFyNtODqNt5tGftAjK0+iKud192JBDk/Y7eGlV52Mf
T1TUq6NCVEIaXuyEMcSyLId+6hEwp1H+0dL4siiY0XB9oLKkhQLwkTF7FyttYFOVb7KLCwgfLlE5
+bAgQsbJhW6euJpkxBQ+drDL7FHkRVqbyARA8m/LInw+fYX45A2ter9xImKjyPbB2LSpX1wg9jCM
ebB14PYuFvnLOh42zuAVZedIJKi9TtK6Ya07C8VE9nsIBe7+LnCDgC90oQdkLcSstvwkRYqc+OTP
IDKMAMncYbqjvKQHjbTtq5JmZj1/6TVCfZK0gWsSfXwIAH/1Cjj614BG8WJ6NbCwOZuwlCL1pt+8
s/0UAxRyPsmkS7Y+PclH1KqBpye2kB+fTP327zcjzJ0OdteRBgRo+BdsNrteiYM982t+HagPVrFR
TGnVrs6yOJIEMtKsVdZ+LoOg24Qy9fKmwkCKmkANocK/sNDhR557guBwCEokSJcNpSufhk9ddyZX
Gk9+KET7VRwBP4fq930uYo69v7xObtvyOMh2nBsaj9t0KS5Xvp1uOXSeuWcM7d10IIegNLaTl2bt
oBCnvRyMR2SQBuBzBlnuBv2lXf79FWaV2TXw5vJ3YxL8/TNhR5ZDrpC2y12is5GGwUQ0nYrwiZYF
NIZbNxb1qaOniu41nOAjgtDA7yvnGmspwlOc4Te9SbnIY4GFd3PFV/Hu2nydRUkJnLllODzATbQz
XV9E2L5tgld3mAmyzVSeZBt+LIaXvrButxX0uRHCx7jclSm/hwtsqviEtPwnXcgQbT8ADtSvhrCQ
p6HK+L5DQz/jNHR5tTUgawEpN/9IAYPQHZ/3av2JfhukLh6VVcIqwH7ji58NKyBoLP5VW2Iee2Ar
ZK0Lrl1Ji9n1lAa+YQO+n22oeMFgmRKkYNomBLtCPyPESDE6cTvZuv59eBxYZUexOp2eEryOCven
WvZZ4ltwW5J68yVMowGKTOsgcIvpnmwjWImQ5rmfuVZFqWMixRVV/W7MzpakED0GbTd7z4XP3qCY
Uyc3w4APuke3YJO5nDvYQ+V/JnY/qCGlRHZ89VGsQwVmzCY+ArXgsmDqopEBH/qkXaS6V4BaANgZ
SpGzHAo0b76tX8UK19NZD8wHt+b3hYQhtSX+O17ebCU99CfzqS0A/N08b9Xd6UsVv6PSY4iyvURi
w1p4cBtXz1RUVJYVy4iR5Mo/5nExaek8xEr3XzzuoEBaU1nvigYXVQBpLi4b10mUe6yA/iytorZe
XnwcbXQRU0z3qtoC5P1It+dYJ/osVeRFYFN7nC9/POgcuZPYT7Jq0gDyoL/rTv/Y3tNtEONDh0dE
zmQ5KcHSFFJD2qDOm+zcLlXGIeDBPGlcZOUs8X/xY/an0Szwl7iBtmykGCf7q4Or2QrM8zl9LL9r
EnFwLZDQredvV7UGgpc7kYxso60jALlB8Ard1MIKnclP1NHDkGIhqZVJSHqo9YLUz/pCAY2NeGxs
/Gw/WhjkO5H/BFXEfvJ9mWCCrbYaeFi7NxhlLLjfCtuhqEEsQjIyxtvZ2ZendrycwMwxDIr5Tvb8
K02khwv7Wj7dXHr/sd9V+SxE87qy1JdUYC4tvJ44Vnxy3neEt88tRKBYNH63Emr//jC1O4FGf2MJ
cJuRRWeB+c2s+xmI6EtJglV1JGOkHouWS8tg8hKQk2kZoe++sOZJ2XO00ZfNnayIkzPJaN/UwywP
nfWKfuNGd21HotPDYQGWwpw12fqBLaznRdj8ALQOHPPQfkHl2c4xeJ1RJhhExpn594E3lbPT8xvr
/8R0WGYYVoPOtk39AtmhmRCieoimy3GdThceyGsVQDqFgSN3QrNzl5XkOK68j2Y1njJragupmnGJ
lgff+kRHFsPKrguA/uczXYrwWeRYDwSBTvI741jHRYXYOHbIw974pjyRpkCLJeheAjdG/BDnMCub
NdblBA6nFmYY7Rn9wu5Rmll2FlMaKdkq0+t+QLVo8aGhYKCUPDFFY+8lzkxaKbfkUVqVFfPr/2hE
utaoGmMkanoKB88XwFmksNSDccPftX5Ib1wF1p7MIbEg61T1eobBglzIDodleO30h0hjC535qVox
qdant1I9L8LoOhIljzaDKV7NKmhjYJofbSW08PtYAHyFXy6rVHFOZeaY1GHTrPTNpJWH5rl1ag11
s9fGXVZAxrpDmrNcQQhKX6n85YM1g83c59qpiBf23gU+xfJJMzYOILLXapRPbtdiqu5YbLtIHVtJ
dt5jxzSLfb+5+yWnndb1UAp81mUc28DX/Cltg4PCOsiP6b03K99wbXJ1W/filTy684I1iXPQUIE/
2OorIGiefHicQgXWXBMcsFYgGicLm/9KZIKDDAMK61MqjHCUVyoeElFlSuf1eNEn3pqmBDk2aMaH
GhHq43V3RSNsQI1lDAyIHknoiqf5nw5piwmf5TT3JlpqrCXs+U2wHptE0SrCbfrrMY3aNVzq/LvM
UE/Sfh6HuFbOhImvjcRz5TylgrnF2HFZPEYUsmRu75MF4hYoEDt1IWeRN9ZI9YWI97NsWA8LXJCO
FoHZTlvRYZqsCj1sSw3720bm7d6gpcOx3JHrqa8TRcIgpn2Fqx9oOuSkuIKOHzPV/TUUX944cOU9
y4KhYRVOw1Tl5pdOJpSeWr2PsQl2GGdeywkFJ9l0CUQ5Uul9xGumXG1OhRs39bKIOxdhUI5sT0j6
8zgSXKBbDp1Rdh3/xHcrsc7drnTI+RdGbMzgfLTrSfXDqXYIG5H8fR1U3+HOBmbkhM/zOXVBQcTi
Atkk/LwK3irW7DOuChFQsB5Mpggu3S0ueGrdXDHbyxGRtCNX3uplSS45B//PJgm81xQFTlJv8mZz
12p+AbOTZrHy+TPPcReQ/wn6OvlriIIcABEodlOKF72Sw39Ox5IISpFOQRc82Cayf87V3do6HnGe
1o9RSDeMEzRPggHfuBJFV+vEJrBIM8hIm/rSF+iGB3AH6mgtQNrRPySHTilrsjWJ6SS9sm2tuoU9
DjeYIEUE/r3ENTLiprpM9kjjhRS3XEly5s4YXeWGRZRpXOApc+CARmj/wEy6E46SNkMDOu0821lX
/naiFHts3PemvAuGCKdoyw3DXe4H/cNjMxJYB/iF+XltNomAZiSEkekTBxo8Mhq9AovSM93hD3Ve
ksBjGDeXT6hOEtSyASAh1YFPxQMHBjXrJQ5d7F0siXkO+BlIPza1sk9IaTGG+xAx7xi/c23yh00G
wP9938DNIuLBTQcl0dUN8EoUmcGlI9Gn+Gsga/5ZbBtK2pE75H8mQyMWoSr2B/d/LoPcDBMO9dzL
5vJdDlOOE3gse5/2u9WDHLFMagBhJwMvSolGbx0o6pp24VXhUXKI+qlmcVUPKsZY9djClyHrZlpa
jIVwjP7RN+CIyoeHZT1vdxlhvgP41s5MNYT86aq3TR/UeuGbOGxa1Iw0KMSPRSQtkItjF42+fDL5
iV+cayYEkeXmihgUORYu0V2MMbuCbE+J4fMUuhX+9jwI/43zXPW2EOO+XW056H3NFJU5LYF3w8Jn
WPjmzpRbDLqO3OVJcSo4Nv3OV66BrZXoGgponLlHvuI6gFis/QTIjL4oGDCbBDwSae7jzYd9R/Yg
fL34ijuLOtbtI1sHGSKc3x8YqnqZci0pdaIjCQ1ZBezxpdvHJ3GrNdiPz1F8+JWxKQ/lXs2J/YoN
XqXq4vk07FQ9YTzoHOjYsSgJrnQDLbq/Aaz5cyWlHcLEKLLNmGlugidTyf+F50A0yfXNkVp3mgjk
CD7CPKm1f8+vxjBcmAIv6LyNnC6+7R9xh0DoD79wHxhaOrnLSzlzoFRnp/c5gJoZ74x69bp1E0FK
nWjnIEconFkRewsZcTuCJJFjhfLs811rLNC+1+c2Wd0IRIpPhzY329OZnzoShrd621DNDlJSaYwA
CaDb9LsN7VNjlB9BcOCjn2C+mvhNNI63FyMQbtGYytG4w6KCLuB8BnwN2gPeoVjhMtw/bcBwwe3N
5jwToRge2ODJiG6AViMoU9wlD2Je8Sjdo/UWt63LP+jzwN2U7BFsuIHnlEVzku9GQSdxfF4nIHB3
GSa+RN/XA71cTk+wV2bdUyDN9bjS7B+fNItyyQo6jl41EJQgXDRMsuNVhbwK0yXcHiTRkHOoRLRS
bHvQHI1UGRH22fHApc8NmYURganQEmgfPZ6is2EHTL2wNh7G7YI8AzLtaSl5Po/hbJl2Z4DReYFC
7ZwNRGg8xMaD179XcO+v4zE8PEOxQUYsHH3X2YtSeO3ED/g2APQqj3DprbdFEUYu90eqc7HsjiFy
5MwLBjtWACdw85zUSdqlT6qbgbfOBEpH71caV29VrfKU43z3FxzrsD0lQ7fVZBON/kUPEUm85I3J
tK8qtt36FWMgX7D4juEMNGZzWlroZ7SSFzix8EWmEnnr8nMA/1a4mo9l3EP9GOAZWm0EIBfllsKX
MO0A78TBZQvUMz8phV1Zzv19z8YHKOKDe+Phc7AQIiyWfQ6E3l6Rm2+amVeSwkSw3rsm8AAczTIe
2tpHxYDpYhp/sNlrmVQFgBEZESPgQqainnAZmnojojWNsDQ2/+STAKorCDkhDVK3Bc/ERuG31S1b
SeYZGal0aNnXUUKvd8Cjmm4wGV4OBszziXoT635nwHu+KfkUNArFeHoQLc0KVANb6wHYEmDYoKuN
51xtKvZY7rERjQFWGoqfF4GEs6ykxUraeOShgPQaoosmtAvsmm3WA7IncVuFCsz0wty3wu84Hxei
RahLCGDUltKZG2T/StbMZYe5kqpuLf9qRanFPxVLnU4WlMVU2RZ48pGwb/aX7jmiX5GmmJ1cQbv1
/h5FO0WLXBpaufAt3C9rNCbUmrWZyuY1BJmeD0y3vuJ0Idg2Um2O3TdlhgokW0Ho2PzPRF3IEuCp
/JorRJzhDvDZHp1lk0lma2Ta3/JHHEOL7kTizngEAtbNYK/6xT0mixda5Nnx+sEJVHkLaO7n0y6b
tcAEb33z3MhKHdawRn88Xs9pHjzZJ39OWq99eCorvvI2A+pIK+U+dZZ5/xaoGiHZ6p7tlqUf1EcD
TIX2ZVRtc65zAbDhdR40T23985OuWuaM9Z/ggbA1yAPs7Kx9MD6sDkpr46wnkuQVeZjG9nVcaEvc
A7dvu3Bc/a849589PDbyu9T5TXIO8jGeng1VjU70e3o0XOoZATIjaz+jwJJGfXQTOCwbVJN7JrHE
i97WduZgPMSCR3aGT884nZoYmQWnZbkfS25mQklgX3SG0VksYzGJoNiepuM2WNBnPSgjwbrXOv1r
hbYh7en/ut/iK2n+q/sOKX+2xxbd8HsytZV0mpzHRZuNgLNaDaMVB5xFt63e2K2ynvXUQYoV+lkz
W5n5aHBYTJvQfhhnQFaR456CeS7nssSMCzK6QqVPKbPAWtaHOvHj6hd9c8CcXYg+AughqigDekzc
jxnLYCM4TWr1Mva2xn6dTtsqEhqrdnJRxqhfN1BSDxb4ZT3D8lyXuImQPwI0MhD+5Zoq6PQnWFUi
CsnPLR/4zsDOPxlCyZTV4HUNobk4yT5xljo1v4hZh/Omvie3sNDXv42Jj889gvXgLAerFocwiKak
dR/j7MRNx93uSutAUSY30bYyldzlpLvbqWsYIdPhNWSxcOSaWXzpKtA8DqgatweN8ZNVmLr/J1+i
Z/0U/ASLSZOXDRVMCZpf90CqzaWqOfJ8NkZ3onD/NRPCyj0NQjSMsR5L6I77W6HlUlaSwU3bh4qX
yPi/UH05f6FC3y3/WPky52vtLaVFHapbSOWTltSdZno2Bx3eWH5Y37wQMWxg+63egieyTgFbZdk2
X5/A+6eYLnvINLh9o4mqVO/Iho1gM08uY083XtY3ppQc/YvHYzbOTHvlwy8okxOO9QZ7wR4KbNrn
axW0JrKTGkPL0oXbAHZZ88cRraWvAc5vDTY1EOgMF2IltvajSUgzMiYDyuZHW01qPuoaNHEfs3GD
JxSQh1PaIva4D+8PUVcRPYp7riUiIdPdDGOIHyioh1S7rI/mSz1oMoDREqc3kKVm+/UjFQKKpYCv
UOHU7VQnYR3P9DKAQD2NWoopwza/VtK33cE6Yn2T20ZSjPScGvAKW3vNCd6gAITmhvZ0Y1u4EmQm
xk+DjeKLyuA06qhfuESJEADb0QDt2d2Kq5qvQCwcjCopGq32bkMRcLDTC/sJgisK0L+us0J2kbfD
PN9PDjRs8MFACRqQjQNZs4OaXQWV7kt1M8xzl0eHpS7GIliTKAjXk/f9ltzFBLNuICk2/put2hpq
cZb92k5IrgM+5dBMq4rhFwb5e1VY0BXfG6V49gxsAtjim12TYoqDMH/6/LJPg6x7wjX6he7vLh1M
+sN69N00/nmQjdfVj7va2ffesGnDiucmq5JiMK7v6DLr6wpO9X0fqUHSsdTl7ApT5ViyTTpC7Ke8
/Uk+3sVRIThAzP7cZ0G1glcqa0842mwGJ+6hZ+nX2SCTc8nU40X4idqqeSVnRo2AiiVCbDEk2x2Q
ooXPFsMb07+jMCM0LRlOu1AGCjflqqy+tSk7+2mVww9d6IplOrK7VPikilVSEXP5CW+VEHRMNfWx
qwHAPtk3yTh9CAhvX1YY3phsCnGO5u0ZtPVUdTdJglKxEDhRLKr9RQeNv/Q8za0QdTlyPtpDdhnS
SS1QzPh9rm+EKYHhSeHgyjcy5qKuVX/j+q0lfFeBc+usdpEiO9I3CPv5PNcKIGqJSIFRiU82qdNX
JyR/8zMI+pZ3D/caBS2aECGjgHy0phfSBTB43jBcfQqrroAIDpd0LB/xsmF24sHBd8q9naZedWXx
GjO0z1d8wZmkJL4xDdDSEBzFFBheGk428mb2tmRM08RNCd0WQ93DgIwuITKWDa45onJuySv8B/nZ
N0ZE4iH7uYAX2Lnb1L5GTJ35dRXTyETUUqCDR4rgWxaNE8CUQeBtg2vNc9lXVMq6zOulfdg6SrpF
qTkEgewX75VyYTKuxHlZexthNAZ8rrsowqYFOP2kCpLO/WilzfaffAX2oywjp8c3QcoOjuYks2Gk
orAdZa0P8TNixS1eh52r2QV0CZsYKCDCx/bbeZiZtuJrQAJh3M1YH/r5kNxDifKYAwF+6XEKPHvd
z16Pdo6AUmdnBWmCL2XhTZp8dIP3RGsE1/pCCV8Ij6vyd5yp9rzNeXO6YGKxT1+WQx8RDonW3a9K
moYYIKAmfpdqYqcfCplO1Jou1CRHOsPHsex8PPhW3X3kaFl9l9smHsvgwcfU08qPrvWVKtGloh5w
KtJcUIfR7rh93ZfWIzAqru7ubJNoMvV9GiU+5uClLCldo2dQ2cT4frpDO54oMDmjStQ/0Iuwn+yh
V1uGGvGXS9woMzhwkn3LkzR+W4DHw9nzUoZixN5edNsLyI70DlY2CLt1z7RBCscpSebwIufaNzuY
NHe0MNlluT6dcfg6Vo755oymPhyjEekSwBRDt0/lsoycSQCqx6cFpeLj74BPkKBHgCVr9fzzcElZ
CKrQYtMZBVfEYplJlTvjnLVKyPvOTo7Rcm2T6+CWk1A+fFhzvIO9QgivXPXqGC73xO+kHLklhhNr
duhmo31/Onz+/68vcCc+nh93UCpGHy50jZOBAoJvoPcObK6ib0so1DVSIz43d82JZWYTwxs7fZlj
wbGRAmKW6nTO9KsqP7SKpMn5fvSglR+G+F7KDHMSImgVO8tbatqo/fzG7f2ImfZx8YZ/Ok+eFXxH
MyuAO9VjroSl7bV4C1Z1ILqt8s1jDF6hZV08Ld7G2rSTh6h8jdiOZG8INVVpWfomTso9+RJLNO9H
1mxgFzH/dzs30AVjr3N55Glie5k/85fop0U+7r2jiqP9NSxbOS99ypzmAYpfjx6GbVkFNszEIHfd
yjKtk8cHitdVVWgvm6iZKVXwIF8jM7o3jFI1xYv1zP4iDKNzcOXNmyApPm6tBxNkOWr5+DHTkNI5
KagY59zyFu2YfNT3oC08RbxCENSmEU3BRQX3SCdyfrQQHtbnr4/0YHb4DEetK7tt75/lZf8E3n50
FF8OQxIIgAOuTaXdoehKEa3i/+gNGkLAmTgI9uPT8vPcqm40a1uDXq0RZzw6+9P3LKeKsm1xAZj4
OsOqGaIBmv7qiO0DDgPScc7SIZ5XjQSsaE32V5H4ZQhLtnQ0Tckae0vhKUU/Xkd2jQUQWU01sj5D
jVJ/wVWFby8V8Nj3FV91bFvyhzGc1Sr+fi8/Q+FjhjbfqlrC2YicfGS/cNbx6yR9bb+RnvdkrF/S
YH0MrCdgg9QOrzzIAC/maDXCoLbY4gKhNEAwnZ14dEd+zhHgdSHpfrgzcvuVqAbv0xBakmLttU+H
7TBogE0Ypy2fWei+sD2I0hFHGk/hs0BLzlKwo2BI3352nsuMZ/iG2VgrB5NjWZwxE3itM8LMutmp
1Ov/6otqNpACQl+AF1DvnJALARE1UwVeKAPCyBts7hwdB+Shs6MVC4LnO0sopBZdu7Opp9djvtbP
EnYvLWCMwB8gvkF8Opts3xwMCrYYRRICj1tXjAACN80ON2YM3g5v84h53P7AfnsBxI0FFvlbA/+O
dC8tV9Y3qhTBkgCG8KiREM6Mi2we3AmclAat/2vyuNX38vAQt+PS/gUOlWaEPfFNLnyA+ykNPZbo
Z7U6mjZZr6YqEleWyqVZQwCC2humMMWKfmNAhqVhnMSi6MymC7FPYWV4nP82xuSFgG+6YzIRUutC
r2J4TpLe8TAGbRwXqHFzc7SvdG6uBXebJ+vJYXe3c/yNJvzmEtxRl8YgRvwuQdgnuKDSmZ1IKx3F
vIE/adBr4XOtSqpvm25+nP2XTv7laOb7buWOS+HvaYNAgkHcXNKSMmzeQi6J3ZpZqS19FMJqIt1a
xxqys2tCNoFyflKWe89iYFJoFueXWf1VrL6NHje0LOQmBR/v4+69pBIRaX4AZ0LBu0uqJr8kyKQR
iErV0SsVy/jQhUuwSMRRsq+PRU9aDTDaA5okfryoCReKlFwH4K+q5EvalT25JLK9+uHkv9rcxBnk
cCK40Z4GbUmHpxavhSCfBkC9rr4xr3qmpvuRD5Ac2fS9gQJ7iYHseHVE2J4oui7rKKUnrS4+NYt6
UXn+qaECqrXNM/R3lcRwVP4HcytG9rIyuZbZ+epjNgCllqEr0fHPVWhLTYnkvAsJYdnCM8ZyMAK9
iRmpqZ2GvZNFHkNBqb44x119Xmj9KvjsgbgS2GwnYK9K3PCbePhjHEIeweEZOP8UsmD832vi/wzr
lhfobMddVXk2uiBAJrEssw6QmXv/VNyiJr05wPgnzUVPYo3fR58RWPX9xaZE5NoXcJUc6JFew8N0
AC83+R85yscayCA23/eHowuGH6khswd05zK2Bbw2HLjGFM51pIPygPdtuvjVWvIG37kzwB7g/O52
qQzDRou/UNU4iOHdLKGtiqvYSO6bSxlcVCsjTFDWgAQY8PN/Sao37AUiQE9M3fCaUEFAj6zCR5HE
cQxk2u6ek9BElA0T2Cx6Z9J/SlgaVbAqchGeZqkLhmVGDqG20IJjRklsuTyJVtGJnwCyCmhIjKxy
a/BN5XHCDpWQPVldbZ774J3h4tmvciMA1LflpiUwU7BFizWojW058n57HxyroKKRPuMYt7ZMjQz0
p2dx6NTu10MFA8bEy0IJCDQqy71KnR7V1cXwhfNiutYQbktnPPipVasv/9fTZClrpQz8Ul8MVC96
2UKcd45wN5q6Rzub8Tvx7feuLVWrctGIfueUGH1pVQDN9ua8e78tvDIccJxD9X5Um3NokBgk75QJ
XFyvGLVfEq5nb8cINSaELkJ1wvw6adZsD042LuiCN5eS3JMHvK8gwLs1Qvt2dHhGKTFjVBH56H5Q
FEqvurys8s++7+yE58jIo+KuAbjmpaQmTtY50C2sVn66kA8MCwySOuCPgSSVLxOMPQIk3+lOifoF
YGh6LxO4JWy5WlztxX7baJHU3VfzPWavk4F4QLo7frYexMmwz2D54Uj2xoS87UqTigdA427HjA2E
nk8LYu9zG4NMj/EheqGQLbWL1OUXuLtTmjry72qw+OETcKJLIdWDUpZnfqMpXpD6xURhYUP+hJEt
VZcsZF63ja9rB030qPIgHePbQP6tDafrEqcTOGzJGL1LHUdEhqEjyWQedLafqHio6KMY2DXC4V5O
E9TciXQ8nPvDlXrfVDGRcI7V3y9JQqWZv3aqZS0GdJy01PW4XaWjo1jBk0+fgK80YwnVccTZHCb0
FXMeK4yHHbU0ymfpkXiJcVsVWjr5eNkzWOtD5gC7wBOreqKhDx8Kc7uCxsiNGVWc5Ibr+bDyBqyF
oUMhEvj5bFsSytdx2IylLdfyF4peH0m39U8HBtm9KqMkM45+6W+jIOg4nFCfwvf2gxhLwDhIlOun
CpQY1lXi3xTjn3wNX4BCCssTVtHx92nYi8aNJCTOMauwO8GAjCa6maK0A4odSSJCc1i5+CfWE4hH
cp4oxKtPFdPRBgaXWvaRXfD9wAaQZkWj17TXKFtG8ej1Ym3ODT/hWYzOdJ3eKkBYtTMCXoi9tCYg
dvlFib/9NlxLh/Fl/tPKGErtHMWiNt9v+BDXIWk77WYxuwdZ+15cxSAaQqYQzyVh6P7J/17wglKs
aTiSYVkfIqd9bMdECEFbyDj6xeESi80DvdYD/YoMyqbXKdAkGwBe3GVE9dcAMR8JKL7nSWvLdcjE
AfKhwrMZ9opN5EVILyKByfT7lXYeOB4iJCm87cbaEU1sUeAmnJvzxEnL8HY3BCCtCjXjw5N255TJ
A6WVixXZZ8l5rOueELx4sljd3JireH7RQIdqpjkBpZAPyT/PluOfMkD23td8Lfk1Yp2yc9dIwdRg
fy7+G0zAUYaiBmFTm9wb83106w+/0Vghp+Uas95WsxdCsj5JZUqyrSNiWnzS0kId0o67GXJy+svr
IUdKWylsvVZFoW3YlADmJTZ6slJ2J70uJAHj5kWLk25uL7FxNvizd9Vj8ld3J8eKznmyvkVJQl8A
QRBaxcyoNXSADfUFpIm7DATuknqn3f9fvZfZVWNIOaZOOqyXH7IL3nW7dZu3M9lOZ856VbWmGGVY
e2xoih4s/+K0xWvAups6VkMfWD3NwAZfqddSpD9TeG6Tt2dMKhO4mz1gwudz+azubD93vfhgi/06
CbgRPHB65OHZrmQmwCfFOtlPkpLhVyRD994xi+/2u7QlR9HcfayRqM7OJFDW1SFYYNFddnOvkUvc
SwbXQgzJgpnVmZ1yWxj+9rMWByDRW7ZhHsOTtXUVS5Z95QmoHiDEZldZyG8h8Ke4jOXW6gUQW75V
02vAKjfq/yYfdzsxL+TYjhYrjy4miANNKDIj7bAUrquz6tVQ7nEGrHZuL7PKDwbHaiuvlALMLJoy
oGBvvXK8cjBLiaHdmGoj7Y1gkl6URlpdJFIOEqgnZQUR7RreFCHgM/aYMWLg48zBlWEjH7rHtZml
KXWveCBRSTUwb7B2uOs7yZuGG/hX+6OO1xH6OJDoawZkOX5RPGUWmEhl9Ssq8Blj3/KZX6SDhBp2
Rkqek2wDD8boykWR2mVSq3vXkpB5kcbErFaAJ4gooN//RMmlluMBIxIPoXHXVzEYiJQWSWOR8Wgd
uDW6KUlETUuiNtvTx6lyWdDqTp3iEsPG3BhiIS4xjt1powqFFfpMmMR1dJ7/OH3QJvlNf030JFHu
J8UFC1DVdwJbo4bhlJxZq2mOOWula9rJXvdROO/CIdMMaWxWLQKXleH/QY9QJoH1cARhHXDdaGcb
wwQ6K+J3EAZEoYjLmjFVBGbIz4fPCFU5ryP+D951yxY9rFcb71k925I9/lRzurlZUujllb/EoojQ
k4cgSrWZd50S2z/jfkwbZioKI7W67jepHoalkNJsVYxgr5fYZLJzt86tNoZaZfWKoZxyHJa7KFUf
bNB3CbHiaTgd7uNyA2ke8bMK3k5Q+I19pujeDuQUuquNid5HOGjYjsujw8QwRd0z+yp55nU4d7WD
PwkPIkJvAvDtf9V5TC+X40Tx9r279lSW3grYMjl21j/xrsRa9d097IMOkmocOKTYx9P9BHU63l73
7vS76eB8335NO0OhBJl1UMybhzuXKTjbm7hqhNp5eN1gi5nV8gNq/siPTmUFGVrMDqlZ7SFfGTj2
SYU64pdYaWXLzS+z2rWluhr4WA3iRP3YMdGkHOsy8jEi1EqdKvCoIKrGan8VlchQDIAtfgPNRUEh
Jr0eRm0KLAp9wMQejy5w30cK8Hy276oVwVm2PvrZRmepsAtHUZKmQlirUmW1OELnTbZ2eEilZM/s
ZodBkdwVvLvsOHLGG8/DKf144RHY/HzRMTdAhIoWcaEWO3ZPTDPX9P0tu+kztG2oTg4jqWmSeMUX
et/Qim5lxjbxp7kZZdw4LOktG+rV1JKDHMto2yejFt4BcalYkLeDkKvZyPaZySI5zvnG6NEmy32R
9eIP9gyLw78djLxDVJklDF92J+pbacgGWm7hpQut3m67xo6u/pCzsi+BnBtr4wdm/XAvT6HNO2jm
lKJKVJnRswjuodRhmNKrRNTbDvbOtQrmNXOnpupJDiemFGKthcRk0dUre4L8b4gBJEMIpvoLiNY8
qhjwQqZAa7Ur45NYhX+aW4BO0dSoC+emvgXS0dt49b+FQM/V0xOYi7m6ZcsHncRKmEyl6Ri0rAfZ
OvQdoW27xTm70GLfE0ek50l1ILRlEDBgd3mY4jzMOa3FM9G20zhFFqxu2DYVL3KOpKeqyXFg0y9n
TX2i9bLpqxXCENz+oXVCGit83tM5okQd4ovex/cRhMKQj+uAMS/6DiSyYh1EV5wmwY6wSHJ8FYB/
uRozIdKHaNlzxbSN3jMw5DSiq6FR+qsZdEiBceIELI51KGemJm/I47ziku9OX4mIt9LEQ0uAb/Tb
qy87a1HVauoUYkNo3fCOaNZOYWFuEo+jpDF26o6IhbjXj0nXJa9sszhZbZeJ6EeaTMMZG/rY/C7d
ak80agrLSw2UMXRFW7ng5GOeG/MfqCSVgA60NfHpDRWxj0IhwTOw+P5p/5D74N6fM6S25hJIn/Nk
cWbGMeqo/q0jK2DnCs/ib1ufwMfG8xNGaceARF6+AAdz9LCx9jTLUv/Avi7CpksRvOffmV7tsjrk
j0+tAEJfrDdqPedU7shZiCX2tDl86gA20cukbavzUflOw0OUWISZMtDjiAf59ravoI2WwK+b/rfb
mk9aIIyjKjjzUwnXBNWy5PJuJBsUp0FizXIdDlJF2Hx+jBZbBjFaiUAOqDNBOxCCNF+A7gbKoOzv
anK6pd5FeNVarQzrzkhNMx7yCDemkrq111f8j4zX3ESsBIqytx6draBjKl8Cd2N9rYxW7dDtcW2C
BUuSWRf/VyxJJlPkQH2SlzafKxZh9HmfotATHxcx5u8bWPeHFw+0x070BG6jQfrbvHEXs8BvSkPK
27K6CqSG6FClo9JURgQ8Dtj1Bt7qdqPOmYc4Vm2i
`protect end_protected

