

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
VInMykl1cb/eyCcstyHEIOqfXLtsMYAK+iioa3bPNZdsHyKysw1sMYrwKEQhbdDvFZxexFV/BuR3
E2V10xNsGQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
cUXIMbq/fNZtj1t37ez/ki7n1ShEuWgIH8yPxJTOO6Au2Dmq6/c17dbZtzNOPZ13Y79JsIBKn47t
AJMl7N429e8DmdtbuhhwCbJ38cBiFdxfH1AfVZI7GGjMAdNcJoTCbcfH0JfWJ/S9l4OVfdRveiIb
dXW5fh7twSl61WcUJpk=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
WHbKIifiSnVyh9VOrHbsAOJaiYfa+g3aWjT672CoQFGtZoHYX7lHrwPeDjn9R48BpRkqqMyy5V1E
kZ30rvMKCifKQNzf0TevcVrl3t6QqBIPZj7dsFAaWjY+3fu0RTcnya994wdnAwJ92k/2t3MWJiFL
8UCO8DDPNY0Xt40qfK/53oP7zxzhOh1lPvsgCruLCaYCAr7BplNWzKtgMfwt5ZUX5jp0hTpI0y3m
TFH3zhFRvsKAbe3q2U7sLVIx7P0al79lRmHpf3nBQ8JKs1WigNl/h+LWFmAr0nyU052Sl4nQmc1V
27CTe4+On+Y4xMsv2u/myTqMuXN6bcLrIAsu0Q==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
xu9pS63o1o+cY63azBQM+vsKaznHACPUqoNT6W0vN2jhydQX/sdcqaY0W4LMPjU8g+1LDfLNYA4a
7f9gcYfJbb3zaKr5Y84jP97vWDuvkp0JSopB7FwosaQhgC9ZFFZSHrzYGBzwuhbZMni9A5RqvV2b
bQteOe3Z+NH5ROjD29Y=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
rwUkytz4o3nSG3lKXYNGBGGd6NQin1yD4vxAFncd1x1HAH4uRN/6Csj8O1eFBSdgBZrbzYpSigyS
irdheULjGWq2hoVKG79mqHugwoJaQ+RWNnILZnDjYUeFGEu0ddu39e4LQ3yMfBCfQxRQcGTVly4Y
EDooxEh83Mu9Wm4Uvi2+2y26u2oEwtbjgdJCVoicm+J7JrH1l744lVTCHFaZPWdZupXmaLsbDTF1
IZL005EF99uQ8TMXRMkzqTgTLlajCuwvHoYLTNcLy8P1f7qEEvcak6Aw3luT9m7/agpHKsss3X26
y4VegtaqqF/A90Z7VEb2715YgMpxzFEM2FzMyA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 15264)
`protect data_block
EOWAVLRwGFTjVn4qIkpMa7Bm70t1h1+/P1jPKco9ucPgLy5HL2SLYrbNZxpSYlt7se0SwywYJXa1
t4je7k3wwjgWbONmBo5F7c4cwkwa0Lw8CZIHBJSTLboLyB8G+sVDdXnAJh/T7qDHCmxyLPMbOdfj
k0n3P4nT5hETuRShfR9LFtNqV41Nd42El11xT6R6Lnl+1hGpLEn6jAaoOWmK4sY5tNjv00qJOayv
+4hwa4YuL+RKiWsK7JOSr2A9nrmudW/NvTc8axO3d8ybrBf4JTzHRCZ2luW6VJ1sv0IpLNfSc4xm
o8+BPvBwWbKpSPsDMu791CRMpMDhJxHknC8tzYuGSD6IbVCnf280vuY9afAg6QGSOwZdZuoKH9qc
Jniez19Cs0TtwSDP+6fkQ+IlWoPff03kPF7O2Fgk4seJ7xbzASS2U/+bkdcFzBd9BuuQzYOp/8i+
d+GLr9H9FZEfIbYdccUqRNhvGg94OpokWmph/zhYquf4yS8IXbQUicOPbcTBW+v5xhO4uBm9a0SA
RHHqO8F6cXP/sPPVQH1Ioh/ADhTfgnQJu+HXh/p49BflveckiZcCXO7PXSBA94WdESng4txlQjB/
F8bnXGJw4Xr7Op/tRSQl1DOXXL3WrrzMryF33/T+LTKVR4ud1sWIUtjt6DFMWqzJFZjWtcigDOr3
l7cOn5W6vnZYsL1hsXI0yG2ZlNg2/iTpBUQnTxxcmhcuxt96Rp2pZtSaHS73vvsrEz13JMzRswWi
31U7R16X1iwqHaCqbV7GTNlCtz1WHY4aO9ETxNn/Ya2LiIPe3ooTPmcExLaiD8xVjy1s4EkTv0CB
ckCmJwh+zXyEsz0ks2ox020WVQQiTKmv835jPXfIMiMTCevvII5SvG9tuRzdhKPnjzM6b1a7Jcj7
qZPu4s48jj/23pQJoxXPr+V63veP+IpFCqRy1bRm3wTIP85HxDd7WGcQAPtMeS+wlqnyI8XRyjQH
smVlGs3izZyK6Td1xz7b76BZJBq0c6Ft65EwVNxAu84/12XwnQEfs15bUSvh1hKuEv6+NdmNwuOd
eJ9jliYLgyPRp4KexCDLoaY7tLGQJMlNlbZbf+km3TdpPafC0JHOruQ2JoqsBNKkK5ktxoD1NfVT
FC8cmJjovD6CGQoKOAEL1jgnNH8VlHSxkBcy46Wnxz2pFiFsJspp4pjGccbZvntSkxw2l78ccu9O
DpKhOJSj4OZ4ZoNp/VIox6MoLrk8CLsBS9YtqencM1bKjzELQCImbMr9NKO2vsY9doj6Bj12AWI3
zVAvSyOyev3a0z/HKZpgPyDW/x/WxA3IkSgUuZHkLr9MlFlQ7Kl+gv0RFXrAf4pmREtZEWa7tof0
UDobupwxeW2CmfkOE4nxLIzViIC0uXJNIwnSh+DyAUqci2hWppnXbUzZ9QaAbd3f0sA5cLpGgPMB
NCBEGoz8b+GIeX5mHEGTUpKXDkRBNqX0O5YWbhTuxR2+OrctlNlsBpIIM3M0emeSSVdFQjiUvIfp
6xnHHNlt1NfrAZqyFdHNZr4eBzUQDoIfJOJzlXk6+VzCT3VQZYcUGCf0u3EXctKE54CJWVwc/s1w
jj4r/RCHnEywVbr7bSQ/W1cWlju1BSq+bYYu9WqIciBTz9BArrBcScCwuvzOqlquOlOVrMhfdraB
/Bm1+2ezQITMg3ZSqvKYsdQdzz8jRPCFiHFktXrnZ8+dTRZm9EvQgVI6glUWpv2QqnJStN7N0UIM
TGH5vpnHAeciYvkjkSTHSbJKlxUv839s+I5t6a6/zD5K9uwpopDynWv+lDynwLSHoBiCR7w78MDT
GLReZx1D0YNhAM6CKpNdu0jUCLsXcyzmgF6lBfZVlUAX4NrrUEGu7L7usYEJvzXHTRPLQJMDNT8N
k/159WJPmcMSJThS/KQ6PwAhd8RcaSELRgETGBZDnvcIXmOnxS2tqRPnjJmW+ImfpzcRkhGviXFe
MT1d7Zq48dj/tE6KLGpDQYuqEEuG3k4Ms/llemA9Y2bhHozJtngI9Bn3EbVFqzoWuTKre4dyeYqT
J3cwW5hHxSa6gTbc5ZK0baH8EDXNyEMaP5S5IN5g8Up6T3Eq8VHKKed+mkil3mZTDiZRqAR7r0kc
jt1YOpgve0HMCLd/MsuCms1YeJuamIMGfnxiW7Yez8JQWfp4cHb/9CkoDiKTWpnkRBR7IG4HsAc5
zJ5h9vn2yYlFrYQb3/7YgzAHK4oIARgrUUZNFGAa/mbvnLv+etAxpMzokxe2Fvujq4+54y0UmYxk
R2n7flYnUpPo96wZFglfzAE9Ujs30/tp2sWGSPqERZmIKB0PIMeq35MWoztQZOjUEwoNyTNKaKAJ
4Z53udDfmAjDNf+Zf88wlIi6QmgKdybZzNZgD+kVU/Eo+e9umnk9ujEyE7i4xtrbrI+oCA0/NOp4
3Z/9omRcjO8s5flAdYQxsyO+OplHFhyicLaJNKzvXoujPKAQi7ztYyBufPjJw1Ewu8FbrIaETJR3
Lg0fmh9ZwvnRFuY5fWh260zDEbk6mRXk4OWkQ9xAWqCyFC7apefRi4M0w2t9omb9zSVPZ6tC7wAS
xs0K9VqZuw5vytjFy+CpxbYQH8O8mHDIvrKts+CgW8N5IH817yQO0vc4TS0NBGG4oklB1uViTdV3
5Jy8DD4B5wMBS3ycwMPwrxBwxxNZp6zXBbVedhDqzndQ/c7I1t8Tn9ofWo0l1zgihdCGYs88uDk6
vs3nR5LEq92DnUbsjyhBvjZj5EZNp6/WGpwlNI4QXgXstAA8lros/Ixk7IaPawsmk4WveeHi0nSS
WbXX0RakFBIoA6WJIJ5TermH13jvI8SEIN6JFoc93sDZ+/pveAkzlicb8KxB3t50wzjWgOZd7c/7
TNYbXtc8Cp4seh5gEVR5DIjSRrRQFUPob2B+Y4pRyWz0QPpiYzR8Ld+jwUx0Hjfpeyr5JUpNvcjE
1gT7cGxnq3F7rsL/7h2XA6ziN2DPNEiuD3ZXc+df1RGTjqF/go4sntHf1TaK3V+tz2KrFJa6JVR6
zP38X2+/WfOoJqHZ5ESJ/3R1m/j6HE47WjJqJydwLYqj7vXyZVO4Y90pGjt0Vqdj6zdN1q8rVkYj
lTX6PGNaLwb5zcW1+pxiBXBkkmRKqXVRjwKzuI783PkZnG8i9HiHS48vkNPwdUywMk+ru73xpQRp
jQgrlGWt3hcr1IQIcDuRHh5z8HbzEU4mp3Kf75XoZeTvNp8JjtqEThDC5qcQ4C8nSgabYh0Ax1ou
1NiOxLMpy28xC41UIMOLdENxFKhObtSQodbbQcBrW2SkqbVH6f014EFQdB6SA2G5Na1oSzuKG+UC
NPndr52TmbvMWGMP/rXg4NMnlbbe2XL6+3QrsjjsspTrPUD5jc7wYWbitOGUbUe0YNIAzKxzAfSx
5pCDPvNpWhwpqO+KCuqbDY326klpvTXcPdbi6QSwUe/L9LKWZDLn8PLCagTidV8A7tzk96VlTgvU
3xFMeJSklac3px7HRmzmWCx6Hc0QlotMsVJ4SvbzfQjsvqomyjP8Pn4xAmzVsfHmU4OtaLkjGa9H
biLK2n2u2N78Xw/ZUiXyb7+tqfmZSnnl95myDRtrjmw2kJvj9UV1Gpqxg+WYBkiBaFRjh3/N8qi/
YM+GkjwGDlS48+84v8AaDz+DUwgAxWmE0QU6uf3BM/dxG5D5dRuEk2jdZSpIFqoVZtHUkxcdJdQq
4VE8pXzf2WZd+NwJDjGCZPaMJ84IojaqkK5pvTkJ1sCSzhzdNCAZGL8uoWB/jBLvQqymiHs0c0W7
G0JzEv3EI3btIaG63AQ2YHr/LH+1WmJSJeRJhGsX5jQzP7PBL6AIvdvIlUzKm1WTni3QEvSklcxn
nnPjtZNyFCcPumqgnGBQFjqG2mA71mwg79X0i6E6bZCL29xYTuIV6zjToaeMq7xpC+phr7ksnian
KhfH1inQ8nufOvZ2pYm1DAl+J1Jv0B57D5kCG/U9FHftZyM39CmQI4owKHBPJK3yLqMXzmFQep4p
k+xmPf0uzXjbC/jsn9f83n5yPLuqx7YGaSlmcMCvYlh+OFE1JqvyK8qETX2AJY3QT/dDd+uDll/P
Ie3jjRFp/t9CRUC4ANQ97y5Tzn1we0DpoNBx2K5vH9WrddEg6K5APkU7t/Izr40MU7qVuce9Q574
vSwAE+YVadzaDRkyyoMnEQbTL5L/jXBxy6m0cBkcpp1sVs8hvyu/uE36k+VbMH9zf4iTY8P3+3Iy
Dt1WqoIgrQCsgg4FBkH9LiEZ6dw57OwcFiS2GI3wWLIntK/Lcv9J//jFxAneRbAOdhBNTfRHnjXL
Pl7Byw/W9J9lnn7YicJfwr9Vy2u2QCDsHpQgSMxTbYUqgaYM8z+FIPHIro86+BfqW2ALSbCxtFPD
gSCw6t4Z+aawx/omylMdk6j16bIm7oaNSrVfEbUslUYjGpGSFdKfO6jF4bkDZmqf4wvqCnHhQ+Ek
I6IJAfqXX4wbw10wg2vHX94XREYd8vQ0YxPYDjJnvZgAg5WndW7PH1grVwg4kwOE0CkbWxyKXLJu
RONnWw+5xC7RzYE6MByG9d8CJUoravwK/heg+JP6EPISWgFPEyroTfOn02Hf/KTSC8zdCjVLHet7
hfv9Y/GVG+rzZHfW0HGuk1YS49dn3WmXQioROAfkyqvlIxhhBwBjFC4aiZN3s1jHh4fCtPVAjNNL
MIwLC7aCdqg8/9I5YeeS0TweM1vNQ6Mei3KvyzoQDSrr+qrmPDK4iEwY+BCtZzRXhfUuKEHTLRYP
vRZPHZHKkmDetbPlLAKN7aJ7DzhO0S+CGazcx2K0LSxOGhWxa9EjjQkzFt0uu9ypaZF6tEB4LMj+
nTJQ6U+xhVFH04kAd8YIpFoxfXlprsEO1ivcGe+Z/PQygD3hZ0kgJ0OILWU/i1ihf4/MC0hCXLHy
QUXHU3YZQTAYuqoAkmR+oPIHoxM3rM9fBLZ5YZNB2Hk6hyPz3Rx0+Ncvr+EhRjxsYWYwVqIHAn6Q
HQdylXNiA1vyXtibrKNfM7zD6yX4t/vBkbgrHSzOSpMZ57OX7s8e+FWM2hUj8bT9/dYBbWdP1dFF
RcRD2RMOclPb+vBoz5sYRTBFT4ASONVTtvm4fkwuIpsOVs0FbnUlaTDE8d6KTaTxqFV7u42SHotC
8r0BF8lg+biFAZIQ1k/7JuvIMcgkEdKXJlh8D+7ZTKhGsEfHsrp1+detDIg5eGK/WG68lHpCxXFH
E/v5nK1kot7vDRjyugmkonkrxMTevu/SzhPrjdLbqYhHFc9JeLgqbWQ/Y7u9gLHhaqN8dARct8H1
sUQwy7dCwgPDRlfuLM/ALjwFYRWQSWU4ud5ZlaUZQyH5SqnoL+eDcqSSStkIiWL6bfA28R4mdHUA
XOot8Hm9XeOQ9OdeqWp5v8ZLPQhsj7inmDI0v7BBhdN9Z7FlnvkByqZaS9aLjIpBbe8VhHLNAjg7
7MHe6pGPlMNj68ApLaP5AgsFcY74ntKBKpRg7f0BUVUjTci1YmyJzk1s22Lo9b7VP4t6gKogS5eD
KgVlbydcc1xL7cC1B3hJxmoRwzSrKf5AW5JKCWGAcfMUU7PLi3MuQsQHRbclGtDWiX7QZKpiT/oa
CE3oyMuJZu7NRNE1a+iUfKgffQcJBzI1yD+If3t9QAGh0BywoyYvBsJqQvPIDBGQRl7ZpOl5Nv9Z
OzfbT0QjJFcbjdAlI3wBtzyALCRD8hT4CfCKQtih7mRV5EVNWWLXrGhtbBeXv77pDWSFPB5WTCeo
Klskb8K6A0CPbbXJx/sijHlcrSXVzaWZIfVAzSfED548weFjuEsWCKL5pa2puvBe2F9thOPOtRMW
sIMCwLT3TQtVd//6r0elloXPTJWGjh5N3nVY/ETu/agwWn4UIUwDImog7w1MrItkuXW/Cfgdoo3I
WrnVdi4BtrE5PpIIZUq58t6ookzcmbdFOjk/4B6CnmLA3eNS9Txbrevsi22sqPpI44YDhI5Nhxli
JXPtSzZZBmosbWg3zmUvdyivXJBVV7LoLF9X4XAkpdOvCXVO7ActfaoT9AUpgKT09SYlpYhUpExO
3qPZkn4EC6yURL2BzQVwV5zKgADf7Rz04t+Y9Kng66EtxhVj5H4cF0g3fxIcGPLIVz/YqEDCrlXj
DimgG9mx940RXbVEzlIq19O/eo+7VokHmn5x6n11XU+Ypybdm1VkKzX3hP1LfvKskLls3bfPqTIa
zi4/lVijwjr5MIFTRJeRwdNXY/EIWEkB9eFu6cd+mK0eW85pHF4SbPW2C9EaJE0K1/QsgWg0vP7o
zIb6UQqABfyLmIxvYDzapisIK7BtCdhSdranDlAVeyy7zsKuh+OMTX6qv0JuE3kKd9E3UyjGevWR
k+qL0OD7apMhMAP/daZnZOmSeKV+TCSNzJdVNfw2yCiHYKwTXFCbQsjrc/qgOZ11Z9JLJNmRhd+W
HdFYgc3M2SfkImjM9k1JHIUzamjN697bvTKs/yRdI9lk4tVfnzEbNVljjsWyTUahd29uJAcBbKii
ZSHSpK7pgHQGIelAoNMm74me+GGKOdSdUsuYRWLH2sjpW9l0YpAULPqF86OWa8c6NLhWFOzRMcFX
ixNZ15gVo6ZfZF7jjLqeL2d1JbJVTrvFTwYe4haH8G3HwfdK9ba6IC73cN8GwwKMhVzuPdrFQ37W
WrHvExB26qg5vTw1Y3zt8Qp87pTvUCD0tlJcnuO7C8tPXv3BmU8RLMoENtZ5EDZfUcQZyO73w0jX
kPoCNmRtrp+6PvMLmg2COmZjnidq6y2A6jaEc9fft/vuUlKHJZmm/OpcrUYlts9NtoVtZz6N3D3R
mT16Hsp4F6bMLMlRMDBkAws0LZMRlUs0qs/bJnwGrLvlyBP4YEx0ka/FFjwR0CAykzoUwBqNgkXR
wx+VPOo/GnM2Se6knLtZgFDhGapLNmGcLhe+ITOZY9gxaZOYo6O4plVQUJrF2N25i2+2oRYbo6td
B7H//Bk+roHlpwDAigf5kxhPJjSBado1/ze6s8Jw/e6+vUd+rV6utTRuQXgXpE9ou8aHaZRae6Kd
8cwNP1tccwn8rir4KG5sxhY/dZgPbZYY3EgX/jvKL6XYXcUStGaG5SgsV3qs/l8s6KSiSndacgy2
Cd6DYGCyVQu1IsK1bppUfIDYzsakK8y7DfsiT/MrnNvA/IMIVe+GxhXicX5OMUMr4r7l7UORvth2
yOGH6477UexbE57jLI0S7/qIckaPE/fp9WvYc7wsq72KcDMvIT84MANu7ufaaiKi4jlYvUI0+Hhg
/NQEeg7ooJcfYIfGYI2HF56JWYxtDTiyikrfaiVpeeaOoOLz0DrIghHW/ZBXiV3z3bk40xhjJRHC
GGxCUL0k5Hc9kyZlea3gmwVdjyPi1LencCwLqRdZEv1C1dP/gmYGFHtnyX/Blui3X0ztHMO3/f1p
hGo4RSq4SXnsBDXJddIdqfYMcFX3XeM/hR476O4Xs0YiSXzZNDoym6+u1m+I8shqUghh0ImVRt+R
+6liyJ02AquTPAMiI+izR5QaMOm6DMcQRXdHtB9urhtr5iqMCkP7kz0kP9ax8aXs5gZbl1wyPasg
++H2SXGlwoJS9XmnSTX6ZBrbqckhDAUWB/vRYQc56LZdFRZ6pRFOrwAHOVnzvxGcIxpcVLVOZoIF
Oa7kbCvLNCF/oJLjVleCUIzHSsth+reg/3xdmchZWSweXm9odd2E6qi/HvL7zJhHtrie2XTqQPO2
vSDUhqIf2iW5/P5Ahh8eqXiZFrraDgGBdA1hXrLjBG/kHnPZLsBWEkeTLaCC8lrtP+yQXpR8GAZM
zfH2bgDQihiFNQ5VFqdbn64X+BOVWGIPi1+ougRcwW/lobvV78lb4Yux8qFf1YtphUkdBQ5MPMaY
dWnOLqb/qhJORtVH8sBgbPS07pFprYBCXG17pKb5/uLqJNlFBpRpQd178sMoenVkU4Qi+dtYiLxb
62zxvp8Kp+i6w9li4RkR/vGWBvt0KTPzrwhRQItfcUEy3cLyJgViQh2t5V960GvahG4bwHSK/6Ii
xzBL+LqjdXsxCG0pn3PTDVHQmyR7miafHc/5x9LbzndTFkZL4f/oy5OKAbjkSid80FhI3OWUvVgY
y6eIRurk6g6QIXdmXrbRf4Vw6W8lWiRto1BWxyrUWTdV0zhEwDgGohrcWdyG7/dmOHQR4QI7zRLa
5FJBvFSBf3q6J6e8H4LzlLgZp2C6h+IstLUTlTAcT5qiSD+3nV3w8a9RDqe+H0AMlRNKekCIZq0C
OjqsayQfePV8Rc/JzSgPlw2IeQLDxsM1/QUGl/5M3qGOQeg11WODtsSK1tiMZBV/NDXqloxoLnQe
exe4FIBqNaZt5rDplj5bJoTrcqs9cg1h9eXunGSPPp1c+mYgBR4bketxTENTSk+vlcyUF9fsFVZb
RwusWsof7e8LlksPADjQKReejpXagSCuckBLcX+G8c/+CkALcu5GWxiLza48/W0vSQ28eYCJPmwd
Y6Vh95ljywFH+c/Kd4qhet2lAlftcP0WOyIw3qke2pmdThaWYQaNDNIvYI2sF5o4MbJpzcpIDqn8
90uqZGREU6Y6ga9xiH8/WBRf4XlI7Q0uOmJuwMmeUmSZ2P3dgt8g0KlrHSr1PR2Lj/w83Vn4Ke1s
MFHpRbgzdWKooKSuzHLLn6iv1CRhKzLcBg+ILTX66V1qlD1QKV56eopeok84bNPm1MpUG1xz0NTB
WbHby+i1upfuzkJRtrZ75YfpGARtLedYogROqvixe6ksQa+8/qXHWrlOEPGzQ7jZu4CaawRLHEnM
yZUyTSgIyZjXG0ZfsgkxeEY3aQZvSaDVErw/UBFebYlvYoZpYRN3fZ6/fC5mCVno30kDE4T0DqFJ
UaW1JLutKdqrzLm5hyodUPabWYxLKwwxSOk9aPCxJuKmA7Yq2gZhPPcfhvR3YWXQHyba6FkBYGLI
h7HaMpWR1mrYutFZwXChyyZo/ZtmCubIx6dtDaPGIzU1x0kx7O5P0sMylKZ3zdWBpGMJkeNByuwG
TCwCUF0iXgd6ut4EbOjAWkUgF5ZxcMemgt0sloOfKO+xWCSpulw0BmqXWXKESGIJ35FfZcWRmZhT
w08/AN1ekk52DAeb0q0VoEdvEq3aGP3qp+MDwRKsU9TNOdxm7jBbwLY1WAAQNSBVoQL3ZMFYY32U
9JresICBRc/2DbOLG10IpCOToVwA2AT2YYMXsWT0LXr1KZrHgBUOMqxxy27q6pgDk2iKmhw/WZy4
hnnbu6B21fKFipj7+LjUv4i3nDJlr2IlVqfFQrDLMQnFFuH92SL9mRxtPZBOSSm2/B6TKzhRFlD7
KzoAm9bxGS07DaLT4pxXa1qmvYfeYI/4WFmjKf86UrmjlyEB3M5biwdyuUojeBEarQQN+pe1YWye
GwVKNNXMEvhoCrKq8iLBJgwzxJ9rpZLSD0pZoyLmuNzVHXpFhis/MxXbQV1l+1Dzwj4Uiv94PCZV
YgL5yeKfr4plt1T3Y2et0CvbekmVQ3wa/16b1pQgG5x005NxTO1si3mXx+43VE0HhDuUmbBJKZyh
r2Me6WyKNHCPPHAxJRZK2AojPMjZJr77eGy7mbuobdatNvjLKLv9aVGTWwFiYsDhqjFq2AM9uu06
nr6DO0yHy2RHuxWQIsqtYWmPbXxPzclgJwtxCm9mXeUr8Vb6Yc0p1BkkxAq05eXbDyCJOyuyYVE7
zavDRSJstau5IsRncf65mwJhDlqXZ1Osbs+TCDG3VuxRZpk/vA5nOLQsL5buDLeTadh14qbRgXbV
Qzl/xaxPhKVBS3T2gz/3X+3Evi5O1G5KR1TLiYPRytHqqBjogzzGsIbTRPfB/nECGJTYVifQlqoh
cD4xUAx3LAPOkoM2oUQvjw5b9EoVgbnjyI6B0AD9AdJG+SCIp6+1zSMKIV0UwqFej33ukc3lSkGN
3s8HUZ1vIDhWNlfSzeNShqsawiMZI5Buu0xZ3s1XOlPrO2Q+T4BVAPmWCu4wMFzfnvhNj2cCkamh
yDwjk/eEvO7J7y1HopKV7iVcj3EH0ypSE3afc9C3G8cJ6JY04l17k2UxdS3ogwhsNnmAyR6FDC9l
KUzFVneL0cRHVf1t4D0Mqz1NrQWFLHcNAauj0s7pzFnWExlL3nIP6165d2WG+HhqrV+r3DulcFo4
fEHhtWgeJmBvjO+tFitzuE8cXwbl1VXBTfU9fcOSVKKV7DE0Wp8HxksxvIWtZmdyXebuUd2pJxji
nUhkRt0AI3SODeELlHQmiy6GMrlqppojqWbn00k0o/7ZXR32mFyL7H8hYAL3yELbocbUbcKGVVcM
EyakIY7vrf7k+HSb9AxfXETGQOgR5s+spwXIERwo6kcMyXPvGYwtZjyytGCuGv7o689VewldAfKz
EmcBBzlAMt9d5mKvHCyDOh+jGYGJPhCpzCaoXdQzF3yZVB5FjVb8ZwJ8TppyatiJ/iqc5Sc9/Tgl
XGPA6LpvENwV9xbhLw92FSlvOExn2qrnzQeaEmfH6v36bp2YfGOho36bjXb8QsKauDDbrZnjawLI
Cwu5887r3sMoTdnm0cb5Y9ssAPoW2zEIwz92auttcfpszsw56eK5gW8uZtV9hTKnmP1olKTw+81i
qe0xFlBn9+k2S+zVaTAvjLB9HGUJZHYp/f5K6re5v9IxNAl4PTmcaD0cr5nMJY4cJ9riVPUML0U4
VJGxlkHs/JmJWpIoRC9UDJ15/9pCDHFN3FR3lZ3FXfx8M6XBLMVEVhUrMltP6h18+vo09yQgP1O1
3YrDuUi/rQ7PyzqDFI4j57rRviqBIAR0am2o/iUEnXrNUbDCxVULVfytIlx2ZW/V+VqwwmUoWKMh
Il9BFVoGxsFHWiQdnmTnN8UTOsi3/VO62Ep3J/ciwIK8I0V4M1wfsWsbFGoW8bnLNCGGmcad7XrY
M3c/f7VMdLKOxJ2Ds4k1gq2rm5RJ9E2Dnn7mLEyapAxfKxHBKClCufdb3wGEPlHy4RDjE3m9+ecD
X4Cfs09vOe+CL0R3IWM9iyeRgDh/LUgBf6mj1OqNWdAbq3pl0Uo+QMvjnAOJyVUB2QBn1zGfKxkp
eDRB8PmmOCPIBY9gtX3cQLJVRFRa/aIwahcy51/dEgA6XeAd52+gDQ97U8s3l0foYSVSXuY8FsFX
fsgJl5EPBffTKpmOwmI7qyOJ8QWcWV3C8ezgW+OOP7XZtqnQiOY19d/MU9dgJ72GSUtOWEsMNFxO
OP9CKYTcCe5oHUvOYkVKfr+fgXPLpt70p+bBFNtBIQL1HDe3Gn7huH+MXzvavyn1WROol7xe1TAm
D0aJddQlSBJpLzAC+bW/xwLkS5ojAZht0FXgwzIp5Txf5qntPskKWbottkHvzlX6SKNfkBVZMohw
HpNP+7Hjim1fQhWjkKM74u3XMu3y6in6YFs+Tv78E/TpOz6C/ErL4BaFSOOCrBP3gurjFxhyNzAl
yEWMdCPVeadKXWEmKmqb0I7Cj80f9X6uGCPGBCt9Hv6AkLrblVfC784CmJQIgBfqqNTMo9Bx7vBA
FyaZOJWw7wu29CqE5o+Y1dMiHqXNSSCyqh8XhJ6X18WoojAnJMLU9+yIs+fLydkJvA/JZ5LGCCLq
QjzlOcLGRDqBVmPVVYRMyGqU/7joauvmKYEEVE0OyfZg7vANJ3mfpw9K9Tyb2fgIqAHzRoEo6hmD
UZuytFLsrfrZLVyUri3wZWlkFd0vcuif5oV+4TGRY3LtcpAjE1nDaSlN4Y/+JPiGBrY+RfTbCc5Y
rsIr3XHCl4o0v+h6hBHMjbAQxDT9JUTz19uxYJMAlT24CvCwe0BNzQGPvzo2vt2ZApgcVkNenCCv
0iOLb0+6Mwp7vIXqY9/HGGXrRFxFcADV4o//d3dBjytDrtbc3ScjM5HRzGQBwEHZzMKZf4kzeIkZ
QtDfozS4FejzURUM/jp4RR7XQGOsbgaUtp3jjKTiE7/wpPKgxXXqxD3vTX+1MTiUJXQY6Gy9JKDK
92XbTUFHBY+JVvaScOKiwZP91OlBFGqWTWcgMhNEpvM4j4NVUYWQfI1gLaCRn44ZA2vuYXrcSzfC
uRGdcCF0i5Sj30Z/aEXq7sqPnlhc5kWIa+3C2SiEVDONjB0ymKxk5MNr0FYjInU4ZYRZtUYpbV8l
m+5JTA33zRWJrqQMMn+xZFA/J175Bgzpb6YZ2FNLRZyJXU5WgL86fxdvNE04zwXQCbROEBpO9clQ
MMUShYnpUaY6GoyfR0dzuhbTgnr2wvw+jv4JD4D6JzMh7hfmSrKaHUMrauuON5EV+juxJLlJBzex
YS+O6uYFe6DiVVBDAJcPEraC1NAj4AgQDp9Fn/3sUNBSyp3RfT9ORhQCL0sdCedCDtri2tut4djC
XOT3FKqx5p+5WdEq6N0geI/wyO6yNJSFRmPSv31laL2xDz89khMNnIFDMBGDtno4FOQUyoyE9W2W
bGnYdmTJaZ+vrhwKn1fasQLb8+7o6ExcSolvz+bPdrh0KWgCIUVLn/jzVEEQGFi7UZ7JuEGnbgSd
cz3sYOyRAlumNvYPUBXFN24BYOzl6K+OwPyTx6KAq/6Fo1IZ7hnFwaj+VeVavxnLtnEHX/TGfTxI
aQ+BEAKThMFYN/yqsacpg2WIKL6kGtsCYDoc/xpFx20az9P1ONB7D8w8A49ENEPa1L4+UTJZHLT1
pAT143HGEeZcuREMgSiWVE0qKBQcTFFMcHRPF+7D0eqqtR3n5NpSl1qY+fOuZ41EXene1kqvM07J
ChNwLaFRR+G4kWRq9pNJvq0mYDmzFx0kLifVodZL3EQrYYK8Jpmd8VqgebdHVVDbbjLkGSLBNKKW
jpPxYA5eJGfbvekcnRrtXmy2NOVgFJoPGkr3cBYA2igjgOe/qYuweJP87KqoemUh94zB3pifGHuX
+VicxbM66HPsHRJtFBsUcFVaKQLReLJwdxyuR4chTFBi3Lxt/pWGYd4cp/ObACXfNAb7uDHN3+aV
qMidS2QYfZOKlf5qx1fRRFxgpkZngnUq0D3hNxJCW6pm4egG43sFh6EXSXccyOljzSkwFsH/O+Gt
JGy0hTKVevTd1dgnImOODeQUzoUvdrVZ8toHVTPlFfxZoOH40noss8UgJfpBX1o+4EeOS+6EnFHV
zimQxJRso6ktaCfpKUIDDxX7lzozdcIHDEtobEpaMFG9CK1uHZdYMa93M8dUoMlOHhDhk+YaGK12
FC0k0reV8krNtJKYh8Z9Vh2vGfqRbmoyn3ZBW+4co2ifyE/ErJPgqDqSUrDGYHmZ/XIcPPg4Wt1s
/4DlgdAFA8/ZGfz8I2pJTD5T+2BaVv8/Ozc374l8kB9vx1t7qCz2GlQ1ok2HxgzgDxuIP87PHvsh
FLMJqyFwOAJevGRTq6IVeD04w8SL56I1vFpLeDctD3gFGmuK32pv4d5kyiInL613tpKt0T4BepG7
5JscoELxR/rg9MV14iiVgBnESA5cT5KTKbtkir/5eR4RrE3Hq0GwewGIqdv0+5TiY1RuvOMeHM0B
w/YFu98ztYLPe4+9hQOc1wJGvhK/Cf+oU6CXFjwN3iQya3dg1CwYbBsAgKoeFhRapTlU/noBqpHr
Sep01yBGxbybecEdlY+Rv/7aittu4Pbl12w2qaCnODRbGqOa+xW1s2BC0Q69WgIrAUF0aCI0cUX1
Yb8anuS78kds78YM8CaNOowCuPMB3bNJMoC+oPkF/pHZxOsQaHmr+69YN+K3XJEfEYQcljwsHRru
UCHpuMWhLHItt6FYx9bafN6ZHBkjr0zE+Yf0lNbX9AGxe5Gkt+gl2VWC2v/kk0d4NeTqlZ1qk1Cc
NhwVNSWxN5SYww0gUd4RaFYkCyt0QDbQLLikbzhcCVGVgKr6qOcvO0scpQi5sAEjKx1aY9VpZY6+
FQva0lKc5QHqtrGQmWJB/kgKt/6/rYUxHeD/2jDtvp5ncNsYTWmodFSl5pj8hNWSNu1WGfplLz9a
3CroUHitM/WV9XpqwLMB3o8aAl1pmF5otj66OSDSd0tXjcaESgNFDo565XxMWgmfK6zq2PuJZqc7
WtUBQcELYeUFiyyGrF9leSUCPkzKGyi+Yf5NBmCoHuG/7j1ifDC6rhHVlFev0TaoAKyKd63E3/gH
3NskgbqEvHHvF+FojDHYjwyONpq0ktmyhbWSckN3wXZOg6qqeAMNvgfvXr4b2YzUhMzU+DIA1Rlb
YX0MXcHX2edLdPI8VEEBJPobPvmk7Q2oGGPa3xzEOE9KkUD4ds7m3E+yT2jTtq3cYB3wPbrPuS9V
M+EZByFrdalkKe8Yv9ddqcVr4bJbwdn+PtQpFDMzKwwukzJQm/ZQI2/PA/Pqg2MJ/GCBquKBdYnK
i9KPJiyQU6lsqRlp5hW3YniLwC73w1ms6041zPlY7Hn9G/OqxVCbZRQ3t9MnVLdOClREXcu0a/Dg
bP69MSfSduwNjJjQ3dxY4/SyhiFxLQJzm4tagWYCOK6bN6y7p6aP4JfXItKBSw5u/0hPIbV2Dg5z
1tN+qS6zIDxefEV8r79zmqcMnl6CKe4Ru+ng/7sNt0bPF6G2kF6RUDqxaz9qlVrEvDnYDz7X/ug1
LF5Ww9SVi3TRTEdHOOWjdYWdWqPnJvX0QrWE9pTsnbwbHeWOYB3lBAIzGXgMKp5NDiEml79Wi+fp
LZIZ83ALerf3YQ44N+iubmHr030vE9Ghl+ep8g8uNI6RORylVLjHhUVqRPh+MDzcSr780HtlULDf
rSmF1Kag8n2tKBmF3l1wE1tmE/iXBAjGPnBgrXJkHjkpMHr7X26wnL3Quj5fxfZBJuyQ0OWE6R0k
kJk5jTftZdbdGvPWC83q2SffsgTdzN8tgxWJb2CVW/S+21462IdV/qq6egOEfH6bBGYMbdiRCjj+
m+a5gvxGqdJeaybUe3WQHmhvbfzHlgugla/K90uRtnhxP3QB/CVNig+cQIaZdziseFH3TDiv2Bcu
KMPx4O7mmC2ZgreGzxXNI9nSMAiEtii1p0Daj+qWPM0g0J4U9d5vR4Hjiq9y1UzUlzi832mm51F7
JnBJeQLAn0vqkUSoWVxpdCfaOXhyArTH6BU8AXTViMaaWEO3Buuk7QI6NQC8JEjQq9bzU3VPeBKs
78CRti9ubi4UNw67iZcgU+NDcZOEWQwx0rYBM5wjQtIEW4BkV3WhmgG2yVBvBgqXaCQ8hnVsjR6K
P+o+LSQvDNcVaIz0zZwjVZ6aX4c70Rte+0zgIRJW1m+fHtD0eQpG7CoJ1AtVPZm4ZiIpiQ59JvAY
33GJ20joYsn5v9iNAuKwLnCjENTej43Q8kVzINk828YMj3Ym3UyxIat7+N+CgC5UzV/JhFfEgawg
RbyFjzQ0wmYRKqsiPdhUveHSJhUnwFGokDbPheJ7qreoXOLrgNyJRBndlQRQ5SA2jrQ5M4c5W17h
zuX6vVGQbAJe4FSvJrVcKWs4BPVjTX7cTnF3uOa68vzc/nEVIpawOsnoMzAkiUyTlDDzvOSzSBm4
hNvpZDuTNhQ8lCVeEyZ+KE1wB8VeJU4LuE7wW0+YsduVMBRe6m+HjM62xLEeXwXxiaVoKx+NRE4A
+rrk1riTl9Z5LXnnJRVahxVAs+zybdsj81s2PZkBZRSXBKIByQw8evpvBocpu26UZiFe/vGirJNl
4kZ+3TeKYEenh3LyPODzLziHYKS/lhdMf6/RSV5MmFo4lHOCTeXhfWqMJNLs/Mn9J8Z3zRl7BLrs
EO5Ee1n7pbwuBQjKthEVDz2K4BSPgpBC1kkCKIHzGeGW2PGJoa3nX8mWUCjYQ97EhFzwuYclzyUr
dKJaW9zTQzTddWvTT7Ouhky3bxrL+sblLHVpjM8sspV9mloU4AD3MrCqiv5vBGF8ZIy2hB0QSgWZ
PxjxQkJT1Wv7Jv/7h4jomL9DRvRtb0xUgiheb6jrEhltHFb6jy2sWxvhr7rMfb1R2CQj7h5sHY40
0D0DKN9uuIFY3nI2/Dyah3/QuoBp/cmolq1LJd1U7Qi+GHLL6P0iInxxhYG+AOxi0q3NisMS8hyy
eR1n+Wpl6FemZYj1AElwSuDDd41BKgI4/Bz1TQOLAYa3pEvVyZ1Y+ITZB9qm5+s1sH8GFXXvOKcv
p5W88LpTnOxxlyM9VoV754oBD/1kdsfCuhrzRG20buvb9EjEDJc7woxBUPwmRC71IECQVjmvCbNu
Lc/FVGFlvTgwc5FW7DIAfpVw4osRM7rHxPzLW6tXRBUIOLiFPa/klA9SIV4ZR6ZHJFM5lUqJ1HC7
bhjhyR9nDWNEJWG/nK9i0oYAtnVZEJ80WQfHi/Wd6lbp180izA7E6vVlolVqOpAeo0xqm9nvb2x0
Bm/TGKbPWc0VaraRppO5A1MTfXdRrCa0dT1uM62deX0qUG5xOdh8DSq0Qsaff8mCjmnHsAPVmh0u
7JRh/kuTSdEhGtXXhSjdVby4EgiqWv4NcLYt7VPEM8ow290wA8AUOvTKduuQr4XMsu7Ty5Vi8hVe
ZnMowiQXjW5iG2CZUPoUWYdETibjitb0m7tHFRutvY9eGlhY2v4Cjf4x6xmjtwxmOxCAbgzkjWfI
cKCB6BgqkPI22lgIkwmDwB38UlJgumIl6o6coNKjXjm9E8NfOqO+qceMuDOdB5DQZCue+ZdhqsfA
YUxmzNv/Jz1ki//9zac9q9G8I8kTh9s4BsZxcMq+HzPkkFHW0zbwiIAr6RFSumb8iIqzb/qAZ0pd
mr75tGZ3H9ysyTIsTTqrUnoOZrMpv1aqWHB88BEuZEbWn3z9DUls8sqjFZBl3uUcU/2jZPCwv2Jo
qJb4Bq5U36vATkJIZds1Hj+5U9ij69R/NyTCZb1zEWCbHPx0o8YSlaUGZJsRXCevTp6Rgc92Mdnf
7OLHvutJS1MS4OeJ9qY/Xr/9qu92O9ijjH7jGmWSxsP/5fYc0WCJi7FmWR0M9JQ5YbpUoC1D4Djs
vp91N+Su8IBuiezB+ZjgdJ4Zhbe5+MnPXSJlQF/qdjdUu2t81ACMfNbsw3gC6jb2ifG7wy8xi8bz
ior5mxHmegO0BdByJO9mnKOvUaOctCa0Rgo2GrbCthXo4jDvo7hqXUK4oBpIUU5q4WokPvF7hFS+
tZvMeRJaYrBBPi8WRp9i06VwmdV47+je2lK3TrJCQY325Non1iv4P1u0txWbo5ntn+7HK8U0v85g
hPiDnpu1BetnIQlYTpxq47lZP7DRjOMnK1ULjdefDooLy/rgQQVrXPc9GWym3Z7R/bKjtA095BPw
vOtkQj1X2b1U+g+EFr4zk2TeKMPrdlxkBC+zb5OOg9JIClRw4G4QNKTCSKLfn8ivE+a5CtJQ31Sh
SN7wtjijypLnAA+Oj/H0A28SmCVsVG55mkg2wScURxBq9yymRpFSODDE24ckHSyHu/kSkP0FFJI0
8iFIAK9iMwEbaDPz2QSVACmN+a6550zA33EFqwmzIfzGiP9OJwPLNOxbhU5eTEqTn2RJrS6ULCVG
9lbW6Yn35v8ByDs/1kSvF7aATXlK9TcWQ+Rq7FRVFsJ0zGYZICM1S27hUdskd2SKygidrfkjhzWK
whPFbnAZL17g/Q45xEr5UKocuwjXWPBMdgLYv5K4iu8Hk1OtsHTLyGtDpoBq+jSPa3WcKGSUD4wK
7YrAiAEAjDKQ6QXNLlftxFweXTsPQ5e40opDSuDOP4almD39lDhkDCYzTogmag5yjNJt/uxiJpG9
Mi7lX41Mkyh5RtOUAmDNjkvGYd/gt4d56MpC5EVWVLkwVSMtYRYGC1dejjUkrMDHnyToNJ1q3GoY
YAPguFvSZoXC4UZ9wXUl+YxndGT304u4iImomzD+kF9SZuNV5UCF34rh2Stv2biJxvBL/lr7XsXq
tnHSG+NXu1ntx8Co7Z6VgP+zg6obvlYTAMZCSHc6A1mIfTvsQCkeDoum6oiS2scJr+vpJP2c/HNc
+StNCxDmNRYce1Xa9w2kHrNiNUk4zHex0nwGMmQHdb5KhyxdyWFk0MEWU7/vXqku27QT5B7R4ilw
eUv+IDyCyEUjbxIIjfauX/TzJ1WtL3NN0uvFI5C/pfEK1xRm9UQiQd/cLaGf5DTvu4QUQG6jj9/A
q+GT9YXcJNgL4aGv4mm5Zp9z0tQwdsXFlL+xidUdaUEAak6EdMAjTY/SRp3j5+tgmvmtJTz6Pqpq
AG+KcGegdNZ9dPQ+ROf2E17BMCVegFH9Yk9WmtYqV5oLV6qFI5lrAgSfOPf9SdIVSVBJDvE15Pwd
hj6c7ZV1qkAojdwmSsJEoKjRYXejuixQs+yBot/st+i4JWV50Hk52cyTkqzrlXgZyzt/cMgLJwEO
P4Q1uPC+jGU7X5vP/OQ2KLtFX8ByRRUbvirjmUNYkWIn0bL+Y6CexYOpcTo1iXfqbZJvItZU4ioL
Bbc/WwFx8bqgq+Ug3A/VcaYZ9yVQIe3VhUVc4DgbrYQdPEVFFOy04dnmyED8p5xCxekT2Rm8/bpM
kQArFEqyN7r8LAZw5Ep8yPNcEHXbfVO8xEn0cFIs+QriqnoErbQeWpLt23Ga13BA91GD1YD/n9eT
J19dtf9G+t+0HyDHAT1UtuXqqJDMFBeruZdhVHK7vB1Sc5/IX4lSa8Z8lLAr0sw+n03zy1tWrdYU
Z281PW6PywctQCOp4IU3i+Rv1XXFEjYVN94JlzQUQeFsup1n9B9ZD/eXmeg6G7pV80l2PTH04VV/
NtTBPH/4fGAdJ/iJwlf8MLQb4Zys3QvaqmnVRASGaSoqSKB507YMUSATw1CQUYcEUJKLm8xICdi1
XgZ5euFZk8uWUYeX+5JXmpFL5tT4Gl8KvRtXwwMhql4JCvkiAREjPKZE/qsqOkAOtHf3OvK/n4Ul
k8XxvGgQl1+nuASCsmcRD1dyuL19Dl70Hs3QTxauicy9PpTvHbrJD60yo24IJpxbZvmCXAXddnH0
dscds8F7SVqUm38X/tSwNdMqs/EB7XmhLNhHYACLG9z8/xLodj5kDRQAtXqShg/7NzbQ7m5QM69Z
8sPBx4DHTU6qFRaiCJRJFDpJVm0cIQf69R6MS+42GwHaMDz1//plKM/B46m6NhTjhR1EC4pttr+E
y0TcjG5mNgalQwV+7YdPi8qoe2udiZoYAugmUdDl+4/nGwphfk+QrAYI7dxTqrH3JW+nBiHluZUH
5XJPVKjGWGA20tgmgZXxPoE6MLCR6s3Hlt3CGai1u6KQ7fefDH/1kHZWYlyVQZpy6JPXliEfpHwL
QVjvIjIa2wmxOXpJlMxCdedy9i/Mxlwa00XNbPneqFsBv8bDF4O7VHAqy2oHxh2G2hfNIZtF/L9q
hsLwptsxGrWoWyt8YWdYIsfKuN2yAoHj7RDAerk0C5zjaIly2LXgaTWJFh1b686VsePnNjYFcHbL
ceFHDbzlRKuTwPCEPFAgFklvkqSuwHWGqgrLSOBj3Wv7SeZtgJqU6uTFlGsVESRkE0xId6uBV8/o
zh4nDc3DJE/yxUrvISu7S7x2Cz6duyg+NA2m0Fm+ZpuoCDegZ32NSR1X8HczgtlM4PSG4zPkB0KN
G+nI/eHxtoob/MwhwftSs+PLzi3b+y8aqvpEDxlnM0cmvVrySyBsPUiLE8rjukrMFREl/oE8mvMa
I7ylPXbBlDWJFDc5cFYMSF3NS2B8vZfbpIm9vBjWmH07HJNOcpP6jMCJtJSRty+r4AQCePFZYMxD
9UzVwW0Tx6BGHba1ynBkp6mTWnEeu+sHgfpyXUFcZyuQm7cEgfV50zeFC/ZyJOadyN4dt1cV874D
gLBW8tPd7CKnaAAN2sgj4CEv1KqecKeHLr5HdZLza1ZUYt00FRJ0WQ1vccMbNWSF8k2bifpMStqE
UYeMw5lPxQ/BKBv2mZqJ5+CNKJ9wUCuq/O2dEtUu4wr/qn0nn+NaWIXXeeN0l+p8Ne+Ch7dC75bA
6YgELHehhsV56HJB7d+YgdNE6ARV1Bo2f03r9zaR+GOP5ghkFYhYzgmerrMtEKmJULMTEqu/8oDM
dkdfQmJEsn6JCOIU3KgCg/N8psT4bKpiknDTb7ogHfRKOIwZ12zEiUNd+xmQb3yHbJhlDEK2UujB
EYYb7Vt6RGUNinx+9eRp8wZ9YAZGv+v+bI9GetTsBnAlN55TLa9Wtvdn/SVa6tyEzJ9UGD1j2Rfh
SUbHRgFZQXGMWvG3zhb5XJawEO94BvyNz1Xejij/9huHu2akzet2y6qY4Ox/0dirMzJcfiibTH/l
x1ShVK4t1yf27uFNLhPH25a9z8l+kLa8fn08Qmn8KYB8MFw8wpZGGLgoT130y7c4yjZOw3u34oo/
LNDQ2db36y14EVWi+CPWcuzpVKuSbDXAtVWHURyu1BSvFknv5RrnDs+UtVru
`protect end_protected

