

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
jPOKnt2dHOagW4dFov86UptHPGMdrE6d2ZgqMnfJehhzqeTiVLl89did3kf45SSrRMnQy9YGjxY6
jqpfslmzag==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
TbXlwhQ0d0UG8+CBDSNOnRgRBfh1oNNVi5QwoMGV3zJAlkTsnTywwNiy3IArHTxG6Niq+d59upyT
QOuldsHqtyc6KQBpxueCYJG7Fv1OIOGGq8mGjrkLmbJVhJEwBvPv4mlhsXKQ+/UhmQDpF2ZyKhkK
EbgpRIm7ap2EmEdPduA=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
iaTK7nKuH82rPJSrGYALVeHLyxEbb+9Rh0wJiyQuCqzY3/f+ne/dT7ytF39Hm0BXD9csWKwQp3QC
vOqzo1FyLi+w9Ik3lkb4njvMdZauHueYbVoku659dslyFGV84Aivwjcg0Y5de7FqsEonjWrVPTE4
0oo4m4QHuK8VN0pa+LmuzTIHDEzIPM6IMp8H0IstAk4VaGHg6wlCrG0u2kbbhcyaOKk2xzxiDfSu
gcUy11TT1zHFME/fHUU4VO3aHMSGacP3N+kgMah6x7bBUjBd2rfEXkVcl+/1g+qp0xW2BzItYrMY
Q1wtoE+N2GipiyxU+AmrXQ4zQNqO11zaj/N6Ig==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
QkbQ08NIPb90+bNjwXDlVNk6WbvhfydYhJZqryulAczmjZMBvdwitIPmanwzKj9BPStsPNHXyOKf
9PFA9l/uvQOwVNRTz3G2U0+6+YFy3j+qj97mRopffETTpncxm/BoroKpRNN1DrgSjygcTkfrt06N
1lOXW+551KWRUPA+fGE=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
LXGnS/C7HF/SjGcWlSWMUKmilNZr5UhJNWaaWr/ybus0u0ctzmNkXcydCyfmEQe8OngFPF/IKSaG
XMrlZODcxs6BdW6TBJGvkBlKfbvIYg7iCmAit8JvgZpuYsROJrZ/IapJ9XCUZT5PW0Y/S/PoGs0O
fXalNP4hoIYlP5OYjMaSowkFFmCMq49fHUdBBmi6thqlMFhrdpbAhfGoJVYkjStWry+O4YcFvpKw
Q8WXsOAh5J64eppUG0x86EZ8HpsK6EGAeT39tAy+jNSSIcnklat3mhXxMF+BE67OS/DRt5H346yK
YrLlKC5qbVgH7HjzWMBFYeVVtUec0iic45xLPw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 11232)
`protect data_block
o8QgSLBO/8wy35cATgA3myUqbIR6Itf2pod6O514Grb34QCPCRgtdG/EPegq110DgzN0LqMvYFPt
1w9laQhfW74K6d0oilElOji2MoplgsKF3+ng2+ZE0GFueMtIlkWth5DfXLz4PtjWYTrNUYSG7K7H
CcOJ8GdrpN2wZEJ0M1np/qCyPD7L1vqrIQTpbAF6VBml6poew06cYJGDDIHZwFJbEw5ndhpY0/gH
O5SYValNS6M36AoGH3QcJ55pHKuHE6mV+Zcf6YFUIwuXOJSNsf6srp/pGoZHb8gjnHoxDw4MMqps
IZ4bvSHBlI2v8M2TcppLdcOc/9xBlsh8c4ktV/qE0NmnXzFJownjWNuWdTys4UHzZDFx7L0jqcb/
hdya9mQY3iHOLs7N0EqeawwuXasY4QggX4EETW6prnIcheiyvPSna92NGmj86M9MBDuRFcjxwnqB
OvhywczZvVxSgtOaie+vursQemB3xj9jrYpIVMRcnZsPZeguR4ekdr527qPRK/i1TuAnJVmy5dGh
Pd/DPigPio66GAWuBSB/MJNMbuo6yn+sUsJSNGhoNh7c4f5Q01IlPHerwReTwxLb7G4t6SWesNP0
LY4H/cIhAEc3Vzco0TSULj4osfnXYcl1L0bxh3LLjVG7BTiCyImYnnKbbXyUoajCKwdghB2XjZv4
iupZVywTWHgJRe0NwPlJ4c8cnbUkMM85juaGB79wUUP7DJ0RVQDkmeVDhyRMXahT6BbUz4u7IxK4
vRft73bn8IhZhos33lodzXnx1taLed0+J9862S5F9skHFA8oGxr/LickKenB/kO4tiIhL8e4eFLu
OXakZ6Py2ZVTWrjmtzcpwerNgqvXB4lJwZoZTqGudooeylvBVhrDys2gI+g5jlsMg/KxKKbeY3sj
10K33uAquSeaWyE402uVLxhqAQUz0naEHvCuAJPATXqcXg3DFH83M/vWMPdlq3B3n2/wWjE3Vg87
V0yw54IqMq0qUdR7dOJavGg8fKiYxbOi4iP02Smusfru4qlMD/93y8nejiIl+WHepJzlqJpB02Qb
BNphrXFYNhi/3dViLzaYtcuuVDKytBpKiLZJJQbDaPan9PTaC5pl+kl36cng1puqoqVTicZWu9SZ
bi7iCRdQ3O5p82L46yM2vENdYyDrjsg2rF0DK9Xf60asCrRNOhCvug6vAwkR8wt8u+h1TfPDGrtd
m01tukSPGkF7/1b/eoQvJCRw26uMoDQ6AZGAc+MSw1eRtTwDZhCPaXnR2g2ZeiV2Mpo2mEBYYatr
BQI03DC1gLSb4cmk6psfxF+lgQ6pcNyv3KjGDABjUJv+rrHYZF6e1jXlxF6clm7skw5+GxcfwzPs
dfE8eUjKmFY4hSUGKDemIIlfkTz1TOicTflSu3v+cajrFUrVdvO8jCq/0nz0tNfv0pMhc1zUInzY
US/WFY57nPQVza5cHEcxvlFFeMgx++qyufxiwn98J/Xx2ZzgNenGbDXria0DSmloJhYsLtXJeYC1
4iTHOpgeAlRizxNwzjVgSnwKeSBDFelQ6WlUG49omtSkKvS5OIK00XeEHvrmZcWvPXK9G/Xmw4yc
wcOJhkhmTzZYSOh6Toq+a60oZe3iMBDbddg+KS8oCIeRDxLMnNsy6bSPpGmnFD8RZJhP/6pgOuB8
kNrIgzLUHSagfNfJpYx8wHSF/dtjLsWABTsmKQd4j4xQzWO6IpiRYWB7yRNi8Uk97lIrjBXw34qo
C05+/Qdfw2aj22qt6mOO+uk9dQU2jldLv7P26X2mT6+XMXoW7sSugAVBkHHmKILRtb07r810teQO
PYFLTskk7d5mzmHxc8TT4Rtu3H/PAV2LWGK5UOuTMFXY5gB7KpNLMVIocDY9gYhUPEDTBnPrWMSw
OlzibtVnO+dvU0MxlvtSPJcIHLxa2FtpJ8PAJqYTCUh0Ky2AQOmY68JEeyQfy00VPHERU2HOz/MM
Fko6pj74iU0XpMrxwhYXH6v4KgLvQn5NU2WfvhUIArCRtXShPAo19GYKng8cfeeixZmNicVMOEbb
F4/EVZ0/3WBHO0z8ELLK/Zw5xFIMND4xwdgl3JXj1k3rbGBNPSgTZvR2CoQW0VXcLc7ovVmlnQmZ
OlCgTnjWWklpmxQc6xxroWYjJRei+4uxeAQpygi69ef4GVRBkBcdHllQ5FFZvynBNX5jgr5jaT5b
rRnKwXHPVXUWVeEAN27drHRAoE17Mz5B7pApJKr7d3cWP+HBkMqOOd1VFZjIFFnklsJX7PhQ4rJV
TtZYtULpf0G4eRLQCMWCtivcIlveBnjS8QGxigk5h1WBfuMyH7uoC9Oc1L3KUSkCMAkPLU2CT36F
kKoejPFFrWEKw//YH5/K3G2AiOnSlqZTE/fGOIovn0JtGoRPDEb9vIC98sjXyH4f1NUsCeh6HyYN
QFRB9q6jPBDDKBxMJSHQoPLSh3gBeraiy87UV4NJXM5MdZTyhzC08KnTRqsKfIQY3yzi5nIkFIr7
bRkP1NeCrKd5EFUsmQq8EN6+qv+1fma3k5oSi64z9pXv+Qt1baTWetP6RYVtKd7/zVfvioR37VCV
KddWRcHnQKQZKXCHUenGPmGJMqHRmuTwHoKGr4vwSgV5GEVdl5PXrYobpR5w4hogZEGrjH5tZwsH
fBgZrRXYYcqVAn3mMawLmk4wt13sU6HDPqiSX2tC95DZKtaksymRMgy94dr3ueOxGLsFHpo1d+7n
8XQvUiBvf7D8+VWCx3zlrQnogezYSbfon5ea2rbsq/m2GtwIrXjyi4NG5DHUoygBnMKMf41AhfPo
AmnTMoBAry3UjgOszsLEP/gJ3T24CYoh8IZW/NEnVRMViphULNJ1SfFoQHypCi62FTwCTEDY2Qj7
G2/JWAWXv69TnZsvSwug79kf5M+qOn2RCs8a8YV8cXYCCa3A2OyqjioURLxhzyBj07VFjrykv/tj
6hGWcsi7ZrJVyCiopy/borHpRsNZSEi59pQ9IdBsEz9nJejJyQEqmaHaeIOxo0VQZQJrIjoZRjf9
jtxcywvuxkT0AIkAmbSRZRbrqp/9ed19vdO//zeNnl9RnDaip0nlGQi3YVYS3RDi0XCaOt1MhGri
H0ZU2b3Kg9OTbJNQIFhSBJ9WUUnRqo2htu4vw0c0ukFmbths0odIKxBJp8vEPUxR4XsCh1Fj1LOD
HwNkvczNv9eNXllDgeVAVGQSfBsjRBdLgvKtvcYwJsNfJH77cDW3aOFQNWAX+jIumK6i2iEYt3zU
NRYoFf6O0/I0T+4gZeUHOn/SEa1wyfF/HvpMpq9EXh0Dhdcff1n/kOp67CRLd1EzJeHMxE6OO0hz
cZn60wpjcptOLj9JHBbjdF1jxtDh4SivJgCeTR2tw3hlIkKA6RXOR/ndpRjjrgMifWgUyqehpN5x
OeZYrk2qVZ9gj9p01+TBH/M0mGhD9rq2DJsrfa8HV8qYtilOEbNSqt3rkUbirBIjOakLvRYQYOmO
6gsUzz/xZdBUzqej/E6Ro2deL3yNkVf29Y4GCFmyNw2gRTFcvmYPTg28ZGnJyMhPcWBGRNUENq4O
zFcb34yGTsvlIZ631lTB6rGgusdLZu+wJg79Ipyiqo8TnDn4OGEjy8gpMQktE1maDO41tNZubD8H
9ETadeIN3l5AuEDUa2vQLqm8UbUZSgtSL7k0GnjEFOPKMxSui2PbaK1u1Yk58SK/Ah55o/pVZ8yt
8ISv232fKQqgKpxwn9SUYfewcJmaBFgTql7HJwfghjFnrQ5xms3U7Z62eFwKiMAnMxdPWRKFwSOW
85KrIVO6IyastOWgEALIcLCOD60rmDNIbO5i/L0KCBjLZpmC/rZi125m0Hspx+6X+rTEh2k/ojH0
JCfXP1z3NE2YfEauFSR5VLrmLe1UvSH6XyPoPiLfDrpgCMS8r5BPOBTqxZ9lrAgcKj2sgurKGezP
JdROcXly49FbcsB79QrqNrFWthiZaPYXwQkwuN1rDKWh/24QKrTIreOFp5MzFD41YoaWyVzre7NK
ITYsJ58ZY3KO7/G1q1oyasgarcoTSvbVdfs1lANx+/7N4844nP9kSmtwOPRO1N5OXNLX+45L0EVg
2ofjoEYQZsB/32WdqwKYHVo7p9TK/5N2qB2J3wz3evWVtlvvVy5eMz5MKNOA9QMx8fSOx0V6TgM9
SM3RyyGgKRy0PHpiRLV2ImqlObK723TVWSRDTHibEdFIoBos66EX4sSEIPnvhROOHOrrOyX3DorG
J4kFHtzRAN8mRI22EtSCxlLl7EE7LNsdH1GOGLZ0d7P+aBovQLevuzs/S9D/iy4byW9nrqCQcXJx
E/zHWlUeMAkjLov90wvYVrlD3KY9LxmU23F1uM5AVp1SqgIYLkVc/VNGdkrEwGTopN/V6v5YdeeN
N/yuCC+D/ZbNi+PB2Ek1S1Lt8dk9C8nSHQFhFqxJ6xY24BLJvUve/IzPBH4qZfi8sqG9Qp3udC7M
pYwZlHrRRjV7I2XxlFKURqDhQQILtwZjScpx51Hl55MUcV/SKLZEkJS6/9FoVxHNxnTrqBR+GlRU
D1DmLwGxGzvlvHd5FaiPfqJekIq+RBR5qfYmKbTQxcyg0BHu/fSsnaAh2kXDgCQqnFWLWIsT/Oya
Bi0Nuyqt7OMclsp5Jcwb6lcpVVW89vDPtn7/nHgwW2aY5Ti3AKx/bq4H+BbLOEpWUzKFNid7EDlK
MwqOZF/OaJYxP4OHrJM8FYTEgzpWEl5CpxB8fyvVIhQbg/NmMj1tyXlHYlPNz8aw2laNN6czLWXj
EMZKqhodnLlRiusaA71QySYfhzcELPwcRhXBqQ8yalW308L9Kf6nVTv9qyjcMk1EV1bDwrri4dRU
SYJWkR1uranFVea0+vX/iP1eqxepKWmwRrMgs1A43Hr698LL9brqBEBeRtgTRFcQklqmCmrUqz2E
TQNEQFdBTlCnqCxE9AH21GTdUfEQ0vle4TvD9YYR2/bX6byoBkCSS66RGhFFEBZcibXRiRIsKUBq
Xui2TdpFSO+PBfivr1ahnWwJtolrAbAe7BSp3UvcjF4ovD4p1PxhltmxB/0RCFScSlH6Ex0LXOD0
wOd7pnsp1R8x48Zoi8IYM8xGPNvbcidIhEJOgWYDKVhP4uK43oWcm8kUIxYvCh6X0YhvZBTrYmnq
XLOjY6oLzfUtBsGSQTvD6YpxKPRqD5++jsLkuHvea1/2TwXygFolOc9bbzwhfk2sEF1dlpe1MKM7
rXfzT93NAKTmivFQlMwA8IU29QeMk0IYeOwEJaubs/nLhXVW8MTYAXyIKBvkHMJVzj5cUNFv6GD0
iiXGRMehZBE0opBfcrQNJbcL55Kj5Xk2ZGFF8W+qbHBkv2k/P/U1Utv77kDDODjkhXhKr5u2q1Jj
cDpP3MsPEicvtKEfyKor318tSdVEdko3I9Bvi9hchTXTqw6Sm9sHR+1TwulzVdqSAfw8Wz3uXSzx
HQLl2dAiIA6nb8XGE2MacEDTKOxsuHFeGUujJq67NMHTZf8gzYj3Efl/pHQ8QdnhAh+ZQj6b3Lbp
Sb9TxdVFX8tSU5SAQRsqg12d2Sp3blReZsyPtRMNuhloMimSTbVDdOGv+DaZ78AvUFzLKCz3bMys
8miL259Sigd8/2OrIWDUZ/PEgXv28FNAH2yVBP4ijMOTGT8E+TfhH4suMz2QkSvVpHXLV6UTLADx
iIocGiZy1SOcWScXzcu+K1XlkW5fWHYsMqEsLZVhhppj8Ya/QM+Q1qSyTMZK2giOmhG9StkxbAdI
oyZmm8CHWMAa9WtcJya9RpJZXYDbWp84NTg6WrFyEiz7mSmgJCvHIYr7XbjkqUyNIBDMD7QT4rH/
n3JATddKmN4euWeZNJdUc3+CeU94pGlvhzan0p7AKHc9NUHQ6XYR21rxWwmSm9Zvmgh8pzjtAP3N
eMQPKcUnkeFyiqY+L/RnpFwp90XYOyC817PxixhV0tuNbATk4qp09R5U2BuEDV9gHGFBvNllAiVs
VK2pbWyGObZ+yXHdj208gG2kUyzoYycJQi5n3x4yTdZ70BA127SxZ8ErLejtKtBofBsvnDNj/JPj
oFm1UXLYO1Cs91N03rdYDGezAZcVb6JLwNSARnCpBy74xN7Wbng0WrZ7dJylq/t1EK9XaoWKH7xj
5SeX/yLvd5t9UzdO94rAPeiG53cQBv4rEPfr9bcYc2p8qwls3PGm8+qvRzjt4fgoAtIO6yxGLvX7
GGAqMYYFhjaG7BET+ddOcU3mrgzYmffdDpg7yl7SqyluAT2+UELrnsFAfp70NQ4DaU9jVjEs8zhj
GUMzC7M+kaozcisu5X16+HbBBEVoBQ25XR8ZfgaTbcdbS6B5aFo/hAAK1Nyj7fAJSI4pXRFmE26Z
OFRQKLOc4BgEG2POZiNsMvsY8f63ggAlNxLQ2xTYdG48mpYjJ+cpBEY8/XaKIeypTif9cuNY+Kpd
qg4leM64F951X98Fhb22SXNTvTYZOagVVPOXYAYWKpWjde8tkA5MQ2H7qdbLKIibMD4T6iRXU9en
qpafVPK/K/vuKFMhIph+dSdVqTbU4vOIiBNhJqOH+WBIP39E0116lpeh4D8DuQS1cPvYU77enLsN
sJRP8EP+YJ6qMMft/c+2GvZ9SI1w/X/hKReqjHj6+w4aQl0bZBrKd824QBGgYf7k9HlgLIGG7Atr
4ynYI2kOqQsNYPWQRbq8bdhmBBO8Clm4/vPB/ePXhkeU+LPF+0QhfWtfNxcttdhOr1tYE+QDS3zf
AffEd95BuAnJJ0kOHFtE8orIyxzfw9jmoDXtQ5TLcoMyZ1ZSbDgjy+6uwOGo0pb2NSGIUwRVESBo
QQquLXVwOaFIFspIqmdOTspoU1E8RK0LcTagkaAizHKFcxV9cbhq8o66o8vd5p+xvXb9JkaXXNDf
mCNuvG6jZta9L2c/C4AsoG0X4xyL0ko5qYhNaS5UigrpYwdDkFSUrWcEyWKx2wCx01Tuywy4By25
dRAOD11HXFYRKg2tP9UkrY5Fbu/NQbNsJPKA/6DIKQAYDq4qDThfWFQ4wjeacG0WYzS8AjhC15Lv
9V2aX4/UYFZ6opjjYlN2KvUPIS6UpRKJdFYobMSQqa6/drm7EkmYlnaxDPGrOksNoaI5JFAwsOWg
ceZ9s7+Hieki2XtYaDbGtUIH8DLE6RVQzlOtJ9GWhqQo/sSSDsqLzP6MNHfwo80vlE0oyIBAdBhN
txd5nWl70fTGW8eY/+MhcHOZgcRGiDMHES9UfQKgVXlR4YNQElNB7+wUXvltWRm8WvUdCTlwXovr
ios9S/4uYTfoDa8J5BKJnrt1rVtr28LU4HfKO5TXUCxsch2+3wAD126qv6Z8DlmEe+rs0gERXqpX
61cCKFjS/uQKiv3fHsi515iw5d14/STvL/MLOqA4hhIOmh4tAULVHqTuXFFdfWGEV1sbJJayaV2Z
mzc8bJNx8ueDCjBlUwOOwPuw+ax9aAV9+fj4QX0IaN9QI0qCcv+i0HVw8w8Lg0XH1k9YxK3OcKUA
bvz4cbR3p0CK9Jso5t1UAmaIc/scJwKZx6CynQ7oU38yg4m+1nBra61UfQwjenS+h3z47kLxlKrc
sM0nYtN0fzjQrp7hywLPsGFFwpeVs8+M0ujshtSDc8mKmGF0YV9Xl6CswEiOnEXzo16EaIWG2htE
lg0i8F7kZf7f/i+BUTemQ9Ou3HNlOgLCu/udDNBr9oNCimx1O/hRzIH41rYQ6vslEJVawC9idyFQ
esnduSekT/kQvejzGbw0nUUKDVCIf0is/t++u8F3Yq79jwA/kEKgNHlSZ+r2kIEeT2lUppmTf+4B
jrwfwkGWhFI3Qv1OLDKBbRwENGRe0bDiI+FYwUBbJD68Axp6Y0dABLhWS53Zu+3HST5Obfy/UBr6
6/0Tu7OHC/2pNdd13LDLgc88sdeRTzkBAPa+Kq1aQQTcOmBypenvKIo+GogunBKv+BAAtz/zH9yK
hrEJzP9UJzQgoLD9O3sQWMA7iepVVVkmgZ3RS/lTFbOYtdZdrPXp5GqKzGMHBd4jXJjXbJl9I6Ih
sFQgLHRUil3fg3QXZ+Lz+uKaEAvuDRm2ojfU4SCUUlAMnNWwpQU7pVdkTWH54DiTY2ORBQ/Uah6n
4FUubiiex+m06ed1WbYKIb0Zc++istO1fjCJSG2kP48gAxtHNYrQ2kgq/geighve5dpdbK69cXrP
QMvY8drGJzz2JFrecbg9bVDjn5wkjZZ3qd56m8NrJHxrWt9+AWSXvz8pD4E38+rpmmnElpBsl/pZ
mpOYuEIq6TTJrKDATGRzIguQQ3tUWA4qHquIvFHvDoVnhcvFRiNPY2TIrpRWUNRtWER8Co/WkkhN
zA3zXiX+wHpCGdTZ2ZG4cCsVib+f+sk+AP0CTXAWVG+m2f1GxapohECsVk+oISCzfqY8sHI+X8Bg
J6g5qTRXeFGxl+u4DuUnh6gHYMohgj43Odyg2bfIKPWn9HK7EyTdGQcxbZextNyFNXlXAUO6wnM7
FWfa9a2a0BsEM5BkdUoBQiGPYYfQJ5XN8rpUYjhiJxl6AaaCUiqBd1Z0KGi6Se0R7z5nazOOkAUS
GWnWwSmxmTm2ZlKlQSAwP5GYdx5F9Gip1GcGXeM2jnl79OkKLc8pUnZujZ6UHYlzSh5LM3DhoLG9
SbnS1gd6MAJacGOtIIdJlQ857stx6/kd+787nlZnlCsH2TJiwW3HxH2InB9YUgzmayvdzWwS+5Me
26krHx56KM6Ia32d5FldCgNJLse4CioAtwo4ubaE28P7iAxDuEU7iekSgXfRIdHgbcsf2fwwloGk
DaoYNV0GTyUcYFYXuNL+G9/5CnEPyDKjH9rHYQrNfSpvxeBpZMQAE0O/2yDc/j121yBfzGI1yXKi
gri3fqvGB1jfjvL3am+JKsxQAEPCKFQbLwkcPBSDkmHS5sIj6w+R7dNxNRlhHLITlcsSfBzbc6UB
lo1VOYuVwFTxF7eLKczvbK7lacO/sn79PPfRE9xRQP7N3n/mUB4G42PETcrXL8FdHFbK9QoQIW8z
mui3P1ljig49QH7Uw5hFo3j5VMzO5wLEHFcH1GdCZl6fzcp3/N7ylmTUli06baqVN0m2J99gPdpm
jQoN5yJf7voZ9D8Zs5xthNE4RsXzg5LjUFcePuTO3zhSykumHcoi9cVDhBZmWeWlpvo5hSMhInCO
YiE7o6V/H4ew6beMX+yNOi+Ttz2o3D2GK/zvYdZ83hXLMTRGEvcfrQVuD3Elza7xJsMDZDe7r/73
gwiYEpA6TKdqdLuum2gxFwLmlVFjmK1gX/F/PAZGTKqDQstNWQ7Zhk6qbBChkRj8KqdHjAoulcfd
uSFMRHSSId+VeOmT3S5tsCG739TOuRAhuAJI7mMuseLhNR5UJaMqsBYcbsJIyXFx+6HimHwc+bAo
q2Zr96vJliPIqGpIQwYPWCOtH+LiR9FRFyd3QLgivzQiQiuPMFXhrKQGpzmWeTMU6cAoSCSSXLAq
pNIacmQ3SrMw0kvhwu52jdbKn1LRLDboeS401xxjjJmfj1j+jPummWnfq7ieIgGxeBPW/GWt/kjY
yRzBFlPBoR62uyfamzzMSdPpZGka5xzxQ5S+iwAlWEVHI5BzJ4NYUmbaYjPWgpeTMn3zjSRL98eX
Q4lAbdML0CNYB6ceeHSMOA0y2OzZQhGZ7lwdnvllzeyt/C33djNmYXQ6BEFOBMGMbr0iA9+sczJ7
w9FyJ4QwxhDMv0GRwXtaiGdi3qqIFNizPffXRL9S81a1bAGLs8bjq3fdVx5OqI982f471hMXIIdj
Htfek7eFNoD7VC9nWeDHKJ+XS3Iyipdp4JejSJHut6jFMN223T1aaqSblvqTx1VfJFycFqp1V0RF
ryOP3Lr+zJ0vsIkERTapEilaRg+2tHG7KSXKpQSl1QMh+PjQbnBD4vAwTOXxt1hLme78CxBb4Okt
HwWadOlU+56oTIs5sLt02FpnDHIhPKMlHUB1jS1LzxH/mZqU9o8ctqRLbJxoroNZ2pPorAZiyGuf
YjxHgjjpeopEIS3yh6yGGcnD2ka9mwW84dOe68SL1QgLV1/+8zGEkJvuUoO90s7pWiZD6/tqN8lI
yYLPe70qV7c4awiZS/oXsR7Uy0HnE3GOOkoIs0fxShREZ6/CCVJVZHoMd81roi9kIN3z4ygL3wcO
fVTkrlaGyfwh391NAPE+ScibLlN0SbXBmcEkIcMYq8zPrIu0MVp1tBtiQ9jAcrGQfV/LYCBb0Rdd
y742RdJIL8Zyue6MnQtYja/3H5DXjjCffRN/PaTQcuh0Y+m6hfwg8jhJ/fmkI4FXbiGTZKYbVNPH
PU2cUJLQBevr2LPY2WpA4rYftBScfKW7yel/+iK/QNQKYbc3PSjRGbWv3GsC1EU/LRj18BRXFDGR
V0/PeFuZf2c4kYOVYMQZiCQtWw17RrGjM+v0viWgOJ6s6QgaliB0wb4wDoU2zpBXAhHO4VcKvQdU
NFlklToGki3Ro8t4bMDuKwlK1+c7QdOiM3O08fZwIDfAcBGoXcMqyQWSIzoHDl253gmEataN/Jzu
u4idcAizwckxauH6al6P+qPZ7J9tyGfnktSo8b1a3r/F6jOM/RRQMAZBtVvsdlLcYwkQ2EVur0y5
EINnE52yjXfkzpDJPpHowDvW1NKGuzgA7fW6lEREDbjOTssS+3OjKNa2cU7e32+TBTHfpDxPhjF/
Cc25rq6Li5j9LTuHWYDBKvdYLtz/Hcu1q3YcR0yGPdJv9UEMx4HWplS5fSpyJijIJtaOo8BfIGju
TzLFgVzRWHPdYzKliNtDsLhrFZThKxi6jvKs7arSFKxo8EfitRc2iWqZ8kcrpxtmO682YQsVfEQp
wEJiKPwPzajCizMGky3aKO2yvTTPa/4ESqTLlYG6aF37zOXnQJTvqHQtID88WcUV6cYHdZy3Avwd
mAbT4CtIbZnh9A4IudMRsSTQ+/cUrMUhU+PwBOd1NtXrOdnjZzD/RxqZQ3ErICQTGeEK7JYy1x8h
ZB+rCRQeXeTSr67jq3TVJZ4JsJb6I1wUrUSdyKkHFhUwCyBsE9yH9fw/QK64dDa6uRTjEe97xTB2
6JQ3m4t7Jh4O5DlTL5LQRfPKBxGeOREQ9ylhDYZ5gRH/86NGJFvf9gXMCYYNaR7dF1FvE+QRbjtU
OXVZ5gESse5zp2LmimzxMEfbzkeSf9RHkugDbpuDEVULvWaGbrmGcac4oaJHChxuxcwRr+rVnwpP
sUYEMDH8PhRZKX1M7VlrPBSM9KdYCPSEz86/0NlvI0QoVqj7h6S5AaOZgnUO3AFQH/8OF5pOvORW
ufeIZe7kFZ7T9aZtPrgETyXiFdkTkyr/NKHtmYBUN2yKax2fH6MhtLkdrnBEzjI+jzvwNpsqv9gk
ON6J0ft1qvAlLyDJ8NKX6EqHMoAZvyNXNZRvJxgUfOp4GGxA2mQC3TsENOtelvYDGu+HGAKsz5bz
JzzAkeS1mvK2Pzq5zRZX8bpYj4BWrZ9VsZ90FxU4LE+7QADhwzSwDlBVyxY3j1yAXwLzMr67D0iZ
CcMtjtzeJbcRSxK/w9PYJ6mcTe8vTLDQrp74qjRjwqI4Q1BNeywAK/moymN8LyjPwoeqdnAyTrNu
A5P6xAeKgGWQT4uSpH3qYmXS3x07hJegvpj2MAEV61yWyVliSCZWlNgFiV4KIqByP2jAPjIDO65j
W5xJmmnuysWIREupxGiguQBCDiFR3poN/VzOHqOgJG7gKHsiqOOnwimDVL0/2z+YjaXYAdaETiKY
CX8zijhkB7NQFvszzpmj3qMvcCGf5tIfd+mZN8P5uUYVY10Sv7HQiJgeazPvA8/PKx0pEdmjFKr6
dTKF5miWr565oaJhN3Wgvih7xeCgW89vyTJat5/MHCEZUhqzjFs14FNVfot1jBe6rsMoBWbLRLjb
GhLYxqCmSvIC5JiyHfRkKnNF8F088JobG9c1lEQOLFUmOZeMzoHoIRVsC34Ba09+ZDSPv3AyOG3Y
Ivt2qP4np/UuKW4LkmTtOxKJLSHA+KqcwcgFaJoR4AM9qywV5eAr5LcUcxLT6p48iT+sRTgL5I5G
wCnKt80Fu8ZJXd2envF7ZlUn6h5/qyMJMvvPDaulUS7qdGVGzh4D1WI/MbgJSuUv4qEc7WDVCimM
Gj72T8wOMr/p0+c8wfXQf2oqKlP33nprMW9nEG+TfVuJ9/WdQoHAK/PEKNjXhRcRRoH19hIu6+H4
j82tffSrsh94zokVcp5wjW7lJ+uJAifatDSnfLyRKT/7z1Y1pIBPg48Ivgq12L9DwWbDRSRTR8W8
2ZqhV2NqxHoQL5c9nJPMc7RxRWp57mOu7JEcIIKpIibqpkBPT7qzq/vLOZZ0ASkmtbtd6eoSeRKu
DytFJp/qYT9x6vCHK+6/HeZxCEmA2+I3zns2TUmI3EpGmNg97qvFBwzoQVRdtJkv8L9cyWlpXRdo
0L4paw213OJAwOnDU/Ad6ap/1XPgCoZA1Id8hPEKxzVM9vWwJ4FFHAznrw1vPOz2qTInolbpYiL9
98e2ifUosc5hh0aQXPwGyYA9CaTuGRIpY1d+TRrumwJQ+YqEcJSJdtlZRNjtbcMswsv+Ywd99/6e
cl+mKKJirOh3VOdcjUiAD01AJDOdEdGx300aA1zzmTrrSTvvughihlnOq3VLf+ty86LijUfNDZM+
hW9saV4GiclZ+RYNjvf2VzvvejSTdav/2vRFRHBiNb2OpGEnNCcrxKmyiUdywHNMyqNus/ezCkgD
wiUQey2Ri4TiP0kYjuaEy8JkvHSPJRPRwStAOz8a/d8jgGbS1K4SF2MQqkcMVfbRBDtzlnOLa4fM
5jnyQuF5Kt8smFMwchWP3cKRaHHb9n2Ew2UDmkiIsk2WbVFesQH3px3/WXo4sewt53IR0oOyyDbJ
BMwcCErHdRcPG6ZCxTg9tWbBDWv8JOd3c36mFzYTGFY3BLXSjkhpcOxu7jFdJdXKpDHqcoH0KfRa
7l4NoJ2tMefEi3SxAgVGjHbsgAnqnmzZl2vT6ePclexyE9TcjSczNZ37PRXekkKa0f/hyWJLaB3b
R8R0+Ufb/H51LpEnMs8hX3FqS4NR22dMjePbwElSGBqZa46Zr9NlpRl1PaI7VoVDolAIJbP+A18r
k/WvVGxNdccC7Ur/zMegXDBuF3BaScp+/u6ifn0/1ydVaaiEYBAybEGFCznthIun558+9zfm1K24
893twrjo3dAJLaUqu/PeTyIamivYQ5UXzf9+dgnMe1F1jUb0MNoeZ+1wplIYSDy0FAYSsD5ptZmr
xbMjjWHJOG6n8grAo3rQNdGu8EzU/eoJuxIwJz5zsPFoLspvJu+VAtm/gTuzIsb9YgZ9Pl9K0YME
jDvVA1SWRO7BLc114/U6XNO5xElOWbnfdaUbKdnGa91h4nnTtSE8W4f5wr7zmhw/eI0LefSVS9nm
Ct4GLA8gGg4qHo1vTck+uphHQ3ONBx7gay48+HSzwhWB6ag+2iNOfsSzkdKd0igkoMMSpnZeIE+R
klZvuLdYOJE+zCLvZN6nLl4N3TPKxPrue3pyw/wwEz5WuVsyF+r3cx/28kYtIAy5OfrAG5WWVAN8
fp2Co9L1MAWcvF+RtzsIyPl0T+6VtzKx8NJJ5B+Z9lwDu7s3XCI2zh0LpO+GXSrs9/ibv0W4N+xl
Pi+uS1F2eKiYZyt6vzB+bBmfHvvp85F8UZqzFR5pGdNIAzuHImGEwK6EgMU5VurIXttWmwMKlp0F
bdOhNBslEChOSXHHcKB1iU/DfBC/A9d4XaAdfnVyj8YkPpidB/KBwUKvRdug4JlccZYXgqSD7KxC
U6YFFmW1NwqUbuopFpyZkl7fLQorshBImbNlMyTQExMvHU3M7TL7li0O3oXaiX1kRXWUQlvlTdIh
3S2nEbLAJx6DY8QK/OTM6fQVgd7meREhKcF/trir2uPEohfSsybjMOABDntTtSSLahom1uG4j66b
KymyZRTLMQHb6JVTR9Lxr8Ow6noF5jvbV6fogPQ2yAHvvDM2z00JCE3kvLWu10fyGvxBiZavJnir
8ie7VniBVwrBBSLJ/pM7zNWyzGfGnRpo2zJuf55hhl5fHGbFtinrcdL8LPqXZka89xuCiRADNbKO
8ryeOwBHs/py9v+E/rQLEKsg4etzSFrG9geK3GjeW3pazce+WeAX5//mCokOpUEVCc4pVbKg7Kyn
CdnG2Bn7a/mbOhSPvALU1v5A19OO/CbOiEc72ddxfJe2+Zj33Uu82tJtD/oMnNty9/o2w+Wwxjpa
0XSMDWzxX+H9buKTHTlfP4FPbMvGT9u77BxeSI3+KmYNBZsO2S5Fu3OKrz4uW2DD0XV6kU6y2sqd
QjIRRXmk9Qj+jmNL2ScJMzjR9qkDWaP/GAY7CpVP2ugTJPAuc4uTAsY+tXOsh2Oj6KlZf+ztaO9b
b30frewgefUGLiC5pe4jZCUDdBA7jaN7dwfcyr89KjPIW/GrcHBUDGXiWI4IxFWAhg3gCDC5hWV2
hnjogd51Gso7MuwRgPOt9na/k3SNhlZSShvdebFJgSKDox15bWTXbPopOexSkHMpI1/zsvkXd7MC
zlbt7wMkcipIH2/1WUkogWybaPzDjdilmrOAuFct1AZSEpV3RbbEKLk1QTNsQyw1dtNtrBBLY5Fy
Z/JrwQ1W79jQ/UfKfbokDKIqPL1oaAKiPq63nRsYwFvZwK3XDuEcBqdKqL6/o+hsKcsDWMc80WJi
JWsTyetteO73lrPlXY6zSwF0o7n5158xnz9aCOBDB4V+NOdvr5Y37G6L/Oo/zagyHTHXbvS4o9hP
7oDvYRL/VCeJ854oZjrejVWTkM3E4sylSkwvTA7zzVfSW5JsVZ7KS0bKXMou35MVZzqfif5iIBMo
NooZFUmV8nhrVafyiQnXxUKia5BCd60nbEKJUZDF0s2o0aW2wY8Pv0cuTQDEidq+EpFfu15sjpZ4
Of5a
`protect end_protected

