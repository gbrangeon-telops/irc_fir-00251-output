

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
jtXjITQ50a0ecf2Im0hc5gDMz+eLQYg/zzqRdEOtUonTsMauUR2I/zDZca/cFZRkz2Bn/e1TcNfn
wKr/p3+6Ew==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ANnTEQ5JJem4BDOpiZXGW1BGnlByArgufttfMLkwemXR407wjOM5c7+DduQ2B6Rws3h4VtvHo6rO
wrBVcL7VsvPq1+tV939t3BGzv7HmeOgz+bF6BolXyM301AxlRkWo/0oJhXt9sAWYr7zYDeoXtQZb
l76HOHad93vrCilEPkc=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
XmwNj23lI8XFGQYG7vF9oV5Kxca20ebqjV8UOZJpCCCr+xVAS7ag+llpfkHEOHuw9tSDfsd4Eagb
WTNoLsXhoBdOAYPEcNzU+W9qGu9/wjx0qrsJ9f6NyxsR8o/IzcMAojV3xWACKEn/35hhcf9UXdPw
jFtFMZBq82H3pspBY7rQB54QzJyh7kwXdtgWfJuR8vKgpz2Bgw+sWz2/D2DHqFf2M9nR9Jj5wsYi
jA2guHzbYFRqb3Hyb8w16e2ODRs1Chv6CQa8J/8jZZjpfNE9JYFfYFbj02jB3GIgpxkUh95YsKVS
nyG+AAIy66AvGO8wjxEaZssb0O8bFU7NUeHAaw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
jhiEXYtW8X8urAKsC5DlhfR1BlhyMUwpr7b+LLkcXXJrwnqMhkaTCeeV/MLdD2fZlxbKcfLK7F9V
JGPVeMHqW/OgkDKoPYInFHgV4dQ8+vVlaEgOkFd21VNxhDMogpMeEu/OUw7EcrJ+uVFRL9Y4CZQe
7QVrICfnVX7/1Uf6PJs=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
fOUx+hBZ6Yu+THnpJi++K5FNQDW/3h2F0eesEGevzvwYAUzmUKIlynhcf5gdgPU7azk/daFeo+yk
Krq/01NBV0vQpvK8q0FHFH+ghuL05juk1koa24QZKqKLJESEoqe8+SMhcjfeA/1/cXTmsbZU0sOR
598davhiRIPeODK4SAJwb2vC+fldvr29ZQPfn7IqVQ1mWsnCoHzWBSYPyy4Xw+6asrFDW88G8kf8
wyRSd13FqmDW+hKwsLgtlOhvBagW21tHVBbEEW2kPEAMrlmNhaLMf5utkD/lTPuEPBItEC5xgDps
hn/cW4ZYOpIgB7hTnFioHxnAEnyoEZ+mfU5gPg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 23952)
`protect data_block
gE7XTmjdasFo8pZCg9BUmiK8aV7FJitDmuKw1CUi50P6EbPh8SXgPiETQbZManqHZDiLt43+Kih3
FBzTE9Etz31+PtpTFLQs7EsbPX04xD3FTfAlfKMRreRgb54+r01lbdxDnGhozzz3BqzrOpIaPv04
th/atQy72RI6P64TVcrJ9IFVlYEQWkl1ZhIVZtR0Xctl2GttOiHT2N+cx5SFqAqrb5O3V0YDGrIC
46q2sTn/zSAd3u0W3lJ47g1y3F/bNeiD/+9FXlKY3+jMwrXmDRTOBK3QtdSz9qBq3nqgmzEt10iY
kj6kjJINXK+6T+qDJqbRP7gUyF+DBk1I14cE8bBCRj/J2zoN9QLh3GTrzIUi4746os8mGHn+VhXo
sfX7LpgJexDv37aRfnis+MDJq5m82X61dziCybAk+uSUsMJIZg6X0c8LH5wqVagMhHrkQQMbujkc
T0ogcxz5eIXE5idh0FRaAfnjmfXRabZ/GV5pjsCH2arOLqez7ri5dNk5IWLk5wxKp5Q204/Oek2l
Sb++qV1nisxEw6urN0hFry7qF8vl+VzfAfa5no8OW+x9SH9C0UFJia2aXAlO+84z/myZbtcdX3kG
0/Vluo8S7PDxfBzZkHkFtuhOVii6rFuw2ceObYtqOsNps/M3ug22XLzOmTUb0v2FwRzF4OP06OED
dLNN/rZxtC2CHAVR4IWKOSd+ncVl1Y5bGTbRLTyvQs3Z+Z8HPqNxA5Q0VLqMq1kD0dEdX7QXjvC5
kF2q2LasDNkAKZNlsZe4uGilMXtP9ubuPZQJVtzwYzhQ061fKpD8mxa3xzeTbV7Rs+kQIyFn6QN7
AAkCGuCOMkM0iTUxiwIC1OihiAx1B5XwG6p8BlzJdg5iBqmxXwho7EsY8gyMvD3Dp4kLgVT3r4ED
8j8HfVm6QlLgen+yIYecPWeWv9qgYaLJkn2ZJNAhumiXE76Hs05BeChy50Vb0WB9UaVKu3FuIjyT
l0SPE8joPojP/arsiA3MZeNk38lR5voaLHniQR6gYWe/HLPQ1I7INsm8uQQ2TCxQnq3+dxDKFzOD
ZD3afliDCooERubC02+YPPnrZmPnQImU2xdRN+kXKJTJ/Gf+RiRZLAPI5owu475Fax8k1QfuVGb6
6jz4wazYB5MCWeHEgxmGvXz/yeBqZvCWuVyvBuyAiZQnbNE/ONr/4lPSD7kR/phzM5OX08DbTng0
7wZAqQg/XZDPkym60TfnpSaX9HrBVpjPGyDc7tUVP/baca+wv2+JKLd0FMVbnFg/5nf9pQ9FPgwh
do74s5mh1UFtu9dUBOh1HJt21JJ/joYlSs1J0C0Wj0i6/BUcrAJZCkKV5e8t9XRAUBRl1CaFAgcP
mHPEOAoDeSxXDF9MczNwvIUt/ZttduQ2PB5xiXID1Zb6r81xSi3GyrRP+NuYhNwWXoN+KX6zqePt
IfeaQckwFIdUHBKFK0Ee3UkCdRNdea5kQ/NBO91jCBf6rDfcWpcGdnHbCFzMsDWkmL2vGKsPcvb2
hGN40neVnpNrY37yBu0Z1kITBNWAKxFfEhQuQ36PI59431bEZD+CNCio0QD9mWzbZkLtPMDUHOh8
dlS3GYNEaiY7t/WPR//8D8DV33ljGqKFyv4BIZxqscmon2QE/HFUeD7BWtUd2nBr0lsdnbKdi+HJ
yQKt7iWNqFMVT/PDUtdHtSm3MiBexhXpZff/nDm8vvGsElKiG+cpGjvcfJ1SKd0j3TqCiGbMcN4t
zO0IbzMxNzSx9vFY8NihlZuAf/mbpn+Ikyqp8Bhdcp8J2Ke/pncGdgx5Qu1maoLrVmVK3aD/oAIc
HqPu8TtDwuWgtRhA+PKxYwX9XMlwsa8UbmkKn5tcovVoUwfOcuCTofCLpR9mm+fhxZuQqV8Iv206
h3UcnvB951s5MYGZ7Ff1AxN/KVEGk6xOwgvEBhiPcQ05XDbXCBsASHM6GV166T5Ajiu2oG/29tbM
alO3bsaqqqCqNKk8jJyQnwkN+/KrjI4L9SKfAXOa9B5DmYOMPQUqlkVqjgEoInoGL0T/z6eNMkLg
RW33ALyLIbmL1pqvw6gZJWllGDQsE5bkqAtYvJagE5+Bv2WQJdRphTWG/5vou6K6mdTgk4TZSS4r
ddURAc794u+TC7D4K8bv9ovu5yOXQWhavwaLOXoblgVXqiOSl8XOtw1oxXppJGDssDIA6RyvQz+i
5fiCZDZNR8D5IJ6lJbF94Wymu4nSyl7oYbwZNNujnzyap1YZuMzA3Ujc/qFLiDlw8Y/fHmrchsWf
/7BQ0RjivU7Hf33zI1B42n0uAmmSi5bUe9Ai7rTJxL0K9J6QixCROUEWzYN5QH67jsEa0xJUcWfT
dXsHpvl+T14+mHtVhEv6td/Oeqi/TOG+sjaJ7WfIocIfBDWkuqE6zWddqBvQkw+4RcI111GJqlkp
C2d+ZNd565hn123XreYvKjqi6CEkx01xVcgDQ2AJn41n4GS7lydn6HvIKCDkbH3OqQmygIPM21pM
TRywdu0uN0Ggu2CCfzGYPS3EDfmpLq1M2ugL8ioed9IolVE5bNAptG5SsMD1fcQp2y7qSfdXtf2A
Gxper6W6LlhqTRPWXi1IfQvfKtOHX5jsqZG/LGaT6vE6XP7DdkYUtB+Wb4Qse/z8oET/WlzdjGEm
QVStA8eSOb7ZsVwiTA6FpqVaW3fZ//5+PwfDObovxbKTamp8TJjdIM6/ym7GNHuFG0dsa8nJlnek
w7zijYP+4CbdOVwhI8vxeg2pq69FDkWxPWZWh5IfQo/g0+enGhNjNj3ODl4SSzY8fQv8KvmI5hkL
GIJGYTnOiWZu8fb1f7IZd10MGBjYJbCXOnAemfT1G/NckbhqK4hQeAtVn+DPYkOLLh3LsM+ZWLkK
t+Gv4GBtv/34nWmxmGS42RkFbtFukseiJAeM2KBw+GkOW92BwfuE2wyQjH6GnD5ct3rfZUVIkMQD
4WhASSk5KO1pF3SiibxfkVz28IJ0A8FX1e8C7SFRH4TyLWBF6XPCYdUPdtlUKTnEVA/t2D8wwXXp
BAkF7tb7sZAvh9l1qYP5OXm/+KlnTOmFzi63ATaQ7gXu7zrAG4DKDdHQPQ8x8F8G+Wf9bXBqmem7
wcwovQaHI4jJghKrFb4asdHrGcmTQDwcdfzHNVoe1wegp+TgZLB/9b0SdhKeGdZMkbSb/wno0pl5
myHkn69FEGtBqzl+nxWaCOQTRYmG2JKL35QzhBpsK7TWQHO++rVTxS8zeK6sEQ/3vpVFHPPlqITv
eCPhrGu8y8Zmw6akVeK/LnBTmnfN3vumXR/w0nN52SfrJl+oTqJhy9UReLb3+3I0IOYjx7RDuNNP
QBYfDgf1yW1khcuxHS7sBaORHxe7VhKp5CU+mIURo7QljaMENEyhBGrJTqeKV1rJgyvPa7YagIEM
LxOT2N2tc9rfc3q7eoHmeD0rAnG4WzxVnFpvXQ83N5C63fxUkhoksdWP+8RXpyuSuZ5XZ1f7jo1i
JOKGeb92CQr59M8G9pr98LwyEDnxKU6k4l44iVN8mKVlw351H538/XQuxQBeRGL+M3NE1RGT72wg
84aRZOz8wOMpedIawMqjkuiiLcnV0mUw5g6vEhFzOt1AVIzP1uxDK7vmKvXoU+YUqymeDTKlYa6y
HKCKf73unnANR4rhRsFIo2dS4n6IhdrW0yxmLZ0BeC1O98zG5VHP0DUsmoMckU2F3MmL+y9IsZk5
ClHU0HaoBj8G5DbGq1PFCXsw8vdRnDBbuWiAYC/NmjZVgdEWPAkgwoFalmBLz3GnRrq46ihNcPFl
ObmblnPKZVZVxZXo5Ns/pYomH32zueNmLxB1zYbmmEWuERieUL4ZrXgZDxUiFPMtAJJ6j5ZH14Ap
ax1uc6NoIR9SdZU/eC3Elrt5ypVGdEwGpSUIdS5JjOQqD8cZBQ6eW6HpB4PlTHlBX0YfVgMz8Ar1
3/2Mai6NQOZ/t7nJNC0uBEZTpXeT5W9pkfR/B+yqg/l/PLIa+K4O60qGrOLAxB/83ekyn3dK88oC
TybrNZvZ9soNi0pD4tePfo7nNNuLSiStA/yr0l44CVxMHMRjq+AUaEFORjSWiYbLucWukffbbeEt
yP/4tNLxfE9JXe7L3pw7vfCCUbrUfAl+KyHVvqAFNGq9TUhTdQXCg52vw0abpijD/ZQqez5+Ss8X
6e8TchHdDpTzSycAXpXmuFyRObI4qbGNVA4lErIOUNP/c6PRARXHWIBy3UZL907cu2G+V4pvpL/H
L9KUiUQtggQ4LLQgeyAS+6mO9lLNvwnUtGSbbCBWWxpOvVcc6rjVQJCLUuTIXUuAoko563cmPM4J
2oOf3bCVDj/M7bIs0doBRmCXaErYPtm2P1fQzJ85bc6EnPQAQrDm9D21ECM+KAqfwOqjhkXRge+g
GKlRdeIodi6IvUa/pKDloKNhfkciL6HWSj4ryDzrRps++9t3FLPIS+QWSyW9ZJ3zsiJv1PbTFwOC
m6WkyrAz6iZNhQr3vLfBElktk/zOgpnZNjsc5EqrLa4YnNS5zX8Nf2J1xB89UNCh1DJDt/X6TkUJ
UYRoyUwQkiZNA1FOov94uQf/xp+qjq7Z9C9OnDwSuqSs4yJEUI7Ba1YDje5uk4V4LI1/QGBfJsuD
IX+G8e7BFouNCIJP2Qknr6BjGoHbHSVcZU3hvjQxFfKqRf+JZ53LxDpkBxgQd4w/0kayCEfDmms+
lg1aFYf5FFI10+mRKoGlfn6GIx5o2LN2d/lN5mH4TpvBi06Jl+8Y8ndTPGzZlWXlKbyODKGDQVGA
YU8bwT59qAQmkgrGwg4gO+/jwuDL4u/j+eZfvJE0XNPY5ef+w8T/y+BSbatwJSDFTLOW9fPR5rdD
c8I7o4yp6R66PeAUAkeA0XkByfYqPo0Pm7AO3Bf9IEa7HCHQPv9Fr3SX7Yl5YY3lYA84+1gw/PJ7
dDCiIucpOStiam82yyvWwOCQdap1wxDXCG3rI7Uc27WbQybFl5zOg2s87D4RJAp0bvIYw6s5rwuF
qgn8NyLfqcPE0/Bwcwe9OkdKVq0K4W8D8B3hCl7RR6kqMHFFREs+EFdDjASq4z/imSZGGwDE1Swk
/Yw8ngoH058bCba7vyj1W4lQgJyorEhaV+3RiC5CZrDKHM4KCWzS/9R+8x2xGiy3UYHg+8rJRQg9
SWgMuF82PUsEYvx8YciTYE2ised4/ko1DJSL3CYQAyx6wd+vO2iFc3h+8n8v7JzrBxAtRkHAQVSR
vL+NMfQ5R54MyzVaB7n5Rby3pfL+hfBuwZdEI5CnEwig+Bv/T40HNSpwoTt2RMF8Z1zXKFfCjEtE
uae5BTq66gbTlFsctEU0s/E0gaJ/Yy6rS4DZqN1Z6LXsMoKmk2GpnLgw8YBDgCPvVkCYoYqzSMIs
eUjoRJs9i0zZaUpX7kGlYKzXXqe981TVAt9rqWoL1JagoFePU8l0jNp1PgZeeGhO0/uRn55goQhv
XmkrryT0XYrELy44PhRNpdeDsO1am2HrHLqO2pjQG4vJtHZac5qkRxyl7CZc5mm+kMmsww/MWHIr
3am5Wbsu0+BhIwb1g4O+rBD6hyfbrWN+57AznootPIu8oVrep4s+GPIcU6UUjkNytYdhfVHOlSHd
y8f9wTg+focwduA/9g5pUIC4u3zYE3HJC+HY8Sh5C8AfAQWNDfI7hJhPNIcN2jLbFB1SHu6vu424
zHHD7CeoUEJ8kcqCPD3LVy4b2oRw6P04m4iuiUVHgYUI3amrv1aZMHQSiR20yNJubQLWSvr015lU
5WvglXkGdiHQTP4zie62dlZp5WbNQh4qXAlbn5uXDS3km/Vs+/FSuhhKZHrphsEfMaCtM2Wei4A9
wyyr3LN0O90pG9FxnrKODgcWjmr7IEXDgih5tBWG1Xd9suWq4XxmjilL3AjaiEjarLvhasGLhNK+
5mTwBvhlsUN57jH1p8HXRwnb911yp+Tbdec2IBw6tXkKddkhsHKnbQ1DikAReFSMpvBAx8CoZSST
vjbAZxNd3GdVwFr4KzqXbl47UwKM3cqFX77A8jas1MNOOEg6WtoJoQF6bnN/8HlyLCtGMviwhmm5
Sf8GE7EMLTpdLACVRk/H0z52a/69Dy2mny8kJPPiljwJC87mhwOWcv+l52uKbLKR8qMSt7+pJQtJ
gRSHsL8NUQ3OIR1bs3WgOO2czYvH1qLDDzUprjQOlfqLro5UFShxThVxgOXcucsY5xhIFCASL7v2
uWc70B9tg8Goas/rsVBfc7Z9pxiHco8uwJIaG/dF00+tB2uZWtkMInQMpz3a1mnJPWfYsvXeYZ8v
B6jSjgL1fmiw4EpLR1JuOQP/PzepOprln/zqj1rUoUw5Z/7jCdSwJ5cNIygVQof4eSDQF26LXNkq
M6mTpRpuHOlY3aiedKDfa9YhDsX1Sc2GY6/R+6yFsE8po1Jss8EBKZGqTtNhtB2rfVdFbSsXQM0/
TfENe7SIj6byb5QPw0NXNr9iBKvHU+v//dDaXZYH/Je09Q4jQoiy8bm9Lr2njzwXGbdacabzLAFh
Q7gf9CPMcLTebywyjxcYc/J+QJg2uqLWbwjreF4h5ew8MiieGv3vVynk7uoyrFj9PWt6JUhnRJYO
TC1fJFh6904qX4Tg0h4p6gmXJQ91K6TzGb7Lg/px6JscLmKdJQCmj//0a5o7FB68NTjNs6KJUgqe
7esVlmXLoBSNYVkVyb8yf3dYv/RduiI2GqQdh6ydmoDo7WnJO8i4I0t01BCQqDtG8/9ce5RfU+YV
krPOoHTfL88WhQa9P/n8CcSuzj2Ya1ltmjSSv/unhE9sZBKFymItiKBPWEiVwMW9vmRh3i2jnjzZ
S6UohNqIrzWbFTo18oqENbNmEOc/u1t2z9MOTsbMq/5qNrwIa5o6kWtakgd8Els0fH9akKaIJyuu
jz5rIvPU4LqAqnokAshhU3Q2lJE/92HkvdxxwHRPIqhXkrxWruxHROxhMVWAIT9sT4rbC43lSUlh
mmkEnia0rbr89sIn8/AW8O6EVNSl1cxqlRJYdWixbGODBwQH0Xp2TnA5CzE3UKm+3QFEtEqmsixx
/sRTLdTybjcSqXpZadPwggXekwQfI9/pcf49sjurxHarcUKwlYM8cov/SaPC0iXWEJplhoPprx5Q
UjKO884N4XzWvyKwBG04FO97HZhJ70GIhiP9an/jXnSWgaT73SBKMj68uqsLe9dx+XWrRrnFlI8y
XcyytftySJd1H6qfd0rswFzA5afJiRrWj+g2QHu10zAEqhxOlFeOxzz1mLWppaq7kK75rtmu6iJ/
D5B0cDzMBrk5eOVf0KM4YaDXhZcrfMTmPtwom1ovhglUqgwcuKtZ/3lpDbkrrNwrD0sPRvqyLvzM
G+W2uRA9Uxk0h2Rtd52aH4sAoRIU/fPqv+6+QFWe0UUnUrGNo5Z3tYDf+RAiqmbRRIIUrpdrz98a
0D+niPEjUcmHaxARF+yyrlZHXn6A4wdrqyq6bmZgnEkrt5PTdeTNdKvd4p2tE45PL4Lx9K5HazKf
ZfQ8zXlBqnuoJ1HPEdcquDbaloLMu7hEkvbHjHwFWypC2SKnUwesZ1M+FrCu/7WKB6qOmmhJc8Xa
ZPspIFJAnY24DW3uJpOkxAnPAMXAmmwXcLzB0uKSxJu81IzkXqmQvOtEU97tnsng7yxst2BxM9pl
tT0LuER16tIGbHGsBELZDuYhFJvD72qK/IhDsfd93miJqzQzOua9ghL5efV2nox2AUwsAo2Zrxnf
gJU0d+vA4iS5y4WZznV842pfQSKXDT2H5+GcNH80nhEf6ZJ1OQ2b8LZwNAvALYrDbwY7LmJVESQQ
tWXvvRe8e95zEF5UYS9xwiYiHZe1IluoyTzqKEgeawWlhShSWfXlIXcLe2qSoaiUTxowZZK224G7
APfGFhoGtu0aNGoNPkgxzFVBJ/CEurjUKzdoquOSKgEQrw0sTTS6bcmSFi0WeSUHsjpnDEfL01qd
vE4g804EvPuWf8DGAQpBX711GwiOp7hclmOghjNDlN0R0hA+eENCFqK5Kvc118BeTfsmQHfGrIy6
18rgqx6ptEwczVaZZFHlOc27ep5ualFfNwWZUIohs7YDD98hLf45WjkEld76716H+75+YLhhdcmH
7S3CRHTFozUX4SU8AxT6sMef+1PYNg+WGw1bemxO2I89OaySyZ7oOhEsbMBIofEuR2IsFZfAWRT8
HIE83nVdI1BiZ3upheL1BWb4tgM8LUQCCgjlXBCJkqfv1A1U+QtCQSYPMuv0fBzZ0lH4j3xlEaoh
RGMqcUYi3BdQ1F33d6DwsA+A9Aq59Y+mh6csZnfh9R+IadqLGnlicadwT+pRuziygCc1DiQCwsn5
fUfYYfvBbKzpdCqGqEuRrjOz5bv/0CLA9lMkjqhGjYeD4TTtrUftEALkCYk7r3Qcc+yABd0utr+m
m1ZNgX1YNrBpOe22DpRyRY9RYXj4rnrc9DTIlEDy07/VbTeBuxRPewXcdR2QN8BlJBiZNo30VxGU
OUIixIIr7z1Z8m9UWxmffSoo9EqI/uOUq0q5cssSxtUoWmN/R4hhtgHemqNsqAe++hSa8HGtcUKK
bE4uRoRjHbUN87/XSJaLs65oyU97FFC12/zUW9OyVEvTs4DXiprenboyzYAIvZZEtGUSQa6hf31K
twGAqjMnOVNddyoSQjTMLTvfqQfp1dUu3wfqoB4RkdFyRqO4qbo/M5F7D2OYi2GM/HEKL+pL0cyJ
DSxIFz/3QXGqQg0EOZXm93ezReOKV0YnGYN6y3LjsRWaZy28o0r98/33AUe+cLXWJPp5R3BLCtEn
Jqm1cz46lhBT8kmXRbgCkcSoBA/XoMoGcvvwV8rSIHtHCegx5oefh4e/Iu+gp0hBgbXzqE3VeEMk
yLsNou/qYZV5eHJVnofSRWazoen0UP1sKwd1OQE0gL+Ow5f1WwaSibrr0wFSWw1/CgmMXJnAcQJH
9VwoR3FkvIVmWvIcsHxn8G+5X3oRDzzRHl1NRDkSGmS1iZLpBGc4xZbcRglbrGasSnbgEHqI8nL2
CHYFDhrbcW/hFx+WLRbQcmKRFW0HPQlBLSsPB5ZbQRm7ED8kA1IyXY9flZN1QxlNmMXMxEGPDMLN
4IyZeKzmHC1WpbKnPAkAnKHeMUyPgHcDdmWYLP6hDHBz5DQbbpq5ls3jNhNyPZMj4l3neGp5UgCw
4gZQdI+ej2gFJsbcMM5xeoy6JfSnnesDBPe91hZVjpBIdKHlzOvPEQEtRctV8EnIZcRwpEwFxGJ3
HFd3GezxMO3ON4anYcMcMfQl5X5Wwiwd6qT54+Ux8l3JITHTLD/euqqf4gq0Z2vhZAcnN0sdxmUi
CRuo8CCBI2A6qlX+llo/4ekJ56R8qW6xGbtMsTtrjx1XHBgcscFYF7ziF79BNAknOTvAu5y/gwXC
6bdCmfUvOz/V9YDdEgZ43Y+9Vs/z02ZF/+W5dq7x0EzdXK4OgfOCbBWTS69iy5ags9DwxpCT+/tb
oVSMbOONHfX9Jnm1MBKdY2xrR8R4tCPPXQhkmFtN9NITgC3X4jlCHngaBH+ts86Ec4n6z+pBKeaI
ryvDHntM+5vVRj4K5l0cxuZUhUkxNpnVcyFl15sQ9XXJ+1rSNbmfSo1DlrfizRaIb9yuyWfzqJxb
bzNmBno0zSXvZD0zjHhpbBbFwsqgJ7WW5bklPd22T8c93DVEAtw0lx69qGSFn3KoEEwqwWdIs4y2
izMANqI9hzOP3HuMmb51H+PJCMDWo2umtyrAXJ3f9USab136wBqCb0+8gBO+MEQJjJd5IjVRQGhU
9sgW2YrJCn+164MVt/I2gCJHfFhxk8KL5sgmtDYyc6bZGZ2u/vQUpgds3NfZN0dnpEepFrnrBSsf
P51kuQQKeVn1pUYu7AQC/l1nT5X6qRRlHRcnX+M9P5lViM9lYTOXO6rfMCwaF3mwYhK81wovcoWK
2twqoj8enjw1YeTAXeuBNjptR0Ri46WYTWrMi0fCjmXhNeBWmJCVt5wv0pCR0WnrGqLO5+kq4I53
fa7tAy9O6AoxyLIJEal1u476S9CyNu63C0DlS42f5udEjj5Rc4/DtM80aF4VZ38NcmD9ZmRwI75c
+kPDiOWZWhxYTJlnBWF0tGDyjrnz2MaXuWgeTWmE2L+mFEGZIedio2BnhGdgT6R9GqNmkywhOkvp
Bp7IB83RPWOsjvPM2N2K9gg0mLhaWffnDzfRra+WnS9uc8LzK9usbvXL26VGvew9JlvIln7TlP3q
5UX117PGDM90AgWf3IcsyxjMy5gc0xUt7hZSyUYn2gxBeQEu62cAWOYkwOt7sF3pA5Wg0RdgEfhD
basxhuQPA7IlnOB4zekaGKO7t9N75jV2UjFsFinyz9KACsWyStGgZ5e4bLFpPPoClaBLPH9tSURI
D9tgjc5FyANbzkzf4zoyztlfFsA5HFizfUV3hQgyReb4Y5iJpMRkwnzxjFHwnAI6mZWbmBcUhYW/
KSNiSVh3svRHmb74u1yyleT+n30xdFSYBzdIHV52ssstEH7zae8W8Fn/jYjJNT7q+mlJ9IeCW6u8
Yk450znEFMTTtwUaCHWJ1eu/AOqkag0A2BLB5LRVHhKA6CPcueOCB0Ac4RxdPbdyaw7DW+JaLrRY
HdWV9YTxbgT3QZMU9s1mPWmLhUH4i02Ild+kPps4qOHE5UtwYv7JjN0Xq2/WlVqlqHhB1bHwYnNx
FCoAAPAxms1Axg9NwYtVZXYlWWjf4vN5xWJ3KnnmzpXlcDA+g8LGSAmBFixw0sMMZzVUOjSqwArd
sdqS0h9p9VPcNrMs3Mj3XMgYV7oE7B2DCWKkcGHKO8j+xGHFHOluODzTkzwBqNuRL0FW1yB1hr0v
9x3b8VrPiv15SkpaD/9mY8JgxFw21YPCumJ9SxouexDGW5BNkUn+TvjQyyweF7ffnanqXHfnzL1t
kClj/a73duQvpC0UCtIm45F78qmhEH27+XyB1QJuAGMNDeJPN41uA+bFCd5Kq2hx4f83UmLxsZK7
MN8+vJel6+8lLsMSKQ2usBx46X8+USrLJV9/5e92RdIOV0z6kAiswNeesdqOnJ6xDI2dsVB8tNIg
5Ai6WxlGkK63vAaaeQV9oNCja4mGU2T2R6brru50LbE7z8eUrj17NKziwmbuJucM5Bja/NOD6Cop
JYR0An6kJ89jx7hhCW0zzGYF3GSOWpUIvyPOFcyZYtHiRZyC5+ObHRqiK0HqgTSidx0iOGuj2Pa2
sbZXwWR2sqtdlYLyzBVNge796bfJtB+Mxg5miTVekfriW43IkDyYV2dWDlXcTWwAbQyv8Zrvqf/M
8Un/i8JdArORU6Wy1rGjxOzqKPaff4a0uPPdAQu6PjdnzLCq/o6Wqv0CN447ysSwgGGFOLutTgLk
pX4Pm3VwihcTiJIpod5g/jN0DvAFXiwa8MoEgz0F1VdebSlrLl8xKXKlREV6kT26raKfbP4tLbT1
f5cGeeHbCnujz6vbqyoUB1e7kJ8qtKMH49TsHNkT4cNI3244uWsaZM9UQFyGLPcj+SFz4FX7XIGS
6j4oouP7GIftP1PkWYpMursqxRwmM4SLhSBODbvw+zKaAjpscgflWqVw1KRaONA1LgQN7ekVw3sw
7X6bjckPTR/76aEizgaB3Kn5SLlxg0gZyGcxca32sIpXSn3ZZgScVCdwgWdWe9dUKuAH3x1zkksJ
h9Et853I7w00KgRUEIYLLnjsbIR8Xb7ZM1DJSoewja+UOmmuIfzb6XILfKCie3oVpyNsW3lu1vyr
WElUn92VBzevBeQrQFHse1AfIvIdNB82FACxt/zjeB2XTeo/tjRoXbYnj2Mk5pjmUPoxHec4VfAk
Z6eSaK5AkfEa/MdvXmjd5SETmHUdoeFu8JC7W3wKLfd3NcyKcaDEDRxl0AMXhrq9bzZrclKsw8yI
pGLWhQU4kr3ZGibIqAHf9PSYXXX3yKZc3azJPovvKBpajkr6GQ2WfqHcKSTHbW/pwbk//zJyJIF5
RjZ9lUuId4gWRjjbok4F1D4y6OJsJ7yG+ApaJGnbjNK0rw7Q/jB7539twydBuOdyo+CMSlH4t+6C
8OzGnO5OpjeFb+NNCC6pYTEKu1AfWB1SZ2fS3sb7VHqYhDwvTefx6rqZDlx8biTZi5s2kU62YQZw
dwzAsgBORO486AoAShcSverrrntZfqluoMCankZCxvuagzq3OzrVD8ASZFZ1805b8cXEWPkR3VbG
c5a6/QxeSH6XtBnOxLQjrSCeTqO3krd6t/wQdXw6zneoCqL1HWgtklLgj79U6BkeS81GG3dE2JL6
ct9CsOhuE6Ahqtf+CpxpvFaA5WdJHf+a/pBFS/VOFrdYvcPLvKZofvjV5T3u+Kr1VbS+ZlbGrwdG
+BWXnd32EDjPx7IGLoJLDEjbqVsKNpX3W8YjNMOthX8EEYDNTB7LfmkQnSVX8mcRSW8ZCVR74OSP
v/ukCFw8qmuQuzA4hfP5TXaxF46qjmAQY0nbbtAIDQQgD1aQbHDAbjBac1qO0XrW8D9ZaQO7tJ6N
jq0+Y6xj8En63cMajsgBvuGgq2BlAdQXIh/qL98ysMROeTMVm3ZUzlT+np+5XS+wW583JRXhQiFA
ScHYt5ekpbrcz+6z2wiKdQNbUMoyju3FlZq8I1+J3U0MGTqwFQnIpF089uqFd0YiCfaqV0YWQIbh
L29V8+6Nh2FeVirqecSJgWNcmZs1ODotYMqtAQobdt/T/vsgWZ8iEty/7vblgFFVjmYt+q9YFoIB
PObuMP6BWq0VqRYbLyHJS967+CN0RbR9tgkKEPglQOrLl97cISYNTdZkPpgM0ulQlR8eeNQ259KK
EKR921apStD+gyrqdFkLPvyaj+MUb8xbLBi736OG5o/9gBGJ40FpAy3FXCWHDgy0nIMHL6gOA6F2
ign2FDrnz25bC5fjI0AkZeJ4/loL4KO/JOl6Ql0zqdIQ6e6IJwLqNqnagRoVyaMCeWqt0nV6oPCw
A7qX/kkuaDMQ+ddyBnfx8E1OgcrMMzy0uT/IHb9hbTp5QN9vnI8YuOyaqko8xdNnpN9U1o+CBe+7
jdBNm41Joa61EhEOlA2z8tWvR+s3eXc0UEtFB2nUs42xpf1HzlNWSdAHGWyIqAS1QVxiWM5cqLrt
M6z/ZAj6gM9XtAt4cOTGsQ5J4l5bivGoDDTzp6NS7EXabg6JSip6rPqaDuyo81gBxV1mRc85Xvnx
RHNW1cOCJbVIP27utBMTwj7uOzzfvNDGqk04/oiBjQyVJwjr9HWOJmnQ9cDNrive5QRwLIA2oY4b
LzFqkEh4h31/mtyAUmA2bdEczJOyMMkejpL5Www950r1uzC35Zj1Z+YARFJDcDJh+ouxP4mUP4Xf
inxL8lysjjA8UX0HNsNCQcrnIgrP9QBCx8UZ8xt9KNwPZGj0mgotvpMpWVfi/BanNcgsFS4Rrn1k
o8d2PgrDKrbxGD+mIoaWzLqpk0DOtP9eYyTkA6CRtnmPzfpIIDlmhL62piIqQTd3BK1wnPJgrNGV
63Pw+6IvVWgi2BZOJOHPr1O81QTGwrvpwNRUgQ5qsANLdsAOomAGxRmnrslsCeaLno7F9tJ7woXY
bq0VXPGEKrOD7YvMUjTKo+Rx4EnSTniuWyWRWn7TnroBOOo3wQ3y73spJibBi0ZGCiXG4uQOX67Q
bumUdt5TlYfaNsbltCm34uqlxHaAdBCnC7ae9+A3Y+lK6349W6NYfT53nLFClB+1+e43DRFvbVIq
vfM0UmOTq0w3XTXf9bMELvmLblYvlnpxuoGhjWJinxZNIDwFVziU12uNfDHSwfvvA8KkSknjBRVk
iItr/Hke4xmb76xb+TxaozpTY/W/wvnG79+ggM6XIR8Fv/n16YFjC3s/CWCvfYAACuqul0h+h9CU
rz/iIPgYcc1B9TMKZGj4OTu1E+Tm7dnKwka4pUa7C5maYJIOWExdaG5BEwzdxNJZIP2mYoMLZwS3
46E1NBY/6FKovTFOejPoT35OuSaQxKT5lhkduk/fzei3ynsfKU32QpYG8oqxQuuEX/JKzNCFPfbb
jFBFwPQ5Wl2EnxMx13WoDnxhf2N0L43XLzATKo1xQtLigeiLWgvZ+Af+Tl0Svr6kLznT+tkmC/8I
AR9NX2wRDX6EwAE7jr+W6nlad2JlDBtQa+mKPUTVYYA1mBSgvsu3EgHVeNksnLOAMCcymhNieTib
fle0trxzL0vS+il4SCAJ47mcZ4i+iNL6GbqJ7rst1YHWq+dIQ2WDjF1brj7OjCuWFIxGRzklsUbP
Y6UYOPFMdOYyd7sXsJtI7bnTjuvXwdtua0rX8c7JjwtDMmRWRMQbbirHi4T9ZLYUVV/NxyVhkEZ/
b6o1VLSdUbqDnj5uMNaoDZTHNrOBFPvTqWlN8JWcohUOq4Tz7i1ku6TVCioe19fesV5vVr4adYHA
DQQtxQ0xr91UznZ3PMC6+KE0DUbflgOMiHbm25SiZwnWy/LCE8lC1v9UnlTjrkmsQrugbMWllwzk
YdXbQajKwYnuuxaraoNNBfVFVURhOve7teuw/5LAfdFuNDcbELsu1r1Dtnyeg8cDbsMsV2usWV7R
bKm13r4RPTsYU1fB5tLaoBiH9mLNIJcjHENq8aEv7ObVGn8DfMXtXCTloqqxq/WxFwPtf8AOOk5+
R50EGKRr67LISIGLEfkTnpYBg9LLcY/1h5bA+unq0kD0bu3Co1aYKJMUHJSu47KI7uyMVMj2s9PX
hV5L6O67uDwWHk8q0LmwFqf9Mx5rxxsk/5kWZV+xZ61rhk1S5Er8sX0Va7hN7f6KgmPN0jR2EvET
Udl8dYnxM4UyFq1+TQZ1Y70HH6ebMv2/jhLEYYTgQOaY2HrH16D433SLnHQh/s9fJKibzxFgeEBI
fNW0Q8+zqK25m2W5U9hzVV/mZv4mU0pAtd5W3wJ8XckKtI8Q/sHOg8Y/VKn6+XLjLfa7J7Tw2CFU
Mw0SWzgMHaCkv/YQmkJBOy1RY+tV7GreCIT2PMARs+kqvcddDj0XDHgJRXuOjSbllIlSMQ7mci7+
hbdK4NN4ZCDFW1e4Eu0emfG/MkF8NJXjEVts5+3KyqrV5OYZltHxFy/KPmSGCqVJwGekg64aVPuk
NsPr4z+2uh7nS/zttktl3i4J31ytthc5rBiOTPM/DOD6nqsxkxXzfvBjw2lnsB58t0oKAfO7yKfW
F64Z7CwXW7AmOvCZE1AwS86QSiF8pckF+6H4bw81eVGQh6JqqsZVexMWkICee2D2mqTNBMVQfbZ5
qmRzMZkBShk8y8V/OGIj8xmT2MvuFDwU1WFZg4hZn8Y1LB0g5u8CPu94rA/3t4p2xds4cap/nvV0
vV4b0me2prztJOfJVuJx38UNn2D3hKqZG3N18i+dn4rbmnb4YNURTcntaNsqvAcFKn7GeZtiF4Kg
7hzAFqC3LrMe8xHkDDr3iYrD8kHTwVxQLjuuhBKmy/C854O9VpNgp77Vme6+o0heDXCPqgw5Wurw
my/b0mVMJyTk/ytttxe/JKdqViLc0uczHVvcQeYydu/eJ4lXpxSOd+hnZpRRv2ly64U/gtDGxhsQ
MPiiB5wQWN8xJ2n0AAPwNhcmlqMF4aFiUVeCwJMht71z46Ce+ar13eE4BBT7aw5I8fUqHEMw4aYd
+5cuPIponS7b0g2EflK3kLtLvxA9PptQEhLW+m3YQjxcINn7h2aTeatgtP+8de6GIZFzWhpL+vNP
ellnUldgk7ZTzECHhzdReRgUW1jBEjHoZXH30k3KM75ihgY4B/rKsQTySbi4njSANHs6p7mxK6OQ
szyXiyHqIKo81V+sKhSG0vicOJfLn8Y+/7oJwyYGnGF5AI+skRS61EnAeQ1Ze5GVmWWzoT+rsF0R
3i8Sp8afYz1P86bg8uj4himyjPJxpJIGhrPo9Q4MqNeXdB6QcAmu5xRVN23MVp3u5XsUFOo4OioB
pnfXD7N/pbdsYe/NzyO9Eqo7yo1r6JZLV9mb9GA2bLGZMvDM5/Rnx4mdwvzrbpqqb5SGtg5Yu5c7
shfDCNixJvkh+mDl21FJztDyvgDHL7RC/JyLce/hvCFHPiO4iVqERZzan0OT0Qi7hR0hySAsxWTE
OsxYKES+hYpTalSv670zJqauUn6vzstgt1n9GdR7jsRuLA4JOuP4Ivw3dVKT0+lXZD7GmNgAmgoB
8o0H0oq0VSuzx0a98A7OZI7jwkbPwsUmnqVdBgZTs124SLx5LQ8JFt2XkCqYqGDJt5uD5iud0EvD
3/91BjRWJlnhY7BlihGoH1tco46ptXrrU5GtQhtG2zvgzq2vAvJ9A1OpLsSJYGoqcux1YFC7Bo3Y
BcspRZZWZW+4imHnXAxEMDVuR8KYKa0nsXCly0IzPeUTo0R3t9j54q+3MmdVUpWf/PlGe/4FcvY9
SzoUyVq5rhrlZpCF95Pn3//ehil7FPjr7riw/wEJBptOUMWpHgUPQHTCQkQjSDRIFE3fqJjBI53K
Nh4hFjhYtJHvi/wf3vTTt3CgHD8Uqim2H2ot8iv9P5SHn3d7lVa09XFBqhu+1YWai5+LfL07cjTY
S8E51N136g/RIUd8xvHIPLnNkay59IKFD2tmR8Hk4jJbdaWvgkeGKD5fVjTL6PAdNSyBlG9GOxYs
G/jy5/xYi1TuzZqEwnufLOTSkechzIdJnXgtHfJJqS84LveCIRpEuDezmPGCZB0VLZqS+ztyu9Mc
hKticA85ET6pPpLn6bVqWi8EknSSbMUMcvHa8p0Kr2AHOriany8fpIMmcBR7XnlG4Qd5fbP1Lc5d
cjfnJGOAqkMBo/8n89OLa+appQXcktLYtp7eWW6Nk83MzDffBOism14m2uHhf6OCh/cAN2x4EXKm
tRj0/5q6LJ+8hhcNEUIPdPq5IbYZ0WFpQL9CxyZk9XNKA4uW96mYN9i8crB+syF3Tqxrp3nKwY9G
1HPuwaiZsAAqycr96zKSwPWERI1fd5g4rdKVtOmbIt7/Cj7rEY9+I5O2fZdAo77ESub+s1CWnjUu
Z4z1puiXxt7wnNZUGosEtdqFwEIhgKvXIVJMNGR1HfAaxXLBhIOb5JyJRPMXJX5x603eZymkLBye
EFb+aS3u9DOk/NWnQzBWAH70YVg4JnprQBf44j9tcg0R/PN1AXiEN2wsp0cK3yby/zdjnwb7CZUM
FvoBsMPTStpTrg9K1rzJGOkbqfvWyq1HXwe+XoC3hgbCg9J381kevWaFy5G3FGmS03yxqtTBjS1n
0j8q8WLK5n1/0Oo6DFRCg0VvQcVjp60wY+gaNCYpH7kzXa8jsiqqgCJaityZVpi0Q4VEsXvbn4/w
WOFjxCLq7RiYm29C13S26tFwxrGVVr63Gs2kag/eapeM1B4Z+199lyerp9kbCqZFxPdSMG+egRi5
qZdSIhYnqMPwkbAOrwBO/zG7HB4iXYK2XPCmuVxTuSp9123uNBT7IPxa/HymSJlmgdFliFS1+E9u
nynvHkIAi1P0i+QuXexBFebODJwHtIlOUNv108Col4doWMUBKqtLtjyoSNAEOPzE7NrxcZpSOvC+
vElNPBI7fqvkDSVhyzQjXO+841l9LbNaxs7KdAUdk6LxVZYOXZvFB5Cm+6X4qimUqTwgRlL3Ad5A
qKHall84wYsqIdrl/X1gdBwR36VQF3NlhbvOLbGiY5rMmuMoSMCTNsUG2LlAH1scP3m0zw5rftE1
8c3P2mY5Y7n3VX/C7F3aGSPd4E4E68rQkrW5el9KynF0pCZzvaFyxR/AN12pY6tfFoD4A2JgHq1o
SPBTXPgxYpgsIvOVxb227cHU8n70fZfGaAd/bBXi6tKEawI0m27frwpqtkkHW4MbcL7hiHnm9+J/
2YpCs5aGOLg2TkJVYqBvSvhwufjmmK0RP/3oeSo7vGq+OdVFWdctu+nu4WjCrmKUGLvIr6H3wfgS
gk/atfngIU7qqqIPkI41J/jQEVG/pMLXCg531XVWhQwb3ka/GYrpGAZ+Xfi+E4b6vHxWEwhplzMx
3wze+EOzhKv+Pwq5F8A9Mr3lXm3k/LG2iW1EUyuE9w0eAvxgx6YVq1/LtbLKO72sFNy2jlY4diAE
fqKPGPCg/B04lRA9ksqatAXAdAN8uADQvQ/Z5R5+2n9ClBdgYRPHj4ZWYKBvX2S3P+rjlhTMYPa5
1b0z6zyxD1KQ7p4LMzXFkFtP733P2cjG6CiYx8FGou5AwHdV1TSbxxpjE7SdAukJBsbpi/pabkll
MLQ+IBldzEPral/eVoJugu33lW2KpT8RGEu8DqeicCGxJ5hUDdmNmstUldLvAdpy1yOoztPHLWcm
IYXx5aTGSXJrUDqER/rVnGE215kYB/PuRdQbL4Os8DivfRU6MS39i6BVePbgCEE6I2T9zHE0c23C
98/0JQ4WU7Suaz0S7iDyhoz3hA1tM0Gsym3xEyTZAJFnGdCNmoA/y5/GFnSgMdZi78xv3YqABqOT
dJoUYkhHI9bc30x9+8j+eKlty8CUDbBhXp+vh/joY7efuTYZFkuL14BG/DlzlARSAwZcrVsmklZr
lFiH69r6DrK5GI6TjioaohM/Wb9MZV8cW1T/0WNdE3QR3QvzwpTyo8kYRc3wrWcYpHMANph+YUGl
LJG/1+20ezOV7rFIFmYu545jnLVAux759FUTNuhqJp1yDEcTh6Senc9g39z3b28gK2gdoVaR/Lk1
f0ajCKjmX7ARgm4DQCdbPsS+9vUsEcjzKtuf/4fjEQOgiUByh9UMF6P6V0GPXMIDPjHjXzvOETja
pOjuTSVto+6Zl5ZMWLlIw0HsiGgSnSCc1agj6PXibpTqCdBl6XJexFNe1bxeESRHuy1aoIGdJral
eAn9an/K61DOEzpso+LBs2/8AAakYHtZXV9pM58M5JuDRA7n7udX7zopLKvdjc6sE0592UkvJ2UZ
v/com20DzoqgZVFXoq3sxVYdhaukFpM9NWJ93nh9HLy3Me1+5nOhR6NIr/g4g3UJ+9PB08WI9gY9
x2TAnbvheJhF+AUdU1bLptCTa38WGHrr86k+OcxvfSbEDOYpTg4zOeiZWyEUQFvzFo6QcyTb203z
N9w4AOEOaydjuSfiUs2BIYxgeSChLsGzTVaHjhm5v11QsFNoreC9+NmU7Q3NkzmZK9cDcOyjoreP
dvR8mUomSPofZxf4fDyw2ljfMC5Ki3ItVBxu5liLTqpldsCiMT77TSwnk4t4AW4//ODM5Wl6glYh
sFBC5FED/Aded//4YvR5reFwBXvZRBTMbTPphuGOweJfUOzdCc3+0sY+a2TX97lID6wOZ7x1Ef56
m00GBc+nL0eF+9zRAv9AeiGKNCaD2yPWooGYJanMZxnoYJj5EzPuydhBR4DAcPjRnkGPFW3Iz63D
uveCyGWjjm9BlB+FmEfVJdlQoNHnDiBAiGMYSddDvmvdz59SIvZLeGUEA5OkaA2YaikAzZfPz3H4
6NnkdNfDWTV9Q99/M81rMQuHSLgjKTBWRtj21EbfpA5ebsLN9kMU9s7VLaDa7/iD+zzlLXljSGuC
rv9I5Fxpxi0A9wFiLpzBUQF57wQAqt9IkPMiRsSEYx+4BQ2fnxcU0GffbbRNjPol/5VykPcl++7L
KRcAiJ9ydpOfE2gH9A+GzBE+1KIstjhYVXEzig/Fb2y0S64uAhwwJgdkOzMrMMCWJbGoVF4F1egy
US1lctpBJegtFzRfBOlm2RrzPufRPHQ6NsHioYDPNGP68mygf/Y1f1gYaPq51r3ldetj5oTHYzBO
ZnMtP8IC5wLw/DtZ86zERMT7IFjIA8FCwqEVdH9XiR0flWpsTQZpsvCe77QbUArABbVSQKOCyDXR
SU+WF3+bUalT5rOGAGYvuBx3YsY9TExLKPHI+B2sPCWyIrdFg4pZV+cElsXHDQ74vDXkGzqrdjlk
1ctQrTJ9dUBl0K7Io+hVc5D0FoREP6bJynkxVOMNIbeT0JbZ24wUw/JwEAmTptw69TwdWSfbTAxr
USm2PWneVYpUQmR1v/8cA2hWDh3F/o180hqwufYAGTDtRMI+iGSttUcZzYUVwF7TRKKeah8DatRD
ctBWfQpJul7ZYpVHJnK/V0YncpQbd1JLFQdZCfMkutRLmEfrSEIfVPqHyEOwB3LRP2hQ3MG4kbPm
/wuVS2fiwTNUJPViA6BpbZW84EfVBtZI16VMj5fRvQDkjQEQNIsI2v+NwofmQsaDx5nvPipov1H8
/GifE2lou+0bwHe9P5PKTzULAjG+TTq/CU2NkFbPw1/lKXskVTNI+SUpb4/7bOascANUbyIw2hZC
+GbzANQebICDpkhjAua81VN0Vnedze8V8Z3zZMCjfCoZYiTBAyWvDNdhiR9h0N7iaxex85yBTHxn
5CtF3sRFT1w00CZ05wHZqE56LgXzLAaFHtZRgMOPlzjRf0ur1COz0ttFmRSBa30+tErtoJt+sKmn
TD2mvFQSHrduS9GjQB0JwVglxspqbWOwriBBmHsUuuYjJIuc8OOf3KQ1HUEu50kHheKkGT3np6n+
Rpm8BNYlsnlPB3v28K4xCyokjNrRdkNOuIgTjKEy6qUaKVXsBsfzmZfupqIcp96DpS7xh61g9Y2d
ZQW85gt98KtKQu72JlF6Pez+vSRMrPr0gLLjemmTKzw4SIOL10d8Kv5XBOtCE0Sl/oXrem9Rtqgh
+iZmvmGSYaJixfv5TPiaeWVotZHrDmHS63Dgs7hpJRgHNUa760+Sc7ncsaTH/q1GR311xrDG+mDL
LF1Uxuy3ozo9v6+QQwJbFaxEI7SesOTWvj99BXxZ09x//dz0dmmx8sSZb/SNO4aOjdhxLtwfiF8J
jtjsp2OXIYVLmjnr3cUC1oEvNCRqK60P4r2MgPI2+o1S3IWY4BF219SJ4lFBfEDR+J3Oi8vSt0HW
CUazpea01jH+VHy0WHZLZLzZsN1KiBJgf2KwTK1nPmqgnKd/F6+6P1FuncCl5ke1bscIPpQgBZKI
CvZhSbCquwLwVVZf3JSXveYCgNEnaePjSc3M6Pjf8oGn5WYSSg15Psy4hyRC38gDGtN70HliXqRp
Ag3qUTR2DNsqPIzngHZFV3m3ueI86OIYC/kTi3sssB7yBIDgeyzeDXU1+CsKnmBsaCzQYo4N3n+9
0Q7re7ttQ8/ueuCM/iWIoH1CoKKS8edMDG9XR3nkRDxWRc91jco7sN9O5lXR71tm8PEaCWjWASWZ
KUFY2KLoMMl8d1ueH+TY23HAPoXmmQKftqDLdtDaTP+nhnQSQ1zAE6qeLIMUs7Tpe8SadW6Btqjf
1A3cBuchvKhfw3CkCJtbHWRKrJOd6pZKvOKiEg/i1WszsJli7Egq65fKrIpXCEnPyNYMJ1QAw5O/
csxA3Qxj0hrml8f9eYj7f/gpi7A1Zhkf/+bcSocBXAHJhd2SzNaycNjkNwM4TJSuLPVZytuZoMpv
u//EN0UDqaBuR2BjiJogGT+KhttFk2lks5oIzEnH45eRKy4cf4PavGrqN5/LxRVXmV2T2kTIwJGZ
rB0reDBNVJVWN7Ata+5+byd9UEE8wVrwzGRvvJFFWOkqcmvMchX4Nn/N5aJ+4t9p/MIeP7FY06Rq
lmsW5VdKZePO3kWl6v5Nk1tBNZ6vQCN+cWtv09JBvEqV+7Ctnixm3IENcQTtTdoQc6AsueUTpeXG
PPjMpAHc5d1+EIZjI9wn/bsF11BOom/xznrsolzBYbdYv2/4fzJHPx5c6RryOl9yp+iICF+ucRq/
MaCpRw0pk2L4mvLwS5l8nKX/MKKjDGSThDT8AfjKwVVpoHyHpZC3RuzLPzKiBUp4qmZWYzL8higZ
VOKSsmORwoIsfvklyG9dHTI0XtcGrk29wHKaAakA5lAEjAPWoeR8qjGZEe16msS25UX0Ltjx50hP
o6h5WJHJK7sCbyA9qFzoVRa5YLXIS94V2HYrR2PinFmn3059Va5IXB3yXPtpG5PrDzlAUPN1dTZ2
DR0baG6ZMMuAi8d6O3NcsSDhU63IaGDXnvQZJzpfajnOfi3rkI9H9OfjeywyuDiQAXAxnjmqeN3A
fRgQgReI7oEw+tAEpV9aXkRDw0bU7iggmNsy+RBOyUfNUd9h783s1qcX+I9ih2PmK0JbVsMDAjFm
TUS4hmAocetognUeuFoJ0eIW4V4AptZYbiSIPAeh4IRPQZkHeIp3BkN+sv4mODF2zZTTuuB6GKt/
569a+qqv38MfcM20hrAiY3RbTRJ7VYgAsGiH87n+HSr3fgCs+GuADwuj181J91ClW7kR00I/0aNE
G4KIg4zRTHH3M2MzHVm8eNxfthK8rzqwCW802UBSDnVjWhHLa/1L3Nzi2WoKXT2z7MU83U0KRSjI
EFEvCgMK/6OJb4rRW3JP2wkRlx2Cio1DR/he5T3vnQj5ycqdvlfXcqaavrgXkUhvzl7+Q3dh8bEE
4EhSRCuH7VSNTGU2VTKZmmgOimF7zqEtvcvJA9guI3yf50O8XNw/21EY+Sp5eFRBxnLyEyM8I8mm
oOEk+NN1e2Gu2MxNvsCRSH2n8kghO5MNMrnVrUJOc7kgZ2b/aWo2xyUQeY9T1zNZpLcq/eies+7+
+GWRanrEn+jgRxjUSv9xAs3tK1RnkfeQ9QWz9zKugHCWXwxQEX/jr/MTcQPivQDYFj6otYHVo0fK
IfUZcEq1MhiAWhBPwCbf1PVEMle49/ATbP2PP+MmKbmspLbIld9OUZD/WQtKuYCD3hLSi4unLU7j
5S9GBBdVdI2n1YZZ3U68RJL9CvIruGX3yzbBOaDbdp/U5K7lclHkYtkVt6l81KGgwfv4y7eUHASz
tNJWlIPtEHLXGuE5p504HMV5CswkHKECJrCpXcysF7GD3boHiGM30bSB8dr8vFhlrjqPQ3+masPY
E9X3gpXcwdPS9E+mz6BJ4cHqkHi92oZwolOAwjSGKfFn5zYSigR6bxL6Nva5/HVa5X4tUP9oEdsl
sKJDejC9TC3wA3kbY9ZukorhemmurM/lgwFYHD6uBvEQ4sj079xnwpJTUgMqWntND9iAwRKJ0a9a
h4oF5acPAP6P1u64VDfpV/4li3GJ3TF/737rENcOQW5v63o7tijkdlTKH/lFFCjQYwXgUD5pO/kB
1p3wb1mkwRPGApipClnq1lwVShgO7cE2PiJ2CjfaPYceIXB9EAb46YLDdtPgvfM9vLvowe2s6PW/
YFOUjVTPHGUlJ3HbFQE1AVxnRoB7Tck1gBdPXEMbHCDI+o5BYTOM1F98qccRm3MhcA+mF7pi3sDW
Jf2L3lr9kBlc6OAUTAWSuW5/xnc/v3eTUSmnW5fi7+gPSJmj7M/cPTkmNatOQetDNPKkOYGUGbi7
keyO1luUejRdU+tuI36eqQgsCyOX7Vo9CBSugLANVV3xjsrj9Bx1QNqzEfuEZoI6Dn2+kfv583El
XNO1V91BrEFtjKzz5fielZveInFM6JInAm/nqiS3y382aFq0df/q6vDBWko++dLTN5H7LxwDrbZZ
rydZoO6moB2F9ZDoje/vtuHTS9EIFLJGDLhZ0BINo1GQOnW28HvtmB53DrjWFE3mOz78iO9HvLLd
dzMu+fLVtWms91oeXl3EW/kWUiuSwBI9CXwpv6vKPG9cBrJSp0o24EE2ItMwSqjRhYLhaPphGutX
Uq2bbzDO329kd6EY9ySouiN21VDBFL7KCrF1qSc4YkKr3zsZ3YluXl/mSxSFvRJIgnsOwQCBRPXO
oJIfiSlH2674bQtMxar6ZEOdHRS9Rvd1o+GZubiHzjUy4TdG5XpYQkSwxC8wHHtEdsEtlkxBtPZs
8DsDxjjlBgsShg02A/2tU79pRlaeTOcdv9L7pX7dNDtNy9o3gs9HYKTiTteYIiyk/2aplkSymAle
ZJWuCYkvTPqNQCdH7SsNjwZbvPGQ610LV4CDrqU6E47+q2oo8asqvyIz4jEEFY7t6Nhzpzc9Th/l
UzHpy/S9tWDE62flmQxgVw1/FiBrIApICxxERV83mfszpXX9eUWd/hN2IdzjmPkskVbwJy7wyyoa
GUL7n1WiRK6gskA2wZ+OvsrrG6VpdwqMxhIQRS5ORb31DmbZCt5Oaa0WcVr44ebX/Jj+NR0T4JEU
Ub7LZhoJDl7WXvT5aDSChGDAJg6TuPRG7/vyufUxcbbANkdUtN8HeNwHUQVi3LRrnQXzbhsL8wZu
M5LfVl9dnKRDS8tDCtBNQbeI2/ZNEk2gGpmywj1ZxT4RSP46NOmMFGoaBOBJALrHbLdYIWZlNhQM
la4XnHBKH/BTTpOR25v/lelNCuRyDaJI1ETnJu9sw2MB3v4RC0Z9AFs8yNnQecwfDw5dAdDxkJSF
4JZxNRmquO7InuRh8fVBINmBe24b64zDBLzR4/8KndLK139FWZUdynw4g2HmW7ukKsW6AP4ezXaF
poe1rKG4O/Z/btX6rvasdP/Ij4h0uSnirKiR7vncVH2FNj6aGiVswGEHkNq0iAsQWqfVDMUymPms
Xj43IZ7Tx2kBqXQ96rou3Dqck2zX18d+mO8Upkfwig18d9k7bkJ71FY+w4oRX0omoAH/+dMcvTa7
fbaw782+7v47yIcbm8ywUVLTLbr6iABFg/BrxKK21cznl4KrkhmnXHppJe5Vo5Uxq2BWUX6I/sHL
lf2C+zyCjxOzFo+KjyI7lhNfF3CxCqOIlEadEbRjNRNdjPJTTGkVYs/IVVJouK88QYHlw6EO3kXi
DTIzNtcKQO5k25GP+0zM1dzo44VUXI7Pbt3op7haD1KadvitsUlLjwWYjRYOs1mkhY6VGwNbpbRt
K27BbHI6R0PXbVNXOKaHMXkxZuvM/J7LzFg6pqtG+x6gM8bQHLuwyUJrMRjbKETMjDZqFBXe/XrW
Fp8usCujUJH718BAdwb71jTUtzer61SsgPa6GxKHNU1A3HXJx06RPJEEwSQxy9hzPh2vTYSTXYc6
5LSXo791jZT6woSjJScJ9vuHeq70jqsd5IOW90SH9SdA6p5mvy2MsPk2E+IdpOMZZd6fndEBEuB+
XReYWiYo6ewJ9askaXhIWceF9vUv9IiOG6DGKgqHZLgPwf5dZMi3aHlj+1F/HFn8bkaLEeUsUp6D
d0xqzdVI6E6cXZNbdjAOLpLpju4Yex+y3kdOF2BoZDU4YumdMPRsL+ngW9GuSof3waMa0H7L/kB6
LDd0kjCp8xhMY7zl5WtDJbdwcSnfj8TuV2+FL0SpSNHw5oc5RvxTjMxIdhVwX3LKnQfVCXRU74BA
qr+QuF+XbxMiBr/0WtkFFkY3oYy9x+OYu+2Prz5a/uquhjMaQcQ8H3BgOQoPAgPPP3Xtij/SSFNR
23Sd0Xp5ynLW7rAA2XDDZqEZoUKhH0cePUDumoXWDcMTPYD2RjATuwIOYG5roRClJpv56sWdTsWM
z1Gcf7gimp39VL+JgfJtxF0ixN8yIQSEZ8cu4bz/10Im04oUM0DaRcCBvmbSOQ5/82fcyXLHhvDd
cRC6qxMLNndu22ldEsdmcUA0iXF5IM0F4uLBq2hXovS8/1G35RBBihHEyCEPHblZ6qgCQI4B3ifc
aQ4mX/+Y7OZVy8S0Q/a05nxJqD45Sm2lgO5B7OqLZrk0KYBP6twtKJ/f24k15n8gXkOBHAkKiqoD
ckwK9bv5naQYl4/Z1Tzi7D/HnwLKPogyXf8HsLU+TPvRWu9tzaogTeeG+PTkCn0X7D/ZpZf1smyA
pTa20QHTe9bttVAmiMcXtQkjtnMfuYcsrbx+kbI8wOw7UlAEJdzkXStu79Tmt9go+kIapXJbZ84Y
tbM/NowLqOxJG6Bsjx5z0zcO44ARhtBYCDOUPXVuUzQxPoDfYFx/8REhzCnQol/CUcrYjQ56wK8g
9s/VPRFEPOgCFnBQOEP8+kS29Siw5xPTlZcB6pWOf4dt5RJDDIE75jpiJigEtMHvhohNEqKgSIDe
yuypt/RT10toqua3tFGfbd457eFwaJNcoE3VzPieWjp8H2HivYreguwAUGT5O440lmyhcCASWQXx
ZTVoxTmeB8nam6EhCpWOv29LvUsgTbiBsl6VMVMEoDfhWc1Fjp9D2i8QTxzvIwTNsIHydvvFlU0T
lPyD47t82jvytw9uZd6m6KmW4+6MzgIZFuZZU/ZFNd1Lwnhh9ORI6y8SBsaNvMglj/6WjcW/hGT7
ui3WFZKjxFrSkxVXYwu3qlij59RZl3yud7n75dMDG5Z3uNU4hMH40vfLNCSKqeQWFHp4uMsJdVfL
reLKeKeI22dMrX+j9rCNRPGcZTdY8+QIf7j95eix2SZR5XTQUqJWtLXzPev+UHut4Kqekqq3dHQv
gvDLUNiu5TfbfXEe0jowIpfzS02KrYNj/lq2DjnzUhKbrsW4B1/1R4VzugvZip7Va/64hM4vMU/c
HN9AIDhBZTe95o2wnMwAUAOqohsZS9IOSoYNdWY27Yf1w/WZFuFg2q5jxU8te+Zap5+k0Nr2hYZ9
LPUdDMbpF5SoYziJ+3v1xRwEo2JAq3+HZ2dEgxrG/vNCL3KlmPLSYP72iIpv2VzDV3N6HxHSWnAn
26s+yO0kfRusQTc3+eh22FtezqyJua9e4aok+txs5w+bo5HmfqZZe69de2w8FffFMVOs5EewYpCK
wc5Muhf/uaSrgE8xV7IF8/AtdF4Mlgj6l/hdvcMurzik8w/r6FpoyDs04zp1lHov6z78JAJVDUSG
cuQ7KdAdZiqm/hBixGTInuas1G92EXxR92h9vy1Bxms2C09V759Ro6xd0tJ17HXjv5WJYPXnaYbL
H3w8VQA86LlP62YkqXUMp7pHdMFtpGTjBziaK1QzR8ZAKOGNn16g7PWbcCk7pvLbtsqznz0oRKQM
tXBsoU7JVOZSWMkTSJ6+t+/xjD7ONHybja02Q/y8WA39P9MFHCvfQwISiE2UkC3VBDO1cVs60642
z/qvNFzqKLoBt70CbHrwju1WQTZeAta/V7dXsukVDVOGJBMuIhmlLAyw0jpvR/xdW0yVwAneLRf2
i9Dtab14PB9pFg+zZxCrC5wkJIPaeuQcXvhauy1W0BXDmPlxytCei+ZQEY8BdW8x2HVMVEL20u0S
7zM8QgisGGQa6l07g3DX6dvTPRPZqURtKoBCuzXi2g05Qp3EpBeYCBH7h9ymnLHk6c/eJUal8otX
vByX58KTie7TUMoTWnVPGrE0IPrxeRXJ4baU4ewJHNbXhxnRDvBPYlu+O2Dsbr9M0rzCAZ7VTllp
PxScKZ074h/tdhgmNjc/ZijWsS7cC/xUNxY09XSTS4y6pUSEXga0UQEPrf8247WPYFL2lW6X8uoA
LlwHYDfJIK1SXcJXhhIIPwau4OdiNPyf/gTjqjCj5RsmbFB6aqzG6otwTSvKnFbrKLmU2B4YwGbM
PV2aN1Ig1+E5B0ecGfFzhoQQM71AFUw0ximjXqTucictf355kLJy1jb9opUTA8o2U/NsrjJo7iaU
XYvZkwXk4WdVjiwpynjHHXA29KaKnGiU+pp9uyReh86odahnLnWRSvJfNRh7InMv46wEkACO0DYg
hnbvlK1T1axS7Nkonk1ir/S81cI9h78To1o0StU2j5bIlROff6g4bngyCtE2xrDXobD3iKFzEx7l
lcTm6SrLovWbC4YJf5OIRvbFye2D92cQm9MxE1QopIGn/YnV+H7KRmokVFrRMJamulLujThPyf69
jlr6iIEhdDDdNywQnQZ7+0imxLZ9RjFtswwZuuWc4PeqJj1HreHvQyZgHM2Z1t5ijReIigRq8san
GEaRvUBRYYnKeszh+1CTrNhEmpKe0EeNtC9XK2yeAkDVs+gaPo4FcyNBZCAVi9t1Amktlm019atJ
JH/9X340lYC5vjV5hSWM7k99ThieGtrjho7JrsM7olrvl9vovnrXU7gz9kr5HYIn0j1OO/+XecuM
BQ2vb9BGcwNOTT7JRG1XG/4fIVh9ekzuV//CxBmAUajefckOVhNvXg1Q7/784GXNnmM52/IMPjnU
GKyyCqzruBffHrZjqyJ22Z51gGoHAsyE5fhpG9iKhacW4uMtmDsRt9fDsfNaUqF2O5/rjGMYBt+y
24EedMghOC3hSZeGiEFutJsmOl8EUf5iPJdmRjzJErjJeZkviPUCUKfQCvKQV6P5fXBZWuA9U/O6
pBpdokUEyhL0/5O1joOZcMlaH423vpnGvlfdwbCF2l5ZfS4OJ3aVqMcPZRmxOKbi++9Uu8juCgn4
1scbYLaOZlkXbGsC+5OoUExQ50PF0vvIW4P1gOEJAlWdtFou8XAuS/r8m0CWQp5gYysLaMa9oCNO
FzfSEzAY1HqFDQKjQd9OB7gayPWpJt9F54kWFL/hs3wj1CicuAkqgZjejFdvL3fup89jfJcjrjtU
rX8ruQbg4tQdRXFOZPJme733e34a5F1CQ0vt5agguY95g8c+peepz3BXRHuEWQkrwNEi0J1u04SB
2EhWtEYXitsf/E9AZXbiobLj83B04ULtPshavc1M3GKZDG2wH6xao1f6b1nYS/djh2sG0dYJK/Qw
Wq1ahuilOmnhmupxr+XoUis8/f7GPGDQG+xLeBs85HYqjNg1NrsBmxZBXrk/jtmd4ca9acY8u5Rv
CXIeuMg6ZwUZHOAqjqm17InvimBpxREk3s2vXaIJ2vAvCfMny4LSNoYPZi4VtkxnBInO8Jl7l7oG
keArlgwD4oLhxmwkqXp0DKbo2RxCRfeTDlA1HvCPpAiFgbaNUtRB0APFMBxDzroTrGkCEcIVu52U
cIwgzPcKF3x1wEWe6DRZgBbMBRGK6n+ZEgxZ0Hula1Agi4RY3kUGAyUQ5iPrIngLQqSbXkYWgzNx
Gi/ByaIO88Sb5xqnM+IXoiGg+jAv534Ncu1+7A9saOrOnYaPisJ3NVryO9dcx84C5XuvcSeSRft9
Rfjn6677vPIhAnf80k498NHOpcFZava1mQyYHQ6fTMVue5hfSoYaJJJoe+QBiCYZz39Y9y6I07aV
LH75QjJP1p+XDdGYkjOAqtrzaJB1rDFXKrFKPKvhQIy7ESk0qNI9gP5vjnzaOGN1JTct2JXUdxO2
Nu0ccTL671uqIal9VQxl+EYlXkxMNRX/6TNZFBchWJ9tolA3OdmvzbijS5U//NxldwFVvCeAbKdW
/u7iKlp6fhpHeW3qTPZx884gRcVrSNy+7ce9FhhzsQRIrgRp5MrbopWFOH6DsSSJno0cw0m7Ongh
CFADYceAw2AktlKwx9ZP214DNeMI8LF5ssDu/PRs4wpfT/t/T2tHjE8aAp//p85ahl/bfBuue4dc
z7y+ugT98CCS3QBfU04A6cRHosv3TTUmwNK6fSaBuiEv5HOVPkQHTt+Ol+WBuoNUp6+vqsBk3AIo
UMBWje2bW6zTzcoH5Dw0YSIqpqoDyv4AjvThs2QTOnZpvzJe8/iH69PpeECL2vuKLMc4JCBTx/QE
vxCvzDj3Gq55F6/VliZLSZ/eEb2U5yesjBE3LcH6pn6TpikjCflkANLwmGevhYg/CK+Y4cfNAI1L
lXC1i6zjPepNSCOYJOLtsMYpCExmp4EB/r1m/Pzk41BECsPRER5B8kVpYjtkpdWiRYgjxS1NmYze
0gd3tahrj/4lwip51VgqbQxd+ERc04eRwqzHU5Ne4bdj+228DIWUfFWam5u20HQXsCJyWUjsXhL+
jcPxijk3eRbqG7IcupSDcJ+cgZjPuDUY1yAz9tdlAWpiAaVs8uTW3ieGKeN087EgLsUZ9bJzEMsT
7CU+WH/Xikk1l3EOGZkCR1C2XDkHR8taE4mRV0oT9EVmDhEtjrJHfCKmcDgJXiwpSoNnd6jhExrF
AeVa17sHo55QXzdtq0kD/cFTcev2nApXR11+nTo6jA/3OmaYgje6Wq0csLAhIphbuqLxjtwsp389
E2JKVfK1jISYYdPenNe3xp1BO0EoMkKvuQ4PPu77rEsx9WDlr8BEw8KwMLsxwTuMivPq92N9pujd
kAx+7kIgjEetVI+FJR8beMFMR+HHKYwKlPV472Z7rsltWMBS5rgm1PBNHl8VlsIDMzudkY0i9qtp
al3FRPBM6LokzOYUlh9smiayK0a1pIzXnm3lfLFXb7XOjCO6LVpp6RDsckOW87jnVKvUp9NGv2Od
PLXo/Mmxf6+WHjEn8hWLPMHqs5VttyaLvZ1Upy6OzK/p04REVjrDhHfVasoD2SO5vaJAQ9ir8d3/
90H1czx5N8eqFPKMuBuh0/2jBDyPLQyfMdjXwLW4X45xUpHeYmPE4YWkMWTwFzNB4AfE8s8KbK5Q
RN+OXmDq3w1LHe5tEhgFwCBAJNTnFudZc3WTKKCPOtw/QSeWLGwBtZ/x1dV70yUEQv4Hf54smdFy
7Y1XyMICj8aQQ9DS563kvIUHcj04X3eowff/MGGmB4soKOo6FGTZKzl1174xJzCnow3RGJYyJt0F
OmcfVbbkPuE4zNXAcnIJxmEblTegnyxfF9DQea+9reuv29Q0BipfMzofXSM4ck6KFLN4sGAGu416
qmBVJ0lzOzyUhG+SzgstFqhJxQv4IhowYCTm/J5haPhB8lnoPAKU1swm9Yb8izgnAHeYq2Q+9iRe
b5qmvx6dI6f9g47q0pjGyZzCEDb6GAhOc1DJtaJ5rahjvkilUhMoJRgY9Naze0my/7BNzMpZgQ4N
RGO3Ch6FANDE05sGZ5RRmeKJXtUZHBawM6FMbDQcdapnSwFH0F4f8dfmS1lMYbFYwAWkkea6poHl
WI8RtJB58iIrONHw3FeZS2vzAeCIV4SP7tsjl5/eDlvSCFuZT8fxu1tZYIsJ5pjqVA3vHfB/Yx7S
Rn4s3oQIYddeGrytAak/S7yJHLEBbVUkyOWsZCAGdlaKgrFhRMSPCJyXCWjpaNpUaL+nX7D213iU
PvxieDS59SK1icYQKpepJzsE5xRiPOtTmZ3RJe0GsPJnRnUs1p4oYIcFc4F8bbuwzFIG7INXn6ZA
w91sXiwZm+FYap1KgRIAnZ4fBEB5le/hLbtxOhbP9eKKnnzhEIjm8rWb4NLXQvVIYlz4lErBdzaj
EO4xNFYvTftuc3SzowFIFIKyK7oYb78CelkoHPGczAcj026zjU29hbZ56mgPrwYBjwWvfFbfcG3k
ZXcSP38jGyUUgyWx1ila4l5oYsznKTMjO8TQsl+2KmS6aZCWpX4Pk2ebKBh82xvqmknidq6OR3Ex
psBlRH1xEjO7yegmHIaFU+CTFBoSD9qmQW/2f4ZGoF2PWnb4C/EF8KXcmSN5YfgMqSkIBPAqKd0V
FoAIelW6UnTvX19bh2jp62iMlRRhhz10kuM3PkxHlDRib512KO4QVySwIfSz2jdeMRSGB2bXIxPy
IN1PWjbztwFaABOOxGcOaU2eK/y1niKn6XCLpG67OqzcRTLmVnuJscvyh6eud7HzMOoYAlqMkS+h
BIH9LOerwNghC023dU+NUo4aX947g9b377hRNGeQd9wysskQ9WcdTjmbqFmb8EWcd3FpyLxdfEUP
OuP74rCWydkm+Nuvxw82AVta7Zs1NwJEyDm1kjOx/sV6sEhlKDxFylmxgJN102TXsSnWdTK44Sc0
7uFwCCICJyOorRkjEtTF6fhnH2hS8VVt0FFnms+PsuIhQ08Bm/FuDgOhedTo4oTzUp50rz0pw1eP
ZWnJmOGV49gINTBdVZH6rqo+OAjefo2DwvWfmfnW8ju1f865Fb+opblym7IQNwP4Aqp8dtfj9epa
6PZNyGmE8pgGtliAJaCtaLosXz5+e2D9Qr+eyHKxxH0p464XU4KIpBgsVkQ7yZHm4FyF0BKR/Wkr
/nmSjlAmZF4tkeqf2sxzqR5a+pYjAO3Ac0V/xrtWxtlGUKKPTLYTqaOX+UNmX+BqX5J0BIgaD6x0
n3Nz2ULCkgO+xQXtfwWAggtnwdPPUpSDXGjBDHikPYeAqaEJ5iiZxDOa9v7/dmag2o5wCXWvzHl+
0E2Bt606CrqbkQrX
`protect end_protected

