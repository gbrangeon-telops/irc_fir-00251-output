

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
gqDFw5NFAM6CTSTQpb6ewV0dkTDze+wC3QoGAxwxbjcNW9/DsOht+2F009+7g6jE2OnhGLtqTq+c
HspFg2GBAA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
OROCzcjj1wgCYlIqlabkGZopoXwccuhDPoDiFwbBlsbzl7flKX8tC5m+07o0XejIs9tQT70vCTz8
eor9UB573WqZyEwu6nS7RfReZTn9rXIEfFTmb5LNQYR53WQufFJWXVGGzbi12Azu0TUMNBykYjra
GCJvYkOLjulS+N02/QU=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
y306+4wGPVAAsHa7Tcr0Z+Y/dNy6G34dYeGbx7ATqkdiT3xoZwFMriTbyxCB/BNDpEEpWtR2x6B5
1geIXl7xRsYW2a/OzYZ1VgC14cIMMrlyvjd+Q0oeBhNwIf7zzOU0YeLe10Ln0VhNNlM9hG1yxJpm
PklN0o7dbe4z3qSMhzdrqG9CNO1AfE0zEYRDe4xK7ci9EcGBPeIBnjhSSGUwaUeKV6BzeVeTBH5k
pFfAdDfvgi3P1VwvurSSAL/VyrhWR7M2OhP7fekXRqEU99K00pFciI0NAEcJPUl8pbYtjc86ccu3
OmuQ0fZKcUeaRlPX6glqeiiehMLm/EPWzCdMgg==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
gSn/ibMO73s4UyV+DQBAOvPjnov0A3ONpbzDn5S1gDHbJc8laliw/uAOvABs0KKAN8Q7GKr5UYxh
qWYO6FhJPBG8V6RCU+sAaoeSnleJb/buC83HgJws4chUKE1EbA08UnkA2E57wCSfAlSkdEQl5xrl
E4NsCY7zrBmnjMH1Xu4=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
lI1FhNfWvnI088CMtuEIyHMeXPGNhtlppeaUXaQvRzrpC6F1bRvO696fznybaYq7K8VPJB0YyXVb
8oCJzTtV2jMI6KoF+McAzbvubpz0ru0XOCjjvcTsZJ3kGxHGUlKh6xdlB0Gez6kASJJe4GeTuEaI
VZNg+Q6ea8OLPKgQf7VICmBv1vM4svyVLDI/pSGiGOmfSMrfWDP60zo6tHpkaDS7uHEj2WN7lXT+
Q8c1SGnQvLeKyHV/kGG66fpNSvILAslBR0l5Xt1/csaBtahK2IV70dxaZkLZ2c3pylf+SxXTt7v2
CzVvxEgWwmwKjiuhBgmVM6qeL7+tokO6P+FlQw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 41056)
`protect data_block
mu4efmmOsbqi88SmXPIHtq1sPOnJw4g6SEpKsNceW4t1KAHKXrj5BOootACoQkyBgcmeeCDM8A2f
SXWSb/uTc4ffmzsoVBSk4W3RmEUJKpuGKM3ELmUn4owB9uVDlhEtubulrScpRPFTk6JS4w4mNqeN
SYTdFoeUTquyYPED/jWMVgOub5Gl6CnRW8JRnNzz7wOLQx//l//ZtzqF7kPCjOSMwTIMPlxIK1Cm
Z3okGQEmKFzoBSvcropQa1IQA/0j1+vA8z+cEYRhWznYLSOIxnKko8tJ/0uynX0Zkfrwxjs35SdJ
XSVKRojuXX50fgfUWnZapoVrW/IeyPPrcfu02C0VniiGdYjWtogpfDQEdA5w2FyzHAga2wUC6Z5l
64hGvGylLYbzBpKb4FoVmgQg2juWH+i0jT9ROzYLCY73VFKiVtocXLGHzQKhocVIUJsJaIJ5dbAf
lMNyVh8MkspIbJL+VFdbIm4vaf6RyL9IL4S7AcByPhokwGmEFrnQRVfmGpKbz+bZ2Z/NNmUx3Xrw
mAnHxDcG8DHGTRBAPi7KfVSK5TID+SeRyKH66aFgRNmzdt94VHZKG/lETCU9QDaNyToxMIgzOA71
HRJU3r1o5alXGNGrIPyls8jw9m0CoqrkNMP5N3MQq0+C34TF5xXcC+otHjDnO1MFjMCOaUfY4+Pg
lSJSjyEdmW6ptRR7sJFoO6rEK36RZTwtkOX1IRbsrj3v9VR5F/xnU7ic8pmmVAA1Wa2YityQRsiy
lXYzahthKxrlMdayY5m/6N7nkaH568+o/aqqyAxkmb9/rSqIo9O4OaNbGebql8rfn3qfxjjBPLSp
U6WHDZZclFV+3RGJSGLXE60R2qTs5GNYRkVRzakjeDq86F92B6gH1uPoma+Jjwnv10+29UlckD53
SWuUiFKB4EBv1WaWLoYUWbz1bwhuNhBq7+XUCqzkrdH5n8ZIFW4RPrcT+dAfR4kk3tlcuonJydvj
UChP5AUpXNzplruSOCaVPUkymRUpjFDIAhhz+pURPqy5hF56uoEGum6te6VnD+o6blWAoJjT/nE+
R+oPwiMHWQK8Gz48AFoa8OmhtbBBLLJm8/ncWcb6tEagq2xYS5wwZQNGTB0ZHyJvkWGB/8utQDwT
QZvMUm7Fz82QHQXP3fbthfUgeAyQMJtsA5a/Lf6BLw4MJZpA0Yz9JTkxhKCgqcrDxATi1/bABs2e
IC842GfgFXEvEB74HFjMmfV8I639hOSHwDQ/wx6wr1yTswErmtFs+c7ci04XnJ9fimASYxg1lXR7
aoEvCtC2Htld84foIj2IRC4uIMmNP8Ye1s8yy7sXBNhGtFAiCYdXh4JIXHwxwbw2vw5lbcJT5fM6
fT5ALA+HmGnCoViuZHpK+uuq7v+YiVej6UeP2cTPEaMjxqb8CYDy5uJlYKI7Zz7jlQ3jUZLRbYZS
hC5zzMkk2C8pFeiHOn1TG8bu7O6EsKhGyolOe4aVRNQ4i4T+uHrqypaEycWm1M44mo8sLO1o32y1
DsuclvLT4INiR+6niH7JUIgs/jE0tNat9GIDFHmBLJQxsBucAD6CmxfoGW0GimolTpQrI6Bk6Cjh
r1/JcbvwW2FQ04wsH4FaoiGfPXEL73tZFOAnygo6hp4TQlvbohBCjAZ1BtNK/2Y7rnBp2RtcWd3A
KfJleEaZVxETqofOAEvQ8lZ0DGJTJpsCc57fA24+pvwP72drMVZBkVGq2R0OsNR4JR4YcO/4RHkF
uy9bX1cJVnSgsHiVRmjfTvzJnfJOet9sgFE5nSxnVmZU28qI7RZdXEbKzde0mQARCnd/9Zh7Lkw9
gGCsufngf/3G+LPTbxBIUPG3VrrPDohE2uCpwoq+2QYzXALwpMWF3hqynRlhBxLaexiGI0dCfhhv
gczfxfcQu2J4DPRWTyklzRSTTHcZJeVnefYl5KRnpx15A15lOxtK2RkJaC2HXCqQVkgVwcf0kkrX
Vhc8DCg1mIShDhy9fx70dPgkxULhg6dkD/gMm+j/vhOnXfyNMgQC1kBTKuKozFm8tCIRiZbNsJBm
SuPipRzwCtTvMbvI73ZEVghY2E5DevLUycAWv8/kGPGR3LwOaW2uYlqeWbx2la0h9JstUQls/hzW
0kp2iMHa4lpk8jw7ElsgFhmPjPGlMwhaNBj/c/o38+0JqsUc6tqEPAKNBaNNsGfqOWeACjM5OI2C
mQuo8xZx5c870quimrTy1yGXDeRDcgTXzsEKfGXgG2OWaAWMxhlujqMinkRz8AxmffOQUXHkkKl5
8A6lsswxg3r4XlcE6kd3YXQDfF7woHDyqqL1pcmtACPY/zcW7ZqaR2njVZ1lq5epVPLY2YVCI/SO
zdGeyjKrO430P/XVl6lw/ASVYgK6qLIp5GoXJczfigbdaol40TZCtZx7Pte0gqY+1MieMkkqqJkT
GSOudESTkmmAra2ZdGgewrcP/WZ4FtVn+el81IxTs6KBsJyOd5HGophVA8w/vG/B3YbM5JKAXHWb
F5LJ2VtKB4GnmVOZ9Ylo5SlYcp4lpS8CefMwzwVZRCI5Lc2KiYcuH8A1+lwUOYKnE81ZUJVWCsGV
qQd4SxAY2mBGPAvWM2oCY+U7FCb4FdazAWTv2oNG8Ci7g2VzAubFoXbsodbVzUSTeY9aJdnz9c8r
jEtJr80dI6aAlXhdz7PiiXedqhL9fSx4eoeKVsREKt32lma6NEPYZrbUKCmqcLYsbSQHcN05JLSF
U4hImCJ76Ps1jDrwRUwMfiA6bbANrWSKeNucQBq24z/UdE+Z1AuD3/IQxjZINMfC8uDVxuX/dYvL
PzwkPo4AwTbdNiG3i9LxVeDqFoHVvPAr6nYeoqmt4N63/Jybrj2bk5a3CFn/irTaJhDGVX8NP6iz
qtkDrfLjP0bYDRRHNMSek+QvtQ/WkYGRGaAE7phF469mumTINBlj3HZqqybe5zUVEDxhNjN7BQqm
eZOT9DeVueqUh6TsSqBHS0vrcpMDjt6EmOPe7GSOl2Z2XkwY/3lHCyWNqatJpNzZZDeud7YALHhR
00xY2QlKwm15tc49ZuGXsXi+1rayejS5bnZE2n/DRZB7Y5FYHFL5WbmeW6Prc2w1Y6oFLr1CJ5LL
D3Kz2njMrRVw16ZfUnAfDBWC5rFtOq4JRt3KTnpnZisCHSOKfaNXzrfxwYmb88lZpCd/D5+ik4Y1
8pJf1P7gttptIzIG4HZ72aWCzF4uW1K9n7+JsF29lorBOUNtbmcumVhUR0KZ63eIV5gR2HtzMYka
hrb5NJoJJAikQlDTXZCP3/8N/zDjKxHEZ/XbrsHtSDw9ti6MP2jcDExSZFFZDDx2IQGts1GXmOf4
vF/SjvqwDBrxUw4ZEzeSvj9rx8bp3J/28H4vn/2qmKtpsQYha5en3pZBAgVaHs2BJPzTUHAa7OeS
V/O7eU/guR/lDu0lubXS0Mq17YsfWfwpyyQvqSCBMaJtQhnELhfYuWt337UrQG9xJRZganvCupKQ
kOjSZeQbjmdH2bGxBO9vPMHpIYlfnTJ8SLX2pHb1Se8cBpnW6tVnjH/iWwl828FvBC6E1mO3Rpy8
Va/uWurBfv4jihd3+KZgR5EXzsE9IPL1Pqc0T75hhPPAS3BSMwRuj6SC3KH0nAd0oACSG0hbOvBs
OaTHsnMDSTpnCaAX3snr9Y+kDX4+fX5RpTFBGLvRmFFalmjfrKVg/BRi2oagRwXT+95x8AU77awF
EiM0w5upf4XXM0VNLgD1kLcCnI/9BkrcYfXQCa0ykjxDtEvPK+o4/7rEkbnIUOlSEYxRegZsRlU0
twYOz017E0p/27QoLUZOsHpFttoZYUnnzEpUeU+gMr99PHVYzi2XAsqkGtsmj5CXxKBv8ulHhtXv
F3WfSTfwXb6BJ08S96L8GVlxvbkcE4v5Yj990gu6DH3WTfUCbIvucA2OCPjkMSij8CaoDfpjZKGu
UWsac4ejPfd7d7ebCQvh2ld0qk9FyN3ouwKvZPefD/8Yuct8uBs0SU35TdHaKmTxdze/Hg67EZNl
DypVEQezEWz9rupfUffQ4huOIgwn+aUgy7yMvfZyNjIWmGNbPJ/pmTwa+S/Xst8AaqN1lLuso/pZ
fV6Il9KVPUDmoHD/GykiJd5Z6oJoMcdAR50AiHRdiXcIn+sDtXpA3dcSvdzklGlExaTi5DLd2v3C
9bt0duN5zj9P/NvHU/6afeKJDqWtU85qQYw/tlGg+FW8EENgQ0lpvybaEQyI9bhuF59ZyJguWG3T
OcQMYiBzwVG/cZLVXUMNgF5zKMqf7SMq2N72v+ipzSY8hPImmk1QyBvwSuiBqiM1bIrMwmBzol46
3m5Wz+4nGc500m8ftyX/YkBEaOapVv6WR6vJ0B7Ltq4jGF1krXO6wtoK9oqXqiQApiKI+G5j8XgZ
X2Pl95rQqn74qk/ockLp9n+jQWWUAmTvHZsQRL4AT9owS/97D1Y7wH9Vad8rxK1YUF85VAkGtSCv
LHXBTXDOQn5hX2lxttK6OJg6hrLJ755nRF4E8bbklrYnWjxB4V81WYoaCQsn1o1WirdReEIKD3/n
MrxUR6jNcH0otuydLCVaYSnYf+LUl3ud+qGmsYLQ5iQqQ3EpDfdsb9kBwDBVQbKDVmY1cbbj34YZ
eeNCvBtkAL6JPkUrTl0nRMdrD0uUAKXV8CA2LmZNdgeRurks06AC1eat40Sh6vMfVrg08d8If8Eo
lPc5Rd763d55iOG78QCC1LaZZO6db88++AP2g7fKz44juxjO4sQkun3Nt1u2vvszernhQDLgpULd
VPsqKhe0YTop52JEtZIgj03Pf6ONsRg+r23Qqn6PuxJ9dCONZe1ZsodUw/wVw2hZF/eo0GqLSdnq
09sNp75EeF7X/Sf7G/6RmZ6Luq8a5z0Z82tHDHEoZ46aR2CwdItCYYiT1dik1pd83cRR7dcp86gx
M9ZeV84ys+arF3LgUapssvRWyTanneavgo1e3OTZylp+raGxHkigLe/MpdHmlRzVRgIHGT+9jY7x
WyaELE28TxxKC7IqegoWciBecZdrtYSjXGMykkvjXXzHWq3i7FohJgBg6cBHkEnKsWBaaDUILzKa
uU60uJVC5lRCUaL/bT/gAmMwt1cuMMQFeQATWAtovKCsAxvIcJaj+U+fH+64UqMx2LS8AAJFODap
2yEMojisTco9HM057zvMrrNNOX5+2Np4EjgneDFzpka7Bt0PDjvDGZkVBXOTleIXYc8BzMu2uOop
RT9uZO/SB1hoC+WjT/tCfuM1sjpbnIyWBISx+hjs7sEDjqzl5g6mDrOp85CEiOnwOk/vHIDOKOlf
jyGc/Uv7P1CScChhxnz4UEtBuZvQzvan+PYRELGicmtO3xm7MEB8TCDppOIET+3LRy9Wgugr6Fu9
tbxIZV9nFBTrzbLyioDOPyj+1Yg2p3pZ+x2CyiJDnvP3lXn0pczhmbOiuHu9aL+09hWFlSrT/6SY
JumeipUJBJ2SlsILYDzncGFc1Yz2XG9fsota0rZkqBzkRGQ8i4/SKVcGRGJ5LTLQ5q4r5w1E6dq6
lFcxb553bzAbPsNW+oLiVucqwop6ftiVpbr0NhrfHs0rGmfSvDO+rJ3b/JRFJDEZjIWuA5G2E/cC
4UvkMGXbhmasc5EVyVXS7/NV2J0npwjw6SoTQHjk26OGMEsGBGU3ZSl9WSBo6kkmehQXqMjwD7KH
k5/FPcnx+79rluGLfneBOwZrNN40j5SLGEmDa2WETrCGsLekb4NEOb/KmdOTVlgLbT9q0aKAU4Bo
kwY9PKycey2MGR3OdgNfIaciz7yY4WcnDniJCEIhYHKALtEnfhcXLqL4N6v8lNw1IyHJ6z+gGEPK
2LfU9skRXRd+aDKBtCA0HW2DHzcWTB5f0RgadANLb99KtWFJsydTTMo7yk0bAc46Rjuft+Y3C4U+
zEK82c6myHJq2C8mjxFWvDznpJ1ZqchucSshimDMoctvbN0i8nX0anaErTzRaax3SlIpGhTGpfW/
vX4WZ8i/gHnP2YFCOIEGi3TsrdNoIxYMg2UZ6xMi+F7zlePoIiN2g3mRIB6Ci/O7mAXAcu1JqMLb
wygGMtqAxRlC4Y/KxQ3l2+iX8UrGVEU4fyjYnkmxwTTI8wcRpnmOanc1ViLE3a8J5aUumPWS0ETP
0Bqc4OhF7aj7JDblw6ehR4tg/NIRaKYkJLNmqFHQjAvJ6EsOpKUr18zCqQloqssHj1uvmysNl+RM
IisK39KPOOSQpcIl1ge+quMukj2ETzL2FP2BJfPysk86dDCiI2rdkAr6wXBpyv9DB97aghVc5QCp
SJDzqFOMTuZRQ8LFlb/4PbRCsWsOMYOX9ZVcyxp6fMIS1dDZ107F195eeZRs6pxrLlrhNhxsKPxU
9r+DobnwIXbovUkre95OLfDx0Mqfe+jeepGcaCr5gcCuz43PT8dFF0zefCUXdMqI31C45k8GC7Dt
bv0ZatE3UKn8NNF4zuqat3UVmONbsohlkI6oNEUW6RNH+Np6U9gdOqUI4g7Bdq5afY4YqlOOA9NE
LYqrzNtnFhD1OqWp0Q5MR2kxBiUHJkacLaKn+edaDQR9GhWZrtmGIPEDJe2+GHVMuuwNF2qUdqcu
wBZgNf3Yfj28pSyV7RjJQJ2R86WV1+c/Yfel8ZKJZEvoWfGSctRx69LHm4pzpHot4TyK6eQicynW
V46LPMFDWbo+En6xHkt61kK2qWQZsWP5vpMY8fFH4TyhjCLmtwwSkwf8aRoS8Lftid4iDfifl7EB
OnUUHn9KPKoibeFeFIeOwFUI2sCrnWJgUUONq7L3my89sQQZU5PeTlvE2MJkrzwj+llZLDUqv9O2
bBrVHEOnoxTGmIW4GPC9lSgLzpJTax1GetXzVSRHGfBAWInoQsgm1FC6EsgXIsYpmHeLkoWbldmI
iyl7Jh3upKq5dGxaKn48CZUY+2QEPnMC7mDnzVx1sJ9Hl8yiVfFrUuosyzg1WH2e0tDWvxCAQ5ye
7lvV1JbjFRTlMsgop2EyvyHdEVhOBN+8NSd9p/sS/xZloRK04pAJagobGjtNrWUfYSkF5dHwnPcg
Jafyt3BlY2xOThPHQJk6i+CPE/L41Y4OTpN+cLwLqpnR2aE7fVweFha/8rZYhxgxdjITG+6jXIDi
8FrICn2ebwyd6yAbGQ53elAH1OB1K+fbLUb3NXCNw5KjlBfpERLcwoyXwIcEjHkgSuETzbh2uIfj
ZP/Zm59KUEPyxUYWGy/K3bpoHoAfSOf+QWNBV8Nah2bcdrit71hsm/nb6zUl0RfkR4IrLvTiy3l0
SEQakAZj+m8sx7+rYuyH3JXIBpaR53rK5TAI1Jn1Ogj0cvRgdn4wlWLxstmxBuy4E1R1jcGAK89x
33XVzUNxCP//MV1Gbj2QY5COqueyYmR1IIQBHCrpy80i8OLf57i3BxtoQmFkIbb2R3fpltTkbvZU
VXB6J8zSeVwcOnktwZG1qyDEW8xhsoYCMkEsdtdglMAxBHKKFCid4BeKe9vNixnDj1kXG854nYzE
+r6gdm4/Xp3sPjCGiqKYsTr8riOkOzLTX8orkTLGkfxMHzxoQMZkwAYUBv8BHPI5b4Wk6NJGlvjo
cyV/78VNnQVQ+1L1Yo+IZBX+YGfUmTT1Xym1CwgcaXjjGXaWLTved+wkPtfObPxo3dWHRqOk/zsE
2GesEr8NNQu6PHuOyRRSBMelH0IOZ+MlX82BGsWy0GlxGPYne9xj7x+c6Z3T/Qt7NUvNNcdAH1js
9tVE35sHbUZec5+hEmQsCN5s8XE9AYD9FLPsDPynHMpEdJrs/LfIRwF+zR9rqHQo+xHxP2WMEHZb
jUWR5iERTb/54TzW2aPPi3CD2W9tuuRduQSAzpuWLFaY5zSutYXVAYjT2E+JMjmVkxtoGVF8QaJQ
Sbwi3Pr0y45/7lmddQLu6lPbykxMsCobTZHOHXAv1ckh5lANfPpRCHVzO2VfR5P2jIAApxTK2YZo
yzxsmFw0O7LWqfEesmMXmWJ0GOztiQzktH0Vkglu5MkQEu1vcjLCKnK0MyKnplEtX/y/SNmz9Rr7
WSZsWgl/mIEtCa/wreAA2Xvn7G7lhTzk2g7oCGuZWlBkEGe184dvlo+EOC/1XzYM7btEq0rFxCqN
/gREB7hs31ztXY+2APK9TEUuPWZfBhjpia1tF2oN4/OxvupiYKG99U6szTOgsPUDhStLKqdAHEAa
7MkjBgbYBeNp1NIG0S2ola/enM8PPbe+R4HgSaMadwloMwXm5D51B06TDi59XDD46TySzWV2a4qT
oPU9I3K5Nfd9rDJ7b/SazBWn29HHQa81u43WKCHqyFDq37Qz7CSXaP96pVWAERa26BNdeQ94/iIX
TqqCUtcVDpnc3t140AeYNzxRiMaldYF20vLTtqRES2kTJVqQclgzGCtkDVQHs+938wmoyHV+1EpQ
pQ9qTRBZ4JVGAKaClKAMQx/5mZDftsREan1EloFBWGLJC+6xDHsnQGTYP/tQ0hGODx0D+VlWQdDK
CuQlSpO/G4MJXQ1SkHuCqMheu0rJMNEKN+XU7QftiFSRnRYgO8lERHaze6jnPgXcVdxNQBTPe1Fr
Q/vPC3jZShXxySMCDW7H5nR575vqW6LYM0GEVCeE+9HMW4BXyzL0i4p6MUKM4T8FKGqdC9RphlZZ
sos1+Ylbwlm2lc6q91FsI8u5cOJuZA4wWYQqQP8opyZqZgz+ADxiRIYgbhvyxWv1HElcrPv0Hr6v
A0wDd+WxV/cMusMMBYJ7q6DdYbGMmAc+6YJiPoGVrYZsPQUH9NDSgreIsIBo7qIALMfXlvrcr81g
55E5Rwq9r1o7GG7BKY4Yxlfux+SxCjOgvkca7uertSeBr7PKuqye1sCcK4F7w7+rhRuolc2DSaym
K/QuIG2QOusJGvJWeQB4QlljRP07YXoplgHfCOuZCYusSyNfnPuilxogWoKy9PwgHgitsBaThyyd
P/Ii7iVrd0brpo1JZT8ERuxituJAa4BMfHuf6hyg1JPpdmOI51U9Sup5vetfYOwek8wme1+lOrgj
zHsmYESPSIiI66hIB1Bf7Asrc8ImxXllGB5ahQHo5rgNs2aavc0F4rULxldOjHzT1CFtJKvehA5x
amka41YZA9Sbr9zzc7MAiGJfh4Wtd/34Ka+RGCAIGekBhh84R3kMiC1ZupFrrbCh1DX1y9NFVvIg
4PMSMTUE29fHiPrkeORH4GlUAVdSb+a0PA3yupPLZo8CUDuNIKahni2YJLDUPk61wVNIB6ow5WMK
ByBhjKPK+ZhEmL9hf6QMrXPw5uImNdwq4iSeqBC63orU+1HrYp+KioRTrg/UtMYN9RkxYVPtu81G
uHxadiZyNzP1gBn6As23539YE5Kf31PyNhOLWW1FJ9UIPUJ9sGiLIKyZcVONHXZf/svGqzaKwPey
eOfpvN6ZZlfPmf4DcYbZ6NbBQuPD7hiFX4MsMHHfQYrzfSI9mh1kmRpLLF37cezHHWRg1I2WyMwv
ocpHC+ssS0me5Y8gEomj3H4lRPhVixLtxi91PoRusPuQ/t16/ovf7JmMvlSTD8ukyAKGz9vnyD+H
uSsQuoSw2/FDbS/KqdFYKBbQ7vn2Ch1stDyM94e3sfNRp2zHnnQPXIhMgKdX8LPBDJtQ6zyZtA7y
x/dqUDlFwRuQnlrspihm7yO+kiP1aDYYRbX/Pg6ZbiSoJDpEreCRZGDCfZb4rgaZzkwOR4LE/tLN
yDlRaoS2rXsxvEj7V1VqDRbm1J5QD5wPX7LBr3LrOskkBIvI0kHKtA9lnR5QV7aLI+ecCx+HKxxM
3IL34VldiHt8kJd6PpozG1jzKilPa8ABKENrgT6MZNAExLWSx94qpzSm3AsrjmvO9/Ljtc+G0Qvi
P0zYngqLfikNv0kBfGOQm/Guq8be8RZoeD8a9qF2V33LKOhKJiTDkYSlqLFCwwe8g3gmDxLLkI5A
tQBNDMI8GUKLnLeODi4U7lZTDkCgBf35ElH58Q2Mwjm85FwwKKaucTNyopdvmM7ASNmPeWy7zsXN
M6Edv5UxP0h6Ha38DKsj3PcNG4X+PZes8vFHEzUhoYpdTERL9cp3VEYrLNe+kxlfslEYWu0n2gBm
rxWLqVWA67/kWpVvttQNSgmsaSJ+PkT+6ivV3tssWQ8o0zrZkN0AJJZw70sBAF4Qv5LbtbBArexE
B5JMYDnG8nYd290xEvGjGoCD1XNkLed3vmXmyTNuZ6xVeg38ScpjqdNfyvcK/KlppnXkWE4FRz7y
SuJG6U0yjGEJKnPGZ8Ynda3K+0uOsVdwTGTD0ZNKRATCtG8ei770IxebZhjjRQe4dhUUp7y/ceyc
aClIKlA1uLnK5sIIXuUqapRe8gLw9NeCd0Xn6trpHO2U/9bKw4Xp4ICY84UY8qTm2ciuZF+smxFZ
bsSZ2nPgsKlhaDcUC8aXb7ybhRkxE61FX5pXXmbuvhb1g8v7zO/XYq23PHXEcJbkJZTzVRxX2k9S
f054msSO0uMFX6ixEX1T4Jf8NdX+MJY4So2+IxTzab5UMbd+sn3uGu5DmAXICU8bJwB0KKnEz5Fk
lQ4K7s4VxjnM+o0I/l13KUnFILfziT/zRgZvfOr6NeNhowduLLSYPP7fW5BefocOJ/H7IS0pJo1e
9kxhevmcOgWVSoUam+CWknZf1WzRsjbIzcFa3gUYf8Vev+ikV8x35h3z52bzhSW7+3D8gwDWCT/F
zoZXsRRUMXPwDkNkwIhPVF1yQiLa7J7qprgEqlZzh9fgtzFSoT8rWcQWrZPe/U4CMAijFebejLJQ
texl5M8+yozsqnT5F4CvQKzBzs2zQO5ddBh4Vr6RUUkczWLIVIEQjhw6ggJi439naZHiwQ+0gK05
xjOM9dap52hlWk65G3RmuyMoLwoyR49z4Txh6/4N5XEqBU0iLcoS1XOioaGvLCPIEfZO4VegkbYh
XKjQForTbHhhRLHQe0Ix6yNHsCXktr3HrBXeT9yXU4T0LFskCoJbKQ/4bqk/+1zyiGOQrSQvQ23J
c6WBoCNn4fvzxNQYBNx18DE0SXpgeb/SWOA20N65s4UNGG5NoiQAnUj349W2fUjN9tTGeQm1rNs2
KmJ6A3djp1AjZC6poeAt2S1ZKhPFyAW4I3nEED7uxfI5tOajCXrXvqauxU1LJ549dUoHz++zcVd7
9rfNaXFqcsjpXDoY7HeVVgCeiVnN9n9jijQQnLn/VVYnr8cYGPqp9SYhYWuFdVdgMUqpjRm1gu7b
loE7v828quvbsVv6PFX0y2OOmN5l95jd8iLdK4pQIgIAssEdfXzhwKb7KuGYxNBBsNvBWmdjnKfn
CEs50qzPWw1X6L339nhI2eX0WrQg5cvkRkpE+BTmqjsUkBXK5mJxD/IhccZESBCDM4c10+XXXo8t
8fcZK4cJj+KlDsaXQ3V8wz1VOXNHHyLyJ1OzB4kGU227ah+8/T4ysDYlzhSs3rflhGlFgqIx2bgH
ipY5HdndW5sdIa5ifF6zXRtYzfU0bRAZVeLnVO5Ybjt3/i7ETeyawyFHgwKh9uR8lItVUoOK25qs
wI5pLaqZfa+Bu5CMZWC1H1f0YgaUdcgu6U9JqR2iAF9WTZDTEvp9USvRPC5ce3TXL1i+Ci/Itsiq
Wkai5Sh+57iuZT2Mojb41heLAGqUlxFb/ynFkE8TTsh9/t1rzonNlxZ8EvCSR0hYL0QEJg11z/+I
B6yuwlhx08XjsszpbKiqT/4OLRGHp1A6PdSn615rUqXQLxspyhKEA0qe9O8jz1fwKgM70bg0rUek
rCY1Y4+KpZwYIJOLINvuV87HkViWXA6yhRVVegFLr/PcUYC/5oVCGFf5rimpnZZ18ZdWZUeKBnYN
b4Qr5Tlkje916NyE8Vw/BsKByErmJdYsNOsDv4ys2+xxEEUu80omiLvj+JSVvJ3hf1j14wk0cPNr
GnUlqPzkSMWuH8rf0G1IIvaWYo+9Xr4XodrfA/UPsjWsv58246EnDaRaOsSawHqX9w5l+vG6HkU8
MkwBUpRFb2OmzAo/DhjSzar22bcrLhzoA1nxZDIzM5H3B6JQL1bemA+xRtc7xoOtcjr7CGOUxLOg
3x6D7M7gAYUe4AlTiUoqp3055wT4jPXClhNbOxyHjhrvzUcr9zwmHzy7kz2wRYwIQHPwTBB2XcaK
oFWj4c41fAdyK/3kUOFrrs6+35OGd9zqlDnLQDbneNdSlGUyiOmM/6M4VJlOCJgsNIunRmZPXCmZ
bfcbspPd/DsrZ0YUMGaPY51SCmUERoGxzm2Q5iYvsZw+n+2CPZct3dXM9Zgj74gX7SUIl8UWxL7q
as8dnYkiuH0YqjQxCagBWZpG7U0PCtJ1S+PM/1aatiSscqOn1FVsULFb+nL8R+vXREF0DTrM0xCG
3FaU/Ubgo6jcFi5LQuQUjkmhXZ4ESab8LAMJ9EjjI2zmkY+1//ZzQVJb/JGUS2HYM9tdIDtLXjN7
/RgWpx0monHfza8vbwpqlg8yInUERX+A4aNxhIB0JkDNG4PuuyvZ6t7hxmDjli0yUdHypntpgPQX
75dWqNqbbWztrt31AHkGsK3QiShRMHvVdTID49Vdu3oM4V5PjlujX29dMfBBfpCLesvpV0X6htCH
EmAubVIxZFKsB/6p4IEtHtRJ4VduRkJVU7ZJevyjf1L7QR4k9LD8E1otp6AYMZhrxpRhFsqRclsp
Jj1UVvlV/xJ1IqUnEkTTdGS3go+EzE87wJpxd1ON7C3w2p4nRBRi92SXbNomEmYm+rlUfQU6M4s7
fFsigyK3clu4fhqOhnrWzJznEDucQl1yW7JRcesCpnaBxtL6g7R82lrOWW2EDVDxRVLBs59V2b3u
fXHNY2j6iQkqyDVJOQCE6QgHJq9rIMkh5mY9BCsTx/H5J60GAAr23NqUs50AydmSRpAKvwMl8vIJ
uRuP8OZRgYdyRh8SKI7jsJ/VZ+WJIPA87pqU2DDrv5S+Z+Gebl3N0sYeV/AkgQEYpjsZz1zKtMgD
2pEcyPF4yRbhEHGXQN3yVu/7mXEu+r752Sj/5CSGcRqnDZUjvYmGil3IieCbb22htYMfiZiCFLgh
px5VZPOcLcXfNGLECrWE7nEkmLovuDjIqUTJgd5R9hZLFRO8Y6r1xo+27tbrFX2AYZy+9/VSEi3g
VT4OtF9AAcQQda28GIxxOzBy8N0GI7KD8QO3DhbdQjsh0oExCLv+8T35W/esmGzdMxlbhd2mVVAK
4mx5BE39vWut0tHf1pMHbrA/ez0AdF91uIaRscZpqJXEEbc2v1uQOBTIyd4Ex4/KpweEd6HcOECA
PqyZUt+/QkXUSu4I9d3p/sQsOYA6mJFUhVYzqP1TvRWkx0iy/vqrvye+5eLngtN3K0tw3rk3ZHqV
OzyzlvxD2Uhs3uf2RzZpSMKjG4fDyQWE7yZhMu7hDa+tDXwZW4KmQV1eFxhf1TAuEQy1DSvhJw7x
fQRbwjEBJE6uSGjngCv70yXST78AkJdSfLAHvMkSItJ04yv3Wpl8juIOo6z81AkF9KqWzfFOiugT
qAd+IzcMnrItvreChCkN21gys8BAaGTO2n81Z7oZtDBLN64FjEbVhlYrbeovSvADkO+I9lJGUidX
YT7vRLPEeUnpnj5nNP2UJWKvyWjFhyZmZRKofhGwDp1AQVlC+UT8I6jT2LIYTcKxrFdF7O22SiE5
3h0PltbyXHEt3EQL8pP4Vm8aUce73Y86uH0ArPmD9W+O1MUC6AtbL+NRzW63fOjeOGqEt0MSHyMr
cj4+RTJLYitXtb1vFnIBflUDU0KBMNSJzmMFXpY5qlGSHrkqZEuQuWFCyVfAqWrCa3LRK200qzM5
ToDrQdRoEEwCGmjvzjB7rXac0YNGtoJHetasbDzWZBznxVu5+0LdqXWoDxcBNpLf77ZoUf2PIJeR
4AlaEW1lALQJFECLU4zanfbFRD13cffu2idMQVmTbg3LO0o35jTYGFSHaQuFki0TAQRQs9lQlLk9
Oa3nOOmNQiAwKbRaKP4AFtAr6vjgh5brxmb+kLGFDDknnrC10Z1r05UzY3sEem0n5ZVnpXYtCt/B
i3AfKQdEshcDmJGC8YG0twJva4elJYOYy2SX4axkFLpb6AloiQZbPRHtAdrvHVfnVCo6ei7a8heI
HJz8eldc4Nzq/nOHgGOc4HDwhn9UOUsfvlT54j9bddXKrrJMdzO2q5DIdRbsUai5G1267vc8g0Gc
3HGRv0yJCO9CDtojDkXZa0E11fpeJcY5itbRCgzPtxoBp0TO2a8y/veh5LUCREyZCpKp5+3khS0W
Hyi1+zaay604bOqBAdaMMwmb2UbyxbyUCHpiM3JY8fk0k18Zf4P+/ROMdsL0PrQjIhrlwS7jcfjg
5FdPGxqqOe2vYoDWVQKfnOYSyPm7K5NxzbDy0ESpTWN27vBO+Rnr7ltPw/IMVwKlCFNtFPR3er41
9KcmxCr72z5fCGeCvClJLko9SfFpEa0/AL9pcMYW19lQvaiguswTYLzSevvSQ8mlDSWb6sSw0sTH
FgO7MCjL92Kk0498G/Yo7pYOjDazXTBHeDQM2//56OPo+tf5j40HQB7ckNZVNgMQtFUUObdD/ZRO
mmJ0OGZaCMX088fmHKTdO5DM1g/048eCtJB9Kk5p5rNKYobYyw0PkhGUElrceMeqKdJXabRtCixl
qNBmu3+JqHYlTwkU2q7qO1pb9eW3Yxyq3jxbFmqiWA6vy/rFyjLQnFYowVI9uD8hGVZggihBcXSq
q90EtngwFIj5qculGGQk/b1eIvJKDcYzjeerDrs2kDsMJpKgbAr2Li2AFIvj6aqTGZuKbTpnjfAn
18PTkOaC7d3E86aBc9vhbdgtiwWf1EY+/IjIrAHbEpIqPFcNbIvWSPt9VLAtkoMaxw3GMtUAdRUo
Zhx9tfBUwHdDRh5X3NwmSSVWtO9px1LnNYxFa/KWGQbEZ1G/Nhx/Tg9NE63+JzmNJjMI7XPcbIIf
pj2jOw8F4vZCp8AH91cnTNAllrP0mPanrVZNr9aebv5i4YzoCmq8/b4K5jh+E2rfHEnPs0hL2Uwk
SeugzkRiJcgIZ8DXpxIgdUrHh2KdbvrR8B6grud0oQAkLuNUpaEt/hzoManfLyfzGEdxmhHwedjs
ZIXW9secyaIftgiYh9uHEzcucr2sYDUCgRA+JS8ZYmxYtkBW803aItzAEZAFSxvuV4Mz7FyOBtQj
xuy+ix7UCWsdoMElofeE2P35chPYNryZwG4vBF5lydX3n0Z6z7L9qJevlCdrqowqOkzbZ5irFtGw
YkcmRCt+sz1g9H3nUlaD5otyLeakKFfxpkSOmx6EYL/8fMKGnprlR3hiapf+wD1UhwPoLvyhD1lz
T2xyu7ps7OL7Rlu5XD91ckVeee8GqxcxvZGepEnYiv5CwdVWuF+0uegVyarI/2JZzmJXfNffmbSX
rJrOmMcAHNTVdRP46y5Yo6zbr8TgeGbi+rL/vG6pVOX31gBOCqrpqIMWMsjtRdAbNil0OIrAJ2mF
gWd4ql4wePdfEloid9ra7r2GWoOS7Dbjp/TFF+yTIi85jbQto8ljfFeu69dI3BapJqgaiqCuAyON
iVNxjIghXjY8sOYlUy3koBBzdsKv/I4uUZ0v81YsOY+T/gV4pMtApaaWNJX2hozcrRHQgoDAdrhl
J3wQqJknPTvmN911B/uzfSGb4JSYsy9NCHXkTnwRo3tvcOpNC1VjNkLgfVtv/IKW22xwlTKldYkn
SoBH3RB7GkEvfCtwAk+VdY9EuSmEJHCYzZOzsbp+5vKbt3pzo12801/rxeEtPm6LswAucgimzkwI
YIrtWqWdl2mWssjk6GeMlLmHO8yc7czfHRNYML/FfTN+hZi7hgs2eTxdN4fZXrlZLcXnF9GWLn1Y
XEZFMRQbCnoMvClicO/RT18g4ffp72TF66D5ncvynkFgz+ZWoN/XK0uW8w+3yxwuPIq72JcGDA9u
6Xg5e2hyPO5j17o3Oji50KuSBb0gAISN9ntbtxuHw9eyZSaXi3X7+3LLjQEwr2PdGIamfLsJE0OZ
Lj9UZE0iZeDfKTBPJZrHNhNJW1bl2nt/FOLubaplxcLT9K/QYaOnoHO7oYOI7dCUmgvBiON/8/fG
VpTrdpM46+5cC+zOM3fk4u8mfWLhKFpVSlGLT+RQlT20p/J8WrQxmgxR4ad61leGskeepOH5T8l6
EjNNaJ0VfZdhAKJkpzx3r2kO5MiH+ya/ogU7VF33UxIqVPdoR447nQtm8z0OWNejaNf3eIcZ2U68
OrbVFgdyNcVEf1X58QQCaIR80cXm4ashr/H2ehYI/A4Hi6mlA9JL7gkcgGgPksgX/2GALKpv/Pv1
BC5U+S0WPfRFaT0lfCrl0GxUSjMjG0mK7axL68D7mBOHUXyMk/Jz4Tq7Mh2FMFNH7H1l1yNwJnkv
xyMEL+bDmD0ZagAo491oLuMU6L05kTdPBMzee456EnA9zJ+OI/3GwIi72DR4H4rAVGdtYv9UMKmz
kf0vUUTqX0rpO8OjXFp5p/CSrMccJGSFgVW4Iqi5ByPmDjlE+bYjLgJ9oYwRLt79jEkz6p+3jDLi
RWs8Wkth+f6MkWWKZm2Y0Ik1TffFcIm9ZGvQ+JyXgS3VJT353qD6jKZUegWjJsFV2XGqN6oToPFi
2SdtD6R+1jhNkuQbr/NrelbcFTjf0PpNwhh9KoG0v17DXrB7FHJolpQOdBbiXdovZTmNtmOJjKwq
03ood3+09YdbTzgukH+tx+UaQBbEwiqrE5aJ2btV/BZAmh8hOjmB3TloRZLiTBJyXPInW/iwWudb
G9hxs5PWYt/wm783PXukcj6DHo0MPAlBxcOyUtuDj+2MIQXd0F22h0fBCG9Fg/k+0IO2HpipQqKm
+rQjbHfLTy3T8fiNCHl+u3+erpHkqj7IA/knnkbItLVfXMhwAQZCLSI40QPvbnpprt1EnlMtoMHZ
JVturlD5FaV9aINn5slntCvYiBstAItoyccQVhg5dQrzXv6XNCzDqtAvO9E2bYFCtzXQvUFEZ6+b
aIP3VR1PvSjiwhxOa1FR1GWlLFBqLKt3skEePdCnd69yaJXiYd+tBOCgedyF8OveTygFwyrSqQyx
qWosnqIIP8rkrfvM5u2etf/yVeJMDpxQXROntVJTFUlyWPmsoWqweHoICTY7qUCpipKS4Nvsolzt
ZFZy8yLnb+cu0XJfOwz6qCEYjNBOuwXiO1LBkeRCrA9+v1v2fLAlft/yTjC7SO9pxJZI006MyEdr
9JE1/FmRuwZDVvC8S9O2xI7Ny0H8TfSngd4V8a3pVNEZdVy88FuOqf3jv+R8KCE4w0s5S2qTYs0A
Nsr8hsRJN3woHIJi09eipNQoXJjGlP0c/oxtqGSCmsHqsIvfjWKuJrbcaDFWA04cuUfVLNQXz1NR
1/n3WWsGQlmuZshCMGGPIw7tmHng9uiSvZ0J/0ThVW++IVm8pbYr+Ah3NHXp7lQGdZKvHrT7WCrp
LQZoTWRur82s5kTDnIpiTgKWx44phXeN4CjEETp/f1T942RHTRQXi+SVtxjT4a9grF3CNYgnCZ/8
TeV7GSyAfCBcihLDBZLDjFr7k0MkqmatMfEaZ7AVgHR3MPfLm3T119Eg3PbgE4Hwc07OKbQxNfLT
X0NkpEH8nvaMvQbfue4RLDNMLSfQyYZb0I15gWqqcyMjIfWhvusIO+B+0bA02RYzQgUH43s42F5b
zPJz3jsSHP6M1SE0iatHqfG4DSqeSTkUdPezAD6/M1T/Kpe62eB8BZ3Dc4V1uHEa/gniaqkzo3XI
EjUMH/PdNo/psqN3M3HmsogaSfVkdrRoL0Og5xHbPjh8iRsF5Z77KELrP0yLsyZFtO/VJ4wnRoUK
4XPf2J7ukbqij/CMFHujb/QRh6tjQl7dZTIXqPP1urUZo4vQQjC1N2lIYSk+nXagmUtujSowO6uu
/YRxQ+tdc4IGtK+VPbkL3/gFiZO5XwT09obR0OG7SoDr7loQTGFR7kWV765B5p0tr78QdV//ETPT
kgASiyn4koMnTsoPVBO+EmlO4wtpQx+v2sVv5wwk5gy4dVlydlWGGMr7ILR85EMBCz436HOkCR10
mKaqHTep92UsGh2EZ25umnWgWfFxBUNAZv3LLyKWNvF2EAZibRHDlY9cOPW9aOKp1XJefdjpd+6m
ujzQTPdE/ZYcz5FO97V2ld0bPBgoH2eazoZ6u0PYi33lq+2O9+KzaOUbTHlEkXbtAyAxCVNYXij3
A180ZksBQT2HKqM859qCu5s10VOUjBQZy6ZlmrdZE1bPRAaZSbiUjCgKnknj1O6TkjZN3J9SXqr5
ZtzQ1VXvZijnAKvw6UrABEMNvim6DNiqV/yYD2LxuWxm95CM4I0Yv9jjOmUGtq6k8YqoeMemaXuF
+Z/j9IgLC2vrVy9emCDCa0kUb6om0vxgWZSE0LYU2bo0PYtDRyIFSLDmnKu+ESzbAS0sFjKPgVrR
zhwDO05Esf76wSMNX8Mra1AEQZyOcKy6T9q9YDSyYAZih4I9U4T1FFAC+UWX8kMLb4F5qDvEH2hY
mHs5VXiyC4y+rR4ccjAoyi1l+Aoa+8DwL/kWmOOOk85+4QwQkXFFjgvdxwoshZp/CLOEIAGqF6zW
CsP1cp5oAPWIjU4/eLmAdvI31XqoDDRXK+e7++Bf7Dr0GP6GAeG5bAaqrsmBCeoyFtumOU6FDm/L
z1hjxrkoBy32yNrtZT5pO/GLif6Pir1mZW0lPGeqSDY7LBTjaFzZSARgaSq5U72YIuMytXoQSXzC
lzIvvBHNarm96On1XVJN1UCUSbbapEk8HSs2AdtdHX/WuPMbphBlDCWal40rAxpwVhQPtSRn+eI4
rT129cztf36v43XLHgbb590avSMNjCap3MobrEZ4jw5wnFfO5xFKfR3anPG0AxrcyXODZrBeV3Qc
JTePoJrMVRAQOxm0TK5LSxSFAjm5xP5bOzVCP443MQl5rGSLNshDyyPgutgkBu0Yxf5dLxF9ZdG/
0vGVGvnEzDLF2B+nEOaaX3423ORdwZehguu/59hF5u35LYuQIJ1bFDUQ2rfN2p4g2oLiytH6zmzC
rPr0jRjNCfpPse2MA5vNXjJtpcEF9x4NXiDUtBAzaE4xOxAHYHUGqOVUlrne+iSGHI6OOfppImfq
4ZDzMVdIWPLbvyinzXM8aKxclV4JN7mbTuwrt7Vpffbi8uJ/gtjbNPjtNleu5sAL1CHnxpkb/OBq
Pu8qjGRpVlvoanbgZmBsoBNbii+rXsa0o481xIEHthc3MyoJZ/ZF77Tb6dQxmPspNsCS+3dU0G7Q
Gykxa/dlpjsbwOkjXGE9NRfBtQdkMDc7lDgUbOnLvSk7VFIbAly84TvBgroPe3kqaLg8hxaGdMN3
DmV9qa4SM4hsbDgz/kKnt3r56lNWr+nOy8FQGQZubTeM8ySBQol06clABN5L1w8NEWcAWEJPTkLT
F0esHWccpTSMASHQpO9l6OwEO8TkgfVd4WIHv/w3N4zhH90taUo0jkDO21jk+/ZdcRoooaP+BuCO
3j4ddTsOCnW0UMF0a679k29iB6I1AOnIm56tfCwFL/7rpUGsf7+3Y3IL2Rf4QMOhSW6fEZfAXGSv
QsWHrrLyAq4f/LbERLPC5N6RQpKsc9WRtRmKtbEvZkzaCIqdY5E+ul213bgfpCqwgB4YXZfZHyQy
s+GZfgS6uLgznyv5Tfwd0hf5VT6MmSt57OzInxPNONxfXmEnVC94vOzqqSaJ0/PkzElxeudmJV0I
VpJ7o4b4zYMrdQbCZ8tUk25w+FZovCymofEUsyyvnHWYWW/gVFd1ExqcO0RqXcSLR1cxcxe8Junp
JLJ1OrgOrwnhBhqVaxTUXLEIx0vzcvI4p2GRiIiD8YPthE6y7SFvE8hivO1VgRZPJR6izVLLWJ+A
jglxegnWOUUdVIjQZt6BiBerdoX8oRH2ftJlKsC22cBA+CquF/dwDYbiryuvwNkr9dR298cQwSMe
Fxcy+2uroELke7Zv7Xi2ZjauyBPrAIDXspE/S5ywKaImK9vNUOc69viqcwsL+ehn93kTtas3XvCQ
XKFwpW+z4nhdD5nGDIK5IItB3OGhTqKzf9OgmNGiWUwLbQIR6otWUAEBMiU3S1Cl/5z/kP4R7l5O
T5QimiY2nHaqYGPLhbgjClQrFtWLTfvQ8M3F4h1eJMMGWkmxBDOjxN+33K3+cLm2erO6gU1Y1P/9
7LijrmbI/Ly4yJ7Ll4q4TU0pVW2Noccc7NsWrl38OBuk8mVbCmKYzUIzT+37lgI9QmcCuK7xKJrC
1hiOHjwMyqhPaXed/VJKDsfyBdjtax4kN/E2gQfwQ7Kq60FoMyVlVcN/PNSFQ2aYEaFJdakOZq5l
1lZfLqzI6bDtODLr6i54os+nQfFPsO7rkPia7HNe9l4tT/0flPoKGeKDkAmx4EfOc/6KawT1Nhhm
Fv4ApU5u+8mANY5rUt51Q/+fS3SgT6DbkiylOxWHiKQ/oxkeYFE2sqBX5cOzgDsMyRnBd/+7t0SF
txO6a5ZaWhf3QkeEoCqd+jWV18MkhFmzRL8+/Je/dOzGJpnP+QXNNP4/Ajliwcbswqe8cvfy8KtM
t+rqRNto4xIyAfCkTU3SXRM7cOrvOmScZXcUxTekGLYzlzL7M/yQinZ6hqtEtTJvlhTUbX1IoT7j
+PmpSkcjBHgnI8Yk2EyA+EYNMFZs3HrENigX20S3glrrrs6YGD6cUn2YS21+hZgpe9YX/gfnwxtN
7AtpEgUqML4t+lwr89JuZQCEblKCYtUZlHB04ySpeTuf5/J6TU2dVjmD4KZZAhBTvTgli8/32syZ
1go8Pe7e0gUHwTMCpwjO6F7ZsDfB02e1DIBSiXuA1TmZenZRHUhfH9k+rqax/a5y1kE4iiQ4wVcz
buRtOzDvWjCiJWRkLYqHYzsDQobpsjyjax5/soSbIIcF4l2gvSv7JUcuQfedS4LFj5mV+JF6eiGC
qU7CCMiZpScYJ/LLWV+tr/zxiW5kftlbfcL6fR0jivzzWT9JZJyiEFZ/NxDGy3SpPY5skUCBYZFb
afKOXklNNoi7N15OD2njhW3dRbzjhiyZpVGaeNwCVxWDSG1s3TJNsjQ/vrOS62PfNC1dfeUPV4k2
vC9Sxc+VKiV5JEwQrxssBgVKVdopRl1yyZXWilQ2UwhYk3eNtaqcQ74FkAQK3HFDyilQOrvHla5k
R3k7Y4uv6KCwMLUOz0ECtXb/3UHciJAPOK5VQLBHQEKR+bCnBTI1k+HcCcMu7OW95YD16fazVYBT
3dyzKpUChXbqU42ll74bCahXKdPmK2HQWSsc5vFBXSKQydsFoeS1FP4gaTjbTkRxnEjsw62UAByF
FVUEsJKKe6J+NfyqA8k7YbQ25ljcC1zT4/LVtNYCoTTPSUp3hsUvTjecdqiGSQkDktPTFI4/RlnB
JVjMTL05hezsqJG/qE2aV63xbh/mtV585WcLROsH13GGP+Kgk70gsLL//XPSJbqaKZqFIbZV+z7Z
sM33K54I0XwbJKy81vIcqcfDzXaurO9xEtS7qxPhB1kbM/Z8Ca34K1kIDToY7S77+iUdASKU06r3
B7MyhiJ2V+fsGUNkkLP/hhGJKPjuvBq/wekmjOaWTaDOmP5fahMXbdFf2FmpXrvOOvbguBJOR7jG
IaU/urdjkQ+nm3fa6WIfcX0ilFAcTALjRbHhS243kPOScOEuLgIAdF5TZ6sDE/Gvj7sqyzysSk9H
zpK25zOpBJCNfAbCmzPIvDiLe+huY9XfSWylw7Rb2sl6lyK7iZlPJVzwcD/JjxKXLI9gLPCN16JR
GdhE7BEulk1zzsYb5lID68Wim1zdk1uSptmuykgt/QFSXZiRRtMh8yVgg1pDsvNYGbxneuQnRJwB
QXPFULH+d/WrIl9TWoWi16UPBckCvTdXJ1McYa+jgAyzdWXm64a7mMihfOGeAGQEUI0bDxNc4P9c
hOGun/tjk3Dq8hL55uL3bdoTc38o2HANQlllUURggRdHNUoWw4yFolUCk72YDuj9aGVwGw7GvOQb
ithS2m8nPCu3iUGSj2TuN1LntrqZgHbYVW4sOLi31275JnILZXRqHqvGoYUT5Xnp9iVLohinQC17
EyE96vyqvY3SHK/HEudJabzwzooh2yKoFaIlR1/KhwzSBxBwnWeFBaM9Mf/jMBHV0q1nHVtl+tgO
6RekEV42W1/G0uHyXF2qksz0cID3R1uNMfTFHiub0sjF8CHTyBwieuzIvFlf388f1N85z3TEnUey
dyb7FpSIrct8Nogco9PrshIOKLp+nkPhbC2gk0aJ0OR65OKmB6atr+3nxQjRM/CD42KmTcHbH3c5
f16BYS8G6yo/qHlwbMY+Y6YmrvbbWAC6eXoUC+g3Z2E54qPW2GZfO10MtyAMJngjzfD0N8aFBhDe
2nqP3xNpuSzf7b48tVvT/x/HFCE1CpWM2tnQNH4rn6HAvchz8R4qLdvrjJpcKJDg31xFCXlU31i1
2xpMhkKgQkCalN7lR3Obn/r4XubziWFSQHD973UaCHeRxUx/aasg2kq/oNowUo5MghDtB3adgZLz
Ht/I89jN3oJnt0lnE7dPFXuJJM27CvQobXBvIJB5vs7YCMm2x6No01gNdL/SyQTjzD0ICjS33ZBB
VXeA/K84KHpOn1XaR9syGdbFwY8Un+CY2Ke7wKmAhSj/5R7s4hzsUX8R/Xjl/8zli+FvNS+dpVxX
4IPFeLElBril738oItqNKy2bYmQAXwhUj82UkY2PIcvnHjBkNUOB1dfezIxIMFmypiBEM3MYLDYQ
e5Oa0w5MMidRVeu6HOTp1+YB0m8KzJwedkypNyJPsXfnETtMMwULj2nVa+ceQcM7dK3iEVPhXlpy
tubY9aUX+wTbpBS+Lte2r2UT23NzRuLSSTLP+VUZ6+1jsk4+Ex46akkdVcsSM5eJX+xOKTh4fbBi
EfaxWBHtl0EaTKazox6Pbjr3vjLmPKPugNG0aYZFxy9D00JWSBV6wGV+Ayg0ahaY0gwSar2nzcJN
brkMfQMgWpf8A6hbuy1EnHyCPNGWvDLYAt0wTcKtulVUEoOz0agOq4cDHGkD3T2eWi9FWFCJ7mru
aZkkafHVtrus7CmT2a5mo+IpXJHeFa5iEwsHZuktJmdaDVRCu6cAB7mRIzRiDOul3WDwVK5qqBXk
UD76u+neRBZo24pL+KNCH/20vgr4mAjIv3Tg3hP54xN9NhEGt216U+pRI1QaGcchBiILjXy3pyfB
Kt9T98JWD2dtbcLnwvgChjBxwaaUV3angdVu4OH91WVddy5xCHR0mbMcckPVf1oCaSvU4yi8wkPf
EkhXyvCoDJcyPgMlfQ5ga/uhWqqEsU2dLUs5UqL8aUpavEOyqVzPelF98l5d2znsi/PJvhOZTDrn
PCDexsWDiPdntlxNCncvX3rkyjZOIa9NFbWM4W3ZYYhmo4kWkbq91nFtAQgH93uiJSLMVHOCN6Bw
aaRqq5MqMjvM7TpVNbC1BSWdbbHwZJs+OYXN+32TERPNPNydBQRaODbsDDe+CbjK2XIAN3NiGAnt
t97dcPFSFvcUakCAlBTCuyEW0iJGFjVAfiuvSFBfaQnAOajfn/SfeHLatDqf/zrIalKCDDDCglG5
5EWj55mGvcc3zVI9Qe9APot0iF7hxyI/cTMjocLejDZNyYwLPthboUyiTAd0jSfTK50qgxKZptbF
+AKRig63h5qdMeXEyZJmIml6tvfI6bRnOOqtwiKFERtGZ5NbM8qFSJ7TMPY4yvM0ubCH069Df5bc
teLyDitAmOBNTTPuopUBvN5yaZUEUNYfkG46V+GAGxiUxWTRTgXs+xZLBJn9zkLH88Ne9F9eBxFx
dqw7P2EB6BZRogrTcJ9JgJlKvtW1F4+78YWm+FzauXSFi1EgeN6vc2YxaCxssQIzO1m53cSzbQW4
8FJCgnlmHDGCTEkFiohaQV90hNwjwAaQ1sw322fDkH8pS2a4+1qeNzGgnbAUrqmNw3MWLoVQT7LM
cA/+QdniCZS1RARitqjhIe8aIrhuBeuuYsWneNSwb2FsC1p4qEuN8wW4rsf4YWBEC7EOhOR7qZJX
mpZkTJ6NancN/xi+Z3VLoH1MhKW+3en3jfb5qmDqRjDOnQ4Jed5BS1xt49TxL3rnfBlOcSuTGFz5
tg9ZQrtJJnQ3MJbkf7E8Ib2GX3pk2Wf0+F9j89DJL39NXnhi03D5wOhcJh+2vDIjvor1otDuAXUK
T6xJ+xnSA07woyYhmc9FzyUh4FlrTwkhkhC3VJ37uWATo3Pi2HeDAJ/97382sPf+idQ6VGUvu0Tx
/xCEjrQ1625hUO5VvQAb+70DehgxXI0XYQ9+W9Zxsbo6ua0r25yaQDX/syJdyeVhBUCf3M/CEynN
H+6K5nJcSov2ndxIUyGASNPYBI82RzsE//Cm49wAB1dQRzWQ32Du5yNbg7dNcbDB4ju1lU9Qmtrj
VnMN3gQMK5YT6x2foEHyloPH9bIkx+w6W2wS26F9WYhf9GUXTJITUZyVUkOhyFB86ngAaQqoxXG7
iti7tzA6XWttHmEYl7DL17z9z8tMGOCug4Hbb2Rc+pZwyg4czWkRX5Kx9EOyiPAb91fhM0G6rTKE
Z6hYzUshzz3eIqEofiWH1HgIEZkKPbdBqYfVH9lmtw/JsM+4cE5Cc/JlrWFe/Y/jhue6CqeMO44z
gMa01dhid/706vHs1HFs6dCe4FLq59o579Lyt2IurZcy0jS8lOU4T4N1k7e75O9TaZr3CrvJnaiD
ayA2IhjdahEF7oLfv02774mmo1KcrGJssu0MDFw1G4Qn7n2tYIxfM+6qrMX/rYooGp06tgi1XoPk
fOwY+4UmXcgmknZpRWrhAHGGc8sqa81ih6btRgoDrKXv+Bl3gi7np49lcyYxEBCsjZx9gegU8iRZ
aDJxyNZsRUFGTTAn2Lyanl9Z0A6X98aKjaOfA3zpZ4RiYU9qWB2kyOootrIWSsWkyyXkSiqZk/HC
Bh6W/vnEVpWyeWkASj2c4e3ACaZdDAWEzkZWXB0/XewG/6JPmHUhhbx0lQK0QFmcgRzgrCiE4fai
4FNvf1CypPuriks+8rOTB3zlryHJTyoPT/iDawf30U1A9NHbAQNJFmJzjAvej10bnRGoNHDxguFr
hXh2Ci5bu79CXLiwc55ZINvPH053lhFuV5SAUEDcfkvgmgHmN3OHVwlbL093OC96UL3rkylOgZUl
VAMGgdIWUrBSR9yEIzzrv1T3Zq6/Ibd4LWFULvUb3MtZYDhGLXghSgHYrvY4EOlQUX83FnuUoMl5
tLmdCdYrqyqPDQxrVZFP9jH9hi26N/OIhVJCGJKRdrGS6eZoD0HdNGPeqho6VGGJ+Ps4pprp5zz1
I2Lxkm/q1Tk5oQ9Wuj7d0WjCs4O94nURcVPM9hdawu6VGdbR/tlc30Yw7BJZkju+ij3ozyrX/8Y7
febsOS72TCxs7Q881uvIrUkKPjUREoK9h4ccEDv/XHgaY/FKfPTRcGKZTbaGZl2n9IhK4YjwDQrf
5ekVJdDQo3HdHV+sDtlQnTM6/x/uIM5HBflwgzw9zvL0fKCIA+uEdaj8QdAfrt1iRsxODD5zZNJf
Mrlgs0nBY0UVngabCEeghKjWunCpvMcc6zYPxKZ3H+af7BA42qZJF/lro7DjBSnGMj8dyx+x1nkt
zh/z5Jk0HOVK3Pfbu0NAxxFSSC6qWjZYYCpG4MGFafk5tv1JE6Gx3nVPoWdY6WiYbWvou6ibJ1/I
GXSNfNNtI9OKoz3e78GraNy2yqToSxPIUUePgXth4/WzDl4HI4Nz0aNn8PYIZkTCS1T9FA/ocm++
HWxi4M85ENSGhvYgZO5axrhkP/zwGN9LelrHmmuNGn/78O/TWeWdadHx0Xq3rK36A2o/v6CkIwVK
00PJNjyxQvat4BY1Hhxs0G6YanzeuHi1ytcIHHMuYIUUjs2NdQFxYP3AmhvpwUOt1paAw+XXBU4L
NOPDITOiT4S4LSQCmqrQuKKtYpf81k3P6+p0OtyBwglorIjGn9/IFy6AcEeMSZng2TezjVPtLEV5
OZchcvgpWdOjIjMvthNEenCUHfc0GZaEO2fJbvkWBhA/Q4JK6Zl0YCVQp7ZLXbLR7CQ4QYy2/hPX
y+XG60ZGvZqj/YJBy0vtQww1jgz9jGDIBtXHYpJjvjPFta6aawDFmO2oowPI7iYiRsa+Ju/uinZQ
rQxNClu+90eGPT/s9X4iRUevEZ09WVxLfMyapZQMhLJHQCkOVExBVw+o6Eq6NwVzNzzGquNfMKn3
rmy4bX1Zy4uUG8tk/79+XjtEkz/bjwsfKAgaLyzLMysLY+PHBwGHFduBvzIeFyikG4rxREib4pWi
0s5m+P7HGu/fjGtZTl46pDjHBLsmZLap6UzJC5pnb+02mPgO5Yg/JIjs48JobqkS+CwyJHNUuI9E
qIUE1PruztfyTWQJxd+Q6dNtRnzGYiEzoFOR+v3J4PIPTfx63qVf+OaUitGXROqBkT/0O+ypIrYT
I7v6Npxa5vq2NNnBBWi152FJyds5XuuUrHs+nvVAyhyxiMuNI9NHmnXzzB6RoyyP3rx/aptecYk1
xiy9a58NjNlqMFkPw77TgsdL1vcjwDnSWDORxBEgAdwouNj74SNTt11PSG4XjMYJFu3RL+7Th61e
Fn3qLOZIxUgUgzV3MLxVgs6m1RMWgg46W/Duuk1ysB/GDuWSBmWDuZ0S85eCr30lk1etbp4vr4Uw
+HY5R+KXT4zldepiQWuE7bzJP4kCqBTR+VbgcwRrwt8aZCcKGK5zi0xP9qKGkcK6/1UDPfwt8o1B
wm1E6saa9PJ9F1X9uGEps2UuPA1hXG/niQamLxiOMh9PZHftV+02xYSKj3q1N6YW/bROjWJsKcR5
X9j1D4dx9Xvu0Lly0Q7jemn4lHi4pH+QffwSvF4wL0UqITJnOBBy68W5iZqfyAAWsadCd3SYP2Nc
wJmW9xCwr/eO/yJVzZPuj3dDAaVQHIRi5Y+lg0iK9a5gAa7LO9pv6YDq49pibFXI/FRyF7jpVSB1
EKjKdMB02V5RTeRBwyq/Q6Dw3+fgXg68K8jc0RjBCdFpHAWafs4pWiekmFH3ugaocsaQC/UO18Pb
i15oTsHmdS8VKCUVaF0OBh/A/klVPcPyDRgNJGFbZaTXPGHG0y7Iv49uKDNg+V6t8g7GnyUhrzP6
b53g2rdgmerrQxoajmB8ZQ8aU5SWIn0jutFvi+Kv3DUtNpKoJo6xuVPDRR/cA/ftsvHN0p/YnQwr
s7BKcU1HRks3VyrtV0uFEu87Ud6uk2gAv9CFrMnOvURi0OND/BjPOm/jwrGjikJK+g8jGxP+RoAp
PgKmYF5CQOURmKYYkRHhuURFJomRVRWJWl2haptbImnYVbCRdr8J4acs4KqTKaPgkDg5CFRyn+WO
Y/GRroA5nw9FNhFHDYm0ie+Ux6tGNXd/ez/jAkOVAVde/4YM0e+ta1ERci81++rWTKvKGY92MQbR
bEpXiM8QNVdpCwxDyPJDiRrlQai/UpWpsrNztRzBxTrLmbTxKV0bIYe+mwepAK4ShBIfmQKvu9x0
GpxHTXpGuYSBF4TC8ZyTXLMpAk4EhzxcVfXeFYRXQHTYAeebnHpXIPzJSI/3hCsFZnlNSuNULi9Y
sRdyQl5xwCrb00aWEYUEgg1Iqr88HKH/+0Q8LuV3iFB4Oj2le3M8Ept2m385tiRIS+MLKuXkP+vQ
kFChXEGmlZyOHbtQZCtZktRcq9oG2B6e3sM0tIq+uH6WRSwml5TmdMt9pnEeGbVKhQqt91caIYls
x/Lm4TcVlFUQeNVIJMMROtx1FH7ou+pUJog2F8VbCNsCjNlqgIpstP/s3XAy55xNsSiBe6QLpdvw
kFP1x+JGNF6n1uJHBVZ8Ig+jopxvZoOdsmwkj2HcF8HXc+K4zLrbaywZLoFUzKepcu3fWmet1cmh
+7zL9GW8ukKtl60504cYcgW4jZbvOvcw+ddghmftmPik/l8QvMayof7HAnQ267XqVayAaCTB0s+9
YCQtt6zxnuFjDwH3bEefe5tiKdhlG9hgLxeSL2NWwBy5vITVoWQXlHQaNa09L5HRbwhcLw7na7u/
PuvUxNQqtQY7JeOgHLAC9dRLNcs6GogRDuRqnDILTHrCAffga7FF1J/jJtb274+0QbD5z9Y0XQSW
zrN4kLfpQHc4xFVtpRKm2sMweuIBnIC7e6DYcLeRcjqaa+baVdMP36MVuCe167+ql5L0urM4IhIF
V87fZL0EuRWTd4/j2PC9i3J/IlTHPNli98p7Eprmt5kYx00xq2cJIYXqKsGI5THAJwPxzMOTGKmk
d8M8O4sxAQKXEH8G1fWJiRjBWmkEE2w/mw3VFVW1JXKKlWwC2g0Y357/gXdjz3TW6E2jfdVcnJLv
jN/GtEHIyLZ0GkIB08slRl2Zklixdt2HpJl1BYssTBiVAEf/Qx83NHXInWSBaGk+1ckZDmTMx6d5
0y0liGZFYrjqr74gRm4BX8iRYyTyv9XDOvaLkIel/m+Z9lGOL64M/aMGqUzB6kEMMrDnDuAkQ1Bd
sZ6EJbfu2KW+alWZc9KyQRxR5FBXUd8TbMG4U0PogJMVUly+lStnccblDaYYez2zQZoXiwS8k/lF
G7rBqipiaLlqU1QQDlAxdyE6l+5Mra4y+1/mCHUnWLMlAuj5WpLp8PcLMZnPJK7yCjdnj5ybfYMg
CmudN2TdSvdLg8C7AFkk1nnRWZEuSGnQjUO8kAnfMHc8d7ohwyUpiIrOC/VMLUQ016boleCxW2+L
Z/g7NBwtqpD5Qtwf3dbrEpb4MPTKrFi64teNiVTjq1EAeE41BDgqOXnzpmIsl+c23h3ttagFl+Ke
vgP3dYdc4xzEJvsgNoark3jB4YWO9DjxNSaxwywA9m9yj4lDqnSP9JUrrppqpMzfdG0HU4Zozw7M
3BR7JzJ/X1GJmWL11kKHT2viC+lNpzPgMasFlSrSdZ1wCg493oOW6jD3LpFDjWwPZnPnLKEbH91z
t6ehROSVQNIA1nuF1E8ufO5dGLGexpa9FOoqemGW9wfYFMEB7pEz5gcdMWb661QDoq1cNoAoTrS2
yvJp16giufROEv9+iyw9Xv1dRffdiufPm0x1PN09GYBlCxmszMq1MthZPe95LCxPzOMY1quwHBk6
KT0aDtJ+0NBY9O+DPaMf9YgatKsPohgBhRyCexIuIa6wkQX9/j/96vogCVQ0WW6VgEeUsKdVYg+0
rh1tJvauc6TYpNMUUynIHrbhx9HNb1+lGI8umN3PQ9im6MV2ktG/tDAeyvQGMT2s9aQmNP62IQZn
RfsrHlCw60L9KlgxT1ip2O3JIOIephwyKMKlKX2WRThCnjF7fxHmH1IFRWLRMqR8AGRsOs5FdZMi
SIlrkgqjsRlwQfYK6gPxvAh/u+S5NSW5Rtj/PcRAaYBfGeKwUEf7ZElITYNxNBgZ4zaVRzl2io88
kzDViO4ZqqPKPdB7bB/vLOSyiIR4xdKzaVjks0L+J/AIiUzjl/Q3VckzqANrTVB4QUQSqAFZIaGO
zRleXHUDea/1bfFbaQY8xIqabc7Q/pVBqUq4Lj4j3jeGXrAPQvmSHL8I8ovz0d5K8gEmonl7sxP4
RAx8dmEHvNTHQznwdmpA7iJyuT9ytENWpI6Ix5aKCkWzHXYHwGsLTOLgvcgVTO4WWMlPyr9btZn3
ybZXnBeC1ROovvClrYhDL1NwmEPndxO5Ox7qpK6ddTnWilSSpN99CtKwmMjTkhWPim+OX8DkbdmE
K7cCJCj52oM1XNC38qz7B6ug/EOc+oszzcPqQwySxFgP5lZnDTyRaiQCRaIBftdWeIoGia7aH4FV
llJAXk7+/l1mxKGjOgVeYdbyzRU0Kt2QQi3YD7bisEvEQhffl5yDgCjC8GFJRYIclQs0fuabWdXb
YTWJhTxAR5tPm7Ix8UWQgGWaKp8JmLXl+WpRujAmROG/FmrAbyJth8yx62c/i/hvgrTw6lj8Zjyj
pSN/R2NLJa8tGGX7Qr29YIl6cNOgcWxZyo/yEl97lpR4v22Ug7r76CmGGHV7fKIBsN28cnPHPzLQ
7yQbSIc7GPOXZc+729yQNpvnwax0U9Li06yu13+5alaoOW28nlzefBPS4o+xI6cn/Tt/fqFKdCs9
Z/0u8b0OvDQPccMq1CO5YYyKQyiRilOZkMhjFDB3VW2/ywP5H20OpxPIAyLaI9NnCt0hKUBq+a33
YRLBqTBTije5g7FVkCd9TiZu1dZO0xQojNeL32la4PeI3f/UL/Ucn8I1h7RLw/Vb/TxiC3+XHHo1
GzKveVfyesUKz7lw9XtmzeBFkxQTAuiGq9tDDfP9JYi5+BzldTbbQjr4rZciI7UimedD8AGVVp7Y
OHiLi2aJlOXSm6ieluQeL7ANVcDRIcSNwwVmU/MyIyLyl3o0iFZkBlJTWW6vDM5nemBMtvzlmV3z
CgAk0SnZFj/XdCvwpQW+T2WDOkHq+xWpUfKjmxD4idx62x2gPaXebhx8J7PwJNJhMTfXamPW2lrg
b7kOy70/A44lAaf7Zk3Aj8Ja0c5at5H28ZOReNaVHWO0w+s3qmH6YcqKTJAeM44qHvj7JFk/3Thf
FSlMfxmu0vQUUEd4frJ8lrcbcguoxfJXrWP9wKIMJTPbLqwtKIzL5/JXcGF97qcC3YUEEfUcuAaG
VCOSO6k4dfHtHI3du7cxm+f2bjztjm3nyhVhQmp3BJmYLfV4ES+LjT+hoTETGwCbq6MuSGj05Fyz
99S+zCyOwMQDf2bygOPqrkuB0JlMIYO7baGuiUlB4kCDxrNLHBXco74aoknc3MX16CVgMDjBJ0Vz
vqHqNwLiTUOvWYOBRhOeYEE+b1kolMGTjTjGLxCCaKQxU68/b3bjuglPiDQENw9XDstvMrzzllgC
72zzxiUlq25Pz5hhMxYTwEn6e0W63XBbjvoPdjAx+mwV/475+Psb+SFyMmi61CaBf1AEgFFVTgBW
GJ6FhkdKTKqxqD6ILN/qMfn3X443VUybAPE2mytHijPLXGeWnfajz4ewx5Vuw19PfG5E5pHi+7Ic
NfnUeQ41Uxu5CGuZa7ft2kk+7RifuYFvLi3Q9iC4DwOlS4onA/qHnW5/JkyoenxMnP+k3M3IzZup
itVK2lC/of/XqrLfP5onuAqcFEiiwykujltcmN7ZrylFPLtdqFYOQQV3bVzWPjeBsohsZNi8FRW5
zXj9FXYo4A8wHbNrIewqXCwnuD3UCwE3TeEufvg6ugzNK3GZvZi/PMRH1/K/BsjZHXyqUjEgno++
9IC8f8fHK6PWQsKR2/lnkQJaiHo7O8TwaZvGGQWaEKokEKmXycGBDq0BL8Kgb3lrwWJZhXOPUXfH
RjHXZxrws6uDzqT+fm8gutGgokp3FkcQ3jwTCmeGVeRvqCxieBibeyAuaVYQ8epFS569nR50AQ3T
gcIAtAuHhVy4QAusw3IUeMRNCECOXiGyD1Nw+7fWj6v8OjDLj3aywbLY3nh27wvUXj5fMmZgt/BF
Rj5pVZ7rO3m/nQ5HPLXyKGzaXTnMe7Qh8FmNgSreRJ55jbUDAYbZwQvOiQiAPJfPcWWoZM1FhZhA
wjy6h7I57N/g9abv83aJ2XFgbxg/kYnGZLLA45ByoTmco0psdJgTg0bsSZTLulTbLVj7UqnXSlmQ
OwylGz2gKyEDJtA6GgOcTAJf5VStEERsU1+dxwKGZCL6V5CMV9yhjQMO1mkrtZsvdcn0eZD7QYrl
u1/NEZ6Ub/VEWpfkN96PNgb74+GK5odKHYy2ZHwboTN1gUROv/K3kvbF3JwUaLDN4XCeHX+t1T/r
ZTWn2mKfzvQgDHRPD51Ff4FmNsRwaw/bgoDrmC118XUMrV2qi0RDfnmec//2v+oZYByz+lUfZ5Gh
6SFJjuPqgXEdeahUsGPSMRZecm6T1W/b+8xTXJEyotmcfS82escJtGxc/J1BPDXmdy+NuB9tm3pl
usRxYQVaxWbwZh4fBpXOBxhwija21WF5RqNVTQnTyRqd7RBSN7pdovdViu+eGsCqlDkT6aGK8LhL
mFjkSjvR8DNXojEWq9Z0ofpU6fLf+/Co+qh8TxIHjkprh5s7rGa8iG86Iym/bAjQH/bw0l/2vv1o
nFdZyVfYrQe9GtN34McHcEj6dWf3d4uUR6XXYjtKp79Z/qus8IUP9cxNoind0LQBHSjm49rtv0k1
Zygtqm6VfuMCKpgV1VCBxuge0463ir4bZPqO4kK2IJ6SqNVqUNmokrs0jIUC6HmaEai4mS7bZBu/
qKIC5cotpO0v4+AyXox2BUNLRT6zPYVmTiant4obPGGKwivzqaHMrnh5AVNnSjCw/lTKIpG2XyiP
Zo4IkSA7bfoa+Vs+Pp8WDd04miod8/G0Can9utQKS19OGA0Lj+D2Gsq/VTkS2CzvQGCEOBl0Aik2
eVhxSl6uVWqr+/copuzS3mBqzBT/4ab9eQqxk8DIN4u4Y84ov9GAHsu2cTY4m29K2k64CtgkiRbk
TKxDxjehEMGvEvajXHxnzX0y5h7I8EQCCwusgZVmZsNCif2RMiyhseHcCXNKQSs1ioAWeDbCo7d2
54QjE5TDEp35mUkyaieM7/cQnEU4EYGMVbE4m4aHQPwOrSirTIRPky4e13iTvpmzyElcoypSu+ud
3yel9s1V6hysP+SmDklehHiTwlrSU2YbcrAprDjE99TrSZy1Q2pEeHVuFOj3dPeA7pfKzjAKfJhv
MbuhWWSMJgtrlZ2+RITEORBLyHDYJT0u/PjPPWJ/+0Korza3AWDfVhTgSQVYkrL7QxcXgo88H11a
ZcN0YPgy1SBqkysvca5RWsNDfInglwYZGLPbnvIQ2lKzBJwqGWr6fJPamuzzVXIQtkVBDTPG2V2V
VbaePsoqkDb5X1DJWHvUj1KPP9ohGP7e9j5KKKR7fZG9EZB4B5s13EeAr+QshUEhCBhVVAsvaWyv
CS5JpoT+cRNjzM/LpFZSQe2FFOMhDv2tKQEF/M74xlDg4wAQquRfEQxvPJ2jiilcMEUJZtjT40aF
VWbNe/0/4SCl+doFi39K3EOIsFmaQqRm6cPtz15P6g6DzScKP6g+qkCsRnsCH77rPoWGXngrCpKQ
URnECdLgeYlVUuYCNoRKRoiQBqlQB/uCmhR6mckfCrX+EgCVleEgnM0kY2eWihOcltwl5YTep1qg
vazMfqNflpOG4eF5dSIgiST+9eLr1Dt1gqCjmp6YosyQugB20OhZw9Z0SJ0aHrrZ3m8cQW873UOM
NBcf3Zza4dewCtVu80Th7ts72sQ04b9RQu3JIMr0p8WPy/UIB3gAS+aS3I3zaZPtSxsXQErpOs4Y
0h/H7fuAHKprMNg5JWMArCR0DXd7OguFMQ+hRfrX0m2ZFYyJ+4/0Zwak5QtGCjiJFSuSC+iJ0dW5
9s2wrJn1uD/1G9es2NCwQciHoUb6oLi4zHYw/p/4MLjokggqgF8gBdu6iKBDhG/2OdUVHRqK8XIA
XlowmYtyPhXItu9/NzOSfkQ7Dhh2a4DJv2jWMdj+cN3XHafI7XDebiQhwPkHR5N+WXSMy6xasAeV
AnHkj9VX1f3Z9W9YDehOhR86qDJGeAxtzwBjpiqbZRo0Cvu/KTqlXA6GYjn1LHoEVUzD5OiKCuoM
a9c6gwtohoSCGK8KbuFpKi4gL3OgeaT9AKb94z+An9QfzHXV3aOTink4FZ+kXCiPz7VCY5a0gQZy
04ud5aa8SFTYbi/Nfk2C8MqRgDCDgh5eqB2wu+Fgph3N8/R6gIFIUuEGrFm8k18sOmWDeVce/VJg
Hruzc23TH3yGO+LdR32aIuvZzsfx1PFSDhjTfzWE3pBSqp91DL5sl/ydqowLmx2u9mAy16ETkd7b
DBsZo/FaYjT2gCgr3kRLR1aKhCF62jpEuFS3IGUA+nEHLbbIhzTtbm3bUSfAZzwWGtbpi2d+veoQ
7K+E5Fby9WLYkCCMur7DqjGyDfVInB2KEnJClNrYzlDUKDxgy8jwjlzIOZjxmWfdWOpWHYOa5k0E
DxAKxDPgfeSdHFJVDT5xoeopucYZopvWRoTD0j1E+1OKvHVkZTedQewu/4qkQ45AagoOy4kqzmuu
s2qYkM6IPcVddzTXbxR50NLuEUSvXjs8fuYuQ7DC7EbusJHRJPBueFj82g5UQFVwh6prgxlbpze2
YhG6Gu6euG57YMKQe094n8/aSIPQF422Mx6VxxHLFS2eDXj9/u+ENbsoM1A0r5s45+vTTLb+rZMh
lyMqQltyF1fKww/Ub6uNhQVZzoxUfRvli51ghLc3/4yC4jfnjF/2RlHNFLqGHGfcFvyqpxfUTfa8
9WC8K4jBDFUiJUwtzqe/VYTLkndjoOVd/PlCdzmMO30k67BZ6F0F86vzWCx5WVxu/3jD21z7d38m
OXy2bN1h6P9RGcijQoh5O1218b5avGp9JFdP6U1RwrYGYTQ9poJuozNbcCJ8G5GEMZiK5To1nfD5
AaQ9bfBz4E4l84ea6XPZ2u/OzSVI0P3b/Y+EnY+MsbJ1b1xpoFu9F2eJxWMKb76GqmZtGb4IA/NH
JXZR9tJotSy4V6HjS+v72rpAW+IYlB6WZGrjFPN730JV2ao5GjfNAmr8OC9W+NJceAzdZJ6KTAzd
GLvC38RfLONfclFP3gWTa2gnGOStYMrYm6tgwMgnmNe4LLezC4ng4EdpOeESCmViActnnj5u1+uW
WeY4lqWgsz9Bn1IJkjVN2CghityhHb9Hj88mREqMHNvj/P9bPmgetK9skh5GGq6qD9JRr48zFfVi
LiwHzUDZMFEMV4zViJr28I+0mfzqfpYjb/raZ+doPaTC3ouP0z8aTfki4u5l5yKqT1/mh6/CxAko
WqthO/R3alNYTNFPVBLVpG810crTgWfdWihs4WrKIgj5WQngHxkTXjLf+pZM7uSqO9lnyRgTSHTW
6eXE6YYVxKVnZOAgtqClHJlcfS6XiiA1Rf9J6+KNXiKuXuD72NUxHmw8rxx52sZ8ZL7r7u6nk/AC
l+2UwXQ7LhLC86pzA0inCVlYKczMaxKQdPt6BGZK8WytuMkbtTO0u2fUPxCowBVMlDGKakA1wZj/
ezAJv3Qf6O+tclBKSqGtKDYJEspo5Ep5yTaqpeKmfJW1bUVWZaJ/ZIRpfcB6aJKgTktwepzwSlmT
yRtqhzSArlOY1qdoBR1Kjvw34q+HvgKbGuhX6XcdXjndGGzSQvRDoZr2GdrEDC0GcLoZHzQfbpfk
xeb9+AOOzYOForRDEDn1/Dw/JDg28MC1fJ436gsoDoekuLqp36o0y4hRkVVvPcmR3D7oM/WSgRnO
7T7yLsKbthyURDeMrcsV9efGZUTUSdTnog5i/cj13mnJ1c1YuSdTTC6kR4gkT7skYUDaaQckSEz6
TJ6T1AcQwY3d0dy3qChypvfRkoM1Zh2YS8HKldwsUIfUoHhTjdO6CPaiMGnVp4EiJ00iXx64AyCT
zEXQ0X9VrfhywEZcKUUJtaImTVCxhX9w2MHaqWC3Oy9Glkyn1qzX7kVoXtfoQy+I9yZV9WXQ/aTW
y90Vk2citPXsRu3KB8546ScPwkjdly/koiBbznPyNWuueyfGWbGRu3RbZ7Md0uzHUJLSSdcNie+l
qFmaDfIofBzYbDatF9OpCFz3H2FlUfzrHONzPfkrbeIFgRbtl914o8efE2jukbIOAkErEz9s1SwR
OzBTUCZinNv0P/Oz4JXbkfEslIC2L5yc3X4V2lqbJWAHgwLUYp7V2A7r+wK9SsO6Q0EIopIaUHZ/
asasheWrzWxhQ5fsvFsDZ+mLY6V1WLJn5UWT9nfRIoqFEq+x1TexYCIFhuiTLfBRDYTkjVbFnTy3
K2zZz66VPapeDNuv4T2PRLYf4vpgtFVL6bIaEslnKZSJhd2nhoTtRmfJv46tZtvrFUR8b47To7Q3
tuX3qA5JCNC754ar5qB+/Twtdxohr4xZCcGCVVejvDOPY8PCCfKhjtS/i2E1u4QD54qmRsv4v3Y/
VtXEIlgHt68Iv7ZjuaGvIPiK5F1qHbIFkOGN6IDSk1gzJYyoi5AhY3lak3rh3JE2aExvCQy/u1cW
IuW1x8HA/SVDpgzXngw2Ugl7/4qej4eg97rA4gRhhl0CBLwRLC4S1udmuNBdnNcT0HqT2bSNfJ/j
oAKE/sc45xXyubktqTcMpytWkYNw5j1GCkjgR6hV6sKOZYWzGLACjNTiadwOKi7dExiygn/GMcTt
9Tmon01wIEmxWAhdQiu8y8luqXhFayaZlxKVDOSEg8hYh33r4HiaX/yeWUiz18h8rQNcWfX10FQV
6OHpNXTF6hxMvyx/lRlTlHF30sITGh/ssKa2NLXdjqeqUOnp1xNCUNO/C5vXeviGmDt7g7f50jqP
1/qKrrSsZmOoi5ECV5haUfCw4d50Th9AxFBB03dzOH44KFjI2DyFyM6NacDx+r8tDb5EnnHKc+mm
PHVgwkjajt1cTO+xUag8vnCRz991rIpSuNKGhmsXb+72aDbbyEc7J9a9PZqyHdj+8Wpi25SwTQts
/3lMp6a1kwBO5zWlKobvTlqXpcZvjCHfazeqmHLB024s/DFnNeXkNWIHFDEe1myw73CXLrxthGxC
RbjnK9uTc43WSGkKbM8gkYBbKLjWDpfpFvRAzXq0zyvPOIBOLyaOiP2JzbYhzqqMbKX9NvB/Op/k
EBSN88OYBixdFInPSleu1SfsTcWl4QI5QhmiksAfVRsnb5ZcN15nTLXP4c2X6WkXsullfsqYFTQl
n5S/EGWFsqrVJI1tNyS+12dJxb69uOCdpuSt29Ld7Sv0qtFCK3aC/V6mlzGQcf1HdU05bs9TBiW1
P/23TuC48RkUKfGYt+N2utBU55Be4YwQ0512IjHhe/OYXRW5W6zyEA9kcTOEKwT6Ye2FEWV+eojL
6wx3ZSdx4LnqV6/xdBBFbdxAhsQ06Ii1kL2lb+xzcxXL3ijqDk0Uj0dpg5JBGcycPIBtDkSEHNHV
1NpfDbjOxOZAAEln6flZxXU4nafk+uBeN7wbyQBYniWdZYUSLNtnCIQebVrn/EfztD2UE78AfyD1
1hE7UnmPY4KkQLxl1CvRPZlG43l+d5x04wmAtr4osTZObK7gUFEvWaYE2HxazV9MnKQ+zpN1a8qj
gn3Q0jtCswn4Ad/Ri1hPUWzUZ2cLu2paNNYo7QMLRlVzm6zoVW7svrD2tkmrA1eO30k/OZY8EzjG
2rjvlYa1YBLoGayD2qu9+GSC6FoVGm2bl8TLzaHo/DtHpjXzVdIPm7mbxPDle/5zRvFYlb+snJkO
pElx5PHQY+yTFhFmyQNRbkETNZHkxz1RLdnMA04d0sTpubN6b9GVmM3ytpAapyt+lFQI0V+w0hJW
P5tHPysiJ1R3xKv5uiKNbqRzA3yKyPbI3vJWxsMMep309EsDK2P3uU46TeBwbdfpINF7p/gb0as2
q44PEpR2chdE/k4/uuxo8tsAE+gjUdmGObY7ip7dESf6rwRPqNjszdz00zzBSa5zJEb9ghjnRf3Y
v9edCGptlyY3rJNE+rheulfY+HJ3UEmOQw9y1hqj2oB508tt8jm384o7XhIzpVOVTyTIubh3rHuB
fGWLZ94UBXRMbauvgG9OFhCaykODq//xS1yrVq/gGkSOrbLWNnWtbWhBu32mELIh7WDJxG5ydSIT
Klx7XJ3vfZ2+VZcWDI22RVR/Fk3vc3A3tFOkWoaiS/luZKW6IctsVA/GdDnBAeMz/wqYzj7PjhnS
HxnP/SL6buPyHPaTfBY0StttHym5LubddbQhLVQ1ByMg90k6LK10LSBvgDaffi6BMfU+yfdvU172
KFiEY2f8FiC7ifVQ1mrYSaI8kT5kg8bc8mse31Z8e98EAt3UHwL7ng+Gw8Kyx+DstspUcQhwnZMt
+5c4aQ9VAUEh9F4gFHXBmZR8wx44lC/x4hVELso7KllZuv0e1uKHmz5ISBt1fxM0BhVzLAUg3WTw
hB49B+TZUy7GpBX8S0Quc1beVaE14/uVgoUF8HX1GtWGeH7q8XDowL30P/EvHVTPAjTedpH98L6G
6TW5SxEDiOeOOHrabrXRMrfXEv2dlMVPFbQfRyFpsiWlc/dC6+5XiAQ0ohPmRv+1/dgBQxqF8x+2
vuE21NQNL7FrCiOLRYJ/u0nzyYTjUlAdo5SEe0IJgLjBj3TlRZZIwG4v4fg1+bnfgSN8fDgaJORa
ibkA5q+V5Cc/NBeuaG2wubwotjRIkaugUk0ZLTK9bRUm1nxesYzTPj9E9dMw20WQlMVMfwEG5rDu
yDUYu9wbfuhDm3iucSLgnjBptJeDDZ/8efmkoNi7LlOg2YcTjAUzUUeJuqN65NMhhXWLa69BNBP4
vmEJF+dXhafhwZr2RK11bCSNjA+PFocHyuQoyks1awruvYPBtjPM0HyCCLkY2t4oIdHctLFENtOe
L13RBT5gLuCVvzqvcV//1neBl6dSiE/YrGB+icj81m17f/t3a6wYG0L1zQFdpFrYSdtMXcm8N9tC
I6pGKgUFdStx455KEbwd4bYd8BqwgEX1Osj6Fbbc9TqtFcPNsZb5c/FrO1t+rNueNcOeW+FFf3hz
vgQuPd9pSI4dlADEQrHARN9xVqY3/Y7pYIrDfaxs8GfcxPNs5N2aLi1ueyo6L2+UdHDdU6HR7phF
RLybarPAcRmsVGnC7+A0yal6Jy8iPc8ESGOFwQ+gfdUAfhCIfI782bsmONd8TxNFIzcuDbvbAChm
UeSNMk+J6KThR//eaAU7bAcE/dmWlcC4W7BDPiq+KEmdb3niP1JP6GUZGhEFFO1IKWHyFJP+n7SF
Bln2Vz3gxns2w9GuCy3+JNF87kH8haRvGE4u8QN44oApWCftTYS9g+5vdzG8+0HrujwofJHEfPCB
lHfnOXxctPtRHtH/Sm1/URQ2AS9Xtxdy//rnANfywMJCQdOCnPSmdchtpcI7SgQWIrlk4cXFwHr2
t90/j3oymuoLfOpBGy9xKuzu6LV96/02O7YjFX2CHrP1v2zJzqlT/lX+BBv3TDk0lDapArdmDJfA
2ty63gh/dlJDhgKVOe+tY08uok48Iur4WWgDtP215iEEkWh7NZg0Q+CMc4FUhN5lMnRiwOWt+NSs
104HCvCplOMO/P6chceRQiiDvNmOu9nnkv42hb1TqcRmyUYB3NiRmHllesHGjBmlbTbJK5jpOfcY
jZgw7cJ2afXPC/h8lpcxv2NNKKmMAo2YihnpgF2PQ4OnoXisTrAxk97v0HTkfuUpztpvbKZgtySW
rcQw9pRYkBbtKya/sNYrMfPBYE37i1y0ZwQ2WgvABPPdCS8oVjKwEKvy70a0Ja6Fosf6RxGKpjf6
9gmjS671+Ju9dELw5Z5KVnch8LSAY/IsYf9aPV+thcTP0lBW2RXAw2MQGjPIFp8rQHT23wR+fHK7
ltmhXJ79IdpcGpb1yqd3q/nNxHIPUuqio19fy47A6uRqHzQdF4GHXykSuzZ+2y6oc1VF929vVtDI
EWTxKwsNOQOZPN9R9r0CMyBN1/ZHK+m3vAY4wgnbRIYOZ6jyEDY4PgnwA/K8Dh1mT6dhT+KoHrLb
hc1YAoUrpinUN53MVvd+aRqgvBxzzBhaVbNGylkJ0qjac4fDl/aolPsLy483rnQmTPl18UlfYOe3
wxsASIuvmM/oPP97RvNN170ndvWVvbXAXt2XzcIj9tRoVxClZD2IwUzURFiVPIXo5IpSwRR131gv
I2WPdH2hAqYRq88jOXnZRhmcVHYHIPjrZogrEmBRB6ZHuZ3p1NprSAwzw/XWu5jbOsGat8vinTgF
ezzW/3SLdRf33dHuUYbDPbtgZoO5LzrYZHiFO7xy5RCQ8WHlyV2DXlSOp9nXLb6DI7E1tMogz4ZH
1/aC4TN17yP9GyU4OJasCyIlJyaJnF+ienG3M0p5dGZSN5JT0uLpx5g8gq+atuLTDOr95QIEYBCl
742UOvxm8Ml/Xf6Yzl6uamAjuSpavR9O3w6uOJ/OmjCtfgeKCH9ZoQD5XsUSiQ2TZ8wlI6m5+8Ag
r5Bs3OWthkua0Us7IX2chbjhw3gVpDAss37+ZJiS2gUWVuniZgPnHhD47zB7DOVjt2e2E24N3jsn
P5N6ithdhl1NHX0OMVx97A8ohGd4edSfo3vCTPDPXBkGxH8p7OJtyRN03jOK3erGvmJWzYJru3Gt
hmL4Q0xgbGdW+9+4C0lWQhi9i13l+Z/sJTXYbsEBnd/FFDzplSpJl6oG5Ch9GW1sgGlLRjL83tEz
iTlEPPYVS4BYswQeBZPq74S1xmy/8jCADztzQgiHIZ7pU/YpmUVg1WtuDJ08TGMlFs0VckTjzijY
dpq8T8nmeBTfJBfEGmc8n2QzJ+kKfGAm9l28EVL45kUqWXY7M85BtOsrtLttAFm5r2hDHzvOPz7y
R6kp9OaeHUSFBSPIf3dqoFv/Isa0xdDmxo6H6zg1i/tf3gksj3vRIK9rrklW8bxIsCUyLNAc8moS
RKf2/7FQ2jwRh1sA2fn7Pp6/Te7De9uZASdN8u5wJXzEBgGpLQ6rKBWNYH7knfusgdN6KSQZJL17
3+AVfTWBw+LY+UoGnWqE/EMxy4thudaiKaJh7gRGwN0VtlqX3Ve269EDKjgf8mrpQQQjFself42+
XZDjDzhR7Yw+oyBwvAIwc5uJ4DTpil0lb9r8h3NlMMXStUViZ3hPlk0pgxp6V5Qm8o0swfEELfCQ
DICI+Rp9IdLqjsNXYiQpHKyIr50yChNMFL6CQOkaaoQfJQQYNiCCZsxJu/5yYKxzQPCF1CvpPwB3
xHi7aHGbGWkwSrv5qiyLe1/7euTVPbKkv9ORJ8iwVdsuZSjGENvZ/2FqqUv4hFVhPKyESGGN+qvO
LPBw8QoNsK5KcNhU+/LO6cv0KlF6iWJheqLTqcAb0ldK2O2CSo019ZmzYR69IsKUKQjTsh6EKhgz
DWuMKaTE2B+OmlbwJOCX1l5U9Q3e50knSY1S6vldSMBAPGR8MHcJyaypfUEWkfmLUHbHIspStbzV
0CkyUU84/cRCcE7laXPp8GTkSO5beHxuUba0GiNYhlYJxErMBo0RWPKXGS/eVEOW9IT8/JntZm+C
lFhzFeKikFHV9rlIB8lbEABgknJAsjdf3d6e1k44sLK2FFBGjpt4y4Cfzx+0EPeocSBkILP4Mmi0
N/hIx2pNIojkkR9rvJHs6x1JBcl98MyrDUWnUvQG6rP9m9t+t9shXbJap/+hgRrfxZc4JZgHdfjl
KFYNfu1eoq4Xe/GBb+C6i346W15QY17IINpXq0VsusERRvmNJ1ygZeBjHDaIuG3WBKi4KJ4njjhz
WIGny+Gk2W+Ma7hkbKLXOx84ZVF5WUW+BlM4E35Jyz/wpxZDczRC3K8MgLMERt4qLtAgCGMVUwR8
vVU79hbRktl9adUAg37WBqO1NvUIE3wHHztCyDoQG3pxcb0DTs1jbHwO4dp71gysSh3UIqGexqSm
UTbbDkTWWm6aVekjafGRHfRXJrq8xb3+BhkbnCStegzpNiWSdP1VUSxzdzWYlNk5BwQbHqBKjczj
6GSoLKjzEj+GYSkjztqyUMfqfevn+/BobmJ7YER1KKK/ix7isUwnl3XP7NbSs7L3lAFs6ktzwogK
pzaQ8HTdlYxfiKeolyo6fQmFNoaTPl/aIphGazA2psfwOM11K7uQ8jIGPm507Mg8K2wLfFlyTSaB
tQ5qDSkbcxTv/nFiW0gFccvAyxsNA0D2rikWVSS6ZmyCATdR4MOl5LZFJ28HC+EvkULoRckxs8kn
Q5ZtIZXZIV2WdHjWFGwmRFN2RgNUN0rihvOkaMLUB2leHg3lh3/KLqyrS9gFaK27pI+sJLeSGMLT
jlPDj3h0LufADfbTg6eBTjAIfBT9IEc3Dr3d11rIEAWIorDXxB2V8soSuV8JodBpFW6+0yaPlDr0
RIRVtoyqDrsc44m8VpGV3xgxUjC9EXLpGr/Ep3KxAj+O1dEBgcyIJlSAPtH+2msRoIZ3sFcNccvM
qoaoGbzq93y47OBIeGJH1kI0XH6j6th8qz4Wsm7d1hcGGBFMCUGkBC1HhiUw6XPz57Jp/SUT2LJ6
EjtEtPqAWdGu878XHW3vT73dEPZYtZ8/tvlwx1LqE5UMcD+U/C+Ur+pDOwk2V+Ec7FAlUYqOFbGK
4sOWPQYSaPvJS+7QIPXoIQ31lo8up0/+QO8+IT6PhdnKZZgNjpfe5CrnmEcUGp79KFPaKYzVmtqX
K5K/muuqv2nq/s1YxIVsXlch7Zel2NAK4NI4P2Uy4ifFMVRao4JNKOu71rEvcQyBzLUOkO78TSZt
fnqPg5ShYBSNguAOoE2gVqUQJGV4ubd6ULv2mGPLiAuTuELnctIpKK2HG6agA0U43xY3JOsoffat
hU+VCCTzjrp8WXGXvcoZQ38xSAeKDBKGhAZxcd5BRJf8iRM3dupfTKJqW3t5vnOG4ilE2CtISYFk
W7BrG3xEs+LB8D/JvnS+vBU/ZI9btS1Pr3up+ZzUP66rWMyADLOgNOyafSw5h9p7m2uor8iRUUOE
uqNYh7Wb7std73G5ocafqYVSzPHekOPXtY2Swkt6gTC/abtdlCTZSIIsKJBGdEKSJqoZMAcS9ttf
/3nhBRXu659ncLj705YDrLUzD8ZiaZGWlN9rnTyXmDQmg/3s3YXcE4Eh6ATxVE3OUlNx37sgcwd+
oTg3V8MBBTJf2Y/KbrYYNqWo8O7bmO9msBjLSwhM9RP9gWUnnW0S4efBeNeD4wVL+qXzZUl9YNzp
JNhCFIUCcmj+GX/QS7Rd6ZHF0P2EjIoouLDgXnUDpjzaNc+7PieiYksDwHUNqRcU5CvZbGrx84Cg
je/MHpcJPt/iLWhouLiZQ6TAv2ETkycxLwsM4IiXuZuKOjmYLNzjYln1puH6mW1oSNb68zW8TPzp
9lXDQr+R64Ll+xY7PE+lJYJLYWmYRjRlcXi5qCrNyB0om3OxJaFCPIjZhKf46H+nK4IbJDZicWT2
t3vNYvOvip/s1xQZqcWKG4f1YpllP65CElnbnmbBb1tAZTSBZygq0rM2Spg+BUs55lhLcBI9EquD
3DVIGm/hP6vIuiq5hHs/g1wlETK6CiiZ5qED7rhlMzWbz5+Dul6qHWtV2cOqgyuWc4LpkIx3MH+R
bi1++zzJHvzusvWp8uzJqpE7H1MOMnP3LRsJ6eK9jr6hy0U1cCcQzRmPSMqqNR52hLi4E1eb2F1Z
x3/Wn7eDKQcL3EYU5RINHq8PKsMLNvk8eAKUtkg70M+d0dAU5EUdwG7r+unKULTczmdOdMkaiznr
wrShX3rrIi8b+eDpLCU8NzBGj6f/pyWsqZJjSXzXPP4uVuzffdBNRphdR0TgUA8zSlRjQ1j91yyw
TI0/IuTTbIqdnLNHiTdbZ29IE5KRi4rz9GqSx4OmgQCUC3/vXpVrGkVAfscQzz7iViZIbo4xYo6D
XcmofcGZ0TceAvgjPVe1NwMhGyC6Px/5kbFG3Lcj7TCEd7cQ7iztB5oeCER8dk2h8f/Ru5dVN+kP
RrcmxzAQgU5Iddt0VJn6bkLPVdlKdiNU62/cWpc3bkG0bxogH7av6iwIDA+4sfj6xXuHTinIPu0+
nVmjpE/8LejqYxp7YLyiPYYD5j5CpIwOtk2lANEUAM6ij3zKvvrI7mp6jmdXhqyCBFEsGOtgF0r1
QVGZhV5wZC05iM87170znIn9OSwkZUtS3zIPc6jncGIHyZZoJ9IuxXz5kkr7bW3I9oPfrbJaxTS+
1gSbUxXx0r7FS8K8bIw6wnCeHH2BsBgGcVud+u50oB77Sd6yjxb8/qzVEiCasj1FBBP1s6hPzhkv
xFYU98dUbtVFSBogMtAAd8Tc0GBE0PCJVDrzW2JKbkuL5/3Aj7+C+rAfzMF92EHkL3J49A/FtVCW
u2sF0mrsZrXBMfY7gRmjuFrGrV3xQX99CqAgvVCUHVPnT7cIIolXgfYhh1dzEKoypfHORz85rvkR
MuzIAtawjEA3Rx0d5pgCpzDlH7Ny8KSr/9kWuaaFWsq460BMN0tmZ4Unqb0+dJHhqtB7Ap2LlFOs
RJuK/CMlnB9+oIdylpDvgoBw+lwnfl1qLC/ZfrcH0pfsjmBLjjRKwowRuPhCzHsr/FYko2dr+r/y
KeQ3R2YvtlIk2d8ZIglG2KaQCn0xEtcKbA4PyVJY5R2JbP0gBefxO1Bppjj7h6w1WVRvCbTb/Klv
JX+tqaGYVD2YSYIeZ92QczWmtA9OiOGK/lObQgkrSO9c6B1VgY2wOxHU0co1tL9xerIOjUHAUaq2
/BoPNEaLRJx9z9uy1ZPyKdI9c0OGbvy+IACjMViSBm7e4j9y/Olbn4oJgV9npwUv4JObJTHyIBI8
WIDfY0k4wn04SmDachsZTaB0C+MLNrwbefiwXQ7BK32cwpRMRuB9jNTFxX/DrLVWzQIchZg9vG7T
KcsK/Ezt2lOaSIYpaHfBzp4GVMVjM/JUC3FfFjlUAJkIdKlgBz4zIr4gHB1pyRQ6pj6MvmumKX9v
NAO+olpP4TjjHu7S/2vta8K4AS1ApSnGblSc/PdWRe25fMAptvGaZtrxMmky2gg0tpneEsTiuaFw
x0ANJE+s/Bq3BIX+b+L+dhwNxSge2XZU++OUwc38U7AG24VLwX4PkKnqEa0V+vidfb2D1UTSHG49
7T7lsiAPwawqOpP4Q6LpdtKq2+9zAE7/+OqlDt66urhfsHfN/z3hc4aH1HWvhSA+yMRnEg0qQM7I
x1dQsaQgXoFETD5rwbBaeENXrLPEFMPSNPjgVYwJnIK8Cr8hZW8ec/l29utCEed5RO9/QIJybA/j
nMJuw0rbgZ+grF3VZxTsSZ4vFgVxaZdLM2AehUgxr0T5TPTFh4BI7ov+qbiZzdA1GC0MZYr4HG23
ewWz2Uaj198XjvZA48Jw4OWSPOuSHvjSPNIDXlV3GNLM6mPnZBq7MoiD2L1VKD35X0D79X7hox9W
MlRv1dsJMKJawrUEU6tDxrxxN7Jv3WU7u+Kf0Zc9vwHw63HNM1K3eu2yh9Z9eW7pq+oBK3WXOzb3
+gjhszupqmLpyL2AXzGENxzxn+JAvgSpsJa50XYceR9eSbhOYmd3/JuZSp8giHbScLaMPUVUommw
6BfNVQ99WvxH3D4jDrUHHw/cdzWw5R+xeyxeFWDCWPNV7F74GNKqhijhYVr+uYvvP7LiwLL0m27i
ZRlp0ueMxKbnUo7ycjgLn2GNB9+4qhuqZDFCi8je61Sxb7oG4/27+CGVWdgZ5vw6Go8+Sr0ZXiHv
NivGAEoHs7chazi8kBITDC1yXMTJmwg6bunB735YyefBevBaNVdvwoi7by2faNFg0To7/Xku9RXK
KGCNMD/e5a1jchpB1aMKsUIzeSXrWN2CkfVzi9hSFzw9GB2A5qI2OeB31TxYMOV2sFg8ISPPfbzp
GBt0QhqH6xCEsDapg7lSh2oLdflddImkhlHHIjtfRkAan6Vp/5s/ic1aJzbE1KHqst3V06Hg4K05
wTeinnn1N8cWrkOVM5ID4ikvU5tz1fEM8EywFx3fZTGCLr51RshF6bWoAHTdDb1ISnaKUjokua19
2+MXojTomj8EeV0YqXjuaWoKmvYb6RLfXwjxvrpeo8RtQ51dnxBvMgX/YhcOQzqiVRkRToqZInhA
Njyo5eCwxjwQMxN3ct7y5KOAcippa3qkqqQITqkE+YI60zifS0h4GMxJYGyNihDME6y2k7s7e0ft
0RG3JMxb45kDn9PoDVopRU7/nRjKyyZhoLt+nXCtPSCRD69a+6oO0AEnvZhYMEgSSrXD8ldjMQrj
HNrztQ2ojUM1wGRXo179WzpV0Iur/YrZd2yKVlYOLbiZX30N7UHh2sg8qr0XyZgvIu+ACKaspmUi
lc+ShnO5h+uuUCEHzHajTE5u35wvRLFlkFgM6JDXPuvpZYp+t5q7plKw7t7oRmubiklY54mTAbIW
8//DZt4LyGloGcCMOvw+kFYrkrM0F6zG3+G488QF4cvclO2JQq4ZwjteR7yVVldFSqKjrQBbzgaO
C260mXMxkFy3BGlhI7qTR1dcZo86n54JJez8BLxOYUtMHBjGrbPyUEfgK9QdI4eTO2hNtuEo7zCN
RbG3Trjj05GVpNMqx7JWbFu6PSmBRkEA6IXJygitd2IDYOHB3l2HQ6PnRNmXHGw/fWPCEc/RhrVV
rORR/Aa6c4Tv9IJ12+EH+x+TWWYfeI9LMede+1WdlMjYXh/6PEKTL+kDM/XCCYSa6bOBHBfiPdpW
/N7Pw6D44F3yABtXYAF/rlouSkjai7CLnCw1Q0r7U4A+BHpUk2ChiIpRphoaAwCLI5IOfWtZC/LR
1vcIG2+QFCeX3ofJYYvjNAooRaND7Vfdplkj96tV+Y3Zv4C+mbdCXt5CJZjbdN9lUC7S6hPOTJxR
kD+R5pkQiGPspyRJT4kA6c1K8fosRtXdzTARIr49SFFLW8MzdtXOvb6M8fC4lChA55bGVMaB8yJ8
b7EpZYJCj+xG/aTFr7ARB9sLbpq4HEUzU4RoI94Voim0YJG1GOSEbrDB5pB78g2qhP8djoVA4l6U
vIctcoiFMT8t7MyW1pw5dzOZUKYf2Z23gqhV0Rmdeb5Zf7PwdmBFDE60tKKaILmTRGPG8DAuJSqE
PxM4zWo719anG/UG3xLawBylR2y6e74XKEno1axa5Xx/2aAQ/EVF/Q9yOhkuaNsbBaKYEsvcM9zV
29hqSZPoYrwL95Hh6fAzo/tLe2s9rMWscQdDDinDLFgVmz2eoTV3sICSMa54WiACv2ZCyi6EVwHL
bSrkddywgoqTwkEL94kDIKxHIym2/5ZJNc8QQGQwZXQSACol8q+30qXo4vUF4WwfhaAftphWEWxa
gGeZkmgFoUHpb1cXFrQMEX2gvu8ffIKCAuPcwjFWlx9wAqdsG+hOpTOeITLzxkcDlX3jMND5ysyp
t8ztJSpPXGHx5+u3c01ymSSS+q+KJYEejEd/9qCR0I9zvX7Pa1kSAJekpeem2Lt9Hv6g8txgBebG
kW2SYhVpJ8Y5azm0htSGlOG8lEWRRZPFDibcHAZOc+/CAp0bQbb6UQqdwW5DuVnSo0iuvL3hovFG
nApMZjVJA5oggjChvoZjQ5DPTlJ3bxVu1pAPMPecjBpbyhpXLdqSELxcPue2Fh0TMMB9Jtn3YSMw
wHtu4ceVr6J0vX+S3vJD3S1awq8yxB+bEd0jnQZ4awOK26P7bPaAUQNbFZNqln2H+HiWxMcKzqXG
mHaoAN9b6VfPJnI2R7iiOfGKOPEKs88ofg20RnQN8JZTutWboqWcWiWlRemM5UJwcEJebPQbQ/PU
NapW6VgcJBoLFiEzSCa7DCbOFhCr6gvamTXzEM0cBROb5agC4QVxE0R8JIZUl8DLKbllnb5/1T/j
hUHt6wScImPkeHTjVejYu+IRkZI4ErausYifjU8rCcBbHmNlGZw0JDxBs+slGuXm78NjHKJpytjV
54xItvmKV9Y5YduUWt/deHG3hpivP8F05BIMOm3xUDj2rYfZGtECal6GewTAkWnr5rvQYTr71OFW
PMYHK6FMo8fX33jcknoWMTJWj2i7biaT6Yhfxyf/RfoUrlsRmUQJOTWeSc4k354l3y59DbWhzve3
+aV2pc7IPXICd3BFDAF+PYde+YHDsnQ+uaFmsC+JuwE8dvQlVMYLVIdxLkTO5VBWaGmVqMdrA0Qi
PTqIbl1Yvek+AmRD/+YmIcrA9cQ60uLWM/zh8Ja6TYY00IpXaggQO3B2vKSZO9zpKzhZfAJJZU1d
dcutTGTuypWV+6kH4/rTUG8FWUT1Ky3okIb2LbGW1ffu0zLEl0VQf98JCwkwjOFIm/TH2jxX7RL0
B1mZ+OmXgNL0U2xxl1gKTeBPlRYuTEqlz8LatssebrEHuKhDf+P5DvUWoXLN+gh7YrBgINiuRVlL
Axgod8OAtcZfOxjOm0qTvoO0gJKqsfPAsJFMWZLKCxmYqaRTSIeIQJ7DnG+21SOP+q3K5hreuLhD
qjVX4G9I04zoCVtnwuVRW2HQgDFBhXza2ryyDIUa5SMi9BTrwdMbXvwBFV67qdbobvyeVtcVOQso
SkchgLJ4JT+zKYLTEvHsYjMs1jYIP3TwplX267NDx954LTBCSaEnKshczUrmB8Q1hJ3+l+aXEAya
7CPgWWNwdC20fQ6yz+LiAJrr6xmgxMX7GJ/eFAO6BZmBYCTKQ7NRKRV7YGF8+SGx7StJPiZeKlp1
YTAQRYuX2OqVnx+yZDKZra3V9jGoH7LPS673+xdqW8OASkGTnAHkQq61N3bOAVr4AIMUMtmNAsIZ
egPrhS9TwavVCB6WwBzkZMgI9kpEmZwc5L2rFN9K5sJF9G5VHXItsKI/r73cmOR+sR8lwJyDQJXg
bjzEIApMlkCNkGSdorl1KG/rA8IJ0BQy5zpkC4Rx2mcfHTJA8UrVV+5Qv2dX6dYc3bFljuCC3H0Q
z6ZHivD1zqT2O7mpQQKEHm75mK2klBQKS/fRFLTXAaUhuqP2eTIP56ex03AK+zgeo6J6gr1v4Bbl
2qYV2DL3u8vQG8yaDLJLwpq/54nx5RaWx5Bd7LOQ0yxqiL/9/GLRxQV0h1yRPepndPsxIKQWno7f
30dFM54UY6MXuzDs0zXqoD577qsSfBnDufvIyS1FbQjc0Pgb3WhrROt8C5TSDa6WOdW5+uFLTXv+
WKsgsmC57ZFIkfM8sO9GhvHpoPCkz5mtZkx2BhE2Hik3/QAbB8zHiJgmJW17F2gdPOK9yOcmX94a
pAdnt888rVyflrzNBJf3vE/wtNlW8v4lyG3RvZwxXUnQVhlxbt3FeRNrukmbwOEfsvoOwTMPYMk6
VeHoXEnCy721sYBjYCExEieVn/cG+4aV9TV7obuotk9PjfmhFeCqpEWkgax0mEmOXvaW/BWdXAC5
Gf+1gwi50wYVtG5/y/SSTSBlC+SU6yLvOAsm7Vo7yNHplhzZg4B38wEhWGvsiQMAVqmDEMPfTCbd
ZnbROU2QpM3gsc+3sWs4FiAU44FKJBWLJu8/SaI6a8ihrE+N9xGC5qcd359Dr/+SDPLiThJvRf6d
F37MxT0dOaafZBrtjhmGZqUQuJTp3onERMkOvl70b5vwv1XpZ7L+eWHV4yEeAZ1Iw7HDBAgBJTCI
o9s3E9vi0fO7Ei1xIzAzZOGfbLigx9JxB+Mvbdz1XjQE8uUrnYRQS5fwN7dTye7NdSi4mb2+8jV2
OuuVnCt84ksxST8Gqk/IGCKAJXh2LXpJL6SfnCceewmODojU2vDVe2ohSGPzuo4SFVfyDnlVsKVF
jNZ/Yqlmt8iYk064BuBKRXt+OZVUlcHXDcyx+r4vg+fKKUDenJVS1ib4ln2DQCUu13/G2oMwsbby
5v8MpMtR8iPpJ/rsQQKbcSu5HVDkPJhM1Yv0qlcx+D7ldqrTQlpvQsAJUdVxuTGa4QwdXiV+uUvW
FKq0Rxghi3fJ/nVeulTwtJmU6rvzbtQfYLcEUOVnLjmvzBzk743rxgvslLGjM+mxDZ0kblqllIzC
c2OMVBn8lM9x4syMEqTSHUoC9SKBKAfRlg2FuUgNO/GbHSnnSVIB3ybuc3VjUBPQojSHTUanpsET
v/Q58FnIhTYYhxOXcEWi+V/xjI0mCTx0LbKI2IHocdnuGP7lVaBF+zzhz5oKeFv64UXM2ZPMduOu
9QK3sbupB+CVaBZaNCBN3wxhOqdmWhd9F9IMX4rBWEp/opUDSrSMwsWuRbm86VIR1IYtHyoue441
z7HBoglV6/gQc9JNTfXH5mNCTQ9ekq6/gmX6O/4V1u5UzWdLKwvKFAi6uCreM1FPfGiemE/durp6
Mf/j7FMIq/F5G7aQC8sakLxSFwX0y8ZFi9/xIeFv4Ob77mW+9kp8e6akRiqDv1jvMX5bNnSJDEyu
/K15JiSvm29/j9Lw7WaR6KE4GGLmOPCes7BOkkYcWrDBcdxXwNgmaiJ7iGqxHqfzz/dRbnAF1cUL
YsC4MAxlRzpgcI7c5E5Cexn5cKQIbfrjpb016B3qnz2cEOUSyv5kxdrSqKQwL8bTYuS9LKJCt0xP
duLLnGANbzV3sSI9VOxZIhG1I/V04z3c2jbbme+/W+iPgejjwE/BIbgLCo1v7Ij+miZZwlcRROaW
smQdn4cKz37C3dKz+NKteFKlxrc/Ew0BQgouFB7DtV9Wjn50yiK6xRuavtll6jFxupdv+ru0mXQG
SNcNNHCQFpoFMfpxrU1A4gJbs/eM0ncCBPLXFh2F0IYu03YQNOHZpFbAqqsoqddN8JL4Y9cp19YK
j4+L6V8gthdYf7gUzOMTOvXvVECW8kIiu+hBpXp1uwFr/ZaNMJiVxAeg5q0kxbYgt0bzE79uX0/C
EFN53NdwEqflWszUJwUHRAfVj87K80Ioe9fnqqTi13fafiSJU3U+UEgSioF/Fjy89tPyb7U+oIQs
p9serFCkH1ofoAdKoI4vL+/LXSrCdiYzqAQpmsI8zRZIN3RSsFIO4dD9gkCp4YOZTgdfkcPNIxAx
65YQe2iXqxP4rXX4SQQQdbsrTIikvs8/kcRDgjA5PpEuSpRwo87FDIoGVWyP9J5HFNJYiC/MsnfG
YvumcOz7cg3fMGNB09gkwQWK14dFkcr6DtTdacHpOB90hPlD7OfdUOgbvhevreuHYf1M/w078xZ9
j8/3C+FhvuBttoW8yfvhzbNQOmg//0tt+6vLDknHJSKUnU5W4Sz8pTidaSyzN/bT17oC1HZMOF80
0HsbNPBLJ/ZEoomS4+qUAohEoQp0VYmjuyGnQRxkz4M5DeMMSmlur9sYcePkvEvGS7xL2qvr7uOd
mfEmCq3eqjTzqgTCKwA276bVPkPH+hO5i31m1163iI+8Dc4Nitxq1/noGs/0zEU+xR4v9jNCSu2O
Uzj9u2d7zjl3iy6dI39btZUr1luLsiuA9xbqpHli1h7v6XPBpbVqIgEH7JzzLIWZ4rEL26didD57
XJS2NiWxytfRtuq8eKlFjWXJknz1IwhBa71HjbPy+oPOznR8i2g+iTqoYXNN7VRHu2/JAW4z0304
GulXfzAvikEax/jLobNjOGe1kp/2HkFYjNazYysEsVps/G5ySamKRaU7kPxGRBc0L+BXEZKoMrg2
ZL6eyGzgHf3v0ZPbb/Bkn4JWkQNfyoHeTwFVHXHIlJqFMAzwZfCucgqn3hc4mMPeh8sDSyE7ov0Q
xORtnr0+pRUnGSkytWQSPce2hWymS37J0/ijEZ7SZVkORLLe9U0pvV0Cwc7NrFeIM+sYty8k6qgE
Dm+hx0loBOf07bAZLrbAGoB3xn8gtMAvP9ZBZKctOtDL9iPwKVYwxSHTlWqT9SDjjbaN+SQdV6NQ
68V4ntLT1nUzU1N3TUKW+QvN4iwL5teiukc0IbBaFfD7H+90ZvRTU2tgvcUlXhg+r5HG4kXOHtwu
SVSp8B+rHs6k132mr1aCJTija1y3zCufJEHOcMF03UihEK8vZut+5EIEW3/30y9i8lOY8EzBE6U+
RRpZSEqXwru2VPP9RCOp4kWPaBCR4QeM+aH09jWJU5IdcMEx2BSpyXkLcYzWy4EtqsId2ePa8M6S
2Grm70rrT8TXYp/uhpuIlvlAVHmh3C2Fdu9Ifqdg6f0Yt5h8Wv7WC9/19zLtDApDJAZLST39+quK
XKly0NBMYoOk3FI3Z30gAnqJAejX8Oke6a/3S/neuscGa6t7qOT1SLO2i5TJItU25HF2ABCttzxP
27twXGP7sA6zNpiQj67P1Zw0qROb4k50Ip3BNYEnfTPx1jjENv31UIZURBUZoCxgyHQDNkq1kCZZ
NkUmueCJMgMS7aMH9VoEPQQbnNagqC5PT0o91FqtuGwGqkDqZJpEo31ZqtDVUsTsl+Rn/QaG3by3
Vj61NFhc/xmYwyO9WUtNbMjPCkVTXLX0RMGSU/KAUkqbW4AlWug9u4EyADHN4aE11Gay+QPntCRZ
6GrGE0CRsjHndbiBuNUKtKNW/eMUAt6A8H9Y7c8HPotvGwDIBE14fA/L894DcWNhRkH9IDjOc31p
spSiQxcUwMeAm+u6B0y6pryfygCfdkvAf//VC4FS2bCMnI3NAiCWf+ykrcKAtrpft670/1zOW4Xq
Drn/Vi0rZ/G4VdEBzsZGG6RLnfWR+BHQV+h57rpJRM05PCJJSmgeem0TySR3rGWQ9ygGsqF4LvCs
OSZfXHHpCjig1VfQeQHs1KFax6PJrKO0Otsw885iE0UhfgxizgAUWHPyUQRDon5/Apcjii6liKJR
jWUNzvHWNkYqEwzDV4qmDosakPo0/vw282MUrjULS5XXxbYMKMA1w5FlF28gqutZwQhir2yVaTCC
TAduUipRAWs6zx+HbERARbHYmwXbt4TxGJnKtyN8xsMfW3eXR046BxQDz6nrl99N4k/72IrdxfyN
mvOG/k2gRBciZqKbgHdfDoom6hAdAGYko1hZ7VD/HvG67sQRL55RdOeMDf9l9+Wnj/Rn5NrlotQn
trgVpOcFoJhQywJsVyQggbmEWXAluUNAaGzbG2I1JCIvwI1uQGLBr6CNhvbN44ckoLi123k4r5GM
/dc4YcQQIYGDXJdGYfPDNZocl0sERrvMkMeaeRXkgCCmwwso5lwowOFQnCQhC46tkWV53u7U9zos
pg0WiyHb2SeVRG7cbQjP5sT5qyymDiTLyEezAn7Ge24F9N3IlBAAe721nWUBLKmVhAeDOGe2+SSA
bcqX8frGgQaogBR9CzXPIe5cc1NpC4kpSxfpCO9XTxGXoAAJIC6oJ/zRGUFbjF7SSTs29484B3Mo
JimFcA2dm49TFNeMwRJH8XuZ6w/KMXVNhQaHPy8k1LQZLEzOLU+hMCg1cnPLMXh3Pmm5FG3eWI+9
MrjwHpc/x8cAxl7OScik+GGTOBIUhIrb/WfWZDDsDiNIuuhW5bW/ZS3uHsfvNBjDBwjiwsPPKvrr
LjvqYU1gh/stAGWWPIBUO242VceVeHKAAGhuSQVQBUv7N1nq605OKOE5DijWjV0nUWSU32SryhC8
7ecLW7FOknChhda7H4VIzBAi4ZY6/7ebpe/tfUsu5Z/uShHtkqXBfEHoy1pjGdV272EuaV2p00Gi
kXdBafxit5pXQRfwq/W+WXm0saaJh28W+PUy9nw5RCLekgDFmP+Lnv8Ev8cCRIAzePK7QCQBjNDF
iuSyavMwzRMlCyDOLXYW3b8joSeHG1fYTjeUx7VUDZS/1SJ1JCKgJHMl1k+/B5OYbJd2O/IwMwUR
G39Oy/ZOCXtF279lARYKjFlKw0hGgJpZG72przfZliCSLHMbE/FTidc+Ma1fEkE6+U3CbtiS1N6t
W3fviEeJQiHV34HcdYV6cS+wLwFKJ/p5DCR5ZfQQepa/mXyRMdI4xZujojAJjLl32ySi4w9JKKjo
rYEuWIgyoptnvHOK0R1qB6vB4OkX5LzY6c/LxoIQbizghIAQFYOd55WuHsr/3RDVCfFL9UY6zu36
eQ6Pd0C6Za/yw3E0qoSzRfcOFVUAWtfZHa48t4g1m9d+Xmps3PKTivCQ5AKRqooxfFILDDQ19nSj
QpzdHsurZg+rQW/NHnl9csNc6Wu5S25cE81QxEgWOvJcobXWRW979kOpeVufnYFNtI5EyNNh/pL+
wYJL1RepLU7WPBcFUU0YgiIiPkWmvKto5XY5hdqs1c5aUKVdJMAmWHIGww8X5f9D9Odx2jAffG/B
k3dOMyz0BUU9W6n/HDnGxcISWJCjMPoUsqgbkNcP95zztQHSbv7v3MOagQkOMjQEQam2x3GIElho
oJxXYAyDKBxKreyLP62t4bZoAfmDxG5JKmeq0KElKQw0nwQmXnIS3t87W4OBomdt91TvnHIANzrj
NJ5uNJbH5D55+IzC8vSqjMnDjsZCS2Y0QZ6xB2JMyfdyIh8DX6pWCKQsNr+dn13VYcJDJFEEXeR9
WMeqPxDTvv9RIjgyks28Qsh5oPcOVrrMkL9gJ/AkN0kihsfBRGfZDoHQ6GvFHVsbj9WKxPlI1lV4
vQwI4Sqsl8xAaYwNJHQbf/+2Jjw/34wBoYMjCl1PO+mykRVllp9c4CMeWtMFour7D9TQrMmG0Ery
0tSOf4RcSfklCLUGNGVVNe+4luHDc0u1eHO7p+xQGvz4axLOSF6cGBxX8odRETQ1OUcvFmeyoBjW
sZ7DZoPT412zj0kj9AorHTLk0xyIRYeKfIEV0jxVIUeslgbl/dVDD02eN5A9Gces7tNrHrZhDgKt
wPK2HHm7epTxNnpRJ3+JVp27gySLn+w5EPZuLCgp4t/3Tqabdw3W7WzZoR5mSemBMIrfgQehB5cJ
7X+j4B2cgL8GkN2yOP5KR/v2lPd+7T9brtrkgU5YYyHrT9Bxrsi6kmOYAdwF3GYdGzgSJ1cN/g54
YtNQPJp3AlXqJ5ybfnzVTG0lLIuBr+1/QrQdPIYRTfFxyGCOMkX/6HDlw+s8c+QooRu2AJ4mO5L8
Uoy9ygbVuHqrfQU909cYpdO1CHVbpmwaN7uc7ISGrRggWwzUIAaUg+ibmJyoQ7/1VxGB0DDgFhGn
g5tKYWJKJQyqeKEcaDMXHhABvm9612fWjkRtE/Kp38lKW0kmQ3q/dHx8OMaJwqobLNtLTyNZdQIt
rSMRIlr2kDpSQLx+Po0aFgEi66Sno8HUqotZ3OosHQC+QjBXHtxp+eVmGKc4ouQYjrIEHMUZpsv+
oDdlIV04e66SsjBeBPdeTw==
`protect end_protected

