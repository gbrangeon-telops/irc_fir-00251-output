

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
GuWEw077quLd3kfu8DABFf0P+6oHLq5R3U5znEygNXmkCks1DFRW7Mt6/jd95Z4sdDaR5vCLL2M6
FB/Ff+rNvA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
jFvcfNCzhBWpeT533DDm5MsDXv4GiB5r4Bmmnk5Von/5jho0+BIo5IwIRMf+AlV4xqtSYYHC3I2k
BVrljYddp4kTGUJvHCrm4WaY6cktxQlEnZCt6LbtmRJq5bQ0+BhbjRb+yhnUtxVO+mqZJ8X5carS
6TiI+a3eiQyqjafsIxQ=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
3uk2ioXVXgv772p2rHBKB55nN0zepBz6/NR5erkVu2PDHMiL0sh4KhStRZxPeDNzjzcvfXxTocKd
hKd8wwyqbvI0xJMti7Zm3ArPWxG9sxsPGJWi/HV3nwjRdbl8Q5i42ko8FFW76K8gPbQTkcXqEX+f
TMDFgnzTvHtLMrE1Xm+zXTsDfz2iY7i6oQ9oV094lrdSLAt80D9E8ysTFrLsOAY7rvOt1c8o26ui
lfC5xFONM+l+w+GytYmCYLC1g3/Ymlqj+CUT7JBGrc9OLEVB2jBY9OOPdBfOl49VdH6n2k4l06g4
tPQ+CDbASlaP1IKOpWeipcMMiP2EcvQEvzBqvw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ODN1qSeI0EeO28pILhOMZHx9bb2qYpmwvyQXvKPrPhpTBylybxluT1/v8KSBCRH/tKp0Ke1TAM0D
rxIBcEp/+xGCTqhzkt5p1fRCsGDy/1Kk5L4fYaTlJRk43uSfOTxn6cMlcuTzjFQ5x+FkobtNDSvc
hzmRwInNRUY241xhR0o=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
dC/Y1fV+mqTG5rOr6IWyGTQ8KnFRPeLZShUWaAXrkw+Ng+xoimVrmPwEeCnURpwc/T0yNbEjCDB4
bGeW47AlClSVksRroIGKMbG4EdH+85GyM7JEd8UxBfmIEn2qUdv8H40fYW6ndPlPBbIsiprcQqu1
BO1TrP+zbizezYEZNLdme7klmciNF64y46dVM3KfXIDNKQvoLTlpJYClTv0K9dc9pDZOVD/5ly4k
Nh9OSLv/jIhCDn0y3M3rX1DyQgZeJYBkDd4IBP3NH/wojvEFQZAcMKJEqADK3qsWu81U6IIzKfXC
PUyRFWat+MUxb64pAuTyWw3derZjtBnOfD89TQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 54432)
`protect data_block
Q+nSGCEmBeAHy1P0xUaGXw9Yn6vA++jPuLHNwHIj4V9tTWGgGj7U8X74YAwnMxFWQ0lWRSvy1pnK
LgkQ6hS17wQ4up0hqtmuR+LlKYS0YnYxDuxuYShb8NkOfSCxkrq65cDEAsKnQzvIpc1VD4qAySeS
UnT3W+c4d0aSrqMTMeQgO6LIYc3QAGsqLoySCJBY8qCaokxEH93IF4+L/dLelIbWK43pzdpcHwN0
6HDK+sI3MGrpHcDpoRlsO3ln/QwC8VKX/8drI956KDFuCldhT/lyDaajoRlKZAznQWJhYZt3Avig
5ga6SyWTE/60UCqecP3+cphf39pT+2ISAum4Y4ClcwjdAOOSglZ0Xldr32Wg8Mau5ZiVAg0dXN+B
enoiMgqjlQ67sqHG/VIh9/AO3g+bW+KnHWB4iES+qChg64PSr9NalcXN0cuEt01eK4WeCSAtCLSF
N7LdPeuccm1hULFSNrQQeRzw06StjDbUUI/1lOiveF9+FzF2N3Eiz+N1DSR9aRiao+8QhExV+00V
7zQK4q2sFKxbwoFHb79iwGByZJoEztoMi+WRYPfXHbc8gxYe6sB/G1L51jb4TvwLPAHSU5Qkc6AO
gBH40IwVY4INWRIqXThHuaXRnbEH/Zb+2BmdDn4Vk7D64uKRRbLfMlUC2IMZGfH+YKuVmVjonwci
Wo1T4W0rbwGcY0f11mIDmLpApJcmTS87Gwt2S+B2V2X1HFJLev5cjJ2WXlFvrEEO24U+/IgUTv+t
H7rvuQXBgk/v4znXldO71loZOdE/lCBy9L3/IXebdRFdGqHs6ktGKvdCGdT0wLBHzkcC1vgD0WRh
qvkI90BZtDsA9rgEu9rYt+uoI47wnDIl9+WHZ3y5VLVSYGiiSMtpYw9pAcwjmyFB0A+AuLJJz9so
ZAMfEzqKhLGOq5Wys5A0i+AfKWZMTfcQOPEXNETVpfhyVGtpqhinLCW91z+FqJ54kGUgNjmqiLnN
prZmknHm8xgsjQQ+Y5OBcPCbcvsM0EUxiMNzsaYmRhQ+K7B/b+YMtSHfONNZYMzFWMCPzLe5p4c2
fYFAjQLMWewO5452Dd6uw89iWLE8NpeKN+/nYdtHzLqmaH9Aba2+Vlru2dV/3CJTIut6vf7PDmaH
eaq+nCOG6KOSnwEBDHedbaSLnamFWXPVK5XBLehSIfbpmiuF9CPuJ2Vo6hLnBFAVVD9dvLdL/3Bz
/U9VQNIRVh8XAX4ZbosxHA/I0AAu54OP3Eu53XKWULf4gk6PlKZYGhRZKLSFcqGMFPhlgK82RreV
w2aVFmqa0vMEEJrNzHrFGigDWHWChKPwFazVHbbUIYMI6ZF3cTvGGHACEfj3XsciuAZZP1mh/5tI
cYZPV39GZl/b7J6LwggxvH2x4bj3PAlaxZQiZKHfOgV7aIZXVFS/wKBScFE2Ov9ZaeeSTJaTwz6P
IeZ0/V6xj+UwDnI61zFWj344F8hoePkEczEEi4PNqQY1De1n75OdBHfMO6tl7oGsd3ayLx0fx54D
h08rzCo8EkRtMu86T4o98ZlO65chA2ShDyMf35zBszykXdLYwa3ey0ox3L08+FGlZ0dSvlKESeut
IiAql4rWRvazu/ssE822bFf8ymAnDf2yWbkkfUq4AFu3A/s0IaDuWKSZ+xTzKxeZ874bVsOjEriB
/YxyWIIncgtdVO/cUJjlxUIO3cKiPWrOYBCuqGgr2tDbzZNaYeBj1PqoWoZBigcNxUbqCZjijh99
XspXRbUTvofIUrLxK6sELPa7rkh/fejQzfSffW5ZGZXcdkKamqMBhy7wGHad2nctN9cWmqMdKxyK
4Alj6JVI7iy3gzVF2dmk/Euu3f0O4AA8a+0JNQntlj5/G1wOmFDBQC6ANxN7qlnY/ZkWtFPF2+xK
qQc/peZQ8034UGFDHR1qyaCQTpeF6zRkPO9NvX5o1ZeSE4p22qIwQokOhAnS7QXgLUL75O08oCv+
x+Q2QfnLuR8z6ibpjkj1uDop7eXdGx50pyuxN3qAjHU7bGW3tI5encQvHt5HfcJlvTLHp5TUNN1S
bVqY2JzWsqW+i/fHnblICk5DpVgblG8FYVvnXWgal3V0AWkGKesySbu2Rok4TnXoGn/6faqO6j9C
LOJs/nn7GTAJSlgDT6GSDeAaoo/ppgpc95dhNTieAj57IZP8vLw1+xgIvbLoIdfF0j1hYkILMWGR
kOMsP/iTdYSt7A7eddNs0IH28cMVkz1EUzMWQyfxEF2tcx+EkjEMeQgVrhDb4xHdZbR6e3iV8nzi
9Z+rPqPdSGgz4dfJuew3GasPwsWWrUZXjGIxGJqYrTun5uj/6DVRJF7veSmVI1xvM5sn255wPrGx
kpmRkMzLQmO5TTAmYawl9o6c0AmYybyf6pqQTejYswaQMQ3m8jJV4oLOl+S4Hgph5gMBDgAYPH6d
ZEuYK6gIXqvsF5hIq33iCieN6jV6N0uiFYszhq3odcpU46K7fHDlS7Yna96aQZ8/+Ld19eWEAgll
DnATp2auLztsG0JtVmwqNBhZlTda/no5A7sMJBOFWCZy6t3W8Y53AE1i7+ans37jXdZDpM9CW1x9
l8o2aOiqTwfLm7KV4tCQySC4C6BMYTGw7CCAAxSqKo5HIvb33CyjWP05lgeTMbgTkVF8IGFvk3Z1
WQ4K3ORhIroIAz3XyPbROTj/loXZT3ei2Lr0gO2Wv5wW+tPdSNF37wYwM3kGYzCZG2/TyP+TPTLk
MTuOOWs5jhNoYCDV86vQAfyiIjjdv0ZQe4qPK1zg2l1ARO1DZBmzj19Fq4LBgdv5UWOwGyCxTNn7
kX4Z3mpV1k792abpTEPyVKx/8BFwv0qlBQIFUsjWT+t5VsSQcIzwlh04d5myR8W1JHjWiMAQWO+Z
LsiQvcK996Xs4ftyqJmtRJTSvayGkhpsEJWq45vkUbkoENlzRlUbxy+gEp+x++JYK7n3xxY8c6hq
WJgAwZYX6245B23/fYMNybrtzNVOHikRgsIO8anfeFDkvQWt5wHPBaKfHb+2kSLPRTvHvZgZlajB
tb0nEM50CY6xeFJKfQwAzTk+Um5msWBs6i97JeTtUlF3Ub9LDh1U4TBaU2LrRUs/GWnNXEZUK0lw
/aTY6VpRYbPUSDkEXORcHk+AeV4JnXT8LXXtq143CrtucNPkWodcj1027cfoIkuQwo4nd1xJM1v9
40SdR1eqPZhHovdOSct1SdQvyOA5QwODuEj4ycmzSe0bfkOySIHFfnD2Zv3B3jGLbUWN+90vUnwj
++XERECdh2DMfHzfSt5b2LL/8XnSXhaCiiTs35amaQtEGj+OEASz8/j0odBfVJ/yH2K3ohIGPnot
CIqP9zJOjBGypu5z1Snw9oTlGAsq5/+D/++vQXHwuNMKfJLTmP3GiKcX0+Jo2dXGNMCYq8tE1gcm
Cq5D9l2h+lnXtJjhy9AZBPhm6bsiA4pmEHW9mQ+2x1mu9KCVK4yo8DDRRrxCSnB5E7UhwIZ6455/
yRk9VtdivVXTjjaUwmvn1K5iv+zqyNy9ynouhM1PnqnO/k/9UG8i6ZI63qWsaIZJyaJCDKmrPsWd
U2F5zIETtUcYpuHpRytdmjwN20J4HJ9pKehTsLc45hIXstZVykHGqp+qBv+osZmN91KAuNwU75Z5
48mgpRiBUlGKr7/jK96hDGJcEtW6u7a7cD3MZuOo+SjHziOZM7HoaKmXgMg+k3E3T/+cndWzm8af
zuwY5jpNCpMIFSwIVcOJpUay4ZfCv1VW6U7g/VEjQG2is19GWzYT5A71furs8cBoc9GXujKSFs1k
pl3LrGYxKhXowlwkTuxLokmaBNX/4uDwzUbUMQa+WdFk4soSM0+U/XCoRJsIWH+Yvq1qZ4lGDn7P
5bkA0O8AGoTIfmDHlZzcOZENFpREhge1U051zd6ccq9vvIWfryKehdq9JBubUOYNIr/lJc+Vb45Q
u/ERJmKKdlG6MWs/c0AUaItWss0i+W/aZfZKuF0rSxpah8c4eUpDNjhfUHBSRC9v4+vVlzt8ZmDO
dSicz/puXXLu8Khpbd/61CRD7OpaK5pngIXpukyQQVXpVPtYCCB+PZU0FY/Ue6O+qP7j6zMVge7j
E9uCkzoesN8x54j+c2Cux6k5DP8Zas8xgcvGrvndr/P0HnGcxOur8A1bbY0JyMgAbnMM6Qk9U+JP
ehLgwWx4gOFp7q+AWDEJL0IVA3EgrCfOU3mP2mG8Fq6OOdgktt7wuhiye+hLwe1/gTtc6/0rSMzC
YV8DyunPXIkDxgriemHXPdCKoQBWLRc4T0ecWOINqhbkBOKkiQt9AfKdwn03IjlwEIwFOCKQWVJr
bltIJoBNlLIogITbaU9TQTJgT0HxS7pMjVcFFw/UgHVtwQ0tqIrPM71ebV16EG7jA87OSsScbwEc
98xbb/CvVMcqo6Yx/naoaV6mP8FQrxi0xUoiiELPk1eIVaeQ1Qbwx4hGvqTZbFZthsM/ct56c3Qo
9Bb8QPKnEsnOl8Yy/VEYaEK2VqqLZV3WuQiXRfWQUDu+kmrWMAsKkeYo0QUiuxw/LEq+URrsnsFW
fV90J4/MVUaiEXqTDQ1o2GwXmSJqwK0fXZ/j4ZUSpGo77PK77hpWROuxO0Af0nmifQGhn/agQv+9
gbL+MepcVXTgJl8KWqWk8OFJDT1uqQuf2jijHmCsDllZcYrpwQFFiSoPT2wa1O5d9BpvblCK/w6l
dzg3Ph5KNl0rTqudGhXoXJPl5bJLEc93ZyUoGs2jyb8jPYtHY7Zb2cSHSAX4mQgZvw0TdNbvOje2
gtu89mzPGZOGl21ttAvN+XnSm694q52CF/X4czzUw4Otf9GOd28MYG1qY7vEoWg5Mw1vCsb6g5lf
4cDy6w3k4V0RKiNphjXBfE4FoZG+Uk0Jl5Co8rY5iK15yKT1c10kkyPsRi9N6QfXr/g2qj2Jbeey
N3LNuauzNkOVM03t0vaKglgF1dxDDgfLMq4d4fx0v6+GmYstB8SGwW2nwh0t0RYsov2SmMsB+2wT
FTmUDxkwAHSUXd0miD5NF8AVmJancBi+CHVREcWtalpTUBQhpWJ1CIiwCaN79cT0H7Wi3HmkBDPm
sXURh08jBFIowhkLpYc2FZcETzRPs7Hz2UdJZsd+nwP0fQPq949/sKm9f1kp9rIM5p0aS/CpEdkI
gws8WHb/4UhqoNU6RXq5V427POiqsCa9mqIyQATygJjfkHFz8XxYjlrGvT/f/VJYMlkKF0nDVI1t
FB+HWHsYeKmmWhp9l3Uxl1vGR8HYgNmBaFke5XLWYMZiVca86vW0Q6XvTOIOtqI8E8TiIhmnt9Jf
8hT+1dmnpbvC7qZxWbS4d6JvnRkFCQpYmPTkn4WVjCOTQxZEVVb/ooINxoN03EAacGMhIXItX/6v
spfNRc9+FycLZrs+9PqS/uC45NuV0pr3z7X2g/JRjHAe3czuzawgNo/jJHwct/ha0Z1aibXu+Rh+
bEtDMhS4zCZlZ7mzyVyyCW8GCpQl98VQnM/Zko6HGuZpit6NUfLj3fPGejD7XrxO9werZ+YxwFql
qiwmwm3oafYHXILO5TokZGOkTGlZYSbHMg5E3GUDgDRPezOA3BZPnee4qnGkdxG15DmRJqmVRDXq
mh/YGRJuvCWAyiberssi+Yy69LN3IVR4SK+XH8I/4t6uCY7Xz+frYevSJNk6WiwGQOjjp2M+Yytd
u1VF/Fzm2uJDSAkVzKfn/nRylNXezQsn8jqLZeBnI/E7TSYBG+WWag7wOBSn3BsT8u9Qp+i/YR+T
sPriJ8zRjhXXi5ZGSWjn8M0fzrvzWDWxiHNaGQzNOtr5y9/sEdEI6xQMPwXDa58BW6jAgo17EWnR
vUyxtWbTSyCia3Mf63tq5XSAe4/zoy+B9k5bJZcpEoDu97QvpchEFZluM+k5tbuoZZO091AJe8sa
ivGzHzlKt2z+uXIMStTizkM62g8jOzPpLwGvl/5xx72XX3OkvZVrpzE08DeXqlkIOO/9ToEgkjPl
EEv2sEupGkQXwpwaoiMbiCmtouRQ9tbas9pbYgIv9tkJGkXPMzZTFrCCUVK0Rzg9WSSCRTl1vhQ2
mzqFvcUPKe9xADwesB8sTqvNJH+r0yd4D/tn3pqXTBrVj50r0hDOFdBQzUZrX4lhbjMp5f2e4R24
CAzS90ZWLHszlZ6cfy8vHeJSKtfIl4qDyXYtzlar0NFvnGYCGxrFK0fCuZHbLfK1BudU1bRtlKoU
rU2E+EVpvSxFvtBs0FCMYtcz1jtBLT7Vf3E3cCmoG35QZ90p9rFn3vJyoEAzPTVcaEFmtfBL8TEQ
F92GyIrK8TbhvtnY6Xk6AtFewnEwCupgFIw4E/H+zKatGBSmtTyzMyV4T8S9TOuP4KNrmaVtSCLH
fc5Lyuy811cQs8ylE6s8f0jr/xBAG9OxoFgLfHEJfgrLlNq3Iwoj4P6Eo5f0V6qqsJEIFBjyXlww
WXPUIZqFfhbMfJoxTyiArSQJnyJKrkxFlC9zWvweqDYe61tL2JIfSM9eQVW8OCND2zETrEy9cPzu
nENCy5VDrzqSxIOlGFgaR3x6ZzkHAazhqWpUhmr/mUMfRLK+pf4Ehnetzlt4hSg1EQUrLKkVt+HI
3wGMERPB6f4jicIGolxQpQIQKPHZuU/XHbMq8nyLilcL7Rs/s8O/VytkZR/cyI4nEk9a//7upIsp
2iKyDhohf6mGSKDRUcWw0HA2s6wXavFXV2U2fSPz8//k6urGCqip+JRVGJqSYQTSnAPLZkSqYEp0
udq8Qpb8EwmAl/ZwZRL+bpvTNzZ4XxXfPCGV8of2lsHd/6EyZrSeR1FEAlUh6e9l9h/SDlYRkGYE
Q94mfwNsN6XoRzJu3UaNSsYeGaNpjGlzR5I5md1p/3k3wNFtwah8LhdqIPeRopsGoIKh24pBaTCc
NaTiD2avx4v5kF9Na+44oBuyRqjwqn7d8t9T6OjsdN1LLZuPb2oQmNyfg86fmTzOk2Q/707oWGHk
wBgBXG39MOYVEEDlRAKwHU2CHIZkbaKLcRmnUX0Xzc5C0EWFqM9waq0pTufrb/zhdAcrNahgod8c
ggt86TQHg9OvVt+wc1/Aa3G/F2nfEbm2dnfqEKg3rxB/4wsowpIdgRqzosbpgKQYZRZXbP2J2G7N
x4RYkAUxtvNoVDoq3i9OXMMA3LHuxvcn0BlO9hkrynpVseNUzrW3MljVbPn3eiDwTucXUFtT1En9
YlQtgzvRTlyeFVY4JqFkstyr6V58NiG3ieGGdq4wl10+6wCeBRabGbi1iPfiU/GK+JacEnkr1KFN
viqQVgDrCals7FMVhpM/i2KBJ0HMAoBkMj8+I7wSjiiW7kQg3buBaZS25ab6+gHCsLeBSlq3BkRs
Ti4P+LVverMXRsmYqqAgtkK7TDCLS1ZAw6e3q+rGIABpWSCWza40pAPc0z+fEwvYWV2XtmeC2Pme
YsvifUoklS4xeQC6CG3K7N9TlC6SuJ/jcZ9b3HFfzvHg/BfzDrd7XqhcmayDmLYO8DnJ2F1TyI7S
iyQTlJ17eBCbOEQ8glmkCXQPjOPc6LbFfSdPwAvLmXegsrCop4o/8JdtR/7ghcms7/a13TYRLLgl
FIEjyeFxzSitmL9sgmpTLpFpmL5+sLXDQx3SYJEkgxJRncCwii2+IAdiurzUlZ+yNQq79t7gY91v
Pb3LWcH4zl1vXOvkTYXKV/o394oqP3kSQe20EfeU4mgKRYrfNVFcnC3WhI5TVYRj/s0MYcR7QxML
dfLln2W3IdEtKtxXe6+6fYsoyjOzLgbS+ewsi/3Qtg9pRYaU2UrJu+jLpZX6UcbMKMq4/9DVHM0k
49/6WXksvRhgUeV/eB5qAgX0/7hjCesHBaihljcR+q/19RjCe8yf2VAPDhqO6Fa1Bac8A2RyFWQk
T/Pg31Y1ZE/fF8IgebKxM065NyiqFqiR0MCG7dsP1+kKgRwsF2Z29QK7ifebrcDtGzsX5WynC7Wq
UhgaSv8DsocxdTxUMQmnRjmubhWve5ZDVVOyitsDW7EE8NupPqhYQWYzUep70RkZcnJQlDtmbLzY
8ChhyCvaR+xDnIoEa99ajL4BdGhZRXva1KFvvqgHrZcnOUswQ/b3zc4FJfLgJe4TkK780F1T5nph
yepzcL0u1i0uAL92Wg3JlUVZmbsCAEzvMAoG3Wwl5KOb10lMEHbSRqC0nDSTstR39NB+ndnR23rn
pEH8VjeLGv02KKZFBPbAw3j6VPiGJJddekXvBUJSKBYxCRoKfIrDcOaRyjTje487Z1uAnsSlKH+7
rSc2mJSyMKUMVjGXw1UdSl9HyObtEnN486tqEfOrDcDGF+qPUHjsLQycZlzAWHkMJ/IqImgX34+M
+VWx++fw2McFDhMQpj7TMYXaxlArnD6DD1k87VYLHQwY3+DaB2CglEGVCriz6+kajxD2HUOze8Kz
kuFjhwtAxvhZ4emlzgYlwMXMjfcKym9hShg5XhbQt65ZdO1WjdtFnfeURsMKWKhnuvEaDZYDyewg
7XyE8l0F2SauenSse0BycaekNLi5R3+uWoFXJ0Rh9LqJ9WWygDdbpajS6hUCXF1RCjaJGaYtWGl4
mRWlfxoOILIEv4hNx5E+iVVLkq0ov2s3rQZwTnPcKqmOYpE17aP64tPaJwc8wGB0VlfdcBur7l0I
s6EGakYPtFtUZLUII++so3wfHH7h+2Wt7jlYhwPVh5FVwnr00mkCWFzROpafei7/+vcqYAOvozEK
dbq19FwiGerOBw9tkMnod9rfGhElfO3+5SO+ygRE4m0A1TkW0rpzFRE9Yxmup9VDwAoxjDAtEXXv
2lRh7GAgN78vhivptAEawyrbYO+R7ACtkVbnAD737Y2a6s3HRV0m5/yCaKLSXhd0C0uzN8jVQ7YJ
ztJyWtuMEUW76PQtKn5CJU7SmZmCsF3W6ihYGt5vjRkFwh3eIKTGw7hkkHA0ni1kcubUdUpkKVrk
YmDhtsvfNErEfm17WypwnIwzom+1GQ2d9AqN50LeNupV6QzfMh6Dl3UHD1mERoqZx2SuTe4oaP1P
bn5Rp6JzmXtjv8zV3vM3LebIPiK7dyxTJmBt4Uwk8L3bGxe6ushrq4E6NsD3FHM2PKRjUydAMDnV
bwBdrGO6Lhyoen6iFHKTMUOD86rl6iCUbAgXCrGd5NVKyYpvdzFxfPHtvhnM8+EVR10Nbk+YBwZw
blXDpr5Ge8O8qijiYSNX/v9a+bxiQSg8NPX9j80A6qAI5xTJ0Np4C+3TXsbCY65I6bcw8Og/BN6o
P8uga0/T30tR9XazNpP0VhqYU5yEkvE5keC0nOGpjGE5NuMbd3AwDWhIh7q+X9C48hDy93xqHuDL
exIFXl85fxQvt1kJ1pwfZeLWFPmwKUxoBxt4Ff0PlDBrVc4sNBd/FNo9UUbfQeeCMAZ7UMvWkCsX
sPpX6Tm8FhyTnEIfJd2JOfNQbRlHomKr3u1pDrN6/2EsBaOhgrZbFEt9MFhNs4gEAyGdYqHd+095
mDRi9SnGEWMUVjgL4O6NA/2T9JiszCvOzPb1utVewzRWthJ7CMNC+pdbOZQCsZC7hNHnmaJd7uwI
Pj412BKRTKY38bBw9CYInJ0q9qnkRvIp6KIoX5nP/M23XIt1DpN9bPsQwNh2+/cl8gh0KhJGU/Vl
VUdO3CIerFHuio3iv5tqz/njeaWv/wEXqnpHkme/MolR0hycg9MC3DaQ62koO4in3PS0jR8lE8lL
ZPDEW4E2v4GSbzgJjxQhcqdFHApmS9rEwSiWCaMuLnwx4e44ak6jQ6rLn/Wlld2h/XLUyVoH963e
vIFwUl/nw3F7eem2bdsVfYQOXLBS9TA1D9E5GsRdYMJ4DzwdNWrcmmA4FTyxkLqw5DDy2cVYSG3A
IQQiw7+PhyovuB3ghnCsN9+yyiGQXhfJhk0gmMkYiDYjy83Rnp8YKrgqgTXaotrLecvfmaDwyygK
WN2RhYzvo4uM97CmRhECIvkyuT8IeYCjs/xpsU0ilgcROlsX8Mm2T1JXHgeGMmFkRCAQZ5eTwqE1
GjQ7vXJMy5dQUcgFfs3I6Hb016xDC8LbnPoJlIz9Ab8EunppNgL1LudOAnpOqXtCHoAC4OTKWmL4
jjGxVxTA0U6h+S0H3yNnIRxYLBns+KQ6x0KaZ6fVnWuwTmwwnYLpngB8o+1ajoq5sumVVpqjnIUR
ugM4ndyTBOyBXSJvjD4kZ88mkKqxsgFbHwUM86XJfLy7UgiYXryyTRm6wRu3yY4oiDms5BPafCtV
ERLpsuzUmoh07b0IuyIeC/fw+WLZu35TvxeNqHsyMI/8CqZ3q/Kps/z7YdYlHMptyphpfHGqpZoG
Qxt/IuV4ZoWF178LjP2nT5JV88AJh7QN+FTLDDUL2Kmv2eSxm+V/u/o9FbxsS0alIXym7HGG25mv
ZyGdOiD65tQR2n3MbyRcIRt9aPukvF3UXXxZTbv0gLwSlFfPuxxO7f/BaLS8BdF+kkUSoxokvS2j
VobvKu43DqRdFGqHIRnP+tHYB7R8BAL32lr9wYOe5swFzdtDIbq813EiCOTcY94atkUCYa5sF5gp
G5c8HvYMCo0dAniVTZgvEvz8gxXKlO9y9DTTOYH7CzXYLZRgZQXz9dNUir9rDxYmOEH08caOEXiz
c4M67x3S+IfnInel6BpklG238cNo1u5JCUM1A/ycnU/3QA0IaHbeb22kGp/miVFyEyfxpBd+1D7C
UySuVs+0EP6hE06zlOWypbIfqF0FtFNGbB4Wzr4Nd8WRaenEzyBVjIQxQnSKyfcPItuUh26832Ue
memFxIP6VpJd15UflMDQeh5w1SRTAiZ9E1DdZfZJ7bvBE71SnV9Lki0jW5pAPwryzrjI8FmGpd4z
e7bQrfVBKRTzf4B5rfI1iScHWD9ORhZtSZT0UbLZOIFQnS+rEdyARpjL66VldZk7HdavHuBul1VF
0J1ZJmP9AxkxGzOhXZLWfOs5IuVdXfc0s55p0+hy4boG4QzjDFOLKlVhqPOAFhPGda256gwQBv92
7QTo2/pNY82ifj+RwlIf7OFg1On0c+aI87XdzoDRzeld8MNypo2ickhCJAvu9nLO51d+GHlDBHC+
E5aOLXp+EUZg247N1UVWnvFmNBWqL3iQx7MdLZWrx3d1qMQfwvaSLGQNlgk2bVPoNxJ9UtcqewZb
JUzc8gQZNf9G4lud8Hi2on9ENtCElTZXefZKtkG0K+TXJ6FEv3H/eO9Y/9g4zeBJkMiiNxj7TY5c
nT+3U2NU3JafMxbAIM0O/I/wVMxi/jiYUnnOfQQ9/cpiWZuPUq2gcfq9PfNAjNlNVRtryo3JIjQK
78EU8RxWx99iDOD5kdwGw7zAHiGinxcvWbhvKtGght7EVv126/KgbQOajZUwltVcgCZIwBqddT//
yxfhVvqI1btuqnOWviT4DDYLsVcMGhsk2W56rgaRC4+9QHNV6k5ixZ3xm372J34JjxVTnk1JACkV
aAMnSeaB86w/ILKx2amgOfmZjMCPRq2AqvVK28cATWP1uXaLADo0dt609AJgCR/GUafLh+1jgLAl
hIZ6PJ+LTkEqveBT4CxQ1ru2ZvkXyo+FuhDvdoj/QC+eXcjbbu9uWndU6ZNHHTvEbmpwGJH7ukb3
XwMOJL15q+dbR8m7xZ/Blwv7Evyn04q5fc7UyFRiQ9Gb+RbBwy0U1PpodPkxizyBOonmAkxzk4Em
9wD4XLs/yXDz1cMCt+b6/RRtZIFdWIxvO6KPGvm0B7MvDXY3alEHlK1mPgjY52xKx5ItAe3wAhXR
FsuQYNsWHlktUTqHvRtj5fi9mGZ1IGIgRvAVlZ2GZnRmGK0waqDd50lrvZjgxZ0CrX9ISAYMXeoT
3RcA5iMA+QwQCLZ/DTmAPT7XL28CBpY3B7SUgbLVifM3UCdmm8A3OGTT/yzhl+DjKTytCsT9LrJc
TSZXvA4rO6Z9uq2oVprxOgX8R4QWKhjiShJi7+7+y3R0z7hZU7MNfEqfqo0KAtKjag3nojGNzPzt
xJdjYfVivMbJx05VCwuOgshDas2gjR6/o9+s6qArAv/54sSsjvlmQt2VEM+gC+3LrlMsjMHeeMdt
Al86aO7+EK+aSuSAJJNRkC96JN2BYBZKrL+QvBmQNgkjwZ0ywxXF95GXjTAaNV04Z2UCZqaizPct
pMte3No6JC9kVcWU3xzwY4OXbQ6HvBpuH7dwJQ9yWHru39qgbovZR/0I7lAR5coxBa6ZD67fsXpR
QCTPOzXXjaoyrq9EPrenqg7frBKRl6zXUYrj3d6ie4+YVgU2AWBmkTn+dT/rppSrdFzdYbPNpj1G
tlXXJ9SMW80hYQOGx0enTfuYxa67wIAmr2RfbEqQrwPkjykGXYQigNiy7hniczmeEgYc6LmofoiF
Q4jaW0goiB0L0FInw4ucAIjBJV40P2dxEG3xnK7bDoA04vAX8Qhxt75sISkA/6LsEWkFEu5ph7VZ
w5JhJZnA2HqHuROoszBspHQxFxd1GQxpVRAikMBuoZMbybiYt4pexstiTHzlHJXGxDIHbX6ANzyW
KqwGr0+wtdBRVTrIaP1zJW2UKz3Rok8dsotShdFB+UjFs2DBJjsr7LFGqB/z0gluRcXt81ilZXAY
jjQ+ra7k7NRXt1/fvc+Tug0QVrSkVRpx7Jtybp+i9ZJJx7FYQ21qDgqoJMMVibbednEf6CiHTXjh
OOXXccT75fB+PoktMDLYuAybFYufL3TvkUnatlZBB9r7b/SuJi3kf4Z6n5VW+8Ak1CY6Ih7hyzOG
3FPQ4szao0WneBKeSMEz1tenyleGEz2EBH0oRxiV91MKBiqj798tazvhwDvMrfFxgOkPjyIi7g9G
1UvEnCesiBBlRaSLHJrmNwCYiFnyKKA3fxHjxhftASsmQSFpkZNswMWhuEq3+QYRM63u6yyyxkcQ
JRBEV63q9u34xHXXRKdqvt28dprH8daJwPT9cnJBmrpWQxIKgw7GtbkWl/4fLLyweITJxFoGcYwS
tUC5fDhpEPZ8VbLsIk4pmtx675MYbQFXdcYSczmRfoHaRDeZeIFyhr+LbuLBbNO2izOnl3D+Rkvj
sCuV+OFKg0IMH5w4F4HBc6J65L/yyVicyisSz9AcaZyHSNeMtU/NhpkEmpZAUpPXS/qpMX5JYyxI
2gUWmanryff74Ki03XtYYMgoeitIWANbIGzyRTa4a+rLIVsDU3+6NBXHIGDdWmOk+oWwy/HneZYI
YvDN/wzCy1KSNlRxfyF/3EMBSzx1quzDEhzOowpYUFFrz3Ng/Ppcihz+/rMTOyeDbNh/UE0jTUv9
oHlxNXBNHqXnwbQz7/s0TkwavptbxbssTSPHBoMJi69HLPTggHzX/PVkLYNrsx7GLUtIOcC/bToD
Yym1LSE8XIwwxwD5SoZ6xIAkXlcAAqGaJlf61NtfPK5IxjJO6hyPwSl02+l9Q90Qt+jG3BfnPziE
trV1XpUumdgFTClnLQZLlVqEZgnbYkKFcN+oBdOwJm2P1/x3Wd1TKGguxplENFa250K/HOHsbtXv
vGBpShmG6hbB/hiWI13Oj5qD6br4FCVs4F/Nd8KaQmMGfnNY8hFt/BsHl4rIU4M/MGii8GWy7RAZ
UGg8qEsaPH+KWl2ccKHfVMESn8EAIlvfZR+J4Undv8F9GDC2TII3vUR/L77rKCoyqDDdf34sftMt
eDr1ItynL8MWsyrJItzhsfblUvRWabvc9egftp4pccanr2BanSNq9jSKgMa5PJL2xWw2VNbX/IuJ
Itct1gnJb7UwAHuCA/fK+bh7CL159gRtVdjxaFRpYGCr4iJVqcL10mHN0DEvMe/oWtAI1dbsxobn
y/h19LZpMfgEdeS/L4k3fHWhfhRKZeK/dCYszDOxfQxqb325oKvuZMa3QIIUIydsoExgdJFFvfNt
1BfHiloE4l3g2BF36ceRd6ZxX3UK5Pdd/4XEwgOSEIhyRKjsHM06aPDmrd8uDvpx6ehlQ7eXgcFg
ZLW4FLmDwPHP5Yal8x7AItiPVFz/feuSIoOVKxzLRy8wAjRnfNTRVET0NnKS+XctRIW7SowqmVqy
EKVXriEpdZdYxpaHTiw/W8wgJSxMMJJXRapjx/6THnn8vYEoEC8SA+3yxaWlUoNum9lApodxjBWU
hwq1dhMAEXG15OLwYF6gmI950R0xn+Jds8GdqVJPF4lVIhuXUqsvaJ9w2K2Fh1OF7BJ+6njD30Aw
/Ihq21aGLva5kPBNjV4nQRPWpVhnBxR3eMh6hSdIcwJGcH/FcRvpFu4Rgxt5c5QI4wSOKDqOjhW9
F2yAdEBQDK3KjAvMJ70y8xYPp5bdT0uVEYC5uoxrldFbTHMsSVjsujbIIi7+2M3vc7vjBo6vxX7c
X9wSWcPv5wACpX6A1MqgsdZgD5lW7as4l7vqkf+N3MlUA4Y2tANqWZZYLjBDfDsWIIUSrko14JUA
YknOqsGxg5RL8UdV8GlxnjAOFuLnz0iSHmj3hQ8Tm1tHjOmGM7eCGLSlqWYG51bwx4gCQbLAs7Ns
MYfZz3pVCTBYuS+yi1+hyllxfNGJkZWosqklpnw+t9Zw0/3eO8ETaUWCmlXlXnMqeaCAuJsxmECS
qZ5dxmtWp93Gz7n445GDrwBSgBY8+zubx6FdKApZ981a+IY6lL+KQhFFFY+6Gpz80NLXUKq4mlwc
uwN3H1nNH3YCH/y3BgBUUXSxUpRr+YNT2RpMbNAuJfDbVLuGPnoDuMiybltsJUStIB+Io0cXXLeX
Y56YnJgv5yRGa7Hfu425Ut0ia+3RLpyHcCC5fewXSOHibmslFqHq8MrWM9O1fQTt0YX15epFQni1
i/xowsk55ZAoUX9jJ6YI5HvArXZgXR5ZKgEwt4auMVY8GH8+4glqlN3QzuYdaZyDBgEAYsgAyXxV
/Xxzx5QRlFAMPGzB/TBeOKPgl0UJ+ZgSv2wLMOC1yDmfJzjh+Ydk/zSEj35jXo/qaHUk44oswjOd
kuRNx0NrsQr2hzvS3BXmMSC4wjCIvuQTytQXX9/g68p9VGN/wUzPuhv8SLTQdu08nJAW3UDEAPyZ
ir0Pcf15fbMencQa3esrgqfBAmi5E4KGdEjUBRzqMXmjBOVtbe0O4nEtpWShul6Fri4Ghe7+r41E
KIp0bzriHLxnnwGQgnGugD4lggJyDh5VC6R8Mojpxq0FmFzoxRRVgrckWWrqZCjEoQa0P7kvUcPc
udul0IPd06FuZowdhmH3QAM25Zlt5ciCGtz9IK4QQHALpTLifuZH27CHbzxujFFnbZKo9mZFpNt4
cBfZZ6h4kUADCJlTJw2dcntxLXzIFQzEYDCnFG9RxK+TzXOoJoOOP2f2BVf310Wn2STuBDTmVDwV
EjmupqsWXyeqPjAplfZEBcOkGg4A9jHNt56haiAE7Sz86qP2CJSIpp+C3/dJMMWJoZPy6aIW7BKA
ypK0Zcd1/C3OC0136xYtZUB9CI0Wtrig6iscm0/FGn7+j9wX/9drsiaO3/OOYi6e02oSazuo1Vr0
1ZLaMUmv991OJP8VL5V0fbDxBUPBGpBqz+w4dw5XHOOp6pkyMQ1F3ccR3+OkHQ74+81u34yTK8uG
mbEy5sIFaHUUsh/sEZoHw3dfBki+nrFQPNBM6K6hYKXUsOmeUlUMYd1tE08nITRCP2IDX8krrYbn
x/iBOgMXPjginu0XjUGtVPNEXHA3KwIlZNW1BStx8xmQy0vxqP7Gfg8bzi1az9q2DYB4MkpTw1T1
5cYh3Cxcw8sLnia2pfwbmz2mnOy2qXOa0kV+FLzrhVIltEcJtF/guR5R2wiOJyXrUxVxLumtxyiW
kAGw8kb9U33o9ggNwtKmPUvtxdGo4AbqHzgtOJavwmBN6SwMoe8QUCcOEDhiVIwEzVyzVPSpiFzQ
HWNGhPeK7cm7PedkBeYWcghnqTDrZDQr6KsrcBAfGbgrEZfZF//jc8FLUq/rY1shjELF3ff/ejUF
2JC4M1z5FS2jXcRUsdAgcYXDeGKfeTTLNgOSC32yw6BuN/2knNVaU1d1IP+N1XvrvGvAqOHQLm6V
zosDUpDl92Mv51LdfMMjUCJV13j6IFP1YJHdaYsYhs40XtQkIPxuj55h53uzECfGmdQ2CkZlEP1/
vGc84+N/tOFSRK1LHJqDJnYq6kinygb97kNeLLC+Jf34LLJY16xwH86M+aVY5+4HO8KK9oUjeZdO
WBL4AVmntNtuHWw7vmE2PjiUb5McuKn+qlwQWoIMSWsz7ZGIkpbGCuypoazEzyBRuJJjJ0YWK6sP
grtDwwCQcfQDBh/uKKwWur+RBQJsUdvGmdg6wqXiq3GWwjTgIY1FLRPT2vABcq7Ni81NkSpEXOY4
vbFXtqKoKv08cs0rQeMphyL23fSa8bWKpmXLsPnoKZB8+6RlunxFPe9lthJ/aJ7L2Ijhpx69vXei
FSnImIC+k2Q0MYtmdSz6TzUFpdf2re/YlGjV3KG49ppOAcMEzl4wJemLhTJkPhwNzFeO54yzDqZI
iO6OYI/COgyE1AEGE0e+Gf++Uf4usP+aC6H2/Grg/q7gnYUzssKXrTkSiOVTa26X4/Y3C4O3bCX1
arPmezK2i98PUJNYDmouO60t2WiepY1Xx1/ZVBHLY7FPynNr9av+/Qv7KPUIRsIYHz0bK/ar47Ge
jmYEoWgK36OjetnO6Gar1YJBibTjSgkwRGzvIWrnQJQU+blJWe47oAXsb0iKyD3cnU+uJmr9PIiQ
XpHGIQfYKZZCfdQK7bSK7h6vuZQGpfa9amV+Dw+pen3pb2cvymfDA0wrduoK5i42paHOL3qPd4lK
ypsdSME1rkvkPuN04iChOgE4jQkbYWcAx73RsMGhf6O7nemlnwYET1dT3Lo9EuunLGPVba317Hj4
csp6jD68X61Uoj0LPXP/HfxWuELMZZArR8Lvc5b7wIyZK5yE3JvXKeOqlfQ3cckTxTNeLSg+m2T4
O4kYN6SSw6MxOOCLjDa9/8397b4DcpgmtsdgQ7dd5ixAS/rlycVQy/KxHNzzOkidPX753pXXQciJ
VPc/1dp3n2rZdeuF2B8HiPv1QRV6vljnyLKhiQlzIHEtDP7DY89mXE2+7SXwlPpN+uDFCLcNPfaa
Vh1kVtEST4MX0cnVI+vbWBmPd1adN8Oquf7wNY0en5cDxq2SfwpJo2MMBltU59CzmnOBwAW6uCaC
KMUqGRmss4mXyUVBDcxJsOsXo9q6KlsqEsxrPwpWhFYdX8h73SJEvFKL2MJlOlqLlz0W/qDn6OLX
3YDyOuoj9EOVNtRBYV/3oW2LhqmB3oRByQ7lUUSPt8MD7oXmltYpZRXu1+Irqv1ZGjJ9rDcM73lD
xYWgffJR+GdpCO3XyW55CS7QCnn0vgytiT/7dR29SkeMmalVsnXCk8JtctO5T5yUmEhw2KtVYfUc
930DroA1q5f+I39yUtaR88CktRKi/5PTh78qh3TuzlJOm9i0k9e+H8EgKtMUqPdwDbHImmJhapn/
9Bkb3jaNICk7ThCs5lkrPCnvj84LmzQ2KzfyPpMzY5lIAfqjHh2sEorAxQXzyJ/xskdRXVTd3aVD
klF/IkHwKZEC1ItntZSzJxuJWrTUC3bSH4Dch9MeUo0Ph9gLmZNDJEZqPIv+lMl8PJNlPyXOS8d6
0+q1DiD7U2GOLcbKTqRxDvcRwGD37vs2vmjF2GvCyedXomELOSQyYSSz5p7te68MzrTQ+Nc7m7fn
8B5mR7JN6hxYg13Ajopd9lytPF1MU/2s4d/9TouiMJ15INfxPJOOGPMfeiG58P68g+2tsJqNeg0y
dciF31BIKbJkCZ43LodY9o+6H28iZrib9oObmUj9eJ/wuCFI+pv0JQSPLLESjpVfPm3rvdBLZs/R
EBGNbrgin/014EEialCecG3M1RFi6FU4aPgoEx/HcqAO4OKnJXowckVFVczrj4V+E4d81BtGIm3x
SEaMj6S1nHU9HOWECEeAThRE6mRrFY46NDdkBgcLt0kfAHGld3Zp9E9Qp8kLq0w4c5Q6ENqvH2DU
gZTIE0QXWI37tfePOXMDTpLUihDu87dwQtwE2QR2ezBWBkNV04mxQJaS/k274+Gup28R+xQkeaz4
34w127Ml3M3AXbMwkKiX95yB7FFQwK64pwDmrBOyA2ibsmUQngHGpRUYrVAUxc2cTMFplKZfAUXY
meU8iUl47VC+GBGQZgDVd2pacjusjz36Rtqlc7AVEiSG8bsP6fZ45Tchjdn0aTngIaSFCiKLaaZW
tFN051sYWfI7Ppwo28XUzmXq1Mf3OLOTJDsd6QsRnXTVao/fPFzzp96YTuOmLLlSTQ1SYmJ4oZ6/
2cLYxdjLLrH51rYV5xstSh4U9HGpYobkY9btmgq6tI+C+4dFl2LGurUbXudXCDGoiBNFbRGQWu9s
9kD/bJcMKf9s5gIYajkMDCl468h7ILFX8aYivyrZmH4rggMOCwro2+iAKnr/NjRnnfEf9OyT0WVA
xk6ZvZnJjsKun+MBq7f/0wBG5/oeMxQDUQnSft7HC+sQclft5PYltm+ycvXtWNdzAE7SKMHNm9lV
5WshOaagqSfxbV1HrgkGIOXlLR9MdGy4rHADAk9MuaEd4ooL6KtXdS+ZwkqW9tvCZZoYjNI4KpWW
uoNUJUwKjmwtyHvMVnGrW7ZhAC0x6RThl/xplnDhgmyKcJQDA7dtJlV/rZggqSDRPkXIlw6HsU6v
WDkjfHfyrGHTIkxFLrRluemLL9u0bVFSfMLREs66wE5uQJG1awsZyFsMxzOFDEOubICiJNjgVk06
l9+YC6peIYZ5+0cS1pc/axYUNqJMGbmytKCxKolDLOI2Rz483b2m3b9bbEYUQQuoTyNWPfgksHBu
gOOlL8tPr6lG2lBzg30kJ2Lp9593EkBlWf7uVQwgKcA4lYCetLD+j/d+YU99fx20BtFNyUWroLkn
xzIgsd0x8+sDf0b/A2+xPGVRs9GwDWtmXwdzfk3z3dyIDXowpRrxDpLgHVt5Ni818b4VQi2aZxri
iNEzinGGUwTWPfBMyoNRpjP2o9jTpUnpMogle5z/auHJiGjUkHjOsKLXPC38D8p2kDZ3rWPJmt7e
csJmVtUeutqmD6jOS5ROt02ovC7yy42pzNVD14hoNW5gMNz1JVHNSynXGkA1tUwqqqdq37YHsNLJ
BSEL0Pt2VLdo9EEFHPTg49a4AMKxOEfx1jC3E+H2dUWvPO5tgqYwbnSb9N6x03kZ25zTunAHMnSF
XcbOnH7T1q+k+aht1Cfvud+Q66Okty8vpdQ/pLnMeSc6Ln7+FhknVm+3/6kY7oNQ6C6XVvmY7pcq
v+lE+ZVHCKF77iW7RU5k5Joo3QdSD58yBme0Y+RBEa1OOu/P/FXyQP0jOifeA/zgVlFKScoK7M7Y
gcezF3j6MnpOrIiAfdF7Z2b0B/FOSypcqMRhD4yp9HU8a+gn4sJnCGz3kuWAacehphv/BM2H3Fc5
ovIy5iIXuvGyTGU03LiDVHCJyXPhAreB00BpGN0JAPsrSUKp2ziVPCEnFOJPU/onwXD5FhxUPc1Y
V21za2xQ4TbHsE1UgbVGJFIsWSkZ1U03iYSbHa2SG8Sgi5nuySBCElq5qBvbELp1XcDYxhByBF7p
a74939gCLgRLXwLIUmFfNA90HO2IOvT8BCYxd7oID/ev2UFWFAA0Beta/v/RKZ5gkckf4Nx2u5D2
2rWKddx0LYKfraLjaCCOaBaVC8EswLUP5GaCXDftB+w/5JILZP9JIMo6ECH4RN+5jsMSschPQ3D1
PvKDPCRJSMk7nHBROuQRr4NPDgB8sWLijzZsYTFVWPBdouLFuOrD5C1/iTQ/1jvF6UM7uDkBUCyf
dKcqSvmuRnzz2fDlxTtl1dnuIcN5yactAnPHR8Li1wz+4BJK2FcauQTg2iAaYsTC383VK/9Mn9fT
A28spMOtD9H92PiLLIgbebItLL/M0cUiZtpkYDGoGBx7WHkllESfplYxWiRk1vxY+SiTw/fdALMW
yl89WMNZs38ZCylo4krnUUXg8NoVofv5jJbJrrfbRCc5GJxU6VYVLvbrtm+GBeXYS4iddpqOMXE0
5n8TL7B9fqvjt3SAGNPLG8yH4NJ2jCabkch8lGd2eLyeIZrhSQKl5QCs8zXqfAG8w7rGEnH/EJe/
4WaTKo1Zel4msxm+ihECOFtdfZhGKhc3YSjAMwCiOKwvf7cUYlj+NmR+iCtJgDVzpKwPzmIGq2DO
ymVgD0vHVEr/Jt9xC14BesJa3IN2qqLV0GtRyxlWc+Z2HHPfv69a263EQ86O7FmdoEkLoPYASF9H
qLzNYo6+EyEL/Egrtv9Jpu0Ofqr/CtleuQLTqZMFDKAcucQqKwBJ3kRiSMM8iZqd2OKZObIefzLt
hzuxmLXPnCV/YPKAZTsKtIZjL6jQ5XV/pelaigl7jXjluPDYR2qIz2am0mSWikiPFnuLDuXyxIQ4
MAGzdY4ivdCX5xpHdDIbnyPr6RXMXHsvZOxizA7PrDgck/FdfhLT6skUbvyWAyKEV7Toh3ZkOHm1
a2yzNxFjtfCL6Vli0KzkGME/mgM8zfgM2++h5xOsO3wA86KjScmWaRzGNbAUO9or4/jhgakc3eky
eFVC/0mEYMMwjGd3Ul3UWNxVODTPyfyEkpalDEMVWfNI6wxboPfBt8jc49jJl8fBAvC/SS5rQ4cH
vOC8os+K74aEXPoHZaoYCfNwV+cljsAlaOyZupkt0OD2E0QkdWb+rRBCO3hSQmjdeK9I80vOJBwk
U4VC7at2S1Ywl54GW4DWe+dmOIziS+/WRJx+s/GrYDVPb3I9vbg31Vph5FgJo3exwNUqStVGA+3w
/zBg0D882oWwjz6qrSucOyHKnocJfDWOq56Rlk0uJJoFEf2F99xshm5EcFNHcsXYxa60ARZcUQjo
EZG5lrvUY75ky98HLN1wUBRzEOScxsGHGRfp1TbpXHSzTgL9NbiNXmygAg/31PaCECvIsL4NOpcI
6nWj7RKK6WcQH1iji2KdGi+BhIFdteW7ip5eLy/ay9wLiZY098GqvwLA5LcJWdL7k91LkrOjrvmk
1jh7q+fhXVOB2qxxOZxTICo/oweneoHunLkHcSXN9psO4/ST8a4fBEB9iFXv/3QIvVFZIx/Io5rh
dVYJeR93PnwcVXOOWPTLijem6C5vkQmCibOhI3Urglllv54sALcQLkoA8uHDHNlEb8bMXSs1rqpT
N6KIDtrlPre1z+fUViTaI2Xj91Tnz0L1zWrYEE7tvhSbzUbPJmWgh5BBP1auQPzglFrj7V5heT5z
9uXmEVqpZOGNWpkxU2SGluq9A0BkXu42Wx+YjEFBFXU68/hob0kf+ITkGsAbPRxVo5UFFPBLu9w/
k0FOc8ysq0tsByZwYR6LQ9+Ak+gdfL3W0gE0HGot8RhPyI7V0SRwDoFsryLt0ZwYQ8q2PipukeSL
CKI68XW6gM/auCwXOTaLIWlCRz4NV3VteuhT1yXZLYIyLoUZHbKr79f/lpI0ixpfNPPbOzexGlS/
g2x0kFQLJKEG3KAaxjMCga0+KxPYR7RTn1jCKDoSt+RuSVsYDMcWzo8hMJK2yVRIJS1GPBnddIEe
oIW8w+QmKUzkem7ayF6b2UqQdfxY1vp/fZocFq8R2zqkw2mlMSYeR8JmUhmgCsCMTfet2zdw/ayO
KUSGYmCbP6n+RUWs/nV2zoO61SoE84lkYIFjGHIGpsDRDpomj0TXQhuYls5/kTsKGAfnOu/qs0Eq
lshSjWmxJZlK5PSnIPru8EIphXQmZ4lbUtMmKsU52+WuSvJ3EB3fWh5Td6vV4MdcmJXrwQ1MV2PF
2sqWIR3BvVbP/NhHB0mfllS+nX4kvHsoCQHiRA/WUQbBSquvVIBcGxg7jt8D+IDx/jbRwgEZ40m2
Z88fSJvwKr+w7N4/tXMY2VwMWflxaUv9cgF66FwdM0/dW+nAlvNY2FvTFgcZBfzU7E49+uCflSEH
0Ip0IaR+Ub4bdZUFbzTZQ9DMJTs24Mx4qHmPtV2jbQdGTVIvqd7ZIbizCV5SxJtZObh2beH1KMhd
8n/im6rPVGp5OVkHF0eTah8vTVc8Id5gYBdIS1JS63UDFzmGQEI+yETm0cSLLJwc7QGhUnUo0h7n
g3ZUG/Qi9wh7caNWW5ZQe6YhDzeyj228dJdZpnTnCcP4lzZV2H3/SVKC79+LFx6o+IV21ne7rE3q
F8V3nn0ScmIbhtW4HbegKat/hhSluCxRs4k264TEbOFkgR/ZAXwDfdmbkdg+v48YOjz16p3dsyU/
fVQ1mpUHJqqlbVcc9OjMi5YoNzca1Wumc58SNTxGM98rAr/aCxeLGm7cYO1nAUDbhEWZes5/z5y3
JVJV1BSwc7qcrO3/Hgp7jMl51JkK/MK8XQNhdtB3Kj3+O3v+KEvCQRjA6p/6iMGQ1z+aiJeItIPe
ITHVoVLI0+qP0chnIevjvDtUPEfSdcAyb/uGheUqgGvPjQ8dCsZKkLTldTV3BC9jNMMMm1NVoSE4
T+zbrYzZCcF6+cQN2ZORzdPofReLQ8mOzqdap8HzCFNu8N1FqHAn51DS/eiO2UFj2bbT/qOddEPW
traSTffah1+3R3uFhiMGL7o84aKKKfOtOIyW7hRbwpQD9G9d2NLMdE094QQEHQ9SlDrDYuCyB8SJ
l4hX88fzvvkFG4mYzamb562fvqDdybNVpjtUEbtUhSyyA+URhOiQ5k5MKUoJPiBs6h/mV2vUre84
SzuxP70oEqV+x5iHqjJCEMXzeaWpu8c20ljHMfQX9/5UBbYVJZnXpRLCQJvmRERwdXjeto6g4a7A
zRkutXMYad7xvB1zERljUpJLNHiK7EfhI7BPNmh9eOdYldv3iLWr/5TGg998H7v/HpiRM7/yJiQI
yXM2rP/qF427dpJBbIKiJLJAubl1C14VQAEUbZ2pes6mIP7gRxy/XJJ9Qqe09vR6GTCCVtRySVEL
YPK54rOi9OYXgjVbhD5G6gurjQjd75HJlleRtVUytLZnrv51KLy7l0ZL9cRmbPCvR/4gpQVb9Pyt
oniOkyA8HjkXJu3BpRo4IGvTnd562cG+lGJpqXV2I6URt7Lk1IqXWHMMCCKOfLk2Rbvdc3aXtCpW
kpDKBGu0TTCZRywn3E3ajkRpv72UBHQXfNeiaciwLdwfYkK8wH6HY+tW7EdtDSsqknvQu97lEDud
y7u0KsRFw/oQNWPz6K8DMgkhr88YT1AjDHlDe2IcrIN2Ed9rmh8TmJvNxPSoDoMP65LEv8ZYWgia
5fIc4rZKdFNWZ0dwyNFliIbTqGoEiuDIX1b2XXDGiM2FcZQVRECwJxU/Ql8yyoRo03Sp9D5CI+Zl
aKI2WVy897djqSYF9ly2LawgTuBKufS/ZcpTqqevzdg/s95Y9Ja+EFvKbsA1k2G1HzUv9zWhYFcQ
H9G07HF1mXsgW4fFiM7J7j3elqa3apcBbIL0RddjsCsEa3e+HzfS6ZEUbPyi+fvGSAbwfZR/6n3J
D6Rep/cwdegTC5LqBxfarwIYlpDrdwzdlpAFtKGUUmiQ1bcw9yXmjr0dMZWn/1ra/tT1pTW9W41C
qgf0JdOqjLj8d5ewt77IUb4YL4NhBJJtTdNZQek5T+rGpwofvsXe6Q7kn1BiHH0p3mCULWlEWAP9
p++9D79WHIzTZlA6k26MAWsx8myGhQhuFh+py1ZoXYarY1u4JZrYBIPXy6b52ENO+xyH2fiMkG5l
v587k9QnBRGFDjEY7YTJ6bvVlI+0DWOHcCaaTYCa2SoFLzrTp4SS6B5MK6cWyM26TWQZtwTQRjIM
DUP0sjdxjYU8woxzxrjpoEznUjgBFDakoRRHQfY8ayY4Rbt2lNQgqKPGnTcJeDNInRt52t41YI/v
vQXkeGz6IKyaJI6tXLQWcxdxPgrWZ5SWi7lXbGZsQnVXz5srAfNvA4k68tBb0RcIk9QxWmO8btW6
e/Ay3KL3c+ymOkkmrXy/83SsHTcyYALDUev8Tfl2DTn8wrOq9upPXtOPEM0Dm2/E130FUl4nOBuG
Ul7lDJw0OE7oGJ9z7i2n7ghhCn2r/JRPgz1ui/WREwTGzCiip9SqB43MIq6l68b4x0gzY/GNqn5d
GNaWQVQe8cbkCjvvDqyk2il2mB5vJJNXX9puQ6GXQ/gUWuxvGsxLZcuLxD6jix9meycsAbf9w1AW
7KHwYemA1ZHWSuW7NAXSn/x0VRb7gfsF0YMod/lc/xVUB5ojWBxSU04IK7fLo4a5UMD+vhYLQvyI
epsfkmgGIkkBekaR+w/wopZTWHVhWRTqbj3+/3P53p/wz6xsxAyLTsVZMaJV1TMCeQaxgyxp9iPs
KyNvklyHMxLhF1vhKS4iG/TxvT45wPtzY93OyNyXmFpOld/g2dm5oDO4UG+tLFOc/T2mO4iofcWG
291bdLsQFNIAuMQLiDuMJYjK9DY8izFH7ZNocL0JCPHxhpYeAfY83r56XkkLlBBPkNhT2Mb5WoB9
le7c0O23imHDazbHJ+/l8GS5wWchJqmAM/y9/Xxl+JBd/qHujXrixf4WyvSsmPxWezK/sMfOCKCr
uu2+XHLOuvM+GtE2OhwU2tSY5Wu9iWthwD+Hi5fqgAPoNEMcJHH7iUsUKMmw5eIo26mMCVd7hPq1
lbvOzKsD/RI7P+kp6dzX42/Wrt6rwRx1mhgwHDYA2LaSS/UMIxZGgXbJgxDC9kjFQWdRd8uPNxJU
AljCQkhaUHXYZV1KsU61zE6Wglf8D25ZowvAnOuYL7SfqndNpbqvoqp6nAirfLNl98jzBTVC2l7C
6PwH4+RTXoBqIR8LoLY0UyjkoF3RhlIW4604NKiNEgd+rTU3asdA9QItMQyL7cba4cnzKN+Nmln2
KG6I3Wfj4jhIgTFJOR/hPBERYTMO+Hp2EL2dkSq+/OeWlC34oA+KlwfNbar8jqV+lb9yQdlA9449
BceDYAvIo6CM353KBidftTPFBeramkXzdRLtoP1v1rz1tm7CaL9ACmR1svj94x1Y9tbDNnBWK/Yv
4vzSio3kh50GSfqSmYYudJewrd7mdJdbdvWHeyWcdKW2EHcQJTlkdq4gWKktZDNcl38+s308giLy
8MjIghMN1l0bCQ+C8OKIV1s0LQvxBS2FNtY2T7+r0QE/shMzYWcstO/3S4UtqJkJA0ZpdcehKATm
5OzmbEXbDYalYayXR/K2C6O3x1EvvTicRCm7MZ3pj2Plc2r+ScG683qgZBYmfexWkwop6W2Y2bPg
rO1YGWqAMk51VekbNlhvEI1hMRuM8CSO3aDXX9dL3ddzn8ZVjbUhGPzs/BzOt2r50mllOzADZ80Z
v+86CVOZMdZ8Mt+g/goAp6/y27uz0+rIiGxTbgKCzz0QsK13QGgtW00dmw4m2SFxiJ93OcyKX0Ez
FC7oyfnr9DDmcLR05yt6/mEgzYT3uRL1PJC7Gn7xG4cg7QiKfiNBS9lHazD/JKUF0lXNTLXwss00
5d1+v+Pxw+8l2HPkUEv1u3t2wm0bmUnOyp/lA6p2fFYTtTBa+kv+KBqzCv8VwRrfd5sBhGMxZFV8
0aS4LjOpLk7up3DwjNSUtPwIFLLfLyPgegXPtmo6fV+xgXyBhKdiNdyYo+a5/7vahrFHww0DNfU2
mzLXWS2Js3yChT+RseRQXGVSohggojOaWTXSwtXd6MzuFVseklY39cyRVNp6J59wJG6FWX18QALq
jmigRwwuRLwsf+dIyL3pkrRdTaePw+WUpxrlBkxQLuSTQJqdg+EnMakiotJq1mU+H9i6hrZoWwNg
NNFwUwq8pQbrDCuN28Yq1TQ2Djd7ptk6FHB3o+XQNMrquA3j+v5WoCaM0HAJc2c+I4KTX2KBTm3u
8+xFvDdUGhJsPFHpIyo/G74Tgvj99OaTY5rqNc9ZRnhQOvG2RyouduFHDXBPL4OUtbiK+cAi8vUO
9jEc+CP1bpFLCS0Og1EGhjaWbJ0u6v04p7uUIBvH5VuC9pk4Ti5yrE+WS7IAxEuapzKW4HabKD3d
HdmX4W72VGaclsZGHOM6fmH7AJRePTHyrYgZL+rns8S1OOEamc1vyRjze5Quhog5IIzXUegL4afo
tWg5NGoe32fjCwRyX365ooW7kjw/v15eQdaUvdiXuK7tGSls3ir8J7q3SOP7GmH0ThQXXa4N8RO7
MvVJRFc8DA18ya9CsoOfGlod3lulMO4YeWBmMfwXW2NwXxJTCK0i3Q4RoSQTBDC/w0QnFhoZO5le
ROw8jMcEwgDp8WUT23/g30Rhz6/sbusgiyICr0W0atEcww7eo8pr/Sz91elYGcYkuSNn3iqoRBci
dyytpIHOaU9ToKb6lKdpy92wRXhxDoGU3Qye8gFuPxX/ywG5wZm9T0b3OZZVIp8k0wim6yt8/de7
CM18Jm233x9M2RTOY29gso9T7eDxyLnvVU2XMES49B229SW62t3rUWjtBuTxn2RT+hf4L7V04Ttn
M0Iqjh0ZP74ggvs27vV209odHEhfhjB0jrmE0njyVdCCfzfkxlsWaJrtNYSREe6VkF1rwnMB9Klj
Z8VZIbYMd8Hn87CbafPMlN/JHZIvlC6JqeABEveJHm59uLtg3UVa2FBoryV6cyOZbxfhtce8Ng/n
lV5ipKF1twfQ79dI14aGFjVha2nIyzvUvd1ijdl7GFxNkoZDBQ0QXAssT6Om9Y874qPhdwIUDlHe
kQErEOP4sIhtdXW7qPEaAnqcFlf98XuynQhZ7kP5hZqBk2A1lKuj0fJjFNyv5gj1ajESM3dVOB3N
hcemzI79A6qO0C29OUSGjoKSfKKevL4xcy5d4nKS5lymJXGicjFT43Xf1NOwvn2YYsCBnOYMFUZ0
b/6EF6+hmHEfiHuof4n1tIMDKGDUQrL3/9Td9qvK8p5i060jZa81mzIijUdoqnHEVQD7s+BOXDiN
ZXkOlD2d6rHzs6IrLhpqIdi7WMIeIt2nfn5J/cnX9AUhjgwN0kS0s8Waubm6DtSTGjgXpyEkbljZ
hPF7P6Ylj7p7FIkAcQgqgGEigiCVlzHHF8QWy6bVvSmQ775H+Zgf7rB3vTlj4TBD4mrJ9CV+pSUs
EoVD2hweOsB9UnvPWPkiui6TpVhMIb7Q8tg+ZzMa2vi/cFW8foTlyb5FdgH/FMNICHtCAGhPiWUc
c6FSyNywz2POeXGbRwee1Vw2XCg5GiD8fbKQv1QWtPPqUexuGKNiIt35guNJefrrhnrpVDGXS6wO
0SmkgXmx2m76m+rX1IwRxHbZaK1y7EzHKd5991zd9KV4L79Ny/G6bdO/y+lr4E7fI+/MbKUxYKW7
evv3Cq8pCPAjUm+TvOFuO9ZXPd3FYN4HXZSrY3VrBo3wAW8oXEuDIpxu5ZytXjrtig0GeKIvLUYZ
91+WJbpl55RTkWPxJWMm9fUUzxsYtznmcCz0tsCHwOA5GxWroUj8Nd0KDh3oZiCTBccVyAFY4eg9
uWQEe/zkXRYK0ku+IFjG3ey6IpPqALCbpgyzBMAEY48PvS5G7EblnSczSyqsB8YX+ewPO5aaOWGX
cuGZeIyeT8I8pPYgfQhZKO2s/7sc8sv016tCmNuyQQWA9n4ZIBVGmm9w5z/HuJUYCiqAFTpX8lrB
j40AUO/Yr0ScCLrTWxcVbTyICXMVxK7BhBu8fzvwu7uLrPrYE/yJGlKkp6cleDfd0IQtOMffJR/q
ERK4ssmFXYIiaZJipSwArIRVj9nikPOfNrJTHhMqKCFsNbcYUIiRt+dTNAIPi9sXNzJuD6cHA3gu
A748B40X39zqzrTA8wnPCzXvp0eKTOPcjy/LXm+VeMeslgDAEtgYEyPiWHDHBIWhn2FCSwUuHvyK
P2yDKEPd4rvBAe4FWYiHr+7nY6hQM1O70htzucSVupxg0L0RKTz2bfc0Qx335aj2ui0CLiibzQld
nfj8A/pvgfdRH/RRntpGhn/aAenLirtRPq+NyXvDcYVXnEJRzTu/v3M9/TzHp6oWMvrUujtJ6+DL
p/EMxRFkeeitGt+Ka0Hkh8LUXSqIGVM8fwdfbY39rFonIPqTOmba3ON25dL3ifD5WmHTe+nF8vnE
Irp718nABnIQab0JsrjdIMdZTGSybbsTIEZfBgA8oUQjsjlhCcJdNzb18CELmcEafWYBFxYk3k9/
TDFHRW4KBnVXDPfqDHSGHbATLnFjX6464HhA2i43tTST3A0UyfgXG6F2bb0N2AW9FHkpLZcVCxM7
Ga0VDyf+5X0Kq02JWWvhkZ+FfzzOpIwi03xVeUTxaz21W1OcPA/JHmFP8jSndcamQRTXy3MFh6Ip
TLO4h22QOaveP631TN5HfNUpqbIEBr2AwuT4xHR5aNoh2PHiENsbGVARDCImyRnkeBhiSWRVm7aj
/uEQdwsqlPUkpvy5KLLFD8vSbNqiCyZO1dMzDxb7l8lp10FHo+LkIYcTtcFDmEG8C6OEmkKicBCv
TwB7FEYXBiIoVuRd/W8w/Ow5mb6w2tYtX3tHtNjUxUwZnM+hNVOdtCtXvShHhxZSPYdR8c49DYKe
1GJaay+3E+C0brB6QELUeH6TdY47TD4rSNO9//ZJNqjwq0eJ7U0QlbmmsfMQ5oL+XoEPi5f/Qdgc
Up99ZWB37535GQEplAwXpDujlb+lLC2n8vJjyOgGJhr6cyoiugj8AURjbpfnFo/Z3TV5H11pIPs3
pWcxRxUo638XPKjeK1EizvY9jlgeGaWRcRK32xfkUgWKfGm2q3T654cDLatvCBtIZ2T371kPMqQm
bDRCz5nzx1spIvGx1C2TurX02qrbgM9aFyMjpASjFEoZ99N/1jcWROvOH4JZvJDrecAxJtj/Ndvu
4x7ayi4JGx9pJu1sdBjCCMAdOzNkN2OxdrpRjjaLez16blYZzafJ+4uizTaSFLOq8+Q/Wh+Bzp8g
TN5GTyee8e3ptQjXQocEdm1ZdpKSNaSD5zPhvLc9STxBN0vLWFb5Uxbf7zS3Up0aMU8DVFND/92d
Vd32zmtB3g1J+Bq3qtAItzT1qRbt9H1dvJSJHXYSelYvh9sQsY06AAW6svw8bzYjIx5P6LSgwZMP
WBzboFAKqB30KDP0pIazUBQ/FqBajx4U/EquOUyJcfwqBqrghQDndygijtASYouZVcwUsTwN8gO2
4n3YscNoFUdAA3fqnzYJldx4d/V2UzaRzh/GPaxseycHgN/mFBBr3Ww1EjPTm0AC5BkK2UWOKDxR
I/ySNwik+Md0Sz3r6R1eEvTKHt1kdBJG1MDflT1lHUS3Xx8ZmZixSxMJF/MoGY65GpjGSbe2GMdH
kEpMcLtL8cnG4hmOA672qopB73xvHWQhAHonO64RjxdXfqeTB6kDsOvzByBiYNqgZwwLZr3Sr9r/
BNfG1d6dBegVikxXi5xS5EnzRnijRNdwPNAecvdPcFGuf9vc+eL8iQuhyiP5MJZu8aT05JwAovnV
u2SIyoQVGuGFGlnzshes7biFYPqjAp2p7wO4PMfT+i083RiSjd9PwXq7HV/skZfUD5fqe3uEH+q9
1FRq8xJS8pGC355yDrVGuO4NHZNXPsO37QmSwyL6ba55nsxzEYYN/e3+tanyIQQmA5LHIb6I5mwr
CFyipeDY536UEIUeENlntqbxD8UdjSgICbXBlqxG7OQkCx+seDevmzIzbgHKaA/MZ4mhUCj5P82d
U8rAZzoANtnKS0ufvXFNeDIxRchC18Bmx1lyz6ItQZkeSdW77AdozpS5QA8gl8ahKoKZT2K5Uvhs
9yjrsaGhVfkQNgOJvCye+6vgc+Pps+2kkUvLWC3i2E8v1NohfqXLSSdr2aRzq1SySxi7ZAtqEkk9
P/4e2PtCLgPnmyzmQbZNHBOeTVGhckAgETsCPcdWfeCZt3Zu2f4Xgq2Zo0sfUIVlfdLlb6mRGUD6
EL5vJZ3iAlQv3PjVUU6xya8Myt293iY5EPoN1oGi9mvrgiLcR9LeqPkogKJzxPQNPI00mPZ1dOiJ
8+fuuF7pdJxeB6DJUO18pRknQQtCL/fX1V3c55uUPdtGfBh6IYc7ehesZD5TH5ywML4vRo+DmgTM
YC0T4f+rLUFtt02Z3O1VFSpQbKyLH2Wp5y7DCKlnOyuQ1asTBwJziYjCMhWlzbCB/3fyfnDY11B/
/sE6E+YhhWgLvQoOK9yhFGkEW646JN3rn/n39vyHiqj/oCXRG/hWlE5RfgB0s6+d9QaSq0jzYSUw
KGQNsCbfPkCEVUMSoIMMZo2ISM4R3PEEha85OqwQR0hLgiItdqdUM3GfTkeIfijKjyXgVC63/jgU
/5TW/dNi6xc+r2O0S+4tN3KcVLKGcoeg2dSiE6FU5MjKNjf4VlSKYNfTIIcoc+t/49D72A4pxibA
moz85FIUPaEgUrN+uCOku+uFYgvPSvtbi827mE5visWhktbuGFyMhWcv12GDcHGTl0IaKupSeeoe
h6XH7QYmNjow8OzBYrzCi3VhzrScGCqVXDmbP48SLUwuTIm9qJSAyGEMiwPmG0lu1zkife4Ipk8M
ERwW7vM8ssuQsRNmoAtHbA6fpY4Sxtvc3FuMeeZyHo0pmMcL9ESBcVtiFyrvxR0OBijlmJMVI5hb
n/nOXHbEB0s/68hWSTOdUUWtoQj47NewlUJUE91KUQebICUvEX6VVBnDFbdPt0IWo3CWjxS2Q5Nv
sHNn6ElcX8tS4MtkMpJpuSw6FAEIwSz+zwnx/tt5XSXjXedKSb5/pkVoJPIVWmSI2BjPfzGyD9MX
0+vySErUY96c8laxU4EJb6bzFYdtb+sQz0kAX0sjOlXdizTaiUr+MFuNaQ7v78qapStvVhxWrc3f
gy0Q2+xNIG98VsT8uK424EgqGpRaC86LpAeYPBwmUlQHMrmVZcKiSLSM8yOnNc1dNraPQtZKcbH8
U0lgLw8RM6K0Hdi7mCv9NPkCLXsC040bjEWVO3tSw/XYh3ZuK2qzEUCV74MZPZ9rdbzEZeQnR3ba
wSpb1DcRDVix8AbAcdoShaCbn6O+i0MY3YQ1u7KMMBAKA713FWHzadEc/Os+qs6J/oJpv0tjv7uT
ND171ET5D4jt703Vzv2UAkgoPVn7/2tZRoC3t7aUGJ0usv0JYE6HrSiFfy6+jynvsw5jy4gFRVeY
cDBKCbuzUXtrNP8wd70EARKczXZRrVDKCmDhhMkYzBLJAL70foiSRKikiRnP0LFSLS/UmpfG3Piw
eCOhpznhuXfedNxRSRFsp5Zmv37+z8wX0xS6EVaklXGUAdpHLiwM2bG/HLCbdQiybpqSSjoAOKIk
7XXDrxZpzZvu4sqCno2/E67Kan/YYOutuja9bF0J0hXjwy2c8oIKqrJlKQ0lMc8stjYQwEJubF4/
iV19fp7rZ/FcqxO+4omwLdUY/N9Dm7w2GQP+I6w72c0jDLuaEPuUuMB1I6EDSwWAYGiTmIKApDei
QHk1hNtAtE5dUEdrqZ3pBRayGFTIyUOs1yVlrp/tAC2ia+iJt4U4DWcytLkzKZ0y0f/rBYlnr+0B
HwKLS8r4NDIkiDMlHZ93Og5uu9NNlBBpqfmchPFrH0HjUqtRuKMTUphDmZfqsSwiHxi+wkNiPnbo
4pc9nHf3ep1JYUqA6NMX5E/Rczo4T7Q0/Y0lVu0DqfEpHypbcWivs206QEFJr/TRxWcAXQ+Pqp2n
w0x9qfp5gZsKABsz2aVcpaDKUwb9PArq/AWUYPAP3b7uS0FVVA33qZC8XwYshwzduHsi2Lhxi/kX
ZggJth8a4vRf3vdK/dZ0zP4hDwByjtWEjg1k34dhWwIgoQj+WNDN27ahVGMPlyYNz/nnpQiVuTZ5
GLCChPFEQhAmTEYgmtncZPrbuCLhUuM0Uqa0txibtbhdT+B5Y3aUmsqljpgqHutNaKHd+1001iDd
XlBbXBJK94pzFNnszSGsx6yledffwbgdwbxMLxVIXQ7oEYru8MFpBhAYN1Kmue0z67hAoGn23EE3
bhSnd1OqXSAbPrerrh9t5r6xBew1SVq/AHUjAviQI/94ScnXXiUVI3i7nUBFmFlAtDyFAdzDkiD9
Hso1gCxfk+cbA+EgPzWd41HEEPvcvCONES9aj/v4dEIofZdjDz+oXgGuDiUS/LDRAjEgdvPSQ9rt
96Z5EqZ6gAQKFO++rEJJpfuF4BvRCnx92tgwmJ+uanMnauj+kv6qBzQwq8Ijbd95irplPN0Z8tI9
UnrHAu/3RSsufUoT8uWOLQIchrMwIhn8jJ8nTzCBhm1zhV9ZfyUsG8nEih3AZfE7WFUhUtwWdtjT
aKMz3BlC1uHX44L/0tGV/O4FNZL5K3lHWR+jKtKdJ1Y6AI51ncmO2/XZ/WkmkK9dIrdHPQf2oQLs
V/gLNzQU95nZr8Ze4qGexJndAbEN3/QX2yVd6WkD9eMtaoROlBdE+cscDCQPATrD54QYK3jeoA0A
rwcXlzyYnHXGxNN30AVmx+So5eucUW9HbBa1F6iZiT+Dse7gHCfpOoSME0YgH2GOSAJ1uvqnLeqD
ceK+18xv8J+vTa+hjhslUDSyRwDwZIN5+GbmHRkCDkRZ21Ycaml+ckS1uIabGJOClXNr04OBdwW1
eFS3Knqw4bqrWSte3BLp5h45ligNY9awyRmSXP9zQQG0/fzihuKlrQwTTSsT2ordkQCg7H11gikh
5Al2VZ7LBnt+n9L94FOf6Lv/rMcQK2+1KxKa5yJdULKyifsEdbX2Q9wt374xlDZVm0ppSjDZyh1j
Q8Kb+RaJgaI6JLP1/sk+Im+jgkDLdOw689TJ/YKxXm0QF/MizROflgXXimLd/4DobXb1whg+2K7j
bBoE4Q7HUN0hDD28V2W5RV80UFGVzoAAyzx/jSQYTLGGZoAID3rRfepVZgQc3X6zo3oqQg+uVeoS
u6V2p9LUy2RNSSJIBnLMCGAJdADfnVOrKcDBmxcCZwT1aUBFQ196I58Es4v6RG0+peFberDZvIJA
fOkEONiyfcptycP94esyH4zdyK0UntLzKZRC8m5U0ItB5A7qA7gl+NjsQKdJ6P36QF75aZUv8bQu
kgCWBddG5s4SJdu6ACPMaEzJ62lgWaJ3P3kThY+UxFRwD1T69VTrA68x+cgkXPo2U/9KPRDVPfQn
plfxqg1O8/8JLkWN/4eY54XHHdec6JhQu1gTObbL/7yd4Ny1ECX7Hw2MP2y2bVrNij1Mmi2kUymy
GgjW3yJBDGcsPaOzzi0KDM/aDc3NaB0y9RQL4X93Q+2nDbDYSLSvdUeD0IfNHsLa/TYSPFnAoXsR
6raDznd/QbK0xuDHKBZkm3z80uFdoAORqkgWVwtQd19GpnYqdc57mJ6EYg6PcvOPq6YamgNp7v+1
t2Hl0YjPH6gClbvIQvFHMCjgUH+AZoBm/ERdPTaY4E+ubfJKMf9MD+/Guu8ya12d1lXl31TtGdxJ
SvE4NVTWzmwT3Ks7zvAcHtcp+bluYIJiCTHMw1akCttrnnM/vTKRojSB9bsR+NVMdXdPLJ7yWXuB
wpk3/TprfAAUfQGHMOK1qOXck5AItnXpMISvXcAriQFWtC6SmWo8ev6Jx4dJpcI3AU7Pb4E4FGM4
RtE8EDVQqIX5gBhzQlLzWvHyqmURfKXA1eZCWnLRDVYYzZ4EWTZQJAS1BZ+70piNwFO056QZpM4I
o2zk2Kr6uViFrYZ1a446sUq0lpgAboZY4JhnrTYRYflRfBQ74UAFba44f7FMyweWOEIcPL0LKLbh
FkpDuZ6VwDYmwXpVH6J9KOYRcIPHcAHAUZ3v7oH10MCdRa1CsknZKlP3HegdtKiqV+6o+fBt1Ybr
HYxvdl0+mgSHLvD7Eb5vBhBA6wR9nSms0ssEweHymBPc96c0hJynd340eicgjzcru5okPKYjT26S
e6Ira04N3lnajasf4razETfE2oEa8ZD2END5K5xKWHAOZqBkHTINERHvGlkqqB7C3iZWLKYQg2Am
LC/UrhFyreVPKDfjK9NaIZGdyzF83MbY2uMUx9187GIHl+Xm40RCgczuANiC82VMj1EZ/fcPGRWh
ufHUm+qIZjXkZVL8wqtZCVQgFZWA+jV7y61Wj20JTejpgJP5kuahAH7vvhircVfVGIPkk/MDJtT4
Pri69+O2OYsr3JII4dx9VoGWvOT0RW1PyC0dyZW0NfDjPB9fTqIcYueKz3MLuCp8EuBydjOnCNyE
GINn4dUuXa43KLLi4d40gIKcrA//YdWTDbHdqPblfzWrYH55ElvIv6IZY0KE+BTCVxuvSFjSKxNJ
t1hs5Aoxur/YqarXOyAdVsHXMGboJ+BL0KosTKkbWP71MCfz6cOroGFis+OTd9PQFQdSHr+VkG74
5v4MiwAda5+Ck62JR6u+TXM0xt+UO3kmv3ZH28gkqSQ4u4bwz60bR3Hw55hGujzrkeK0kFI8DJOc
08ZVKyu3glKXgrTV2t8w90rpYQcbENQb+aA5uYd0vcbUJJHeeuW+GMeeSmKEIoiP4VIk/DMH3kfb
Lcc+OuCjT5/8PKFChjj2ubcIeKbsrJMx4Ins1oFg3HTlRrTWPzAz1jsTm8/uY84Le7l40ginBNt3
VmTCM/Xy68+zSNEgAVS9Gr5lhYO3ELeHe2AYDY+TWZT2XLrwdqXPJFRrW09KHxrx1LgkY/zdZSQZ
BTAEEJ3nzYRKU4jKl8InPhl6h0kaeY8z09dIAYZuvQEwIsg1ENsyPcjBVXAOVeJiDUGmiJgph0AO
sI+XFVvGhv/bEb2iSq46BATWvO9WGcOmC4kZvM90m/xTE8ii3kzVgSTHaEm1POwxqlcM54GVXe+p
ECqj3kzcu75WGGyZ0VcuDbhn6f5eCn9pmv68SEXsAvdBzzWwz4SOQDf9Fiq8P9udD6S7Xnx2n6fy
9tLTylfG/w6B51eqLcPHvnbcasK9B/dY1v73uzQ/04ulW/EVP7pmBMSnXEaKhY8k1jdlfrVmU5dd
XNy5WgYgNjRVZ3XUMh4sP3tfqar8D4jrmSDhkI3m6Hv4a8a7f6zxmdXpTNk0HTBdAyGXYEdJ2EH8
nG5UxCi5qzHIjhIb6WzUs7DQ8olNJaS02/lgUwgzxyDsL+Ygw2Aclcd/YKCFMvS028xr9KN/wF9G
vzkW1dOkYMHM5Z9/C2Ecw7dX2j/DA/k0dOLnhK9solmfhKZT2DQA+gI3eobkjhUr/U0w9JI0R+3E
NgJJXgsvf+tipldRf7F0sczh5hgx+qoXcRFDlQOW7n+5ZkxKmnQqcpmCpii3hJwCnZ/6dnTFHNM0
wNaZHMlTxt1zRidvAVAcmLD8TdxBuQHfLVJRD0E2LqT+Nhqkjy42ywv5PeF7MNtygv8lvvH2peRU
A0dH9U8xfSw0B6K0BbhO3PQ0JAnqzOGnmv7sL6idlwXtTK/Lbt9X960yV89oAKJ8BHR2ZGTUGLl/
3XpYZXW9OO3YUCvALql70fOXos2IWPm0WzwmRbanZ/BVGTlF9O49soufeVSRw0rGxYlTjFl6l/oX
XC1n1dt3KKQFDN/Ycs3OhmG/pRP3UAYjlO+sc+0/cH7MGwwHLCuSqm3eEwrZBWW7LB7zzu9re5mL
J07f5r+FI6FozJyz5/O2JbzghDhCe7/dSj2cyRPm0Ep5wVoG1oXjd5Hzi5aVUheE54idt3QiMNHu
+M8RR1ZvxAdN6UT22w1thNzcT7G0OicE8gtvfWt2jGpYqOwU/GSeK+jCfFp3oAUZc2STc/YqI8Uy
CCcwUFsid0yT7atxHytA/0fQv0CUkTkfZe3PbTXHOcMZ06uMBxFI2oVX7InqX+V9qr+9r6vpomu+
/z52JNphJBTTWC8/PN8jA3wWXktjvzUJKOjFaBVEoh6ABcvWfteMZRGE/k+Cz1MxkWGK98Rdw24E
c6D8i+G5giuaDgfCfEBb/CwMUt2fU5evJQcFxL/2t6IyqnaO1yRUeqD80HqJ/qqFe78T9CLOdO8r
YO9e9wQKrmTCjhqMaxL4jjxu+DuV6gK2GY2AhBhOVk2s3cf/RYD0rxnksqE53uvSOY9hIvogfniL
I+BtBujGjRhkzvDTI85Z7QPhnAkaCo5FFFIoYA6GBtbbuJLCFoOn5hCrp9ILnearI+IDq5HP1af2
zR9rfiZ8IL07+lu2ckCT4oQjWaQdPXBs/FhDEdi2ESmZSchG/sJVq0nsud/e9EPIQU8lvjmjMI6r
RcKbm+LhFdrb9tRfOwu9byqdBqyW1I9MusCMaxvEC0s9gvCTgya7yCRElyj63kRrARhqTquD9N0l
ADsTjUXOXvYtSPkb3pZInRcBP07Oavn1PiQLPVYjOWvOZqUujgDtUBA+5OSKUgRimKMxgb+lKv9S
SgOVplSddaqAV1aVHXY0Au5cEM1cNqcAi81cjB8M5v6UFTFsVG0cJmrVV0lPxYP/dcrXkca2iMXy
dq5tzVFDLEb7p6KcWyDEpyb5WunIx/t1h6VV71lXeJh3KsxtUrLEh/6gFYfuaFpYvfrKSPlBcVej
UlS1ZGbX4J88i8+aMVrNiNaDQm65vcQ7efRwlsBXj+ThBMb5kTXqThB9t4j7VK1SUKh/ZAlnqFhQ
n0521yQaE3LIOuI7bKaoR0aq6gIen7hDROt/+nT9QFeTM3xWuQJM/N8I22cumeossSONd4iVlQKM
LnDSt9TDfDhkBgx2yxJvBW75M/QNgRpeXn5UXW9nxeBgIq/lN30Ti3CasA9nfknZy6QNTQcFhFpl
a2Nv4cNODcLkw8/fPEiETn+QhIKjoKkmzo+VMlGW8sMJD0XWI60IjeXCZsZmNmf/6LMZukr9pdQV
57Chh05P4oI4O5l6nziJy1/AbO6WLyPyn8SUdNXC492KWHiWgeDP9sxNAvpnwI3lBovcOaMGAd0R
EJyuNUuj8csDjCTp1X/IDGENrvBSslHo4U09oa1QULY548t8Qb744AsfhfPPtpvhRsnjQ3Rato1D
2348PJrqopWjdEP47i4IIZbt9gO4AVUOUBOhYNCd2288ImiqLOg1mDlPiQjBM9jsTOKXl5GqEc+s
1/ZHKnwgZyxJwsfiCa79onzBbjTq4IEDs8e+DdXMkQsJJStguWiHsvhFuUgDe2cVRx62c2yadVxh
iIKtMR5P99x/PFuaTs3htJD70sEtfmmZFi0FvsbMZpDjlaN/yAlPcD49hrpIBE5kna8tznQS2z8M
wCsZqKZrRJMTh4XeafeAVmjbJbnvO5YQYVgVSZZTU6xPKbUTXvBg+YU6oCUSA0Spccz59HykGaQN
5DNy3CbECTcAJZUQCqZGq47uh2AdMSHIB4hm+oKsJ3w6bdLj1qSs1i/Q+mmh0Oi/3/b+2PuOaVEw
/DsCJwCJwofUlkDNLTjoiINCl4OGy4xaF3WQnnNHL9HVqgBszrkffmmQtf6xUnN+JSHLdbOMzo0Q
1QqWeZa7CaKqlxyzqcxEUaJPP6e/SKRH5itDHSyC0EwKW1HyEGpo8mBBpnVqThfKjk2J0BlqByc1
63wsaYEiCF6OoRH1w0jRpN6wKuY4+cU+0Ul9TdSDDPGoVz1VNcZdZNeLjqyNwXUV+ZDnq3uSqtEe
zUdTYyyTertOmVJgSaOEVXZnchswNIdBuuFWJiWvghl0ohHlN3Z4zsn/PaoV69ObhWOsKTDbghWT
KQt8MQu8y4Bz4wsl0If87fcoTbCPlUSTPdqV5zI6pQWIVPmIj5u1rR8RDukjPMONlW2bV0Mg6Gmf
jZ7/ih5f9BzGup6ge3sRCEA3KWToEINHlMAhrBDSiYepk48/beXuF+P+1yau0SEwrwXrfThqFZQH
g2I0qPzKfjmFn7BeWsXsfWW8W4kWiF4KejzrUWjZCDZv9EULbGPyA8HzCWUw0BLEOrrRtevThwQo
i88Cx/wxsVTy43eqbaxct21WjYZgpOBBL20GDX92VqWtc9AllX2ckpKBHOru6SraXig1JGlht+YY
ZO0YNWzmWmxGyJv3CFEwgrzw9RLkznlN0MAq/jh/DzpL/JA1MUNEdeNLjNrj7bBwI+HTUD4yZk1N
OeqAkBTBWCDyFrINVdH1dRLMgL9BxSTTTrQ5zrdBJG+MNK9IpL2htbUbTOCF6LbyDamVoWTTUubz
sRMyMhDRUWNtZZwQlOxn/eBz03AHD83ZH9veCImMaDcketo5NFRzL0GL2U6+UBrKxZdyJ2DRyGNL
2J9ysejp+kFFsw1o1aQ7qZ/gAxtMWXIXPPcT4XQcyo5/QuSViuGx0p1pf3ljhSREH5xG2FiP9Kbw
IyCgZ1GVnf+GOVl3QSoTvPFK+1vOQ1J5YWvTRfhv0mzkuNe9tM/7D0lnL1E0LxniWltjjyGJCJX/
Utv1nxUz9k2Q1rqEA81Ju+pa2q/ikO1wMTSv1TwaWSDvD1cwin6OTlFPDKjxJrz8XI3LDko07zL9
X0vAP0g02pWSNX4eM4UxmjgViZYa9Udpgh+2Lag85uOVKCu0eyVzkzjo5dm9oNOmBOd7Rg1+oADn
aiOJMJcpVwtpTmKVGpMEUGf/EnYY7jALoBd4/4EEcvY93+wYre4Yutz7eha+Mss1qJm3u110twW8
yvr0QW7uvS19MKmfohFxgbbLZ6DIqZal0lfvI6msRs0m1vS06P8PaWhBSlNm5iL4X/UxOKtyeBhi
ry21CVJHIyQ1wszNuZccHIi+BRQrGzXZUQoeZa5wO95NqCgALkHk5j6jWXjiuigs2KkdVdeSt/Wf
tBJ1eSYNyO+0FSGnutk3lUwtm9MlDtYb8f8zJbDU9Hj+8GbzS17445FNtIqSVjB23Hy+7KMTAlEC
oAO0L2/R3f7yWcm3PYkV2vOdKktoX7KQWehtq1gBPa4zT5wY1rxldWeKBEKHRzW3ANgYRmx1sW48
Tb4ukudYye5KhtxYQwmSkNUYja1u8bUx4X6NrvgmINosqwhkkMRe7LOfPk2sVmIshrAdWG4tT1bV
OnlhdHJUgvNlIES+vZtJ+mPZY59lOxoQiYhUmt/l+jRqnMEQXZB6IaXn3Q4nTPodEzUZjrYovZIH
dU7hX/7VVU4nvG4Lfdm7CGsChoeP9IB5AaD8EehCKag3GSEaIOlG6vb0xK9JAuZuI8fwiS8/HTIq
HlFCh2k0URP2CekXePB9PztIxjxVbcdZVzalMtYh9PN3l7pA+bi7jUeqXBX+U4MeFoSivyMKKWq9
erbfgpUPzskD2cK/dWRQrOV7vqmRJpiIYa3GSkpnSbmmEKGQJB+qPyfLIlDiEp2wV349Qkq/9E8d
NLpHRpLb/22tsaN6PxnFzNfs7BRx5gvIw1QHrFHUpRxje3YTOjaVyrypU2fkaRjdUSDjwsCtNRIp
Pw2eqoyS3YSB3ckAWKPXy9wgMvvMEhOqvqKNXo8t5Sb8bLXAlBcTyePFVA5ZOR27ABZqyCTL3pz7
aVzTsKTh3yud0reu7Qux0UtX4/2UhRQWxlZdLOkWUfHy1oZXRys4kdqokDi8hfhBn9Yu3BWVY5sE
VVJ/Thrul+5u9x/ACujXl2rzRGjZR4PEN052du0lHASRDqjnls9oaVYBoJg+bPJ/9EHtXpfUUsZz
eQLZXzJy2CcFENiZ0nekrAdWqqQTYdoqDzjm8Hh08Lx1ESK7ofoTfcYu9nrPjTUxjimRvb529Dno
f/WbNC49b8+H2SP1EsolVgKkKlQ3J1nomn7D8ZdTPfEXEfBepS0fFl9JH6WGIxmo0y5PsA0ovyY8
cPENrVidOYjogDSP9yC5WAhNv1zMHFxcNonAMkFmUTaOB2Rh/jEHVC4WinAr7ulPrmT6JhUR3iKO
YiSzAqf9G7m3lPWqH5LMkgDqFG5WBzFU1ipI5/qlr8Rft6+OryYBB/TodzaItc/gu2EZvNSDTiDR
o79vpc65Z3wjMR6oSa9tV2GeMD1PJWXC7U1IpFwPaerQiV9KfT+3w1nrH1r5Jsp6AgWUarMvf2Yw
N78Y8A1ct1fWa/M6n1vDGxDCelR5gS0moc0FtbBQaUtUwE+Plv2R8K7Vxek9qDricn+38c/Jd/4O
pHyuQa07BTh+R0jWa/264P8V1MsPZZ4NEmSx6vDj5CCd9QyIf0RgC+4xOgf/JOJA4QBLjMAzoh6Q
dUID253OwHkS+2+U036FlVGOWUgguE3zKiBf0VhOZulAwR85hgt2sYUQfU5alExdCXIN4rQWlPg/
UAp2x8U+yMQcr0eYJAagnr4FCNtMV1ARGk3WT7g7MWAz/i1EOEPfvX7QG/76chxDnggSKoPPjWHw
piDXhH/yu9HCwe2nDxgYaO5zRFyvuxVxEcBkm6J3HjwD20AeGrB6RtLpygzeJSgEB0eLONI/rGB1
Szpvp3CZFAFuSFviqOf3zaonAmNDTBKa30qP3vdjF/SXPqOh1dv8MxDHMyCcmLbdfuFXh+aJMADl
Mm/7mfTeBaSpMtv8phbQ0p5ulf5Tpk4PoyqXBzLAzHsXiA0qIkVtalwbYxNFVbHvs5jxtJBdSOpd
R9DObPhoTNw66d/s/lBuE9DX4Hsq8evQGqra6LXvFEz0bOh+63S37yJU8yu+Xxz3WpBe701ee31K
oLvOwx0jComyPfNNMv/haWoslMyP4a+YjssyajPCGt9jmc0+EMuPaiqdAKhbPxozodi0RAD0nut/
+272E1WtQKQj+RU4nsfaTZbJ5eyB5AbAozUfPxthqHpiYYfDJ1etqiG8ps5Hk1FSUdRIXOSigbcA
jz5JHaPaf9kuSRNoFXG+olWkCfDhNwTv8Q0EotOla+3NA5KxNg0jtHv1R9UutSRV8W1yX+HW+4QY
I8LUJfd7xfiLik6ZCLeOG4TSOKlnnG5JopWQZAdICGGAvQMuVX7BqgbvcOgVudmVEZ72PXYrHAgK
WfdhEjkv4vheqGjO0uhdk/In40vbgVk+kgum6jasdsUA6wif8jfwmImFY/uFL1S+jlLbSyyKMuYq
H2kJwvEvt62sPr3mAYv+vKzIDdo8pQH3muOfLO7EtcK0R/jNKtr4jqT/SQ93AXCBsccXxbnPkcfG
j0yEZCfAFGBiSwQy8yC/ybIwek+QzJTXnC+A6ZmDEM8RTGvQAU2Wcm2ulyWWCSEb7seNS4d2ZJ5W
rN1kQ19qK4dutjMOzV/KX+yEi/fQdcfRz/nCew20FF91OyhpHP6shL3J8nztFyoAngB127Gecq9u
B07qCjVkNI8LUSg3CmF/nNs7HHcyCBc0A3CSQMkMNoIv5bGiI+Pso3WcUJdHLxQ4wjE0oRBLy2zV
uOpY1GG4dbgp6eKDrWXesfQ5Sl/9k7dHciAzWlww+Qs9rAms+z86By9w2p0sVv29h4ViGbTJT6lG
H8n++sSuNwj67osayV/FPVAb4pDLFnBTV0wP1Bar/wCRhZQA16qd4XpEes0zp13skVTKLhs7XpkW
fiSW8MusZjtZWVwF4cvxQjxh2BiNy7biUB/9XmNwpJ9rnu+bg4ui2njoTufydLAA9wgPpinU5rLO
wSxiIUdwP0xJAl6w5MYfmgLCjEAhwjgvVJiH9CDDA76AlODO/XnN+eRNzRjwDqLcpnQf05BD0RsH
qVO0lgjxHvX0y5pUF01Dt2T366z6lIhtUr87qtvzrjnV7MSFaVUhZndLaNO+Eby/esQzHmChT4FC
pFH/quDhytHmduG1RY72jOijZUYbNKd0f3OSzEN0X2cthMQpaLH+pAtoMI8aTQ+qWfBFCRgzjO23
k2kNJ2cc4X4Lq+l+jRFg3fPygySovsVTLieS03kxmRoIys7cRW3XyN9u2ki5CNuTUs5WgRR63L9N
JP76u7+CjUeKQEsbx+b8+S6mD/OQhH8R1QviPHPG5O+NwFoMN/eY5+bikmqC63NZbYTXW4OTvSdi
oEVVThaiQZ/o8NA4HDQTf4Jd9JBXs7Qc46E2hfeR6r5JD8jY7+4sLLCP9xpjPJXS2K4OlvnRIyjl
EmCUEeAh1mHbCihfLm6X3X0oOL8mAEyJg8vyKvM+JJdwwW7ckPmF7EsyMPA7FjosEJTpr6tmcjIw
zrRp5iBmomM2q/Na6OmmlEme0qLJFT6Q729fIayXvJvnns813LJUqrcujm6e/x5t99hyneRnsZjj
5pHdA5X0YD1qHpQVsAOCffVO/ebjN0/FXU/WfixZq8kix+rinJfC98p3nqgcuhGhmStgwCw1knCE
8hVrn+gE/7FYVSLe40PSeZaEV+t2Qlevy+BgidHYY5rVGO2Thr76BNN2qFO9pfjKPf6Plpzv2ZZo
DyN2kkBTSTNl2cURBQmJBnjYXzq9LG5DsGYVVaL1LJO9GUn8WayZ5LV3oHd2kmLJqdjKqnoXU2sn
tBKbf5911gZUAD4Svmar9E6J4wBSEVaEEjvCaEVgTvt4e/G6ZYY/tSHPSic7vKIyghDS1nD61pUc
BgL+ZZzFzq4ydG+/91BITAjn8mVzmK7Ztx1f3BFRIAufQZaUqDuqZYlta1GhV8IwhDeXocFKuLy+
tvdOoe6ZvVBUlLXgGLdPW18tBp2SgUVMZQvdTR6Wgg+B3LtDaNqNLSE/2p0xS1iI26XxVirXVdol
z0ba92tuNHUFVhF+6Lwz1LX3eBP0+mOA748tu6m252ifcc8UHeVptpTqLLnz+3SvE9YU6daGLqeK
kbTKniPmGg2Hc5xi3MlBHXs1kg4ImV77lJ5wk88L/dFm12uZ7o2yuQ1oDkCT0Y7EzOxwngSuauHx
9JO8JbprxhUF+L5BeYiEIcWzFj5AwDVW6BAGMGo8tIjjbpDfVZo8m2VEnQbN3LPADEoHVttC1qQ3
h7Fur/IRbqEeDogRIfUlkZpschvUMDTvXYeuwC70TaE2HfS2itih6aEfz2Ec8nS49DOX5dZAL2gG
autcshWBB9wZR0T8BPWxZYC7tFe8v6yQ1ohvULsqz/ZurNPU5fP7igEmtZ8O0m3g2rEGsHomCnKe
SqF3JRaz/BqSmBh2d3tuDQw3X2e/8o2/oSv4ZpWiaQnm3p6g6CAMHB/0HjIVuK4HjN3rLq+yrkat
DCp7pl/K2Sv1tFCWPPZAYZ5B+xakTFe1QE6JC6k4ZZdwhOonAHmyEz1cuyfd/Q283he9By4b9Y5r
QUnmHm2C4LwG5NwSF8uFgiLYATUTf6+A2+/BRDJISLunDBqBqPEJ3V2x9Zy7+NDk+/jTJflC+0aP
iYUOZOwfgZOtyKdflTnIl/tCgDcNBTDn0XPCqZWv7krxKT9s03L0l0T3KQ9DWN8Bt37vDS1irD0u
mp4jw3MmXYg746ma/IANcnKS8ZJ64jUa6uuemPrwMiNaiTNLSxIl+sxrnF/uvypRaKXuyMY6BvWz
CJS0tHVPZ2Qr5F/Eqn8wUEy+dXuBZrf0SJz+sGkz8yTF58Z7O7TBhgdOlcEuClrjtqGMQQIP3NnN
cCHn8I/23j4KTiwBOljH/bRrnCaB73sxcgQWRUognw64ElMgwU3ZPLjAIYZqWb48CPlVK5jhdGLv
FziJh8PRT2iZ6gDNz6Z7VFmFamM9ZSaEexPS2gyxCwil5Phqo8DP0+jC99FUiFKWkrBvBtX21ojx
hZd0JdjeZvuZzofQERSIXkkhS88JuUJzmf1CbMxQn2dhyeI4D7myyqoiZWWfo8UJbgpNGMsZ8pIm
AKWFlg7s3YXAE66uiN5LIXbks6j21Vn1TNiADUwrgvSOpjSfFYRvwmrZO7Tz+HW9iECp2OAd6ZCz
qJbGdteIgXMsbm6bEnORxwWyx2nNqeur5jwrCav/0/YKFRBVSMcaqrI7jJ/o3/Cfopqyb1sJ0IlK
cXR/ESeuYfPY51DYLa/Dfbzoh0FSBbM+4VMlsGJNvUf6oSNrSi+XUtSQ43dpRJmJWAviyCn0w8fy
L9g/yjyYBKDrvPBo/QBmIH7LHqmTDeds6/FqhEpi/o8XSFV2CGGBSPjioWTV8wa5mUMvSoc49H3A
xOTgNIwqOlT9yaacFH2Fg2qzNoCEPFP5aqiIkrB4FxFbtZAYuYgU9tnxcCEaJPIL99dH+GntpFmV
1aK+x0AFWnOc+yI2Du+NXsnDr8k3hvZuPviBsPNmOqBrtaYpNHRLf2glOc837sj1jLDqeDtCb0rV
JewJoCqePrLYRtmAu+7BJTCw6CfDuX81CdDvSdJolMD+lfy3B1bPSyzfGcV245fJWMIAfW9xdb2X
BmNBpoc1PEGqUa1akO6LYyDbQ3KJehxfIIZVGuqEbPUfU/2Gp4M83hxHDoz8dZdhTNSyKzWcX0gY
bJ0uqEUoEYkxaegdY8WJHUWXMcnMHu0BZeM2E0kkTNuXdPjzfPcWJnoYJ6zG7Y0Attc23D1Jp+E3
oGthb7IS8DfeP7gtupcV8kfgDKY/REMTiAN2orF2FiOr3sFHNH1RkTrVxTgU/CgTvZfAPjOe1sMD
cavxwBWcIiP3GTmbdO8YEW1oBuLoXjYQSWZxMlmai3Rlu3we73u4BYvP8t52OTqqxv+2JMdx4hSV
TtgPgVr42FmtGfY/RBJocJxguR3skrvkjMOXX3GQiCH2H0AZby4qv3OKp2fWEWKYRa5P/490wG2Z
s6IdJ25B+oRPH8Z28p7ft1ssU1q0ydcduLxxhWBSUu/YaLo2hdXoc40PqCrraftH66qXXRXto12L
YDZz/wLnqFxUyMil5oKguzeimBVSG3cX+RzWdj4lQ0Xf4Dsx7kWbBIPnwG/UYMMH25ofJ0y3rEf9
4FMeV5t6wuVYhfbuQzl6ZerYvCUFfQEchcmeke509L1g6qVzwfiVf7PKTbNdXhRSjXp6DNJWe+TX
wx/1b5kbxW/YhAI2PGl+tpUK/ITM9BEDWm3akOfCY/geAem8uUT9nvPiSQ4o2oqrQuwjyI7But2t
Ofnd50FOBlQulAD470NJ5Yy3Uflc99SrAizWegqQQd7ZjiH/UyqPRHiJ82BsCKfHVf1rP4XCmcJ1
Zt7KENTXU45q529hFzbN0mX0QYY35QLXG9Y/RwFCtEi19qmhrLuO6/KHWioDR+7L44j2DLf/UI+0
UseFOmFcKAMWpx6r51iX38IiW/+8Q0bb7aFB2KXLuKv7ruyby9v+xKnZNwLj8QndCRhK3kWtegxm
580Bac5MrJwMKPuszgixZg1i0zbb2ET+9/5M9NGNidudqsQVk8ej8t79XR59T2o8oS/yClqv2Uqu
aGpPYSqErWP/t83slRLmrQ0OfCgxwCpM1bMv+Q5P2oKii/IlNQAD+pBBQDo0zsque0QumsVm0ePV
9mjjLSGzSjhu2T95Qufi7LCojSGOvrl7otIFaLHuq8sASXcvh5wKjr1sCD0uuT9hIOHbeiT7uI91
ooJ/Ip2pKobJxshD7OH2ZUnCpayw3tAd0d0LkJ5Qes1MSTH6Nol6h/YqjzKMSfQ7H1Mo1WKAYSkw
S5EnW9I9+4uGXN7/5Mzpk9LcMiDDt3PrmV9eL14LJVmFyQ5CcX9rVjj1CjuKKOLRpEfTQRO2NBeC
c8ZzqAsL+LX1LiymEkCa7xuErdtcskkcw9Uo9/d5CWRhwG9S6CjgH3xvjDPnfcdWgvntZi6pr4vq
E6Za9RDYXqqbbvwnihCcgKTkeMg6AEZbw188NtOs5/Ubs1X62GpSz+ZX7w+9Hn2OzTLbqESjckSW
kFtxWXW9UNyvYH88IjRI+g5qNqjGytMCBfos5nwrXN+tJXnMDDRp5D1swudy5Oy2B/Q1m2bwRg3y
nJ+WkcGXA/84hDtDMXuD+dDKG9aF9o3HXtldYSTIGfS4VzDwQo4v1ysjeOziuSJo2ER5Y12qKxD8
DDnAG70EvhOI8IrPnN1Th1jfz6Tugwzly9NPX1J87x6znel/jM7lJbnnfC5onq8z+/OSRGYmIZPL
3jqSQxMNpmf5gIvR/mPaCBg2/Jcil+iJOxDpdlt5LtPvQ036s2NmpJjeqM+SthVzwK2LtzFBwlC+
l/McY9G8TyObC7gRMWELtvGFJs5GAYDWidxXGPhhlQ6mUBkq+Ug5re2Jwx7SyNeW5QbxGD/bJwhj
xj9pe3Pow4Lnfnv0Yyw/JgcOQ+LjrheyH9qTcOuTEl4AhAQpP35q4tahHSfCikCuEze/7LJDunUf
J6lwyC8st4HByU7iAVZnKtJxhQtzvx+7aO/epIDZcwmuv2VOO1rK+6bvk0sHm5ZgIP5prrLC82EG
n+tmNWkKHPLAqWu4wKD6h4kLFfJA3z96w4Dx9W5N6us8x/G3eUN1bB5Xsk7QXzM44U2E6pIvlVgL
Sep7YnhpljMwywMqQ0xlTagiUlF1LBinisPm6QWwm5VxXtdKpGcooI3O84GkNR5TsErkp/H6TcrH
JzGl5bPfCezjW6BMRd4CvtQ3KZwzgtRvI3kqGsIEP/tVIt9wdk10a+Vz9IkLsfTjrRY7TmEO6jeS
//G2cQb3sgnIBOh+v7t/Jrqa6IaQSiJo7EjxeVM1327AO287xNqJnlP9xmor+T9VlJ4/PlSp9ZW3
cbg39i0MC+YZuMxTx7+BUfK8E2sRkgAywtxMigbqT9mtgbfNE09y0j+dBqDUdIyTFX1cqsR5wxS5
nGYq2f+H6+F15iDt/eppPJCxXZva+jrMxUCXsdRlI6Zg5O6+vSQakFRhn99qwamSKXFB004d97QH
3fBLfW0ecknqlETBzJHWkCiIEh9klF9oj9pCuA2bjp+ewDwcpmgavJQzmhOqghMMVgYYzuH7NwG8
prdfJTzO7qQnYceVlt9xcNecmsTsGJehH99WrVJofJFdiFQcNSGMKvww0xo9Q4RJRh11tti8bR8O
47IKafWWd88monAKjJP7ph2bbaNP33SB6bM4XrWrKFeKcrvzBRRoIVX2FLHMbbwKyG6jVUpQTlDA
TjBNTZkO6tWHdIX4XjuXr+FhwJvBPIlyB5MU3pbixA0XnZHfh5UhZjcKwY/HtwelFE6BZjg6Hrtv
+BXzHqTtfDVwzzC+0/1MbGyogfV+x1V06wQuWb/DZQ8naMmUFFF/1cehqMpNrqJ1dIws5cTwR6nG
4hHizITrstdchH0SkR6QMuZJvl2LXwS0MfdWU/T9ljKXadMq7jkRGm2JCD1dfoQiziiT76QY0xAe
hl9ucrUf2ebjEQcheBowX3V2rHuPNG/a41AXpuAVY5GQ5uHoUyCi9eGzKv2RF9Yua7sQCzDFMryS
Aj9M1i1/U1TcDMNxANmHpgt0qBfPfVcH78aKhHkkgaENRW2NLbhM+TRZiK3Ksfz7Jxpr2QwkjR8f
O8PasGm/8UjXTzMQKOBpMZCWydtQN8o7raksjBFuE+Q6tWnwoUzFyskq07bIb5VIGNF1ADzKkA8u
QQ8SH/J/qohP96miNWSwqY5C1AMiFHieBlYMffyYiNj+dT8QcQu5wfRfDzsq1hwFN6ignbajC9W4
gCcq6LCNw0nQ0vmZ2oXwO9BXQHuaaFbXcq7GLMv4UOXXYK907uqPz4/W12K/M9wc1h4NdJEF0lu3
se/3KCH39VThTWcHVhpa0L6+gKcykbWLUEz1tfIuq597L8p/HV1l0IPLNfj98ivqqamCjYVDUw9o
7xEk54kJwXOAvoLNnO0xbZLRzRwqmVyC2O8q5q1+z5byYFFv+wgmz4nx6hLBHNTKsf8IEsyE9Rgo
XHB7QiIcPdGPia9p0L0457l40Wso/tOQO8rceBAAFm2wyqP6rJPLm0+eCz3jjU4Tyt8oeutTT8qO
0YPD/E4oiHhLPZjqNiDZQpsyv3qZGEYzYhelY00619kTt/94HabMUFCTZHS6bMuY4esyf+2Zy+Mi
zg7yzvLVqwfLwxkRwkh2oeRTkEGEgMcTvwgYrW74IfBCXH/7ax0foH+dCTlJo4wMjohJ0sVCRV8P
JcYrVG40aXlucO5BYcMhogBsdwxJd50xI/t6xNaPRF+PAQ+YrL5NLsWuGGi1qy0k37zt/lAnSVMK
mMC7UYKJcuhS5U/tqZY/uomEK4YYIeV5Fpbx+6l6vfln+cXgTQwG9gPZD8ITpWB1WwDrPrOlL873
o/kjr6TJFC1lFtdcSsWjMiAVdkfM8Fe5pGzymh2d9Px7ko1/ZJCujT2SRMHHNw44YEQdys0a2YTL
xK5jrs07U8hGrSl8WBG8fidLW0Qx2hYY5VsK7xruMey9sQ76RMxHSdapqZ6dn4KmO8R8scDwlUet
fLfmb/Gv/AKINnn75pphuven4kwlX2GqMAeXpRR5cQ+5Ds4/cAXV+IXpzEIeCqioZk5Y+72Lc+kh
fP/bdy7tZMSVWUqYbZXo9r3ANpGONX3L8xpncGCvuiih+FdM/H/es8UCHKpFA6PnBCDf99ezeTLX
WqZMKtPuXZ6GtD6rgN8qscpzhkWOqRYELuKJUvzlhM5I80CcaLPirSie7aurCMPyMrgCsmfNjPxM
+eKLnmHom7qT6TEgN6hNDqxuSwBmwod+bXXayg0MW+HSZ4KoXqd1ArAlT1C5Y/Nlpj6ZHnGHfF8f
tYMFoKc2j3mQxYZbjSt+5EL89zW8CNcSeNuj+NNOXAIrgH+NrQYKy5wXen7fvh49FNW8t2vy8jvl
Tay1PqMWEljGlPsgyC4NXN4eDeEzuPU/V6k7Ax5Flp4UCQI5YAPiO4Pu66vX2mS7JHpuAlElw4gu
JaZ9NWWvqGwvkWkoaMZFT/gu4xUsplKVsuxGdRtp35AQLfkFGaVK0cYfE8NepwFfJOI44X4G04oe
Fe+DFNK1wERUQlvXXVJl33JO1uSR9qNr9ZON4a4FciOiKO17ZDSeoBZ125SHaoUkkNSqxHA81qpl
J5+Uk/b7S4lYEiBA6oSwoJmaFi6mtplSq7sigQJ+8SqAm6Xxb3FMfMVEyVlOSGUOx3H+u10OLkzw
rY8rpyDZPpegrE08Ylis15Qma0A5BlTQu1c72oBt8mszAk5xfMoZlCg6H4LtxsDEtuG6IrnseJTi
usKlmmbTa2g8RGicq1+J9bGj13SNPhtOaH4HZx4PPgKhvl0S1ibaY+tJrTehqOkgAqiZododJnyI
YwyB9N6LHrnLXap3Rs/tCZkrqKIq5cHqWapF6RGpqGDcwxxB8xJi+CyvUBOWtmTRJQ/f7/1xFt/f
JJrTpaa03vV4Gtkg6mQsJqzbke9ZvzgTmFO3Fz5zDmdyGoaRTK08Bhn45Gk/CoRC5JbFG0avINzI
9ZCbfELeVrOYqoN65/yDlyx+FcnSM1xhxhccQN/OvtIYLh6r74Uo9PfpOfAs+mTYd8VcweKMQgX/
P6HukKT7jVnXyOdi0np763ICBx9DO5vwPDC02x/Bab5mfMmyaZK5rhiyJdtelKjV7agfazRo2QZF
UaS11itEJJtH9kLM3KdB5R0fDMUWmhKqr1AMw2vZXBS+neC5BkqYB87o3Co4oAUdBvSk8pL/9Hnk
WVuxJorz+XUJmc3pcBQy59LG/+maVuW1tepI3NwOpnCtHP30ECSZLCN57iwBRuBNOAsH3wQaPy4e
NkQWP4zYZwAFgxRTAlLtXF/cvhCF0uM+sukQ8O5UPqFFXJ1cO0ld3kssGRkxkLn1PHVoTkax8hTN
bYhmjwj2UFjhuQzOo1vKmoQG7qCWf+a5fsztOUhxJyaC9fqdA3D2RLZMKaUkWPtxA9yyPs6EWSil
HCX4Z7XWJ7N2nFW6KF1BHTXsKN2o8ifqGsZavM78LK+UBlB7winzo7aZh3AUrwzfVAjMEsCot0fk
XNqgcHh6nfFfgesifOXD9IoK+Ustft8NLUqERYrvpqGjPtit/V6ruCiM/m82w2t1vnF2noPYrhXr
EP/YVwrlho/qbX0fefaN06l5aS5jNSKkXQkOfO4TAULvbj27GHhDlbyEFXFwMLh49CheKuS0xBoi
mXsaDLqdE/7mBelVgAlUeFDnbqSMaAIMmn0tWEvPpIZH7FWyYZkvSWVmJnAy7XCOPUh2+RK6Yh8R
IypClHR6uszVXkTigkHkYkGiE6tlnQpkqDy82hwCMkMErQtyCCkvYNedj6s+vzk8jctQFf16aoE6
Ijz2yTfZHerL3m7kPoyku2EgWxlZLdUV2AH0XzIu/2ko+jnf4kI5X+SiX5Uo6XV9PN5WuhlWnY2n
wif8wrNjPecvs8ksgMfALRFc3GOuoGuSk4ad28OPT14domG9o7pUp+TXUvlBnBWVtMN4Nu7CyKsl
Gulc6SOxjfAkG5UUmjNDlzNDZtcckD+8yBz8RNR1/L1WTdTxdyFR1QjtLPgmlMIcdkofqJgJrkeh
A0BSSmqu7VrhRtgG4pfbSn77I8EmLgbyi4dcyfbBcllgMuqBh04WoV9UpPUM5Rr9CDqtraKlDSt2
G9O31P8gz01yGIDJr1HWgoiCpoMorWUaZErOmaSWueyOKvAbB9C50oYNDvCggyEhIYMMrDUbvsXy
DRKfDA2IKOAbfo98Joxs8SLY1ifndv3lwcft3wzEl9G9qrI0r0tFulJRTOaKrv7XvttXilo5hS3M
PUrwrPY4K2tfXRI6LZJD7W2my/phn7ByUtAwbekpnLkReN/OWh8sRZvrFFnI27Dj/kgVXTpO3zPh
m253FDo0Id7CHTuJroEijsEe0sHbM0zOoDf/4EnH5aaietn7Rx5nXwCyaqwuvdlYNVHa9Fu5cotL
AH8sJlzrnUbLsPvjSezU/eh/vWuqL8mq+dmyW3UWMvnOyA8ztbX8JdINHdtnBIY7Is4KfWxMNeXj
RC0F1z4mxs52lkeFq+Z0nAJMN59agT9iXn/N5mir3gqS9m6DwyJvL7nKbFlBEQK/0QCmv1LFcZen
9iALDj1ljVfhV9JDc0je8IjEW5zWVBq7q3lGAg7dF0HmtZZKmY5mxyCLm3HkFMMNcEfpAPR+c9Bu
O2hYVtZc4Daq2/xiJ1aDR2JpLRkQ+GwZQqgyY36i2El8mR7YZ08kZFZYlT33XccL0gj+6LpVwEAb
Yo8TzqkspUwnZF4kABJXOICYt8X/37j3fOXRJi8QcSWJUfgj4BJ7Y0wvJb3O+GwaexG/bhIqmaWI
3EAsJvZqp0QXDriKTCHoltqtW6FwbpLvlFrd4teu72l0f8g+WAdNmEdbYx52IveQeSqRyqPK38+X
1Nc5jw+IpFShxTuXVUTSndx9z6UnRQ/Dt5wlh/lb+Gf9sf5hJ4VCRvjYkx+kSDOOKdfLvm36EQq9
dFPpdgAbBj62wxp32VHhzTPB2myv9e3iOcIQCTozoMMcXZoTa1xtu3TrnTtOcd0Njx5nlJXFpY2K
PyJmAVIvqiolNHYMalvbs2EJlXtj1ySKRfqQQTtIVrEMvK6ccoxD5OrvD6z7l0hO3chSN6v3fUxI
UclnZWmHcI+CtuKAhBFjxeP+iOY77B8HryZgc+D3orB7ggg9yS/iWsaRoImbZ3WKZ2BIF+QO039t
DfUfYWF0VzZR2wiW5bbvy/fivy2HB5k0UE51JBNcvqV5QJAxzn9sZi+vSJQaN+7wXBeEIckhNOFD
y7VwnDJ7r0YlS5wYBHn/f5TTsI18SiZzTAfEoyOEZi0MhRZfC6iJIXwTYJ+GewejCF43L8s3syxS
lYwtptjbqr9InZwV9NZeLwvEFIDbA6g1z2+6KObqG11ZEkp8mi2/MCsJhwPva8CUh8DNOV2XZrF9
6FB95vGPzNSwTurws2HLewhekfW3NXQO1KYFwrFnyfYb+yQOuI7eQssYkgEyZPWRaPr9HEOK4gNK
+BGbj2UZwaLk+SyA7DpyBbExiJxKENqKm9jAjker6myvMZ9v5aIy6oP5LHvRz4dpBFEs1fY9qdYP
tRY+qHFApGqeO98pV7GCRhIsInaBeFhvbmH2XDOmXwk/ZInFhAQK891dtW7gA1KKzrmE4rY+fFm3
s5t3OSJsvOkm6Ac/PFbHfiw9nNzneZODkauXg2uD/UR8dHoLLpWN4odNnpZS4H85XIZwNYg4CQ7E
wd81NFc+mntHyF8ZFereT4A4iNJXgDQfTkbj8/bLLGVohzsDw0z5phFtPSA6kpYbP4Ghm6+voZj/
6USNUkmsCD8tVTAgFJ/IEdBGQXduuWAjcYPwqOWqgNxI31mSfcfnreH47ulz56eitvs/ajnPS96J
ii5gPRQpD06MizmV6rTXdxwHV51Bz6R9asyGJaCTyKsUlkGI4Jyb9U/seeLKNhoA5HeC1ApX9mO6
XRu9HHasA4hyZwerazL2g+TahcfxiX8uHql2nEYMD+oGova9uRmArHLwSO7k4Q897XGbbZVLyRpJ
23tOYwSiThmyEF4PtjhE81d8Vn/qWP3mBvV1rSXMlIhIuYVHj6afBpQO7kbAAGlF5X68KekOIAzU
Y6CVhDQKBQtWHWexG7pn5oTJ0gMMblaMcIISw2ed9xcYzB4FJH+IOzc6kwq/tzS5E3L8fp19ie9j
1Jww9OuC4th7Rpam/q2+LmNTJn+ss2jufzVHWHFjTntOXOUk2aha1Y3rFk0v900CQS+jXYZ5UqFf
iTjgpVU0lMjztuCqlWlDyox8eMNo8RFgDq/g1n63vr72vcpdG8Kj/ChQCtGhf25nY54A3o+Yz4c1
/OzO6z71dw0/9ms0R5+XHyKW1eoZyrRdN+c09zAu4AAiD3cGAZIiNdpfUcofMsCYIJV/NvCt6uv9
Galwqh4mashmtYqKpbZNk76nEseQqr0OmDj/kecPDsIhy7XT19nKeXXQ6nYLoRBrCHWzhS6da/ID
IsFb8II6uy8CxamqxnVFA5DwHx8gVPjVKclWc/vtkKtXZ93P+XJR9dBEFdzWPIZkZKp+eLn30ZQw
zhbLEclcbQuNIYz+NebWSnFVfr37bImWS3dAp+BNOoEIOWEpPp0N8G1nM2VnmT98Jaw9n5/tyOy6
/E5Mesku3li3zoQkIJbo/Bd8f6ydGvRzGKbB5uVQi7R6c+16eXahDbx2GBLVrcKjKRmGu0WsqIoj
9BD/CUBWEMOcR3W8oYGEsWYRMEls4ESkNpjN7tpT01qs2gCsHBuAwBxRu27w5Vhlv+LAOn3FV/cK
Z9ooRRhTy4hVQoDQREZzVBX6sqNdUXtefGa/o2ZCbZ3Lqbi+OSvzS0cOHU/O68LSBAOX6/7tVxNd
w8ov40zxlQEXQl3L+qyqGIlO3iLCjgYxsF+G8UPVewfNrYPhnfGMCHH1K3fbcRMLN5sfPTG0jU1U
Fp1XYNuShei/7QoO71GCR+NwrzQ3GQxozirJo/6CyHZAnVR/oGCLCzqHN/gY4qyyqbJ1Jhy1n7OM
m9y5z6WKrv87QZ2g7P49pQoxUgicNcYd1e7CKU4V3E0bDtsdAbjdE00vVbJX8XnTd3sHYJBoe4PU
xyy+mgkQ2Gq2dcC/8+d2mBbmrNaK1ayi00hFOmwYsplLGil2SYr3LJ188lJDX4c9/Qvui+w/He3F
aHskaHV08fLDP+xGVswxTSMu+T11VVficUp6Ikd4GF2w6zgQUmf1N7tGw2RZkrQmi/CspFqc+zLj
y77aP6DCCC5zqqXR4NmtOzwfHRJ8w7Zz8qcB1G6ln4mIHaB//ipToBALdQDYLy3C1A0IzIT2S74l
s9+UQUuciMEJ65YPfjgdph0j9/mu0S1bhJfhndnI0V4D1czIZ5OgWioErqhZzY6gaOJLcUS/S02M
t2ktXughlv+rSOEtA9s09Lka+8/3CMeDVynCRojYA3i/s7nSlDOeK4Mp3yahAV24oKTKNoSgFgKw
Gj2RJKENHoXd1AKyqWfauQXOyECqbh9wDkBehI7oG6xhg0udp45caT79Mr/E22MOo50sFrOmgx70
BZySg97Ae09YY+lC0G6th33jmqwMzh3iH8StgcbcfYN+d8PqfjWpRrp7wgYsiT0Rd8ZquJN9qpHr
W/Jf97CQswW57dcFdYqp/i+TN6OJioTZoAcNsS6F7xwhXCW2pMw9neJ8q3YLRBHFZLuYIehUO/Gx
f/E8IoEq5tZgMxttE5MhsGQA4JpNkLWbO8Vz531cAqEnoZDrvmAJfb4sUh4qYl7fa4hmzMmJNeAl
+Imhg217gnZLl0bl6/7dRj4aEN1a2qaCYxvK3VIOzhamm2t1pgyuAH/tN5/OKleHx9A9N3jlSvLX
KjVzFyUw7nVTDasSA/uoLl9Xsrj8VvjjCSgv9NvcGijGoDlRScDHC6YtmJKeyu0wVLH87K4sX1cT
rwgUE7MMyBCdAYDzH2aERlCvDCpLO7CTRdvoE2+/KWEQJMCxz+od9RUW9Tfgy+r6R9s4iZXls7xj
zdygip5i8+eLpUi83Ub3Re8Hwb6tT1m8/xq/dmddZjtRnzsEyDe5XDSkXufUwzndt9cXzRPOIKVW
flons5vbww6ivy/PtGLTWEGokbPvaM0aNEDGJ9UpUEO3lNA+0LHa40eL+l2VJT0nSLv3nxGi94LH
mhBadeSbABed4c/7WoguqHvUx0KqOWhal/46oXG9Rfd+r9hRNt6xwWZIgGqQXI5KeMuJaxc2ZjFQ
sLJoojmY0mOP/NxhNuI1Ehkrp1lsMIINCLo8xWFHax5te53VQe0xZW/3Uui+FT45RwFkDj7vOoPG
YkDSYnQ2EI616jdAKsudxL5Bx4CKB4dldtN+000Y6vpoUsICk1acjy9UrsBW5aRI0GIsTmfeDozv
HQwS4iUUG9d3HiuaaW4GjnyxPYFwe00zIsrICMuHa7MdNOo1TgErrhzGlXA4rCt3lfCct9K0FDxu
aB2szr/YoHHVRO2qcNLe7rEtrbIUpXTpIo9enBDqS1SixqsaygT2T9T1nVYrFhmJlanKvY1Sf+R4
rEJykjjCgcBnrCJMQLMWpnyNRY6iDKmQ7n4Gdc8rP9otbH3vs2X0ssdcCu8uM57/kXihOoUib+iB
F5QlvwlkLh8BMd819wqWe/2dFcS9RA/BZrQvv8tW7fEsxMvddm79ygF34P/XQwzpxPm4ALT4kMq9
lngvVqzH1bC4bKIWqb5Fy/lAeg9UXNn+6cY5LIhDzDPGyamR1Shs2pWuT0sonMRpJkyD8arRNHl2
WPE8BWlNekE/sxBNayQdvGSxCs6jeV9/ql9vLCg2hieph771RCvh5NeVkZZ3yq9HluQbOwZMM1Mh
lS9E1enqs1XSkFWzEWaLmHlUXOktww1w2bAvRmgVXGADu3/L+foGrRcrcMXGsCBnjOmP4p6G9Dos
ODxjpTMuZjry7XRlRZ3M1smagK9KCoLNlDyDVfhR1qVFswDHgiyzxLQRvPsgz+ropKc6rEHLG7v/
kyGk+hIjyveyk4sEs3RDeMxvaQntyss4Wv2x8Hb31feEyKf3kwXyr4YwyPoo4LeIZYDs6xgBfg1U
iZOfsf26nYn4t2x8BcS9BPY1j9h7VkuQ96EwBAkcOaVoH7YZyDKNH5kYyeJyPwzqfjGndf60KlRu
WKNG1ZvQE4h3orsFn6BblVdMri+EtXwtvEEsX4Noplo0F0Z2IsfQY+ajmdyooXvBAXCrsvhH2rHt
6i2Um4Z7ZEob082P9MAQ3FqAwtOQ6SnGohxnM86Vym+4jsVHcOUfUoQ9GxCV2Uzolm0vtFXgaSkL
futOD1jVTFxbZ4Ej4SFyt8AiVykMBlBOpvvuvhcO1ZKaCcHYBpXzShp2YVSFeMLoEJ0C7sIVxbdD
5383nIyCnON027iTlO6jQKVHGDdO3U2SCXCzKUhS1OJ9hrqiMeqzPQysZmWGl0u5usrzysgZYv3P
sbea781yU6Mdh5Dbbs9yR3I8CLpsNxUWtIFbj2yMtROl4iuXB9FhagmAshSNLxsDJZ1Ee/WIqsQ/
8yC3DX4hQ/MvUOskERoc+wPwNAMVTGWRWgJbJLIy0I6O2mvHe+AVWRW9/2UkedTxt0SSCLxFX+V3
Y5XVWGjn4oxPXbbhK4uz8NdlGH4N4uPup0wXsXrDhIJLs+HAWpB0+zcAKtxoRPipsT8Hi9d2IyBi
Vf0J3boV+YI8O494SX73TnmcP0gXAbeH6or4fDCosEcKlhL3rZoswBhWwUgiGx2+7gOKDRsOt6oz
PcNFXsYxE9l221UASR6wxnPPYseC25PQZOoN9KKh53siCpG0BxeNqktcZNV3HiOQDb8HkTBBnksx
rnR9vbVHX4aKUpdwDGOIdwPVHnYRXBmZSTKx+4A9NwK6s124Ml+XQknY0rBjSepcvr4VBGQfC274
H4xWi4Iv4Hw1GcYGRjggyZTJzedJNI2S2DCuwXxNzy/xLU2gLyNPMWPuf+2dw0b2dKK2ggpbx1KA
7w///4A3tPDfgA+yb4A4KKUyoZZNhEFQmUI2bc2f8k3FsbW18ar9YgVI/W9YIPSts534nqL6y7/5
HE3O9d/bx3ezBVlLN/X7O0/UnnK1PObhh5puLBBYeybsI3scaKVe7YEsUQ+RN17f3FxKGkMaQjaw
ofq5kIqyXnN57X8PvlVEWgVN7/IWm+LHne9sYCYJ8rCllOgql4F9zzEOCszr262O8mMpyCspH0cb
1hOYDeK8Oo8drC/XvJGEIrjKO3izw6LS0VLjujaExwP2anWij6YL91MW8IbvdWqkyFtqpdXMnS75
6OWsDt14EUHUSc6FrXHqVzshqorO1aY/CQwUksUEEjDaMvugGyPwiPXlkDEwP3g2CJgBf5omtz2p
7H/ABn1VKBKlLS/Pp2I/+xf20FSjxgfFD/crdaIwhpuLZb6NV1fN45hrLO93Kf1DptVpzFRUX6NL
KvenDzfnDAhy0vhUKUoAv4NBDNH9bLuja33rYuEHwPg9mAxAtUC8BVMMHUs+RlTT1vaISH7kS2Rd
xuzlIfINXV8hT0oI8YVYFqY0znUo6vuM5DCEPDKzCGuSeTJCRzNd1NpLcRzVrDwkw/CQYMBD8MCi
QAIoWGArUU2+FgbJb5wzddHoLbMr0noTM57vFo44HMiOQJzKL7P90P3SPOUwmCrp7L11PDg/4iD7
PV3HSyN9APTgk3GoLUtbYYVQ1znrr++WdHV6RsZIuH4+dAbnDrRr3w3Ei/rT75iDPEGGjvt/kGTg
fNGKPZP8KRnupynIlLNuBuZLipwBGuQ3SZX+T+IeoxmCH8j79kKSISaPPmK6Fdc3481gdlVZiwd+
puod+UhekBlq6MJhfa3/ZV0qw2/jv9O7Wwsra5ixlgEQ+yVLxJhoUTw003HFIdMyQSNrTgFAQfDk
khV2xuSMY233tgSlS/o762ilDg6LYIIHaJVy2Pjk1NfYyY44TjEVqY5x5uVfIzNQJKjiKce1ufNc
/3gwMfvataoRHx195PPOrSgN6gekYSAgOu1uH1m3mwNpZDtEcfLU0rXLgxM5GCnBVJtAQFVoC/Ro
r7jLoUlonP2gUKuHQBMpMP4vQhtuxoYwyAmmCzhLjubH4jngWz6edLOSQYQyQbJ3eYVHHmCu+QgU
4N7i7YdJphz6kc1dlnbzvXe9vXSHYRRhUZ08c4MxfGS34sDhYvHw7ZhBkuiHd64CiWA0dHfWuPsj
mPIb9ij3kCMVAY/UT0wvvsD2L0LGgZQcZ4ybcfoURYVfgB2vk61JAH0Pn5ChRm5TO4i0Re9MsNcO
mdKodCr4F3T+DzuHcmrCNcjpSnBi1Ttr8BzbBhDKfHMVNfgVsMeOGQc51tdjuKzHesPMtp5wtDWQ
MEve8UtWU7r0yv4gheZnOQ+8sJLWIAUt7oW3042NYtizvsCZRkdKq60YEqbEYMKJwBX/RTKRY40b
ZDi+PB+/ZEaoImhULeZkyzprnWe+pXD/AkYrEKr7F4tzw6we5YhWyNX1wwuN2fT2EW8AjYq01fWV
AQZXFoMqJMinGZ7im44z9CCqGpAgnC0v216uWTqnp/Tq7uNg1heIGXpYcbbGE8qemvXULQSOJK4n
dK2I3t0FKy/BHP+fxcmVt8TPI/9qRdyIO1jlScFJBOHaKb00cHiZqM0B1YRf/L/ToUGVrdsoyo6/
KlEuO//e0IDvYszRDEciZg9Eask8iPYzuCO+KkVbhdKUiCXp0DCwXGAsDInL7cGhsPTdYM5+kagA
au8k6Lagep/kOpxu9MfxrVtUiO6VQ+uYDLKRlaiusuv1fYSLDvaW7001lhjpElg1lEyHLlWMyWA2
VDs6FuQbDv4TeslqVi8zvmES0lhFOW1fZZkkt+CqOXZ2N34t7WiwDaLfJcDpzKVapPwrqqHcUbp6
LaWPPmqPcI5szcxXWH5EwlIQ0we/NjlNwNDpQ0qyLu0gmWAMCkHrEzylKFfPdL4sxuKYtlkeEnPV
yaY60cKczAyMq/ty4DIE82/A2gg70HcJCZy5v8g0nCv9z2inARIxT5oE9XWVOePPzLEIVz6Z0MOv
ad7NKXC9PN3zLF5ayAW0fshCyfK86lWPTyBnxF9fT4aOieisTDu1ixdzH1bxS/7Y9PhrY6FQi42M
Uq+mJooLVKOznomsdJhbdWUCnaBPw7QkPRCsH+Y7HgoN1cALlvu0pCuN+5SBR9hkwSmfzgU3uY4c
7AuMko5GhAPBxr4b1SbZ+wVa8uL+HP/42+cSz2e8cqBDCRiSKoLDWVnrcvp1WcbmyRanZJQTLg87
WHtUYFBe37IqKEanwDBTM8JielUjJrQf5mcwatGMdhy48PPXQz/cfckmUMMs5Hetyb9MKJAIOjRf
f5TrGhEEP/ufGh44QuVo8MKLLWoB0N/BWUXM7y/09GdMuUo6g6LEI/l0aIGlyTFVN2pb/qCIanHa
n7arePCK4Des5XyZO0QMYygdlP0/TDjlL7SVKc63v00V4tuc8FGwD85rwmniNI2Esi77LBZe3GmA
xE+LFdWIxZgkBVV/hkmxlkhTwbV/6yF64jJyI+4tdXHVRi2boRkd+J1tdiR+gYVpRM5g4fcXQinR
GnWdy3JkVvBDGiX7JRdaPrAK+766HyIPqljIwhkpQrPYiA9NqzsdK+WqWmf40GnsXdA2TO4lFrbF
23wbgmRv4rkrcWHTLPNh/3IMOTC6O1qtvjQfeShTwTLhbAKuihfiIKCB1Gtt4V6EuyjvYLdoed3t
VfMAoTWXy2sowzb27g1TGTO9/dI32LKFMyZbSI++W8LWdClQiVtuvyAQti0flIij3dz+p9r0pxMT
EmBfmwODVqDdoWxF1lMeaGp/IKJo4J4U/bMBI6xShCQu0/9cGHSrcponDnMYSa+VDb+ONDzv2cfR
AzGD9Fi53hJlA/gfZvT8HWwGIhYiXBM9zuJUT3BxOwAWWKAvOVJzmQ5y5m5WTW9NLpdCa+BoLMR8
U94XySUHSUjdUnvi/XXJUIRwEI6JZuvdanBp2JFLgF7/C8NBIENN622XX4tmUoh5f5DWEA2JS9cG
naTH+WFdg6qcdcyIKpDPIDvAWkH8wsMhxoCXCUjDomEcLEsuG5pjUeavaIJAchtC5zB+HfrDZCpj
qUxDKTZRdVwwGrH5zYdXlzDdWYZ2hHi9EYaLejfKRBeWCiBagEN4rPPZoeQcZSMARqcG6TFraXxk
aO4Xc9j+Bp4lo0PFRRbafFdG3evX236E7tzSFJ7C1TYpCDBLVDrMwBvbPHxQJxsp0BBWpQaQarFa
hy+l/npK5PLn4k9201//PtjVofI+BMXhZshX4jWMKXUDdwV7TNpQGItmHqhL9zLBH3pzAqW6LRTE
eoft5QPpgEAhdhe/aQAx7GViPEroE0pFV2u0zrduGPLMr5eqP24PekhoM9sqL/5gEua5mszmPxyh
Wf5vOJR5hWDjkZ0eFWyJhyqkcZjW3bE//+eh0HQ817A8WbbUDrS1nKbl4uLMmmpFtIYSxWZUYLY7
d5nFR+W3S0TWmJdBKMBGXBM7/YQF/o9eaSCX779SwaVyiyQcRsheqwQtdvOfyZGKVERhNSce0rNX
XaPSRhV8mLS1PzdFPKi+vdHKhMYexHFUFJpkkLmrf/R2HF2GRBPoPa6Kw+OwNtgbXnRtyQGm9+jo
BcwF9qq9k0C3GncBb7noCsh9NiBfMoZtfzYd7rF7FKj10kjjPrW0Y6OP7R0h37jeFwm9WbEIiGvL
wFlTpxyyETAl/HqMtwen7dDerS6x7v6iu/blorwF9wkMI3opw0kQUAXrhgmwRxh5lv+/HOIakcLs
jg/jkZ0mkXhMGz6V56OC6PVtEPDKsocnMeZCGJqas6ieaOn7XwRlRNES8yzQzYvPfdOOZMQBqEDB
oBF0m4lUDAVHPpv1P4iCuWYnHZYVkuU0jUoNkead3QbcyP7zpM25GECim9gWbJMY4gQZU9pMho1T
LaXRMBkMlzgOE61D7SW6UFyPltuU1NT0ITIWPz+waq2rZwKXAklSah2wKlwL7z97YhEgxCrtUS+R
nUF6WIrO+RLQaYd0PhVwENmit9YROTuzSf0x22v8/i+RugGhg6y17wDpKMcg9It10JxmsIPjnb5o
qbSIFfwJceYpxrzl3ShHXm7C+0yyQ0geSu0Rm3RABrx/bPl2YNLrl7cKTYnKrHrg3tiCUcWqOYnO
UcEUkFd0IKvdZEOKSTbFNIYiMlbIPQaWg3/yz3KUryzp5QWEO50s5dCFJLT9wZGNpWNrxNVSNX80
RW8qtZG95iisn7WoaYOplb/zYWngJKeb9TufrdIp/MRJ+3Xb9pDJ1xO7I1rOv7k2kp0P1izpDMsh
pXmCmLmfHNZSaonI8k8++mefXdZXPG2iBufR2uLMHsXmWiWpJiwoEM0zB9IzikBzrKnJR9N75ZRS
QEUkCrXNzafqGgQ3Qd71uqrOVmKO7u4K4ZNd2V+H07y1i47Si5+NBNFX7YMYV1evHm3EB5IduPvu
s/7jcxkEOL5Txv3VQI8KQ9Ek8eHu8AVjCIFRPBsh54MwWmV5e3QD7GCoAxFswBFtWu8gZlhL0nDJ
5xHqGEQz9e2vktUUp6enps94wooVZFb3vpumjE7R2WeQFIIVrh/a+LKRmVO+isDG2M2L9CYSpwa3
KwXU8rIFNiGvstU/l+VnhZ4HcOVC/V8inko/N01j6KNvaGMrcjXSb/AKoRVi2RXUFClMyPiVcN8B
JViW0CORH8xJzF/Xf2XAwcpOXZWqrkLBuQ2UEOM9Z9tSoPFflbMRwDivNxYXvRhwVnrifpGieHTF
Y1Fw/ONUcfRrpbdvB1wXVsmCIn/ul2EMsZPIsR9Ebgmh/a0rtaseVpC7REpgx4CF+vsWxYCTq7/K
2SEqVC/uENsEYXul8DyCYw9YASnMFg+JX82qE6MWj3dj20v9H6lh/+T7NPkm1xOWe52H+NmG/XOj
NY4c9C6ec+XXw8K5TkF8HNVxoDC6q+3piXGylYnF6mxTU2IInCss86wYaVAQBzwfk9+zYge90ACY
ZTbXfLlSswjezcPlhhwxD97OiwpEmfh12zw1T8jDuEdMdzNad+scg+A+LUEeZHa1cOINYECet/rt
YVBIfZgGjp6s1gGUk0UuW8WKibkbyiaKJqZZHgBBeIQnO0SUv7Ndl1Yua+EIoDLWEjtvtPC/XVur
Ug6CoMFlwcILN/DrGYeKy9iqXE+j9d1d+wGMm6GrjnMQozaHQjoFpEKijqFRVC9w2Ntee2g0y2uy
Gcr93vjucRcPs7eWSSBfkHrlKh4yEZP7LO1k642aJwvxcQDRCCY9mjRw2wA376HKKJpBglB6+dni
Qp1rHHYZbeQKWwX3qCJ2LsVFWxSd2xkMeRN1E+SIEAc/bOtYyAQhtV6hFoDblzEMFY9NSFDGZxGI
/tIVDQGLkzFHZ2gAR2cPuO1FSz7W/tQ8P9HDL9vX8y0C0sZWzLJas2umXK1mkW/Rr3lOsNrI4TDM
Fayg9dkb0+U7sokBbVLSs1RA+eV0Lb5PYAYy3sDh227kYe/tNmDT5kX8AeUa671odZUl1+YL+5dk
P5vg9KbSImvZ9EDWFFW1UEJrNrx41Sq9fjaHikfTbciNxktZcAQNf/98riOR9YBwStl3Ki1IFxCI
Ju4L1Vv6ia7ahT0ESjfQgWNzE7nGoAd3T6BMMg1Ab8Ou23NSRmP4itd1BKF0/csMb+zSZVPx2RTV
TpPjJ6JYYR1he4ygxWKGEMuKB+0LxgBAwxFRhxwAsJW5a0+Mffdyfw9wAxpcaN72l8CGhkN67MCE
Wi3u4PBdPWCyzRzUqbgQ/rBtPabaj2uezQq3aRQOzt6Xi4eqqlSz5w2yk/XyejS4MrUHFDONdVXB
eP68r829k7sax/hw9TR13aadu0uV0RHbYydLRAX9E1dWoU0CwsIpcFqMRNZr1AIc2KnQDqaER6cH
sr3g4SAUHOM6qClFebjp48JBBuaa6GeTDyLEIgjl56WmGYtyTi5IjrWDjC3lkWpzcbN24y8qJ2n7
COaPpH2M0QOf+xIpXmu+ZIcDjTT1FQAqgaL86nFoxtdzOCJiQVbUA730HR/I+NJuHqOcCzRqtlH1
/yZt9ouip55GqvIP/4ChqYZJfl8ajjaxv2rHyyjP5MZAoL8UYPHMITfPb7t1Li2dO/IfS0KpqMXL
5YQN4h0HXxFXBy4lVc1QRmFW5g2sRxrC5A7C+dYtPlm7Q9yQGqy6g+p2EnySCkGfz0N6dk2OicrX
U0h66Y4tv8zuuHWUXpg6w9kQjKAaZBdPhU2SscO87hMZyap0FTtuhwpu+lxqjRSanHgJ7X+awk1/
pcBXsAdBv9977QtXCEu3M91onEjzwwAyVYQpaBjoR/N4GI6aEDzIFXlSg73WNqYSzYDJezE7LQSj
PV+Ma2PwD8PoRe+7e2311dNqeT/2Ur0WymYrqvyCG9SOv09UbxNjOqWY/bmZe6FL5BNWHBilrisM
ZLf+oksTsrrb12qe775iuFMyiMrLSjR9brcjrECAt8v4Y50IWg94FwqI4/AOELtHGbnXLPFtmbmb
4ZJ95Kg0LpZlHcJwGmfL06cVuBHLLwYpyXGDwWZtqgzsFmFrYY5yg3RWwqvWFGUyHqDNm8CE476x
oZytspKHFNmANDVBEHh7IK1Nt5m3X7Sbk32q4+w19P2yZOwujHrfFv1cdn+N7TO6NKpts/Wn/xTq
CisLklcVkrTlLBF4oY/FrelE3DSKFg96IhvWMxeHcIUFaosdOZGVuaVnXqDy0T8FC9tST2hv2oyF
OjOKBr0ooMCL1IB+PTRn5yRkU4gJ3juG5Tfk4WsGfBaUUP+p4jmDN0GeK+lLRb9iFNfx1Rr+u2C9
o4KKfhlG7GCjL7c4EBCqVrn85oZsqXxV9AxHrIdywbNhi84zFTQWoqWlrUetrxUsFXmHx/KgMYfV
T/y5uHwDaAVaWB+vlEVAQpjmvQC4H0mc00gI+3AJ5lgv/tr1V/+A4wkiskk4fjTOizwMPv2B/8il
FhsH0YHeUvPTTzdfwA9NUOpTv9JxUJL07Y+QzArl+qbdKu3ox3YURJMFJkce3rx33U6j/Em/V1JR
T4Cq1aPvtSFm0mTR4ZB23ed6+Gyk2o06Gvh+6Cmhg7YmjlMTo+J1gnZTyNc8993nPatyehbmehhs
fWQ2jJ3WhSgs9+oH9eOsHKK6KVFTcsfmC1Vp8YmvHp5Mk1VK6JKt9SjN2+88sAkgTAsV8x5RceXd
3QP6IYnHeFOVaA5U+SOdB6FR7hZH8N9//vydoMOqMZtXadRekrY+mAL7INHf5RQf8qVhWsesKOFZ
m4/NcLrevdASvDe2I/ygUyiWQSGMMacGFIr8xfVw8vZKnF/u+PFavZljgQ2TnT5Oa5eWszszOXdc
WEc2+h+OwhzaLLW5r8gNma/4+INmymh9mpchPFr5Qe+a4eLbZkO2AiSCc36rvNAD0eeGigZSC1xX
QVgaYdJ0g1z4ky/E6EsvXNwyyC5WzRXTEW7HiyL3d2WeiQOkogmRXumo4nbjAC2DbjITRPt30FVC
d9Fwfi5OHmUwvM6RNkw6yeOTCN2rL0KvJS/t4yAXQ4qFxFp0cmZPqsd9U+e+QoB8VTAWIyFbPW/3
XoCMgRcPHe7wU9Nqn5tprXy42HebpLLFhoxtY3Lzk3l6jMudDzg+eqDt0CFtRwoJcv280gMx9tQv
lE5HHUTJwSNvaTfhRKQtZ29o0+BQfiGQzFe8OdO0I3Go95qSTmWqXdTpSjX4s0+8d2vv0VIO/PYH
JB4nE6ZgIYBz5rjMPfVM+gkkAHIHp9ecG5VGSfLwQiiF3MNqIm/tLc2LcZlSvJQUaJs7Lf4EQIox
8Vq/S8ey3EPlRq30flyqD95dvTGAQFEGeZFqDjYlSg/MBJ7s+yQkZI/diQHkszBe90dssUzwG7lC
V5dGIbqIi4Kaev7Yc/S64uDvsx7Ad692tKeruCt/2HhMqLFm6NDktKL/T5645RA44vq2cmgGhUmU
TcgKBOo7pQWkHUUOdJje6RYFvReIwoQTrRuliFZu3S7Ou+Y9tltjkhTAdzKtocpYctt2msjmBiw3
aPA6iBYYqsRdugnatqOhQZhJ7JfP0EbEFiCnYXGvk555z8eKd21OLU6epzRpu7aFeZq1QDlTnC+I
1Z0bbwwJs+uYFVGOiQx0W5+AmP2mjo3IttK+qzRTb0CUw6axJXKz/5HXpP/WqIS5+kefIr3bw71r
0RbKYtVDS8hFNE8fbB3GbNHm1CdZ6RjauonKmI8xFuwqsAwtyxpJOe5yf/2+YnIgjXUew2xyr3/D
1yvNY4V2re3hccAM+FyPjemNs1FwJUou0gj1ZI9Jycfv5Itey4vR7Q+xrVXaT+STJqTNbbfaUUAs
MUN+opc59JGCFknHGfJbLmwiLyeOfWGHXKQP2AjObNcVdoavuj7fH0rMRto8vcU+y9DLwcx3y9PF
AhKXoyU5n6r2P7G5GNWArUywDJ5x0Wk1LQ76zL9E6iHrT+yZCJg3IvN7OEkVO9Ls7dkTjFAEzdG9
QDUc43PnzXx48bEbu34ZznrOLBGU6fmssZ2fCXd8RM1ssECfwU9UnxtKBFeCgphFqI6Us67CDLWB
ntZZ/SAnyK0tcr4AsnO7t+qqHLhVFNO1VKzuqCEustW0H5hMXo9ZwQ6s47fV8H5ik9hkgydWH1mz
YMxHqlL6a19+PQ+ZAGRv/TBEmBuWQGfJexOvcbo5sd//j9dotJInrZU0sSJ+FXRIj2Uv0WJ2GXwx
OKob3lT6QpLWNhU7VKfdVzMfCGZlf83ibcj2RWqh6qjn79mlbcd+/C1HPVVBT6p6jTKEpyve/M+2
TO1dyFnFr9PUDVw/fbB16Ql6i4/B5wux8tHU1WY8LtQYaWO2IzNa4OMgES+zBVxbN6Gte/H3AORQ
mtMs+g9CGIHX+T27se242MSPhCwOjYJXI/GhZyqvXuXCmZ42cHUtgRUL0dcomB5ZWtsGrsboOtgX
F9bmrRgnVvngRbZbVgPtSzVUhU0hIrj0rhzh1jIwjsxCyYOU5QKmhT4mIxhwH/00m8r44vFlqJnX
bNdX52CpY9ZMhPPNHviIpksqEZ+vfA2sRLGWCGdRi2Z1rRDSiUbgdwDb3xHR/FVwfDvl9Ywlj9t1
mmj30Wc7TBK/1D07j9nL4FefuuzQadLpYEXuNTgsgMlZ7QA/PjSh/nmQsqkIL+WZdF/GZzo/VN9c
2USM04NHTpuq8ee6UIgtbLafvyo7rzKqpckAIdRHZ81g/iPevgI1F+wM5M7jx7o2oLA6mYfkxQ4V
GRu534HnmC9SEe42vFpQtdHFHmrf2Rcr/ax23F7zTJWHs2DanGkLBPlFgUoHvPQ3D7TIj+Cq8d0M
pPzpYcrFVM00zS1MYBsx6ZBjPZbGHKRubypOGHC+aT3fsj1HBX3K2KtQguItNm2LF4VBBQa21//b
tJGy8y/pn1d4b267IeuuqpihMYXT/WhV0b7G5AnxAyUV08TgVVTROUH+i6vxIVwc3OEu2LtkxaN+
PsgFxWW1/3yWoeGbYXAPYLqUEglkfQ3ueKDieUQ5ULHGcvPP/XS7jZ8RGnhG6sVopoOTClkbfqe2
I8nGdwU6IfYK5K2MOBPIOiOGnM0m+svZlknJOiORG5bYSbCxAHv4JOykCN6T3nfTrB+kgLZRKQl8
qW0eCrP3gqRlQC4Uh+WDfZ+dm7iuwMoOHckJtM1YI/r1YU+94Ecv8Nc60pHgNhME6y7aGr7SOmlZ
8CcxIoI+3ObBEm6nlVBg2vG7+MZ21FyhGslFBmYYcXjT/ubiPMgP88nRA6V4CyT5Aj5zgoIhCiCK
cM48objaVc1krQtoPTknyPb5s1xJTjofGoQrkTbjAT5mTUtfaH79rDyIRDmpz8f/bkcmDyKpTgcr
k8GZ2KQjWr189wj717QcdMD0pVki/QykUypUINqwMPDbogoujoV0Bj+10GvfNPycd1MTkED5JqGh
/Yw1ejJgHhOcABkuw9TcqDQWMlK3cF1A7KN5LX6CvrgP3Hn3jI+3JZRLx8Feznqx+wJ7sfGHNjCa
rcCaAux63DzqFbwrpPXBcTGucHoMKBPjaEW1466Q48G36cCArTLrlqX1lSraELPDPyqPRB4CsYe8
CrS2XSkrTD0KzufLOjv9VXsEKONnz5nudr2XC92OH4MsCYGoSyJd58gnoeUb8PvbMPB+rXuzD2UA
CkOsK8ilng9XA30vBeen0DzreoO3ekencpG9TIctyg2waUB3ZzbC8HLqHcMkFxdtvAXK5wk6IyFW
CS2t+xvhvocnRkVGH6MfWcFRyA0PUJymqkWE4nCp2cboNX7aWeZJIGb2XaPY/UNS8CmDT5rqKz6v
1FpepkL5+79SIZ5K41H9945jA68t38FXqw77+zbyIlFYLxLy7epus16ifQgMGCZuwnxQj4hQp1Ba
qNrGvVoMQrJSBdaGHLOEpzpXAQ3qTP85X+TLS3xgd0+Ok+M4imu0YwYT87OSdT1GiO7qys33Tmpu
Oo1MtNg8mSyrjXYogNjUEr4WKIw+iktJJBswL7G0PkjyOiB3V2gUnXHplbSgqtHUpROqxr+/Vxb+
BSMSDtuEKvOMnQsHRnPf9uW42q3GStlFBASMjKGjG2KEjcXb4wG+qhB/xJteLxNJBxwixRw5waln
q0SeaRBuA3gWPsGUhTIg57P5Ty6eM/+d/HlIen9cuqrjkMAmitoh2Dk88fqrdHSh3euh9rsi4nJS
rferel0L5z7LVja2pFpW2+cd/qlEFfzDTsDF/DmPExtHVQPHb9ATN63YKzKwUknOOKoX4+2ai78w
4fHEar0QQKD8frnvA5pzU5DP2vTdvBoHt+9gQaN3mjQf1dkBa/v6uteIrelRkdMnftvxFpPwOxAX
FFhegR8UTrFH9d/fbZhqRE6qLUfy4JJWSmtUrwlsKn1d+SY/cqKJ8IL691rA8vKVe2bdKjsrDYrG
Efpg7JPGBWfGnNOZmfyPrLmn1CWdRF00prCW8disCVpGgvRwbSwOhIllquL9aGU9zQamc15nhSAr
k/gWcrjC5L515RcIDppBJIxyKNCje+cGaQWiW4ZqaHW7IaX6ZfNXfOPlG2CJ8mUGDdrF393JSCHu
G71JAMZMU8dTPAI7dVEqztdVHALm65IDzyWqi1pIePdFyZAAu8nhLim1fw/iszjoQhMUjxhu1HTH
y7hRBfuQ0A4PYy64xcuzYfkHPa2V0ZPHzI6nNi2oT9eFGV/U09VetnzWFUpPh1KtU/q8/xkzS/xA
e3istTgLaLPrQwrN6f/l7PvMvr9Bmj6j8mLqF5A5/yrMInpwyVTth3kCCqqDl0QMVylIzJSFQ9np
tQx9ozO8jCJuYvPgxphpIynLDd0Zsrgtagw2fazj5b0vhmqsMfR2Shfb273hh/nTM6Lloo5m8NuL
JsUUD2fnS1O1BNOeb/ldSH5F4mZOo/7YqF+JdJl3+ruCb1utFVy/FmYgVeeefmuWrVkhcwqNx2AA
YojUHST7DDBJzmL1hoLcE6WfBcZlJKU6EZSwtlnZME2bm7IxrAod06rO8ejAA6f4Zh4y8FuhJVZ7
lCVzrYFaj3iy4KnePSjZ51VyJuO6Zod2ypENkiJjZag/5jD4nvUuxO4+BsUvQviRZKnjfK5PitEb
aTG3ZeXu5PtS4buh9ILEt96t5JpRsY3I7gUIHD5J2bO5zp3uC1QmHsaQbkdnpSTfEp1RBWdnrx5h
qAY4S/MiU+RaE4seM3//Rfev37tiJ0gj9qFiNSAPTTywUvupVulSleBda5VJgz+HrHFKs2c5uTQM
dG+tJdIpk52Gp33Xv4TGZkrkg0IF8DMJdHIIEnyymGJrR/VPL7b4Th2jl/fQa0rEzOdCWUffqtmW
1b7dQdM2L2z36TH1Mv53J9KBcDuoQ37q1NrFowbmuzbJO7DvJ7iYqhZZ6OOwtTm5XQYlgWXMr/D9
uH+v19KN7uAcwAg/V0OOBOJeh9oTD/QiGFpSI9LWBTSSNqslAD7UCbYMypedjLUJwILbNL1oSotl
pgcG272mzCQRxoL0fzBMy8Hxq7hUmYCOpOKMTkfoPdqzujm2YEKvi3uuqRat51dh0ZCPf10wXeKD
KoqzIpHI0uElK3Mn6ulg4XtOSh8UGI6qubMjnXjgdLvhwej8PcSI0W8UzNtEqSP+hjzzfIXkmYsA
0kw2HIfEh5r0hjdS0VhfSThhwbOpHgFNkxnYDrYwBO0+qMxkW27Ssw+MHQRIk44dmIddBdguUb1E
zViu+rFYhfKBx6d9eJyit8DdsfTJiZE1I689ZHCVcnsVk+ROuqOAUv6Waj9OvK+sCwaO3hxIQ8UC
WBsYKSUaB4J9oK/B/VRQaAGooUnx+Rha7jA7jbQedSoHacs4Wp0vIm2xyxWEqaA8eOdpybeGTZtD
KB9riGyegh0JWhnNf73fodfp4ia0XSaM95SgWIQi8ZmZZ0+katkkkjMOMnf5BGoGLNnQl+GqUPfm
L1dsaCRylresv1k2xL/MYszy3dqINsrRrcb059G3xUmn6Zx1xz0NvVuKHhFPebLOEQ6cGW5/4Nha
K+gz+6cwWJKFbBRzzrex6OcRlW0uUVsujBAdQhZhzE4JZ5ZvCOWodpgnaI+fa/4UokHjHJia2jG7
47vZw8MXLNr3ClmzZDEj/Y2s1I/nuzUfdFFeiHT2Sn+Hi+JWRpE2QUU7pBjc+CwMKUf1S6TtjSKF
3v5dFp95uYxn0ffQn+3oLrw+CM1Z/ZXNfgsU+GF+j3Amln/MqlAEPaXUCOPBTMEdxDCToTtKm6gc
/D7teamzhMmOXvc8tao9JUHUBrb3OI1N9ZBrg60dMaLSN9kn5neSwa2BmEUI8MSGDMMM9t65eL5i
4xBigt193jg7RqgV1hAGPNofPhsU54deXUiWXXM0OlLkzJCwv3zKVuy/6lsBFEGlaLuBSr3MlK07
Wlrxvb5/kDr7VofVWwM1ueX7XlGWIZ5Pf2RFPXITkQIcMMKSnhm6Q41x7FpKVoiEfHEw59fH7W2A
Amjqm/g+cFDnJoU7PMUAxVqgAC4pydPk1ou/wB7zfRh2+G3TPdxLTTj9RghLva8Winr7x8by8QwT
g5Nl1ixkSOJz8zdnOVmw52lqVAXvEKhOiEMP7Xdfc/DZT0Z1q2G8GopFhbYabVib0BVw3MDPwY6P
WXAN+57ifpV4xRw3n0lvPtAdRfIGbIFVCiR7dxVjUDAy4MdSYvpDVx2IqY9DZ6dJKou7Yna3/9eY
jKfrjH3pyaFMuXM5aLbMm9L4S9gpKrh/cBdlyymVz8wZbfIQ/vNTJvgyYVW7TYkV/uMYpJHh2iV4
ENRnrRAYR835M8221NgbTCZiOKpcEdHIDMwbS4RRV/Yg/6T67AFJMz5YbsyT5RHPrS9A+jvfqz9v
0A73QEJXZxmKSSXwQfS1M8KEnWf2TYUwqoMPA38vf2Zow3TnXshBPITQUUZT2royHe+HjgYew1Cw
X4BiH96kgeW9GFwxCCEt8dAWHY/Zv7J62tzCZ+e8HATu8nvjBqKsuSf+p0XZXTDnUMlaN5WXRV1J
X+WFgPqYizm5OOnP9DjuxhQhnhZMn5i6pxoHAZgwm/4zQbziEDjzDbvz1g63Y+3yjlpjZ3guS7DZ
eFMYoLlScdsOpLtFVnpJfjL2LE4L4Os9I5Go8n8abemdanoR2nVqL2fnCUsCjM5RRY8DC0Bx5kx1
jsJ+n9TBDxvYzxKi+i4yWhwXj+WYJvRenMS7kQ+F7+rhp3yLWHzyFkqk4c//ma0/4nLp3k9C1HaI
R+7CAjG8/yKRRRo3xj10kH2SGWMu0HzusiGmayxaDhyet+F3J5n/pjcM0b7/iyMO/DcKFqBZ2X0k
6CsYJvsMUIy3xNeGleVurSYa09kdlj0OMg2FwzBoY06wOWjpdvnxlKZSdS1VvdP0VmrNIV79RdJt
lJ38kvzRU4erfYsoxpt8NzW9r0tF1aF5OQVTvcAnbiwOodJpP+HCmpYi5e7L3sJCkhTyDI7x0gHJ
ioDCDzdVvJQfDhZUaYYgkYw3hsizCtvy4M8gYlJCjB5TvxY2ZDbD45Q8eJgPf6JIViwztLTeYxFr
txGKYiepaXas3+eC7KVuEVl9wCnh+maD30SfEtsJ8nRsbxBq8XyLMb4ZIoQBxstpXkJL2sK20xTu
sIJV4VNcR0WyvHzPKhQZYXWt/kAyFign+m5/IX5Y0/1wrfRWGuBiA91nZPGxI+xaTXp5Fd6VrGcB
q9j2sGdw4b4SC45VdN7TNqzDlLirPBxy5/4CpSBbelfBWhPsWPCB0fEj7ttkOboc4rExGJJ7kkWX
k9I2pjsEAE5ez/760oP6LoLTHEGYvtpSrMqJkbAOKMHo35AyelOH8mQYJc9Ngj1Rs0rN7MfyvokJ
hlxGe19tOFaII/lb5gnWwsDEs1EheRjrzRtOrO1BW0JN2mv8Q+89WidjG/b4rw5KQYZMC50dAwfZ
Bw1u9EJ4okjF7DHozY4B31mbamgSJlaRY9RPjPC1gGiq24OnOVxXUW2CIfoUHgpiSFwko4n61k1S
8QIB3utMILB8HFeY6t9d3kX1OAwLkpbKQ3N1B7Qh5PXxi0knnrSIFkRclWIq1+9QE2es1++jO6/V
gA6ioFNZnpiwjUlhJcBocOYjMWZUk88uO4AItr/V8K8CvqyE6kedUHZL7S5yuaLT332BfqYAvfv/
zoQAEEDa0xia8fUycS23FDWZCZoVlvQxZAlJ8GvP2afTTIIT24/ET0uRwLtiX5jLDJtZZVDnFDZ9
Do3TI3YQnjG6tQtPcbcNEDBBAruwwaqpOQNQ16UuFSEh/NQCsz1t6qV58ChoyYRPsZp8QDVVANly
IeRkTJDyGXTT8gbwEI+OvZ/8r13REGWZk+CJ+FBFfRemuACQgLSLpbnHSG7HLeP+UiWJWZzbStYQ
vgLszCliNctet47cSZXcl3c8HCnaY5K9Tn6t8x/BO0/ereEh4LudXwyhblRz9ieysx6z5x2i9Md2
xh+CoK2j3DQmXUqoce36GdZym4MMj+eQBVDOdGoDj6Nc/yQy0aGPQIoegaHa8eu3CMKVY+LQbt3x
ahMe8Q662eYl4DGHrl75Zh8rbT4BMJRlL/L8iaogaxyVKNcEWMa/gFIV+G5GNepRIsyUp1GYY1kC
nzCEgQyloi3QSHTX6f/ZnFkfKJkkGg5o4iTbV8Y2fusoqh4Asyjj0imXNyPEhhxwjUbP4Efyl8BE
fJNlcl51tvwde9t/6bezeEJo3tw3SrUHYdcHCyx9QlsW+OBvX5u/xMw+Ku/tYaDKaHSH8sljA/Ic
69LcXz9fVCVsT3x47s+f3TiTmpA6Wfw1h1UfyKyimcPS9s+iGh059+qDq1Zrsag5Sy+3fDXXyGPZ
4taeOIvtlkFPdzVvhQjIysmm5uiw58ot3sNuPAwisCYyduomRi7BZ+PKJWsaqA6exR4KKC6nPdN6
xhBDgZqZ+4M0SWXZ7aHKLqyTvPto5MvKZAG89+ORnIp8XgLmKaigCVBw1z/0/ZyqjV+YY7scuYcD
8qzkggiwtCrdVULdc79v9lTiYSptC6VQX1aUpAWJ6o9Q3d/RCPucvpFhPuL8+phlI5pWDr/IGfv9
4UgGtys5jb+k+o9+1Djcm7Nio6Swz/CFJxTYgTTivEXd2RI1F3gYaKFzuEnnWecHHqKJ46BbVLr+
PglcE10Z7yifKjNg4ECEgVx7ftWUh25B07Jc2niu7ODh5WtRt85h2OMMzeCkLOL4P6w4hVHxUDbl
IZxdCJwJRppQNpG75kxH2/Wgvf8umgLwxRZHWPYnC2UVXkHjntdLPq8r/6Ep/X2hYT8OkMI+WS7k
vv/7RejDKgWiLGPx0wR05M6h4NSJUD0ODtYgtPtNsLrF5MYjlR7Ft11wbxSuJuG2OYaV/GFnr+fm
hCKa++uycy04ifOz5YSY8Pejk0YdCeppvrh33BVlB9jSE5bnQlMW3AcLTlnopsxyuMW5sXb1DMbz
a0VPaSvRSGphg1Xc2g2ynrp/Gw+p8LuMO8Kfm8ObNCSar1mrGT5AWC1z2uuSnPQ1EKrcT2113CHr
j2aj5cMLF2WVJvQt/7AaRHCVLau08ot5sRWzaRSxaHAFVyvVQABqe9y7kjCDwe/3KRpPui43t57O
y+4O3BEAzCF5t+sd6M8dSBU/bO3ozZa6KODi3UO5ksSUDWJU3C1hso/f179etar9k/qJKE0biqfs
MNtEaXwig3kOTOEUGCW2IcqUX0z7jiuI8yeRWiGgGdq0lnNg4fjLbBTo1epnIpSZU5uetnd0c3xf
1GKnGs+DkNm/PGytG2wyd8I3tHQD/0yn4XbAFEYWMywUyZMEGee/heBLmImrJEKuV+LYREYUo0sW
9oFwaHhAVq4cmymVljQnuFOXCUWLFSEZq4lJVgt27bzdWnhbJ3XVFZT+1mYuZQvPlxgNn1zsWV+e
eKEl9gH0nkEr02dzEzZAopUBv7puHi6pVgHQthF2rGreJ1y1ZTSATB82XonL+U4l5eiGhyv+YV0R
L2rt6iMqZ7KjrYxe/88JswGSqWpEsT9YNSZ7EHTNcEOLUZ1JdBml08t6R9M+AAfw/4BhEPQoNdj4
4hlGtnaEA9e2y0AMhSBjqIx5jxV0m5ZmbDiB8pqHQfoaIMi+zo/CR04CNhO5V4luJ3wzm4wQ
`protect end_protected

