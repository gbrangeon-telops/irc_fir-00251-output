

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
WrSZEf64fUAl1kVl9HWWVm9JOgHMmzn0fv0uusEaRSoZ0YHKAX+sj6D4gL2WXWrV9+rdMofvPwNs
9A6zs8psHA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
R/iTmfCVAo0uuZTRynJ9b5Z2gujQ7+Xxv1u+96JME6mwR6F6/MPV4ayotodCx+xcD+9l4Ktib8Ml
C05jFwQ5vFi+09RjQvyvxQAR5CtE87QE5Bg2A3Gt5QmE+m7ZfJiQZgi5YQHL3kAHS0jfaofTkZIU
6VFVSW/fcrod0Swq7VE=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
RAfB7dvLyt2uCWNWspMeHiLYPG4TlOk+8Dptz+NhWH6nMzYrNkf7IWIjXk3hEVf7lwT/X64pynoh
QoCCtl9AW1iC77VMTIu5MgFRizuZMUfXZ0crSPULV2aGonx9nQ5JKx8TiRv5BTWxeAsuh1lT/5p6
2v08ZCt1Nwa8GPmEeFnTZsTB1B0jFzZQMa3GGdV0nEcSjDo4bLIkw9sMEBW2OdUuvE5yIHF6Z7++
/wzulmNKOqQpmeHrq3r1VKkMUHNzsDpLkGo5HMiTmEUJr/s3uq2EhCIq1agWSVbcEjS5uDaYcwdG
D4cRvgOxtT5sxpWA4fivRX7vvCyun+C2e4pYew==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
MsyF52v9pEo5RpJJtfhlgAJQ/9a172C6pJMP5S/aXQMuRuv2+JV5wCeynUZSXHj38Ger421EXuQd
EmO2OIKWiz2pShaEh/NwF+InGDF0QzD16vAgn24LAOYAOX1lcCquf4w2rs7e+0dn2PO/GYRn4rxl
E65F1qdRiZlUeVoRHdk=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
klspBE6zapxwDIEksFW+V3vEj3afpsQxyK1CWGpsw53FDriMhZB4hONIr9yRSN9nitmQ+6cnlGM3
S4Cxnkb334zdXXX5YoppEYaAdCcB5nDsYhSpn4PyPhd2ANmiSIXxEjiEJ9MDJlVIobzrtkNgFEWA
QkqC/Eky3QLBOqPuDJIgkf5UFynGEkI3eWzGSyuNAHTTYXfoLlYBh8nelaKS5vgYh7jpllyo5l6k
hn08k3sWZKuN1S8dwb88eFGM6hwg1UoX7pTnUY5yGPZZS0JEiN6WVWRmh72r5l3yyFZOFNcvByJJ
z349Odlh9AHKI6joGGP9sLtbKDrZfmu9y/SSsA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 22384)
`protect data_block
+PXvzHBx4GkS8RtSnr7JxA6IhWp4SLBChT1G+Pel2oI9CO5+4dv8D1TZPZd3Bo8lZuriDEVvjBLG
EM6NGkND8y/lgH+JA8+9ufcRLHVqW/gGO6cSe0oZaoYXwoCdKkxcu8wLCA3+Vc0EX8Rp4ECt56KD
qF7UEDpi4ujQTOLYHPizGrrV4aUJ+Pqo3p9fkvIXyimhin1kxDtqlvtyi8Mn22Or5+R1tqjkpH9O
O3uhOG3QrveHVPT6TjdSfUZbP5pbmHyvAWMIS5tbfczRppVLlF+zNJfsotJ53bpk5AYzcY8DesMa
7evhdS/8pVejSvrzF1lhRF2i3gXayzWDjRJDeI4JvyBYvez6VvRiwV8IAlsKj6Wqlwk5xGnwR4VH
t0w8lQKinUgr79iCF57CjdpncQIOXiBXXkwdmqgMyeEe36mlbNChUeKponUY0y1+UkvyQ7P/FI/P
9vpcOrM5EyQP+jB9yBZiihid3AW8hw0Bjj557bleFOr8aIu3cu6CXRHFb7k7LQYsnuoveM9qFQOW
RfKwmpBK+on+4zdumYdG5MiF837u6CvRdzxafztYJVsLInrzBZnTfyldUanuDRRGYmFdzVJcPqb8
wQa2o6CE4h0PWYSQH34zvYD1oPD5EOHmtqf08yTdx0ixdoWembwq1VwB3q18cZ3BIRTPB4k9jUr+
rX5ud+7hCuqxkkGSSc8CWPjXaphKCnvklpSAuu6asGf65DOEuyIqZ4Mbym2f4NCof8fjSa5F4etl
rbOPdj0wpPS6ePeMJJTvvjfzTBYtUB90S4itcR4tC4h3iZ5EoFZ1SMb6CC9HJwq+r8ALv/2Fg5ey
fjHOAsM0RD0Y1LS9kmcpxWbQV6pQdT29I5f3pLy4/G2swpamT0jghjOWwQY5zBTDydt/ofk/R0hI
5u1PP1bfcQPZT6AKxRNfPCSo0I1gvFFWDlui8Lr1ctE0SFjsIahJ/MH/KD9COW5BWNJDOeiLP2Uj
PLfbHuAgn3o5dL3nq0XyhslIdTjiAnliKvHWaXACQ5QGMZQj9Or8Q5yWsW+o15tj2T7t+FSZzkF8
NxA2nTbVSQzihocZ1I9lBwlEvCY925hvlLxiqCFSMJZs1QlaR7xr56mRyvZfQ4BPuC609xZe6m3F
bG1i9eYsm2drbAagdlgpl6n7JXV8b9kGKYcoZM5GTMbOzsR09t3LyjMOjygEUZDCm2jnae/ZP13b
S/TEReVuJn9Vm2zXbvGfxms/L3OPHdZb3L9hxfeonHUEMdtE1mwQHRQqxJ8/T7pwroWGldH1husU
C8q4NVh/H/dfmRPF2f59RWrjdR8Yise5ua3I9hqI8CewSuBfIIy8u9XHzSuUZYuWljyMT4PmaZce
DFe+a2HbkENmJGsuvMLT+UGDFdZ3db58MJZdl0D0KH2Qs5I835ISJpNTaq0ABrhRhypGrhoMYbJK
NPvWdeUg1gs0F8SiVuC953+PCOJ34QBaCLYlu7jrHpMW28NMw1Dph4EWtBoTVe5/W3Z09xvmI7sl
PH5FVS4/1MGRUfRw5xLS3qxiQVczzVkCebI5CKSd1xWIxcHvN698MZYwYXJillccrFIwiZVW3dkt
5ObsHwfJX/+0phqjISBM+Jh4d1dnkpPDk4GMlPj5EYR1ecZI7LtXlzlyAGqLAU+GrL2xTcjloOy5
7TlJE0KobZyYnq+Pu9OLmzyQ9pNfdkBeLSE31HDjl94wdqAv45T8N4JTUl1LEaShLVJK+4m7ouvE
zRtkaAEWJac1hXMWiN2+c2TbtWrpX/GjBaB22wbh2dkwyHrXd01gDQdj4m8xhnCsNgm+icv/Vu4L
NeY0RAxXSXpxTEDdjjyLXgbklNUkeb9VuEI1KRpuRfjNsu6k64PGzDPVO2bXLKZQiGIbd0C91eAH
cnXWYhW1HBiJ6LFhKBpGNkWnBQi0r0P8dqFcL/ZlB6cobnoF17dcpoBwZOrfNf4aZSrcTnnmc8wm
xVWzh16ZnZAKI8O02zYR5sZ5cL+cF73VdYxnqWA1vK6honBc7/uW67UPLCTqWmJ16ScIC03+J9hi
c5QLlRLiBsUde83iZXP8lCr0Z/FKZZnHHK+Ieg3dyCSoavsFEGLzno3Ha/nNIs8xvTlMWCJA2aIR
RSJhWlJ81TaTUIusWDd5R2Za4or+YNZPzDDdtq8Tphnn1jElKXLyIdPGooCAKV1aY3ibph7/5MUD
N/5KqRYYGGa6LORFmbC+yMDylb0f/jybhvjnvJ221Irt+RBF4BPxYz0TGkxbvDjzBjGUqiC5h+qz
r7qK8K9eIQpyWehLBfM2SwSxtOOtgoKXr9kwQz5RcUeTMPzenfWLZpfYlpGkyh/CGGFxsn1Md9Jf
7lPG9DbkaT734jKEaIR0YcXi758j7wdEcsp4WGzKniPfqL8byXRsfmxAWAzXcA+xm8NUhpRbJYQn
kpOpI3GGvLpSwpANPVDbyrIaZhGA/2MDJAy5PMOsKAlRq+QrQV5RFEXDIiMeT4SGrZ8vW/CaQNf/
2DJyPbmwy0zzwvLMskbZrVJl0d102G1sorR9b1kNsFRzyEYElkokS05rhzn7wKRRQ3WIq22oESvI
9mLCywTzoXoqWagCKHb+hh2YQt9lqD79nNVaAPlcXMxfSBOr2OS0xkrYmJeHGRj/UpBfj8BY+YQC
s9fEe1e5lm3pBXeJBkUWdJ4a4qi/POVTa6eAbjZoY80Jdbyad381U+1vkHyiA+qPgpV+hI1xTkN1
uy0tGhlKMDFaX7AFHKiJl3z+DTzU2+8VvY/ybD3itJPuTKrDrjxCGhWcTfETbAioR+PD8EHm1i+r
VaS4XV6J/PfLxSYKHNRZ3q12DyMsjwHE71s0T4gf2zNOvKujo+WQkFMZKm68C8yWiYjhGxgqtnkG
Ay1SZWJ292REBMIv4u4h4b9UUZrSln+Ct+RHtNIT1C97Bx2uUyxIIgO2BZF4N7jMVnlmNvqy7NIw
RpLQfx1mq/q8JmMa6vJlHDLv6oN0IW22/zd/WqueexDgHP5zsO/u59lu/5Z2umTKVhx5wgNaBZ2F
LHZMfjFCanKdImLHxzyoiykyL6EVYHIyptDiMErFVDU5P2HK2HFZ+IooayF6Spgo1Yg2Ncgscdqk
nNvsoPZct5fW6k9f14NI73G2rtYVjZ9EVqP7fr7tMNZeF+DB89HlC3P2UytpkX5N3Fn8nIf48/F6
2hSLokVP2KGOgpOa4wX1Qg781mi197mE7QTfLGmaO8pl/TiFNvXP3xyMcUYiAPOyc3zeJre51SiC
FP8m3DEn/HgcnDDq7y6aW9//zU0GQBx1P/dvZ36B3yjbjUs/BrHPoZgao2dR24MS7UPx4p2fLuR9
JUryD8vE2TjCHatWXMSmoPhoNfqZtgyY1iCl1L2TGbo+/8Fy/ybFzOXFIU61TrnK90CIDyA9DHMJ
hFNYJQpTjTufODyeOCI2IntYIkRPme2oilhw+p+3K3Cl8izTlnoFsZ5PMzEKFfX/mQ09oeiHqTwi
9U5yVASTa/w3TiWS6fbI6JQfUaYAkdoL8U38YhEU+pAUh0mSMwbH6n0VxZCXEBy7lv/G4bIzN7J3
A7rMHRVbtfvgLRhXlhkkQiGkROZWGWJOGO2LIwVrUAAVk0K4KyMt8T69Ty2+BeOwpXrsxmew98V7
x5AWs8Pt9WIyUPdlzRKpIDFWo293Bbdeq8mBP8pIFjMcE2vegIs5iKBYo4aeLPCfgSuXu7OZiNd9
rRqQoH0kC6ScXcnw6sRrDM89rylX6F/DliQSD+II8umsLrYhCZnTujm0CRirBwvfQ64FjcOUZK8x
9+mrdU/dOu8LeYMRtukAClqP4ql2BbwP9VCSMSK3sHbfrGGHfIawZ3zzT0Azmy+doLF6ZzmxmBtm
otLxFq6XqD2aRcvXF84qWqWzpCWp3DUNMBlBCsUZ1GcjV9ID15tfH1YnkhMn0cvfhMei0wpEHplg
Z/pNz6TRNxTfpT/fgjYgHadseH139Gz90bQU9huroie94tESPBIzJYrUNYAMkImgtGIOJJTcIuad
spm0VBpwuBtYr4OsJFbHr4j010nUtyZMoffToSx5YVdsZfm9Tg7oDelWG8KCbUjYCz/j2r4XukMk
U/qjPzEMxRhTtShuDhfWM7GbZc0JDWxmUCr/qx89TxGRK4Yvs+6O/KEH4VoDXSRsYeMnBGLYVpwA
NXDxUfiyBQGF+gy+1Exwsj6ZeozZvuvahy6cSn7VfB6t7GXh9wwOuB2kCAa8F/oOSMsfxSuoy79A
IG2ynvWszjTdKB8wfHWA5KWyKZxllBuHCZgu56VFMoF7drEyGrp0gpkTiJMAnrZ5RJHa+HYcLpMW
0UTKNPrP+TXijzJ04T7K8T90nmzFBelSqrDr28kFoxBLKcwXrU0Qy79tfV+ee+7mIq04T4mG+qNw
gpvSdH/yNpgNslIBAzooJcoN2MM34LWdEeJqJP+UVnjyLFsh0egu+s0OCb/ZPKwIL2N7opz3/ZFL
qNSmG0yQHrj1eSEQ4bUsXmiL7EldK/RGmmqIWaRkHYCiYzsOs7sMe41KxSVG60Jx0iHGzf1NnJaY
jwfhIj3yTmfALvyguo5VxpguNKgXr5A4gHoU+ylimgWobhzwCVXLNu249D9o4QF9dXXK4qXsD4nf
I3Xd/Fcvzz0hR7vGGKtW5MsCCnUDqSXN+01taIuUK4zj5qjygfhnDYDW6j1SPPd/t0NXilqSN8aY
FO4qQEhWpVi29kkTenGuxzbsHZYTF4Ste9fVEe/sGNncmeHyFKKOmrvYMqVmFV7D3uGjkIyvxRM7
Ax9wp3Ms6zYCDx0aX5f1D8JhizRrq1jwCyXOlKQ7dMQnuMfjYKfdk0K2RS/wNfR+VYmipWhC1HLb
04RmaZfxiTaQR/A4jE3UvsUm479SjMlpa97nXTjxYvd/G9zh0HXqO6Fy1Vbu7y+25ET/FauzEQqv
CVQHvAg5pBJg1fZRuf2Pn6x6QH1K+d1F3oCLiVFM3XTBcY/rR29U10zSsR1JJjGYFWAcYjb6dia6
meCZ4ZSWCxZe7Kwsj1fLoB+jNJrPq0AWimXLJ3/+9nUoTC1bnAaHytlT+7O2J1VeLmCvxMjZkhGk
/tVutAyB181kNZs3n0DUwskq0dkxzy/wVFNAKez+YISLi+kBunpDyH2ailZMrs16RMfTAVDBRP7A
wdV/Qs4IpNEmwR7OkOMB+/wXYfzokFLQzkCiQkaBGJ8x6M4VZDL3AKa+RxkTucDg+CXM/LTiOpPA
scLh9LFbbxtFhFapVB9mHpyDXz2yOM3X5WJb9fO871UGONb0cDr5DrpYdWjBrfINVtooqwhahU6T
R3oGkXsq0fEzAlT7elrF9TJsR0ZG1cI1aXWKjAwoIVt7ou9sSS0WtvG6dlOHvnZU+DJR3za21zM2
ad7n1h1wH0W0OPHzxR+5enIslY59GTp+Yxf0z0lhyRkzCbD9uYzIFrETuIcOII4TX69aoxIKe7KO
2ULwAva7qUjULFqj/yxhoksBl27/JzoCG4ZGrrQDWnlvjJqjD+VrD8knpf8BU6B2Kjy/8Ndtl5ga
9SxU73IEwl6anckiQaWz+bZQ43I8a3vmxqbiU7N7qZSgk7kQ4cJyfbcnWreSwhNX7VjiAhxHNSI4
aiNdamtY4fFsGse0uGZEtvNOb/6spaSQEJGJ6TmIpxqoD8yDeBsoNqjCUr8/eaao+VvdQLJFcjbz
HEnyyAse+5S3o1FPaVocDE/UQWTlU9Fj6wE+4haaInrULT8RCN61gPpKMxHo7EMFD0NlIJKpK0+S
S8Ij3eLQAW4Me/8lnS67St+9jCzw7M2nmiHjIRAALKq+IIMXQAZhiLL3zohwA8HTVDexeqqYgofj
pBh6lmBrAmPnOQFdeO1ZnmzzJTHrmCJZw4+Mj8/JJqri1xqxk+zUuaxduJPojCuRM7r6Cdtt9MRz
lgK2RvNHI9V+YS7JarlUP9Lf8VTy51ZG2L/vS9GiQg1WMYtFwZ+PS+jAEajcBqi1ANsToocM8Ai+
CLtRLcS1B33ah6iI3bTyFSBou9OK7E0Q4IRhopNgG+FmZfZJzeotD6OmJzJSMIHo9kie4YbU/Q3Q
2P2EvayhNb6rJhbqwTy9tLhAgDQWqAc6ETo2lemTSL/2+HfhrX+DINIAQvS+JlKPnnzjgf6aV996
WUJUYSz9wimhPZLD3o+d+8oCPmwIqMLF9YcVQgteezIK1PtPQGJmzAM71U8eHqI0wh8PZ1uMruGA
v/vnnPghkEKnh4coihRYQ+sc+HiU7sW2nYAceXHX2dDHVorQwGHOFq9rQrDw+3eK06JB8ZoGBxYw
QOZAY6GwLhqaZPh6AFCwBsOzAtt1Kc3oG0EDJzSPTvjTCiRRcMhJnfApiOr1ddl3zYgylm05MoHb
bTyYMZt7HMGJUoWGnjuX1LjHqq4Phv+213CXbEVfIoidSRKAqDCjXPuhjc4AKIRSv4WdB5uzNIyZ
2NNDxCCZHnLmSS3rVDtv0Zpfsf3qpa+SI4NbkBqrze7JtbfMBvSUbx1RjUW/5+czk2v5xaB2pT6a
X8BUsuTs1VSbPR435+UKLGCPpDbDa32z9n4imedwyXwkBeAnHXaax5xYWXtEh3pHJJ3AuttCn3eM
Drae9uo+tp30LTpYAxqAxt6apx8LLShydpUyOf+eiZOO8IQnlp3b2uSgOiba5+FLBA54dyLLiycH
Y0B2NYNyeOKfaxcrSv0oE1SaWTlS2yjI+ThAHdDuEfKZRAwrhH2EJkAD3nuhjUqgpXlEJ17gZGxc
64GlqVvqpmANln6yX4diky6McwNCZo4hKd+b23HXkm+lu69x+ZbZBCb/fF8cUha79SDAzkvabLML
gXsU375e6CDxnPiFsY34onuOY+ltB0k+EzOVS+7k8cDpl6UrK5VF05/Eb9MUVuzizdTwA13jR3tf
YEoCzMwDj2nGdYnoLOzhdbMjwtjqoOxLYh6DqCOIbJvgg5eFkR4/Ix0llr0TBD1MypRtyivj/Au5
NTqP64/09ldM3vQ2bSJUcFzJRDKxq6wPQpzyw4wsspQYpH0yGlY6Kx6XsI7eYsHZZ93UtmQrFMV7
GhxFmUFo0J+HWlftO9vZMA0h7zWO0VrkduPuT4I/Q3DzJnd351DnwfmQa8MJB14NnFd6qzJOv3tA
FhOEiaBd56rswBqhmo2S66OoZDIRafKGP6TpbgNoUnI5hSVBKKR7A7sXFHaPs0HKBBFehmO4P2mr
emphsvaGUneIZNyoFIyWVQ6XTYNU0LYOo8KPSsmBYlBsBqCXQHpG2Q9W/GGhHIMSZrBIYuyfa5DK
PthKNbvdMBR92KGQZAfe2zHDdLCtVDt4Ii77arNzb9DQeuh1FEHYoGA0HyhsV/yEgxOPJYDvMAW1
v9IspK4WHPW/XC+kkf8VRWoZUsH6sDHvpaLxWmWbyiHt/LwkcNmyjgglhTUC9WJd0LgKKiExOFMt
+WLPMsQyIYxwOONMT+0qJA8QY/6RxX2VXhsntoGIJmTxUS6X0IGMk9zq+q51W2rU3Zm+2SblkRCo
mXOKYBbbU2hz8K594ty7HcZXiqQQ60C7XrIYs2nK5LeCrn4Y3mrJnB1q2Iwa7xE5I5WcOCwxoCdE
di3WAhlbqPT/oh2cwuPMUp1smkmAVqvsnjaFa+OmkFxlj83GnaER/q55wbgUf8Jxv154qc+iOl5Y
4uFR72CIEIGkZ9JL2jLWUYfG03/GXH/LIyUovzFEAyC9kn+xp2Oo0KCgD9TB9eiEZhw/lqKIdbTp
GzKg4dAP2ViUcIwGT0qHVW1uM9JrdNDaETtT19L06vejvARVTbqy3iLUCUbkPyYIfl3DHe89/SvK
SThKGI/CUVIbIqhoUw3Z3WnC9bCh6t9SEIPAxYVFLx+bfvrBt8NQVyRqB4fkwFIEmPPJTwOo6a8I
9PEiTeBTEXIXSnFV206Ep5A8Dak2HDugpgcETfgmdPJXuuRE5UkM8hAvtudV75gfZUwJAFchMfh3
68kpWBpeczO3a8gC6qRaRlhHFqxwE66seNRF5UEhRgS2Onw9CH2xumnhz3LR9LTCK3ihp4sU6lZ5
jzUKIFH7mMdij4EbEOFvyC2NeSOtkbnJpDvGi99PblX3m092OKFBDSBSOuPlDxQsi2oN4cfzmUCg
H9ZlebqO62gAPQwfVKsb0QAoDzMRL5u+hvV3MJGtLZix0nPhB3apVcVmcvCMtbDDzGxFzc2Hcr4U
zAmqov3ddkpj2wFZU6ABQmhL8WhlHKYXhowdqGw8VshE6yhgQN8tfMrHXQ3RuywU1GS/xHAA4yo7
RGhfByqjvfdKLGEFlDp0E2ixNI+kbbZYiZythrJUXa2eRril5qnUzwmuMngmzpAx7GZ0w1TguzFk
lrVE3537M6lC/olAV1hiGEYrKwILSGJK6T3gn4v34VQkhQXcVLDgzpZJyBbd0EWY01LJmKEy/0sY
0ELZgdAXQaV6fBTyj8IH7RZrm8/7EOfjPtDRNKBejjGLTBaXV/cJ+keuW/1WBSFA3fz16oxsJxO+
3TAXc+vCk+epdxnvSd3Hx32JAdYUUypN7IYJkeN9uhRZ4qvgTlDQ+X/7dj4inCP9zGXeya3e50GI
Y5VayRZlBz21xYQ2M5alRIymtJ4QlODf0m8f2Ab+YaF67MM0mJRdS0Iom7lSjGt2SGXRGWg0dSqK
MqVv1DZIj72YLAH19QBJJHsc5TcmqmE3XioPjMR0fGypEhXtUFH//4VQvRxSjnQNj0SXEvein8aI
v79nDRCW1JisZzuoTMHWeAYwr4xL01R7Y8zUxDcou00UPLELV/irXtmzurXcpPszJwZdg0kt+GXv
8OUxIn+XMvTQBIJNzV6bdJALgLbSKP8xZHzVgH4jFN5g4EcfL2lzqSdGz62IxS47c/+EHXXHJJvo
xQP6S2BRHnN/kDQ4lhbspaJOIIGAffagFIlzs22WIxEcx0ZVHbd+AhDQfHjXShfaecwVuSV0yVz2
7qhzkvIcgpxk6w0xs+d6+/8hDpOOMUjr1Wd2TTYTCKVpiptoF0XtBrspdGwORJJtQNC/cd/m4+hP
7Acs+Ikf9I7HzHxv1qObSNZaqgZbnPgIxqcVTkLs/hjV1n87woNCpPeWe8A5vw0F4Q38MgGUIx+t
IsyIJhWrX2A0Mv5vVlg/j1btT0Q4EY7qq5n/uoKb6cv9k20FPS0WuW+BkHQtR42J0Rz9UB3X17wk
ljvMFzQN4LwVwmGkN2u3HQck1gHVhJ2PenEQOZFCsdjLUfylXXYs1pyxdMamZ4HTRKRG40Z9mmFV
03BkQhMbsX8+XLIHKvuFjw97BnNptkGA8AkPU6fazzEfCt3IV4CqtQe6FmJJCJesXkhOCPdfyhTs
+IANlEP0giDdxKCOiO7GBzpnj5dG71OITeHPFRJ3pKGoHWhHpXaun+HYoRlxdEcx+m34d4yxuuAu
QKf0eGu4bVa9f10HKDw9ZhjGMZk+LATtmykAlkWEwNnSEHhhuNXemziVeTmS2K5bieOf6kZWA0Zg
d/10pLUYo2OqyU8VxBQ9gOOHwzEGBJO2+tih25BsTwHVHlOQuvTwMs9QBL38KNPNByLQzBBblo8P
8vrkb8w1pO03VXlt7mXcFsMMsKz8kVQsMmLOk7XOoLfleM8yDCCq1IRI80kQUiIcaLo7TivAxEXl
100mZnS2uG4DU7Xf7v03iSPg0Ny4o5mtiiIEzZq69GDLatlWIY49Mg5JBZ8cKmaJoGvEQhqEIdkp
ej9pua2V9GGBhydkMCNp70FWAuj965h0qzuDc7B+JidYWZiHMZRDbOZ7TkBvQfm4/kKQd3QO+GZB
Esf3JGAZj64lpx55P+JUFsnW06TbrlOsbtU+ci/+iaerDtylsNQ4nDepMPn089EBvo9mLmeiHYn3
Axq6l5DYVPE0nb2gtiC0Eq+gcdugSq7IU7luAx3divOMh/+j4UN2ZyG/2Uyw4B9YU862CtYvlJl0
+CyR1tb9a6i8KMqgtrfhqphNAx0qDkUx7osJLR/aPywRXUv89YnYcGZVRQ5jfsA6QdJTC3Z7o8Lm
FVL5LIeBFrkFiM8Y2V1kol9sgKjlmJqHYWBzKbrr4s4g9pfnBlKtBtQ8qFIqA9FryIGAQPjQtJ6A
4jYgzfPwdjNWoz4wDca9H0sMYXzcN/oON9734WzOLBI4k3leqLdGwzY0/d3G8i3AzC3E/mlTTCWD
2SIi/VauWToZULi4Axl/xZHS+O1Cky9oCMoKm4CtATrZRr0mOl/04UT7U9WlaeRm6YbEIAtJgmj8
4GN9YEgKTW8XAcw567ep8J+eadPnmbAO7lT4k79TjRNegNQPAI9l6MyhMybqFw2M+JMUEhXCTrXK
EGp/njakXOW9yO6CgFNskOXryksWajodJuEKxzO4y7j5z7gAkreSHSFWWwVBOjUKt5ApHF+s1f5y
aJ61m7Tv9AgJOkVMr57PctS2OOS9Fup+WnnXDz96zfmrHpaZ3+dZZRqNYXJENvEFqMbHjDGYfvs8
99CTrjl38qRC7jsNPfH67U/APo+T7O+TiFF84ZXTZChuly5lf363kj2rEpxpqUzCSH7NWOJjV1bM
/GFLt72/J1BgLEQr1eRqF8069u+REDzec2vf+dZnxxrmbxc6GAUEmjezpY2ENqN49NnD+tRdz5F2
X3nBf3WonUm528lp0h9KYgEHuIFlVDVwRGiSAgqoqbu4o8c0HJIByqRiu4Wzq6afiHUZho627aiX
sWh/eQURWaY1NvWqwGOHY8nKOhNaNekS/JLJMm5KwJoaIGMbe1nZz63RxPfE00/bmMcbiVp7P7HC
nxACCCDAXd5oAsSLC/v1TUgeL1awesjI2BFFvd9KHGKA2ohhrIBvQDlWf5erlmcPwcBXT97dDlFZ
RYIjcfU9xI4gA95BHYx/lsWaYIZjumPd10ludY1ydTJJvwyzR3kylk+uHuidP+L0ilq64rcRVLdR
OGGU+93GjweJvhqsHjj7qNS0ATbUEWz85iYNh9BuxPdwZuGzZYCSj7ZRy+fJI+KWOGPCXSa4pp1M
CG5i/5WquQ1zec4WUOVWjf2QNA3+3vB6tjOmfVZ1CvcsqI7hWsZNR72bncCi9oJRmV5s/GA0x95D
Bum2kXVB5ZjMSHwbrGswfau4F5K40YZL+Wm95e78enXIA5y3byKxfkIwenV/LdFAU+q+1SGpwEPa
LRcHQ7HTzF55KJXuLQzPZYly1YO0K9FM6WM3NpcukBCyeNCJ7/hcU/K5wZvhiJOAq982CiP+JkgX
2BRWK89+G/+QAlR1kPpFKk1bQFOqDfIjtOOK16XF7WbD0SJbYsFMkayN2xENcpEqRU93cLYrymg4
tqJSdavFc9ES9eEeluSkpwVi+ronl2N43EaeGsnaCYtT+LjRVZWKol9xPI+FTA22xsaB43lDGJ7s
4rywD4gqi51rjTnnGrP1S6HE/DZTmNEEISP914/VfIGra6OGYhmjqXE9Py287NXcT08vOwTyMWid
4fFpw+yLaJrQZI3/L7XQuA9dhsiBGAeE89WrCbbsnC/JoKkbiu+/5atIi2mn2fPCx4I/5fCPfNSv
EW6h0S//Y6+n98mxaUKA8RMh5EzvRjIRYyy/pD9iX/3tPVwkUDbkdM4t58lwmv4eWx2ec0/Z81R7
puBFpPZcOh7ek4bSWC76DGNKBcSR033F2Ug+al1fLCU79DdoVNkkeDgGPEsYx36w8wIgHXcNs7bE
NPLzccxJE9ejPd/o/TMwpXJap/dI5M+GrGmrlqZhVe2d0pTZs2OS8cwO0RdQLaJxpVLSio7kiRDh
jhaHd+OI1iPHC7F9QeJ0CcVJe40bVhWp8CzJF92D1gdteGpquXPYw4o3ovMlQUTAC5+Za0s9Rv6H
Dm3wmYCqXK2EeQ4WHG05mWRGJ9N9L9ZrjrMnZK+5FuFG9lGbFVUI+/N5hTd2mbMXmu45Gd70m2S5
0+ehW8PKwJSzLRCKMgZ1XZ6Ti4ulvKTHdkZbYc1LqpVvovwzAsiChwBS3ci1uvVnRtyprhiMXsid
yNpeEYUFPm7vE2t8g4akriuJbzp+SKAmWLckRWiwXyMUDrkp/XKSB3xL0icXpVO7JCzQ7CFSjZJ8
89yr/A1Ad7HEAXYsqj2YsPd2HqFz2e0OmFBb33kgZKwcqdMWR1vEhFkIFr94JJOiwY6yxc6DrolY
mRgP894bD3MlqO1TX+xQyejEynx9J6ju6ghVhrEeJIgPT0kQM6CrLoUgEuFR9eq81Wo6PAvcRecS
ZIj0QiJUx3YLgKsF734z7czATmJelrnwGPaoFWaLxOEz/zoHZJO+sGBEhRGphVz9gdzfhpLflnX6
WQyM7n8c7r/iSET9QFDZnpnHkahJnoHAjmhBdlTQHNrpNScJhPa+T9yji79/MxR+Id/Lca9E7S/q
pYMwN7S4vKyy4+RZTu7BTAoOqHXyQu4Z7GdKFxphTWwa7+4dkg963h77U6MNtoQ6wY9xnFA1E4nx
hUBoX6lStrEBP0AvqhiPy6fsaYs41UDhOs7Z15XhMsVpQkaFpRYWPNJhL9dMA6BMANCkglFJ9NGx
6DnPO7oGwROVNOy1tzR8p1CMekv4dzRxtPF83ArIH+FrMMQ36Ahx2SHO62/0GspmsncivTg8c92m
XpBJ0QqmsJg2KpU4sHgKsdoJ0MxygppDn6hJt7FWihDvslGyFzDR6Fb0gKDSVL2jwGpH8xHc0xWN
vePdbnbovsC6J6/mNHSWSJbG+GZE6ggqX67SmTMjf24td/TBex+LLUyd9NzkTGVMV5CylizHTsdd
Vk5mPMX0zQrGD/svRWPHJs4z2u8jC8vtCPQvKLdwimA4n0JPUYZy9Rd5s6eQxDfI1G2H+7swi5c6
0qi9nK/sAkG7s9y4wCB2WJ3LDtkCESbWelLpS65TOSJeR4X+Rq/nsCbF9jQkietJJq4Y+juMe+CM
tEhBOjN/PropaYsSaHJU8QR7+kf/voPIUFKcqfsvyX+slKjVsiJI9GS+iGJuE0CeqBIUeap2MSAt
6C9+fS2VneQ+Ce+bwP7IqOf48YAUOkVqJYn6rSEa7Kk9Jm/nMtA2xEEeDMGPXMW50OjOJPzqvurR
c3tnw6JMn9YDhrKAzUCzL7e3cEppQClsS/UOYc2VwQfSgZBOJbzT3N34waRCx/IN1xe8in+q6LgK
KTNg1l3OB0QBMUhzasatmJUjL6q7ltbdOWil/9LqLEd9TlhJIpMvR0Oc2BHPN4evTjwGrjNwPk7d
exhUGTe+R3gd7aYbfH5u6D8Yf7uTcwLKwiSOdGYytsB59EUzaghWDHDx46PWJLScsbh+NDggMAoP
1ZII5D0t/ZVlj4u1F8/XDwReGXxN7kyk/pv6apYZEuRFSI9OpFBVjpmF2DDHL88N1LRylieqxkUu
ktdAN7pKJBSLKeTZVNy0FViYDFdBl8Ako7A6bsvHpt2Q7kcA9yRgrbqtkMr7RT0dfwlzdAhkgBwm
nrBgpEx4jgDev/qSn7KEOpn+YuKmvK/bkQkElgxRRmmZ2aSeedZvhr9c5eXZ00BBRjKgLJOca/Ie
uhz0sCL9eicd16jLF2tYDY7YuLIOwgkLcMiCDeq4VDz+GOUkj7t5VabC+kf+FwAKFCGA3GunLUSy
I7gxPVzQgqJnIAG/jVzL16cdQ1Xg/cSTMuQGLOsvmbPCBSinAiD3pIxedLRjZCtFdbDvZBzACdeY
ZO3ckdL760hw5tROI2jA/pXOkBGaFt7tNjH4oliRj7Q3WyB6UMbHCb0xuLrggaFMEl1FksvQ6gbb
06bcCmTrAummtDdKWZ8/DGdtSwSqJi/V4l/Zi9hGFRf5Tsae98em4U590t1H4plzIR0QZr9mmAvg
3saiID+ndBnuj6qzCxoGsrvBHNPGlQsQGSSvwT8UrYEQIXMwW/w/I4yjiCkE5bGpccGjwiRTcOvk
2pvZr6a+9gyDBmpuj3gJgKtbMhSTxl/++nwILmsyR0Y8Fp97lKof5wewatRLJyP9mKwCQP+eiOCZ
evwK3+6ldD+1tc8oxYefyio/apatL8iKDSTbPGvH6Kmi6MyhTXPcARdVw4AIqkVXeUqAFrl8L4Qp
BAKsnSQ51ZS0bDSotxURzn5LweRmPcJEltbNsDkITRnc5jJphypNwkVeFaoersJFNdG9k6ZqpVDL
sFfR9ZC65N2HE4GCCraRdkFX7BWZ4UvuklNHRlHC3PRbrj7f8n1pUlonjzTy4zUOr6+1zGJPmIZ4
AkCdTS2KzbDubVQhQQE0JJziIGjcEBZ7I2xz/3d1R94+buv4UVqoytO0jhn4lp1D2n3CLWiH6IrV
3QTl81I/WLp1MDKyIQ4gdEmKJ79MgzDbh0jWA7WGG2KqW2GPLuwV5+CWsmTUns+TlcWer6KiGNKP
TOZyPIMxK+JO5z5u7jbm7fq1gOkVtg5QVnBx7gyE6zsc7KjnSWOULoqu0ARs+VNsQN1ELZz6GK4a
9m8pPkLQjNKCduxT+LCcXwU84A+v9RTzj/+ZHov+x+rC3ae9urnuJYwViAjlj6HRkr+M9pZc4kOn
LPheF8nVhXG/2SYtqf4gRT/qC/W6znXj67witTxVlmGmFiVidsyW9MsgVrcG0YlE6xQCZM0DxVlp
BkT/t7RNFttKZbBTaamnD3qYbvK+xwBGMkRrLkaLWn/9T3hXfkcnCwKVX5QEW9oQIwweLKsdIhNv
+Jf5cegz4qigrqo8srP3ATvv+BS231LRVqvtPTEGV0gUbf23cSPJX9zSkqF3NcNNGgLU0Vr2NkO9
uUjmpXpd5V30UzpK83a/e5RO25rg4O7MvxP6BM3CNkBsejNUpvHCBBKcP16CUQCsvi7td+n01m74
7mIRtZVx57xSVUbqsy9GsTNtwM2v1L58Lj4ZLbjvhO4Zb1ysp4iZs6e39RQnfknr71OJGUtBDP8Q
OomqOQiEItrKwLjQxCeSzLChU/5zox8zlmbCg0C4mkkO005FGzAQPzzrSP4CD0PK+HUuZ6nzVp3Y
sNh9miD5C9HtNZ0orGk6Yosoy4XdPmHF5Qjg1uNj4PkatSSqypnYMgFs4ZDEccoXhrUlczsQ7mBD
xw1gyUp1Quh+5HuyMZbljoNtbJQDnNmONbfZPNlZYBewqFec/mmwNfcCsdAxTb9EcWWALSn9nivj
IyiyRSlLzDFIwLFNSZsyrO/5jUWXtxkKh6npByVU92egNxBnuu1QU5SA+ocm04owvZ6x4A0f+h6a
y38UQaDNQMPzYNPgwtX2z2GfqHsRnCDC3fb+iBpJUjjRf3YyJKHvDDNIHBN0uV9cbjEZNHR+aapS
UCLX4bIyXWjfPIDo3ywhej7d5GA2E09ut75HwzfWSBZwk1sfnBBFU7RRo5EgorJBgLpduzbMXltB
sV5ZEZ5iUlMIm4/HtxLzEUNnDS5BxnyP2CahGtR+RJtbfWbppOlxaAp8JAoHsaF0pjrqHxUCQCJK
u2ZSvZAYqzJRL/Y1vu2fGLaCKKZf9EETAwYxODLwx4wUTHI8zYv+/v4VW45hVUpHZSX0Wx0hx59h
Ollto+ZgrRnZoM4D3CFY5vnQDE1iy+tgneAxJYL97FXqYNPzVOBpFtE8q70hqdM/gprhKOyU9BLb
zjqit1zdGi4xX1oD4JlW7tf+45kBaiDFamkWGxv0tb9Mi1LdKUHD5cRy1szSH+SutPKOjHqvFd/m
ZXXVIi1cE8HGYJtX2eivGB+bdHjehSkRL4bNQGqYJngEZHivfD5VFpMjbD8NVj/LElWEnh6jomES
LPXD7rA6jRYrwjNu5tT/+ZHTc35IEDA9xaNBRkQ0x62eMcVKnJyHoGuzNonBAv7m6CQkWqxTiKhW
RF060g6l+6d4vZ2pVfHZz+DQwOB8D7KDtAD789vDtbESmhyZFLs2O2hUHVMv+IGkdDx+n8ZJxinV
8BtppbYHOvc2lQNBvERAw52HN4f/uI+Huf6YtG2QmQo1d+fbdIjnCeU0jt3/XOS/kHYPqKhpDe3I
WBzMy1B4EJ5FF5EKjxhXK1Hn/JYK0aOFGz14DHRlm1UYFGp+ijXmKdE7+z5EOm3m9f8ni+AGQDA6
Ex7Fv7XXnCaCA4QzmuOtDQBag6z21Nc16zp367d0gbDEHmNarevyC8G4R6+3KbqZVE5xTwsCKh8X
s84VCzdhgWqguHT3d6JzFqmLshS8hPiP/mY35+6VbR7m7CJjpaJfN8l0TaWdiaN8TlyadEq5dCCF
m+cy6rM7UCoc6oSzja7t2ObieJyTmpEnCCxatbFF7LCBsnr5QDPSfScTFL1H8l+eg/hr6Mpyc5UX
xB2isfJgn2RS7ns4xp3pKKKQOuFxIVv7UeYFKa8GuppTcb+eYovs9fdXmMWsGXibfEwDPmrPkfpN
4t7IWbPHFSarSyEJBqmFa+tV+9a+pJiOShttiypJTUzj+PVJYOM8Oim8j+inZ4hTaGxvAhGavvS2
fHqqvRupfWjtI7oxS/2Fl4YgchAcV+4pWmphe/eqQCJBJ3vz+4jwOPMg5HkzZ7G21vNg2XXlG9or
luqRKBhYXwADb//1OgMtKbosrWuU0+5dUVOCTgj+qycjRWa640yyUZ6NMLE3y/GOL9Tg/5+93uli
Kz6E3c06KJNVIogN3bpe+pJKDqDtRWrO5r6AjRSyQtnyMRTp6zeyNntPjz6qBkhq7C0ygoQpQajp
lPcMZ1htobynQdLZpNAbV+rJ523K5knI1ZmZaNjw5iRKz57QvdbzxdrjY0KdEwWigfel0VGABEhW
dIjSGlmtJwFdYSPlAsPuxxlDEnN9FVCy9okMIrQGm/jJzv5/BlOHoWH0i26VYEJa0DN3RLL6bm+h
p66UbhibL9yEW+sTp+eYkTupZCdTAyT3sRaJrLB1JJXVctzJsPtM3j/0aT0ybuXH6Fkgrs8n0rhO
lnZeqmlNkq7csAMliUE2OUxfEhgW1duMDrU8b0MIDqySUBTg4+k/qsjzNgbzKdFWMFkJB/8HOfRg
Y2VoJ2KkFl5rdC5Qe+p80rQZq6DgLzt1DzciE1EO8V9DL0YxcTU7HNK7Yne7ylKl6c6b47fbl0Nc
CjV+FYttbPmj7RQ5QFcdiZDbfTj6/MTSnO8Oq2tOstnNqD34qZgE3f4Y8C6kfyvKlCpbXUzLZ1bm
7rvDJIG12X8g4dGq/gDC/Ue0QJbObqFZ/wztfHDPFTjcnArqOJLQLGaitOJY9ejAf/t2o/l/5bMa
bC7MWa7Nm0rboHhgMOEK+WJ/l4Q6aYCVIKRoccbqb5zLf35Hr4jhrr889dH9c/CsrnoqGyx4k0po
TI3tJNysx8YQzoYS8VrJso4hThoUJEv04gfSHW+zl+PCYk/zkFeuxDZOS/woOcUjqhMb1Cvy1SjT
9AJ8Tph8vH5ruXsbSvFfuXslGVoITXY7jtQNIjnYorD1AbW640ANPoMqPoNpBRJOAgzezv6QfxQg
tc4n35ose9OtKh85Od7s55XgliL41hopmZdi63mfXBa/UCAfm1vqpng62ERkXJKVuhIt7rDjekiX
CjyBBPSqPmZrEUwZAQAUb41MxuA1xMe/yTLeP6owQzfmNzWfgaP8As6dv9rrFcSZTTRlj3Y5764Q
JqlzXOdBJHeJTBmbX4hy9cMDSDncw7m0DBiHLfTxlH0dmCAuZv5JGSaVIZ9dAyGXouBXdcEtT6CI
t1aE1jnJwJpsRtTZwytfb1G1KXwvKgMFLy+CHw1qhcGK203cBe34g6jFr7eMxjqNc+dDaNQfjmrG
6Z0DkMmja0fpXYi9kmKnluOJhIb/FvQgQNdIyAc4GKFGriEzu5Nr+IAhAZxzrDFciWQCNcYhMH24
niEJPYt370zOm3B3L6FBDgvRc3aBJobP1am5k2eA1c16WX6hVUrRSoU1ONeK/SxgxG4iulUSj3nX
W0IUnFLSJs6Yb8ijvKd5/p67m9XLtQxdNCx2UdeTxucgJVI5PpxoZQ/Vp3u9rs2keQCelX2HCSEw
tERqC3WotuBCuH3YHLuAAgzyNBYMkmazGMA5e8wZoWY26+7EVwkqya5c5riiHpVmBwv1DghYAi+v
vq78hTzrDOG12ZVNl9bPrz1/KHeYwHT6cHT/rhG/wfdcmitCtI6FdxOtt34KRwTMbQQw0tYJIc5D
TPWgx9x1ImXPcozAdvW/8ervhU/MbWlWXsStCu66sKaRSMW+flr0uuGAr2wB3PwU/887Ca+oF2Kf
p5hy5LjeI8O86Bl5GyAUasTCFj+Y+F9B+zLKAqqN0UbvuRBj6P7YokN6EcO+p3nr/QR6L4f4Ejol
iQ+Wbj+o5qxqFTALnAJG0+sJmjq7UPLXCicsRP86Pgo3z1AvA//RmCjIYS1lHG7CALn7DEvqqEX0
Ypw69qK1WmYRsPJo805s7wBzjmt5aQB4mwUm5SLvEs08wL09NzE1/aFlDoH6VgMW7/v7lpKey9tD
e/j+yyfBrU9s5MZsK+jxIA3nlmpe36p1NM3qRcc8h+x+3eUKyArR30WVfP1TVNFynyXGZ56pDYTv
QaYRg5j0vig3m0tAwPkeTlVDqpY0Tj4dPG0Frqg7Q6E+iLZlkgB8FZD4q5vnGxX31i56e6ACLM5U
QnABkJzgKuEXCO317GkfVMxV7YiW9fkD0GEvAtYHrJQ/dsxAHRaZ2l4zUlRZAkCnbL5a4Ajd+Om3
QWjc4bHxQyxXZeOcwEN0lkEMkYTWuWnm1D9OscGej4NIbXz5LROLBC8cd6o+ObaE3x8fpuRelT+i
ib7JEiN3gTcLuTpa80iX8RwY619pwfT1gMoQ4ecGOlRGi3zyx1egQjGzumbrauM5MUEw5s/r85VK
JeDIyusbLY54tw60rkdxRxZjP/hIWx/6IO0FcyRUkw0FzZGRjnw9HN5xUubM7CFV4o9FBmC0/aZd
n3w6ASiglbV+eFUxxy6np44tYMaGYAwUnVPmzMwC2TThn9LQEi/fIPK621BzD1CSpTB+y+fQG7a7
BfMFXmgdQNgNJh8jQV5oXyjjdhX6AbA2io0v3bxUzQTwBAEwELQhPuHLBw7DIF9zYmDrot081VtN
uGz2N56lwcmQ58fIu6i9E+emadhvR+FgRh75MPJpyxBLehKI8Z+2KoL0NAoxr0vwWPjIdbbYZft9
of9SmQgnprFBjvET7Clz991rfY6Ww3BA/0AMcNZvKKx6wFMcjWbUuVcd2LoNKQbBMnOKfoMwyhva
VgcD7d/axeB63YrBdoNopi5tOqZSrP6NacbV0BNLNSANM6OUENNC+bnL1YzZjI/KGVII/gVkd02T
sPeKaKMVTAGAGxCuA7X2c2/DiKmu8QR525ksyZPAWI36RNnQrQc2MkfNqh5WOteUwrV2ICuFCwsr
VaYXH1oKSE7MCF5xzm3DQFgiNKLb6za0uFXMEbJEHqYD0Szei5vMyWAM+t/T4z1etEqNDT7RdQNS
Mg078P5NtEoT/exL2u4jeg+6ojEfz/K3nCHf3NuJsVhKN08x5Qs92e/K7QrAp59Dnz2x++k8dSR2
Sn21TVPqaLyYgXm+LrecYdjXq1l6MdXMFUOd/bPzVVusIkoiohqphHB49lp46OEc+hnaImEslT6P
NsSIwC4pOQrKBm1aI81aljMy8ec2ZJo1FiSZcjUe+z6zJg1SdIkEajAqzEYMAD/KoYfvD/K7bUfL
jagG507AD3dlWEH6KKumXCu8NGHL9HQ7TTyKvLovR2mnzttelkINfcUIU2zjTBnFow6lI6QgrcRI
srBtNlSRKrRsfGHlZV3yiwMuSGF2j3lRjXnQNwGo/gKCeW4T+wSvZmtHBtwvO4SFdRh12xTI19GU
utflaOtNFOaIyniq2SzXBGgj3xNU4NAfpWpSdfAti07+1J3WZaCvABvdFPHJrFHbqBazD55lqkDv
DfxQ14hQaeO2c+Hd1XmNEhsBz3e6GRnxCpfqsfOx/onjdrhXrUcVQwRhAEl/hxvjIxBuJjYqCMXI
YuN54tnmFHlKHDG2NhgzU+FDKuiOWK+P8J6xSutM+Yj0oqOoPKyXSen9e1uteK82RM8wAaZJF0v6
g8iewdMod/ayvWBXR26WxcnMowOtl4YiFQ/j1gLta6EsG4EmBN4BOJvCguo9aixXn7YGsToJH5nl
mFiNF/SnBqaHjgTncqAQiAAGVYKUAuT+gbNiIxFVdpTYRtTjZ7TkwGTPzzcyxbDtWgFBvFJeApe/
9S7EZnTypappc9HI/rzfLjfIOl8DNKa3ZqdN5FUoffZt3uUP+KRYZbNFZj7Q2A6NsLy13y5etynW
DGVqBTHIsJOc/T73Npx5d7uGmgD+9G3S0VWzI1QUGHi41gtkRH8xGuV/qnHLsr8CgRHLzYYcfCp5
KxAtfEq35Tnv9pSHf+Flmzf3iB84SJNRHabIlMhO7k4t1tVCnzpHFiTI/UXbqhAcvO6PeMCYcvwT
rApvTZuSvkUXDM/KAznpYo0odKeWLgkNsJdjiOGCHb7ciNnhH6F7nOatwsRTxGEYWqJS1D29tRTS
qqI7hGI5OMkeqzItfWEMcINMuiCcrn7i7GjKNTddu6zf330UhlY4ENz7dfMW4OxjHxSgTXwMXElX
BEBnb6F0qwqsDJjPPvJ5i9n+kBCuceswqe/BWDrhfr/wQPfbWWeJmx7IPAyebtv7JjOHGHN6stU4
FBQ1Q/0C7zMQqeglW59oZhZnO2g1JSp19T+/GtKDAzwmaNpSGNqhxxQSQU60sGEsEiyZ/gf2J0B/
dM3/dta3dpzh3E3UYd+YnPtnhlruAwwkJIuxLYhV/FH/tyVLTGI9CPfvYmRYTAvKyJuwsEPPJeq6
vbxrQq3B0LvXeS33eks3ZX++G+rHaRo7owBNywkBCbgGs/8PIwNaq1jncI818g8gMERcsQJ1/zCP
UwSF984/5dIyMc0B2vqoNyCyIjlqm7qbXeprRJQdHkGOrmofHCHQwXfZg8utmGMQxQLm6IKu9KQO
T/aHz4SNJ8CQgYcTpY323K5r1IkGA2s0osdA7DGp8YI8EVFNLO7WZaRc3/vu+lz7KIsrYg1S9RGQ
0B0+EhScnBQaxEZottouczcu0qx91gVJA3QWozGl1oTHp8RBfG3yIPn5I5EXZmDWRWeJCecBzTtB
K9V2ONcH+gvhcb2bmjB8sUbjRpUmuD5c0/CnKkLQwYHGkfQcYPXZZxF6r9uAAhrezwq/roqWP1cn
xc/6cUnt2Xm8I0YpQyGlVbYT2ri46F0d5k1pVxxHTI/mlApz7s4lhyGH061kGPJ+ciA5IFJCO7hl
rDHQRqBrftcowrmbHp49SAidzs5YPp8Q0V1jbCrnGKx9SNlQ9EgN5hd5PCAGvisfaCal4RUvyy6X
aERfymjgPwpGn5bYwtXN80h2rwz5Loi4TzfWim1kZO/K3JLYzJD1N02tVcQLJln1FD24QQzRtwVf
kftESTHfvxueLB0i1dl3W7uuhhjJBOzzvLETKo6r2zDx05+nTOlbgvT5iz8SXmzkHNdYIHaQnQI7
FerkYOj28rBX/mEbDvhyrV+NSDeD7IyXA706/GwzXzCAjv0zQs4Qj0SZO62Kb728n2g/nNUdKh4X
2/CGO5gEVRquzYzC6yyjhGr5FJrbAKjqBgyebvDmRgL36HjqsVHzODmtoSYJUzMs7lIWzYy7QdpY
pPvkkjZ9DrPT+yqgfUnBzuZeo9CTIyVwR7qiuznH17e08J/U4eYrPh+TXgbyf/W91Dt12hNVIcxI
EK74mZ/9n7Bhojkoev/Ji8Dl9r+5xgtVnGgommcO2g17MZyoLXj8bwKHYmT2FHMCLNsURHs3BA20
vAJdPMsImzHDr5LZaKbCrMEaUKPiJHW4J3RL8TfT/0vVGqSgOFJA7QkfCpEw6OE6DIeO+KB3aK3g
Tr8VpGFw7x6ep2zVB8V9eNK7432twe9+icYYx8FaE6/qAY+A/+on8D5lPmClOchWBoAYiSVvg1md
cK15ROPHUwVmN9yb5jUPezOSm1/gL8B5MY0yT6bFD0tHgmfhO2E9kNagPrbvDxFmutqFm8hqjOyh
SKtOcoVxYgZ+H3Pxd217L9SZ7x9c2r3oYq7RgY23Rv7mI6nF0d3G09co8JHLttb9zSdXdVUJmiud
Qd2spHBxgL4mmq1mnZZ8dFZT6qYiio43jbfF8NwSgZ1GUZIqhSOuHx0LOGQi4szOFLhRMQRsUyZe
juH0zF9HL2Spf3yn8ahDBiVr1katmqFdNhlhFtZkBUkGUZPYsmFxVJhfRpum/ll8JASsKXKZFk5c
kAZ6zJFU5yGFrbvcLIcbC7mR27FmDNrpYgQNjez3eKQLEugBteD4pYmLf2ePVV2GcsI1aPYOQJwu
ag3F6f61hcBYplNCMpfFs2rUqB2ErtP3A7ZKViglsx/oUjDYa7yQUHftywp1OkJV6mBFJB4FWIjZ
WAQprsQk579lEfPlfh89xGsNF/natiJcW1NX1+FGWaIbvGNOOGV8GT8VOcYToo+ZMVJnWL8jNc2j
v0X871lgz8yGR19FBIFnVW+e/zraqSGjSJWyl7IfyFfNOnzhUIrL/iqV3qw5hPl8f1r0w3Cy95c7
RsCnBMiKARGg8tV5hhNATay0JdtbJKPPsYMjUaaonTRnfDgjuzz0psqfY/p1g69bEwLnCxnS7rUJ
4h+4BDmupJoHc8AF8LtbaCD7xAMTp2uHFKMLb1IJhwlyRM7jQyYk/MAtRYkTMAkX88wPHyVb7OJr
ygN5V1xr6VTAMQz6KbkwYB54LU2dt0FuptTXwJnN2Dre42ICN/CDQbrjXFGJnt/M8IYYFLjlzcAU
LiNMEr+dgxsz+IG+mzXWr3G6N/QZRlk0ouNuA7SN4xDisHtdMwIiL0iWIn2rB/sQRHNukKYy2GmV
oSBjjyCd9A0mD/tzBbmhKZeRAejgjr1Tg2kR3jDWRxzWM/uoEBSb/27g6XK949A31XWg4PsPpPJ/
aH8SHDBJ9cij+YiqDgFsrWsBWiE4vuusofUdN6CtwBhSK0/gYWaqVT50ks1JIaoykoMkHOzkwmfb
gmy1YVveJNgOtK4LO2oJUEnxmTx4dYZ1bDNncYB4ghEH4A56ZQ/DpJlfJLo+rxUTqIOUcGerhuNn
lGvQ4Szym0YhUfJj5yYczRw7F+9x/3aUmFNPOTMZoYHLMy4l4yNTTOAnr03mjAO/fjtcBfwRvZHd
V0/WQaNUjPcmGRbmOdu+GOmx+ZzZPb8sJscyZ3x8kLxxtbKH630fA5vsH+ValrDS0cbxKHXcdbiy
VItWQcwic+o9g1zyo3z2vLAMrx6E37yVZZff/boVc7/ajpy5C9T5hCNsgimJwMNRblEmKJXy4sUr
kfaDlPHWukVwFp71njloyzinGTik9io5d3JUs10rXby+TY/X6nBIRbZXjSZk9gvDLain+qz1PCKX
ZgujCqqeUHe/AdsWaAiDTZqpOxCKPxu9RkdcTEvxC0ElW273NSMEUV4nK6l8RVzQaw1x2dNncD+o
EhS+5FaS7SY4KIaCGs0/Qsz1Z/kgZLXIhwobkxT07ZL6KUCkJFQAvrUQS4sGJNTK2kogyoA5i7Z6
mk5vu3Pk7T/8SBm37XZqOTrNQN4nl5YmoRoqtJTAGvlsiqWxDZTA9qJcpW6ah00nxhbUnHXrR5g7
cjncISB2UoCjhGZyqyEgXlUUQfHE3VE+chxaN/25NDp2q1An9zjFHpqc2cPt3dK5/f4yX2OxovHE
riP1V9iQa/wi98MNBmUUza1gUuAmy0Na8Eyxg6eJpdCML9LsU6nVyWt8IUXKYhdGJxzx2ASd6SYG
Jma0uQ9vnIk6+SowLFqz5sueMU3+gPwhBp/mkDp73KjN7DNRJwFA07UigyeZM/KejFNNxTXOBHUh
YT5lFxbewU5kzWhEox6ADItKRX7uE5vOTJXWkRBl2/zqlgAg4O4nuPevt8qcgMoY9oBqUOnL/4u/
l54CojSoJikAOrV37lrEiObOy4/2ZEQNpT2yrvYwHCSHEq+TT4pqU3MiGdqFZ/lgS7HRAIu+DDgg
28AwQPLiJ+hX1vUKbwZFuKsUj9b1D8GeKg9O8pGVx30v+ZHGhJ3QdZHiPbn+sOI9WLUg/ts9u0XS
NA6sDKT53h7C7e9aeYWO9lVThQ7ycqIRWXlhm4RY6WhW+LBXe00lV4F5AN4PXKUvTQYaGLXORkar
u9M/lI7o2OQCyWn5BiheV7f4tNEqcbvAcuBdzXgJ+bZMbOpsCPDTyY0DN9Rmq/EfPWKDr8GE3d79
K3OEzg/OXBvQW0217dIarMe9LWWfE/YSqWT9HHF50Jw++NwQ16P+AUiAzWNXFmvC0Pq2c3vCKZZ8
iWjiDzfs61Fcs1iHdxuOwTKMaiw77/8Pevc4jnqrhwS3NVLAUlGIvVRRkyq/edTyie5jDmE2ZNYa
5JR2SLWeqg9MLNX5WXUQOHTSAsWo02Iu3UG35kdn0JXXnpo6fA0T6JuHcvlILUEdo4Kvk0TbPG9f
kvWYr3QQvR/CNJ58tvGnDITVhZPiC9guxQNPv3+X/w8ODWCNikWUCMx82tfXUt6O2jzAy4eSDj7v
07n3WJAUKC3187yshN3nUzpFYGlm1gDuy3ejrOduLQGslUahLeIBReHyjRfg78rsIFdctSGRJDiF
BEMsiAVQLmCtqASbZCDJvB2b/KKLJC04tg1tZak1EKHK86hQql3dFpU2rOWgmaSfVi+u/VY2FSdX
i09Gbc02hFxsriG7eMc2PPp203/pjmRVarqXbdtd/XfWA/K+OniDirGjOt7dUguGgSeaKfRnBZie
fWw7sURLuCQiKRjhMTvc/yvcjsxGa7a4blsvNc3l5cOBhgcQgP1FDwKCg0F0LHxaKxeTpkazsY6U
KF1VJViplOnbqfLvX6ncuUW6S2vuukFL6wZ9r96k28sW1PdWUu2qSbVhDuYi+rW+jDnxa8mvlscm
S5SRexlMSQ5sGscqk21bXm2whote8IZ2QYTbTtCwmsfdCu6VtSuLs0Z6SugM/yGdWb9HlFcUfxJF
4Mk8yOQh0yi3qZYOIFbcwHWeRbkC5sJ12r6tbONQDhGhz4aFPbc4kRCpx3ZLC3i62JXpbF1itiDf
f2PJMjlytHOTYCmefON8k4rhx6v59O7EtnXz4pyTXQdsd2huu4CO1nify5pxbeSeVC1Og27eEHvg
SLw1WG4uVs3rruiWXWRIf5VWMVJI+bwnRfHh9M/mH0nSLc+mB02PckHN8lABgwt1KcduokzeBOVy
pY53H9Sg1EJlLV+uzzeZaC9NO5cC33TWBVHvc0L79Gau0JZ9ZqEhv5xIi8afrgi0kf5Ak6OqELFi
8lVMi4XhBbAiiLUjYIfH/nUT35U2RvJdYQ6pDML7uV9yV2wIAPyREG1N1YFgQyd5njjMqxo+vIW9
ABscpbHtt576sinAzbJ7TT9WZvUElhQ5R3iADzh9N3EoxRpeS8T6c+bLO8qiC9SkhH1x4x99CkLx
BHDXEi9IBdPguLliyoBW/imqyIMLtLSBpTxuOIPse6Yz0LaKmATpIoaXN5ZJm9IyDigsgnvfcubg
YOsZFHtelfNkacPDc14l8jzsk7tpjKBrG19721pE9IclpygwWNBId0Fk3MRB1vKR2U8pnNHJvMC/
DirVKVH/InFg3mxPLkY9djC1CsWOXM+s3MfvA104VZPe1Iia8DETQoGTZVhtskbJBO9B+Fec5re0
Ga+eAp8yy0ANQScVX0B6q6lRLYdIJQQ84vQp98HzojQ/cd/bPpzdaajndqKgoOnxt5fRt9KsNMzz
k5VU6FHpo8zkx0xz3j5g4kXBvNIhflw/wd0IFHvZUGVYAX1IqMGS3jv0g2bLIhI9BsznW8r21qy0
UhFtcgstKmV/QrnldpTJpLFCNfVJTafNg/4Ool6MgXb2+kUxPBfCU2rrbXDuybnv7NkLWAmfWRU8
1DtlMSoQyXMKTqd7mdalkXBLMKFqTqURdaIFSxBnYBpH4tU6/LpvDAYKP/vNpsYgMCZeUN6CX/Sv
oUVR9icM6B3bEQS/goNB1uhxlP8D1+k60xvKbZzjbDPLdSEpmyv1BycUARKDL1Mo8XYec3hpB++w
yfz5sR5DMcSC4/oGraZi/UcwlhsAh57btm1CWiRNiQZYDqODlK8bBtae1HTjWQ7rCafN5yIhNyuL
wd5hlGIVbdMjkY1+pWGPlCtsnqWhMvtfm5L0JBaOUhwwiHHUKZMetjh8SeWcu7ZqJPIgj1Y27qWj
a6wt4KJsJuPnljMzX/4uIsE5IU8jVzcvDI+q33uOAhzFLwCP/JGLa3AT7bhJrK4nBM/9UzsfpbEC
J3Wf9Aed3T9vBrSz22tlZd88DSncY0C7x1oDQuawEKsfgeFRdHkkxfUZsxdbV1mdjv65TtlQry2b
16eIos0MMLt6HeVCl+aXDB4jVjmgBxUWFvDn+p0zDd97VuAWEWKJzSPjS+4ddZVXlXolzHxo6Af/
jG02GYz64TTBbyF43pZmfo6fsOP0bkL4Y0vMJozyRDdvt6T2RrMbtnP1lm0hDKizxf3QlndUs58Z
ObQn0Rwohvj65RMzctJhVlc3kQzT8+dbZpkYtHcXsYHLFy/bybgvx/DUTLm12nqO/7ecpDW/cybl
GOHiGNQqghXLQ/chUNH2lVmDcV9LLPpeskYCSJaYuIbbC2c1atQnxazEoISmt/JtBtWfZBy3Po7f
x6Rn5hYfkIPGxiZikGuCMfJCNXc3EcSFH9ELHneXjYCTfpVSaul3VSzmx8oU6QDrRY2l8nW79lje
YyaX/9u2+KGDwUVSTofnjcNc+huRXBXPfWfV3dKBKpVp0+5fSog2xjgob/bIW363iO2R5bXKxRJS
K9H9+GxErsun+SxiK8Db3NHQMAtnXeZOaitGo5bFh8DS9tK4TOznePlSPZhLaUaa8vi0HiDywgIb
JZqylKW0E9EXQf/ba4u6EpCAYEwUvGeqGg6ao9h6Hz0WhV95joBpVdfFMhZvqthASyNyGKGvgdZg
KxJimrW8+35HH4zj5WR/SD02/YXLx+w7QC2ODIg7R5PATNWAnos99NMFfdJa0Qc+UL9j3qGd2fkq
1HTEEUbDLQscfGJC4Z95a2i6dQVmZmTj9Nv7zJvj6+/8bFs6V0TNuJJxYZIJDKb8Re2HCtwrEAyB
sfnwbQXi746usFm2sTZX8I3IAaGB+Jj8iXe+81nmtJo2Z7DCHg0P1XtHrs/AzCS8Vv8BbE+OI29a
N6SAZDpYsrKFhi9kdKqTsppjBS9lxkfvKkLVYppeLmqZoqQ5H+sFDw5kg/cBKPWh4lMT8/lUV1vQ
hqnL0vZye7Glro0Yx512jwszTVVNxdXcsTNMHQjAaXUzq0NElJKgowZCdiuCN4A86dE+plPmknv+
ORLgOJSTUwcJWiP/fz+uY7j/xvHwDQF9+IfjjPxXuMGyP8Dv7oLYTGkBdzDqXwrcNE1FnIuzLGri
DQNx6JbfB+Y/ZVnJ1jGA+oAgZsy4vHXAQzIJCDVXIbAN8a4w6uvXwp/KITSulq9/nWYO2+ebq4zI
BJQv8K+el2geVxPs515AymnPWnSJumFCv/IP8L/8t4LSwjp3QxUtycDtZxT3NEmM4GkuUvpgsGuK
VrR/mEEf4VeP0I9i656Pi5IVpoWIB5GEYwjqJ8AHyxwDJSZAtI5b4RAWQO1L8tKvbXjB1n3U/vdS
Q9U8cfQ6vjxgIFkXCMm51Mt5M4Ga3hfwDESPlo/PVDPry2Cxt3tFesxSb9cQaH/fv/YVKVLqwQKO
GCuhSajMS3qwQqeLSMrXWem6l+WJTiEmcM9N3ifkSnerwO/joSvgVWAL6Q3HWPQXNNF4gSMWjtlJ
mwrNEfbQeIms+tMzi73C4CCuzr7jz5JSHn5Dxs9ksJ7nL5Ku4V/CIxWC0VawWkKfFM+Y6YpYVWlE
8ED/frIujpC+p6hMP3fYq+oEv4E5xHekbekBJ1Vc08FEXXsnYMfgqzuyEtECtqYF0pQ68he1DfJC
w7q1aMvA0O1wo2w7i3iU5ynR21NsJzkEn85RRE5lC5BDg+pAC8wpTjS6azENKBX3WWC9lHzJAMPO
I2wkTlHTjd6eo4OQkQC2D40H/nsry2e6ndMVIdDO4+BG+tYP0Rac9MY7IcXaQFZ1Qjf3cpbKx8KH
aagZrbxL2q+2Qhm+vbeCCTjJ6CVS4Jlvp41aW5cJdFrv+aMTSlB6jJWn4aRF3uGq+32hFDmW0AoB
Q/K4ofMqO1anop3PLvdGXtxzOzXRZUHxtgj0UYmsIVszB2Om0aaE1zlPQ6EQvYJG0EeCEMcfbiCx
t3Kk9R77x1NssRRBUX7HfYBZVMYQL3+JLgK/1hYQP2lVBblpZYnFKTPW3kZ8rV6BC7Or76tSYVkE
PWaOlUVm8mAp3LbIDcMhlKMm8lkjzel6eB1gI5KfAGSc/wkg5OcFfjefrSqNLsb9ODhgJgpUBo3k
FnMlFO1y+/lFgdA6zHuELm94uKlRF/Z6O1CDMkcT5CAqqksv3KXneLMxRkIE7rwNfIm5sIJC3W+H
isQ8rnipaPtAkQXz4iHV71iHsM2HOi5U6tLCVHgdunkCr3BlOVyO7ZKqcahZY4KvCFM87GLYtHGf
d9ZwmsMINlYid8xlTQlRCWl1ELu5r24y9UQTJwwJ9/1r07Ne87njcQLAll6S4FM1UElogLPNDuL8
ZE1dTA4MZF6ZjVvSgTItdc9EIyMhjLuOPgRv9Ex1+WOkUGzdNJgBFWQ760QKocnmBB2/WNH+JWD+
tBp45rLcfbAW74d5swR1DOE0ahSst9e4HaVCPnHsLdn5JpzMTxni3EOh5++SnTva4olZwfJzdSAo
5ZjWgMrmeEF5r2I0fBmuyo1man4ihSAukaYT5FAZnATU5kbEmODFXitRJnMRNDXa1U/aicM0ns3Q
9JGL5OLw7j9wuQxaErJ1YUo/S7XHs97M6caGSQZmNOKPmLsv4UCMEfA3hY46gKIoEh7KuJTV+FVA
I9Hkj/Qmv8A5c8FyrzrrgMUekNXA2vamRbOvAFnu6RUgzVcmEwvTxqigi32mEzDBjlnhdSVBiklh
kHUbu8w7clZq59UmvN76lYtwX0lZORqDzgQlERpS5d1Lju+ClpctFSXK1GuxAdGKOYYORKg/h0Ts
mwYWq5pvVHCiDyoeTVXxg/RKEg4bFD7mCpsK+n1EILG3WZSH4q3MZlcnjYVU3A21yJFrSl05Tt3j
9QqZHd2LaSz3DP7HdAWmdgT1GmpyivCE40QkwkXbsewPSOOwP/wdlLH8SWgJxj7HiAGJasm9afEq
jemBo+sbfO0q4I2y6w9dGNFJjO0vT8a/qlXH3l67QsD1/VCmdxVLEcat2AWOFFD2FF+uOWV90Rbi
3+wImEDKIhGdwOJP7i2N93+CODDo3UbBkvx5Eg5+kwJPoBQ7reSYkHEIISt7qwb2DX/DEijlKTV2
jqpNY2xeJi3Zh90Yty0HlJr908cyZub3lbwEPhBAF6BWz5Ok1M5fkDOU5kH2kT9YdHp+nUkX9CFs
646dQ7rOdsW3MbcpftA1G1bxPfzo0/9qw3xHWwuYmueJ2aCH7juR3ANnWluVQHEBkwPPANI59GAH
eiqZH+vcWZ7AIw8owaIbPIQYW5lMOSSizbnG4+oLzKUlJIYCizRJ0SWxqe9HElbJinTAEgU4ulYS
/R+86NX+WH7XkpQp7+F1V4rZgGbk5eo9hpN+SsvRdB526bqzZn9oVJMJYjEbAvhQtZK4V5hxv05B
y/X0rPP3k7ChBos9EN+cHNryPv4KFghmXT2jdajJ+kdjSD0ayxZIdSGy4p+6qs4HTZt6P7R1aiPI
jVHAn9EQRUi/fm5q6Wx+4QAcg1rVcFMMrZxJkQix+nMdzGMeZC+ky6PgdOeC2SKc74mRiwPPYg+8
AtuwtEld5fPtiPiBp70NqnaJB+uQ0KtCI8H5YbcamVX06YPXn27JZQ==
`protect end_protected

