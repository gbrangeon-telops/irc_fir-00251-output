

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
JtfK/+1JKYw3I976gLBlwV2xqGRbyVsJ3RDvlPNJRewqWZOfwn5MuTyc+U7c7Y8NUZJKZ6RY1Q/g
uXt328ut4g==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
SKJFICLwrmXfYqYNdiUThnnX5tJzUEdqxXF+PdKpwSGA61whpH8w+itTbLnn6xyBye2kcWPZGi5e
86BY4EjHm7kmXxm6GHfc5MWAMFduB72GxoAF5LRKlUMCOdVsZag78zFjXdMU64ClBQ4zjB8EgXvA
zXBqthWa876wjTEo86w=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Ho0WiFevcJjvoEEaYGtHkcW737RD7c5clzugQBBm9an3ZkyNmpivYZbh5x9redNVt0HOAIz4unf2
BSVy7qVCwKIsJQlB2q0JzVYTIfuco8FlNbrUR7/BeLSPV7XOk/MTxR/0Dg6meFJjnWuC3OrBGp8S
Ul4C2x7zg4t68SLTuFe/LzPmogzBzDfD3+nozb8sS3jX7ZaQAm/T/7eoy3grLVkFjUg9uj1IhVTP
59FDPnvyx1zZ/V9kzMjvM4XKEW4i0DGLbDEkqT5cZNTgcxi+sBHO7OnQuIvFzoIoNFONwh8iJ8xI
jfha3bFVgIjIJWFL/KzL8e9Uwq67H4YDz6GAsg==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
tPUgwDCRFsMzMdJqCXSx12cw+CNwvndABCoiKOSYIqrjgxTgSZ1CAyY61ekJUz6cu1q3fnTmoaAx
Nh8wOKV+UbnkqjbXLltbzNbjSEawEnAI8RSn8gStXvDoHe7R6pRqYg2wbvEPk6N6UhaMjVC8JxUE
Nl+LL/ApnNDqgvTWrcs=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
EyCeFS/0OQO1er1RAmOJ0VIpIQN1auXP1dzcGUAOeSe9eyc/jA1mhBpZ1JPfDCNxALRFgLLGYZec
wCmtwGwTJ9NXiyrouRmXyaKsTpp21jNq9KLTxpWtw00JZFdcekT3NPcfNHa7nkycvsM6yWSUR/cD
frws/8FBuaG+siAqTh5qClTqkxCmbJ08Qh/l3c/D5bCXbr8wXY+SVe6EK7TiYFpV2oOMuwWw5VVW
3m3/ZK4knJ1G5Nn68ZhcGx6rqQE9ZbHMigIgQyt/y7vXemBfmAZ3xkMsYj2X3k1fFfReGPYzTOCE
6J8z+FWVfzx6XMFACHDbKayB8gE3RAvjSqIISg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 7056)
`protect data_block
Wx3XCFB0PA1oiuyqmwIk4U7F5EO+9e5YStBclEmCsj0gEo2DW4fKWjevwuF4X/6pP13oSfwOxJbZ
vfT712MSBTIjIgi6/QPjfbfjOrYplBWfNHARJhE9FRocaetDWnFzJrNan6g6y3rcd+3hWf66xh2/
H0WaZm8Y1N06NSC8wtn7EoCK3bG1ifBhmAkS3YQQpHcpvGfZEI6nS2TEs89yo2KsGCmJVUKF2K7V
5i7CuKvaG/WN3TkjA57v+S/2sNWyMuCFj30AuzwG55nW2UlPEVhQEk6Y2UhN52GESorvQ/RulJvm
AakqDPVmnlHEJ1zSXRONRtmcBpTg4WCIuky+ReCiT7yXghnA/F/+DM6zaoKEvTya9FYCkyXjFKQ0
XnTB9VfxQphoMJComY8QfKNhoWz+ku4assN5UfzWi7Xg+x/9Evlo3gExC8LJCHnJWOyGG/S40FOP
vQuMOrU+fXCWyyNdxMXinQBjl8lOgapN05pGp9feRhHb7LrNMH4DSTKtM6dqgzoAkp7TiSuDFFBq
9/8lTKv2UejzwaRpk667VD7zl2ZX4x7cTbR3H4EHCowcCoSb4nm1ViFXVej028khF9p0ljBF6kfb
4ONmoeCA6aUJ+82Ztg+KFQ2FW28gK++JzMjE2PQ5W1XLD3fAfn21sLbk+J+5n6HgBQmVgvWCZxd0
7T0x+6offugBNumOpqTGD+xQG9guYiS2cdBlkGHe4aeZE4hw0CmVGTFpyw/B8p85DPUmMj4bI9HW
F4+krMRi0bKJGC1UPpav3L9nJu4l2ZLPm2yUuWCDp8dNQbUOBieF04cnDaemu1/DF2rqSyLfEneV
fYkMqSttVOPFVPfePD26IMfHC7NNVviZy2KjD9Gnyp4ptK3k3RrYW3ignUyzsIaEx9lrVntJ7ZUl
Iyv3bCP2e7gRsxJRoS15G4x/jvuogws/gGn2uVWpseP3lsGPaXXsFuv6tjGMBOK85DtyoyoV4OOv
5RF083c1b4fybH+fJVN98uQr40PSlxTQ0DhiNj6AoNds6PFaEMNSAsSBgp2U5qCKByMAOqroowKN
0Kbld9DHDFCRKilZ65N21FKJdDE3YKUWrti90WQqYERtdJA8qm0bl+AViYrs0zwRK1f2s0R7a3Td
+GMUXwRPDMPK1tO3m2MvvGxjbbhGCIogJUdHpRhggfV0c7bcjWfSNsew+wm2g69tpKMg8D46RGsH
oIgaIID9JHTknnODm/FBUymEmDLg43cSvjHni6P1z1k4QxJZhkeLEaWZ4pDUKpkk4Yb6LIpMO7eT
cx4SmPtOOYdvvPBsCXVD0uWGujtOMCGQs6A0CXOMWRie7JjcpdV88IDp/ZtXDajGD/tCNQURPTmh
kx4X93FWZfUliGWpiHmdBb7Qh0bykcyR5O8W2VrKGHIWKLHrOpVIGFKAf0WIGSqMgyfJMu+f1a60
HCeqIJ8g7zI/aKuaTrTdYkxfcHzXbLYrdPJlahajYhYBLPxGLdXpbpiint1W3kdU0RTb04qQ8cMr
2XcNBPcXcDhJa3z5rGn4NOxwRvLNrgyFqlqjM35u0X7kyjT82k3wXnxXvUpzTZnhKQChLoyQhjS0
IC7JPMmA8dS920K1RWAOuRdXXsLlBy1fAwH8yepO7+ifkcLlQ9zcPbZC07TQX47hyLdmGbyA3m8J
EMwWILz+39cIpDbgIKZjpQyGM90KQYM5nR5Yx+GmwOuXHTYLquNI/xzWEESbQeOyqOmDuzrS3D17
lElBstgwIixx7TgHOfDTELP4BMl2R+ZGTskda7BrDu2DB3w2KBvX/kiag1VEIgUriHVopV6DYCEH
1BOKNVvsEDB5FSuPn6zv2tqY8NLIBXuMthK4patMDbbdd4KOS2nKgOdQkR1rO+H6pCBOieFSXmj8
F2vmFZ0pIUARrhz54IfemRg2I8RAeG/Tq/+msf9WtLzJzlkKZPjh7Dk7EhMZTAOm1SvSn1OLpk00
eAT0vZzG/PuEJD9MaJupobIw5JLB4BeR0z5TY8jB4COV7wTbT0uiTmO73Mcwo1U9OduWHp4rtLTZ
Ps5+tbBnVYPiWDEQVvHRZ7cW+w9wiWi1vaQfWfxo/2z2ZktN+UE+x0YCj+pOYyMPfx4JMc2jv/dY
AgMQDg4sHK/1RutpcYU0x2Ydg3j/xh1yy00Rq73VhNzQyY8ZoF7COGUl4Q6qZkmL8j8ojKb7Tg20
zhwmFE2bPPNxjeDRQcPITwxaHzFsvMZOhqrzphsCiZU8yEcNOk+HdwI3MMkcVKj/fGwdKbfThwWN
GdpDA0hYYt0VkPEFqIlSxV15ZfaTP/EPd2Yrhbx4EX4k35yI6FVhBUlOhjcihIzMtLBkuwBSx1CW
sMFbQ1iTgKqDBuhjYron0gZPOa2mA5WLZ+gcijC/9ugvIjHqfYr1EaLftIIPtu00/4VI60l+wfFv
n73ups2XBN3bd/ZKSZwhErOkyma4DUYgmFdPcisFgswMLUF1nMN2U9wrD2uKsMrlUkFFkByOXnQ3
GZyBaohEBE+2QWLr3bMTZn864wdwCRC7FyssP2Xkh22jAslaafjP+QEF2Pqfd3Yd+ern535N0HIK
epaPXuPWZkcuYfMA/wfbWAkWsON5ArkeDZQQjhZ1Cm7YmFAjkpnWQC1sRB1L8bs2BhOF5rT1NhV3
fKdEm4fdFTcsTOtk3Q+4tUXztV0m9y15p4CRqpjD2/TKlKVq/6n8kRB/NKDgOsjDbjiY1BqGZPQK
hGXraXgN1hIVxSL7bJXWJjyShiGFvB7wvchjH8b8v8OgJ9amBPaMW0C9slzTxTj1vUUc0jTzVNG6
6w3DeBG6hl10Ub82+Web59ik5MQyeUaMZtrB+T9/aj2SQoTzOYHOW2L4eG0kdCxB1L/PzkuGiInZ
16/F1B11VsJqQS3riuo9ub9tlEXpCEXnYRWpFU62T15X6briujyD1H4WhlSXbTrUo0xH5RYtYBmu
WHFpqIRr8wtzRs6BuxCCf64vllVbTfD0pHL6PzxbOh0oILEwfBKcM7603SDDT4d5/AKbpRx03p5N
ywss1saguDxEqYwwt635IJnNjHdZpvZHCi2Jco/b50j0IbmLZ/D5MHN+txSB1IZ/tDrYdqm0nydw
SmzaH8ZF9LkQiczENQX8D+IrtzYnxJ9REGfzMLUkQfg5h5Sz34FVreVTFNjQsMEwNtFDIxrDWbk9
9GDxPq3eS5GbpGT05jJCT852qqpKKtvnFR7D68Qi612tLvWoQqCXdKg03G6YvPGVi39wBvITshK9
zCKebZw55Mk5Y1S40xnNLgnmYCGaQbW22TOeE8b4HkUOElI9Ir9xkTPRTBqnOQeGM/VM84hdAIdz
/hIyB7/mg219lFt4fJMDUe1hfN2my9JbtAjog4VOSnNAKonWfqOWMpvUM/h4SNb6cSgj2zZWHR2Z
xtBcDyW6ngSMnddbBqluHAlHjwPnfA26E7zOe2qYndW8pIX8psK7FyzKCl7h4vYnqHgmAGyTuZEE
TmJ34Bn7dLlccW2iXvmvBiylyidDnludOueG3vveiBK56XIjww+TQeidCOEsLLoQXRRkdK8osAgS
BPAu4Tl6dasT113jtO+xQqJwBEGiQBO5kJMuupkmbDYs1pzhWPRvIQ50SSVTxHxwCcVhIYceE6ob
+9/iHZOsslb6iQPlpJIe8+TIlt8KxYCFsQZkbjZIhQhdC1tgxuDvfSvB75kRFlGUa3Tygj0053a4
NvLVDiiHGO8q88e4cbbon+g5P7Vd7bu06yHdvWnkBkQsQAnBw6jaDfp2yk8qnpQH80nEQI5acpQF
yEakUcC/4LHkvZjUzwDmSiTbJIyfLSStqhAhb/hYg6iOOf0OQsy5Bk3I7hLnN55lm4kzesTKKvAT
peyurgfE3Lx8SMl06kAuTUqEMbHHcNpJdX2ih+eTmiTG5UuXCdo16sB3ObhEOlf8uvH5zAjvdKLU
MOmrXxflWa5Ln8oFeiVdcB9ErKU82xIjyO/fM09mbzaq+39/e8vUf3AG4cYGSdZc0TDUq9cX44b3
hE4b9yTBdOu5aGg/mnA+jyOHWMLADBqbv9c3k0SyHzlvBk/C14hGQU4454cmUHNBha5uO/+aH3HM
FvxS2+/ybnTgqj4SaKxwy6V8ipHhawtpumR4pOFdiyNmRUUtrYJ55IuI0ovY5aIhUmBZRnADfprl
rmYzNSl3Znnh6qSwSsdL9asDAZoh363uxAV88PCZnJgYoTzVltNskcoHRMorNV24OsCC6HVu77lt
MtbWxtFOxToXPzJSSLg4+t700ml2DQyxsQS0mOwLMbcba/bmP5ZyU/TOhv21HLAqv0rA4g6/nNgS
vTc/Ky58Yf9AqmPxGxc2MgXSjhUIrtoga6IgjYiqqQVw7i4KTSdtsknirg1i7T0RfUuzH4WWbCBh
t0t8okdInwmBG3RbZFOIcFJyba5Xb92tk7gNR53vug+RGXokEIQNqc2V2dfRKo3PtcVaJWDI+CW7
Z5KM/XXJUHsW8Hw1zIrXpQLPV3vHg4Px/vVfma19Zo2r8Mg3ddXaEWpwJrsE5eL3FlfXRsov2EA4
vTTT3gC+NuNA/aBAshmiiGLa0ykBWbx3sHOmf2KQzoEYjTBF6AY9Cwqo28dKRILbrkHQ8xwNkcoP
c+PT/w4OvsysjNQ1N2GT9UfpyvzXmjopX+B9sPGyIIB2N36Oqo6+575z+hdK0YoL/rDG+1xyEJfj
Ys6DvZMKfjKDxH8zuJx5A/oJsnP3+lt3U6xcSi7DHk9vbOXdzM5grou6cORWwWsmwHz2nBRgZpNn
ZYLJlLIxmsIHZR/P/98kyDPwPIndvP3/LpTX5oKFrP2H+nWPdmqMXiuxZ3rdcSatPVV4GEgV5Rqm
9FiByXqjifzQnOdp3U7ptbeHbLzZLVW0j22lP0wrOPYGbmp4tm/szi5rhZ0NMinvJwTCkuhHM99G
lJdzjAC3Suy+b+VXjv3prJyJUcGB8dFXsMG6SdnRRW4SZ3KiaUELVwFERjVbpgZLpMSrTit744aE
KrQc3nO//RvpC1lFsU7JyXFbFVt9fydcqTuL6u8ANBRKO6KyidVoMODxqPv9RKKe0V2A/pjb4jq7
i8zRi9mCqvsy9LbUIX5TQSGAmsRqENh1Eo1nBFYRQhTMlU6qb2NZgH3oE4VBscCwCgD+GPmgO3A+
Bp6rp/m4rqkte/mcF2QZ9579DhNhMxbqyu1s8FT9b/clUrRRPt7CTo9QESYUFjdVFP7TdQxYSLfH
boRoqxZ5R9nRqLNL3WbwrVxUu+6c4GsZGbwgozmy5ZhwYW1lwdJqrYAGABMhMOEllpaIDa2+C65K
9zYZH7ubMxHrXDzuJa5PEA5zGa5TGmbvjhUhpvTeyYVCUEjSby7xx1NfA7IQGV0/rnv41wJvxfCm
xrCpYZm05PH6EgIBQkHLSAVreljLzIPJSCOfGMYKsP2fxSFPJwi4N/5z47mG3+n42l/+h2wxLtMQ
D4jtHdewZfcmHHNOooqk0VQ6sh56Sx3ft247oAlZOS4M+EDkhcBV+yhuPGyZA70Ywxuetd0A5nDn
ld955ZJ1nAt9v7vqy/udrJWsntsX98Z2qBxETzMSqWMHSdUdqSJS5fwKEemVwa4J0+xpQ4gro85n
MvGX0+QKZ8q+ipQtDFdNUrq01XmZTvQwmVP6faOJonHjIDd3UVTSS45ziOM59KbkDBluaLBQ0J/k
3VIGISbTg7GRdp2rzZ1SheKqn2hVt2Lf6gtqcAwOtPSul1jcrhDa43ozxsHIUYdqLoUoNdw8zsWE
3qwlIihDxvxhc+deA+7sKVSo3NGyGjeDIb8C87uzIjXW8J08yLk3M2Sbnvbl7k4f57ezIUCKcMnX
hzcicveHgn+KqldPuvWCjtgCcswCYTKw6+FRaMTJlZr1JjupeOeUSOAvRCoSohfOsiYQ1zKL/3YR
NOHi1HP2PScbqo77XcryzgqZ1ZycXMZyJUn19LCsonvIkmkhb2yLiV3W3Cq/6zmiTfFslNai8KjF
Hx715Z72YkmR0XLVe3O2Wwa8w4uejG1Kx07beCFsDMOrW8HDn6fRib2cjesZ+umFg/xGEqMPP/ZI
+WRAelC3UWggmzf9/f6Ro5cAMh/usnNhZrum9h83QQqyENNlND0OKFPvZZD6vx7R94xYrX5wHbem
oLN3ET5TDHmntedF6UTFeNyuKf4jzhk+5Mjt9pbzHYm2YeQXEG/Oah7mZ/So2tIPjT7AyGqiWpVA
11ABMg5tizRWsPOV7aNw+0DnM5jUfvYk9MUq03KfxjS4JSOjobDt2mwL4YZ6aOOic6CVTwB1XoOk
o9MkzrQn0XfEGZonbJFgcu9XOVo5wvqELbH/0ba5pQu+5GQXiw4ow0UiMC9nWnGOt/3kr/YptA47
f2M3oOKpw1p7Kra2TROH/g0wpXkbfi/4NbGflTFEP46qaL6HYyp4yZ0xWVnQZMzNJmp7nMHC6m39
JSL66qH9LQ3Mzx1BVFikBINwSSXTAD09LlzWxcStIkSWCSX29TCq9B6BADQUmCp0UYqBB0DHg+ZS
JzExBp4xG7lj1x04BL7x9mU69eobx0+YhnZYHTJq8d8MfvT7ZAKqeZnKC2LC8UEj6pzKFyzYGi6+
6BnLNGs+j8xWYxpgrDhJbVOmTorVxxOGtNZGBCKUhtxc1pG3kE+CQEfzvSroihhZ4QmWSMEV2bjl
j6aPUlTjLapW7sSf/FwO+Rg4tOfU3RJ7blfhPOER9UCBKQ0BJJVtL7WgwvnJLc3FG+vZVxPa7zui
+65W2WJIPKHRlwQqGgWUcqwlEOkaYSHWcmB8ln/EOYYsprLOAYs1SfE8mpa8zBf24ogCWzxbUf6q
TyW/0iXI+YGpm+HOQGpv0HZuQBSlI7TMJWseO8t0/M8V1f1E/racclITDejjwbuQvk7DyYsh5PmN
tgDPTv4EIp6kJuTjgJ2j3YR/q4F3LY3qWcgw8rMOdELzNtlDHqAWISo0RZPJAeH7RZrb5HAZPnhl
/Hnr45Eti2we56XzVCKIEW7YvUqwH/Pu2PBpOR7GynXHpx73E425GN3bObcqXuCZxAnbRwGfl1My
qbIL6CYa+oRVt9XJbOsJxIeWj9jogZu+x7b0v/cDuemzR76brpw64FMrv0M9DjKAzztvGPAAVd9A
nsDx3RQqi6qruq0EE7qrqyrJ783zuRcLHythfpgWAwVAMT7qyGBcWzVO7TEqp+rtb4XmqXduEgY9
Fx/WIryFfKaZI5YXIbJ7a/dR+f8WDIuYqDbdEPPaXbNW5WSiqEIi2vClr1v6o+jXGCyW8PS0gdPD
dhLIWgHnm7JFN4Q0kq+huLAchMILTtVLZN+WJJIu9hpw4TV8iaWm99ZTBfAC+hXmUbFNZgwmy8xn
ovxbYPb8TrQ1RzkK6NH3gnRFw4decGMl03M5IjuOQDL1FvlbaiOXR1nuDPaME+3pGk0gErryvfqu
Yk8AJCL7mA/UZSWmPMFXkK+qagJ6bHJ6xNjbz2PvwgoNxazJgzXoGUgbaQS1xH1QkLCkXFx+5jt8
2xMYrT44lznHxIJ2XnJe/pr+jm54uKlxAvCtHr1GHSZj1IAG4HMi+7KLUClkvONy7W9NG2L3HbNb
cpKvotV/2H08P9S9135Ie3xE3typ6dYHpXoRhvSDpazLRFOK8J4w6duqR84Gyehd6Z6lva0kYV7b
kVa99pGLF5kYBlqojkMfKvfXAMfXLT6noKzsgU4hl0bEcoH7zmyzmZTQt1qqme0xm5GH1hAP7J7/
zxwG92VYSLG1pu60TZy6579iHZcAKtBp98TjH/9EpqR4/SWQTRBCHDZodVrNSnlesbdMoBh+zyKM
I/PWua2S/82ZEzC2A0w87Yi0PNjtxDfaqulHzV3awlhK5rn4eF773ueOPfgMsSZVw+M9G3iO4s+C
vOSB/olWZ6/+mV175BTxVciPQRYG3Fj40vsRrZiFSm6zJiKLCiw7aUk6PIaR2QFZNG33K7mk73MQ
a2I12TEXhEPdBH0LR6kr0ckpdpAYz1rQkWTw1XOTzaURwfZ+x4LlcPmJNkY7PQ6mh19/laCMu7Zj
RpyZS2o+vuYbgafrxnJ7nHszkvHsdIdzosVCmLWsg81m6BPm3AkNDT6G667BhaNt5ujFl8CDOVPG
FnjQsepqE2jB+IA6ycKw0aifYI+zjwJF0DdQ6LrkorScOpV29lYb9LRuUOVE9FzOJd/9BqoPt4Fc
LkhmS5KaYJz3D9Y1tsff9ePQPLUF/VsxXSv2uBNPywTB1n+c+HMiaODlAKJM1Piv16IXWz2nbpKB
DVmvTCNAMtwtzDq1hfVEUxp5/jbEOzuPSXrcJzwzHBon+dM1IG6q7+inCJjgt47eYqq8D7Q+sK3w
slPjdIrYzCfvm3vWoAPyErGKptGPH6zWj8ORdGckTc4ucAI3Z2FU1+VGTJgTV8bH3hyAgePzeaiT
HnGqRj7P76FBoLEaW0oTUacYZB3YnG8HhRo8PjrzDlvBsJ1UY79kIqldiqYYn+TwGELhTDpGKYq+
dkZgjpaJ5Tk3y75IRYQEib3eK8grzxzt2O3FZdph8KQYMYDkVDCUOMiN00x0am67ALLb/4249Gls
CrinsEAi2bR+okE+QHIhOj8EWUEs5i+H6qS8xwPNGJFXCtinOY6Nm02WrpZjI2SnYQwgN4WvWWOO
y6iYhd8bHFjzui77WuhDuZN19lRLfl7x1aYOXuTjAU1DIafwDjXdPRGpXVox5xK4doCr8LESWTd8
VSMeD0+UCOUm8klQffHEVLzM6A7SYC7o4PSAMzivp2apYuNM1CwCOz7T7Dy9B8pK+dAv8Aa4nPOe
9ZIWzifuAxf30hRZCPbsXYkGiFYEfyEpzmGw1s7I5jLSqBKfVtv0cMe6UkLG4EwfQtX804dcoLL5
IaMOPhtEBHduzp201wv2i496gYT00wa9fWE5ne9DJZsj4mKVId3xWYdhGq+HfwOUzMDtTyg+UA57
iQ0P7SYN6hPopkeLwwHLpwnNBGYgVfGuMmQNtrfw3oxOj7oMPYAqXdVPfYhYFT01PSpM7h9l3ZKr
sT0sRXEtH5TKOgGwvEPt0kziKFkPpRX8IBRMLyCUslPpwS5qLRWf6a1Iz98dX6ZR5u6MQH+mAP9J
X87/70YcAzY/w54oPo9equ0kN8QnzV7pYg2q1RkazHecXQZNP4c8awQZjJ8xE9rnnVrGzj8ppQWV
YMqrReTzhqqIdS6HrtoTFfEkgm56y+e7q4wlKhCJ45rnSsQ1MoUS3h1iFjWospPojnU+9wGLp1Tb
Hv168a3/I47zTgY/90pIADaKL8/IMxsKNVR0VxLzYj3vAzMAVmlYQpQBdVPErDVDGa3OyB4QKQo7
x3O3vngfSK0qy5GVWWns1xSr4gLBUi5bNsX2P6WJ5OzZzD6XOkJbUCKRiVu2
`protect end_protected

