

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
WOJX5Fv2S0CzprysR8KMEndET58Nnshq5G41sUF8nyr23cEOOYS3xFWHzDNrh0BglAkKcA2/EcsL
0Mi0zP+UFQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Gc0ueCwDN9OX/N8ZykP2NxXOhHr0aqi823TAFhXP2T3sZajOBosaRN5Om/T8R3LfwK7+baNKGGz+
UJk1ogy8JwdYWmJV85/JpyrrDFtvClJsQxdfCiEg0IVlJhvJlhs6FCZi5Rj8qwlvbn+/sc8hT0BX
IEC/9Hv+yH9f2HZIeiw=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
gOAtaUsYvJmoKivS2pd7kBeODY1Q4VX+agLZ2/SaxV/BkQgGuuCLHYg9eGdXBmjxTqXO35IrXGnw
8lzEMm8YS53SBgfLbyNKtLJ5Qej5jTli3Hhz2BXRqoQonahfpMOh6WT/32Mi5HxamPl3+Ad8Dyj3
AbqGosJ8LBJRb65Babsp/E0dGGngj0nJjmmY8NHpqNTG489434uBxC5ykK4ltOheXkVJtXSHoR2s
c+RXEPDO94CZYlHnY9b3pUqLafSVqXTeYuw//0PIJQNmrXYuvkdozgm129vQnlKXVGzYsK5DUlRz
Q+VO09C3aal1Ga70326sWIG6XdhCFEnAfQoucQ==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
3INKfUgfMTydNk3PjPUP24H0r2p1C85cOfDxce4LgEKtine/HDrFDahWRWORtm3mNUVaknW/GXSC
5KErdi7NyQ5+CFdf2MMmaC9h7nGYKW8O4nbf09hLlm3blRBSd2i3h46PihYy7iaS3Q+Z7JKvWuiD
J79EKDKw4Kqn3mmg3iQ=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
YHV/PdEXZA1kC+N7hsk5uDSJPgfJRc2Sgeu6l1dsNtZhWFmXeBe9vCszID1P11I6wOICxCc/uQgT
A2JL79m9I3kuY9Ji47hSGH6+xG4kfTKsYaTVdl+16SjuG/YaIhBwQfN13p/8IGQ6FysnYNYR5siA
+0Lm6CwAYBXVRwsuIA3R9dSPKgq+Sbk3MQCuaqKXbxHiA5oAAI2R3Gz78f9hrvy4Cj5P6dJ+TbkJ
j9bOdpZE4W6tXHasCVI4EqJlfqQQ48uWK076fFPDGpd19w+K6NBgkvxxlXDC1t90ZvbdFgDD30L/
SOFjS0BafCCf2aKaRk8VIdeBs9pr4wj9gMwZYw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 12496)
`protect data_block
o8nOzlNksMfrz2RkUYX1YyaSce+36qw5/njbWXzJ5+V7nYKED6feFJTdw7Tnv+ih3LxFpl+XAIvz
JjORTieiRmO+due2ie72KWJ9NHl9CbDMraLiz7kblBdMldJY+ascg6cLY0w4wDzJNTU4V3yJ7WLt
UPAmCa3UGrtKKhKDumVcIkGKFMpOoCEPCQzbJI3LTdfvaWIKGxFqVPZOOYkuXcl8Byfnloji4RDQ
DSuJbG22W41OfPoYTCx7/IO2hKbd2sMi5um161s+KDMjtBXeXKv+pyNRmOxTg7IbWZ2dtH9Pv51Y
5YlXwGLKmMdcb+AWZ2cwo8lN2s+x3DhtU59qBB/i2hRlC8tlWxapJGbcnja5FshqX03Yz3jJByoF
Fc9UomQNNs9dwhr7Ns9pps+dAvzEWNAE3dw/GUpu3Z1dhfMxnKeG5tDeXeJ9okNU/xzv7DWoUPN5
wmR2qVxJX9H9hF98D4Y5Y6bak3xSlvs71Ay2lJynFv/tYEZeM8ptBwogqFOzLoZsYS/gzraZIot9
/pB+/OdbRJR3oN4Ptz8i0I+7Yy452f781nfHgSE/HBFazRskHJVcQxhNCx4z3hqjE1JNoswarkAp
uxMf9HrEt13aVYtkHh17XWKFQLb9fxO2/K4/uBFIVOb1vFgClAWPH/WeS91/runNTPXxVhjY4z/f
on4/EfQC3ozqIRLGb+wRwQyekICQDLg3rZxyfL+NZN0Z3N+3j6fkJLt/ck4mu6JaWixKnPjjhcrN
0lF1uHKBpQMIW/kPSYAefNiWNNmnw9/OUAGQ1dsmWyLsH6ISyGX7YZVYqWtvsGZGfzzDnBr1wQbO
4oEkLEO/B8mQCnKdPLdpHdqVuj2Mz7k1v6OoHlqgj3IyXv6cKIItfg0HXf2uCwltH2igCAL4EQSi
p/0fgG/EdFXx98isUHI/9WEx+fRtnt1fv+YxSCmPtJetnAhkZAionbX1Fo56PWjy2Gm1ggs6RJT5
v44EDXcZ52FojUkzVG9w7AsHsp47otgipcIIOSI8jhuQFSTI5lANdJ6U+A02L260ATAkaH/jVoVf
FKys/1syOAiiHc+P/WLfs1Yu0JOiKsneT5CnT5Xz9E2tedyiBpe4BG+vnpm52SrPuzTYb09SC7KD
MQbAQOculWUAwiThXV4RW+QY2Evm+X84uQnWajOeqkLa/aUVIGgdxtwKiU0yR362DEgvu9XfLZ64
W7EBjcnPvcfQMRPhtyiaJrQRij5TW9/2SrniUnfNW8w3PUN05Vc2go2Ssy3VtW1ect2Ab99yDB4O
fb4DgUvuIvEVsHNhjT9LRYy+5n2x9Gwi6DU1ZUGSoemqTCmKsxZsFxPrlFJ4DFZONY2sByc95iv6
UdJRn06p1ofvr3ki/lnLZ5bDUh05UGrj6Yo7By7jCo6VK4HL/bN/o7AKrsCNxWYoy6a5xueQd3i8
QSCEg35ufkXJfrIK/sbc7H0y08wFXDrYzs5I6Rw9xY0UDiT6yNNGNCKCP8We9M6ANCe/7pxr1k2X
fhX5aIRxHU0vI5UJ/YmV/AEMGTddHYRtCpAT7BijiUoF3dEOAXhJv+cHoEn8gB59HfnRrhRumwjI
Pw04jOq35FUeKuIiZYF+BAfaZFbl6ezABJjQkpz9BPfq9kvl+Av/nb9t3YDK7cATDElR6vAXBXBu
dxJutKjn9n5Kvrf0HXrZBqQfRL9lYZP/bUQlkeNeZXWNI1N1ej1QYYy1Gw2K/O432GfBmRUId4IP
97NU4+gZkSApDjtRMd63R+n3LlOxCMHSL+Gw3bozG5uTh4FswPWB54snPedZuFgbJQZXVkHu64tc
0TDbjwTmkZSeYr7B81UJaper7PCeerDpEf15TzWRTTYknyw9l/td43sHcdomB5GBZNdg1XFlSoTD
r2TwwftIJ8u4Mkk6mPVjTfQvmxBaqj1DICVKUvcP86+WTIHQrltolayBP90p4NW/wfM9/EVBSfOQ
otghaGBRE5hiOsZVCR/R4hs/4SQdve4+3Irfhz8LNHeu3nphK2wGYCrSXVztXVZIHC5R7liSC2zB
tDGWXvIjnOLpHu5cFeGQcq8s/V5CKovQqQmiIjx+nuaDwtq4p+Pc2Rtkkpm4QM/wX9PRVLFzbJyY
muflguHXAU8bny0VFbm52n9YZWhPIFFBkOiHxnQP5A+5PvoTD0GvwyOqj8SCniuJszfB3fFbnww9
2gdKHogjYGZMGvS43v26kWSzYobM4oNS0YWKvdVklWctYcOv2MONkf4WKtgWZ6iHxd09jx4NKhQg
/0Z3DjBeXB+2lf9fuwiWo9AZZaMiUGYnHj7DvBRD058K9n/yhm0VYL+5qMjxbBVO6N9b7C+bSeNK
1HIdTqSa6/Hq319XAnitIIjeo36F/RenozUT9fs4PqtGg4UQ292ns/hrJ2WraTddxQFxheQPhG2J
gr/6SF2hx81x1UB4N4bcy37KeYHOIIkqh39X6nzZLEFt/vjOrEymlIcfmRKUmp2aZigKoOhCLtL6
6ZYwKDcyifF0JNAClK7xSlQrkLRqh6B+qERzEgQvToeJt2XLdE43R9+m2tO9rpzaVGwVGVbq106Y
nKs97OOzB6PUedJ1+GDkxJvRCj84VlDymZAGbZRTKjoorP1aD4CvRDKFQmSj38hMIHuk8YZmLGFo
L/+8X2Yk+f3kH+gj9tqy4EZuc18isNdVPaabGJkWFFsmhPYRZCPuWv/3DT9tF/9ydD/WSdlB2PC+
P999laWxPJ7uRbwtWF+07I77iAGNNbVYzD+zRXiGWIb+ryRaZUC3hKxW5ZkoUVigj1q7lpo+arxd
VvoWPK9VVqF0NHwHxKdnAzX7n+5CCgWZfOQWnWjVrAiwLN+NgKb3/uH0i46ty8BcPsm/P8dluNVk
omzP9NT1gbhXWiff3UQjK8/NT+SdSsHriBSq4AIE552KI0uwx0DPOIqxBqRKAK73xgnq71uLDvHt
ZbXzrFEywy0/+Z8gnAEOLyDlmuZQj8CaLbr5hnX8Yrh7HZyZ3Lz2RJPrYoGzW44XiEHP+DS64WD9
MX1jPbN7hvQsMk9zS8N8xtZ6m1ui9569fcDQjN8VHgGAips/f1squdsadH+xoOKUwVEs3z0g8ygW
lgUWbOeD/Y3wtjWfhpjdNrsF6Wyhoh3RBuzsJzlsHyimOV8qPsnLYes/XbX1xFL+tqD6Lxn3acSx
SFA3iFJQNXfnAhh3HHUdrDszpQcSpmqWht+PMCBXecCv0pDaSINZh7rwwhCL3JVCVFulCNJMQww0
etlOF1Y7/sKNayXzLis5YW7jFgdSkF7paXoJVeVoCf8QPKXho9/2o4fmHtwR75BslxlfXNPVXTAP
ACiviquu+6mGRoF/ZAZX2taqaON+l9khaKemGOfVfeC56L5dyJNGqnfpp0xfvtoTwckY312wSj6o
0qboWskGVf/hfnhTFbUXwPioS0S3/by8Jn3Ocl46598LYSY2fDU0CP1/smH7K8Zw4wuKBcO9v8h7
1cG7UBHrQGCYoAKJBmY/euQL617g+EIB/LJrrzYc6QKEpk5nf917rt7luEJXKU3XHClrHzmsReY2
Bm1wYmDCUPKMoaBrkRCD1aKjAaIyOu03fwiZ8QUAFEEfTsL2CiqTfHhMQAqgN6ahBLDYmBuVQ//V
RPCjnDevmHsrdX18JDrRClq7iupacBTGms+ouxrGXMx2xOtJDuMYm2lZmi1YUHLpl8mWIAIa9aJc
ZZrhhNO0i5IsWYyzq4dubZIXXXzKOQf6RNNjl/wTCj2xD9yKV0CCHfQaq0rVV/PLPPuMVwdL41xo
dAFJh41Jekjdok4yxew1Nu2EJ8rn+ouBuKhYZtTN4b4QhMc13FgL1pv59olAVSgMtSYZs/yh++sA
hW+NB+BaIpwwPOnFSBfI5uKhmfUC2slMFIxl3vDt6lBLuVjNXKiAokpRNQLISUomJ1sZbIr4e/Ab
hkQB+uXnctuIpMKDaa8jbBJzCAVfdXpgeiI0GI9z+KvDWF+tZEqPYzJXro2gtmb2oKWZptnKJthl
ZU4zGGmN/zzeidC/zzYHsEjJOZ3tliGgnckEDLOKiE3ZKMWsxfBJqO9pfn2Hsd20j7xMvUTIfYm4
iDQN0WiCYl3TewEZniO6BpYpf58cI3jTD1RHMWWnD/8ULwI5hHssYKqhGHlFMGXZE2/kJ0cik1o0
hPkciqKQdIK+nwgQvlcTV82i/xsb3OThy4HJAvPQpj8yEdIx2Mb27Vm3/k93oli62iJTs7VU+Kdu
RpGC9gLFtlWYR0DbzkalUEUjMKVDIW7qTSVtbgNv4mqBiu4Bq1LaIYgS+UxZUqlE8I7EzKJA/Q5x
OSvKlZczsoDNw1U34D8RB18AtjsmlG1witcW2kI5JYG+Dld1bEn+hDeQYVYSdKpFI7V/vdqToOIe
vGJUCagjtS7G4mLTQdSMfdFdUYgmjEtcTOR16enXuHDVnrL+o0kiTURAiOUaeNRfiCG47HKLoyLm
kuFpSJM8OaQDzbNBkF9p36QCtWP8uk5ap0hIz8jQ6FMu4pv2/OyJbOFj3lp53vqa+psOLMpUDTMQ
n4wqwvfFXqTPaZkvRlLNhUNbZUIatz60QRDgU+wfaLU/zcDRnFFH9YQcgvOoO82yOxB8S+Qyo9vj
B7oXV0veDx87YDtomoIlxGE1CC0RVQgnTqGAyzeu/AJPgjVZOxB+95Kekda9TNIXGQMEzMk1mqsB
KKDXtxjnyxpsiT7dMwH9Ar84utMfskGvbe2q8tV1ooF49LPsZishHKcmE8aHJIpH3Mlrj/oZPih0
UySGKzwShSBj/zGcIB+RzdDFJSF/zOSAz2mfNOnUtFk/LOv5g1mGu4WSkeZUh4Oxdl2UgEjjlyH7
45Fp+8kfk0+KgF/x/VfxgOqKQV4XGOw313CWl+g5u+qEMzVyqCuQkDV1AnwjJ3DTzON1erAoYqPo
AhGUUj+5+hAG5EPUX17pnZWOmG0mgak97ZZS9g1FphZ/vFJFoO9pFoqtgNY6VcvqdPC4DTnd4T1M
Tti3LO3mTSg0F1yUp2mOJdVu72BE9dN2r1Xo02eEZnpXVRake7ltOMg0wl9LkPMI5txeCp3sTDI9
aCujESRETxZbwevaj19Q6Sk8sdtMD/SoVcZkLYI9Ht4LDoVwqJ/AljuVgsQTB3lPPyy6FjwzBXDq
Au8qOAHkBPN0z1tNNfNmBSWl+hSkqBmZgCqTjd2CKziH2s4yqUKx+DcIhjp5jJKsfvxefWzYDfZu
LFxzTNWk4lPi7bKyHMg5FmdFl9bb4RzdmF0O97pnQOhhB3txfdStZ1NArEp6pnIrd+VDmgw1ogSC
gv1zl8+wP3II3NrVhbWENNkDOGpMaPlgzidOYIRrVxrK/mSHADilaDM75aZ5l0E6Ib2GsOaFHvWd
PH2zl7cZcUr/hnCysxQWYs4n7WfnhWEtXk20e3914XA4TQEgk8BpJvomKGGJO1ItO/pUXEwoAMCU
RUv/hNdhs9ZOlRCifhh49YmWmnj9i4Ba4BVEInb2ycH2FoEYSaGSYe/9dAZJkHeYPjHXqrVz7EPp
RjfoHVO7a9jBEAI1AKQIHs1lEE4Ym6bE6dvHiW8wpe70dbRy3DgkmEQrS7zTg+NrSfWjCW9DnFip
FuTYKxPJAONTsY8yjkackLzdeqw8z7fMWauk/nnAIFPIzLHaGOnK3ugVbBdZs0oPSK4/zI4eCEGb
loafWqZlujQ8J+WHBzIVC4HlxO0g6hvwmsAjny9Gvd9wkjM/DDzxJmUcoO7ILnGVqOLjeJ+O5woJ
A2zQDoaqQKYpM3oiY3rqS4uyacWspJ8HSudfsiVwaiCrZMYtE7kfwItlMtn/0sv/Hgi1kxaP1ie3
nOmmIWo4hmnaAT+sPV4J+rXttfrPOV0aVOp3yDDPk2L+7AFwJpNkazRTicurRnu2oXcD9V39Tjxz
N0FCbUaRNj6UgAeKDMH48n1UvQf/OWaEGJpYFNU9/8zBTuysoT4gdR9aEujLmM3dhex3zCThWeXz
+S33+DSGYb3KXwQq/LY/xfNONouqmn0+JqkbyX5MLovdREvKZAmuNYasSY1juvmeiAw8S6rYMgAm
1PAum+lSvqAaHfQW1qh6uv09xLQn6rol3X7xQy3HCOB6QW4u6bdLRfNZYla9WuhCIVuhHlmluhk/
8vIqnHNnz32VUYS/c0CNXg3XYaooFsZb+2jS7Hb5ZSLwyEq7X1bEZUySpi/ts8EV9Bu9xONqCnRw
aEtsXAH16tebrNAXNEYKtaCpOh5oK6Yjd4zCrMwcQH4H3CHD7XWLHqtq667MaItbZVAizIV+BH8Z
f83L2vVLdErPzzrVpLhcOlm7ja406pz36RxzCQSeUMORHw9XZHn8fBsxhnJrJ9jobW2SL7KFwsgw
8WrQ7FW8+/2tLAvstR/6JsGVMjKTbQBmCCuKuPuT2dCH/TY+3zc1q3x4kvEeZBM54KHnjs734wS/
Q3LT8zhYWuTBavEKPWJvH2OSnqDYgp7dzPTlQ8999OjQQwmV4PM1pwC0OjBJMKAZenu6iXHjeP/Y
kTvWenQlBMM2pFMYT+SEUqpZCMCnIl+kimnR0lTU/IDHPA5sCjBCxoOotyWPafRg7DIg55ihgNfo
t2975Xdq3x5WzPzx+so5nhLIBQPEjqkSiDp5TYz82A9BS9xCXWlCibUdey6n3o9qg8sHS16lUpta
RdI5P5c1GalVoGswMj159mefouDEGnpGL/iA7q3QZvyT/FwJZhpZfVcJGgwoj4XB6DQTIVZQ6JyM
L7Afwfh51EbIkaJbgwVH4LuPCdAU+FffDr25BsrZxu6PEHwUXmaoiiX/G105Ye5u2b7jF+E8yLoA
V9KhwjBoitNARuwczz6cOcJ7RtYfiUunJ/zAXNnDdLnkP3wtA4VaamnU+3eMtagRmbS8Xe9+bARh
QFMTujnpFbfEAG7O8S0KdYkqg2PBaA5IvaFBSXssiAKtpvxbMEYO4io2Ro/ib7KO/UHJk7Pk1C/p
pAgbTHG278GcdAk2BLm3ar1+i9dd7lx4gjNktTczQ6F2LTfkUfkN5z2SPADe2vTG0AghpHZ6RwtD
K9LzFMaK7Fjurt3IZPMcTNmkFJbikGoH7hHLC0JXJ5fEYLApvgo6wLDIN6PJbi7Ug+1hMfnPm0ZG
umuQKa3nSUbCFLm+zRek0cIPIEvdSjsX8Teop7tY8Z7W4iEG6zWYwc92L5BmsR0n8orqYOU7bXYx
ojXknpncki8ttt0JtRzOaAvYRhjmjPU0G3KCHgk5rznnUk3KXwnONfO2dCVSX94RTX58CeG79wmh
DhT9kJnxf3si9iLhIpo0INqJz96pSSf50HXYneC7apKnH9wdJJYu/+NJg4K5QPBKH012igWyRalN
E1OWadX5yipozF72FqbJ0URPL5/PDil1InGRuoyTEKHPXAAPrgKrKxdsqaIU8GKzgjrr6+P/hYkE
xuq1juetBmr/GSIr/exT2BUwoQ9DXVK81aPnEf/I6TCpamp7ulQiSSVb1dteRStLH49cPOseV+C9
YzgtwawMSjTLp6yb2AkgN+Jo3IcapyKz3LfYwB0pGxZ7ooGhfxiSayiNnDsLWQYwX1EYAhiYVv8B
Y6mT3TOUITk7AyDkxO3mneFywttJp23dNPjpZrEQEX9+gDTlQdiLfUZOpke9vHoNYsAm7JZgdo27
xKH8YFX3CjdV2NCDumHiTcpY30INo22gFusciTn7qViTeUAYyBRNY+8GhUXD4akG249WDx86HguB
pQZjnbhBPcZo9YGg8961DY3NbV4oowzcL6DVE19+uoY0BZsbTSpvHeAmq6CTBWkVE9UA7lPZ2xpo
s68Hb0RtuWPxKSvMRPZiy6UQPr93SnfkwysMjMA0DlKxEsvtY1V0Vvo2WINGCu9aD+r5k1kvAVjP
bfesIR0IwVKnMzHvvFMsrjCWjKdFCE8mujCjZ/NB0078OUjTZfHR4hZUqSpgQoMbtHsUoEsUtNQW
PNpE+fsMdZr9WgtjMIR1y97bNkuTBzVATOV3dKcLV9CzM/js/+s2n0tgw9H/4iqCy5EGFmWsaDLe
J2LiGqsi+2J2W9Fm9ZzWtkrteRjEdiVhgx01NDSH+rC9bYz7cD0yjwpcgpW1Ywes5kRaagnRBXg8
YrBtRL6lax410BU9aNLFBTZAHJ8JRuqk806//Pq1YkTdDVNOJh4/n+myQa1jHJ/hRCkPkd2kcqMU
SIYGnxD3BOAqpDHFZXfCIxehzB4QJh91kfAkomH/w8v+191KByvc/5HCXGL9OfNhlP14CNWikrNy
6PCPlPg76LTploNWQyn4E0fo9CeSPlDDVc4BBPKVcPN4TXscWPtpthaPFA6+kHTQbtmkcJ51F3kP
SoIPQxHBBIWgG76x0oI5k993VaLGakHKe0UvFPrNXYYZKuYm0HiVSjC2eFbtQAw1rMLFDrkEvpM0
6ai1qqhQS0+Ol8pHK6YflW/GrSgBkZkL4MkCObUGcq1TlxLQnd8BVtdN+HPOfJHgEyh/qR38IIIM
ZagT+31c9cfYtinCHuPhi9h+Vs+64A/R855YLWtQjjwX3gYIovgOlKKo3Pgvao0RmoM0JKrfIJyF
GOGv0bfvFfWEXyVm/YCuNKBCY/7pZylJWWmESoG9NqCtxKvsQHY1rKEo3lEEok1VVbcE2JQDCpSF
dRv/qeEuxinRi7181pmiY29XoBMqIFKzfZzxhoYPghwAYONLr9Xz6tBaqUz0qoXnWRrZupZJ2e9L
skqc7GOWTyPROgi2eYczijVzFYPwmTNbJyjLu7yGQw/qpJMkmf3zSV824fNsWWuNVcRPpPOJPMw2
+AG4phU6K8AvURqVTSs1o/0y/E0W1l7A6jlVgYOpOGisDcS5eipaQfmH1wQm0TXYcWnsCIOC501f
rehb1fIuand94QRP178JguP0xXILnA9bhjvss0lD7EOqPfXfwq+3I+F/gSRnof/vcbeY9PhUWjIF
cQhUdp//R7/AXrxaNAuemd0Dk0uLmKxUdeIMHAolvCAB2s493zTxMZ2QzfqyzAxIidUJpZjH1nGy
IeUh+tpCP3FpSXBJXyq0J6Au1Shp3jJJdvsSTnb/fxvjPhPNhBobPrIyCI2UVQlaTFaX4jXWB/HS
p1eTTNNwVXk4TPZZmpo4BFGiRIpuJQrE/zKLMo/nE4PEedh/+iZoMBrpEx/o9dJLIlRPlEh+0Ke+
j6T+F3sfp9lCCp6nZ/7pVRqbIW9Cw+uKwgEUU+ClZmHGAgd5n5ELaq/d0fQNj385uEgPzOzWxkcp
8D0S7W4wHq6jC7RMrxQfP9DZwC7Y6zm/DSNAZtQb2QNP0QYi6Lzp9sBQGIpAOR50ghpMgNiOi0ek
pHB6PHngMjPRWdKIsc71+NhgOE3NuwppNdGY4u1o4swnmjEdh+fdQK6H3JMKaKshr+QYJkU8eKdL
RUmwYoP40khd1vwP/saLkw3DhdEApHi+8+Gk9OHaxnr8Q70+MUhTOhraHGcrKoXPzWEEf1SA+PHW
HPcCxinaIHW3xWa5DoiSl3+EEPnPecxh0K873rmzO+MZNPV1BMTQvSe2vjOFIOyxQOF6zrcdgf8E
jn5jGqHwzLnWJS7fIwiYr7xpjSp13W2JeIX0gQihUwpZZ0cMti94291jC+Wm2So9lfK07WXAMxQO
BXjiEhrFZo2vTxemSKIpzzCjG8yCZXRd2Y46LwNJUCdfPv58Xvma/vk4MsQyV2MyUP4DnLtgV1Im
PEC3yLQXm7QDzGvDYWHe9E12r4uCaPfsPDXtsJPhrghrvr7Nwwskw9+FhNPJdQ4fmPSrvT5vh9Jn
B2A3AAXfYqUloUNsGOAOdyO+WCA+YYiB0Qxt0VY3FHC53d8gmAIHqwQuZb7yBLxL08BxlyUUGuRn
WJ/8gpvr7rFRzbnqH+kLBWME4aEswROYSJyPBpyQAA8/qkLif2xAxAhM0iYDumq702pPc1rXNUmS
lH9950yj+bdUXmlkaL2SdqdD7cqgLRvMDnhskW9OwfNx6UXNY1ft34Ym2dGp4ZwhrP4P/NxkkW4S
7ar4sa8vnahf7mDqQCckXwPtK0jKLLMNhMe5iCRvUrjCH2BnjBmqZRdZcn93lYHa+3S3Yo81gFc1
ro7FhTgNLTJ2a7y3XW5EhN71k6a4UCfu6jILEsdms5jjPSuuSjsLj4sQpfdnroMBRVZwiWmW873X
Y1KaSutQdKf8WY28R9T8YOmAwd0mu5Hj+BP1DL0lZbNxftG7kCkMg3oaiOdUYkYa624HWxDVvr3d
t63biQi115Cnlw6WsmQUTVH65O30S92f2FPUqMDLPZ8ChwUm0ksMA3q9PVIGKngemmLJQIK8YSHs
PaOt3enMjhk3qwen+s3dNx19R9MIsp7GHeBNPmF3+TAqswQfllRprG6JD9esI+6GN/M6JOksP2BE
IOT5Ny2J/51NGk7nqCoSwI267Bbr6TQoPxPUNR+tl477qjCzys75+celv7U8l59a7gWazPeg88/v
izuAlGnCO8iw/gu2wcS10bA4nzB4NSfqyAxuiCl7Gk7I2yF2YQWoWHOQFn9pkSklsVdsbIl8xfGC
cq0Z2/pfffQGPZ0sdNl1QREeAMHXKnKecw5kpGS1R58bxgX/AMp/zchqUg6Y26dTo8LDaOhq7Om/
VCQeaTtb3OiJxEWN+73/Jc0IjATHaFOo+klfN4nOg9IrbX8nttvWvI2W6NdJn/ezS2aO8Clx35ZT
qKFerrHTOYpEcKKudzNfYm65mAiMc8OPc1jzMwOj93LXQAVMxlT+WMun/MY2pm+WoaMySA6MR3t3
uVaB4vY/ou2XU5LKMzEqyorP/QgDVBmQ/gN0NO3MW0OpUcGBcP+1CnyZ+9Syi4KJ0vUocVWnmlls
SOCo8mr0LLgT2jgIv5AKpSGwULzV8CSlyqmhhvgrguOGdQqDnJo4g2xq5ubICVx0E4vMJ9MSiwmo
+5wlTYbZLNd5sQFgOfy//pCdJ/6NnjchcM+rhqDFZjGWLZX1nmRVCXNnXntxO47FSXyK5OEQvJLK
uEXwOmTWx06tLX/4+37amQyyr1Lx5C2wAFBl01VhvBeAIZO4h3/lHdqlMcVC2TFC3EdzHlfBvYn2
nkUkGjpxhBJPylk/zO3eAgDPZtyM9fVGZSbCivdTiaMSleriu+IxnMREVFtcdKoyfoofK298IMC/
RIJBWZWqFENzmWRHBngrxJeLvzv46VRG0OoL+rS9hstxPtOk0SeAnX+gpAlUwFAM6SDsfRAhvhZw
u9xBLO1x8RAAjVhko4B/evvbJl3lJ0n9B/rDipmBe1Xcg8xAo5QJx0QE31p4TY97wDHGTABdi/Ac
IVuwDd1EnyDLxPKWiEHK2zYlaoYNimO8gO0cPwtpEMSAw1j+8X8zTybMTJnrXdKZzRv6Zfoux5Ja
LJipP/o2c4SlpkiRVPs8kwXXSC0+DSvnFHj5TBuddR5abwzKRPkXkc2sxNiuJX/usVuXbAyEG85Z
30wG5UhWBppFvs4z3j1zSoXTCKW6KuwssCy1TLYRdRBjasTUlfyht2iln6nhh1kC2btjzbV3iVZb
eRoNS0vH/K0HTD+0LbpkYM6568LHePF2ahbn/xSiAU6SiWBewXhjGqc/LLsi9mNXUuLrHGg5oKqc
6L2uxLk5tDPQxez38yFbw1JCtmhI9b3X29It3SqVvcY6R6XZUCXq4nBOhOHtnkZGeDRMvwL+290H
rePUNnWI6O4mrf9rQbrf4Wu8Zu/hTafoS2S7ilLiitwCOvn3U5FPxEJYk3w7/wefTZINiWqTs++w
jEGWyvBUrUpDx+SkORMxLVaFZc8XX4TM651vfumXWEyt8jd4HC0yFCZaHM3oHd50swfn+Vv5bDrl
0QjI9mk+/GW5nJ1N17s/iLHlGXK+K68WfqItLW+uPgHrSKA9NZciwhdkngiMD8V4Kb85km5ZdLfw
JuF8zmGwCM3gIjpNvvBxEqAfRz+RElrl5BjRaTygWRXDVymVbVyRf4tjA/6oObJ4hAjXBF4b3vvw
lxxsoZrWrV51uqzkOh4QRr0LNGBsHKVH7jWhYg+LwjphPmrl5991ttH+ufXvqk7GQkxk0AqCyA7i
8mLRq1zmpXVj5f5rN6z5QXwU3Zots2GS42h53w3HvovuVyMg327FzrsWbjpfgnpw3D7O1S7ntxiv
KH/XD3btj5Zm+r1jOdBioeai+1ahHwY5lLT8fYPlcUV3mMNo8qDko5ZsFFsJBIU8wg/6vj2nXXwc
BZGIFSoZsLUUvbF6Giql1T2jTcBtBHITqVH+IHFniC9Exv9WLJ3fgSNHAZAyt+ohFKfUwZg7qRgP
dx2lTL5d+rJvSwtdgDOVmEYvoQzfnywcBVkohYgENX4wGTW0Z8i64Ld4dLwZekEebelVjoFCQb/P
Ibm9ecNv8CEqm6Imxixi956mK5G0D8Q/cxyUy7sKI0H0mh240Rq8QzOCJI15O8MI57f0GcnN7ruV
JXchMiusmnK5wtfrwe92z39gJqT1ZPuNplRiEnpKEh5xD1jUnfo1fcvEB6znwu6byyK9j5K6gTJX
xbEVCV4wIQ517pH28v7MgAgoeBi8tkA3b/IpdgcZ7eg6TbBOqKOLSro6EGqkC2NJ/pEnK/4jCyG5
N8RvPSjE8eRnEU2NI4i7lhBHD3sLK5o84syeJZqVdS6oQ7gtZOvinT1PgUVdRq4yqo39zssN287s
kYz7xztRkzQQfn/iCGKpm3cuRk0kyaRKUk+RqtjhJwIjWtV0pNup/9AlD0LkxXONQM/53jvtmnyU
p/l/aum4DJFbgyJtgrxY8anDDdqHsi3pX7QR1o8ortlbseKuDGe/xCHElNCY1uLZTW08MF27gj66
WP65M4hWPc4UqFbzRczpERBZ2EAiIfrfroqIiFqmYEmLBfV3iEFsqjrTUOxlUFCjAOekL0+dm9lY
U6Jd8Z8axJjvitvadFGTlUi1VyQcsYLAxjw6qrJ+h1dDOUKvZRwbzboJfhvN4k/wfo3efM3dgeoE
G+PH0tHHUoU3j+gKUaJBpcFOSzbWjkw1Q/cVPozQhauvOtFqndZKggO9m8WaoeIRnEF5ozaBE98V
4T0AzRxuisIk3bKPBo63+wf+E1YFXlmrQ58xpEpOEysOQ0RCawZ11cxY0XZ0dDTJFKD/0FoueipK
MbGcT3ldQvBHaAmOBzLFgYRBkPYpQQ2smA7Bp4szRaKNWzgP2SXJCL5EBPy5PKHFPkGZ2RuX1y+U
Rul13dt+9wwdWbCESmOkH/nshErBuTXbfCqs+T6CBpEqnlytYyalmlIeyhukVhdZ9m4ZKL5Qrg4i
68+AY+6soCtNSUt5IJMz2ywdMEHferovAizSG1WC1x/5ytLKL9V7C7WXigEpMwc5hoRA303oPWc/
ZdvB2oKMmdXp9S5nN9vN9x4kVaDJrLk9s/BzGBd5TESe08rLkK3unPHpW4Z1S0FRaYTdoXrVnFug
AURlDifznrCtWYXXpt4KIt6ba1g86VIR2OZ/+2FC2qeivfj2BJ2t/4vsHX0UE4lg9bSNvNGFOHB2
5jDVjbUuRQNuz6VaqKsOBFJ4iIQQ9iQ8DkYcj2EY3PFwiQdpsD5hFGysbhjK0i5KYDioiRp2QZKl
0VavWYAhEzQoMGiyL6B426dvIsroZKNXhImbFW580LxWGnHuLm52CmZH58IHqo/xd6SX5xyl9Sd6
YDxv1mlyxQBldfT7aUNMqBWhjmoio0hlcxc9ycZbLz4nOVmTTWS2vBdc8ZYytP+A5Pn7aOFyw2wu
4QNRNYiRS/p+OmSXNaJoyZ+7bzQFWyjSoSRN2u7XCASXGGmGBv03MEqpNOH51WKP0l1Ndu4SbUSw
ZYMq4L8s8m1YtgxwHlw0WGGMHIHOqh+CgfvDlahIBkppSKBwYYJ7/ULByOVp8kv42biohKc92B4q
l6pHSO7ox7ba+pZcQdDAmcycBxmjcCmki2uC2K75Thxn/VefLF9Y5BLkk9pthKopcDgCkn+TzoDI
WKN7DDN+4RuC93Y0fAvV27NCTCKbQ6PRNCDBGmmI06l8ScbK1ppor1iPGaB4DqwFX1G36pIKWQpg
Flh0W5DF7ikrWC3EBEEnOBstGLERSOmNUCeVQ9bRLSVptXt9bZ2WJo9STYe+DcD1jfiQchdrTvds
Tl4Pn7MAGyFkXOXaoPd1YgZDo59UGMJafE/GPOfsNeoVh5VYdmcJmqedkt4yPce8Rql3t+IYSxZv
SYv8wt1vwWxZvMFOcH9LBVvrZhatiG+0jjijnrtX7DsxC8FIMy2iEOv6bGDeYopc6i/NsGB1IXxm
tcMdLznamtA9TpUgmZcu6mjaaFcb9WpMmmc0X6IVq8mnDOCk1/E+djotOKcdkY3u5zZ7uh9taagw
5xYLe4nR/R02cCj1P5r3mQwNSyijUbd9nJC1VePHqdK8gmwhrMroDEupYPdHJ6pi6lufGER7m1IK
u+JWZZjxxHdJFnafqskK5PXrXjI5jRp08gamA7hB+wsFUBBHi0WGwS2ajz7mrYEYwyxMYxCvmULh
AeYqj7ykKxECfu7n39+4f4b2S1qcTRNF8pc2HdWd4Bl/SVu6p+SJnlYMD4hEOC7UlzF6yLTSV9CN
xkEBlKUz5GOu7s6Lv3JkhADddkBV0Y6esP66GNjfrGBezoSUzsmo0V5Y3YIddjLO870nks5sMRR3
a9DMJJ0EeeDSbUu30jGym3+6iaThfAsQ72GdMtkbvGJVNjSNyWnzfYtQJeEU4EJnubNzgdjd/mhu
U4yHw6/s14OVhOHMnLUs4T8JQVObSyD1qH7olkKDrZw/ujt7KCclUu3ZHLMQssj3dhXSkMMOE48X
N8t/xL/xE4Z6E/CV3zG4UkXTSARjSHIz0pRrzKd8/PZ1z1wQKEYPQZO7MkOP3WxSZsWb78pHPQXQ
4EvjRmE607uSa0aNuZp3HBESTPacFLPlhDHG+p2wBFXYPeG0BHJ8bhHEc6KZiGyf3mZ6dsBrKU+a
nrZFHUyDUM1WEpA5xwN91rA3CVA2a47y8yW8wJB0z7b61Jc+FLOj2gfnp32C9E3aEpcN/8dGlM7w
SWvDMicfAKT7PleRdqpLYuDBvXviDmyH3zUfiXBeLa+N69YgT/3+JMKM1tRlvDWO0iOxxfeTAOxc
n3ij+yj5qKZSW4ADflwK6YJjUEjHU818DNtIz6uggxUplVBg4qx1b2OgqsHngDhPy1XlutZUdMtX
UnP0BWoFlkm0qHoZE7LSiQsKoHoRLEJi3u9Z9tipmSfYOUtku1X1WGHyd4uktTX/dyt476SFT/nP
MCWWqp2/AvuffufWEcVSkdIHGUec8bbVNAUGcEvO11YC0oJENtWMfWcVErHOw4fc77PSy5IEh1Ie
fNOFWmp62QikvlIulc7+VxAykrDEVryslo8nUeslU+fGkF//L0hJiovKPNa2DQ0jecClhBjqzBjI
NrccwyX1sdEnfyxjVog++wm4VwElcnfSMxAIeZha2AGmAiR8O3RhYJvIqa5iWOw9cGDfWp/GDP8l
BtuxUAYxOFzYQseRrmQIWn2XOfeyG752mh2nDxoerqIH5YWMaYvZCoUZR/ysTRQgka54JGDJ2XWZ
Vgk7mI7kct323j4kvAs449NCEF5Hp0LFyOmjEaHT5UKSIntjT4ZZkiBor9rutnn7nnk3uoGmwepO
iksXNgBGq/k+MHBmps3WlUyVP837iYMdJ1Tj9nIYyno7qjBHB3xyPeS14U4McUVpXlIKb6jcdBqv
LySDrDm40gg2fFGqOAiXUd+PFwX+NC5kY1BMrg+CcSnoziicOuK1LxJ89fZ2m1c4s93BE+fjaVK6
jpvGoSrcAmYq6p8fd5DRlZymVQg0C9gH1e+rLNpf0qrBUXWUQvAf+e/EYT8ANQr3FZVuGbiawacD
cc26lLe5VC2DpLf6s6/kwwaWrc+TeUhifr4Tf3aIiAdyurqs5YuNYuNHPn5f9Ewc2yWKh3pZ+PX5
mR3JdUjJ4X8Twe4JyvWl4UjLWoLNw+Kuek+Hj3+hcscfUmNaeVhDq/K1Cq3/tgcRWf2SYeeIAzGC
CGO58WINnZ0+IwPU4Ftd1J70wUYPmCQcaN+77uJIssfDg3+BjtGHpEOSnNNSGssQKFyu4rS/uLST
FFw7w1IeNcQXpNUjbus89+/SoxSNXmaHjM77kAcCzge9jsCRKkuycOxnMtiuanAk0O8C2F3LOVMW
JolRjDgie71TgIoKdlDjD2IB6CSj2gQaYS5ZLZSkCUhT7ZifuZIbYXSIFPTTvpsn0wxfJmTBQKTM
ZBFkOQZa81J9vuEDjZ/BHzXzsI1wKvoF+GSDGAfftDN4fSEli4j3yi7eOmaFHL9Whzl6XWQpzEJj
oGstWk3KrLd9TYJ3PaCXVPyFvJ0XgDzdbiM20gsl+YHXBDjHtESbGxZJp/8p28SYE/Gp+kCotziI
ZGzi7JD6YPriRXAr5eeqQ8rXSoeX2ry75txvq2B/vo33JJKBazTxJzUiN4t2qEwKIG8aEdVP0NAu
462rA+MrPGTu+w7UcDuhySXhaDZRXajBStjK2m6QTcPAdw9z+YLI0U56kotD8ZLRYFE+kpC8DR4l
bk/FPWkxHVdCmHkCTkiseIU1wm7133jDTQKI5eqIteg7ZwxVRolJZGvD0nAi3qSHABv8SHRPSwc/
VezmDLHVVQMKavPMbQ==
`protect end_protected

