

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
WrSZEf64fUAl1kVl9HWWVm9JOgHMmzn0fv0uusEaRSoZ0YHKAX+sj6D4gL2WXWrV9+rdMofvPwNs
9A6zs8psHA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
R/iTmfCVAo0uuZTRynJ9b5Z2gujQ7+Xxv1u+96JME6mwR6F6/MPV4ayotodCx+xcD+9l4Ktib8Ml
C05jFwQ5vFi+09RjQvyvxQAR5CtE87QE5Bg2A3Gt5QmE+m7ZfJiQZgi5YQHL3kAHS0jfaofTkZIU
6VFVSW/fcrod0Swq7VE=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
RAfB7dvLyt2uCWNWspMeHiLYPG4TlOk+8Dptz+NhWH6nMzYrNkf7IWIjXk3hEVf7lwT/X64pynoh
QoCCtl9AW1iC77VMTIu5MgFRizuZMUfXZ0crSPULV2aGonx9nQ5JKx8TiRv5BTWxeAsuh1lT/5p6
2v08ZCt1Nwa8GPmEeFnTZsTB1B0jFzZQMa3GGdV0nEcSjDo4bLIkw9sMEBW2OdUuvE5yIHF6Z7++
/wzulmNKOqQpmeHrq3r1VKkMUHNzsDpLkGo5HMiTmEUJr/s3uq2EhCIq1agWSVbcEjS5uDaYcwdG
D4cRvgOxtT5sxpWA4fivRX7vvCyun+C2e4pYew==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
MsyF52v9pEo5RpJJtfhlgAJQ/9a172C6pJMP5S/aXQMuRuv2+JV5wCeynUZSXHj38Ger421EXuQd
EmO2OIKWiz2pShaEh/NwF+InGDF0QzD16vAgn24LAOYAOX1lcCquf4w2rs7e+0dn2PO/GYRn4rxl
E65F1qdRiZlUeVoRHdk=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
klspBE6zapxwDIEksFW+V3vEj3afpsQxyK1CWGpsw53FDriMhZB4hONIr9yRSN9nitmQ+6cnlGM3
S4Cxnkb334zdXXX5YoppEYaAdCcB5nDsYhSpn4PyPhd2ANmiSIXxEjiEJ9MDJlVIobzrtkNgFEWA
QkqC/Eky3QLBOqPuDJIgkf5UFynGEkI3eWzGSyuNAHTTYXfoLlYBh8nelaKS5vgYh7jpllyo5l6k
hn08k3sWZKuN1S8dwb88eFGM6hwg1UoX7pTnUY5yGPZZS0JEiN6WVWRmh72r5l3yyFZOFNcvByJJ
z349Odlh9AHKI6joGGP9sLtbKDrZfmu9y/SSsA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 22384)
`protect data_block
v+LLgeQTsvV5//yUPlc0KNcJ9gfCk2sPeXkT41vZ4sp25k5erBGXhbYfKwuEBVyezdXQKlkO0ByQ
ZlMybsZpzXnO0iI3pp5iNWb9wg+k1xkNFdBY2mozBMKDrhboqx02u9d2hv646J5XhX7Gjds/U5LN
1t4bcWmSbn4jQmADXk/VXgFLLImBIVr5cd1B2qzvzamOuip39jcorBqq3VRXTl/rIh2vEv8tRivr
I9al8pDrQGIMDG3XixFkHQOgg7I49qFagcw8e9/5pHedeRMaDLzfGEpeAqOiZpk3MNsgDy2Z5VAB
wD7iaZwodrD9kubcUesUDGq5wCGT1VuE1MN3Mb6Py2CKgkQHpSb2der+LMM+7K0WnRSDMyq0RVr+
7WSHvUL/yfu1BC4vfSaZCLkf/TcfJy/2PeUOGjJmr5skdkmRA1rVNTOcql29+Jo7/iO82JBr9CPC
rUPQ/Idk+BYg7ELPKLTqctAYoXdqaqX0jN267dMA0NzXs2ZMjlBvuzQdZ3wzFrnMCcuDCexg/2c+
igWP+HZIyFQ1IJZ0JGlnwg3SKoSZoJ4f+D/qAaffRq8iwSqvdTbdM+BR7Z2oRQxs3SeshsjSE4sc
xr45StxqVUC5sI2wdt3VvXn4+yOX/pNsbTfRj48xPFBOH4enB+EAtJvAkuHutVXlW4IfW/E+9kFd
vRAhiYLO3czDYcQCNvmF0W/YzhDxQo3GsJPvv327I25+TpSGmQJRo+84OnW1AOSNB5oRG/pNW3FQ
OuWRn9H0797MKnnXjzBWA1OBrpfd3w7NsRQEEmervgjXmXCcxQ4mZ+NdL/YZSGopewmVMCbpy/EA
/W0QiA+p9HJY/r/S7KsYmsyqBJf0685ywmCA1S63JO8N+TTROglH3yeYalFmXXevWeRD2nH8rIx8
g8cAWbd66Dg6GBtXVGVpUN0jZfbiSOfgFpsfLmZpa9HXwOOqGmD4iNYse2gws3c9HpAYYWN5QCmG
sZVKvKmTGiJHMSfQRRq1SAXuHmFejJOzDzAh9QqwNVKQ3a2wdM5lmmrj8XmNrOSThyGThi88H3GP
U4F8JVhSmHZAL65l7xcsl/pxqbx28csaOgplSnnXFxbi9qPEo8f+kVvnvduyUqFcc8Tl7W8/lsOP
fOjQpAR/fhiUbEDge5iDp9r5waheYgi8e1SXjS32TctUmJgbbjH5a05ulJuZsxFVKvZtxstNsA7R
8hslOmxgqAUewE78eODDDB+sv00+r8OMX5L1DG1XRrf6wl43N2heZhaYPbMYXg8p/lCp5RMip61S
H+l5SVynYbhjwatlDguDTdWZZPhPxsoB6rBLH7J/mD2d4Tam0GGAyIMOwfDsXDmjdNAUl0jPOhsO
DTO6VmWPUiFnWmkZ7uahMrWEE2qCqIx4f2WOpVFMxX9c9r+yp2sKFemQMR+GoeL2YorJBmhP7KQ2
/vUXTEwn6lJTGGfXfsrUofMs16EUZawLrU44ijXaZGII0/7uHJS1INkLjl+tyQXO9TeBmKUADYCC
Nq1EPlNKtvuI1TUF3CN9jMaxtpqWZ5czZAAMtNjLc15k1HRyHHmIkJuaccq7bUccNU0oS5TMVEIK
vG7R3YW8QVosLsq7PQhmyAlq2eDYl+6MABRYArT++FmxOhlqiREATcUYJGa7EuXgOmaf8pwUlIKE
YQPNC6DRRPJbgzYE3OTHUr4Q1qEjX8q+umoD9dOcn+aljsEtULXTgUfwOR9sOE5aPGzefPjSQyYM
SG+PuD9gN9dv3eGY+HpCiPFk7J5pkOdcJw7dz0Yi/R45dP4ATtTLp1apzXCY9vG4R2hp7tCeRf/k
/XcDzwzXSdiqGOD8kfsBrJcJRjUmsEaqMNBVh0nkwi/ilqDXZnK95sKIBM32gbVdkYvyyU8p7pMO
eugkSEo//sWiCxWcrsMkT165lIZJxZOozAdodO1VkRtmzhT74JOfL6QGlbpjp2tAL4X0uLa6rs8j
PUGe+QPCJQIIe7sTtyjAmPPDJMp3AMsUUfTLriSSl7MBd20nNW3e/Dcnjs4jBwXHSTe30F9g2AkW
DfXcYnLjn0f8HbqLKuHZicpgq2f+oA6gTYCyqqaDS0uZOVCwnj/GEMHsxMmeGguPj1gQ1sR9Skmp
VTEXKpp1s9EnOQhZvXbuPXFhsf28u8UTwcBIZrdRCRRPbqwOgQ1hQH7+zJQk5/eQ/GiM6GR7/7Tm
GqXoxgMZNcBdBBTcnEm8Tgw7OWLjnjpYo22OgSPmeqBgkOazCIk+f/2JJzANtsw4ecDPkVoW/nSh
k4uTWqhfeVDguoT21yQAkS0NpaeCN16ya9VJwI+skeupwqqaI8tXlnt9DFKTXX9pD4dfBvmYioGH
6ZBVQT126ptzr7sBAzkR26cff/yzVrpZ5gOo72A1vTNWU5UeTEYw97NnbfGQ/K198Mz5vt/ull22
hQdXabM/ma/m2MeqVrnbZ35sumHyrkqDtWIeISs7hgL5f1gqdgzS4a2HN5JQljzrRY2xLrJDgucg
dTA8BwiTgcRsCrXO1/ZRD+lwgVVt2WjjXNN54rWToLZ2BEOcEG5iZM2QxyWqSsjC/NmmSB9oemXh
qcU9Y7UZfpU0zftgqgErVRlZPAhNsxPIwYIW64jiEAzldCfSPuOsMH4gEpqZ8lHTntOiwwAozOvO
xdxaRq1ysxwSiW0eLfOEGPjVPrWGYSgAl9LNv2ATbZ8xM91XOMxLZ+BEkfbjPRHqhJHTZxAbFuQY
wGV2S9SYKSpEt4aUHnBoaHxs1xNIgPqEmojc4WOpATAVJYMNM4cZA73Y+uzvrwhtPLNh6GgUuUZT
QC9IrLHz9lqtro3poFnetPQ4a9okQG3/kQ6CEN9jED5usK0+d4NLp5eDhj4lu/oTywOgCE2mDvz5
rYLW2gnlxCUpFvUzC2LiSdy/9gmKwhKhzaRTi92ZtSFE3dCxgMCpLNmmA8JdtFbQoOtExSH9i7tx
lIXmo7On0pDRcbVki0LvTcx5j5OfWyFRoXtnqy0k+uz9Xgg46a9rQUZGpiHdbxtCTLpO0vidZHpH
fHGCn1r0FH1KBw4cF91nY7syFXxRgVPYQy8dob+VlP24bismJ6RDuSaEDqQaEPkCYX7EmWzji0PD
yVBkLep6zWywA2/nS82gEvnaKlukRS8uK8kU1Giz54HgxTdddDgXkLIfy4utAWtZQNPmNtNatztI
Yq95AIdmaaFbmLmwV4hPkgfxcJAqNfie8vgMmUiIkQ3C97Ty2byvk9j582JWdVoIlDJ+CtJjb5Od
J2hhMVqqBlseHqc7AOwtsBXaRUQe1IPNxkDQvAACxP2t039O4sntq2CuidtHE4VrJAoK0fV6qqrr
kG7gTzzpFy7l+hjR7QayDcwPP2ZM5p6pfOFERD5j3eN8odlhJ17dIA6vsnmiQBT7rjCuw7FIT8NH
swUy5c1d2ubD5B8iAlFkpXGp/P2dKU1W4y9AwcxI7C+ZYQkJTwmbPln3oHdPVQPKvky2wzDInUo/
JGrfOQEfABxeUdDIHTFKwsz+IqRqwdwS5tpYckNOTcYaR525D5DFRdR1Qd3RmIh7ZRSYG5Vl4efG
Ey8zdHui4Wg1GD6j2xAqVhK5rdjo6gG3+bgMkDMxQLN/060klzgn//ErgojNWfgby0z25FTlKFTn
iPJiEggtXqEfDNE3dDvp0Ab2Uiw3bZ09ialLw3l2+swdZah02EHAMeioV1tUb9U6tDmSgAbGGIiR
aKnv633lTxBOgYtWDeeYwJjSiSbZeXLP3pO04BpQWAUk3i732UChar7RCeucJ0VhS+VshJu3Og+z
rvf0YkRMCRZ2gIkhLN434QC14mOlXV/K2/AhBfmyxw3nms2HUOXNTPxDp5m0sgGDwMKEr6DRfabg
VDzB2ns+n8ce+KHdSPrYA7j9CPmWrlPfyVBxWIxPKiaul5LPu9BENPhzWGRyWJ2gfgg5GupGhKTx
macRgHaXU78iFYiix4XrdWCMU6sOeQlrvcfg9p/bd0xcBeTM3z1qHOdFabwIBfilZwCteMCTO7HE
ukbWszYYfa+wNm7CYEZfZiaOnNsDhdWGoDRbUq8hOiso0eoDfNWCgOrvG6JlOyiZTrpH6NPPsKaR
zX7t4yshusGrQ+ScVQc5hyGtkM0mWsu4zlhyQtSmC+cKi22PmjO17imZwEmFwLWOedTLZ1GgvQMr
jCQ+kYLCy4wsSBAXwK4/wzhXlHg9ffFw5goG0se3ZYh09HO/lUm9HtxRc7qDH8m/adatN74fdd6/
Tjme7ceOBP+pOydSq9QrxXc1ED0CW6d/2zeNXzTHVW+eXILOW2OGdYVZcHr3xbq5O2mpqw+ml0Sh
aYknQbdpCp08iOTQsEV8Tj6fhmVCvZ/zXxNB5pn62KaS5+eJrnPlDkMcK2Knw6TS5KHo0IEtsQDl
PePJrGnYrb7qSlU0sBR7kJshB5k+Bt8RQq6+sP506Om7ZDokDXcHrv7x3tp70mIyoUxOafOJ/Ajg
PIiwhvMwxRy47RfUSgLwonZ3mm9Mn5gTbiznOjzazn+wvFfYSxgk8gnzpvD3ea+6lyagd1se+/gS
m1fepc8n5gz1c0IIj+pIY7SzaitC5XkiIp16WvphEzLbGiFj3swP4FZUp6/+z84r/6yLVPbB9S82
d/elqhl2T8RyHvAFApI/6fgqsJTn3QrVRjufNnNZxZGIveyLZcv5brqPoMPwX9GB2ne5Q9EN7rGv
r9bkmUPzJCFt/w+6rruiuYXqiLQ3MYTecgK3ObC7swgpe8w0jCVvxvqEKTjLQc5WrEUJMP3eSRq3
CD1+bBDrU519Pa42NzER4yW/YItdUhEUk4iiSbGXKFO3OvH/ZuJoR0VDAC5uAxyC2kCY69WuNZJW
fEUZBDg0Vi/K0N7iAj5dFRx5YVRz/x2KIrBJjfEVjCsGCATdOGIXcErkn0r5YX9l8DCQjFJ6omNy
4xC80XH9mxtqcVKDpdZSWJN696ZRQrosGfkN4SF1XaGYZuiWxGQdzWjWK7Z5QnDO6/jQfaZ3nri4
W0BA3RxPTsZx5pXE5ZNdWALYhuXt2QJYSkzbBs+zyp46M0XJ3QTiDHPrt+CKm2kgk1K+ujnmMW4c
0NkCCcyeT5YA1UQ3DkfMIP1Wq9YpCzhEmuwAP5H+BViInYPheV7oLytoB8S8yLnZ/8CoPDSy0cLz
s2hP5fmMIGfWn8TaSdp7lZJlS9Ut4JLSLM3FA88NAV2TzI5iAf4JnKHJ+gqXiapUq8lOk1xF69q9
q9ulmXGUYsP3jD7X+uUhqFgoz/MzG2IdgCUUs3CTnfT3aTiOvqKxoQ2DZ80YiBfmyS0F6vGFTI+A
sDg3sNxaeJ/qbmsAouKBbCdNjyMFikVehEZOmbtMb4KbW0Q3HfjLF5oaZBtYPUv6AE69xj3VfvWQ
xeH/aKalusVwaAgohDRWcAXfMBcnIBW/y4skjpb8p5FkLqMLG15czEmcmK3LoEhbaXl3XJZBDwfp
Klzbu4JR9QMAMBfMeR45J0vT3YSWcXJ5Ixtk5tgYCuVdEl6HF8/IaydZ1UxQ71LM0HecE0dlpge/
W+V/ndaxjPbMLyFWip5t82mTo12DWWuoAK34Ac49IohHkbHAz6Knm3JOczCd+6dt83Towe2RikSa
J3926bqS9VfVbTPowwi2OqjdxJfb5KeqFun32R/o1JgkD0slPsC4T2jUCw3gqxiigAeRstUgABRy
zhWu4e42Vo1RzWG7qY0kPf4mxRORGnzNRbboA4ZjLgvOZp6T72U9J3nyABLqne4mR/a9XZLV2cxW
nMOQCMaottmCHVfnYbR9fXIByzw9l3RdwJhBfth0XlPtEIhxf1uod0BYSBaGJ51TFg64+xKRLUFe
yPt08zLsxokA8XDS5LIMi99v26QlJiKRS9riWqlG5aC3v8vRW0FcXpVkxWQ8dYRAp4p+9dCXdy+X
pBCdUS2vC5wUlZOelRNZue912FeUhqCMeHfLpKbhgVJ+HpFNxNnz+MIQ1XGpVteWdcKtkGb6OlIG
XaCcjsyke7PyBQiuLUFI0alJVuttAx8j85I0Y60JUfT+pzkYfd4+j9zhZYEs11Rb4q2Ab1tsLL6B
yUNwYqTtm8NQP07SUfh6j14BOCN9483ZRRVFqMENth9JIt8n2Fa6CRt0eY1VEAFdjLOZclBB49Rv
zSdXT98DXm4Thy//PvXXcsYJBzWOKiOluo2t0gfLECD2Lo4ZJFBF5mBf0OrNIVN0QCSS88Evxf3L
9ZH6lQAvDIyiib6jdUdd3Npj6dqEkDjY3rzyctt9+LUD6sMq0c4yKxe1sot1qv9CElWWq5sS9EJw
u5YCmBKRmfc2kQZW6c76Wq+9d3gJPP4QIzqqiOveOPG/CQcNKlJ8INwnFulVCFTfmPyQbgA0ni7A
Hzz7Qc0RVmJFCoL5d7diQnoQk/OjAP7kv2/aY6/xr4X/ihmuLQ5BK9DLx8XKFoymGIFv6NKuHHdh
Z9qp1Vpvy2B90dwva4ewArppVAIFcRQMQYZw8q7kjEc6d6Sc9z6SSmbq8i2X9IEHGG4amgIavcTr
GdBxW1nkXw1IfGj11+jtOdnw/pO3nJSQdM0X5am/GF5EHeUkpL86oa3HD2cbxMlxK4FGNXuvungm
PTBw1Ijc4xs5uRzHzL1MDGCcRBWuzqJVLbgu51Wq0A0qhaXIXAIGrpYoLKFxpRx6kbndunA+HPeQ
XSWV9DQPG6QDCfk5bUv5TTKGTV+tk7vsm7cqvfvJCPcwVZvrs3cQXoFofJLjfwTS2MlRYyvAR1kf
gIGThUxIwt8NTR85VVlUM5NJpLHuU7LRPVEbalkZX2EWChDk5sLmdjWftn6Cj5ppEDs983yvEyS+
2zFqqjruuPqQFedNT1aIGEhs6SPtDjSM+3AkjtGJ9ggW4O+IkN8ahZa5G2UFKjRyzwSwe17JYBI3
+BRSFTyuZ7/NlkWBIbfNKtjtQmh9uXPqFGWLC03rH4+sDybLBtMKtKWTWKeZlgZldATPjhGR3TZc
9qyoa8KsHqI3uWF5TUwg1dQj0T07g8UjHlcgeNm9u+F4EKlDmpnVmR1ok2HpiOZAv2+eKqeU341+
fjvSCKcsOMNc5li+NIHfwrd4KdkcHEMFwJtsaCME9qLVMkxURmVkgxp33/0KItIR1o9e19caua3E
FZC379X2KQnnAaYLuJ7uhObVg6JxBmklfJwo53cmD20sC5YUyF967/YyMZVSHFvo4w0rc71YgCck
WyOVbBp8ulai5MWjLqC3Kds54Seyj66s/gNpx0VvLuRYFjkFAaJEGQkdoFxvmOAA0YqFJhhq38WJ
D3YzqhvsVaAnl3EI3MrjrmJx7aAcyNvUfFqRD/7AspZEsNu5GOITamLvDdTiRj1Awn0Ks099/Nph
Tx1ZQYMplAx00pMBaiFREVRpIklYiZg+PshpGyG0L6p9/wuUQQDFCXDiqq+oGeZwcMr5NQ9sFAez
tm8UVGlGh78fi38RdNo7y96+40S2UXokYwPRB5c5tBVEt5VXeZ0XZmvL+r2rpUs9Kf7wxga1s7Jv
sa+chArg4drRDFHqM+0THda4Oi0FVx2YspVtDhNIgCpEi6sgauAzsKGqJOe+7Y5b3JDzrp06dKTb
2AResasLO5WEAmnbmWs/cfJ436W9bYGqb4DgKEEbZ2SZ17ad4dU3Yqq6BKMe8sTjyDnt7jWzJJP+
jzgf4wRx+F8lzRgKEU0iyNcMWc5CBNeTBZeqwZYAbJqx5GBLActokXtFmh5l8H0H8VnzgJQ1kkod
YYKYjT04rl/Wq9+BymL0B/kXfSLty3kLzeq7rdGKcn/fOu0izIBMjWUgFzqG5Fp5BO1jAa/7EB4i
qE/X1AxJljZB0jFfzVDXLrfzh5p1xBm0/hBhlsaYaI9ryp6Ckm1GZxK8ky4EApSs1qqzqHOCDyb7
d/SsYmk0de7Mgz3N+SCp0v8JNUNw3Xc9QwXaIrlyuq618Qq7fpQ/N0BU/fXqzHaR7fi0NjiXk3vF
OlWPJcXvAmN1NaLfQa0Tut4jTJO05aURHeO+3BAkeOf/j/b8filNryFncn9F/H538MfbUVEp6Pb1
yQQVISdfRurWxAjIz70WOtwWam7DOEdUHZ019jYjnsPMhbAJk1tV4FeMba62azR8yMj56uK4k473
NCanR+HScF69ApfXzZXy3hCYI9KmPIwLrvMdDPCX1i8qHLeyaNvVHa4b25ZWcQb/LJ+N5VTLPjxA
ujQb8oCSxZO6gjpiknYx108e9Jgc4DeLOS24Bkf7U2/AXuio1SX0khWxPaK/ySOjJp81lx+SrsJs
nWgNTV9prlOc2FZgTZ6klU0ousu0GFZka0nQ5TMrPcSHzOWXiogxyg83Kq4eQiEMFTznT7PXGtAO
bD06qC1m8Fr/3nlGGWzTeLwbwSivGMPxnW02jElVfbgHdo6HfPkfvFlIoibIxbGIyicuec0BYCov
J7vxqvh1ULWc3O8WtwD6Z0+JOGYWZkNQRyYo+loHJL/wD3WwPfoxD357Sq0O+QkDaipzeHFMhH3R
+MtchBjPcqT5CuuPjhrnPRqjWkxkfFuib1p+6aW3AhmuvG5POs5hSiVPKBcuPFxzqqRXSJ0ZsXHK
0rF1lAYH4ixVKXo6uleI6Jm5LWs1ZWiA1Hq739wj0AVccpiB+P/ZrCWgL4YiO/reNjxWirqja1LP
h26l+vGg7IucAn88sDddylcnTThX2gxBhrakbmO9Fs4yGv9j5zYjeOfjhgo5GoD1dCGPeaFVW4yZ
dwDyguqEUKy4oCJ5o1GyxUYbAo6yfApiE+0XkliY96lvPfowG393N6fyxxxFdf/1CKbgzU0DZSU0
NeuclmFv4P1LMY9V7rD7jivkFrwxUC8liSPfAJLn5u4N3q6VBzdp2igcJW/Hqmcm96ydYGnYOJ4M
bgHQI0yZiJ816uUoFkIB1CIIzBNTRe0/tszsVcor/YxZy1xZEmoms4Mstfk62oeqSfF4DAa39JQm
w6GD99Tjj/kY3gbHf6Rma8VmQ//fS8TMd5786clbbURn2Cr2D7/xJ4iG5uvbarDgm9x2pLevAAW/
Y4cJYbDS1xPzjzcn1buFbTbpylSkOnAqMzEsHHPlYiMFI93gY7KEa/ky7cf0IjWcCTfYyrKFTYkb
QYFIKO/ZtdrZ2vtrElRrUWipiBGi9XcGlowk1pFICCq5ymgr9PzsXVkME4Ee+7IIB7Yh6UfCzyRx
bXY4FZLOhLrimKpyZFu3TGPxzX13bJJwY/7ArO4OObS1I3mlg+On1LIH+NXGMZ8A9e2ByVyySl+R
Wb0CI0w8ZxJHuOb9M1xSMvqgAqfpvUWU1Nodk+cniVEnGJe5L8IcjAQiZa4PTFh2AEPSxR5ZrJcB
GRQiEUnt0m9DIjvs/DyVFKXCP0UWnItRN9VmLuXubFuoyJ49RB/cArGYy17ShO0XZaJqh/o60ngK
2ydTvSqhOxv63IEkd+Hi4MTRugiIWUWvZruHG7ZrQ7V2lnEXi+7qGCyl2q7of0qYlznbIKWZaCZo
vFXB9sZQQVHZLTJBZinuBQyM4KxgwV0okHBi7a3fUiNahJrWo53ET8k/xnA7y8iNI+oLFdS1jpz0
l+hsu855PUBrvCRbiN/4PBru5dZuQWUcf+Flw2NSBDAU+V+KoI8AXmaJuSMPY1ovX9HMuQsolMef
jXpNphy1sR4GfoSR3+yklIcXLdFszjS3LyP/BPaBCGndNgDLzLTvrs9nWA3oYa+JMMEGd/zYM+C6
r+Ui0mHGd8tSFy9h3qEOLIygQJ2QS3NL4in96MDsQaaBzg/RGEDLIOVTt07F+mEQXuifE1XJG2nq
AnxgW3DSJyKMBc57RdYLjj48otCovaQTjlO22Y3kgrHiOKEc0tzPIfatrsNjavlBvUURQ5lSHpi3
HDODesGBer0VoQzUrm02dxvFdfSa6jYuyGIXuvmN8DytBuKsn2xDc+AIgMj6mqMwP1LRqJrfN8UZ
w/Ffdcsm8hPGSu5+hXWadRDchKBh8Z3JJ67xqvpKoPAIa6aLKAqYDxzyMk2MAcIlJwQQgH4NH+Xm
u07Cj58Yjm6NpFMmcSeuTmjQYVPwzCl5pWGaMcivHHKqtRzU8Y9AqNYt0lEQJ+6NghK/lL4pDCcV
IiAV4pxTfAb0XME81bWf0HsS9uSoGdmzgTwRciplTRq5wcrzOILi+C2sl+30X1CtmLdjnY9Hdrz5
re2UchAcEXxIF9G/wXZS2Ss0fUyyYaFINSqcu6JPRYd7FcjyqKPKtNIYnBDxy0/hUErkaJFLLegl
aUk9Qj+LE6MDzb3TR5g/v5TZWcgDgOvv9JRhmsJU3UxR3r/sMKi3W0I/+xDkXixnjFmXH2mna51k
Xt1Ek7KcrKFH/D4mPhhHvbgTtzFjbdliOJj3/W8UUCIuukJfcv1v9rkDJbAbrbqA4JCX+YPS5ni4
JFDM6aiRxefsxuXO+tXac9uTa62Myr86sMTIK8L8kBoO2TBedipM1gNDnmfras4ko2bWTxRuMXgq
YpT0SSLh8WQpEVJhWfYJ6kyrW9Z/qsD0nyHl2vgK6FZxf+xSBLzXx2MH62cO9u82yGMPTz0RNpkg
79gbEmiNgmTWp/eeZcDx8XVYQWPSizIdNs/PBFInqWcQF84qsxL1MSgo3rRGAVSiWp0ncM5bEGJ4
fz475O50uXnHFpqPnyIQcdoyjUeWz5XdJ7ExCQGnxE0KH3trpZVNHsIxMIUHZ84QedXuuwgcFfex
sVBPi+b3dpqGxi+eaeQuHaIxBDHR8/Xek932FYQbh/96RcbuG8R31FebJmwHgrCTpPM0QwNwdBxU
yZg23U576P/mJryy28yCB9Q5O+nzC3Ky51ISK2O8oe4IFI2VvchLCAkg6J22vbtSOAnEfTyj7obe
t4ahwYqzKoM3XhcXVuOjr2yG2Xdf6h2T4c+FAkfr2VLMlMZehlWOUD4uKK9StNQI13LQumYfuJ0q
Hn1pn2lS2eZGW0dSq34rK4zCogufU8oCfQFr5ufVVLKpiT2vociNZNBQyyy2H9j/RMKETbkofU4L
ELVsMtKsQD1/+DCxYfC2Z+/N+lvoTvQQXT3xFIWU7RYCqTRenib34BgKeggKVdmd/lmQ+tXDTytl
/KqSt2maTSq+DuxtTyMiVvFAWUvQWPwZZFtygOxrPia5JYBWL+7JSwEFOAfI2qaXQ8dbqhYZknfo
XC1i8XzUBuu9ZrFb2ZbhLIo74aDrmY7Dd5vdxxs0qHZq8+M4xhxDWNtkEo92udwgJnLndHb8FwYD
YmhFR/h0/z0e7Cfhb/d7OhH1xROTKCTi0XKwecpCLJV36HjR13zqlMHtju1mp49jvpEkG/htx7K8
g1rZOftnkzIss/nZCdlS4Vse8lrGRKivj5mUdAbfcGHoqLCgVn90xx8a8jeziLjMOew8aruIZkzg
dTYeJEvLf/Op3m8p81KdowNoxZnNML8Tgn2aXiClmR+dPqeTTjZzJ9MApVb7HqA/xny3K2mL+gH/
lkPl5IDts3N8lDHmaywi0cezNEOYH1wgCzxRIL1wk3xs5vJAcnXvbUOlao17ZVWdZfpmQ5CZPjf6
xOTI1RFylCy1bVJErD6zi8OpnTAqm5ChM7/NL4ArEfpn0/TZ8q6s5a9ef4NPBrnz0OHoV7zBRRKN
NlzfyrhCic+6sl2fFg1vbvHofdsEa7W7yujweCoImMxFP4kGI6ZINvrjQ+9OwB1Jtxekuz9OEHuP
MtAAoYnYszJQYxUcPpOoBlnZphj333OdwURRlRLB68NV3PuH0LkQrGzBRxuVbM01OVL1n0fvH0B1
SNiwZ2HZUu+2VqntkhbX0Y2VLJ9wWd9bMMUTt1XOI+TjDf4ezljN+nvmgEywPzsvgjRVDFjvgeWi
I4PeR9Q/DdMXdse/wiW5fmShzfiQ4mczG4xOhnT9R5oqXPL26bHW4vFRzrsLg8MnWd+gwwBUG3M+
/V1r68Z6s0S7NNXygNJjujZ/JvXzZISQpoq1/jbOKnADPT4K81q27LSHwkzSU5oljJIqY6YtvZJp
r1SDzcH5AsR/EBQaBDJA8P2Tqnoj1fQD3meHogCMU1bHESDsQ8bdA6z4x9dz7B88J1/vBefcK8Yq
uzbDCsBo4YrMovWH9Y5YANz3NfyQxH9DCsrz/FgT7eHybMp3SXj5v/PQExbnjLjhTHdFwu7rl3ga
28zSelE4PCgPi9P8qLXt/sNBs9AZ89uE5nr3NXSXXNLHd1YOJPGdf5ArwxaJXC+ZlzCS9KJNubuM
YjBNajUHGv2cppDZE60CuwssyJvVZHqBkN2dZDvqQ771NgHdqbRRv9okB0+AiPBCUgq/cMz8E4Xj
/gE01hKRNSVBGQBbNKZ4MsBfWE/sky1sIo1MAwUOFhz5JYALwsW364QAkhLdZlMMqVkEMdf4/FcK
ktLOiLHPwt7NYc1xhGnhr9sxsbwj0eoTG0B6Nkfg3Ae7eaIRMesER8lsIavy5T27PbuTbCgES0Hl
2SYIChg/7evh7Q3TzMsgd5/NjcND4vsonySkmeme6VX/HedFI/K6mDPQrAN+ulkcxE4wsYsCp30O
VGKxMbTIIPUIvBSllf7/bMGi9+IVpOaeMrkM7hM6Xol33xmArMzD1vqz27fUi5oNTFhXPgYYzo+Q
TrPsLrU/Ob9FP7KPP8YNkXrCQIcdsUrM8Pcbd90/H5xFlyzVuVHJ3Ni/CZKCY7oY2VS405zciTAb
RzH7ZFice15PD3YLE9OfFLAcm96nr3OFwCRq6N2rbKEe0haUGwPW8y2SNd7/HMWuw3LGeJMpP7uP
qHPS3jZ74sAgJq73FdUv0TCMg6MGNP64kZbdJr62VrTCtZauTn5zRPW/S9KR47BKlNCZQYD19q0S
FRE2eATDSUzxh0X1yzhc1xUoG2CJwPseODVpexGw5M2s58J7KwRf4Ics3PlNDchbNURU87iiZfq8
Oe6qyav6EugNilV//IaDmTK33j7nDIdMG+1t0+N93An0R2mvnmtz2T2On/+eAkT4VwS55vDGVvoN
ipSddUP3hsRHPIl67lHasqRZgl2xGt6oUqHCW/fvZov4n7sZQEh2bt0M+HuyXwIzH2rYvshp7TwW
vw77vhO+4pJOv3YlkL7/bIZ3isW6mse8be7SAakIdTh0aylBM5813jqOtBAuwLF/6IChg8ndiNKl
5sKI3Ga2MULtwv2NL8Gw2c96VYxdJCM7Ori2m22w+Ox/l/TfCMe2gL7J2YLhEcK602cdg2Ko47DN
tB+n6cKMkhPi5MJ8qxFmynGLZpQieKpIUsRHtvGqJej2fQ1VEK5s8w//5LDIubHHnbTD1VcmzEyS
xJ6UPfLC5HhI+RO1jDKR2Mmh9h/4DM5izCqTU2K3F/gB+SMdvET/p6LbzEF5K4NDMeyswp3x/r7O
4syd2xuqHTvDdO7uoNwubs+pXGrgBQVsYNAXlddr3U12mJlCnSjw8+sIG2fd6acmmmr/AxfDUnkX
WcQeiYZ/eGkxVbEo5Xwg4lLJGLvNBByAwyTBZ17KHXVSmXzhU/fFJoSMQSfVGk25mJ2nwFVSZpfA
iZq5ocLDx++ymJ/EaV4l7o5fS02ZwfQo80DE67X/bCrsjTaF0VF2RQqWI5thPIuUzhxldlqsWtXa
wI67dncUnATvI+/8KmenwswfH2M40KsFy5PySx4ld51LcaAMwYq08HYU18/hYmN3BM0HuCaG6gqs
FZWv2Bnl+q6kTduoX8wWpPcAMCe+Ts7xPfHntl238pSzh8qmX9q7K8jo95EmmFeSdb8zPCvgyxpZ
w/aR53YWN1RByETsYnvAKCpcBLtWur79FB5rpotOI8t6e47r1APR/F2smAlXNPr8in0yuYuD83qo
wsV0ZgVZXLeWSC3a9EYLB+NN5PMUbwdqe+F87meSaBKZ01HnvUjwIFlQpIIceEkHPbav8emqkcfT
uYowSFl/Sf8pNyyEpfTYgn3W8Ku39lzjLzkSrwWin1kQlVPXHdCJoTq7HDa7Gf8+cwHjKasMKGfU
OuR5wR+K42WSkOJklyrBDmPdAlHPqm6jyC1C97WWdyoVl+yQVQbDB+8hiNaLiFp/g6R6eZpEViWZ
cVxNmelfVEUkVBUA4sYKxUiYp68qXc9ccVbd3xK7VpUX/zFE1/GxU78LrEinuASKxETLeXsbZzzz
YUvycd9WkD2I4eDKkjn6WYORzgthejmaGaUgqGoxsCZkxoiLG2E9usv2D0acwfQXEGbR0Q/1tKVb
yKc9Aj1u3rE3P7cpwRy8ZICU8HpryBAdcQ1Qo4grsXcvTfFgtvEvrHmYBfs7Vij1o8nCM1AUqwrt
acvhLQbj+fxhImbdIVNF1NL0+sVjQn272w6Swo+6VVAJ29r0zWDXkFasFYuxuXmII/3MZsHzsOXj
Nps8nyyWdKomw/MxavfatdsSGmKkI9H9anM8lbRPe6PjR4Z4J8jB3jAZTZ5Mxf8A6tMdeVDFRjC5
T63x1RJ8Iw06jKUgje5vS7HaiAfjZcXx/WRRC6DwEueAhbNy4RIvl0TpQ54FqJrdxDhXlwI/n/IW
rWFUzmFJDXYRzG4qzDHQE6jdu08qFXhjbAHlOLjOjljunhAHniTxa8FOdodrznD56KNq7c6iccCK
UZbDwdzo6apekSnLMUNDstFb4ed4l6KrSVZPp57IkpL+wfnShgE5jyZaj4apBFXNaADGBLqr5MOY
LOnevLaRTXszN+n8EaMYeJip57RtnG+azk4LE+zTVD0PBurC6TN5b/WgxydUrgvHMFxGod3LSbFD
Swu+y24UsOGvkGsV6Q+wAyg/LCUujhwBy6+FO1qKR+DdWWbktZIu0N6NQdsu3Y+o0uHqMA7yECkQ
hkCr7jC2yJn2fUeaVCFDy12IHN3laqpE9MKKbt/IHHjnvkP/S6ohcUwPZMCYz/wjKaBhjKvau6Pp
TeG1XuF2oQzuCrrbH+t+s5Cmgqx/NZ+MuRTMJ85ymNZy0j2J23tkXzpuq6fCDeSXzko99EktgLub
FfJVn9uw4mLjuf5WscQyHwNmQhQhusi1z5OKrB9sPvdTDYBtKd/24Gz7wih8gi5WZ18ci6xgWfir
hD4Y4MBtuai7hfqt2cHt1F+fVTevrdHYyFb6jSB4M/kZqy+bt4WdCXWebd4f4hNGtatjzTZVyFGL
Ke5TZLIbczJqsz2sSsqFJWfbGGdI16HgnaeGwXjOd6o2RIcUP+urtVDUpY3BAUw2oNHsQkSCd/O2
JD/0+iwjXf7m7fojkHgjMSk0PtgbP1jT7zm6dTooGjj33EqH33nooYz+geL/5ExW96Umg7NAC8S+
KqSxWc0wpBl7e4z74hy4hh5ctQXRVYC+jJ0N1jiOgedY5lTb5ALXgkfEHtzw5JDzbpvgvUH5g10b
g9eocaBRM9z2N4r8rSJ/VSXn836lqMD3bsqGW4nOCWryPQhecIysaiXrd+KFkh2pz0QGgwiXzc+Q
khP9P6k9Hrw2WLzz9Xa8jbKgGltN+S5nnhBgBbZadvZRZvCMzi521twGIJYL0UQKarPC61JwJlrM
uVadXvByzEFuw8F48yI3R+CgdjjOW0chw+jcj86bxGQVJk0ksL9ZZrwUgfF8NkjtTku+ufUs6eH+
cZSCGeEm20gqQfOhi6RbfIFdIfgYfM3XzmVtEygnmn5zX/Je3KlSNABYhpTzwptt3O/AtPWEM04K
cmVaHRP/pxBXrmRk9TbAQ1dSP6Dvf2XXKICZVPXA1r5EpI7Id1RoorfqkooEBk9AR/lMoStWSjDj
NTcv4s9kXL2wc7Uqd0E3mc1KT0qgD3BBHAIqHv3EvFaNpZgMSLVbw0sgFwQ5SDXm2OhlLh2BExBs
Kt5rZEhMRgTwaS17s0mSoimKWX3U3MawpoxiJtXawK/b8eDPVmM+7l6cKO4sDNzBdMymk/AHonno
bPXOTYFrJAFJitKE7yEHQ6uhC8TndRsyAIR2VXYszb9VrQtrjhDO8jGxTEd50/S44vEQaDbfOigC
hV5v97mYwJTYCEc8ng8S6d/1QvWx0lr/vc4J7QCBnhEEqJcjrUAoYSw+IccxAvu7VKDkf+cGdu+8
RBYuMa42UKLzPq7hRUqGArAKq7KuE4HZPIDfKUEpue+3nPqcDJiYM8VGcep+540oyOCJNiWeVkub
2qJDEFAdMe2gIshXNKguqG+9F/BfV/EiGQ7naWFE5mi8bWhKNBwE79z4EU2mIK+UsqfKsm5qEyhI
cns184/mIgDKAcANAUFn9Eow7jRJ9Sil/0IOTbmAtH9q0uhNq5ZWDAo4Kz4MA81CV0bh2b87Xzsp
gndI3OeVcvVwNtWn3vfKCbRWyLehjQCEyr15xGVqdcC0e2K4RNkp5ISBv7rvd7c4C0L8yiQnJGiq
oOSMslxE0mf7Ia8fYXAdfe55xyHEKaRgbXKKAFbvyTEu4pvEzhOjWljJ2cKHmBggQK/o9CAGdV2L
W/i3ZgS4FSRlN7uhtUm6cJrnXjNpnxIokliYO5XszBsmurFaiIXHstq0cgPnNBKF3XOf2KwY3Svp
EOJ8gpVFW4ja+70p4fyrCS2CtYasAFZ3C8mHFBwMg1bIl6dDlCUYN1EbUaL482zvrAVnlm2SKVEm
jjjGYGVEYMaVcHEMVavjRrU/tALkDgGVqEm0eoUkmyNtw+ER2d2jS26ra2euufvvvWqlJBledwzt
4E/ucPzYcDFn0n9nDWPtLXv4e4W3UpJ4OVGgn6Vucom8TkhigG85a15o2QbyuTl8TWgPttnFL3WS
nVPZUXrKF51wjEjEn53XP0XbavgwI2RPu+7VFYogExeKfy8clRM1swF3M8fWmYlu9mDjynsT9/84
EL2KSEKZnzZcxlIZQHxKDQg+4bURKf+Fs+PVYVGh04TKSOefjeB4AkljmYmUoaiIrz+r1fgqyhn/
S9Pz2wpiBF6oWfS5vkNzOvmTS4XiFQOnVcQGTqlhhhFM0yZUEC8udGcBW4b/8NZQW+vYkKXG+1v0
9FT1ofwzo4v4wkCP7Z8sp+JrlWEOXSfpxEn0cg5Vwrz+PqHPIYG2tpR4toPXgSYgn3NDsuDFokps
U00+yJxBQIltWl3qLqbQp9SCuMmCTlJBkVWgRCX26NXFRjOvL+WMer8tgi4egb7/e5labD7DYghW
9t25/OyMd7lhvvKRHVAuA6H0TqZ1yZOoWmqxlKwQ/gyb0sKfi4r1Gq26MXEvsqgWNaafR+Rc43TW
1WVZutvIIDucF/d+WCZfG9CADvMob/ZvfRtr4btWKHZ0098R7Z+TedAVuROWGcSxPL4WTgoQj+5S
+DIA9MxStyLpENGEhaOhm++Gu/0taQi2GMdEa1GZbb8ZD1JpaLOV+IkNXXpvegZ4vHXreWObW5PQ
qp/Z1akN6g3f9nLbqi0q3oCiQvPzzFuxWRcZeCunXVdKnqBBZZkvOyjg0W4vjTynSUKUUdIux0NH
ZTwY0l8/cr9WKeJVKCzMo9EBe2Fd9YufJezpSFCf7FcwLfF+Lu46XZQ5hFx5EOX03KVvY9/6XNb2
J6iqfBjxAA3iwDm3e1a4NNdcPx6UVTZU88G5w3RsQcEDuY5of1CBSnGCkjS+mYfH/EfQ07maL33i
uCS23VL/3xsP6+XL7K2Mbn8Yp264XCYdmeetumHZ/2myptQbPDxwgYk4hYKsCjoH8nfrTY+pvYxm
K+by4FTgNjrlfWqe1Qt+iQxXt59YAY0v0tILoYy18ZZ61VXL9K74eMoC6Td8VPFjvH0Fc6//i2RU
WONAawZAiWYohHLGZEq6dnj8dGuvY7aWCFsGHWlVNf7jXDH3yPMxbS1ZOxpDVcjVDDw8bt1vgyCn
9CDxz+HTJdCFb0ha7G6Xs0XK5I8TuRdsV2aki32pfqUaNug2A+igck6ivHu0A+0/cPaLcuKiPbP7
B7ypy6oLwqfvoXctHWm7OuqhpiRVxuxMblSgDzo5MUVLZ42dvSOGj5k7GJ0JXcrDyltaEUNJ+W28
muwNX0znjXfeypC/Yyh7YGuf2IKoVXRm7Vipzpsd4GL5I12ZSSjt8hWKZMGz301l6cOXJoX4hr1X
neZ9tKDyflBiF7oQh9CpQ7t97NNZ6DfpBh95K6yIXc05B+DzS2meDSTL26uv9JVETVAMZBUkjOcP
YvsPS6y9jVfD3D8o5uJdvlNeVmm8Me5vaWYnOuTUWNdysx+XTlTfYvu00wbXQWjo+D6AkbBGe8S8
ssgY5vX2PkTK1tnzKEDPDiXSS5jwmgSe5RIKvWdrENInU80oqK1NMBlus6pY/rnPr9XdY7uN08B1
jJu8uD90wemnTOC1Uf0j7zi4khmMvNmCrn6rNLua1QND++UVJCoGD5AEByp2iEyifMFUENwfZSG9
V1jpHAO4CmxelhC8SJ5COjp9jYWmK9InbxiLdb8frGwQ5AkissuTjUZGFxIIF9RUpJwQDBXMshga
KBQBXWKE7Suln8HUlJe0/QCcznbtjmCcmytNVKpaFsTwd4Q6a9JZ8Iw1POq69GsCLcidJ9jz9xH7
1UQUZllrYsS7vfj13i9w0ulDrJiAjjTbWJcPb9uMHeGaKNDxM58zfr/TYW95LxlRziAsJBQjkzys
bY6h56YdVoUpCEUnqvlp3OknYvd60LB1VoGPgkEL7UNHG4qDpANJH5066/D7E138WUXB7a6BovmN
sqo62Vd9vb6VojE3ovgtmjakBC5+ADMoKjgDZuA3xVKtu/hybgZAuUxYMq3Ew5cyq2OE2+JTUd66
VqkFLPrjwzcd6gLGtdN1LoME8qyZLBghSe74ayY7NSxbi7TeotIQSNBOQ6Gm0YfpGwlJhiRnbmr2
vMnLv0i3dpglW97fB2q15U3HEEFpTieSfyWAOtu4keNAdCK5Yg73ecXyRgclRyn5Mk8fm0Dsm6yr
0zBZnl332rsJITrdOaCYj+bhVbdTgts255gagmU8tErpBp015dPgIpxa2YsHWDDIjuCY7ucjCLat
X8LsaIQ1rCMA4/ImmjPrGgShUUa28fvGBbi/ui977E44l856Kim8nkXXQHjmryIWEk0gQTzB9UOd
8IttBiKqHW0sjNTDJdakWVm3w0JNXudlKL+QDtQsdR80JGLK1GykkltBHRAJ6XqcDA4dYISfDtln
VaLF0DJcKDA3YCBnzvfn6vtT2NO7HPqe/JBeumw7OQoBfVMHhTxAFjPJe53zJSAC0AddaEsycDbm
vpk44ctESNuOFtlsAwkC1qLxhazZvmK2ENvTWzJwUC73Kd95kbXCobRKNBYehCEVDGVdZA9CvRqf
tbA6xLbPk/q4r9jdEYXhMX84+LFOyCYv0+lIqO9N4uMU8YcmzZd63Q7S4DMveUbxFi+yRx0r3kr4
SQR6PWyw9/tvkC/++TAlitVCrYRZUVczVUpm5IL2lZ56q+Vw15hu+2N1SdTppwBk2K5RIDJuPZib
b+Olbzq9vSxaZ3urf30oWGkTnqb6U4uwPOZyPM/l1oBT6wQWhj9ygaYrXKRFpxGRN28x1vSVT/Y1
Hn6u6rFWd3no4GfX+uwxsWkyUo0ZxNWvsDHdM+l4dqMzDPPwgSel4k9Ksh4GRT/ix2mDzotclHix
RW2dQDhy2NaSNCYJmF7T5ZsWTuZTnPwnKcQbXHAosMF7oJ5Z+weCDr00YGuLx+i+m/x1C0maWVNt
uVJEfhgggE8BpinjlSJK/wex9zq3HnXUuKuWlXUgibqQO2waXhfEPCVTCgQuXOnKBXcp9gYMQPHQ
YqxFHl6FMSh/1kODXeEH2Qy/xIhyN4WDFg9ARfiuRtJJeCFVzvFrNEunfcdHBK/GNu/t30OMk4JC
yg4JwFyz43nqgDwFcAGfrTfQgQbtekujpPCfMWHA3kP6ybtWEhWkrZ59Jne9jMt9gyCNPNHL6obT
np6vGmnPq/nv4Kdiyy5w1tXjpbp9s65qiyVWkjSC7ezi16OGyO7uMqA0ENl/4TF1lCemk9XmC0jT
QbYzMDg2KNZsnLfDYVl5tMxQIvPNbKvGjK4YfyJdMj8VRVrwFdcsjleFbDpwcArE0flFsL9X47gm
qzAfZmSTiiADAhVa1ehjQlNMGl6uFcQroajzZSWFwnu0rLcibZGvgxl8CdWp48sg64wd+HsSAUfl
Kr3MLXQ4mOuOQLly2v6QMYm6lIZ8+KkPwHBoSUuR4Ws3XpZvRSN9EDlHp8Po8vfi7KM/r2EdTtMf
J2c2YmGWIdexrNr6eKCSZg22USiN63/CA0vLEE1vORQfGNFYh85SgGAvozmWDXwJ4759n3X1KyWS
L88ijPJO1W6/V1habAp7Ji1n4rmH26fkuodsiAiGhkTHscC+xF9htB/s2PdAcrCnUskSQofMI9ca
yGZuLTPRpITwvTNJGn7AvwhPDbzplh4AuPoXjSYY0Gcpl7aIzRjofagjQ+fLMOp0bj4BXUHv2UNH
wgefZpRvKobkAr01o7RzWotHEzLjxLYOhavcy9favLdYdRW1rLoHp9N+TXC9x1vu9FSab+aMmLa6
7RV2bDkA6QDCTEg1WPdKCD6iR7yKPzW38o0XAo5gN7G1ZUy2rF2HV6bEZDfdosWMKehx5B0vw0R/
D31CABbgGAGDYKP00fieT8Q1VZEBBJNaT4EjMqrzbQs2PqHpN0QIauLZMozNCPVzLy3VdQXOUhCt
8u1zL8MizOg7g+28tucniUsyvbCmwHxUtTRo6bFyDysCAsAGe/A0nEwL/Zd3xjFyjqp+o+LT5LvE
S/ja89+becbL8Pd5Yzhw82tcewP1mYDi0+Rc66oEvMIBT8GImYB7jyS3gaaJzbdNdYpQtzO1uG4W
AjQR5MP0mE3C2maRKKrmP60sBDCwJBjHzMzp4fwY5mCHLNeR2OREvU8iI7QGZs5x8KHOroysKOH1
MErphNPiP0OTbMr5kmVNw++5hLV6wWpA0FVIXzxkK0OurRE0fuCdciTV2m72GO8KOUG0WEVMAqgv
sznCwzbGY21q5McHinHOBZ9cRO5KCU3FXc75csbTGtrAVP/5Q3ASwuBi8TmkyHTnInbL2hly+r4r
0bbaDr46Sqwk5u0T6gsX5ZcYtUpQFrWG6/4IYZpiKVTiobw+pmQQ7LKbkgoxNsNcGeOyxVXJzF60
PbyVX7Ps2TWsxA10R1lP4/hD2Q32+TWBx4Z32+RLvlTpphwlfRpbTQxTqDrnt5IdP061v2H2PeuZ
xPPYO+ZGKZhTc8KBvLB9JfwPFBuPD4W9N44bemM6OQzv9x0o0INWLB8oQVwnhSVnIVSflo58kpy4
LErV003rK7S9Cgdh4Z4mC1uFv8oFprWwfw3nDWEUVs1WHMvU5wXxILyfJG2v/gx7dUW8eSz2avjM
VYRtEId+R03tbresMMxMIuy5Lx5W/ev9628meMAf2Gmf8U60zmKNQhxqGtjtunOSn8wsG9EX/SmU
WB9tHWUVdG9MIGh7j+3Y2ZHf2SjS5jWlx+IHkizeqHAz9VQOVkRuGCdvbSzIrZIrm+ibUy/U2yp+
dCSW/E5CNU+tGPrOcctP6cugMKV1YR18DTk6P9fcXH/Nhxd4B41Sar13VNJwosKZqvg5aSW3XORu
yL5jNYg14nCsH2dLodEmrKz1X8VrKyJRxRcWWK2wYDIyMgcE74uyjCHrBLtRYEv/STo9wn0tDnll
SR7tfff846V1gJfOF6FsaLaIdJRac39CbkFHlRywtKw4nKIElftTsS3ypqR0vnJe9HAByB7Bui44
GVV/zPDzf9QvW+NE79N1HLPomXwFjXM6p0S8qi15nypAkaRDQka6WuoWRt+kvULC9NQ5T58bpGBK
WY2VyH034DVmcgWcnngBB5Yo7sdCJjloWDFpO2YLs9/DzDh478tOMpzt/AJJQlMfu6ZPjR1fQhke
5zVhXuDMBqzHKlKnpaxsX44pV9DYT/HqlpJuaJzMqp1ALVE0ulho1ApIAhVxAqTq3QTr11UfrFz/
liHHXEZqfVzeCPa0jgxNz9Xl1RJ+6YR8FUIs7MC1NSZwdfVTVdqMUwrZfqN9MrUrleL8tQi1lTzf
FScTvNuy9aN2nZNuaFelilnP6tnkSKVYvTBgWcQ1Vp7uqyJAHH6nfaV/fmxexo2PwbULhUu8grFC
B8GGwFc8S6Zm1gMKIhhA+pFQgdWxqlJo8krz2c9lchJSEMAimIOmz7jNMthyyQtgYF06V4LhJs4f
AKupydqQGLcaFwB8QWoCGccS1DTCPI3HYpP+qzZnDUmowng/75C9nqdBByI884qflJxf0xpjAVDt
Qu0qmF9cv2nLksFGrpbWp+LZP/PWMlIEPXd9zohZ+HUdjClFBghZl6oMlbg/NSC4yQpzu/FvRZNN
Xuax2dhrlVb+x7XwVHoQc1JPjU29xIg1/B7R+oYVl6rvcmQNqjw6JvSrdoQCb+f3SEbpKhFWGEy7
Hv50dZrSt2/XhhyEIgPCDbj6EuJe5eybBPJBRObd7jTfSUlS3zMW2Zm4H379t5Z0yGTsGpfdT0c+
vBAMoOWDc6VeAx+NJN6dD1toj6b7QENiPe0r+Tu2IPTQId1Awm2+NINnPNpzjD+RoXTiPYA2PoFg
b+r5+zXGfWuyRDv1uaUTp5vmUPM3HPRPww/t+jjJFDC62Zi8mIB21r+qHsgjyderp1wkKhyOUgcE
oOZ2OxCa4KPsyz7F6nkHPkiIbnvnX9KYgkqGMaFy3sHqfjk/GnnbuocOh+JkLNDBbpfd2ARhwTbK
QPZTjoXyPnx6ia6orDKjd4M4W6w+ne0pTNOMQY4gKnXpx4JAaeEaeynsyMSke15IwrrtfYg//7PX
VelF+GR8zM6Mkt6KwNt3b8U1JBqmk9riPyFvtoiE6P17tsm/qTVyn64DNHG/HouXjv90LiqOZxg3
VKSHnYbVFQhWyGUcoA0LoWlsoBOkdlV6yhpNeSi7mOlbSlVvgn0gdR876wRrFSB6qHn9CPE8Lf2o
+b+8CN0e9rWd+f1ALnAaFN44mDnCgvdOy1au9W9qN3FyDBsYttwnV07wOGr3Rh5KGdAaIa9GvS1E
iQFExgTsJT0CPoLthsUY9/mUSKC0NEu4j7vcNVFjqwr4SWHe3o8CphGjUUlm66nr57DuXgVl/avs
r/u2X6SZ3cvwbQ8Bn0nB3o1JUSiN4ZGqwnaYnR8bALPo9e1gX0Lc60KHdkL+54u4AZZtDb83HJmx
uig0wH7fphCYac0bgFKW9zpmV0j19xqucWgvAL8vDBqSgjd4EZqdcgwu/Ga1nP5kKu2hJt+Jg3V3
s2uW2lp8eQwCz18fPHie10N+P/vf7zcRGfWgLCXITzKv5XMupQNg1KYPxxUBg8IS7FF6UPtVIxsu
t+rUQoaBARCuSOyryGXt5zT42YNO8uO08eL4Lr7Omt9DQBq7rxQgW9jbXswOjrH14ODLnVwDQpVD
R7FIfEPcR14mqs4e84vocVfvdLoinCAz7NYVD1PvFTHYNNMoeWfndnlpqJmKX9gDSSB39iUTiNTF
8UC68kUFrn9rbNSx1of+nVxC6Cftat4rJVgNKhPnoEMwL5lSH8/NsFlc9ML0EM47+kRDIrp9tX+C
WNXp1TwK/9icUSprZUuWkqBJlMm9+SGZ5Luevqg815On/mTYaVU+3a7BaMerGb4mR5tDC6oLgH+2
IkUpo6HLRLswtzk/PCvOrO88O74PAlfvq3zBGj8WdLSr0tpeX3Zhh7yK7JGCU5NfT8DkbMQxq679
A+Za2Y/ZtXDlKGon7AU2s9wGeQkZA+3J3PgOT3g+o8Zy/tOLH5q63OdPR4wYBm8tLzH+hpehO9Tw
/hHUxKch3c6OsW0HEQL8lAyDIIMKMStUyO3XwjeOsF9sl5onFJ0E8Vlcf5Qb7Ge7zhRN2XNpf/tg
OVxKG/92nKFJbNM+FAkbPnKFezvfiHiIwsGKiof8fmPs1l4WzjElADgWMA9SFGUplWiOPbK+LzHc
QWEggVElX5jJNo7o1K2RLppIYc0TUFDmgd3NvcoRKdp0iOgELQ90VAZxohpHexfY9jrS0MNEphth
E7b6XdmuFyb0N8bQbpA7CBLWWFsiX4sne2WL0H6sPZkwc0OwBfmtzv65CuxFmZotyOPZjbrKmR9w
1MKBz7NLzeF9lfr4QdDDod61ZGAbh0vJ159QacNMq7ZtiOUjKX8HBaPFKrtON2ehF9ZRI20iaHXV
l00XyfwD3FQFMRg9OEb20CFzSMhz9Gj4oHyQB6cTJ8JPLTS6L+SgVmW3uK+/wC/2klpC+9xqABE0
s1IGSq4JAEs/ySH3gYmEiOnWh96My64v1svVM/Ag2HS69CWbEG/WcL89mNVDhDVWK642guP01g8S
o2iZKx0stINfY/V7tmzUlPWB2lY0bHOuHjeL1f6EKxgOL+ppzoE4f5uUr7aZztB+uqT1NswrXqWn
ZVJ2a7Sn8SzflAfdfqzSgNVt1n4e8E+8C9CPwLVA0+ECgC/4QVTl9WyiPTGSetU5qFa4uY32i8FO
suLxsUUyDX5FiKuZzGsffsOUAxZI53FTTA7eP0xFa6eU4KP7T/9m60N5wc8QR3Wbc7yTsxtFvEGS
zs8yo1I3ok7oG9pVJN5u03Mp09jjTZOhQwLwhW9On0RxSiGEkhIdxnteYu7XHme7ux1lNtKm0L81
kc++/xX7Gh63AcPeZwowQyftxD/PbmjLQNvGBE6XtL/Pz8SgksGlDU1sZIH7H7JT5yNbkCoJE874
ZUyYuLqTZs7k/XFO8ChP+4JeP4xtO3HNkVl3csukUQSmPOIeCNNMtoEKK8G7tBIvS0gLoqWhyGNt
TwnAV2P0Keka1dCS7qjZje5G0xLlG4Vnsg/IihGhqQFVCUSxy9V5Hbpu1M4RuBPTYLraDkSsB6+M
xbQkrNR7qWO4k1Nw68TqtkAKRA+5uEA/ib2pGirSclC0mzX+ltSLntfnIiCXl/4fhVIlOfma4Uly
pZs9iXRrDG5w9+apW/WZheISaAlAAeumyL8mpe2ZI7drzZGvbbNkWJLgKJCnr4rp2ClZeWzOPcRx
eNewT7jHFCN953arQbSR5K0FWFVRS9N5+B0DfwjvchTKhe3+xzRs28Lta12/S8vRY9r2MxKhF3Db
c1rhhV9P/7m+NR1gyNkrr3Kpot/DviA8VpZzR5fmF+SSuclFdNJHgqAzo9q/ot8lkJGJ69iA/hty
DgGQwqpKs3+/2KlE0rhQXB5QWkz5sE18NFO5RFOaCxugGTJzGiQn4cW7ihMuJ1zPwvAEhkkm0XRl
w/w5qxJHusO8vau8O82L4WIYsa1+Qctj8uBkHw1XDzfOS+MljtuVthl5JE+e9JoTa81OgyVo5i/E
w70Ic3uG62zifypkXkbFVIk1QSdz9Uw166hIoQ0G8a1sNuAgH3gizN8RQyOrOZKJKpePKZrXp4Mf
lyDsT76zMuNifYxvnCZk0yIVxyAUKHWibB98dDbkoEqx6RpIuCBFhwVZAEEq4/K8nBUzgTqm1teo
fdwt2qBOMPtzHdouu2XyhQ8tnuTTqWNxl4z7D2GfDpIzrDJKVvNjEUsmVVg8GHJdHKQm2wRdekJ1
7igmQ464NR5e2dWUEJQDh5uR0Pv57QLLaLDuXiqYqxS8Gc3/f1Qsv20l9Cz/IU79zebBWqBGimj9
0OB7R9sxYPIqfRlPeNY+1w9pjtbXO/n6r0GVgzdhv/hxlwBPQqq3l++lDmzPB5gaLb7OEizILSRZ
Zbs49BLX81R1zSzVbbTdsRePPDb/7DCgMrIbWGyMEPpw0iuwZmlzRVIUblfoJvUnYOP0qXyfR/Jd
2sg3BsHFTy7NigcHSzuX56ZUog84ookvxsYm9I/bhkda6pmoxJfKNuQnjzuhMMyFk6yPDaLgIiZY
LenOMEaIHtfqHhmol7gkJbrkxohV2J2JpCRn0ICCZ1tq5L9qS7ZTThQ93vX9Wz++lx6bURqALMYA
MNtQ+azAKXJcCUPd9JNmQAasieNVMz1idfGSv9HTbJ1Ceav2D53NtohJE2sJGt8xheb+v1BD4Gjc
ulnKXSNKJxc8I+/neVnLdfb3Y9YsFAQ9IedLar+CdTwvTGUWzP146Mx1OYOmq9AjJV8Fsa4xiqIO
zPSbsl3j4Wzv4IrpVH2HI3hR385ZjrhSc/AffK4tQfLjPtwi7DFrVa3T6CB8GN365QWQ+UbEP+Cc
ZxxLgWL1m7Chn21rLT1/DkPIU15oHqbKoO86lQ5171Ox23RDvfgYn1WMR8YVN0qfKv2A9SLZu91G
sL3wm2nn1xE6EQgtIQx2C30EKzjUQ92xwQKzwD8bVYrCo5mBlLtCH5f9bAl9RV2hUCwaCfv6IvFT
cVyJZ9vmyeOLJeLRWZnfah7pbrxXqsjhgPmlIpFNx/qT4H43A9BVnFXZ4XsZDf9yF8C1ZertTkP4
xr23wG6GNHbvbYNAtMEdnYhOizSpnbCjA4vq3UwdcUigb6YG1gnhG/40VAqwR2GJaPXavWc+ZxLC
d1MISehGhIxUeKXiFJuc8tcvjvKtGD0PB9b4JeU++5iUdhXdDctI7yaspUkkAwUs9fmzyRJFpVgc
HOEeDAgkG5ugaJKi0M9row/5W67h++cA3CaSi+J5nNAttAPPGivTh3AhomB62kwFvvsoe/TZRzMx
+TofVdPR4m0rQB/YFASfddddOnc8CgDBlEnCzFlqPnZDVadDA4kAuridJyXY77jhEMNvFKUcLJAp
ZvUFgulIEnf+vU1VaHv49xdb7rJMiV6FTn6Z6Lx2GuQv8dF/4+WRT1VJlEYMJtBAGgAeMRO16/Xg
XgfcuXoARj7wSEhL3jpGVUoSB7vJkGZdorNjeESS6OP7VRLTaeOB+ginbXpg0bYReNXuj4YaEW/I
OwfREX/T+mDK8UQapMr/SmlbYWprZLfmnM88LvHqADKaWttndi5VYQawa6S3NNpTEEt051pC6pod
pIy/vZu1Cjctp5Z9BlBmyUpCIeIcoo/4qPP7AVlRYdp+7NZ2ZqXn6hJOIVPigzbIkF7qupOj7qYa
/q9wH9TvK9YQH5Q23C968bYycD/5wJpiH0iAeXkf6Az+2yjCNRVk/fl3LNdp0/Tf2fV7tAtwirCp
7Ygu/n2JxVPNF6AeE19y8A7mHBigJ/O3D6Rdn+kNVxHYlFsR025iQ7U96uh7A7ro6s+Ib26c32Ml
nBlRKjEG9M0SZMnHO+ywgrWiwwbUFprBPS0hiptDsSNHftfsz/00vn+oOvKmUy+98wHJPAT2iHKk
CSLBZ7Jjc7ZUV9vL3az1/8bgWodtDd7KLn8qvTsQFaJM375XGiRTV/br8elLuWThAHveAAbRzfij
Nbw6JxMnEA0+M6Jsbfk3zgHpD6YwrMJBOrX6QJvXZmAr1AMJCCTBl5ypDXftlBaJWhoNIzkR2eIy
sQtHaSLjSWR7mfg8wHIWmQ0cOJ1Z/lcU1BYS/8kHj03SKU5hWll8kBjcQveb/RnLZ/QI7JKVIDgq
GiaoFFxKqqAiRwqqTYGtisDiWviYTs4JHrhfbdtxYEfnhVA6oLuvo3+RpBriVHDhHuTKA5hFD3v3
RuZFQgnRBIL266cFtoRvyePQa05EJWicR1C6ohxz5yOKTHurLoOEYqczQtMmqqxqIIRa6duCI5pn
ippml4ZaxdzBr4WL4K3hfGusr28Kms5Cl4q2B7Vo1g4dqaFRxmwHvlU6E8nOW9lws/4rP3aTKsbQ
dDAIELZB+pqPaN1Fd4ILGcU3lvc7e953bmWWkBorkV7SvrXIojFYuu74sr/Ghq0LeV37EfuWS8s+
cRPzfv2I6lgqlIvTm/oVUFQCOK4xsa9gLNOy23017V61zrQQrhyuvHPSpds4q0ehBTk/8GNL93NH
5NfdW9Q85w3Sb7cuw9DRzYf3PT5fsHBnd+6Ow/Pmrh9+Y8Oz6YdfOxcuEQT/RRmgg0dFrOYW40Ka
aZjY7g79Yh4XJSR1xSiSHjGn5JlwScUdq+5tWjMG02AX+ZYH+BtoVU2VDPTkrYv5xUFPAn+QaCeZ
DoU4DakCgqm5ObLubeIXAKCU+XUdWPQTaTMe7jgBFrJkZIAtt7o8VQ6HagghjHwSLr/a/S0g0Re7
RE3+DjrkfXBduErN78KLhk+xfJx02SyGqipJZqwy8U8ZvmxtMXl54glFALeYiUcRlLFa5ogkYaua
jZ8ZMg5vyxu7U1EUYEDGvvGOK6t8sBQTh1hPK0NbBkgIW2OE9PYdK1KRFXxsGEVY1OKgV5Tvre/K
rCyOyLj+8EQRyIXrPsuo7Iwf2EhZBkpjDbCglFepurE+71oLgOy4ZXx+c9U3dZC0g864xs5jZLQK
AbLppFR+sANaebP5KjmqDrc+RmivPomug+8xzQiFhptFeFIAzZPYRruUL4CUMiJ+j3sWSEd0YfI1
QFToW3I7oBa0+KKVCf+C5rS2k0IdwkmmpQImo3aTzBFdSM9cpbiurRlYtLRITIt9NUzfHb+z4ZC6
eti3NO5zD/DDRmAuz9ZDHgYPMee2S7wYHa3ZKAcAOsEd/c8y6sgBvT4P/oGgmz0qCt814vPdT2Xs
hzpPwKv5vpBlT/rz0nD14iE9EX6ZnTD2gMLts2U3Uu9hSoXFXS0SM9+NvYaYy7PBYgAneQB2W5+z
tt8GXYhEB5RkOtL5MwoImGmMxsVhY9WQWBCT0a/7WiRMx7FYoZ+cBglNkEgyxDNPUL4g8uvQN2dh
1hNVToaAkl6P6mOT1N8hwWiI96WZXpBIXm0Zcq5+yvX3uNSR0n98NE8aYlyoyvCovwJYrPR5SXKX
i49kfEBJwzGLMf6oW/1reuN6ROQ4qrnUc+do//YwqRUdvEJKPGquHMFaW1VrHQXQAUAh0kZL65xC
iVRVy8gdUmwLqKvtn/tM+osyT6pTeNGVFBL6kFa9dRF5SDp4YXeNi+yGuCHtwQASezDOYVYqH8AQ
vx7X7nVMKqjCu/FejWq9aPC/GQlJPD3LqSgppslBbsUFbhghpSf010qYsUuZv5AIqtpHuQdPdKcI
OhdleDuduC7hsHPsFW7+N0ybhgWKPvOqIs2nuwFzsJfS/RZO0zcjh/ElYoYvx0cOgTUhnn5kwvCd
Ot1Ts0VPrJTqbE20+DgYNr5X06ZVA8LALE7jqtdfqfiGjr/0uYlVInbGN8d5k1F0Mil9fkN4Jx+E
CJAjmcQ4Sjt0Y9tUQgeRwClMRL3W3ADlkHTEFM2T3F3XqUtntxf6YeSugZmNZfa7GpoG4UzK5VC3
LNX55A02K3mjiXQHLh0QCa8hZ9JraDZIl7GzQPcIEqTPz01i6g2Tu7TpoaoLRtwc9w3NWU80reEZ
6bXkc+HF6gBWml505QrYrHy30758g8Uqe6H7FPy3SSyooF85f6c2kCHK3pHEeS4AVxaAJIFM60tZ
9THvV6AlIXoRoPIL/a2lNi7eMmSVwdVuKH9FLgTGU1cDy0UHe+6ewb/jchrphTr35VQgx1E/nOCu
sJoWdch8LJ0gz2kDy/PFz9yEHmY8tHl+eb8vHcjCneH/U3Ski31XAD7/boPIKzSRixfs2crcdmLI
35cP30rpsQIWcoNYhHHTioh+x3rzd856PZd09gQDkZI1LVyAsRLc09e/mNYL2Y8GBLxEvwIJcHPs
he73wAHQ9FUobVBqdIp0Po77H+zLj4tbz7Q1mh6OmCS/4NN1CTpedOqNI9s3CtXrvnaXUiuxUawZ
7a6HWZlvQG2kRf+KG1I+WJTrPewkNiKW8b3nxIOAJsugA//XQcjHyLBvRnrPPSZ0mhfctgkli2GK
tv0SBfyFneJqrQAWmYjDU8yJx/PdndhdKZNUlb17u+4poGIDJm1slTQY7VrRMtKaylG/oiT+7DF4
yiskYfWRV/6FEIoRcCpJt2PgP1OE0d79f/ZdMqrVRiRmJwoc/CGhiO9VryGk4hTtQlVM1ddvcVHn
v6xmoI1idsuW3mCJpmCfUbRO69ngShooPhjGbgS6hhsc8ejcgZVx7g==
`protect end_protected

