

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
qm+ahCoXbtCT96FlU7osNjp8Kf3rDAFQ8vMBTpaKgTo3EvHN1CM/XiHNcIsmMQ17hbL+pWxo5SQe
TeNJ1GZN0w==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
KB+ek3mkpx3N+ihSLNljgKYzWfCbUQKXGho6dSjrHEWrzL9W93J5UQjcPdLkP/4r8XQ5AjiJVm8G
O0+WgdiO6dbDdWggVe0UZIQ5qp9jotaT15XQQVVkD2rcK5wquost1xsRm7MTsEsCbzkhqKPM6ASZ
mpW7GzuYQ2vDPmY/r9U=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
5IFnCgXf/KjXBNbWCJPfF+u/Xe3PWCvLt3/lqQEWvv6nS2jJ8qz3O+bSiUUxyt/rlAZZm5DvQ41j
Vn2wE7il4mdux1L3DFueP8Ob6UEbh6yobetr8hrEOpbRcnmnH7rXtvR+yuK3psDEpqbW7d8GyDcy
T6jGK5xIsUceYrUwudt7lxYx4bLnzP6q2c6uLhkxaoLJTWJGh28se0dzlAMX/BnMMfjK0HDKD6kp
1VwH2Gj4iT7DvyBkDmISaH7LPSlLhe+ZmQMkilflhi03bS9w9ABaqs6v4fufe3/pEUeBrvl3gRH/
oCU4QtUwSf8qfFsWdX+C6Nn7mzOb0WSGIH22+A==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
BAf2bWZTeSaPIqnT3j5aNO9C6t5/rcfC+/QtvmxOirWtcQ57aHowXlt817D+9PTxe4qEx5CjzmUg
9oMYSESB8IK4XXnHzrwWEKN1a7YOhI72J3KxmNssnP6jdEMx0znih/oPMXJaAdPPRUXzSczvXVqf
S7AhrmorMi/7B7tc1xI=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
dVk9aS2pcwcb0BrWR4Sm4FSW8QQWqHH7xHbqUaQTDLyPydXvHmrmxiDqUJWu8AAmbDSnHtBnMo/b
vhz6TIedlqcgp9o49Jh0CEli94frA6kGx65vbdl7q0c/R9+UB+XDf9B8tq4xwdSd4Twx0zVa9WGD
lmNliqJyvFk+OMbS2OJJyBNqK6eZPVzKMFkUG0UJu6TERfYV2nuxVMsugR94X7JoKx+W2jEprOdB
UQVXsqhudTLpaKEQiNqzDCaBK0P3FekkJJMtZNaV6veO7wX6Us6tTDs6pxGysSo4e6tLocXysaO7
1blW1S7foypb+e5LTkDXsQjIPmjtBTMz3Y2yyQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 47328)
`protect data_block
PAl/McOmyjwhKu5souetcF/oPKgKvu37P4Sxi0Z8PmrqpIj+n4xKFpj7Qrz2aIkLWOlSvgQesCFC
tNnpdHApOOWd6QtKtnWSMNg2sBopoBzB+SdnEacyCp4WTyImBdmazOHaHaVLkpMBhuPYmYcisod+
a14YWI8GOfZYUM+zheyZVu8wEk8pMxkumUtTJnkZJO/qd/5cxWno8sIaQCY2umB0H6V3BSKNke3i
VGwsDVz8GQPQVUGi1nltgAortYmBdlikt30Oc2EFD/BsQuGKdXFNQkr4fLqpjhdEWm0hACnXxCz0
Kv1XbTPM8PF/SMMgPqlL9f9R4EDp+CZ861FqVGSnzWbI+6gqQjOu28cjYj2583p7vi0ZJtQgDlG3
qe1WEG0ReBQar82IAdKmfoRGN8FP9gkV6VaKzRXSWFocewUjqinRrtGsr4Ghsk4a92z5XJXR6mPf
4oZ121/eFzRk5FgFbPpfXusL+e7iELTgjSrzUmztDkXTuGsjV4ZptMCFvrhW3WUa5HhUHc/8xhC1
f6J47oNaTjCkuhUa8WJLsvB5QiWa9GU4Xo7aSpyq1o9j0AxNJLxLHU83Q1v+qp7wTYxiGVLWgiLR
/vZPkrgh3lXaaKV2dOXIw15yapNT2nDuGfhrOTZS5bu9z5imIVZ+5kSRfHu0Sc/44w8QHd5X9bQV
v24iLym2yA+WILHR1jKsxfvXmqJzqXbE4+TiIDzBJXF2gSraQAuUa/uCezfSFPzEheODiivwMZBb
X8rYtG+BnpubhLor6g3u02OTv0lRNS4UPkcChs9a8gogpOzA0B4SmrvB9jMRI0SJ8zRg1RcsnQ94
h/y/Id0BrMDcZsZmyx1QvOsXY5lwH8QWREFVmkIFADHgvc8Vmc6HAf+6LsHGKOyRyV8MUpOJFB0i
AVCgX4CejxsNgz9V5p5fes0si2Lk5G1JNAbvSOAmylOoyim/H06uFFIUqRXKBZV4VYJZeQhgZNdk
aSxR9+ldnKQ6E88/otYrfUvzDrzROzwj1UQOBhRwmUPckHascuKMrCkTF79KcxP0dMt2poy499nt
lMq4QcRIF4YBg+nyE1y4lXTNahx9nnd5GpIU2AQ2WDR/FJiXqAQnSCz30gYNxqn9QCPgnXb8j6oe
7KohrcwuuJyZxSWVYRRTdSVocehcynCMFQ2/dTaptq6reO3ni9piXe36SZW1rdoVdtXG5RRQHktS
tp2fDQGhdP/mSh37MqGf9M7i19C5QagNxUbYmdKXt908swe8X7tGbO/0oxAqY0H3fW6FIOKS3tVS
g4NH+NkeWdtRHtdqsm3NPuRXtMgPJF073XmtNi5SSSH9uAvp/AX9eQ5Xftl08O2/84YbK55O6v6R
LAsMwptUX30ntQyT7D1BCyT/5cYs5Eu+LaP8yqhdyuHxBmSOTNATiuXHfQ+/FITA6xREEKp4QS9f
FxsPXZTtbNqjGGRsFo+GGZ2t07f4Q5tEHgGkjym0kRAQB9/tshVXNsyXVv0Bq3gcoveZBWCmBszv
x6v87lez9eNCsSZDw+R1N2zimRvcn0duetFgHKlq5XuW0DzmiSxWEcuBBbpIndA5ij6A5feuXZF8
bmjjEHT+MCjVbt2VjGwLtLtx1iFOuF2DYmHzf/bOkPmBCUDAd/mV+1+IpDVXJmu4jrH0O/dnxp1S
+I602hXqOaBvC2GAox1XtLbJ08hb9BJIupOc1i5Lgw9NeqONEKxsL4/Ary360Fm1ET9qMDxfH9ds
Y3PO0MWcfLwOkdS4fhDCNPhDn2fSgj5P0GlDes1SMrMHbqhLvKByllp7ewvVREQyDxZ6Uu4KAuF6
HjTwK10mjY95IzAIzH4Xc1mzaXRHi64xcko9FDU5X0BEtKtdNwxJAGkYKSzxmMcYqq9hnh0RU+Ho
Q0HlYc4XsZo6QIREjCNxDto7u0SU66vGTE70fvJGDReFo5PUsKbLZg4FSE77VwnFU08WPTgaCJ0r
ze0GUkPn1xCLNtpKNxymPw601S/AipOuo9pKc7XYObnbwMr1j0QH9QV3r+xp8G7uLztHpMjf+uaJ
LyLIkvUSOw8154RuLxYnOlLTlcORGCQU7qGcYV3e/knM2o3exvz8+9axKrc1CsdD1+txKQw7kLRD
cUyvbUNgu3UsPpUFtD6QdrqNTeDsrqS9jamdqwAqLJ54dOs40Upi7MQrdv6q4SPgEs9JsnmHhGnA
vSbr0dFKHH4X0wUFP4Lb1S2weRRcR0Dwo0TzGE+NQgI4EcfV2n3BoJD/IUuDyz/Luz8lha97A+rI
0+u/pg6R1jWUIllvSHZ6xVH4UDXwErl3TVPA/JoUwpmcOQQ62tfHVxqgx+nc9GMLZ9TYpO5nj/hg
Tkww7S+OuLvJ5QE9/u4K9eyuF8C7Xm5GS64EFTF3HRBBc3Yz4gzvsdNfWnlsx4r10vZnm0+wMcrg
PTeCUN0/sBlBAoEQukf3EmEachOAS3xFv/p8MGDgmJbecO6WQU/8NrKE5XSQXn26v6uNZUxYKCIL
kBkiAx5ABMdKZRFet7wW0MGwGINXftWFm/QDMuOhdE72Mr/DzxJ4xce0KhXXId7mFTtEXTaJx3CG
0a82WMDTGAwEzwTgJGOsDdnEfRnNjlDuQulF7Ae5Kub+nKZbkaAYS6a2KHsdeGnLWu0dM4fabgvy
ykhvuM5WFBAZ5BuyH5bD7Fmd99o1YUpPfRm5iXbY3bbM+3j3bHIBSVahW4u/BExtCO0924QFlGns
1wyLhsrgFByobuf8JlwaLuk6BMy4DZwn6N8yMjjjhgmrSpGQruhlzgQv1TjCPJDLCWGCDaOy+0zU
FW7F0djdVy/HUvjeB3oET6OgJXPxDt9rJD1UahYVNxUeO6FdDgL5dkF/KSsYkjgciHmiqHKZsqVk
vjnCNbnVWCBl5iW+TmTdqbtgFRRGmrFn6AsQfrjavMduDk5PnzQR9UjbD9hmNGQxh+hmtIYaXmcv
3atk5D/KkSFx5bph7au9nJ7giezaBwzZLsBe0G9T5O8q7M7Yla7mFqst5fBlpwKEH3QSd4eeZIkG
J2mwgRNNddv/xp5BTHfLgV+Y5bUcnvcY/9Rdtxm21IR82pqy5cGRV0bbiGw9MK1OQgikvK/k1WsH
dQ58reccjbO6GDvdPLD9sSjBcPyghta4ApWqnpQTCdjNgxQFIR72Q3elO5oSgVEF7+sM5NAwEUFA
pRdCN3tuxVeT5r1auaqCVkaSh7dQb6PvK9D0ENycNKZpCPRdyGxODynlLVIKimwshr7XhoxAFi5v
WRjJxhHC9N5CYyzbwYbXEggsSWrLxRo5x1t9g/06/LMVmp5idIrhsZyjUScep69loGTMEatFCr4S
57FQdQRdtx5FBsLBDpGFmPcQvEV77MoEktR0GoqD28sYE2o7fvl6HG9xce6sVoKQT867X5KOdbjn
LwI6xf4gg7FPxd5KIg3wHLhy0HH63uY2hVb73J8jKkDvGRpsegHkU9U/dB8nTzkkLzUsln4K+4L3
2BcQ9jeZzhsb377L9wqFyKX3cWseqJZQebRETHV5xmo0dYbFwVOVwsIxZyK+RzqqJ4VPoWwuPdTa
7HAudtcJgWwGYuz8szyPnquVlfUW6Rp4aIvTdp9edzcim5HLcmdC5Ud73vX7eWFXu5nT8o9VYpSB
pwzSPKPycZkI4gma1aAFdMWQ7USwrzznnzgH3VnYEQeGIjkalOQZmWdwhAravUJOBQ3zaI0mggu3
Be7X4xoGBecSW83Br22PrbvXhyltcvPYzBtARdlKDV2zkDptleg3GbHu3M2bDiJxXgB/1adpN8dJ
Y1zgSReQJptl6d0MKrOIzlLVEGW3G5OV+W5q/eO+RNKYyarCYNyw3YRyC1CJ9fe17IbdNcpGU+iS
5afjRt/kcDi6O//Zv+CbEcl8er/9LzY+JYDQjKclf9jM89xHv2LfDxoAgTZ9N3pmC7L3FGNHPF9B
Of8xgC/Qjyhpm5AQmD+JwKl0JtL8bSbxGKDJN/Rys7RML4HseXTuXPdBF3jNjRZj1/cgvnc7a7oZ
EO2ogSKkkB01yLtt7FKl8183HZ2YM0Fqwr+oIfiNbafgIYu5zuiaKsw2wR1cIeNHLdRZh8CFibRm
fK3Q0VUzh6YpEi/KdpkN9lz6uCwmoZ3GA9jIMdp/QqmvfPu+IrVBa3At0btJmjrGzUZqhTiX+B9E
dUAgEpgFIk1vvoXfld0pcvlXMJvhRtySY2AR8EOx+bjhRvozmGDcJ2okY1W1lOvTALAAvGjspdSb
J8thSSjh0vQrBFs85a4sjrBE5OEuXEwnTNy/NwuG2ud5XgEw8zcP7gs18JMjf0zCPddxqFzGImOj
w+wuSbsQmNvNvbdE+MzrTJ0SFC2b6jlZfqSP/Nplwehvel4+9hviGIvPcA9KnozA4k1m6phuxMmK
QlDXefXgeoLdEOOtYPQAerw0LIDmH47Rnfm6QmUE0fCK2OZ/QV1HDd+R4Lb6aAOEMU+Dq16zOAzN
rARJDyLErra7httkwKELqFgpGWAMlg2os8rDyPYa7tzaqPjsciNI57F9lKFEeno/w3N6TS1R28VI
GLw86O2z46hIjlTFKj2riibHSkeFNcUW3+B7An4I2AkYPg9CoT5+u8wskWwRIrDoztpfz7sEM5MV
WrHlkVYk/AClWkdNhT9fq8ueh0wqOpw+dxc56NGiGYQa4ATTm5NdYJdz9QLIi8+6AOYe0gybiqDQ
/4e2obdLIbZgg5mB7/fTX+RjkzdJJeItzamvUhfokVjo6GFMWZ6bqoZdhZdCs8E87+mlP0sF4LxV
VvOJR2ClQhX48xIgAch6S55Z/Ybv5r6aCHWQ5KGIScD0vdOYPtINbg+Di0UfqVeZrFV5NWpdoBDf
sji9x9xN4+S7uqLPzhC9fcXiL6bU0HZ2wZNSnmUdZcpdgjIqHA1YrbiU0pAOw893n8sg5BfTKg2C
5xMb4Y6MoXPhlJqmwUBqga4Xy87aN6YJEywnwuCMEBS/9uTTSN52f0bp7j+uPjgHovx9A/EpQZ0E
czSFjffWQKH9C0kTr5lqrkHFbcUzwpbjrz8WVGGIcV68np3hZqjKVQpEP+WdLdVJdAE30RowQxMm
Z/mhZS3kMZhQ7l8XMg7yzdy3OQK72jaqVx8y1V86kCzASeUQ7BkDhE6v4Jshe25Yr6511n3PdYpB
BljknwQdpKolR96GXjRbSv8N5AExkAflK2t1nDghbZmd1Ex0+OP6Usa6YyP8UfY3WnpUC5mlz6cY
yH/oAbFJ7vdoR+QYROb4Zf3B/OFyZwaQ9wGfjivaOBSAUxQ4ZXpFdGKOtcr1vw8tbypuqKRBDMYY
2Ff/tn4lkLBiXjGBdRtZMQIYw9W41t/YEk7GKBQF0ch+1RaJ26AKJ2k7n6QWoYCUIFwUGew6TWJf
fP3WvAUa9JshMKpcPIrqJoNOuGIjCL4+yw9CTngisB+Lc2qqRwvD2LLMhb1vRpQNZ8MNpqFsJ+Rw
83QhZQultFZSOK8BlhCQp+sT7tdj6mZ0www/PWCNM+ssMoe5yqyFxmdjUjOo35/nUPlAhy90uR96
8tgsqxRDgQx+jfHLKdU0tQqI11LPt0IGPDz0GlbxtIlxGdvYBIdWG1yzBgcxzMADjXJZZ0Vju5Ma
RRtF+VOk5n0GrY2YOq593AZlVAog+wGngYgssni36yyW8qMLdqzv3JK+vCoWdq2mxiwNRFg+c91S
s/1RBFo0aRsNbb9G9u5sTAGRIV3rdHhcmc+kcLqa9MOraN+q0o7dwphwjqABy4aCJSInCLTMR5wj
U2iBVudlw6nfoNozQEgSY/2cNWqYr5e8ZlPCeg4gT+rePcvE+/Ty/u0Y6v9pZkVgRWzt6p31HoR6
svR+TnTzvACeldkPIaeGpVWpEHdOwIdtk7kb3QFmN9x0hs2HdkoP0gvEopBtoD8c0upyfEF+8Ss9
b8NEe1qtK8W2eRLxUeH+4gbE8HpqbUvhj998tpLQ3nPS4MPQ0vFbZZPQEuy4ZRrkWtaOOh0AqB6q
x2LqwIb8/7MiiOU6lALDiohqgCA1TssUTWa+AkloSencrTLYapLC9WkjvhjGzM05Kur/EqXa+6X1
uvox4a0jpBBYe9ksVmORv5uvn9GMkIyE4NHX8mnWg4AFHwCRz7jsVRwqS0D4/2hhFqvPUZap//rM
o55H147V2naHy4+8z8NbuQazEooZe0LK3ObUNvZ5SV13rI0EeFhFXJxsApQ6J0m6xbJxZa+RTR8p
bdeS/pyjTHZh+9c67sTRXJx0zqCaCoWdtuCD1xXtmpxWNceVnRtM3R7VcS+BxfUYqYU18BdlVY/m
ZTDNSP4R0AesBTH4wAMEROI9E2+A4wvOjb7Ot2jj5+iXEE5XTAonyx03lSGlCmpq89qc6Vks9fG2
Fc9eAUd10TB1prAZnZlJAg+DG33kW/BqBW1OSNM5yOOLJbUyHIj4/hfftKp3HKZGMDJruSf/tvSv
c8qo9qwb4WAzeRvfFnxOxL+xPSB9MxeTtyBQHQQfuLvv14SSGNzG9gn8D2zUz7R8odu4NaIV8DRx
l+teuBqw8quvJEd7yTCwYClGX2dCFcrIR/Ny02SNynVgS1k9vOr4GRkA4dKtQwxF4totVEv6yOBP
O8yv0WAUONy/lyLRT1FhuMyRtjfAxoOdkC4IoOoSzM5in9XztgZBNR63aexUhcU7zFXwlbZMqUNU
sOBY2JNSeZ/IUaYm+K/cA5Mn/FEQWRBqADPpzHTWvPADGEBZUfPMV3Yp0ecVA1UQsB7QGrhHl12t
tiM14yXeHsbVkvKidvPD2sSr1+2EqW9JviZdHJh9U74tYwy7RdEPP3jpwIkGZsmvc1pGqt8Nu9SE
iy1MON+VnvoQ4/cEpbWrlXijKu1NXsH+sjT0Oa636FaEw2ub7j0vWjqK8GJAwb9WVd51NkScIJeM
aZrYKo4+9+DKeOJMsads4AlXNGlrLmqsuLYk7x5DBOR3ohQttqWkboYwwTstO0MdBnBW48y0BLOq
Hiyc7K2MbIIGnNOCUyXHl4DKX5jEN1jLMWGFpAU/qnrmhrsMU4876JQky5Upi/KMUO4ubQB8ZHLn
U2S30BBGhNFcwMrabPcC8Z3F/ytrgdnX4ZYSjMrROzWyOaDPGC883FiZF3PEoikU85BoUF7y/feJ
/qoXc654lJih5mVeIv5vYVb6o2waZXhtJayr7oduKUwBDgIH3592MaELpu9dtC+RKbQX/8jHm0t/
QGJXLphTp+IWFIl3AHpP3mf0x6Agv9Tu+k7imlR3zdAQSTKhWGx/Jm6+OzF/crgOp296C6Uva1u3
j+YqEUaZ2CJ0pt8Fjl0oE9exwxHLAD31621jducH90AEuzjmgeE/hDhvGIwAOh4/s4oYvYGL+VWv
6Jq3QzrOmMXE4O3W5fKHcBHVemWWez9wi7IByUhXwmDgMiv+jKv5EpBST9z0hr26sXJ7iwHm/YTJ
7wiI9qKg4z3Rq5MQdXH546jNRjS+z2MJ/Nfp8Sw/Kb40G6wUJx8L/qtsh0BC1sZ4rxB0E1Qasdao
N/TM8vOa7xCxN8BBE2PHvWrtuHZKoJ62NphrqfJ7kB2JT4zm54Mihz2a12TBCHndgWKgCr2xtZGy
wYjeYR1YT+E1QSGhdgirQ7hT4ab6Mq6WrN4+N01rT8wmJKnTy3srIevE7OXGDD3+iTkwwQefAy3s
ILetLCxhV8gVwHOqo5dCAbPf3U+BQf1G8I1w3wSu4BB0irdTcXB4qW25SSj6KYGBaWX1N0HVncLM
BFebdjbcspqMpVxa9wEl7ASNM/h9cSExNyX35lRj5x2SYjZ6zMo1eDlFsya9sseP72eMPJM62ca+
BTOcJ1DMZIQnKtsMbZB7du28Ur577vH/dWThtnKwA/mw2Zj6SYgyD5RTouPORf6pVwFW4kyCzKJP
NQnvqmtf2uKpeU6YxBzjF//O4opkFnVHiTe4uByXJPJ6jO3aImv2rSzeJTocB7tPnlcCZKywo0Nw
M5ARBdJo/BLuxWJPShXtigQnVr7ONuny/Z4T2JchPKGW9hauSVidgq4WP4wH2yuprozy6S98Jrlj
z6Y9NHkAoJyKZKSw9b4dbUUvQb9hLqkpguHoZadDJpLT3GgjZIGwEC5+IFwZRJpIQYrWvejIQXP5
jJGAnECChwJuQ8WVj0Gl0kTJtrnoTBW0JlHgetiTcfV++ODSt8bO3YVSb/QMn63JJbVi30kI7yeJ
pEH4oYc1uG8Q4iun1idC8bl2lNDzkrUGBwg7cM9T9hz7v3oCAGSlbFZ4NzkkiW4hzTpCLBol70px
a0H9bZO4ExYbw4meJsyCh2ESA4y8BQaeWlMzBqmS1XkwyKc9xMhDOn21ugT8wdkqayj2d1vkVWpY
gg+oUflLODWDco/Xh+gBIrdm4DHR5zAz3I2EDniiB8EgHQoEh/JpkAU/Zp+e2vs5pdWvL6KKaBRD
BVmvT4g6VVsZ/9mdDW8iyPKmSIgfzH9OSdXAWuj50oBRWMuGtoYokSvH+YpxG7XwjEigg3H4aur/
WNAPM1kODpw8u6N5a/Q2ljTfDVikCM6M6k+PYToZeogSvcyMRiCMkMdDWPmuM3aLIHw+PqTxkr0n
wMQ1xmmJvJO+1cP+KGEhto85K3NdSnxQNX9/p4Ag5ietBPSqCzjINg5hJnKvZO7Ll5DDm5yjrlPY
xueiA6GAzaiCxQbwfP1Q31dlN1b1QkfD1GL/8VownOw6Lg0FZnRg35aENpT+SWyQvG6Hyoe6KdCh
SfjltfgAhJhoooDaCwwoM4kMeRdDDQg7IPYWb2NMvqOYdSVFkrsr8OvG3oT/8xAkF18syjhKy/G3
LpoVOlJh+nlV5rsoUcaPk0nv2fkHr5uDFEitN5plwStIOGo3wQY1/nNFsiZLF8YNIrA2K4YqfA9n
7pCPpN7qxB8qzrrE5mqlbKKF46BAHyVQ6RTaSDqlWA5vpy2ZB6iKtOwjwkoLw3GXIqz9d44G5XQ+
RKY7i+ui9D2JZXwQN158p5G5JvJ2gP8vByBG6Ilw0OpeIMUPk1ePL4v17GCDAKRAYr0RDhtRxd4p
mVBWQvjP7bWysJyRKHmv5vC8M4kgtwy27/1sr0tpysi1FmmgP8GXf8KjUEYln86s8HExIbP1LCya
boAIS8awA/dL0wx4RG8EpbkET8VRmQYL/vFwzUkDsWVPOPyleU9mqerwS4sy0p/UWCrw0LaD933W
6gwfvL/m6GWMNehyuNqqfeMUOTlflQuHOmSvkUV3e7xEJPbTCb1jQVyQwBITbnuwxDoS1rU7Bwlb
KCdyeUgC5JHUsh0rdvJVUgyEeAEUwkBxmrPW+5r7Cm20w8v1y09SIEhB5MNtuN3f0YSIQbXK4dh1
3lCBNGcmJNreTz1T5ibimhHR+qzFx7gIUZKW7fYHU1wkQPJ3h31rMBjtYv6olepFXJVXecx5/3lo
FPAVMLJ9mxOArf/2bFRmt3/Coa5riz1kVB8kzBtesZs+cFYamCNvO2w5SQ0q61OmUDXHuL2GLEwU
kcFKv4W7iJLi5hkbDsj8842bXa5AGojabmwjPSuh+gbjlsDQzNAswlQimX4qCl1N5l/11MqCl5dw
+V2vHC+O9dECNoT4/n1FqmU7Us5LCAqnyCAUwdh8wgb7mLHXrisGZyhsYV8StPKtgJvh1HzcSQ5J
aMIsbuMXRRkohyHw+fRTFY9BTnmLaRGfCWNSmWKA8rcqBFiCnuHuAZryZQZWvL0+6EXovA07mfVi
9KS/Q5TLrTLw+eAFAtPThgrCi6JQifnzBn4+8ObnmsKcHXF3Mf0v0cfctTSlO9PmzpeRSx6HQGUn
hBmZ6Nx7Li6rb0M4WIk6IpMUM/y9EFNihAKmwQ5Un8n966OB5amujWtkjoH8lgBSahiQIf7ybdXL
Z4RHjcnfVgXzMt/D+0hrsAsyysKkUya/DVVp96X3nV1fwtRrkTeQRJC+yn9dF6HK9FC3TzEyhF72
hxQodmJetlzxJ3Schz0YV/ncp2d/+tyhZ/VzOQgiIsoLnTXN+Y2XXrcZKe+SjbeyCvcYIm2NEotv
heaXN4R9SxbZLaPRjTmc4qPbHB4lw5u3TDJsSwWkOdcbVuI2aTD3dhZJlWKVOakroyh74I0QgDCq
YNynDEB0Ptz/HLNpBXSGT6rxISwqzcbe8P7QZbnUtt1sRQTrv2dBLm8eWj8a/8Vqn7rTDsaHOp2Q
N9ng8SR8CFzXper45LEjwaI5QCh/LlsBLD+DMD+Y6vXNeXEumgQKzpgSYvBsF5wKfbzbjjlUxVB8
h/M2ayMNdWd0Jhw4LGKxY6j/4gXK5NQNirm/ryGO/vsgy7W1T22sh/TGXMtttn6mETQatWWWKOYW
z/sVbE5WVPjmVKs6GHnT+oI5o0AdJLXGt84C0Yt66y7G5QItO8igx6Lrh5gVx/LyQQLLrGPXHKl0
KJ5T/BZxzfMFAKHtBq97i+dvcZeA1WL2RPeZGfUqIgh+s2kzqvLkfryKm5psfB0CKoxyvWE4ULFZ
4IBjmQVYlpxSIxwFI1j5W2JoUT9SVrTEfaoi5YLtRetFKCXLdG6Oo0CFZwt3AfDxysAPU4rZOSyG
3KcpkXmnC/qkbdXLYT/oKaRfiSa4HLoBIrf+oi6rPmBHaRBHux2p2CpQTqRz2IVcva9QmUe7RzFP
1z+ebEOoken4iwu/KfPcn/c+e4lqqxrT6S6OO0/aG3kfEggoAk6n2UR+AhKDLyTvfO9j3qEdQxMh
57WeUBqlXT4LXzEyYh6F2xkJAhaagWDgPFJNmjUYhP1jGL4MDcbANDRkNBEcxKVFHinP4C8qyuEu
1owUb1WtgglUNOgKdAlAVWjYtUglKMxeew5swvHGy2N8TLWq0B88VPaXIr6leEIMGCunHOZfOlwU
w0HHm7uosJg4BGA8hKD8L62n7c6Ny8P/6MKwDPQfpxacvEb/hKFn0742Dv0KzhUX1O3nb9Q5Bii7
CNLtWS3ABRgWTeQwyZz4thGcSRLQWHKzoYLXEPuyXCRhluh/a4nBt8DvSVjt7FoUyytqoEsCl9Jh
ai1V7m5T6Crh0xam7WMNFiHLTahUMsv3Fuo51x/Tjzj8wRFzEGy78DzhkCVN76UC3ysUCl3TklTX
bGAXnNKGG5FAfdiompnH92EPsOVTNYafFcCbvu3QkOO1xHTMSxzb8RO+8u0iLl95kjGu/drQcN7a
zqY2Cv6IqsH77XRy9WW9c1M/ohW84qO2Y7PpZvNRR47kpQECgTld7SP+NUtKBG/CiPuolDVxE6kX
Pirzw+ZobBtcx7JOzWvN+Rju2CSP7FKUqX81traM3UJEVCTNa+SH93ADgZQ4MxJqwLdANlMU4TeA
YEF3zce6/sFEwjL4R5rr4MTJixC/2eJea0PTtUYlgg1FQ/4gS1wB2Cnovq3CMO9YE5JBHvm7Jwfo
tfKfgMugRyrdodHPO/tbET3pHeA34b2CF4nZODj+MBfwFUBb9b4Y3AcL1/BcffteQCu6o6LEuCWE
MHkAHTwL/ZdxUJd5txXRv7zgSYU//aNIZrxaNdQJ+U2Teqa8K48EPH5WhdDoxVQ+CfmJ96kQHufU
QLZak3jhM3qqU/IU1YDJrxuYyH+eN+UX9pyb2Yha3ct6CR9N7sVAQ1HIrYOBOejlXqIsnTvfjWO1
raTm6/c3GUM3hb6nlkljGjQ+J9v1CzLMgTlwArEa8W67Z4FNcVEbrMHsi8Lc1HxknL11+JP6bFBZ
3UhOcJuFgEcNOBfsE0vzWRXlCQsZLcR9oEWfVkpa7b/42SbKjWQcrWoM+XTCkoRsYainrUECeVew
BQ/ynq6FunpOj3RbwaI/+bG7qgdwmAL/sEYOaJXTXiCWWznNwJsO+9eOZ33xSIEqM/ek2Kah2mFM
As7bXADTN1B+8kDirpZ6B1CA0pwWZ0lKJSnTFKe64KoA83Dh8YCTlzQL7kUZI+BDV1hOq/ZzipzA
Ozmt1/vuFDRcq7Jz8cfVsjLuy/5LxWPJPfzwmSuBHotMO7RW+mUsWItNNd7Dhha40deWVQO2e+/8
31M4hjab3eFwFVJwENIuUXnGOIjsEIYL39qPS6rOpHlCuCijCdv38ea+7K1B2ih4d8q0U69eHT6o
pLiFduo82E72w5bJSyrSKeTivGy1H0dvEor5Fmf+zdZvXg3KSkNSe77KhflOgm3T17lN7PBVuvYw
T8zQyRzY+MISIowupM1Vl44IvdlH9wGeqrUc3rj0zwuANuUXh7AVYpve99p3X7rI8fZBu6R1L3xk
S2Tupl8wr636MEmZHc4i/PRv1q3mjtTezoVclXG0F/yr/7asNg4ryyFkV8ee4YLOpaiq8E5v0fta
ksULqILALkAG61rW12iq+9xSToVgjZGzjpRU3Sa8Bzaywt0XgZBP+mjlHkzD03vkjv3jexrbIbYy
Z+eL6LLDXRzJg4tpPBWI25niLKQQnuQ41oS9PBfmymb94CGTEtdsL+4oTTYdFQ8+ZYhx8HECTVql
TAQJZaDM4O2r5phaB5V6XL+YvC9KauzGXDbr3H5t1v1tAyQWZsSe3vOskVXXQW4V+Nqydg799zxT
pZB4RTrlB/r1g6KM+Ci6rFD7ctj7Z7bI3syGiEcougfJk4of0r5W1Y/F8H0T2B1HVoywfIGQSSRh
aa2mt09E3K/uCUvGo+vvA9gNV8/MTHOQennpJeGOLvGZD92yIZpKjwVimMwfzmZW6BFYYaaXpgOk
hmLZ/oLXkqWWRPHogPZj3dK2TjEQek9EKD8GX4fJUvA/BlUvjYPSgZpd9kVBTxyLIk7H5EJMf0+l
QBXrlW69/GvNxhVJTr35K0Ps/HwnRTPcaSl7Nk9Aa9JsMTb4R5N9qd64JgydNJmJmylZtbtOO4Ui
AbmuJyiyq9vc30lbe/SMKhR1jxKFU8V+SDHQSZamFf2omLjEZu6h9XgrU0CfZ02BWRboG1Wz1dTR
j5MzhXjUTYRC4llQdY7+nx1urXcYPPmT6VQjvGckD85N5UgBjGEsQBG29cqjh1VMDeLbkNaiLEnu
L0w1e8Re45eW/qRHGq4Plvdg0sZUyTVNLEsUE0F2oiqqX3lp4M6fnWOb8zFoRMIT99kQu1ugShfw
2ou/DFUiVPVNST9mdJh3Lh6HYebTW0KdvV4cBJbCPmCHrbWSAilE6+mE1g5Qqj+asWGXfq7zenM0
cDRd7ENsUJy3WCcnyIbTNglj7vHgacsSTpm+Az9yFeFrdCqyuEwK8CTSYifNvWTyeYGYofi7GgVU
fnJ93KALsAxJgrEu6+lQHNSaBCVFdZwFzuepj66cW/WG5EMUHTjuVLKtXzccICJn+wPpE6IDuJTk
g5fvivQzY7dRqroQoadtlqQNbyEVNdnK/cGDePX4pkcMjllnBNNHFHxwWzZyr5TqGRdTLQVFHrLQ
xgDpt92r8Plqbd1qSTBpi9dXsJqyiZEVLsTQXK6UcZ38b3YIFmRS3U3+smUVR0UzaflqD2EDCaxz
QoA4zfqpabT+RGd+emTtE2dWkCnT81NuVFP/Ey0XnMNwKIcarA2kwvvt2WMzgPhbaybpx5/mgEgl
89IW8ysfik93MPU5A9yUbEND3jTlYoD4ucB8ENeJFTdSkOUH6SwBdaOB2ONXR1rTiMYD+OuvXxmr
kV0BiVSuMMw6peh7JS1HgyBHGaiRHKnvX6+mJO0+TPp39cmnNxE5sBPF5ZsqBxEW8LcftKHwye5/
gskw9IGxWe0CUoziItjhiVcw04+PzvWfW2hIQoKPhBagil/Xu0Aih8x6oqfPVgWuw0nQW0oCtVEZ
bt/Z7C83aSq+RDGXc+csp6+/6R3mvwTf/yBXP9uZ96Lax91jtrKR3DFUBnxkjIQ27TdQsElra3VY
XygH2JK/2n2tiaF7vWI0mLtrNbi+HAF2NY19kCa+FT7RGQ/dsPFvHpbv+Aqyw9PZ5PwfjhM/DiVN
q7JL/8ypaLW1IYbcEwRBlBoafu0rAdAUsUrZkTOlloGzd2GTP0XPC5R8uaW4dq/5fIpWjv6IaeeO
aOWJjOE3br7xcR8k41tjNcRFm9qPvbBdN7qJfCzaBFLoZ+sAoPeGXWm3kJ4QZb+4srv7MF7dE3xv
M2USkue3mwe9KWELCniOekTHXYCEt1T422icxegsd8rF44lgaltlfh4HBWygMLOLsRLA0SNnIeis
xBb4AXJ8Qf9eLuGD5OyGwhllX6IM8gf31n3jw1HihuGYlDGCYHlBKPbSDsGkISwSGVm0UFW/4ADv
xoHhjwIVbIVdaDs8S1xuVpzfHGH6ZiPWDrWGJw+AvJt2TZa/bKFo02jfDqi8QMoU9fZ2GSAegX4q
CJj9mv6FRJyi50tSMynzl0A2cSKVqWDXILIvYIa6PdH/N7WRNAQHZhhU4H75tXqHddX7+5tKTTOn
kCyGNnCa+cQB8tPpeN6cmstki16n/cVhIpIneuL6xPhu46XdspUX7lCQJjB66GbtRDATwlJMnes1
P/jJuvtTWI38kNcRvflA8VIcyS/qqF4BpfZT97nJ61Z/GKnv7smlpcUOvU/qWzPKQmtX03tyMeLx
WGwt0dNlBZ5rO2Ff7D2jPGGOvsSw/Jn0DDUxTJwCVH1ifDs+2ExQeOBjuO5NoCRSzjTxIRD7sEGS
cpIf4gUmFoFWdobfL9Utlqg8iZV7fLvhMX3/TjmFY7tusSfgoIZzI1fC5/otqw88lKb1UQpGeVJm
DH39Z+WbuAMdGRntInI8HfPuiBDpOJW5hCN6jNDBbpO/QGG01d74bzo8zBkHdPR5Bc5F2oq5LN6g
2ptcamWrmPtGSb4l+QEvK+SUbbTQcFOE++c0O9zPZuC+EbxCL0odmHr1dPFWgLYrzRiPvviAkicn
RIyS3VGC5tlmmAmcr93+uU2rd4IKehAkJbnruTPdTuw04m5+rULUxoRxywVTu9LWc1N3QJnr/pVN
TuU28apJ08+Jc8Hu7ZDia+9yLKU9Gkvwprz+x24KuLDFEN7QavqVzY1p0l8zE/BvgR/hRr8mFvIY
kLGt8jwsERoLXi/q0DwWGshthdAg8I1Sh0E7BHQi8QwX/KrDFDDkU2Tv+NMXZ+SLTQGLauBBLbbd
JKYW/hr4ODRaaqqswV4cWll0GXgsYzM3iwwjfifdrsUeNVlskV4OK1LDBplpgBwhWiLEssnTT2Nq
PPaOKCHMqwEoVkWoS0yaiHWOn+jSvcGhQshCN/Cs8rlFNRiMcHQVSMk4sgG2uAzmn2QLEQX8u/03
MV9w9Ttw9CDjF46X+C3vDoxpiRwHlKICnMsh1Zwm+oixCiCYfexVf7amDw9nzLkGHA5Of9lEJU3e
Xoj68ux8fzMpDHJkolcy0IAQAkaOwC8dTPx4zV7YSoZgoHpCc+ln7N45SGt4AIUJvBzvpIcOioNf
fxIROirhTcM4Qkx1eZZ4pidyG/VmkrbAv/b0FHBLKewFimY4J/vdiEXmdLZOxCgK0yrDmu2UhNm/
w34aWsM31l/+ltl/dvkAasfqlBMzVSji6di+Qjnpy5EmPaA1unsRtaMaOcPXniEprD07WtEsyzXm
JjQkRamL8JoBU4/Hfj2ouhR/rSfAIsumAeguDU02wmJNtDeWph1QZiD8rgHJjpczF/3QvljEgq27
HFCh2kBFk6VbgH2YxSj3mVvcml4jMpzyVFDUEeGF5g41n7AMkyMb+uD5qqCL2Vp/JbEfbglqjwfb
UFKvYESBnIwe+/+142x+xaKUHtIXY8Z3WbxZwHT8MicWqncYxJWSWzsPfdCxKRFivFav3hJJScTu
9sbwsS8tn+lpUyVGwN/rBObSMYwL9mXclYAebSkq6CVEZQu057/1NxzgprovxgO59Suw+EXAGFBs
fJPlmQVsg/hQshtSKu/EA0I7sn/9bmR0uKp/YVcd0Y3c9UQYBGvnPKTKl+q1u5l+eltBZTmGDFZc
fn2QfP0MQgKkEQGUQSjaGgQx1SPulizIQcr8Q2sJU55Pq0NKvXvMp0BBhao/ZlVZCRt0HcYRFfK6
+nF54IFusyp7YZhFGAjYGq6jazqWkKAsvwXGQMCBmwRXz0Q61OZCy4+hH6Ow7AJzGfdQ4z3zDRfV
yDj3b5V+bVtHYJga7mfqFG85XxaE7xjzByAgxfW3lpHRED2c4R3Ri+YRX1V2DgIsr5dBx5qYUPno
zp06bB2azI8nP0XfnhjAb4F7jl/OZBxaur8ixauWSHvp6HaZ0JHqAhD2Y62r3+9RSsaeBmZwfocB
3Ibme8dSvfRpHRRlL6jnotHk0oEZsgpJhXVjxBONU7ToWDGb/9caGHc4MsAlb+l42GEPsxY60HeJ
Kk0jKc3oxLzvZ7dOEoc6AlPfdn0HoHh2O/dELmA5kV0b6/qD1xst32MlM8g/P3sVfLQ/EW2FpapR
ikuKKfaQQbrE3r9zWAyQXeKoKNunfEbsI2iDdi39hlOUpzaT5KjRr6etZtW0dd0sEbBuoku66G2S
cWBQU9BJ1YasoZsNcuy7eIFqe5Zt4asHnrY8E2kiJ8EMOSHDBKWM+zBS+p0QxrJVAgL/9zmergQe
Nw/9D3zXT2b3kIDf++oWUv0b23X2PqOSkttT0yw/IgzC6Z11/dlS1xDs6Vp4wdtAFS9BTvWVfQF+
OSsrY6sOsNpL3gFimInZANKLcsXQmyy2YUgU72bvQLPJQEOFAIaqEC3YZI8JafNDrX9f3xbcZlad
FgrcCOdUgqKBBP5B4wkPtx31ZHjxssbiRES8nklp53tuAyGC/o86i7jmu+y5+1rOfofcKo80AeAK
DPKRV8YZ6lzhGxbXEEmnZ+Nz6kLK30SB+fiaQ5s7zz8P8hwb+K7RZNU2DDuytbTtRfuqr6vT3xE/
+By8/7svue7hkI9dTabqj3CK3NPKcZvgKWHe6vjRX5un9+Xo74bsIzU5Mf8DRXAGIIWB0jOp6aEE
M4PAW6z8VVkx/XkJkdTVUwG1Mpml+faON21FIqdd3WX3SVoz/RjjNIqqVhtm4QV5Bo/MifoVliHp
pgHdSzTVccqUWWgBB15DUFJAIlnFJXAZJCU4V0qL9cXPOSaKlgbxLBbsMh8RvtApsXUAY78Z+Q5z
gT7QKkJDmt10iX50BNYTzSwsg3rvzBuweRk6e5BvBLEYxan8wkHLpEcuQJkWtlz046I6xrJVGelG
sIVEHUSfBI4mb5RqMMtJFTH4xGGR18+cQOOvoa713+sVDo5nVY4o/Vkx2Z6szGGPx4ex4kmh59k/
nn4WAeN4Y0S8btUNXnZDxQn0me3K5atFYMepn3TCRHc06XJOgClXtBzBfETRf1zoaEyVA8kanSfH
uPhOWpsnizyFGAFMV/xL8w0OiKMxOI7olDli0AJMFpLw30/Yth6Z3EG1h5julvZh2Z+b/oZTX7Ks
7BM+YKWxgo840I6cd6qf1SLxiPIrzDnHWLJQif+fcHoS8xjf8KjdGpIB2BsTqKDZnqpJQZJjtJsn
/73D9VTNPLCT98CZO+mWOkiJIm849apOAdC+Hqe1sYUjyt8N1DieWrx7O3MsuSXQAyrJPHjLaOpp
vBMo+jDOmWXbNz7y50LS4tvrSCSbMiaR6EiJe/G1FjSU7WeH9UP7X6mblQI6WadTBo8/Hl8CXyxX
WN0P8Z3m/MFImkS9AQD9u5cSibQLGvmqMOhZnw0jEM2JsZvXutiQAyhpLOLfe5k+cRcmPcNu+264
WSyqbbE6nV8c7e7j+c4PCwKxmZ1nrJkcJ7+saJz+SDPX+mrSZx64tCGYtVQx7Q3FxI8oVN4PiVW/
6nIHAUJ/lFX+V4dSUjRNxEAmkA/wU0HneBONR5CE6vyxA+lzAczAKZHrgn9MjPgICNXNT1Y/6sjH
YA7aNJ73A8NH2vJUKxxARoND1c2LEDsgsh25dtTf0TN5qTwkiuuMQreUXZT+LAZ92msevWQuFaGR
xleU32GzdlYSlVE/Fospdbke7+fv+TconxwbUCiLFdE3ZdTU9xd3QDkinBD0WHBqG8+w9YmRoevV
bAwphHzbX0U/VCKqmtJYcvp4PGzWaRf8aFte86ts1TTP60949Q6sg/OvZJDz83FOm5Xw7H9w6IkF
yWWkBuRrLNxFXSabC59sZtn4M60cjHHaGK9JehM35VlXVwJJtPwZaRm17vU7y21gR9brhcFzWGOf
OM6fp6SiqNLKF4ao7WVCBI4pSOidVQZ/VCPTaoV7zjxTKstKvEZ+7qhHjyAal7q5tU6AALdcKxt/
sJz8r+vEtKZ9nCRqFEWBxzLUD8u0uQt7yPqITsG+YU6gI0SUzYNL1KQU08ICFd2Xaoeg1MmaBuu3
97WcgrkWTfoH4P/OmMU24tF/AP/njFelhqw1Zrui00cIL/yf8Jzl0/oy8fA9bEW6qtlirN7E1+EC
W4+KKjiTb1AzgdCjJK7WdAhNMsZLWQSjr+gABC+PdLtYYHW23ivaJSD4UgbFFcUbWXUiy0YNA6cd
OvIxwnMg2LVG0NRc0gUCLPuXkkntZHNSbkVmXDIYQslbwyGEq6Ig9+Mw4ZiseD1h5DCvFZ5H0A7i
B9AiIPu2bTQJnMzzOm+xFceRtdNncULi2Q/8I6xiwIeDW+OW7ykwLvZJaQ6nm/ocXXMlxkdx5J0D
6oDanALjYdQ7RhQOq5/gOq/t06KddwqCNYVYL7Vqp/vZfOBq3JJb4C3LBioXN7g881z2QYxoKIZz
sSQ87kMmQI11DyK7DQvwLprovUx+XyLzpw80UGqrFpOJG8xM3RwT/0F8ozytKfRNMWoJjoYuo128
c3atMl/kBYGFirqjxs985leGWCKXpD6CsHGkGp0kSaXuCXBTrr+TCvipSsvmTDBPCJgQyZ+NgpIU
RKatb7Rjv8PMo5RTfOGO9WDhTih/22FXA0ByH2jq+uqTNmfNsmjxhY8iRtfDXboLDJfLkrCPIT54
USv4FQB+Nu0WHudUcBvmrH6WyYJVPfUKtgInCtIVFyAQ7Yyt77mMwpJLonG+YV0It9jGVhUFeV2J
49e3jpBGMO95B0Z2+ytj7yQl5g1DM/ghgD96l8cmbNb0kBRRm4ycNvIW3BhG0yPQvXFEfsJLZpVW
Nyso1Lqe6g2/9J64oHqdrvm/Y9W/2cupKsBlutOeLMKkqUiJ0b7Tl//WTON5eepcnYlalrAMWpMV
N2dQfvOf+0nBp/Al5Fvgz3jPwYwNDiMt9SkaU2pbiX2nrluTr5BCCXyergNY+mrDVEJaheLImBES
rX+dzCkHg4QimH8vfVlh3FjDH9z2U9HHwR/5J2k9q9ia2Y29fHStSJUFwrKPqkjnvpoVRWakFoHv
ktowfWAvM+sgzmFbb7VhxdO+We4q5ocT8vWTqhou+FPoL1m81+RnbYCnmVq3AIv4v68hwcmtHX6T
Yas80y93q/OW8i9xoWXhEUfGEChUJh6/HQ+23dgUq5aRgtJtHSgtTMbWb2HQMcI9teMpmAouct8z
Tgg8xiDcgKQoNtBxBgQU1p7omWpOyMAbFRH5FxoZrAtTdUHTa+htbfzLZTDxNeMhUbgnbmGjnb9S
+6q0+UyW2CH6kqB5l8YHeFk9sODPKL/MqSrwH6TMM3voBeuqJjOdYGQJn6s/a7H7TypLTph49nsx
TRP8QbJSVEh9hY1lqNeSD+icrcT+6O/oTl7dtTQ0Wfi36d8sgc5CEiT08JYjapVRNsn65jvK4vjJ
m5J6E/aZ/fFRn9kkXp9Zgkvt5thXtmIn8XtM7J8d9QB7v5iXPN5P+JnEV/NcT0kj9mi8iWJkZ7o/
X0VrlS2zzJolBRnOPYG6SQqeo0hlAW6i5xdalau4RkXPPWciXvarWRfkiPq7sr4hW37IUwlvjdjN
f0FLvHAzeunexSSzNWV4Y083+xjZy5eawSdT95nk3s3UjBWnVyRpvt3Yau57UvYkM7XHgrbXgLcV
eGsDN4T4fLh41bjbvzWeV3bZSNK1nBE/g+ewXStRgVkL1mplEohQFazjLvoV1MsyArg2cZfrN/cn
sUk6UuOLWHcy+QWSOuIVUbu1pIU+UcuZ+E4pK59igsCxpfrFjy63DC6oAJzTb7zopo4SFr9IGjo1
WnMANfpTZgUzgJvlqLUakq65TYM6iVjJ3hxzmqC8SzwhtFp6YtqBVlqsXwH1sLkblkOHp/GZLyAJ
G0dRV+14IdrhanMWyzlZdbg9faKHvvZZuDytuuGXAgvrJKeH6/VQmFuDPmEiL/MKqW+yBHBSFd+m
LeT4l+IEah+j00JV+gYb/XOUua94IDkSOjS1AfZSXNl1S+Wk/gHhmxvN75CsX/J7gv+b5EbAMT7i
/sTeIIUYst+xmRpEyeOxdv1a2m+CZdgyQtKpOQ91I9QtZOJyFiw2vGbQkLcIWDKmkB46hDqrzR49
RP3alcU73iT93zd0vHsCAfYsNEllUAGdwtGzGTmzZH8f7SQad/Pnp16NITg7bwNMGShPJaHk1mL6
M/qmC2UAvIV/w2qF+lMNtdOj8XVTWJeKaK5slJCxAjJ8ethi9uI0FDbswzUwXJG+Ot319IlbDH8o
NfpgCI2GRDsvimb4TiTFb+da7wMhkYlO4Y6nwSFd4oUKPDdMvyeFmH5jo+47UlalBtuzJe6eiY5/
fZEuVGbx6HcFgDlN48w8SWIi1yZGGe8hmvnUnpA1qP/RIi5JdWlwm4OEp5DT6dvAjYQRlnQnRY2O
PeoWeIK1liwstPf0ZLChpkQujNZla2QO/bmtuK6VlxesH//Disi5YIKzve4SN45B+87m63B6+J1r
JkHSPZQE/+egCZnjCWi7wmQ2OkxxAawGX2SXIlRLbwC+qWilOAqInJ0qZXJdNYd+20WPg/IPltvv
53Vl/do31VjQvwZL5kLGgCj2dW4zvDLJwZnSB5GYXhRg/WMj1EROWij4YVn8ChbCeP+hmATyZQEa
cXVD4D1/PVuGnlL/qF6Wa2uOPIKQe9RkEkq0rzu8DphxM1obb+mOn2OsLrKadRpFZ6K78Ezo527w
xCtedS+4c4w3mL8NbcqezEythQPT4dsgmHkvHIuIiuwQEki7T0f3jWr/niHC9qRuEsBPSUgJ7mqU
PXawrjjOYs/ovrRpQZaDpF7PEVF8ymRwfNFGoefGYqRfWPYnR5+FrdFiqaVUjvAhxO4JEd+5I8T5
0UmIRDFByaCXhYSZ2gs3wCj4m9HC31VhZ/JjSlT2Ak25P7jya9uoGv7a5CdErgDkGU34hafePFPQ
fyQM9tR7lAcFg9LE1fahfjeebMQMd7JjpWg/dx2ZFYmac3QBJaC6Uc72+hClcAnxeQGhbKB99LLw
mmizYVWBbkdYsJk+Nx/329MFyjzii1T8byD5AooXWaujOkZs4GN6fHvQuTAbGqOjSQf2LpZbJO2a
dOBQxtdtrKnJ9TzEuaKXspNkmhPFCkhojJU0Ce+gdgLk4v5DL6eVkUVx1JVVBOqPJWRnBb6WX/uc
d5NOTzTvnyciOaqrdArzUE2+AprTp/0iqZLjs3LkPyg3huF+OW+YMkupFWczAyBjgMbxRWVDXrQk
ieZQnnwXimFjm4usPdzEQkUEAe0ZBlUujJDA+2BZUDJ/aPpbMd5kJbqniIGOAg3rNN6LUKq7XKjY
/BtyTKJGZ1+op0h8QrHhUu7F5qMBQiFEBvIruDC919Ga+JQ5jdSrhtMmjSDKMZc7vubqZCao9QTs
769UnNaAVP06i5+nPI8JJIr8+FFdVa4Jahh5UEd8zAd8rVgeHtToKRxqOCFqgJ/xKw7IfeL58hbU
sFiHkkan6TnLslAmhZQ5FDCvELirv9DUS4eNgx89qHqf5hDia5KXvoQ/JCW8M+BdLEabnxwqx9HM
Q4NbfifGKHdDijVlbjbf5IYtAkJ2zUCLKQ0OqusiHXDm6E9x75iw68qXQOWXO/ZRJdUY/LvpAWem
CFj42tOM2t+6Xqkq1euQJU3F9BK42klaD9NNkPnkA9PEXYCV81+h1ZHggBOMyAsPPrbN7qXxfl9n
imYs+IDMcFRMifSIpKqQvQEmNoUwuzjD++ClkTgd0vK2JiaEIjSn2zR1ZUtMOBab3dwRW4z14Ry2
RliB3f1YenBtIYldWa5jDzFL8icOYaaClJ8EpxpRn+G1/XVR3RJkKmLM9kMihZQVJPwDNHMGhvMS
1+4G/Hl1IS3x3s5JPuXgLBQv797porLEkIi2fy1+URIGMA8Uz0E5FpmfRDBFhmUAbKtVGTROZxq8
Ku4dGpD62xlb2buQk8TRqAgMw32xK0Ob4jkTbB7E4wO/9r86eGwQ9oGgHVAVYH9RktQbkpnjEe8d
+J3PY6391ocN4vF0khZ+mvUPxUjoEbWbIOGtO6+pRHla8P+D5u2BHTyI6YA4TgmDvTFZoNKHd0fn
m97pcAhWaNbbqb6tc95GZ/Ba4VIPQw2osHKW7UCpJw4e1Op/DKFQXqLcsTTuAmtO+4nc2rKTVqLP
jD4z9dlAty7DoKDXZTT8r/qsJP/j3dXN3DqLuN7XhpzCPENNUd2x9q1PDp1LIh5gWGxaKZIFQX1a
uCXuwnWQXFyJKHI2TAC8gZQJmQ3zxT8J5O9sWzEO1pMS96OfSqD/+jGhB9TmZMZs+/RZxjv9vAQi
gHtTOKSJhmWdGI+TGG6Buf4WZTtz48N+yodO6eg/iAhp5ReTXxqKuC8xoJG7HBIGUkEGNSrS40vS
qZ73jFe9EJZPSkDC6eBO9mZIqzs3kwXSWolvx/4mLVs+yjbifPKgtv1tXt8qlEGYsHQJr4R/4pky
s2nGqA7CRLTdvavOgpTsGkgTZ30+cvFYSIKLBcUWO/N7CO0rW/y2lw1a5gu3PNcEJpl+KyCbsNsT
YxxVYskmbhverpUvHXEgkJ0R8wrD/wXiROYH1DAsyQxpnlIKrfqMiFoViwQeGWoY0RO17OEvpHYo
qAe9diOVLGqJ1/Y67SY/Ogl0OSVKXwhBdnTSpnV9tkxg32MfK3t0dA89cXwIjKm3ywoLhJ9piaPY
/vXAzQwnTgi+OrndRdATFIEyqKvAvzXFmV7vn7t1Gt0+b1erbXTzTfTIqgM5ShajF6j8hs6/jkpE
0Hgo1A3uhxL9+/njqaNDxocrRjMLFhulEeDHvUUMQbVY6kRHF1n7QLshWUPdKY4mONZFVtjrY+3u
OKNFmy3k/42892Ygte7WTFku16ttC+NoHW16ipW3rWp4iPKDyS/YudjIvU+UXaL4xGTmp3C9hKfV
NCQCtUBVscs1rJarrNV/WwvS6IounvvyiKoa3uDvyGmTQAys2p4K/iJiP5SESBEcnx/0Bov+t/2y
lVL8GNTTIjFelbbjkaXb2V7xhaKsJVzLZ3hqSlvYYkcMRXTWZQ1zIuq1Sa2lvVmKzzBM/odAJ+du
RNZef0oCQLIqUBN8C4UedPv83BLmOAHOmovP19nW+viYd8y2jFzasWrPa+9JbfPtrgj6FtkTcFJE
cJKyJWsYg3Ze3RIkha88z7/dFRpNqApbe5o6Y04WDuL32ZjbjUqW/v3bOML4BxGMRv1p3IZoDmNj
vfkjYDRJM4SXZk0xCFg9cNHwBPPSCNKhcXCtLJULQH8q4RWujvzhhIHNYU+qYevk41vS7B6rA5bv
tP4u4RzwjId53m/s0SkkKRgvYppY+FCnYIh7cQ+Dis96VuypEPXIed/jwqpkGijUWwfLW1d0oaqv
9d3FXnrtSSH0eVcG9oTbVtbdShusfwu4dYeYvtiKw8PSVq+SXivSbvfJ5axOdYLy3qi++Vfzb3Js
Td0eBllYNyFjARua5TullAEdttvFXOP5SwKqX2duZpZLfCJe+Ifgl4QjsX61216aOCdEiEoLg2Pn
+xkfFA6NUeKXCKzIlY9ZG7FZs4qy5p7Gh2EPpg+ojYyqsFHLd2n00Iy78T25/mYwJQ837o/u6mkV
c4zbWxhcNIkwXBMHNqbv02LSUU9GlEKpC+HkgRJT/Acs+tAaxncTu2PnmtMY2X5Ac5NKhEMrlUni
DBLyZQN6Eo/rpLd0kWamg4JQQpyPjPggMN70912QOCft5D+W32eIpC6ngHbR5pS2KrGSEmOjnDCy
31P7MSbgrRDf48VpoyxjUyuZ7x28bPVlxPpS40hHVzEZGJen0jqJ3vzxMIrChgcitWCsnsimkv/2
6nOCFGP1yCfpHn8REtBDAly2hY2NswSikvgN/Ej2YaANwoW+zsqF7mzUx++evvDJHXfZgnFrIp59
5SmQ9ncPgroYjGRvB66gA6Cw5hVRbVwyMnb0TFnehIcegj5EH1qQeRBvSxBYbHPpIPIA+ST0SlYH
2WbAFAb4CFEqG5e7Fj7bCaIAY4OUmRI8bkfIx9xb6E9AViOarELBxiAUHchIq/pEM+48f2ueWLRi
gVxL55fbyQVVXnYfwubyBr6weSWHS1cNOikkvZcEEihWchyKBcb4JhfZh+oJwhAAJ/KMIVd5/FXu
CzMFzLbYeexVRJOCD3DzCGbE4oFdlB6stpGriBymLrHsJp5jZX+qpTdd3LvzkUeBBBwPjCBjDZz5
DWLrW+1I798L0EC1v3KW/oCOscp+rljYZQ7brKyZCtFX60OOMR4Y3oePo3tMycKxXub+aSPbbnZT
9UOX0J3RW0fH3HHeCOM3nmZ0eHEtzrxYqdmqxQlehnSVMIJDciIIXnbyRdtoW4KZIDDwmJS6FhJU
qBhay3wCGeg4aN1HYzeF4YmD26KoI3tJFoYIS4E2yX/S+lC+FUTZK90pnssozhjBKgiQqX6N88sJ
16QWV0GRqXMvkCFz+Gue/KVgXqZVYbyyQPtK2T3JN4caJes5AXqa+ZMeb3GE37pcaNXKVysI8iGs
dDTpgKoyZObFgikX4G05QH7TAamonRsQcoC6iawKzGRVND+Jk1VQ7QRQh6nEhZro7xb415P1LBLa
cAwae0bztUOMnLdbZ8YnW+FImnKNpLNQ6hMJB8fw44Cj+XlYsAX5wYcGmGSoW2uUWhN+nAPFiTUC
DRgq7gT9HpSPSQXYzTBID9KPfEd23VTMr/ox35Nk56oS/REY/BF+fXFVwBJxA5YEua5R46HD3rfb
ILerI/IZiyRJC9QK54YRLmhSriRD8Xgfq73hovCLkpOTSCzBzXH11NUvU+a+n0v1wQQpiPFxsrep
Yy0me7iNXqGQW5wMip9v7k8h4raO+/PCbXQ5KzklFwCpfoSMkIcXyfAd5+h5Fy33KFpqvB8lvuwO
Kxri/g89Hm1twj//DVmkLv0AFzGqDntDnEl8VrrpkH5HrA6zPPesZNk1SyirBAokSwcvAGK62p1t
jy29EAKSgPapi0VSqFx3uJlvF90rzGU86ZlML/ZViUFPpmz6bjZhQpJAUgLh0Fkw2ktZvkSrJ8hZ
2y2sYX+744NIlbYhFnZgcJC6HEFx7JM+xai8yN/FwqDJ8jqtbeM4xlIIA1eA28K1qcpoBqbMng9V
Hq8quAgx7zzRWDY6ZR4MRoECEu2v665sYobFq4SVY+izn2opwkoR3/idTufUfAXk2CBvTYpQ8tt7
Bnch3dRWhGXwtzfWnllN0psENJ99+ClTO6ejQOiWPtZnk2AZ2txaTrdHdbnHR491lWDoV5hVrwcR
THc+DC/RtHvmXQQ3RK8sYXVBj/Nm/R0Q+Gpd8+TZ2ef9PBaN43GVKUFtlTwRI5EZt8a9rojEkLht
BhWaPIXvrPQPvYHqvYNswP68g2OeFPMIVLLGQSRj70i17ZuFNwo4+JYD/eE4oThGqY7hhVJFqKa3
tzjJ52LvkMHhs/M6WgUb0BpfB3D6Ot5S4Sg+OthhEnIXT7qC+pxy8wWrLNDX8eFfd6jON1y0cowB
segN506WQYMENqS2cnLKPw+VKvTfj/IQWhwjg+O1J6r24PpcJrqbjGs6uVKn5z0YAi7h229BSfRb
jbshdA682Vuv9uCM4PE7JNFE8grVKdKx8l09FTmKn6QesfZleLm0z/6AWBz5u4UM/8Y7VUsKpxHi
mCFPYMRwAzPsxX/g5q4TiHyy5rRABbnolETVn67A21CE9EEcyShJxkCr4Ral1N/VsI6SqMekocDJ
T9kx0prR0mLHE+toF4dg4SGQTZdvkS9BTVErwOquu/4b74+BUB4ULsXGNVvndfV9PpOjs8qFD37M
JmGoNhyQZH9g/CJEQvr63JJWmdIcc8d9hDCy6/OM448DByFAAROxO+zP9F7tHuoAR7JrInxh1dt2
r6cMwpzw9X4b24Hep6PYci9fTGMdUu2Bz4aYbHjHV88kUkjKgi5RtG5iSoUs0VRAMdBTn9mRviRI
RjLepeqSMA+yOBonuOFUVErzJQbxQ4Fn5VKzuFcKwh/p18jw9G0tcW4lYTgWTAJWgidv9R2M51Jw
YLdDrDnOpZ7G5y8sZgChQUiLLhW4k6pC/yXGpq8XADNdLOCkVjziimVqMSJVDe4qTK/U9lM2MYvc
lxM/ZmGzNIlwv1BYyngoklQ16Yj/M+oGBDfJhrwDSCrY7xGqsIDGeib3SJcuqvSAQomySJoMfJxu
dOUd0iSdyHTxfvhQRI6w6EJ8Cq3Z5SUpC474JZcE90Woq1N0oa0mPlFjdPoa3u3ft7g2VZfPz/El
sHmTLb2kmgeRIVUmj5hM/hD70KrUpG0lHK1vtD+ylqRzcFPCi1cPsTVqcP4eXpzJbUWFhmLGRhCS
Js6k4nyk6OnSzG5Gq651KLPUOT/WHHJBoFSAk0xSTU8hn7v/VOEBfVLZS+VYpYzGo7t0pIaTdxNF
9K0/XHaEKlLZNdmCp5UCQcRa696le1LaNH15OIwWN2ccdtl4LiV/HliWmq2FZMo9R4R/iy9l7oS2
lFdHv6LKlX62Tt6gF+D5DZwHpGko1oPrt8S+G24U/7gLHQZ5caQiyswamTJyjtYvEklykSN33yT3
sj7BCrdJabmDtGM4+KlhU9zW66yNBiQPH4GxV3h+ZKo4eZSJ6c7BzF5woN/hMGm76MWaLTTYuT96
SChMVZe+SsOPpkGkbeaO/wibH2V1UC1TKPjVi+juYIrBN9mL+56DUIJZAWbBd9mRuZMWNK6mU7AE
L3ZflD18lCM0SN5tet2THc0G/Uf/FklK5L4hL3pJSKgqWNNuq/MVsZIAh14eHQGNt/BR9NomShEM
DGCGVHdLXjCInyGJjUpsuwBdGMZS5D4D9Id4tZVA9gfOvtzlKZ4gCCuwL+yMUED7g/iOYwwxjzO8
PeefFmes8RrShhD0Rg0ZNY+jP4VDCtCPfV7dt9i3wHno3qKB5Yz9hnjUXAGpHCoWpK+dlW3LNfBd
ItLwBwPGikFKiuSyGNt0uJTdr0p+O4VikV5QGTa3e3UXn6NS/6r7Yyqf2Jz0eNLwXBnawYxs74ix
fNcs6Z3ATDJ4y343MR8TZkVk+ewR70JTkY7em/d/ma4jraOkoYaIfCvtYALh4bWSJzJpz9UCOcAG
KkXC8/1f9v/rhbfhw/Jfjfj8teX+dj1f4lgHpb3Xee+P2/+AtK0AL0juOWMXoF4TEkCOk+KyuShI
JaBASPhdgNgNx62L8Tit6++8w7a1MeBz7SH/9JlNeYGLk+4dyta7fD1ghp2xeO1QfDfiDIqwNE16
qug77bYiBJyqEy+Y8qplQMGuiFgP2gyrpIvkyqu79ByT08fPce5MQ1meEaR8fdH8tyrkSHY5qqat
+uF8yU9FSG6sE6uxIS+3huJxOzyTZEWpXv44UmljP7jztuOW8e/+1h5VmOWsKXZ6NQBrbytscfOQ
dChYciAHEtfM8cVAZfNENGwhS9koPJ8wiOpQ804eX8l/bJexvAcZxs40VNwiggAG3Iypp4wQ5B/6
CJ1phQrM9cV7RKOyquScPn3wILQXR9UMeKYNXf9bkE7buykQ18yFhYp4RrpQLBZQ3u7tQg738n2n
+bak1MslS7Zc7gaUWv1k7/ErEB+6YQsoF52aaRPYPJh1e4IroD9NJoQtZ/uyoRdRnKVcfjPyd4O/
k8vUj+J5fm/sgsiL0i9BQkMCSk1o7OPefAR0INYwOJcnpK0ZGHzbZupwXaP62ZxYw0ixDkXC40m5
GgL0sx3OMbuwT7JHPdcNN1/YDFwV+6UnfW8Tu6M7+LJqrVV55M5OQUFAPMNrbmoWh1dlnWUXzva+
oB+kGdOP1BjnSTEhDeHC864xD7FA/52jFHwalUglzBavwseuIk6i4ufmxGrVVOj7/20A47Jjguna
KfWy7cKsPGZZ35Ji0ko6ZinRGPbJJBuTid8xEYxR869ohEif6WoYkf9JdBBLNLDl6onk1Nc+aH6c
rCQurvUPpwXlJGi1n5+ICZNtJtKoUqZCNmjRiz1AQqmfN49rPaiaVdD8dmJG8IwNNoxoGB0wZY5A
Cn2VqYavpfNFyatMxFGF4O89/p4ehr7FgjFsSeqOoVjWtzqvPzR2BOFsScs6va3gGMI6nODcwLwP
hJ9XypRF2fpeNclQPKOYqiCmEhNLek1MkOUpq2pW5yyBp3TdmyiJOZy6uA2yMzjIBYwxoM5X+41n
E9XzSvrmyT5YbkvRza5II1Hw1rDP70JZk+0nRp3K0jOBQRQr48jmtpxVIlGaECWLxoDzqnVsi+6k
QLLT8BDwaU8rai6pByzQnl26cEQiMgyhjrOiY7HX7dJ9ZyJfgjcxJBo/sldVL/zYveiYEY1e7Xeq
aSmAut1ByXW2k+E+qlYAZwawqoLFAcJZrl1mKqeymCglCNnSc/a/sbEK0tsE+FqSQTeR166jbT5N
MdgQYvQftBEfCRDB/zOD9qoitlZO4dsRbM2TtUCszcHsgvwPjGNBB1v6wEUDGRQJFbAf06Vr2egm
MNeQayxGBE6SEwcfIwUiL//Xw2Nl74b/Nzu+TV3s5iIrEV4RgHDcMvjQPBpEprwecw9IX1P+AwTn
kND6nayxqLdj7WIAPGYkBGH//uX8egiCewDaq5kZsI7hIpySQV2YpLmzHnpkqtFquSmJ1L2A58Rn
P/fkY5sUld1FEQgBbldkHMv5yrGuGznHo+arZcCoEgMNJRjUTN8PAGILO0b6S9LqKqfjlevn7l1h
M6nfAzhBus4Z2Q//z0xYfjYCtiEAYRPLbXzIuuJna0r6g9s0vVfbdm3yV1A4Bb1ZQ0K1dM6GipJt
WkyYsmsyWWo8JTba9X3J3517wOPwga32bYTc8iBrT1WGkl84f6bzxYfurt4K9sJc0fy86Lp0bLV3
itIimdJQDb7dHjmYxZGo+txY7R0Iz0a+tkq9nca9JRnqezX/UVQKNKVND4GUfDgx/b96eWUCSe2D
8RMg58oeWF62xheR9rUR7TR8SfwMHUVNa8x6ygb18zsSwSR+odcMV8L7+Mddc5v60itbHphcEcI6
f3ByigzP1a8osaifPH/TNtE6ogCO/5mVulCm3UkgYMv2JRS6KbrosgE+65aAAWOAnWQpKsSz36uT
oNVinTy6Ig08edRJFcxAjTsHLGlinHKeJsWMkQQJQCcsEaFEL3GoBKFJDr53iPbb68/d7RYRsj5i
3RydK+aBdEjRU/65sz4THNuiCi6H7vATTLbGiKN9kiZU1xmFK8AhYJCamBJbL9RkBk5yYciMEysU
6q02mWG9xw4PH8bso4pjmh5+jrgxrVX/hCrBzIxhRW+JM2YmLJaEensxZkyb2hZiRrrrTZPULj31
l1crKXF7sMs+q1u7cRkC6IRY0rfBVkBfcEhu46zCC2ogMf6EZvQvYbySdvN4moOEvwGxKJbuDerq
7mlgdAR8d5NW93LfxO19YngRIgdAE88qOTuWVcCR8eUvI8vSeC427agzNO646FjES9mwD6DQASOV
/8+cmPFoRhut2F4JwW8CGcYsWPS2JAiJwJUDVVwPLLnEOoO1G7tcs3nkPhdrFXcsDP7O0wv/PVmh
GlcVqsZuZ4zxowTwsBAXIux0Q/BPkEyOSThI297Sm9IrDE7Inl4bpIRoRL4nciGL2WQykYbynx3D
/yXV3Kc0OQaWoKbXiBb050xR+4PihXMreGNW5Oyi2SGKxGIZy7nvoFG64x7kEK58JWn5PbebeDJJ
/mhHReJ1//5PeZDm72GCPq/5WGSUFfSyuqD2tezi+WmBZUmuY4Ojo7jwGfB97yPWs4lKTeDQ05jS
fq1xZnALPOI4pQj3YC1fu/Q94myAvNCR99Zc20BRjIf0r5nzEU+IzLfTUp+5ozzKK+ytsSo+RKEz
g+aZsLtOHSYt5b+d4QMGFaQNao9pL15DkYuuANbbdKpxgmodlRlTpK9sRdvP/Z8uh7r5fju8x4tB
c7eK+L5RuuyxCDjPznrZMH08D+k5Y+FCqGUugyezn1DIpz7SoqHJzW3+Yoe92ccdnxFyoPWyN417
SnFKa/9566Y82uqKDT/caH9wTSSvXQ5/qfPhg5aDzxKY12AVqHgxLSEd1sWPKjRZe3icUZAfp5BK
dPdqmlJHQXoczQgApYFGqpLUN7lw5ksINp3Rb8VmLXo9TzY4rk/HZxR+wXdDOsBMEP3WW17Syu8s
9hnbxtbIbZouo0oFGG+EDkVQELj7y9tE8DWox/w3Wu1Bj340vH8e9JpeY/Uy9BYyd+Myv4Kxl9am
atsYl3/eHX5MYkqFpxkrKBIyHfOK0PR/Khdpg8PkgI7hV+8XTHQhRSpF14xZ1H1xS0PqE45HyJqJ
HjIHqGw9IVj7hkTQIUnxCByVaqEmp4l0wTESiD1m/52DggKUAmeIs+WuDKJlORIAXJi0baADhArY
iLEMviz5dQlum+9lNEPyW5NCKhjBDAV1KUAJE/8PEO2LuRZl0qdTryAiJePysz419C/JPe+zRv+Q
EJpQo8L39vN1ByqIcpo3Alrxa+HegXJxyQRTXpKjkD6jo2WyN+Q3irNFFUIlQFetwCh9WyI7YyoD
scheWwNlbLbE9dV3YTzkkC+nbuZ4kbTvTJ/QmtrRgixwgZs9OB9WesI1z7Bo1Dxi2o3eOH4lrDPE
FN8oyuywaIsSR9mTTvnCb27poNkTCSYKXNni1Ubjwe3SgC0qOtUnXQORukqNcXzs0+DkN74/RGPK
/sEAvu1qJHWLHvAKDcm4FeULNTJQ1GEJ1nA/dxvmsOSdEG3RhS18afDNSTt9dzHgEu3ESigSJbRm
J4eA1NgYdCrSkZVqjiKvNLBJnLCvMV0Cd3p78ZzFG0EkVdvGLmQOkMvrqEfmTWnicOYwGqYNxmsf
GEOeq38djZlzqAmSwxZtR3bMI4xsOwGXr65BNbl5FFowQYudWg3oEpZF+2JHG16WHvrnQLybNAz1
DyUVzMa7K5Ffj0YWYRLNC3L/s/j+I36vt+kWsxowzssVmvlp3qmiwECPeVc318aptuGRyOw11avf
aF2tUh1RTb4HHl+Qiup9OElF1f+KnTk/Vm8/uqslEEfpHvlUv8k6XCxqQ2iEZ8eSOWYjobUttI+K
Ssb9kzVpQYj7e4Zu2sc75hkQjO2C0S1fg+GhEBMPFBo9vQOc9Ks41+4BviexVRgxkdFyNKXXxkNG
MYVvJfM3CLks/RFyeerViSlIk8/q+yW11/gbMmvfAIX++jh9GLWlMAfP+cAb4Zq8wJbUjfk4vRRt
SpTxLWJ1OGworhsYyv1lj1imwqp49IyWeMI1XyzTuwP1+fMcOl+rpRusnes94JhOU/5sAFgo1dgr
sefcKgzz7tkbcb2jp9C8JBGFYSdE7ZU+xgRdQMOrXCpZWWwOipaeh0HdNzDgeD3X/fSKxJUA/p4e
iSfkwfl1PWf75PzY0myupRKC4VcQ96JWsAv92XE5VSGS2cviVoCnUvRtb77JHB59sRMe4qgQxI5V
A6FeJTQJyvd25hX0hKykC84ymU3mTwTcHO+Zj2NyQrjMLtZ28BOKl3FvQgALkCcnKplNmC2GHnbm
ciYXL32XIFehldAXLA5mCZ5gPIWD2WC4msYYT80ljtQXmFtVnuPsyEbcvk70OUD1BZBVWo7WMKPb
JFkQ2wW28K5QwqePbnwHpXqSIoS3PxrxMW4gjsfUvNlP1hecKZ2cWDloQtrFBdcb7exTEy/TPkZe
2sh4TtML/DHff9WgaIkLPI3Msx0BCknjxZJQ03sxO4vDbL72a6t4P5Cp5pGhA27hTkmYRG5n5n9z
TKzg6r+GJn6hyyvTjvf2XdC7LO2D4ZDW3O5UGfjZqaxXjZpAZTT2OnMm74iKWqnRA4p7GIo7gW+A
eLSeKI/v6NZuMlm1rjkxfBalA/Gjd202ySMC/w9KIrF38Ez3/y0fWH1ayJs6P4X7jI+ql8+ISt4A
ePg7kzemtI5Y5IsWi14zMyf1LyH2CbrzrM/vyBQmR1Ow5bFNZHwA86nzapvjFMVr1Y2Wxh5h70SA
QKQbGGxxU0BC3JbRr2Io6aX/OpHeHvnCZRQPiY7lBN0hdB8CqvjkgxciEBela7vqk3d/91pCL3Hf
tBvmoigiRH71cc4uZRPXNlaGh7pTeW8JOy5L3g7F4FYgyA2ZDRz0mhJ6IA5h2jgqBA/9N8OvXl8f
X9lbPDquOlKnvWXZ1+pR5gF9y+bD4v2c/FM2fJYTwTu2ce4d0weY5FmfKZxplriRUUzadKRUmuEw
cPoujoRe2NOLuW1jWNwm0ORfwzdSXqlaFR3YH7qHbIDskv5fZoHKcVa4JMIF0MA4Zg6rxM6q/qPC
T4PpCLjosie9emWQ0uZPV7IVDDd90tFfCIo+smy6jzHgpovqujtUVd6lUhKiZ7MnM9uHnf1dULLf
q1tlaAEvaqDgdRtmWbvnANc4WNZXRotLO4dq7K3eExO8RZxEsZ4o/I6CgC7pHGOLvs0RcTdMFvwe
zQRbnJjpu/JQpXqF6EjbbxPKECd0BFwM0+DI4kl7F2k4HrSsCq4yZJfqLhLI3niAIZWrf2Fhi3aN
ok+2GLXBEIA1BlIrLSEH1L36WdnKdEs0hiwNsK9+jbzduEC4It0h3s3zkZauCR4J0JQX9pKM7NDE
Ka6ZtU5YDuAfYUSsEVK6Lg+o1NdSF/cpnkuMehuOuqU/TQ8zdWtaVXgu3Po229+93XTycLJcGVE0
Rw/DslMLK2EK/tkn2SZcLiiiqwsx9ZPN84ihGnIlNMuN2EE1iEKn05u8Wcdoe7qj11/Zfu2lQEhk
yE4AwCt/63okvo/0KDqs+cJjWyA3HYn2xlheGKbBkkxJCyHEs0hDaTXfDrJkhuZFt+HPHfZIxhvk
VzVfsfZNa0YWi8HkDiAh8azDHcQOIMuzMTFL8XdIaiHJXMpLQms2gHQ0uDqlMD4WBf5Ob4FbckNX
Ugy/0+P39pRPXqSnNH5GuVWAG3zztqwX4p7BZoc1BPNo1JXEJfKI7KAhmCXm8XulhjxGmm200MRb
nRMTnpQ+NElGXTpENLArQ4VBnSfRa+QgkvQtyH7sUjdiRl4o5cbqpa3ibdq5e9E9w20D607GbxR4
F53XEUfg0PqlqGngsurC9HtVlYumKq965sYa5Em7tyJINF3v2SK0aQDe3QK/g3knCGCw4USHfX6Z
pVbwL11tPUsBQi3grNLnyKnxrbgmQQjozfiGHzF5BoqHNX4C0Onik8HSWMz9FXkDuejF/wTzjptA
mA5yxHPZLHWQMan1jWl5OGODrAXqqLeB6F3D9UckxddsnNUC8IarxiCsps/6T5FUwBiydKyTubfK
jtKfUxU/3xVOSrPS6USf8fN+bk53xzH1hQVC2/HQ4uS9cviwMKbAMKXtZ5Tj3AbfquUFQLw5tR6V
I6NPC4e5EDFy2H9KX5fcM1qf2kpF9+zyGN0SC2X9ohcPdkn25sQlsiwGoa9Yf/QdfiRhpDgtqLHW
CVyjmYfgGNLMpzMznZLjgI8wTiyzsMlCMmRuW6gvyi4sPE+L/PPIs2QEhpu8JVwMzhSGa+xcp/EJ
lQhczvIesrEzCIRhLtqRJSj78rfYPAZc9vdDNhjjZtTFBtwcxAienzPvAmj1PSp6yE2OlYDW63ah
xeHOsqAjFZpWQdJy27Jqms20CZ57S3aVQ6Bjl0ODKEi0JPfYEYMmDqPAcaExOqBmZMORWDZI2XBb
HC6a7oEyhb2mELIgDfpftJeu2ttF4p9FSmm4yJR8JqQSZWpe9xSrZvpjYHfIkegzBF0m0J5kXJ5E
P577xUD+ObLKBTHZJ0PETkq35NXYqrFlXk6LqyCfzuecF+EWUQuLWjhL3COMWGYX23A3q4tdbcP0
0eO4iIEXrloUqXMUC8ZJCUnqEr5NdXqPApsRWfFXW0g/uT7fWmEyJCZ88V63E989foYEpBaZIp6H
2YbsTe2B7ikWJRO/UFDRNum8OAcXBmPSZWsg5FZoTl3d7np2EaND7lRWVBgWbbqthQ3e0w9I7Vwg
2BXj9/OQJCrxWfjWDM0cRqR5Jwy7irmYz/FMw1r47LDRS22jTDp0VPoE/W5iHKeic7PMfF6VSHO/
VBCusxjQHdPWMzxzx0Dk/sJJNdO2EkqA4KC0aukHOd0ekzJg2skp5ujBQAx/fr4bg3RG+wiJMPSg
LWeAt5RTK5SjeGhwzTDpfKwrtAdh6W5V2nEO4+dW+Qo6kqDGGK6AdqjTiQg0a0yUIFKYQoTmWGlP
kwVCopDNpGvx3IQmX6DG891noPSWX9KxxNvOTW4N2sK3WwWuqaBu0DakCQbLPjl4bM2lz0aAWUKe
zxYDgy1aFfcTgScxZN5BOXW/Q9fasncJT5fJ5jQ6u2Gyd0SW/gf/hqCcatF+kB45od8fWBEC1u1j
9M6u9kAekfyX9xQemysmt9ToCFaajYzBhhdbweN7K0zBqCxkMhAxs9n8ogEU7zZcGPOHUA7ojMKQ
r83QJgM7lVMDHhBRXvYH8fGrQzxNAe1SokYq0ZPXqIcS8R0pHZQ9X9UeiFm2ihnlqXTKH9MJJCq5
ZrE6+jAig4myX4berMDp3HbGF2MYvh0tJxzZ/gPAmuB1UywtzHAVeN/CR0ku5lXGI+zMRrk2haL7
QCAZzCq2WvLkaYLp53Jkf2rdEMsxbOmG4Wa7MeHGUWPoqMCytjZ4f2R4BLI1iRdw/hhrZf0xEesC
Z3rmHP+CoGQcmlz9tE4jdOrivpwkeHFKneS6IMNYgHUdGtX+XXQaqEK0gPZeeGz+yABO3ObMP8hE
yb8fBwsnq82+DoflhW9oFF3QvhmyR88PeSwZ9O9HlNJgeP7+a3fciWu3RMq4Qw7zvAg5XbhcyFhB
mlR76lnXJTN41+NIGCfQ82Ygk1CmOIcDVKmRue1BicmLUOrXLfq03X/806vC3ae2J8LX2j3ZVpq+
mZd/IqNoJJZwU3fi5SafeUv20obWRgsk3BWGxVDf3EF/Pvvpia47CeNLCTXhspD4B1TRxloJDT+U
UBClGL3sF52rinFIYrxxcZg9JGnjj20hjOZ5C6l9IkEqYlBouJaGIjdqdHF6oLiD99Y8SkhAYXaB
lhpdpyt/7wSkHeAGZNTChbYE+4aOtu3V9nha6GXd5xepZDWdWqwLzYkfKwLxIxqsEkbiEcHXdNwm
CqWiBvXbYHab8bqVFckcXaapo3PRSvN23QngH1qgW08NlyEX1EgDqIqmj2uL3kcmLc1fycrAkOI6
Fuw6GH8rtO0iVXWZxc0OGW8VrBhtBifM5Td0mPLQMHV2viBYuMh8qx5z4uJOMZN4iHlEQaSmP8D9
LGwqp5YcTuYE1gtkXMAfsLYP099YOBenj6KnBpdXvpOUZPH4dg1JihhirPq9hDciwBmCIXVFzMgt
c9AH7jpN+dnoLOeUEZVoLKs5Z1Lf9HWLTyzGaROK+mIbAOfDmLsjuPBOHRR1mjj0EWbiVwuD+YWM
wCOcdam+UGODG+Dh9ZYIBlSC6AImF91vLWuGN1K5I94UBmAKFOGzf5N+JXzn72h1pYAyhjIWLr0C
RLotUuVFXU8yURI9187HkLw60jjdk8fo0vSnDF2Q0zYdB2hMp5IZm2ykkUqFb+3pPqwLc6jVGTDg
a0xmjjEyNsPt16zyxCBPE4QTsVhL6geU/KTDkRXAjH4mzCgcWePWOpvUblEBzlzjbVMbvAFWmGbx
uu1Vey9z8dNGMf6RUc8xHZb4XMXEW/ne0z187kwV2prapYpOKwL+j5bCpjhlLjiiyriwTOQjdGSq
4hO5SDf0NCviJZYRBPVGZsFceLtvjkZ2nVA2Y5dqgHSdKDZo6Mt0+phjpQ1F7nD7+0FQ9pd4LyRx
2AXvdXl3BjrkzELq15xG/idC5s5diK104lfhNK5r53OSdR3O1nnlFiGjsT3vYE1gq+PfhllmHkq3
epD6K13FmVcpbWSBEdO1YabzdFHBErPQOhpi2R/XpAenrkF4x9t5+hqJAXL3VMS7GendjrIWleQ6
UCMuF49xAzMFXMEr3n7h5nndcGeR4TSlirBIiLScuP/4rYnVkkX/DK80jZPbf+JAxna5DpZD+Z8m
04hWVFiVZcKLtaUVI7Aj4gGnUtUIx6mFd4dhnyDB4r75pVRnJQAmFLX3Y0sWoYMk1maflftPLU6O
G2PEn6H+DX9qhHJ7PPZqAv1Q3D2i69Mqa7YjYB48jImLiVAU9CKI+887HBM7tsgEaG9McNErlQO8
eHgJbRtOcp6GU1bf8HF+qmPyROi2KrIA+EoggHld3e2DiJ65yAkU8hMArl41AX731WP6t35BgBda
XhP4rPf2uVu1y7VInlzoNp8weNqkal1cD1bt2hgiycc/DwfvR5lhhyCZs/utlJQvBYredpS6N7Lz
aipTvY1YWQp6jxYp0L/UMWEhhcZ0LZNTbnjyRf2BPh8x5b8OQEMw6qxxCfxFZcZDnYhLvhDCWUmT
rsDJNop58gJm8zG0vxZZd61y3wHaZSc5OyqRwWZR8/2Sz8MgvlGHUruBGNXK+Lfq9ABSCNvS/wqZ
DFP8RC0jPy/nWx4+8zcvz3Smas0ECooWAksWP1xH5IZsD18yfMt1K4bX/hVC6xaegEnooqhWk2Xb
Z3c6feMa3VQ4m7IttCeVahOeFRdegiQcTLe+XrQJpxL9O9DpCBkpPWUkoFf0mWQTWcKtzxPdx+d5
LB9sSlI2UG0P63HWR4182RHGg+SgmIYMArfYGCn6IoJuVfjCVWEXYEjJ0wHSyavyIa2RrirAmgIU
qS3ZUXnD/9UXioWGzLtwriZ3cCtv8M06X+c6UFWg8tioONZDO5jw6MMDF8NeS5pXK/uPQ3ZZJYOF
iUzKUCLT6uyt/CPf3TksFZnGTt4pE/jeq15qyNBWlwBOexX2HAdjeW/2aF4EseJ2YEH/69txJJaX
6r2ZhvRPTbqISRGgCwiEE2ivW3Cygr/2cOwWJM0oi9G4mvqC0RcEBF3GkiDCyLhBf4WiG3ZWWaJn
mISOi3ToWash57w5KKVZbx8Ouwz1iZU/0hjDXAyz5SP1ga0RFEa1Euxl/FHZ6Yf4JXfyIThnP8Rr
w0+q8pfFeECJcjhg4AhGe9eTWD5AXydQ9O6ckvMKZFsazAsxWF+w/xatbqjra54af1Jn0UYXdwhG
JhLHpVOa6UNmZHxOZjYtmWKy0K3Ua4dNIBM2fgKn8/wBCyg4+kvuChjnn7HvgNveILgbJvKKNZlB
3Uw3G8JL+XC4LbhgZV/8YigHZUUAw0KG5B7SEfZKbGVebDP2lrCcOLbRiuWAcTa+UP2CukVMh/pW
Tp7jO3dr+exEF0LxmLrnoXcF4cdSg/YC768QBT6rzXjW+s/9YCZV6HH7gTN0yBq8sx+ndDYcTG5m
gHqzwKPlCcUDz1FgzRaq8jNdYWBHDQiTuUSKHprMrejHZMSDF/Y29vfPXu7c8BFSQpw0HI4nfRQ+
wPvqNphxKHOSPW49bF0zyWNhM7gpAn0LxC6tFaviJqERq6wLfN9So6QsemgAdc0ewGJQUH8OjAGI
qtKqTYOvwmTq8n6qBVRzoXWh6Hnu+5eJDh7AQK1feGum0BbljU7/CwJRWqDaGZkvpvQ41okwoQ9L
BhTjNbK+QZ4BsHzsImflrB42jA8729pvplRY9p+2tj332xG9WL+uNbcueO7gdD7Rc5tn+A9Juit5
sg4TP17Lhac+i3EYPuUi96+B1SpayfLYjNuwUclgMbFab3W7VOi6OXZog9NaiunEXRlOzt2z/hKn
qqBXx7BOFZ6557KeiAxX9ef00ZV/diG16EvBI5W6nxia15Yp9BFZeuvcFNwoH6qhi9uTBZG5OgQq
kSa/NwKcPf/3NkZ/fQnMW27tc7/8v7aPBIgOsfdbQ0MKpnGySFeNlo9Q8BoA03p15okOHopiV9pA
e2SJX5ap4TI6z7Voq2IHnbK1MAA7o7i3o7WqOI4n5ivYWXMY1rtdUdhkAPlTQcJS06JilorItIEA
PXqxGviS0+fBCTzBY/2X6J6XiMGFVWIlGj2ls0UR95BvBgOFJ8Vi0p9yV9+kyE3/0xWhmo35caLH
rWmTs1RRt5aRWpabSm6wyODocEQpD+ylshGSMd7qs6ex9MkOmt/ydbFcy2GAINYbYin8xb0tJRAs
xegKUSjnREfmF4Xw0ECHWKfsr0+z+e+m4WpAhkBBoPXqqgBtfwSPM/KCasDlkvk+zaSl++C7kPSI
5AIELYs9PQjAzfz4oGFczo8Sx4yR6YcppB5+k+FEfakZzZjEWQro/KgYYL9mYITG7ggUm4s1Xa4z
JPRYhfnnocTLRNDB0cC+360uC87FTynD6toDSYu32IPfgmx5mBhgN5bTdaN+24XZ7yjnxbEffxg2
Ih/lSe8t+rI09+Cofg6WCoeDQv2vAkUVc6nUUOKMVSa00jZNXhxQAoX6w6nXl1dj18tBOgDyVEqw
uIfyJk1CGZPzs/b5nDHzE8PQp8Pa5kzVV4ccAf6hMh9b+BdeQewEPq4GDbweaO606r42L31c6q4O
UNrHNDS4jMalszSjFU26smxBNWWKH1h8rtRgDqiEBOlmuS7KWzxdssJmjINo4AhFBtETNSeMe7Sv
7zXCKz/t39efoBNWkTLx8N3IXUOQ8uXv4LPmIJrVk/QKoW0Aufgx3TCsZFybnfqGiLm1JtSvb92c
bsQwHZPgkWI5mFnTASWTdkrpTEmonqMDJzv3ycYUH1PdJ7mA/gD0RsWSS74PqOFg8W1TsLJBU6gw
Ol+/HF1eubwj55VJpKZOD7oHHvIsAV0ttC5ivg+IVmo2L0UjXWttHihVX1FDLkgfDcT0qbXdNGl7
mNH49MUhYM1R2ok0+ajaFS5Mq+ksANHHXJf072pkqpX/S8+MiiLNMdmZBp6grikzMvv0iyErrYBZ
PwdXcPUn8fN2X4ri9AOsQJeiWW6Cca3sRIvVMmDF576Er4tnFp+FL/lo7PO6O+8TH78y+kCXBbqu
3olFB1yfNRP7fLpX2M32RZKLShOIz3eWe5EVYn4QUIezIZoVr0Okz+oPd3KnPBEiO2ELuHfm3Bex
4q1Apt7nabrHhF0SQUGRJZaIxUBJep/3TEN0+CgXMuDUJ5lneaZwS2eumGlx6kxKzxLO8L+cI0HX
Gh1pTYnmcfZNJ7kgYuxpWhhTRo8YJhI+F5RkdkzsjDyFVD9FJL75nqKmn3XyK64XPFpizp5fF+83
1RgdZ5RlZSIhrQX0V40hPikMpq7Y1XGhj9xIPTlDlqykUzfezaRBDcg9rCQIyqdiP4MolV3KAtfS
e0PbhFFLaB725xERnbyBfi6IFrTpQOP4kz2ca6zgUq7MIdOIl9QIBxnwVEwsxySy0gyaH2zbu7uN
rX4nTaBCACN3s6Z+OAWu4xErsSpjB1chFNrvjN5IVcXri7+xWktI1+k292Mhvb7UY3h0cc/KCv31
RUzLFCZmk9ggdy0+7C31A/4SRFm2sIBBqpejFlRGQ4V+8xks5U0FpsXqs4rFDyy0VV7GuVB4oSvO
iZvKmQCrQAaKFGXkYr9CgqV40YIFNrVUO1a0ZW5wQRdvoJy7tZBBOkfEsRXrdYKMF2Q9y0ChxOvg
hvIg0H+GUrCqq56D3jfuzDCk8mJangbCw4AWwzRD7JzGTRsiY6jpFsVnYOAZFlFsoLPcQ4Twbvdq
K0C6REvCJTWkcDIqTcfxeCmilsxbqGsTM8JbJ3qSKH6NT7iSHkokvzHlEkX10Ad5ZTLahQsDJXGq
0/23lHnKTjBbH+rB8MjYkoT26Wyv5IiAO2KsdKr7zWwhu1TjWYWWbRWhvD1yv0CE1RodOSOVwXIG
fkJbdVKED8jhydlWbrQQTR/+922z0QdK+sO6AE6sw3eM6ycAT5nnp4wzfjrJnpcOj30dF6UOJMPK
qZxCQUML0du6dIdLMyRCZfSqy0LGNUZfNeGMBzldBpXsoAlBFp7GJPbd/UCqT5ADNN66r+0+UGE0
D498KLligpI6McheTWJ4ftexj3g54Pv5mZ61aL2557XPl6kBsChOzuAvHkSvQybTGsbji/Q11HIZ
mTkOoFrSTU5xoQR5yt5AxvOTrg0Kmm+Ji7EPVbAZA4EIgrwe/wK5Z7x5OxYMUO66OA590S7v8R5X
jmzH4rbTnUKCJ9ECGyKMYTFDnDqwPeTNJwTslOOUfUDf+dVw7V3gGq1HBemovNT1robdYoCCME/+
CQwInTM/mLnuF12FwtDvOFAApwrfQHihiCdOggegUeE1AMSH/APTN2TfAvXxWNxVAF13LsiTok/A
28O3gsoDeeHeQgABWF8iE1Ov6JfCGt25CYFMFN6x5MdI8Twht14LA1D+7w7orgxmNnaOYeX3BM4m
vjr/B3t8+cYDuRULGyWkomZprfrYuUwe8wIfv2R6UOVyKVoqVH2FDIUlF5sVHxD7tu8n0MOrBfpB
sZYE2ePEK3kwuzKf9ph6pVd46job9NNz6AtJHdPT9vTz3vN5jUwBHKkodobJGd7vWCzPSnQte6PQ
QfG/C3S3v2++VQxXKzgyXxUHfTEi6GDLs9bfw3tx6fFG0DS3uG1TL5vpkDITcuHFINHvhPrvVaNs
WT9t4lYNeYiqERAfvPBIbAYDea2wfL/Wui5HkIYYXgkEBYfIsB/wDmgYa45V5VPASwa129ZnI8Aa
VGZQzmma3CsNAbJc4ZWe9fE0LoXmC0v982kD9OgeMVhw7Bn0ekpaizlwgIBQjdgWc7iiK+SBHzB9
+K8Qj4zFDFvC+DrPS8oTjoLoPBHEWM3shMp8uxCHFV6ZlENdWNl/cvfWJL1oDPiAAwHQ8mKspZtl
nX1h2igUKwIb0FeaoDSzfHGIYVGLSXuZibCamc50cqyzhkvbfyrd4jaza2MJ7pPUzG/oPNZG+/rP
AtsohbMKz6MGM8C8lkuKV1khPdTilcZ51zpVOItzwb+6hrx88X4nnjhAhyAQ84fD0LHgLKjbvLze
U5xW9hiEKlCL29eBZp7RXIADn/P31h8lGv4GsLRvE7hETZpUDZW3LLLF/Tw5RXIrjcKeGT0Am+ob
6dXPAkW+vW1WK9Ar3VH8ZY+zxKKffn9mca+KZNWfYY8wVs7lsRWkv9aHAQnbSO6Wco3G8lDfh26X
jJSf6fakWaQAh+pMNI/Yl4FigScfkYL++3ROlXUodQ1FeLTypVFrOU4ImrrY6wPzXLfgRqQzVDtP
TaPWvqL3ZDyMBWlW8/OO1uUiSl/+qDegSgZ+y2V0EAqoJ4XlcCUQx2J7XbFyw5NtykVEnQoAHEMN
NBNAUuQ7gQTIMW3Yw7+DlcFvJ4toOsHxxGH9raIjxM3ypt07e9ukU/wwgYggOuPc5x9/EWJe5RUy
eCT0foX1yMXBhabitNFdsPTV8T6z338pfn2kOT6PvVNfOpcPo57utz8ZHDajFIDHfCW0RAOMbuSF
nEu+ohGEWd5fPDcQjSf8dx1F10ohIpNpn5PxipJFiej5r9XOpx16V6253BrZzpVDgYdBEWOpTS8G
PS2J9UUu/9wWmSa0IXCKhKAtzNZkVwOAfGs+RNVsbyfursV94serZeJuGbmaEiDW8WdDgg/RYcpJ
X8JkPO9EUka7BPDxqNNkwzCWSMUEyi6S971FYgaIWft9tC7TnHCuaF3+ulNdTIESMRbL1f7MFB1O
K/WLGvwlJeKPL+IxPtWU4DtGp/ddeKhcpsPW/bj6xP1cOcSItjXILYh8qrvdHqF/tNuZA6GGkse3
fX7IYHPWfcUMnrJrDUYuVm+ZyK4j1m66Q/Ps89WQXgWFmO08pmi1FLIvGEOB6pdvhPs9yXu/g9tM
O92qibwlp9Glc8uKZOYX3WySsMzQjCQ6Fpv2DKKTiKPHQKGTzenDoaUNu1ne0vxoKeuabMGs+9RG
uTW/pEKNh5Cd09zsD0A8RXKleG3HkCBPxbwzej73Yr9Cp+aocBdZVilxDjalcKwNLwR+FTK2WbVq
0wKYw8mG7EBN4zl/L0xtMc8zieC++9yOUQm/g98crrJQwvq1DeVHPBG6IXG/JwZUDxGNMMgcBjBV
OUvvhaMXcBGMnTTzbIZN1v9vNXtHjMHJozR3ZoycK0muPhKat6OHTWccIK6zgqpYd9T4rcJzb9hY
1pnU5agoSLngU1wIkYBCg6t6npC/S+hLAIFwnctrPb9YnJLZyORrINlLFgJxX+OykiR56RWLtAvU
mCgqu/9m4KpNUyyNecMJPEj62QP26ArITWoY2pDCSpgwuaT5fsD0RHb6TS6B5oMjdHZY9zxifzRV
9u7U2+yJMY/NHR63zFXX/DHv14Kf7aUywO+yqcBgK4iPWqdOv8YvqWC0Krl1m26bHO8TfL1/WFAw
ZsKmvVJDu5ni3qEadcLLyYKWfSCAqQV5u2SltacGQIQfaQtt7tZJG15ylQ/I+rOfDND3dOImEvvl
utsIKCXrgbOVZpLxQgWseKEWs248RqoPQSvns38nyL3iLdGYfXEMcF7i8LXLlu/UYNjsQevXh1tA
qoJojBwW7szQUexeM91hsFAtETb2mvVT+ueY13oe+r9d/gslQ/wetaQnvQXakp5gDBSP7oIk/5ZD
Je3yTwIgTRQttp8G90/9+hjAf5bGD3UpeF8U3SNQvwVZDnRk8aiv0P/GMmFjceErh3zhCBTkn2rt
eGJHLyqq1EAgH1PuJUMa33cV4RwTrpd2E7/tUWCuX+lzOTrruMBe1boW77fz9BC1px6AHZn/E8+C
dk0SxnxtfD5eVS7XKsKFrBKij+J1TZAAdAnOH5WC9lpc0py4drJgW2nQpHX1HGdAEa1a+S3RcMzk
gXF4CCOUsEk/Yu6L+Tg8wvoUdvR6nqg//TwZ4r/TQKFJs3Rf5+OYb8DppA/OLIHrWvGm/hFClK8U
0vdpwLilXUvfAdb7Z43OfuzijtmuAsJ0fgJPcmC1Z5c6uBkKj4LoHXcToRcxSNs7xBIhTe2dDjlw
ssiQHjEeuUMD456I7U2viQOeP1q6IRB7fOiKgrPxQRFSHxznrQTqTJ4A+luWzLqK0gx6xzBL0UmZ
rSFitzYB0VUoj7/TnsV1ffUTaoe/j2G5Vj4f8sRMsGYlbXt5CTk7Jqm09U+IdKoOWqKbzn4x/l3e
nuUYkv/gP7vGmA0Ysb04WMUQLsI1adRLSrF0x8EGQlzcqL50675LwS3rGpCajoStjs0/fvFbxEfw
lpilE/NwbkFFEptBTnL0ly4hnXSxKTCOddunN1TpD6BV2k6SdIMqzyHqVNLa17s/81k2zB/hfsE2
XX9niE8g/tPrKSFNlkuNAuNlQFEmPLu+/f31vOB9081c73Hc1kY3HNIQQvRAqqk7BAtRSf9C2a5a
O1B+64ZEkhQNOHRv7sDIuhoRv7yBLx8fuOnaCpaZoS4Mq9juj4i1S4/SY+HwFLTAQyE1MrxoC2rx
NV4QLvtXIU6QY9DlS18LuxuxU0pErC7u05h+DYSN3VRQwlc8aq+HEIUjHn+PevCjBlJHJ6DlmkC6
k0OKrpllHBr7wrDAi0qCB0414+/zSiM1LOrX+0dQCA71Q3asvCW61MtzNqONXzvrPAL6nUWb7wCa
pvbwY4Ne6106mNSZh0EvEQd0SFoSaxVqRFWPKOk0yLQ4EbTtkBUrZcFJrWPqvh9ZjyDFPk8g7/EG
PBQG/87XoAb2tMXVgSAFb46HYF/7Wr9/HLQtB7aFxnOjwXLJRYoxLqGFd9F+AupXadoWLfjYBJNn
uom47AihSbDln34ewj+JXVYQGicnN/+OyMx84fXNI/2a1Bk362R++6Q6MjKG7zCZ1GA+lYWGNPpF
XuL60YwidR9P2g0R622x347C5Q7157NQ0FdcOaLxE2cjVG4IKl39BR9tIHnCwjCNR0neB2pviQZG
qy2lt8PedTtW3ms6P32ELb66pAQkfh9JYZkidsAhfqlkId8VhTvk7HAaFzZkFPHqzrRpL2kLSgTE
RQu3HcbVgXbt29rWdz2yLECE1J4PklIKN7IYfOLaaOH/LlUdwU5cdJHg1LZ6ScqxF5A1KRv8JERC
6YaCGJ4vqzZBE9ujXYzUBMLZHAZ/H0BAXggo6ISRJZBGD8rVpNnLxXBzDY/g/rP2JcstE0Cx+pwG
IFTvhCdiJJzcQIyF2ogiHxoU4wu0KxAyMzMaaOxkvtgnPjhOsWjgw3ULv+oWA+nXbP5oZDfFwT8U
H25g/VrMMW80KwiFiIWxytqrbHO/kE7ahaYzZd/9G9WpCmH1rPfHVbkOcd7HR3SkjX2LSwSd4ki1
Oq4DMU3+4FWf4fzr3zo/uD8/ZeVhvdzXo3IbeMp7ZNS1Q/jtg53FmLfxtuDcKua9Xh+QBxPdWYl2
orH0dTMkoK4+34GddRRBGStuKX4uLZZIELX5f1pGDEDupuZQpXpjHlfTuzVVaZAEX5yMDoErRURf
IF5X7BaLDi63UL13WYTD1258c866kqYqCX6BWWdrppgtAY5hJv6FIvi+K87VXFelZ9tQHHSBu2Jr
EXBQ9wTSWW7/W1fiiukjKSFM3JF4gpHzB8tsaLaAfei43AwkRujQPE/H0l8PGKu5b517Eh+KVQeA
5KDAx47e8FmROg8Xj8Z09F2bu+ZcpNnumJi6vyJyz/QDtQh/g8EVci/5I1nBGzKLWa+RUP9brs9d
nf70iX5CDzQoo626JhtaVnE6VZdNE/yhD/4zWxgERvIJgnNP9Xvt5JtSksZ/vDxOQuL3VE90pTCf
QnQzLjY3v0yDzVQl9Nu/RQgUYncuO91jXIHixQJJqKJKS4Pqr78BpqlXcw+w8eZXzOk0cigRKzrI
K5DjBuKwgO4rEXZJ1wPTgpZLH55aSPC4k0pt/errLHjTamc9rwp1WzgtSVxawmzdStfCxNXyugRr
+4m0NlsVTHTpQ1ijBsJtmO482ne4FMKidjYxhnquxpMYVrgE/XeAaHan9zD6YQKJuNiFM6ahZzTJ
Y7CpCuezuTfHuToZBiU8TEumeINcr+CYr1uUfUA656OM4LOTkLgdpStRmC83/HsBUu60Qn0EXucW
c2Smxh2Hm3eMFvb62PX5LpcJY9+lqjZ91YiXRc41Ew1Dm6bZCQU/Y56Bcap3GjvRoSPSmrNVTUfY
et65E57MTuLISzcxPS880X6+/lLXK1Rq1B7CBUiqwnNdH56mUDcrCCsMZ2t1vlWEJbumI28aA6Ph
/qzQPFYRpX8Q/be7tN4UD2gYEjvEEsSdvpMzMHE+uy9UBSCS/UUvf8RbDPGO9LQp6tzg0/GpEDJv
sxm1o04dltoiCAgY5S4DLkm+ze8ofGFJjcMzlBDTgIvVYQDic7FpR20aIdH/j+nLaewyASspUUoG
QjKOYsXEvit2WVFujvvKazcG19K/htvaeWAouBsd+kkS3YX6010T0JnM4ETtJrZcr1tKVqP32kJD
jylPTC345xMo+YZ1aN3W52NRwUIDJMXpxc0AM+I4goWX6EIUQ6cmWLjPjKXktcnJkETU8QJ3Z4/M
eSqtO2r9XFSQN41TUCfrcdJp6oZyuAa+ItqOHB90Pjf+T3gYIXEdiLxP6XwSEjA1K98CKOKLcw2z
aGfvVCGLltzMdmI7yLv8tEZw+YBoJlKtNLxpl0mvZQs437UERyCPd3tdAUKARGD4baLjUpLMJo4M
kxs9KaFGHn4/WMuZ821vHiRGrfcf+d8Sm6GmKIgypdr7ZOafGFMjzPMr5uTMO8elWim8FqAOdVHu
FRuQNtcOkpmKSJApKux+wu+OnT6qw7qEAqJ6uciIrehmljIaCpy9QGYztGTmZ36K450k8FqzceiM
U6IxJf5/l6wjSoXT1Y4SKUhR+2XeNI4yCdxcM8ho8ie28nByhel5iAnOkA6qNoR0bEBzBpNndyM6
ywsQIIyghn/0xl/L1Q4liRuWE2H0pMsvTMBakzw/Nnzoc8V/0j/LLNinj6NTF0j04oKS8woyPVuc
umhOzycCpYZt+Dx8/+kxBVRQ98BwTKUxOoepofSIfjixuVKkRGTdjwhW7WCrVNNlJ4sjrOoPSmeB
R7DvPWFLZ8CZSJEurGEzx3i3Mb2Q/zx5lPre555x3yTkf5Dz/9Ai7fHBdgXITOvMoLmnha3EAutK
/eumUxOA2gnLWxIn0N+xAzau6VdPFTBAU0LUGRj3WWjdjWWFAZMZ+SuDaXySXcrAfL4TIsGqS4iT
P6LjfE7M9dLlK2cRbt8MSKldxfUVaj/8QvwG1YuKS0XW2Lbcj3HeTrdKf3cgViP6/yV4yynDx8Sl
tZoW44Tkb0yyY+ltcu/DoCQtgqs2dZKj5qdJ3vtyB6dLou7aw/XP0/ZFuXfht4FUk8952dWBlcbf
QaslV9HBfdiHx0jTkh+IVNpw8DTQarMtxypZbGEv3x4dCipF46VgGXsb4kuHRDa5umqfUxNsrQAt
00ZdhdDrA1H+VAmbuBxIgXRZDoSon7XQbtMm//19lTg3LmDOaVR1YqU7rRCcwPdyZg6dwbFca3LY
6J5grH2eirpfyfKg5ceuUgQItLKU9Ue+BbSvdvEy7u8jFtNdkSa/TDvFj93mZ+xmS0C3Pu58OUG2
y9VtpVfmx4vK+iaObuh9cdOWXSE7vx+q2I+uACxvMYyCgxExaVnFeug9OUxUdxvmlZQFD8aVlvY6
mtj92DS+qIarmhl2eUnoroTND+QILj6W7obzif6k816AIbMrzDwwml7bua729/UfV/napymWcfau
E9+PuEpRaiw87mjXP0Yf88+HR7Jn4FkWpvQLJaSGRzoCIYzVDb0w0k1JBPNAtNyuG04Z8Ty2dhai
KhiqjAQOyAd894ajmErAX9pyjIvUg0n+/Yg498KJHfZkGXi6Vf0yPBTnHZqBAiNXx5oyXwQA09BB
8jJYxVzy+wrbA8MvDCGT0YV0onA2zhKbwaroiqi7pKe66TkqbB2KAaEU+o8gfN//2Lb0cM4K5E6j
4e+5vj7a2FPXZTZe0i//DSJIU/fFp4y7vPiIU8sAsJuH05PRiu8f4U8h1JGbj1lA+62AHTj79lGz
ljDi9EmecCyRA80gy+LZdulT7kBuPaRtbo+2Y8iPfy8yBoI0Nhl/TRlKkOwsuM+G4qJfpUnysSeK
DbqDOFoguAcwQrq0foYpeXMW96RcaQbv+8MDz51P0VLMtMr0OCMPUg25DOr/GMsim1ro7rvpF/+N
kgGdrHNOcnr097+XHuZWs+3TQFe4dgTmwtbjzPmQ9BdwzJLGoGykmU+MNm+mXzIwRXjbmSNp356A
jJ6e5MxA4JaeMiS7xhyC/pLGMgk5wEQsS+M3HDHBPL7g0I6wN9xF0d2wbgS2XPir5wpp6WE9xUEM
s1ZwYuQeitRFCFgNqdgd6cTRWV/KdIOiptHBch44NcbXj0imWQza2XYCgWLNY8fBHcyUJmrGHOdA
F75J2SC8+6xOc3/PqpjpS0yp8BoL8zSo0RWrcFMvF83qT9pc8L+rXoOQLu2NKOVGJci5N5reIxvL
nQzW+VXKlJiFnC9uGANawTFWRDLC+jPYgCWX5d+fJSrzkaUomv1tcaNsiH78Sq3bN4i+XBYQKCyA
4ZSHj0RzZBMMAbVNp5Vv0IGs2k86VM9BQzKVEKF+j4cpsqCdEDqpLThh1v5Vbbvs83sCiGDZDkjd
vfeE322XY9xKDgDqBN/gG+9rhfVpwt1OvF3KehEUYaz2SmXnjrOooml5fnhkZzpvgSQPuheDvvEV
iSxq3fcNFsWe74vrsQenhFKTsD8rb8Ilqw3I8PJz+rE3ibfq6kJI4bsf2lGEz12v7eBC0XyGVynP
Hyif0SrEDh2CZd4VAmaP0C4O5aOWUdDMfFWGGR4s7qFJ5WlPVwe4p8OpDGAntDLSePoaVLXWV91j
+VglYJ/QTahhvzphqnuQ5cCAQfxiA8w0F2guVfW+jtNv76Xf3peF9xvIgMEuRHKoCp0rvlKFy5UU
vENmXYt5I3Ml8NxPEIBH5F+GdPtqiDmFGSLb2Bs4yQZjdsMt+nphs97eouyUpwxjVpfIKYWl1SvD
DTQe3ZWOMwqOdtnCxQw+LcHc42S64QtF71/PFY/nj3bBK0QLe9FDvNrfQ9xMwt780bEElrSH2q56
8DrYN9zUOntFdHeHzEVvpoBRQ5a80DWWqZ8f3lZm/kXrtNdQFW9yVt9/pepb8KEj6ExVYqD3NXpy
tPDlIcu9Qfjc0GalmGWWm5xlmjwAszJ7EEdOvVQxeCCDE/ya1uV3l8VR4J/P1X7/zJmQtXVRJtHb
Z8Yaff9ExC1aQen35XYu3OxzFPp2nN1PppCf4HPOu1d1kxj8IKe6Umjq4EeCR3/Xe6fJHTpsm0Cc
J5r5/391ohW4ecrUk7SH8S6bA2cVmK0dnQZcWJkSCRlXY+Tz6p7FlKJfcLCZz3Lqr6g+KKmKhCkJ
ndCEG12vVCvDozLPiQHScWn1nWVmGy6zFD/W6G9eADL3aXvgFOhkccFOcI4vsfVXHSY3MnXJtrto
2JpQSocR55zujorhp2UWuRxy+M5B+V61VxPptxASSLKjbRHC5ppQXkHURfZNiRqDDCSuJwTEgVxe
6zyLp6oEG4Yxq+3i0Odfhf/BSR4igpTErPJyXTFT6MDT3ciBllsk/ShLzSZ4pdHFog0Uu3542bof
uzPy3oO9g/IjTdRQjyGhqWg0PWD+9PxThZq2u10xenUh+pFF2tRwqr+me1rcSGO92RxPWb9U0UpZ
JNav/H3xF/x+oMrh3lYdAGwbMgv6oQn+EIx2RIO6cb2rdIw4Rl5X+4rM5X8raNTnAafczBWnV5Th
YE23H+ei4Rl2RUdgUYUkZ66LSsz84jMwwemUNtIh+yMt9eaz3FQkcWjXyVx4zjTjgPTD9ZIrMvKm
/IgLnQRmJiKY/Y7gxnBg9dvg7lZKV9Dw8GQ0cd199Bh98nIh7wXIBV9LTrKCoECDD+T4+//Zp0Hm
Y2MTY6Nfq6iXayXDK7arOZqsuDo3s8BFk37hVJ9I0gUTz1oBs6JaC4cyIWcRVv5f6mDXEylJBSvG
iUVKA7xic35c2OY42lgMyBhIUExsxrErGar1CYTJ1z8/Lzk1g+uv8AZBW0GPGLxfTISXInvGlriz
M2PVxtAD1SwqVpzQ5nqsduEzc1k3ZVIwarxhivNrGrUhT+fVxMHnanftRQ3BG4tzDJeq65qKmZLF
w5QjcImSY8PfyOhGcxD5mh3QX1P7RDjtHX8Nc9ughZYB9ziAd9TrukXAmaxoNksEZO7wIQthVZhH
o+rBD10Our08wm+BbYreDS/YsHMvg8qoL05nzvu/Vm/L1zNaluXTv+VS1FJZgk1AXIf4nypPzCKQ
iXNj3+xbgHrEYekF7X5E98XFJzyVnlaO10awGfWVmVTmdqVRK/URFhF1O98LIifEBdHIy1foJJIT
8tIac/Ps0HDnIwrORjZaUu02oYy+5UQ22FE6EwQT2QnncL/1giffafIKOuVaDa42xMe7PDPvYvY0
Y3bJzt8P3vpE+YcRl8Bhvf9ArPCLpmPC35mn7JUlKOUGrJV/g70h/NMOgE5j+JLdW8200Cu+aGFr
3Mtkma1gZJIRIA9r+E7SEptRhndjLoTE1gRy4Efej2d4TxbmM7yi5FI57OjlrmOvwYoOXunvI2QH
pEygnPMFcVdnmDU+NtEQWCQaranPPcsgDDUaVy0WBIutG4njOe3YUFSocGDPnLlG9sXQ7ls95ByX
BdlHnn7Lb22SObAegwHV7V83e6IE4Ls52oJBDa9NLxvrF9Bh9bpgFPe6Xiuj45irrPPNNTirh5/I
mQu3GxapqSIv77Tztg9PQmTK1MKfkuUqjCbyy1MU3oVqnkSwQoHzk9C11fHbLjQvBLraYMYq9Ooh
zL1/rWLuz0856/swENRKwtenEfEunj+rWcgvg/m94sb4N4bfhGowRj5sSvJSGUOrHIf/YpS1vXoN
UneyKrz7hUr/4TO1YrB427MxSre45hsFOkS+hldVUDbC120XB5/pra3vNojj42vOmgSWyAV6RuAX
gnym3pQgnaT542mAfN0w8kIo3IFiCbBTbK6EgACfmj5T/wPn7RfcSxm8mqmXhSSwdOV4lCp/LxUs
GrFYKMotWbaFBYFkd86ajVA3bPfF4cfqqrmaJNRI2VsXUx6QDimc7mCGmSR61vdqGYLXYqP0QNif
m+93Xoomk0sRoXvef6D/JTxxSrUSKSFG4Z+smepWqKtvjrkt/hlRKH42OMiEHmibFeGkshhfkrfC
ILipt6rOijeapzhNdceI8YMX1g2xTpawwTpBIvKI0X31/4QhTTAanFBZlYCr3UNzP+jN+RDe5Jut
phnsgUwXULHRRJx7WS9Mm1OAy5Ssn6KWjB1ySIy3DxsFfRFIA2T1bgTB1/g/kiRNIkv1EZSLkhj6
wJ1WuDQnhE920uFDI350UiwC37Mqe4f8xboxILMf9RxxYnvf43eLVdIh7DYNGRPKJ6U7dfOInQW7
/iRWVO1CfHKXJWRlNd/DR/CIfaM3cQVOwvY8SzxtfPTWzXnQDm+UvvSvPCCpthgl890F4jZtIHlI
dJtWdKc9CMrAUAX6724iHD2pATjCLSszTYxtIcq2IVmyJvtfuaq7k8IBMxiKrLM9fAmDl03wWbTr
y3jELT/6/5KPdzRD8r5PdANkjJAMYh/4nZjTrL+Nr4FCLWE8i9faByCgHLG6tetIbIGRCjCpHH+2
kFxCevFhssl31j5nZQ0nTXk1Gco6XK9Ss+xWubg8FXjOj1zgm9W+kKf/g6yQ0S7aSTc623QC/6Zm
2uLBgDp0UZnaNJjO+U386VV7lpWO7f1WySAxLpmZ4sMhe9YBrFntjpCkVlTa4G+RDJEnPuuDpdU3
IEHPWRc7hrE0U/9AZp/0eJ8w/yae2JgfUcYrA8UCGdd9lMhkGOUUkYdMWADtvVYUJ4q+fNqunQDD
kiD96JBMzPX4Cct3VdvBnso3wP9KNdz4RIb980ZceInjhs/aj40C0aMquKfXl55zqubPOKl+KlM3
So+EcqavzEDtkDY2Oz15glaCrJIFamkseOo7m7A8/j8Ac7csxIbpUWX/qNaNQtagnN3KuOL/llQA
Ot4gYmFdZTuQExvmpzt29kZMaidij5YGdNH+WKs3aVqgVI70yj0uqdGS9QtzDyQuvAq3fsQtzNUW
MGizv457U6SPavq3eNJHkr3glLCoDr1PmFE5z7jbHshqpIdreFiqkuxzioQaHc11FaNXwUMbzit0
/6LMIS17pMzPwIptaKBu1KBc9YDD9bTeNK1ufzR3N/+MKnLDEQ5if5bOQFxDrp9Rg0OpbdNvupI3
3UqSfsdY6V2yj3YHO1vpB3Pl1rC+yVWLlRG0h3cHXMRHMgQj7exFdEQ/UZRaJi/3zzQTWoDcIcJ9
fKyQU3JBO+Fo7He4OUFuq4mffWt+dN1YffmW6r80+Z9xf22ORTzSrNUx5vrxa3ixvUbKX3T4YiBz
Tjv0HKuc5m5JP5xQeyVnxjpOqXkcJ9L6V2S3f8I+NDAWmTgwTplVgDh0j+bfGmRgzAtUgVovl5/W
IBg47HGKVVsFFlmaO/J99O6aLUuG83Wr8s3jhDEXsVAEL9lo0rvR1G14Uhxr2f9AIYjJpc4fuxTX
T50y93Zz24kGhCMTBoYWEXqy/pvblJIdXD4/JR3MBHgmeqzDI6jkvr+wWGnVuLmub0otTsFcmw1u
XkplJmu23TiMZiTZopKfAPSOVV0DN+5WZeILsX/2aZf8E14jbiDQNTB4PnMCrM+GSP3axsnD7EgC
+nlyKU2HoTPMyxRCwYrachcGAXWHDvcvX90S5h8oxhcK+l++Tk/aNZu9oG5qFqWNFEvnRweBceTu
7HxpnltPjC5nUGu1nC/QGJQEWXJzMBfEgfJ4h3SKylAPCN2nAkLzltBZ0v0xtOmb0TRIJY8lEUVg
GRxbNCdmJlrfnofs+rSHMw5BlmeQ7M61E1ybDr8TvVXKFDkI/2TBbQEKALKglMwas33f0VuvG31r
Cn86y6K2jM5j62n+Rne+SiV3yIAR1Lfb0Wqgsp9DwwYufjLuGeuNOPNux4fxYniwrLvotvfbnwkX
+as7LlujoUk2N45s+AKkar+XffodAdNc7Ynw6Tnr1RoQX/FCiZSi+7xVhqsvBbvF3e9k1AvG4pdc
fwKy5yii40NJvJNFUBLqnCUb3znaDeTPlsh2X6+7vmHNOAIKH019qviNkPng6kOZXWNBsMvCkLBg
KXrqoRT6R83rVNMO64j5ItXAEH01nsnye7k8r/UR0BvgS08/zJYVKoUIp5/uGj8XGTflogW9G6Jm
a7TWgQaRTizG9qJJ4GDA1d9CVA6YJNp6HQBOm00irt4FdCvZICcbr2dXbaWigl6Qxa8osUA4Z5ta
QrQEwsjsfu4syftFDeuCKIOnmwuMmEdMd0p9Z6PwVY421X0lD4C4UOY1i5WtRwJ40ZluxB0qw2FE
sfL8qPgteGxocwRBzXpVRaEWNbnlbif1/ly45M8SqRSECQ9nlXESwkRZNHnekIZMDUS0CchAM3P5
uXQ7/FkrsRVLf7XKOdFl/5SdqWchufnhNQ22HGOPtSzmyxWSZ2udHveeW//AAOMLJZGo/9ZBDr2C
8Xs5JUJ2xB2ALyOZzd/Zd2/WfEd7nTb0tG2AalSvu9GMLjxlYJ1tY2qFrAsmVgbffk9QKnpwKt5+
Mx/VrZfseP4ryZfOOAW53F9QG7y6u8QdMi6gGZIQXIogcnkt2uTSJOhJu4vGypXYlCruFLauyEa1
hJb3KI5uc1vpTU4wYkPk5YW9lqJFEvg050kSj9CB3q+RxjY81YIvzhEKC8pBLqAm8+SNYHseVe18
VLavRuiVf60upaSHUAQLGCtrYtLjPOrWl3+WSK7q1pCtDFqkn/wejo48rOEkr1Urn8K57Ng438Bg
UMO/xn8svj5vAG7bjy+dR5p5yfLyClpJ32FASono7ncp4/soZ7d51Ojf4LY7APB/ZUL7mQ/t1a2R
huAerwxZ+zOAiJcqrNmRZz2D2WslPcQ3JWnanGVrMUY5wY9kf4kspRehiEx6Chv/0amyX0W6AVb+
167ntIf3NOK191vE7PH5fMZbnw9Jkv9i4LpE90CQ2o6kqwHIizMJMbfAgD/M6HQy7BrmN2rBoKeW
j7A8d4W+FruDWhh8cR7Kqu/WBqPehM5RiFdzRplDiffrJqgtRqrhkaRJsK2G3/eI0sQqVyyG62bB
ixypUtJSnEY90Fe9wWrpLFEUxl6EiRqXCgu0Knn9It/KLycNWTn6+IKQazUTSSlJ+q9vrPD0eJDh
P5uvrJ2eTdkEH9C6ZZ3kOU0vwZtdvBk3/7wiFWd4WcHzrxvgLY5PtDP2caTeYDTS3mnOKde3j1sI
6HgSTlrL5s6i2baMa8awKAy9Q/1IW0YzKOMWEepJ2Tk9XGXU1uurn2Q18oZ0ENdAxjJAq67jdpq2
Vu2z5d6dnfGJ9L7xYo7n1dIyRzKQR1pRNZJombjhk6CMBBjIs2tTursuwGadoctvQuI5J0KVqW3E
2dy9eppcJVKSgmli1TQExcuCO/joONOEtp5gVKezgTYcSzGaG02Cv9j9fxx1F7nWcaf7xvj/Kk+1
Ql+TLMf0CqlAK77M6v4U/IWV+1Hn4aWw03ZfCQxRmGhWdNDKpm1dQgwRiGfDIWCdGbalAh0Uju3A
yjXXI4S2ODkwdKxV2kaCd01u4ZRPcj/ZEyGXYWTUNJgvuRAL8RZF0By2WupnqgY1PLIGcy1Ws/Z8
nczEuSztwQmOrte7cJSzkj8ozj+ESl9ZE9OHmCe27JtWf3fIby8OuKautn3nlcisPPKhxnKUnkIM
XACgd/bHqSVYpzw+9kHJ3eNXRHE14dQJ0lc8h8yraPZD+Cc6mU7YKBdvhQUgLhN5HwMspoIFQWlT
bH2GTri+I1PtDSpmWlOEoqsARdhsd1F43eY4twuozc74q3/JnbZkq5jPf2yk53O83hG+rCG7txp1
xzQ8/RmcOA6xdDnZy6GTciMInpX6CWRERISCjs7b1YCuOlHQvfGWz7agZEZd/phrRMwtDoUfOeLY
K70h9bHo46VIgo4vBmH9ab4TyVVK7zJCEAFz6KLEeHGOTgmi9WUlMEmtesnay+WWaQSDN8BMHatC
l83pIz6qS0+xUADh8AIdSZU9DPkwLF1Fq83GEpPZPBS+LmIeh7E33YqWio1Gmx8vVat5+lkjjupk
/qEpfbF8SMVFBozzW2yuTz4gRHVhq9it/KJS5PMj/j0lm5UQ2UCuTSBbiFzlTnRusyij69gGrLcK
hBC+dWsnEcDZRLZm3hZdYTHsv+oq77UCB1ZpkZLlk7JLyRwuFDv18MSdoAygV03wV6wHyH/FzYTu
CScUH9iwHH+wIJssS5Eg6QVXiQmBoXc5CHS6SMsAB2k4SEetbEveETjiqUTYmA9WIJa93vXoiipf
6JpAKsBqBI+imAYd94uIGoc93T5q/YfYLWyI8hV0CnFgcQJisRNH0kqwUPS+TZy/tJhCVbmwiepb
zwzixDFclZvmxrA4vX8/NX1X8QaEYldG+5v9h0uKwis8rfRM4c9b5BFG/w5oCjh1nKjyaSDWd/bm
5R9I/A2bJMHDJdExtzzLI8g9pzdMQVQ776I0SaZrHe18OXZVIwTCtOC2Vfxe//ielbz/0lEVviBz
4yh0FjY9iuVYkQQIpRMtF/bcpHWHlM3N4LWQy40Uf60zKqcZpRejQ7merN1bzytbfmBKaCzFYBUY
2NzsckbsUb7U4wSKfUfEulCsvns1UE6RhsYXkLoOCDxzIwdq3KezbR18AgJcT5or+dLlFrs2Pr7y
8T1JcTylGpcmW2T7LL3b+mV0PLJcZRDPHzzpzku3QeRqgsjkoc8Gp8O3h9SmR1XFpwppNgGz0NRW
YigMs1fMJ+aTbkGNOavXPfPTix6NPVPEoevvq8xNvITI4iUIQSURUbx65vriQSiP9TKOgfV7lhLs
MP1lKC3/ESxY7G6g6DnjxhrAmtt1px1uJwStehRF+0I+AV0r2yqUoV7gVbGLB6QT9kaWs6kCteqX
N+aG3FgtAQj1JeycHrEeUVxXLHOGZJjADGoEYeUH0QFZowVt9nsvclfnY2sX+rKlYZ2T923pgixS
PlL3ECLXXfM847v6lnsdViNbcYpQTf+WbGZk2tKMDJZefuqXdq9dQJgmyh3PQwMzwVhhpd2tw3IE
cXHmKYhQBez2tkPv/cIEuwrWGp9bBGDK7CsrGqItRSN7rMlRY/e9TWMH0layvbvwd9YrQgdMidlJ
KERiQhRPuYkEZq5/McGq7eyeguGJ+eA1TK5qP0Xf4WQjktijUF61RMbLhMb/s2LcRfZFIhq1aSBh
7fCMxfgcUHf0UTr1ZeTD6WPwwOKGH7fVXfEUFDpjybt07gGDi6AyxxEdueQnSjBrfEw4ZJdOBT7E
woAqWwiqoPCSTJld27a81lSoEeq5NmKyeU5EdhLd1OndpuNYCglxtjr20vGj8nORfCW7xDZIsdrk
X8a69ZmuwZkWc0ZXz+x9WpLvPNAo4ZZipwcKmaDPok+CYeEemnkLiWuPvLjWvdHOlrBiFp4b7A7A
gqdn7KFTWdKepkoP4oiZf8N/3ovvPgkvE0AWleM757zIn1/40BcaC3tb6zTZy6v69C00+VO699sl
n4FvsyDKfOsOkfhdEmAkW5WG6EudYl/9mdSZEAmm/OCRHjj9LsTDH052t1WpsQzhMYlLiR6rlVVN
KxuOX3DHX0zUAiqEMMDUR1Zh2aDMK/aQipUvuGnzA7EwnnPU5S2cg+hsrroLhZlf9d1fsF/T7y/k
JQYPG3hcs/xqoLYnc8rHqxFlv4cnpGf7Mgzm+rGV40XOobDiROPKE/tkaLhmSCBCMb0G4Ag2wSLB
gsIPpboMaLKcThmbZ5T1+Cpfx5+TnzcGgiIaYWqy3PS7PMgy8GQqGOC2lrlffqDhSIehxue6Xeun
yE9DHJe8se7Sdce0lIGNjxNWjdrGyqTPD7Epe/iSvDxANgCPi3Sqwqx81hFWP9jPEFJ00hxd8gT2
G7r0yIeoENarMYBAV8wL01xG00hFD/vv0tXvbkDJpY6nChvkt3YGmX84mVCVV3iv0iXi86MZ/lXY
hLwTfeRaaUwKyX3Tocn3XBC/PZglCIWM5hdbM9Rsny6B6eNmc9/4c8109iFL6N51FO3D2ydvzHS8
T2wBGAG603IUeNQkswanqqor7538Ti1H7PItyW3IIlgnOxGI9C0OwcvEIAXA5Ibt1M76Gpl3qJEE
P6BUeND9cH8Bd9q3fFctztGciQn3Bo/5vbgdI+eKHz06WWkxmOiFTQCqsZqoRjJcjifr/PR0PLzo
RIuBfdSOjSMzTZJOv/HBlMgVCpwuILl2AsSxFc143SCJ3xU0vDnphZc4CsL340ySON+RmP1kR1mf
z+QAt3tIHbkv0eaKcrso7kJMb4rDwP1MdOqlfRoiXNqWOknOVSCaavkywUoA0ej1vJeRgIXDVqYd
D2x5zG5TuAyIF+esy7cQtnevFM1j+Cw4QFDxJaq+ssoYf6GKgdgAsWxnTVrHyZSdQKwUQLu26cE1
vgzaIKw4PCeCZyQJ8DKXKzF2OTz1nYg2Gdu5oWjYZ80Zl/BmUB3BDybr9lsELwhMjj98mQoKuPtc
hTp+RUgal1ApSlxXA1ne7ZMIJ2rjVTO3TeCoBsYEZkjgOyWUPWIIimMkMknHlLABIb7mqSPRgXjn
l0wGZlGqDy98q36SOos2vIEmFwspsbgh1xdtuSv8C7FheYoSjTC3Jgwlv3UPfLOAf8vq2tBh2Geu
KUkVmdt/I4DNebB6fr1bmkE05Ihh6HQ7nxM3jIvSWRm34TyL/V9RgMI56apnLSA6LvQVREXrMjSz
q7j0q2Oxm0dS5UsZjfziByt4NGlxYbDnIarERGCnU3OpsNJuDbfwUvfZnQRlEasRRO2QAgO4nN5O
vM0ptuumWwj1YgbVudpqvJPK5hvH5jrKmCEa/wJvcc5uBK9blKMmBov+eXKvPfYVtZ/23hVo9VJs
TA1wt0Lgw4Y6PmNoMYAWCoIFWUPU3aMOj+ABQbcUc2YgCmzgk8Y4zwKALf2crRJfBeahLL0mKZBu
y/WPejux0Fk1K0H/PHaZvhsDGu/WvX3yoKNXtuIIynLP2SBFagKZt5n8cmAAFUHACw/o94zBrnG5
gSxqRP0f5wxBNoHVRfcZEcwBO0IoeB3lzIWdO6MKMwU15f/q0L94aRwLTP4G5LXLKKJRpHrxAIih
qBFdpr9tpanRQHQGJm3ZixnswaOZ8sg6vbrGPqsGk+lXI6VxCLe9qYu+PzwpEU0rcALHOUgQGtm/
p1c6jlDGK34j/C2RJ3BXrD5IohYTnqkoV/6B0KLUj6GvyyPKB5n04MJZzRFc9Lb1nascoJ8vNtVE
n0W3WEcsOjRzZU4YGcK46c6e330Gux6hQ6HwVjYRnXCqaxVQnbbiTfL5eQxxDf1AC5ksJf0NjNND
tEUwd+kSYZSKMhnh9mKYB10QFm3TsQ/7TLHRMuBwVOE7Ot0ZLnL3z8mzK208e+OFsXkglxBvoHVK
XDrSz0pm+7C/g3heMew2gdsGKOFCecymPvm24gMFME3f1OnnmTybCc018aNIr5zgvx3nmRHItQ6B
gxmX9HgX34rfLBWRWszS6+6VvM6rkLzI3agwlEVkPM0QjC0ABn/klKRTkNmYp4Zj6LIRk1nd02I6
mA6Ac4jHMzXa7ZCiNS/BBaN7Vu+1/G8nRUT+eVngASOBDQT8TR7LEaKSudYllhHgewyU2M2eHzlo
hniY3qo7pD5LvkWSx6gE5xySqrkeLnx+lXm53zGcnfCZxHcS0o+jYLMoFm/CgmoiPHQ8PJzcZgQz
ocJ88C0COpaK0z/ZeLtXbOurYJzGQ7zdZkCEdxFSpqjGI60gvtm1di2erGWqDvgMfpuT+2m52zC5
DQlnozfeCtC7eQndzvBwcO7euVNbn3jXnFqIuNbbSRZvpmBiB29Ly3/sJP6exggCfFdKeFDEVG2u
Of6rmWInkZGzFwWckiYcCLI3v30+dnR69xMBNca0QUyjHWuZb+QleRlYMyNTp5EFP/UV2t1oIdsn
MZ/RQk7vtqNQf9hG2ReFzBmOlqBbZsevWQekiNkrAMUtCUnOSzwkaewEH7SVjovT7GHY0Szduj9c
eH+fHkyIpTFT+ffAxlWTypl5veuLhSIrWkrqYXyPdSmKLIxGJMWZGqkfFoND6eX76gPnNq+BXzTx
TzKFUVLyraSt3gdNxgWJNA26m/wrn53VSnzT28Ize7Yml041eu+wyXhkNz43qYdF+CUzE5sJGEDg
zZ+I+l6BpP4ZMQfqRNGso6wIqxKr7O7dz8XrMMcPreohgw9R1C5Ab93HcxkGvShD9/JYXajz/tig
RlgM5h8/NYmRkT1mowBO45Qa6e1TkTPh4gSViQazZDQNXrAnIhnfgTa6RJUzXjzco1r4ZRd6kxmw
P3vO937z+P3jKoKmHnQjvtE8UyOJbD6V4vVAfh5Fi2DFYW2bQhsF6FLpdr2UtCF/3+AYN+HQTkyC
/vAuUyPxy0zHKs2u9wX6hTwy8z2Vfmw6W02o0nxjaELAHYjBGhbhlYQaAkneEuBm4eAvlwWAdp8j
129Bg+VQ88CN+4fAol4p3Ni125bEQNsF9ddx4vBb4ZT4q4fbaeCpAYWWC70IyWSA002Q6oZXEiTK
/8V7MfF7to/P6HPuBZQneBil7QjsU2jGaXsQYEn5DslW60bY04OY6G2JVBlKgsBiaRRjoxHycAdQ
HXd/pXOZm64ZqPxTLFjyzq6v/QvDoqfGuRBK1vEDDMxwPqith74nE4mk4D9DtYhbnnVsthKwF2UW
OsXWmaVEnBxGAFGlmbXrywyVTZuf+dLCNbntYEIGWn1hSw/bwzJahZ0Ae2HCHFlnmSXrPK8Sn8vt
R+O497pHeh7qgzidZRgZWostjj4hB3Y0j4qR2kf1PaDXVcaDAesA+1E2ka+MyCfrlbtuRBNpJ6hx
LkguT8nrPwWnVJOz+QNp1gKUCEmBVe8BDXHyRhyuT3obabcL4uzK3g+XiyUen7GtaMXDHZHIXwlN
uSnG+H7vFwmieaFNNrxALvGzzJ7k/15Xtx42k+0qoMLLBPHcbfV5moJ9STjbEf5z3e+i/ivK6YDP
9XTNZFQXUTlqDKysUWxwPxzbEh42C+wcAPQVWFawj91rISQnfGbQe7AKMmB4CUAOVilDFgE0AqLO
wbp8N00cDscPPkb62M9/0kTgRVFVEtgtGu+OtPwTQmcKnNI0gEaYQ3S+Smesgb6COgYiSDx8pQst
BhJaqGAxy9nAoQfc+9E/6xUmUQTeybA7vxzeMWcj3mMLPufFhi7++Pgw2BJjh+zl4GapVj+DCopG
wtxuDAubbM6DBlOfj9I12L/5BgXfVfCHlJnC4wSTtBOH/SqTgGk3T9hmmQEUujHrYiZHYV6zKj21
vuRIg66p7aMjksoewA+DxofkNVxk99S5h3YQM+nmi/9LOntpiW17v4FP7qHc4+n60M5NLpGTgxP4
0P5kwAAb8+JdWJ+NWtiOLDP8sfO3E+wDetvwk3BRjwVBh2r7Flo18LkDUCTWHfjyaWmSG67fY6Ui
i/MxJUhkehl5t38CPXAdzWuOfU9r8dF4oFVHYrv16nwi/g/xGti/O3YX8CmVrO04MivqCG6MkaY5
fxIsATITaTsC132yotDpoyrdmmXuEzkgpr7o653CE+wUEbVkXqBmfC1Nkw105KHs9nFIK/AmIIUO
M08ANVN/4i6K/aCl0xE6tvfdCmPl/8zHPWQ9v28h94lEjd/d4rIbDeZFqH2TReLdchXoelbM3nP/
74DsN2u7d+BZD37TKOA8QmHGP6ZUG8mtV6N4J+2kLrxcv41kZbWBx7oxw/occTemUZrleGcq/CxF
On/6ii251Fy8gswFgH2y+//Hgfa8NDzXridU1X0Wq1OUVfeWsTksapdEQg0sfXHMbfBj3KKFzQKN
cD/KSgfunOWhkP59/P/4eBN62keKoLg/iDl3IEa8mFRznPlDoHXBxc2Ce7DEGdJcZPuduZ6Nsein
l1GGm9DuuXY6aT7SK1Nm3z6YaqXVOntElviGVh5mpvUxDRlSIWo48ek5s2EPU6aa470fPW8qkTIs
aqP2qHKyGTELSTxNmv3revmxZdVFRkrqXl51l+9h8LZG57pje9+B+OZwNNuYoKxXGvdq3uToG2QL
UsGjEORn+eifwhhmnwOKdvLpu7W9pvkHwpqxUSoaORHaJd0O8RU/avTzso+FnxnjUkcNLMAQ1K9N
Seh4heIjFppdvn26IuMhTPY2nx37Gz1Gvi7j9iv0YpTVN7eJnQZLk6/mWgfZ8Yx/V20IgwSOWReH
9i1Jf/4nOvi+nDM+3Si+jNRAFoCGqeENNhDwdesw3KU/WTGel2cs2hnJbvX9SB1z/6uC8es52rxx
57s/qxFC3B15bAUjoXN2AR6c313Od0jw/0c8I/5BzsZLt2xmAp4+/kAMzQJ6UjT1/y5AsvB738iC
MO+zuT6eG8c1QIINj4ksyZNU08DWA0pt2CyFzu8r6bLIr+iRcML/BLqacObYrmTpR4t4bVWoEIME
BtCPtut/hepR+Ydv1YjWgHNtPdALUmbiFEuc7bYi5dEvDt7sCzx6GKApy2pBehPc1aIsyH1RDzCs
AfdphsIkSP35x4Bm6nujsyAKH+2H3pbCjIciXkGyjDHqk834INBNU7sse6TWjo1slu86wh5mucX7
ainlXP+5rRzWhOnok4SnawkCvrwD8hq3ZKGdtxD/zq4qApjlW4gPC3tCiz01WbJpkS2IsCWkfI+U
w8spym7bIv1czzG2zSdzDU2Y7cDjbBROm3em+dlQT4F5Vjmd7vGTKqzEyVZbvJpRcB7FwAwbjsYh
pyG4U/BDaWClLD8+k7cBnY34ZoWkmqSgbj2pwWBndMb0FTu3V/z9wcfvJEa9g3vAwDKW9TZJgUsX
twM/i/hfb79eH+LON3rYQAr39Q8buXjcYvA1B5oi9z0gdmn3al1ejRUMn0Xo2dXNZUx8rDv3VXvE
Joa68rTzhfnklU8kD1HomYFSjQyQdOZvWTkTgL0eVcj0nZ8TbSY26kcsfSM0tUURBh90dD9vsZuq
pOwsfsDjtJFApL/q+ev6cEo0f6SvqCYVsshprVBlucbe0+oZNmVHU1YRCHk/ElqMevAwJvtge/Wu
Cqfgx5XcZXZvE2DBUrTd/Js4Hp4uMwSMg6zbxvMTFja5Yus8vYCBbTnx8ORrKTGQFgMlTDVHA74P
Gi8aR9mpqooiLECp+RBUKqgesP/62mfxF3G6ZaRLnIf1bEL8igvksj8S1aMxWknDUo/+6wEa2v34
OUNOL2otDYSGu6Brf6et2ckABc/V9HUlkM57iB0oX04Pozd/YqASxfCBzjNn9tSaGEGcHlJL/lbF
oXmhnGKOso2TBzNxprQ84PFFcbmfoDj18w14hRoHBH+0Weq57LLkb8Q3wDXssQ0sbX+1ya4Rpzcc
TwpG9iJ4Seec/uBN8lwCkgMjYfXQFuKDEwQiLc+V2u5FUwDB4Y8iCPT3GHXCcM6CQtD6vVe18W7y
0MAuKwETL8rrpL4LgCvfwjoHNqlQJ/pfI8mp2Ssw3BdA6f4SCeZ5wsjPCBB1ubQIrEuH56XnlIk9
4TRJmwUy8VjIVJBu9S7Az48x9Ysz3to2RWsYukIs7kbxOUCw+2En0b6TfzalavRgzQZPMzUvzKJO
JDZnp0JG7MVUiuxoWF1ACnot5ljTRqJaSq4zUy+BRY38AK929O59SXvNeFiIZZuXhkiOI8JFkWlr
39ZQNLZgoH+FD3fZcT9fI06HLNObPuOWJB912e6CFh6kafM07c1zI7HINta/INTfKgyAQsysZzXU
RO/Y8/9/jgohG0w/JmJT5viZQxvNP6X82LrPqSJYAbYDdO8ZBexBM308UPQ1mnI1ObdM0CI8ycKk
GsgUnhvb9Jni9PK9Xl5jeo/xVRsQdXOdsR1g6iKK0i8XLGzXjmwM09Wh06/I6AhA3JdAaq0JfD/R
blK+MMD/US3Am50I/AXqi/TKP6GEUw4gnE3Kc53MW6mbmTTkSpq3e6fZLKvybFashnpH+Xj2w3Ly
c0W0MNegreD3ji7C6X0XohKrVUYOifce8qxYatAfcoMPJQPREOgGKbmHrqD1Ycpmq2imCHzCZb45
R4UtWdkOInKbY5CDMTaQU94pjOZWYI9ZT3DjEsy4kDo1MQiXXdf+7HiumVfMn6mxRowec6zJHK1o
b7qR7P7ziwJQX7kJDFHvvn6AFrgm1NE313VtXOgR6z9Wz9a7zABTG8AMGkzQKCzYNulw4sWBo5ui
KPpZloFF7SS/Cd7/AebtQMGaj43Tw7/PFAFmyfXZf7RZWmdWe/w5DRcfwPcmoYQ/7VibWDfd4hxW
hYVnGEPVjXb5DHKShfxhH9MqPPjLhQKFx8bYdKtT1WeseLxHLqGNBlqXfVphvQeyU+l1YYeX5D6E
9TpOIraI0y92nfCCAAbrdfzkocqwEv8LKcpWVuaJRD6/XLVmuPSQank1vhdpUNcCj/WQ9n5RQAKg
D0o9Uph1cZ1hybrk3FlNbS79mzult+kWwflHaSzCCV64g+cxjy6wf2MPWo7FY1yf8wJFKRGpuHi9
25ZlE6tnj/Het+8292vlHkOjwV9WQjA65reVAKTBcrYF2Cnqx9enrklHF1bRunHG8olwKIP5nx9B
JXJWkYWzkjNcWh8zk4fe7HL7mQsTsN8fTmW5e5k/eOQ8Tr8mVdb4TaiUIYqC1AuS9XgUxgUPEbrz
52d9DVztm33qRXqIZ+8XFK5825orssnvSIEICJ6vjCdE5hwrHtIOvqrhAy13y+fRxjbLrDL1jd6a
V7u6nEU+qRxhZtZxEdb5YRGYUJniSXQt1HWjCiaCRIznv8kjpFcwZJQ9byeBLC2GVboxacF0yMlY
yBvTqQgBGq2GVnoR06uECIgU1w5pFFMsBLFVTT/FwpEBD+PIM1q1240SSY6i+kaPVn3XEgZND5t2
PzYuMQOLAc0oM72TLktB+7UHwKmUOWcAJb3ouT6qAPx0vSFdYjCVAGwaMnO9W0X7JHpbhSXIUa6p
Mqjo0x//pgsZl8bOxFui9qmg
`protect end_protected

