

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
jAc2elpDF3eoKND1/3jp/zR+PqlylbAiYUxqPEeJkonmmMj0p4wWQxczZkP8HQmv7tuBnI5hb1Re
XvZ7MbtjgQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
NcCSQniKJvfmu7+yh3FyGy0Ym5XaJUypJ6Y0uQPsa1akcjYi0ta/33mMsV5QsYvu+JmAYVNroROq
Kz/qydAoj148DuSUxGpr/Dh6K6KFEJQ68T8sjkHECM7M9i1ksK/n3u+J02M+jecJiy0HOyxQBNjN
TYNC60RH/oHr8eLrkFk=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
bUAhd9meaxo49J9KB0t7maJQYPBZ/miilGsGpP50LlxHKsJESMzras37N6FY41fj0BrwI2d8gwNc
EAnUne+xYMqJWaUJpkx5tkU3/Cq7YHGk19i4FrTEgtDQCfuJmvvnxIjd1KLqJ+tz2Gc83+JpCcen
LoaQjHQoa/X/vrkqv+GBi5yvXYw3CmPRVPihw2cyPAHh/aKqVK9U2rN3QsJFh6K1GPjF0J0zEoGU
HwvENWUy5CJqY+RhFtoI4cFMx4zvZ9LvGAYIaSHNcjGEuPxJtjqEiRDoZaxAPs4fPiQgVWKDuDze
FLb5NkzGHVW3Pw1VKV9puYBInovkYfTC4nb12g==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
yj/twyTkVkmohkM4L+pOFWHFJL5INTv01+xvkfId4SWEcQdYpyZZSWwRohyHdzU487emKgHzTSTy
GFDvnAvaZMJxmURlvGRprcX/FxMbqrYJ/QXjtyclneLv8hDwZCLiXegIMxugiwW4gYlZjMaOoPQJ
gs8ya5IBC3x9kMPV5rU=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
tu3CqLR7y72d6lMu0BtbwhwW0WER0YZdVAODwj27MZbWzMWHxGpAy3KeDW2xQMQiri7N5lQ02ec0
GWpokUjyJkcJKOv6cAVA0bMYymP9zM81k2IaifDaYhtB5Ah8VbDj/ArIWXDmp920Nuuu8ntuPKBS
17ifrJikBEgCPNkkESl85/+YxK58m3UimCI0iHmw3WvHkIj/sAUsakbfIOXt9rbFyqcIak6vi6kx
Gi83B53duhddmOvXqbhgzW3SRCCdyG0CtC/tlZjBXsJNv2kpjQBMBZf4BiACBpRjP60jLswfeEZE
bWRI3cRILGIwfm5V+sLTGxa0jiUVbd3TzGM7gg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 14464)
`protect data_block
zWA+lYFytXEcDQxPXMUQYASbVgyEr9PFVjumIsXFk1MoYj9t1of2Zbgn6WY26dqzN1LPsfTWPfrh
3Qb0t1ekhlEBA2WokIIkPGhotFbR1imDb5T6rnwwhpUjdH7oxHQlZ98I3U49+FN7xdt1wFyj5McU
A/MgBnoV18k5n/6MxKgMmzaOc9JEXvAPP8LyPUfPeK9KoShIxZ67hmtwgLyXDuI06v95kstWKlXW
iDWlrsMXmgI20XGcxLlCqjaClKKsnZ3bR6iOxZI9Y/5M0yfcguOJnUVe1c8Dq9DkVFfCZrPwfJPZ
//i7URlvMjkuTB4CI50Hb2OCWEIJidLt5b9yx3Knl/lgC8M6gGd4Jro2kxD6+iOUJMKm+Q0wwqAa
y/mTFrizaNU71KJqdiFj3i33OvkkE+RqjEiCmyP7NIyPRwhCZzkeen11JJC7OEhj9seodgX7aG7r
KnEmhcdpbAfFvxSSKF6yiYxeJfzPzAIBVOR2QHqUUacHu43USg8H8oqq6CKcq3AIGPvYfgrSCg10
/dhfoZZxPSJ0STNXIg6Thh8L7fXWRJJkn0bZ24Wo11vG8Imzc0e3XIE+SDXuZpmSNhJgNN+jAMon
2v33ZrjGHzHrKQ7XCASt+HO35P3DGihMfe+ijGRHkZ03i1xVT3ypVgVPa14pTJbWjg1AKDhKBdMY
UctpjSXR6nlYrpNjWJ5I/EatF1D+zIuuyuUqaGMZwDirgoUjCoIwcmV7To6+bi3OboJq+10qJbsn
zDFE9HVlPcdkeZpQZjQ6H399b3BhpGitPgX9D9MQgl8UxWDQzxbUYL6YA8tynFwLCHfc7t22NsWu
XypAymvUYdNUUM5d/+Us9Gc7glgwh0XjpeyaWYTB52+COKVq4s7lxv7X3gCnd8xMhU9GQj0wI+wA
GJv7E1kYJfWbjg+J4lOt/mz+DDCNi891knr4ZbyCzj59eqjWeSUoPuuLdldaLa1ouB/a7/wuOcNw
Z8pvzw68U/woCcYSksLwh28Ci399mnCQnhhC6Dxj69QuSi113m92ruF+t0MtHm9qVWPZIBZLVDSL
OmhTWczUr1DgwNsBBVZkjuuGHUZwOFcMDaS+buAD5pMpyecxsjzgv2MBYYlkZ1VtG73rgOMqBUwZ
E6nk137AjRoxGckhqAw1LbDJudD0pkfSeKlW1K6Aps3xQhZiBsXZKBxzWplteOT7pTzH3eBihRQh
MbZauFOO2UIQNrRdK/Y8gUqK1l7ZlohKd70+O+WOo6r68E0Y0lmFaM41JKYF61NnraqrOMGdGXFJ
LWrKB5kMrSkO81oKlWLvwq5q9eL9mWo1/juavVpptOXULMjfKCAUht9xBo9cie5Lox6D+yOWo+FY
AKuPlJmhplsSD7RlrG7ZSIaWEw9tuHJP+FtlnXJYewoFDV3McjF9rNzdHLbEVfu+UFBQu3Od7a1y
qkwcjpZKRlKVWKOC1IPDOQCLSCR1eohKKkqCbYeagoT01vIAz46rT72HYjJa7jdofDAnesOdNgNn
YtSBG52QPdouKZvrdKIH3VeQEDodyklH36zw16lJhif5zpkvaZQyYI6hl4i9DMi8pQHzXrbluYpW
pFX35JGrL6kwL5TaO+l0H9CKrmo5OgKF7W+QtIsX28eqWr0StX7fMXfAxLbi+tixvjSZNqR3C803
MYu94hXl2hDN8u2uhb1KIQit4vKcHWVKM+uawp/LD7sMbV1gZ/wYDd7eiErD/fsi9gbA3zFvwyLT
b9lr+31Cdf4c+elLPSjQnD8jxuYOuyUw3GSE86a7nnpooy64+xwolj2EyJeP/cbz5XS+7ZI4XJO6
Z7sScKHB3pXUR3/U+F1KHbUfHCXm9X84O/etOV5prC76LRfBs8605RRtrzCFzVDlFI5yv5Fvp/iQ
We2aFjjZU66bMEH7lCTixBnI8Mucxu9py0a4qyWu/WD1WUD65EI441glv+B8ncTc57N+Y6HynKsl
Cqkic5/vPsXo+yEKXTd63UIaVGS96cI3c+NA0nJzvUeB2GvplU9qHYUK6eBKDc2zutpv4+/wt14x
sfDkQ/QmbyJhMKlUyFiGQTydeB57sg9AnqwxWl3eye4lvXG24wRAq5BNZL/TVjnzSq/FkLlVx+Ni
IRbqNafKA+H75HgiaL18mjB4kUVJGEPIMLjkcDYds2w6XpNL4QGWLZtX76042jFTIbay05oSnk3F
Mj68dG227k6k6l6tBC17PUwJZe1l+G4HW+YbSnXYZZzi0ah57GCU6EjphRtM5jbd62qPrAhX8e7V
TM8TAwYFa15UKR9+ecsi5We9P5DTH7SOp382EdQsdRIHEy0R2iKiWMHnUaEAlk3npE+UBRkk8TMD
QuGKTSU+vSXQjR44vEfz2suWCXIKMItcPTY8FUvOU4+rjiIFjlPL+3l+/dUGVXTCp6OI7FZYL9c6
Rrub3u7MzdFoz8l44OJzsNuUgJ2CM6gwEPf3kbrH4Ej3TKt7tBEu9GsetuVTfF+ybOIs9zd0TtKk
j7oE6MndFC2m3lsVmz+6awHxCCF95NQqvUh5X4PT/uAv3fe2bctQ54Daj8XQ6I6A3EGkG2YzrMPe
7tSpadk1XVg2WPb2qzDrtt4xSVuVnYJvgMKhqlIXWpzCW9G4GiR+KaQTIECV8tYnkUVRK1D7H4y4
Qivut1KAvVfsCMw9kNhfOxos9Ly4s3CkL3AQ7DGZGSOe6ldla9Hkfh1HB1y5P1+PIbmCTQs7PSik
cpJFi80Y1IhXtrT8K0EeYCBL9FbDEX+7fKhH304I+Ine/PMb58SoMljcB/pRdN2r0uWVEEc1zTBa
WKA5KRMNNgUDXo8RcWf6mH4pgt2oDa8SSf2O+wMDMb5qFSI1ZOMgfDfGFsN3tqiDv2yTcQ6avnYv
i910GK3jcYdMjCSGtfGRS8IOsp//lKPzOHOD851pwgYOqXvim412i1GOW9MymQk1m9LdxqITe4vp
IVFwQr1gaNF+viqbl0p2egoKQZYsi01B06YahUmYjE4q2n1QiJcZhzYsazZ53qp2tw/bDL9Vk6ot
XzleI6NSdxzGQKd5ABYV63LjxMLEllhtyVgzvMtMv+Iy+tOlmFG5wm+gSpRU6geIeR5tmfWhWiZ4
pQ6tXFgR1Jkl8iyTo/XQcx8U3SjgRDAgct+Ql5UDgFU/FH6/M9AjhUyTrSS/HaCuZhkn2jUnr0dO
A629X7qYuikDtsl2Gl38s04P5KcZiTn4771nLag4PjMApqruUuadqU8aiWDByAs7XKKdHXtobGaj
luKZQMwKz87sUQB/2yhHpXQaWDxbNMkM6cKzISEqMUR/okjVIzFpTLnAZI9G0TPLcIjZ6AhrLKsr
k6dP8c/pjLoUlTQkBiYihaJ4YrmtfrI8UPjK+3tIix+2Buxk0Ys5GErtW/8gRtqtXpF4d1lLIPB1
iUJCErNydcr6q+8Z7M7BJFN5gOqR4H29JBRMmB48u4lYumIL0Ec8wW1PDBUV9IqF2NLhXQzXpzrH
V488onacUox2nqSFzt2tzcVA9g32zdOmR/Sg0hPZx59yjLeAEB3ocYULoo2TmVJabAkfo4Ov69pN
25nVLtEnjj/tuUPSVcJJUYa40XP6YQkbwgtBPIkuMve5woQMp+loIHZxKcVa4zRHuSiVUFu74D1V
mLr0iyy0zLTKZ0UNdCtCmbVIIlYDkzqfwNP1ya3E7KcQewygIQezmahrYzNHtJ6MUN2fYMpSTx82
gv1iFiAs53vIXznAm5EKu0GKLKR9WbTibb8/r4t1HHIfgWQCqBdvQNjcTWAuyYrEDsPZ2wDgjFav
MgYDRLCmrtmOfB8tFG2qWNAyVeKTSLwKXPu4V2ruK3g8gZshTYg9UxfJQ2htbKhSe5ZkNj8ciDB0
riVPGZq/M0YAxey8H92v6WH5FaeXEAqDRMXa6E4rhh+MWvS0Kh9nc928ocJtZE1/JwEGiB8lgbNP
8rrUs46avgew54BdfcFRzG51BoPa73ClhP72/zf/1t0qBTG+M6vmrsgGhuqpcYiW9uZOFf2OEMkh
WQjCdEaRkxA4PQu8JKTffJhITJ5KiLXToslHUD46mqpJ4PSArUscOuPxmJHMMNme38hUev8fLA7p
wO3uUocJ7wC2eMBjHARgdSJ68gVNzZDms3dsnFHgy6PL230oceD3Upw500oM4w0BOFq4cLnVocsb
ytt6DY6tUE92s7i6TWgTnWMHMQdUE901ZbpdrVsUdJViQddSoiEzPtdjJQxelm3LsJM/MVcbSjTq
OngaUojBpMyAg5ym0n8jkJIUGOFFHl3Io0fSihUOnyY+q+odERA6g0DTOoYYRw2XjQDnPvaCGKD5
CH3ayyyXAFJKcceowIYZSeC9wwKcyA5LiH5DtErXjt4f6TaYV+DT60aKH037Yf/7l7RNwuAcKM08
F2I1aZiJvtHBkA+7HrtVgB8oITzTXZ4Yfa3E1hAhRUomOsGyvWY9aHR2H5Hd5Zn9WB24JsOY87h3
RNXtOskxOr0WHMVNXddDyUiRuPoBY0g5BYsHYtP6FowCkyDjzloRlodvP+FFZhylN0VfhdsQW9E5
QzDREBcgPu3VAV5jbPTFPnqL3CAJfDkSjR/rcK7DjQezTzbE7/EjLFCQR2rwb7wP9mKNaOY5ZWI1
6jKUNIBuo5gzbdA1K8fzIiQWvZZkNMdtS0wIao0oFTxdvNvhke2nQL5XT7V4i1Sjj0UCzP2cc/oH
IUDCcvQSLrc7J2gUN/WPhORxxKJ9CVmcc/PmXu4k6WxWf5WW/LnoZDC0sPX3p2j9T73Zpmgv2M22
jq63aVVYzCf3Ax9xIubb1SLOD82jwEjwIoLvHHEWDjHDAt8aynjM0Rr2iRjszIZqSnIPu4nz/cSU
oR80rWiY+C5omMXzpcfIbdcGrLHaoeEeINZRFUqKywMkmaWMY6nxzEiDNUDbRco57tu9kmBrYDWU
KpxiHZihC+vRrR0EkHvr7tm4+x1ofb7OHcxUFMunw9/8p2uKEwxv0gy76K0PgWvqqwYFCxFQyTzB
rcDIgLgfG2+rKiGpNljktRyVKr9xyfIXgZ7Z0Gkud6FNG/SHFvyVdp6VaiYh5PP/ln6SwH9uwlnw
M0Qol7HFnfDD1BLJNLAkM91Atbo9bL7wLVzFCyoB8slHWxvI7U/7g3dGGMXlPcgdLyfrbR7O7Vzt
Xy0LH7yf+eHPtKd/O+LkiUzAoTxPQF5fAztz3tNLmUTgMF1JKILQbEHbq47BQgM1nmX/9rg2Xm48
KGiGv1DKd9+LRVuvQVpaoIa7Pf8lfNOral2uwgZa/wCtqIOG5lsbC22tto89K2wmX5uV003xoY9Z
0ppegcnITdz9gcdvpNKEssALJZK2GLLSrPG6wn8unR7rB9FhZl+5lMAujX3sNsUb54mL0Kz36SoY
DNSipPwTJ/6jHi/8sa22NJx/nEQiQEeD3n3ZLnLEIZ+fEZO9ARzT9ny1bXhTh4pjl2s/d8hIrQSd
iLeXDigCvaNcwNN0Z18SZUVrbCzJQbor8P8BMZFoxr3e92ZGRt356jdqdWOL8da/qBpUReHNs7mg
8C44mCxA0yUUJOmkvUUG8mWTYZFbHj8LKYeMENQ4SsjmciptgtOPcKZrj7fIBiOw3pbTfjis516B
5WBmlO6+J47Aut+wY8enSZzHI+7idQ7EGQPPv02U+eNPAW32X8okhChnzmYYBsVyyEI9MfjRcNc7
TPDooymueICLMkOApNFSXDxIUhts9HSASrq1au5V51ypx3RaXSlJlvcO2bkrfdr6pIUHAMpmDO3u
a7k/UC/PXufxhYaLY5JHOivaj42pZ7ap2jiMwLKRs/ANFC0qE6j2+cfONSwrkzsrFiw15EyU+BG0
i02TkWImqOG+NJd+02k8PhOHhnOiG5d+F6gId25gbbXucKssM2rIK/1PL5MIMcylU0P9wXFRO5lF
5DFLqZ4MDWQizSIrmPUQsrSrr2BRVH+PtblHiQ38QMKh+skDVPbMn7Ufp2y8baincH7hSgWJWs2H
3k5fuPayLhBjTat1yl5r/P12/TYAX8ygFga4TDNhqtovws+oGwubeeq2q7/YXTGuhPxywYZbmxJk
dXhT/pFhPux1hey1MMRk4tykf3uPbq/WuOoOMnNzrRq+d26yIIB7P35EonYLIw5SFFOArk26Pk1i
MtPkEMwPg9ct6Kg6hA8nWzx6u4yQaFuqtia6Z8whMGkHTrZR/6V+u04frb3GL17gzZVhI3AcsiMY
2tsVk6ipFS+XyuzdQoeCh7Mt+OnXWNTaQGypXluoCM846uAsND2F+eTZ/bUhiRF2YgQ876cuSagN
6rmZW/ScXUex7adbHKj9Dc7IC8RpT+JdU0b+aKSIl8+gqy5SUxLVyr5VHfB4uIebTMThL0eWo5GN
B5d6DG0D1tVYgVi06II/SZBBFgR0bTwdBBp+yJsBe9suhK9J7sK1VRDVG11MrAhGV4UWGa8Uw9On
xPh/EgBx1rGI3AYZxcQuOujwQBLn999l4Gj4tim7Z0qw0iLT1ZGrEvvIRgVuslyZB/xEiMsEHzI8
+2LkCRn4JM+xfqggAvawt8mKkNcqejOCPVZsVQyC7pZFyo/Kcd/f5J9MqmQr2aP+yk/ykPAnK9ro
l8/14V0RXxUHnz7+mPvBT1KmNgwCcWH776LmzJA77bvuT4aZsLoN+MTja/hZiisyO1DTOXWr8FYs
OUqTS8mfg/FJm2dgzNXlhc6AjoQjw+PLlH7mGbcemJQ3Mrj81b4juehQfNLag7V8QLUkjUsF49JJ
NF6nVaedZlKDplu+8rZoyyJKSYFioGkp1N7tfO1GvqU0vNmmdIZHehJhGNpWBl68b7Rvb2qoubYl
b/3TmAzQi3K8tbOgfnAjfsYjHfvgD4o8zpn605BPmhd9rfriw75oZgQtvFzlq3hv4MdWzr1ChyGf
1SwnULj2dIUjoqbV/Q78kkFAgg2SyxUPfvnzyIxy+VCiyxsepx3fV38RMrHnXnARbcuOkJkEIylQ
MXnhXSdEaUPl5N0/OrpQQ10BkyMaFXgi4HcSbKC7/vCdYBuCj4LyfbYWfU3w6TS8ffOZ5YO4G8uq
6X2LoWmYDFjyoVTTA80fKMIzrZ6TrtrHzUXW9woJPGzjTXHfuEK1lkJzoi6eCk6FCO9yvvMSNFWx
1v/6zAIG0h1OBneQnGyhN5jtLe7vfAS2RNvIzCSUryhRr6C3ZXIIP2Ylr0QoUW3dGv7Vjn/hmqNB
IsdM/fY0Za3n7h6dIH03FB3fCFpPqosjUAxRWN8MlOtbwXRxnwz+j67h7YDvGFJ43gRPBvzNAAv/
C8LfixVw4UZ5DC8q6FyV10wfK9UWkbTheUBuVqKUt4AXCmbiJp5M8XURAqqeCKwh8FH9OZQptNr5
b45uLHkaf+2sZuCOhzBsdzLG4gXJ5rntgH0c69Ff+exsTdVNHxzibapd2m83yL2DN90LsUlWCaKA
rtwimIulrBzcjdxQ+K00Z7fMpmdc0Y3THp5bCfXObNPLDCmGAt1gHlnQ/P82eQSN0SD+hI8bjpc2
IMKmad53CntjIt2fJkEjuVwJfmvvbD+4e4qSGp1BYA0K0xi8LkUo9+PpPcBL8LByRnwvmwTX147m
691YxvsW+EC3xrNtNFSdOhQ+Sj5Yqa+r4pv95MEn4iEjCrLtid2NlAZqx0vYaWiBlMY1GJpyL/Kx
3bFyKLj2iTZMAPkoNgjEODQ9qHxpnlm997ii3DtfwR+68QPNnFkyU8KoAna5tcy6V5cUspfMvxtN
UfOJaSnOjk8g5AWzcqsX2e+yhMmguFu0P9KSxNv9rpPZix8QEsf785lKLzXGdz6DRtIJY3m6gA0s
SLe68ea2FQTamHWtaOFw31H5pbA3wdBqZan2YPu6kb7HTH406h4qJ+bsaluhnamRY+iS69yl7pTU
jML56XGUhJDX/wiRH4cZU1xQ0ZcYt5pN0KGGN/NYvnlTddr4E7Jli8XQKVFOrqp4nAd+Vq2iUGRd
G1F1TfXNhlQ1DeVxglcBVjz+mKK8v0LTaLT11JS3ooJDefXYzACGCFLvxThP4A0qcOKcRpl4vOxq
cNt1imQxSpEQOjZzWFwLxjjcLxEgNYe88asuM5lOi89DLGNYlt6q0BxAscggMT3wiYFjYSz/TotF
xNhQL4TBDDlLjhfJVmw/o20gRX+hXSmYKi0yy2ATOSB9hl9wdFYeAtnjV+dby4GimcjM0HYD5ix9
UYmk9RAO/WCTRsYNDT2hpmbG//qUg7RS0QEsX7mVTvDXmf8jHecrlGOVNBhK6+F8hSrnlm0EKC7v
u3KMDa6S7BhcBkB3xIH1kvgg4/ZPIh1kdFP/7sytMqeLqG5oub9nxmisL2/zac3MUIi8nxe3WTX2
1V/RHs/KIypn++XJSTJx/03TUHEIVvx8X4b580NYTPRx2MpDiWavWTdrbF6GKLpWjyKaKgQXNZqf
nAqiPMzCeyWBX8R8TOMoT3w6QTHohYjT3oaJs6cO4njucbe/33NTSo15n0aasTvE8TmUMBT8Gm+x
+yudlraJ5aOk+4+JcAV3SsJBNxuxQD2eW+9C03MJIZeeyxmbA6CQtB5Ph7V6waUJjn+d2uZTC5Cs
WVIdeTx6IdnVbMLY5Ky2FWZ2YM6zizaJdrFVAX/tRrpi1RDHqBWrM07TkWYXNHBU93NwKHqZUNS7
lqWn040eeljJOaiE0+uov/zOsUu+KFfaVqC2pUHJLYki5oDMqqjDzwdScJJmOi+Ryg5VDZ0jR/U6
G3d6XuZKxvUEdLPcO1hDMfzSRF0N/XXW3BG3zoUxcfpIByc/X07Y6A2DXCTd14UyjGnpQ25q4AmC
/rovMhf/8OOpMyVhT4tsJMOhvppQfQFmYNfG7poFYPBaV8uQ9fxWXf4LL3LcvRdylFRwcGlbdVMt
zCTVanDTr94m0YZfmvyFv3rLHvINd52o57l1i+96ZA2bq77B2XiEyn/LKXwuTwHsvLlM95XVnOJ5
BJHZ994962py7rssqkDAraJGD0trOTyzMHBqgrXIYHHn8qpXPYOWs2RuXYHJhpcENQAoJ9r9qjyc
VBmuCDLQzOVduVDB0Vdp/doM+35/pBOn2ttzC2GFHuT2LUVKgnigJxSjmwi7vs0L6YyoiBtg2ygH
w8oGFqwOwpewc/LOsSxVFn9W+VcJfx6PTxE6EA5N9fK9K5PcgyD0AxOPxpjlLuUD5deki3snGOwn
q/8OzaWLYOegQybCGnS2edfpOwTRKc6M8oPsgprnoBKM2bMqnTBfSNx0UNw9o83PXHfyzyASFc+H
KY50ZfJ0OVRsnLUU6bPhRcl4Ht8TlGf9QbJTh9Y5EGApmTe6WBTQL97fxPriv3uWxDpJgE/g2Yg/
IeOKLEfzQYNPMXsvk2ZeXvBxy0HeOTb96Bu7L2+oiL2ZoBRlW5PxJvT73mkJnzqyWI2b+4kxLe23
xr9A5/lHZ/ysVyAOSOcOQUsM1W7nj3Iu+a85M4X10Eo0yyhJKYCHCUT8ZFs9DEHfdQ0i36Crbx5i
TsLJVib6BSiZgbPcWP1HH/CDR/nWMsXTTYZbQqH1XU4gKCjzbZfSGvDY4barJ2meeq8xSytMOQXS
JDVwjE63aDlXwzQLO25S85wonzgHIMygmoBPdNi7dilNCfNI1hwU+TUrReUWfWHQfKoh295L8zW1
4hcJvHP3YL0eEmbck01HSA+mRmzNhOqwrcW/IBHDTZYrwgvBrkdTAEV3XtAKCxE0n9bZADfzzMpR
SwlIlPtRNGvss8AEPDqOb+BQ35TBoFDt5CjtD8KTP+4o2mQeeETHdblryeRGOZ6thiz4O0gzrLxc
q4MMu7ttM2OftaPjY/H/Tb15H4qwLng8fEeQcy3WaH9FSKT4GFOeu/KCtGYf16DjOm8qlTmD2mul
m8UX61ucasCIjtOgpg2wHSVYzvUQXjUrVlllYDvparq3E28FGFs1lD+7rqlrxplcB0/nlNWYRClj
JGvJgG/ZyuhM0vufUIOT+U3C9et93/msIWxL6AY4hLa4lPo83IA7vH7sYj2Bl9p/4+2YNQs7338Z
z+uQIVEuSCHWmYoRmj7p2mkZWHDeHzpSo/NnxVev885qiMkM7aCjFPBoKTh8FDup0dZVWt3ZuvhF
BGfU+TFpHROo3LsFWIqATn6gCqR5kPLELD8HaNPi0mirB1DhsHx3dDPbhBFf+kv+tzi5imss9YVV
warbyVPgNm280IU6RBhDp7D7hM5pjj+8JSzaOT1DNIB7VZCI68cHDhjuzXKaIHhjMO8QGO3uvQZe
l6LTLifv6WyKyOHtA6rDpzSVP7BRcSdpaTMc6MlBHv8fcJ/Dv0sfGUZi2tmijqngdQ/idViU6M1p
mX4SV0HaerlIX3GLPYmjYFaUCacV/N9pgbSgjrBgXgV/uOiV3WTKcfe1u6fjpTogmx6cwcu8bIdW
LFmM3Oj8uGErHcyJ0xXAkOIy5yg+Ya6e3tEnkeSxXYnt9FMyy8KY+S7rch2ihiqtUXxHOQwJdV37
geZDcvHmS46hF+f4sWgLAMfvaAFa1RKmJ93cGLqf275pTP+yYrT3r4P/Ra6vZgr1ZSzacN2JXyJw
nPVhjF4KqPup+bdh4Cs29JEJQr0UpVAveJ2f/udPkjLdSSoXClZPwDJ+fqGgJLQUyjFbaomM8KLp
TSVhMiE8AAAzR6f3lYDhTtQeJQ2CxIx/oPQ3E14RE4gta0/hiX1wBNOccL/hM4bfsBqTY5u27sl6
4APevo2Ll2ncmYtVX9TIYai7o6Gxy1txMycEI5MUn8z0RPseoDXzmDNU725m1m/9FER4qHIH6ojr
C8sfNMaeqr6LKmG3B0rezhLBa9DcMqHQWcbbx/XlKfrw4cVFAXpNHxiUgJO8QwlBVIYDtMYcrHK0
ckeJoEIxMAyz4wd9CL85CqfgM0FAeNahvzxV2KJSO4RBdMCsGqK+IQTWcmecf9vKzyx7+Ak2xnmF
KvH5n/Iy3+IU/K6cT1tdHbH/Ilxkytcq2x5y4uJYacIy2s4bdeMMrQXp9+WP4RBSmqOFvgltj9jr
jja2m4Dd8pl1PDTm3bDYbD8jMiXaTXL30f/fWKCVrWXgEE1vwHvsIm3F9gzlpdQZb0/TEi9MSNDH
8s+l21i6plm/mnP/3E7YMJnxsquToBDmGrqoPdBq2sk1GdKMzICmM4fEMZ82xBCjweJO383mx7My
gC597TkWIAAm13DTcqL1ERqVwM6Y3bOL5NpSJHgUcJOB1G/6J6bUR4zUpysVOZuaphq+9HW1tqXI
zspxRFydrAP2ejTnvHnB5z1NEJOzUfReopV/JywH9c9ebFOCmzEtLgJ3BUMmH+dIDjjURqRr7Gu/
bq69SvGT1JosSG47pXAfVpwWvc+BmlV6k9oYOstMhJJGIHnp8Faqyo/ZF/lCTcJFSK0Jp2mhSM1M
zZUe3ZitCwYazHzXPXJbSE1XxOgcGlpcFTAh3MOEyzbkRgvzilH+fG85qUNkCwxfna07WAs3+qUM
ToTltdiwvx1sbsdFPfWPD1QSiXiz3sXTlV+jyN9bp9CwoptztJT9MdTPmTwJGvDgKTWHbz79zjpH
/mShINVVGza/0qiswapePZh538R/7vx2UOWBLQPWfVGRaBuZKrkrVqR4o1FMbXKMx2Ya//g6o3Re
+u+PWd16kijgavuAC1CBqCIRQl80VIgu7Dp0T0+aWuumcCRjybaleqi1AgLdIpkpUDncylGyEvtk
LEYBKwgVV6RfI0StFcLJgETeGz6d3twuwrtmWtRU7mSg7NoVwyUvHy3FxrBc3EYUPKWLLOyl0JuG
88zgz3RnW7JjLfBehS+bi18Ao8XiwuVrMu7iJFjSDuPB9Ge7T1P3pBp8rkX1jMbLjRy40s9X0krC
W+lGkGiplaDKhOnKaikTXc9fgz//t0viOzM7PnDQ7cK8ZuEyyBRjT3j8Hp4YhqcspKZEF1wsEPSL
meMfkonV/JPILwULxsTF9HAZZ8OPyA471YpodugCttG4kcli/Ju+2toQD6P/oBmKvANfUp+Ux9GX
ATYa9dMNgzeJAK0tELR256ZouWDagZznzduTyBvOcBXI8m5EJygH44zP9GLKQNUgQY16VoiDVZOO
GH2FTdAil7m+mBhMLk9A9Wvt5yqT79e58jd9QY0iUXx5lLmzwVJxAJbx60MuPsnZJ4f7SH7DP0Xz
T8S+EahX4pRoFQwaNhKy9eQo4LL7eD7Lbg3wU22iDTgzCF+qx+8FZNgR95hqJ1cgxbrqMIWpSKMt
rMoWwkSywlBAkbxqEi3HS3KW4L1tQ04FzVeug7lYNNY4bULHFRki47PJAL8HT0qWlywyd33iLnio
ZSF2f0HcX9RGl7xmfO07YcpAniW8CI6akSDMpwiQJOx8u4mMVOxrJDD7xCwPcF3YyH4qaJ7yWwnJ
4atfjNoMnDTENFLGF5GKwXn4ka1Zy1IfKI9O39H1PDFLx9dL9H1aLZN6jiMhvS2IjRqdHxG69Fnd
/GS/HUDl1L2hfCcofjYptkIS28D3WkodwRNydTZJ6IZh2O1simE6rBKMmfx4PenrLgRGAHFpYp96
cs6Fbyfvi2y9qzjuXYcG/WJBr3NW8LLsyul+TWZwTOaCyl5YN2CTItJhnWJ00/X3F4/ewcTOzEvK
uWqyxve7beZE6UQzGSECoPqLnpjMsUQUtXe+rKnYAZBPilmWvi8U3cWRMc8rkNcRwEJ30Z8wd6qL
Oz5itVFikxpj+l5HU7rPrQtgY+3Lk8ejdu4G2ejDAH1hA3/1auOpIi293sY5GMQyZj3tKq++QmOa
HiUE/1y1iR96fbi/CwSTXMW5qovKqPPXEtufUpXSxZQolnkTNNEh26mKkoFYnRwhCLeHpqHNkESy
vL/6RhzVjSnF6eD4+MC0JYop3B8tNo9q4tB0WapArK1UuBsXS4tOJ1FespF0H/Q2WSxvlYqJxjiQ
8ksvv+VrK3La8PkbdN+Q86TxBCDudEj2CiNpLqTt3lDvaABLogfcq/+eg5fIGUJPLFxWV0spi20d
f8HUTlUBvIAnC+kdxo40sTeKoxpUSf6vCNHr+Gbwiynbrg6Y0oLhxlyQB/iz4PzxBdchnLaMEyLr
7hK0Rj0ixJMO3a8IhLwhyM3PAwrKFUen/+OL99iCYjsSWx3OvKBs3SZ1G2nWsaWs1Gyn72d0agst
iB2oxFpeyO4oU7LA6B26DHkDpzdHHQwhkeaNg9paG3Ci4NUrLNT1n8ZZEU82dtNx0Luo2dhkUaBs
Fk2DKSYc23vfbP1HMiSUOwe7d5R0QlXIMwRET3D059vDsBlnEeoOo3gZFc++0v5D38ne0kK9f5wx
ARFVg/KHxKqOukf8uR5HPK/ICdCDKeynvh57aQZQoSGJdJeygeaxX/YfPp282TmJrqMTOdm32fwn
mvlkkgRg3nSzsHour6hZaxf6aUX2B18qtGz4ac9ThqNbbrGG/Qjp630XwNkBlU2CielxkXgCThWM
9ZupygV4v0Ieozlr2GmSgHSm7be1E/HVPjnkaQ0+66WK9a5T1WjIAuhVGfAMjtCcBvce4EeKbyhJ
5YeoSF5pR04ZGBnX7N/JXuXsEt4lub94mwpYXlS9WpW7qaYLbg2+X1cpLx149c1hqqIBO8U3bR2K
Vxhbmfk4tboPaRJC1Ev1+oUVLPs6FHlU9ZIjjoTlBRZ5coJGQSQucB7MAHCpBTThw4Ax1gdwdGDh
4XFsuKmkSbudnEgkJbbH4wvHk/CxLcw/A/UwgB+n5nFnrFpCEFoas2Yki18b2ml+Fp+OqmfWlxtO
29L1u84IITd4TXJq9p2NGCpHfBUoL5bdm7FJF+yV8uctHVaL56fDP8n6d+7Nf+59uJDyvHC87EAd
90qwdBAbDFHlpd1cXLI+9aNo9IvM7T+vEzmJuNpXu5FPdEjgp2xx+4CmHTjoG/AUMpIyG8YFxyID
Rybni8rkZKCAexGuvo4JD/dbGNCPqa6zdf0d3TNa73K58k+hihzFBgJ0UUgt9wlBMBUbXss2d2XZ
ugX8t38S7XbfmhbYlRozwelzITO2KrjsZiMdc5oWGWebclKk81inom5FQhi3QeYRgXfA2xYWT/XK
dyirYigOWhIMKvI2filV6r+OKSvZWMMdS0QJ4xbqW2vf8owFLUg/gyfdlq0Gjq8eNCm43/jfIevV
bdXPli6DmJZPyjHIzGp3YzR77NAUVWNbn12HmfNVzUTASysxjQnqfGMzmaZQkc6n0xmifjgUziUB
94FRRm7N85iFsMik2cUJf2KAUeRH3yfs2FoQIiOVkg5MZNruA2pvhWZ2wo+Q/A4neQSf+FWjiEvl
7zVvKsOmUTziKwB/vWmxDdQHI2qrLN2s3o05XcqRgyO8lxZyoEWVAAOrR7JQHxaONUVeOxgd6Wit
R0aiizl6DeqKJ0NGZYH1nO/xsXKjh1FoPhI2FuTHQCA4qDXKNDDL+ecBJyAUfSVxn0LiF9JdzCQU
qI/Gkdcce+mxsF1w5qwnvRTY+4ks+RCCWt2Wmm0np1TWsdKr1DXtz6exU3i0IqmOq9j5/i0SKKxT
DUkxHDaxQmJXRs2QFguLm+0zUyZcyxhtBlZ6peTYNv9c8lGgptg+sIvHEGf1rQeZH567ovsQTF5f
/yRbiYuef+YsSr9Dcmg7yrarb+mccmb7XOBWcgBN3RxfVzJgDvKHpP9qQ5J5d3C/0coHA1vsqw4n
RsHO8kLqWgeqD6/TLbfG6cNIS/19Sn+2PbIX31nB404rzncz1jIUF1PMUIgOFSfVg+A60maytefR
bLD3Ap62mPu9vwgQFP81xZzRV+tgLJHWqANBBNUAXIZVplatPVO8Yh9hNngilLlfhzMigvuZuwDX
V27jtnvbF0qeiEZeSNPSeb/peylTsnfuOUccjxjwmRF/e8NU9IfJYKWPJRhQkqiHfJxHM/pSoywR
48GAix9FAI8krIPaFoPinelj2zYwPcNT9OcekxIhAvYjfB8CZq9z8Qp3XUBkgFVYcTVPTP8XrW49
510cY655oc79JF+3vXfXRRhBDzgR8qGC3zP/dTGgHKd2PDaLih+nfwyv36orXZ773EKKZAg6tq3j
jIjVp9b9aGsmxjKN9Xr+JrlAPrJtYRgHAUIjg3Gfkb+PlEyRA9CJ0qrcEmquj9V3E7TAaXYxUGW6
Yl/5ahPxPuIhpuJp2bHxw6qA7dcYXr+OmvjW6hIg6nvsvoYawOhJG8h/+mYMRfaeI3v1aP54jxn8
aABx+kvGogtpgTWSBimglv0h3sxO7fBoKh3SfeeErvrTf2uzuWFBYgApmyCJARp51H0SNfnz/YXg
ZDo0CRBk2nqQYGNM9XrZ1Ju3m1DqvtA+SBkxGdDkcdtXju6HP39B17uuFV7bkdFeX6rNpLpLo2+w
ydYAirxfA936s10PLs4QWd7x5wuyK7gBGGWuDfMHaXADTK7Y7Q5X17Cte/iiG7Ky2mK+nqCRtRzP
rouK3BBf5DuKqF0NnNU4Wrj1lrpLQP4TkeP/vhxGw0ZY8sB5uwd43iVf2k9sjTHo9GilGhxTz5HU
AC0nAnC4YYOAaFJubsmXGQKqjqpCsnUR4Zf3HVmuEUaSvizm78p/zEkpeGAoggZmcehB1X9rg9DL
Bp6uAoi4BZdXBqd6eb3910CSQSIC1efYjxe7U/IA7YJ9qhKRf599Fp0wwvkElnKVuZq27TJrFGxT
L74LDS1CYYPo9fTQOXpNRhbOpM/RCdfcVBmMo7S3pdX2d1RGtXAQH9uTlt619THsZxl7yxq059LG
wJjLiFJIJ9Z8NfYECRDjJpdPxI0yWuXZKtdgdcpGY0xlEdjENbEFZrtWC4eXXv9x0RK2G2+z7P2w
MNe5nYFfsZM/EnXW35U8M3n4ZYF9MPB75rI8Pq83a0JRBHvfH/Jr/eU0L3NnBFeEuaVO17JW/o/d
L2TmOxnTUyl2ntJfGJ+aD22rdOKE0JIgeM2O0Y3n6KXnFO/7+4DcBP1A2cMwb2MWQ72WXQptWrLn
95lDXi+91ymH1qbR37HJV3jHLwRTK5Z8z1M6CxfC7TN8/X71c9596I7PiIirbMtT8k6jVSFswYc1
cOL6RaNxqVL3TMEjLBejacfmN3IXlt0C5rqKRHM5CvDeezfvzNtRlG6MO/vXqVdGkNCr9e6JAnXv
nEoWo1uovhbYD32jp1BYtf0q28JY2xs2J/tdkg4aEk7+jb2MPyWQy7AmRmGDm01DfkDMjhrcUGsz
i+04bnCcEg+pcRVdfDXdVoOcWcx3rzY4PVut55eyAbQ3tAFWl7PegmPhzcKqxo6pV5tr3TvNlFT0
qKC6M4mrgu9jbUwWnElSd7qn9dCAMakCA7pY7Ek91BLJEDJSye5t4pTSclm93kRPvGnNmoaW6Ra7
kHPznM+F9BbfqqkdfSXzKJfTSQjvUfIoP9GG/fmVMkblJsCKvnLkGYIFFELIVPLqYoo5k6jArKvw
g+27dDjJEpQ8G1i/+hCLd2nY/iPf+TdWF6ZDLMh3PPX2wF1fs2wZCigfVmNiVsh8bj+CotBFn+XQ
iPDEuM79kP3va5eLKxUu2LRanliF0F66mOoYpf5acKaMf1bGu3noqb5c/nx9TBP4eyQb6eTaZYJC
4ivQ1PrtyZz5O0Nj8MLlbDwJdSXS5c8hickAFeKS0LNBtInHub6gifaWicIQ+vzsXBWp4dKivwAr
ChFa5HNSXrpTqJaT/P7O3RSa15st4Axdr1npeGDhp8t7YIhZLCfnYHbQvMrY1FcHUb/IE2q/mW44
euhBSXeVLuyoKEdJBQLJoFDvYa/TtoWvoUzQrC7O4eIpoeu5/cHj072KBqitWkQCAhzwlQI9JiNq
cUPDuw+CvrZfqrnztPfTwaNt8Exinkob+Emc+uL4JO/n7Kmfvfyz8GU9Es6UenoDJ7h5XPdcCHBS
4hXWhFqp9/J3+GO0t5GfrdtvGKwBzUYuxQ/j02HaM2ehWBFN6JYPNM9Oduw08Vavw0+RqepPE0Nb
sKs9VMjjiagflzMRhoESF7/3a0LUXrLIN+vFOnTHTq1SNTj9J4MT4PFrKV+2q7jieWt3EB1DXPIZ
Js7J3/JoKp9igl59iF3gAj9BTV9oAsZudNfEBDiXfZ5z7/7V5kKoQ5jCZEoVna9rv/HHL8hSVoTd
QtT4ehQm4lQCXnaSOo0vIv8mRBXMmrftl12Bm3BwKS84MypoeC1rp1keJiLvzGS70Ay24zDeifMc
S05RHcgqpm3qazyGN5CdSxOQtgbrd45GCm378EpOM5CpcOugXFQjZZfhF5ZT3eMlP3mqH/Uvxahj
XQSMp1w5kZ3hOKhDAtmidM1cqJnAA24Jm7QfKWG1mKnzLNbrMVRyiQI3WLzRiM0+PA2/fgN162VO
n7+uSfNHvYOxksnSiyA54i9pHNZ7VVni1/mWPtgKeA5FIpxYZM8kUGU8F1QWW678AuwOO9Sxa9rg
m85D2EZ/bl2kpXjQqcLrsKwW8XUN/4E2EOD8sf9wtaK8LFUbSQEEwrEph4rWXmuWCD7Eal/W1nxt
NbzZ7ol8fN7vKAemAFglllfHzuSdQnVwq75RhdhEiVouYvsh94AATQL3ZLqKRc8XzuiS2ZRLpmEy
Yxjo/ySu4zCIoiFUGI4TQWg8JWEGSu5lXn0oqlQkw5WDL+dqoJK258qo6RXgrCFdZLSV4gdom4E/
7+bgFN2Gr60sCMIm4jJx/sN0BybOFWig64w7XHv2F88fLZWyhsxQpzvSPP5kUFEIFte0Ger07Z3a
fnSY98AKC3Nj5ph8raaqBXDdZG/0ThkDvsl0Qh2yMReTEiDjTOv/ZMq9bx7YVy0M13rl+YslgMu7
KVTnNc51KnQcHQBd7jApHV5PjFC1N2F/r/qZpokSiA2QGpo4cWtxx86vBhUQ3Lnr56sOcE/u4JNl
02vGKv5Zp41OctamQYmiOP0ZcHkOrv9GkyU6Cue+uMbpiwLkq7H2X1qD+VoLz8GNPKAw21FtIfI/
9QH8wyTg2fMfB2TpNdNcu8F97a+mQPPP1bwJHazxTeyt69fcXIbIi2LycVEfElFmfnTQ8+yh26HN
MbhcQ1Whrbmq3vYa7vBYLb/m9RhIbUvgPTSsnOZfIlc1ssVhOOXJZhSR/YWSfcq5Vw5jPjr6kBqv
6jj/EijzXWHAXnH8uKV43tJCPbySaA0u07qY8Vd7Wh/Tv7m31dOWw1s6zxZQ6ZlsqmxIUnK2af46
0E2WDXFnLpVtnwKDYgbO5gfAlE3G/YzX0lJ/7vlYiMu5hS43rkxJcbc+bR2KC9qj4mz6XtUgL3mQ
Id7TTBHDkbS4vCIFCeQa2HEGy9piapetUBW0vZRwd2ILt+WgW1iyTZ4q5f9SjZ17vCPVYFLa9pWB
zggWBqFKTVxX4T5cEDsw8sTmcT8DMUM9E8VKce61Lx5anQyCU9jfIsYPY325CR+t+iibKndbA2mn
VxLi62YcGBv9tUiZ/ukvhTm+sQ8Bck4UUEAqGtJZnmhdaDNCCBFZfqjlefgooI0h8TnyzXphvwnM
ZGyxVXmvc5fn/7zK8Yt2D3HoirPYce+f1WrjXDSbNuG4+U5NgmDuInc2zmE4MlPghFuKQjZTueQW
fqg93MjyRHXHX/oSdJmCJn0UnZL2u9lyXqoCBbDNnaekYXuPeV447n09YUIwz5pMD2RZ/AVUDD/T
RqbN54RfhXN83uGvPcMb7FM4olI2IG667obERL/QlA2o8BFhbuyWZT5WaxWkkt2LnA+PwQ0NsrNh
a49e57s+w2Xjj+SF9JOcSJ1PFkPHnQHpKXJZFjY9D8m3mmiv8Px7BHIWmA0PUWjob4P6nbltt7MV
If2fq4F9MR0i0TkRRmtXRgbDipG6yRzNE/cpnDS+EsvMk88cyIdCjGimmMHK2yTkOiMbQmipDvkI
j1px+QqrvdYttGReSDm1IJpul8XYK8mVP8o6GVglraaLGRk2G2Jv3Cc5dfTQXTJcw+1exRocG8jx
MpndolPB79ASZJLfXTaLv/ayGIbfB2Wgv3S96XHZd+S60fb2gu4Odk07OuH0oC+Ptq5mRQzpn68k
2QvehZclF14I3qZID9qkBIidaB9i4MRIY0+/fdtkChP9zNEo0wi0CPw6cEjdnGxY7X1QtfaoK+7f
epx/BisH+llRyIDuyrCVy14RCLqcl1BrVBZG62HqlLQeTlsPfdQDj+W1HPRl+lgrUkeQhJrJfzS0
XE1VFUsnLSmeGE4GDUYGT6ljsykhqpOHnx/JFsKxfTsAHVui5sh2KZbGORFCcy6e9FvmmUv1oT4E
EGZUKHRBJCAe/zKrMt2AZw9tPf00KZoRjhrE/v5yUjjRQBXKJWMItskVEA==
`protect end_protected

