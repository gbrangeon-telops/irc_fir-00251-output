

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Qn7IteVsnZ/mdHCLR8tB/KgmTn8ijcYuBtDLGh2oUVKuF3qoFWhv7eC1IOCXLirwb60qousghfg7
0xqsSbRyrA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
VgzxfdCZunpPyUwqbYGeC3ulpMsK7w2LNEgFOrFKGlFGTp9v30dyUA7MsiKFgCrzzKT+VrIPwMvw
QxU3GQIE0b38WJ5xx5bDenrFuj9fMfRnJLJFcG2V0iBV/hYdVoEecQkZyqCPVfkUdjfKW2nQQ9vE
YSgHM9qDx8fLqyQ6zAA=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
1ig4g7vOmzvtScDRtVb+tZEnSyg+feSk/Z8usEB/u9AljT40pDkFhR2JxLDYn3XXgfKo9dhNCFm0
whMJYjKNylxxgSFkNtQwR2XIg0BWg/XJdnzmvhE+MtmxAUvbHjuEhgVFiobIjRufLvFlBirtf174
Rb6IlMY8DFzGP8TNtNYlVuQtzXS4NvjPSDwmxdLLBUryIvh8XgTaS4XKcRx4c9SU8usSs2eZmKp1
PQzsFR6KYhbJsoU+KNdgC0qr7WxKSf9E11HFfNp3O241b9T36xgfVJMNzGcu/ZHXpRemcPttjJFK
GMln0o/DwR0gidlS+JLK6pgrPDgP5/6nmLlP6Q==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
yE7rDdP/qWpLchJqOpJirpc1zOl8T978Yfk6G9kBcFGYD0r+ZC5agvccz99iMwduJEgIxwFmjnzG
7g7dI8mK6Rjj6eLbQ31Mhsmq+p5Y7KQTNM1pfCzFCw+oJzuBbgsBggo35NClB7Hfb8DM7OriNRWJ
U8K86UkzA2Prba4TIBs=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
BN9F+vWJYtgfrzbWbiAE08ecWOdWyzeeA+i0U6sGshkhExwtl0R/3hfy5ttqQZECat07SJZlP3jh
V4CCuSQw513kvIfiNR1n8KZK1ODiyg59gOwmz19wCVgWfDfnfDXmgYxf+0derYmc4F2n9+pXRhDQ
enznNCCvV1TM+SbAXbMWWC77ZJDkWposT7aeuix0KzNLkoMsiFOvzPJVJxWsxkGPtD/xLXraVjuo
/R9zbJjLpYz0T/O/R4G6FwuMiIZFlEBmhA8YI04Xnb8Of0h/udsHa/BIz80Zs9KgMYw1jOPT6P6u
7aYcNrAi7eu92a51ZSDtMllbDqQBzVGgrUZg9A==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 15376)
`protect data_block
+19ksAR+wVLBwT1T53h5WO7h1C4GG4hblNbK6IHuRp2IxS6iX24eNLloHA1LJ2ekvb0mvbuuQtbN
C5SRtGRfCZKhgAA0Kdae3tX2eemiSOH4hpW9eaT0CEciNavGADQIE3xnns2qFVoa2sAOhPC6Ess1
vuuZBWJPD1T6iwb93LM5fnQkm8iZiEy+MvKOuw5qfjkIGJw6hY4zwziZPXCJb/81bgKJp403x9gO
NfXExAHnRUPPrlb0saxKwtWIaNQAoaUQx0EAZULiG9xQSKZILCziHY1rmH9N1M16F6vkKc7e7Pjb
iiGkEt8slM7Ykm3QCeGuanH+K/IHyjHc16k6yexdn1bVTLTAY4IoY1+nKKawh7zUnxHh9//qh7aa
ukaLga/YpqPtlwAHvgFWo0orZZa2aOk14KmCdfuYkpXSl06EiDe5JFiIIq2c3xCMzv6Qpn7Bf33q
JZWYdRyA+Ilv830bORZHtCJo7APZnoQplx0bW4pFKhjeKgOqYka5SzBPbPJuTsLBJqqctIbppFqY
gV7eOD+pDctNjpQaV7USKWFjD76qIh7SOqajE83eli+BX9YuCIAKNZRuqKK4YkUN+1dZ4M3tljf0
LYPminNUkiGJIK8MdimIHbQzP3XuFR3vkufKjg+HrQGoHNaZoeM5I5qDP63M/sJK/1aru0041dTf
WujXG4W5fhB63KKi+kl90jecjsPRMPHZnlkhWRS7cEr+cHT2cWi9O2e6WB5oP0QjPNcVMJXLNmbR
Ouwg1m61L9aj0zei/Ew4YX0hqY77oONF9pN/ptdQmEdmplABYAJGXOfF2dJTRZ0O6yYq5CYFc8u4
85PPO7DIIKbaFy4z2DfR7+5KU4+sHG3gI+GBUMNeTELkFMFbK3/OuhS0xPo4xI83cGc8K9gwQSrt
yw9OeiHMyMdl5PhVDYJ5EXqZHBWRgY7KfF1UOSG62NpKZ1hhMk04t0wMWrF/vXL/C5Fx83MGn3W6
4t+piMWjCYPrGXoB3rQMtQrG1NFJP30M5DiYwqdEGG/ucXghGSJZP3lvs9gQuzXlXTMA5Ahc5Veu
YYzVcFOpWIE0uDXQ/t3Ec6X3yiQTeMiwUD5DjxKg3cGkotzfnWZ20y6JS80Y5E/ptf7c2E0Jjhtb
tkicjJ8Stnt4r9FaNnLo1byOckXV0glqpCdYi45QuEd1hhYXIiDXL/0+7/KJzEpgGhbl5lohWMB9
EZjGtu+5sUkblzfeyuVoX71++kj+NuUcX71234HEwZMA/7b8l6Y9H5fMLwxaK9ZHEkeiAMJACA5U
s4yvot8kMsspH+pukPu4xMfJugy3LCpUW7RgGxTFGSJkoRZEF3dHWj40YhGZy1kZROseLgTZrLm1
7RTPv+vL+/z7BZO5jpX7ZWrvtZSd2Lv2qxdl82EMSdEkXyIKikq4yMRzfDPaXATUBsRyxFns4f06
H+5SIirAsKKfWVzKFv+gGaYdn/WlCYQ6YX8L7bFfzeGFgbO+oVbhmpv2S0IDpVHcqqbrD9P8e1Xa
vdiI6wdD2MmIPjCjJ2Rihohe/ndyxAveSyaZCP1Z51udJr0uvRbipdFB8aLuvv00Tb40/p/4g8Ot
Q+TRBXOvNcyUYwf8Pi7N+BOE5M1vE7+GZ7CuW47n3JNpxdw3Z65DC1nFbyK7Bal+7E7sshjjfN4l
dt88bBP+udTQmra64SW50pWCdfuBXZkOy2Hz37ceIx6OAdrXoFs2OuZhX0xlfWGJOC9v4cJDXcpU
NwBMhq8CFYbDRdXuAxYPCGFBszn/pNNgjjWvK2WYatunUBFiZi8QAWHSiTCmbvIoJaBKGKbMvMuy
2tJMD6a7PbHJDDQZr1uWxJO7NcnlDj9CdML3MEdhBo26uiwcPCzVjJcrCwgBY53zzrpiYq6jplBR
vTDHxNPPhPea9x52PSSGhBuYXQ88l18zE6M07hZqSQT/rS6VfmDEqYw5WX4e/iGiK1QpxnDo0G26
re4J+xpmL2TLpO1pOrK9dJEycIbJL0qXeja3BwyvyGioWKu5+vlkqbmplTVKDyhb5ANGstFjQcsL
nmtjN2X5tIKxKWwb5pywrElFk+g5L/fYOFA0cSAY/ZSgx5ck6dbjxzEGguq+/pY4hWwn0ii64ead
EDn5fKlGr/PePTB6hg/Sj+4QV8j0hUpWeLwVzxr0DZR+CTUXOw74SK2fIsZr14Luu5q6aWcbwIE0
jHnx8M7jLzCgE0ZcrKO1Wz2P5lO1eE19Q2JySI/uRYaZyYxHONM4H6wBxnp4l39Zbrumu5GccHJy
FE1oBO9t3KxBbc6rkTBJq8L4zdgKxa/Po6ooFWrjMNlb+bp+eJmTb2ywkO9fynrNii3Gn7Rxavz8
zjp0divcSv+0od2riYv5PiXnSR9ZlOyoGbzARgsZbM/9bwj6o+yKKxkqfDarpudZRGY76Y3kWPEj
V5llLEmFPaNqUI38IwqFtUYnTbfwx69n776B5aQFXDvpGaAeYa/kQhGKnuGvjnc6KqMxDZiC7AHr
becUexooy3j7qnwRV3lnufdo1vNtOhxQdKFxWO4+xRI3pkw1juYR4OeD+AzW86TyM1jvopjKfglp
49MnrlIk2q1vI8dwLQL35hw6xek8B0/jgt7P+jGW04YzfeitlryNvJb1Eud6wAfTC1rXrmaAdDa5
j3Upxo+MQoa/5GuRxK8gPkdQ9KpzKYvZfA48InVsyOsoYbldtF00kEQCC/YZ1LCPZ2WHOjovy1p6
Y+6Jr5zJSoKDHD5ED5j6crm4DlpkBPB05YrVjDTCMEMi/Hyx3h2BuqlEf0NAPP0RCONiOQrs7rM3
kibFJn0dLBplF5lrpEGhXxEixtJpFDhxSVqrEO1oZllMUADs7p+Tqr+TaUIH7HLJ32IReozTzdtY
kod3EoHgUEcVjFGOw0wQ4UP51Ox/B0VWWuo+JfR8k9maqaICEhnXTS6WLA9ZqdV0RqqoVlNIJF2n
CBi03K+EB1keAZNK8O8wsTDCSXieXCbmeHYFoibr7CnTRKXUJAeiqfqnqfzQy6Fe4u/MimMDzCBm
ObFrte2wO9SGODO8dop+ra1rtZNxyuSjX/Yl5ts/446DCTX2F8+RxJoPIhpI5J6I1T3RiSUtNq7T
KREIgadAsusT+LHIP60WvSnlxIpZYW2W38rGTuNNCDz4X0Lm95m+2XkJsMRUxDz4PhTQkczKS1Ha
hDjy54lfSkHmvdnUVBNRTYWG3z2CMcClCdU4ip6+RdkwRHNtI0O8UKGhwOJI9ShC6QIkqhyJRksJ
5mP26YoPMjEB1zGvHFxbmLIBtQGZki8affcGSZohwgGFw/bLQZlV5ebDNCDvCSu3L/zVgr17arf5
+W7EZzz8J+f2QEPzOrscgwU3kDaLN25zzlfyh7D25zauzEfR3Hiq1PEX0zMc6i0B/ozpImt6uzWg
ALO76L4zVURJzW88vwSFV4xq7+w8mq8LJ2FnvYPEjQtX2AAhm0ZBV2NQQcWza41RcdKbG8IT1IWd
KA0yR4rjUbiW0Lj3jrLZL+193d18BYFph2gNTMBtKDWyWR5/mAsLE9LHE/cBzpEgGXhyoTyPhKY8
mBpmIjl+MRpa/23jC7aLySPzmJVbt4SChvICez9IDBSKWblsNo+fJd/4OU1xPiIWGO+I7/xIFPfn
yYG5a7J23zztnmAffgkpLqovJvnPdrcbVRv4hI/uQ8HeEAieQGBmDzSNBcV/PzJrlAL360Vtj40j
t/44lbUE66n+kb6cN63opIpy1T/1oPmXmu+LgTUUWvKwpurasET2YqIXt4neZGLTljBlRyKIdUud
RqHyiZJECE9nYfdQdSBzVRZJW3Eb5V8x2aIhCRbvmGibmkTcai+xpveViVXAgu0Pkx3Sm/n+PzTs
MJJCfSiaK/h/N9Fqyaq7Tlga1LJ/tTd5Tst829SpX5DIvuxoFxh04Aq76wKR/dUv09A9d6sFC35c
nruyHkVLOOW/Hn68AAVTqDy3y5U70hiPLMWgO8qswoyF/2uGMhS8il5H9yTONvqRLt3dskF7B+fq
K+8SLW41bRnGxFBGW4lzRInV41EyIy38oyeZj2M//Y8pZbhsEqMw04bFXD+2LMYryvHJmZzHW2in
xJFOBkpVLEoEsgD2ZTXNQ1d9KVX8VilZrkJAzlav9056KJeG+hirX3RfJpri3gcfIdQ638wcTS67
+Lexnuiq4+7zQA8P4SoURezoAa/O42zcc5pO+qjzOIZd0/ngt2xp4n1FqCTE1lNO1XLQWq4rWJs7
ISzXEfYrylTy3dTsX5zzXMkXgsyqxa2p9EeDrFNb0swwQdDSCPpmXglKxm79U0UfPeuzCbUMPKPj
hf2BdaEpOIYcKAJF1I7LA0rjPHW2sEshF4HF6yhEmPmwKzFJrmKa+rHJjdg1AJObhA3z90mJzI7b
TAuCvBrhNXJ4T+A9ChV+wauMxaXaLPg2yS+b701FD7r0Uu3yX9M75XC6DFR70NrbmOTVfV4GZrZE
TViztEpRvGHfc1/XnsC2/Zs4QcPzqle5fNW8gzzFq2jruIMM/LOf36/US0oHgADjY/2GKynEWHyB
PT3d9QqudwgKqH3r8hF2IB3Nujzt5pTTArNUoyWNkjW5w1kAcc3kU2pTnTg0P1o1Mja5EDBRpqvt
dVuR8H63Vft3bW5FxSKlbXDq+8v1EF8IXzWIAN0YUCgM2mg7ZEFo7/7sgzxVCq+jKy+cMk9y8JxP
DLs3MH0/C7OCHhAwfDv2o510tQk7AiA4SKQk5CT/w/Bk3v7cK2WcHqye9ayjRWw4FRPmYceBYE+o
kKL/KdCXxloMMClHGSNdlsvcylwb2NWZ0YBvWexqCg+q/Ol6k6jnyNxLyhopvNqgjOnVEBopAkwm
DCoYG2uZpAtgFQ3Vc5WhRknc3LedDhxI7XHVQ8Oncc4nIGgCC55s3XnsmsCUvMeRbmS/2Eipj2o5
2oF/ZlFZGDJtK2H6k+osK7Gfqr18wG6TJYkBBTH1vh8o41qxwBZIzFym7tNDF9+5W7JD6YakV4dq
jOGIXqGWbGxS6VzDBp6CKYi5XFVCdOLmoIbLJ9tV9BegpPwUmXu8/loYpSckD0LF2a2qpCt6w2FJ
TJ+JD2tGyTwlVKMtlZtyfd9ATbVRZdN5+UAqe/CtXsP2JE6Dn15/uBakV7wJ5z85nXw/XWR3Kftp
s6IxElxYOohRx8faJgAf55LI+KfywFQUyW4DOqPUYMs1/xPSR0iTOnNwbf/czverjDDtwQiBoAYD
Klpd6Ua1pKk6p+CKTFQEIvF2JuXX2JdCR9uk6CrPntivK67AOj2YGpoBIRqpGTJ0W3I4K9TXJuDR
CD5gQRknbc1V2CFC+GG1P+xBVSWKls9ZuQ/KUwsNKq5knw3wJCovjmWZUq3+7J5UQNOZeZCnYT7H
Ij5lIn6ObVNKf772LvV4MgxB05FEIyaFM5opf/j9kL5Nd3QYHLa1zYwf108dkEwbt9teIj+j8VTO
gKn/N04WGOlrUuAq7fPSVTTsLVEh3m8HbYNFv/jEZWbq2gyYhnteCtRvUqW1kNeeGUQb6C0I+CSD
PlUkM0VGGCoRKQQugMPb/hI3B5dpPtRqCFbjHy6TleHiZXnAXkWVBf+qkAHa8g5qZ39zwVLLjCK3
UEog6cK3A8Ps4XHVzUR4K4sNh5qMJpPK1PMYbp8kPG/QZjuHvpBFcf8WxO2vq0+GKRMUBUvcdEad
En6wIo125ehkgY3MMwwR2MGD5+rI5fppeGeY05VQpdUBhObLRphcMOg0DTJnxD+OcGetfiYbRoJD
oDKRKZWypws7ZMaW0/WH22cqfwlXioUnwvFYeULG9pGfZUTrqlTVVLvLCD58QcmQ7VPgqMmPg2aA
mD1fYY23Tw992dIEDut/OFcQtb/oXPs8EnpgdxkTwIYUqfNiK31OqIzjXaolme7NkW83z6qa1R9t
vExUI6cME7XKrxlbY5czHomcQfPvYXCL2h6p34hyqUoKIRhZF4HqHo253/zXxnYIRnte6Vy+Y/AJ
y00EUVV/yKLcpjXKytMhi7LPkHGu92SpoS6tOiBM4RgVdkD1cj0hgI3dFHxJIlUh7p4nvQHExC+0
THnjnAxU3N3LVq5JsZPdClZ1nrI3m2UbOTSN2GnGNBJVY5FqHPKzV9zZ9v54mNmGKEs8B9yNuO70
vC/5ou+saWXHEMv2bHSJ9Q/wm4FJdsdW+ZIikbtDClnEi0gKgus9jIfo2c20CcQj5h+DsJWg8lNK
16cfYQ99Xy/MlsOfgejXzxTqA0OmWELBRiE/GS/tGJ1ZO0nl5k+zqoHGbxwkYZWJ+wmkeYDctCO1
OMY35tU6iHCCn1YLErHk1nce888vK/OiX+vdYuorpKiiOdm8C5Z3qbgmw9Twol97V7fyZZsB+A5p
+CTz3dApb0lofzo7kC4ko48Wzh6MzsDx1tYu0AM7u9A+FXzh5hriGqXPK2+XZVBzkqE/CSG7hNvN
djJc3azwDmCMTU1Cjrj5+qph69Eyq8+anxGpAvG99Zquml2eoW5e24CdMyjwo3Oq1nQJCX1Oje59
4/cqkUOAKJgewYAjQWh918n7B7gDyxXBB1DO5xX7RIkGQIpYeY1Rh4sTPN0ABj1L7hLaZzFwUkbK
/mVdg4rgzZ5nKgqCxkGoE/P63mbHcnHF9MJLBEmKXBLO/aBfLm0rp24gExo5IIGYm+VOde7+6JfG
bSzLHOOmNQkO6oxYcMNNmScJ17PcLq3XVfijoQhwuBSYB8CChaxYl4CcbIPcpDBZjJtxDLpOLFUN
p9RE3BBkDJzB0uQreRlySMAIqAwPl8paiVx0WUNn/57JJazY9exhCsyBVdrsYHPCaXo0/2g4WGm1
th1X3YDYxsb+/LhVV8Fuvl8a047VkTH/naIbY/ZdsiMIy3myeDqG8w2cDJKh+YzH2G8ADOCoC6Gy
sNtkjoi0eeeThSLyGmTEskel5fqxT5fyxG7j8IsK8AbdsVWZ9tH+/9mFpZFHliDggFzfKens0Pts
S4rgfy9B/Nnn+kK6Fh1zsP7Ru+ergy7i+HWXs602eTCWpj/mfBYcssk0tjbMJT2tR7k3IL86A8/J
9am9tPGqPYxTEbdecBPZ0y7Z1NIUGOdCGwkpwR+3TuM+5h4UaVKZVasHQagA/nOy6nFItEBjQwto
JanAMjuaYJmugJa6OL4mVUChqUInwq3vkCAJXyAE6WGU4DEGVirfbKZhc8zEEn4TcoJIth+Jl7jB
m5NrpavDM2iIG5US616BUXB249tWTLu+D344DDdvgdNnF8A7Y7XUIP4yqEL/UGX5M8y0XIAAsg5R
21GjrtaA3RWyjh+cOXh/O+rOKtKgcX8TzcW/yzYcZiuFa1l0t+1XkhstDaISbs+nOZYadHsynBOO
VbOrOYkAPb4/XUnH+ewfvrQp4up6ZRTItlfV9Y3gQeinGIgHNu3Pw/VCRxIN7dEqwh9E1Zis0Kf4
PCSkPWXNZ3BiYFQXvVd14apIa13+Gx+0+crNNUX+u4UKa5mmN5V2ttke/NT80VazmhyKA3HiB2QS
MUg6MJAJ6vrqol1rwqwxroIp7bA/7jwbHFbIDZsgXoZeeZWR8cnHrJ15hHqqFkcEM3soF7zwoqSQ
Da0cyYVHMCP2QSE6CFcjUFSoy0rakrlPP+/oWHPKp55M1BYcnZ9IwiDG6Br0ZeQJqNPwZA2zdkRL
hqXmaJ8qH8BIP3R+c3BD+TJim4V6v9dX0II5mAWZzbFxvH6pFoYZbOtJ9fxdld7zsfOcORIp7h4T
x/yIedZWNKQvoU7wOf9LB3nTldj/NZ1rUhGjn/n8+CaJLnPzW0KwQx9RQXOk3xpU65TZx33/O0W9
aDzR7g1keEFdqE52fAgf0qtVNNuiDqBK3Pk7I1z3VZkZuzmwa2Xp+whh69NhSvPg8vvBEnHxvN32
WnjX7lQMF89Th9s9I893KhTO8jTD6tGF6lDO8DKlQRs4zNYFBJXcKtIVImLgUjeCZZcMzXfrG0R0
t5txKL5G2+Qi3blAUOJMctnprp9seY+VX/mWG93t0VB8d0TPFOkQVHpgenOTeHLCGg9fhbACHvrz
yn3htN4W4077TB9XcqqF9LFmeb86zu87D5ga8AqgAUAsKWdZGvOgPAVt1qF/KStxSg9i3eZldqDA
V8z2y41WrhWkL3ypW6FyAry9LiYY292q/z946E6aQd/9osgoGdytMvi121+Dpahe6yhobtk2Il9H
xMJvteo2PyWB8caPV+Z4+DpbY1cSRfTSlU3kNVtXmgiXcHW2hz4qa54RBytFU6XKw09Kx1jpfsZM
4Q0lorVqx5+vK6iLHGh3trGm2eBWu8izyerI6uiR/SVXLx9CA+P/OP/wCucJhLJbezwe5K4bR8x2
emZ8HeXaUldZPO4Y5uBEv2RFU94jZyBQCLrPFR/wRDUQ8NcQQINNoJHoUK1G/lBMOtu094xqqCAG
zruA/RbIU9HkgJVLHhVv/NfxYwCJxUzNgP/0smdQOZ6ZRky1/mwuf9L5iO9ie+UF9uWJEPQjGsxh
eqs6HvEmnDoJ8mgwkbbj16z3wcGv778HHCt4yr08PCb9M3Ub9+3CgPc4g5N7ljCNrjVGHDLOz8KA
qY3dnEhaIs7FX5uvD5sAAMfQNEJ6YqhR5iPjuUdsn06EXmDb3Iy7bvc1gBuz+N5TDkn+luY4Xc4n
Z6ZJiAPWuJyI6KLZDX4BoSqVUagidSVpWFkpJQpPp/oKp/9nlQTp5BRZc7Dc/QW73vcYx+8eeZw+
VqlqXYM0RKQKolLwaEWbzLDp4+Kzr2NfE9xpvM4oZut5uz1u/vISRbnzukOt2GS9gRrChqDZJgkS
CILyjXausHrwySLpw+tHYlMPV9za6Izw7sIIrRE6ScoEzdceYB0Ipv6fLr9niCgzSS+SoFugRbOp
U6tfqjJbNCiXMEx+N/QgNh2rq2bGvVYsCtQP3Dzl+MGIf/qcwEBZgni3IsWcwFvgPJBmYeIkxBNK
P27KdlkxaN29+Sr+IHxrTPshENFFAtfys9z/SWfVdfpJwQ4Gw+aELSxmIKjSzpfJzYTxIGqVtuoA
xXqMWf9OEHMKXCbx8sJhcAlA8a6kYFU/kHdY32V8PDKUVrrkgMnHavWfDa4w1/mNmkgwpCOj67AR
dz8LsYM5y3O9pVEmGELNP6DSBD0EOav0y8iiktiPSJnDgqJrffG8IFEQelM3XS34vYkLij6L7+y6
bxCgHCc2VIrO5wEJ5v6sD+jBtqgAfnxupD97U7Gr6O3+PDYToEoSI93JYBr65quRJojvCH7oY1j1
Vu1X+bC8UFHzT3nTkshtVtFIgE3b3gJG4nZNS0AZAJzvbG/6L5DBQIB/3ODrV/QEn4WqjQuFR+fc
NNy3cj5xgMpZiWJQylagoWqeIDbY342XECtudlFu9IdNDxsHzLHDLoAp3YVqpg++v9LnakYy/9MP
ZZbJ7VXyj6W4eFJfxm3AefKm9DDWutF7+DIOpRUxzHB5Vz0MP8wx1rgtx+R96uLCvGf4Wlbj6+BC
eadC37cjTmrYqTWAus1H2XiuAyFLY4ipRHo9YCpNIV31y4BLxOagnaMuM7lIHE9GvmrK1ua31YAj
nkkO4Li3fSECOQ0rNqimv91sBB56RsEh4uMRQ6NiNs7Vb2ADhmAYpYX7bgBzVTjBRSyKKlGeMmL+
e5SsNHrThJ3RqDPM0hCjDAjreWgW7w85oSuEPf5CoocOEacBAgqNDZ9MJK2va6UNA4Pj0rYn6d+M
kpw6qrkUJsj8BAhaWZX3yG9B/gcVsuTtS4u+2W8DKIUuNHzVZyEpQ9U/+P3Yb45t1w9JAcKNITgA
D5Mlc0+qJ9JL01mh3lz3YjrH2slegLUPKmiacNv6uMQ2eMa6GcyU1RTRs4QQWdvgK53Sb/QU8rLm
ai77sZKCIJZ78g6BWpq/k96eeaPZKhbIO0D6TTcIhlZzoPcEKikjanc7BFjrErlFrnlleF5flAdZ
iyzQCBVKNXZ2UY3VM6l0KKEVe/EOMaXoLdlA8Qx8wMWF6rYiWumjmsCVub0r79kagfvqazaR8UIv
q38YSHZk9G2LuXllI0CNB29vhIQ2JEiDlaZhkJn6ZlrlQIiMkG0lQoHOI2Rm9DHmsUyHymIPwpwt
FH/LK+O/DqNlUiulhtJxMsckSab6I+taOXLSljiNdSbi9EtXX0eP2Uy+FVrRJrDzWT3TvPckuj+B
af3ldFTwIucPUWJ+uiObDmphPsWi4b4Ms4vi66Ar7taIwEBHJn2GjO7UKXVEtYWM+nckbXtbTUXF
W90x3jssN/HhW0g1YIdX+IEMv/lzGpG6IDkcR1VZ24bsU+realOgArhjqKf6P2i54GqB6VGduQPK
xyzSwP/UIa2eJKKkEihsTqrH7djMqPVvc/futMOxjqc5fzMyeyyGLdeHSkzAGkbLtnPP5wf0QRCT
nc5ZHFC4A8JIpaIZC1ak4C7QBkAXFA5FgA+KhoDB9JHeWWeXIuHZ5eEFpa3bZt+UH3ses2GofB80
4HxpvW/oe+TA2gTCJdxFNLFBLZs7CU1IrNaPYngHAAba7pQBsnCql34onjMu/JHolkqFN9HG98qQ
lRvVwGDP/ZNMCZO3ci2Oe4pUhmx4a31zfzXI1P8fLVrODcHNRMl/NrsNCK7QSX0eGmrad9UYjj8M
LFO/qfvJf8N1gP4WClC0xdlL/Q+jjF11LbuJ5VC7TU3MB40ruve5mK5z0fko7fQU8ie++mfUPT6Y
QpYJ3pfaduNPBniu5/1gdVPowTjq+9w/qMqvPdt9ubDJH36LR9qfx0AgFthZmk45ZiAl/3rS9h0f
8QO8IEekX2+Dk3OZ3pYeUqM0UppXXPWcT02HMfCL/2qNctM/sG+2FaPL1zi2kuqjqKQBV4zeFU//
ZcyjDZ9AVB2klMQt/gwqF9DoIpfCEs14IYVBAYbBl0lnNwVDHoLG7zqh4g2BtdFhFbf3zrz7I5Fx
hNjky7bSeIuP9HH0tMAzkkKCuvJfmZtmZdIqFjiqqnrvPfez7Z51f2OxCusz0L/xitN2zGYSjNHl
IrOpu2dH9m60fJlxmHPdQeUW1W1FuEXNRcK51MpbkiiaLjLpnCsnyBc6NWeBPyIEmtjLwBQ01aY4
Us7eIMDmzwFoGJNx2YADSMmDmpOuwlvOUpkhGOSH6Ia/6k6M72yI3gZeftMhpaZC6UG2egv2TgMc
PgQz4LnMrmsS5GkNX/AqTEXYQf84/Znr2TqZVaw5LmG/MvTASLAb4oaLCdHV4RtWqw1RwrzP4+7J
eK/VYQkiY8oDYBgFCeNuhJVRpbeXLg2G0jH+yLHgN/l6E1+vF0udWQ0hNIR5l/LtuBS+RUZFgZPZ
igfB8CBW1Fz/ojhnH5qmX4OYnkjb8CQR0zsrXt94Y4KxDoMssO9BmJAgED8Znzclnzq8/0rVR0am
Pt3LdXWVIza7eg4FC2Suqyxazjo0yqwpMWlWyxt3MbjWcUu+1a0hyxZdI7W0g9EuLRs7K6UHAO7m
G9Ly479WhdNH1gbBohYoObhy6dnyI3Ooebh1FT/aopedHV0DCYr0llVfiFbIPuuC9eMRAFN24c+u
GEICqNvXLrgkAyUmMlp10MXzHFr1EbGAi2WGS4ARS4667TgHlqTiBM0U4O+wBw/JMwfnykh3W3Sj
ZwnVXY/MGat3efO5hBJl4DwhxQuaUYw54KHRCvJKyQCx24P57Dn0lNkrv/3YEMPOT1xmBRtvNhbG
dqElm1FJNZUZ1PAGT2ajZRGAaVV0YUVoSXJ1v6hwZBAEGGkTHO3t3h1FYvvKeEmp2Hm6qd/DgftE
wA8dpG5aNHeIfkxDgMLoJgrFx0f3/6i5MmJ7tPYoniBpYFNoXDtktP3ztP64gUO6zQibw7Wv3wYF
IKEItGSdxvR8xjG1//oj9X2n7MAl3KTdXtr/R3YsxQQeFQgV9g3tcaJKFcmMvhskCbp5sg80QK9Y
OeTRjbseftv8mf93RrbG13iVBV70pEj6n5XiyrscyqraaQDEljepEQjimRb1DJBixZbTZQj5IGtP
jlEQgJcBbI5Tfr1XkZmqiD1fJG23yks9Yrbg+Awg3v1ya6neeLNpSWwXQAIXTqMnnTD/TwiOdGPD
oN5orcEF0YjM+lCCzw4yryItUfB0ydvABbsJ4+9hwA6Bt/nGmrg4k1TiSwTcuwW1zjw9Ai6K4hbs
xwLbDUu9ZmPuM/TnQeDvDyJNJ1YgBDugViOHrjWOMs6Zu+qKITFTU6OjhRZIxmbcoErzW4514pRT
HhVKD6AwfeckBPvGhto/2O8ayTLgtHaFPhVLFtWJ8AwCrxzPtfcwRTF9tmyiCgfqBaKJSK6KjNGL
LAdsuMilzOeC7cj3m22V/UnZ18GD/Mm6eeMfHzK9yTATx0IuhCjbeSj3ksxNNZfjV6yVHmkgj/tK
wJ2+qSfv6dSOwYTKOmXhcca+mQXj6Vvc8rS8PZi+jx5C+N3MPbedP4+V28HWfK9IcfCi3pRASQ1N
fvTE6HYzESTR2dpYGJFuWQqaU2DuPRVTMSaLhip4HvjbKk9RsJZzgRf9xSvlm8CmuS5ckGsYb3S3
yGir1pTl5G6P5akJP6LEj/KV2W9Kbpd4ywGdEvlfkStBWffyxPSmWK4F1/u5SgoI83En3i8jylJZ
zLnOa1o5Q2S/PXryuFPcC4Y2sCHp0qsGfm9No22dSSUQZR7uumrBkS1ZrjW+avSJKgzSh5TqoSpO
hsGyLFohJWtDKxpNFcUafZ079wB2jceoJH1psPYY1bjuhAFreKpGElwruCURa2QYKaWLkHTeHYuM
eSwRMz+jWzB4uvjqMusAlI1eKk+wklYdOcMOJjptRpguw9JipVCEAHP9uuJCiM3ZrxBXaf6mBa2T
QCM0fd3of74hTTkw8VPpC2GrkYuHFPb8Bqqkp7BL3q/NiXkhPVyqY3w1lg2iL0kEomtrgNXYfTb7
ialjxv9WDOGK7gJfclCA7Ioa5bIhGcsTXIvy0QEPDP/VUTas1Cxb+WEyHbPSVlgnGAj6UapAqBuf
xvf2lxaOBNErGMqGQ5qLcP9X1+7YNvcX74At6Lz2ZYJRu3Khrpp5OGl0OLvzWb/u2v5xnn8MIw1h
b/G6MHvjvFEaqeedscrSeRUIksOvuiFiy5veNXaP+tognvQt+6fJqjS42Fc2cE/e/LMyqox+sZRp
nFk6d2fVbpDJ2VRgeVgeQ1XjGPyV6Ke+PhmPUybn0seJPFrX0cz51CnER1Jly1c1K1OILuvp4Ph+
F93el6iFrMCVtpHX1y6Z8B9efYATZ8iwk4Gt1JRZAxyum0H2f2ktzexFz22CNdRDJDN8rpLDRWGi
zkdEvy6qaj89MmMj7Sr1N+nZfcTlCCKN6eBDQLO6CUyICkud4+Pn1EtObbuoKx7Pfn8W8GsJ6h+p
0yoo+6/YQhwbcOBAqy/Q6gltTHaTtqUbKIodcJ89WYeB/NLwU7xfB6OCJ5zM+x5kCelQR0iOnuZM
aMWOTr7/wQMRyDNQpHyllD9WzWqfmswP/fQZ42NTIjTU8ku0KUPUnm5AQrLyelqKe3Vg0k/tn3yN
cWkbl8z4IqYwy5ivIa1DdxSusQYTWLORqCbMvUrh2lRAa5mc/vg3+eY/YjgyGxyhrhlu937RpfOk
xws8T4+P7BsW2XUDiYXsrTE12LS7l4jFcRUxvW8Yx6qqm4hYLS1Jf09mtR3+TKeJQumiQI+3VDiP
klvwgHctmTvbZ0AVKQkGAU+wEi9UugRAFvlgjEDJYuBYLFrx4mQiqxdCd9pQz0ThVU+XQqY/oadx
mV9IyJOKyJwa3h1QB9GvPCYquXWF4hUx2ZnLPqI7s0+avU3TKCXew5Crdp+WaXiXyAlJXyShndJJ
H+vEy7/L/j+svCmUhiqsRMx7Vb6exRZaq6ELzawgOJRa2SH7KXbuSm1tD+P//m0LC+Ubfqem41oj
1a7JLY4lhYV6wXSkqcp/AKYqckl036dH5+5JZdWpGp+XW0rNVMVitKoCDBIN7s4EbBzk+BsfbuFg
G947K57yc28DX4N0ogixhrC1S7CyhpmxDUjFGeziZdmD4dEHULiiI/Uqrs9/XiI4iYAD3RMY2afy
/6iOZZOw6zRyWxbuifW01e3ecTKBnozEjRiNEJ7gmcbNuIilJStyJ8xclc91CX9Y5QyDgmUt0GaN
YGVJObJtc5U1B139iJRhz0gRfGADnykkxX6RsW1QtL56xJHjBtGQ9nhotvFrA3EqSVB7l2ZtfCvb
QcYWnvwv82yb4R+gx4Uie9TaT1VPyv4tDx+wN6Q5pOeMZsHtukkqLKwfXSDAYTanoDKVjx2mrhaj
bwECYWuVZiAPWc13kkG8lO70H+MSZXbnqTv2v5Wh1wTt6yj2eRfRdBvU7g4KA/s4fhCfhc7xkK+m
hysBY3BBOu2o3xpcfz4RcXo3u8uB1ZqYLcbi1iwru/4t6FxyxfRwqE4Xe4HHqeo76q4CA8q1xjYZ
Ji516QSF3W//sKHoJs/XCsMfjXJ2Ur/hAQ4XgJM9SK7XdDgXQ1/EhfFJjmErQ+ysebCXobZ6pHZu
My3rek79g/LXR0ReloGTQDfifoDlSvi0iKrndRKFk3cjbuETNm7z0KXWUbmrPyzhy4VNmGHo4xeE
bosrBU2fVGSZz/7/yX7jYto2YasGVfuSTwzbycXJxeal819F/vkVwtRJmsI5pCmFGrLltWy2TkRq
NdUoyEDn2A4GDgupeBn9JBZQ+b4b85juGEKrv5CXjobxrcX/67Swi+5J4DtBIkRUGil+tBWLPOK2
fwSlZPwVUpwHb0xkarY5qeRZyxkS1EwMNR43UBnL+pjOF6lEObd5qE7eZ6pk7idsEdnl0aD86VJd
+S7pRwUsy0+tAxpOZ8uzFPybWoQyvTZDOSYuIe3nIQra8s4gMcqwvrkzJWSbVyDu2LP75UaiPA1Q
GreHpURFeob00G/5f6xWfC32UZ2zjw1zf8nks2ljvhUb3JYfOe6C9lZbNDBZi8Si3tjUB6nlE4NN
iIM88Unjt0CzV4Kik7mXJU19eayJ37DCkknvQ6yxmdpoOqafbFMq07aIb5ZzlSgvawKq64yu1A/i
dZWwskMDHUcQ782g9H47f5yDQy4dBi/VZ6cC116D6VYG/7x2TNiAt/odreSMFKSdIS/iAFgGwlX6
dIlos6p5jtFJDOvne5ZnlDY+UE9HDPyeBcmcgIRG/+36l3bOIgi7OMZGbx8GbO7K+PYG71MuILpJ
Ttb36Gq16IlTlrRrRN/ovanjhxLFE8PRmNI2A0CuxKzA8TxdG55A19t38UHIqLubCoh/HG7zLrjd
36ZzRYGkj0LXglHySuAcXfS6t2hX5uCIYymahr6AWnj2QvZ9PsTO6gAQ9pE1jigz+ZELnIp9hs6H
i/fCF23+wAcy3LrkqnsWFtyJCbzok8EdhLpZXnF8CDlMjskLWDawpysPybiqz7kMEdASE0GED8cY
mO3gnJY7PPpfU1gEeo0n16phLEcKF5qHZM2DcgodikkgVv13WtAD0lH58JO5DMAR+furXzeayzNX
pbaOeSSzpG1rNxn6purBWsZgnqivjcdv/Vqe8h1tHWz4VHps2xavwm4lFJqC0IceVU7P3wBqH2F2
ceUhQRcSNEVyTyhJRpdWXg2zhhQ13NXfEgkIbgdLQ/XbvdiAhTpjJ90d8amQ2bZ+qs92dPJSWQVS
h96dHgnVgFmX+QyJHiKu0lBGAQkhnE4FktBtPQSuIcBGQQ6Ou+YdInYwt2C1maw+dLZcgo7zQFRu
VGo32pu7TPTTj2IhX5dLAlj0rkclg+RkbKFfh017rc9xMbTKeTZ6DKXlZsfgz1hD3FanKz+MquzV
MiAJl52lzVoqC6pWs6DJcU4ni1rUpkJgY4r44aHddtFaYlFb9lTN4pqTr6gRBl233VsFGH1uJudo
EogcrMIY4T4ujRonJ+pN2g/wFkYVrkQjGuS1+SbkLPDygWY+zayTMiwJvdRRNfVaUaCH5KpZ8CNw
mLL5mmdcbfeBrkqiPNR5ZdNcQ5T9QqT8H4jex1VoC9okLbTLsEH2JzL2IpEp7bTF6WySoAKSD6J1
EswsSLJuT2Y6w81999/2jlefYddgZVfFW4GDvepmoRcTdxPa8PIlDWjsiVzy9vSUqDdm3lBgt44T
2yHsM3AcqkUvWYKU+YSgNUSc5tuafKODDSe8aLczlOE/VsBZc3W/4s50w5B2/oGaQy1KEd/dQkIX
/QxY3E1SLJFF7dGZspgxYs7vtkBfW7P1rn3OHE/ZdQ2k6ljKgul5EBewnu+yemvt8piJBsq3qa9F
MtLCTRPkxe7H+r9XfXu1KcFvvkZQ3J2/MK8Btmc3ID7LdnozY8GprGU+/EpIX35ewc8nkRHa+65Q
h05gj7bbZ/2e7PmGQB6bJuCwAnkZqhlFOmXeuFLSfV+k6XULnbg5SHPgkj8huY+XHFyWLHjAO+Rm
ZKIidGehfvfdNkyQq4P4M961ghhiI2GA6ypX71WzxMl77sG2ieQQpSn/4iyxFLWCKXInjsT8by0h
2ePx2Rygl1CYZaVo7PK3yuSAfnMlr69p6J9pk/6YhdFkLQWenmqXoIRFQewxh7+2Txd0+X6n0D5S
cTaTfh+CqzfGA+M6LR7/xZRPEDpfbKRYnudib0W6iVafRgaxRxpKEBh37bvCWoc2kE4YPPIyVGQy
0exDN4lafbXBiEFb+31viHn173JNmqnqzmujW9nWFOL4DP/bbqdZnHveMClb/0UyUlxy1OLnNtax
sR+Gz7khQg8PhFB4O9w3w494arLJQ+XZP7aLgnTfXRx8REv10JW2w7wvC117ZwzWxJKa94IjMR4G
yNOYWpcoHY6nu8sLt1kUs4wlPelPx0fQKlnq4XeBYAeB3uYSSdK8KXNBaPgDi7V46yMgTBEZJqE0
pSayMAo3s8icfYv9EePqpO8xdTl4tUKF8hQXMGHws4WEoaJVbg+0XFcBnimfbrkEPqDjluhx37Af
a9fG6CJ75jDCsZ5Zm0EkFrix6l/ewjiTT6mzyyn9jL2x9v+L6f8otoF19dl+G+sS+wqyMC1uG2Cw
sRi+Ta7B3B7dTHTw82PpOWCTt+5pDWWbwOCYKRZCCZUG+fsOFGMzMbgM0PEBIuX6F8iFsguwDTyx
xZmLQKWSvkjCJifuDDtrawcknqhptithlL2pnuc2k2ATbqjZ1Qn8LSsyjUnWhH7Smzq7UkGRM2j0
dY5FlaP2SsX0M+LAOes4xxrP2gCQeauuj9uBWM/O2a+7QGs9PfuTOOfypJk6OyXLWS2r+SOPyMaa
Rqjif9bqen3IdGSrYbwYOzuqqH2TOuW9lM5gQ00mHtAWpMS8SnzWc4+TzZTZRxb2T6+kqZdHsfKa
OT15x2RMGAth0Ixem7XPVv7Sj4MiivlN5VUdukGmm8rlrWyvN0xaohMDJ+6x+JPjImJvCIzTHyGT
xKL3+BOip4M72pyUFsPZPV6SAR7N8RcJdvhcu5N5i6JM5nE3R/gszubsebuzGhau0pP/feieSu2Z
/VU5WXo0TWYaYlMYeB5Axb7TEg55uXapl3WZu7F2pnSIveQrDaYke0la8yDmONhKET+tMPgB640O
UI4DHw/OGNyoDm7D4s6XvsUioHSvYeI61fNr8NVXmKkkd3MoeC77o04G/dIp5oAmFWLUpWwuUHFP
K7ic2LXtFCfaVG60XKiRCNSp2CnqK3cZqvD5gGMyCnK4x6EQsVN/mz0CWfjVNp4Htbz7yVL94x15
5V1yJPlexXXnS5OYUInEwaSOC6ORaWPoW6RYviLuEBl4TTRb+sLX3IavY168Q698WkObmLOGX/sR
oB64GLKuGRS8htWVJnxqXCEypD6l482n/+pPTivWVZpwYnIuJu8QqZRSq0ObbTd/DtDt5lod1Dmz
t8i2U78plR/9a01W9jWqiVk9Vxq1dgmJ0e3vVAHuoHf+1OGzhfs8MRtuwnFMQsxFTQBo4Envxp1i
fmj0flS2XV/FsZNEXwlKSJ488VccAhGOMYj/CKBY4CDj8SAOVQhYAdWpOa/KjBT5QxNkg/8Xy4hq
6cdVPgmSpjr3YNiRxz1t8wwYR1UTzdrzZz2U8VrpZHrtC43FcmBniFxAeGzyjQZu5dcNamBqCJ7R
Z3yxsABeZe32G8Bc1dHnuoc4KmsrUS1U5Fs36MX2wfFW0vZnwUVGO0wgCh2QThQPqIo5iiHI2rEK
/sCwte9682uK7ZTTCQFCARn+WV1oKOlpdxk4Hrwt65Vo+QNuP5LAi6zdULFr/XA7IRtFxHj/UPaG
55Wt5HPwwhppCazLVskdaITzOppjzcryJj+aN8tKKfgfyj8OB3sPyvnnLcwn3EFZUJ+mFrwcpDlk
JBGgGfNNNlpW1O6l6PWgiGuhRkiZo1/t4UcFxwTpUt71VtOYH3g4/F1PzepdEqXM01sRiaiKuZML
u5QSfN/82Vn2eiUDsBUlmDmr2wh32wbliTJdSPZKg9AkECR/kkEvok3NSbHAN/sSRk9Dx60gLBC7
3Jy2imgyQ0M/MYWJeFA3eJqbKB3/j4NGSzH2GqAS75q/RJXmw4qYbOuP5jvzPbi3YyYbJksmSRVs
qpF7vn2h+XW74lI6Q5pfNUq5wWXfJuJ7yl4JN6J3k1j8jj/8JARuwLkRI89DwSSFyugpWX4SLxvp
iWK1yen4io8NgtUslZFjk8A8lzdWhDhDrHgTZPduNJEs65NnpTsCElbOD8DpDICshSSis0z4ZP/D
oPzC8lwnC2LIOSieFSXx89QhRfktFjkQm+wyWGRjCSAsyIb19l3jiiulrmsEUBW2wX8qm433lXyE
JBqfHjZWCTDvZANa0V0mWHvQx2cJKXaE8ygmwBZK3U0ABJmyR8h8qd98J6dCS9igabZI0M/C+Yel
BE8AEQsWR6/3PWbhb9OcqV8DyzfU4+VNN8y5m/pbVO56ZEY9Apk+lSepWM1mp9+1bDyyCwq6O+iY
dFLOzAou+iBayOWEZXDB+23eP3S9UmTLvVoqxU9rVg2xYG6a1RljJ5wF2oQaZGwNbryS6omtnk6I
htE74RcmsmvVPrcrZb+doUUfnj9GavAfTUhEK0gqc9crSAOOSGU6X+Oj6JncbS2V234bQmujkpM5
GD6FnKD+U4gjzLnzksNVxbUYDD65YH1XVYCcjWO5w6eFlM13fW3TZ6HFCL682cc79t0F2r9+xtwf
WszkJdsR5xIPz1SE2zVs9eXVekzL2KY5RA19a6D6uyoNTdqBL6pK43yQLuXk0p1jLK7tUO1iRjMG
zT2yiGLFYBoOm+LEXF8cSkL7TX8lGEUN5jwDRHS/ucp/oPqvRxnNKZlE0dIQgw1URKFsKntfC7Wz
eC4tOk/skoLBCbym/QzqNcrW6S9YSMuO6DDXu+aS2EIes/svuJoqPv9+S8EYFXsxUebp/GiB6wL0
WGYKYftmCe8dLUTqzrc5Y9WNSkePNqyM/83gjqwGjR7IIm0sJwj0qyYSamzmjAHC9HHx1bxgiGcO
ZYAQlRMDIX5NcvFvNQE7Xfc8ju4KSB/K9UEtCafaT5FT7OehQO0gIC9GrbaNOO0aJE8xBWnh4wY9
sGvg18t3+zi9xm9MGk21QuR1up8fTBhwqksH4Ia9/Qexh87WxCmAd6vO7G9R9lyv83ojeurdku5O
8IGkyeY+OFUaf7T/zHoDvUkyLU+WP+ObLmbcrb+C6tPo5n6DWWBMulcA7JOqBMyA++wlMDRCEp9K
RXktJxtSDKwoE98Zf7WbRGBvLQsmJJrtE+8bAfUa1YNSpFwxE1MfofkT1pzDqWmG3ex3T44bLr9h
ob5jPG1OHbAqN7mSn9yHQxKoMFgSBCG0S+XB8q9aE3vK6p5AvO9HeejNOpZw5e9898wGk0hNzW8o
G3Y+OvPU6DAhAeWwvIV66O1WIeFFl+AIz9k7JuDMYo+lrRE9XvsJHG7ZfdGIr3qtY4T3Zl61w+fv
UaQqOMezV/tL5GZRGD97cjJk+dCiSPHeH5D53Q6T2KcuevR6MsSAzGBUb1Yy25hnxoVP+xzo25SS
IpYBBnULDHSQ7M/hsLsCBSDhw7kPi5inPko0OMxZDn9i5RDyMhol4nFWVnX0poEoE3meGzMZ3Cu2
eKg4Jw/PkI3S3HpY4r4o8QWIFCLH5uEjgnlxgljETpUiCSGyc2Qfdlz+8K86zzKncHORZNE40haU
vINr/0y7qGpdT/MPVa0olQJLvujbh95+4KP0XdOmcW8SJJplSyjOq3YQrIgh+fhqC5e71MZTzANx
mqy4wOVdScscW/Dy1RpF2hHU/4/ZwpyCTwiPM9BcnuRijaCwES9iK2etl/XUyTfSpqnkUp12yGfM
bS+DVIuVTWYSeinOQMZgIXQnyFue5TAwatJeAtKZFgTrxIBQFBsWQM09/IQbbfbq6LxJxF3Unldi
x0OL8fJkLDXhCqd9sC+0lzAtT7grI9ZWvoLjaJVy1R30644gekUvtFqnrXuKqCde5wWovCcpb7+w
j410/O0W26DJ3MoMh0fQxjAHq+3CRZCQ/yxktxFuTO/V5lrYkpfH/bsqhA==
`protect end_protected

