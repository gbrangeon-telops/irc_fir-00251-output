

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Pb7E+qNVEP4sE5d3TkwQJMYKTR/FjAPrexB6qdDJcLdscPV5w27UvNCqw/kg86JgS2hNrfoEvTNF
uJ9eNTpy4Q==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Egq1eCtVuCp02bpffloqFi7UMw6fphk3UOZCcejhe9NQNeC0Z0b1+S1NY8yEfAVY74l4oz8pZ1vA
hbrAzplanZae/BDY57rCQ6UjD8G9keaOwYv6mG13f+m77D7Y1nVpXOE4Uujw3cZ1QgwXR1H4YfYp
ysjb+lxmo0pqYRikRIQ=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
KJqrZ5TKkbTlecBRrKRCsxKhAd1omWJvIin7DNafgTE5a5N2or7GsTSawdWWjYWHESLBvStvRGQE
jVUeK8m63dYVJN98fa8T9iAHTDt9yiBRki/VqfvAejvDOEI+l8row+LhhHMvCd29xmkCeQKiq4Qt
hsdsz+jNufnCYY4Y1CVO/4preMZeG5Ow85vRd/341CoWEOBji8o4pk0XyIttBBgjBzWO8JyhLpza
R+Z8LgFoZ5OTfgpyTJ4SjYRWp9IHP2HL9TShNo3PmM36nFNBvQSLoEjLgk4+rUr657++ugJH31/C
Y/QScvwJcbqMK15awb6twj42y2gxJSFzAPzSGg==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
KxmYEF19quU2lnDIx1hLVbiBV1iU7MlwBSbpQKNAVv6HLtZNpIjv2UPtz6sPs9Xac0T26s1Kjo2c
fAw+uaSeKdgWE1BMMV8ya3nIO40+wJlyaPYGp3qW9dt6kM+FZZl/3MCpgIMx24FXg4CPHrHNKu54
/3DZJ7o9x/QjyM8WSeM=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
n4InNydlMoO1IH7Kq1VdB5tuRxM6d++erhleefbfKU7rQGdfSjRtqcQ+h67LKfA/jQJYdDdZMjd3
Jp84+E2i9v4ovZP9CPOifgPGXKRtOz0XzimXarAjLF+OJp3As1WqoTrPJI1DspdbqtDWx5caLezn
hcZVfRSFpZUoLc9H0HW6DXtxAWvJT8e4ntjJYO6koEzzHlZPpMhXvbbH/rbArm4iRGWLOVN205Pq
oJcFHv1n/e24XGuCRksBqssUXd+D0UgsxKn8Hy5kQi4Q8xdFEXxEOVBI7ivvG+HKnJFOOr+UNhLY
+rNFOKSwlDtT8tPfpzjKS5GdaTuv7j2GVoF5Tw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 21824)
`protect data_block
vlB6dj8SH4JNshs991OLofCmcy6aKxmE/aUeTjGCsiyVJ4LGYbBxciXmjWd5Xvt+YX87c6vGJ8vk
9iAoQLnaXKxbPR4+S+PZoNfwF8Uw2oq2oC8LYe2cTkDHoI6qHukaYx4j/nV4xPjJkNw6Eo3BoymL
MVpThxuvsOByxGRuH8/X4QvBK0ScwqmBgtDMcLFSqoLsngy7mF3itsgzcJMpCDEKrlBx/bxY+OLC
9PdZuroVTYeo79CwNvVBQ9WZiNfA4XQwgeyBvWasG12CE1+W/rXIgyb307xT3D/9oIZ0E9z2gRSQ
WCjD0wu4ptBgP2H7FLvZbivhYO37QW2hgabuw1/uhQg4Soigx+e/85y+ZPk07WL+yMyH7Z4dXEwD
NGZWCUv2qMxrr7zA+aWMgc0SKTxDg7INAdh9TsrtYiAJK3r7cAZPYJ4f1dMuTBkbG0gZsVmfuvsM
GXoSBtDx3B2jSlPua0ZDsupjXqbyP7E7NFABFsGIjyJEESVipds3rd3EXY8jbg1KeO97Q1zkuTzG
uQz12OywOCKt2blzZFYbGXmEyKDi8J7wdO8R5GyxoiIzTrVl98CdiBl6QGkQbyQ4xZDozZ1H61wT
+6k3lrPzit22Z+zJFDsdfp1t9AQSmkBZ1Y76G3MVlP8n4bNE8FYm5dTq3dqzyfAKsVRz8LuqDPrm
5EAX7BW3bSgZvdOtoPWBrV1l5jIEMhwPFQH6Ooxe+EtbC1DI1SLE9SBPBT7UDwP2VxWand4X67Os
xe23NhKNG8eEb16zcZ+tSP+ctusWTnYMrAZicMcOgnKbr67gTUIduq7ewZb0ojZfUDmHiTzEewzJ
sYMpQU+bfLPo7Oa4Gfi+IGa+LTj5F9YjN0GDx9Fg8z3ezxIJadfP8ZgGtmY+qdsi/SFcCXczhCkT
v9ZD9hetluIGC/nQf0t41psX9K12TWY5NeGo28zPd5CEKMNHZHidw8lVRnhns+J8MXrUS0GafJkK
Ywi4gsI4XkMDFscM3SuSgKn0hE1Y5w10j1Fz4gMD81Uo7HIsqe9WFoYOuIgvAPIU8GxQgI4MgnLW
xFXt739jxBhS20xqRjB+WnhFG9jYA1wZEw7a2zvyIhkhoGgTRXjwpk15NEfx8dr3djbW2gmb2cwr
HVBnh/CT2WRPSca7QHR2g/5mvo6oXLJot5SRi9bN7u9uMpxvQ+hU2txQEsjNcBn3SY9psock5Yd8
U8kfKpV7bHFDlv2xvav7G+gn7dvf9mO4TI9IymP0D5Nf+PaQVmYMpeoi48S0ss1ttioK8NzYDWJ+
ytuJf0Hh8gDFMG0lh1inDKZCIuUzKISi31bvCjAhYd6Y7+pt3OnUFezwUHIIpKZa2rEn9Q6s0rnX
r4GVhYgm4J+Xhtfi0eHazTvOytJz3PnPGSbNqnaZuMX2Qabg2GNCjHJFrueQEEBQn6dfhHKaQ8YB
5o99908azCJWJM0fVvTqEyrJYssjDdjX4F/yF5Shmw1wrftt2LKHLZd/J8OUCIdr1da26duJ81ly
XOjwG7WMJ+4dGqBgG/ZVS6QmGVfsaWr2sM8AnrD5FNHlMhkCwelz0N62iDWngYivc2/0lLatWyfG
2bF1jJgawU0lkeSneZqFKWiQauZ/EK7YfFt+FZFmkRUzP0yP8/Xt/6HzaCnlbfACjoPotfG+5UH/
g3r7A8dyIFvgtCMeWFV5NgxnWbZO9dMVpSbTj/mdDM4xtrCV6GUPO/pD+MPvUDhziagmj3jEbGDA
pyAkUVPyEeWOAhIdi8NF+T/5D9g5W1+75luW77wuV4Wz2cD8DSaHd2xZJP2mfzNi8tWQSFbM56Nw
Z8D+gWO0EM8mcAAp7GJmKiJzuCTQWP3h4pgPZha9nDViBznkFAn3PTFkeOPEjBq+2NNvYPf0dwi1
wWW5X2HKxNL14F0QW5Gae3CJFCIPOuKv8sEIyTCVk53ZWNo5+QB0lxicUFfxegeHrg9aARXRP6e1
wLbm0rLzRHnIoQnZWDYO9a7irvybv+/Tr5I2k5ASdHezOHQW5XMptiAmGOqoGhBEtPTHh+QEKB1v
fzgz5p2msAIYP29DpmhaYtfLMnYz7YS3zZrGb7T2GO1v52iMBwtmZqxBqX34iPb1BDy4f+jj+x3A
3T4KLibssAWLatjbzQEHMDnsZvN8Xz/EXCX3hiAVKjicldqQHr2CwdD9U3rCNEOtBP8aMrrt+HbR
/Nhqwx20Gb0CRS+gpcxor/gQBm/SBNZO/urXBd0OX8rD31DLECJhhj+DaSmmassh4yXWyLXLFRYT
SGUoLZ7HeqKjuiD4b9NfHJ8K5hCpB93K8t+xIlaoG0ZGlEZi+Npw931cHlRZetf9LXMZPUzl1Wyw
+FrEy09TE0byPRoqzd8ewAS+3NCdniV1L5dS1p0EsT1BNd4SDonKKymGSqGZ1z+m9uoOPIQqJzrd
+ePxPCxmSr4VWH1Y3SJy3kZiM3rhjWEutxf465JzCRAoXaVyMJg0eL4VCf4L99bYFG/IIN9JYyDA
8cE1SBPqHwCic44mZO1YM4gOz4rzH5iBt6hmxXMTFqcaB/Xnxc797wfacexTDjpYgG0WImE6Sd3d
C3PC9F0Qp4y9mMfZkvEnlOtHFFh+jTaVZsZk0ZWTfFvWjW+x2mvgnaHsQ6UlrcozHWkkPf2yOB4r
NbOha7i/3jgrAqN3yWVjfu9AZV9xoSJAnw8wYboDBatTYlgUEI71Cos8pO8zbuMsRqskXg/4FtBp
jonMFYl7V/eyVGsluNSJdMGNhNIlSZSBp3mJqcBeKF9VvglGWa9oWm+dPzp9dgcJ3bJY3cJFBTq2
OopCCvaWLLzJwEbb+zfA/98zFfTm8oDzH/SQhEtPj4Akc61+WzxxxSI9KdDdGl/q4gt1Zxo8KiPf
/mUvQsHIsOKkGIXI6QLqvYReTO7OejhTz8PCw592pO/lBNEF4FJB6gp1pK/wAELcVXTVJrVOI5sV
MzIssOrQZ6WzMCkaDoNGseNEeBytyEFAERMWgTxb7AUOQmRsTf8Zoc/7dDkfWICWa41lMU23GCIS
4D4NkFmpWiAO+K6OmEAiisZw0G8rsXmgKRdymB03WfvXN813yrIpSTc+i0irxWLOR5+1/OZ0ZEb/
zBtmjiGmBcg7UIE6/anPRFx/yhmLsV37Ynpgixx4bLQpiGs8Ze+GmU1Bym2UJn8Y0kyQtneuciod
wMMd3w0t8QdP+4HUFf6m6j4IHrx+hn9hC1aoiAXFn4s5jxiGYSPBmC8Xm+5dsIYq9wgnsPuPua7N
0e7JAq1sH/OOoN5ToaglCxyUsggVygHDcPygi0bctZY9/pZgsgl7kUitMYRppoLoaA+iOqRnK5xe
UA9u2O7b4TSJ+y2NNBEAnZcvy/F2jejbaOGjJtXizn3K8QQzLcuCWdBukMtYEO5k48tUrAzu6DdG
ssAymIiq/0TAE4dLQycM+JNQ4Xx0qiwHCtIkT2JDq7P8oypPLwvPLohG+v/TXW4ZwUBFfyhPXDJN
gCzDsp/2sss7UQAwZuMk9vMma/cllUOeq3VonikcQydPqBgoIPlPxEdTGPy30zIcwKrN2ibhyU5K
OFssvmJkaLX0fxms1O3tnPEAgyWfi2MWUyA/LHywDZ2+Okbv66D4v4yfUzAyePGsLddpEeMabIII
9dQ5XIxp2aspoUD21bQVgYkvK+AyRsCwH2E9Gbzh1ll9Zd/Th09LY0PDwYH4gRT0wOsqQwKk8zzy
CYE01e6yqlCuGg37kD3zHNisC4B1eFLyML6uGlYGmkqCIDIym1GPdsjkwV9D+MG4AfRUrN25H6ld
lmYVQ+kYqRMxLbv1xFVdbr2+VR2up0nA3deicgJrkqgvi/10vqJ2chtoUFWeM7puRCuY6AmzPHmK
QHvKE/wtFMpVi0xwEnXISo1VGzO3hVtDiYKNPW4EBanaSh0K5QMoyj8bnS/W7ZYdiddkkf9SFUSe
MSA4UUssl8gPh4Mj02goXVCt2kTNUzxJYYHKJtnoWKw9m4eHcUJe93qc2Am9BFVOD3dK73VI5pTA
b/n/p84JjPHyq/H0vQ8+vCzkSAXrUDRhuERc64x+BSC1uQKcf8/7nUGoMc4oL4vdOBAseWU1wlV/
bjQMa8CksUGS2G3n0onIQU+PJmX+6PPaWKJPzSw8obgH6HU5QcR1Mo7bEPo/4ED8XHK3NyX8zFif
NrphkUGJZA9vX2cB5sOVWAMplbY8mvPB6ZDrkXpYLroj50v1ePL8bIY3N5B3bda2B/66rgWpZrVG
TzjWr+qbhxAOyyavWZifjZXvZQFpKt5kTAt9kOIwOhrU+5w542qqp26BMLIziGE3nKOEXu27HXE+
YOh+3RftYby9wqjc5CHyJQQjuXYqZS6Pn9Pjv8trm3opanUlLYIR1D/DGi05LFEKmXqd0+gp1iBg
L7Mq/1uRMhtOJlhlmTT3fLypD3j4KVIRb9oWIF1g/G9upMJ+cujMU8p0b676Mf7NkokkSlg0hTXn
QdyL1Dpc2aHFvn8YhY7M+hpBnM1PcqtMDMlEjW6q5Mu0NLxCj4G9+yeVHPQcNcfFb1gAtvHeBUck
907pVQXyLIEmVmDGdo2fytQZPioa/DjfmHxkzpa+DFFW8Ds4ZBocHgQ0gFv91QS2XzZbvDDKvn+c
FvVZMNsoPwxZZYdS51fNvV8qIZXXmVY7brp995k7bhoLjna+UXjP/SbeWUKrFeln918DWQbMydjT
M9fy3x+x3qDoZPVeVI8itIq102n0jktWcRSr01vuUl7P6Icg99p/4lc3S+6DBDKGZo5jewrzU5sR
FPYWB8zdWvfHwQzcsUIXrtlKbl74alJhxbIsiUcGdpoiqsT0BXUnlHvR7tGYOuOwK8DrD/ETr8Rx
3dAOlBXjYgIihquGwWc77Eza1/EjfQNDVdgN63FecSmefoD0kvzf9NYLxHFv8FgJBZY29zXRSLwU
vDcQFpQkQEFlvvqs9cL9OpnNz2XyOW4CbLVP4q+o1rV+tLhPZg9y3u0g5B9UI5czdHU2q7PxbpBz
Aj+EQEzHnzMDHEevCMuQZfM0P1Msm1eP8ffVFb6/sJRCXg0v0czX0NcxVgulUzfQaPVuEZoBERki
oC/IVMiXAAebZJKY+B3V61oFQxV7DB6ADGXfQTYhB64mFjig3CBhaGUNKbL6AtbUxV8xFPfWK37I
6cdvSKVkzBRxmI7Wb3RClp4dpvTAaDO5R+5LH0keD3slTSiwohPLKRrSIz94NG7rbV5OhQGHuQT8
OUvVw7PBq/IYU9zhxRA38W9bb5tEMlrvim/xCWXTIEPY+oVX/4L40fblvWs09S37NGFRpCHYX6+4
QUtkUtaU+gTXFcPOUEAuO6MYx/tppqwhTmgcBcPz6VJNbXRJdADsEwbqiP9dgn8mDwt+CXtHWOaC
s30McTBSwSNh7gcklMCE3y56WKSGqp0GkbdxH/zhGA7ht4SX1gdv2A/RofK/hmCV955oAJdVSZIW
FAXbmAvAxsl5ECDHV967bUaUGyJTzw5+PVGABBH/1zoNnw2S7m88okGcAZ2a+f9uKF54xeiIKH77
WtShA6uoZpDGKZY0+sjbepLHRcqkIOpux1B+73/BKsjvxIdk0HN5jED48A4vQag97fQy7J10ryju
l9Ma2gPz1OCf5oxRE/5tbQq2GlnHqL7spK4JwrD3QXaTj0aMS1a+DHx0SaEeskYPTOqWPut0JzRK
VxKY3i7ywNk7TeIfPYYH8EhTwoUgNidclezrxQCb887dnPhQuj3O+nCuEttwUCf00gY1ANyEPFqK
fWDHiqwPzitpCDMFcCFJRnEEAEYpAVNUmH6NpNGdhlwVzbkjX7QHPudWheZdVeyyCUeCpQEv6BJE
8bErikwgdUprD+zPACMZ9cIHna06KU6j+gUw9OlXOpNoQNvEIw+xMBS9r4VFHAH6J6aRHqnUOZMV
kEhFLAZRlvIC+YM8+ZGU6Rh92oBoxFyPodI20g2ZGlIr4nxR88eVJQBVdj6meI73w+gB3OguN7kG
QAZnWamf6RzMoQCYr2uQu0NWC4cAQS2ViPx6PABfIiJgX+S3rQnZ8Xx4yntAwoRkoYCTrNJlcyhK
IVsMJ07Jro6qa4LCfeX0yEIMzxcyN3Hg7SYMGz/bHpU9Wp0wvjwOP1TZyA62Im+Iy9qv5Dlb4GDZ
4ABle8Sk74zd6h/O1W3Ys9TAeNH0Z8ZxxE7gWlI03XMO+fCXoX22gdwi0mafXLPpYqenmwhWglNb
LsE7PutyJcPc6i3Y9JwucjlLNLC/cN5yIiuFLZiwZ+EV2wgKsyJZVF1EEEPrhji8JXq2F9obYsMn
3EHAB2xlD9aiHKHQPF6IfDJD9e6FRq1cQ4/y//K/tAnDwgPcsemwSoi8H9Z90uo0U/ZOIS7Vidzt
INJCaWwri9t/Uewv2MWXU/sSYZZG2EftB5ivFCTQu4GlAqhvhdZHZmBN7Fuq2GCGaevbMp7lCFJz
cL3GnRbnLNiVfdWyQbmRugY9ngPdWcZKelRt1ZUjjApFTY3WiPtFdlRYWzl2YaJx9Sk8W4ym7Tir
4qs8CI4eaFbHyPPb84b4knYIzkXoHTF3UEq9mwh4cXAlx4ps0RRrhyicXDsIvR2YEcb7kpNFzUzY
vUimLHPXzZwLnjWZGtf7BuchSLX436pGOvvxFtj6HxAdsG6rkwRC7atRDUcsDTx4KpeXjRCvoFqV
7cKpG0N33ADXMmtkRprQeQuk4ZXWZpr5rjXNsRH2RP/D1aL7kdGxa70qljEpSiKEQxn9bnF/TD3a
47CffIkJoq/dJ/1cBfSl0/QS5BqVBSWovzf8iVQd0ZgsWrOeOSLzHF2ErUJ7qu3cFyh2jGeJqBxl
ZZGDHjLLfjFnP9CiCokkAGvi/ByQ3QtwFayTS8LAngESOyxeQH61xCIP0LkHzu7uaPzpplVzkbxz
QTk0TkwdnDjv8KziP2oTYRE/9e7dpeC2DC5XOp2F5lvDK2MXxJ35givRpEx85UFEFqqO9dOLR7yi
ug6CY/E+YmJwKdSlMJd2l9O0NUJ4ZYkgEjKaEl0msQdiN8KVWlg+Nuusr4qGXVCgHy9ABsVtqLp0
jGkzt99cLD9aa7u7RNbBZ9pLxVpxbGvqNHGbGB6zb5+F4eChRarqL7FLsAN5pjgJgiGpf6V9qe1m
R6uLktk0T55vPQFl0T1P/AKqOj85XFJzDaTHb6ZNJd62J/Re6/3sj+3K/NUB5WAyxCr7dmgkdBGH
b9R+qogRdEO1fezHGmWNU4V5Vs6L2xYgAadH2DjfQDrcpllHeeEjv3niQsnzNaAT6V201/HyTpZA
18FxEtdEbn9q7QA1xFJt7q9le8pzcJiPs75Kd+i69nlgJ0QCTQCSx4vS5u6bg6z53cu2VgYs3BQh
titrXj9ONg95Df5yHsSD6z2UxcwaIDZtBZdVaCZjTZHM4rRNylMQnw9s1Yzsp2YfmzzAIwbYTYpk
UxRNY4QhLjO3KftPH5NyjKsEr8rDv5J6pmPQorpCaSwM6fY2VZLIFkVwDipC9Zer1NYEpYloEuI/
sBXWK3gUlc9syfD60MKsca4aQ3hYZO6YoRq2M5ZVxhPkEyR/Ppuisj57x4yniiUw9f2DTrv2MMNs
PMq5Ws5jk/L2WzgqQzCK9FxODjCDR1MzlawQmJfFaEZzgcH5aB96Iq3jT/u+dbOpJgeznFqA7+aU
6jEGiSBMMl9jA4ZCTEjjwqB9JH2tsv7KdUYnSga3J0yNfDbRxrTCRYJIWFObmedGbhzCEX63167i
lHdgq6oh8QHJrgoXVbvVag9IfVRraj26iAdIvnhOKgeP/WEmuOqcokyFxIGv2ocaXFehSY39AIAk
jnQWekn8KCec+Pdyha6FHiYEdEpVAVmcBhRlOjzJnXr35E58jfKdXtnXbPJ3fZTdcepfx0gnW5i1
zN8ak/an1spVvC//bNoMRNsaBBQRkweOq6LF/bPqWg5kMxW63ghfw0R/JAYm65G6ym06DeWq5hTs
C0idkrLR+FeBteNW0dr26avJHeGzL7HJql+uJIjrHueCfzGjUUnSpDttnYnIHA/GihJVI8sVKNR8
df5rf2DAAf/vYFrSOhGqyHsASzM83/iuQv0GU95xFVZxKgQ1vl+MVFpCXPNNxPBacUw7hUdQxx3c
E7KdXjQbuq//TL+1cbBA0BbcD/+2+AZ8QiTpnMmuQyeHenlOeR5CPS/jksud0HKBxdXd09Rg0puL
PWmqMKGwYuJJJCNOs3+Z+DwQoNs5MnR7c0QNSGeSNcx35SH+KO7PS5JCvtNSknOZgXZFzFRhHGx/
nPuieGbJ4ywh83Ug8gh9FgK5aY8NQFQyzpVmjPIoi8yeotbt5cGAUys9GGbX36C6uEoXt6u0Y/GI
k05M3qu7Igp9bJNi4OUVPSb6hmJJOUyz8AB4lfurhGl1XCkiJGjQr2sP1sDPM5BSQTh1KvcXuErM
/U3krcJbNm6a/6lwDXaUif0m8G4+ZV+EMnTeDIQ/YVcBmCzKUkWklF4DOSUAdnjtG8NhrpoR9Btr
j1lCRAKIb0AttQu/dKyoRRQOxSTfjeAavObAlDM9/13iDOWd5R+OV11Yq5dT+n28xqsteiXbwGT9
sgx5IWYIfvgfoNaHTR3PZipI5SL3QkypmJawE+3HgkWvFczAZvgcvcWRA6muPXjJyrmzAzamn/48
ERpSUFRdNtmmQ8bhN3ualOeCpA5foILqGEodXw2d03CYo0YMCU8VkUytmQ5CmAB+YhFl5H5GaJd5
c/sQJfr1qssEjKcaVa6y3OujWCw5EdLvB2peA4jvgWcGbjIyOI7VqPi08B0Rks50aqbuv3latFEC
+w9cJhlv9Q2xBrz31iqbx51+KUHxWTgh1QlpVcBiWz+BO8UCEX6hffW3b9cb1NvEgwVCZo4vHm6G
Nc020hRKzAq8JjKmdIenCOw4HcbKM0gpno1SzdISSBeF+CF04CJaPBSK1cfpzY2Lgi3Pbpo3JBp6
szXbpeoPZDMlgGki+li5IX9NEQdcFi3R7Cx62RldusvaCGsNj95Pgs2FFYc2RrL5Xo2CsdcOeRt3
4ryYTsxZk5QANsCPK23xgE99xTMtuvA/aFxDPxPRxQxUv5wNCBuexgOBqhkpoaWnvXo/efwVgpqT
BAehE2AnQu8cMt6mvSzlIIxfwI/iwXVpIscHhWMk7zapyk+nua3buKr7Reu2x79F+BqUz+hTDlGs
UAVxIvZTBKz65iBHFhwyU7xzn4UKBPf84on+2QTc0n8dWTvJWYoBnDy+xwh+szsfOB6/vZ7Le2m0
JcgEz5mJ9+swGvQWg1zfBhRpiY3aMJDEdzsAjnCg4hTGrTOMCj80zE49FHvGg743Tsube+HpPFzf
FAgqan7ar8wUpdYdc3WvE2efQl7wuDUsJZVaLudFSJheyxhJvKrNlFQmtqbxCJD7nMZjuFn9zLgO
EhLAGa+6gfIohXTMygIGMKGjnLY2RLOaNq7jpwAoVkQrtm7VxVfOV0Abnc5fA62+NLjbgGQ24TVw
x9qPBhoTuJYBWwR+YpyqdsT/ZsoSGo0ig8NWSZW4n4yLcF9FNmGyMb0XqpyKh2z/FEJKvgouigmU
r19mQycdLE3gq8HKzpJ5rz/QLMppAvTlcDF2Qi3NMwtknaM+xJBXTVd7Xh4k7wX7zYLAg+PhoxEc
fbCXFpcjzK/EpUVTNG+lrhts/HNKFtDgpWDNoUVqZQbUV82VoA/cu5fxUAkZKozMkh54DEfd3eRy
g8XfM2ElLGR/DpUM15lCKWQJFZM8Onnlcyf10PJdXByuo9cHVaiE2p9e+xp5JzXpCp3KLOpWxvHL
yaD+dk1Ktn4TVd5pn3zF4Kxrx9wq+5QGGPiZ9fcphcaQQKi8b3JncRKuEWMcvkZmmVO87Vz9ua5m
mwUQEKh39erx8W3oRBcVlKlQ0pP3YfcCCfZMFWB331A3L2q+eOBWwrY6V+zAlmWnSZ6x8CDDEcWY
qQpPiNkutGL5YQrpb5fSvZEjN8RT+GuLpJ2gtJ1dSJbj1M6FoAYAYQrSUK99Y+hNMvQmDxiFpwBU
AJ59AMQXmhFfaD4MxuZUJnPE2bmDLcIbacF/ZBuhKBBCAE8x8Ef8R+J2PEwiPP7sxEd75I85sGOQ
zNVWQnSNyz7qjKUMXSpG6XPy2fcQSzXoqLrews3AukAX9CxoH/SghE/VGUZUvOI6L3IHG8dUBumK
8m+QaKtJZo6dOLJ9lz8liFJu7meAeT7+XXsGqBg7Jol7MjuAiEAz9MMEE7cbXKsXaHZ9wWUjs7ki
yp6tqemARaxXhJ+vbpaOIujRGMZ10o6TrUsl/5r3HjUmEmjU1U94alHfW1FHj4rnN9S51I3qgP/i
vBWdziCX5aSNNSYo7m72T3GdtNeskSXxvXJDbE8Ohd8Ywr/CRJl7S8ngXmKEhkFxRRJyElqwRfoz
U9ZJ+SCInbsaxQp/xMvXjAAaRc20gljE3qGNxhFaVWO6aDWU3pKW9fITO286070nm3C+WW2qgGGU
1J/XWj+NAy/12Bpi52eku+OMe5PAjqAddI6+zS9oKU5ZjGlS5m75HQhRsxFMvWVDImeixSpB0W9a
FCUWTLaks4KI/XdgofQGuYaI5409r8JaB0PQ9KKKTL6PgBVSmUjXXGfiVbZ2Fd8JK0DrK4CnibRD
JqaMsy2hgZGGEgs/v3OdrzNXuYvUESFmJq3evDtFl14vsfsrFI8NJ+OYXo62Kw1nSiHHaxTnrTgZ
Jm22JcFv+r+3pL2H/eE7mfInbfGqoky8FEeKJGJ6GFK3OLbmdMIKCRt9oHC83IzpxjX+UUKSJBaC
7SEHEIb/P8LH0ZbpKBjdfdoiALb/WKsLQQmue61x1LreK+W99HxTdJCZYqYf/v7I7f4KgryK5cMn
Q44KkUMusLR9svZTHwkT8dIURI7B5kB6M3uzf/YusG7++5PSnrHvrc5p4Xw119OlAazQOK7FGuA/
WEYJwv3Mm25qjbF2uNfMd65o82CjYcSdbk3+7PBQkts3E6uNGuhOIFvayCB3dFis94R8McYf3Z6y
Q+4PY/9sxqcXFCqpXu2iYBRivY4u2RgBksQ6c6i7hvKxzUnfG9hIdVIxH8GdUxYYE2bRHSubYK/t
3EvzytCEIUuBGS24Hb5mhYLLUoIHqhMqAbfUA3DM3V0GBCUBUtJPnzFGLX3Krw0UoWycIyhbfg20
HjFuYtc3kJmr4VuT2/j7aDR62SZS3hXX828oGwWFNV/XMqv8aKropQ7sZwlzjLmmjUoQZqF+vs0Y
UrrM8ykIJSsu3KUPoxNe2mlq4o4BOdP4BWWiYchLHHOybr2dI0O76nqif0rHGDOaDlGo+AnHLekR
S/FxJYoBx09Ew91iw2sX/5ivZ42ZVYOJhXF+V6dASlvGJSWkoFU0jQErXfuuWAIL1IiPzBoCLwWa
pBDqT/Lh85HpowbDyYBI9hx+iDuhLnY71WqlJOdpNR2AfdvgaYTbob5UWQlL5LUrtLiyLlxPPMdz
/tPrFgVh+Yw50JRZkbFYPxS/uelomdDG6LR/SG9g7VQQEzTFDK/o+0drLJ98yjJnFHgokoHYGuCM
v/B4BUvIwd61IQnvCtgU18lSHRndg6CrSGuxlRUKFcxURqQdUrAR0opfIWgj8wWHSDl7NAlDrnSW
I2zah1coMK7xPSdKJJKFfiFnncqZxEw63Un1vIKb5u/L+59eYrsbzVsdSVtE9w8onrf06xjifk94
HlGW7x8/TKTJRkbXCVLeniiv115BxRiNDH38z4FmkXD4OhJHFC+D0/5vUnFOny1n5GxCMvGKeNeL
3ATy/SfjrnZ+xm4YbWYvtmy3g4NRcBjNqHJyHgg/X2OEMHnMexxlyIau+LuAFTBEjyLmIaACJsmM
8gZJb3aH19EIInZNOtnmzEDR5Z1P2pHV/VaZClhj1PHelnBCG2ItPXA+dFojeHXCaOJmcy2EjzNz
YanuybaO5tkc0TJ28ACjwk9WCV0FSG7LiMO501iTOPCGdATnucBntoh1RN0UlDXD+8G+GFI5pryt
++gN/xVwYA2TIJmLyfLEFYJ6ADj5+xOIX/UUpAk13ZjAiKKGRrwxryGfufjJCbhvkCzNXXjM9lp+
NPrsURz6HtSu4pbu0mTClil8PdpxOh7x7rH8COZvfPr6G7rqAGWb2cchG7D98ScGSBgB0OFUKnDa
tn9ZpvWRycWA8wXYPa9fUs4jOUA30aEdmCsp30b8mso8JkqiT0Zo7QJf4FMEkR7/pBZbWS1fkLks
STDvtwYxnn9qV21e4t2QsMLU5JlULVPvM2sp+dr5PEoHryegDyK5BfW0IUsMyiIpC0gBB0/5zBVP
0505XxO8E+Wrl28ECj4FkFikkKwp/5JlcmP5Ep86CD595IznJYxOFu+IPg6ZMTrDYvl/tcsDprZW
A6gtSWVcdXfUXem5BGnZ6xgsywOkauSP9JTat6PGzK5/Jvrv6sbn5ScHdBZYIOb+/mYcD4f+gY+r
n7/YcgO6oS4OYMGRo8O9PSt7OdkmEZUjD7MvYbx5RvZ999fieq1C26ZsPTNjxJ9MCTLIRvn2pHLy
r0EonXh7DMs6NM3mYVPDZNBEQz3d2H6IZAiIDJ/zzMe1uO3tYBeKj8iLgCI3TTyJuoICXzdTxknx
D7Ju1jdaRGRCdKLbonMpjuzuA5ezK3Zyvv5hUGizCUFjR4SgNMiNCHUZQX8FmcA3rZ0Sp6rrlIVh
j2paXG7TQHmxU+4fNMNLWtybiGQoRuk9axfK8dtXmm5CDjAoYY5TgcwoDl+GSwJldI4C9uAlTjCW
pIvCoARREnhsad0SMWXqVRxFKNkiZ0iO73bX/646LhRrjj6qcaj5jS7+GpiA+haQQYA3bk3Q+fCb
Yd80KA1HJt0F9kX0M6JDZzv2R0SJWERdgt2z0U4kTEqII09Ify3oEV8BienURt79usdh/qXDrttq
ows1nq095Ey2ShmgmLl8vZWCGSqhxdnxyCSGGceMo/Oo3k8adQy6ximgAbLWYQK5rsXqvcguGzf8
OPwX5uZbSLie00DocNjNmEs8czCoj8tvDJZRYSJ1OYpb+punDjgEQm0g26YzwC7Di4W2UhDrd1ps
NaNIBIDHt6cuZvtN+yaF0USgTiCtSkhls359ta1BrOX4faM95Frv3k3ifB4nEnpzhaqcFMshFlCI
zmK07LEonGYUJfp4bCF1KtA4PfkG4tnUEj8Q7Wc9V9Y/nRL/Kt/FVQCArDLMfCc0yZcOuWPhwHKn
5YverUbe9QCx8445IM4IaqP7xOKf3Hc9zuAMLVVdvH1g64w+uQoY5cM4bcRbGFuHDPc1FZjwh2Y5
5SyWGVeHUtljj0VqYCW/hjHZqjCzlwTqKkh4TN0W2cXlxE722zFiMiXY7+34MDPxmeJPvZ46xxym
smR1S3wZkhkIhrmozXswzLZ1m/l58sXts6mmd8cEB02Y/A0SS+j1riPqx9qXwICVq69SKf4fQeIy
i0TTJwXpGhS4rMtXcMJ2m6Au4XV//vVXX3fTedSlrL+GzWNZEH3r71UsYxNz1J7c+0tJjnnBsB8K
eyP2Wfl2LSpJri8yxJsK9Vpjk//ggSFpScVVdCKwv48dDDnQVziXLLGwB1sQ8xMjrEazHcRDtOhT
33WXujGJUizEFPCCqiqlmTe5zcZoN4T9Tre4FHmf8ak6UIMAXGLfxyZb2g6URBdDi7FuWQwUc4/D
uVGsTwNIwyggkHFWXZGlac5FbUPHEKnQHn0FSUmISYDdpFp4nf2o+AQ9+ZOcKvsq7jCMXZOOPQPX
Fzf/q0P7XN3Lz2wtbdimNUzssDPYK7Sn0dZA5J2iNB96A9bjJTIODmy91Q/Pb1bajqEuu0lTTnva
jpHmXFga+8U1cHiHd5JgNksdv9gf2uWF3GqI25P8mhhgD3oZNQpxrYGautGOVnxAjhKn/DN7zXqo
lvm+WIncQXEaSYkHAt5OKR0CIlutksxrVHWvgnZ0pEBOZOhuXfHPpF2/QvjnfOAPG6Qw6SlrEqIA
1JoqmppclY1xjGVhwXdzai86DrXlcRdhNuaTyEDHA83qEz/FHj+HDu9jqVr5c+Azy3xesHHi/8OS
G0KNcgzmck81jV6QHEnhELDQ1T+MuX+MaFCA6Z3IGiTtXLp7mYv+CprQoTwb527vG26CWuTSMJfj
ATACUwE4oXkh8H0fCugN3JNigs2SY8Y9i+Z0r4jJrpSMKOVIf0WghKUHtpWUe0kC0kP4/px/f8dp
IYmm9JsWKhUnfVh/1gtavGNGN2Xf2QWP2fWvUEboT94EG2ThZ4VTt24FQ8v7wKcFWQFFcctTKSC3
vrcxxCDgtoXVOyC6M27XKs9hgZhyeBWjpbHZQa2RP74dfEYE1lrCj3Hw4iNy3ZG7i8Xqy8NhgXXg
i4vem7exy+bNcdpjSrRY0cSZCytTRZKBxgMaVBl0fGWzvAx+3QIbkagV8OGQaNRcNpSOpiwRDN7P
poDmQc2+A9zrT083kifN99u4Bukbv7zl/vcFUsrXEKGAxOpTq3z5M2+NLyWnx2nWmq7DFEb2RI2r
ygRsX2F23mEnSXOcE/JJriMMcCSe4weiX5cHnfZEwEWscxTyzHpscpcWVNeTPS7qzUk0ih/vTmjF
BLKPSqf8PXF/OQMxmSZ+Ht531DMGoksIWRA29CGIAyRz9HJaU8bNK+0roGR/yyVvH6BD4NHmqo6h
WxegYW+c/ExKZiuIRvxTOIgLN1RXT0Uy7eOw07kepxkaQypWIcF/mQy5GGaPlxXD0j1iQm8ldOzg
SEigpBReC6CKyukcwRoPa7lnw6O6CRYoCKPiHsI4SxfJIt2Luzsj4WOZ1sU5mG+Q7kdoPedWCTlV
Nd/qSFDIw41uJLCGYawjIDawjiFYQW2MeVjnoPpY0LZICfnL1u0RfntS4+4TnUdKRx0OPvbfF6Iw
iUaAanx/+deUqyhYWiGVEz7di52OC2Ks5KAAqvC/a88z9SQLoSfjPbJKDkAEQai7t0LB3oVnioel
g1qwx0vuIpCg/akj62V+pPofg1mfEggsfH6Jl522eMYR9Sk1fha9JqngRqYIF9wrxnCkyGDyQhZ3
M+7uxSqJ4RD19eEW2dlxDE5Smx2E9xbtOgvW0MtX7DkTvWROQ6Jr/OOHwZIIrPajXY10emCcwA8h
SsVhmy94A9T54neIFlmJbLPB0G+NWZ2pvXd6VHHBPKfEBUnPI0Esaj9Hz9hTZGnldcpF8hNSoHAq
UmmTeG4HS2hjZUjbxdF2vxRHlvjDc7p2FGyjL5NrwTLr2t+r8pkseEUDWWFHdbAxZL2gkMHmt3nt
QXu9K0m5YtsOK7AYuyiALOpwmqZLoM1KafNwY6CAawYHKR/U4ivS7vh0rYR0LkRpK2UPpTpSKCQ/
/bTPs3R4PQmy6+qleirjv2x85XmESNf0UEOcqdLWycY9dO6qxDmItrCjCkQk7TFmWSJpCZGJ3q3x
JneJzKUvchdT3Rs45SkKNNk6azEETOJmjccqcFDy+TGEPNaNn5Y+gTj/NbyUVLvzQ/ZGvD0wnOfK
TVV8P+LFDpwMuB0b/Wvg0AMm40sXF9DgpWgEnfrC41Si2GojVlKI/9bnYOInd8LKqV2ba1embzV+
eddWQaDnr5r7tk6kPR2DxyCmdUkWcIZx6hSHggikG38P2KnPmti7Lt8HjHV29qK9LjNmdMfLC1yW
s5WnxpsIhr3OPbThHAx+CzEgSaTBWeMXKopTpstDxLeHilZ9ndxwVJpv6tNd6qRceKyqRHW3EOVC
M1w/ex0ZGg7l7Hlkj/WX0tvKxkmHptAhqEKF/XN3Jsk7RtpJn9ysPyWD+6oC5/RSqihFZ6oDegKx
sT36cEwfMFwViqZ9cV6gLkilRFHNP6VLEIoNAGYVDVJY4qqd4AO2hzK+yM9UtqBcfFSfb9e3TdaH
LjIKSoMVc1rBMH4Vz9dwY9cGTvo8NktnJvG/yXJVsDAKEWkGqAQDbT5XobKG2yotWT4WpI7FkE6z
QG7N1I+F4hEltwB0x48hkeW27ZPR1OJGbfPH/buH1BYxKgjjLYNV4NWFd+Gd3wCu0Ujr9fxnQV8b
SYGJxPN7qFU5ggBjLQTvSB14PLGW6EFLBvMh+AS+731IEwdlkNV5DkXYuFuNuKAyA+EHshqAkAAF
0zVhgUhQwgHY7ApN1C2VBuOUf0DQRYylC/Xgq1wMZiDveUGCPiWczPRifpLAPJStSDyARy7gthVW
gsCBrh5IrjLt1IePFRl4DaDMGA2RLBkdVj/o6rkcU4au5HLUYnIixBJOPEwr8/Hwa7IOQYVouLTy
4SaSHyWys6Sq0AOHxk1jsam+phSAtDr41z7hZTpXS4VNcP3g2YjldNLYEfgrMw5PCvmqqxMqXh0Z
tjHqMHWxGutDSJxeLb5Tf+u5CyCQQxLkh/ne/QhX7veWVaQkn9uJMBVkE4av9QJc0g4Oe5SLpaVI
w3fxfvfcu9z6hjwXLNWsB76uz88iRwD+hJXDA0Lbx9krs4LTSf7rs6XzTQl75Cr3K7UWYjnYtRJP
DQEutt7+1iYs3Hi3WMHlLZPjR6KQpSJTcjk4G1iWmnXpBhSKhFktBTBT+N5E11EEaMcaU0xi1miZ
iZ81SGyRasdhHIR2WmdENZGuK0G7nLTVmxdEFanBl9+t4T/8ZA+TRkCzcS/42k0f5/yXCWFN11kk
+hsjKzGkTyrpDSi7f/dAKiXD/uxFJjIytYSBzEGs3YDa5oJ0P1GLGArQV6EGo60UVLrzt05nVhr1
amm7PGk4jZz6ErlxgRyTHdyIqcHWMW0H6yaD5gKZ21EFVlyeTvZEjOH02dZpu5Lbfx2EBSMW2evC
thq529f2vsa6wWR3ty31jYTz7IN3zIUsJqfYea9kA+7Y0hDrvVXbnuxU6ucWEqsp2ijexUyVEKWF
KShKo05o+aMjmw9OaO5KMAcrjapwejHjwRmJmj0Wg1UvaVtvgH9x/DB92IvYSHKcyzPMr+cHTn/J
belfQu8W8dUR+PTVTqAi8EJcqmELOt2FpVx47AJymFsrjAtaXi4sadZuuA08DdeFFZkO3HFt9ngz
1a/1tbAEbBCxtMCSVf25CvaJmueohxtmNqw0qWlFnlBkf0QQWjlkLIVeqHqmnNRYmcmXajtTrR2X
H0s9zeJxhqi8GJJxiI9OOWbOofpivdsIRwZJ9yAqf1YlWNH8pSjrNU3xuwMuXOstg9kW+9dEejpk
ZiKbSbwkTX//3j2d7mOoyfstyTC6jWqgnivnFSofuDL8UYxppx1Ro74UY1JeHjbhV5At/Xf8B07h
vLDbttaJ9L/l5ZaO4rAZdCqJk+vlrZZtEtADXJJ53hhXmePR+bdc0V3a+GelDmS/iu+FXUcv+mdl
TXrP/REaE8LUwLQKlfxabbLpriYcLrJEV0pOFA547Td6rP0IN5bqaGjqb+D/3KgSQY2x9o3n7gtJ
xkgxz8oYLgLyokhiK/rkP0D/Q+Ygstxz62Ha0b6UJ1HW2v9XuOGzlHM1NisKeR5dWlH3/UsYnH0m
CjWy1GuXyRJf0O1pUZDqac9hHcGdNn9svnC98f4Ep2iYt3/AsuwGQ3PmdYtll8p44MxeIBUrACQa
o7WOr0VPWTpFxyDfJrwxew/gORhTMGv49nZZdCQ7YI8ZIsKk3JdBheYQZaEeWA3RJMnfDBqQzY0W
IaOg+z7wSSMefmEFJ+zv/L57UN36M+tQmYQBnNYIFpBO3ln0r4CL6/Ar7BAjNMYuBwncdbqLHlwW
eYNKmCC3CVBb3MSqu/YZ8SCuQ2f5xdZhWgvE854s6dUKC1cBlIqj2W7RxMXu4TtBSHrXS83qHiLc
sVyZHqy4mVpj9tDi2a88xa27n2UNoMwVJqOOvDYL6AC7pTeM/fSexR6NNqz/Ax4x9Pa/bbjZbjMs
wm4U/DFCT/jSIxsUCUBKpGfv+1sKorlhSMWdma1d8kl2Og6YODa5TD/k6yj8dkrf2t4YoZO2p7Ki
RbOOeWAitRGP8scY0BZuWBw2puvWCOQPFCC3LcdVsTYUErDtteer2basiuXOSLGussisK0K50oTX
t3YUm2x4q6KVKmLoPGidr58MYZeGNLBhUB9LBBqcL+duuoDCiZdRsjjGC2n0dEn5Lu4Ke379AX7k
KoVCe9d8Cwa6CvdMhm1K7XPPmfqA60HuxhqC5fhujqLqvqZV5Q8rT++/y4Aqi2fZsBCqX8HhGQQI
oCOKOkEfjZJhKZUp6gq9S6Z1ngkBH59vITHpahbXQVp1kmwCn0AdFYP+KK14dI9NqecRlEJkw32z
26IRVhimzAoMMK7X+ShWmpIGzJYnF6GE4J0kqIjESAygDKSdnWbQ4DGLkplzpZmp4xPXAV9lpgWd
Lt1AswxS0w14nO4gK7Dhin+msE3btU8kDaaTA04B4o0asZlJhyRf2cOT6LMmC1GsuLI4YUMUSyfn
WVt9aynwhS1PI9S28bsh11PBDNXzM0cO5DxXgablLM67oFm0NbiipSteCq/+KTpOCMvFfA76iweA
e0Ul+rrmX+/zBOWMp5pgvN3ez9SS0grMo4xpUfuh9LE+Sc5BXLW0Fdhcm6Pww2hCOdCysI2o1KxF
I1zvKiuiZVtPIYwYiEq0dpX7XyFn6kMkoK6d222faQrDfwOR02japr0DM7dWFfaSVY4/6U79fkyx
PayJASpOdZdUGz+DRBcnFbg+jf2Xc/WuzJE4lNnaAYIs4ECMBTwd6W16VvzpJf9MWgqGn2tVWG2B
1ZxgzXOmf0Ru+hgGpIK/nd4Dfqexx5dlZGDzxVfCpRvLkKsQLilrCadljU4oSc8ixR32baS/xFbT
3mz8BozT/ljeK3KOmgcX1DqGPyo6XxHLJpEckIUsOwMpzQoTU3Lxa7aHdKPNWvQMZteEs7PCu5C6
r8sRsqS0rJMS4iLgbB0I+A1O4duoq27fUYXLSJI3wFko3rNdh5uazEo+cCaH23KqdSudAViE375y
cxx+GYR7EoGNK15QvtGhucY5fjAeCzW5ZrEFIyy10fY7+S5ARsu22Ta3W8OF40xYUn2oeBRaFbvc
C+W+yb5xX7pZL/nFJdbutQs0WvniJnnDrXmMlXSWSnSaGJyXwUbxYcjKvNmxYxOM4bUZFKtU6t1S
iZElwVcfACekbyZnkpqunG//lpQKcQrknroosyVttXbroBbLYPuZ6Q8hzNTVH/jS280pA8NdzX+o
wrZshhcUoLn0j32QXAOubYvXHEQ38l2WEFzYliluGHHiE/K5k45j2nkTn/7jOyqL7SFWfW4wz1fM
npiT86bf8oIwFU1CYd2OmzVFRDqpRGv3vHqfvZrvLQqeQ7FyXrxB0gI/UwvwTUJVcQAqDi/tBHVv
jGKoJ0Jbe4ZjgQoJTk6bsS5clxN9Ow/tL5PK41j105/0+ZTLvOwtOUDn8qK53rmGGVGdeR0Blm0u
uoU263abw3DXLSd+fcOC4Ex/LGhTqz0LSZNAeFGCqLdXhfob4edjDAfR+T+g8VQkukTGAQxxtOJ6
si3ogky7fXSliMltCBtw1HPGP/ExYZ2hl6u+GSxjK9ZpRHmI+Dx+df7yuEJW4A19Y0u5aDApNnym
S6oCh1y36g0fi8pyEPUwjR751Zeo0vp5XWWL0Y2RqjJPAB1BxQRD3zNNTRVuqh0j27NqgeqgLQro
o0M+q7/fwdOIAM3PXxWOWoXEgL6r1wFoZ3qpkGi3TlBfKXlLhhcaseULoxqD7MSQKyrJH4vPOXr1
LR0JEXlPzbfUODBwwBsVgsDU+hU/PPNT1ToANM9Z5gbr/8z96ForALzxlt9d3lcJwJQFJu5v+EWH
CABMB9G/QBjqnw5tpz16i8njPAeh9U9IDSghvli3fXhwEpE5k7WomUE7NLq3Gto+BMiO5SgNxUNl
JBJF66jRyv6IvIMw1JcjQ2TZcFGMA5jUhOOvCQDClNvuzqidwamVZILHLPz0Kkl6J9tsPqPVsP6i
JQlMU4DWrVh2qSwZWDYR4C5FEuhzrWGXwfAN6G2EKff9gHi7rxe1i1x4euGxeju4UHHWrbVkOKY/
1BH19OpgUkLSfShbGryizFxNVcsCAfPeL8xXF5JJxGqiJs+5om2OtI5hcrqaETsFRTqf/N2CejJN
gyPNn7w6y17eGanGM/SGFzXDijyFjVip+m2wKOECYfjWFyHoe4sEzUt1gglBdtcXwMsHBk1WytfZ
jUyAJe9j2xBRioln7lzrQKU+8nOO8RMhcWjGUNNgBH3doky3lRSq8knVmkGj0ZAt6kDaYgf+D+oC
xpLp4CqErNVG6iU0fR6CMqp8PLeHjON0QY1ucQpDvrX3qoeC4TPQdDlA4jZPmH1uHcXD5SNt5Ewj
vdsOIedKlUngOiuMULXbCwF/wwcJsq7XEuwnqZT1UVNRjjshEGGwibbyF20OVCA+CmhpmVfT67hu
V1x8dZzmzthRTHarklVgwNi010k0JY1JpHlwEMCs6q44wglBmeu7XTMOIIa8vK/cj4IPYTxGZRzZ
KQ2j+I79hfB/IcbRu6FkyTSYL9tjQgJkJZc4zUQKbUADC4TvJ2i+n3wQKmK+ZXOe851635FG7g2c
WZn9a1y8Mjh+DjjezfgHsy8PY5G/lU1ks0Pw315nceugdgBXRKI6ZgbjQzkxdncMp1QJDMN557ot
W+FALSsNvMZhHUMaCJu3SQJd8aDCcPzm7V4gxRb7hR6+pnOrvQAXNxSLGzoux1OX3+jqqx+C74uJ
9byP6QP9UPT41kZzHeV3JVgC3eUL3gMEQhpXiNIdYq8RhZ3GlFEcOq1LVpPyXoIyRj8QfHHXwhKZ
pewzyqH7SNTfuSrUQwp50IBEAtDPrmdQKdzs/qZu2raC5pnHs5/6SSNtgj74AZM5doOk0mMjnFUD
U+oLnB8n9p4y0WZGSZSWJytj0gTys6iXcAyFHByzhNUeT3p/8LqeVAOZ5pPpahPQMfMtfs0gkPGm
L5ll8Qtdde7ymP25+dtONOLa2y8CcLiH+OTCtzqsGJqHs4bWcPeNuQD5OIKT+iIuu6FNA1l0GLN7
6ZALAT2L2WfU6sG/Dl6YVKs0ODXVH9ROxxwNobq/eE2xIQASAGBifKB85GWWSDCIULdPtzd3kBRb
QdXBIiFoKhME1ZX8W0NMRj3mqwR5HKd+6zZQWJpggn/Z0Dp7JYOllwaFosRsRtGSd3vk96Ib4ZaZ
4PwDeTjMKCmbxqt8hXtPhm6r0qE7f5e6RvHg2sX+tULsCO126v0vj+teXnv9fTpdgct3gKSLXvRr
LkHsOfW3n7qVLOiRf3T6Nopu6FK5+cx0ygf/d3ILpMnO0Xm18S3LbaYc/XQe99M7sD8caEqVrQGW
xh2c1nSbXm8r/XhMFOVJ+leFfJNS5gBL3DHzHXsc7RDZVnEeeneLIPeqmzn/izA2CUxj8XaUDYQB
BrF8p8kdmhUGTlksMDbP6SAQ/ZG/Sax+f6R6T2hqJuvQZ2B/YH5ls44saeLEEbjKFQoLCrfRAsxx
hBRiJ8hvvZcTWSylYUDio17vlzY8V/ZsuwuXdxYpkcWauMs8hKtr/uABY4OAz+rDhiXklyV9dEGM
aV4y8WlobgbHub505arYmoJEOAjaUuBNyEecwdR3aeEFvK9YNy0RQU6nFZOGmNba/CW3taS6H455
wr/dr42beJfAM/sXQNXr+WDm65hTRNA9osVfpzRsKI1IY7q8exrd80WyztAFTzjyp/j6tvmjFXVl
zMiHxS5MFpcfE0MxhZD8JSPg2aofsg+kV4Se52vi6VQTU/Yercz7pr8qhBXqkBWmwGSJqZfJcJ3+
CVHotGLWAnDnAaq9uXbY2yIt4MEfhCSfRV9+UNzJh3ZtDxqwEcGuvc9dGj+5KG3bSQCjWZxnt3FB
Dd5P88EZavqaCdqDbh7vLM+4sUXbVr0OtX3D9luU7Yb9UEm3RC8ZCDVVXN/LpIefDJ6vDN4YS+lw
qAnw/G5gKhgPiJP2lNbRbvj6OCqrc4S1GPX4fXKJKdbTcZR+8mcJNBp67CmV+yMFMgpz799QKaPi
QGYNLwwgt5z1mr+knZfArqNGdNs9e2UV385r1ojy8RWv6ELhhChzccASKCXybWBt/mus2Nji8ACB
zIyeKqddaon4F+IWOw140g+5GHMe057eEEQGm5IHzxZCaPFa6eEnUOKhoDKbHvUnPLbwteoP7paZ
DzRWTogUk/52NatPIRbR0zpb4mFMk8UG8XJA6T4v32ES77CLy05/CcOfHQWD/fCIvK2yu+Lefm0t
dgnfQ/a9sa9/9l6sTOjYmVoo27AoVL6eYlRCpxEJZMFPsPaPKsyCst5FYMumRrZKr9RwEng35jHI
h8SQ7WzJCMlklP7jXgdKosf8HD5maAKRyhiE7p23lX+8T1Yva529PldcLA7Tj049KrEtWA1t6vgl
4We6z118hQlugmemgLwH18ae2u7ZapQVBO0jLvCXs0uGOKotY9LSLZUm8LHSpZ3mQ3Ho4fqWZgkn
uwgA/0uROuH6G+karBpYbEOmdhpVsqsCpxQUDy6fGJIzSsse9evBeAQoNFnbotyDmUWlFLmLTJYM
9BAl7n4bEjwMIByxjUJm0inrbVUOIT0ZWqJnYRXB8vAtiyBconXuzGpZ7R5T6fpm5IEJoVhHiCUE
sIIzhATiJlsicG+ua4cTv6vzGU00PLolS13bJXlRo9NSLnac2yHozzuhZGO/Yvmn/KRTyPGVSn1L
y/fcJ/2yQDXvArcKz/kqb/3FdR1rkiWZdBsZU2sqOLAe9GJeum9M8pF3072JFe2uo+I7R3jeDpxo
3HIOuv323N6OFOS/CKJUmA7L/9bYmNsryAqCx/v/t7CTXdUToYG/afrzh/q3L4Q0jqOD1/gv/Rqh
mDciI51FW4InJOesE6tPO6pXCrqQ5pEHkO7mWQnwS1smnHq5PIAFLLdxcFtBrZdl2hJ8tTaqvkPe
gSRwvN+Gwyme6Z6W7j1ezDktlbA1zx3T66sglgTzT2RskBXlMhdRcFZ+YJVBfB8dqJ9DMRT/lH/G
jtCI9E7q2b530eEGJi3J3PamWQJONiRNchN9jgpsqy++XWTYHv5WASwAx5ANu8vDFSHVJPxNXr8+
n43b9oCYT/Oni96e9cxdGNdv3ySfVgkjVx3ONqP2oJqhcK3rQn5bxW914BbA3HPC/TueeqBftPC+
EAPQntExze1Cr2VJGOyKZsTZy0i0GuXH1F8ZaLd5JImfLukCbMetrCOz2ShFhCeMQdqXfh7zw7o/
Cv0/No72JfR0vchlX65Kmt6aMt5pdhfoqr7aX984DcKp1oFXfqmFJGXOGNCGQ0EQ1M+XLwypXCrD
04IWd83Hpv06gg2Xeg0eoR0cdqArbOCsYcY02IwJwAwr3kB+Mvm0UUs2QwzQyolmyDIbAegxTOxZ
6Bs+gzPJghAWYpDJfO6KvsbKVgJshA3p5w+z0VS+Gs9jaKVsI4fQkvFO/LjptKscCXjs66y0sCuB
YBmO5D0EabR8PyY+wn0WOAMmx7KW0YRFtcQe+8R6iBQ3Dr8FRy0objqMD/eGpLQvaXBUZ/M8eAPV
mzhoUxg9XYlLvesciYjQBLRip54rRgq6r/iHRGgz8VN+pXS6i2Rvc0FZ1WmGG+aAx1168suunwaP
dbEph6EYiRPSwEfycbKXD5Gplej8i8m1eaOBQwauKCfOeCoAZxuAQjoE/8SSIxY7Qko3P+BKreGY
kWWyDObajaeIoa+cyOVSKfUp5+lIO0YWj6wJlorH0p/Smg1uqnEOhrlXFCaxVbLWbJuyusTnMWWU
QQ2Z0CtiTp8ZKDNbjKMBfozJr61em3FvXB1s4uK2FG12vSnORWcY6NuXe2ClXGpGZL6S9T8J7Hu9
YylEKt/32eozhKFi25ZGSWaHB9oCZQ0jurXKLxwqCy35nxmx2uXjEVKN2R62XRB0fCgkFqteN/cj
JtMMA96sG4yUcJzXLNIfhrHId5pDygMgWM19uhaySjp8GleML51mfRvJVfxn9CHTpBHDXHoy8HOP
FBWgHC+fX/66fVacE+6CRtWnf2sX3GoSct6R03FCsxwn4VywwzaG3r72gnGPyq6gDuVQOdw0zeCC
uz7+2J1J6ivuHoLUI04BkCG0HKJjWckFb8ssZFPc7LJSshkkQi6cBc7uNw45OyQM1JuFdyhTk/H5
GQ7q11p1QBKL8136t00qvS+QmFQ+9aUZ1W/Sz1VQRkYq+vZ3QqZdr+pcMZNwSvJMw8lmdo3m+yjY
W7AadOihU1qrTA6MnyETHJb2D6F170hEaLYrGpWYh+kJ1BFhTyz//2GxeWFqXKF4UxcrjWnPrwy3
Z/o8ae7L/TMDoJAM9kUE/y/2uCH1y7P6iKrv7YDx4og4h+CrVY9JdTASLSqKRlLNDwud7CiXgOSS
PcExyK+5IxgnMeLECznpItYMPUcXetmC3xZP7yMMiDWKU2XYIKoNDd/y4s+mv583rVjgdCDJOeqq
WsUJAak82EBmuRB7C9fwA+8hGaEKdmeWP1EPVkZyGQN3zx9hkiZxtURRE/ekVQQ2FK5+ZH02LBTJ
yQzwiKFaCPNwtuCG8kMqzSNDROmtS/+X+tR95sKu3sPNcDzJaNge+ChQbrWZFZFIhL5GBCKOpY4d
pN2Q7McsYAx+NLJn30OFhlpfoL2zJ/Esx2sXg57+6/e+PvoUqDsxw8hWnwu8FtLafKPvxnNuzeFM
vSbtNPWRWzOpcmRgXJw1ewrqKAeKpwFQRXlC4imMyX3CEqE2ESjnjKlpRu6Zl555eRjMzGrnt2X0
u1clo/NP5wdywQ3j9NCwDwJeEywF6UhdI1OgiiHvmN1xjcSNJG+LJwGzh2oUUdtAiig2gSSYcoBk
suN9MRRp+mzkZmI7ELmfLVzBMtPLixl+OnmYYvK4J2RLJ6HeFzGil9HW1oXMw+BGn8C86dnHTXg+
3glmugwrl5XguZZRX0WSr0zEPHL4CbkGCjm7iaNisf0DhWq8YsqO417pO4ewW3plTRaXmgfqFdf9
ZVYRKkQlI8rjen0zsoy5UpTCyzWXIKK0b162VNiFPgtlrYsVf/Tfv2wWipSrJNbqqt66SNePGyiC
CXF46FcbK56EKHi/bHslRFmrzGlRuM/2MTc2XaueF/8Y1uW8omg+4HJNo4EYS+ONfOwbKaf6frqE
G4JAqr7l2ZT1hyktTD24aTZcaVMdDZw2NxboAPtIBSRSfudW8s1fYa5ZzXAfdDT7xcIoSX5GPtpU
L82z//mpXAgFUxcOJnSO+O9Bs4TfosAs4azEby9xHsS4ZsVRK0m0g2F9Ez8mB5awwYekCEhMP2Rw
gBzr3x4qASMsj50lP7WwbhW/XDr3et4M7BmIYBMSH7cZOOitxTCzKNhydi1tN6P1cqbsvLK6FulG
mAQf46mkymG1T8tqGISZGRX8+lXBS1u3vmyjobKRGmZyFvY3JSkilDW7U0JacWgaj858DU4wZmC3
+fsFew5HGGfwCfQoGRqfssUI8p+9in7BNqiiXgDLPyfJ1+PmDHYc2L0tzwbbUP5bcV7Whu9zsucD
ICnglNhL2WBMaX1WhPbesLB6Ex1CeMQKk8bf1XuN2Iv6eed46la2YsfSeP4mR5y+W83ygvPrIJ/x
1TCpFjyhONDfafPqSACVUrw358ypPw5AA04Shvh3hChdtKLnSKz+/eaPBkYHsqyzvlPMWR3z6ycd
jhJ7ACJNDWENAPB7Arq7Hwoh0vc0NJ1U12lkNdVyTJezw1JZNjoUFLHUgHKIDjf94qvxoVJWTu+k
nc7hv7siwouVIjrHgFgRd1/hCCIEGBAwdpz1qNd/9TQ8pHoNXEUkeT6bTVA7Kw6wvzXqKmNrrhYB
Cy/RNhupXabSVBh44QJ0OxUo+vdsl7A19Zthxer9Hv5Y8SHcbdvcKcStkJowkwH36xMUoEBKeaap
q9xjLA17BUogWmzlf4ceaLBNXAt9BfGAtKgJ3CeubwiZ6vmGafA6IbYZOzU6kZ3MOBypG1K6TxR1
HygsyuYrsdMWR2aaJAAY3QIA61xwDurmB5Aba/dwexV0f/+TvtVos3gIKfXgixWOHPrwX8X0j77w
7gb4pbEo0H4mFZV6MjpWAL8cHqIa4O7TV7aw79QoeuiUWYjFj+K1PtaWkJ/ahFfQgBgMNM1nj8+M
rqKCYEnLFzieZNmLq+m4o74VRfRgDJxxUx0nzLyGWs04cuL7wbPDiPLWZbmMNiqwPBY1Qb+VG8iD
eEH0umcUbidGVtAaOSod0K+LIlHkw+HB+P6ZyvYIjVaBjuocqk79tYNJwuLA9BwpihXZCyB9DX0a
xNFD5RIPvlKfs+dCCEB+5sS3QEwdaSCUtOb8s6WrVx7SRFpUAhZQ6cqsQosxBNOeLwpTCzBsQILN
TZgGLC2SlW1MCgP+L1VVLwvzql2AtSS1IrY20bUm11y/63uM2Gj+I+FbbLqKF+4qDLf06cjlMq2q
XltmaMqQ834iJmejm74iCPNmABQj44r+x1o23xmPOPYH23jqutGMRDjnUriA0lPe922YBDBRW4/+
pejwr/bGNYYXc+ypvust7DqTaex+NVBI+Bk2ZVwv5mZL4bOXB0BD3pk8kYFC+3xlWhoLssNVxp4W
9qMql7t94QWFqE4PGIcIZ1b1q+RfVE2xrPXyqJ2XLfVj5ApDFIMUE6XfJTSVmaCZHihDgGXy0kuM
RA4ya8rlMVTXiy9p+w+7VijdSGV2+fRjcq4ERDJ7bHOO/uBOXh+aPAv3L8au/HHKh/Zbl6WijE3T
lFT9tFAUIMbaImLyOyZ/FrYmf4KZT9SFAl15sBVxyAZ9TQORiwpkb94PWEdsbkt4mgzGpuUhdbpP
f2ezyonl82d9XL4/hI8z30PUQvkFb1+AVp/CbdNDYAnMUN+ONnAIDhjfm691XtmGS9M3In2Cc6lp
pkao0xkmOUKeA4g2qmJ0Zbp8JKPNh7lPb0zdfEUN2LF6kX2OrfJPXdefnlgedOMpVBvO+k7FmoUF
P8GxUeSUrKoCU1c7AIxfrny5niO05jrpgoGSsA/QraJOmL/WdOlaAY5R/m/MvrHPcdmNr0+CqxYm
d6HdepTRCRQJKv26uidqGCM8GomGVArD+MUkajsYXnhALy8v4Mcmg/eSwCvBhYqAjjGx6dZxEGul
xvoqr4vyq+1NYtR+wP7HRacJHKTNchrIRJjiO9Fn71Ka1CCHeHZJvSLGZivdsGDAbfe6B6q6gR/X
HFn5EetNwNY3WkPcWscaVpOoUE1s+doTQJ98ZNiQNBqwy2e7ohaktmLMxsgZBenIox3FB8It9IMA
ljelkCDAR72Sd4WAScEO2V0lk0ki9oXF428b7oRkqIBpBNZrCec2Vqi9nEzU2zbk+O2KBJsIQ2LE
DmYDEsYcTALKkvp9cmVyyn+w5k0UCZvgVqXXIG5cWhtDedemhE92cQlP0+/8XjWd5rpDqg1nVTZO
CSp7gikKTp5UEyRQRYuoQycYzJPoWs6983bJN1lTNL6Ws9qu8Jh3WzS/xOHP5XFsUNUyHlLjibmQ
NC0JWvytqwTAo7hWHjOObp18QOfm8/4E8uEcgnzmbuUNIO06IpvmUXRXI3sWKjBd8pL4dUJu4A3l
KcVdgIZumuZA//xsyN4XFvWXFNXrQQ6h/L83+C3xyfEmbWUIXH/1/IQjz+Dt4QOw/1CfUtYYDFfn
lNe5JuRG/qej06O9kR1zg2v1Q5nSd+pkRyOMVFP+qFEU/GEeELBWar3lq5VPpa0DyeiClejHHos3
SP0Zzuk5GaSkKrK6eQJA+QWhBTxTo2obaazX0RRan9EIdEA9oB7kqUZX6YNIqQKY6WC+IirlOV+o
GD5A3vqoUlYvuVdtx7FBk/ilQiXDUQ31cjipgaso1pTiRsToJo++5BuTdj9INoPL8mXI/KbTGtfK
LGTheT2reUZWHoE45dMvzsEA1WXuWK6gf+yQo0gt7One+mBjKQvnStrBIgbKtRxFg5PMJ30genyh
BADIHLZUm87YzcNWByXIvNv8jSzIjdD2OQHykSNu1lRLH6eVRcK/u30EyGSINhxcMAhFSJwbqZIh
lAqKOKACsbCKoEZT8EqKT0DxxQdP+dSutBzIamllkBANFzO7xTV1aAsVQVUcIt/Kil/QRx8JMsPW
92jmotBNQT8R3N5r1ciVakAc/DQE6+1E9TDOQG3pT/+/j1518DFs7/+M8EkHr/yX/7Az/+N9BRzA
5yshluK7iLzvVimol20LFV2aQ27Rucm0wns/pHevY98PQH2LQw2bYX7kvEjAHF+KPr+DsUJhMDzK
Qjm9MlMLFMQHAjZ2DYzZLZKxoUE3T0x5QAVrG2rFlQbYL3Ubgd3IC6jStQ37LZlBnXGxVsyA+tcW
YBldL2v1GyjxR52Ou2My68FGIVzlOUx3Jb2XuZXz04Va2pitzQk12d0pmGUNzBmG33N+8Kq1iNT7
yhwRgHxOmZ/ri8GuUgS/QM731+18G9eLgkKzRVSNe8q94PDxsmqbqUv0+xguAs6EOYFl2h5MDYEx
OO1chSUIWDj3tBsbVQhVV7SKA9nJl064eVS4KK4xGCPq2mIvkhdHJvuk7KkssrjwveIVQc7a8mhZ
gd5W90Kxct5KTB5dMu4B+k8+/iZDHKzvZg/23I+84I2ZizlgF1FPJE6GtEb5VLQYSQYqVvmnQ8ms
ey95BNbyEoexDPgbgRW5GWpmeZtdIHXb67K1BisgWN+Hjjh1ohW5dboBbBqonzp0MXZTM3qm1dpu
t8oMI7dBU5D4c1ZaXATykKftKRtLu+THmL5+Lo58xe9uKrd9csSt4vSIbVIXEikJty9JG0aKo3Nu
aMy4AH9TT3Hufv+chYOvF7cTVrc6CUyt/KWTqHwcnCABew5rlWAE4dRoHNYanE4jges2o+tzIhSj
abv11U8E1RgrZfp5JUE09+5/Lej3zk9S/9UsMHs+TlsWx7mztxCjKKtUGwgKlavD7vxgY7t0KpRA
xwAjp2peSlNu6eC5XvEIWPAAtWEiKx7wbellXk3imF5H5QdDs7Tp73bKCg/NujYYan8CAkoxcpbJ
X1EE3DCsr2yP4qSf1AJmmhL1TqFn88kuUihFnoA0w+34M75Fd/9UpVCPpiLC6VTZ3JZDupFLHEc3
HgwVnrTG/YCvBSHpAOJUu24qKsnQJRvOHw8X/OAUd+DLswDKN/o0A9xgxQj3xdQStfM=
`protect end_protected

