

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
n6SxQ4cZpYT/ILbURpz0n7m3/CtPg7Srwf+5G6B92ASMc93ahDGfXsRmbxfQ4itjqNp4bImRWGHp
TxDOCQa4ZQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
T+03ThTlMB5LbidY7dBVWlYp0mNjkvlbypoxh4ls7n36ZTLkklcCR9ZkGKPsYI13rJYYLwxb8HQ9
lAxKeG9QmQNzwwKufgYFwBDRimvj8pMxUUa5UvV+Um8vyzZZSQmIWtsYrZE6EEbBovwAJw8AOtaR
U6gMXGczY3zuLvGCvAw=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
xyeO5Evu10M+3X2Afou0ntsX5ZB/pwkUmxi6MkSVEZEp/q8vhRIBXtucD3zi9CwKskciGYDIN3V0
Echz03lkOALKA28V6TwxpTDjOCcWnPUs+SbNU9hrNos5LOcUeyT/Umkuwxvon+y1+GmmTNBs/HsN
LDp012R0drMTXSZtr1fQtCR1xHLj1REwEGmrPANPbJm5g9t7g3uQ7e+eNRUcylifmDkL5SHkZMiP
o5a6WQY9gEml+rOEV7XkaZKFEUQnZO3nxTVqbYgCz7Fr3B2jvSfBBfXQPG0AKW9Iz7aUGng8TS33
LFSc4gt02mCKBH1NOkwuxP/U3rpVs0fnK6xENA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
UaJ6dwyNV7zPNxnKVFOwTBNM7GBgDixNLEFTEeGL4zxIus/wUjUkJRcBksOgUQrjesNLi9rSamfz
a+6oBrRU3NMz/a6LqvgLX0FtqLiIT69wj/tO+121sBluFxMRAbLYxwtNx0oswICZG6ot3kY7wUo8
MIP1BRyvBE7h7gUe8AY=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
iLkN9pn78C1qipOzfdJflxHJTY8JBXpf4rPYSCaQgqf5yt0IOulURCvwg0EGtXIXYL5OVuC8GGss
Cxal0AVlk6DQJUg5tnhgoani3XqnRusVYV7ivY3j4fNdUj8iyFUm29wArxnau/1wGXLQIbXlD+l5
Ze35HAoJRWjnvYyl2fMDrjYG0QtBEQHUh7moVIQ+kI8DwofjU8zFsu1KHGJsBje+80Fr1j2xEByY
nscMu+13hzF1cQaS+Ce+aroaWDuHJWx1kJ8/T+29qUQ8IgrJDtRVEWayMxcA9x6qrZ8JHoIeOcCa
xCl16mCCnpbqxuPBt6lvzV/n1cAzp3w9LmCffw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 87504)
`protect data_block
AXSDAAENmhT1DX2M+vt3A9dX7gzCi2qPK7U4THX9lKzy+8Nh60GU4BZWa8BySI9agr1740Dt6fXH
DMUh1czMgovyRsmAgPOSLTn6Eu0upibYlrMPCT6wh17vq03hcWCHdj3q7kre35aKko8NMINZ3juM
vMyPrlH2viSn6Z0UFMJQgIgPrH43cmJnM8Ce4/JMEj6gr/fmx9tcLYs1PTdZevRYM2KcF2G6hD6u
o3Y35wQcUSrfP3/zpSSZ/cfQ4df27DmqAFxlCPDOaoEPCbVdV2zIfzZ5X4gGa/bHosiyen4ElPTb
vPiT/WIMdts+wF/uXURX1dvPjLfvpKeL5bdo9+itgLLv2GgFMBhnVI50z0nfKCd9fwOLgLy4xUrO
pmlw9TNfGoVtsKrtBQKBUCsovQUvfd4La79c85nAyQJVSVWP9CX4uRqXq2f5O3N+V7OQEgT3V9fm
UD/VKzkxMesZjxLxQPvN9geSYar7BcBv2jiMs78OBWoFOCayz1FoqZIVm6691gAHQntMfzWsQmwz
F3hwbGwPdgdBSKh8lsUCwc/Fk4FpjXbKNCR3WvkF+PWv2qfqOnZ7Amt2+8HMEVjHouE0nN5EM9DG
x+b0Ph80vPZ97IbiLwpPlN2TWAl9XMJXWnd1Qta1uYsDVCqi99NaEa82CyuKOQ23bXLV5MgqbvTj
oCGZ80Op37rDXgVtTOZd0iugZPsG0Nxp5M5CJtqmJIEtpHm4iNc+7KPkKZz6GptDPm0PZBxAPUWe
5jN+I0/RO+C69kRmyCfj3RYrl9CX18iNvKF/r8TfIyAkHhWcvQioXrdcPxJoUq2ZB5aIgIWPXtiD
NDg8tULinaojw9bkccpvScMiN6ELOdqYGTS49SR3VyV5PeZS9I84SHmJ0T5u9MppUgBfvV3VnHO0
leRk8C6Cy1yV2N26zxzWxqE7vbaTf6LTBpkDKnb5fnF3cGLab6xojkulJ/9k3bRWH3RtJnpI5hI3
o3DtGiqL6OLq79t61JjMzNOZuIvV25L82sZnDul0Ys2SScaC6fq344xEluZUpX9NWLliqXy7rwjL
UErBL1JDdZXGR4/TmRAaTl4UUi9/TCv4W7eNuGS7F6V06ShCKW3KOZaoqHRPiefbT/5sak8qqC9O
1Q8QA2K3Wl0HPR722mXwJ/hlvclPynmOJuf9IcAJAeybAJ+j6X7p7uwppE1hVDdDbWMN5KrEBUgl
v7u7+5JbbtolcOHYGcq+/rraU4tp1Zta1zck9+vKN0CW/AAc43EMk/zy6P7TzYb74LiEPvndwAe1
0NuwTFhu3jg/kwGWT7FBPoHMeqT+PXBH2tWYRko5H8Hq47bF54iIU6N0YqXy7y2BxPqbvBL/YC2o
Outf9d1Fl6zkzeFFDM6fLokysKoiNzYSYOtU1LTGWee10s1lSCQVMWbV+VVOmz7lCbKiO2gAFdEn
JGTd4sFozyo340Gxsp/rMPDUkGxwLieICZUQD5jdK0HvG4gpuJ7DLCUdZymOGXigh05mHj1VLokw
BZDs0RJFooWJ1AGIDlOXL1axeJlkIWnSpMDdPUO8hs+flv4WU0Gj+iz5nOEW9yr8rfTxjTxc2e5A
syV2dxVyAvK4ya3moQOCSPOKJXelH3hConpQdBrahuQZ/dXIpQN1ZYHUec7EAXxtykYkqe++hYLR
PpiNT4s92dNXZ9Nwh7LFFve1aGYAybkCQf4tsbE04RoKQK6QuH0GHuGbCnmZ6aG+SFApibCUXro3
mD2VRwl0lMdg2Df9X7fGHQeX+b4En2cSfP5LVZV0m0A1ClMyFpDO5bLVKRs0hwFBrZjHSEhRtunW
wyQc1zlT6FDiaEDoZScMbUsAPAFKiKUbvJj7RC7bcOan5BwdSq2TOI1N22fSjB4H5s0CUIsSKEHM
HTf9AU7yya6cWDQRJBAQBQa9e/a7zcv43iNCBJfvSCy7l5WurIQ5OwVHPutUMeliX9oyuLZhg6/u
dLIDeQZ7zCsrSYn4wwyYAka2f/Mtse120GG6kNHxdcvWmS+jcIG+H077PlU9EmJIHfoB79ccad6E
Iao+eXfZ6oLAoPxQZO9rIZivyHy/CsOP4mSQ0v/xmNHJ2dHAFSnqYin6odvUSi5w8baqMz0EbOQQ
y+l5RfRBlnVNKfJuZsuK8dkGplY2uQxcjnd6uuXrK/0MrqDyRUTFrQlhlGW3RkcEECeV928Jmc3Y
x/9HqwJgNv2uJd7Ja1NWp2thA4Vn4X9qWM6glj9qltXkostO4Zzeti1NFHAqfVv5mJtpKe8bncoP
c/zmtTo4lCTTKUN3dtPSq+w2g6Ni92HxVbmFiKzLsaS8+t8MZLeKAEmaQopnLQq/4vEf66TRSrd4
p77w4UEy3J5aP898h1feMwp9fB1CvrD60eHlfgLiq5Q0kpjSkg9Ezek+uMz2HwjNg9U690qx4dPB
KKUXfnO74IbIpMxCMEYPlS5dvKQvWRRKQZ9Mjvc7aasooG466335SMMDzDC+ON+4rfNySfXZlTG2
+9UdEuwJgwQQ4ZkeZAkZ18Y+WkTCHVARrcl4BxdgbRFo76ULCIyzuVv9kOm9DVGAvtPYoUTXpMLk
5SQhJU8liXBpvJN4t03U4ObxuVPjXoDpyJk43mVUSQJZTcGrhSqz2rJyc4Vh5doNgX8gt6XMnXYx
Ais543vk6wxcOJz3qJ//C6xHgGaNdT7jfdSAvQJfzjfflXZMHrPen2/0RLJJkV8awOgJuxI9HnUq
aeHwyDosJ78kT5JyJf4cIpECWk7r/2D64O+srAL6JlxltEKB8MlrwfGlFjkfD+ShhdLnhrsaIdq4
9CDRwIlNj3xNYvvjJOe51ClElI5WSUNzoCBoeuXaF8Uq8lg304Q5bq64HpCIWxc/w4IdBZrRxzIS
8ZdxL4Mzg6K7r4u+1dZ2TsgHKs9305S0dhW9a1jNC0iAzhMc3I4Aor/cCH0ytCB6NnhNABMgDo6F
yDb9HNJHYt+tQBfBGI3MNKiAsWK+VMbUvVm6p6OElwTo/NMl3FIHXYTDLDaI6E95MjIKu6Bxsm2b
snTjybljbRoHhtFNMx0pP3+4oJ9eZc5XJStYwIqlvcPbQf3mI1rJANH3rjl/G0/taRZ+34f2+KUr
G1//10gny1DEz1Mgw6a2MQMAXOZ3az+nfjm3Vk3G6frhaOGzNFjTnW8EAE0u29yxBFbOzwnef/Nq
vfPv/2XWEckumCaKKs6TN7BcRunh93civ58wkkWXGs4tRJ5p0CsQxL/05S+e84NuWY+/ujpToJ2/
ZWhvMyg3C9ye1LQnS8k2w/lwnwi/dnVKcAWxInUkXAbmJ4KRHt6h6xqy18XNvip7Gp0QamupUuVK
Feal1xgKmr4cBfIuCTmUxF02G3KlJE5N2EbcoSGOeLAIWVcTV7SyGzuPuwrp1yLuKgBZPOTxiRS+
d+5MrOllEVEuEg9l2DKiXjFoXPMCOf2yzv8Em50nzc9qu/nKc4GoulS3w/+NdpCUMq13Fyu93j1B
uhIpaZY/Ne2Z4ig7n216ZdoDTT0n8BrpWDwNMqQB73mKqcrovAzlnvwFguhj4RUJcUbmCir8WcsG
vRh/exVsCUkOjvTv+AOlTj+3S927WYd7KuUerPfv3v5sHyDq94psiWFSGSeJLowxEXmnR9gRKMU6
6jSZ4W8bqiycwTFgaE7urOalMZ1HYeB+rDh1t64u1bpXnl0NZiKHz7GELAkcqfjjlF8BKwcATgvE
JXk3wPTz6crLYJT6chHg1Y6yyxiEf45OJ+kYQDHMxayJNIjhd5TmHenEYvSKR5ejFHuxFsZ2ALrw
OFOx1BEAMZYSC+ssbkSNZEtt3b8vH3e79yCj21XmLJ1qeBkkkUUo2I03iut5ACv/ubXAyaurlo2g
BxKvK0ppvGp3JehkaEqB5vDpjHCNAOu+RHdD8a2Udek+NgFv2/dO9fpHebUHNtS6y25FbuZoWnYF
EupaynXX1PBjpP1L8R+RlWaqpUTXIzUzg3HjzM4lLwwAuq64jsapE5DFAjCafOfEaFpnYNVqClhM
XXiHeUNsNzkGEzqFFvMbeIo+49rsC7Z39nsgR2qNEl6/wK9qW9WuF6abL+rKihCml1a7RiizAOu2
aos5gpXT+wORgfaP1DuTK/Ml6keg5fX6dtjw3bLOlGC+b9t1sNvG3OGftpHkjKD3DxlmAbEWBEs/
8sSApOE/8k9p7rz3skI4lqYByEYkh4YGjg2oCCXbiDrQT/ssJoeBoEo2TKGsCnsNcDyhCIRAjIbm
oW1mgof+p95XIYdvEIwGexIGxV+YbYKKXLwrSmg0yoIvUblAnKXH/7Jw3fWjzqjP3GPU+JpRhvp1
g8MWRWa6UowrfDgfJyydepJ9DGT2JFVEY4DSTigGZfRfE/ZRi/rCnFs9Bg2eR8q7k9zHL4ZF7XN6
zKGPfQGVqQHWSq1tZHFMsr+z4LLvfHC1EOW1M/Z4t3w9wB7cWSIkQMXVMrBx7d/4op4oYV4/JtMt
4FospsKG26Kx3tK7GqHE4hJ8/9+NKihztFm0XMltcaPK/tbwQwgJfl01XTZWBvSRKHQbd0VRVgbS
4fFJV8EQs7cA4vAyc4bil3TtMPR1JxvJfvNq0pr6gA7c6dneKJvgPY8CksZm0lx2UWCkJwag21yr
9VDm2Gcp7PEJMkgVhH6yxbfTQZDfvNXR+IMzSDTsUjB4ujv4vd0S+yBgVvqJUvDeov0yKdbF9B6O
oVSBPkDMD7ljtQZa13kU0qGnCOS9HDMXGCFHttsHTBB26s4lHBJmlxPbHQYo/Ka1g8BMf0TckvMx
00gWOzKQBLCC1DOrHzvVJ9xFnZQlg7OQiKVPqGeYFzoCcdFSfe3tZyd20lzSGlx+0MCY64rWem/Q
91SrlG4B9CylusuUrVDDOlDmMVnfcw2Iory7bznxn/5mk/mT5UuxMDd2BWzv8vjDk9MwgSLYAdyo
/RIC3X6giS8MbUyPhAQf8Z0DxSRI3HMW1+DmdM2smBmtM6AltknctH8oXyRU99ZS0/yFQK5SGEMW
WP+l7mn+lxGhnYboXs/mZBZigKUw2tx8zV46259so6po1kzqD1GQyYDuQitSLFRcU+sAegwDi9Kx
8qOuFfSJr/HbEP2tDZzLtyRFyVqfNiUkVUxgztB0j/EgxATJOvHZVlfGYQm0uPXI2TJtYpl2WkGP
GUt2GZZLzM7JdsU6fC0V1Kx3R75Vn6j4H0w3BQ9HHKQc07lMSbcoPYr3D0CSEKb3g3P9RRH5AqSH
8mUE64cEuLyjn6Ie4dTeh+sXjZoBQy1jMbsm8NNAH29lh77y99mXJ1jhQJHI/q/sFxBNPPKbOumE
ekpnh2x8hFGPG1ivgUhZNcO1QNDdygbvxnKy1obcxpt4ox9Y6yN6WjFwpwb4d/F6tykVQik7Z40g
bs09RaJsSLk05KwQOixj8Zn+p74g7GkZUhy4QG2M4uCAGHo/9Bm6qhsF/1oL6Br9ixIgDnCunTme
QsBj/nKrrqbf4rclZzDvUiA3r5tsSxfwGTxzAZ/rT8d0p+Rld648Ogmj2XglW58rc6MuqBy9wEKB
XWx9jPbRb5DG35p1ZjuhskdsslSopdoWIaoXHhko49Xq1qemFIy6dPXGoF8qA7VS0cxI3W3TCdaS
L4FC1Wb91+T9X45K1QR7tA6e6h7JDgem/JRhOX4c3M6rOplsexVAaEcKaOu1dwRkScKvhJRViIab
ye7z6z4DYdKxAIRanqEksZlNFsPvaiWNd58tKuFHKwu6ImLj3C5JYTvCjKHNsx+h8cfqYEiZhMo3
yosXvHo+PSmW2HrrDwlXg9y1uYKM1/nT6U3C2D/gE/Di6geifoVn+CFfPTd/93x5MD1LI0WAu8iQ
bAnv/hRguwYqMnOK+V8fvK8ENuSCmHYsc8UhCvLmubC8ODhEzd5rF9O2yqJ/zB3VwWWwOG2NXlA0
gBDyVDbKB4Zj8dKMgAcw+6fWXbM19k1/Z7mlNEsk5IaOYVUCHgJ8tTGmgoavAQv3q9n/PH0ybKsU
vSuw6IUE/m0Egl2Kqhsx+QshlfTsQXvbjaX6iq7bg4b0PwVs5ttsWcnGc3BMe0VuG/ycpU938lE2
OrgYJZ0GW5wRMkFPqqwruQZy/56EA07Sdh9aMpxNEbKekhjRherKYFRhRlBouf7TNkpQF7deTkek
mklJS/3aNpTSwXInaKtjMo82ifZzWNOTmbGqmFqjn5m0fpFRIk3er12wGu2JCL7eghHCbWqzmetW
qNOPMu+XczJzOxShF0nj7fUDxZKHjVIe/p94C/dezyM29P+P0m/UTh9cp9dY5UmMsIR6sT3vP7Dx
loI62R8LHunv8flWMIgElOlPYLmZ9E/o8jRdLvHwK9vNCysBkNDy6B2lg6AHFvPEFKUXWXM4YyHB
TvNngctkSL633S3fcgIbKys7CAemmYMtJykEdd6k3XgKdg/NmrlziAvOClFqTc343keyzcRKjcyq
pFfYXoY8tGKiy4yYfnVmr0/4bdSKii5p8bc9G2z+7qMdMnV63M0siqsKoBJDxX3Sh5TGrF9bhyC8
hGXGOrBfsA+eSN5KjUXJ5C8fwBEXU03t39NozrT42xiA4aA6kqu2uj/QqRoAcZeXqqpba5e6Epyi
T8fQVgUENcE/uaSdby0c2F5MHp71q6uOS2+NsGE86CGqeIrm/FAmzM3KycZjjql8w51PtkqObKMz
QNpQuqznxdiKxT2Mt2R9K4P+nm44ka1bJrldDD8kqoZ9+J1V6JZa559Dj1xILA28OgUkKq2Tim5x
YMPQFQaeJCWJbDnjkJ5nBRM6Jr5C4YvsVccINctYk16ZDydqONaC92HdHYksIHxrYitz2fsAU8Ml
Le/ilepzJLcfclEcw5lJJzb0JuAar4TEJEQ59ODwu7ryaltSKUUc0jFMDy1Lk9z4d0Pl+cqQFJVR
/SyUmVY25h2QFkxHdLz/Uj1jHe3sDD9c7bUr1WtaeHhitTtQktIbvw8iwuONqqPPN2glwZ0Zpi+7
aZ3vTGiKDko+Szs21pN0n5STrkreM0FzTTNOhXsVwceejLcl//U1iqruuOPVVEnY6Dk1xT84y1Nb
OgiznLYtAs2dDBwy3kOaOuavJ5Ojxs+jmBr4aJ9smxFItBv4+3+btL/oiKHCQN8q+b2o6rKUOb3y
pSF61ZXV1AZWYBV3lqgeZg4YsRVzo/8QxFf6JYJr/jiF7a+f56wdXK0jb0w9gSrA2VSKyMqLurcl
o8va+PcqYELe7DNwls29CEZFeOf7gDOvjF71M8kDqyt7ntSAEhBGNc1jEmVj/W6JGNTQnEN9RqRc
BLBBdJMJl1Yhsrii6EsmsjWlRvd/D++JHBa41knrxyOrW5aPxwLwOiED6oA9AgheXmzhyGPMctZY
g1gL03RA+kYBflrz4pWRBN3eAjF9WaNwRQz1TUNRfkfPTKM71y/EtxcKmeA4f/qAq8L8/2ar9vWO
/SheAuq3xWqArPLnOnrNScji7GTefGSRPiiBOxbkBo7/puozhpAemS5AsAa+MQVF8/fBq/zFkCXJ
Qy2Tkwc88vLZO8IsdwSgGNF3igWUk//aYxxd9ZxVMNwpIsnMiIwatX5IRCPIGSqafLPo5oMFhTdv
JKKriKVkhAy3iEYq5gm3p6gtnklvYmSXhmXiH52opKkvMdgCo7EmnZto9vXI6MLXO4cHeP8gj+iF
63Cf3cLXq8+WXPSjVhF6rCYEhFdkjzzKiVObM7ffDsH1fpT4lLYpr4LkbPBmP6685K8ERsPk02t+
5WZO9f0/JSgMulpnQV/UkI4evjxy5E5rgU4VKMm0CUE6wq8WtghP3c+7iKnZUG8rXpVjgh+VW27u
Z6/ll5dvhaBkmgaiYhpLWcTdJIR7PY/nOejyxtE9K0OrTwth8fK0IPlOGYRMOyI9IFrh6TCiHq45
J3iZaFidtdEHhPBTypsM5HBDfUQhP1vsdikO2WpoIRiWHg8y/UBKJDtNa4rg9QODeJbeJ9o/VXXV
txTS3quFdyw81g1vTZwIxuT9UgLPK4XTHpIDUskq11XYm0jLxbHDJDeaWlBQELtDXd3tGKMiFQlv
G7w9lTpt5UwnHeUCpNXeY5C7afF4NOyY9XyHM/Pn6CLEGKB44vLNQPo58VTpdXW8rikBstYklmWv
wdxT7VqvU/qGKxeOYw/lN+c94yiBO/p+Jsa6X/mHoKiK66ZjNEwo4YPYuGFLz1jwsgj0rxTlFApR
FPVovaz7LsU8ovnT2zIYGjeI/ohm/1GOd0pq3J31yj4/scZoGUypRC/MX9jdepeVpy0pPytPtVV5
GnejE770wwDTJApOkv6E0kycZgx2qqLpkFvvjWI3ZJOQB+HPN2pm8uDBJVlLMcpxNMcVudfgpD3Q
CF8YdSGYAdSlzi9yesYJhHi9c6D4BtK2kg4REEK2o0BAj5IpKYM22yKTfXteimkQlp4SCXImAOnW
gpRUmmNBsEqTRq4BljWIvq8Lm1TmODQ0lblw9z2v5rybhw7BudIoKYznIbOLZE2FZidWaj67NmHk
SJPX49BKOVqW4rUZqFZ2MxpSNv7HIzkj68nhPU5Vfnl9OCviDlfLxRgHnHKtMbLQYP7I7sjffQga
rSOmZZXekozEbsRKIoJuYt2DKTf8dcbS/hC73gGtswcquUYNyTf6WusDxsuSbpCa0+lEUg6KdG1R
mVjNSIy0Nw0igxekOZyuD4dbqUj13WKh676YjmzcwForjAugK+tQ/hkNoDqyuq+KM/EzNRYDkkC1
m20n3MNxB36iqJsorhhhhYV/qBssg+3jgBsbWjMVOE61d2Roh2/C+ldK0tQUa6DvQM7b7cE2VU7t
/I63xC8/eTWq2+GLOBCE0id2scBTzJUxe1o6+TKtvSSITzI3AkcsDO8bmi/13gEWkPZb/5qvlks/
A8RY7juuWyJYOEzwU/5N8hf8P6CTXSy7T9kgQ8gwZ/hmm5ibM8h9uuJEtg+Lyjy6LgjS0aOEUK6s
HKxmqDGpVgM0FIv1aKP/Ln6mG4DF1W3bVxwMTzDiGBv0/DeuAgZ1v6KlLSRU3T1SethUHeJf8OEo
xEdrcevkKfIK/kbCAnNoQCD/JTvonNb9fvFRMVMQPekOs6btANXgVyUlI3c+9pwRbVhVTT0FAps8
HRBSBmQ5w4ZoWnLDsvVfH08YlGpgK036Q09ONSsin2AkFYIwWR7xAVIbyHb1eV/Js9LzsFzcXJwM
XGQufCTif1YtpjNmAF79NKOWSR5dKinB9oH2stltyvaOLppZEvrRwKzB0CNBSNlRdOWNSXAyChNg
8xbezVS8J3Z5FVkz0cff0v8/cKbsKi7EMaNWbx5p2j8ngAK4cPJO8bP8UgBVuug8UzxxzcbL70QK
yNNJrZnrIkEmLnF3XK66k5H8/xvEmUyEkWLH3hyouP4fFXBidYloM74g3xtToE8F7y4Hl31cfBY/
I0a0PJ5QRIsjkeedKDqvLZv8UWJ/mWBnj4sdM4KTd2kipVGIXUJNYIvkyDZEkcRheNf5Bi27d94R
MyvUocyWyU2NAboiGGc91kGxj0CpIegxvvFL+EFH1Dd0hh57rErjERrN7E1OJms2dxmdipJYr2WR
NRrlcsFkzT9tisDRwkZmOJlGhk8795uEnveCOS7It/tmvjHpg+OWXWgF5qCVdkync1wnxoB2MrFv
Y5VGoitANasbCI4H13EK++eaRDwwVhMuidWbB7o9vmoWe3B1jZhSQQaKRdpm2Mt4VTwozJiRMQj8
1LHtJxR0iogurn9dVo2AGW6TvmgyONi+eaOOVEiTRZIuiYstgNrgtI2/2G0xD8w/h0BoftsVBc/l
6TIsDy1sD6JWIo14A8nzrpcPcvfYenHRvLdDQ4YYj2ebn6/P+TwgWTOBG42Kq0ugzP5qQsGAK8Df
0+rTWNicwsQof22Vdpc+fmXT+BGy8hB0bbrC+qD+INN+Rn3xB+nPLuOEslwKKOG1gFjtPf/TOsTe
ZKol7gyUL1+i9WDfP2aysJTxSC894gqER4GzBMfBY6ULcgcbAs5I5YBc1JiXz2f92K25d3M1ax2a
I/tdM89LZw6PRb/3vT/qywUN4gVBQ34xdIUujqkfAp0+vTtr0OcnQY+2pmImY2XfovBDGY9+b+JH
Cy2YcI083+0YoKpYXwYYNJMoCAlYheWwlz6273sfzOJ+tLDkUh+IYztQX0vZD9KTPJjjFDOKuRGq
L/Y+eXwaPkrxt6oRSiFf5e0plAmhGK1JeLdTOepCzTy6H/rSU70r5U8RfCimmwY3Hhb9f7kyICLZ
GuQquNvm2lCGPDbLK9+JB7nKtY3GpYHW9SBt54aNr8L4RWtFzlseP/oOJjbBsWw0JmIUyC2j9+QB
ZcKJdEHFuXXcl1X1JytG54rWqa/iuKV+cwe+OcDqhS6MpG+B9wVf7b6RXl5eE2tbYkZ3XCgosbRT
aMsGuC1udDSc/RJAPPPMwrbhb7JvXXxU+xwxbKkbu+I/6WTfELUUXQJZzhzp051mgppqA/mqP5CZ
QM36q2KiTd/kY/1ub6HtciqHETQ3qGPfZtB1y5YNGQjQmIA6hj/Rd+FtwT4UOHdaWhAKBENlKWQM
rW8On0V4Z0II6WAlmL9jN96C6AB6hjto1yjX48TZaoORZmYyreYPI8XhaUYhq8qv5PXrdeaG0aol
4RZXnHv+yoNV4Ep9CC/eWPN/vkOXcOL2W5UtBkqqcimCbRME8q/GT0vEPFzTAc2679vijIKI5RsK
u3smKJ8N+byCw/7TBN7K8oX8b2XX4e9UsFfnW8SWAbfogYztM+YJJBC6GTCyeNurJRT2emHp/1qD
WBQrq+ymlOVodJMRzuJ/AxYHpBtR/4DgawqWmHDj6zh57Adfq/sfQZIAcS1PxkT/fkPGTsn4GDSv
QDBxxEnmChmU0E7cgiyfGoqmxTP3oSkNc5EbTB9CGO4q/uMqZaf+TMp/RSd6bue/5RDNZaGmcWCP
C5OoOLfek79apxF1REFOjxMqEh1OvdmdOZxTC9TJ23KND2Z7lCvIToCPfIAO0GQzNRclyUQTFhzE
AioYEx6Im9xYOf9kibTJD5kWmVaYTorfxWFoduyi/PY0f5yuqPSD29rTcWpKN6Xg1QFZ/RBIuIbl
441eL5j7D+/oWZe5O5/kUOthbcho6jP2ZmnVeJt+rxNDnjjb5sRd6776RXedNxsHnPadCZHBpvVh
WVrSIVRHLvDGUaJP7mr8us1fHQEyS41wWIB4ZqcBDzd5+28Iba+kmR4lbg+I+OsGIHh9zjeIJh4I
1hjS9PeW16gM9vRnse0O98Du3qEL3NUsBLcxlYI95SU1o/6bFw/8yBU5MP59XhluGvRUOI/yJ8M2
LdZO6Wp5r+iO38pR4uxh5vCM7i2g/+RHYol2ym5K1tTgMWaIG1SmDcPtLfJlbbSwWjxwrVUryJG/
Ob+RHoRjKxb/f5Gk86pTEhDCXQP6uKPsrrZmjB5so4gOeCa4zgJyavQ9SEIE3OYhRHb++02ykaf9
6d38D4vMWAfuOXact+ON1w9DaTKImi6lnyZmvr/H5wPmxxUxlJUlciuWLGhhWe24222+5VoxNcSL
OAIbICO3xvHmIs4lJmBVu4hHGTq6wsB3LXhnQTuO3PyJSexl9lo/C0g5FVfkVX4hKJwvFIcfOIpm
fYp6lJc5JwXqR3pQ3LPdrRdxRqBAlDCGHrMshUJ4NyRqIxo4Cl8UYBmyNCzcHJyG5A+T7LyQorEG
bjp5Hmai1+EuupI2IE7iS7PcJJZXkPL9UTdYJMxTSW97Y8rSdtCYqnMD799U4qM0gy1XH4v+NOeR
+aR9z6Sti7VkwKyh5X5grZJVMHbBPQE4UGE2jG9IZeT0QKtSgmDBAAUXMQsppeWcsiLA3DY+/6ks
DGuSJDgloSN/qcrW+0Ar/T/AiURSLERJ9KkHh56qmwd1MYjQqWBo7U3XFAy/8I63tCQ9U9aFJZ66
add6uO9kAv2yhUCQXKEq+q3k4mWryWqryTnHFOKWcpKVX5r9X1ng6KtImp7aHP68+8YF03pr4f3u
Tuvhlo6hAczwnxHd5TAhbbxOq+qEDHPKvfpOjZADAfjmsd1TvOSHW62E0FAO2CixYKe5obtTB5WX
DcE/riu8efCSX+aRsVEesM7AzmH8pVl5FXTq4jRvZZijZfW3C9XEGmBgutFN9aGhgp9hODqC+FVV
zgH7auZ1dL1RFs4IJzdvwPEkfT2hCuhOWZwJXc5BQ8ilCJfF6aUj/MpbAwpsTetzJeKUOhcPKQEY
/wKYJiyPmC9xb/WXLRH8eOziA2Fs6ECvzrGddqF2dt5wDlvra3e++K0F9NIbmPgW9vPiIjNcWA+L
Bx/pZhR1dAyuAN7sYEXj8DGAdaXmwy/9bNE/1NYpCwN2da07ydm5+Ym1rjG6xaRjB639ZYod+kWE
2g9GX16Ox0WqYxNnduf7MqrQoZ5C72mjqxOSq4b6agvo0hdsZs62O5fIo8k8TZqZMQmS4dNg5WxC
sKJ4Wt1ywF6xB5YKweP77hP/ZpoHNOwpOqJWpSNGLUnrF+XGLUAyA7LOrjTcWZdQ/GoA2iRIG3On
Koq/XYfFJnsb6RoSSry0c76kjlJFalvizVgI68ylHl5oCCT9+3Q79vJVbiKJGP8uKr2HUwduyIwf
TFzr/3ssMTOVwTjZojW+mCiZ9seJHeeOmx8c1u0jMJSod4cqoKdL6t0lMjn/Q+qPPfr620RkEMRO
wHoqcYZJi9dtGu+IHpkXVWC0R+P00eTuS9Y3hsH1pLWhKRnU9i9lv0Moafs3EZy55xrtTN7IZtAD
o+R+KiNflh3gYiXomv5y+HBvBAutPQRcd1Z1jm6oHy9L2wMWTi7YEL7m3c/iltgMTjEoSUySjPd9
uu6SXL5nDAv2xDwx+mXGF7ECZHtN9prUrgar0tP1zIb+spLoJVUefNEKZEwY/Sgjor95sA5HBdmF
vPyiQEI9Lu5tgkQGpObSJoSawwjey3YIRZY9t/vh383Sw+wdYv1y1dPQiVI6VnSWc+/+zTJOH3jr
GYNJwNH12wdFDP0UQvoQCrxAkkJGobipWcx63IFY7SE93bgJ0jQjbmxhlztvo7OAf+WH04oeuREU
f5RjxYvTFLQ7QXCGn93N6vBlH/MG9OCwcSkiXbMal9qdHb/T2nrT+m/zqKHIxnwTORRsrqtFenAw
1jYj1+cWHpS/TlaQTZeVUrNhbuQl8xxZFtlp1ZRtlxEJymS1wjEbEYev1mQKvEVVnsfE8ggm7qKk
VzvkRIeBjM5C79PY34IHOLmm8Lmtu88eVzkOVwweBF3PV9qiQsSo/ntTvPBME6MIf0TCvZI3vl4u
ck8CccB6VAG1CQFuS6Mi8enZ3t3CUrYdtU1+qXWgGOeryiNpxHwjGMsVDGmU5tDy+GE8+U27bTlr
3+Ue5GihfGuwFeEI5QtMMXmBXhJDjgfEC5lhGNw5Qlet0QQwQ4GM9cGBucEpniPeOu4+PK84UGpJ
0gamwOnAgRUgcGtYbUn2Zm6j9F+pylJA8eeTlSi5kPuFJKDdI2Eawh6vOihv0Vrn3yglq/eUf5qS
UjC8W0adDZ+YKICLniJdor18f5SPxhQH+4Hng2FXUsovVgwyBH3sKKIxFeO2goaNYCVVs4qVI7U9
BO2v1p75/g0Q4TOlzLrMUIztg1dFFAEWKQTC0j7oICRuq1DGakOHRpWavUT8XkM2sY3657w6nFw2
ge8CABUCdSynkanuFTwMmiqqV8iP7FekVKSAtyv0ug9ua/vPiO6XwftpFyMZw09NsUoXXRtl4Skm
vIDaadSrNAJgnxx1gGZwuTCnTWN3ivC0SQBCoSDr5C8sZi5Bj8L0kygewKnqm+eVHl/joN8wNKAJ
k72hk/69paFLfWO62DPPRZRyZv40/HBbV0clGEXReRC4ixAmGNA4DEfNWDx7g2cTSiQ5x2LZEXBq
SbONYqHt6bknnopuBotabzO+DlTu9gSihhVIML2lAIZPw8nm1BBxdQu4kikfvDJRwiyY0OfiRi7h
ZImxJxRcq2+zRhdpUh6YzOb5QoZ7vwNKFINVDIReEF5Xnqxrcf8PQqy0kCE+gDJeHX+FtzrRTNQo
mgA+qKg6j5P97/p4uK+ODDWZopuigpVhUapI8yJ/f0WzgscdL4l5qxkn4Cct6FX39Qx7GRyqy2Kb
YRpTTsFnIF/7OUeuz697l9R3OuDSF81ZwMoNTqdcXTWvBSZCy8u4L9m0+zTHlWhQ4d4t3JiWOFzJ
QOI6wABWLRRDqvYSaAhje0y6AjwlqRGJf0aSh2REoGQLhyqg9G4a26G2rujbiRVNyPxmxGPulJE0
fw3A4dxugpIo7NHN5pbe8eWM8wXWkoB5QcFRa7h07a9v3927msU/bP20GkekQ1CSSH6Aa7BMCzxe
z/GDUoQ8ACz/uClW+5OBbbKl7f41dUco/A0fhQZIb2lmcgp6leet0ucpk1YVoE6yNSf2JzCTRLTd
ugSB5eNOvCd+hOIWFyQJ7sk5A+nVsPisQ/QuEOsrAxLC1A3Fc2IXAqYZdn6/PmsWKFoimMsrcmeF
Z0fZRgkFONkp5vDvxB4P/zYzrvUUAJfD0ae9zUc8608WM9ZeBZCC2Xe+94r7OTzh7jEpYr/P2Dwu
zzWMQB9XRt5h59T6cGuZMJghP+bXmpp0eM29JqZwImRc6ZwsG9RLzdTapAW1jE+2SR6+FFVmRPUj
X4oScE1UsBXmBA+49h2DrK9LyrPIYqzeCK9ZhdiZzPMG0sU21X2SZPFWvhK8xMJDABluqxfMN1du
/YD0qtm0RQpZqD8osLS30Qz2PG2hrlEHgf42+2sjS+foHwmP03HmPZ3HIIXAiLHLQsOiDZBXlL05
TBhJgT8mrsE1FKe2BbEq+i7dbqUlI4bTmrZ2x/IeakEK3cK5aB0KmoIWvjJaFYgQ1rkjtgQD2wiF
Is9Pced3gJLyHFVn0nByCv+D9eX26UQidS6waPYVB+Ld6tyzDBRhgfCs30MLUb9lT/U4N4zALn2d
/tmh1F96k4He4JndcDLYaCSuGGQm6hdQiKH4pKfMPDWvTTupJ7FpvQTcsd+VYErN4QWkhvxWxqTo
eJTziSr2BXX7IU8dfXLcay5gSPevvTiMHjJTuA+E4nf6/Vn9PMQjeuCpSR8k6dLACGk4kvZxtjup
5EJJNdw6gZ1YWTf7w/f+gYGoF8H4lcS2InrGMKMTmjKvpEwAJ+4opV5mIgf/kXIatGTueLsRjMup
R54ijVcmcGGV9zHar8bakRWuHosAq5gxu2iokqH7tgsmVRF4yZ9L1K6Ks1lAFUgDFY7oxPOnn8Rs
RStXKTr+Pm4q5Jx/P7tntCnMaXc/mWP7tl9oJaBsJj8xd55lp94V7dMAn3ejAxZ6B8f640EfwUuL
EBGWLra30W88kIP59SyjxP1Dn3++MU8P1VelG92Y0KOX8bL/2GiNVZginbtcUKOhxtjJ8ZLpQpVF
7rNtTI9zmqROqG5WkP5mzEQAX7Vl94RiqYBz0wOlwhxEZ+8blP+bWShZYMSSaG900J3rPOR9ZfgO
2pttqgrW1V88P0nUQvVogCSlYoVkRf6UN7uPtTkN2H6Ui4J4T5R7fXR9KjcNOfRkj6vAv1WRWHzG
tPsUjihy00aLYV8RoWgmSjvD0nuWIo95VwJXkEBO+g1H9pm9Eax2WnVN421+NmcWv0g023Zcudbz
2Auy8wyczfbvolfHqch0Bqi2/lH5l25o2iYwZExU74Ggm/KW7ih0T6iASMN4W0nBD8gR2sb3TUnJ
U8b/1PfVQi8JjiPPdjZBpQNowASgKZTOS46iibpzfZ67q719QSn9U9Ik4g5HonAmtAofgxi80q3h
nQM16dC5NRS0OLJO0o+sWIK2EzAS5/LAmOWNW3R6oSJLYesHxZQHZf2nMeqqqmZJ/+LyyFJutGYP
cWsL+mfrItULoI8gbrV6ImM4VmatKO7E/7XR+/bBu2+azgO/6hhKycCyzM1TvabxdhrRUzhAYcQg
TI6h9S8bYyw+GhnFy3bFoVVNVMVESdI8j/7e9t945WGQumOwZ94s3NqbfuAmcWkbOJfhHpqiHB62
Q6HecLS+qAeinmBbPGqHvhSS476pXg2US70+ir0KzqI7p0frSZYn9tuGDSNyWkCbInH89wUu6vkc
uIVnLcuFbSIzLvF4oyDVvzL3A3xhDLpGlJP8++Ec9rv7quoeIqDgqpm9TwRCj5lqyPhXaibl4/HS
totji6/kJhDm/94mcpW/hFxPy1e3OGPtFuUMFYnPboo1AYMJyDxCLUfDNjVJYWOES6ZvN9FV9IPw
5FW1zsTEgjcTsaohdyUKRneRwhoCqquyE3CIKVyV8cORrVItQC4CnSQ5zK6A/n6E4z7Pjd9cuq0n
pGzxm6hpW001lf2aNTdPo8Qz4PrdSMx0nXrDhBK6Xs3We66sP4n6qgcErKAr4lkoFUkq7adRdWci
mXGU4Mrot2Ed0N9uGX9xgXMOQzd/r6FQD9jhst+GCp2cfpvuoljKbTLTJo0A+f0xXbGM+b6bb+tq
+YlwaYlNP7zhcEpkyzhq0uKGmEQbx1qFN1C9chrQ3ofZQAcCCSRfkL4cgBxofJlPuhvDwFTgbeNQ
BcApcKvs0dyz3x6hbRPYl7Veu6xA2O+R07Nxf10C/fzVPtezRpIIeQgIV6FtrEr4m948c3op+HYb
SUQ6XB738x8874iIGAZn7etyyvmXnGZuUudV2YVxFJUSkkDV92cnALh5S/FkNHjmgG6XdRF6zd+o
Kl7ObkStZfpesJPVBe+WpnmBH0tf2RMlctjFhCd1BwLXQTKP31CiCnzEf51KkDLicyJA5MZfdFcg
UD6GzflJIqcAIv3XRr+T82iwfyvY4AiRfGA+IRTgLmXN14U0pXLdwvAx3zeFS4UFqlZxLTbG7UEI
s64hCbA1J8kNinBgTH98QG1CQ4OFT4pghRLPkWHY7r6E/7b0QX5ka+ORP8/K+WD/gJLtHqEGKJap
xdosVWI7eveZoXMGT40Gul+uzmYVGu4ez09qHVQfaRI0l+e+A6nd1QR1tA9pY9NxXkAAUZbWtp2p
PfV73xf9k+2+bDx5IQRWkk3koFbou4rcbWSwwZh9bzxKnDLtXhqJjsXZgK7UfssC30jSJ3KvhSih
ZTIuNxoGlSUGmJbvITPf1dEbt3vDJs6but6EEqOc7Ynwv+H/YMPQPhZdoJQvC5Gh7jfRWrNd9MjB
/on+J3+5kiUHRd74nWllEqU/Ur447bhZaVTFae3KtVdJooD0kOEUUiKpEi9378576GDF4Vq+Tlln
ZWbsrO58irBMCqPkS8//54AfdnzqCx/o2CJKbuF8vNUq+iwv5bX49uDHaRvg5i5NdngXRoySutdM
nByAHAtTjbSmzWty6417s56TMPyakTStqaPUrS8zAP8ouDsUUbC9KT6HuQjs7BpEpbQpGYNJRRjP
TmXQ5D5fCH3g2j2IhmTbb1CueHllqp1/bGu9eLrueo9JjMvun/ho5B1bGfk94/wthbtdVw0/FX8V
A/DcfbPBOiWqMNCCS7tXDjKmCFosFenGmKk/HUDPBNv6D5/bdaEf6KYoo5ELY8vE9q7EFnulhCA+
nqNWAiugHnVBgTNTGZ9v8tc2OBVoH56PRXElLZMFv2kx7BdOPQZkQyUJnH9On5jDTplm30FGm2tx
5Y8RKXxlug/+U68LWZr2xRiMo5E1ps9bye3D1eYHgy6nbaWzZ2LDimcIBqK0EsF+vHrt97+6/l8x
/1dD/IBiSvqHUGEeWtqyDsstZ7Alj3K2peO+GEfujhUkI0Ux565E2yxjgN0M+OOS2pAiuZU6qIjc
67rcXvOXQbyM+zRUERH5zLrY6AhIYBU84GhdZyq3pgaa83QPVVq5xnm7PaGMQQrCx7iHOeQBmPCW
zIFDYYsoyVvltKNtu6v+cRuObKJnD0ZmAPFHyjIh0Axuaxre+Z7JtAzrn+cCg/YfUjDi32SeyKIS
F+z7IPG9ezImDu3ise1JLgbz7sOg0BGKkgcIsbjoMhJ7lG+rzG6sQcP8tZf8KMDpjsoptFwtuc8O
GQz94P7ijgRt1eSLkm8iwmlNw0ps8uFtWc/5QnajMOlmnmUY3ycR3Bpumb5ZeCLAT1POEK679EtA
Rdahg0Rc9f7GCkzdEJQcwdKNDRN4pYjOMi1ypFPUZLh5+Gjw+xRakvYuP4USC3vcS5Q641B/Mcmb
P1ebxaYmjCXiBHVVHh51QSfuhxbWAf/XCQumMFpyKkxnR4oMyamFLAe3XggNOJ/r8AoD08N58Qy6
9GkOREHFJaCBBwUG4/+S3cx7N+Zq3FYCRHm39K6ruLD640uJeXDjvHcioQf8TUqQg1JB33qRzgOD
Pnk7/ZeVJFfdDdAim0tVK4p9l9eiS/itd6WN66BY/lrcIMBsGsaggXafmp74LKU+j0S31VqkLXsN
hzB71XgYIdv0TTP2+UQhMWvExdDfJ7JwBn/6ikU2oHiZYPhlXU+eFfHmpBn8IYk9jXhIk0BWmYdL
WyV4W60zmgk1I0dUGFtcLQUxIgq8CFztqP/5ypCMaAbevMO7PI7hLc0eSr9iVxixUQ3uBG2n6+zB
SN84wm+v2VuGKIxL4dAiy1A+rWPKekUGY5HTocwhwowNh5Qb7vbNooshbelK2xM2/An9kObbREBz
qEqYkPxwiLeWCImXgHJv+o6CU+DKDIp7SinMZifnLFqjOYq9aLg9Nj2oonO/zVLrypQoj61DchEr
lw8El2B5WfCDbcT3r1RXUDyLqIFqO4nI6/1MiEvppeT5IRJqwsKQr1KJbxaxovpJRn1Spo6O4b0z
D17/XucWPMk7PYc4h9IXjoBBg0DG/sNZpuD33oAvwIjbix939thIIZMOlvIGEERMLtkIfZKQyIIO
DgpPL83RDGqUglt/oMnTHzKR8l/OYkSWn3dH96HPRcAKPkzGSpTPuoI9gnpKOesPj1f+DZL2d+za
YGKSCMADAnri7LzJsg9mYjI0gcmLHv5g+KzjhEVZ7/WkNgiHAw0PFMWXudQTDP0Lw4b1Tajf1YPS
AlGwE9CfJp8ELB9aeZ/4JZkeAvSfEKw++JVD75BnbkGyaf5H5QJ0LovFdzH5H1JeM5wEK6CMwAQZ
ceWl4FZvrzfqY5XnEoRRorD8l3EZ+zkBz2CoJsLaE0/S8mPi7N06n8TpViRjo4D33dvgyOBWV1vS
M9dErJOVH3Y0elOdx2zmUKsqIdGCzHWC4A3dqNTrAE+XP8ZHz6i0TgsTleI16PvR+HLUrc1e5AR3
9dAS8jfLe1l7V5+0GaGl//Z5OaY/vL0z83yOuL8OHDBtBSiiS1RXcpGaYJSbztKp06jRyYpFvkNV
Fap/vu/Hc7QGv3ope5cVoKrZuTTufbMgYcCkzC6Rl6K047dKVhF3omGEiQS2JMPNEAUsGTdKNvUs
sc7Jn7zcbJw+ldaO8ZhfQoHhcjG/Ej/3u7LToXvzL1ObaPdLTAfFfV0zciZHOcpAA5fmCeNwkza7
xPpVPMLPebL//PkK2PMBD6ba77JWdeMaSCWABaWahfjklr71+MbObZ3jKhpTGhCLlUvY0sCCv0AR
HH6f5r12A1rx+OaIvqzcLmYI1XuDiflSNeiYf2GMWKZPVnNme86j84Lq9DcDtQudwldCRDjXM8Z/
wQZRUmw6ERyDfUAqk4Ju57pg5IyhpnhbjYPbaNoOz103uArnYWpWZiMS+qKuzloFKj71FeVa6kzc
rH0EgotNYMU8G94kRGRD3cd+KuS+PTUOYQg5vFB0lT79CXVcyX1AIdo+rE3YDoF/yHbyN4smDYnY
vlmzrPCDFM61Nd2qA5GSm9yfzBcNIqrfM5odC7eGtz8tRtqwuA9BtJw11fy2DSUXeIzXibdt4iiN
6QsYklkr//PcRyjlc6etsWcStIZWCyuvpvZx4/qGlskPZRrZIvzADlw4QHiKQHOw0G6OdRGK3Wqh
t/E05wlC4ytq72iK7M4atPfPPbf06BK9TSCPmKV1Rju9iJjLQ6H3nx96rWu2enEfVjiAm52Z9rbI
3ovU964NGtb1hXWw0lpy5NGLftp7DeV/r6BhI7Ll/WZGs4mM5DKOFrFFFTbTmHKXayisiK+hkg7s
LnXPzmLIAsZgj6BiwoFiIdKE7nqC/3n5b991+hgV/71mHiP45WoPQkSeMmTAGqV/nzrGf3Nx4QU8
Cb7UvpL1F7+Vjq1cjR738CY+DTcw6aLsl71zo74bPO9hCax3d5OaWGWGD+/zwBhuMjCUI6zIvMtT
ama1dQrSJB0BpDaqXnGao15g2ddVvs9v2bk5wPAnjwUwSXA69V/6hHSlddjw0wekkIzvXebDqLpG
fxa6vCiXV8nnhxOiXzD8Bxe5PoNuvh5x/T02szb25ZQNUrJgTLlYOwF6GD6aYyA3vs/zW4FDJe7t
Z+ZDKR8BzyBhRjjt0UKjzjDeBAUQnWEqni9ZEWCYd9gLufu5/ts1lD1a/6dKcBXtpjP2/2+Mkey/
fUVYH3TaWqDQlYC2Hx8zSF6cf3Cr9466B5OPg4PzHBbSlImcDwnplzdRgOiRQJMTl1wuv0y3TxD2
sk4VhLw4MvbW5lC8+Z/xdCtEDCVjOpScmJ/qe3C6QLxiHCj/aXq2U7pHBCnv0bnxc5RXsv2ZThti
GhMyE1tHel+qm/FcWUKqV3JNG5ZZQ/0fAFFQ6/NhfYxBjr7pgspglDYYjBt7HbNhrEE1VjsuzJxv
SB9EUO6tJeCZNRqHw49wQVd57TnOeuJGFJRb7JUS6udDTAlTJL7TkVCMP5ZoYgHnXNx3IFnLi86g
hRFD9CfO3fUsPLzPInu7XZ+wd5JNo8ZIrDwxLgA9mvzw0kurmF2fzQJx0XEf4ihWcBrM9ADf/iTF
ZXP2YKMB0hKJCmyVY3kskDtTg5cBgYm87Jp+muitu2lwKW0K7TPNPk7tKHDKxsylKfrNsw+MxdH3
tcj9TePWnO2+rCkt0Yqfm6uWk+OwyYBGy7TmkM5cUqZzuS0R0Hqqof361YRhiuKunlviRlYv0VQY
BCd8gLkSysso1ueAEAt8TpJGNcJ3kv+DN/RgTule+e9ZMzqD0oZYWIrXJU0U1zVZkz++ixSy3064
xQ22+T0ZW8bE6DOWzhwe220Eh99O0x4LlKCyl35eWhkVJ3JDLvXbHuUTGcOzdNNsPas+7eAavd13
CZzBkNxBAHSJYUys2N8ew5YQ4P++IIM5KeD9FvFsDdTuJBefRoLNdIk/x4GHi/TdQqH0zxHF1Net
11nDFBQc1M/hWcUJpgmvuOHKSRbk5qdPD76cls3t6DKEewcypUAcl6bjYk7J9rAWfCt5HkAxCjce
LzOuRYpEjVCb4mWm6SJ1zbSa9tL9kYsR7yGSHNMKzwCwe2kuyjvs0jkU3tisxPdSTcISNKEMDwlt
4r6DiF6VoFh1ufDyXUD6lEOpM9SW1oChNFx/r5p4Owg1/Z7Xn0rL+XnjkGeDp6ylfQEZG/bZsVJ2
vPYRIHFP2RMn14eC/Qi6g5AnwrGwiGa14YpITuXuJMa1TbmTQWqJUc9T+wbWysPWHFuqbPGMwPT0
dPxO6T/XGMtMEyd6ABbr7bncZRRDQL0V7L0Im3N6HX3zgT8RR3tN1KdDhGiPdCRkS2dnJDjQ9FkM
x8GSW3YVAIUhy0wAmP/b1fJScLzZNcp2lWUfsKMyiR2AcrI3a7JhWMyE54wiEIRUwZqRfUO+lUXg
fGNPBEohY815WdC0l9aKc5yFd9XWkiUDtoBn60ySOO0jNW7IF/r+3ikNK6lCxYYFLk1T58EegtCa
KYqBK2SpfzErh72xZPKIC8zW8Wl3Vi/oC3ncyn7QCbscljvBiNx0PrTEWJLJEJpbBlEEdNAhnr7M
OxohwsCjzibf7SaZhsCn49Fm4408jNBTfmsumryUqJKul1/Oi60052/q5Vj6uGYMnY19ipYyBdTl
5TEa7bDsjpoWzfWUJmJfclvtg0jy+RDrpnEkH4Y00jd4tVR4Y8PtVu3uX/MRgr7Mx25UPFC2WzBd
N2zXjOCcLr5d6wmgVfDhAppFJmLH7XcmthU3hlTMwKx/IFUxyWqJPrCv6lxF7S7nfHxubUm0jWty
JizgFLky4GTA9PpgcO90cXs5lL8bj7/4DK+026ejjBXZfm80HhjJPXuuWnMGrsLkd4garmEeRN0/
r9W4OBEJWur2PlBaLgNDz+U8E0sTUIpx0troceLZ4nlgMD0L3m76SLhkU1+zCUV1435JrzAvD1E9
NMpVjbr12LBt8N62lE3zLBPshV6aC0ElJblJAJWupdFXI8b4aShe87F2DytrqSpXCAHp5q+vmhCw
VnbvGde1Z7X96IxRE/g6hX4lQQgtde7euBjALHsjO2Yy7H5ue/cE49uQGkxfYf64vPunC21yV49I
noAQVbVnvNs6UgNwLzX1d+KOHG+KLCDHDb/W7tAVKS0bHyeNrY7Zfm5SYNQ9LZpk7vhhw1Z8RdPa
njpqTq4YwwprY167WNHqCBJjC25RwLeyTPa8hNvG02ZxISi4oC1lWpA8jJG3bHf6zYFWoCir2WuC
/ly+NcB9ifoXvx4vMuwa3/ww2J1t0LR8n/AHN0yvcFGb8vwPDKRnVd5XKtYQsA7wKlveOES9h0yA
Nw6WXdjYzWh0hYQwDjz6d+bVVr3VkKBNRcWcM8HNzFAr19ILj6VR6RJZj39Qn9DsLwYX8Ogtdo+o
38w8KIkrXh+pUh9ed+orWsv8V24TBlFI/yVjutkGg5NJEprILf/Dv/QFbkoKLvK0cjB8oyndzh6i
3oYbBjsAiLeSuDWeYbykHi+OJXmsh6rHuftBhyg416DTnk+gc1v8pbH5Q326qxmU5iyKdEyknVxP
kuKw8FVSyB5w8B+EE8vvCZ5UMg2NpAdpgG0PQfCY0eS3jSZBudYIzb52bQc2UeQgk0mgStje+TJB
ve1jheMb4UDBxwztsgbCzk4nbnFeaHSTFulac8MxggNJcz1YgYKjn10UCKmNS0CR0dN+5LwsR7wl
d6N43qMaX/1RSlFN6QWewY8V+BfSeuvh5qKdTHRB/D1ztcD86tmfNewZyHAfQvkTDT07rhNOmeAG
4LdOSNAvoMBN9zvJgqBb88rPQMR/n5HwxghQbekOpaznT37XjzbzCVW1iqbY2y5kXRlqbIOElCou
msBPEvN5yszRwzGkeIBIOdjl0j/7RaO1LT47X0JN281yXvpVy/pGcR+kOIo8uCmEN2qZ1l2udnU5
aZ4mn++alMqpg1IcAoUtzYZix75uXMcQOocX2wrmfRf+/BRxP4a7yS59pS7RK8dKPfL9nQyCLzY4
Myg9bgiwrNNf9hXf3y6BAdTp+3os8vfzXiJko1zkLPoPuqM+/UEXPNG4u6zUUA2Ce4kJxJ+ubhXh
gs+kvAn+3EgbS7y/lj87Zw3sUCPvFdQ+V3XGEtSgR8pSIMQXKXvOEW7puqWGYmxUCiDC0qlvPWvh
XLdPNe25gcpoiqhno+4U5hnp22C8GJmU6XNSwZqe5vo+nVIYEYY4sv2VdkDs/lEjbqVM/pFh4jrE
gpsO+73HgmE5XV+MVWI+H+U53BxthPgwZvoy4QniuFPij0du82iwu93cG2qguyrWGfKI5gjAHr4I
DSX8uAmAxmPrWXs07XwjUt8QGTNfaDZoYkn9p+rn3SKtCPl0h9CwZPLFAJzLDJ0J4wtf7XjCHJdm
7OoQ83oik71QA+HEa9b2xGvAx19xUOfA21/mTIy9A6zIXr+mlpJ0H7ibOcpBjyp6bmUQOfVjtmDj
y7OvYQ0nTQQNESC6jhelvkWA3g3qYinT4WZcOSyxvjnx8oU47E2BG37j4GCuVZ/Ywcq361ZOG3gk
CcUhm6KTgQZw7a0OmLhdoGyI+3sYWC4/OyzWy6UKlrhaHqB4/0KdryEfb+k132ZHBOx1gCUS8u2f
2xN1RiMSRHCLtugbVr/TIobHDybDvoPKsUiZFaXtTICfC3NooXUJkJWKrgaafyDSuw7QyPk2DRe+
SD8QiWC0sw0Qx1xxk1+ZEKBbUYUlIk9KAYzbFEyxXjy8KMqPl4wd18UzgBz3TOXXESw7Z9mUHNkS
C6mNt5fzb4PU12R2c8GC0dv0z8GmpgW4MzLHl6BTR05Nq5eAlUF1ZHyT0iU0uUKUlOfJ9WUe8vD6
PMsgnac3MauANxsUUCheSq+VX5RLNGMhXIj+W+fuLPQ7k1zxUUzrVDcOuK0cnULm0fny9mSlB7uq
Ln1i3jd/sCA8lW//Ewrl+ki326PYuBaWuw7juczffMTb7g3dxCgxIG9Fq206f3hH+/CrWP7/Sk7w
8X8hMIhYIs8Mpw0M4lkaX48Pdph1CBDOIezi6+H5jPVF8OVAqOqONGW3UMB0PtLf2C379prk3A5N
PT6D2OmaT0q7sA/H9jd388UoONOsaNXjT2zI7Zz+/6JTPZ/1YxwlMb9J9i17zxUncy7jOk6uSQh3
Dc0YTMDoBPFUyonWg6pkoriR9lougweEXw6k+ukK+zib4UMabmFC1nEPN+/AipX605w3ErKanK75
PemJD3ecM4tjHdL/0xmDvt73B+ERpqX26AuKHsIcb+TiOJrhNC2n5Y8x0Bsx0qdAUT7dcn02s+kr
OiuphC3x2GvCtM4fmiwxeDO1n+jwYvJHgyxGi6BT8WnuVHGEHMc6zQ02LRhQfGhVrlBEMVkTq2zK
J6SeJ+MueX8BPj5lsxNCQ1aB6Fp2yrFFiNyMv0XQKjpxOMzSNPTnYU0jI6LJBE8jCppcMQkZGNuu
RGVZ77fWw4H1FnttEkPxiq8MyQbhplS8spjKixzCT19y+IUDmpbs+nmP1PmbrbLBIVh17Pq6ma9N
IT+SVj0xVs+kGIfUSxsdH/v0TzjO2uR3Hyocd/tGDX0L8ybkLPO92xwRuvbDsZTAT8XGprIu2Db0
7bX5QrMI5iDYZdVVSq3O4eGyyaFd3qKuR+DbtsDRqJ88cN4WUwlGw296hwtQrhZzJj7umJsW3tfp
m8ZwOeAF38ooTWcLxQofCNpbPZ4VdPZ9REZA7YHXwoz02W+xWMmhGFiRvq2nUatLGLF7VzAu2sPs
4TS8Yrb2gc6uzPkxNPz6F8PAxBmUd+9X6cmnZM3QDssD2nk2wC8mbOxxYDTA8MqsxQfGHwirQNIg
FhEQNkh0JxpIjztpl78Ngc6A0WUcRdtWktHqk357hOoZAsk9p1uYs8Pf5TjehIBNSpbwEND1K9k0
84L6FYWqefEuyXyrxIekyTeBh6N1UnseTXf5xti1BzkropM48aZzm5b04NlxVo7R3L3dc5daxrbC
vXbpOfkGUA868928aoofCck+IY6SKL6aRr2XwPBxxUr2VCT6Am0pNy4HVtKKkIs85gnY0yckjK3w
3qNsiOwhNRHErNGq+dAu+IuSouJ1ifvKls7pG30yPH+gS1GPdhpw5CRf/m07dVHPYVr9lojv76Af
AD0LBXwCOABwo2bi/aeEpCDIrwHEeC8j4ab9vOVRPoOVUlCUJH0iKmmgOPXDcFJZ5lQy+XgPW/Af
G4PcpI2lL+QHr4Dm60g+5n++vk04tKzda0zWubdtgYffsnv8ahCuPSyExD8R1S5Kw5CMM/c30j1z
9Bc2G1JYoG1Ejfm56acllpHqWcK3jNeOf8v6rd1bKBNZvBGO0GL3DsJr51RjCwSklcD2VETCAN7h
MvCCEcMK41XeNi5HH94ypAJFuczfltYcVS4q48dbOji4PMkkc4eW29GNW9+RdXxupIP8u1kIBzdb
4kYvQ+EIzkySpI+V252jYrIkhjHShAq/OF2+k4bC6KwJ5p6gB7vLqAvMvwGMewUHXG15c2wDdr6c
xRymTb3CvPZViRIuRZyqMi3BjWEV8jVT+7G2LWbbmZNIQ0jBhSU57ju6SF72zSDrfv/oJwT9h4zr
8XTgDOQaH6tvUftywV9NeVreSHEVfxM6W0GAvNbKiYEL8bfmlIgmFAmBcUJUL4cALxhSgF4cM9Y+
5xgX0mjZWGC68lKPlDbisUWpHxyEqTy8BTeiS7Bu567gP8dKcODRZSEshZ6pj+Nh1aQkrmriZVTU
5ztJ+suGoZz10Qsy7YiJfsmz/rB6SFuEDtNY1kH5iLJDqre8HrEx7qydBblwxfP8Zc7gXjWK2us0
/8hA2YnvMNBjcasAAVNcQyrpXvHLnF4GZD1G8J36AxTh+BY0GI/itKpD5QCNvlU4C4RvzpIY5vMp
w+Mxt/FOqcy0AZUooPETYGK/wDdDXPNslqyrEOnrH271CREDIb8/GUKVQrmOOzGCFb+8m9BmHS9/
BXVpVSe8Y10NxwvgMd9gaolUMCOdR8NT92N1zbjCSTFnX+tiaAqpaQN65VAkBeoTXrlBQ5SVuZKS
2iG8qjCxb+l/zadC4N5myIDbtfdRslfk1qBbe/I7H9dqoHmkoQZJNe1qA2aUlFPBTZTJaA0Lx51R
tE04C5g8yL9K7NaIrUyKC10eDs+QoywobrfxtA9Slby5/LL5ISau61861JcwlZLaDKZp9UXfQNeZ
uxpyG/azScIIs792ohZFIyYgvfoHSLfoo0Za4rTzKCeQclLqfNnuOFkfHm9SisKdXQzfdhRRqJI0
6eLHsRTdVp+Sow36dnXuBY5oJvGQNa0flvKVcXO/l0peZX24fWsm8qG4TNZBw7D1niVDQVgs15Vz
xebsfer3V87tsOunmUBBGQFCbtyiO10ut3FkmzG20G1Tfi46k0P+TQJNiXLevkw+BG2HmEGkaqg3
QDTMZjkPSLCQoSdf7O/CUF+t2vkFKND4L2xyi6Bh6el2jqKk5tvXCsEGlhEZHl6F1w2wkTB8CTTM
QHbePTlc5RpA+lUsKFewzMNewCTAThgn4AsiZ4LktUh0CZthRqu5uu5Nv35MJIlqKyqeCx40trv/
Dv1BCkqYf7C4j3khmu3ny9MLMO+dxlUfW61fAb3VQWoutwKt5ZW5BuqbNIoWHK2BJWNvVChlW00r
VntpSmLsOv+Se72nkozKqs+er4urdyetHJKL6eoe4dZemLRVXhTWQsIgFVfPh2I37ne/OZEk0eyz
lMO/HR7yYK8/gFdDHtMtOAuO7VJ/MtadPx35W5OY52mA6vyxK+hmKjsG84ve5cT4WF5t7UUApZDz
cAtzDSWoqQ4Pd+gRtKxX4HPziQJT1OjUF41rFwLJkTE8BEPla0i4JVnpXs8dukrD5WKKOy3pchil
8eNO0iYWvV1BWBmQp6MLjGcfCTObxDsxLhEx7Y3252kCGxsi5jpjp+YMyMDGZiAX7JUJw989jq/h
3sJocLurVXdt8tkunEdqQCuQrnoIS9eyQK5kpnvqaUnepmABKBUuTo/49ZdRqmHkIDSamyG3IsQz
tVgGrDgkuaq6oz8Jkd5lgrf90fQ8ueFzvwyD2UxEafZaS05n3Xq/FL7shbaZ+G5DkoeC4hVZzcu+
jvcaTlrFNmPtvDbeAxgZ38SzmSF02BuoU9rimG6WHHnv30BWlZ08OGvKpA+i2Y47WRDQvAW3Z/0+
OYsXviWakdh1rzWKLmTfWBXATjaoPV7RwuEqLcPLto388lDbT1Nl7UtNRsSV1uXS06gQh4lZqXHZ
NJ1aqo+Xu0xIQ7cWSeJ8/aa/8l9gbA+57lIrOnB61UOorTBrb7pThEd9QjpMLjHaZwYuwZQ2E3j2
NBx1omo9MnajKEIwp5OeMJsjBTEKyxV/o6nQpoikXoVjnxWzMRju2ezLC2I7gtRGvhwkeKZh89DL
gwQdXbH09QN28867SVReGkYH8LYCvR6oIQlVufzw48CdbW9X9NgYi/J/6HkqLl5yEw4GsVjbZZKK
CxifFAXIe3pjct/SVjH+THlfw96rXIdAYzJ6TWmi0Fq24ahK/mXf8gjacfoAFihhJl4diiuQpEuu
y/7yhMhpaLaeN0BGLLtDparfvxeI4Npxmx7trLAtEQLwlYTcLkC4B5DjPWj2vPvrqp7uH8Ia5oHT
t6ogK1imoC3oabGvNATrScRvOjRpNIQbN5vhSxKERGEkost2Q7wIx+UT44AlCBQfDDQNETLAJyDf
nJ7dOPOiozk3rIzhe/wpjBTPa22H5OyC9p94KZkFV86CMeSz2InUnQi4kQVC1+T8k8v5hs1jGfY4
eJyRUTgnfCoJRh0lDOQTKl1K1VLaCdF6RHIhGSd55hLKc8kXyjHm9zHQCevWfdadbm8Y5DqDf8AC
CO3cs/GaZlJ9gqSVsiUrJLJoMIpDGyioZXn+GGHQtTuDYcMSXtpn0ws2qpGHCemllZMukaOs85eQ
D7u6IY+nKmUexoAP7wYUyeoXmSZmo53xMX8DC8sRICutgXsMHu5R8oCRyUtsZCTvJzEVLpVVCTPx
dIugNVOnOA3oRuDlouUDALoPTVe7sDGtzRr5zmOFsQWxUhba0QpXMvkgMJ24sg5X8zCH8x6Sbbpj
YsPKXSi2iVCE/t8FoRXOEEXdm4pD85S4cw4mSndZjwuzuXid2x66xjmcfUc14zLtW77N+5RixvfD
aWHCqZlzyH+TjatLvfCkBPDwTgY5jdbgt5ZfN/Pz970/+/rlA171pf55oyrm3OgwUsQbF1ma2Q+0
ZPBY/09/cLtO4dcDoKwQH9EFvMfqkT0Av7RRc4gemSPizgPeskaALTBEc2+2gWLFO/NJfRrf954b
VK76dxrvBfLc0NQJ2fyr9FCLhERHBonJkAPN9R3kDzjHqfP0kxm4ZAs04u3KZkpgYGxZmZiSmMB0
vAgIKFWhq7w1EKHjIr+K6uB/y301DWMQNC8EKdVzFIaQHqyikfbQo/quJgexrKzuFWAr+kHFMZyi
z/JYboUjdXBYT/+ALYzu9jNLCvb7+JbmYaYyFGxQfzQ5dWgLFnjWn8pZIYkNarz+VjZEIx2+dhc3
62+WaxWw29URfyx8HhMDTdqdKBk6L19M3GnjBQXCHnTQI/XVK9w4DX33+g0Nm3UODgVtUabiGyHh
0jq969RW+d4EYesz5EktQf5GdA4cNTmX039qkPmLOkA7cpsXkQEbU283+LzZPid0S8HKyyBCL1b+
nmjSrWQdF7yrgByM0TeK2XigW3nzCeoUnVC/ipNllxy6vwgqtYdJ8K6OzKUgFo+UFLUjIjkSG9Du
08DhSTT3uhdlz5ZB8nU3GLS1hLeldh5smM1OEJiCwLg5nq8qV2cvDaY+ppElnD650S3XjuEyyESI
SNqmOva3BQgCIaDPSK6IpmXYZrYQP8kjS2QupyqSIfw0V2Cut6cLpfqzQB5k8k443yeVigYxpbX5
X5gIB1DLRO9D4L/zYRNhcBDEkvUWxIvjcpEWRz79ELVTmsDmO0mnbnwD5fVYbeGwLgLxcO7P8Jqg
vQ9gqX1bsmewDxsw+zS1BX/XrRvSqU267csSHDmj+PjWynf9AGW1BC4pQjWDl+tTh3K9ph6/zD1q
dq8JfDostWPOAtFK524Kun9fOt24KrzvtlxCmZhKfcflmwc8hfJI8Z+gMtL0eGoXJN3GbD5+DVCE
Ka7SWP5D5+hoAdX7NluYxMiT1LBXKfpzXdK0GfcHgnAXWKX4ZC3XtCQs+C9N85WjqJuE3jvZ+PsR
S0CulwMLoG+FJl9jA74kj/wnfawKUWTTaujtXlSdw6h0Fiy7MnuCQrslNuXqzudni6wYsmHXUqiU
dIoIKHbLlj3Z0Ki9txxYEw8/j3aLpsJrzzAOe40qCnsA1LI0aICZRa4UZCMBxldE0Xau7tpDJaYr
ccBHa/MYiPiQO7KdPK4DGSAvIHUh2spcJ4zTjdNJWp3rVWKga9xO6/oN2TCnEH96scTtnYibCAcl
Wka+OOa5ebWLsi9lKDteJ2wFMwUdCWX7HWu/KbDjCql0/yvk7fyCg8qS7sBayjsDOz/lDMekZx0y
27Ud1w1OzVSySi0q733sBpMrvF5PUQIH6pk+39izLKi78pjPKysVr84PwOZgk8pRFpfEwd8ERRlZ
4SrMJyGn0lYHWjONiug4tZvV3XY/9KJ7Jci7+lyu4El1EzZ2EkVrdN0PZfAVNhcL07Nz8hQSI1E4
bfjDyA+hEP32I6Y+bR7lSfBNWr/fo6d1hvGjGCJzu8ojLZ54a79Q53e0WwCPLT8EPTPkQtbLximp
MUmYUz9DIFZZ/YttdLD/q4mRt0NYtSDXUaaaGcQ0fsC963IdJhtA8JToQ07eOflg6YTkzArCeBfk
jwOfcCZWnHaly9YkaNPi/f8/fRSDvyF1dOxuwWWWgwpxA4hFzXd48xKmbE2YXTEHCZUX+ANXqtY8
1pm4JI+I35KvBvGl1A4MzoBGtsikABtAgziI0nuwgELk8pW6jcDqAZ9/q+9aaJkAkf4AWXsPs9Yk
QxbS4U5u2cPwBepvwO3viJ4FLBupwPTwmB+DSaMuaAj3C9Ug+/FIQs2VWbMVg4QDJ2JBMxsY8oei
bT8SVI0Ke1dJuU65nnvr7CKHduebPvwVPi0kGJ8CvauEpcsm0du4/j+yV7yaMGYQXndAHGcMEH1U
OoqvvDmN+nVU8j6NIQvQBHaorGgnXCjS1xZP39IveQPKBs6lLYlFoHy9S6euSWMy/M0vD+nr8ZZF
tMAphqoI4rGet2YEfowSXdG5//ZYmbqgIgU/CmyKRjqjL1yBt13U2+H3c+MylCS0MhI7fKH57RlN
b4aRk6nlNbF6plhN6e7SGcvK7yY4atgJy0lyBGRHSlmpAGYOHlsbGLYNDzebjj3sNjg28ryDylT/
syRp0GTaH4sC87CXuwOxviNAHNTCn0Qysw1/thZo/b6YKiGLwso+5WKVKQJUdNEYtds5aSP0fTlp
u7znQdZCPoq4zGsfWtBE7+S6N8XTySLphIMCBBh30mby4OqqURLQYRwSoiZ7GnoV7McKWic7JOcq
zXCBW6xW7duJKX4nS3xm2yXIDp0zS2fZEgJTZuqoZiwL9A6oqHPhBy0lCN/yWlszwD7BK5cjx1MO
hbQOAurwA3kfut+WrwnHe6QOuherAS/VTwDUis2aKbxO/0K6j0NdLuJwnlGIwnHo4otwIxzxjQS5
OvrqtbLzt7Ib6bZGz1Lv7aSpxnt5ucbO7Ut4LmYPBWAmulZ8kfkPkks5Rcwqpx0B4Ou5Glq64kVD
vPJRFk5c5Hl541E6zxhvpIjuO2ZiS1hKA0jzaPf5RKt2AtAsc0Eql5+gdv/bERaaaZ6a3J8lM/zi
hqe5VBtqUCA6S03leg2vwHeWWdzXxX4D/e0obTwC4vH2G5fJr3RShWaL+tBUCY5vDYisxpOvw7pA
AviOtT22N0prKyeFEj4+QVKIiqWAWhQNjbeszMG8wmXZP2iRUhNFJEoBLTI0F7mCkEz1Aoe9D6NL
EXFqvTbP0YQhnBtz9wZd/bOo2gBF/uW73YLGQLSI74znEJgW+gYrrqrSmQw9j21X3jOofwl0B9kH
87R4xERitfKKu/E3xJe2yMTLZ9BVqrx99KOSYBpIQwj2VeHlZpuAs06LXs6FZLrJsi0mg/Wz0YNv
lUI5ivFssAO2iZ32002rLhG+GhanPNX1WvrjT3rkKDhy5eNcBqKPpvvM1wRbtHCOnzRfPL2FuQ72
yJ4AXPdoPmknGfitSURWUbc9CnwDBWKk4WZDm6Su7f8VRVi0uefZA6Gp9KCqmiBittnN18m/2ov6
NwLHoxDrqO2fY6v+flQcjokxuIl1rqjqWcMs5AStI3FNHR/sbt3Peo1uyRzHOtaJ03Da5B/RaDa4
9d7EnAgEEmgCl3LFOd+qQRk7/9vrObVnJit+R4kkbNPOoLxHJEsxbfDVs7pBmUqy3HEbfBycJ4Ku
NIje7AOPk+1hInYK7hDD7Ptwg+77EDcIJFr8TpiFjawkSP+SLIhmWOgCfGSQwMtnq/qyuIXatE7r
rU5j0ReDJddSLtLgsHjECBe6uPgu4Zg9SFsHnNSr7xgYZk3ggLn7cORnjJRE4wMtMCz7PFAitdZ/
/pzDP4r5anRpwh6dC3ua53ZiaRQFcW5X2Hlv1UeC6wtftKVGYmI3/7rEmzw4Y0wr24bR4Ri7EmLr
1fb5cpdLwQ0DuKdD1I00idkLjSJB4pyfgx3kt9I3HIHQ5wqA7I2JtAI0TeMiezcsKAEuIPbbcDdc
1NTm896tlZYIlLB9mpewP2cL8pRVFMaU2cH+vN3/HnLmB1SLYduokz9Y3qhml6SJvtqpbIPPYoJW
SXTXzFGm7WrTwNJltX+W96RyM4GE+8+kpP6O8in4WAjk0mL7n1o0x4sGTZwaaNv29OvHaXDiQHEM
OLkpCzEjEB/HJ/sogJ7K7Nz7gfGkXuYUmjKMUVdV5XIuFRPrBvcZyvnQtcyOjCi3UIPoqHbcoLLt
jglgxoQ6fmph8Ke0/RPW199QVY10VccCubIKyg/4Ro04OTyhoQUBzvYRGhX6y/cMEl6RiYERYlmk
fNXfDJ9pBV7kF9sNVnHU6maZLuvge2sU8i96PBg1I664NPUCuyIl438gqKquVGKwyM0O49liTjaT
HSTKA6yMTLFveWUBlHl5zwcKgy4Y+I9s4RE5NLVuSP2RxNrfttVi89qNLzm/6m33nmj0uOS+DQ8e
ct9oIU2OTUuZQYMEGkngC4Kt6YCwaSOCpqGkJk8ntiDPfBG/eyhAA5at42J7Ca66WQAuyN+RC8iu
MVZuTLMeNhHwVkQcIf5Wb0tkzlU/gjPl95gz44g6u0v8yTn3b02x8Dlv9FDZe+rT+wR+t6QR8RRd
vefjEfVQxn+gPNuwTnH8tsl6J5kKEkZtN1UHqlbx/zVOohb7zbuycxRP4AStM1KY6zcrLRH+OCB3
pSuMKdpeAgttUjC72xBwfAwyUsVZSKLxyuIwjldM3VhiiBORv+Y4rejcc5yXF142474x5wCxEcjN
47onEenskf6mPZRCWg5vuYzTZJMwBPsTXl+XkR27cNvNZbDrK6iACUk7BgdXR2VNCbWaChXeGwEi
sQomOmPm9tAYFQ5MDkU+WS+dJPqHtzvmvsjqiK8lmu/gW/vFq22z7YPMd35tOrPN+/7aj2MxS86A
lywrG2rhNSlx4YVUm0+7TIwicBOyiHnn6m8sIpsOwxqFD2OEiCFCyX9/59x55hVW+CFPnSYoe4qN
ndJKH9I9SjpzkApH0PkiP26YjQjo0AYScREJYOtKBBQyevjZYJ7lC/xZy4FQcKx7S+Qf3NC90CA2
xOXJsaugwhMEQj9ug+TozBkRgIWQVLfBqXpXu3UxXyx7AYzbI2Cb/0R0iLBs9Km4fJod14XyLq38
m9z/hG9V8qzPzLGCrJaRKBmN9Y/+Cgz41LGow4IPm3xSCTuZ5xIk6tgfxcGnuc9yrVQ6mDKcurHM
uQOh76vT1t6OlYU/7EcjMDVTb2XT0mxfod/RcptSPxBiJ8ILIWXubnePaaH0aRDsDZTzO9ZwoBE0
un22fkho9QEeZ+4OVbqm+XAsm7wted3b2XPqQ/KVXc90unSK3ZoD6q3faR4zgVdj00SvUeNSDhOG
PTA/NfUjbVJ3yUKTvpmCPF5oWOosNQ4zoScXt6SLiixoeYbiCYnpudx/p1IFkORhIxfJHnrx3621
yd4Y7yg2P1Hcrpn8OWoNOtbh1lbXQ0RuryeiwQm2msnepQL4yDof0festwjphRCNevMFxAKF3mMR
RNX94ZpjvPdwTjsjF8CRlP9m2/PYG3RWsQRdMab+dJ5Hb3TovgMIRaq4QFVXo+4Mgizf05LjTQ7c
U4KsM45hqmJI4s/YQ5IDFPqJZww/AWShEwNy74fhnb4UxDhGYRVucS2haccslQ5i8ljLX9C5vxLm
IrXxbgaB6r8MTU/sOUZRlBjyR5WN7gj3TDFCndWzaHNnFtZ6su5EFGLZhK07cqN8pXH0kVX4NMhS
RA7BhVqt+GLCnmUm56uKtXk9HE8nirHKCy2eSPl0EJ55GoJDlcIY/IqdLSA+5chqygGb7onOM1zs
Q8MjuV/Nz2QHBA3HoHEMJ8Np4mjbT7ibOb52UPbfBDiTP7YmP+BaKpHMgAMiSo3T6TzaYphncGdH
ZFjj/fh6hGSBQQ2wC/5AcZ/BM7jfY0nTp+33y+jcqPVND9i+2EXoGPbtKfNTO4YCkD/RyCS8iXte
cHcKz0d0HM+5JC/MR0R/qMuih1SA+CCvCPTlYZSIvrQtSbHbZnBhDjSCts15cbjcjstmYiGL4ayU
CM03VMMJTq/h8CvVvPg95d04QG+3JsUjlwpK3iZ4WRUsba/UzfRTLLQjj9vVHrIJesWkMmjoXPwK
Q3m6YAUKWFH21JeZdNM6UQHBt2fu2vXbEnxtU27KBzqK+6IkJgZRNcs+F2Y+nd3P4m07hACTTyg+
JSGNi15rdBh29n8j1aBWjjh98wvukQGbfNF2qF8kBKeParNlPctmoK6FyAGzLr/XO9Zm2rvWmlH4
CFxpbeUOsRfvf0eAXY2DDt/BFDp96yH80wCED4NHB9n1RIaaSnf/DGA2UXBwUUucw+ZKUmi96V9R
M7KtnDkTj6Z2lbseFVgHqxRbe9XH2LBt1hBftGWckxYc27L2qbCHAygLyJJ6/9kTYrkjbBf+fUzS
l7rD/6R4nPriE9G+15A63fL6RCQmblH0Euh5plC/4tqbg8ChTlIGyJc3z+LwDrL0llrbcyiNy0LB
vMxvbakausXAM6EVktubUZV3ZP0QY+ru9G4oHbNoE8c2+bZ2r5odO5bC+eW66Uvmg9vxD5D0GlSv
IpP86AK+NPm+vmQ/+L1wPEwzz8+495kwIn7cbgmjQTc5DeDIXFeyPrV9VAV2a+qxmLoyUpwvct5s
PvpczMljJIXow3MxPnH0btFdT5BI0krpYkW03NzbBcYgIiXjwhdcVQV+TvYiVZDg4+jM3ZpoDerl
AyxQbsFkL9QHmXBEpvlq6DLXD/FbQNLw/VR3HP3Rm5Bh/DppE+znKv20yXm3D52OBJ8m7GcSDNKS
gb7/E5nuDbGYon7ytDz/i4AizEt6+6yolx9YfF/RIZA+Tm5IwdXhxBG08bGD4jogb7jAww+yLyp8
sQESG9MMg/cLrFmNsCwh5nidx1wjHbYGq840LASKr6fS7czUs5CUXLpeMMNIB/x1nuub8aQmDVmK
S0YmiG7sb9GGDhzzmuZTsL+hNbqXlb2pjfqi7PZ+zkudlj0TdMJCh+3bJjuaHmeNa7G3KQ+OzquR
s0TYLr1Ei5VTJObWRU7vtZH87LKkrAtOMFgqSfxjKv6/oL0xq3IOAvACMpyg0NL+70urCmkqQx/a
O9Dp5Y21Xf/vmTKrzf16fnpbotjCMiBuXRCLcVq9abgpeMTZXsYBy/MuSex576Jfs47EHLCiV09Z
hhIlyFZxPKTmTTp19fBpTB9+Wol+JxiNC9gTv1/WL2rQe/4lqRKHGi76J0DW/HyAs+HdwBvtACVS
hQMf+zukAwzYxxVBQdaWgvZfjQ9f18DKxXtLxqWVPvszImXy8zcejVU4sGb7gR2OGPyB8dzKseuQ
lorKkPuwFB9Us2ze0EIKGpZXI4SpFhYQcm3IRdEBCLrpdqG86IVYDOGl2CYdqmJiaBQSaJ7T2W8a
kL2ojeIvpEPXXqThYyU4PeLO/k9N5LPXnTqSat8ry+M+JyaiGaezuQ9TAJQ0qYj5BkbAJxvvr3hT
JOacztXPYgHT67vzRUvU7CvFvJZ2YnOoHqHzKEerTvtpJkCu5IC6DFsNyJms7d8mTFakUswGV5Lb
oClv0Z1Qzcf2s/fs1wmPUb6OkTVLM52MyH7IQYPQB+PFtKWDX3XsOLVxZk7KedTMRJZKaEajH/0F
b5RPiPc9szUZwlu/YE3eS21w35ggUG4pdNM/mRSIs7NksKEZnRrygy1C3RQrg7wSO8R2soEavBVY
3NmXXQ8sk2lkGQqQaL0cFZTW27vJXHA2+I4WnPn0V4UyOZRnFjfUjiM+JL0M+NbJLDv7ZieUpyxI
J90mSOtDmty/hWkN0d3WtHul1QK2vgMc9yWXlsRh5z1esB0dX+dzKz4iivX2Qu/6LOV0XxNg2el6
WbluhdsayfQPdl3C7oZ7HnpEwnkSX8amsEMBCJLXgtJD8XD6cv5waS+sNOVTeum7TJZhmLtKHWKE
Jv5N88esU96NyGVOssS+KvB1t7e/o459Izyzm41F1g1ar8kVAkUxoipOAd/VgDwKH4PLLJoIj7YO
yOpXUxQBT5hncpfDeiGQWGb6nwrzPBw1k5uqlyDmJrYBIH7BZmdgDZ65lBbGOZQFaxNWGDOmeyhh
1Cio9+X1XKDkHDuXfiBw7WYkOfYxM4Rcb4ejjECEjK86l1u1Dj67aHUiEvcy+W60lFLfW5Th5W+O
q3nmST8tM76hG5OTaxqmyo1fLfuu3gq1nFxumLhqyfLLAFPhQMHGPaVhxde2xt1YKj+KI003nYm9
UF3fiHseY1ehKhaEvb5egtbeg/6yB32lR9zA1VqZlz6quF+DiFsiOwKSkXgKXW+TQi3KxmJS06eh
TY0b8KDfCLirx+COgz+wzHVVhxQFp5qMkpNJLIKRy3yLVL3MfdZLe76vfS9Lc//ZlT1TnEpWcYev
kxsng9Gtt2Uy2haeUY7BiXlPHvt06GqNwOqLWj+cUzzWpuvhcj9fp0Mo2/ix6+O3X8wP4oe9wbXk
+bJuBPh07NcTW2iYNZn9XkdoTPD6Pr3gFoK3S47eN7yLrWQ9YwOTFPtSODpmultEYbZa+ECUczn7
0GTTL9mGZN0pomr2yjR3fmSn4XcoLroSLfSGmIRrvwP+kX+LY6PqlZPX+gBZIM6M3xS+B7hBV3tK
yj6E3DEBBgYu+59BuJiTIy/Mfn6fBLb8DdKFcfFMQrUDzs6RD4OMvYlba+y+r2YT4Q122mSRNZXc
zSWkXivzFS2PYJTtrj/4RLMtcVHfVAOAZKH08AXBeri/tqjODS6lHyrqpd8oul/46fM4F6VheSvA
byNQHbxPKpBRkPkBgZWlCVIFCw2waeDk+p4WOM3J39y+iqjq9LdBpoKg/VdGkrgxQ2R4xaHrAest
Y1IyAxy/4oC1Hr758E6PcOSCtnE26EIHXslVyx8PmO8x+KOEkItcpgyIm7UHFU4iN+vZgHe+G0MN
XVjQMhEIxX4ZsAnSV9owj3eZPWeT1fc9z3KsKaXTnfctR7AkmZN76Preeb7T1Q/pVbw3d5qycbFu
iOtojVFBUjkD7adILHvf+M94wb3si+UICK3I37s2NtJ9zkrc7VQdXsYYgU/xVo2BHPptxvkUpOvy
rmQNzGqMhzq0OzBsPLcnkkgqGd2CLYPIm/naNE1hwrxffZMWa3ylPK9Wxc/8qnHDfnnRo8y4hCrW
yrC85h2pO50WTOyh9Di+cn/wmr1R8ZSwkmWuMazy1lWpUZ8JGDaBrL9Hq1wWwzOV9gCGipWblbnH
tYKiax/DMx5o3q/qvmvchGjH/gB/Y+eta/R2ituf2vjGdcRh6iwMy8C8BR8JYuS7MBZJNc2enV5s
B7bEoyTaoJ5Knk8wkeKlkrR72FXpjKpdToBuaiTbMOdsiw2qzhUEAFqbH/bDavHURQ38XCueN83H
bty1o67M0BwsBSTFPMYE15GQf9zhQjzK1aDblXYUjaKCSTlU/pcWZTur7tdsrSS12DUo3LZECYNs
EFmASiHepbOTc9kZyO1JFQ4TmXK8k6fUMLbLlmeKlXqX0C2tWbXDWwBGxuYtQWvEUuz+JqAcTxP0
q+7d+2xnxUEOxwJcWwK3csu5z8mPoGWQgKom3ladXYAPsyxRI25tS8KlfkYLn0aU0bZCBmkpOMsz
tIZMPusfTNeToT2sZZW6A2ZRQueGKkCHXe2hgtoTIACpuHGUotFfQ4hiSlmAv84KhAFg32RjmQRu
mXCU531LmLTk2r2Cs96ayuiJLUcUMX8XjfS6QY89eBea0oErJ4X1Gf/C5rOkMb/o4O9bbZOY2RKf
gAPcPLS/zMx8oV/pO9WlO7kuUMu67NX791uEb0OYjpZ6oyMECTsNrd1eSgYhA/jBqa47+eYj7jgE
RU+MGpoqacMyLO/fYZbgH74tRTBYbd7JrWzLctSK6x52lmtm/+/bxPlyoPOLmDGtW485/ckKVNoD
6YjlPJhqmI5mup5bTK39Ys6AszoukXFNbXJ45fCRjmeiDaeaAz+ETAbiEZ8aXTiE42KMy9qvGsPX
5/qLsPcyQ0+OR1Qqni7dTRuo+Z3mzi+dMLvrfoVW7B9KZX5+SVe6t7JLp4Z/X7EWuFYPSghnlEwN
5dcXYjkLGqllGzH28dN/sm9A3keWPBP9uBm5ifUVXoufpe2LDlqycD7E/MwDbYjZjOr9b4TKDIjx
MswoG8L9qA9t683ZTGiZ7E9/y2tIShA1r9Y4c7nJg+UK9ng1gQszHZfitt47mm4kIWEsYMRGY3sH
7V4XiAcMwR4tCiWHAqZgFqSwLwW0xsq8f4S25QvuDUbnKWt9h1bQ+gzfJDgJYdI9u/h6LJBYG0F3
iGSHiP42E6nVMwjN9eOkvqbjRzd1sCTeuFgqiy63zbuVK13t4YP382LtiMqfkdyOdNyNyy86F4NL
MyQt5BkAkzrcZzQsrQiSC8PcNM+IfrP1OnNrwIyW/c8eaUw3aRNZO0fLwGr8PYmwZm83QQWxtfr1
uAoNntNfPEtR8SSOr4+OOJolxYTWi7OzwCGIrjFAOVdtfxNqjv5eS0etKxuDKgUNdiTccPHfeXfD
SBLzsvLa4R4I51GaJ+i97X6JcT4frfpN5nk+J3E7kajKyRBBMQXNRDRyNbpVQGQE67TfGwOJX6Xn
TGQaJTSC5HXhPthMI85RXKTK4G09jHr8nZBMzN++6nVOhin0aFQiP9C69H3mxro7pgpzt4/1FtcU
jrSUVU7N8GXWGk7kY+RMzOPC3hnTU4D5WbusItCAhPV1Jypneh9+TyOpMuDFIhc0w5rG2qofwMG0
a4nzjvrYblmjBHNVJGr8ailgfDR9cWcRjSAST8NF6gQQOMmB0ywz+7p1D3qsHRM7DiHuyftgQU9J
KHoxBrnW+eUkMc0Jp44ZfLa0HhgbNdHAVLmag2dmYwI9ZZ+LplhkYY6BREatSs+ad6+v6pysoxb1
qo3v+V7sumxUyc5mI7ne9j/Jqvirlvgw1uxO9lxfZuk6dnIeI8MVhkN8/+6mQ9aFsU5yWXHiQjKJ
V/y9xdlEhfRIyZiaVytH7c4sZvDIrfpgvovTKVvs4rSzYkGaZG2eOsnrRKvWDu1v5MeWF/BexZny
1+ARwdJnK+432X0w6GyzkGyzpQZlMalEsprddkFwk9uzjqOFfxmIqz6/Tf3hZoghjq8IWMOELa9A
Vg8bjEAQj+9Miv+VNfjaSWJ35IXv9vZKZZmYPdIRswXXFOlKajKTG1cw8JsXkTzUpGhWmbLrRRd5
Na1npscBNGCfMH2tJQelNwREZoR+juCOFWqIEpRf+Uo1FjT9Q2Loo/8cHLr5kqx95PAo2ZYvBGqV
z9xV2av74o1QnCup3XzJ+GCNDyPJ9fWEcyA9BOei+oPIRSP4HvTntlh4ZatEROXt+71Fd3PqfEAt
E5YlLBybcJaQuvwJLpvdTWbPjaJWRPeag2DX4wpaqLdd8RujljdLeh72gqexKwt7p/0s/jh2VpFI
AYP6LLTViFD253oWaeKaWz6cb/pMRyijm9RPjtL6/IFNSZUkLZ7bY5i9gzzUILnG3WRFJqfz81wx
vyW6FRx8LojB5NdZbiQk/NiFl3gmw0Xfa++F2+lNOyNBxsNImx0I5n0q4CwyXSK+wY92IuGiDntZ
riVPF/STG+WkK3atE9OGyfeanFI0+sh+R6JdbIU1DV/bwFPHJvCPlt4UHDZRcxtyVuzvpaxPZc61
smA21iixr0x9TBDENtSZr2wtRMc5YK4E/7IpFQ6O5VRUUkesWPJSw4VcsC1ukE+3qrRVFSqIvWFn
VfmrHrF2EuYjG9DWdxVcbwfpVEmvk4dOtuuQGpOJt03l95MKWVtQ7C5LlqGU5d9GWxJ3P8+4HyIM
H8YPCmkifLxEQ3Bp6YaGxi+4J0S+26cGf6O32ycQv7exYm0ESTs7dSltJEcf4TWG9cEU0mrT04eP
T5JkI68QGgUaZsbRtz13JI1oMpM/FW9ysv0/qG57atXxPtlaeLWY8F1q9a0qqc/IV/j6/on2p9nH
pgJWXV0klaOu+C8Ttqxw/tGhqCmI50r1bHzehGCe4CpRYdBCPR4wgSsXJYJswxAMwuYc/DvSu2Gx
VjFT/QNjmltkwMAGufmGEMrnAJZsBNlE0qqZeL1gCnY6v6Y0Y5/xRvxVjvQy5lyvEAaZjLqC4xQL
MReGx380xxPaBaDcHdYI4WZgF2TcIqfls0HZbalCXM0QD21lekosO+jKO019hWJcz87MCgh3BsK5
QPsSmLXSNOmbQTNKKt1qqZEF64h8l9InMIvdvkUVK2BWE1ftB5Sy4WCaLmsPNsTYxypd8ZSjQ0rq
E9saKs+xkZkyyjI0MbQKo8sp5uzgWMq5Qa8/JQ7AppxwwpABzeSRUlSusJBWgfN7ZqRPkSsYOl6a
r33BcE++oXl7Gmg1BrBznRN6HPOeqXePr8Xx3Mt7yFMvCYDirQLaKNr2ZQhClIHE62S2X0JlIn2p
XtG+W2v4wym292ht84Zdo4QCwKgkYEjzCqqLx39dLofOLbyztQW2STq76h5FFowH7EHe73kWKIqC
znLh/d+BvRrm32LnuGfMCQvlBAQHCLbDV94rxfWeZfdHT6Fg4v5DCoImU7ETjDQ57Rdx3WBvyOcL
OvYOJatttxWS4GRpX4RcF8nTLdoBoDYHxisvxfGV0SzMkwsGqQGYafMH0TbvQ5iItFl3uhLavPoS
KxoygzXq15K22Z03WhhlngtHHrOVfwKoK9eCCtrvdvG1SiYvawiRE3EEg6lTF5avKGQHAHyQZvt3
5AgkMbPvIglyMroVyVIC8dnGM/vz5Qjzqmday+KKomroiA3TciQuxoz3zrRdQwG7iw6gI0J1DWHL
ZVnwbLfk2ba9E9fyfZ3/1MIJBUzm+ThOsxgUAtKeLpXqd/ETLAAOqwHRdrv/fLJvTMzcsxu7P6zR
Xikg3HoVcf3H1DxByVw/15i9zO1tSV5/gYMo5wNYa7LL2k6al+98y3Vy9oDF2ZrphnSWRDEhv/mu
tPqGYqE/d3kLu1rm7hvNfjr0jjZWgvEg/SIKGRLoHs04Y5xHMONUuSxBG0Znp+5vkF4sZbpwrILj
5VBn2S4BRQyy6vIJd+XE2NCjBxSr4A3YRPH72cUQBq+08L6pXgDsjtRDUQHtrVT144ckcjmTxNdN
ix4K72sQkmAyrtuDjwkogA/uX6AnKgcn7w/U7vEXsPIwv6TNdU37qsMfklSArGy+12ZA2V3c57yN
Tof1yTBRODsJrryvaKM731jiovdWc2Zf4hH6HBj5ZjvWAejghr2byYhimtxmpNRfbw452PBec4BK
OUlyxGd3Qe10qprnQGO9dL2WZxw+h1mctTYLuAPXNsY6uuBxWbtSxiKi++MUXf7v1IbGl1YIqMVg
OL2j79OokkDVodWZpvLQvXL/2+1Y2YwdGhboFfW5E1oNXqMfUUcQqCD+PbsFrWDtkj9Ln5Qgysbb
gI15yXW4RHgmLJcUX53g7GKOOufkuee1ei6mxjx+ABAwuPJ4JkHdMquSYSraVrq1qA/W9uaYuJ8j
l1CCBQjbSf9UUEWW4WX8Uv6QNvLo3+39NaPz16Kq5D1S/3Y88wRID/crTyqgHpTjnqybZkhYWmoi
igHvAiSy8Xe4I2snGIav3yA4R7Tely/I2D4Ur6pj8/IJbRJ+fDgRJHhxCY9RJ/rPoxuUaKVQhJbZ
oMd/t0qSdDhQYJUk+16c9mBNml5jd285sNYE5/2fhUXEHNpcy2WxbKpxWlmzv7B9mAF+8n6D8Q3j
U0FnhDe7dTZPbIy6Ahx8fbbPDUiuhlJ0CcGtGegVsknCOSw3EKl6OH4nV8LKQDLcivJ/p7EgyLmi
GSm9ciDqf6aQLgXDZNCFtW00BK76O7nedv4YR8utcJKY+FsEyUoUSnRKGUf9bhfkg755z+F34JvD
JKwUqK7iaedBvXOG9OA5Mv+jvdig30yOyXFUw6iZsfF2S5chccnXEWH2nGOwdBvulSQGcZOvTqdw
vg75LrxgF+kZak3+JHlkKtiXzGIVS69y62BD+spsCauLOoVNn20d3Ix885D3P8st7eNieBVlPBWF
bH1TH38UBjI8gBpr1qKMmn1/YSFIxPEW+B5eCFurUo95aloS6hhGl5pidZuBlm+RTLNygP44ExNm
lpVoqXM3qIaOUgZWjpmyICWxUMwSmV08HdL1Y2jwgsm69+ib6pfT+yjAVSTmgoBpGy4lsIsusW8a
w4nBDuHHUoZbHpv85xAn0MDJYfy01Qqx7SOUAKguXHOdwvcHJ2n8Ucg1oRFLcOBsJyG+KAyuzBLy
zRjkM1BeW73Xx45VWwHpvAtF5f3Uk3b+RQ0LO/NxhcgVSbQ9kMYai/V/2igsFJLL6VCnPboTeG6G
WfGKkJY1ZT9HjqsR5DPFQ5LFyLowdqPCrLBcklYUr+qgup/RpCqUM3Eg5gRi9EXR8oSc+iF62jCE
6mkDJLURQeC6rfTMrrp87qQdgQpUjU6NrfarXlHbP8X9r2EWi2rsW5b25BST8bzEf0ck5eVPl9KR
i4ujC5A/32w44dCBtN4HhmGgI5dBcSGMAe8HBVaAgO6jyel93B4Wqiozwcrbhv5h+QPseTGdHSkU
jaMSI29OExPlAaU5qdB3rU9ryws1EySzzrA2t9L7iXQ56unbf1sL3Yu+A4IDRCY+bdk3epLZekRB
UZYW46Zqk+b1fvxC1bPwoVQNCPOzeseJgmopF2wT9BkA+aZVlukhOObkCtuetU6af5+i2nwSuDqe
TQ9xlqaS/KpkTbHrfekixjNDFhiEmn/YJ+OJntUb9D+tqS/+Zi1cV3E/IG1s/gaOcvlPtM/+ZtOG
SsB8+9DtZO8l3u8fvmcDdQtT/R8rAzYS5nGZ1CqKXutBJ6eZuokfe7MvurTAI6GEBd12Z8pq0a1i
6Wrks7Krd0A5VwjFwOygDpUP35Q+/HEGT1KmIb1t++tygWFvIrx8Jy6/bWEYy9NzPcAr1/xnUItH
KnbkjH34Qw/ktAYPVVl8xF56RN7DaVYQ8xIxg3ZlYHW6LK/y5xLdL1IZxY+MFupsOuCWriCDNFB3
hjK4NgHsq0EbOhO1MjT88OfwuuD697Vdb0Fz/wWfHct36wfXNO21AfuvnMIrYRsvC/kD+898mMly
c0juvlxn7zyq0u7c4fyStelQwjQDAL87Jr0Y6k/XUmRW56fzfZH8Yh9BTy0C6iI1kksZJONTqo97
UO8QET4emuz36dd+nIBFZt9nk8aNTao1cGkcCq0CHVg709oPzUsJkAJRGh3T7EqDlpdIAjTlP3Ph
yeZxy1X1DN2wvCFg9PSOT6LjigFqc//X4VNUTMW3umvSCm/5Qav/BdvCTHH/aq8xYKk2WHqE7NDs
REJ7wvJIbxN1sWarPJ3Lb+0bdfNzYTgG414HIiiM/32gKxYGd8w86FZUgTEgwZ+V40rP2iQBs3I1
SE/L1MEWxWu0xhM/3OkbCu5U8AuNTVKpebCMv/F0JlPiyDqUuYJMmg3TrjaKbtFn6gNtQv20PfNG
JtqynApIYbgmEAkPO0Ol3H1DGqUlJ5d9byk+vUIwWZIiwZ70pdl9pcUSBrUa6q9I+enNq3fDy+Jw
NM11D4UYXlxmVhBJjOOgM8tPEKq+waaM6VXChiFdLwt7IIRYicAoXDkQ+tGXs8PiY/VXJu0f9H0R
vIbvvV+KHtJJAll/9ih361ehWH6MKinc1WqB2X3HvZE65Vt69O8CJsm7iL9lVn9+mj8WCvM6/YZm
uJ1i4KHusm5miqow65Okyheg2gemrrVg/1eDmoMwOGyY9dtm9kFHHZvwmK+eStvZU8ju43o2F1HO
0DI4YsLe7xsub52dVJkIaNIpYPPrpLWUxbXNd+C0SO3RI6/D03jkNYAXv7EV0fiBFJ9vU53BPanQ
+zNBdWDoxMvt0/e7TddAXy9bwzYiWSKPavUD21pXGVc5DOsmludirdxUp06iGpqgTGtsNnk+pl2l
U64tDFxFqIyzGbcGZkMVbnSQVxSwixlmc0+jyfm3yLF73Qj6m75jd/8B8BpE393Kc1Sl2tc5NP84
hOB8g/vfkyex8CwIU8G28Ie3Cyo9RlVZm2k0tOD2UKG62IIq7Rindi6OwLjZootnf2/B1ofci09a
9I42ty1/bNLdOd890PexJfnlGPnUlcl8kX5qEgukHh+OzSOqNDFtvm1tnQfPiIQ7r2U1c3d7C23d
G0rnXXTBbETNI2KVM6oLyEUP9CJeIwhi8AQII4D290Eiz2drYEPY0Pw5oZfdLPCFr6/qoAdZ5ZzJ
AXtWNz6ji+0pTcJLe7C9WEc9jxOiX3RIE0h/ssM1ilaxW1iLygCZer1o8KullFJSuS9cLKB/6pwD
FfDrtMYQ8lrvF575ohWAYv2BOPPFBw0rQVK5KxYPDPxEnfEpQd5FQmlmctNMHjNIR+YALe9Zou+y
5dUgFmo1T3Z5hbooe6LJZnRLgXWnF36v69IGYEYRczGVoJ06RvHtmVEEUyYJbVcsnrqQryTvFWMq
ixWNeEk4aLpbMiG4nq7kRvKSlMvn7QXX3CZkbj8MniL8BpfynVHYxWxSITHlzfRva+ZtCNRNpP+B
/bjDo6u8dTm/T/Bpgam7Z/IK0i6wrZmOfG1cHc4Yk2C5LxFYwsafU5GgMvJFiwWCB/ga41lkyaWr
fRx9lt0t37G+jD/6Vtzd4ODeVtAdBPaMdzVzE/fZ97NmgxYMFPlHMNu57BznMjhwWKihyVNVVvWr
PDLQYD5Zf3sZvn4sRNHaFz2DvZ3mDuQ5Ux79tvBOsskHTd/94jXIUAsTrnZv7eRvicFFY43VPJo/
D+VEYSXn3J9Xx+VH1ym9XiGiPR290Dl2Q8urfBIOL+ylfwq1L3ZJAol98Gue4mgYIDj/JKboSzLo
vztb501FzzqN9kIfexyf63n8brzcQM2BPc2KN+LQl15Pblp11r+TVdXp85DZhRNddQLtQbYE1Jju
PkUYWH8CQf/db/iZ0TSI//93eI2nIs/NKWzJmjTw3hxpWZLddNwkWDUKYZrMYLvKblsbcmkZc9Pf
c02J7MB2jPDr6Tb/sLP2bFPk2EBOmv6oUri07aNG3he5+wCV06Il9Ab7WX1j+OPn7ZadVidHd7Ao
ra+xb5XZHF5n1g6viTtT+xA/EFZqAyzbf1EguqiaBaAci2iKzhyUbCireMFP+0Ypwy//BaA/B8nl
+Y7pcQkp3OYA4ZfN5pWPBnqSTAYS9AsMRtD910rt8L57kwGjsB7VubvtAYFDK81Pb7yx64t+7obQ
bjLGxN6GP6m4zSGDK8dTPv8ScpAg7LD7XekDJxYdbkFTjXTeHOxCD49N9aJ2ejSzZqwRNn1eilBR
NF5CEWgR7KA6NTQScm4Of5C69YOxVZJ4BquL02sjHViRZM9frECkfDMJk3y7v4KEZQs3VX/cciub
lvGcjNxq7jkDAVDPbdHI68qywJSteo2Z1n/K9Htgw6Ui29qXuigYePg8LMDxVR/gAcQeMJ0MGOt/
F7nOLoVgvovyWZwA/hLxVS7fi0r2jAK7ih1jp9h7rWV9T2P1flMqkaZRyEV0MWTho7nouXtDdwrs
isoBP0uhSKMr/mqh5GjBSHxl19qdgZi8uh456Znyb+RkrepPCLFYDqsDlQaPQSO3GYaa39yvS2Sy
MD//qnD69NECURXQiNZskJnbRLbMn/ERFLWrY6sYmaxM4kx8MaqQ5NF+v473u5PEV7DHGfJhelSJ
AsTr3N8+u/uN8b/iS0acALrHht3ESNSAv7PYT4ucXxS8nVPlACFGKjxs9Km3W5ACw/Avekac4/Ac
vmsGtqnfJqpLPjcjubwWQc26N3IWkyFO89GHPqbvcfWWnlDEGmKRb6vz7DdjXLm0sZFXlFJ/0ix3
o786fMtS+lO6uA6gi3J4StuOv9302lul0vQNdYs1euRclIniB7tiyfxuITw0Xs/i+4XVDYMPiWsl
WyNZAJOXCGWOwdbtTTAEEStnM+PiJ1hxRPvOiL40ykK4ZCrE9/D/oLOvCtm5MKLw5DxtSWEXEmi6
drxA7zQeud8Vg9i2cww9tl36oS4tKIzmXjsIEJSfXZsnIm5HesGzY3y64ZlGT0tLPV//0dYCskT5
55q9zHQ61IKxaY4Ij2sj4CwBmAS9StzW9V0NhPuBNr9dSUTrp24UoNknElBzSz/PeOE4T/FpHaqd
rb9kf2mx+IWIxsRzbvtTBlAqGF/S45MvBFTHptulqFmB148Oesu58mXoqg4eRAlcESk/87WsuY6B
aho8UDfWNZ0kP1yEpQPNM0SA90lJpdw3xwEuuUt6BI444opLJvUgLqeeOpP1vhHnoiqblB7AOluJ
UbtRtleIozKtcZfsDtvhdABC2Tk+8GKqg/mdOPs+y9zlRkGYW8SqF+qk8ZxxtKO4iELOEQ8JbXK8
87gwHxrVSbLJh7plJmcnGHqMEAUlLancmhKqT9fsl4T68m9t/YVRcXW6eTQ8ATdxGS5bwbB8hQnR
8F81gGza3vql2E2PknaQ3u7W13v8FgdKQ4d8dd7WVcGlzMvawXMadCHHnM4D+dzkX8ZfJhQhkCMo
dEaqE75ONgm7F4z92fWkuZU16Ghq4KneeEIQRvKkqXSOg91/UA2LW6vgtDGE7yf1eHHoMiIVMrNm
wBoi9ETJZr70rxLQtkiRRdd3GM94s+YIMAfLVvGM75qgR01tsUfx5rhYU2mQEnQ+hk8pMGur2iYc
ACyOQY9MkiGHsjSH1x0SQ5/Mh0yepC+398wcrXY1Kn9vXTsXPJ5qIuNWNqAmAroowG7d/q73Lg4D
6/dckDY9vQU4pTvckboy3ky4Js8hDKTkFtrZe+L3/dOAcrh64rfSh5pMk6JnE7WeoxePxD/OoNfA
zsGCohsQe7vPKnXei5yThT31eWWSoaPewTICkD1njl2WT+S8uqI4cRQGL/S5xrVrWC+z3m3yEoJQ
prNPSlgfHE7XAaGRAI8ObrFFrWWYbQKELKr0IwNLhDI1UTu+moSHzsW6qgazWuA4AQzYAuASp4pO
hv5bk8ID3WlLGAYjRZtmf7crokLOveWnEYAf/XgXpu22UGIWE5Egp5bafbt5Ai2o9WKeV841My6l
Qe+TVOlmlP7XBKWYdfUPXXD8NggOcvClfnN59eY5splCkUtmzEEytcJsFZAs21QAYhe3gBqOaflt
Kvsfd9Gr9+FmuZWLeyku+Vsu6+nFWDX+MAHKCuBvRdISt47RXoAMMYewl0zSk2V6nAV3QVVIRupq
Gqt+tmMYv0a/CnHj9U6WPb8d3EBw+SGKtIPNoO5itDhGSMVLoX0esxcEucL4mOFNx7rAXJo1qKnu
RfuBD3Uvdcn5tHuBDavitcwdsBshtdieBMZDCz9OStJU1/hs1Vxmb//w5Cmj5Bv2yPSDMZeo08rD
p0hNZ7QQPymDicaKADF27C0EHCrjjX02VgZSbFzMiH3NDHSTsCXyk1CSnKbjAQsqjIAtc8jGfFOo
4mQXOuvJG5e4N8g6hgABdubM2fmhkze11H10U7UJdCg2CrYcrsiG/aY1qMq5ffdFzl/p/Sq7ZTL6
cMixlLie4QaeZWzOuUEZA2r52s0nbZQWBn6JgedoBPCuAlHeY9i8SA3GF9C3vervbD9q9BwFAQUj
rrFx4h8w+eOqHf/68sQv4VKWzRsMk9RcXH5L+Z/zQxyuHTcrdF1xt4fHA6bLPCxFhAZbKz+RGB1o
22vMD4yNC8W3rOkCa2ZIoCCEhRscX/uOkngePJpzJ7Bft0WWY+2agCdqGarEXNKRA4CW0eh/UQez
rwwWoRvPDIhS4D2THVEby35yOyRG4gcNz0P5EzcjOAqm6roZBDxALk22OlcsBMcl6tEEIv7ruOP1
VeffIXhNayPsC5qC8IR7dvBvRXuTs6Vff5FxBfXmZhiOA0SXLZ7YBlYCQOuHXdz8bKRkpQcCEgLM
CG3gZRlMW4vYSWDBxqPv6e8wxAxVj6/aefLMUlNfNELIW3koIA1RCbV0e1gwFRKr73DyDv+d8CMF
aUMbRr/IFpRbzs0X+/VPLNZzss4MXkeZPxKd5pWVdJd2C0PM8ZsGm883V7chQ0l4Xr7EHdLgJC3O
g5/ZcwOUmGAYJdAT7kgddWGnFz5f4Ky2D6RcIwj21Uz+GJ3fi/qLUVkdL4eHU6WDvhSAOFN4cV8a
5fgAbrauYyfslVH1CTRG8wfOSiDad7wCMT2uQIBdN1Q7ucCgPnBF2tylBN7A/qlMEYIbEeeG3FbJ
xxMc4IkaLmUi+f+ZtqzU7/grggB0V+2jpgiTmGEKbbRMzhdO9Lzx6YfBVsGx1W7BnENi/a5ZS4ml
zdaJ0NAw0EEPp7rrxZzuMBxY0YutU+/a7WYWlwpfr6avK6FgQStWAwi6ruZO0z7hDlpn0tD1K5Ae
iP1pU7Czp1WhKbAmgtE8kiZivy08rNTDbjN77XzSejuecSIqCojQ9qwFbaoAusAPmGZn9DrrL9n7
Z8eJiA8s0Fg8vmWvC999C2o7QpvSP6BsTaSkitTQoPIYjk7xlU6y12MI0mxGl/Tec6Qeynl4Oyau
vmV8ppZarmYcu8o7gDKBRKeXmO7phYZ2TdNWC4wKWZAGKa0w6j2W1QvlLBdsj4zZBLrZdL9mD/2R
4KAnp4iQKjA4ghIVJ2aMtJUyoS3NlyhId/3Hy6Sqlw6PEgjPqmwJRG/utIDWA6xD1junyC22fgCp
D7QK0dOl1XrUbvr2axPDU3YhkRdxo0tBIT9EHsY2bk/riTr7A5Kem3NJmdERREdfA9WlabBuxqL7
XpcrXX2COLv4eMzBbciKK9WSrdRUOVF8m0vRTn8DfEyGbPvH+WGWJS91YY2uKusOX9i1jLVQxIxk
6KQKY4BXsRuXPCUGmMYJ5QFXR0/d3jJKuHB4nnDWbQ+SY95m0XbfoDu3eadmAtDdpf76Q+toV54q
uh8QEfa2phP7CtA0vxW7q28aqpeKdjP3LYxHCtESzamupkVAiy03tB6/OdhsUDM8khOFXU5oI2sN
myvQzHdhAy0yGQUgfHmZ/9Q3FJ/Kg1UYPQHEAE74Ck8aI5J/uVprFlD6uGGOiIawiZ9C0D7QpGYG
dnMiNxOeLJ9ZWYJ7uQGyor/eAlEmr12BL+8obTM0ZrfE0WWSgrW8hefTaZr7clskVKxdMoUjgFic
PDdrrMOsj1eTmPbVxk2MA0WzyF5Xj2V5J6wvQL1Rx+QhKp4ryEO2zysqTeSCU3ZGF3q7oo/Z+7yy
D98Hs4431WZtwzqs29LQPfFC6eUk3XO6jMkavwY1bXyR9EuLuLqxQAdSxtlg5dTEm+w9ke74TiId
x2d1+rFpYMjYhuoLbKefXiYPJScE/r9mJwqLPkaLvzgooL5BKPDtZ9WRqG4Nck0LJLDlOCbemSoJ
tmO7orBr6fzvNXaJxkNSGgz9yDMawHAUTaRt5c1hyDQxcHcdtD0kn1WFTjp1RSd/1W/nEIdIwJZ/
olsIgHbpSHS6OvKV+l/76q2QSCksyy7Xcl3jTMScb6Jwk1e1g73uN47qIxHczkfWv3+/F0ZYQojf
dKRV6BFlbdM2mWdJTzrEU6o5osUZ4g6q95AQFpZxlmda9ioUGjzeNggVI/0jhwdYbOjhajTO2+iG
spOpNVYaexrg03qrRZr6JaOeuZIa0pTllL/7G6FLlTODnJYqHNrkUuuAQL7sfoS6A7P2Xc2OOeU8
R5Z7JnWa68qhcZ3FUzZLxdYwWLa3nO+QrQ2/LfVi3BSOBnzEthOzPmRyJShZA0ZzXcCP+OF+OXpN
BqPjLvNg0Tp26OniJ4MZ7PgtItPBtuSAGlupI/eVkChACSWtSmYq/hRpbmPNTeF7e3HZybu28AK4
jLAxCDxlq5epJjJ1yYjjxsuKI8qGrrHN/KAjhTik50amSuC9Oic31zr/5bhGrovOC1Qwh0OUnxQu
CwESE11HRYzDKzwIOescX/GgQ4gBTpdHYEIiFNQOF5ARVy9COoHXH6gJvBJm2TTid/Mic7CFswTA
0lupSXWxzfCc1ixQkbAPb4Zx29+B7ZzPm4VW5ZRWyo/V2qMNvRVQXAwgCZ1fM3OAAmYi9mIFgW02
vLkb01JDoEnvbEuOc+WRie9zDt7y/ebOeJxdF8/9FYI8f05oYGqjao2iWQ7ICNWyF2Jp9cJ+8z0A
cYKeFfUA6vAMBEK5No+LeT9uX09KdGifnYGl+GD4N6fbXkymz37Ofbn57f2wjBKBTS8/SD17ajA/
FCZP5RwsQTjRF8r/ejM1ilDz/21retVd3FvYpJJQbSMfFdl7pLYkTZUYi0mTf8XYsKp22XWumspj
yIj2u8ZuYrM7Q3Azcbb0RUUkOFFkEdiF3H2dpH+z5cg2H3Cwe9tpFmgKtorxXXpBhHTw8hetRjye
6qEyFdbGNORQoM/uAc5gyeRJ229G/VaVxIQHSAvFu+a6G6hrA+iQiaOTaHhuCS4DL0nNmMbdceJV
t4mrfwjzcPnlNrU/v8r6ReiJCHXSpqPRR0V7K09cS9+aTCawcDSqz5uRB8PMTRqbB5ISb9nsOVKC
mHKPGnBNQSUPSoB24f8lswacSRsDd0jqAphjtGRsDJ2uHY/lvI5Z5FgViFTswnKH5bgjrtQRSAhS
G52nqrORN5p3M9DRDoBmRpizBtqqMiQVBs1dNQ6rrqZAG45jwCMxnzBYIwBU8l+ei6FHsx1SixJT
H9CE3myGs8r1pjmSU4BrtH5wQMDWMw5xoPdHOsC24Czs0yerWtRP0qyOdox9KuKsagHb/jbz+onS
CKqA/TljuqZqv7aISzBh8uLhCRRvTmWRwr8Auqgyuic2yHLsP5tXF+3OjmgkXhH7EGEF9pib9mkr
PO4j2mIk7E6X9NgcWKtBJKxajMhawdy4bxwV47Q9rkGfYkrfF08OPXtCd02EGmwPoYTGbbQTYxv5
K3phZ0Mr3ko9VFSQRLZEOAS+pfpK7h6UJXilJykOcTh4dkG0rQpy6y8LCtD6nhMogdJfBgV+2/Oq
2h92DYjkzzKgQT4wnNNe38JmsiTJYZw5ycsVPwbwaj++UY7sGNLzCXGDhuc+IMLYDscEyqXYxgrl
fh+R54EI7N7NBPni8vTN9WC4xJ/Y7BtJc3DMYUiynrHbJTQjjmMmJ6NIsqznFuEYZB6b88iBELom
SwI4ww63cEw7NTtxqoh37cpmCg8Xocipb9mr8xq03tdg27skGvWNNDsiwpvpICpIIKMx3yEPAkVO
cN5IUJ3EOWoFAfWW8r+dE30AxRfHGmysbDt/KXDi8t0C7mKl/SqJg1OUOYggKEfV7mXQRRPzYXbm
IEs19eQCNpeI3zq39FdFRf1JpZD4xMR7eLBA4po4mGHE40uRyuMBj72PvVy53gYChziIxNA76iDf
git1NFqhIDs7xRtGkgyB3r8fdk48Eua1etDLg+tgrCLp9MpeX67RmYLtjiRMsqTm6PSipEPGeD5H
ghrBn8SIj7h5mmcJVJusDjTCzwHi1VmVjOiJJGd3ChNUl5x2bFPsP+az5PcLG5SJ019bjIx4jwPN
KuIaDWumrZjIjBhaChgQz6vlsRI6A4IK373RfYkvXb0oJ2MPeLjCXmCjQ0d0eeqNWWseqSn825T9
TiXpqO6KYC5d0RhjGTqJRiRZfzTK1BfgCF9ZSjJH/2JyhqG+wa10ag9f4pl/wJO3mxHdgjYJwVFZ
Y1zVVPje5r0Z0//4i703KMOmQAWpFG3UOg4ZCRjKn6N9MGR5JjXLDb+BXqnBK5o+RNlAwBpKyu3P
1w35UmsQoRFOSxteGLwj5kkahiInnHolW4CMiB+jw4qW95p1BIziPauNy1x9p0eLArPXVzqDriqF
UesDLbk4CJqMPEEHTdVH+3reU1mOZHPx0G1QOS+UYF4ovjD/PwkRgV6PmsAp5pI6r46ft1X3qPui
lZfPF6Jt8eqU2R+44kGrUi7P+uCRxzJ7HnV/GWGR/yTJfLt/d7ep0v2QK0b5SsSgZ33pHJU0FHXr
23yOIxFS4Nf61LjNG/qSqU3rIwJ9hxE34+q1FePLfle2OHINKJ7ZbW90xFrBlI8SamI8/rjOo0gT
t27tlrjI0jxcNWP6YcJeVhT+/trpDwyO40gFLFOlDAkhUAXrEt8JDEr4guhrEW5dYT9r/Wv6K44v
n5vzdvZlMZBZYyOCIfIG2vMsK0wikrgo450nQQipK2raCesEC7zNGsRPbMa94LYBYPlZI2dd2fNp
JRv1mJq3GmcVcc7vxUbaXa1aWsLrEE2oeV5RJyosE/BSrXFd1d8yPKxIykP9IG/qrgbMLylID2HZ
eylWzFDjupp4HkcRac/xmnLo/ckL+IdqrzDq7PoOqJOh7T/2z3IOBJDHHQvoIh6EIru7BIh/BUCr
eAimRp4txSolhlSly7MFEjibVJ0xV7aX4fxQQhACHz1pIQt8KQb45/FCPD1UxzdZ8LE0XYgq+EB2
Qqx8XsR2UFu2YXkR9R0JUyt2a5mAUxzTRr3D9SfV+1B9SNi/r3vuR9tGrt1RTgDB/8xQZIsmtU+z
S6W/QCGgl73t19FamccAk4QCmqiQczO6cLBFOrvj9SETocwg6VfCaatyc0Lrk3+shq2cqMrauyDo
bmdXDmiVeGF3KBWjU+TWDYHzGA2WuEl3owke2MAMHMSJYJFdEe0iPpNuzRwQxJsy2VjXG5K9qga3
NDOH+T3r2dSmG5tHnsqGb1Nqvc5hV6MDLsLsQK0YWtcmIhzRXkeG0JTTqoSQpYpn6n1nDpsq8Iax
8ngngywR3m3A9z+XHaZVIFI3IoNLQmxQ9gAcLw6S8a5Esl4khelYF3I3Ek9+p+aJkHpvJGfsIv2A
xhYqcliSLUqDIeWP3uneSTchyxVXSM3U8ZoApzAipYuGvnGEkhkZnswSFNebDwnuBrd7xTIKVeM1
lJWpS9KoL3OylGruhAraW2H7V1Ou4dOzIlExOFaDVNjSCFUrtfjiz6HRrqA3P+DG8evOe5GJ9WfK
wEReQtTsM5Sigi2U1A1f8rfdoWldVGzvMWYJnKOT7857vbCM1p6KaW6uIEDCELuFetNtqgIDTc2l
IvKQGvukbYRu8zo2gLEGCMXzqVv5aW23Jp6uGyk1s8P9XqES17pkn8nCYZkCczFW+Lz3Bk1CnXI8
ZbX/QahEmCTAc8lUCHbTROLWME3lmI/tHgzI4OqtPw67JbG/eYRWSrbhfBygovr3aHP0y0x9cRXu
NQ4r1cAZnelHrS963NVf/l5YlGkF8+0vLCyZmg83Vs2yRPKgrGQhCSn/rWLqRWNDvrq3kZTPpJWc
xzy8pJnMusKYyDVHQ/G5apgo4yd/TpH+hdANLCzsXTjMOWzMpH+9xbOXI68DcfF6VMzQ8zijoCx9
HPPn/NGwGmVfFfBdPpjn2nuMGyqz0im/frOK8JdADa5Rh5SmORmO8k57Sq26TiJ/ceD4tRjKFfOr
qJVS8YT+5+4qEXyQ8f2IAbYdCvSkItjWy+ir0ja+L+camanYoWp8RHEiEKrummcguRXAxTTk/g2C
kHnfYthl1lGZAjbJmuNdYwM55Z7qIWL1xJKDApf6tyNM3N9Hst3cxKA7KBP5KYd3/ofIe07QUwqR
30FAkFORsIsEW9hf4dwepvSPTjORCvRYRewXQ369bJNGcGTh0CXmc9MjAdVno7kPRODdF9s3pdSy
XGlZ9nuxomwX8vKT7WFQ1vfHjsLxpbH6iPIUiPLGRtrv/560dsvF9RHQud5NNCB4T7PjsEcW7Kdy
SF835/VBMh+y34rGupfFhJm2nl6wZGyA08sga/5BY8bXQF5gIkMNWyUnnavH5RevSEraDYH4jW+T
1POnSq+4nrmBskGeZdi0aZEcQjJfnfe2MLeif3VfLrkQA+g1u1JHxilheyRrx/saJvPfKB3sJypF
YoMeMHB01s4OcGP06GckGC2g99yp4D2WP9QCRAH0fbgzmjDPP70gu+cCGwiLOD5FhszYhsdiAaBI
CcwLu8tE+NN6Bl9Jh33v6CVMEHt07rrq/ySC5udkpLKBSqvWauIz7xDh/W7QRLvRC47F2pU34f1Z
y3emPKaYtxgLpea/g6q3crWtO/d9YmvYT65x2cG43l3zTqGYQWKjgCMoo/GV0+g0yj4TPnCG12ZT
fYeWaptSWJFgBCpCqUjiTxTNaMclxAGbY0D/muvMG6fXumD6WSYBGhyA3ow5Edbfb/+98UwPOjvz
NXTQdls5sfiH9qKeYbg1SPxUCr2Kps4Hqi/mW3lr1EZkJ+R5d4rchiYXTnK9CLH6AayS4xTTBTAU
JU87S/A1UEmKI7gJBW7alHbOgg1wE1en9yLPyAr2lW5z45enVJmmQnMS9nk8tDWxZd3W3xv/TR4A
+EKVdPn5JFuW1QjI2ohizftrIqy+xuWERAKUzAns9yRFb6DmkI1BTYOYqZmUiMaq0WZ7vPdZSO/E
Mkyhy0GHRw6FtO6lHb+EKz6YCiiYX3RRZ+qNqyZlrTHJgQHpbRLrDXoytr/MQ0TwTUc2hKigg64d
ueeRHOgK/TjsW3pLcq3qZ9Pfl59u1h4L9H76xTTQCFgk6AlFDx7nXtvoHijmtneHLgJlHOXmW8iP
XH/PTxMvQl7gZhpDH58ATb/JOgILJyqgMhtT6aWcY7jncuI3LAPxMAviiGrkmRoCUNAOH38P8K/i
N0X1xtGGxhgXomXPk/gsxCfN+0Cs+KaFpq1fATWATusn+Dl+RaPQT1Rb7qH1S+cTkt0v12ZmkV2c
L3xQntttMj4uYgINmJIQIN1OTJoOFMs+H0wYlU/Bpy3i+rQJS3/72JeXmeDVzb4fUQbJEtDAsLs4
haXiN4+nYww0E77rpUgm9rm17wzKW3F+paCdhJE6pqOR2XpBEOK5K7cHVP3bTwkeQQtNdCeRfVgZ
m/bzQGCH/Qq3BBFFhEiqj6UAOFLQhjjmeJsifr7zevMVVhl413/olPiAJsFDF+TGIPYp7+ntlH2H
RpHDxUIqf3OiGhfgxyHQ6letBO5kjfftJ7s6GIaB166/uUAFdlpR5DIiKCkIkaIRIT9pAcr4cynS
82kwuORUslEYmDrKzlqiGC5lghX6W0RJp82BNJuCiIxscvx4tRJZ/SKwjhH6z3V34x7vhK7JwvJm
/tNBEG9ff/cW46pYBjrXhNfLxrA46gizp5DiQH8hevefA+dcefQy+93goWsRn8uOq1jhWd3J7XYf
D72whJzXJbs7RuU9PeP5sTKsafCKQbGu7iu6qxFGfXHj/4R+A1jlX9j6YWUsSN4scTP6BLB3DsjD
eGECUctxTWvfJIZsAtYKJomUkBVzWo5EE7aV4qZ1puM+9ga9sWA4WeX6Go9O5+fGiPBLUXuw7vPy
k1bVVun4/7Jgau2MiV6ePdWgSVsSqpjKePmpe7pYixAM5GX6c8OtN+f8S2CD63FORB8jM+qvtKTL
MmUGwpdLlBkZ4d6ZUIUQQ+pOy9B9Xqtg0Ji5EO3TgCg6vTaRnPzLAVtqpBb9t70UW/dJ2jrSAPru
yzUAW2Prqe/uYW5p4diWNw2Fc3SivVA+XdRtVHR1AqOoqa/b2UhJn9HKL/YvdAV0fhi5ZkocnVXt
Bxo4OYXyIE6tTGenlMad6dyN7AEInZ82ABgRanAjNwMgGjQysyMllVSg7pyerCAaBkvnnwHKC1Du
cUY2mcInz9pBmqzUgCW4mkzbBIbJ7tSGi33QuW/LK4A2Jix6OmD/NTn0LpEXS6e/hKVsF7VF1VDu
SKabH64815xiCSAjqDZBdT/ogxQIMKVSB86I9aFKodQkMcCAwo7D2TMZ4Depe8ZECzVoXQn91V4y
lBLdKCa6bXJ28ZqNtvFZW09/Drp2R6mnY/eZejpEAImLGq/G4/OPVu7va1SDIkfN+vvNyjpMlTvb
Wc0UecNYn+zxNkejXc56O2BB5UM6bj9tmAN/JSnA/fr13VLOE1WgF38XGNHvmZFhM4HTiesNCzRa
RKz2vdQeIQcjBOcztRLKSrfCGKmtkr2FDdTkur0/xEJYjYwEXI3cI2Zh9KQoN4qsmaBySmMs2BF2
SG1Cva5zMa+6NCy7PJVX78la8ERmAGCJBo3ruQ52AHFkzP98yBxRwsqsDoUYb3ZgUnO53vOLN2uo
FlZ3YG6lQhqwPimRSNUKQbLXchiv3jbenR/xa4Xp6qqH2b0u18OVkeJAIJTWwPxuEu/mqWn6i+BZ
dD87Q10AZQBMJP/trrHUgT5tn5+y6b6ifT9xlz8ne9HAaiqu7bsPyyEvGC2Dn/lwa2uS29MJViZ0
Z/JKbcedcirgQbwUb+hOWGDp/Jkhppz8C38a32yiVnXr5tTiO5U88X+x5E8xgtUZCdwAaPBjDm20
8NPZm/DQ8VzqfKhUtlRuwTfhnA9vttlfzqiPlzKFh+dXoiqXm1ZWqsd2rkPmTYgt8/209bERmRPC
nViNA1hwP+Jz50wLz0l6QtGtkTZmKvZO5//ZMNqboZUG9gl0ayoDK90zGS7tHpGHXhIp8XQyPBVp
vUfiqXPmsOUh+iH/bjCqvdKrVxA+Q5UGPaLcgFIWoj96mdn9io3OrkcI6q88Mj2x+Nnl5qcAppcT
ly0JLDF+ztiqLnoGGDe8a1Kpdiap6iHZE3JRBzOCD6vwoEEzLj4XjvYTq77mv2NKqGky0KUX57Xj
enW63v0VDBzyI04YRuCBM2xfFzEelzVqA+UcVHb4PFJjxE1DoTZDdY+76RGUluyodxgDYqs6pBlw
NMs8BobMylKRBkgkUhKj8VvSJR2ECAhXJbgY65PQVppF3stGwnkXE+fGCtiJnkOVJ75p70BNKLDj
pGH1wHU3M8eBq9wj4NBxqxWOr1/tADEmMnphyD3okFr8JWXlbNSKXhj2uJjo4/lSI9ugXrq0AeX+
N5resHsaHyEqMT+43VKNFCAmBIMsbT23cyjuk8jKGeb6YRrxwBbcYKHKW6Cyilx76e7rgsvTkuV+
I1FL0Jf1lEANfiG6o8OU6LwV1WTWhRrr39BTjnda8fEELWaVmiw40r3Brb8oR6iTordyfqVPobrK
Qm74aClx/VXEMURxOKcA4Kr74qBBeIjIbkoWKr9KNpwBlU/3orEBpp1Ayv4Bvlh0TDVwcGbHYmQ1
CrJ4H1GjUQAScEOnAYkY+dQuTY2Wab6KfS+AtXRJ4gxedRPrsR5ON2IcDg3i78IDGvImrPUNCo3S
wWbiJz5VeTGQ9dIRgOBKjFhIFnzWUglJvEC2byBl2lKPqB8d3MQ4Ed8IoMBG/Sv2qzgT37cUQm52
wwZKcA0hJSyRbG0JeSQ4Za0KFAiL8d2yi583DI01hXoZP5bH3dPS7Xs1qjCZBomj0N2lH/onCFVX
UILYcy6ae4QIqft/GsBdiIzM5bXg8RbJ+unVPn3wB12SHF8lYABhwyXpeXixCAv8f4TGttdj1p2C
q+ZuuIWisaB+f4D4OLdWT7tskGyITciSlFKsoQj00DBva1Hs+i8dH+l625VdNUE5L6GMnb0/GJyJ
6ybeAPO4VVtDRXQctLrpdQHHok3NKzfpqkq8D68EopY03dPF5wjJvnqpM3tbqi2C6PWB1h/cB0Wx
luPuLzT9rNt1uZZC+JvY0CyOU5iVQQYuhyED2rx/FUtjDKCgEHkaklMUoHFIJ/92rHM8WEacCyiA
IuB/bl4AOxPPE8xrRf3m2lT5cPskmBLVGdQe8tQsgTls6dRh0ulKN8iiKz2b12b026eEuLThQEFf
rXiNVnK4evuks+57vjhusVzVNysGhm5M+i2q9mQCGvC/OuOEx53CYNysoji91/zYEldUyG/QwX0E
uE+qxleQj+G4LlfnbgBN1Qu1j52D6gxlfgSP5Btqt2nlZJggzzKfCWtyVEigXxa1M+QvU2fRKwCk
uKvJmjVsBFVutdsyHiWgRhLUK3/aVWBBA7ouzX1GYiBuV88tlUCXNA6rspdiw9TYNvlmZErFKIHM
RB7WdDDhoCdeJdxJ4ZshDkjfiAXspt9A/RxHdmuOIsFybFbDZLtycr28rwPPHLoFAt7ndEH/3Aw5
yoV9Tnt83b/44M9X+A0glsscpmnMxlWq+eguOfMIbqUXrCqTHujapazSjU9WfYiFVuJuZbuznQrk
ehL9xLy2mS7kLyb21BkTn1qj4B+2Vss32gGWu0YdsLMNhKdAHIi7nD2f0gBLbHVCxeuJmv4gTGKV
bdSVClWwCWxLsGN22aLmXWQab0G95NWbhEf7rtA6whH5ptP6DA9E+qyqcDpPqi1H7gouxTsYEU2H
IBNVeApKwQbUhIBGe43lVaAvkAAxjT2e/hspvuBq0lzIyx29HGmVB/iG48S4c3hdLhqyaPg7YFGL
I4MOPIS+pAWl40DknuSqp0DaKI7BOOqsqN67s+kb73gxsEExYSbpJPD4EA+OZJoXVymzOGEj+KSe
a0WK4kNnC5fhw+7ihSthW4Q+6SIKS/ZJqb4gnF/Qu3wkL4KE2rTgb0SjzfiZ1QTvGbHFj5XogLDG
RRcE/T0oP+0Az3OPWAWr/+s3o4xL3O4D2/tk4ezogNQBz8o63bZkkAB9R4VSvNmUc4t6AxCYtan4
zhxn9jMPdCwPAisjvuEKkTUpiiPDLzgiPMCK3f+0fHrTGg+d9K456gliu7aHvxmFKeb6Ardg3rhr
3bJxoSF1aAkbx58LdXFuxo4uGttbDDaPRX+9muzihLHN4A6zwPJ0r+uGzax52bCTAgpJsnAx0irN
DM7Tk9Fx2ZCOIYs4JXmfoVJDhC3AeGw04T2TFj/0kAoTjyTpDr+ScwW8KP9y79Ehd22XzOwwhw4z
a/xpwD8ZgKyWEfoqNN8ZMdgfl2IYSJYU+7myfgC2OSdYpHaLdOvVUNarq9DPZo52Vl/vTBuaKp2a
I1OqYr0qjRy1Rkd+AaQd8/ePm4wIU7jZ7qMHmyr50kBC441KFDEhIntjD132PzlRUisWppD3LCsd
xJ4wEiEo5kaNbh2QsuNVS2gUBpTEJfzYl1dvggFYb5Ub5Ii11SfBycgj8Eeb1qlCGj08E/+IlUMV
43QqEEgOlgmFwQUrpqoz+RDvCfKWanpsoUhf+93LRKvsl3FI+2hYwC7D+5k3SRq0kYqnY9TzSK3Z
6iXuHukvnYPkDlMTSybUJZvqjfyCMoGZX/yS3HCdHRe6a0wZmF4VKLvoD4hwRJvIvpORfNpGUVP0
ddT6MNWkqNfuMvXopKR0aQQHgdzaNAaG8MGJ/ZKCbyAGAT2dS5JqXmAfn0uza8mt7jCEF5ZeCq6b
xMKAxwFSK2p9YWIuGCzrqjK84Sb9ZG9kSB2fhXXFsCvYyUJlqUh7MzlbYpiW9v7ZthHm6W4yZeoh
IVC8CzFzTN+bGEdoObG1HGw+XAAixBBDOwG37UQXG5UGT78uvGCjASxKHlrTZ4oG1Ig3aIxSw2L9
e1EnQ+BlCPr6zK0lXu9KU7jB7NkBUR2ajoDqYmq1GoLixcoxee0cFy1EdrrHJTEE6TFeI7ox2Wgf
keAZ0wxusBBASrnTejsh94RUEzVtZt1vbGX1tJ+3EmUnmbPYxcuBYy6MUJuMpEv5aennrNc6vtJF
RDPwh58rM5cFbmM1pai+DKr5z9eMvM8Neok9xdR+QSPe9xadvetdtAxCBffH1c0prITZZ7tMd/8D
NE+PMdP04QY4bIufwaQM6Mc3nA0DMOS54MHIbrjYCdpH0iZ2z23MKC+/nYkrU3XddD3bShIBuYhi
ja1VjWOh29wSKrHV2j9zJN9Y7CSbM7JSmeg3ik7DhQaI5YDxnZG8ly3cDXG45hNRNCrYk3J7H3Q3
xtQqzYO/+VcIAcKi4SVTGQhiQNPRxRhu+ruOTUYZLkYnqTNjzcx4gy0H1vmfbRRXe+FHGjN61AiM
zuAeiv/Gg6gzFJoNJDvX/5HiHRDusfksbvEs2O4APH5eTP6/sdZZhcEGciSp4Aw30RMHgL/WQ5fq
1SfFtEM0FAqIA86KhiXpY/HKiMzPr4akS3p1BBwJNGA6K1sc8lqdV1etb5Mp8r3vAwamPNR4DEMb
Mp++jQtxkI8t3/eFo/YX2PQvmej8BNvlX9k7P0cr8Vr5zj7vCyi+BxAE5EpB2JX4Y6a9kKDernB+
JeTasD+AXBSUZcaChbPcXz48OIr3GhfA8g02vCndeYBQzal2JzNiB/N1W0UF0LBmkBGDLFR7aCAp
CMdQgbwGFo+3yZtTfXvdlt6HwYHjuESCacSKArYltrgzukOiQ3iXpX7ZyX/yWURl4SfPKSvma6+q
BSPoDj56cruG01fpuaXFaBFzhkF3jgZctv/ExrKLgXrsx7BnlsAMH+v595qFPl4HdDtqLHk729pT
iKUbMQAnaUiuXKz7z51rVMTgfnR0pBNzDj+7V/kVSBZUJpKZ6yU1FH85hWcbRxiRvjrqKwl8GKEE
ksrbBYbwscOd95fjivAarSRzDnBNVR/XNLKaQ0EjSbsxOtRfpYbbSJt+aQb30OBbxUWgdqfGqQPT
4UyT0S53YqBkPxLWVFvodDUG3fsh3VLtG9touFbIjTdBwmS6mvti3+cUBrxP6yqBVQxb+viILHBs
IkfRlWAaQpStod5Pazj6XiejKeTxruTp/1vJvb5YYcLVdtZ2XWznjiRCFLHfzJdicJm8l2gVYNQn
Ey/uGrkSqFJuJ+z+mLOp46zWqO4vXbeQ48jyoBVlhp8/41vMe7NXKUPl/qUdlVMB2tygscktnwkJ
mv0tgrZIgla5mWSKwwGHYnZn7YyYdrarPLzLBh3y2lCThsnEGIZO2kfTh8PDuuXQI4Fr6DuKXnwq
ZGMU/6tukkpj3PTNRCQ5lR81cIY64WCv1ZrsTzbVQURvs2331k+PlTwol1iXHOV85M63Vu+WMFwt
xhhCvjJlqLUAX+UaqvV2fq7gHMLm4QD16oGyXC3UL9o15fRPu/tKCXxg40+ZM6d7m3W1ClWvd4AT
rSHqdDwcjJWsbPAsajfP8Oo8pVDOIPmxYeTg3GCLo0LrswsLNYNK1dUbLdUpBFstkVRhIkMY0N/s
e4mJxqLBPkA6PNNtdmon1g5TULAD1PIP1Wl6GFWCUAG3tyaQBUs/MWNO+jJMS64cIsadNXaNkuS2
KphofxTsOjkI5Q2HszlV8OOhCCNHh74PhTYibdKFSqg3CdfMZJzQLQoBpK28rbc+GU7kYu3CgeJ8
bDcOFhnB0gPdi/OHU0Er9Td+2NpAUUPIbIlw1wxWUbev5K2rPDUsE7Ez+0Gudwbc8QR4bw/OE0J8
zKZTziyBIA+kBlySEIi3Pl574jONeK/bUJPAN4TituKCibUEAsMvCf5nPBWC0K4MX9aOg9lGrFpq
I4JT8al/7RblQnL7OTtUTJRG6975KuVskVkj+SsaYpqbCVBBKhJctam+ogjXHEiBeS/GOinYgHl4
xPLClUWHmcfUEZrFJ4ISGaagZA7dIsqYZxeiTmdVoNRaSGstFNiPaDebFbcKehVDM7fN3Eo8e7Na
eBAJtuyc02Hd8vjOgB6JZOt/H3mIOCRChtv4Gb86eK2Y/kBIV/2yRoervpFOqJt+kyLIETBzeZHy
ZutdxYhcqtYkLZuCDH0MCOT1r+71/yecozBvg2AoO6ECBkzivd4ML51oBdxuA9vpNXT8jzjx2koG
4jOOFkF0fxRxTMxyeOpy3jBDYUCTcEyWHHFigTpKcCKw6KxVOO83yXtiGZdt5Tw9Oqnqbw2x+hDs
JdWSa4lA7wxDSMWxwuRAf7nOOQzFNW0ZzENkWbi2pSg8O1xR9apbwtOPncyDh8RKPBgZIiCHw6ve
NpRvVH9WaMG9HQyc+2Wua789I9Urk9vFbGAFWhfTQbYuswrPfv8J0KX7nhR2WQEuoIH0lvQvLJM6
O9MAIdUGQ3nnx7pI498jLqYO9plCIxUhejvs27lliKNAghJ1idKcrC8YcJLpzOXfCrKUlgwBEHqD
GTKhZh05F5KBnSxwQP85cBdRJUrM3u4dteMj35/S+DRa7qWrVTFQlPRZ4g0hqzHkAqmNstDnLU+z
RkfNVgN3PWn+2/wsjmRKfQHyoglB6A+qYNl0sp0Rf3XquV2eY/IMI5w7qciSCDCyLfjmAr/q/aDz
leKBMBSTIZvvYB/0JFo5HP5+zx7Qcp51gozYNDiGhPTgMqpegFdmcKk1Souat2Ja/ArWre5dp67d
/SEQMkTBvApfR7F8uZkwy3HB3VR7T3sYsgUn0kN5ZQj8OWJfxXARVy5Lv0qgwBl3dUEclVb4MAm1
jMz6QtEIGwv75fs4upLu0nSncbcPTuxUJjd97miPPsHymMK4zsqnMkQ20+FZUeRcrVUcuYvulqVY
o5R89nxag04ufvFYq8cHsOXWLx9SbxMzTrvol7XbQrSDyGtiO1W5a0Win5FKwmUqmI6+YjqLwj64
bxMagUJoxcPHro0K1boJOUe5joaBHY98QQSL++L3HDA6oXphcZrLcvaNwVUYTKDM4H2c0QS0gJZw
JRmH72QFNnnGtZVlkMnn0CNxJkxLtsaKaW/GDdSXCQeMtglbr7risBWFSlL3mH1q/FA8CLiO1OyE
90kabtKX8zqfyMgLeK5Dy7npQcubOr8i4f51UtHHS4vxOza1n6v9up7/sIhmMYb9tQ5l7N/kFQXP
53vyX9YIOJQlU6tRqWBfOmmuQq0XjHRsQI6Ayt9P3+CWo2mQvpZ0pYHdHDIW1mFSU9ES08SYAKme
XRjTvZrk0SOXHyUc+3a605oEwwD8fVWZYSdYsuDcPZWUMPSgz2hrw4WyZI+INGaudVFUxriOpTXa
dyVS1Ea1k16J+OhpophbbJuRFk8y9HLYOaJL4HV7yaok8GNXAs0zfREwG020yWoM/t4LUA4Gr+u5
WbcDpaAllxGcIS0CiFxARsPCINmqp8LL58v+nAbkav9RcHn7NzuC1YhwNw+1OLqH+YjYAwlHjlac
X6TzYAhdBUR3/A03Ho7z3VvHxwVOOWATvjUAFJahn/P0gL7gFTjfJYjmTI0c80YdE+/wEC/4BGvW
fmzUSR5N0Vj+lOOsvnxg3OM1DKXooWRte5BnzBcBvHPf7S4ZiFsAZtHuA1s/hKdCSj/MA5KTN/p1
5LoS5LigBQQsuneKfz9sgctzQVzlWzjJYPcVSI2HETtYLKkIuOEw70YswiE8bzV4/tT5pPbbfd0R
Lx7ptZSmLTzzBuwAFwzrdyRir8FFC9+QsdROPbqBB1TCkFLbdXyJcUay9BIxQABfpePq0dOc1dd+
QkqgY92Y645eFpivjKqinxEZHXZ0fsdwi+0KENp8H6Jk39GAxVskUhQBqyuKyVZ6+TKE2IVUg0zS
yBr++0cp0lteL18UoK25xuvc6TZjvlnYxUnKLiNqhuY9sG1H4xAmYUH5V/sohnRZ9OQFCJx+bL/g
MhL3zy6j5Fwcvh2tLiZMQn1k9YgPf0MsFlSPGsF7PGy5RP4tQVP45omA9KqMZ3MkwC3LTT5Cwngg
Gkz6WxeH0qWdgKmkuvVT/RNoPqbNYcENv9c1LuUAXFv4rMORzrrhS7d+Yzxtxbm+VxRvc70RzEqF
GVZSor1T51HXI/ZgvPLLjGgMQWMpCdQv9p5PXvFP2QkTGAmlCk/dV/2xgdUPyUTEw9rM4OdLE5NZ
OH2qTu5ia00p1xYf6G4eduLrdVPjqVbFY+t4vgaQVAesWyHgFlerHkc79LaiiLIOC9K0CE9xByyJ
ouMxtaB382FEVTLGzVD488LE9l9dKuzcjA3BiL9QIrjkqOrMprhQjIAL9ICXsHxq8JaxOhYB1D8X
Zk85st+PJAJ6PdGXj9P3Amo/5VVzTOIOVSb3Z1pcOx34SiFvbUZQzq1WXspOIrKQ7gVyY7a7XdGE
8ws3aGUnYtWGrGXBpMHnocQj9E2hLgUrzzIxIsvGLVKaktVlhxhyLIv1TnX+C0jjI1Jf2C9C8QQc
41lsq5Usn/o4XEF21Np4r5pvX4rs/BLWgcRBAHJCPbIB0ZrsgK9OPXdRL0F3tButdsJNP0HDVdYn
NLY+F8+2Z9iDihlbWJH0FjzWuCmfY33sOK4cOZKlLEtr5Xmee95CC+2/2xxSiT1r5g51uhtIguzP
AW3x3s5B6eiz7khRrwsPD4CvCk4MYJ71f9XbkCXk4gekJJTOqmK2CMEMxiz/4HivBZj1xdWGF0wK
u4Xk1A9TMWX0XOOTjk4sdRDRRKozNK5WRiS4iNB6xhefLrU4xluu3/Xlpdbi6fradbjF2UqqofIY
+9vPLpq8AvIQWsvkD1sqe5TwKWa/QRcAHGWQsQ0oJ6X2d/zWi99aP8d93uXmHUm1OB+v1Pg39ryP
FfslW3TWM2xoeIQNDg2+XOEQZYeSETZGqCWteu9ybg74tZ1TC8B91FLhMJi838DMwgwXnsDEM4ZI
88gh/HpEsXkC0X+mDLyZWl8Kzm1b5TtvEVlzfCDUPq79arA/ifBt6xtqNNZzhKd10RjkZVck2OJZ
YorR4N284J18TXULMWTxirLEeZA0inJlHzM4Xj1cxK9by78zBqv73sB8P+PswDE+mzloimrAcFWF
DVe0sZgnACw6HQ5P4LtqOFV1jbCfAtPmUnqpmiVNrs9TOMNNrmkD9cfv5jAE1pcRuQjusYd0Wrll
cYSGYaBSOEEOV1ulWQ07icaMMVS8sYB2/aUidBuUsa5pMORwjRciz6oVpzbVOITEWo+U+upvODJI
r3ovO9gBUjGEYaqaaoZ77LOC5uwq/Kk54HhB/CnDXzkGw30moAuFwhGxFjGnrJDbjccSjP+BLfU0
pMO5c0bILlGQLL/OG+vFlRD4jHgndx6/1ttoyy6FIkdeg9YjAdyetSXysnhicLk7jy2o2d2wgJ/n
10EUekiE7PSaCsaStdFU4e2fipgtEzEvt5q6uNRtZhKR8cRDBLZPiGoe1pGLGgsfy7UId9qqrT4Q
RQCpnWinC0XBAm3bBRoEfvV9i2jVikbqUQvwDacSKdLB3esimGaCbR61lBB8cVQsdek2ik6iBv2B
3GGmYQ4u+tSvI3RY6wFQUqzyVTwussVpItMYH8xcPamkz7xd610prsFiUVLcSeMdguSUut3R2+2Q
WBo+cjW/JkbfbH94vjAf6iNB0ntuS6bqpY7TPb5E3C2YJXMpvyA9gMmc13QABjALx/isTX5gV/my
NmnHrdzlGFthIFuzl2fQqyzGKH/oD+SAVr5jHbOi0eBqw9esbbJUFVttbOnkSvQu3U7EQUwxpcDo
FGLhwLKhXUEt2kVW8ouvfEvdlnqQljkjdWm6+SAs20ayfNZ6THiueTz9SdiWthpnrDnC/qnDpQXi
we7GzolyvMUZ9jMmZdOwQNQF7f6JJnno102YJ5B0p1cpsD6ubXphjyVyQOTwzPyOBU14bCK+Fxc5
Bp3Pwdgw9ZyomXwm5dLcHMmoNqful7Q615GtpqmnMIpGnrfm5NRRxlgDCgr/m/J1W8wLffg7gIL0
9PqdlZNDCRl+XiWTF2MofKQ8ZnNzWiqM3G3v+1JBYpIonu1YTCsZM85hnEdYtsPcxrbiuNLpkEoV
9xxUKKEFCrfZrpGEncKNsfss3a841zr1+m+MjwpyI5vyfy2sXS/zohxFlHpjiQLFZ4OomizKmr0r
7v9DxPbOVIi+Q4MZX/Vfiw+daBkSm4tWM5KdSCXXkl1ycz1nJtM4AQQnqJamKqtEAHl18e4o45Wf
07SilmxVyasfms1up4MDBKc6+V2c/6fcCzxYGgw1qDkSLVm7c5YG3EE4C/kV1ee3IeKi4NMXpQmE
HL4hHyKfwU/9OHq28jnsPY8VdVMFxYjaIVP0+iegr3CcvPWa6kYB8x1j65BshuTqSqXt3avSY/uB
8nYv1Qej5jdhAt0oKq1CWtvFA4vznofnbuv5bojv9JJaqh9ytztS2w0G3JhwcdaV3QxmneEicpT9
13o/bKRKQjJW7jwfM4f+J8wXasOuVntz23+8KJOQlPBU4uH7l6hSqNWK4QkuMb68ddQ9ckVBrymO
4a2zmymYujWSufbbSAJ2YjiPp+J9JyUrI2d5zULhptXYxd2CJLPRVo/5jI5nMVekDl0BIUdybLJY
+MryvGVBw/jVh03u0wU2R5irP0LVbvNVVa14r4VoyDdR7Y1it7dsIbddg0vjsfpSJh/cUTwM3uXM
+MAV/nc79UyMQ4pKDty1QPMndMB/mrkOgWCq3sVLuQcu3e6MkUHnIo7pN4CHaMvugOQvC0bGQduo
Nre3iBxlYo6sIj54aVCw7IwnKAezyFrhbFntSUk5yDYwiI9QhP2erPbdJ7p+POHw7jU7smQzQeE2
x+kD13CW8i0/KKRZm18wnCWFuwMyo49EA9nND14qInnRc7du9K9zZ7YBH8UUjlJ8ZHUN1EUNQE32
PPtkdCOggSpbNL+xUiuCNiF9ZhLFC5G9/FMI90EZtTt6/dsQJ/+3LKOgCKsTYePOR/C6q2wzZ3ui
D2DAoV12skKKfPBmUsVoaQ4V3sm2IbbDfvrhqPwb3v1vN0SpNHwXyRBjkZEqRrXeUSs9ZpMDbHTZ
nFe1U0naoQwVP4RuI5GNepax2XS+pT1fud+jYMSiMJGjHf+fPNGZekWnkpf+lr/3Vv6VAWeq+fNy
9NwBb+0tmMAbuaqO9D62uRxFFCKzZggbo67RB6Bgq7KTzu1ZqMyA4PkQVi1blrySPJCuqq/PgEMR
tIKOMFT5NFNVlKzk0mVe9Om/RmQKkZhGKQaGB3GV/Bf1vJEAARCCQMtf88tUqc2g4JmuVDf3TXsx
n8Vzbyzhed2JhJ5nxPNbMtMPenbepaB01hgXJnlpNldfIv9qkMevaKOQ7bqXCIQeuPw3if+xk2mD
66yBIMA4D6Pdp+E9hAzSHQQAgBQFsUE83cucwpcdy0Bt0tdOSK+qTdGKVwIsZFypvka4yaUGiXlD
cIOhW7VvpyVC/eWJhNWGwqBKde3Pj/jAEWZK9iHW8GYYzYoI++jsPDTS6c8h5sGKs2g0398XwofV
uXqLpyBM7Rv2agTt1CKKd7lM6IeaK0YjNWI4PTd4LyodkWETEIeJx3hv68f7TxJGZcHCJeOCj+a5
KOfTNZi+5tlGHCmuUpGCCVM7U2MNFN3nfUALwNNH7CCl+sqfXTDQ6EuIAo/zeoVtyT1hGZGFJz74
VwWbwMzutcWwiRzaZIA7SHYI0FUWKUQd88/L1AEZhA9uJ51CrhU4Xqj30NT18kNWo8o/5Ueo6x40
BO8yM4awKVkBZE37dnABfio+Z3hLhUClsOI9wSghgmuKA38IxiM2bIEM7qXLjrKoUgl5WSNUFF7R
3Bsc8ZrIDoyQYglxZvoFO/kZmpYXc/PCAvkYkpdz4NfnGgDw1XibQDa5hwrTWVJkc7RKn9lK7QiO
5P32cF4mePU0VQFc2xF3vQ/Mi6CzcmqqLEnOqoj3mhANOTDIEhEaB9NlufyNc1Dv0X+/CFEy6FkK
92fAQsH5S/doml6fryvEYJDdglClSH7NiSTQp+1r2ZiCkxHb/S8+MGudmcX4dEPbrujxnFnWwAea
C3G2OEki5X8q+vemJgQjvRSnG5XBPqyHl9xhZxhtNrcyxR+fPEiagrnGMw2q7KqL43wRgZsK9ErQ
EQ8VWc8lz+EsoOJxzyIM75zlDJXx9Lz66oViKZH2k3bvVAcphG2N96ovEu0hqIYaWQvIPTCyo5I5
PMW9b4WqG7BJzX085OgDjzdLfRuKIGMkUcEMhl1QDuwNUCKYlfK90gklvhyHw+xiUOK5lZvaPJk0
nGSOHa9cGVLNuo2ixJ1VD0GV6T49m9aP0q3Cy79EvZpbUOskERVrUzxvhH2nB0aIDXhaTnYUkjJ1
B4qEerFn/8FoS9tVM8zD+d9BMAf5fkpbEdWqU4zdaxoQYuKnGQzh49yS60mjgLufYHjTloZeh09S
l7Ly81kR3OOA55KEJVvtoJ3W662nYL3BbI2NTRpzYsSZBXcAq/Zbpi1rtTNyfHNDAPdcojWRh9P1
vVN8C+dG06E8YSy6gcnsTYB/R7Rt0VI7c0Anbfs48VAomDzAwpsL3L97HtP1405Rd87GKUlnPRDC
xy1Eeky8Mj6l5Qf8d+J1O4PvAlcfDuRZR++QacZGP8jTqXI5KDlwNRgIDZVU1FF3k4EpJLw8r/8C
/Aixh2eYn2GIDSUdLae6rWrI9GjX34Q+XB/r2iVM2IVxNXqsSB/q1IjdswPV1J6JCkhad+mC648n
NuG/iksq+skVFukx1I2p9CDptTaawmFQdAMAbCaEba/cgd9YLGCn72VEl4LspCan1Rp66RGUq5Ia
HkAvDPRWWnflkzSNGXgShIy3+lPa3GZ0gAJIUb0NmlyxA132eqJjDqBByr2zsfOf+CRFTmj21cqz
2TScgl8e3lpRsi80sSltoRtWcZiLRTv9oAMC+n/Uh1N//AOMgXYzY7eSU1eAM2GbZ2KKR56RjVOc
0XLVA6FtN9rcazkf48PYw3jQg1Zlx5y7UG9IXy9afMT+/LyceFy0o5A3IeWgwd0HhVViAFUXHI30
alPHpXGoqfKzPUOH3xGunXRUrNwc1OxtFO2Ep/rQwEFGgxBu22WcDVAlXHfSje3lfT0df3p6/d0q
GINXbKbSo/jmGfjElQ8S9kN6M/iKOwDoF6+ydw4Qul/26WqCJxTpj5KVHdvri3NsdMk/OynJokPb
R59a9jcyD8wfZDcl1dhkFTZO0T+YT1htv4qTdSxESz3cRboAZcpKucPm8vT/LF32QIrgrq6RLgwB
4MM0AjLzZ7/7mgqlqXD5yZPRQgKhw6xqs893q2MxvLRQUapeQYm3N31cvjHVJw3hKTzCTLu5ffND
Z0Giy/wdIbVGy5DRjbD8U/8C3UKxLVt8WnV+ZGM0i5phQNryTL3giUyNCK7A3Rn3BeXzeKqKDI18
WSfQkxdfED4J//UOjXLQ1rODADW+Gbf7haz6RgXrft+dnqpIUM5APKFnitNMpZIaXVvWU4UzNWKx
GQ3pLFRnKxh7yem4JBG9w7fjtgOfNVhdUCK63WjIwIqKjcAuLuGvjwdUAG5tgmRBZhyt4XCak+cp
IpfKhrwB/Nr914SDTXIgXbre8g08ibsbzA9vrCn66RzdT8gkzpL2RUqoOmVJCnfDa6DhHYRfG5vs
mGFqyEu2IC9KGkbgzjacBmRMlMAjH6FJzVxLUuShqOMHEr3ibpw2wt9OkVd2T+U/6taYiacPvSK5
jnmAVARO5s8+b7MG4r+YZRB6nAhRTiaCKU7PW1J2aOsf1QOmhlUFRw1/YQ4qDn68vFxeH5S3Kv/6
hUEwgX28sNFgyuhqpUftyxUkGrCXh8VLwPPEe4f34uEnrK4+aRg6NpdzNcSsTN6m3+T1T4uOomlE
luV/OXHAefIUhj81ClwWnTYrbMW2hzVD9KKBsW8k4hEFHyrGMOqelAycg6PVUS/W2igncp+y/Czk
Glf83BNuS7e0N9ioSB/wOvrLBx6ROaYbZdpjVHsl0bh/Macs5Ebkq58mTElQmGaaBX8fHhiwobjA
s/7uv0wZ5gWoKV8QK1a+KZkk/5KTjqxQ1rj3dalLANYHO7bERx0XIH16uRWyOCqa8wkxuebst7UL
D8q0Tkpfz6YEDZ0jUSmsRRViEOpmkrDcjSNlyEnkUFwnwSOr8FsxBTEZwlAiDnayFrqFhXhJgkJy
La62EiSR8HkyeqKhn6FLtNtQbiFmp9lnFlwLn9YNRkpslvb3LZZ1VRu0AIWIrbbCo9qNsKjI5LrE
nkfOSd/NXC3KpMStj80RruWJxUm7fl8iYsJGHqhLZwU/5aDjB0Gl2RKCRL91Skj1V56G8wZtrR80
u2OPG2uCbTayBzJ27L3ILKd5MROq0whpReDL620utuwZDI1KY4DvX3VNXZbFtPQqv57t4TE72VVE
UY4lapBB37l4cJfQ7w2/PA8dsPEIQ8NxTSJovGBXTjOk71ZKoKl6cpafijEGRBwzY1lo6c+HNyAP
3xCHtfHk8g4KcPHlJ4NKkTMUTLAwR/FW2mpVcKFhXer/O9R2nqTl52pes19zwu98dkFa1ntHebJN
FyPS0bJBgxaXpLR60keF7YCiXcn8A2I88GsTah0+La+4Nu6AOLmCPfJsE29uPj1PfXpqQzaxaa6U
3h700eZzGbKNavBbZ0dm2hUbVaOg8nsdSEx6AsuLQBuViZF8v6oDGAB24m8MnN7E27ubxiitUjXp
ko8fSK7Z31bdKnnWspIEeGg5mrJzNrW8CEZicc5sNHPobDJEpyvMOgJ5uDHTvQB2oNwFaso32OM7
ikbvjpKQraMSPdWKOFv763xeJQLmszeKeq3oNDtNo+/naHzO6sGIM7SgQVBDeMwTbVbSLsre/7If
HPieNGQbDW5nwbUKtHSX8jhdopwT1mWes7TjMGetcs3mJcGhpJL73vxzcGue1BA8pR44N9LA7Kk9
1Ic/aakNDgs1VmwzvEpKnFRLD9TWbZNSOzRu5LzDaP+LVcY5yj+I66BVAGCasw+4XYTJxNZR9KzB
jmyukvex0l2fASlFyXtmDc18tbEGKGRNP9uCCTZ2MJg7o9RzVeSLJU0tH0j0yagNcncEGo3TBe+r
rwj3gqvd0zKZQfYoNrDLW+ZBzqKDBxj4tTQdX1u5FXWtwbm7W8muGsMLBLn1c+3fg23DGwPUNfHS
HymqGxJWc1gsnXnJ7SoT+x0MBFBwYrJKKX6qjmjGO9NxmYS9I4Wt4cZcNJRow6VefKRwMNtYGc86
fzPffs3ICf+4FTl2X7KfYt3qr2do6dTE2CMX6tVnRq5KO2y3qSAcZtleEyIrctq65qELQHfix3rU
6QPvbVAz2rW2sW8FdFfVJF3oTN7Oi2sXNdWh240hxh275C1S0lZqs+qGdwo6++l/TVSz2gU5bBeg
54Ko6eeOyvmCm9vKGP4RgvUTGKrLYf/HmcQ4s0b86wM6Fw586D8BnV4MJl28rBzWZwGeQH4jORf/
AgDhR3y8TYTL4PBVyIZiwh12lmrKPsDsL044uN5Bnj18Y7TioKL0odW3MGHIxnxmISkzsTcop5ZB
YE36H+oa400sAUE8DEO/WobLexz2zwiJRfh0idfPlLIKNrBEk2amMH2eC2WCanJpJD3iUh2upFwh
vCoHulG32Pq27RPnEDSSg4jJXD0Gcu0MDe3Lbh1yaChxwABgT6sLm6xVRtRMj3uNWwM51t0E8JUZ
vo0l6s4mGNXY3LfqEsGJX8lAcRWCfw7iZ4W3fuBzE4cLtu5jaHfxp4yWFHka/0kYgG7FWUh3/pfo
vXd9xaNuxYRzX5GNVffa9uuH2pRJLYCz9/WFp34tDVL7kx3iV/F4BZze0cLGDIEDuyAKKdTBf7hF
BOq1iM9L7vrOUH4gAM6uGefLceKBLHOPwnkpkveSROegQUP+LjMwupMsNCWOwjDc0OWCVczhXZ2x
d64BlBnzq6WtTRoepUjgyHYqd1Fj1ABRdi1aM+KBkLkuU9xLsfeO+ifKPRwIiQnW5GS6mZZXJM8O
/66oagvxpx0D+EKa6wEJmE1zSNXLi0u2+U3cU5wPwwzOYNmQgTDLUhCYiU+49tT20zXgU0sLnPz2
aZVNQ+beZcMMfgIM9e7YIp4+Ij14vFJyI+zKau9MDAGckps0miKH1y6lalyqW7zDxJHcL4opL6qY
Tt4Z+u7Rmnics7B8nio/7o1/66zghF4teeAdsZ7bv6sCofbhALMFsGa36AzkbQ503B/UbhKxIflf
vFculdwJ3dyOKnNaRn5koTJp2i7EZAXXGt9ReHizlSdqMlfxb78Np/gY1Ze/SjJ2k4IYYaJfCTY4
AnR1m/un2Z02v9VD6hgdvi5gUO7YVm8ufH/Qke69dsSsz8lZzTr5NvZokdANVhCXgag6kPBgN8u5
W1h7OmSpUSyAAEqEGG70icOhxLkhG0ERqY3aL8NpxOZ1Lz/SrJqRzQB0k2rRVydRZdWpbdpAcNlE
0eihLfhJvqx7vBiZUyLopzeskQwmfBttElDRvaCpGPYcVNKLUPWojroH8oGJt5PoVZKw8A/ScxnQ
IwCT6fP6F/U3jVdlgktGEQ6cONYtHliQlyhDvTRqka9UJ17MYSGhnRwS/JVgtbPK9Q3Hr7jEsczx
lqFTELOR9IVkKld3LVQ+hMznyDKNWZI7kuN36OvxsMzdyMKw3kLtcunpPy7bGuBgGoULnbMADqs1
KF7rEcEmvGQF0PJmEYGbEghbpJrIAsI/fMvuEmJt+OkIBuzDR8q9wKPoIV4GUu5QwSb+wMvKfKh7
Bl4/ec6oszgsue68tlrNKHRHaz0aw1t+HU+HePWf5NBOCfZzb+NgjJdygOpAIQHh81xDv3jlTo3B
AvEJfSCGm0vy/06JSFj/m+Q+LTvGRrtiKZ9/uefe6lBVVm1kAz4I9pHFuwfSxgjDB0WuCoBLxgzR
dbMwEJOYDlDcXuwhjtl9b141GCMml0GvIbCfLQwFqVwOhGvtXMUJ8AHbSaRDOm955uFi9aKRW3nG
f9B9OGecTkqxlBzctKh+/e3DnmXa+wcbvWAI7ocDvfiq1VSWhTcU1JpWvep6xi8Sfx5hbZB/ligk
zXLBXp/jQ4dxHIHpf0MB3DPkFA9rv3YmEMqilVUXNUjlL0VkqA1TzYun4lryXfich77haJKmL9yv
6I/P2+dzjzFjxdFuLEL4Vbu5lx8PVwJ3mOj6+yJmmsZBJoDROsph5C2lc7U6n+p3WHD8ESFZjk7m
bTqVFLkvTQFD+3Xp9RZnsc2DBntu6kBdylGLtpl1DsbGlSUZlzWnNQS/tXCVhnrSRfSpDsl5vocv
L8z5OZDqBCJTGMM+D/fKbbFjW7WUS/72Y9+JKDTYnJHWTh/Fpn3hmaa2KPTcFrDyiDuasBOX/ep5
mMB8FydEkNWl3iAut0dntlXkkZSxNETbijoTzwGcPFilTSosoy+2mJbnb52lHYi2wqKhKgwOY+l4
QZyEtAW2QCV3Dg93veYZKpq7WMuxveGGM88Zuxqi6CCIlyOvk2y6Z4PEYOCBPBR+1BgZP75j181w
ZUdvHRXTnuTZndn2bduKB4y1dV+1q356gTEggde5ewfA7cf1MaJaE6hF6bxffQbHBImEoQSYV6t4
RtU0sxMJyRDiXgYM/jtZFtFksJWO/9v+Hzpq9M/pHBXLawoO1ztxhsty9AzRivLc0MGLLrcmGWYW
8i0k3xAWjCeu/X5l1dtbsFRrcpob0hfhNF1WEvwlFOO6oHGnAf/Czn0qImoe3+jxVR4ZIJL0vpmG
+Fa7BdTz/A4bNrHoS1IUpElQCMBdtz4AeT/OhqZZao7jedNTEbwDssu3VVvLA51tIXuzmodhOuF5
JYFKlRTzcMOlCgxAKqpCchSIqhlttGGs/8cGwKM1I0FW/Z+RBnHEVZ13yOyYvpZKFY/xmhdllaIj
Bgqx4c5TWHb4dNwNAEwePmF10APZfwywUhGMrVmwOvC/wySUq6cekhSWFuua0f18FIRzd5r/qwWq
l2SMyVtoR/mZPNkk0Vv0DZzOz8QMN5TTIxy4jWRRn9zPw1VpDS9zBa3sk3XXkj5to5XXdHI9ojdu
CJa5RkIu2DnQ8t6GC3xKD3MjJoEIccx2YPparVyuFqobJ0efbFT+jNly1do1ovgv5x0GCmZFb0MR
BMZoS0IIfXfuB9iTXN9DI2R3MsdIgMpm6J31GKCU2+L51Ww2YucYBorqtKL//033LrVUlQhUAiNr
qQW4GPOjHk2XnJpmr15/h7fRtOAhMq3vnK0O49mxL3iMV9YDEXpp4PThW4mfMMERa2NTP5trkk7i
SBndkq7A7l9Kui/fFbnJT5xhuwv1ZTj8SwdV5FTKZEjdWOroQCVJhiDsB4DwVYJBMwaTWqeU8wye
ATXp4SDcB63Kl8+BZhfZDdv6RMci+uDHb9G5oZFTndqDm5TVtPhOKrHOTx0tqE7VgcfD9oityoyy
hwFGd7nhselVOcSv15R/lqq5RUhN0KUOqORdPGq1ikqev2isEHkbsUPIYy21Cwzuy0aaGEgETZph
HEoLQHmbKn3atgmV7iB+jYBz50jzaDp6zL7mFAxVFlf2zRwQchnqXikDPsnlCREA3vKlrwIdt9A5
zdvqNFc7rgNSLpRJViR/T65dm+eVJOy9MWL0xdvExl8axU1xa3soJCxBXBecQR4G2QWhVST0c34M
V3zLwkKzyY02jOTawCjhghOQ3T+KOqk6S305RqWS5Avgudxy3OqQQkrbhBkmKc0eAQ09w1OiUu7B
Jx533ULbMcv1t+OgH5X/8iW8C+HPPJ/SKSuv2cIAL3/Arcsf0ooSSeyd6p4GX9DZB+pjRqJ7iahW
g1bbpb/i+dAgB5fJ67VbzjiKElf7k8J5IOa/5xZMp6F/JhCit5LDFAjLi+MkRGPI0OwMshzYuPLW
pMaqz/CB5jkE6Ab9Bg1s11A5W6485f+N3qoEtm92z/MnfyaTk5q0gWn9FELtq7oJ8akCAWv8p4Ez
mmZg9lMrJCVrH2BLLaKZfifQpoko/G4dM6h5wmod4WaRuaslkR7Gf4LMQkqOH+L0UKBxF3CkGQhR
s0TfVHRoxSgz0YyWzye+NX+Epwno5EchTTRvKmbdZz6GU/rpxhMAc8+ePhGI/TbXr8c3OdQ01Btd
j/naqkh74PPut8b/XpKRLtC5Oo841PkFChYWAgKaGb/eMyOYcNIVjUHDwNVY0GYAs+OSfIScUQDO
prMT2uOn0hjQi42NutmkkwTKGrzCWO3T0bh3aENWOava2zGoQsPRduP1GtJMrD2ZXXgKjiXiV8SG
OnuJct/z4NZrysRU9dPRVEpYrnl4YJ2A5p+XvUnU31SHvsA3TQXBPhq7EiIYXDm5WkpI6ksjKDg5
kp4ii7UwNuldkdl4ojPJVV+rtanM3UFuKO5790++B9xNYNDfyYqe5dbn1RoeKABjeab5Zsre9/bP
m1T+vkQPgTJBXJ2DnNmAQF0tis+1fg+l1N1tNl6ALTsCbIuiBimOTAy+c/O1QFsal/cwj7Ga5O0K
iHFSj/pnour0Vk4UKgr42TdjwD0Qoo+7iUJuqtTF/t71iGs4YX1kOq3hsb2xLTix/UCtB2w5Ehaz
lkkbwoiVQHd9h38TCj36Uk1X4HfddSMAEeofyj0Xrxt07ZfiYDLg03fCQHcsX2uLrWrwne+0LktZ
J+bQS9NuZQngkxYwv9svq2RttbF6/Jm3hiBJ9taWPnhRe2H+vGvuPSfUppP2ID5TO+xAJ1iq18wD
bEDajC+QTgIon4RSWYzRZLckbfEleplvOszE1iMNuVBCGO74zOdn5RrJXFYxH/zUw4Ktp728L0F7
JeOpjUWzlIOhhYqXsEcb/oRGMnndQc696gpB1G99otiEXCKwEZNcptsdXdz2L9pOYdKzCXKtQG7s
druoYsRNKcCiRf7yuYZy/2rE0PPeIhx0A3lQYN/4kg3teq69Pq4a72hQl/E1MXm9PRDqMfPIUmBp
RdQsWWmiHixnZktGrQ6xihtDZyMOwCqU5vVfj9K61+ALTaJwDmGYt7yFFr/3rHAVjXMEjEsr5ubE
Bejckn6qdLGrUiX4TQPPtjYaygOsvi6YaPoVogMohR053UQhukCYzm9DBF6jJUMfoxwKC0JmRElA
ft4TyICpCiFqFO3GVimA4oP9g2Itz8t1kbuMSpEsS/PjzvYc3TuKPEjvZjuROs+o67joCIgttO5G
Bv/HGyIPzw06UC967p84W5cwHbfLrtekznVi3RGv1GL9ifHefbKEtjuBvH6MvdBXyqwUwlngVT+4
CBeclokWRxJWf1NovNMkaZLwwuE21PUlhx7nSTgpUocoQ5CBAFjZrXVRKeBCLOjxHbA2sR4Rjs6K
NQO+qwPFfnWhiWa8UZ2L8YmXnci8QoSFjnGbh/wJTcq84iiQnN0323bzeOdsPKvCYVXHP1Un6fyt
AaFISU8M8gRiPfwdybDwq48Vo08DCOc/Th2V/nH3qzoYA6KkXR6GgTkNCB8wqzDm4pxRU4hP/Ccq
3fBwwRM27TK20H0buIKpmIk3IGNTr/oKnF4iJcA1jcLtrmu3gbmeJdCTpbN89Q0b/vtw09ud0ZP2
TclauNi8XuW9AVQ3Hv6zSPFzih3JKf/NmfUn6kiPJ0PFGIAuPDNJZiT11cSSuL0G5Thlgee6/t9V
FtLGcZVW6fTXBNSleH7GpL3u6C30ASdmD3K0btjL3rDaSFQ34Gy8szIG8NCgNZT+af9EGlMexNVT
8CVagoDTgkInNRikpgOCwkEWYvzUsr4ni749bz+Esjte7a3ozJ3NO4vQttyy8W+FyplKfQFzKM98
8w7SKASfPrJvAUrTfqd4Vy6XvPZ4pVn/tJBDR8YHzBNApgerg5JvFay1oTnvG688ruB2bvhACvAY
JR1cF2roYq8O5JU6mx9ZFE1IEHfDqfWiSR+CHy4HUWHn7ujV5HQ/J8gFd5haGVU5JwjSQB3epjLQ
mRe0EQIZ4iNwhCwpnWfOQBIGndB/BLXChCN93LZRh+5VGsGrkLn2ejxJv//B8jTvio+H13x4Fn2p
C4muzCXITiWS+ZYO55tfjpNZt3DEjE2r1lenIiAk6dpZNX1nLda03sI/1G/lNggc7UXNtyu1LhmL
xkZo/JjwfG89XHt9qiLxl1H7LIJWSipIR6r5xHtbC6yEPuMVdpwDTEIqtGYXGW13wRZcjUCZkJZh
8NDra8uijlaxLeJ/NEGuMaxD9cREpDtvoMZ1y4y91WOl6ceSv3hdpOmoY4+dYKcUCxBr0r4t3IwY
I4HN18K3iK91WK68nskNwA2TMRuV9N2e/mFVl64dWTgcxJV0Vj+ppesu+697+7yx0xhl4VlBpTsT
yBAV4Tg91XxJz7+338ABSFw/fURjXqhRMhPWFi6n+ayPLX2Q7j7Dkn2KfNypGZk3H6/feuonY/E+
rh609K8zqP57R3+EEGrY4mm2Y3wrNvKxhtsK3s+qxrEE8AZc0+funJ0war28PWlHydksvkCoE3i5
aHBhvglsfY2076/K5daVMSo8PN+3IoOZq8BNGyuuj7WEwgwrMC7KdrBDD2fpd5+bWhtShfW+OxQS
ZSTyrzQEm7nMdf4x6edMxkh8dOgNBmPSt3RCCEOHduSXWeJhte5YKnZWxjvv9HutjjzKUJdzCGCV
LJBMXmBEZEeNRlQCirmkhz/7eezGG0V9xzvFwt3pju4NLk+vNUwl163RgMU8ifMT0fkV6clO0rP9
SBTCq8tx8glGa5cEZi3zbQ1gMvcJrsPRkE6H+zG5I7Q2td85TAmNEOLeiEHuAwHGuKS0bxlp1RSi
KPTBsOSH6pqtW8dqunFcNEH60oGJF8EGTQHgo7w0qC0ZnddFgzXmgRm61HwOo8HIjCvvFPDzKvbd
IKA97btAys8thnNLcYFQhdY/IK/GFMREnWysCsEo5LY4cv3aUQHpgnElbZJd642HzDd2PMZGQ0Uz
BVUe6DfXb5Uwn/4f21YYVCEUh+Pbp5+6cyFI+Rg9jnZmKt0oSWkQq/c9glj2fcCVyiBewbSZFsu1
nN0j4oiZQRbCNhfmivsBHmGZ1kL+NwrliBMIe8WqBFpXuUNcHq1zClT/DOGZptrTjwzFsOKPJFo6
I1l9DgstRrFkZtewNKpvfsWWu+FchzTXXGloxI70fXkEPlPOfgQczJLHf/hnKaX0tJLdST5EZk+H
Zpf2JYVACHZpofH2Udd7ETbc1TsPFthn3fphWBMDMZ5Xjz1GFWHT0BHgnJMYA1nTfEMqiX6/VM+1
SLq6lZ5uYbrw2N3babtOTbVbcxh9QMYUMWnnGT8zwmeWMDdmnU5bgBDEiVJx9cdQaxQdsCOnLICN
1O/KNH7XrBiMsIAwJWsY+saIiY95QQB5uqJo/8vn2ZQoVyvvhriA7IOU03vXVKMXl6Bpe6Wgsfmn
2nvdgpZxWoUZmbEdVAusE/NC8AQuDlTcXYMNXlMC7C6bC5RhOX+uKiXrXhnDsa7uYoNH4dghGGFx
9YrhbRCrGGPdp9rYG4p9eW8spieKg7d+TQP/4pbNnc7xN0o/TlaZW2IsuumVbgzExttH0tyGuBhw
6VpS/vz5DM2PiPG4F1nawieZMubqNMIUr7dw7EBKk4kS3No/sIzI8Xc+UyRW7nBYv6B0hk0dl3Vj
qDBCS3UlJCG8i1nLIb6VCLALSIf2xgBWFkIWbBilCG9wes8GGUVueEFwToehDGZfgM5qsDub16XN
19Q4m/OkpqZsZoINBahoGsF+DXqTHjVDXDhkuWUxgDVKXJIXRZqOIUSw6vmzU7qv7cRj/pazzZsd
/13A/MQybW3AxKh5z6wdsdA8Z8x9Q+AXtUlNNxn1k7CGmRBUt0zB9vwOthgtlMueF8qDUWM8axyK
W0xsuaJHOxZbuBQeKwGo/Tv2GCVaJDAvSrQDnc/ZMqCvV8s+63V/SeoZcwCb7CdPSsNonLgELGJk
3bftpfOfeI3YjgUJJ58muQQ8FMKQVGYmEHpZFrwTsNlla39HDDEuiz7FW2dOraamZvtVdmxhKwog
54aADJeEuDFa0LHsA3p7BSsCGYalq8dzahV1WbZWM2flltXo8lK8HnSpJAUuYoBKaHmX7e8fh3g8
iyo4wrIHjqaPISqWi46TfpiAX0yr2qlklXnoutFaBZopjBcgHKeTEUmjXpvBuLHEj4+eLrrzxxnw
wxQyxp9ZgvwxB9mNOy8zgTQ6GaUBc32Z80AuJl1SpWnQqmHmNjG27oNU0GC8zIh/vcYCNvEv8uB3
JfvcKR7uBPFnIQGDZW6IR1Ou2IX0iAd6MFOm0ISc3YxvG/yvxX6uS+niU+Ct/CqLVGBQjPRJB0N1
6MJCRpkVTgPef1LB3jd9zNpx4jilhH+y9r/5xnCwweHTjclweGD4B4yXaIpRktLwc2QtytgFVyk3
lqdCpHObrqjaSIWBfXfsLNXHAGZfPDefl3GljGINO5RjA586Nw0ndhhcV9tp//cpt/1a/i/wACJW
zwyGlURWQqO7GQChMg8GjWRCoX/H6L9+WPekCQG64kR6jjbwaRXsxh2Ovx1ddDbEWjpMgv+w3DUr
31d7yYY1Cg+8x5vlQT8AsPWYUTYTIf5LS1TbD5UIUSOQQvzXWUgINp3m4t5pSpaQ8Ngaz14ZI7N+
JyeN3BcpfRCOcTLvAeusqzjfqtO9B9Lk1FDHS6OuZBHCQ3ZHBCCxefAVVYbcia9+esfyrH8nFYu7
SzRF3v92/XPxOAgi6Xy7nJdTrqUyGlY1+rb5jZc/BttFJ8MTwpHUjf0MnlspZ53sFaxtYXp01Dp4
DoEKvUzUSEedKTHgHKmuJhaNbJJviFRAi3nQ0i/hLUzRqs9klSYpTyviiins/8xHghP80aLSfdng
IRAj8V6gbq4E8ys+IjWyu1X+BS58hDVf+Ta37xIW8Yvg7z7pfoRXaorj/k9DLq+usUekJ8tuHh9f
/J59zHngR5zqy3LsORbMnIf3pTnwHszMv1nUJ+5bFpwZs5jv86MlVOwUlvzRFvRTYG8tuIGi6lZ2
dyTiHy9KsdqmOyLVC5wTWuDq0znY5I5MuA+LyuL640wAezsYvDL5asxBwYlZSkqBsl9Csi8j3DPW
YGxsnC1uedLjYywGtqrrcONeAh0JGHsThkeB25SRdJ/au0NFuECEinBrHB1PAMdL9L2oB2a34uXh
qA+4UQXe/zighVIjK4zeSPJsanXquXMCDAYXhJndiU1B5RlD7YOLcFiP+CLi1G4FIYo4g79sYNwh
j7AE8YPCTFfwy0B4SRx3vHZCjYkwhvmhwDbfBR/gXBk3BXe6b1JjfP48N6kdIeOUeXDpJdzgADKC
92n987zSNnW4hDD2joxt/0s7NXzJ9JqEHndO+Pj6PMKSU95uR9oE2cppS5EZVpEUOZQgQAx7xEdx
GHQDojapryK4mssUwiFHBx27kLojXAIf3djlYRMESZs5IdUZcbwPuyo/yolhAR/C0rpvDRRZ0RDd
1qOrniLnAfN9QOIrjicKCPpQZ2XDLU2rkJYVAXHnP8C6Xk+/Z78xl5Scjpdk5XS9KBaFoFYl+9/g
i0KlZGysybW8enRFZoIUeQqcHaIpe13GH74dZ1AG6OZEtIXHSbuai5dybISPXxQus+lrTxq0f90M
U+YdKnmBSSNTDiIre2TnNMMcS4sTtN37RqlY4KGfFMu4X9H4fvtmv8uWvSaU30kYCT0Xxgbefm/e
JOzMKQQ0LAVt8X0e2ZXGPV3nk1CCDbFHuOgt/dTRdgsT2eqTwMaJlqKTskqZTllw/oSRRN2mozn0
2NXWELwkfi4V9j4bpG8M63QGLN2xGPFtrT7eUkm1mt1lithdyN5VYXTCvU2trLAqChCns9M+ucvZ
6NHOJkuFjTtEd7ztnGXRnX0DxjLHm/c+8Mpw4f4BKbF8AI8erCefga059y0lXFSL/2avv4cks/PJ
IxITTo3AqjVwzVkgvEB2ARToS/xwvdfSqRWTsPHbcFlckzD6lt4Vc85qgQU/JaD7VcRhrJQF+Fpe
+HWKcO6CnM66SvzfbVLu0EFQ0UTPF2XO5Dk1yrpUEzf7Ux7aEN99ycEFPym+Wnq+BiS1EZ+zZDQD
UkoJrwNw0HAqhe63T6FSJ9+mkFjBvPV9ys9W4IkDR2IM9FNSWJCptBJTdt3nY+W8hJwoJ/WFU0Nt
c0jceJn2GUvmzNuGNZvVHPufa88oy33gnBUUybGIAB0j6p6r2sPu3pONBPls7RcvR05gqiOyQ7c+
knchxbtnws8p+ifGwdawsc36+sE63pniWWXfqIQXbQ4YYP94dh2j30CwAE+bfHynauXvcdhEQ25P
/xxaXhuKiM+EeTv3ONkLX/cquX2rB7CKqAxzaZ1/rZC2qwYjvVxA1n9aAinK9naqbHJeDuPHJkWD
a+okv3EzVfwfJ2vqvRx/speWwjpEMHobEtFEG1dbClu24RrgEMhrFAVDqa9XPHU47N1COprAFTql
VEOsE2D2r5ZLu+2ZgcPF1yyECOtFNF31xvhIKUKCGvjVewmLdEO9WU+1YQZEXLZnQUMq1adVDhcq
NDeg5cUQILU/fnRM6+BL35gIPrtpb8wczUpuitD2eysE4nAys/QLsNptaQnzdP5O4jZLNJZE/2Co
94SMGOS6P/N4tlzfiAqWUNPyao/lfW8rpvP8PgoaN2x/L5rhw5Zi9seI5B+ih/BrYpK2su4C1fQ8
4/DtyIcrsBJE8SAGkn89KGhfWNYdHNBkicwEBhZfzwQTaLkO7ykK0kWaZiA14AGYbaWTJSIBUJ83
54mO8SSsTETXS7loJK1iI+BPdZahKDy6eU0jxdwQnDuu5rQvD7CJ1S2bKvuOdludSH75Zqf5w0hy
zw+UifuOAi0aWmMQyHHAYv1axIemmN7eKjK8dw++eLpSK8aGl3pS+6eqE3XDVTX7A55bRr55bmqh
BSHgsIa9nuKUN8pOedHt3uM8NmpHz4rNP4psx8rqxBELH2XyS/Trb+B0QE5Kaky4z3YkdksG7+Ov
8gZQuic8+cPinfMSF+KltvF/IbrhtVn6/FQ+P03UKABzDbW0HBSMHWiM/qonxQrr8mC8pSFgYTtC
oQCGoF8i4hUUPgj9nVTXr1+x/rm7rWxLlr0y4JxuVPicsQkFr2Rus4w6vRo8grlHv7sG2tJJ8ybs
kXxP902anT/wZsUWBKMR0q8+hDrSte8a9mC6BWqWE+fpAHHN1RoJN/T+NE/0g6QA05LHrGieOP7K
6NzEt9ARrWQnSs07nPBJ0ETVfQBoMLxOQ+Ppw5BxeWd0K0UBCpyJyOnMrPlB99Sj7wP3HoKW68QX
76TlICqbFOZLH6wpfjD+IEZEZrNvaBE2CFmt71ATMzI0owPANWTqMd8ihs/IyLT48T3mkCbcC4Ec
VFRK09BZp53f+8thnlepOMWx6/ep7Oi8cLyXfqTf7N4IWzIx/4KAjV3Kf9od19cnO/rSJcSiHQYa
SGmUWM/ReAVqfCMdSDNxNjY9POKDHsCba/8n0n0tU1fKhA3ULAtY2UISIsvpenaE8rTlzmp44Nb3
ghZ1WVPD3Fd/pZzceodMfOTnPwUUGRYQYQWc2az7CvzK/40t2/NRmKKAmrmsQXy4E9oTDMpUnRg5
cOaN4toaScd8CDNF0/OjeYEi8UUyLIca2A1TIoDlgKIypHRD52+KUU6GgALGLkMLAQKYwE3LM1cH
xfGhDto5S8K2e8KBZZcw1p3uHW6dmHMAyNNXzzcERoVm0RASyuXqz00fOViwYyq8jiY5/6loS5Bd
9zW6lpWFvCyu71IhgQ65tiPgocL9//vAAFwDl3DPbE8oAue3O3+R5kpGNdjJ/1SsCFfpeta/kDWD
rBfNetGbw7WCBQKYSOeA2Szv7WsChkgqMQ4jVJ1uqSKwg2AMOr+OopJWg0m3INQbFFvMurkJrywJ
wjABxUNQZsy3jcBtUTXPX+WjnpK0mV9mRObCztTAmwDlqBJdHmsY8JXfFG0Gf6khpzRZZoc/UuBG
XYV2nNTcsGSKF2szSdRAvpnr0gsP/FcRuwnEeFaU+Dn12Vv/iZyx5ZaZmUZ8LCkjWXy7gnmo2Y4R
l03Waf41AZ5TnMqtguZlp2y6lcmA9KYTaSoyu7pAe0wFmzdMF3xsJ+nhZp4V9Ns+kHzqYrZ3hB8k
ZNCmqaqZ098mqzKNG5UPhtoOg4OXEwYeb0i171dYzTZu284S98+vyR4aCg9LZ4DzV+WCQSjDapO8
8sOhUrtkNIxDZYNbXkFL0Acp14bsK3uYIAz4GBhofDM4FQ2KmkHPqGCAxsYWqLDgJmk7Hn+QKW4S
Ma8jxefGkCYMga630Vo911pKeOy7KG1rLNrX4kNYhwpiDON6tNK829THJy87+KOGSZ8tOV12MtqK
XaygyPzBAs893IO2xiKiTm+wLEF5NuHTiYMRS8EfmGS9zqh20/o2Gvt4HGeNkoQZaX85F3SYSWxv
FcBOeWBFXZlzxQYbmv2p0jHklednDIiTnK/v8W3sRLEZUKb1IOtKXRmJVAQH+T9QO1lprKlNSOeT
zwUw/CtACFCzZASWinBNwKUbAD5XZhBDA0N0/ZGcOkSlB9Slg898lLyuePXZZJHk9zdPUwE9krTS
mJorMnPH/t7ajbH4SvngYlfetDRWeUQWNNUi85AUz4DEULFhdI1dTXEJ8yrY6JZQdGN2nSNKwhoU
U2qlXspShbwJ6FSvOuI55Cfj2KKyX4sdlh/af2BBwzWCNL9rhYM5Nf4Y4KqW2G+jr/TygQfhWDwj
2VOjveobWAAfu0RUpaR181cy398QOCLXQbtOqYVd3c7cpNuFC4nGWBOCikoLzDx65wOrRLS5a7tZ
BLdG8a4F1pr5GZVjCznxKuduLPycBk8Mdk+9JbOzjct/NndzvPo7TGq2djS/rk+wafHYgAJiGf0g
NHgNgCA0UVFhv9gyRYhK9CaZLW3orZmR9L+IDPyop13htKdkUao/nS8jz+qATuYg5VB/bcGOkbbW
dh7hCNPwE3UDrJ7aDUR7OZudiPwfd/L4o3Z6o+XnX58pngFK2EOX9rbS4tWsMkA3YVXRWH1AxrkE
BVZobSitcmgx7EfWiVKj2ivfr4+ZbowERBBFEkdSYc0EyA4YF5yKWDMXU0Gw4mXjHWJfVL+Gd1Qk
gTA9iVVcVQ8Pf19K11mTBAep4jPxD76UPAV7pBEiVg516vc8YhZrLD8L3GK1vJWz7dmW2i14jgns
aDIoUeC1JEqfEE5qkSfLJpSmYuSFQq/CBN6MFUwEt/uTngK7uc5vvX8AIL71KWefnNkDTXuBx6xB
hsXR44g3lYrOiPtdi+/qc6nppKxx+BANhWRKWNf0Syvxhy0dku6YRIfmEauCTkxmkEI7KXitNJFi
80H5Cz+QAUJUABVGtL44Z9YLSTqWVPPfi9sOFPvyZkYfB4Oo/ftYVQw2mU3V5ojqCHiwsBXHlpNe
70ejSTvdwGUOprrvmFskuwVIZNPwc7cnQ215hlQu2iJmrLdcm+CIJzkXt4jkXXe4b38z1LdF7iT4
Ii/4Eq/dcu1Rvee3n+2SJ3Q1bgMfZshrAKSDE7sH0kQ27njfnnjBmOZSZyJWKQAKEv7IEqmdGH8k
/uLt0wSHEQ4tlJsOuzushA3/dnOgMZrn9yiRqk1rfsw3Jb0h6btvlYDgdqBf2HmGsUnmgG6Bznc1
hToDPmWWgZwbIOjFhqDOCL7YNRg19gVcP0zTp6hGBvfkWcflSaezfgGcExBix7MA1P+3v0jFyzu3
VI+OmvTRWrQG9S0B+LXttBShWLUYzZ6JQosQc3MedIHpjBKtv/WSnsb2HBYY2cPNIGxPDqHXfrZS
Hh6Q8fPyWofTDboaUKoKEf3V74HWKPS3qmPgCVAoie2D91TgA5APcBqvQU+h7jxtvfT23uAZq0QN
jifyE7IJCmOvOC6HwGQ6Bg5z48fEW8K5LQZBKooYGGVfcOgGqm1xY2TQXn3CCfsbTEIlPRDVn9EW
EZ/u2LJPcfsu8MXVwbFWMEcuFhmQC3Kc8jw+6305g+f5i2uht2LBBCpHcxDwT++382jDskcoLtVf
2IIRW+togL49dw+1er7BgvdXmFLFXhXXVDmRp+TQIIAJUtKnB0L2HbSdTteKCicBieHSTyfBBncQ
FrTj6wlUwDBNuYcA44jNP5Xml38AvxDU/fqZnL+V896CWT7ThNR2YI5UL164eRhBv5q1Pse62DmV
QMQOIyLB9xQ53K18RDIGjPonCZaYEXRErrGjbc/1/Rq9tKumRmWconAVniyl3uICpVr0anw4WpZ+
AAXknma99kZRZCFrx7Syhbwza+JFFQp29TtbllGhapPxUZHo284AydUlEgjpY9YV7fVGmqvTFg7/
9bQ2SlP7lXPnMuDX6o/JLUSuXYrj4KJWU6v50uJt2q+w2JrW8GoVSJW50SonOoWhuKsUVbONouOC
hT2Wjc+ext5xSLr58wQtS2515EmewWhzLGKlGbg9+A/aA+48cwSngH1W4C0RrtXzOW8Ydcm0oeas
bku38hdCXrXNZBQHkxms5gXPWc+Wk2vRfp82frC5IUnaEsuQyPiyJOWrctLInDaskxhDo86RuElo
CM9WtsDGRkTXskvZXhkIJZeoLs9ibVa95eDBUMduGgQQVnQGFAF2aT2QpdhxnszKMm5pbOGcRfUr
8Xe27xmsDntwCAtTWKI9RM02lpW9zyPTe8pVRZX7NDCnOAQ9rmyGL5dKYOnwEl7fiL8wTQWUYjfc
/+NW4oNzIX28fr4mhGyYknTcjhQmzU4FBFvKI4CL7DyN6b2AlahAfaZQBSy7nzkjEXmdeNgzyXg3
H79IesRYzFut08EtRyl+MUKTaFm+6TXVCdZnLIfymxDH1+mmrKPJscWWMEh/4pfiS5Tyt/1NZEei
twkuRB0CtyT0ZHHUZ4EQxQ4IXXrRtMdhwK4EvCTH2JCREBX/gaBTJtuw1JMaU6eLFV+LqoqP26GS
3DZhpmu8pt/HBjilHrTxiyg5XQ0seftuTTsUCDDvu8Xk8lIcDdIB5VyMJ/X3Oypvu3Iyu6Q4WiNn
GLhO2I5oKnaTdDDzjHYu6M/6sEXFoyLAXlUkql6bEjj3BhjMGP6GZKo493DM5OJn5mxMnpA5qPJP
ukj0prjqxbU1BVGr9qtDueAHJObH/+QI6FTJUOLF7GJuv5rZ3IZtmueb71flrYY1JoPMT9w5iHxU
IBIeshZyRmU2iddfphAChrjm9Prhj9LYcH0GmtYltfE+jlVADPfJf+ZxNfOEeb04etSyCoAtAOPg
QyFyRRRek1jvsqdCSpxYiMU9nQoO7R2zHXKopODvg9ZzVS5oXxFDHrzQ+nZWGwoqKc5xD4HQZrGq
cq3aMJLeC07zRHqi4tEWYOR8C8tkW7CLJTTt8qd6Nv4TaSZGt+j/FLG16OTrkKdNBC04KPecZdKD
w1ZsadbT620zLvLBsCGVr+PmFWKeXdKdVP4a7Jt+/I8qSx2MZAhvwxwRI9eKasFGi7LRcb6jp4EO
5qH7xZI9A6ELBmdX3RTxlYxFXUx6+eC9PJSqVQ9z4JJ1LOGrGyKjGgu/ozeKWUOFw4R9bVuP2fP4
rUY4gm8KGQ8n7YTC4QiESg7FKhnLoCVO/ElPdcPGCk+HFO8pm5e2u0PbSzd5tURS+8xKf7hpzJ16
N+/EbhhbR7Iky9oCOUeG8h0B+PgJWpwpXlsRrEAUqr6FjmO9/EsrfPlaypbIR1FloZUlEWnSmQtH
F9yC0GMawqWv5257Jux4Jik6WbTBt/dNuq1geRWS499MzNPncQmeBOKtOvR9kb/pGMRVPWF/fHFp
fy5oRNFtoRg02WcYmOtoQFbtK6pqjOOGAPDHouDkpu8AIqERi3goFVBXgK4eEDNUWI5AsY3VP1wa
Ex75F598Y7Dj3dq4lru3lHNtIlZzYZSBszUGy/t4Jypl7vERSVmjmlc9Zfr2085V87eKvM3I0Txd
hZiLMR2AMcPMMsbwKi0M9n42rFz/KC512mrFzVEZ/zURzZR02OevfKbyGy1zwiUD2mPqhrPMkYcX
u9sEhuDayo1Dm8Lfn1PMmq+HadHzDRMMyeARNfEVz62yeLWAqpkeCIEpEgok1WQ5CZ5mqdKAhhWi
jW7wfnoy/UEp6YHKvaFiLfI/3rJ6uAOvtuSJfaanNLS0lgCtGPudppOxeH+m0kGLAii2Kfq2TjL8
5RRknTZWdZLB/vVWSfbUruzbGbBqqBlfES6m/voLzQE5Wv7FU3/e/5JJcyD9WqrB1j/EtPWVLfTM
WPZRDUD14ktLjalOTFN3Yk/gZWaHszZAJc7PQZHbYgiJ8MCGXhmBROk0QqHHpR2QMT6WyX9O5XvN
T8jrWFdyjoJCDK+PjXB3mzkCgSrj62vaJkfFhTRY5V6w3axYCvnLWb+I4/aauAlCuoURC+hucpKy
tKX2lptId+WejT5IGrNXaL/tswsWO1H9zsx/UdBujLp/DG9o5FfpuKUn2H/ILyP9MSGU50CwnLV0
WLMxCM9qHkDE/9oO7BgwuNH6JURO8e71C8Y6G2PhUzHWt+1kJjpd/J2ch0jTuqQcRMapGCxHpDDk
ZwFLEzgyN1/Ryy8LWfIvBz9jSpYUSjsjz6AxIjs2MJgBX97+saixNBA5zLcQai/TFEzXOQ6zTNxU
HJQQne0E4BLxuoezDhYEQcuvfR38S6r4o8e7TrEAfHrAq/5NgTWGx54TlH87nFW8Wy4JSZKqxAfY
manvdpjJgxHbYibBpDadyAWE+X0HZ9Sp+mIb3mY2J1K1UjaZAiR2s7zZUTcS6uxF8MX+hv7/OhI7
ACSzvTEwHpKgv++4ZxG8i8fWIst8oPf4lfgK3d7PCOSD4DXRV9g7DggUYZbADs6nCNVi5O58k1rn
SihrHd8xylEECp+G0pk8ZQ912HsF+Arec36WdF46bSxe3N5d3lrepm4u15c37QRvWYyDlKqNEIpg
7KVO0u/C5xZgjKVmUaXsLxHorMa2+FN49AZQdHR40zCyHU680lZDmM6lHawbRgQXAVdH1fjbBDLW
qTCbTfico+kNVxQ1sdwjbcebOojK7RpLA7iIXkMkpsW9GYpsTk4UwmP7R+kUCPAVfB2vTnhRAabM
X+skkrfzxvFH53CJIMN2px0Eeos11ttmwTbrVD+RLHae4bxD+LY4z+kVj29EbULAyyfb8NKI0IpI
aJBvDQbbv5Agz1Gv4mHzchPQrorBwjDYCtvhvULT2XjH2u+KgsTgHXNzIdDx71hkVA69zacVoQyG
vMja5N9Q3/J1SQYmcqF6NHyU7rPpdVNTK8ThaMFI7wkqn5i8GXXnxhoooD/OLK4Z9emxb/57c9k8
msqnyOmHVgugbheEBBgfxWQ1skjYkyKPe/2okNk+bVLEqO9jFkvp2gMLEUx5POGwXb0AGK1iU9yP
+x5IVw2ty+zBVPvpmfegxsW6P0O6Oxgk+e1u4MfbWX7cUickjDVZl2/5DPnr25piI7vQkCjA/xyA
SNqsQWZUkrhUocofpQgIRLLUMYYHO9EHchvymasGwcxxWK2w0HxX9eoWggEyVYLn6E1Zl69uLUNj
5RY0xRuBrtbBK4nsW98RhxjGVXaNxf+MJSA/CYGlqd6KR3G5CX9e+jfd2oJjNOdZGxiZLYGckX3w
9GHTPWVD9Zvh79rl+MjFJjY2wk6CW5zIc3CzM7NIZ5u18CSugDZ8wj+s2fwGdyG+CysBB4ePFr8P
0/S3J7Kna5eH1m/cgnTfo/bpISwKptq1ofjQBkBYt+UyDYrplwm7wuSVVV7Kj4C4sI3htlemo871
/dq6DJaD3scg73eFs6jdcMoEumCHVFPp15nlz6UBHks6TldDU+5uJhSUUJqF2PEZLDc1UK/Ou0lP
hkzddUEs7X8/fQZLOGqU643c23ZKfZAuqUtl+IUShDz0Jc9n7u9Jr528LZtlOHJ5oT3xv9Hdcerj
sRZRN3uHmTwot8xgS5LeTnk5S8md3Pndk1D7q00Nz2oiPfWBUwdV8L1aZQzY8y8pDVH6nA+LUus3
LeMi67/pw9jHTRJz/Mb9+ggcqq7p2L+8L+lfwluKk8ix+cHcaPDptFFAjzJuFqfxWyX0cwNFI8eM
s1KY1E5t/jap8noyVqw2oHmvy3bCCnnFqiPsHcxwQujJ0XpGh3nGQ6VhVEjHAG+ZE4q7sn+6flPW
AZG8ay/tjsP4MhETRR/EiBkOXyovqbJDk76wVUvGLEv73UnZZbVDf90UnA83oWO36o+Y4y+lsjgR
sBLiHs3/12Em7DP9memla8Vh96MFxB8/Wjoh2HHyc2Ous7fwiO1Fe3rMXJI/tu4GKT1LrBnfBju8
jwvVy/eV+MQmGeLLJ/wAvkVOxat79VLH6VjZC7uHi6Sqs21GxNwFM9PicAeN+UB0j+anK9D7R4Og
kBruR9VGPsnnnZHkQRqzDcuxwocYS+S0HVewGeUD+F8J24iLngPbhSgAeQde+FKhjHXbMJkyC8dS
94DqeJJb2K8PUWtMYKmEcW19nnCzlsH9z4Ya8QJhLO9bSFrjQICGlCO3zsSTizhS/49CoAJnE0c1
zWVmhDVBV846XDv/mLR8+dUm6f5lE1IMhlh6dh68uU8tWtFNkL1Q8+ktdJxhaLnbAIF3k4EZl2eg
71mvlUzeda8MrT9cKQBvlnsWD67R/tnnudyrnHjgXVBgTyV7HjSjmLhmrvU78vJBhZZxCS8KB0NQ
MiBroNeyyvogvGIn5/9hTpWwkcNoJe6/Z/ri+cq8Qx/Hr3aUpy4Qz+YXHDsbeEJ7QyFXNuFdxxFS
FhL7RqTmBwR/cmNEUnXi0YMD73TpK9X+w+m/LxEa7sfHDOHefhM8vEbLEgVjEo4DEHhcZTQWSTEe
wFKIRwQ6Nv8kANmoJBzhOuzsWMNvEuHu0zuAzaTmqFceHD3t8gwZfklVgkTRRnNYG57WTRI3amcV
B+zDxxuhFkZoCEBQ2bsmzMpPC2klrjRNro27YtydkCZ9u6sfER/Z0+p1A554Dxd9D5NAHgyhzIq8
zHeTAAuxmPe9I2jgowKwfaQf1yU38DCq681+dWZbN3hXNoqZ/DFhEb4v18oPqHj5IbDo9HbxeNkk
9vY1ZJKMwwWg3P399gr3GoLMwxCiI0uz9YKIXvvVZhYOQCGMwCMp9i+a7Ntdo+bnfsNcuSbHOG4T
05k+Xl+zpZfHSXIRq6KEqjntY2KWIUA6pS00nGCf52XlpG9KhqCBvapcQ7rl8PQY3du5FfrFdvvM
P0AlBKdtlPeKnQ/zO9BwBQhp1OK+MyMlEZjhZYmQw38UBcTlGGgBBkoYZIhdq0w0gLT1W2sMB/Ue
QyEZCGqeRVwYRiLFwe/Ws1WVXV5SzgYeXMlD+ExSsRmYNWndOyVaDFu7u8K7Chb09h8S3BFo+VOG
a88RjFQsx4B0EnBt6i0bCw7B2wDaVzZ45tOfabOQ719lIbjfoOyK+pJ0j39wggrtCPogl/da7lJc
T7+mZcbpZSxwHOxXmrAcDey0XzCtLuUKqiCJjQ/maVY1vg5Z9f5X3l9If7VEqkDXRkl7tS4a104U
EO/xssQM9wCJOINbZg2UvV8+j/6d0zc9CccHdpj3RCGmE6S5sBUTUsOYxM9u4v+/u6qXnz8tRMWt
SVrzU0NaP6HeaW7lm+wgYmz2IOg5F0GHlmsMfLXRG4p1BlapKcVWw92LIjlIYGEMeS05Ta+AP7kv
bSZbLizIqT/97QP16NhZerIBwCaIrfU2yxlzJ6LNqMLAUHJB73mQxZY/e4nV4hnuDNI7mxWgHeoY
vvXe/Fc3gBpmMKi/fFIu2DSU/euocEeKke4YzeFWyrvqqVStWF3oPN+O74b6DCqzj2b0qK0EjSyl
u88SYs7V5nBw786ftpQg88/anuVIIKuAFJk9qF82VcJrnZMfX5qrW+h9V1I3qlyMlmyegLl/h0rI
Q5fBa98GPO+h3cZ227v8cB52zFpd3wtaIJiEOBp8Dp9ZgO0EfLVqQ4PMH+Etmu1dXiJdGL8yr7L6
JqtFzF4PId/Nv/gVH8JovyiW64NYCOBaFLQ0yhVqZYqLf24Aa58/tuk+emH6mYyEdUaGYLykEJ8o
dC0gfAKFaB2E3tdWFwKBkCi7zTBk3LpGFsw+HHb+rXOe/9/D0hh+eUHb6vOha0P4A1J0tRsGdSNE
esMTKok9CG0nH+UryyFM8MCjhLbXGjYQ9V4vkvnOYwO5WtfNmbm7WH8ySZdsbQyRT0oe/D6zGv/Z
y82kxWnR8bO9tGMwFJveDyjx16m+saoZS4HiUGFIYUBMVU+3elL2kZStc3FM1lwcmX8NK21Zb8Ib
n2bcVMACXOoORnrxlK1BUJaWdQXTe45SqulnptWgcOhhLwgX34OUi7J5LDo8+N23zUXkk/Ei3uGW
E73eEEbVlIzc3ueTi743ciI3QCb4NLXCf6fRtlmEPOhwvmBfExPpiZzTdf8jISoORRVuwngSWl0b
J8SD0gH9Ob4xPWH9MrQen1WYu0io2++7ta+DNvp4jK99hEaCTDsh5+Yd7JbzHIM1ebJHgUZ+lKuV
Z3WDPsRLuGWKzyaNp8hRI4jVB1Bidk9JZ9+DlxXQtq8bGiTCmw7bMQxS+SXa9k2dxC8eVdyErumu
FFH8E5uFsmeNS2Be/zP70iPhfnMRVQvkQeaS8kH65+VCWy44ZwXaM7td/sH5p8dHz/1Zm0WhxQ6I
uZ2EwlIF9U80nNtOif/Oh52+WlKt7rzd0lAKaPzw/ab4dwQsf55PdE9SBHWi/mCXHmRhfyAG0dM3
H7rQjO9PWFYWgAWgcckJJdBu4FYZMvsswdsXx9Gy1VirVYXipgDWaBCZrNZwMctr7TS0p9XmujbZ
8GmCQtK2cv/fpCxmM+U+jzljjnM0C+sTULn6BhgRIQW7c6z4Zd0P89YigR5TRFZWLziP1GLGpC84
FAWrdb7sxzK7kTOqX8ch40o/tZGCbGr5OEiR2Vwr16PqzWIeR/2SHIJ8cFS2Cmy4RCYblPe58jYO
03+KH+qboBHHwC5t5sF6JulVmelb2RgyUBWsPwMf5nlbdqiawryPVOHLqPPZA94Pqd6hKv91kmff
XPalLrYpR1lBWIMtS43EiFgHyDAoGH/p+su+xoPTuxhUe2o7OhyUIbxyGgDYQYDiCR63pIVJlIZk
IYPBfaQZa6zu6WSegHf/IOpTunL9DgS2/4z5xkxCvvy+fyd56RNzACXoDzQd2nvICKvVusfcYe6g
Zata4BQ7AKLqPLcRiw/slEZ29tcu9Ij8/bbkkRM/mdJeUUjy7Q8TweaF4SW4hRLPQTBRY84ZW3wc
2HFABHC/x8Z5kLHwLC3wc3jwhhXPNwXWIgC9tyR1594PLtjjCR3RjuW5xYbBcTO0M4eyxrizDSzW
DopjeYSIHSzkjbObVqk/FgIq9UasxKkOUOciuNrpbN2nHY9HSlN/kSqKG1VqQ7iEWfXVdUoHT3nY
jrpAsJDbVVmAtbulA6BkxKua6tSSIVVFVnDUnzOKYZryeXWWpMNsKijmgFg3iDbBR5IMPvu38uF6
YD/HcHAPJ0bGCcxZFdsA9w0AL6sopKHvgtiNgMycq7JwJHaUfUL8DHOOHEEebUyCYESKLDFfJ9L4
34fboxOuP+qIo/pHfRAWY/KubxkGUDk68wgAP92pINCczvgXNVAyCP7t/LiQo/5tw7DgikUA+e7R
9JpXknBTKY0G75D3c2k+Tn879Ec9fpE3zT9IafGDd34vE7Z6IOn/riTPEGXtqOuCXJcUg+j3rG6V
2gZ8cecDr375SRI3p/06tk29YGOCgSU4L1Qau+wTub0zcqoiLHx2pNmGZjlatyQXQMiKVEeMhefm
n47MbPjQTlnvcdgbnMT+I7QZ/uLv8LLyhpTvEAWcesWPGYCvgwyouAcbdVv3Xe+//oqaVz3IqMVZ
QYyVXyyuz6PqTNhiP4FA8LSuDzA5rppt99WwFzKJjnuxGFR0bxqkQuaKv5lM8tI1y7kj3q2vbPkA
URBZumL2CB+lOy29b3/Oe/wiwOmJowhSJDuEbVB1hRmXvzM24SJ5y4QbckljwGGD1qKnOPI7oAJQ
ctdGGIloubxd0SfpWNCEQwjrohYeY9g3UKeWLNGmoQ87ex6j0QzqPO4DWv2YWF1ZNZ/pbhNO7K95
RZ+WrX5EYdNfHMh5RXhb6oxcmTsx/0BZrytwdfCZ03eHzwI1Fd0+opK6s+Ly4gmcdKC/wLMn7xPx
F1bhQHMIhe6F90ZBaD1qXms9znmqW4dA8fdyVG9QmqibhW1Uq2mt4LKhIfaFb7UBwKV5JiXGQsoe
woix+nppugjE9joyYJEqY2fxf38YRRWYEV0O4bQtRlL9JD/OAeTYHknyVbR6MF0w/Oe27tUUH0i8
0YBblb93cXcRCFxwvX4aj3MVHuO+W6zX75HxtI0cR5UOjCWiakWlAaiXDYZC4s6P8XiHxqT0i+Qg
+9moUMO0wjud8iggS8i4+7/gJ9WSVyAWkyFq3QN1kiXAn5eN44jtni7M1Ie5B3AYfyST1CHSrXWa
beDgbXxjoRtVpZR2G86HS6aENhzJJwoQ1QrZg3kGBWsaJkVv29T5xkR//8h+qD7fXP5NSzg+Z8vN
klPrUxypkUM5ae72OqVx5ryn0Dz61wGSQz8XRpwgsVBSFHJCKT1pP2p5YYBZhdUPtgKmyHdK/fh3
DgdLSIOcRaFKumBsf9zE6+ilmIWevt3PpCe9Tfd6ABiDH8GnFuwtuZs6x/UDbsAkGRYVIBIhwnTU
bRlT9D1YS9nvqrc8WE3bG/N0NVwn0b/BlEPJiHyvH45WqBZABOz5FsBuPMZPtxKJSspDE0E9Rept
PkpTg1eKsxG5XJPd8UAJdZdau378Bi+QvV4R2Fx/nVjzOE9R/ATu4DOyFJpoFv2gLnqrnQiay83B
bxcUsF0SMhf9l5IMM9hE0FSAvdAacA8BopmGM9MrgKIgeSmB95brgISIjbuIQJeeNTcdTH0Ox7Hm
XrqUIg0+ZuE/FOZZr5WgzWuS57t4p7cbUfkII+YDz1fpvjfjWmfWCCix7m2QsUXEHxX44Y8hpV2C
8+tfRmn6XdtQoMrL/3gdgIXMTX6M3omzGBZ0G4716QKWQwUEFog6WYrss9XXwM4phaOzOosOb0Ej
ohvOZ2kRxTgF3TYpeXh/EIYSRcwgT1uZ4Ich3uhJ0jwJXougRb/aOk6l96Eizx20PGFEbDoFLmDB
Y9bb5KeulLP1yWeg599YWZfPWvQJ6kvpQ/1xRxK0oAzQXIv7ebie/wJbDDy6LsxU2h8wKn+FdC/o
f4WrgqHOv9y5dzevSZJCmTd2bOxzWMuiRW9HXgwFIi8vKZ2r3pnb1BDcarxbTqqoLOx4XNSzs77x
9klt1XFgAAXwhEDb3JHAR6ZBszPxJNL7koomKPriRvkZy+RmUKF9Dh1rKAKmTmCM9P4oB7hadVtB
PQbHpoCKQbcX1SysrPX3Clcsf10JoGadAIX6eDGvvRuFDjYqZZAXr3Y5gL2N+1qBswnRi3wXNpD+
/UWRod1Woth1UmvxnCdnVouttDTroTB5BaO2KaHt41icqFuUz/LrfDZUqAknL0eEQ6XP/o3E3FIv
LFC/FEQiBB1BTKxq+i7Yuci8G/G5OFvrHIUdMEYo7bSCLmAh3uH93sgQWj5ymhdvpFFQjkB/Txv8
i5ZhQopkBWi91pn6pcup051dosXsk+Cuvtcu8QgPw4XD3mHhgIEHXLAh9LokNMWUhKiAEKLp8LBI
gc/kE6FiGgZnUc1rld0dR8B1nTs9hpupWAw5P4/cvAqX3meFY1gK9KIFYznHzmkaKA3FmpbnDxt2
dJraum8A6W8+p80xCjDStp/frVk0pr9jvLrhaJ80FxGX6O5QlvgLNL7l8wabpONd4WwTVvLsAt5B
D0IIIBgwGDqh/W24bqtohKFhyFb6A/byaUZR2XnElp5lDdz6A/ScNUuoxEZbRn5P6Ilf/KmN1UNS
jZFlc6kO/ml6vSiOO+68oYKyez+ZztvsFKt40CwhdVvJNyhQ4tfjj4BBSw/fsJSAKZADsy30j8sx
cbWW88B97aaOB+h9KzNK85Yv/uie0H5VIj5kBBAdfHoonQb3e5soHmT1swwkELPaupzg24EMZV3q
9kyz7Io+HgmhofSuPAkZdzaLol+v+d7x2rXQAf9LyNOuDA1Ebm3HOmW15qkaKZ/pCmPt44JWXxvE
/V5D0TT6VSd9r+6KpwuYlaWC49Kg+DJEM1dd9guKp+oO5sxbl2GD72CTHOPubu3X7MjU2tq9xOTT
M+7Emmoob53iwizf3no44rlexZEf+uLvlpVgs5ZJmvh7C+B1p5OcPjSn6XGTH1I77bPMCbM8DVNH
t+S3kafq9X2AElxFbBxXZekOyNeVrPCagxq6U0kFkBW24ClthWKk+9EgT8t80Nevm3XDrLOhXI+h
0ce1nGJF2xOw2zWC+hP/SWmoSDXiBmLGOT0xJYQur+w/YdkWtC0y2/I/2xMdrHEcRFIigfn4GPok
qitp3VA3bfmHGqIYCERP1dgbYGV4fl8iLOCOwJS2tWLZN0P/N3uzva9FO6OJ0hq0HY/XIgwk2szV
KV2rCBClsEayL3Lm8Fc7N4cnF696v+xYb8fRVhCF4Q7EGaQBGMThjk5IXasxnB4R76nVn/sBItZA
bhHL9Hj66UU1z5ZR6qlFinKH8DaqFqNlSQDCysZumDY7SOWRioHrWUNMtnea7PatXiHqZfVUbT36
25z7QDfTeGbY419lOTEzmXzCm8uGX1oDavHMgl/2j6Kfs03xAxKm1CUZ764SrKNtvZlWEBz6GOxG
i0b6I/pUewCw9d6bMO5DHzA8jCnU/pH71APlrMBCLQF9hv5tK/836P+r0Udb8MPqYoyWJ19blJgE
4CP3igp1bcCOlsyTh5laCvh/6MR6lDeWrm8Sn8VrNcw662oeYMGzF633PD2mTGu3DavQTEH1ntYX
fvC9YXhdBAK+vCXvHCOTM0GpPNtHC+2k+zbUfJsHQpedvZTpMrdquY8aTQY2xLFQBaLmUIC/hzE9
1yEkGs1sdGCicT2H/VXd7JQ6+hrXHwkYPqGRv9sh9t+m+E4vne0CTjx3OPmQHchA++D1rxdzX9xs
OLS6KVc9oqeCyUzituMsgAN0+6bHHRifQgsHVRjqRsJSBWfDeSuRuxg10zyS99Na5EWdk2b9SvDH
fNSwhTWeoz5TiNQajjWgPiNpkwunogqoTD4h21WlGZiuhLoiv5euWVIo/0SQ4XQiFgRJPRaX8SaX
EhM9xeFj3GxmbG/lUsdJKWOubmFMQzuc5esdq29BlO7OJA1AEToSUUygwYWE4y7nnUDAAHSCvVGF
bgh0CChHzc9R8FPc5doo4qFF7HOzzM/4+sjsFdPI75cEN2Va8kLZ3uVvahXhAoo3uVH+NSMNhfRz
G/xeLuorGyV7S6LgaYd1CrupVkpn20AF6BLXvnmGJjUs/z692ah0+yRgdXDATgU20KhCKEQrgk8B
AkMXyIiKR1fk4qM2+UmHSxiq3QMWxc+AdhWsE0sDK2NpB9F632lj2U0ucsLAU1rErew/AFM+/2Tb
PTjhRLblg86zN1k2qtTg248RJBw+E9BHiU486M3/6UQMJrU+yH9l2lqXOJVjJUxLLX+l+tcUDf4t
nuJDJahX14nCKF2cckXtTi7j77Iy2XWzgH9HO8sx3+KTcfeTH+2zLAcfGgXSKTOhhz6b3C1RpTrT
HIa73/AD0N4vpxpnIWJAzOlDJZqAvMu57teM9kMJVNOm+Ek0jRvJMeyVoEgSZSsBslbxVS2cnyqI
Mh3m+56h0Jj7fTkyBITkJF2ukGTc9b9G0eifTAyFOmaUHn3Pfe2IOSivMpoTzkk8SuTJwBh17H4R
16ZhDrl0WdCMTs2pnhce0+3T+wJHt1/tHv3ZpY9tPmPHfkch+eWWeepzC/MOn4EK2a0kSo8KlYXl
ZhlUcV7B4UBnLPNrIhPud/XbDAz0T4JD2ucYFTs0cB9FvNFBDJawQWrfCfN2bsbI3SynM6efre6x
+2C8ETQIUqchUI2GUjBwkyk8WngdCDmYQ7WgwkByU/8XUl59f/ln65hk+PWJwEOPgbmB6tN76DqZ
86j+Q2RX9N5J0ZeSy5WaNaRtAl1ekO9h11EjOIerlqux6k7IbJdFm5o8NTCjV+SOFpF4R3AHF1Km
lSUDgCkMZKOm9g6pYFYpnDmBYjBGhxa+j0NXvuqUN2FkaJaJveqX1J/aM3HoNQlk3zCuSM32p3oX
of5PK6UO3P1LbF/EFRepthgomRO9ydUXQLj4yMa9AVNa8SZERPq8ajyxF5lYsoND+taM8MqZCnkv
j70RcaIrYLONjxdToOUIDC3Y29El7idgID7ZRni4eMNMqz+sUenPaiJ4VgkveIVKIswO6XkBlB/d
L/fw6MX5OZhw3UqMU1CATVBVAUOes2pidQNs0nw5WYMvsE+Q46BHZoJvv/OhIL/MwRphKIN0ANtr
4sqmyxSeMBMdak7pjyAtHcdVS/0n0QFIRcwP+BfCtfVmpb0xdG1ymzBU16v4IBKn/MEL+Ib7Estx
zkfiB6VnOpjqUTSGEVtnNcYFabqtQiwGiHDsrD1gFsEwvE4lbhNUlEsprWGCZjc57GOfo8kGafwt
C0wZu5au/yE4N+0jIB7nGoL5kw9ymi/YVzLZXBCd+/7JQRygzE6haqT0TeacqLKGXfaH8XGNs3O2
+QfCm8IUDU3vvCUtRURI+X9ah4EAclbyxZsx1uVTqJRGCfFgTiBwjWGnCSmWlqB/AvStUSTqce3v
u5oHSFC920K2wESYyWL+cB5sPtTwsbCCrIjxVZeuFVOq5yHb7hDQA6An4Bzz58c+OJP3fPzX3I4Y
rS+nuQZJishAbZFF8keX9ZDuRvwwx/EsAms3u8XI8cpb5wtPF0OPniL0shEFNxbCUhtw9K+Oa1Ig
RyM/xUWRloWRgns1B/SCTI+uvvvPex2xBF9UmzjjdCC8Wc+9AXPz7mx9hf0s6aql9ld+2ys24ZmK
1mvEFINDGmoosWPd+xFNMWQPify/fTfFQQP+l4s8jCQKpeunmA6V7YNenkjg4uzNSerQ93smNnR+
RINa0RK4Mkimjj5y/2BDZYuwzbgx7cYqRXaUKYeNzlYoOc/d30tcVPXcdNaGl2E4Joj3pUZvluLY
/GmP6OeyF0orP2seNRAKxWId9HAlIMBdk9lfV0A9L2MMnOqVR0H1LrXIg2pCgjwiI5sFQjTqVJ17
rVOpMyPiHlXhPN+CDVm5fzDJ22tiCyRLJAn9OkJ/Mg7rkuiECPbGPPuxT6lOIypq6h6UvXfOehif
ETb5SSUUSSTBvSunD/n6YjG3tp+R92KTaF3iFZ3RSwsj8B6KLxgHJfr02VRI46QiTCv5jylfMPMr
UzK0ZgpwpPzkrMg/prIo10Rb/TfPxSIGqzUh1rXvdmRNMdeLvtk1JrGF4X7kM9ojz5WOCw6APpA1
zSQwEcFmW4dd6LcZdn8NMFV29DxyWUxnZENcJwJPeqRzqndwgd5tYjfyEB4eN4RDwTujqZub3pYZ
pitzM6LeswMXmsl6jBUinB27mIxEQyOucTDy8I6FPDPK6wQlMrQFcNQUchs7hK0rurWdBSeGqioe
auwvL/DE9/nOQ5MNsfBPb6KXpGOQVdfXtiRa1yp7ioyuexc3YMTwFL+7giiEcvcRNYtrCxRzm+1v
UmDxLoggkPGgwApfRXrd7xivN8BFmZoPIQCfTufVwgTdWz7fLjy96hDI8J8zJPPAlKHTV6XmKtTX
hY2NJbc8hRn/wEdEUMKT0308ocPiDt1ZqScYuze5tpG2jd4PEY9AoBJWhM5IoCbCrCOUC3ZRvbLS
QGXt2JhPi5OrPpJXvlbkiuehvuAQcG/Qmu5wVgT6BDL0CHpXbUiVMkR/soKdVSw4LQWawX4bLh1Q
VkSEcEfEYzhEZR+QAQBFtke0DvQpP90Y7Q/oC01rQkx/JYMvKHa9nFGKGyQEPJzfOsdoV4OZuG6r
akuH9xPQQi1G7VHPa5usFfjkCw7Q+JT96YHiaK53RJVzQRxDOyzNa4Q2xdtO3nhHOLSqKlnT/4gw
PoxEfxQZAQ9I9QiqUrT72Kfjy9P2tml7P/3bUxrZ0XZ3U8riT9T6HEPtJFq8tCzEPFvpEjUBOSAs
bl4eVMpk8/SYJfIb+W+5xIFtjbPGkAM93+rwukgmEWquUenyQE0jg6JLuRirWCx35cIe4+i/hZbs
m7EEGSudUVnkXxiv34RceYmvq/UtavuztIwq84L9oPlG5nN9r6nlhg9MzXyRi1s4/SiUA8XkffWS
osru0h3LK7u9NV4bj3mEcKcuXiB/gnRNf3zkEnxVG9HwD0YcrzNF5kB3hJtUhnHdq0muHC7HxLKA
itRP5UutsG9OFMzcsIGCybmf9wHvs7iRpu7ArejXMpoV/xKJXOMeZWP70BEv+8/3GzB7I1LHT3tB
dryO/P17LSN3Got8DNQ9r3N5ZNOdeBnzBdL+U18lZtfJFIrV6/8j+dpOpV66Ex8nn/In6bwi1ski
lAiJsk0mu3WeiHsbj7rGJ/+WyCws6yzjHHfpzotvKKNucaX4xAFeJUWrCUoQru0ZVQYyz2Ysv4gN
M4WJ7KG3vZKAw7lU/Eszzs/LHLxNVrMadJuLgJfJ+oHYlYBI/9VK3dhamQG8UCA5t4r9lElKrvAW
Y27xdeFh5+rvUMIp4e3raI5O4sn9B/dba5BQq4q9WPxBDb89ZNBy8dZKlbzF499TvS3+6kwKhzn0
oPlif3J2jzQgyjxhcQ2Ox1Y24+db8GR8v3d6BXePQLbD2NZg7dxSWCpf+rEaJAE6mBFZILeA0h3w
yBxzg5iqd9B2vae4EwFaHVWor2MZ/HBrHY5Mofd/qJXu/+bnVy1t6bA8TfhM2X6iH319dHkvjBvn
teLrJ88caqBfkCqZkXaeuPXS1MCc2gn1PzKInjD5WDyn3JC7m1nRkl7baw1kiyJ5T34hV2Lj3bjp
RXvG1qgqkfCoxCVSMPSXeoAekDR0zxkMjyeeCw61hdvq6VsrMabP0OcmTU9ROhGREs6pAFZi784f
A5zm15DDSi0Rn3lwdYkf9nZic/cPwlJPSISCkinXV0yC2R1Ob9eWeW+mee+xh4zntPmMhMzFfNvf
dQW4gLvPxUO+BOFopDbBiehIr62TIVNz7LhsJFK69IOIT8jtrIxLPwmmuzWuf2FYBZj4R654jC/Q
F8R8hXZRad0D0APuYgiAd38ayTY/faPVi1ryFxsExz1mhRraJgGk1JwI7G0n+5nHsNVx9TXpRMZ/
rhNj72/GZ4tFlUwGVs4kb6bhmtsa7LrJWWYmMii0YnPwi/9vZZairo/TRFiEwKpt+OEnC450QRdZ
jh0EdQKlFvM5ryU6Hb6ZfEOKmYS+1HYQqEaD5HWjear0QSUI4udttMoqTn+rwb4AkqoBucEW+8L0
Ov7f7trPFW3CjoQM9rFsoKfr1VQT90b6Gj+iu+6NTxpwsBLN6vv90MnpigSfAo8vudQKBW7C/yTt
4NNXyqsR44ShoSOeauua6PmnhY0F6Mde5ujbEJR2pgayQqZmqZmiyjfRRKSXFjppK+Gkr+hmyL4X
PkJFaKac2fpW2f64E8vrHdsMZT5SJYABZPUJIQpZ9r0TXJom2G/Xp9Krg1WQcAZq7uNSCJSXo1eH
rohuxUC6eDDYn9l/QW4bsj4T2h8qya2LM+9MWfpDva0HV9EzsS9xxK0DIaSmyYHCNp1TPQx8JWdI
z9a8f4RrLtEgLvtIBWiXzlunCc5PUtU6BC71DrRDOuOFtNyzciZUGresqoZpuqcQXX/PBLU0sEhR
C/Ttc2ejkq6GnxY0pJSZlzFqguyFek01sUx1nHEy9SYseoHf4m9HjCPk3+oA0WUc3MKISy6A5rt3
FwrhmtQ9Ynu/SdaVihgBvGSqEeHz/mmojF0UYmJqNNnRtkVTm2OtGdeaOSN1rOmFfKnGjrkgwDE8
lNR/NJIGUl86XD2kamolYlYidrEgFt0H1bogq/k9JjclLazFn2DqkYcWXfVfXgznOxaNbDoEU2C0
m+FLgASC0dlrkJ7SKIHmqFwpHKNdlU3q8+Ijgm5OEavtZ8gHyc7mlwfnxjBSIyL1ddax9Q1f9dUJ
1O98Yis14AUxoxIb3uOETaVQZC1JCo8hUDE1Saxt0Zr4y3nKJ1xk/vEM9Nb9qRV5GlReBFes9abl
/STDPc2ggbNHVgfVFNQ0zETmgu0EbGpSyiQ0EFRuoDNRMPHGAmg9kuGUPUblsg6FZnVu98XDQPro
pDzK9F4ULXZf/ZlA1fgqs+4mZY4vizqhBkrU25++SILJD4Io7WS/skXJMq2lboMZTrpYUdaC/oUR
gWolSFSxpdDEOOm7pRaec3DE1JSVmf9CgiN/G3rA+8i+sfDWZKgMPVVFUsrPlcFLvaKvvNj+yzpd
RLOwAoZUklob7C5WG1Pseu672TSVipSAeVNnMePMzqebGI5wNYFBL5ThmEXqTbSTbCvK2iYoWhcp
W5po25mWke0iHchTPwPTMyttrkpId5+Jw/CfAKqi9S4vaqX+j3Y9NI0zIQIh0q3lNv8fJFeVxwdi
v9WSDqeos0w2+yPCtRz/i/0EG1qCbcER+1LcTo+8bYSV2dQs6xrF5xWB30JYwDNa9bHeXprTZTh7
lRWTkSyC3floDQidFDyIWK0jG1OkmgiUDVPwVn5vnSh4DJU8aAFHFk4zpbgBjv1kiBDrLprUb4fU
EY7FHea9UH9/IZIaKcRty4JWC1PJOpw+0rM4t5n3r+EMEIX6mEX/0e5AFhdfIuAAdFzSUa7AWIy7
7OhTckurDwJ9QZJDc+46Ngcla3WGf/fgPf+XFlKz1v1VLOe1FgoH9Qwdiv4o2kRCoTinNp+I8kO6
Png/43nVd3ivQwYeUSKXZ7tWX7e0Apnr1C4XLCRf3OvYdKoPDXjpksmEk0nLz2caNYuoQ6yG/lDP
t0+usCtmq1SKs1aMA60l29fb2gNL3+ET7EgFoYLmJYxsMlmIIOMH7Xpry6Dbgv4ZFDPQkaCBHJs/
LQf+tO8IpA+xVr499PlzeeBIP4dpCOURRj5gAh7+Puf5IPQGagcdKIkAn2gXDJMN0WOR0B5DrXfh
GONlwYNaqcDJ5eXerywLvdao3Zs4ugPzjlxJUzVvFVPKPc0Ls3QHWVXHYqB2WNgB90sO55ISZobp
BWmyb4+V0z5nDgvWhZrk0KaBYzp5b5wpw2lfMjFOsw0wZPYfP2G2rzsfcuFLu/lk2dKpAUwTPmCx
Hpla+vbigQ9hGmOOHDRL/ldzw4iWNwErUZLwyAIC99qjIkIbWTxvH+yOYUAx15zK5yI0fRfcKvME
wX1apQ2auu2icxXOe94LGVhTkOHtfoXX3eqicS+ceozSBps2/+J6Uw2diF/bMJIaXwGLMqxFv8gy
FemJ4z/Lryjp20e9nd2GSDGFg/lR5hI6+WPeFMjfxtXGg5pkOvGkHqwXAXxdf9WYQAzYwDmr0bU9
JxAcaQZYm/lW73kK83wW/A6HpeK8IOdgORqOwqX7P1hvwVhNpHCTL4g2GbVbeaXkodl9vYKx5hbs
zvOinqf040KPgN8CntsYRPO0Z9iIPXi5PPqbLLxbjeDvq3xsD91vX7dEi3OeWpTPKaX3cqZ3qNwt
XVeFZ0EZsRFGC60oT6LFAEaWiOp/gXTjN4GA14Ll4GjNOM9Oe7PG0le39IZ922cSImeoBdnTRqyh
nOjvgy/WvduigS019tZMEvy0YwlxzKpgDEol4bbQk+vx6BcnWNXBqGf5NXrZ6uigB3106lg6q+n8
uuk2ILL9qrZAifW31MpZj2bGHsTOggddNyV7IePNCT2+ZogGlM8pMIWCphSLXlQpMgYmRdvILOfO
rsnisY18DAEPIlXW4bJUDOlqw0nez7qSCR3TWn8z+nDZL32yyPYMtXTDGdG5mXWKMEHufTTq9aMW
gYkHYqrI9hueOUCrTka4xW+5qZOjlEU6mKmqs853RqjG4tdCk4kR+f62KKi0KDVYd3olfOBgSKTs
oxDI5OpFgqvU3hG0SDIjkYnxlyqq+pdhX4vvXtkE2Ggq4WAtY7hGNaFIwXrv/DkFUedXOhoVCIOZ
ZCmEVj9Q9LC0tRJz2vtQnPhftE/RDm5sWhrMVHiIqnIP/VAprGJeSfTLopF4pgrgGzttux1UJ62G
xFxGExmHPDkAD/EC/+psL/p+R6VzLEU3nCZ4McP2gZpHMMlvaK8u7vfzHuhqLO9sYEKwnKk6aTQS
jAM4BdRJMmV8cQyAa41gHmjj0zq8WYLB88XlfkjW+BacbsITGCyv+CGogTgcu41C2MauHeU/KJv7
wFiwh0nG2E/0eQfQ7O8Lqk5peJWe1tjLjkeOhEUTtw0bsoR2ApsLvzQY8RVgVj4LyYayL8hyHzle
LS8OLE4O7LGlZvtYuc5h8sK2QOcO9Bgu0mq03/RHrwyVkoGKwJx3S65vXFgMGPbGdaKh0XtATlYC
5+dbmgvvf8QDW+MwLX3bzI7nBNHB0VC4ZHIorWS2QekuBFNsdD9zIw0zHSBuUumV4SbuOuqzmZGn
RvImbGexlR1kSSy8gJKV15JWtZgNl4Yk3tpqkemP2TEwx2FcswnMaFjAczev4Sr8Lr6pinT9pJsB
uvarjyY3wQbndGP1jkChVntp7oZERd8pGu6G9XkQWJCXd2ZKNiUsbPVmCFzou/x7spJdrOPTGX8P
peQRmFLrkxhpR8AgBt79LWHV5g23s6paKtnqmPLlCLAgIExtlkBYtU+ovHGyX0+rIJJ07uyloKS9
ad1FHCbyiUdNbfsLzASnt4FbKYtnKVHZEvO8pwxkURSyun1/S6hxlUvYfgj09D405m9NWkaKYhW7
ePjmlwYzVBIteovvcuCfq1kJX2n3LFo0slInv3fxGOk7vM3yGaMbQW3XbMkd7nSqfCUBn5gD12b+
Py5ztCAZQSL5BFwKqN1MuEScsh+qvj7EMYk+UibiUJ9ljH+ojH/dZPV87T3MUnZ0i05hl0uR6MpM
LudWAqTThPXnAtOrFNxL9zMvgEs8JLw0g006id9nb+VD70xcRBMoDpJzktFN7lBxhCNgZxAPcPln
/gvU3UwptrZ8WW78v1eJiZavecCfq69yDyov81rO8PA/zxFbO34H5BtN1b884par2iT/Hyot1jWj
jgVl23YUOoTeazBhw49R7ibFzEWwksCb2PynqxsU/Y7ZHJnNeLIvh677sFBU9iDnWz3SVBPCiDS3
etsPauvWiJt6BE/+fAajlBgsYdb/A/hzgeWl3mORQ2mvOQfr9m1BOxx9THXq6CX3FzzFLG3UqJkX
UJpG6TmgLbPrQuCb5uUNWWEBiklP5nyop64Qr+fH5Tlnoi+0WNJapyEaFF4Qw1L+tT43+qUB/yUh
ZtdcCAA+Kil4HJ8V7CSpS92FX6p0ozisLO+yeKpA5abbWXsLcB9DcYeGTQ//Om/hi/6XYus5AiFE
35hMB70hP/JKt7l21AktGeGWLoo5BGAkkAWxmf3nO/wHnGyqVR9FXCePAq5i2hYj3uCa6ranQd8i
nYpgXkCpktpTYzXkOPBo0merawT3qPGyr7mFD+RvFVLm9Fllm8xFfdRtoVwnQtxt56KEvVqERdcj
y0o7MmvOQ7ZrgsFsY6DWG85tNThCE0+cE3sCpsSHKrErGX7S1jZz5XDEhIS9x6/6jNL3nBDtf/AO
aagp+XSbo7xFFPlz+7IdLkzU4JUFt2k8zAwURT4zOySG8aaohkDH1U13aDHeXxmvMxGnhXKiay1L
GB7VSgs+L9pe61EVztd4bW93MKcoCCYyQhjmy3TyqDFOUsYfYRGpxe/ARWSwmAUumrDRqATf2gN9
IUTaE2yP7eoJahBWf1ZYJlUglawjst2cpx9nSelDrNOrTSqzJLtHpFwI4M2VvPklusvjybaaGpqQ
eMiSi/MpS6iCEHqVIGoJUojN/GTzTeGPXFusLfInrRYzTxg4L5OilklmoOvIeUdXBRhOX9iS35rm
eJx8uFb7CHR4I3LFlKC6YjAlFJUaGzlyrcgsefOeXD5L0YwI3YwaPuUVMUjxAMgPPuEwsFUZ8x9j
lVPjH3/5zbOyaSHhWbCJJMaU45Ox2LPEG1XgkFGSATGfHfHiH0N7WVmBnQZiiGSM2cjZmcZOU5l4
c4NtZyjgVVGbiRFwoOq+OVZE8i5a0+TUMyCLeZZnoynDubkRgSvwGvzvLNS4neKReeNQCnD9szmv
dePgGHWa6P1GTcBGrestdrYHdmDCDVyqwMtZU8dS6c3s6HEK4Yldx+c9oRoMgri+vETXGXpbRpqL
vbWCQEm61mlmWWZzmp69PCaAMPHY/9oz9JWxGAMWQ4V27ZsOiAks8vHqXqrOssVTjjkeyxs6XpDl
8mqVeA8FIGEmUcRUwTiAlmnsjKhGqOpOGwPQyxtNlFJPUUNmHX4wll1jkQKKostqrtfh99IP9qsN
Ax388D40falH+kF26jjgYFZXqiNfDrr44u2tWy+BaC3PD4tQGKxvbww/c1pRzV+35jeWD6d8OgS/
d3mfzxtZCkWMfNSvJrrwMCDyvGV2iTiwGBm5waUUcvOdK1OQOqQy2+LVthDjzNnRSbar0+Ey8yr2
wsMcKx0hti6Ui7nnWw6BqVLZ5F1PYAf4OlZIH3kta0tnDzAVrtENQ8ryKnHxZO+lPlxyWAmj9JlD
XoI85U9hGs2CGP7mBDA/GMQ/qkblKYzOWFXZOVCjPoVte0CYUhZFIYp38OsxJsZkyZPFvJMU6qXg
iyC6lx0scyTdQoT/vLl/S8KnHiiIdphrWII267WuKksDKDoCK0VZawk9n7RyZRfZjhnq3uvu2nTD
BGqMts9CoR+7QHwMQqqMgs3hNHpjGvSiFj3/oiPOOjXCgPRRU2kK1hE3eZYlcBKwHxgT/zfSqIcG
jmDyOoiV/yFPkhP0rRib67T5LnVAKYGClneDb++tHqM3zA3wkpbHvMzCB/oOgn50CSEMYk3TicP7
JeRE/i5uB5G5WTFI/kgigjfAUSyp7WoEGjgyO9oAgYUsgYY0KgPOe4aqPYGTx8s8vi8XfRFIzDHL
MMBn6JYhEoiOZtBcXsLyKKJcgSfsOrR0N8b/wic/J6oziTHeLl/492YHul9+7rvcrdO8FdVqezmK
6n01C2LndUuO11h4n3VVTR4aV4wV+g9SMvpAhnmYx9NIfuLdj01AlSZox8UWJs1Rvjj9oMSO9T2D
7IWnI+hOXjRqOuHToVQ3oZDQ2kpiDzUMqk1DwAqP62VqZx8usWZN1FWupR7OaHJk5s5lN/+GtX6N
8D3PnzfmiqyZOjKHK+ycjYx0AWWdb8EneED7NOgSa0URVJv2Eq6QonZSIFvsxbE1W8pQ39GDp49p
mo9U07AviTXQ9whsld42oqoCDk8cSPRD0q+js6fyd3M/QjKgwNUyt1LEbxgSupiwjoOxTsKVENzs
AKlfCRQN/y7/r4/f69MbTQ1+ylDI8bYQf3yOTT0iT2+VOKHazIqrqSwEeWqlu/oNmgZHBeprkYrG
IOhRV7xM+glNrZYXOiBpEb+O1PyCYg6WAklGFABv7f4T85kDB8ieU8pREqM7Y2MypwXqF+qMrih6
zDupUyLJA6euDBz/25gaC9UgCxqmXx4IdJVBSmR4VU0dqVLK7GdmYXU05rlE/i6br9LMvWLShRjE
x5kYzNKFp/Q7hhP0d8T9Ipy8atCBpiDRGjBA+KVaKGEYqhcYj7JOpknpGNM7Jd7GG5l7d5x1h9n9
eAPOAdvIy0EuJpqMD9yB1k+i7tcMyAgyb3dAHaHdQ4zn+kaJ7Z10fkw+I5cZtPxR1MjKY7F66mRc
ZhqivsHI0NG3BCbqU6Xa2L9wyxpmSDkf2HpTWW07nowawW6I0h28VmgGES+oBeSMUKiRWUIlShGc
YBsZnY5SFY8kEga+hI6UyksKccmC7nWSPeRgn9uGBdDOK8tB/dtf15uvg8UjQYZmKRu3qH0LqwHM
7CGKIQz2RAoJAq63pGaG/z0OTU/wW7eX5VlsKcSyeaFUsfhq/pn9pmvJwO3SeUNM8OFQ/QqmfF2E
QrqXYwSc10ymZqqK9/5Kbh0vtLwozSm5HvjXDQtJPvxrO25gF/vOG/4a0lQhznHVnv5hILAK4CXi
MU3MEt4ddxGYdVfHqEXHdvkBCSPORUuDjCiUsWzHxe54Zy8+e/hu8OZGUO+bld/4e1b5allj0LQi
zZVi/AuNmhIZkxw4KpLNaNsVuJGl8fJ1c+TH1h/tDC0Ky/h81b21Mdar4dG79bVxN+xDWTYp53S/
boGK6Bj8nioW+Vgtja3XqzTGeBMo3rK3+DQvcLUBQR5D8kkdzV58biHFOBBsYV88OTsu1ecSmf2N
tCrL1YGZ/OYr9W4kqgzg/P7E3Qu8mfsMrdn+Q0H4pahs4CI+QAkL5I+o56aXLkeVbG5Z4FjbHmf5
zb6WjH4QMbS2xB9uaX6CRY92FtPF3nq10Ra8MY9fd+3P31yvUuVIKG61N8rFbiuZVgUiTfeJ045n
Au6taQPnaFk1zqWlLTNZ7cOALTE4LO2ChgKwQKhX8/KPzY254LQQqlZAwTab00KgbtzhHhbiNgMI
UX0Jn6DgQhVDu1UKppIF33tRwJjol2kD7iteqlx2zEvCKKVODRDM1eQpPdBFhktgTRRDqxf+5PK1
z6g/BaADx98m4xHrxaTH5r+M0fOYLYEMjhiLPgerapUtA9AojwocYBHlXd90RG0MTznvJyDL1FRF
WUjItbuATbaJD7K3FXUhgkVlBK2tyRQK9sxyyGi1yY/Q0cQj4qJqwsxq9ev/64X9gy+WGaeLI3hi
PeAmXOCgT2SYbUtDn1cBbkQ5q8YWaC5mpmi6249slwHDCVBkLUQdSXY7OgBJaawFLommB61M9VQZ
dWT4GdRp1IkL9xfssTV9xulTiRwxwATPg2AFjJRp/2Si6exaT5Pepj7QNAYrqK9NpePKkWz3zLbI
1SI1oknhVPQoAUOXNFKOqd2iS1nHBLy0Las7P4WRG6GOxNOCeAuKizW2yqgirnS7STRkqQ4FrS+r
otxMs802tCgG6EQx3iXRGPorjbK8SqqF4t+KQPQPsqSiF7qMQw8LpNzCWHSSfocnYaznzFtuVNFx
zmqK92xiwRZI6fHtj9tN6cqO+6tG6xzDE/BHRkCHO1ZLy25aKXJ/M7yXz+yAnRfgAInipqD/olTd
884QxAbZuD96jS5nTP582kggqys6X+rSVdOg1b1ptS8W4TZNscZcY8Ys+BstFmmoi5pfFiJxGtnC
TMfa3mSLPu81JVuhOFmBMWyagMiUc09yJo6aLYz12O1J5V6Z6SrCajEi/2pEPYdVtjiODx7DbCAs
ZqBGUYV3CTKHGV0iKwheqO3kORy2FaTgbg8KBbFgUsMQl/5CWPHA+pg8Z+ni1fO5xlowFb6KbDC/
Rk5Ps9Nt9um8Wk4mWj/N/+jigebxMRzR/qVqg3PDgszsNpJzO8o17cFDQ3LbjajQLEXoCo/PV4el
pbnMR4TcOYus1IFlebGaz3hsqeXesGJy4JUfjVQbUNBAqw5zfFoVVGVaqm7ub/qXfzHSSi7WLZP5
PxxxkIBQK0J8v4DRlpRhsg8vtsjUlp1YpHKVDRKW38kxGx7RJxXGmzzvSZoIhEMa/Ht4wJbFC+FP
dYibE4EHnKqtiZ9PcGvY9x6SuDO/9DZFOXKbZ1vBLufQDTKtyH+tFa4iepXtHytPC7NVn0ObgsOg
pmXjcsJi8g4rhdZkfL4E02orClveTyD2RQiR4ucbitKJuhBIpUrhSuPgsFsIz3CzxEPxkvXRka0c
CiGMa+XfLfxyVXcvTfQTv9WeZzizJZaQJm9CX0r2WdEcfCREsAAvQwniMrzuTxpiXFnvmZYNrqbj
dz4Vf1H+x7z1+rvA+z7x7lnLdzWgjmeQdC6LhbIrR5g2Pntu/B4V9pQt+y68wGOjBMJe1chw65Ik
RYlcfrSt/hrthGx1NL6tlz7hQRthtGwg8KEpLKPi7UwD23XfkscC1lYrzah0pmkuSxJzcfl3e2lp
LVBFPd1lc3/M4cJ4lIy9FzMBKZW3YGSZb11a+oJH/+AYNJw0Gd49/9hq3F5+nhINm8TkS4Qg177c
yJhrfNlWjCxc3R6GqpYrvw9Kwfzm6xNqPPmlUI006P8RnDdLRo37XAptcpXk002Woea4SDo1Aj4j
uV26fw1t34Qi56u9qJ9ucAxYRGcNYC/gg8rzaYdleW1C43xU4HHRyH8ej3tqTYB+yUj449tNLPsa
2I60c9mgXhhpHkl8t7OdwZ/YqyEeuAxRsbeNQnkMQ9Vezo2fc14/KvKGkLhwJSHQv0wIIm5n8/3t
7QRLThz1HcjmJOmt8W4hQS7vG6KGNtxawxKc1HvJ36F1vP00947RUTgrcACnj+wkv9W4D7Rer+z5
PcK8eXs4eOv1BPMIIStf6E27b9pBSEvoByVku1IhNKrHgWRFHHkeXxCG9J2gBm3t9VH4EnuEsY9V
QuhKkMba3cHEteP6hTkhHJFkZnmBSCIVzDW4UiKCr5MTuHDNjbAcST5gpLaEampQql0+vkMDUufP
7iog/jKLnKGDgDxWDbuyTgNep0UmDxpuYMCj+Cl8mI9Ax/uppAWBecGWh26YOCIGXJd4v0JJ3rkK
5jC3D0Nyn7c0Lb+sTg3Dq5ZdfH9FuEmGJg1A+VCdsn04CgelpVxUwAvjlNc6iBipkOxBszHWRWOq
3cWKNNcSWRPTEPeoHu/XrEqkDmp7jSUk13lokQtjghzx0ubFOWetCZ2RIzbUEOFqp2/Gj1x59HEM
jNSR5W4psEhTMOVzbZVwXCa5dDzf44yP8AKAMBbTh3ymDAPSvwfEWHGfquI3LEJsWoNkb2M9LRri
jqKIrS50pOT1WolzX5fbYjHAfVfoWS+U3n34yWyl/WgKJwk3vTByZk2UMR/Rymgo9Z9O621R9BLf
jM8OP/sTmuy+I1/bi7FOszxuJO48cz6Gu1+Bn/eRntYmfDHcB6I4dF4g6Iqmp07gPIQRK5E98JaR
OITdqCKhI7fZ/b97XPQd2biZ2lBNu94Bz3G0ACi6VR1wvX8GsLgSdgZTup7tpfHfrf8qzhLXQDDY
U1SolY7nTQbi4pAsCsfmaYY0g02jmlxWCFb0dlCMbsf1PK+XV6X7SOWZUgBlkA1ePHz7SGdyZggY
qobeEfZPkuie3fiD9NuIHwlaEWR18JPTq62bs00UlmTfb86ML13jUnw64QytAunCnRXW1Ozxr6FZ
HNqdldqroz/zCZygW92FZMmCBGsPU2wylpxi8vwSs1AjhGGPxcPF0cnAU3ja1PQgDKlDlgjVf5Yr
VmY+zzXJx7Ppnuy5ygW9rpRatfvEMk6Diusuc5ijPwfdSC1+TNnDDkYS3eSCo29Rh9BvU3k+uvuJ
bOTk+MSCHAbcW3idLFCAeL4G8DGJhfICRbfBtxztyMlPjcTkn83D8fv7BY2550hefF+vsCmJs23l
RzS7siLAc9H8MlpJg8tq9QF/P0Xc6Bma03WWowx0d26WrLb7ydmFBSPXlhK3QSLLvcLS9aziZ2a8
EqtVGx5CjKpTLefYilLw161Et6B98r2YjFk+rL2pz6v884KlHxHBEbu8aH2AwhFT6EsE6uzOjohv
/jOt4owhJlwxGjYyMvm1WNZYcgbdQSmE6RxKcPtMh2WFadiuY9n+3L7JvZx7fnfbHVklT1nf9Cei
Htg7LsqyAuTQaQo7uWZ9a5P74c5WDvQAT1MR/Z5CZi3FlI9qeBId2vvHT5VEUDHJWo124JC1tmqf
W0PgB5tILSkWKSzwOZSWSvOBlPivaP6Jy/+I0I5vDktAlFVV0zLfzrbTfh8kygog2tA92pQUgdG5
jUZjZSfUBl3kI40wJcTEi5WYYN52ZlzDUiupExf7kiGBMUJRQ2ttygWnXDFrXwdVrcJtyMFQR/Jr
52FZjVb3E3JQwXS2o64xvAEnGGptS8xhGjmJo/H82Rv9z2EVx6I/61LU+oDeMl5+eCVuzXpNGIB8
CcFpMfDrxwp8d5GmmYv8zmaOdTvonVfbTjlDS1S+grgKseZgzQzl4o/2m8AkvhlS+eiJkr9Djt7u
9UtWyky1xjc05V8YdL3bjeODobu5FIU0ZkVp9Vpzp+MyqfIvGJPjlVKZJtyVTJs84J5p1DCPWNVQ
DRaxCwxscW7RCmdddu1sQiKShSACjPyTTDYmGfjwvRP1ix20ENjYiK8Z/3diGRyjYC6Nyc7dbbtS
A+pwCzHXc9f2ZZfz+qwmasSnJykyk1Mo5eRe834i7AOxx6W6v+xzfLDOFN6g17XlJ1icNX5dY4P4
faWtJ467aqNhKZfk+taN/Up4WxTxvnwQQCTWOSKWiRtSdQ74RyN4rqOqCbmrh+qvcwypV3mI1byk
RRGz2N6Y8WCo18aZfueWkl3o2e2/rDHbu+7+UPjmDGamL/sUvlVrOvvhhPiv27laT1y1EYd17ydL
omQuKeNJzeLg0GN++11z6xL6FTJSyWcPj9RO/TZQ/fjxTJ+ttyDJixs1whwwDLJNba5zqr5Hi/4e
/B0wwb5S2eg2J/6bA5yDiosYV8TBOYCxvZ47PdcpQj5tzFRUKKj7VoSjfXASEKZPq4dBQweeXDBW
cuZMSsTKfC7ppgcIXT1/aNdWZg6av/mLu07Td22f5IAMqGpK8I8TmDM7BocappGZOdSr4F9to7xv
YdpRgXKWBCjo1zCJGhodVJadSB/9sgkOy4gcNb2Fn+kHuRN+REwh320h6dRvyye0A2eePTj8gnTL
TLy6ySPm17NK2Q7yBS9ycKRrjVmzsibr+reN7dGaBQIc3oujDQgEKwh8vSxGGcP25NgNEOQ2D5W2
5mFNKq3HtgaJW4p5kcHZjlwuk/bGA8fL9PngvWvy97o4JEMJzu2be0kwCRVsbSDHGjhHwthr6w/p
9rDf44zaqqr0sgyYF5UDL7iMT9gmGe2x7MW4Qo19NLhvaegiP7OuHhWpnwjF5tOx5zn6Cj/95sCg
BG4VbHRUPElBqByUCu+BbqnycQY6dx6OIRxa69PxWzbJgx6emSCYGK2i9dwHMwBaPrVdyfDGHHex
uuDlcyYjmFH7nZmm095BgcdAsUNErxlNKIBX9EBA2NqVst/t7i9sxEqPZQquDjT8x/hF5kH4PCoH
glQVnj7NuM4T22z/pKhFX6vIC8EL2Xlsjvbagc6c7cqzEiyMMrT8QtsHzY6xoMoSaZ1hFc+bE2Y0
0EJmMlTyC8TWVmWaNaCzhip/5J7JbWnA8n0cwa7/TiuQhscLuq8Hq/kWCuvAn3SPdbHtsX7d2o8r
Vdub7ZDwqSriTkMIMLkdCKvlHsvN/9q6Laj7GzS4Dhif+1TsSGFXlbaeTx7yP/T1lPul3H9pQ/N9
klWxDkEW5mB4hjn9o1M5V3oPLgsEqN41C3mI2LCq9oLRSMg9xkEVqGjjCguhRbaiavAJfpQHYE+w
CODszjyHruzKNmhIbiW+qt/dmk/+Xl6L4SM5uNd8e5eExs7g5fvxD3TdwUaR45Pl/rBJGAcm/T3k
8OyU9aOzFkvlD3OYY7XnoY//T9VNl6WBaHC70/KPOYhi43ojZ90H/HXtBZF/bgA727cZbPwIBOHH
UJJ7KpmNoNtZh/PiexCF/fhtULqzZoZkBs0Wfhw23t8TXVXFhXdW+fI3CUL022z/IzxOH7O8AklY
6xvraAjxgoBBIZE/+cnLAjdsMXnhG3KCIqIsCYyo9I/tr18RkE1ST8CD4Zdh4wS8pzDhIhL+h9cT
QEUFvT4LpLdHefnPk/eTLUxwmDJ43VelZo7Ad16Sxh3GKyM3SQXMigGIPuFoD+3eD0ocW6zD3nkg
u91oPs/GbgBOkKmMSoDrQBh2+p3iClo9Lx/kIAr3Im7V81GTCNnYQXM5JYwvqtVvusvbluoD/voQ
EoIHkseDdvD57GnxwX48Xo4w1rdAYXeTGJUm44o72n/ocLSxJjoIVI+vX4+8Kq8bmw8G4X1AjLic
fRHU7QNOEvJf3wi/jlMqHWeMBFivf8CDhdZ4/DCATPAWeMqzVuw2Z4uAy8PpQJl7BbGENAtPsmjW
oSNsDIcAFwYD/xpJJlb4soxl8QzV5F4dDMS6UgdBYDNIiGfeQ8HHH9rQaH9Hmlt49VQerdsd41ho
7u1InsKh96kU3GM8/cGTaD5CiLUPEsxrs/BUwcDc0Ju5MwQYoMtN0F0lw15Y6Wbr0RE4v93VVxvv
UtzVjJdhc1E8cEKwbVVxWwXDaSv9odT9d1mjhZfeHMSKi+2OLALT8lOA5QFBKSf3YJNzw0tZj06r
Y4v5bGwyE8i52oT/PPMH5TDRNdZAwwchjTCq8z7aGuRIFeFhkN7oR/TLjt7jEAGMTOR9iYMv9M74
v6BrodwBx9sd8hM1zr3GXYPQJd8+zLIn4htHIcIY4QtCl84/TV1SgDDwX8Rme1w8awTOLrkgECpL
33RABJSiiO2iNGZu7Oi3D28p3/2jj6/kh+fgkbt/hK8+Rl6DFQCAFWa/88/8OmqYd04xXICYzP44
IvXQCD0fbExvGrpVnAVMteojn17gtEKLMIFztsL6RkSJJrzE3HAIz9OjeaVJJz2ElgDD/jrxTf2J
8tk52wtYJ0M9gLXXFB5EIVgOcOPcjb4lXbWfZ8bPeef5t+ush5gxaXMmsnzUWrhHzZYPykqA3DaX
0MzxtK0Q3OGBHyRGuZNj8YAL8z0Jy4Mli+97bTYQbhmeYfSG/QSsdly8QuyXBmiQ46fIxZkMh0pJ
Le6aLCHlD6mwdiQr/qEmIIWMDGq2y51rnPsRozKzeHHaDdwbDHmNYXY5FSrM7UlD+1cAGZV4e+pb
oRYFe0VDOujjGVUywXt0UFoWGvjtt2vFx80wC6eSeoHPXWfEGMM3RTVhtot0NVWMnnrUOAV4WBf+
aV2lSRYmKhOwR0kiX0VRqpCKoqmw0RRRjKaR9BsPifzXARam2ee6eW8aDu5VcNK55iw/nvU2Uicn
EJbN/SKPV09pNDlck6vmSiS5OSw2L1C+/hzoGer73nIhKqAvNDhcCw3xp4KP5PYdWQdosmiZpDNc
ZJ8pKTsZL7n7L1v/hHBXpmLIvxJ/u/5LlV+6PM+kaRjwuAXNS3DipHJ+0wZPvcfp6fu0FEfee/dR
fJYm9a5IBqVUm4zyt6pfXpgHrsCCweMGBthm3XyA58ic23M8F1GqEVPvnKC/TAsGFivfyvFoaXSs
8r7bA+y0mOjcV+uLNQPqEHR1T8ucLiRTqn2QNWczvmf2YE+JiaiIqraQBdcsNN0cH8IQyE0/Ag37
O0T9rQlw9mxL7gx4QWrvVh6wctHnZHTJDRu0sD4OwbT3sDodyAfR/hTOffeWDnKTHI9EumD0z7Vp
rCL2r1E5oClsrQar4gmruKEGjjmK4HA5ByEFAxIkZdcEELmxTZGlLF449IpLmLJni0Smq+NTCCKC
CYdg8ZJPdtUItpAjztmnbSvhLeFex8OpSUNqqyddG2F7fTfPYuG9ku8bnsUF3PvPewmZK8GbJt7R
03MMARSJ3tTjg2+jFr6uFQI+8pvJHbVi5Ha5GoexwGk3IAIYNIO3zTbMDfGx98ClBU/Ada6zAWQ5
nL8wCunqt8vbIoVmjyjNkuN4w9WMq2wb37/yLDlG8Y0HpZxuiGy3ahs62q3EBfBqXcQKtUcTR3xU
V6mfrLh8jGBDyoKu/7vvJBlJKIBtrUw0D8GWtygnG30Qy+0iZW2LVVRpceIpUhsTQcbj0KBv/D0W
xz30RcboNhR+K3EXp/Zk39IuCfCQxRFQCyu5B8mNw97JBdX8PA/yPVJlzWYLKCgaTuMf33tNXgSI
gRurYYUUGnjVnI/eCU2GTbni1bzDH7Orgny1/n98UtrPbIxYK4ihV3Ereqrg5bp1XxKorMAs4sDE
q2QvEcAg0XJE3Qgbq4a1yoO4exQ08XFuNpYtUYFn9IEDpF94anDr06PAIPbft6ZYC8Klzybw3VO7
8dNoCwZw3w4aSQxIVQvx/Oc9TnLZGZMqYHOj/odIrgtsKlSctEet5988M8k2gJ8mAYX41RHhLzac
VROzLrRN549O1XZZHAifi2gnnIR8nLKCHs1lwZ3R2R/ieP4rk/GIgbdqnVrPaE9eKUMBD9X1Xwns
X0mdTtHDfKr78ZGzYVgSsAjagfrzu1UiFSz1BXxKU6gTB3XZfH/jNjVYjQ9Emq4QPDrP5NsqgEKM
xsLt0uAZicQixP4jiRvAC9FmRHoJ6USOjhj+A7RSxPBqNfs8kkxZ7tNnM0kwDt7Gf37tbhrfSqXv
HUHwqqe2bLKIZ+JEJtUzZ4ha0WnvKRZtKIW0xEFr1BrHocYWNvBbMG+atC2Oqo7rvaSbzexo75Qp
t4a1cy5gts1kMPMdq6iH7H4dcQV1bpmuv096WJ2twmaMChIHW/s/VO76i8Cg33M3vJPhDwYDHM+D
Y45jXXaaj8MIJOqReEYrfm5u5SaxRzBIqWc44v+qPbtbT+c8NprhkgkZ+l/u2QnkdoKyf0jW+jtL
RjNXTXxUPkX8jvNRPkugf3i6bqQComhNVR7bfz85b2xnA4NG0Dh7/0aJHwNvizr9mYS1aX33MVRy
XzwrTha1GSULKVX2/S8kSvSt83ZwTtZM4POz5LsGKRNy7Ecci88Or3Z25xOjt1JU30jTVClfj7Mb
tdDNOWYbr5+UejvHMUBfKKvQH0YM9S6OOd/TnJCGEZCdWFp2bkEpYTUEG5fdtbC9W6Yo67mM6Dz7
kEH8KVcyelK3d4p+J8rava3qKLr+J5rx0Bb6HsRP3KM1BBeUyMgMoQrZIm9HZ494Cdg2+36eI5rs
qwuk9ZZyi/FjoXeV2lMenw2CHQ4aruxxXSwRmJwdv5st0wynHzr8I3IR+fRVRsqA4LuXGG/2dBjj
PJmaWddFPtxjyF72RFgIPmWSK7pljRaXcTNnP9gCzvZqOt9OPpCGmDJWn3QGEh8uXbstdbUmlzjk
LHqR1fNDWF74uEJMtTanGtiWasmeUybBK50EtvTwZ69jX5rm0epXfchNITzt/SEIQR4N2bJ3ELZM
OaDNZTeOYj/QleKqL5Pv6F45HitxyKsV0U5R3MiSKXQM3kSCwZbXUAMCtIbUnw2miuQt6vlxdPPj
DKEpZy1Up0URmrf/kshZqI0LIlNHx8X8RuIO9jG+2MpmZzVr5y9eVXZntlWykVBpVywQX634zwM/
0awkWsS0z8ycmJa5kILIUTXBkJkNNYTQKV5t/h+NDgLT4zOwb/WDK6QMtr6h1ls8sS8JvfwapIcx
YVjVxdOJsVvgATDKpISsivYNjELj2DrGYgiuhJ9lQ6UzpRBBIbCEaQbSd9M/zm3kT7F5eAknpn7J
A/5Emo2UU9bWuMH7ldE/+oP0kAV8Svz+GdrjULJ9qdP9puakY5ukepa4PcNnn/Dxyqou9mFbCBT6
L0mGL12CJx1LGLiQwQJPoBBDrkxWa9ACFdUOCTGpowFDZk9AT4o3RLWyTMkj5b1uCYXGaDBdBAJw
YDSjKmbZdpAC0wacjHM6xJhQPoqtt+Kfn/iRm7WWArpICdL0SxszazYWfL1VQ6TXBl8wYDYND1CY
Wa4PQnSEhQZrvJgOKIxenvzI8hOB2uEB9deITdAnIN8QH6I4e7T32qhaxcDibpFcGGdZN/129iZc
mwVy+N52CeQgr9m/qQdLGpGNpdy1RwDjyd/cA/sO0Uc1IcGChOBXfryUGZHKhK5FfGYxs7i3Le8O
/k96b89tDjA8lYvqObWSpqS9Yj36n1WrC8iN6ueEKtvTPd6aqkpjmqKTOy8CppE2SdXo800Y7xOy
sUqDmSS4uXGPkp5bXCyAifpRP+PY+oJCGSyACsYTeXV1N/q+OmHumYcetvp/xtGq1jQ8n00tJ7RF
0ifT8G+Clj8oK1M0nYRQum+sQz+Cg66ov97NfVAzMd8GgxfgHMwazYxWX74EQnJ6xvYmhK97xevK
22y3OHjbSnqGHSB59xgKzA4tlHhN0yRFVtENDjXN/Squ18QvURHvzdbvJT/cClozSAvA+mmF7ici
kZkG5KWn+69DGAPjCeL1nTXO1CVjrWrRwd0M3D92+Qxoztm7al1gNVQ4pidDYBtYoSoKoGs5dgIi
UVMmLwe9KVXt2xyU577q8mc6VBZYqln9WjE7h+4w/ugZpLpvQe10goIsf/Vvfv2LB6Vs93QBaOPf
fIMmkWIqlOCdKGLfq+yiE6WNIw0rMcqLUlwMeNJPak2bViOEQVbiMoTOW6sM5nPzSSxhOvtMoXY0
h/z+pUA96ToLnDh5iU0uR2erw+GH8v8b05qWhlisDgH9n2RsNWHvtwvIgeORRLXL9X2/8oQVKCNf
Y4VqSbwwVK3Xs+ux7JAQOpeco+O2pYCFYa0Lh8xU420f4BKGraDAN1yiX6PYkKKlfKboG85E59YM
so5Snp0b6EVFVou74otGK1hzwgI1g6a6mdo78DBInL1PzRvd6YLW7lOrQ0OxdRYBMKyuIKiQazX7
xhC7ccn9f+2I
`protect end_protected

