

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
L9EbKuxxzV/09pnAb0OGW9DxPQ+o+m/MvX4x5f3JCiR63+KWt2eYB17k+9mGgVY+K1VLxoYz0z6V
YvlDefublw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
gJD53XIM6IXGcoGao7b+pChhlJwhGxOuVwSTI1iU+aaEVIG37JelabzUSiGlwgboK2Zv8N9/EzBK
Y9pDSGcMvhlTABOa75VEGmta9QvVzRVMjXtd0b/jrdUkZar600zvkPbB8+QESNshxT7B96klkdIo
XvMdlDR/SEQxmh4Mkpk=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
uMh613zg14bfl9MaiMXKdALr5q+gvlBiCCfJpnudkmj/VEzNaqE3gABSgWbIJEk6l3XEblsHwoSZ
2eueijgOoGBjZq9eDXqLeir52M0Z4RoybrJFqX7YgYE+2quggoW8XJjUPK7bExWH1Wd6un6XRwZo
+XQ53VUhkTgctFKNHRr7bEqxJa0qk8dm+fTRKVmCc1Tr5X6rd28yRrr4koH3+liBwEPKquwcMKJL
zK5B0g+bSiHJvGXlQQpKzQNF3+4MebcveUUQPOYG2FAjfRJs1t60dgE73q6y3I1DMI/3MguCuvoX
78TA3nOFRYGLkISVFXDX28xYA0EnciH3BlzGiA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
2ADp5V47yVkwRII2+UsRY3zvclviExupZdil2h787eVOjYg5odQlZCOMnldkarIbxDBoj52vjMGc
rG04pAKa/Z3oDUnDkDe8ZMmBI29kynugqgc8aGxYPVKp3KD8EvhnicB6/4Tt66g9A8WsjHtxXLuC
0ImlGHU3T8u48JygeUs=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
s5k0DDcwk1Yhkk6mc4rW2ITc+jBCojX0QPFrzARjmvIjcmc9EJT8pAYSdJK1ykoSIGmT8u4U6vaF
5pchZ1NWV4+0T78Lu7ir0M6lHPYDFRgXZTR6CNdPGqAe+Si56W7NnXEM0Yylf/w4tAQ0u+05yvCg
wK+mPCq/91Em5ZiPcvKOHOdJBSTTkSYC7/n0QNniR1mBmd7+dgsFr5yshClYY/q8HngDDE/aNYfx
P9AT4ECjL+OzARXCnbTA6RjbHEjVx1ewIc83WIXkwbZjUYAzp9rYNjFdx68zjq8U1XW92RXAEXCc
AYKv676uVGq/WAryucxGApaihL/izu2+HGUsYA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 30640)
`protect data_block
wRbnTFBAZO14DyPQCXhlyVz+c5f0avdsdbfoJ/wD0Wmv3FgHvt8C99rz+iIF+qXydkzWu+dRJlZv
c7XK5ApcnhZM1XragtE0qUbY2VhVX1QuJKGoqNCj6C0IJsm4ExlNCxu6ZlM/TfFfrY8gnTSZWZqs
36aHZZQqNHbZHJmqZOhsYTQKWrkVGCOyQMmuCoEi1Pj7VnoGTtQbwVkDTunrTkDFYXjfODPfBfcG
PfvdMoSma0OjtomjVLd7g/2FZcs7+hxq6FerZqUrR6G3y4ViMalmNocD23YVwGKY6Y+NQAP7s8VD
/RxMZlkj/DlX1stuu3tMKRCzkmcYErM+JQV8lGsPSWtzcHTFtzApCBmfjNP01OFjOxePOZOSsCCW
I8frF4Lz72pmnDWwoAJVB5jVdb6Erm04fp78/dKInTuIjBc/6fyM8jhwH4XKuiz8tExb9HAwMwEE
+CBK6q1e5KI1U9GF1FclFpWmPTLSn7XZJ84v+Ha/AE/NJPvN/teCg/naYtcKKEuqFoNMxFJixxZl
rCppzt70ut1Hi8bc1A6bCoPydiZ4+7b2kRuJ8gljR8w43YH5SCLMEX2aDnnF88ofbDiQlW9fCRUP
SLvKTX0JuEvDhDaK3EkB3e+4PG60EVDCOL1hMfy9YhnuX9ZfdonmZew5+UwfKeQ7HFKmdOtzMDes
ma49tlyzcWjnOpNJQW7j4vfzIG+EiND2Izo1IeXXJ1LCKdEYl0NAeGuZpvBds5bIKueqvQQ4MRqc
ZkKnoGtwsPb1rzvLA34SkuUt/92uAwiVDlr/IjPjT4K+jb1PoMq7k2UZ3NToppQFdof0/yJnRgS+
7xapMa9jFc7MoXWnhMhK8OgI5Veu8F96KaVnUa9x3AVch4Cuk8qgGD4IH8RbSmJB3uvZf78uDvtI
my3/8WEYg2HRcu0N95KpAuTx1YXh1sQ92xUX/dhyxrSWDMD6BuHLelQskd4dTrcZwpZ/B5DtKxaO
x3yqhNsaeEwx9q+eb2LECVgVVg8NnmOZn6vqj2AgMgj5hgL+NSdfY7BWyPtGGUinn7bL54ZRHfUX
lGBtWU7PaIyyVMZkD97MW8guDLMErnodBEZ/R1VRosLCMXLlYmbLHfxHlt0wezq9c1lJYUMNb6BU
ayFHNK1+16UZ/Vcco9dvZsYbXnSArMOQxhckqWmzmGQt1S5J6aOPvbhWuU13C5D6dpuWP2XugTKL
tXuqDNnL7zo2frOrw2GTZ9lS7/7ShuYozS1MyQki7Q5MYhybBVSWSyQNR7z7HuDTRz1zV/jm4TQn
rm+1s0TZ6XLUTuqMRW+bLVzPeFKhkgRrpLffxkoVcA7D0HXLlbs9GyK27p3RHLJo39GjuhS0ejOi
h4l8wwDk/VxMFNudK+7LNKz29fVcTyDiYT2z+XsSN+J/LJlz0T0Q5e7aTbALKqpV4CNNrMvcxJEY
DTuW35WNxRSfUwhr9g+sgD92d70FBGXRvDojGelsZXFUtKfxRkZda3M3ilpBZNe1HSCJ+ZID0kuA
RtQJJG4ef62TNNmbU2X4MdRm97qUM067eTJLqpCtMamh9zSVcCFkM2JZy9NWkQX6DSE9UgLyKR/a
4mB8KN4FImjgm3KxL4Weykhf8ZHfRzF2MaATIWfVmRz8/tuObUDswIb5VT4PrInGqiyGJ5y9I/dc
h8TH14cST4o0MG/lVRv8jxto1rwGqTUcyPVl0KbuT/FMaKtiVmI9xMDWM02mrJ25XrlRIekz/PO2
vvUeNRhL3FlYOvlNuxzKCft3Ao7OuXZhvZMOc3MbipC6LDZtl55MfIi3XySlRa+UvK8w4oXm32oz
rhDkkHtKlWH0Ov6ddyCHNonFgVLGR38cyz9Ags/o0F+F/dv1NFOebp5zgcK48w1mtJtK6op4wRIz
yRbDQeIj4f2ZGv4BWnWoVJvU8l+sk85XJ7r5G5ThxjceZyUgk4pyhOgPF/PdxLm30nJ7SPwwhtpg
eMx+Ppk8dqIGnh8SyoyCmrk1AqMH4Ch8fxBEt+0AracLzmgOX4+IatYOcj+q+VEvDsfteT3hR3M9
SecqBOEXV8W1ZQirJmwT7L3IgmsKNa3WWENkisA5SmbKiD3cpKKMVwdhaDLTDSWYakHP1YUCbl88
9m+l3ecNalImgcWwXVHWyB281/7nTL6/krFtC9Tagycp5QSOoVGsv0aD9rQJUKadxtqZ9nDMPN3S
jqIp/udGmjl4GwN1RRhJr5Ynw5/YQex5V4wfyF5DB6O/ejH1orMklJwzuTvvdg7QB6fUNJrXMlp2
aJFB3VGMn/LIxEFp26jOGr/kODz/W/3kN8Xe5FBDszo/dbKOSIq5rTGX39HgfF13+1mL+cxjLnSw
/IaH32kp95WPKC/RFUwMTHmP4cq/7uEKLkVipNjd84j/kn7j9qqVnlcN6z9/bsGUJrZ0WCP4zWa7
IQwl21gEbLFz6mxM7ng8Y4HC8+MvdqB3bidbA+Bf6YFE1uHTZuoCQWCQyUELytQCi6GQoYJrWEX6
Far7KGgUlGEJVrU0IyjJ4FfwrRp9I/0btbabM/Z/Zc4SwN+b62eGal6Rf7CLTRJTUDrC8rjzTivw
m0H7Yul+h6nbmcopw8cwrcL3vfSScFTxHY+pgn0TbRyjO08SRH1RPZYvoHNWKu1CZLFqGWZDYrIP
1SzLyqOV0nDqTPJyj6aE4XcDA5PbvNJaYtnE3JGPsuNLg5ZtWd1Uk53hvBHId4IUS0L6h8pXFZYO
w6SdiqGzssfgBSzIlYUleBvuIn/Nm23Mr0qLPLEvddbqAjiOOo1NloylCUHGbrRrkPZ1UKxDmmwD
CzIaElrm8AWMjnRK5dWf0yM0un9lFlRyJ4TaHY/0Utgk2NmHWQcT6Fmo+B5//YCAU3h2bNmXjSE/
E+K+3enEKPsean3wbZstet5io/Hgctht9oD63rD4I0jPL1PSQ+wgr+ep7KKjzPRiXrlucSN3MtA7
JiN1BQuyMBHlAsskzTHHfulf2RIgFQF6oL2adUaZrq//Dsm+FIXBYzPVob0yJwmqZIQHJwds8zaC
xAMx/JyDOPJu3XxBL7YulLRlnOySjtfsOHTBQX1P3b/PJsVhq55lIiYXDij66Iu9NSU778MUIUxL
C9CltOiRZcVEs5glVvPPl2Ww3m+3j8M2onyprEoGBnroh6ZhxnCOD58AJNfMwmoBWmLVRpw1nzDJ
0Cs2GXm2mB1FLrUh73geK5197Cu/nI69KZgr/7R0f6tqywgxU2Q29mhA7ca9EjNeq4PHUnJi0Hqr
zQQuX3gDzqonwOLX0Vl+Wf4KfH9S77c7e/EXQgOKnRiFG3VMvW4DjlW+5xnvQaVUQcVBDTKIzYlu
Y3vQwyjqRu9H3uVPKnb6ofjvrM9itrFhuUci+DdDdeQXkDVgNZvKafM7SdOHw+GcnnmD0oRVSPBd
4esJw1NF/F4j/cRDN81d01vlslfT/U9qliZ1gqD0wnMXd2Fuhpfjv4NUNDys51xBEyHqHu8OI0Q9
/FWEbKhpSnDi+9nmnJ71oXsoqVjOhAciz+A/LhvTn9TgGjNNd8hLvrnBO3yOStHRHgS+C9hhRI3G
vuK7y9qw7lyb0kpGwDmbBXcbTTnMhJofECjUJ/J0Vf/jKudMgggvPmzgAjr7adXfQmzrJy1sSjLY
2N8FgtLjwTKBV5UEpWnsQ9BAR+DhdtDvbce3uqUuIB/QuU1TzRPpGmisySFV0Q1vgn/6hwpfr80Z
3LsDrSZmHWVYv4j0TiXMViP5ExB2iaTBoUgq20zKPI9TfI1lDdmlxJFEarYf3VAl8PvIa0w44As4
kXNwf3RAlZqq33ifKQdex80YyRBpOpaPMpDYgYhdqeEK0COJGRT4ApkSuR6AphD3sgMhs0nMdnyl
/bTdMxlW3DiZQdJ1qvyv/hPAxXeSnPkCcIb3zvA5aoXbRy+PzFHDg1MupQ7s5V1wiQtuvu6BaAyB
lDR0OBQqo0BXGRdb2obJnZSJV2N6L0NDNKGVqIIvOoYBczJIhLCX74lrypw/PSypXUZjnQ5pOBEe
wqvilFcum1lIp1lNKX1HTiyGtRgqM1aWTTvlg3Cw+5V1KGPeSdJ4K21I0iuQYDNa5k2VPDWos3hJ
PxQaTmFWDx+NjT4Qxi8O6CY9gxpFIOO7aAgdsdNITWfvcyCY1VbgAgsDndPKQI7Vi4ffQoQnIoJH
dX9PZRzBM0PP6FR6FmJKP5YnCs325CbMCKIMcy51jk1oOzIOMgnVxzl/u/GFNyguY28qCm2/q121
s5DvoIcx++sNCdwnznAZlgowixJ6Z91nJZz8JQU/eJgQRrwlzoMgaYhl+4kS0pRo/jrVobMU7aiT
XT2KmMiAl/0wsQdNIwDt0xw20HNFCnoGWM5euZThUeujv3NgrTxIuAwj+79ejFYBm62EpHIb85gY
6NbvTEQNOMMkrreMSUhQJYsd5+HO4Q/2sDyKW44KeOw3Rmfk1Xj7vt9ib7ygNy4L0SM+jaixTGnb
5uFb/3DOpk69Xx1wKuPLX1hFE8r9f+lSHh91zU1iZ9XnTehU7j61Eiil/oS7SfOSz5RkjMn6DqlN
13eLeybuuqAk7OIRbzc6lMuH1lG9sLTyeGzUursk+hx0TV9osv2hkdMVm7X04UJgiTZw031SxN9W
KZ78AEAOkcYsXBUGcqgSCH15M+PIN/WJo6Xfrfx97DvwtzIu6NZLVYYuxA9nT8Vzqsm/Rz7FA/Yi
4D9KdKjXQdI6luGuzJK6WG3IDODrmUe+4g/07aL9Fmxsl8Lg17rP2OJBYN6KNPRpS6ziUoNzUjpo
j1cqtBUZPbk5qhWaM7yXeRmhl0dbdEMkum96PX+GtjLPj/DXlP4wvJxRKNnGoSCler24xiFkTV3P
FbnOSaopzTtCG8h/2Qw5qDb7JGaiye6DX15lscCcNb9fg2rEStoEM1mh6N0awmmXA3/O8Gnzm2s/
bBOqCXJu1scCzHGYhRlXPCs9poYBc8+yHZOx8QTlt95wxrmjhMcaBBGL0V19hCqwrcfax2hXmCZx
c7856l61Z0kRdC2G+wl4/mXsu+aBWL/1S6J/jU3tGQYY8H3iFfqTMN+eDv6PAYM2sGhWCYFSV2UT
gnBmE2mLec4jD7wpB5jE7Y6qRc59ebawaoTC72s5BX2zVNOpl5BLkinlWMUBZuBYbkclnJ+91x9G
OdM+dBTeP715+WGFExwtb76J/dGCHU6xtzSYDBXLE8e7ZtqSSjq5ZQxBKwgx0xhlBHVb/eJGB3F5
esMSmtoZhGntMe4O9hzRpJp3WYz7yz9plQ2H3w2laM+8evX7SsiEyEvI8xOA2SxSiTGiwPmJNIi5
IWv/FpYXvYC+qfcVoaWGtN4p6oFWB70qA2fNVFLH9fouk4L9SCjJG580KM0S7RIrb1yX5Ff9hZo6
XmNlmL0GRolAjr81kvtcOdyesrTKETwVp9ecD/IhmaRoVEzGEArO8PaIBJbtFE71zEeC+UC6iRF5
C3B+11sw98UgjEiHMD4KxPIzJnv1KHUdyqWztsg2yc1UyJGf5bZB3i/FX7VZ1GAK63j/M24s8inY
ZfpEAZkcwly3TnbLan5PQwWYKRmwRxDFF6GUBDJm+On2EGn+cWh6V5B7Q194z2Vz71TdCm1B8++m
pkQcq8GzN1SEOIsZRA7DyLwl8s4QI23aE22jNgl31RzrIEYNPE339816ja25lFXMiNgoDQ4rZFct
l1StF3LDQn9hQWkOBC/YbRfgxnhQmyvYbG+FcVtvEVK+VyzWTyFcx2cyyohYABT3CKrqpwcl9Y6G
eMloeNtDNas73camAOpVqBcCW8ZkGNk4kAy2e+aVlQ5t3ey+2QZAbfQ6u0F1StYCt5UsIfgsPgFB
JjaA2XVlEAWL+dnvWKoD+IvzJdr5mpq+9Dfd8vtDTPm8BGiGkEdAnOr7LD1CDp9jydbwyDLdVYfg
FZAlF6//dLFhEC+IVwBP65mL8CnvNjYlzLzUvaj77VjK6zdlHYh+zXyDLlNPkD85PdKkFR69FJI1
Q8g6+Kg0EmF8H1KL5lnnMnl/Yu3oDDR5gQBTWmh2F2Gz3lelSd5cJT7MKKJLwycSqZpGs7FiOfeH
HUW3Ft+phqgRbkPJIFKYKhZHS8izFsy7TjcO3knSRDnxReLiiVrMY7254yrrFaV/qwzPc9EiGUHK
4nen7m8BfBWTPZzuNL5BYFcgqnDzOddmxof0hKcm6kvDfRrJIXIXXs2P/goPnGaGVzvIO4+HkYpi
1j0dYOhs5/HmH8CkO8ezK/t6tf8h+GwQTkBDdNIStEiGyP0CJRdBeKgxctOXk50IWI12QyMbC90k
Mefao/4boqFhBcOAcc4SGguUhKmTvrvfqIUDzxmGd2pjfTecsd7qtLsl4z7gZH6BAaNrvoeWbh0h
JstyMDR5xPZ3qZXbBCZbtV9owJcyodCV142JR71iZw0lXI0mmCEScDZrtfCjAb1ZA1k2dxLN43Ay
vWdZcgq7tFxfHViZLDV09qW846ZY+LeU9aqrMXX25frsEz75ZLuWNBEAvqmmuR5jeKQiWyOXBufd
i1LUfNyzExC/BSWpbHz55GA5O0MntTGu53INdg7kSF21/4m7nYT+t2/Fm7GWyLCdjJXFekdbdpuc
cyODcwbvHoSqW3gs46XIuM8dd1p5IQIEWoPBYKp6o5iyo5YxDOSemI+6L8YcvxCyv/0FfMdF1ncr
GWOI06BBCqL/HlOHCqvXADaOh1SE76c+Na1owrLTacuO5XjXVOvhDXVPYXxCaqAwcapI1kHrkjHs
GQvA4yuiQ+mtfSA2BGi3Q59Ebc5nobW7Oy0/FC16scrKNmdVkkUbcKPC+u18Pic/DzFiVfSv8jUf
LrMk/DJeyJBYeqwhcEvpgraK7Mlz7WGNRSu8hceOTjEmDONdOFaF1O9mkAZNQ+hSyMAOwzxgyDKa
EYwGV3X1U91CYMwR/zXJ23xquzt2nbgcC2LKsfTX4or7STfdMuiHYpgkB87fMOxwuu1+7VgzvIVf
9gsgx90Yr+ujqMpgBhh0Ry4HHqa5Z2/kBfjHfmybquettkwBlz9rRVp1khJab6yxSKi96cPxJqXD
hnoZWAde/6O1GisBm6au85y1QYLaZFPoDsVnGyVa4lntyEQ/CL3NFJPccVwjpH3pQp0jsxKcQnLM
Em9jIBqlWyLQAE9W83azyfT+ify+QL/QaDojjtAZStWYoUc1D700u+k86499D7WBcY1qv8KURNTi
Pzf4X8r3kQSuUcyNZkygnKsw9H6xAAuz5LRarWDd/qVHflcx1MScZyiZkn1WHZbNFJMMqQQa66B/
wQeuujP8WWhu0K6G3tmPe5YrF5p1gvR4jOn3YcMUs5VO7y0tvHLWSBxqbYIwg9IudvL5jng5bFXY
LKFbBg+tCTTLJeSbSRbx2QZXdmxsAXbTZLQE39F5MO25QJaUXUyQW7E8LEoR6ogFJPMgMPGisxSD
UzEYHqeFkf3ujX+nga6d7hUxzWXX6p/uFHYEAfc8q99Qm5/D4uRxJ2xBCB8dYVuKQ6j+MpGvXVaD
hYRRwo33qO8/9usTc5vabk8LUGwz47XvBEqFaVwxyNC/SBGnF5KL1ZbthFKFDJGZug+5CTD7hMo/
JbGAcdacvFgvRfAtVDnyftpRiNAuk+uVWY1gokGBVIF7faykwplwJ7i6rrT61Ag2EnIWEto2uy/r
PYApwK/bkgr4tHzwyN0RQUdJvNGq9JvOZRlH1c8vh0sTAthW5N/SG4vfmVoeD77sPsd2//w+iZZb
nReUt86B1jXTrik1OAKT4fH4TVYx7D5rTpYJA3zvBZCOeFIELVYq4yUIbYaHzhIh6DOgcJ3mCvFD
vTK7ae21+OEAXig6/r/RnGhHGm4kd2JQQCgHSMrfou6qF4P31jF7uWPuQbWOGsoN10EgsUzTWBhg
vnGLkCWb5f73jvIWUm9Z8oeyZQAUogmNHJtn6n7tn3dPe0Rz4eY5BtPFCGmTJFUSnAZvhOKaPbX4
t0ghEXrOzDmktEsSQkqjXk5Ej7OtaychKmpuTr+lFGdcKzz0KKgkWPRoCGDi4/XGB8tQxEwGsGa8
VQX8v5KKtDu7vootkahqK5JUcbo0UUypqdYggc3qXcA6lohxBPS2DbOECQy5uAF3sIsQv5oqAWN0
7S0G179GW6Q7P+tssxhjvTT3JA0xFNOuzbn5eSvbZCma8BhM6wYf36hOqUKG4/dLB0/Vq7GksWgG
lRmUPaQRBmkWCr5GDQfmJeA+V5jArbzpIi3YI0M3m3Cgh3eSYEePAzZaK7fAYNKdbeGuA3epqdRf
TKoIOUCI9n6NZPKtJ68qIQEZX73nO5UujDsDnoDEjqwBLk/wu2h58CK9cGTGGmjuXuBkpB5cf2OP
sfCwCFqoOKZPwTqZLAMCFWzAFYIF0bCJ3t9k2cDfZkmllAKwwvVhP4liXDh+GPvKBvNSOqLJfdso
3yKUZS4HXzhD79VXOL0iPHHK9BVvANjjEYNVk8u9togsPzpL2Bb7oX8JxKySwsvn4K906aqQKLaP
BcSc23fXKno1x3TqFfUETkYHXsczrRNNyXnq8tbVtVbHYbou9UxqsX7FkC1XAnapLa3t08yX3hpi
ad9QDyKnRPypRJb5qutnykAJlHMRwrgljlgvU/j7+7Hzu+cbjZ8KsBmTBYJ9cmU1e+vTewovFqXt
NNoFrII6NDWzsUfDWA++RJOQuoDXERgpchh0kfHhTtE7Nn2mTsmvjidIJrVGaOJi9gd7l02EMG6V
1F7GBApUUIcB34VprptDuwehF7dDsxJeDBlONOwAOKHJvmWuWcfM4uaQYkgn6FUlrKSqYV1hiAHi
Ih/WpkaEjjd22lN6andCPH3+KmIwRZuuLWTUU1RtV1kvmMzbj3dg7blb3JCLMwydyg/dpkEsQRJo
ZshCqINaR8Sffzg65KtSM1moe378E/pY4IrjkMgo5i8NkaqnGXjVzGYUfa9B1ZWH9c3jzezQzUyN
K2sWUhw0cT/ErQ88ASnPrsSvuedcndD3GMqti3jyHRWOxp70+RDaXn/lng1Uv6dzYrq2dDbrHHjT
pQMsqTSIfBqeyFq2oIBCzNe4Xb+06Yb0gOJ/lHpf+5LkooXCSxMoW1xPD7xCQxTyTKfY3Vv2PpTs
e1CpkNenDwyAAsk+c1F+l65e+R/pLkwO/i1fVnZEWXW8JltOFnv56RZ4f1ZJkD8TXEUbviBMSkLZ
XpZd1IPu1SznOomDD9OHeh+bJrUI1B85VFfd2YpuPx0ftXmFy0otqgf/5DdpQBT9C3RS0N+oahyn
mXiiop7h6tPtHj4r3LGP7AVImBQ0kXqyNZ3k4LQaqpRuvwQSl4x14xjDbbWVXlOfSItG+zE7kOqQ
iKQ03ezp++lJHsAFSe+kCkWABCFIQNOvT6SpRjxpOmSmyyfWnQP35k7WNcs7zB1416Lr+B6JWn0j
zTE/rmW5PxVrJgUSkAYQPDXemr6qcPMNuD8ZkOV5XFZxfUhWCepTRpeqRneZYRTCbkGBgmPD82co
EZAT8bXEpDkvuWilL0ingqvSp6MdEvcGVtGo1bgteJ54RXI6HVyzrtXyjnPSR5aqEJ7djGTsY3Id
B1Mrb04WWfnyBO70XRX7C8Sll+OFKqUcmHS/obq9eXJYmZCFocOv7vpBozGT3ovZvrRTfMJ7bbJK
0hhZXfJoX8S7PsQuofRZFd9NLzD2NFTHea9HDKZt2zvvjbSYYIAO3bjNt/wUheE+2o/6BEkaa1w6
S84h9OqGoFCaytODW7c+ysVVV2jHmufhk3mpxhGFnfmrm+fnZeNOuAUM6afOgszIAdPcx65Hiki5
npbqAjfFXbTNPkpuNAjgXjjn3LCrH1A9G0yvqsM4n0fGo8Q/LCIk4O/GkYQPa9oTLJtDPnbFHooe
sZar/3hPyjPqApUS1Byww10CjYtB+n4lDp6zJGzWRP4Pfx8PlpbqzmmAc0suYmdyTZhipHI4MFH6
Emzt8qC/0dhF+Ud8AFVCdwAitrdcW0NHJd9HpXPZ9HOoPO8vdVOmgMpUkfj1c+mgB24YaF0RBFBT
v+LphIi1Kzb6QK5AeuuRsUgACgj2sp4SdR12C8Kp9wLy6f/f6iQnI6E5KGAuYdbyVMy8mfdpdbKU
xODL+NKecaG6k6qPLUEsgPXoVvcWtQPndeDib12uggf0r2KjImjfCllHqkLcdUcmCjvKljfV6QMq
rgpBlsRKWAunswr9ehh0VrtD6+YwjXHX0YcIdmKA7zVuBMnedZGOu3pk3yiULPRQAjrCk4C1+GEu
ZbL5kV1ZQEfYlTLYdv2meaQrSeD3jC8oPPl8PcTqQ9UgdtMMM1HjA4EQxvhsCQKBX1aNdafk8r+M
bo34zg8Muu6SGjBW/Z970cH1NOXIpnDEi59pkikZbApB+/GKBgTvT474qSZtxZPxRnn8Xl7ojURH
/nME1Jhe8lEBCGocE1tn5hs8g3T/6mie4E7+8WaX9HIHhXCHB9fWhaG1/X45qvhtl4Efa0FOB029
zLG4msG4Ei+6c36ZGO332AeChF3WfX3gGU8HXGpjhc5gRT9aj1nu5yNT4sO1H7j3NGhz7vf2LE0x
1or+ncURq0CdrD9tDvY9wDhTx7LwtksOf4/cRU93C8uzIOqpSf800xoGsvbB0gLItoIG0imz1rr4
Gp5iUmNMbIjDgh410fXsuVd6nolUkpu9ycheswHkhEB8He04XVsJa/aE9kghhSCGx888N/x0FBdw
U4C2+oKo7jU/qmiC1KffiU/zQR55H7nXy4eTJiG7AnJwb9mqQ4yKGPGswR3k288rV1odkqmqdebN
m8SKooo08G40DaTXAeqrL2A6A41oCsXJ8oEPJIPrPwfLfobVjGUZKF4Q4NvvOF65IOio/RsG9f/3
7f3tgSCyS8ZVNdaBgAjyOEAcP7roZpJ+zGTvorEFHOQ/FrAtpUsX3icDZaH16W+u8ZbNLF09hOsB
cYtthPtlHd5cxjW+PjL1aVJDh6ndnEYBjWj2CCoLX2GrAVQpCA3YkLA/mBDplOYhJxt39EbZ7BVh
Arm+Hlkb6BYu/gwk5ahbm4UkRxelBt4Mu/GLauBV2tbMz/M2KfRhTu30dpPelAInHTizoZNM8xDm
aZILuaqntirFvNM84RlKeWJIgrDKVVSoq0vY4gqyf2nbiLfNOCFuGlzFyJKceikuDhEIOyLvnN+b
bUD77RCZsHbVACml2nIDU5JEyd8Wjl4f0LjwyUrbiqb5s59PbBllPzJU7JNo8JnRoPRyyTjJnCMn
lAeg+BraXyx702GzNwMPbTLIC3rrGFeC9ZYY/mUEIqnMILUmRDVM3nJt1maJuhmoKgHOfPS2T3la
Mh4QbtBdsfjToHOFib72kRflnK9T83jG9mORsDZ5WlPnbc0mok03bq5XLelFoIOig8zdlRy2sFEa
UyR+vbA0lj2JvLumNaY01Plb56vFlh+1pnU0Dzpmw6ViBbv1KY+ppB9O6qop5oelMuNEKCzPuN43
CrMykBMaBboNaFxoqvquhevwX5HmYUk3IL+0mrq6I+mR2snPq62dwC6tMucCHA4k+NsJoRoItnaY
kVAv5dKBbXjtwQpVo78BxVqsMJdwE2LcS6ZCszVH3am+AegaTPxxjo9TQoo/MpogvftTI2p39+eK
6D2ncnYXpGAtBpJnKfW7hS+KH7SkAgtBfdnmAAOjW+D4FknXkx9r1ElmdSSWwMibI92f65E5ur+Q
MxBBzaXXykhUuYOtEJ9Qjg1UYxQQnNW2pxC2b/YvcmTPufapC1HNbiupWx9+VtoblDGIZogBUyZ4
dv6JttEuyCW9IsDH7LGXiT9SThRig3kZbLYNwN1VnYUaaw/y/r+mEiaJzEITOcArIkAmSFMs9TTz
+J6W+YU0mqol0BOfYsFEU4dXcJcDacqt4ZO+zbDh2PitD3mpO826aIp/GStotsMsdtMifgFRX79I
wDlZwylMRDL0Zy6XvS7KfaOGUSleTgSzB8eF3zTlObCDM9IytqhEjoGhP2LABRaUSu4jAdahIuyk
eMBaVXoV6mCUJNYV9ejJSLrUc5fGn/wv9a0HVtrdJ3mcwg1WGMOk/E4+gDIdaIZe6E847w/XG4vg
2aytZDbOHyukF4RhjXKxVy1OERhHddZueAlxziuTU8LCI09zz7iAO+bIdOEdvmlH40ZkXIwd+dsc
fMVkPC5aglfJcVDbY66wRBWBAFWAS60FmjsgKs5WX4tGCemYQerUfOAf75FMwQ6rLszfpBFfaNnB
hLmpCdRjIwk+jAsJG2kNCsFlJ3l+Zr8OKWy28ZC2wsooI349M/AoI8nojos2JerZxagKFpWR7UR3
aUaHrofo4YQxWoRCcz9qd3OXCbB7qBusgDltaAHwgy4P1kSmWtTS9yl9wsKq5l+xM7jKON2z46tj
Q2a6FkitvAZYZ9QGmEXi/70GbJwIoMtFEn04SJdKXskuVAV11U24TwintMhaNB87yxaivvSx6s8D
/9KP0wHoRGrBaUxFiNlFKPWQKcevDJaH8ptgTAdxAnBoBPmwZ5ci97S64kR1XrqGig76skpOk9F/
h1lnRLm7jR4CQwEawqjAyON9OxevruBBqgLp/0HVeb9+YkBZ6knDllPO+QZvk4KBkmhQ4mRVg6Ge
7YNu88hGB9f2e3/3oQQ7gg4cepjfCweSMbfha3Iu4Pnu9ycf5GXOB6WwdvNZWYOdTIMLeCT2iUaA
t4Iro8qeQsUoeQA9rR8ApRJhSWIJ5yVL16EeivOt88a1RDZlMAyFNCCrXZGpkqyyHVieV1IZ9UmZ
JyqRM0JmhwNduM0u6ng7w+a49QdeZ1BjBNZsghPA7HfyaNze/mIbD8m9kw81vZDs8TlKwjvMPRbD
VW7w0JDm/x1RFrKXxEPHs7N7jzDJnuuvMpeWsnVISLw2aVSbPPAz7dQOmipvTZ8Xl3AQFUGIJVGb
/I0OTlITKcHZC423MK7nae/aiGMp0GPr3TUcfbHNcR5FWfoxWZOLqF6PZNx0k74XQuuZqT1bJFxS
gDJ3fgXZSfs8L/jx4PYMGuZfDzPiceZIUrg3cXAg6eFDvxo7x8jKoZZT+6A269h44KT5EVOrlDER
mtYbfdaDu5yOuWxW/pqn2G8xRr2yuQY199XjHxX35nKaC8ETIVyCL9/urkvS/0W8zj+QShh6QuMd
z3beHYZrA0d38XubI2q2KcYG76NZoYWZzgT7kzcDeZAWRUlRMq8j+Ga8uJVpRtaXt0Kyw//NvtIY
bpau5LPYD7D7jz/2LUqxzKXz8ET+E4dtJRcz6P8HFewkTKQgrkJdIO6voSmbB5cgYOirK7L0bnHA
eHA5jeLG9t3Jq0kpCY1cQJGTk95jc123kIT464dCBEx3BXTiGijqVlqaHAg9vY6wcRkDKUVNeHTx
OE79wwoAQb5fTnbduRy0Z5s1S6gYA7nYtqmYUt1Y4jG8qw+M7KCaCp3BHJVwKFJGsrpSaK9FLvBD
NR4NRU4icQWCEWU/VgVi5ejXKsy1oN242GUTyuzrh/+h4Zvc5E071I1zIggE0Zw89S+og1G+RGLw
We9NwrGlERaKUNn3CvDNEyP0o+LD+fh8kxtnVmDW8wvoknr3nE92NAWr551+vbnTEDnYxnzYP4BJ
ckWBaK3WvJeF/Oo5kmNq0Z9wFCN1aZ2HudI8GtCy3adq0wCx7vnb80uZlg7DXOCTrEOCVLHLTzx1
wXUFhckYAH9DTU7fc6cjiJtvJEncNrRcpJGXz1c5t3J8f9I1sthMwdoPCdypw029Rfe2sXgg5CFS
G2rb5/72FGEVu6pBIe/qB9uXKaiokuvAc7YiihvLMnNXqi+9nL6v9Ihry6FLjFxR8Hh499YuOpbs
4TKeYl0qAnCYt23lP6YoBJOMArNWomUvJJox0qUOGSgbnEMLb28PJxucVBF7cKpGGFD/lUeRmR/b
HHmU/QjtwDbyJ7gcjOVDx7oJpob3tCJhlC8zIqS/NI6hmT9tSAkxMcL9hnBqclALYuLG4kMe6iWp
MaNpRMSa1jcklKT3TZ9kUx9QyTN/C+Zae45dHGQvA8TPyQBBkyT8mdHm6VLLnzGHxE8rzciKlfjl
cBWptOvd84BFvmZgRuNO1Zeyl6PGnJuvYOCLedCtVblWzcEN9Qw743/Ls6ok9dxK/ErDnTKxYDY/
bgewBPJZ79L0Sty6rODv+TYPD8JH5srvK/zHn6bE1q77xFZJj/c5ZiGoXy/clYKod8K/jRgP6YQd
croGmTRPNgngNUrSOS4UmZvXQUk+yR5ADVw/lav1FPcX+FppdJ4R9ZIw6uqvzlixrlAZEWpzfbey
w9Q1aHlAEuTlaBFhVptfM4aKBlG5ZZvm1fT24XAYdz3HAMBtXKiJaT4L6yxqJOzQ/5ukJIXjFyY8
Ca4nqdzsOaay/nRF88M6CR7+iq+7RGs3nxN/CyCzpNg/1Wokq90sHZxvrsd0jCZYJbgWW+1LDXwA
hll1XEqTt009JuB0PAoo8Nr+4F4/BXYnLH4ljkldFOLBQvXdS2TJ2bVaegXKpCgCWbEYxT5zWBGa
9BNkr1PwwpSBpFK4IMWffWAljIlb43IFRZQ6WskS3pBEiLARGwFlYQGMeyUcuNuYIZg5V+tf0uXv
YnSRwN4M84j3wIndrA5ARDMGUbbwQ+QFjAlN1lJNbKNGKufk4UIJKzD+vb9hXKRgNrCiBD36VMr7
+9rL1XnNbdXaoN44bCSgMa16b+zIdiqvJYAFxFpXarZaQJNslUyx2bQlDDRf5DcJgaXxRbwMtUVO
USnWycEsL/BDeqyoqBbQws2Gvwt8jDyAiplbgAoV1B0Ph2fuWHHzVC4BCW0AuGC+uq/Kl4u/Ten3
Q20O2lBehH4VBOMt63pDWo9eX2i6nXLfmeQTa96OlPKBLNO22H43Im2Xw7OxHbC6dWNHyLiO7pcF
tFuxJRWiSPy/bZd2BRiffvUysYZIf8+K9DUt7jRMwnnRFZQjmQADZSq2fFJKhoZZMLlSonqoZC87
UqrfAW7EWRHCmcRD2hh7VO4wuYM/xel5mQRoHWnS7RhCY1Jh6C1XPFfjsLejYzkJLKY/YBqfDton
/OfMd9ZNV7h0xXBcrvkCJdyayVhWCzkCIjUBSp0GC/ydFCaszruXuKjYZmoGBGhdoWeGkR5P5295
e1u5xSuqG+68wdvO3S9wwEW6Va/BQzLyAYWuVXDQUyK52ZEHosJyNVGDAbxgUrjgum/W5QEAFsC/
Jb4t0CYuA9bZW/mepFPgmOdpNLm8z+srUJFCw2wIz8vPC7Om4Bx8uCAhoHUqjz3zAG83uz47WarF
bY32NuOOSQZfZd2mtgQb0DRvLtXQRJB5ppGTy2QmJLgzuYn0FhmT/uA9AD8Sx728Q830ABf3CxCX
rCWP/va7L3jmYZ45fcyPNJqI7LtfotjiWrNDZQ24a2jWQdqwGtXOIzuZAXsluNQq3AmxbwIk61Vm
T46zqPO0r9F4H3aPad27mwCQ+3aT8F9O+E6EULi+W1JeCjBabH4ydSzRDyUfuF7EtwbE8bvjjFy7
tZLSNf36zXfGDG+pIpqzwtHVkLbaJ6kiIX0hYKb3YWnBH9kMCStGCd5NV1fEzkOqZoFV9RgujLGS
L6t9Sk+3sCymBg8W4KxNRy+JKDCycQo6y4vIuS5vHfG5l5yHjY0AaVEEJZM/9y5xE5N8zggrIzWE
f0KR7iggrMi24BJ1S+wBZdcV8fGYXQE5WTQtwfJlqIsQ8u56bWDYfCKMwWvlEHZfs5u8dvBV3Woy
OT2D4YcAFtI0Dt5OJ/U38TuJHostRbRCwKqGQVQcFWUMiAz39aSVsDSl94nWHLKpDVkPhCsrS7Is
bm5MNhVrQoFlnlBzM4Rmv48WryaF1j4mAU9CdlW5fJbULo6VTWCu+Gwc5fMh487nipc8ZMJW2woK
EMTKvM0cd2GteYab+C/8KHKg4E5GiYKaXI/skkmtYiKNBG18Wr8XCuZv9vamGM2o6VeqRmhb2m2N
cKggXxSSY4duw6NiQbn3oHqFwWUnziScBuqBGeZY9VN2gv+0XKTLSykVqE/RPNnZ/fizUoKCFaxw
URQZCkNWHC7NG+hf/ul0ithDtlPp6mfbnaX9VYACO1y/AwwUcfqls2wMfP7ohnzhwvOBkjSZJupY
vOtFec4CqU4YzXsTK5cRw6zoof64rm6Qsri4WiDd0zVoT61hZgXlBfjkH5yuAUjApYBw1eURQi66
bqII6Al1/4eYBOrqXXPjZXa2tx/vOSMskSksjKmLLvwqEruLTuGvWfirAaDjSkZXAPX6JJ2cmkVw
PA6+SuW9NIPP8won8nMKCicTRX1hNfU0FP06XLgmsXU05DTGaX+mM02r2gL5qQ95lEAHo7HV7BVF
uvwMj+ZRtZ3SqCh78plJAmgt/qaDV1Jvz/2CD6wLHs1yP22jtXunVT4JgbHxYBNxmT/AzspTOjCl
Ni5AFl2zUK9zrXNkiwLlC3d1L6KhGlHpt831tu1GxcwjsjScJRs2YjwHwmQxwQC5djUxldgrrqVu
iEHSN3AYmkyM2D99s4fXci27MJRXC4XUPVyWxYsLzO9T7mS+QBn1QLvSksOIApGyMm6bWXBR6KgW
jIpSpQYiT5rsYa4BSYOorqABBYIS04MjZW4cNLrrrAUBmCww6avpYLFcBryCktNb1cpMuOcRepKF
lpch/BIaEFU4yuMobR4NkiduK4u3Zn0uhOw11xMjrqd7sVt7S3TeoD9ChCa3TV0u1cxuYhWwD4pL
nyW3Ft3RmoTL3EX75YLqmOFtBgNsX6rEFVlEPVKW656MBms+Z4hpvTR2eZvONMjDzoR/Z64G+Fne
XMKY8CDaWL866UsE5GsjmPPMNAw3fhNilbIjXTUyFJQih+mPuO3BC72vkiFOK+wqtrxbWfXCvn+L
up/1ap0RWy+yEsoCQ4x1xi3DKZnBPQnM7PJbYYwuLVYSBFAJVTmGejEoT0ONiezvDcPtvK0FGbW/
mn5WEBfXj9g1IB0oK6wEu+7vYFY1SOb9MLAwuZezsoXi9KocSpDiW1wKrFNBD4omeFhqJOLY86a7
GizEeAP+JJywrT7TRir1VvQ0+R2jXxPbIK/DRHmjuUy/BBmN2GemMdj8w9nO/hhgCkGnztqVYKj3
j+BGRQHn1+4DDsEs8xwC5lVKnKn2qgH6B1VLMVLtxowmSgplJg7rLYtooZEEdxjnbvYvQ3HXsqZe
vy1qZ0gMSS/Dgkt3bcNKASSRKrh91WLDXVIz5cxAgssPfD6hOYtMgbQKKGckPUwqIJvMPMCeZSNv
+fZg83j0hY8BAhmz9rQ/iGNPHHjE9PoQK6FXk0/XMOBsTmMqauvSSAPRGKB8Cw8wfSbSQWUYVUV1
VtRXwYd8y9LhJcpqWLTeAkMjCy4X2WMRLni4Sw6f+bexEWkYJquM8w/OpWl9jCKNRbnDKtU2tKbx
Oq5qFYhIqHzHBekZt46Nh3ntO4OwDEpkpYAtvKjV1f5JJHtgTePpT0fPlCiR73bdfMtIItMuy+am
xYe9r72jPSQ7/KUskb8+kgVolFb/6JQyiotVw1U3+Vl2YmpGXyz1po+wQqamRdgtq2TKTIiTFtDU
ELsAW2LIAtotLp5DLwwFaymOGmtQ02uomiLi68/TVz7/sRci3ECcWxE//VO+HJJ2FsvuHxUiK5lq
9riwe3/tdoVXHqzLjJWP8dYoPJ3WVBEmRkdPkACUlNRqB5fuCEf6HfYP4L5ET0YRdIkwBiKUc1qt
HmRfLIWzq4/JAuKcoVpRJwzDlOxIywvs51UfqnjTx7hFohn1Egz/Q6G8b4v3p5EyuRDeBJH/ZR5h
fVAyb0m8bSF0IPo6LK52Un19dgxryyc71NCT7ASqdzoN+eKu7QcSC2tlJVqRORJK6NGkyuj9M02S
1o9ya2F5OI+HA/yyYTHYNG1fWm7NFdNdeLtV9NbZPr6fz2L8Jj28z2DTYhDOlJZCIp/2lh7rxc4v
SmfapWH9L1SpPj7SVdNntGdyBvrUQKybCLWsn8Bx8LKz5p2x6JS5NCkoG9UcCHX4LeGXk3En9DWD
d4eyv7kpqJ7s8uj8toDYtIdenv0VcwCTUiD+ORGeyt5YHg5J6X4r6mFD+HsbCC+DRqmH3m/g13FY
exA0pogm5IA/pcDgCkoNPIOPf7gddnmUU483kroFBSY1cUpxah3m+wYdvrPl0+GuCj693QvztDfK
IZ8HdxCzsrVpRSE2apVk5bf56zgdlaJiaBFjvbjdlB4cGh4SQUvC7zrbJAtKlcutmPWqasr1DHpx
D6aNYB9XK5R2CsWrlSHhpLnDmoyQE8SzW+kb3vzR+yQnLVmxYQjnxHu+5VhXA3GZOMQYqXyFhgnN
9YSGXJhVvbhKJsaENS78oc6sjkYRU5H3QgB8Cgr9W4/FPPukzUnLNlw+PvB44MUpbRI9oEeA7zow
PBtW2knolitYrB2yhfxLUnoRWS1MQTwqYpAc7vpCOQS1C87zmxylZyD1n/XF3fvPqeUdoK6ik8lK
zmNUnTscZ/iZgTYijHCfPIU7yzJYzvPV1XpYkyjOlEkBbvA6ZfT2Jh9cquyvGE4VlIP5CwQ4PR1d
T9BZ/6L7LdpAX4bmPVxOIC2GbJOARICUSPrtxaKQMCuST7Ns4zbBipWuB8O2p+HCYx5CiscZovH+
m80dcQBulML9dRWhqD3xfe7r1kUqoLykPlRnCz3ZFbGiv68H44VtFnUKLPlUi5Fsh5Ked7Vq/HYf
GweF/oJpoB+IFTPpOxxLKoTWir1kXd4TWIm7A5Hx47iyV5U72BXRzVE6AhWIMb0zK8s4+2nZQ6Ly
5R2xgeV3wSfst+tISxxz0zXQZxbJZilo0EKcqov+0kj9jmty2mo0MkNBBM9ogIZEgNKTK62+1ier
aKYhml3D2agG69/5uQOLzCv9MR3euSkks7qslMsdhqHduBrwKLNSYFrgZJGhd9pCx+pU6GEMD/+i
wfV813sswZrEYD8zoAq7zVpq8zxD6Oa7v+KrPedegRgsX9KKZ+2sHsBeDg+07qXO+dGYHPl1NUbK
b5euqfLwOsSQSA5dK/e+z4GX+oWuTUfDYeKIf0rd1coSNn9+VopBG1kPUmHvlgBib9A0dJy1K0He
q+oWTf4hsdJxcWiENDbbKANNK7HHOzWt+QE76/WtXn6QtcarwA41T/WQP0YFNIsI7wZT8rvrDCFr
oP8HkRvu4gGXdcic8S2G8kEkuQ0MqsZfABZ65ZRUUfVnBjvjvHqgpuf8JtfTmTYbtcqqDg2MsFJJ
T/OYjwWREVMrfbXsFdNM1C1/Jv3ef1WhNycLeivH6d33EbB/DIOLldr9R8oPBDZMi6sNqFuJeFRd
ufXkNjS3C/5ofcVmtzjwAd5mO6Fh/ORSh/33NLqzQJ6wUgxTba3XIc9u1tvKFP3BMc14xBYjhPTp
Dd8X2vTQpLrBaVNDW99aip+rpL9cXFqrw2/tOReGuuz+JVtP9YQlTwA8Ddju1MVrnukFCZ39K9G2
klYfPSS6ozKHZ/j3vfFjq4krxE3Q6HCQ3lBZk/7f9DO6uu3Q3AaF/zbIGcVC/Yt3ymMjkJmKNfWw
FjQzLquxnjqX8G2v37hxTKaYu2h25ciU4VLRtAajYlF4rBpqkWr4RQdvdw5JRrYRO4wL+FKJlNUS
LvwJ4fo8LafupK6ftCksNCI4hSRetllMRyjEE9bwEBnUv+pauNbsCSlxhD/cO+rHjkurZDshePeE
1rH3mTuLkQuXR8GS7HCFMtCPkEVs4YFAkhJMW+VN0d4qyv/d+Aj/XpzlsnMtSmzOzCW90S+RUQOU
8dsdq6+gxciuF3DbroE93MyEtVZfy+opmKgE5ZFs6YYwnbHQQh7cyNmUxS2c6Isw3ZmcqWPIKy6h
h2BWdx4lZvI8w175tt2xgbtSooQ5OHfGiUKroKCV9FlBHZcI+BC+lAPof7hHMTPINjl2R0TX9uiM
i8tQLVZQvT42Kmck/a9CtKSdPkfZPKB2sqdrdCBXn9mbmxOOA9rd/Zodl3vg9XhauE7oD7cDXPTb
NEpiFATkis55Ipz+Y/a2N7mjjjNNlfqa8GU9gzDbE7ra3FeU2EWTF51Wv3/3Z1mNBcHdCky/KP4W
TH4n9oWB7gj2e46uUYeKG6B70ZTgU+2+5u6Cssng5h0Tt14u9RYM4Kr9LcLhRhtzOnPtiI4w41Xl
DToGadXRr26R/kcFYfr6vdgPxfWegMeoA6shyjAGsQAUOJq9eRLFRz57P9Nonwp00u0OTVs+svaM
MeDlDXchL52pAnmbMqGwFs+Ot7bUG0skkGe4n3V4qoavm60Hm6IhVuPTn/0TjmwyG7kM/atDuM/g
4VllH0dgcVWKpIb95NizDhYtDYBunFIyWOlxhBvJpdGE5ESUTf6pUhjnsE4Q6cOXSGP+YS+cHb4i
vdqy28wk8NY9Iyg4KDq3PatD4mlN2+tM7oz7voSFHPWP89CNR3kAd9nv8wgpPD1QOkmnzH0Ht4ZV
4oFgYMDvY3iUtx1qZ6O5qj8QElOF6a5WMIwuYFhJ6wKJ85pLQql72+TX0/FWP77a1D8+MaMwFGCK
t60Hb0V3SoGKmBEAmG2yxiZ9LRc/GmxGC15GPK7KUjOO4F5j0e3BchphZwLTNZg6bcuma5K2Vlwq
aVwFNyS0WN9KIt8UBYoH84rPWK0he/X2UN+YjgPD/45ZNI+MvGs4gZr+wtnsSlmE5vAcx4LErBVD
117deGMLBH0PmDnX5hBk29rPpPe6WOoUxsi5HzOfi3X97IgAalfJtkTm3PRAidVGG8eGmIq16t8z
yVATUD3wtn5Uku3UM8qud7AfL8mVcPA858Vt3lAuhwFSN+9hjoJ2gnCx10TXvzQ6pyuwm6Voubiy
LCg4hdvXm4wj84ornSKb5bikwT0Cbo2kZvQv0MkzQI6rRFDI13r+Ulv9WGxdxvihQpCi9XoscDat
f8EIVo+jLmsbl3OyBXxleQY3ZKs+AL0Te2dNcQykBfgMs4lPKgsSxVjv/gaQwpq4X3OHu7CLHBkJ
+gZyvSpFa0HVWL+feqS+l1VtsG3oarMUbTMNmtMkBA6+iRM6qHDGjMyd170XdwaxPrNp64UtwOmf
194X74UtxehhmY6C61r+9VM/ay8yIguMsNcF47UAEFd5ODNGy0fJgOmGryR4RxmONOY9R0j4oRt3
w6Mo01Q4nqsdbipVKZ+CGWWZzSNuCIjmJeMCx3jbXJqXoStO96tbMfateAmr7mqwzh5zYIxnivTL
/G/toi6EW/nTGJw0VrEWetz72Me0bW4p8c3hZUFNomgqPiqlLMkueCuds8xKT2owMd+FMRpF6xNe
cVbychnGHUujQsjPJov3yPelA3d1jkdiFZ6TE+jH/yDlokZGWivcBK6Wf12JvCovpelEpS65mWMx
I2n/PJezC4eeWr9WkIJjBM2RD+faxePeVAWgtIx06sR51H1xjqufNbTqqIPtFsYieZpxtMQKCQWQ
TEUltV3G107FJrJ8fcrVHKWQ1AYeYFxbQAkWbuwCF7rtr1cKEvqD5o2E4FJ686fgdoDgyAYVjh53
l4vrUBitd22YsHP1BtraYCP8Od4rH+MX5yQQCWXNLn9h+133CUV05TgR/hkkIyYAmJZwNNPHVOuf
p/mazQa5+bO617qL+Au1GlJXKjW6mg8U1GBy5pJV7TdjPjQ7bbyrRJn6pED5HGgndYut7RwVlNx0
K6vcS7UgVgkUZQwy+mPwovJ8d/91DgOrPLSSSN4SsuZC6ejSvZE8CIBZJWF8oO7OO9y5lttHyW5R
EndDN6G3/Swf3wc4yLDIdWOuK1AQpYnNwfRvoTbRtuQKgp9ChY3LbqPA9ibrlA8uBTRwyxgq1YHa
PGRLG+X+SHcsba2AuZpf181dtr04n2wfgqnO/pk2d7b4YZB+gf1Fy8CBPIStN5/eHsloFM83MuPd
N5JRQSB+HuhG37MuzG2bfh2qHl4g79vC8QF3p6L4GZSrzTHZziGl3MRTvv+Thp0digY1oi5V7uaL
+a5lFC+0AM+AYnd6HRV2gEfQ94R1CsTowACO0LJR+QUaRXshHVPoN6Ls1vMi+td829D9Bgk4EU56
p/P1tS/dEHJqOxiOwvNAzIpgpUgpRUi7Q1sTEu68y0wgyPODlTaSU64Wuli8uixoOMKX4yG5GDmY
N7+hAVg8ZZ8x1OzrO3gfy9oYbaQP54k3epxuJetCUz7Yd1lLfk/P89WIwiMZDDnKc7GGVNHFRxM4
9qiDbw7+/uqg+zeIA0UNX6lOZIePcDQiImQT4qXvMZclZXfGJFwSWFY3JmEZK8rfQyC3TITpMfdv
br+B8iOdkfIZ9S1EzT2TV/BoVaOamBsywBov8NY4tq41Yw6q1hGSLtAlPIcEIDqo4P3D2VYPG76r
8gGdjo/I6ugt01IurzQMAc/IbmeODnHaJIWMoq5VHv2nfyi9Wl2cnIdByi9bdhd/7oy2gWJoz95C
89oEfb3sEsBpn6Gt3JeVjoOJ18NP/RgLfJfwihpjABXJ2HYdXtZtwxrBiSGf6GXGjFd7IZrCvG+8
14utcDQpEqrT3U7bOZsRTkVWCxSHTACrDA6W3ZsqHOvCsTG+poRUrhdRDE9FzPKi4dxrQec3XSmQ
bJlJ/P9GuLuyz3z6S84RpkORNxDOgzvmr1WLBJdkcdbEhflxvOeE50k4z+SBKSh6WhI4XRrd3mNP
yQ1PFmBWVFNbFipKRvhFNHtnAuyoAyWg6tsRhNbjYRZsBh3xmioeVioEdLp/im1APszhfxbW6Ye3
hqz1jT/9NhU2bouS8eUB/aYHkxa9WU/PIS6g7aheAPMpnbmkrwosKkL0eymVYKpoged6JMXTLwdK
puSDqYql/x6lEPN8yEsDTprlv3hVvC3oFdSfxNkkdLyFq5NvfT5zQrKgIKZ8YLd5mCYT0rcNdklq
BKdRYdDLu9adfLI7cWKm8egEi2Sz2ZD4elNbFJMpElHPcSCeBQGsI1Y/glb3MG/sDC9SinFKtYMo
Vh7k+BDMnbKS2T/+UvK/ngaKDYcavp9ej+LtH4hir8vFmfNI8n8XZEVqVTM9hAjbDjIeTn89/309
GVBNOvaa524f0kERoYZLRi1GNeAHjjzvVUAfDJAFp/U3q49R+Tsc+uH6Ym/MqaNzQDoNhjQyepnb
qFypVejl9mhi2GK1gIZ0roIteh++rXqDkfWOw3eWzo+IQ0cBKiypQs4Ez/3JtmewGkeHwwKxN4Xa
XGDyu/crGbdhfa8fap/STx13iKVUYcRt7BTwl9Y4nxRgkWuBsbUnynMMQr/miwWQ5K6jC+Ywmqz7
/c4F94x4N72mJFIDJQ/g/urreKQ7E8STqIl+9d9suITrobn/8WYIuFcz/oJhAmT8Kmbj1G4ChgMl
/PhZ2V13+njcLjvKhjfS4UvZ3gORBj7In59aUzFH0W04VWFQHdRQfuRNZyhgG2wNJ3efUZo7udBx
7ZRykWyyDZdZsbHii7jMQUwsgqN9LzAF3IrvCVg7vSfUbpUzAhESGjd1NLbMfdQygpSa84ojC9bK
+EsqWgVoHlGb/JoFPZ2qPl2dQJz1S9Zc3zaeDwuE8/GwkFyLpa5dJJKWDpenMaoAId5IS0knWuMm
JBE1lcQ1LTrACh8rRDXIeLr3SfSzPD7LuQLzw+I6AVQVgtRlKlAItOsb+4aNbqAkKylyQFUjnbbw
njnNb1yoWT+ENWyGAk7kTVorbT8+ltWJZWBtD423lkpWzw03e/TKWfRwu0qm8Sb7HZQ4FxwvKFGk
+Jd7F/UjmM+Xr7UnH3C/T34gliqXD0t9JtTxHhasZmhBDBn+bBgGkoDDtxxn+AfSC2tYIBZiKVa/
CNdC3H5Nt9C0Hsw+8Gb5eNz8BnvEtntLxk5qQjlDKhhuMNs3MJ1+XnbOowCq+SYYfkviNpUpOEnY
WJ9QsM31ruvbl/a3Os/mN0hGqOJCCvlBzhEcqLOF7YwYZsu44FiGJkjhYNdO2F5HMmliE72ddxTb
uf+WyFZyKPCSULBgk3/JgDtafiNsF8tasId6+LwU33zZrGMoXYRzBKrwdCjxiB37NsbJcutDaYvX
WU3eCRDDIXEBuEwNiJ4b3ObUNiAR1WrvNcex0uXPQXg1rhR9HuvKC/uI5X15MLFIV8d5Q3f9+8yn
sZmOd0NWaNNZemdx2+Ba0rKq+cd6oHmco/tYpIhVgoUJxYwNn271RM6sCr86tkm/T1R7BDyTjjVW
mMcrp8CZe1n5fqoFMVr9ZswFUCXki6jpKLFwFeQ2fcpQuiGI5JmDP+YrvmbqJiqlSbUFeESen7jz
kaGmp0QAaLssvNaMUr9c1P9ZzHEfC9obEnZo7o86h/oT4lZ5d/232YBnUDzSBY3Ctij3us40gKlb
qtfv7YEaOz93ZMJqVv4i2ZSR+JeewCzh/WoaGl4gzLAnaE/Mli/4vQt2dAnK1Yl/SUQ4lNOOObAf
cw6+xMASEiaek4cUdVpwctUy9oKMe55Oaf2wMsqc852FAyQFLuGWsspZ94XhvyTfxVplizhYf+QT
+ni4CHgp6uhD9qrslyLANw5Zk2yiCf2h+p2j5YA7MRghuWb+yfzO8wkzm9FYjMXgHKr8AbCca75N
EUIIBk+f2BqYj/bCBW1I9TblMtpjO8LetuzmsxdXK++c0mZMcma7iU5O1MqzU1noJNdCVcVKeHzE
RbviJ51vtkQhvSJEJi4QXNOTSKuuzHy4GqPnGOxNTMnhSMb3hPavENRdUIpTpInvBqByvoydvC3t
XhUvhHcM1F72eqz0dbbSDzgDOR3k2IpHpxutB+MFhLT6ZHVUIf0NURqAIHCKW2FZXUcwtrM0sajN
NncZ7koLsrYumFP+u2mNH01UldbAtvNC6ra8d5lcMSYwWwOqGod89luxdebA1TpAiqcJxJfZudME
wiAOXt76EZRROCDh0nMO9HuzVqg1HQmOCwftJxHASkfd4a/qjKrRakxoyCKXFLxXHyFXCNhzTaXF
L3hchELegeHzr9TLzxh/0XvEROUhF1VYCrKqPdZ7t6RSey95Hd24WHQIW1xFbXYSYratob4iFKI8
gTLHW0eg8HbBXT5PTPN+wvxIL+GhG/qkdAim93Tz/ZyfH7lLd1DpRHfi+HDmUi2mUJzGhgEWnTm7
2/W/eS0xiTyOy571o1icht3n3nu2wR4hFt70I2dR9HLZrEhx7XvsVeYB9YRcYLUA29pXP8Pr4pO2
gzUJxMR0vCuEYFZQrwimCUNs/x+UtGoWqFLRvKuPSou/4MGGgtOMGRo9hpYY0c5GMfJMbtmhSej/
O5eyAjt6G2fHGtJG5UA36C006lQX35R51+22y3khQ04Mf2YMn8Zh6XHDmX98VkoU55VRZ8epudx7
Un2YlJOufYaTxsdgUug4Kjt+3FHczIRYr6THsv4Cfn3+HT9ItvzT8Iq9GTpnIMEL6YX93zxzFn0S
7sjf8bVFQavhAAVyIMJudnm+F3XZ2olpq/kji0RyKgVyWI0ekN7YpZmxq+TX0e4ZmHVU9vdX1hO+
jjGPoAMuaP8HlaqJh3T8OXEfPJBWzm6b0+aHtnwEUMS8y/+EACfkBV0x2nxLgpNNhwW08WwONvaD
Ge9ust2EiuI7o1n3W3xyzj1XAfota2V16y2izz+/BNEPisrHoHg5pinxKilQDyvRvXMOwMtwfNB3
VwdBq2+KcAA91cEs+wUb+zH8RsiFJ9MOTUUC65yLxHLIk7ruMswlG+EuoqM7UgXv2FApz1zSUjcv
5B7Df9EOtiDOl4VPl5uEtDEACruMUEJCveaBg7Dzo87mGpmNCnkgBQvroOGLNN/15qldGlAp/qQW
ZV7QOaUWzO4fahcYXSEhoSeolR1kb3KmtutRl6J+zcslqzjrZ2HcVHZmebVIiUp7+Dy5lb70Z2Ga
LXuJ6PdKj2dfim50qsVedPHrn7iM+lWXDm1PWylV0wneW6op6WPIskdWRgfnuPGidodDNRnqQQas
mXVf6tM1cNCNn+zN52uTIchIkkrV/TjJpoZnc4nkb0wuuOtj6tUX3RIK5TCM8IFcAPJcVFLgg2E5
vcf6b8CEylTHAVnWLWRIyjWq3r2NgFR+bj7isuAugnhqGx8jzoaTATBoVtTPew4V/mvgRyD6O7Wa
9xX7R1+8azecfijBoAg9sw3OuU8kDjdsSbpddkgmrQNbsa16uX7AJW4fhQA8GCk8165Kt959QrEO
+v17ue/TqhRdz27jn7dz4TBwwlFDgbp6prvQURkYe3esqcFKF3cDElVKtu97YUVOc3yAKp25f0W4
s/Im00vla7Y+gtX1bRieNNYBnBGZb/T95ePS9NNfGJgmQiTehFHOHUJBBPBcBec0mC6ESFU8yEh4
9ucMyExv9exPrNu2T3eiRlZfCY+dOLw88nI0s8WMc8GmQUT/tQGxb23AilprIWyyU/hg2TJZ0u28
oOBHH08+LuLlX3mDPjXlDgYLKgzY/IRflXRQ6ThlnHEfL8v52O1vnyX3fgR88Lyfwv8ip+cvumjS
g79yvR5CQiwpLrIeFMKxlRS9DhMmxuedZApVzlmhQLrfggIaBScmluSExeJalm1tIBPAsI/GxIVi
W6f9yN0hCUO+9H8Agtsm9gnTrU5J+bmvmfN5GwIkMmIBUNZmA+ZaYWxHGZkkDdl8sXR5zefyRj4S
eKzAvCczLXjuWd3amp/i5ARIKmu7axT2QFwB52D4/4xiZaq9uPrcokY6gH/N4mvzBX3y884Z9ClA
Q19SU46WwsuBxVhlir/lGIidxpcBMWXMviO/JdGJYGsWQh1mW5MjumYJ4IkYdvqHKWE44qp7akOJ
uK2XWtkRWc8IrxUGA886rqIj5SKdrXdhgFM7WRysQ59o4qjvtQBJDYwSULqGDNA0q4KXaIugCv0a
4HnxG0WNTjSTAdF5GTi+gFjccrQILdWkA5EW+iiqPYKv4RpyOswc6LnkLL2Zvi+ZW5cIHp3RtyZa
//9v5Sp9UlTehxl0TR9rvXqFgW6qR+XpwhT/QlNx8P/k/8ZHzWf5WOPJXCkKcblm+GeG9fg/fbkL
dI3v9i13m36TuS2n9/QiJwxrsq15LLMlAodY8sYfWoUw9IzzL4CBHreM9jRClVgQW9ClqchhaqO7
weIKUsi7qOYEh/iSLDTPHzb+l9+vqzPSmj1FnIe9DR4OagnksvgdQZzD9zXxGnketu71fOlY8HUS
tvn1oJtlL5VH4ajF51AwjDukKzIhavB56YZOF3TCDsutrw3jlFDXDVYVYFsJ0gqppCgQAQbz8+Se
CmEn16KrIsIrKlFViB2OskvThOQY6Y7g10yQAQpRy6jAQ4UYEXbZQ2YwKkTMdkstn97z5SpeP14F
PwEXosVDEeR2p8DhFVUGZeGcBuH8sc93leiKvULit0JVaWV87XSz8F1yrtrYGP0XevH0MlS8R7kx
8lWu6ZoQX6aBWYJIHkUiA7vdye66/zhDylZI5nj4S9hjaXwgAoA9tPjLV5aPnQ8XIwzPEOtGMmC4
MbTOJ3r0v7KAGe2l6hbHtswoNjans1WoJYYUIYfAWKzes/EJiFd0TuHcIPM7Gih2h+x7otu4v1lC
roY+oVtr2olEDu8krKHncp1eIrtBlUewkeq+vlSvWVSPfwNeSPmvY9dmbOJ+b2EqyxD4HnvW+nXD
vacOj1aldlC4FtGPlkkNnPTUVw3wLiulDt3hThwpt4xpVJRp0Ci41/re9ohHdOAAc0IjZSfVAIKR
EHsJ9rzGPygahRBPYvxjHi2vZLNJ2xx+w6KJvVERJQnKUFqn6QR57n2nTGq/46jRGYFEY7uq0aPx
YT7sQncF8OvbXnOC+oANJ49AlgsNWn9wTpSvc2e0PBGVRdvJZnfgVCWqI8ag2md6BZR9wBrP+qZa
glIodnFyvvsOwJ64pQODtFFTAy/B5XN4OgKedpqkR77IidZB8UoT9wYP/4q7vjMZUmyjMQsG1ISY
IWDDG+n6KYCSdaj3+G0/h9f1ADAj7M/RMi//FKuFsULjve8+2HZYIlFOCsGaGBzaxnpI2rMv4EEj
iSFVeEASjEqeNTN7Bd4L1XBw+PvAB9ewhwtIwrzY5Hakj5tprTgz845tMutWDMnSZgoRV0/1Wlm5
cDxe5KFfu2ZsifXs+N18Um7H7d7cG3ljekDSs9SEguN81t/0bQcmykzp/ZHty08aiv2g6LQ1rZkf
6jvv5hhH9MKaIobKGEYq1EyOmemJJsvAnsA6Cgh+fEqOmiujDrD2N+FMAQYOOn4X/EZhtkRIDodm
wnFnKkSZEyrk+DdlrmcfzE7xkv2OP53wJ4hLxgbY7SVqhVNmGhQ3GYOHf9Cfhg2e4kqpLjDoDlhy
SQ49o0rzuqML/1xReywNwRqy+xguYNcQZb8dabF1Qgb8xrBhYagj/Z56lV9ZfB7JkG5hP04tr4Xs
r8bM3phSW8gY5IxyqQpmGDg6Eu7/puRoyr7HAtgNHZCQQvgkUSb+WH0ONJ5C+rOtfaPE66SZiPmx
JPzvyGsl6hGQYCba6dr+i0z/DpLSTGFl1xuUXmkmZPuuu8YnFADzpQIuaqf0d+xDz7RSETAy+Q4E
bD1CJOkNsMgfdOIut3pVRWMY4pMuRDqAGlMJRWQV43htcgu4B3pcf5017EgFqVpoUgZB3dMIEB7U
TMKWwRmRgYD09nGRSFGFtVNy4DgrGDRpOcvc3acfnRJrdR6zsd4YCtNx5nKXkUwnEjM1Ttd/Gm6b
9Iu1RSdoC+oeHrOE8soOvyQ00DMmrPw2O7yKlrZuUdTuVl8orsYI0Ej8WlLqwZQNw75c/SM/fWR5
aqaNXZA8ZponDw2qg6SXeME09xkOl9YqJ5rN9eHF4Wli6mctns2R/4GtFC+Zwz3xTtqgSWoaMbmF
UuSymmxDe/RPL3fWg2hOp84hC2Yicr15a9palcuV13gEbXZVjg++JFrliJUs0QvjheZzJqXnikH2
CySkXf91IGo69xnI861nXBfNnTaA7E0kqxQ+EpNz/OEWcfaYK2R0jiwV6iYNgCfSosfnUlBSuKIZ
vRmttYdDtzd5rSP6FNYAFCu9C+O1DVlODCmR8S+gYde7Ss7k32E/5GauHWo5eFi+NbZ5KzDpYBoP
WlJgH3vqkdRoU3ZNNDYFG3SZYEGeU9WesfOGrvPzNorgIGLdo0jKSQlpZGcT2VqOOX/uf6tZkCyW
NRjpnlHYy9c8PO/XmPoPJh36DECBKPBKhJQxt4XOourZLF0oQGoRLCQmuRhSnVMqENKuVUKbOeIo
TfC62x/sKajO7JKzQjr7svBgQbQ+pemzXHBRqLAjVOL8Gz8+sTOkSMfjqojUTIW2cLrvl1juv/1j
3bYxpa6KJARg8zMroUVz6Hg0vEMPbN9g+JWa3r/7VOC73w4h128vEl0W4QoYxStshFGCQD/DSAoA
Wzv/VSdYsWTRBabTlSB/ztQS8CmgZSWfoSklB1oNO/MTHCBf9M9IJFO2iBm7xX+a6P78OZjLJyec
rdiyD+VqB3f3d71XpgZpAm0xBspRg4YgI1O65BPIkhIkg9OEAOmaXfNFW4+SdqXbelpogRkw7S4p
Qr9epGW7/cqjTKLHY+RMFG04VKPVT8bifemBdavJ5A22SsLVF2f5JOGLyaI9smZMm5FwPAIIJxjh
Bpam0iGVMdxg35NT94Nl3c1OGnNED6wrGwWnHnqR8cHWiJ7vrWRCyDdVZCONcauxmaP5sqROhZxm
RsjRzzXDUQ00TwGatR6Y0kyx5mynhfo9Ew0PSO3hsBg0kH4IwTv92yinPTRClbYl5zYLrX2wgbea
O93HcPL9Etr10KB2AN6VIvuJ2nxP8nbXrKjDyUA15M/UEPWJEunzcoJ0EPwhdYKxnzM22rmqkmHM
GiOZPK+KO7v9qV79SRombL6Ju/KPxMjqpnS0PF4yjBbmQCwRTL9uRhMAfx7M9C9Ps7y2jWJLdEhO
NCezqDol4p6/qxADmMmyE0cjQwf3Hf/cJssnju3k6NXFPkycIPhW9123dOVUW56UV1aVlsVjwTfm
4PRaVwG1xdV53Bnbr+7fCiUTo6Gn9ZBOFlRhJXL9pL1DLPgtVbyZMbxtfZcUzQ3VDDfcWsgfhqti
/26fV3q1iJDDhG2uN5dgU6DU+yIpmgeXXKflg9aUylpCu8wadIXchyEvYm1aDXX7zFqz+TTlub7z
sKvtOIr5+36uWsZuZF6mpqZSw+SxA6Fwvi6QssNdycTF4YJGSJ0vnXidLxq0eX6Ukngs8c50YRyf
FwNCGw3WUcwntl3rbwmoQnPboOBqIMa4enytemB2/31msUPB93pE6P1hJG5kqhGkaaDdGNyBca+N
Q40wjLrExi5E6xU+L9kvOdAlWl7MNzv1H1kb1iAU4gsB+VOV1zLLoXNbdk/xyfHlcSY5WqP3blQc
DBPxEPQYkscvRyQ4JufqtI66Gfdkgv7X2QD7vXl1q9g/OFMDI/EDJSpcCvbkYdAcHmKgrlPHYRfR
+LbHNQrfPxPAHohZpM9mM62Dw2eQrE0rJ/Ai2ffTEppgbLT0+/axbl3abpZf563xAON+YJKNRPI4
7c6fcPNbpLRQS5PQXlOF0t+3uA6vuUb85eXoAgb3ijD9ks6dqCm10X3Aag3G5gsXBPvoKdnYn76Z
S8ai7zQ37y1cDxWk6+qtyYKsvbrzh2c9CmhawPFODzCLZTwS08e6mcFisIi47GvBa7C0EOWPvae5
IzABG9aLYlWuF6c1YjOcbd7FbILBmDdc63m4WmeWZkyaEDQN5zK5l02MzKOBM/fgnKeV39iQZSNq
emOsmP7xvkpKPsLqKZHjPHAlyAgV8P+5fZ3xziCWKIT47UnZgUPI9Qlgyee5XYq7qJ0wRNbfHPAy
C5E8Gip8UUUONca5+20WD9fukIPzJmoauOszrM2FuuJuAag/JjePUGL+4rx2g8MMF9Rxlv+crWq4
9CRdx/Phvhrs9qe0i7n/gUjVyhhYUmsw6W1u2L1O1GLta0QAuQMcuQVCPJY9TQrFpeWcUXZQVu+w
75ypFj3j1LiCsI1TQw5fVNRD+zADsam5hOlsO/jjac2vsBLn4ITin9164DOH+UxYbAsR4OPGWS0B
fS04jH5FHeNFVpduNK99ipCXQA7tkz+1aBc8qfUPYrwpDPppZVA/vpQ2QP1xux0z5tUhQoP5EOax
IAG2NObcZCX15qmwvcyPODIEu9VVvK6nBVOANbve8npVdLiQe0nxk6mXuTQcnU4/JuLvdtWE89TR
1te3fPly50Uhc1iyzbgca4BIbaKDBHK4syUvWxo/GdpxlzQf4UzkbKAg6Fi+BDWqs8euggN6yq2G
vaC/tpkMbu9rgNqYnsznvRyoINdHkpCFSNguP+7IZ+05IDB0bGi+Um8Hg4j/XDy7YB4xI70cJFpR
XjJEFv0bU1L0bJHGNNCe6ufjpqVETu4AppDQ36PyFIlbAOQWccWU1873meVNFeeSDjPZcWcFxSpJ
HUIkmpdJdbApcrmlv7cvbeWiVL03yN/o5EP+UoGmlQDgVi7muMpo1QDKbJmb3ogxLiC441KOd3EM
tlKrol7WP/ecZWzJc6CvavRsE2Unq4N9Nq0lnnWuI+V4+JygF2FBO3Wmf7CfK4dBbaRXrjICdjUv
VeAxgvy+/EKOV3uUyIrFOmwIBIQHThONnjzU5HfYJghlkI16vGqvc2j9jUfEUzXmLSufyCA6pLdV
6hBh/UQ4oYvjJLahLtT0Q4e2JcMW6i5eCLMqLQAePcjCZYgntTXT0jImTKJoRumwlIJV9OJ0S5v1
BO0re1fWWe2NwBdxjt7lAzuUCK5UmdAYqFlkZnhlQnXP4kJHqO0c0uAIzeuqTTwSXfjdaYKEkmMG
kobkPaVp9e7b9X2hr09ksRmSHCicS9PpwuorVLa8i0sQpOuU3wzg7/PoxACwPI8Qo3cPgcYNWXU2
AfKTTlEgDv3JxKr7bAtfQnR1CegOIqhwYVY4Q4T3sqIbiyRrd1hcM6WTENLqB8aAAL5choku7YuS
BqwjIqJ49CbGpZDApI9cT/O/3mK3J4gkh0R8BvrRbVsASrXnKWSifEbHfQOGYxuiAfMqLQ+VND+W
1dlkb37KIJ8pAwNdHBJ0gTY7YMw4v+0tV0rvUj2MSRQzFcvGPIMYzj2+fuVb4o8HPtYYsT+Vv5/K
hxUk715xVYpVfVMmc4fkUEQ2AW/Hx5xb/qUn0uTqWyAffZgfY4H6ZDUKSPtcMnIGJkm2qKNd6569
lGVBWypAmf/d+qz+oQylJpzcMsd7dFVUjF/SuZNNpM34uxq4qM9YWVpXpCRDENk5UsMe8ln/dxln
EBWcRFNpdfYTEdmhfLpjCFQDkOWuViuGotplj4o5hhBPSNX3jgsV/Y93Llf6DqngzNudSR7rmmZS
XQ4Vg9QhAAWICzN8EXfWdtebb7RylllxGLPps3FSxcLUOvUgKkEcFq5gL9wH37tB770RZ+l9Nj5w
Kth61M7MP1ZIdJ2HWc3/Iyn/3AAe/VsLx5y4anX4Zif8Nab9jXiMZbm8rWuBHWieKdpGdmhFraBg
1Gg9NS9icKZFt5BEWHsUqIehlALYybG7Hkp9FGn4OQBbnT8nIZ+wA4T09vPSj3M1faY1iK8Pzauy
3ZLOF6dtNNtrlrv9mF5uXgbPDQyypKPSCyHQ59+vfflillhAUOtMgV7PwK0ppfrPJnetDoTuBfys
BjL5/pEnM2YhQ1fb9unEWc4RLjCqgo31MH+e6Dj/e3DWVJAogQyuWQ0YHwLMv3UJV95wELWwVF3L
yPiV3tboFLE3un1232J9SF/07JJJBmskZIFRI6xN7zJvyWqUMwqtNNL58tITeMm1RCpz71LiUHfs
XnItb35umn7p0V8NiP7rOC5uJzwpMeYJQpk0seYihx7zAAY1JBBakkUIqhfw/dZwN/zd9EGyLMOS
r02bsKKwQ3u0e82j80QHCmSqR/a31r2gGHeL5xx85EaIAQI8HqbaXhNTeQJnYhuPUH2dtXOVONLI
UWzHjQnLe0ROKZToJqMUyi4GKD3tACzxIWBp8DEao5O0B447cAUBQrrGiUb42SyffZALmIv0sJ/6
1prozGXgshsBLIl8a+uctgf0LCphORK+2O23OEX1IfEMiVmDLRwINfusYrMCGJUZ1msMf31I6Ca7
nhZQ/vtYTELyRPN9e7RKSXPXpAqcMOGmicF5vAsV96U6iQdOOLIJ5Wl5q14Mzizv7sNv2znWN4PV
bZhlEmnMUfrtqOm77jaU0GEYVoAE1osAXomBaVWAxvFAsvgz2kfsn9wnfp75KN+1iOuliXYDBt/a
TgcrtqOmv58x38yE78fhnaBPumZ4Vbjhdez5Q5WuA0VaQeb/Qbqkdulvqvty1fst7qi6HDiWMf+Y
Veb1PuHBECWEBHE7EL0T0G3EwqA6SwV8z0/Lm9OtmWVxXZCUHNuUHrx4RPx4Q0oH6H8Lr9eVz79N
iaxEb6JBkwgxabGR8hABwaWm+k6Amt1WZ3E/IgQQouhLwxPRt4Or7LMmacqNUBw6p/6uAS4I6KWL
AfCvbLXfIsWqoFwJLHmdS3VbRfJSLNvpF5gVwbyY12u5+U03rYM+2BTRo/1LnIdIQriHQ1sdA58t
OA6DMjAg7b1Xv4GMTHRxMDzPkHEqRK6sKR5+s3rp4gsnYegHMD+BNAIEWIKZbcNiREJXCBvITJzJ
R1zlSDHcaR8GLklaHC6+ehSOMEusDelXXAGsy7i+Cf4d6rfnPSlL7UvFZMjRQ4I4qHX2wxuSkcgD
ttMKkr0eVIOBexmg0Nmtss1NI8niW2Bsuabhvyf7iy5QOlD+Rc2OukhP+KrgLNLXY5mO3XeENuOT
oEoK56lcmW/9xvEbDSR8eVQK9mtFrUubUo0S3ATgI6Hx3mdw9NXFhHoyL3U5oySLGRzraZ4cleHf
KDq78AAitKeOpIryWnmcoYR95rjVWck2k/IHQappwEsCiQC/L15EE0sFwe1COB1R6++NTgzH/hIO
750kXIIpAJGoO5pjkcYPJGAKKS8eYl8UOEdmFXUQqpkIt76Fa+CiQB/sUhKJVGrgYXXPNgFLewuF
Da1QvFXEh29Nc/+vF7K5osKEW0Hcv/0JtTtXVzca4iJKIEba6UShLNTUCPxTpYDLD/hmWc7qv6a7
X0nIMrZzNCxRUed0SDXhN+ARqRLh18pVcxTBpedhVtZlH9c0kr90KXmFaQj2mZ2vXwdx8gH+Ka4J
5HI13L24in/iH7ywX90dy5Ehv2RCpC43VnIiNwF8s+U3ElsHyHdjf0tDf0U360mq0tsn416hVcK/
R0Xa+gYmTuROk7skH/K5IDOU1D/EjHHmWCnUQ7dxPzHWfz8e8lVz/7Pf41QRjxE20vyvILggtgr3
4Hb5NuU0wMBbjImtDmNfrt/tBwvFoZCenU+iYxQyREDqLm/habYf4cSi0HJhcKtcKMEsclqpiEuF
6IA+y45Ix3Juoi2MmgOzGeM/G3O2uNV0ACUj8DITWv2w7Tau+4RF+vwmpIKc8YUUI1vvZ856KOYJ
kOKu5BZHUT7PbgQujJx4U9cyPB8+WXSuJuHZpBuKGJAjSHjQijG/JYZifkZpgT/KF2AAVmqgxpRj
Nap+pmGgGiASt3vZaAc+kzN53asbX1roGBRXS4piadcmtUGeSb9Fz3//mcF3sTOxBUQ7xjh7Cp7o
QnY49rzOHoOFOjv/TjggoFqbIZ6gN54rWL5I8Mp0FHk23e2PK8feUxWzQFeoXhU21OLAptl7P83e
CsNifM/QOeoiEW5g1ck3d4SRe9ZtQscvmfFtbTIosVgOq+LL4j6bHqMlu4MzhknXvHZDazxo7fTk
hoxbbEfqx9kIlw+CzVZOgP11eJgs7A8dkxSYkU7OynDZpatCAmCF0SugAqJd/kUbYbD+fwUxpVGM
EHdroYwd54s0xeKYBkL7xFXwgCwagQNm5jJU57DM5a28lSSZzaRAFk8MzqIcG95wJG1kXFwoyjv5
QZJAb834D/F8st9pJ3g9wC2UQ6pHmw4zbq89u/+QBc5mU6gL8NkaJbjKOZ+UApIS52IlBbzv8x7p
j+mtCbMPvmBfH7LWoIB90aM1VmR58/A6GDR8OhxfJIVgc5eR+LTJS+3yQY6DrnWQ9lEyJ1mcYa2A
RGUDIeK6bYzTZUHhPo153Vi5Ti2P7QyAg2IHGna27pmWotYCXCrW7D2e3ePO8ZxDhsAr8GHXVLn5
TKngcCVi8zay2rWO1mZrlhlfokUXTVydVNb3qPHHRnx6oelmyo0mOAQXMWSoT9H36E9WqVM4SH9g
SAs2WK4AUUb7RvSP+PzNGrZf6+zJcj/QWRG2U6LCcDA0M28Uf67zWthJAxNxLo4kyeGGeAGa+7ro
hnhjwL5gxT45O7KT4nP1MH7D/fB8zgl2FD4tYFPT5MWZbbAN/WVtFOxKK1iEYUIzsn0HR4OuX2+S
kViiF9mdaSFAl+04rzVql00Nbxs/nTrmD5Lfr+84gR5eZeklWchYqVIIqE/mN+IWVk2gkQBrtjzP
JIaAoPqHIZC0MQSq37J06M/1EUfS14m32L+girEPNJAqd0CjdLns09h9AcXBeufa8FbMLcXPsWCh
cL6g+Bd/MxJDOqCvMAIvTx7Y3U4ACBdlVQ0IJaXZU0RWAtiVh6GUYGrAuUe0b20FvRWFKN7ABm4z
w5qNpyHqinlZPcp3sJ+Dy0C93EZVIUMvWVkmlupci1XW04qkr8mng9EjchzyzVWvDT2im8i0kZbZ
Fwrkoly4XBRRv6uqLvJEyJW741zrxYKtNw4FfMjZQMky3OohTkWIiMhWX4oCOE1xU/s7RCjiG9Fk
EGXUkSnM2rcFxPRndcPnzNRLS0Ge2CDE3CgM2mR0BYmgKPWZ0L3nh9Xf6iwm52GNtdeNyqk4dxME
hzbXDZO2YUh9faS91Mbi+lLhZ7lIVLXGq4CkYt2Rvx0jSPLOCdagaFCyUjyd2mZm9U2QUrXV/GA1
7ii3Ct1LgInwDyj+2t+cP5nmJdO31uZozNP8+wEz07pDA4nUVxAaLodpYmGgyvxMWvS44tcklcrE
Lxzi9ZVE7z40hu2pF5Bod0qzM05mTyUz3Tgeyfubm0inEGda5Bf9AczYSPun7l/dR+pbp7nR4871
y8QnFcEkzneI8akYpDoFLjqwfStuEqFCqIi2/yQNagIiPfJ2wndMOJRupKZpFAjqx/TC0/ToZjfO
0qOo8mRK3ncLmf1EKhrrD4gRVFgdbqpAOtjdvtpSCp+m07dRIk8hYFL/6YtGXKHc+JdmjORH72d5
WFaijSK9at3+0+DyFQJnlB5T848xI25PGCVBPGZICY9Vfaj5t9TyFqmGz3yM6YNQYC1eubeFddE+
HYzU4CkMwSA0szIrL3cBJurK/KObp7z/OoAPcf2ishTPyzJL9p8er88PJpgkOrjBKGDazMLP+ySm
MbO7o8Y+Xl0QoVzRv/v8EmSnF+6/henVx3NUfQ+E0nHNEH07YYG7PB0Rq/xN2f/KtfZcvW7ZOQPU
Jt4XzQJVG/7R+xTZtX08Qay7Dcf13535W4PGFbMMexa+2jdqSXInsKI0lUwOvT76k4f/RaSnUVyo
cC+EI7csHmd0VsDe5AwCY1SQazO8QfVZKQSz+cCfKf49Vrxa6L6xmeIrly9KYkoE2AXEmR8xCg/d
J//anZ4iqAF3mB1qZE9DGh7rUGUEnjN8KjSyq6Fit8TXMGQrrNCPE+kOS8NZazqaF52My8NJl7xg
0demwtOCprphDgJI5TfDl1SqU5rDmdJgy/US+UTnZUe7vTtAVGTRpnjGPtovnCklyZBBp/FiUeze
Do1Aclk+TwD8Go5cw9pV5bdtgXBWFqt83kBz3nhtNB8HsW17M4EAv0gk2ziHpTkJj/KLRqLuW4cn
WfYREGBlmVzjbWCV+J2vWMazTOsUNuFzuPRjG0q6ZnSVV4w3zwTBCcIoLvM2cvCA4qdCLe2zIYQ5
XFwHlPkz49n6vrCA4MICKq8tkY6q+nz+tlfzkwVZG0EFWh6dGcRquljMt2csUihE50zQX3M7lC1l
PUaqZuyOxcdsOCAy/Be/SscEcZ6pNSENcvW062yArqrxrhwa3reiFuCB+HOSHms5+zZIjkJVlScW
7jtFxZuz6Gv9KEZSdqt5L+s4yrsG5bxdO5WgZiecwsOzFnbTPioF9XfgFqbUs/03yDtyvUxqE1Yx
iuYRBkME1VrxILKEDtbdT6mvZu2oFmRHnTYNNYlUFR61i2RV0epuoRUMYZ7yKlFG3w056mxmVnDY
v90mArkWZAAKDYxzMraax3BDrU8LbSUQH69ju4HVm4C04bR7jRmmqyGszAYpLsUQOGxhADrEFrlf
/6uJhmEWh/XexWVvRD5WnRBLW+TJpkSVWCsq97n8UoZ8EEyPcpv4cuyUMiuN4FXRUrIW00gwmZvH
YGOV8X5TClzTIQsLt5nJ8uIyxWvhNKWt4ESIfYJMecCtsVqOTD0Gq/5UlPvbHFBLgAAbGMQ1bjDZ
teXRx1pPC8OM1CcX1vB/44scuVsFnhmJsrjFNUNI68skWlGHNKinM5WWSwtYYJ1ffuq2faA8OB1j
gOIckvbb0dRX74jKR0OSNLltg4otUrNMWjEgn+fHZFjpkduYMknkRya9LK69gMfp/jtkpr7/R61p
MZOgOf8a272UrC7sJbHtiEpNeqUai31qsg50fiwkXo1ySLYf4Nt09yhPs5rfRU4hgKdzEw53Ml5E
PAODt+K3WCfwpinqwnYSLeU3ZbzzeuxBZYkwnum2cnk073pO84IwSJTR/UuatIPi7Ogi6tAqI8Nr
JlqW32LaJkM6kVPwvTurh5tkjF+cKBgrATjDXSyDnDWqZWONDdySUU9h8Y69Gri4M74zdwuABqFQ
qDI0trLpC4HP8nV3vytUoDPyWggNMB1y5649BKasVOaiBAuamlGPCm5LXVhXMmRQIjPbrmj3sReO
fQwEnK8/XOOC4UfFVmbDgxYhHxrbexLE1hkd//B1BOX01LZ9vIjL3gCfze0t8d75H6EJQVv9WtkH
kD7kvGeWIbhVZzTj9U9bfu/k7OC8LY5T7B6vxjCEkuhsRWfkOyGkgTIVoEOLq/PhKbNWOYkTyX5N
z/fdS42OUcGNn6PMGNfNPHKPNykbbqiJFLiOjqD6+VXXWT3gpgB6MWYrM0rxTQNp8TdZlVuRx7t+
TcpKpI3qzZP2fBWuLFjbxZjZ1b2Ijvpwg37UZSDIZlA9a/RGOjgSImZZGSp5fuTiUG89NhcgDQ1c
tvAWazjuFmx2roCPg+VRFmTXpudHi9CbsqO9hkscWFgK3kqaNkun1os6foX1Rt052+IL3THh0nNV
Dgp+CqpPyJcXu+JHJAGEUWJWLDduO8VXyr04Ya7KhoDtH4iAS+OF0KBZlT2+slhLne8cLiyOTePh
T6rnrrZ/U9e/zJe6cjKnEP9sHUVtBbzbNdFsRYoR0kj+1pxHlJm5cj0+Q6mltuTtmWpLm+mmdO8y
Y/TN2zzo5Ilr782pwnrFT0G1bqDM5CnoJEsz7Bt3t2nuY/WOaBC6QBAAQZuti1QSGuhUa4gO//fV
dn3H4pb1yLQnq/A+FDX3w+i9GT3AzFOAr2Ewg7oEWYBmfuN/k7M/FbnPElU0qE9/qBhJHKtNAgws
zteVKBUdI76x0v4NBeCx2y9j8CJYuYdnkX/s15KP5Tgvp3OP3JYGM96iCXyXg/5ajAj3mLw8duh0
ET+fYWwwLLBWgd7YzRxApfC7IIWfZdPin49aWmXJp6YlTxHFXR6FITfuq+P/jE08hSsmfZYYKh/Q
G7ZD6DYAR4kSL8c1B+YpCG2sWdig2WhXtdjhgMsL4vjAsq0IEtgRk+ApyFK1HGIp4ixuYm59+ajO
PB6JphWvZTyPGWFZAXNk7SN87ohsYVRTdUoSNqHd9v6wfQivXPk/5HYy++w+CpmGCRYe2FFTT4O7
Td7H8Smi8u7Msh3x0xeX0XVy+2OGVyK3ENgYWKqekh3hyYyfH4StW9HKp0ev5DOQGeR2/VaBK3Bq
qrFV5MUCJ6Rvo+67y7Bi1//oJeSsakw7BjYHXkAx3+y7WnLb/hz0g96OSih9rMTtp4wx0EW+vnvX
23XzA0Z2iYnm/wajd20vL3f28el+N3yWQKqF8IPEJTA52rmlEtFj1Ffv5dsPs1aiLjmYEyRvqkrf
S/3JStqbclQ/i6HpZro3qFr8NyAr2TdxsubFRTSuAw97+r2A0SrCSH/DxGJ1q1vv2tvagzDMajOg
FF7ELhOLH7g2enHMmMj+mD/Eu0bhvBosN5l19+OBVP0HAjfCoY4PyVSFTA4MycneSIAunAWvBjJ1
jjxAufEQi/ZcnW2/aGMCfi4oyUq2YL8rreoeu4gubAI6WCH/zfRsiqF/834jtBz4CplhrVNLBm9L
vSEAWR3NXDQYmKkHa1v4Md9cRj+w80MwaLnxJq7PSvREKMm+P8ljgQs68gCgMgijTLuWM3/48yo+
03reYXLu+xT681ZhaxgNFOO6+enAvow7alEIeT7dw5MnhemOYQ+Yy0nETozuHYhiyRDoO6FJHbnr
AQLdlym0cCHoSxsA9VlGiI6uy2BE6y0AHPnDxIxRp50cmpdHEiXkDGMvj0/ved8M+IYRxcyDmmZ2
VH8KxkEFybxwQMPxJMb1SYEhd/VV+44KqAvIxESElRK8JX+iLiV11l9WBk4ryaVFyKpXHBGAsyki
SvavN9Xvk2iiljNBiW9luDtAsbwWGKHCNXNzn6f1Ak45PWgqbRoMNw9VneRTUCfQLu5U5USqTENB
8HhuIM/wMLwyZHyKvp4qiK16FLh97QRQlaTQFhuqG4vommavk+8rUjEIB/gwYBX9w17zZKPDDpS5
PDnpRO0sox3O1KZg5FqUaxZK7xCbFZvPYx8Db2mxLC/gA9/wbnc/XY1GtkNl/+BsKfNfQ61NyBPE
XCGtGQHaqcG1ROlnma/spEuUHUE147eUfvhWyPdDrFmzTGyAJ16NO7oE8UuvfJa/n2pjzCQ6DNd+
TuQnnbIgb44/xU68moscNvkA3IM20PZNZ5hsAFhA212FyfMvDT4SpzCoYYNRrF8jkKztsFmdt7RE
q8JfU/7T17M4LiATT2+kyo7n5keX1i5C8jx1s7nL/lT7q+pk6QfNH5102kea4wCqVPiql12x/IOD
R8AO0JVZBOAhUkms0P7IAJNNCu6fzIBGcHikaJFvsBOszBW+cTn2BLL6O8VLSb4A4wjEFi0Xyt3A
6gAQsUS7OoK1tXQBelFI4o3LRO3r+6U6h6RCzIkvyecAZ7Ha3SQxttvzw7pmLef1O4nlYdUGDre4
ZYFH9d5plT4AKIQydOlUSCVXgQge1D6G1Kfxb9RP3rwmmUow4iHwps2hasEz1xfE+dzE+YB0A1an
c9gMfZ5zplzSBaUbxhgVDSydPzW8rrcSwSoerHBQeM0ZqC3TYFADfgh7sJM7bmeKdrkExkOXcaJ0
hPngorTdhDPqYnzjJm1YmG7Fj7aHkB0gtxCJnJ2Mks/vVa6TaMjpHsCnibam0/7gNqH29TkW2wpT
0ibDQqXTxhmvP62ws+lPtzNx9Quk7npAI1DUWSrMUMT2bFGwWELJDL/qEb7agHB0aZz5v5Ti6jq7
4XtE0Dozi2IGyV2vSr5vPilwwXoWV8bh2792DJ+cwoiFBzuafYFoDPgX8tgm8duUoSXds+izOX7p
GT7DwoCAb8X2NrWDjI3lB6e3Bl0EoeCrw13u+8DqB6vKsbmnNePY4pQhss+kkKevp/A6y/QuojPF
u8mv7/HB6Z5DJnWphHwNrHs6X/8WnFJ6gM7nyb4Pk5LXx7PcE43ojHZpAyxx+bW8Iae+TrJTY31D
boyr7Wr6Guf+ak0rvHT5yTF0VSZLOExZ77ZUcTkVXolyy4H9Z1iOgDay1iJPKc+SIF6xFqcHuoco
080g6D0tFqj+x+aBf9RZZ68ZPp7V5mg3lDOLDhulVQ==
`protect end_protected

