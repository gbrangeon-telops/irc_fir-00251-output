

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
e5xVIDBGzQkhDoQ5sfeAF2q83P6A1Z/qsmlSYQJY5xTravGd4CV8IrniJyUa6zNomwm8ijfsSBDZ
3Cv5fk91Hw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
JTncam9YaU88Ye5zsiMSZerKzQZ8ndV/jFOlVBJ2+1NMrth4ym5MZgOOJUn+hqDs7WawEc66qp7n
dAXASYJYn+qFnCtyUAhIyvGYbamoaDWo5Ex6WN67wq/uxVFQHJyQE9mBWmFUuyQbfWAxdn0X8Ddd
XBKhuVWHjadjfvTndGU=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
WysH5jibOCiuNoaEF/J6UEux/f9qwkqszrQvmOG1LAQguVnzJ7+cmZtEvDLaeM5SMkI/c6AvWtXW
QAEuUSUqI7fc7s94OSdoy/EO2eWxzu/2PZr3+Vm/RDQkA2VgY92Mk7iTSAe4nvupzjwLJJp7MPFn
W0Qp6hutV366SMmocbalqT6lFUEm3BdJRb/waOPaQXsiK/eXFOfDC+OkXBIeDSI4U6bTS5BbTI6J
pFf7UmKKQ3+TO+1O/Q+2hW5WOgJzIUFjgYlL/k7HV9GLoiTkFeWQv9D4PmITDLLqEoJBQEH042D6
w9tSjJ90YaeXyJsQBc944KHiROaj7JIGL9ptSg==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
HfnNrIheX+bmcZCjcmnXLaiCn2W6T6H6Dp6dScskVGNGAylFhqrXsMMXHrPiUKf5LFkT6rGH4xNt
DnPlwzwiCAkQpMo27mNuJmSmEL1NZn19+z1IhIkgUjJMK+DU6V8j1HJvLoBzdBKXeOfEsIha7CfH
SYvgpUYxukUrvYeSdDM=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
FcdqosqcEEFjwfToDdg81IlS3kR13BUL9UoyGE7K0tYyJxwBRWvuEZwjlqyLvEdW74UEcoL322wG
MsjKrbrYQdHQMnu0VAIvQRAp+YUu8ZY/Amts9d4uoKQ4ceZKPNKKjhA2gLCTZlClOnHdKjhfnFhg
C4vFlIgGFFvgy7hYPvMYgUjBeujuUeMJVrfDQoBe2vY01NCaYs8PD38+MZrB1yBWXtoIH1Kudp5s
6rfzNC3iiU875HSyCH3s6Fgf+5qupOBLk1FOGYXDOgVB80WiCFsXlSgDSubN5g0HTJQJ5d2+rdH3
3+ADIpk9sqzMVdE2qp7yCA7kfUMNWwWOq2rtCw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 15872)
`protect data_block
876OETtVR1ihu59n4sN4K2GRVkbHKAgLcHx8Uc3gnNBFQWu9joveNwmF9XLaIB+cb8SdE2ppnAZH
0bwGhIpuSfUcV1pI/sqVgqwgCNKNitgs3kK3rVd6RuCY0IDm4vzb88WuIFWgNV3jFQqU65O8h0M7
eoC14LWdzl/H8pYXfaeQYNedziNQ1dS6FIMFZKHq6f0ZWKkZcRIoLzahnnR8mvrBil1Ds1M/PYLv
N+3cSozkCIKLeCbMipoOhZgAftqoM/UZpTjcbjIVm5ilCax+anbFzXFEdk+cCufTo32XIlvad1jN
fn3SyJ0VX7ckwgFmj+L3vTBBp6jrctaT/xm96DI/Bh2Mct5vNeEn36QHQLGXi5BMPF/SvCcGBDRf
kPWnCKgEIcvonhIcjws2EYzII6BXvhTRQPdaN/8lWIAEGhGxLOgwdauZHhUFMnB8FMl3ubvtQcXI
EDEukomabmctSG4Kv2SpBKZgmO3lStBFF7ibtB3kS7ad7QT3WvSkuLyARlr4qwiz/wU2PSobaNRs
KnOv+hxlUgAuqNL4i+yo3Cp6/q0VSEF74DIFEPV89CG9Rp+4HvQphg55AjPmjPmW1/FAOR6xK0NG
ZIvaZ/sFcYLCd74J7Ci+l+C7a5Z59NMRPjA2s26URbYlIF4jZe2P917Xb3QS7vlIuVtu+I7VL0Qm
6yCD+I4HFXPPPKneuzBumc0/OV8awxnvFS2UfkU24pYKIf0Wi7Hzvsg6Gz3paGwakBh7lNJFqJ5+
anXvqeqbFVKRIOhuFpiCCAhWAGKmOQu73tVdT3x6QQqTl9XGnrN37VQeoQVYthrzPJHY6GPsliRN
SXMG7ilLD1zZJJL9NZ/+Vd+/JTMiUisT+5Zc72imvPWvTg8Xukb9JQFomNCZBIWxUErLkZGTgIxx
yfSynRIEcF/2Vf/zGZNXRBrblNAFx8mmtxwqCIk0nJYQ5rtSQYV6VFbtMyWdZmkqqCxScB8FX+7G
72+R6utZL+85do67S0z8hCeJgfg3TFLlXaE/zlWDkpG6lPwYAXuuGAcX2esDxCy3mSGTXBGZrwxd
JEBD6AUhfUk7VEDRTETV1kMo/KiY3MLbyYZVxytxsjkBXXfJV66WcWq9yM4q6L+QT+RZBph3H9FL
DdIiboAwH1IRInw89/1fARYWBD9kJgUaXnPh0c0TnOOHoYdMlm6CIqPN76EqBT7gAC8sC49bbxC2
/j7HaeRo2NgJEdqKysgz0CvCU89G3utqPbqFpH4I3YK+o1n7kmhvCLM1wibTT5gldIKUmKeKQ+wm
Q0iWe5giBHlcGP2a2/bFdp1RSbDTWeAMMzLRkU3UTj5OqZGLb/FOgaUMUqiQOGIS3slQYyBKlHNs
0OrDGnlTBIfVvM1o7NfR2JnH5MhWvGJUJoXc/+2CGG7ZsXGpyp+kbXrEb8eliBCeoUOrZV6KCE/F
kN24WEIBgCh8w7R/4EL9QLmjF2ZUDZf5xcEIlTh78MJiLJqChkFOBrYKdzkpj3qHODCVj8jkzqnf
phMvTdIJglZSQwbMjVzQ2LQT2mY40y0E7r+PJvPnlP5cHBytFadcvvqAF6OfGw6OqGO6tUfuQyga
mK8/ZC1DqIzec9ZwXaPXtOdCErBnrGnuacdeb8QtUWvhCoLEQOxml4ZdCnN62c1wnnwNKTc5JC0D
FDGON4c9Lv7gYnqg/dPeUn2KQeRm8lrNUWnUccWOJPlf3tFrrbj280Lvm2shE+Y5RY1QaCMtl0sA
F7PKBM1o252+WkBVup6+8TOn3heq0TBtfgybz0JmaZW72tTJhmKiD8p2f9GYBe7DBd7oL5cwedz4
gAjKmNWpzF6JNzAjgmNDmeuhn4uI/7Zf+Ox09Np+lv9GrjfCvpdC83kB4QaGlWW4fsTuvafVwZji
HgzO95cLjIAgFDWY/xpLUy5OLFqC1L2G1xfTg52C2z9W0hpxCUAZcGpPKv1EWdt4GUk+un6lwwqK
a7SQ6TZ74hkoSwTPqt46sRvBbJfCTdZrAYwccI1LlkhGC4QQhI64+x4B583sHrORji3+Mrzw367k
m5VsHqME5WzVNpYY6CRTf0jzVOECyx9FyYyIM15/7uVjBnTgGb/CGMeRQ9lKM0/O/LD7MqDp19XD
iwOUZqBp8dj4KZgx63WA3tCREI/hlBKtr4GR1ptwuPmVvgQCCyo/t7ZGAMuo1JC7XrUiX3xfy17s
4uFOTKeUj+iVB7pogXb+ppIj1Y0SQjupoS7VwAn7p6/yHIXoPg8wAIUAR6WeCR0ef+v0sDgJOsiw
VAC1oEK9Ms1mQ/dBwyP9X7RF/OK1R2vD4Q7TQe2bhitXnoD7pIBzO5jRrk67sKALc638DTTOJjhm
7zUu+Ab6I5WEAaCTXUeUzLGuIbODik/Fw9yOTJoqUpLskCGHB7zMGKyG4DWN+iBT3wa1SSiC5crH
38kY062EmuHb6gaWZma7HzuiRLHDb4dMSKwCbkicXH0zpWEnVSnZRZ0A6MR3GYSA0VbwBFpN6mqg
lgaIF+7eppWPPNSF+o75BbGDc4JuXkWYpAbvCvCI8nzSuud1//CbCuvVm894PlTrgxiaUXbno5pk
PxvL3nLkwgl6XIPir1/ixWTZNcUMaXSlSZZLs5sulSE607pyuiyfuAbEEq6x2XP61cz6RvjXaPPn
W/7JnY1tVFhn2eQ5F9FBOkjUutEsACQ7dPNKNgIUmodOwHkgWxjulDqZo0mYWVk2V1Xg3htp0x6R
yZyV053i5MW2eH/p7S4HyEwBlrYny2Oav3D7VEhTR6VXwndpS7Jj7513cjDnMhCuMD+o79MYa6Sm
SqKq5wxWPM5PdPtEqqlHCwUAwSSei19octzens33sheybI4HLodzhzsOxTd7MNhD5xe/gBFNef/X
YlKHSOjxf1by0nOy0sa3NjBIxvSkeO/jCJZYEZPce6/QvoYhPLrnmZsl0lYgew0xUWYKo+J1nidU
9OlBFR8itY90LVXtkmfRRgymMidYMKSRrZnKnSLFRIYh5rQKnYqLA9tfhYbPEdVpqFB0/UppTuVL
woXVkNzvuJNs8jqh3K6ZwDIhK8xD17lIzqFkdrJvWiiKpgNcMmvXXiycC6R2f79cNCzb0cF2X9ds
PhvNhu4uYoIWiBZ7QBi4BFO7ErSo9fScsNgqNMH3/DS5TFS4lerLEoxnqLiDfOYyv6H9QIRzhx0q
H8nd4ePcBJDw2VrD+Rg/Qxe13aGbfSCZ0sJxK/M83IzkqQMEYnrCQtQ2FkbZey7a9GwfhhuGsfTN
naxi9137FcLvLdJKa6DTyc/g9R1GOLXtFdDbDaCoOXF3xbSvSWpc28AGyqS8K3GMu7c14D1vMGX+
pHyM8s7CQS7xQ5nkz3ZwQTt5TtoAhMc4Qszqs7EAYhJrMRDJxa89SWCLXGvtMZm22JGVpgaoghL1
wM8aVOECvIlI3cu5B5Qgy/YzvlWcByHQzdDmbal4r1zy6Xq4MBVwrX0+ZgSXcERnRhLRrnPO0qcp
51Hp+6aPlPoDvsEPCVI1tH5ddqeUSrMkJXRHrTotvJiimNNpmSr/pFod1fU4iuvdx5ywOp5uWTwY
QLA642vUsnX5U1eVbr5fY/tbzwJw3A/+0teK8Yz3SfEKepBk1ahJGGDSFMIY3AaVflKSofrQU5QH
aYAc/6WWHZRcy2Owc3CL058iX+y1KQTobSRkboxmP6cpyhVsRXfQ75PUQwbUnr9f2TdcH8tXcvZ9
9VBPS58U/2tfllAC6fUzOWMdnuDBgw9MHDpAqvXdpHntosUJXYuBKnBktpOwX1kyVhBm8qjG77y/
xV6NK8G7XrLBhuiy2l4XFR2fSR9TCw/vnWId5X4YOmV1tT2WvpzUJ102gzeqDIvgzgWLEkZvDuM8
9pD6Js0jCP2hBDMzQMA2DxdQfOknWdHlGia9/H6pCHepd5tHUZT0PrC0X5gmBzDjmzmuOhW+99+a
VuxA63yPK2pSxCXeHMp0wpnvW1JEgjK0DNnCJvWUCEFG24VuoODWGjhu9yGmQyJRQgbh/LeWp+ZP
crawqG+1T6G9WXDCpPfDqY6ctl8ia9WYt3LWAeLxCFWYFGok+Tou9U6ciJ1jORtuJ955MxwA2EU6
RlM3kJLd3nq5rwPNpIZDj49bbLnZjk/t5LyGdt19BDPL0Cf5kTNQybmiAZpgZJ68h0tzvi2rRet+
/WsuJbuhJNH6tip8nBryYxnSYoZ5Ax8Tc0wG0IYJJ6QMJoZJIghiL3mTrRVTnwXWjpk7iQ7fC5xA
Pf/itNnvGVAd0MFDjtnkxmi/b+8Z5cNSsGOixUbBScmT9jBLxUVkLbAqFF5qQkCA1VQ13hEBnIWl
JEb+YVDLPi9e9BQYy0zPbYfiWE3Dj7WjzlGmiah9OchoyrxAhnZYvm5Yh52nKOzHCEcQSXYoZ3Ds
zhhRvUOYemR43qkS+Todm6n7uoTY7c9Od5UOADW/zFQ2Bky5cAY5rNtZjbGZ9QkE4cB1o0FkpZqy
g3dohatLhsu73MbngpTYRQK+roZLf0+9/UJjS++wgfKgqkWAxZv27ErI0CNFsiafr93ZTXg7iPzd
RHJsz6FpYQ5hx3bey9udixuIvU6s5ekW8UipFXWlsyveC5a4SpT6qzr5T0w3DVDgkqwS/foRtGwO
NaVv5+3+Y4hr5EpHsrSaoEKgUKwOAuZShV8oFdBEDzU37FdkyMl9YLZbsI9eBLZhY4AQ4Pt1dO/e
2PIwBgks+tiJE9aKoV/pmQ+uuePYKvXLbW0KF/IQO3HOFMfKVB15H2IQSTuRYOvPAY4eFq2U3Mc3
dKiGUCWa2mG55Ns67zx55x5saIat2zZl1TMsJsf6tWByz8ERUGPIk/y5ZBixSQ2fEeHCfKeJAeP+
O1aBEkvXHhYTwaTFCuBy3KSkswnjKIun+904Sxpj5WNEOtNVkrMk8xKnuDt/bcayjOic+2E/tH04
YQbBV8VB41c5C+f1PX0IWl6rnGSpXJzVWHqY60+accZmSONWqiIQebskEkVVVLyCWkpEgQ7ZS7Un
q0UXJFIYqvQMg9s/SKNI23/3EpN9l58awIfy7y0uRjB0hk1qyHhMs0kg/UVLlyQPBbhrR2Ck/3fI
ZLs6xTRElfzCXpnXzFUz1U4CgTxnISUklHcLLZ5qmSq/2HwBD/Yxmj1TdG9EeV/D+Cys52/tzKVL
MNT3o8azvhRcrE61USjIWe959tvFt33Pm17TJWuH9x9ybO4wQCHei/8iobf/VsyN3i0RDx2RaGrb
3XuQfO/S2Ij7UfFEpnGib+9AfM6svv3NVcvL72B7yWYPiyHUM3usjPlIVCjIjYV+fBHx/2M/xlMm
gSPQrmAD8zyCPoxi0slA9n54Q3E5FQl8qAyo2izqNpJx6q6TBtYMOVcD6Wcj0L3KulSyRvA4758W
L7EnnVntZ2w8u2fN03nTx1KW3d4KhsSO+L+5VB25AsXq8FfnW20gdLbIGF8QnG0wGTk6g+9PtEa7
VTfaODm2V1tzrlaSLeEsSW9f0AQ4947CVLv15flUJBhDIZ/dfJZy0NkESDmdAst2pqNkmpcjgEiC
6BByMWbFPk5Y73pjFh8QbAdvP3V3l7QtS406LJ705QsTUev6cCe4mnLv3VYcyyqh/Tb6XatIKAlr
hCq0ir2SamJFL4sxWjqu0mp02Eqd26ECfdZXSFxmUUvAI0KsVwtoee4ir8Oxmlr6BvSze9IzAYWx
E514QKdhld54l/aPxxvVsa7gkKuZXgRkKEW843HbemLpXnrl+c7h0Cw5KqBjYgy8VBMWmE0LJ97i
EUvoNVAkkAhYOWpZ7GOLB3yYfkDGOVbyuPSwTbwg+qAa10BUwSHe6SW4iH1+6fDhZomlLFqnpZQk
vuHg84shDTiI+OBcogVc1UOU3hrON966B7l6sKJfm2VSYHetDxCj1wkiyoD5YUfvrkpRb5xK2A8T
BoSXmA4xoqR7h9iSW2TI/GGrrDOJjenmDiJmw/3B3eF75NtfF13PJ24WGxKhvj3XABEUcT1ajhqy
PzYgTx64Regp10gzNgAg3UnwUmpklhUPCtOxGRdNx/Lb5CITM+B2zPyfDzQX5sQRfhI3ZuNR4xxw
8m7wMFSO7VO5s2Gtng5OstnABEq+t/jNsbDww3LEFcZcw3uKPvtF5pHi32raTt5k5SjCVyQdlYbz
YJT57IB53R1odjeOvhuZSsDEuAFMRGDGsU8QYEoRh212evckeV3jN4ZmL34FwJ8TNERypj+NkYcv
lvb9n7W7qkm9BtNPsXLtXTM3rK70FgvrUAnRPoaUaTmGVUnzaltnre8gLrGSQv2gcnXoGHpuwQD+
zLNcNl6lE0Q8jDEJhz2KbiEbjs6ISmjOvYISKHjlU+/o6vdMvL11OGA8a1Af2zCxIYWXzPiGxKcY
xVq1lN4ykjboHbuKwTJahQFWg39PwiQ/z8+s/X0m34OXwNtLTeLCmnFsPNMbcCqgz+C3AnqlohGb
7/Fa4vJppPfbefEX+w6nWpmvtYCphk8BgAG1r0riMhf7reE+c/n+QAHzLKJbC2XZ7UImhVIJjzpC
yFMHx9bJDSUAROHm6x+/NDb8O2Kem2p+L87vXGtSt+0Dw+/uHRVmyRUDJJVYR7hPk0aSJE+spjjV
BRou5nsa2JEO8Hkcwn3rKu7GlqkeFSJYi3ZZFZqhgoAxMsBJ2oOUDUBlmgSpWTVw3HrumAGDuTJH
z1p7wHW/h/z7ZEwpnntm86fFWhM4vj3iRn1lACRe4/6TxcHoNWZ3snji8xlzqhFSQjE94N/tyn0c
vJR4g6RuflLMcc2QD3PmeTY4/s9/LIBCvCmIgzz48ALlRIJxUdwGRviW6RoTCJvHezdtLMXuZnrZ
2FCOl6GqduiinuG/a3lx/4zBnO4EJ5TyQN1pBCicd1BDCuWoXgjMj5TrF+nUM0Kn1wOjAkS9dQnQ
kYtXaUgHE9oR0HoV5q/5R7Y86ph+WST5TZ0CfqQ6GZ1N75JiKSl4xZ0synrmVfx4ujCguqEUEp7J
XxDx2DLjreIO02R1+ufAcxg1BGMk6r4qZeq75uXqENVIbgeYgLG5H5BH7gr7jqjqblbyf6Azuevu
32jcSnojLTko8oigLr9NZrgXg9b+Uh3nFCzTkCq5gErEtLnhpaqFYVBUyrvsz+lBOYkv32baupQ1
mI091fBMNK7o7vQqh6pLSTca4GHQQCmU0GkdVXorlPGaRu5L4urG7m9VkCE/4sEV/g1mu222Jv6K
4DJxik2PtzsjDwaGMReZLZZ/CObDh/gZzSRUU/XUFtAQfth065tq1ahLkztQiKRBDcE8JYPCw5DO
6P2IRA1JgoIxydi1eiXz/elQRIH0amjcRnQEnUMmbjgsnABRw6YXprF2jwH0w0qlN8XU7hyZ9GBn
UPfvKF27IoXTThlyxZcYY0EYbGGgd/RqDTQaCb2H2vwsCehnlm+KFK6jsJ17ZZqbHJKBLqoV0DkU
z4dLjDhvD5C0/teAW98E0nZBq67vwCfs3+ELNBwGKbXMK3jZaQRPL+3XWZX2i5BnVx2R0oHRW79s
GXTMXkwKJnuuNSU5gXVfgYFipkRNiYYTJq1JZ9VYs6I8BpkCkyJ1dBVybABVZtmf7M6WIiSDZ/XW
Hl1Wacyj/uQKtgvVSPXyOUg+KwGsoD8bi0/yHSWe4oTNK+Kfz0lVGD+Wzfa5UxVs/dSUKYp3mEia
ZvN557VArbLOtNQt2GEOvVvFEGh3col4JQjtQ+uPW90xsECOHkuB7Yu6eL0cSasSIGrqlcZDuCsI
t1/+P2SvNS1YZtHC3ZUEr37OTC/o/3E+y7yPohvHJ+mtllalmdX30ArYkKxP9ZuUctHdBjpUkC+r
R/C0kDHohj+xNAf1Zya2Dk0Gd5drTjz6DUCFMmtD6nLkxoCgnR8FCo0MQWtWgYUPsUHKF2a6ELEo
0W917gEf6YzVV8bsbfb/srHGyUZgqA+sSusfWOzUaaN9cG3zfPx8ZvkyNTXYsizH8EAtfgO+zYOw
TqtWwQlYQXv7KUyu8T/HG5V2Cvoe8NybKkra0lbZGPNWoVhh/VE4R6Hx4jU93Jp02RPVGM6m7CyK
w/ggSlDcQvU8InideCt45y6sGYc09manE8iYm7dCE/Mbmaw/uGbE1Q1Rh1SK7o/sPq+ytFjPsm73
B6il8wyl0Tj8k8MJaHXZf5t9Ctz8fgUhwEv8FQKYhasQfrntsYFtH/KxHm2FhysHM9jgB3Qo/qtY
0UL8O9Wv+g82Z2+JklgFPtjbnR4N8534SwiVVwdeh8/VcBUO5AU1clV/jhAyKFbYOidnbxH7Qqdb
Tw70LxmI82QfZSHe6Fn3bz/QPZT+xTYZkHvoGdUSFPHLk7wUZc2PRpofAek0vChrmduDBaOT37Cu
kAJA6+fYNTBZTdz/HaUkvt71T+G9IsamcRVFR7K3RYpmEHnKVEQFkefaI+ygt8DLpJR8HS3vjwuf
Hsah70dYmmP/aK29zIGKCkVZGzO2W1YkTi7vy3JQLlD47yPMq9mSperRXZYkuD9ixc3xxLnHodZn
sqlz5tT1CfRhJ1tq5sOKsWp5XSg3jnb4eHL2O+SgdrJCZsvDXnIxeZUdi39xA3GeR+0cTHxWRBmW
Yyqc2yfJmwCe/7tYEMDmqPJAmD2vZQ7IMiNwPjPvDMM/qrpYGdF1mFfq1jbRu4Oz3zV7YhzYyCvj
rS2TnF2T1TgiUK9AOH7Rp6cdo13CvQxoFqYzULc2VVCwTuAdEevvqYRA9OKIyWJN01RCz8JDFd+n
rgIiw5ZhJknEBU4Y915LId6iUKWybqy4kzYWZ/7CXVbR2QRtlqeW+gxfmVNJ4g8GtUwjiY5xjfVK
lqbucYkU70MHe607khY7sh2zbMg/oymD0Qaa4G7ijYR9/x1YVmj+YFrpE2qsFxsPX0/F+oKU3+4m
/wmKnpOs+WSBgV56xdcMPsX6by52NLgXkrwNEuu0cs9t2U7GnS4TVA+sDa+CD5yymMsLKaBvAdQn
9xE9CW2LV+pXhLlm1uZOcDBwycBH8+3r9iKB5aO/Xi2KSL/YxwpFoV8Pb2sg7dWO4CyeDOd4ZOqZ
PqaXAtJwnRfQQt3+O+o4pnZK7oYUVWQED/kUIvb1ujxp45W3wd4EpdVL+nL9LOUQUEllfL/ossGP
AuXCf9iwGaRrsGDc3jdVKXVux2qOHkJUHay+MWxo4oUkp2h0/lShIUIXzbOSl51m0SAE4/7VPhQ7
0Eyad5kck9pOcYTQ9rsXqItngrPinZjW9AF+0zeI+/gmGPLH3J3mPZfQsbY9RpWoCPv2agf7oG8a
Uv2cAxhyYPEU5EqIRNRSieV39LA21gnVSlLOxGizBXfxifUbD9ztuji9vzETR14yQXAQbtegtoht
IaZZQ3PpyIsV5frJIhM5NgRbRHYdWYI9mxF0Of+eSMsP6zLEqR7Q2Ij03NDNguxnHEN0RM5t7Pv3
kKK7nnqrBwZkavqhAYb2er1vYBsPhVHz9so8DaW8PXOL1WgAiUvJ+xLLUgZ0UVFs0FWmDokMuURI
A4rYc3rthRRhmGUAMGCifzmv86VT4gc8QatSP5Ps8YNKksaJoaIKWrZ6nhdOToStMwELtfrOJhCg
ZM6z8Ff7rJlu7gEpXo5Lf3X0C/IfjOzsj3smJ9Xtg6TNTp048i+qPy//ZEw6Zjzpn0mFzEpr30SK
KlJFHAUDG2W9vaSOLZfj11YLShxBhnYVdJ1XxJmLGmztiPFyk+oHgCpAGxKK3V+DwEpOXJCW6EF9
lRDsyDmJo8W0VYicUWBcYK+i007cH3u7EeJeAx0zs5xhFLmMNBg5UV7bE6+Z3N44gYNtoab03NdX
RQ1CugbZxBKxHMZxcVGPt3D6Z808vx34e8/PEyAwpQ+OKSXhhY+Cp5yjl+N9jwAdh1VwLUvazHx+
HIp1Voi7viVc918St89K9jdiAwRi1mFxZIUf66DNzKuMs8ckBCsGakP4ljk/kvm1wclph6WlA/SP
XBAkzbaJlBZFAKscAZGrtE8Dyy5bI8za0Rg0x7vMFiinjoD1J9T1wDiKTkkcfgkKkfaE5cw8FdtN
4ICgnWScOvUXAKXfNHPqekWypMkiG7ihYkLKWQY/tWclz8W0yKA0Nx1Fl8gEDpHe6/AM8DAqeCRG
9BaUz71TPKwSyjI5OrzPvRmkakifPcFoUWuoy9t+OeZFcwF/6oAh4rMbR8vBT13TcjeXBeJD/biT
kgsFr1sjxAoH+DZ5tVmFAncbU/miCqK8+pUA1mqlod3sfjTPFKXajmSf6PA/21Kz0FlGV6A854iW
kYhbIrVuU+W8keYm9LuLTwXZhM5zD33u+q8GKU0PYn26jmyfYkHYBITUC6qys7/dotlZ3v1HhZt0
mBD6ORTQ0HdB20omMwaUgzXNpSIJX4LWlY0k/Qv0RP/c2EEpEsUTxV1w3u5sPjbdM/k/5svy3uxQ
LMaFcwr78EsHqX3B5tgfKT2A/4IjJ7L6msAC3rPNS02rJQoessiUmEy8QqOM1c87scenzz5qsi3q
nkMjsI8hKt+CKfYpTnSOKRSYymg0/IGYwR3/XSV865LvUKoOdLLsFd2DH547XVybCKYcASCa9VbI
2dSuSHJYe6fuVX4saM/Y+QAPGYb3m2LbNkTrqCCJD3LnRHZ8jjqPV2dWHK9GsLLbFY6uS1FOnNgz
YsUCCXtpJ3PqBxMz32gigOw7uUCdz56Gm8/BzOK6hVTqhq+N+chUm+7KTduAdHtJ3bDbCbJIgi5o
peAzCFM5C4vfDA0q6yWa+4quw6ZypkAP8rGh7ZGG8SwnpmvglKpkuunQTU8QwrX5OZbVnX08SBe/
aB2k/KXBxZAQqrtN3QZkcFXX0ROLUB2mcDlHvrOET17Q1pw2ufl6w4ZmwQNwzK3IIZ8UtFHszsJu
0+tBQ1zLl4PNhqAZwkEYG8qKE0plgBWZ8tTBVx+jLdY3VQ11Ye0lXWZ4PS5U+aAd++Gv0BpGJIDu
ovZcAzwYtWQsKUJdUKuSkZJFexqRWNEk/J9LwwwyhjOJbyC5qqMHzZdZzEXMohQcEWLegLPu6Mh+
GiBsuiHIa5rTkOrcEJpNMI+QNzJVa+CQSh1Yot6jwciA5CUp/03jB9NrLUNH1PuWEMHckAkRhC+e
62TtVLvmxVyCiY3YaIyTCCVIQa1t0FvM2szbBNdlkrXh2+Zzdcj9UwQxjdjtGcYrkXFhV5J8ngRf
HhLtWHusXRtzau+b8mmeB7eEB3oR1rrT+Nw6dYLRBURfS5wYQIPVhESN4YE57J5D1RcTqjKIP/C9
38HGfkcUNMOCZa46yUb9W1lsxBufCbhdfpirec5hVXFDbDcrPd49iUWiKHKLe2fPbagZRDfn1I1A
wDZbh3i195MYorsnVzjZTAVUTUPj1Z0Z0Vl/pinVql8owj2VgB8dpHJkgYPC+KiK2Mp7maTjOJar
DVPZ9zf7Uo2wh8NSOajt6YNa4S/totHxehsjeY1IWUlhd11qW5sb660bVX14vNFQmjGUCCb5+ts/
ojZMhJgOzGCf77BZT8ZYb4OU4ppBkirprNDbATKq/nf81bYWH4bKFJ5SGqByY6RWUWVJsz0YqJ4x
AJwGINRBbK5IqnHU80FaM6Ds0xv7Jwnic49JgkL7IWrqI8mRVHH73BtRWKnZ+lRUM+kKDsiAQW2E
a4s4dmOOlzg2YxsI60sNWV/xeTNcp1mmoK+7VAKLGUiRUZi3a3im4+TDjq9LYb2AOqBMUks9NKxa
P8GJMDlGxM5NJsyQHfFF5zcI424mNTAJZ6qawS9xrlbrKSAZEo20JpDrM3P+Z/v+HuSRU6bNnqMj
mpJN8xLLc1rUpd9Dyj8X3Aq/cVEYiS3TfPyw9G9YxRL99IVqSMS31jkyLnITSt7d/4VlFmCIYQ/l
2spmsYJ0PP2z14voFCVkW+0UhsmQWrMEBvaj7xrzpLsg9a4vI1Igb8jnoS6McGKlt8tXoCGzfo47
VhSvgt4gX3GjyxSUkC1G8kdIa5y4Ktot9WGXY/COlUUwWsGtpYtSpImKK0sZUhNwXMN+2h1PDBm4
x0ZSUMI17wFzxsbgLMuTG6WqpeUCimTSKv0KnK5hVsQDjQ1sMBv+au9gJyo1wFhKcY1eepjwCvtW
EITrk3835uKjruc5ODlKAfKNosUgkDmJBnBBCIeEtPlBOwcN1IE4lkd94RrEYM5utA9fr2cvoeyi
/U9t+tw+sBb5H2qv92GhqEaNG8cA+0/njRlSEPSYSrv8leQFvqPdOx7k15Gpmo+Mqs+L7vXF7nps
QckEQBDjsVbDju0b+YUExs5nGBVtADVUEYNrHFmemCTxV5GbGi/Qv08A2Edr1lvc1NzEhEAt1rhT
EjGCMaSKM4GD7Mr1M5b7NI2HJ7/7WhXj5r3D3/hDmzPdvaxyZUrPTr5IaUvYW2egOmj8pm6ri1Uh
I5LU+bV+OjyWvKczOdYcOAjTD7URwpiVQmxRZ3fwvZgpIa1d35WFejI/EfCND9bAQwFRH9fE9VG3
988r71aZ0q7sEMhKvzrxKm3H+f3jd2eCmdWgx9O/7PKN5empDhlB8tEnCXFaF6m8Syg9CuR/QkD3
rjmVXjb8BA8XKizogmshxOXX/68Y974QRj4aB+tvh29RE149uqGV4NibVUZPvEByD3uF8aPHC9nm
mTiIcrOr5y/zKqcxxNPagNhjfoGKL9IPZOQJMGcVNYvi+rWAcsjuYrH61sd2Ed3rHR4UqG98b+2R
6ii+bq8gA5bXtIfn+MeMkmC1cUD5LlmCgiBqgQZSdCmlRfd0FuSoZ2TZcVMkMeqxwSkfLqKVq9D4
/41V7b7ZKYKY0ykvENOZ20g364cTfmysPSCOTqVAsgkj8qqsrVRpp3Eq7TsFkl/xvRBWl7wZ/NWl
nQPzgswUDOJZPHiWSwtlWVEdJ4AkMhL/AOqVYckFpxcN3lpGiM5e9anLlX2ZZ0c9cUg3Mdn2zBTY
6B28ms9fYda52U1+03tgl9gf8qiOCpmiYAhTo3N1YE+xyqZBXVym9rXIo8aENljrrhxWWQc4gmvU
2Dw5NRMAwlSGUZYAyNtTFTBYb/mBgYKSgPZpvf3zW84jyo8zqGtfkuppy2KJ75qt0HVIaJEbr31z
kXmgdpVNRpKHawHvFC66ptvVZZ1oDIHepFNhm4URdCl0owTfJElJylZKAwqYmTL/M4xEb8QEMnW1
wSmowDVlBUqkkaRiBYUPh1cTd7Rb2VXcqSuoDDkZRUPG8GblD+cKcDgpuk7b3YlhYLthTpe2dunf
6L2JQVgePZ49zF36w7Kk6VFhu0XxgYx/SXSdD5Yqu4ku/tD3v0K0NxE2RVJVuAQONYDtYt/9UJ1O
DQSxhWEVJw+2E6mHM4Wp2vDISHkrMxN7f6xW493fznuG3vU2xatGy2TSrbZfetXcJloqngWcat7a
b75xkeLdKt+3exhOTeCzwV2XTH1NMWg7NF+R6irSTNQJFJu/K8Er/PLqWaBYTVl2dsyHt/IiC0qF
tRbPEbSsjEIbCnD96lhT0/Zymn+6Rr/Vmf51+DcMPJh/RND1P9HdL9g+b3Kgqh9hXnfr0MtQlM35
Rk+6PSo4Ld9QAje4Vk/R5mdI48O72nX+vxTIbs3UT0TkNRRwUC2nUyHru5l6dBI2STHKmwPxzjT4
KOvJHooF1Ku9VVuIUhi4VJEfIngvKHN3rvjg1Mb49OfW//ZNPr5jbYZLKXoRBncFIv/ym5feDBJq
cpDippIMXHonQVPE19MLo+BtfAMtx5j4jOk/ZTCL1E2vtr2kM42PNvYSQ1+C8QFlNhaIltABW3dR
bttyX+UMpyY2bm8XrE8/Qe2lZVn67pNv42LGjaLRBDs6F00dFaQ8KLIOtJ+HxS5t2E7V+Ak0NLbY
o7434DxJ4OhkC5mIR2FQHRlkTtlyUy7QIslq2ungUjwCX3ozoUUYGVzgYG9R+EvMWnmkmqAy94et
FmMabzunK/sjoYVDdvXzbrTSM6aeNurqcOUruT6WHgEkAalZMbzdZTIVqU4NfRnDrBKo3dGUSjW2
Ov8bTdZSfePxu0uKe9BqooAx04Yo0ydu4+9p9rt8rWqvmvB4nKGPy7APofo2sJK0IZMQgHsPB5ze
cpEBHERtS2yB2ynv89r6u0Zu8pLt/xsP6Go2AY8VyaUUVl7K3Wf0+J1XgzWmpM1PxfOCXTytMOGE
O46huK5JJtISkYA27QEOm7lYSuFQCxgIYxMl6PP9Vx3kiqy40520+9HKv/u5Vu24uNpMY1v+Z5O3
gN1cneReU/VIj9WYIl0yUJx0Xs7Qa+uRPy9Sh2+fArIgPYHhttVxFM5itlzHzqY0BPO8Ccl6CTIf
0wu34rW++kI0otLlxsynwrzVUwR8x9HyQoUkL4JqkckXHPx1Jpjvg344ksuPn1AMnyYad+KuF5vW
lx4ItegU2D/3dP9an1W7JeBLGE8Zm7ad9piTPLMO/jr6yg7w58PbmhMYVpWSdLeO4tb6wHV9tB1Y
D1tKD1LBl/ZWfc8fUOIzi2QeP5KfdzSqn/Xhqsm3M4z+jtPrJ96/PmF/yimYKvCq+XBTfGQNH4no
E2cHMch0ULZRsWg8MTep+Mt7Jermmc/HVZFjsJ2HJRbFi0siVtXG1scJ5oQYXRFxf7SKUL5GCNXA
/Z9bTThHoZFm6mWviT2RFqa46rWy27nAKQgNwbPaTn//3DI0HLk44C4XIzHbiyEXV179Mf3tbd9i
OTt9x3vmTM+dB48MDU6gKaSN1LEUb1vu47iWMv8MlhdyVgvpd0qn7jwH1CFmMxstKBfq8ff07E/9
SZ71N9xPw/dyA3CtGPvC/vbwAm/cYPWK1WznmoelLGyZXmq1lZI4206Zt0/K+sS7OHScvHzrVlXw
coUveG9rb5j8oAWyMi2xWJxq+H/slE3b0jeBIOKXj75cPFkuTaV02se9Rgg0nuehLBuacJMA5QmL
i89C/vHTBSlcA4zWmNC6LnnyJuiDtFog1DG+jaj82gkfho0KpGQybsaQf6H9j3s4LTytGLvoyyPm
GZeCI7Yld2SSe3+trIuMxwKUe9czk5c49IWqUGSomP9dJCqHrOu2gdjTX8MkixZx+KU8CLdfjvr9
cSVGnZhCrqY6P7/GIm54NHl6Md52bgC4VpZoqWgDhIq8UxD9D9IBtZxs7+3YaZIe+P91/WCPrDYf
bxwG+42L+oOooe04hEpCkKx/d13/plF/SSNOCRVI6sF2+J5jUCuNH6DSUL0zVt+5qelXy96ndSNb
vvY0mCvODg4mW3gfOv+tFgpk8VgP3tFdQIsK7XSJ5ovH8/XfUAIlEMPkwYUvbjj5mjZLAcaJTa2C
QQBBKFjwN9YlUMnYNpak7PMtKmV48AK/uKR34vYg1Kal/2DBuA9mo98pd8+TD7O/8ib3e0AqQvPi
V9j4ntky1TEpjbchGp2Evg8sI9lheBmDE98W18YeiYAIA9F4DgDZGlzzn+lNNmbwMegytbHM8XY/
sLC7uD4eBkCyQoMmqAVIEYa736n70Plo4fURqWKdMXZtMyreTK7ddCRdcXWE157fAYmWyUeoqizY
2rizeTO6rWnMZJudNs4kSR1exOg1mlxG22WqwCoJM4FNpzUl56oSiCCx3+6vYZeGJSKTcxY4GqHd
CiAECJLZYrTIyv9yL6/dfV+5QiEJICohOpIS8/5vbFzh371XdvD90FiGoz1o41nHqQAtCuNAPjDw
qQJ45MeeweER8wofWjyZHLtku15uhW26kgs1IjSlGn5vwZEmB82L1dMCl7huWkrAHVsR4ZAHW5ND
ChspdbTOV1s/4LrYNB/GRQ2BA264JFhTkBJWAQ5+IRqsVq7GSC2ulchSKsl8AlRz+ojZ1zRRiWuU
/BOAfMVuIhJ/Nfe/KQPRv94YytJgWvyGAiqRDrN/ttnXw2seXAwMPlL871I6FDfMFUo8bPJevXUY
Hqa1Lf3NYirBWQjROo7gsbVLmA6frGJwRfYQ7H3cPQrUoEipTKsmpDny26HO1/k4WLSp2gC8H2s1
6Q/tRRXvAllnbtFSzu1TDWt3vR2p2V3PN3bJgNZ4S573BmgvZCe6K2+SRa+VsKnOGGLa99yBuT40
wKBMxO5LmJjJI9CKxFJJqyL1vm7XrZ2KfCXOFuHE15VDwwIcRwqiBZAoMqQcAi0Hyh6gEoSqEfqD
6Tft9WSmto3uYy5f8WYw9MjEmvKOawaqHFVfTE64D4k+LIbva9XdvtSxjHatWqDhBgpzaX2tM21e
83bvb04KPYzZG4Y52/DDLAdQzMXAOdhuW/OxQ2DgcVgDSZryvjua7DLb8Nxnu4rGaRh923wXB0Ya
8WoAr6ZxbZTYPyxH0JqiKn2UbZ6G4SXZntdJYWU7XxEDoZvjJz9J37EtVTDyQ1JNLG0YeaoWX+nk
OZtuVW8tXN4oDfZFpdxmTuMJCSZIeR3G8Zm6qwL/12Oywz2FNP36uwQY3SaZfAj87yE2dtEO7v40
N0O1I9mppNh3y7K6nz3YwLKTZlInbukKHef8MNTPtu0Di0KeIYF2HhI99eIFy9KtoGgSqaxiKWsg
ZVVZbv6bRD3JNGore/hmnNJJiESJz8atMHPeSNjaidXc2hmmY58OkZCAhlknnJtIzZ6K8HaYjBbx
Cn1HuIgvJ0xHNtGKMxnlBodLkF/tyWrYmYlUNMu8NBnG88kjaMZScBLgcVjR0OmwbrEopS89QgDL
zw+DHWvNnfxmmkNQBwkuGv5hShhZjdyyBmFcHnMxdTuP15u6CGI8Ff8E+TKEZczf33AqnRt94Hp+
LnabOBXn7QzJi4hs1TV9wsz8hacl+oS7iZMN2/TLlDRz5bXj81sOd22zk9ftuQUVySy6pX7jK+GJ
Z96g//wQDfTq33MHSNuAhwIVUQdtVmhdIQXCoa06mcOVKOXizfD2najBpG8jbzE4wMruXpzcd0jC
jUzh7komTujvHvDaaOJy9MrAihgKqZ7hJ9Vxih/FDSHXh2g5KK+/eh0uP914S+ra6GsWoqIBbOOC
Lqef7HMII1KPW2/5j6YFTu+3K0v+kKjS5RK9KB45mrciYlIXMWpuvOuczWIWbiOuaNHdcZ0mklf1
Dp/4frmzOyb8pT4SeD1AMTXo58vv2Kfxvi44nKSqH4mWRNpwt6jUIcKd2pKQNHWjEtrEhaSLPuQX
rUtGx1V6eZImJcHGNLXqKGyaDeuxG5QMr657vxZeflFcLYljcvdsmIJJXc0+ad+oWpPf/SdejkCr
ZHAbnVxsPuhIKvX706dCLhPQEnslczpwyyrzVVa+GzlfZLLfOUoTU7swcmqqHT7Wsi15uBobqFk+
isC1F9Sv+6xx4aXmiI9fscB4CKUAzO0wtDDKShqF+8TRP2eft5FpyYXqzEErSTDYKOAjKYS9+lgC
6gdSd+2sqLaqINSrWPRay/jNhQhgTwjluizobk4gvDLe9sjWkE+MjqsSeh9/mXoOgNwUs8iE9DxG
/5Fb0JDye1SHhRwM/k+lp1gHLQjncqHanxcLLcKyAwzdgVUy/x67IBcm2UudXIaxDnphXyd4kwLL
lTH+9+y6CR6qXav1DoIRgVgh+MkCeyfYscKxXaS0+pdO3G124WjTaoy2V3T2kgoRi7j4gyoq2d0V
oz0ItmgE1vLWKUVQzJlXoy2M+JuotuMxfQ/nFuYsAv/LzBp4/veNQj6ucxV+lBUfufNvaGzamMlW
Nk13t8TTCMVFsD39OE9No97aNyk6FWRylhsCBle5K+yhrvZrHEEBzNgYCieVChf5gK81UWUOkIM/
+sDPijScuNGod8zdYRBHgx667vUYASZO4jWyhciG/6ad45wx2OexLU3NiPxsTY+f6rODXme8PThl
wFFaJtEPbPb61dtR51ukVdEOXKAmF1z3FqTwXr50SjyVRc3S91sbYhbCMXpmDbF/df1IUp0eFPn7
IRL/HcjbfgVuFP5KYZfY1a8ex5V0TouI6pTuh6DjM/f64z9bcN0qGwb6+wgLzavJSOjj+s3GSDpe
nvUCz7xAtW3TZ6ulDo+b00Sk05EptfAS5B2XHOkbGxHp4ZnFwaksXoK4wP2AMZ9xvcOJnce7+UMa
myywh8CIPndzp7EWGdfb7wlfAnWx7eKUiPzLBkPRs9z4JlHG3248/Pwy0Jh/scNDDjrgULkQVoal
mX5gLlznUXcbR1FmAecq93Z1CFWpusnYJJrOVGGzo7/dk6hq+0bmggesvo/PIHhbEmh2emSE4UEq
iTebrwaoKMn5qzQ5fwbpvIUdCyfOH2Su/ffN7N8QtfG6QdyqFbvhli68IWzaEOmfiF8zu0hGQTAS
UWp7opplZprV/kY6YoHIUjl7BmTyF0p7i/rG6vcQdkOnSLVfWBe891fWBUnaUnaBgXz373qIxz88
9WBaYkZlK1cO84/04wh0QKSIMqVOHOIlIiZli7yqwsOzj506rW7k7VnQzwMpF80JMgr1sKJ/pQlZ
XEp5gmDI0GoKCZnJWgf1v8p0U0gYJWC+2wH1hnD3S4MRJany9Q4ih2NOyLf+xYg36wx72QSGMIxV
N/ZsX4Vzhy7z0YSfn4El3oAd15AIpw7g7UrOCjRK82tkl7TOIL8g3b4mglUcLGsmAWCUzIf6buYO
/j+VT7iCcBvrS5x8cgVRl7pMCzkEz/T/+Ctw92kJ64L0Mcd1BGSa05JkGV8rlewU/5D95CXLrC09
HgrWCjUYgx6BwJd9JdKYWU3S07WQhPxYZxnHN1SkkskesxByu48dKqucD0II1SVtoc8UNwIlqAgt
1UPRoATfY7sec/DST1CCCcClMK2qWxV2haSPTCM4j8MDtksmEgGL+dmts9a6+dFFF4unFC8LMdeD
PhgIJ939GaAvI4+OGM3AwtBfD6zrQ2ThC+nk4rVWXSslTxX65aw2HpUDtmU5hPB/xXtpHypClYdr
LGoG5vVnz1k8NNgH5L34TYK80pIbMAOgXe12A54k2AgQwc5q7NR75iAJJ8Q2IgI6GtGN+H4tGCHN
nNM2QwKCJuXkaQL6xpYThBbIQMiXmDXQJmfghqdx647/cE6T3ByysmFlBPjoHZa7C5kj1DA39MKD
WZpo7XvUxcSLBnxbi3+ugZJxwICwB/ET+jvN+pM7ZqIj8uMLQcZYq6QxPl047x9XA5rjX/tH3C9N
sl4goEZsge8CNGKk8+YpjuZJCtPMRyriJSDV1eZnDbiwEX57Mtp6Ny5nQZoTkQg1TN3/4Y+bdcT8
HOO1lxmRR4Ty5z5pOz7LVl9nejxpN7FocxBvHBf5k/NxfV+2dvemWipf/BhYL2cW77OoTkoQb8bX
ImDVOFSXcHPZLSJMQaqFRwAX3gypsYkUmROhs1MqV+rBALCQnMtign7wnOrGQUxL8CXhCz4jQ26x
UpHIyA/4ZMyFRS5AE0MhkEwVTUeUYKsRhBTzLKs1Gl1hwH4Bl7NynkflVuZhvO3Zo03yFJNb7IT6
HuSU7oq6qMg5cLFERbyhwszhInSgDc0b4qPL64GqeZOk9sP/nTraAsGVOPM6pDxvyf1ccKqvj/BX
hXvToEDetJLq88wdxPCfnWRsISuobJOKxCGKEIgsNjNHx5ke2ltbKP28uN0Gj5JYuVEXu5Ws8yZE
k7drmGArtNCOjSVMCFC+MJJ9lGL5SkrpU+k0CLkKv2SR4ZRkPK35OPwOVR5amasQphBAKoTz1lpK
IcyDphZJObfVDW3j9H3+qFLsIsxFFvwMN59vJBNN2Or19Eh6yoDGERHkQEw1WN6nWnBsqD+iczhY
D808sjxRXa6e7goYcin5CLzNV2PXbW3BeuBpQIckr0Np16RnPxLKbLNtU8F0SFQNQbtvmz25lUhv
LYqTDAOEFx8v/K23hmhgmlvcy7JzaOEhrUKzkp83lISVlcZLQvTpas2sJYrCbdmfxAzk66PZ12Xq
qm5sjUTvdK6wCTRoBfUQhwhzjHH8uf+06buPDBjJQqo/fYgVK9vmWhrWXXdvKeZ8V//JsPsdjgZp
Cq2qe8asdVimrU5Y6zxhaxuecLIxafo9hOaxxlS05yV9hHroKVN0VI90jaMljn/mxVMwqW04AjgY
HpTfnQSxWdEiOtWhWZffzIOMdm16GAjw3ZC3h2zOR9jEpDj44I+dpJD4w/mhZftpclA6VOitzbRo
CfbhXGiIMmAjaaKNHRcbjAsz5Ha/X0ULCx2Nkr08eQARlh7kNeJJEdUTRMMWcQAYh2qUe+t4GoFy
tOPmOpXxJgKSTqbbAVeQOXCAgsN6leZPmZ4jHhj5WmrApQKSxQldAokiIwn1Y7/rbpkkXCrYc1sp
bbsuaVHSOjTYUZ2xIOyn44it645SToh2Nw8ojqlekz4MVBCL7eyAh8rTKLgQKslHFkPRrRviZzRy
s4QrrVqdn4eJvJcU/0V/i5srOnIMJnj4VilCoknxYpoACMxZnKNvzRfPFqnPoysjNqXJf5H/n11Z
CTNrYdi6k4MuVgfUF94GVH+gf60dZ0XxilQhvN1/YfpcSIBPiWJSHTPvx+crBogQPNf1ToXBdkHA
rVhEMizdeOJX+Nx1l0R+aYZBlm+7EE0znw3gHVKnhFv7liKTnEzcXjXewh1j7Ig9aXXrt1/AFuo5
nIiIT2se2CC4HL2nK4p+A5vy0S+WA8FLmr2oEkiRVwtCFPkDalwjukW4rpBW+twfF9DB1JIP59+w
DRTd2ffeKlz+ijtt0GPkriGogZhSp9RCfTS/Za6QOLFs/xkB7nfsNLe5atwjwRci83oF9/IKQOgX
bk6VhO/GQJrvBikJt5N5fL01EwbFP5/f9BgeBNtBG9RiCnbBuFEkNz5sNd8X0rmsH6wC3cPmvztU
7Fj2ceyJbDV7N4nU+LmnnAMdCcLS2qEk93mruo6Qp0Ees3nzMfF3+ZN8AQLpkvJyLBoj4Yreki3H
OJ/fLgsJL5o93dUfM40J7si4WjfjodUO/kElJO9dMoEbLEMqQE9Yug/Zj2R7AkVWL54kihCaDkr1
FkHHRmktnSLrpIOatYZ7D8dHL98eSwQQJ0G0n/GMonCYBVSGQSG88Qb9LUlMrBBmHPpu7Q2nd8uw
Fh24no/bob8waIrwnqGSpmQuB7niWLx/FjmJgYGe9aejvH1C6R4C8ECikwV0fTf4EZEbrl/9bEFv
ZPQaxb54JQo5abJ8rAjEafMEBQT6n9GhfA6PEv1A98cEJr3cyYSBNv1viRwUJvf5+/qc8YZy7LuL
xQyGTXfojJHRksPqMOYL3Lrj0pMQrA3HHws=
`protect end_protected

