

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
e5HXux03McEJscFg80ZeuZznrIJptNO1SFQrz1pWkRP7P3QoqpS2mJZRj5k487CXMg1LSvaDqmT2
OL7PFCCTiQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
hgCd2yd1Ey3kW4Xi8EYui71ziVJlfu+yPA/iSZYYtw01d1xCQQbb29qdxk14t+CL2ulbT/AG/Tph
KVRTNfPiGK79TWiKACghNYtvZsEbOSiWp2tzfhZzsTJKt6Q/Tnk5KS0q9lShCg5S46ZxNmKbnoII
YTwtWH6VQAWKrWw0gQI=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
tPm67AAwZoJgqE6aGdH3UBgFSYY0hEjWFTT4t/9DwITm8ODgcytWQbTKxugKHOWkwgxnsfouuhwt
QO5L1ilTy6LqSek7CTlbPwPy4k6tJZltW8YhAKZe6X8IJvIcPyG5jVx+6vlxM+WibCk/roITcPkm
9mxr1ZYPG61/YergLsZha0lMNqW4wq3ID24jQg1utjPuifsU4f5hPPbAaCmkiuYhwkMNuj6VHmIU
m/hi3cIAvUetwb+LazrLlZHRjTpygeOmt1PlMgoOOBXow6h7AJvjUUWQmikWL+0eXLxGX1SKnX5+
Op5qf6RZYmh6jR7nN97PHzmxB7CCeLZXWlS7Bw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
as6iakL3FcmLsNV7kgkV+92olQIBIL1+cbziWnl5Jjo3DH55nMZNZI73AcIS3DfwFYnxJCqB2SLa
SuhR2kAcUXkLjAVN6C44hN7PokTEYbZ0O/DrWDwmWxnool0q47JMJkAhu6l9w278iR2KPAv+EoYt
+JQKH1y1F/+RNrZ1eYU=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
BFKuZqEfqjecGcxpRGmpCDvmWO5m86XHlx1Avi4sYpYvtXIvQdg65YGdV1jpIV3rjwKZHTLGWY/h
WohbbV2nhc+5Ruu6dAeqtH04PeCXz8zphv8vhckLjpwnJT0GWHiaXAcncvq/6wuXR25ASAvhi3Ai
lvDf+vNs8eunn+yE9uSpqndZXDEQrdOREqbbPaHrHScG2A0wHmKCr+QTb2IHKcEfLgWtjt/VCXIv
5krerkdmS143EXlDVZB7mfDSlR6bwswWViVYnH2kDpeepoBCAgyzi+PoFfcxhkn8DGVtdsW89QDd
rLaMLCCjYMVnBfrYxBWw0Bz0mfZcivLyxd+wbg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 18544)
`protect data_block
jsSFhpRRLj353S3HUifcO+ZHmDNk+o3aFfh1U2tcoSGvPa4KKQKNRbngIorUrH7Gm/eL+33cdDVD
BUAPkyyyBTs9yM/qIDF+BDUArMVPJWDpK6Rp/4zfUp6EmTB8CMdTbS/VhwAW2k/ACKwobfCYyCqx
2Wd/NmDWEOviS7N1YNA+rmZr4QeIXdbyNEnVkV45HI8gi1oBg/upRTspnLx2Au2xRieFCKkOkFsQ
h2mV/QdLMAwbAaxzS7gGW3f1IvW2ENarQ0dduOMRYBo87QSe7r9Hs96IrKV5hEUua6DHSddPwqs+
Spaz8PhchcaHrsvZ4jvL1j2zJ+qgKnqIye6LrnLwfbU+OvlRXfpcjnW5L9gnyHzydrpNW3ZecH0K
IcLHKALSSOscB1mxXQfcz1XmCnkU6UHuBkiFTw1E0d39TUHlEi421osIivXHmxjhZI1tYodoHlzP
IhbxlFs7DidjvNDtwPd2Jda5AQwxtQDJsusm/oFoLLFn5n02ZXWcPSBSO8RgeqA0RHwX329rnhtE
Ffyc5yyoTgy/r9DZ5nUGv2SKEhIl5NperE5TbmXw5CiHvGjaFFDBNQA2MIHTshZwddSZ2KWzCVL2
7OGOuBBkz/0/2Gq4J6hJnvI482PkC2XLpstOol+YSpX1t1CLIES8dO1jyadW0m2ADgTcJP9WiDMy
IL54Wrl/eXZmM0FoVT6pc3KbIrLj9PGnrI+NiZ4mQsyRx1zmh4oVw9AhRM2DJ1LSY+/ErMGuU2W9
1cz3XURHMyMq1sLumSteodRgD96/zTz5NCBcPYhuJ90cFnUZZjh9qjSdzK/mch6UN5h5uqWwTs1J
gf9yh494Y9gLAMpaBQubf7afbwxxYDOV4S+9+qtQIu6vPqwSmjD0nXXCSz+RHHwJa8FCA/2l/IZw
Lof7W8ORyXY24tAePbqjaJZDkMBngaTf2MhBEuy8Z3/96/xsmtwWhZrQ8/QJOv3sLncrLohzeEY8
06TZBnfgN206VO0Iqq1kVHg6ONJ7M6n6WZPdjjuF6Ln3JYDFnhJTA6TuKJcttQ7MYx4UCPmSntJn
2+Gyu/OmhsiqS0klytoNa5b0ni+7hxfp89He+FsxKXXOMT+IPpyKawl1wgMlOggcsM3CfL1fW7Sm
rwYmQXaNmH+Nr/h8wQKULcKOrGvWqRAYdLyskPEo1N9vynGgpo79sw4bbsktTQEyKtwRPPxX7/Me
hJlWPaNT29Qj7swot0wvl1n51zC5vNZT5qxsAGh+YJ0k/ngOYyacvtdkW15MvnMk0l0w3mVB/76z
gCP8tDDXwq2tSMHz+Vx4HE9g6ZQMEi7Wdzrav9dqYj167Aq6lSNVu5pYuJ2AktcQMtto14pKm5MC
8W7xiBTqPjP4GONTj88CKgLLkMTQVuC4PYgPe65VIq+REHS5UqWkrumbRNYQy9MP5PLkKNxE4TBk
imBPl1MzsPZZtoDrnly3iCpuvIy6PJ3IDJ1RaJntwJKeweB9fU4ESgeDpM3LR0n/8H1CqIt3EgW4
wRmtX64qZEfnQBJN5nPG4lL/I8Nop4eKvWuwjdLy6/WlCl7+qJtqVRebH2pnSu1SipKpdgdcaqIK
8vEkk8DHhRjMJQ1gy+TQIELESf5RXywQ6pkaGvuqyVS0TnHln73SwRkVCt2+/6+efhnkKde84ZIQ
uztiov2ypvUpwmJlCsCeHmYjfx9euSGMeHHWe2MxTGMFI7g3K8+fUHCFvg55jV+qURi1bON7EfB2
C+NboZ1IL2BisRbagWrgQZa5a2hW4HCMXTYFAu31Q36ogtMlotCI3yC0Rh0Ydoj5iZeuLyMYmq+3
fIQMDKQr9Msa4nvss4Q4GhIfbpoOIT7i0hcreYLKpQ9/4p/qxtApHoG+WVEBD6RAoTHxbYEZrCUy
GwWVF+NTTe41lm2fvZe6Alb5Sg5Ji4fU4Id/NppFMS8grr7xVnmfg+U7SpznxzNAl5ikyAKBoQN1
rqEmSp1UFoZjcJ10gRm0dBMSsKP8gAGi5/wORGu0CBIeOooSMr8EL+1pWojs8exhUE5wfnAhUsEF
sUNv0S33rBX4MVTYuSesS7/bioSKDox6oZruJbTiRjCl91kJ2nnVH0SbwlLWgYdeHzwZKskSiTCF
wEdxIi0SGkj3eGHX7rlsgGDt1neH6GrYoNwBINemDyoiZDLjmbfnNpCVWhYxnHflYXTkcmCdq565
0yMVsv/4zWCkA9gKzp+eGNJC38uxQ6LVfJzy3ReV/XA7UA2fCVNHdZNudW7BhAPbCavC+JVlMfi3
FnDwBarYnVi+BZSnBWV7fr6KwicUfpd+VMpRXu+DXuNDMxrP9EyDmTWVv6VBrfzoxUt52vUecQu2
a/vZs+fjlhP1rJulzLTB9O+DzTszIUluj4v6xO6Sa5BVbNVrPyCWxVahWEF2ZP5vXN3jpqgdYtio
PDMwDK0dME6imlUk0YSv26V52XxAvK24zENyojZnOEln08mm+mS7Q4kkxNoTm0RIT5E3umstP9uH
62iGLgOX/jtpZ5dCffpt8hY+2Ll9SpGXgHajtzNLqvC1g2Kux5mubRatvWWUKewaXa6Xbs0dkRqe
+Wq4uEmSkk8T3Jk/IzKvvWT7jQJkuQcmD8tPfApOpHVh9Z9eSVg4j4CFsShOdUbXZ2accR7mELsj
/w1TdWKub8tLZSQluYiifd8sYq5d/tlx8/i8TMW8qPyhS3wCUHQSu1lge7mS3niWTJ2EQbPH3INm
+vcL+T8Yv6QhqM0cIQm0bvXQgys0oAE2hHwCb0w5eGRJcvHX7NtkpbXH+isK1bV7lOivgUgIbgEr
uAwGk+7GYWAOdOC8K5/yk8QxbaFMMBt+eJxWMLCO3vCBhV44H7H5ch06Tzq79hjEK4BekMX7LGZG
ZKh0h1/FaYpTgSq1dzfhHGofVRlweCXCzXu8X1wRPdSXL5kN3cec0E7gBKGKLko0WBISKWanFoVj
jMR0pMfeqoTCdjU8DJ8T4C1LkcptWsjNw4n1gUxJVWSz35BnxemyK8DNdcBu5mM+u1NDIdAyW5gV
ftzK0PogsamMkOG9ViUeuLiFkno+cIpgwdvorVcQp1II8xZQ3yw6dZQ3CRjNzTsMO0+oK2NCFwwx
L+sPPU4rHrHNskC0gJTg+DMjzfMIbfsCUJSsaMPunyo7LQ3NcJJ/z70N5MFNUOKybj5TGSyK0nEU
eB8nxgY2E7Zk9SkTvMnGqGum+Cht9EOvokM3Rj5nFL72srU+jShnOS+yRZ7/l+/vUlsKDFLNqtld
S/+8EAtoy9AJn4YLuvnvDD/tY+2CXcd23maqtBnfgb+N1H2DnNYbU92PYSWXThhRHLa2ZDnJMTWJ
J65JNX4zWsbCgv3XCnKDKqXx9f3FnAjmhlHihQt/rHMKpMqceqvIXMxVi4ANzKbPxTTW0bJWZ1zf
yGqfOOKDmfUn3DONGZ6drLaD6l7SCf5lb6ddZcxmSxwKSAtNAagH2E7FDQMpPn18rN3bLMAm8Lic
PT0tit7b5iMstZvnQY220j39m23/Ni3s+8MIPMgCocNE70J8RIk1UwIxOsuBOwOP7OfWCMqCeFYG
84Dmcuf7dcP6Y4505uKV3Lx/p+2V6kwTxtZa1eatMWE5t36SV2bx4kzIEKf1MmsPnkP+2J9/uC9P
mw/Zywhr7i0erSo1lZoh2ItCyB3LQ3XkZUZINZlcrZCbMpoDUPTZHVZXiHBHhW6FHSKmAvAe1S5G
wt9Qq/ymcRWCBRAfumjEhT9A1xoDwkzTGP6DYXw/osH1+fCB2bjREFe1cAkjEHHy0OWzlUD4iiVA
k+2I63nh27foTpI8Stz7m1Be6GEeb6s+KMQzA0XapHb1NpuBxy10oPOqp7VtHrNFtOgS3p8+g+Gm
5lrjkpu3LP3NcEHlI08wyytoRrN0537d+fbMOEBa/gNqtpYtwnXhZKo4qMCfhnWES3ZvyLLM7v85
xbXFiQbcd84t/byQbt64qmKYvWAhAAdpCjz5XH2Ki5HRsB++YKibcRywrQRGI015Zv4xw7EuDLzB
hHkLcztXMXSOBoJGSVS5JKk09F79FvtKlWcVIZOvJwnIMmt2+iHL9z0MIuyNp0Y1WA54D8W3jhiN
19WKqeC20ww5akwEUBKjmNwGJm+nZCFeGEiO4zGeeY4jLSakgG+Ih2f2wDoQMXxbLIUIupLAlP6G
Q9JpPFlijnms5GXtLWTL4Ni5jVOJk33ePMddwhXnGf4qwebFskz9JZFKI87ZsAeAApUjRRYwQmXZ
pKz84+gae54F24hZurpVU+0ip/iCJB05xZ2nIGS7lnv1nAz7rFahTRYWStSMjRaun6+qtKMESzH6
I5j/uJLN+rfThORHyEydQsnB+JPXR+GcFG2xYnxX7mkv1xP02kVfh6kc4u3sSyE/NE42jYY0VKnz
bdowJI0bUuNqhwO5nVDm7ZmjO4M4PEdEDYCP3m1RrQHKB3Y8fluIQK2kKbgsYq+jx/+06w4v2yEd
fhVvKRfX4RGuGRz6uLjKSykHpFfWyQzGJb8ZzccDBiKTyn2OcggXB1/dmizJ8GKUdnJ0z3+mZrlE
t5Qp3G7S66ExrHbxaQYdIAB6PEfqvz2Lp8xjawRuCKSkOcdGSNEZss2NhPBdF6tOZBhsyRuWN2g0
PXT6wdB8hPl/UIUXDtAcsbMWzNGLF0s3ysgl/kJ/ukApxPswVFZeE7nlBgtYof5SrZcWiCr9jsS/
8RJRFSUafjOsa0JNcGYF2tEJxpukjRT3HvShqpoJnDSqX3KePSxWlIUZohZ9dFR4dOWFMhEJWiA/
j3h1i4CDNsX0GPBlIRjtv7T7cYGW4HnA5tTG8GBBh2iwyYPyCTxSvWp48i6uOi/ofgfPYu+b4Vj1
OcY6XUovfJ/rxKXpvHRPk+Q1UOWBp+S0XuO7c3ZCRdgT5TNcc22s8MpkThQwSbIpyOQJQq6O3eIL
KAEUKEQtOTaeCJMYJHrmiq73uHhg3Y9yalVh43QLQSp/IRQH81s2Kul54RRwTuLy6DnKmzX/7UX9
/vQENNrk/Tux8/gYXsGEhpmIkVxULGq1cDC4lkZqXymAr0ZKhHm2KswEmhZKnBQ7HwCpB8/cVhTt
pMtN03jA48AdW2zfWNc0OFoTy6F50/kBs38tuhC7RBuWHHnH/PpNTTru0wp9ySBEkr9O4u/cJDfG
00PAB+h0luvw/2aKYmsart1IMexZMePSaGmhq+DTP0aEh6LOl9F0GUwYzLz3C0he85pMo+kh6h2G
rKpF/1lRFOyO3G2un6LvKDK0xD9Zq5lRQnYOrNi8XcwvZPGiCLWGczDoBaiJxksjaIrgGiK8j2ua
kn4+U1ZP19C77hJx2hCrd5/Ltez4QAKR5sZgeaJAVg/Phwz+Dpb2n+L1gPnCMIO2RZuXwGQkJq7c
ooQTKHeaM/OvqXY8F2AtiHV/hCk2VklbSlis2B008ow2uxJq8HAn31D440SCVW1XZrpq89schmej
qIxpoOE5+R7+aOjkerryUcEcfHltXbR+y7vuUFJ5HZYk+sFq6BjM5wxCVJplX0J6YQuu3ftP6tsi
3zdF7R8LBrASInYEvhn0B/MIKc31t2ORthF1/79CA/cAnwKU87bPJHaPSjisfCNmvk4dLkKf5e+g
cphd3cSmitlJhEir4jTu0rksboG8I7wHHfNmt4UPbf6Qa/X7q07MW9Tua/HnObBzNqeuacaJQKcn
caTI1/XT6fpmrBF9OaxCdj4burkO+qgRa8vYb/FgFMO2Un6zyDyGf5F5VCtUYaKD4aWEACiKx5Dp
auITkRn6pFg8uxG6Y5hgjp1VcS+PqBtby2Vx7HUQ6+aoFWOLUYWFgTrH/jrCUd7YdpGDB+bV/HNP
FoV/M/nY/SYElN3JKD31Nrr55LljPPFS9WK1Iho2XHFbXFv2pAUdqbkE12Bv+nUFn406D+FMqGt7
M9cDMyDfVtviiRqyNXiKk7jtBgLi5iPGL+xR78O0UCJw9KY/SPiz+u6omdeGtuio2N9yXBid4aiP
D4ppB+SCt5Xwlma+FLjlT4OoULrpQqghUpOBPqSmu+SEzmUs46llAJPbu/8xWyv7gviy7f7FC01E
wWxQbXYdJJ6RvaLpUtehFnyNNvBPhXvkMMWWIwBQgApf8Bxe2Sa12Ng4k38puxXh9TXefkZt0ufz
KQeihgEnq/nCdLR8e5kxSKQYZ4ScbcIjiZLxQMFyYoDBm5dF7QLKMKzOsQL5uiibf9L+lIMsXVYh
YlVGL0Sd6GleDr9lLqCnosEiTfQSCjdhmDy5Wy1Nra2oIlvSjH/MgM3lpUUKJX1sgKI41/vG0LPm
c4T5istqEZ/N4dc/9FJSw7Ihy6u9JspoiuWGb3coSE2AFJa9KqjAgI4rKsWlXDXeG10XNDQGcuux
pMIZg0LcXEHbxE1M9t/uXE/p8joHdHH8Fpsz9J+ztnfi0qZSczeqSrQx8B/UnPGsq5mqjDz7kGbd
NqgCuOCQrs96om4CE1xDdhOIr/V8CPOyAyNxGdhee6NOtI1ZwshjpS0/K9+IEYNa4PL8J6WOq1uZ
Yj5FO2twzIq/FMnDJ9AHFclaFLReC7S1aB1a3ZY1GirXZRQQqreQkjwVPN4QmLcGYkiRvzjzqcby
BSglAwqO2nskGAqOkdwzr00oHjrVk52Ya0B0gLqa+FOAcGH2bp6cZkydOIutWD47D0fQqcyqe4mf
prWLzTvEsNjK/2Xu0onTwU8Q17zwM8nRRRm8lX6dT4E3qTS0NomMHAnY56LHWk3K7XwPdZfawKD7
SzyAPHppGt9ouLJC7O/MHEb6SQsNj6zfppbTBOw8J1h1eYoU8MG6wFQOYtPSBiptsfSv/+8bfTJW
CeldCLR+FLoWNwHdWNHWFnmx+VYp8Z4DXm+Sd0CvyGrask84BWS/NqT3wV5CIfM4Efjx1QjiS+8v
Bz1Yz2mmyAJIJR7N1VRAaTsKstkmKOhz3dYBxz4yW/0XAIDSjQMsfr+nQ/keQ1IkFphQhovyTa82
XhppPYjwiu6OthlLmj6lo5PFsqJxB6JcAjfSNYAWg817+j0Vrd4dvcUv6l56HuNOBowdsR36gmgl
x7iR5qboXfSsRNpV5ut1bXH1ANvXzwQu+Cnfon6Ia441rfW6qP/cwWt/OXuEXNFmYeNjhhCC5nV+
c1t0MlR1ihvw9UuzQ9LZbAvVV8Paz34iFpfNbU4GomB6KH3+a/pcJwvWKRl9x1PLJc60YxzRx2WE
WerU2Ag5umxq+cwa0qauCIR2mV1UH2RUiaPfBJDyjmc/H2V1r4oaNkR8lBfSTXUx5wl2eLDkys+5
YuBWq9vBMVJlX7dmgBHLuNVJ39uYMmotLUsdeii0V3O4CvcXC1vS64aMPTz4Dc4GgQdNLTw/X3dy
D4kEqtxeOETOwIxEFbrYZwFCYv63l1jOUGQx5dcPKUwpoZGxi0JivE08wO903B9UueOWSh8uxi8K
UcjZnZ1BndGHYaD30kov4STuuYa8oUmJLcT8acbepPrBg25t+LNgy9MFp3xxYzjtkT/78Eq+Sab/
BLpTh2jAsiaDUmKXFgJPW94BQTrKP5IUzd3CjWxjbBKhlJiaTANjfaJgWJnHDPL5HpDuBJmQ19DM
6N7b5R2DKHTha2kmz6OI6QR30y2odTBncEQkYhbnMDRB6UZxlNyMJxbGbPPFfnka0vR35TErIaHD
Gc1vgo83lXuKb39plzNEE+4yMf5l2NT2R36s3g/pjBcnFDmmfxBQKOG5wBaryO6GVGf4MBMTVU8G
kJS5LsxyuWbihbDNAqiZRjM4oFznlg2Edm65CCKBPLyZ3EXpVqKgvC1DiJubFNv8PEe0nuODGyJA
uiJXT80X7f5aOYmwK+JAjmX0DKx9W/OsaYRvOKfr8hmsG1B4ZNbF0XxTbpeKeuOgoxMULH0hbjAy
suJpUHWtqobRPfO/T79E4H4lJp+VtG/AvTUWlS+c2wcg9T2fZPinUOhoH6hiS0wGJ8TOKa1fuqe3
2oNYsbPrhwcPeJfQGxO0k2BksIuO36DQ7REf++OzkqCzX42tkIoS92ydsmCLr8MefqwdELsa1cZg
slC7HAzDfcNh9dplEGhXepqcIlgK9lP5fk9qUH9CEs4HLhkDAxs1WKnzo+4bga3trEqG6mIh1wav
zgQYGQdxhUU+a3XFftBWwF2OYv9e6xogEgxrMx/kqYG7izXTXdoUUsaxDYVBMssnkQitcYAhSa8M
3B6zSdJ9M7AghAGjaa5FPxEC16op/6ZK39Orra83oR0YXwm4RCLWL14wizf6NsjnyQOXkyXHHk02
A2J+dOaD1DvRzjTi+c6qjiwiExK/vOKYH5d/cyH0rbANwLO51QTUerqFCEnHfMb3UPj+Mz7qfXGy
eem/gJ36/IsRQHy5mtX+EawdaIYvOoX7ndsejdOE5pPcluMrnbPeC0Sigw+XX7qtVLP5b4SUuuhN
7SmMm9WNjPRyGIt/l7dS+OEXfAC7uq3To1FTxUG+Nn8Kr6g8i4nmQwNGT/lIio/UZGABKrRlKc5P
z/HzRJefOaVqiZd2e1tVKN+3p3uOqfzQ7SCrIgEop+zVXoptpJwmpWVst28sQGFxyovs0HqleJyU
oT9YKYVC4t1+uVeUtGWz32QLLH5uhrliqA19YrnS1gNGJNFnR0L4jV0bAmsrjb+2wQCivL60w2mv
82TIq7UPYOBM+zQhNivmK3zXPT5G4bMseEEtvJGpsvg3oG5fAsDwlEwjc8P9eZf/rvhlJ06pNKeK
gMZfBITw13XssCxXr82g2faJCh+VjerEgLCEmAGbRzBjMmtTPrzvdf1rHPdOroVMlAljjANSu3N5
OCGagcmLldV8/DaginZSvv0ciDv49CQUQvelzbN3iu1vBqZg9HSLH43iLAlNxuA5OchGU9XP5iOq
SUCOJhb4w9eUwLJF+XEomt4QISr55FkIjctzHFRBPy7nbEyf5cVmJeTLDpK3jHIWvKpL67aPEdjh
JHrHFu7Z784R8FjDw3hbZL7s69quiFsNCuIm4mqgeFa1dM0plkgGgRVCRm8NAJqzxN6GDnoy5vEG
eEaqVVdCFYv0VwMsjnD173feUf8gOiLLuF9dwNTc7dxLuDVyG0cR8JWQX0zeN8E03zRDmii7V7xB
bkfkEjzzji0+EYuM1fBSM1eJZH09SmjMEjw94kUFg7EtdIJi2VERG1wKuQQoJ7NDfj0oRg5zcTMp
MMzSrdM5P3UxtnDN95cX2K7rU4XV+xTL1r67TUY6o21r4v/r3dL7eZ0xjAEOejKItsqeyq4f/7Jh
w22/Hco6a4KHDPBUo6escSvroGlOjjPDPuiqCZ+t4VqQF5tHuZtxsPjPVQKq+UuMzUBNNYn/oY4c
0KM00vGOHnsMHBOe/NOXjUZi1FVGywuTwiyx/kjPaeMqrhkn9BtlUIS4WBzk+6qY9mGQY7Q/J1aE
BVFG90a4PX23HUtml4QCCAG1dDsQfHDZ/II8dXq4JpLqBc+W6rYhym21ECBl1854118bUsUPk+ju
6p8KIfbAYuVxSKewLG49guyzCbBhZJ1KhNuMvaD9frAGgMs9X0JfUSq/rNW0vMOET58DvR+rLccn
fiqKd7x7KWhiQx+bJploj4rTedKsmpXPzVE+mKeXp8pUit00Utz0Swc/xEfMegKNlxI1eIBD/SyZ
OtB8R/HtFD34sn0UYgMlpiBZciO/hT5jsGGURE4d78R2wZBqnialwDOee/4DXPiRiCk7nrFaJoH2
MukyW3PalivO6zQFeLEvZaGTRpdv7Ey/ZwSWNbT6R6OU5QR7UStbbKyoN5qvb6EtULopkZV4GJw9
mGBZGE9udvLSGCb8sh2ylIuXRysBnqlDrZF87BR7tAU75VvVsN1HiEkmUrPhc49MG+lI2HyrpdQf
1dodtXANm0R7vIwZdUA7avfMsnkNQ3UQTIdGhbX58k7MeYkk6SaFRFzkHgz1uQPGRi9TUHVFRjGh
BN+d5Hbv2T+93XwdFgGPVUSCzvQ4+4rjlh9yjwnhyntw5t7v4DI/MOpVYfHzTu+WoAfjSUjZSaFe
ILdjBDiVwNLuWYZQVM5/iBIpvRRo2vtig+UbGHYdH2TQv+L02PlDeKWx4XcUQ4ElfD7D/kSu+P8f
fnRKI5DG0vmndNBKtp4zlledFxcwe0sdqtnt3VJzTeI70Wow4C588H1QawsJ0sr6ru1EFlxCqi0/
JYUWyY35APaHaJfCLRdcvIZZWBPocGTdgQ/o3ZxcqQ8pUcVWbskx90F/ACUYrj2HczgHS+rO8WVB
xJxAmagj8N1/dHNC7LInW+SRSSmONXd1VtAwiJ/sfRGLGpbUdxniz9a73LgI0FS2b5gDA8Wv8iZZ
wTj4mWkXZRVZgoLHTUplArOBkILCzDCkL38z/LKNFBjcY5xLkepESUde9fOMPXNz9tNH2HfCvjZD
AoyqBUg+ErWOgRXGxgX8U99aMzfxYp4UDKweqLyG28HSNp43h/PcTJV4gLksy7WMmnm4hr0B1/2f
wLXxJuOvxRUq97LzZSGLWkA/CjusRSNwjcyfQzSHizq5CeG6G792oEwS9Y2Xpz5tnQXPQOrTh9u5
h+oI6AhOqlyLI4vhyFWANvATthXIUTD280HC8RST8hpNle6mDbGvRfaB0jXNKPqU7kcLDkUqRy9+
CrttLUX9tS4e1m1WF2MdurTbScpHxIx2KyMQ5cKQOprBvOJS2FI6V6JY2L5nhbjP11R056aFGN9K
LB2HDKoaW+/6T/KofZBWOHWxYWlccx/PUmSllGHxzJcCf5psYGgv0UTza3az5GQqDrC8qPA38Xh7
pDW8zbxleq3aAb96ParqyHs+zxjExBJLdavo6uGEvVlLTO9NYxfGPcrctGA9g/OUbHXmK8ArVVC/
+P03CR1ZrPkSlf6ZHAAcAJFcg2UlSFZtuIPSB5xCkE34trFWjwjH64NQFtDRCgzNaOjTq4w5toxh
IhAAByp/ivLI65vygAT5pEnu/tzhiHqOAvQv3srblAY84PpDc8ExMIlmzeBOQjYnsVbF0e5jZkOm
KqsQL+NCOVm2ENL/uAS9SoP28+0Z8q72PKFhv8dFWsMRGvU/PZm21wEzEC5L1ZK9RCsA2633YELm
jQ1MNR8VvId7Zn+cU2TznM164T87aDzMQp3QQb04Y460HompBfLafGxDX0UEtOuwSt292EKKeQu1
nLzYF2yn2b+nig04EEdbuyIPUixgcQlv+UwTTqAHSnO/2MKNGk3CRSyUde42RnnVykmoKJ4GR2YV
R7E6gE3140ZF0/mpW6o10LfYSTMYQqUr3ttamsOoqwsLyZCJTEl0lILN88hMq/GfWqGFei5+oncr
FPUcdMNZ/B/oRXEMW7eISsxdVM2DhQhMxxkJC1of3RfiH8WeEnpdiYhSPTAjeQiROG5mI5upcy56
IPTm76Qd11VIw4sYi+LNxSjpVqYVSYnUS1Fg4oIlB6EWb8o48mCZfeuLhs92G91ce6/fgcIsBVlU
ac/WY91FkIVTZhJCvmx3ph10XYW9pc2olrGmaLRLxcZ5TNtnP/p+orWodFY9QAyhNHLTdBzFVWBp
GbB44ZAFxj689CA2jcwmNay4Bm3Y24HTc3SpBKcTcNeNfdlExXiYPleuipBhUiWHzP3M/nqHVT2k
V7qVr2xXGDSazUem7lwlCDDBLly6ia0iuda29uZjNj0+jpC5IIOSMFGJRcoLmiFmBiJzDTUobv0y
4tH3SIygrL4PdvkfbtUm2cDFFpkttiAMNM9LoImW9hLDbGpJ9c0ERRHWjJcIKmPmCDasOGHNBEKu
Hzd2jCROZ+qLU+PKottiRLSqkEItifw4D7uTaunGgLySHllzRMIjYewSUZPJyS1qMTcL2eEELktu
om5CvA5snJFGc9pcTtY/jwWhYyNK+RzaEPU2BHAcAygwGs5t/tqNUVp1yJo8hcexa6DdCbbw8hnQ
w4se0lXYiztw8i+vUd/aIv9jEqHKeebpjn1mILY2Y5hQbcGhTHK/peRJD6YSggTvEoN3i6pTteuD
9qCdeEEzLz/M9mhkN/Iu0qtGRt01VA10BLv9hl3WlPjT9Jj7bey62+9Fiw9WIRqTE7pVQxHLRqTM
YLbxngftcxxbQZJSbhGBtjIPwyKAtGFg8N4sCPDLn/19eCYLsiBURKq98l/jvZjn4EBWDFZuDdMa
JbHoXCL9iBvzKPQ/kwmb3AVICZ14NDfhIW6apgpVAEEvbN+evNpJ9wY8CAhaba1V7CCniUBktQoU
ca4TEgODomtdMPZnCvg2aWyzu7+UrXgDAqrhQBjaO6BCrIWYmIqxL9jJMMjcE2wvXTw7hACIgnSB
jtsPNqEormBEgjdEqpcmQWSge5xQ7drekj9f3Gg3x9GK+ulqx7AXhQZyHWSNxl1jn2k4Hz6xgatJ
e9mPjZ8X5Ti1Wdcdlon/GFH34jh3jue+QEnUY+Iwt3vDQB8If72fJQvKaFMWp6ORXr7SnhSvJKpJ
YYCrjufWD/fp92G/GW6Xy2dKMQQ7Oq6rpDPVTq2ax9m7SQs92PfqSA77E/sChtCxYTqG4jNTdi4Q
+8OtXGL9veiJMHqnRCgK1YlM9973Z84A5U1OGYFP1e6hHk/4ZlVa9HORr9kMVZx7HQ3aGvVanw0X
EeCXmjd7Ujl8uW77lJ01iWUKmyUblhKtZVuDHhvKdGb4PfrPlS4NpjxNOs+VS2L4DqfWIjACuLT/
A7tQti30yj3XL6KCI4EAR249tR9nLWn2aSsRVtmEacOLFCOJpaRH+3NPKTxmUNkBooQ6BqLXT4vl
l/9tN6DLOaimSY9DE31X0m+9tNwQIjdNCXlIErqpU0kDFcKXahRXJBDr1KiwQpyzaxfKifckLU9s
TtGSApLLk7XNT3G9p5S/opf+fKllMmUqOet7PTvQD+Ux+gHUB6LERrHb+XuiYU6TJQLqZSLQoCQp
EOFF/cuFRecFB8aZb2d4yAOhwAsp2DtevVqlLyWfuxX4DfG5jiH6k8wfgh7d4+IUks1ZK0NTxg0u
jdCDJi2Thqfq204x10OZWL8fl6xRdkkXMrE7XJMAI+QuoWyDGX6PAD6vocR5hqMLbcdfB+GrS09S
ksm4AtfYb7pZDXmocW3y8dtnMe3DMaN6lKVw6vHw2tMB5s5EBEb6fOXD7BM10WXiNWbbJw8GrDJK
cC3Cz2jRJmz1ICmfoBE4dO+OrOevLSrXO14hqHgAPZXRDMMVVCbK5/jwa5XOXB0pFYWLtXcmfYHW
QMWE8u7f1TfnfiJQihWg+Qb1FmyIudn+J8rL/cUkX/N76q23BPekQ0sLNpfK5gXfqn4RYJLB5bGR
4zsv9R2fFAVfPEnzSv5aLhew0UFaIu0Z06JwG6TuwVnTRCS3QfV7o2Uj7WHWzatmbQ3IDYoldRmA
DIHJvkOFso+LFOqyyb4vIA2maUY3LPlAWtJYsnjLmBL//XnmW+vkdMHNsY2KAnfrkMeUEFqte9x+
Ba6aBNzbdEvnanvlBpSaVemS857gOHAPnwGLGx3CiqVrHeMy03xyt8lJ/Gnqiw1OFQBAw/PA+7qz
OBwiikez+h6JAVaakmF87RcNzB50UMVdLeiORQSyj5ZOdCBb9SI8BoD6GqzcnZkoj8sDNoVChmiG
oggIXAUEnNtX4U7WzaJMPeGJ152R9g4zdtzPfFPecyeOVbfUxd3546JqOe6RgXhy5hP7HHHeJvt9
2GM4gqF19Cw70sJqUEX9HvvGLg75UQFt+ozb9uoxAvLtON6LkwG+7AIiWaIbyFWVxw/nJMkqwFvY
2iyQkxgOd5rxYcg1x1jopSnGltVx4KeqwBRrKbwx9EsdeJoFaQOc6Vv+8zF/tAqlsbPnapYU2erT
RWOaVRhrLLqMoOOu/1guzO4OexImF1ir6+R7OlPP3snTrv8Ctzbnt+EL5OuoeVYDXy9XG1oQTsGg
nl8iUysOuqtUdNR/hzCLRWrKMZgrnMgLU0c7EGPxxasH7lRaBTzNMK5KccpcGUse6msd9XfJNkKe
QLmPSccOe0VKZV34q8yl4kksLzH3dAwvGW8S91QfEtLlVGkhBCFc2QieUsEWQ2v/1S+x4Fs6kxC0
lCLNftz267QLXtr4xsJdL6ipGlXpBVlkA/0AxaZW4o3YU4G20OWAa052nJ5cRIkSbQhEwGqWsN/j
F1+lMa4qgdzxVDZPPd3KDxux+3POzrpuBz0r2QA/iWqiwtEVpow8kwzim99tMWDxbvjcarSLB+G+
8dewFMkO0JUfRh4to0dYKWX7aNsRHRoMtis6UIUwYvhm4Kop7WbmuKCLlfcdzZ9mDIykpd8tNIWq
b/GKRdmcM48vZ+XpYIBDksMXfnnqdjSWWNDfQCsCENGoj8yKqYev666JpMCzBfRLAoV+0PPZIyt6
UfGcZKYjGlhWBjsIaOl3eJGfrMsjhd14dDzIzgMG2r8cpFuPnEM6AEIn04qK2eR72v8iBGR9mx6J
QvJR/Z+W+LcY59xszgL/5uytS57epUaVDKASluN+YktMcoHkcURPxbCqarxntYj2DMmkBJG2TUC2
TTYKCrhRuc97MUsgjS08KYClv8XwBHVNxOrOgid126K4xWiBeJ6KJsY8EUIGGOYmFYHU7oXuUp4S
nAUK0sTUhz7PQSXiNOcvSZGUU29Cs7HPVAwDwFPtKk3GM8Q3DY1y4JdEG2oIRYK3uS6JH8ecN+lv
vyZdQtqGXTwDDlse+RIR9HkF80+7Ksb0xBHhpO+2E/40wnVLuao60G+9e2uuIxBE0a310vu3gK+L
sm/xp+94ffHqRpUMG6WCe45RdUZwDuP0xlgcywKSLwqpfhVzqOQNLZ5l9fRbKeGXKakcsghUcnuL
9OEcfpgHok7PiZyGxQ39vEirgAf6drt6ZsR1kzlRZUTOZynrhcQnAYprUdRp0WioZObEUA0F66+s
29giNcaxULtkakcBFs49zmO+Gx8zDeEs/5mIojsKpJajpqX5h7g2z0nULBNCytHzEwEwbMrY6n4W
Gu+tGv6OWo4B5LoFUJq+QiMzWqIw2YDJjWEF1XeQJcUg5O5eCqd+87NgtTfXbKI9+jl1YU7Agkca
+Ts6jiAM+Z9x/g1YPtA4YSArJvIH5JnFe2KQQGwFRuRUyFik/OtuCVcNacj2kvcKpTNhN5+K1Bh7
3T9lTU1/BvQthDNWUpBITvm6XQoxvasAfN51mAJnuv8aVkv/l1T8swbqRvVy2HvxbofgBzGyK9CQ
kSWG7Letg3l4q6YAiguYMF59rYLxKHTVBwLnhsYzzNV32vIcse7IKJriGHV9gHxCK1cGwGsd0Fiy
cCpgWE8LUIeEU3GUq7pRVEAmTJxGAAONnss0K2wb8chNdL6bcBlA7T/uZGJLGzi9EHes+iDbC+Nl
G9YBkdFBO6DOb4PWxBCRAPEcR86jTyv2nZTdt50Tg4CsLerL+RI/diq/xZWN6/NNBuz3KoZAaYGA
2txN3KarcUSSci81UN0xlJe/k1AAE/IFhn91O57T2HueMpko5StoQ50mCkVYaEPernSLNK+jUJid
KHTfGEyVy2xPWa8DgcBo0kAbIUYWyzheWPj2ytmqKBsDDcxPZHl9nVFnEKBjb+ZQH0L0ZGHp98t9
SknP1hnSwBn/MJGY49E65aLONiBB5TURnaAmVbRQm9b6N/yOXBTtbkZdEq87yTqHoCF5B0NJ6hDu
cslO5oIdVSBKb60tjVD4BQk5AP/OxDIuJ90HdI4nOZBvRiMPrDkdNtT9htjNnJju+hQzbH8Db8LU
LJZsWMz3KaCa3pkseGcwpif+L0rox/6XayKa/6wJxmyWQBmGP0DkIsc3ZxBGkoxO+Mf30lHMqoyZ
89rw20zvInar702u3RZNgGJKT/FjLl4VnSpYJo+JPr+RGkxoBF2TEd1sDQvxSUZU08av4D3eqCyl
R01Lx5viBIDOrPm0WDloP6fMWMiR2QIK1EFW/4TVFi5OuJFgERF3SpWbst1YwezL3mfZ8y19a8Me
0z30+eb3JslFgiXsZ7KteC59DlP+j/PgIxf9oAYn9MxxV7bJMIMAkv72Gu+xx+MGTzk31Zg/5smk
YXY7+F8RbJQ+eUvpKv4BuyUDstOO5cxM8UYtRETF4y4P0vY6HORfFjW0YMZF4VzKkGbkBf5FdSV7
CYNhGM4LNkd8cKwAbK6zkZULNYUoNX5BFxdq5rMG8OFy8QzJ+1+pWPvcJUKBrUefmA3DQEbOpU0L
odUkRer5CIzGt3Q/7VHqmaKuVqAwEa1TBCoCvQ+aGv7nzfX5ogOlkIkXAoCtLBbIbADQlIdOspdM
wNyUyAKQFp6U/ptOgg+R6Lvdk0ZOM6a7zNKCqB2tEPBRPrcHJ7ixt7WY+I0qMP8hc+0CWKohjqoH
oKqteVZ2cziwzPRtB4+HvmK4C4314v7y3VZ9vEn7q4VgReSDgNYvb+YdSu6xrLOn/+Je+RbVRCJY
ovy0NJc3gsctIIT6z178okwK/vT4ZEakBWTXH4MVwhQrbuEYWAcSUSdtVDHEjwFzf2/6Y10d0acu
RmhWhrUz4//Pp6ZJZsOY7hBmvgV2C5iFFyK1p9oADc/l/8M5Zj6MQ8VDBHzAVGakqgEIE57w43CK
mcy6PMMe1NmoxQYRbGjtMf9l3mshkXilqRnhyJVp8jzVUnlGeo1bpUt9txz6pJ7iZS03NasipTEp
CZ49i8YRLxL0QWGet1OgMm/qedxb3kIvvpMRVKDpLyZEhqjBKwpojN31/FUE/xgrMtT8VUvgiAoh
ZMXLbRjH/R6PqmuDAjgvy/XJfkYSWiGo2aejveJKhGAJKO/7yG9f2ncfeZhPEUsplHLWyY9OnZnd
75HH4uITEadY74hUbAhsJWkI6DvgeQHJKZDqEqQG8OjW21ae2uDHFvipc8QxUNEfX1VQOW0yXU6+
4uqjSP5LcG+NcnmB2OiJPH2KNgiEEMOVg046ZAmpJ96AqM5Ched06jVrHKjtuQdDXdxMGtm31fw7
Iv12VJTjel14ZBRc95aqchRUiZh29VrX6nYwXGVetBQHYGJmgN7jX3ypFqxVaTBZhz5ikC8irPJM
QOz+wreyZvib1513SV4Updk6f7bi5dje4SZRNnLcH/kC1y+JGNIpT2TwpjDStU/tPhpTK+rHPnwC
oS04OfEQ5YcbVDQrtPVBQPn3GjqtMg0OOaOd0ruxsJwPfyqgF+EMO/cKzGzZSJo1F3Cqsg1T7oVA
8i1g7bhIQKEUztEuAKVOFx6q7KrVSyOpp8DD1+A4uBow3rbQuhgIIq/zyPtz/GI1FOoIdpaTBoqs
Us1q4ep50O5+TY4i3ffVfBeP4V+xeLtUES8rtHg51VJGWQhzE3NrJctPo7jkwIj16ViqPLUgE9G4
NlNw9LW4we0AG/Yxx1V4d90w/enBDNhiF0XcXXEYjzaN8SIHKhOaFYvMBPhaKerS1ht9MeGF3SEb
vzJoV7U6PLNhXEHlxbTng/tcakBNtnhKWet/AXQJk2tOVzZS5X6vWshYFW3Y2dE6eOSntmwWp1AA
pZ1UUKUu9fwnWgcUGwenYBfRho9PJq4O+JJyXaRzfqq6HCJnTNsguCNR4C7gLKBKDEU0cN1BCMJE
XIwQvk+c7RI+1SM+tUQSw6mGXdBpJYAoMwDGGJenBxtrrvh0o0NLQl1j/ffFObmIGAyDmBqSby9T
Jbjk+gsyo7N0Ek9SJqDIOKQgudqupqilV6RKE5gQcW+vmGB7cYOv1/yoqiAZ7zyU4rZ5zlKL8kDi
Z51I1s5hN6fygfnLkdDv6t8uKnNs9Fd7ezqUvyUIko320pTSqUJfsOpXuVF+0BWQoAhPJG0EEhGc
UXcDeMDV5b7VmtsShDYwiBbRUiaeDDOvNSsZNlbbXO8guQDgx2w6hnTlBcL3IPgkSLJbBmPHiw5b
vD6p3ta5RxAuOSsSltX+RvG4ZaELnUcIGoQoyZApoCpw+2mHJpxUaNVvBrPjAyAiawjCqO9KOXoa
ZyPHpwP0EzSGJjO3fy9LaE2DgUPXfVWfPFZvK5Jauv1jsJkxNldOBV3+1Nki98YQe1lZbsnOvCZ0
E0O4Cfj3MMDlY9J50mEZ0HegyelqYomrkpFLhVGROhfHKbt0zprJYrW85SBnSQQ2KNtlkxpTwcBK
VLrUMVjYr+qtzlbdMZDywNKS7MqnBEa9SxEOMKXtMl/+fRLOdkU1fjekq4DHwEdcrChkesACcbB5
Naun/QY2ToBwPeGck8LonSf9k43F/I+glZswWLIBk5th6ZF/oMupQKNmJbgiG0uNLZDH5xrTXENf
rnikEf2x/H2GWwdtge1zVaTbrxTlQkVz1xY7Uyq+OB6gWz/g3QZFX82O/7oc4Nu+zveZM+B1jWbP
jzHJLs2SZf2VIiOksXndOOpcPJrGAmmxNt9i6sxgb2h922Xp8iSbbHAT2qWYxgyBC40sSo6atmr4
M1qHBWoGvJtr7hmm6ew+8cc17zcrR+ttiHAH3+U1GoWMw+edrsOzrv5jKovFttb0hWvnFXV9riFm
mnKlpmeHWp/pTBwELeZ2ACvMmrs6MLLEuuQnTPETbzOWYYajwl3sTsPRKQ8TPRTsbbq4Az30dxI4
XoHJm9xCkFaxc8GavY7KDiAZ/pkXAXdZaiBfEbB0SYktINaDnQspy8r+rYOBs4pEwBS6fxH/13Oj
cSp2wuBJZqMLOtdAoo5tqiMuQBvN3CAwvMOTfb8g4GLjXKM7muZz2252+lzBgfNex3S83hTqDu5m
T3Vew7Na6R9KuWaJKjkGoAccOfChyq0suSSwO28J8FE7gQ0Bv/q1GzlGL5Ny2cwmvVpbhBOvIOJu
axOKOLvE07QFvWEpNsWN03Pmx5naGGeXaJ3gwF+d9uubhmOOsfZQUGJybkIRNtSmCb6RmwAVOILH
2XLt08kWXfVcu5FgguyWpk9qaSorwn6R09noYEf1RYtm3bfbfr9sAal2M1QirLSNeQod+os/z1e3
eN9O+EPqDj9yuxpvwTG/BwTdvOkyR9lgVlGZ9FYy3fshtizmkLIE9foOwfY1wwgs9LEaQ8WzR5P8
uWmPHUKQDdYY8yoLdxMED3V/5EI7tBqMC8jF8m/MOlYY5Lj4omkxWUeIoAaf71L3im3vHsSC1wvB
uP7BarzXiw2z9hJD6NDbwSJdj2u0T9gBFjcQjvHHbKYLSBc6NizPw93V/mo3nfBcCAhEpyH3ihN/
C8fn+v3eieEvPK1gNnBJET6VbZcIWqlY8sDnWaBbYJKvcE/LD95D6tUU9cIors4036pE611MAIep
m9TQfOjt/jCREqGOEi9G5vaW7ur9hEZ/uiMNH2fUYWW+8/xEOZUp/pKxm+MjF8xIJD8sr5cwwpmp
befFHmf75iQjdXiymYd5jHtTGifU8hqOeEJkIFj/lr9qEo4ai2W69O+5ZnYQCAt4hF8TWYtP1PdL
Zs4z1wmDx/YdWvlSMSiSRgxqHMIRFfblBicWvagS3Y8UNnYV42BNFSNzMB7lUv2Qg883SdFjWESn
UJmJDsAfsvCoYNpqG0+YDr6Xa2ywgo3SZx9WdZ8bjsfZeukmuCQs111PRKVyiH75k7xmB5HxUavb
zid7pNO/Esk9GKr0AyZWCgSErtS9xNLilGp5SurGNRTkwLEV6hRRDvcuUEBBTcrIYGRFGzYpZgrQ
aP811LkaxV4KIDIL7G6VyKASTQGz1x6xQv/ASKgQnd1YhaVwRjWOem3cU1onwRCEJUqukFsFN5Eq
cVczMIws0R26wyhcRfBd69rY4hNxwH18gD2BRFHqAC4OOyb62ZnTaPWj5Iic7IhxnpDjaxqVQZIQ
EdLl431Sp3384wB78LOPk1Iscc1seWYcXmiLoFMJ8skmdbOcjWnwRd+dFLXrRhMflS67pIaSZmN3
WzDGU5LxGkD5jxqyVc08A581f6WNiUEQIqM9ZK0g3IRW4lv6iR7iz1M/fFqm5bPZIFEeSc5r3hTX
Sw/0hFtb9CqrGgo4si4CP91L5pKRgGIIzdeONACbjioigfXELoZ0U2lYVH1+RErKnGbz9EHHygRS
xbE/6yEqdaS3825zgvQpT4RfV4Xjp+syN1A5/PccV1EqNIl9skKv6LuGg+6bCTvvKMEtCthqNEJA
9TgmBLZ0xqh/DotlWyqV0c0sBA6KGWEm2oEY+OAPYV2j3TaPQJ/D81th9KJgBbwC16tJdnHkk7Ob
h3x/tiDPLVefyKF9Va8oNdAgItyW3AcSi2VqRmgpJEb0xv9feHRndmIZ1L1hCiQ2+C7O7T9ic+Ia
KY8ctLFUhZA9BX/Dyhidkw/qBjtkijnFitjl5pginHl4CmRtcNAEPF1OHTS1sYgsDCZWhPkiEt98
V52GJrrjTBW/2Qcm3Lwm4DScnR/2imCmCROoAfa0iYN5K+3sgO6yMSOoWu9GYT02r1lX6av2wEgZ
2VlibkRNZ8WwO9LTJqOgYqmTmSzfVT2y+GrZSISn2hxYCrsusOPBw2iFNCmVKiYkPg7MfdZYjlZa
k9rDqD2nlSi012Snw0RUW2PgpJqBVEYhwPGdC6oi40UN0i6ac50oCXd7YhL3ehtQMax/mL0Ibv1j
eH4vYIP/8CUKMxFVz43pfRMW6frvgvt/2ZGIuufjXonPUyOzSJfGeGIY62Frnq8D0VII6CheXRhw
Lnkel9/cvv0UtswccmznCRX0YBYbUycjNtxZdnXTI0vE7350jG9N8WcXDuvnVcwPqJrxaW/9TVet
Pnb+yRvR/lBCYBY4vGLQhF49Z5pKmv0k+v9iipGVzxvNEoe6GP6kVOxzxxcm28dDp9zywxD8jgNL
2VnmE095q1f20kA527YyCjqng+etdprnWMGsFUDAjMWFyUMiLx0rAHcddZi15m4GIAfSfNuhCBLK
9fj/Hube+K+fsHO51xVH3QH8w4rySHjjWwrWNTHG4jeIa/L5S9tJ3hj8RQ4l3XIqHNC9mlvbdIS8
+cRQyJTe30BWwc7/MkSQ1IYF0x+aS0d0lFCch6gUzvEkSQSteLHsUNdayocinU0Jyfop8SNK9pPB
XCOame2Twtetch9LqmYoZxCCRxyRsIcfoIUDp5lfIzwxSl7MCDlXtQaEzjD7wtA/EuY7kBZQIisX
AEiUGvTqrt8gFty0F4oGW14FrsE5ndGYNdhjoRADMkC0OVYbDGZS7X3CFzBDIMO+AKv0ShTQ8965
tEXeS2BS9eZo6i3xv+WgVj+6grCSDhKudVYC9hjhbPojVbg8ZwnW5uMHWjqzeC/xLDm1HogIyoIF
le0ylrtgFFBGpwYXvKi5VMZx/0CGnfz1Aqg63bAAiK1j6gNsYdjGcF4HiiCa9qcHgXjA7XN4DxbK
OEaaAvgTqARCNmX3nRNpkYDtfuTk+Df9lWC2yLpiTWl1smWyU9Lsy2+ETIfE6Lgwux0W6bGAXoYR
HyQLqNpsEC3juqkLWfMtbE+8Y5WH+FqKYTWOpy2o9RCWSxb5ksuXHL8ThU/dEJdbkIYO2appcY1h
cabbT2A5eG+Zb/V6QrbeaXWqEOsVXCjpXBeU9Mz3TBPyE5lMRbAkbacNazFZTzxo8EyinN/qGKAm
33iGXaSt/7abEgLw7V+k33073wXF+IG/sZRhNrfpYK2lqyN4t912Sz1CmgAxTPEqypecOHwKPTU/
QP6nlB5fpjmFr+k2HPR6Iegr31OtoBdx2+roTjZVIAdiyL2zvWY9JqIDJr+DtGiF5gIy9Z+/0txn
XWn3pMQRaeU840AFOMTctzRkqCg1bGTj2EmAuLkfLz64qrUEFPMTovobE1jnMLfNErJozjResy1o
ba8Mu+JPXtHvHWeC8+5r0U+jO8saM/X3gYIC7RNhcCL2cJBl/bDQGoiKiRoMsdBeyZrssnp+kOkS
KZV/QH1S2meFovBeirT9hqicMZ+hEauwgMy4AMbtKNc4ckIEe9ypvtAjt4RjfcSMsQkXih2xtR5H
I6+VnZ71/FoKtYHx0+t147it1xQOed2zKDhe22bgUNDkjPikTDy5kszlCHYIdHVWX+AJ6rRDtm0r
NhtPHxC85tq+wBhLNILFD5Knx66kUYUlGXKdF89LkSA/WxO9hv6ScowkMwIfyMV3+x8tR6F9GglT
FfT4cu9F9A6Q57GrH88IFg8pxZzy3w22TBNwJheJ+u1vd2IypuTsrqoxJr4RUu5tsWy6yKiEaHkx
1BfkH//OgDpEBakH796vZSFtq0nbtgj2yRr6w9v231CkirtaRX2t+ojtbJ2TYevkrxGrQKr9N5VV
cr0Pl6PG8LduudyA2LFddp7+TqO4qtkiNipe1KsurSNGAGwkPLwAaU4ifFQIHi8OZv3iGaqbXxBk
+gANqiBRzQacqF72v+hgHiekitwZm6wB6ngQuQxJ9URy0QW1Wh0I7vwCIbDumNQUJpW+qsZpcShY
8JBn/Ij/T86cRYC+o8vzrM0B8VVHX496SSgJXHWeM05FDCAi8xOkp79YLfFyVMrl5bKTHGWwPmYp
lQLn3CKC9IfQHIQYFwaMLCF2R86n+4lbi0r1EUJvPtRj5YPdKSdODGUKhOOmkAyB5mJnig6NheDi
hOueHqqafCLliFMxE3GG8qdctt5/WorTUgpw/DAEvTJnyZFHc9d0MdkQcBrX2EXSoPAtPtc0Q3Ml
Vuq4H/XlJ4uPHfcT0JDdA5t6GODevzYeuCQ+fbw45WRe2H5Znux6xYxpURyePv7JX1jo+MyUX7PJ
KbdZYjNc7vfJrbg5L4hwmUGlQX3uyjZiApfK0uNXpyphVL4ns6cnVEfKt5JATkW4+IvtGyE2u7f2
S4y/8CalJtczhDakgSgDBasJ6DgixmeiEwG6eJJNuVQRFSEw7XJB1BmWD+t8WHhCnKSdVYtHC4jy
JWa3DtzWbnOkbOkIlWQFUEqkjLZmqYICI2sRsTVVl1CE2MjNIkC8X53BiE/xJdIoBxsKqKmRqsDX
zHWuLRxQe6vTnkjzfovh096c4qHNlyKf96ML/tFmALL9jfbnhv0vYMcfBc41IrGVtrfF/DU5orUu
X8+zUAjIKR2f2+3nd7NTuQvlA7RGSsAVpafNAPjlkvwYzuV5J8eRctyQKWIK48Rib9RydHwrIkLh
GnkSV7KUrTATiaVTc4ltqkvgpNBeff7sy3uGEQtQPKidxO1V2MKtIDX0tx/Z2dw3THqFURT9iToZ
JEfnUnR6EbRAQWHASnA0by29JDS4wqq9QZE5kQUyHqy5gE9z7x1VVZQZb0qIP8ByWmx0GXt8CFBZ
vrKlbmr18J71kzs+72eFn11qpcEtWH8Q0186VnBTtXJb0k+qEZzRWyn3JvTpsKFpNEArYGmkrR4I
Kb3+T98vRzmSpn8oJ8wPLsx7lyyR73W0JRHoXFRDhsD1gnVrGKhbwSEOHURgjFAfUCzXSe3Lz1n4
hAySqtC6XFXhQ3Rnp0C/Z0CqtlJV8P8MS/bBLSgQpFXftMByEH2fzkG9VJCa9pz/lXRmh33Xpj7f
dFe0TTR59dQH2uxKAIISoJxgd6tsS7VPxPrb4CNrWtM242tSfyvyrlvngqW9kDGGCe9eRBcE/1K/
+z53hmFimAGUfIu9naS4pT/LIr44rmbSSm59YIRW1P3zPh7YNJvXPhmHiK8ESOqgC7T2wNm8ZIT8
s2sM3RjaUZ1sMGflGiV1uv+pTjWp9bflhtKuEZBBCjUz7P7JMJRElG835y1uTilvsC61ZbS7MG4M
oREzs9UzVWHyJDQLRgbfCRAO3Rsz1Z+M6mOh79fe8JmIlOIXWhBOYvbypWy5b4MfFl0j8+A4lz+X
RbKsNViee2zKDuwgRMeyL8SU3Hc22dRQ2/2mFRfCBEibQjjNMvegTqqXbRzjTJxry8jZ+48DpQOA
YUBHJ1/5Z+ysZfSNA6hgv8rwfu6ko3/zqDsPRQFxXkrnOt4OTjv0KzFqzi2NWc6S2HzisF/RJPfl
EOEwG67l4PIne9bG2o7gyAIK+LyyveiFXxqlepXESSgyegajG/bPY4qy6Lb9QMTCp0D0hbZEwhM0
/CKGbniLiuEc8YdKQHfNtUi/Tr1FHMA01kG8SQwbr//M1Fht10ru0tz0piSghYkPYov6mpXVGXVo
P4uXy03Ss1Kczn8AUk0IYokuwcGgjjHeCUPTqaheQWfEwuPFSI/4s7LWEPgW0CojUwLfx3SvRMf+
+BGkxal3PqWWc63A19tod31YmVX99WdhggJE18UkYzh+uO6hBQduakeXYDq28R8kIAZxsO7NR4RA
EvlHTFoA+HEmXVvqAYcBt0P+Gha5gN3GtEpWnCH0J7aqVM/O4c2qEpcAGT9OENYSEpFBBiGRcpmf
viaysE8PR581PQARnyVcVwVqHtbinDSD8IIQEBakzu2uewE0WMSgwTo+QDFJPYr4AEI35U+ZohYH
XxHNpMHmd9tPXn2rPkl1B5cmRfJLBH8XefL9QGAQ0MJKjIYqa5cChDK9mOFFUnvcE2TasQtsajDj
Wj/7I8RwmuQ13vOGngh0rxOUekAw06kiS8kZm4CTCfpIiSPD4E4KRK4mvFEmStshDg6qjCQ0YITv
Ue1kE+PYB+qI4c+fiwMdVjjvAWAIfqa+AJeOHBAj9y5pRgX64BZgANqEwzrRz9riwplrIeKhI3wa
OE03i8mAucku84IMbg2bUKArjhJaktBV4vhVY+HOvt7vaxMi6GDcz9btqAOFUS1RJAjeuZQwNz/m
MOzoiVDeyMsovTBOg+s736phLE05Y25exnqoDt9/ic2oxRxKKCq/7cUH5xuUczBVHY1Xq/DQxRtU
9ij0Cf6yTYaviVr/eEFgE3lwVA==
`protect end_protected

