

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
iaGK4Vux1Zzm9gBS3KKNmBXNdPq+lSqE3Nnx40zW9JpQDS5U0+JlSB5O0czPvIZs1e6N9M3JonU6
/VRFISTQHQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
hnTIGD4PF052NtQspkoD0qYNWsnDfk/EZli95x6g3PoDiWDo2i9hfthnklZPOTwcwwB/on/PGVLy
LOGgor+yT4ZX8UGtoSmScYDFDjshoGWHhtXrHczoGSF01e42zFHCzF3p+Kqif4EYEFLVI0b3qWfo
JoBwVA5mSGa7z6eKZ08=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
jM4x3jcOa6ByCa1VWDPoU4L7JC2eupLAavYhTE4GTMYrnvE7xP73g8zjlwq1G8Zy1ODZ+0DDopVA
JY2gdvefh3SJisXvlbuH55643svFB8C9ZXe+EMovXErk8XGGsVfWZZ9248m2dlrUXREntbWGdORb
Fvho+MXYXuv0DV2DKImT+u2TQDacpvX5e8ltSYsMmjYxEdkZrVMF9C544bgDvuCE9PfD8XjA3SZW
m5oOMSMtDQabvtrFCxaEG4NyuxA648giN43WXdidnKPUkuB/HxDMEcw9NxHOVNuLeVs7mrwTNW8a
Y8nkGhyssdB7pA+UlWrXAfs2U9Wpi6SjK7D2dg==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
l1zDcM4+iGcttYyoR8HHgtSyP4Fiyy45WEsaODDzemrDXcJaURYpyLa2UgO2HmqSNgBK4XdlSO3S
QC2s2wdlVLq0nr6twxtavd0Mc90p3l2akMlkawzSfWC3lR7JsZexWZNEb6frZfXhesr8/8i8wphW
9oH5nUnhDJDdlXi2xk0=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
pHbCg0c3yWoABGhh+X5xmKdWu54K0QNaj8yiI7dbYcl0s74Nnt3O7DJj12bDcjZRfdRoiT43bXo4
30QPK3Jr7E41USUv0QfI981OyCHaIYD9DzkFx/42CQBEOSHNBrRTW/rge+4hugPE8z0ogrEZGdei
kB3oPw27BqROJcBQEhzDTOz6PP5L7SaiUGBsXkKo2TeQ1sLfd6VNm52eUhSewTFcPcdSylZU9gjA
/KlsPUnl2PskRWTiOzVvvy7q14ROz/8yTOqbBslSCNrDfBQA/bwCsE4HN784FAGU2BIu6GH0W9gV
ySlMw5kMiPDazI4NmLxMcJvTd4Vi8xnRt0T8Dg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5728)
`protect data_block
Tz4t5q26w30iwd3d3Nhca9S4EXkWKA+yBKXZbNrNHjh66sgSnMrS+dU8RU3COw4zji8fe9VoNJ+e
CbVE/9T2GfwU6ZCzcOFlosufiJ+VbFW9NJAS6E46/gRSdRl9C7Bw+AqBE6Em74tAE44ZinpWkYbO
FEcUObWyfSSFJjWwP/ADCgkwFmFnI5lfLyQGz3Kw5TChaE3sXJZAe3PgiTFEv9AqWRGnUBTw1RrP
4hC+XxQBR1Oy/Gi0RQC4i6CwbylxhZs8KrMACqA/O0/h7wRKsgJmuCa/miPrY0wwIZD/vAJRa/X3
PhkMzZNPvolEOW+HosedVJ2/KM9tVRvRM5IcWWSmPKygTyvJFpEomGfPmAvms7NcEGxU0aQuPnPO
sfEqvs5D14joLuafHhZ6Y4ClxyA066Bqj0I4y45RafXMDnHlcUpXBh9vyIsxc4FRQFBWQ0jL3AQg
ilgbHgOaqeOLlrtjayl6Vd4cVv/mPxnl8pY6iIxqZgtPMxtlp4zCadYz5NtJP0zT5vNuco/TEeWJ
SH0d2iATjCTv6OOccqKSLMlNYw22LNdNAYOfrH+3B/TyePLSg/9QW85NrLYyRtlUl+g1hFXieqh2
ACCD70mzCLXX+5uXCbz8tRlpuLtBKPNQqssFc5Bh3He1L+uWFpztfZqPwRuBnl62qV3tqgCDeFc5
Jkm/anYZXZU5Eo1N2noIYVHIup3T3iyRjIJZzNZ95Pr/dG+PQcW9DH5fvNYbPX0ll6uc25LATSJI
rVA/UgPRswb27I7xEXBU7Ha4fef3s0x2KtAXkyJrFDy4cuB1N9FXgQ2dC6AIXi/rYeLtGhifX5zR
Ijwco+vnERzSO0//au0rTIUrXg57KKYOAL6K4pijV4tyIEoVf5S1w0Uljww9rgNM0P/DC9MrSPHo
fUQKjBEF5YP4QIqhZefDDMstey3JI3+/EsLzO7F8d52GC/FmA3UU7dvTVXEK9CzcmEd1FMrfldv7
t8LOIOVqVHmF0sDl95RCYh9YjaXMpuSpqebCg3nBl9ZdlcZhwBVcfcDyThDFU7ecYslM1Z4mH5hi
PK8OHoksN4xWiSZ7sVxNP2fFGosx9C2P/AfJuu6DXmHYyqCsSUCkWHDZdamZG7vtoy8iN0UyUMHU
L5zDFrcN0uibXZD7PKcysZoVBu2hTq91TvapIwZTHELCUDZY+ZoEOPnV+567jE9vuL4xjSmWNPum
VHNje7dI6wwQF2jrxgwWPrVVyu88qtuO7geat2B/fhcKafosGj055PiDXPQRbrn+hcMrxuSXYL4E
0GVqrpslDrO7/Jz9ZwjlE3DCvKLxcHyH4JTZC1E/Q5j5XUc3P7gu4GVowe2tOHuHFTRmQ8si3FQY
T0Np6O5sXghzT8j9jKVLeVJysxrL6ymO6IkUeA8+aiTmOng5HefPOL444BNrC6L0d4n1NHGQzGpc
LzvA24fLM6aZnA6qT2dZIL8yvrGwKjIDObpcm+EYU1H1jX9HHQ+iKyBK0exiBgU8tzm4en+gS87/
J+t9pts4BDYryJP//AfqFUe6nPOZZSrGC5U/w1qjhKsaEOqgDqnmTEft+4ZqwiDW46Myhg/TSa3I
OQ4IgrJY6AZp7sTadLh5yHY98WfLYvvkxz0HkZZi5re2S4R+l3qis8TeA/fYGDg7M/WDVckcJQCq
MWWvpnylS/5XWmN3AoDBH5JV7RYVl3aoT77Rn3ZK/Pcn2mI1Z4u7Okz/wFSFaCiDLvgiSPu8rmVQ
Tilri81uD3FOGkJsMfFfLR+PqYq6jh04mjCLQk/6kaugBx+dkOvgn0XYRFGac8esYYEoLYXbSCWd
T2Pv3KbbSja74BpvTsE8avFqfluK6lvRJNaSrdNbH+4pTfwXJXogoUpwyU8mmxG8VoQBZ6Yh8fCh
FlkM20ZE8QNIxwQvrdAiL/DUQcUq2qEktEOJ0Gq2i7Ss/F5ReM3xmTCsfE7ttXGJ5Tpfr32LEzYr
yzlYv/fjJGCcMksRfWP5nGtbmKapUz9FIADzUfosWREcOFr2pzW0FQdQflJ2JF8E+HUPFP3MPrSu
JnsqWy3xQJjlYM55dkQMRZwHQIfHGF4tGs7oYtqur2s22/aIGzWGBfh3aPWtmcMiKTU+z+suA3GH
Up9jYMOfffO4zHsxd/pU4fSbJgJ0XUlTbxhDZm8RVXWfLc5AgV9bZFO+7WuRsg3OLBNKAcdf3LxX
jHMAaxpUU1gSUAypMmrOZfcrkUeQIAxtpZtXiGILxHWOag/lev1L5bn4lPcAl1Aps7DEOkFlSTC3
UVhWOji2HaNvKdtHSoqNBlPRH7kN5JYGbB2i6xoLtLA5Tj/43D8ay4wiMj1QBwj4nDz8rYyTwbpw
rTp/e72Gr4/yZQUjQGnTa2MVTXaAfeeiZI2VthVBytCq4Dn9Q12vNnKf8hmp0cXqH4VlIUZu3Yhx
3aLxn9kytz4wV2SPp+fM56hMTQ/+pkgb1xdzT2s9wA86zSu+JvOvZMKL5BuMKY5JXd3kSGnRZIsP
3vHnVIYbWZyILjRXdvUZ9SZl39092Be9brWT3baQVLIj6SCeQP6Bcno9qrGZlSIz7jlQJ7Eib9JQ
h6h3vdFFJXOmiCBaXhjs7sEUxR8HD+J0Gf9bbM17uklSlRhHGP9LgvaVaXEK0x/4yxkCbAKS0nxe
xcegWn30F522oqWdqiqInqcHJrJn/SQCrJO7AUrIKcGI8neNumE0rTiTR5Lln5NKqOyxxFzcLKwU
ZnqIhVPX0pvEonbwipgSb53LK5LiWt/c/TgUH54UnOF3sOiVD9ngvDrX2BsfYnieFawO8F2ErI1l
RCMbo3jdZOJQJzgq4zk23WIN3qRMW6aS8q1yLDZbhTevEsclORDaKx+j4GTRyCbozoH4gaFCQoaZ
0P4/V04PH4cwxWFJcQ5u4MFLhAXxDOvYLHJbURjofEM/oKeYQksHNwWL5HFXVYzRk2I6oH+YQiaU
1GI6uMZ8G0NheJt9EHCpgfghz3Hk3B3cNi16+2/6cvQT96ZJH/XNsCZv32nQIlC4Am+P2k5Q82hF
qdXQgvnb4XoFOm6U3dIuKFZWjfR5gawb57MKBqSxcAFg4DHk9QN7VqJ3iKcz9vip1/j2cOLjFowq
gAr29n/TZfkLOb9vfdItSl7PouHRu1l6jWEzMq4TXyusOanQsfqThjIjvcwgzl/3oJNqTZhccALW
TE1Eg9/vdQcU/70BQd3ZviMiSptOrde/4wURQXzmStxjSYUiPUhiGaMytNo1/ZnXZ6+1pWwMiPNd
RRTnnUh+uf58K+WFj2Xsi0mVjdFHIYFWqfri5IzXNGA2/Xpjw4K0Vsryk7OK6x9Xcb6fmxAKQQ0F
bVTJngud67VdGA5EYwcj7zVZcEVpCOcdzNW1pPggCmhVGA4ncvpPStpwtdJ0Wn4u+Wq67OZCnnwD
kAgbvsY2KQINT1X2xIhVZXYNDEkbE/9HJNABwZdEjjrrnN6ycix7GOQVHnt6sNz2E9Dxuz0rrVSx
cvXDqWXHXOoC9IhyQIfN2K+UhgiOpcP4v200oEv27Bp1a4f4ESOsMSFdPEcTCep2Au/pFzHlhDYU
VxaFHB4C5dQlCtmsstChEUoJrpJdD1Zq5BvDLry6ULodXptOHcrhfbNE+d/k/5NWNxDssjT/+kFB
oG8IN1Gc+qI7IkbTodSGoAqV2Gq6U7fa8pYRM44DPZK7a17W5k9TQ/tvjgz9qf2I6xHSMg7aQAW5
tWpVAyS4ImKuWHpCGwvB3CmqU8zVHs5bCogi2cEo4VW8Dz7Ue4tSTjc6uSwnkvTsMB64vt7x+A6o
E1d8uIgSOfkJHtRIeTN6GTMj/K4B0hwAazHPDBjqEqbqlBLRvu4PtTWw2rYt/wYm6pFdiY87+TW3
/djzxbnIihPupD9ZR3bAkWReeRgWEyr2BHBNYagYnT5v6OauYgxL8pwF7rLhQhznrmEuhFEmC6Nr
F9rQq9yEvoFyhpcZj/ZnyUoQaPLJFjx3XR22If/V4lE3uXP7OuMdyyWCf8nBSgIYbO0ytMIhnypq
iUPfFPBTBJnYZLw0i9BiOWNN+azhVIhziy/hK1plvfyvCbCGWCyKHm3nLz9qbDQj5xVtHydvjSos
v+Xp1APLNQO3gm/2iaxya2T25QsldlPBYcjfwBu3oUzZS2EuUPdCDDu3zDHOtqpC3H1zn2kYTZOB
ecAmfYhKx0hRU0WdxsLUYOscvDjAq0BvaQCcKGRp62u5oqrheVG+tpOsBMbdVfMdsONx1IBXeV5E
fjX7FroT/RmzgzvHCN2OYk3DAxJU9/524XmWn72XCQNy3QV1n8J8fEiZt+UFoeRRTowJgkVf73KO
HtV3kQBQOMOd5UwjUGfIXDIN7hNh8kalL7R08NMa1XRJzamRBSs9Jea7eZHZ+6ObnLo6nbcEWGWI
hbexHxKGaR7ocZm0oUuOjpfsQqmfmuxHQWCiIu1N4OPEjdxebSOCkILaUJ0zWc7N/UAp9K1XLl+G
TnNrmm/PHQeAV9SyD5ySuDH4ufGKoHGxpacg5WmjRAcala74vyJKuzrJuBVcvwtB4GQvdMhuBROu
zElgXh9WSjyxj2qEpklsr+vjyJ1nDcidOCAyJPuFh2cnDadxT9X/3rKS+RLgSYIOT2T+kS3gDCTG
VUfnfhW4guNrvYRhkv98cWlmU1RlOazyF06ZA6FG1CTdb/jzRYDsJtzgGo3kEoT2GoG5dWqTvhCW
VvyYZXuvpZDejelgM7KYgrVt5BcuDI1jE3wHEscwd7sQVnswBqt3RBwbaeyETnW2mo/IruWj0D7f
Fqavim+kDDy1QHy5jmzB8QxNoay1aL2Bz+7rt3PP/F9C6q3fAD63iIqpmE/VHp9OCLLSYyZVAoLT
hSjubZB9m2pudw5kIRN3iwnUqr+cwcRJfUHkCTGkrAiAApF60wbZYUOR0dy+fukH5X+ZasXfW10H
Ym9lGBQvYdqicIiwB/J/4aM67Y8AN4vuGO5JfbfMRrsSeoFftS46a5G9smfgdr4Dnrk+ffIt/FTD
uuwN3HM4vS7Ewk1jW9M6/ybDiCt0AASaQwy8sVEBS9H+ColGGxG6NZkbVQ8Q+OCNLjdIZDtQuNxM
79aftkIv9WZ23ok5f3Y9RF3uqeDUvMWcb5BGJzC8SLuf0keJV4fx3oaVJmeC7MFVbftMMyr2hs/3
yiiLbYq+l9GVtkEVz3vnoZAYaI73h7taLwoeuV0mLOV9Wn+1xfa15Lmtg9JtAMeXtCiLA3R0Xhvh
zlx+bBZnIlQrzTy/o+zax4qYthds/IuLrDN8uggQo5JzXL6O2taZJrrFJA4MaZ2MrADMEwjfmxeA
0F21lT6hKaGvem4KK/1ErKZmTxPqQoa4sMH6AegLQhCmKlZsGC75z9zDOdV6a6ifgVaWNr1ilyhJ
JiLEjs/dBe4+bNC2LlPY6o4T9HdCxq5KUR1xrlu8USoXQSWt+VJB1so7uxdXRlahABqwLRCYanMk
QV02tjAEGzSkiQmWvEFqh4/bdPss5tksgECqhxOvOp8n1LbrGM9RGtLt7oKUxWWa/P0BIlY7fWo2
i84eC/txkpnx+RUYJo6w9m0JWO5DH9i6Yi018COML8gdI4r7sursNLGNvnbeM/HwQ2MY/2/ECdFu
3/xS1/S1808bTnrBOPa6CVTjJCHHPSgZ/AZlKEl6gQzGICXNKdjTmantXPp0b6o9/p874S61cQ4C
V+u4ljSmHjMFOEVW/H3COCPKf9tq6K3w1YiYvSMhDTF4s8jRhV+DJAWbXaJP03JR+FefJj1h2TEg
kkxzAevbAE5POTisMaR77egFacZN1JulzKh6+Yg68GBdopzUNGOyy8cU3AeXGq+HaUv8NCrLvRii
IgikATWjEqV1uCKi68JEwkX+E++cdneRHDpbO1ydoJNnA/T0hnqwDWEtF1gRTtxF0I9tQxQ9iUD0
lhMh6TnYbrZl28qvFFew8cSz+Yvh6rxky++LXe64JoZOI9DV+hsN8eEBuDyE7oqpR8ulh2hnLCdl
gIoR+d9QalgQoWdYpGLGwG/cg90htPHDCJ3ZvdxwZoH0QorlZmGX56NXHxbWvjD+s6DQtFqASK3r
onTmeqEoAkiGfFEavJaJU/Q2lcAERMBNVOGu+OxkHpMiFO5SopHtZeDpr605tmuFNlLfLY0wKaGb
nwDvh4kl60ZietL//glzdxEemN3opbefTT8I/G3yeWYk6CKpx8WKYApIiKvg/5Hk3CeyM9nFCw4I
bJ/dJyx1/7rGieaZhBuZb8VzD1MJTwvm/3J0JXXiGXZIH2/TytZtn+ZxTiEAzaAqEAApaocaQqqb
ffKgyna9taHb5aKTDpdhnherCDda+lHsksUT7yAFgvrtPbSbWbUwtskhaOoAMFmE8woBnh6BaVZT
5xWdiCM5Tm/H6upAZJX+/gR7VUDhvNsUIW3yat/t016a+BwHC+hMeTpmAfcl46g/S6Goaz8yKt7w
B3DnAJcblifufF8F62Xb/x2yyoz8pkKg/8U3lipP2WcnV9oFtWoWmYqWwG1/uVQO9xItkGePY8sB
ApLeL2HoMkVMK1SXDrYejXQY/w6d3Mcs0SqRsSVXIXYXpVNvpvT0hdgS0jV0+SNx/oC9VZDHHyWz
AxCUNYgHM7mpvqE2njGp0UZRlP2FfDgOI35+QsXNObAQmmxUWfol9kWSfUPLZldTDkhIv4iTx0Er
GIfnWQJh0d2XQzoMr4P7edjXRqOSAMsf85oGBr1I4cdPnU/yF8UdbSeiO9F9sLj9KYVVrX+BsAaE
1gPS5zcf1HL+ff2AEGnQaK+j8Zia9KJLr7tccUoLjtU3mRSiPqR4FCEiVKZji8IjeY1YYeKuwRml
l0blbLLjhoP1FP4nPlNXXtqG7F1/J2rJ3qfYI6efmp7U5BZSvxCZX4SqpkBW+alAZ1wda9YYhLGB
tBeegGxeDVdxW3jx2OrqzVakJkQzcbmXE8clBVwXH4IDWB93VDqDDy5Ae+y2zfWG09USHtAKZ0WT
km1pIehMiSx5YYZEgWCDzlA8FsisinHh7MDvNmSRecNUOwAIPt2LiOaqijWnaDRebWlL0qH02RM7
5B8WkFksPpt9wLTSvgRXLOepkgEpi2bS2qRATrvwJ+8YfDY+IZF4Z5e5zizeXcp5VVQWsnDZM9fi
DkUrfmXK6Lr0nOBqVjLB0Wya9Q5JD8LxKJmkmRyU3HZvPhQIeglHqRSftderOYzZu7/kJNHrXjV6
0lqFZG4GPvWyCSJfbqtkX33v1PSb3fL+5ANNWcnp5URY/8riYJeYRuIFbVoX037QXGOKR44Mnnx1
4RKYXWREE0fJWW2oQvf5ACtiH0j0gRr4JdaPSNpx7e6eo8gqG+7YEY+nU6M5tpkxWN88KV/OMbkw
3bpk3QT4rMjElFKSlJq0u19vdYIqBzdk+aWIWciWsgM7Oh1Kb4IqNryRmrhUmFiMg2Ml3VwA1OVl
SPXLUk9m9XCscshl0l2cCOaNZgVe11uqxJol6HcYqviPEKeQvQ8mRpIGqDDlwlkMiBVK25iLQKiM
PZ5de3F2V2RhHDoMJzIX1/Wlr1dx7fqcONeV1RmzBK3G4/t4nMclXbykj/RO+bz5vZcUqGdIdlu4
TWUS0TmzjXfB+QSWCWcpLEGtHv9JBASANDz2zA==
`protect end_protected

