

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
MPaacDM0TWg8wcifAVW4jEGylx4PKrqc4CLboKEk0r6t7KyfUnirQwQAphZDsR83L059CNEzB4wD
M8AKmBfOkw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
XUT3zAfEi3anHP5UZ9Q64SRw1RnMtcFX7nJsXqsc+jcNnlmbg5PdhmwV7UaFs/PrWKFdgim7UZCy
o9NtHbXd3iHyUEXXZiWfkC6NC5Dndoi/rfKSxw5AtxtcCSaJ3/cb/i40IG38fEOD0mldCmJ0WOZD
xOW9J2aHwV12uWmmUBs=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
5hB2z6qFvCHrfde+xOJHAAm9Y4Zd5X0rYu4ngUzTSYyHrr6WAc0PuLxe2Zog3gNAv7DFoV1y/Y4U
F6T4flnTjzAqIUvyAW8+maZzCAeWDi8VgmeKHRbLydt/JWB9Ri7GcOoofnS5/hxq8wRCMMkoHbQF
kNzxfXz2j2QXU8RR6+E7pvqcJkK5H/P2HIhS88SnGwppr+eD2lVT18h0s/QB43BH12kpY1JIkQU4
LOR3Ej9QoPTxmx24xAodMjc6qGME333306vLcWETw7evLQ7fHCoyGS8qVr9xvwEOuA+HtAnx7p26
Z/azE34tKzoImCmpb36r638Bv/NLBk+b7agF9w==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
n2iw7CqdgxuZ5kdEH+pm9NjU5keAcvOSKkOt8pim3KzIVtdYby3hWhnEsC/F1aUQ3kkgfoeHTv/o
nwfMP+AVXxDoH7hATDu0iX0A8s8avaGhFp6novk5xXzwMVnGP5Rbk3GwwADpRNWqzKN80je+JhyS
o3J4z9hQTmce/KBAfWo=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
sR/mTVuOveJs41YLuqwkxNe6mc/KV56Pt/6c0cIYmcRhmwLHOU3+/VfoPpEClea5ISswKcgmSmEA
91cZp5XMe9E1MxpJldN5YBxK+3XVJrpKIG8b4LM2yC+ZTp/81AZ6CpAKQXOcZAota3bpWOVB7WQt
kPn3pALJ48nc4gaIOk2j5GO0g6BLITkCLwe8Z4XOzYZAEaEB+5dJ58Q/7AbNKHr5UdGO2UVVG5Oo
7GIt9ETizL/sKscnCI3CshbxwDQPtnh9/CAQY2Ci2Oqc2ptOmylUrV0jpazJ/ulKvyLMe7D7sjb1
BOUUkYAI7NZU4AkYW+pW9jcllm96HEkuSjkTDQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 50560)
`protect data_block
fVq13XkSVaN/HRQ+5ExgRF9p0oZe6gIHSW3gCdDM2FDpVDEuIpLbcud6OxIe+oAo6QuBXt3VzlCk
h6S09wn+2+ZnfQqSdUSnCPiyJ5tgcKNBEudx5Zk2EeTU9dMpwVCnOLHFRXa8siBmwkLHYIcx2LGw
Bgoji52Bi1oC3X/2uwJF8PpAF5X+ZfkLMr84sL3gRCAzSFrpMOsOAJGucO1A+33W3qYy50xT+a0n
a+uX85HtkJdS6/4SbcSmmj/z120vP71bOKtiVgxR5/UQJXCd3jjEYf2ZCswDr6YKibjfGB2RJjAf
GxcdRSSSGpoUByqRHOFU0FPBb4ii6LRJvm3g3WZ4sF77F6xDNzVl5kZFRoB5/Lm5vIV9f1uMrOoU
Un2tXU5nRNuBj6QeQMS9FNiuyb7D2HRkTgV8tPnhcpTj8W3bYYsdycBGCS7+U14/NYMXGKMukzDt
aiSH0GMYZPuiJVFesLONmVtFdqMv4a+/l7Rc9j2u7vT0goOIonJXoU1UrmPgMfG/7RLdx2qJBPq3
3inwXZLGqfn3FhzchW82Pj56OlQwLL7vRsfS4P6A0xtJ4cjQkj7duKfL6TcLRW7kKc+LF1gxt7S0
gWR/Nnj2myxPhyfYgxJq3B/StBJdLUJlNf9woqaGGF/s4dqsyJzjdC+y+w2MaIl3td5vpca2lggm
MglsDjWFBiJYGI4ag7eaKAxlCIU+iYdD3j7gOfCW/ZYHbcHsGDF0OMZjdZQ/LPPvfsB5bpkXTaGr
Ioc2ZQO/mHACgY8if5WXfNNmC1M37ftODdfWjj4L5xBdIJJsKzz3JDwiKB0lEp0eslCkxoG5CxB3
BQnNbubYFX1YAYCqMdAB9QtHeFQtY19cCIsLL89RExLlKmuVVZ13/z21i3pzXwSH62cA2Fec3ysX
Etq+8+fs18hmkvSypAgTzv9Ie91GLW5v3eOGJUmta9DV+57u7iuU/H2yV1YbukJ3Bbrw4GBR0PTv
0HZd9KgHEVz8RetOJ8+WfL5ioM4AdSYjYeVk9iHtzAK+aQ42YFsh6zEx90ropDo9z9g+5paW/gc+
OxaqnEGP7iwmGycL8YW/l38Ak5h+tjQQetLoq1QBVJUdpDzvCC7QSBpm0FKabn70Aw97ont1nKR0
xlPc5WSmi5GlEcEM/cG+Ey+ywPQEO8hlGmiuZ8ru8Fgp7JwKNKj9YxN89pWDo6B8CNkv27PmFqCT
IcAk8JeengdVfmRSu6bq4/SZq0n7NJpqnvUz8uixZWxlhqQaz9UbQk5jTVAvH1d7VSjmiCl/ORKj
tZLZiIpOyLPyY6XcgKoEEULZmJLSClzoV0SxzS/6jmUEQMiogBqDLdf00sdNh06m1nRs1RAJ4hhb
2ar2rXtmSWDYhY9AHSpedT5KsR0EVQwx+E6F6Ph8tPFCPwyrMH+NWbHDcg6KLmqoYi6UJtKwVewT
vKPzLb6byLPxw85YlXkdXx1mYJeBfgHeWCD70T8NfoMMo4S5QhVoTq7LWWlSyY0DgnkbuZQ3AIGQ
0l0bRKnxNa/BBGlmrsj1qcl2NiRB7YoY4VAeokFw6Jot0X38aEmCAgSnOK316BQDrio32PewJQ/Q
swAhFMAx3MapROl+F2IFv5No89bOgA1EsNHFTkkdtQXnFrjZwErRp8d6PTDjrNrFIv/gfwmoM8Qo
txDTcF0l+5fwvzx8RKLPPCNN4BHd0rq27JttzeZwGTtLPeTglomF4olEzIV9s+JXuWORa1MjDnag
Ez0Mx1iUo+hwsbuMmH0l+9T6gtSHzJDXa+++cj7XS7bj4QTARiZR08sWlhq2CvFdF1GFYnahP4qh
JE9vlXr3ZLT62p4regYEiPrT6cLfaB28YZstIJS1u0/9g4at9ut1n11x5NXJrnRCh64RLOo9ZJjn
N9jEohiB9fqPj/Aa4eY6Tr/xDoJGdqLHHgu/0JO1+hCUgCQaB2NaKITU/ptaConZUtG/Ntgi1lLk
TxkRkK/O2da0SgjO0BO7UxnQuBUXVXI6WTaUVAyAdwYaL/5NmFJoeKtH5j+ajguc9bG+M04bllcF
M6i1SNRzOhvhmmBZNLa9rQ24JnCVbwLr9vSCygGEBSCbHuKmk0fquX7Jc8ZGTCXErzn/KX/+b2Vn
6qLA2D0PVJhuQmc38Rcaue10LQIeokIkyO8M88l5Y4WuoQ/fz4mG2/MVGEHp0zoUcjDS3xhUT10o
z5hSol2hsgmNA+l1qWqyK21Mc+tuuQbGm7cI86XWG8Spk/6J8Z3hZBOpW/uNmZu6pe83H97w/+Km
PkQBktAV8CEC7A5YasRw6DmU4Ro4PA/UpC/xwsrTelWr2EhfM+j40/K3o1TtVDgOTT6xmiIw/KNb
YshxODM7B8fcmx6BeI0bI3Pznl/3CBfTCg4yNaW2o5LOvifMdZuZfPJmoK/BzuzHcV1kb7neSccu
5n2kn329TsH8Lw1AC6NBVgPH5G/cwLwQC7ExdvLcQoW9PJWEX/OA5K/wCSs5G/CKvphss2PkhTbE
jS0YV/s9e3w4GBJZXJn+eE5LeN59iY1LeSpQ9rfShtBZCYq+mILWB4qVDQ6vJ96thJhKrITckJho
U6W3nCrxmK5X0jXIpo3HiU8q5bt7GT62j3Xq+VBUpjghpNxxySE91lj5ZPDMryKcliT077iJy3jm
PPE9X9qENifjD/wBf89s1NJKGND76DDiuyo/i2xFx+mpdacQzK8OiegJHSmLBCSquVCMjC/f4t6S
eaW0QzES0lf6PzIpaMQ59pxzZzIFV7xyi3kOfvRyjFvB/Fqx71lFt53+ZcpnRAL5QENscc2gPF2q
PMg1mOXcXW5Zfu3QCxsN5DipPXqwGoQDfKLYv+dC8hgzEhf+yNpQt6PaoBgcJdRdcjSoh3KpI/Zj
paMHscPIs2mv6DCwfEveYESE4YzlvOF2vsNbwzEQSNSE46O+WI0YFIwZOsrqK2ylh8HvToseoNKm
LVw7SI7rGEAR5TFan38RoNvXOILi/ldv7rZ56egGIcYdv5NW+tV4PJ2xnvhZp2F1lqmdFREp/WWO
RyN82JLkLCIdO9gNf/gwxgd/1LkLNC47FSBBJ8MggQYBgh0UHKpBVDxucZTtp0xeahGnGUYj1SkT
29FhJl+Y53PupjHbfwTQaL0X8XO5GUJhIZP+hZfzo9vYEOCaIshxquLNNGEeLiSrv6UgKlZLLNho
QfZTOfSc+z6mO5cfzAH0ZC7mVH9PDsHnxexwSSVUCzT2C9WGh+fo40bdN7WgAwT4vZjwmWGBObij
grWQnPbTZzB1MO1UNkgAIZO5mcXlvR2t6NpY70rRT1R55p9lqsRuZ7bIW1e6wg4+S6D1BozgH6mp
ZyPKYwRZir7szucbO+hQyCVVDwKKmYRIY4ff7WIysdeO8+QRTWjoX4gYd8rKM0AhsghfygiudYNu
VHgb7+DIiAIh4vMpx37l8HKd3wpwimmxCLyF+wmxfPe5ZL/1Q41zOZ9Lw/vVMyH/DFQLl8AlQzFH
b5zn1W36r+RSE3K+GqC2Cd/Z4gQL8+HO448IUjVvlTECWJtALcSOM689FW3+ok2dyw0yPKet7g3C
2GM6EjYupC9fRjP1oh2fPrNdQkwxxg8uVVYk1kFyTipC4jb91uyWOH3JZ9g863YJV1925kfcfYfs
BVhJfZS+S6b3WeqAIzEtgMMjo87DXO36RqoIO4w/sG22J9hDo9lDCwGjCwUKZ+07S7uEWoQKKft8
Mcchs4fhW56bEsO1MQGOu3Zd1LG7OuLgJ/3HbBQ2vkppgJlYvcCMhgybUdcUmuVBg7CXKALzygCG
qRWqL09I8YeM0P+GJ5X9hV8XfOPk0PrK1yWn9AsRfB59WnRHzLuNsJvZIlWuaHBbhWXvX6qSlwgf
96f2zRiYpvT5vu8PEw0halTJI5agcJa039K55e+jqP3T7B7F9Vwh9jTZUZ3zPT6MrzQQBP9jWMR5
oR2Hh2rWJkJX0YgGDu5sEzHsTIwvYeBkEVHxSeSPqwhLho3Gg5h3cY6RCtQ1TzEZc7QH5SD3Uvah
uqkaAzhaovlPbVKmbv+/TcXNQuRDgGFlHR8Vw72bqVj/Be8yDUz4VOCY6FZbyaLCjakkWtjKaYmv
o2YQAqIfVh58l9inxEh7mWONsaPnuPMZ2o5i8mm4GdxbwR9fjTTqxtym98jR47PJXBVux+F744sH
k9N2mvO6/d82M+bvwCouLIVg2d+jrHkr6bn4i8gnTSAr1yr3XJWLuzUv2geIzlFHrWaTv0C26MH1
AwYEWYk+jikrS7XUGSymzPKdp39/Fs7+mOkCnGOFLepfykJSpfnt1A2i9KnOPwqyBP042o7kSt+m
MzXUrWQSqqWRONfHiBj7CEj3pBNGLqe24cGyqg4hw1UpHlwoeNqC0o1K2+Mtn1tGGqi0/wNuPEGH
fa4yVZniFkWGQdivw0QrZmIY0Bli0NUn8PV2LagU/wXYdnX8pPSXQctFRe5XljvZgoriiDjugcnO
oUIsG9tNEd6DKcpjuI0D1h3KWoFFM9hKV8yKoUj48g1M2PAwKQkQmsYcViDomWoy6tOhcq5PsHtX
pxna/mG+W8veerNaFcw6XVt/bJhc/kAozokC6qHTmFC/KU2xbctvo5sR8QORBuS9iGSH3xXPLMXI
BYKsH012HnmP5PLUSS2GKAPH/QD6Mr7xMlzTm7GXMEsHjwJAqqKD3vcE63y6coQhzs/U/vaDWMhp
p0PUronhFFQNkEGhDbScdp1Ajo9oDuaPrsode85FI7tWu/fQW1C1ucYWX8i98JC6i5vfgn9ZkAgN
8vY+JEi5x8qIwv9vhd2fR+Zyr1Z81GY/e2BM3e+WbuppZEW2Rg6poZhjXolTPoPFX5kAy59SEes8
oLPrWCKPtvU0g7fa7HdalJfcuRF4ScP6xY4a5n2yWW1lZwm8DnI9GVmw/8DyOfRWkNQqynSj5ODJ
L9mDLahF271eFS6k+TzAruDWt7uINIepwOqcRSKPmPyarfEWIS7qDqmgR9EZS+qSXQBWPRsMWMSj
fQ9ZXzq0UHHqDLFsUJx9oQwiW6gfntikJuCEVvgYXoKD+91SmCypB1TfLpBpytCI9Px7d6YQCXl1
tMB7ey/nvpJGHHABbDWPA1i/fEzfMq8GfQ/MCZyvKjxjXEtSNOcu9OuN/9RQlW6SzTWsnHkQ9FpD
27qg2pxCIPxkTsRAZz2zqWTpDKyPEQPAobGDKC/4G4xxcTVoQlMYNiO2D8zYqGK7qYuL+YypQTxj
9EBD6gP2dBwUjRHRTnrfGNc3FOobAVCcvkqq3xXX2Gk01cNL357flQoHGl8JrFqT3BtT/FsbN4q5
Zr2cb0hzx+906TRhVnq/9pBPSv2DdlWmc/z1ABigmSSwH7bWDCQssleketRbbzjROOxnwtCuZIOq
PNB+IUJk5oxypIL8nKfFyU96vJW1W92a4T6C34/d7jE+7Nt5DR9fmUPXXhNvzud8sdd+dqA8qN7j
i9FEHXIAzlom2ZYODesGje51CcWlW2beYPQ+1YX+e3zpvabi8dzvL/+fhLXlayXsadkYsc64YYYu
V8coVXiFZP4Bf93EChOQvJq9hZ0DeB8s5WdBYWpdirCiYoECXwfhkwr54wJt9LOnyaTQzr34HR01
BXwHT6LbHTUS+kf0xXemhcZVFMlkI1wBfJsKksrhsg7mNikevB9sjCu80x2pN1HXE4nis4nLWE3f
zOQy4KskzTwSmFWRYm5PDdnfPHrdmcnzemY6qseZy7rkJW0QbHelEC1LsGmDFmJUP57kF35rT8Cj
cepw32jHEQfU2jwiafp11BnKYHN0hmtwlRl39KFMB+tgYEzqYMwpj9bgyzorisl1wdZArcVVW1OH
9nj2JzXuSkbvPDadXGTEFxjsWjxm+kuieozM82u7+0rsl8eYmiUngR6vjZCnR0Hexh2cOHkepf5+
ek0MMsDq1ZRTjxGNRaNCf4txCeZAPDe/AqP6Dw12WAM+9nKZQyyJQ1gE7+YfjIRPeaV1elueGz5o
75txVtiqmGoX/2oHB2dO3oYciDCPq2Xzhyw970G8leU4UcodDKZUYJf1DXnUeREJyl910ka6SbaL
4trWOjCUiDFSVZ82duawFVVO+p7+0WbhxIuBwlTk4Qe5jQX+QTVFPqShSw++fx5SfNBtB9eH07PU
jDrC121jlhVtbk0OSAB/Iw2A1fza5vx311PAX5fBzpxr6e6c+mrpHIizBNHZk98LOcIUnEABF+vc
N5f/8A7uGxO9MbQIrfyonnh5VdInCv0IiWm0JLVQUGLA8gSzabcWW+0Ew9GjTm2sdsrgRPcK04uL
XjHoQQrxFi2XyEzWEI7VK+rFLFP5IBJPPtYsYcmMSswHTI6IRCyk6E/Oe8VMirVh58I/UCFEtC3n
2hIqDFZdDBx+wWV1Jr3dxdtDpyhAFtxQcz2wM0YOjvGonF6JNx+4g8KNSsQo7W9m6u2Teqb17dmv
5OPNoryzRyiw0xkw8lkupfCiYxk7bKOplK6YRc1ggK0bKya/O7mu22onpDau2vBmGK5U5LX+tFoD
3ZSU/5eVQRTfyvyrxIfEizhKZiouwNpV1AbhBfb6nKvXTeO6++XLt5du7cTtZN/7zvL2JmTTF5YR
LENeLIK2zWkKYY05fe8nNHyBqagKn6If/M/ZEt8vBZByFyH4d/Rc00c5MDesMYB7uh+3s5xHaHm6
skx7T4BLOoh60F17MXHZommKwAnA4sKT9AMDdnfRC4pX/2leNwaNPnGPPwQAJvI/e2Tq82Ov/Xkv
eM8Js9WTIOqO9F3BQV77dZszvAwgMJCLKCqrj8P42O5lohzYk9qhHsGTWdQhf1VmJCquVhELRXCO
8Ui00qqKnpQ5bOjmzm+CgNu7RBnzrZDUgf3sxs2fPzrNVPE+NLHSKH4F58Qk+RfNmoIw3kf+gAeI
vQv/UNNK5IBJycOEc8+jzCKXQhd97mxfmQR4SlVs4OXOvQY+lmPJXWI2wjZabuiup0JLtJJRNcRi
sq+bcQogJLaprizGn7iVR/tJk7NMe55a+iZSy7sKpJ6PzJJF+5LF8Ko+ELFg/bBZ/cJFs0MddTd2
mHowBQ5yDNsYQ9ld0NTwRNpwS/8L0Gj4cU0DFwt/SDEjWXCBL3cmI46uX9T7Nn+9f+gYL7yIYY1t
3jHnaBI8z+BxynqtWUUAhRA48ZBFCzIVWnjx9OVAAgeFXUlG5mzkrjJur94yY2Ib2xtCYVkeCcTE
My3DsBgQMwf4pI7eLoZVfqFXczJSIjsmkVrjP4RXBmMJvycspywC3g3wsD78zN1S8k0QGX1uWz3v
Q0zHuomuVOFpYIKx48ZHTfMCjx1fJRf1C4C9D81CWQZBi1IwvD13rt1MdMqpxljdnkPt9wZ2rJTv
jkaVAuRRt1jaoNoaykUKo/y2KCvusJJ4/F2EMzDNDDCbn13bWU47npWRN3yJZkHKkZ5uAptE935h
YToJnXUJLSzAJZlJOyAjkbOpeiRrZ/TgUGFgZ9Ubez8lnmSXdPJT7BE/JXcfeyNepgMtTicPwzjj
uSBjnJewc2ryPW1GtxvigY5/Xxe7Q+XUQdEFMrpIAuvplFbhgKRHwccsUJl+QJIqlHQYlR7Mk7/5
70F7oRKHUbgy5sojJH/rxfvEyqlJhlsnOGOLCEulh7tBiJSz7E+raDw4BZQM/d3MGns5374NZ3s4
303P1AYhB5iLhZMBDA6CKshvLd8f9rikpcueqwnupryPEs5bFb6PC66q3ZRaolk1/0pxsfhNVJel
85bCp2YUoEiMTaOhyz35SGJbpFx3LXg6dCwSl3c4yu8/rtq/31hYOuRfaCvI8RbQp31FoqcZvdaB
QWErHL7s6geeGK5QmXh1LWhfsf5chm7tWPZCQcwZE6ICot49XuK7l+HcXuzFcbBq7wtbdiZsxgNm
eMiCSy8LpN+kPGu1OEX3TiO3XazKGJvE2H3b3q23u46+AnaxRLI9TOflKdswFMZ6KmwZ6ds1ZzpF
t8Yizt2ppZlLBsfexixsLY4dJAl8Law2swPLWU9NoJzk0LMHYp/C145Fb8RfjAwta8nCWut635h1
8XsBhE6QCGcg/FPF7GyxpvhcgupaYiGexmqoSX8qPu1OIGeRD45tW3Lk65zwz2qh4oJ2pAd4A4dE
zgCd7reeCovfMmdcVVlzM9ZuO24bkHJU4374CVAwJDEBlYPFO9DTwjjepgGOvT/ttBTotf+MqG2T
GEp4xyYARMu5YU/GMvW2yWQiJvvsrpr1pUhnjnqqefOix+jLTR4PsOEaokIzFOxnipd6vmNXfyL/
vE4ivTc8GOR8qUg869EDLl/uxa7ZrlKH4QTmxHvFqIOx8/UF7HNnp+TqcfR+JWr4HW75N0I8nk4o
qP5IxmXFUvD/AzoFJxOV4/cPzlncYAvcgo4Jy01buMAvF3HDm7oTwLWlPaLoneVSrEpkSJgovgJL
7GWjVz7kwReGXBFqXPkeRIaz2gDmKCofeIqpHHbMK9lRc2yvslewtBKgwDtnYplRPZhfFxn8myh0
1bgzZYVVsMzZk6hEOv0mTMF1LocEWhYGlsYucUIV7+byYfSRaHY5bcleIurCslpBKrMriggnKLhk
Y8k1hUwImXieO0v7fnvW4rJD1PZfpNzjtrsA6xGl2L8aQdwaHuP7aS4z3YTx4bji0BftMO79Zfk0
WvbsSWNzbMczb4BIv7/Abv/coPBBe4IBoCaT8SGlqdFUN9dAri6II0/ExP5vLNbKd5wfglsjgenK
QrckuAPqL55B7t660lex5NUHG9nK/ILquPSy+aLrVFoA+f4+sU+s2dNeTVBnXhaWETR8xg4dNrBU
VaSkqB4Kgve5Wu1Zd7I8DFNpEbnB9WmKccmlwNeJfiaPYHUHzjLmssBJviaKOLY8ujEXJNHWmFM+
UjrhU64sFOfXREp5cSDV2UwPhEFwk4Kp6F71nWlZi/PT6GU/xTPeg7iG3IOaWxWBN2VKLjLbnhBW
07BlwY7xjtEhXba0b9AqAEgz9NUXhRsC1n+tVOhBgvMrkebqqCs53xW29Ic+Xgl2+58av6tmv9It
gtuWswjgT+yA6AkRG1E0aTyNO1Lf2TxPTn+UBvdocnfl42CzwfeA+fyh9wGh48ofjTdkmfUNIZlr
G3lFdY+o9KaKiVoW913BsBzgojY3OJFZOPlsjkrNgP/KsFbOfA7xQ716M3PQ++GVjCfGlEuMc2C6
1eQVV3Imx2fM3eJDNEFjC6uPTeZgqO8RzciBXCmuI2pAkLhXirviOqIlk8vTevq+TJgEy+UFmzpS
0VAOTdF+q4CFYoQ7vkRRPRR7HbvpGOMHLPXPuIK3bkjAQ+EFaFFGr3T+xgIPqYyPZGuv2jEaGS/c
f6KBTHjIFn9+Z0DAvNZRv1rj1v04UHcXc9e37DzfK6xgz/N6R2jRMjb2yYWmnnhvinCTYPHLmUJq
ShpVpnhbyLU0NBF8GfgnRzwsV770sw4829dqt5ngh8ng7zxSPLiAFBwFys6Zc6nfWS/JJwIAvxhl
XQ2e8e1NpzS/exqeXLMPjIRHy9VdOQ/APsW/15OZZEjSk1EH3B4VoJCxCWAcuJY3hSJwlvM+ql/t
P70TpHbeDVbCghEpn3Umh2JeRm2jpVEytnb32KfplpWAV27ph06zpC5iLKBPbuez9CneSk4cjaRS
sMy+qJvBI8Q1LPVmzY78AeszP9GIu0ASK96cOiruX+vpTOcKUzlzlJQPMjG3lDJBbfL8SAHqugp8
ylk4GCsv0X2KiKgCQFhwYrpGiD/HfVcMhcGY/eb+5QlrC5l10HWrAHIZbQT1sphSm74HCFLoyR3D
jG/rWM1Y0xoxCvk29mEvwNKb+J8EpWlP5HNT/jh5IIXHdvWBsJs1CFH8jwnf85pZNJjj6nbdJmdQ
FnCF2//qx8W0eyJ5qhMoylReWjXX12jGTTu/TsosdEEMSbzPLV7aCqakhQIqgg/I81gm98+PF9qL
5iD5FbA/5Tg299BmirVxtTvCKvDgi17OLpZU7NC8Gul7DzUwIf1kxquEI8YSd0IcKuZdp455xc3J
KYy2oB5PY4uDJlgJDdp1OerCnB9p4pUAovgGxT3qVEQoNuUm6vMHpZKEQSJDt17V2kZGwdUq95qh
ZMAzVsDBiYr4Wewr4+9S6ohOeiKGFGsnyvhOGf3GBwnVbvyai9SYYjwybcAOVGx7iGjOOa8XyeYd
xlARTCxHjypqF5iarYMr3z9TYxGZmVjwMf9/DfPdqYb55Os/TMaJJC6zNU5fjwAZK/hnAFO3i575
mKqhbSxF3G8cft8LpF/Pwdy6S65QyrZXn7aVHTv61WGEHTqi3KbJc6K7dQ5yc/Zipl+r3JWAYhEN
iNvh+VpkN9zPWcr0PuAFVa73FYAOhIxLBpOI1cVClWxQdGsQL8xwm2vHGQrgovBFndhIw6VBymYB
zaNan7aMHaJlELl6XaYkYVjryoU8WBFUahUEIJFjKBR6rzRe0xTsHd1uw6lxDuUG2ZFbRxEusDOc
uzSd43DM6AW54pdxbnQeuRrzgsgMJP3cmNllSTS5gGsyCo4aKV7j2GBeWtPqoCQVGIt8a9SwMAIA
IxMOkmBtuO5reDaOLzL7kiOJxJhLX4DGIKXUnF9fy0aM8184oS6R6f9DqsNma+W8Q+BGwM3Wzzsv
3F5kysRCFmTR1TdtUUBXMWOOSCCWp7qMVM6eQEleMk2xYst4R2zBwaqwsfb+Ahus8RPfEEAw33B3
ZgZvjiDFChx5/LKLKk+GaJtHgqHzK8LZ1/zTDqb4fa5GMNVfVQcRVU/434D7AS3R0rFatMyCehg5
XMBelx9p7OiMGExEEDPfnHWM71Zk912VEhxgkezV8sVM8pHYHjPE8mp6Tvf9vW55metMLsbI6eW6
97MP59pfOX7P9zhtfuKdIfjpcItbgeZaYJdumdCdAp1ksqramS8XG6e4RSJL7JXfuqDkT+SXtq3E
aQs7YkGuHJJ0xWu4yCdbS34HYdBME28anc8RyRsPOtmwxH3NHi5eTOumB1RmzkSGeMI58iLLBoTB
wSXs/RYkRuww7BKuhmAeR4Y4BFitBzawc2WucIAXXS9haYk2NXcfbEPqpOggUHAYK9MQpH8yFarQ
3TA23A3K5xwpyGzYhKfDFR57OFEwgSTgY/sSHrAct87/pzsBa9c5iyAiCpTE/JTJdo3tDy1w0NLp
EyxZTAkQ2b8qrin4eSwkiq9h45IbBboR+3eGSp6PZWj7VAjKDdDFmC9fy/djGLMvpyqkbmUjz7DT
tTuQTxPWcXWPAalkMDRCwUPuCpfKczFUbDfI+696FsF1bQHBrN5SoSRRF2chBfF+8M9Vous01b/t
LiZ77tPiY9HZOsfcUhMn0N20Gztz9QCi6GVsfEa0W4v3Z+VB0SIjwhbPf7zFYh8MBgAQmSVjMW5f
5CzEp3YvlT1901/+pIRuyeTpLKfNRlpdCns0k+dkpo0WOUgGEesG5NpX4x8dyMqvurbQhwz8NIAq
9eAe2guykebCAryoJVRKRAVYih5I0Jo6zLQXIY11bpTOBywPdVipuHn0hFUxFHrMMvQGd7e0NKFX
2Rb2r0KqdUJ+LYn5XO8Rv43Iiv3IQ/f07JpK9GRIWzsGfyWQYysyG0qXqZb3vfRvRLgmNctPiq4U
ujHstD/5959rnrroSC7zdNvdiqjetiym2u5iB/skDms5STdXcz5WF6XxFMaWKtIc/whxrtQGOgNT
47YpXWyFtBFY/1RQLBpxFNuUdN8TRjuX/MDqw9ap1AQ25MOaOc8eHe2gvntCq8EDhOR7bnWLzndj
gfEFhL41aGWNJ0d+EGV6TZuzHfyO6MkH2IDTxiFyfs266IGrYdOE+9pVzgURQ8WvhPXHYYLXUPi3
j+TQwHQLZumm5WzyQVh8ihA7iquywxv4flZ53gmWkS+TRg6Kk1OSExC8QLSpEaL0QQP3yWSNqzzh
5gnHIhXKVRZ5h7OVR5ta/sQt95lqe1ShhsmfU6MwrdwCij3+OfPufjV1XAg9mfzSu1R/nuJnq0Fr
mpFu0fjSNfAg8yx8BB5z+cL3Z4Af25DgyAViTuI5MQzmcgVW7npbHiodhMVm8Vk4T3azc18svqAq
3F0hGblm9Kgc6ERL2M4yt3hVe9RrVdR87lk9XM+QxWeyyYvpRBsBbmz50k4OTdX7urNP/kj1j70y
pw+nnjjD9Zcm9Q3ryat1b5sFEGeX88g67Z2E62Ca7ikmD3OPQERmPssJKj7X+AAS+4rT4pmfBKN+
L3frfuiJiLi+3zSHvtJRsTva8JAm2b3plc5xGOu+C4qu6yHssPXyvkE1oJ++p+zRnF8N5NbhMPei
0Kh6r3q6lCbzj6HZQH4mlUzoQD3HDnq/b5cKG1lyIY8WBuMcziEJBQf3z/w+lnaas0MzHDzQgTsk
jVeYRzGJzJEa9hoGBwzwaPCMxipOJjOLG1MVmyhDaeSe/vr3+fnz6m+lHpmsfqXAqkBLnPwG0ugW
4X99yPf8tzfkNrydo4swjNH9d/Cb5jGEoBiFvkdDAa9FJmyWCBhQ+ff1ICbMA2QHwW4ulCd/Y7j5
W9DG4oMU9j+IyBkOiKNKr1jxewMnkhf94hktVuUcr5hxX1X+W3kTPk5wNcDx3+I3SjkrMboYcph1
yJLbUual0ZPBvfk+iSFcWzF1tbIuPNm91KtX3yLMjfbM+4p3lKACaPDoWKf7PVzbftWnRZdRqBUb
Wn2CSu/hslaeT8Q3uLoSPusYEU1avWXjNK7OjgmGhPGUdViwJ7SBsBKcHFsFJ9Jz+goqWsNw37sb
Ee+t6czi4uBI8Qle8IAZbVsZ19XSR/Eb12+nmfV+cCRnrONAgPRCccRaPZDynRXfJjnF0ACTRi89
A1wwArAUn/WHknYsVbtq5n+LhlnaB4qmOFnu73jG3RtII6SeXedtkk4j6XMjX420AeVhlHipH9I/
WUxNa4qnJl0iwyDoIJWSlUjzcobEXZiFw+v9R34cOTSQvvnRP+YUWdkFvjIxVvdBd21GK6mxdN6F
b61QeldrfKxCtyIzOd69up2O2vqnIfs+a8+pymuXAL8ROfiATrp4/OtZRUByLIbM29l1zHxxMOu6
2yZmOLlU/jvilbO5anCR7NjTRrtvqj3goX46qc65xpq+C7orME++ruxJEzAVLR4514ydrUwtChyE
ZYIUirqwWuH50GlCwZ6hOVHh58TYa7bw9hGs6co0EdvZsfp5oqHRgJ0HWP9eruSANOVCvfO6JJQd
QdCuYgXJlu6tp2bGNuTHQGgagHXJWj2OTXOoLp+uxP4v6cwYQ/HseS2a5AmSrAf8JZ/Dn/vZiGux
FtGytKj4IKzPbEliZ60Dch3a6WTMA3UXDtzNhFkOYauf0lA7SavlGu2B8VnINIxNkhVS5CA1r+hL
v3V8iefVbxEidi2e24GrdXxokALJ0DYuNdsGSK2KkLdz8kn4oBGsQ8dZVV/hAPqU8fFIRRZTy8UE
aUB6MviYCytqMQYDEbu2ycwW6dAJfyZk3fayLsIMxIpOTop6nnP+iqtKHGzOmwDG21D+Fi1qHmmz
C0SjHSOwtrumJ1Jk3XYluDqbGF3VgvwCw70amONCpIaJkTMkobt/keabp1ZZFxaiG30jwDV/SezN
n6a5p2xM8gy5ITLcxF367Bcpz4+ZbhRHDEsn9XlRHgx8LH5Hsxt4zQnIfFQOVt1vY7SI8+n4gnVS
17yiS8RMGXljEkTvmRn1nsP4+yOcIR+4KKAMP3M1ElGdovIAoaNwc/wQctPoVFvxIB4S7bHcUpf8
DaxcUPziDay/lmwDJDYcztaXWm8QlS5iXz6GUKjWrt9jhO6a2PNW/HTuwGBqFrc6cv66wAsLsHiq
ASsxaxHnwHIK4aJoev45O3R7IVT2kc3JB8NunO/3sk0c+XpoqZ2ray2nL8HSZ66ILwN5oMSePqCO
vWTyZiAtNbFhjPIrwj20bH5U/57IJqxkIHGiTketbWOn+J7uyK/IhGhsTcsMzaeiX4pdkI03YJ73
SeFqh8ky9gFBfyCXHVionhyo5hTmWPuWNJ5lkWd7794wgvqxvXvuRFh8uA3G6dvwPqeIxttzQ9op
or/PuACGglPWrcap8PhZpLM96/pgyQIorCyRUfpdp0Ea141zJBGViOakWim8nKmE0eVyHscIvnhf
lfa4UZxIViFo7bibraJsapWe+nd+HnmSzgT172A5jujS0nK26NwFeI9hVQGdkN0Cg4DeFcPUcym5
rPT20t75zmYszXs1K57ScnOT0tGI2FE7i1Ztx4zX0vaK+CjHqnuQZTwPJyP6nu3oxl71yYF/tM+K
WtxT3SotNZ+IikDswooIjthq2ToN5Ec/JXnCMSDggPeORL8OfDW4lqnkUmKtl92PfGpNwr5PpXUW
ARl8O/RUhOnLTaigcN3iMcUL5wt56xLOh8COucO9TbA3dwBVd+xB7d2UgLjOlMRhAw4y3qtR9kVT
PmudeReYroGAJqefGQWWsOI8Nst7aOzNjchO5oZpa885N+dyaEZ6T5VUuTDhqn5CY3bnON3EBjCg
VCzqE7yVBLKrenGd8l8G6J2Jfrn3TOte+wAoYh21lfXGKS/nftonCm2y4k1OsQFOiCh+1yxatywe
ZMd+9eVl+JsvS3Jq1VfE3L3TyOpfuR3EarAZpdY3VAMrd+YQqgFgwC2d3iT825d/RdidmTO6gO1p
Fdc57TUcWmGEPD5q/HuvDF6h71BJVSgQXhChLyOxxvo2yTqlgjTDANTvmwwQgPZYRoXm7h7r4A8c
WfnayK45XsvKJdu4QjK60iDzS6JY9Az0IMJcftlndUqC+owKeE586SiOChJ3NFoLkv2Ue+j/9tmM
mDkqESjn39d1trQk/Tv+JDquXBDozeleDj7UgSGh8Zxmk2PlcDLaQyOKXznxn0gjHFnOS5pPIf8J
mjCDvG0v5TDw5GLT1LvACPosLGQafK1NmdkclPtnUkE3jS5cqtvps+Y4Fre6w+eFf82o5flBPU0J
vN24+TCqfJMcRzmnWqoD4vjUatEMziU/RG3nehJnOF+w74QgXBN8kSiMDPfIbKJzulN7K6NcxwgL
c5Y9jRc+uOg8Ufhyka6AxhXXUCN2D5DutxVxOLCT8EPVw4Bj15X/S/aco1pvBIOSzKu7xj/d1TMq
YMP2T04wI1sYegqS6i2veHU+nUv1Vt/xnVaWbzON1plU/r8tgnZy3hu7jDQaN3dZUhQfkZ9NenE/
2mOGZt0P3vXvy2rAw8fd5SyQpgtybkZVpbJjxxqTWeA/ynPv3kTfbGpIh/5LMrPUUp4duNtJ3Ieo
LU6l2tOm8TGwYlmNPlOKRqzKxVrNlqK5XmzoP01ltpgvkudT81q7QPBNXJrOaXFiSZJyq/InnYG9
umVd1K76t/h5lGcmn3mb7D4oYAauC+nwJxlQD59iF9l2NWOQ6VvZhSiFYazyDDLrpLKhNOV0+2oK
8gNvv5lJ21QfPkKmbiYy3k4zJYJ2kXmpZz1ItcrEpP8Yc1t6nO9pfBQj9eiaCV1TU9AOAbsxVzyz
XqWTLqenmv431BjNPuFY65ZRXJOhOhu0CuV2I3fJ6KMSsy8hJQV0VMY5CCGdrGFfUo9dGF6JO5fV
bARnkCaG5V9+lZpVG6mwruTc29+NDzBAolkaCoAJEm4ZIoe7Yu741eU0ftiHnni+KMmsKSonwsyz
OXvHFoLJel1V5nNhqyegYXjgyCZ4VpYcDS9LgLzpZTWj3528m0J4Kf3qM6xx7FCjuER3XhEUy3wY
VFgA2rXA4gCNzpqrD1824gNNC6mr/MvvhUCHnxnoEOnbg9aIjkHtkAOrXhBJn7J3N/aQNsw6JUga
86Mt3zV90J0p1djw7V0J7EoCVeV0Q67HC5ekz8GGa782cEbWVvYVZIrNzBgsw/jGIXR/dDUqkRuJ
xBWmgQdtN6VNlHYBxBIGxRYSSdaNhGmsMurN2Dr3DNaK+94lohfiypvZOcOtNDZXkDGgq+siHe70
1+kRSNMPTXdype0fEKc0wS7EsrvBrly/g2OS+IFvkcrULbrUxuZFfUQqtZzuB/SbTJmel/N7D7WS
vDxg2wlSM5cdwCt1Pi3dfL52sdL9lIigOgeCMDNYAgRkrnw7xQ/cAhC5fpZxYzV7vMC+YpJePk+Q
fN7UK/U+z9jNNTl1tSn/2txiq4C+2OdH0PeSvSAE8onZ/ZZTiR1ojaFLeAnTGxrJuqJ4efVVFgW+
Md8DE4ZDFvkuHNu11z+3s6zr0fjYkzWIGB+SD3m/1HhzpdNuTwBkHHiJ9MDegEcrSvYsVSb00Z5G
vThaZo7xBKISzBHRKdm4NZCTfz7ByH/W77JPq6yviz9Df2GCJWYfMsxRZn3UdIOpLE15QsAcpNZi
L8YOiAaQ8r0xlOval2W9xuabQfRsdIQRcX9xlIo8ZyItxQ9cBC1vgsBp4ZkvL84VvU1YDRgaeBdt
QajjIDe877RlI6lFv7pT15cnxWTnkHWZ7bW5LrE7AR2/qoGNXNrQ9NQ2DU2Abwt+kIvmwM5nodMY
0xCLoPzbpO1hrjnvon4C+vDjMgi69x44RMwPir/E+26/HMf6rbSIFldidIwwf27ymsX0NYmMMGdl
cjRwmPKaP6r43Zp4XF8yXxz4dH2PQaUA7MZ4K7uPEwM3chrvs37/ICcNLVE+sAGY17WBcN+w1DlR
gbjeE7gKrFrXtyM0FLzQft3R9Nv9rcKRsyZMnXjgxe/AWWLHB/FaAtbj/rlM5idLF5ha40H19sAi
jkKT0aYhDUXYQVX7dAIFaw9TpddVmZZkRDni2cyXOeTNidiKQLn+X0iv8kvoWpmTeTtQYUVansu4
vrAw0lAwWRhMfalu4688t8OLdPMHRpwMvZVKvPzCJ34Trx8ry+1SwXKlGKr3aGEJ0VrlHv8kcmlY
xcLsgovLYY2DewHJD0yX5pMDkjZk6H0ANQqtwnAj9sqkzjDS7XYbZlI85oKdpOoE3mG5eUxDNpek
zKXI2MWFiInvqqo3QmThuKgrnBjijO7/50BAEvNYP0yk4t+9An1rw4XHjyxCKy16bStqFW5oqmt3
Guiz28lkyt+2ed6rsH+CrdZvJgrQTyf6Rl1UNZP1fMyD6ZpN4CFJFHwm2uRhYgh1H7/BkVcY/WPf
hAOcgddXh32r6xYvx1wLl1gg8Z8kGWV6v4igA47T2yZaYR5D4T4PE0yw0GVwhUuZAIulCjS5Ysrn
Y+7ShBKAYGge594IUAYIrQ2EDLLc5faSvYYIDO/0ELvMdrp0Fi1zLHayDd2E/WwUb4QBdr4z38hs
ST1UyCiHjuHxCBwRiz1nd1peueMgwJfFHiLY4MD19ycqA1/f+Zc6pSRv4GHxrINhTNDKlLrENPaV
WYJMba9vfD2wk7dtfFt+SOlNAVVqBXyY3vBZT+0QQII//gIbmix8YqAlyEW9cUszuNdr/npCDZI5
XQVaSyphrx43mq2wwzoCNPTi2kZSKn97IAWV/8DD0Oe1ybOke0mZwtSM535zbTiqEhNs/KNZJWrt
9fT4nIb3RYvrTiQtg6ruoapvoIKRdG8A91Eg+BNIMHUL+SN0MI99kd6YdqmVZ6deEOoSqiBpvs4r
lA0cJ+MovfVtvQ8NsZ/BdE94U7T2Q+GTIMzJGm9K8pzrf+ZxmK9N2i/cysdrCVjKiMaPvUuhgLVo
dIGkuNlJzi1Yyk+1jsEqdYlLk1uIcOKv7IZDtWg/rGAJZ4UDb8jkFOSUf2CVAeuqZ90EXS1I00hU
kNrlg2qhiiU9iP2mde1cIXleXA287jKdosWYLRfmx/9Ls0ssDFk9SSB6M4EyxWhuUBp9zY/tlvhC
mLJ6g/lsQRDjXuQibNnCE/Ng/9JwP6iaP+G4UfoLe+Dd+gnncs5fMjuFrER4WG8h6Clieod2tEF0
4lq5kg7RrNuhU02PYXbztCnaT/ss2HCSI2sQe1jPo/TSrXPsFN+nvBs8JGQ3roGk18kuCjVnSUfx
IE3AD3VSaV6xyyVG6AGbKNVnaL1zK5QyMBFoXWpeHmC2HPqm6qA3pIXiXvJ5n6NAaD0VNgigyt9K
fLNgYpAGLllcSre3J4WM4mGW7lVZANKGPKtF6rz+i+JejkcbPRoAMVVWFTe2+OX1GfRX3/xuSjuw
OTTa6sAVYFB7KNuqK2wH4Dqz4DCXnftiZc4UYAYi9BpUBh+ggrigezLcA+17nHxitohAvtooraCO
iDJ1POfgdXMYqfyCSFQuF2gryufkEbyutc3I9elMdp5PyTzWbi1H2Hj7Hf1MdbsuUq0z8IyMYD7Y
JSwhLX3+14BCM9F6z0IMXXam/5pNHwzrMOlOWzuD6N2mDPswanlBml9rFlMSeCLehmnayc/MuKfX
LxGEVfsp6QGR2+FHsJMfYH3PzISY3ODASwbbo5ZNektFeRaGXveHUmP5MdDhagRjKARR3SoLMKWm
CmfCH4VlSPQf1ci06iyzoes1pp4hiIKX/cVlHF/0CSBs+ck0xwauu+lQvoMLHFI7D0Sh0CoWrgHR
2mjs2ZnGYR8HX7oYHwy5fZ4J3upP8tYS6wIVHxe8cM4ylGMNEhI8LPLHoANYZZOqrLRKhH3AWIrO
teGsf0/UIWh28Y2Owb25mshmariK787BfkD3gV9s1tKK2PMdSgI8YQSk47GLldBsNMEyaX1sHESX
ERwAk3YVQInSFodpDQS4LdzVaVUvOr5PVA/DQzxTfK8qxsQOaVuE9MXyIyGm/knBY4jC0XiLzjqH
RkB8RzDlERnKWZh7E350yZCom5VRZu1fgUdfPjLSqN6BFUUxzeyjlxd3CmWtl7M6VJwQm2+87geW
qD8CIRMT+d1P/SZDXU6/+tqjVVC34sJQ9OTUxYEotcShz679f0M0n+Rjv1BMSBlVL6QLhQsva3fj
JnPwPprhvVzlQtt0b8QKKR74ZD8T4ds+rJNfR/JaNT/5/UTL36RKhVx1XrEIhcleFioiRMSsQhWZ
zanLAYe/i+54muqkZKBX1LDvVX6c6KXzRzrWxgc0PKzzk3VqwrTvfKqI/rf+W6kr4H9CUeSJBI0U
kD/yYvD74V+/Vr14ar2QsI3uC92EBLUSM+9neNm6CFVu0qnzgB98H11aUIRSeG+qSvlm+Mc6yDLE
tFHnuJo6U1JyanYanW1iTan+GXw4tu21RksTS77p4V9A20xOsDvE7h5IDj098U9GLvmdL55h3myj
Ge2bKh8O0qS3KwqAFcMBUQqpb3lbwFHywyyJ/DDanDkhkDNfP0IXEIkMFNa4ppZW0Wi1PS3yQmST
sIL/r6TL3RBNJl20IupBk0GaJboGL+6yuFKN9Ag5IOz3iYFddjGIi1viOQ6Dbfs6pVT51ornSGa9
Xbd1CfvSwHTL5m1T2ZilayCpmfAaEuLrY5ooZfO6BCGrevenQZXkz6skICOoSgUcrz0GLXWZvvaI
KOOIb5tvqGWLtlOILzOqFzhYrFCSAeo8+obrKDt7CJrf0daat4kLiQur5SZmooLn2EdtlDn6/REE
YA5dfz5ODD52y8zrMstg2MhVWypJMc4Mtdtwc0H8NreRi0MiaZ7o11A2v+Hvj5QzhunWCRMiXuLm
Lzrhijo3ikm090o3YFFA7kgfurWbjmkg0kSJreNfEg0LbXAewZc/8/tUu0JECAzTAAfbyjoTdYzc
IctmQ/fVMSQjHd8ToolO3aCaEfsS1lZlFVud7vtBamUov3GGG3w/5RQfCmVARTB7cMO2i8cKpMLC
Fg78bAtsUwa6a19w7FQ1YbkiXm4ea3vWguYBG76OHkVZDwHawFceZOrXWMGa3MOXsbJUKAxRacqV
K9hw5uCzpwhT9rBO2ifjL521uhlK2onqMM2eJPNgMA387isUwhacII++o9wyfUfrzwWqAK8GLIn1
ga8gf3KWEPSOrtMrnK3EFIYndbx2mxvQlVwYqP7duRLvo73mCiVmF6/nG2/hc4JUU0NcEFfS+j4b
D3G5avKAyjRU+Mc3stsh4r0nrudNGLtZAEPg/up0hXIGx79IsOUlKAGNwBPeqTDvLcfNdZ+jT1M9
atTckCwU+IZRyHOLoCDOumxeWFUrGQ3kL0NThHqE7DszT+XmC6fSpZ8tAs9zluO1TOk0ZtgK8KWq
8AQGwxf31QNnb2DistDVMwvmfOQeO0YtNcg7+FngeC7SGwcpg6rCnwY9G+pYKYM+Yaqjz2x6RLMq
jTZzJYGEc44gaxJZpVEHlkY9Rc7LoKJPqH9LAou8IDtAGUnTDg9ar7Sgu14TKLbpX4n5HkRWEBXH
S3/KyDFDzhkMg78SXrUiaqYiNwS7tAPk23Vxi44t69/+e2mVRBikVKPCMB+lxFpkQ06tTYHUtSQz
JiY4NAvaiVhHFeAMmo+oHH0KLfE0c+qTffiY289ppKxY9zfcFeMspMtMXzSG7l09kFZFKGm6wJGo
mJq40SvpcCmMplzXwfk9lCRmbiOvADooDVxDPTj7qjonUOdifk8+CSDVxux6/qnNYkaFNA5jiW9D
jVQhJx/8tP76Tr0KSAu4/8n8b+mBUMmVCVMqawEujxVWx9gp8StlZpEqHzkZRUkyUUWlMK0du38C
sUQhh2wdqmAZKsmZUuIBnodNJ5eSmmTJMvn48QKq/i7yfEMYy8rGHfjK4SiBLbMkjTq/cDdh4L/0
EjIE2w4bHwpJLcovmCpbzjzSWgQ6H+wiqeWkyjABRszUvYOTV2/XiUnntrAYrRtzrisk/FRwLWke
AR+aBthc0fBxToXdluIl4qFnxUrmdlWvWLqlqK8TLCDPLswcmTzPxFZrJPq2ZqS8IQ7azSMfx686
VM3nQ0hZVvHkmhzjyLNrOuH02M48juQ3ebUH2ev6Q6ZLN01zpHP+6whyMXSeSqyv9Oigg+11n5E6
tPelYaKqyN6AFQ1ahWnYAlyMjDBw2r1Zt4vFxmb48YUWAgv/y2Go3UfFvq/jIc6w+1G/q4/ZP+aY
B28aj97sX9zpQBTDSaIWe0f8DAP+83wZO75S7HcRGbNbKLIogoFirtof3+Xe0UvePjICNaKC7hVG
u8ZkirR9jUh2eDzYROBEvpgD3RwYS1tEx/9i6+B3w+HtEc/0thi9+zMRcHTV9SqvjQQ4PYExHoJG
n49ySuBJe7OlxE6nDS0Q4KBFgSwThTn2ECXsz2byLXqYfA052vPBWQVnCDTz723jUzNNDzKh4wxR
9kvKLWZDPM9XCoUVYa+ElZREDTbSv6JMMK5+BSKVacZKpOtJT1D2B37kDmbfomN9eSHHOAT/fxEs
EworqUUscXISaA/j/pL/iv72NGUKLfHXdC898fjsKeDaVwfjeAF4PCGNLYwi/yH/nsPkGIncH11C
c6K0XX0leCN5E7TUBrmMGi71NXtg3VAQohnOQo+fq5Kxh6HPEiHE98yCfSpya4ZY49D5Ffes+zU/
J0Qh9iqS3JQ/wx50HMUitO52SctCiQHLo6oKP5eyFXC7SXeeQfOZ5zKUkcsv27/i5ZBMwf5pW7W1
pEWmph+5JVAM7LJ2CvMIbMW94LBSsjFg2mtZz2mguM0a7PtGLZKK97RPSXqnnzD/I2qsb+IZsk+S
webxLNVXP3Vnvnyt3Ywg7bFylXCYI2eDC3O4ZiCtreA3Z+b9UTGAqn44cb20FK0kNhvzRC/c4f39
bCKV0VUY8TEYs3mzvMSy2HRi6+QJNyJyktP6TyXLh3OA/JKeIiInNrz1uxbYxzO0oMrEagrips5f
ONc/6BroWTlKGd5qizr2BZBrrgcQYG8sM7MNdEfHldW7N2nNY1tuPRT+TBOf7XWA/N+N1FNmPini
FaybQ40h2TcXrsoibMmh55GGjb0+otyAX7h6HOvkFV4bTWWtLeKiPH9e6JePOd8OK0/8UJ/1H/uO
Ny2tZ9cFAMoPqsU0kvQmoVUzShq0tVWjatQ/xNmMjl1+zF46JFnUzEUrI8PKdLkJguCgMrNeRuwW
FAllZD+ZMoG6aEBQaaxj7DyYgGThC8tNpqz2tGD3XSfvBjKy1tqsuGh5bH/ess0htHPIqtSibyvr
f1iDyIcHSFDEmDpObtAB2Oh30CD48ICd+QCXML51n7iF+2tyXHk4tbAp3Ecis1EP9Ua3NBA24VOY
FjMOdKTtJbMdrvonrJvxb3dTCits52MwqDEQNHjYIbZWijHoUpaz+q4TZKyMZys2oU7lY2orXmBV
uVOW21l8Vs6TUPlp4t2nCppvYcZQNAWndW/qeJMYDfpM92e7bOfJMQxilTS4LMxirSu4rNRV0cpU
C2G95AuO03uYixLVam+SLGsBQk8RacElDw1iki+VX58+7YOE+EzzaT3l3mDVQpHGUstXDZI0JNe3
Rc9I1CiLkRE0wVkud6A1+LtaoKtZnM/IFADD6SCVsa5keROwkmIiEs5np0Ly7x+3dZWJIYd1tc4+
UVKcRsoA0eTGpdajSp79kO3kMRj40RHbV7ZtJ8+Vjxu4GBjOLVSxIzVqHXqXlTH0joxBUbaNhbZr
OJVbCD5gnqS5ioxSs+/B9iGrdjRdN3VFb5aNWEB4R4+NGllgYSeL/z+uzW9fSgAghFsa2lbi7lGl
zKW4ZslGMXW6DI5J3Xh3gv6NKfCR20ElY868euJVOjxwzMyhFQ23y5r3HsjMeSp0zoQazW3OsBwh
hPsKx/qydq3/FP7MCaY6Ovj+Hz9A+4GhonCvpqI12NfdcdwAEGkFmKIE5ddd/jzJ+kHkESVQmG4R
C/mMfiGUkYFEFl7gM0c4xDe05sYRl84RpcNDGL4NDGFIBrL19YY/t8girvFHiDMbs583KlRa3lEk
7iZzlG1Ui9ElTCCle9UnaEC9Eu0gmV+yx5ZCXfOXmhPyTd7tbI7swIFhxt+3cL2wMPNaag6OzqTU
LBr1vWu539glago98yiJng10wGWJ6DqdXOx9tRJTZRJmWlzjcsSZFlPmqlygp1QHVAqljaiX/Eqm
pAw9HPt/4UKcCBJhMCYsYOLWbYJ53LQD9wAlpxBlAUfwTbBN2xplnq9KdJiEqQWL48gMf0AdCpOe
zUYHpc2i1ik+5g25ZtQ32H78DJTUUvRfmXOJyRs4nF9dx8+625MJAZ5m1/DMFnhK90hON1R21NhG
d3g8w7bQVYdN/OaOO/7gsnQFz6CAj01NkPXB72FGq/FzQ5H9MxhPjScLo0+X1Q6KoCOU7QF2yOjq
9ZX2i8O/U5nT11dLehjRskpjvupH0YVEksdx5+2RPBuPa1zFWB6Zk/HY/SKhz9ByIuTET0ownAXS
5Og1Q6o6GFta8pZ7KOdamJoNYAfYGMNdANtVKvgkjWORgu7dILaOwmASw56HOxQxU1B3qVFObqnx
1YN0n4nBhoB9fl2LALbkB2wXR0U+gs40DJYps1W9twsVl0pLbto/7nJL9/OnRK4tHB3ySzzGetkh
0GyfpzdE8iFNeU87WSFZJu0K8An0gijI6AUcFU3W0YqxsCAzReYfCEOUE89nrQBfA4yI7lVlC84n
Ex+wf0LzrbnkCUd6BXcYZmcnrAPlBcOmHV/kxU74etvsdpcSOJ+m9TgbDft4C0q3KHkkbCWeCPyI
q9rm8PztJrwOgiciPpMP5yFXS3Y1v+B6LnwMbYQ0wxyLLn8QWp2uPS4+Iq2zpklb7oQa0OcXp7x/
uySHNBO5Y8xBHw2CdQ0Mp8fuQJ8qR3u2tZVtde3H+oPq5rjFF62EOymUbCOTzknchDGLiO3BDEbH
06VIGYWoOmZ3P+lZiseho/1kqtX1D4gLGgUlB2z5W/yFlZv4zuSnoCDxRuKiZCUWMAiVGCTNYJzQ
WKmRVCjDYciLT0JGM7jLqCwfgfCuh7NwJQemxeUPy/e+bm+k7BiBHqMxspaj5lPrmtesIFyr9Eea
tm3g0ATuofX6SEyKinhr3KC/T0SqWjK0sHQLkjno39tIg209/ySt18yFuacoEvSU5Y0+pX7ZNJun
w+dglDeDdKcZu2uJmGxO+iMzOyjQ2833teZ8+R8Ne1imF3pSZ0N8/B15uWrmi2LkNIV7UutJcqkN
KoL1vVWu+opoQo4fnZMMVCCXDSqTzSplAYmniahD1c+uUceQmd/YEnFVZbXIkkVa/PWXMVTjMxWP
4aDMFmiB00PI7xmNwDS+Tz9nENqEo2NsqkLeagURfLIgyWPyWtY7DMxg4GHdzhw8ULlPnpF3DNRc
NksqANJBh0ZgecliNWikKTwcw1wNoss/XcVxlRjV4jjHrk6cHEqgrE3EMrbacG9BKValV8QBUZfP
OQvQ2Cg5t8FlTXvJ0b/wRDkAAksUYNnmWwHwtM3vELUw4R2jp6cDP1pcEbAUJn+76lvQpZ7MYKSg
tfI74/I+ZvNb8Whn3l+KUFkvP55197rsJ87tVP5B159jfYJBXSJ9V1KhYtWOJp4B24AdmUnfJUHe
1n8NMNzay7i9nWjQGsoV0/7vJI8cvPhi4NrHSsemPNLOjXyTXlRnryP5IOe5SzJFn3J702yRdLQE
knKUh9iE+zCRsclOwq6bVBI0U0mUOAVqfeF0PqiUYerWkv6CEkMTcJl0C5G5InQX2l6o6F3bVv5T
0gNapT3k6N8Avel6URQkdONnExSlS2ZvQyMjkzww81M2SlTKLlbDjKh4kZiGHQt5n3EyvH6JeLpT
JL0X5hQ4cOpVaHuyh85bVwwuOf0bZT9GooYbS4k5vPrAWpjNmATNfQXOb8IyN220HbqkVIntvJho
aSAKlTkNQX18dTHOY/XOgQqb+fjMVQwfrWaT4xB3KkUbOMZtKCPuKF4t+EvrbT5FxgsKmtn91fDN
WRVJj0oM7yFqVloMYbpVv1C2P6jYMNbXTb4cjPHHV8c/sBiiGGOeEIEvM1Yxh5e8Gi2oJZUBx90d
ycR4OK1wFVkCYzfd3cfYHJbK8GpvTo6SUAcVgaaS6DcogCAIZ55YLhrPkoPOwW5c6sTZlK8PwgJ5
3RKrhXK2aCysttWtb91+Ennnt87l87V2F4EbFpZOZ5NmZSouPn7WYcexsSTzdqcG4SmI1TVMMraj
Bga54gJoRJNkGoJfSaizft9NqyhBfdQigLDvj6aOhN+Qs4rwQ9M3wMe4zNGg/suFWApCs9qZzsBj
pEEuUVrWa5NSbcZqH4M/VngUYatMvMJ7GuPS4/EwIHtLogTRdRmTApL3wDtCR0LqCLoQ6IQhbD/H
M+JjUyXxFSjASnvS7MTRH3IAGGf6SOKaYvWGZlhBvEF6d+BIrygkDSBkgFNHALbBriOVNRCNmSSk
Mgy7Elhlw1bmUbAx/6Uo4n/h9G4vJUk9vFGbrlTQrwSyIYe9d3B/nmilWmTy21E+uwPF1R8i0XmA
CAx2HvuxYgORcD+KXphfkKtvBypUSRoAJEbyPL9XmOURjJe1GOGuZqbQX5XAQ+2xNNOTRD2gBG0P
lMDU2H6kBbTV/w2aQ8j+0ZOKilq23wut9/f6oaQQ6rZI1T9lAR+/T6bTneb7VLsGL0bT6SnFK3QF
+NJmGyDj0D9QOsGLe4wI6tvpWdsxPMhjtnDMwYMtKutPv2PlgDNE6CHBuECcHrIQIvamrc06maTC
hIXrnf0rKMNyYVCCPhT4c2Hs1oea+AI2FRGfgsMLQiNy1GQOEDg/o3jwb3HGxiJ80zt5f4EzybnD
xE1Y/jfULczj+lJSmIXHQemBmpGvUHk4j7YpGo8nFJULwb7A6IR4v3pHx6yr+nXNQGrlMzsWffn9
tNLhqvkgjQWgJk7UNm5zJSiBuirxGxmj/i8lCrxg47V76wNtkVjyZxggcsdsusAofgUu7Anug/sf
SfEyzJh7twxUePHpxrEsEBEtEWyf4d7iGVhI0scb5xLTOlCWlctitXePUuSfBT1he2zQIQUV4YWB
7YFsWCccfawBL9gwdtNaDyIL9uYfd0lLPBURDgvK2UyaCbh424IpMJDLKPoSGyLeq1/Tcic1Gzw/
nGk0IUQxiEqu5AKDF2pZgnXDpOpsYmAe9LbBL2aZMDJcREJBoWEaF8LbZK+jpFzb5zQgnJ4MY65P
ruwZI1s+trLddnX6lFXKJTivdRygURs1Rmgc3ICOiTbLkkl2/tY7P9d/4HV1vqg/5UTUOenf4PwM
wvjF5F0GHx11FwHfC9KFejR2qUGTApdRwQNiN6vmZlUNWlEot1OyRvYtxB4ege2GgbI0j9ZDijJ0
hBDXQRjOWLVvejDbU2ajcoNytkWv3ecsZN/eU6L104ZjyjL4XoQzGSMFAApaGz/WzNF3VrkOn8jY
UxLUguiW8fYDR8yGIQYYU1lWTJ6YdFfP1/X7FfYgHLjPdbSMEXpn0FojRvOb2IzutQ0e0WvUc3Yf
AiWQpCf9+pdhQ9Qe7P6sgNh/lJKClu49JdoEocLi0xIHuxmOPFH5VYTkV9gbi6VqjJ5nKktGjDGW
wGfZZIA5hznuZ+orbod2b27zBUNecxKQziGP8LVvPUQXz30ivtzbf5C8YUmfwCw/Z0zUFRRMTxD4
u64EhTIfBUYlXhE8DN0eV1wMsGdJhY0Xmw1oGJy1+Q9VP1HBKbxmbmwl5HmbKmNXFg+X9uyEcwSn
WP2duSlnJS4zjVda/9tHzwLJsSujYJzMKy+zvpSWPWDAaDza79s/9Sc1VavIZGSs8fJEmZEyY6Vm
h9LRXf5qsRH52Ha7iIBolJ1qHfDkbwrtPXcASxYTCtIjrfMFchomYw8o/PII6jrDLniORgbloufJ
YR0LeXf8VKzu2vq1y5MlaS04MGZy+9R3S+oF3SKrIuZtsAdudc4aqu6gIu6Z4EujNfYmJNoFqGw4
OflIQx3orLdC22se6No+JqH2QfvRgx0VkopyVHiW1e2BpMgZbhQG68jxAv6PJ/PatXhxScaJ8N3K
IbRwP9GCsICcVDuXZSc4vG0KK5GLgsgZQv35OrZXNcFJEJjb020cxRMa+9MrD9GXRsi+od6jObBC
gDqIid2u+zkpiSqNXlZoBFERONEc9G3XjNJcSXe5WsV6aGRXT0qUiwrwKiGqYjmxN5vYc69C0JeF
HckWYQudiv0g5R5pRlKiiBTbYXk836JgcdMJkhaPwwtK0CxjosK7IErYrdeRHPCwa10bg/1TVIuB
jAfJpElYaF9UiD6eU6riwwJAlOLGnpCCBTsMeg7q9S5JcUa5melYxG6JJ2cpvWrj7lqYtJfX3PO6
1ENFovcVdNiiBI5y5o7txUxj9cYR1Og9ghKxDd51Pyect5nBpCQnebRyKGwP4qp3jnUq3SYKIJ/l
UTMO89C6v5L2HVqZrQ6WaYWrHDj3OOt4mmaOyUYqwvfN/O3RqXMf/scgU6TZKW9bspeN2nOIa3bw
UcAH1xJjYBqsQyV3kHu3Ex4l5VGTsfV9Jya8N7TMWpwakGWsDoZ+s8SZ4UriPiNsaoo7ddcRBCli
Qos5J/VXDZ5eAh3HcYByL+KSJ5EsF4wdfdryMnA0EEaLAehTDxIPMu/XTiFURESThLxouAM2lInE
cdle4kaIpSfoT45Ka1wONhOojYdTwVEsRsYSa7pHjnVR0md03k8IwR5KcMllK1B3zzWJizHab9u1
nyzOuFUkQXKKESmmlw/Am5GO9x+yOv/yxixQTXp7D/2o2P+v01aQJ+E5Ldb2wkpHmLLgQx2k4dj7
iaO1pt6upmmzBl7b+gUoFiNel5YAsKurTGJv+2IXY00LGzF2GPUtdd1/JkQ0GAArJKglmyPKXr42
IxR4x//R5pOO1kvH8sZSRQNw3wNWMkAVshhoCOu/YFNp/fNd/3MUnYAfpERWf1yD4YDxnNtml5Nb
g2adakf8M/Zp0dzprNj/ScXw98KLlNXWZjFZYcRpAWm7xXTCAnMkkaY30qlnVdPVPcc1W6caVAnV
YNlAyggMQyg43DiuUkTHsMCQmrKadLTOApctecVdJx9CB58NT8LRT57Ilm2/P/7cf6p577Ca/Ram
AXULnN9reTmtVUHpggVyKblSKEHFDzk4edZIqf/Dyb6uia4g5QeV+7U4+Otf1xop74pu0JWtZsUC
0Mf7V7MPcf4gpOrout4rpVfRh3eXsQrfd/w0fS4tUi9cWGO7eZILkAsPNeSdndubcZOPD27Cp6hE
3O8fwW492y9WycqAq9Tojnt8Bk+2e/N7VCf54kqtBZxMOPwS7EV27/CzjIEdxBHw7W2/eyeh42XQ
F7/qItF7GRxD3nA8yT9wcZ1UPjxd59BaRPy4S6zjS5XLnMpj0y0rkqiQcqE+oHy7O2mo5Zf9LLFk
snqwuG/x5AbmWgPqUb2kBxCsvBIb//5KhPGf3Et/6LydKvi3TN8at+H0uyH1f8e++b9+IQtD+66c
rX9H3NClpjjq+RrxTCR47/QnFZF4itXgZr15rCX//mlrX4zNSbpmUEcUDJb/G27jCzt1ZY0YPSMe
iCGDp7bJUyd0dTDUQy0fxwTGvEgkf3cX63Jrl8UDQxcAiIV7t8fJ3O/U8jrqQtwcA+0fmGDpNk9I
AUlfYtnw7T0GYEIQ0Avu2Lmn13KuwFb5a8NCHvPQfzxEv0fDILz6IkkN5xW7FhaqpQA7+Ior1V9o
8iPf9ISPqnRxOgEreboyVmLqvQuKGIfIMKvDLMHGhj+3qt07iWpD9aLN+mvuhuI08Tv55NcylMnt
gbOQJcKbyzC/mkPY73WIHyLf2/1fx0JwPXE0TCZING2CQXd4/erOsUPkI1xQiJImMzn9wY66L1DN
R8sdZl+YkeCHa2gEWdRtUNu1AEtvpf/XoMRRocgd81cgm+oPTpQWf65QLUJfaKCTGxKuCxVBhWlV
ozd4BaGMbdxCEHHK7vEznbpq92jGzhgSMj8glxN0Y8qZtvoiprVmE6DEKmQeVByG8ME2anoWZBwm
OwhkMy/qmqaNry1nqv49Sh3vvMEOAh4D+QDW0QJEpFIqGvWN0rQcvQ6zs5y5bt5zgYRJSgb0Vc4J
gl9l+lx1LenL02GXXDtwNih4IJc/+wRQLAsNW5xPwRRhS8J7iEiJbm4CMEKDqgOAWriCpYG5Ev6p
NJAdHb7elVHX+enydjSNKBXrrZyExljsr1RrGaZJfLDGcvkN45HW87QMBTA7g5RM1Gq5h0n0spkz
532UO7ZsNrjhMexvQR6PR0ARV4mMMqWDZH4eFps/+MgcmIIDG5WqZ1SgHOSkH0fuXwMsf5B4VtqQ
G4BR2Afm2+hyAOkLLn5+zzCTrhv4UopfVVd4ntaNLGSwVTqiYCfaQepepU1V1I4y6KpLTffpuaZM
nioZLE+Dzh518M+qeS+o86/3cyPWRwPA4CNdqTKzzTJ1Czp0v0Ga3hHNM5PExD9y3evfBW1ztEhP
MsoN1QoTWGbhSY9VSU+kpxWod7+Q9XmoNOLyuE3GIu8f3zdUAmc0IF3gJJ8X3MO0GSk/nBJK2Fup
7Prs3qv1RtN124ya6hrozHFCxcrMZXzmgzKUSulZzLZVFk9w52XVSfbeoK99E/jHt3UKXNX8B9Y1
eUpuNlL63NAP2pdArLQS+przh0O2v+daKfVQ6H2lIkANCPCgN4ZY5cXoHbTwl06U2pbPZ+14smak
hiPf6esn3nxfenmRRHCCM882PvzgFjckhaVT3NaVC26mTgLSYLQwA9OLWV7SXMdpMbDOq49Cab+R
RF8IXa9KZwxTT2ODojWUCc899zu6XVy5CUj8Pib1TEQE2SWxt7xtdX2kHJI7hFbAnpuEKuCOUCqq
jo0mJcAq/wju5qxfiycq6/8p7DqAabyx6rEf1M7V1VYiAHSd4V/A95hAONGYHhYEIW+i/HDC5uNf
ipdYNTIUPTxIgl4gCsZxmeZv03DSn8HbK3wg4eZvOh9HnmZ4MBiiT8Rlg6a3oX9w8EbOqPmOouKd
EecuLrmAaHOGDo/CwittnjbuMzW6uB0hFt/014b4W0odElzEIYKfusc0ZMNeEtWWL2Xg6SUyuQ0y
7hXhgJoGy+cFMrJMduZxFtn3stxyuf6hPMESci5jxvQruXDY9kH8xbKKaruIp+Xp4KhADF5JhGbn
bh5KwMZmNXQm1lXSNKwlLhRRc52Svyk8wDzIUk4CtAw5vUGvAXKB6NBijd1jAJHUGPUbLf2lr1wL
bCIKtePaO1tudFjIkzxukDHP2s2V09G7AQ4jyGwr28zZkjgJKQmudbAbXj+DwwNJ2M34yVxLQew2
56Ar8oYteohVLThT0W99NstlPPnq/8LqwSEIENUWFiVruQ9rrp4ZzwEoMjbPo+ZEbeWaFaEbaloS
l6J5ulaeqkCMfJ58G7JAM7iTWdM34PnkavLG19BkjQyardATXa6vaj4+ohiMfPgTCguH3/mHdEwo
lTz9JIr3CBhOJBqGNJXIMhHrJVlIzpHIDxr+noJ/9wLjLQ4vBOinje0srrgK3ShCAv5tJO+CVysL
xRFC2fhOw3cUCy6eHhhRXZVCF6cVhi6WFxEwLoy5vIf2glSIus7vSUjjYW3/zE41Ouly3NQKXYVj
13xH77mnx29XoHbWon+zD3H1BK2Tx8s6SmCCJEcBOuod0GOWjxASX+l4dFY/SVA4TUy+O2xrvdy+
KiuGnndrpZssxOQdwVlVqVCsr3PMW8FeMQB8br2XH+PI9qvlBXiGkkh2DG6qOgl3rOy8mVVRldSl
xY118PZsHzFVGL4FbHVBYkvjiZCI0S3yXVK6slO4XXJHlZJU6brgyqy8mo7agEF/74b0wnb+N4rd
gac2hYfQMfvv+O4870leInWgWrV6TeGKHSItPsIaV41wkfievtJdy5/wZqv4o/8QQrdgdCzic1hv
I+nU2F6HumX6+yji05RbWRljMdJpLR6N4lAmbSR5fNN9TwE7ZRyPbuRTBl3916VRsyRwU8RqcSGF
Go7eJzNvscysy9ETuuttZ9Mr7M2eiR3PfxXW3bNjhSmilQXQ9RrgDiGlIycU1JeiTuKc2Eo51do6
s7gJxc23yR+0Ku/Bt5VA9Cw5OTmnvP4hbFBJ44VIEFMclSRLhk7j1pKGGwfROnMICqgWiAZvH43A
FaT3w6E0+2ZNjlMR8t3vVa+cN9RrBQ2bKulZuFnYJ64ww5TyGWbgD5+mlw7DYjTASCZhxyxOhIth
m1r0qMrFVQQsc/1MhN6GMbxHD/GS+cBZBxINrQbEqicmIuPtAS+onXIYSuZAeYFFDp89ae6xBcf6
brXlQkIDKj2CVVqryw+wdXqZfBgVFDQM7PwGHR9yO5fbYl1tvNRYC4pnIM5H0bfvFfCsJ7QxEmBK
QWdYQ5IlbbmaUpov+SYg3X1guZxS3CvV8+oIzYRgMBgHG31VujrgK3+pUawRwuOTkcAe17bemva0
YlVyHkYB0w2sHTnqtsRTBgLgZGp3S2BNv897HPP7rcwVfBBl49zE1AbNMv0zJh6PjuCnp83yO147
5RVBWR3/yPaB+gmhnU8HgVwqMVD5v+B8cBaybdCTuCHuuHZ78XmmQiQMFR0JcUEIVHeeNU2ODynR
SJxhdbXDBdPwEi9QSo5iVmLgcCiPinNTUqxtfNJDr5w7FVD/8EqkP1xVffqLIDcQpaGWx1SbSkpP
nIkiHyy3h9kbUPuw/S8ISh0CEFZkiktqHMB+tTNV8ZNf7viillbmyT0t3Hw6sLL0AR7Cgx4SiuBL
OrkkACYvgsAKer25JohyCjKLjAWb3vivTibijnikJIQ6ABW1980n9T/oepkC7HxIWBP3PLOfqudn
iawYQTgBjqzfp/rHDboGuMdS9kY4UP/S34kndCD5k4Sx59NLy/opvkuw/+hOOQigF3ic+4VKsiE3
x6D3xvPyM22DV7Otz4WIqzaIxAzi87U7vShNH7CTc+vGK2SSU7nsfQJgndfHz31Oso5xeKNvviiW
NsGZsBYTjtpeACkZH/DGM3OCruAR8JQ/YzDhkuPwP7uIdUTy+0GEkvxxNXoI8Zd6XzG8gJIKY8Vo
KT//q/dp4D5turyeWesI3wHb/0/YPOCzxJx4X0yHxMb0PA2FNOlFKNuM+vHSVjTsFXiMnKIEdB47
xjuYL/ethISNG9u5NsKEwxPCkZaqj8EYmgkeGdwryHpRf0f1RHu8T5LjSu1QTjWVf7+Sqar2EQNV
F04MerdupYxCB38Rx16H8ED0xWIrzNdlnyS2qzu3zBCMMOun/Ud5Kg23+zQV3V3h0enq4wqDTJg6
Kpj6tAJPl7HyhZ05Q9ZaUXmMJWdhmkOgHgg1HQOxmkzGMQOQOouBvh/kfpJwEbO2VPyjd3Xys2VC
Flu22kWmbpCqZKXxLwvXBefBd81pKmKCUcwEE3nfi71Rn+kW6LvcrZK30hvZsVwHb3/MU3dieqDN
pXrx5IU6Q36iGz+geSv1nWY0qRVqazMsnL40xsCrqlN5FHUXgdd11vmGAp1+3p5h6HVUuGQF2b50
aX3BTgdi28k3s5NOPmnNYzR3w+qNin/NeLwI2fOxGHXnxMJ4jHxUjGFalNDbLvCPgHxdrCo3124l
2jjEsU3rzs/U7uLdOMA4np8sfDX6FqX8iOVmG+QX1EFCLuolBM2woaMRptJ25nacPuaVwncTKaW4
TV28YFoyadRubAwxPQ5cHdecsuAc+NXboEJNOQSJOjumetm8MJD27i8cT2Ke/0sdM+uqBxOl4KOm
BXGK6bb2H44F2p6KHDXvwkw9qF/uLGksR5I7c/uO7M76yqFG1FVe5EB82O29ewAc873J2f0jRPhn
sR/LDtEgQ6ueemiNg0FFM5d2eSQcletxhPW03gMzfFaOKZt9hUKP3+yMoDt6k1wcxEhisREVUld4
mTzgy8dNIY/QArEXM0KVWAAgWpUQEWRHCs295oN2aC4QBnWwkHvAMsQwnQUSFpSbqCHzmMB7HiRH
RGZSbQwd2P5o+xKye0fMuZDCnjJ3pSp56EdIIwK9/vChUW1RRgjQaDGnvp8wlcSG2aurRqeh+wNp
khPv9h1/mg35y7xEwjSu87eCeFtYJQSyQQSRMcWEHcbeyD4z0pU3EXH/W0tfC+Gm1uE1jkLniVv+
XImNq9wRgHYVPVYtrQLE0U0pH2SqHzaO5h4QwpE4nsJ+tMRJk6H68EykC5E6WxYDMq+DgXTbz9eD
i0zGBdHYoLWbCUq/xmYadymdcnatFOILJaswDY0HhUHgVd8FNw2gwhIho9HwZ1RyOX9IzQjc+GQ1
/ZMoSiy+oLlqju0At9u8MuPhDKuPy6YgnBGB1DQEFRJy4wdj4uh+JcxaRuONz+yGbwyXrk7fdaJR
GB9hIni3pkW2wyLxzdSl78Tpi+jr7Wmi8zJFy6HJ/ukqQupkCgEoT+Yss1bo+rlc0XxcCeoOfDA1
So+tbQKFWDO0oTZr9axlM6yLsZQp2Y4oaVBcAqIevdJ1eF02PQHI8bxxl+EE35stJV8qMpYC9Ylt
PPf+n48wRFvFgQ8alBRuZJmY94VV7gPjHvjFWeXJO+4fDnRAurp9lVDQvzB4G9+tsdWX2VGVR2+w
4in+qJ8Do4vQau2u+lTIXO28wY6LNNLB0Agcf1vvDItu7PxiKOqfyDJ8CNmRSaXWUlfGv3nrofWG
hK0061eaN+DONls27FnY6VGAwICALqHWl293+B+lqSA38KrhYRfeF9HDnLMJuXDtskvHo26BoUz7
4wrNQKDvEm/w2YFyFLguCgNePAl0/wCXh64haeV9iEF/3pmjLKNgLm7bgBYKv7zEdjEHDou+o+PL
9N0XsKkN9KDX2F/lJkvkUtc/P2UPVW1B3OY8SzbVJQsZso+n206CZt2lQam5VNPe7zVQJ4KB8DUj
l588oNoaKVnsJ04Nwj59tzThrmxsEcr5sLRDzSjeGIXEpOfqDJTMvigDCqL0cy7iY0Vf4j5tpR4x
QpJrUx8HHBROrERkoSg6XLQfDiy7MQKoqz3YpUu7bjXgu8Dqn/54LD1kVANJZXmewAxUWjOS7EyL
RnqqayRbNqvJaTV/h2aMyxGQEZDXJz6ESKWlrmoDfYST28kSzdjNoWXxcxrfVeInVQjQQcTGGDO1
p+dmnAsmtTapaWzovV4zBlIwDNEtiDncGHSKg3GDqHN43juNdF7EMQmrR/APULZveyo9PXcDr7hE
CFzeE7oCQdHQQFwKfZWxsGmPRRpzy3iO9uQ5EZO7oWdVy4o72FeiiuFIFQrtcV/kFQBPGlsm+ok8
p3HfY6fLGCg6+TjMgqPNjODGnMZSAwzNbcUCS6VBlbj3VcNj2HkJT8uZZoK9KRbgINL8aPB7sMCi
nwjXgD11q+m+b6G/ULmpBi2ilRgZChFpoYaBiyb46F54hxMdbSHGdIle48mu9zhfnjAi9ADEbBQK
0MvBYS2yliQA16V0GufYsxvha78WM5lDf5f69tixIFUj0PHJChhem3zFprhzRNbdaRb/LN5fvGHE
0ta+zW3MbR3ZerCLka07rWYJz8lM/3MdTnav+FDCNJ9IFRz9/2oTZkeOvo0vcyvI9JQb3t1llr8b
cXNaxzmk/I3XWiNE8nhuLpKjbDG25G5bXrhp/ay1xvsl4rquv3ldQ7rVoeEYEZBnAUsjrcTcZ2gJ
R0nv1SEZdL3k+LD5uJce2Zkz3sGk3QgNEIyRYHOoSJV/gY82ggZMlCvzX6MLxFRBzhLdVXORnVFl
HlxlJQNH6yynIzGKsQqsjPnAZIZT2iNUBZQga4vZBO3VNhI0jQxxckuUa3E1c8T6cf4cUWvF4jpf
vPvMPnmgs8GEgzunr7g8hQMy4rp3BKmNfgCPdE6aQVJAfUoo/kcFh8kNwfuh3ECG9wZ1jQwGJJxD
8vzUZoMueiy4hlwxgUzTFZfbYPnzwnaoWLdFp+YPyQPGe3TM7FUN9HLNH0WJBbIw1v617ToG3GLB
ZQ/FnOGzeml/o16no2U3Rg7E0tv133A5k/wfSNMf8KgQSA3aVlO5YuBUAUGcmR77wQDwoHIsjWgr
uZ9E0daEWfZJTVRZiMoElFHpXHvfii3GApMYMcZ+092dRjdrtcZ6ymsEwG4lTrGRyK1d2pFxpUxl
6HjpvoG3qDK0EkhyIeaushLUAdIhhWHF7kleEHsSbzvFeKO1sGs8A+zSkjAXswIVSVki2jwPV1Vw
obsNHqPSZL/5kMWqO5NAkF/l9I/FCIRZm0OWPcJRRvMZsVLZLdSMKBdbTp+XL70mKMFVZaLjdOjr
HGQ3K4BD8Pkx1y/V3iedRho7FQN+z3yTIBAaIm+hrAXiLp9FWgJdOLYHrI7OXjrl9eea10UThs9P
YoT7uTf+Qc2DB7KzDF1fC1lR9C6eEOIWV9XtNUiNccEuIaCZXnOp+TktaRphmV4UmsCYZpbeUIuf
4J8cn6D0Nu8mm3rEkwyw+5AHrJ/h1j8xDn1Ywpz5LXFCk03YTOssQXZKcdpzIqIjUHceIXDyK7xp
y8fmRHiYq8aUMEZ2vySxEkR8hogRSv9ZRrzheBTAoDrZ3+7Qa6v/Th0zajOeKfeJqnvFN7tlcKbk
lHsw49lE/jRBg7TvLfjnQS3q+0BEAy0c9bNzy0Zzi5/HMRmTqkCjd+3WYqoKb62Oee335isS0wsE
1uVvTOGQcsafVFNC8V1nokFkeMjFDKoUebFhKVNJaQssfIVXWCDl/hHg7NzcYZ1effLdbjjTH15y
tQHSoZt9EoozINbSnVBpTllrCuRWijTo3N+daYVR8UR2NicFEm3TnfwUi8lhtYwdwNi+2NveJ2/Z
vac5IheCTxW9kG4cRFzhimP4eoAaGVt+6V6Nnmf5gjaGCq2uoHN8TVXtysG1PXJhE48YH8ZS0eFC
JNKqwASKhgoMHitvKyEYBNqdXhZgYym6ezvJlY96OlTbc9bJv2aoW6vVnIuhtcyTQOxtErzViFWQ
Z43hZl++X9qSMlD/SuR7e3SrEHQ1u4yBKF65bDNrBmtskSFj9KKbbyJ5P/t2fST2AmjZAr1dQB+8
NkOBKcJJCzoF/fO8puFIEzAkL4bxSOkk3UUv1zFtj4NqldZmuwjrMwxQCpA4SdPZBycLOJM1taky
oo7djr09DPJW9FYBHQ5MOmdRfEgIqnr7SDk8j1FeKPsbqEceUKAM5lHZrtx0stoQZqevx3zRpPZH
GRlndIP5plQUkTuyAKVYwDqA1H8SHVE7buUjk+gj3TAGge9R/dljfDI9wzoX6TMoIMd7q3GliPyx
Vy5xcyBPZo1hQ1KvUVBVrJDY789XLAsJcg13Z/kY3Nz0WDDMrSRtr9VHo7WFCkxraZNH0z1R4H8p
rtU1Pwu/x16XyDB151pZkkfzXm/flrbp20TU0i847V54Bcr6GZhKq0vyMr3ckGs1TQNprlL2Dagi
p82p1Qzf1yMCcOotyrOBB+mtPsKz1VqKVFgkOCpSTeb83T5qz4zNVIJpK222uzAx+FoqWZ0pqPwM
SlFbTKG3rON85YYIXQA+F6NHB92HmXOd/d8n4DdSOignAXNJbpGBs8R3smqEp7OsdKibwIeJN5u+
5nVGwe9V9aIt2tD+wbuBUuOPsql6nb2n7H0D7JZYAuo8ZnNM5JySoALsWArRcPSB9TcVOdBlwpyk
St/wubgzvUMJFGQpcCmYYtVd47kRug30V9xOHTqunhW70hCF4TMt5DlyRNChFVm+QohZwLzH+IEu
rdW/eWFbroTYdNlooOfbzjxfP9nr45ZOh8aZ+UZlUbZrwbiyf+2U2DJbpPbKSJW59nrwkAOIase3
MUCrH5mYp/Ji7lntmaFIbVObfmYn1b9Bs3Vesh6xMQuDweQ/i3CCEmcO0irCR5d+X1XkXkBVVB3W
tffV675ViY0SlDhMwDDzGS8T6XV5mpOGVqle3kFiW3THeBDsjzKqT7R5YSOwrd08GM7KCDwdA6cN
UsJ8+V8lEZMK+TKa+BvSHtN57h7ThTr1qxvMKoOzZVrfgJgw5syxBOOBeqtX4ABPjvv9M69Vs8fW
DgD8AbaiB3XuHJdjPOrtQfKVRRlNEVJ0N0qfbQ4yq2PEX9s3qGMLWAfeKv/gOPPCY6iVKOkTVpCX
bu4+jlOHszmG0qEDW/H3d2pvB1lwLHKWlVcf45mkeKO6tjhnxYYXOeXZdn54/zhWMFAggt7kRQI7
RRioRq5HeFbA+vPDeZV90XGq9Tfk9KOIy5gQkZCg6DSRr96d8MVaQMwWSzVzgvQ07NbAlbYZozNJ
qpw292iywbpyLAcdwaytvlfWa9PlwDmNUFt0bQk/75QAXZ3FxcGGDFzNke/BNlY/bR9GMf/pjwRp
SD7HveM8fpbZI7KumUSF15QvF9982B+SVIhPdr4FQz/ibVW4/LY06P89rvTkrUPCZqWL/vTE6hIF
Zut6G02KCwE1JnCef02McV7CNBD5VvJrGP6diaBxH3Km76wbZOn+9s3nsDK6XVUCId7+iMe4JvkF
KokVFJs++YiEToJKxK3y53O0EqufhhXjAoRP6Gh0iDfXqtYUOmCwyjOwWrZJWyWuM7rZRriheb7+
qbDW9f97UXddpmyWzBrEChDBrbVvVcyTU/qjeCM8WIzM9HLtSn7390ktHZ4cYTzLT9N59cDHLtc3
e8hljTHWnOE4zz0XzXdm4LPDwoCWzsSlqzxhAsQZx6Z37fcZOen/T0isJ3DHVLDj+0BIs11gaB/u
6tN/HqHjWE1u5ZNPzCVVLQQT9ejH2EbrCiS4O/MRdu8sCUj8OMzg7Pylt089XBDNmMb34WZ1cgly
cmkoC650C7CGr/FgOnyHGuXjNJx/gdX1GF6NhveuwBEAPVVWTTrpMIFUfw+5gsYCJXIbs5qyAevu
J+lnbL4Yeg5ryP0alLqNvEtXVpYWleTc7opMTLGMWGVxsaSvr0Q7Ckwze8gCvdLccWJMTwHev4bd
PAD7jq17b2DwAclSISguJfWaZ4HKkSwUOrML77AaS4sMgEIhQWNKw8EAsaZbsu4nQbzUBUYtPORy
EwQZlvNP5K+poMDADcsQOO23o/chQBvBSuyWyOJAErxPlyYXl7JXrcnQnveL3xbHUoGecqIqkD5s
mWWcRly/SqiMfK4DByjQ20N3xv+DXCbNybx0RFUQF3yJ0QOriEtqXlkVjzDkYXk5q4SHf6n1d/Yp
w52AiMarFo/tmTvqqoOzlVOP4vmAsPjTy0PwXf9o0SXb6gVgk7cN0a+FKgU4/UgRm6bvbOjntGzF
QtdZldud+gXJcW24kzkk0zWkGqBCL3YMHAAUnRNqOnO4MArSLNJ62w6w6MLcWAR0OGHqq2IMiLI4
JrtWnkO+ooRSguzLvziPY6G742s5ge4YdPVPzu0+tR3SiGSkVK/LN1DOJk2gdHp7JKpnNy3nnPjR
viRmjP+lEAHpyTeuTjDS5bQD3ARg5mqPv+UHDMjtQnwVIORIz4+PFI3vGx4FGO+oxvLBm2merlle
s2LcHl8sbcf2RSru9MAnK6BqFYM6pRdepOldJoqTJPL8LYh2rh2Aa0rBfWLvSocb6NRRV/M7foie
ZL30xasChfEVhtbyH+0VdqCU2kTNC2QTJQlCjyr9DKbyNWG8zARb2wzu1u5w15kaAZENmj7SXQ4o
tIeKeptEDFaD20RjrZhjghF+4aJHQj2tb1IvIgHwidvqhUN/qscVW9nwH1B1qPdVscTGG583yqap
BPXf0TnlJVfRPXF4GCGqzgEBhEaV4nfm6Oz9mCN6T1nwwe/v8WaNFd3U+RpCpVE4QE4N/IKyFj5p
0Fpw7j1e6nTy00Lkb1D+PgGI8s/CNvgeIqxtymVFvXuLpZ0G1ihmtNh2VJXZ/poW7g4tsf82hwt8
GLaMssiZoq7BgegzhQOhtAUafhoPF17BYffTo+ef9XfmBXuhBwnGfG1YOnJqBtIAvNYEGse+qHrq
tQF0ynG/T3cWQOZ9McO50Sj6PoWW2ILKzJiTzIg76pWgPZgDRMgoGsJ2WQKRa1CyESEzvsdSwDyi
XWvrxOtmKh+Wtj12EopwmwxZWarVZ3lo9CV/HgxKjLFVw4YioqGaeEsYJ3tIj4rVlQk7/87dK2gI
H39Q78QrnjDLrNbuwzZR18xjc7DLD4iDmPkjIKUMWC12lnUilDas0XaDOIuFIrxSUVYfsWp1pEwl
Y0pPpnwz6zgBONm10bal8yiq/T0p99xpF+zoVECEZBoZ4nbXrxhu76M1aGv7oEigutK4MekuZ9TN
cX7WEQVpp7tOuCkDaFCzCwFZ1h4N9gnbHwL9SUO6roklHP6wMBIeyJ4D/7E+ej9L1Cvmo/Oi+ZS5
hv4JMsG3gwJPZHvjPIvwavLNcnR97mqi/4FWqsrzIf3R+UgNZImK5DGpbF839I+pkL2Sou3AGdop
Ixycbp7WdcDp+cA8+zNHsOsFxkamUhMUp0syf+XyCpBfUfsQVgNehbT3J2XUbbsWYii9Ze6Cl3f8
/OkDFaR77tsoNxfElfHduZLkdwNnRwUZRwswZUp8yDc1gGmuS/1MWB2YO2CEZ4IA1aouJfwXsliF
5bzVxLSYEVp6vj0V5bQSp0TzuisyteZfEpbb+PRruG6GT+bAOnnvQud6CD6mmwg8sjnQGGrGTea0
DU4jgk5bSQfLXp326uotHtY1w7nr5gabrTKoj8t+18/xWyNn7pN/MkNUutAfAsdVl+XOIeWknLd9
oeuGVg0hdg8/mefjEwKgORcURFz+32QW2CJHcinBX2r9EUePTof3OBi8tWoCoDLZATsIW1ZwXy0t
YWXktXtuO97ShVgM+8LJcktA8kwEensCuG9B3OZmTbZV0BIyGRVuDGYG8Ujqzn3aqBptov8oVR89
VQnCVstEHXgoWEazor31MT3/lvL75ctDzB3e3F3oEqgRePqm4UcTxt07rYCv3MIRFyKJYpcCwZLx
gV7IbX1hB75VO2W3cMcZXDN0V0hKoGZ2bo0Mu21n/VMHKZECJTMAPARezOP2OFhFvP+mcP0Id0xv
YzxNTUbLJiQfmCAx+EBeuKOWPLiK/WlHiWYoj1knpIzlm8YCtDfl7L1VRa1hnDMfGxtCeD0cu2Wv
pA3wbbXGBqfBwsr5onmnWDw0+0Jmq8F0On+zasHHQQ10IMavP9r8b9TSwGy2PqPuA9njkSNg3a3I
An2ONuKWRFgGuNPvz44/G+KtVwDsA5ruP0omnTe9w2xEozUKtzHUBf3AOVeIH7hGS24xWKk0xn6Q
Ie8loQevR21VTjkkEbLYl4nDgW/BggApzIzoE6HVMxQt+pLgWh3EjLOAnxHFhKsap7TEaXrnGSOK
9nzFyTBDd7KVf7zTdrDQ8BejUloPX2WyXo/IyEzwaqt5p66kB8gB24Qjw69MiBZLUUJPZQmMm0G0
Z5YTAruc63/eE1J4MLRcDWZR0O5V2MQuoZx7zppDb90rx4VCDqTousn2TQVqTWHgkFVKmb7fa55E
hSQKtQpHKGhrQSLwbQogqiIbLQIFIw9PNbh4qyvc0QwhIGVpHqPcIILoeuNYlF/gs41Kmn7eeUmY
5cDvM+6uloiEGIEHp+V6tMEyEu6S4KyCIfRZZSDMhVZLy8RBLBhNkZ2xUVkZTqOHSJWIJMA0VSLj
ao64RMq0EoajWJso3nKUB2qlC5XeePYvdQ91ZES24Y8mTFVLL9q/koA00ZiU0JHJ94hFl97hOsNN
OMZSJNKJC3MMDjKhR0qYowkw11ITpbmCpvdXjj1LGOpBBuEDtej50s4SjrGzVwa/kdUjCNG2lMCt
MyGWG2MDsAqed/xYhSM6AQa4fwjSNjZg+3N8losyRFdgUQoRljMWOUgmdSo3o7Z14Ksq+aaVp2G8
T0gJXWfwOtNiP74d9asW15rao1aLS6ag3EfJYVS/MaQD11Z8n7uNsDGtpp8qpWiq4Va4BK261Qgf
JmP3MJGw3422XcFRx7Trazx2NTyPtgb4T7EZW020Uxu7PCqC6kuhBT0O+L4lWRaU7tF7sDi5E/KL
h6COaxRd/OZVjS+3VonXVtEBThUXMLRZTyW+FqB+bshkQ3F4IGC/vkXMi6qYEKwKJ5PAEdqANR4t
N2j2OBbufp+mkybIs7OMTuYkoV99SOdeiolIkGW8s6GyxYEDNaQQtCL//rUTiaQZLTgA6rpBbeY4
ylqjBMLkJ3k6/y/JuOYkP6sb6A1X09vcndHCI9zfAWcfERkP2v3qCRIkDQ2eLxqD7XaV+uBaV2ON
mNJRJsiLXmI3R/Ql314cwnKKExwzJ3xmv1vGDNtLp4UfmS4Y5y0CMXzV6RhVmwp4OKPnJXkpvcN6
BhsUQ15pP+RCqMU2GVZTU/F7Zc/n4VBr8IKp23wYz2mLJI38KokI0egg7m9VBIJIWugr4OMhjdox
JCmGtCHziw1J6wK1VFk1uXFyWlD1fcG2TFA24IFfVgK1YzxKOh22mc+7znOTdqBEOMRN5bnDUoYD
n7BtIcVXwuYEq9peDQOuhbtLF1JUZi4VokZCYZ/glbwiH9AlNmmcUtk9wimJash7ZzKvoyY1f1ee
92K0ZU7+A7czU5OtNj/OhVMaGjISGncHBD2ApDnmgDrGtL8pC4OQAULYbp7wleajlde/QLlOsWiZ
MDjxD6ekSuBvNTVC5vXnqCKyrzJvdpSHb2IdkUUuzagbIw/qfdQidhafFSy8KmQ8kZvXrelUss+k
ungFJfXPxhRf/QhOlkPkPzY0uxjvNeEW56jtghGeqJK6KFZUKc6Gq6kEIYgAtMraN4/FnWuiUzWI
dLRoOrOW31TmP82QzIqhwS2UJvTCc1W2OB9Bv7oEXbqTPw5EYQHb2Pzl86nPgtW/zOogeaCEqMc3
1id2HPGDnO2hwPOVbIcnpwebUPYf4A+pstT3/1fSC2VAFASszeX/qPv5dGfYb5aP7gvFkBGtHm/H
bXtKKf21HRMuKWoCfpr+lPtVH7hq3+qzYAEgWkEcEooQDG6LrAQiraahzMOa1kE531lq0tkqdTvY
7+A1NdL6/c8eL94I+ZMSvi9vsjpoBLmWYlhshy6NJsiITi8Kp3T69Iq6ocoKw/ywa4nfOzS7ULAp
emi/1V9SinMztcEgJdsFbJx1eS6SvEBPPav9ZOTCbszVNjxTyJtJ5e/Z634qMoRs74AZaJu0Duom
db4FNGK5CkdEUe7Z9KPOiwYNKp2hDm2JRjQNUiF1QgjGiGFHbElQ7BkEnUbyac+wHfl90jt5hP+c
PPSO4PqKbBQpp1CKHrWhaGXnODZ0ZEDem86tlpNgIG2oHNYMkUYAjb+CL1xDbggnPCJ+RIMcBxhC
+vrhME4f3i2gJpHSSwgfNModYW4pn+LziSGe6nqaBj2qENYiSatU8w+SWG8gpgqMWwDdaOOxhBww
alS5Wactjr7gbIAoK9GkPOvBuItUS8sufc6TsRQM1GKptw5vO8rbNsoCefdMglsBIjvdYp0I/KbH
uohkhTAJy+34RpEo2+tjTnUrzwKo43gvelqYmmNZdo2seZT+UzRLkhl/244QfIYTfWaxzCVZR6Mq
+idfFaMEtCHTR+5vpMIQA7yz0Kif/ep3tjVd2r5bmj3p18c7qbv8zsKe+Iklk/OGQD8fQ7tzGCL/
BNjRCCRLUmMpV8YfT6aR+ZmK0W1hjBWxI3KX90dUC5FmPLRXqPuwqjL6N3TC5LS2Dkc0/sZ29Vrm
yeMan/BYZS4n1FPSbetoQtgA2cbeMlqXgFs3pQjBBs6bBrerTrJRgNNn6n2Kf0gQ8qGUularlT7c
eqrK/w1ls3fOfAqMiXB09sV7YRtrnMnPto639Bb0JWjXcpjSATb6CMZXrjR5WEKr+i5EHleC5hWs
oZQZ3f5oKziHLPet0ZkuTaNz4hFLX9dUWyOgRbaRkFFokxwbOswN3Ebv20lexqTxW6htVoBFfnsQ
JwVFrB2HPEQDZs+zuv+pP/QCTWIVHp0d1cenHYi5fwNTOSbiYWdcbQwdS+G1rjSU3FCXdQmmI5HT
C9IvVZD4gn8XQc5UmuLX7FS3+7RdEoQ+JsH2kFSpe5N0PGUdo58GuBbQEQkkbzsNO2Luh+Zc+rG6
8PAL8Ie4oYUWd0n2Q94mtJUIAkgmWpWjcvQDrWQ+ur/f0TNI+1U+w6idxiHcfD3uto1LZKlSvJvR
hyUx4lS5NwlfSU6Xer0B3JDwjsMBzB3YptFdgxUzJl6uUsNcvQU/WDlSlY/e5YNDuCH3xMuZZVr6
qNONbdPrZFtad3Mjb/GmNL5bnLkJTB51ldgso475RiJLIapYZ8R8Iaq5oJzie7fFMXX7ceC7EHQg
V8eD474RwdbN6X+mtXn9Z28ywxB1jClx99+EQHZu4KN5aEm51E7UhQm0CY6mwDqG8wYOdQwbxoRm
M4B2k/vtOyLcTUskR2Ech6YX+B9lx+5h4aDKn5bRATfuT4axmhRsOOz7BwIadRhrAEihlC/jlEX4
6x5m7mvyablAR+lhh1FNEoCvBvkycsYhg7SIZOqG5vRlebHN7csXS7qO5zpafQtH8X4C5h3gflcV
YkzdwpkjqHyU4Nl5TYTn7RmR3fOSdxC52SdFoEMvpAhugKjoJs7eO+6I+0wx7G9IVCt5xu1JOHcJ
3R4uUMDscPo+wfNaDOTNm/MWlpofTDIjB9fEUFF6jCASGibe1VjIe8AMaXqD7D/VfyOOH9fPhOL9
SXv4e8uo09GTno2utehU9Eg1N5G0APFLYONVooQNGVqSicE9ooSwWp0Xua8xuSDASBPUEvavo501
WoXubPmmtpOACLV0VCxgshx5HqyIvBHEI/WX6padEBbzeXSSq5Zy5K3gJWzSlzWC+8Ai67APLvfX
vORQ/iSKQ7zVEUKDgdEuvWOydw7YBKiTUHzD4Ywh4mDuE2heyJqGFh3Wt2Snp6VirazDSlY3Po6G
SdzMDFj9lmQjCmxcgOp4/LBHJbreNLIm80Y6ElfvctcU0dF3BRs30aOtUsWrQ0gGhuwem8hJr8ZO
Sc8oKH670wpATThNyqEHkM+a2RABU+SYAxfiwm/ebNBGN/GWvGrlK5DhgAF6Nf4DLkkrK6M9Mqc2
i3qaYREAWEnv5+F3vBEdBn3h4xsbLqq525nG6XDnDQHggIQLkeNCqNKK5k00Rl515k6IkWpMLCEI
w2u6JgztlhTqT4pjz4iNyIH7dN1IfuOSAqVMwJpx2X23wfswM8BeUGDf53hOwBqYkEPWAQY/k+k4
xT6+HddC4zciTXIZp2kRIzRZWsBb4fk2PU/Q660218c2FLYwfzITE/WiKqhzQLYSh3FXM+xjZ1Qq
wlT/63W/f5bl3rIRZm1+fCRR2p7ESVL+dfktzQwvaJjUh9nHyCna7JYN/NsLOKKzf+ylghfn1yPX
kZ0n6XE6V6MYEixY/BQjJ6foWwuvL1wFQMjJX2ExGLNSFaxUtKC5Jk8s9gJw6sKn0TzYXFmBOY/C
mRangALVr2DHjMdKldvRaR7znCRXWbhgDTX3RYtb4db/FOdUfgCl/xN5xu7N2IcsYRkgxL0qLem4
F92SqP0qhIJFhMdMP/3441vXCfVDAYwuvxr074tsJ8M6/K0yJSGKcta6K9OKA3+wYn7cD0CVoWfH
+j6AKutlvKxVe2TM8AEBkdwT2WtB24/LMcZ7za6E1dy9Ha7Eyplfvmcw8/zglYlREzRyrgOx9BU7
AsDcvgr60GdfE+pWZ7/PBEm1O9PyocmS28LGCPLh1ZqdFGS7ih/ArNfWpD72/2RQtTaWlh91skFM
n/vvwPjT0qjT5U0iGcGYWay6WhchucSP6FA2uXdeNwwRAJzaDXSKQLCwvA4ZRHxaPXRxmtaU3ddn
Mx9Uq4vxxm7d4kH0qUKxolknicVX0MYzTbzvyheYpJvQ7c/DC7ewrz7WLSiWHQfoqjuk5DibhXk1
TP0ZE5U5/wDddyTG1MrUN732r+0G4/Mg2rUnTsvRiccClCFdHpkfYAp1G/QcsQPR0gtjrXPFk/sD
SwbeS0h/JosqUwWNsMdW8XNm/7onEsFVZ388DIUOFnQZEMQqPcTxCv/A5HCHLn1rLrJ0+aCZmZ44
DQ9Fx/v1UNQ6inb8C1NgyE8PlBcG1X53ys2HIj4iLXxckSodgNNwDsF0Rsgq7QdOb1TO7KYZoz6l
6EpCQJeLQx9v4xrndp8pQXD7+ramcbJckpVzTV9ZFPTL/w7/Df054kiwQxCEPWLX5qsfwrEVTOuf
AghpM/+yvfCAtj9Eh9ma3KD4Hj6SaH+EfR0jghh9LwOf97dQctNYiH2QJKmnjsCadTZ/ooIHLQLl
JiyIKNcEz8sU0Ip9Nj20MnPxa4YOeogOGlbio4Q1tSJ8f8S6y5E6jArtOvMDKi1cI9ImDOQQkirW
EE2Z9uZTveVE+fZJTrCiFVQ1sUrVMikSn9Sk5R3sjM9jPdLBEKtSd7CUECWK7O/XuGbqKmI7TOCg
MFPvDJLDupNHwJYE7jUsu6VpddOtxOieETcat09xvsZqdNlw/+3blx0blJT1x3g6kVM8EB3SbNmG
nulU5XOM6cuclJJ8UxqmTJx0cr1rfQg8sHNdfsgzD9Mu8pFb60eO2YcF8ioC97FZZCvQnElMeT2+
LLBewHU8rtLxmQP4pFzhviJvpyFdFJ68K69iBxskyLqROfYx+yaCDLlw1oa5M3XqWRPsiHNvvFT8
ExeEPM+MCUX3n7boNHaalB03s3800uyIg5YrTeSz4Jz4Clb5zifTf3Q5gjapJyktYFFs8cJF2+oi
9e/mLJ7Vhp/qU79JE+tbe3GKRI5AFdlpCYiPwgDyAdbBQqJy8Xcv6IHioL6m4dV790keWJ39btuH
5VbHaHQWCIcIOZgqeSfUy575TZOZ7JlSZHRL7Ur6xqzox359Oya+bj5RuMIXnvEENeY2zPNG+6fg
dhX/iXt+0GXqXbTfKSz13TuK570Smp1TrfBmbLg1W6xLJUoY+CdU2MGVm0HIpLJdDNsr8yZtJdTy
OZ9hgz//Qte7pqySGkYnF0qUUcumYzhSAO12PeGEY/KXtqt40Alf2FmA9yeqXYaYZkUi6PVWbxNw
v+pq1yWq0apVO+JLPQW2IxKGuXPAXuIXgpfxPNCketyM4MYl7jkLqcj7WcEh06EdntBSKYBPANd+
CcIQwaGOULPtHk9Z+TpNrlfYe9HRcB94rmdb/KFD9VDAK3t95lmQ25ILn/1/bx272Cc5B9jgOx8r
4K+z4c2Z1SmPmjmIf/JTd97UqryEWCZI4nCgWQXxvVj3Uy1XY+94Hb9o4QuCnsJyg6oL5oYnCG2+
Y+WCDMLw24es/97GZrcM2LfnHlvPhD8Yac22sW4lNVw6LUqpeUf8qYfCw2FtwNJFoQUqY5TeKi+L
dVc0pbhhex9K7PLxuopjsSY0H7gCctqgOwckkijdbfGSiEMAY1u09sskfx8T/3peSk+TNWyD4IL9
CX6M94zDjyLGMCnU4bWiZ6C/DRZgCRXKfASt0S11YD8WkW5x905C4CMaH3fZO87jpOViXcaxrm0O
Vb4TURa2hLBnjjkVuw8o65OF8aUv2x3fFCBRFdY8OWJCRtdQ/FP0Hvx0vZ9IbX5wWlT4gwkN8x8s
a0hqUyupknyWsKztf7aMMW7AS1azl0eEwoQ8O7d/XYYcPsd+R8N4FtkhkYNemuPiCs510YQU/CBj
1m+K3Wi8M/Jr4zFj06ep6vM+Q0Ccefwef6jRlsO461xCi5PjjYWMM4FBHc3PPj0BtdJbeOVaRiPA
cnmoNWWlT3FsUYkn4ukkI2Ss7IWWmqeqz/jbEvMNWEx+ybpP3K6wtzVMOm2ljm+2f0Yesrn+kdog
QXTJ1GqM+KjVu5v3rrtb3Fb87X/v+WDh+VptcTFBurpUBicj+WMBZophYvx5gUfkZFzNkOXrc0wl
7S/pZpj5tYkAvBzhryCLW+j8spwlGY2QKNxU/+iScMKqUXKVX2VboOotp+djvVPFoY0S6cAmDSRs
xiFxaEjpumAjsfKj9MZrOc0MKSisEm1va/YSSO0ORnpWr86gEfjPdS3Nu5+72S64hehF7xVgp8fX
Alnm8xGOtPBcUz9mzM4XYxovRkbZgFQrfnU9WREwx5FtORulxucKV4jezHGAsg7fw6+tdk6tG6Nv
hJkyxZSuMvoiee8rf1IBVRP5JKK2E2buli3v6EKOYUXR463diqOCffD2HJHg2WFfPgTyor+5yVru
NrzY+fUdAsGl8/X/cnPL+gQQI4Z3b4O3jn5QL0fExkRhiKTnU8KD9nTD3KojBSnRCZvgMvTQgthO
+WaWEE3pXt53hnlgUmCPzKOKL3ganUloHlElZmw1LvbbpJGHmS09QE12dsYPNxHUKO2tFkYV0otL
uDaBZ7ECGhG/09H8diYRkPxBoDIly4guXGJ8yXoeP6LAWDryrVSZSz03vQeNmsua8Io0Ysu1NHC/
jf5ZZ1Z5d36d9zngqY8T74OzG13ANVHcJaWxH97OCR19ALbCESoGkBdWglxdiJW3ltMa+1WhxamI
tFhXV7uNhlC05GSQ0Bi+biS7iRZgcHG6Zo0j085QhdxKmmjIJ6gU18P8KkMv8iVewbfbij+CKDgY
wz7YurBikP7Qrrx/k+OPreDAbWiIivU0AvazDaZlW8guLDYCpXOM4G0yJDHCzHW+iXVdg9AbA8rH
O48dleItVQP8zJYBar0dMpeuXuxBcERHL5E/Yechjp1VlvXMgM/7qCYZZsP7kcbgAZ16Op8Wdek6
WhpvFSGDjJqpHsUtpI7IuRP9mObtGRV1sM3q9X/nFQ3qd+aeyWBF8OaLbH5s0i7SsSkjNrG+t0J+
D+n8E00HsObZb1P2pJ0IuMEixcLS8VD4sq+b+k1yQCtudT7eWHn4c/WLdCGjWUB9DRq42lsdoC2c
yRoM64e0EtLUpCZh/AajI5ICnCVVGFgrwL5MXC5Gh/dp99vwMFvLjypc5X1Swe6oCyVhInQ+tSUF
Rj+bkc5Mfg/eMz3fRkLbYYM64MRWZjf7ZnH+bAXYTGe6LuMdwgVAV2pJzlKFMWwBijLamPu55njS
aE8YQI5hwEvxWs+tvPv9Xkv1XeeFv8buk7Sk9QteDh3Mf6WN2DlkEns82uRGDhs1MTzyrF+GvBQa
IMbSL4pGRhtZQXzRrWNghyDyD9t6CeOwUvh3Rb9Z1jM7iueJocjJwBXCGsgwcL6rZOy0OwXa3nhI
fUqWw21Fy4fR94MsyKUoa5PRQSZIQQMKEpYSx0qev+gnyPLJeJkVD+HwVS9Gs1alaO3svozrOTpY
BXizzM81VgEYX3c2bOlWSGxtn0qRKSKnJrIMs0C1IUdS0riFnu9myemhtyMVfy0cj6Q7sD4EP7Lf
r0oEpmlwzOfpwXtPbr16TnZ2A1F/XRXXO3YKbu4GdovbbpNBbcnJ82AkKQZq1mgjKt2Iz2XKYgQY
oCpzGZEXtHaX2t2a2eRWLLxeFts8uOSlqH5TEnamiUaKxczsTcYocee3Ia2Koe7TyI/mf98A1C7R
jPdM7RK9vFMOLLzJvMiObQuWvENABcYgDNZzc0ePYoKtJn/Fol8QznG9q/KrMDqj0Yk+iuMfEqrj
aN+NneILZPFDJ2f5NxtEJneg5bhgOn64CQXNDio9DYZh8UlPvfXJV0+HDAhQ1v13v9s8z7wR/fJx
KTHkF9lv60wG+kanAcAESTZPtrdEptvClhKUfQHlwOHekWn4uGn6yZrTJhDhYM12c8PTUNFIj/+p
N1PTzamHqY8VP+Hc1e2g7eEi9JIoOTEmQWJwGwVLWOiOeSsgmX0WKTzogJrqLqa4OQ59RAPBQzxq
VFCxBA6LdPEUPmynX6OBpQNfuOYmrj4eNEoPYPQJLH2W8L+EiGmTRL7tJBBvrlYhJ40fFp0pw+86
hHML26P/Oum0/NXEiN3J4Di0aJR3UGV3CyOVNEDqOor0P39uVA2yHsVZOTftf54wvlllj/y9XsNQ
/gmggwTRzFC16BYg+4zdbq5QTSpt0rrXIpDwlUR2EAdQ6xgpuNBHTsCvFEn9A9npsmZdmB05RnLH
6OoyzTs1+AwfxHPaDkyUavyM2FLwAGdZ8/H0pLI5obPOHmr0w07YHL8UfRumum3IkE1Q/27C7Ovk
qIVS6vPKn/cdL/Ve8Q6NssxX8rH2QBZTaSrMNdMzaXl7KJsnIV+08zcxJLUNF8IUV6SjK62OO+dK
nPP4ytRMwGxjfQZtfAx0RwvxQyzNlsEiS6rDRpPERrZkX8FWaCPFA3bsg3R2f8cbTrrRfzekEMJw
tZP5EyBpXezornHGsZ0V+Y/YbGE7k4AA6uxRJl5EfSTl5Xz4tHNnG+a/42KKJS1NZyy72rv6p+/R
5omgca2ADEDdLmwWeDFX2POJY8rbOBRxuiG6EfFBxHLzoaDpkKv/ySdc34FL6jA6kuc8WOIVO/KY
ZzNvtzXd40ncVgX+Gmi9zNVFKqq0KFjUx5DKmM/QNskUBLXZtu23ujM3LDTsLlrvUdGmBH7EUtfU
Wg2xzpCEw0coWdUjYSGqBi8xif9+13ftvp9xtCBJEleSajsRXQA5NIw8YVZ5kg8FNO0bH/l4NHcQ
eZ6fyxOcPZzixFSKop9NYtR3rOVfm07d1V4OQdBqagda1jyTQjJEeXqdl6gwnVY9yFZDaeUDIsPx
2GIi+/SnYq3RXa0ZQvU15Qx+V52VIbRj5byy2Tc1gDCf7pQI9MPewqrUj5W+qVangLdjjdlv/PV2
lms1lp6CcFXSHpT0UHHa0Tn+rGdyK2/cWAzw0MLoQwMYK7Ah4sPOfm5G2HzjVTS2E0RJjxu8dmOk
/VS5v4ImHA22yYqFWfda26NilNP6dAhXFHd6bJ5PY0RT3JTzWw9yhy3c4UUthx+LW2Bb61RokV4+
RaGZvHR3Dxv3QuaTa6hD17QmPU+fQieykiQbCfogrruaZFk1p276X+9/caPOzstYcPQtTMIBbCcB
rFjNHh4EDLWl0cM1cxS1bLbRfUyiWFL3PW1YZaY8bJtUXMZumoEFKGssNu1vf1jAIJwwPWjuAOCC
9xXjvzpN9BQDPWlWVfnweB2CvQ31zbV1A3892jTOl63RLOa19P/Uh2ZKGXN8JRaCz7QuEqbT3S3R
eN8ToRV1gvo7HuKIUpzSssPAvW4ECdOEhUHtnpmex1T3FyNXUpE2bV5IjLRCRaZkTztgRe7QXEO8
O8fS6y8g+LAQXms9zDhCVlpO6Nk3rFb73qOSL6fvJfnykabHPgblgdwJ/kqU/N6K8wRxQAVxsbfb
aCFRyTdm/TszwOUDM4uKoexaVLFdievV83hkQQp9TcZutwoB66LV87YSsno59R2fC1ga8r1lZu6N
w3M6ohQGSLAktTuzmQOzqWFIWxzwBz37+qzzS+wI/gq3HfSEmBedh4o2I2v4rmyByhEMK/FskMj/
WObngpBB+J8woG3W3KcSPI9lusFqyORw1vg2xGQw2PZkramIICQ/JvTd5nD68mSK+tp9aCzbKcA3
0Bjs1NTWC33s0IY5AkZxEYdwFPEpFTHld5Z5K+fpexhDyUt2ftacuxe/KmZ1MMbcsKDoUz+wbNXV
V33f44aLXJR6dVwXVQZ8UtZYq6opIPDXdPUNY0J19wHFARql1+r6eGOs5C0CgHVs2LKkbPTShVwl
H4DHOQA41INgiH/WAbaBsYQBHUWzoc6D1H7mc5tZgrKcWk24VtWufPN/Hheec9BmAKXsq2EleuVI
o2uynjteds9pG9WjS4+PNHPI9yh/0MfcaDedFBDymZHaKPZycWGagolMhO6XKtiW2Skki7Gdxnq8
2SDNoT9xzmRdVF1UcztaME5iK7gShIAg2V7IaEi7UDQ+w8e1jTIn125Atbbz6pWxwwU4z6uz/tow
jA6/27Q1Mhpe6Np0MaE0MSFQpXKtl7miBU3EUTHv+QZ98LBG0Tbc/BcJsGUiVwBTAkBAYGP23N7k
2Z8oyKb0cDwrUZXw/ngdhn4s6sxend6AWlQZAIXitmtw6FPCX5bCgTJ7uP8hB8Vrbw2n7IlzUfoe
w26v7v20HrOD4jTTIW8Wt71t0OMhnZ7sNwezICNlpTcA+dzCGsl9o+kDHgP2zYXn9LxEy/U87SCo
mnnWztEwZepXPzqGvrwWKniel9hA9g+hfdXk5EjHlf4aCOgiX8VfSRMCyJHvbxqHtKbqBcJIyZY7
fgXbBSpj7jEUseiQXmgx+vLDALCYSgWYzvAfF7B7/ktu4VRrEGqC6ECGqhgnFIRDKCgfrIRfSzwJ
61AcGPF/aFe5eOl8jTlkQTwNXWSydOjpb3Gf6bZFoWjdyQASJxSAaZzlhJGegKjT6HfMEtpIs2i9
w2zsg9t6dSwpyejnsBGN9AVUnDguajunWPlBeEkuW49CFadPms68WH95LLGDMeQtg4AfKgpE9k2Z
+YwAAILCNVrqhD0Kl/3NHdXF9qA+O5Z6r1dtoUvULXKmXQPXkKdh6V4imkd5JZgYyrUCLRZwtaOm
jak2BWdwaQCFjwzUgUHiqm5+Kikmpnall1H4x2xy0Hp8WL5zEc+iVSf17WAjPq8AzQ1naTvrvEOe
gcYqxjBkcYhqEk7P+BoUG8mUh54UNIPKnjpiEuK08mLgv0XCfiY3aTV/VT0uDAWCQrtUAQWcsGOB
3OtcnCWbBIdcgKftmlhcvAyXQeqddiNhOI+DE941KUB6K03LgZJQOInPji0StU5zhlGYJJtFI+bV
RvgysbKOXtgPViMJB7ou3joj28Ea/OAsnHkkM5Ni1pxpmZa2EwReIURhuCTkawNhCugzXXOWe3fu
F2eSXGVgjoavGHWkf/tugk8Fie+EN3siHgnwVso+V8WbL2nOOp17VBTsDEHL6YebRszs9PP+KrQt
ObLziWgTHVglOL21dqTAAeDTuf1ZwF1k2ojoiNlHGzKUfuwlu1j9vQVULL8Vy2WV3K0iEU7Po9nk
SnmH9POSdtz9NlBweBa/EbcR4W+8E+VYXBb4Gm0RN125JHlWZx6YqwKanHwuEiY8y27zvC7UTCor
sjae2cuLXvEqC9zNdKnKJI6FXW7dVA/v5KLxxXKyt5adX93fins4cS9sl8jbt5nBFG+3cN9MYSx8
qhsuCJh/tyR/p7bMlA4qbvew7/qmSpP+q/uyvY+GhqYEusb0HRBL1Ilw8OzrHWGsDhyT1wpxyE/+
ZkQVCghqAJwhYnvq3M+ieGuBFatZcybX6HCHAAeEZhje1LnNSwJkcgBy5IBvMFMQzJqKueyjapsK
qYa48NGszAmWvDat9HyzJ+RzXVpBw615fSib66G8HdqLU742sL33OG1B64PBR+cmQWUK7FH6tE04
07WiRH8SmThVtNPuc+hWGm/yWVlhuimT1RrDmBkPYOj4GPWQCzsET1vVsKG/AixxWy7w0/3QUkj5
hcIcFKHAOzZdpXOewwTYcar+lcv1va6ukSQv5wwUb52HXjbnTxWI3MLmRJf3PQHViCGeqrv7/MM5
Cie56oD2Na0Uf+0NgXgzXb0VIrJ2IHfwjViKcflQqtrG+4jiUU0AGE2NwGINPnHTn3h3bjy/udbu
g8RBU7r9V3hfQK1TwtcXQcVQbuCjiMIPvXm5d4kdFUQrsQwLt84M+e/Xlx8lZAQ9EbC/fjO5xLNo
hwXfZmYdU0TLr0lHrGJ4m562CcbgJBnF4LIQCDVH9QyZJ7MY4NpSyAna6/wxqMM7/bfXaZufkpuI
fMlgJAkqX6vFjZgxAHbYV9kjEh8VxiAId7vZyI9/hh/B54DWrxkONagNYfjD4mN+/zV0Gi+hRJxM
8eErz5S/9enEeDqejVXNmXa69edflZWZ/lJw6WXl3PwmBuBmYL4s/gNRZNyrWIYLWRSts+YOZBi+
sH6pxySA5n/yI9+Ha30Na1m4FVX172es+q1p0i8xnm1A8Eis7s3Tk8nXN5vUz9TkZ/SX2tudHked
Go9QwtqVQFVnQxk+SL6RMKYw0sz0BcdJzLllz+Fd7f2Onl00L3gfGb9aYgLVNgAh/IQm9QTj6Wep
egoy0KFDC0IDgt5usb0OGcpG30u7D4RS8SeUKTDQynWzl9nPzqQItERKMN5MqYyxpTvrMwV3xDaw
FPT/a7ZNyoYL2HSdRQt754/wJCTo4TrtHhZJHOjdiTsqLykHJ+PD7cAUGJ1uQakUWTKwtmKUNFnu
mcLM/U0PftCSSfHqHrI/aqLzBi4t+9mv09YAL1FOjydXWfI23dfY7zLCpW3RxOUxaX3SgudngiBV
KuJfBRRqZm2vttWNbKIZEol9k/bRImD6tp37ZGmezu40r30lVBROkVuhCttXtbmWnRRBnMMYpSqw
az+3tl+MCyppihdHy/LhNn94UBRRMNcZYTxGcxEQT98a0thdCnbLL95Lsue+uyJd/RcDC0Y606Tf
KdkD/LGvSLkfdicSPJzndMMTvWlcJdRZt6UPIopH4caih6wVTh9GuggYHU8SyJkMQ7lKsyDvTRLU
Y5cGs0eI5Z01vsPSrb+hfPj7mEHzpq6oH0qS054UmVgMyWoeBlpKTgP/EKbrjj9a9Ryt17TTIE0q
L71Z88ayVlftxd+88rFE5nCbJkWKY/qScw+jj8uvDTuWMcu/Ob1/8U+x1OdSbzU6Cpl+W+PAOCDd
TBP4wd1lXv0touMk7O3glRz4Vo9Qc2IpbjsuDPb/MknDYpwRcYp68ieRBx/tUXNTdbQ3gsoZdmCd
hVy9jK0xQFcZbxZzLgP19MNXGRFu0k8VuF/eVjxR0WRR6rCcZl1jIckxrXye9MsaKzO6WKzLIBh8
BH3vYwqjmNvjfJjUKrP9R5MSn1PZGek607ksai4KONVSJXmKbzzPnO+xTdIEFNFYbpFVGIw5n0KJ
iQh6eNhlfmNDoM762M+Iwr9XGswBNMd4b0xYSAGiLubB2J8fBI4ck+jQ/45v1CMfjm1xLYVLFKj6
LDqJME7uADBhNibj3dy0nS0ZxSlNHok0TsMfM8RlntJwYmxDru2WjqOTkkxy+PfEBRGe6lk6lDb3
rGM1KIeo5ZMgzsgEE4p0iB4trBUoRhT6re4Z4N8F28Bn0HrmQpaZG41a86F/CcMlc7NwDV1Opn73
B4jomv2F+S+nWSQPsOHyAyTNkybqlT1/JSZCd2MeBbVJxs+oYKVKxkmMXW6WVA0rZZO/aqzLmvVD
7RiOZgfAd2hQk9j6rZfwIirOvjkFR98xHNtYXvjKAVHIwKvXXngD7DF3gv5R3mgJjssYmMOT7/1j
vfxP3wYqUbXIY75XZlsVTjgQzJIkez67C2mseJH1pQg2gUMy3fvO/yN9LzxqKXPddkYjBqKy7BHP
UMCdyatmnx2loSWVWKVtkQ7ChjE9T0r9fMTZt1tYLEU9ftZlJ2D67SQqNw5fcTkNnNTmdu+tGjBG
yQWOBA2IDptUcjnAgKkFoSRUQrxkw56n4U6Vg+cPTPIwkjN4zWPbskz4GYanyo4AeFg1CY2Tg1DJ
9CwYmL9FzS2htx3F8bm5JTlHIegbd9IVNCI0o0l7fO3BppNok9Ebq01mVxqBuohLDF+/dodhhRDV
brHhWvDIA/lc+1tX/K3pSlEwiT6dObL6I4P7hTcNbh/JE4evFJMc2/UB5dwnghtUu6t6XlGJuw0U
xS5xG5xOg0gyz4vVbVX4XJkjzNCQBMxmCfWMbmxP120xTRJtlei86aphqTRZSEMP80nhjb4IUl9y
HSJdIbCVCQbgTf3bYGsiW2AE6X8PPcDagECtMRZnF4gM+rfxyTd4JYbhgvT1p+DghPkSqASkBszG
YHy4LloyXW/3BU80xwiuuS6M0wr5l67QRDI6NthzxqBUc7csSkLM9f4vtJ8Kws3zfijzJrerGguz
DmOiT7E3pP8CjgG6b5P3bLU22r9tVEM/mQsAmK1hm6dbCKZnGZwTF25ZAqVhTUGdxk1KEbRF/Y2L
CP3VYC2f2OK92Ha0jRy53jnh4qEC0Bl04ISKIIYRAxe5mHynN+H0/VWEgTLPPuToD4XTr6fE5iGy
uq31QqKHHBeJVLu8FncsaTsj06yPoCjIm+PL1/8f5nSypnXhtrxysGvdklYBWHmSZjO4jZ0IciLv
XlUqW7Irkch8Adbaf3Zvwv0UUwIo07EHmbQ3JPAx7+y4xBEa08P3JGYU2G3xduHHLMgiA4/p3mEz
btBHST0GSkWeaDKHkOXUxtR2fXEtmXJbmp1H8wD+K5qMvrysOQ5zJ2RSpR4Cd3DFa6gDkaCNDLtp
6/KPbS+fx+SjNDgY8G4cepwNQGrn5C6xqryZRpp8kcfFUCbV/ZDBsWwK/ozuxB2yTePJBo9QP+y5
eTkPE3HSQ4z28YPyues7lhAcLcWkqcTHwx4E7FpgQoXZO239YIAaBlxH6Y6U+FM6dGklVrbz85ik
hYYPnNrD0fz9ehS1DV6R1EcVWJJ9ITF2RdY+YE9Xavsixrz7bs5/DFSBjITjFCRuBrmt3GW/GINy
Y0aED47nmSo9EmugRmdHIdPyAWLVrLumZwzpuBkxR5/goRajETLXwxUuxvUo4M5InM1CxVYrbIeu
XVLCarGSUxd/Zj3thhdefXqdHAogtQ80MHg9uPB19xvBO2zxluYy6clhxpEMjVRUSxjsW8uT9nYf
kFfnVeIk5DJylWDilIYJRgC7+eldThg46RooNJEUn71Gg1rQvgblW4O9JII/Z3IBYuGF2bRq3aJD
4dDnV2GiJu2c6a6FSEgAj0CtIZMv7CjFey1Cnbi+5tdk3DdgB1VlpUTlgZa6pP7RWTyxlv1zkzaD
dJm/0fkQpfV5oOmIz26Y/TufaYGZa0wAJxicjYavtL8rd4yDlu1xq6jfGv4C0mlsv48MExOMzR9O
ogp0C19BQ9W7S8rW6Wt4ze7jp/iEbCzuS4iYOlxAzziDcJ4Av4Yw1EBdeuS6WMNzA/NVZMUsiUCx
7OqZVj0ZzZSxsBM/qB64mQP1YqfQkdGlL5Hb/Fn0+HVhODI2lBMgEeg05SzxjFkp1rcd3CfXAlak
fOcv/eZXW7CgOAhCJw5KBY5aoRG63wgaxBniF0ymKKlANJageOLwX6bogl6zZZyAWu/K4AXrCObH
gtUDWs2/94bxbYazhOjVMN7dTxATIUzlVGemvTTqHaDOsdERBk3PFAHnzueaVUJdRAzZmbJYsYUc
4veFApsWeS+JgLRV5W5R4VlsStZDrTenBABFIB70ET5jOOsSqgzmewjt1McuMF26vjewV8P8KUU7
WeBU9IOsfHXPiSY+7vCSKFE7rvFiGA/N2Eemsu6CaRBdRiMLSHG64oNPY2TJODTkycNq8/57w8SF
ws87IbqrCeALcmz9m7rvKjgHO9hdP3yusiHDbaHGQT06GmKJACEcaMd8faC0nbKNfpMjNv6TWZYh
R0PCdZLsGfsL2nT8OA3hIWW5yiiyQeASTg01KMGJADCieQ6mmwIj6WFoHgHEyOcEBQ3e3g/ceVkm
WXnGuKaHWC3nAFMgVMoBWvsONurRJnZjV5LXYBrttZNh1hfkTrArA9xuKiD9IKv8BROH80K0TV+P
hKFtdt0UP4NnoteO1WybBFSd1w7SxQSMrjGKFeTheovujT/We/q8bB6XcgqtyLAVWBfygwZcUdPp
/948nahqk1+35VHGRXIpIE2rcrSD+6SSpUJrjyyEntwhZkZajPjP57WMQErHDceXMGIjEO8VwERq
pBYSh5UPOUyB0SLLXx3AsPUrxMNNNoBAVtQbnVlV8yAMnuG487vHu1Qqq6FN9zT3URF/UJRuWxpD
66s9zCYBWdQZlNnT6CBBYALoCzXs8XUN3kUweV00HjBjNoEE/nmutrTNS36j0rfrNg1+to5CukJv
qzjcF4IrnEtRWRKvvyTyzqj7e5+N54m6CKvQnUB3bUJI2lNnVpXxX4vSimibJCHX0EvT7MkdDe1X
GzOZn5OffXbj8P/ORjdTcLH08ymoKkUlGaH9xcdijOObHr6PmpNRECL64FJ/SxR/8LKPcb0mlIVA
zRmwQ9CRwQhUHyLSA1+CA5QrG6sJ178FEKVxSH/j/JrJaAE2ZwavVIZ1sX3YHg4B8aGTKCa/zcDg
oRXESlVxJuxq05K9kzouI5vNs/yk8eOiugmP+u4LmX5fAQ9GUF8LmYA22LSR7KbXvLFYHfCdv/qU
kxy9nlDKiyaZfi5vMq3hQmZWIUDkYlCzZfDFbHlLYhkh1JHsezAfuLAJNKxmZkk1dMv8szOv4T90
IGKgmJXncoKHQoPUCNNt+4qnPVT4Pj079++Binf2Iu0rw5P/5GtRj8gas4vQutEbNQAwWETzJ7yt
l9n1HWuRnchjikkLAB0NVtWOu3MnoABRd2BVYzQ/Z/6t6ChVMKpJhkldJWXCeomQ9+bebLpmZoMM
lrjcY6ZDRY545AyjGhz9uOSR3w1xlKw2sajK8gmIPJ2c4P152oxGwRH1x7O+608+K8A5FpUdcTMY
tOU+Iahca4z+v9oAvBANwUD7hBdUfHDMLvU4kRvp5djXOeUYEYzJIywvykfaVPPgHDzgUBKGU/g5
9TfzggAxO7wIWkTeHjqC46jIt8BBZyyYjjIbjs3+76ZO4WMyv73QNr++F4BSwSe5wGhQOWFOnAn/
4t3D+Degz2p+6DJqM0Bz5eWPjzfeUMbKGcMz0W05wpnRdVykqvLOh9lasCc+jNkv5PyN4FrBlf8V
ulhBynVEuZDIHfV7Uni4Zj5qEAycww5k4tHO/H3omnE5rFa2ZPujqpOzi+CjEbZHndDJsS5UIJYQ
1R9ZPUvbNhTc8oOllujTg/+sK1Gwt6dohjoCmUtEI8Q8/urU5FZi6rEJEvUPIBMqaXHqJWLsDCmV
CkC1/gsq3VCbPUrgLcspT7VTiEBWwC9/b+/rJZznTtlXy8Q4F3SM4of6sS9Dh/g9zJGQ0cW4Axoz
pB2mDmhiosw2RrCgOKQ793CyYHEd+IHG58UbNWEOEx/Ek1bqRpPKT6V6Tmiovd9ti3MBvdlzM0N8
poPrSkuP3sBC39zkqqmm0l//A6WxVwQx7vQ9lr6u+ryMBBHWi+ExO/xixSiPWZPAiy9Xpp6UlU/F
yOrFFXYy6he4Usb/PsqMK19wzNLutAE/9UGDuIAcbPcXGHbo8XQJ3F+2U8hcKgvoI0bntqjj+M77
AEX3xnIhV/V9gnH7W77aB/Gu+i6ukBlpvsjQBO5ymENzUwiRtcaKR79YeRdAwug7c+wrnIMYdq/D
uqYaffntPVG76hmpt8y4OE7Uwhek2r2RBgTRbL/TzcD+8w9xr/BKPE5KhmjbzDuyqz8mGsUJuPbk
tKLX26nZwkGjyVlynr38l9p1QhmVTfhEDayjkaq4ofEYpVwM7+YzBApe+mrmdnBNR37lLRMZ0c8I
lFXX+axtSL5gOZieDtQqlzK+cibUYP+2iRHrclbF5iK6f2DMN8Rq3f3RNwklDBLftTcQNpNV+X/a
twlBzEmE3UsMD/pVEpzEyc4vg7jq12Iyf/O9o5aPMCRdE4XDH6X+HHBxCWKvs4WVEmWO8K7OCVKB
CfKBSVOkDuku5W6iJEiuOF/yzXLtVRqmLrBsndtGc0DnOx6GLnqUI8oRjyFjyoBjk7ZHG26+gLne
RIGYfI4cexj01urqloduohB9eRTnrMDKVnIP7nQGebgzjqa+IsHW64nAPBJIAKFiHqnhETmxYC6N
HmCAF1KFIQN+qI08B3Ty1Z1Pj3uPQMOSZ2HvZLeoPRI5jIoe4WOLN70i9Hrc7fcVLPUWEm1i55RL
/XJijBmPvxZQCBvUr784pI4mW172wT1JKqMUE4qOWLQeRbDO+2UDoN7L3kFRwCWSbaqpYy/OhmqN
G7/3wYpxneMhv6OjtLXSPOhObchBQIg3xK0TVJNkqzeHNfkBF6kugX7Kt28bxzz1xeNKr6uPG+1W
KK/H6Z28BgFagG9gSgHFCZE+EaRIpqpf4tU+wWMtkQqbSGRY5xUm2ZTkMFsgTCygmi11CJvCHUmv
Y0wDpUOaQ38YT/vme3Kw8zcqs1yChF7ds3Y66oLu91/YVm6L3WfN8keimYUGRp+jop5ki5Vdfgm2
y8pZ8bqOeqyiGMc+cicP3+x1KX6EeXL65rfxc2umxBPsiTzZ5DAcB5n/k8dkwZU5xUjfOTc7syuF
IQKhc2I/+yNldV9P4gkBKmA7BL2UzkciFmBfb0p8Q66hGchy5sKgirwRdNdHAHSF4b7eGKhwvZsV
av2fssRwuh8NFzeiaF6yF9JT8vWID7UaGWkEmtJoXMbICAGd5LEqQ3ZMllvGGcdQmgcMZ8+EJb/K
JbDfzQifw92la5jdsi/fOo81glNNCNZ4pfz+0NO6iyE/u27RrOUDoeeAE7dWZEo3/1/A80qIICpV
twkjhIffkIbosGuYzKN+e+ScR8nOqrOn4W9eKcLWr/qz6klOeNzvj//gApzeSoZU+qDPHhI4TTWS
8Nt6wxMElArDQi5vpRwYpz8nBPFE1tLfK3ueIUoKDJtKt/zycKK3Y61Q6xH8e9QEkFVRaytSpXM/
i3LIk5c29i+wy1+bKIBywc/mRCJL3TSu4WcsT3+emMsE/5/yDRrwCewMWX8KRz98lh+PUYtOEDWg
eT7yGmZmIlIOb4WysBJZmY0PgFH55J1J370ABuDcI8xlFj+rK/XsCZrioa6R0nIAcuVIxvCGle3a
Rm9vd3gk+7FWXpzSMCIRuJC7bMJJGaPNKT9pidfUZ7znePbFYYzEelERCm4iM/AK7cTi4PK1CPxP
pEihWix0VfT8s/5nyrUqOzUeVhI0G5CaJwFR5gJeiW0yCD1bzhQg8MolRXvqmcuYV+TM0eXhx4mx
W7EUM0B/b/UJCZDPCHBOftoluHkbxoFnmjDb9Jgv6NAhgkPYczCDjrfMbIjtW9VKxOquHUepLIgv
80qzEGG51ZmOBHBsyLkFcvwIm3XakaWx2/DUhPiQfw4t2zgYmDaP+5B3IoxJ2OsbdXSij7BgEpnW
aIr2OVc/eIypffaIIWWsS9DXeXN5MKnPcfdpK9Jo7rT095a31Z4OFJ7+V1UUggGxKfvZ5N7vLwRe
5qzS1Z+xftPeVE0aQTOak53W7QJvIh5cqF/ykywkXmwSoUrgXAZHCzJzOMdD8hzsLJvREByMkJFc
LAYUm9mLHWqb0ASvc8REB2BXPLQLCGNH1ZPzhwAYda5csBJzZbMxs5sQ3LE6SD28MAdFfsSZue98
5vQcM2fa2++HRPzg11YtlaLgcRReV0RCTEljJHXtnw8sy3dV8lRKw5lffugYvBld3ut9NN9/4bHv
5LxyMj0GbWYatOPeaj2XadqCM4i7kXSrhNQGaLzYcxB9++URUv8NvXBuMhCIXdRnHsvBbpd76REV
c7Ova7H1dljvikOkcySTugTAs+qA+NYsktj1B+WgFwz/xzFomKLM5JNNZJMMHFqAA/wBoleaPCwl
jjeXhVDmF5ELaHCqBQ4wPS1BqREfihZBySnfknha74q0T01A9fztB6DEuVvB5l9kSP0wHZH34tSw
wNFhxxIsGuDVhqLZ/mhzcIU9inJwaSgUzlyxP7XpvbhSRFEQA5voASLAalyyKQ5lkVeh25MDV2B6
cPygZZbLSnBfnYHeHnMQZOAtDIzs8+hN1Ytx3YoXtRdE6VBfz2w9Spm70iD63C/cSunrIBAwGAyu
/0jbI/QjcNnT/PCGypia01EybyRSlgDFHHeXc5kViS76iqddXlGOLcykg+BOdAsevCR/4fls64e5
If6fx328rrL8Iz8yLqH0fcU6or2b53FgWURUC8Oe01XG+iLX+XVNPjh0s2Jln7oSkUsFS9xa5XZe
9eUQ5khDdUE3WqWGdvoQrOFEEZnBYIsldt6ACq6uze9UbVq0RwG4f26h3/2vlp5CoiX5r7kcVd8M
PfmgF+jFJVnyKkBjTUg0DfzvLIb/V7/0EdazwX/jel+qI//Ob20lZZXDredM2CaQE/WDdcwbXcOX
wYN53YxJ95OksvFfe4rMxKhWavu1kgHabmIE3FZfb0o/1wfPLPDyrlXtHjQRVPqyu3dvS/R7aqbW
FnBxZcwTnH2r/5s2IwjOz6XNYa98Jtc/6888nk9MaaKfknQC1xDf5fah/WwpZQodE9fiwSTvB4TB
y2A+7S642IfG2Fm5xEOJ8cnnl/EekQrX8U9Tm5vz4+1KFt71xQU9s/iLZH7s3QVWOnn5aNfOhKK4
CTTNkD1marq8xcGSwdSc+vhbeHBp16aNjD52IwlQCM9MoJJ5zIPCmSEgg5RZA2E0YC0AiMQyAJtE
tAzIt7aC+Qqe6IBSXwI9FQtiFLqu1z3BeIP9MGl9XQwjSA15+8WAM6t3KOsYC+V4JfsoefY9lY56
xyFBHaYKw5ZWDo5BNYje3DGuzDOhDemJSLQRMZUlqPsILgDqusfIa+clQulDl0yJFSsJfk0Z2juJ
9dTB+bjA/ZTiCwmnVN3OOpW6AW6IFyO8d4gVNzEmcoKtpsPpcGhFgLDTHjlZYzeMEYW/CBp7Hqxl
9wPREShyFKKJ4S5TsUFze8l5iJP+O/jb6EomWhp/EZmt1vs0edij7xAZb7D1qRVzK70+M/NPvr90
jPwYl9hXpjueK21O2yfcP9dH7AsdxnSpFHsnzowKCvdWTNIaQ/7fxsjYgh6UkRzIyCi362ODIcxr
TyzItnO/csUcZfauI1DyfIfcGq1x+UM8/AkMkFE9Yu3XRVrK2sLxpBq54GI7Tr+Bv/wGpX012zJ/
6I1i9EkUYAiS7Zv30hM0AxBwKCXDF7qbiAX0b5+RYhwaMOAKTCsOkcr6vbv1xvHacK6KCldldykk
vRXqt7bucIYDwDLPVjQ0yExW2UPVg9+VKAytW6l4BkUsB3AbNA18beFzLsScyyppKgvn9djs+AED
EXzct7lLgcs0ugnyCdUA/LmN0mgFSDkbMxEbIgO/hs7bdfmvAtdC7YxIwtNNIOvdo2L7G1u/6f2d
m/GQMBT41U4NCstPFdG8Kp81DYovKrTrYStJ5wATcEFNjnStDWHJZtVgikaT8TNUACLAkdV+tqki
7esDTGrSwo8TJ/znStNlHgN19u/sqoZRGEN+D5fUbQR9Fp+tfWa43LyQg05CJs635FCIXgOxTGyN
RHYfKFOE0D5WzHdXLcedMXsl9RfFeqe+q+k9PSG/uFIiUN3qM1ZZdFRBCtsFoSF5eYHXRIi5bUrj
ry+b2O/Fw6yi68E89ar+z8HdsJrFAmmXV6K/tn+b6ISEnTT8vl9sKQiaPB4NeOq7cjO+o3rdcGoy
qT4Z2+U3wbnIq/04nY/oXteC1GXDqHWPsjFqP8MJYxpFiXMc/Wq+Dodi2bm6mVzQMO70HBtuqSeu
2h2yFvRz/MR6s2wvss7fkRJIhttUbl3QTrqjoOCCef4EGCPFG7NfrpdwA+NGnH0SodngduLrSKf1
Ei8fRi5NeWP4dTlW2Ue76+qE1Z7QaHHRA5GmKQDspiXdlRxvDD3HCzFTh+sYgwP2EU/XjxcJzKP5
BkBGR5g5+hVfpynZLQhXLZrU5E+9YKfQyoxWmzeculS33FJnd/0rZt1OO+EHyT8LZHXMfTeaorhf
8qNwEBQvW5cG8Zc69j3ngYBCtZ3D4LB45mMA2WNFKQwKdrVmHkP3wOcOT4moDlJCkONDkoB6x8Es
ngwmwriWfGQLSlLl0Q/mgHyIpahBbMBFBqF8EHM/XQOdWRqPkeIVZe2Cvkymic6cfumhYEsZ/Vq5
rRRWBO7WS5GZ982ROHjk0hrcr/+RvFauv4dsvNHrlFgcrD+JfQ5yhd09e7y9EFymB7BtwsiDs+W0
g40yJSRrVbkgy4NRUd6reZ/4HhYCttiRzxjMJQS+8UDkyAxAaMrhTQToFA0p5ncyMfgLUmg8uoFF
jC1E3zRqme6IfxfY2Ygj9oNemj1UFJ/2vsjCjqFzB5l+PChTI91LXNXxTA3KY2B6wVS+M1urvQNN
aWXpGwFzQYMYXG7xz0pnUhAXirDxVdvckzfADcZDjhpVyxy6w6oJSAlQf98Ifvpd39hxDRiA94OI
76R2JJkObWLWuxHL4dU4ibYkp+L2SFMwd79vU9tk0kMHvM6nc7nhySSeAiDNebTMFM/yumz/g9Fr
NtaRitODezBAQAFtnjIxomMyBS+1ERG8wQ4/Mvvdhdwym6x5l5DiMRkPaGyLhcrWMGx2iBJBCNjx
iklmv7CVBmwkcW0jdcc+CoReWBEw0ppCJImkNMZjY/ucCzq/s4lh6t43LXN3HVoc2xyYoBW1vV3T
jvpnYQziWCsZ8UbdxNqGbSDjz3tDsSIpziyI41h7dgTrPerEEK0XmX0y++QBkLFY1ECFYlg9ZeI5
swHnbH+/FRzTUbLqLDZRa+WE9/VpdMBGInOWXWjuO7vI5iraeU97Ysd6PKQIRATzzhkYC0tsBgqQ
vibU8CtoU2/dHik2I48rN6UZnUMADYi8gVziZCvMJb878Opl23Ju1i46pc0e03/KRlLtVFMcfP3/
CF7f5l3ljgZy24yWRlv1joq050baSpcH86AT+areDwmu0KZtEJMpSMEWhynukG4qzFN3O4VP5aj/
5I+hXkFwrOnQXvvpCFg+AJHpzKTpjh9+1JdZOsH0thpeCQ/QTa4LFiU+mVjpf0/fnQBhqJ+DTpS4
+LpZBx8GMQ7ly3ohDXWmUyiqAvel3v5QppgIxiWRIbeYZV2+kMohxQPfMKnrRPrSGgq3MkDIzFR2
F4TCLqqcOOtY4gsd+t2e4bs0Ufl5U4lVV56j0cga3UMnYXjt/0SwTEPN7mK7y0r8tDE6WhVMbi8A
Tpqa88HPvWcDByOYgE3MqWbemXH8d/HA0kYXHQTtDqnqhdyvlZh7ElZMO8REnBJRQw7xFofwYsEQ
cZNzUsJMLatAfvVKyUdvDCZ8YpxNc8Rem8c76/WcM2gOXp7henAytBTVyycmMpMmFXKl8cBG3xLC
/vG6JOJylWH3CXC5VPkIvrxpgLU7b+qS+Io8vtKwiwy8uM8fZMgt5LRc4Cuw6hVINRFO+Ef5x4xq
RpbIE0xLXLSLvisBASjlY/LwDreXQ/AyHTK9+Dtx9U/KfrlscLKva2fW1Ms7RWdgN8oRkFP6pFZy
x20K/8L9r4IGfbI3e3P7d77UCLCpf/sbcwIvIfSENL15V+tM+S11u2rBMt58a3fAmJVVS75wJ+Eo
++PgAwRZEk2Ijv/vQILmWnsK6i2cf/9NhpwemGZyG6IL/mrGmoLM3RePjLcECZUtw+DO1JRucv2X
ruD2MHr0V2KHBiDFrnNEnAWf3by6F1ZQ4hqQdglPSD5uTN3Xw5GWng/U911DCi2E1Yx+ZOvMpPMP
K4vu7xgeDV7KMpgZD2bMUrsdavvBLXDigg6DdEuQjZ1aS3QBOlM9gxGQ0kmv0YbJUnF0wHKtpoeN
XGum9ySP0o12gbQQK8lwuMcwI+13Dckp8k753MyfnJs9pOr/sgslsslDBRjp/3QbXKvzYYpSuJ/U
owLTOxOWGumg7voJwfbTt5uc5nN6zkvAmiDdCS9wfgbcdCX28V14/gINrpb7KCcucmK3+l5c7o27
fhXVv+THRPWIt/UdTp1Vd5yKYDl4GecnerO70VTJOis/dxXGIsy9qdNrZKs/sgSwqoL1inbjbenb
de/B4Ge9yIrrTobTyhuTqQKT7gi2M2UHKkSF8vqaVUxY3/UEf7+4I3CMsisQgzAllJymIpI+iNZF
WzIHz5Ojicq37jkFMr2Hm5AKiPs7YWV7RvMRNPf7wSG9S9mj9ZPM8ymWDlzKPOVEJV2BqjORXTwZ
30Uw04M+FL5etE40irDp0sLUVLrvHuVhda0Qhu1ZtOXFWe/fAAfLTrZ0RDqgUWrlmcvPlOp27BvW
03IyF03+1kw0di09U4XcQvMw/fQUOQM6ea4WDNkfBydJScI63yk4mXuAvMBe56O4tifESwxqi7CH
HFbV/xikhB8JUnI9ES4GiBQTqcCg0kGpUBX/NQg35afGxmG6n6iK8QCEks1hd1D5rB68Ho32x6h1
gN/U5Uy145cD2kxdimCLrDvdorBEwuDUzKsGGI1/wby7kC6Dm+L2CmG6SXljLYTEAe/sL249zLly
SPy7HtuVL7d52NDfkAtqCxSsjZsUC1/6K4gtCFXa7y0SHgYWFYzp4atPVbhtKjzwkjEJtCL0MsEc
0M21IPhdaXrW19O3OOuD1RtA5itIQaed/TzbiP5tmWXWggSu+ScmbLya3SOHc1H0B+2btg74Tx54
EyS32y1tzE26gu1b2lnBAYTvezNIMzx2/yGQFX6slu5KX3NVESff2u7jw5nn7zoGI8LV2aZBKBND
Bs7RMWw2Q9DZoUGxVzbyryIkO9ZH3KBjAWOvq5Cg5l3itXbDDUTMrc21Cdtc30nP92IkAaAlwKy3
neyrTg59rSkviKCKCrXTG4ZB/aGXvnOOaLwfFrfgQYYqfyR/UpjKID8htzJSbNfe+vGRgGalY/tQ
to323+cX0fbxd//gkEmKvKNXgQz8qZpjX8SIg9KgZ3DQbzAo7T3l+X1rrDPfTtp40ovQRfjGiou4
+ssuZFjZxSh/LbWo19JiJZkIUuJwfovF+GTx2LPaBZbwpAwBn3zsCgzS+LTieFqZrldjM/381CG0
JMDCb5vnH1Tlqeek1i5A1XM7A9ZM0a1UqL8Amd3Czk/5B2K0LCrenrCTMzhjjCExPMUrlwKBh/tu
7On0Tnxg135lKZKPURmcBHHXk/p1NQj6TrP5WNHyNAhPtniFtvlLNZaPN6YXcXr+zhaDva/yOViy
/n+S92wf5XlukrnZKPFwnIQ979RmE7JxbS2AUUqFOnC/pzNFUHOhLbQNXSq5dkz1X1+t1p9cg5cw
lsplAwHGuiTsuraKFkHpm9dOHSCwemcfpgSEP3f9DA1KrwTxqWFpDbmNme5TFD6MEkc4eZCNG5tM
2WIjP6NOEBU0U1nqE4QTH23WXqf7i7UEI+GMRAfEZUGQUL6xxm8yBom3cz29FRqucITXqGGFFyRl
6KcOlmCDLu9zRrHndBvqGDslFpscrvAgofo17sb0JM5wZFaq7q7ZMpvhDlawsbT581IrW29txme7
NPgHyuo1YBv19ctJz4GLIGTV6i/HfTAF9dK53fomCuuQYpTTM5+SJtZByB8sNU70JUiSel0jvrwU
GMXn8Z87eoJLP560cMr8NKwDeUdRvIZ2cIha9alSMtwBJdNKhDFe+IEgZiMbj5MmjRq1oY/wcOyw
4AQukXJ5lmtxmNN22tlN9JY1MMjcNp38NYAYLzVqVwOsSRkqbQpgltuZiUpzqQjLHPZcU0ccv7Ln
nmVpYfFu7a7InNGjVLIqXNW4i6hO0ezwTCxFMcsUE9wasJBOPQTKnxBBg/q3luTVDZOytoCKfP2G
yHs8zyc+Mc4xFE7GTzkQ1kJbHyjl4+nYFjEuCZ+SJkskoVGXsef2D+A7oCwS8iRyCp0sACJnMYlP
nXHTkqe2Iq75ohZAJHR76T0rokpAGvjZCvTpbYIFbO8qHr1udO0Sq6RdxCx9LmgvzkxF/0HGbPEq
hf5yfduXw5aYxd5cJ96YLHvLjOSitIfYYsTGx2nOEq2disUJF/2KIs8o57YH4KAsRMmNXD7S4f+n
pc7Kapt9nL39YvsTXk31o6WKnMA0DsGLzd4fogBIQsxhMdvBtA5PSZdAQpMegkNDP2jytTIxv9L4
OFTs4AptgHM+aiu3krFSvfxxqiPIAIFddFOwkv8aQWNEC5msBCPvKurOLPbcLlkV3RWRp3uJWD5C
Ol5kgySvcc705fGR4t1VQEhp3tfBrFhRx4FIrAZdNs6VUlzRFxL1XgPbIS3vbGRPkTDbWIvWoHBA
s3EOOfTziFBRZHAW+RkDzjYXunlP6okeXHq2wrBpC6bv59K6Wsbika2fgH8TzcW2WjAAr/s2oGBf
1V+hlrdo9ug0GDSJgd8F5svYREet5CuPBCeQrNHN1Bpy+B3r+Le9fYnQ5uinTjPx9nrsWt6zLFVS
MxFhlXBIOt7U4bAn7Zfss6oZdMq41b7PAqeQvDFm9Vkcj1235sPip4lFOkZ7hV4F9xrw1kcGTS4U
H+yfPNhJxeQEI2/qW2X+d/qaxO6PnFwvYwOL/IUZhlfYxowjWs9p1l5iUDyQfoha9GlS7oGH2XIF
+aoUPE/Y57bJ7r7mmnSElsy1hezNWzyjkbJ+xPO9C5ae5jCPAen1yUvtePSJ+WpiMXlOsxKaYR6E
9l5zynOCr4inrI3YSHZrCR6nItzjwOLx5W/4Edq5CDyztQ/yYrehhxfO1MSkyP0/oHSkAd7A0NQ6
Vd5OAp1cbbBD/dMWGZQKOv3hMuh9zDmm+CRgGbxFMql20KqcJRJifgKeXHWYHm/u6Jjtpoidb934
ivy0dXSNZaTm2mkH91uC0ty3zCLRVZU8sPheDtxCBJZ95CPm8kA7igAk7a7XmOoVzqPtI6vBNLM0
1rvoknD3KU4/l8vyqDLiAq0b8Hzt6IYXXsJzdQM5PiXHYIlVlvbkzxjU3ceoWktu+M0Rt7KFoErc
oKaI9fGwJkjyhaHcBIay8trLYgQttif/Vyp7MiTohxymXyHPDdkLqcuk6q4HbJm24SyjP4fV01vX
f1AWb69iPj2C8jw3xy+4uDlRNqi+QTFwg9A6cPX+pA/o2PeVxhiNjFWUca52QydPP1Xm+amni1JZ
8RqHgEot4a0jwktcwJAFghtOxPbT+zE7nA+ND6SJIyIirMIMwJ3o/A4g4gakjfPZBnE5CFC6++kG
yqxTyuaMYM+9Z5oobqWOmtHbFtAY6Nr6dhb5VHOKr8yKT9MIJzif7zSXUjyVk1yiEp/Uve5qIMo0
dTewJzAj7K8mP2CJKLyx0Meu9H4GspDCZ59jBWZQO9S1+vpL10mTpwOuU72PJSfFfOqlK89BLUcE
hw==
`protect end_protected

