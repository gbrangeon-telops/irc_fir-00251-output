

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
OJrNPv25gxVf6MOkMLDXm9qPvzcLiFn6cGPtPoJyX0DRSMUs1CiCHluul8VfoMGYUnRu9NzC2pDa
fD3Q+Cro6g==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
OO53+YxV1fz+fdQXiBafTL0TfU0s578DnGOkBDgcp0ZiS8qBHyL1R2PISafYfK37QZ2xP9F0gTav
+sG2DKzZYRShUhSDZBSgMOYpY7yZxYTXlswORtjPSorUAG9VDaJFPSJUqemfgu4AY+n/BsniNBx4
zqFaZSDmDQebEViRgn0=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Qtwd1yFLlmEutFKAPe2eqNz2v7W0I1lWfaUYyRoJyXavTq0FDRoJFjh1vw8Id+dlXsCh4QCKBOe5
q6ztRPULauE2vnffEDrTLD6uStkKikAcWpHaB5kHv8W/IU3+JNz65HQM8j8hOwGUzUSaTQzI6Edd
Kua78SuOo2L/RNS2CApKLh4UlLjlkL69KZuDAj8Ds+wPTUwjY2h3tf4V0N6PH8lPAy9xJk9S3EgQ
ni8vjkjW6lK8he+zqjEtOf7IEGhelGexSOLg0dP3NDhMEcaxfcI7Zo8kOCl3C+GMy2w3TEyTZkQr
3WrfN9WllC++Z6rNtRNAqHVgNVA7hObPvyuA/w==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Y5YBoFz+YhLFw0DE8aie27jXEk9zfvZg7zgS29dcVa80RbYJrtSDIAboa1ixJiDhfiME1gY5XfYR
MSxbx3I2ZAkTI/5DwNAjKseDEksXdqu1CBQcg+U5NxNg5wWuw+vr6DqkJMxvZoI9BhjAErRu+2EZ
DgyTp7XS17TjzQ/Lk3I=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
amEW+kSm8JLnUlmLoRCPt0pU7eCAirRawwzTZA3XEOaldjEiNg3FqPsvTGL5ScrzO4MhYsVv9max
1PQJ/lU1FLIUBgG3vy1UPm9QWkUIWp2rve3mDkSCfvDRku+GIP+/ziqovgiDyF46b73fS7Mrb40P
ha2QhSaORrSFucLp3v+D7rdh8lKmMq3YY+qxM1KZEpdfbausR1NP2yVxQP/t1g0w2pAjiWQM7wT5
6xmmRvYxl+7EuZQkxaCLozCO1ELg5LiuQuDVfKRWPdTIjtVbbBvnn/eTARAw8sh6+JXXfmhauCWF
cGkCTU9noi1D4Z3I/hvgJ8IXztgyejVNBMRBwQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 7392)
`protect data_block
X2La9kkXjAi190k6By3eGphhSyPHgg1XwkdAViodDqcyJ5CTP+WhFQZlvqG5/Zd+2ggtnMwRowOu
q3ZcWl4qNHuP2SQkI7kPeq6IVTPi0jqSdvLTRXEQqZsBlTjyS63FlWrQHyyIiG66PvRKMjL73NBN
peULtexdwqTMMWNjM+Pg/xey08kJH5opXnU4FfE1TJn7htCx+AMK7MOkFTo+q/Q5sA0fU3xyOxcd
WV+5LjC3ERg5ViFefGH93znfbj7pi+wuN1wNy7nzzgY+yQUIlWqVY6hMhUIacQJ9t0saCPsFo9F+
0rp9A3zqhz0BC/zhcg/hzR7jlnZHaFK44GpUeWvXKpnq4K1Hl4IWxKAmxDgLkXw6hlhRC+CbI/fh
UBvfGdwF65DLRsiFR8t8rnXFmxZQkvYtEeMtGqGcRDaGBaNkDZNBVnqf38S2Q59yTelMfQEZhcVh
iTCFUK0GcRAuPmN0SLQCchbn5ChNslP6OOzBL1lACtFrT2fC0QwFlJUnKBHqY0mEHENGBCn41h05
oRzbVeeYAEjWR5bqXVFsYNe56lHLOKLgU0we+Wof7+r9ITNHEGvuFvt02wMoqiQloxscb4ri1Djo
RzveBrmLT7PFiK3H5peR7ycX9a4dkXT7WDCv+KRAuOKR2OsMG/RICWFAe35/CrFxpMCTrT3LeJMa
ZatZkHefdHe0G9w/ztg9RhPhluR96eR3gdEnCYOlrFHAyFJZGRpIpkdMMaGEFqZpkPGkneHXOzl4
lQtRZVn8jh/xtUF/E5gX5MFChICuPuDl17N9me9JbBswnB0LUwaDJ9iuA5bDqKOsEAQ8vVGX62j8
yFdkJpF4xB9npkVMvvCcBhH5qPOQlAX1qHccAFmgaRTH+M0V8t8Tqno/OYutWrKSpxw22Hkprf4u
pXUU5jqKMX+kF64Ln5aOfrm2NBvWg5aOCGX+2FQP5Ey9evKJQF97AkjvfuMHt+I+WHpxiVM9ghWM
LdXFMdb+Jd4kdqKSM6xVAxV3sz5g6YWCamXqRyEkEXuM60h9Gkje8GXwIxqUnvE1Pc1yhrmbYGAp
MVavVqnoUJRjfHi0WcTNQ/ZstbmOuXppssOQl6buAAKoDEAMnDa+iNi48VTvjM/popqeA/tLJ4nd
Bw7+3nOTbJ4U9tEeGniJI9P30+q8Dw4sUOURmaTIY9VMSbvG/pSVn/KxJAEudxTkAhMFCCp4QR3c
uIicKu/g0NHj9pnx0nsO/jxPWZN9sK/gqBrhfemH5tlkO+pHkmeNDo4CRW66756Puj/HgUvmtEG0
RBV52LaboXT9tlLnjU9AE3+OQNcooe5qdXjnK2aeIo+8ZFHNk0vuQQcJWJ1XuRB+VsEo0JHf/9/0
Tnsu3ROHHPJiwe0DZ/u11IcMuhHdWj2TxCZdvzeYIeV8JQ+4nTmUIVc3BYvx52q7f3KXOlv31Rb8
vqYkY6MhqzMrrbIa893mpln4c4M3E0Db6x5ABMDWecn4SA7dgtI2KMPeWkZe10G0c+UrOrWThAlt
eEGmn1htO8UZfynMF+6bzSlu+iODU+PkyRSt2o5ZO+Cv28eNPFU5tU8oEduf0MPtMkGJJlVbe2bx
vj8Vss/VDuFJzJts3tjIBkqSlBEbADA+Tz63+9qVX0Wp+mUo0ahi4hxm1luKaz4OlEnh5It5GeZk
FMhMaxsf1bU4ooruwW3rcb+esDoHhWiCxsWJQMS7tIOT2bsVlztQ1fxTVM5CBbpadQ8gFWZTHvWW
0OUWB9ewBSPHv7/PwSG8jrl/PioAePT9raHdfIhjQ9ax9TEyqwxkeFzbGBanQxd5ze0WhJIQT8hw
UcUw10OGLkzSXcLZWP3lbZs9MH+pI9gYK+6UVN2HBQVcHuEZhV3Q2kbTxBM9bDJdm4YbW/Cq1VsD
vT8Cr+z/D0X5lHv8ZdH/UoHviGS6+4/ShllK19vzif4Hp/59T25T7Qp9jyDdopHOJu9ncBoC+HKd
JYOz117nWgoFEvuONuqPAouz3qmNHg3PYAbWMTXL1czsby8xjp5Q5vakrNoLAffVP961K3pK5AVa
kp+HbIt65tWVuAZecurShp2Zx1AR3cZS/7dj9a/Qedm/RvDrfSV/WR54NKCikfNdkDd55XeVw2ov
ZJNF0VlQl8ArfX+xidVkwQZA9JdTHv4qfxY4bZJM4ZiNAswVF8G/yVdnZe9ayzaVSdj1rz+5zytE
aEeBwZ6/QRbHbW1uJ7Yh7+J/r5Gv8YtNDsaC8nOtB9LRp5pwzjMno0Wjr4VjDV45Va04uZnoCodP
ZFO/vPDtFKRbGsiZfg2THesj209IcwvjHVuFeRYZxwaac081h80EcyOmhdDmrlPhBnmuP+XPflrZ
Kpw0ZnaLHTmoE//hqCARTYwWv59XX7pT7Urt5PwCXxzuLRUmozIUG9jdVJR8LK6HriEOYDH3cG7Q
gfWQe/c/NhhjwYMDRoQRh9TvgWPV0SMF9BoJuzG0iiNOCaeelNwjd1Fgb+zQBYHZIoM3+50SG2FK
k7FznwFkrfH8AdIuCvb/k1IFWBXlZWfSMd3MQXabgd0E4OxGQDk9x+ccBhVa6FrKiy6iYZf7bT2h
vJbh+NQx54Ua6Y2u2IK7NM9SggBfXvJ3dPfvO9RnET2hHh2hictlAjSrKhg0sLKs7qEVGDcFMSIs
nnMqTVdkjqsDDlgPA4za2UWpX1ysQ8Fl4iSztLxGtH9WGFpnnTVNp1C74iTCYW/qFiSnJN/q1xFC
b/wPawjz4M3Oe6SG3Sgli9jAPGdjs4onXwfoTbKHVRgKoa7JzaZhvPoG+/1PCgiXLZEtQrTYuumh
LzqM7HCD9c5q+MS7vFbK7T7IikLuAbAu3QaLuU56iDKbmLDQ7cQjbowDyTsh06exBowphG2mEMRn
GG6XXbA1LTsXV0e58c40sydlDxZU7YOPa6IcGVpPKGglDUfF5NUdqXGHTPM9OSaKDu+TcqO93Baj
F9Fjsmm2uLm4GqURSYTWzzCs4BYEiMOTiWO7B+I+3k9a7ORu/jof+HIi72ILUhecIn2vo6ue8X5U
hWz5Fu2ymsRXv5e8NXosCchU/jPWlM9uVdL0bhhQo1HI2fnDYCNtSAd7hKjQaed5virpm+Jdn/DT
YfgPCvSXGfzOOc4iK+A0LjxNLGcvLBUjc3GcAHr4tbGotfVuBqw3eaYIAqOSyF95e08a+CqNeCFW
huzDpyHsBBQ5kICma8XesEMBk2KgLqGKNKiIrf10/cHlZd04qRPYXOmFIasCvuy7X5hMDDbdSPjY
CW/3YMhUoCUqTbAr+gSltUYV4XQxQGzJqKVV+xP+H//YykjGcd4E1/ergvEB5PRKL5eBvxf1Nisb
B0PD+2KO4GUIcU5GVZgq6foQbRunKYtcki81W/gbpLehGwFFz7uwsWCFWvMZXKMMP+R7PWQP8LVB
+1e6CPuIRvtjLofMQRBRdkevShW3k65/c7d1UQnB9+vSOGCS0ro3wSekcaXUpp32kc5a0mD6b0O8
7dTzrAyr5POOA1iDJZL44JmRrJjUM/ZC5PIIWOG/URdpYmo/pUk5JhXmB7Uqu8g9G7K3Lf+RzWjC
izi14eGe/b3iM40ZSgdrFiJSdA4GOYp5xLnhlTgeHmAGWiSd4K1ijSxBzxC2jwt29zOkRwl4yHdc
rPR9QzrrbN2TdkyTwX6cNZFEVOTZjS89OcVcvtO92bKGonIQLcjz3eUOPEXcD6TfN4e3wQzUYoQt
juWHWo7N08ETsoI4c2p8U7o1V02xdOfdVkXpssBMKmtQb6ZCTLq3ntKOch7rGnyThrS7ViycxwMj
gOdCRPHbBahtDxPLAZgdH3AP78nr7E+a0fJhFNYqBuDTXbd/GVJrEqOsv1DlADff0Tt6DytN2aEL
+4CJWNT3ULT6AOyA3iaxZSBeTmFfoFrTsRtTBLwEwvvBHc2q6HjixCLphX9+GuOlVTnqulxXfcMA
9S2agdO8yL4YczlhFGjc+vsmQXNdLsJzl92KgfsQlM/m4oPK4YUcPvzNp/EK4/3Hu4DGh9hFBxv/
yQKKUcsNbL/ud3XH4JyqmhLtj8YKabPEiowwtKrhpIyiJ3ja2k+kgChI61v4nl7kHQ3sZ7OAd5oC
mrTBVZVYDjH44LeSS3FMpBqYijDIkvBoSKdbjzvEFjI1+jSdgX0md8xh2lFIbVzH+fI/6FyDpVGt
sDyii46+/V2PCU6GUXYgJItsvzhRJBrKtzvBm8p6Z56JyBaOEhx43IrGQ0pdYBxfam5RFy/yjWtz
gCUTguVKiCO67qPCUAzIjr7K78+d7AbqBPpXE83GZvaMeqGL3c8utHL9xp809LBQkLBILkoZ21Pi
w3g0Lt9bw4qVMvshJCO3RORNVfmNm2KSMeBq112GMryVj3kB+LTREOke+5AZo/1Xxtmutf1iMYbn
0XG/XoP5bkmWsOWbMczckSmtgGKIBvG6E/YjjMTKVLn1Kn/2oKAhD8Jz+S8V0Tsitf7w/q+1NYFG
SYG70ChZMvmpRbz2hGx6qsJYkt/b3Wk13ExwCscD6Pbzn9648UyUF4yaw2DMB9LybitvqY3y+5dW
ITV7aKO9aN+0okTVoifcvL3jwe6nYf/953CP25fUCSNq6mZZOhsIymfUsxDwFOC173EZqxFfa17E
3EBL827SMs5UBRxDRspZWTX8rw5pkdxszXEe1doQJrFRDQ+0TcadozNCFEuS5/KxUhWUJLICWrA3
T9lJmRuPaw77CqW8pHUHDXahNb+DQ8VweuNXpr5wYZO1H8MWu+2dXmx1LTjxCJpAht3TcuHa8HS5
tUrzmQUdc/kyq/3wv2edqSI5vCqRQ1MN5wIZW/pb4ASDo/10Sb7OO9hDx+VNUK1GF1olSTI7p/OU
4enhP/ir6I9oSSIYEdzJEh70AcPCAgK/OhBZbf47mpUSswM4sqxoxlDokQNaiZ6Va44Ir8jOEAox
DI6P20SnT07FoB6TcwEmZoH6GzaisYw5C8kFMhUXd++JWDhoPe+1LYiyYRpTRZXZDs00hbJu1p7d
KCGuD8FgyhkSrevTJS3IwE3KhI7aLaN9MbT01CfvQ+K0zLqlHQrvpHV6KuY55pfQCl/HLEb+YGll
zUCIBZ9frh7rzVY65m7kc+XbWppNebWgGfHUK0B8RMWDDaNV1vOK1OBnlqIW0IN10jf+0lWzxvex
aB2XEgXtLuNyWRyZ1HrCbxSxiM4DToVLiuJnJTzJ6MxxDrvxA+GvzvfsMk5KlvZX/7wQVjrEjypW
qk55MOHKx3W/713w4acxQznoCpaTvcwbH8cl8psywI/Hy4N5vQJSy4UeIAyCEWTCi9h1+Oy4NSrf
zrSo56Aa6vXFgMR2MUilmd23t8VzniC4KNRgJuJynhUFdVAgNLBfqcViLBDiWrZ3dcTANNkM91pr
5hgomKXjUO5zh6RPx/Pjo+JtFyRGThg9MXa9CAMZRb1ssgOx7fADD+aUSBC+PSXKi89tfo+WpR8e
NPbTLxZoMkrokSaInEo7gLrisUJ+rO5lei5SR0jELVwbbtqMMqZPuiAZT7iMBxCj4h0R4IiVBAcY
PAgdeXUH60lp0aXv6ooOsh1NWBLhv02lqZ0YkrEndK7rvhxEGrAObLSdjNoGb7VAEclhJeI8JfQa
oWOR7R05kcIksJTLxvEx6SKmd+0l36wbORwu5NrITCqLaXcxCwBBd90qc6sUf0KeNn360iZCKcm2
cDZq76DetEqXSaxsELiNNP3wN8pmM/O91frq0qnimpSod8SaaEX5eZ7+2IgBdeW1LXiePQ7iYSFj
te30+5FR1hej9P4W7EnkbYTCWTW5iG99nhpT4JDoLDXOa+u7w/d/OPFo7BZ2X8/1RnQI516ukK7t
nM1Z39X7JMHQx8tYX/WT3nTOMrYzs2abuR/hGgAbKdNO307HanU4xuc84Uax6FSfaC/oQAaIPw8P
FamILNbrunXOtyI3Jv/RzPqMXlZsfX+Ok17qwMB8d6xTGwu/TCW2wWPTmiTi9Tf+0mXOt3LbBhnb
DVq3Fh5zK7PWGPhrRJIicv6m29d82krr9sbifdEbIjC0svRUpWO9rObSJ0LQiT96BsNLrbsxU4uo
Mha/K7w4ETipG2pCqIvh9N7uwLuVb5tH9nrhkzfpaxitx6egTRg+00+bXlW87jyKH5v8SHsWt0o6
QvOY5SUyobJWOSxpU9Tu/KMHHPeLPwFUBbSJrmiZBrKuRktNzFwxq/lg7bufYMhZrNuWa5kyTNdU
DA/0FRenwTRyLtd079kKHNEEKWdUsdrtx595uZCSy5DiNaE/mZV7ZgRnnu5nOxzVWdyhetFMmtrZ
21wI0Tdw/rACkM2YyY0ipQrUICzwVw4anh2w9rCj0qSrE3QlQvqWCpRpTnD5VnqwkocDIZB13x6u
FPSr3Ppa5Opu/OVR5mbHPe002gxoDBpDEwmaISyN2TT3qdlrSLFSGf0h4Q3tFXa1NXdtA//0JjxF
wlghQV8z6GymmYm+z8U7S2QxueX8rZSN92k7b6l7ye6nCi2n24rHtyWjN0YCb2/IAgWl3sEGG/ir
8Bo0EKYw28jPbNfE2yYRBVbcfsCSl9R2R+eMZU2mUFgX13X0Emg2RkOyEKgfqlF5jOLYAXv8Py+4
hFtrhtDNbc+5EC+x3TWjE5BCkWG9sPQJexDnjzyEeuB9RVGGRDC//5zgTrDY0/E3l4woUcgvr4DL
kNfMgu1WNduEPq7+5YpY/SkOPoHinTwUMxIVMumZiutMA0SlH4Kj+AUro1w3ag/TX5G3zIKilbqV
MdKywitptP1BQgQjFnoAzN2zm0OyN8pWJPNsjdPFvBPtuxKWETO80qzARaSOKVZys/uMzlD/uTyp
FRxDKdr9dl9X478d4bi43Gj2kgxvAZ4O1Og7MiadvCbi4/3MXQThJ3JF8cVusV0rRBpA5L6qf4fP
XN+LOOf7qvzQPq2PUY9VgrXMk2ONCVZuop4Eba0Z5/Y1zcwJhR3G9O19D++LSPM/mSHokCRZNNQV
L0rU7AbN4I39oKTc0BVRenOAzpZl7hOrAqfDYxgoY5IkyMsT7dWei9amFgY2uGPaGPftGVA/3VFg
qbMkhucfT/XAyQyFV4TtHxxI7MwjeBsIz2wLYd4NMjdP2qxxB10ErhO4ro3S8QeaMGd0Ft6HL0PD
mbZbUpJ8cEfxzm8ovKIOJy2uH8+oHD9jsnQgYrftl3ZtnSSprHS1fzwYkIk2ItBweRtU178iggXV
JqnWo4sFs6cr+Mvz1rJn+e4dUDhTUaLD0FzcPuFyaVefvn/e/3rreaT+KNXIHrjVujkj/lyFDBcN
y21CjWvQpL5gdLNFJWpr41z2pNVERFmXNXF/E3cAJ3F1FoX3Zsbbc8mW8GL08rLOLrEOagQ4KPYi
SP1ht3DOehRlqNJeBPRfjRJqEXbwyqOG9jSXPlKMK/vPbtkwzRFi+AI70FOZzrXD1TPp/qpQYiCf
eqlXlhgErrI1HQIG6TqRWvUxBz52F3lCrt5jHqIdXI6LIXpM83SzzmhW2lXuU7chcd+y8ovWKAaO
L/XFkVeR0WFPfrSPY2ScJuFbFCUdHKPNuHFPK/GsXl7/KfNbUqk9H2oa9Sr75kQFpFw1hCFGR6Bt
3NTCaVAVwb0SI5X+RoqBqhkQnnVUfpvOmQA+ACuhHVPtg6HuYk6s2j4rGNO0Kt61zeAI0iukyqDc
0Ie8Adzm+ce/HbpquUFEb1oX+40z02RrRSSNOQdsL2IGYw+k5xmolj1bo0QGAVfZy/f1dF+uAjQQ
rvk4e3ePiPi2c38L7anY7ojFUeS0C/4DYfnuWP+wuZ20XUFgD94ObbArc1kL42ZRViGZG5D/j4E/
3yS4tfE2XpnGH7uPnFze5Bym1X+FtF+kQDKmCaJuw3T3lb8AZ2KqvY2rBHHnU2mnIWgJcgYCC9cb
oL7QuNRdlBxV14jKYRJRd4xGECvGC9dUd8n/ZQMBN77D4mthuxh+XVUJYtkGgTs4jBZZ2HVIYzIz
fm05HrMkunKcm+6V0QLXQnqH7mlgMfO3Cp3DODp37/KpjvxvenAd42BivE/FsgDsYv6443yFJV2J
nxa33tFdaEVVFjwCL3OJQT31H8JNpJ6TZRyQDvsLAQPFc6dUlV11w7bTm8XnEPUPmU20PTNKfm/K
xDQxus09Ia6TbXDc5sh8qJb6RM6YeRO1Sx2HcEZwK/Ql7ptLKPp5rj9hznLSi4aDJVV1DOrNWwC6
XX2NvVY+26inl9bfW97Mi5+lLzIdvRWP+7Ohh+aINL7ieyEh33rjaQIiIWUh/43lQZqq+IULq2XN
g5LIX28sSHvYZUDmbvREEUPIuJmoMyNjXzV2MbIwWHL6k9V+y3OuuLeTMWc+/YVE5KXtAVQPbhGE
htHNm99ADBtHC82go6qMRX4HrnDPFOO4rTz2jpc5jtRC6/uRmOMWV+9rou+OQKtw4NAdLQUM2pWD
HK5JpU1Pw+IH3xdScXCCXPf8o9bGvLYldNXppDVcDSVVFKa96iZsoMRid51h3i7Lk3Bl7hzxvmE1
UlXP/xFFt+HBKsEajZTzH/Qhydmhw9ncguiEOs5ggZF6JWf2alTmHCTed0INuhksji5ko40k90Qi
nLz8KsGf3aEVG2j0JDCO1vgIqKsQ8NxmRnG8f5dsXBvtby+qzhb+qUFVQTH6nxZZjqOtRn64HmRW
zK5SgcLst3Qay4znH1ngEJIZv5LpVvDjutAYgjzUjnoZM+xqhd968dxY0G85fSbINo/5cRQyXpIh
SjIa2AOOYbHuNphzAHZ6m/QjXbA+soBliI7QJBM8es/ff7xtA88THxpWVz4xVf4LinN2DkyB0Y7U
Kce1NuQKLsnPs1s1rHTpHeq6dCAEZv9/bdOSR1sOOMSSFYBnu9cCxrcPQVDrBn8qkLl/XnOvKFms
4bReKjNmb6eFNbDyIZ3BLNbX00qIJMhrWa1CS4OBmAvZ655cgmA5lWiMOgFd4bqFrCPbaWMRwtFO
ZXiw68lzwmUQdSfAzwDWE2X3t+9D7ru7TUsqFnwST5iz/IcQH8AJMLG/kGe/3NJVs77xX/dWae/w
TcHXcVj8ICGcEpfX1hEWtIVnDkoHe/Gwqq5IPmYiSnaum+e+ebWgsBJAYGR0OypJ35KpptiDIWaM
d/+7YE6GfbhTYHpmiEWyJH3QxPDQHHfrkXwGLGDYx3SaEL9apPlE62Gfg1lia4k9kDi88ZEVSU5Q
qQjRl572WC5Hify6SJd1vgWoNPX+a1QjDcikyVutU/j3PKUBvlm32ebgBiJQCHO5ui0dc2aH5ltt
mTFZoxDlL/SauZvTCRcldF8Hf4ow24jtoTu/mv/z3UeZZzaW59UYl2tLlBVq+JHIE3uQWWm2AGzc
PNcwlv/m9G+2U1dqV1rQKCIEKaDS6IVna/TysCOZUodi1sbAAUzikgKDEZMalkmJZ45EXj1llxlH
3nhyKBYXY5ApZjLIWXCuxKV0hAJekSrhdlt+lJuIgwz1PlsCcnk+E/fZj5LKW2KRm7b7WRwTk/V4
SCht1WqK6C/dj7iHD7CAh/4T6DKKv45D6wXB1qm0PDM4O6TdNrVr5d7bXY0FzOvnRrslEhGb/NkR
wisFwyND6iEiP3BkXl1amk1EWXr9vGrtyk9S+WAkgy58s5et8jLxvDJz8tQrsEpMmBz5BayTrQjZ
2ic6gptgkFzhs8AofVSRB3/LT3lijORqAOgZ1nBi50lAFabhfnnMZt0HG63ddcSDMszs+8i9Mzt6
+aNKlldDZBuVCD+TJ9XsLw20bJtgoI+FFTg8g5DJGsM2l9pt1/Aa4JWbkSm3RMfZmBfRcVrE/mmC
VbRW9FTUYEMdA3Iu7ebGy6AVyk5aiAoXgyHfkS2h9cNWNfbXL4yy
`protect end_protected

