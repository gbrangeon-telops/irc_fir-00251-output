

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
eddlQ1EVBhLWIw/V3Y4jUv/9vIqrPH4OG//oOzrJzxfxJoDe5AYwYtf4Sd3VIdakKHjGWL10tZxJ
4ECEoEAvaw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
eigFAyj6GpLic/D0LIryLMG9xQfLbNW2aTMhx8nk48gxIwiUUV5O0RCi0c3WxlsD0Jm/PNvkmU9f
0bvLBoFrSTxK1CBf237YO6kwoV8FPGCIv6uN0rXS9lJQOPdNh2ZUFAvoavKMegwZ/325WocnFLGE
+YU4kz1iYX1mmK3UsWQ=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
mnusdFYP+cjTwVO+sX1Blw6b4HVRZgRv6yA9tZdzqDv0sG/5WALWkeGj2iueXjyR4cWjsJaH1ItC
lJVwVFFXjpYvHwJ5RnZSqxv5F4MQSqH8KyPuaWJ7fxXpna2BJOvJUmLpfNOHHcM9ZtydeUw0FeC9
iaG6qychgs0JvDwxBvcNWeI54FWlrduydqedwrfELAOgz2Hnkk/tLLl8ktgdmAuHiBSlaAN8i7/7
Tmw44CbQzhCNPl2j2hqobn0a27C2ELHJlqNJpm8TlXqvKo4J8RYyFeM9H9JreJ/8JZ5Gf1n3ys2S
lY+Rp2WYXmq0OKzkZyIfymRWl5zSUC9Q8owcqQ==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
uySJstuqi1YIYxsMDiwNUjJcaDIhlVqhon/QnlfUo3RyDfx9K7bIKjrz+E5jMqOrIwDUZDswr81x
cRDaji9FXOgh4P4INZOlQhXe8T+6WB7arsOA8Ipz2w1V2sV1eY1zPj1AXh27lapbQpMmsim+eCnE
1jY1XASKE/xreD8Glkk=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
l0UqkRkbyGn9mj0GavEkdTUw/Zw8lL7XEPhtCkfsrXvwKb+1KR5+77+E7EhE93Pmbk2awJRlXYwm
D65p2I5aXxW9fMEUNE0pZrhuaqpOOrPdC2bw4gaCcKb2BQm2PHu1PwR+8skPqiaBAqZVoUwFCZE8
LkMHYL9PggokRGZn1pk2O/ghNvl2eJ30v5gmurH3kQ5VEWU71s2ecSWfrCtyS9G29Ke80rPgnbMP
zifmkvX8s5FcVU1LeIe337473lbGtzk/tTh1neIkyiQD0Lkip6Q3stpeftQqI/864FlzKS35OASQ
wgYvGQgHNq1FJbrpROfsgNyTrijicXvjvpG0Gg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 37152)
`protect data_block
E2j8/cGOX54sQDpB9wBD9gu2n4z7oNkdDbQt5enU8zjK0d8QKVMFXCUVBi+V0lcjDAUeaUj7OaP1
Xo1ymzPk1MbUvcRR21pP4AHXMEgXxMfvhfhIW5DNuIXklQg11uDbSUpMLx3BrvOT0uHkaw1shlMs
496eyO2fzhBPq1m51gUtalLVMNxHZiVGPMsmakoAI6GSusJ4WYtTiBVBsVktq9AnI/Zv+DLlsZbu
VApKXIdB5xjPQV4aqyHZQs96EQDmKwcZ0KbHkzo86dnClB1X3ENZ8YNAkgx3LXUeXVRoTsUkXvv2
PXuNPNSAhtyRNku2/x/5VkgkitKSsLRMYAV6sPob55rnfiKxpW4MrSfZo2oVto2/JvXjGw6b+RzJ
/SIgZM8pXbDgzjkBFd7YhN3Ugtvk7+bJjlM8kKhrnRnFmGPZOAXrHrgc5bAAc+P8L017u6iCJefY
N1xiQhLaH9SNu3tM0bKvygLhWUs777iSB/PsedJxzWGin3EWEq/HnN1+XFedaBFUg/lC6JeOzbNP
4WKowkt+7u2A/u8CY8RwB0bMyqCyEyXjBSTJUqWOrMw0hQHea/bElR2NTCAI9DVxZOJNT8uGOPMM
NVKsVGYH6OqNo5dcIXCM92maCbOyPJ/1Q4DBSWtlACSKdr/NaF1BB5uXtcSKy2pvj1pkqu38fQTW
wVvBNqHLwqwjCI/jNlPEmyREDVqbNb1ANADEJzc5CFwQQRwb5IQDdb2jVxdui0xTLgEXwd7UWuUQ
UFipI86hXp4+0i7YP/CWiqd0ci1/+UqEbqmVGjbGzjFw06npTrrpqSQzr+QLmg/+dDGGaYqAGZr1
0zOAIM7yZtO2k+pKJuV4k0aXPlGPhcRh6VWO47mL1iinBcFhPbJC2RZfOF90vE0ThJUIoozoVeDM
DK21BuJycWHak4pKeP77etB09tsBADs/b52VkyA/UEQLaO0B3/grdg+KcEPgjAdUpTmqbOabpnkv
A49rRpl31Ef1zmwYq0HlDiatMkO8wuSjk2rAmJmSmmcMJhKuEFaPCTbzen/pu4acssMvGLtAZ5cK
kPIPg1b276Oc85wvCbo5leidrhmzbC+IwiZhPRiKXunDOg6zbvLJJadnPACCd8jl7MHS1DJEYPME
hQF9c2Wx4YkVADCOqnCwN6tH3tZXeWN39noQANjSf5MgV9NwQ9M4s9cy3oszY0/9mcdAMKBRW/ah
OJ6gBkSIlxuUbfEBhY2ls9udMbmCroAShibKo/eHG/uVNADNmXsoZtRn159gSA5ScOS5mw9v/2in
3iXYkLdKpP+4cfSbTQ6FdV13Z2T1BcUlP5taBSFChnXt2EIjZfekh53rDQp+1Bn1Tk9YbnyoFb5C
XIlK5zjsFfG6uRUInEK9OMch/J9bmmHxeKsz740KDtip7KGwmU2Y5TFYOm50vkw4CAXZ1C4PStW+
Fc9hbcTh7JCXHX18WxROZiUDmMIxSvwza7qpHcp1BZPovAGQjAHBtdoqiq0gm2UrMP+Ih/n/eoeg
/rkzNYjNo7Oz9Fztv403+nxdNjJcPGW1BAJP9/OrN6U8QATBPTWy3nAzyK8kUszXQDWJ+sEtKB80
rafALNYJsQCZgOdMCt9EL2e7G8yB42jv9pRNI/ShUQvCpHUFrNjkcvUis1QHilKwDWYbasCxB5YD
cRdz8ejbea6b9oSn85df5SoHdsUNUKHAHx+iTydY2qB+BErGXMGe0MysOKqrTYtwyx1ExnSGfz4H
OkhApw1RpQuTIckO8cZKehB5B0Ze7CGqXHGvM1xSV2mxIUn40ZcaJc06HsPW4PU7DCYAFp6Hxg+G
xRWji+C6UvNNSck5uvOu8TP1UCGbJP2J0LEzzOT9Xgrt/9rXbSfmPRsu1SsHL5Y0NkDxXWGw+dX5
uS7m+T+Ckkz9z1DaGaj/LFPHZOl1Y41pyeRsmXDpzCzmiNXPSXmknP1IakXlBTQpAVA9r8YBtrlB
fs5Kdmo42Ae/IYffl/EyBcDp1R1ZtJWgFFj6lSi8O86t2o8AI2S3G8EKVVq5MzIfL+prxcWYWVis
170QBNk0qoo2Lk/0Uk4MDxQBWsGEoitvFQVseXd5tTVK/od8XQTIU+mX7gPwp8o/SfsYwMQ/BfEc
WtQC/xYp/OebU3fjA7PHkVxOdAhYySjMp/bqLmseS+mxeyKrdPVWVoyPQ8iuQJjD7H6iDpdNFHRn
otR9ng/wKBi1lSzkuaQ5Qs4h9uNRtU3212/BLJKM0Rz/WHcoNw9gheVA2PmV4wPsMYk11c4WY34Z
VsKArKwnguBVd2Y5dKC5154FlvNRNOzcKE/FgtqST6RrDzenaAmzYqbNGNwzc2rlQZ2hV6TgNhZt
rMseF86NSJxVxNPNpdWgGEhdluP3+ojcKv2BQMsUgqBWqyl3Z1RG02ay35k88CEjj2wwgnO/cnco
Fw6nu5P2bRM4QU3GcC/wmyYZYLRIGwvy4jv2pJb2+SmCNlUVdgfy6B6mGiqj3GGawiTeU1/h4KU9
/TGvKEHeQio36emZ6ED1wfI8sLFBwCMmnUWNRGUZz0r3N0q7q5nYmM+X/WENG52wVSONniKfTxTG
LWoszVvYYpuXL1xdZqvBgQMFM2hvKGIJtIWowZWJBCJdk1WUUqxbKP5mHbOYx8TJtwzNY2go1ncD
QM0mLWKHQxm364OIhBxpEKuuMOK1SRwXA9ELkosixoxuSz2tPyjjlIr95fq/XJIuRGD4o4SZKCSm
9d4BCalwsVC9oMFxDaJ7gHSbQvRSYgLRiSfEfdBU5psI4y5Z1h4gT8VylYAKOfCpzmawwmAQkyXR
c1YdEtnba/cWFDBwqatj/wh1cqKfHSiGyeSbFeFS+lQ/NkU509dPhr2/3dwYaroipeQnxnOS5jCn
Y41UDRshQ6L7jARmBd5JwXkelKlrjbEmP1tiBAbnLVhzlrbe4SqfckdjPWHtWScq8GKokp7Waupk
FQQvArslxWUBxJSYg3e5w6ySZz/3lfKXZridaeHINV1I+4ka+leAbBXo/4B1AzLmIxnhMhfYVkXo
s1e7tU7dWhTlZtwUa+4nXWhs2gyaklgFDXO391y8ZlyzmGVlnyDHzGZR5cd167Z0p6o4idaRkn+N
a1iAh16NyjMua2qrvRNH2Bqnpp/Gq2ur8KoxEz6DGZJbrxr9N2Qg8Tvw3ogpn5yPPSHJaLzdQ8S5
Oqpd7o5SUldrRfPuSSsiO5YtfRKc2Y8G/7JFg2WAo3gpg0Q5b+5H0BOu9vxZMaKD7+hlUjjMDo9q
22OnMii1SMUqlPmQxGlfyS3YFc4IkFbXyJDOb5WgTXsIQjQ8zAaoo9tIZzgGDCz0ojkhPpXCjuUt
aiKONFRdnph5kpyaOYNiKCAk61rV5zFBA+iG87nmypnT6PNdMbAHTlJIJ46W0ZjoL2lJs4+/ylqL
1xVA+9B17U++ucCDSR948Fqnk7vxm8eno1m3e2P6xV6z1r30eltVD0U4HJeyzqexG1BjOqkorPLT
B044RS1RJfXLmwK8HyqStJXw5Jdn4d00Y2kQaJ1XNjmApZ2Nwf6cnpsrJHQbqHMyzluYaK4wtTJ9
2A9JFKh49F5h7Jx8Dylk8CB95QuaiIHV9YgCt4fl5j/I4tCU6ZicYoEJAoVYdp2ezxvHaY2HDzuW
U8EvSYyDhOEnb9GU/9W3cAhbLyyZRDG2bAveWygMvFZWC8viWlzsVTF8V9/bEjFKicXXObcfLnlh
64gZMP10mjQUNOPAMzjE0uc/PlsikfvOifruJE1yt75QbDUSVlB3mGTsj/XUqP2NPGDPa5vOB8aI
wXQr8+A2Pg4+QeM37/KP69bXm3Hmlr52qwa0DhaDnFTyOwjALdtEuPsTO9AbQGGmrZUo0ElusI5o
tHIC+2zzhRZiJKNHej1ZJsqtFhIwcuYwHREgCVIydDfEUKvlv+ZhDpGcmkF1MM+jAIx2IzcZGTLE
mhgwxYFDbLX9SUL1kjJZMK5rlzHu/35QDkVB9MyDJL4RI5C2qvu1j9KcfcaI8VVzQ6BLSNQrNsYT
/wyF6JhA5iSkNfFJFNypCkJFMLFUCHLBcHTEzA8lT0U/ow8lBqccIchkq0NlZ6CQmVbhSXV8ImsB
7U8bDS3QGpdTZfAT1zSDYsrDv5DYo86PCaE9mNVOvz8O7lw4BRAk7kV1eGgcBe0XLkZnaNP2A+JM
wLHL9Z+enEnuNRVhmfwfuM+4BD7M2+lFWiIEy0XRUEaT5LNkNrDBetJSUUk6fhi+X+AT9m8DSCvN
ZWzMC13qguad+CzFf9SAsLvATZ95Hk6qlu3e37f0iGvNNCi8MfWx8xPB1toqR7wQRubTVR3HdapZ
/mEN69A89iUaYojB6aDDCTwnAGFgf4iNx+3sI0TOWwc+m5VAohSmOMCGMl9k3FHSEc/HZ/lpZlb7
u4fmC9JUoWZci8n7Xj6hNAQhbkGWEWag1dcgDNM4ZQ4oi77c+t5bwZHiT2HPYGeqZTd4GaLWccI3
XbBavO4Dj7tLoa1PTMe+E5Rf3gvs5bttnu79ZJehcsuchX+Qx9Po86F9BKoBIeQeqhAQuH/TvzCw
xyhyRuouLLngMWarXK3UN+nS2FeP+VkT+fKFNIBqHSPCAXx/CrDHHLsj7lGTs1mtCSP3TnW5eW4L
+nTamtJEcS9rX6URtnM3IbuLIIr6rJtlOxWCpYRRRJ3woCCYAoOMDbMxWSdV+bGykW+unriAoUN8
gwlA9p6w4neonlEoMTEgE/6B4qt/hLAJbSzorWfJA5EnSirp2z4KJNEbXT074YxJ6EGUSMhjUfGZ
NVfX1ez4TUaxxgGu5veIl0Z7+/DVQN/YiUbCh0JAfbvWUOOvpXeb3bZkP+5v6mcGuEHR4TFdVN2r
5NHfuYLCnJYu/62PMnDSEzkGn76BwmUd4eFPt2I16+NtJf3cEECwI9Bj/qJRPf4AVdzii5nFZ+OE
tj3D75KlZ6BzQsbwW+Wf9CK5qUC1KkicTHSNM08q2LaoQPVOdMi5Z/oW0z20+HKPZict3kSu+e/J
vBXEvq+oPS8AMphxgQsWWz4iyGKrkyww6metWKVq1LdjL3BtapaVRT3XKzWPFjd9XyTbnZO7GCvr
UjIZkh5mBRRzR3Vt/EJk1UX96HUJGniTNjT9kPzvISaAV710M0t3Bcdgcl3Jq9hr6HUmDkjDQrCJ
I2IujpY9ojddzloGirXcSxPNUmvo2uJRSTd6DEqw32EZPChQdCqE/SpJwdSNKnB3ENgfaRjW/45S
CWj/dPBWtmuORp8wYFiQR5qINnxfewHQ4XROcn4HRbBOvZU0CetzGiWN1buOaaZnAwozdQBX/tPG
Xz6pokC7GDRAdZ3ACP56rOAAT/m4EO8W0uDPkRV0pMyf5bSX2M1oiQ2174cmGF478SjglxlPvOOm
sYb5nniFGNW6gCd6M75YMT2GjPvUuKAVyXtThDhi3f+w8huIubxhzG5GnKmE7/3WsrueKuke8OxV
eLkvPXCMppPhFg9KrtFYd8p95kzwwgoRPn3e+ZmoCSl03llTdHQA0EYSZWqv+PDXq9sRM71hTIUh
MTx4HTi6Rn2WZEyMNYtXwoZQV091IjRQeo+JdMR/j5Z6ZVNdZ+sGOCM3KLlUvXDste9dUal42jVG
9agX4kLhTmiW4TlG4jhdRq4nQqCHWk3JGJCwXYL+JRmKS4SQ1wZcu0aCNzd3fo3IW5jRnJuUKnyb
0Oilf+CCFMLMbJFjxhK2toLX0fCgSHm7WD1wbEclYgngMfoWSvOKxlVcj++qNsH7bjYy1/e19Kb+
4iSqMB21nmrM2aa7hrmwBON9r4YVG04Rv2KZQqIOOCFYK7hxQ+7RXOBRun5WKLy9DFdTENZfpeiY
hCvbYnUifDZRq2wotB43x0FYUBjVtMm3+VXprlgIdBhTquMbR/IKmz3OtLFGPMA/SiVvrT1gjsQj
0bEYjNhAU3ebkAhgLs0hVvHZkCuU6pNwrHiIat01IuwgkLCwFB+XkfeX0SrFwun5y3QM1S0ZK5l9
9Os+7CZpO7oi98/M1tJtut7Rpr+vcM5iDIo8g8QvFn1otTIv8955eX9335IgxRCa1v7RTWwWbioI
a4CIsxt1SwSmOmrT4iyYcVuA0dzBhbI2Gn+FunD/YkwvZK98I9uuMr5Boj5wzF8CMKUsLZVdBHe3
YxW3QdQpRo7+pY11qia6TiIWSS34BpDrQyi/Z7V0O+bKLm7ckzjfo1VnKsUwEme9zWNUKQdNdnB/
NhznZitVT5bIE84io1nPOtuWaG0FJNByS1nDJq3zzyNmZpQSQNh0zza+gMZyR2WnBkpNS4s25WJa
iNbitZtTvLQuTXSu0FcIGHbxreuenAZw5G8wM9mZC/Qn/6O000c+xZdLlClbgsqJLrIuY7bYhyiD
oCQ0NFbIshRIq0kpRduDWhsXFRBCcdoIU4Qt6ny6t1U+mSrTU/bLlx79hL4xQKciagVMdl+pn76Y
nCFsZbL7g93OBV6dC1XX9gIAv+SCn5cBjNJctmEDZYZUUcjqvKL34LvST35Aem5IRT6GyHZYudtx
rlMwrjTEV2ACIC7ZAnzUwWSiqXyqm+K8j2vdYpv7qOnPB0eo0bGplgm4HR/ZC5f2Fl8jQUj49VtG
88DpqIM+qbtfpDum25ncJTD1lKlfDFnEUvfve3AQuBXhtu7u+WbHVHhZBOf16qj8BYjwsedbMr8E
A62iGVZhgc+jMi1iqO6AMuOcBAShALLaz/0+mEK1b/hJ3zEM3NsZdB3ZxJjjajsWn/QEb/906Z72
Y6oXFFiyNswYUlqQn5kai8YLyhZ8mLQlx+dUhKZWIlMzaiz8s8VaDaTVjCFVONqONDgG7bAZQvVt
C3vX+MesluNtikKmow+z4Shq0elj+ln+7/lzKARtUIX8WYyZ16pq7IDCM3VQBtmGRq250cUhKQNk
5aN6tEEyvY8lGa3bQoSkPvwIMfqSv21Sqp6WB+p+Ht8Cw8VepEHHK0nAtiPLiMPB8ntppVxpJ4+Y
8NTY7RsYKpazqTKnzFrzjIgj5adwd2FhhXMwJiCenXQaQGcgN2W5qzgxwTvmFTH/k0G+/kBGFSM8
rMRFr07GemOBbMCVg7Tyd+ZFlEsFUgcd/IowD8HmSf4uqXgQ+r4abwZiyCVyb0iv+9+buAjzlvQR
1H+qNpWQUPGOpzQh1mCABTaNcJ8wMu2rK5bcbs2ai849Aj0PQVpqY6IYxj32xx0gTm23cfK/ew95
b/17hVjvYp8iZS8OCJhjOEUg3AcmjqPCu9FK0rm5hVJ/XQTjsxPDqsHjxsbwcFiQI30YIa3vu2Hd
7Q1Bqrb8jECcQVjt7ajBVV/J7DcoQ5cCcjqLdqX+o3W/T7SEgjU+ut5vqfltC+1KVcg99RpY6qcF
JWfeUUS9RyM8DiZluxdixy9A94EFMuQZAdPc57vPn1k2uBEWmua/QOEn8oEqHyL7VJYUDzfAHkAl
NfMvKMy96l1EgQKCzrWMbNcNdQG4/lgQSZ6uCpzjgvD5QtHrzgxDoBO/wCG0da7SeDSpmv8VOBm7
Wk1eXpH6EkQBfooQU6H8LRgbGOtSubEN4eclnvrkFp0SJ5MjhMuRsjW4QuJHHgImlXpYnHCGlwwf
0J3USlh/lA4Mh1IYcNEQF8Lo7T0VjVjGmn5hFDIiW3L0f1ze6fs6U+J3XS/3evYn9nYrTbQh303c
Jy/5kfLODA8Z9X2MjuIPYU4coSGuL82WpFptPNT0rgFUhRXuPxQcRBkTiEus4nU7xYSVRO6TPs2b
XBzr3Ilcwa+euaNn6nWyuSFs/2UTnq/g6JTBrCGH2Fzj2EXkZT3DTxLA2oV0kPOH3dp5pRw+smoK
l5atu+WH8PfUveR+fXUGQOhFg85y/TBS6vZgHQqIKPWs4qGASFCs9c50kBlmSJa75qzOP/XEeW6F
tN8aMuMNYRZg9pbwE7TPNpxZCe8l8bsc2/N7DHxdae9Z4s+ZmlymJPTzD7z7F1ZXRCIwpObM6pGD
HL8rGawFA3nI9xTsr0IWi2yahKNivh989YFFJF8s/brUwC3Zt1raQ6Elmded3OVtGgtqfGRtyMna
FteP5T+h2tqNxt6/4HowT3MTS1Zoe5natM2dcD2WRe29yu+iPaHhyvS8n7jzyyf9IFK6a5bOEw5/
O6h3tvDY/D96S9Bg6oTH2ErtJHElx2rID33JyTXngHDjaNZInyNAphHsBC8TbBIYrUWOefvQRvDM
YR63HtdJon/9TKoWkiOn869Soq5uCepryBXwRbCz1snsLkgcMfVk4Tt9B7lt3ZlMRrNB5qYe61LR
V5hOSG06xdP689AGPN2RIkKsupBFjfOjNiS6xU/S9cTPvC1SJqOBxnnzuRjJivZNiX/d8DSLHgEs
JUafIdDP+NOCJXlOmCcKuuDLXqNVASAS+yk/h1yJkGQBWdYZJZv5xjv1ok2fqbbzYmpemU5T298C
2M9XRZ7750cOnOfjVK95G1HqJZS32LwlnQxVbUI6Q6E8JRhhslDyBq3fxJIwIuNadu64aL2Do0fB
I8rUgMicqYWWLDGKxPe3LR7J4d68AEzxaJT8YAbnRkcVTaxtaGEzXoc4dIJmIJ0wutV3/pA6zdcf
p+Hl4wcCvTGQ/MK9F6Kz/K74ljDicK9OeTIIGaEx1ikJZz3ycbhV9bP4j3bV3MpFH8qaBN/IvyPr
zZOT91/bZlwwvE1YvFJtAe4NzMXhj1Yyn38PyCkOhmKa7hriTqYc1oz81GZYlL5Wnd4X9i2UZvwK
Bsc8A6FgEMLz10D8o3245igv9CZui1nH+9pdJHCaD3INbkyiPd1Lhf7Jgxdg+FYCkTEo/ylAsep8
E84ZNq7zDWGUnWR9bCWm1N14muLv/YAubapW7Nu22Zx+4QMOVJCGPTnGqsa65CvLIGZkNeVHsrEw
egZUqpMT5UsjnRJXgaxZ5wnc6Dfr0sXLXU8qNxrJF1SrdcVegnWZg3NK9AUlGcoj9tO61VbMDYoZ
zX1F60Khy/koMbRpM3Vn/g3GqRI0VJ+DaRyqTh1+YX2q+Y2ajWrIuoH179tYXQxYx25fvvACZC05
vz8soaCzWTtIoDSjDvmUVCBYrwiHEa6LvJVLn5aZluKuDFVUkNnwApRzu7/W5EaSDRYFj4dIzySt
S9ZRGRWMtOInEEV4eAZIcl8Pz5h9SsZxPRQB3KMU1KlBuGZahfEuxq5h7Ug5Ps5b+wMhuuYAkzI+
UKs0k+nmFu9eaCGro3+Gz77C7K/ICZwvBzNAU3/tVfKMgqr2+26V8QPOOJXn6I7VPaHLfLvNA+3G
bb4mB9LjVta9oPrXlqwAseTeOEnlEwDzSOMJ77Z1ZXbwi1oMx3Knpk7KxEPAQ2i9eLDLXFo9Wga3
o2J+mZENY9zU40KgpLEYfnF4Lp5R5661RokDWA5GYde+yeA/DOpu6YpSlQhGYMzZOCOYuQ00nMAF
oBaDQNvYlDg8NvA7oR1VjmOgYvlAf4MyInuujXiS14uhRELKS6TFEp8jgiBfE97ist3OH92efLLz
Cf5P9JlgM9+KZ4M4+nSA8MSXv3S6P3eDv2zgHJ4QCs0lJNPQc8i4zv9sHQzIUhKl1fXSbj+3LVq1
Bi37YqWkNXxA/dOZJrKZ9ikZHxDeB+SHq9xcjvZHmKe/GBEvkusvZVhMjrIKJL0wbZqljoO7OptC
PctyJ9z6JTfOoYwPM0W5dH87S1GW2ps5ZFmMZvemToQPmvWvO4eDt09OO7/SXME4ji7+ASgX+GhI
RhWM3gPTcP+zD9YfYoA+qaTye6swJII4/e3h99Di93s97Sqk2yMv0truWjJfes8YgY13EAViNVFa
xLFTF8XW5feQnCz7mQaBVf8YQtHtwLf9aQEOE0Obrlxvq2LnB/defURgdQ7f39YPeVlYZ+U3yjmW
gkUwK/qkgNl5QGY91qc0aRkLyBc6A1v8Yj9vyk1TP9GElDX21bvSv+0JtocaIHRgBoyc0oN+CTR7
HWmS9QMUx4V+mXmBbE24tU2RwD7xr4wR00ThDkk5QwLkTqS3WUx+Pt0Xaez/w1ogYFT0dlqC/zn7
0zBKaWfYFj1pb/ZZENzfWCI5kR/XbZ+j3Yz8bVTa4GIctbBs4VkzcY6YPCvSH7ht5NzVnHAHu2H+
+GMzcf0FxdKY+csgeO/DEyr/LpUZ92SIv9HyzHMuO1kJSLMj+Vx7SHmOJKb8j9TWrkKeoRXytqOJ
Mux8AZ0x2Aktw+p6M2HJNYTD+i/X9qfXwmuoXtm/ezm9yor2asgM7iVeHJcLqTJsGCqI8OZDUnkm
EjbfI9u6fprx7ECvX4qy2ZDc1gQSRZ1fnvkF4qVwCGPqcgrZ8BLd5o4NzuEHsGR6SJe/QjV4pP6N
MabYfrHgndmjaeM8EiGIao6RFrid6FJnwlxIx6bVfC5buYXBJFb+8Hk0uS+yKbpDSTkkHjReCM+h
YhqXms+KBSX24Z4d1sRo6p1OevO2BODO7MpUNb2ObwF6F9IpaPV/nDnencAUOO6stnn546Y/mxMj
g6YCZf84ehuyLNwGiwqI9v1ZD1EhtphAeo0IJrIk+kKHESUimpNl3RUjQOdqhQTwSH0AhHL/yPPv
zFhHBJtMacNRU8sOXgSU+9PpcLPVUFalb5l8hQlpRCSl6OfMuvkIciWOD0SZ0ilraFy2NsVb0T7N
lVCwu3PCDDH/PlPOvCxdreGPsdZ3TJ1IICp3cNfJOYYy2a1e9Ux5P1+ZO9ta8qiWhuITf1pV5QPs
Pe66AJtRO513XG6kCJBWAfiP4oI6i3kICAPnsLubaBwbKPqsDQHVoryRAylsCeXahk63WGUsrz8s
0osqJUY9/0MbDoPfRyKZCqH7iLWduuzfAvY91RJAPH2z77od09cHxXWD9rvQp7sMAq9iBr886C+L
XNtPau+aAADopd8TkxxC+lpBuwF2UjZmvLaRo976e8qBF1xgDQbxzYYhjsidHWnEtIlzkaz7O2j8
WSkJaDMJFQq6hvo7fh88irboYqYbKcAP0KseCWNAk6mPJKu3fOEkTTaUuVbyTwG15GvknGB7ZFFd
FtfVoARsp5XC5r2xR17ULfMLnGWmi0YJeYNvFpqp85DY2k30eGO4C/R1ilAhAgceq9dfktpDTN08
IrSnJgpx5uA9rJRa5Vmo6cj8tK3bEJkXx8VBJGArGskkfNF60RGE23sWMOUqBrpBpWg6AH3eokXk
up467Smycr8krmJ79WU5mqeaJkDEBzl9MbWGTdWOQSkbhH+xKhtfIerHyR+a2bjvyyUtm4vhemwy
U8VlQBP9H2b+j6xPytrAJKkFPYbbx+rVRY8/IJ+VPA3rXEFh9qLnspq17x+rt9299NW04OrGF1OI
XQJm4VIcewAi1z7UrjipuKw5Ad4WLTQDl6BW8KLHFe4tEjmNYihM15x+980LAPyEWQbd3mBjBcMr
Fjva7JsfeLxmk6F1wo8KiMpfQ7u7kyETOgDkMpez1UfItM3Oo8HniJ34xy/xqlmL9wXCHep68oLg
+8UGJlteF2rEDfXy6zvbIDkb+0hIqZHyQVjcBBetFW8aRlol5sbM1O55AmdT5XXT6iKhpSHMR0rZ
8KSEi0i7OWWnQsPBDxbkBjbOefB8Hy5J6rkbmJgnTAjmdX65fydGIKpxbEX7VuSNK0JYz4HqtMT8
O7VfIvfzKQJ86MWmpcK2UaG5V2dp5zMuthvNHfs9nS7qGsxEv6lA+qhjXGMrkj1d73HWaUYtCUnJ
Z3GDrTzQqRoEErRAaWMYy7+aoEf4NlYzhHJHuzLLXzi40F4GboRBWYt52Mpf0tkS3qIFMHqqlddy
Ek2WzM4UO8xL3dc+U2wKpLMMzXEDDmAHmSuQHzBd9oLjumJ2kmXU3VdUxcBio9aSHE74xloL9lIl
KW9/vH6rlbE+8TzmXpGVj0aKSDmR8HVHpNyBnbvIB2mOopnhmO4OgIg9TREvLBJws4zB9kf0HkqA
cOAa6QZriafJik/cXG3DR7Oy2zfFKUSmdq/vHgAPCRoqRxYirjzsV6SQ60zwJyHZe1C0JeiGhdvH
k7O4fHKQe6BrdPLmJozqxdLdB4ODA07mZbrVMbUUiLbFSdHiWzYY/JN/MqVvsIKhkcW3Bg7OOrre
8fEj/RQoQD0ISJ5p2tNmxouN8FC+4VJjv++4vpE/t+0rINzyNEeeIWOHCsjxWACxL930vmtl8xxe
TmiNq0mcy31sDaLBfWDOFw8o9WnVBj+rxZnmo1RsUcEodPwheFCnugj2Cjbvw4GKPWH0IAP7S8GR
LOf27/RQx+gC/nsmdr/n1PTYIddtY1KFn6F7aMCo7D4uU/KYZxb/vxypbBHujgS5S+rRk/yYjAD5
vknN6CO/7SsXjVE9YBMnMkaeEt6uzbVpjlnJ/QvNhdIW0LSRAv/Ccu+/hfaguK8fDO1eRR9Pk3XJ
oIqgHRuceCGglT6XY11XoQVioUKrZE3ziJE/IQI0GeETBIhRs0uiAsAgMWXK+HOKaeGp4HQc9Mh1
93Xnjlmv8+h7BLHSEdqPGSCyMGsMxhZQsF4cyHPzJ9HvwrQOydLIpqe8DRg0BmF8BrVUHcNFCGgH
kP216R+2xERRW7ovd62EFd7OHQOsxylbjOPfZvi1bK8qWeUfi/XWyCpQvCgSwrM8MUCVK7Pidltv
GB1c8U2K3n2PAL+AaFu3/Oj69TYPTmnP/2/A5E54UCCuxuTFhBSI6unWqQykHGe6KuQR/d13rgaO
ise+eQ/N7KkP73ZIgJHtGSaXMKTf0ZO9sto/xy2sQmCZBDgGhlOk8HKTwYsWb10UVQn25tER+9dN
/B/fOneuGJo8QHQ0C7zNf3NZ993hXsbnTuvjx60DpDbnHkSP4Yn/H1WiA3k5Ubn7ruNoJyCQvSZk
7GsAcLm6Rr7o3YVYLRY+g+5JJrGmpsnCluLTa+zPVve6ySv/40TLDRwmm33AIpT5tSDCT3aexnGx
z6rL96LhIuV6RlQe0+boxTaSugfpbatf/iKQb1erA5tgvBjAOVccgc4Vx8aNZyW5Z4wFDtCcSULq
WAB35dd7Xi/5CJJLsaa/if9aG8pAMr38JB8E+vtdRQsRvE5ybsQrehVpeDCyIIcEvb3tFQjys2M/
I5YOapAXCvlvSfOlZztyxYXOqs6cl5Gnxo6pACUCePWA6ukg+cvvV8bXr1hIw3nOhVxASbJhHCbx
2DPQr6tsrM6H5hiM//rZvq7jvkg0xix5m0vRyftSGICMm/byOK903fKkFLXZt2oMv96SssVdZ2nK
L/zdzIrt6OgTrcILk7FwdOtOGOb+sbEPuWJAXp3/FllBWa6hV8mWJE/4PyaQtME2K6wur8bob6Js
E3vUb+q6e27UQqU8Qa4+bOQXy7/EPPvyj0ORHHyWlMFDC2+A0ho0AYmz5fdXg55Mx0JhlcQ+Ztv9
g7mTrXKLilKLzBSfRQwqBJC8uAH6QubvTaQsV/aVFccNdBbaf32kLbYLG/NVGGU6LsDKLJ9A30a5
9qvA5TPv61bt7Y/DnjiZRm6dp1ENMtw0CH4jK85mJv5F/uzjwDqsrgIbeD5IHTNLh/jQ7MExoMhI
yxOTDiNJPtv5mDCv+dPunz/MOylPPL3UBI7rgKFpqpGAi5M+spBnQWdh9JpFFHXyHW2R0qbVp6s5
tooH8NCSRDopCg/kHaJmm5Kojt8xTl9pg57r4tIQLItqag3JaqLF36HSTxZJc2HIVh7LkQeYn1EK
3F1632hjjQpsgrYSma6Kv/JBroCQwJMolI7b1nEJZZNlvPkFv4D1Mj7leTfv41cO163R5PNbObes
h4DvhAyiHmbS6NpPydD+e1UOeNlNkIHdpz+/ym3+MaxYu2XZ7lfeX+Hk56/EfH6jpR5Udkf24ara
rUGI18a4PvYhXbWtH1X6+vUdSUdLfWyts279o2v/sqX2blLgAxnrV7jG3o/nJOzZTM4D/pIWUkfi
v2uCCefk20fx60Kea5heXGqH78LQD0rurz6kMO6hg1OGK4c4OK9cHOWDvgOTXtXtiAcN0TE43Fvw
B3e3+xGkTla2UMqhT6r+3MYNTbiSf+qryTTMthgrl/StB0TGxbqYuZEdk1lxy3b2nJefKHPLlWhR
eCMLMrVm05SWBh40gi9DPeYI56gWAf7AAiTpb1bj0WByEpCADy+mWk6kNzQU2t9W6kKL9Z88DJZc
CcF2KGuSc1l3btbV/JwO3JVrSUcF/xX1ilvg9+5RCNJfD1KQK8bjs5SLfnheOyKiOG1giuvhNp6e
TbLpDfIj37HFbGLMUp1zn6Gsgwd/+yHp8Yf1eDN+8i+QIVo0BUfULHVLJMj9dvFxjdcQmFuZwUli
gKgRoADsuwuRyQXpTwcDZBNNixxNSsMtTKFW6GxlVWQ+Qf22lQ3a0WIuIN1D7AK3JIYcAYFuZS+b
2zsQtJQX/xXSvA6UNYgWbs9jSxQQe3WBvRkUpCwa3s3WAu76z2YfET3L7DGU212DuB/7tzoRpsv2
p3AVEFjHFopQQnNRf2zBEijdGtx1PsvU4bc1A1FQqXeBahNIDNvjVcYh3PbahSQaLZUVwaxuiRXN
WWxHAx0u0K8N+6FJEp4fELUGWGdP5eszXGBpYnnfz1em+lDxz69AqjpKaXSJU5bFpVs8/fL03TC8
MHlKYzmM5bvATTeRKvY0b/7ZV/gHUA5QecrQJDaszgD+meSI2rE863kWWxr5QSssVqea3owLHHnQ
OafaRScli4UjvvsWlsasv7pEOWWjsnb9UWMjPX8zUMJFwJUddzKYkoY2XHtqXmfxNK5N+oyzATJq
ZyobzLeM6hgp+NsKY8DBFwiHZ0G43kBQFPdVguz3Hfm61ywl0j9jo27oXimzRjO5inBYpnKqU00M
omUVdJBbs5NIpLp7Fph7QedBE+3xERmP4AEyCpV/4PAj6vloEvq3UuWxafLf24bfeGVAhDC87kwq
msUygdOUDWXyEczpBais9Ghhh5KAhebNAuAQ0Qsl/TXo21FgEhBkYryct96odIQ2Y7lzbHuHo5cs
o5z9H3NaBMM8AyJ/oNPwLXfttbEaoI05mcWO0YE214I3gB7DkqkhRrpYIAiWSnVafMzrpkbeZ+Pl
FAdijAPGW0QFxNEAcckDvjBN3euvm8e9v95CRtj3uxUam+P5cZo/vmIsh+zZ6tMK69NA2R/x7NHm
hODzzRLUiG/oOv840yN23XGp/GcwMAoXV2jKO9tz7g8mZwvX65b8lRM0PoLsX2V06DSt2G1Bgwvv
Kxgnvlz2V65Se7iCwXyctgm24xVkJWPr67AN0Rrz2ASv9SH0VRQEXDLo70rKrY2KV9P5MtAegD7S
KhkTPQECQZUPdS1rnJtUz1dPeNmGnpMlP3y+6s055w2HkeYd5t1k2BLRT7Lth5mxfnmoSkHd9V+m
waJUnVsPRDQy07xXnZ5d/9GjabRKWmdDCRZ15nVQvlJfoAVZhe7RSXZ8EWDYKflBWf0GQpP1Xye/
X24Ham/+b8qucv3WgQoZTwf9HSNA3O0HDIkNBjZWR9NoQuzO01gIxAH4qFt6u7hRm3kJjyF3Vv7R
RTZXeRQzqzDoPSGrOcLfiFn+SwQBiAYdh5zgZv5KZJ0I4ESZtFypOHNoC25q6nc9gOuLZlJaVuzB
lHsWEqXqUBqTFc7iNl7yyWV0uj/3/kqKr61+v/fB0Od9RSeOB+Y1PK6wfprxhxdUy+k+z5UGfh+A
OEvNZigC5ERCr6OuXqKIGftZA4PVsCLcwusjpapCnzHm1KsXFpr9sAr3mvRj2Ckkr3b3f0ELlNYu
BrXHeheIMxOQHJ1NrzneoIAjfqOazcvk8h6Z0ER0JktHSwznrXWcBytCnCrQCgHqS15RFn40k7Ts
VS23/s4Z2C1p35+HkFH9vzwB1pdgiPaOb2A4tgEH0eXer9ReAEXdvCdLKPL4izZae9QVdFMjo0/j
dyso4RAEG7TAyFtmqXGGRZDyitZYDErK3BlL8sYWLlnzC6dPIP81jC74IkXY2LSwTX8d5QkP3L43
5rSbETziXid5bSC/0D32oaPh1Owy2Q7VihmOBMhGXiXz+hirqR/BtEWL3RtsrmrwmYqIvnDBIk4D
kHrA9/Ch06+8Ac8saQMXXx1xoiZnsgpYD7rFpWPLCokJIG3on6s2dvoxRN9aBXZpEefuKY4Qexe0
Q+cugVjLytKfEA2OsI580Hf/YRbP8xIOVsnyuLMZ4AJgZjDu5J2iSuX585aAt1yvPrrH//XxxeW4
fhCjpfucWGc9Mkv0dJYwQhopxvXFVWqlsaBVeoa+Q+egjjOYTVviofjjJaHouwjUu368UwkKJo5P
xIkaQTxsSq628QiPW2Bgjg5Kr8GLuhFkS7KnHWHn8DbKXQb9Od5tW4WzN95DS7PxKuJiYjp6QIGV
RNEETaYFZDvqKEQ3sgQe90oJQqO8qrMeusSF0oSC2/wwC3VMQsX2ZUmiNzDGMVzrtFaGgKHQ2o2O
DbzOOA7bu7pd9MYQXR1XVwC7laMSi0DFcnQyf7isJSpldBBNCAQAAMQ6DAwEtL9f/+KouVcafVxm
XcxjOwwkd7fAiS8cEHMOP9gh+yF/lU9X9IGAYwF2fRobUhwLPZiKNFi/yRdbLw/e6u8sU/UlhWtP
EmKSD+kJNyA4gJ4R6YBdFdzXsglXncb/L3Ce6+jPhcYhOF3NpVoLHfV0zHWVI9T6O3Q/TWK/Xt6j
m7npVxxhSsGhoPJm0H6VgEeEl3C84jE9bzNHegn2NSK33/6jodRGbLnQVBTolChhmCQ2yN2tAjtY
2zANDK6JXs/kPvItFXZ0txQjxtuOE1GXJIlZQicMOXFeIN0bo3DOEf/80Kicfs3RZTEr0X67WQtI
dXe/5fl4t9Qoyo5XpV4gIcFics87U76zJFBxPue7fb0GBTU15dX75bxJhQz5C60EoGDGz0AVcp+M
XZff9aAHmV4sJRJ9KgFSmYbGv63RE+g9cQh5dy6svme1iDrhmMDJpZsPuNbTlLy9xia03LB8oBlT
w3urqfsO4ZWTw6VhNVOfdchsPigHAzPr1LYEwV3APg8TT/h9le/we2vaLwG6ISJS3veYPYWKeSm+
t3Ka3cJ26FKitG2ubI/uWyzJF3n/Fqyb/hiG7ufFFZC5s6stlLARsujXoRZPS8R2tCUz8iHsevRR
7xdU8Ei6Czf4KcVN7NvJsycS6wp4/aUf4FN2t7CEjLsMdd+eUDvX/T1js26QtDmT2Wf07ycMPpYq
JEJaZVuVVhMEIJvkdvHdsl5uchoQoJhWo41/IKty7JU6Qw4JyQrgd417ce4QTJENQEjIIjTKQIzz
UcMzHbK9LmeubZar4nGYagouncFsk9eX0WffemaA92UGw5lT6aR6uStu5m5zjmauL3jtSs9n8w0B
GPIPqQHgvBMtuRX6ig3zCvwBRn5GlvP10/Zcq/+apEUMRxV0sskYmPDd3eJJ+Ve4lU9K5YC6ume6
ZfbEXBQaNNfp4UZBFw6n63GF1J2KwaYaVUBFh8O1VM6UFkubQpc60r/JRPxCceiXkLIcJcnViMll
QLAS9XhAXtYp2XIGUiknXp+Ic4HdupZt/u7qGPUZZLxjdlnh7eQaxf8aVbMLUuvWTZL3kYkB+hgV
GnvkHXb98UwieDAjHa308UzQs8LPS4IUieXwwNGzuoDqpojAu/LTljJglBfkq83C/qRS9HUt26Jk
ZXptkbM7HrFawu6E66/wcj5rLwlwWBVbpjT+7jP0GSYHIDI+e35tbyHsWBvRFHrTJdEwC2ldB+M9
e6kwQ0vlo0PcCRXF5m2pzrLFNsg2fU6wTHJWmLESG4dPYC31Qwpkv4dh6/yJrMuAFhyyyxP5WT94
YE6JQpDtaUiJye7eMnpmDMSbXdl1W1uqZpnOr6erTWq3ZXcy3+PzQa1eo5C9qKgr1pVb8yuE+5Vq
LZJradYPzJ5oNWw5fCaWpdL8Fsz9KngSRaC8Ms0lh/pdcaL07laJhaktMvn6IXsilwi9G5GmC2r8
ErZdvp1OSYXsnPbkswOxC6Dj1oOSfHVyRp1S0v9unJbIFwSk6sY4tlqcUCqM1+ET8xep6jaR6J9k
qs9ravkdBVGydM69r0d1Zro3RrPusAq6D5HtyffVZNd6SRRk5uUAocmVthM2/eVRMiSQM4FGgPUD
NTy/59uGvwEOZb5akCvZqHkgQGBn9UAPz300wCxo3xs9yAiy4zTAmPcVldEdqmIGgmAWWJsESHWy
OqvBAWSLby7cPtnwrXAVKyhLRRhT0jN0t7oFF9vIvlCDFLR0zUr5rXNpB5AIzMNH41jStxcH9o3q
wuOnN7dZnSxxDItfGELmCniY2mYKFl3EY1ZNuZVmxTvmhZb4vYimAvB12qhAczflm62lajilxhJX
VP94CN6Kc94o9C9skiMprJoUsmV438WTZ1V3OmVundIIyOshJjURF5a7Mu0j2n3y2TPL00BWbjyZ
tI5JstVTZ4tUUfYlWLE8PitxOQhrxotKTY/+GVyOnpCy2aStPCjUHzfqwWxJJCbvJg11mb2aO1Vu
HfXjJCmI6AEJPFhRVfn2wn/100NV2pQLur1tB1P52vct3Hsn7z0796Ah2jaGkTqsGmMYCgE6Q7E9
xqLEj7Y3YzU1tnKlniXa3eOV4B8TtLx5YBBzYEYBZRUe6EjAiKy6aUzui78zarqaXIOJbN2P+gGG
gmvH/KfFnW/XR7J6dvjVhuayRvfTBYBXQnQddDnMNDdTMbGcZOD3dbgBxa41g4X4wsPZ1coA+H/e
e0zp9EEqtEEBnQmek+U+qFSQxPIJ2ur7zZWjzLUXhbtM4En6h4ZW7SDRlv5ph9ZrfQ99Ve01YqLL
3KS9DLtSyGzNl5ugfpVWywswfWuMl6vjjfV3EzBXqrt+ency3NJe6YyavZ/Ni+rz9xDeQr1mW11C
THvPeXkOtroXwBgJylHBvwmB/mZvr4YU/4EE1yJMWcRRnlJml/89ogny/Nf7yTHSGDBNIBsps769
UVYR7iOk3ds5R7Y1esUCkjfAK4g55U/MNRVgh9OQtn8sAPTms30sS/r1AbnINaDMyHgCKnyxrBwC
LWQfxjE/XH7h1bYGtLWu02pYJO6jHNwWfY0+8HjZDAHIh83kliaMfF98drgrk9m2E7SdmIpRkjA4
5nXKEFw7hLiyytsCwyaMWa9U1on6eOktk71OyxPvheMeFdUFVweHf7JsQgskq+kFan5hhCLcytTp
v2kcXxVvwkX/zrqYqr8mYY3smGxuP4HGm8YuIS+aJbKMEjUrrlnVmqOTlq1bxn+V5X1e+bCzwZ/C
cobbiSqh88ZTKd8s1YzdhANkGdOoa3yiQKevZt5dYmDnZ4SlIYPbLCt79HgcbjJVck3L8f29NShh
O69NHUEEWWY2bCV7YJ/aX3l7aS4TggJyAFEANdGHnwdeABBimkTKI2MYsEAu6Su6mZcDtnZ4n/yT
alrS0orRkzmLhwTjixy3SFOjeflqaxvmN6iI2p6uzzwUYU6tF0ez8Ls6lAqj8k/AhWvLMh3tlE52
e0+7E9Qh6vP8Ob20NWqSGYdJ59mv4lSo30LBdd/0fPZJebBfEsloWUuUAvWJmm6UsmuC8M4mrM/C
HOX4eRDzvjL6p/tieD5+foeDYMQXnJCvg+8M2vIuuqZv6XqDmGRqYGB1V43eEyQaJt9NNdDrRzbN
fDZ4Ydhkmfecjr+yNPZ4Zdx2cmdpcQF+n3hH9IhAYNjN6APZyzYocqWNZaESdhvH3PrdmE311Mum
PrZnT5mlPfiXDrF70+wOUkozWMCT5w9b7I1ZTp5cKFamDDyAMFJwxuEAeOKeaOHEs51Hflky6BBG
zOtnBVpThkFa+hyVaO5qrGa5HiFtp5QTkvPr3XTrv30IMEqTn4DT3gBMap36ZBogXtBCQ1dYcoRv
wTXmZOzNrrnHjoCodi/fFCLKfC571k5QiLmvIrXMmHvZrRs4PjMcKjQeWFShFlT3SpXhCzxB4PKw
fBs0SyXPUedbmTxdZzWvAjHPimooduPHva4KDW/xsjPrzHGMxPQrdm5i6+LCUOsF5le+or0bFAPf
ohsprteJvxrxxFVRwKvp2ft0sVXc9M+K5XIO29mPqVua4LY00u1j6FiYcM6YbVpL6V58X25vKS+O
BOWXuk0XhXzz4lMB+lzfAI3FB2583cyPt0/dou8DYvsZ+1ZPGQNXj8RaUdoO/uBBEKk1WCDkAsCw
9G7xnMDyx1r4mHI9Dg+6vDELPJnwsEm3HRtGQ9AVrS7VyQh2KL6cWazMi80yPZG57neoeBfefZ2s
5w6K9exx4qZhns281Bgxm4WScYZmz4iGWASERuJn+AWp0vKcGuwqRwVmAZCWGX5g+eSIH3PEa/kO
szzN3vUekgO4mehK4VnO/RwgMsRy6SkWXXqYlFcuf5IJgPwsqZ9t4kEBRSgKCyUy56a387T1Y073
RUzrWVjdt1XqtiGzPWI2yeXjDIiDPslVcS1Bc5BYKlWbsQYJZt97Edl0j64D2hUXFMIj83G75bKl
alRFatA5BKf5HYskUU/b8NtHOkH7rdGVq1+Utn2u2PNuPmv7yqqclqqfawCxAahMjwRVLWDrp8YZ
w5bQfzQl6uJn6rjxvtbDv+BzN0D++qanKvkzKPTTxA0tmpSZ2xSpNmLssotSeLhnkWQQTCjPzxUD
CAZot6jU9jHiYSQxKFYHonUDwzrAgpixrvSetwWm5u50ct4IsTpVhLxbaIGX4K8XCtuKQohTZLJA
SFRMMREbTIOfYQtMf8sSY8r6bPE+a74BzB3z4oq8EkYZuFbhrhWw7dPX7hjDAHN7CGGveJ9ZTDF2
QlWHQptr19fWKThrErXs78PnqVHBU2aeIlO/JV/Jy859HDaI/IykD8cwbb2lk8Xn3TpD2LLHGPQP
XkO/eIWqYViNOuTOgCNRtT4rM48L+6umGhiXkSA1GKCS5R4xBFdm3NFQuiCniNO6QSq4gu2J7cKV
+dLwL0r7AL/LKNAkgxH/M6ytaURPYPm4J71rh33STfKzaehDhXqTn3Q/RC2eZgHir2fearJneD7a
eBU7fag+lpV0QPVfjGj21nnAkOijVwrPLE/4i1A8yz8s9X8dRLGIgcCzlATfj2mMFrRX1KpfJsr0
qWIoG1ZLU5N5J4gYqY5efY2tzeDOcHJmdrdCEk8MrLE+AVGMm5RyIY/wtZo5I7BWIwuFFr018WsB
9y8vx+YNfqWq7uTlq8cP1+LzXqFAoBeu92EM3L+OhQuGTk6OGG3yUsRaDY48S3JtbfPenR/FSvso
bnUH0HboYnLNNd4Cky7fXx/B5odgdpjRxnSz6j0s+Z46ssSxTzj5m0L6tuA4q5f2yM6IH0XI+nlQ
82BxRFQ4kNMDBkxwUDDMS2c1FX5PpJYB3DMgy+uS9E9NjPi3bUg283++vcDncrSIALn2QlTA01iK
tGicMhIjpQFV2VrnxLOpIDYkEtia7Op2fUIuwnADYL0qdd+yByyXTy/EkupyZlpg/YD2bUSiP3Xg
VWKBrFDYf+hLG2EjH9OwIlotrvMlUZIXSqNpVfHYWchW0xXkUvadXRW/m0JESRrBUvOxzeqcxMvQ
FzvF4LEDAt2d/fX9DsE2eWD/IUb6iufcspVmRMBGASzp7zlvup+7Lg8BQMwcuyPlWZ6RqtJDdrzp
jyJns3Ux5fo2uk+RUkfVELbEwA3Y0y6QKeP4zNB+pHhPvpIRIT2FHw8JdLlC6pTpgHHvo2S58dX4
zyWm18rP6IVjQCblsIEhJ0F/C+cbiDwlhcGtmUKIrYqbUwN/DgHqCCTMafBQlYKUMnnI+F9G5aCy
TvxEy7mLzPlY6ztcM/Px3YT1KrUije6fZ5oW1m/sUN4o1QcxCP06OlkejQEydgg5XfIcA/uE1+9W
eqqc0FMi5wPcwcftQStKRYWttcFaijLvf4MgztV+Z/D+8zU65tG+mlUS9bLZWqZolZVYpP3IYIsg
WGTFDs4f+o1ALsrJpIMt9LRrrRvtawdhOdEwlfFwOzr0BBGmuyoJdBCtcL/XoXtgqpuiglQUG3Yn
5fw915s3CtKJF7xDvHjSY41qed/B3ytGDwF3rm7AV0nLDaS0iPqE/uvR5e1nE/h7gvyU7qCv7dAi
/BX1Wv2UBGtozaoFmJMcnRQQSTUnf+dSPoe8PSeK9fxJaYkKv4xnccpk6IsTZaOL4CrehWQlNMRB
Tsh/MvFRL0CCNxjGH/G9bAYbOeSXYB9vw9SqKxG7WtYA6q9G3rgOPPIKuMF5nJh5axPZ2EgvJ8ys
Lcp8kH8CFLotraK2tS7l02GHGO+zbAdFdgZzBaMVdhgjRkyEH6/V0AsKOiS4+404+lMuCih4HUr6
UdkCpoub+ABVKLCCdP6YPX6rFZuohF2U8V/MGvpZZ2ewUqaNFbWW2zBY4gNS3dzrwVHzzy41oClx
L4+AgnkocJXZiw1MNthUndEtFcsjJmpqdHx+cQktTevWzXu8a1FCOywYpZeh9MmhkUw9b/1PS4xq
twx5/yHFsuRuk8vOU9P9mEaMV/TaGOtVy6p3kYK11xXyeaJNVplL/gOLf457pDTudVy8B7/cEnJ7
DNDEd0iW97IXTLPNiu3LL9jcuEGFrcOzrNFqgD1NyUOOnu9T6CQwyUvgsoj6VkDbqIZW99xXJkdu
muaU+NWM5MTlCvwwvczgE73UxrSFJT47qy+ZN2OkVc7exuj1vWQHYG+NKtLURVYx7zw1lgdUxf9F
w2BFaR8jlUpDBy0yxFcJqDaKsGWuiDrWdSS6S8iuuRiSLUS0ANFFazUBdfIkWQhjUQ18AT+wP8MO
B9VWTdDoYdMYwIeh1SFjZKz3BxyArdIMSo1x23NZP7xaXNbvvWG+7W4ow7vIGjxYhAzAG5cBJ849
lFfeGRZWUSp+fC9fL4LJm+rqGn08KgFABS8V0F7X2qCSK48+QVATaw96AHYqpvJFX6kjNxMXWCC0
5redF4C5LQndtIA+FsQJqUMWwvBumF0MzugOz1OCNooBLHeXxtHxA5Ow5hmFiI5qphJ3DyFvUl1R
huDwg6I5+pIo0p56fO55Rjh6ljTKMrN6wOtuNOX7ud0qkg/o7D1Jqv8ULSB9Bt4TjkHjmF12WSgd
IZskX5gsqUcf5HW36HCHvvXhoeKVhhab35Q0+G4f/RaH7fyVxGzr92z4hdZBo6J93Ml2YnNAGhGx
WslYvxQma06wDZExxWc77hVdyjv+ZhvvgfzSh8yCvGKelz+Hd8lzV8HQhEM8LE7iUwe3+u/cn9k8
FjBz+RCK4t0JmK6RELe3wBxNpirqnYKnM7qef7CAG6yQaLjRVjHgpiPFbI/EQjy2qX+5TO087dBY
toPLaAMDsoez/a1AbA4A5d+c/RWxMH7B7qLnBDlrcFjltwrOrLpqWa8Oc6N4RP4H2er126A1Ncnl
ui5EVXG514EJuYuc6vmHAfD+t29pHBFChUvd8IV0P54HUpW+X7mEazvIQiAHNGzs38Djr6+4w74M
vKw0QZ/pGEiQF/7UxjVP5pqMyvBH8t3IzghI0OPLneZXK5XW/4piY8j1kz+Rul2UAXQcZo6MyJyu
ozFqthPXymXW2dG/XXgraVzK12z51lWMuyVLrnYXW5XMZFb3Mi7WDFVyq+jCAMcDnznMLKW63Fr9
qeEoh6ubqiOw9G2hQG24k00HY4O4k2zmETDrc/tjp2Ft10MURSVWF0gNLPcWt+oYCQvpwCfbYi1u
q9MsaySssreprr7vidhPqF6PD4ULhj+b0JNsnGSRCLCEwKy2fKBqTUsRWOu1KGMei38PqyUTRR2Q
mnQZrfu+hquCN9eLQFBNE0Tzuhb5colMBjm+cAYMCoC/0uPGpnXejFPXM3CCTkB3WMowOC2sHYrZ
qTIHAmroloEGXYrsxKCDHesIUdHoJkeC/PKU6rj+YjObJNiVPDivxAbdrnzbuwj3NGR/sQUGOHnx
Z7hC8IqC4gUsemiim2u3jT2R8EdkfDILE4uABNwFj0fgJeMBGMltrIA7d5QWJyf1lRVipgTqNzzx
hOIRdaAO3mnusj/QvPJrJA20RU2zA4pqRW3KesNWi9Lxz6mtEdpJAgB6iO42V2vIwfEz9xdiHRST
Qf8h4YZWx8aT6lPoipNEgpip0rTUdymfEY/lB9LKogRxvcq4dtaqPoif302/+ROpGnGkGEJbyeqv
eah2zjX5zOjW4oSkx2FyymS6XkRz9oE4ODNxlVrRD/PAbyDiZytc/NPy1GcFSjcyTk9NNqdWImaN
bV1ftSm7zdWSRRPyLB0UrM72AOilBDr/9+ZbJQBXfzuVSXMfk7/vTvDK69i08W2k95bwufXnMLfo
BwEuZpmu2ijBE4TZmXpEt4Bdj/1jHoFR5+FRLPz2T1dwv6kUW8GmAO4mB8TwQN27Yfe2GMg8StQs
BTP8GIV27+uYGby9epqOJ8pH5zC5mSlkM5vI+VKUNH/i+iOi0wBRw864h4xMDfnP3tU24Q2x/S8w
9ICHgKu7yC5rzO0mKdw7AlUi2/tkz03ZaQg/NUr/RUbvvDjuS8r9IlJGTmkHyzCHVC7EZJE2z0Dx
E7KtCd6/jnNW7nnBLZXFUAkPgZewcf9lv4UIVukKxR+RWxCgT6j3JV7uZ4Bw2yY7uN2wu6JB2F4P
Pjz/qRae2H7vas+/UfY9LZtcJiGQKPhDsyA6VSz1YGjWGye+U1VVK/2UT+K62f4ZDDfvHu/oMBY9
9T6k42Bs59+88nMAC94MRhd/sIdn+Aw+MPlvIl2PGS3bWrHje1QW4+MY1jt2afTQEKm8Ayf8Itv4
iy2+zPt2n+r+jIkZ+S+gY6FQV4see2VD4xfCi8ZrWM9LW8XatHsOjfDun60CcoWwQtCpIXMpwDww
9yJaW2Kh+NT1GVAyY5Uad0a0TIKWXRZsfjV8RGdzcuw9bEKDutjL5LxmC1wYlEzL64YksYW0gLeE
E5H1+qOuw3A9fgcLFnmNcduTXqcTBZNwwfco3MGo/zmi80bylMpgIj6bwvniUzUshwtvPoOCe8h1
+r47pZwM0fZBRwDv8Qz5cvDZCYbFQcp8nLuZgBI1rLG26nzZ1djDZwEFIArhzwfjpZKlmCxbGiJg
PexG1B6+8XJcnZW6+KOcVKu2C1Sb3hobuwT82wOSSJHsoDmKJITWAwJH5SY2euYHoHLddDbUHICB
7Po5M6/ceYUgInSP2TSGLR9d4M3yjYTJ5Zuc/Z/kq/vH2cEBDIqZeFPqhiPL04RGDLO62O/+gftd
tUgM1mF3pdFN8BILLwrfr9Rhbed7/wJSmWMc3s5IMQeudCVwqMML5eEIQXFhi3SiVFK6njidtyv8
Gk07fERQzhNesRl7ffdO1EgUNfoSsx3S96YuIOO0ATu2hCmqoQi07Fq5yuXywwtEx/y59z9Xgg9W
Cia0lD3pnUxzhAy+h6pEvE+MPky9HewXANqIGZzMeMqZm4KFlhKSaPNSOKQDTmmgydb8QtimQMkZ
8ug3/+1VJeLdkM6TXdIqfJMnhb4UWIauoVPJ1CMRiiE3XSmQ5vwkbdjIXjgkvjETxfiUi6Hrf3oi
OZ1DyyB6sqlUuiY5Znf5LxDT5DLIQJGS1LCleJnYIDUg7uZ2yZinJzjfsoAiE5anDj9NqwjFPEpo
XxScEHBRdnQNRyGLTIcZX+h0ktjPFq8aEJXkSFoUchRltoYNI5K7T0KF7gyS9fs6uXEndLKrpfP3
X1Rjba8x6I2KptQNNvgqqTVw4hr/uM9kOQS4V9B19IqnJzdccyE50ucufGYxge3zsu9e0AU1AXKO
WVvi1i/MNamPDNiuy1Lto9gGw/kIvDIWKoVjn0RzAw6Ks0qoJ7ERp9wvcvRH5u38gr9G4lMQbHqj
2t9zw0WFwbEIPrx3fVG+pjYjeJCH/4SgN7kPOTIv9V7pV5NjtVtbR7dlIHHGegrxr0JDVHEkEBhv
DxQiAo/wV9BKkEfUgcB4XeZ7jQOBQUAh2/3F5D/3DzOHqip86UriO6nyvqmwRQG8ZBFTVYKTSJ6c
9AkkH7By6I97uv/mhVwKIDIXiyKzSqQaLN4ZSIeQSxTk2F6Uo+fMPyMB7sSxIjOYkMHwnKVp+7fg
FqdgoO/KgDNBEW4dkcfOC/kvE0q2hvcVgRmBFi+mtHhGve0jBc3aVWsy1ws7JKWzvOhaCJuXgnT0
kqI3HLX1qe1hn9sNr7Sjj0GBvPzKtgDBm/XsZpzcUlHvBM8ELRhtcuWmgwqkZgRj7ZBek0xttbkq
wLBU61lIhW9w4QG9EWlsQ2jcFH/kifTgoH0JJCBX7KplZ8MGKJ5mHK/ALnPEK9+oJeEMm1uLLC0V
THMWt0PSC5gceg4lLtVVYqdqBXAk4RNIPtqTlHaNNFUE0uEbkrUW0Ozjvon0K6wEwO6UN1kdPDq/
wSDc9yggjqzcX0y29jO+dMYAUfwkwLwMhZ+DG0SZsZjF8VTIUt2qextpiZjcb4PQEVjEptqr3fhk
77zZhEkdfud51HJF1kkbZszx4dCBanmDE1im2GNbF/ZDJbhEZT9RhmTd6M9xzkpfgwVBJl6MQ+eO
foPvwUnRgy7IL4Lbj41Dr4Utp0yqcqx8xe6Ut6kfloK15l21hslJlRTxCYgj3oVQup5JZzmOuB04
Zh7PH0TLV+AFiYxsFe7B3WSVE+8STDdRC0slMAJDctewXeOWiRjRM5H1WREBIvKjqvlGYfMveQJN
0F4zuY5ltkbdzZAOMnSY2eHsT5GJ/rERMqAoGUZiIOPHvLJ7JuZq9ZB8zF9pKxheJuWQkhMuK1QF
NFXvLbbefI7hMa4MPBEKkiUXbNqTMZA7OqUpo756sEAOkFrkQDuWmzhVZALoBRkgY1GZ0+EKSoN8
qupOiv3b3eqrgwhkKXeCJgNSjBMg9sEnbXyrX4a/xg3zxTE2n1UYtiONqFWIFOVCOhANz/XM7qHk
JkS53Rux17XjPgDr1nwjHDqkMI2DYjo+QQ58+yVH3FK1X786s7hKktrjS9WUU2S0qAt44D8/iNqh
S00AwabEoqxsgyheJfz88znGYgfTMIU5ONhD3EQRofS4/w4095x1MdKuCrkfA4mI/Vs/6Quux5rG
oGW7hke0oE8otVJviT2wCxAPFjau/BMe6W8PowZA2dO3OSpLfbaf1GdgoC5xO0wJV9tR1yD36xnb
FPMINMIXAojc2KLLXLON2sD1+muUTvb2M7hZlKJwk91qKsztdwuwvWjCGNJguWF//YrYHWS5XmL+
zwuWji5Ow9vy01RXanLp7LeBgRq7/mfK6F4QZaXnC/e+3C3vSGN/1qnUeMYmKNtc5LXEeVYLuoDK
YKr3ITZDYBNKiiA7BGDvdZWdYKPiz7XNbcrSuBHazGQgc9vuf6S3weGdABpET/ZmMFUiJ6K41nQP
SsMQI6JVc6/zu2Xe13M7MLzE6B5y4naZx3cS8NxmdJmKJw57xxu9o+duZIsRX2CWeWB9D/zUrRIc
1POLnkb/AusBi9cl1baKBxOdi13BFZ3xxFHd10a/G8t/TWjrh2cNTytXNP2dxvVSeqqFaUv0J5eR
OGOzegtL/aFZ1aBAW7RO6/FElOeCKymyyg91P29OkkQIQKo9MC2IoiuqRu+t+KuECTSSaqOVgX2a
ecZOcot+Qk4m6AM0ezm4RSDv3+Zn12jDRP3WjNlSPT2VaX/WmBj+RAB0YPb5JTrf/WBIbXQcpCaL
IvGv0gQuGKr45C42UeZiF06KRwwTCLbJ6vMqfuyrNf79rifDcdbgmWknrYbPCbFzXrEFMD8e+2wx
WKren+yN+YX5sAiJ0DpyjkUcgTDORRVob1knRGcm00x+UG1Ea0KPP3NuYBmuTzzCLiDA3oqyQTtm
U1qcOXJbnD1KNvkDcKuHUbGQ0RA9leIudomlIjM6dWNLjDDkFXmknhfT01WNlPNqxgV8Sm1nBwpA
UwFisF03x92jMewHhTMvJB6dcPCOiFXIWuNGTpIPWvKG8/njnV61u/04VMmkS6Yc2TO0A+S0E6++
tvOwnshsdnvRL1yiz0vA0cA64DL+DdajS4k2zGgTWEoZMgshH//ixHcg4W0xiyDZEvqTWDbSkv8C
Vw1hrVHlNjYq/lxNkrSR1QD676KdXwJ+ZIVtTrIWr2gJTDb95RAI7Wdu1J3hkStBb91ZF0D8uy+3
JkhsQOaH6lg9GbrlCA7245SLtwCd+BKst4C6EwFkcHCBZ8KVsOjdacTS+IIiJrySypValigOl0Z9
7+1lcHMXy51HSOmcqOKjqkOMV3pBxkaqS/UEhyG3dPpTyt1K/5mR59joeP5lQGSAg9knbVjv4wHv
ItXUPnOho9Y1yRb1mhleei6I9c74V/HUEQwhBmHSReTnG9EFQ0borGug9bKQJJfj9euFfzsT2Y14
XHBpQwlxFym/MpubRzhnR/jvQHUhLyQX3l8nIRw5kQ799c9bNe5yuQ5pll0s59w6Yvn6v2sWy+nE
u1rG91OlbNPXAVb2Zub9GdYKj8D6dTWNax6QHshMd+QuhTlxmxiaRP7s0deKhz+kGvfolGKlJekB
nZtXGzhNtx7hCxWmiMbM67c2x1LD7E0L4rd6wSS4kdre3UL9mFsa6nGefB29iaquEkjm8vQ/xhru
776o3C27Ix/kX+uCfUkwJw295UNHqk4NKgQsbZvCRsDf7l9qIfgSD50Dvoo71K6Hz74tv0Q3YAs8
GROUwjjgfjm4/xjypDFl+gjPWmcvRdzIcN9QcicxK8adSlsfFHh1UilP+vgPkBodbNIqj2+1IK5A
5K1ewqfK8hBOMlRxLjBwndkLgBWhZoEnEOlM/RI+wwlMhGSbHId6Ua5cpLwC45jjLaYiyXjsXTZs
IEIEq6xRIB5WkPdpJKNiSzlGobAzcbZ5nUYtGy4jk3r3MkjuA31yO2F+6Ie549Sf7UA6kU/Vk4Ch
izhCN5llV5wzIWRrNmgzUmLoAsK6nrVbOuQD0xCm5DSsxli7u+wsU2GlPhGEgAMH3aljghFjqYEr
Ngnf6y42xRKU1MquLz5il8VY2jf80dRMYFlyA3B/CeaVtsxd9m8RNE6WLKQgbrPH/eH5D177g0+I
VwkEiuoyP6sK+qgCiSaanXjwn1N+wF6q+lLmKMBwTBs9IZDkCeu41sBh3N28O+/xSTLCo7+1X9bz
FW8jT4EoFcMCfGNmRbw5fEMCI+9kdzatOG+YYNv7ypbl+zIw5eDF2XuJIjf2OP0DTy4Q+lyIolGL
nOPIhwyweI4F5LnGDkOL6FSYMnfXdTUt2kejXplmiMRT6dQ+4sqVXZYr1GBEftiy9ZcZ5azeDlSy
EFS2O+FOjPEUCzSpEMAm0DRqfljsC15wgAmwt3wS47nSOSLdNZdoF8wGuaPgy/OIUlHKLSfT8FEV
hntJwtZ+zmrlSNHpCItjPvskeY6ofRy9JyzmPoSRTi6tdcPixNhzqtIbQTEMgkOhojw1xhVF6wPB
u+YbY/Vqa0k5iR+XZKVSRQyM7fd+TzCLJL1p46jYAIbdRq9E/LY+vpUx8krOdhVgGzhiaVxzN7dm
dd9/mZel4/Qu5RIqra3Y0ssTZdhzeXqyf4kAn73wIzsSR0RQQA4Ycl9G6yVePPqEzHhiQHPKt9L6
auRMwMY7qEF3DuZigzrvhaCBV/j16wD7HqSloNRrNmg7uSUkPn7LR7ndH1fH8sCxnFjB+SW9XZPy
8E9Y6AhldbNIXad5XKHUuhEw18kd6LCiSFwzK/iF95ppRBwZLlcFZuyui2nrd4ZxHONUQX8+mU8J
0czMKnrpZ2BFajDzGD0RCpEyvKuw/TrdUriFNbDn613QAkZmYUpCVkw5OM28nKeQKnea2FssLtAK
2E3lo5BZXCKgWTo8XVzYsDGf8WM/ht3+I5s1F5DsIRsabtXw+1FegKhe+J12irVepwoWyAnJLy7O
1fLLrqOv6DgLptKnIohIKAp3m//Kmmqfq9MAtBoPPFN8Q8FyenwURVPodLAAwgYhs6CA5ZovsHnn
q7dk2pbwRBs4wnBzZuli70QC/lQms7Zu/o3O+EGTT9KPAY5k2jcq2uYr3VkgVmuSePfbqKHt4I4b
Yn0kze531+PLJTgwp1gARIcP1LpnD+D+HeY3vMAylPmmVainu6yNhp2ET+2AgRt+XQDC7PoM2lth
aXUxmNE0yqxqIIofHf39iXCutakNgxWmrKrNyDHCBz7OowlOpAjUTsVyzR33FS6oQLqM0G7gmxVC
XG6nyUSsptl8UvLY5Ec8AwWBQIRX0o9wasv8aROiXx7tmbv+rsSUbjtpNTXVzJ/DC2TV0et6omj7
1deva6a9TBG5Uxg+v/RATcoomFqxL3ApHqiuKSK8QsdHxm2UbYeR8MK5+UcIKiepENQMuLLl0GBP
3J5hG8X09JNC96Eux+slTYvBDiBq7w87mXQm+P0lpEfbb+libA9wxPiysvuwG1ghzMoJ1hbGlXMQ
bFYYj4QhhVBirQHxMlhxI0xvoIA3UUKWCKC1iBRyeXs6wgklEHmgdglxzPHvqmx9py40AQHrWKRS
eFQnJKpNaAFcd9W6MRKS1Lfch+naPOt88BsT9WN9YXe9y5Ndyqtu8Y2BGryvWPjatGwwH13X55/h
xhXCMTcbHINZHLTG27Y6ryZv1dLFvY/Pjw3wXh1aB1OSmIrIryGFdcHD0h2vXTTn8LefvXXfhgd/
shnxNbkUl5xj+V9iCYeBwiCs5KUekwzkvLfCxIjJed860bERDvo9b15m3rZLjhJT5gg3zSfOumwo
jlbHr7mozSiw6C8gd3m4pnlFdoHIc2beDKZcSyqNeBP3bMD091aenkSXnj4uloFfGDiEzX7k/D/z
GLuYGoEYSsCnUrNEPhsPXt/BXf33UaSRL0/hCj/rvQ+LTJaBwB2riTytlKfWGZ9893v+YrvE1h+H
SbpBgkgoJT8oq0993E75PkHh3N6JfuhDm3FfHZunK/qPIp1Zp9zs3CuADYmtWV2qm5s7wpAx3Wa1
dOWVfwhHfbtaKYAQUtbq63AB+wTkS4a8/q+azySaDxO071hk8rLY+cn2PQiNPeOT53Qd/kL2WMYw
jyPqVdcD7AQT1sYDiS/rCEazV8Rbkd8LlW9uMtQPWnMJpUpKaCqi9tR+arJfaezO3YZAqbNW1764
kAhO/5qFq0FZtBRrIBJOMKC7w6ZjuuonGbWYUE6K9lVP9RwjRYbZFqFyNpAmVa2lh96vc/Jk8bGW
khokDQz5yLU1wiaiPRRUvCvo3Ct8qXGci4LWstCh9gY4nGg/bhwHrrfSkSe7yDKeP7yECSg8M52n
XNslqCLtKSXThcpGp+xODTTlDEFQFrYYP3NkUYJLiMm1mMTcknEtCHsqIcY2Id5TImVplyDe0QMq
DXan4t3xXcIJ77UduKop/SuRCJeqkHzEC4cc++MN1y/ZkwiJiwHDwBtYgmMbydwb1mztKALSSL/y
tzu9JdY8fDEybEF8sJ57f5IZjIktdHRMiihss2RKV0FR/G0ppjpetm3SWY3qpp0c3Q2sgR13dooc
9MhdIjHeXr6Fzlbn0O4teP+36STRG5kj+6ela+vZ4Djuf3v/EV/5hGAR7KuU1y+acJiZT3AEPNNM
VpIJTEEBQU7RKFGhmAMrVL2IzXAEInUIFaFrL2jDFkK1VpOgc1r1iyavendpqaMY8VTIdbcd3CgW
TTHeEvgSgPfJrj/wmIVkCjCADiJZEBdQJnSq/IpUgVfUFvBH+mYwrz4t56psVBX8vHGd9zi3dOTX
0coSE8Eq+o0KieDGnYsMWQ2bGZL4mr0bbl1RR/K93jz17wEQ3vO38qolijrK+bbl4i9+XzaPAbFc
TYLqs1YZDoSMbVWBf5l12Bvq8ehCvijNnJb6exOY8dAQCbBLKQx0pu90Qw8YjLNgwPD61XXcFZBT
KCdPqbOleTf+q2aiEKFWd4Gh46Yqp9fS89inqY5vmfUi7Xtn19pLADB6FKfNV04CjdlWDQ2C6sMR
ci3XJB0OzyarA4QFt+jk+tkgJvBxmoZUTqiRS/wIXqBNGd9rVHlm91uUJXHI/gNV8SSLCci3ZfCa
3KAainSFeIp7n+nxIZDRP4bl6ygXrUNImgS7WVFagv+/f4UMHbc+bCHuxP+kMXu0nSagaW9B5USL
wJso4HK7+WnGtjLB/JipWE9VCxhwd8uS/RcjahIS/HMViPNHUCa2JfmNMJftuln2H9F5zYwyLHrA
55/J2bv8fDyBFS++HeKN/CPkdtkTTvEw7szCJeJXXl3MZfO/9+GXgTybQOr+OdBSoViSwGHvfivk
iv40xJeYatCp0qipxnMqXbipsi927SarmQ+ZonzrUnmE3Ydpt4kOdokeig7TgcCxdd+z90OHxa9p
A5UeHmbzNShw6R6vnruZJ4dyEqidJKozji86CXt0kmB7dNFEkzpXAo7TSWlCm+T7XE6PkehQYT6S
2OYz7Al59gkRTFFPOuQav0HXs6Lum5AcKNFfwECS4EYhAG7TpIGlCYubvK15LDQWHL4T8QcAs01M
C4RCeCLiIHFvB4eU4GZg1yKRPg1ViYqqsrUdRlvL3rb8MAaokcfurc/cXz+aMKTxQRdpCqHqyUvL
Vf2/LJjNK4erLzoSLgwRZHZXuZFxSmEfRKXZ7xtBy8/joo2bdq0jcXcT7LS96ZQMgk6dA+qwuvSC
Gmov4dP34PGMHJheTb1pR9b97+QploA2KyWUqVlnihxI3ywgGherSXq8DoNB/Z3t4wxETNLj40iV
sGuKOCCikQ/P5LYX/CbqTvJu/Bpxkl1qSlVOzMozsii+Vldx5/HJ7m/YhWA/5pajWYJ19b8q9Axy
iqjCHgmBH7XKdC3yHYlHzs/H8W+eUIxR8WJ8djLGDHqV4x812OR7zcMFVgmRjEVCcViND7AqW0hW
qGDuK8XU6eb3/R7CzEFrR5sUYR9X6jCbsHlhp7yvAoAeXbI15M312R0rZl8F5FcjAN6ZgR3i0GkW
Rwl7DzEjPXoFz3yMsL3q0DINwoOP+oFP5DKiPt4puzQ0ng4VQ/w/wzKc/FAaU1O+WDuYUuF4JfAB
uvg9VvMI8g3ljcVUZHe6wmosiDcSvhOcvZEpNjx3XFZzunp+M9SdZs2g58VHvx/v6QwYf+mKYlv1
3DDYKfKcxdx1uxxQQOidknqEO/GVwy2zVMS60K/bgHuFA1P6dQFRqXeuzbnpUXn1xRAf+XwzKMZT
OBVozf1qkyhx/i9ZiIZ0uCPASprQaixDywyAow6fUPktF4PFKR3U0NtHZpfdlYdKeaqPtWO8nLwV
HPAuhP1h0EfxQDE/6Rp7wL40u+ESsIagfVDO8FBS2tWbXTpX8L8621uappQjxkoZyWNrhO68norJ
BkrmvQfhXg2EU7Q4TCewhJKajI9LVA/NapP7xsp46bP5lJ7bvt7NbZIo1RldA+YWc1CLAKTva9EC
r5LsBjbvf+aMwSPpJJi1dIuzoto23OfcmA9kyMSsYm8vt0qdFD+6ugmcASOrj8VwV85VA9XRm3ae
mJ5GMJ7GHaEnykRayFCWQ5EF+DRtqXhpNGg1LZa2vVbm3qz9U65BMjqM6VjqRJpZMp4pUcEGTjqi
5FnirvORc9uCdO1DmNIZt2NMn0fzBnULl7hHErWgoaK6RLBkEbqJQt2cHfuVK6wPZyMav9TASCnJ
GPMdVV5/kMjoUn86+xJqmoU9jdAE6RbLrMwvF2mkKU6OJNg7ijbrvN6jpAyVUE2qxzcAU9VP4Vz0
sY2oSdwxbp1F+OKUvY165GXGWypU8gbSEAq5s5DHLnlz4+vU6S785GqhXDUvJ72wWZ5X2njVyVnW
YufsPA7GyS6zbrxuxFa5rXTe6G/XvVRqH/9FKy8SkSdg12qwl1/IxSM777temQ/vSgMLxuKycz75
yEZ4s3leXFezgiJ7YUtxcjxAx089naSyGEViHz0r/sDYUH1QV67DWKoTpHOMK5hrEb/xu41TDKWY
WDFOf8hMB1/VjNQ0dXpQEQ4I2tHfga8bIoF9v0Hn6i6yEfPsGw0BWdXqJgiY48Jh4tpouFSgr1w7
4gdQ7R8XorAfShEYugp2AYsjEiAsimEtmf21utj4imCmDu05iPotd48bEEdj4tnh0y7Hiw3Wgcdj
j9VJ17ARNG/pcK2kEA5T+1kQBo+JU1CRD3Dwf1bSZ/ZeotZtuiAp8n5+7BBNLNybkw2+m3pYKgn7
xN6DikdDaOus/GR0dDnR6l/xWcjVtrIQAHTNfc4JB3JPP24VXnWGIPyxgESuEcRMkqa6ExJtGhIX
0m9RzMhj9d8bgExIT5OVJ8e09m2mk8xv1179M0/0Z5dONm9nlB8IwpkmlzaQfsXMN1vT7tqw3C5K
U09ksGvysEUVV09ws3uCfDQQ3lsvC3AGCmDZtqmDewtGPonizgU9u1F7mRHbptYYoAb8WOhcSj7/
DMzLCLFKPWQSeWAFx/lY8Nlvy3tMgRST3nd8YEAVlguAfJMWQiwDnLqwM3iELUPgSnQSEFWYkvgm
eoHqwkr0dSBooouygq6TPUaMdyCbXL+Y1abArSlTXLTEvQ2m0ehfMKqwXiooiEJtZohJbCd06PNk
DqwtQt9WQSYz7vMF8wmjzuAQxZ751wiYRlZdeCx6GuN422EIdza74BSPqNrJxZM/Lb2XDCa/4bTb
v/FR4oWM/AgEKh5lBQVsqjdBn9clFAsOaqePFpF6/AIJTMjx/jXRv/xY3hcYCHnyoZ0Uu2FeLJ0c
p/pzXDAiiG1V/Z8NiltGEIQAybIz+8aQZqLeBmzudIi4LWSfHYfhPxXsAEqtayu/t7wYra2PEko6
kxTiawNx1ezbx0He189hXZRgreQ40MtiANix9tRHyhQcmABOG5ZJQ3IvwUXI6fqL7ELvc6+fFYms
7bkeda2SOSXPTAvcDg2V9IojVcVo12FT+oSLxQQnD5J+BPg7gle84H/cJiLPvpNbtdofESJKVTX0
OSMr5KM9YSpJ044HQYVMqCM1E9zVGKSpxlA2Rn2YdzM3OWjxzPWG/woxYOcEiLxf6SBt7FUSSfYF
WZr9g7gTHOheN15nmNqQkRTf7BRpBbCBeo0s8FdbkAyvoDRsZY/gGtO6gwRcvaO2mu20LvGECqon
mjHGrknNVLg1p2kiJptEB7lRWH/tM/ps1z/pmksS83ExEhtJxVclxzh3nUDSEnlendD1EGzErbXS
qy8qhCyzBVfJdiAw4UqhwwHDvGB440cSQ+xUQfROL4T/8m7nU5/M0T8oI+oya/yRpXmHYK544MCU
nIZ/GEYLvghElXZkIEBLLgDpyDwBUkZyc8tKujEr5JgGhH/Fo5ANgP/GqAJbOzT+0duMcCqQdCFz
AI6fH7pe1jZtLmqH9jJ6qMn5XzZOly0zcKi7Wrb4SMvA3xYvOEpD+L1SS+eedEqju4Akd0+1573M
s4HrtUq1hQm9JDonTuSxilN9gGbmyS97mF1+XBSW/flTAx7wfPITYQpp8nW4+GuW1ki0b1NIw8cI
LiFWwjkIJZP7j4s/GWvto+7BIQOvMonyCx5HMsCLzF9wS6jVl45Geg80y0iqlQ/WeC7lcZqN/qMn
1EuRWTthhPU1GhXH63I5g2gZlamggjPC52Zv+O+Chu21e4Ffn77J+SRhoBMqcIvfhdzuGdlcQonS
hYLui3j17Rn0LweHvvlB2rIwTtwrY/08XoI6TD9jdVbRVKQmG3M+EeWwDiXv9lMes3VcggmB8K0b
sBFP+L1dZJmBhaMcBPtGLNr99rZy7Lx4bGOMueZQsAjwkN/o7qKEj0flR+u9JONF386OWrth/AC2
wvqfPgkZj1Dc5nveF/J3l7qTrmRdbGMHNNZTgl63Qx4+N4vCSMwo3JsUzWE8QeU1hk8wR3yNwaiN
Kba1pjqbyC/IJ3wje6vVwix4Un2IyFDr/Dvr+fuYnQMc1U36jcDcha0zFwxs4UgcZ35f3gtNmm+J
UOr+VBcwJo6EJVn01e4XE/oEhodIBFWiBSwuIPQO5mC3vaHluTOot8AJa+KSCzl+SXgPUv6nVdz1
f4qn1I+ipWkq/XG+n+tVyWjE/H4vNV7ZxAmE9rIbk0f+hbFHceyh7nT7UvpWWwTSQHiFlKL4g79l
d3Fr0zYUbjqCTvDMR+bNW4iSibsluY+Ugj+1+xwy/PON5O8mfcA8rU/5nTCemWfxtOjVF1Jx4MUX
5KwQsVuUFu+SJKUbXt88XW9yZrcOGRktqBJD1jFaiK+mwEWIXhwevKc0O5Ortf521v1AhUV8exIx
WGMZXOxSAzTIQZJ48EirGZP0gYP0EWMYnjT5uWjiyMBU7fHkfddX9AhQaJB/vm2jyXuGr2eDNo2d
qjroYApIq4FSROdOLwUN0MP7xiUKgiHNqvo9tpUeRRBdoTvVlSrSZZpVNuA2M1rSQTM7UOYgF95R
xJt58uAygXf7iceEzo9n21O0cgJHXwjaNkyaG36Yj9IeFV+MYHQSiGl/mK8HtQFN/cXz6nIq9bK9
Bm34Mz1GS1yglDfkz2tW7H6VNl39hAoHQBe54FGX6+ZJ/VYC+aJn8vlCet1GDs+0o26Inb3i4PX4
pQikQRR2yZr8PCdtZbF+PSCKuMlJM39DMIiCXKdMw76sHk5UYYdSq1nV1yoyjJjDxK4C7F3Cr6rQ
W6mOskrxsI3H0FjZstKGPn0PzzhE0orejGZfp4+7MX7T1RvQGBjRMZABnEz40bzFbUtwjowzYIzg
7JF7oubYkxeEaUYkMfOP+2oqjqsGsXu2A/Y86tGXdkezKUbk/PGTezQlaoxLKA5mpjrA6tNW4mZX
YKRgYkSndi3Y6D0224DVmNHFYm1qiVGrFIGftupPOdGOm9tiBmucnEJr0dV0IMYC/sbMX0sC1oxs
ZOpHBWgZMqa3KIBXJPk373zN0jlbHf4zyeTySHU/DQmdhagdrl2ASBCromkR8rUvxSfewtp5psSW
I4GRgZ47HsCrPA9CDLrGJZSAnmMAfbrFbAajQLpadagneu3Fw9KqwbkxgiExg7KV5btKBB+3llXR
7sMHdJJ3yPuN9vZYpO76oYMh74f5v5iAi4QPw47ckowTuo/sCAviN936uW5881kdFBavjjT0c9Qt
IzmXCOqGEPvpUzUstERafUYXMX1puDEzK1/t3w5bttqlkh/wzXv4jOJI5A9eM/cyZssseWBpg2F0
fppfLqP7frVW/pT29alwtbKAuMOSnS1dXbAYpckd0JXmt0AZdfXMC8bcokrtvl62TGmgEtBdPfng
nAQz1xt7yINaVPjEklq288wUU2sFncO1vn4CQMr965mchmuWuPDX824fIWKSK82yTcS8b/DRdYhw
oFWLhPfDIJPTFKL3ICzV7Eya91qz3DxE/RrFOPlKBjTGdcgT6aXYxartFkWseARLpXWTYcLIQPRo
t8lolvCMO25qTSoNskf2xfGO5X22tync+IzNHluwu1LqDWquyO+VSxRjbD9gcQE6wY3UEd0b6kmP
aFi6cTb9BxNlfqiBi8uNosh5YnCLZ/Cm2On7nxDfSSLtM0cqQo1pDfjUiWhvVPmDYVpjs9FoCMOZ
byNZXTnAM4fXm7y2aYMiaQOs3Pie0pLiKpWIBeRJ+BKS/CVBhaFPjA9cbOa7omkP5A2hry4ELes1
o84G78MCR4NF6Wud8PubjhxnUfuB3niG56wZStLnFIPeyizAtVW/hZK3VbBIuysqegT5JpKa7g6M
tK7K9xuIfSlPIcRPZtnQel/sar5iJrlbKB1Q3b+2bycR6DBDE7HMb8b0GTrx+Z3cFPI9Nm7P0Ja8
rhwjE2zqsKpm7FaOWYAm4x16iAMasscf9IQmGEqM/+cJBTv83ETnSiafPWkTjsuNb9OsK+fbqgfe
HjgDTaMo8iGzvj/inc1SJpW1wX85sZ7uJ+/bvXMCigTA9ZdtTGqtK1uvj0XIFdKH0AYIl57j+9UQ
BjE2J4NDp98Kb/+WVwhglnIilPL9F4sb2sgF+HUvUOb2rVuvrTqvyNogbK6sVJyt+22usiR7iowC
CAWEDPxa0+uGiURZK51a/hYNawCgOjzibLJfSsiY2aEQ+8+sVoqXQ/86kD2UxQzVcznCCxSeoiP8
py3fvDSkQgLf79Tb1hGFOwbTYpJ1WUk7vPEnnCxs5FOzNK+TuGPjt886xSfCEH11T97UgIL94l35
aZdjJCAcIRaxYG0Ys4W+7M0M7vkP737V6TVVMjm3nJsEZ1jbnr4wAxIe3TL5qFtXnCTGOSEkMaro
EAwxoAZn2TvqHgAuxoy58utunjhOAfy0sC1v7z5/dWkKO8N5nriVoqMZaS4DT25p94xNJwEgq2/q
ZwaoLvC/tzSJy0fYhx7rKKuljdlUqUq32z8CUhimc6LD7xygwEW6TLpuGgydDZ8dnd0m9Z9ornXk
2ik0HzjsPbAD4NnlqbxesA4Xp+xIn9HFKA0V8xpgthbqUipDJvW+M2VCaO/RDNea7l3kN7Z5ylek
McSGf14ZYFsThqV45msiAPBR3bHJoV51x+SY6eSLpYPB17NGDU79Lh2HZ/9oOsMtcMhbML/1qwRP
ZErigteYTydNpebuV0/K1YComupHzXD+7O8+jE2a25o28n+ZeVl9kTr3AkxDHVaYG7Owk+oVpIUZ
KAWBHWuantYpfWMEKq5UNMTLDrDWmDXmiBrJ1MuZ4WhWc5KuDNkGWVporXxL4r/NPfOd3x4xTQeI
oA/8REQ+ENMcdm0jFLzjsTR8RW3YGEdoFmdBpl7WyBvlAuxdRv3X4qC6OTKPrwUHPtViU3U2UWTr
UGIeuz9JjmvHYW6ExT8lL+UItF0KNfrLIkN9kgjxeFVqTwCRiMlHJLhXMaQpG74OyVrzIkg5ZYWL
/asvR1sJvt1XlGW2g+iiIL5BltDFErcl2WfnvUnlnn0Qb1+imCYc4TLR2AFYOA03cQyZSnNqKMqv
DzEPdKd1tSEHqDKaBxGjCL6UWMWYlD0oIvepsMgcFmc1lc9kR/2StscDIItTTbwFZ89EVDfoF6kW
XMMJ3FpC5u+7z6KGNHDRC9QWi6JQiHPf2iJ2/CLJODLBCEnUf1BErOgzTl0R/WvbFCg9xwYIrE95
aE9isx8jGJw2z1hz79KredMn3nk7EeCUN0Hgvxkyf/B4q4kDEGPrG9IVyRxtFARe2+eZah4VlJ43
uGC4uwCd/7OarHkIBs1EMfpqGbqbY1JLDqLRN2rZbA01PObThnVY3eTbea4OPGmM2HDtzgrdWJV+
WTprIuZ39VZpNS1mcQH2HhV7Vp7d0keX55Iqb63ObJpMgLY7Paz/WnenbfBY3xWJKHtqRoENBXkZ
Dqp4he8kdcEzgvpMHv6ZPonok111qQDxA9TWhfCz0uvZW18/96lCMmMydnkS9RNpVaQZ5zP5xoxr
TP9+DLM6bj6XtlmMlVvpIds/BYoqfQIU7cXxiutEYDlAIb30CwnCagjkBHypComm/pcdwpYkubT1
yy3AUko8pd3PN2H2CLrPrchmbq4ZoSFZvXz6Us1CDC9sSyfv8vMYF0CgFjWXk4oLkgf6Tywwx9cl
rSR9ccRRYHNQELMy+/eBxKt2ZLxUSweHICsKNhzRQJi/nv/uJ5lbapEu6k6AwfpsqI8CqprDwmiY
tWDh9pMyy1NMLVcFJHUDLmyIwi+zQh4Zu6tZDBEbbq6I+nW8O0Dfqb3QuyDuBEecGuboRvHdsCbC
OwNdRw0cN8maY1/w6iujKf4Q8hO1WSY0J+Bz62vDF2iTdzGUj+6KXFSg8QHQYLTAuSmAOR5xd/ta
YGO8oLM7zNol+G3hK/gTcTr6ocaLnO+ti9liykiKY13cj9xV4sm+zXg/NitX9OnlPSBymHZlq1YV
zLl6ddElmJgC4d2yW84gdLa6JYHgOzYrG76UDSWSt9T3ZSf/qC1k+Y7V5L47yhsLSeI+KmPXQ87w
7jW9+SsTgyvCA5c0NFcVTo3jDx+rFoCsT5fc/V/BfJ60i6bIfi6d7aQoAR3ndUmVX2NN6+ZtMosu
jH9JOVilDknC33nSzfrP39gZnoLfsxUHg8ZyCKpXoANpmqbTHL0w8GlFOU9NHO/6nbg9ys9nY5Tr
EzjnJIS60Hn3fP+UE/VlRhZ63c61x47annUlOaWsUzO+sH+pmT5NHQCm8tpAS2XMIUyTvSieZduY
bTAVqgUC6PocFsRqudcIrpaiwaAFhGdiMkp3Ymyu3x5CYcJ+RsDujLybx4d9LCa2WASHkcTYpYWb
ipX4B/F0Y0cCdID1sH+RtvuPdtBcTWiFsweYoNW5vSfxEP9/MRI42e/maBVrxr5a97Ea9X+c0P50
jcw6sP41VvDEnQ6pc3G2mUlrlHddzVhoHwvk+cCxD2PpzmH30lDo8p9leqkwB2VTlqKBlTt//97R
HNQn6Qp3CDIW+6EGYKE8AEOmQPy+QYz2rZApPSwqU7fTwK9a3AKZZhY2WUpH/AC5Zjlx6uWu5d51
VKFwKAZJ0/8YJdBavcvdHbe++svaEV4tOHDVK4B4/NdbU8dLdYv869uTrmbonv45AD/y+KC+M35+
br+azYi+0mNQhOzWXq0n/bISsUzW1gUyWuLxTZV9e6iCXWchpamwGA7Nl7jOSy8P4I1c0X7M0u5u
GkvB1kzzd6zm+i3y8jcsBKMi83d/vnDeF/Kj0r5bTH2S0yb6omNSVJ+0foYmcKBvdclZbBDUHGvL
jksR2ECuxsaqXs3xjNo14cKqu3W1cvsBu9XCaKQtut77AsPfClf5IV4y38ReuAu2GPikoX27F6yH
If6UJ4BiKv64MQRfAFLNPUhcM89/Su7vM0i/iXdqoaDfgyAYxTdtnqejVLTtdkkJFACsOzPHQp/S
VNwJQWLvG8Sp2HuSScrbzIiaxJTmIK7HU7WTihmS5jX2FbU5XVtki6iywbW8pAflok6nL8va3yVW
Fiy6/T3weupNjh6JDnUIEGZj6wwZNeGtzwQBOgAgEb/jZ/nKrdST59eeV8Wh4HL/WlaRjJHztCCk
4ymNIlgxMPoQCRZQcw0U9y2XufvH7m9MWZOj9d/3l9R1Bsy8pjNODG/YOyD0RWVNQWds+MMjeyLE
131wka1EHcGBpFhlEdw8Wci6bHFH82Q1CR6TfBKDqvwcIOvPlqyoz8YtED+tfi//0i+JJMd/P2R8
Ymxf/dXYTQNa69LAPKXAJRiVu+q13AZAaS42hksH9ubw+J4kIcW1t7m+/pMmDdMuuhvJoHG8u9dh
v3VCM2DC2aelIHFqqVtQMt/PuxSlDdhOumGdN8urRKZOwEBBlraAcM/vtlzVfnPQ+VxglxWdSZMN
3C6xXDIWF2nGo1LhGD4iXQsa6fRvkj5yI4pG5tYwlylqiRNR9vmi49cb0cCZIvMETBQbbEBDOe3o
NKkEi9qRj11912gcT/HYi3Vut6gIywT/v4Q8+3VBWYo/dEI6ES4xBLzQ1crrOhqYV4nOUfJfEOVU
Z+cEd9O0t0iwWVcdu2TNIect89VrhiWBrx3aaQkgR6i+RA7UxCEAb5CXJr0gBz1ywkIQIXtNLoHC
/3BKAvsuV2cqcdn2BOUFI1taHMuxu+hzl7VRfnNOPz58H7zbNKw/jaANpaPWQPVeu72yG5K5/Wan
AB1+KY/xJxlr7VFQYdgxIoFJOvCHl0UbdcGYXqUxCLU7NX4EHMNmh6adNZLsD3MoWxrBLYbnabY2
y8dY1CvtDsaraj/fuTbp6uORgqfZ0aKoEIbqotGhlQGJUxx0hH4qXojo7JzcHK0kCBf83Rw31GoW
aTyqdiAVsPd6aB0/oUCwV1rxrVIYtN3gdEhA7BSRRJvcGR0ycwsukFfQJ6hrCGZOHHi/r64VzeDS
hCN7TRTDEViRnSo1VDJdnXnGaYfsMDgTNap51fSj9fhgtC0qHVcgQLIvxCAAIsEBv0He2s/mVCMg
x3cczSAj3RPIALwsuyNs3kG7rNzbB4u9I/7j93q5hnJvVqsm/3a5Z3ieIQPO0aK1GKDiAJUuvkYL
grS4iLVH//JzcNjYBjtbgw+JKYo9teWP7YmPVUHVZCVc4Z5eTlyVDNsianeO8RjsXlFpoj9VQHvu
PmbqYBIqpI9lcfbsjB9NOOn2BZ88J4brGoOrywEsSvuWvuGvdcvd8uAfhCh7Oorr5fEmnxyfuNpF
BIlNL9CKeEWBwJLjA9Mz9PrmneOUe6CjDJXQvUzAJvq/rVrHBm8Zw1j5PhNBy6nYDAfWQYrLde4Y
MDmonBBaURXKW+zc5cSQEHhQkCcw2O0h7rPIxZFuJ2JDJdJOTxW4Ju0t9ewtQw12ufIwtcF9j2Se
NfGtWRmENWd+eDNxla6hB09CU208trDcwbF7FNQUU5zcbNA71V9yRKLpxlreJ780e8bbUHlRb0av
Q489Zm+AtrR9gGH2lVe6nykdMBZj9yd4P2rQ1Mlva0HlVMvh3oH1Ko6QJrfxPrbmBVIBaS8qbXYN
eocrUPiXesm+VeOSCjL/OLkWif/F0ZvgbXpqWu0wJZtBxQBa9a9liGY4QioHLbZ2YkECA3pmhZRm
9HFNmshqd2CcmaqCwyCPNhpNe+sUZJw4u67iz/u8K6e3WivWiEC4WN/THRb+2PVrbFPhsm1581+G
yYLkA98zdBAPQtNuMU8rBIjaqNtHZHJVGevNWj65VorPLDQR4EuvOBov0UL8Vi0pjNolxOYx+BLw
1g57mtPVQ1NUwwBrdKY1StqwikHiPmv6C2tXJWs1dqo+Xn+jljlUm8Gk1nwZPj2rnyAxktZPiavw
6CAgDT7LdBsnj9vemTOCA0NsAT5AyBmC3/ym6ZmOGq12F/nRKbWtvqE3TqDvTp7GXAua7TeWLLO2
/6g2No2eaXJNsOknDkaemUK5tZ4LKusO/bvGuAMc7jQE7FlqsMwcBNvYyibPM3MgW834lRcal1se
D/tZw8NNOqJc65hwIlYDdWc7Rsyo+Sy8eToO0/vSHhhe+wNA5kjjmj0BVCIfKW13wnlNkn9np4LT
gzWZZnrgfSzm3Mpvef50Fb5zBcPaXU7Vu6e4oJZqLG20tG9SgPhP3nQjwC2WdUhLO1xtB+LKayQq
ASM5Phc/10zHMmnViRzB2eXUo38Ptda9aRuA/fSyilKaheC+AUlWJRmx9Q0I1yNvdmvbyokjpwGR
l2qyL/nm6vxxZR5pEqOTS5/h04Nui0jW/IMO2zV2BPSWaXj7HoyKWt2cBggk84KNuoOKD3lr78uJ
Am5BV3F2vSWVaeUtRU9MELQJ+kDsMazhoMkWb0Dqkjz1BBLiR1I8kvuwP2kdr+F3t4sPnNZNGDAy
SbXAc1MUs2RSdzFHQf5Rz1clTDqBRM52xQKwwZk1NeI2QG43NMaHMWfMc8BOVhCzPZ4r/sw5bk/F
S4Robe7wI8UAJ44BeHmXdU0QFKi246YIhzxO+/xlUQbFnX9yrJaI/Pp3tLbJvxK0d6d9xiIc29gN
H2kk0T3bezDR6a7tAAIdLlL9nG+aX1P9qNfBYe6dgaf8WC9Sk8R2K0Bd53YNXelEpRhI8wlMl7+P
9Bk8Xy60o/z9tsJSv2OpP8nD1neWRaH0u4YG6SIXUaWxvxK77zpUgIcJeWqsRteUoFPFfo21Rgkm
JyRGfoFPambGG8F7EjK5ZMuWpOiyk69jm93LjEHqV4M20HQzUJunI908Wuuti+FNbuiO5e/9kpgi
7Ge7KsWHuh2mjhonPKgWJNh4wJRmcHP1dqUoIBWaqHTQHG2GCGEXBI4+Kl7RkGd1bFYEn/94f9uf
9Y/EJk5Hz4ntINEQuNJG2HMOLIuRwzCnnUb2FiBWJbAru+kqCccyP5qDrIbJdBQw8SpuURhUYmfH
+/xsqcGVSSpH5gPIcueVlvhg5zo3HWMYA8HnvNfpwZYmd0IUWUjY69NMG5PP13nILWM/jtiWjpU5
jAyPj0bifJI1aXLMnPvNm1Tf38lCk2pMGrXvYD33N6sWsV2e9NCd3pfzXyFal8TbU1wwqb2Htu6e
Op18H26BxjoyYnZRtlhhZL/bBQ0lA/IhT22ZE1wak9dhLClplBhzX2lIlPp7YvIG60EFz08gugDk
xxlfCOLCd8+TqLJmHJtFJeMHVZhcryCoSsgTUaB+LLA9LjIYZbXERD1V8OuYrX78kv03nLMRK28n
MbD2qWeFZL/6WivXuLN5k3aOvtHVneUSzK+lWPhiIJQR+nMkA1zcZefGdhcBHY1YPZscI92o9wRP
A6aZWAlb/XfVLzAXvpT2VrxLXHwGqZjVtdCxa1cODNMdXvgtJ31Ik8oSIAw/aQOjAvcv3PABllUq
EQle+j4IZmkOO9Rf7eloXGhr+VdO2v/e1gmXqSmUfss8ef1pMwvxpjUwCOr9Dd8o9a/tOQHqlXXO
4eIE/npRUvvxEsX+wjzBT6lUxfbKph5nZ86pi5M2sgFsGRGy098APhJDA4yuRN6dOkT62gbuL7fh
TWNpK0e+hq2kYkKYDktQj0FE4ig4AzXSh4yN8aetKe077IHM+CxJWRBUyVtdB15Fy8qzZl3WfvCj
kzhtb+6sTJZbwqL2o5BCvni71kkhDdOjyHxyWd8JapVSqLOmTRo7vZNAPWbN4Dy0uDsP4+Vap7XM
zfDNyoaz4lXnEenUUMVMPQ1yHrlt2exul8p48IUxKNUiJ0Mgf+cykjukXBFYXglwlxsTbqNCQAk8
RzT10us2V+5qmUk9C1dC5w8/UktFoXi19YQ1/tWStG3qLw9rirmpWqx2BkXcNQmrZbho6KsoC1lc
ORkSkefwZ282WlPOLM8UBB0Bjpi59UGuWcxP0+n+uRtOggjV2pfbuXtH/rnW/U/HC62bWihcUENT
3AQrC7B2E0eIZLkrwSfuNvthf/XMKDMpS/70HGRd/IO/uU7dMtGZEdCWxKteyJRyIkRmIKDfPu1v
ClWPNtxSpV8NKbEU+OMiNXQIBkyFmly6NatxBVqW2FKQ2Z/Kd3ivQMLGEdST5gJVKR0i25Ei497n
vWVHtlGfgxgw6N37EUaCP3H7Ovmo4mu+G+cNdtHuUsdQWCbGlQSeCp9We5Ky0DW1DfwFm/lbdJUX
Gu5k033oR3Le6L0MVo+qHEa8UT4VK/99lFHu/vHnJLoGk7qrGfWrDcelCtVmwN2M06Rki8q2T7kv
LwhfUJXgl+sGWeTMLW7p9lCgY6nkWoMiiTqOM1SSHccR9gHL60CwofjZA48DwKKRfs57JUS/LhzT
hUML5/nIDzjKpgUk5Mt5U5W0HkKVjVTDY5NsYBCLrtlhHlOth9mKru59g5rMP3T8UTNlg9TUF7DN
nIdTTGppdLPk1Daq5p9RhvrEHee6dVsWe8sCbS4a0K90e0LHNJFlGxZkSUFGCvdikX+u3fcX+5u5
VdBYOu7cD0TzWD1t6uPwrfVanVcZAkGLnrEtdRchb94id3ZlowDaH50jlF/F65FG7g1nK5hCtE8x
Pq8GgY5cyCW0u2SyokHN+TLJ35fjhKH60u6iza3jO+M5ybgifIj6tWUJhloudFYMtxKdb5pakQDF
7inR2NcAV9Nnlwq9cn1PP5U4Yu0CGIWbNBiWFRnIofA8anVIR68P1faBKoLZ/h9HRqJC63m5TMNX
UsevH9tYudQR7OA2ZGqYnCm0qDUURYKFrOyIQJbLeJecH8QVy3GjCV/sH1NCI3/qXe9Sj8elpbLw
5T+Fj+7k0aDXGeFJ/+R7jYW9a57IJO6dHpm9TKfEuRgD0hDZ4UAuLWLjowgxliLxqZGvmv/IzWc1
IuWzOCQUUHmQLAPz9b0CpNLxK/R/rsmT8+9LBjx/Ho1zx3I48SKMmhyRZoQzfcxUgkpCqWgMTnIN
3g8mJxUy6dtDLtNlm9l9xqFBkTh0o0s4YduBqFOv4brnt1aclGgFpdUlMNG7Zt89FF7u30jo4Nzt
FOMG0Sk+T5OFaBV93KNz2rKzYL//pVKJ1X8KSzoDhZvf/hn9/uS/VuFwTdS2+LYmuXBltD6QqGGO
5UoXLuNxZzUGdpPYVfsUiusxldXYqxfte/Dn34Pa1O0ZG0WgQmH2DsBbQcopJonKUmvl2H6VT7vW
KuvU3wBT8jpwDklVM1YPea5zMJEgQ56sMvUpMpj9CQJYAwTwjShnHvFbdqFJZBNDfAqD9UXlMeRM
OdFv4GbuN0Z5uytvsYUyeFACmE3gjkvk+MT/nofovE0h8vUMH9LUnHw57lyMSs0lV6PecxpDY+tT
AUHCBwMmj4+JLyPmwdGQsTSjjkg0drwwUqyW1rXenw/eqpiVI4LsELx3fxEV035LtiQB75I4yyie
1TYTR5lcTXJ79hkDHHLxg4ppnn/fR8ilrQ9JCYrXUDk/uh/8T5tKPvRLLlEbeGBEyO/Q8dfqKTVC
Zdm6NdcXRbGLTufjkfMw8o4lzHVA2KMvpJUDqBHswMoG+WkXGzbkl0JZaRWam5hlyocSopQpP4Vx
658/8NLKsDEKUArvC9MiD0mz1zzILYJTjxntr6njJpBLJ2Jv6U8xNeAv1O3ytcinvb7Xuu/dGAGz
rgb+A6WQ5hJ7S/NFNF68BdVv/l3IVMWvOBwp7a7RAfZeJdUcKlkElTQEpTJKdevm2xufkOKzal+d
emHoZNaAFTlxB1gvgNK5504HpxG9cqPiulMX5R2RUxOA6sx2bYQWqd3f8WzSO7XhnYTRw12xSE9l
EvTmuGTN1bZ+Kdq44fjk08fcrVU1FqxhkV3NUYbrKq/oLdxm9uee79b54G9MmLxJf/6VqUo7/FD9
ukl/Ik3RtOBbGCz8xeNIjzRF504aYaShErMHyWd/tdNNKnD4lZ6NkuYn6yi4OF8LfY9CO2NjsZxl
NMgXukR0M5UpjWzIOTZMY+/QlJ4bnlTBwL/0iMLDy/+cwR1gdrAhXcIrSHkKPAKUUfw2zQo+jifX
Oig8L6lpoKsb1qc95K0tGloA3o2rEHmJFvrGTUgr1MmPADZJcS4kafKr0eVAX5By34Gp1UzBUJbI
vOfJStlwtWHgKU2iCyTq3Yr55zM4HggqA695RXtkDbghcmPzg4feORg3k5gwqkdvMVt9bTXgIjtD
DUUemv8my02wolp+wGiRO7Tc8FkCPD7S258poxx1zBKdHT2v4oMJr/xrmxgZr3zVo1HHJMfja+i1
LWK18NapMkqYWcZPFbCFMjKcB0Iv8VCCLH+yaxl5Ff4uy79eROFRTrxJFkIuodj+Hzs2j6rlSAP+
h3Y3053Sc2Y7sGQeiuIqtfdFrWl/dvB7VCnFzYgUmYhlRciX0ZA1bYdoqygrXNiaccFvd0wrFqZr
acaX3w2OswiHRQzZSMS2Z/s9jI11cAn+NRbAetNMlPWw+Do/NHqj4Kyqy8TcGpXDJ74b+Mmetz4n
OMphBlsJz0w6jcO2QIJf1lqJw5hTjgxxQApWlpLvSzcDX5J+XEIZ5mQi9fOoeVAJsBFz0YJGwiFV
TLteFEGafQ6IQxF47GyHkuoC9bfo+Lzh+cpejEy+1G60SMOB/0qPfivrdnPKzNPHsy96o3tGHmH0
fi23fk3SoQPwaKKAKFfdbLcVi+26byDXWf/TeeTZitzXaTiSPYEvUMiOeUAmpBiAuLeusiLVZ+X2
epeqwT9TDTwbNbRijgkJCQNXRIBO95clLhr4ZikbZIQcEq6ASRYY9/LxbqXFHL4GHwhjZsl11tKd
0InVUy57VVVrrFnW8AnRpJ3kBGDgOZxQgbhjP3oIdmIuFqX/HEsQG55+MEaNd8jPciwhKxqXUF3i
dboV2f2AFO1oB46OgrBdWGSCncpA1bvyDqAOpEAjYRx2QwYM0Qj0jwftLcw10yoOLAFOkDsW1ay5
YzGEQvAB7ME+Fqkic+RT5Toq1Ei+gWZrjKPKvhN0M/lWplpYC5mljBqCon4hd4RebBuJ2WolCHc4
xNv44bgRDdVZijR9XWn2afS5uwUj4VIl29DeOp1XYEFqvw5UFo5qHEw7lEtzGYNWomCCASjsG/0V
q7qxvaa+oiZugP1tZPpMwqVeG4hrZm8yPbx1SxS+E7ibyHfvHKfACBS8RwlTWvsVQk//hHlbIYf7
Sv9MjGrEI1vS9V3jvTcmxdZI4nDKwVui5PYB6PHdZgk0ASI5RsvvpoUThECI6I/mvQVdMnPzj53E
uEL9Q3yBE70cqE/XbJuB2hK4PiAvlzHWUygiDRoO1M1mEde3v9xq05cOH8MUFsgivL/Mq+azxOVu
qC9/gebrQ3VuMUomZDqv01WRaF9WnpaNhSKIhK1W3iWZ0RY4cCwaWfUWuAGMiToiYhVqyJ46e6y/
qWkd2HSCxoGTKt7FybxUl7ovM4Q7Dv2j1/RDjy1sMG7lXtuU3rly82IbsAWyuuoUEGxwCxdRzF4f
YgDcqoUmFenS1ur3urH9H6kvknKNTssZp8b5BZ/4+xeEjehNofOV21dot2i0wVfFQ/ir8Pq5bbfF
omhhgF2nMO76ZRB1zmEaQze882FU0MvnEsHl04+OM3DLb8S95dDn6exJ89hBMomH/XR6N8gRigqY
WFgwaQ1LM5YkGAZRc5V1rsG3zUHHJ2oFmy/IMIR1TI7y74FBWneoCEpceIj8YhYrDRmWZ/Sl9Usy
POqE650ls/BmnaSAHCFmuo2eABlw3IIMuSfY6Of7IjTz2lXTh96xFgzFeeY4gJ4vBUfWnzkBrRZs
Hz1NmzCA0PhIcKXgE13Mk1EThbX+IM9dpERm2bLxRXnS55FDHi+22MyxAB7/m8YfnNIw7OEUiw9T
9HicC2ZSOLiRAp1k8YUMOYu/11GijFCmoaXRsG1LUGe2Y4NeyKTG6t67hHjVGiRt11AdL6K7Hydl
jtCceaYmSyKLCXy3otpsp0+ujPoRDMb+o65dZDnhG9djEERfYvs2zPv3e6DWYj8I8ivQYY+Haw3B
CiBAwNwS7PzgF+T2VlV/QuQ8ruOaFUDKuX9kn72834em6SYfP9lBerY8t1Nj3vlAp6KC3M5+Y7J+
CVP7EPKMBsRA70mSp6XlrAr5ABQdoRXSOWqIHe8gAHSXjGS9/u/dY14H/wDAr1xPia2cOAw74Ycm
yLe3U8AOKC5oK7omBAWv5BhRMCKkHVWn9AYcgz9THX2MboC2roncBniFMJ45TpI4JVqSREfzlI3M
CYRA4LqPTotWamLsAOPdpyTEP8cICjHM4pwww2Q3JwZlLWFjjW6PUL+EBa5io/5r0VdJo9xA9W1i
fmafTag30RggqiOmcy1uYTE6f3L47Zfiyr+CANKBYDVgZHCNjNYRMHJTncs18Xjqw7M62W3SZprV
c1vMMy+VOal29TCw40jWxz1jV7pbVtz3ekiCLdXOcIjiqvhyCGyVFsj/970YoO/r7ZRtVVcaG4SZ
tFOab6rNZ12injwpI63bRFn8SuyfHZ0wfzUZ59lzMQw0NV0pNZKPVW/l1AL4sa+Tlw4xM53m4fia
fgHm+7iG5mxOwI0KFJ3SsWj/ezzEBxK2m0y+M5ralY34KxmeMkdGRL2Flt1ERZcoIzey9CT9az8F
boegZbBGYaCj2LrCQ3Dypd3LmxxFPNb6d4ul0AH64qVIeWvr2k9SHFj1a3bWUlM0yyicw1X7sPUb
AwRSN1kT4Jhc+C323qlmhqy1Eu8JRipZaFm1DiVxak1oeJGaUPuY7vjVfjcZVPJto34GMWFc4ESk
q3tjpokTYGs9DRFbzwZpRXTOk0nE+RuNjOvzx5uZdeM8ISVoPlES819zHfC2sPJ7MMOj/DQZmb60
EQVJDMm6FYS40su1VAudIBw1l/khudSgNKobQZHwII//NaC6RmpJ3VmDi/N6
`protect end_protected

