

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
DZrqnYwqMkKoBvgXgaWSB1Gvc9B94Zr8xHWYvXS3Yo2in98iiVsrSf1RUePWKa7hVSyhM66u+GP8
6zam55ovJA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
paoR3khjnzY7oR+WJ9YkW1A7ZzfFLvvVEXiP81AieLlGnfQuqZTzy9TqIBQ7d7KWJF2u8/GBJ9gB
S/XHVoSTyo6Jte9XVVsqnnFiHxvEAnWbM2e9+Vyqd/Q/lFB3TCGyLNKIFNdGxyml1xea2Gq/DUf6
P6PVaPylNEwivSbuc64=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
IuseMdZSknnKUME+O/YmMG9MKbslcWjYg4y9t234jonRTsM/8uUOZLlJPdAz0Ojsb7gi8Afg71RU
Er0Jr7fpQJ8YMMDdLQ9qwRqf4zAR9ZhntG7zWMIroK9jxtC2bvBKKArJREVpkzOWU1g2+f7dJ4FH
ubSzqp/ur3VRiEL9rSTe80jSph04B3Z7vLg49YvLUGmYKlwP09xV4/46qike4zQtuofkQ8/u3jTv
rlLcM6RtgeLWfD/CY/EWIIuhTxeQiucCqPyYilV1cA55FNKfdMv57PsY4PVV/CwLFMYY9INUTcQ5
vlvEZIaCBXiBH5TWThAkm9erewSr/bL5DW9PTw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
cyY5ZPlO3Eo0cmsRtMR6yuz2Eu2e6S2W/D+8CcC8VsHPfbx1fHUAOMrMRz8rOeXuKPOa7h1hSFcJ
XZ1TcAU5VIvCkM11jW1o53hK8qachmkkZZnfj8JtjstmyVTyWri5LmUnPYRufwJmQUQ0xqMJytkR
VTqDp0ZVnyDWp2/qKN0=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
WAcKeockg4TPNpKWNqCVvf1P8zBdM0HIqALOQnRkxsC2RA2Dy+P+XMiOG7cG04xrgm5iFejfnqcO
5lDRzw1y2vm9IxrTgVR8u92CBfbBU5si2daX0ciu3+tUaMvbyjjRBHmWEJd/+ZgwpEBd4jKx2KQp
YmRUDFYL5WDDgF6aGgbY7bniF7p7fSFQgxz06UbHJt/aNGcXnfge+DPA60LgmbiAZYAbqv+bSmqg
gA91XQkI7oyEKtZ35D6ZzgJ25i0EzUAy/u4ctGTC1xnExC071TQUx8Fakynqcki4h3cwrvs6RbsQ
1XULS0sNZpYYdAavNOXALBW23U6uD7bNRcfAog==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 33936)
`protect data_block
/ufI8eRNu6YjfHZno4oDvXL7P5xQb9ErqwyhP/lkooHkuMepFJZsF81ylhOoOCgmghn3R3gW9+0t
ZIM+mAK4qHU2rieXc0KFb2M17M6CsmBKgo8mPKBdyhFEfwKxzz+28vu8u6ewBdTg+OxwtY4Z7eTP
J8WrgxJ/uxdimBNfP5snnJPi0/e7P/wCWedXGIK5rAx3qRVGdee3PSJmpx4TNQ8ued7CZOMKOesK
8Ive7inuC1gx4Od65SZ7O0nHvxiJ8JKnR/bm7iGrfSJ6B0lFzhjmPDByYovNUcYViocTSuVbI02F
U0cpJmDo6BOFrE4O6RmCbTHYHNoT/Mns6J+CxCQra4Gh8oDejo/6jEDf/4I2WVsPKBIlAdLhLc5Y
BKtNdaNL8tXMi4WZzYmez9wLikq59ihcgVEGpYe87dAsMst3QhB0IRAP0jBSTcRZHsCZN+yuFqcI
3MZ/HWYa9SxmblmXyZhYqN4z/5egIaQwZQJVrBUl9SpVXHpiY0EwQw40Cx9EeUqW1GYJNqp25xuJ
j8vgDcpW2zMngIZENEifpmQF1LJTymxawGepT3yD9HwbmCXImkeFypfPltHvffrcMNdpJKipibg4
4x4Yf60xV+GhSQxiso1cHGiCzcQc3896npv/U7Wt2lERsXrTUXH9h8YhahG/C7XSYRbXldPdLRka
YgZM6vPbEpt58I+/JUO+vO+G8MWbdwxcb3d6gpqJfZQljJo2iEd5KdtE+v78XKtbHE0lI8DqH+I6
Z5IsA9jiSD1QSyglsisqNgw+xuWY+DrcpBokTrt1vj/dD9G60D3sx5P9EzZx2lBwH2fV5xLGGNvF
Sksr30ydAWaR7VOjclhKKoBu5nIsMUjbSVq22Y6O3179jyyJnTd3HVLx2fxGBTGGKXEHJOgh8oUZ
quQuPWRlJNkiNNW1dbGeoBGtcyiE5K6PsZFak0B2MBJho1a/qzIIHnl+BvYsZ2n0lBDk67bvoPN0
rOvPXrZLQ/FDyE4Zl47txg6OZmkmweuDQhMKElC1mML1zVB9BVtXfY+BwUUv4PriQqv9HgAUcv6U
EGKzK6G7RfbdU/o315dIUl2QIIoAVUwWLFGd2JAZqsBR9obanlkByI1DkreE5mZqvjUv0LLpV+YW
zDyTklQIir0U1tIlQJuXLSsLAF4N891Oev8kYR6+X3bzq45H0gWqK9dujam8Hsa24U3QJcKmFKzA
yBF5X6OTOGNvXGTOtj05A0tmQyjJXHvvkt2Cjv74sqZFuLN0+3EAC42GRdYW3WWP2P0BPepjrTgh
ec/aGAKquPQq+0B+mNFh0/oFMrcF9DmUcjzWyqMKrM7b28n6MkfmYo5oG2m2yKFsprMEqOvPoPbC
8RH6hV+Zr3iDa3StyG5AWElXfXkL23zStLlzK5kH4QuzsXklTCY3HBNVFj0U/9k/N+zcTV3/Sp62
K4Mm9XrgFfdfxjwD/JbO7DJ0EchFJGLj3L6Ns5eb4GVgrJyU2O/EjJMTC4y7hFip7GAp0m9wAjvS
JiQ9OWT8CGu4dTE4LZeGgw6d3N0KjbM0hUBpRd84wxMb6llI+Ufnhkh/PBYwXSSh8iStZv39qyV/
6yqS13RxbsdlumU9rxDTZpce1uU2//JjGbAf5EgNbsavXZvjb1SicOmykoIX+skzssam/7O8gEOy
9JdKnFcxwjMkMz2l500IiOIfPIo+eUFQ95yX0NrHSHgvC0AAp8JtjWoq8HkYGbiighnwV5RtSfq+
td9RFbUvBogWPsvxvACP5mq3FyeyxSHQ5fqlgee6U0sylz4i2n6QolUc7ZUMIb/cFJQAC/+Nx+I/
k0GRB1MeBx2zdFbgWqSeyKf6fBkI/xvqutyD0sDvwOa4POG3pNEHnN37m/8CfTViQPdxwcde9SEy
PveSxJNglLtgiTrPgyOpeOTSu7MFaTnbAo0equCeFfPzPi7q+pugywIr8g/3FeQim8So3AkzA9ws
Wc4HsPt4iGi0//LkXrvQp5H4a3iMUDg1Z6KgXb0f51e9A3TncQjTnzmKHNEwh1n1ACWPTH0Q4g7K
tkK375n+U5VlMMJm1KR6Z9ZK5r/edefrPfx97t7BOO7qln4o9zQtUA4CBpGRyIJdKm9YLtAHjdG7
k6zRiLywl6z6h2fRHEzZjV1mqdTyecPYSdgExkeGJPW8PojbRxHexR27sExvS4hr9ZgIfCuc3k1z
b95NdLJZ53nrTyaSPRdA21U3+wyk1C0MhYIot3Nj0n6IKz74xM4GaOAepnfxaSabJXD+uLan5zYY
yGa+Bdf8HWRiF/iCHapZfWL7c8Lws+YcE0V4qXrElfewMVwRhH2o7Bb89fw3/oSXe1Mz7Fy6X2mE
R4Yb9jIzFmL3MKurAC51o7SHclkbO8DAf9gIYsN2rY3agGiZjhkwq63MnHOvq7lxAWxBVXZNF5CX
QkKdU0do3CW58USiHarfrNO+rh3Gh6uAvl6OfzREIQXNBrtuN4OYQ900IeUsLNli2nBrHcpzA+lZ
06N/Yr+HUwFh1lSlq9+HzZHb6Ud9Jlgjw0HNN67I+LadiVfMreGiK/OtIX+Zw+Nx2j/7vUyse7ga
3d42XstbDHnzO/sYmHTNDOUy1mNWpblUuB01WJTWnkrPiqXGPvI2BruwVIkO1T4WTpI4dyNohKM2
Xd8Ui/2Q7/l2pRes6X86pcIx7/DCOpNfb+/OM/976cbyQo1AokO9AYlpowb4Dwa8RoKI5lLq3BSL
mSBpTVtsyESULh8iIjTHi1JICpn5njKH5qu3idy8+zMMltlhfgX13dCalr59XRQsizuOQPH2WNAD
IOUBTLuSHzH4U0hjfBa3bR0Fcoxik+rX4Aryhsf4vcrv9sJUZ862qZJBQi7eI2hOFp193NOhHfYa
ZziCwt89TF7gTz4GPvnA+/pe6BpfSXGu3NxhO8xd2tJApuqHg/sv1dfj48cDD/jvoG9rorhF5sW6
EuiBLypSDpArXbg4nZDfnYv3+oxt2xDXigCu/32Q8VVz8HN88hRpvupqrYlo8cQm8XagOrUgKYAy
jJu09ae1/VzT3OiWD4nQwjYlmhD5RkHVlS75MnAFLDQX5DEoTO7kVrpu5mm5S8JqF2n/dCNN6EEU
VmdqIyQvOFNzA7m8TN6gq4IB6X6yz9heJClG5VqlaK3ewnlddeclEg9MeEnnIyisehzxG/D+lEur
+fwBsODhmaSwaDvwmxynPYQ4EgTY2ozkKSHBfUfRQQ6VjIp/6zcjAmP0iovR6GoeDBJ1Pfr62Pul
rNz9wZjrKsNEBwxDWw/2GmlWZs3TV1RTWx4MIcSuM5V9pBnj3JY95HEWc9xOkfuwmjBMnIWJSUKq
kpk+RpEyn+Oz/1pOau5Si9vaYrcUzyhL6eVOHzZbQkq1cYcEf4ioGRvvrb0K63kqDehkAlZM46s0
FI2H0U3Zg9i+m52LkUy04SC2lLr/6TxCnzQoVW+scV3w2VEKvFNvaC08yD502J72hP1Es/kUtvE+
KYVPw4NtU2p5Ve5w867udTf2sagv1Rqj8vtkThaYtoi3N2e2MMiSnUCkx0p56D2asGE1r/Yk6igJ
I7TFPdjn/tCie4ofPcE1mpoOM6l0mlOGJJoDdyQpPZEJpzxyP5NjxW2V4qk9DsyLiieqCzbmiYi6
EtjBOhkR1Vba5aIapM31qa0ELwbsr+DeIDynKimZB1zxKbROWoxRl1bZ5PTaV9ztsG8W+kZkwL+I
gQDWsPSMTgGTrk0rGIR3w4mlSeyzlOj58wRzONolwkT3mc06Ez9xn184w1VguIQ///an8vvEbr53
x/ReDncFGXbUlv8IGUKovKRTBUitwCBP8CCDfvLBusgYb44HaOfJRBECvaNF9JXwHdIPJhkO359t
bbSlZM3i50aAC78WLPnlplAkPSMOsCtraY8D1bMnrxGoqWj3c6Pd9YKe1fpMJlqxvdpXbiYJY1zw
+y1qT8B3CpMom+B+ykmnkaMPQnIQkjbGlXEYkFVYZyJOHSMOEEW+d0PRJHAx16qg1eMk1yK/06Ml
iHGzGB7eEC1Q6yDnGLUXWp4rpoEYqTgRtoeS3/iMeD3r/VNrWjZs8013hPkCceQeExlAdgXs+Mh+
xwhJCEO/rYlgq570D7xrm8dt7gGQAiTxOgjCRxiaz0G1QmKpHqnOVoO984cnw6/OIuoHNUl3hTVL
vL2WXUeAI6yiw8NxpMd2FhQ0EECkE5Knd7BZxy3orsECs7SLzYZ2+OpC06521sZoMbdmLCdC6gUd
dQGYTj/YwQ/X0uagCOqaAhwZNRSEQIEVC7AuM/waNYeB4Gc0MaAMDblUkwLC9v88QRrZS9N4+T9c
v8vENxUHN6PHo4gExPU3uSIZwgaIqrKNWsEtaGYv02jIr3CXJK241KI+CNWAIBscukbJXSMDIa3q
aH0U1xjeHTD1uMuqxgReG7AP1SxrVFjY2HpcggNsrzTfBpD0VMIhwQ8u2OpKAFAA/650yZj4OGd+
KMAr3jthVK6+oLgmxIPXC7elymrfAYcg+rblb2Dbxa/Awldt11hEGJFb6mAz2lY8GRQJHg4GSa5F
yeF2oS02NlwUylWYWBmXTnaAvmOmrwFgUoby4PxEEgaYu0MmPZAXBRLtclaZF5Tiw7HtyGq19xbP
DhzkDe1RNzZeWR77tjwvufDtueZ/OMQzmFjYvXAmcx+a4ZACkW2JrB4eUom2+1gI6OOp1o5fWy+B
G5KTk/JDIhS+ozDvnlColLH/20yKv50nhv0/kGK01KG3qT7HI5zqtaE7gtWBg3MbpmbnFkpwxVfE
weJuH9qSFDUxPZz8PFKG0r2Prfr9ptUlt3IUjCu7316Y5a3rTb+ZHX9m9g7i6IV5ASIvyBUpZy8g
G0I5f8AxbeAKpRCXMgk8cmwcJY2b8fHGN4SUGyKoZAJCQ+3xckwUq+zfY6mf/mmeALy3FKyfptVV
drSdx/PqePJpu0tO75VOJLYLuc3+DAafSs9RMQaijh9rFoiKI+4h6l4Wb+6j7CckDGpGBC2kDp9A
sy8PC6Mc5tsT2EfF2HI5TW2wo7YGWhr0ap6eeBI0TSmrG5t7SFmI4PNAtUX+W8CgdeN7L0ICkKzN
C7UpdPMNLPJlg9qf2S7Mp1V97fMkfQG9EBPNMDEr7lHsetAGUygC3ARdddqqH83oIgqCNbVhkcap
f40kwnNLJZXIywKgluNPimqIj1RmmU1G3m48qdaei75HGZEkuQGUPTNFp6F8WNDadNHUDGxA7P9F
NPpbXvU21RUBWVr20LM50Z6Vc0LuN1qwa1S/ralpOK2dklnCxLaxuJWwn6eQOXy127y64LA0yqTP
2EDC9eSmNmOsIm0zQ8nhDPeqi+KDNKRn+AqX5xDzgnMS0Zj9abjM2dCIWh8tcF39eexd3x1Mjzzt
cw016r7eK1Wz6Bi5cFIn2a9zc6zm/63sjhMCJo7sjAs9n6DQhVh+ddCzkUw6XrRmGS4uQHHVyvig
ChIQxg/OmXrfWjkMNsfUy/tc46d1xw8UOMiPzMjqwOhqR8GDKBxjwi/RzCU30gsoLXxhBchEYbPS
D125qYxOL981yBmE4tgKEFs6VTsm3WKjqC2ZzCAaBB93XOvAvhI9j/gsd6P7bfM1g0DBzdT3iGAw
qW0I2c6bJKSmYgB4FS9Z1yLYGgc2XlOxd9nx7XBt/5mONdDvH9YSLJ9s/OawngQXg2nLA/zkZVvx
wRUdlxRNJR8eVUVThML6jrrWCVIr90D3eBa1vrj4swjmg8QzNb992pcP8S3/Bhw/nQ2nR8LUhQi9
IKXDWMgYVQhb5RPk6Ocgj7QLgYkklTbI0R8/HtogRC2OHc3MZ9IbXfYzcKrYO5y+A1U3QA/IwE2R
ORlHL1yxHo9vu4t2PzksOEOZx1w3bF9jFMkQrivy1kn9mQlHSGt9vOGTmz1jh/oO2sYJSF9Q1SxK
xR3M0RMzSil83MIl6Ckpx572kkBpqgHHAot/fL7mafkk4PD2YKH3gT+9JslwDzgaUw3qEEHOyesm
Q9LIHcCOr+IohN/UTp2xkBkyABkdifaohsLyTPhUod6u7TxIhPhvsIH/75kGTAVVJ863vfEsD+QC
jKpBskf6OrU80E1JsK/86bJfVzI3w3kmsFGzgrKZRVCFbCuStPOeuzzwnoCTaEf2/OkahEqT8HT2
ThPJczLUKFtz3nbd1DGiCWh+mpqDjDJ4K+NRhm574adxbTS3MQMQCFXcsiovOTCXTRVlSOnF2TB2
508T5G8RFncqT/BZKOnU5MR4rOMLJKLCmLYWXI7VcV9c/IKvqt2/1frAhmeX1qyRSXH/+MU+3621
Diz7YoBkyTGd8gPiiULUyuXiccGZnhwKA7I1r1gPwuKdbN0pM5hcthbElaHRI8yv4yuXFaTcWE52
/csVbFDthUGF4kOIm5GYzg+LmMrrtDnQLXHFd9vPUU8DaBDfM2uSMIjkPGKbgSkRtufsqyARa68O
c2nDmeLUJNAOMowjiS7w6UoYscn3nRSkesCwMh0Fh0QHzR8mXJbT2BPWuWWbc701XcuWcH+NJ/Xi
OJmLplsPxdZrm0Zj+3JbbBNRiHCZXNUztU2mmhnWYNjSDlD/VJjWEKbEYiByd170yrxrT+6UucJd
hbp9J1ivNNWutthbJAUDwFV3H+Zua3hm8CJjthphhu3Wc2nYMXEDNP940dVELnJyUKhcUPx2d/H3
/G7c9XdFnd/87TZwpukKzOSBJBG3EwhwY+DB0UPJc/8w81OqLXTWzrCfkvkIyrGKWwkM4cgLXGNf
sJH2ZFxkoT7jNVOq/4APG3mkg/dTv/pcccTGlfJMasmqm6dq3bX9XGWxM4xL06+lD0z+YUuEragO
oUyRfzKVBtyejF37yanPiTmiGCGiX1acyG8dUdhKhd8e2g8CziqI22R0pcbhDzkk/pDTsLhflnrR
7mNxWSZnQCBfUG35av2uX9VeD3V3IijG3NIClDl282PkPSp+ZXWr8LVIdOvW4o+gbpZO8kIgNso7
Pu6Xbj8+3P7f6m1I07C1FXKwkgssQPjgcdK3Fe6zdDaZhyNmsFQqzvznEEK4KW4XbSGGMkLVYtjL
XfDJE50sSNRzgYY7bhEhSgens1TfUfxWmbnDRqg948XeRux2/7k5VNpp7dwomrYyn7qcAComcDNM
BpqV74FJJmcUCkVvcfrijPYyBKnCGO+55o+ecpwPkoclbWjDwguME/Eevsn7UbQpYMQYs/yayXlK
NqLk1+6em/uLXueNB8APiVgo1KcSp7aENP+Xpl1PQEmK6y/p1ArCb1NQ03e2mNWJ7RMS0Oa3vxId
YsdaCCyhf8PwqlLUSPT8PEMngTuI2cdsuI7UmqyOMZwI+AMYP5UUmjOJuyu3QhvMj8Ur819h2k3T
+l+5wv67dvS3d7z/XI4vxVrJyhJd7Y2kA35tT5d7fEtWF5/5NF4FqG2MWEf4tExWQYPc6HMDjnRw
oQn4EW/xCI2ny5A9fR90vItu7HIgNlOy5DoYe/oULZ9NSQxyWOCZzBLVAg8n0YeXeTQnKEunoVHq
Jb6VLoAPDmdeWgGSRRDyJyIK7i4+xTXGHMx9RafTjMZLkcuW5l9oYoCT3/U1vSl+WXOAXdB1TzqB
+9EIn7+dyZs0wJePbKLSlPxhDKgXMBy9yIFSKOxh4FBT/NYb7gL89XDOYiNFENKbwM5z4HxciguD
uQ6M6QEUfA32hB3HkFt+xGMU/zFH4Ja5GltXigMYgozYAXOe17SZZdNmJK1vtzofoGlEOGerlh+E
gSe6Wfa0xJ/QGUjiwHxv8CLAmUgvzeWTUtfsBzZYG2qXmZVxxbqwIBsfFwIjndY1ECFRrfB5aPex
SDypMt/jeqEfhf3t+2JQmhdw8IaDCVaR5srXNzLWAzVgCcjhonq42AOLRQXCps13ONRSTvMjrIF5
8tmEuo2x9kHcQ5npQskJWBT5KxE9NM0BWSsp0y4tikHcRqDC48ZjWn2Lc+EnK9cROKaNrf2XaGgK
GIpEMmcU0qPz/BgsB7AAE1CgTt9L7yUfYCkj2R34vr+OrhctTm+UHlObT+aDAv6G+OvVzyjQo7o2
FFR8pFmzf/fiWEK3bfHKx2rFYd4R8T2tFsB+wnrSv78MBw9xOrVDrllsWtPRHh61Ufom/nrCJMVH
Qs7tre+aTGAN82DWLffVaSNeTa0OTgJztS6fb0S3dLaYqvuw19kXg1Uzm12kbqTHDMOt0SaUDZmv
b6BrM5TCmtgxxwoAkt8MSKlNFAFGLBzS3tXZJhGFvtlUzcvLTSzQhZWp6Dm9boUy1ENMlC5DXgUD
UAZfYU37JbTAMcejKMSn9mX21iqfErQskQxe67H6OZU5ldnnl01WZz+S2+UgkNCdKkOncTjGSsNP
njlVohHXGOlp7mAdg59V14GH4GBKjRQkpQjiZOdrbUymE6uvwvgloGLlahcUnTB/0L1gPpC1baTo
Ycj2DH1B05ugUZwjAUAaL9Q5IbCE+F33zhc7WqzDZg6bgEDJFwM6o5ye+zMaS42DNI6PloCBwavL
B2UD5o8VgMHcyRfRsWl9Jb8M8mrOhV1mWOTo2yAFxn8+jX8DfQo+ORApDANuk9+cSeqqj1sHHOt2
LmQgIONwBvG50AMPDbMxmWF70CymZWMlHLobdByKyC+EWaTvWjrM99SpKhabgQwUTKX2O/sz/BzM
vhIRvsuUlYoumZOZ+86xJjOFas7YloUEi3k7C1uv8jrMhAC8C90rSZIgB+wTlDwBEVDA/FMpd7bQ
9Si3LmllCmo4uordpp/Ng3zETGutdGJun4mmRMD9Mw7R+Ge9TSTGGqoAhfxRg7NDlG/vrGxBojGm
rs1V0kdVM8WvIIbdmIG/OcS1nApL7Au7MFxBAuRHeBMhR1s8uWQQTfL0Q34GcWO1ZFqXjYAygmK+
EWINwbr1T9aiu6FRpvGIizEIElTj3v+KOf714yFHcaGCGRKYt6uvv6QKMLhzqXuCq7NEUbdrY1BZ
S3xlptsUF6Ej5jFNN7rLwGGNx74g3QFG/0DHuZ+LdXACPUNSBj7xum8CCwbuRnsX2Qf35cPy77nQ
zLggphb9DkdedOfTrNMGvlifRBA9CKdewCRIASN6k+YqTQXVGLrdGuxDGxoQb3kPzUIr/GidFZlM
hntvIiWwOA14pxN6cLgNdS9ctm8TXarpaaFrehBF6PjzDFVyimEH/RTmjde7mpYkbdjBaK+ZGkJP
nf2ce0YADlm6HqjBHn7ZX0ng14xp0LzFp7YCjhR0tgc5te76BygewLov8AUSz8dOli+MhdXO6ems
cK3KG3KWm9NfTn9Ysw/Css0hdJ9yHoBeOWvW/hp5X8DlGBxKWE+e9YC7QpeITNkr8AYp5gbJrrHb
X2E84dTqmgSDBfbo94dJEgp7zFI5wTx+rQE9EvuJmIDTH6bSg9J8anQjIQ9d7w9NAVio4LvBrdf5
ZurE+PweAQLrn0b45usFWGlbKLikh/IV9IVPGKHw1+kyIlDt6mJBI/qNAFWh+L4anMYX9Ll5RW10
Xrodb9vtkyfIhpxdR3Ft4wnnR29Vdl2WjdQzD9vMXMvaMMZvGmS0TG//KL7SnDeuekz2GaPlNKrB
XKraQY5SaN9uRIWsFAQcS6LPkWJSYEKfiSXYh6SVlQ5n+0rrpzMvjoz3dD9wyJ+oxcNs+kCpwWGC
bskumItiGLGzek3vuib0dkxG7c4xW5P3kcUyvPSKWeK4xxc0mof9Ruxbb9bxOAevSxunBnYcuA8p
3/fS8fczExr7erEdLTGFzjscsh/Y2gI2kkqiJqHhjjAeHwEE5qOFyN6Va/1+oAT+uGZVnWH/+/eA
MJ6iaUDPpMk1eluEFzGY/kOWpPNEj2eV3O+VRDFYzdxvH42M6XXinNoh993i4cuN+WnCeS0pZjX2
3VkNqlm9vVZ3NEv8EioLI1kV/lYvDOZsxdagtJk4YuM3TMxTW0Z3u+C1xYlqme6tOMCE/tJBFyUS
M9njULonFhSXsde0oXfVb9jA5soKbznOgiTbbLIbyIqkQhOqjA4FNZdNiGqXo/qAZvY0/AX5vE+X
syvyV/Hc9vw8TeWaX6VvDPvAiAKU9sDYyfUvDl45+h9gPWTrMpeTHsQiuI2hOQ5MzVjEIgEBW/yk
BwkPFeviwI4cnGqO2aleWEbC/OCG0yJ92Ph+DNgx4JdFtcNetxl+YOHWmVcXvB+/ACSqwh3xm9uh
po5lHD+TZZhT2xAuWBN9jqc1v0alIIJa2CQ7045ZoSi8TmMpJpO/WDVC2tQFwRdszujS2BXIlUpp
5Y7YtHHD4LdAbPkvAJ35kn1LfnF1pDUISedRUTeQGYzWcTRLhbM7bGRnFujYxl0BKbr4Fdd8vL8h
bEAEMoE5DKzdLwzt+nYyuAj9341lMbB1N0BvcAwPDj34I3Z710F6dlF7UBzMPsgp90DuDBBE+BO9
3Zo2D3OrQJWvmkDOijgm4ysvlRm/Fo26B5FKYNtK4ySX1FCKZ5fU8If0vTfTUNhlHGbDPiiHn2JS
ZDGrXZY6FDOW4I7LaVzYdh8UKC1W376SRheUPxubL1Dll/HIzrPXZ012CjO9QDUZtOc+aPCu3ziF
um7F+0DgEJbfH4vBf3FFOZ15q9XkaWLxgCEN/SCcMIXPpO1sbK/6OZVr0r88qlp+JWdA2aoCEzEj
Zq6QGRk6kagbymRgXPtUxhqLXnN4xAWT9FzM8b2uMQQ8zbZraHlEWsIHtcLTlI3QNT1yEUEgWFDt
HHK4/kBbQzFWk/KNOgPDNS2Zl9BT8TXTl8OYXkwoKmJhrMzw8AaZCOuXtOQ/va0vX+xc2PTDWMxl
IKvDvoYS4hra0C8vaphnq6FYuf2eorTB7OqmO8lrwWG+plPsZhFVIYmJn2MJuipZ5Dtwg1zjWKrT
hqrPdy56VQSgBuLk4TwO2e0nA0QSnTXvWqsyuy7KTfuLz3eae+BZn+bamFnKw6tpBOUZMexj8PgF
x7rpwZO0P8mp8tLFvvhzCmFZUH1kvgvR5JAJXGUQVqKVuJ4H9iOisbIXxKq8IaF2BrhXgmR+tZxu
8pgq2PLAP0ddybDHKI05ytQheLTW6ohWa3Bo9p+HKHcLslZG76Bvn2pBRW6Qahzd/THVB6SjF9/i
QJIQT+jdKmOlqq8YuMu4lCGD925E4d5Bvur3cdXItt5gfoZfefrj/ntLpGtVacHwTsYaioTI0BcF
PoZ5zXKxTvkpx5t40vI/XAw76PW/Ml7rmJzt//SnAwoFEuSXqHOg/MEo4OBGvnw6T5uoiOwuhgRy
T/a2+ESRdiFTr1RC02M8JvZlgHjFd9E4VIEfZ2I0EeqRnAclvQzJi1P4/T8A07o9Lsy/FSy93TKY
Qtgk0o+S7iXdwV56rPJSq/cb8JA+l0LbIDLPVpj6jHE0K//sRRpq4HfspNtNfus15JM5gS+O8CCC
48EI2lu3+SmmEasaJGdHiq0I7r9w6PP+x27m5/Y4+rblgc0dULJs33BluvSNbChYitiXr4F/h93m
Sfkh4TPalPGCH3YQ7rollMmCbSQaqJQfq+TFNwUVKgC/JRL3yrxEjyp91vb9FTGMItbttky7KIUk
gDpTihGC6j39XnVl+Ow6x6J8a7n7A01qTEe6OcqHjUu1Um7eynRwur6WH0FefhOLVOLq4wkLYxsM
joKDZucNBezrlsJ1qprP2bdkYFQsgDhLIqavWa4omRxv5w5NLOxEARFIArNdAnVf3UmKdKRDZGcQ
23Z6wgBW+pWoJE9S5iktsiKaYGVJJG8wOer30BXqPN2ZuJROOECI7qIkMIO9hsdU4WF7Di4KSFdc
gUZ7+kgjcJSP9mia80SkOJsSCPEKdDcatIs4v1zidvA+ULfWRUJJb9jfNlRRXGFzUYHWcB1e5v9s
Qy7m4HXWXXTKAne0+rhxyVvABNj0X1QpYTkVuS1FaSvdm0yygY0DdtIVeDkNDyjztaK9nz8CaKc2
DmuBf0Y0hX1LRWNHQLIrIpZvorMkbPI/UnkiaoOcqFV+0+JM0IorRRcNxzmmpjLeVngRzDtBUv7z
YlCst1JQCknXbsdLIMX48OQnsrpMWqDvWpKdvjjcjWvaittviYX/YHp9L75gjnrl0gZ18bR1HdV5
3EPAu866JM6GVvOENlOUbfH5MLUN4UllB2rfyBjJEAyxE2btesucx/0GZNDzxsJZV1uRH51KYXjH
s5TdXrV5a+LkuNGxWPIdYQjcdCWO75hznBUmstFkt0+swQSbt0DGWf6xPSYFXEJNCimJJKuXg4hT
TAJDaR42RKQ497VOQZrcCwaGusUajsvbw/gvWb0ADWBkRQ31a3od0S2lFIehXsd9OGZy+Mqgt4a9
B6COq+4Nk9ElymcsT5TGaggjeSiN0AeretiZJ0tofjxi58YqA3dGLODVQ4XVukTl7DL4lK31+bBt
SzlTEwDTqXP9Z/IujCFijUaBUFjVH1U6eIK8iEY80kPe55t3FSfYyPGCJBlEYyf9OvrV/SOJc2gu
aCAHpG2abrI2Smx0Ip+0D22BdgrifSDCOfULI9H9+kyj2tEYSPKlMFQJRubC+DsgtT5SUTlKBiOc
cGq+/GkaLCe0tMRLIchafA9ZbleS8lo/0PKcJqQe9G3i78Gq44zKsJsbSKqQHwfjQi0WlpQv1OIG
92zSnfKd//65KFfJemlzGanv82mEdCyxxE3/wjYYPkNaBQIFl5p0HZyblG6+Hm4nRSqXMt5ZT/Ww
JLrKElDddTBV+Z7pp9KcQC9ig6uCoXukGKuFv+N+tsLIxeZEGKWjwSCd5juhoIoWaFy8dVryoXy1
/ZSHgWismDjV3hlsldTCoY6ar/uI+G2DrduT6LPc2DiAk5vOjFNfPovi0Wp48poJi/GlXXnZeU/m
NJUmRaaDlcbbwFqLWHgAWUp4G5UiTvEXN6j5xbbXET1cDYWmgvIDNG4FrrbkU5l08BkFKkWzsH8s
UzGxYrpVmoOc8CAMmO5NRqkGMoWjoYcAHU3z3byihoTvrO27BtbH86LgRxuTq85u3WYW8t5smO9b
veOk8yh9drSOKwVCghckWzFWr9UmTRCPTqsStdaKw7hVNMWkVIapU2Dph911SyrO0UDoe8/racdw
xcYKZT9hw3Zj+iOeHi6GoSAqLt3DGYvGdoR7e5VQjmWoEky6yWegmoQ9qn7ZKh4fX2QEzghlhg54
q48S+KWmtdbZwT+CJPqRmqNh/tcpzSOdC4rATSe8atb64H5/oljoHxeXJj3XBl8XwUeBPaLnQxJM
GCbkwWGid6+hLaL8fQJFbU+4ZkP9J2Njm8ajs1g5vXax/imK96vw7VLQIvSvL2JC7yxDC0DjB06j
jFH1Tstq9BPyXJX1qcy14A9iFbWD6Loy+SCNDCb21/WpfS3DTdjk1lco3bITIDLRafQXlRUHVnr7
voHqcuRnQRQsPazUOFUIDtH2SUv71k/ak8y/5R96ewlFh++kdSzZOboZTRKDMy5sFPlsIgdZy/qT
J8F2RFcyNBsGVg5pqf6U66VcQqnh+ETcNwMN7QpFqjj3IklWWroIGHviDYTOgsyiBIZNk0qB7+me
DmT1Arkl/qePyAm7wzGcpVMW1w6Gh4PAybGvQ+pnntIZHsDCbVnTGkY/L4zzQYdBkTyiukLZJMYl
ap6qFvHwwr5ECb8QfWByoQnn6kEFgSUhYH8n19X2nai8RlN2YSu4t14jee1EgA+1Ui5mPqmYAidC
4AZxxyLK0hmj/i814YyOtRpLmttCG6/mXZFTl7uUyuha/XxRm145If0UGqXnPbcawlo2N1cJ1RFr
xnflIZhw8alLQXr3kLLR7q/uRJHfcbLH13Otsr69uY0nBEPwCPEBbMiJZUdkdnyDnFVE485K/1ql
ZAId1hD3lvc1+s4QTCjDOHfcCrB6lBzqM0lj6inDI9eJ1r2+cOb5Pua2CE4j4iNxZQclgTYmi2TN
KaYbXVNHOcX4J/Aa3DmMfeoH6mu0Cah3gsLW/JZbQB9EBiQjL2jlllaYcJJdCNaY5MbyixoSwBXl
T8BkkbNWsMAs0OgSPrgF3wG+PdpUZ8iLRnZuDuu2QZzqr+5DuYOo21RdiO7texyMU5KZiG0ewHsv
jw9iBzerGlrDG5zXaWIR0b+x9LHiK1qjOl3RpGOcjceLW/e7SHr2KxqGU6B0DcuvjvB+YLPOqSfg
FhbqZ/KcDVNwRTr4SmmEMGetsBqleLdxiILtwN5zk19uHS+DhxNpscuMWPNf+rerlfgjNbJ0UTl2
FOcZr7cfH+wGSSfeU6T3P5PyLbUl4p8doPTD2UhWOWRZ2Mm/mfRb7vEPFVmTY4K7Akn2VnSDfZCw
vGsNN3seZTY1jOvvCKE8sczlDbydaanqzbFOZHt8Kk9Q8SSr8K5+7JmQBGFenobrUzVverLnZ0Ey
F4UD0UviOshi8mvFmwW+Y8tTydKmiw2pGGJUZBJv4WJ09n39ul8CyRbRCLVE3kxZEC6nDeVvoy6U
DH0u2mKBuRIMk3rruVzpsSQA053tgkFQsosYpGBuNrnGqnGtby9n3Et8XhFobT9kj2g9Zl3erNQy
AJNSeVF80i1gILJuZhnWjym5npAQICodQBq58Mw2xvqoRjEllCDoLW1zacSx68D9GUCzz5FP7D1L
8Kuz+vXv6//cLFJTTPvr6SDMQ3hCEMPE8aLy4mvp4POWwKxvtmohjM/93S3xitRBOMGsCyqv9QIZ
7h+PDm6w4UH8VMmqXkO2wQj7W20CaFTlKTUTwNjm1950rEmT5PX38H/rz+l+oEuSQBhxTp13Gw9i
QiPTkH9aWGckspboEfKAKwV27al2hwx6Nfv/7fSHAlF8EIoaZiRvKRa2J0f/sQc1mdzANZDPcPOS
83Z0giT5P9Jtmk9+3hjscwqSinlfKGHJyohPM8sACGimTT7Ve40Yef4o/mB6hx13xNkuAitOEiki
t7/nBIT64FL+HzrT8INIw+hmoQwW2OmpZDH4mdeweZ7C5IASS4VMFaOc7zqT2eqruQMS0HLLJDNo
zbwwMPwpJ5eliDEBQIdGbGMf/sRkliWIlKaOwCCof31/ZXuM3vi/9IapbcO/ucHRpk69xpebmKvU
w+wsSc0Ayw//WbNRDybpkR/5LOwJUoM6kBEZgtgBU1wODdAyR3EDmF1XshPOPZHBt8mVlguUthJw
MgCtMzJP4LaxkPUGKPPFo6NCQbTUZE+G7pvlkwa1e4QDN+7PgrlklUgE5XDUScristjVbgNO3Who
XE5cpFvekoG7QKcTXFW+VkGfx1O36EtmS4Dn3lnMreKC3nMeD4zs21EUEyJwjZuyqqpAyCB2nK3f
cPQun6WRCEQgv1lkRaaIUciu7AoSORwFwML2OcAEG1VxdDhPocMGIHc2Kht+cVx8BQ4jUQVdvkjP
EWyi6IfxWojR8AuVFIeHJxM1C4GFMGoOx1HER20NUb0cyYwlA51EdP1J/XMbv2ygvww29RWFyQSs
j9cOXl/gFRY/Ep1Ye1xLcmYK55z9VIHf/eh+xFJGHQ/kB6Tdrwik6DevH5snaY9a/VKn0WuUcTvl
2hY5F0pKzn1TzI/XJtzk+DjBjan0/Cn1xmCU5UDnR9PbBSQ8eTevE0Ovd38oH20mTBxVS2JeCiKJ
bhO5v22d6Matn6w9kb7C9CFjxbg7zP3ne6soTgap4Qb8JcmmpHuon1MTKVPNtQaVJusjumd+2bNH
IVrlMqbxHqi4fISU1So2UEIuXJcSMxV2cMVdHi4mv3K9lft8uVb5CSeOZy8GgmHSuEQOCBt82faj
AzVBFTd5UzREsaNnNVrHKgZREV0pzBYaT5zU+nKe8bj6OH/hCaoesc7Wh9uMdfxxnCWFThwXsvkm
S+OjDzRNZtafcmxgcJGQhHAplHYpGOY8cnYpSr4+xg275CIxUBzghcRmOI2ggFdOqK3D0DLXVTWP
KlyGk+HMH6A1KwpM7hW9ce5ZO9rc9xAkZqmFelRHKKM9kvQb79ESNtHl4rmJSrU4o2H+c8sxfabj
xVCrtDacq4xAQhgdLbLbQFzToSqclr3H9yMfaVtxV24zFyjWmH0w3GmbckQxxZ19atZ+7trySYnb
pi45QgefuNBrqfZ9qjuYvhwxBTL4DHorPRkQbwfWpM0de083tJlSbTDL4TKrQArTpWtBSafGCr7B
8kYAmeITX6JH6tHnwslb5BufDpp4MjCm7VdxjjP7vcT22O9GxCK+SLFmQmgUofRb2VRIQNXs7uY4
KWdYncphvc0cueYvm3LUYO6bFsj36T9gZVfS8FJjvV6QYbFPTagqdXue1FW05IvI0ERlThXlGMRn
d3vxUAKOYUfmRVE8f0+7wNVmJRsYsPyn4++BqSuDcjih0U/f/uxa8PFMVvnNrRw9PV4pOJLZaUJL
utCAgEIrcl7sjvN+FRXGqWV4BF7bST0J4uZqiwATYT/v3fab+RhaHcpaqqJl0/TUBAVnTYh2MXyX
vnormCuKeYVRGes0dNeTnBXy20pUYl0u9y1KMUGpVE1Xs1657PGLe8u2fmGT0FMNyU/eM9KGUBQY
k/qqkYN63qJehSLtiGJWUY6VtJHST5voFcCvbjrM9Yem6b6WREeSVcfZUXNYUzaNvgEwWRemrbtP
7Zu/ulLV9AYhwzJ9TimS598BUzMdUPyM3HXi611/5kn1VXuwzHizvHOXRNXDchYFhHlNnguDZ9Gp
ie0IhD4lswFJbmSAQWyGnIRZK4aaMPUfVN4xM+oh+177yVx8a9sOGeHnVfLErby87dpF8nKcA6MQ
2Wwxl7+ubomvoZR9AqhcUNcCxTQASQKyz98I/e4kkH3fH/IM0ACBtLA+Ms8zn2Mq2AQyIBxwRPiK
Q8H81xxqPMtCLjNJdorKgJjfLBa6xqEcxkOPYWY0T0XYLIHHUAuA2EqkZEWVylYj2DFat+eM/ESn
dYpHi+qxYe3IdqIxAA1E+LsLNroCg8R7QTsAt6SX7I6jYlEjcUpbg47czaftCmKXg+RsbMw67AhG
HjpYchr9M/1CG9DWNW9Lb0gsD3tFdYME1R6SoFNkP5vvWY7cHZfeErA8HOvRWp+wHOXwKaIan+pI
S3OaYTVbqVIsqn/uV9j6Bf+FyLhsZsu3G6Wo2Rox74mJhlW7UuKSi0qPbVU304FdDJZL07w8QdmH
MPF1URv2PGcKns3JhSYx6V3DNKX1PzGSEjpdfyN15gfhEc3KMoymQct4GjysuYgUGxCCdhAIlfJt
KyMKDDLCOe5nn32hMiUjGofZ+4b1c1YamJ+a7VwuxFs/ZlrHlU0recFVmWdyb7CYQ/Tv3OpNva/2
yoD1zsUV4f/zeArKoannxOu2GzRVuBbAcbsUyhEVeisW9XzCGIB1qD8FV/keiNlPWvOVoMesQ3at
nwEA998OrWzWKmt0+FDJ0v8cwLafQekeCJde0unj2+CXGXhCNbyzC5OiYw7UffuHp4E2W3C4V9zi
M0xPUM+SdKlKaLhBKyYnwCKn5PLjefeN2VxD2MoYyL0HvrHRWwJZPx29CIZolXk9hFu/Iq+bPJua
+Dal3icYJRIQ3ki7Ljp9K/+n2qfzjKfZ0HlXdSTCNybOjmnK1NsrvcgCgpq/zWL7CgyBAS5QwI3y
mg28t6qlIXN2w9z7HObmgWnAceBT+nhNidh3QPaC4dZAwcBVzvyny43DZU0y1BYBFQbA0mYfuggs
d8YfEH8jpqy7Rm2GnCTyo69O8q/VoLuwzwB/XayR4yjm1ZNRFV14F3Uf8hKzrLkXdQotC1Lkguo2
S/oqFlQ7XZ6Kt39yg79wCpcVS3Eb4CLYjNqzKdn/h4TtM60aRtEpsRthD0kJP1ASDwW/m+sRUsbK
5KEW2Ui9ZGgEWKrLzaLmzCPG9EMvYfqu2w88jMdInw4izMB7d4SSEwrze09viBoqV97aMaPTAOFC
OP5CGgi+ndgxv2MHlaIfyfubfhr2sAZP14yqvT+O6QVAXR3bdyM4eXV4gLSyQ8r/Fc5Ib4r4nQs+
m2CaIFBnz3XpXjGcE5ixmI/t8+zQmSwunSAO9+xvMpU9BK2O7lirnBuhlWbZjQgZecIqCAK4CNVV
Ra2yZF0JPyFgvYpEH+6tD5nu+IZLNspLuzcO7mvYQtKpSwkvSUOXWmGeg5VaFJh6wiPhQG8PCCNj
UL7AEaVJ9OfNzPtJgO7fGPoKtnLycKT79kBTP1+jo2f5H1fWb0lOvlNR+S5yrWVN5Pexh7dQcbg5
vbuPS8DwUkg8jrUfj86HWpaNy1HdlJTKzh0pRLezMcPjDWVlOHgu2XOjEjCYgbYN8JvRBGpCNVYH
8U8HxfNXdNNoIX+T2vBB8R8+06siu+iZjX4E8++urNgCDd4yiOpy+3I/TM5y5uUoh2qDBWqSniAs
bH7EiDE4lK7TnkC7+svv2do30huH6DM4+NEkK5U0ROMLkkL6e1Hcqj2vg8W1Vq+CeNQL5hB0cGtF
3zseYsOcHHvBe9q/31YkDekKYcD9wi3XlE8WGvrzcAfEoQBvPP0HqUERKkjLz531kkopvuxwkZRa
f0KII1+bS75X7UO0BOrmAlVWFgK0fKbeFKqOJ1vsteXZQWGV/DLb0QfJnexQhx7wGmc4yiEJmow5
3NcVGFLJsGWWpllG9+KfJ5ZBpXDYpMNxAuH/+sHXYYuDgg16S19cjZo+cjZOewNdCIyEKkshCOx6
/tIwmTqKiIsA331SK1h6OX61NCZAiiwVhYkUs6tLBjMTxRz2QhzJXyPoFVnZyTF5g629vP8qzSGY
sj3VD5r4zNS8EZUX+/xv2QdpTrqlrnLXz2TdUdPDkkHtaM/n+wvpU2qMiBfmSt8gL5sQykfsC85j
YjT05K0/4ttMW+m4jhoFc7U1pVvmVM/xN5cEaCygd29zQHTj6iV3cc89VJdqBwt2sS0SyDpp3Q8o
rfgqSipp0uH8jUupXnGWvIUJIbibOcLLTXzRxOiL2uPlbrhm9P6SZokbcpXu6xCf8id2tNfyJt12
Ltwr8YiBXBrCJC7YvsFqCqQPOQh8VFa3CD5oTINhgZjP48CpH72a41z5A9GamV+Sem9i4+2G41mq
l3w4XOAwyITpOfV8uaoXK4tWFC/R/rKUuqUM1iIgqTU+Bwh3pHPO1pc5hGM0Pp0nJOteBCfOwB8Y
Zlq7d1Qc8jhJUvtSQ7JF6ZDoCsmhqMbiRXG2TTRBMi8NvsFHleXU8AtY1OicIyLFyMSJyjwdM6qr
9NHKqrDtpc76fEXL707Z2BGpIIHC4iYO99XRkOu4d3nxwadkNZqEUPf+SAsgZWhd0jjrRng5m+p/
0yfflO6lLA+6I/c08oGtXoMcltneUzL7ky/HS+cYMjl4O0LUn4WiZT96MznCxmuidHutOoxqUVgI
NgHNa9gE/ggH+2oh5dJPquY+34Y7GdWfSXco5eTKMMTzwB2Zy1slmatADyegaezQfZVRcyNN9WwN
S7GEmM7sxdah7IRC4dK8JjOzfXESv/iafBB0+tsygnivWu9CrORltyFX+zFTnpFsElMK5/fZhYdY
k/D0E7Ri/jaRsAZeRK8TQWLX6sgb6EhyR8ECXR/62SLCNFDEtcXg2WfqbPz7e922CK3sJyX+G1EA
sQVNZdOxmXlzaxFov+UGUNtWMDXtk/I/6cBWrEcua72lOtHZwoI0DdyPd0BjqXMkRnyDHzbEc09Y
Mw+8iLXAfpvgKy//6C39RcWLoZl4MwJHFw41ZYycCw4gH1Nd57vV3IXvdbhWUUrHi0MObL+iHhk5
olZqT3fhxpiqFjx0WgXiqWl7Ek3AF2fW1+UreAiT+4O4L3ZZ1cN7CsBaOzGmiIQM7JXjqabP8n6n
3BMcM1wngv/65tTp6Jzf1Rto9SR6WFKkgwD4XmJ70Lk1CNcwImzhL4K1hvzx30YmYLYveLcuKo2/
zM/hURMVQ2oYclE2UUEGZSnrLllZXsGo9mEZLGFpOh3N9VYc/s5Yd/McWS7YvNBKNTL/T8Z1Nqd1
2drNVNRqAY5MTG0OrtpYoxItYUC6DFSdEHJS3qBKevPFHhskfOQ/7Mr7cHuz60I3uwj96foDBR75
vGphlCFydLYKN38c27ssBNqhhSDFJcnl0IzSEKzUahO6Msh26k+McXI9UcrGlZx9EM8VGuv7rfh6
0tRe2qt3ygVNji9ySkmePFMtIaC7SkDpHOIwX5JcNqz+Tm1UJoXKLtpz9aNMEBYWufJHOKUb4a4b
LpEIGxnca6N1DnIM9hc2uURaEDEo0pEPGjQNhoAQqGwTXv0Td4PgbN/oeoXS0paZ6MbEu5uqCNLT
BXkrNldfDYagQHxmLfijS6j+qMpi435z+0lHFJ4zugoXGIRt7E2Q4EKxwULCeKBpcQfxKyEvul7r
uS774VON3vwuTqb1hypd+ErcvExx81+NvLvpikwdANCzOjX5aw93Tf0yZryk7Oi2ntopK3GrWUqM
fYHVoYgdsY/TFNjo/xXZvQCcf9iI5cO4eotOjV/JjDFJ3WaG9Ns8tnlgzthhhpGk8zbgKtLz7bBF
JInDJ/SULddvmTRGqs0a1KKDWZPPbK7vIykTO/lcQLTtnRFIYY20Fm8BfC33i+41VHlp7P1LuN+U
Ke2BJwmK7JcNO75sOMeP0IhcNSDodZTXkAhX3bk0qDcFE+agbbyDc0Ub/sXM0nuav5AI5D0bSqWb
Xu/I9pPXra2dqt9zIYbYH6DfwAg6BmPcbm7UbgIt/JS68FBPi315b9UNgI5LITYWih6tbQ0UCA3/
eN0fFmc5OlEDj0lt0DeongGBK9VX7z2uiQLlkAGJl5rTcQXoduchce2CIYxTySfGSJI4+J7LvD8n
GHrmc3vwKubSFO8/lmdBwlp87CRRiR69YfYv23k6p537ILaAut390sInZhpeOhX49CP19rF8+KSV
vVvbwUvqU9/6aNGZdYImCY1UOkVTbR1+bh502KRQwBte6NGUZ5DJ4R6Oy6HUxdzStMVEZPP7X/J8
5QLnWz4BUAhst8uzkGmC4QmNAbflH068+GZFSUuweGwqVaNw+HYK2omqoy9tW5o5UrlzNCDWjylj
TUGnbruZn9hp2lEEPXS5AzLAFMitQGMAXz/4TdUAEo1aJ+vhVBm9A/jqTPk6/0RbSwIAywqxbcC/
x0D/myGs6IiIGvm24hxbEsMuStfS8Q8tJ2nK8kzrh3P+CVDFKpZWeEyAOL7vYzhz0sw6HSZ1aFdW
f0uyTHxpXki/SWbDzzV0jHNqxO6VKjXEuqs5GFq3P7DxcyGjr8/Zd7OdYm2wsCwVlHaEgq39lr7C
rHVl47l/jGHCTCDH2hWH8SjoHsDFWt0iUKbOu0cce4w4f43B2E7grSK8Z4gxuKw7IMoDY3KzRQwk
FjO17QQDBXIM26p41XpnfD08/MYEg6J9I/dfaVCyqS4+lwuXsRVjFe58z5FzAsShsckEKk6rL2Ed
uB5wZQ4gMjnahPZYSoWlMk3XsiTmxO2Z5EaKdRfGSriPjdAhpG/Onwk0jg4NXArm91UPG2VHvwjU
Bd1sxOF7/LkdrLNuzkiDYYXYhz2aodunwoST2RhsBSfEM5doWa1OwmMyJV5znCqdAV/+x17TpIns
hwRJfVVXvXJJq3E+4NEfY3BcAcjYpRLvSkkTpMTnkGMz2QJgkJjXgNwdkJjKRYt02FsjUX0tCUNC
YoROnLws7BCMTHkXEKym62CxdViG8ZkxsAt3dzJ4PBj2XqmJSYOVRRpfpiLZDcYePdrhZDEykFrH
Sysl2I1491pIpGgWfSztedTC2pK9anNd5GqbN/hHXAgQPYpQpvU4o0TskvZ7o4VO4DXbTcLe0LEx
KctK1XTp4VxvnghA/ts3RJ1/tagSClGLB3l3k0MwowVMelAEisOBaarr2aXk5MO7vPytd6Jm9v6d
zYrVKYCxs/2LFdJEPFN01j6ym4f4asghIfWBWFA4A7xaGqppcOWCvB9p/Ysu9v5XyRDbfr+dcZej
PH+3Gmuz6apGsP4LdZqQaEdiJg4Ms/whuDCFofOcF60qVUp9KfIIK0JMVwV760AcAWgK36LGs9a4
emgZX42DeGz3UblrNxYCTzD5YEB9u+2jamJFsGtxYw0TQKFCwyjQQ48T8ZceErrwa0NWkPcZYSay
QueKeG9jXeWh71FIcTBj1BtRSmiN+OMoMcBalXNk9XQSjjKCWNDyp7vmP1xfNT+tqrb+QmavZwXa
krIh7BJTtuOAEC4ONhjKcb4O6eQHIHENdcyUfYZhfVFtV2v2e3J4WAeBvoEasAaqll/phmNJgTPT
uZGFoT+2DaeVkpHkw12P1ffthhY8Al1Mzhk4yTOKL+Zq2FOBYXV6Cd1jwNKunfjzsqhXPE/9InbN
p9ri0cKZXrBcrSoGAOh1ZCpF1ksPZt3ZZJlVkLmI5n9xdrIM/2ZPcFTaR1nEoHt73tMZArScrvF1
GQ8Za13HvBjmh3rEz1SL7AoiLsW7VxRlsO8ZoGcaLh/SzpQVgGj3uwWZQTj0IapEvZb3aliVaLpJ
FauZDAF9jsIf4tfIrXH9OW9NG9HOS8r53tiR/Lhf1U26+MylpGg+B5FsCE7aOOb3jO5KIzM4kSMX
TvMmOdIcCZFpUX25TcY+xlMZtzWW7jKxIYjJ0d3ct4xt5qzskFnRylFfUKfEWK117MORThv66+gg
7ifbXrNh12N7dbiMfzT9YpalRnoo1ZXUZX+CDO6jwxAyr0LkpWVWI/FqIoktXwwPNMhPR3R0sSO9
etauW3LDhj6zmrjUDoeesha09iyoVujN3NG5nEnxg9BRosz+bPt9H16SSq8sPU7JAgO5KvD0RZKA
EXCHNZnRtiABLg49nQ766wZSBE9GdABBn0iYofTkCZ/IRV1z8lumB8sM8ixiLZ0iPqSL00QtBIlQ
xjbW+66SG4U0j8u+1eg48XSwJ/ZcrJXnAVnhLWq1cETamlxU5sMHmssdjJnuVmIBycBe+DzyC0Nr
ae4Eas3UIw7iPx7wifvdyjGsyYat6/iKh76KCOZHQFcGX5Mi7Oj/m5OFRxhX0q/3JiVUpcupudsG
tJ06rGzNwa1kwIUbf1nfDOZAHyfcBJt5nhsm8Z74C3a/ae+SIOba9goIdud8CUHVdnLcYP86zxjG
dsmFCFqblf5Xh9DiJRB3rGwuWghx+XEl6qXF00EdV6ei+OxKgbLFbHdBlxMPQVjYg+lCw2ZireU/
1qVeycj7SvJgIArxzw2EwB5xqTJDiSj/IgEmHSyDfvsk/bjOUI0sydF8qdmPVdJBtuhlU+jbpV9p
78cY6PiqDbSD07KBArHHo+AFWeXJOL+jO6SIRVYA/4l3pAd2HJuZozofBgp/tv1C7UJmmxNriokC
9Seq8Ok9mgDx596Lr0+FGGikUT4+7W2Z0kI3OTD8T8Bn0yupvWMJ1rIQpv5NT0HwKdujqV/Ag3H5
WiuRG8EKycsIRj5vlHPxq/4zm/QMBIrOSBOf+VUNIqx/6yHoHeqUbOEibX9ibv2K5RwIZcgr6c6I
zFLYvajZKmlsyvrfk9bPRf97egmsmNuEre09bqdDldSP5A4Wv90wT6wJpRvA3wMnMBOpVj2jA1Ea
sgujTVggTCafXf/IQBDz5nWWIt/6qIHDjELofdSe31zmJq/l+zSOCyP3MaE+D2M3Re5kuJzdWCfs
nT9oQ2uRuMUIIe+mrpF2qMnY2DYlUOqK1qw7AeQUm3c55CDhV5c8TKnkK4XA8JiYWgs4E3BohcX/
pECnIm1wAVbjOv8p2INd4noCDLYFYTdjzbhjvQnyr5dprCxqtwUUdFRn3yuvhak/NBnckJnpIsgZ
J0V5gA8e3jUpsyoyCYc+gQxNbylI2lVtEd1gUnDexuM/lF3v+qxK618LlBM6RBngU0yq5f56XPnI
rzRkVmZb/mZIMk3D4/gzvIxt81eG+/A3pCK71Stwmib4MEKOPYXpKbFzu0vjOXA+qs4H9b/dj4Wv
jv93Q6UvNZN3ESW3bMCltQAMi6FxM+uri65+xUB9sy/Hj4ess50xiiGxLLvk5bEGKZ5PTwye6Vmz
svo1gOOvn9zNsy2zkfXO2ed1oB+oIcXN92rB9QX8Ila4rfwev1yiRcrIzVOVo44CGSK8emhbPBMU
5W/62Hf0aalMg8XsT3s31e3V4s2X1/TNir0U9v3LQmsPWz+KFBcUHsflXAw5sgX0PdXz2kPSSZYB
HmF6Q1wX2gPOsYBBUwjdIzD6u0kRfphOYfTo6vZaa6mY6FYiq9NHku/I04+UA5DKzjDG4tqubb+e
wiD35Q1ZeyaZ95sUupsUO1mFu+Sd8PSXlFRhg5uco6oSdMtq0sGAGgHZWNCYXg1OyAyF/4Tycnhu
roif3PZxZPBQtCarNlghZyLrAZSjF1KFhwz9+5QOowyOfAFsgQdFFAAwNOSwuez59ocaVbyyHHHO
PNXwFjVhLTeJRRnVXOAsXwh1JICswQ8G3R+WMMme2j72a/bhDasIQJQVEIhzLNiPwxQyxpwFgWzm
bBPE9U9g6o6o5dSZWx0n2j662gW8UyCMfAdEzTi0LummIfcBZyBa9hqFkTOQ2no5NmTulv2xOIm+
wa9ceN0FDGIvkG5OBgs5l1Ayaasv8vJbMbK/1ufvyJjNxJEfdjwhDxD7U87xXCVoDrZo/f4edTqt
UGLAbU1IJ0sdrroflGx/5tD7/6DxzNHQekk2y3SQIryGZJ+CBFKJa63MV5BrQ1t52f3CeRtVJpuk
vdamMDSAzzXAkKX9sseROv4ziy1LCCYvOel5EzDiPfLRMRlns8QyNdUVYlp+freE3xZYxEzR/HYb
2fTGzDyv7tGUZMAJW38IYde191iFJu891+T17A9IK1GxgEV4JwRx6OMuPKEWgHk2B3YdqgivbrsG
kX6JuutwJZbdigfaETjB2pziQETGMtx8BPeXiS+ihddX2hVu0wTnw5m555sr9umciQn9TVrXhGFq
6tUsk79Dsbl0KUILdUXMbLbMm2YjuAA1wISTpiih83Hw05iTch31qQg2t6vUxszsMuq690awPvR4
9Rlx/Z8mW3vn8zIEv5mngUd3auxYp9Ow9zddk8U5AehTsZ5OTJ2QGjnt4RuiaigzimpkipxgR/07
9/2DhaJkn4P+4jNAicjK2ioeShVAfvQUiNLkepFR+YfgcvFr37IjXLG7LM7/3VPVjhKI77SxTI7g
z2/3pyn5iJWTRcM4AsQ9PcH4XB4B3VChjNacDclz4/hDrmExGUHs1RbjowJqxdpNHk1lk0cyy7aO
miG1HNGtCaiqoRJZYgtajEgjnttJfRT12ZnAIfNKyuZElDNwSB7yjsw6C8VCajF1Xu3Fmun6zUFE
okrgmFA3xcz5L48YMU5NENS0BTFGmmhcklyQ51MVpCVkpzxgB00zSw11OkaqzEFk+gudjXuKb0Rv
ZSzFGqyJ6sznDYFcZxr/slk1EsmpKzwUGZFbB/L8DN6VoRCL+Cl9H/w5Ph6KL7JoHVe7lQov50xR
Vj8UQck+AXBtNXdF8bdfRxSapAxgodyrRF/4llqMl0VtzwEpZvhokLep9A2/CeLtNB6DR83dIZZv
69n6SBXFCRBtrWSLRVjcTWMajXO4mCrkDkXa06wMDYRcBsqx+LSCHaEDMAdFxlgZW52DeqCSANf0
qokeTmnGtu0GWA5Uq+DmGRkV2as1jfV7DHqbg2zejVJOqvVDKsra17AhtaIJvF4mUxG/cQ2BVqZP
vBbNvKE4V67mf0BVWqKUC6IHc98iP7oTmn9g6b0LAT/E5vDOxzsBPvRLF7qf75Q41zwuzYQawqB5
SrVfBHR8IAP3iLFt+1n2b8wptQXC2CdOgQIJ4QM4iiC1PeYzAbVHHweyEaFDFFAKN4klaOzKszrx
CijvxKtDJ/EuUr4OSOhqpoJ7PHS7t+SCeBo6SrvHFQKIwgwnpPCWkb12awqZPIKwxUTnaiZG/JqI
pNB51myemcyr4BqoX0+NBvrytXXC2Evti4Ymz7Fr+8Okp7J7UqBTBclSrLmcRy7vw3ZSq/sD/ByP
ao22xh1Qecw9XsGxqJesNMevlUfiXJ0MYQAbN9VwOq3GPDXCgYVj3s/ajZH23Apm4EXnKCgSzs8Y
Byv8F2V6wGImLhhfeeDVwPQKfoO/Ed+YGNMWhnwj7TRZnfVOnSNIP9SAJFBg9bgnJP14hR6xW1pZ
3iv/4mF6gWDoDA8mB5GSkO7ortlTGY2alUETgnlLF4MlLJNTvQnSiSUug+G9qERKQeZZ4/GXjy5h
YRCzHfbn66R4uwehNueDQt66FMgLC2ujuDg5VPnxtSsly23j5VjpWTO/Lg/kLhIzQcfP564lvum4
CURaScS0ZaUvCv5FhkNT7CKLLNg3lesiaygnmJ8b/d9LxJXNtggA0rFBzclEPYt1M5E/recfOc2k
1VXYnL0Eogc18RAPX7oDqQASGYxgS0iF2gOJQ95wOcClxCWAOEwRami1UyFEEqQsrxEWrsL5iElq
YlC9xfz9OrieRPWaMJ2xQ4/tPjysmGC3BRX13wdSCEhG6RmNA91lVHi1kWHy9PXq8VDHI695vT7h
ccGvt0UeJfIXEjV6QvUoCKO3LGZamvIDO+8tzRu92OTofqoG0SMY7m+sq/6sWawVOUnLXg56H/33
nH49pbuUvTRbYC9p+/yE41Bt9yasalQLdKNqYN6TTUxKDA3eN+fSifA7i6szDHHqbQ9JmYIjWI16
z5OrGoor2fFDVEnrWIIcueE/ouapcX1zUFOpbTves60by9jXqF8A/R/sBFlqkaR/emKWUOMMxUhi
NC6gz9N4mPO/ClMeP71EkBL3tZCqq9Ndssi0lU6SXKivdXyo8VoI/Yw11WuetptanvIabzzYRGyT
D6qIJQy/nlnyR6lt7TZ0U5kyOwPVGXiVzm2lGRZ+ufxsmGcvxykNQOT4RNcXv7VtJ+kXh4NBi8fq
eG1N9qzY1dwb9pVbUFE9L5IsZlPL6Ynf3dbz6Lq+A/UMeJTFQ7Tl+oNmLBbY2KnX+2vbSXx5OK01
0aqujTt0aM9vqAfP1ZBenEecen7BoCJH8Tr6C24GZSLwK9MH+R5ROsfPYbkVPiUAzGwWYxfUW3NV
uLxrxRXSbb1TG4hARdf4m6qcF4DHpC2vfO0VZs2gbU2AoxhgKa+7mDrhdya20eQ6+7ZrhqvxK6Lg
rnvS8i4dNIGzj+PrpASQ6u8FjJFYBRvitCZs6Pu/qMR4EQAP+NpkH0V6zVCo8kA9sxJ1f15M8MWY
0tMwIomnyONzGyypKEzgUQMpA/yt3tz14dZ7K5yxgqpCbtZAIH5ZggVi/U1jkDDaSU3oPnvrBfFQ
z3qhKYVt2RHojNtrIVD1TJvPQIqDS47wzRZvW2QSMKxQuQ5qk0zug+zstr36yRXI2d/MQsa6suAY
LqhgWP6FHjo8u//GYtBe1oF+yxVKbIsZYFk2AhGTXQXdRDL3L7lOIhXSO5JXUWrwCEJWxymQarRQ
H5e0L/SCsgzTErMO8t3PxbDLzBy+EejKnh5H0THh+WbW+kkcMN7fxtueLC09coghEs+8OPqBOemH
IIG1nqBZAoHNwAA0ke9q+vpgaI5TSPvzj3TEUtFPHv9zvpW9dX1wJIsmL5dm98OfhyU9SdgCXTyw
Qj0NyVeZFY7MhbdyBHq0/CLkHFMjl56Y9gSxiBYs/UFiePCT/dQBwnpo381mF/wv46IiLykjKl0w
mLMiHC7s94TNQEs8qJGl2EqqsZnJPkGzq7NAYChLfHrFEQomKyEBa+sv1T4cltOewh9pb1cHaytu
Z4Q+ydA106vvpT5d/CTGrDUIhPBibbMBKmpg2MQ8Kuj4EcftX4mzYKXxPaD4k3LLA5kTt4USXN3i
MqXy/WD9vqlsH5AStJZ1/fV26hemVIysvm+DY+ELRZsrWQugdU7WWuWcL8VXnlETRKYfo+6vVvF1
NSgM7Nh9byQbPTdad6dmS99gbaHQ55H8Ar0qkZXV1/rT6yVGUcJtBEBzWBjp9Dgqeq8mzPRViViF
MQ3qWv3e+faXIyZ/a1jAQ4GVW79URlMLx/BceWSryzu0DxFaB4lEDukeYuB4AVm1kAkvRoreLCZH
Yw32QIbpiXeOv7xpcWz7g9kbMK5Ma7tQCK2ipq3dxBZQ6rDHNA3GwvNZiG6xY35Hr00TrVJCDFeg
mEKjQasHEKVahfyj6G6D4vsXHiWuVkd2Kw1cXfTy/4xe2o7fBBnZmj8pFb33hP50sPJf4Nns+DE9
8F90SB7x4nr24zKvpTtGdXPY2qlKucTt+N5YkxQ3iLCO5nZFGllFE8s+x0GPW88R+bsfeKbm25I5
qf8lYasVPYi2ePQQp3KmDOyzXFXS+rqgWJ8T7Sr38GQtW/rqVccr5x0HcFjraRGwqNJnvwzZWjHz
WrgmSMOqeVpUy11aNk3W2CVq23lYT75SxJ4YN+q92EWmnLvmSKCdb84zQWMoaAh59Nqg89PuBmph
32wCgXopKzPxqCpSY0m3TAKxvGYHylo1cY2HNe4qAxd4Iv6/DN1ESq0vu8emBsIAUoZnolyv5bSS
IfHhA14qxlMSxA0LbmjDs2bzVddF7mBGX6lBP4Xxu5DiMPe4kwbyogKzdUC+8yqrJ8BYxdSX2XJr
1tWnZ5dk6lvm1kWiPR1mUfmfjguMJTxQjygWoSweEc3TzdhFIazIEpgYvwwMiUBkohUYElhtEbad
EKexvivbYt2PZa4I4Srb8lbFhTXE7zXBpsyeUBhKqAcTjnCNJfMNoYN4XzY8hotnr1SC6YaGUeJi
tJ0Hrn8ZPSbdG8IwvxxwXDMvTcbYRDcayUmz7B2QWhhjyfe74vwF1Ru9DuiSxPzlcYlfxWc/9Qwb
8lKtZ6mxeBQWZ0S003JtwPln7rT2C8YivIH2Gd1m3wd6t26vhxDVNnupFgvTf6XRQssdkCvZ88mC
I9FTTzzS9Z30qvVcCya/P8hMpn6XLkz4xzcxIJ6dFGXkinT8fGAD0uZD0N2ezK4P0Fgx9w4irWL5
IfKevedmDWgJiUwS5DZ16nQ0Ok8NRNqY9vMJN5OrbA3LPJ6JBf4kNWLyZyO5GmUaisdJcpdj6zz0
vqlafe4XWJD5pqMPYBVYTBkWL1JKlRRnVGxD3qH5i/c84hOZYy7jdO+8y9//E8MRcQ3HnQfjbOHf
chYz2dAzdYQ4nUuvUqeTu/oEJ72Hft1Rw7Vtk1PBaMAB+jQ5KxTghywMcd2Z/uRiS2aN3d5BPpQo
DX1QRrrfHOtZMm0WHwbR1ouziecGvA9KGbpU724UjHnV9qqM7Y+rWYUqxSmDVl+bLLSeZPYxe0MY
vN/WOBzq4gtW8nrWssQsmkK0O/Emcu39lw+vhsyZOKzplksdEWPsNO0xTmAHwRb738qV/HR9Nac4
LY0R5kWzcHScZ9htU4q0NaA5QLJQfVUT7rBQ9dYGA2mTXxC3QmjQgl+TRcv7x5aB/WKGCjW+ZW5R
2250o7gN+ompfnYUK1irLPh+v7HHSJaKsl9UnpcMj+0M6RzCH001TlvKEThuUDIM6wIFEqJTbu38
WHEd6B6vJ4AGCk77qnV/girhEqj84Ut5YlI1QeBPfPf0gIcc+kLszdJ+FWn7hgPelL4x3rzonwFE
UTOTnItTCTwHgVsgMEVxnksGM1X0yL9nt0sA4fLodZfthpkyK/tTrEveDsX9q+No70uk+O3DQ9xu
621mOWQ9kYJhCCmva1JaqNGvjgk8C1MzWZjcJUy432SRIVPSZDi150JDGuMWGPFft73Do/krWv/C
m25jZkPqUeIdWnUiY2aH8ipr75Vcl21WNvBvTQNWv89dxdfDHo9+QB+HdulhZK5A0nsjpV3eqkiL
r/avqWsOLXEfGY7b09X7JWTOUV4aVs845uodZvmJnM3lrwif4RgmOrc2xXuJ4M+98I1nwWfi2RI/
f5XOGbsuojQzM1NKCyro0QaOYOW5ptiqE0IWQJr375uPsmGSkd7YF7VU5u28S+qDV6qI3dqkb3hV
aFvZyla0CO4u0jNLm92IGNVLGG+n9BYR/VpaqctqHCZ+E0S5GBJY2fbu/zAuU4O11ZxUy0aSNoRR
rjznF1qVR1FKEVD0LNt296sgLLDBBKH1mCBdBGbCUEh3qGYzwJDbmDfHrDC8gtMYuTmrpSl7hDmx
FNXxA8Y8CEZO/3xIfHqWQKgoPw+ibdOoLEzTkw62V8p/q1UjAC/5FFI1/wxne6IqiUTYnbqJcgOc
+ix5e5+qsxCVwvCu4gviB/cxIxVGESjgb5ZFaP9yfFG4VHNtUbWZLWwAlLeuMCe7SIHtzw0Cx1xd
fpssN98qUgfdFSHJgIn8RTvwiExoLu428/a76ZXUKHbVK8GlmNKXtcYQV7f3oIZiCCkUoJEqFmGC
O/DVqrLyT2GQhI5mrTmPIAFNM2y6qH2J1fF9EjtQtMgrjiTTLS1rDShLooHEgjEUY2QYlHjnxkyT
71J79o9Qs7DjJfzWK/+KRkOMpj4rzmIUZdsN02VF7QZj1xaghWuuhp4zZMXaN2jSpNE+OaPy5tEu
XBzhYlw/M/GqeNQ0UY6NZ0qit2Q+I6oazB0PTlhh+KNtzqPtgF890pvl4PVdaD7TNE/4ovTxmRsQ
93fbFef+/ndXno+gnTyAB4/+OtH6g2R+s7yM48X34LuT9et878Waq5efeeCk0m9dZ+Sk+Ln3AmrJ
lpD3+uBbY22ra4+uQumcvWkkbgyVjyjdvrkhW1CUr5BThgBdkbSN0MUN17x3+KXeS28ZyMzolxvh
gOZEXr8tbVxIocbv8S5udeMunreGnQJ235nbhVcFux9RjVbm7ewpNgN3WklH80r9D81awjjnIC0f
3ZTkKrnR6/a5e2tMwRMi2MDwMe9mknaEhYIxpCUPzDyScfe4oRzC15kUb6ONPgPins5J6tUhoGCA
A2SVN+3xZ+FaVdtU+8yFwjeE5hNESmcLndo/QJda3mOK1W8HFJ0fjPJB5GL8o8y5HbB2XSQTAop0
GvtfcXiagdC0YWrKmFkYjXqgohtu6cC2i/cWxQlznrKKfPTyV8F7mqvF++lNoypUJ1P8SElc+qRG
g+zhuk4ocBzn9W0z1ScubqjQZn6d1HgkbC0GV4xgkEliz27j1dy6i0zXSezsNbF4iWw6mt4RckZb
eCjijxYPcymQ/EFpdLkrl0EIYieLx8DeuMRBeFFVil5NnkxcW4t4uOePNkt/MlSWmpjJ0ys96eab
TG+gzBJE0q6u76R9jA+zxxyOTN45zDYpGNGa8yz9X2v6CS/amnrYo26brAETa46gdvUU5J2Ev7xR
GoMsvrpIsmC4Gxhjoeurr58f3y/Qtliabl+nYnK1n8cj7AqAUUhW7IboVS81mVLok8QlTaM5PdpC
1CsqLtn+1uH30LZPqGfeQdZXIaoluymeHD51Zk6H76NdKOI9mtF/on8F6P8EA5qzdXVWl8vVAQnx
2vCNv3QjvcWrQMO/0jhca/xb+axU2d09oBVJkiTQNc3b6D0Ou2+QUb/HJTi4uCswm3IVsfXewqxP
6ao6JjHMEQAj/yB58PckHxv8BHMRsQiRFe1NATuPiMzdoXTDB0urikvhfxj99KQTLYGR2CcODDR3
THtWcXdpiRoLGwJgsg24UdvZ7T5eHqO/ko9JSZTelVfWAz4jiPx0pjRkuobfNyV+3HlnAef4L82v
69BNCBDvNhkt8/23gQI+GeUN26vtB9ClBQB8bZnGQ2Af8h3nQWMWGUhJfsTKW7dmu5qAu/DFde4w
9zpSqtTaUsx9zBC7sDoVSMF3q4xolTm3aa+LtO03RnDGyZ1PcGVZalQd7N7ozyb6wmIjAfFMvAiL
6iOU8XKII/xY/K7Kp/19gMEJNJJ2jdNrEuMCB5RcgRIqSYr+X4BKVpjvzDXoX2g73n4iKLnJ5gwE
RZ3MXKAOO7QR/tLEwMfvqy6mRG1XIKzR9hn1waECi12KKEJwk4AdwDEPlvrv/WEnFWvIrM4ifFGN
107NvPUbnCsg7A41XgCeWKN+vHI2dRqaqUprcegIx1Xt1LI0D82QeczY7Rhb0TbnBKrQL8oPQB+9
HqydWXuIpFj6cAxfLamb9dFabYIlupzPT8StZ5BHw4kHyS3CXbOquf7WvIjRk/GoB5YarBTutjJF
7Hs4FPuYafpnJ76fRNzxZZCYVSseKJybmjkc04NYWa+DwTJm4hAvotic7piBv2VbnO1J+EiqFNgm
EGvq5tKMTxFN45wS1BAZp5qovoe7FnhTGISCE0VhrkDYH1+yFkT2r6VGUCQJeqhZDeysVZC4E9C1
WMPmyoiF8X3bOe17Ih2dvA0cFMLEjBfgqKz5kO7FXN5U987YNHtBoksEhvfyNu/MrohJEAG3SlQu
/VhdF6kpgRVbMfXm3WOXiokGOJVLmS9Nuf+F4cvkyixuXJqrpjzyXWMiejL/YuI8eB8k0YM1rsXg
EPk4ep+SyYyNULLFBT3es8Rk0O0j/s9ESpxv7lMoT6DiCPeWNdVfBESL42f/C68tJFr67nrujtmm
S64Zu9Ocvn0xLWiN3rVEZ+2qVhklwdjUrjJaLkTHwNgVRHQjWYJyIWLRdIJW1H0TW8h4momXFneX
Wix0NOjN0YviqwtTVhlMQ/ify0lIyRcxdiQ8TaK5q8cUKZnEaF7o7gjxhdpaECnyWxtXnA5cfitW
yX6eQhNQAKc9GGuRdoPemOIKCeel6oFTP/485kjBPSnT8NFpzLUFMLREhJ/QvfGd2nlKvMWTTeX5
8bs8ABpK3hf65hEkPRJBD+I4XA+XlifMDHNrKQj70MNdA4p/j77ut+n+gIwnP4LRLjQgoOb/+sbP
68uPNhvsrruR4XeDsDBV8T1UctetREEzWx8L0kDNoHoAFB899Dq8R6HTL2liudmWhlRK4fxuGItx
jtjh+dLCsVNWo5MW3fy/jyNk7yMbgpU/akOhvnyS0djOXmKYNGJ+YTDwmyvtg8APritwsufFqXeT
8dR2X559soxcTL9D2iKOR+nzyotnsbgBM8/gTrdqaTw22tB06USwXwoj4tz7eaeIvxVkTOlsCnJW
ihIiQKKahNmgo6XMM6c9cxq+YWiXI95hrBA+IwyJsImipehVfNff/vtv0BByycY45PYLBhuZF0pb
c0ZlovzGAtnSoP4kGclSxw820vozqtBfKBNGPq6R3mnuXPPnHrA8jv/tOjk2A1r5mjcu1eKd2H5/
PhgqJ7on1Bfuh7iTgroPcfjDykarjRyfwe2z6jvb0YlOyUMolZ9/5bv7SuzKR9kHKUU6K/oVQObp
wTM1l6fV1WhoH3tb/IGMhApJReuJvEQb43p/XfhuVMsM+TSgEI07lfD5Umj/a4qDl7trExHAXjZJ
ow8EdAL8NL692Ayz+KbWVXr20tluaJbhil5+h4Wam4lq3pRCRrdBwvGW2jqIukVwWWsMybI7dnbl
u8Uo3ynWQUGqqVmlGRORLcvGcE9i5e2Uoyk18gjIgm9iSsDb8mQa8cPi+F/sHm9dLxO/5KjgCJyc
JdTppnnDZnJiyFp00lPocxP7qv+AS6ZlTTSBU7FCjVI5+/NdxPC1tpkbLcO546JoRMXyWDmk+zIP
2XEBTkYVlmTPBU7FQm1E4eZmwVoJXyBnR/yjALIyMNB729rug2X0IZMCFPF7mln6kGQvWYakR5XJ
Zt/7X92C3PIbrco/nacvHR7Xwv9lX97jqrzU8ZvhbquMjyhIDhKA5GS0UgmXs8nuOFBZjrncilhn
2tsqIOUfI9DVABF2z81Mj2hZlghlaj7HFAKPLaLReRrFP3PoAniE3VWd1iuuopoW09Hl3LyjGkRW
TN9p7LVvzcpBh/wGDPjzMMwYiGxaXoQG37DydM0a81xOeoZb3EZ/hrzH94Lv0I3MZbCLtsywUxRT
nUQ6Cfp+gC3DswFy5aW3sqDUjCatdKY/vbX21jZQA57UmpsXdPRH80xTQdHPLKCPM/6EgT4HoYAJ
tX+Y47eCdsTUjqtC0ETyV1S8Ad8fzDe7p4hOfUM9kHoecKA86UKAkuoAvl3DEaMoybv+sNbZL9qY
ePLB7ndqugpR2VPaO9CY2J7S5OygZAIxAYOYNGTxb7zK6qcERFrrT/8bb8mo+6vIRkJZBIcIwBPt
qATQvCCkLXKhvERlqihQ65G4BviQGjjZt8uGvjl24KC2az+bkutB7Gik2fYYGZYYGLLT9Z1D83ZH
Z5bQxkkrYpR/Nn/6us85QR9PdX8px/6OvCvgxU35d7GFmSamMp+w1RkeppS5q0ihHenKN9WnjppS
eSSN3owr7uKUEv4p/prr3x86DTVEwks3ZrP63ffF7H4JtMjRi1UjfyQckRY1HD3FAKkpf31gF4PF
Umtq4N6dxClNXRADWKQU1CuKzAWYIh7bf/ORajbXDxDL7C02L4YH8LYW4FD8yyZpNRRaTjVs8NMG
36CXuBwWeipc9BLFpc01I3vHAbQIX8Z0yMdL8vcVLp8HOx1fHhtRcZPpNI01CmfHR+q0peGcJ215
RRgIDGASftOQowynq5fZ95ta+CHEmR27ObZsb1CVX4fwMJtDLjJl65d5DmtwKljkENyT3hCcAEjE
Ljf1TTKaWzCIgbQnLfxXQF6GpoP+8lLWaYnZobtR13AyS/wx9FaBmoaouHCNVeO1jWXZceXOhtgN
w6MYTOWgpKkk79tON79PZDZliZ4kdb2rlW2G+fmXPhAbv67OXdFRWJzsF4iQk8Ud11eXRqkzJpam
hzcFdtsHTvDbrQIZ8o9Joen3Z11NqRHXElL6/Zs3q7LYeZkvuOM9VrffMHMCaAEwhoxBZc9cpoXS
I1gTaS960xqO9BlNo8QrHiB/R/IwCm1qPryC9gamZzjYcHMy7crylWbcl+hrD1z+UknpNOZhSq9Y
U4c2WZ0+WjwQ4vWwc87zUANafQkxlxCzo1IfrUwfXbUAyasb3im61h7G5D95oB3G1bDRwgt71KMS
35pMIEOjnXzonznbkIXUjblOpjppd5dJsp4NeiBnvX2HckX/gPre/nNijvtWAtgCFf3tDkPwpnlU
azaiCSBYnnKyFVxL5nZYV1ZVyRcak2Ba3LoygJjwRthMEq/XK7ngnLjqjRm7tsJRO2NQjyN3MaBf
fBeel8Qk7FnPwG/xWV5XgqxAJE4ZAYG+RAHDlwYM1SnJhqYubFQyTB/v6OXgGJD1Od8xh1sLYFoF
v/8crckMiXOMJzBp3tl3OicxJAR+G5PJDbl5//R3P5kLhZs1t5z2vEkU6ceEgZJTuKQX/o9RrWlo
kT56YDYOVRIuZDnLJe+XC0A8rq75saUjoSwDZP3TI5gZD1kJssYPvS8X1SMRZaD3Vj91mY56JWLE
iw++cJHqV6dxYp9pazzFBXSrxobUzN6tgyiLgr1FjH1gJus9LJkCziMHKCfdMavofcaYUpihDQkG
Aa4P7y3xPEyv7KTJhOVh0QjvcqNdtdDeyKWIs7irY1vy9QUsAiPfiVZivqg/up7dsNJrRPmSLfQC
NE81lu3cBf0ai0CP27/XxLQeFjMKvtYhCW5+qcJ7lrnMFVscMBP6MaHLB7qCheyYIIJUdkdun6f4
Po+WTgfSn6swFfntn0ZmSPXnaK2If6YDm/xYJS7XbdpKBMqYLyHaJ4DTOpWwuwqY9nuczP2gDtd6
TxTcbfiOfoCv6oQcS8t7eM7m2TjRoAxqGSNwI3Jmy+oL4SdunzlQpHBLp6SkdJr2u3TuJcyUW3FF
wRI9kEYqK8XVhguyRlUx/TxanFxb+ldk6g4IDYVzue5WLieyZwvf5og2O2QSjvcKsktHgbGmh90Q
iGgcamVWuR3tT+QFFuhAByqrkP/k7f+CxT1MEB1gZhrv/o/Q6a0F4HdFyytiF1OmnprmbPp+SWzX
WuIDuaUFCAqHtOf6CL6XkFoFi89kJmpO+iVdYPyQrjgUSbr7R6PGYazOZ6NuGatqE0wdypz0H8v8
fX7UEciluOKb8NsWHlNl3PxStoMSzFUFWiVFvMR81cl3qOGXkUi70vYTss5q3dx+6TpXbsTm+eXy
E85IXF8XJGG5cTyCJuaxqEQ8DHAfkoxr2t4ZZsMmxxx4Y2l14aSC/gLlHp3zHCWsUdGXda6g0QZt
067lW5+3lvoW5khzeGTm1Y5R5+toAaEtqedWx7yyWrIgiyAMHyl5dYJ/3hAcnsV/FHKnji15YpKw
AuH6idbo191cmiakOzFFFIp7x+PCAIc9t7JrH3q1r17OQqKrGNaAkkCe8jsU08yVTyYOOFM/RMet
lto0es2QhT2j8d36MJYAiWjxGGZhr5nLDunddCafWx8hXIMybX0XJl7wMvycocypaoVXIvrxxYvf
Mml7YkPdeotyNO6Ex0cxzVp+dHtLRdoZq9Wyo0ZFPwuHnd7Cg8dAMdEhsHc3qk/dKTKRWj1PeYjV
85g3KqNQTl4c2lw+GIsC18Acnh4C2/DhQ7EPV6DHfTczBWjME832yQ997CVNnlDBwPCOsW2HMvDu
pOE/4e8RfeFr76csfjgzbyMiZXUAHPLAWuMDyfzd/59yckqA/zMIigRC3rbR1KS9ghxW8YIp3Wsl
KzgGuo2rcYVc/LoKRlryiwjuNv3Z6Dk8KducnBD0kdRsMisfwq80IDRMm0qmdM5Qcjtmh+7ingue
G5nGh8hvUtCwmz+fKkDngob2432hSjcN3cXegDd9NN1pyZhd4O98RWfYolH/UOpdJxho2DLgLt9e
FMk/d4EcrB9SoYmZ0suK4eQp7VFUBnHE8VPdAy457TCYhcaYODhjK85UNhBrrPRJ8cmnR+4j8KGC
ibD3yqpqPzX9ALygYkJOsrw8z4JDEkBJkFBvsraPfyDkK96O+fW+VzmUNdoQcRQsZqXuaIMCdu58
VDscMeERQK7+NrOG8R8JntFp/nLPpoFWKZfPJTKnb8EWBSb7dPhntZHzPqn1j+uTIakOcnd7bCJE
Au3XqeRio4JJMddxCr7hD35uoaei8aD5QNpnyr6vtUOIDp1erqZaOMdKV90LdgTyYm6Ed0eq6NHz
poZ5ELr2c4CA2O7TpM1VuDBiNHflta6JRhzzjuD5uJWTH6HGcereGauuviynp4cce4xKcXN/GqVu
IVHJmd+83ftoDwcwrkBGRaPmIKU362zX2GXPCaGb5DaLU3rpLDq0ma+cslUZDtZ6BeTRCzROo1iw
vnlG7FYMsQ/gVogktRIzuJycLtjURv+fmXkSQurKugcQDA3P5jqhYvlfDtVrPrqvFrxOdAKJkmak
qHAcJvoWCNuJRncTLIDICYvz3L+UfUblxXDDwAjom6o7DhnZtxFYykVXm6qSBN07Vy0wbHbJaVzp
Cbc6V13g54Y+BqTD/JokuFGw+PpQm2pWShOXw7wvGGzQ4FfC1MK0Gp0u8kbWm8eyk0KXjkQuKmRT
WPlErmmhBDPtBDspVqmlGK3fNU6Spa2Y6ZIjyIOjVj3gfGn6fY9aZ5Wkx+aumTwxXEK3UOC1l3Ss
vu0jHA2w7tQfUWoQqzJi1u8SappnMDL4WbVGaq9WhEpLWC/tRo0Pikxu9LLhDgvORWz2xKdg/onM
3Nlk3/c6N0HWi2oiVucu1icxjWJg3TOv6z98OLlaPpfj48zZb/ieQMo+ZMSnW8BSwv/wT6m1NOFh
FtYQAQJNwjttJNQoFxuEnSfyy+BMuiCAjxaX1KLhoZxfBivB1JBCgv263FAPzMVijQmAcm2KxeYu
RdE8IZ+5t+XE6iSw4kL0f05DyeJa6ndr4+JDVenB8TEunE6xhXkKf9pM1jGnbm5zpbMm5vP6X27v
aSk5sNpgl/9j5RnYIxAMuFfMtJbriPprx8bPF5LjQXsbYUfND/lUUhafWlXC4VGjxmB4KSo73O+N
iyt1Z6W3eIl3zD+P8qBBJ5tb2oNAxX3og52boR8xNrFxIYO+gi1rkfQ2AmPM3tRLFrTDJKtRc74E
bqPy5w43Ctj8Vzib3iRVyi/nfJTj5qVQUjlVO/8lSM/NdCiO+uqle78A8RXZaIsGXv8PlsIyGusr
73CZrQdeZVmA0+aszYsoFtjHv9ZFendLQiu72HWwLjfGoW4Haw+LySpzKwauvH339MuBhTVsVoiY
oseIn2lt7MM3o6YnrHKKteo/+YrKQ5F8ehIjeBMmkNmF9u4XyQTfJ9ra0TF6P3PlevgUsYQWgDt+
TrrifYFjf2SQVWjyjNMBofwaZI2Tqc4Ah1i8Tz7lWKAWq+maEiYQckJFsCAfPKdlMha2D/GgPlBu
XaAOpk+ApS/8WmgZ2rDCZMiyDj6uL4WMOT6jJBbUj5lsLa0oytoR8faSnJg3tY8TOqJf0TSg7don
7RiFXoj0aYrczVTBoM63iqNmn42WhjaSZ/xivP8a/J9CrAFe0MqTCZD5yBwIamTMCgJT8R+S6C6n
rpXFOz9upLvwpkZKGn4L2AUB6A1GVJZ2wbZvPugtvRTXclWVzUWmI4md4MUBU4CQReqctFr4nyRW
YDc0QYe6hEj9VrGfVca/T0XdDqr+iXDEEdtdWYw1jCivW6tOVfkcYqgd7/eaooJqBw2+gAxTbSAa
tVNgM6BBh5depQeaLvgbJZ5uN3dn5BuyfyI1tKd447qYCNhErQA9qYnmMziv9ASFbZu26XxwlAp4
dDqB9+i2u1opmnH9ELUou4X2Y2HJTRG6rtQ5zTTElxp1Kj7hb+uIzicKRsgnOykxi/Jo6JNtSO/R
xR3XHQ2/KQWq+BXwjBTYgkAscptboNQlEyDjtdCoVnmuDDlt/hXMCzZUJ7qBrlVGomnAhvGunu/K
u8OaYG6VjF6uHROeXnddkRIB+STs6A1slJG7aTamFft1fLkVLg62RC9XDViOjpxQm5tSBblNVlDy
zsRW1NJAjM+NS6E4XxCk24YGmqc57FCbaGSehyGLzD32O64ep/q8F4TdkFkOKXvs3ex0B/yR8TTh
79GtITyCowwcOWhwBmXJ9VV6EdJX47oqt6GBthadxuWwwxDexbNd9yHlTEOiVUdINkmVWXAGrUZM
/E4kz7d0Fpta7NyeK2g5jlGIrAAvej+IPgE87I6DkjPXYK7HTMvuMURlttsu5aoHvnms9kGRyFvC
aduBr4oRjMGY7P2XBxrUJkMVtlm6w9xldEDzcjwRxxmdgPGSd3d18a51f4LX+Q6fmMiaWOIA4gyl
BARKkPeQv0kolPMU5Gi2830XCXaL4ITh+iCGYAqqhJW41BiBRshnyIhwOkd13tm5HBe8ulbVimbt
MGUUMBRHPFz02aBr9D5WzKLnZB3s8tZzGJhDhWtVsohVtU2haBlgU4gY1q5I9M6NEu4Qi+d/aHnY
A27NuvW/gl496DJk0FFLfUFq2UCDucs3lc/vAob91nGnulO4nzvJJmoi+tceKCp11YRw2NOL9GgA
TGfZfr5InnLrLa2lDzRya5dtHrs06xa3dZ/YpXmWkPgn/caUejZMJKyUPUuvVVnyMKlZEw6P0Ay2
3b7tRivOSJCGQcACohJSGuXPWswJc+Elknj813fBoY9cPtszbmchbbOepeHorhwr7BMlzCH1UUKr
V/s6d2fU0Dywt0UduvJBPGQ3Irxq34363n0eBhghsyQLsjq1Gn1UymiGC0r15cACJK3IuFZyVxrj
nLrbZSjma6Q71IqNxqtPOE+033Ug7Oe2Z6tmpmeuhYug8XZC6YUmukK648z/bo1dEonnzn0oENGm
ZYHdkPVMJyXYgWpqQx2g+ic6yIMimSJx236CipYSE1ufLKirA4dpSRP23wApVLozGKTHssyc5idS
WCnt7dQMPzy4AGGWJQnz5ElwuZEPDc+cTDH6JawmaQ8+lkOOuZ/eyxt4DY7jm+As17FotfAyZ6Do
4vURxZZ85aA+vbQtIwQ3SGaT0EMle/yIaDLAGO+upV70Z+jVXwDWB2vDE2gO2/8qycIAW62wGE6T
jOpoBasuwQrV5ftUbsgtu3Z9k9Qz+oBRuMLGL6zLWiGldXRcuBFW+NkegcUudviz5HYcweb367Kc
cwNqG483NizGZD/swnA+8aTFQ/kpXAEkBxD+dlxbepUCGfy0EXGnRuAAN7YS0vEVldWJCWzVf74U
MvwyoJdGqDR0Wfx0JRy8URkkq0iAhRaeOd0wyQ926qpuSxRGgpHRU7BjKOrSzuqS62ugRkj2qQvT
nrV8+po4144iSOBrunWIQfcPkRF0OnuWQ3wVdOOU5MJCewi7BceCcMR+l9iGrgaY8Lz8H8TGT2nz
sN3hFnH6UjSpCGjjt7X9q5iYwSf3tP9dNy33lQxjTV4tAW7Hgy/HlS0fIP97YYNlP3W2jnKKdC5r
LG6taO5694mrtBD499Gb3BdRDT9GR4gHCExGF4+C5QTtLbqC7UroJZr42dgw07MH+fOVqqf0M+B/
ao6WGdq5NA/gkzX9EjyGNhcBT46X8WPr9FKMGMhWfzwSTrjUOZxcL9UUCmumTlGuMwPou+bPHubj
81w4u+QbGDbsBrvpWCO9wpxKctQ0yyRefERRHHwwCEwR3h0hUDmL+SbE6vQxWAXyfMCZfsadiuNF
uNEloCanIEaNAuDb4wSX4NVmkr27/YQ/5yrnIh2VdhWMAE71PucS+7zv5tde0nhhtBQt0BM4k0t2
0h+M7NWNeblKCdhG9x9muozrrrsQCKejQy6CiW9Jm3bCYehtxzk+O8TVeu8sUtcoxrQzRsz8oLMI
8wyVSJ7XSmrJQx3shwPPS/4gW6SOLjSoICD+AcnlhXWRooy3uJKBNhjCoIjCUK1aSOnGSemvAkpK
VZW0NFCTX5pp5tLkEhzG8B478j1ZBtuHYzPhAGK0Jk6Lai+WY5YzmvQ6MnCG0xQ4Ar1Ky74w7tIT
Ym3Uz5WDnl0az/VS7bN7Ikvm9cuE93G3QP7ACbVh3pm6CPWtfZrKwxrlcpCmn/hJaJ1hwe8YuEhP
aMygLOO7EhGNMUSsWq5W5tbbq5YGaa3sKO/uu4yJPifXoJ+dxFWC8+B75CR2QlRcRIDvUqItKHMk
5HMzGAamyJ8LOvPHcl1ZOKSqFELk67LywZTKiItyrQrOLr6mdD0GAbUyXJNDxHkQJhnC2/UiWrHO
+9UzFIrqQQ2szKmca2XG1fTNQEVsMsavgUimvJrSSU/xB5SS+3k5nsr94+FAAXScyuIb2gwD8f7k
5NYJmHx8CEtTcOHGon2GfAK08ah+bT6A5SBTh89LfKMvPtqxbCWUXgrMsTu6a0Akn/3Zha92rcMj
BbEqR8t2nRr3He4EouADypN3C1L9yn9BG4uIXTB/+w/DzqdwJdVm1MHQ8RhBSEnryAf0Lnz0wHoR
AsK9nKh/aW08QtlaM8eH3EfgPN4jiXOSmBRcF5hRjAD20NcLRSV2VAoPkEUZVW5fivpiweH/rLMe
aM3Xlw17mHQufFwRpKWrGzQoq3br+9QQXo04nLiOTPftRSKjdY33Hcunhv7M0GZ8Gc9NgvA+eKII
tc9t7wXijZqoZpL/ddQak6C5nYfwjSylYyJQC9ReHvdoKYbru2P8z7phQgHX67DEzqbAfB/AVQub
SlIZp3vAy41svdI2+OpSJzRwTRLzIU+3OjlJNPH5Fhldq6Wy4ow8zaaKdTUyqxcJb/LwKfiQo3i/
EG354yJYcTE8TLgP9UTy/5L2MoGRvNQgsiA8Vmbcc7aVWS41J2ZOWtWRFlyfsOzVQfRl7All19Ym
s2O5YiV5uZ/XVo9SpssOA5wytBpIbyxn7iHEzhi+43a4L9h+MKUIFqrEjkwymTdF9jWfJ3rbIzvL
ek6mOUZp+JYHzTLA7TuWLp8ljs/42nXedb7vFZaVSL5ykIkCprtCzavCmVgblDmL1ct5mNOrbtDn
c8GO7Lf1Av3gzGhBzuvbPCbrZvpU+9PMvSeDczMUpU+npbtJ0Y5ENIQ5UKmM2GIl6q/IHsRLp0DD
GhP1zDorMhoOeXMc4QycdHNuY2U68zmvKZRy4H3HtELv9JJ2YimeThemivwFyr8No/eEPE/YJegU
OxLiMDhw6qO+OfdmF8CIlq4PHe74a1LsBIv9q5TbgrHdFgRtuOwpl3lS+WOoHEIMLvKFvVRuSI9m
KrAuguIzvEjyyGyKpXgcxpD+lJB03PbzmRf+TBXwhhz17rBgiCflL1mvifE2KtG0TH2PjFm1LXGn
cEsx3Y4fpXNs1lR/zkvzqs359wipMOoUrqL0PItpGJltlbGE7GRuHcVdPqTYlDCL+PR+8+xw5VNS
cJ+9ZsvB4IdqwvgkHQu/l12+FKm+r4mqjJs7DektHq7NsXAF9BXnccbDZ/qu65Ja0WZHkyVVOUde
hfADneZeB6iDDSjm7VwiAl5uG+izMMb38pk+LHFotskCuPGca1Sh2BpOechd3BfQbMiNUWmvhjHH
iSDSqA8dWNCvMWLT6gS3LqXMAxiGLIbRtCtrX2kCnYhUPvDHDkiTP6jJE4mDy8/L1ceVWvpsavfu
kfkIor6gCv5N5hnuCgZ8mMLjfmVs5s2ATCsyaAveq9SV2+SsmIWORcBwMlo+TV56OES3ik68aE4O
gia44seSQ0a9pEDx8lhKdHwAJzXGgY6YK+MYAIWlwn45Ot5d+nLjQfOBfQeHYsIpPAQdGBho52wx
DOP/tIosNnwPAz6+rdJumBladR8A0CnWIDGEky3Pkl9ZLDuvNwCBY/yUIa6AKqackUYW8QnCIts/
219DDYyN+vCRnnuGSvXaWVcI9QOkp4EVi9Y7smhtViNRuLen9HUknSVzntCgraM/MD8VIPIC8r7/
LfuiVAfAab9dNny2w8k3QFGqxXjAnmYV6PZfRrnBqNWox/cM/uUKd8DNVoSfppsad1myXTzh8lp1
n7RaWbcSKM6+EwAwbhP2jEGz2Al3+MoydDBcCu7AgqWHNRwilerkuSja9SIdgROSZMZI0DaZPEYW
mvMLsCA+EDX4kj/krSt4v+jf+VV+KAybY1Grsb31THX/+f9MRGuDX2QbHp1m0+Rm1p/YIs+1laXq
zquLbpvL5MBAexdlFk0i37+JbwZmoFDnhofLeONjW5kAr44uGIr0W1wAPNhjsEmBGaK/WRFYl77O
g7VN34Bx/gyOR60GNhOxZIDx+Tg7rmQUzd205UZH4YpkBkDW1+g+q53g8+DqyuOP35SitKZxWtxt
fK3MxswpL4m5bApQINbdypSoaqN5ca4qmubQjS0h9mxzEATJtWO0ZkzGxMdHIZkkf37IyaHILWmD
09SvYLSt16j78Z1hItulTLhXvAIpaDI6pIVGOyNbunmMfRETPoYLsP0DG03eERy4+wAOdFpebxc0
JCDXBIFn6Bv1bdiPTzYSahk6MnzYh6PgDB866JNpNp2Jd4sP2lNsVbx4sbVavpy7d2Rx0LguCY3g
lojwORoDuHMKosALKB6wgDQm3GDYYJA/YbyeCbPonVhKf3v5OkeYtF1aVDgeqhkgeVFRN9SQKGrU
rZa6UOdYTu083FcQpdadaUHXj2wAdPWkToKXtzzuROAVJdvi1HTlvIYrYsTmnzj1hXiCLGtUWRg2
9Lc9TnB/4EXh0l5rhn+OLOKmc8SCCGMfQZvaGT9+kX7pXLLt7I32vW0OmHI65HaEbaGrzi9sxsg4
AyfvKnolsObmRsUmX9OWOV7T7U5IaFogT3cuwy+JCOU2KH6R2XHzGzJY/cMHJF+m3sFplLCkgvQA
AKwEl/ndDyzeojimmR4piUPbVity4rSia9Faxj4m2us9sDRyOfJBLAn2fCwAv9JP5vjG5gLge/AP
5UWhSWDU2d/ihHzO+vHIZ5MaFLKxagHoiNp9apsGKdNjKTIdwAkkX/hWwpjLdj/Rfvux0Y0/jaJj
SF3x3zmO8i4x4wUIMLiEbDG8QgBGyfU1PzpyJI1650Mhq9IpZcqjHR42OZZw9VN43YvJokRdiaCZ
WlzvFx/nLJZLr38aEe2Z9MHjYtG4QppnIe88F7x3kw27pysizkq6A2rlze+zUwiG/X5+/NTJl+FS
ltGMHQV/OjbnmyH9heiUAB+BouX1Wyihz9J7lwILVdPE5evBTCUDXy+4v82hp+o4E7CNlENsoa/E
uGjqFrp4kWv9USmnk3HBVicKjBwGNZ3Wv/Y6n3oMlF7xs26URfvOLfXagfyJksl9VArQ/7q35Y2u
TbumUCWmKuKi3NFvmwWCxYqHRKRX0adNcIMRAK5TPprngHdgE0NttprkP9EkIHVhjNSPNci9kmAH
dvkuW74LbThRG0nEnGXKuZUZk+I4NAgRMk+XHHK6wok9+T87iSDtJMvJCAli+C7ihMLA7BIW3sbB
omudjZh75W251EyoKWtofeXNXCAaHaWy5ndUr1I7OG/gywzX0eW2J6EbUCzGHoWhmhP+Mb3hJC3u
EtufsTMs4kOqgMa+h17bDeqEF/ioispn3+HY14GQucpjvu1VZ0LP+rl3ZAUy3+aJcHZRQFyYAmmV
GJNsgrb1VsYZu8dwXewvs8h/e1mtjo1u1i7/dG3zoioueV+NP49TDq6FmmvP3xutFlLi3S/N10W8
6MUtngkKyKuWjFpoW9JUCkHDktzooUzBDoDsjDqt7sWEErBIoPrQ3PU8gq95a0GLlnBJXOhojprF
8VkLR4P3QKDXnxFMB14GZdEHDBLWvbnhTF6a5WcQ3lL7EChvlJDqgTqvccd68ggYuaIZhP4jKuRk
LHQGDakXpGH1hZEOWXnXUTVjXNOlwsKbue3jKW7eYtA2GSCcngNVPNHuZBlnvuB+uC3ljyf23dRf
EfyjAdxpNdm/7lLph51nKGMHdqD5H6OBwoSnm6bjwVjAN5SDQzbR15y81ZkGa+jlTah4q33/mvrU
Bdkvtgxq5Z4Pq3hk3mf+SAplhfjwRzt5PKrsSEY0Cm05dLAysmBIbxhQg9lNmUO2vBt/4cZvwffu
tVho4kRtNYmXnVrDYSR7pOpyewLSsvixlJ4Nx98GCB2+8K7leVAHtJXLTZRHb15jcFGW2KeVpBY9
jld1AtNKgV8F8pazEJb6Ijedn0ZMW2LMPXyF9TEPMCBmwMFtudFkh6DnZ7dlkG5g0tSUM8j8mHoY
3tPYQ8wDFAY16kvRQPbsUzi3DpgG03itLy2pFc8LjMO0DYMNbHLud9m+kDHfRKdZWoS2uYXmRyxJ
wM/1NjVMGT1w/Ea6FkCxkv1FdYRd3JdOCqC1cb79KpXkmH2qvE7QClZ4InMVUaSp08Wip+xvVki+
O4+29KM4D4XSIrcbFfF4qZbNJBmbZraJY8UF4/ODoi2IBD+1++lBMw7r/f06l/AuiXvnuCPCo74x
Uth1e18hKg4PwnUnvPeeQLWbW7kSZXqXpVVb1gM4SMT8u4Zc/D/I0H/YnZZYw3pBEv8DnLMcpv7b
Q3HJjWpzqiFHg3Mo9Vb8fXGPxyRx5kT/iSkQdEzen8WWEww6ErqEngFJqssfOZllwnEtiCuKZUT2
flSWTsgGxKgKa5RPfllFVfgmVpMb
`protect end_protected

