

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
CZom0vHERP+sM9B2H0IfoDUsJRy9riNTVWFr3BZpkrcd8N+2GrPBLGYjWv5bwWNFs2qiaRKQWIBH
5SL3Ros2Jw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
RCliXKg9Iz0QVLqI8b9GfxxBU1GhNUODWipyNqGvNd7T9Syer0VoYCIXvffp6DiDgM+PWpXEJgNC
ZPrITDndrkqwjZ0UurJqd8Mlj+O4jokuol/hbGtnMKDg7LMTP/mcm9YRpJxuqv5WE2ZWUtD1WAlU
7OzpzsPnbliZhM0CcXY=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Kq4rQuO4iRu44woH6WSrRyNcsAgSUJbnevjDngvc9cypuoYRq4je1NTd7KtIptAfdlUTFMhOQTcF
fyvMO0ctzr5YXTPO+6ZCPBMymjnbHRykXwGANIGORUKHiAy8zVrLHGA2Tn1n2komEaNoM+u8Q25L
d17PGNi2LYc1A9ZX79yuNo063Qy3QX5dSU2poXOWXHho+u/vL1PlOKA9tvs+dS7HzKYxYNEywyjD
k9FyesJcGgO1rBPy+iEmTMF3cKMWOg5VxnjbUI6qOTjL5ZYgIsb5KR7Wy+RP+kUhXE6TZP6qsxFC
3QU0aGkYLyynNyIHyyLl9cVQHtYz+x8w0KmAqA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
3w3EGD6E+efCt4Fs6HRylWTDMnbDGksrBmK2LrIuuDQNpphsT/R3PC062rFGmzFuJg/bLf5Iafea
N+aHJBb97H7ueY9YF/kPUqJvkNizbPUPQpBP/2fJ5zOg61lddHncYUooATB8NAF2hcSBgU35x68X
0+ZIEJC/w3FOSQwJ1Hc=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
sL/FJO3bDIPRCCsg2DyY6eC+YEqAvN4pdWi2+bTJiJBIOsoCbIwvgrvycADXfLHet65F7sNM/rTn
YIBRQ62HHXK4AhEPCYJ16a+GWujel0mLrgVipEjZe/PIBzOTjqR8RXDwI8IW2xOJhTKtdJhHoHnZ
fRLpK84QgF3/ft41vG+L+M5INzunmmeduLlvL3yJO7PaDzNzZxm4Yb6qxrxT22OrC7GODv7eJYeF
/B+o0KrZLuu0VxgdWTSijA2jO6/yo3BIW6TSbvbn1C7fQYmUfGWF6ssH9kJPORZ7fLwb67UH+6Wy
MDlUpxP5xevODOWeiaWV5Hs+S3v9MGrU5a5myA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 18352)
`protect data_block
pTK1w17Jwm1RJAcAVwn5Mw6Dw1ROtcCc+uOIfoLiBVQb6WSf+ZUWiZjkdyGG7lltZkYTyB/8o12R
eiPbU8tHnI60Aj5+a/nSAsxTrRPqhrZJ7AnQulAmxgBsVcFRNx8LbNCFVshwCLqYp3Z9QpzrV4Ee
fkcI2O2Ga0C4IgomNJvRpSedFFLRqVv1/r6yX47/z6V22ByqxpMLx7vCmiiOlOAbOE+WrDt7WMbo
K+a/1fBnumXnV/eHpDZ1W/vaWZ3CbxaJsRlkXgXL2XcC1oC/MJaTZR/Qqe76x3HOTs6BGFZV51jZ
hhze49fS5Y7FOBt5UYoqCDuOSxO8PUMG+XA1ktApelr4vr521U0cj9UzpqbuJ5w66vjbuAZYxjJ0
jP23FYsQDExVIJkjakKSl5bTri8TesXRs++pIpbx/ypqe6VJ+F6SaqUS9C/Zibf2Ubr2lf3HQpnb
WOi3VpUAHyD2uFOx5yCC37Z7Dta3mZmRre1E7jMiExepee6fgPfdSf+9yuUyTtCt26ICIu3ri3I5
8Fm54iwhLRBy1os13KsLntDJUDssUjX0TNV9i3B3bDd2cdYee0dag+q+XNpXxM4FeX9wPHKfqP0v
XPL3dLnDk5oUcnfsqg+V22wALvaDxMPsX+9jswlQ8y++oajSdqHcueUmmR2d8oRlllQfgJmMqmml
ynGM6x8+BN1fE1QCiu3fiyYp9uOS/M+kYjpJASqBMFGvGCwsb6CSCkO4WHH78n2yVK2jI0sHkpoT
9aDBgWJbU/Zk+EmfeSJN7TWaf01YfoQ9up2IfEHs6XEDvsdculO++VYPD9R4Gflo2mw/qJbcZHVQ
2SYFUGoe6rRKo5W/gAntgTDTSSshJVvcpZWrqXYLHKMosmTPXFqYVqiEBDoOPnBJl2zyGxXqaiwq
XqP9vhMfVcrZhGcVbFCFctFMiLYlivBdQyGOEitVTExH0vd4LVl5fLX+4gGGNchKhKfox7A2bxyA
6/LL2Dp82G+t5ZQNWqkErlnEbZrluRrduCPCsLvMBx2BuVqSfktZonbAyKNsSJ4IyB3GBP0q8LFS
MiDOCs+7a483HUkA5WNzENAFjGvFNcSGUFzhPsxAEhYugd7mJIaCiRz6c4kwOrGvaUHOA044uIKW
KVR6rpqDSAs/gBqtuM/c8o8Ah8yZQUZu/d01CeeqNovUZyYBJ07kbnxPEe/KPKc/Jsl9qWrtN2Q8
iyGhO/hY29xwUmWVlFxBEEcpnLYMl3Iuf+uQtkiO5kXjHJI9Ft1/zmKqpPU7yJsLb58F+Lj+jOUJ
zxLuqT3EG26v0dtYu2VYUjQCBDFpbKN/g0Z0DYaRurn9E2J4dc/N5pBD0eNSx/qYKJgBL09/lumo
Rq+U80FNnbewVyM0yfRRuBbE4LDbBXWFFVXx7dhDlQvWKeiMcb+p5ZqYO91+tgbTmZXIP2yCS1gj
hd7BARlX9Turi3g3eKHIf5UfSkMi2C7fioPx4vCQcRfd7BkE2nz9ePaOb1XXpbIE5KWDWiN92SwH
DAZyHHBvDh12cSAXn7V2mzIgYgD9Gjj3/8m+S+2MKCIQ6MFsVnG93zMikzwkjgvPRp1Hb8JEsFTF
cCbXZfN2gYb+PYgXMksgimIiu8UgRM1H+JHkBGOWt3Lv/OcUD7MUv2SCOeuYfD76Qmlm+tcqK38g
fAa/0CE+XZolCpt8buWig80RTKV/XVMhICWET2oUZ26V3AhD92jNJLhOlm8vVA/FMP/1kwQwScmU
EV4mf7gG9S4/N/J41P1OkrX0Kurk+yXIvtpYuxB15ZEsmYonDPHsrPL3qzFtxuCENDcBxVvIi9rj
saC/scVoutRS5smBYzoKtvpiSvzfSnmBNWw59W8eNZI/jgXqh4XTrq2YADhR1KeZnVHRVrnFFInF
rruKSAH4b8Xq3K+vT+s/O905UHctUw+rIMyOxt1DWUkU548KDfo+iJLJae05YYoMIf1iI/eOUqUh
cxkA1aQW4e9ADnJtlNGwXwNWZU0Z5s0hksdtE6EWs0aGVRNdXXG/lpZ4Eta4x8Ga4eOwZ0MfxOEQ
M11fj3kijS4Ks6rNb56BG0/LgcqY+Uh2u5f41kpSc3iLIkdKxxPMnsdhxcug33yjQA9mI30wcFGX
SLHJ+sgN2P6Bjlyuxult85eZlfxz4af2EATn0w1lxXpCvKkTXnoQk+cm62UPRVGfqW4AEN4sTOVf
lIHpyQ0rGvJ0auNGOEv2/Q3ngQ/9DqpKqRYKM8Swcw4uzPBM8sHQMwIlLvd0h9VZdtmCPuq01bGy
nTzpCR9JbE8xUmh2cnMKlcW8FGR672+ixzYcW5GZ4//xod5b5Amb0xktAdLUaT2hKLkB1c64ze1O
oblhATZ+JFxOcnl8guSPaL00By3Laznsk3pkK0OW/4xbJYDUWfh2uf1kJ/P0xIRhoxWhiJgYjT4u
EJXMyTQsiJYkJm3YxWiKaAjzx0wQxJYS7IyAinH+zvY8X/cWS1hSS41OqqtLGL/4lN3XGzda2hMX
TxdO/Rhr2zxzf/n4w9KsB1wXRn0Jb9ZXY6AHxtE1YSupUwdVgTlO7oON0La6j0F1igOzAu0GPgm6
mxk9G6tZ/2OwULYIRhNEdP9GIo4qqhVvR8wRuKJZCpjIG29ZVReQYnHUQ82gyIFwFGcizvBez44O
LO57U/24sK12JGL93hqBHcPLuF2XCRLMloAqsPzEPBFdfUpJ7wJqrxLTXUM3E2Zl1qJaaPJC7lBp
31bgLzjTvmdsNQrgOpkyCPs4Fl1C6834rOD3VJdoSxGJI9kcDfFGMvFcTsLiXeygU6rztH5xxrQ1
PmyaqRlNbLNqq2aV7lJ7WJVCyXMoWl5mt2qNtKNSYxd5I2o7Z2ozL+2SBgyOkYp5AF2Dsn73ZojJ
lD+pnfKV9k/5nH8zk0xESEIv/yuW/KkA3KYwuUnsOs5hGveNpP5sat6FPGKS7kyptj9U/09HJQkC
3EngKLrPSYwW3fBbH/L6+XbP28aMOCZoRRngLZPQyR5gg2MVINlmjAJoQNLtwjZsNrZKb+agAAFs
WdUGwgUCe6q02AXZkXolfe0ulzt9+WisqA1kztzPw/jy9KAE2vN4Dh8jLtln4bXNCKZt87Pd+RQm
R02sGKUFE3jEApJzo1xjpQqEzm9cvRSxEor63Ch+eitqIoxUkn5ldfaRrrq7mr656rk8XA/AIMJ+
t3itrmc2llD8Ptf7g93Hi9r7Fi0aUo+zKwxje15zbImO2U8CUAZVu2KysNCU1EeFchaKrP34djsG
0ekwdgb6hWeGd2ufZl3cw1ks8fW2fxocXn4tg93pzHc9nvNOHyLUGsAvAbK/jnxeuivmmnQq5Q4N
umI+cVlMJgbqpTOvTX8s/1IEEEn6RqKFQBs/fKiBYe+V529RA9oGXOfuByfAvCb08X6gHXQKXENT
AYiy9wr3rdscRDmutV4kvlK3qkLuUrXFh2Url0Mnkcs9ToCH0WD76+USy83SQBZfNQGs23OBBUDb
exMTJTqTQO7pD4Jy08reiKWDYAj3VhnLRqkNzGzvIFnGlBuRQCWif6bptEBQeSDhjVchmKXbr12e
BuR9CT2E22xm4/DQrLQyF6BGvGpX+EpD7PPI9fWIWkXkHXX781ZfmNrLWzY/scNzvuzIWU80f62h
LX1YJUltmgyR6+e4SzWu0MSQGVSgQFzlZfXytNgGyQI+dCbf0uSqU54xxNot57w6mFqYbbDbnNVu
UjHmvXHrlGKWgyHbjhLLBPqLgq4w54QWysXZy5G1sphKCmiAfM4N/Fki6plifAUqsK+2YjfccqgB
sAr3lbXMjLVT1OFbTa7XHnu6kgvNPeqboclPoiPHl9QtyEIsEv7wvgXoKgeeX2LNePNwuzJnBK5e
xiMg7h7sojrqIFkwgdnSWJRI6v2xDhrvrfPc2r/bosMojwPLVEywVgIeEL65T4Nmub2z5wcpD6Aj
NlaTjpe2L1HK8X402N9gbk+SnEB3aU0U2uXcJODKTManqd3xUb3s0ftxfFerL/yMQJyMDEKv5Opc
0jL8sKrk8R8X1chJb+rihfmdEiJwCPVkTfZjiW5FEMKFDmRcfW3w/ROL6dOcT+xann5UAL/btPBB
qe84gYvwkA1KhCCJmN70Ul+NEkpVgGsm70jFOaKRHYzEJHU4KJ9Ty7LsXxY6xEJxSPXQMqMnejn0
0ed9piru652BcV0D3i8oPfxdckvpN2y4w2aFFKIDVmBY0U/+746Wta78rFUDUiqv5Do/u3j2ynKD
FcMZK5H73BRySbAb2w2mei1kaPsPU9VXZ4h3aaBURacMBc88LF6UoSC84Y/zTlUuAqg0TjMMhIlK
7EUh1j9123uKRB51NakuofBSB2RWdIIKrjzTWhvEw3oXsasR4O0KR8COttRqAvQ68mEln13BB4+4
odF8yrK19fHkuiB4VGd0RH6i2MQTcJZLN/JxZ5ssKlqioMul0bHUUqMd3xoVNR1DSpoI8ilTG3Nh
C1EsD1lUqrcOdinjXQtDvrur+rorno7pE6bjuF6lwidKbAA9VBOVCbpRQJ5raFfLghDEpvrPPCBh
BD9cgwzRnv7DxCauF1hfsLSvhVJhX2AKEmHuenD2bDHrrRgfJqjA4plEApqQVw83OgeOvyDpt4rz
eoJVA9gsHfL2+qrEr0He3EJXIiC42YJJBFOQzTXZRbsnfto3/DdteXO35T3PWx0icBc2Qw9GFteW
A5lLIEvmyKU8UiMuE8LpPc79KlrhrUJKkwiQVIZFjvvRpYJtpg7Npjbzx/R7YJ7svMoVp6zXGmSR
uOBKI0bgtzMb2xwXS/5WaMpP56ItySBnRqP5jX4fv6XCQ5Z/Q/Pg8x4gDzM0nSAU2KLk1Kt77gKV
w4MUw4QeN/K5f82w422h4U+qfV1huCJNi/BJ1Kqx9zDw/UZmQ05Z4PK2g10ecHMZS+Ok7J3ixNKp
i6grfALpcPk4kALdBsLZnW1KK5IguwJpHeuLxEpzhN6MRnFmRcxgPHtrgzJVNIcaD8UEd/mhqq6F
KVG18ktblHTNPlh65nnCng1AmwocEyOxbrvjISzztioiYQlLxh5zFdgRTimIrC510t0jDyXTg1Q5
/lrtbyOWwaquhPh7u1GcZuxM183UMpvYGymI5S8v3eYrKvWC9olcFmo3w54bXI1Bmjvl7zDEBr9c
k0KFM+WuvqSgyJqJ1D+O3LQcpYd4gEdU0XiVV0NwyX2jV2teZc12q2ikW2k3A1VyzkoYuLoC6buY
rbp+86IbRD3Qv0W1LoPkuFKsmWTb8EJTPizn66TZ9fABPNGwkdx/Z5HObSzqojiEgaRObUu0w1S+
Byd17855f5dLcqD7qs+CBOhXsUhqF5LpxJQc0nbcR8jJ1Mo0CAx15s0ijIPmicXTxs9FZCeW6aZR
NGdyuoyrdYJCkyLiunKOV4g06qjR7K1m57Tl5/tEnhDrUAyVDvZ7X6hDvw4DFTII/Bod1GpOmmrm
XMFYHWBCli8jFz2W7xnyVY1GfpDrwRZXW99N1simLyCT2ORqYbCtzNQ+qeYcYCYg2LgQDR12J6El
4uZnZHdwL2Y1KyFjLhk7G6gcteFEkWnktEC3lDhUtBfLWHFNaWPYmASj/xPml2OKIiOjL5HNdCTq
cGpHmy/u/VT+FcU04rHN14CVC4yQJGyPBl2R3uJsL7ToqaSc6RZuSnLZxO3BZqkwi/KsiySri/CV
biGBcG9n8Su0lYVH+4v110Sj4v3SoB2RxOC7u7vNSFnKYbHoB7M6GJjU2MpSnodXJUP4SQkXZfir
eM6zyE2ApLtLKNhXsiGJLtnOeayFsUe4y/hJkSHlvRF6MeB662uK97o9FLpXA9zPXo/wX9E72NrP
lvLpdQvtMg4hbrOc2hOCdluQQtN5xj+s0SV9qvXDIZ+BFlVyNk7BRQgoY/aFAHtyU2svPHSOA0Ei
rcS5Ix6MFcgAnPPUNW7+DQAIlRfF6rCV71hBCg0YvniVY1nQtfizTHw0n+myTmYc/h3CZ1hc9ET2
e+myBwus554CV2YE2txtQjVuY1nMqdY3KVIgcw0rDq19R0MlrQYtXXwApQSeuvrEKBpGYvfOYA2s
XyKxPeWKcwumHxQeNiQDiuovC5OYtA4gSlFZyqsJDEVY1sDs+WRxAGjOTlsVGZ9/HHOGNzHl9Wpx
MMlbveZi0n6f01CK9m285/3D6R4Dd6j9Qwcp07JE7+J7X6b/npS+wpIyMHCFvp+S1exFbIMH+TjR
phSYPEbqOl/T88BDZxi9g9Twt+t0cag1qa7t03Bgd6Z1gCZ4rf7QMHnIqXXa7ofln9JtWe7WrJfM
XXrTmU7ktAImTUtmuJagyrzsniOFkhzBRhwH5iCkBu5+b5bmryqUdxQc8/BxxgoLIqO2339lXgnY
6DIVjMq+KNbhjV/SxQeTlZ3OuauFMunlfPFbjygz8ed1/fs88yFWxxQc2zZlIoEY/AMjiFl3+5zL
9A8tgqZO1l1t5TRtCJvhrhvJW4y04G/tLGw06ZDO2My8+tNnPjFpYQX1GIoP9BY0OAxZY/c3Ho3j
2gRDsMOqkmr6XQXBe+88aCUBoEnfmiNl3fjPeesX3A681dYiDyn9PjImSNw8ZsMFgL64BwQpB2Jj
6PBNKXxpxld4l+bpiMPadLF26+VnWMJXEPAWRMayfyQs5jlJyd/s00+y7K9CihXaXCbfzYGszLBl
+L8OKTIBpCJ998N7S47pIfCjpWk+XM7kHhfOnwerUphJ2oDoEviZRPj9XwlMhGcX2XMIV/Wf4fl+
ruxJXqstk5x0yQeLrIoJi0Z47FrDIgFY+/Uf/KDoMGTaCg07eOccUxmZwsWuODEyCZWfd+yXZ/rM
RS7MyQBYBQNuQqPVlT8P+XmX7JhrKdA0yRPwCwYWHWbjyuWZYS3RAqu2YDEIz92C7edb2gh3dtXk
8YupCxctkEZ1WXhyhALJvnN05N6t8dkoe6bLq2hvTXwo/nBr2CptNkzpiH/GKCfaTd46CYo4tUNU
m8QDjw3/vh5feG0aawaurFIX2SWKTvbyaTh2pSbj3TFMQI49pYXES56/zuTnn+RL4VewPHXDPCjW
nSt5RLjv8df/GczBTc1Ltw9o7m/2Vs8DcpLVZsonx+YGMwDHkaXfGyvDeVAit7GV33jAZ/1UuBva
liGKUEYFTjd00U5pqvh+F2j3H1NQMB0ctVYe3LzHAvn9YKhO7X48bUJDEW3k0MRUByYQsFoUj0TP
ad9OejbVnR3Myavr55+5ZoBxPu2e4RtYnYrq5Po/E0Oa6JsCAJwYIKyHLeq6KhiNa6iQyq4P9PHH
kC93/V5k17H4skTBu9UyCEzp2t8w0euVFiIGaYBbzlsWp3NvW/O7U6nU4enMlfWs8HQZ0ShouCRp
oez6mNeY74h1MStu4kv7F26Ra/hwqWi6HApMy1uc7XnvafNyzALpS6A1DNYwde8q4Ba+Qthhpckl
2xJ4rijPcdinQ0UXSvhDFeqss/LbaKL7tPAgIcf5WaYyt7ocvrEMx7sIRKkhZ2sjVjKNTA4ZSHVN
5ZawU1tkNtISVzldi9sULgbay06Ry5JuK1RQloM/RecCccoPRIvak2pXpoKW+wnxzzx6eI8zoMB2
5YlnUjAVTuIkQHV5egUrU42iMiX5lR5GwO2Gxmv56wzYXNYqzN4Qioc1JDuCj1dtlfUXJdEpREOw
tBqJWNnI1d8zjHmHVlb5MIofOn1tsSkUvm6BnD+T1prYFNFrtMRg+s7WihJluONH+jUjjaIRVNei
2d5XlZ5i+kUB1Y9YxRwHxLkpotMM8QMqo4F0NH7FKxfxXYR1HFerqxX8pxZd8kKv1jokulCHWTuQ
YvN2xIfMTxSL3ifrUIjyQ3jmKrq1T7zfbtn+bQDCiLMkZDsH/b/e/x8QyGWxORrP8RrLPTf7YkXl
Mfco6xlxGCgfRYf8XYr7MqOMSNZrQ4eyjqeom5YIARowbFkrorFVpZCvLbhlcN8M521RaXPvSDEB
tgTZ1cqKN+qkxvVxpNj00t7M390+uPkZ23CSq0xuxKmLKcEOnj5PUBMjh8woOI//pKL8yR1Tvv4b
FdIrQAmfvRworOrJ9eeSKLz9/a9JTBGIlIu9gUnzYehnFVl4anpoJ9U4DVw9fx5CmVKeyze5C1pe
YpQMukLf7NaCIawx3A47CsT1i1z7yOO44ZvPzjNNso//kRqc3ndNaopXM6YfTV/oSVVRcvmpZBIt
sByiaGNsHt/ClG5WxSyV9WbdyG9CQ3G3BZ7A0T+xiJgTh6noG0dk5QFVIh4Ot6zunFyaQOjT46rg
yEiaKq+ZI45YqNd3c6WX2TE6wrTlcvK5IR8fc9fXmJG6zKVwKsvew4phMTRPb16cT+s0zii7IVHt
6lH6DNbLMrbw+iW8Mkp2Nx7b2eCQAp43ADwPAzsj1QFpwZpGB7SMK/FCbS3ImYqWRyk2pCQFvRnB
+mXayA3gGBW87HKmbK33f8Oi/Lvh2D8/MwtXx6NzxLHgMIkxB22SsIlubWSRLIpoHFctQ/+QImkV
tb9CGCBA969Iig3YKSgHzMJPitMrs4sHGIgJC4aXzqwG8CoFatpVJbpaCWzevLrlowmfKToVh09G
BD0KTN6MKygULW/n2NT9wug/PNsuedgzP8I/LVx8dp7w0Cgq3OaR36xPwumLZ6q3emNh3V4JHWsC
QjpHiQe3vc3Sr9lgSOglCA+1Npe9qz+pBzrmubsFg4tFPk0uKuM+S5AjHkD3D6nIIe+0b4PvX97y
idEAS1pHBlw8ep6Plj1qPtuz0p2oEzLxyjFER6sOQ6jdolJBe8I1ZaYWDURtPehs0Hm7RKfieBQR
0Ka1BOyeT0snq4o5QUgVDWyFj3WI/pz9gy1KZHqZ5Xu7jn3HrXGvOVyuyrM3CDGMmVB9E9oM8r0u
zV/0LhwG2YYWfbBlKkyUNx9TX+fBUMtaj7YoAg0qxKwLNk/SKWdKIFep2bjMzYlPqSvpnmvzDyb+
lJsw9ls2dpSIkK2YIfsBa4JPMB0iNTMyFIaWVngEgiZCdJNsfEfF8rz7QWn6zAbciqxR611T7Dxl
zs69hysyF5+Ur2BnK3dyEpzcR+Y3H+B8zlCISMv8/Q2LlGJtwu9lO66527mBgNpjQPaqg9Pij9QE
ZQ9aoDFtczPw7NqHWk6JTbLJjsimo15P9o8WuF1g26CNANquIL3rtJjfOJdeWt8fUv7oAp9eGug9
d62izL6BBqttbAEhqw+3A7z7TjBzGoFekcL2R1uNnkYMwgB/UrUKktmKL9oLu+JvoKFcv6LN7eyN
enAsqvmIASWXtIdH/X/P0B3LRmit5Q+CBiiwpw+1LUq98L7N6FxFCsLcHIGBXGwdCksEMhPwdQzR
Zy7Zr2a57FlXYQRriEu4DD6MwZoUvaaFtxbenmQ7qL6G/NZkKZg7iKt4maPKkypOxlR6IAeK5ohM
lf6KnCDi50b2mwpPEk5a+RGFX0wU22lcR5SQ2rq6bAruJItwDizqBCZ5tBbQnYyoYICGcjJKyePJ
gEzIIWwUhy9jw8tXfteR92/F5vMR/Ru3BLW3+ovOIRwqakaCpKSH7U1VsHUUcyGbtLyydPNtEvIw
Noyu1pREaZW/A4n88fvKd5gfmt/pa82hATa687St//sdKI8pUtoO8PtLKbJDJubRRrOQLXfxvBPh
o8Wtz8LAI80v71D5aUN2zHRu+ZTj/rhoj4icszcv/QHnio67oeYLq1WMtSR0bBZf2uUww1e/f/lJ
DyxAG0XL2or8oe2zUa6IhcmCQEz2CaJVlmKwC/0jae+NccouwpaHSYupLWrefcBSb1nTSjJSPume
xRuRp0/oXMHVXFOtKBjPixGL/ts4FuaESJdO6jisVM8Yp1ncGANgfmQRIWn7EtTbb/wIUczpAO4P
mm+kfvTcvqP7FcxHmNZ5SiOo47NvPaiL4CsFylfwvBxXIzXZn9Yi8Z1B9aXFIhJIrhA29xOs2XRw
aQil9jY1EnCagRTCmfoiXJsAZU25PwNNdUgPlaqHR6/1pRcwGlGgCUA2Ojnnwl/InvGIosfr/L0z
zENKOIIK6QszAxFi5muQ0yaOAprQpKQ77rY+GeiaC8wddG9n+ja0Ttdoc+3h4DbUnRRl3XBTga5K
T4g/zjjjq8CptgSIcH4Z2ZYMqfN0CAS6JErDjMLYdg2LMafhLOXz5zoAk2SfgsNL2agIOgBfI20O
//Th3SKck3p8C/2aLS8dCmOmOQDtNtRMTIem80ylyAsPOV6qwWeX/BxNeyc/eDJ5xwq6gOjA5ymn
hsXugZ8lRpm/LHVGLXGQ+bDTzxRfniIfLj36Fu0SFOLxMDSBA7PA9cweYKX0k6JbqhEET6mOhLlz
MjZ9YXo2L2QezkCHuuf34rzMOIBPUiNEe+jhwUpmVu9srlv+KFWWQRcnUhTfksB9/3mWCVpPdu4b
h7g9TE+NDxTJEg6o0k2bSI6uqu4P+9ToFD1oZSEcUS8MonCvUsyqrO+sq66uLb4POtvOVdjQ4UG0
UbrKDkuTcn2C3uaxK30KOTnbdBgvzAHxiCIJZZc9kIVW/ud/ZWWOvuxaIgQznw9JKzOBIfL2C0cr
CH789RUVpbBhzdu2h/2ZCkDUfS//dnwWRfctijjGynw5vZku6IC0rqni0CIiqyqGgfsu97Vs0F/8
FNjQyWQr8P37yDKWOPdAYG6h2xMeBZFAdQIxSe97lPTtaD8L1u6cLKEzSdyFFYSG7YNGVCCre6J6
e3VX7VjhHLzMWMubKZeDFuaP6DOsp2c9fw83yNn1NBmCcDj6TULecvMNlj+6A4cZZRxwAfbNYvze
VHC2BGH7n2/3p51Pf0FF1YBh6Mruko+piw5sQonXeYNNVf+1dNe5V0n8nsdfrNMAsdaHpxxA6EC2
t3aulLJOpcip5PJmLoXovsCkEt6nraRoA2/tuUREpvl+sF8jRX0OzdXmYvl1ofVCw929ybdc5Pga
Xgu3n0A/6lj5O2oWURFy2JX5UYpvSYBo8iRiozV2cKe7N2BtTma6mWXbgkqj7aEcTnFCtS6fA9hw
RnpQFOyPE3bLg75D7TiFd4OquqxtkJ2ecyD6Mw3P3KlMd7pLHa83J5L87bySCnhP6x7o4W5L3YIf
arS+luy4xsU8+DlETCX5fJoxO/Bqf+irQ8IISOeUkstAqU4+UnYnbZc9rU7DCJhOYiEbT5HSj+Ek
vaHBf2TACynla55thtAiosG9slKOzMl0Cn1LfzxNSWXpBQCNzwI3b34CGqeSImtq/721++HLD4nL
ZS81TlRa1KBsNtw/JiJoa26eLTlRImuNX+ces03auNiBmk9CcTPc3uvbmG6QIqKNxDe5sAJHthMQ
YM22l9nVVm6UHDlacW1F5m8aUFKdLmW4xYHON/C8ThGsipcO9ElUR/IcIQJypeqjq4MiOcUFVf7u
ybiGE9B8LNEINCCMBR46Ku8ldN7sdVIRcvLTov+l4N7JF4dVgoETYpL59q0nI1XpO0yKorXIRqma
yHasZ8Rg6NKVLO1QmPtgpb0yH1SbweixG7WJKolgvgQthvgxoR0e8NeFgfvBFX70yoAoKw16STu3
GIwgocTJTWM6sSpZ0QILgmx2J9U2EmJV1yBsYcQKua1zd7CbK5FZXq9JdxidtpW+U7dr7gdcuO2z
FI/0Xna/cMPcyoQ13ZKzyc1hrHTd56G/wdTWTdcc/C6B1IAYx7TLP4RNxuGWvM1DOSAZBza/DqnX
heL6NYDwm9nOhnU/3T/o8zIDhVrl68J1OK2ZLMQJ+hvwRM2zhkllggIgoZMaJJGsGvKNfEbtlvlL
ht6uehuod1bK4uD5NKhNa5toR8qZE5SXTPRCzTCaAZsmVe7JOlByKCU23zW5gQRB09Rljy8REd+m
GL7tnd6+nDXOD39HXQVhvfjDQ5XCc6z/7PW+ye6S+USzFalAHlxFDvj5Z9caU3QTRLhpI/sXDfqg
eLJA6XDmdjm8V7bYL5zXyk7P+QVPoOvn+cm7baHzAQ/xG+M0O4yyx93VwWrLlorbPD70ghHLCP67
e7ZmrCIb9fhaapdQjTDm7ThzaENn0p1bK8jnNjUBeN3zEFsRn6HAc2ZaIcJsWgg1W3145FmxEJYE
ZndV+mBRkG3KO6gg4rPgeIuarOBgeXo46iYW8AZ7IVbbrjQb/6oG3YDefoQIGV2tJXlAx/bvnAky
kYAGpOFF7kCeV8Dk6jfM8Up2tkqtwvkDrYnvp2dFQv3pr+tr8tLUFurhuqua0yk7tLS+oxBrDmhb
7qLB8UQiS9Q5CxJGbCMyozri0e7UpSmSJrxuk3UG+0L39n1uLaPvdXNaEp4iAzqGpLf1F+kCzmsO
8zV/7ofNpbHNy/cdsloXvXCblG2jrqLfl7VDzO+ZOtpCaluj9sBdhA46anhTRdO/G9ztcP3puB6Q
zvulm0B79xl89Cco+AF4e5AfcuJLlHQYVg7EJhxeSAsnbrVhDxXywezPvBxR8CaB2gNYwi3cr+sO
/XPJzLQgVc0DHZsTJryvbzrmhvqvqkEoaWc/lPWk3kMuDv65WQVwK91B7f7Mi7zrkEaVRSiO3GcE
Az6mpdAK6WGudkHjvk3FAVmdaLF7W40WsD46cawMULAVaZcLMHbl4HOnBFbTXOHnoMLiD/JtBOPa
RwX9xhQvTR4b+IuXulXSXjAo4xXTffdycCgRY7xxYWHyGBGEWqDh7ORwmehhY3mmRXNXRchbzXQ9
4fX326YM9OUG0Ltx6iKIRizWsV63iRGC6z50fqlRTkFZ7DIgycSJc9egVxrXDIGv1zL0F05UmRgS
dVs9jLSgAEK+FND+BZqyjZWY2GOv3fip55TXwskmAgj8AXY84CAjdb9KaFPSdDdQaCp6mM6LIcUk
wIZ4AJtF12HFubrWpHrkTVouHLEPwk1EUxslOJVrZvgOT5d2wa2NHm3aA9QfIrWlnGrUDPLuzN3J
90FGHIuyxxYbnEwpaoowBN0t+h1LqB4z3gTtOX1xEclwCUv/+JtlpjpZzOk4RR33f3LNcrDoSFq1
8JG9FyrbyQzDtQisj1BxaYRMMb4cg0S984NrFbvkDmfMe1AJg5MJA4j41seWFOMORDIHqvGcsNGP
op8WRFhCfK4XR4eXEB55Fz0ARrJOtd06HsgMX/O0JdWw8VtyIUxiBejlIJRlgBjDwAAgmVIL9nQS
wUFc80QBL4gNXDyDYSr6G7hZHYIj+1m/6xpyXZUrFzwk85p1rGBr4A5kyb/4ptyQjLW24bXSsTVK
OSVqtX2VwjtXtQXItNOBXtFcNsklpFH70ifW4YKzwLSBtLtBTF/4EiiQeGFlgl58qBU/8IOxVIij
ZmKc5p+YLXdkxyDQDj11PGjdJC73NMzlHK0hzrqEg2sfZ3k9Gt+1xLHUQdwypDwPq93Qpx2NyKMn
sC0KZJ5O2wse+3oRte3HhMk1BiBm0r47aJWxKsYM0uvvtCsc/dx4qtFO09zYND3KrnTr1RqzvC3H
Wviw4fD5yjDoubhhdnm+626ld1J6hGwe1p6+hKTKeeOQck6dTSA96XXv36c+TTziMnrrD/joc/Uy
ZVYY5soH8iGsNksUtaevprd2k8zeVSrhmEEXBuLpoTJHt5AkC5T5mko8hMKfcA6T6D8qQpcT6oXc
8FfCXRtFkAOTdiDmYdUPQyMX1RevZbDqVCl28XVHC8k/Ox8tjVQkpTvmIeBfI4I4jZESQrxZZjzu
BNRzAyf+yj1/DEbNX1zVOygEvfjVdYEkmk79mJP8PoSDk2/RhftXYhKerUenDvBWnq8Njvn/DJ82
z3WEahgfWlnXzvlbTUFTgnffySpdPClYE6tgkA/q1qRJ/WjqI5ziaS27nCJ1pwFJ6EadZ1YmzMBG
v9uVOCF0YhaXStdHUJi7xLU0w6+Tb9e7CerGD3nytQhnOxCO0g7T2ufM0U6gBMpT6D8pP2WW9JXd
mr5PTFoyz+MkZPhs3ScVe5rc2+nfv80M+uoAlPIlyoFUOZEIl3QGZFdPRMQN4xr8IoZiaDwsWFLz
OwvlKk0ARfTVTZFvDbsa1M0CYUoRexzFjmfe0ltIaKRw84Js/no9MoKRa9mqc5RxeS3Kz3CBzfpb
vNnqqn6E6uo0/J5hNRZ6uqUwSUysHSI11Zm1FhxfZi6bmgHv6BPrXwe8qJZ2Elt/+kW86tVZ1a2q
oo0oxj6O5lF6zDhH8cX93XDBsUx+V16mxi2HSQXJ0fRo9OkmkF3uCIlkwU9xPt9LFIwYluIqT6wH
cXjs1B3DtKrnIY9ROB47siptBihdvvM9phvV74lm62hA4THp6Of2pGUT3/zRdGRs56tVZphFGb8d
5fdu7ANcXToyYq+w7alHuYqGWhqUzfKQFfbtRNOTiqtzIf7/1Xr/9DYtYCuBGiVdGXeDX7y12Awf
vQQwSS+wRoj0hScVoWjaeBgxVdEK8J6FWF7ws41Uqgp3TZeyZZ72TKyE342QhAfJmnKUKxorNgGX
gLLKmHHaoWSexKJtej/d75zAJL7VwV1lxUapGHBUQFoyvOX6/q5tynbd7hA8lvOHC7foLgBPYin6
ArFbVizUrd8CcFK9y2fFBQTCqhJYhtHZdR7FinTII1mRRgSQGWo0eLb03N2xL2rG67FUZpO2GdaG
snscJShzpsqMoZOhV49fdc6OOhDN4v2KVsApCUHXklac0dFpaJPIjZzHEb1aO1jQIDefhbHPQz5n
2Wh3/vHyxWSDwTBJYevCXoX1pJYfkDxaTU4FDEpMqU0BS+WUl6BfmAWyWVw90p8K64aVfDiWbTWM
s2kzRx4vfL37lnKudZokEOAMimJQF5jFAi28b1qgtdaqPQzubPc+rxdzkwbGR9Gl2OqamLFtG3VE
UOK5ngFG1dkaISwEsdPO8KAfJLx/vz6U2tFVHv1TXq46OC/LOsR4mCGWYemzLeZnaYamEudeEqPo
83//n5v6OyUamKDUXF3lfKv1k/M3I30Se8Ef/bF12c3BuIfd7J/FOztvDx8GfFafjfiMlYwdJ0x1
UHYytZ3jwzUT9mZRTI57YGV+3d+vfgMrHHhe7aNaZtHh6jMgQgycOOxkSFLBtmDDl8TCuXWd0lQz
CpO+WqcTDk2smDXO5Vs5Cmh+dupWCYcIueMM0LyR9arrYJIJ1/TTpOWaPsIsNEi49evb0xtKdzYd
ZCMgcuf9lWjgagvH4tSNzeNHdW1e2NgvyXve+M7+Kj6XNrP/myQ5b539XEIWiexf5MrYLR3/P1i2
DCaIM0jT0DWiAVBMzhidi1NEawCm8fNDgbuiPA5X35XaRJDg8BEauFb70cAZoSDJLgtMWJ77DyDJ
fQIyPGFZQyOged5yh+xGdFaiu2CeP7Lp2aVYIBI0jElHcgRPOsE4B8nUIBpFjI65dbo60nz50sri
jbq4WfqXCew+jWKfqQSqAX4iuX89+m7/uj6CSmN8Ac9DVud3Ty7u0mu7mX+hSUmPMRrUJWLFfohn
t5qB8sF2ky3l6D+vljTBh3iy04oyrWZo72PQCEhuTBPdixRUAPVzwLSrrjybUd0XrObqqNGsJb1S
hUj7Jn2C7s1TRJnoyVKcpvr0rxlTeA2xy+NJ2ZVYcEPhz3wRLHkSmoOTtiakTnJS9Ad8DWZt+/G/
X5F222/czkkg6rIByZ6szSYTEvuDVo006roWhFFlExwzvSW4gZ21mzDwu/goApJF+SChzIo1Uin2
JVie+N1VvxGoVR/Lsydb3KZWu0CLYCGFuU6qWE+MXa0rMO/EtVCf38PLGdgpo/JuUMnTJaFgb0A3
x9jEtocDpiDj8Ih3COFxbL/uybykAh1jn0QpK1sIP3tZBXAItG4rQLZpxNGJEAJnHpU3oTJwDI3B
zF7Iz0gpyJ1yCTrwdG5WvCe/ikn83lPFmQKaSkthgbYrtg0/fqFgEvkp+zkdHIwwpXdtb1YamQY1
4rRA5b2o+pDiNc0HNPDY6NUyPo2GbyKy1crlABeMo7KIhF2GAhZNZzcrzWozyQakwPT0p5v5uPgs
VwmXcGbGBi7lWZCVlenfv3+flgCn0lfirFB5ymAV6qrLDO6HmbWU3nqdMj8TouQQMB53v6swcI5q
ocYxGKuF4VS07Rw4Is97gkMW4UaPSZVjFv9amm9Iciie0gB1+QagdoBbEILyP3ns9gWDbVIf5XNl
amJ1dfnOngyEhzxB5R0LWiLgoii82P7m3GqfdOJqKvTQY8d8IdUfR+dwRPyJmlHROchGp3BSh5OL
eFRnlT2hQJ4Ba770Afku0vucEeHaQoyY++QBOEiVqJG7KRhlEuc9/NhbFkCdXmS3n+1bMnv8RwqG
ORpUlaP6QRu+cfMUKGKgKfj6gGzX1cUr19Lh/xoIMuIU/CVVUP9uLK9qGT55EaZNTzh51yoC53CD
HgndDwca4ARCtZzPGe9wNjSqb9m92ZUijzggAehU0mSNXgX17Uxr1Trdt0rsht9+7HWKX480opXk
KZ+E1Vh96IGyySwlbZ7KqJd1Y8uhnkmhgTTp3G7h+KqXh7lpU6jJO1nn9wOyPQePDxcXvasILmk9
qYYgiqzUs/iEcELmXbSh9Sv6kUyb4YbkulC5FIcDtogjh3hZyu2yMxRnAym0D3kJUbRRx+2lHaIt
F6txGV1zqXI4o3a6ZX5VLsZetYZvVWxtdgdGdk8BH+c3lP9fhns+82dMyIBZ6AspJzzsLJGyV2RR
9KbghSCEOJsQ8iOIQAfCPhguzPe4w1gpLppSlE8qdPos3Omo7WTKHlgV8hcXfMPsQqUxRLVXx2ud
EY3FSjGreTMnF1lHATRlq0lUMsiQxXtzRc3HMiB8TZ1juG3rRQfa052k8YtZSCnL7sBYar2xfphN
/r7DHt+/cupHJxhKNjjlaz4jii+jLJ3IJtNpZz+EWHfSNi0lgtfNYv0fsyACVenK9iI9Pwg1lwIT
CQN5glW/WBrtrS0fdFOB8u7ROpxqz/zNzGulJolqNR9zC/LyNRNyIliCb5E4jd2eHKrRdxbeIVw/
ttoDEtuVjv7012muqno9lE3sD7J2zokeG3Smpho8wxW7x0uTEYDAKI8V32u/+p1tFLri4o/NbLxu
JsfkZFpeHr635qNQiFh+4hdVHFbCUTcnBSO1LVh7nI77Spwcl0evOUUYpim+2WHc3Iio0m7tv9Rw
SqU/GRWSN6KxN4kpqtMXdhVR3516kz2OTvzLGnddYWtuz0YYm76AafpLZZOsMexFuuUe86krO9ZX
OWhH7HLbqTfwIVFnvj2baAedWGbbICsXiCGpFHx/wLRRe4MvLoniDRx3ct2GQaQMVp3EH3hfHIy8
fGoFWMNROHshq19YaeZ+Us5gYQWMUmzjEsZjeVjveTjcMvvv1GHcm73FjNLJPoBu+n/nKFjIt6Rc
Q5EOI55/onGI2XK+/l3NOh+XW/ly1aPmIpMmY8IowHifaqcPPrM2v2OCQ3fEtCPWZJikxGk+Dp5V
pWUEBmm7yLvPItk/ua2pEXOtFRUaSEByRH3Vh/o20pdjSjTcAhrRdt1wS+BldZnIfmMqFr5xddJw
ddB3IlFGw0+14cd8F5OuwRx6ubS6zsKP3Lv2mvXL4jnm7LXyHeD/PtZJvrfXoX4HoH70P80adVXM
9jCItPEbVTUoBlpvzufDY8Vo5TC4yLIqptSfdHEyP54TGiKlIEFVb0TtTbEAsN5LIuhNe7dF2KGt
ckS8MJDdkKQ8qOoW172iiwoGhr6e2qyHmt+QD6QedgD5xl4jbArZsGgB1VfUMWxYfFzAYUg0514m
TnjixokdYA8Q6yucm543OcVRgtezllatrOLieCnV+X6NVmj/0pXicMYKXJdhcsqZOuzLLDaW8f19
xYA/LSFwN/ly07sqMfHrKUyXyTyUhkRUIq/i7QxVuuTkrQkewRNfO8Lg/2hDx8HstOM9WVUEgumV
hv6vfWtoXHOhGUlM8jj0M6x37+DeCVa1g9CShzs0KlFjE7Z9sPyuNeRtZNXVq4fO3hi4clngkRzz
JGkwdEW1zPzYwS+nta+9oNh65QVXZ6zJTyaSF4eUDVJauIrL6z1vOcmjKFfredwOViz9HwpVfyDU
hYCtvTgeAn+EnUw0KlsJzrXkuwhw60ksmretDWPsIgr3ZcmWAUNAkfDBhlHMI+abBAHPpdGUblH4
4kRSo5B+wwRx+Q0seECB0qtc1xG/kixHPsbHBcH6SLbQ/qsbYRt8AGZeIYGSZlNoiKHMqiad1cNA
qtMUBbMqIaj2uAGqnLwmNl+ENEF8zrtwDCR9Lu1XvoIMfzcfaxIikp1YWR68p9CGOpD1T7DFC7jg
wmYUts0BZsIlC1sLckyriTPqEHA5yO0BE9Z6ypUjHlPNxamx3pZPjrHndQ5IQ38WLGfoA7F+J65X
IYF1e55j4AlmDVgASbtm2y0TbJ1+Skq/LO6ezZT9NDlgHM+JbzTlquqYs6IAgTihNxoaeTKwDwPS
uDnD2vY0cuOt/8F4ytPc8yhV86yCWPJTql2yQFTHZK4UwwAwBqkuNmzY2svgUqECxUiWhOxOUlXw
orISch0RoSX2CkafMKItDrmhZ+RaHVLxfrg8YPt9gTCZ5lEZuWiAunv04OV6SmQbpZ/neBqZZfHJ
UrwWpbimCwTZ9Hwx+mtcXWxjkqZx/tEFeufDonE2vWeVvoac53FpwHifx0sozTnAn4bZAxmSVcmp
XDJyY4rFp78wicvuWnWIHwRbFcH5pEqrwTKgIFxqTGD8EELZNw1xivtkQz3TuRqy1R9Nua2GA15/
kuh/rg7f6i3MRUpMjUv+qwz1cGyXG4MbofKWQlk8eGwG9P+MEsLmULjQzD9THmj/nPUj+FmThfir
eIbFZDr8DlC8qyfrcYq6dUOTRnmyRK+/UnPeVVeSvnSwpUYUgpp60opGCiQWTycalrZpVIK+rFlq
zM27lEORgJmyArwc5pW2DGMh3nflNOvpI+CMboLxtTICWmQFLDw3JbPkNmR0kuJXzBt4841rq7fO
4kn9LRa4d2yR7rStYKKzqEPB/bkA2oFC9SE5ul5HLezLDPyea5lfz01U/MQpGjwoDaZlG8Yp1bSx
qbz/kETo/njbdxzpAm924bLzucdguUsHmOAEB6sW9yaFcxraYdO0j3/g2MnyEn8W7I0lNLHZCv/H
DBXZCRHKvObBsgjXBbeMeGAOjm8GEV0VRV7tsZ9oP0kpZI+6z5vIvX1wrjrmoNx9T6NyP1sFVJvt
NHhctaZ9TTrrOC8s7uiMO/YFo/pNvHO+6OTl+eB9R1uwarpwtQAIm3RhIA5VaK3dX33+vRW2CaZr
dR80q5q8SnrhjXkvV4zOXw0vvL/ch4si6ImBH7L3jiNBufmcTcBCNZpzdgwCzXhePXCa5mL7dIhv
mkj8VvmgaQ3VbPF6k3MfI+a2aub9mQolhzF1fRXpL4O16cZvSjKlOPbp9L+UkouzT8WCqoRISLaZ
AhfSHvVw3nRb0FWsYxXOmayA0HWF3QWIrmxPGMul5gB74pvKQ310m98LCTeN0OOpoPk/wBtVD6OV
l9TNrzqh7cRHbQQBjPjpdE95janlEV/jEdQvvVH0HAascG4bFfqKPT7ofyCih8czpwmvGazzfCYO
gBAtcS0kDz9Jh2X8hfScxApgVCWFVybLVf6sPmfjZBFpWXOD0jYNi+MmpaK2M1xUNaLacgH48hkG
ObtyiuhGd7CTElG1eVAXRB1iQfjtwjrxnaKCB6x5nsyrhVF3haD+YmXpcKd8DjfHXkMOY0OJAkdf
FkxQSKZByrkXVotFl4OBkMxTC4VcyYXkXBURdtBBw/0CCX6AHZt8MruEAylTnz1Ag+59vtN/1f8l
hX8ZxTFAfus230hyO42e2z7ObmiXws4dOSLZ5Gpvd++t9W/Ak1cBJJs7HEAKJK375ACup+uUyBlP
CRB7BIcAFjmD9mepezshN17SNDZ3RtwNyyRZIg22+2SSViCkyTa3GSJ4knZ00IEs2kpOFdgSwetg
OI5P5F1z31gLFudiNtT38YReF9KMSQeGTqblhJ9e8sEpoXSf9jAulcVfK8XNR85z7ocOAuQBN7iV
XbXh66G1biH8M1wuPEd8DoGFVSflCQpXf63r8B2sz00m2/0ryOMV9iT5RkwAf7lJXFi2vCd2dLCB
cE0GeBfaOxyPq1Zci+9+26Q0LW2OgbRxr50He+ujV9iYZfVBG4kvsdLqQpFQzPmi74MOqHGFLr4N
hmFUmQXBA2ooJPmBhqNP6ylaBm69FeOeLPvDLdEST62zhX3QQQvfRE5tUWodJViiKfGzL70xjhle
mGpvUOtfzHJKUTFSfAQ46e9I8wPPtgZmqtcNrzhCe6TCCvj4IYf23mHeI1/Y/2rbOeQ/SxdFtpbr
7GCEFneHveo24C4LaqrmKP5ibZig4eweqoR6v398v81U9D0+DWMrOKHhQQAoFRzPcSSbKaqLChTz
ajxgVsBhXZfFqrkpf0BiUuw7itpKZEJqJhXM6iFACHfPCmJFFmlToogrJdVTdbIDX1B/FAN07/IS
obPfpkMOl1nks5rWvC3cFuaBr/b1v+g1SJusvij49AslUhwBdltNwemvK9G806Va6A4e1fZ0dUGS
2KN4eU2Cl2H6QjKMOKzLSfruoRfulOypi5aFI4EAO1jO2YD4SCnfGI9aiwCS209G54dHEJSkTTXV
dTZLNdh1LnRgwVK+79a2p6poTVOCHBDhMBGNu7qFOo9zPugr7phzLT9wtpO4NWC/uUQHPflKumI7
17RjKliVWZbtyRfeoOGRpRbTXtDcmTecM7NPcIq4sAwj/0Ti9QBSVbEif+6n/8ukcbH/VAQYcnV1
XxlsO7FxqPDgFl190IyQ68Tt51IFNC/KSQ7mZOLbX9WG6xEynTDKz0DUWZfXOnMGYUbwDY85l69g
Sul34Jrdx/KFiBHu8aULT3E3YWnNVmlfiQrR2DZ0vH1yhppA9QO950pVhDPqlq1qcDSDfxD54R78
w8snO7B7J+VkRd87PSGq5bV9fum/01ZaOKGigmT5Kz7sotnaAkngnDTH71kf9vL9dKyOeKBbNXea
qHXHtLr7ANTLd2kNCUeRRhs+wpN1fhUBFD1TrE4CQy7tTgBPo700ULoWnoKeOgVIdcAT0J01lL98
d7nYpcBmNzFsiGa3H26mdCIysTKTlTmyLhdBymS8wQ3ZRFJwnyR6XIbS76RU6MEboN7Vk9x205o/
Iu7wT4Aw7ypGyE3mX4VdBTytLEiH+0daNaD5xubTcFl/ZntWX5snojFkiZQalfMoh6VrHT+EzP9N
VQ36Dwtqt2EMQPlkYAMSfvSJJKwyhGpLVdpXWZAID9cm2uDRI+1VEy8NDkJP9Bj5DX0QQ1VUJtEG
jeZs3KUaH3qNV2hE9ykVkh9/B6Y0UUeXea3RHjdNKsmLS4HIFwJteEwJ9dNkx23m1y2sMpBrWL2f
Ky+c0S7FG9J4GmO2semxH6VuI8xyzde9nLgDxfQMLDcOEIsbnIKsFe2r6hVClodLoglx91t/U/cE
9ZCykvi320nsjVyMCrabGyV0jZYNnHWuAaSFZ5wZkJfaIx+4iOpnDq6MX8yUFdniFnF4EI9cWhB0
0gFUL9ABCwsJMS5Do4qSx6wcJWWfyoSu08LUU0BriXr+pHZGfHUAvn74agao89edwEH8zPldrqxC
3sOFw4uiCaw6f4ae+BqDTWCbS6E9msd/cj1aesrAY1u/TiBPw+kuqXtCg1hzVLm+StH3CGHriIf+
58nvEM7myqBwZlGwIWlNjLT2XYxwMP2W1waQDBYhh+r4snRV2K/h/JlUfAAOcFfQi9/iG+a46w7v
fg/ejTGxnVUrcw+ESvLY3LdWqqedRchMJ5Lsj9XNepbv+0ccI9RtqOMAuLEP0wYGwBPZYrw6rAAG
PedEbFUnuqNVYfHPjlIDDPxkNAisYKebVBKtePheHsWW5jEfknQfU1QBwSh0t9RennujGBarCwEE
5oCG2uBi+2GJVy7CulrAdy7fSmrgyA/GO0owRyQVCZe5qdhtEfEXCbJqLY8Ha7SYuOXxL8DeJOx5
gB97YdrR+02pGsrqR4Q9g0d5C1DTUD8btebS49e2aE9ptmESw9/Qj+hGKcIbtsnGeFw0B+peOjS3
uF+Arwrhy+kbpJAykTDolHWbpmX4RvBwgJFiP/A6ZbgbONpBsgxaQtws0+v/CdBjUgtZjzgGhgDS
zjLj1om0xZO6oJRCu2vapSLuyaes90+ykXdcixv52Xrx+3R8q6sPeoXG4gPorDSkrwNyKhufrJm1
BLZ66K4xnYIuYp9V07RnRfgqzQAovqgAFajEm/OAo/BkzgacQ+dQ/Jfu6Uofim6dp75vzfRmCPAa
30RqhofiuKkmF0hBePVRJxVHZdH8+0f9vJY2FP4FnH3FfBfJmaqtp40WMI0BAjtWZCmvPkeHMX3I
B5VlL1cxka2NujMWkoSBb9n7yG+IqOUMMTYfKzdyT5PiKLDSOZYq5xeR/jItEbuV4NuWUXppCFMY
FzGgsxVU/+kyamXI8jJWTEJq7f8wxhYJCMU881bGhJwrxrTHvUQI349lAyNPG6APpJLlPwZqiuj3
poXmxFnQ8sjYMzgJcu1Ld/vVCJ96m9MZunDUmMG9wE3lYF7XwUS7+Vz/c3aKtPax847c6aYt5nvS
TZ0J+lFDHl9e0kulTWYje8+/PtT+QqHJfZ+VOB7BOxIaHy3QSi7JyYghqB1QWcrJhiouA0Bz+WRz
0cwTv3DhN+iTAHDufvr1pElNfCkYUR49PDbM5D05zbpazhkkZM8hTD9lgZUOwGZAqF+Z2KiZmCZm
Ldyp7UBwk/X7k6DWuj9ldd85ILq6s1nHBoR2VVu2PRUDFWaM9mKYOSV4yZZOftzYoTvfsCRREG4G
AqypKXhcdWFxmJdhe0IljzRRiNyEMc19l4YoKpXrfUQ/aLa8gskeyU2t2ixsrjO0O7eLPYBNvbgd
VNMeO3d4hS/VJFDN63ZtSRnbc1m34l2O15TfvhPbPDOEHej1O88+HUCEGYvFbi5ngICxBZFmccXJ
IcQ7WYynwpRK2ash2wBg0E90GR8u1TYF8n9zf+TNl+431hBJOu4GFTcD5vYVy+W2q6NdJE4s2e+X
IWv6voc3Ry5d/tl85qaWBT0moWe9wadBfoh1Ovf6U/2b1SxcYs9Mx2QolRyN0Ph/7vrWCJAF04hU
veEL9KRmuWdbaPbR0xD9aKmh+xJkPp0msrwhgOCeYMUoV8to+7rO4J/530kFsAnPOiY03TqX9sfs
g+GrupSTDXH0mtdEPOrHYiZRstgayZ2aaEyuX+QbjWueZ79hh6WnWvWo2hl68xRHxjgmQctntuUp
oY3z7JHEC7Sw6v8vthek0KwQtTvAx9OeWx94+uKocQKhYdsM5WnZqCOtDaetZSEWZVW+1iStc/5q
4FV7+TLmIETGDIY5O2EVJI7wKUn9rmiR3F5aBefKpLCCv9N4PEzceOGVOf7hfOBnyDtuphT9YQR9
rghJl0tyO9QnXaNkJrXXMneXA8dgMww0JMcYpJABzT/hv3e/xwe5w1QJZsaZZScGoG7xPidJ70pb
Bua0vIMWwYdlwOALBWEvXbCD4b1yh7zrrfptaYwGuwz+eOn1gKImn9S0Zpz5oMqEv8FUeKGEYVXS
XtGvr62r5lF+EtWynYGAbRQMA9SNApc5u/NSilcHYahEjwY1VTrQEkMRxH1ELO8tpajWN0pFc1qN
4GttWpRXqhoFqfddFj3UNJb3YetauKlMfSwou2zE+6N58EJmKWOXRSm0N7FAPTUpa7jLo3lKP012
ZIhMHtX9W+YIM8Ro/TusNQBEhN4KeEOg5F73bEH0LxOu7KzPe2zhb323m67Z/YnMVRy93Sxd6fLD
d2N2ZrJ3F/vfuZZnRQ1fd0fDKupXoMEyASFMh8UOOY0rdpulLGXEk5Vlv3WC5K3sDravXARg3bWP
2abrA/DqZtg6iKM18J4f5aFurH36VSmbXU+DbMJsh+a4EkB1AcauRE3ChAkrRugolhG3c6mkrgTX
ve1fYlkmsb3sVdnLTk+fvLcybc72lOUBTrB6gXZ1twmuAcGbwe8DlwFUB6/ig81V4ZH0nPz1JFoy
9oIRdrS2f7mvhqPV0oNk1gPi/LYhbU3G774yoeegaOq152sgenOwgyCwmLlcj8AspUm83Lfq5rvS
dcoouOR76SCd2iml05Qfqd2lNcIlM8JPmJFWFlWgoxbFQDwYHzfGNI8MsGfGbK8jms47uD14aq0p
U4G71j/5tE+kXMxhzSdtaPfeZvjeLvTpaDYGc44Fb3dtX3450r2UxvrYA+2viDFogGA8g7i0eU2F
WbEEsDEPCAo1rMEgpAEqZArSctTe6JTJP6E+TfDnswJu3JpFuz1irVKiugH7JnbKq9XedgNCFnbC
XK0i2Uz9owpWskVqfIXYuP2ufPqvTUEcAz05Q1OCRDdnuWbkUELYV7r8YbzQ5U/hnlkCCMSIFG5c
iCDtt/zNo7GC2G69h+5kMlxrLp74FwgB/wf+fsy41/9ofMlSAERYLtvcgzkH1Si5HmqgLGrmoQ==
`protect end_protected

