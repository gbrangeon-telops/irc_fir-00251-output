

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
rMj+x3ocDbJ+0HvlMPtFLLYN4V3iOWmu0i3VYcvwPU8r9dUqilqv5BoOperD1z/j12cu4ait0bNC
TvgieQY6qg==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
LiFkBwHJvbvIRsrs7TuS9x+hbpgzWqPRKAN+86jD7W/DWOy2HiTI+Pr3kejl0F7PQ/wd2Tf3u0hB
l5PFI7Uciy5uXiQA7fDmYLdPcNoMNQWm9hohp6Q8wB4H3kSwMFgjlrwYcv97jBF9K/DD+f6kjMEJ
pjxxREwM6oJfyPhyhBI=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
mlNr/JQ7BAznEw9Lq2hOb9T0FUxDG5TxOJH6VJoPGS12EjdrVMK5Jwy/CrH7dSOtWY2eUHhpsxFO
HZJnPHkoY6pnOp56kFqNAyiHJP+z5BexlWOYCHMzTTDXl5ecpknkEs/jFqX2DjV6R1MuxPdeXOjM
JpDfpA+rd8xFCgAvhOcvKEKjw2lJmNukB/NqmGdLZU9Yd/iDC6mJcVuTrR2gzFDMoFjQUitH7TCG
r1krtYbVQjkm691WyHmxufh/qSc3KdzrpZqycBevqxjmEqCq0nMXCiMyQRHMFNk9XLymhnx09LIk
8Ck9EeU7sTUKIMhZ7oB9NRbr0Jmue7w3V7zoXw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
jcrZIuGwyVPSe4eEqA3CjxEN8wKBf64m71qLvmqrllZ8mLFeyFjj3f796U4fol5LeUOSCUITklpk
5B0LZiT34IugfACCFG6eSa/KnYkpqdaiyFEJag2zBthAbQTJIoKzv4hrVDSwoJffRhWS6ZAZmMOH
9HJ1Z4KODhrBj2PMMOQ=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
He/hsXsp9htM4v1ezeHFxTi8NbCInK4GRCTZh00v46syUmSwf+mXhIjhLm4sHKCSUqmWt1TLUp0m
CWcpoGxiawBF6wEpl5GgUNyVTq+T/CrlV9Oykyiw8ESh1/7hqCFXSES7D6yS14KOyEm1cr2UmC+u
X/NTzDDvOd9e5R6zaiks/z3Qdqxiq6f6jnMuQiSiMBsAMCHxpq5kEezVTATURKXvDebBjGkSTomU
Wve9JRKQPSiMHuUURnaiqzi8t62PeJzIwk64jI0DQYpuyHeGDNIZt8qQokGYPimAYp9IilmsSuGG
FM6CnM5XioVenoNWDUkk1F8M0K5I/5eHgYEnkw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 30400)
`protect data_block
4N/FPf85bA8merW49n33ELdB5S8Oz67vyUmW2ciW6AXOsCYdnqmCUCX0XXj1fIE1xsq+BM82hZPp
CPZ55+2zdoPd2bENl4u68inN/YKxa3QgdkUanFZXp38H3CXyrR7GjG+PK4GVcjdy8pP0xhmjA/wd
j1PZm949i+UC1rJnnM0bD2x1Zh6hzwMVblDLcB61p5gIRKuG73ep2Wq/n4Ck2fMZoTaxr78h97Jv
sYy7pANsnlVcMmBIH64ZV/fWZRsxc4Qf9zoBO9vvnYHYmDdUIcsxS4Sfm1qXR4bguCf8+Y/I53qL
3PbJeM54/xRmTTdLx42GwdjDiLX9MPU5yKsOgFyFdPd9HHuINVGRBe8n03Rq9qy/dU77kCZt4xIQ
zcoB8TrJ8Rm4xql8yW2AaZMG6CqqhjGuiiYw/CrE6aHbGDTLBfsGnnkJmAYdg4DkCWkMGi+D/g7l
zHncSx956HwMioo+Y+rgHgOkAths0MXKlGaeKZhSkjiCn7XduHyF42YM1JdA+DN8ioYY71WySLch
VgnlXeHtzxQaGgFI/5GHRe/ZgwCguCIkOq/iHtkm7FmRiofnkmwCPzeF6TDwcJQ+cIasn/CXd8TX
jMnQ5an+c6Hoikz+tYEtRb5xCyFysGHyNCtuGCjxiTiIB8FdNxZB3SPxrF9oZ/HwNtvZZ1MGlWCL
HyfIod4svAfKbzQUT84ZEcguedeAQF15T35sxZZcZAg2F8hPTRW7Jg+Esh3RZNbN/U3GUGGsPUsg
juhaDPL+3xmI9UgONS40fPU1ptDrqX1qwihMmTWtv1gbxSqtFwoTYffwMjfa8Tad5Z2S64Ud14Dr
O+cBHCRVyMvC66nYz/a/NLDNeC/vtEDh198ovurlnV8559Oeu1EbwHUZqBBwvgh7M4Pgtz942Ez1
wkmRXd3yy6DARi+rpixs1idZYxIoWwgWdhom0cXaXQM3WMlVizmCrJ/2mcYBRyzOoFQ4exwBwy9c
f6RHxThRaPeXy5/jw6610K6y/x9qgfmvXC4Z8sR42I++zo93Ig9t19W7Dkn6iO5bSDFZTDrUwFih
LCG/deyolhteEWd4/JXc9LWDw6q0Rm4w5jxLsvE9a+/GIV0SYev4BbMpGNMGIk+oT3L/tsq8AlfC
dBrfGqY+91OhpbEtsA961wGra3BQGj/INTrQgySQOcQ25n6keykdAg+75v59B1HGsn1a6rqnKmoL
Bs6tprIBcvkzj2tYu9Dd5p+ipaAHPziHTl/Z62MX1U/lhm+qvRYrkgHcUo+Q1AUf/tE1JWqQmpJ6
FwPTunGoJ7HEyVRA0UyH1iiS9SPK9zYp3QyLhJIXtrVGfbchZ7odeaqONg4lMG8fvHEc/uqWhCCM
xYCQawROpx5uJIk1qErJtjVkasQsDLZHOqjaJGbH3mIiJNTZF6StlK2x6470qWtNBJHCzaXPXc+k
YWFBC82OXa+UbbF0vCBrPKdzm4Eif1RkrIkz/spH30D/6Y7d5uv/3bqNuwtDabWcPK3TM7hJCQhO
VTa61DCgu70x+dUg7P911/NsuD3cgfXYh2w/no3PGAEK5gUvN5gT+urMVWFD3SefQL9dNxxsQszK
YWoBKm6oeZCjMZEvHWfRbFXyIY9ZD8O9DiKhy+Rdp6xV0O026L9jXtbK9rjxfFOQZLi9zP47EgOs
uYJFaLzmCI5QvvbFYlhCvHr3+tyUwx15Oj3LhskqbMz3jUPVV/1ZsSLpM4wQDXSo258TxuGc2J8p
NKnTcFfIymHMS5D/2pwj0TtUGWSCQ46gQrvOp++BN6DKXkNQ6LmD8l9QW/28QZ9GXGCo1/ZboiYl
37W916k6gPBwWih0k7SYfudlNTSDLU9ZqC3GwdMwhJfFIGnv0DlVsmmYQNr/lI9xnNaSok2yTszd
UfMgi5DE5kL9sk9RPPiTr5tvyqg2gEYNngyB9oqpSHZFfDFc6/hnUWZBvVYUG4lnxJ8ol0G7UIp/
nIgO/JUni8gURMkrYOvuJZbp2di+Z03kVY0DCvaZEdcpXlGwN9gtk1M+1z1FFDXbFiBGMDBMg3oO
J9o9sA+UbZZUdsjmvsugpoo9Qx9f7KAh80mMZ2+idFAcupYQrYo00N/Hjz8G//rF+40fEHv+wvRz
RP6Ta1uWpz/jaPmc9OkMOBKVTI8PrO3HVwnPbvMdCRRJXCTXoknZ8tvD1fV7PZaXmK1oizth6xUk
wX9x3KNO/kMNB06eomPHFpRWBB2aTMPGld812i9CrIKwv3RbYbZe8gycEMaMN+JeajAJd3c9cJ1b
YStweWHpZPc0aZWgLdRRT4pAestQYF59Ppa02sIBmxRVIB6D3uLWzmIUq8ckd4dJO8lzl0x9+QIR
SnJI7NpMcqD/GhawzsbqFHwhqfIVsUftMcp8DbANnxYMD7vL5gptCbkkqgqDVpprZ1/YQI8JRRQ/
emzwnKSEU74j0Dbe61kXUi+wrYRoxCnWcMdD+Rftr/b6RqPl4yY0wWyNMCjBU0E67Wln9J+R5l06
W9r85c8aEei61x4mqoHapzguv/X2HEDCmjr4H4d1JuNiDaMiacDJnMRET6bxltHhUf/n4ZdtKTAS
tPvl5LYtQ+fAIOz0mXWWluCImrxDx9EK5cTGET+IEvx7ldPULGuHCIKYhWtI5pCRHH6jRtPHAT6l
ONUKpQMc3+D9sSoTrdis/hLbBWUuB/sQH/SxMnuNdZ+VoZUNERuHcGgLGIyDiwGPEZnGzWUDOmbZ
rNRDGVq7kyIIoiwmkTpGwBfDIzC70ZjWY6kgpBpdMG9hPu9UeYrFFGzkoW6HqASpK2Gc0s6rVCtR
00NpHd8nS+ZQi7NP9+j30J5crs2xS90ORDXq/AJ3PvRV9/ZEX7crto8lFsDCXQTlNVr/TP0w2bUF
C3mtDEeRJKLR7iIEVv+P/zOaY/jGCflfr4XeqrKwU6D835gLRKrX+eP+Rv2puvBSGWBPABXnhhua
s5Guj4V3j9Z3+tvAbA2pNrhvv09gO81RUOD0feuEB0EVBGpdJLW2zbps9yqt37Toq0Y9eSdOBgME
ya/VWH/DhmNGHbmdKX7sgUO/FhjdVOKUUirvpg2/K1j1mNel44i4WIXs8UcDmi2Z1onsc2bOPOgY
Q3u2xXeGlAnyHr9//u1NFfcUkVJB6ekW0MZv+eYPOjdVryT2ls9gbyEBXG8tBrGTvUd0UJ4QfABx
oL87Jc2EjkEhyLdCh+TFbhYQjRgXYtcG9ag37yHVimh/gEn1aO+l6TGbJy2baVEuTKbvrbmLsik1
97yqfroA2kYbtcKW3fFeib3Hi90zw/DTQG2/bF8HIu40fJJ2xis0cVMM18IBGqLBEV2t7Ko+5KxA
w1KfHoiNc83ZeBuN9GVRCs0r5Dp1MqDFG0vP2LphKTcaUGeiZ8jV/DX8o+aNBTuDIJyW6nGmjvp1
HE2E90FvrhhTtc/PBQVNAkFJXvOA8pokiGlOLBLgzcAAozGWXR188NUQeG+ldaSXPk2Lm9tKM1kH
lIuJaUGmkUGXF5fjlbZzNOclNKH/+F2j7nzKLKzHJ7oSO5w9amrWPscXqCSUk6XusV0U8wYukWP8
f2ZN4iL8OMn+nJbKyFbXp5ueCoo1U8nAznpmxL9XlMcU5WIDs2NXsQlgCwvI4nQRWtdsMcxRsrvu
u+LJQOJoUTKuskrKDBVAT+cGf0mXxnTuOB760z3NEKjt36K9Fp4w0OpG37U+NEMddvam6DKOObmH
yaOKneVCZvH7h3wOASkjDn67SCwP8AgdJQrKzBqU6nKnINheR6hp2inaMjCU8Xd6M8SvFqRWq+DA
Znoj7clPfNomdc8kawbKHgJgUboUhu3BVyRQ3ZZbgyLS6u9bDsh0QcyTwCMvhafVapLo3Tz4zBpc
/aOrgwUpUFGsS6XasJb1z4tyJK7yxyCVlxfqB9In2dOroYL7S+rgIwsy1qKNKQcQl6dqDehQ0w4L
iCWICVv6DhiTBcjl5/HBmAjmY06YiWhPoV2eQiDrkwFSkg7j0jToXHyRKWWnk9sqw8nJcLcf4ZPd
3+/72VVbWtmZ3k3an3MLQYjADvpCxONnjOo8vNo9aUFOePgQckYL81n8NZiu6SzvNirkR6EmbutP
O0FGtBY9FuKNYhHAN487kX4tun8TpN2cm8uXbxXi+jnk83GCl3eHegog8BaVESB0E7LziqeTM+z+
DJ81lpp5bop4lvQclHgNOVgh43kftqWlKBINCo53nLvv+OmMqu1wm37CKNq0gKW5zmGHWjbqfeDF
4fJIVC0wPi/Ow+vsf544LTBFTNg/6JgTDkK752208NV89Gk1pb4o+P0IH+6k19sF3On721np2sqG
/ExUx6Sd141KHwVXDqUWTmVt3TTfhaT2bkOJSp4zwzHvcE4VFmt4Esj/1LMmvtKB28wnHzVsn8Nj
auhy06JsZ5knA03p4tWSQf5GYJXKQ5QJhDfsmxbEcy4FTrKRsZ3MwnFRyAaOZE9RjBelVMhb1NCA
XsSJgqrX8VlhV2Cdnq2JvUHM00Yt5UM4MUYKmvLjFux1SqXUChaE3+8w6vLuGIGhgGRT7iI7gdDD
5Ahz5lXSXqXpTlRLX0N2Cx0Mcdsygd/R+qsAqTwbTkasDdGmBYS9hW/tRFEaQ/J0mE+bMLrqMDa7
/c5UD6z8b4AnQlXgGBHiOCr+1CbLRmmFibkdlpx2HqUVu8DMBN4wgSzwkfpM1tW1/lttGlXeqzV+
zpgwNAyhIh1XfANc1Lv2fHMsFN/jOU0IML86Ez/YagXXVCHOM+xfTukp9XTQHznD1JOkqtLq0kzU
ZVpDHWlbfGQGLnFRxMdYre0FlwlHpfkpn1l5OggkA7kby52CRMtJ9hYwXt0c5gItzKD20B+liebl
OaFluHeA1fSL+iejESc4v3P83QEKWnwYdJHVgeFfXAHdeF3cFmIlA4Kce2VQ+YboUqk0tzpGGilh
Gdz3+meoaDY3bixBhffDQv6xL3JoNHqEHKghcwq91EAy9U2EAT+xQyJFaqMmpEdmccgmvJTp9554
Mf56zW+DHLCJN2m5T/2lxq954f5JwC/1bo4+N0/6OJ0PtJJfGEp70s+s9341FsqBPfwyD4JfF3Wg
l08gR6e80blZNyeBHcna1n0vLuZmWB6RF6sGp1Ej9Az7gsyqmrdslsrs/3+OxKTkQIDHx8wv9r3Y
FzjAhnHrhydwJTplxmwtBdQmbEXcFEcMSrKUbmOm0AZywq00fUKMZs3+rWE0vdaTAVW47VxZPTjr
K7VFrPeoHKhCApIpEy6V5oSE+As66sqFvrav3wNmt9pAldvWCEf8aWyjKMOkRvU84slOTwIZ6wLK
22nijLXfxDIOcjSLhHHqnaVvtPa0f0Z9HvvLrO8niwEirKXkn6BEE3kEwHb0mJsSe1uETVoNzHdb
KuQ++/7+TalSg+uFLsM6iJcZM6L53amitbUBHAjSoRoyMWT5hCZBB9Ljk44f5Rd/ZWD9kJnE4Qgx
sEfftSN/KeNZsLVVVOzGspfukyKtcNjnAkGV3FWMNCIS9oQldIVc34iKhw0x4OkobNNgdvGC6Jcs
cK3e63xtNaW7PB2m4mhA9b0eDVmhv2zic39ODdLrd+Y996d44J/2WxfT5qy4snDsGN9wxNUxSroX
vgXrfBE3dKFFT+F6H75LT9VxcJktoWZ76kcL6fIols/YVFBtfeBosnA95ry8Q54GVrxi8ctoDspz
KUGp/gkcGookJPnmeZ8eoDwC83hzwJIBjR3Bgqy69BWp/irPJjLHnvxklQ4ptGgH3zEx6iJRRXjS
/sSbwy6jTxx5/W30AZHKTthKoqNADCR6iCJ6hrA0r7NgAeLNoTZJTOLe5j90eqB/TyhW8dSCg1aZ
m0lgGEU++r4k3g6GzeWJITxF/5/l7mu1RWSMy7YYv8jjFwHIN//6yxKDa6e/OYRqWWNCOq2nx6Fq
ZNopyjZ45fzjBhHtYcoGTK0WbLKZ1cd/pAC2XI37gZGwuZgHPZhnByK6KBY9hsULbg8y0cjc866w
A+YdSgQvLVf/btgv9gy+/8LCBC4NvYES0TqC8REERx3onU5KIZIrTL6x0o0Wo3bAgrzY7SlyIgpZ
Ns8TvksgsWYLeRAYcD+BRn9KWTSFby5j9cGHuejj4ZiU4H+8SaMk3bEDMTYG47YTYko9NKDkCh7j
Hc70InzRz/l8tXSqsaM0a5lqnX0mUmEd/M0QiXFToTBVQcNqy0Zp9f9WD/0QFpG0SLp4UlDYItfn
B0E1BEeGZLcgAL1o4QJnSCcU7EjmqXJhiX8RI0orgZ36OHZMCK8qCClZGF67g4N7/ricLyEWPbW7
c1HnJvHnkngAb1mz2IA3ByC7c0Fu4hZc81jD06FFrsf7E8KJImKc5y5VLnV4nLnT11Li8JXeC+oH
AMwJ8SPf5zkoG7BiZpPCWCsNzfV8NrtCqQ0V7zait5QtlSoR9BgtpuBGlbG3PwOyeRCzpa3MzDBa
mp7ov1MixMuBQJWSA3j4UgNMjBVqk6B75LbMzqpdqe2m0FP1Q70jACl/hiVGinrVY6qUB+46Bn+y
wFDcKAvsc6nIS5iNlQSJGJFhxM4flyuqRkW6WrJNx6l3dEfWGFGVSH/tOYIMdcOTEmITsP8TTLP3
yjr0jcSdP6ZAQ+t0OUj8NCezYqpeSVBmoOAde77iecDySpihyqnRR6DQzZTysNrVYLewKbfEPcJF
iREGPOXA3U1NGlPpX5jBf23VHQgaeJ7gFBP4Okqk4OgWou76VbDxvDxEdC36Kb/qfscIGeINeJwS
ihCgygS35Awd3VzWYIBPc97K8Pgm1ooqCE2xV3Blo5Vj8KqIP8yJt51g0Ow7wgdN2/0cdc2utJ4g
P5NB4A15ZYSnswh3sQCqXqnGcoiI9RZzUvieQCFpXf4Qeksgl18Y7ul/BL/14QBeRkhys67vE/KB
nukhf7HyWlg9l3CnchA2LDJh5gQdxJrQuxT5YYOF1zcip0N4vuMRZyXIsaZVwzehRAlclYbE2Sax
6SsQ2CcHsPKoe17yGR0DwhiFZ5NMEOzkfM4DdY7lpXIEAPeZmMSSOASXlrccEo8a13hUrIP8fcHB
iPO0PiUsAhVIiszyE/dtydBkjLRLWjJdbVoXjxR6z7oO5ewa/745yXMFmdxfjn/Xefe5tUq91w8c
fZ6ETe8OlMHmY9E6jWGdTKUPPTZGmt4oIehA1xZmAeDjoc5x3aBoUiIOH+BjUknfcuLBCL1ax0Qx
uFnI1cuPsmNqe6RkuiRwhvB+g/P0douYpORWu01yzuLcVySCxnzKGBBFIfX5MH3QLm4eL6d4Nyl+
89P3fonFhMqByHUi1CAYoajwfkOgt1D8YduA3ikW3FaFletF6Xga3an1gHq3iqrDIFuQ/0cWQRHA
QIAwmBUi05wRbx0iZtxF+83HqzxhmBqc1tW5v4GgdDMWi8uUuP8GQFfD+a3ciM+KD9B2r7j1jmbB
KmdTY70mrDyzO36uJcwr8TONnQqBbriFZflfHntwRWc6rbvV7NpE0KqQDb24Mn4zCo49hACzG43r
YF71ABb/iFiNj6mIZ7PdfYug2u+737wyjp93BJM5PmdIW91ZeP5ty40ZDeMi/jT12N8tryLFr5NH
XkLyb4UjmoS1S11rtoBvHOwmW0c3xpnxHSG9i/oFClmTVwTHfQ3yx/aw0rZqXJzMO18UA1LXNAbp
VEH2DuVqY1H1fNXsr52+Fu/ExjY/goOoBQfqDApLBH+iukwgGMGlJ0wR67l8n/Ydj285haRqUco8
eyOC4Nx5Fdg7DV2VMaAgy4PgdGO2Zo/xs+Yq4pvVvUPF3Po65A8zOFmjZYYKKEmum2Qfur7DjhsJ
yRyEe6ezkR9xXUnRlqanycQhneNRRaW3kzTO65EI0bc2P9hf92F24VAnKS63LsqP5yAm7jKMcKEF
X8DbBoO8xA5jkcW4rCXYe8rHnjo2LR0r7+KKbxo9T9ReHmAQcOoeKB/wik1ah+QDD6ueqIDPker2
B9g3r+FrPK/+0dwfEzl2FfYg0yD7NyfKY6mPvQS9C60XR++Yn9vMqOD7vkvYA4QPEl3UgRGeQzce
rsBHgo35U60j7Kx5KpuIiO0tWoZpZDOdgwlFNLsQupcg/org7ga3lGLwnbJaD3Y75XLZGir/6MaZ
d9DqBStnAVjAKCjXTlLLCpIQ+JVvSXuEQR8dMOmgK7PnAMrH+hKU3mU8HNKTuyiKTaAaD86TjphR
crP3QCEm85KrY8uazdRWptKSzdB0siT/MqcElR4EcGLK66g5dhtcQZeZ227hB7/APPtEUsj8oISt
atc+w0dIZCHZPGKRy2ngfjw2DIJj3GH6NNSaZRvd97lPmTwh04XNYBg0hGcaLEb1wH6ojiKajWZP
uNZsHzwkme0mPYGHSqVfuIFsB+GXXM4FgC5Bj7uPV694QWo67Plo8i1YPJelM+y0QIUFgaiKqteS
uS1Lt87ab9U5s6FdsVIRjyvXIdyWsdXgWygD8W8M40dGnr3e93ZQ270FVsGBWd2FD/wJWLePKA0A
l8F8zoqD8LZ2lj5hcadX/+2bja8Ms8Fdylg88O1qMvcGWIar83NiXUSNUnlUEP0VWvIOMlHQZsnI
AQf3R8fX9iEorwXFz3O6ZtDYwv5eZ+xN9JztTVCpua2XDLzNSJvVva+UxBgOdDdB7JniprCVrKYN
HEaD0RcM5EdYaafArOHyPEAfjTugWiOwQLzRSjdV7jIfG5RrMqh3n/N7FNnrCRcQCXco/gBpBWKh
3iohhq/XTFuql7vuXuHYH3kWPoHW3LNTKaY2uT8Kx7vVFaABnaM0a2q06PzyJJRz3uvdblGgWU7x
0LVm49ktK8GIS/jzL1++Zf+msGp231R9iBbjJEt2H+e2CaTSJNuvNPM/hyCKCbT6IpmIvOVZY2Hu
57I1zKFsiez1ughH1Wkjbz/fl+VnzH/2KEP3LZGEui9H9sEtMDiM2ytNDrlyavJRtAfMjF+rbau2
q3Yfkgykw3SIi0wNCyySuQ6xGZ5GO2M3CYEdmqNX16fq+OajcvbUHM1NhzbQsU4mx6WRClSGxvWZ
la1XsBkY5GhpgXGRiWbkiXm/OmIMsYqu79in4XloxKW7KzKahDXKTp7J+Te1ES1QO85LCjFVQs7e
soh50ayAWfnDMH7XFxNJFbfRH7EiR1lRQUwUpJT8kz5uokMf+cNMlkqLt2FY4jKZp9KRdOmsgyOy
9FQ86tnAEj8X1CILz8Z3IlkJ1hTYnYFPY0nNG5nPvpYLzvWgwOlKwkU3J1oTFUTCVQI7PXy8enOD
khcRjtSB1EnZRLJKKR50Z5A1DOQLLvtMMMAnZqXYI51iXvaZ+hfABiH9kzCJ7pbLGJTrF/BrESL+
u1ZRjEbn9i9Ig7wLkP7nywUwv4ZizrRlLFp9Lqy/jwQWOh9q3Tgw+LpmOxTQKgP8SIrwmMEdNs1z
dCCt7tyBOQflbFHE9/EyKZKC136s5VV2Ch00fHJ6oyjy5Jaw+7xgfbkKrOSXw/qx/Dy2J8snYNvb
p0hdDTTg10voeqMQ1kO5VVzFAdgZCLKrZx0szKA2BYfH7CYeo9RhelzBqKCaZZDa+xZxeds4ONUb
6dGPIxz//6MxJndYQOCpCLi6iiaSkg9/B/tQE9KM48lqYu5RPRmwpEg5RV4GYKjMlzGrRfANHgas
tZ30ySfKh7wO1l1mIiakw9NdHtc3jnvStMNx9BtpJg1eERm4O4kf5NlAdOqv62jQklAUfO+du4th
B2xF72okTMV2JYwFa19WyFCE5fmStSgFkTG14zWlBkB9CjFqG2HmWpKXG06Zi1K9+S0656EZysik
uTTxXRArFwrzcxvBtS2vNlzVeiODprOMtvNJ1sAfo44B7ZB2/65mI24mp8nOdgdM7lTFf94N6X8I
CJbCuODo72DZ25JiV8FLuE0LO8eP0dgVDqHkJouvAsLFoxmzjtRKnfjtFv0Vcr9P59UUJ8gvKxl9
+oMB5mogVXKWVLWgd9xzG0kfgSnPOaEPVdgnakA5QuEIGg3VUBq5PzT43K78RE4frqVUNTFn1M//
hZd5ecX1eiZh747X5KCsFNhO2e1MulkZ84VGKAeklL6ohfoO6t61WdfzT0T9vw9A8uohcjQ0jPTO
642G6rzYecPOEe/ycecw7bEXEDYTw+EZmEWtqevT42FfjNif95RDreod3Gif8rUrwnd4IxspTCzZ
8sG+T8UoVDg4l4dShJwigsz4544+36ICtYBWI+BcwH8AAJkcKoznAEOGagRZZpy9YcuX9o+CfyGH
R5C3RRs/KKP5Vr2j3ekTZNRNUBXcoQJZ2Z1z3kOu3tOxyt5KZocBr6345zAloic492/7O1TnYOy8
TD/uwN3WJsPdiyfmNZc4J/o4qoDsj0hsoqZoRRI1j4osceeaTnsmoAN6IXslr7OEsuzFnQA+VWzg
vDuwNFWPlHSsOvzz99LKI2l4TeD5r3Kg8vqVQ+l2IQecHBBdOA6Nm3rEtsyxksJ0dK/ZFn7YHKaI
FIfDbw4/3g0S34wcRe5OC5wHurvZ2ooYeROe0QmWY9Fy3r40FpqKou8AD9ptl/jemsNQ3xEmz7Rf
I8xZODfOKvTsoKCz0+k+L3sZBA4ciL9qN5GbNC2QTFzNU+rgBXahkooBAjPWZnbCHBbXm3cBU11f
PTANcjZwFYo8vT6AYhkKQOUlSiZAcNIOtvYVGNe4XaWAbqjG6mTIJcQ3CCx0cF7TsnGQES5lBqV/
0D2U21N6y1Z5mh5dE1eA6i5itHmiRf+R4EaFQAYAVs7zW04euucUDaPUCcpAnFGx66i414h5Ml/y
SA5Cuw2fw+w8R7Qmk2ecpZxI6Q9wZ+jFqiVBz8a821AOPVayk+C/hGMBrJnDVBQ+NC9ZreXDABjH
KZEW6lKl5wHGY+wZqqx4bayZ/QmxQBc2SmdmQb2ZNRFg6VP1Y2wqVxr9YIa+HEF5+SiBMEZuzcFg
zKFzktMGtjvzg8VtfmuIM5p2UGiU2LV/SMNXYacUjiNYQAmDBwSS/gs0+j3F+j7hz9/5oLeXWuZe
tLEIYbkvJDQ3EvVpYGqW501IWhhgzy3EOe1TxCS14It6YoAQn1+WgQ7daS+SlcyP0xoRQzNu0say
Y4nM91wOxemmZ3oEh0zfMioWFUpMpS+rd2NYeMpM6j3CKITkN/QXHUfQzeKOPfGq8sbu1QahWOfc
q8Ht5EA6YOAjJZs2mx+doIup9NPY7oxEeG+R7Rbvhi1YWtppodYIqKye7426B7UpwYjP/0HngUgW
dGPk9kwVsN+Vgk22G9k5SaLzzF+hfy4ag5BRgVkgtT4IbJQxCIrACfS2Qq1SVvr9y+2H2Gc/EB1T
8AMg3ANm1iFZlmHzTjEMhczQCKIaU7wNcaCjPpfNjcwvspx7XNKH7Pv9mBS6AYor2g6WpD33RNz3
1UUBr+8X+vIGFqmMESGtqfna20VT4mLQop4ra61cgSFYoqj9c6BBjrqJKIGdqovXmK5YUKi2H6UI
7wxnpGoUXBaHBY0anz5GDNuNcY94gWIxAJSCvFGn3NpdHV08Qdyo1Jg5zVbd53FPCSRxuQ7ApPp0
n/i5pIt2ldA9dOSzxEHZzAJwM96jcLF89WS8/c0HNnGKarvuJf6b7b5LIOsVBt5KsKmbso/HUjU/
mVVka6mVFIyjpIc1mRPIdgNeFja07LM9TUibBtflTQxg6B7HeC7Fxpdbti7awaEYXD7kTGbiu4Hs
qpCoZtxHIhu7crjqR6drah2Vht3g0FTsFJc46nZSAayfFNQMUnB95GrKdYnx5QhL6rNi9pKH8o+g
QTTGF7GgiXtgW1bfNfGKl2QsmWEyRG9lyDTMZLdnAYUfHwl4j8Y0FxNf5Vnd3hMtrMMjXz9vAt2X
nycTEfoLJxP2OQNYMc5XMmhoMGHpsBMUcgmGofr8rrp5zfVnRESQ36m1/b37xXsEZH2QZtAGJdvG
FI1xN3NGXqU3bXZz9yZ6GmmsXiXqUqgiG5kzYgGSxy5xyTvhRGk/Mmdm/IM7NvpImEornxLcFbEs
vPmyXb9UgtSIDy7kKz57e88QkiwApMHXSlvmz37lXIARThNvD0uNxKi4LbWg2ChwppIh8jY1IVJ1
cWRz5b3ojgLQca+tGof2hfhME5F4hD3HjKcmTb8zZh6xmhXy0oN9PwAjaJB5yNPJTfDhzIuTEv1S
Iz8eNWTGSvu3+9vHULAh4WpsjuoWXrbg0nZBjTE5llhUtr/wtU6ZeJujPvw7rcTC6tZLk/3J6xl4
p3J/57LUZNj1Hn/GngkHVikTZrDaidI9lF7MIsPIpfs0rBvcJB1Scj8r1ad8jr/DDoQBhWQMfqPw
4Rc7uMzw1IqFv297ul6E5omQKIIYdiUeL17oYZSDB6dYvWzTXB8OVMYz+HzxBbVcG6bvh+8D/6/K
2YkA7aEsGiIpnULX7gdzmaoLwZNSxVezxUeC7bCdWypRhnVpZEH2FC0g/J5EaaVwoH1qjwCNKBAs
qAIKsxh3td+RYimusNqDgVuiROZrLL+Pi2nbw/P8aNOSL2H5yuLbwFoQI7UVbagMWkf+Q+rnJ1cc
pNQwn0C0G8MOxnxa4l0MecMwFX2Ufs/CON4f+REnRt/yO0317IM36hz/3sZ/hVwzIeMeEwZmJm+A
1/0zVxfCe3Im3CF0WG80SQSSb1udHz35vObVpoZ9Ea/5AZudf/s1oIbhm8H8Xn8NSzRgfpdNVAHM
+/spg0DE9HePmY7Ly7ZBKfNJRkxFfnNP4TWpczy+2KLJTvtrLNFy5EC0AW/yH8BSV0gYCIEBJWwr
DsnhMAo/v6Tz1VrC89eApI9yPPN9ivaElaai5xghvPxoFFPmHNz1vUX9uqGWyvf3sdbSToB+nsxm
/H+GghkveH2AgGs60h4uQzglr6i9VjcJiP/4OiveSJsY4XgLobS8XurYDRFOGSuaeNDhr1aNuZQ6
Nrj/zpQaAI6+VyAfDizVPz+KOhHEVUOGJ17A5TCAf9QOAkfJ+O6p3j4u/raVZqUhNQ8/Hnugg2QQ
ljKG1NkUdLk8JwY6t9jEuoo3E8B/WobxfZ20Ll2dfPegqq7wXaS/RrwBmzGDausbHaYAeafbkE1o
mwwlSpxcigZ+19sf2Wgt+bJ0XRztty6ziorGFo7a0gROyTszcbrLlnAentaz6VGXc3BCUHDibY6y
O3RaGyFFQPy7hA0N/07Anezh2vkoTN11JX0/znfAg7Yz66fMr6EwtfJX33Kd1iKiJfNLGU+zsvkH
hDrnZ4BbwsUt0kWEMmAcalCuAoFhCp3vFZg7EPtdzB6hQFuLDRVZqOd6thXxGKjsyuNJvLNr05KJ
qdQAVOWHDWzmeLoHkWx7zFSNIPeZh9s4T5ux3NFw5b+PKCReA99YNfLebYh5l4lpvNnRVAnHBHUx
W+5LqeyagGaAUVf7uvPOLXBOzjJ+/gCey+dPO+O+yDieXt0TuCC9F/zI56MsRGSV5JiPSI5vWeOS
g7hBpcMo70+BpMa1b+4oHgieIUnHI+x+L18vEZqbFdPxjvy37LCXn+7IG0hIYfp/HhrWe1Sxxn9I
1j5ZlIEoiAgzl7geFD7kRcyjekvxqy1ncOPnULoN6Rvf9KUV+sirLmzrB1kh+/xn4xTm7T7ee4vQ
SUHSxkxOy3cGJLKxYZ3iCRF+ZVfJ4u93lupj3VpQ+XQoZd7uB4PhDuLzHMqc3+Y7MCH51wF73E3S
EdrxPaW/K+nXAPA5ILci2pFcbTAWwHwRQlPmG+aJw+wUKoEJKoMvxchoCLsO9VUnZfple4uw1LS5
BKCOjxR2Bg93cX5LjimaG+ugmvnUhxA7HWvuuIZ+GkycysAIWOXZQd+gNezM5AjxQcBFXjP4UxHP
nyyWRGAIPrF+754yBhbBPq6l0y0h5cRtYwmGfEupb6gnvSi+dWvB2zPB9c8qXMqcNYsNqyeiTgyZ
TVeBkctR4L7xvs+n/Pm1FkJ2btLw4gWk53An5Xvu1Q25VkOHJ+OW2orf+6cJYb+CGObZMMb/wzmn
jOCJ5mSLc0zQEJtDF7HVq+GHTcBKyra4ToEavIAAWH83tpnqj6SwbPzZZdEKPP9xGmSxUYZ4d/Cw
POLsRoVuAaeH8HtclCDbFSHAy2ijoH7hVcTiKzNqZ3lc9S2Vl0EpyaHL4Vxpu9tk5CL3C5NuCskO
mQU6xetzRwzVeVA/B2rZXmfzWWu19e/85zYXLS9THu6f52cp5gS9guyG3w41AOL0abZfLlM1YrtI
77if9INKZknKFoS7y3IkK7N7iHEoyB0qOL742GynLeb5bF5Bph7hYc+RnxlQwccG4SnWcogRcJu1
q4qpw+Ui9FB2B/mPF0aBPWh981QhiQjXf53tMK/hOVYJ6VwBfxHL7lvreZ5yud3srHVkrGAlu6XL
HU4UB5U059a8F723ppTyUgp44RVQhpw1qo0ezHoqUQHiLuYvOoqxiGh+nu8p/9aU1isziU+MqVn+
Q4t1FKMn3Ii0GlworqxxT30K+1PJKrVkZWRUayAN6WOfS2fN+ayTkQvtareqmT7EUAcBoAwbqydm
mMIXYYP/ON8DedWUn/aDGtJ0UsbvIhqa+VlOtEEOOG/Kcu/pK0YuB0MeZ1IsFbrQYjmh3CoSnTbl
0AtmxBhDucCGf21RE1sYyaIcK2rji9m9F6Hy5vjxYgLQhL+iDBOHOp3bC2FEfzvRPtu0uAwAhkK7
plUt/fsV6glRETkkZeyqYqEKLf2NECQn6a1TzrHuSEiHzXyM04af2CMjUoEUBxiej80rZ8tL8b0w
Vgy+TjfvFjdPnhS4j5anO398wH7t8kAWqAu5iFGX9iio+AEyMcEZsSL0fWi0QtTmQ4SInzAb0I/Y
ECa5u3FM/7IzxQ2w+CvuWhAUz+jxTXPB76MniLNGddnyHeryzj93HXZrkKE+6bjoPAVQwfdLMAuV
nfJjzgqhGnxW15WQD8VwWosJInVuwOxM45toO/fqzztMT+8vRLzd/7jO5zsIcypX1s3DHHy/tbx3
3K2FtT5oX8u6HmxzbqtiTDDcF83VWYRCARRmdjSkEuba7p2EQ9Bgq52sOc5m1UN18EkyfQtsvSeb
PuadT2Ejp1j7RNueYTeeWdrEZsb43Iv1L61ta1q+ioH8ZkVHAKVvnPSZeHgqb6ercoBLZlUxasxV
KjqiW9TwyUchQ5amLYOvZ3jCRaZ8k0tD1DSP0Hv9GD8x4iWGKp9dps2ezoJf1vdn5y1KmzeE7meG
QwPhVJrVO9aGriXJ4yGoy3Zr/a7nxJ/D4XOt9FG7SzvuSzvIpnxcdy1Iak6cisMbMbTEnaExpCC5
zLBGq/F57WOA0GjFezwxhmf7sReRlRIUA4CAl+0nfA33g8HZk6aoAkrI7QqFmNhLDG80wwBUPSg9
1K7/fCtRYVCfjMJwm1OdJduNz/0xHDlQI6qaYE5tc/Rjg5ZtMjuAG6DR0/TfAJNCkK5P1VsxtPci
wqx4UdH8x4fCowKx37NKVctMcpXoUBF4Actt+/44jD79C01p+FZ1+OkZGbQ/sVkOSDcjjNkXMc59
UCvzZmOPHPQdylasVk/EAO9lvwA8tlkYFWPXQrEK6UJQqBwk1lkZve6tOqKEs5FPdzqttfV23Z4M
q1zDUUazPmNSPrbdfO5mePpcAcD2Tuzxl77CUgOfHiE2ybgfrrze/bvbbNtVGTiAwa+E0UUvoS6Z
iFoUQ/o+m4t89sJXaOIAkLW1DKwK+qE6fSiswFW92EtkwqxZgkoBKOBmBck/tjb0L6kfeBwHi/2M
w6Wb1aGq2QpS37ZiX02zY6HPKMNscQNMtFtO2OSSWk+X9xaPpIImsZ1WLJjLiTWEvsLRBVDuoDcR
iJlvFRRDgrR5Rw4tRzQ8t/eosCmWnjGpStwbBG4f5T24e9vjTNAQcgnPl9fAUdbp7zvDf6r5rMiD
QrYPJq0TwMhMNDRF8rgYajWYA/upfWAs+duLATqi8Xpk7Kb4dos62LzC7wUdZfaPcU5oHyu903vc
owO5AZivyqYS00DDRFfAJnn2rQ3FTcTLA2ldIPLpKKxjoJgWlWjgZxaaNDOG8pc/Mu1oS/6/S0Yg
fSYFZHPcRUbEyuz4eZQj+pjQD/+EkcyC6czCOrH/FfU2n6H+EWaxZorTjJ4+fO+bLLqCco7s/MkN
3KyZSxbX/GA151IB6qkofkIMFvFzSk87zgW60nln6tA2+qAhlTQqHUGEd8PdIMZJ/mixf9ux53oI
/Ffdw9t6iHzfVOB7InRyu7sDFRl1s7iNZW6tBtu1awRzTZ2huMIm+rrHbv6RfvQpmEk0qUW15yPP
lqD3RqGlC9AzbTxOkprY68yCOcHFiJmeoZ5vyt2FP4yvzIXB4xZenUAjEdxbKgLwaE+o7qhAmTCQ
Q8WM8T6QypN5E6IUYxeqt2nPv6u5APd2YWH+LV7dXG7lWQdAs5EVdD/ZvAgjq2M4NIwIwIDkkxbw
odBfWtJ4u+eRy3A7rQdFlsUQd6foRBoaC+sMMmO0WGsB/RoNj6/JJpTz0IfIm8ncm5WkxgZ6Yay7
7NRcXH9yFqokaT+xYC4ebap0pcTakyFxnlgu602OQ3Ps94sMoTLNV9fqMHbppxogmB7w7eigbCGn
L/RRlX2Ii/VjHCpKeBj7ZEehhIg7O75uLbF+qqQWkH9LM6n3cXvlJpqqzEkCsHMapDZSxa7rPgaN
ImbxJQoeM6OKfSs8jrC8Vg1syWvD7e+2FwTVIDTZu5OWCalt/zbfK3xH+K9gq9Fc+kYFJluKeRA9
swh/akVOUjYLTPU7nnwJpyA4ubfFqBmuQwa+jWE7z1lUtjGtPPYVTvKQQocngsWgla1yqUYcau6r
QS4GebsX8gbr/NhvacRr5yQkgDvPXgQDsrrWI5iIWrVtHXXFoO74+Hcsmxd6YUD3P8C0WQjTUf3L
SaU4+mpGgWqujuZbwoi7PlJCkmctr6AHuNBnJ57mr0WV/1/KFbb/o8d4hp2fBtFBjbkcZePXwNIV
R5uMN46BSUfXYvW6J7xO2BVUBvdWqRxh/Hucn0huUotWj1EBVPR/x8oS3At2MnZHlmqEu5/WbI07
F0vM7iKQBCV59ymcfRMegujy09SFlacCCVJVkJlM3ouVLYgQ02wSqfuQbCu6MEawszGEmaTzkMbQ
q04CdEB9LL2r7gK9AYzKbu2dgwf+60hj49a3QfR0jqDBLjkFDqlYRswxTzqGLIoOV3z/Fir1rNt+
jsVdDIaz5YSXKw/Owwfsb1fcGs+dZ+JuBCj17J2HFTodLF0B7QW/RdkRTNW+oeyjWicRR7AXQbq3
qhPz5aDR7QQJbHQv/acrhWCyJenz8dV3aMZZkaHRWE2Sz5uy7gm89KYI1v0P6LRMWUUV+NpwGt2I
VIn0ZiNkLqxbw59zWClVRgr2EoRNsK0PRylDEHqn0EMixvfPI8MW2DapCKkoL3U0rfktc1itMjhl
Scrp0xOteWWXhSYYQ5F2FoHEVAUVZKiHoVJ2WGgOp8LFIbMeY9uYzZY/dcCy4e/8lLmG92SRGDr3
nnba+dc6oh1miOueSVvf0STHsepQOGWVi9HkYobeEcEbReUQH5gMJsdTNZob3s/1wFM4pyUDrZbz
gfJSsmEXsGgkMQdK3+y0rHIWB3cbpJCiByBVyrF9mkG9Qk5CQFOtCaRlw5qfRN7Urv5o0S8BG+x0
p+8yoeQsxST/5xv1XdcCoAOR0R6gVMDGhttQUFfM5ETGb0hJoAC/XpPS7a8sH+4Si0AT0vbOD/B8
UkbBCPiYa9cq+GOel2MM4YVDQQhOvcIoJB1i+Pz8BcnEw6QrMfn1J68z4IouHO73sNFOjLpNSmOp
5WexlmMStEzW4oifOcKMECYRSPQZrcO/4318fLXtD5ehFRwNJ9F/wviIMJRg55Q2V88vwW7UpUWs
ecMP/dKmqIb3SeA64OvxC7Uhf270wvTv/rirMHByK4LXMJ3aI6IqWrv2IZOu++xdJppi+GgpaIEW
FdezRL8JEZkgZUxEy8EbBXdbil+8iivsOv3la/7is8rrTdCBddqkdWJVU98DOvKWBn4e5gQJloAN
kv6RIdBO+AHLjYeRSFCyCjMVbwj75hIfrgZ6W2NhRVBodcoj9+nwXLPZiKzun5NHl8uynzDYM1OU
9SCye40AjoUM2nn4Xt308Hhq7FAaRX/OLWqYUgrEAiBV903xwuHdSkOKM8OkZo2Kqcq1vbP3gOVc
jN+fGchlSWdNU7UxCXCgH4hyAlFGI0CIEx7SS+q5GxBQE83erB5uDYP2YIWtVh3NQZQ9uiI/VpOL
vThdfGNts5AyWbhBruXoZw+lTNDVX7QKKCDJhLvMRsI3iFb+xM48LJIlkFFrD5sfalM2BwI4gaUW
UnMy78iwJZ+jHmpkNROhlo1lVzPQeouth3rRqrWVDxnIwgtDln9GT2MHoZkRCYrEyu3KQW0J4wUD
a3bNFYqQWBw7LlRHBGda/7CCaWukDRyvQv6dxsKKdOeTjnK5VvXtkMk/9trbdV4gnjH7Jdp9zUrj
7kSJ5GZGWrV0zoP/fqt/ToNlHF+62LFWNec5DCKTA4192EI47rWBXwVEKP8DOJEHKxfPyStp8pVB
3qNMOV3co29F0wn1lWw6tXseUDsL6xhMcANDwF1Zh+7v1x4OHQEatdJxWS3lAKEaKBISVB/11gZY
NWIGVE9Tn4kzv7UoaTz4MRfS7ANl6B9MIqsCDMF8L4ExtibWh67kToR2nDJ5OxdxkGiTux2eX9RT
NeRVrmmzOGnl1ZBJPZLDJoXN5wzuAU3wBIeT4wvBGRSBDNJ3v9cQaIK4DrmiYLWf/5r8fkrdxfJA
siZhEyaauARrx+0OIVfThEntroXshihhIpNuO6REb38mzRnI8mSPySUCB6e/2THQvo0YSbF7FBx4
bmp/m0vHiZ4fpt0bYLAYa4pvY/7hGiTflqDpw45OdA3wRQ07jwgBF9onCaJCNjVIAKgyGhlt/E8N
zGQ4NaGMs2IhPF4wKV/b7LkXKUT1jkfrmQEn3N95M4JhByPc/5d1hiMF6e+1zGx8f6TaDMYsibDb
guLexPQg1j8hYBShF7wmn1Ac/nziyu746vwdktmf6AFOmBxlp6vsold65JMuPvA5DUc/tWd/6EXv
/4ndTmDzhyWp+Uy+iAmDFtU14DwfkvViiqj5VwSPtk+wZXCIP7c1OD2lzcjJQIEHHYz0MV3PrHNB
8xwJZLCeoikLTcRfKEEdCuYa7eT6y9/zmQZuzVMr6krUogvXHzsZugqgrNsONLzaF91Qkgqhj66O
JAwyh8wlPMf1I703D4Kp1kYC483InUbFw6mNj1uRVmUpMS7YZbV3nNEnWQnfJajZVXwtQV6O/qAn
ZMIpo/ArColoXocBuQUajgtsXrmk8FTcFQtRzJQ57tuLYrOaTE9ge/VxqVcxtLrbIYVYYbe/TIO2
hJq7cU3CfiR5DhPBxBPamYdhU2v98yAi8cfvIgtKI+B5RQ2JKKU/jSU+svoNjgUtqs/evJTSsM2B
pRW2G/B9eb5K5sXay7mXWKsOShnpO8+HEDx5qydVwyejUs98lwbV7z9dC4MwexTMQIqAstWFho+K
OTWppuiqKSMYXUTnCmjI8O/YHek8pV01EfciOQ2ePhGYEtcp7o8ZW9mRkQYBdY0aAnhBDkIg2Vez
SFRzeyxIa4VE74FLJFJsBGIzVuVjjACYwYQH1Kl5u5UeyrEVEVyQXW4bGCgiIX5GPcTXe8JBR1+g
FIuMzoj7ytZK1HXNppKLu8BrKptieydZPfv/RcQ4/fBo6VhEtYBZ0KtW9ZPlFotSuEluQewgNFHF
7axGuLRtr8yDp/GVEuZ0G0521WUoCqwzaRps/YoXgJ75zLAMUIRgjX0vZSkOtPgY0i4VXdkFUgKP
tfUd0HjS4ldMkGdTCeXGiaP8Pnbx+bVb2xm8xZJLDl4+1TP7yXIsJyeZWGPhuYuEsysshmOoIxjk
ynycKfec6VZi3vym3U6O27eLyhpexEEq6S8rEL3nT3GhavIya3UzIs/Qee7RLVYx790jbX/tjN7t
i2ia+3758g2O8+4kM1SsztSHWfQJblj4rk79ZOCUHQiQbcgq24mQYyD+ecMastT5yRgfgF5bL/ax
UvtPTjovh3mJZ+i2tRClRX4pWpPISuicgl7SDqKVrBKNzzIxZPf2vhoc+1qdCse8cAxHIRLaJr9k
Zzrmboi51XWslsR1aVDQJaTsdUHTyv7nIy20bI6wB2xyC7q/+1fEZuzipyV+U2mcxMeakkO87hta
A1swH4AQxsqGFK2eHtz28ovGa+0QF3qqMBvZMBVw0c1bx+8FjB0HSn0gE2I2PAx0EKhBJpVdIxaL
WPUizt0tuMHh8HNX14ILohFfkvvICi8xdRLK34aFAHujhTNxLUlp2PHO90/TrnkAYj+3ilPTempN
cvVrEg7Qj55nTz/kuuYtq0g07ERsm5MGTMdBLJLfS+EziF9LSDmixt06burfwvwAjPdaTWFtAhSa
3PGrvGD2nizem2opslXj3cDaf3sCkQhDUrs0LQKoauZHQ20Lk06c8JiCPK218FmBLmnINlFcIWS7
GDCzKE0+8R9q0osv8p2qfi184e1SzRFehbkF3U41RtjN3F3beTywoYI8caaW7vaDljLTik/RHbf/
6d6Ja5YbUdRUdcdUDjnCTTvnElEoeCtzhzu8OUi66WlueisVHRUMV14jGjIANtSn2+lysrY2Gpfz
t2dfOezHvI1qW6T9F0XHa0bnDZVd94PKNVWeImIb9SlVKugvfNS4fuf6Ie/GKctzMUqkYxrUueQO
OSeoKx2ESSDn36N06dxyPJ56WSJbuaL76UtQnVOyREIcFeGADNXIwDyJ5ouK/YRZ4uroU/XBvPUP
F5Pe74a0zyF/neXTv9PhUGxfY/jBjav1PAOHKo8UnOJpyJQdpLBRR2bpt83QOYXjsSTPAJe2jTma
ASTtcbbH5l5vLJbMcWTCxYFgz4XDcKYTrWHVrb5o+nI5zxIXjOqeAFPMSs80kSPGA6C1VFEEGEUE
9OQLQdKa32pwkJ5Yvmnh0CV/YFWOFeGIzr6m5Fs3aX4rgQnrVG3tL+vkZ1v1fAqpnGO3qGwm3L6J
FHI53fV7078WpFs2nMr8lQ4HTnpvvTme1cchNC4Uc1GClW7xCYZlkUffIA+JNp9+gEjahD4Myidp
1/JhpnUooJDuFjUBuMIHvqn9SzKyNlDirhbbeoQaNj925gVnGZaDXZ1Agsnn7TpJQoT+Rz1Hz57s
sUQWQx2pnGwxnE4uqci+IDtqp9icYp2l2VL1q2hGM44TMq7UK0nc7Tn6zRDWth5oMw+zWDoFwHej
YPGrshaThLQU6t5TCNDxqCIEvrmFJjP+i5KWgYjVshezExt3+f4X5ZUdTP+/AY9qeKS8dBjc8XCG
vw/85tOOOAKogCsm0L7EeJsEzS8GkEA1bg/OgLhpjIibBcxSEQQxkUbGnJHONdizVq07rDIW6vJ0
KRgcN1bT7D6pr6fqtxKoCPZ/gtrDBxZSO8uoueQSzJ5aG74WolfE0EBfeiEBykwkw7SidSPTj4xM
S5cteaQrn4bLNnhXJ0UsexdJiPMm/sulG+hUJnyPv1eMdVTn0lAUXWdokvH/WQk/zx4WfKPf/93Z
4ONQF9H+K0R4hA8Et6+sK/zRoOZ4aWb2WUSPeiTgbr77Qn17GFedogHDySzPPnJOVUQIimSwf2Go
zQfazAQr4kt7Kr8N+b7HqOGyFUzADxyv+4jzUB3NmPdueIt7GEHUTOn2sEOZCtb6MdwyHJYqNdJf
XO5CdJ/wJ9S44ph8EZ7geXjD2ew44ZofnizStaDQYWhjy6A3IzKl0krm2ZCdChMJu7466xbMzGcL
O84xq9aWM+nS77XSq32f8Wgt5OgtiDuD77voSozRyY5ogZcgG41F4IL2yp8a5k9KqWRJB+qt5cWX
ZWK/UWz7oaYCln23kNN2EgUgSg7RrxUGM1vExYj2NU3g2fmUD6H12d77klnk9VzCBD6+WB1GpkGO
Li80iRyBXLUnqgvTzXHmlF5nstNdjfUj4cPlbeDlZzpg8tukp5gJhj9nIhS1cbefkXkQKBETaEY1
P88JvxzzDIbvlfEO8VHu3HhdtXjpFY7OO+XwLx1SqnGtuXk/ub+ITJlUXvUHPwDJ4iFzMbWMg0Xx
7YBBfuyOksDQ+N/vYcd6H4UPK4cy68m86M747GxtBlpNWVADboDKWx3wvkpFu1O66dOf1zUFdRHH
ezmIjfI2BZPDh79Udd+UkSZpkR4pvBIgoYob0awyWSUqpDt6S0FwJqUcGY4fhrdJaf1SkqR0R/HM
VW93PB2VN4y46zAz9dXIsKhRFWPMoHM9FPAMSBbT0AxjAloDwr0yaWsEVjidb67JOg8aDmZdSSOW
PD9CR33GsFZYpDZCQeXs86W08/X3yWdLQJF5+11T6ibnn838fEpQzNd0/Ji3ySCkNKo7jdfoey5P
bysKrJUpQEAQTLH7B5o6ykeraAtRVFB978E7B4McAh15bju2MurgmGxBsF6rAOsiqFiQe4mq8fh1
ipS6IU2ndQEvNev2Ol9emwOcPjBGRDZP05DubhNS/GIRi43P5kYiuMhUf1QS/hVAQ/ENVedhmF2i
BVSH7rndIoZQiGZoBbQOPFHupfsSLxqOeBTDEr64qbfp5TyyQZrMSOIyCWtrQCdqAJ/aaxplBPGz
3REnQAy8tIQBqHR+pL4KCerTxdBQomjiJW7CAlGV3IMBGE1s2cuI1wcSMruxOPsCb4MTJ12gfjGM
xxmY1HCZKs5l4VfV/5Pl5hRhdP/WgFoGEzl5TI9XBtuUkrxaZN9/VA8LQFLGnxFvZRbMtMaLig0n
82PCaM+IeRQWSFqb/94k5o/2TOZqG3LUAlHrsSnGdSdHSSxVyPt6UEVrBOS9h4hxvHVhc+zjM1l6
+R9ovh67HtYr3IudYeE5XjrDz+fcwHZJ3Tb+dS8O+MntjrX40Aq012Has14GRHu5v5BPpGnc+rBP
vGjii3p8EdelcdWYzRXwpy0GZhRVJG3quRqnID/8Qsuwnp8Pw4gc/98FW17yfGMlh4b3jylR79nd
L5iVPBfccwbibcg+Cu6HB9ZEtXk4Acs7iNLa7ua9vYUDDlrjRCt4q8uxIDjbyTO1nnwBk6Mm20Ln
9sjIxLOYi1P9WYIuLPyqfcSiiwkhv4WAWKrtwAkKor2H3kpfww/V+P4fsrIrGSm5HU43LUIMGLpx
D1TaNfSYbjbLaNNXqQwn4P8GJM+SxJuYsi+vzAlyQm9wZKjFsZvulUc5paAM60bkiAnKk2DhKRpk
A/oJqBsJy/3dYPfFBXSi/zWi38r6QolM4JV0zWRvf2v2PqEZ9fpd+wUVuycwthzemufMQ2eLCCAZ
1qv3qebMZt+KFih4G1P8j38gkT7nKK2p2IcQb6NOSAArpLkEClqA+/33naKpjEDlWkDSYJ/6s7aJ
WmliyVDpjbdYgGyk7H7jLACPru3v+pClaL8hTlamWZ7bjYY9kBAAMwwdYTMahbqMqtWkTUYZlznq
njq3hGzFAgUm3FljVVtmg6ksMzBNg/4WffRNWnwoI+NsDDGLabJrIbfyZVweXEcQRYNBuFluI3K6
PgZsfHebLonbFseI74fh0cmFddBbGJbxAMWe6LNeFqcGKho2a3Kp/JzPK3SeCMCb7ehXV7v/sgpj
9I8krT/09ntdfsKJ8QfC0iD+3G+J94qrQtHG+kfbl9FGwkEJgLSadkrMKw1X6DMQwVqf76dtjOR8
e7DjqGUUoq5Xsc7DiH0bjtaTCtd9RJHlDjpNfO2Iq6aHxMhtl1+HxoSObdX/sE+xYuA1wf3RtLKx
aqdSkY6FvcvJJmeQdHZrqeBQ+Ba7FbWtCL7EKhqrdHGU1YfSgFqzY3pCZIBRXzl/F12xtSR8qyHt
m2+GyvwsuW+oEMNYSjsiPEg4wpssCcE4FtRjjcwQacn87zR3mqGY5HOBGOPmX1qNPS67IPeqnlJw
05n8k50tuJVqo1vY+gJ1pLCxCHEYjpIEWtn+vIWsyINQx4i0tn3Ig0l//ZumOyybgDZAOBta9e/3
G/KGgkyUmN+denmJePEZqAVStI+DEPb9mFV6/WH9pRM2ZfOs3rYNBSBCV9FwbCqiLBa7dfc7R2FM
auY838aLtMbHRNVQ1rSCO/hXT0zUY/j6o/ejwwVSTyis0frxXnVhoi+VsIN4NuSkx5FmrC7km4WE
aIZejMT5jOnYbJnL2r3gP3naAmG8pYJfxkbc++jnG76Fh8RYn30gvJCRCpVbH4JHU1P4ojuFx/JZ
dyKtUTbRClYcYq2nFq9jxgedrwsriX/7TakOgndeGj90poVy3Q7gOdUJ8M7EFZCSbBFKhpKWyBVr
i6ERnZxw2DcUUF/yPCk15aiMXnzauZz6OqwThsAe1vyRU5fBfMMC2ofni8yUxVThq7PWhWyOp4I/
zpQYk2337drWASBDQjuBEyXgmsoEP4HwzsdHDgZJwtkfgTlazvDXV4JfPYiCiVhdmgnFA32BTbgm
s67/vxrW1cBZd6Mn38PTZGZB/nzNUqj1hGqT7iTo6IUWqYy5FeNNuaR/EM/Z3oMfjscm1j44wI89
RmocJzL535pk3SjcpXOUZqnFFXsfJRC2opMejG1/5MOtsOqLkOdwnDvsuGQ+WJRCBuO5oChp4fcf
1QXr9pMSyMNyHa/HnYPNzKQcFE/Ieu8sLusHXKTjqI26Ql6lTy0HDMReA+ReKd9uVNfjskyhZ0x1
Brrm8VDeqKJ+4NCr1K46hBKfDYWfrHyAOXwUs6ewKFn0ryEB36xuyXUiB1CPNUmjyy8kAByKE5TI
eUg9oJurCtJl0AnJQ8hfmcfd3VppvlMwRul6ZFqqxh2NjWsuMWlpeQFzRSCdYiDId5DpxJlks79Y
XM8fBSP0FIbWZIY6TNVqHpILVyX/7wl/UExRL5X9dfD49Rx1kQ83sH3BHycSm7dfy9qlasjsySS1
VmFYn2HBlMzPvA7UZADRYozf020bzPQ1dsJsD433oQY+qjtInBzEcmnyCPcusEbulIXBzU9Wu2Hq
AmopCZIE4Gbg6HVUacsDVm0qF1lZ1QwhlbtA02Gx1v1zy19hvnKf+QsLlf3Le2ITHB8XkJOPV8y4
ahrg5RBc66jId5pAbpT1N3o6bAJ2zMiy3dHloFv9jK6GmxoIlifwLpoEWW48yCFMIoedxuam/dP7
sPuB9aJlm4db6aDZ0HqnNzZyHuhAOtL5slodIjBXMiPSYsjJlwFQBOVRT6WqTP8VWekC9xNHzpKz
2NtucBNAd0PXPTLIUuULIZf/vmhzRC8KRlyAO65nA9ChXWPUiYP+9OMXIf/Yolj08lyCdvJyWtf2
epbN1ekMVPl4HXkfHW1qYInWB62lESFARjUPKfhuqIyfHNv4QRXYa0wicQAk0im1qzNR/ssdtpzv
AwmkMd0TbB/fQPd4Tpd1gWCje56vaaZNs5dNGHoSiUmz9iBRKQ982Viaw3+/erjJj26L6F82E/69
ePNg1dMfR8nq4U7kXIwSqLZvOsoWqVH4828dF0xHcMhSv8sUlizFKmaqu10KDlDQ5ByrJLR8D+xu
LuDz4yIVPhNcY6rZGvEiB9UZ2W6rmxuo6aWPpbtByFww534kaIH8I6NO0A6UOuGMIM5nIjFzn5jo
PZWZaPuYNdXtfumT4R6U8x8Beqap98mi6nD/TMOtO+geVGr+hZVzMV2RfQh3NnLfGNHiPglDPJgD
CXnnpFo7mkm8/VHvTTRdDRvuRKmdmCGbU68Ygzn7obnCVh+HcSbnZ6R0rcd9hWpa68/+FW0ID515
uQpOxRftsmuxTTmJjnJ05GdlLfNLdZ+Y/Ut2NwJaCI1VNsmbM9ytcqTpXhO1PPBdNRh6yqkhRoGW
70tPBwvw3Gld9f4P8Pxq0WW0/fP6xh3D1XCjZvfo3WabClIQzoI9oE6gyhvodGfvWFbLbPK5iu3C
3YT24jSyA8bMoNsyjEqkzntyOv81SmQ5iF0BTIkD9RHwoYCUWzPc8TcmLypDkBUiYBAdEZdpqPWB
Jn2CawEtRBaF91BDjd08EEsPr0M3M9AnyPzY27x50xLrpCs6RwBfDICS/rFrniOB46TMIC+P8Or2
9hPIzgwvYagMeaXxTUU43Dayy4y3ogBR+MGLW4e5xK55Zp1A/RSKNCs6Q4zVIKBv41tSH5r8fgeA
8d6vH0kY1k+gzEv/2tV610DxfjMtUj+amkpXQS2701nRAGxIl5b3ZnAfz1x9eJw+fWsnz1kkRgoA
2T4FKAhRLz4k8KA0gBFLzSi7wnpt8sbH16yItlAndz6UUtupgPqZoBv5mCEpk/XXzlj7iKE79cIs
qZtxmB2/8U0e1vknIt6THhBqApejYZdyadtaXvU/qwoe8L3yC7dpvre70CTvj2RzG7xmcKcj06wG
RBBo6EMU3bJM7ETAB9/C/cHk2b3fpOkKcbvmh2YuUUkQfFwUjlLz4qSpavxNes58gTcKHDxlihOL
CZQrv2XcrWZ53xbpOP7XEX3B4YoSrPKPxMfOM3z+cAfBAT4LcgDvQOLOD3SwSHAGyGQvBWXwcTZz
fdg2VfpJYzsaQJD4YQ6xNgXAqHdZezpGVHp8Ptgxm6QkXufQVthGrmSctszoivHjTPWErSNkI+TJ
RxFumd8h09hIbxX+XqFYLBH9Ft5gElgJDDAyKJAP+hPSdJeQbWq8dxXBvBL2sePyiSS54KR23F/M
yrcg4Gs/HfJMNnXzytrHITeXeMhOx2x1O+VKwpvY2KrNMYcZvEDINLNhbl/7/91Tc3+1fngkJH4u
q+67Nw6HOPr0yS3zIlwaUa06VlrUlLgcX+GVUL5z50Ykdt4x/+BDO01dbJZBPxVTpQHevNQJQVql
wEmDKROXav51rxAZxvqSGnb6edBnPp5MShWLV1meqE69KgSEYpYrMEtL/xdbu2ipSBnoDUg1Ng7/
VOo2cYTCWI3XWu+rvU9RpB6p6EsfWzLcZwo8/2xGt1yTpcoWvY6HEWmmdHiHeBYsm8IeGRNwmfVq
QSbxu3Qz/YG8PrUtQaZlwE8tjKnFja8dJNlPATJ0gGn9tahRzZa0wh0Tq2ca2UnOzf/scb2lL1TQ
5VLDxQfVT4CDIQsevnhHiBvwO9gALqtuZNthZyvzITWawE62icP7h9D5nyxO1CYW7PQdp5pCtBMc
x5r4FBkbVIYC3kQCXzbQiCq9GnfYxAdUrfoKnbAs4HpQRTm4gNk0a7d302laJ7iHA2cROBbs6yu6
WdUE9jTrkojqghktFfS8eNogCTIFdLzc0oWu6vsg85GKJXgQJ5kol/i1v68dU9iTsTPZJX2HEvh1
IZs6L0cjNRz5bbII2jZ5IVgg6+u4j+gWAAlS0C99UO6X2hFTtaHGXrVKg/kZJ8exdLOPC40AeE+O
5Vxo8OfZr71XOL48ipiBuNwsJ0lOp3Gpagi9jkM7pqyZhyOtb5ExOdgt+tJz/i/id5Qzh0Mxh5gu
Usjzlc09M8xNNwMlMozRAW7TqDC1U4MofoiVmzMYUuLsd7swdt8ws39NGxXKXQ1wYjRgKrxQD47o
8I9Wt/ttKZRSLxheXMPV0MsqZIwgTRD7sIYdZJLTaVt+K0igq7wElV0YAhG79PI8BaUj1G3LOIAe
3zqEsrrUklGI+8iplyR+CRBKKsMmnwMghvaJl1Z4BZV7PF4UBV3VOEJxCTafeoWu9sm37zeqBPCg
6UV9AuUQamkbp1HLnZM6OVQLX1CimsF3nZP3PvYZRbFzCcGCwoRg4fexFRQ/N0IXU73zZtpQuYKZ
j4wfqxr3+rud63xLNZZe4CnqXCwUWHngthfyeg0olgLdDC803RDTzfPo5a3evebxMP9/aaJi5+mq
J+xdEJdjRmQRK+R3345tGohrg7wtaBJNjHgdldAkLsSJr7wAq6nKbhtgu4z0tM0QRGDBuiKcBm/o
1AJydngAAEjIXCCczvKygb2l02QneVL8sXiGJLxBp4431WVL0bMdhrFrCwbktSg2UtPN49jsmORv
tYn3os4Mbxx5gWbRtqTjt2PnOt4dTi/rkxD/26MJPaqLm9fQvXd3vl4oc1KXBCk3OxRzbSNgZBNz
4U74V/gwfGKILgKvoJ5x9bD2WkaMMSyIZGawXbsYrT5ZQ3ZqEDb6s9QjbRZORgWAD4O2VH/2mDN6
3a8h2KRupaPTqtcQngzQQGzNmqyIBOFTok81NFoJhPIZk2DSrgtMCREmUqqjxi5zEr9m9v5NdY5o
VUJ3iyLXbjBRjK9nYpevENFadf6s3VgdZlGmk2ZwchUilpubuSroMOU65Nm61tRDRK3lajnFhZKz
SkWwnWLyrX6tEFmocyOv43R1Mvi4F5YVHy5iWsS+7v7NpMldQNIcoUbwSJtCRojJPAuVHBKn61Oy
12N6EzBUzuAIrzAWxMqFQOLCzWHcs6Q/uWbgLtK5070qya70XHQGDzdU0CNdezoB66QEe5BEbysu
R+qku2Eo8uWaqTVnNL6ycnWUfuhfjJwadDhcO3hxrxEFzLVfjgRrYyjJY2r/4POcFKrwC64mUsIo
azpt8VcP/X6rlORy/sAiQXMoaC306VHWo4bRY7Nn3I/JTt6S5rDxUba1toN9M7yecDJfgUHwiKGH
ODkzuOF1F/od57dXk35wE4Ji4oSAiin8YH8CSn/hBIS9IhSVOe7hhXGjY998gG0+8DNIl344ebth
KEFVfC7irOuOGYu1CE63FGqyyKYGtFGr1pI2FixTIp3jA5bDzn6NbX42/Vpf6Cf8TCG2/9HE19vW
JTdF9GiyuxGR1HShkWMFgkFiuGE4kiaMPTx5v6vA/Yd9yGvuOURdAHQy7eAV+3dscDaXfFCX4aPh
in75UnD6Wgs80Tivk3l54VM6Kwky/Drg7K7fznBMyazwZ2BAiXiaPgiVLgwrcsofgZ8v3yMEQEdU
XdmaoHoL0afR06Hqgwpgp9aMtlW0fnESzq8nQ0FyqGYbJNSjCDe4W2SSO+VRNd+1jITJL3OWUoFl
QrIVRlUnv1pvWGmu1oMq67qlpixVrE0WnTaoEeN6MMibGZa4Gh9nmTUbSRntJvCjBMUeFJIqF55A
DsCYGT/01YQo15zJjizxuFY/2o86tHroB19dWCwmiEPuAdEz5enDyQPboWOF9782bejP6IYL3C0g
lC9ZPfHXkkZsOIestudF1DtuyFReeVcBF3IWEoQJV4QXtphFVjLl6+m5dA6tLGK8xQjJczESnPKW
6WgK1Sg7LbflD2NlCre+6bagK7VP//qQn+723rikW2noqrqqtRlMHGSNtVZESiy9zuF41k4aQGUV
uFOoSv15iBmmrnrvDKyMG3d4x9ymo4+T17x6m21QS1z8jEu2/o9pLeehBXY+G8Jtbx09ACipIpH+
mo6G7z5Jam3sbmyImvrXirdc7ynyuRv0+eXapa/aO/CQML89BBxJ/k+ZvoQ12Xa4yTW5aN6RpNhN
6F5H1QKoQ8isMfR2Zi6sqXHAcUMTbKy1Zz3IRz1iH6feJD4xZVtUl8RFqUWAmRplqo/hMuURQw6e
CHKK/begBvoLSCj7f8drl3/VjjyXs+A2k4s07X+qduhKHBfkhBKQGYuOJ5zq39BNg2rc3pm9Wkg9
j62QPjDm7z3+w+ypsWhuAIbI13UjPOoIzamCfCn8zwGeCxmiB0ZCPdbYrE+mgl5Fs0neNCX3whV0
vT9rRw56n5FYMy7F6iZgcJM3K4v1cOQkacuZM2k5P7Z5q68fjfcJrVuxIVJkDNc1dF9aPJKow/64
uX/jqk2cN3ePmyzXRB6QR/kWztO7UIM5HBHyrop/d2CK2/7Is5MimDfw5uM+FWim56nM1z0l1wK/
PseGn8Xparou7vIXK8UFTxSTRFam156CEoO9Rd7p+GHoxYEIrRO/LTorCIxgPlMn+voBD5CKtzX/
UohU0cuYPloUljcJjZInxQDWFWXSy1UknWEdODrCpb+yM04KxKLj6NQDsk/Tnj9LUWuJ0mvLlxjN
ThIun54PfhTW4kozsc3ZHoGe3z7FCW0mezg4eL67WVI2hhfE+CuY288WXbvhOU970W7tQ1yldpK2
COnalI0ESZ5j07P5EiBm5SU6LpEywA7lW+VQu5lbYo2R0WWSIV2HrXB1mGNMBq4jGyf5C9WB6dL0
EgUWy/oXh074NBxqo+dgs902OMtuwE9+fDgAmfRosCbRym+cFnZBsZIfbkXSrs40gQx13p6VZJMK
OePmXIMgq3F456PcIjSyA5e8Q6Cm4B8Iu+DNt+DQA9tV75K1v5LglJTV40ErBznvVQTNOQzHqAuR
gJUvyxPKgMrsPQ4Y+XXs3SzAkhhO7ucI/gRmo6VAcSBrxkCUk7kXfFKwB+P/FwqmAo3oGBRu3gtn
Ux87cw2Gcls1+JPCk9Q9iNxwZu30J2KnhdDmvd6c26nFFhDN/cL5j/YWJ2qHLAO/1Ku3L/OMxuUL
OaA2KEAiXFuN7C5tfVu0zIXcRSssbeQgeGDmxqygFrU2kuHLTAvRPmLokZ2o0suQACU1vAz4fJLt
LP2eN4LVWZTSJT/gZpV/5319yT+ispDx9p9+iBRLJ5QTi7tJctKXgLUwg4J/F3PW5in5xz1afFWI
eRKDaYDbdMKxAdv9zCi+v/fgAPmj1N/ACNo1nUkA7ycIXnBkC0X0A+IWJv0x0EnbBXe2mku2pQI0
sYA/2sZ3JE7dlOghYnq+GQ/yfoD8jskyEpGIqblJxgDew7hUlv2RbC0DcYGfiMxEBcDG8IwC9yQ1
005OdXAeTNSM6BuvrfNvXtJO9bcMwTc788XwbSqX++MUcgPCPtddCOzLqgauSoC7hpiXnZ6aVX02
fYtM0LZq9c5IKxGwchK3BgOzmEMmxeqyjky8jN5JwVGdm7VByNFc7yMVpdiTmguomEARDvg5B9M+
8xc/zbhTyrdBoTFB4hISzEGv5Xn16Inj8O5qAsxyN9yimgCfvtFl0SUYQ2RS9UGdmhGnrzgDCWea
ggWZ8bJNZGJp0lGW668OHBvGOxRqwv2dP3VKGtWaj9G3yRX3svFzeEAiwcnfmuVWrWdBtSzTcybw
a99rLUu1rIO5jyS/DvwGwmhc7jNsLoTTioZWuRlteAtW4YV9aotTSgC3nunIlKWnJ6PwsihvASO2
dRKVcggMZWwTheBdtBNpLBI4IuQzRmIzgvo5w+tHMTcQ5u7d8evBevEOV/rafzCkGKu1zcLcALOZ
TIrXAkYT3tMkS9tHVVBRDfJavuTL976lVfvybXcWfWYpacQkq+l0pjUyqHdkS86qYRuJfRgSIyxi
rpl5rmCGuukufNNxwFWVH/r+aruCeoM0ZZXMXenlV/4SRjvgOlmb0nEn3QBzI51VwWNwset6YlLe
GRkooiIC+QclASqH5LNpzWnYgAoBHygVZ9yopgoDQoH4bYJq++7NuCESyei5Pk/K8RZWevlrWwnm
2RxP/LZcONs1ua9QOxdZr6f3ygLGWMAiciRh1TGyHBPcxysICxmqev1AtRNNGq1TL91tduJeBqcr
a0PDGBy5u3pQVJRfXgpvzPv5l05c7CNODOIi5210M3D9dUKrvlWE5/CK/DjXh5pnFClbe8212TLH
7/W4MRNXNDs3eqxGxrWNhspBpJqBmjGac1Bk3hezbPaxdcHrH040PIe99PXwsV5Ca9OKpANrw13u
D9nosyV0vEn+sNqmrb6JIzo1HF7SMhODAALh01Ccgn8IvqU/VRCajp3g19WsoSuLal3LYMX+e/vH
iR7CKjMggjKuHq62kcBLnF408dxE3HVzz0DY2vCnFZk1r93wBoWWfcX5Y5L1H0qhsPwN04CUUseO
uCX4HtGAJWzozj6hDdg+7zDux+H3THSTd3l5x+9ZQ9g3Q2mkYL888bENrTYFtQx6APw/uOWOetnU
1SFu999d9GDIG+ibFpFjLdB5/tAH95hAq/czkeHnrT0QVSL+JvcGomu9fb/r3Ei8J7BC3AfDQAXF
Lb7co2Mn0+2YQZ0jVO8ha1v2+PM+6tEqTKe5HJ+A6wCyjeE1H9hYKf5cTJIj4shunVYKaFXvsCZE
F+ZvNbyT2dSCu9mMUFn9dm9geBAu1irhNrLIBibFj8qslNTv8x+UD1QbZmwMHAaWIWU8aPMirCH8
MOpK/4DIxQ0I/pxsZBZqVOaUlknjQ0CUq81pAcCccxDb0CQsmzSqA4b+E/b0PP5BC2p0XxfGWVbG
N77D7TtiLfVIluYmVT0wib9JOa8SPrmnJ0FDchzcCFJPY1YABRdJBmuGyNsU0yURCljeh4HidGBf
lKrEAu1PSrN2vpwXHYcCkMJCHf362rnc0nIp4NUFXI//NlUWF4bW2cbMkZWFjQckUEnh5B2sBbbb
4yAbQkXqVRZVCLLdAPLLnnAeFfYAYIAPx9xNPZE6iB3QPr+xUaNH+reygO6Khli0lO9O4Kfatg0z
tvs3+w2ebhTKuVyW3MpvmHl8JplZFeHqV3i3eDFDqbifJQ6a9CFndVnZ8YARwc1QNpsDqVTjzdzo
iTuRo8WkgshIkAn5yiNgsRMsuZH64h9+C1WAaxAHv20uJPZt/fEnMfCTPqTvF5OyLg1nAH3F7iM+
/nY6VQqA99JXhjXrcdqEWdcSLa2LhdaszVopxTlGrv1r4R8XSPXFEQlVekCO/HlQpTmz4gHd4/a4
KLHFJsChsoIa0pHmZ9yEpVkQEZzqmlrzt52jsjsB28BjzdzIcar8Ot6xdYhyF2/2Q+2YUtb5bJtp
KgHHBWeBKSMdWXs8ri998iaxQUIAMc0BHkv2vPegXA+mXpC3aNzZrfFvLIiIGjdvckIOu9MDRs54
yuYadmBOmZm+Rvhnf1hlIKIdyrvTnWk8wPE8NvkB/NcvcwsBT4m7KIOVC3nsVyJvE8nYyb0DmDKo
MZpQj7kQqFxW3/BTPwMB2JdI5xObsMo0hDX3DnBDl4JJ2dO66j+L5bGzyBSk/R34+4ecypxJPB1H
ILz/gYINfc59u5iIIbrVVUgckoilHxZhTAqAsmR73CuydfYvs83xVL8hC4Dz6Ztqea0cxenzLiXl
KbOLRTwo90MxrmQk67ebIr2X4dsxHpPNnG6XC94E5g9hwdwoVpACKIy6DLEnbYAnbwUL1V2sUoNV
3FqT90dsxa+Bex+K7WTsO0Ky6cHfl8eQv7rdnEI42L1qa3tLnxyoUfa8EJnItxFQ2MlxnO0e8Fu4
Oge7953OQZ3aNsTXyBavZ2vMfstr+MllLMQ1jvBaAsZFcqSEtILQ73oLLrlXb12eGAIxu61qzDYv
eWIycfYjfzcHYCOH1GUeA6mta10tEPx+DvKXcwe4eiI24ZqnKOhKEMFRnZz5Eia4TxGzyScE67Rd
0dXlccHVx5XDMKZyFnSx1OVBhbMGJ4QI8w3lRJzuX/PKL6KvcNSdnsBMGdz8hJIcWoUCGpALW4gZ
Xz2/NzuxmVaDkMrTVzCi44Zn1PWLVSYf5i7y2vSZAsV4DEvC2fKgrBD3mVxJnAgqFk29VBXsKvdZ
UXFy5Fw9Ye/zriC7Iroo6pWEYmrK/BQ3JY3W7yRfpuHy0Is84XSrHrsF/usgOvVUdw3SNm40N0Z5
dn0w8fmfmV3dwJENUk0xLksJUvclPzXNdL2oSzrkBDsvodpGlM2VLVEHtnAHqVyzghqoqpdrfPP+
KeonET0a+XognFzyUb0ED90xnjzAQoN+hR0BXAFKrtm+Ti085cGp4demeFk8Ookkm22ZZ9u/I+Se
9W/44A+ISlQwQknUoOQx/H8WX2zHT4ifaeEo+ly3wngJzxUfJC9uqe9kiFksWLzhalwYFLj36T8S
lr9PBXI+7iuk+oH4tdf/vdbxuHXWovm0HWqrP0TK5zpHhpNnRPO2H2L28r4JG02iEFOjyut+/JV8
fA6TzPpQ80CShoK5qHyBE0xkbDg5bbZeAK9F3QL7kHI6hQ65IowLbM3Vp10TKSDp0/l9DJ+whiVE
OLi2LSTJWLD4zGCcPVLRSKMIPa83Iva7NTjwBBnVpAEvkO3OeKDwqdciu1xbZEcd0vuyUiYDqo+V
QHvabvJo6Npc4nSGgZsIQrgXF9kfRDVWP0rGlB4lAZG3wbtp56JsS5Z48x2UCaI5vLtIwI9nDL7V
qYS9JTT6wGZEKBZKaHb2VeetTL4ouIogwGARHwAjvjd6MT6CukZxgHOCU/tMyyYJ6HI/5pTw9Q9M
Xqb1biZvIxiCeLKO7Qp7RUQd+yP/oBAZ3OmedZk6q92aDqZpLXBAcZJSlq/MmtnK5Rbob4b3cwLM
3838rLZi6JPficbuZ2OKHSmdztXaai95YLY/CIcCIWNrXnOb6WRhf8kKS7waVuuJ5mfdT18WJe0l
kZ1Y1GLayTycLjxTllBcYhszaaEYrbx7UvoDq0j3byhJEszQTwZo+vX07dGvY8+c/Att/ZPNBY5e
HNInegRvNjR7Nv7iwOqHZ3ofOBjkNno6TRjxN7eUNIe/Aei4Jmh7vmMpwVPCHas0wHgHDA9JRHno
wyRMu2flnPkn6dmLNwcepmMGWR+avncwlTymVMpeSByEVuFmhY2coASoQpE8y+PN1QorKIC+y9oQ
RMGxc9TsGnxcP2vhWVcY9/9KY3DRgQHz9xfN8CD3h+OACoR/hazMR3WESYnUbvGu/GBrlAHC7Y3m
V/2/z/mxKwYJHRPT/aWePcmthNMJyHwFs54EpIXfaJAIe9ln/bRwI21P+eKNWp2qg777neaJQPX1
j9oq/8iyamd3lmcdpMaIGHDSxZreOAOSQEvsW3gWvORpq8HeUXG+VcRxWq3KoKqzSvYVXMADwrSO
+Z1JVNdiT9Gd/PoByiDc8UG2GSb+pZwB+c4bmfhw3FSL5UYp/DsZFp6Z4xs60rDSoc/cItlUo1zg
6OyjT9BZfGNb6B9cfC7MABYjHsY9B8alqDnI3C19j4wuUUjvT+65JsnxRrroQgX4HZ8xLnzP5m9a
avZYLupbMabdj/f3bfFllqtjl5OHg26W/0nxOb97bkioJv76OGiJjhttjznU2IQ0lm92C2dnptgC
ZhWo3EqzBd5tOmNW+OTa6DLU5Vp4BMB13rjfMZT2I+7OOFc7nTq+XaUt31BXhqoN6xuY9UPXOVoQ
XOmfJBpHVoelg4q9xjAdUlcsrNVP320PASYRWWzoQb42ccYEcBKlZHckqpVyQnJsZXzIljMyZdHe
zKhF8vLHe0arGteHK86OR5Vw7qelK/CrMi0h74bYM3yv1MYaZUC0gqgwwJTP1GOCAJEeZW5UKCkK
uug7DMGMw1BwoSHMFdgR82GqUl4/w50Ih0uZ7vGC+lUOpJAn1hA4ua1PXAK4gk75mRyACu8FzaRJ
5+vdytRjFvfMaRRUO0Q51nZoVOmV6SP8SCEXeoW/PgNIkzNzZqWr2d9eKC2g/EVvHZ6OOAzKg1kk
4n5H1MH9fdEkysmxNCsZBzz281X47lvtNpUnCab3rjf60gRqAllDuVO6AEMIjiabY0rUtLeq5McX
qCQX37kWzU6A0AzFnLNXEPgQleJ4vKq24zCLL5DKUo+ZiB9Y9u8rjKqUy0EtRlJFPgJCmoTMFa9f
vLPTzrenQjsjG+As5JRW45EmBBdrDxHzrpANulNa/zmzwkk76LPsYp/iK3XIikgY+CGRZdFMhWNk
Heidzos0iWbNx2ASAX2l4DXJ+d1Siris6jhcG5e8MztcVW5WADrptudiXHhsCUaexHFeRRqMqPoT
yD3pkJ6if2D9VSq/3rx8XEjNVcdokwuk7Y/wEnw9rXrxjfcMZyxMw2WBU4PxPLm2qqaUJ5Ngm2nP
2IVGJ51SvqaDhgx5zx/Ojvpx361kkBlMEBxdSQrM/luGk+Kx4GbT7gXX2+hd3TbZfx/HLNW/M5b1
ypxOihZz/6XzXVuCF2RUep9hsrX2iBV2mDTaoAdiTR/rIA2LYJf79RfjTiHLX9CBJ+eq7m6EA7HH
0xXFcGQXpetG4m9Oi0csefL5P5XxH6SFTGTGwNjQNycc5iGEbfQ1Yp2VXX9a13cWr4fV9xbd7E7C
4rC4Y+v407yBsqaceTHGGLHrYmeuTjIyDwpW37TPgkFAhicUOWSUH+KlRfvYLSqWfRHgop85MbDp
/rJDwRvertX3gb6j03hh/Glp+4R3kD4gkdd5w0znhWjeq8CQvMlGzPJU/RJtyt8JPu+V0vIjh91Z
QWE+g8r5mDz1IO6iMNipMr4xLMWrHiEdJuYjCyPNm2N8MSVsYXz/kLpuWRfbdJq1ZeXV/zAeFTT4
8KBLtW8PimOXN86DfS0w16dv0acLU4XJGN2SnTc1OdUdj4vdevZ5Ok8clKK8AmyqphSPHGvYD429
qJdfU7sAO0QpLhx5HY/FfeoVjMcNftfnhrPpL+i1FAVYO74/pAUmCAmQMeFzeVVdsk7OtPo4AK3l
GOogRiJiZW9FdT6lLYbT/OWN+w3VS/TJsc293cJOH1F0hgsLqx6E3GmWfBINlfhfklhevsfOXAKk
6ptX8cWAJ2EMiXfzGknjsrIEzlaOYIDRqXUxpimBad75Vz4tBa00QiMs7/S7zKpaKg0Gsk4bGh0L
/fP6Jyq6Ccy5wNMI/vPPW29lMjyyMgyIWb/CGTY24hq8fPk13ut6zwzu9obHSXmyHudzFNMUlvkO
/KSd7/xPMu/3/NFW2gYtQDWlDPDAvCpkDGDGSyt56iec24TA4KO3gPFN14Uo75hV1l+YyfoU8rQg
A4qC9oWU9sijq2GcTt+zQKbbwr5p16OxOj3T66Ii7cxXrmRUjLEKDYi2zKaMUNski648Cvl/XE4L
0kCtv6ZY/C3QvYWfSE08v34wuh6YyN88uESQRTbAR/ZX1Kj5aksMl/I1khBug+MMBr6/o5iQpiF/
1bUH6ihHEVYj/pKCl4HMYVfUDDEDhZJ8JB2qrKLdv20ky0mLZj02YsbN9n3Rm8X8hz3yMCIvhWBZ
hfUlEigIKzQonRMiGDmgmD0arEdzbXHeBvuMClgvvty/rv2wVXcgmoz7UQHOr1jKrqpTpO0SN4d6
dfsjgGMSTKxYNh4cvWQZjfJFnGE63/UCvb9f7ykFO61n6PKu9pC8LXh4WBzWwhcBduWWEKS+4Z94
VPOF/VkNyUqytqTlIZRfgEnadHptBc4zVeS+gRA6Csa58ctJZpScAlgt7p7KKfBsxuhcBUnCou9y
CajCWeFeChJnGVsgaHlFJB/D8nmygM/93q5xBuE3JzATHL7nagZMJFIC/XXQIyZWPEF58uR9JcRX
j4aIXHMjAclmBa9tsnCw3RKnsqHPqrmUj9j6Rrdjlz6nWV7TvfwVUDIzgbPSMmWAz9415mkY68lA
zJS1rEfHWLHLVBaH/N2MXGG1eltMpRe6oi19uNDJQ4ZkOZtWR7F00dYxiLDUZcv/D3CHQdi4M2xh
Eyl1OA50JZYaiyw/8cPVm3CFHPdrGUE4ho+eIwjEJLdbyF/kfs3mfWfN2M5Rtle7tCHnXxlwbf68
jF+KEKa0snCqNmcvlS/Iwwl34Ff05hrA17iSpXEVVQ0aRNbh2eM+X2GndDPNA/jo9dHEP0tey4E5
hQrqcCIM9C1bTX1NwjZJQOFOzopCD+1lVCagAOf0o/fz1du8ymhlHbHR6GSqe/b2NMeShrCr+a9b
xApac/G3ZQyS3MkFNCaJ82vMDDRduaXwQEPZ/+nsSXfp6K31o1zFRJVnmE4rmSp3AQYBwtxEyBo6
2ycEEBMPakQkg+/WZQR7tknoJ8SK3WLfqTCI2vwDQ/tAaLPC0+7l5BilL3+f9ndODPRzgxKCwO2p
CTe0qvp8j7+fUQGlm+dwxdKCPS/83tCYlndANEEKWxvlssCORvvsI4UkAzYHGThUbLgcBTW9ZqOM
B3JmBMvYEmUlRSNosqhFMiQ8QDygPZD0+Z49dznHjmepaYGkfxGRf9Hk7rJjwEZBlkZwCGDkxE+G
imYjEXJ1pE5w2lf3a05nIsEaC5aZVdeJWjYHcLQLziBFS1kEpON520hU7Xp5OrqcI/IfrJKqo5dF
0xU0iUTITSkAUfniz2QhIhhcWt75bDzcvgwAYYjMZy9GOxbyLm57nI69LKEbnnGJS4n3oEuKxeBy
5qLy0Hau9xjKgL19A1GamWYBEbg8Evnc2lMYEif3urcJgp6KWK0KUdOG2etvucrex+yo8+qCrE2z
D08MhKjv9qnlnkRmpPJjTvQdMBlOCgKQk+kXI/yD1HmNzLv9zovuB7HJJgjvCA3V+aoZKyvcOnsR
NS9kUkb54tvLMqZWIqQhl5GmKSdkHufWWH/z8HQMARashI8NWTflO+wxnrjpSXF5miZ1hDkSFgnQ
pTifjFmsB36NxQNNPtPMPdxqSBaYQ2UPnUWSlrkRJFr48ypJeNp1cL5uyM5fysjZCJzbO0ERAuRd
9epkccwnlRnCGfFj+gTxFDcAYl1ekmv34rtKxA6NqR5PBcq/DAuu2NB2l9to/hfjOJQZGG38jCPj
nGY1cP12/lyW5WwKUWl+/vZPZME4EStCXL7i2YpRX9ipy+EF7b0igG87i1iGrwAN9Z6GaY0Z8UNP
4MFw+LnL8KjiTcNqG0fesqhVUthZRWqQj7x9nlLABXm8AkEQRUZ2PAaKRsSXAi4bWLpkI1mONKlp
rwhy4AUt1l17ei5DUHkz7/OQ0NUAkk+nNCrpOtgwfHf2MQLWKCPxJUr71tcb4C5/qFXfQLDu5OpL
Jz3Ph7YrHT9IUrIxfek2ZIQ4k0KN8gsNd2zqWxngEocEfrM6W9StHdUfZOMN87VSW6gLeiMaOLxd
J+mpnX2rSaNKxEDgVZPk7/12QSa2EDxZO7EcPwweTow0f4SXiOPQqyrUWWbWaXi62jpN1niCK/7b
Ngx6LL1LXUwXv/QWC6zM2KAbXmj9tblkr+2QdGd8cVs4bNaY0AC7pvjXHqfcEuNllX7O2VCizk9C
3wwf4aEOYLv6pbK/UVYqJr2dY4MaOL6sf8oi+XbiFtCwnVkVWw8UM4K3AmlxxcqEClclPr2R1OVh
4mTYjGpfrkabdDE1Xc7B7G3s/SJD0WFvIFF0VFg3juOorhDePdveDONBY+lzBRja5xaDDRw7OIgo
OhtiWsaBmGFyPnZidbOMRVu3w/2+vNBTCLD6Ud1CFyVM8f0gqJX1vawCUUp1piTQ9/Wt4p0CUsDT
T8pJTEJlLYR90z5iyijR1yr4FbZiB/hbp/S1sUGQqKcl0QTod2zceRTmz3c9hg7Q/k30psq1WRd0
1vU1VJ9W3xs5jWyDx0MjfWpMczElOII8T6vmbslljTbZDK8etUKjNsc7tzXSG8eVQ5PnG9DnwDxT
CbOfmAGsPis2wOJFILQ0RNcm9S3Y4J/ufM0hZLU6SwdYMDqfyHufF0R5au5uczI9QOYu3UY3Z9ne
a7idzZkKx5crF/cPcIaUUw3iDQ3IO8NYus3ZeeczFDgFt209DJAK6ckLkIHKKL3qgHAAy74ViUoE
nZBjTaooqeos110YRgMtOwFu7lL4AXILdncXXZzOr3yu3wmxpk2xJ71o9XFrGoKyrzYNYe6jkLy+
Y4SiJr8xw6a9CYXLsoscigQm79uowU0A4uqVikAaXR2tEKyXzdGu3iI6azN1yv5/urmMNFI2Hqeh
dMfVw8798O1ZK0EvY1F5AgrbYNbuwWxasRrK68UUksiGehLCCxDSKIowije8GNUb2suP2QJHpxwM
EJB9HUIhZ+MNYiN8D0PgRDXTB+e4Pf1sD8yzsmSPkTXqyGS6Uuk+VL8+ZJzlBcJ7FpEWaMMJxsTj
00EIASZppCZnx96vilTpYeKA9jLOn/6Qn7DSxYAApK9HPN7NeEOAPFPyLHlN1Z46AupypLRIXJP6
8Y4sryMfUquCTIMtDlcqAVIfheFgoZ2+3isQ6LIo0t1lpZ8HR61bjXboWn4gdHNAo+fdzSFDjwCu
9rQf5raEJtsDVrKdSJxYB8uMOnEMrAzx5Xqy+5u+9thgqUtzzTWQBo9wFqfhhjg1asKCEnQ1h3/y
k3lCNvg8dpdRajRBOv4029PUqyOYNgfbm/M53S2X+cZrJo1ye+EuJGaW4OLSCDeDQiR+gURekJ16
kSgTgZv9RelJs3enmA+Si0NxBBTok2K+ofDL7W+m5tkK5sWl8FqbbJGr4jldNNr/87Wb8LHFF4/m
6OCpgECunqZq0fEKcqA2ZSwIDq1I2RPBUEpSKS9FSpRe/c3fTO0LGC3WbqmuLKuVnTeJn/ZNGKHe
tVfdI34ARi7QKWs1Je5Lr9ox1QhzKsFqR3LuwCeNH77Xtblp1uGRJLmlWivfA6ccIL82l3qUn9oL
wKnF9ziz61BBLhR84Nl3E21FR9CvOf1QYbCUxkl9k0OC+z6CmMeGJjyN5Jg+FAP8LdW3l2vHX9js
olV8jejGeFtC8ihTapsLV02bZVhzZXmWKmiGmnPsBW9GiuJFO6FhrnZlT9Ym0Z6okXwSD3DH7k0S
uX7FKrVGTdZg/UuDV5pg4Iq5LKhpLaU92u+J8whVOSJJ5wfmXjVONlK3izfv2umQun+d7WjiaMff
K53eWHpf7242kuhZVNTcpVepuYxJI5QXDBRcKyRNFwP1I06XjGmCbPVgEVQsGzNjz8X8G1UFrRG0
77KpHvqXdCR90qmIrjbMQhLB1A==
`protect end_protected

