

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
g2RN5TBir43ECxFrT/y2GRXX5NGDYpjq+n5gxNTYWsuzDCjF5YeYUisYseKLr1ryeyQynd8Epzt1
V06LipLPYg==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
eJKP4nowQhkS+sdlDJ3aF081jbTFWdzdlOBNNOlq8qkrol2Z2K32WIgnl06Lqx6yc1xJY0X0kmV8
eOkRE5vog2ePPioAy86OAcMONOPoHTqykW2qaaCPwvHqEP73jf7t4R18PaTf0PZeg4kzgW5BQXqF
THWJ0viu+pagUeVYQuI=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
MDIZ/fTOzwhXm05ObJ3zkVB2FpJAN9o34cB0jHfFprFQZmUeUQ3tZW60svZwBPLmTXGm6NjoSEnE
d1b16jr2OvP7e61sGc1GOIzSD5lAxq6KYGFDCFGlb2HKuXZP87xm86ePu57tT4ld2oGvDNavbknR
LLxhx9ZyBV7SuzGo3PKuxBA2tnF6vIEJkp4n2dqwXnKJw+xgySn5xCMvJuNm4ghYOfBAsNQGJ39j
9OlCVz84SN0I+ZhsnI7KhLpJBWOyFN5hfdsD0RVsTRLOBu1rLKX6200sXAdAwmaB9xg+3o0vilh4
pIPe6hkIVYlfHVKU7Znj0kURPqGkJtm2RI+CaA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
RvD4A+WtjqxHYEUrji4gUWEBsLfMuiFWzgBi0pzOF5kWQsF7tHiiAC+dbiIZv5TBKh6/SeRqqj5f
up1ybf94wq9EXJ/d1afld/HRqNac4VRPTUzPBHt4z5dEncFPVDK4ucOaLAd/3B1aieNd9xn+mBS/
wR5gmSxp/s9f+zaVsS0=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
NS2iEv8S/DLjr8oIhLcaUy30De4W+2t5q2cf287k87h3kSCMEoBnjvcyRcG6CE1IFz2i6ewnJ0mb
4oesPU8Xde+4KmwGSKnw2OpNx1aFtJHy7C5xPLKHuYCmY+9zM9y9RMguGvxUNsPvXEO9G/4BQZtJ
xHf97YW4qiiYtbOsAO8R0m9UHVOYT94pj/6x0Itkq5yeU0YXuubMwNfZ5ZRnrVKNyxQ5Ilm1kGqH
N2bcD8eyFlVJydABBBV388JKwKrfOh5ZHUd8//7U9+6XMFYO4OGZzTYmAvyyO7iRRKEjPElnyW25
UoL5ziiALbB2biJ+eBPz4dgChqDQ9nB8HsYg8A==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 16672)
`protect data_block
ahFrAxi+wZUlxFn6mYwuYXQIx85JUs7Epk/bE6/h0+U19jMDEiGtfp5vC3/WTlZN7HDvESAp2/lK
5I7CU40pOWUtbRhP1tiQqZF8/+poB8hJgekzrR1TxBNf9C/1Zd6Jl5Uo6K0btotVLZkZfwt2PbMl
p9QX+cZW9NByiAzUV90NVSHVyR7wxkEGe7ZYIaJHHFTSo1JYCDMsEVL95825+8IBa3u9h/7u2CaO
+eUcDll8Q6EdM8Gx26z1U6unaceCKZL3oM2BmTrguL6gFCtHLpr+dsXyjtyAnVhaGH2z71PJR/4p
TSgv9BHiu5sqvf0U+Gk287Rmd0fppSlm4s9STSMJpOKfN+4rG4L9Fw2YtPlwQ0bczTSeaK5QDQS4
xIBjTdINQz5ElezG3uh7UCt/UnQ9ce70g6cUQmJbh5VKVhcPNnF3ZCSRm3dNKO3qLWx0Ha36lkYJ
Cr214WpHDoBvM5e1mg7xdJQQVvKvlBiurnqHHmALlIeOSSbErRlFkY9UVSxQh065LYChkmnNkm/V
XxQqXMX6L0ht2wWFRounyrT4RoyKoRRmFDfyCuEPgTZumWIMov5qTt0OCp7fuX+HA5lCSXvDh86Q
gf3/yZ8RLJGo4sqjgsLIbNVUwiMBasfRkjMtzDSz4ylu3Wdy/ZBCiBOycij9dyghHagP6TmeSaPG
akAA0ONrXC3zky4ul5FCLRg1+ft30F7zofDUfTIwlGctjwequnXmu+lgOX7fgTqIQQJ+wjo3AknM
XbHhvxZSgz69uD1YxRSeB3aDZRpdXBR0wSwEliNHXxM+QKfxu7V8HsZewJfsIb4iglTnS8MKLcP6
y0ZPftm4lM5bZgbrJUC7EhxrtbqqFHCWsmL3OoPSHrw3Niq54yh81FLiJbEK11MfLWO4G5doLzNa
t6FhCiRtwAfAkeUTBcjTpDjI8WzlKpIEgySxSwJGn1e2A7pTC0iopsI7x07W8R6RTrgPe4l7Bgh4
4nskPKFZrcH6sgIQrAqb38INrWjb3nQ/1ay5e+x7qTZmfp0mo+97OPEDajj0DbY42ctmaGOtQaYo
upgGDV2x1BFYCyhAx1BKMGQOuAdPpIGslKkiwxN+KBThzo3CwgGpnvyfbOTYE2TcNRYl+pjj67Ac
uTDiR3NmVA7zIZ8YfaXv5SzpUxXr6D7vlqzJ4Ht1ijxwuDsSLB/d+j4hPyX2ZjNzZ0/iNcD5Y2GG
qdWuwhmlTL7tMnOiXEPBI39KOq4zlNoviYBfTMDBg7rDcBT5+dP1/qLd7MquoG4gntMeUtWFWa7j
1eaIyIoRSG5uKivXt3gey+0Exanpozm/UVzVPrGXHJlElIyawMqq0msS4GAan1CUH+/Qo7Aod8ye
H0p/vrXzFWsBAOjJm+65ZqazYIpW00Nyb8iq0G/0Qzxz2TyKgob2HrDuIsbG2E8xhGm+biKA4x1q
GghO0HVQXXe26y/MVx9WUpLy3DhjlbcgKaPyzSnlnVAQ2wlGDfNd6DVCfBqBGGCQri0xZ07EMc+u
Q1+D0clVKed86Jfd6WetRwOudkHBAJkHBR+jBvPoMTQJKf0KxvS9mQPOnhXIoXkzAzh/VTcgugMB
Sxrb99m8EPeaLRpBVKWIkKTwH9yCcWxwOz5YtuAGnTvwgVHft866s21CQpKa00f0289QzQLa7wY/
/jgC1OfnFR0VA+rhzDddL5Ts2BHpcSPv+WuWAeOJs87lIL+gtTXK+NjBNltZYEONTcEHA+TGCGaF
rMZAeKeTlfsJrX8qfOL3QCcW0LGfiU59RtMReUtwuJN2sh9x+Mu9R3YFoDoPnoYh9KE/vNvS/hc5
XkPF2FW97rOD4Ic2W7NhHgPAb2P2leodFypxvUPtDe/AtpvqvHWvhCH+paxaermSEPU2mm+5gVq+
DC2rT0s9xt/97dgmerG7E5J5P068k8gRLX4Zvvv34f2fcbtyU2no6aQR/g9XyJe1sX5KdOSrKVPP
XDIZ4CvCWLB0E4AfEy0Q/CpPW2qs4R2rdmxZ8ktY/W6mT55CEzjDqHUpd7ocvZyL5RmX9VKfK4El
2h7KMigBpXPjhUXlAUIxekM7ReanKO2itCvG74Pv8tT/vIYIn03QSaiciBnf60d5/Fdfqfci/xNC
B910QrUIN3i1necU96/Ybxb/8Ree3yg0tRFpu6d3AisUiki6ReT3LcPYMhERiit1CLkMWG+L/0NP
WhG9RFwCj7sWLmBdpZDqZYBEz1qhFUmwpbxCO82Kc7FGoL3Ot4xvSWPwzBQiLiF0oQ68ueGghul9
zcRUw5XAEt/lQIEb1qrIk+hgS5n7GF9jjNRsiHtPhCiOmrJTAJUOmonTokeULto6/LzwEP3bFESZ
ljoF0lwqQdNCDMTA7iN1E0u7y/uBbLKHGMSiVIs128+0a9w/4HiOYd9K5jyB3DrHAYKcEWWq673h
/SRbgox88LJYVIRjVsq0ZvDMFB5VIko3yFjP3IZTYoyfXLYeOuiS84GNKWxttNWKXiW9MIaAmC1U
Cou4E4uQAy/Y9n5ohuwJd66gZRD1Esf2Gx8/sARCGyRAGCV5a8o0a+SZ6WEJ2rxgnkH7QM8vry8a
4W/8DFAdf3n3W+72JqmPCc0l9Zi0uRo/To5UB6mr4z0bobF7waziZNLF8htHn4eZ4xw4VWi+7TXa
THyS//f0OT5Gr7kLwrKMAD7UP2SwN9lXt1TQEFcmY2so2f7NrSJXntByupxoW/rrsWLISdmmjydk
/tC0R4hIRTf0ZwXSqtReHG55JYEwomvbSEm1D8riO7pXycP7/jLFGtZfO6udwuFVX2tv6oy+bPSR
15HIzzch/7a+XT74rOSv5qxC4J4ZXNbRw06PbzMkmm/fU98pnoYpG5cuUaABORJJBMUuXAsUhAJM
VZtybfr9OzHFhgx4wkykNPxmOMuwPMiifbgqf/zgUJCH40Kze7lahEFCxfrrFtDb2BHYgMw/S9Qc
aPaVvvCmXZosHgzErFme1JvpYH0X0IvZbOaKDlkp0tnd2PECtJLChEovCqlrd+MaiWmPpFMA/ClL
1AiPiUfWQtC+ovmPlBa6dART3tgW+c2P9e23a6g5LqQcF633LAshW7xw6FsUmdBXne+DGudhOn0l
AaP+VDjHcgkCwViCcPsZoUxvtLg1vWXEp2iyHpwhlUokhjYw6qg2CYdzwfIB78sECK/gaqskt3Ns
b2fYNg/frVppDc2g6VMeezRSkEdAVsNr5jSIBpl24ZtOE4wX40k3LvvK/axcCK2siuCn2fRkSssM
hcj2LP5jJxb+0dMxDYTKBPh+KaoaeXSb0ahZwXk81r+eZg+fBdeTNQu4b2kx4LuU7eF3hvkRdK2v
ZJGw93t9ZdXIETSMISl5GxYaGOsk1uQ8pqviqLOkDK35lEcyAGYL5DYr8jiQmkfevOhYqKjxbcPE
bRVp1NGETOwgCn11TZHUOXD1dmpmdNJbyIhWJKUxLgXZfdLG/YGDpd6iRxxHqEwaZmJFpctGW7zI
b6e4Gvj1m+qgDA5f/MMN9SPqS0eM1C2w8i15NwmVaVN0bmfMIVnV/Aez2AZ2FCbZsSxLTjoNfNQc
Dc2mofzGWPmLLwTERkAGeDl8aiGuqrZ2W+bZwVSDT9jFYZ3mZgFx7mCFuNEfJco+7M2NP0uz/QGa
Xilkd+8PNCt8yN6OZctBnKMp3VUo46E986NIjmJF4RNsWi4xJEEHsyBs8vfUMnntKt396OJa4//h
USIqHq14fUyYg2d6SW5LKEQEyqSy5onN7BlAiJXSfhDn9Im9wGcwW+Ls7NvPG4Cpm1IPSiODDcn4
MVGV2ds6+UYwlElToe0aHBX50B0ipDbL3lYCIAZgsElqm4uBNtDT2dwXGJXNVVQzEd9LChsZ8sEj
+R3+QOWEmI19YkcsPSf5Qo6qBZ65ywpW9bpvLLX8z4kLGVWzp6lWWM3719OqBdteiAyFry82AakR
CpZn3tVbChLwi3N3X1BxpG6sxkYU6H1qsoEfiwSPpkxFS+2aAaArWWDs+GNOtDy+Sj05TjUNKN9W
u6DuIohSAsh41W3wAlOvyrg4+8iP6C271Elyy6ikUtpZpZgL6TBJBm6DfmzHn0yk9t+W86/clMqi
zx73cOEOqgbhS3p+sNIIjoNM7WSybdU4GuRSYo4M2GeQ7RlEYWdenD0x+P6R2qmDtw61v+rXvgnc
lFu99nfoIT0mDvlpXjxdmp88Wo0EOTAg/dvr62LoZvtIsgpQ5JXYpf7Mzdjppml9P8Xilb8EUYMo
2+PkZN4wO6K5E4GRbIvsbgN1ETisnepVqreKAv9/Pm2Ooidt2AlYdQChG+mAXEcV96g2SgfzMj/+
7l27n3YW9NrLPQGmIVPyKsel74gahYiMHiqAH1jXO6EncCzxZ6Ttjn7x/okCTFOcQwYQIrB4DeCF
3lWyBBdUu5xd7sgsK8iPxi2iE8RPutZ8kL1cBBIgiIfAgGHsl2tFWVfTlgoaTybQrLMOLeFUMrk+
Naqbh35tW3KIEq1hZY4UFx1fkks59qKAec9AmX01/Nlr0bomfeE0K42a2ccI58mThM1J1V+NPvKD
LGDoBjmTwC6Ei6IzjKQ5+sOKvuSnEooScDQqRYODJ/K6KyMdADzdga+jeSL78jYH807lxb2/MXTe
KjAvjAojNK/toUvozasX5VF7lN8SMnqcnSBfZRiQex7N3+j4H4CbUvyGKJbDkkWdeqlo4bchlfE9
T6j4gm0G4/dFVgU/QGj0cWNZGwiQoc/YJtJSm+jn+soRo6T9YDAkQncGr429p1u1XnjefP5pAg/L
6WKRb+Gu6HMpV15cOBV3ZVrprmgMLOSlFThxGFwxT74bG5HO7o5PdqccDYX4bJMn3oLbnALeHz0g
dw36Z58sxQExZJ7zALFJJdPrtc3V/F9mszyYbTKdzL49RFJ1hOVxXttFTPFG1C/SUhjg8ZFb7VKC
ky0xZ8JxSV9YZ4g5wUwGngJGoJ+xseXRRH6ioyy3YkHf+aHWMRtwH/4xp6jSCdnq1KrMJmXberVA
NpMF2G/OYQ5FqBg7F5dB2Rr6nJL4JD19X6VDUcc3Y+0B7bFj05Yy8apLN02JTG/F5v2BA8yBtj8n
xLWF/D9qJz1j9MziMVO8VBDO/7AY4Ifo1wz7N/puzw/iScsug5QRewe3gvu0amxK/coWshDKKIm0
R4AhNAfPN7TA/7SIEp6VOQL2RF3wVjZNk0NCJSVWd4oSAzJgcPSV7rSXNNQjesyvQzQ9uCtiB4sB
nfX88RF8M07HrQR2non9/MJBxKpRY5a1FBpEgGUWN3orYhYUw7Rd2Vpc+ReoAzsVRTcWNVumS2xY
jqctIfj76FCCLahgrhcmHznFi8RC01u8xSPgfoYcs08SWA/gCUzBPriGG4I2lS7jfjHYfu94tmrt
li2si4996Kez07INvqw+iYf3h5MgiFeVGuSnFJZT8iC3y8L3OEUXjAOxfarB/BuZhSRRZU32EBKD
ufsA3s7cp0edoEHYfl5kVQdR2pvVDN68dPc9tErfjlZuRMWjD6kCkyPqC4CaIfOH5Bnth2vvbZ+a
yLYLNInp/0RfBeKnGZMQui/a5Fi5r5TaMK3wqvhFbWKfr//kyLywEbooph4dZjvUIwurAvQWG2W6
jgIUirjmX2Ozv5QVVChVpEL5umhVAfpQ7YWsGrwu3Y9+aot6Qxe0mAFXr4wc2UEZbjP1+jGilLW0
IaqboOocmmsn0EOpXdncEJAFanhPj3UpiZ8Mut8NZiZgIKjq51ZAU/0uNeYWRs3QWaxWKOHv1ia0
vaCnqLcHwX/CdvoyVDKA0m6LZckyteDA5kR/94hjCAgtgr+RzZ/L+ZJTrXQHaGaLOIlXAAG9A7fA
gXUXVhu2iuWOAxItEy6qnSe0m2rPUOMADLKX3aTT5iJ2w2wRvcBIl1bLc1UL1moScIRropkg1N41
gk5k70D5imgK4ETknWlhnSx957rCEYxjRsST5foICgEm/9Uk5BUwBLWOYqHZzILiUE7zVzPa/hsY
7VwL6kGoE4qNrXdxjm766QnHBN5VVSqAhBfhk3q5ERyN2M+aCnV2MUN4KCFaSEjgkF0vb3DGEGtH
ilTKoUgWXm7b86nwNMUi+70dBplYldbQb5xdG4tMND0cvwnm4d7UizDSxdOTzBj9kVXg8zjiKAJ5
Yu4+N/zIQuZE6morYBnJF+2pbo2Va9Pq/HVsPboWaHvew1hzvCY/JpNbPqGJ4RaQO8xFKKNeVJnc
cjtzqRDz4bHhlzdMzdmCzKa0UCgXJEJ9wXDIf9Rb075nNA3IyM7a2l+GwemFKa6gMplBhXSSTWpr
OUj82PVJzoNUbHVfGvJ12h+9o9M6Uipq0c/Zk9XcZYXDjFkePGdAgHed4uhs9mXIzJEyAv9S5h8J
oY7TCQLgOTPn+MJPIdanVL+Rhe3d1BWAxKJ1+L1cbBMzv/fx7jacl8cHuRRHfxCjE/Uwn07PtHrs
fPpOjvNRTatJ+Uk0L4xpV6QPyn1OC1Da5I+TPRTJemn7o4ca+k/jPtsR50JKpcTErfO3YqoYRz+6
+3ImvYnN1YXUQsTZ53Hy3xyci/AEWuXn0Tb7F3410G8D1E+oUFPwerHMDVOdwlblDLqAOxWscfPp
97F6bp8JndGyHZT+1GbEgp7PzFbIB+guCI14NUYAlzmKve6vLP/c4AIUNhW6+EQDH6e9BmOm00TL
XgZk5koo30wnroVau42t/jo/DQ9iooSk5x+n7NJCDPbLnPGsULjMFk3A1I/fzuoHDO2NdlOK/DTI
CfCgrGirvnGifUFkmToInc1SG5VpYOrB8jRYun5n8AwqzYnUp9LWZXkiJbhExjlUdKmS158c7JOP
gLpqzBR1Buc8PJAsJr9yX2YUnIvHAontNru0ng1XCWsnNuHHAizOw3RObASlK8K5rorgjGBx9fhM
PbfVMPVIlpAg9z2BT8tUarvWfVi4hJGu1id4UULRdBQBJicJ2OWviVSyy7PQSkEKdjL5tDvCY8SD
vUurrUgmO3tcHwaqzQxp0JEROyw3tD9dDjPSqfe6bXDjLrTKd8e5sddjgxbRAoSPJJ4ObPvKdSID
PcMuDHJE20XcNVIeFhzlINgGZoa/2aeLYkeEB1PtY9H9i/Tle89UWnDPD5XIdDdzNBmJ9jPyFLo5
HAagtGRAfifOU41vpTHo6H9lKCKIAOxqHOcOY+12kxT9R5Ho+3nkzjQBZLVqABZ6uuZMNllocnR/
uwalFQh99YDHlEQjdcuhyoaYeb141fZ8I3aSzdmPA7/6czFslkHH4Vg+k1X9ckJv6i0TjGNPd2fl
8SbnhdAdHeBkiKXDlCyfM2qQU2WciVMep3qt8MjY2Pmacgd1U+/sIkUeMSABUqeRsObbjjIiRSpk
uL72QgIWiCMjixp9VvZV/pN0YDvKNKJDkDIMsOOV/HrYikkblj/9mO16NJXbnI9LnnGrVc3xLuF/
82KtOoQNW5kY0ppWgIVftIKJEZum6ebMJIHnKzjQ9TkW3tYww+RPcldnG5ziKVw4MVCQkJ6CcfmG
PXFhK5gG03w1mu5RIXIrIwEE10b0OHq+Ehu791CJjhN5JR4Q12070sCUzzHXc3rLYH4fYSOqDYjL
YP8if5JNaFy///XJx5WwEEnBlrIFJ7yW62oDrLVWrC7ujNNdux2DWRaITQdLTiEh87Zu6m1WEDVi
W3HksTMq/f1qKi7vRFj1DJw+n1/9FPU/ySGsfg9IrwP+W1+faK4tiocQZrmR5nI+qtsNoVpmByV/
ll8UscW47FXR/OxjpeNcmeRZCHxl2UDYyTSjN8zuxu00la2D4hYgAOU0mkVn1XLFyCIFfS0mPftw
ZVLpkMygFoBPUAswN/15CFG1t4dhFc/VWIMDfCOg8soxg28W1r/+sF6jyfX4lSxMHXbqoN9VNdEg
8GVhEUAkp6AwAIjO5fCZg35O9MjyOI7Bw3Sctcmbrva3DzC3G7jDyoqOgKpOtm5v/IwQsV6/YZ+B
41OSArHZhe2O8qMsRUOJ/75TMBAG8R7Qrg2MFCCmJ1CnvsJfDjzwikwP0Zs07vj2i4iFrDnUCxnw
71YgW2hFX9SgU4+px+aCkZvnz3u64PAi3I6ddhzsoAytXgKneCD6ztmn3BgVAw3qeYlf5GSIDXzW
h63wlpNQD0wA2S+PBRowhdNiDCaVbvMgYsbzprN3mW891YWjjijySH9MDXe4xLsJSd8vLskDbwlb
BP77nuaBXIAnKgcPx+alfHxLB+BLpJNkQD7gQGCrB6scsOZED/prkuwcqQRWbbmy5c+MwyAfAAri
KBsgIUV4rS9Haj2wY38wcW4KkokMt78rC0d22ZK0BUSQu5DqsLVFUbXaDoxwjeiqYPlkYnBs+e2g
lnzhUQt+Fm8bSxtMFcFg+xlIKGKDif5o1knLoSWPM6KlY12WcXvWQYkv4sv9Gj8+pp3AT25NEKd6
Ty069f9zygr8W2EpVmLJvxDFTz4FuKVLVMP/z9FSuEL+7LFDcYlr2azbyeGHjpRN+GucoCvoKT6A
AFPJcW0lSUpSF0l/yy9mdjPvX2TMyUKONFt7HTJ+Vd71h44eVPbYYHg1uosVPBpJEMiJ3EkkGb68
09u1reDQ8LPTy9A2CzwNjgDUS82BdiJyAMOgzRQ+GJ/HjYB5lcwjxQaZ5voS4hdbvnd6rxtHQ0Cg
BZ5VNbz2xn5m1afC9NW//mzUQ4TAg7ayI3qKpr5hBAhzT/TtidpPtN4vlRpJRhALjcOLbi083Kms
d1u7AcDgR4Xak6d4A/Zlj6AklM7mtp5p6I4EJZarlme1/Rm1k3r/7HIuXnX70INMnE9k3CIKJeFb
guZj0DrlSRX9iiZwGkp28guwdpTv+m6NyWir9aIrE08MA76avmKd8JJk8TfGSC9MBuu+flF0jBY5
Vge9gKj7A7ueMk5GibxRGleRjuUAYd/e4HiWj9Wke9FO8FjivIUXTtDPYC3rhccCsdb8bjR2f+ZZ
aFBo6OsFLjRik9BzPQ268ZNbEgZFWNTuC21eyfRPW+dJY9j4Q1jca8E7phEn0FV9DutIddqmgYMt
goxYevQNrp/oMklVZSYIHxQut0R9hE0nbEL8MMXy0yucg6pSQO4syfty+4IuBmhuIhQbXhAN0dD8
wBq4GlLe1j1txdMjs6UHrmPq66/cFL7QHALgnPoY67QUOAkNj0/LtnwlTAtYtIZG+QKu0qnvqyuu
BFi5GZdp9/r+aKMIhZxmg7RFXCiG0wOe83pC4/AD/emtfLoz4NlEdMLhI/YdF09GqJVpdm8+8cOB
0WLUlUtli2YGFZ1leehms9zzHQMrBOUOuLn1+oWPd0prb4EB7Fx7JJNGICMba4DBeoc9s9+LojES
jZmzrsf5ueevYQwDV9G4JlGLhqN6QODddzWOkIZ3L0pLbVuB7lKPAXnRgZAHXV1jTSvXXI5YsQ4V
APAiXJq7ewCZs7ekcI2eqqQ99MOjGghHn5EZWDuUBtgljYUWC/gJl32x+9DAK36V/YuVVTW3EfZE
V6pamVhCai7/4QDRPf2UGBTqMvTs5jcq3Ez9/IGqkD0XPB9z/CneHS+v7jKONEm4WKAQKQ9Y5ahG
fWM6GC2eEw8YNp2b7aVFgy9iDjc2gD5Vo8VU41tedl9SRmlSU0mdvkZbaSpHf4YE9AA+z1tPpX5f
YZkHNia1bqZJPBkGMaA5DAeI471zs33Rl3gQvS1HMfsTbP4Q49lD38W4sCrGZfsJtEUQpOovtTMi
A8pCEAEvKTrG+kc1a52yjpd/oWqtOpDHUgUcqUdi5UD+0o87jkXLOVlwI8m5f2fj0GaAi1smxAcu
ooRDZTfI4YmnBzuS81MCyANdYrW739PkF//cMPpt8aIZRbFdMkN4TNZUYTkDsTuEcy9TVhyXJeDG
kpisi50xKaZrxsr2Jtn3wtpAtFOkSmpzfuDG++ZOtdKHbMjehcmrIEX9SthXr9jY/PiwNCx9ehe1
q+OklY3bozy7Djdcvpbq1B8DzlRsVKZTYln3YYfJWzVneGeo5tMA9byrVSYEcD8qw7iNdgiedy6M
KnJL6c3HSqTvWQzcAJJxu+f9h4lc1JHjGuzIHjIhcTl/H1Gy96QKA6fIv9Wx74n2zbzKrk3Xlobq
akFadh1avHaQR0zvkATFvVMIlqnz99g+X7cGz9bsfJ1ymRfZlKjkO83aDWIeax/it82BAotSlJH8
lPxgxW3czJAU0Tn1QrBRo3j5YSNDgaJjRXfjihtHPYJ7XIjvLzYq3u9YfdaTMlIopSj7HobaTyrc
4RjQxDXzPUePkH3dk93JjH9OUPwjkTQeVCf4oN4pDW7SLlJWqdouk2minl5LVWpo6DAef/igZLEa
YWsVgmAFfQdymzh0xIUxQh+DCBN4NsskmBqY+P4k6hc44nop7owv2dvharT7crQp1UkKwflVZdln
Bi+eCkPXDu5vWg5nVfPWSfpk9/WmzsLfaAVk/tA72Z6JugTZptdKyOsVmE6Zd7ZhN3E7qCZqc5Is
2YBIkKv1hdwJ7o2OdR0OtGNDkF8FOm7MhB2pmDX4vdqcYg2wNI88XBg/ymtWmBFzD20Sm1UWc48r
wQL6xtZBsBR0VdpYom110uJR07Y+fNzkudgLHfHQdEHiPRG0W7w1P4lNHgKCAQudzwiqyxUOTepq
edXU/HEMcVg4Q/LlgIDUESgNmgQLn0CLJPLb7zy++N83cN5qpRmn7iY18hkO2y3gETBUHLAdCaXO
IyAaohWW/8YrbgTaWPfU/c4sCRQDc8dwHLSwR7ITbjxRWab9wQW9QZP9259ziR5P2zF7NQ+M4UJE
ictFo+Wx304pFN6nRrFT6JhX+AZRclrYfkxmCWbPSq/84Dpro0mpi9dqZMjTHiJus43az/7dsJXP
2VZaK52D3kRSea7tkcFTCNGz2nQ/H1fdj5k0ByYJL6KuNDJryj/P8grV7bd8/4h1o3TI8vfECkPF
gwVOakTPWz64FZwvZ5JuYcVmDQl5+tRjIhkVYKIV8Ez7gL/Cwuj/Q8hr1yGBC19BdSwC4AUvP0XY
3S6CV2nEHR/n8MBpoEllQ0Ici1DqVfgJWwg+mITeF2Z5v8fBDiSxqMtEHqAW/Yjoa2hqYT2Y4Ms4
C4LhIdI/9PTLRyFbXUfVcez+3RJQGlidHR/i0YjE8kokaEbJ850rbqEwXTnVGcymF6zrMODj59aH
vUf0Sjc6sYeEgIStjEhSjHLQ4o5B6CBVmlVulfJFMCwrVZ3wn2oGO6UWDJLOaIZ3pTMOHx75O7Es
ZJ38RFKobiN9cU4X0HoSpWXZXTdlK9mYPkLS9jyZxwkIN8VPI1EBj/kizogTmzb8cnA1S4LPN1X3
dcGIqfyxR6Z60T4fY+FKpeL5REkxDwIXJ28Aka/oMdPb2BYTfInhqO0YU7IT5zM5OMR4rGfEL5wZ
+yoUM4zLn1FfY3vELzLhKp48HzxTIXBfHQakc2T4LEfPylpcZbm836citYJ8f/32A2wpEMJUEScP
zxWETUM2CltwmGH8S0yh3huAygoO4oDnMFGaTqlxsaIhUTiAb3UjvkMxAMOY2w1jso62KcEeKiZ+
LQtj9j655GgGshgcI7FoOgOENVwVN9wAd+xTlW+G7OsT73R2I29jnRhwsWnESrfw7/DTHwnSqGyS
LTxRk10BnKxE4WFrA2v+tHJgnKrutECvPaxLNOhjA7r/FC05/PLz2RDQg7eOfwThet0pacGWv6kR
zB9PpSREovhq3MxUtagu+0Czjx8FwP6vszllFta8CE5TII2JetFYx/CUeQZRex+BqyzcmuqBahm+
p8G6t22YDR0ubtncp7fK4K6xH9MC0E+pVqYkObc8/jh1XXv9TZkHlXL7bOJGMYm+P6s7RP36gS5D
X/Ya9lpt1GZtF1UqZqb4HORkhlR1zEp9qcKJoDgHwk0yWBQHMNPlz7gjJV+CeGu5A4V90dF9CGGp
jAZwpapYMF1Uc4f9mUeLDQvQ11JBPcjCeZSdgjadUXT8EhRkhlP1tjv5Z47joggkWjUnmZkMOAeL
vuSxrO4ahp7KxE8DnPXxml3yeWT7wD76VARAyOB3jUyO6Tvh4/QvymXtNUx5BWDKuXKWgMEvP1GQ
ut8Ht8GyxPTeFfd86KqICwYO/IUBTjGAXz2xZI4TlZLwA7ATtVvy9kFRQLZ4SdnZunRyaWSCyijB
oKtpJ4Vftjoi/smUMa/iA/hGGhEpDstPL/SzBZJcBkJULJFheZuaVlGPXLYi8Zi6VsowXDNG8pfB
DKwfFq4X7T9DqQYBgyD9WDmLTkQUJL1tp6LO46lJbgSftrMq6P3KQLMrBEm/v1QWi6EbTDr72EhY
ewFJ1jMmwEIbp42xQbzH7p1pOLRL6ZB7v02mQ3764cEJi7pGGetw6ztgdwoR1wvq9D0qxmvYVkf0
EQTWIwvJS2riPFMV7jRUTFPgzMTTWh53DT4leGhfD7W4wasVqsMAO3RHMyy7UH3a9TNmJemr3P8K
0paAvZw2zbRtmN+mcXSiDn1xL96F0iT9gnon68bUYgh0vyQHjLMBnHJ/suBRZpf05mKkza0rm2+A
AKGXYt9+8v89gL4LxVDnfbtrY+tjmWU0LkVQ9SMTC+x/BQlxheUTY6FIMb2RyLR9phFdBtCBC5S1
sgID8HJA/kxvH0aptA4wKW/8HTXFi1jI2R6HRvWE9HLIq4JtGpWaBSyx4JIVxLfOEGJCXK/FZf5t
ENBSWmrHeAqOtMCdfXnQPiTsJKlopSST8OQozkFB6S5ILeROoblESouS+xbrqoagVWYxph0gAzQp
XfSLX2LXflPEeEQygWm3BQGITboTfW8dcs/I1raQjB3IK1TO780iVOiLBeWMTdHznIHME6poWFCi
Q58xgl2Y1D3j6xzElGii4A1QItC8XF12CKbd4Y8HRaBMmX7zhUO0CVgIfuEgdVhxr11wX1TK6W/h
VEW6LNN66ejGOWSSyLDPaG1mx8hMWN2dZKRBPnBbWLrhNmLn2eyw3z60hiDP2SEaFbcPenIIXrYJ
4EYHKa8YUb3ltsrlwqfXqv/nZ3mxjR/jMyVCAMZxjYhFQhQv+5SHiarc1KQpzOKABwdTaW+QBkUj
ETXdtC89qAdFniKoA9Y1Qssp8TqP92AN11nieWQrbs/cuSmAHzVgcfp3ne8xMigFFC2C+JdqWMPZ
Q/kMP5u9ixK7isOE/lkx/AUvSWFdonDAoV8+PKkXKSQXLgNdtIP5f0lKqRvvImZwzNUimf70WDWd
gKfmzWlYVXi+Iw361kWnXR8DaEE0Kd/Q0ism6VGKeEViv7bzRgbKVsOXtYtZWGhIVjysqWQ5+L7o
o+MyPwfk1b97XiMxHS2Tc89oup8MU3cIOAcN1xDpkzgeAmwLQnk0l68qyPUSWJRCFpx3uvgaAowc
qv32Hez/E6AlqSzbdPEUiPf7SI+sPBGAnZQdZOqNliP1FnKxZVY85MV1mpdoPkgPLA0MZ7+Ehasy
fZ17B89jRqTvPP5nbysMl43Vg/eWTojHrfO1uuXz8JL5UwCWTrOOTNqXCUeg7F16e140hEAN4Vva
uc6far7tIku4vHBW7WxdnaaSlUsLTXwTnoD/ZPmlozCmjo5c2PSz4qDILKXDCOG0potheCMAsQWn
svSimGXJlMXR4ON7bxx9ofCuKO21CI7KZzpbTvjz8DyS7ngHTXruOqXhlMofK8bUivvlq4LjswCk
TCj/vztj6loVKpNu2+w1vs2DivCa19MxQrPx9viUcCrAx7aGCAVgPmMPOAx88n0uHyE7VrM4RYIb
KgQAajXM2UDhQaaRMHJPLEhDfRxWu/KjNDbxLXOWsVLMbuRTgmyM6Tf4Ldr8Luj3lTGLjCrz1hyT
3kAfPYLkaFebMYvNYjViVvUH6en4g5+7iTGrCo9Z92pbDw4EtP63KuAICenfSxDX5yTsTWx2VHQi
LGxOJOCoBGrKXZySneeeTBop7FmAvzWCQs1BLowcKAKC2JANXfSg9mEOZuyyZtUgUPCB647Yk9lG
Bpe+gqCeaF1dBmYYcZHLINMbiGhhFYn2qEJ68/e20/NKd0Ew6G4mcRNZmqwIEKP/CTJ6QVSta6DQ
QKdLkcyjKTTH5KWui0S4QPRR+mb/ps3HQGQ13izRIxdrhVxBzyvqYBuOSoup0O/b/b+R3l977lI+
LBEpM1y1RjcZjocqdG7i/xVYlpZ7heSBRz86OMX2vtQOm5paK20wqCyZdzx1I22pwrIsfnMBQ7IQ
z1gSShPsyGvhd52qfbxzzar2dQ45OQZfbOHxn8Q/7MhwPviXYa3grsPb5yEYROn3sNA+jtq/YSlm
WLMsGTCJE4fHs+RhK48RJPsEdNVRV/KiZRYNaFljhmy1UPI/P8uAaOSp9Z0twpcRkgWTzQ4pSmx/
CrqrtW8Mc1coRDEtj9oQw3CPG8AAEFp7IPBUpyDh8Uo72am78OwrUGTWnWT8/tuKFO1TJPXWQXxO
KK+cCbEvD0zAN4AJfCWdcRiHQdRlEjO18jZ+WMhKFjDPkPFsWuX/OY2d4UlQOl8o/WAksJffulG3
QaVEP/EAMshQmWYmJtPu71UGGGulaeYWSjoP4LFf+rjFpREf8UDdcgSlVT7NbtEARr0ViPWZ6FtC
emyhGE5dfh/5IqAHaWiSFovT5tovjT6oFNy0Lec8czaRlrelqrUXmJStX+fiEM8hHCsvlM80kKBA
gKR+nfQyjUGugg7MiWU0+xzQXsRTtC6l24vIfoIAkkxUAFg/f+edrRPi6CCD/0GO6TIyWrISaSzj
BIiry84przHLoDbuK+hyu5a5bQGPPJbDXS9y294NEve/aUWiU34p0Tb1ExYjIEN4jzhXWTR36/XJ
P/Noh0JChx2ubCBUMBs+pHdh75pnvgbHgdADGbZ3K7AoJ3c3CGJYHoYvZN1m7CtD2a0jymFZmDfm
gPMObkuiAhN6y9mgcjFsWE13h2Q8eLzJycjArAT338Fav9Pa5iH80+/CAYHrgUprDNSA+gef+l4r
GqqZnh00AIYbknGkBRwYFt8b+NoPpwvZrYZ04qaBAak0D7IqOBmM7Izie7lPqGVkwwlXsRCmIP6A
pQvz++9gSYcW54dTDDe/wdvWKhKiuISsodtCeLJ5ip/zf9emWpwyCeJj47B4Vuswhx6BK+1TKwac
mELXViRvFkhIuCq/3pBtFVGLwb5lwEhCf+i/5dT+U4GdnaA6tf1RymrwFTVHZFs44P4RUGejmlCT
vOlqNbaWtJuo7zOY+kXhL5igo4BCyGVzFkjdHcZjLObk7KGQcu7WxMjlWh4BzzHzb94snHqWiOXI
J0gXrPh6RYIjDmDw+zsSvUHBnkIzRjgIYbKGLTgmweUOPebxFON4986GlqJ2buikz5lXxagQ9xhr
M+IoiuNXq0w4IBzHo70sV9xTiej66fRDDVg4L3lCbgurMoeO+avShvyedJa6VxUk9buC/zqwxYXL
owcO3BlDOgeOR5GzhZfjNRYAt7Jsi0h6cZ7YhQF/1brnxslmJKRv2XOV0Qq4KRJEjE8QnRdJPcv3
GxwEgVMKR4jwsVunA7Ky9AXoF/Ii2m93pL3Pm9HkYHlCkKHFkvVj81NGtb0HSoSv1lbSZKYxj8rX
iIlMXUw4OfuRpFhb3gvDChma2aOzvmoFwlbtgOv5hSzkN7f46sfcliNe0eGH2n6x5VoIJ6FLet35
vl2Bp6q557v6vKki0P3LZP9i5rxrgJ874IJOEgI+3oCzdT+Ab8M9roK9h6GalqTR3WsjVetwubqK
YFo6W+OWJtW+vri+pXTHGW9Elaew2Wl9tyso8dWUMfDI+q2ffP6jOZZSjtRH+cpwynJm+yhiTmBe
s9KKOOkUZp5pYcJdStAS0krPHlRlDTcRDSMCiPPGffFKhXgNMfuZNgfL2Px0ScmOv90SEBckbHCi
waeYZW8mJUbHqwrPjoHJHz0xs1VV48XbIN78UFTSBAbQinW/OOw2DUNIPkLzKMeX9yLkCxcCC5dW
MJhUfLuoyUuzrn8ZCYkZ0VUf0Lu7FPKEfm4intF2jtddjspGB6F1LrLP8Jb/jEjgI1XhGNlWAQt3
hqy24Onm2GX8LUbITzRYoQZI9P9y7jgWufhBJlbLS8VNr7T+pGZOV2BwgmKZx0ZmNDP6MaY4KIx+
hC2aYPxVILc9+ssMZl7hPsVbwHm21xRGdXRmfDXGiRxeealwE/QrIZfb9qa3HymRixk9DGIkje89
sULqMOCvOCdib5sztqj0F/km7YJdTc2bYM5NXnJjc/k2Y5azN1btsgqs5I2AFId0Jo5jOBCxZRcV
tB/0jY0vOGesSiJT/qpZVFlgHL1XAnKLqRjqK82PgHEysdNNprpvuBgdDai67NbHGTbbzGsJT59L
jUHy+HyY2Wv9uCUEQlmLqcd9Lx6hn2HSbx/LLjPgWXn1YlYlRBcbv4SfoJjK5v3hcJJieRZwMBcF
ydPRwjS9wTDdk4qGW0+HP9TJ1ijx6f4pJ6KXcB48pDqI5ViKzzy1BNVv5adLiX4fG/YXSnVu68mn
V2C/FkHuzys1YJemy9X+rqy46g7pE7KKmKRZClfh7C7sT29/PNloJfzkquXs67qCP/PWirajuu2B
1NxzqsUJByK+LBt3R5uAqf7CofcI3dDF8XdbQNSOWHLm6odcoMW+bOS7sL1A0uUlZmuqLMAjoCYN
Et6LOGEAGrrCgVEHbffB7nMSnq4AbvAIF2HDRfY4v+lJ7IGJyMUETO6AkOB6zZ3f5NSdmIIqUiJ/
AFPCzEccPAtkPOo/YhuhR3OwyPdKNU9m9QczLcyXRCtOJa6v9AbqafYlZyrR5vnPFGJfr5iyTyga
84vhiUoEJ0hRSFJFxA+f2PAZCztMyAxnXpb+0HF1FKldokBsW8OH4M8+oNqAULauto1Ae4uiDfiy
iiubSqPPZytsMZrSR5xJ+8myOI1qN2EYa2ZWL0SBXXb9rqJLGGeud5h4P7pMNEfnRmWrT2wzkXtR
W50ZPCRdzLGRVLmoR1VMlQxKMySPUQsyAuSgOXv4PmOcS4e6upDjoPPvprGNlquF76abGqS4Y+73
CP2yO5DbsJH2EmkcObeUnjx9S7kmyucbP2QZpFQbD+EsHPA/Rq8lAdHVt0v/5F9S2yuioJl3TJpj
6II0U7GlAxL1SXWBL4gyeCJpyNnY75GYOMrfBS2uS3rO8+EzVzyrdTQgvDxZ+paU69fXmAGR2PF9
03kNl9utdSBcraUIte7rM719ZjmEc3vMYnEnYNb9d81zd3sb19WBwERKnYAh0o8Piw+KfBHnBF7h
VZkEu3dCBqbfxtqZIZbxKYBiPNqEC2f+6vIi5PN+nQe2wGu8AP4O7ngMijs7D6QXjkIktHjhAK9e
d0EzF/SWRHDhGvv/p5/5BlmWQ14iftjwvUByCL4ZiRzP+bwgaqb3WrtlCx8mtoCTXLSg7hyGCtpN
FgdGwURgP32vHAfOfo8L+vVM21ItRvuT4s5r+35UXLF7mHnUuo31iRPziDkTsoDggS1SpwLfJOtT
5SRflA1ozsmK17J5Cm6KUUj8rOMFQXdBOcfr+PEFAG/AJ7uRC7JTjGvLp6ZHWB5UtjEGlFdhMdkv
6V/rsnAeVr3aKPtOBGhfqof6R5q7Ndp9N6hE2AZ81W1IRqvIsJLAd6nJG6eQn0kZ3+ZWvhktgSHG
kl3WrCuMaeeJqz5Ax8AudL73dZf3AOwlICaEcjEUnWPPJqf3zuWTVnLSD74ZFKbkzGFDkMLK9sVI
6mv53EKCwja0X2/yrtJYPGGxRSIonE7kyWUzHX5QSgDvgT9MGAUrBFQDmZJKZFh5HW9TsrhlvfAK
ZtHcuLK4T5V3kQ0h2JzzpHKKOWaf5UXGoaO5Pq2pQM0ujp8zHIPHLMo9k+ZPMNOTg3LrRh+sbhs1
LSJokrpfH6DXZUgSK4Mm57d+fk+0k7P8tKZALvWqPm63bbvrb2nbhqyUVUgKI43JJ6w1zHq1ZRgZ
nwGxnsA9iLWKX6sgoQO0Y5RCgAFaNi8sS1dvq/eV8ihJEqFA12pFs5pLrz96Av2avRV4pUMb6+9G
FrjUkhlGWLqJ/nXCoBIxKWpep0WNeSR4/T2mdtxt6i/nHrXK2XVGc0/gBTxy02p1iPQ7vQvSrR+K
5vJtUw1zujHtYNHAqGyQpmNVzmWU0kdLi+KGfkUeTfEO3oXAZQE3kNh7SYgWrBNoFLTou8ONOcRU
M3L4zLPBmWWgzQaYcETfD70hOOyKRXn8QfAiNoE/Ay9wPEKmLZRCo/JW2nRSN1FejRS0gfp7jCn2
Orl9u76TLdmwyAd4RZzTSlUNjfgHNUTZ1HEKxeY7sdBGarPgmrPgFrjq8oKXUS7H+FtD26+hqoAi
+DzgIeC4PJwrKDBHi/RSEyfq6w1ORsOqkgNhA0zIDYIJ/32f90fUfNvMSfYFT/Dy8/nmiSuPzNHU
ONgmuGBlATxsym8HcfEwMfcU5QrgoM6IKXUfVwwelDHNXHg++YgfNVCmeGd0FxGWqGhQDfydmH1D
e8kHvDYGIWKolo1isaOZsYs1VQDnLJ/68SbZGIH2Q7lhSE/V3bU/gw289hSrTQaKsa4xJ3MZCnVb
u5Kq30QeKe92DSr3CmVGQwLN6q0QZmGQYH05ZF9Ucix3mbnwcKtvrSM5o4UQf5fU+0Q4eiyAV+x0
Z8KKdLJ+bsmtYG5rxBaMBAURfnKS22wbhdJWZXy1z7ZzAX7IGMtH5CsN1dr1TVIdsqXDhkVxKige
57GGggLKTpFKsbToHKUXAvtYPjUbCRppLdSgy7U55ckmbXgi39jqesw01JZE1CHDBAgP+Up3ZWDU
RlSquZ1K6LcuHyhVKDM0/FsY8wrk/DC3mTRfxLvTnyHpia0RTW/zxUS3vkZ8dgIPr8HN2JELXwZb
51vDkA5F7QkhCrIrTVkUvtx+4UnvXbMOxaKiJYUOBs7ZjKPkoat4W2bxSSEQnMCnDKdztlzuYGE5
jGTOj8FEAftuQ2jq2Zxf3NjGKD52e4FmWhsxmVkf/FJpJLm8Q2mcLgoYfmSPJ2E1lbOVns3VVKwT
jZhUV64wFqpyoGTPwpvthrRaoPJYViX2KVNzUKKth7AHZbhszQnwpl4Bzs3Eco3GDo63LbFCXoyJ
D4IRj79rvxt/tcFjBgZgeXwOBZ+ISlBfsD9Wlw9Ccxd63X0Ru6ujf9uyjczBSnHKu0KGFtRztOOZ
NzPxpUvgbkgquFNcxJ2aOf9fVjjUsHITKuhB88oc2rXPUwWsC6OUbmNbHnbVTvr6xofYDoLbSLUd
Ta4IU5x5YwLVLVuBYVSYXzKEjbhSPwJX54byaZBGH5mZ7AaxYhUsWczPTTjHFVK3vI+LUANeeiAV
sr36/DeoedFtYr/hjRzkeMBguYyqvcCoyXadis+6QJKuqxTewcGG/3vCu2lUDEMcCTZH2KsZmlt5
oSen6Os1IoJrjLiZMze+wWqgb9ma6R9jXvevf2r0OJvCQxI5ZzKu+bVFbxFfKaxeYxsclNdH8jEt
DZZB9tC+A9ZIRFMxH5M6CBdUWYAPf+uYadrPXi2+07C+GCaGddUkvw67Dtp1/zps9v7QuQJB+WWg
jKYDfhDTtofTUpUlgIQUN4YTfua2XSVWKFXFNrXoirnNlEFREHFV45o7hb5cITWmL8drs9I24DsA
1vTHhRAG7JYhciOei0pcMPslGMqLmkYWK/rngaW7WCnIcE74RW7KItcKrsZlrmx0VdZnLCsrLwYw
FWR7JhRppVzW6auJZLM+wAHmjgBPKhdkyd3O46dXHAiFj5PcazdiR56BKF1n7lxArd0ShWvjZG4B
wCVU1VKaJe9xAGBBbQF8KfI5pfpY2mnZiSROLO3x0XjgCO9TEu0t+nkQjjjSQ+O/t0pIpL2yYz8O
q3UwCKxjX/HU+UDWntCdOBwnb5c26Y+s/XsV0+cEisbj8Ne3Wdynll4GK/QSpv6v0Up2cNv6Qov2
xVELuOoedVXPtKeyjECh/4xL+x5u+A6uT3LC83JOhRiD0PDI5E9s4xPByAq5ykmqbtg62Cc5twOP
fe2hqWQg2t4AkpR9z/bhSzLtDhUpw8CH5hZAYI90R/VI7GVg6mb1p+tR8vVwtGSY7oYavayca2Bz
lRqlV0JUZQ611zB9NrUEAgZg40YYcs10md3kwKuEL1W9gi8fvdj7Dei0lXFfsGQSGYX9AEzMnME2
Gp3r4L8enXzYYLbC7wzlD/wtL70L10n9Lt6BN5sQo3kAhGL+EnLr2exLvkVC0I3mcY3lcdyHu6fq
zx546ca7kxFM06suh8hlfn5cym+v1jQIit9NbDTdOtWoyC00ZpvbtwOK6IwgoqVOm1MblZ07ZrMP
9Y0xxpFi+cUGjPFNXH6E3paEP9de825QH++1aDiBxpT/TlLzfMjVwLUQ5E3+0U4jXD8XznNdNMAW
vrCEaKNOrpJtn6N4C9UNs+ce4S69gE/Z9bhY30P6TGwA/GzuimjixRrcvcKIISuJpgk9splHPdjr
v+Fmi4qj2TOX699KXlugDdkwWPIVEuDPg+JXU0njqcqdOGZ3+48Z7HL2Lx46yvi5wB+AQY+cDyLU
8RZFKwvqh/Vo+ERaq4bOAa8wHOcYL8bQ/jXaOjBYklH2413YguORYo/nDu+CMWwyXV0wS3wtQNSm
DONowQ0jC2Z1fi/TqR1wF6RdTfBrk9b1mEVhAcFDUxwOY8EbLSz+68HhvIEvOFZFhw2f7QiyI9Dn
INIE2uppZQwG5TRYr1w9tmqgvAMLokNTPZrySS4ahqJnwIQPezUZWhUFHNlhaGhuupP8FUhDax3F
ceZHvbMng1Moy4ja/3hcpkrpqLFTXOzMiFZhPjba+rHzmfmQXijCFTEjFbnOz7UZgERGJriXYlCa
dX6MHrb83bUfc542iPwcSM5v5eA7cbkZkir84X6H/n7GKi6KbUa3wAUiJDkGarVveCn87a/Yy6TD
kV4RN//4e7ic9NsAsvny5H727komoWLZJEOWv122q84oj4ytIXen8pixaFQag+Y1ecrw56fwlL1w
3lnOu5pvobvHPYJ3j+xiE5r+atmxLPc/TJ02Ljx2B9lQVN2XSDq3ZcSgzXxmWMije477eUy2rr1l
5ZqKRpPvD+Ap6kbF5+frfvJeooAp+NzY/G7YOmV/qQlG1tBNutIt9uQwsey2W8wl15KaXbjKtVBP
Nk7/uVTNf8nALGf2QhScfq2cIiJZN1QaJ0pUQ6hOT80vWmN65is2kyTLpNxRALfnWI3dKla5Zubo
ZwjUidceljon+Ejsau5CSEmn0JHaVyKUNHg/qQkutvXz+a0XT4L7pvDQYjugVsjIfRi5sWctlU3d
S+Buo9HTf9yXpHm+5j55xHa7dJdyFaQUkKtRdhaI72V4fDoqct36kjXvpK0maPWYZcG0AMVNF4OG
Ag4FCk204Sx91r7o2NvtkgY/nrWPZN5DDjt+tMxUf0UOBecTEaCN7Wzhko0qb+pf9/8qIb7bs1q5
f0PfKQBkmtazPGludmMMs60HP/cXiMjA4cDmkZXGAGEGMCstx+52vbyOl3umx3wWeWQsDJI6w33K
oZELiFT7QjAtyfQDNdPSe0rBxmg65YHjqhYy/84bWoHNJuFlpj+UiyYoP5zlNSUYgaM2OqodNUyR
VfyMoL69u+M5OkEIh2ss1wPjoX69CQT4g7zieKb99/MbwkqVbvk9MTL7sEUwKDRgRosEvuoTIAK9
I5ApcAYzJW/nx0tXcWve7zk2eenZ5Mczp9m9tQ1Cl93ls2wY9EX4OdIG2UeBHb/ZOEanmemG1jvG
+qn06apMDzYM4/uX1jnqyWT2YF6u8rIKhVZbGBnHUaPrTGdyxxaocLXkHvpFusad/3/AGXMPD7BI
2qfqt8wAHSVxRANSZec4H3s4YKm6LeERZPPJTAMN064SXmhVwPYOQ6q6qAzxl7giR5ZqP9R2pZ/z
SF8ldHFOv0vrkM7WHrnBnQc65XC5RjrDgkpdV5V47sfBaDCSfFBsWdUSBe3ajPeegUvlrK696B76
uscrjttYEe2hc37iR44O/bWVQB5rdzknD5EuDhe0dsK5mM/QMXaNgj6GWFVSm3/t54aeDMEppcnd
UCwthh2ssH+YRWFRCBu06jEZo5DIMgGVO75VuZNhzTIHhSnRyvbAq0Ni6AeO5LGD4JNLRjQ6m9NJ
kqEDNCySbJ/h5QMfJuxdC27IGahr5dj/1Te4ML3Za9ezSTLQRZCjYcvMQAuFuGbFJinz1qSrR5Vq
vGXihzVXe8PmCJ6FQXAvShTKEZXrvleKO9flnA==
`protect end_protected

