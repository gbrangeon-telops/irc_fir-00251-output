

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
qYvaWTl2dVn1UYauUm5HneGLdmTNfKYL2CALcG7YBWzuKWoXlk0Id+l1oLffyjtPstUkcnB5XMcQ
6NZs7JK9Og==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
QYtaB7bKNbwxVddRWt78CWZ0keZknIQG6IQKSIZ5COH+hNdpgy+tCPVsEHq4IVZzTG1P1o7hP4Vk
F8E4xV3B+P4d4XumR2TMQt1O3p//18K5GFLVc+tXegTNm7nDlHWB2EseJW3Comce24tPY9JdBxY3
PqZ0pdNcJu1q3elLkyk=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
dcPEPRyvFmW4PpA4iDmUUiTH0W6w8Tp3x24VnlLzTcuDsG/S9IG3GcyE78eNrT/x0pAgwHhrMrSY
yZo9WE5CUIc2230lFJdjwqsu1GfylgdJvImjNnSRTPzlw78/vxcWd8GQIKrHyFhACpS0FlCWX80u
ir6wyey6yythPFMR7YL9alngEab5jqlcDLLq05xFb5xa60ZtUm6H8H/kSZM2WCTQ/2EYo9aRaoyP
YNJgznw4M4JlCmjNGCsEEMbnrUH5XC2MOkUpPSJ6HpAPhZTjHtmrQy0MjGpBzDrrGJZmxlIzL7x1
7fFFHCW51Ue16QvPlxZlJr0kCC3nTtDv9f7xsw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
zhiiGh6iqBtYa8uvzkWpAts7vZ/x1/EV8yeLKnAXP52susoGuPOfmWMYojIG7BJlvNdJsqMcu4aO
YgpCERsfm5E2WNcFxUppU1uIOa+cnCBSZ6N5aebRGghJrQL1tUzWpRnQ2slMJ8Q+gRbsoc3N0qtc
A+A1dAH+z+hdTGoZBRY=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
lbE1QAVb48OwhlUCQuKav8khO5ghQAvoWa4EGI1wknY/PAoHSz/mN+mHHLZytFcumXquM7gAj5vW
FkPYXzAy7xSUZBC0WEUc0yo4Xa33jDRDxY7cxGlzHmyb1RsXl0duhVMcX5rDmM/+KiXLbAmtS7n6
pXv5Z5tj4x3AoNn90rxrYgdqN+pxQ1GZhPZPFZggV3JHWj2LJUr0U/7aGlgZSQCcdWV2V8ktlt4l
b9BA5BfHfgn1UuvjTl44uqXII+j7cWg72Zy7D/yYZ92M5Y7nPBoBrEiv0PrxnHLMrIv8+jN76TPm
TMiyhLNg8NAb1xNexvBsDmGJWQnxf5cukp8uDw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 60368)
`protect data_block
YEDQuTXkIKg+G0nE+AOxp06mCl2VZIj6JqxJQOnKUtYD5uVmDJRGzcpXdrfO7hRJTnLr/OAxsxTp
u5A2MZul7L2upTaXFoBsijiqPnKRBHPpi3DWrXgkUOk1VRk6nMPgs7+M9zV8gxk8drXUQdDvYtMB
GuNDInzLatzZKjUPV8oG+wNAIjd2d+HNNHL/5OuMl6U3DURSqw+T44+yiEkTzNpTd712W4f+pRgP
g8APcx2OV5XDI27MZv/vcdHjG1JMYycBns8jetSb6WsAK7TAwgos4oV3DLH2NzUXIGNHex/+V7W+
FZiFUT+YPKQYnj4HbsZlB3RpCIyBez3Ig6G/7TfJTVsWTSNyHUEkEe8a0qXLVhJFPZvGkyVL3zDT
WgiMX3SdELeSJcBLivGjdYJT7BnognhcJTN/JfKSE/4igDD/N1nRVQ/JFe++89aHwbkZmaPi0B8z
ACEeBBe1xz5YUSjv8lSBrNH8vf08oE8mxyVsPCyV1LTkTU2IOK+mBwKIFa3bLXGNoQPUyI2UhN1z
Xq4YT+fEzoF/Lo+HJPRV5Rc16QiRyWrAPQZWEbI0DxcttqEHcqCOV2MkM8TlKr04dW6wNTEVTaqV
6Zn4DGwktsaZ1Gi98QSi1JUTUZtU98D0s/uMW++0vQ5lscwMlsYXuCdBvGzTH6kMyMu4XQMD30y6
l++0hYsrzc8bb8OGgzKZol7de+HFk69NXBz48wLcTON99kxGIRHwAXFVIRDxUj/LgyOvgi5ml/5j
Uv+ega+MhhJGdjezZoSXJSp/cK9LGhWbN5U1jO118k8rqil+Cth06rgzOicqp9lGX5PETjbHOz+6
zpDssBBWvLFk8EQDAg0DyMEeljGZA8N0EVsxzxsRlSi9DbJzPlP5Vu4TxG1HHJ4b9fzhiwOS/PrA
xaDbYCFnOIQvJ5CZysQ1IYyWMu1RfRH8CSDGCN0lfmgYeGIZ0aDdIM7bb56HYGhdIfzVrsVbke17
Y3rOoxAflNuVM5t7eyoBO7sWshXA2ZMhTaHp6UXd197K5CDnhS8oNCfvT+3l9/O+guMQmIKaVLNv
Zm98tHhgvaO5X5l3/of6LujWlUYNTNEJ7FN2hyM0doHyBRv7r9xHzpgm5JhccmygzQ9hZKQnZMPW
6cKvS3rkWO1pTASNAmPTIkHECT7RVEalZ36YoaeDm3PF/3USnYJtO3FZDS53pk0NAqVpwj1XjGgt
P3iYjoNJjSee8tJf4PR0LMbd89ihtOVmYyvGbol5gLw0gcuj2gOyQEhAU46sBYW5EOtn61lqyIQ3
t2e5gTx6HYBS937ObVMWuSW5p/WsGkDB41krgA5dBpC7sjpj1TeV1/5J5Q4hY8mVsllI/J5QqW6b
FKWyFdMswc71hrt/2Q9Ify3T9kUz8LZg7+qY1g3Hc16uMkZ7D+EA2TUnEwpiCg66zClk32piOGjh
XJ5u0vrUkGy7DSXzRLUj0X5epLKhUqFiGKDTTL/kV1RKqf0DHqk8LBY7GFatHIRs24+d0MH2cbVm
NBS+tOf/DkoRQwHUliCV2OOn+XVBXQ5sA1uxqbkQg1tZyxEHWD1oiH3HBZLCFLbZnhscovwkwtdU
IXtgy8PCqekZJBrIO/iz2f2Z3JPTQVP9akrFUczchL3QJyXn2C/lyINw2SiD3/uL9oDnCX6BxhRV
8Py9sH6OzuKUEXfXX9Mvr9O75iRrZj3hz/2EqfVQoB70/ZY74iR2RvOZknAgjoiehck6x7O7yERd
GNFfHPcTguCg2xjUsvZ6MDf+HUBXU8WWUu7VkIbBprKea3Pb7P75rVcfVpfIcnXee7vohk2hYX9d
jDqS3JfPF+VAXeMlmk5+jNmcopJyjHry4hpn7q/QQjvio3IawotHONyoywrkhqmYFfRNMWJwCrPA
XsUfNAvjXeV9B4/9DFz4O032cMNlkL5aXNJQOriXUxtSuNMMs9z2STcypvwSxOaR/xRxFWwbJ36L
aqdtRhCvHTYeYbw9zciLcaYdP68qDZo/Wu4OyNC7oZhBEhOvd+sL/qGyGJwUjmtSDlGQ0qVGcADk
AdEpKNhBqS/njLzIOKfuXvzO4mgYkXnzU/zR3WHi/IyVWAkg+vLassXDWY0+2p5xrS7/5XZQmhMx
f1ruS5Bh8hs1gzjBXD+kkOcuET6lLT3VLnTSOO63dkMU1foaYLbbmRiFAl1IW9DdwgsNGm4hEYgF
uUMy/i/73m17PTmjiXzhdkQjaB5ChP9iTlsd8926dXsdXtg+VQCc7XGyc4V2k1Y3qx7Nl8ZQYNqo
Y713Yj8qr7FeddqH+7LIPkl9hC0Ut+tOQ6Qojz5BiBSIs82tHexQZKQCCnzIh7sOSeJnB1///+ZO
fWjk9ykgLdnGNGd1qBL49mdSlC3DKvOJwUGKxEzNdDFTdwOT9ghoW5y9FbxGUDPIWNIR+3bOcBEB
v7eNe5rIhWwHRSqcERi9U9y4TxiOntaOXtifYyH7mnBqxJo4BSISeFNpSDYDGU9NMHFk6VJUB9qj
Hs2tZI9muytMFB94fFzMxguPXR+EW1zxW7G3KTUheJHRqxiTY3bUJvOYvMIYOk8YsKPpM6Z6jBHM
4RQEDKIOzMg7GDraJpSXgG3r8Eip6du77eSIu7i8+qzbelfE+wjjUpwGhgV44emCLHevsY5y2u2K
9csPqC4EF5AXUlLJqCxXZTwIjm4eKHTLvJp0txsqLqZ4XEd7Da1PGYz+hWw/0oOoJUsODW+5S/i8
7ycuv3G6K23WYwIlrUDwMEoehii/xzlfw+nhTN+rNtwqq8mtT+Q/+a2HQCIbSJFjWGSuAneXMpTr
g38myT8uYDEy+2VSDSA0IQ6f+4ZUCMG+OE6O6CKyJWSDLZuPcWf7KF2zHJzu5EJVowGvyoLAqpKL
823OP+1Zyd4AbE8FCvTB918ae9mwEe0R5QafZJOn0sUboy70Y9a7p9poWLb1Jk9Sh1wW2iufjL+O
dhn65Z++fCez6Ij3fwK79KLCQqgaQFWErdwUKUuJfwHHO7Cx7yemJWtj51JmxHCLyom/xVJc2Pg0
RC/tMPLI2mxNNjH5/v7rJHVHqa7/m6YoQRyRDGek4A+33H4I95qMrmHzCP7Al/31wjsH2dZ3YRek
mPsat0XEChxJffuWfrzVvL1C4UWQG9d5BnD3rfv042nfUBbiNJCx50UHqP7s3i1g1fFPt9A4U9Si
kVLsE4SY5PxKYbcpbE0vi8RffCMHCPUXbdkoUvvw3CH8Gz4T4SDLeSer6jSd47NmhGQLPF2j8RU+
KUBRDv0unEt+k2Ft5FcuKEQ6XuA/RWUGH/fw3DbgGmWvkkmTDiim+biLSCvZH1yeP9JU3DfJeSyu
fFIkLZqA60JYi5vHVe6alEiqmtLJGKgsc8a4ohPo+aEMivTGMMT22cBru5NCYshIR4RzzLRRb38T
ZcTZ4BoJmvocD09QYvsSG17NsuSlTT0eWbT15lPvb4HEl/bfCDZx1PbjMIXI/EURP4b54tEcADF4
Vu9vNDnJ7Ox3b+ioA/G0AggzT1yRp3FkGE067aep/QcRYJvvZ/YRGkY2W6GBJ5GKph95bp/LPPTV
cPMg+YPDLi1E+3TqLHU7c69lUf0p6USKoIApvyZsgl/ZkqYvBbhIwGuLVif6wUbTxQ0WjkQpAGWY
JfbDgJ0drHxBQWlntOHnCD3uY0zlYFx7AIwuzKRBi9Oz8zjbxMtYTAmvGiFex4diP6HavvjR6g7/
BAYE55uYbkN6uWvaKfFIhEmv9bUeM9J9zgV9xQADFgVhGAzi7ynv3xf42WcggrpxkOfigOaXtOjk
BdY+susAmpcmAyFcCoGKY8WdUbS5aGtR0IxXb+kR24e9iUiwI13bs6xfY0T2dkjgLWz/ODYSchxC
9Xa5DXeRDwAZe939lGluzpsCNMCooy2nByAxA/uqAuZf1nsg0QjDpSPmX9qaq78zFxItpxnGsZgs
sQopIgZeY0IUNGzeEaZ1raErnR4G/30gaUPmSSf5chJKTFsg21xFR8GDwwNYjjU1fFz1dS6194Oi
G5ILEBPX9uMnvNvdAwP42Gq1BBnaGcpXQN0L7j1o7RCR2miJrmCrjRIHa4pJWOt0+1CtCQkNhzjy
Jyh4Ue5aly1+t0yqLFjD0Wr8KGMNwpPqwRuUhGS0wZiLPObasWXwkK2hlmwnPeLgR9vj9nOAhJRj
CievtDTSlgfOrs+C/hKZbPwtEOq8ff2E1JvgNIZ1i6cldx71xRzblQfl8YO12KL6m+JBDjW8ctRj
HingtXloed+icN17czzhOoObVM94LmciSW/w1XSVZuyS7j5PeLSHkVnT8ans4r/sQ90GcOztZdLF
Yqndd7Vx0fJOy+YEuktk7WK0mk/s0UvQTHqLqV79vs6TUr0DEjKSFJ0w8jM2D9+CjZVo91f1yPbt
6u+Q54BMkYLQ/s4HFYsPH1Gn30PR2yti7zRMGsnRkv9yDZw/0lrTIehHEhfPPHu5/Lx7PyqvKoMT
+KfpTzquICErwkEHYEtg62TWdEhVxHMqwg3YeQOsaUq+gessTMJcyxRKgidQHmhl4ohVs69QHtoD
w3TDgNt3bgCMsv+l7KMMQKU8LHk/Fpwm7YSM/R7GEmqGdnS66T71A98q/GCU7XvC5/ErKQcs6uDQ
xYl/nyj2qflxS8nOL9c3Sq6h6Vfb33rIR4NB43JJL408HnJ8ZyCb2z8NcT/CataV9tc43M5whlW7
dlEQEewZm7CDSmm5mzgN67UPLHc2jFZctFVxdOKCsmxdDGnUfGnL9/Z/OlVBAy7K3QfwLAmPSRyp
WpN/a8yZSdRQKTdnYkPNqqF5viGd8TJKaJoTI96OD0gWKxCh8pfcpa/rsT//krZ9mMN5HG7T5Kgn
mtFgmHKinRGJjk2o6jvQ6auiLXsdR2l6hx0cu1G8Bk5IX+XlR+lqsk0msx2M2V/EjJzPrVAbzesP
ZiVOB62gsQFfc8bOxgR7tGUHLabqwALMo7JaEKdnJA3FRm9iCMDz0L2haEHTPc3Qxvn2sheuJs1G
x5u/SIlfag/ve06iUw/Skubi/as+eAu2G+4hHO1ig1q6xVp4XyajYqnzZfm2+s57EgWHNzq1Af4Z
F01OFzOZfNKrSxmAj323nuAXnSmnHishmU/yzFRZ+etO8Dd8J5D1k7bY8TueoQkmIRHjXH1SQkTJ
V3vQ7tUabxHk6rDEjzbzEsKmg9U4PVst0fNM1YH06V/lIn1qVYw4YHo/tv+5GEtEipCJDq7YPIJY
sftPvKXG0x90uFcQ9XYjCUVqRJxJIYfOMcpLbG/f9G+97+nzRUbC8L+TJ/EOg/CSBZkMQg3p3qs9
h56z6a5OPceThfnqL/j8ZDHnj4Wx5dm2P3YeYsDOnOFEJ0+jOO23dSlXaxAZaVEudMThUbbeiLOn
amQdTut1DKE8HTlSXF8a8QB6rxgejQoV++aqnFsZ7T3QcSjGGjPPBxJa+QV36qVjWbOzf0/aXa8x
LMc4rrUM0BS1ZYL9bG3P0Dcu2uNUNaLEpWfWASaOIwyxaNi5TCN61sVB6A6ig7On2x1zEnio6FyS
ASCe4B7BWXgXz2VDhhlG96XxBsiuiE4Aq0m9ln+Xkz+OWCb7lrHBGM57Xk26ySuFZTFUhiV/lzhR
zGBUJUEANX+ggq8n3icr0LQvr1DOXCZKRskVCHFzjBLCYDJDg3rhz7Ua1QWUWZUaaX7Bcf31TF59
Ebvij9DQS+uQv4Hi55l0rMFPm+BB8XAdsi6MxUpA468bwhwWyb+2zusZ7bqID6nVHwF1CSYyLpR1
bicU8atnk1RL+PSFJxlucrjZhXhKNR+r9vpsUhx3iaeCqTWfEZuip/PCKrz721eXWpgdEt4E6d7R
1Vq0mnyTs4HXUzLBa5n/6jfWAnL78vSAiRx9ct8PiWCKhqRk7E3rFCV62b8sA3VrJX0yQNb7EZw7
/ttBzmz1Z4zMA5EGVQl/bD5YGiK6VT07lAa4cQKWLUe7omD31oqD2ELGkZwLFtOjGF8WUStAiezH
OVvShB20Dk4FrOnSSsmeJgZlf86aRsvm6G6KP8rae08HBeCwqz6UbYVu+CgneRvM0QNs3caViZxj
dGKoQQb6ZkseFLTlX+rQ9pCB6lIdR3sb4tFDTsvbI7NEsaLCcFGJqP165VS9uA0MY+KYReQMkORo
cHPdUJZWMKkcrNgZUrKTtmW/GsDuGBKE0Ih0lS1wBrX9li2qN1fj4DJ4T2JysGubTHp6MNXtSXI+
L8c2SnGZShzx7/dCWLmJE/uh9CzAFWefaxh81/oXlrwxI2UPHdBlrTYIp6acN+RkMaxHAuTejVYR
k+s2GdEUpp/VjsTJXRCYb0ao2DvypdB4kpH7EJD7xHbHdTl+GK/By5Evxwj4vZx3oVjMKWULFMpl
FJ8kUJPvHPM1GRy0vxLRBLVGXKhKvK+GLcOSjQxAN6+ayLVechK2rndsFX78nCr0r3gXSgJA7TO6
iNR+cOVhEgoBDbHUq/eBaeUqvrFv+BqanqCL7d+VW+3Vl3PDIum75ky9I+8wvVWlGVkt88VwQ8O3
hDjBfZNpm/9Cp+I8jshJQgDAbs9CU99NNwQ44nG9aHkgJYZQsGaNwh7vQqB90I7Cctsv/1AyLa5H
2G+YWD+kXxYgvp07Dh0ovcw3vARkqxSlAh48hZVGLFLkyZBNNJ5cWn1QBOsNbUgAoa2iD07Tg5Dc
VxwrG+o4QebL259jqGsyNsSZdS92MkT0+4W/DnM/GYbgc3+pHGeV/7pT3HpymlFwasUQvpezc/w6
ltW3Za2RD8M6huFO60uSAWQb3sgBKIfKQEVMeLAFM+LzFkpLu01s93q9b6jremx11b5G7vM1tLBk
e7DTBmoJK0i3rQ1n96BEZzOF3abGniqPt8jhKahwPQVggTc/T/Rf3L3p7nMm1rfduC9APyEddWsM
AYXPJDAjll76WGBjS/MlJWF7OX1z1SeQcbNJTHBCbMMGUT8k9wXi7JUAGvgt5VPkOUcm1bYaKZ+3
6S2ZdznObHiQc2esOTLVpGOLizyE1PRH1MgTwf3PNH54tsbDjAoN84xtpiXmTlYFuBh1jss9YY1T
vx2QcZsXJOfGHk1zIpLXb7N9vAwjAbZOqUTFbgqIIbUftK573XxqEzetSZvleOAF0SKujducGrRX
WXS7aj3lkOKyXRvlPywdzRvn6Qf/8w2VkWiPatjHqvMICpNPRNQ4O0s5LpzLZudu6/JimPxBAXEG
JWW/h0kWczVXbIzRMYqgu27EBqkV/tZeKBPi+HTQ8t5ru1rXWSeHPziw7JUjy4ix6ZoM0Xisur+w
xzbPvV2FenfLXK4Jr3Skszu24SGComkpKaY+jKUHvjYuUa1rXShrdlrCjiXYc1fAAm4C0z/Ce2oZ
v2QJdRRJ7eV56VNvHC5+/DdrkEQc7/SiMZJYInCc4L7Pdj2rXKvh7FbTRt7uSL3RwQhuM2L2z654
T74gcTxw7BfxncfVrp+rZ4lP+hLlCPyyhVaQye/Ot8WPmUErRtDapVjb0XRRTkU4mrYwGAo0b5s1
Go1aBxnnqRKg4C5QKJdZWtimdaBu8ieH2uaBUwvUYMvM676nN+uoEHod3d5tAj+CBw5YE1TIxd68
UY2ux2ZHhX9QABKXCyx7ZLjxYAxAbtQXwbDdnhEY+xXoQhzV/H6loPS0rcu/2RucrUgsjZs/KTC3
4AXoz95xF0necoJUW1aGEp7LhJkFA3VkXjKz953WB8RYVQE7sBxvBv7hviQ8UDt7+3wSs6KH1LlC
9CQ5yrtOJY7IKLqNCbHgGxLNKaA93sTbv61qPkhGHY2CKqbFBwB71JYCvgnhzRpbhdxV26LJEEll
IerHWf4IoGQ8wp9XwEJC2XlCO4y6QV7Iwspfr7ZZF965tuZ8fqsRdBTZP1OXB0smOuTD0T2guiNz
3ASYHajnJqtFOxpU8zg9mhfQFD3DDfZqaS8mBuV1IQ5MkckFhpemAQH77u1/1RopZo/To5h6jtWv
QB1iomPKyanOSjPPbn8scpY/iXDoRRt7+E4OCAYriH1v09qn/BBDaGs8Kn+0UE6DxDszdSu4UJEX
gmGz2mzhnFgP+r5UFf7l/VWrolc7vOtsbscj39ZgM4AkQQ8FWd7CoEi+quLL+QWXhiHbMUD2xxMk
7KV9iPndJUXn1/E3Um2RYWniWXG4XAWuxvwCwjpeMvR4RFBkwJv0tdz6rOaIz0+9Coi/FYWlDqtu
mFlZbog6sj9V5TwbvmWAKamCrLANw3w3OUV+H+vo42YjIsgWpgkQ4c+aIsYrRa3XGwLtOgpzFQ7c
UCsqdrk+hl1GL9QEDg0sY3IswCCTO8m/YfV6b6aL2OJUBgrWUj8CPZI/ABvOWjpbrpHw24jUzCK0
GazAvNhzFFxdWiptiqullfd2ajxFdlqIw2pG9bGEqdGDt5HNr/R7xlTq12Vt0AOVkCKYuT2yIsXC
mXbVhinlt7ekaY6jbySfkh8MLtb9X7UTijbFNYaVky2T8NP5nF/e9ufH6/xWfGQDdrUKBkm3OVQX
vA7oDmRwYIsXKajZEGAgNKzje5ZUDKlGXviJ5ddluAVATbi5ofUjoHOIXpfBNFQMV/cickM8XDGA
JqqvfxyGxJCiSyOfqgVkhNjQWIgWVtsk4XNULRlWN+akzMK+fTlY2dLOq5erzG6k2L1VasbAcid3
Rh/y7e4gWLo/DuT37a/UclPkWhETMxFhbsaNO7Hv+V80qJZHh7b+L6dAclonx38qYt568htd4Ta/
ly3OruBmAU7vAZV5jVDeaj0FX9xBUOTLigEYdAQHUdg/A98r/jOyhgt8/G94BY0tFs2X6ZqoKIpO
Bc/992AFGcSo1Rh2E4D1VXypIB7lr7l8vjPDcxdIv6KwJZDyzhFUXnS7W0qd1++B9FK/bxtRWwYq
t7xXNkx0Xme7HEfRt65Vuc1aeRyZwzmHiW1Zib7Br4/k41cKfrJH0JyhPcLjtfYypc8GLfSMXjkW
RPHc7vLTCQhrE9SjD7Ov5NlwkLKkTxvW7bzw/yeSmLDGE/2mSm1lzxVJQfEG58PUPw8R3VfL4TmH
IBOPm5ThcSqAGNxH3sSG9nby6/ArJxErDblrfLKvGjHrAvgUU9qlT49ZRu3Y8NxdJzMIc3pYb61J
BJp9ukcGkNrFuyo4OZ5m3amvdJSbx4WhyXQDDSVK90AhTFXHlZ2fbstlIkncI82a0hRszebzqerk
HoFO/oXXBDWbNBD2k6krBH0vZtJL+BNt269NBI7wMB6HbmelqmHsheth2EKJzrHtk0lXuNnqkbKi
R+KVvz/R1DfdiiJVBIKkJrQXyAMiLgWVH6oWIvksPaBI5P6pj44doDxqBjRADkg/nNpMCyx47OSO
T9g+aG4dQ9pAq9JSdbSREbitaSg/z/7vUEvpspDbagz70Quzv/qTjd2+VOE8Y+4NTCtkiOvIAXAb
h/z1mkxDgohmayMs91T5sgvWpp0UBWM3K1A93BEerU+rpQmsbXuOFvgnuPBTma7iWs9kd2161aef
kJW1ZFsMi1eqZsh/BkuIwda7HFj7iRQ4kKw75P4oio8oncV1wqwAHPqL3hJ4A2h1MYaO3hAsJO0s
kEjlOEoxhoQoe97VCQpBQIh4ld/e0IJizEPveo+KkTjBuG95a+6AxafZo5GqaGtsmLxMqtt2x+AD
0Esza1crLnB8CA9ZCx1ZKSk1QfW+oV0h29coL3FFGReYoLKQZJYJ9yMR3EkYc15GXcJSwJpPES7d
YsWwQPEAYfuvBPg0+HFuZeiYcP+5GvMJ1XRZesP3RMGnbuGi3KJU4/REegSYWvki+j8vu8dx/Sy9
hTjtTnEu5vpGd/iCA6+JUDHu1sbQyD2QHTiop+W+NvvX4mF0zjZVSC2/zsoHZLXSBZDfwYYjDjGf
/kz3DK6U8KyeHq3hjDv3stbBW2q9fM+7SX/1GcZ15noryMhJAnQag88hqTJaogEPIhva18lnhT2D
cnMgaOvVPWC/k4IlH+z/1KlWCQnYMSo8hHsEkZCS1MXSJGfhCfnk+sKSBqCatGFN/lJn/49tz+rS
KtciSbo2AUgQLnWB0abCHpdGWdkQg+ieKStvZS7C875UYkicGaurUPcwvIaJGSoxBbnDqys5ROkK
bWjaLBa7/4RP4UuGHU5K/u7IoFYXEdiJn8tFGH2pL1xpwyu/oxw66HPLNRqT1wKuAfAD4hk2XHzi
B0PlBasPdiKpCVWovbXZPvKupfIA4htZ7CgBsGMBmZ/ZAZcs5PC7a+tfBtMK9xVvpK7x3BTrQAMp
dc8WCqRNRfFCRmCsXX37qQpxHqlCvxTLBqOpNP0uuhz6DbaoJZU9NfDueCkn0KFrlKz5E372lrOL
e3sS4eThjaBdjpbxgJtqo5j3kkakBfS82F9mk7Tshl2NbvQfIFuTlPsM5gceaw4HPMLRkuSsxJOV
OtlFbeczKJXZCxQT33ihHOXWUfkFKFofTcka4kccQAfKICCPpn/U6PUDlSm3KIRa9P5pHPStFLUF
9etzxTkRkyIptAHuM0ehlvBXisM1TU4m1j5HIicB24NOJa9DrK2xqfrMrkhyyCNMQBKgUBrlsdRi
US9UdC4ry/hBks6cIcS6WQwJO0jygmzpMpg//cNpQ1+/ByEE75ZgQ2jlyV8XUT9H3esMEmpkDATR
b3glKsB6DZSl+MoBIKGw2vL5udAuUjG9RJxoSJ+nGhCLh+XX0QT5qCSLdl6QmpTtUTsT65egykvP
1cOuVsd5c8BGYGTtUeuzJrW0qJ1+1zFzx+HahSCFOEbJ0pQXEYXPRkC1P4q9tKojrH0tWLcdvd27
knS6rmh47ySMTZ7SoOH2azDQTxT8ACBI/S0nSzWxKkZ8tPA2AN9Wt1meICc3dAz7HiBlvIVQaLUV
HLEbfxld3X7QFpTUqIFjC5O7AfDOuM1bNHCDBctF+prd59ilHtcwKWEDXtl91lsAXHrduElokY3v
BtnakkTycD3nodsBDH9y7lVaWqLE2wuEqX0duU8Bs+rtCZlw9Y18sUtWXV01rFlFXMTYylfNr/7g
SC/B3fMLvYFRgpjB0+40LWUI9mgKYl2PaQsBd61PCBjNkFg2GWZQn7SedszkCuBuCpojZnOmaVjt
COAtp8KI6I3tIpnndeVKEWlbkdqc/YL8K7UI9wTCpTQxBMPh8AjhY6n7r0QMNt7t5MmIvacG0f8W
ett9xPRGrNOiBBdXQvVlaD/HiAFqlrWpUKGVzNsL8XTf24kLHH/RonKwqocq+WvXuH8MsvKou2wA
VaaKqCQPrm122tQMlwrTHxYwdm7WAaNqMyieJaGIpSOv3JOqqPGmpFl7M7K+Ny1br2PPCV8Gfoov
Kv81vqVl6RJHULEE+9sCOQ8jAkdZq8srPcYoZt9e8X+q9tv5pblc8TmAHksvAb1FknTZtyIeS1Wd
0rgbQxkSIomDEQMHFypCjPbMsNGI34OY2dw46BgY2CXeCAJCuAA3w2nKtlRkFuv8Eu/b5CU1LzNs
oPrcYgrvMaN9wRH4eijHx/DAFk5Rt/psTGAG8SaD/HJDH1lLksseCmT2WRoX5JIyZNJxC8+QjWsa
2UxuIvT70cpmy8yEL63PFw6NBplx+ct9nNgi1+22L1qBRSYa5pR9xPoeZDlJBmb2h3ZKxVjbLtTb
VQYgfA47ouZ12n575GlkUpurDawa0mXHwjLJGqDJ/bkMTWrKZlvFhHEf+Cbzv5kZse8HNBzXjV2f
eebPYIVNks58g60qaa053frXZPNtQXICKz3O94ltwyFYPiF5srWIom63dsf8yTPBT+P2lsWcmR6E
/Bxgr2VF9dmn3Qu3p3ascrf3lqkI6BNrYxNYX9CKMSmSPrTJpx/rksfOaSiJQ50IjhMAT4I4PeCO
3fn4NX483GBIloBcV8mgdem3wMizx4OMcgsAK9H/J3qgGJxFEM/JJHEhqi6ONzaU6q3x8Zv+jld+
DivmmWYxuEkQNvCqW1IMFltguLktDRmWna+wieF0q1iAsqjlnbX575h8PwoYq9HCzOXWHZNDCasN
asJXK7Dz8iTVT+Z+EFmcc7rf+ImaGUQHsVul5LXfU9cwcYwl4MYhLv5D0KRKj7lYr50SdBBJC/69
G5JwdXrUBkXjhJlMeJ3Vw1VRRW6SH674tzYfBQg98/obbRUge4o6lKZjLcoALZdKSozP5R+CYSW1
qToiC7d7ofRgiNUoAnsQoE6MLhLxnaZaQWL3lPy6ePhe3WQnK3AC+CmwVVahXCY1HJlkc0EaWR4A
9xmmI1H9NuvDCB05YidiLFqYT/QvM/qPaMseC61HHHw3Qm+e3diO28ZBOWVAaPIKtSdIvVFV9fNc
WLvzYkSyJHQbmcxVob4mGNIgKcvxvte5nC9rvQZnrjWlq0bQZLil4WcX8vE8mLVEvYcZKopnLKTT
6m0ed+rdQO0Z+/tzLq0WYwpFpILmJQyoWCMxDrZWxlYwHpZhD3yyvAkuO1Nxs93lVPg4vTggI2yP
O03LlkXUIRINeCLoPXiEVpIwNKA9O3/szCHMemtWT9sKGue7P5Uz7s6X8SZQ4uxVS9VOm2xwgnlP
tivY4IgANsL1hDsnrHufZ6yCgVfzxvf/ZOq2IAkBz9IAItM7g5tmzguPQ0fzQWEO6ugLnDFMnjTn
lJKwHRVLPUqDHB5jyUQXX7X2VSo5rgyp2GcirUwyxyhOueNSA72o5sZgPHNYViHdU15BXnVadw0R
jWylo4i7z4eb25UmURxAWJwCMwnTRRsMnjal4/Mbi//Lp2GwvFY6r4JTHbXq5XkCuc+2XzKJ29UT
pbpBBRyrR0F3N38csVwdrcFQp0mrlvBaG3kGYIeoojcxHhtbr1gdxup/wwGSAMCVOYGEE88MnbhO
hCSfEPhA1iwX1KeTxR5ZF2jBer/R00Fe9JPDmFk3kL9fIWxjlvMSy+rSr26CieePQKWeV/5r9bXC
Wg89NXOXrj0BA0ODRCnh3o495et4dmq/7FsdYyH1n5N7sr43Km7sH2TP5x7EKtfOS6FPyiltJ4t8
hxX5Rr6kXq8wqajKBs0R/XxHj/Du1zE+YbvklOA1zX1GpSGIEPm3r1Uxo8wXuqKM6SLwZlA4Su+W
bND7/PtkMjbjAQ2mIfw+a3ZOrayfz9/a8tFW2tuqMUc+V0dkpbB2xW18WGYnS9N1uJ4hVvXoOgSX
Wkyi0h40r6ohCjubr/ZxAjGr6Mpu6vMA881mRGhIawk+inXNkWWqNXX0vcNzQj2VaUlXc9hoWOUb
L//5TOsR8QtybbY0Dm9jFqdUHKMeLHZhcvIcg3vlY+pNESkcQOFJ8fHEELzD8JyL8W5C/IhorYYk
xz4bFq/kcLvsT7O/2rmei8PdG9tryYndtHqxL3OFgM58FIx/MkEHg/ulgb2tHtIzvpRnc8KS0WDv
+JJoFp0BpsFWj1c0G4ZzHB54Om9KYz8K+40OgVT7dtxjrAoAfbS0iteM/bF6MdNZt6XxL9Iht8yb
oj/kCwlCg/V2aACcqF395T+2gm4y38TKFb93FCipv1E7u2k5pumns5VltQ+r1V6/M6B45OKfxora
v1jz2ivgYuaG6cdrX74FJw4oMbNOGRqfOWp523Recro/aWEgO2/Q5oxNOEWDgV/4cj6c25fnzDzc
guTp+4a8+Gux/WHVOdH++MIKQKKeYFLXwsXnXoAqTKOn+neXsWDp2Pbne6r61QbLwe9aD9mHOApa
RIZCd3Jv1vzg2BPXcyrJH8Q4JficOExAE4MViGQnT7Pb0KfJfToCtW0L7bYV1XP9uEY5UMMItbmF
/OH25ur+5hkQbZmWEfmYHiDhNlCgbTaauq2ERjG8Pzvm1dTnjL5Hef5OikOV779Cdz7oY4XE83s7
Iidq3zuyKNe5NxRBZrBjsf7qhyVDVlam1w3W8t/D2u9bYaSd8pb+cJ7I5C6wwmfMdgXZkhOFWKv8
zO80bxyFepqUyLYq0TsMwcFwQgBEt6UEYG0XVpQ9IXKMMhgTcQwiQov5qdtjSTcVjSOc9+W4rSa0
VoXS4u29U3sU4YPuZralysPtMLBotrd174e8ExvaZMF7zYFSS8Y5lntkHJlfqZFnliMcS8LT3qUk
nnZNQ8uK70XOJVEDnfHxahv45lDb5Udlw8mKa/F076y30bO/yONPUJnb7vXm2ZhUNUkW6qu23WzQ
v11XdkNZGtyIhBaH+0wX7oiFJnIbAGikepph+8Z+o4bSgm3iXeLpHctL3Px3vDDRGZz7iFETEtqn
rejaJrvSB70uhv3kk+4Of7xZa6QPrr/WsclnNRX6Xkr2B7ydVqp8H6pNH5ZeOkgLhaXhGLDCUEjS
TAnMIBKdx+uD1pUVv5L0i8TvYYu9fJRTwOupnBXJu8UGXNWaaLCpKm1qTdEmxCSrsOk8SEIrOK/N
ZdqxBZCfIRIN2jCL56Q3zVhq5a5fHUd6xhNIQB1YFoe6PYmNs9s8Bu8Jzx+pJXOOLtPZ87DCqDYV
zI3QSdCVh+HWKePKOz1Yd0iW3cMjekXKAtchm60ujhQV941F4hRHkZlDxS+jXzDtaRCxUePufkk+
yPwgzqCGOPP7baiH6SH9YBbreoFWN5AfbCOJMBxfRLPfdGOHZoCuY0oLYWvgU/JrmxopDeY6+EIH
0J6kaBygqU/WAz1UVmZklAuVqxqXN0lD5fFcCdK1XOwqAtm4egzxSRbHiYmF92N24TLke4hwViIi
gHIb8m2Pj2ECn3WiQPkMhFGokEQ1UEywEYkwWxz13Vp2cnDvwC8XjtL1qfrhWAI1j3qgaONtHj7n
whVEiLng/qYLb1BrSOB/DWDDkvxEoyYx3kuPmqd4GkH+XjmUZ4yYcObtceJpV57Z3fUSl55aeXM6
zgUfhrAzkeVyFIbVnsECOmkys6LjXOBnBxZUEQJybeXlbMrI2I6UxHXBxTsYF77C+Kz+x7e/EJHx
LLk8ytXrHqeni+jNWbLBIuo40y8t8ODHCj4mbvmFb2EzN6zohGBcGCWJtOnnRWLJWbB4HkUMJmuD
jMxw6BcnyJnS0yQHrrLxEuqrkpcQcS1+qnFYUnyRs9hZ5k2ncNFxvExWbvmtAm9Vdr91qiy2UCPt
ZybH1/3k6kj3lrHcEnoVzSKJKa/Jrl2jetsUxUIcpEd1kd6NexMhLoGL7wwnSxgoZpA/Xx0v42NS
YRXv7cX0qRqkY8zGu46ViPf8rmioMFF93veem3i463rQRD/8ENMP3tsMIeU+dZtZ8X6A1loDVG1P
NuMtuB0PzwCi2xn17X0ICPN13jWPYqpayyvDZ8YXXpN1p05YRnvggDh8sswRgpNB3VvmJ5lGrPR+
AaS6w0koTg3aJYHHGAP15GWgYbZRX0XzXk8labjWto0BsOs5sHOBypjZQPJNNPFrWS79SWAgRoFm
sm76awtbvomDTFOmC5HKpkbjfQ0vyL2/vxpRVBl6fldNH3BJ6tZwyTqvzzNIj/GRpLTu+C/P/lv/
+Fp2VUv0UccISTa7NaLMRnEnFNYO6eVcuCCrj4W3LsDv3Exdp3a7uoueGsqowzhlopP1llJakC4R
pWwIP4VWQLxMrtXEI/lgsJ/GD/ERrfcDIDHd6iZCCySSiPmlK7CESVRM8eCaJ2VUhrM4HlNFVsM4
pqOjPvEAu81M0SKJ+BPcVGkGpp1oxiNMh9/QYSEeQAWpgrLjXLk1UNFOiMVshaSgzUVV8so3qXzR
Up1FhrcagifsTRStcKUOKuj9Cx0HFXNcLJdRmKuZjuLqufEWN/D92rJ2heR+rfu3zivqeqORQ5ea
KfGgW6i6toFFQJHo+/R4Z7fj7jvjaNVurIZqZ5mad6eNjcjwoYZ4bQTA9jq5olOpCyUkeYxz0Iv0
5968Y+/Vsjz0qJrWV/c8Sc9JlhNBcj8QVfCw0XVHUT/vErPMboZJx3e7EqytWt0ia/+POqEX2gbU
J1fzAbIID/bRV5T2iCI+Zij+/vNqpz408ybxWM2iT70foDnkqKHJFLqmj2oQadQnex0bJ6V4P+te
rTxa6u9Yk75dptoksBgTu4smn8FJW0nwGZ26NKmjvtSusqfN5n04QIA97vaXeldmrG2SWohUHEyA
1TXLVcQqBlsGw8pfsKWNQZZV7Gl8gvKoKSqCuB/b5C+JL8h697p8Ie8xCXTFX+cU4Q9Qm3gkjyiZ
ICww+movf/V8Z3F6bStt17ZsPMKKbG19TkZPyL7tRdqcr4lHqBt/S0+LImFvYkT2tpZee8AEzFam
+3Iu93iDAXiSdlaD54JOM5fLSTbMMMgGurdLKVlLxI3oqAp/DnPbH1HOjEDox+StNn3N7Ij6dOlN
fxPnnjNpRs7rfZiTrmRlEz3huIRu4KZdZBn4hULmbwJBK8+R5Qd/D/xYG/UnHasBkzhmdzSkefb9
6A+mmZaiUZKb8yBnH6GzbRmOlBjrLXo2w/QJr7ja08ErSLLdeFV72r1Z9+duZz+Xhf3uBpXo7mSm
DDN9TzlGkdvu15BftbhuO+tW67V/Q0fSCtWqRBmeBJoOpJDq1o4c+HZbrc7Xt3ygRcrhOcXlK0Wj
/ucAMWmurol4vNssJw6nCKyroLIfrt63vFwH7eC/ivNZ2E5CPY+MEFbjNPD8R6Usk8H4XHjDqgYK
kEn41X949cMbjd5wwF0mbthX57fkb1qgZn2qSPLry4CxTkbz3wl6xW8I3vMzEqxsSvB/KgFS9MFt
4Dx7ZHKix7Mf2ddV7vRMpbWOR3dCfSXpmiEeweDZOsC2CVLFgooTu1sT8dBXf4dDgvpKkEJ3IxyQ
lJ6IPHH3cL+b8CIDN3bkC1GalOw2T1svJq1gOZ23pAX/sU4GGHXeQz0wmSQGvCTvkGeesqu/F6U9
ZAHzTbeRTOnFrMD24buPPyGpiP0SrBJdAJSehu19ZHaIVWwBMx89fCkBUYJppeYcszWACNvehyoR
EvSyhW4/jUBvxtkpghYPO8BgX3UDMU9P5aJkSx+D6z7NWe479PVn5J3q2rIRV1JpfW9ezkQTDPyx
aJVgroH09PTOglRO+586wvRALEUfLPNo8uLMkowDlLpZMU/+UjtXA8K9uNvppIlfGeWGRb7npyEo
bnV8o0Y7X3nSUgZcUWwNe+zdsM5ucov7U1T5VUn5jbsQOcZCVqimKsz1Giv+z+mPMh1J3zSSM1D9
w+xng6zaU5ac1A3+nn4Ppu69XkZu9qR4kUe56YTDyAX7psTuWmLQj/vuRP2gs4cocktz9mHp9JcF
9VchKbbzRNBje3S6W3aCdPrdQ0NtWBAVhqGSE3CsdqPUwzmYdlYiZfBfMx1h0HzbyShrWpJ9WrPt
tmU0mdbYIQ4Rs8iIK+Fw75nZG0nm4ZzAMuFjbaNlvI8z5jD+L7D+jCnJS0EnqTvalyUM1HTp1vTx
IBYBoEzGBBrUCRVWPmO3mXWcC2Q/NWnjDp3ANErZdUjqE1y7LdGYvKTQxu+DTSDQPxgk846Ik3wV
GFMmomrWv57AW7ELqTPNitMf1X4gElfepsCdtVEcqGDnQjRo8UGir08rxKhRzKMvUD0Isz7Do75r
IdWGkcmueAYzMaO8ku3zi9MRDOsDk3AKbbaMJ5b2H2q5UJTApc8syzqTuOLSM2g5M7z2+yRka2at
E2D9NJBU7kdPlEnjaF0jT4dnAt4BIs7R3oN8YVYTsLW2WoBg4xQJd0dLsN1R+XUBCCSO2/VFd+2M
orTfyeLPybwoIKJP55pNMQvPUiZch75LxQ5JV6N3xlOu2SsmxLprMjLBesYi/sk5GRH6rsOPG685
fB2o7g+qjCv0oxsK0cGtA7qsAIGJFY/bsoTAOL5Cf9mm3eRx/2ody1F0MXYd/2J//9WN69pDkxvk
vqGc5hYE3JeXkP1y+ndEwGpUi7vcjE9WA9LvCWBtOc41457W0SbP/g7LyQDwPsdYy1lXUcAJWEIX
T9oR3YdgQsybk4nrmuKci2rARYU7nGo5oXJ8CS81iRCxFFVa3pdLtqX1YGTmnmmjMn0QcWZ9K0He
YDJAx5x6pr1MNGvRvD0ABirktqD4tBKGM5g4AlhfYBDzYSiN5vipgXX3+UK94JGyWQjiaV1aXMn1
t7rgF8Kklkpbfc597eBh4HIPx5RR3qvO/HXx24UQJhtG2AyFBEhufUf6okeE58mdtSHiso9boaQM
XWyRM8gur+yY4M3R87nYgcyRLXSfr8vY8hHpiG6aimG/6DNEpbyNfi8NET1DZ2hd0a/6cHCNOC0H
s16ld/35dtkTCBfSsEWdV855eGb8rCYRQkgBQFBb2kV9bZVjQPTXCX/tTrHi0K2yj/eodWeSbxF6
ZQJGwPmmaijhEhmXqPcfaQietLR6GEPSpcDzuesuJlWpwiN2Xkji/15LNUcwwrclgcl3hSKvrItL
Vvrq5G37OzPR+yaT51kilQTvpG1BbaiLmP63KsLspUPlhokZ5mLDF2K5SI8/SfasfkLN/UE6387G
irHyQXSmFXZnGVUHZ59VpawruB8/GIelk9+3zZttozSpS/JCwg+dIT2RIHWhxa5IOz8mvXFUNOmY
/6N/5wIbIlFbwELb9L8cMbMUO3t9VV2Pz7mb7EvzrYrvwsb/NyWES7eFKcrQampPctr7A3sFm3cF
I1KtRN3roxTZ6rtbFNV2EXd08QmKFDGAgWoDum9+3n6KV4NmYJbmlQAO9ZIZIYB1SCZY/RsvLcrV
6mcbWvyD+bH5Jnr/7ZxrxSua259qpX5IQZwPHDPP5DzKyXTbPnSSid1AS4hFlN3lOjRhwWkWXVcY
HlrMzIqVBvtPq0sczHHUs5reaIppX+wArup9sHfOMLfmJ+aCEKnbE6cvV+co4g0czz5RWnwuPFE2
q2A6C+VXvEKiACENOqc5WPmZ3dLJJJmPfuEd9Wkl8eNBNsobsxbMymc0w99XIPP306z59CUEsWkd
lplFRUacZvUx2xBPwZ9243ukJ3vrsC+A8g3zbd5/MCQYFgEPuljq0lkaK0cap2fkf+w25pTYzD2w
TPxWOPUZLiL+wtzRnNZE3uAkgVlIA/cyJcHTmDX4y5DZZ2oabMOPn/r6CUFgH2YkJzSkdIXl2t/j
lVjD4Mlx2TR56/Gr9avSvv6TbTIJfJlXhrKKidv0Qt+fdRwEnj8Z4NWgfJAnxTch6mrvpBjdtJsn
ymsgB0zAHyLtm6SvNZXEfXauz04e2wGHA29QPt4I3V24Ou/Vkf1VLDZPIN3jm13wq5SFsmMojElL
R0aw4TxHrrNXN5YRMEDPbQUDmf+MfrraqB9aeyACo73eAtMO18aEKfOWfYin4qQijSnT3UxDZnSl
mkl9G2tsmVdBEfIFpTnws8Vd5YdAn5zwl3QPgXUa7Yrwbt+l/ytAhWnUYGT4CWyCZ/0Y3ii1U4Id
HiA3vGVawBMRH6D/DPYDi/wMy1nFqbm0+iXeWT9kpK01sk8FU+AvuhwRPvkqPmqCp3ztc7bCJVyK
j1qUNsMwn6nFb88M1VWGuuea43dRr6J5EHnCIsMdVHU28DFH336PkdmQiuecUOVkoL8HBRe/PFbQ
6ImTFWaV71I5XRpVoGhLxlcCWqr4pNQzvjulvsLBADIhfa6YCrxMw0WnEfptRuKL6suxUD5lzF9M
R55JiVgKZ69MI1wuBxnpYoYH/Qgh04jmI1wYKtmq7CrUm/FrXnxJnwYOmL44mZHtKJU7s4ZoxPvS
zyJMgP8sfUgYXvzt+QT7oPFXY80iyPGhiQDkLT+nSIAFTJbXiRMjC5dfu6LlGlV8rnkvHRxmdjxp
RlRJGzIT/9rkJmL8L5t7DQvRaHB2GG9Z6FSEgoB9jHuspy5c+00PWZRZXbyVfg++sObbPxuxoO9y
aVRzZkKvEMK4bb+LEeT1oEg8Gb8SPU9rl2/4xIq43duVSo1dpFDqQ3a1bfjutL8ktdFcLBAF1WdG
e/H0600v1x2fDTgvmXTnXfmQ2lHYf7CUni51/0mNRCnIYU6dOmpHzKRcVsmgRP6J6jsfMpfHFu0a
mW1BRjMFFEtyzOFtAYGLQ6U8UxIBH3gBBjQEMyMU/emn+lY+RAILbOAySJPUZ1qqcGKPm6z0avSJ
ymr8AOn8CkGm7UC6woixHrKk4eExNqrZ20JCCEmFGNL2fMRWz7W4PIarCpIeQXQ5JISeydFQTUka
BO7Z9BOadS/dVbuH/16EV4tc+UrMXdluIJmUJ3EfAA7Oh5tYeEdvCKSbKBsu/eEvMmtyqpOjF3TM
6s1A9XJ8+mIe5c+aN0+8rW9WmxcynyeVjHnpx++XpeKuwf9Hq1uYoP2wS6AlnroI5BWLsK1u+zFa
FJoXtS19fKIWX1lOMX9ITCceKG+9CnSdtVHp4NREmpx2U9PJ55jsOThbPWXUqQ3TW8Rj5vt83O+K
5bwyYvYb90suCZneQvHmwbQooAZM5vCHgGBuUELf6APIOXmNxIgdWIRc86UUzlu3RWH68bcNQdpj
P42EKjkNfw9D8+hf9eV6VZTYQdXTE8EBrAMPtFoHdHQz1KDAef6y/02pXoYBIGIyt7O5V+YntV2Z
UTubhzn1J7WdzLudM9QWS64JnSTqu0GJjkOByaCchDqzHgtgDaOsaF4/mn/habLG5o+1bylsB/xE
IN50xJUfEwb17wj70jQCxAwDs2P/ZH3GJBHjF8SGxAaT2MeWTWfFMi8tUr8bffY50q74BlTCOpfY
KaRY+3U1PNqkDcIEaVhb2z+ybsaVVzpF07sQQps/rpnm7uAY0+sDae5Df9yTxTK9bzW2rKS7F3Pu
ZSOjXDGVA8PJjmUUHHjzOvC+Z3QjZFitb8Lw2GjI2ovafVdeh5jmr/1sD6wH1/kmIMYXAb4fM5hd
M36/dE8vMzFlvfvIFGLT6DLOVYTyILvSaC5M08gkNX7aOG68cu7YtR2y7kklwxMnemoQt6bZyjPb
uWXHIQ6mUt3UmyYwyHk7UvOGh6/sPOhr0ofUnOjQYqlcYGDPfJidzM/tIjUlQ0Vt9EAIAf+w6h9f
KoLDXnfdxoWZQ93myF1OBF5QkApcPVSYimP0iEASC53BM6MdO23BH9h00X9ELqwDgHSAlkxqlvEv
z3TartTATC7aFumhpvM6s2z2CKKZeWLHBFyHxCrlXBEF22gJ78u12eOBEEnFeUdM1ZrS9gVUj9Di
sP5mWkR0eFT8QyCBsXTNSBabBEQVypUhrFBYa04qkgEC+I9D/R073eneooz2Rdf7DGujsjPrxMsS
quGUyWu47j+pMENAFSb57neE2t5Ahi/FsiHeL4lpQ8iy1m5uuCL8ZTxZ2CgrJGcJtZcO7IkBorXy
WtgT4F/9YRBuF5Ik2jKJ0BxsJ9/2GZRst/rXzVoOR3pQgzQ6/JY2O3L1dJhxiddFhr02H3Qg2nTI
kbNIWWEJQ1h9vCWiypIMy2Rf2qX1BC7HJhBPOquPtUvCMcMUXbRh1ntZ3/H+zs0CzncyLNIeLZ+V
TUnTiHgeaThVOL3m8BXKICXktPZfxEU6NkAMmXHoYknNqGq3ZrDjC8eHpvIUINN0RuOim/sYJYo2
Lt8fRBiWZ1Bcp53lND1BFchueVRKl+zjDhpACQROEWF481TjLuQK5KsADX7rjaRviXWpttFQArnS
CGgw4kJxRRY3Bma+UHx3OAda9iYj3v8zo0GhKqBLDmKxhWSCOQVmxvnNyhZArzfUUEtpYKattEPP
J+R6QpjKl56WGJyg0v9LA0dJpPk2HS0M2YcK7QHnQeHu0cQXoKO+hAQwVn4Jny6l6xVZW03sJ6CQ
Fx4VyzJlQyRaopHewhwvP6I0d6Q/y/fHBTkD0B1O8HeVpysH6f4Roe/U/KMX8UMdrXb6merbMz+k
sgk5AMOwJhyKn14F3EwygFB6GKReanbQhj4LHH6CKVg2TZgJYzWKTk0qT5/1Rwb2BuiDQxBiSMF8
DxHwgbhJy4UjDJJM02onrHk5SEF3ZF3wRbAj5wA1rKh7jrdsVcIoAzgf1LwNfmTFU3jqOTuPEswR
xOXW8QzZFI2ULxZL1qH6Y+kPFquUQPHHoq5KpDRue0AKPHr6fl4pmhtl9JIGSLKGLKkLkfMqsSqZ
wfvkgoc3zFLPtlMTa8+RNgOVSk3hT6L8H4Yw/cz3j9yeN7kFDWsdGWFp37qIfwMsMUwyW9AX+/34
NO7XSDURS8Gbqik6ywkG35k1G9FpNsuIG8eoLwijMdDS3bZpyRsPnZU57gisNb8vlv+AIOFLJE+D
D/vkUeYFnKfNi6eqUMazNvTimzJ1mahoAKuuT38/G6HF/3g1QI9M/pIhLeRLrV+TyWn+YFwIRUW3
WQUt7DjvmUDBELFSRu6UFk7Ys37lb5S8QerYCfrsNlnMjyz7G6L9kWfM1d6axupY3f43kJR66Yvt
os2j5valHgZGj+joAB8/g0i0XRS4OByA2lKiVrdIIwgv4o3FIk0v5ioZTvgs6f2wKNC1cIQghG9z
A7FrqWq00w/xNFJrRBSRc4XchUxrNY88ba1F9p/hXZ7yY1ZaeqU0GzVRlynYifA577IqsaixFQ/y
SArv84uAsizSx87xkopP7z7MP0tFTQHQxnWHaq1BmZDI0/LF2r6hFDmlNxc+qL/gtjOSM4SRobkw
SFKFzqw1SDMlvrR+GhFBMUWyV4gkARHHr0p8PqzE6/tPa3B+1kEn7ZGqh6kuxP479tuttWAJ74nY
teKulkHt9FfG0X/yJqvpgBRA5S9LVA5qXArRSozQ9KPhKp1m1WvOBI1jEcZgijPxIkkEg066NCip
sz+Q/a4DP2V4OqgtTJxpDjhFD9w60fxvaqH+cZ8o1o4QgN6f3tKUfRqzyMU9328A0RqSOrMB6JFq
J7F19nKkvBort38sTWgp/wOia9SsUlowYMzq82tjLjjtII6T2ksXnxz3yTOjt0AgtWm0mwZHPu5Q
TWTYoOG0YAJx3BveLLZRy+XL2TW0ZLW8XXjj49RKeIu6jwJ/KaogRZUrk+jUVWkYEPY1mAmb6JCc
EaT/PrBszA7ocdceyxSffkzArfSnU208cllzRF2TwCHdNzslkiV5wKhrF95BpLD+8fN+qO6bu1bw
jQ0Z+VlH3d0+qRiVENNSe4dwJni6UaoAHpsmRihJY+KwqNZHCrfrjgQMIRRJXZHBGhWafkRP7S/y
4uRH3lO9bKxnDpZsW8XrtVz9K7rbtzP5SF7KIV0bEZhf7fASV2Wxhpsu2BbNceWZwILk3EzHqoQT
WxVmDH/lvcr1wEBdEqfblP1JboHE89UY5e+HSdIdfF2KQ8qHChB1x8J0YN/4fqLc2zx5k+0TtJO2
j9Kn6FkBoHoAAcx9LhtbvaZhJAteAVYlhWFOaNV/jwF4cDcGwhqA165sMX8A+jfYKtS4UqqiTWcu
FhX4dZKuBsrShVN+0N4g7MVvmjm9a78+YHiFzlHUJDCSMyp8u2NjS/OewMJKifVu4iWUsbueLYDK
fKmep1HvJtGaok9+gKnHNXa49N/Wq3ImfXGnE03Dh/wLpnXzsQ3jNnv4E+1EltTCpAgQJm+IlPzQ
ASUCSSMI1mgf90lVfxUaac6C8E03L1tIPtbkYYyTSLFHqL+2Z/7yS8RoGOFR/4Q2SyaqZtHjabcd
bpq6pkcDIJLr9V/NskOC1ZMwdQLHuj5rvguTHX/w4US+OJMNHDZKGl2DFmw9tuJ60rO59RbzBzw9
muVlp5eVyLJrMrQOFnXpZxZYPFTmHoj8b0owees+qd6RHD0iPoYfdF9HHPKouq+Y4j6MXYR1J2he
ShR8dzHDkTLK3suxkPrje7Zp02TyAd+q0XuL+uv2rN1uARIY+3Xy9nPsyFcAVPGGuNIqzXQTlbhQ
fSI3TtVsO9yqgA5ndu9tbCcDd4EwtHhWfL9clQVOcEE1rLNtGEp0wmS3z8d6yX1EYBgP+UtG11lA
9jVQ4Ieo0CbKPTa8eYRhIeO3g10LSgTlVQZCNPiJKdurqEDnJK+6wxM4KANGpx32huP+y02otznA
skNTsSdxFLfaOTDrbaaovkWwrj36xeMinGW8i6lnDEfxQjnGB2SHcFalmh3plsM07nWaq2IyPz4R
rA+lyzvikt1iT/Xoc3EvhVTSXRaYvBRNeDsxl3TvXa9NwG/1Tb/gUI8syCLx6F+yvwlhzcuRPqid
lhQ5IlmsnMvI66cB0xAr6d+IYlVelPQqYAmGqgLvX9cw9FpTGLD9Kp05DZ7FujlQjL7kllUhuJeD
RnbMzJXx49nxjTwGpVoGp4iybqT4n+JV3C9iExlGG+7Z5McB45zObUzzhvHcDTk1mGIyZFG20uqC
kwbbJ1Iu8Yjmcpwn1Sw5hTxBh8iJ+JbKpOc+m2hbQym9yqIk6xdBo4tDVemEDkrmQkQ9/s1XJTp7
z3MdP/WKrLjY1NRdwvEr07aDK2fW6iDwB04a01w763dW/0eZu5FmqMO6Y7gyKCYKdJmWy7h8mh+o
FJ2Ck4+U82jN1HHPjbO3coTAJatJsmnf/3IRUVxYfaTOhvGXWtLodR1PLqbDJfdJoVt2URZrfbKx
v/fkMmefhH1hFsvQ2IhpO8I2kaYaoMbig3B80//q0DaVbqPhFa+ExmNrBPicC5UNs7wX4MbQ0JD8
EvlYdhyMmCLrNI0T534hQPGeIPXplHBrU6VGuFNSRorP+EkVjCDHogY3KOuLoNUDIJIxk4619sDa
iqAuCUYi4AKaSVgI7Utix2lMRZj4XfvF38EIUrhnsvopkTYS2h3LKs3PVysxeDsagaJ2018DFAE2
KcHgc2bGKdlFpw7p9aNGz+2FCF24Oe3MYF24Em7kfdDMcHPFKFYaNcGjx/1ie2E1iti5JY7ow0qQ
XeNgErOl7kEz4uIm6HoLa9ila7GPfKwTL+zktbqouTGvkGdvZCbSggVF6uB3d+XxYGq0xIcDZ7Fp
Jd1Ytrw5UWsmq/LCJe6EzNdSkCIIPCKYAghXX9poAPnnFiqiQsbPc/+3UagwFLB72IdXZ26eTYCD
C+mS1NtnXE0ppvBx6h7VAHg0CTv3XggFlVgoZ1Hjp9YlGMXrZrnOMdVtwA+FKMhbDQKxYMzsPNu8
wMWFnXFSILkoRTG7KU7au4cmNqSs7d8d0wz6xVP9x9IUdyKilEfNGb2yLaYDJ5JQ+G/cyinZq7aE
eoQS6jQsczya8FujuXPLKoybjmGB9XLBx6LABzmtS98pYtnkTFif0IQtPhdl9vvpoB5/h1uGt5kj
WUoP+6Q/sRGiyVoYmntfyTKg7tZDE9grMT+MMXfvR6/RlqExE1w7vU1aJbZfLsQDoX3jJn4hLiro
fx9zkBmZCUM5RmwYMfML1Gbpzo/i0f5KW6WVbKcf1Nd66S7KFKUWtJ5jV+JF5hGxqvyVM0p+N0pv
Yam4zr1Qz3KP0jAVEdNfGGa50WQBCdlVJQ0s/rFakIZksNxNgHLhD+cnG6ynnq2VhhxobAuCpy/q
UYqSyeADlyzuva40umu/kRFm5nlt27MuJvQJGsd9atFuwDaN4YX2wZk3rw0l2LMXO9N/I04HoVgT
f1WNrxz3RmLzT8EkflB+8KupPhDYtGVHnpscz0RtT6iOabgLCBK9Wjs0vpL3ZSs/GZ0nDHZimYCa
rl9gI4AVcajWKl3JQ+BH1fVTH+2uXfyzksJHpvskxwVT5xi5VLnrlycLpGNnFSIpnNud9nJi4RkK
ZojaNhjriRVyiMDcYpobhjvTH2LjSSkQ369NFj1+AddQhH2COEZHXXfeQZNaGcPrmzuWHY+L2KHO
CVPPplWR89dP/uv5dL9MIYiEBNOgoXOGAB+ALO4085+AAiabLL8gDTLgM3qoNlZeVq1xhDMqXmEL
oSiKe8Ju8092G17dt8iBWVFG3gNYg/13Ph5/ztKiD4BK4TfRQADVoQPwioBnOGmyDhgo9LFZIdth
6Snc7ysPFXPQwNAvOAaojZPyQpfIVRiOD2mRla6nnHM+M8iruTk1g3RtgUpXTn2NDqFf/dZ//lpk
cn6QRidXLa2HgsplwQFBZ9qzu5Um4QOwycJzUiojykIIz7P6ZBlNBCfs/A+2PzcBI+s2f32VOGQ9
rZ/WWN17T5uloWgiwFXjaxqvK6sVO4HZZcqGW7bX/2Z8KTN1vY7/RhDOomsCi5NhyTDlQZ1VocPW
OnVqhkjzO5t0liuS0u9vfbx7Iadw0lhHyNepQOw0VNzQfYs4e0k6dXmBQZinYmcJAQzFdIQ6NiSF
3BNkiXMqSNhAzTvf+SqRIZq0CJ0ADm+8//Ir/CTGAotaLS35v3CDBTLwnk4vdXzfU+6Itoaq/Dby
1TrnvxSOHzKIMmi2G7zozQkST4y3uyeWc9saN3C66zkXwXFm2Yf/67B92lrV302kfqESLCRu9zWe
O92WzlX2AOXvFuqEczyOk4oA/Tx2ozdjJ0VOW+/3P83ACQCGXmcZo6bArzW8d6eyv4Bpyd6LFTTg
kRY6mWKozpAse7g+dWCU5TyfVNORFwJvnBHyWF7l0zdm0X19vZWRGQCZybagq7zvnmOUUMxF98A9
S/9KBKh7SJcf0gXq0Fr4z16Ui4H4nGZP/D/+/JWzAm7kNYl8VWXDarG4zueguq0xF6+OTSEzOqQF
0bhR2ywi4PfNQTzVS4dWM6B9N3CH4+wlES1mmw1zhhAzLqwst3RANh4GW3bdUwiK/N5F7AVA9OUR
TptSZCNDyS5zhmdbWnudPAazI4i2Lt8Dr0DquRtv0H3AnB9xE65/PHMA8B73HBGwNtbKP0zKjm1A
u0Q5D52/PL4qETH6c7vL/ptngA59JqWpmQD34T3R89TOjiqtSF8wiJrC3O3toioDOUOibe+waqIc
pFK3lkrtAL1qVKXqlIB66u+iGf/R+1wZUTSMdwFZXPPfqmXlLcSonPBxlYuOjFWL6sXZQwOF1rew
XKS07pjYW9nv1r2nDM8mTpF1ONJqzReA3aJBsH+jY4cUMwPLWpptQq9idR/a+tOAZn98Hianf6aV
JS2/KHDks0TB+90i1zguFAyBb4hoYMBaTmYZMVvhdYaK7EEhceTxsWNomr/WN+R2i1w7Hen8bYwn
g/n5FsS44Jp7zJcEpGm9buo0KZBWS57aF3afm7Tq0dbR2MuN8BEUiQDOZw+vqWjvMusQ7DmI+jmK
PSu2YlAs8sYUj9IIEeNqvlAN7bUk8d0YP2M1rrnvftLkjbnsJzCv6SVnvDNLa8I5Ro5H57HcxIYJ
VnCivb6+fjySXyjULVlloeG5DuByEEm13BujqV7UBT0bvlnQuJVfu7GA8tIlo6nMl7JQIE/jOlmM
zK9OV8xbufl53Fb3XeurwXafHt1X6w04ZpdmG/KRpVaIw+HNhvvgjpChSFAUDkvjiJP3Hoxi14qV
8uXARzFKI+9PV4+cV5Gg6mrnKzLlpsLxxAEJfmsgLzmVFe5zRDXLu59S7IwNk3YJpoBFmrmk4Zjg
+KNU/oxKF6orlWXPfGiFEDlYTzAuQQGhxyLKfxGzQlODVmIhHTyYQ9vdeE7jqlqALwZ90inP5Nof
n9DJw7gLzYQr7dbCQl7L3hKioHhIq95tUbBRqWEbdOt1VYDZxaAF68m2dGYGVEFsYFALUf6e0v1M
NpjqfB+X8EZ69WZEAdWFjXlhQzYTUppGjNcgZaXbcq/gNhMGlbe6GDhDYiVCJLEto5X8Ifi7bpBJ
1u3q41hu6bH92oBgG5cYsd4RgN2MGPts1rCWMBfoSLPYdSvOh6fm0+zkhZ+wnJMImWwjo0tkUuzR
Fs0DVoy2BRXa5dfahMyGbvjdYKx9eG/i46UpTEN0GH+ezj50/woT/lmqJvlxI2pZq50z2fvk6Tcf
QOmai1ZPv/YBY9uRC6zBiWz9okZAYihywCQULpWM+zZ89C8MEG1pLJOjiHutMZa5Gua4q6ODX/VX
G6LkhRE4WQIX31MX4yGSsdBH3/sFl07AG6/aQTC0X5wBPd0XwuWDFdeAkkE9Sw615nba9qdvuzyO
4dUlrXUbCSJnWLqgEad7UL99EvxNjgGCpX42Olog3ExBf13i0NyZRKzKXhsxpgP5jQdiD3y7Hjws
KxP0zw10PH2K6z1Ci+kBDtHy5rTgYHto2XZPnKRgmDeDkSGAR14OepiIBdCam99vAWacNLHSlFrv
ziKzZP/C1R71hHew7ztD0tMVDC791hCn/daP3LBZ9Uugr2psGs3LVwdkYriZtePmv+lOSXMa6Kbr
l9v749rfj1uaGe7/YbWOJrEQ6y7IOVEJD0yI2mcKWrF0i2i0DoL20yNI/aT0Y8r/mSmhARHxdHSP
OJuwXU2ZaLMeMilP5lguvpQH82HZULVwKBJUI5mmsYqWcrYnUF/3UVXGBOgbnN5sTvipRBUWfGYH
IaCBmC9JfO2fIZpbU6JMc2U+K8L930HQPd4CrUehIslBCgyTc2jdk8/GnbuzhArWNw+YJF8Rqr75
+27n94GjxkODW0zCjVY1JnSGRa0wshPrA2fIL6dV/5hHj1cVvUN76+MMn8CTVJkF6XbG0DOWNqE0
kpfx+tw87higX2Wb8WxS5oyRvMvKmVBOY9vCN4Dc0bgYdJUGLEGSijOPW6Nz1lPz7HUuh8iEfeh2
8PxDCX+M2TjpncoiG4pdy+ZCDbvT0Dd4uhZggYyILWlALdwplI/bVkpoykK4vqJkgfMG/2Yy3D+r
d2uGfIcICCV1CRjxruWlznTySFmcWJcsQxCe68NpvN0Og+Ly9gPYk76vp84FBTSONxQFPRe7bPn3
PR5f2hA1J5wYfpAslO+yndai5Hkl6kO5dJW8e4A9HI9nkdWMGRHBYVjOJA4b7FmX98ju3P81WG7s
Kz/IBAV0y3Dho2PZ/h8hmY8Ko8PhUNV+rs90JYb4U/U2Wg/iNkOFWjv1k+o2hs0my+Jb3gG3jSB3
WzjancL+YRJM/Q2OhQ4RECxZE7dOXTd0/ctcqeTLEBprWl8PTIwQc6n6s+FE98TSo8rzf5ZsDQRM
uwgvnDpqL5ecQWphx6hGo5jNtMdsYlrMd1zXyGv5INVoad/rM0TWXegRhWUIm6/B5TOZTvcRye0Q
0d6cUTm3qw+2BO5o3Zsmf8r9eiw30DmR9LQc7O2m71b/vjvge1c5VQA+HwPjfpQ6bp9XwljyepEP
78AS2OyfaooZypBZvCHQaomEv2/dOfrrvb2qjJC9gAZPRXSQ0kld6hthc0JsQ0mXnySW3VbJoPDz
K4iJj0utOLWqymQsD4Yyga8n0lrWPECnbhZ8FQicEjhiL/pZ4DihVE/IdYG73InK4+4zSKKdfaRL
2CgXbqj/nFACZyYu2Av/8fWKgtDDOHTAgKIWQhnA00+R2+mDHF3Brl75HaEdyNUeVK/2InsPlis0
rRLoI12KDsB0ipIa1jL7lITkfDA3hWwMxIoPnNmQhI85zeQKO9np3JP2h8fkCE5RSxv/IIlN90h9
vmb5WoSSyiZSYiRYLE0U0yP2Rm781g0BGYYfHT8LdqwWSq6mpZ2bDmPRSeEVjvIJXmoVoCZqVMP9
ArY/6ad9R7IlQCN0r0565dEj6Ej+i7dFPV8V6HBhrOQxuM1sPzD2Z40f5AuBL5Sjy0nxUifhQFOk
z6BKR8M+7JLcMzITQvTwLk9HElfOR7aBdzwpFxC6k1GQLlOq9PmOCTmI+IbM+fQOEpyu2dgizO+f
0AlmhdcB2/AMmwJ8rhhvv7jKnCgAlSZUC/MDVcupc5BC4FJ5Rwe97Se5JZ7vXeFcJkhQJta5hc9a
1J1YRDCOU5F9pMQior0W66wa9GmtC65OhnZmb4/O5YoF/cshr9pWfN/J4jvKPF/hrVCBVDldgon2
ZDrwr0QltVNFG6AqDLggY9nKS8cZmvXYmMYlXsFrNiCmwB2gLgOiE4Z01RpAApwE99EMZAfwIFYU
ZMCm8b+As2TwaXZnrtcx+AGReMudp2rwXdnJ75oSxh8dRrwskwkBSg43bOE3tmooQXVpN/3mD3Tu
4GsjY0/FjgLx8ziH6w5WixPVXfiCIjP/wHqBd6iMi7Q7hz4T4pzcLEVMFgPe3QpurlGkzgC4Nknk
OVbjM7TifAtzG/F4afauxF+F1Oum/RYDkCtfTgYAE2WwaDkR+iy8j5Yw8LdI+Kg11w5FvlIbvLkB
7JrusWvOH8kAHaipfWcAAtUy/1y9r5S7j8spNj8B/45W5TaG8iRMDAiVacVEQvOg0h2kT5GrWghX
9wou+8df5n1R+A09xMvaz7guv9T7Y0oY2EUCSOMHBJViGJCNeBzpxPR+hHXW5ESE8grmRtfiTQ9G
+nMpfYvUkBRWHYs1nI99JxQBmSS6gxkKdeObtAtbs/5pQH/vXhjgHHv1G5+eHE17SGUVF5ZtAvPs
q6tml14If5IU3oWl2Fi1dnUhOY45TsCuJNSbb1WMS/rEdSGKJCwQbSBLvGUv3OOSXF1l500u2Hje
4316bZKK7mEQNhrcfhMLzraEVJr5bsbN3epM3jKN5RVfXSWAXfm4LWBdbI712xGKu2w4VyVgFVuA
xz2ncpYy6+PaRmnGaHo3QkK+9Y//G9cmE1zSK7iMicdCP+14G8LDxckIDnXzY65ly2H+5ZD8J9sx
BhvUo8br6tklDuegUUBKkx/BkfHJGD3g7ZElRYQx8rwEvRWT1wTQCN0JHn6Sus4vAWswitOqjnvm
HjRQqSmW0cT27xcxIvaYFmxz2kFKeK2hCkpmyk49bhIOtfUiVN2umghzvXC6mzptjl4zCKvFb+eu
d4szX4H31Ylvtu2nTL9LDn5a8O6SivOQEIHifK6iQx66RBLyoEnnTAMehpdYgt+APYyO+WLxG137
gqLEQ6mWWIBB3rBuzLVDtFF6K/YQK0n2cJ/+IaUu00Q+sBeK+U4kqHDE2uBG0EpMx389k3GSO/9z
ioUrxzAwNY71uPmHbcGImmodbfk2XMpsrWhgQjZW//lXUdG7/W6qemqvo7OeNDKFfOPrdipzI9qv
5OImhppmuBI66UJpbCGSPB8AWVJgNkH9lSDuuS2Hz+QPN3nZB35uQTlPXkvySPuwDhkOdhdV9cNW
UOusoqfOaiJH94ffixIqtgnzm4i6hBFsF6Ru0dx8bLEq00iCipdybweMKm7eEQExz6ERTOqFeDB4
ZeR5pTV8vx1zLhAOb1pjWP3Sh8fzgwC+Ura0hETheJMB8bXcBlWLi/hQZegee6KxzQk0A5ZJxo1l
MfU371y/vsOYnhos+xWjaVXmvOmxYUiJRkzO0zntWzCfv838VhnwNGW7De86RHx3ToscNsElGw1X
R+8nSalonWiSX/l22e6cvyDkFXj5ZoLslbLZSmqflBpja94w7iX+QfSKoKH+LhdWk/j3RrU0g8Ov
5ltw/cH0rz0dBza707i9696lyEbaiVvvwiIwlxAr+HwCEHthLW7W/HiLU0pIT/f4WQPuFGSmNxUb
J+rqrIvnkOjNornQt3c/LWeVeSfOqh79u7LLxHrx8K6XCReKmQV3QDekwjp5+MCD1uKmozLMX5Bu
xw60jliHcyWBmDuLLExnLAZW7rMn+iUx7uMIeTM9Uz8rMlkAyOQNmtsgNyvaFCdsTBgMe/hcwqEA
Bwo0ExNbeQeFl+DKhbYMc4Scqm7t4OMPdUp6AhJfN6Rs1VCgG/Rf8lkvidVCOOoUfcP+MpDxxBLZ
cEPjJxGxyasu5WpjaM/dmRWI4pH+/oEdFk7YpKEPt5cI5DqHHFE377B4fxJSD82oaT00WpEEqdyL
+yaJ6PI5Prw4RTnmFLqBsUgXFycmB4/qZNVpkkUH4T5d1lx7aTej2OJJNZK0GG8Ys+ex/azdp9+m
GVX+/4V5FkIzJxnLUGNEhAvoqyl4zHuxQRaK9o+hGFB/j97Tv96LKwEj0IT/F3ttr+oDTSn2F1n3
YCyafH+k5xzm5EN/LUwzrLnpaGSwRxmLA439l2Eo7N61nC0fRSMLhz7G3fZoNx/1Xj2tW6nei8fh
hbJPfquTvYd2f24lkoi8fnJMHHVIxtILIEB9PQKcT5dyM2SHEyiypSNes1cUFKt3tVDi+XzNHDKk
GsFTsnmrvK0EcFKIn8Gyt+DAmdgnTD5NHGuoSVMLb0s67Eg7PF19AfOapHar9V5KMCpHEUm/fl/V
chQKdOMf9cwXH27WeHrupErsN4UOBCA8pobJ7RmAyp7UxXmaG4NxguTx3KnbsSIaq+/obtcfnIOA
sYjSTGrfnK9/bDvxPYDxvyzx/gOgt/6ZLqd5V+OkX/faCJ2behnBp1xliUhcNcDcvuf6cUCdqIA4
zMj02EfQz6aZocjLqj1aGUw7M8ypaLb4UOb+Myo+U6sUThHd4pDoK1UmxRsB4iufPOFZeJwB+kt9
74ZHlFEyvQCvU2MAJTLnsf9/fLd323gJnb9Ls4DvzmLZlbuvmFEmJIPHoe38v5wR5XKEhxEXM7/U
1X846bBvDSgIiFCtKNaXeHtJ6Tfhrm/89Vfa8RvG/Jl0osVnlJ7+TZYO9LVkSQ+NM45kNMiFS1z9
FBue6/TDDFAHZJ+hyIoHITUbkbQ/t35Fem0uQOOTYumywXKT3b5eCa87Yiyld+pEAXUghCVzoG/Y
qg3BI95Y2bbjdrBgewre70HdDXoOaIvfJz44oeN08fcD1V6VLDeJqYcw8Csq5Q0gqvoGf79WljZ6
yjeMJnQtWR8XvRjyqzlMGQBKiTrSUnqwDOk6noaz1jHo4Evc2hkf1hCI56B2SxZiI8Y3qf9Qz7gW
QmZz0La+FzHgSgr/bq4fCWG0ur1dRZIYh6BtpLIfWpNrsPPE3mNBBlwVMJzTFpkGnEWbqXeCgMC1
2R3cSnaHppep775EGOblJL/xQhZCR00vfcqHwGur/W2fXqsnFr//VUW8BqQGhVQ86IuojBFDN+mp
RftV2Q+QozkTg9vLtwRW8+5YLxitoKtGMSvJBomEEHl4+ANxvfRTaXg0uwZkELAuFZJ+QvEBoHo5
NJsHPPO3vEyDqBZriHqzMjrtMWslZh4cRHMfqQbXZhQs54A+4A9Z1ZgUXmlUpv8+1VUGeByV6x61
oAWv8bKNAkKZ2k13HdJGyDtdHFhjlJV/DHDhMta7MbWBkYBkR2IBGDMTlPl9w8vWkOdaLJgkQcEs
y0Bmz/M3Cm/dRUlrrOTo8RcJOXnguq1ymVzSnyLF7YIvwz6mEgrtQi+LxUSXX7yShRG+SMT9zULc
lEEoBnkYuBHZBcv+VTt29c0kOQFoD5Rb36SyYFedh+mr+Lb7wb3mYzboF367RA0EEUbcVoGVMxxW
NsJJ5S2/Wft7yaywkrsnDtYkhHkOXIEDjFiiV6/mDgRftO7pQ204SRfikwsny8Xx8u0zvEICkbzR
nv+Iluboru2t9jvaSZ3IwTWYa6kaEYRdV/I3ZPVRBFABkzOmSrpkL0+xe0oysy7y/FfiLHsLYKLo
uiuI4QaoD51BhAbAN11aodmNJUNYJ2AbKiOc9DztlVcNT4Z6um+V56QIJFQRbPFNq7CayvBMQm4E
BbQoYWPv8IxBJf+rV5sCJfJotmQ3L03IeZQ6DnG3FrtCFaI3mfE6nhNQFs7W2za0JxexKctxs6BD
FaWBHISO75kzZsn1q7PnjO5pEJXW8+9486Yt3X45MyT1HJ+4QnXjEw6Egz23NvsItUKbYdM7E/iA
kdQ1s5aA6DcdT3A0v0TSyVsO+eAHduJ9nbJuuMUnPebaIIyEbFlHBlUJcMmUZPiSgvBuBSv7kTbk
IXW5jCb7oZLhGwaqK1ULmfJZLCpZKoO6JZgG4o9Cra7rPXVCayylfT7ydR9nnCWg9ZFR8ThVkkfn
oQJP7X88xaW0dShWWeUxT1Ea+hzeBkboRAWbNYKSadL0Ipm/oDy3ibYgn+kaahfyZhdmMrpgmcaZ
yq84RP+g1j1Db2bh5Tov9yiGNfSK0Pow9B7HwYiW9kvLAQwnZKJKnNvAbiHHykXS4/Jk7rxucY9r
kH9PUbgqr3u66CKbJGcITt0FiKFqzEbmxGjXlmfVs/13AeYpiWwf/T6pmr/TNrINOhIfs8a3H5aq
QmvfOvAtlv+ArBkvBz27HjtFqoNZKe5MoslCr/1tbzPeryNNQtlXpXydxzFyZ3yLulPG3lB8vyZs
Xywk7r+KkTVvJ9Hetx7TbL+mxBuEl5f+t+mIiOS3ISgLourhpjT6R7J3w7UPYClBnrpQne8F6107
D/n+IvTqSmPLTC7YYEi+2yeYuPP9V6eOcN9aTrZ//RwrMVxwzkU+/I5iZaVnf8W8Z3JN8KdEQO1o
30WvnJMdrchI/r6oL84Ay+uqopA7esSKK95bshr+fw+0xt55j5V1PZQmDyLCW0oR3FUmo3vPIr09
GuBVCC0ImiloFaah2JCJ3hoNC4e+MwW2IN14Oh/fxSR8P/p1vjDIjzV77iyMpVWlKqaF87YdRbf+
QHkIdbjgJFeyLgCS+LLqPmz0zFyn9htu9I9Ps8O/vfbs95ifhmExqDfF1Qw7N67N5SxBKmQEMOG0
D/TgB/2bMZoLTRtd+PGaWY/9X6XCJST1txxrANYoyyIcR85aKF1EasUTH1MS4nqv6YolFqkfC55/
GbyLMg9D9f0Lskyx4FgvPFq47tXUK/8n4F/dSfRbxvFdEDS/rCHN9RCPeA0LQsK9Na+LIRgHEBG/
BxOJHjNNiW6zA+V09ouIMn33y3B1Zw4+yDK07iEinasKUYwdUYMT8Ua66EBRCO0ZNrldoqVFc2q3
eoN5PezbIWxUGJuTIhxbtcXrgbWWcvPLbiu+mIvJwMmAoUTkJFK6Yy8eitTDC+8gNHHoZEzJYuVG
xtlyUYY6TK+u+KgnHJfU43I8XlDUZ4j3I1g6mcgWju4QjaFbRcVHcfuFiYroOOdLwnvnQR8I0szH
+nxVXm1/djb3byoByY3eS2T0vG0MJXoznbaOneMXkoaOhFvw3+oDEysHLTxYWwFjBonFU0vtkF2D
WAmIWVbp5mbsyyKoDTe7/NoIvtN2KmLkaZ8e9f+zSOhWH1hxAhbRnJo2Taefz77+Bxe+7wHDZ3VG
V+oncmdqoJ0Bz3QSoiZVLH+jwHOZJYe6fFqBdqiROZ/TYMmNFjASW/fyM/qEDM5RcSPV/yfE9m8M
8hHJjjEpEx1pFpybM9p9lclQrGZDAaAEhh5kygVAQGwcrQjkbTPZr6MqJtw1YQ0XCbqvDa6xUZ7G
T+B9lCX7oXgEClAa5wcLz+aaTmFd94K9E1td8/nmY1xFyDW+jzbxX1eJXFb9+zjcsUeHXksMxVp+
p5y8yDFNQs4cWbDQtUrQkv2s4PCSPwOjoXFzXtVDWKR0FkaWSSLiQpGsqhqZduUiSIqjPiPADP5x
KCYYeLccVWRkvGO5FIDbh1kZZU4ktKKuJiouFyMq6SDdn9qzjFtp64d6NwBP7LvpKu+EoydQIhT/
sqPLx1y6fXoZs23wGZx1+Dcy4fwJSyZuC7cJFr0gOkUp7IJQHRNkpMEe5tlD3bWyBAzGmv08fN58
/GDuRyInpm40IIMeHG2y7Q4NecLda8BatVjPVFmrY7hh7xLVTx6cbc3lkUir7TsUvEOymLQw0eHz
uS5fgwgBG0hUROgXjhhHeAdd0X7PcOA8zLmezySbd15RjiXUdpsUR1TmucF9fAjtV1PjmclZYYiH
epL12+LRyPH9unXiIZEU9bOu2n8yHfYzlnjChHTqsQRKZWTyO+v5a8f/aPdUgzLwXBo97PiYnetG
RHB/iBL9NaQ5KbR8ZbkmvORPa7UrxvfNNdt83KvyT3qGOOcpSOA2y52mqPN07NOvJhEfIYPyP7QT
kjO/vBQejCMhpsfCaREkdFxQhKpsacE9kDmEy4W4kk6+Z4oOLXfxPXH/KRPYbySRAkiXELfVyM/L
ntcOUwynz1I8iJe558aThwmPGIOa0qDuNEiO78z2L4bz8IhWxsbzMWT9Ej3CCvXBzCxLJT/BzHMC
iM+/+9IudOnfHD4tBkXDn0Ip+PIZV0nic2imxM3KiKj9p9Mgy1IbAwnHIMKrvbQSUIFyO+lI0I9n
D+iTibUex6956rmDzvY05jX1uibOClkjUvTlsiIEZoWZwEoGylW5DE8h1efFA50c9TPeIULaRuI1
dxMeJmzZZFDicFjilRQ1BTuVzQRRsWdzxl2yun9yMyotQhx27K3dHhd9MdxLSbjXsGiwNdKoq74E
A7HLL1cOs49n2pKzqVRIGQfe7GGmZlf9Xrg4vGnvg95s4DatLDS3+sxljvw59rS8mq9cHkKSqI+x
RuT8Qsa9t2W4AbIBYwuHJ/7pQFEo6HbFGwWLuk3ek0+PPUz1sTwk3H3zE/0ilFE1sOm/fCsY2Pbf
6xxr18X3DMW1k1X075IR2XNc5v3DF7tH6ccQ1MsUgvy2+cdUHZHuhx46GotN0pHx12BDNyOxiyZw
bJNDWd8w/IG1EvBlbfQrhH1Qf5au07ropJiIa2UivNzWPXDYTqTR02GaIqqvWzUKf+3FKj06W0QA
YK+hKHxLVQTmKRcgAp5uyqkB2Fw1tn2kVugf2egOSIRP5qJ6+VGLtGDHAc2nVFB9jV+SjyUth0wv
w6Lkj5iSXxWe2e7G13u3u+NEiMHv796JlBY9Qp63QHZIG/Fk+k73PYJSr/3VtCjv+Nnrw3004TkX
kSxOQtFUy58CXARPq5/1wPqDIPzL+F9txcBIrnWSYTfHMAt+WsFt91SXXM0PCXu0Fl5HcnePHZty
NEcYrkesebaGnhPTuSrpHkfZnlyFvLiH5pmnwVTGEwVFpZCpdMZVWDGeSe5x7tjLcy9JAl3L4Sq+
S+hTt35j+Y+E4gXDzKZLyxNQidgCxeSqIwhRKPzeYXW42Yrx1OFLuBtrAUHkrq5JISpp+2LNRSwZ
hetrtQvZEVMK1+v5jPBrRl3PQuixUptbH6++fiAAfXxqCnFYEV402XhESz+bwFQngnXCDRH5ODjK
lYz7AAZu9Hj9IMDWQOwwDcp0A8j86xFTAe5r/IL5TFoSvXe6lbnskHmR7EOSXLUvUNdbkB/hOVZY
qTh1H0PfFhFVdYDcFLII0rli2HwE2UPcy3gHYTK0JjZv0hQ+bF/5rCSsUPVBg9nBHT3DS+6vW3PR
8k0nCem5DCA3zF4d+emNZHdR7PEbV+LB/X12/wQWd7X9E2NfyHPd1UmrtBMglO/ufK6hxhmLBqys
rwxgdNPNKJC+lY11H8KilxII5VlyrRyzn5q+GvRigpqi0dRbzLx7sP1MzBy9D3BJDwAJJl6VmKwD
G86KK+0k5qEfEbEUayxvy8mzDsiYgZRdG76dYuVQN3lkAgqLyafgwHR7Rn9pUH6KqMvhUFiIKmKl
kHjgtYKfXfnAJX6mSrI2VN8xrU4Dpvx3V/fyYZWQTmifyHSsD+L86l5VPZu26pf5OppDqvrYWJi5
uLWQQCs+bh3ortIMnORFiUIanAGtTQW8LrVwGh5UzgLYPAMoPg5DCHo0B3sphLE8WCxf/XafqLfN
P6I08T7XaL80i7yuIfK+KgjylVlRZ30Jc8V+HZcFUSNSWoJCHjty+N8HrmqrpLST/z3avvPABu9P
H0Ia3VPGVL7bNHBKkip7DwQWiPp83/Cn7HVQztJoRngJ0qAeTFlcPZxdr/QjN85z96twzjmdI9LB
Bp4xi3xSy1gQwCCppocllb9RHs9DIgAt/iCKmhMsWTnZLKshHUm4SoJ1BLrnrJqQLBQYFk92xWxm
VRzTZgbor1DkIR8woT5bF19WpQzxVHyfD4bHWyFmKvC5YW/SHahqBg2KxGjeHSVgfIibAbqKQWwz
p2U8BpOBE+qFnhOJYp30VDNj8Yb9sDBltcuawnu4fGd8do1t1LlhGil58cTRx603iZQTeFFMRJVA
/dKjddskEN7BFQ8xqQV9qKZFhoaRtSYiVL60LGtxXKvDY2rIOfO6FkDFUzEcLaYMMvJMUDGWWLdz
cGzYe0CtCa9j7AaV/s2UnpGONRCu/AWXNaIYLlP7hArL1DeN6HFRWs2p/HAlYrzjF1+WCz49/5Tz
Ow6ojzgC1MGaC+BKmXdxw5ppngLiMe+9sKEkcObCLxFSiRdn1+FS886DCLU+oYKBfqWtOnwUUU2P
8nbbmzrQ6kmJudosDoInnZs/USMy5+X1tfB+KsqxLYk5cmV+eDDuQswsms3Nh026Y7wCWc6MLcMq
69sHEi1BPZA6RPr0qDXgVohOnhfVV/hktRaB2rtKjvBJojQnXOiQdf4V9JyWWO3M3+JMttjFiGLk
tWONSrOTaQnez7ueGTuwffHx9D69fbI1NActifwcYj3qHPF3LAxVuWfa9TSYlE/p4ZyeQXJ0BUww
LOan7w4FT0X/yyyVO+rIjed5DhNC1nqYjrlDLZlX9Q6pa++ACdfJHBNxuJ5YG7eCqVrvcIIA7NiP
lYxiKBPB+XEm7W4Qd7B9MT7mcbL+PYN446wvxnBHJ+szvWW3es6y+pqZi6ppLftaNPq59tecJI40
4hdyZV8Q9XJ5xoSLTrHr4v8/93TfKcwmyCoOg7WOZQj+arUroE+R5A0vUH7xPm8y/j7F1jH1KjvT
Jc+x3LA/fpLjd4UQ+QvfpALjRJLMrSg0TAfrKqWQloK9gdXY2Myat0igOuH+261tvihPfbvRWs9p
xv7sswkSNYq5PW6LjIp/wAOQnWKUwVwa4Alf6WM+YDoKYN6U5W9YtoECc6ptn038MBJ8zJkMxQ32
7RzZPINX6g2026mRAeK+GzN4rBDxyQrbFrKDbLPzcb+cbxINfqOu4JOPQupvCPsqODyekRzdEoEU
0iPPlEHtkEvazErz5dbeawHf+1Ey/9ZOYBoRY6csv7OkN5okdQS7oKee+vQU2a/8EW2A9MTzHnLv
EltKQZhBoOzjyEiOO438U/73F5jtYrf5duFj0IlRgmStCyNxSiQpbsXCagv17zclQzUETy424IrN
2ZGbRbhdYlGu/bMR7+i1AfGj8usZwaVlTTQzgGnn+GLR5MqXeRQgFgR9bk5CCqIDOg3viVPjjwPn
ylPRju0iU0beOCHk8V/Nz0lV1H2yUvIWgKTKf9O+iqbZWPNYtH7AmMkDhpltFVbITo8xxAMsUkKQ
csi19/D5hKhFQoYRVY4s4mcVL8xHazsZa5sAEWNZNXZ8ys6U/5pga5F5cyYMhkG9plK9xK7TZsmO
QIsoWmo+VkIMFQc/q5jkWWLk2M6fjfX3g4cqUoeCQezuNuNQDP+mGaU2jeaWtMyrbVcr6hXC6gmZ
rfkoDs6zdjxucOoSqDI7qis7CXe43JNImPU6Wt1eLKTNBO3w0uBs58TX0pM+1o9V9cAkgW1gofG3
RMW5scKAZ10rgasrLM7iipcM7CwdyIhrRCdt0CiZCIZVMI0eMdVdhmQIrR0WFrP3T7DCTsdwt9IF
NeZmqAI9Cq1hBhiqTjzJQfowf48Teu3NfdOIV5u5RwsXTw1fljzkwGjnS20pCJjIIOnQJU+79ayS
kO1H3Vf81a5F+Iir++p7fSxWm/Ft7Uuj4PYZ93z5hUIWx1qM7SIAf+7lZ/l3Gla3Q5JigrhCdVCJ
kS4hBw00EMAtE+A1pCm55Nkrrl98BrIVpDblAUSMitMy4XzSm4FrgeDueWslmAAy2rHLHCBMCkre
QAsdMfAXLN7gj/IpeG6yO/4b3ZERw4wOTSG+bG5W18R7oz5WtXItW/Qx8R6k0E8E8i+ZgoTLrVJD
pIATnmgF8XgEaK0gcmD8ISs7ge/kWOvowTDn7KPy3tGv/VAcGlMy/XHDOK+aWC3l1b6XO72eq6CH
bscKiBZDrpyF9HdmiwXTZU0Rr5Jrk99tAhLqgS29Jzt9cTCKpAM9RykGScerQHfG/I79KAoLxrCq
nGBx+uZTr2VOWO7hH/xRedWDXP8GzeqUZTRbQjbg5qPoKYeE/GaDv/bzS+soD6WYhTdnbsXC9if/
Q4T93ClyyNXN9mDM+fcWWMS4ArcwY1FCI699lDW4fwbdXqWyBVSp5/GJT5PFng+70L9W8rz2J/Dm
Xf0Jetwknr0UrR4fBBwFnwc5CcKtxiL+n4Pf+GdYiJg0HzrFzqYfaeihw7/AcEFQfeRVFdHMd4Rf
tBkL0xmHOoaY3QdMRzXrbSq7P1lP5kVh0by8HpujNcOqxlUGJI4f77A4uBSpi3ttPi8yVPFISEwC
nxV6vaiaExAc3aAUMoYVGL3fFEONfdt7eFymi9E/NAdMKgTpN0iW4kf7FJvSuIeR1+P/nUuMRveK
mXSTGMdEH4X1j7mZG8x7ZY5X+duW/sANjqZfPhYLnSgie1y5nNkYjelibQrXntdQNEtLYb7oSTPf
V/zzE9I22vBO6AuP0K0M5LNb+3Y0203dhoqw48U3Lo4hLJ0sJ+Wp4VGSljzG+gz+fWrg5YMiBqWE
7uwGTYeXiDkB+d+nd57bvCTyVxaXeVL1Lzm4syQPk1NIRyxnrvqeyKd7g+iCvfYNJMhprAWdlAQv
CT+Tl6HpB+cQscSHTTc3ttdBJS1fsdnLqyGR6vkHG4Jra1/z/1DRtLpFOpbZHUCU9hxm3K+K4H+Z
zKqP6SaNuIlrHJilQpdlhDV0Bnl0YcE1PSmpAUagiazdDnRYX5210wiiZ/EhbNeqHqv9wk1/FvGd
hORlT9z6w6UN7ElsSstZZ3Frvw11PwnOkRRyP5DxZVmK+FNFtomVAkUaBIixJ4+Mgfhh2PuhcuQf
MTwfavYmagQxUfxmk85mPFBxv5zxZ81/Wo2idlcqBaHdC3pr3J+dtFCLdl/n56wuQXiUmWU9KyOn
ZaNbMigVSM/n4HhUnl07c+1P9tSMdTnPBi8sdrQ5LF5GNtXyJvb/lRBVoqYF2zXVlXjBi53uo01c
LbRgCNs9ZAZ85HTATqWUJXY3cbzMW6NdSxGYAn2WbzHMGdRtaabcixyE2866qGezcZktMAvtByek
ZymMujEQBHVhVW25d5xL7DocXWRB2ilzb3MzoN0SXxj5sr/Gav6rmeGN/ohyHY3O2nBWvJUV+FTW
ctEysYIYPpXKZwwTy8lCeCPHbF+bRU26pQP/Hv45Vrzwa6b69foGu23IatWp0+0KcrIexXB9wn8l
DytmXHi568MPsdQL0ITZSAh9zk5QGE0XuSmSzrwxVgcRopLIq+d/TpYHX7gwLpDKL/adA6SFpsai
mf0QGVPbkqRrRYIhcKy0/JeLOEc2yC/0lsioa+VRdRLnZqOtY/yhL8xyhFTGMoeKuol1VdJJw95D
rZnbDtCnbBIWkND6/swyNNkqunhwwWY+PpDRDCVWLc5fPg5leTpduNIAsA+yn+w8iTW6wWvo80wf
J3ufmj1XZTHzS42ceJu5iA/Ne2+sukOJIi61Z+DwHraJ2SuzRtK8S17ZrtZwJ1QTCK5JaSLa//bP
8BKY9cGiunRBLR7OW+166SJo6ECrE2IzfMsRxOC0YWkkB4lz2TU77hTxBlM2sTNwpB1etqQSuEvj
wbJtTTS6vhSBVml1y+ya83GETtn7AQtnTXb+WcAGS6UaZZovBwY8o/DCA8G9z7NmXl57Rgs7v8/3
ilsZ4H05E+etlAbnQKlLJ1lWRUGAetgG2qXOacBRuEkXnEVejT/ruKJzEDeKs8sehUmZhLKXabQy
34WHFwVbxsEbkjgBb35pW34FptUyq7UGiy0gyFXZeN4lmoVvul/wJZUW1ZTL9h7ajYzV5nXTDkYk
/Sj8yIYz4BJ0cTftPWDyGhXT5qCdN7YL0jfSpkYD2S8RIg9OJhV+WMYHEQtgknypNo6tl5y6v0Qi
UtGnXvt34kbr8oA35Ifl9l16SGVvyXE5s1hcZdjVxS9NTMl23O8hQrobA6wt58aC35X3XgVCrdUw
QoY2w7LPr9TZRxhOY0TbMfqxOopMwJSAOVIpcD39pGNj6uhVQHcdeWqNcmjE4y018myZlj2SvR+/
/vnIAu9Dyl/Gfj1BqQWTqJOzo/lwkXme/Grp4A01opjUH4dpgKIQM4/4TzTg6k7LIlW2bSUg01CO
OI5QCGMjHWQNoz1PSvcVpPqgqXGuZdMA+gUTO1jThWMgjDPGeMnjtFOnDyjrT1ppwo9bQpFm7Wib
TL/Lr4mV/aVemPZ4N+bQlaYmtmf8ffpyaRGbE8Tvv1JJus9WLBVwerUCTzHVZk2zVEjXzJzvwOlc
oD43e1XNtyewerU8blRFBiEEKxbAq9/zYJu7tq+zRTn2NsBh43fdIqYk0Lj9Uarg+4REPVdGMDMr
UAsk2xowhGFOHIn10cyeiCcVyJq/5oU2aMaYCTxDoEt0IzXrAIMMsaUyFwMwPDIi9NP2M2lmXZSC
tbd0U4tSKAzF16WKhFoFORANAQLP7V96MOB5nLOI1uzRrMr16FW+XkFDyeZcDN9ylO4y6jsT8hot
dt8nAGu1jrtRbpqeVnOdp4U8d7mzBwKiAalrEJQeBPvc/wuwsEgICVAMeTsD1WGEQ00VvggBWydQ
kAVcR5IVKe/y8/Mi3fAd5gOsVX5pzekO3KOZQeggBr/7snWXDspLWv5pclZsipicG6f5MhAYnTSC
03RUi+m7cLM+vCSl4eeSOwU3vhY8e7xj1idNUEvV1kJoHjKXRiUqlcmQwoU3whD0foXuXcDESfRb
nIVDuN+pT5kL6FomT5HE3a4BXjzcszjmYzJBheFafCXqbH23e10ZwByIF4kUmLDG25ESweX2X/M9
CzwOkIvgCZnMmqhp4pQseZtheHQK4UyN+EKNz7mtBQ0ObxhAM8HzQVlq1LAXFSroqItkPxZ8s01J
VQ/4TOZarH2Mtp46zwudgGbYPfwIE2e9esGudBeRGP421uBBpAHs8DVupScf6S7MqtEguOjE7yhE
D5aAzftPdYyqzT6s82p90qyXSxZHBYf5qXCrvkUzXRi8/CgzsKNzSfg5Vur0cmZgJBCmC7I1gH5l
WwkJrz4BSRcwdzcTTepO4/rxVFpVUWw93PojeGYwX0SWDnsJCQ0mCTkMAzJiDufausOzbQBbzsf4
V/ozekgL3B8KOx6HK9tdJuyoCKaktCb0GIlxxu9xVNXUOl27HHXrD0A0cvXUkS1UWPJBCJ/IxIo3
8oPnB7xPteReeMVsdoP1YN6CZKzLHLo3b748qbt+Tmtzv8f7qGBj/e6SNJc4EINZNZb2IH8OnXu0
RRuZnFehcFIXeTwW2TijRIMvgUTFq1vL/1ckddDOknErU8pioYHUCamFXeIPno3PXOpab5EmInSs
QE05z71bvstLEgpSB+N0InYbDYn+mYsB2Lxfy1Q/LR0HlKBpZu6GEAp3NeJEiYqHu6Jwl/MRfIll
g2ldUQ8Uq3ajRnaRj5SGDnCZTctWE9m/fkhH/ntQ6M+BTuxUMIJLIMHBRDb+BQDCEt4+X80dS4h4
s8CSHnNgxoXp8JYPc5qr6e7Rdwv495rFxXEH2nCopFdu61v4Tge709bRr0XiqVmgmyVeqzis/2q1
seADsWFt6yZk3EawSlEsgtBKz9h4F0NDGMf0jBAqmgFwbi8rz2QTitm+RtymXcEDXDBdFIRd8+Zq
IX6R9pFe2a6Wj6hLufX5FGQpYl2bwhttad74oxJVPL5UlnNVVV46rbVEZjraw1YkcayK0VJ143Bm
Qz+jvik4mBgzfAzlfnouqSgg6LRexU8NA4qX5IQjHON/F8OHkdzHnA72J6gzmR6V3K1o2xgvJB6z
rNvMrKuNpo28rrLWTmmXd+y1gs141nFLZ8EFhSCPLyh8+qlQqrKwtdgwQHe8a7+LbYnksT8NWbF5
EIgDmdaUbq12sPnebo7xF9nh791qup9RPup8PcH2q5v8Ejpg9g+BkECseE2z70WiWZmf7LPDhE+L
fpq066idXUaGk+jv9wgCSo0cHsyTkFKiihbkgvFFyq+O/9mrahWSO9xAn0iJvSORVS56vjccA2Kz
dda76zSyqS7ixKqhrobsOPTXe4+QgdT1jvJfNq1/+2/Gp3kkrKH8v217GKTj0n99tpPJiiUzosY7
55mMaFQmL0UB38Rw1rjgBT0nRICsbXa7WqoQ/uTprRu7yRPCJIyPUKml5VOBa3xqmrC2Bs4QLNnN
ZmMfuzs08iBL5qIuXiMu2B4BtjEMjUHnSZ57zGTak6EUkFyrgeg0Osjs6YX9/FD5s/91aeQAzyw5
s78NAYEdBkLaXjwh0vIlV0jluFh4wylA/Jw6QngkrGECa3uQuUobs1P5erUe+rN1IMqPpnk5U1kv
bB3aZrRJIzn0k4HKKsms1YurKhTaczIMvOTFX84OjU+dJ8ZdSZJ5+Am4oMkwqcm9SmKVLNsuPEDw
wiBz9dO9EHDXYDsaUf+eTLcm2dFs8E+FHiouSu5GZDpTNwTg9tcs/1JmRgIq5XbLPrXiTlAAK1k/
xBqty9YTKm39wY41QTNVvFwHTeo1apNHYeYfz9nWwdbBupU3492msJDXS075stL7rqAP8v9cHH38
Xt1AsqYhYO3CivAIu6vyEoKoX1FrHRS/+XqKRvOpryge4Gm1WXaES8prP7ZTMvSc9Q14eBS3ldcb
z/QHaIeaVeVROqG2I4i9AygPd4Iu2RCiyNgMmfg5XhdrJepm3K+FwO9x1TzeH3vKZ+5SXsUJqftm
erMzcLJPdL7wM7+0BFtLYcfDDocN55g3EPAhOk6rqClh7Yf/kFES2DCad4oY3vdUUsrgYrDDaX+R
Gm1GK3xAge6R3QlpNM4PGfjaEXrClVFqb3/ix+E4BC/rUpWdMRR9bUl0N0Wj0JXaYbnrYy+A4Kt7
olUL8MZN5wmCM9dfmPHR8hFCsMmp/ZjlkHljUYbMq+lLYcsTgxaSAdDsLTeiIxO2FVpwVqjefrl+
qUqQq1bbicGHehznUCQsN0T5xNroGAQ8J3cxcDRRUZxMCdGx6770wEHmqvcHI9mDz5x55R46NSAw
pSwxYs+/P+2gN58bMUHH9BtWzm2owLXbmit6BT5/yK+sKzrQ/Oe4qCnThUhfv67OW3wVWm0EmEv1
BmvQwXus/b/6oB4pn7lWS7z3AsucmGqbXwJEoR9kayBQqNtbZrI5ohL8YpKZEVlLlNdlS2Cw4D5r
O17gliQdHIq9baoU1/XBAt4zH+rZigoig6JIRgF9bPp4XwJ4Inxe0S0TThl7YnJDTGEGgqikBrd8
46JpaMKqhpEOfisla7sNmhCTIX3XAnj7VSCa92sSYY/Jzw1CEztNqbDDktUOsoO349/4kaLINWC8
XOM7XIx+w5CEdhnfvR6iKP5mn3SGzYFHKymNwDOHeUpU+n/WP6eM1YFS3T8mMvUe+rIaIOSQqHQM
PlJnjecH35jBNtlnLsOFmwEI1GPJQHlNRmwWFj3f3gWaSBaN23v4T7WwtXDuxbob1JXrhcruH4rE
79oyP91XBldT90Dqyr0yi/3bI2s8zQicDYQ+5QwafwA56JmXDm5yM/GB+pdm6R0cenyOkCKDDARP
KCfSjNLEtwFZZGBRygicYaN5EK9ZYYP/dkhzzGcUGjyt9UD26SwmLycw6PurqAHckTQFV+GMG5QJ
4Q2S3RJdAYWlaOGMdfFu92X2kNSiKwLVM2rhr7xfY6BjwJRbIuAFTeIcWTwuP4tJ2qLooxJ/jLrA
zfh1d6Fq9ko3Pgs6VRAx4GLQ4DAioJm0+zkVOxpxU9n1yOmZK8UVT1mY9kelYU22lw0+uZ0D3yH8
3zXz1b/M9urKTiE3T4uWnRxWodWebwJZ6SxJLTc+Agm1s1ZoiGhMv5dyItdinLbrLi6T1McucElh
MN65o4Ku+78XGBzsWkWcubg+NS9SiLlSdbQkTI4tOCsetWK3plY9EIRmlSHKs6u1qUy1GkiMbqJ8
cQAYqb1QLbDPjDpqvCSzGcfQdFXRRuUX5shjlgUdaj7iDpTYsa7MUU5M/clvWeqtAdedPolCngf9
sWiHjMFSPyXmSqXmLXn0le69wM7omKixSaFXrNSf4XkEcMWw36DI/Zm0bn2MpuiiMORCpSBO7yHS
XwkVuFfWKrv1jEPzMJsPuk0ATaXHFrEoUAOQvDSSkZYeXdJKR2+QXcp/JQkamnoCCLg4Y3/J6PIk
7X/XO0wrgtskRqcnvfHmxTtszJzD/91m5tFv2sZFo941Vg/DL4w1jVsB4AHi57fXIBUwtfdD65is
9xgxXZY3pOpwOlafXvD4VnUFkLWNtrXa6qgUtJWorxrTV9HB6iKLVtw+5ZLQgclRwq5sSWR8ol3N
y4OcT4v+H8V3Vz+WI97B0SGJAugVsRYKykg07drwQRMS1sauSuDjBxnU+7a8/KvDMCBCP3gMrYUS
V64/w1CsmnLHWSgHW7s/TRSwSteXrC6AX1lJTg272VxFk3xm8QnN/UukthePvA6hT6XP8v3s7Z3Z
x62CnXJxkhTVi0t/gL6kqRzOgWiZhcCxXVmJfHz/hRfa8tVtIsFXnJggNPEs4B6WU42/xR6FbMJM
yikrsSjVxEdGQPU0B3vTcyaSE7R8YzfBLCdaFwTMpKh5VRjbYUK6ds6PV7QYEjF3QAnNzeV+v2b1
5pLTEXuliQ0lBTdGigh63tfiDmDK/GJi3n03tXcNVBQiZeF4CTx7OqTNt4hiT1eqO5JmNhbt1/2k
VcU0ilRhQTdeeHAjvfjgBZgGh6/+0ptTf78azJ0mFvDjeCU4l780YwG//2+RXzXO6Ff/P+Eyr1x1
Nx7BFOcdP/23FIDncMZcm6097Czvl2OJ+sZffQPGJYe9HCTv2PFmgyQTVPG+1W3ahVwN8fnfW1Mz
sTETOllrUlphzrlwhR0vfP1mxXRcLVWZSOT3Y4sqI30ZHbwOnY1mYMU9P1omRHO+2LCmuaT+NM73
3PrzoenMhv/Dliy1RPEe/3czFccIYgzLCnw5+s5mRdUwTBLvbrDcEzz1Q8EpbyVnpAUVS2vI8RiG
e7nj8KY/4055e6weDOkAVSsbp20tZq0WdXm9AWCN7vFpnpUWnpCDza+s31If9Dh6miMDgHCGeJBr
tqevpm6bGQJbzneBzlsnwXMnbhbYUxMS6/2iLnHs+h5JScnEds9TwLhngBLfNIaYV4dI2yRaa9Qq
vL/mzk9g5v63ZbYKDotyyzOFf/6VtsmX0HfNdliaex4C0uboc7OTm1Rh5AXlEg3jU9vQzN8o52Ol
yl+wbRtfUo8O/3YcB8TS1B2yYwqfNfoG594CWg/HzJzvpk1izk6Hp2YVVVclhRl8no2yrRzEhVtg
Tsq7dep1qyeOTiZZkVhBVvbSh4fZY3h0/xcQ2ezjKeRTlcienEZ6sbxYeLznuFrA1cv/ychym4KU
aUs7wjifEatc4sfF5GGryV/Q/rSy7PUqS21a/AmayUEQHhMxN5UVLN8IPN8RRQ5jJNL50oz5L3Ry
bskspM4Aleu/S6uFdOHRWIfPIFv4pFmcWmLM8tG+Iv7bSr6f/kUWhZG4iYDYEMle/F6kfmq9FanN
y+JYyNZTd6p4R/yJIJ1GKNrcKww5t8r1FfUNnNd/OJTNNx7Yo/gJr/wqJmH3xsCetwV+b2Ao8y8t
KWyGP7LE814ucbo0EiRZq6eWkjwRRlpxnYpsV4qsAs0xh+wkFKlk4Dyf0TEowhp/vvAEKYfdq6um
NBtbGKKl0PgjMMPcQerNLj9ecHUr60VJsSKI+4MF72JvaTao7foJG/foKiZaTs1/75vrTPV13qLt
nilOmNAcpAaVx6jB/CmqbfHxiaQbFWGDscgFcpcemoW+0TVr6ElziA9JGsgFyAwtMCSsuxZ8Exr3
m+lz5CXkG3ChMP8ZJ0sjHEC2jY4SKVD+GA6O9J7pX2uy7o6D381dDeeMH9m+7Vty5vzSH3m5qPqB
c5GXUdyW7+t+9D5f3yE95DbSTi53PgzJoXINnJaRhocfIfS5mAm/6bHIKErUu3DeS/91Yo43fuTK
59vYu9PvfhyDvIM54DlJVg4SJSk6DRPyYFmWMsQFPgRfCgrB/o5nEhTs5shMTpAOKvEU6XL8I94w
2MwVC0w8QmkMTjU2Lk7qoHtGISE/Y+V4Z2roBiEXN/mfKoiNCUv+Dwr+ucvYHw6aZq30qB9MNAOM
tU5K4jxt5kComoOH0VRUwHGGZ3HgDtkiKI4q1MXNDrtuVZos4P23TibHZhr1LVXwRBG36WTlmjjY
U16Tuw/jU+AukCG9qJk6ijwhW2ef5uOUGg9H0jXCda6bKlHEKYYpJH8yee1Iige5SB+UKSvSV+bY
Ttv0wfTyuIacTBgpNJLHn8tT8lsmCXHV/mGV+SIeV4YVyzSjI5A0saCtfNSFoYmc18sG69BoKn4R
KWf6UyfFhJr18QPrIsWLHIbVWsCqybkoqOrY3VTQZgpFhCWVYEQnGdnOxr8iBLIVi4BSIfK7DdBY
SDaAj8JdC3nrTZ+hESLG9WtIVSYek08srs/6CQM+RhVxyvDoC8XPBEEn2KbUsxPdDkRWZ0tp2H07
hqQ1ymbfhUml4UE1KoXMZbE4gxb4NztuaPu2fNhAygyt5+rjYVOj6SVBEeDBiIr5NVeowBNU2OPY
QeB88GZz+pcp+Enr27K0gs3yb6eG0ptH5uSD/o5tN+5OPgKa4XT9BVdC5ta+cw0l3C7sFhm8DERj
QiVcrlKtbyGIpIFiE4MQHsFC+tb61M+fyhO0RkZHLcvp8uNI0DWxKwpJKb4Qt13/rHQfC9oRG0hM
Wjzn49Jtx7BflfLznA4ylvi/kZviGbZUoPLXPZf4BulCuhBOVdQ1NEfUHEQkRrHUlDEytYbPTgBm
WKAhxIgKTNtVy+YYITFup57my2mIQego+FPI7jpoT33a7MNbNdi3ZF8YI9i9QKJVO4Z1UljBZzfp
55G0aEp8aT6iTiU8zBzxZiEh4dJuDks5mcQ3kq2u2adgJKkUehXqlqMb6T2c/RtDrLNeWt8/gL15
SAKGTykEbnqnHyhCrVxXErPErY2mEeFTidxoYXDH3ZqEsyaIlUEz7MKqcmjwXdflxCsjR5GPfyHS
1WKjwyMewFG28nRP2nUCrvrw14AelL/4sCQ71ssophm54ZyRLOmFtNJYuxWw3nqbXED1J6lqyONW
nIPxeTcQ14Vu7qNBQrlfxe5uJjfbI4xlo90rVkRVhH+iTL9Z0hjOAqeifdsDNB25k1qyMBaMdHH1
PRrbHcgUgwQBabEAsMih8/MVIF6rpCHFKItiHNO+yA/14IjMV+hfK5FGS243wAzmfW7/0RkNw11U
tDPK62ZyX/cLVztjPbrchrvcMpYfEV0dp4s1HBGFiT0ZECtUaDAOdy5kD3t+qCb3j95NnKvfK9YQ
mpon6nkecLSE75PhNKJ2CEAvhYnXHnCAnyOoN2AX4I/YDy66fm4ufGrWFhtnSqXTLbb606QMfLd/
HpzjIHL9A0rJMBD1O8q1J9ZhfWpBeR2O5XuetmbwRMu3Mov45BoceaGmWqC+YSmv5S6l04qb4jzK
C3J0/NzLRRNjCZHDwVuiCfWyUPWlXMvdGcS1swpkOxwUqoIXIzW24Flr8K8N/1wU4GrU6ZB4kyDe
z0vIHoRSgFTnoXekCc4+6QPa8BXJKeJVqdy4Vc8vLfQIXel+a0ZT+l72OoCP0PFi3IslUdIcBRJ8
BY5SPF9yOQgMqfY8Ai7SVkwGhhWeVbbm4jsFUyV89DBQSeb1FUEfWD/+WxJ0ocvwqQkaPRd7pyz6
A+YJIc7wnsKnUPsGqRDqjY3qX+Kiosqm/ljRWrN3KWIc/3ZDRmdN76L/ZfBycBh/WEspknfTkcO1
vraLd3wBa0Okw4WDyRVIS8AAQ7XTZL9yEJsEp0BUrKQMHQk0hNqTQ2mjLN1ulZRXpOLdwWXOcqlt
aIy3KxuejKcnsvFqf8jKh8GBXUcFAUUMrelM40pRDC+q+0Tx93I0DhvJZMZ6I9bqSGkTRMNnaAQ2
+b2rL5uRPk5mCQHs8UU63otQRFPQu3rHrnW6xFck3xq3PqMBJNFAmQI6dgf/D5gVM3E2G4FTnisk
uDRN2n3OvJeiQSldq2GngCTpYzNj2mIRkTb/cE1kPnBSj2ONXGGvYtoULjVxx8yY35oZHjA9QuYo
UIlMvucDV0ve+GzS+8veef3XQMGJBBBZqeTGXhzssmADG8nVkDU3mP/CR3JVNZhM0qvNfC0XLogG
0+guoL/eVSvarIWBGENXIzKuYGtJtIKw9XBTiX8E1mzDUCy1f8XxB5hk4tGMGrnNsYN4WsGi+S5m
ocp1YQ+w0/uryP0slGqNgOf/+Xr8rJxKUvtMmp1zrJ1/NrgkQNYjdCpE/+FV9OsBezgT4ujDtSsc
+7vv4n6gEQJMU6nVPTd0wrW9HudVXiZskr4L/2lwqMZEkpcFT/LS1wsaSJgE9jXdk/enY0z/CN+B
JtRYVPvn2DK8HjODK9cg+kqbM4YYkSinZR6ySTFo/ocZcrLq9ej/lHB2gJ2P7vcnh7wA8JmECVhC
Ge8ubA9Nw+n0efr5ooLNWwJcyBqUHyPLdscc3IWSnmqnbtxBZE6/yK2mR46mADIeGlTEKqd5fhav
1Kw4DgXmuKzY0WAtqitaODAhSjT2SbY83ganDTjoa14NyxrcGkjHMUf/vKCajnJjXbz7KitKnffc
9Pv1kounP7Dz5gfeN1vaiDWskGo/8vfU+mI2YccS2NzMzu3Z1sKKKjAli7F8HYGBv+kvndDa0anv
8v6wSYkHrcFATiTq8mnYfd2+bR9mw4yKl+NVzeW1DgymY/XHBsPtwNvADMMjD6CFr3aDAlIPzrve
PUvGP3vro09RUfdmOe8NNw/RsLCXWhddWUhuZ7vX3BWyMVji5vTNKSbhC8virIv+YNuvBCnC9NnL
b5HMSk+4miTMa22/02+qUt+osALHGVX48npSywwk0itdc9X0OYS9o6T6ecRx1zMQ51b5s3djc+G7
2ExhRdiql2DflKlMesrv4/YRTo5bm0JUAJWZxNweyDj3JBrSQR3rZGG943+fmGOTlPG8ilKYjSkd
+eXClnSIABl9Jkcc3Da2klZ/py6fe/KOheK2PWbLRil0nrApZUa3s5uYRds55j09DA3/gbWxDZ+E
k6sn337ZZAEX7XNvFLMw/q9e9jepu+QogZcLnrygGjH4MQ7w8iHgFENXtlxxXJbdBnf2BE2IUnyY
04CJ7kbEzN+pW8xsTrPZJG2KQwp/5cYekIgtN4kiPAAc41VxUopu9FPSr1fqhhdbNnnQcxQKNZr1
WgZW6mvi3qEneBpE+Jhgd9KV8t+18kcsggWgMqh9heUgNIEXyfH8eq3j0MqVJ5DVBZcwn7lyCJkj
TlEjPDRwKIgpVVjiqufV9NAo05d62PsKlF/esTx6h6uEXRyWB74ZS5wBxhpEfr1sOTfHOzXQhNlW
i39MQxfrq/gTAEcMmbMSfjbCcsGs2f6smhtdQh8VgzAC3wWzf7vzKwhMDfe8Z3o2ay5BUolKf7Z/
XSeWC8Vm9uZDPyBWuBqzmz7W9mBt+uQgbsn1UY7iGhjRwUh2qHPTrloFEXZTwefUj6/nhOvFiMxn
P+WST0CBzNc5qpBnDgzmItO3w1EQK1c31kktqrjtXW6sSSuUCz0yhpPr63tkzleGgRenvEQTUCVi
j/5Gc8I0kAno2vG83yjdeVoTb/+FN5q7SlFj7TtARZ/c2YwarbR++aIa1dnqK/Z0ntlyYdc7Dzsv
BeShic67JUBp4RL76sBhUO3de8s3djjs7gHGyiOVZgqfzHf2443R/W5+T3Sxpgj3VI3DYz9UjXHK
27EkahxvDKLBn93wvSv/3fSn6DoqadgxJVRo2IPC+7R5YO20EdMSDXXUxE/tqudKZOjex3Up0ICJ
Fg8eSgx0Ancuty/og6/zKgBASZJR8UIwSx/POb66WQvah4w6bCT9qOTEXaGRScmB6CK2ZSzFZKck
CY/r8k4/CYLilNEwfrW1SGVfOICKqRVXtEXgbkLQQfOYJ7WlAM2xOly4gSSmnsaXXJUeRBi1MkZX
ICxpsucQSLd/zkvyJk5lsWRbjtrbdc7tsRmECb53GGNPP4eSBofhtZ2OG28qtjbVC0T6KjZ5bTeW
potxrBsLWFnK+XytITRdArR+X+TM7GJ0b2o+0aSBGpSt0KM8udrxb4M3Ks7KbUbPz7cVeIkYF6if
SJfSU37CcHNE1spAf2NqS1MPbJviX6o9AK8qmZYaNb4/4pqmsn9f/7p1PbXPIfucRPpaC4aDRoig
jQuoU6RNoENSqRgsuNXrQgelNxRGPwgoaVnje7T1/0x6JKWl+HT1qnYcJhCChZS5qmb4LF+Dhq8X
772sPTW5RiCWP7I5DyOrTn/J/hP2m9lluQqfi4UnkLmCT2i2FkZ5jQjhrHdFQgEAAjQzXZVVkM6o
XRSy5G21++fmc7IKBxo8A9HZbQTrxo9Q4BQsCO7GA2mwhvY50Pp1yht7pTabV2Cr+IPooUryhpDq
x2Bbki/Ao7z5DtXu/0L4nbIzOwJy50//VA5GB9fsDIZHTprmSBCu/DFZfJ0l3slsCjcwhKzNnTAk
zb9VOOP0jkYYfd5wdQ6lrCo50jPJCMG/zEHw5DNNXaLebqtP8JCABm4YGFyhOyesiIYghAkR9gG4
PiYbep2QCzfH1HLb7sbT2SipsqyZJgmuhhsBGSykmiRLU8gyfC9T4CCD5iAC4Jvh8jbwF0L3KoEf
Ya8z+MRcVuH8IbFb8CWTUbbs+jA6rHamGKAIQL6jX/ih6aW5KFDilORwszwPwD+ZobiYeL4slktu
hW9N1p12auqB+/3QHSJw6Chc1bBm+cyECtehNX8p/f0a5+ScpmWtPh5+6hp3UnXavH/L/tJgejFZ
ZhYqnTHcWQDftEY5y/06OL3pevnljLRC7FPxDr/9XL0xr5GjwJ8d2LoZJFudpvXAYj43GIoATYmW
zfWIgPPduv4SgABaUYwh7c2Pd3GdyH2S5myIvVtVwBvcGZ/v94mml3zaZUDU69L5janAFmuXPLpj
OOTb9HHBk4xLdGDt3sq8RYif+jKb0zf/owQjIB9tkTMawinNAHESgL1wiGBzB/FYl+wNjF9ZEitG
MG7kFMXd5b4QfHvHZs3+qOvcCM6FsO4Ne498NETgQRsjZixinrw6UumHpogkwWS8SB7jCH8yHv/v
a68ckqj0DC03bhgdpKhuo7P1dYyOJjfzcL0oTHlKqfNjcWPkrhaNkNV/NYIeV5MXBiNBVlqiZmGd
n8r4yjyqZEoxucO6X65mgyKxQ96mufKfj9JPAUGqr8Uq12x8uAQCWXMlyvQH2iZEB4UdJZfbUSa4
EbQngK18mrP4ukMDXS6hr+QrmiQEXfG4q35fGo98tVVxTzC1484qgdFq+vpEwFffLoi/e841NMVf
IgQzdYQn6ye91iBA8GJrDnp1fFH6Pn1pe6GFA8nTOQd0/0Pd27akVbRFCrzfQeIqz630Aa8nZS27
bZEh3k54FxLWFYpgrFttXUpUKhejk3xUdvpvCsliz1efXrFh0TemteU0RgsuqFrKIOnGicu53P44
ogh07pW2shXFe8oRxAvExri4SFVBE4hIzk8agjsDHHGkybHkMAP32j0zbkykfdv8wl6QlPhm9x4+
AoUG61c0AkLdbLZFva9afN4biD3NNDikUs6cSG6X8qtjMuuS/CY3Q2zZ4MeuVMRqwzwC/UVwkktN
H2eLaswIHPBx41umc34oru0Rzedt6gc0HL1SR/QO3vqm7Q4r0OBwF+vxZaAjvtDgoDB+F4ETPwJ0
8iS3S4o7gpKoDrMvID4qRMqFlBBH9DFHxB33C3Hfe82CF1pjo5WTjziOfLx+6bgYZK9mu6ViW00t
9NOv/68S8m5kjMM7wpK9Owm4JqlvrYRx6q3Jcr99Tr34VurQUzYUSo+vC3er4RyoewHDFvpJhkOA
18pEHvH+7qGYXihJw3crk0YgwJ2F2nHdqfEPb6mJWD2ptuiTWilRmHLRozWtUriuHEfjk9+9Yjyu
4Gj9jOyVNtD8KUX1/g/BP58d/BMZ/HWLoy7cyuKYed+BobNddT6V+i97DBCfmqAVG1RxDS2hET8P
jz31bRPR7D9Du9oJS+2CCSL2AoZTIvKQuuFNdcwU3E2rGFpgI39B9qe48QWPP6O2xOk9K7qiSIoR
NgS0r7KZi5R28mYkdjWy60WJszMe9NWHicvDm0VbBfWKik0JfOJGLUoT4sHaHjsvswMMkci2qKrQ
DUtoPWPV9KlSmRFPxkecuIDFFdnYhBK+OGmreuf/0AM8Hsllg1T9Dr6JAyKyEEUP3EEMtKiC5jtf
fQSAUSEuPQYP1H5JOrd3fPqo12pSqDfszybd6uZ0Ob1Fv95iCukpEHlFt2HmyurE5pDux5GIGNHE
Od/+stjjRImVsBGQNtgQfMvT1VlqBWau1c9XBR+94XplgDPHkBKRhb4KSCj6zCyJd0Rz16K6rlqy
zDvV/kkVjL5y9wPUAl/aWmvqQOxJriy9s8r/pWw12DSVhBJoYxPVfbcMACyLbirAmxDsSs5KyjKh
uibnqTdf2C5+3eMuGDhYljPxw8qHUhROIlljPnF0UrBJ1hF3w2n/MNEfoY1AWTzP4ftw2BUoWC/r
cHp/O1Z1PsliqeuIfOSjixn1NONMC1qJkNMWq4kY6KJ+l60ibvqizGZQcwgK08zwf/hQt3epmlil
DVW2eIWR4v4HLOSoPaOA2TA9wk80d9RYzQfUtJSy1ARg52EYoy542Z9BGMica3/AwTiUnDRLMUz/
nPMxVUljBzUx/GABbnf4JtR4FS4qBgbeuaJboKn/RvEvHXgEn+OMj0V01OuDwfMrbGa30WqxXqYC
mzM8/ZMqHzUYMoQ/bXKINvTgDpXPDipMKx0H5m5YMZU0+kmU/Gka48mMz0eqiVOLjev6ZpwfhAl9
37MTk9cJFyarftgGmZprKkLAS1C5XKnk2vEQziHXTmp0jl52yg7Et9Mq56GnIehgLgjDqqyYuO7D
2ZkmHdmfFXo3Rhejc9R3g4PUvHZ58/FUubda8sktDHJKQn0G0zBH2BKUFDmzWmP87QUc9FQ4utv4
Y9r5uS7bf75rhON6o/HKh8FE0wUCcaFLeLi6mx9FbstNkt8HqwtRkfROoWw/MPrynCE3/ROUpw0u
H5QaghZQAYoFKtjwwhTEPYGSce+Lb9udo3P91rqirGj5OeBvs5qMImiKoWGDZlh/7QpnXX8LYvAu
+BMN7fXGTOBrhdfMIrMV3XVntGPDdKeacqxT1db7rCPdUO8riDlETsYvY3Cvy5WReGaRiN6SOXBO
FlN2OSfpPKZqDOMjr+NYI7WYyKXrNpZAxMYjfoWI/bOi8+JRWA5ighxjAQ81lQwO2+QHqM5Vt2Wb
1rwspXKi1CgQP8GuG3WHEYCmfcMvr9sTjUiy2ZBPwa0gRb29NAzoZ6RP6kYc4nljrFqhV1jmwAOK
yMtHIF/Pb2gDW1rajbvH6h4bLrZSoGnhOuIF5fMNyuNhb1EP7Hsn/q6P/6AtPQJDUHwXQeK5C+mK
Ycvxt7jwVEscgYIveaQHxiSs3yL6RX7eC0L9ONxRW6Q9zDqbwYUQDfvLaT6AwfvP1m/WkMu64buO
q8znny91BODqVB0p+v/awaGWapqexXwo/dQxW+f9QFjDcrnxhSevHVHwy20+DzyoLSQ9skt9weRv
M4M0Xdy+LmhmfnCJHlLUmJ77QL2fEV5kmwE6maW5vJL53vU1MXIWTtct7q+ntzOG8wQIqqeiLZIF
DNdH896Vz/sWYqlDrf1c4TT1yYBmKRPw44GDBm6brA+Thv8lFiyckdsKPY8/clTQJPJ4y+L9+LXY
wg4PjObBOwT025jqrMpp94PW3PbFJwTCXbcWJX3Dy9cXoPPNHlkvfHO9lxOOPYUXeqGwNwc/yrmy
ABe4+jYHOWyvqVxE/x7jc8h/sfMhp8G5/rn056H369MORCqk2KV+hF8cyMm3WTJWD/1N+AEa2VsY
kKvPly76Y6BIsiwjy3UXAR6jvUhP/SuQCbPTOgL4iHZQr2O0aO/8GC4vlqROnmh5g3Q7yVIa8bDh
a4T8JCKMmoNWgsER8ggCcvwnYedvL64Xf++DNwnMPCcrKHEpsPFlR4wQ4N0UxWk8cGKEUZ4Zs+oF
6UWrqtjNH/FHU/SE527E50fOxt7B9t/jBwMCAZOtIL5lMIwXwtsauHACbTsonbfBILE3SylmGowV
BnofijvP8PPuFcWMNqA/s/+uqe6/X5PfD9E/4lPXQyOOIYSCZMtzTLsvZ7xo4Vmgr6pUXr27mD4E
JJA8Cisj826kAOQFyO1FB5eROU3wGmcSbPHQhX1l/xqpSXLkG8f7FQzIPRLZZY8CyE0G50mzjIgZ
b6+6r+VzkD8/u6O4aRPrg5TBiI7Zfi2ADLn0M9NSxbwZqh49aZGl8M5Z+FOLTW+LDzvWGv78iEqv
IYYk202o5HaU5mvf2hTnuChEL5KTHWrxW/xfayS1oUcHcI/jFWHZqFS1y3O3KNl7G/rgexy0kzYP
Ehwk298CURObAFUGKteOuRI4nIwfgMpeRhLAPOKUuPpsnJTmeidstDx0R+H3JBu2EXEndgkZ0rwC
BCOTQa4J09raI6Jskt/TJjLYwrZyecWfhcorQS9AqCKIgfch7rld1AYdcYCzG+DiU0Ih03DOIdvv
pNEnPIsTSvUMxPzlimQDZIpn/AtLZmg2eAWsAEjGQAToEjYdwXHKHIiG0eafe4Eyrrnz8uvslYhy
KM9Pjclfs28jCUSP8w1YI+Wn5oHjaT4nTMxFm1V/UXrEFP8TLsMFYm1w+CmHAD0aozuKClGmPLas
LmfNlEpuKewXYgswzZ+5IX8D/tfb9Blm5aML56JXY/Ax+F3QZhVjOmlioGJSS1FYF29rLRTt+wE4
Pwowtfz8rgijrQ7GnMELAkvzJjV3trMVgb/cWpjoqgMaN3Ik4uoGf7am3qXMCncI1hyJGLwnkb5r
CXxGY62+Xs1qiSHcRawHtOnctI/GgzsTHBz/Ow3oBbwX+LGcckb8tzWRg9f63oQKw6X5dnspu7VM
XbDDgGYbtIWr8xFH80DG4TSEdTh6vvgTwfseF2xBCHzj3+WOTlm2i1mbPHSdkRPogIQ6bEo2itc9
JpNJqwg6+cb7Qj/fsCrK/WrVtCGu6LN3+uf9ELaYiNtKUFJq27WdG12zZCMpaiGmDNxIEG7m83ge
Gf4IKasim5PseWgNulRPmUePt+sxPKn8EynoIoH5EJwCBEpa77TNS/ET3zeWhUaik0zPf3KNQkvQ
cAWRPt/A42OMAXh6RlD2/Yp+fd2VEMrfWdCPVYMjvOBFBRrWlGtmg/yWpOoyZi58UOd0s8y0SHnl
20FpRAKORBhufyNLgTr1NHRfV1JcVEBzpdWpcMYLbeVP69FPRkvi5LlyW5egvhiayP5K+mScQkqc
uXnwNgPM5+4KXGWI5W1Z1A5VD+1pwoCZrvwjmZVQN6I3pr0GVWPy8kkgOO1R3iPPUjKYW4m4wyhh
Wdk3BHUYSmjxflDGM9NreuSDfVYdnlPy4hu3GhcTEISz6nQKRLHn9vZBJn6268lV2s7PAwMqKeFj
ko342eTg/3zbpONz21EOangZ8rFGanuQ3NLOC8zuVzHcYxarUwt0e463E6dDsJovMhdfsx9gJ1Zs
xY2n74urM0vSjvp9jAjiSnVgheWAW7EtHW3l71r15Xe2O8KGL0Fzxfek2xGbq5LbJAsPfjmVMVyr
JV8/eWgdUWwF2YMuOHOYZUDllb5zZQpUDtQYsptpM3pa4vlI81Mz2g5HKsU61R/HkGQFL+cMqgUO
o2PPAw2dI5UeLM49ChHRpc20f5eKl3FcI7GQgF4lEZXeuXt783utpEyAoQF/PJED7ZBYfO69yKLP
kPLNIpdRZp9qdrgMZTXKAmdlA8tXWL/n7z0Qr04rNrLVoasPF4d9aycbI7catm5/vdKvdwj8eQCF
cN3NXAgrn2/jMMIq8XI4NXylMqkkWzpAObD5drjla2KPcX+lvk0D0qDgI8/DxwrbN2HPsSQJhwCC
Ks+fNy/A8t0Tgw+tRhkKWE6rIQakHXHT3b9jP6vbIoVqvWqKlKPJl6dcZUpIoVxwVKAub6m1GyJh
wt+RTBwzv8jZbxG4VhhUGDoNg+Iov+oLHOtAs14z0C0DQHVuHY4MJNSljO63hFvmmivcUCMv3f+G
62NnZ275Q/mE6x8qpXeZYIitLQPwV8gLdfSG0dc9F9qACVC2CWNLfzLSwLSjkR2RLpFWc5gaz3fB
jFSIcTbKaKBehyyq2Q2etqdfV/0DSv9ndAZJ0P+ckihAU3tlj9vg1JzqtlvcmiX09XiBkFUw+ZEf
9hDhke6iPhJhoaYR4OnUawM+UfvLp1uxLSOEKGv6LEo///Zsm7YOuJN6iFHmUr0XVQB3PemNwLEP
VDrb23aieEVd0tl6yIxhu/8oVQGgyqHFS+4IURaHWbSfc7j/wUAUaN38LkYnXqJVyC7pC2OZgabH
io+AqiFLZ1eyRlUK/tOIKt0k63AYuGYuIDXIELVL/azC3AghHuNtgkWNlmI0TnC23kPExtGCNZ6a
ADCoHzN4ho6KGzjzvB0jAybqfU20FUGnuCN2SMD74KxqmyRq7YS/texIfOrHuHd4LrdXmFxM0F3Q
Hjwnm0g3ukLJK5HCHXgxz/Fwvk5Z92k9Ul/P6aVhP5o9AZcIXdk2EUC2kcAqxjhO/10jCtqctvUb
pBfie76LuSAhj6whNWJIOiMwjXhMj0oofi/mrr26Vt4duvLiMKiNdDyKiyt5oO8Qe3wXSEXw3Luz
9kwJBCk5brzQNCp2psHdyYUUFRd62be0sYfml3u144rFBvMJrfk0gOei3GdZMNyKOzkoHBom2HLU
l/RSx+qKLXpYRF/ClKE7Joqem9P15FhOSDbFAzqMyXSazurI78k+35XVQYWqRAOzNjSDI8LiPdSV
AmxqXx+VBfRM41PI+XJSxjA+iKhabqIUxOG7JKI1hRypPhwZjsR/ZlbBIzYKqgjBKPPkXMb1qyOB
8SKrMHIiBDaW7EeilKFJu7eAiFEgKfKItITvHfPhjnX0oDaODynF7T9YKrqZYSk15uozUBwgMfmd
9ED1Mepcp/F4u2UM3RhgeJ7msAdy/dtfOzem5FWe91FZgkajycKcbNwmEc+zmY4fSJQAb1IWAGRZ
+qOPmsPuYaWxJ3YIvFEmqTm+7fReEPXiILng9GzzXkoO7vWuo+21sH2CPjtkfMsSqvaMHGJxhIV7
VLyifGlF2+KmjyTXHaYEcORTh0OVhQgvUvjzb8V33wiu/alOYiUlN83xEuKKTYeNUnTfaf2cMWKb
oS0SEZNFYubalLgBFwCod6eXeimFs91FgtmOfU3gEhUzLqQWaRVwBKiXuuaFzkn7FhL9E3TOFnOu
t/Gt5vnBjic2jC0jDH9tK0uZq13+qYj+XZp8xvwDc6C/Vq8zeNTIJwGs0fy3dX0cTfP2vnDzRdwp
BeN8svx9rqjA0dR5ezwk2ppU07AiY8tADXa7zklX1f8U4fMhmtUqdvb/eYKdvrT1+0IzPTqCDALm
peSsZq6fHlQkAqV12BwPpEakFNdiI246X/1NgDKqCivyFW6g4b0d1xG7aheH1qbffpPZLU1JSFdy
9CZccSHqLr0w1YiZGGIZIsoXxQoPflwDNpSm+cwx1u7gl1jZ+cL34vJLMGK5s9QltxI/mz61LdaF
HqEYkI9q8Rvs29z+lLu4aJrb0oeB03Jh/lqO104EOwrjEEKtBH+4TlbHyjNts4PGd7/DD5dgZG13
jzBMJkCzsPoWmC/pYGxUBmsgaJBK9/l5p5Hy1XDf18yEgRhBdn+vjQuvoJeLhNuZ30IYErnvqg7O
uv9x/XF5696Ea0wXAok0XyzF4wjdBCBluZyCmYTv1i4qfbZvzeVE0nKZ+nQIAVp/P/MWudohW81o
nrG3W4/KRrxwtRUFzX8u8BI0pUFjDIjq5owrjc2PpxNh34ccU2uEFvu9qQzeKfsiFAam1rqVx6NP
Qi66e5/1EcIxuZre04HkZCLby9AoJyfranQAkQOCUq8zKxX97linV7m3YnC08vnf8T3Eqx1UJRUz
IbZQEt/Af0dZs8jopOnQVLYjo4gySbzjgeTUX4DiW+GB/hiM5sfs3Ecjn1DkZUn+bjJFxy/xpDoc
kV6kzqFPG2OXmaAtMUGTAve16HBn34F0GG7Ts4jP9iGkQbw29ZoIEAZrR+4qKxVX+T65C7xY8CFw
2mxKvJNr9mhZhfCuiUx/6wKVZxoFu5wdQA+oSXXyfF7YxvpVkwsmVZwL5leoWMwJJT/msJIRR5d2
o9Tcir5bopCKLeDBQ3hVh7BAX8W391IaOF9Kh0QnqZvI6MPYRshl7wRGFPZjzONE6gCb1ezyV9kw
931mukL96AwoNKRqRnWI19ypFgmMUTCIvjs9UeQyQfHS6AfxgD53nI0hdN2grqjcyW3XOLW1/6HX
wGikZ3nfT7xVG2Vx3uu+mgTisO1FQMHoMIyqe2cXR2eC3nuGPDMZk9kDJeVmCTRgqX5XvvXnHfg/
MZBb+DWLSqMPuyef0o35Ora0ojM8YKl5kg0xXDEW/OnhE4qNW2OEnzi/dIoQ4ZjfSDtf9sqVhiQk
iZmOUWFWav43uYLqlpLUGDYQU+dX5YtxtIbtZssXcecWClMr15ne/pSwUHa5WMLmwPSis6D/qxbm
74KutNL7eDunzeaVvqs29qFr6dPlhJ3+E77tH0td7i2AeoxbiU3PaG+xT8xm8ZEDOP84V2Afgctr
R39bq/mA1l29T4geJZRg28H3HxQbX1STKJtRU2QtC/Qk/8lF41jhFl6DJE2MBVV5lQkcR81wdmHb
5El455hpGVaUElFo8LwwwoPHAPbTRoqKXguazRA8WYNG2hNbSALTLeRWL7y4shefIFLX/ij8BmFD
y12VL6qG9OwryDCUFinfsr3sdtdQgd8u7PYPROIiojXfCdfhtgEdM9XKKuVSF7ZjtUox0EpuaLnU
VjXsXi4grDw93FD7eX8p3lcGxVYHyaf0+3CeypMJ751zvsJyzJpBevmVnqz0nhISp8yM0Xuu7vhL
pndzwozSjlRCocCNaiAWRITG1eKGo8dUhPMFAItqt/9mMJu1ompM1O7yQQIRPrzfzBvivgLu/+wO
18vlTsPI8hKY9cek/AOCpKzqttvqANkNZvTnitjiyYRrmKH+AZrqVGBtNGabstIq4GgPF9lKC1Ng
rr7XitGu8xU6DuF+2ozzfP5/u8H2Q6O2YK4ew98V30rimJtUmx73gNVVvG2sEPopTpy9aMso7wAm
WD0L/vQtX7481kQ1jHu3GwYTg5uB6RL5LX4wr9JLXogwX77Yn7M63SuN6YLSK+qKdinH+eM3bl8Z
xFXpiqo27vXXshN56LJGbWki9LBQkqGFqcAOvK7SHmP1JXm22cZkwJNitEAfTJFsKhKM5q4TnxR7
GEjuhvyahAZPm0ElUNRRpSQyIi29DGl+VFtrzDn3s3EZiOT3Qr+dFH6CKWRLhVY4yBIi7AniEE6c
E8jgG1zaV1E3fcs6eJPfwwqFnh3tNH58pi1c0QsqjkpNbcqXMoDWNWNNfpu64Z1ADqgHKz0UhgKQ
FRN0/d7tJ+UVx+sn2PknY7JPpzyruotIeUnKLtBQ/yWT1g98F1fhcHDk+B1XNy5JhWXIqnUv6OBe
jtYQ1/CEN2jXb9IrspN9ks9L+7TIIeWUBakb8i1rISEo+NSB3l1ScI234zsVfu/9AD4/MCEIlGUS
YkbQfE3aw3yPXfDs0Q5N/F1QS/Xl5S06GizJNU0S6c99svBSSHfsdeCoFXK0Hm1BQmP937340X2k
1TP5wxVjgBXvcPxgdi3zSxQDMJ/PexBuyOYsMu3UK0/LfMFg67/FwwBDjyOt0AYPZCeXQTXZVwxz
+KuAZUsld1fnV/tRcsofewkpOWIXbrNbTpZz39bksYYSEwk8ODXPSmL2mmVNsBZs3LwHhxf9fhma
k2bDClqpMSDI0xndy7FHNCzpLFDfJnLygaSDSd0JdCE4x15SuIYEznZtXyggKRQKOEU3PfQUbsQi
mwq0TC67pldDQoHvPUKpSdsZm8O11v3LmBM1zxAqOdRAH0dOWGzwkIq6nhfDHKxOjC7KXixkMIjl
RTTXrUdKqK9I1RLqh1zNuInbXvm6QWtjp6O+dd0+a5DfSCmDJefpJf2sDxQDBRsJ1BHVO0FNUEc+
7fyi8vNvVXiw9cGyOXZ8HNPgkeFm3zwQOJX0YylwRFr1uHQb218ScQlykc4BvcSPMo0QCgGjI0XV
bdGARz2GVZQ6t5+XLF8kBlWcNuwBiu6+f+7+yfyZiF0HMszJb6Zd0J36Ic2E0VuxE2hHCRE66/9J
vAR1JvY0qUdzSv4FGcSMAXSV79kxOsHpQtDZp+oiRIMKkShfFOHPkkB1FHrROIIR14bCDl5y8MQq
AqKKb0RF6EFMPwA40Q0oIV0NbsVd+EFhfU+bpWqcGXhLbUKZfIZkxtAnyAiDtXqv1ayE3QtEoQjT
6q8h1SRMuxZvGzr4eXqeEUQnrxFbVZf1POUH2ZiAjGzkFEtNLfUtNXmnz7vY/Wirzt+xKGX9z6Sy
IZTZxhmJAB6fxhEcawSR9J5qAv2QHKwGB8wftXCSKfd5Ugwyvm6e0joJcD6R11RwjMcaDXayRzpb
CeSzB1FPPmjZZ+2tj1M4d8vM68Dh+66f0dvTRSnXP0GmTBroUDwQfKNVG9iG5FYn37Y52xGw1LmD
Ra8+dSIy+x9IFWL+8AgIXkveBQecgjoHFIJxQvwDN/uzqxGoEI8DGSlEFa4XOZrLogDnBNdGl/mM
O67Z//yjVvJYYYrto7WKvWAI4WuSr0BxTLg9VXIgjt6XMa+0a/ZJF1mIe8Aia2vzEE0SM4Hhny04
x9dkt7eJ6Qn8w8BoPl3PYalkgNQbXuYL7eldtW51nCZ21s59IR1LzW3+rn1RUIXMBRWEzfLJ41pk
RNMIYnLim/ICGDhS6Dv5aYXKU/Zic24eCcqjOWycX0+miZQnDViM4XQ+N3ehiFgfDL6foWFG66uJ
O2Sj5OW+hzipwo+ejRhVlQU/jVYrV6D2kJiOjFjDxdPwYCO0tz8Jmwb+Ud4zyZA9i+yi4QSy74K6
EiE/kjFQBKKmVRuyc/UCoDSvcNxmFDCZn5dADECEFVgD2MsCf4TpdubnaNKf/PSmvyomX9Jbk36f
NGrz5zLhwDsBGplVQPcYjw/qHvjvwZOQVLHE/awINScjuqrSCRmrn1yQullZntnimfKGKMyHqjCQ
89/6ZReRocrdd+SjqKz5UbDU5taJWKX/X5lg2PDQCl0Tn8+Ykd8qhP5qvTzUX3jhwQjmMObpbQqs
NDsepHw2PL2wq8HKp4qBCpmwr2imBHrbEhS/cWkqckbQb96+iY2wZ/U9qgDa8Azm6O384UsUhU90
QG8fL3rLw7j21DigughVxZwXjzCXxwVeyws1eULPx1mq2AOlVr5sguAEXhOw7uFOoWMmbVvV/JtN
sy5ZA9UWnj6QMQpeDlIj4IedsuZyWtoy8cl1FbcKlyC30Ucb8d+RoX0+QeCfPlU23BfBgLMIdpSw
HjLWxvS8qyyC8FxouOuJmqg190WQ5c0XJZpUlF6yOiJ8OxSDVEbFrnRVN8OXRKy/zVgmRf6ctxA5
jhQN3LI75EsbG3C4VkO0BJkH1lkU1x+taSnnxOECfRNIuLFz0Tn66xE58iREg84Zs/LGJQzUIESl
oAp1Viei0qTWxjt9AqCGuCJV5ka3bPSGRoCefkDb3Mfg8DRPJ0aZEfz7peYKpEU3cQfbTIR/YisG
Sf8C3JmlhbvUhxMjig1wtxXdKKY6NVRlr6r2A/2Slqm3VYrcucSdpsjE86sAECVXG/d8dNAArt2D
zt+drTl+lAJgmhICfYOstIYIsWYxK73btbeNmEJZIXpihtLz1LLGHEzw58B6VYCHqZqm0DYHBdui
EbFu5aFDtqevGaMG1ZRtpdNbUL8+wJ6SI67UPBKQD2VNiWBGARVSDZ/XiMN6NZo+ahMi3moG5I4N
LxQHdA7rEek284fX+KI4Bn8NG5hF8ZU+QhwlmYitxBELhBsI+gsfoZ+ADGmwILYdGTngzLZie4EF
jaYl3hGahySh4l0mhE3WdfsNMANqGw0r2lxOCxFWAXIzlmxA+qg5PQu87lltfT+RSTU4AwYxGCIe
tsd41I8cKJUI+iO0k4VyT//x/gpF0JBZeNgLoDbrnenhpmuXLMvJklOqtoqkNGnbheGW6pg5fxkc
YFfl2sQBUfVgTPtmhqbQCvEiUJt2w6vFcEy4QahyCTXZHr+Zpk+V5bugy16T+4H7YEjipr4Bc3I1
q6PmOa5TXQJCA44P5Nw6or1pKu1zLkvC/4af4TaCHEVDTjs9BqmLIY8Uyy8t+O7a8PFUFHloDuab
NfLfJKuQjSWS8v0Cw09d/JOAtp/nPXam+sIYGU5LvMz0mPSqP4KgX0WRbk3ERZNdXYncU5WGxI5b
YXB3Oc31AcGY05T9Fr0RF93yLTZscLLER1Gsug4qldMcmy5HJenrBQjkRDkIag+xGgdIUsRvVOJY
wQ47YLwDyL6+wqZw52plTcIb1/xhEFJSqx5zsLx/LLP+g/Jj3d2PCzlde/WlrWyDFHqT1hHBmLAB
SqCf3WkvwETO/b+Q3uFTkn9O06Ao51GBgiMPv9CjTAhGB5tDOoPjFY7PPTMibnmDMHFbDmc25iXk
s1o9eI/QLNsXXw9H4xR4Xjpv0nfMXFVvOPHuqdiaIo9A8y0wIHxdY/Z+31F7Yyki/KAd8P2MmRX+
pCtdw8MawdJuWbvNhyzjonCkb6tvpEKDQYjFYHnDehn5Xi4TwRc2ROgvXYa7wXKyjLmHmSG/Ftqh
9tEUP94lQk3UbPstZxWJJRd192ZuOqe1rUj1PDmK+aSMnxROp7exBGt2wbNIEtApWOK7i5npbFu5
QWo6hRS8geLQrQDNv8jJ+YqCbYW3eJRE6XVdPtRw1OIwZX4STJJwB511RfHZasVL36eQkgGjMS1V
PkM1vgI6RPfPwWL+xaXk8oSgRJ3aNFdegblGw20d5w/lTTpRNZkwJhFMlsOkZ7O0x7wpSLi6DLpR
g8LENcoS52hMXSK9ASsjR8jYqbomkMTISpvjR/MCcKubmMh8vjeP7DOyKDzBvOFmTinqbrGOjJ/Z
vMztXY6yHZKRtAvKS/71cg7MJ4bSzNU/mQ/dKT/dD4rKg3z9Ifp6rmtL8lpnMcc9f/RT2uYDBE3b
ovlKkNMebVkevSTL5oBkaVns0Cmys/I9ErJPiJzf6V2btsBPW0P7/fXxdjPcSqQxC94WNQu6gK0l
SXjCuZYY3dsVbq3m2kxWa/Ua8EDIp0VRdsNi6dezt7sKLL5O28hZtTc6ecSFD7KCPPPLsUFbP7Mp
qsm6QQSzw6tPfITQIJlr0qH3ggrcAKMo87wg+fl97JezzR5JGcVNYyxnzf98fs1+37p0Yzxv360X
JF/WfP/6KTgd38xtrEZvyJVyumIlAOhALrBb8YdDKSSVD6lQj+STeo9nei+4hEPwR2HtdIedW3O+
vqlKlf/7T4xEUKq/pK+h1Q5XNqrU+etAN2oZ/iCtQAAJxnXnk/SY+Sen9pQDdlc7JS7Hot1tmiHe
eIUct2TgTnwPOeQ7rERejuygRZ/fYFucw2dzzKN9rNAh4kaQ333axO9hub7TeU+U/sd91ZX3yJVT
sxULcp/sKIox0ZzeymIAIroefe5Kidyh4WliW3MNUeNndnjLMAlMQtbQFxJnk1DVfn5uUwEaa1PS
11el09rPHD9xbggYmIkFf0IaaVRGBQCv/qMkH+89lpuTm5NHCHlpBS9Mq9lnnb4kBC7lUD1n96ew
gmasFWuaKd5qUBAV15K3v19MdsKYbygW79NYOVo5cAykAPTgkwsT8vS50lI3VUKtqYhJve02P0ZQ
KCAcWGhfmaJntOcIzOwfsoMwhWqDMk6yA6XHXe/8QIkafnHIL3FMAfeKEvHodPtF0+s1sO+74Pba
yp/LX18EO3tYxudx7ckzUbZyJSasWGNECMQRegx7aKT9h6287AZ3nFmxQfpJrxb1UyGkKkXLAVKX
FQfD83FoN0LK7y8+z4ueyR5stuqP3rsFnx4CeQogLtpx+3XpFmb3XGdsxqOj9nTNZHDm77XrCo22
WLhAQWAiDv4i2ng86qNYhvRak3Q4VKvY8iCwTagVbrXNTyOiHG1PPntvCJJoX+D+5TzJYIed2e+C
v+/SaeCrLlWDM1UijavJav0t9J2TAm9YaNmR9YV5itzuk0HLaPDdrlWGZLaG49IhbsaebCTmWCYX
T9XDJljrSmDAaEwc8qOX+fMYnh0eZm8pRYZX0Xz4hbzz1B+2uo1N5mi4uhCIo7B4jzJqJbgcRVCW
Y+F+Uu5+FDSlGsL7xfpkrZ9DN0/wSQuLi76mQ7zYqbBggC1W2Jark6mxZUFESiwJkLe9h8Wzae++
GaMpTacBA8A3zEyU/T+z98EuaWj/RmCk7BcDnyNwjVf9ldxJRulo3EyZVFhUbBJE/2ZuBnBNmFPp
BSJl3uoDSipnA/BHUIqPqPrCHS9su5UUB6aM6QQ8TOXbLxwbsxbclG5twj8PtNAUJaNSjxGoN4QJ
P1ygugQ31HekX4gwclAhrvA3ic2ibZD+E8sZhzHxK528PkAYRyWCRPBeicV2ss1VsVtHz/086OlX
4qV0d1xJnJJXCBVgHUjcAl/ihjJ2IWONV6SEDv0A0XHhxOnbx7BYbsxfiZzHV5qXsgCCDFSq6QbD
4Q6xzg4EvOEJGmSI04duEX90+UyvY/5dFbKJ0Y00Oec92gia543ofuBHShfgLfbk1p/cQXisefjK
mVR9fzx2AaR0gxZH/AfOmRlcnu2s5B7p0TLwMpEgUnIdmnGhdWKAPimfJeXggHzCNsModQE33lQk
FEWfORPmMK0XNpZPXt2O3GPes/Fw1KZNsdlddcs3n0R4UwZqPPeNmrDXiegu/5//jl8EIrSXpuNT
EGfM9Ry16+C1lrPmVesUqvuXDFbUt+i/n3ksQaYYaCYrUJ24TWPfKDclXZPqtTtTpc8aESZFldqE
uWzqtQ/cBckO84JxM6jRyNnVB/RBu61BZfbJ1an85CYSNFnonKjIgx+cqdeHR2AwtDpKnyE8Uyn4
W6ztHHG/w+kR0AvGVAbgRrDqpkbC7undemtPM4soi8JXCLWp7Exb23POFQnQ2caM6RK5am6c0emh
aDsomZs96HSX9igU5Vael9smc+iRVRU4vFf/dT2SMZhsdwAZoczBHFL4dm7y9SLIo9POxlCxufe7
IwzglJiNrqrsJZxqpwIjdKtkpM8wdr5MnF+/Dh2D9UZmVNo6DUnrl4vVy/9S0WeYBoC3SKDm4Flq
JvTjhebNL65mV1AIkzfPVOBS0ADh0M3kvpXY4kCi4h36Lf7e5zaXniueWCwHpfhtwYNr5ojHPIlE
l+K9Ns5BdJ1fhIkA0fXknJdImbfeorvi3gXRIq7mbYfziUr8TGGcxmbUL8i1i6FpyQLw9C57FPJL
DWpebdcScxnFTIab6tRRX3vl4Fd8tLcCtD7Fm6kGBNN2g+IYgYhB0T+8K6anBCSDm9pNdfV4Ikwi
DDSv+fPQpy3/1lV+d4A98E32QYOYYF79fLDsS8O6Nx1QaLRCz/eEyCaKWua1zrYcj2UGw/89cfQ+
mSMUj1E6NJ+bdKLelkrJuV0OpCzKrUB2Tl5lP1KMyn9vWBiQuL5brrbvDavblMDcSaSgITISHsYm
19T6UNodyRd0v6NHaQ/zbdb530Ngxvzj7ynY/NfrRtZ32h+bRSehRcNdgyQe0tnqhXIjArPbezqT
8rbg362Lb2JD9lpdUWq43ee6is/VsNoUV5aoJAXccV08i4E4jzmL7p1uppuN4lenBxF0QOr25aQ2
f5zytrtE2yDB57GWD2SxXxv5JHN6euRA0oZZVwPcDtijo30AOjkypBh7KM4/qEuW135T4sHothDv
YPnjX1uj16HzrJjlZSVO4uBycPku7i4GjR80s1D+YgJiGEmRQuL1gXTiJk1bWJ2OX0MVnxfsX9KF
Hst9q0NCkj5sx29/Hk2oFaDetpQ+rwWLB8jO7OtGAE+vFlxdQH/biT0zLd2itPNnSfZkAzHEd3P5
E3ozOblev02Z1zTzSyES4le2QIl0tRvlX/Nsugn/Gwvh+Ho9SGnFn7VGoA2ThVjRgmiHmQZv3R25
sm12zBuc8aS8E4G4tuvYGq/fqejyT8rHfT4MWcz9l57MYb2E72jGuOSZGGLZ1yZO9G+a+O2oUL7H
bFYgEGiB7Lp+cqOkAuBkdOobR65gjxJ50kEdjOYNA00b2UjTZsURDgI6TRqRk/Tbsgzq/33B7kcX
iouMIyQDfvXQtDw2aXD/DcCYfaTKOjS8xL1367l/F2PpN/Pgk8bxroQZlBhpLkJgF8OL1jX0pSBd
h1cBFT3bz0Ysm0wW8rEeKUy2kMsE/K6ihMfeZCF3zrgoXnRRVy/aoRAo2Cyd1+wfuHOm5IKM/nWN
0ptc+EBvIMPLYlwTjZ8m9beAHsZNXCZMWk1iXwM0D28BEpYVCGjniGfjUzTo+uhn9MYXYyocLecY
sBCjnxweFW7u/3vBOY4x71mW06ycVoV1L0rRlerOysevIwS0+WOhb+JMNS94r/hx7uil6p4P76kl
wZUSzoCb7tizD6XOiIv7EFd2bcODRBBVLhtTq0DcNr/lTO13Or/QHUuLlM8mUdiYIPp9bfskoSXl
v6+fdI35XrAw72KixfgWXWydFEhkhVoBGUo+OLq6F+/euEQ3SfxMBcmIILunZoNO48ZIJpqRzarc
AhhsbFeoiXx8513wSOEigh4APsvM78sNv7qCS4bIb/Y8wtzZ/c/aCtl907MANorX4RuwSj5sfsh4
YOo0lqdZ3+6ki0imx2LvNCNQumpTTZLxsPGskALmkqUl6De8Fo3SlqN51GBnY8D4YTRHu6X4wfc3
uJRGhjnJAhSfL6Du5mIJulSltr+r5sLUQxW8Ys3LSt9JsO0jkwalhFIbLpNKXkuN8jJB1i29xe5g
r0P+r+a5ZjfQGJQrxhnRKLP0dRldleErr7dvokZR0N00J4QBfHzLghCWQWiLkIZYYAkAPlvR0QL7
NvJg4Em83UQu2FjGcLuRxyaj0+6GZuG3AtQUgw+TrWobKe2CV4mKrPMCGiEXjB4n5amHIN6F61cc
4UPa/fF08Y8QsmkOEs1akGHQTndhy2I6D43I+2EB7q0902BDJQvFGLCg+ojXVUnTkgCbEFQ7kowF
dK5K9g0nnrfMPrXA+qKp0vPedbr+d67ql6sJ8lfAFOW2ahcZbsLoD0prqeRAkJ2ieVsic6/VLGJ5
0wWPfhU08lGPHPtsaH/RUtlC/zkvwNKmJ7idPVmeW2Q02ZJbmHAmJh3kMXC48eW9ldplaeRveANs
icXr1cE2zp2a6lL8gCkGKSViPdGIfiPXg5HiFZGEjhve97MBJx/g6f5zyU3o1CcPzBXr/2ZItJo0
c2sbDYYue3LuV3n3fJ+LE6B76zBh2l0rf/FgCfg/3OZvrSfKKgV7iqS3TqkRCLAppw07T/sRYG9O
mh241EVZgGCzDLkPbC3QCJxfZg+eRW1kHc2VrlyTxd7ibCqW8pRrBqBpKPKE2ziB6p+a1cH+DR8v
fZRfg0MA7EAiICaTgK2piUn0LiBCETigbwuMp4Ibx+3OMN9otbmXodG80LhjHn+Shg2BxjxLxfvI
Oaigd9gd/ivffgqfA0DkNSJw5VyGU6FNAaqRY2hEkhw3Dng875ulQnrs+CQ++UDpN/jGnRPYt2Qg
viyAtbvZ24xGSvHli0sGZA5CsfE9hqgErbi1ZffHeekmpt22aNFOv6wB6SeLKXGFWG0hTJzwKCS7
PfNbL0e2cAgtTzj3h2nfcVK52hidjm+wWLv3xJGFEcwMiVF/wHW+VoZ5A4fvZrbBI3+1BIy6EigE
6EvB8scjwO/gR2Euh3TTRUPiYOmVK1kgyBe05GOymuaXzZeUkF9rY+N8VSVgSlSDxoBoSooxoHrv
tCb1Q89IuSk36hL0JoQgiVWkenfaoZD59W/bY37bih5AeONlayK0qBYgrRBk3Glw6IupBO05Hnn8
OiMbUPq/JoxpEuNX4SkVTnoYOvbfuyTZ4aw3fzYVmKTyowMp6nEXmEm1/6lT3IsV8oWjbHyknBfj
aBxg4b2GRUyVTnOCrkVLSzULQqpWQdeOyJksxZSmd6A49e0Gk/TZDKjDolbnH/8vtnRSd5zg4fYn
K8LfxVoaqfgci/ccxjmL2lMVIrS9n0nYDKdksECxuNkdJz0QCcZsYEluhbIGORmNvUuEaI1+gwPh
zsL1Lp/TPxf/pBoq7RxSxrAgh9SMXM1NM9/1Ynb3h1D+zniLvKyTtA28dJoOl1zrBBY8FOTE1qqk
ftBSaji2hnG9KEyeL5enJylW9FcHXDXDvqTKWc5m54ufDYeEczEH0HKm1qj/n9rjz8i19tDr5qBc
vNhN6VLiUJhFvzrZqPYrkFR1VxmM7/uN9wRZDgDH4PjMmB2N9jT96o+sb4Gta9feg/+e7K1xFqqS
pY+Ov7S/Y60aUIPWLelK38mPN4vtSU4JIwYvKJ+oMSWO8L5mPPWdfZzIUnyNCXgMcI8dFMDv1mb0
zX16/m/45fZTsDSJO8du8bajairMNC/sZEkruUxss/WR8XTFy1Q9m8vuCrckE9mrvvBDvXD8cGLS
Y3zNEYwUd7tkyIPbWAwHupSDsZjJ2yRAfQiOGDknpWQzk6Ltr60ZgvDMubTE6TaylzXVtwZf32w7
EEvkm6fT17BLGePOCopOYolC380TizQf9HLvpoZdUDcmFM75JBGNgmoh2+elwuA6Kk91ZbGLZqHV
Q/1mv7aiNwFHeIQKwstg8qsryC+6rgqwOeLmDm55otnLvV8YUMKuc1nyaeA8ucDLgC0ER7Vkizix
xjt2JE+F8fssr1iW1zZ+GcpQBO1BpvPCR53SvZJ5taBrZUt0ywI6D8fSnksgPUjFmMvkQMiQQg7W
0iSPU8vdSfDAS2GD8zRGLPzMl9BSFNm0K0T8BeP5KrPG3RRM6l0YKhOiYyUfWa7PNhgmdEAZFXCd
CoSVmg7KVnOnACyVa+Rbak9+0tUsPK7Izk5p83Mka7+TOcab9o0dCMtpoiMQR7Be5/x9r5QaE4xu
6jL52GyDuwWbwf0oexUjEVlM5Z5ARl6dtO7TbPB5RSDmqPs05OOSwJgNSPmwI5I+3it9FVJppdmk
pW2VhFSx/UU2kOQJk32MVg4oU7JtvitwqxwrFW5lwv88+jzW3oEaUHWOoHZ+r4LO942rX9SHJl/t
vQHlvS7OwrQd9q6rUhwbeBauMPNL5yHzKaDwONa0UlQ8PcmXe+hagaLCLpLRbQQzRv75EG7gZoPU
lLzL90/+mz+sWXy/RZy/8+ms9GP83olW7ZvsePvkpqQcYbJH04sf3q+e0CnVOOvGc5nR07UAZjr/
q6VvGPtR3qwSsOZbHjjrDBkjyWEnpPcgF8BFIGb/Sqj6EDIVRXXAyBzNd8ewWXUgdf7CPbzX9zTH
fSZi4Sx3wh/ulT/Ni+8in/bGtoSU3iEhIFTZ61wYiLV2EO0zlraz5YAmMrA2kYq1IcLiRlpeUl+M
+kzAaQLlwI1IBKJln+Gg0KqOvD2+zdUBhvJGAG1GJqvptaPCmgNSD2aaCwPLP9UCjYAf+vXHS+R1
DM4OjRwRd/zS7HIQ8/o7IV8Hm3MGUwhM89JXLlNYZq7wItytk3HXeqsAq3hxnSjxYvafR25ct9Li
Dep9sls0J1ClielODGrDZiAJeFDMh/wBHZoYlARHoMTJIUOVs6UwSX8PZrfDIvXl50afcnO4ij8m
AMYPIf2GEpayGRbXC+Pylsi2ek5/ESGTPsJfyOhdQnvNmkpCVXebDp/jqv0tlEyKhENg88dYVbsX
4JVjP5j5/hxRxAFNOGJVaWpu4JCTpVKEsx4n0oiIAQTmOdLIvt8w0wkS+G/mnYAHn5N6/fk9+r7s
KHaRiJrpG235gdDcz1bqWczim/s6QPQ4h04uwyNAV2+UEMb8mfFqw1ET177MThX5k1ZOV4xv4Qjd
1JMA53W5iRYe7N3K9IzY/kPt2U/7LgHvZ4ahVLHSBP5Hwa1pEuDDOoURhaje7yd0CCme8LoKEZsO
MIZ8mM04KnuKYXzX6CIBwDvxcmxM/k6xa+gnFWcRyW3bWBGBHAVnOlWH+vrzbt1YLaKB3NQm2x7E
sQCL3vjKNznuaKK81i5WaZTzmarNll5zTbEjBN9qW1cD41RKg711O14EDS3ldjSugJjFlja5WKSj
OjIk0N4bC7EGShTjN9j2SDn2L03wETWCIRKsHexNHx8oLF5avljAeMNLJNz4r/OKVJcQC88E09Z/
cSH76RnbeqDtXnbSdXcIXzPzv90qThcUlgjzqpDQ6/IqpjScrEsCQEhsTWOfU4DHhEcC7oWJWGTy
wzwShtR+BMe0iULVqnZL+ik3rf7s1/IuwPtCrnfPmuSH3tNjdoin5g+T84BOcd7sqQFs23DgZVb4
qVHYFezDLZ1ky7dz9oDdhoKcS6JeJzUOeHQbOgozXc0EghbYYPc5gtqia6Jt14lf9mwELjDXcWfC
9SQU5DrYzTR71cntiFs18cWknHbXOQTeTGtqig4ZVRxtZ9z8mBSbrg1+4lcef54u0Bvcxdzpt4gV
QX5my4OYPciTclGlKMeaA+3aQzIjZJk4VnUrAWXRbfoYaWP9Xov8FNjFgvLqgd4pLP7bFPAczD2j
kVcA2I2GAKElP/FrWPWu8zKQgczDlRQaOO6fKsczrDosKgZkYY/9xM5MtELr99DC8iMuBQADnvCj
4dG9XsbwPLF1ZK6eGJZi0NJLaDDpOAJ/XYEi/RL/JX4LUGamVOzDeQJ/llRYgcfzBKbOvLrbdrlp
1RgWdijT2QARzZG6uLOGnkFcZCcVoenao8NQVOq44qXZbvcz7/zHehSRd5g8P4P1qPHp9+siiDi7
V8Uj3QKr6f+zcwaBQSvoaP5nktVMiAAcJXVNsnoGm886nbIxnWu2wVQ4alLBSKHoLSM04uTWBmCd
3T+hE8mdiUpuV0x0miCYTJOthoAUiAnri3gN2deaHSQx2HS6kKomFom+2XH2mljDlmlzdprnIr51
7s4xOwhUKDPAb3VCX/8AIz03aSeZil6ZDke3ryOjb1vq7dt2nsq/1lnAqLwMA7GUZCPDDrYu3WbX
E2KH+7ANKDD8L2jmlkhkPww7NLMW8cEXzcyy/AaiWZ+D4EFYBsiVICvTHbST/b5sCabTPX/W1x5D
uexvWoHFG9Qn1R7qaMaeht1SJCgReJKijicgTcZ1jimFIvkryG/XTo6V2ZeW0Nga6n7Seg8LwXvi
xA1TPlWVOmNlv4YVsAftERGKamNeIHqGQ84d6VZMjnlha0DrvyqrKU3KMRHIFBKMYiwDNaTjNMn4
kE1hF/hwivtp9vmgtmFavcmZkPG3RXxrzbmDOc9NFdW62QxoqjZ6D3dT5N1VMcvWhhyBfPs8gtSm
NRP9NRjgReYXZ/Fqv6xMC0cN6nyDoG71DT9ukV/PxTc9YT+EAwHLUFdJIjpRi//Aqe4BP2ylLyxr
mGQclOzzVasLrdleSv/t+hQ7T3vIAauLUP7Czb5iF4vNNQ4y6/qtRlxlGizRN3M/MEB3FrKFaIzm
CBpTOy3nfK7q6vavZTQ4MpMtwKy7EF4x3ujYD4FRiaWtuqjzE+Hv1n3xrgs45JWlCp9JdR9JkmU3
BSkaTiBFn28mIH/gK1TsKlUjkt66oRrj2DtS/sc0aYDXDI/P5h433AZi6N312+o7MaNznCv33Kah
9ilRQ5KuGs+2v709ZjIpQV8O6UZXsijpJeXL8xXF/iwbDGm/qD0dCemnrdMnQcvJ84Nq24ae/ycs
xTbHYrtiGR2jrhWL2TRuw++1gRpptYFQGUvWdX3ReT/SOBUBrH7tbQtrtjYhFkwbQ0AWusyEiLY9
x+PrnVtPD6u2FC5Jf5ukC8PoWr4d2WESqnosd0Uz4yigqGqrMY9tUDuWchcvTaSPlOn3NEjMIYCL
vZkS8gxbfhjOJrLZVMLfivjQLiGqF1Qxx4Qgs09vl0HFs19gVrhrzKoOS5i9RWlWpdh/6QC+uuCs
LXPMhCTkg3L7exih3EJreaD8qCj9e9CwGvMSiYG9iAJ7vkBs5mBUz0ix3q2xfKWSVnXDfo2nWTJ+
YjtZSY3Evv7rh0ak1UTT1h3xPUJimy9AoXGcImWkiWDKkwsL7rkqgcD33lxCwcvK1qwd5mLuC5Lp
KKusF7L7nkkuog6xTl8zwcgVu5ZkNrhbZ0vOl98JyBG9Vxnz/wsOQjlw5SMrjpG+gad0ShUZGo6T
SPo0ZgbNeA5GE/BTWgeKk3bMldY64W0Fv22t1Va9EQxVGPsXPU/1oBFPM11+j/ZHBlMbEGnecePF
NR1kMA8mxTV00HRh5joOzyWqDE7dCPk3vde8hYw0jOLJpXCle3XJ3MHREXBEZr7wsM8reRSMh68z
i8cCcRNGHdQEiR1UU+mNzJX3BxbpK6tJlpPNaNRhMYh1CRzYdwvNnQ85uX77GQ2JoHoM9gf3x7LG
9HJ8ly8/Mn8gemBAQy7mlDRH4Wqqocy08tiDjPzFRc2HEx6jTSkG/lA5Hu8TheAAO70b3d34VnYL
RBVElLvfMYi8hZazdixYk1EB4hImCkGqoFadxOqK6e0x6svm6zzBon6iSUvhiAEiDlu/8DZrIit8
IzR4pl4+0PU2bf5yo/vJlR3ryFjvAh+5Jc+bDhSElpfwIviEwvfpjinrmrQ6frk/RWwCgmBdBBcg
1eVAydTyl75I0plYbxdozqd0rUsMpFQNAu1dpA+7gQ7ch+30uBdzV2JTr3og6INrRlfvROZGU4ZP
/+AlSP0G4kJNiv1mBZHGVYiYrBc80Y2zT5JsmYmL03Iy9I7FyIkGCNpKz1wHd5H2tmSmfT95aFzI
P6X27g08DChh4chW34I98fqSeEavoGWen8MTa8K6bsm1RymKVlBVvVQFYRZudj5cguCih4JPV9I0
jmsW5yNKNZMxgZzSSLG1B97jcpsfwYu6uTP9uY8KEchDUtVDpA+pSwXxcp+fCLEUMnH6GxeiFAVs
RG0YCPTPWzKDhbX2pjXV8OSV1vlE2AaVBwJ0puB2hflh5fdus4VTPTsDhN0YELJ70K0YKjewST9W
4PVOo57q6CbPpbOpGNQyFHUoJ2gmePpz26NkBitggpc1PZ+PWh+4eYfB3ynSZU7WaqO4kIK3xmqj
rQOX4FloLQO8vJDNMiNjhli1WGjAOlwFWHQnzAeoDjKbNfayouQbMCak0mBhWyVsmVezkqfJT64q
35XWBVAFHXQG+/IZl/VqY55x1v07S2MbtK/jhMmn2o3AxaqMPLPaqEw+DU6fDfyu9kiDciDvbikm
R247abeOTv2uVyhxsiu4uIYt5/xS/VeePA+uhmodNmCRN9Kx1uTPDU+qvenRqnOLfNnnRwVMcviI
JAzUYarJMQ/+TABcEv9sBigd9cBLBHahFYC1zkpGg3gRE673sFwn4ztI6AShfebUbyGOwooxBsDv
wO7hp9HMTv8A47xYftoly/j7n5RpCzvoR8WRDFiDbIfq9B5iB1jMOOzZo/ctkb8hpABFQZDT97aH
sU3ckwUQpKbjWIPLosNsjuA0olXeN7CgOSZ8qvRWgvpCPnouRLHrI/Usd1L1oD7ebo6p11rXq8nr
CCojC/14AWstSGoLvmTQrC3zpd5mEy30V6GEu2Gl3Rqnw1ARf/sl6lFs4jmjNUZ0ne+lcfOiaSmK
hHY6hmfGo9Uiqa430DM6YNSehZ+1TiX3kBqMvKyAVhRMcHE3UXCrbuM5C840LRXppw4UWaITi4XP
iyzDg3tBepoOORd8AwbMUi6t5jqlW0mLhqq4jLpddCEdtszrwGq6F0/mLVo6eu8ceS61wUPHKUIM
7Xco749zvOVOq6qC+HYMdnyyNazLWRQ2YcuskDBuYZJVXIpHCz1CzWLfEM/N+enHaLY7aSa0D0zi
8qhZH3P+bQmhLwUxtq1CuG4UkQx8hsYKz8oGuPvd+4uu0Jmd9/asfGYm/FnZis45ky54YvfrKKu8
nTH/N+2W4kH1Phg4owkHY2CP6ujjfNOP74JRXs1d64+Vg6DHNHAlzPbM7DkraVtmgDSRYQeseHYC
34c4kr+ZxVtkmVKnZNgDfu5WHLFzbvKTTvnIqvP6Vo6fGpxq67y1rerXUMP9rSkswGUsEkQ11Ep3
s0VeWF/5PggrDeuXW9fPg7uR+LzodeiRgrP3CDyr+J9WAuG7pdOnndTxMRcGJWkcCV92RxmZaiI6
wOmNwtO4MSUg43aVLD03j94+8QGhK0ANA6T9N+p9hdf2DlEffZDHnDtP4CINS2dMj7nMTBS1VVGG
qAmexk2LbirBZzpBy2RUrFLZPbBTIFg1UhseTYLlvQ07rtvthfTcvt5alLyOJPm/SWM69VbLqC6G
XNXjhXYyav7vg/M8W6y/JgsBfuOZorZBHWP0LHPPH2gLiYuoyG/BG+1JknnI0/UnKFhSq6C6/wd9
4vb41ifpcAdQtovkvyWh00xjxl7bnON8VL5Pl9rkGoqkmYvQgrSom7I/xj+zE2frFf1K+mXgdeBg
bqgS+tkPu5PPl7xPg5o1jb5nxUoPLw1lmZ1APUN/7zsVjpyZXlefj1z2EJmn+mfMjEjL9PlOfGyq
iWE2VoVPYefUXVCae0R4iLJqkqkF64lTstp8XMknL+x0CJjDgY3/9Pe4f4NdBUTpbH8LZ5A2Askj
WSQBviekI8PG+rF9YNdoXKuKgnRMpBfV7nLudkQ/Hu1m2CWMoBmKP7W0wRFR7wHWGb8ZAuLBhOMS
u+xxCyxAhenZFOLlaynqMHv9TKJWTyNnrdQ+9Lwp3l5EJLiyUGG9RUDe4FzuESc4XrnVTFqPtpph
UXOWgX0FQHj7i2pP+xh/OcUKU58jd3E+EFn4fzoNosZndHkhHJiK0WYsrK1V5bioFhjiYEQjdreA
8tODjqySNX3aS9LXNyti0vJxpwEY+mciQ/DIhFZZjb+zxNJxiHmPp7+743qwJyNJUPOmhngxH2vf
2UVj85/D+e7teyoIdVR0iqS8q32WOXpIHxAelJ2UpEpMzSr6aEZPUDnxRZJJzYm/NJ9n8kqZuy2a
IQSRzar2s0eE+WPqEwk46GgpZR0QLyvIP1t8HmDaTbOehPfmcMRP8/Zop0CeI1QL1Gwv2cDhokje
Gb1Tm17EHDlqlhmpWpwTPahsqNix/RfqPtD+PENKVvu3QcY1nlvgwKu9eHXnuKm7EAANbouWBdEb
1fRnfdnemg8aXmFR58nS65vfKBRqj4ulMHKVlcaw5Rcf7V2ixevjSQre43Tm/6mlD+zYqc/eB9n5
dSK000ct5d9ucDP1Irl5ne9D2Muk4KoIcd4Mj2vX2EKXsGomKWimvPb1hmrOQlqTSYWPmr0XVAIy
2qCTQI2flsVtoBr9DZ2cyfJvBG7dh3A8aBSgmJBeYDD94sL6Mb4Gau8jt7ff2f3esJX6REAfq60C
jdbkvlzIc3mNZo+A4z4RLZoC2VKn/4FZdUHrH60qujAJ1oVdkE+nCvkAshgjOuhhhoku4HRdgS4f
IkbYWCRtWNDyA2dY1Zdt1Jt69pIZNkeu3/ocxuVNnLHrTeMR6IfDym/XltZCdD8fZINkQWpD5JXg
a0kHZrhg+trUhepcZy6mQw1OLBlfGl1nmPWr36//Yptn//7Z3DQV9pdZ5fq7S2jIAeE8/CkH17cc
glr7XliRigzB3pQ3aTQatuo7rVb8nRw6pHBCGfSRJNT//6sdPw7PYw4REN0Ia84WieS9j4czx4wb
LQMrvbozZyDNIKA6H16TjqugoGtTS8QxXTEUkyRLuA6gZUhdS5r6SMe07iR74HfPis5MhSb7mWde
8TG80izES6qJC65q+4zZsWK82yjgm39My/6uzoQOLNPvnPC1b5yEmFCN2ZHsKTZ/ftbKN2Cl6Klk
dCMBeQ0R23LcIHhG+0l/G8J5b3S3/120S0ep9ge0v/u4ghiL4H43NSf+Mn8T7H0tiMZlAqgVyXEh
3/moi3dceT3nzECGhW9UryJpCqbOCXhyspwEPWbbVof5J43AXYcCWPvYierCogxwR5lIxHj31LHU
6W1UC0t6U6ED54tsldF4akQc3h6lcwNE1lxsK8zS6s+DF78vwQwms4CLtoZgWAwokfIuFfKVhaTT
CvNqLSGfR+PWpRSQ+IZ5rEoPeVTtFG+rzFOpXQVhgBYfh8lib+M0N46snDGzfMV6AF3+9hs69I7q
j8m+nHPRhhgE8Mq43x5DIo8nV8gl0GZHuLhYIcvue326Wv9ZAds2n/qrOeIDFg+4BOHOUTlgws/q
NqcFFEjJGJ0RVTNflhxrQQ8EyLiEOEsiJ+8KsWwyasRWaTZfU4/JUr/ocR/WWaXFqK6WhHcbYFME
19i1yCOtaDT9Dv+vV5w9CdQxoWUxX/E3bGfXtWRMQWT9dfurRZfHp/CwX028i2F28TyysMPLdP55
ntn9bCrWuIy2UiYshW4CZ8Gsf9iEAPP+ftR/8HNrMFXMql7P1SZQBFLtgS2NCPgS0ZTLOeTvSTkq
UrDDa7/84Xr1Y2cBmFk7Vq1kaSDVqjstQD2r9A5mRHn6OsZtvoPrcbsClGVO3SETr/mG0POAZJCg
UZlRmNZiBx3PvzvIIrAUJzzz9Q3rvOSK0KldJAawt3QeRS97HVYwkrzk7t2ozto0vYNrOMTqGTkn
fHXt4RyJTRo/u2Y2VMhtXqeRwHGm5/R7eBpw8b2B0ZSK+TcG0Ma+YwjK/6GE6fwUZgj1AcbalhUR
Idn2fKxpm2NlDM/YwvrMpt4ZNkxB7FBVIhJ/N1/7rfmJ1ESoagxEBNZpk3pG8BgU5LvSBsKk3miP
qyV0kmz1eF1b7spDA8LB9weHGNigdi+hDBlusJRP5Mn/uTSR9BOHaBa2vWctbOC1XORLMwhDRfKi
eQt8FO/Pv/G53/gP/u//3GpYQQ9w85WzR7VDBclmHDei29QuG+F6G5DM56J9VPubLBr0bLfvFW2j
JHX3IARR0QrV+V/xAe3G5nYZ3fj9k2ePVNrcgsKVb5bWhwYfkn/yd2ndym4/fxaAKWlKbRv9+spZ
x5zHXmJb4VzHXwKQLUwGzdDeQUQOA36LUVcDe8sp6YJd8my2xIi97LSIvFFXMBsE3In3bdJjEcNX
Ye4rUrI4q3jIGDW601GxfHmDaLJpqF0YV186fjeM3tEbGClmdZMG/jEwM9F0rpXIgNUiQkE035DJ
f5kk8qcqPErnA2MSOm9Q33Pt9xfkgx1cROJX4sxKBQKjBURVbH2z/QbYTAm62Xm9jHXzPnpqNxgt
VdQFMbSJ4NA/epXrm+EHY20OWefYuqMP7xuzSrX3AhQdNLfYl1XIYhwajdQotqpnRupCl5tuA2UH
1yuvxXwRpK7wZ6w+i8zNYzq3fYpm4iMJNv3HEad0VOp9fsEeCppiQAjQozvhvyE3LjQocserWN7o
gxBd3tyIHbFS74zhYfXZZxoW2nXW0WqB6hYWvOj0ZUm1qU0Mto94AklNRv8gJ6ZyTA5U5uiY1uLX
ZeH7jUmIWKkFfR9/I3ahZeJwsYUuJx3aqNWJeL2QQxMv9NYx0XBpR9jrqzMlmKx88B06La3X84tc
07fm/S/HGzHYLp/pGT/9yeuqQiSkYtdXrTJsLeUDipuoI/87048/gwQhfHbly8sviG4pcTrjrJF1
T3PsWYgyx+aUto3TaooBD/OG3oLc5+KY2y/1ufz/G++bPu6vusSSa0kMXn4Q7SlZxZmoxCSDN2Bw
JgoY/ykDfEoLi0xrMlOjwYYhe4gGWGac7H252P9nkq6QKyMO8wKyrzZq3WtyXstd2df5Hmyjf79T
FoxSqMFylc4wW+TJ1eOMcghpXM8bqTCE2WL9J/6zYwke+bbpRaksVx7RvAljLt4cKmSX9LKtEbTo
cg3vfEBozyiemwIfrkrk3TniZfxho1EMqCX5p1uc8IrTbZkLxE758VyfRC5A/RjwPdij0xn7SvcQ
FrS5rlP/IdAsawMTIVgmd1ktf/z4oLveS6iHS/A9QXUGTTRwtn8PuduMwqf3QecFv3VeWDAfVeXX
NUymXKonUM9/xrBMIaBwyBGSHSA1sGQDoV9hvLLk3FRxCoTpAvB2NLn1kzQL/OOGSKnlHEakXl7W
zq2v52ZVE2xVAx6Q20r6Ydqheht8lCloIzccSLErSJUlHieEtZtdc655+NtGezC+tZY7WXEFDcJ4
5K/J3PAYvcxA9siiX9BA/ANCyeqmuIbEQOqh+FXP0hx4S+2xGj4hr+09hfD08UTedFHC+1GgTfVy
WomaAcv6HAuh/CX+Lj3liECswAP9YAZgb8NBlbNCM88YTuGLsA+Z0hdt9Fb+FMfwMS9lsWOgO53s
fhKedVr5dRvXyNPDpmPNLWYSQn60N8GuAZxXm/ZpIjQkPJYhgdmCwySDFHi38DX663TSiUHsrNsx
SZISQ95Cu61bewMsa4MTQMte05TuT0sNyaQ1XewLIZikRhG/P0EmsRIceRq/J2ox6RgjVx2T9rQB
9/W8d4LEQ6+c/Fh3iPJB6oQGhyT8xjKwwVjifBYwngV0TZb3wMtyLRB5rIltqAC4FbclmLvjIh45
HYhp9O64yiSyye5JPa2XsKVqZjaNYB2yjVC8VQRSXEO64I3AljVziW1a3Dm4CI0p3kT2KgMpbVXU
nUVcS+fvLNC7OCO7z7ALyJ9Yt+bbdegU2vAQKyXpP6gzvTQKExgUtjf8Q3U6YLmKALzq1Sy7gmOs
6hyt/bNrI4O8pybwUdAkrraJh9GJzSD/Nf/W+LcJF5EuUNWmMrFccTkKqJKkNnyqBIkHQC4AN8PI
EZZMvnI=
`protect end_protected

