

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
L9EbKuxxzV/09pnAb0OGW9DxPQ+o+m/MvX4x5f3JCiR63+KWt2eYB17k+9mGgVY+K1VLxoYz0z6V
YvlDefublw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
gJD53XIM6IXGcoGao7b+pChhlJwhGxOuVwSTI1iU+aaEVIG37JelabzUSiGlwgboK2Zv8N9/EzBK
Y9pDSGcMvhlTABOa75VEGmta9QvVzRVMjXtd0b/jrdUkZar600zvkPbB8+QESNshxT7B96klkdIo
XvMdlDR/SEQxmh4Mkpk=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
uMh613zg14bfl9MaiMXKdALr5q+gvlBiCCfJpnudkmj/VEzNaqE3gABSgWbIJEk6l3XEblsHwoSZ
2eueijgOoGBjZq9eDXqLeir52M0Z4RoybrJFqX7YgYE+2quggoW8XJjUPK7bExWH1Wd6un6XRwZo
+XQ53VUhkTgctFKNHRr7bEqxJa0qk8dm+fTRKVmCc1Tr5X6rd28yRrr4koH3+liBwEPKquwcMKJL
zK5B0g+bSiHJvGXlQQpKzQNF3+4MebcveUUQPOYG2FAjfRJs1t60dgE73q6y3I1DMI/3MguCuvoX
78TA3nOFRYGLkISVFXDX28xYA0EnciH3BlzGiA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
2ADp5V47yVkwRII2+UsRY3zvclviExupZdil2h787eVOjYg5odQlZCOMnldkarIbxDBoj52vjMGc
rG04pAKa/Z3oDUnDkDe8ZMmBI29kynugqgc8aGxYPVKp3KD8EvhnicB6/4Tt66g9A8WsjHtxXLuC
0ImlGHU3T8u48JygeUs=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
s5k0DDcwk1Yhkk6mc4rW2ITc+jBCojX0QPFrzARjmvIjcmc9EJT8pAYSdJK1ykoSIGmT8u4U6vaF
5pchZ1NWV4+0T78Lu7ir0M6lHPYDFRgXZTR6CNdPGqAe+Si56W7NnXEM0Yylf/w4tAQ0u+05yvCg
wK+mPCq/91Em5ZiPcvKOHOdJBSTTkSYC7/n0QNniR1mBmd7+dgsFr5yshClYY/q8HngDDE/aNYfx
P9AT4ECjL+OzARXCnbTA6RjbHEjVx1ewIc83WIXkwbZjUYAzp9rYNjFdx68zjq8U1XW92RXAEXCc
AYKv676uVGq/WAryucxGApaihL/izu2+HGUsYA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 30640)
`protect data_block
b6o28heSIHrooY8Xxacc1TSllSk3azlj+0oruI80Yk7KXdGpIrGXi0koLc0XNsJZuj2Z5B/o5Upl
gaVGivfsK10uq4wxqY/Q6ACdB3kjKYJ0uDYs85yjm/ToMKSaTelB7p5JyhA3hWvRveJccWl84Fsb
bT2n+HoKhE9Ce96rZbwDmbxMqwnk0Cn+5rM2eK0XbxWcHcXKuRUYsyFf5rmNM4H5OMDbxwbycPTp
eBxHHM3qhLRYhIhGRKVqjuWnUKx7q5FWSL3+1tIxtuUKv6DdleBy9t4F61hIW97Zt+79r2eBXVT3
/S7QrsgRoHHP3v+GfCEcAmftQXcM8iKk12vyr69dDA+ZG9bduZTvtXmxFkTp7K6yqioF68mWmGOa
oh0iySQESyqtp9oYk0yexutdV6JhGkIvzr2yroPci2jCmur75WtcJPzJEhR07s8wo+8Ewo9i1Z6E
w81ZSKP4IdjKx23cFrQlvBH7Q51lIL7FpbrQWg+arXnrSesoELEzsYCxadYdgtYubnmqNOviiLt0
AnKZpgYscKed6FhmygqSa9cgbD/sDzvJ9p850yAd/uq06kYu/4bpBrgrgW7dGTy7VYWnMssEq0fs
NcRwpJPmSbXkqudKxx5wxJcqT4RnKyJ8aPDCUEBQ83e3BeQFoP5nE9IM7n9jRJk4HCZy5DaJfqyY
giUwWmJaGD2c9Yxuf+067RcXkOsowuQJROzXQ6TDdBvPzkdO+/TIEWv3Imp8ReQVZ/o0furpgHDi
1Bu3ZXjTyzZZcfADVYUikWkyRnsxg3XnvfFF+d4eTGir0MZmTNU0HCDu0nTPdkNzzqSaUwbAKjCJ
KYP3oVFuoZAoSGB0bgiBdRTOKJnrGyy/uODSDhVZtgR5IoINTePtDRIDlCKuNGY6DLfa2j+6/UoD
iV7VjP92bO8dDZHIb4a7wCZXeJJg4X9EsQKNnHZTg2FutrL9KRco1NGvAYV3ous031uPMr6n3TM3
2EKjq1DHsi2faPKahxLmofRB6yU+i4BXU2BV6xW+LTk6rMqkkqvLudd+Ymp2mfPclRvDUSOKmHGb
/orajRoyP0pEP3rqOENfbRXuWolsSbrDiRDc8975n/wUqqK0QlYzXvd2xKpecuaKbgEzPAJZW/nt
1snJ4pfZlVj47F7lN9g61phf2/EMOl7tvDP/GtXnCWlzQpJOCbLIzOQSmZ+JKHciwDtsKspIlsBI
alSpCiuBN74Aq9sDrUAqw/Xpl7g95MmmME5XaupeMUY/4D/1L+jZpGfECEJZQVz/b8Elrm5pCVXg
I5f0fP91A2j/ZU7nOmJ3GFRezwBmSMpHJdsqI0AgshyBDojoQ+gnh/YgHej3s1FZCvyUYHvpitVN
GDEo9Pbe1IxjRK/Zbfp8BB7fGeJHF2Dj/fLw9y6+sQTtrvfOxoRHogMr2U3jCn+/UFk4f2Mp1VFJ
s3dHNY+jwVp4WKpJ/T/1ScOwwmafG8dqI2B1pkEWS3dM6VkyU6ESUcCH/VOdRIeV5SRtv4nfdSmy
CbXA0Vtnb47GCrUMoZ+PnkSdBn4QhhY9/x8GMtYM0fDbwnNF0kt6a/2doTzoRs7OkTfwHhC0SQL3
Ki2tlOwyTKuu+93rXdSoTJGBCYTStW/f5MgY/2pPC+VYPDZvqk4JGR+yaCAEcdgUSdjxyuEhCukG
y3KC2fwcy4IjN9rri5JYPgnDgoR9hxwSVlXt/G7KwdoEBluCdJ4VMN8V33fXrlZ3CaOdbrchNL2g
/wN8eH44k8UzwrgGyKwsCj3Mpa/i1xMf3EbyKoQD26ff6qDZedqPyOVsWX5aBq7x3xSNuPQ1WcTT
afHUrldunlyTE3QMkjPJ4LxC4MECPPBsWS8bj4iJryfs8rlcqWD/3p4Pe0VxCvj2zrTQPqzIeCrJ
4N+YgMGKBKk3woOec1rKV+rj9GuJxx6NlupE++qANFTX+oXFtynYNXUjfWN94VBDpteIUED2ZpjR
JFC2OSeJrSP63bHG7dLFQZ44wdz8rJILre5Ia+5H1qvRU24LGzMLE/5ZHQ4KDbkWnoxRBmq4ArBd
wNjUQxsgF9ib3nHxMu8ZekBYrkRQUkK6foAypzZrrTX2/jL4/pcOxoi5NP8YKQpFMFrht/QQCMh9
DkweMmCEgMQJT+0t20GvyX9Vsh8k3umYqXXzC4EwV8Cz7QhSF9DfoHfX7/vHMrDo7G+k3cDDBplK
WFb9cKS1asMRqYEJ71yC2o+Wu0y1GU00iopfVTcGLJfeAD2Y/QQA9zwiSyw/XJdFNPgq4CpupqtU
zQZaFgNuNo6HEzVvwRkxoxqajjH0yDHMB1W3NdY6m6XSLnZDztuu6QVtwTxUyWkEfLz0GVnw1Bap
UC7wZRSrNHv9AUdlPap0YD8K8xW7ykRCp9663dEInG921vJ1OgjwA7WUOvUcLZtH3KXpJKh8iFPu
+CLj33k05E4wrvduO9D7QBcJpl7aREXyTAnLFbkZ2+TuvTubzpbWmw4EhPOC4oC1/IDMfbsOCUl0
5HXK/FtePom1cKi68SdIvQNM4H4ULgI9/CL/2hgvtirJskrUFbR6Kn4TyxlkVlcM0mGZj3b1/DzX
/EtwPTm+D6MlOMfLqqmVn2ADCQSyiblduPGang+/AbcjbOFKyfGnLISPm4R6fiUVwwDmdDDYY9Iz
sitFbJZKmS0cALHuPpX9c9d8lVn7Lsh/kwew6g/qvHQ2gDGojxEGmHaJJE9oK1GBpCo2eT+tpe1p
01dvReiJwYhMlhFTKdndCEk3SBlXzGJR3lyESyh7/sni1Bq2kHy1FdrHnEbQXuLMgwdURkvpkcXJ
DJIIHasZ7z0ljxh0gi0bgebdlOQnuQ33kar4k7QC0/2ANc1LXvDT8JSyzVoNElGgbEbrsZj79knS
vivBZrzhQBhxESABSiY1XOFogmXcirS0zQyjtlbzzfzUh8bKk5ILRVS3PkpLTaNxTEOV99Ic9kAf
136IUKeYpWI77y27TGlQR/oTeiFI7q3riGdz6w4E1hVySdGxwnxA6Bsv8mmxL72y3aaTBiI3epSr
9ZA5uW9WwBOI8W1BZiMWEtbeC7U8DTxOCoPWelIb1yciN9vomxMRjAY289P1QHVwVS797VnSogYO
CipA9svdNG9rsf31WoLT0jKx0w1LvH5hn/lgYKjEn1VBHa795oOS2EUnhdsou59+zB68Etjyujkb
vbiN3IkURd+dmq6syxTPHD92SVOpt0/wfSpg/JD/qUpvkdwKJ7sE25uNhVuFPzPZTbf72CblOos+
9k1en9N4KKZKN7ygtgeTnWYvIY8IG1CRcWuDe/NBbGqvuG6iI5qIFGoWcMSLOkPIDk6YEgVSYzBl
38EHi1gjYG+v4t5P7kN2OMhLn8+2bKR/4Ji2u4+MJQF3sALP84b4qFFqxGL26lw2JzdSgiFJGfex
uCopAcZSTOgBdbHcdyF2Y5VmQ4wyH/7QCW7qgMpn9qapWHawHvxdSO35HxeKbOyX+mTe3HVniiiu
vnwQ6HdesjJ3eTmzzKaY9La5p6r8Nn8+1U9BZv+dgPD31xB4JYAA04e46SyP5o9Rn+J/RWLHUEaL
4SrOT9dQgodnN5FGcFS+UQuzE4Lfx+/bf7saKl6L67d2aMWD+lloCyzuThyEJH3B8LP1bIIs6JX9
L12uC6I2py00Hy1ZeP+7Hbz3m6+iW9Y1OMsizN8O6c3AX9PwAzsU6/L4mtFGzd/ZpQA08FYSo4Nv
ySq+cs/J1bQYeGQzU3rG3e/FaDhLYHHm1xOlhrO9Hcz5KJ9NcmYJz4O5A4TNSPFoQmS/p/oQLv5a
bavu5u1tFltgRfLnD0GjGdkFbzcxc8QzHmRPatlLkVyhIlyTB/e1tzNrWsW9qQbl6ZFyH/74O2b0
c9nOfDPDUMjLn5jcjMIfxVmgeHkjJyx9EucLgPyFwR8C0SS3ZnbbRwarcg0wl/rHsNdsmnH+UKtP
MoMmya8GjJAldekdFMmLejCPPpWuec5G3p+sYCdqipxj5JDYSw5YlNuAY/X3xM2ZI8jc8R/3/2CJ
1VBBsvmjm66QeE1hQyd4/g/8J3qZLAVVX/gqoVM4gjJscwn7IaNUlBAiI2+bvdJGOskBlCyqFa+p
+p47y8HXg6OmRZL7A5WgjcllAD9QeYiL2l0S1beBYm+77Em2IMZpRhCgXH/44poabUEhTYdNYQJQ
ojZrkMejwkdntv+sFOMBM/Cx2mbi5IO0NDah/KmrWG3LyiLtaVwI3vw/hVkOApKWnsmMeERCQyl1
8+Vobj5Fye+z5x0A9jmqwzcMOlQXsT/D8uNXtTGJVU0cU150kZqqP8Sqq/71O6Tk3wkFviYsfQtj
DvLW6VbfVO7jA42sqUYhnv9fnNSLwgw44pUEurzpugVFdUnUwiju3EKdLguKkEb3Pviqj7DKLsVZ
bs4PxxOeg5m7gR8ENEyUiJe61Mrnlgy3xCk/VQ8+WUihi5iHXeXUJvHrpL2RtEH4QmEJcgFJOjK1
hgJIEU6xT7oPb8eIOAwXYyXaBePlgBPLEtMR547OfIuLk36yNjEa5RZTOOB4grz92Q+Kt12IHvm1
SW8WRJ1hoIb1pNv3nXBVQ5eTrrdlK9+xKv+9MpiVvEhrFaSxGBkJtG1fHSAtf7k0dZnzDnMyWNST
Li63/7sPbNakwei4gcAL7S7bQanpqB09BLC4BXgUWPeOjp3i21BQmbu7t45SmLw1iKdscqS1fD6E
jOVvadRJS6MeybusOlVWp72Qn6Nd6XjM+zeNozvVHY6yxryt/Bykgl6hko85D6CmoTtTjd9DXUfW
1BW23cu9D4fSK+of69V6LvGNwdeTFbNmP0F7DPY3Wuq7nKkQ4QXp6dSfzu0oWgzXwxhyEipCVoPL
cod+5fKlLRtBHBpTxDnVyOwC7jHTJPit6NIq/l2nDjVW7Ppo8RsMq7I5pwDku5HPTl+a5+j93gZ2
SqjBcFloYOuyZFBBGgqUvAigia5k66oOT2YXobGtymc9aIw0Co0+aqzKBlLJxrJ7IWXbzffsFdP0
CSb1MrtI46c+8jNUnRTEzNrBMmjP65JwWY1eN95gQxMiLWOI+AyydfgE0JFH5nLTNS9Gnkzvqay6
V3IJ4Q+shUDplRo/A6UClSzV3WF7TQ2WRxhcYDBBGJiCPUPXlhmGVoEqZlKsq89vWM5O/joC7fcZ
CZRo5DpgWAoPfZzPnFlVRr88SltJUvKR2E7VxqYNMi+vpyWHul5HeupkJn5sHp5yQc/WC7FMbQk7
xBdfrDqhAoFqMC+sYHtXnz9AS6rgD/4ihCrAZ6ZjfBEl9v4NyBQRVRZ90JIC5I6SWUXV64Ov0HG9
GADA+a787zxz/kAs2vUV43wQgyiF5aYRw2T5l6TTgb4XDeOpcgmk6geHn1QWaUkYbp2Lwe8RgQt7
7YDEsL9s79lQ9eAG87k4UvJcFqr3QERfUp1Nemw/AoShY73tBnuhBm5vsp649zE2KYUZ9dk3OOxq
/tJ/8WR4/aDdI7ZGwLLRAPOn457hO+9lytAuSoXC2SaGeCW5vYp9JEu8et1FbHTcPY9wQzcghKF3
NikYr6OtLky0Zz5HvJ5p/nPUw0X9Wag3RSquJA1WbuyPaN4FdERYxUw+aPXkB2LqEb+L3l34uQQv
LWPo0VgryKpvOHhBJNlwaOO8IZ7L2d4ipt+1MHp30vMQQWgAcCPdxH9/KEkDyzNr3/xzyvhG9TD4
OgtXAO+yE042H60lTeKM4d8MFxK0PDl9dQEId3Hy8RrdjZFOrBrgsDVhlAb6d1e3T7e+EAHc3I14
qLHXJwwE7s4caCxZPLYg9GQThSHSZtJ8IK4enPRC/d/JDaOvbNch1fYqeyJVEYxA9xiYqntMQdAc
4p9pGv0mWRbNBZIxovBsfrhmVsZF84cl9FyOl297YiSdM6tJEQ43NLTKCdQi9hk9RDSl49BpdneE
ouswni7wfcFKaqpWjW/lVQJAvGEaEa3AVVM6SQ6PMvQmzFIfwacXlhEOtI6Ml3bC+XbOkgg17w9x
OqBGHQtcWgJ9Yexwkn+zmY8bS1FUhdGBXiAq12mXXPGouiBYEjBhCHzyMTJeTWTRbqVoLZ7adHgy
VoSIFhI0sm8oF/htGG0xyxB7vFhA7oaffdYA5SCSDZHnhLjCd/dVbjxyJ72DlCKsnKh0Fu0ndnsz
N46Nj5O7YQKOmPNbGFsauge/Iy7EnR+r2H4+HTfnhDEaefMLe427RLvCV6TRjDoMBks+n/GKYTST
+9ORQD7rrcOVuhiXDkPAfKDzdY5Pbxg/nzjrOyjqwtwFWdC8/DUxhjxP7O2c8Q1Rl6owV7vUDVx8
Ofwf3CTSUyoFddM0JI9VCNFwkmI/MGTjv323zMYScFwClPzouzFqhAqF1QzpAnYMCJFpCG56lUaC
qHOKJyneekxZJD3tx3KHAXpdDQ3RQ2eKi369vBzWFGMtCupwFXaK58eWqDxFenT7VP+AD3wpD0fV
LFDQuRdQHrGnZW/BLQxNarElJsFtoHfgASLS5vvpCv+Gg9QJKx3bo2+fVbw3IMOKoram4lCiknEn
Q9GEpyUlc/cKf4Eu4T5HtolwBHu+6YV1GfafBKoShOoIINPYAUy0Z6ooLNX+ATnL2Wg0FRwSTl9B
8CET9jFkohTzj/Ap+TRI1YVxUyNcb5KAvy9AcJEUbWTqrhMG63f4B1mPr83W3zG1lnZwyMtDXrU0
Ss/5Sr0r7e7Wh2TP9PRPJsEqElNoCnVGDLJ5lz4ZJ5D0MQybcuLU11C3V6eu7P9Ev8R3Ill/xdBt
W0DHFBMvKxCJ1Atopv90OZsi7hFTQE91aWcICxGXVdZUgHNKxb6J+NkllSONnw5ZX1awbkSQMpy7
frX/ncrtreVUZLk5qEsXeeHPRsbdAaTNI25U/0EjgwFSoW3F9eHYOqd63ImPInf/k4CcfPZYClMC
VUnhYXeyelnF06ginpFZu9TyFpNmu9JRkEYFnbKO28/zkBpvDu9kknoN7LtEzdA0ZjSjQLlrUkL3
vJdy72ScAMKnqd9UP1lAAo5r1nje02gHmhMMkSjH0jhCZDqT2QMeswXDrPDiHT6ZIh+lZKhOzHL2
iVMu/ezG1M/yequ2zhYFrML0bq5vtclvNgIG+P+YeClXQCsMXU1/yT1SXSGBWN+Nx4LsD0JrIMi4
lqlc1lMWJ28d7zvCER/Wa9s3TPPPWLpKmbM9k1RobCqxZ+FtslAFVsxXxGAEAcvimb+dhS/rnCMq
4GzXn9VRCAESkaBcySQBU+JnwBZlx8WzoMUqHVLiXVc1wjxqQEPni4pTNtFNgP3WOi1fejsj6pGK
Ap6fjPJAvmFh2rbrXYo0H7HTkOczK/kh4DTTTgkItB/hCRJGoG5EmJLOIbNdMbRjjI93T2BKgclt
e6u0QSQ1WdFj/8HQwQt/8+W1vZCnv8xSYpacFXqcUX1f3o/8DChNG3LhgkVz4mjPBK973qhN35zY
KugeTCRBfMhGhOvnPjWOdd2cIB6lpqIvl/oKV6EPleoeT4raTfaGbgVsMUI/u6NguLBJtsqSGT5y
YuLtm70spKLnOMxDpvX7JEnEgTlY4RNxwim27YDw1wu9vt6KHJTScdHZUeM1DJyiQLLooxAtn+mK
DvmSah9FMv0wWv47dcJOpPsQh7kUkcHm89meGyt8CA2Ppw/zd4iyW2ppM5yr4mgv3wp252OMoGcd
ysN31CeA4o2MaCncUOdkNOGdsQTvIAFVHkHx5HafaD8TCmVVPXIlZBIGtu7yvXLYOiUQe9Pwk6ov
LuId/aw2bQuW0Hapuq5WDQa8f8bGnAP1Qugo+KuCWZB2t3tl6tNaZBXud+LCLfzVbWgRHj+7K3l4
B9i7z7QzKG+BD0dDyEsA7w+WYad+3y8YPn0Tjosr5NpPFYSWRJa5/uOBg+GwPzHHW8dT9sG6pKma
wqi3zZQNOQlBnSHVwBBNBxHnwY4EtKWldlI3yOWgbgvggWv2kZ2hFOr7ZJKuhBCsrg/9kcjTWZ9u
4cupEH0g2IkemIOXV2AdTYZ2cDnUj0hKTlMeg8R1Qy3UnTBjTLmqgDPH/dg7yxQAEaHC6RE6Iw4B
96BX2TqDzkEck8EF/F7vCmgwwRJntkrdKAtg/WzU1iyr/2cNY+/BeusINtNZJCosWwWLZWD4cTl2
jcjJBSm7WGxDgMtU7nweuXRVTSy0CeSso904jRgg6VSmxshJ5/k3mhCbUS8+4uOsZ/BwdNMh97wU
+Oh4S/z/6uaf3RycOzJUfeg0LDoKkQIc+Di1+6lPWS1SPy1aBLdthiRiv9WOQ6vxp6P9oXTHG1SR
AgfPBJNVNjcpR5kQ6QAJLya6+TXwBPnYV4/Q3KATbFqHHtplU2tQTAQW9jLLoKCBYOtEJmdBjwCC
IHW7R69ziDGFbpMa8y4wxyb0qlzrVEbCYswBJSxs4uU0rooL9EtJjy0vBzGK2VwzCybM+3S9gfTv
A9EuukW7sknyT5fwSIHSt2zWwdS+srjYo++8WppTnIVR311D6lc9NEN1K5SOszbKZQ5Gg5WU4LCR
UvNhWKa8eeMm63U+AhXaSqtdEwGXD8e8sKvFrByVc/Qr5duYLKH04z8INGRP75KEOzWpcuFqNj1t
Kqa7E6F/AVkylopeWBnH7NsenbyMieUz5WFo/q5Avsskva6WKBHzscxEeybQPChtNU9yUx++ODsL
Mw4Vrdfq5NKuv81KrgfN9qGCLbQYKZo95cQKNoQIfPj64daEkSV0lQz11lVwxcAFnqhOWV4B2RWO
ANSvz5JtVblhVuCgvZ121lfcKaSaRdeaCTtyi+q+SViKvggP5n0h4gWv/tRpXykx1uF64FRCwSfn
htC3FIvZjTK4qtuQb7WIKdSj7LX76vDTuvB8g1gN4dPUlbgq79byJSYq8QTa+shXm4No18Zha5HC
A13qscc0uD5PjUB2iQ0DqQ6oOKn7BIu9DTh8PI+pv/YJxdtM0o4hYqkJ5ao5NrQwT5BDc8CGVahz
Va+mEHnbgWkYhcKErM/2AX1FtHtGoTUuHQ+njtESfMGy89GdOdyeY2yVW31j6PHJu7gk3zoXCQde
beDxbCy4nQifW5QhZobJ/wpeC4vi1XQGe3T1KEvLxQ7k9R/TPCtmRSkC0cBqKmTc0Ty/rkYrWixd
iJvkf2IWUUIa8J1+TTSlTc0GViWgrExdfN3rkjHj6ADTsLEThwGPqZXliJp4rzVr0hDH0LsCKAbN
nKdwZdyxkfFvA7sODJSt6zKLpTAwJbnjB2NxLegNPXkq2sdk+fCjbCGlFiuhPhRbTJSYkqZayrg4
/dVsLnjia/EFs8wgiE3wzG6E+NT8jS+EaasAYLxzJI/+gUE0S4LSpYbgKmyUa2ZS6AlpiDTR5zMi
Y3Vv088wdvq4ixYdRgZnQ7VP73Lf4u6fpHJzE+lZGCNxmVNt5CvM98xUEV8SkiaOsLgCtNEg9wYg
s82//f2GizifLbWGcgE6/OleJ7I4vHjp1OIPYWOrBYQCI7+Eij1MO9nifBjMPM6sUOqe91obygSE
vxOW80u4yhijiKUgDD3AS2sijbvOMGjfM+vhfqLFMlp4V1DG2cs7pordKlJD2r/daY8ocyULyXy3
9xPZUq81RZv1ZN4Eg++nfxbaqelusTZjY12ftmqs70ZKprU4hCvtxBY5HPME8DV9w/FaujgOPnK9
fm1qMrBZqBQxpNkX/zu3pq/xI1BwdTFWpVI2xrt7E3wQl0avo71JVc0co3ASNpVx+zUbuBNa4vR0
qQrpg1dlHroBhwU2NwnK37gYvQ2ziyzGTK8xCQuJSmsILc62U4EKT749zO4iLjd7tJZ7Jr+lZUxU
I4g1ECvTNQAHF1lw9p7v388g3IMvPRbUXZRclNVc3GRNO2dpR7YjEja+G06/x4BOPFxNqd2039u3
e4Tj11t9+3bhtMgxITZUbzD3cK+V2Rnr8eEyrCma+n2IfSr8+oN1rM08hLcOiufmnP4y+JwqiTj8
qRdEQ8aSJAw+bru0E+5MSW685rWRWGnzNAU5/JMAufBDysMY/jwyG8BQeZiigxPD6nDal3LQ+VRJ
ak2//i/TR+5km9I5ObGyP8E3idDhnbH8XZsETF4xv1lXszhcdnuJlBMDIFNiVq3yF5f70szzKJya
oIC0ditCQQQHb8sKQmUD5f8vAd3+oNJ/ajWDwhGyVP1E6/1lnyMgtbRRqDGOb9ADF65oC4TmpyJ5
oiqqBOaAcZSeUCTsIpvsiF8oKuzH4cmQXCo8prkmsbtv3815vift78oQgdB9Ao8rDpkOEVeBJ0MP
lt/GHcjl8pKJtqAfqEdX1anpYkWsTsBdS7nvGsiPRXmowUsNYcT8OSKa/cWxh+GNXJjKDfGgkqu9
dwDQeZlX3bQNPrZEJUx01heu228VxnCJbi+IFf06L6uQ5aXYpycbMYHl4KlsqOB5j0geoTNd+2C5
LeEln4nnpjuY5wQli024FdVVOCqZ9U4i6pP87o8eE9Aq5f8n73+HHmARu2niJ5+Wp4Wy2zedEN1w
OiwldKztFNXAx1oU2XQOwHxG/nbh2uGKF7qatzWxEvYS4phb4cxiSlPZ1tclyk+tsCyu+oFCoKLn
rYgyb8oArunHfLs3/qkfvJDsMdeZkDK1VALhdK1wsJplo6BEnaRJC1rOYogfFhgWY1LhM4j1ib6e
jXI8oJ3G6vrpOgVqmJH/lpdGU5iQxLTfmaGxZTkPq9cD02vSv365aNtbzJELr7GpiIYJ0eRUkfkY
EQVY+e8/ZvjrHW0PE7HIwN961zHbc6Vt05QwCEZ9LKKQsWNyRmRmsa2d1IURf79PYzUB3TY+mPO2
WWnUR6XA5HLI/ykOuER6eYSRMBmzI8p6wq/VW0a23XH0il8xUq81DMC+LH2aa/4zavW+MwDITc+c
Sr228iamSUrvNvY/q2449T2bYDhdQ/YSwSm0INRcuRBZ1QUdnvr/IXL9Ys4SCLebrV4e0nTvAltP
NTGyqt9kujI8/aM/j6l1XP9c5TrrkOR/QeLutPvPEGbwaPBf13nrUfjOyY2xfhqxYoGIevWgs+EC
NDvLxxClcUyCep9K2/k/jH28KkrZ6owInA1wuF4bSN5tWjp2M3qxgZLa7e1Eys5R5iwU490XkS6y
G3DBXfYEm41YXjo3DnR5jB1bngw+ib8xsVwiA7wcVmQ63pQwAGAmu3ISFB5mkzNN3l2AHflJ3935
jMlRlOgtt7KLy8CsnFvrx3qSTQIlvGMLZRCAyq15BZ41BzipzgcozUC9H2A0hDNoo3fQ1q4bQYmK
73JPKq+ZKwmDOCnQOrK7M1lpnxQwZR909ON4JsZpG+0FpuTU7VR3yVb+mSrl9UuCy/Y6vjd9CGvt
20o2lY8ncRyQkyl9r/VYT5Cdz+ba8Q1ToStvl3jicB7SERGZc7HVeYR0x8hooqXsZQ5hwkJqhxEu
fP4EMj027yLiR4phHL57VC0Xzqhi3rGTVfGKKNWTc9jxahWvH63OJC7wQ1/qk47ClRiOM8y0FG64
WhIwGZfulrUdDmN+W9XqqmH/00nUWPw6mOW+4bcg9AlTvydvwi8q9nb7XmKuD1jy8OxMn9eWafQn
HVDwQBycHlsLwRY9wDpKqXU3YRTKBtRhIRVD5ecGrznU0fcqvl39nWkQaBCYyqcHJ3Uuq+mzMBU2
713KeR40Cm5M34Ffmw47hqQDvt5AiWJaYnq73iQW6zY63A9bt/wSNn9c7n5qJk3bGYhY96WlT1UQ
qFgdBgJ67Y2RktGzsXt/jL+3PO1kwBIfwTESpQvOKaJmHyAvLkFYgJu60n4lFMylb9bFDeUyU+i+
jHmbcN4IV57VuJBQSocbAEAfcI2IjrzTGnxhLvzCuzWzPfEPEZoZ18jVYTxnb/tWhhv7p67l9o6w
ayeOb4yLM9HZ9wx2wJeFDDxpBPidBp/4U/leqm/4fYeOhJsk3PSXCnkKMGqhoChSkVsMyNKm+/Cq
OB3PoFW2ZUSR4bKtqk4kpXLNk4JIdidjpo9t3rOyCd1spKCwUXxh1FwEwB7++Z3qptoVtERqMLLM
5sIryFok50pUjdBXkgLLPUSo2eD3U5a1P6pE+giwqTKprRf0o8GAdklIh8UXS77bi86nFLLvVe5Q
vnQkGfPQFd/OBHkW5hBjBazD18xlr5McvPFUj8V10QkgA8leg0o9GLcdFe6SN37GDufJHRL75sB6
6WXUyylP8rpXlx34ttgMaJoYagKf9HnupRlAmXjadhMirAhzDZMiZ1Vk6FydWjOwFrme8k6Ha0xB
WYNT/yqOEqShI+N/5C2d5IwOr/FHGQN9ZbamBi3CtLSI382jpvX6KJbO0exjeJcenb9ged9WNwNC
1InpFSPaPc0lmOz3s2VO8FNkmLhUhPEq0pTGDs4MxxktwiB3JLH05wXg+jtPfbgJVhSsADzthjuO
QvIKhZ5jaSyuEyYEorGi1qhprhBm0nybGkuXn96zIUZEiU3W5W5izjcAFYJavhO7eeOe/QqZ6lMe
UNdKC9irzbRS/hH4PU9HJNDS4oc0frWX9JTZzPOBL5ZqZTJzLFwVRmNJ1KuLfyG4SjJcZmLFBLn+
pu62rwl8/At02zGvudWMlwqVwT5a5vSy0AC20VuyLgvbeaXgT0ttjaoVqYCRZhIBvBC62wDBaOYs
6nNkv7nKqVqCdYuxE4ff21154OPssItyArHljqsCqGhLP510RbUhIW02n/2Ds7jsLmkVamWTwcH+
1DgtM7UhyYbcjwwF4TyHRSAnVLKDCZi9lR6W6266kozfltHXm8cO/Vm4J2NbEpTZCJILN7wnWjra
xPy6oZ6YXzrkwqeKINBPzwnUtN+BwmLWE5uE275g+HMBDofgJ9dKRaWNmqFXxoyhZEC5da2+nndy
uRhJLs7HYaC65evKBzdMubLdpcG/WXzorEd6FuKQHbqDhxzUKX+3wyRWrD69vdhWitrY0ENVPHLZ
pQlJKbVGAjC5iNvy/4xcXNHEcRgXrLbn0afwTuaPEWelDI3mvPBnyIwG/h0K7tXzU2POOBwmzU7a
ZNV3FQM9GOzG5i4vLaUY+YSKYzmp69DrfTgh74ou/Fbap2J8wgbCY5pR/mJ91mE17dHWmh/HOTd4
dFkgrFV2XQQ8JKjQGu/gdnoDuCF9l+kSWE0YzXqSHa7is4UlTP7M+IccJBmbZTWTLGrdTB9meBcy
qS8P/dPMBvXk8EyYQgB5jQT3oSjgcZKPojfg3ZqRN8CNN3Mf4wu+KZ4xqZN4GgugO5wa38dIpPdA
pQmbG8bNRGKIC5wd47MTm+duoH2bheRW8AA78iv7jvCafMmGq4/TRcal0ut4RsCUF4ea6eSgD8Is
ryEU8CPI6H/o2ZCrz/n2ppR9wfwVE4qlkoHIu4+CVmiKQt5fzdmf+RbR/GBCDtOXb8ecrThPrlwI
JPO65KhLzmOzy6JBnaRn9z2yr/mP8ggXX5SPquvQiWHk02AEBbCKsS1ChLNJbIuuYaHgDTXatNfx
sA649Tee+riCI+/T3e/yqvus68k/4Ooj+w8I6DEbuu903nwhxiLOEBrZK8isyAXKMEDdaGQRhMRi
UBQa4lFC2/oMpCx6aU0R9bGY0ZUuyc8Rn+BcSa8kmx5AhpvF6TaMpxYBfOoWM8hOcQG265Yh428c
9vyXddyU06nngrMhx8phA3c6dmBn3hH+1LMOmqNlFp42cvnqHsGsuXsoPBm8LrlW6yFGW0SmdZu6
9uxOTSjq51HXx8fGIhStoNmlLRf7o5mBsCJ9kflfFBMY5a8WpR3S8t2ZFcdtoCtCk7a4Of7rLPze
gpQAISCsX09x0BBBCW7CND/o5z9kSox+8WWs+bP1gm0A0WUax5TE5HPONGtCb0CjyJWLT+P9qhMi
QHFhy1iV4JcGQWMV56kkXIXP50WftQVL9MZ4fag3vEq/jt1/YpDADr81CivT9AuDMHGKBEhUsrMf
2INrXMlyr8hBfz4wOajUYREoA20M2Z752UQifTIucnDTX37bJNiWUiy85SEknoSMW8zWCBzgMp1Q
EfyNMMvB5f2SkEVDxvqgQwtXyCTHuouWsKmA+usarYtrKgi+on52DtNN3nazzswD8HsHYSxALi3i
s2HYyCVwIgM9d0YhdQX3Tbgh0E5nOEakF2LThgXVnA5oqKj2ns14NZmGhjH6fUOCCtpKVzTpO20G
/ETwuVYP90UPOc/WgB8dueGgfJaj7xvtz0e6BZ8gRJxBP4uklWuUmURQ29SDKClQF8mgdj5JIQ/c
6KKnkXq5ICIcIzQRvn7+GWSAIjF69ajevZ2trciaa4Doq8OMuLu8tlFtixM4c1dRrRczmC10yyx1
1YArBHbcSR0D5D/H42nicLOaFu//xiUn2w6bNJ6NKiCnOsqQqlO6NzUkBrUNPVxRM17e6y9DOdoF
7WeMXxzBxc9378qxBAC8d+Q5S5bBUvDy60HabUKYzspIKqhWMBpa/nfHhCGnGxIOgp1xf9L/n8PW
VMzASPYBJVhlqevZ3sbvlZusK83kv2AogX3sst0HUUjqgtyPJmkl5NbzSWodVSXSBpRFL0ta9HAM
voS7FCnlt15mF3DvEPgH+QBrPo0FshqCs416z/0LNiGEXzdkoQe/zLpwInkq5y1iAOL1LbH1wsP+
95YoIifW8Hpt23BRX0s8FwG4+fZjPp6YrsA5/pwxCs1dbGGGz0H/s+c225rDLsxHwJJLDpmBQ6Wu
7/FoQpboK9NmRrjkWWNK77CTPUH47RZTgQTz/o82DO1MjV9IT1YepXtibSEqJ4DU/CwndBE6lfA2
T5Wp8rhNY0NrCHTrbTHKF0D7/p3LYz+T9zEPaI1LXHEHwrJzm6TSFbfu6OWTG9VP+StDdE65g3m4
B/Ogrm0hTFeyXtVDP1ltzf3v85U+yJN6zwHIwHbTgp5cayP+F3bS0Nj9jEDbaCxmu2WwkkoVS+zV
Vmgaemwe2+7O2SCjVTn058nTq3Wi8i4scv9lLcPF0Hrrev+yVzsIZKzBdgPw4q33bhkxc/9N+O+E
ygH76tbf/KQrEawIKJ4Whd6JSOe41lyF7JhVbFh3/9/UN7wMidqDumScijv9K4EFS0SHNzYrRsjZ
oYk5I8E/iECGo4fIMZM6232qYfRSS1R/MzGws0MsXCl1KYHrKuKD6VUzxkeWY0XCvPdb/+nk2/8x
AaIg0JA11Yp0t3St5yApqYW5vKTzc4AVAusE31VrbNsyYMvZvdFgXlksRj93SdGf8NIDuPn5HA+4
FgBf3jVot9eR1RIki6b0n8jii/Ak9/KifVb+v50Aaa/61RdDP+cSsZEZdw5ABaUo1L7j6wKTqQz8
joMLozz/RaQqozQG7Agd0lXgd6EKu1VXc4cNU3ieddj55u63Ug2iwlqHlQyzt9gNQW4CXNzUT5TG
0cDl3IdWnEhcAYtiEveaVW5S++ipv0TsFLGP/ZmT+63+Q+n2H5I+a7PjFc+RoQtJDQX56HYyMjxn
/qC+H302CenNErBsur5rVKMp+BoWhm1H3cxQ015kzEIZd4fxgOWHBf8Hudih2s1IEmhWOuvP7Q00
LvAJdZmIWcWsxIEb/8tuP2q0NEwmEe4v3/hfqFD/u/H/BmwtKQQGLKQy9kGq0YX7oBpR/ysBJ7I5
ynIqjUYg0IAQDSqSbWzSDDp3VGhaqHTGrb9iN2P2gl/fZyYxg1iPkq3HsR1TAF21Xl3enUaV9ThD
Qydmf9W9U+y4OKArgZ9mDUMsgvK7AQRRkMUnbn3AgrpbTbDBwEOgyt6r9bJuQZnk7vkPQv8fmAvz
2Ju6GtxK2kzJvPwOaN0AhDLHOzUs8m/GB2wIm/+tHU6kqRm8xgiR3Ny29v+nQ96UFg2fTflFwX2o
E01wTzOwOYfOqiObQUirC6WoUnl1YXH1CbWxvpyPvnTtDNAO4Ezir1VANcuUFgkBcZy2JivriazX
dJ8UuFz8IRurtDm1EtNSslk0Fzj5OFTnNMNZQfgNDubAGIJL03vrNueq4PSNOfy0AIIvB9AQMZNZ
LXlcEE/A6B/pvsDqfLP/529Wqg3OJrdXLqMEKCAm7r0h9CVhsBbvdiaVsF6raUKjg9y6SiYNaqkK
wNZsNyYQ/rkHA5eKhxOfIaDc/80uq0Y6oP6eGgHuRcJ9eRMQIG83Th3H6FlVf0YTkKebXszxttJ7
VmcsWCmXeOjCL9d/m6d/AwkwblXi0toro+ktQKMYrxrxFlZSDkD08NT8HWEBewmfnn/0uP+TU4+x
fEGsnOQMs/Zpl5CCUh3zgbAd1xi5nxL9lOntAlw0Kl8gReyHBKqOJvpjNB2pkiG3R193qeN4vEiO
W6jGnSCtaiOgolCyDDCfzjlMzZLmNGUxKmZ7bYXLcTSMbresnCwLqOTyEjPnzEeQXqqV6NvFrJzr
pR6Nc5yFd5R6dyc9FvcvzXkevs01DEsdojYDrY10G/yZYazMPhAOQJFCpVgRd0/qEojdtzHgRuyS
tXoelFA+KMSBNlSOleQK6Z+VTLy9Cv5Tk1moTGYEip/i8DhjS61KicBZT0ftP5qp7/hDlQW9QZV1
D4ADGz5EXcQ5bSeZj55QQ7UaHiddwXrLGaC5tmsEKN1GLacbUcnBDXYY4kuH/rZ4p9r3MOKG5cw3
9RR/RnuRAIJx2SNi9a8EQUy2KiwaJtWwWZJC7zM1X8C0VivdApi8MAV/vsv7fStfvZ60oaURhtci
iJ0uPSJfugrYEY4lwv6dW5gF789Z4r3Lwu+T09q5efiEJieYyn3pqp+nDZNj/hINOLig8jcw901A
Bt1t2GmKvu1W8ASwxILU/d76OZGHW3rOcy+tflpY+4yTPd4DSixxEd9bdU3vp58VH4rIX6am+AJ+
Umfp/1O8BahAfJuminhlqzd5hAQwyfv689320aO9jtjtnvlEEVU+QSevfT4763G2ETp9N3mzqj+p
A7+qqIBQtiMnMBRteKBn8at3UHB5LIF7d8fnoqymCB3hE9EwQ+4pje0zaPgK9VEwhnbA6ax5YbKx
p+HaJyE300nrywrMGEZCmtAPqpo/8bV/epnKJ/yHkIhNl69e61VZ4eZNSc1yYKiLwuuWlOdSbrdO
7h8kvXGe9/w05MsST+4gB2xhhWs7IZCICw4uDq3+SRJpFy1fdxHxy0YOot0yfvyM6xtm3gz3B//1
aF1c5k7NniE/e1j0GTBG6levX3tUMAMeT4aKQvCiDr07XdKcpfo0uOT0G9d3B5UNNuJwx6/KIb5D
OnIv4tiTky1h8EO/y9pWK5PIMQMDOkVxcK6VT5ib5MUw3MWm2o94YzPeH04c73QX3zCgOu9CPXf8
9hd2Omsv7NpEEAe1hEoOts/C22UFD73mmKzYkAuaueTreV0brgNhS9WuAw/mE9cAQAIHAJKQk2Ov
YpswR2KB4ZrT9QSNYNOqB9ngP4UoRuKip5ox4/xMGjPr1pEY2qVjZu462+YsIvs0PMNsWAZZPhEc
SxfiHzLqdubYoAfW0kPyh49XzL5CxPSBk734NLGO9xeZhgRB0zXFMAjc+2SI8AZVFTPIL2Sbr7Nj
FkYDE4RCG0s1flwm4HYzpi+52+7ynqbHlmk4pL7fuJU8mKWv+KVTJsEPpjptSGAdnqU9eBfU3fsB
W+2GYgjpIZDexzXiEQ7+FM9+jt+tYZZqLwIYFj0I9T7A33kIQxYhyUBmbSkufZiEvXFIQ50HY/hp
FWaxDPbAYBeQluTuOjFFrICwNROuBPESy3gv+80zHZulWeP2Hcozh1BDCTLICONV/i9rA7XPaYoS
HPyuhTixKBWOw/To3uGFNLxtbDLAHj1F3EKSSHDsq4F+TYO9gZd0hiT+8q9gb6icCBfvI/cNJM2h
x51ZWHKbwypO4fXjaZjrBDR0Pcjou+WEvSKh8CFQQL+SJpMhvDADrkWxqAsImqBAbCjI+Zz0tL3U
wgTnsRoes8Gc0WxADmhcNKHUgFFU4wuGQS0hiyrKHUSRXADIFdp2mhHpGyt+MN7VXTTBj4QGwlb0
UgvtoGb8X24+9cgzAwjnd/gHN/QmYPdiyhQfTFmJOHqTp2eKi07yCeLBqDjmSUhwDqxpbxtrefYi
xPH3Wa+neQp0mWQhQ0992xZag+2DryQIvswqwn5HKQr1gvseKqwNFVoA4TuYTQpyybX8yJhzW2gw
dQ5xudPlZF0uU3lPhLcWcLDfTDgOcUC8CRRpqB+sETrgiLdniygLn08LE3vCTCe+dNEZUWF/LAqx
x14dwY1JhOh4notteZ1iE93DH6KBWbzbJOmivlJS2fgjaTnHYKKhr80KwHCgEOSOTeAoa7e+nM2X
bkOGzFFWG9sW5MgoU385okI55CL2J64HzELNSP7QxtEnzM9uTJcm64OLjj1Aig+MJ9GoEtVP59tj
ZEadkC3snCEUWb2OMZ5VlezZcqpMpzf868puGQX2MDSF7N4aaMVcq+PGd0gnVQzr/cxsprta9+ms
hjUqsP5m6yHBM7T7q5NDlcyuCnDhZJzvRzLeB2XRkdGBw0ZTg/jZuHXcouFkVOoZdFbSO9hNubgT
1810NI0+KlBhcAnJTz/XaXFODk+OqLhotC/dn8dgrOw2CZDp3yqYMSysJnrJS2BFU/h4D/WQyiY/
XNwQq4L549ih/bKPb3xrjK0MrctzrTS/0OH4To2iSYxIFIF0X7hRVyMe6EjEu/yk/C37df5Udybn
lEdUYEwwKkCtmK1WhcM+S/DBTKsBpdGUg91A0zpKWZarzO9WIk00sFiBd+WWw/p6g2oXKs+63hCv
QaFsPJiB1ViSUXwUiIUNO3kfts1WiF9/CpZ7l+UXZ9S8wv1kfhBXC/He203TTWrj6+zCX20YT5e1
mOc88xrMJ2jEhqD7CdVacvpWoLoSyovosvC++UPAKMSnyg3znE/Uv7Zvxytp2pqr9ZSXHUC0BwgG
tg4TJPd6+VZoAHp/jeT06N0tmKsdWXz+PQQjn9vmX68hciem7C2+Hsl2TIEOjQ8AUBSdo5lXdDTX
4guTSFkqi2krY3tMwmAvgKzqKP73GWDIszL8jsnBsn/cyHvmKSX6S/RVzzHZ7HLI6I/f4GgEHICc
3p2xYkrE8u+pBARJJeFWxxB7430eOR9gabmp0I24mK6UvZ/55O0Z1eZEfZy99XzbiA2iCgkI+DmM
+4+uKXGEbsosE4hif3smMRIuF/++7eKgmQtoL2hlAOX1TLtCj+EcGoUEfblRGgzH2itx0P44OlZM
VZ6+5N0qHPGXjcf8iwD0fFd+BLGCmSgXmtfUvKV39XJOQo5Z6fD1fnZf/lWAYIuwiT9HC/DwKz0p
fUZb0qLpZKYNOdMdHdpdUs1ZN3hLZaoVMuEQQ6U5KbjenC++kUohHhdYc4GKRErDT0kLJKV8vm0W
MbaanS5Fu1QkZMYZ5+WOJfEI/6vWKGm2/JF67ZnHCXPRhpsIp1eBKh+2UxMqriZXexwoKn5G4wuD
ZGjZ8fahexOISRpPfCuMlUiyosQM0Dv3wXYfuvSdR2MKZVaLx52SKXSMXwMSTc0XGiIDtVvDvK0v
uu2LYQ8266oGekeghwJBJbhFPWs8U4Fdg8AdyiMySEOFjoOcOigojNcEfmGCaGNtXTaD93D0VN1+
3WRvn842eJfdFlmjRGn3/Waedt5pz471vTywmj78nI+hDpqE4MjQ8j4yQlwj4X5IxE1RpmuQAHH6
MGFhbYUV9Mual8+cDh3R2dVyNv07g9YVms1jUjikjohUHLXBwNiM1H4yvkr1Is7Ee2pIy5RYfv6I
zlruoZRjvzLBOPH14yfDsgk+U3PdHGA8f8ZgYQX7je3uOcoyWAfxVmsg+nZVQaLyggbvAO+dJo+Z
zMBaEBhufKUfdkjTbUuGjRMhhTbaYWcAwGTcGPvQKYJBFwKD/RspS9sM2Kac1t8ycUGSYefkhdyw
Om2NyYf4C7aGDzE9ufYhYCRCcsULS36A7gnQlmNTnksyX6tKIhc/mm5RjMdU9h1fj0Ep/ZlULnn/
p3G6qZxptvS1VGzyFhCKNmBkyntD8domwTPcz1A1CA4DQsnxzjNJoFJRi89L0EQo/fzw4vQQWpkO
SSkrfiH7Irb5dDlHgtSun2Z5tzqXNraZtUpeq3Oj/d+i3CKWriOrAz6bwYvoSgbNaxrgQ7pujMnR
UMXgnByNyoYeXhaPHduzaYJQY9DLTAn0i278GauNKuxoKEFle+vgY69wWqtOcmlrhnZD1XZVqNMx
c+tTaorq96AaWfUfTU503Tv6/GN1Tab6NyxHUC2MfFlV5RbPdwLwQAMe5FDlz7s2XnOxva65wD57
1kaMLkPW6lceYcOAWNBPxl7wxJAPFmAkKKlJSV4IxBomB1hzVlwIweeXLKwAJk14Wnz6N/uctxPf
sz/t93xXTXHfjo4/M0GcL1d0yLTGoyjmNLKs7C62U5Jhi+cfKvWPVunHPwY21yMc+hyKZ33YZXyU
eZvNvtHvxAWH1aUxuk6028UFqwIJOz+cGC0aTW7tFS3oZDO8IS0QZj2jCaTr6JydQ3inKHQXRAG9
v1b71MocWeKwiOqYEH9+6EanU+nazBW2z2vFH8qjws/K2etmwFryX2AHsIyacehP/QyVvg2hFifo
zZ28CQ6rr+JXSWrzLMdjRaoFo8Qcde4AVH7zdRFUX7OmpZu2+qoWWt+T8AODQAtVMjIcYKPW2pYb
mq7jsLCUTpmszHfXU1G1IoIXsGQKcx4HbuzZY1TRwcQX2HschaJHsjXF5XLl8dRsO24bNJJBqqjT
kKNbXBwkuSfAdNb3mUon/znFRYDsdS6B6YFhrdfzPsrHJ1Oryziir7dLHu9jb9IlUFiEf/SIdmXC
uwbznPgI4zbI73OQbKyhjwVkBdKBStmNsWOS1adAgVf4p7eYPVM0Q7c5wXNdKbWAP+RoZoiePq9e
sY5x2CR5o/EnRCSTYS+z5oadV3qTamuNiM0WIwN4ybXtUd79aBa9eFCV6f6E8QwsedvV0Juy82DK
5T7+S2t+9BefkKbrD5+FgAkOyLmKwKJIKGg/57UFUpzE/EddubnjZIp/SmjP3Nlt1dH/d+It/PJW
dA/wM7WNtN/v+RsHZnWCTwNmCJIejaUK63A9oEjjVhBBkrRjyEjPO5cCxyRsGmmpsXLW5ZGlP2Lf
yq0lOGKvObbqxD6689EHI/xmqMpd1LM3CLPhmKsrxhgxaVsuNxIm6TwNIZvZL+7dgrCZ6mkF6A6r
vHpsqAqQxWRJn9zY15cyqFGEaGj/EaWghxurjWxPO8WvChITktznpFoX0DcsJAqIHZULtN8aBfwN
ylhwU9c2gORSd3fkzix1Ivh7J1x56Jpxhvb4RiBdiEsR0+Ncgs39ghXAACnmT/CnbMHJwkI0YZGk
MHQBDdBlygAp4VWHYFmEuLihmgfxY8c+pj+jKEhK7zGs6hvoa7iw+sbxhdHG7FxkusCarUPVNfWe
DOL2iR8areGRHso29tze2ZKo5LrzCsVN62qDf2FxlrzwU4+Tz2Nun5OXaJ6IDKgP4DPATQmDa8w+
BrVmWOn5O4jg02E2JxfSZCxq1/F+4CZXQ4CJ8jP22uWwCPWH5LhqIBFuYjklFPbisnjLl4JM9Bmz
XCs+ffNrGzmt9jWbA1ZdbTISbDWjSVpbVrIG20bSX68wklHeyI41Wnp/np1gMJd1MLIadqendNFF
aPJTE9H9OP7RRatH3RWxHPGgOaAbQHuGwMJmlk2j7S+zLjHVlaL/q3lzf55Mhlrp611RuDidD2Ls
BQEMptjvqXtT8puExVYWs6iPVeN1l0AI5OTQjRmCdvye3t8pqsMOf0vrCn2Qn+L3pyRaGYkwV1d0
UYWSBhFWBecPXSYVzkQUPeW0KaqztpZU5j1Cl4sU58OT8+4X0HexaIfvt75HPMrVEgIX5Xg76KHm
mfKl4vwvX8FhXmbxgIyy+nTe7fBsqzxUBj38hGJj5TH6aWmoqeo9CZGYjrnvCPTl3A5mE9HogDRp
b86JN13Gr4v7Oeta81Af/uAAMS7NobLFSZRDmMnQ3WoTswMlGpSGJl9CBBLChytBk2t754ZVhCT4
83jLZ+u6u+9HAnUo9WY399p6Ozh/52hk1NKXF3ZkKN/8rRiZNB95xkS3nCgxVVPgh3INUB5aNH/B
uyCIcvlzGKYz1k7cvB4geWeb3Sc0Bj4J0xu25bSJ+wuYZlWLCLsKZ6A/OQa6RKfaHj/hSkrnL+4N
AWsGkSTbUEF6PopHSxPTYokSX31gUacgDdEXes6MeccH0Ef+ur1y5LkpVUcmh0A/TbCAeL8ysO8s
n5eAeVOocBaEX91438VxDVMl9jEXWx4aGFnCZSZ1FSroU5hQEX+nCKZX0WwrKxAvBa2tYLzFfmuc
igLoVmeYayesz3qQis43f3lRgwhMPj26vLgCA2RddrdiXbb18EEtHH3TlBLCvZ/bp7TMH+V5u0kf
oVz1xUfpf4Q3BYqXnI3IvfgiPOi+/Xv7zbjVH7OvVird0mgWjJR18XVIovOBGJIEPWul77JWxnmh
WEUoPKD5y7wodQSyWWuVKpiznvADUOkVF/1nTdKfwoACcXqNdfi3wKzwkmQBcPbwmq4oxcWoG0bd
cqKMSaqqw2GJaVHkfTM5rmV5mfXaUE/kA5MbLFCuG2zVhff7LXoKEgD+n+/aUq3AFAmQ7tnwJ8rW
FGYmR6kE1lg1420GNIhxw0E9xRzaMV+2mm38UqpYFx4xeQtmW53tXa2W0x8xiou2uhj8QPLXzja0
9NAvXxxZ2t+D/a45WW8z1gPXQkPjE5vwolFrDNEfs6J39PI4sbQWM1Y69qbvtDi4qQzHxfRIZcXv
QnyQPGvS78TI7+IU2KlmGhq7MXcwbm2X5EToLn5mkH3hQ7v79gg8zbNKSw7iq9v/nRoguhv1G+6Z
9RiqbQsWRvkfw0shY9aX+IJAA2qgVmtHtKibUEBuawne9/kgvL6zvaN7NkDKSt4bs4wgLUGkov1A
wyO0XgovotfyMgtNqTvn6inM/SWgVy27Rlx3aRfNe8g2mStd/qQFw/ZdVWnghd4jnApmoUfenMtX
RXWKC2dYK4tuZvYOmZ8zNPJ+C9V61V9g05wwRZo7W9YKoC5xeu/ap82R4fyHYhtiTlKn2QGRRia4
zlri7opqtoZl0zGSNgdWUhTtFdsHU1uGNhV846D7PBzXrx4mxRJgWfjjQyq/57PPKGfEqNFedQAh
GtUAOBf1EneMHvMTzrnktXneY6WcZP8KSFZgdQOw1rsRbAFrS/5ac2uixqsOmFkJ88QJA5YqANTR
oluaq2Yw3sFDroP2XLSA4CxO+MWxs8CuaIm/P+tnT0O+lpoQOkJlu+Q5Lgh2bGwG1U5xsd30cZ9J
jWQDdN/w/bnPOe3ZZ5ETWpHGzCPQ+qa0FkYKTaNbqojqVq+l81cQQd0NI2VRGpqI7sCWnxDqjoz1
0e2/XqD9TO/uU+Kqa3Ix3USlokWCBCBK3WCgsFOnyknaU5zhpkt+OFoc9z4KGJnFEx66WEX9n/Nt
t9SIfAZXkArqircSo1Y82M29GCL9NRm33meX6Gu1S9nIa0S79idYWYxq0IXfi/YuWtcXXkGMeEM/
7N8xhyZQYguvYGaa86tr3I9/ZQFKPFN8OB2CsL3Sx5vB/+UHSV5/+dfL+4uSIrUfnDPd3frxO8yg
xmg7jF23EZ8Lf0AORhGnjsF4ZzAWzMB9LhYn0MjPxASmcHkQgogQCEh4cge/PY0udKb8McsyGiTA
Dk2ynEkIHkqJhvspc0jWH2kSEQDeBASGNk7DImGRq1uGatAuWuCnb/cSIit94uNgVShRaY0kqSJD
FLHbAInOPRW22S7pnueo+jI1kmyZjP6cdemquZtTqtoVl+032ZU7b1jCG++pbLYpbcbIFKz92zLs
0Ufkqr6BBCUuvx/77KrXC81i75fxtezwfNbunyNEgOlKzjwliWBqUem9NzWy8JD8728sd+A1XyQS
hEZPabsTD70a3TSg7sR3MHhNXsYcUivUVJbs+olWK1iUMi0XadmcXIAuehuXxwr7KCJ5aYJ/ss+w
YRTnPo0X0TGtpb5YzLDDvKHgQnru50TvHowckm+Db6/z+KfOjJuXPnz776Sn1l0hhYGwT+wRbsi6
DCRySTREtr9IG/PbnPbF3v83KnCYoW4IZBPP/BcmqcghPKTWyKH7O048LwieIFd8UZ694M/unMGZ
RgJLqc37w1Ong/z/YOWorUbi+2TWqbG2DmfJmfpyAGplV5iLZIW3qj5vSsJ+CSR2w541wFZiMmDD
gQuZKEf+0Sc+KCCr8LxCpKdoM7WFx24WDNDqlwMNFKeYB5EgMbUZ5+oJN0aP90dy2DVeGD/fPm9x
MLt6PPbN/47jEBxjz25Ai25gTY0+gYMv9cItBQBE7Vw9x23bQo35n0jHaxHC9DHSLaNoB6Q68kyA
rPTZDeozqfx4U1llcVo4dcJ5jAkJP7/au80+7HuzqdGlSRjfc1efXNOntigUQcRRbB2XRW89W9rS
/Pzp6LjJTk/kmA7gZ25dbXQ0db7TaUA6UvQVWq8Kv90DBZZSioaLVFxXvNbbEjHlWDCzG9z5maPo
gHj30G6hZfFuG4o1quusyUO87Ki9FzzP0nX7qg0GRyQGnHz6s12HjEzlSqK3qIZp23Sy4jZnkkJ9
tbhCSQqCPdoG1Ioo7vHDBZtIshhwg3tI+lNjrSi0DVJNpKzFyA1VZ/VacXVKiPnCNQhJndsOP8Ei
tKIGuSuISzu7TBzFFC0qDcyq7rvgwwQhlKbNCvdKCQ1gDDcZTOit2MNJGx+UvCbSGZJvxQZQAbTr
xQG1TWoNjk2HSBmz3MFppXw1FN5kt0WrFQFFkS/+vRJ1ElPMm2miQ350gN+OuPHQpTcZ9EYVMOJ/
nJSZ5kGTgIyiMeTk1RpVRgNo4TaU8tlRwr2D5bsXjgTXoVezkJXVtbQtuMMXrLqadTeYPQHjqYhD
blNSuDn6fb93eyDfhwi07znAeoCOiVxn61T4iVv7C0aHRL1PVEVSRGvb35BDvRXtyuZm1sh+GH6e
rXfGqF14Wv0PGFfKiv9h/RWCOiYzEsfzjH2Qujxx2VrjpAqPBAJsgwnx8yzEmcmkUdGSv3JVJy87
kqSSi6+3aPNiW3fkOKBzfDw2KIng7RhiFlQ94M8LO4tPRimwaq9QClWj6oY43TEkzDz2C6JZvun9
t1LTdmwe92FkwtdLnfhZCF2K440816KWYg/VH4ph+XKWY1TxYy76cSvtuunr5tUi2UIuKs3rHJdS
IHOIrI8j53ijWBai9AOkbJZddcP+pWWxeO2KxDbz1hKIwRbYs76XxCoCqqIymr2ed9Xl1Fm2JMSS
lcFb4YUo8tLS7kO5OKSr8Vca1xeW9jlH0xC7oD7H1TNK8KX+rcbVXkgPIv1M8JewBTPoKewafWOD
nnVaOqcCA0OKyKiGC7BxzSdITDu8dLDyeZsQFY+GlMXx2qsNi9Y8IV8zje+HGEWENKHse1btbX6Q
R2IcNSdnDZIGgUjS+RA9t0Bv9Pswpb6yGLf3AZZw5hQwuKgZdh9erNq3QxU4tqXgmvZfaWaCkL69
w7GsuNo7eNP5UQjyqwm/np0Eio9KxxirAYasbLT2eVno95xtn3SEuqGlLndOpmZy5YNIB/u3MxRB
8XrRygnKtwndga9yJLJ/oGpcaK0lh4/aWBM5mLh0txlwBdi3ppERL/YeMsvdJ0KdUPhvcCrQhQix
aYOhGhmukh6+k399hUes5gDgwmAsw434leN4XDIlZAD+RRqTIXByGLXkyoCB/Vo2u7ql4M744G2c
mzupcF0nVvwqba/PDx4cQ1BWmuWjuu95Bo9lUqzvk7OwFWvYHHZSNvtXfbNcwuZVpQe6XtXfaWfW
e/qXPrKR+5QjZUjIlioqW35RUFTiXJYQOKMtJLZi/DTwpvoSeljyLAx8u7qwgocA4LJJVCCmHI9u
nrmAnISeiaj+ydUh9HXY9+pbdBWIEv3wQR313ib/MKSy3TyotRmFBEGH1CeudOQtheKvWmbOaJm/
dnijFrAxWGj32ERqXdITJbwDx0hxhz5WrY0pyLkCOhlPLPhKkXa3PgCwVggi/7Jzi9J0LlwfJwBN
GyZcZXLS6RK3adzDVZ1KLYHDgNNvF88QlA6I6HyX/4bfqExbXdjcMYhYRzzLQ6TthKGFFHoHqFUv
TzVGhmH6ckyZr90so9b/MEF9cj82CdU8iB8ejVbh4OXFrh7Uc5YxtEyp5QWchB3A13sGDeQWBJXV
UquFf4aFMxF9PsLSgLqWocJJzxDwfzGNQbanrGXHwz05XmSAzUKId+BfhoFGPk6EpqPfPab4Fh9D
JzlpmnFvZ46CNCZW58+EKS/faXTXx6t87Snq8QdTtvwsLO4WlfnDkVZhKg7Ftrh4v9I/HgnGpzbZ
AEplqRJ/uI/ffa8qIO+3dD0vt7HfcjeAW74Z9FuunnJdYsMqEtNSFA0EqU1IALHkugvUrj8HqFDi
B1eFFGffNaM99bXqWRE1Pr0VNsIb4FpJSyUYdH8ETK6bw80MrqPyQJBcElLm12wunw/yfBPK4e5D
77qgZ/mpM+fedr0oO1uL7wIoDf+TB1yYQO+iivXOiJTl0A73PZDAj/pIjiMFuOksoKWY3rVlwGGG
yw4ntSWY7obPz/JYyAJR3pp3R8W6BTI+XLsSEMgnqHBkJUmxXbTTxxEocki6eJtoQr14Pum6trKs
FMdzcx/BY9iyKQQvCOL99bFyz30s/Axn9AXhVORjqV0jHc9E+xyD4U3rNvFPO2mSuzMLK+P44Pmc
2gqUYA1eMWTTZWy3PGgPnDRMnv8TFera62b3fGSmAfzwfu1xJdK/VilvfpUvxZ7JfE5WGKT0dX9S
fj+R4tY1ANG6NuX8qd3yONjvB3sxT68XX3tV5Tvfkas6vWt/1SEjWOZgIhvK0pr3rs1eTueiFapg
JnEbzcJMVIwL6/fricFohJnneIpQSZuYcsMKy7ZNpPNabr/5mfBUlgGfDFSCheE+46JNPXJ7QS6R
66OTLrKiJAXHtTgE1XvWOVznJWvkEWo+4HYkP88/ovm8HZEgYzij0LhxBf0Ef2tAHjjQsKnmXqg5
+vQ2as8qGtecdqAlrOMDynToRzDKmeXm8mC9fgbPYYeOLKPJHRN2WxckG8YXlSDVYPCD5aJ7qW6i
E4XkKhw2fOZF0vbGJ79wkbgbeL5ICy8peKrKPlH6wFo80igMKm/KCLv3ZJFTgHt6iC7ZF0ZzgClD
uSEKn493io8mUXj8wdGFmOx/CH6LqdNcbLlh/7O43asPTrjTdqyaXcGOd2Donv5uuVQczfN9+PvY
zJCBfwUlOwb7DurPaRPSYY7mknkRncmeYObHQk1DnsurhQUk5oj3sYI+YMpaqCrzRb2ocxvJAyg5
io99Rogy5LDlOL2sAmKA3BKRRJ74PLChaz/b0fkxarTK6JU1QephgnmmcLg00stTDzIEzB3Svyq9
/8DqOjVFgtpAaVhVBXE7qXvVvIAzTnyN0yYNExP+1UN+MDNZUfG4QcY7WD8t9g+ejCHTWtTFle08
v75NaTZ6vdbCDjrWKY7AWgz5Fa1vLfCxMjmWQbAZguZKenG3v2IUO5JVUeiXDoJ5MOn3LCrfrSH6
NNCp19H50CRxATbLU/k8bkZihU81JZ01TQM5LUvuGOBWXF4KRnaUgy3VoGoEVMa3Zxajqcpx4FkI
+1nznXpwUHFcSAru+Faa9N5WD8cqmI1rqQyyKaAtoCPwMye1REqNSaLG4E2/0BUB9vvZIubNcgPz
7U/DSIavRgjeaJb1JOedLKhqLQnJJNbTn4q3PifMHXd8VODr5wNRkG6ZPmnj2scPCCWYypHl6bt9
nfd0E6CU+AtOA/1h/4pxLJpMXVDOk6Iow/VTsXWnk+jTauLLuzajhLRItFT9guTQ0Zqvk+munheM
kfiYwUL3Yy85zosw/eD+VGAz3XCyiWvwgmguwMftpKtnOn4ideuKq1jONWpxABbtu+prEbLwMW7Y
AWGBLVoXVT8pR3yW5irRTCfcwQMpgJZi7VdoZ36O737NaA28gkf4x8psgQENGPnVj14ojAtvr0cL
/nin/OqXsfysPJCd120m36Xs5jXGlMKs3QBFwA6f4cIIEUt8NfQ6WEuogwRFfB4fayOZLQQ0IvsW
3FlV84QOKQGBxrL5Ki/SDfZQ+b2JR6R8d4lPv/jFZhaofdktvJJDKHiAlCGGo7CguSxDHN+3QvtJ
cijW1xQ908BnRQzg7W+v46DYJDDJ2fN4z3mdp13ZHuiu7yjMgYfuXse987EHjKVEkZP0IYBiA/VV
PDUxwfgoO+4X/8JJZR3WQf7/9AwPu6PTSHzLlp/qej0qLDq7au/kX96e9WMo/IW7IntK7Mh4CBO8
SOc9z2PYmK+rrApn1YqYmesgTgj5+KvILxK/u/mJSpoR5ArI9/oKxKNqikVRjkiYqF3TG4BAKUOz
cqBSaATHqLkMCjfyEdxQDuQcFSq8sHTVDLXMr0b5Lr4yQl9o7VRKvhSl9yR5NwWtNhJGTQQ+FnrX
tTEjFH+GsWh2BxQla2AXt2mlw3FM9qw2Dmav0oj7/maSXWeGE2LLawCEwurXlaB9QwBz9mTE4pA8
5kKwmgCcyg3SQPF68U4ysapa0Z99f4E1x4nNBfr5ABOeZch2TKQqMTGe8jZ6edGGGxF6lWyIggRA
FU5h6ru2OBJGPH+D8Mm8rvDHWM0OV1M0KPvTTJTYeqepZsemKo8sc6sHEXWeNYJzrGXs/neOyg00
mNOjIPs6IYgXOsrPmfSC1s4en2EdpwqTxrpJ1LRbRexfRXSQ94WXCda+gYiMX2YsPCTwo1Gi6duO
zsofsFUNVF1ebwSoTGFHxlQexNzyCsb5tTiiVXtDpS936gNHpUbVlvS1w5nppCgRYrdz6+fg8KkY
x1Po0hJ0BzK5Cd6uqzRrex238UuB2S5LfFlfRItDNPpw6YI9lbzUN8fvLZEkmEYlGW8uv3nwwYM1
B+jUW+ePsGE6k6O/f3lizjvBHJXcrWf2pnPL6qzNwmKixByUgjTf0Hxn/jzoHOyDI2Han71wE4Hm
t2n7wD3cFJDcqeQ//M9w5wYDQeMcvunJ6m4uOj6HLrsOKG0sNu8/hj/lBmfT49e+U7VEcLtJI+B+
7kQznRYqDsW6q/DVZb+mci4z0R4NL+OBRpKUUB0wyS9sb1iPaO1FI+v6pJr5Bt4T3Z4bR6OZvi98
dtJPpYBAW5PBg6vkp1MQJbnpdIF3AYpPNH9u5sJxy7WGd/uFjYPZFbta4toGxzU1hd1JzXV3PX9m
iuePZK3gkMVnSj6zuRwEnXpoGHFcb9LbtPW5GiUm+P9kIoH2JsR/QAFQ/HjZuEvifbGKmnozv0pC
9WpOEAJztxbG1MeKnu4fb37i27OV+TCEafSOW9yitkuNnsjLaBp8sBKGGNA0x5lROnx4PNSAnCud
01e/fcjXzQoO7/rO+u1XOQvDcjD0E6MnpCUUXwdCwUtFkE6y9l3yNuf/7cU3wR6RtvLcEdKZcHgF
i28CX/BPX87By6GqnJgm5/3Bkfl+gfFqL6nMIrMjS4tgXSi6iMrdTzeeHKXpgGGxJCKgMPXJRMbg
oBLCmOP6+tyJH9H5PLkaMNG011XDS6s0NHNjtR3R9eAUznAfVEXaWsaG4g3HQTCZVeRP2HPQfgiP
aZXvQbF8So2MHXnSxSLFnLGHYkS3PHBqGkl4aKx3rM2PHG5JP4O4UnVLWAXxBBtvaisS8CiJmIcG
O13Af87c054XElPPSl7eWSbqsze4ZVwCnDOOnrnTpOWeCRaAs3ExJjtp5yGWdxowDqj6N7QDlnX+
yWaxBktKUGnfd7JQzK4B0Y1snLSUZ0T1fy2nhgteEWkgHLIgH5RWmqgb7uj5PNL4z80EaEpweah2
WKNxaeaDI1+tcGqhCcBVAevwFp57b9zxNtymcXKZ+K71BUeHauempQ35ja/MkG82JbG0szh0d/E1
91ZmMq7XOdqkWcYWNRepRjfauf+bOl8k0omzcXYLrMokzf++6uJj8vzasl9EDt7+P0Wp4OXuMAnS
CUKgDHDKmbXuv1gA14Hy1dGz4x2bBA5gHMUZkv0TbLzsKXS82Hrn3xRswqrtyC9pw5V+eaiUXoiD
pNUVdPH5aui+G4QHs2ehdzokUovPe7ED55Hhy03hjhpBBIgEydvgBF1nuxjM/Ms8zqvR5AN+wyoJ
sus5soAlUWdaF5BqHLlysAiXBpYlFuDFvidMxEx9vIz5YYYY20iBb8JCt2/REP6mCbjJSh9rGrEP
aOjh9VhzlZJ9PG3ylDMqGyTNE8IhhxDRiu3bjGMSgYwXg2tIYxS4L8lvv5zsLGP3jX75w2jqXQbG
6x2+fwqhKpbhBgWdxFX3u0rnhbSCm1kejq7oqtlTUUQ6hOBdT/9gZ0Rn8h0ozy0yLn9GkNPp/Tsw
0H3BWQ3qv23amYAwQip9tbRyZWlChTMTK6nAfzsAHqNc5P1XQm+Ij3D1K6TNOEZG0AGdj3u+DDcG
ROmrr2A9HE+nywfkQYDkoqcEyF7snggMNqcNiRK+zTDyWuxZXIV/wPuBXUKA1aj0xPJ4uBh25nAx
G6RRN7VD1VS4OI6DZ0oZFRhBdCaz9AA+b3O+TC4LkRC742KHpmc7EhtTzScakMCjxLmFTY4C2+0K
Wdy2yFZr+LYvh9JXATWUg/WdrYP9LMhDAzSlReaFsCMNVuUFZHkIVSPSaNQkXg2TSP+MsW92X1AN
H7NoEy95owg79QcmU7TYeOKEIhFtCDumJbeWQIGexgWfk2iDfuQbfuIpdPIFwsK9aoPsPIYb/y+y
7j73H3OZKvdWipwfkMiDqzKgL8cFNuYdfYjVmSAoJA/KGRJseSGuiRhMQ69V9r83zw5fuqL7m3RQ
BA0ign1CgEBfTq4TEjHpDlhhfvDgpkWrQlP4HK5UItgp1xqAeql/wQIc4qnUK0O5kY5F7UNZz2mA
sjskq3C6UD82xFJ//QkYH8PZb8FBDCr+ZbNxEp7VGBt2P7gflewy/7cjVGpUDzKAwFUIbe76xlLT
FRwgboucrRKaqm24IWa60dWgHRgkxr5V/ht9LPUMhy85wOb59ElL1j9I2Ki2ssR6oCjg6xaPk01X
Bou37fxXWmGKOpQobpZfCKfo4rZHzXsrbTOCIEHPWIghWBnq+Ymep1w76ZVsci5OT79QxGb9S3Dm
k26ThqwuQ4elizOeCdfU/lVD3Kat6sV/7+Z8LsCEr46ShWcu1LemebSi0JpmAfyfzQAHA8w7Sxfa
tVPmozcxqNuNFGjWyfEGdx+Rtq4X1MMOE6/0NhgFqeQQlN5KStZBw3eT7Y4RUR7gG/+Oum9YMrMB
rC2nglPjGZcExIdUiGOuaNN4/skf3xFEk5kMHnP3Lu8DHWOF2pyXUQY87Osgz3T9GGvVVc4j6Q/T
E6j+Cyfdiyy5QLh/4Oeotmx0DtUZtoFrXxgQU8B3+M5eSI//kC7uJBUeW55w/O7Yi74H1tzrt0g4
AQsALdRPr9Kog/cJ4yJk3MVj59n7Fi+aaz104Z5o2FnS1J8LKDm+FF3wqZzCxfQOG/RmglSLiR7P
L21eWCVzL1J2HHVHOsNCnZuAoC6gq4SXYJ8O62SAvRI9ANnsYk6TItPn/Ky/q8uzSplIrE6LXhfG
zUZLZE6uQIyN8PnJZKRlfhgNmXqOoteD2+vovyg6GXXHYrm4Tf0B48YXiUnMIsAyB5XMUqerATBr
N4m97WqiiDoYrONRUhrnRsZfeyw+VuXza39EZHbFoGgfacPpaTwU3vbuqFBFibvVHt+K81TcF9Hl
vBXO6nv137U/qQEzfUxO5xrRTwNogifKIpLegx7SUJLBo6S0hFSvIjrh1MepFap0usTt5Bk8s9fM
Y4lsY6jiqS6xwxac22yJI19JWMItLKNqWS2wvfM/p65flqL3K9GczAuv3dPQh0nuTapFNaugniRS
dZMhUpXr0YGbvMPFDqAn0nYpl4rlo0IITZkMJGkdDArui+6VK/L29Jp0NAIbkHWvy/Ax77ypCpsZ
ZEgyVNTOJ/LVaNFwCAdbi+Ifah4YAe/QzHCSfUsFOFY9/VLrkT7IBnpFgME8UZkN5XeNMTNUSVBy
XbgnMownPpoQYex+vFMtlQLk2IJoazzi5AxL1p71n9rQsO46Q1S/94jsG3hz7MTnqT2EOsE380U5
xwNPFjiV/GGjBQNblAuaqSaGmmN4jIvHtBDwaxiZK/XRRZp2jlBewGIw2U9uWV4tqHrZDjLHr7rM
NqXGfBGCxG87Vb3G/wsUJdYOO9/DHpfx3vYzANfsV2YNgb8AcfbFoEp2bym4t65gja8MJkBem70v
+DEv1L7B90LLbnQ1FhpJGjNCwBkwUzcU8xUjrkqM4O9bqd5Nfioq1ZvD3v+oio73iHqwSYhX1d5j
rgaOMwM/8JXwV2Jbxqg/miL8h5CSU03nUiGX2s2iPvaekjOpF7w5yp7GV//sDZb8nERQNUwCm5Db
SHQqqwGFOOwrIwxNHtLUAAkRKgjqW2zg2Qw859/M7MSgZ/8vA2QXPuFhNJnKqH2+4G0v6mcUCuBX
4DTtILZC1iOD//tChWN6e7RLo0/kJ/7Kmb6n6B6g4c3k4q+zsUtHeqUGsoAeZ/Yvb4Cf2Qho2kKq
2NZ0bzemJepiRaJ7ItW0TZyRj+igKSm0pXQOV5SwQ/XRMxOffkHdzmcgwsbUEnEvIWPAoKXoN5/Z
3kaibEKsbGEWAm99dGP8BLphYpIjwl+dov9dGHHx2WeRbhEjfPNBNZdEKgid583TDfsffi3Pa84v
HFG4CtBpXsiFa8F7TtYVNQrhfLnX4DutZIucfh5NdmBvUDKPuLoOMUcaPzLgTAganboqbkiGuCI1
hUsWfZXNUQ21pw+ObfMR+4rLKLnq2m/Afz5deZpN95KntXs4Rqpe+iafmxe7lRdj3RPI5JrYzEb8
U4WpLp2/2AC/w7/USHbkjCwl69SKVZQ67dtwW6waTP7lOIDa5BImqhwPXLQvZNTRf9i2LLzE6gba
RKugU9iO2Mcn+mc/CX8HvmQufAvXBC544izmk5A1jdx/X72Co/ZGwzhbGlkjlIxjYJxfSVIEZlKw
3uVXo/rfcBOxuUJERgiElwOizIwcmeCIovXlVLiQsyJuDFbrR/Ho49F8y0nvTZvVM2mDmSIrzH5A
Me+9oA3JOVRPhQGgKrZDyDWx6entf8nQNkXGUIBo2uDdOK7JJf7sCXWRu7TI32Glj5zUGyt8UX9N
ewYBksmRtinWUW8FdA/9S3LS7xiNlAgO47BFJfX0e0QeOp5O8U65WzdTQf8qBXm1EOp0sLNiaOXe
5ajnvzOjr5PXbfEHCjr420lxzWcCyloWWARZW4XdvRZjkWKuTwC5mVYLhPOXYyfCVIc1dSA2cmip
k9MoQ624c6SGMhazL5baPkm0bRqIGklCObFybslAiMQicyp9dG9R7jmrfkcLcObywEyQcaZUzf/k
BqfCFadvpGOAGFhx7XKkp2Qc6tQGl1o6eDUsb9Q1M3ipwmR79GWvs4YoDYvtXmzjnGpZC9pXmHVi
iJ/eaHBU2n6548JbRyPJ6M4GXqSCINEAgnT5GpKR+TTcqvld1bFF2LAp3eUH9tVBTMk31cmV/wT8
Mq7aQ8Z6tKceGW2zcfvSfmFv3i5VDoRMG+ydmAm7LMiYHvAc8Dbg2qfas2g7/f2xKEWKuTnmK08+
+E2IbCXZNebgcKTMFpKYpdqmq84XA5GPLy5aXwBePVG0EHqPAW+VMGFoZwnDLfWMb3Paq7yy4ccr
/l/2iDGuAB/iAV/0386g5/S7+TR14kdg/iXnIJ4VNwKVQ3SmWefOBut3MHe+u2B0J24xege4/mCV
OnRY0w2h6EwciusfSKJW2XNCB0WtqBgucyMxHGxx8ivh5p6eaUKK5KtIKCMX0M0wpolLXNFA/yd7
T/rWmAlINUCVuwDXC7k+QYFUK2UL99G2Y744bgla/rqJQLNAS0liGr+8It8+uxi+pK257h/o+oLK
tifpPfwSQUFeUG+rSR4fTFrOt9Y7kC8yz4AfafZOQ7U37oNxN7fwvs2fvjLfXUJYqUAKERm/QuLg
YB5wd+LCTJ9IFIRLS5ltDHALn8YSf5ZQapWs3fJccUUGxCiIsWSja+owHPwchWL5nGiyFQERYwkP
EVgUP213mPU3bfcz1Tvl0AUjPz2tRA3eSvbYNXp+M3FTN567ut4lr6rqQisqKfLxiFKK1USA0SJ9
6cdw6VFi0TpFgzbJ0OOxaVDPBkYf+yhFPZ4seZwOfDES4910BCPJJKhe9kQOIdJ3drmPM35OrL8z
zc4qM5ljXtZkX9Gxt7j8yWNML9f2hktGZmx25LjTdeEUWYfpPrOAlqiinIDOZETlWRZVEdZYJp68
g1l2kiPT8/XQAdT97jKiBzVBxEXZbvtany5XQLyL0CBNEAJsbEZXPQPcVYPbx+efwYf8GSQ+1BeO
LbDNt33nB+gU/pby0pbMh5TLUU+zW/dfTS6brCWsfjW1jrYa8vpnp750Ciyk0iYy860ALTFXZF4m
HWH+HhdolwqX0E15cz48r0hMISkWZUgYTuS0JV8wFGKSMo856GXZYuhFMVp919RxLjAxkk9Qzh2l
k/RB6+mlkH4/E2T+ru98sWQPu99MLxc9IQmLIli7UW7ZxaCNPVy+kDKL5oJdDrR3ZLsdvUMlpDy3
HmSPkJ55+AzQdc3AcrAs8oo2fdvc+Wg5wkfNFx9pjBnedLwoPva8kaa+v81m8ASSpb12FkeQW31h
ReTRWAEokPQb/T90wS2CspkwCUiCaNiTxziZbnl8NE/pIthmxc6k0Vxp4RpBhz5jRTKFKSqiEX2S
tcoOleBIv1hgC1RRfiNPCvwocgr1C9xYd/4i+QSTIAecQQ/hF3uEmYaxAuX6g/nSs7T1DZdQaEqX
LG8n4TOBgYYjWJld0VxG4iyxsCblsmok9Hiv5407NL4EUswruZVJ9Ajt4ZEc4ywMf10iT+7TmAt3
0Nfy4M8hYBvXMwO+mDwIwVeez1/wNB2eogriLkF+T1w4HiQnJQNA0va2SANZJE8cHQYaU8ZY+HUh
RViWLFKmub/6qR2744mZ5xcETWQoM8q9GO72uaTq32PNdu1BNuT4J/brjNmDiN9gZSB2eoD+aqDP
gWBh9YaTzHCm3Q0V5gHXZkkVJjOz9mkxapHkgOAc+zDCbfIgz8xE6W/f4UNweDU6cEMSTjbgqp1D
6nUOLhaj4AQGwnUmhZf3aQAHidwGx4qaXh8g/Nd1QeJuNUKPdcsIOsfl4SaMkxoNmxEe0WQqzRc7
a6t52QGsWkESCpi8jEAPgWsmMb5WFe3bxbQ0m0x9k1P4C2KnBnhMR1xj7DlOxfGQZ+jxm9k3lFhU
1BAofY92IVBeM8CCfj63Hr5ohr4AttVshwtDbjo1xDtj56AgCs6sJTwULaCSrAs2ExDroqbiuZxR
MO7vzncih3c/JWCNYnf+G2Emd2JFJ3skeEjk6l36o3qJm9uYtf4ACwoZ8hVpG3wwv7huYIRJ3Idm
QchM4bBIoe9FjNjbzpx7pufBVwGPueLEag1a4Z2eAl+dW5nG1Bta2Cp8207C/RRHQVX/81QT8PAH
OZWZnrFFk0jpNrc1bRAiSnuu+m3BtXyloT1NfKN5d0T3J563DSi2azPuE5H/VaHwSK7Slq4mN68Q
LULb+li1zROV0wlDFZ2n1TdgFn/0s9+aFWbs3TM+tEMbAFqYn6CwDrNrqEvTQa+bFNKjqenRTGQd
um09Ar/vpHUgMvY2/wtVleY+H0ougvA9Ea58CwHYXP5gbIzfTJyT5cgv0f+e5txoj1abGw5/V9sF
RRY/Dkg4Bik17YG31oFEcKAguwre6M+NSUvRwU55uApV04W1NDt+toqc2QXWjj04EZ076NbtKI73
0qfZ9yyUm8wxuMqlselCS0XhMJxZhG8euGvbeIC4IyRbzaRBSdL+WCsgYbb6MLdssHtFvoGWoBhV
aU+uC1K6uQ05qYz+01gTfL1g2a7lebHWXf/qn5UXaeuWx3+hjbM7b5LLGSp1SInq6mbfa4K1oyeX
418j2U947yrIENUVrSq2ftPq8//qCEgv6H36hVOjEccLJhz+9Y5LEmLBhNKQFDL0xceRBEHCU7Fk
5Zmcogxie3jsjzoukOb+xgJYQl8FHChRUItE+OUfWTNBtzk4JLswE0A42l2xCwaGdqD6tAzuGwXC
cKlfxX2uksjlH4ThreNgqJvASooRfZZURa92o9hpVzJxThDvjLW0coy1h32zlJ5J5dqeMvocHzRb
rCcYB4f6XB9+NSQho9i66xRjYPuCfhjBDklh+xoQ2sypZGVMh4lURt4Vm2yCUyYSA+pKXI0+P6ou
h+VA5ZQwTcqxv7zbTYwPBNKlmVGxqFRr2erQY2xZEhYA3zZe1wKBE42gcgIx72FtCSUInXzpYnC6
a3HuN9tq45EZqoBHg5+4N2baDsVrQFuro4HgyEvVZan/kUj/GarqVJvV8ud265O2wYbpIdUVExcs
d/HRcA62l6BJZCdkCTWmQxJNlWivKeXunaYIb4fs5bFQZOMSvVy+6urUTEUwnlHWHY+zkG0zCU+Z
8AV2G7YCccad9E+s8Ok9KYrd+hass2ArRZhgD9Q/rSqnCXSJ3+I2Y8O/nDxbxS7fn91SVNat9L8o
7kMNSIxdrp0BLX6OWqTvZomIzKOpDPgqdFbHqeHj4Eir2JkGjKQdUfd+E97FOq9M/O0qiARisvUv
7nt1pS9d7+yIJmKQcHQYbW91qQlrRwvXPlNQtHTXlerQ4F0iy/Wt1KK2Ozz0VckblFt+LDEUWsA/
P4PkhYW7xFuExWn6CvtgL7DU/iIX/84Dqkf2SCNuIbBfwNCZ9hbS2sXK/aRc9Ct7oGMUzlMM2+PO
QeahnC+/Ae2Rp6AeTTq0f52whEx6dQXKl5vI8+t2Z+tD4dBOgm74oBoDArvBUQkhP2GA+cjGezi/
FUAQznubSI7eUDqosp550Vhn4CS1EagApYrCMoaIB++EIpyXGQsmwn32Guz3NKcmROYxTsMx5zkK
PJj62A4aL0sbkQtfGgfqTM6bESiWXOHflbpfToWgqh/rBvu4oXuxG56Pdwjkm1eno4RhcHT9Wq8e
pcT5dF41nFR2j5jfbChyvJShqSFaKUElKvcddI1hermV24msK3MyURv4Z6xo0KY2KQVRqV4x6u7D
CQe/cC7dofL1hSlGXK40/T1PBwBexhJHOmo/7UBJ7fJlV/X2ula3o1TuNQj2vlIEqhqmajm+0+hn
dQTUUbKL7lo6GDo7xQ+IQJ/DEgD8HO/U0cXYVWfig4NHyHbwp32NXVDSv7eeVkAEGNpSKzxnjD9A
EZIOaSV/pmDk5yNjf4WNsfRGJFoasq7v5LY6AjLKviVVCcqL+HgtA/n/3YoAXDObZ5vTL3OR3ZJL
YxePq+ffGZl1UY5ljyuE23+669oVJZOinkS+kjB+6vNkdz1658Vvln859nh9f+m+ErF9bDidA8f9
t3YOSTus76J5wUgoK4EADzJ/FanwIiVa50YuVyROM/ijv5ux2cnN1BGHbW2mgtTQ5LDdNrZ7yRlj
OutIZngNHqmq0V6/5OUQcxLgTkN8+exHv6GSwDhYWN0SR0MXyyw4WoSQiWB4L1FWIAD1fHxaTweN
Z5d28Q29TFxn4K8r7vdKdG8QnXSnixLBqxvEngPk29zS9cH4LDWXrFT8+g7taUt4LkwFYv8hD3Kc
FRPQFCLJWZme1gN3NtE2IgTbjinG/nXzfK2HKkvcD+ce608KDkuczC3VAQVHXeNFiPGz+VGJFCz4
Jb8xaMGj4u3DhIMw7FVK51uYyrU93XZDf7/4IHm5v/KYUnY+g+47Zw6/WglfaXQLPMRzY4AkTsG9
2+LpXnU/ZdMGPmSkYMlM4uPxxjRrWN1cNJhgmts/4elfYkRFXtIbysRrFk2VEJyNXIKDo8FW4eCv
duY9fCdhflbft+P8RE+M6ZuXxtwdAYLAsCNF65ey6L1S8MxhGnHWEPy+oKsBons+iU6kGUlZSMJN
GQ89W8rBkIBwl9jpFlwmWf3gNofVdrrz8X3g4OEVxXUbGQ5Z3odMmB3B8pECifu2aWdGrSxrMWH7
ikapYbYWPLALxAgCPvSK9w+jdYpzegX118MebnWuWz7ieLp14F7zJ18+VYh55F/n7cr1aRPgFS7y
suKHMl07ZNtV36xMC/TyELVyypL6ef1Xj/dmG/QfsPnX9r/WJscrZECwX9YDXiAvJzVaVJk41GSJ
f6Qg0qshgT6t5xaJ1am8udfo23f2WUFf+ukaFYLm7zfqEV5ZhpQMExeJROfy1u3m0mISgmRgPW2S
BQVek7ggUnnO0mE5rob+GlFO5a1bOqjZgGCTzGEk9QpHMXJvyRHivfjCE8rnlSD7MH4ceQhx4Rzb
y6QpX8rt8CunXV/PsBqduorTbYpQPjvzYQQ0h37H1Jjvyro/78JKsO7Ocw8li/iTFSycMLi5w6RV
axVTLBy7B9DTjn8UasikL0cmVSB9Dss66dg5k+0XBozuRNc2jSw0GG2Gy3P0dEwXrNEjfBYoFr6D
lGzTygTEJC1OV4UfK9mGpLyQPAobiLeFbVKPtaCP3BcgcyhZN4+RWljRTirx5O8E27t3u1RcPxEt
zvp3qncuBkoIAdvqkdu84iUagAJAL9+aYJLUO0PkGFP5pJ4FwV2wuvuM6QrUKOUDD/0ZW6LSVBYm
E+X284OTL9408erTqrQAWNtCw7rAhtApMgfzNVEDcnmkYmcU5f/oWhJMG9FeWCVOe/eTLykESMuU
okH+fDZQbYepNAs0W0IjUW8eGD36XpYTp3GzVv0OC4fIoyPsdY8eaR+2waHb1EopZQgalJYXOzzM
41opdjjzKM5aeMW+hatR6M+Ej5ZawDrAYK5BMILkS8DtEEUh+Wbubyns0hO9ZM1KsUKRWCHlkm1l
XMt0aPBj2hiXDdFnWKp5eLx3uHFHn+v+mjyLm2EMFblr39uWBnl+IkFmVFO69hMCMjqk/ytYAkPn
QVv9Wm61/JDaiEdtP+pEFeDSdepOFncM4K3Uk08nxxukIeIlGJ9yjwaVxjGA43D+x2wRP6wighkC
QWjyZiawDsTl1/5bXgdHG1FbGPioTrchE6MnJEE9SYZ7rsZiiYxPd7lwNYrdQCTuXilrjRRZL4/w
vnBpXaRf+7Iz5PvKF773BLKyQkmhCOWwZL/82PYiH7W6x/tG1rznoHSu4/mUI+x5vcqYg1hyrAQ6
1H5qOWX7chQ85bQ3k3/5WWyw2Ke5CWIAnOhLfTArMzjsNU9/Xjn3+eoWToLYq2KizIWp1ZXXSQbK
FcQ/TYQMfOVPaCSbZd5//TguYi3J0RGnwMr2rfiNZQp5v+SNsE/dRFf5f36zuh30Wt6ZAtQWTkf/
RK3e5vUSOyXNoYTsQ36Yk0zdL02Tcu+4fKlKmev1jhmZg73OeSYILjKWAMpvmSrciVOPPiL2fC91
6oQFDul5gbCtvn2/k5TbhAS4YJjbcTllM7uDnKMCP4H3LEdAFu5z/KX+AS7JCm3gAd2PPqroQXbk
gdWEg0FIy3+pcDbPPPbN5Zkx3wUHuvCEfkIS+VrliTEEpJp10MmUz+5zn1Y2ulCn4a3Nk9GixOGP
/i3DDGvq6VhGUzefcYlxvJJ3Tgd4Z4Zn4k/Ol36rercHna0gbanLbBiqg+F6YBNd3whmL0xYkQZM
s78XGCRgV+kYKL+TMtCj3FGliKVoAgrgPPbtGNPsZ7NGOvH+599YdslYvZ5zuHg9Iv/CB0XkPRkJ
bE1dD++gfPrFS/zJgzFV6dgHKQfXbG3fs95lOtj6oVOrhkJ1k2Z+H4LsqeC8iJjuE8IbvUn0Svwu
fDJx0jF3gqcmYb5/+ET8v7h+VOkwsMp2zggs5plL74ZdXcfj+L4aYiym2YD7bQznHyCKG+iM2je4
TN2C7ZHWQLtpXXelY2HDG6oiSzJiY0YksvOBoQ5DLrJyVtA/IPI4NKkCPm1oSzD9N/1MFXMRIBg9
CEc97XoTqbxHDr1so+cbpjx0qYOpfUi2jd0RCTng4QUlIkTnA18ouW7BDS9f6YihkW7GBjs1kjCj
Dj/PEZpsI6p5XUMNARAiJunjVhOuHx0JSMg6ko8ZIKYhsIVgp0HAU2cbHgtn1HG4fI19TMKZ5Y90
MdtmXnvnhI/TfiCGiUJ1jXcw1EsHHG7Iinart4+eOx7STJjWPcv3/j/McZrRg2TCCxQ0rSzTzoct
zQNOtG3p3UKRPMzWX/YGzo6h7tywfYHAbsLnuAdDOB/wE14cGndHw9SSbNlIz3EdmWUpCxRwL+PQ
jSxIEp7ZKpYZ5BZH4ydRbFYkJ8BuYvpBPvzeBoUQInQ9hh/msm0p0xrz8xmXiIxzJl/mIbPYePKs
bVB9jlyQX8cZU9FduDSpCorJisSVIuBx98q5LLxsWeXNRMieExeioJMeW0FnIqXATFLcR7pP8FNS
buAnM74UH9+1hELtwZ01abgQGfUewjmTJXhe7Jc9ISZbIq6IU/uUIPMhnjWX96wdNKkXxeX/sQ+S
044qCldNKZtEK8hE8T111Dx9RpG3bGCPxKEhVADdf2skzJSiMDA3O7DRFTi3i9Gevf9TrDaRfCKi
f+dEGr2fkGD99brvNNmt3xCrtZ5sCHtNzyt+o+WAtI1nlZGRKs/juAG3q4Dr7u5HvWOuzNBVK7my
fg7+hGCFJsfR4n6ZGtG/m5LeAxf8Xz1ZzMRZHQ2R0DqB2PeLd3T46VensvVr+Ex1lchDhFTrq4Fp
rZPs8eo+n978SRGTmL6OcmQncqX/gmvwZv8I/9KhMSi0emn/p/qnhA/GAG/hZgfFhZRIbFM6RfZ2
kPXdMqxcNPbSbzLh/RROClxcwznRKh16a1Orj2f4AlS9amHOBaJWyv1QRQkMmDFAlhvtYwfj38OH
ezuLO4UOljjnsIYN0jAOYt9QPtAty95yvMuM9wlBiQ==
`protect end_protected

