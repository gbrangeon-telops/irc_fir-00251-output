

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
FZWxslbw+U6Wgup1K8ZmbZ8ZvAwEdSXoQX5Zxu+YDpvGpSAvyJJdij56SPMVKmhf+X7kxMgvbsEm
5B5AiAyVHQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ntA4Op0vLLt6gLQbdMxO+e0Bhjub4O0zQAgtU7SVthNE2o/5St+SvTkDoJ1ve5MFs/Rgt4JL1gtd
IBaLjbwdyEGV2JKFzmLfNOLgk4U4bgeRTGAx1e+I5wKQlcq6qarG8xv4yuzAX6jRFWecgDUKdkZr
uIZCcXBmuErGbIdhFKI=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
I/9QBkeb84dQg6xWUGWLN64S2R+IIBcNXAJuDMwqYLTsejjUFtntzi/OgGH9xu74CzmvMnJuiSkZ
p7NF+AufXfE0LUxVeYNmvB8UnCKeswDMIWMuVEpX3XPk8OVFRqBWCRJ5c38XRjldLuPPEii8dq/d
MjasuPQowI9n5pgL7s7SczhrYfNu0A0XEQTAwaUPGij8aO4+LpdeoyqZwdg7p9EXJlysFsw3bvdq
qHiouBqf7MqPbKppmCVMlrH1R0q5YlTlllFEZblTUq4IO2ZWi+5zgGnEERNaNBZQ/na3tnrwOTGu
mqAR/EaIPbn2R/AR26ZYNuBuu0Ym5XtWJuqzJg==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
jRGmdT13qAzfiT1K2NPIFkj82nI6QO0hHDoQ7U+cF5NSt11k+3KuVBnDKOWta7RjBJSeiJs3q5WV
MSQx2R9/yJGRUjq6DQS8PVF7sqUyuFjNc8w4wdPwxcG0hsCFj/tEGyFHTU90BhMVIeVjf2WlERXd
+UzGn82C1ATZxC/M3Bo=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
c66DzsXEGPMNOrzYyBeymw4AV+RpL9x7eTO9Hf3l3y/JxC1wwEbipw1XtleybcrcOfKY/ACDBUVi
s9qFxHBAPyb46Eh9l7EGLGzxXJTWMed4eJI910mZ+WMPkBgIF1jvUqr1JGStUHDdUjBjqP5Bbe3m
2g3HBNLeS+8Ciq924vg/jBwWCA+G1zUvjlqI48sc1XMFszL+AzQf3r5t6tBvdkd9goSPiuISrM7C
eaSWriX/kCtr9jogh2EYVx1Ud4JT59uRVRlS338jlkF39xoR0AXtgdhjpZa3Qu6PtAnEwyq9aWWk
FBo+MHknw9HNH3v+t/wWSpyyW9f8/AhQrF1o5g==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 12512)
`protect data_block
DB88D7EnVct18vg3yK9AbpMqZhc2O+/NA3RsLOx57bY/t407ISqsieyBbsIsPPIgY3sa3aR+/SK1
fgDdwz3oD5k1ZncyvHUTK99KAcqT5ll+R5SIX5x52InECRwuVl9CpIbXAWxH7jSuyIHltCYfBTup
r76JWZ8oCEt6Wiv3DByPkcsX2XwxzIp4uc28PwvxYHMkzXqUpe2miWhNzbVpd0+hzDcNsuxpqIBq
90C/QzQuHLKcEuZmFo86gV6+o22ywZX34MpoKi67g2qKwYy85/WvJSlUJSkIrg9Y0Qky1beUn/n1
HiOFzYcrxgibhOtEcCey0iZJ2xPDXonjaanZR75ky6rbKfk5wtM4hHgZNfUesYBNsxVNKvru15Jo
9m2pMHGl6g9CnQgAnVD4qMApWp8yV0Z6Vpm8tsJp4xnnj8D2VK9/wRYrOnCzosS0cuBEfDA3qa05
Y3dFrKzkdu8wt4egL2Aq5yb7reNJnjjyfkd/SEIVbBl87bnwgo+A0066ATDBlSvdX4Kp6cF5nDG9
+mmlDtTvehM+LZL6HSVKa4TYmP09bFDLoZGfBuHEnyMha9uukWe2KwquT8AwHw23c94OQoI154pG
dNEA0EG8XKiRAOjwUjaQheYTCi2qBT7f1v6xdm/0Cam3Am66xobw5xpyMMnvwymKhKR7M7SVMK67
Hl9QzcsQDP4mQPBVZgOqKnUAKefOJVs7XBFuoKE6+zPwbBl+8680dOg0Qk6l9OBAqSkHqdUk5lDY
DMisAXp8udkBT4yuin4ck18eln98obzS0WgfP2R470PvuGUJvIdK8hf2lqHAUcwVW759D1izd+tQ
2kIWheBMTC/tX1++15UTcJSH6aYDDNA4UsxPQn63oR2WjwJaXIAklryb+9tUajFTZS55a/juvFWb
NHYv1ubGIBfQOTDDtGXCPZJOHj1vENIsUKR+nUufC+rK1AY5zMfDYsvtDZAqYu3hFH/dgUS3ckLh
lDaQX72Q0Qe7aMctoykEFdu/tApHOhZnFZyX9OttA2yk85CLvB5TVj8Z6PW2hBGzS4cbijQ5mKx9
nc1k0IIwWcy0B6xaBN25i8h9m+Ee0KnhxBoCOLsErtfVYkw9+9ssm2oRDDJzkTc2+/KPlSTfqeUw
HwXRM07uHcgGm10+i4qN+m9bKvOmOAbUvL2e/pi+BISStg+R3+WC3ra74c7+q+8w7k4Z3CAUzCTU
F1DIROIkCEv+U+6+fZlw0ls8mUPNN/qhJhD1tSz63CPvVuQ1JpqFyZNGN9TJhdqt/KHkoGAILshS
BqDfOajZT2gOKMz/zdUuedXjIoaqe+emJCn0VLOz4VTZRaBgmXy3ItjCCeEnDsw5bObAzuaMW3kf
DCizfs++mYMVyO2HOtHQ76zk/nrhRZAqL6JGb10OTpYOB1+1RK7YLBbhoC652XzgmBMi3DAeVqWD
ibQ/WkGNVkjC9gBxlNcb9MPtYcT0z4Jt020W9E6Eu9KieLb8tcfGienFDv9FwVSxtMgKAQ7pxdrd
QOhkniiHH/VeroXMe4eDuENaGpx8BNlgykvS8/FIhMj7FmtjpLTryd9dFQQWxrhPyU20DcIWLaUU
WeH+TNX7g671qxWBw5TOG4xFFGrJFVYibBxsZeB5Lk2xU71SjKEISjLYyAEJapZp+vnYrOW22efx
EYtqTPXXrAPQ6QiZTNKm7J8KalciDAGnuKjTXTOFI7QsP4hJ756E9klSE6lyXls1gQ0lysNxf4TB
ng7T8c0uIVAVq9Ep55iHNzYZc14vtjewBbm2CgadyB99ObKL1voLgAg1sbNph2cYlOCzkatRiuVx
l4pQ+EPGffbmz1lY9u05kH9sGheKhlNMHAuT6tjYKoi1RaSLb4UHb39UWpZEQX3pBJQQdDCATF9Q
NgT4On2weSFOaGXrd4ts3VjRfFRC7K9ELAh7PuPYymJX8sK3UtwFYm+mUd+pJFsCM/NG+CWlppC2
pXasn94JDIX8IHBDETFlr65HLz+Gir+TYSGrM4jig+ws/2czBA54RDyoOlFX73F6eD205ZRnkeRx
q0UJVWDMr8WQ1cTa1oOkTN7bqM4e5xNEIO0DcpERbOHyKcfjXbCyelJ6kHnX3F0Mr/luqH2Y/w9v
0f3ElJEBUPJ3Awwc00rbL0+8wtHRGgGyd512U3yX/Wka6AaoBMhEDmBp4Odo02/yrjWmK8OtmGqA
vW+cYgqjeBbqdXezZsV9suttadMDsjLdqFt7DIQ0oJDFqhp0GeabPzNLAyVGmz/Hoeb1vhJHb/s7
brAPxrUHZYjDjmMXD3WxYj7xv8UfvxfV5iJGs+p9zSi2aIb5Mg64hdgyR7xT8930izfbF2Dn3J90
tFd0JOW0VZNXuUtPmP0FRY1ZKmQrtdQUkQjRZreBH4JvF4JR/XzQq+Ry0htJGslilyHbuQeQnB3T
DfhqM7QgF9umNVKIsPDT1yPpmEhUzuP+h8AESdV9eASrGETqqWpNJqYeNQqd2K7qkDlPfV2fGQb3
Tc1zI31jTSJYUmDhstGHo/a2/LAwSNgZqzn9flqJovsxjpLQLPWrhTkLfHHaCzKFl96qAEr8kqSg
DvN8uLn67IISjLxdbCdngpIMR+I+f2i0LC9AYN2P1MIrNwXt6FLF+D9VC4liBnHeoi4vo4M6hHSG
uXSJu6+34fhmqvY/7fu3AMcbDJme4GwPb+FiihNsjj5pgMjk3U0dBNlFDAAmsCqJlAJu9JWwcaNy
MA62KzzXDnSbaekPk0dLIXvZVcgYhEgGB8AfM2eD1quAFmWTiY+tVzsTL1ITQuIx+1eJwxol1ZX6
71Q553aCrTMe0P93WySJh948eVS10Wb2BTsdY2EKYxQDiRvhhAvu6aXUGT2735fMZfveTYNkARG/
h3gB4Nv/9pCqnTIpkuA+tv1zQ6xdf9UkkoU77e69ddLW+tpcOz61yH5qwNeTE8lz7yFbuXpekEs3
ftxOl+LUZyrtAQBHpmB3XUkL3O4CC5HDHXEKlAcCY7AfUmr1F+mW4m8Rybs3MUt/VCCf3nLNBJKb
UPSYA+pgGp98KTR4TM8TZr5JU1pDr6r30SQ/MHVO/caJcjjBked38siAbt4ErbFwYtj44IAfkFFh
DGhxKYmvlu+q8vFO6kG6fQu5tzR6Xzx+pcUZVSrpezlQcUjG352EjkvWJPfVk4BhKy96zi9+jDx9
FG8rvK2T9SLMNGlvfgZgK9RMPtmksylHV5BoqF6xJhcF+Bu7fKYTIIOJrsAV+fuBaiLRW3gEHIJn
G4utmTl2WYaUGa26IpH+lJdhOvf0dEWI0MU2kXtMLYnN+LzZ2qLIGluNw5OoBSQc80hqcr+K7J5u
DBHxxOEm0ifjaklAHuSeEVPe7M9xI8KvQSaRff8EyVhkeCGkw5b9D2ICWl5oe1dnXmCgFCUwwbs4
oRovrbx0+vrn+ubHcrfOWezKyzXjVyBSKrtHcG+WagGlERhN61IWYAUK1ZFyybkaRnnWpVDFBMNe
APWrdP7SZa3l16J/KBN/f2uVxUey0NaA0iBj8PbkRVWMepJ/1w6o8ozdOE1b7RK+PEy6fOus3TRX
0upWCSXnTmwTCSarrTrp0gmX+sxNJ6LtzAI3MSDSxdYfJevO0ANAQmoFMHqDDSqUid+Y5kdMFVJj
KXCOURgeq39jybXSrxFfCyqMWtHBLBhDaQTAH7R5u8uiE7B+18HA2aCJ1CL2oXxiMf5d+ZDw0ppZ
gwZYcXhlvQjB9IjSkVH+St4zsCPTZmR/ZcFDbfnLsPyzSFSdtNDIoTjL2N1mr6LMsB2F62QL9zIJ
XzLdIhgX4k2cNWDB9X/6xVDteaxj0e8oL+Ntf/4cAzD014I/dILwDrWXF1lh1Qm+NehrkICbvK9R
BaYyVSvXnLLgqbsyhWSzyYbPmfHOcCa2UfuS65cHkZLslD0DPMlfrOFETQTnctogtXKisozAaT/g
kLtAWiCbTGz3ru64+5/h9/htTrRnfsePL0JC5RflS2J7DUWJenmPXgqQm00VEq6Ua7uRBbjTh/cN
NCDbYRAtRBzL7X82OXhNLioUpFShAmmw08bCDCORZg/RhVXxJWyUzY9P0OXEUTEsCnVdqrGQFpGH
EAHW/CAujnTr5Zl6s2zEJWS1/WJeFvJfimBGgC9g0liW7ZRmXf4VVbovr0CslzqVRqcS4itD3ltm
D0lE19djubRbjDaXnCufnu/vkoi4+V93mZFgOgRBFymZDlAk5LtrRBKpcZ3lEnRpVB0LAq2FR2A0
WsKZZu4jSVQuEJiMZ4IhT3MwbV7u0UqEFHcYivuaqei0dYbx7vBssvQybxg4s5J50ovmyiMi889F
c8KQoQjRPr4J+3fmOwtMTaj7101evOu3LEPwIuu5rwO3N6JeGlwPuHF/A5+GbHbvPGZ+3Lula/sd
ReL4w2i9/WJrnzSsLh+1YF/LBgrCz9eIne+qrPq9XL4XcHecXSkLzAYTfeFagEzQvwq+XJIIFw66
MDGXapUh3Cm/eIKdaQHR+7UBaiL1yKq2Td1n7zhMYlC4B+m5dmHrvyx8oCezxssUAaog8BNaDGoP
qRsxEhk8wXpvHPSSzkOxg3WLlq7N6xxKI3nxyOvohGW2v2fqfVwmtk1LlRQ1aZ/+4WeTXhPkxQsH
W7FnxordGv0dPDPiRmC+6kBtOLtK99ChT1obYw66JBH6XieSR5kG4TMq98cqNIrhpQHy3kzYVPMQ
QuW1xxqn8V0bAOALJQV7LkuE8RgeqqL6bb1CYFjaTKubcNyBQJIfQZraiFHndstG0+l8MioNYW3c
86JLpSdEOJDBFLNqMGvwi460yteWuYsPRZ8gx1OQL0+PmmI8e9uO/REymGnCnxh25zCYc5jHhQJc
RmjlTO2vxUL4Q9Rv5CR86QmLsohKL9XtKXB3Do0BErvr5m9ferccNOrybOnNILmz6JQAJTpXfW2c
l81jgUNR0tFznnNcOTVttmIiJlLGJEcfhowtxJLXiq0j0nuLgTosB6Iwetv61hzeifeluraZSKKS
/9VjFRdl04WNDS2vpM+D//MFkkrRORKudRe3KSeQg1TEay5dHvOj6YULH0W4yw++E05RObT4rlBx
qzlYYmgaFKKrjaNBxVS9Lx10rpg+3xhrifleB9zlt8gU4873Truoz04tndYBENmKwxDYpzumVFYs
HDoVsYCWdkaxj4x4stNvQqX2P23F/eWI266YFcZ1IA8GVFUxJ00DvEZ98FQ+KFBBOjTs5T6bE2YX
IZLc4KJ77+ZMDWtugHAlbrIxw7oNEPzndxMgBhbsEIq7yuWSdUa5U1qf5OpVboQQmtsrztTRir6e
z/y4BuivmDVHL0OjfZVXAT7Gehxr/UuO1xsF4x2GF6SdPTvMjdQshADRnvZCGBhGb1lAstIEWeWo
lw+mo2lzE++E3hlslK9wreAsl1DosVriVV5mZbFM1GYBBLtQsJ+eMM8o+JpLG/4sgTXYbHtcLC08
St9CfvNmKGusc+KXolIb2+FrRRoNegRLeorv20AwjIdC6rbTbcbjRddNZ5cItC/GZVJil+2VEe6B
cb16WU9D0BjBb0jWUhydpIrxTySD4A87JR+8OHutSWvRCrROXOsqp4GPyvdR75D3/GsrzvlZQqhC
/0OhCHWP1bNR7B96frNKRU5pP7xYAxYOVYrWW/knDlT+xmvgfSuVUGqsQp7/eNbA7Wy3YCOodKgv
XwUAca1GR9Nif91Lj1JAXQTSC62R/RSSx3Y9THIbp8XhT1sG8wur9j3aBf5qZDjD+Gq33msGWB53
hM7G1BgfTbrVeN5RzKT73WXbI7Pyu7vAZgCEV9ocbYiF5C2nbfeDcULprEHPjcR0XVgOrlg2XM58
jSXF6c3VeBa2cVhiXoOo98Y8Q+0JRsIRFPTK+2JuFmrva7Ae3H7EeyG1yFdKNi2rj5oiJSVF6cRT
9Uqxga8CsSWc+5ZOmYmc4v4KGQh8J7inSOCbbODkZJjMYMZi1FMiAzUqKC1txoWWIoS5ehhtwD1d
Nmmy9/+6FmPthqyzwA/rnY6+FgNiBx1GbCy3DlpiZP2PepAfIH0EF48eOSLNbc42azWWtU6yjyVw
tfgaZTIsqS7eabnstSdY3YY5oq7SA8V9eO4RgafEz6M7LDP2lJPhf/s2tsiN65wraPy31wZ/28vf
Iv+7KpJMr+aRV+pInpu6/GAVV1JcweFvsmfP1x0qmq9Ybk8qVJyAuJNe7Lpr+uW+sznZNU5Vx8bC
0alnZA1q5iG6Tq0IynGkBxaEad+bqH0D5Ln/L9SiHWtTa0ZbXYOpoQdbOORzgNFzMarJZw0V4E/Z
5xQcu59sgGUILqsK6ybES6tXxTmcp/97jnXp7s2stvdjchjfRtLsl+e/a+2CnF2bWoaAPPvrsknh
VUkUCm3blFVP7aQYEp/sASG5jqyz7oDkjrLsvH1TZxOhO5BVPYP+LhXIw8t8oOsj2reIhj1Mnydp
NH09tAQTU6grQ0c2qcK5SeudRUc8vomGnaVyr3alJ4Sw7rZ5ScxfphAzDpE7Odw3JCnzOmq01XLx
EnRvTA2wNh3jyBbDYgXieo2RE1+v4AZ8gYM1mULf0Q8KAm93ebGd3pHVlsFfCneGGKxhIcQwUEef
wg8tq8gFeZrMQduD5Qp3yFJt7pnPnn9jkbB3zzHq1jv84OxaMXLCr2qu9kv6NMyL4xBQ/IWTHqXH
M0JWqll2V19oIIcJ7nXxsD0zhTjGgIHM17vmqIzJFnxAR51fJLzlKKQ29b+79PYhlDA78yflypWS
rbjgT77IGwLcLc1C6KEWWoDsGXP871DoX48WkJFDn54NCGASvDLtBZzAc472ESFqHN5Fq3b4kPuL
etTlQOncpVSyLyrLcuDa4Ecu0SHwER7JC+ew2u9WPaeSakH8c8s41GFc1nFkHbFnkBe78TB5A6wn
qtcLHOi9LPapiQgSs/2DZGRYBbheCInv0XCltHylTq3jVpkkRIk7/8ZpvQr7DayQ+FIUheiwF5rY
RaOflGrmfO+uEyp9mnMKUFDLqxnWTEd5FjUdYrYnBgApsZQk7yPepveS5g9Vb3dAyaF2L1Ug5uth
HlmSY3HQyh2VwCLOC2a3QT4IYvWcBr8Ai6vObLpX29ibTMuRe9cxP+2hQL2Cy4x3UPCFkyliJQ//
NGV1/Uxt5gHFWeXK/RrVRH8RIZ2pmA5eIE1WHHMlrH+jRC4mnIu+f+qivFvEoDkakTQMyy14VrZk
7DxklpFyUPXPJik3Dh2iQiPRJchDEjUnEKQzHaY942a2RKJEi2rIp1u/mIOlWROkFOa3Dmi0Isuf
LYG1Zs0brHjYv18mllaioBlVb//PIsElTcZKCAbnzvjmA78b+vDH5Vjvuu5dAbflS29X8PD8isSj
YM4jz0n/NDX5Bs404Gr+ODH4+YvahJ2uXnbUKp9B87dzq+Un+fGTegKoi6AyWhug2EmkoraFPWZ9
qEP5KORKnM0Ga/j+uM2yOSmUCHNaNNgPFvDHhxuPcWhqermwPcABE3xhpgvyaSCRDFWb5vsE1/Do
DcPj7foiw0ja9U0+5OMrp42IFhpzKOs6vtgW7XV/7YxNrfgKr/mOq5Idp0v8utWH3hqYb4VqF2cf
EymoG8iSBnUG5NxUwG6xbAwjUZOgrVV00g2AhcjNnt+dEUyg9qlGzZlk30KLvU0w7m29v4rLNxk3
aIKeDm5cCtDnm1wTATmWEWDmgHQYfWTkWcqKNOfAbPgsb9IF2Bfq+yWTB9jkZXs7ddmlMOGQCn5R
9SdhC6joLLEr483VnJrZblDZ5DIXMpZ7WN4ZufZ5eEjgvHmIyznRJ2y47iFR6bupMVXv9F6l5gr7
vXcHBWRnjwu4QOKeFHIPwlTBJhpBeaKxIvvOokN61N+s7C8hRhpjyNK5G6hp/lcP7OHpOPvdW8R3
78MXXY2MQzYAZYHYyH5LMybNx090OpLZ/o5EV7J3qRoHW52b9YrIkZ5NzOrS3uI3YnP3a2zYTiCZ
K0Qs4vT5U5dt4HJuTsMg/QrC5V0OHuedt5HVHKoY5Q55lPDr3NDyQxnu7+2c4nc19r8qb57VaCHa
2us+vk1f2Uj22w0jxkW/R8Sd+suoBrH0350PlSH/BTXrnJne9+uZSHkz03RZ7iXoGTXpRuKfO7Zq
Nn05Cwa7yj7D4P7VEmxBNQT1bs4bdsTLtc5enazoJdCesIJ03FSSC/7p+rJA9o2J6lpWU8x6+ASD
HSegIKJV5BD8U3VFRt25XeQveAO9s6ldbFj+gLm0sLnPHxSL5TGIDTRkopjtAclOUKWOJak2VmBW
sIxWxM9IV9JaoJxRnf8W+QNsyxt8QXo2TpPWFpT5e0+6zCnZb1kh210BcMYvJrLA52308VHuzh6w
qw2bYMo8gFVrRvQ2+lvVNLmGIqGfdpEC6AHs07cNW11IHPC18mbVRYxK70PFjAGZ+1Z1i7WU81ki
A2kBkhPNLfQwRRu4sJ4dJSdwOMAbIaQqMq+CLl6l7ihaWOW+fMrIWnASYTtnMaU1L73VcM0t9Wou
uWsoVdDMcIrpZW6mWz096p+Za1jx3WVVVG3JX8eI8mu9Db6bleRb7FClRL03XnGdQ2lFYKnyvpW/
XW+U2Y2RA7z4zkmIEyEisIiCJHXXp62khESJrzoCcFbSBiYqZiWqOY9SUc+yOPYl9ryIhQX/pDIK
ol39S5F53qKSqKUyE7mxRjwZ+galt6VgKJBODmOG+gSqYcxCRCZ9mggD/jjhuK+RQJ4/guAYqrdY
Wa8P3Jmw3hdC7bV5HsEspwSwUcJKBhXDFsYNd6GKI3RyI9LfJFhq3r7omq2JoxSTvuXOhXmPthLw
3V70Y+VG95QsKV8O3fjBO20Kbii2YNUJX7ydBB/ZmxiOOYHIBNjdh0vMGrqbtvxZDs4FNkZn5PDD
WgvK30YBkJDWhzaYslan3rz6qnPqUguvj7DJbtsarbJVZOy+KXK8UIpjXt7VQJJ2qb5BEM1ylzZ+
PuqRwKzVUcfnftZmtrMPFIuDyN3NHBFmO90Iw+5NS7IdYxTyl4oPwxrYmooAQtO3mmnG/eDu9hIE
O85blTOOUio8kvB21CcWMzHyPvIlkT7rclhxCSRLc7IlFNC8TIIM8Y8F5kUyVMAS9NajShyoKFfF
/ZyhDWFTQ969y7RyMRdRGzuOD40qMRodikxkRMntwO0iFOZi1eUwubo9VyZhcOSDHJl7zFIWsfk2
aTrMAh1xidQmIsCmoi85nCygSTym++04ua8pK1jnxG+IIQULH3TmLkQHzH2qAkqk+xp32u5w516j
9RC8ts1i3KCGJV4X8QkyERi3pM0TO8WvPsqdHKR8jDJSBM0PALHy59Gw9QMltfUnmpoP9N35XnhT
RPBQB8QjnpxTK9XjFMIU5RLXqA04m6yqNpo3fuh4B5ApPv5FSq34rX5l0EFrddTJYYncaXWsFTRc
nKDvN88dH+45gpITDMffQYLLxK92/bsws1IgHEKVUdviY4TpjpPOw96IgMl25AVXRSWXvpALNSvz
0FUgYD9v721ZULZ3lLLMeufVQ3zjjx2t+RZqdq0c/66HX9KCmeipb6vKmkMqAbP+NhsY8ydLdab6
aNeRhreyu9wVnPqb+tWAGer7I/hnbtFss4L+PqVZOsxn9FSFr8SU9osqYlMy0a223/UvSeLslAlA
obRr6wnXP3mIkVMdHBIsHRVfN/kECFls/Xl8+63fPBTnExmMJLm1tixAVoh05pSboFi+02ncl35Z
54tcH41U6xgFUABmC1fyk+DiOV9poO65f66xOqNCODmTC/RCfJrpDW39Ni9vy8Gy3/LkAqH0x1hx
zwH3B0Cl5ivB6YX/TaW3kh1DyPFmFCZD1MHoFf2ZUtAMwNy8htdmSgnOMbT31OHLu/DYuoOR/46Z
LoLnpKipBwuFO/bRpiJ6ygeGxuxpjd8tn7UxRh3xP9Hl4vysPVc+fHhTKUHhZpFZrPANYWMk3JVm
547Dj3krRNrtG7uW5Yrb+tAmUly/73QESh8F2sCjYRzePo1pLtbO/ejQgy5e3wSVlnI51GvMV/v1
kx+h1Dd9AMoshiQUrU0XxM5N6QKDwGZ5+OnzjlgD5wHhvy4mzZ+qUixYdiYV5FCtorXQFz+aNltK
SW4IBEgyjNm/UvMknFfW2pyDVt1KXsAZlll11iO6rPdp3S9ABTw6uYZFk0itgGpDVs9R/MihzVn0
pfzLMApxi4FrHHhc/NqQy4Fy+nAUaslR/FFB09t1ijIpZ+5STcrOOXGHj6Fh+okxywWxzD3ShdEA
wbNyxKGy2EOXP6D6l/5dpyjEnlMG5UV12bkVK5O6RVWqg/4BT4N1CyfZiT+B/tNGTHAGNfuEVCcO
XSqaGOS3jZREiEEen/cZc5AeLZz/G27+KvX2v6hkw2+/INcPLkOtnaKfw/X6sllDDp6RFd2fsUZk
+ZJnGTbKN8MleknE7DihPqEQp0ivdWI+hw3SGBW+Z33Tc7T5K+kPNhjnUfKFR+3Q6OKWIp/uES75
za2rzHFQkb/WAurpnQiKsd4SsbPXdjdB2+OFskenkiNakWUn79x0+b/yTub/6Jbq4LW5jEoGx22n
BYZOw2r5NIIdYCBqzotXYRs5pQau2DcdxgkOVSom1xf2dQ28zLWW6p922+PBnVwy9IAWwu8mlTtp
bzzr+Qyu6OVoJ2xE1a6hwFFWcd8w4P8fa7KOcu9kOiZWwa7SxJzJNN3YryOrk5nHzjDyDN0z9Bat
uGDv0art1Ng4FkVmQmvVMgftRsBlkYNS9OlPHtijzPzPnK/QTeJFUT8xRbkI3FZP8RtJRy7ern22
Kgun0TG7WMRrFn++jmQ6Kupv/0x6ko4rE1XDhBhqaigfTzWZ4cWlZZc7IytiJTns30oK+8xLUNFE
U58dV/LqoqdNBVLQnUVIpPpyRDO0HzH1cZDBticiPGJWf9dMyo4yFhaIPzQ9A1W8jraYRSIgSiQo
pC9pgXOKGYuz3fmIY34NNH73Yxi1IUQYeo5tuCNuz87dOpCXqfHlylvaXMA8jKW0pzBavZjH/Zj8
C+ebwJWXgf+yT7KVJqJ2Grqq1vwou3D8g0lc3nItH1xeEsxw26qXdGphDEpNSikOgZ5ereapLrO4
3cwAxeBYfMso/SK2NGY10JTsD/hTPC4KVJYw5ugojlOIC6ioUFfOntRpyGvZ8hY5F4YzjSQ/5044
QRQ5qiWE1PcwpEH3dKDoT7s3mPPiRPfEXlaC3W3F5fBcKpgO762UE1ElYSD7LPQ9NqFKuTdsFRdQ
8I1fQwsteiHIMFMkzqToQ8jBZneF8NvQGdAeHfqelbobxw9rxzHeAYUT+tygJc0GacBlemRosMev
fs3rxxFMKjOAjCZH78d5gK/c8/mbQSKYmlzogKzHaVVH/tu51rLwSMzaDJRFjov3T6RySNCdLCm+
SpnHPU+mnh4lPcfinNNtQcUcVea1r/V9wH4WlKRyL50QNr/rjNBQ8+65nXLfbsTvd5/AY2dmej5m
NLRlIxiKeCUvYuMJwZHi7642i8Hg1sfftqp1YQ4JTYQhpdUYXFAtPkjyrRiB5nh7Ryxg0Nw8wnCT
FB9K2iF68F+BQtXxGwnFoST0QoZAlOKfmFR3qneRyOT7WUqlcFCktUxJLbrHH49iX6mtEEgHuiHc
bq61vDTOSKxhZ6iOHDLp2nexvaW2XFYXi0lz7jUrrPaBFCU8HIbxmauT0zj3kaqg7lPL7mS94uAv
95l5tk5xNVg+kaTIait1POnfZ1wIBbbjB38Aq9x0YcWSQi1JMV88RGauTbueGLDI84JwstRbz4jj
/KFf0z3pdqmeCG4AQ8Abz28/Td91kwCR44U4NctC0fy+zTxqDRUkgn05ZbLZxXF/BEb6woyYye//
woTT8V8riP+0YafaPd6ABpBRdPazpeZCDD/1eJG03SFeZKeKaEtEu5vUFgMBEXuTH+j9gBUuUZOP
oxFsch2EMpycr1Bl0b7l4E8TJwAP1hu2UWierfs9qDPugzCJScOHPDQAU2gJ02qDQZIAk8kqf4jr
B9aiyzJQId/Cb8XRhhkb3eHwW/wxInJW8EZT8E647jc0qeKcYTNWvhi/OOyAM2/VWEF500nhe9sK
Z2s/ueyo1KBBAjTRK3dozLikw85+5LLvqSyhig0UEgWfu/jkCem/2uneMeqdmAjV0AHE70oD1Rox
54asE1HHtIorentykTQ5M4hw/ow3U00U1E+gZ2Uthn61c68sugGHL4mntqwDeLxbsZr3pZpL4Z4d
wwY76IJXylZh4nyBtkk4QxsU1KlnsWa+bPeO0lHMDCNWsxzOWsbnSdcbM4DtFk/oiTdlLGawO5ZE
l3i9oasNI2pThE3dcq6204m8uewHdwwLOvUCK+1I/594m0qe7EJbD4TboGfbsybO3ALk/v5MopDX
+JdXHGrjUpGig6E0dFIb+oKwYL6bxAH50w5XWJJFzanoEGObzKRsc0UmoM+xjBtvi8J5kFj6GtTf
EbWvArLkZf3NMBHYr0IXHs9AJSFoeet3Yyrcyz3uhXDMXlcrwNDS21TszXwhXPlM6Q1x+M6O3KTu
1b9mlLEXSJVzLxSWhS2LOzA47bGwt3YJ4CME0Sq0NyXhh8Oik0AjgwYq0TNKkRvs9jmu5FgqL+X3
Tq+auP6bFyIlP+ATIDZkZmgqqXrVBXKnEH5/fqvdLEuqyFXwPgc382AQGGAFDuasx3fL03FS9/xB
8A4dV3YHPcLfqN+jcPktqCsOYNUVpowduWqcTr6koboXKVj38YZP4E+x6BypG2u5W6ToRgvkCJSR
P+wm1e+muYBVWR3JN52yHHItVsAJ/ExDOFb61QKUJZOYXAcreh9sbQ7x18lKz9sk+Z6OEve5tCw1
FZa10kbaTalWHZKZrS58FVqsDuItxsB84CYzI1zf4hWh/sOc3LibpFculMR7YfNYd1VFthwRWDIt
Tkz3tIZZHpX2Bsq/D7/F9LXcbBpx7NNt1yjzoj+Un93Rm+VAqei9c5qFf6N9TEQ8KbI1PtwEsI+k
rxt2JaUDx2CuMcXr3uaDn4Xrp1Jm5z5We/r7oNNksP4p2s9i/7/e6eg0mMoDT0gF/n0ZcV1zJygn
8Q/QZ0Gp578P4agpdj4aSEtVSuZJLMfZSW06zbLT1JcNjglQX1qhTCmQDg6zTXmyagh65YvV/65J
+aGetVmWf5KDF5TQr1x9d7zR+QRTY/Vfv6jmbYamz3stM/r1YSGz7CSGRaQ16mziD9ckWAinj/8Q
8L+/2rJ1TNBXKutEX5YOnhopNiJ7v3Osf9ow1ylwQ0qNmzPNAbPzBP4ESYkzIiWnGYEUFPgbtong
j8ifhirN9Gy54qGBrHAa10oSnlHeLLAluc+ajT7pyiW1L4779GZCOI8W7xhnFTlw2FLMtmP2gADH
FzOeNqiXYG1Rs+29S43DjQusrdzmN/xoe7m/iJ3IzNVeUMyI5P8W3h+VjfYE7X1nqh0Wtdtc6JfG
cMHUX8CC8w64OJbhEvIorgzkia5dSW+bZ3/gU+I26tMiSm2GKuG05/YLsP4/8d0QUQg+7Gr88puO
DIGugshtcZ6l2gyHeBYCV/sYXbDcYvUnEUcmmQGVK8FdLc66NcheH71/yAujIEx/wrdQhQ0Y9NW7
LglcuwQW0DRnU73luRhxpZeIpx+0iKX9MlYS/tdovPJqDFuFExdDQJWe3BWx/0uoXGkOi8CtGtjd
HOf2v5uOSN5nYsCteu4G18vHMVnNiKit0azvvfmL5DfikEdwaNYSYtBc6lyS+hhDtWsF82VYIlD6
lwSTYFVke3aMT8CBB4QOAqJizs6NWopLmJqHpGZ1+PEohDY95Z5c4Fm/+uPiKZLjibOPpwdyiqQV
skR6LOe+WJyPqwY6R8tdVrbBGmB7PPfR1ZlvLorWdhpF71KlA19KRfEeV5qbWfh6ZjxVSzBPpTch
SjBE+zQNF/RXrcm/g/crt5hE7i9hqAWADTKBO3y4R1my/jUgWQYrxo8WKztvqDcyExg8/AL46riJ
W6xu0GskWDGg0/m6MUS4u3Yp93ZAAiP6LyeDFgLHUEZt2nX+P0+X6F35/pSEMyAQYCXMPS43s/T8
/arq5rRsS6y0sMhV9FrHB7ixBPuhYu+hRVCgu7cQMKDEYnPENJ/nVbSpxJg+Yo4SNO2oZpcmKH3Y
7ntI8htGN/YK+IImvdjJ48vYtOtjYN7iBb2ZrUrgY242VGkqJuG0FpNZ8JBmcm6QVenziHv7LJel
aXpW06zKcdFX6jjh7Abp68JUiLMC3aRFTDwMpxNXwmXhIV193Ld+HS0wMMazYZes+PT7kd1CYWFH
b+ed6uoGPTU3QaquDWNrn1vl0PSAiqXH2eXHG7hYwoxWRWVi5AmGRZ2qLVTlv/jn4i7dMVKmyR8n
IWA4H/SY6ZhPOfFRWuOSE1mvGSTyOggwXhRrzqKmuBp8OZG1tsdOKP1e2mSLqXTE3cQAf4TYODY6
VUEukQT2t7CeG7Gd6t9sYDQqd2GvGcdLL+14BBZWJ6qgpGiD/gsIcLe+jalLpYsQfcujs3VmCGPX
rHl41K9aqeeJ6PsPUWp2HiKeKzHCveKLRLsl6VR+gSNlzR3Of2dmw1w++U072c7GqVEOKjPDGVgb
XCag9zMD9rZ4X+nMyOJzt23xF0aZmFhzQjgucw5h494j7rhwACh34VhKNmA/3n/ZmdBIYMKF5/Mr
SVjKCoaLvgq+nyxWuP6RWcWRKZh4w5EQLuizIH1PItsAXJkRUl5Epii35KO22P/FQ/SGDg0akABV
grJqdgpgdNJqvt+vxw4ub9y3qCf16tCeCcArfgPtD83Tjb/t7VfcoBcm3aaYC59WcM72TYUR35QT
PfWxs7DumxPLCZF1NlMGsjz9k61lKcg/E7dp009/soA5SDLzNeJZ45uLgquF38k6WvGqlyi2fXZh
6PrQpnSoEboEdl8TqwV+50C/7ip4wKYnhUwhYWRfP15ufUXf074oUk0SHJA8N4MaXxed9WRQ+yUC
54sd0N6O1MKFSZ2m2c18SqHb02qMoRGF2GDAM29ofv3XATQdozHoHfgL8MY/UJLjm9Bd9tWuAWRW
e9ybWtN5zEpdzdm0nf2UpO5jljjugpiBkONgn2FizSPHT1KMEtay2v6wDRiVvqXbi8YyxVijdJf2
AHyQw6RuTS2XJ3FXdmjAOfXgKYyxJL1GEnOjjsNI/zsstkJqe2/EvsfJfXmLn1RHq3DZp5jmiDSt
oiyvObuvbHt4H8hc2E//t5TiLXZbGKy8U4aQV0reVh8Wzrz5+4p4qc8En+y6pqGoE9/Z2aP1rM2n
+iXZsIWXB06cAa1U437gsJE1aiKt0uiL9xGTf44h0q1AW744I5Soq+GW5y1S5Ufk3RVC9vCuFaRC
gQoSNZZy45M5bRVie+8y0FPH1KZjy9WmwVUK83OcvLJU4lA5bsV3d/+o5AOreU25uzu/9MKmFmYM
tXoJb8ToqDttFSgVjuAeBAr957eaVvR0faHP27LX+b0K5PngGPxgvCXjzpxdiqlivLaO6K57YGUy
UVAuhlK7LBHXQIaals5g85HxSboWz94SBwCJd7mmceQkMFpYNjBRU+bUKJfUMSUgvqpRPCbDarun
nZmZZ/2JViW0+INsO3V0JIjnCbB6z5O2Hi6pGxuEfSETklB93XVaxypbwdmMrnAvvnt++r1HcZXr
JSINyKv8KyoUlZ7c4uB0GP9NqQNnxv4XpFPlMIdU4yFF+VbpLh8tW1adwwUCZqOzajD08j0xo6c/
4plva2EFs9hc6NMOvEHbGiYZpenABK1pZag7XcGR8ijRiVTG8H4DA5DRond5l7TSzjEAHllj1ruQ
3j9wJJuXkzUptyNZuOuuJrCKF3/6G8ipcEK/+eXKKWzFgnWsOtrxFLso+SNtIKRMInud0ZU7afq/
Z+sgGL6sfLt4x5VGRcvVYEh557g1g/sWfgNnyuZQRrhQq0/1h8VhH564fSo72bkkD0o6Ch3tFXfo
YhnG2xnL/NcQw5vesyui8OptfaUQKochvkWL/n3SiVc5BGpcpgjwwozM7Pt9jrJNIQr3/n0Tomqt
HWZcbMf9Q/oVzdHo2SNST5sihpgzQk476SmOvdp7uIKdkoLnEq/J/win4SHJJCqUoLGPGPJ2BgRr
yE3NbjlzMK3TlMERQb2HQS3HZvsdwSDZgQM265AjKjqGO/ajuBA4W/vzkTEE4l2LTjLa7wZ+7t1+
Z9wA9N/1ojZIzXWJ4gZiVm4bu3Vrvnw3IAkNaGuYsTrNP0t+TbrUHhkZ95Md32egFMYwUZDif/4u
NBlFuoiPQxT51zgZMwCyZ5+B0NsOmTi0A6dPLF2nsilLRtiuFtZrO0tSeA4kT4pe9SJE16b0kPCg
WXNHKqCTnkCROhByRzgvctm9GVp4AcBALNzc97O/yM5VQn/H30RzKnFf4xFRgMwPrcTU6xSzj/4Y
0K6G+GITAuSuTE/q8oTzaPfYqE5X9j6t/6/SahMeZ5Jus5camZoUIZqVXzVlE1rDPEV0FZHBIEw+
wCrrTli6vg97tIXKvIipw7ATNNvVXArKTZZ6WIgGeeMS2hvD5ZAmW2eJiT3Cq+PmLMoF4BICUwN9
K9spncj7FYSyRyfTb+IdJCLmjgPI50RqqPuo6KkdtgvDCjeuO2QiLAgkKnn45OZrP0oSHLCN8gZK
tN5FIFlb5I6UjoB6UhtW7zxtkCVt5Ofp3XAMQtM=
`protect end_protected

