

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
YdpNuWNv5ANxG6sesr+pii9y21Kx+NVDp0WoJ8gKKxKHNSppxy07GkwBsVP2aDgHIw9l2ULLZTNZ
WthaAb5amQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
kEIsWLqGmgOl8w9T2kPb2uPP5XenCQ9kpxljFoCEGisg/vUEuVE5EQlDS3+mxviS53p6zH5m8hA5
bszDfKwHD76EbEoDDpJWL09MvEqH4hbAV7G0A9Qe7ZciYDi8os/DYZvhR8zjbLils1MINgQgL32T
+DXtGPXNuzJTAMDKzws=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
NxGGOrhc83L0V7+Qmwb6+Gi21+qsbQ+hA/5/9jysqY4QYAqiXfCrWB3N0NrVsGWuuTvZXoFNcxot
Izvlkgh5KOucyz0ezFvnhsYziU+FkvqQYf1g82Syrsz8zvyVWXqii6aXcF/WSMwXtiDjm4MiGpFm
yTcu8CcJgBMXYGVZx6nj+IgO08YgHCC4sfTqmgIgkxkmBrOsiH76g2hPxvXPgVWaBlJF0bS/hLIS
Glmsy0cU+pqQlcfbTEV79W+sXQ5Q3KPQFXj7AhMrHHD9esRm2Isg/tuzcRVk1cq3LsMUN//vGrfM
OKoYOozZxl1/IflxrtIzbjclaBUaFr5bvZYMTQ==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
dIJ+Oh/ID0KokdCrmxnp1QfFJ5QZBtIG4FQx5Pan4DTwhUxDWY/BQobSBBDXzWh1TT07UPg0V7Ui
zobKMfHgBNkMD8/PoD0AIDWLDLeXLvIJje8mGtE07uncec5mJ2eGa/WSy5sFj4M/Vdtk7C/Ab9LC
9qAaWZZ72ZUoEHuysZg=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
VglxNkzPd+guDL8DGRWVtgWGTdJbzbKKn0hBXJRIK4IuLrtOeezNwjLTIb0FIMSJGqYYwUrPN3z3
TVnjDJDaG+HA47egpMvivRkbnfO2/EAJtU7n0hK18OztWFzW+yXOUsOuQnFS20EGjEAN6HCMCAXS
ralqFAJsvMtY2y3dJNuE6ytT3WYkXmZUpTrJPPJOu2l9mCOnHkBU0dRG7RNYXf1tEMPaZrHSYyvp
XKWW5CTowIM6jJQxDVSVfwprGmWFUVJFtAmp+65D3ADXiHMcwre5cI/ty7nYS3euq41mrkrZyEF4
iH4/gU0xN9mM3aF9hBPzu3xQrdML35ONnUZTzw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 13184)
`protect data_block
7oWnNFlwPh1KWuKzjjICo8IaMVbWZ25chwk+X3cIfHUqIVimxR3Itt/wvWabsLWQRNHlpY0e8xDW
BXEUwb3Fb2p/pRSOnfsVRcTOAWPedELwamZge3Nti0tiz5OPMx9Ed5S4wZvQdHLYEBskjPw+vbl3
PlgD4bRbsZnBs77ER+O3/9CQVHzSNDyYd87YIRSErL4N6mOkQplG9DqIpIh7h9ECye2AQaAjv0Yy
kO4iNzPp4uEXD5ZpQYeRjzSG5IkFAbpr2TrUchhhwgNd72RwjrjxxYJFG21B7ucuDfsksrzrW9o/
Ox29BnGJM2Rd/VSOPZJ3rAwm2wvs6e7ZFWfCZv86iqbBnaLLh2iVRgd+XfnbSPqTiJLNCo2OrFtQ
IDBVi/0O1RpTvbQmj3Bkl0v8PaqfHU2KrZ72Iw/7mORv23MsN+ChOp/sHyPZZQiQ7tVzWSdapJ+Q
G5jVWyvOYoXqad8BMTg1Ftd7tjQeXJcxWPRAjKFJjpAobm/9FAsiHfhpEzo8W/SjS2OBHwOHZvC+
ArQTnLurbdLjGPUTiYRvKvyXe/3BxDY5WEE1BCl1bKtfYzWPYi6B42Oo6lYdh9bRv1QQfoDXIU+h
LcpKTr6P2xrKfwANdOd/gkccalNkTodCMvzxTy5SKsJIhR1pYbDcyAAlucXwBuy3CjwRUD42T+mP
jRof1jPLL3saCXgy3HWHGwrcbk9RBiL9X3LlehBSg43dUjjnZyuTLWwXr6a6aGiscIAP7O5mWfny
H9+zKrbc81qoxMqsaWxi8GsVoqE+rRGTCNjKMCNZ++ziYaVTAz9x8PnjrFzKdXKSmahVDt/bnDlQ
wIauggHP98fGfjZLYKirKuq0Y7vqKlfh+bEpEW1M69tUeIkCkkE+f/iCZesoU3bNiY6RK913rJ6L
QT3fpBgzqtV8s9E7IDpq29UMyG6MsmINoSkNOB/IjHMFSt0DeLp20KaYs8EPIGkt4QZHBEhoSiun
60aopJ0mpSRbSWJUxw9d1C50wheDy19BCINUCgMBdoSzW62HwIvL19e3PDUk8Y0e2KGw/POXH+eN
sfBuJC+CzXULWI8oRUavo93w0bwNOFVx3B852irZJBf2YImWUbwE021M4JCHac7uhHltL/JvotC5
FQXf4gEVXsy4zqfwInIBZXiPDbnXz21NAwJgs/7gdhzumNvGAhSVBNBMg5JHhKjKuiaCfNCifPqd
lD4KHsMq9QhSjlebfk8ptK9X9CtrsWxA8EUSCzm+bRBRDwMi6RsX0vdGQPa20+q66QKBePb7/xH6
Xh/haL+fewyS0RADh4tEjwTGXJ5tgOws5gyPxl+8NbLkfwUH+9OVizIaW2U4pi4zIZUk3MN21YSw
Q4VmlOTtgLVylBjUddfBNWRW9BPGJ9NqT7RuyQqIL6TcxFTEUvQDaZouydzQd6m6OFrmgksbzdpd
RXmL2zvibPuLvM45NTpOKYm1ZFP4kVUsG0EM5CbauCAn6wQ415KQ+yvw9Pawy3IUZKBw+heMu1Vy
DNuPPXRRNKlQerOvDyt9svRJHn/B97Ya8pH6bDN7bWahm7/Rckty9E8wYcP6JAASK48/e11AJreX
eFIU/Q5iUExUJrnB7c6rCUfasQOdBlBNs+9ALIWqDgdEZTi95zAGRk3uUtxdwdtYgnN2lLif8A28
BkySPAQu+H9kqHEaekNxKsBDUkeOSxdqP6Bi1P+RFp7PEhy9Bu/GJd0qjUgL0PnKdjSJuXnp5PTq
/KtWwYw6Dd/0tfsVZhjwGY7yfjHB/yhaUW5NXUxUlKU5YVTcGzSCcM5kQlxG7A0I6FUPJHFbb/7+
+d3jp9Epy9w+sC9vtnPAbPmzdJnu6e77+Idub1UQr6b5dArJw0QKWwiaXjRqcbrxPE6DHWDicK2G
VWvC+ooR8KnT5kAggNdy7t0ZMwV2Fugt2CiedWuBSazHxl/Gt2e0qHRrUC2eYdqlAQwFTQ6B1wl2
E64yypO3215m+W05uu1OOpY0K5bL22Rk0Wjpv55vWgh/qBzuAAnTAsSd07qcZ3n3RBD0R2nyWdeB
NoGNiORTt6uVXUmCosIlU8qb7dsjan1cg8Kk63Kv4s7vFG2sp/M5X20viasyYoWFOxMommGfIxtx
BRjL77+FnoDYxfL8/GgjJ7kxuke2mxiRgZKvIxYQyKHP2xz1aXpBZl2bAUFSGl1UnCteK9sqWYMT
o/lsSx5kw2whOFQl2anw6uLajiHFYwFY7rLJsA64xUeu9cCiVdI9y6Mb0I2IyVe8fXcPiHrHE3ny
UEt5vKeEd+wizpDQwafDQfORFJm3zHr0LFiMq6dekjjM54r3UWOFxSMl3wFQjKIdXHs0Yn4Y5Dfj
tXDtl4f/jeTJWxUaBJmdU0IERBdERbOO0a0V2Eak/g26pSLR98VyIFwlnGc4qjqaY8o2+qp+UV9I
JXRwQy+bQzFRSmU+xOT0sj//HoH39+l/gF6wVO5h42shVUn0I45eiXZosixFcVATvymgMjLOarVR
XKrbZIZN+DeiuiMbdxN+5uJWxC1SMfGLRnmsi0/2t2fCNXU1JP4u7jgWDJC96DLpgIA1jFioXzRI
fExGSHXhVxIRs9333VvgXpOcDOXUQDVVHpvDAjul80Q4Ili/l2HrJcZGPDj63fLgPyeSZ/fNSfXM
q9ucGD1atzWC5Oun2aFB3H2C+Q/NECgcSujos2D7ZnjvzG9pIL96nigbMZVAQ6EF7dL+Sz6HtkqJ
n5Ppc1vo5ElV88eotKqkblvpz8krrUO0qVUqkVqU3TvwyFPe+uXNcLW2PHzc3c8Xs70v07jgl2H6
mpljF8bzT6r1wGHvUBDjX6e1YzzqusfUnYfEvIq8KMG2udrB0zkihWbR4y12xyI1VFkZgphUuaWf
6jVV3/oU2ep1LrwRAzHe/e19jD9LZ3gBPw2ogzmgWuT2tySNupxZ4ny6yl8WJRI3znVk2mOGm+Hu
TWMtB3YPDLNcJRP6xn7IB5QiyFNYuA7KJHYI2aZ6BxoH5CDAZFWnacmuu2YgG6I8JsrMdmiroxGd
iUttZqGu0DOrO+qf4VvPv7k+KFLOW+4zdcRZ8Uyf7bWCN/AL0zP3u0XXLpnreW98JW7KiUgxyJWd
KYeqWzM2L8nLRQL7Z1KKPGo1bDfgDKBRu043dBwlsfABcHFhH0t41IjA5RypHSREyHZJcH7Mmt0L
PWcJnlk3IDIXaJmIQkYmM6SOiRMWAcDoAzsaioFMlbh1xgivxXCXwxHu2ca6AWzsFN1qtDjwiqg+
uKN0Mxc3Zf6vJqvPMmyZ4UseT12tzXuSEAw18cq7zPdFnRdQyesQh4qxL5BZP/H9B0AuTClzfll3
vqXyMRrkx3a462M2uocHWvB1HsoJuNlbQVR1+IOQdpYvRKoW8Ei9q0SL6c3Sx4ms5agnsLgwN1ON
cis19c9E1xALPy6riSAercULDViDXt1CrzQ4p14qlVrLrN8ReM5EW+vMsUQ7ZVJFPWe37isFc6Aq
/HJh3IQ5GvP++iPq8wVYx708Wy7tnW0cHVCado0gYnF5pLDvNYiSQSJfo1JhXTPdO+DvOnRZk8t5
FegFxYXfFQEO+LHo1H89Vxg2tlmeoiXPmnJ9m42z+1EEdrVZO355Ow9DK4vXypL/et1xkEszYRMQ
0i17FrsH2A3qkx+nu4tn81OPOHfUjJS5loBmjZYMLztaT92DdlCwGWuhO+6Fo/MzyMoKYgm7UBwh
NI9X8wW0lBFHk1VaNHFg6QGR5Z2BT/oQqDiB8dtrUR/Sn5ADK/43BhNrLzumEgHoxO660iEDIKNi
JacvDScPkrFZwI6q2IL88ApFAZuOQj7qhhqgYunyiex6asMYdcPZcp9y9BywKV/xLN/AC2Lx6R0r
2ICq7fN/IrY+4hlKkEQq8SU3Kn+rb0UjVcwgZr6DXPLmAg/FGg7Z1r06LTRUucFNFvBQRKIN/r16
CTLbnDXgxP7a8rai2rlEOz9vqfb9E+zf5euorvzBwtdfKoUVzl7hcmetVYpeQyyjOKBqscD58RiD
6k3JACaaHYmN+fx38OX72QBo7Syl50fbEGb7COTdHo8RgHgeNPffgSHmM0mVQ4cS5Qc2sOOmhedx
uVp4o8WnXp/3hlonz4Cu+2bptsiKVNceI+QLidePMhnn9b5U7q+1YTFSoruc9ifv66z36/25mx0A
gdI45kqjKDz4aeVpvkFTuXyp6pDIVZ2qDuwmicsGZVGdvAnRZ2yD7wuHd3k3fFbFAg7kgAlyDnX2
tfrbK4Wgb7CIWZhhg1Am3uYcCUbTrO9Wp57cDWK9bco3dDABGEFbMS9gU1CvcU5GbN3MZxy4iV8I
XOI765IltG607+Vi0LTski9hEC+JLjP2zESQ4z7ydlCPA4k9dokyM3hxwF71r5sMlS/jjh2X1nVg
r7XIgL8AqtJJWNbIRkvO1G5lNRpjs6TH9tXKjvIwPxipYK0MjUMtaozmgX4WJQ8Za4ub7EX3R9Ms
8+xEhdhx054FXMgER3mE1/GGEvFDPxBkHr+JxtR7a+xxR+PGbybzNk7PK24oZKni69f6Bcc48xvi
B4Z3qOYUTzu2MbKz68yMl/hpoCWxIAJrGJlroWykKXDj46CLiVUfvl4A28Fbx7X7uWMIShTxOeDS
czN7gRqdgjRJ2pL0bnA7A7OiokrjvPb6VGWrisHuKzuSItORg2JD6WQipfUwGvgxw8mgraiudLFj
uIrZiCX8GLgfJ3+gwhbAqu5nocNasmSGBOtxhbGgq+id17rhs8hNyyuTS9IyRzgVXosviWlnkVL2
+qn4+2oyCYRhOeb3M/ZBScsuVf9uA5EU1K2ofX2Mqn716dJJ2hhUwDqnRPHG/rasbBBXa9PEiZrh
/gfIBD+rMVHhZSCCPyXurRaI/sILeU5IrDzeszVZBrNpaGjV8gSUsXshl40/7418zNkq63am7QSu
RThmGsY4hctbz+e4oK937QkAzRqyd/pyxqTcU8VEInouATgVaHxEpl7dqmeH81BOxRnHX0+bmgqO
ogyaKFL/eDdCYP3COceql7gGwskz/4XUkOHSSTRYQfrRCND/ZBfES3q01cJkwCvgwscvFqX+Pvyt
3bLr+2/RA2aIRqQYFRl6anJpBcBy/uFxJUyy3uyGaOIMeO7JLilHzFeAtX3l+g/ZW+4XrzqNAw5y
ECjQQWySAtK+EJYaSGsCgCz0ObUOBqzOjgVWWbmRlCuLAv1QWd4A+sgLVPN2dALDbGv0z1y6/Jhe
pH67YrewU0or9Nz8JDjaUqzyV6dastZ3i6p7Ezho+BEbvRV1lXn9fXWOaSbWxUmI1GGdoOsP4yUh
afndxTejzbEibXhLwPYOGtbUcAZcZ+rkDwwf6q9TPFnQkp7i2Bg/bDMgayT2SR4Mu9/ntfeArYu1
82HGEjnKcy2nYQnfs8O536NCFjf2HAmGZ1NHafOBnTlLokTVdSxkaVVozZektzUQL6zKdstnR6pS
gkhVTbmN5+uWhgiVRcmUrGQtNUFgOAWv7Zu1RQO4YLNaQtKsvEw6+EEKD13JFLtq2BojISwCQXVx
3SetRXsZgPNT5AlcqOlE8aSYaCRMO3IafBkcFOA2nO1N3HQL4C54yZtLUweTndfzU7MPLB7jQmzk
BWUkImMpW+ZVOFNTC2pWmiVf1Dnkjs3nPc5IaXmL8+GcU1oNRb8XvgsvArz6sEJYWuXd/jT5KD4f
a+ZC+nQm++bQSEgaIbomWdAgLIPuYrJ0jyYUHc0sCXyJiW/wom8Ocvo/aJYtwb+P2xfdHHnTgw3k
6XNnO1NkTEzM4kRWZilFxtl34D3KNOPnYzuIXTLajJdxt2RaBMIqOzKpnmJGQ2End3wkIF3J+6wb
QWn10Lv144p9ZVjrS5d7DfAzEp2Zjb4sVeUkd6lBORLeG0k2fMhaAYTkfVkjTaKkqPw+x9dGKL09
l2gaJeguc9AsfYKQMgY0Fl4spQ7eFhjm7P4VCJ89kYZTaWpDgWMMZXQdRMtUWSij335ASX1rBuZa
bwNxbtyxnmhNvi2fsAD9QNF/Ap7PkXhX3K797A0ER/Jg53b86WHA25HJub7ADy2Fv+Z0TWoZX+OX
a+umx13z3WG4K+yHvKP2mHmenBlAeJTTPbEP2YMezxG4L8IYil6oS8BmwIOj7Y83zCXWVyKOeGIf
ssW5QHUGqRPkAmQqsg6VQHrtCZt5Z5zZOvf3F0ZHMX0Y8+ijFkI1AckFa3A8NbsgH6bZJGTDudop
cM9ulkE94FGx4StafgHNzu/pP48p4ZYoyHZKWXpgIqnQjSPrrThkKcS0rTV6FKd+Z+XV8ODRC1Dj
Rsk6hqJJ9fcHR6PV3GC6N4DGqYzttODq9VNhsbVAxQcJcWJUaVHIQwK9TbN+wW2e/YKNivM09m4u
5IdH9yYBO3CRo0uTDKRAQGMTfe+KwEMCSh9P9Cr8nD0BuxPfUJg5ZROka0RzkEM1X60jz0UaH2aq
e38BuxtAq0sYIi+IZG/2NxCC7ZS+XjGEXSe1Yh7er1ynRg7mt5QbGKM/Lpk8UvqJh2J0DKLhPjFI
63wgaH8mfojKfTPEx7r+0X+OaExKIzapijBIwS4TPMUYDpTzv/R3Rhw4gjKGWr9uzkjXhHoCAcXK
wTN5pLUvFXcdKCVtzVx8hQW7HLDBl7fFZMtBWoAv/bsBsgj94GMgpCwDjVFgJJf9osGPE8sDo7r9
sm1VMk/r9gjyBuq0mDfsaSqM+KdGSf3IhWk7rXZUrWPzl7E+ZrEgfGKcwG8A3DthM94wnEkeaNoF
NcDGYgnzmlYPfm7FuwN17a1mJC0rAdIFP8kYK0II9O/gYMNAoFiNEABM22FRLTUScwSN5+XItZAs
Q2HRak5vJGO4/C5eMUILdX/c8xkWGD6ZAW7G3V+A8yn49Yi4ysdQWrxFaeHNGtSSOoWqXPtUPo+c
dbmvb95UOH5GILIhXO4ldqxYhpOT/hcPL+rZimiOahTWZTUImZuWgkYQe2FbZtLCbmr/DrWnK8eq
xzgN5fo/W56Pl+OKgS6H1lEMQxtivgP5GdOASuN0mVT69BNgtpPZFtwJ0KdDxEyFECa/TKYaXQ3y
D2DXXI5QIIrvCsV9lG2Gb+92KoeETtyXNVFnrWQ5yYZTl/effx6zBonoSIpb1hrC/Gkle7O2Sa+Q
7WhBCX0zSDUIxmlaoNHxOHoclmcKMiZztQd6Y/68lHlzkcBnU7PylsKi2VGlvMT4yrxOmWy/iJHl
VXCzJifgiB5s6ZYRlO79NrWlMVS9wv3WM9QzUy0kl8jVYLwVZCAnz2cp9HmFe3BbaZaNwEbIzG2I
p/rQzKHO3J5xEBO2BOMnm+cmrgRGJxjdNokOBQ6tzyh1VEKsg+dYsmdocODKdyARNdnlu1lqTail
aVT6M4y+ako40SGWfj2TVjye9zXNkS8FiOaTqXO/dnLLnuKFHovK6ABH5OZElTNZC49yrPAccsCj
oCgouTiAp9xoeWYqYxU1GskvUjhuPQvJmHhhS7ykRRLPOhpkzLKh03DC4BY8CV8RX+COuwf60oO7
Co4AZyOrtFhwqWwa3wCWcr1bq6E6vlUFLBSSTbD9TU+5Zu+60JHGviE+ancMrPbeIvy6sf6U8s2D
pszOXOPT1zGeFeb8eGmJCuQMbRmoTrKfWgc0EEtirSRmRehaj+GypUerk1UGo0TWZ606vrJ40qop
zS15wN11gJDcb7OkVWkUPAQWlbhABsFQAoYzAcUsXvxzTJY5ODz3zf2495K4VX8RLCx3CsHIgekK
BbvYVsa26dI0MQIBBWmqjNb4d6tmWkWc681TgN5aJoenXoOFTwS0r9W/DMoKMScZdsnSntUxMUwM
FWxso/retkrq+wztgSer0NOP7a35YODHaRksSQWitKFaRkwGPPhQenmUeFLpf7zEje0zge6GYgv8
3RKRWJYARDJS1MYMsn5UshsQlUpZRMOzD3qDsS1NOarjasrsWA6HGrTX3UDEOvGOVbuYtNZ9ICwm
6vYQZHQtSYbP8evdEqUn1E8rA9u4KXNWjyPhKuyVvAb059QwmK9WTKn1la9bvI4WLhmOzrkQnxRx
mtAdoScN2Q8IyqN9vz2mNNK2f8xxFEXHiFwezFkfVs6c5ZMiDIceKJzIPIx0jeoPJ+RFP18XFN+Y
UPTNOL1ZzK+v1OU4sMQPimJMQH0x0MpWCTSv+AUhSwZ9jd+6xD6TdT7trxhsy2000Oun4ccFPYzb
3L2+kOYleQLWmRurz8TxPw9RIXfYI0iB/rQ7jNmPrfnfa6qTIypG39+mFdOGLdFFbe3/lUh0EMSQ
RdUtw4f0yLeIxQH0NqribA6/OWC2IALacBFhFcjEShlZDPRXlcCK/I1aQK41XV7ZftNgt2pufzd8
yXaajTnv6nJAYnKF6exhea4hr95lUdyOXi9siJ/rT67abk0HrCLkAX7THXuKywIrZlLizEp+w4Uz
Dk2Td3cV1q0wLJbiroQaNJDkAl+BuvXv8LOEHNDzp5NNdmKNXJWs3mnBPfy4QuR1s0xaxJfc3T5M
m0g23mrUGiZ5p35tCpGsJYOtFZgzGf4P6XxvB6hYTP7+XFcQ/kr1DAapYTsRo7e4GdNUphIjZYYv
HyZmIRqP/vlLO4H9gCd0cRyaDIYZhp03IKshBOg2K0a1CsHu8WczmwzgsaSMwAC7tq5u7+khk1pF
uMDojq4nLJPiSOitNB5uJ8nVHs1upsyrHpV9JqTtCMle5RH9x40lfK3NGYIyUH4hmkjKZi0pZhOC
y5C2kgvfK2e7EslC+aPiON/Z0S/e/rBDKFhrT29YydpSyRqh0/ylTagLu7ptQmMaaIlSc4MZzP1A
vjNO2nGSaSOXIYb/wSBEFdsFSJHdAXlUyFsaQpMBFLL/wtg8J5eY2NdRfCiLotSN/jXim4GyqlMr
HCUMA4khUmdilQ5aqhCNT77lSeuhuC3RNHipVudpUL6TrFmtc4/HQHeEj7LGqldsbBw2q0PIKc51
wXBVkCG+YCdVX0er12SgdjxDYu9tZcKwVZwO9ehRkoo8NKoRMFtMev/FMCTsCDvz+KQN/R2wQgN4
LWosZSfcXwhOgvs9zmjqjdrM0N+C2uLEud3tHS3b5pWWKrxiEqr0bjirt4dAZRqwB86uEtgOMz5V
tR0j0tO6LUH88rqyjbnZMd9ezyQbhh/ARyn+odd8oMLvpcVGTJ0VgPWoQQBqwQC3SBl4o9UG3aeY
otpNHGco59yE1LMUZuia1kOBY99GUYqdwkOZdpdkybU22KGOycDQmLoKYdXgtKKmGa+ukzpeC3D4
R43/rdMqKM2kMjnVTZboQ3neLO5JwFNg5btxL9AIEBpBt0n20A4FHFFKZw2mmfrUDxCWwPAoWMfi
p4th2Z6H0kQ1zSqyjgkR4FpGM5DFz1Iy0uzgisbSi962UTsMVh1PVq5jnmeuRcZfstc4KXf19gZs
vIbq9s6SXMjrXlBT56eIxBWhBWDRIxTI9VN20G6cK/bIPQEUMCGkOTreY7IzNRT6ApMZGgSOz4vr
SQkUXawrShqZaxrVrJZFyOESFUVKiceC8Ue3t20654eIHEAn883fR+RLRvhEeaK2asnPIdetm3L0
tcuGg60NP9qEyUMEEtylwv1g9o+y1u3VYsRZREotwOqIFgA/eRctjV2NrJow3FFAjZKQYeeyRwlE
aOSxvFk+Z25LGAKlW75OeG4I1lt1VA5ymKFqr8LI05UodCONVoI9NK1zcsSsJAXVaWSBGMbq5dam
la8x2LVmUC6Q+CD/MfqZyTY6f6tQtcXXegkkgyAfyxFWJR6f+d1nTeVK0qaP0ySUJChmk/OEjTVa
WPomn1pzsoLfc7yHt7XjHS3la6tZpnDsm13akS4qm9YZic3k5zJtKy7I8HPKv0ocjSpIk4NJ0FuH
9m5x+A733GgxewyFsmVWCuiZzUePk6MbJ+03/8Uc4JSlqHgSXPZBC3n/s7GNRnSYupZRNHSdjT5d
ajE6DuS+N6Me4BIGRPr4PelbmrXu/UExTJQBzDDn9Ft9ni/AQIsp6e8mREgUIi4End3mwRTAd3l2
LThHkcM/VL/1ApZg3w5LVvgkRPkF/snuakEto/t/+ERHrhzqhEvaoqBJKUOEhYvmrA6bkfwLoXbo
syAinWgVk3NLOJqMmI2eO01cfB0+M5MGm5UHTG2RG/yTsYMwcPl07AbDQEUq9pzKyg1YdCsVi9+h
YhUt+rqfd2hxIPj8IoWt+USXmy3xI4W9ReZr1asurcKokeUihr0nvxE2cY6ss9JpA+yXCHup+923
fp3L+q32Vrhih1j3rjYYDR3lEUIEbqMJ1fUBpYXwtJtIdL4VfNofME7lKuCe9LWnOQZV7j6gh8b5
/SY2hcQvzvcH/2RJX4sA6LhK4C9EKcXdQtoypNPkf6aXWhhMvmlDbPBNK7QihFitJgNt2WcqHWzJ
xAIpkSAIzLpZoVrN23DfOtTNm54yo/7C1xPbcOPAaYVEBKQD7WnLusdvvJUcvNfoY0dsMa31pb7P
JUCPC7IFXkSM0FCkE8UJZPYPprEQRlRdZwV0+jPWC5HRA92mU306cEvDxtZ8QkAYKIiyYkSiV3oL
gk9614jxL2y9WTwSWyBJDQXpo/wyoxxhZaJhCz25CGEIgjOnNFO4Ybphb/6BAGKamO1m1vvTxFZY
P1RAa0ix4Rm2jXh+NIY7CbazhwgiCA47sM6sQmFRmC80ldSHE0I9zwPuz9kMpO2GqhDmBrJch1AN
8iPfCP5EJ3jjOYx9+naxktB6BNJM963MGqX7RivdsWvRkJjsTnncPUu3WbDpd80wcPxLrQxmsM+U
j9Q2zS7LV4Ar8VhyfU04W2wdie6/ldz/6fDp0MIkUlpj4reL6m9+cj1/o/lorsDRJEJkE2L7Lh16
PxtM+BExcGdD5FnJ168xgpZeupVqchFKfnEg4D4epSC1uNRiZN06IvzCe5IwVKjag8I1Dwuh975B
8FvFJr9aEGWrH9OLEY52oooJab9yRsa/mRegdKyuVBUtheJDqLRqpgIM6X74gKFPD0vUU+7hw/nN
gc0KO9/Xf258lGAw6o+jOgdU4I/0rslS6mTolcttYR30MK/u14W9xGfKsUNGMabMkkUqXdQj+Byo
w4RMiIrEj4NYBKqGrOTHfmP+xtyv3sQ3IGU2fqr4K0fugzHTkvKjHXqnEShTfK9XtnZTmAygYyJA
4C15mpptmz7ayPXR+DtLBuAIstyLJI75bxv8FJB4jP6AszkN/WNSLfGOypJPHVSY2DaPoBwR3LEZ
LqrtRQyVG2ox0CEZlxPhpXEe+rdSSreYgP1MRtzlrMw7szCYMNph6iphtFbhQHBWprNL7tNne6tY
OVLBHcE7AfpGT3p8w/jdlOBjrRAe7nL7503qftVp0GYKfmH2U22cWnCzZSqT9mC0UEF52QuKUkdu
WvDL/heyijwhGVuoUJAZztIPZE5e+5CUQOI+8dY38UznCR6DvcINLTNgyY4u0t2bMv9y0Tj4wNbB
GOGrgdigXl+kw2GmXQmf8/4B1qKtHAuJ7by/I7jkRcvwo/YUVudCy5a5BKRFv7HWjI8N6nSEaPlD
SxwisRf2X37iajN8ygUtTQC/TtGPpxd63LDD80ZT0zMzFo8NTK5fwjufCCrzbMQjd1s1cyG7iUnr
fActqoY4ZASjZkbDF+AyFF847RP3ojUB1qLeCRP5aTCtjckGmrOcptgwIvKf3dP1cbQWJFLeLBnR
Jgnq5545zSbDQzPgfNO+MPYVFMtiWc05iPhKue2DALly1gobGzOBeiPRMNVPLhcW6GCKeSFfogwF
hHya9YD0+ETDYcg3GR29jUNZ+PteWklcEQiVjuy7HsPyquJ2R77ONj38E/09fdvJE7hpySqhtLGh
5xfv6oi7XxiIUBf7QqoU8/Flm5keLcgBH2oBQq8vEpKK7DJXREHBOrnLzeS9JXgvbmkUzlt/YoNW
d8ykPbXyTRkZn7RUgSwozS4FLUJlapuvObE8cWkn42wKBLxw9pkv6tM/gfacttTjaxDj2K0wmZCk
h6/I0znEDVBMZsZ6t9UVNfohbG4pivMT776nZDSttUx2BraUQ/CGkm93/LpNeugiAAVha9/qAXfs
nDCx44uIa5VaoxHzy69z61/UfONZ28yb7MrS9co8k6Px+DTsCioUHt8i/Ys5BYUBI4WVtRzlanY7
2PHYH4ZLDNsxKXyeOcnbbNi1spYBGEuXllpy9vR0Q4yuwDW/vys4BDrIVy5IKEh3UQ7Qwyshc1mE
p6cYEKgh1gt9yZ2BmxEjTLnKGIxpZNcqm3bzruCKQyl6gTMKhEYeRUpSH0mIxgD1w8tISQcc2MMk
5GurFn/cSBizLZqgKbMutSGKfhQnMrLyATGBM3p8q8Sn3u2XjWJw57ju6P/InL+5ue3OLqfyZdpo
7A9h8B++LUKChNtlU+kLeh/7IkNMcKw3O9feTChF4KxJa90yK1yI+2viPihZkIvVK3AhLaNBm4n+
EPHH9YKWSElcsUy11Cee0w7IcrwKij3dYIk0KLXVSGXELCiX6Hu5NJC8dnYhBc6v7w5Ek+yognsI
FnBnWLugs2hiKOb9cG0Bj5NUFjY30HVNFxhmSQlTF8QT/EUkmppsEXgj1PAHoS1RrrXIOXIHqqaw
r2qeo+Rt1VwIeYFxYEKZucjaNC5hj/vHrQd5ZQVbn/+0bMbLvXeqDbKhMIndy9CwnomkxbzEPOF1
rXcljuUINrxv4aSgLkC4sWYAPkyoubHX1RTh8lRS1BvwgT/LwQpNxRseDoia/eV91CB60ytU65D8
Z9YEOCorYxJZhKVO2RDsTLDMnv3PMqFx98qz4bzVdNxIVIHjdLf1t4CyER/hKcNMUFFGEYo/1p9y
L6CmHuhx3kh83rKjuSva0psovew/fZtc261f6flBL7Kg46H9I6O3AKiLcfl+tdjq53WbkVG9Th+u
MMihxztJaVKRb9w1P8duLB0WNfsITIob7Ttr8llZJnFz1tEdCDXKPuz3IxGoU78CxQA3luNM0XvB
bo9PnEcdH0SUgMPm7h1uqOoMh9oyxf0rBH7sV733hsLQ0hEhw0GKt4UWIk/kuUrerY+zm1ilLO8G
/7PKoE5tfYVYyGbygJlNDlNMQTmn/bdOWjnRUT1DqIVnXeEhGipGdUv3bL7yuDJ5fQ34KkwcX/7x
JO6zJDfKyO4DAPFItuBnTTpkdi1kyCmu/5y5TuN3GyRqENnhMLI+FPrAYNTgt9MZ+EiDBKCVPWBw
OmrTJyLQV4EccOnhZHWdx6hvxxcQ6E589gO3+0LBzlXigKf9llylL3iDQvBuCi/vSOJxCcgN1dfc
6mSlMvSXvlqm7C0xkN0pf/zqukTb4rYVoA06B2RsX4lep1FqRefs8N+OjqWeYN7H43F8M+vCKiaQ
q21bFIdwtEqA3h/mGRffsa1uz1c9lmdsaMf7P9CS/c4JoAU4+xUS5cFvtnbXfqLxixR3F+aGY1Id
1WxPSRB9EFme9UwFXx2o5Y77QGcRpU4lB7NcOtP5uiUEzg4V9KnXBLwWZOK7BrWExFGen+LUR9lT
tuJ3YYzUyD/VAodRzR7RiXb2MfAmbh22pddIXcTlT0FrpA3BdV5ekR25HXF46Dr9CjsY2Tt1lFfG
ELkqBHRi9Sb1PCuNDcC5IpriRKb5e6CDfT3icyXRX+C28/fGchvd3Jl2dvARypbpH4qyNgTmYwTC
vqFxufUFeYqzA60JwaR0j3g4EUq1OBvyg+RyB/wTQ7NgrFxtUkNQAVswO2Lp98cHO9vEuiRCVv85
J7Ss7n6b8IuoW59nwxv244mgIsP0zdltuVJ9KqqvkOTmLk3fSokKQLBxbKAmy+WiKmePxPmFPrqz
NFZ6R3geVg0SLu4ss9zPNnPUR/sms4IIHn+HeCSLZ91iS9Xy/9yWpoXMVkySpgooJ6s4P8qR5p74
K1aUFa9f4dM7g4gikgwJMOCt+0UP2WEfsx88+htwZvk6P3s3dIZ6na5Y3w3sHRymTAqqUNwCoJnY
iqUx5QW/DAiDnnMUxO1CBwi7hEOZf5powxU8XLhplYRSB6GnghJ+0W9K7FhmxFt1F/narPZgyOAk
ywD++mVMVJOcbRKX8vRlzfZ60t51RRo7jiarlroYaz4LVvsij1q5UtXRsuoLiNa0+XK26qZ7hdcq
/c/zVRGIwoz/z7xG8K+R8CYmiWRaRZbyNuGUsrbxpJvLw3CjSYpbrYGTtVAscW0cpecQGl77T6Cs
ZquP1MfHQq6BxbTTUWF+ww3Ab/VIeYjdSgKyClZ270yMYzSZEnv5DIQzpnO9IRaOlAY79C95GGxK
hcF0D94AR4G5ziW+t4Q5bRpr/RhN5RWfBwJAYTF8Erc8Hscjh/VlChTyWu4uj5GodAI8lZThA9dg
/SWVHies0xbdfgtkit7iKfCscOIupaWIpbWyE2+njF5FtmzEP7M3SLB2LbxoroXNWVgAkfkW79x4
RuZEH2X9IIenfADiEHDmXAu09z4ff3B/wZy2iNxR3zWQ7uOr07k6mWQ5IiLMki0ZVdR8ofuEEfpG
mBWEMDp+pkJ3bpnOvPkiUgi4MRva6831VpS6JxE5zci7HvoIW2ERPSNbcaIHzeGFa9g+rNqqkada
JtFWZHJ5s/S9EjRMCj6MfZHy5lciTN7dOzzzUMmumG0VveVsL2v10c20Z6XGUUM+LEqNkx3ns9jC
dhszCZq/PJqTZ+WbEYaZwMuejn6Y02kma5fR5MSsJcw6fJ0o0W5usxeT2O8rXoDCR7eslq83sI9k
dVJZsiZDJyR3ZOHYDzOzI2H0r3O4CdhavnEDV05eAvKc5siRviLRPEqcitMsNenWziRlSCyzaXIp
ytoiPgLsPgRe2XLnPL4zkR6MuyIDu2rJ8C8fpeE7HJ5iuyzk7fJZGecf0HW40+/ppKONvqmDR00o
qBfSh6en8eu0YSHqnsUKegmNK0melEfxW5+9esCkb09dqCoGHofS5+wFfR+RXd8U9mpsWc4ayTEz
o98mC2EzQ+ykqCrHtX9z3BW4R5qwwA/x8429TCQcJN0jyhqJF6KRm/khSxfQNT7nAfspCj7QDpOw
dX1KYK9VogNXXQKZyY7Uqzsej/WnG35n8eNtb+mU+VqWVdshKCXfL4l4owlc3pkGOztYYw+DE5Z1
ILNVk98Wt39tBjr/XaJh8yFH9Ttk5VcpG/B/OcGFWL6GZ63PymzP7TKxvGts/pVroXfcr43jqzZI
CBkzIpbI/IYbsUJtfK4R9wsZzmiTDiIN3FodSxBYV0AUEnBbog/EQ5SwgS6Fqi/iSIWBXL7PnL88
KT18kzLLMDNjzW7Vb1FM2rNc6k/Hk2JUAuyMk25BS83+WHRqTyBjocKrG53sPpManEGknrPpPaUj
JUCNVH/hE3vQQqNQ5OIs/Km7ldOfNMCrOJOIuqQDaO03pDHQiz5ihHRdbdKEcF4+W+lHk6Omml6i
h7iw4BncpZFR3uLLUwqi6RKXiORj+4e722U1uPo49g0n2NCCvnYgh6kYExLzAlYBFTZlqlo0O9+b
lOvz1XYgqGRQMdzuOoQhro6cHNNo8f8vAMRdnPWfv8BfqsKAmBEnCAoSFqChnSZbJ9qi9Yb06iGQ
88wnnVXoE0Q10M5741E8j0qTXDPRV473T04gM+NCUjmbNx+Ak9wTA1wTV2Dl+0uIVsEkZ9L9ynnK
vpz6B42qqccmnBoikwXyD/PTIuM/nAtiY5aJRDyc5ral7KziNl89bRQCEQaRJ/TK5vH14Sa2ThdX
JQwL8MCqUdwtn2s9vpWgJ/z3Qt6nfO24w+QM6irak+CyUPt94ctRvMY/+HCOExaUfOkT8fH+LauM
w2/CWLELAhpLXMXT8nhF42FmToZzs/q9bYVbdNnaSZsXrJnqMz08R8S2415nqAi2se04EFJA6Yig
4O1LecLuTpJl9qP2sVDNrejmWICXQ0wpB0Phhtpm4XZD3AguZ5d3njvaftMVkFmWe/b8YJhRIgij
VZiJnVkbMXwNJOLpKZxmryOuQaRHw2NpT6brlCw9jD1Sc6KrYT3v9fZMZ47TOEHg0ddxp+yUh2Y0
WUn1BZIIR3FqNrXcLeDuNR1V8uTvsJsxh41h/CEVxvcw1GufSkFf4OGxldsstOOb/N5VRrODBi68
HPO45sP38mW87Kfl1H3FtttwI5P6GOofW3ukxp/a/csWwBG+OeO9asQUAmEEZ0astQjKMlTPMYyY
LugcyUVYRrExD+Eeozxq2pnbwoY0bMOjEq2MGkU+dtIvaxhtNx33UUGHY8X49qqXqUNdNv1sRxUF
uq6bb3TMDo4ZxyQcI+FH0WdI4Ht6G5PdgoEw6IjvhO4rolYhwfWs6oJcKLFjH3Dzm3vHjVJN3QJ9
rEMD1HhIqhHKrTr3MxBBvof4HmtNOOiqoWZ2/cBiPNWToEaexnJPJ8ONsTCVaOyTrxl5QZYZqeUa
WafWPiyGoImgSIDgdJabtJn0UW9x2qAQKuEYexJl7wflaw4EoNr0Dp1vFX7dgc7Pkt12+0ba2QsL
fGNCJtIprlgnqw0z8n1BsveiePW9eo7X5ZvnC15xD9VhsBh/o30aaf9Fx91x0ZJ2TLlETHPh+1fk
i2o57TsDXceg8yv5aBneI/nBmX4DNjZmzaJL+yH87xcAACveZpZLqdvk7b6UEKYOj/7k9P89aLdM
/5qxA3bHu4Evlks6peR2sB38Uob5oqeyoGQgU6GXOSP0Im/iWmlDUSxcGrilRueEUBuaaVKve6Ue
oZSh9B43B9KxchHylYcMJDzL+CKusV3Ta0PRL3w06Fr17wQVJFd/WaKtz2wvQ7pfhCeg6Q4utqaS
U/cpLL6Czu073sODUDsG/2l/uSJdNWa0BEQKq3BX19waMZambXHqrsld5M/JqdN5SeShadCD4LBz
cLmZFlDGZJ50Z8tN2iyVKYW4Ekd+5krNt/6JcXtJSWdkHhmLakYD0gI+Yh1iTBv6XcFyhHOqcO62
NpUxFc0ZG383dX/XwgEaQVJJ37EwczlPetyqneBX+SeFLVVVYQ4zpHHheTxaZmrElZjwjoK0FhiS
QPnrlZVzUOtw6IIhLLHiHfgz1f9xrbE/64GDwIuXsF5ztf3tyNYYkukyvPkae/5GZ49Q99jLQRJC
R+uvCmR+N65kIqGOJ6BwbwE8b9BEcnfqo2GZRELVAZaoot916A3Dc+jEXCig7D/s7B7+njzn6Atd
vEiCRiwgE683J0eloE1BYNr+w8C8xourl239njGYACaRiVXVV0vU4geFgLpatJPeau4VdWGiEoJ6
B+aMXi52DEIGbwryB24Whc4Z/gb4SqnxRPYC8c8uHhSqLJdkRK9dvucEDTvc2/d1OQDwllWHmcNH
Z9MjaYU4MaXjfgOzBkHXMPgTRVvTTaHdLckiO4G3WvqG/cGvZCpPyzush5BgDQaRtrwpXvHKwsrX
SBmrW0DD0Dp3+1nm3o+1Ffh5lntNWPmBZ/QQse3H9k3lIMRrIL7+VTVJfV8RZlOVhSsMD084a/8l
GeZ+45JHS53XhPSV9MnbcFxRfnhUInxvzBQzmmAvxALt7PuELXTgNKtmYlpRwSqCiymNdnAjAl6o
y8OqvbYnsXWI40OkqKjis+M=
`protect end_protected

