

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
dwCKj5yWv0+IePBqJHT08eVU+DwkTeU5oOrKTCm5D5dLE5fjKonyT8s7ehOuYqmaU7hbrj8cK+dG
v6Hkf9vaEw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ofPimz6qWDPfdZmLTvO15AJD3qAYPdAcnxW7u3A5HKCVeJi1plo2JwW0CBkFgjSMPqG4mB4Hkwjh
aser6hfQcfNXvJ3JUWr5ZS6ezr5tSrAVnAOcpabYJ2vlFEce3rPTiHxnx3vwSLvA9frZJO+K8rqA
zTaVjBo7aLNhP54LcX8=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
xVx1mMvfUwlXTa88EF8IX42tnG0cXSGFt8ROQqT5GxjYzkciIVjF2lg5N/iujDWrU+m+Hq1jVN/S
7L9ZrnRgKz1GFQOxHGVlrNSRcf8Ej88lKuK02N1SzF4b1/VUH6ht92N2p/ROW4dBYnWVBpIxhF08
xg1QHd1cs9lodA6VBrB5Eo1G6aluz2m9EBGHigHdWN9RnmtH4Lso1/y7QElbZq3E4/diAxIYh9aF
1JcFvli+iX9S3ENdEluRyVweVryo5jTYqJabkRWFuo9iOs/Ic616lgSVONZ4NUl4ItIqkTq/gP0J
z13d7iJ5zyP7sku49PKKDfaHMGhWx7ug9eg68A==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
mm3ysnbGmWPGigjf3cW3nqCJ7td02DMWAwGM3y8Ir0JjWwms2hUSloczYrXXwus0KFJrOvbcp8EI
afa1rxF5AlIKiPd5moyH7qLa6s40f+FTseHQnAhUIfuaGWVSTafXnP1rMlydXotX0OgXaf8ss8Rn
aesy7+qw+4loCzosrzM=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
quGvQtw6SKSqCyA6Sp/eeM9Ow8TS12WLAPu5jebLdqM/ryW0A17A8N0thkaJZco15r7Owh4nFU5l
KZcrcDhvn1UKmGv+3eWd84UW4QDpY80dJTTq1XGSt54iFPTL0Mo21C1hbrKXm36H71Xi6xWsaAlk
nLsOCKMEHsujeF1naPb1xFZWSlnfCp9K2SB7wEzz8xUdktOS4rqm8CvHN3HMePG4N3SsN68l6nRq
sed/9GKEvYzA04tbQb5NASiphn6udoZq4W1cZDMS1xzdJ8v00rtDdh9Iinn05spY0CrdzbMqalEN
NkRAqp28PSG9/FiSfEP/QtuVq+XzCkevSe/NZA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 83872)
`protect data_block
Ml2+bwX28Emtq7Posn+A2rezU+/S9rXmBJ5CYmzgUChXySWt6K8uQfWpdEMe1vAZoj+pwuF/y/mr
TAKlEjyy/HiW+ta2KBgJCckHdHMRWKUaHnq20uIhnFaTVPe9CyRQUUCpBo/7DOcKJ5hCVEFwk2bz
rjPpHbCgcCddJEVeO7okeCHM2GuqDvQjT1lxdxZsn3jreg60O37GT05dRxnJj7V9Yc0Eu0LhP7S9
LjcP/nYB4iCvPcJ+8DjtK50FxlE+c8lxPTnxXAu5l2/AXWwXWG/uippwSQ6A2uGZkjt3Cjtcp3XE
jJPA+YhvarqxbKQrSycIQo+M6mCny4eiehS6zZ+gzFKeJPQfnKMALXZ5rpxEEDseId00K06yP1ah
TGEr54RX9WYvUAQFuz+ShR0H+keqDNWD+Gm9JYjrQqbTkdqXePao8rYFLW7RuRyjqkV0oeTeHhEj
POBBxv7reY92MKHJzwLEdgkoeBk85RIY/UK41ytAqqnL7iT+RXluMj7/air/e8g4LQIREYJM2aOD
Nc779D6bV/6XYVDqa19Xx6YOTWc0NLzhD4vgjlG10oru5AGxnwDijMsmVBwze8BCW7ZRUDOiuwPN
DsCuAomrN90IyWDUgQZxINgO5r0Ss5Oi7Tl8uFDDsV4A3su+nIg71GO3inDGkytd/ITN6eo2ip2k
mWs5hFkTkEmCy4I3TMSM3jo83bbYw4HH2Pn4F+3eMoMXVHbxKz62yD39r44p4rrs8IxU+M6akFVI
hTo+TZK8/Zr7ioXIC+6yz5IKENou428I0RwnDXVa3oDPrXjI26eLLQXenyzHvl0y7qMSNJQdBtlb
J2y/sR2H4Vh3y0PbTJG/Gx60HuPh+333HfopvQJzqdLajeCLI3dHytBsaYw/lvT1ErLHDSsFBH10
HTCWQ+Z/JwCrOMkb+uEksGlo/1apH5u3hRvIjHbJcl6VxlPDTVpjbzl1Sjv3sFx5WblKiwYg7X51
OSg55TJX4IO0CphbqMr7z9NkWpFFqBWTSVUNuyGVrvYAQsO4RROK8AK4kHJJSNk83ad29BrgbXtY
rLiva1PW8lVGQrJPx1cN9chQcT3DdhS58d5MsBRZMPdFbwJtxWCfpWIMfdJRQOO4tXwSrFH75mn7
yJXddt60kw3iFmNWmJB5KIt+7qDMk4+5UdxhszMzXxBV5rU8LNtot2bp49qf9a7Kfd7QIUbHStV3
RUCehoYn7DtCfsHPOzKffeAN3S6Vr7svy3BM9xUmg5dU5ZO0LdAl3eOvhDtuF1doL89pxhQGr2IS
Pe5tGrgcIuV+kVgZ9lNXeMclEIHmVZdsD5EDsooEFxuRlR0v0YKlyFx2dStNgsVXq/Wg9K+FTPQU
VmzEqJcbBFIo8j4Y3C2m0MgQlGa05YMbef860V1SoDUM0ziPFi9KbMO6UuiHbVVAmYe8QPEbCYpY
dSXva0EYClK/Q3mPK89XJn8NkvdRtw0kc45utq/0zswKnORPcSpLyMceHrZF6EffKLwv8ugUuwXH
+CafLR+k2jrn6RhUNi6vn64odRIdSaqDv0l5+PP4mbUTAOKPDBUV9Q0Eu/KlXC0VwkOmfuLoGpSN
NCi+ZEwu31Ag8aMduwOpCd1jkUobIXP9Ui+d45WfUp2aBVJXxod87C0BXf2B5xAl/MKdqTk/U67y
SgIaK5aN6VOA0qxOzP+WuSqEt/j36BvQyHASmW5N3Pwebx4LBaRUP83wLBY3xoRdmVOqd2x4t2Gf
f+LdBoB/Izw+wU9jmkfht4d6AkmXW8LPGb7nuWQ78CrBN1triSkS0YBITNMK5k7zBG0OiEP7ey09
PyFM/8HinvMgCNpBSxtn0c/bH/bQQX3VIDU33dFoCTUiYtCZ+/76RCB9eJYUnvslx0tLDKYInYEW
LSlXbUPPZQP0vjsQVP0FVFkkfpGUu/o5llkPw9UpKX9sN/rzc07JPTwkmUckuuenOXARiGUPo6/a
KmGg4dYxIRREPLvSIad181U8QBotBnddEGbbKid0VSG6uyNpQWdQm4aNJIXnG1XoaRXASCRW9mT+
FgqgOfNFZHVeHLM0ya8bf4HofM+GPmOWbFuR9tNyzS27KnhWtYR0jep7hun+mFuJgK27d13JJZp8
9lShfrYknOVP05pfGaFXIHiBXN6xW4sFkHxe30jUT4uIOK5rh7q9XgPnMFv59Riv7l+RJoUHxugR
fDpQ6PPutTGsmKHHqqohUQoMdx/UBapIbeZxjB9Z4PwPRvHdzm3Sa8HEUGewrivUseTFvykjJqnn
DUD/4Ih6r/L1EVewr7942AfRVcMn0ZZYQ6toxiEs6SqppoAMSWsnRvmgq0L5RJZfpzRI40IfiXko
Qrgv31WIkzhPIOxIXY6v7BFP9pnJWbnclgNl5BDWM70hXy8+4xvcPtVrHNjZFG19Cvj4Fne8CU1h
9Je8k0DxDXBPy8UHzXOBOqTmITtOU5BteZEYpR3/PiXiW3dKjoofzNd1IOrJPKb82DBL/t7Nvg7L
nNv4ZyU8eSDpetT5npzJepA0miFskQ0YsFTOn8fH2VrAJLqF5kO14KTKolYujzpIQoikBzYt5ahC
zkcAZllwfW3WWTJnXGaJtLFdevRJMk1Qbbr7KQLlbSQlK3SVXCa3RhHJYfgRD1Vnnl18uW9HZ6f/
j8bmO7sT0wL2ldaWoS8URFjPv8NGzQ/BOVdbxUKc341TwuOJ6hyP1CjC4OInZosSbF+QGadORhYw
IA69/N1sIUCyprKPScb0jFq/QtQ+f5u9CZwd/3HFEZULcxnnMAvL3wOBNMGLwWf7hP1xrjpd3zLi
biJDwjUK1fj9nhWUzFj0PK3OiTyqXkvwLLVZuiqXi9niGKatdllQ7wn1ZZhCeCaH1uHoGW9aLACv
8zROMV64llvfP00NlC+3dMyl6WnpvHmB7W+aANL32tm6xZok0YP37+Mtiimy9S6WiaiqJfeJ8hs1
WPpo7bMDTo0gfuqBGNWF4TFHsUkV32sO+klK1DKtO8mBgTERz2uKDzeOKbpMMZ3UQVzvjRw4ZSLG
h+trDOJ7BSMKzdYUy8IhYDDotoveJRSzrHs9ZB0P75Eayx0Q5M9oULqnXP+wi/deYbsmkANeUcpP
/l5gCwGz67qpsPiQsSMg8iPn2UiUDBb5ZqVx+Le+6R4WtzzWS/Jl9iOmktRhY/IpMTk0ROQ3KoMS
Y+piGEbe2RB6qLKYkeDLVM0oHv5e3OnxlVuHjdkJqj6TiCSkIbBBe1Cx9SPeIkUuFKnJdJSf7OxS
m7YJ+e9eCpOX1kiMyG7ZBL11nFFeTUTRgxid7sI8oE+V0kaSUOtzl2Q2jbxVWNvzhrKlaUW7XkQJ
QMt2VfgCvp9TG32uisfGVKmD89Phh1Tu1wctpPp4jQKzP1NlTGlte4M47ns6vJcyWL6WrvFLeYK2
KaO5828m0WPqVznLirUUx/2W2TXV2UL4/EJIZIbnpokr5g5GoSAoQ9yZM1z1m/Jqkge4erzTGXEU
QFmvnMjZJlq9nVuG5gb9GwhA2XOa05IN4F7Lwy3+ve8MNYLwMMzNeZN/gGhVng7SiCQwa5KK8Q6j
hyAb5kKJbqPaFUQvEU5TERo2GOIqUaLLOEW3j8c2s43dgwsh0K1DCS9SdBZipB9MnsepFDuvarbH
x4QkLXBUertMaSot8i9H9YNkwasrnp9RapEyXy576usQspOdMZYmbr6LeOqVaYvutxVye1HiNPCT
hBX2n9pzGnuyuv8sBbQsrZ0FPwtVRYV5gGgF9oLwnopETLsYZZK2NA/y07vSgShNL06RWxlrlSpf
TQhNrF4M9FGjHnDgq9cyAxcdxALB8pCu1y7KV8Nrtoblb5mZ/0Zs0/ZQTvJQB7Hs1OtGoqQBW4Ul
8DlxnW28I26w7nt0aTbteyUZsp6VQUV9uUeBGNSuchTO9Ko+XhN4gZUkbFNaVZ8qTwuEdKlYgjps
w3jqeDzX71lvSh0Y/s0haIMP6PX93tN/WUoh29KDEfQE+5pAo4jvlP08VtzTBqPBMzlMKJ6+xJoV
pdSr/0akDfvGVHEf0SodaEqs91WrYjxpiqenh0HX//UrIGXeh9tzEhzCwwzCMoYnD0VLaKxv6d9Q
yBKSvB+3Nqqz3I3y+etIDkAXrZtVkyNRqT3/wIc0Ket9DLiL2vYPiKdh2UgzfT0EbAG/Q+ObSvtQ
sFQSCGOSqD/HxLqlXqyZHQLO1cs+UrrFQQEqy8Mg1maSRKv/PTd+PPgW089WsZnWXvd283MQhpag
W3Qtr05sjI/iU7Nou9R9epKU4AEFwXClNj8ogVstIJFxd3iad2W8ECBy2Qy/cdfAi/gkXJdV1cwz
/d27Z9QGbMtSkmDIJsLJCO5uRsEH1P3OcG/pVZDWkpKVfq8GYXWkv48OLAKYU+amA65JxQL33GuG
7iVN8qW/JJhiZ3MXBgeDFNEQ5LszULosMTppf50yyin244I6CBMWcqohdp9pv9xcE97R+tYilboo
um4+mFWES40WoY3IrHxA6hnuVRtuVFQFpTAljfIj3FqXIJDi2dEu7C2chZSJn0UXKfK/evx+NnAL
tFuH02e3xUdQ3iCGmzaJZS6IsBb74ovmgBI8gqrh25LZwEVreB7utXnaVd2I2QKzpBvFDdAiwi3U
vA2KxHetnrPS0eNFOsNK4gLhJ7Zr3QAGYrSq4HhrdY9/SEmXWNbTVbiLNeyM58CgohxSJJy8Z6SA
ROuAPzM3LTxlQypJFCZEpnX4i/uY3wsocSeDU0PAMai672mIFE/0/J3TONkU4TA40k7h69CyYAqn
8tr2pDGKeeg4pljujCEY7eSujoRUTgTjrIeW52xb0Ul93fntu7DORgWBiwD0Lp5jEdSbX2IEs160
nOlhRtx4K9NcsMXprucXYwm/6Sb3MyfzT06riGf/PKdKwaqKmvb9gwcEnxJCP6IacwzNJQy2OHJO
csXG/s1Qe8T6nqVqn3aMJIFD3KveCPGHIahrxzbQ447bqhwQnMWeoWrNtfqmSdfOulF8p+6Msm5T
ubHZ+Xq53EY2oidKBUDY8wrmV1AEHZks7zAgznjMbHcIfHbJm0fYiTQ5m1hEVBxlYy3FXKDkyEZp
BVfTGufcHxF5GCqvJJi7xvtKBMaarFpD/AupHQ1+raEOWzXfiAWEo3/G09rm+QnXXfNttjWAy3xS
XZd+wck7sHUgS+0yAq36wHiK8dDYRrsq3iW7JKxS0w5CdnnpDZut4lb0uMDVzzdeZ6HzxIxwMLWv
9jq0n+fu8RhHZOrHx81ZvUZ2j+Q22989R/GkZJuRpYC1nNh6/BP6e6owYMw2YWbswqQlrL97MbJc
OgpuvTxuRDOaCW5fCj2pKLJiDLZExVpSwcBzwTtS+lxYXDxoebJiV18Gok86Xaxjm2lCgfo02wZP
qRHHQnokM7tXcQLxIo89L/louYzjN01XsP7BqcKyqNjkmZGp2LcEQ0osagWT6rQ7EgxQSqbkSVXM
b2sxD1bEnyhEMQF9DRktfEadenSZSwnxwLM3rFhv5gbB3m9LpZIRlDbkhL+3cPzn+P0OJVbEM3i3
HmXrH2pwjaqlQ0/5vwkX6cxOM+jmHCfNtEwa29T5xfQkhpR86FhXCuIyXRj0dt5aWuuRcKlZOFup
kswsdsaTx5NspY1LvdFhR5SfC3xaY2kUUq2fzfFjtvVG758gmLyZ3rCnHK0OWVcpklmNfHX9RLi8
Y74B1HNj1pJ7UyVke7h/nHu3Mb9zb3tR5Rk125Hf13uGZj1qnWL2KrHCp6EntKC426kUXDSfVTBX
DzBanzPWYQJ/h4RfDizDun0X1A6ZsrubyW4zRDl1IhAPxUbaOYtBupMtVVFoMUxN0eXfAH5huhpi
8ZYlpFkh3NT083AUy3BbLH+zsMVcH1Rv/mEYz2itUr22UcZQcFd2v/bMOi30NpruKrEX7cET2Nxv
ROFh0tQFsKlKjFy/gDs7g7II2kfzp0If735tI3ZCgGnuxd09x68VC5T2JwAsWYmxvI4HVjnz7i1D
VW0KHrCmUwbHl2izZxrWSYHsGSaNe55wz224jg0wZ6FKwDyY6s3hoE82umKybUMWAbPsznFw28+c
+cwnp2WEIDyI5dfAh7PHGfEak2lQsyQrd5Ijgv46F0In1482XZlRtQOfV7q98a7JA9yIIYzP8Sey
UeludgdnkpEMiVXRjuQomub6hlo4gOBBuOXrv2BhBUyxD5DB3sJtNYYFnKuF5jh1Ty3LraRHQ4Kv
AhzJZsPZkerRVcSlMCVDUrIKGnXFWb2r+Tl+HmZ8jG7qvJEFjuNxnNWUO4p9VV0EKdU/yqLH8l5e
pe+FtcfoxZxV2yiSogWkLB+REqNe2jeIlr5LVxHaogBy5n5p9ycIO5rdb0idusUae6xhDYxMm0RJ
NUwgV8I6thnOTGUb8A1KqVsOzIvSPWefO1xSMu87qbOH+PQb6+09ibTk8O8Adx/HDx1HMreD9HZX
kP7RydwaWRaJgXm2BgHtUR/ohzaDKoQ+4cXuNgl0HAVbMvF5S70XYmYRWPvPVtWENX+ACtncAx0J
zqLLXE7jgQO0TA1ah6Msz+FJJc2Uk1dY0ocqeFaRvQFeeA2tINYtKmBtq7pEZM0Y02+61KmBgpKG
vw23jHip51c04+Lvoi8ZtLyH4wTxFrQZNOGCEnd0BBI5AtdJ5UklT75mU619lIHqN2Y07N8egygt
+b0ePMnUlrDmz0mpN6kY/8dtT4I993ruhiZ4lJoMFKJZT5mYcPxCg5JD3TPRc2sRoodhN+9IdtFY
YI1DIHvftKmhcSBa8+S5H3ahINV+5HsqDlskYvSQgR/5P/YQiP7sm52MbVTytggCOel/hR6m9aqU
mMqEsOEfE1/j4uFXqBFoeLTHj3z08LxvSW6HjlGOTGbbwnC6Ti2FdW7GTFKJdYBrp3N4vOZTw2XG
rgh8Us4UUsOs84XTAmwrqlK47jYrjm55kEKX7bu601pDng2xmSD7tnOzk9eUUBnESiFJuMRxyPq3
NWZ/kvfIwcpvSIlR7BLTd5x450Qg/aUCJNXZfTtMeC/fcy0gIpuzdbCgWBVRDKskSAY4s8dP/Vwn
bRSfPspmy4n2DuJVHRv4F22nQmxk+wClrdGvjUCTSpYHROg/NuyKo4q+hLhaUkAskFvQ82yGpvY6
WjSz1v+UvOHKzQIGVAs/iGp18R5y1kZcdIZdbLsaF3/WZz3TieXsjCqY8dDYipB8JGpnHguQ1Vvx
1UATMOr27dElmpgDAO7p/qcWebsy3+wi/PqzoDnd8i3CtQHN2ssktLbGzvPxnKNtFZjbMmoIyrgP
PP9gS8FMU66A74kJJaekNgnnoEF3hE3zHut4qAt93tTA3ilfbV3WzEL2eqrwy1oWtlsm35W+bBf/
ElxN1iUotWwe1JmfWSxjij5NHhg0TBp7HFXPmD82/FES7dYiojIIcD6mEKUGIddH0vgGRQHhAR9e
7hXz1VjDBYmG1liFm17JdjD2SpainKr0PPcCsbberzPZqwiRHbLgiZ+0z/TAw6eD9gABBULSlvOa
AF5IC5Ay0WwXdvuOXCMgSNVfSDCQFHTfejHAhsX30HOwdrvvmu8tyxvEeXntsZj+ivggL/z2xxdF
fB1mVpbPUWIGC8Ts6BNhkmqAKtLpqssN3U0kFhO6lsMvnL0Sx/1Lv0CW5X2Y+0EYnkaBRxE9wCHB
NLNl+A+8lWMlWk1S/HXhMhZHZGjt+Os8zIW7w1zxQJx/8mL6XSEJdKH/TZ7zaKaBk5zhvNN6zNHj
ZvNpzJSnSJ1LAyc8Dydr2YDrxtzTpX1ZO/4wd7H9NSCoPGznYdOpQjMswOpmOY9BFfaVzm9sBm+M
vA+qhjXXETDYpQzNzvdZd5GpL+ZnJQqfz3UOx2RQ5GvEsuOh8kxkv7saClz7hPqJhmngyUr1JuBp
nX0dFFH19KT7blOgBNv3xXWF0jwOS8GhxfZ0nm7rl4a6f8FdzbZZSP2CbvyNp2ExBHkznLopwkCM
Qfbv+ADPABiqFcgM28bzJM3kTbqhZGRAX9STG5j2uYtpCZGRCxHIMcUei6Kv27LLX6GBGtyd3nkd
KYUUVS2OsOCAP00pTf2LT5H+WQ8KfoFWtk//94ApLsO2fIvg9+azktrFJn7SO8Om8S2+bz/Dxcmv
r8bCZ9ZJATj5Uq2ZU4uBwNBItGRZIvzZ3O2l9JuiPXSFi7dlrrET4X0n/8bCkk5LPMYx/aQSVVsv
tI/9J7X3Abb1/e5d9KRZ+xgBDukgSBLwfFkxsdsDpZbdC7MFqak97MOSW9nAatqi/CYDNnoXqpjT
tSS4G43FEQ7ykKomvqQwl7zOmTBdWUX/Qntki+TBtUK9iSNaMAB6UAshAs+yrkBg0iYaCO7v3/BT
g6XkkCvHIPTfHTA8BcQhJ19vSGpBAC8zO4ScaG/lyZuK/OaT7Q2EGYaSn2whipcwR46KPavxWZYA
mUQIde+zwTV/iumFYVATKwMWROyI+LxFgR5f9dfYZJRuD34braCRx5YpMZBhl3juYmxjq3XV7Htt
O686vxd7ORct1EGrNp66IZMRcNjCDwv2/zKVFppv9DhAz4TdBWVwW0fe2P4yJCq/hdfz5wJPtRdx
bShpbsPynpWtstkMWmqxn46ysDJReWEIyYzSBTVwWRZjYiPEcbbRq5JLFnXFGLx6pVIRkXS21Ni2
GiQOZWpTtrZ5wkTLhDt56IMFKLcD5neeID29VNsszEnKgq5MGM2+Yr1hda1C9HvLNx+cWTA5FIFm
O85Y1eHvkMBjXd9w+0zKJinmOcqK+P509RXOytcvOFAPht0zBnufNxQtSPXsv55DBUdilK3xDtR+
spbwLSBZF5EVu40SF8rEeB/Pa8FXUiqkyhuNFjYuKjLX3o7N/FCwhNmxNuXGusq/dwxg8y0TcI4d
J4TudAcWu1Fl0mLAQ3g6MHH8vIlaQODhi/HV+ADIu0pn4qgJRU6kQQS1YJxCg5rlnYQCMWzbwd3W
o0eUNSZ9ibJNUomaraqpkeoCcIdyTBiOis0aCRx2BSceO7M6CvqzzRtAxhwc37K2kq6NFK3QbVwV
P+jNyFJOxRZh2gCrFYHAFuaVPdUq5drkK+FUgNTPYIxFpjaqsJxHg/0Ka5CSTh7RPDp/wGa3mmFj
iwMJnel/zQQyYJAJ9/Gd+emcZ8X2b4265nw84+hfx7zggKUOrbowxCZ5fcQSqCC22EF4orRPD2KV
Wcb15+yOQdYWk0xMygb6C//0vQVF639KJlqiPu/N+cfW2uJat+lvtWxqM4uTcIrwYNh7hPfu6H7P
IDchPDWTKRr6WjP8QuPFNZ7mcILWNMP0QGWM8lki3AuNLYEfpdkJRph4+oCj3rQofIoqKm1YygiQ
LWPQ+ohF/YuqolPd0b8oVOeBO8TODHzcEpiYMyrlk3945PH0tMxXigVeWduKlPbnQv/9uVtraieT
i2V5AwGlCP9a4JuMPE1nJWMiQI33dp5N5Zx7ATNIh8PDvphw8UKUtXlYcW6+aNJgKttPkUg1+vQg
nTA9bcmhUNpAGvMz2FridH4/DpnKCANbmQa46c1NJiTVOlgfRk0LUb3Wrl4batjWxFlTfRfi6DHT
2lOkGYLi2uiBFJXdqsa1yNCQK7Ol4nhLKH89d1VxjPvLmOALIvddeaAKj2nQfFTLEksnzFekTBWi
Jonn0aYcnJSeTbAU8O+PZvR4Xt1vhdZqPeFQAInesDqDR6VvFQSBCi6eluda4W/4Qt4VPRtsJqqV
xsSylc+FnMSQUqtlW+0/V7szTfSDC+gRj/1Z20rr7dOLNrsn0aUolJdduDl28XnfS4ujKLeSQs4W
J+qf/ikgYbEKwtpGNDWzfK8sdJaLE9fCgtCE2GqHa7/PFDR0zub8fFNrOWX1vv64f6OqZSFb3wsV
lgNs1wtxg6GZLx/pPGl/RjQ1hIz70bNU+ILeYi2AzV7q/zls4Yhpd2o07S54iLzvLYHzJIfW9y93
pNMP/dcOkzs6DTwl+5/2xkMlk+CNsPuemEBJc6z2HQGp3PTbp0YFSuqjgYfO41EnIqhwJn5Qjvkq
aSIrPvOi5K9WJUFRXF4gaWfsX5dgiX4eMnz7VTNZYsfT02eVpNL4svdS3IqdsL8J84zkS5htJbsu
s6XBTWDWF1Hq9WceOW1xNxO4rxzkvdW+7Om42w4ZIrbRmStF9+gdrAFkH/A+WMiqxMUUxiOIad7L
zi73gAQaW8FgT82On96zBm/nnXEF4LSEj2EAqKlwOI0v4364ht4rhLwec+28LhpRS9wLF/oMhWFf
7/lI4we6clAIXM8pwgIErDU653d3gYeQysjHIm7JDEjlvMdPiC72plf9NL2D/Glu17V5FJovZkS4
jCaqo3qPr+SbtS7gh/qNHV4RfO4iyGDh5Vs1vkmgDZU/k9juoHToIR3ywXnICUt9CSIBdijkRhwY
KFaa6hj0Zaq3kxtGR13EFpH4gkPOaermaMQvwibyB4tLQzYQKllRA3g6fs9BhVB9AvsfwnM2Fu3e
CUCvkMxMRdIxpm79rvXF20WkeQj1i6YL/lRKI5f5VA/l1cE5kUkgLo05rCOvaILxwj9VCz8s8q4m
OaN8sA0UEQROmJIlhzxk1BKKGbTwpSn8If9ewZ+o+XPzaziraAB5CPi0K8w79fzYiohyUMRsrPdH
A+qHoecGM/efDzOmS8u25ZIhaN9W/UCZ4uCXnrmJrRi27qmOVBNL+IPtnmXI/UpOON8qwNA3x7Cl
R52qW+8HfZ38+1Z6prw2Dosgm/Q2h9C6PPcnwozS+ceHl54X3PW9F4Qx9NFPXgGt6BUD4uLC6fef
tumvZw7tW30lvuip3aa9Sq0al0yWtHUQ4ESsQ4Spmb3nDkwOnoep3zWu/RinDCSzR4+ZpzQ0oeC4
Vr/Nw7g7eUV2ABd88m+MTQNmj3zeWhi943NiuosMxvjUsHUKZHF8nfscvLYQZtw6yhUwkQLCCEoK
RQyXC4XBZR5Ltzfw73BvLNUmSSfpOK+fP3rScCwNDBcnqpAPwcOlaTOcMBYbTAFJsaiu851WsDkJ
wa7Yx3jhFQmxl9DqUulqLPgnSU9s4/5iZmGz8Q/jzk6uerjcUHH3inn6U6dMkPWuou7Zl+taevLI
DjbyTntXkWS37hCawFyT84KDhj2439V6VL6snKkyu03XGg4vZzKl0qtM3tyLnZnC3NYeXSQ5HZCC
WAt6nMuS8EvcU9LwcxaS53jEJN91JjFxun3IG8dZzNA5Bs7lI6GI/9eA4AAXmeYo9MOc4TGOck7A
293xQsKS+rWDL+zYCeInQv8A/hIEwEOPPtMOmXssbJyci8zrR6GSPOOelKVAuRAVNKOWc3r7ecLh
SBf93Z7Kh9aahPHGkOtlW12BX103wlfSDjl/1nf3c/vGjlYGoAV5c7bwHSxiDFqbiH4xFvOoNPKZ
xVuHQBt7zFruwiaOlocZl1WrleQz6JWD1a72Pk8l4h1dgj/PMVzjpNHPu6HX4/Af0UC+j6dN6Xyk
qkMM9qI4fKIvYS6BDBRBhnU6siZ2zHFrWfRQHaB4UfzvD3pi4qDwDdqoEBTjduoU6gbV7YQxbi9m
u/sp5K2MbOxySr5sDbdfdgxCuntCjWayIrEh9VMSWGoogE1GKKwXFAWgCl06rF5RDqx9+M0TfN3W
+W7WvZBTcgp8qmysTvX/dpbI9CIjyE+19WJ+hj4r35eKRrFp09Skjv8NRIRye4gBbu+bGP1r2X1a
QNVPwyNlHMshXbGSqcUyP4c3y3yBuCSTeuGkZQ3nehhR3EtPZJiCJT1891uWr/S7X8/Qy/aovm5j
c2VEZrZlCVqK/3LhqFO8igxsX/kWUht+aRdEMhpFyXtm677rkkDySPCrREx7FaVXkt+tvCviJp8r
BluEzH/0Ce8zhAHdnlFUGjCJsA0xcaF3ZFtiVCzrAEMQoAFLz1ekyTo7rm1EzYFPg6mMhVsVhi/d
CVM8dlhRsMbVHFxcbX9341Sj3dqCG8db/VOpgrvzDgmJea07ool80zc2E5cUudjYXiHGlyvYlDiq
j2Os/6j9PCQNIpuxUNKKjCBs/wHxDJQBeYp3Om5IRJHW2qdjESMdRlZh4FdyQm2iXe6ziVeNwcOg
QLBlX5BkLTDiGn983NCmQvL5z8cFjZj3pMQjcPKT+9bZLIFhY0YRtSlI6Lc31P11kz6MLbE5XFCQ
PSgmKKeTrPryRPR/wo90a+HcD/ew/btAkj9DwUdPd/xVKaRL3v+i6XB6rALTm0Ibx9DOx7B2ksHb
R9viODjG2Tvzl31zAvFjhEFZkPdO3HLMRamBzjnjMJ/M1I/6706XV4gAfMY5rbdulc9BBsyUYe7o
Aryej83bzbbQsiNpTlCy+sjzauXQSSQ3B952sgkYlftTegSMLSUgQ8SVYMbphkxp2flMbzccNQig
GLumUzTghqeJRMz8wfaHW76UNdrrkp9XCRPol7fH7tP2iBz1feGBgIlUJVkDhN1zJTWTWHUmjyMn
jOPUwvkHR1sTmLqjNbh81mXOz53pxD+rIjpzsInD7XDkrSE0EKe77rzQyWhHQ7dn5XXKSkXhHiuP
dfRicfn2FNfOYPHswyOBWZP+G9lydYLjRDlYOuoOZGrrI9ADzllnC4vUVwBl28y1aH5RqmqTvfIG
U7d8sQOGEAAFsfc/W8prQIcIHAxLBOzOXkkkIj5ERWAQS1FdBoRGwiI6ePhYXZ2ohCIGogrBhDsO
08OtUcuElxlmvz/6ZH27NnJ85wP/bciwbqiOKAdnD4v51IDZZhugskKGoP7dhg5waIhTo4D7ATD+
OMhuWi4ASMdD92tzShIn1TMgvOWYY5zEgmfbaMjkS4lQwQvZAytiE1uglOQ0429/9E3I9UJkNCqs
rdi94nddB4+rg4j98p+zeTq36r+wK9m24uIRmgRSWqoLtDgGTfVUCjq/yPaIbkEXOeLEc1ZbXSIm
NCvmyOZmdPvUfxs9QPkTdKvEaOzsxM7d25a4D4Ftn9xMrRESv93nMpB5CvXOb3dqYZwbMXwViW3h
cU7puQCZ0f2J4hk1rCiplwdwWOujav1jPwx+DgLljCl3oQ0s6/rcEHabXAT//77TCOoGcqREfeau
6usUEITDrP7HI+j42YYGqkxZwG9j4qC7vv7kHCzAmcFhsMnEuUnmfVYLl8MJy5WbdKagoV87gkgw
EoRKpqdwqM98A7Ulk0b1OjflPDyaUxRE5PYMAvm25i+6frEXNxz88qI+NQu/Ci4fUoaQODt8DYYT
hB9ykaxyXZEbuD0vMjEfqo6ypHHNOOvocAVMVuhz+pI/gGKOZUGFlQ/vbof06ZrPRjHheSWCI99C
F7/qm1mZfHRFaeJQA/RvbM+Zhc7uQx4HC2s/vNJdJ+mE7vHBUAqvda/nz770ZCrNh3ibBS6PU4ZE
DujuzMVG8pTR1018yvZW1hMA9EvANWnZfZbToluDzSbS0TZa5O2y5x3goED2os8/J4Ctv6075y+q
xys77vPiwfLan0QWlZT6z+rntkyL3HB+S46YcTYBT417GG3eITy8MczC8mfWqjncF49gP8dDmHNj
G4RFv9G3lUNwMfUqa3UCspzYyNtkjiZyQp0pje1jUKY8q0H79p6BRrpm38X7SWTb7IZjKe625+hu
u85cM3qMTkxyv+1hPYxPo2P2XutmbnYFR9gtL9ZE/Wg5w3zkhfAxe7jGFQoWbTYIzTXB/PDqhzxz
V2E8DKSul9HMO2hvU0UOAFeVmWzZXx0ghA69sKcvn2mgZf5mgW4g66GzstUNNdldAAkUYvZ70Sh8
f1Vm6jC/1PLVsPeaXPsiJknAJholsHfQ9QiHw2crl2xnWO6+YnGY/wc9RCEiT/X9NgsrJQJSre5T
Pmm0AxVQWEuxfMhMNUF/Zx8rAarVT1lEvqreJbe1+6cE4r3jjtq1n4XOilBzxtAO/NXVhXwp/Ysn
vMdVQ85qDoZuv1vV9ROaZq8slM/TrsD/cnf/588L30nB4Ah6JXVbPdqako6lIyDVH91C7SPX6Lz/
voXG5TlUfcWMGRCpiF3/UE1rT0DW9ihAhjwHkNr1KRCotanyOPhcU7vKdK5CK6qccx5MC6BVpJl1
OKpnUhEhqWMmMnIp3Ty2+7l8frc3Orf3+4meUiwbXRVwcigoVmnBPMPhvWlDBnbICnweGM5WUNoF
H8wlvzFb68CBG9i4ZMzhDW5HaWWU2bBqFHMFo+Bf1yb7pfsXoB7MK/AAqNzscuuJ4ITdpaLNTHQ6
+LiL3YuieWs/VR8m9Slc2P9wx8mIKK7YAQeehXLZbZfUJs+3ATzmjMr0BRo0QezxRJbvb8IlBQu5
wULsEgjo8Dnzj/zHWW+aJtbrdVpLLY14XohZuFo5+GFMcLI/eGWZu62YfSLz/YuPYji475bGMVmd
QZL0MPdE8TK/VO7KdBpo8OOXXQ3Ii8ku+ICDQBpLL0Cj+96B1WXkWsPsCZ2E7qRDVBnBeMDVHTl+
ydnVEGQEcjGXDfZAP6qbRNCwX3+4Uw2Lc7TlX8AlHZLa9ZXcKiTC7RQeGtv/2EzTzFyUYd0qpSH6
Q1ec0PP48oke9e3Mlb36za5C8RMYmgI9S7TkSH6m0bWLxUqUXdin4SkSJA6q0b2fhdgzeo9HjRVi
nUaoLb497RmVinGOhj8DJsx+vnGVEu2dbt2fAbQxir9cA+tJBjxpF6VT3fphVs8oum3pAkAHzLLf
g8oqFZdV0+RfgFs59I+YOEzkODMLXcDJMxucvd0I+JzaJCstqIBhoa9ONSUlx/P26k28NY4Uxe6x
ytmqpufkQ75er0MqztszSNYeCeUtWfjR6OOO/gEE26PiB0meMEojZvRtfbdJwZVzujbW7Nen/B61
j7X2yWFhy7u3aYSv35IinOLiKl+Tfc+ommfRA6hXP/m8KugqYGNzArdwmkA77RVC3jYYSKLViiJR
OXaRFBW7iqsreCW0EnSpRFiZdyp/cVdA9igh/OL5NMrwN1QmIFmp8PEYwOD11NG8zJMHVkxj9crW
8UNozXmkyegQEoADV9weDo+0esPvUEg+0S9WBKVcKcANC98OWMqJPGI8bi6p+QmkGwd2BmRhTvbQ
ll5af6XQ+FkK8EMTXfVh0dcR+LrNf/ZpIGEjC03nEJ9L40KaD0rjS/F5rsBTwUPpolndmg8449Ot
SRZKt/RtCGjP5JbIuBHDRnjmrS+clEyK5frpSscLBaJ9XOOpiFSC5B0KQeeHPPbL8FH21MZR+CIt
iwi4kDA0UX37J16YHw1uQtHVlV5bE90Qry+Bwd1eE0H+T2J5MnY40bKiHH/m0FQPwaNdQ84OLK0r
hjaCrWzH0BVWeiUXtA+Qxgk5PeMJji11WYFc1xQzzljUAAVVSGDoC8yY3Yxn5t1ACB5SPX3msiUJ
v0WrDPMSNghI85P4Oc1JtoCIO/zJLI80uiiwN83/V/tHHFfvtz/5mrxD1LgOohLiqtaPZIQ1UGsD
tSiI6Yzsh6sDaD7Dr32seSHhpczmA1zlu8nDBZgZVET14wucnTzKNoOdOdaG6ejH21O/6aKfQNTY
wyPW4y7GORN84kS6ZHuiTi7k3WjCLqagYe+C5AUjAzzx2BsLl/55kBkm72I0/XaIKkkDuoneru7V
8aXmIfDZhmJyKsFqrLQMfOrGYKttmBXFSv8polYU58JGJl3OSSA9TcZ7r0o/aXy+HKh0CUkmT2Ao
EgDk6/BLgLGTrurDfatN5Ly13h3GmfBkp7DBz6KNv887QXsBSbtqCIaRj+Trvq4m9p86Vj4mZE2Q
nv3mIyrW0sSnsn8dyLxO3wvjFqtdG4gPthwESPbf1xCKz/ApOG3YNZCnUMiosU2BjsVl8bVbjVYM
hTlwIer5aZNapDa3OsQ49Uu0UGqn5iMEMjTZaq1hcQckTkbnPpzUTFTzXpZaD07GEWcCbvvbRsAU
NtBkVtbfu1YNf0wMqabmOpalsjI1Qftd4AUVfrQGXnDEHg9f65gBNCrFVX10aqvy9Wmj5x7hkVq9
3xIcIdTvEF2LdutTAAiY/Olh53GpTpj4CdZIuxcsTN8IwF/FFMLwGyn7lRn/G4KuuMmP/3WWFSfz
GKjpOWk/gtryNU8i+dGoJ+NlHSOw5M63BH9XJHLwiNtNhQDr0MNhHJtj2GNErN/6lA/qLaM3zLYE
rXh9S4ip6rASrjtqxr5OuA7fm0kS8/cDREAvHtE9JmW3W+AQCBzwBSFx9LIaAyY2sMYEPH2jaM+f
16irpguipxLrqWk4PlwZkmP/p5r+sltDdhu7ACt+ZGGGEZE7xV6GrK+n96m/99jP4YuRRRLdVCPR
kz+gSKQQOBiuHF4M7UYK5HBUhl83sL3O6MTRjSaw+Grfmi/yovQVf7+wq4RMjgRs6SGdUaoKwrkT
0vxVWXfE+/5fMQGY35K2xkLaOYS3S5nXee3VWCq81ETyHSO7s6hhYTsyjhd6iRbweUmPY+sILviM
9XWsTnz7EcRp5ATUi1PXRQUFTjAXE88mFt9mKmqfAnRw1c+TgBwxXPftSHFvXGZk/b7kuRZubmUU
5tMIL6a7Bh24BKFfFZTbI77yTbEEjiBeq8nShI4P475cAK2hIS2n9yUpUqs3awQvC5ObXSwE93MB
OJXl5yWWPyyTWEknN3oTV0kbpulUf5l2kJ88iMrcPN5CHVdblla+7fFmgFT/hgOX5z7cra09AjD/
5tcOMOUJTJOx0WLEK6b7Xzy09LCbAoxcPTGmi8dpJKgTd5RAfgusxCfehc2lkF2mOFqCXHotjhyP
oQNb8ciy+VL6Wo9nklA1s3PzJk205fWMnGHE66EgJhj30z+j+UxCEq5nwN6vJwQGbUDLvb83X+eN
/JzBQKyKmc/JrzGotFf4DkHzFMTS2QI95ZgywtAxnOXACMI5Nqye9PFH6mEMpKXokotXpySD1c04
4T0vo4QehzNVaIfrCctQvigQLi7P2nETf3bWmRvz6IlYonT7rWxODnfK/mtnUQOQ6aUIBRR25Wis
3wPvtFTcC/VWRboMDVT7uSQBObrBGQ/EN44APkpe2hYbpVyL21Yg5IDyjo2CbUmo3B4uaGHaFXlH
Q8DFu1BbUZUtF0bRCF7SYU/rH3O+ruyVDNzm1B3st9069QDV0Ila9mTbyu9//HwJot2sfzkVodcb
vj6r6A5ZAZQf9PaPqAyAo4PCHWPFYEX9GY+gPg++KzsW5GC8wO3t/C0bAXkTQxyEioHz9GPGj3r4
7EQDfAJ/GLHrGvHtm74V8eI3SLfjuLqosDS8fHS3TXYNycs6+JeUe6LJyG2K2cG55QaGoHuQ/KSc
Jw+Z/lF1YJghJd+eH11hH6TIwEHl1/nyHTRnBNP2Dn6hd8C9eCPGUeWFi1YGZp0nLrz8+kRWgT/g
zRP5sf1piofFQNkefVKQK951CY9c7dvBtDEnrefDhT4TL4y2fhhqhxdxJp4NRLl76J74/a5a6eA6
oRhXgbkVKFdC17sD4pr7B/BuH+LjEsvy7gWPG/iQTR7avhhFT9GDinRz3r8UBQH/mujV2m2ucPv/
pNBZIc2+8Nic8hATCTIpWinvfvbHeg+dtAN6hwBak/0okF/Oyjqg9qF3MUsgHqO9qXeUvqja1Cel
NsQiiPX3U3jF+LfSlK+HrPsBgQ14Cej6BkfM9nh3kH1R5ZLMOub3fwmzMkjSXkz05SLRjSXtrlTH
sZj6qaLb86rNaZqQnkjMyenPfXSvP/9459DGMxkrCd0PFD49lXBw63Bhj7EbNynK48Fnhom79kDA
sdvNFH7oZ0L2wt2/V20I61BJeMczMjGQNtzlyGkSlH3s3Uqf56Fd4JK6LLpsmUepvVg/HaZ9v7xq
fDWigUsINiBXVZM+N5pDoSCS4c1tx54U3YLVd35RNv0OYEHo1DSyc5gNmZoG1PfuqD6JSKBEKbl1
enVi/T6cU5ut1n5vjG6Nkovct7zkrNINs9vgMcKatmpWwdvimc6u8EXe04rOIx3aWDYc2Q+O9Gz4
//+S33i6FxsLqE4OtNfhAbl+NzfVcm/cJOGeYb1C4exSBKy84gJj3rviAFQq9c/+jxcJ+wadIBmx
qWgPCQoOtsc2nb43dZICTYiD0miuxpLyWIRKvcwnIfuTK03l9fR/aYE21vPrKzBCe05EQLjvyaBr
jvBY01QgWZmDpBIi2IAY0Zo+5M6S855zB/A2vgdbUANXn4kux8QijAj7fDWKTT2Me14zGWGWBy2p
g4udyoy0TNWwOaEpS3tLvOWLkqbOi5/7TkJaUZ7tJKz7whJTOurNyLbY/2AIyV7h+Lymt5TvXqcC
LuXLvHcVM9jAMkdr0j2TmTbhPOGM/JTqfHnG68l0Mijdidu6kZuLe3gRTmHyx1OEQTh2hPVayKiu
2stZ14H0w/SqMRMmLaQ827A62Dm8RSvgNBqDk+C5/qsD+fM3RcoDTJxenegoIIszTYGnQ1Q/YJhL
39QtuiUn6TesTMMgjB9W8YwrOhRWiGt6ThVEQpRwtQXXH5pITlisntLdVcED9vRrnJQahhqFfLO7
W4MxexqLsMRC+kAdpgrsL/I4xyUo+A29QqvztdrvLx09XOjVPbovv6GWv8WTVzQWpbgeOWC+5Ct2
RWcQxl0rcKSQW1CUdgVGEbkBoFfMSjaTpmqHNq6GMLPFIMW/qVzomx/q0rffAeCLKy/U1sVdEjE4
OolSpZkCX6hTSfeIq8y7tUEdB4AFvnTe/uJH3w6D33CnJhwWeUHgU22pVf0G1tI8lzSXj41udo5J
cAfOwsYsbEo8BBvwOnTfBnk0dF/cNIbPB98842p0dDfuCaGPQ/iPsO8r5ZFLIdCrMj/DJyFNxnyW
Ozf9YGvrPJb6tXROw8W03IxQLqHZatu0CewdADFOR2vQ4+Jlx6hYRDm8b1p7u0b8zI4qdJZEJgaj
/4SzYBPADX02aIaA65WgJrKjw9xeYt5TZRzVRaymIq28NZUw62r6L3LblQDC/gQC51hC+9L0xlFN
z4Y+/dVyyIma+JaWILT/FNAl5bTB9vNVCD2gRzC40+ZdaJqs1x7cpVAm3nhUEzXYOv0s3Sofg0Dn
+WOXyyLViY0EyLIyeD7eQCYbyzL5hl9z3FG65Gs4NVwk7FH470A898pUdM/+krsBBaNpo6dknen1
tSbVdv/hQBJ3gKuW+fwTBgihY/yIt9gRF+U/0bPyQNwfnkG1ItT0RVb2b4mb77pswOCxFjljhf9e
bC27fmDphMsNnmxznIbtxqIg18+Ve79voZ1BZzkjUEoRx1enaQu9i76R3jcvmrmDB7AvddC1YyVW
3XudOB1zcu5KUYYcS7ZUjQHLNbqlgFVlJW322IICM9YYfTarG+Ej2cyOFTyVOmIot4mwRYiqQ3L3
hTJuK8bTP6nY6uYR9bmgOGJKg62tN3i74UE4900i0t8+6VCJtVF0vHCiC2UvFlYy8Fc5/RSmMT3a
bbI0yOgQngHLrnow4oZedNJkhyU2wG/jiOSjpKM5LXCaBHnj7PVlONpzNRtvi2CuCpklhNdTDHdf
UnHbmv4sk1iAd+YayGZfx7C+Odz6S6KLCjLgMXSSGANE6kM6u8uduCmXqp134QBSG5rmaPGEM5qe
r34ckxsR6Ce2rH6yVtHhIK3x2sQzC1G3yl0pH/cTnPnOiJOoXvIVm7hCu6sswqQPq+Sex1bX/31C
kN316pKE4dOJySjgdbuxpdKeGofkASkybKE7OuPt6jEr94RciBR2lpTYx1bniR/lfoYpQmXYdkMx
m5E0Im3LOsoSXVCTOxnnqP6e+qJOLIQn8AWgg2Api2gHohiyStinLD+DlCd8EhHrbIBia/2F8GPu
RESnz+fIxoUFYTLbd4b/qIEMPJ5zSlNjaqn5qkoVBMUQaS2d0iVgz7O8P95V+CMKLh6r4306Gwtt
clmfC8wPHq/DXijdj8GaseXRsED2zlrlHEC/8EvukwPL7/3YRNVYCzfpTwMn5mY3NQY3hGqOOt5Y
32UcQMJ0JnrUh9B+JndQLP7eGNKbz9OVTgBSNryAFkNHkDc/YFPoqbSEvIRfc/xfDhzC5LlfFe5Q
Hnl1r5UXY2d8xermpUASDx9ILWUfkRKKC4PLfxeEymV9oi6y08DKu582tItclpL0z2K5dJZ9FSbw
15Qn5wNXNh8kKVJJmwxGiDSuI2pYQ64TRKaAwvihyC7zhLuTqm2XXRFDO/NNKtGc+qhHUgXcO/K3
qOGMzIqzEHl6fiBei3U+Th0pp0jITGsTxcil1qbsphEil4TJ78ZP/lgGec9UCBR7ij7v2RKs927r
e42a2rYCJtRQfUGK24Rpkd1E3P9W0pJIct0cYGhh+WpxNyDOI3A00+Jk6yPdWQRFFuRAF2MpLS6v
lQyghn15CLTZk40tLd10gyjffVPeTx+tfLxKalK1w773+3HBePLiylTvN8c5cQgIqP25jzi/Pk8T
C4I1s7aM932eXDy0wXwzwPPv/DQ3oXfzogl0UId7kA330IoLeaSq8xN7vtKeA37X+fs7DvIcWn7B
mIuoCXLaZ3lfvYksne8qEtL4mzcHztbzzu7c7Y5YxI1bEsH5WtXJocI5FguP5100KJ6WiuNqmw0z
p5bD5BfrHUaBt4/Sn62JDk6UIB6+g544tTUOoqMkHzPM6vy94j+NMXADTLWzJeK9DzmEkJ7lOwK6
sXg3Z5zarzUz14wUNLKnUQL4/xZdsWdFLbjuxDsEoIy6+XNQ28w4QuuFXqPymoZ9oGibESOTwTEe
2x5yn49TN5arn7UkY2YbMoY0js3U+7WcxJOc28AZCbBAL56AaFMBd7ZbWcTYbMcpCRRkFiunCwiZ
r0VRgsoWiPygKZiOC0i+FtRSeL8bZiK9OBf/7+Jlwiq6knpZl9P1hZ9IdV2oMvEsxvyzSDRdNN4u
JpT+6i8+CywXY+L9D3T58SmD9mZizcdA7aajuROLc8IYEtZnvtfiIc5pX52cuQ59MghgzW0AEU6S
AhHTt/j8t03VDVxmbDV1dpHcxhKxheV4/T6ncfALulHS9PkLxTD6fejp6jrq19UbLLXtw3A31T7q
ga4vxF86J4o5qrjF+FIbrxS4V1u7fIX8/+NxJxyLIgJ7L0jHNyCALidWM7/h3PS8u8cZLQNExO8f
xtRu3axeolvReWj4UV+DhAUB7xWSLj5ffCVHMMdCpAgefbGdQuiQzkDlNjfB+a1Xb/SMJOmmnLUL
NLLb6JrpaSk/cpnM9slTbcsR846EtH9Et+ReH9I1CWqNUQXqZM2DaDJrkFhV4cjARCZ9SB2g4PJ8
85oXNQak1pJdMIMOK1V3twtrqhhyfOjejHkMLVKiaw42OwwLfAYKCmbVQqsbSlnhV9Ft5b+OZJJY
xFdYB41PoOulfjEXe/HgGHYDzlbrtJfVbScl5YpgWgw/R9l9p9BmQedyv9LEhtHedJkRPJyQX4sd
kiUTPdjWz6wNMgbO6EuMZVM2FhOcdkArLE7NS7rLsYCMVNvYIAL6GQ4sxtasFQS871aI06psrtXq
We8tutgT2jDTdAOvSR5mB2BUKNKNYy3bW6JKeoFlL50Pthqiej9AGfXtGEKb3suyRmbCdhQ/xPhD
5rXP5rAOjATPFEFK3EFEYiD8M/9urHuiBOmODct6Mgugth+SvqPNSr0OU4L0as4d3gknsFqS4xWD
lbif0nUCaL+6kWEBr4cSP37D+uMLz8Znh4O5hKoea3geqT2m9I8Xngl+CD6OkzDdP9L6TXPQeRv/
11JreDsbVS4Lqn/f5IIyXewuwZ+V1PelwVY/SzwApls0UjZH15ivMtO7MQCWRTN9MTKASCcw6bPb
E/7E1lRG9cTMPQMrGqQgMZqO0bLzBA3KiqHtEJq4zoEfAq0t55HxNV/tTP+ldzLcctbGhWgetYnI
cfvBBqRJk1rtmMQWKZg3RiMZkxUDavyQdIWw2wU2FOZusn35fb9OJMbmtVoKZWYj/NNH1l7paj/8
0trgL/O7n2YfU4VOp2bcIZy+LZIixs8C+bKxyGjQ84/v05Q1A7IDROq7/EC3EfSTtxByyzse7KZy
VG4ypY2yp4+B78rIIs8w3x3G7qcMrWDupA/W6GRiljK3n+rC+hlvCdda/TTkU75IdwZvhDBGVZWz
nh13G4qgIQNPB2rbHHWolFdeQTCVt25X0lnzVg1ZW84kGrTiRQ8d7r8CPfyE/qTq5vQX6vy8ALHi
r6Kt3Ytwd20w4P0KHwEBg088aWsFEgxx1Ycmz7K1JNQky50wq5wiXc6aUzWVy2U58EmkFCOpnNL/
sPvOAvz7aNPLMmtGGxMV6qt97oNCVluCeBMe5Xyo0Mbr3GZ3+Y7d8OxMq9yjXcaEcmbKVholWRS9
oKo4ayi4XD4tnyA5Sv1SpUppql63kFGsJT0SgU0lX+WXW4vmrRdLwz3bZA7mY5BIKmn3W9/hYyin
QDXLF8eXyDNDoNyoZCxPNB+gFiJP/Rp48r11e1yasxP8PLZjjxUty67hTcaSXa+kPCsMGY56zHUU
yNKpSNtYy2/TPY11khlM7ohkoco6ql7DBN6WD/hcOkrA7AnXdfi3FTXOGwW9WVlRsRB9lkQwYl9M
0j74w1ZD4ryC1ZnyQG/E9ljYhM8FqsfgJygxGR6qvhHOnH0GK+KAp4z/dlXA3yQc8OyuH3qlUVJY
Z7eRzMsaVFNFNcEsvpReJyr71034KGM+HpMgVsLbKJYv1ySwJ9IwJfeftMweKFDYwJdw5B/qNfdw
4PIO7rbWNURim3v2owkgUrwSpJgRxx5i7YOMxA2i2vNnRa9PKoiMg59+v2QEaFKOOMmOCCbkTmqU
ja1iu1Hm53EfyZvsg+LgtvSeyW9GCKbLGlTcGpWA6H/+TLINU0T89iaeqDm8tznz7NSWsYB2z8o0
07hsSSOcYD6gmUh7z/2fND+v7bcbQN6YoEmfcoJUcph/biYHjeKNTxDyjoc8FQyZuLGEGK1p8puL
+SgzWQH3l76UuBH6SV2E6VqqHI6OXIBgi3A2Qt7AthWJ3XxybuwxuAaEO0sUDtqtfBmqewU0TGKW
d6TEYJQxQdKI8evrNDcoZGLFfAQyayXtzOc6E9kXLbNUWVutIFIPRD1oJ5IMpULNmyKLA6h8D4Vj
XI3sWKAy2A1XTTE799ujWpTeSwbykTZN46bbFsSc+bmvjaqfKlTlcaAoyFwplwq7xnv/TENumTFB
8lW1clWJ1gKa8K9zOmTdht6kErcIIG6cy4/RNoy6RzhAoNn6GrE8bmUCmgeAk7OgmUalMZPXn/L3
+6hAlC+ODrnZmP91OxHb0JtWWztHYEvGo+nlJlv/Lm+wqgMbQmbsBz0MB/JYCLMqrRacco/deJq4
aowRk818Fh1vPWN8Dv8Ndk9WCleX+zK98ZJa+/DY3nCV89C0doCiIDSM4hvV/F3Gr9uUd3NNvWgi
NYDjpunSQRYLOfJnJf4Yz9TLEhutiF+2sCatzYA+ZXcpatUEO9X5HCNVlO5Yji0uc1awAaqcfTtB
Pt0Db0uxkQsfppxkjrAMpb10pHCV0HYiXr1iDG5KNhiodLmk90Uk4mQKO+sNpUBwHkml0WOO9xec
NWauKevmYxBSrZ0/e5K3/r5WhKb7PGtstyaNXAf6Wz/Q31+DWaPe2i2kDgXu6CGKVv02QAxHnWeD
5iX4CeWeZa0hRE2mQTenotJ/5Q0P2+Ch8YY4iJ/rDk6BUxl46nuUK9dDdVsl53RDpU1k+R8c4MVk
Zx/x2TLCr0i0JrDnpeIe5iqgwdJEZrq5m/t2Yyv/CiTWYtZTBJBTDy8pzlRXuEIg7B6XbOoWRcnj
gIBJw4IdOcMP8mrO7wc6dqEJx+PDnPrOKTx3vXbQ73VClHfsn8Xtt4KaOJCgTNq0uSrpmPDk8GKY
ykdjUUbLb6b8oSfoHG3Eu5cqv/oG8Wzi3bpYiaoPJjnuPrGGMYctZtKT4j473qjK2DU/D4DpVgvC
/IxPH/O9JDRCi2VKwAQlMA5eFTkpTs/BkSrgYlrdGyEv9DGKqZzJO9BZSQignc72uhU9QFtHHUyx
2S8t6v2ul+Dn5Xc3lRI/K+wxIK0w+FCKJfzNCHv6B8wxjT/Vgb9rf2hmcA8bH2uCymiLtCt+32EU
iGS5t+gKn/3mg1mewzlwieiGZwAUd0tXYDS0HBOptCy+PkmsrNzcT82nNB51WpBz8voYcCcqJ6/5
knDyeK8gTMsZ028uUSmq9NYWXqTyXCmSZTI/O61JPa7qrfd80hsfqmcUCsYdyzWTACWHdVMeQNqD
HLh4MjIZMq9tSW7J9KHMxlIjzs0wnh0ksKhtDuNNOKugnIC+U/qs0EShm22+OwR6JDDOpULgRIuH
fR593sSM8TeGZ0KVK/DMv9mcoLr/fhhgdEKxZQirhLwZwkMaPJkh/2jkzt6r5/btjrIgb8whVDP0
GoQneiRbNNdB8YIRo/DzQqFVeFeHOShOkROv+jeHGBMv+tEMuY5bDgWoNExg0lMYx+WjyIDzTDDV
WnEDaVE6L4B7VURMFVAD+eYRrPWgrOMI7j2m7qIjvzqRChR+oAfrf3rKhp+0+2yOBX2Au5xTqq2+
BhumcGZoGQOMBDdqIEx/xtpTtQKd30Pli6Azs0zjBxN8+kvCUAYfKuHVNmzmw9tqM0oubmCI9GEW
soqlUTyQsYz+F8tNIQJ0ObxAW+YEndsKPPd2Xs8Hjtos7lpG4pY+kbYvO4PYUdOf+G/v0jheXnO3
fidbdXtNqP26RtnsSCOzsouVlMALWO59XJcyE5XtloRaRBYtnsbpKIGntleUkMyD5AvT70TWWYE1
tD1RuzT5VW6z3uoOMShsdehYaXndjebvUeyINT0scQ7bEkkEvuWQEnagtZr/hfmtce8ccwLQ5YOx
mueSqoML+b/DtGBeDopNP1478Dm39Bg9J2A+P9Gk7WgfqGW5RB946FC6FLpvsi/BpPGcVWACNtTB
23m9E2lMWb5uq0F3eki+ADmal5anheSjBzOwpuQe+HdPe1t2etX0RRGv9OxZVba0fiDd74FH97hi
uEXxx6A5FDe1gS6HRiVXdR/GKBAUAypBYeMCShIlCmZFOosRRIixQvfzlAkfBaARYhdqFduxnzki
64v7DZKal7BRAVy/SQDofFUcVJ/A5+gVm+69yFgN11b1/Q/y7tdyqZMwjxninDoz+Ubh/SYUBtn9
mtm54LfLiIX/UgAGblbGAs2Yj5s+WzTpRfnlEFOHhu0uYdy9Fk1z40iuT09xilL0EVefL5MQxLJh
6GX+89nMw439i5LZQpdlPfOyGfUOhY8DT4F5SiF73u5F/IzpBO9E1yeJ6yiDJtPP2gpi9mStXTsI
Ls0pA/+j1XP7bPUe8dunAJvqn02cjStaXYsq8kbDGKQ4PQxMff9R/JmF3xqowmG3fT4Jw2QTNbTS
WcT+FbGEsUKwvMjeGgdpZBuQnY23CiOjVb7D7qsR76xwlVtULH+SeQlryU4EUERahHSRM0TtgtBp
nBzfPRqF8I0nQx5JGMQeHBsF6VJhZnqyMu5zjvmgsdxlmthMf8pV9ndZsHnaDvmA8AggL76sk4/A
1sCDMdZDWyeMnrPDrm18C0mGPT8GPfzAkslSE8EWGbPZF9eqp/hsa+ybRWd93/QnhpKAbjn7pFHF
H0WlXEifOCf8oFJxgI3CtLkIq5F9geRlPf7DG1AN9DACd52MvxKlAY9wt3Q2KR3CNHyWyhPLgb5P
Sa3CPrcMTilSgNohnRD9ZqAGbpAb8Ix4y95AEyGyqAPuCyC/BGurLGL8pkDTBc1fycYHXo68tfOv
yFGIeeCCVzpP98UZmWnx1hk3mvSD+TSyPS4glxQvdCpWeQt8ABVUPHEYam6g5rotXRr//K7IxAWP
ler/eKOQym31MPYvBqCSqkN5N0dSA8/nXT9s3BGCHK3wuSHaVfrT1lblK2dUtl+7hGX7avLzp172
zK///MPyOAJyt3yPmplWDrpsOUXHlhwdS70UL6of64jGjfZ7/AZZ+RBkAa94R5KbhPR9swnhlbRB
av72Xs6yfAwFRq/ftGWMX0NFcq4trwdZQyGNvttyOK8zTroDIrtfRf0gJdKCnaAYu4PP4MEPdlu/
5hmBMSE7nUC9h1Tk0yo+8NRSSrOuXqq1TAIvNuxSmMuD1mb8iUwLL1N2a2NiZvAN0ZlMYBUMnem+
iUfCxXyJRPHzMQPRAd/Z39N3ie5e6AVaV5AMe2e203WbJv0SU+k7ieDpQQnqWm+J5h4n/2n/U80J
dL2hZRUFTsQT071GoaQ3ZhbzvnJmDp4CD8HhM2UqJxng8mQfIYyh+u4eaQVQhBWNAYVNFR48upPh
uOpfg+eYfApL9giywDcV0se7KQs9sgNvGvzbw6qKZfeAAi0kpxsE60potddYB9DlWvLwbovjc3x0
3IPVMBtBR+PatXhGMPhOjP8vDzRf82KL2js8SAlzgdQt6C9zGr5lUIYQY0uMAmFLxURIjtfpfYIi
b7pGBvkJFZ4l1uQZ3zv14aek6BSzqAhDZRCTMDetvsYp+FJYU0rV8jm1VP8Rtr9FKOmI/H+1vaAC
39EjLV3awMBJJ3X7UrdUJk/oaVQRMMlnNfVZA+YRgyjkUV1gZt6W4+bfn82RudsNcFdh2NM1kGH2
hh1Hkwy/H1hkc26JQBkAd5JApUfFNWzjZk2pAg3tY8pNjhQetnoJJZ/865Bp1fHc8YFL9afXAjY8
Pqk7uG1P877S0FRNpEAhXHMBvzaFwHqdBYPx2yx5bqW9E5/ip59yxL8D7pznF60aFF5WJJvhKPLb
KqX3ZOcmsNBiYGMSA8cipig8VgInYBriYStxpp1CNBvrXW1ma0tazSz8uILe3IOGRiQsMW8Ot8ez
rrOdnConl5OUFPXLbWYfb8QSUSYphBMQ4pTLcUdXssnZPGdY75gOqSlJ1sJPHcGfZFpg+cqmlkpZ
TxDn7r5rVtsnc4cAuHLkPoTwwKBNAazmWs0odur2EG2d5Or/zuCLnJ1V7VVnmdh0HPLYNQ16OZxN
QdSlFJcCebT9gD6FsQKJUD1JwA2YaiIbCpq72mOQFnkqMGDO2PFckzMjclsGlTSw+/dS2R/J3WRz
3zky1WNcqEJmqQ9R2JC0dXyLzDua6Ct+fJUR0WoO+LSmBVND8AxdniVdRNc9V4I16j/YPI/9+8hB
sYT1SanuAm4KpydFaKuyEU9EOtFzxxDhRtRVDI8BEN7oQ0QlPohaKJVb0tWkdMeBkm/BwrXMoqQV
DKnlB+0HJZn5TmEKIEupMoDgbL0nLWv+nRRmpR7Aoru0Pr/CATBAK58mWPsHfdzil0bb7s8soNFr
t3VY5IRRnFL6Qe8OPsmfPUQqbS//+BJW043bXMNDPrys0Q2FUHt3/E2s/uNGmUFzFZFqAik+sk4i
E3dk/xUJfyT151xfOf+fvX1icQBUsVD6GyAOIhs+tLcj45vzq/JNBhgXX0hmzl3cEVr8P3ofE/Lg
PjSBdJB6x3jSbt1PRSX5HyMkRioWAwdiYrg2j21VpsNKU5Oz6lh0Bk2LLfRvvKAO2KsxFr0Ribx7
hzManed8r57im9cqsme07yeWJRgjdwDFA7mtyY4/8smZXI4z/FxA6kn1P17UdIHEE42KZLADMbXx
DdD1fmsPqCM6vCGK+yt5bwQ8DCrIor3z9whBAl2NSB2yUQoHqfPKvQ4LQBTvHbF1FMsNqIxId94e
is9Tca2AvYk6POWxG2ZorYk81i35SmHAiab07pW1DPDfDavMS+JRcg/LzhS++al5mwvyq8IcY0HD
EBIts83JnqwgYdOGoUDt5U7IpLTA9/CBXSXTpwp39Ma5H+CqjDwPZoU8PNLO+b0JWLx87vyw+dus
Se3BU2uSNmhPPif9h6lLuwkGW+udPTHqFGSJ/CXfYmKLzEK/xx9MqlanPIv16gxOc2tgugixqGWu
9ttp7//TH8n9BUTU4UM+XjtFaS0w3Id+KZIFTolTQVhJDJDSAn1Xhz1iVvTi5RZ6QSzQrAhWthLc
nc0A3evmS6CRb/Bq6jNsgcHAWyBzEY1V4+OHLkhBhB+nmDDVq0TJZeau+JaP5mm+dPW30WtR9dE+
aPKx6LBWB9PGjOP3ecsl+t9CuYTyVRiOA6z0Ks9oZSjw8geeIrgrQlSjuEMV+R+GVrpya5Mvq2sD
Gxrer9Pz3Shg74LF28mw92QWkwn+dC4D0vGYqBx6cfz/xd8Q1DJFLJaO769iZweS1xFkeJBOPYtF
iiRhMCjafY6uhlbQx/ZzFBsFACzdVZxr+EBMB7rPZmXhQvCuFzSeIAgyUrmpLV7S/v7DCkXnvPUX
TplW0MRQ9/BxkMiOxGYYW0OQ0+MSIoMZR597LTr+hVfnht2d9y4fXwKzJ/d9JKwqG78UUOnf0lWd
Dym+OLLOH61Ae+gruhCnkW9lK9YwFPyEWZnYX+nx+Mx4P0Iaxv8cQlbAnUIvi3ol5MzJ48MPCCJ+
kXXAO2gmT8P9pfRXNoCiYLGRkhUO7h0oKCIIgEm2PUDmQSd2U9nj2aP70ICJarH8N1AEvHIByEQI
gZ/9xD15c1fNlAj+Zc8CTRTOMp76YxNgblG4e1c58cmAUqJw2PW55bOyE87iMCafOWeCEmu50r8C
IKSO8FsgA3swG4m7TTn3CnIRkBN7RCOCr9+WuJ5S7837du3MiRFCBK4Kgkp26E/Xp5AC4jAMyIK9
7ECd21EIv+vwK5SzK9KRAph/20y47abrBnaPk0jJYdf80y6vJQTD6sYlqGpPZdM0Cbq/Z5aa2ef9
YOl7MIyKI5/qScdkhF0+3alCqQY89i4820WJIlBsWcLe0OYmgCAh/8hcP1yaSOcRrRmHOYdK2QgV
CvP8AGoGV6ENJt2OW1XeDFAjrDpxP6/wjUfYxKgwh7vL8xm8sK2XkZ8Gl+0HciJ7/UPOt5qCKfF1
RfEaIK7x9rPOiiB8JFXtqNLJGi8eTmEN0eT3ftT1lCZqyf7WfJ57V8n4KGu8NWtZZN84g5Do6yTV
nJn6MMp6cuItJ2RSH/rwiThkV6oLxZUrnBeoD54GxrG3xFGdqig6o1gw5Ddp6avZBD5ARfnhhok5
4y8CqdeRN/hBhOT7TOFRy5N97LmdYW3C2ZwNwGWkziuw9kEOijxhq95OkLDYUiw4lyLpGhTlFc3J
2lmTHt3rHh6p/iibCzpFkVZZJ54hYuBo2t9xwvvLu+km68ilPld9op0yvKXyU9RBMLT5lUxBkeOi
cph5D4tWIBD8ezTJcgZ9D5MwTP9nNgseTwoy3s0TDjr7FWf8Lz1ENC6k4j4Rqi2tkIY7xmoGN93b
shQxi3e6XkBZ0Y48ZneTC23prU7Wwf2tSESvaC6g2dpAqXFZPxjRgmVzSKOnA0Zhg1nYpzWL6NRs
nY21xl8qgYT94AZd0C7ds9bo+mGW4dwMQ+Mg7jzb+pzH0YGnbXXDgB9Fj7gnrD3a2YxOPml9cG9K
uId3DnheG0WnRmGNnU6nRTyEO4oZgI8lhjgMh7qyqc0SmfKiGx1Q4shpqPO2MHNqubFZIP//7FA2
SILl0tyZapE+iqiFjI1QPgtoi+8uKzKJF/K+Kh4M0XrmArIibi8TYtEomxBpk9mvRyA8Jh8BZ57S
7pBP5yaotKRdSL8mlhQOk1SWjewcoUgwxnK2s4PN/6bcrXx0dm806+19vExhFsjD+nV89TDNlADa
wTNr4dR7j1UpCSd0z4RFpYzLEB2bB7Khk35u1ek5h23MGY5a4Ux9mja5gxLVVVmEkN5024qqPeAn
K34c4XlsM3WyL/3K1yCXOsKSlZ/TpJ/jVYZH7+OrbyLABYvhURDpbrMQbdJtkJzNOwrFm6fp3B0X
xcCQ63lYIOxMriogGmYarWHMRDmoZhB2mtBRGZBMr7E6hjLAfBgE5iMABAF5t7YYhrcm0mhEeoSN
Vk5favAlyh82NOqHwJIW4+1woWKl2zyk23hwzkUqq7xRKVlRZWSgebX6M0Io6G4EZWtVGJGYMtuL
4osp95z4t0Kq36eMcrB0l7TuVh+WrffaWOoHVtvaZDpBMTL70qbnYRZ6SWDzcJo19LbHg+thAuWa
q3Kl8ajUJBvwG9DWGV9PeSc+gVcjRfifi6OmG6tHqLd8cieDftBMNC69+H7ZcvURyR4XVZ5yWs5F
lERloEGjTxrupHXHsHGAcAJDJswV7iyoBW2uY43irCMLv7wrhLGxCXPmI/Q/PBfYGPvqNUmCyQh3
TWwQoJPhib8cQtdFFMXbNwYF06W8ax9u1/ZGC/C/UFjimn22Z4VR3FpAl3uW+1pXdDWah0C5wjwO
3q0ip69LjP0pYUATvCWXGcd7LcM3tvHsFO7ySBwsaEr1kQE6Vz6OSONoXzBNO/FSg47chvX5XiI/
6jGoLMxyO4NdFbUg2v0A0YtGQI/+FsJK4AfTWvqTG8tahoofA4d5107uGHOCpGznZ2IraPb9GGHM
3ipSh8nSYhnRRnrf4GItvZI3H8thZO/RJ+l7G9LqBc3TJvJvFMjW4dYe6W83gNs3joluCg8pH9jp
qRHr51zfGlXsnKocq36I/AdIxcWtY9v8UZC92QUmrd+goeSjK5k25WgFpbsVtrp7EYPHFDF+8Z/I
m0+vywhSz/m/WgebmCtLNrbf9ohJDBO7JWvFLxxv3neGcwRmqm4INK4PBeWwFsOVNyKqHlyvvvu8
mQjaAB1NCnxRNjMh/X0yRk520IMRpnxZZt7esa4BRkcev4umyOINdpzMPgiOwsJ+ahqT2rovAQFf
bJRIJhFjz2yCYpJA17YlxSl8SjMrXUwcsNSRYqDARRzAAFdrtsykyRws2Zr0poLTHuHDDbxq+mcs
ZBudslLDgTe6ZyYm9aWR7+ud6o8ekoi3QB2d2laLwGvhFfdga0J8/NSw66naS6TLrlAYhcL1Zi8J
ttdYexOiku2TFGPZyKxlgMpFPSD2hXzLTq49jO5RIrbuI+hS6cmOH5D8K74TbcZAvDS3ylRsf4NX
SPmAhOaVLMwP453/OJ1Jp1lL9ZVxOJq+9mxwcm/5hEeeeMP8KBhyUqxtYRqOg3E9Pz5WSo49+ICR
R30OO7hR5ewKbYlxxU/hvmzD+R/rQFJUDUpGitPt2O+Rr9qlO1FATTc2GGsXJmEJn7fHamGjW7VS
/CWwZgiTEHkBQGn+vAijDYBb7uiWvkZKL671LrX2YdDaPT4CIve0TGQjChw7y2Q1rO+nDU0s6y7t
f5jMyBC/lOGKDtgvt4Xy0yGl9bVQZDT5vnV0e7cr0K8QCnpD5o/o/XIssJPP0Hi9onUQ90pbl4Gu
MvPLLiKyWSghdlb3DW3wa7O5vgOPzQpWRZT3KOC/M0tUs/WTtzyV2dZr/WfAnOZFFIcHYAj84+pl
KfnnRtyIfO+RSLvJDQtvyseFpp2cvx0nipm6lPp0VrQ8IEAqsofqbXeQCy8afypFopO1nsZq2S61
kT8LkP6h2TQAj8hhnNh/66VI6PhmEwhMGEa/0IFEYx38CvF8e5F+QpaPLIvfJu0fcEV4weC1z1vQ
88UnIQ8oqAgbxhKXKR0/xphuBQkNHbdwGKNt4lo8kH1Eeii09RlwLzMg7FH8JJr0xe+jnN9b0Pso
aSrUoaVy6K3ASp+flVNbsxdZj+5WMNqPU4xs1Z2D7t2BjlrY45pZ9UPl9Lb8ZomPPKIoRtfCVj6s
x7jNWgw19YWnGlhu3yOrV8RkEl0FK8kFbkJHudyozXiG3RH7KY+1H58O1xYwppsDakstNFJLjj5K
4DqcMba9LICLmggy7ashVsvj2czR9arbjfxR5N3UdR6IKPM150H6fQUbV7dbw6pm9Fa8UK8Mxfko
1CKKNatBOsL8rsQg+OFRfQv7TWZqiAXbRK/K/7gydthx92wW/guNm7jEvF00o/z+7Fng/TBU/VhL
tHY1Jb2ZSqHP4CIAPkQLmBKztmxayCgbmZ39kAW5rEgcnuhqfca2XCTlYm/sSkJDFid3JmRtC/gx
bhRg/WOPtkS4R0rZ+YzkawmCnda9cFDajMd6lYwkJdw7zf/C1cruitI7zX3AIiDYiAE83oE7Kg3t
MzTk++u1LGZARv4h6yla1z6gpVwmhlp5gL3JHMyMpxSqkbBqLiMZpwpDIFkOPsYWPAZrK1L1f+L7
23pSJH52LlBAPjani/bOXaDpvJhQHI4s7IzPbkX0sG0OiCxneyaG6sXnM1F6hYcye5GmoenRaP40
2rAN6m69kqnrlJXWsUSUik8Gs51WRCRJq0bY7Rui1v7CTjvQhIlyUzcKBJQHZv9CowiaOpIbgZIE
ovBhcO5l7UufIzD63LHITa+BpvVp7AqQhhULuLGA0NcMteVnymke2nm4hmCKPZl3TXx2tkKjGnuV
YI2J4n2/SXYOm2tCNe6AYFvu0ESs4PbQzk0XO8p7cOt0LdUWIO7nLo4bpD2ojdMub7hXHYgTmt42
50ZOj2PSuBcMDogSnmQ1DawQpZpQ6+MtBboM3mWMN5V2tyrpEl1dmF1/3iw5aFffHJlpCYxY/pPu
CxYjZpBEzY6iaAAkIzlFnRkuSqfKK7T/Bn/uZ+eyJKTb7vSACS6s6d/GLSZZDxe9E4viM1t4gY5h
m4Ej6ScO9+baIGHb+1aT7IO+WnnCR6d7h9f/uzkIKuVULk22tUEeAwSBLCUBGm/fI+KzeGojMXpm
pejnzm2QBnoXK05roipaDLNQPaddeGjghLiSDdIMzCxS2AXcOiUZ1t/ZFkFUvu7qvuXmK+YOFTOU
L0pKMWi++AB2z97OdYxKYvuxXCsqMglKyPNSF/qDVuW6FgtrKnSwZuLonBtyot4GS/Q6gz+Hl6mQ
XwqOmIzF1FZSxkl5dJ6JB4cc8keH9NBtF1oR+8OP+SArmGvJOKzvQMigW9WncF/5ZAJphB2rTWPq
LQZ9oeohUH/5VyqKlbLU3tZYUxB2GQB7p2DWuxMR7KtZvvq7Caw1fQAxTbCq83QBQwBjbGQbmmOi
ybMKkSAHNRMd80OJhmODczgMG8ya92A4oZrnNQ7dlqHtwGJ4QuGAA/P+xctR40Jwe9Fyk0UQQkyn
qOUTE2nNLaRxlEucRkG/hgGper21JOOUYbR805Udr28dwuTiOkmI/pAwkouFmHK0V9OhfkOClbcs
mdSZxbGvRMyvscq6Um44ube+uRY8EuAVtOZ8kVQg1d7sNsMDFLMBvDhJcQ539skd7+fCZo+ui/ij
VDoml9WlXiTyoHBgpuf56+nFOVJm5UoOn0UAU5qrADq0cBdIqou+tzuX8ttqE6bpqK4qV2DMFi+V
4cpC2aG7tiHpK6gs2apa1C2149BkpjfJkuwGE5zY3a/+8ORXGiB1jpvcQHnBWCzT3uSzDq4gHwtR
GgExFD4syjl3RVJG4G65Bvte1Jw8MjcWTUZ46DNSkbDcItlvHqM+VtytXthBmmJILmAm2t2Hjghh
okngpuPbmaBhcYmp3O1m/BefLtAIQhuntmsA3FBajM86j5GYJiHuw2B+txWNmBOh3Mz0URi9Y6ch
p+TPC4LPlM9VVm+lV506RDiUXpSs4r3eXsAPLE3g3pO3drbkm6leAo2CNBFR206YKfoc8yQ0ykDu
ifHQR0Lk2RrMUf4pqDJquQCte0SNIigSZ8LoobH8ybxnn0xo29IPXetc2rMBsux2/rWcbzG3v9mK
VjxecEHwdOxVmYYD9AoscaCMNRo3mJeK9dGEmrW7ljNzLH4A0A9WpjCiUE7IHbGB781sfXeVfDNB
4FG1FHGvjxb87pQqVICS4jmpq9SH5s5GjlSet3i62FaSlNfFz3KWDYThQZ1wTu40ogsgf4Le2J1e
1C6gFXwFART7dlD6aC58Qf+pe9Zi7dt0RKJDM8i4ZkBQVOasq6OG3I9z/62Ww2NPiDr4DnKezV74
OgCP+Y7BKnDR5F/YPfg8GHCHnbZ97BTNcY+YJDOkV7aPbWBJOfBAg5SbCkg+yeeIjLaruiEUWpbx
x2Ls7cNL3VQodSVT2LvYW3eSh26egKEHM1ptmfh0+UTw3+gEq3vQ+IqaEnB8KfUFWQS6rwR5Dkou
xIpCjxizBVYflquJLNDNnfXrOTIrgnF0+yBEH5X9k0bmjEtNsrwmoA2YDtzghZI4gkz3Smv48LsA
ABnbsDdF3ToaJr2qISZ678S0vHItUatr6JzKkehI4LO7fpkyvyebgChTmFDWY3j21gCDtGePg0v2
UBl9Gk5PVRqcMTUHoGZuootoFbKiZclSSrwSaYOX1J0xzuoTf8Pk1QM2vY49qpSZ6ZNvAcZ4qxiS
My6EhhOxte3XGpvwrOtRm1ARaW9SiIhEs/wjv52GT1PTrWoRWV2hrdyus+yO3QeCND5EcrT6oqUf
mOi60lGAcG1Fk2BVSKYGJpVyu8CM6VMEtBSxi8eJ/GGThNzfisxLj6nmUOzEU5kS+sfTCaB32Y1y
D3mn9mYOhr8nFZwhMhvehLKKMU2oywsT4ZjOg0azEPUhTQovKZUFLn4xARdvJlH2yJvHfiDIHKgM
PrJBNex2ikM29APGNLnTd76Yfy2A74FGlV59ws/vstVIZ4nhNkk2IKdmy3jS7wMFOrvUMzbP0Jpd
9bqrBbTIXa2HmxPyA+A2nq6faQEAE+WfxRQu4URZgNERE8UH6wMXFwnpQp4unS/dAQ2QdtkAEKg9
1A5J54WjCJ6qV+c2mNm4sXDqx10jUGGtGW+HUq8zSdFeMco+ZoMjrDpn7zwwgpKN8Mxke/huiLDB
JSRSqTkH4lb8H6qH6brN1QHDPcEVoErynPcF7LJt1gl4AcrXczlzgmfiPmZRXbeXs0NsNb17B+TF
G/L9u61Pdodo0zHhlMe1eF0F3xOjXz8IrX7jG/BuL2ydjyPOTVgwkiYkvRXrFAmB7KuSQ16Ql5XX
SUgdCYoucZ0LeYb4/vT/TfQbkn39BRermeVEJzxuqjsUkUBOKslnUT0bwNfRrvmjAwNl7DWu4v8y
xuaVKYcuUW+sVtevSY9IoMfy7tYJAXx7CQUnckzToHT/WaASlo7K57iDVAfLSOsRLT8m+nlVQjQ9
luGjtszIDAurcOxDMf3W5brRfAVzeHQ0AhRAMKLTA0gbLMnPygT0S68negNI6H3G/n6/DTcEKTbj
C+DSof+JupuPohNivW7plFlbTxH2VaxY4QrTUc6lMqxVWS1RXhh/CQdcg9QuMybcq+G+X0IQ2Sum
nUqVEcTxaP12KswSAN3qXqbJuDp/L1j2JEB6WaAEI/haRllF5/Lr0Dl1Dlxb62kZIKvhCWPx9GZx
asdXbLQwOAeHKTBbu0dR9UQ+JHtrShRLpHzXMICpgD4JlEA4lAh5GWK85EZsF9GUnRqbksnolBPv
PuqcfqHXpa4M1xAso1t0QUIdeUa9hmAgmEcSnkshp8PjgAT5xdcO/IbEw/dkTAQLBQdYifWOgD5K
q2w0XLRKAV7tqxpZTynlTfuUpOsJ/fcEMMcL/M6OkCo0Z+blw+Nd5E+KD+suqV1Mzkr0ERfTYmna
HgTmvhkBYhp1WuRyTeS9zRc9z0l+aQdUcMrziSbpGOPIHnvBHe0qyQcM5ras2+5qsrdBWljPpPnm
CAyV7MW48PFej+vzLQeLn7AxtApLAydgpzMHXrZphkccg4Y89RkMoMG94K742osdsB1qUVDjCisR
b1t/oi0QpvUAlL1o5yRvWxiq/7m4Zr7rfP05lfvr3R8ZYbh7cnvTSwdZoKNRgDyB7gBeGIfU+sPF
/PzeWxgj/LeKNNtoKIjT2BPBnxu+iyRKNwlnag1WEL3n588Z91Jvay7j80gqKjlMJvoL/6q4DljK
oaFpDeqfhVldz+Wd0R7KHeaChl/bdoJ5M206mHJmDpykCDsG4G7vw7ozA8y6KhLUQ1BgxPTwCYRl
NJM0Qe521utQsJvAtsZRcPgB7yz0J94UJEHkd+ayYXRftsLj5ictWr37MgN3209ikOpn+cLOYow4
MD8j0j/So45iwrDAMvwyruQkBIiLLP651hOw9T/9T1iTLpoQEZWVrxlh9mrO6kNJy48Cpd+f7LvU
y2wZ6thVVwxEt+VoOwh78naWg/LN+WCBqAKJHXYG85YEw1AOeNrVT+83EASqo6lsAJeaFu8qX0zN
mgbrv3rWMc8v/m39PocV0zuoScYH9wp+GUSXB+3KS6GG7wkbZYzwTSMLuI1m7vjVOlw9xdH7euuG
z5pKaqHyk6UdVOlpoHkndUaGeXXudb3ktnSV4SD2vaxkvon5OsCRFB28g+9XKfN9Pl0wnbp3gwL6
5b7xKWMIYMM+d69MRqnCzzzWp+tP5mcjDKOLoDx54lCc294BumebtE6LNg+7M4aaLDL7aKTG0N7/
c6Ojv7ajYeZdYbm03XTJE2av1pYoiRqPPvAwyie1zHgDxuuBJSnKG1CzUVjju1xf6NBdbh3hoaoL
3IgH0ckcVJVjmzr23ZOZnouQ+H8vqrMMm1Z5fzBTOldQZIHmnP4vxt33fdshJpkJXxnEJLLvjNg2
RVNdNjlkmy4WHn6kRadRrU2yO1aLTDp/w+qDK/iXAJlaobsHo1fCG5hNDaJNNM890idjw5rfsWjE
OQwq/hL7CcueAOQr1G8jDRN/8+bDD0RWeYcOaZdYg+EPgGMhW5j41FU6njHbW+MJbT13vb0T6S0b
Ki+l13MzvD1gGIQSRNWuYgpjEbMv0cdKRjyNTvCNcg42b7tp/uTvEIA3jlQgAgJgTEuqpPlUydxe
325XfjSioB7c8W4bu5rXNdYMssn4PSzg8sC299Gm/1vwUi2fafjcGDSX/q0ts6o5rNd+5NKHWyRL
Fjy/BYFfRIiOd47YuHZrW0NME+QfcJeDY1PElPzer45froElS+dqeDfEmUBQyO5KReFeM1o+JP0z
ADIopsHYRhTpaELdMxn0yd+O/4og8CSN1o1ndl5xLmCw7DxjPjIsHVcZX/e+8EGVcAPC/eX+eco0
lMzVucqkTSvcX0MyxHW17B9oxI0W7qB5xuJyk/WbuJL0rDQ9kwZbxBxs5za50O9XHmlogOmwhIOP
JK4ROM34S3ymO3PWgCbURpFlT8i88UtE8r6V5kf+oegPJsaT0fsMOosZzoGQV8YxqZgCF5zuqKr6
EqqJZEAFrBzynMJDvigs4jmW8TuW0ObET+p9DcsPdz8pAtGIZ0fDtg7S7Q7zLbEkt28dtwC9VeY5
hzf6Mqlsu1fm30zd+S9FOrevJTCbNSz1OUMv1NosjF7+mRnIZCuqmQQMzc1a2b+hzMb0YnTBnlGt
/2Af3OAyhD7nrboGENG/kJXOZfwGKiFISS9T8YeW0V0tdzlsNjzpNJkSkf+tbWcl2S6BKxqz37oG
x0PZI99gtik/tDqHQ+kX/M81RKpxmTTwFKtefQ9WzjXFdgu1AQTnfqjzWV9FhBMFNbRCS838o4Ud
KTmMmq7P52LXH59exZOdidCRcpYqRBWFHrwtSjwbmjZ9pi5+w94s7GSf0i/xZz5VgBB49TICyEHF
gZcJub5BMijZjvULK28p8tNc9CR/caxogpUa3mWi9tBtq+k6blozFrtvPbwAKGlQnlam0FwY05KQ
yGXAUShwyo/cFtzailu3jR7OqP3Wn5FYiLgj0Bl8lxfU8a5nKuD+fa1wvHSnLlk1xXGALHIkaKsu
65p1viCDiocLBkrV0pRhmaKaxD/mAfL5U1wKHmky3Hqj5T9ecyicKnAG5efyHE/8uhROHdmzyWuE
zue1NSOIHhQG/wAGKQqXFpL+mLIkMboZsDUPn8kct+SypNk/0YY9BC1wB3WizJLzY4eDv55ek/aK
DKGEGvcaQXkQoIsqJtzN951yMmyGVNzzPFdui5r+2/JxTm/cERKkrF2jKYaDxaTY2nlbN1iW+7Lx
7iWY2gaimD/MNo2KCWYZmgy0rhZlHwyZuheAfgIOY22oDT2l9qriniF+2xrJqSUPY0D5n4Se9f/l
4vxiDENvtYaSrQxDOW0NcWZ8SPXl1gKIGBZ8/MmcsYGz9USH8+Qsuw9Pc+SiofOGU8BwlPDBVTT6
w2dUsZpUqxRM81oUvOyivWyLDiPWQBP1ic/DsznzAS+gNNjuEkIdZz8flq6dYj8bmSukgTt5tNAi
7X4d4xzgG56M4Sz7IFGVoqKI3Kl/BZTtpBB0hS3j/47TxzNI5uYlkFQdF+GoKztfXmKDtmlxQpz6
9ViOXPZWrsaaEtMwcJWIcYG+0YFW6WY4V8kOQA/dZVqaHCJbbKHWkQLiWMT6O9IB+rBf6C0Fnaqn
AYKcL8XSOZOPKgHX/LPeeZKTH1VEvzxbsdpX/guvtcjh1bEm7BY9Tf+n3jec6QC3nVjrSgaG3rlV
x6d2U2tDXPBg8lXn3HOeD/UGWj1ehYcYAwKzME9exGMcYwadTS+ygWUvVsfGwB0dXty30uiK9Xth
4QgXMBlK6g7fpTQuIr37KdmfhfD4Q8hyWctR5Zn5xTKJBTcW4fRJdFhMX9wIpwAlb1XgTEc3SRhp
a1N4rzxKJt6AZfuDI8x2xB60KkV+4DZGR6HvXYfVVUs+fHvR2E1azbCF6KkRah4GxSlBLucpJL5Q
vmJ90BplgIb30GJ7aadn1ei6EYn3tyf7iAjDfcakkO6/XsPi03GK7gEjY4mADUM2wHyC+c7GtQX/
1KNT/VHTmp7oGToZj0zp4Ba7ayEGaR+z/YBfhanG3kiFI2B90P9UwyvzaHz7LHXsuRmT0+JWY351
mfvlhjv82vHaRoxr4eDdAKNm4ZWGjLtrFF8RVBZugCo/4gSdJBQHoArnD5gi0hc3tvNTOMg+08GH
eB/S2KxR9pZ58liXtfti/Cu7Rnl0uFRJqweDs5Y3ZQcBsmUrVKjB+sfMPMZBleihYbR+pAJ1Ev+x
0Rjb0XXCTva06Ql79YaJOnrg/aUqh3z2Qgy99rOtfwWEExTeol38iAADSDYVIyLybxSpUBgr3TX1
7B7uCbat4Pd6MIrPD8ZVrFcwQKEa7mwQDHEcaIZ33ZT3K8WHx56KsZ12EVJxz/miX2IYHf7WaPv6
0xbWnW9ttunwxQjO8O10/aXyLz4QKSlgwHIFz0B8qquJxdxT7ml7unafss1FF8axjQe6iai0vMgk
zRnIx6iCt6vs8EQ0OG5mvz4cKIMsnhYowIsqQJeU+eO5WnwaSP1gcoxUQIj3o561z6TuWyUiD80n
YmIxTFEs45PPmDo0163gK2VHZpi7YX1chCunp65IwzRM9E2dfO3fE+7dGjePgrVKNk8mKrBgWt+S
sbmwVewrQrtGe7FDx7oJ1+Nn1l8Qn9JAkrKbDazCp1Gs8Oeu5D54lPwUXfUVzcq98wjXBogqVNlE
PKjiw9wrUt8VEgRpbFjBsfYW5xNppLtZ6zeVPnb7Z3C/NEcIMwh4+FzqQIFS2YNKnqwWj/s9UEWc
blxAwue2u376OpCNZC/xlaCLC/QsLc7NNxbVmsvpiRmDJ0nCjogPDI+h1jJ1XNjaDuiLaqeC5iBu
viVQ1iQrkF9AV17G5hoEsFKTIprthbSDjgWA7ooSx1Qk1Cvi9VN0Q4GK6DIUWheTutSoS7jOOXXT
mCKfOfUrR+D5sr4Hn9fzWkdFillLCtXWvhn22s99hKQEZzhskfKHrUZyKwIAoFIL044CBBCVM4Wg
hns8NS5Ev5TmeMXfkUflNK/IO3BYvywZe9UHfphlazTBCMGKGoh6qigcNWjl75BI8WXYlqYGf5BV
Jv53ckCvUDuVV89HoJLV/oClJkr26uJ+OeGEvwGtEho1SFUUQ8VgzLZW8FYE6ztFthxwSuEDyDd4
CR2Hw+L0MXu3H2jtb3lOr+5wdd1E+kBN1nEnnbr1zofpg2pQ8w5zOrDDLLTddjP0by8OKrhX3Bia
NzTuZa5mQ4B3KxuiauCnhBrBpBr2IK8xw/5Vux5/t7UdOH9o37elZ8qFjaIY6KhKkvY8JSfOIqXZ
FvkwsfkrOB1mGstjWRUIJA/cqH9gZnQpbxpnVfmRWfh1ZYLq+ZVXv6+cIvrtM/WQBEy3FBi7OZYH
8U+SpyIHDF1x01DHREamQU7EBhf8sFerMRJ+IGRuLB+7bHfYBlp2ZUxVx+ne9HaNXjsqgHm+xrZS
snUdYD0d0CDrDSfYkfQeOl11F9REiRt9rYCIWKawZ59mNpQbBWgtICuBVBnoGch/aYSGeroIEe4n
OUxz7GCW8gdQYQEFrmttYfE/OY9cftEnIjuHHvPEWEYygDod/xHHRjO0yQHREH/JLTCVsirSUQik
JJz5bbLo1bTYdzQz9ThUQ7XmkcHr4bet70vd19R+eyTISwWqxfXk2vEOT0xHGUbJV+XR4/diQQec
YiYMEdPMgezf1Cua/pKsexefOtpfm5gVQjJ4xJwSDp0RvQQxrSE8OZ8M8KDVZzFhY0t3h9o/gpjC
6Puh3LpUDcZBaTVJpBrb7qcDqG0dw1ByYg1lHYnJ5ivS8uCtH9BoDWuHfQc44yfJtTbOWYcuUKi3
FYDO92UMew0pS2BbhcWKdkyO8xUsI08q+V29kIaPeL+CcQ8Sn3j0uHIpEtqddy7pzy21Ck9JviwA
E7E48lBnE1ejE57AV29lnsH34FCJZaOaG6sXBexdqyEpJZWu21bvXeIi+Xi3DT5YVTLRcE85VQ3U
gS8rLLqaQYhgrOqbL4EWjJxzi3Uxr1vM6ASrBXoPkFjFSfxczohWGoRzwUmLRu5NQ3oC1KrP9BPM
JHPkmy/WIylGHy2MSONTzs9+5Xmj8Yn7bOcGmn58e5UNlQrjky6e29jiZwKl9r6gwN4dwHCWrQOa
ZIZivQnAEdqjkOpK3ALblgBwl+RPTLd36FQpj3mjQE/8DkJSTxhWSHrf1rcO7FrsGNutGTRn+qjI
IA0HR970ZnvoBIdDMg8VcBdfjJs8b1XNxMuKd/tM26GfNTAgQKwDubgyDAdgu7I77l46lYiqqAgW
E7cRG86izb+R++dUjXG5Ey1nMaPhy4VsOBBmXXGSj2rXpb4MX8lbcfjO7DM0MAslbt1dpQAtmsVU
85FtKaiUna6UEHuic8JLB8dHO9+Elq6vRN9rQmH3ZMja5sdRFBtdx8omwJvQSH9ix/XWSDhTiqJ8
1jmqkMqaZJT7dQCR9cgIgiU6K2DHv42Od/XZg7x95fjTkV+c7Y9SvFmv8iZ+QAOoTZofg1VzSvnS
PYoYW0I6CnqDOxfteOIyKGMbwQC/AnxwMpR+pDNUMzrriyc6MH+FWzS1CBBj9a47f9/Cm+P8lCtc
BZ7d2Bxcn/89+SmaMVXm3pTpbJaaMD59+lwpUYIvRZKSwinRKuSe4+rV9f3OLtD9OQlDrwoItlR+
5qN5HbujyPIGnvr9v4ZlQfYjR4bTcVCqzIbyEDXLcidV/ForxkHDGTU3BUMl289zKCAZ6eLJb2yE
AxS8LpMfOMxenEn4xQs0yh5Z/LXT/tYGP1iik9jUbFMQbG4Q5F1zFQ83a1iw4ZhFp9DY77jSNU2z
5T4Zsz7zDbHm0Frrw6fgjIfAFqSaVEeCdVpkyJiHylXtSDvFL+okKZpHToR1FhCjZZTScpSUCsDC
kcv4SCA+FoM8S01fYAsIJ2dFL6TzUFiH0e6FgM45cmip1tDjGz8KDHvwhExYZE/POGxomNuAqwP6
/QsvEmdqZ5PVN3Xj9rqbWPYasLNqGSGt2GVpey0GkpEUx/RmSUC9AinmbjoFdCNAtdQzaVCGsH7M
NvkS78rIu7O6F0QaE2m4EUYSN+OBs0eFtaWSDfJUykAKlmIwydilPGdGe/WtAij15Sy73qDiUALM
9iHoRhEdfHWaif8KSDNbP0N0D0duwU5cfGjmig6bxNos6EpbysIzkvw3uX+T8fZGi/CzpsQozRtD
ny6uMU3qNIixuNIdqikOT0JP7spmzN/5FsKruEpxqNVAam8iXpl+QxSZHVsorrNWeNuw61lVspGg
ADyY3L6P6CAjUkSwx/jZDNz+2/mVXANgUSW/HReBVLG7Tlg3QfTWJtHm9GMG973DTNVw9Qw5aSbJ
fO8RzRwnJZUzmIe67EA5gv6kGnHzUsFY4NVIY8s70YVmXQGNq56VWtTTc0fYc4ijQA10jO0/aPNy
HMdSp6sOZt7BjfGa2DcNVzM8Ky8wiR10/jOCXbs0pprCjLPIn/qlWYipDhjK0j7VV/MQhrwf7IuH
pSEVrxeghZIyycupYD1SrEEXQPvtCWxXGjhePVPFasibBFIeVamQoiCtFnagsqTJalINSb9Bpa4e
8v/A5I/gneD9hyVwFU+g8p+pyocU9toZ2dSIS69uEJ/aXy7Q8WWy1+RKIxACozrxb4kYg8nJiPw5
eWZxX+kRwN9f3GqsbNo8+cqNW4MzC90fyAei5opEtDjVntM5RGw781JKbPuHxG0km4YGVR9CJTiM
OV9keBzI+GzjK2Jbw7g1ubd//venTE3ORJ/rRc7aS+i9Dz/WK0bfpd765CLOr+hlMRUcmT9ZGzTD
yAx3iem/Vg+eqoPPUSv9FLQZEu49zIx2bUVZlcPhpiE+1bdGFRmYWMnCtvsJG/RBM9SwYGWyM8KK
3EpgJQ+iY3wyYFkcnIohR0/lJ0makd4nAu+kI0445kIiUlSD4PVCdKiYTnqfKMe6R43OmGvD/C+D
5BQvuL2SW1xpXH6XygPahY8l7G4ob7xsl3ljK3EZgUAM4tizKH6geUa130fdCOYIQ6cub6dKTBM6
hLEIIHIc65qMv2MmYyvo6sS0JxPdiYC/T2xxwfuTMqFDI9m3Ec34DFoThMjlt5DnqvH7SJjYr7Yf
8PQpFBeI7shap93gk5mlXJhDJdvgu05mdDu4e13aths65etoO4OZRrfOwNp7RiN3iKnGNd22c5Lh
KvZQYZcxOd71QFbCb0IMlcXvfpHQw5SIvi6G1ltO94thzbv29jHavKZ6YlnIDDusi9fK4XDX6rbH
lHq/ZfGOlHEdCXLmRNuEqRDHNTAzFV/jBW6EuFnf0TpCUDnGvlVTv8NdTuFyvQ+aYv1QwSUmWY34
Uza55DGc4qZvCsXzKpJQssSa7jnLUuQ4rpHwzQwVEc/c7IgPm78mRxnoiPXVlh6NESN7ogCIXWes
Y6gzTHSXv5dH1l2chENaiDZnhieoLLSeJuT1KIR1ih9aqu/mKvXC1tXnH/VN4VrDnLSEu6fMVGgT
nbyZIpcMszS5tV1btQDNSO+Z05IUMVnKG1wGW8pKULdsQ3kGzOHxrgHdGYN2+dl/5iAAkKanHaHv
AlHcH1ZCOJ33jbHov8TU2wAK6ALnKZPSkxGwQK2Af8hFX8ytZFzvAdn6o3nEyDYYrbWJNiWu1ZlI
Ew4OnnnKM9rVdKqjBLv74w5TWLH3g8VG3mmos8DJFtoxYidT1KfV+AZ/9P1FwIFsIHwfRYPjbZ6P
ojyDI6RWXIxs7Kqtq8gMGTDV5sUNVjqTxR/DG4TYCkwdPzFgekrplsige0HEd2zQR+BFcCb3MCSf
AcAv8DObh8nfWejV8wgHZ6PisgHHv94YlK9Q2+zUcBHk+EoJMwUa/PxeTdeoS30YfdqGxUp/cKH7
pd+/9/3Ntv2klgmJ+OAv8Hd9QS4UQVNdnYWFYTObPPfdLMYPZKwnxBAxqV1uDp3jtl5baOCgxbEt
Zqj1iAs0Fbx6oTv4zoWjt7/iVvJocK2FmMfSmUUK2GHo0W975l+6n/J5eJPnKyKbLtWc9EYTOLgB
Cp8AISiR4wkAWf5sUlv+EGlUhbt7eEz9pmvLXRKOqRHrIpCtMG2icoKd8FKBoU4Yy6EkYe8RGHw4
h6RuP+d1lF6xIGmtKzg9Ow/SwsgyiNMEOdpcadUUsm6nIUvcRIWaU8Eabtw/ORed088Bxf2Of7Tx
wRSv4AkWF/Gl9/C04itkpXNRrzpRwvYvJYC7kKgj2cjynX4Y1qoDTJN7+W+Z2iENb7a/wV5A8+Cq
DsJTP3dJxC5s+Z2Ri3AuehSt/R+Zz0fEBFe0M7Xn6k07z+gMPIMwl9SRNz5G8dyWfi9M4Xoswvzn
yRJzrZ0iP+l0MmuK8rSgvA6R4SDDuz3mqiYOi3xfm+xPrtbBT5FDaVGqJTLm1BKEV5GSP7DhY8bQ
pSxrNBq/Ns5PwGTfvA4Qg9tCTGUg9T0zROIh2K6OfFGJOfnFzwlUWiqRxRwy3nce/SCmGn465Tpu
cTAkPLhBCfFJYhtWCOJE2wz+T1BNIe2ZTB778tcQScj9vrSYM3nVndYQsbgeGDuXBcnbTfYxkeRm
7wlhmrdqAJxr1wU/7GTqgvIrUKrqe3ZR/qXs2pLfdx8yTHOAsyd3FHznb0g9kovu0znjSQqU9ipB
GeCTCSizCnF07NRen8oeRQttncaQX9HOyD3snWq5mBgrxNnAuHkEG+HjYIwI9CfgYfv0Cr1syLpZ
3WTJdoi7jXKBwpTQ38cOrMG/1dVrHFx1E7EEtGnui8Xqs6ptRHICeaHf7rK4bCnY94NUuplXOeK+
y8M6VNKzyrk5ck6XEGrI0ZMQYL7PIPbzCbHxf2eY3viGQaiJSibSYv89mwrSf0kNJvbZfUhOB80W
Fu7cW0BAl8Ca0p6VcqwiiLtcutLv9wQ1U8qhH9yJ7EOTuDWt8U/9/amksQQKoN5HyPYWkTnfRYSk
NiCPSA0I0/p5mTWSwahKzAuyTqOKEiJTWEozqF5LanwtYTFwgwYaNQUPtmKNIbpuNKOIRePSEEOi
dRpy+4FVBG4tKnjFJMKDOzfnvc6LMP5Wa0NyaX+VCbli39sdG0O9Vr/Nb7rFF4VLPKvFKvMMQG+c
2TVta3QgJ4sIeyD3V2R6OHyZFDzqlUvqlFwnZNqqo1PeYY2F5er6s6Y3kId2cgeBofW/8/1nvAdr
krxtSL/EvOpZcjbPlM0WSgyQZD3E+xBzRnZbAIiNajqVbxcrl4lfDG5m8WFJorY384iH2zRCNtOS
BqkH/7PicdexerRT5tkde181kFFNwA0W/H8b/6OCwEg6MXrpxSjfDcWAbaDZTOwnszQpCTvE7wXV
UJHjPX2KUISJ3eQP93gUc4OvUhwdkvvGMqHbFKC/zpg6hjX+1y4U0MMZ+lzwdPkX2fH6yXnokyJ9
ucm8bbIH6jqyS9MDvCSn2UkHnbJuP8hABB/ac0q2pRJPcibSLBYeUWUL4NE1Wts4anXUvjCSBNj9
yg2exRCxU2F5kDXzMqxe9JuipBL6HtkFe4CFsU6hiMP3p6IoqiRoZLYdqc4z268MfZ0rm6Q+okmc
cFTaAn3jAiLUbRTE4spIVTguv3k1Rf8lNS4f4HuTQz5aJVNnTbSXcFOAZGOmCHx1siMDTXHjoeOI
WhjxTqu8D+j8nfkOfVghiMsk0vfQkufOmAsNbx77ShVXcMdtZSfyL2CkOxGTDfZpGg5Kr/bopkur
+En5++DLhM5dTNWq8dm2jZJzgrRboWhUBgFbv+G4076xDvoUpUTMYVVqRXsf7f1YDh1+JoFTgAUj
QLWYmuT5KIJAQsLAD7nDnNCNooEtGEwd0A84cPZpOr26a3zTezGk2er1ubgxXMqmPei0STjcnfJY
ZkY7hXZ/HC1BfcJDu1FLA5fFOyD4LcEMwWj1lH1tkL9EyjdxiK+Q80eBeoVnPhDfRtXDOPgeKgL/
s7TwoIHQGjwNMHtI6kpet+DnYVrO4+YrgFzz32HyJ8lqg9dlYLCT4KdnP8Vq6F2bfcYpkX8mFTQa
npzbGdJ5PGOTriF7zavJ40pDBcJBj1ke9KKe0N2CO5QdJDU18iuvZmQ3Nuxyz7wG0OSLe+VjkQ7D
YDkpHK6NQqUmgjqRx1zWz5/gfZdfvhg2YAZ6gzZ0d136C6JOHQ010q2N2sBgzS1P5dI7r3h24tdJ
wkqJwOiB3Sv7sADQfVOCSculID4YQXFhid7N8tdnBKg4Y6zMQPXgmYxIr0rKLcDk8UHUl9Bf6iuV
o14a+OGNEvVfy7IocqkFR03px4zfvqYlyVaMcQLFI9hnJxXTcwOYWVLjSm+u4R5cSo3JGGUTP3lL
G6I9dyHEWgtcc5+H9IT2etLeMS0lpW2lqTVhq66hPfQK4SLL5x5h7IvIX8dRQedZ5fgjl733O5Qv
t7dKN0jSvcP4H7MUS1MZfNZl097MuOsZBtuqSRTNA1mtnKQ493OAozYgP+pevKF7gloRjpwnRdP3
Olu89KoVHjntOSeqcEw9b0mXenGGfpAaw2jZbdelNNec9J4A6F5hauSvpgcDrwXVJ1GmBvmrhX66
eMMLZ+f/yTD39/q9TAeXD1cRxNogAfwTGbOWaYMzhSxGswUo3Sph98+8P3pf1H97WhNpsw1xHl54
1axlm8PPrioZ3x00dMPDLVWOFt1oLrmHV4I2BLFOhkWJMs8uBqZjpvvwF7w+mrmIPo2nmb/sX+y4
eHzJGjcr8lnlva4HzCvaYxxmFWkirMn1ab0Q3alQwqcR41irsNDyFd2UWL91LkWzdkGtPIvQLLJn
d/gfXDpNWNZ4f/Q9eyhNtxotplTE6RsYN5kuEgY+gncE4Vfwk4X9AGP+OOjGMbJ8DDQTvQe+ECpW
Q/rUMXj8cG1xBKgupSQPGpuUk7DS2MQqw44RxJbGFFIo84Q59VS+oxPbiIa/irrKslFszyD3Oqxu
Ram6/d89Ew4J75CO0L55I2/QGmk2H/6UU2ZTZOBFhk1yeWUFbgkfQhVXdDJqCvDQnBjQ27oNgmkt
dmDAEBkVXJfB4vRVSrIoVD9wBcj6h9RgiYOPMjxkP0uXhPVmXx92lOx+LzIheoVgST5blsnX1vn0
ufHMqkvMgty5BHm7JJM+MiiG3D6Z3s3YewuxucYs4aMZ6nvet1KDAtE7VoOIbr5V8citrVy9pmpn
XCxBVL5zB3BZg9oPYssDqmvxaxdXVwieug1nJMk9v2BlzqEjw11qu4o5UK5RpEiOQRb9tAAEPKGp
VAx9+GKuICc5nxgVnlXzSdGOr0aYjo0G1zX8VBNh+am6GcnIqJTICSrZ3ujF7VAp2+121ggbfbPJ
ujAdM4zP+C8C1+3heA2cmRTX5BM263JuG4ZhHax1tHOrX58FG4c0e6g9ktSGUkk68IIVnACUwNKu
i5U9xlIj7QN/dccEOXQROdWa7XZdQqjuUdQ/XksAlGXB2YY1nkSz2Lp/0onCBtm/R0mpnDMLtWpi
v5Gs8VljJCD/4wypAFsXY3iR3gymrK+mMnFWmKoXy1LycGhH5sGEJs56iFUwBcuTAWxJEVXPx2Vw
sR3HkFKpggTexmqUviiHezg78p1domQikIKoMaw+bn6mWPl7XUxqFtwS3s3+Rn1mNcudC27D/+Fu
NgpzaHhy2GdZMqA2NKZu/a/2kcQLRnlct+SDVnhBhB2RmkRwj4WdKlImFAvgShP7jOyDhwIl60tl
O3FMM20q6yAtI+XDABwuSforBQVuUYS89Z3wFf5rZPfHk6gVOIaCTHj8DG1K1cMgpHg+rqJCtUB6
k6aZP8ljQuQHAJ0DTi+3b7ZmHm/v6M4GvcAbJQcLl0pQKZmSRSG+OwsdaypzLZqaSrWRrb8n9T8k
GUbGHE4T2yUB7k0HSB1kMJYTZ26YKU2OEFghZ04Ly4ExnvxWJKn69m67cY+3+m9PoqFAQfx2Tzmw
iBCV7MDE4y4rfeGqJF9Z4TO2d4wkDkJdX9D8y12Yhhlp/H6Wk1/0qu+CQYpIzwUms4wwgGSre1tO
z6i5bEM4USN/299NwXfSS7xZ1K0CgCzER2U6cCEHeuE+1efVYWRPBVyWiX+X+f1lpA0HdrPYFmpb
eDxEl4RybhsNgD8FmNllqOD6YPqykGhy3EkIjbIR96hMqCfMm71Cl9o6m6aby8ECLdJrlfwRzEAd
7aabt3zFT/Z0MpBBTSN2f+oU3Tx2++Macx4ZJeFpwatQ1lRZpnFZhPbz6n43u5zWgtic9J4zOsSp
TitE6pD8HwMHk4Nc3bbjzFEZGshTuP8EqLlNRkkRJrVjNdnXg20yHwpupQxYlSbm4kgPyfAVXtmW
+dgP6+V4144fveHsAm+hCmddB1oeMJJr8iOsG3ILARxMtRDD0JM9MVlm6+UvF82/EeOmJpd1yXWR
44b6mlPciiYaM3jwOT1dmVUskrVc1Q085FxiFkMQRlIHX0ywvVC+Hp7mUEY0WQ0iLyjBWkQuCwDJ
EKRGGj9LRx63PTCH3oVMyDCZSmEizCPLqJckOOQaX410hDFL14CvXVNeUnZSspylR8voIMrAs10x
HSRo2OSN8120sX1UnoYsSOdYxgT79uvIECI95dD2nOEeahHkEtLsywG5js27wYbrTLS29VQFeKr8
fIgxEG0Xf90yll364aRZuQhCMGbOaHF0clUd/2wpfxgPbhosBTclG+wzXiDW5U8Kw1ANeO6LV0pZ
btmB2JPOSYRyTrau0rLlNUgyTarVAU2avGpiAjLA4pktEczG3WWWBWiKnFe+CJNfEGchpMeU07gq
f84jIfpGHwlsy8xYSUkmMqHtXnUDkHaBZLcnqxVmC7+GGbaSgiBh1GLgaBHWqeYQyMJvFN94H0vZ
ajimuCDz4zGgNuysmsqCGPSPChtTqg3h8ujH3kzjirYZSCSp/5NUbEs8VXMFl7OkD5S5tgeR4S3d
DKcBiFAgDw8oqDqcZSreGLyerSdVrtdnNBbsy3XDY9WSdakuWHjvZU5fuqBc+9qzwLZsU/vmG8+Y
fYmSlgZbzMoOOg7JBDuHHzEemOJ2IhBXfJQLh4ajlJqtx1ZVzkhm6Gb6b51+rVkhAXJkJfx29jx0
O7i9S4G0JSIseATToZ83s9iqyV9r7UwkgDZrjo0m6uU6Tg+RcnJ8un7ayQTU0XqGP8yiLaDJ1woF
9OUkf6QuRFGqAmn3o9Q3unyypYZpOjyq6n266e8LukL65YS71ffL1ktW3CeatKz3/y6TpGTEjoy6
B690UWD/OMnZRaqRJ3uD1IPtn2gFP1ubYJvFRPo7MbpphoTlXlmoydSO/fpEYB8YNBQeROBKaFUL
/3q3cch56VvQo6gpnWf76g3GY7yIIroliusc4M7eSi9CfEwHQYJ7lqgFLNYq4Z6PDQ3LrSRrPvQD
evXr1RTi4MTEDZTvKo5sHwdpSKC8IdxJYOdglBNg+CFEsAHAaQ6Pyb2tPlseKvgNc+dl5uFXaHYq
7QIQ6kSfwNRszrpoCcqQ+9XTqnGjAHFIefp6dRXQBlsJEo5RVr+1hZQAEnON/T9GohIn/JMbDTBu
xpsOIFzgLJt4yEbWD2unQksIWC7TTut46aTPNTkXew0lcVph7jAkUFF8bHvRKNyG9dAWF6eBipRz
mXm+k43J7OxC7uJTRjubluC5wmtXEvTwXOdHPtt1rGb+OOVFodyYglL4Fj08Y77EFzlO46TVvF9+
rp+0F9oYLwpL6/E8vwT/h9RauQ0hctmvv4d7Fb7vfZsFz5Co+6i17oa+mMXLd3UByVvBCijQJKX1
5X2bE4+KjzAIVLx5YWEkszJPNZFTh+9HQ/GEkXS9OMVzSRH33U3IhvylIAzkIozC7owub/BMcUk5
/mTgmAKDzvZ8Y2z6P2pAwUIKyRGWjq/jPvGY8DAyRQ57l6l8R08DXV8cj3AEKPuy88+sW5lpafaE
LRLbuiE4ew3LFnQNd6hVR0sA+q2PXEXbED7dEn0L7PAxeynGmvVyoNKujqxSo7U2vYfiEr+I9J72
BFTGH+/tETRdg6SiEB2gk9X08DhA5qaiTCuwxocb/DSOTliUH+1GGC93SU2mWGHkbzOlFtfWAz3K
kZB9AYXAdCn+WWwdogSSY7aNYZ6+H2N8HMMI1sajTrH1LdwS1U5nB7qtmM1IBkzDIBIzSMQOQ5+o
WxpuufUb870fu0fqRqGAmgBnbriAjzmDqD+UekJ5MQ0wHWEh7MImbR2gFtpY9PWZHMy7/6at4/B1
o+qIcCrBkrDZpyWH9r7LcTQtrISHyFraAxZ+LijhrZNpnYnLgqSPx4vGtfD9QUnKN+yhPmAHD3/X
hkLHmcbbG7pesxjWeGc1QJDg8AC0fR+xF+s1q8sogSDTAimYFRKAfNCeoNP+ZxaZMPS1wDlMwQ1A
Qj0L6l+bVUWIozGMrfnmJnlB6xAYl05JoKd0PyDJKsd6lzySlzaiJl8xhbPa2FiHxGgUJNioaw82
HxYtoXSU/6k/OzukkYr3qPItSpy8ZSr0u6FraLA8G3+C1z/ydP6qAMBYH1LfygVJ4t/QnPET92K1
0BmLNWIsJCl8bnF0WiP6a12Ak9TYcru4HlkKfDVucCJEleegBgo9x69H9AtTdzYlWmNhVXdy0eA6
QvsmRKjnt6toeB6eKar0nvJZr+hWB/4Of0z8uZw/1wNt4z59U3beSe/VR17wXsJXkQurvu6hwd2N
C0hjsPS8et7VOXLsoMYJri34+V3neBRWPQofBLgxct3bXLx1l6YnEkvBcBrO3kHzwyiTYMCZRlla
W7Oci+Q/O5Gdz8qj6s+UwFSSac/NDyP1u7UrCET74QH+72+SS96R3Z/lfYqiiTbEQHANHPVXzQM5
QD6fPI3zjy8zNNgocvGJMKPwBUqSQBhBnoIGcwv9TZcxgy26v3OBZZvR4/h5nnMtZPF9JnaORhlV
CgD/5mkQtej2uUiY4sKodN3EKMabYxHwBBBFD3qZ17/ZHVNH1HDrstY+3GT+JjOPOxkHKeaVHlV8
0cPiCzc0lPvKhqOxfm/jnOR+tUd14mNmgmvKHvgRJKLCgsWGIi89JgRC2LxNBbYl8JwiRf8wRwjS
RG3SQlpBHnRfKA4l5kDVJPQbP9SN2olIgmQQSGNXuLvjgE/tk0zDZrn714DhmSosR/xiooiCqDgL
90QNRZKkMwB50f6zauEE/b30FeqxRwQUEND7bekxNFd0NYsApY3BNSk/a5w71nu3R/YScLIcVPsT
PlYiU3rgwXdsZSbmJKg6veE5h+v9zwmrtafOXzVM8Uya7RnGUH8S1wOFXC8BOhCBCNHMGINZrPwU
VuWqj39puSrOdbOp7n/j3YKyy+mMbinMT92wdUo2z6G1OdHRj3EJkDhDoiau9pI4Vl1a0WL+TDML
xrOMwAC4LvV3yElKXcYNVQjAA1h5aGnR3QoLOdBXVHDaDvs6LBLZlXZdmKEybsceGNs8uK9BbdMf
6+AolXf1cp6A9y0WWUPv3nAjEoC9KHAPp4taeCQ8ler+LNdo+d5WzvhtoSkTdlsgt0aYzBb7edly
MwhjfaT1m/2OwOkza5PejBuKJU8iC+EKz9/it+ZSMAc04yLqYDvUMTLL4DcJlbx3Ni3dX3tsrzB8
igU6LY6VIYcmcx8S4wQuQ71m966P1WgY7Gbm1OKCyAJRka3N3PR9dYIfUoL6Fm4HIgxV3kyNja4j
BPwMMFsKEwXmz7xP+tDoLlWGrZIRSuir8JND0U2IwhmpHlEckf96vehFfNjDa7DYqvRRTW4tv6TJ
qJRklA9zvIH2bwHEz7o7rTOPkm/ihkI+brJkxSetZuT4OOe3lKT6EQSKphfkGyipFXhZ6eYTvs7K
Ga7JpwIulsRySccFyP0TmpU1Ca3CXb3PKE4QrAe+oGjBQp55NdxpEW1sV+EVi576xqJ6EIQdAuX1
euMR164u+dkv7KFbSczXKj8r4F0sXizC0FQ245lwZneX+S7gAOu+mONaIGi0oj8HWoIenlSvq/il
kfRyhWsy2xLgAIeWm+IF54C9p+tFTIN84at4OG6fr3vXPRjoebxsfuYkXdcSxPFJJXSyDdoGR9Oi
wRYM/lIVL1ebaOdyK0RnAuMlpSuuUJYqJkvsfaXj1C3j0O4RxEmv4FNLwVFqU8iRoL00uRV3Ch/s
6q7pEt2Ji/m8+FFHeFmTCe3/O55u6Y9NFeZgqLS8MFNEUWrfxW2vuUxHpB+tm/7oliMi7mRvOAPQ
h4XbfaaUlnytu76WHjtPKadYILpAumv6wCxt4kArXQM92JpqO0QLu2gx/NoiLWsEp2+C/f3wgQxT
BG49IuA6BcONuZLi0FqCQghU45t2UuPP59AbCDipOrD/kDyyfLTbVzudoYIZkKnWABukEVculEhb
wP3FFhJk45O16yGGldAkvAmlCeB7jtCOW5nlQFcdN2APnprCqbdSvfjlTMxHeTdX+6pKBW0h45Yf
bS1cnK2e4zvscUn5+tqprKA8q0doK8K+j4BjBXOSQ+Xvv77FN9E83t0XZnKU5KAb1tU+zMLunb7z
lEzz1hnEoqdyl649cfX7ekNpfpdlYmJZSnenrIIC/kRi1bsm717lqrZIoMcPOwVTi1o2IvMkQBW2
MUjZ7GSTFKRnK7k4DBsYoVohGuYmj0LAAdIPVeNwt4NcoB2TsXZYwOZ4PQuSAjq5DisgjIcu2Rn7
NPqDoeie5Kw6pjbWqptNDzIvwFDyanmQRHoewLwdBmoV1sqGrkHxtv/SNplYb6sTbSo9cBI5iiwg
oDeApIG6IRbkaA7LTIAN8Du32heZEwn40Y2R1dHroT1wglDCk3g1n0M24wpH4Luh+JIoZRGyYYOC
x5RprtL4TqNuKleOIbIam/u+4SR3vnqYQUI25oO0Py6/E8Qf+FMRo60LD9nspsRYZylZiNIvMy7p
SZ5RAjrw/Lk+5J10Or9unWYC0mLpM+lpo2T5SxiEYVHRWDFwDbEB9HWez4XBsTqMPyBsqfLyHt9y
0gJB2iNnbWIFzmYnWfY0/jirjmWeXBZkUozRT1uRDQKfTOo/0J4cmpQJPDjfvoLUEnmIdvtgYI6o
ndmhAC9J2cPm1lboIBITgrIVzqJZmoRXhAQ+kbdvP90IiOLMZHUI1MDUXNgXF7qz2K7NTj2QzazA
GWgThnoqg/U4iTpap4F5LF/gwvf/k+4XDM0lRk9TcjJbf6PHh0jDjjf1vEv3Y2IZS1l0898uwtwQ
HtC5xvtco3SfWkrJlSJbocqd/+DC80FO24OCyf4SKdBl1i/Z1QmaLdkai0l4yL55YiBNiNxu5AiF
LABvfObmS3CXZqgH8EgUSpB8TQwRpkAcPN1o43rYMKhk0scV6NSkG3XLYabbfwNDWXUuiCtN8chZ
evMY7WznRUmwe75KRM6C0byMbcnaV7TvJzt7BVHWsEpIoAtfSqCPqTjtNpo2W+bFDVPIu4BFDcpo
eoxirzj+ImYlV81cohlgeg61pOwBGxJuiEUC4IBpdt2HO/YoviuNIjLguINl9EYnigffbH4oV9QK
9FWvSNs4KgYh2Mvmyv2KiWKEwSdw0VLvVHtgmpZRCaI/5A36JDV+TLSWwRwhbefKjJZI8eeQxipW
yBciTfks+JucMROA0UJug7FddEc9Y3+0zRAHURNBkIG77AF8KdybOCl0fWT/rWnr8NSlioWROsj5
Y3nViQZns6daueHf+q/PPrGuum4W8xFLxxysGuZCj3EmJN3p8ROr0XHCc044VSDdZw4T6avTgx/0
F8c+Q2EhTP96Liwo4CDo00BnSKI94MQW6MilyQ8/edYEcMdWQ4hc9yLIz4IoVNUPXJyTT/x6ACxu
61Lu/MsGduVQtJd+3lAFTGn4Bjet/Z06Ayo3JNjzcc+R1epd8P3jyb67g+sCnYkPaKOa2Xz3PPId
OqiT0dL6RfBEJHbvn/oGXM/858jtizmoo3Mhcg2Qnjyxui9NinyC0t61CLHj7RF6IBhYMBNMgIfB
egJHJOPvvwsJbqptPfJlyCmfuZhCtAB51QFHMBgK1I/lhZItXzuiT9KASVlWdwzczR0IhO8NNKnh
TS/2Si2rpk2mEwVrIyTik43EPMSvMEIEqaGnePTgzbQpFxU4JKnchVmNByZhT94wHsIzICRpAC1c
lsjrG9C/6jeE+Fj3iBiyThSPJOv57ZHmCCX7YurFS+OFeLxqLivODp03QO33z1sJaGlOygLHmPSB
D62ezkt7Nmg5a3jYp5q1SSZ/sR/G0EVJD1bwXi1zRtZxvYF7TPetNRMAYyLpKHafhHXaUr9SFPqf
hfS+IMvg/69evw1aJlcH2G/+XnlSWyqMRJM4UDk0Ey40rBLvEQkKHHtsvsKCwCwLx8nB3USAjIrg
VgpXE43IoBIy4UHt0PWJmNa2T2XxSdgp5AIf4OQO+fAZ08apFzS1fQI/FkuAc5lxt015AEHQUdih
Hh1R46Pq4A57W4jDeG1T+LasJhdrm0+s6Zbqq7mBA2gig26atD7WkKjtdepfoyvzifdnBG0wR7j1
WottkF7okXfgm4OlacY9MABBxlDZ4Ft4CbSuryydezDwNIcN9+YWFR+NjyfefzoIUDriE8m5bmqt
Qeb28R/pA8WWQmdSppfuQDqwnehXBYGaOEwmrEstTM5m+wtKc3F2SrUR2OcaTvZLTqSWN39bSRld
ndp+9kOaFStNTtRbi5MtIcZbH42sm0bv8o/7SIz68VZjOoL+RknHzRldK0iMPNZRmN2tEpHFiVIz
lGPNsx/eYgUs9HiO6Obd1jRjHfCTZPop5NgXqctx8E6qIrwc2AJ0PI6mlQq2KbLfUKl2bpBtpmcy
FqiAdj38SudFlW7PIMoDt48cWWfMt7kjDGVjOdRd606H5l7sF+B+uMQuvwZ32kz5qItEWFEaPTfO
QhN6kvEPMxsKO1zbFQmvQY7uy6IVgg2mNkOu7IZzXqcTsuGwM+yr/OaK4aRroMOz374M7oyGjq7G
b8SImLRg7MGEZZGgo9BQpk+3WY0KWNzKMyAf5piZfDrH7IotFzWzeYU6np0SXwL85//3PJfy89vD
8pVJel8rv3axAIa1kfitOzOO3jHFOkwzFA0kfVShqNkAJacskxBSjI6FpjMQzaC9IlNhw/TI+dJY
3fhXllLgWCn4asEy6+VjXcwxJaYgnLWRayJotRj7kjbQUYsZe4kqGQSNL+B/Yi9lVYAVwIPB1u9Y
hras40T/7qCHojYwytRtv791yyl2eG+5SwdTI3edE3XG00STPpi01qaPHS2dcSKbkIe4QXAKx2Bk
rhnzIaixkCmC07y94CGG0gaJrhygZ3no83KqRNlNiPuZll4h4sGFRQC29auGv/IScicowdSUdf9u
g9kKzshd8f4KnUpm4JYt1CCT/09jXZmpe+66qpl7drsezBtuI+1JjofcBDNLm7J7rVVQBAq+UzCt
xUyzoF+WrPFtx9bZXk4QD/t/1hMTlSEQERk16h1juuP2bDDV1pe9eSUhCauJ15/LxLBRyzJRU493
UNUow49FRkeoSXaGvK9U3+SPIQcYm6WntKCuR/0CS5bnudYYLae+vmFKD0ImLg43mZJGxPMRg9wE
4erA01FXImaFELbEaQEE8iSepaiM//WVQyxx1YkVIMiZS+TYNXj42jV+Dn2rU5eFaT8/raoEvhr6
TA/A20AQ+BN0fsZgp5ZFenpUoFPCgF4t0xDv8T1jZL4PlKol3fevfcWgzcvrtrX0aKIsQSr5CxcE
YAF7EiLPVnv1zEHQS/syoMpWFjYkftUdPCKn9VY+m8c0EanKxqAWaYQunazgR/X6uKqDuh4ip2yT
jD+R3pkTDrDeIwk1Ca4pAuUd+/6CB5VS0Rlw20zbBoRjtdt2NSGTTn2rWOxWTAp+Iv7IV9C0ViCR
nx64RYrTNE+MpfTbBxz0iOblviJUhIt89HE1AcG2cDIGVA8gaihCWSKPY0U/5jr6/abgvLRZMYRg
PrRZrL9IiFUV/PuEJHjphH24cVboDzQkHYSdBSTu3ekYnoDheFC39Q0U1l03K3mkKEBOyLPSLWzU
CH2JItemL6moXMpbMxU4bTuf1VrC1TOsGKJjXZgi1ypRc7uTbgRnxAxEziMVeZWj4dvMzUZ1x+oT
mtV4kO5BXBOzXvye3fygmv9dEOx7VVdxIO0+kiZEZhZ9s2juQ1ab3Pp2SjZwcwX5JRj0s0AflpQV
qpAKFwOqIxvSUHL7UQuV1KC0f5YyKWea/FLi9HyhqJn3hZ6VuCSaVZrDd8dRMh2Ncp5PX6qTrMlL
Q+a3nSiUoIe4/iItH1URuBoyG6ZKW+ZKhQZ2mBf12DLgdgvOI9iH1VrRqSY7C0iyMwscR6+BkDYu
xa+mgmlFM6edvazLfMHDOwHY6RErNqzjfkOlelvpCol119gP9qwd8iFDdUv9ANnr4D8JyYUQ1ER6
gRIwbEK42d65+PoU+E/i7pYnlY6/SuttmgHv4mDeiwSsowh1X1U8utGs9qI017fTVE1Zg2IsT0A/
K2Hn7ERDtIwJOuCnfZDrSQtMU3IBALAxj+33kLtbYj0X+gdBWp5UpjlPjzxR7zlkiaWuBkKX1/b4
2el/gEyfTLG28ZYPuFTkT476FODM1CBZ/utOPV9Tr6AvRMlZklzyvkrqmVOKyw67NQB3aee9Suju
vcwqLmErnAJEvpOjGLFzeqnxKSGqCmfEpmEgvTgyZUKsr9q1FbX4SMVIUfhoNiZqnzR7FjWc6MOw
NCxj0qzEK/25LfWHmWEranj/pRZGQZ/7PYerSjx1eHJiNbDncFNbBclbMgK1hu6JSnmsAh+mR5p0
4r1SwtXMTSsaVemW1rT0xwtEqe73nJ2R2XatyCQn5kaPmdI0igVpdEMvjAUQSVZJ2Axuyqtn1ESL
TXR/oHTOhZV1yADhzspESUMtclC/fmmd0mrTkS5mfKxhGl6v9OScrzQNl/iQldU/5te3Imy/Of8H
5jPW7uoSQzbenk5TUqoigMBrIZxeKO9yFDfT/l3G3Ps4f8brXE1JFLBXE+OHA9d8TF7sAnGkjG9p
FC7EvSMHha57zWBsb5+fxsTVxuU4zXNL4iHqBcaTsNiVL5W/e3r4niI2Oikeq9ywIkoWwX0EcBzA
11OxXXS2s6+f0AYAFOyn5I8g41eNzm+eJXkRTr2P1RsX5kMvDYeM87IIP1KemhMSHKLIAoHNBmGQ
S33GZcL6FiATvNLU0OCBnOyLgRPRy5OyPY6n+a415wIf1FHNifG4YuZWP8iafusKV63ixE0BfoMr
F0eaQOK+OF8JEx5IwvFRJbktdoEJsAQePoYRrsZn/vGCmKfAAhNBW0C/XXNBk3I9YUjrovUklP2N
6n+S2qoCBZ3NLq3QKFuxHzuZfuR9aLz4IJBQQL1CAufmklFAIe/GSoadjMOvYxwcXBS+c5zJjxA+
as4Le9WyOuzR/OnTCpGHXJX6teAlO0595zUvS8UYtvqGjGDUimjL7mDKaZ6b63gUFHzvb/5t9oXt
TQCXn3QKo1hGjQJWkMxkfAr0nDKQWJu/0ly13g1Z7cDh3pY3j0IuR0if41XDLJWtoxZxp4gqT3ci
JGx2xrevk8e6Kdl5s1xOFTi6vDQZcdrx/cphMWq4ULpSANy3/qvyt/G95GizMwPl2IlXvkgvdeB6
GI0O1Mjj9r3Csc3KLKTTeuLz4FIjbUguzuZvpO975t/CttGKPISLBfJA/3OWAkBjHzTOxGRJoIzq
x4+Zd0HABXU/Yr2KbFfJC0u4j7/b3wP/SHRIr1knlikLO7JJvPR5u6KPiUxkvtAmsazLlOFu4Shj
5xLmbPdDG566YdEGQy19RMe9EHcFDvtKRsTYkBXD0u4Wx+QzXiR+R9CKoUFUpVMK6rE4CkT0C0S6
JxPGWHXqFYUBhCdrVoZ9nCMHNfWO8tXDcwl+fJ3GjygwtkYImrR+bFC0bDKKMrQiVBFhIHlxcBkf
Ss3f2OLagVoqnab+UWZUqWtvoXXytaj7XSy6n1PkR4xfa1Rkdv4b8y1sliW/unG3TpxG2xohgx6v
zJIMf4vGTCtPDvZNZC3/vb9uHtlz0pH54dT8rog2AcySd12WbXzkrg43zgVMe+4EiJRPQWpQ9ypz
0YSzxW9D2szvioDfXRjGUwvsk0ibqWPuDAavfyFjAiygEw4T2U3On7GzkV/ziJp+0JR8hAtJSrYt
213/7unBwbeoxriiLRjrUZSxZUNkZh58Z/CAed0ysbtz1smZWJiYpVqBIR3tdaaClj0FpCJqbT9X
XBp5+GaVvPm1Ra0MBrCDTSr4Vczdbl5cCIFePc0/qGG/PX3+4uvYN0rOVNCrr3aiR2U/GJscoZCv
HU+Ieg/+1EEE7wgFsvJZ6jkbLcaMiM3ABfMLtf4bPbYmviSB9OFUosfBdQQ0c/eDsb185s7oFPh3
l9nIWWcoEOzDK/dMfhG4NaE9r+cQ7khN1Le1FO5mEA7Yh/8mWbmsqyZnYJUA8dadG8W308CGeR1t
Ml2TLMK+Qf5pIJB7dzs2Tm/djVcYOMmAw1tLap+CHt2LVq+Ju8grLGyJ9QxHuIspn3vMWkdFJJru
c7jd/dmcwqw0JoUC8oAVZVroK2lRdsfnVPZUuIMsb6XmpLDbKVCmfolZlT920kppr2U6W6gcxMRc
bila8mkgTkiOqT7Trz9mD0XiPuhXkt8ciJeZYUjaYR2UolJPoj0DiW2YCKUhDxnGARxEwwOALQrM
XcOojAULc/9pulaXTH+enpWeCv/FTEyKGB4HMHKObUvZrCAw/5HD3S2ozwgWtV3OrPxmrbq5H0pD
TzC9Rbi7EAAa2FjHco8bK+3bZr7FbExohUv5XshgrNTYMVuc2vJk9/ZPTZeNvJf7CGWrg7S17hYH
jGkuZrG/TF8/194m0abpmrKIOs6bm7Utq5B1gMdYnBB5mvgQ6DhTJlPqgZYgWLHbehXliNGWGboi
i696vrIIvrDkw0jLYKsL6b44zpHdTg1GSKqqh31H4YskwsSkwxhZ93e9GEiQhpu9Sp8vtm96HAvz
CzUdjML2GpUoVwpxpFCsU6Et1UYxCHJy/bAYVU48MCycttwXSHAGk5wxF3RYAM/9J5YDM0zbPHwa
OfRgOnfnSgw177II47OrnDHQ3hTkfThAEfBnVNgncdOlDYKYGAmYujh/LCxBzEOn0O/mnjJ/ulGO
Qu1OBKm4zgxfFoUXbd/2N5bHNI4QQKN+wjZXDLpbO0ZODIsq7rZQNxvLHD8GhlNKgPGp8OhxE5nz
nOE+WabgiCyZe5mzaHcqJ4UOmsHqfKMtbkULQQV7UxexThnOK00iT/MwyfqUs7jPRehFcBdd+Erl
WYET0jy8aSkExuwTea3qY4NDcG/8t7I3uUE8cRkn5z5JNrjc36No0HykhA4QAGUkhQK0PnqJpFNa
Eyk+/dbB1POl+niSJcOqVMi1ghHaxHyucX0xM0flp4CzcDXVwoiIPKyqtTwC0nUg7GonKshQ/8io
IrAIADk7X/6WOs7PEu9lCWGp6VHBzhbDvlEZ9sWNKwScW1GUdZsx9qJDI0ZCKHro6H+NILBfpDz5
nGhX6l5vsCAGYRCb9YnDoOqWMxJkArBseBOqq5BUGNiW9u1wMwq0JzfWVdYLilrK+5UkIsYLy3vP
Bth6vg8t3RX+NYMACEAflJrTPpPRtWplsFnpN+pYULrbhVccAGRl+1yjBSWBdVFV8KQQktbs+GKQ
BCIaB5vwcpR4zw37b5e4dGq6lyXLMahpFpFa4lhTy8Fp6AWDshSiURlv3Mr1h+b5FlwDeUINTWny
Upn3mFAKKKthAw6g6r48zrNK+109Y5kWNXEpActGK+q5KBVnpU7yoSuWm2744FUrQp7+1YfsKMXC
EQRPudh0erYAYDPUcTykvH1v5rmIiZAcklypMYiBjw3OneP0qrpUHUSAhRULU+ukxGzyImGewRe4
bRlMIcQrkgExr2l8ZwuDbocA3h1A3wgWHZW7Jnez2jRpGU9/xgmvvNaXnY9rRPt5Najfv4BU9Ua7
ce4Sp/5SQ43X6B0XoHEkpDRKUvqnVqootXTi9bdWi/gGIsDY24QZKYI0X8CRjyTYJjA/0jHzpFwv
rQhrfuKIt/n52tDUypjCwIDB0TD1WfT5Spm9XafM2rDYfTmr0kKEEiQzOFM1/+rhO6ezLUTTIvd/
rLfYNP3a8eOp9bBHdUEtsSFQONI74NZW3Cp3E4zD1IJMdGf4AONckfhIqo/hdOujIZeJWvyLdD08
jKJFOdxeL3DNC4845qM9gGxZtrDnDxym2Yo0hOBNveY28rhpp4PmeSDifY0naNVOAXXjDC+tSoom
ZBFJMRCasJb4MKsD3nySmJPQHLCQDJKXYIwkRsK6lL/yOYVw9ssTaA0a42yuvUjnCwfjZ82Xm5qH
8zAT45CtLK7+cQa7jZE4UoILaMj3MPfw/nSUMcBv4FyRfkXHGG540yPw8hl1VJQBOfXCB468rZct
CWWR1vUsEqduftMMkDPYKu1ilcJHnB1niEzxsVo7Ltifk1llxbz4d3h8/pQC7cnrVx26zOMYseZh
K2J7JdAiLXBA6ZnLzMqqJ4Vy9StvgVW3eFlKIVpAHmb4Hnnyw4YM3RF3YE/tFaSgDa9y1SGbP2Vv
3HICROgn62V1/tPqSAtv6sCU2EKQmuIK7XLUYdKNj0QYcBHXXMzgZ3T/Cdl3ZwIPZ75KZkPTiiRu
/+z/9N96m6HuVHPueIp8g61qp3+vf7GEP6Im2AV+Va1gIGPirBwv7dFvfovyFOL+FHiQC8vjVsV2
3Iw9vojCCce9PCeXomH+TYUS9diIofcWcdUJXSxXhclbcRV9jwjr2Y1LHXLwNssl2WsQMOUE7IvU
yBpYMwycJsG+4rpN8h9ibrc1PMrgMxNk/HYIjRu4bGNR6tjKWfPFXEJqOUXAmPCoYq/aP4WKQ4yC
4I0Xt9bRKOq0jANXWagZdkP7Sl8+ewqlvseVVu/+efh8TcRqUVMrm4f6v7Sy45YdVCuqwAs022Fr
/4Ek3QLBg5IHZEkpwvrtEbPK2vmvBCY3d5TlQNbB7Kga6CEgDyRBj6Kjzws4aebgqWL/2+o1c6Rn
ntxm9NZ7i8a8SfW47qf28kgKbakihOl4UYtTwO9UQ+rAQhlJ4ws+aSJvs5q9dCBTd8i6dBho0pdS
xejvZlGG1vvDqbUdt7Qv0kDhB8Bq1RDaXNMIcuQx9wV4N1j0egdXrx98w7gVyhm0Lj+YjoKt7nD3
3Zc1dB9qGSw4pud1Q1d8BAZr9DwpMJ3/TJHG/1tFW6mwMsdwYXKHXyMK9k1xU/Xu41c/YT6MDx8F
Pxsy3kHPArr1wjVmzj4ofZx0PPYtHuFVRfdAXStzczXLTPQQu2uIkOM1tI/ac/lXjouGrSWoYSCZ
W6tkUzHQMmFtULQWoo9ylCZl/Olt5GtEblVzODmVLnAyQ8/8SdyulaV0hGsFEEQwEPknCdWrmKbC
kCyqvilbHFPjY0BeLWDt1vOPz936xCvGXNQ1+bdFHBvORhq07hC842D3Xf1o+yx+icelK1azgY49
f8PHYO1CMh4dc3TnntkmxLVnBUZaWBmlgcciVy/ZYu+8gahiWSzZAH6mcPunWXf5yeFxPrlncdM+
ZJdsB6tXbEitRhTv3Jzfc8HgT+CqAAEqJyRoNz7RXjzPAbP+yBsBcXYXmUe5GDrUDAs0SUsQzTtx
8UnEXFo2riIboi2HHqFlu9qtqq6FkyDsySJdmoFqmWddVU+ZUfbPcnxcqlFo+kleGSmpmmSsgV5i
9BUIvOl9k1Uis4TrsjCH2wOZgJu+xuKnwzEadm0m5fyNwsZUwpmswCbecKFat9/kn1zQOMI/bYKP
a2AG+iGgkjr6czGNX5xuvprbUEB34mVx5I8eVyo2VWcGuHmNsnBbSlFxgjPW8krFzNQUglI8tUKu
qbRD+sJ7NZn0f4BqyxPbzsgKoFVzKVChg9P4IZXjYxC+XCQUqxV1yxKRspE+TcdaoTCjwqEZ2+HK
+yIdAiMiMGk1/7G28zwR4UrEONhMjxFbq+CDc/nscGWMl3W/jhebeN1PjCeRAfVmyCbVj2IxS0az
NJ6HiZn32rVPYKwLTzyKmRl2CC5YbarRsApym07cs2e8LTvE8TKNwCpi8MdZoWBS/eotSJBri4TD
eJkbUXQemhpj8V0uasFBoLOv9Q4vi8+QVI0fy7s/GvQ9fnjhHdmIaIpc2fii5xg1diYRdZL/3B9F
XT+EnKWRJudorAjCLhLOeopq1JvfVP0Mln0isubQdjpH5EPYdY6NKS9x+i2JLGGZqHZnNcT62527
VPkjRn4fA3OlxcISldZSlrlein07lDVLGxojNxkj2hesh+hy3K8uP84RKfKd22yUY7RvgOHoSWT9
IpeQWoqWBJoIAA0BIU8PkIDppFYIA4SHdKRfNGKRwjkKw4ZO9OCZaGCPdYyx/cE2lExiuUlcoZJq
uWzrK+kIj5p+TCfGmbiVt/FfvY8bZYh1IjdrCHL5BVTBxD5vOtamV/Mo+8xTNhWdH88UVn3xHH9D
ftfCv49apNUUEqzIAu291ShNKcwduBETOv4LGWSMxyG2EPxNpkyB+GnTQvY/amYp6cF2f7eH8zD6
8qVHcjOc137hh8TvpGEFqjsXw9b5KlQtgjTp8aoOaf4F5l1Hc3bBl9+Y+vCGVUkWYh1VnR8Tj+lG
x76c/Zk9eGNMN5SliuF5QYHIaqqh0xmI7zN/PlRsmKxJg2v+HDa4cS7dPKPUjszrQz49X98ONKM5
O1tv/2GIxkDsEBjKF1pJdh3q0R+w049XOLbHPDNlbfJ6cJpXiGpz27IVLyQf5bCOqmtjpH6yCgqT
EYF+w9h/qe5fyUwQPFe65xPDSJjBCtmK8+xeNc2csAUtayImG6iTgMTcVrLLxV5vqgg+W0qy13ok
efhOUDw13bBFM2i+RcvnzWV3r49sOczsR2kv40nK5ZXCX4SsKMom16rvzvaJSbvznzuXAtkzLTRW
axbBlM5Uky5RUAoKxDg1huRhdd/A2K/ZSR2JKGf1Sj15xs5eUm5+ReOUZO2Eu3GpyFZ5K4HlNiS6
cnXDdKzJpy2BYe/5kKXWK39tS5zClSMXY31eGSpDecNsG+KJXNJGH5yRdMuhpoNZVaikroc+IWgK
+3w6HJNoUgFI/O/17WfUu2EOjrXHzzCTTb453Q7NxW0mRlFAdOSXdZskhdxYYKJpJ4m47wTfUqI9
BrX4PuxptPHyVgPt3OPZCkzr5Moyx7RcGeTzdhD7zVlADrcP+JFzpczj5ucA7iXS/gO1pH1xGORk
xygxheVPAH7+mOUYwwJ9silv+bVOwQ1kja5tYkfOh4zbeTP8XCfDEAzmyEmjeNCEVPtNmI2bsErh
vKyYv09RZlKc4qp+MZom1H79nqmojWUHXuoEPLMgtqfodZdKNPSi2zHqmZk5ml662J2vOYLSRemk
WxSjAdeNqLPQmNj3HsEcGxAURaswBwLp3En67Gjd2l2mhGwr5aKb3mhhAtKhyx7/rJT7AX0MJcau
iHzV8qNsrFeJw3gqjUmegg6Am0M7PnlWE17nyd8X58ptxqtk1iD1hwXvfBPVHJv2MrmmLmVr1+pN
HbHLMF93JnO1v6xVcI5UiMst5fhMgCS/u7LkTLh8d2MBYJKNcgF3NGn9VgMC+BwDFoGHrOmVf9x1
Gcy1uHlF1mka6T9m1Nhj8KiPxqWXEv+WffysTT98ivaISFwS/bZAyUXGhy2nVJu9sBvLruNeSOeS
O8NDAPscivKHWLLi0JLJPHZ1FIjy1jACQjfBk8Wp7wUy+r1E+hpwdl+8s1aNQA2rgIV5emOXaJ5K
kCuCBiouso9FmrGfjllINlZnXxU92nk8fIRJ7OkcHbDYJQTL7CPrkwqr8hTxlGIwe5UWVoqu6NTQ
5XclMJttQiLM/RDasDgOwbFpRv3XY1ZbOEDBcCnQGjOpusedw5MCu1d7Hzq2bKdmavzUSggbNx3w
747rFTwJmrkntT7mvj6KnFIUi4gl8J1Gw5H/9BbwCuYeFNrWy3QA4J9RQ/CFzpDaxRqJRr+NMl+g
J3dC4+JsJDxVxrfVORdoyAjHoXQC3zyq2U+gYVjJRf62VD6OsLbRoZ9a8IqCus+8DJ2LWk14H/g2
ehQ08Eg8lVXGtG6TD/1KuGBAKyxMBDPLrxHxNQYKhbmsn2f4Gr43EHk8/BKMyzfuugIfWpRd+0Rq
teHemxyCKV+9hytPDsRVMAPP8qk67fMuAmBbQVEooIQX7b+RvqL91fehl4Y/izyYlg+Ku7Wa7jml
gKIBvHIyjHdB26ZWVjmeB2WeJeqpInlr5VDJD6rCvv7iU9LY86v9omFxWb92u8BmoXZzgKh9Ydvs
ozgWzpyWWTvX+rw2crdvv0PkaJLvP4DJ86UTNhKlhKhpfd7B01iZKm1b4NS05bLhdxSnYCe6R1JT
3XGoOIIZdyWDIE2xVBZYyr0Wk9ojuS1AImIyNKtYLL/prG03QDKe1BDXgJttkupTmmhRwcoYD1tq
JqJj0iuNzuc/gC2iP8cUsbJ22gb5Gww1wb619HHveFgYW62LhZnKnbQSU7KpNtGIHxvLl2veB6D8
AWCmvMmvyF2uAmBkB6jGGYAmHThKex98oivtiikk9HHGZ1NLz8hjEAcM80/Qe2cKZwixQmsk+U4V
pNrh3XREmoJ0VKWwQcGrox60ZHhHcHpTvkLxUOa6NHStThUALUse0d/pdLM3BMTCvTs+lTFqnP8n
dF03XrbyKZrI2QvpYpVv7mkJ8L8oiYyF24vsARxJnEpAqXnysJl6056ydIA1j1qIsg0vTSZGswt7
HjgHOZOhZc4E2whqkgS3wBYofx/PtkPhF7eT7xdtb+3p0gg6qPpAD5wMqTQ6kYgZtLOEP0tQBFqt
zeCBFjaz1lNi+f5J2OpqiWbh9gPBamTIsm9qTpkoQLPxstUPbMhDl0XTGAhKt4TprXWTXCaggmkL
pxjkImgvmQ1EQnRTYWSbsmz6i4Bn2oAXmmO15RcMY03ZjhA4AGj9RGAcCS3Mdu0UGJw6th4bibMN
fSqfQb65qT92PKqTc+b+H9gweJesIoaX+VZM3mACeyWXRnUB9pUJdo83e3ArAKTXaRLaD259SrjT
4Sx8ctomGb3HYs4u5jTiz5+AS5Tm91oZIwqVtQ6UssR0RrOaoq824xTuzUs2byrYwtXIchABe5e2
YD6HfAfahXPtXvvqZhryoRT4snmYksl2nyzvDaCzQB0OOshTzJn79YwaDpppfUYk5LL5EUCRZ9/M
alnnJaaOf+0Og63jrGY73Wxgtu/aNVI9lDRHu2ot0QBxLXnNpSIll5ltIFtuqeqOleqB2b5xGciY
9AqylOxR4mvBw9jqXsSuFcSJBo+huJlaB507yu95s7n0w+tFBSNpP40H03wiLCevjnufePO3YOpe
NZ9mlG8fXLHprQ/fqufFlAgLUR8F7OAWwGDRwXFmYNS6IVm3G32PlEJ8mD79gdyM9DBETKQttqoe
ZLbK/Vmm8yWc7keJ/9+p0NzKfRrVKjek+BCoOwk7ZedgNoPVtXTqxTEr4pFzS35sa9oD1dayDsqG
gcQ+HkC0VFX0ij9aPSkdqq+lOy0WmrDcmPGpCHBEFrbCDwH5fi2lMG+JW4P9z8hQ73cKWA0VUWNY
C2P+Bm2FPWLETlx7LOHiaS6BR8GkWaUFgVaAFQA/nMsHUAoWDbCDrwI2y/EGUnKg0cLMzD0wbVjz
V28Ey8L51ak6esAI3sOBieRkkjVtcNz3py53tXAri/MF2hGFKQWkW1PEt6pyGzIXKsv21HsRL2dv
5HjPP6ggVvHvpmSRDiKkvtFI9NA1t9LF8pqF6JXMNv1QooWmy1ZgiuGejmx1Gj31zFYtohu37ZKB
06YPaRiJjQCBf6g+D7YVoOsXzEutB1gn7C6VNdgy7ni5gPCapFqQ7Nz8Thd6pVMoTM7yG+9rG2t7
2I7pB64YpLmZyoP2fFQCjD+TFkMzgOmTX8scg8O/HTLqvQEJiaIbTt5/vFYEpaSOnatsD84+4KeP
n38LpukNA2tsgd1kiLKMZICGlfq2NDT4QSN8FfHonCSzU+7rSHR1kQ5B11bXmFDWYGvrpZwbCfAC
+iSKT+FqBPkLHpvQFdptZbqbpB90J12LXl2D0mYWnItMj0dQYADeHLxwJKPLnpQFzyO3OQ2Lzme0
GPA6+G+wQiVg5Fou8sCF6VcN8+tX6KiFhWhyVFTO1ZskznfUQ3QgPqzbrGNxIrwmyIB4MxCLy463
QlvD8esyYvBM9Auf/tgy6jZ/i3oSXu8mG1nX7ekTODJVdIYL4nJ39iu6MtcnCxWdBwlVaEeoF+Yo
tIt4yB67GWqACOXFUTueUFcSBMERIZF2y48pi3mGdbuecjXdWvKSC4Vl5bGRSEwuqtr8mnJw8RS5
Ez5zg66q9QwteTQ8R76B+Lclm21doR/NOxQyvqSnVu+MDE9MNGTJxXv04PA95Fvwl5ZF2TCxFPC5
CHISqNX7O3vMcydoiELkptikYF/ZQdHVMQSd9Y84Ea/iIzbxVlmU3NAvrUfAhafU0F5npGpGq7EZ
KIOSgfGaem2B9MJtwnbbOZ7u7jP2CvC4RW//YyhDXWN1RB+5Q8tyZbSroRhVsxij3nhxqlz5C0SV
5em/UtT1J8z/8nNmatEN01o9UMA4MS/zJipvRMmaXGYkXua+8Pmd9aCzFWvsa1EGSAjyo0dZIvtj
YqpBL4yuQCcjuDIM1DSBeAST3xffbRLjjLkmpUJlsej3cI8at8lDAIy7WrNtoQtaBH1I673zi/U1
FeyB3FEB9HLS+LFzAA82qHXZNfd6WhHgCjZvZ6weE9tfkqC8FmV2FO253izXypnRpaf5HvKwSLtT
x0pSb42r6wlwNIJZOAUd6gOtLX/CjUaINZOYABjAuRGadef++DwTl6HO5631pGyzIEJDWCt0k2qS
xk89FM+4CllskQDTOdSuk83D8gdx36XG4Z03y/cwyw8QZT6VwntjJN8quYILmYjO4chE+BkUlnSY
In2HNltYMDPPCtlyjmc1+Z5PW+48Q8qT1eKVLILIzPr3qTHXaYBecGe2pm5rT2K209dw2QuPZkzP
hdu3nqIxjWvPlPkkPEqbULnzHJRBZQMIdJfHQoCfyis1GRNl4hWsXCCT7dVm9AAjzgNF0Tkz/JfH
BoMI195gCXITzAX2uw/uOE2u6I9XdHp0lfwPQdjt9vxiqXKM7H/sUZUk2GkziwqXb+cMiYuTWzvW
9pdrV6i/0FsC2Nw31blnz18VBpWt0wCq1/2DA6OPoHYVEtXvuZLrhUxDlKg83q1pEfVkq95ikW1f
Xr27SlXJI8hLInoZj4RTqmLLT8SlcGJokRORfI4QnR2msip3Yx++VZuzCkc27OfLjjDpD28s5gQd
r1NDAof6qVT5/rwTwT0mgR/Z2sHX8NrZ8CgZ2jsNWslcZX9NHpeabLAssboTXALSz+5TR7pc77XN
lu2MkCAMJ0vSvKmgJdn74Jk+5vkQtmng7Mw2zEQWMJMKtRfxhy9GcF4bwbmM95oMPL7S2L9O+YY9
jGbtzX3PIIksXR/QosftwAZ581rylZOOCmQfJ6I3RrFs8iLEqBKvjs7Ow9fCYav/n8QMNkqJrhFb
mzmD/D7pNWF9djf39YQ1VETa6QfSUxU6ClPrj18kylqdvNhgo3mmJNt3UGtGuRyLSxc0enqW5Uzt
JsWnxT1W9IkuMD1HFMzohxm91cB3oomgk+FqQ0pfFzqka+dzJZYKFWnLYfRaztXJ/99IEuulr24y
II3lKyMQLd0KrgyP1ZxfFVCV0KM24TLl5mFvad/zOwy2OAIMbvaFpZnPei3D2ObJF9YMVqjo3jCD
Ijasn4k963FDHlrlQatsfxOGBI7mPuSS5ps5r/fvvuvMOSvQ44HIitCpaNmzyNQknKupO/rCM6yf
ASZt6BeAz5v2gmpjaT7HleTZxNZUs77mgunMU1uPiLiVwAQuiGXrin9Nxo7kbfBuU+NLOpDHkEuC
v8x6zG5QnIaajSotk0+gOyNz9IOgUWHXSfRopyUle5KEjherU/s7y/uw/WclW6oQDrk//0NN2xXH
Svomuvwa/gP0aGsHJQhqADcEcn6ukdTK/y/vCJyimFg2pAI65CnsYaUfI4T7IWpVI0YBPmwZVZuN
TZzrCRQVL2MruEKm5PLxgcIuZ+8HfXNQXDIEXiAUp0T+C8Z92b9BsqCcmcxwswag2vlOkqjjz/I9
zo2/Ji8K76nbfHeSg0k9kVfDUaUTe179veU/97yS+MSYUH9Uy3hCN0WbuyBfMctMgUXdLYpiyyoZ
7b28vc5hYczhqdrK6ZjEG7bPF5fkj6MSHkIVfIGx4PzKiwsdjIN9yCAInVuF0clrKUqG47tp9N7h
DZmX4m+zFgsRC+c9Ul6Sh0JOmaVFqRN+q6lzqGLFcFqPu8i0ZL7OFUHK72ep/DyD+tFfpBePb7AN
G2k1WqjyucJIu/sZ0IIECnt38vigwaHmNaxXEFSg4Ug7HtqHxSJr5SlsvIYH5HPelr46ZbfpXgGD
Ixk64s8EB5HScRGK5k/h5JmcsFKewzW6HSilrzE/VnVfY2WbBCGd+5HbxEi2DTQamkemvAyeaWqE
5FNpRXmUSCUff1gFMfQb/efKhJ5zKUgPL9ijZrAt13sztpD38YqYFr2wZP6xllORjz40HxURhfrZ
6l4Ol58Mvbvui3YIQdCVEGR0Ej6FbEuBgL8awKn0OEw8dWxzdlJKvlGwR09bBDVx0tIQuKadhuJS
dqNqO39z2Ltip9HNEvhODkA/OnFrFLk1oN8pT1bzujhqGdTHUIAS925PEMnlh66pnUcyJr7rYZ7f
/VmeYjQCUjwwur4Bgt6BbezmU74mQVy+1x941yH3ctQzG/13uU0BD4jfKsxXzp0A95K4iYCzSjcX
ONYqbSTs4NYAVsCRPu+tzsm0+sy26w07WVoZpciyUxOjNauTssuWEa6y5mzMug40THwAHmrGKIm7
iX2J7G9GOEkS4JZtxjVdHE1C0yLT4VudrsK43eS2zmGaIUBimqu3vUCvBqtyCLoOM7TB27z6CP7T
iq6rFzjPAd/w5HftOe8Wq1CVgIo6HwT9fnJn5yMO8D+R2vstGvPJHJurjmaCPMyymBuX8bsxjNVq
R7Jf4Bv2DDJ3QLRI11fsm1k1oQmNfpLQfjFdrWQeKa3DJdIp3na4omBW5BNjrT/e0ZkykKysX6Do
h9dSqD05Mj+Lf93SDtB39PNLI5bCodKvLq3gCu9BCstXTNzWkgeGjiU+hajTODaSE35f+83kfBp0
aeog9pB2SVLKnmt1S1fXYF261tOCGN3BKrDEQCGnJaXLdiPNFMa4TYOwLkFd3fdYmcX6WlEC3bpG
BAIJIGEaxXCLLYLltxb30ZTfk/aIcL3x/2OmCscPbA6x3lWSi3Cif7IlI0HZG2eIP9Rw05mGzGZx
eP6fghlDLWPE0j6WMGEPW0CMaltSlHC8hG9/iy3OkAGR+rkJIxvIG8kBFQSegwTU2MU8PHQMsHgc
ntFDvh4bzC4igGp9rIJi3Dxi3DLGzP6h6Jo/FoyPwPP67nJm6UTZEscLyMrvtmHPDrb+JE3xq2+K
uBBQhhd6y+oGL1Cit7g3rDkc/I+Rqfs6DLyaEIZafFXM0aU8t/PYqwy7WZSAwVC0nTSkNI3MhVZW
iP0cCyLo+xbUskeC+kXkZpMo/mFhmHeHVxo740jGEVikYMv+So1EvP4gPo29uNhitcW4g18VKUCt
rVNxwEUzGSq62kM5g4PPIP44xDQK9RSopUTYLZAHcOh3aPRWmfCptYgAeGEnqemy2KOWdhCoik8A
DDuy+GAEo+44jBD4Fsh1yFYO2fYUlzHOfNrNkoKlc5+mz+Zjod7sgrqvN3Nm6oBL/T4FAzq2Pn81
A/sUVPB4Blv4whNvM99pQkVvIQuPJdB6hv8riCOIZyFYT0iiq8OoEv6qYOiYfEwEt2wz26YneK2c
HuqINuxgDzXC2XKv59V51ZKreZlj0Dq6a7btaeMwYbETWBPfhBEbKAa8vZjq5FL1c/3yzuVdprFN
jhRFIIAgA5skRjo9pO3JTJ+YHbm+5AG+ipfqlWmohQYoWr13RNu0wYMPrh8MyFbKzyg3DR/HFWeG
YzHiKUX6zJjSJAKYQFepfsI3xvT2+59bbQ4xbTbzU0xcZQDd/j9IH2e8znCzHAxGLH6wvnufD8RE
6Bt2j3loiT+xyuL2qvLAjdwfCnDoRgpuXIEfkDPNOStco0K5cfiLSqKnG3AX3ce3uF+DYUlskQdw
3z8rAVbwP7XC7X4bONe8f9PHo/zkqCH4Ii+4qDm4D4/HV+6PB3zqxMWVF2TZ9L9pNmGXGpT3gFfW
O82/+yFv1ptCBzS6F0j2qxwJk56lsTbqrJorWfsn5N2n1Ves8dfRDsOxUABVZVbi4i5AG8G+qAXv
ubrOpcUm0bxEt+BmSRUzGq1X83DCGksWPj1c0jOv+tHvfZz+L01fSYS7X7t/pSu09t2pa3GkFXVF
Vd573QL3WSIca5GcHRXarjDDPciMyaO5LU630BWv04+gfj7G+hmmCatprzCuB6BRkS+QXcpmpA2V
oQRMhJffSkZet2sim9gLUKy1EUzYyTjvqoNqkFkhxQd08gDouVQeGFEErS5PVZ+u5awXKSKVcMPX
5k6rpSRsZ96C1FbZyMp/VJqJwD1eH3MKLrBd6KfM8f9khlNRxaoBus/3p8m1XsVio/WRUkSuBRBy
M9KxLcoyV4dm8I0wa8ic3qxoUsQi5kXLPltgD2ASA1lewbt72pE3TVWsTAwATVFqdDm/C23xLgWu
c6/QsyWqip6J98ByqVKTvWoRSRYXBxLH7aauHdBGYD4RpuiMJOrinzIT6lcZT/YGCLBCI9NwvwYM
5QiOPD1tQpbTapqGQnUOgWhuIEwfkXHsngx9sjrJ2iIDB49qQvAg09+RHd1gZlJ0bKAJa3Bl1C8x
1S14HbWaIykTH7SHVmSs+hXK44EwOBHg1012PXhHW2CthKk3KxRhcrFRXgblK4Mt+DeY+sNjELRA
hWIlFKHbEXcF5YcDK7ggKckWjp7vP7sKqYFo6fgcbdroidlDh+4EgPAKzamIFR6wrgW794FNbnCc
YAOazqgXzeerjaa2uHk9RKlAxIg3D4ksOm19wbZt+oRa3bEw6aAeJfCpYe3k0AJQWJ6xytOaJ2jp
DHbln5LV1Uo5dC5SaPY2+WgtoHnTmoP1e1MnEAVAnhsqz+uBb+TM0VkMA9syb56+nmKOGTbCh6JY
11vAsM1XWDZeG/w2i3u8BorHh6sOEwSGcnY2/ysWzd8PUZcVC2KdQB/CTejiJCZUWeNrVPUX2Gfz
IeyLyz5+vWbZIqbm+a+oVNYRxRjBvQqBTfPtMYHag2w14cdWpe7uk3ZEgdy1s3XMUQh1yOTxpPD+
ubW7RQBhIaSjFLfEFRufQimB5ogkCk2M8p7/13247WixOliwscuiylo/nyuzWlg1hnDI9LVFe6L1
5t3TZtnATcKL82jxNzaF50VyTGSLHlPOMm84edy1BG3MDPf7pR7ynBQec38zgIEIxd8lvWWjfZgG
ZWohyQO0G2MBgEksBo3o1mVrmuunTBc7VnmFjb6+FJ56Ykkj0TG8xmBWgHbku9RFtSdqmbFBHqPP
Sj5KlBNYlPbsC6bj5XEaF+mdb6WmZE3+3neWEYSA9w7qjke8ODiqZs4SIEbvXecpHnWqSOPALVQN
Eu35cWMfClD1njx15V2zxtCqIUlBIdvkbh+W3YHNQCtd1ixMJcAYxK6a/FSh6vmWVUeaAsK2+9F6
I7gzVGj3YjTxPIzS+AqPEL1JDqbgqWDTEHFbvwzg/HJ2PTm2o2aZprcBGVZa63cfNHzph8lh3n+z
VDcjPVXnFY9grlPtKr3druICgRlVuK75kCqqaxEROvp65cascgoQ01wcvQzjpBqS+6Xvw/gEvXRH
KeaSCIiANAYCy0SnoSbSmN1XdhfzOcqHU4PsI9+qvco2gUyj2Zp2XzAvmZl3DGP72oO9khv5/uPZ
99YCDZDmXi1G19OaQxebc1Zkfco24ehv7cXhAahvQtwHFsWcTOIGK6Sa5VjaTtv9zYIht8UjOOIb
bHhfrENR8UV4o3lNtOvjiIBVXG0oKKSE9SReCrGOpEIJ6uBkD7Zp9obkaMtjNjZW736iGng5Tkvy
FO1C7HevWTyHfy2VWpbdIa8rt/74js//VkzyKDjhZCKTxfoQBuS1ZuRUzlKBNJGrIFeqt4xvH5Gy
r8Y1Yn8FdeWYE1pCQx4zIgoq1Nr0vhYhUtunD+5PxyCPPHarTHSodn/4YRBu/nb3RP6M+3PKhHCp
DrzYQBqaEiAYuhE96SxuSRW05rjVZ90pQRfZR8N+oTpssYoI9rWHeuzHWp2fKY5b3JRXRcpruC5q
j3w4m3BAXel7bYT9k0jRBZY5U9xByIeDNzdMrqPCX0Q//IOfH2c8ydJMmhge8OfkfVHgK0JqhVR7
gozv68U8l491CWA96Ufv/DGoI5zobl01IJXNvDAV8W/HBylvntKMh+AmxfCusnhHLZJR+1UNVKMy
GTh0qSWvVGXin+JbrQ/KweWyLS33ou8F3YZn25pTH98qE+y1LwLqYRRqxsu8UCZzLvh1cnhAfBx+
j4vz0YNfjKlZXsPsru/VpYySTB+/ZTZACGyU1GAGUaXQkxPUOLItBX2g+cDgXgPzC5tX25FBf7ng
6//+0QKQ0N9ZX7AugcwBMQtoLCAXHpaT+NBj5/qklgQZa2mkagXzTVJlwyC398LXhL8vGvuuCkP/
zBVny8ZGZS5smYcpajMx3fQr7B+EDfgwxF9/RInJIo1/EDiN5sD6Frzr5ltpWvp3y7AmpNQuu5Bn
q1QGufykZItqP91ZxSSysOX4f7gsDpJGNmj5S0gKfXOTdiGPCP6etPUbHqcbynAoUjnmZCNGM0tI
xGBLh0Hc8rtqsE5HpjMj4Pfw68YTRqAo06ce53QZBSo8xRsgbMFMTnMF14YdP53pfL+iwCac5ZyL
PPTQ4nOcLCTS6/07ZFBKvs6Amgi51Z2thyiyXEJ72QoDT5/6B152XMsnHrvi3ett5daxS1BLy+0T
yMyQnfB2d4uGkPox2h+oDanew9iIUDyF/tNrPW/ZS0hTJEOOcKD6y/QBB5YBZTmWF6eQfOigirQz
H5lnI0prwHc0NWBF49kvR4ZUDCv8/nDUXSOapJXvA1RjhIqCIRu56nFZRE9hDQwRnHFe48fNtZ31
QTrNoK8s0IMLSVL3jtGXevUnxpbfJOqJdzO2vWDenXR+/hNF1psgLNUCdofqAhJQLZpHLkHbTElh
zxNpch9fAbEjo6LYHwoTyBNORS9FNfZHKwbWNd3N6BdHaJlllN3gRfxjU5FIjy+QVl99xe0iucAI
GM4LT2qOCMfMAXFuGuzysrHsoUIQUhV4nTs8umXL0Pq6vBnm4PEf+GHwHg4ZiMHl691y4c6ARbrw
/cB5e7gzsusRx5tv/If/NY96RSp2uF1M6V7TAwLh/I8WJlj0tqPnBDvM5kqSGHGRXImZfbQ0b+wA
PPss2R18Xk8hEJnhKNy5mDsSObzDN2TpMgbjpa6kio0V+TvhL0I+4B90uiMiJVdKDRYN29TOFSXA
ddY8kjj2uo8cM9peKd+mcFT6VDzqaMhZVx5hwgiWLiTcdGXNfR4BNgQNND2VB9VoHzHql4523Gvx
lIYuMuFTbyL/bph2Z7vL4IVERDapwXK2XuWLfbKZ0mmI/VYs7HPXh2giHPhvLfzCBLTCgLYUjs94
HgXy9kCUg/HGE2Rx4XysXPNwiNeR1gep2+INGOWYi9OafbfRz/5l1ZcIUULYrLOVStQiNDWeKQPi
ds1cVyrqvNpNi01Ko3V+y+PwIoylwwedcQML5DigdxCMtJ2KjbfORy0yDk5j4SzDSVTfbMyyyerL
w2NB8c99q2O/SoPDs3okRId5W2JI8S/k5u9gGGiYAeP7zhssf2GMbRoZEGhnitRVye52owV/4IUn
8LuDlIyjztXpRqEZ51Ta5rSKxjc/EamBlpxNPIA0NebERKXCvJrSZxz6VPhcMLcbRTQMlT4MGMpw
5z7s3MSC32PaYt8/suoGfW5YV/QnG4Pdwhkj8bZ+iy3/u7MEfGUwvyNdkIbEJmCNkehf9fduhKfn
sf019cPE45dJGScJIiUQ6a3ZNE8yB6hTjVFlTmVt7ccFMSkqRsv2UBkm+h0bSo56321BZ9e0cDYc
ZU+Ojvcnr21DxQ13vV7neZFfaaCFuHsI4ysYXpwRv4FLEJI7xQnC+0iDUAScNcNXbtTGPqqs6MDH
5Zr8d3/4zHCqcEcdbVoDjqtJnUPdiC4AOM4/u86PGQ/ikgw3XN2aqor20U9BT5UlCI31ZofLqGgY
n3h87jggskb0cHTjnCc7aLUEk5EXV5MZMZ2Nax0Iw9FbJ75+Suca9E6Age+NS0NFfOVOpl5pNRYp
9O3kDh3KvgcrZ9GvYIT+7I2uCV4qEb84o5rUCNXfJauZ22xB513gTiQhU4Obkhe7qk2mMgrPmasO
MZ86Vi5uXEnr/dquhu10Wc4yskzSLoyGwRysuiMpMSW7AQkgqs+DA+ddgZXhx4fYmuoAr9eEBmT0
n1wsVWkw4FOauW3xY8Has/8j3/WXfNdGpqgf3Yo+b5Tz17gz5oy8jrkE941yYhsmbNcRJWJcqKCF
xr3d2/nqIv7Ud81Cv9vOC5I4SwOsTKrw97ZR+Rgpc0kHmdHz4A41HtfAuMQMvhHCQSsSX05GXYhr
nlSF1g75wYgke788fBnpg5OJIBxrdcL4CFrCn6GgBpBh0JIqbAYPYJuUo56fgDiMcYH0huGH3BKI
aS/RWfEap4/tXyHj4yIzJDSv+UPHl987e5IKqA4lD2M5S4FziJE/8pG5v/o5csMre7gAhsPFhVq5
eE8ZS4OtusS5YSVdz/GFA+foioKd5vzKljXYrmiGmTrZbFcfrcs7E6gxkhLFSZ7LnE3/7Y2Tw1HK
+ghRitPAV5PxHSpiYHtUGLzhy4h24v+aN5Lwnc1Nh/bfW74VCvBcjPb1i+o9K+0IPcEqObEqombH
SSl2J2WQnhVKmMGXEM6wj/CDyf/Fy0GTkJCLyKUMSOlNXLZS1FrBD2frb0dxVZEdYcshfpUkCRiv
FI3g3euFOiNF3Tgj0OQi/GaZFQpSobQWRWPhwFARG50hkaqcuExYyHicPC4qPpT5a+yqeVTXTZuM
bjFEfBnal8yiajHG0mP9JrVuO56Wt9rq0FL0x5VdEbPMbVjhPE00j7llNrBPhJ/W41QfZeR/LZ1D
dWRoA+PnkdzB1Wcippfo5ABcvduaJuMcaqBuHYtHUj45PmLIM/nW5XE0joOVx+t0kamPgLNBf7Bi
LGE1XzixuhIP+GbBiM3WfIZsHsPq5dNXaEnNlpGa0cm1+JvtgVmHwOvGPbONrzf2mcxoGZhXPpmT
xUf1ZFa/KFdqDo+pNNUwOXb/mTkIGqTXi3GDDtp71cwUpZ6YaM91Xb963hY1/KXj5fCne1ybHVpF
33+8HpyniGn1f9lP9m/7sClIidy1k0o7MXz3N5OErNIJVbBjJxzL9inV/JSnERQmlQ8w5cLVdFdc
CsrfuudCBslSaiYrN0j80v053Dm0E0f42CN+X3+/AQ3n6lep2sJEJUsrpax+T3aQEkja4wZwv4fA
Nl93iCGZKT3tztublj0HimvDibo7TR+t6jaRbHwIDhSxzzpsZWu1wO2/QsG9GShxEqL2Kinzer75
8Pc6JttqwNkWIN3iHXJ+jPqYW5YxMXfZwF945a4Y6Lkjtz9V409W/49fu2dwEiCET5nQgi7YeDwX
VqnsxYJB9ZWhQksrv+SfHVDob5frhL8s+gjpsU+Molff5nam1lQLXRhNg38G3QzH4H7h4ZbFhnOc
Bx5W+CI/90E6/SAi98py9UneULmXyEMfOuJmlzS08IapZ5O7b/3FiwMkvgfkeLLipBNLTFbwU4+P
yIJosYsLKAuuUBb4DDv5GBQ6wB/0pzgLleVHPxIG7TYWJcidPGIj/uQ9bqF+bVOhMdyCi668L/Yn
B8gD+ufdA6jFQvN4P6yQizcKpjQkWt+uYO/GCVwJ97KfBPb+KGRcEd3tlota7u88UCnkCIu4+F9f
FoK+PppUBwnJI50WbPYdqwu+K/5UaYjfgsMtbUwRU8aAYqn4zF4okgXIGovm1c5gYe5bq82WUwcv
JyWRFPo4EzuVywo1exyWHsCcZAsuaLbWU/of3PkTvnP80sNWsUKkBFUTIR7kMgW7VPLr+OGXDk9M
016Bypxq/pHeU+bsx8VOLWqYC5KayXa0ap4y9wxeVuOCSAh8OYp8Sa+JY+qCKQkoBTz/Pqoyk7Bf
ar811B3Zzm0VjNj1cQ320JpGlnqmxgCv2KVSaumI9DoIuo+89E6OWsUdsA74Je4dF0DcDbqf78xw
61C088wFrc/XeCJfXlBdiLDG/oEqyE2lhYhAiQuiPctJmOEsC8wWZUZZlr1v/Lk1XEbQ6fNuqdYf
9FGzywQnfdlf9C/XXpyotHsky+zVpDSny95mwOCJ+v1ETsiUb2V2JeucBzuMlI7tSixq2af5A3Gi
16baiiuAGs2RNrMh7UTPcSAN97q9u92jizANxgpR+HYtsQaCnkxy85fARymBPFyYPpxbKF27uS20
Eetpz909BEc3cbLW2rN3iWa5f6+zYGL27o4UWyOmh24SaTz9Qi5+4XX+lU89d3jqYG+MY5I7mab5
xHlrkafsN++tJHqBtULIUeNGWgKAsl0Q65217X/FpiF7qhRX+TEuqdvlewOzfVL0rsnJaln9D26G
EJWuVE0rdtjXNWcO3XKAMHVqE1Uyw9Cf5cK9J3cQO1os/Z53kHn1g1YCHi1TNo5FUyxInKN0MN7y
nlH0E1/vtNgRhO7yBjKepKrjNN1dklpnSwtVlSUngDYoXRMpwIjBcBoW7Fo1VaNEGF4jfK9C8Vhm
fErcFbIWYDiNjWa//SSA7TR0GY3OyFMDmth3+t9O49Nd7n6B0+G4YrM+Hyix8pMQqO6rI4sXszQ3
3N47rSs60aQncvrEaa2tzfZGwoBaxlhx/8NrzVkk6Hjbg9E8LRJVvnVBhQfylS0dFj+p/3UfHx1q
56O0dWpJAH1LICIkJK7eJ2zuBbXyA3roSXKcoPn4Jsf1Hj69zNtYQLzK2eBUlrpmaqBu6eUf3Iqv
AoMpr0VoUwua33xyzITayQiwa4wUu4BfO3mk6/duEfdLESpZbwVzcKAWcxMtDjrlhYRXvnZRHkk/
PU3nlSmZ5PHOJ1G5Kaeh23LlJwxBosA1vzzxioA3iaRrHTG55err4Q5nv4XEzteefksWXfUjw9wv
hOJB+dO/NZx8VlK+kArmAEkl+GrWECf9AhLkRgRgb7URupGIfzJidV1DEQ0m2zNvLPguBmbfCPIj
Lbkcd1R5Z9R+6ekvkg+SuPUjtqBgEWCwhnoTiMede1y4NkGg4sAe2sIoC/MO64+gVp34BAcoBSh3
/iF7DIPja5I6QM6z0JdAPEDcaTHUMCU87cnaQShpGngFgI4MqLX92qEtSkGUQPuc/iXN6QIoZtU9
uCGiYiU3rDMOAVqamljwGnyYLrWhYiwYOYzQ+mV2dGudECdlPOqBy25lUm/EsoIl2LM/6GKzRHve
jv+vLbG2TfivaJgcNu2Sb+IHDIYwv6nPzpwq1O6s26vMrbjKtYkfZXo5l52dvyubPiHU4SQuXQir
QNGWisX7nvWuBtF9YUdbCRIFWnLxSCMR9tBRN/3m8aXFGzcObrSTopNJ1kgzzjs/noYkALKDwpmQ
2T9m9UbzuQzKvdjbGLxpV8/6QJMeKlugS5NnqW7whjhohxn2nb6EcOPW2DA2qTahf8ozwXsnA60c
7WfXsG59tTf6GPNwLau5Wel4MjvqrGxw1IwDKctgKYSs21r8nmw+inzw9KQduKFYcMmyDyD2VBWM
yhMHQ8n4xrA3uU6eFsRayEilzRps3R9zTzSG6r6XTRW3ngoyGHMZ6DARdO8fR7YyT6OIZD5/hox5
VCY6M4hNsPKKA2u8rx1RXkbFE77mJDz4enRQXTSBYVjvq6+TzBykrDeyPHWaUkcLNq77PwzlL0aD
BJApjboAkMkv16rc+X/ouOHoOKyxiFs8QuYP+yWhGZ/YevzPstvkRKhg3bRZOKGdoUbyvQ2mQ1AI
tmmMxM0Jabe7mk1YQ7kSWmNDlqcK5f9xOMR3vPEnRS5yPSqab87N5VaGm3UJQ1PcdoYH0Y5NkIgT
KaBJ08Q06jg4XS/orl2hdaFoIWUTxijye0YR8YGfiEQdCv5sZL90NzHj0jpZ2FWXER6gxV1DCbrb
TlvKAsg8xvbe3hjzVa0ToQUmo7dPnNYPWvaynhUD+pq6MUgUzImpMW00M3351OrrG1M+9BaMmXEl
1mULk1LIkicZd6vrXhYgzuTaDsu9dhlTvHsJrGII25rRQXxyNxDUJ+SMpybmz8KP/u8SUyEXU5ZS
AT1/Gd/Gp1xBxcWEJvBn3R3O3Cd+XBldSyoWEuYw7tU3wN9cF5Whexa8OZr1ktaVXdzpjV2rfBvy
usH8nlrQr9zKWs0BntFKc11qkFz3cOg3DW25W/STeHK1e/VV5GFif/Iz23/95VyhZnUDTE1r9i6l
oIA634pM8ZPhbAazOBEW0M/AEn2YsJNIKpe1QydMgRh8VER7GgmmpzGfhiWYBaAUAufMg/NWO26l
OyBgge48tqS4DPWm1mbtazBKwSVabsfAhTCCXwCRUG1vECqO2Np1cu/gubJmcD8blWHHdKY/axtt
bI2MuyqbDUC7blPxVQYl6pCKeQfF7wa6Dvs+13uulU1n1H0twjgLZyW74VIJPP3B4EgzsPtDKyc7
gFSvnlntbPreEQcM8j5j45YRedeZnDYoIMgMGFL6qQSCFvhRLz/Jze2KvwY6DDgYKVSxyaNSQ8p6
t0H7uIUM3sFDBGtki8XPdIKIKJ+n7OtOaRFEQ3IYGcUVCcb/qPf1PN4rWMeuZ8qWHF4nHGX5zVS3
0ehHKPDVZUCZKwNAiF+D+J0lNMsEm3QF7twT34tBLoJY90op90O9RNH7hIdpzbymK5cUwbVCu2WQ
MvmK/ePUS0BW4OS8l4G2usaiqevCUIvMsVC626zvODiYBLDqzzybOq5tXSPOrIpHfKcf2A5Wv+y+
rkoTUeRv0bv+TiyViPbgq4AmJONnDqJl6IcY8IzJWdIQz9N/+FFfnqhfzfj6Es8JGfMlJzZskpEm
sr5wF1yiM+kBrHDYTRb6Nt0oc8YvRZnl2mDZ/2MHCfIOxRGTcT62xiSSDW2JRLiTglLjRS49H7Ty
CZHvIKj1feCYXi2yPT4DOGYUfuIObzEnhORKwCGzZkE+egxawJLVW2Tqe2dbTc3Lyv+J6PF/4sJo
t63TL/88fcgI7mjJ0nxqQD0kWjWvubgBk3qNpWtYNYpykbz5gWGWgGKL4B8UzX6y4G1Pnt7kgBL5
rJpar8himjOJDtDYnj8szobBmRlgM46V5puSBY6wL0fH0fpJrLUx/JsQz1DdPA4gJYCBw6dMToTB
Ejh0UBekXGqiQ6qku3QT0zoJWHy8v6JCT24Z4xmqT3m9SqRTX+3nJMlQr8FNzzaCwqMNzgVa13YG
IKMV0z9Q285uBDJSSVdonBdMqROP9G3vyBxbmYsUbunTs/XCL4m7ci3xJW1vDiZOv/PW4zhlus3x
1hurrHgmiQ7wQo57rPpxQFVWl6q1AsvOT+qwYYVeD2GOiL+K+W2pHZMMZeo19vENH6uNhA48cp8O
eBCEKG2o9cka3hISbIALuUOfIzRWdp2Fn2ttxCjXb+D+ykZcN+qfhgKO7F8E4c2NpIxLSoHF2DVE
h5RoKBn8RRxz55YzQUwU+n6ueY60rFbWMjdJzjQEQneZ+/9QFpVE9jZw0YtO1cmhCB3zGj5Eloi2
O2Pf3fVJy+xn/UvAhGMNL46ELTDajdqVOdEaGR75UcDEoUnwIGVlfAhgehc8+anMAUYyfKZ2vly5
A4TygFJ6PZr2YK63+uv1UYn1mS4XsH4Sn0pPljcmIhN6qmHmE4KL+nhb79mTI7e00dRpW+CZ9GK+
E6UXrrcajWae8yRPs0KepJC0dDWK6rS9j/bnjX9iYVSaSyf//LEfKhDwlLJdORMotN60lS7z7WgF
7TclTsl2WTUsAUOlsD1BkH2/IG4cN+wlaia0epn6qKlybEHvBcztBswfsEorgt6EL+yOpJwOS+6E
Y5/+MA184479xtA2e/jFIKrbAde9TTZkCP2MAM89Jaf2PcpOfqiPgIEU0pbxAEnSVYCfFNrqt0Ya
1RjqQSTzlMQr7w+IcE4GpITUvIRDF/Khb1IoE2kHfYyLKzIO/wZn9iwdPKHsWsSAU9cH3HB4i5YU
rWigQHD1Jnd3YEQyHbNmXVNW7SDoeBvMZlGwd4pDFUa8OMEaiVzb9YswkqrSf0OyVn5PQOLoFyK1
EOB4o+H4a3ipNT8AT4cf6AyHSjc75+GPgWjBP3bFQzkIHAv3M7o+bTQRTJadtLD2swnznuQe1ZZW
1pec3o8vFPv4209V9RcvNS99Q1Th/jZaOBi/LJnxv0sE6mORgAR/+ZS5CcY6XkDBm1wGZvdmuz5H
Jx69BKdAenSA7OnAB413h78XqZalgeunGow3F17K9IYJc05EQa1dmejyGIsX4v7qNvbU7+iBB+se
leVf2kkNx88lJgQ2MjJCCgU+KK2jxA383SqMhGzdY8Mc/aQPxeeZCsLwzRiZ7rQukHj1ZhXyOzPS
jrcITWqOWOWF7OyJ1G0AU8/Qhd5bGc9UNjrPYIecnaRdXkNZuXKfSoiKvg36ozxAg1ypQpJzD4Et
I+/lN09nziet2wGzhYNDbHYrVayLzl7Mg5lL/HHkREcKQ+gsaPTS+C3hOhPnI8FKT74LRZQdC6KV
jW5pOKxuKdd9aXPTJ6bgAtamCROr9DWhmpVkcdiJTf9x5Fi7Eo1xfxqpEdgT0qRsRfEGgPhGwrqh
74XOckggRp4fBs24nrTwYDWICzo732Cpj3LVDfZXQhcTXPlaZ3UykfOsKQdnoQlkigv/sUUiN93m
hjAMWc8JXKy4kVnpSzs4Nzo2S2ea63/lufqKdUgZm0Ne2xUptbzu4iwXFg/prKrs4KJDgDEa7Olu
H2l1P/wW8fNtaU3YHE3qv5cDewG3/j2dFdSZI1r3D4lpvoD8+9pNj5KhwhrJCz/8qztyVhca3wZP
zWk1bwRmDkHns3V8JjtQjvQvdqRp0oihl6VpBZ5nBfPzvh3ebgRwFZxpj8a3PgMjKYfc3C462M4Y
OmoY3bFeDK6rNZLjnN7fAiTMn8oErQyHIgO/2uJbWS9n/oGuLkv+MhB+Bo743noJXR3SvSuhq8E8
UUurrRVWGfffF9QxwrlaZ0SzlI4772mHzRePyjnTQlZgoYVzysAx+oRDqct4DhxcrXNaHjjAT0BR
56okLmx0Y6F7KfBAEsXCE6uNZ4ubAUvHbZdsIZqp4+/aqfxsN0M15vPEyGc2j9+KOo1n5veosYiR
DmvdDkIrmKW3gFpuR3pYWJfFd2GIybf8IFn+9OH96Nl9gkiLqHQxylC3rpAaSrwy/yK0G9bV7DG5
SEO071BuEtvbW6giecY6/TZR0wdGabjR8QBZyc1lG24APsq0Z4qzT27IrAjzNGUa20j5VI4+/EEU
3xMl2g3SONiqcjHPxjmcA+OFD4tzF++Zs9VhJQgRBUk7bnRTkWxTsKxkbEQ72A9hx0J1WNa5JvdY
FMqpooaSOwq2+B4nLe/PsRLmW2Yf1TDXFKmapjxejTMyr5WubjgyHw4PVd1Zg6wAllR9MCvTDqeD
dnHrDrFgR6T9qq3aV7ceKJtbdj4fpcf1S9nUipCwI7xiCimXNIlQWLI6ntbdnoqukrH+s+uyPg1o
KsdXrdt091LzDcNbyTqN1a0D8jii85ROa9pf+3gwxGb9jxdSoKy9eu7v98Xga3h8bIUT2ad2zJOC
xOV9JhuHtft/F1vZ9wpuSlZbsqqBrVxpMN8Lw8OG8TgcGtazHCZRpP6A5NTrm+xHBe7seS209VtZ
q48GyXD5Yqpfqz+mug+9Rdvml3JhBOwAXQ2GWtJ/PYsCIiURWRgL4HuQMk/jLXnNdfGWXcGlKfQX
DzSAQwb7Ed1kn4+3IFgbChPKJxs5afA2ihRiV7P+lWaTz0uokZFgunM5cNDzDX71vZaJywTE1skr
ZGugHIm3TkPBxv5vU4fs+uUxRfbi4DH/JWCQ9QP/MRW9fQsp/9OParFnt6C15dWOXwJlprDUqm+P
BlMGsvXDmZHfh0U81x98IfxjWaIdn3H+M32LhyqPDdzb4+VNXJMGQQp6kjVpqQxQazhLX2j3yZ1p
VNVXQDtwaVw/4V5nB4f5xnpDBCkxVPfPn5ZDvccvRIPY1JPrsSxyme7Alig15cKGNainIqH+wdlG
Nqw17hhGWSTX23ZKmEK59Xvc3/L8dOM6eOxuSqUdwmKDeShIPqJO9blxr+7zEavURk17Htu+CDKW
MwlGsXZLh9NBRDGeYK7r3zU4AHPoBy8wmqpOeitpdHrkfEBSLFz6W3mKQgGLAxuyUhM8fzQm8fjF
tXUPdrEKoUeMEpUyNQQDOx89I0VqDLU9pSRqoHYc0WPPBTTqTtWx5GjBF9Xx1iiC38xrIfrg3hWx
e9O5SN+oeJ0Ookg8GvfSdw6Dksee59vqslS4ZmJiJxuWvxaTwpLBoUY+lU0dTlazqYJZ2PMCwtPg
ca2vDteQEn7Ael0Yi78igcKPGsbZ4uutnTBUl+EuoKWAmzFP4eQb3iZhCNTWDdmj4BbcPBFTRGt+
3VDNE83Ms7CkGIZSnKQNLiZw9uTRpYd8STE9G6kFfJFoZzxbBLKMCZ4kNQidN8epGd9W8q3APVBB
QWlrJ4w4KRM5h0Y5ywHoE/HhQHTBzs0Edad+zuyVUWizthi6ejpck07/TgS/+qf8zHJbR3InDjjt
7mbQLLNay2S1Ptyy6rYgegE8oDgmWrmv2R7153o9HUwCiSwme8KFdubs5877KYS5ZrpOGau/FcOZ
bKiSQLkzmQHP14TFTKZyFJTGaMtrkJrb1QTV2LGGcajfs+8SU1vDvjdZXiefoZ27za3R3yaZnrqn
Rd2v6p2rS18K9KWEEQ+JyGTzdUgQC5R6xxy78duJ4SIf0AmtSPWXbEDgoj5Q85l7NO8vgGdvbT8c
b51CO9CUT6s5iAPONTa9mnUslIqxecT73KLEf+Iyhoe15utjZ3GWKvlJYtBH4DIIyniw5KaSx16f
BHiAa45ZAB5SiE5vWqoDxczf497hZ+EK8hBw1epYq7y5oaf0YSRSxQHuR9r+2S0P/qYUAB5FoS2W
6N+Vyl8cH9u9R8ZFVWGVC4bskMoL0AZQffuVf/tgVHTaJzRQYJTgvpXeWHU/5fQhhyWeu9dOR9Hn
CLMIlGDNJ1dTei2kSue9eKz0r3naevyMeC+7fbMfRsth8fl/Z/tUGmMCUbxuDVfYxO9tynEJYmX7
k/pGGhHtUUq/zG83IAYhcIqx9PWX1kFYHLomFOqRcRazh9ce6BzHHEBcWF+fYq53oLpHojCbSTgA
5V67pxAno7xKi2ow8JHmCE51L5HUHZhz6/dUoDuaOdGDXtmpzBwHwcv767VdPghhiYzwYTygcKQm
tJezDoi9fdsK4bL+XaGuWUYxw+R5UzElfePgEiKru3VTfyiGHMdfAGcY4bUqkhtynjSBIrE+Io0C
g1a/dLYJBv8C5BOcFdxmhlOgS0iHUeWFBy0l0WA7cZdxHfB82mw+1v67dzZjwJTZ3XlAXiY8CqZf
BedmLlj2VSgU1XHbt65hgJcNerhk+PVT7DXHQVDLVs8Z2jbjJVQvoFAP9wNKUQBlXjLvf58xlnt/
PSMiWue4QDlfA8wyLJgwOE/hD2usCbsH+BKKq+Cw5trA7Zr5ToJLxnN/Sd112hVgL+Xy1Y3tvGlw
0UvtawquKF9SkyN7DsGLN2/FmzIZ/8zzNMWWbwWKGU8hm1CLg4fk3P88dv3x1lK6LsxYojRmHshM
EV9XcJEDMzYFVRG4Dlt+U+JG2IJYU4U6RpmBnq9CBN8g41FdMXZfLWRk6dexqIbLzDp67O/5fJAt
fWkOnpFADhoHj4NpOZKMFSYirDUslICNcIe4g+1Zesfv+2a7JQecrx841JtoTJDzqz6RYk1WBIYu
t7ICgQKLQ2iloQfuyDetttQUI//QKCAVyGFygrSLU2KmZER3PZ2Qn0mVgrAuL6YOS647O8vwgpFO
JlkNmSvAs6jEa/DZ41QUTVcNIUYLOy73dJx0+Xkws0l6PVueF7S8TOQBAU2HuGP1Tjsc4rGk+Wok
KFsrj1AzPM7BY4C8MQTZizZXZZDbGNHA9EioIk/80t+pnaFz4H/YqAk5ifYyZh+HyLV7jhK88vse
vNIEY6+RuEFaJgSj5/yYYQPBg3AA0gYz7A0lw6HZ2fOZArSunvTDtNVj5i9OAIIlHpyr9+2OzZKK
7+c988n9NRJaeRkE1hgsV0YBEHNMNZa1T5KF9AVYXRf1I07tlE+HEqdGiaUcVSEjF9JG/PeVH2VI
UvfXavjYnfef/LFnqeXrb8Gs7Q7OlcHhpM+HZYE3O6QchQuBM7Xq1VHKuzXtnO3mT4oJ8vxR1QxO
raqWiJ23kngbRIz6szNAIFJ06AeUvIuK1e3ZME0OGbMJBUN1/Fyp+ta/v5fH+hcBVGce8TdfPREy
r9pM8FXaRROhb7fxbgmJbL4/U5hBe8m3QP+6a7ooOuiv25dvH0sRxVam5hHMDFCf47LAbRpymgis
tcXQCkUcjRqgm0kyoPd1g7TAfoch9LJdObAjn6bXw7w/0hSEuRyUIzPDZIugvNjc8AnuPm4snUDw
10GYoTjoD+rWWu1uGk9u4aDq3wZnZEa92AilRPmmDC8vIQQsdPeEFNlZoROowWSlC1HetQH/BQSz
1410viP6hggXN4G+e55Ou/GDv6xakKB9BJq8Ry4ssfDE22B3wWFtH95ikQ4VdUlxZsbvgzx0VsS5
M0xTsfkL0VVL1pAqJQA3bltGYjiBbiKvg/edpGVxX/2+ldgojuh+SxpS5KQVTH8Ov+5SLOKCMYxr
rHJMDhv92PLtmoDUJaP2IO9hgx+zPn//M1l1yRFAeXCZF9BwGMij8eIaUXOEer0cqBEe0r57X+nn
OK6VMbJFe0sYOGmrv7aKwMLWKd9bZ9NStyQHpOm+eMvdwK8q6qH2yTZKmI7qoLrKTFjB8NICNoKN
U7cUbP9DHtw12/xKtFr3+3ApiMFg/zCVhbfIt6PNIPokmVpTjL/bOOOfY4BRTE+uPOJxgns+gNet
dZlDe0z7x5vM/GG2yiyDWrWzyRsZ87wb5nNRt7v1l90KmT7gxLHRIP+G1bDiMKGw/cLKIGbXeLwa
7nZB6C3IxeWh5OU7F1mdoNvhZA0KPQY+mWRX+N9ErU3VjE279lqhfVr1xFY6QTshqO/f4y9VcAN/
Ml2ezcAhOfa+VyvoZxM059wk5I2brdHsoiLd4DDqGKpGTmjatXhvWLNHObbXnVgNlfCjd9Q8hWGe
/M0peOY9apW8va9yr7VeuP7Uan1Id56qlpqhdFu5uNozvocT8Mpq62ZCAC59jV6YvL6l/x2FEcL/
7oDxqD3WlR7pKuFyJ1c0yapF03NOQ3lNGmHjzmkgqRgryySP+GxbBFFmD1VTfFOw2ewAGKsPmBf4
mVF7sFWKKv6sBV8odxb631fjNBSihtcKv7yGt6VjQZUjhJKJPbfEFpb4GcruJJ+VgaYn4H8H8ynp
2pv5pNbf4fkneB1NmDNEgYjj2W3UAojzT1umSLmttDqD6teWof7hD/OLyS+FHHMrPGRNW/oBHJ3O
RZZcYlBoI0M+IizGzxcK+FlMBamfXF7dFeFLJagDOaafCZPTrzd2n6bKMshaqOeJMZoUsFGb3iN4
Ob+V5GyIACWGo+xtD/ml0vJzlb1dXpawfXxn/LbyMqFOw9M/YDVHci7eTUzuzJIw72CImMaXQKaY
6HJOsyIfNn1YSui5YA6OYIX41+NhG5Nw+Q20bdw/3GysnH9iuSZbulBrun9lEhkTfypbZMhuI50h
lhzZEubeH5+tRWaE1eLFle+9Eovs6P+qD5HZ0I+qVx9proaKRglSlLETYXtObCypnWpjJIrBJFwR
J0pTuOAZXrtQxyPNx+6wfn5XCaC32Qw+9aXmvqNesu5HE/N/YgtqYYwkemntzgJ+d2klChrVMf4J
ZGBhZAgv25RLFP/kZmG0ClpPQW/lGGtZWiK68VU1fpWfJfQ8M1WDcCE7p32BF/BamOXUZU4veumy
53nCCiFdBvv9tPWMMn1ib1S2FdYvZzGxjlV3hM6QksB6VKIK0z30ZvcQrr/NPMbjj7Na82S5Mgk+
lhqDt/VmGVgqXVhb/Fyn+JXPGvPMaApwDfGjzzcbmdIxQCBvttkZUpf7XINXAh0EwkV7PQ5DM1GM
Wdd1X2e6AroXTyqpt4RnlxVMBADBreFghR/4OX+/Pc44UmR/YpPmMhmHOq4SfIQchR3jvl7PGps4
m3WlfBeXBWm7olmX/F7c/US7/YdRbagfGvKGgOjV37cFI04wqeuWU2yint3xJ2qOcUUbfQwIorKy
ofi0mDsflJy3nsIUAuyygmFAQqvxUE5EbwGjN/8Z3e4Io+plsp7xBV1NEnFvenyTeUQr+/Knfr62
TeMbXn6y+O63ArU2QVtL4IRZhp9USfhyR408uCStFQgsAoeNFFGr544GXNlGAjrrrDSPa2PR4I43
jfCir56QUMMGEyBZLdmVptfyCDJ6bsRraOWvGLpYb520PaY9Dx8rr1t2g7bRu9VWvMiN4EXIon40
hklo4fDpahqlCdg7zMk+dleCiO7MqbPOJgEfDJe+08r/7F54dLI7KLGxLWQ5hdA2lszudUVnEFY5
vqbs5Eptl0yOY02cDr0JjwJqvB5QuHHWTiOeMpWcq6UuvrAMdsnRIVpjtugDekc/AbE+ozxjebBT
JYv8YRldaiISGVtUqOnOsu9ANqCqyTc4hQ/sEO4MtxACaDNamJfxm7dj1m3Nynfwh7JtFp39Q4mg
wS/xw79AuuCxJGQb8PKH0IUiKLp5vHCIl0g6TP7GhJsNUlMAp8Z3spWG+IkLB4RoEjMDX1GcwWJa
6ODkrLKQRBEx3TUTOrYX1IDRfEI7prWYVK9zgYQ03Gaxw2dOpqkvajqXKMtLMUqRdBD1jU3zTF81
a1kL1KDcTITYavZon5wloAYuMXVc0Sa3iA23wtJEQOwKw1uO1koVRNHQT+qyDmwbwTEcYWPpeoqy
2zM/lzDbuGpuHfhZU0xBSWjoDRWDijJcv2o/MlwTHLaCWEVr7VMafIDFlhQCZ5SElSNzThEWYcv2
G4/a0gZjZI/dQed6wZY1qwfXIkDX/aHTOlfIO4I0SQx2RryrTcZFuC5/7R5ecBxTNYOqAri6J+4h
XHy1wkQKsBMmdgWsI2MkeBZNu/fgPti8V0CTVBgqgGbDG6ZTJ16XD9ZsyOPY7/QW3QeKrhVXu8m5
x7MDYHm/5KZqgdPd8GWchsa78kADo3S2s5/tiPlsONMbx8f7938JdVl39Tm7IW7luCwW9Z7KEari
JfhuR8zMJlBvRVF7DmThOC9sq664iJU/OZlR1LZtFJDWs59prCLu/88B04nCclaAOxv6xTXLJDiS
2U7/ODOzA2og4dE+ECH0GG5w6EHOCOqmDJeXH/FCVlofb6FdMksMlXdI2NR5kjt+an3hetARHqlB
JmYAiU17FKw98xXs/0nedRdhkWti2yzEhKlWDeDCl1bAuieQIL5XNOhmJJWfNaWmgzdSwuIbQQLe
no8RE+WBfCdQ5SAYHTmUaR/G7S3WHZ0ukSEd64RinQI+thljngb17A75dhWqrmk8AIsZ25NZX2DQ
RF3dzs0t/Q25zzAqs3gLTFrlwc4if5UPCGuoA/tRLG62pGesN3Vw0lmFABz1RwEIZs35rljCAEbF
ZaWdilZL4y5n8tdP49bzVQy81dWMsZRWP2a+Jq6Tt3tWydC/jvdSFVYRUtEP+/Z/kHzJDPW4BpE5
g9lp+0y7HdKrvAx4re2xSh8cPY7VOwKLOY0//9JAzVSkzQ/hSFOEWzHLREy6c3oaG8HGaleJwTQu
aCpnDM25UrSl0pdlTQZG7sPinl4e7ZzWq+w5wwrwvrMweuAZhJ4Lq1DEjJ9nXlV+sElw52qQadML
1zQZbYiQxMx9nzKsTLhgoibUrmh1cUE3lTRIuxDBg+btsWo+TVyy6CyVxRxWlUmVLXmWeIPgtvvl
7DVvsggP8i3qgIAHVbE58UKgGjoYx4igGTuzTlYSa6HfTfLmBlIco6zJ+SJT5+mCU0a8SDzxgc05
sJd56PxKe0CFuP9PU7zeLfr5NMJhdPoLZvSloXOtG57GzWgtnrxn378sciJTmNocIhfFY5NIjzmM
4JTEILKBESlFONmjUlTX4fuOPQnaq0+9e+JMkE3h8ZPEgkz9WRgiQNUGttAw2UKYq9rrDzQHY8EV
stEoCuNGZs3LJh9yR4Z6ub+eGY3qzDosxR5zvmYng7WpV31SHQ8RfT/JuC+RGn2CcdGCvZTeG6JC
0kxc5IUMcKMX+2hdj+pMtNtXU0Mbzi+3TpKWvGM4xPvZx3gGvmkAmzicFsNwxboh9EDfZjzye3UL
QVv/PyUKMxcM2kRliw/8wqcYrCMht4v9hacMoOwgjbJ5GenzeEME3DOgK4spma8Q/n0IYfBoVB0q
ZR+Kg4GPejukpuHKJ/WmAxmchc56rhCFJ5z4N47tJdDQteVvEP8TU6sWorFbyMwIkH6KQcsHtwKV
EtgPZgw/THQfOhs/IXK37e7JJxlfKFVPFme6BytZ68XVoVNrys9YFJWeaqIKGikd8qg+WcyLo40i
DLqF2nxo+STkgU3fu5IUNBkcJrW1+l0n3w79eyR0Cwqg4zORQ/6rShXLmxRrXbHP0uTCn8n8gdJv
NyduSLzTzQGouWuCfDkjKToRJZMJlmnxk4mIDith4+YVp2E0Z5p0/CA9r6I+1oOUOF+ilVyqfo3T
uOffiHLoTsI9makSmQo8JQc94nOZ+R1RISR/XRHbj9eNH9vsBaOa4JywBOuVdAnTNMUsjWWLqCed
nJXKs+ayZAjvmgfRPant9rB0hWQvUNWxLLdbpjdCrfj0IvA55S0WKnqamNK8aFvyvJGw5MMS3C5D
Ycbc/jKXW/YHGMXdY6ytHzA3KiSon9VyiNH7MVEo3IBFWEYXfK3BsBIgqr7J76WwUnJl3VaYLUdJ
CSU+/Ux1AKgL5qrOdaJ7WmCqvCVGd5ZZ6g4fHXuQ8ik5CnK78QS5NVfUEI0v+EAEzXS2P4eCJ8Ud
kay/UYNGYn16+9rzYPOHs0Ki74B7OGVOhVhLNlv7cNKfN2okqwYHbkjpox7Rsy6Gkjg1xQFIZQ8I
x6Q0184JJpdhOG7YtFoiO/dx940Wmef1iYYH9I2+50geyH3pxzSw8nKKLEHsk0OgCBMrT4Si1Jc+
69J9chmm8S4bCdbkurTmwvkHgsOQI9IkkLpU4fjvQ7DhWjSpYePcNmjPgfgyCoz1Mzpi10kEdQtQ
ZJlT0gUKt48fX40qgmOGWz5DsNdT5eAfZUYXmoCAhu6lkwkdupuw/RmfiiBll8Lka93M/jrDWHQr
fIsRipuqk800OAdQacaTdBVuV8oaEgpirOGaSL7IyrhauvwXHupny0XZWxMHjndhkdH5ABBLYMfi
FxUvdXLz97Bg2XrG/JTtI1kgVi+aAgHsoLnDMF9IENhy5bVq1SCH0Jp6/hewjbYgQbgiRxrtyIvg
dcDFZ+W3BSbLmc9MuanT36prOIz4EQImt5+EtDGYwA240w+/mFr/IirQPYTx6YRCLJrgAFvlaa6p
8jWk2Wnjnui0XKt9noWLGh/bxqSHb0WOkFoOcHlTrvH79AuRM5/CbTr+2eSF6tqMplZ+Fngjfgzu
6fdwh90wqee5MjGUYZsCiUrmyu8MZ0jtd/ml9NudlMMb97qaYn3vB7M4pg22xY8QOm9Cod0/RyxU
fDNE9FL2MsyovsvbRN8WrJmA5hmQ7q/EqlqNuDpSQmfziaR55qtsefClB1vt/+Mxcw4IAS6MAIJP
lQlQHzwvGIsOnVB45YWxQUlhnvRxZqn4xHlcaOPPghl7wNvVqGNX7Rx3NlTB25WfPTV+ZMUwVEEe
Ps6R/EXqjBKk6JS2BgNQOFY72WI7a+8Lteq7oiISa0Ko+ZdEToJc3dOjdT7xbeQj4pXUpXMIMbqo
tdZk7tUMkwgvVw4acKD/CdMB/8g8sT0N1KBQn6TcwO7fNHJr5lQqZiLH1OHZtjqNcK5Xb6pm2dXa
Kg/P19dkaO+4kCM4+pXiTxMTSPlT3MDJc4qwcTkYAEiTUBF4drgTkvjKnb0MYz7GH9rc7JaFBUSO
eay+1/vi5UAfhegYo9IVeZ6PmTwsLjnCkBt2FqwB1CI0Wm2ktAMehccVEX3blntnsmTCccW8vUaU
VRbuG3EtQI6cRiOpbdW/F0lOu/MZQf5apfdqD9sZDV2Wcpx1n6Yy6OxJ1+i/pxIRByicER8Jyzhd
SND5+C43o1swpHurNvRn4OzzZpIhuuV33nNSzGpEtIXlBlPIWh3wzgfb+aUjcZ/CM0p6Yk5mXUmB
KAN0lwC6MUx+J9hzY3pQdPeJD6D7O2W8YTMueLMN3EpyKBOXnV5Wh67U3ZUucy9T3iHtX4Dyhh/y
QsGN0SkeSZZA61wUJs3IrR9MawFF/7ZhRdoGGxOq52fjTI6eJSHnyVDLuC+LPM9o6evd1EbcizWF
R+5f9zv+aPnCOArSxVFpfjXL1VFcrz5vkTYhe+mQOKg/wlHJMzOULgoRaTBY9G7qbHFNNqLO+YIs
j1Z5MtZHV/33WgDtgZblvLGN7OzqWNqpbU/YJOZ14jNZWp/NwfbSIcW6PA/jwOVD7i3R/hdRD93e
tmV4psaHUHe9eZ7KykE1nOLhJ+cNNtvD9f4cuboyWfetC1ZndHcpU128RJYgnaG4XO/0OGbjdrcr
BWLwiVEzGccoZCCAyDwzAKWvkr4uMC939lhD6CFCvBQIkj2h2e2vegYwSgfEQaqJcDHQfzbSsBtZ
xUreVGoLrZWKNuCynq99IhDABiaJL8lWeL/BT3x08ah5Tmx0FyuafbpzPFzqrah5Xcfk6vGSLjwu
szpDTK/34Pwi72ILAtxo4616QUDOkEbJg9mXSrbWhNZ0PdSdJB0INLl0G0VTdYnVCxQpS3D9jUUH
Emp6c5gB5Sy9a+M8B5qYgNq25o46bBpQq4P0RsDwYSZ0FwtbiXWxf+Xv3Jsil/Cp6e0C9GXoRzrp
Z2hOfperv+2Uez/YD4swWkftCAVoVD7SMF3TGgIJBYMC7//Yv4d2YfCunZTAXA8bvIOo6bQkV101
ErL8S9ISY9y8bMdqgrDwyx20EShK01Gctn2SRV/rxhei5SV9bv0eYjepxkSkGGrHBPzHjYaiiDU7
4tmGUFS1oXDAIv0qmiGL8QHSVnF02umaVeV77gwoc7/W5rff7n5Z80hUXnrXM7FelAcd5DiVLmN7
bdJzzT1mz30xYul7zGls1wkVzYMNGSX+GeaRL+ueT2l5lmCFQZ/rWX2XuVAbncV+thEYkiUWB84v
zbFQ7hKb2vEZGzU0l0im8WUnydyZPuVCCGACjpcsIBfF5wYXLdWaZmEhKH6onqgPFpp92x20H1qc
BTn1/Itg+/tKxRGylFTTgeFbQflUuaf70fbPeZFDO1AOYcUCIvntjFun94E+y0i+XALhHONY1GRr
S1nKvspH8hXD+sWvCfdJCsgV+fi4nHT4oTSwJpDkDivFrbG65ZrAIZpZEpswgklj++kVsUbnlrWL
v5n3eUmZ7FOe7aKr2B6LXiVkWVnMamJjl33iLNgx4wvTLgEHGP3cCr0OXCq7rBVLr/AVP1+3URDK
LO97D18C6dldVIIHzVlpyZd/S5UEa2pDs1rtz2nUYN83agK55zvFYG2GO3gDLhzpbeVKeFA8noIr
INUIT7YNpy7wdT0Tgo200mFN1vHn8fxr51fBCqa/yy4a1mUjbBaR8nExZYisD36yY6/KphzyDtY4
gaaeBhsLzYxl+SUYLzjWjiBR2iO31GC6ndClT3SLN/gTeMtCUSNKn1AxE8XS6+A8OmtUR8yvjxwu
7lFOvl9RxW11EbaNEPsva5jw6OwkZLmftS9UFracwUv7Z5D18JwcjWn6XGbTTVCaIaN+3Oj1tNRY
aObk2iYMmp8/AkQ/mQPqQHFILnyHxDS5TPCPP1G1J3d4V4n46ccqrQuzoVyuu35wm4og4XBkDxVH
zxpbbWiALAPtq9UAnqQ2CjpGn6U8caizFdI6YqxW2uSxUohBhmRYqHUdmBQPPRSuSLZpikgCW9/A
4QuBDR48Lbst6/xt4E1wYIg8sADzBHr3RqD+GS6/njYmrVwNfHXIolLSpQN9tiH+R+ycq3llNnSC
MNc9frKR0jSfhxQeQ7ipWgv4miFgj7OeaXBaUyb1r0oXTmDBx34vbVKo0arB92ZYFYQMhoW4CXsg
bX2sbUasLCTmCzIQlxD0Ky3jh1olRJ02QiQXONISa4BsRRhWsmxjwSTtlICnKNlHjxbvAvH0xu88
O9Ll8Lqdtg4oIUzLfh2AnQHr4OMtXtctz5XRIwTyXqI7m3UWnaqrVqsB/r5mk3wtdManjY+1Fvo/
Hi9oyV++hGv7oBKRGXNISC+pYD43jN78Vf7SNt/V+NeLT3ZiBI6Q7GTzmC0EpaYOAk6/awMMurbD
BvESRHWlDVgmZMhXVoW+EvyL2CwyxCLzDXCkXGU64f32I4Af3+8kPIUuyUtzlP7i2bHROPErmwIT
x//bbKLIjKQTgCnUJtIIgpWiDlh34p88WclVPCpD/KlHgfw/eN7We3RAsVnWiZKjrEmxqn1NojcD
13pW11C3Sjme9Yw79gXPjj8H0JBjG9uo1RI6LdIeGRgguz39apy3wyX0yNSXxTNonHe6FtAzI3r1
L2AATW7TqIwhx65Ym01FhHzkw9DFyf7efxSd8box0GKGLRVSKw/MeybdXsmZf7Dm3hAAqVVUfnG6
/q0sCJwxh8cu1Vw3vaAuQjAji7LmsHC+1nuiMDsZlHuMPhAHTwIKUBBX1icPXJwtu7X8+HFhTKHO
BgodxwvBLPUvjocMxQx4SkMjvPokZkbcogSKKGtKjfPrKTZoTXW6NLEqgfSwDPpIbZPHM5O/+YFz
kUJEpJggAVzgUmbGvtvRZrqI6xz1QH+k7IetbecM194QwgkXji4ZOkFCEwTvW8xwE8gSvzH2CNjn
tVdOHi3zZSACjr4NOfsoJoKymypWG16qayEW4fAtS9X5mVajKgD1yGVpmYFiO/vnk5xC+++gFKxg
5mpVzcEyB/5UkS1faYg4g12btG/glWairh7hhX5go8IwEAyglNq9Ln3tnUk3q4Mex5DBoJ2Ha/Pu
VlHqrLKkhstTsrZjtQzOHBMDFb1+vdxHagMjgojGZWlGNOyCPL3J8uCvlPGY39klqSWWmFgiQU0B
3ZbMMVcvhSiT+ceq2rrxKuyUTxtDBPSrpBJaCubRxJrvX5nbVJwxAsOnAAJ8mx8svLKz4DsJo1VH
icDQ+vUFes2/MQNx/7WBSFC2tUmYEZ5EZ4c/L4QklgwZo+LD6lVlaf8zbPNfCm8gj1qwHr3GFVGv
RRSclI0JCfjN9P2oqlKgQYhygCycCzxBrMQy/5fS89e/bJbtQFb/J3VRreFXvUrWZJirx5EKXppj
180EFBxQ4K1IOTBqQHl4ms5VF+LGZ9h0TrDhAv4SEn45bIDAA83OxH9Fi93Vfn7MzXsa2let3A6Y
1bl0GxX6tmPtymKf23UHX+pYqHXaRgorcnzLHPWZyB1JAGh/IptfTqImk5A+EsFkg+DJFgs5cK0R
vgr2OKhYBuC0H/he/UT2hLcclYglYA1SwTG5kOkbZKCfxLCV4OL74sbrj1FLjm/Uq3eNDtgxXU9E
aPL3Bp9hRueWNp97bHaX1rHM9Ev3lQBHmteZEGrdNlrJr+mBvPmxshT+sRRZSdZZvnqHHPcT3ZjI
k7DJRVFzShSC9hwPAnc4pdaeiTv6FtXlqb54USBoNeys4/qztEdqoxwEaik6QFDzrUqTjxGcNOPw
FfJPGJiZAnKP1uIn1nKHnaoqTO8goJDRemfMpWTUjsoAiloJxvTNugFeXZGFCGBzxePAJ7aCBDlN
2OC+9MzhwZd4HZ5FRAMfhQbdtyaL7G6S8696GLAdNYjTp9Zut5M74J/cuNarCvkvEl3Q/RMP1D8q
N0nmAIJLJVZSPDqsGD8pQbDPa1EzsM7oaJnPkkZcsae75VLRhXoEq/BxE6Eb0hWW8ot0opKsPi2j
q7QzC+McwdRIhxRt5AHiFHNuOzyMn46sopCo00oksa3fhcQJpbsKID52glBRwS7XeZW8ErkGvOWd
U8yiZwmHpiSh+qucRukQKQ/W3eRY4byOFqS2WImShGItDsZI+kxUEjLb9pT+8NqRlmezo2I2oR4r
zOzlMFAtG5n2dbE5aSixc6efjHewEF0FUoNM1qzazFTNGyGEwf2rwj/UlUqnR6SSRTORUgapW6BS
8Lkz7ZvGrKO3yQFmYwTWbWIAOK/YTsq/jUEqgOeyw4OR2hdxeTW1JF8Mw44nwbygxE/1A20Lz966
RxhxZjCSQjlViSDdL4N3bI+yOdBNtysjFfkUBNVcX0DcAAIPah48Agn9UOSSIm3BKO6/Bd065Mqx
ZWr1tkxwvVQcwJOw1aRHu4c7GkQ2FBo3yhNktSnR+g1RrmXVwdBwBB3dBMZVqcJqQRIw/IaQ4uE+
lrvCFVJlrlZbtJqfeQBpSg+Bo3jkE6kCEcahj4e9Jia3Hzv0R2YWnOiu8up1BTwFC0GdFLYW633r
E9shHloi1WUlrSWrYNCgaZq/A1hhI6uWl5c+1C95j+L2Tkk/17yeBD7Z+BVrFbrrS7u53N/s5bbp
lwraSzRcon5t+rmamfs+TSHJa8pOm/ydqDmXAJqjah2oLl9+L2uus2WR4b2jWVX4/qm/mtXTZC6Q
rC1a5JmBF/DtbBJXZMYiGIEC3hjodRb2wCCowGaK+EpRIxUb06TVlvAqO77Eqfg83qGw9sohMBjY
6LfW5nrgSPxvT3TBTPF6OKZLRmvFz84fnbZ979gpPTm6VmzlOjgblEjlQ7ziBSvcL9+cicKTfYkJ
H16BmVlPYPdVFwA3RSIQttVglbaXtNpFYcAM+Ia/jUS9SgpjuIYYn7RCDeuK7pwX2qxWB2kIY+iY
Aksce2qu4JRSxFLEE+iS5oD/Pno/3njeoPzZMcWk2OmhKeb3lGGz8psFwPDR/FEO3UwhpYE0j7ep
TmpAr8nf/en9SK7QLOUuuFm/B977DrGv7louAsEyO8U96uL7idSvlSIDXl/2//6YbwkajQxnjhTW
BDVTxPB9qf1oDqbH1dpr/M8AS3TEdOKGO19rCcUS1LhfILuGxWW9I/Sy3Fd7Pdw48zHuugPaCiPi
inQ/58WLGcd7HRTp42DspjIN829xFQxHPPtRAs2+gRNT3EHAhaefBfpdkgiSUmM9g05ChXWlXJQB
whsUyKe+bkfMViBd1LEbNOFuzoz89ZWPCNajhjpO+Z7BNvsgTlHotwvduq8XV4fXbx8hgW5Ifeai
0zdzBnfPyKsS7Ebu/U6cOFw7L5oLOPOZcVGcJgUTzsviowgaFRJR8jJss6SJy6iU9dRoNuPliA4a
rVrSL0edCCdgfUW/5gPl13SY8vmvn82JHBt2Pw3veeRmfMaX8pN3Ze+qIhChjLN9aG1PHFt1ZzGC
+NcBDYdGg70gZnW1UQ/Kyr2FLXbpGC/h9/r8uvwVQ/x4EWun6GxgRLdu4F+gOn3tr+Mf7QlyQNw5
12S+PioveOYXMZP0Oj6A84sJjS9KUdiir60wVsKEx3dx/D/I62Nli8NDv4dfr4R5tYju2ZTsDqZC
aL/NvvzsZOwlPT12oC4lU44QXFRDUQNXLF3DvPN6//qaBjGfBFkb7L3oRz/9JdiEKS8PesQ8OJyh
yHQxJfuiV1f36VfiQes4bnaS6uNeyFPE4C+vZWrLNQA+0m5lK8nDnyAoFzC6KBfFN6yvJIIQT2MC
C+IPtu5RFHKb/O3ONpqAiWPDh77Pv0s+QQcKDxClgVqMZf+EyXkVuMvLfT/G255+FKKZ99XeOHJJ
erUkzE8eYS28yvqGYnjv0kPGlwPXyAAprtcXO9CNv3UHJCvLechMVjIby2OnDW9Z4or/PIu5wSsJ
31aQKkX6iZXCqtonlriwJbDWH3CzxFSgy/yeT15c6w9auWstK1kguDvMqq+fbvfSMieotulhBpt4
7KS7U5k8C/jC54FsOHLLTUB4xHEaxdWeqCRN6A57K/eSpKXR2WF5WM9AAKtfQwqzyNpjdEOvnrY9
ty74Vm8t3ah3RIC39vruD/EOvNUuCqdnRcUV5Vy5x4R2F5fu9/Sxd5nY9eSW2w+bP2m1xyBo6aXs
66Fc3qjECHxN8qEIZDzaMlJYcDUNH4QAbVhXzNWCs+S7Aip4XxZDHsB19pOKGmJMykyUWZgHfKta
LLXSY/IIrHyf7Rf5ilVT7oDwWldIdD0s1LKL/a26FRXPal0ipptoqNvgPNQbxQWEEHyaA+rzwpVW
oKsKiZrhUqZF6L+2uoV3/lacDnrTTbETkUDbjRbkm0jH/kNZ3ZxqT2Nu8gItIyjJW4rGtlanBJNV
9wWt1iCwdwlFBcKgFFi6ENVVsd1shqhxL6esGvDgId95bO0s8tbel1EaM9ECZQ6I9Q1HzyWl4cAa
XvzsVatB12JjlXaf7+RAFZSIiaHCoqGGZYXGxmg6ySz3CPUmsn/qPAHHFgzDG3jZNAaqghInDpJs
WGw5vZe3VSEx1364RHoe2R6NMJ1NwpZPa8ZNUQuJYvC+QtmF7ZKI1osM3oJct8gKnAJM71coL/us
E0nIsx8dqGfyFZxSQQ8n5z8uauj1CY4gnim91/5KUGmeHMNf/SZ1tSWIQIfulaHJVYI2cNVDdi4q
DL2FOyafAjkUo5dZ+JZKYHxvxLB1sar4sNaKeuLyL80oWpWNVSJ/PfAi9f6ZIOS6Fm6eClOApbKY
S9P5DWXgCVCn3oea0fst1kPeRq/Vsjxg20GP/ukM3Yi9pYgdScKIw5fCNuIROBwzBtr/pWDIj1/f
X7D70d7K7ILkaQ5Vy44GD2lEFxCI580emy8nYmobhVTtMe7jKarMH5BxLpQ1RwwAcP6IgbvVyk9b
TRqQf9aLkqGMCfVP0bkTumMdLpDHO5OvEEHjOyNZ6Qzi0wo2j6j1drb6nGXZU/BjoE5AjVFKT6lR
PrYT6HXO+YSXL3iAU7UMT3rGEzP7YCbw2/f4E9aXW95X9yndzFAQBJPMwFv7WdGziwIDislT3Rpl
7GpP8kvzhHHH+pjlbUuphrQYyazkBD13/A8MKK9uOyQjKuj+TG98p32BBOp3A5j9f/iBML9fIWI6
7OGBjzSSi6fwU+RU/11mOQMw04CFOzzfHeJpvlhy/YZEDF8FZgAS9fv/lmTKNWcy49FVInXpf+eB
mOrA6b6LeBcQ3W7I7KRTKPDoPOyf1Gw+uFEpaGwRR5mwEco41+QVNO8YZPER1Y4RW1vhWHKhvpem
aPHMJsbVkV4O3fhX4xmd17RZ0ax2sYOSrZMhfWN3MyCVOwxN1OsD6l4EWj5fX0ig8bupTM3fWV3H
vm3qgO43tCjB7hkRuiFGBdwn2idJT0qwSAHxRyaoPpWqgZ/TlCbgWJDSUWtYx7GQyF+tU6F6Mc0X
OZkIwIBkWNnjS20/Gnq2Eiueob50/ERpuuRakuHN8zQjPSwQN0oTgTT7ASFqtE0Ni0UIo3o32+Eh
pjzZ/bbC22O3ufQ+IElXXTjbSV9v4nqzO6oW2lhrOJqE6g3AnM7Ub57FtJHECa64URwxm0FwLPVP
kesNaj6tReke+iqQaKFBFdJQxypZTLUQQBh9bmaibc4/y6DGUDjRLz07Q/5xrvobiSn8ND6D2azM
Gs3aWjAj3mZHe50zvYa8hfiTTdd/OsQUzOh2CTi0jBL3xU9faF8zWg1xgzHFPX4mjr4eCgKT8mPS
NwyiQYTITG/UakYd0ZB8BLrIS9610KxgBNeIH+ytLcF9z/uickvMq6ri5vzGWCQhVwcuVtDIWtHH
8q5bxse16mJpOt/E7zHMqk7V8q7qwBXoyJujXkJkR2HEXhX2VEL8SZqYuN6hkdXwUSJMi+gNndJf
0FRx+IeKqMl9muZ7unU9PMqQDilR4lJrhcC2Byl+zZzkJEUvgAw2oWPQ5EBmQZZgA3H/tUA+sMBw
6rHBZQUTKjqXQCknk2QYdnJvLgFuTqjZ6XXqVVmjyz14UOUIKc1huDAFN6ePVJm0IAGO7omA8v7E
YNHbOOOFaeiaZTB95myxk+oPjv5wwoR+/Xf2ionQlPyBDKrrfmKDIYYj3hu3BuaeNcWganYNIlSl
C7opLDFzIycXb3fIC33sq++I+BT+wN9ruyVCnQOj/vms/32+2Uq1E0zAZmWxKa/0FHsYwj1I7abQ
gmSfGu1md9K87MMw4bCzZbVykYgyyRNQULcq1bd7GNTDYP7OX/v43tRqA7jzzx72eSccZbsmGZS3
2ielWtMSUgWaAM9sY8xqSn2qfkrlzkleq3I/plvVJc4hQTSOX8aar9+YvV9C6m1hXeDFSjQZox2S
gM/qWd/6DDxPnYrOoZid0tU0OyivTLmxx9f0pWh2S3xjdjPH2nNj/ekh4FQxBzO9fhuFCgAZmYnv
wjc+ucqcvOyB4eITjlT5/ZMcNXLA21ky9IWO+4AsPwE0bXvsn7FlXyXB64K9hWa2jecLMS49fpxY
InVA6RhxvPKyv4C31UFNRWeqCHTghOOo5xSCx7ygabXFohdPm9DzuKJcbWE8y1+bK24teMg3Jo2q
jHroWWJ1HFr4jPcSY9J0lFAX+SNxWM82jUwX3taM1xaJLjebJQDjerRIxJYRWW4NSoHQbAHqn6Y8
+2BwRAAgK0Ow+3os7CExJQi6cTzsxsr5yXZE1mpilbLz2aAVB6VzeQzT7IPpL6L2/XMdr+phS7qV
6FXGlKdWnlvg7CklqPnIEra5eaQIoDsHigcmx6eSoYKQrOUXdgB79alFR6WLcIAjpaZ9V/oPGIJd
JyvVZSsqUikXVRHG1pQG1kGeyp2uTfBzi+DoRsk11wuzy6gSIdxshNdEfeKWw4t9zyoawQx6lcte
zLd9vAfIRxfDofHu6A7NuIzOEsu2xlX1V8vE+3os955U8Fz+edAoX9vCgkEQsupz/PKszkMiEtkc
96UiP7SVy8ny4JTNCwVCaoppFO+gtiTesRHzIXRVUgxURzNNEbqkHaKiyo1EU5hhRwX58JRl0y3k
czjwMFYDBaxUj0WAgVlcdZT//1k6MlJz2h88VNadNs+R85gjnethhK295Lq2Uy6bT+QI0zxiI5iZ
kFtdzfap5E8iePhWVVHr8qnqq6J6LwQDqs0D7vOAzRj3Yo4d2fx9SKHULjTgI1u968FkHrNWEWng
97se4gj7Q96LgCAVoqUWKCIlFEllGj2du/P8j1qB+dcKEGoW8uvO9Ad2KhO/C3sRgrXAwValDqoS
o+DT69stg+r6pFpkITh2vrN+65wKJTIbaYWslxU7PC5+xGrDBdPTLJkV9L/EmE92if2wmOlmGRjI
8xoEr3AscsM30G7h1S6SeyYca33AgaLghDrrBS+/spmQrwbY/ETmZKT0Yep8ygC+CV/eCP9KXyRH
kW02U+cDiUJ1wmoNnpsezmVrxxnPcepX2tJkqXJQtrlZGgtpEZg1oNuQu2NHo5uRU40nwzIYU8dV
yBDIIPp2y3g7xU5HpbaS/33DRJf9pf55x5LvYVOeneSbl2GM1sUoTqBygEC6I85FlD2aiKZ9ZNXL
D4Tfj8JZfTMUMS2DYKht0BBU38gDyzZMfrrWgyVTCRTqgV+s9ukGv6KOG6WKD6JPyxw/nwDqgbr2
E02wn3U9p71ThrgLWR5eNQiK/E4Z88aWHDp3VoSM0A8x91NCTSF5L97nKo4qgygKk/47IJ0Hi6Tf
iuJCppdCuBcoPZPIOyhbxPrnyq3KLS3OapU2sO3FefsrWe/fAi/DRXTCMSkxblOTYlf7sYIpJ4Dd
AXEF66pHVF1dKd1yesqTUryRvRk74DjAqSYHfafxXm2+y/GqE6TXGxQeDNXH3Y9UL5J9nlF2cns3
JVjTnhHDaYxA0ZZLWEj/XFvir+l3P8xs7eKEAj1Bc2WiJmVgnmSHvFpavAN1g2cd8dB+8XgNKkTU
M5cGJSmuxNC+s7UI8qAUiDtkVY0VNiDQt3FPCpeSG5giZ04TK9XK6f9KrdAERHiWio/7016nSPpC
ydLG47DpHwH3SYVtbsqh2VXZUkby6TDXZfxseciQmu475WS2XKK7MUx1jNEs5KikGRZMd4FFa5Rk
ztFha9umDMcpeuT/ZbcQg9PEvaFKoaIRTb4Bwa63zQT0BP3XPhgQ89WyNx4IeB8xShlZQqUFZ1PQ
kCK+HBRRHZ5WGx7TNrbNdYVOT86Q8O81bgfIha/jFQbXQpH/mYfngpdlgynsUsjdjx8ZUztVaqwt
yeZq0ckcziI474oaFdzJuMj9+S9ge3vajor6eQ4cWPF+qj0wNAO3SOLFXG/sDplR/7cQu0z97vTj
jxdSx9/VBbN/btE+DwWmPKzNvoms0B8dDbdyN5xLy/CToIOPTgiZPGPVzktaXpX/+gRixlvM/234
R7JCSgmo4hL5Lok5m6QadIWJM6zI/d9Sc8F0fyJmze2S4QVDeqJUumawfsXm16A4QKANEpq5f/vD
J//n5gONzMwp/ff0E34RxTiX/ykRRHyCFiKytr5YAZAhwo8tp1uGTO9xSeGsStvwgcvTg15uccjD
Eb2Jp9eY6bV+AbxINkUOfwt2vfNUywSK+r05cdp/P8k8n+JzcXt1Q/0bNYnA6bSzTT4/oK7u2LbV
r4eCQrDKqg04vO8pg7pNBPVfZpgdadcRt4Apoet86iPJOPbEIZPOH/r+SL+RsQfRvILyZMgv4PpG
Cd0cvt5qgQLRgAEbOHzGbqGaQ+PJt3bP2NfAqc13waxY6uvzGBzoAb8vmtJOwDfz/pErY9TuZ1To
EvuDxrskJKOp51tnZrbxCtLb5iAhcFYuThraJCUqeWx3Xs6SaM81u7PF1fr3nFEOj1tCjgBfVEid
gnIe42Ovi88dVZrYC2LehhCBhLe38vgFUDP6/Hz7TIG/1E0j9jZk3AZOaKBrke0/ZLrazhprZsU/
py2lwi0PF+Zbq67pv0+xLRPL2FB0mbX6PrgY6zNZdwzTurL8WPVxwWfN+fwi51HObq3IFR4PRc+9
1QshRm44+xKdoFJ4OuyYfXcZw09iNwouKjL3sQ6cRsHUnj0Jf9/WQ9f8xeAulJXixuHK1Mlel0fA
ER+hLxYOU1e+aZAJCIOfMXPALTgXk7Y0xsfly86ZU01BfxooZZxNEVBUbUjMPyovrwJ1Rtdjn5nH
KSmyV2TQj4kGgoqsV2CKtGVB2F49cUgMHvOYlGZrE3eP1MZ22WDl1Ct+l9KIrmFQE430YsKkyDgo
oL1DXX/StS8bOXulyJch3KbJCoJtzWzG7Yop3bDdhxNnqmlUksBqFioWXdAmEN6A3ituXA+wppYv
ZRsX5/K0URq+sN5lhlvqvW+uUXWPp90zWM2he5SzGohG3QD7WAmYjPHIy1NyufBjh3YaNQyNAlWL
6jdatlT9O0Q415DEiABlXAdE2FvSdlivFqPHhwBejQhgJ+wnNoFs9yC5NsrWvkQnOrUFvg61wbWq
99Z7KT2cfr7Gx3T76cGQujnNVMKTyRcm4mkXX2WgyHvinYF2lve72j3s/YQK79fpeK9Ym0w4wKFe
ChBiDKu74FzMYNFJD1CZXyBQfWB7/HaLYaJ10U5PIdCsUrOQWELA81/ES11GSmq92QqD5OabXemp
4gSpzDK+0QXM28Khq7PRv1iKW9eg19+dZTENydv7kWm5um+mHFZGEtUjO4zQv8oHjT3liu1TU//e
8bsCclndtmz8oS28ClwvqHUqmkm1KzAKVO0QPLWasPyyfo6dPZ3pXrfHlTprktsnmTipyzKsqrZP
lYqa4gG1d93ix9VeSj2QFjlkGM3Um8KMidi1qUQ+rGkVdbmancGJtqVHO4hUyW+yXwiiFB77ZSfV
S0pOnk5LBDSG+VIyHeLn9KITt4Vl1RF/a43KmIDjQ5ilAbQUKUi23DB5q3KehlYF7O0cLAITKole
IfPEceHxPTBYhxYrcwdA/bvYz83GrL3tCHg8QIfe/Nhp0a0M8V7t8yWtacbtpb41P+luTWfm/Jy7
HeiuW5ItXxZTqEO6/TZbnui0ZANz37pgN0j/6NJ92SGa0KlM2uQjcHnWmGI/pNml3mjwGbBCPLHs
aiXiRFsH1FBJo1KCa9pEmNbcKzMf2c0KbyaqKaCCgXnV3UPTQYiXiDv5mpeHOGsjdlAqJxwrnyWD
lpsGBwRj4u38PM2ORiuKvV+3MidTsOabQr5Ft0dhKNUTOZTFcLUem43gWY9+RgdMRhd0na2tT5em
52pFkr3aSUAmeWylR5aO4ORdeoJcv09ZhaaYigmbz8zR0xxAIHd6YrH7nWa5OM6PCvBX9x2qaL33
eq2LbXDSJCCwPYW9oZCFjuiVdYg0E+46A/KpNCNaP8Ab0UEDkCghR+/0W+EkgXR6XWt8pMJzWcfH
3ws01soZa9YRZwgiqDHsMUKpRIxh1eiXOloBe5J2Y70Jg+HFwl6apSA7XKzb2gfV5nBInGqXbQsC
vNK2GQePYQ/Y2FXzquZqBelQRZ+CrcyaA/g8RbVW1CQMDYka7hl2zhpsdCHpPwuoZ8Qw9djwnkq5
bsERmHRydrYNUHkqIzIM6oPxGlWZ+TI+VjxcdMLqqEyWxqB+skPo4oUWkvbEOalnDNt1US9qDOYF
xxAyzFqOHDuF7JC9UgunWQBTK94iT1u6vIr6iXNpU7wK6JzUbwqPXd9ML0/Fr0gJY5VKPj6whKf6
PzESY/J3bPEHlf4z45JvsM5XGoHMECDn59rxwDPn2qJqGf7/rhcSVj7llf6zdkladnOY2wQk1QbH
oQdQYcgsdtln+g9oZreskPpZ98aLyIphGoqZrw66Ebp6VIYnZtI1fV78BclPJ9BIKmGbWPvo2NvK
idtEO4+PZAeAZnc3IfWLGc9gdWy8O9Xcdj+MwR0pAXtA/HaGJKFLOfuN6XlQ/U39ZKSK16a5KlNS
RFY19b/b4FxuYcVnRgwRSr1e2bwR57Ji6ipQtPO3gu0w0GwdiDcneh4aXVkHZWrVNCwhzn20OsJH
D65vTUW3n8Tum0j4ZlN+a2Tu5O7zxA4ySKFXJ4WKhmrWlRPNZVyAJE2opNcFu76u7QpqxzUc3MiC
LLtGnGBa4FYjF2jVqHE/mACgBJWkJH6IZOhhcsZ6HbxXDsTJ+0CqsU4+huZDbq+UVXjtXTiBCkHp
V4QmTip7AjZl3Ar45EHdQMOsgg1pq0WHbRz1nmtEQYO7+gfPOBqGKFt/V0iim4acejwkH6OGtdOB
Sa5Zs2s5mUpQ9UkJ7eCbg9Bel8JG6SNfP+d02V25dGiDjopWMHvXgoWk52chVcMl1mcR9U2ZKwYR
waKCFf5tMei8FpzXBHzlX2ncChdOww95uzEXGffL4h7gTpM8r3RwIEx1ppsYKMMSOjpGe6/k43TZ
eu2Wyec11m5nTAEE0qj9qIh9J4X4y0Vqj6tk9/M91gwFIIpCXgh1h0j8DgQTsXsQDaSP2IEVDvSl
8b6CX9dG0fUIxxHZKQV19vNvT8E61svdnXZLwVE3fVAObeEQyFa54/+jolFYsqi5aIYYi+mmiiv8
0p5qektioG/Rp28OYGHPvKH+x5CjhMantsBCBRjblaYlCzJh5zkW/Q9IlX0S5mcAFSOjpYTOKIEm
O2517GG3qDHcACsvUzp0Hz4VP9pw4+n/UZhHwX2t+V3m+ayTPSmQVqkmLXUOltEW9egT7K6DlWVV
D9KcKcHmKGMs9LvCsqt84vVlkl5Avg6mUgcTmRwhXdzmRehaVCzKooHF9yWQqZ6wle7UllckIKGT
3cKw2exD4WR5CXWgqEUzjmWDWtDbTS0ckyeJO/K9b65WXkaI6gFhkIo90+kOVEXJV0p5AaBCZcV8
0LU+t2TwtASeMWdoCmP7aqxwhri1Ka30SaJ4rsce2bBeucY4pgNqKK+tfhhGHQXtchIUMdGNSF4Z
JYa44zhV1H9NuPI4QcwhrzvZRUYyAKcvSdAAIj2RV1T+dbCT5NbSaHXzeV0vdDuKhaEao/h2x8yJ
EmPXVah18yWD6GfeZn073Gl2vneWkD9D8cJIDcdG72oM3KWZZeSO9s6MLXUep+8VRivbdC26xibs
BJMqqNcLQH5cMFjOSWo1xp5dlmQa7p7GmS6PEJVjl/unXPGBuIcsOdZ6jLRmKKMhZ4im+/MnpnAX
bXG33hKUVgj+MXNBq4oeBWxux4D/UTTsBrwa3UGcQ/+qEYuTbbnOBDHcfnC7bqO5LJ8EiBaYXTyu
xnHPOkgGdoSGsHwx3igaAf78wUx3rtMBy2BV2kk4LqRqeahLsV1OfKUOcwJZdwm2K1xyv5H59WjW
Deckp2J54Z+J9Mnn37qVxJpQX5LpF2phT4xkRAM6WjtPaISUSKGUCUMLUaUagBV2s4ayGlXb3v8z
GkdDEqht/odfw11E5AjBoiaKvinGatxCOVs9oJQOJWFlKOcS+KFQS/Qyjj8Aarx4Rx5VQkOSRzI9
ddpQTfX3e9AKE39OnCyTjVDD8yhriBDTOSj5orCZ9qkJbxHywIGbD5DbiEa9gssv4Xk+zs7+m7Ku
rg0NCcYYRHAvao5L4cBlzfqewI9TXK0XaqchZzIO/dJYhiOSD20o87XQa6aGoFTD+n0L1ebtab7G
HJEGJsh7GHzs9u3YsbZoKII1u5ATBDsXWWQe/NCee1TFZ/fkoIiW0WBxHG8m48e5V/negHMrKsFG
qTa1ZfJhi6vidECdfdFZ7sKAjpSVdq5QIK8MQIlZtjU9gv9hvsBvRPUrgM3H99lSldSpXpLthcRV
mTu0U9YZ5WKE2G0xSHHs/jYEKDykeobrRsBx93Ur0pcuD8Xytffyrx/F5VmQ23GtA3pXwfs8VlLF
lnUmBloMNgXwCD1DT/MNdHBplzPWtE60evB/Ti5xyTnhVPt2ZavLHhQxIYIzmOhBNsLq0eQ+kp20
rH6HvGawRHMxJrNm24+kKRUZC+G2ndkUemvnBj2RLg2+b4YKK19Y/Y7MV4enS96LRoG1EuDhE9wX
fLqNaZ+OUhtTfZPU6oHLmnN0d8FhBDFudlzMgeph6tG6DygUBeEf6kYrEt9OXICt+aMzi7IECYtg
Ik+JHJMlcfEhiZaSH4LVEgo4RxGQVOTpW4mdmwX+8mk9d4ZaOapp8Sfdzqi8MWqtxxmC4fxB4nnB
8KkxG7KLDLbv9/A9sOO7YJOg/ILw+BWfHEvIALL9Bo01DpGYzprM2OLpwKrKthGWKInnqgEO/L82
BC9Z+eAc/PoOlWp105jUw+dQTz/hL0Sbgk65g6oCsFyu90qwSyTAPY8Gt8cBtTzAufbiOMTnQvZY
0Bm7V3Tl5LMC7M+4itOua4au4ZVFqGiWlRP6RnLieIw/OXJFCKzK/M295RKd5lUJij1t4ZmN+54j
H0+pJm+fYkfiDSJleEVfD3YZW7v1dlAF733OcixIQaoPTwbtpkU2piBgJmuj+jNayJh5fCPZLofp
McT6Mon31FYGQ4o9neVGrWXmZziu7EBH6WDHLgjsGBBD5pS/akUEfWh39xF2d1nthpR5IGEHP+eV
q2JZ+3A/cdq8rYG7K+eGalxJUQijpu06mFDN2hOMP1psGRopSrQevUg4D2rlFT/Bq9ZMQi0d72sk
9h3NfC3P88eEiZGxHGsdLGIUlXJ7NLjA9e1SCKgNowZGnBzTgF0Mmn4L+km29NRndMHRbKc1J+Wo
nsNnc8bzv7C0OXroCxK0dkY4xnpXov1Q4hVQA9bFJ1lMxMj7LXi4dmzuahEKlH+72GaWneH1iYMM
/JgRfw26K4miDNq0M2ArCRmGaA25uZVo37YJ5iGMEA1Z26a6Qv2Aisla34dnK0XwM43xw0JdS+Sw
OkV5sQOZQrQLRHQ9GxzWeRGdKfvEmwHqgLsdPuL4WfWj8qdnIM4XvDHg0FbgjCqL7DNi28Dp2a42
Ztt3PxC1k/ThWT/TceUIUg7XaLFMkdfZLTasyi1ES5tFUfTdQaU3fQz8+QrNLeT+53LNNJ8BShcG
GCM7Ectt3EJ6SyXhCXULDG3SiQW5N5odCiFawknATHODNxTuNkuglnELT/V59gqyDCel1+60ENsz
JFJUH9DZlKMzrkDUiO8+fxIP6tmW+4j9tD/H9MjYmKHU6AEBwjSK1Z9nEIFiYaQZ+YIW1gLvw3pF
yMkY20cydIrX8JF6r2zq9ba1JYuZMBbYMex777+xsZ9ZPINHlCQcYs8eFg1aCFEhR5LOFoDoDstK
9MBr5RmygnkSDVo8A1UCwpR/TI11QUMae8gZMXaiPnJ8iJf3RI36DsHyBfBON9HFkXBmFtMS4xbA
JRbCjAB8A0lGpp27TX+N2CVswYWFKfJVItck3MThITbi7qTX1ylnN4RpLidgpnhcgWmcU1TBPJp7
ongSNsCzNkMKpivwjNkD2QCGOoM2uMkQKgL5Yn6QqlTY0ojECmflUJJSmOWQZ2Ddu/8JgUOnxFXF
35Z8CM89GJOHrbYEuvFYxokHsVIaaFC/olfBzXreHtLsQJJF3T9DbryazgIbDw6ib47paQKRwH3j
OcTjUvcuQN/+Dc9BPqpsWZ/Zgt6E0TQHuM2hjyMZel2G3KEEMxoV+FuixOEdUA1rIoJt5lqfwyK0
fP8OesdcpTv8wLnt+hAoj8pcdlKgxdXSLWHulOYWtI7xA72VSVwHFg7aZUoKmzmpVqWEK0zY2+Cx
uwPRifD6SlgKnpyZVGaO7oYH7aQsSwhJMcNdE3tJkm1+yLKAK4y2vMWmd4aKoViGWexaX0epYzrS
xGYeQccYkexk7LajpXizWuwWp8njFIt1j+kl8th2wQIy4GZgYL4m1DwuD1ZXwKwgcbMSTQyCnlAH
TpyeBuDGghtwsJpaMNZw/yzZBkTd8i7Nhfjnxsp9Szp0Lm0ysJvH0MHCS39sk0IYk9xD7O/dEGdx
w2zyuVjqnD/tf1y2l1hKe0wCtYkTb2YXxQbXGyVoyFpyCOI93Y8n2G4f+C2vBVigls5S/BSJGmW2
RCYgopkuzUJVUwZ+m0VMtrWBXlgsjmXUs7yeyUA93UcA70hVX3Hg86sqHkkW+s5ZhSGg8QYAjIYE
VUEqNLy3zl7vzKa1O/85i+LmlCOz6UzMq1Dnv3nsvTEnwpN+lZXs3dnqQWkgO6SwRdET71ymRkgr
FA+MN0mybcPC4e2xRqzAZuV2I3Z2BMlvZYzQf/kuX+xwOgr1akqH0nm6JkrLptSCJTgk+AY7c/KG
cS9N23xKwhk3rJpV8lXaPZJMhCzEvujxEZRxVGR5xdeJxhOs801OKwiFTPb+0H2qd0RnR235pTZ6
qhHVFV6dsk6uabmovCRvRr931jJy9hYzS2e0vEYt9gnhz8UGGgHvftw7hZ6V3SPJz7VQ8LqsWtGA
78HmK8sw4wpXYtaFVZtGLD55EdPaEckv9R6fDLX+cYMTpIvfg2WwhT1DH3mHb9CB9Cf/e2OZI5AO
EZpjNQqcAXYctd3gRgmq0dsj0xIlZEd3z5rRqtCvS89jYOpLFEioLaaqARpLMKdItKoRGlLFJc3x
3CvDO8o4fb4gRDo9JVJwcRvHzm5jDn9W6/z320PowwGPKZ7tJr9tumJ3Eub6189I4Tq36Sploc0c
KaTF+35DsI709YAOwl9okfKpJ2qcl8loUSuvUc/HDmVgMfLQMIoq5oNuKYQeUt4VpzbDY1ztB3J3
Qe7wfUwgzuQqwjQuFljIoGX3XPMrTbYjWHWH80lAvYKzA3kHI3SSCtw3IN2rx4f3na1VK4MfA6Ut
IvxyIun43i5v7FV0stVXFrqEGkB/JNBlxRinBZUwtGloEnxSuY5f88wYyAL1w968kOgzcHuNlSVA
emnOFqd9TFZ/Tl/zHQYx/CcX2TX64OrSj4HA1HRVN6UpmK9O08MAA0C2Ydi3zfNHhziFJiuzfpbW
9iePxROisSRk8+YGkrZpZPtXu+exEf8qXgNxh2botb0kyqoj/WZ1mfQW414s3lVnfqbrdKycQNsZ
OoCV3JtD0dzZ0RgP6xY8RP40LvVwD5sQ4/dYpRrqjFZ5DduxQXynKEjhXhm8wjoYtPI1jOls5DGJ
jgRC6xC85t1jvULV68W0E79DwhXstFv5pl2ndQeDpNRFURRTK5KRzTjbnyECJy1E7MRNRuE8wBKO
uVusiWyEXtrhtGjp5ZG8S8B9n31h6Xz5wQAS42KvJ4uuCzSMx/zm6z/pNH8okjDTODFwz2gkF0dv
6OdEchnUDZaOO0C9W2v7l684jramnnamFI8cQ3g3Ji9nt9BpNmbKn+5b25nHLxWaZFrfBvxVToIT
bsOSXmYdKW+Jlovn9DkCOrb62Dyyo5qv4nv2iXL5lMw3RA4hPYDExQ00lp6t5B0nlZQj1GDqt03D
YIZBivBqQTw3i98uGXGDiKSQLTB3u6UKXJr7XHOdl4soOcjeipBM9kfB4Ff13JoP6mvIaC71uUim
xx61agOdYZnPHg9GZBPvqc9Q9kL38zTVB4dGg+FAjXRwN2ZDyvECX5ez2dueHV+h84SQ58XI5Bia
lUEJD3e2gSHW/PqUfGoIkcC4y7J2a2zVsel02tUyU1hmovbQ0/fE8e0nkowFjIUiibZ62dpOwFYP
awqydRvqNBMaDo5wgeI3Gjr61JDynIxTZvL7KhMmPubE3JdcgbBnO3LqVx3tbc/7uwFS2lif5IHi
7/BwHGSokrcaJjh5Evm/aw9r3B3jBU1pcqfv0u7v5ohCAxJ8jc0TIQhEbsXRVDAsZkeLUw7MLhpU
gNNUk5xLJduTQ9uB+gCWLoj5oePJAQpt6rOmJ8pgXlFSZGkZlu+QNqag1pC4gdjyYHo16RKNILQG
wy9fxAu6ZKm7+d1Jn3y25vjGdpN7vB+00rdY1dfsSw+7SDcdz4Pt4jvfsH0P3H+KUgv6eapXpoNM
M8s/uE9G5jkA7KHpLHyxNS31Bu5/r2aW26qfFQJfTqt1RPqAtA3VFJO8szEA1lo93QcRLrKa8blq
nZScDfywnEvSZ2NSTqZ6mOsOvbETdp3o9yPCFb3VM1RAv6+mXTykTVZg3v+A6RhRfeB2fMJiwzB2
FUxjPxS3xZQEFUFhXV8sqA9+K9t1IFmjqF91QLOT9IkjgoRPoslse9J5sObOJfF7TSKXwpm5uaT+
AJ5IYkA9LIXaFg1w0fHC4aGvP4/4oUCXaZ8zKSg785FnPP54NtrVnTrzjecYn9abAORkM7R7JtLN
kUA/Mces/hneXiimenBwkyryu7egN6zyOJ4qQYAlsdQ8yG9ufJf7jXYTBS2R1iWbF6An2gIdpbxu
jbdit4juHVg+aTYs8Ij9y3EhesQdse1dqqPs3ZwvFJ9VCZQXJS2hxUemfGL2ed5rb4q1p01PqT7f
ICxPXiALwDFG/xWGCbiKQzKquN2mfwqt4OI/53FiPgKcgXE75LXu4LhSxsB8MZXGkf5N8jttJPHl
mTgI+ERqEcKsneauGTN84s66rAmH0TyfcJrXa6SkGKSIRG+2VHthNh8eFBfx/AL3MKd8aAdcnvoU
/ERXgr/AqvfSe7pZjoMaqLmucmD+uX2VM0K1fCuKpsCvVNQA5+vM+LaVLwOUu7x/CrgZgUPNcAhn
JE7ox7VwVAuSNTWA4+dkubwa+l5zCc/xpLPje0YYbUVwrT1p+Q8VZngbFv3s3Vbe6lajJrS+sSxD
qse2TwxKJBnZIj3EIRHK/+kcjvlo3mIxLQ8A1keUCGHNIzrIbPHctSn4KTGs5urRAQr69m8bES6l
2UJOE16RYM+hAfOOGDVBLJn78fdNnVHdDQAgjo/I2qzKGvIBVhvQiLqquVfG8IuClLgDhI4twZLH
TUf5rBhLFLrSG1AwhbeuWo41od8YGJaq/JhnGAIKgdDHpig5QyMvir3BiGXfVJ6RqcH8DaVCgor+
QuerITvBA62DhCj2qZwJ9AJfjgaVW3YGV0SofdQ2n2sxvYlwlETJ0uHvNX8tg62Q0+pcU7MD0gpu
AiUS5Qsrp22vfvq0WvNj71m/j7MpIzQXYsWqJSIKsKy9SE/1SWjNytS5QzOGbBMl/AvjESw1cnX+
NgqPPpcyKr6UWvCsCTWCoWCIGZ16Np0v+7T/OQTJeTRXfRB4X3X0sW9w/Y+QRVMMpwfU03kKnT40
cu2eyAodOuNNwT5R/xT/v9MxwzplNT3bgqIKqEuRotKLM+GrgbTbHG2BPyPgTouRYw4Hr62g6Ubx
Mhhz+Y1fSGs/DEXzFR1laLhL3NAauumAu703hyjvEEKTWzOO/PT9dJ6IeA/yiATCxTd1uJSDeGf1
AXwVeHOszjPZPe7lI9JOUisqzLYetC4NF/xAGkhwi64u5XGUJN4fyvfDe0womiMD58IwkPfpQcgH
TVBqDFoFUOvy0C93un9UHk/nzDklwHLtcWoSZhKOqZWBvtuWMpA81tbTAV9ZU0ZERMMxDULoTs2S
sHpwZMVc+Ffi4nEX4Nb1SM6fadjQcOkJ+wmjUfwLjf8ntvQbAF5KWMlIsxj4GsK+5Fjd0FMB4EKP
CwwzCEkK1GBZE5JcWbq0NtZHAOKzdldJyrCJTDcXGdL4FjMr2XD4FYNUJWC0/kNoekG7kW8Rl2hV
o9eOdezAqCSavmzs8Y90E+uS/iS+WzQ+2bBjuN8iVvK9HAp8yFNq69wgXZ5AswIE3+Wdu4s6MsoG
fT1rxbuO4X0OTRlfbfVXF8r7HCj+5x9MFg0qWUr3wjE4QKO8SdeVotxUImyx8bcqPQjgb9Sv8WBL
0ToW1ATvcnivUlEkV45vzz062mCQi/SVIn83MBit2Ij8N+FlGugjlDANvzcC3vf5roLUyjGW6cYb
hEasXHWzd4aIIJUoPiG4WPxcjKkJiIgyHvr+Nno4PdEu18Qrm/lzSzLU8ZarU6qtO9mUfJ5rjxCP
ppiPhd31sQfMNGsTHVtyVCRTBt7kqopdj3ICeC+8r/K6xfRRw8nPoWfa2INXjy6DYXUyoApTBce6
dBF8OZo6Ealnok06vT6+S0ejOnkoTDXDD6g+9BJd6TBV+tsi3nwAcTWDo+ABUF0Of1hiT8dA0zDq
BW06mI7AUK3AG/xx4VKxZf83aGbi3QTjczSzayNoFhGI0axXNFczaeEi9G4T6yfqfCkwDKZ4QqXZ
VkmGpoo6lWvHUv/jRQwjgsah7WbEpH3CM0FRMECSdkgKUqBUGFV3TcqVYrF1cHXw3qW87FoAGCza
i4cmKJCJynrlGPnXMCS9c/VhxjdDrLOnm19cUWvR7iSnjyUSoYSjm8kaOGxC9CnWD5W/XgLA7UJQ
+yTsvi+fWvcv4BwAWKyoGwGuqrvgXYoP8cjAFXzA+FUl9bY5SPEk26TD064qPOFur5oA/HDq8Ny3
rYLiere5xJLlbpyK/KMsSQhCK2V4EuPfEKDtpCDLkIb7L+e6AKH7I1llLsPo9Jpfgv7cGUm7gQPt
IaMnpk4hFHttlII056E80QrwRVS9+qcgJIYuFq9xqi5DQm+y+L+wd+gsuTUfjr5DSixxqWItWdDb
a62AmoHR/ETdAQ/tv9tFolBMlV3ecsHpbXVOx8BRHqiWNQGqKoJlRQiYhKasp1VkE7BWyJiXRWi0
/QBiB4QsgfG4t6QrZYR4+q/gGC8DtZ1fXuP93Vc42rplbFEsGlz4LrdWLsATL+btAZ21iLh3+PjE
4iHmuYnqf/nBeKsnqEglvjIVQhszbesMBP9UMyETnHG2IbnMOpT93IADHQgdXOaCoiN/i3LZRVUF
qWtTnoDc9ZIRl1AME1ADGE9rNdZ+hZOi5C8F/5cYC33cJu3r7sSq12wh1DtQrrF3nXN4zCIPV4PQ
PktTKg5ItAG9xs46BuIor0x7ogbGGn8BAeRbGrrVihl1TEpyzGJJ/6ENW3MxS8+G07C0TPEFiO7k
eMCczNLzdu8HITmuK1sDM0dySwfa0m5v3vRJw1IFBjMS6EAgG6h8Mze5UahL7Va0EamQVPzqKDgo
SaW79fwHg2Oy52uUZf5GEAl/xQzxDPQ6g75pYXmlJtzsovpvDlCuDmaze06drELsCBeF+ckSOVWK
NgqkS4nNNNdgGTUtBiOC9fuUIo7GyBm13LoWBcH2wx8Te0NBgu59L9VfKdMhpfNHUXA5KJUWg6nv
a8qeCwQHYvz/KyKXs9AohjYKLbrPDaqaCi1wtmlot0Yk9G/Yn/n1NfY6A7Advj7e0gIdtl7CD53Z
eHhDelqAWA9tMnBG68pWn5GbNiZHJ7feTQ==
`protect end_protected

