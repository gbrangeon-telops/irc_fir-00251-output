

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
PT1CWY3UnkDDUklMeaNBhV6BliNbBJfbhqNG4kOV7Gat9/z6WihgIxC6lRE+3ldfsLvMpYhy8uJ+
25GNPlskPg==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
UvJJPlyuv70VHT4mYaiqDRKTOeGm/bTLqTJOIy8dhI7h8MQzd+YE6IQThFVGwKNg1149OMGabrJO
oYkVzjNGF4B9Aleco2wvOpKfvWGZDwt0GGcY0bPwCYhgwzblbjwmCgPjWkv54osNVTW8DzqpXiHT
yqTtBlllC+UP6StZLKk=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
IvSnqjuvUH0Q1DG87naNrsoN4LstR88Fpjj6aMMwh+f6Fho6xAvTtV8qJudD702FeycqdNzlt1ai
QXhCNPnT2uuSCS75+mdCpNaXrbRjxmX/iWoxCnzawaHjNORHnFYbE5ycb12Je0b7xDgqmfK+x/mm
Rr1i9nWC3k0y2ultNBrqag9B7JWz2UiAxNLz9gIhkdjfo9uuq7n44on8tD92VMcRgnjXzhfwsV/R
WQcm7g2SVj3bLFjNpwKO0qkV9egUmW/eEov7KDZj0D4B6HRqmpo2DevGwrEmNSVhbBsv+hYHPySs
vJezY6TBoybQdPcPOmulaKi4zQJv0qMBHUSRhA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
N4Lf2o4qQIsZJ5JVKzqV74g/C10RJITmHA7UkLNDA0jMmd38lQ4sUVhO++1w0lqqkNK7gbVbdw+5
aHqNf15gjyNPjYW1ZhVXHrYiWWCWKhn1CmdTyUXz9OVBdu2lqmPJnjbOZQNbhaspal62bK34xeW5
H7uey4lH4qjMdyRPWyo=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
WmWXhlbOXU4TrFQt6FbjizC0tiQugH2eLLLRZI3zQRGusS+51Hgzx4mz/p2wkOrjF/inwb9EGctX
9EIb301sFgIc2+iI7RGNXRFy/HDMZa7bViPHFvPX6IIbSblSMhaUsZnDGZ9ShEIypX3t04pywLmp
oC8cxeW8KJ9jku9s++a0XQ670LJrlDd/u67e8zo+xwxrAToVkNJSGwQcgXMc9YDwrXqUemdrJGhD
qf93Ms52+vFz6ikE9Bpwux97WA69cn9Tx5Hhj95T7V3DeqQDYaa0G162sFOeOncPAYjRFsxSNp5b
cwcMCxbjJE/oLyWzhKmrRPek289fPpANZ4f0zQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 45744)
`protect data_block
bIPSa1N35/0+W2AJcOwFo5/+TzlSP6NK4WjvPed2U19A9aScI0mAwK37PUkCKxTUu8FOUYYv4KyZ
dbbIMj6ftN0dX/c4lz3KaTLTHnxtp0z0fXdP7+Sh6FdFnL2pYGdN4P02MTO2qGKh8O6w8BnL7CUN
ymPYzHOX8aE5+j2ecLgBvUdpIIUwbu8Zog5be4uS3dwUc1YpiErXRaYRvDLEiyyql+1MoTwJiW8l
LVbiqN2zIvtX+F1ZtHMgjBkroC0inJjdcK5eEwTeJJnCW7oR+MI8Dp54DU6XVzsPmCOdQwuJU5s4
MHUCm45VDouHk/j9M4o0/C/A2svBSdguk8GiX96nDyPQsSTv8ycFFknG3ihc/8i+DYGIX0eZCWX/
wiVERMzmCMLxBlhmCJAlRFwC64jfNVc4h53/JWCpLFIh+jfxFroXEt6NvkwoFfLddiB52Y9GzFH7
2idNkfjRai9cCbM75hR2/EekrnpsjhbvbBhYw5eI8dUJ1Pb2bSI1PLDfPKOhUucRoj3hJTLvT4og
+TPGqeU0m+Lxs2Gad2Jr6Be8zIXM5Kk2xLhcjBiLVi0WdKMquiSx1LY56f8dFm6nTK8B66ACKhIe
Rfofv6RA+KfWBwpQfr5Yp9lpJ6kSdJNXVzw5rUHILDLqGFhW/GAzXdyIu9CH3+Y7s6XJarV+Cf4K
tX7giKT9MMnt04sMpJfET/B8GM9JeylBu+rF4pxoUxwNkVNYnGwycQdr59vkNcocRU3obfctSkS5
8W8b+SPgVg97rVNus2jHYbmMjybT4wdG0q0S59rORXhwN0ZKucf1lWIaNeKhodwPohjFnnrjpiy1
DIImJ659/8z5w3Yp8uvAC0y8zepLEcG2R3cOmh9Yrh6Qdvv43E9R/RtoSkztm7gRnuL7Ktk8sUZB
9tiJS8bi9dYImvSijdC0S1U8UIOvAlDvOmVTKu5T401K9OYpOE5sH5RJtp2MRy4UVLSnUPf4CnKp
IWGZx6MBNA6zXfd+Z5p3CM7jscSEhzGPUlLfwazNYLpiLtRRNdiQaJwtG81zffm7hvQ68ld9mHsx
WQvvS43KbPR5uVZofBmzxOxeiio9+1ntUsWaVh6I4LsCYQms9BHwu+4+e25MdTR2Kn2yO+rc4k34
/jJrFIJ8XXCc55LbkE+sp4QlLx/U1+n52poJ9CpDxptihxzPhOW+UHmoVN9FdSeqa5HzH2u2NpYh
Wi2O8KumE8ovfhtuClvWqmnk1tEVfcfIMyrTYfw2laA7pUb6BK3ym3oB0Dp6zxjZ4OiQb6m1ssj7
IqQKG9JMjlPaC4N7T2ytSBkcVFOlb/wXgWPxq8xgQj+nunwDY40UHStX7AqZSa172XbjM47yGV2V
kM049Kf1QrY82oN5kMBO7HWrjlsq+ngXUTyqkcCjePhd8yACGsFFSjWd5Wt7NrkbORKx2qbNAdK4
44qqxOqZpijIVgorNClUDRXlyzcHftMn95qykn1te95P/dYwH+NVnadDDDGI3zMEhhxKVmJ1DjTO
QW6bFAWAgyOOzpLYnu8WtfhOH7FabaaCxWNzzF3JTbD/m5BpvBj6118XZPDuKXfjV6DjPjTdQSXb
X9+4P8p6ieiiDNGFgA9E7GNLCRF/kzDPQjKPqJVqEv6+J5hg23NP21MDJz5RXgJZvLglYU3bBsOe
j6QEmHsUFIna849eliTcemOPphuYxvbFuzYVj+w96bc16ajcA0dQ1Xi/ABM7nUXFNSUXYVV8yKwy
fiCv6Dy9+jnZJD5Us35CSHUw7WMk92VSPQOVI0xItrViEpAnUF9McdFq7dV1Yg8V6/vWU7fK2aci
oVsAtoqZBrG+0KcS0InzRuVFl5VQUPBpR2DligdRlfawLQpN4fAgAiljsOqNIDgs4lWznCjOGS3X
wzNmzz6TvasqQ0QEzyjeohf9ODaOdn8tbLgShpJJ8XklhiB+EOSRaY3AmC/p4jdKZq82qnx0J3uM
7QJkR/GAivoQTyINlhMff9V886jbASYgjEAp28TRJudu5EXKIUU3M8KmTEOb/x0xUa2C8ihV/ZbU
0OBlpVRto/l9gtunLfklCHLUjtorOeRE09bu6YM54MBuVlzTX1zpLJ1kI34xWkEVJByebiO5P6cI
FjEdb0aXw1MqA4kWc4pNVtitW7dhcEpeP/GyFSR0mesq1ZO/QKcW8F0PNou7FkGexugb6AXstKlC
4XthVb4HRS98w5R9i1PNOEVlTEmv+q5UVCFsujEgNuj1anE9hKc97wTX5TojC7kC7ibPQ5L/kOhX
+aAB5Rgr5UDFTo8+rER9QVW5W3lyveaj2gJhtReGPzKGIrfr12RX++MX5GWE1LHOOOrQJri9uO0w
shHsYckhgNV3hcjtpBQayXfPuJLa8h3AKgMy89mQsIvAY7Z3ZfN1jmbZ7Gornq5YGLY/wKCTG90Z
IqTCf+HIVUKhIKfUYtCLjIRxaZmKFJllobtXFhK6oZqr74WGkzi931BSNJi5hEMQccCby/ZdMtx1
WYqM06svwsAbZW1M5JBBErFvFjbOlbyE+1PnATzezbUSpDhpmhgjn6nkRYNE80F8soV0kCzXjEbp
cGgnEBh+aVOFwCpI6wvPukMmFOXoIRVc+e3RHaDY5afMctwp/ARuUQtM8xN3fGHWVjdyMrA+jo+9
XTYBL5syAxB215Qs+6wWbf1uwxx0bESc2FpMSR6doPYbyYS2edlaBxRMyHNE5GXvtC2uJlp32vAM
QNvpDvz6tOpK3wLI6bxoEndOXYCx5p0FeM6kEFCKHP9aEtqSzrRb+qhKGLRM28H93NPiLwgewHkR
gp9b+vPqJai29FpCn47TxBwa5YFv9RnSsP3/KrEdqriHwYKKVyp2tFV7FZMRUWcE4yHPa9rtnVvO
Ms0HFpqPvDYZHT1XbY4496DQ4amXl2iJWTn6LXr657Uku/b31nswyeSjz5qLxF1tP8bnt1Pjte60
iy7lDjmZa0tNi5u+mujWUESFdHRrSLZWJQ9sStH2MIzCECDh+yIXZ+sSs4veDA+iFITnMuipUz92
q4sM4i97C1Lxm08PIqAYvBBB+JhBGbZF/WnhQhDe1qehoCoTvYS7ejawLc5jQjlcd1d9jb3EEu3H
WQJdK7I7LgHLEY8ZJxIxgvXehLshQWS/lNdYeJN5sQpx6r7QBmFSjzRxWl7HDHjw+DvYL3dpvxqL
9z3tj/Y/pEXVQoUv9iRRHsRilmHPRwjvktpwEe6MOdPLa+IXiHBaEv/7V/kTMr5hvyTQcQrf4kTG
NpoWpbLlA8FdZ6GYEyjdz1hfxBAnhQZAuVvXHEmrOc2u+KVUoVMAA2T0SKEt1Mk/vw5OUClSPpfU
G/m6HwlkZWbLX0HxcaS2GCHhsOrTV5Z28CUm2fd9UktyjiBMHI7NntJZKipH6ItutIRgHoqrhZi5
FTDpOF4scWOIWDIlTgBF7G5AT34anvlnCLu9t2/Oj+Sjpq0b0At7MwP5yKBliOErMIsUQpcLpwgw
f8ib2Pkr+0jpPip8JST5OVbyuWL3bufOokj0lqY6ULyhVrM0fkmMCuDZiAGKQ73jJq+kb7VPurl/
lmiCNUlICcgOk3ocnMAAZGDp3eZJ/Ce7E1TPwBpXi9vQoUMf+ckbm4REngfeR5SsDPqgyX4lwInQ
BchPnfA0jxZGS8U6ii4HJEakQfip8mPUFpLHNpuIrbGf49k+R1GD6kRUDi3ONpQed7MhkWFkb4YW
tELi3J34cuYq2gbnmlkdeJd4MV1QILTR4wi7j427ulKnFEqMaCK84drnLeOTXySCugzfEinEBCAw
IVLDRorq2f2p+uPKMOh3iUf2geXL3zZttbp1ZV5orlNTGu1u6QLuLKYwVXjbOV0/kzSpFIM6JY8i
+ugfSmA6wfIfNN98tD8zahMPcYKt3Z8c6BvuUR7Iqa0SZ3jKg9wOiUdeJ4TKQ+EK6jYzD17WALOb
Npv9fz08k51HnzZCNWEF8u8VGZr127cz8MLqkvPz707YSqTg85cN6zI5C9kKxb61qgyQehb7Jyn6
UDZ3p6YMJ39TIk/xE3ZKUch7IBw7yI+r8BDIUpGLHwjZy8L3GP+9fi4Vhn7vuFKu7OnsZ1/JryzC
hVQ63a9anraj0ZxI7wEUg4Qx/aUq31HL7YEVzjwdIYqIvEcBylUXQMCX9T0jXqJyuhk11dLVbKzC
U8dFZJ26F/bTrAdM3ze3pAp4vxdLdHKBwNxyR+Ap18crT6XxLff5mZ6qDBdH8ViPDjUS2lWk9b86
FEbdDrM0TrWt+PBOmI192XJRnVdQoGxQAAdDFaZCCK8Z5S+e7HLttRcsio7085z5JvB4ZlynrAmy
mUieh5vMFLYdMie+vs6EzGuvivnSNoPcGcjBm33FUOVB+CX2SHvGOBCeYBD6RaVtQc8dr4wPDFk1
S6t2HBZu8jT1wqLK3hRcOAjWGlsvyusxdFVKL+3/PzVpZPe0VAYAqRrqXlipk/yRx68m/cYbRung
QXatltYiqLhWGXUy4J4PvwL/OOoNSdAF1OedK7j+QBWSse0OFJSsoNQ27UekB5a5nIpV639WB/Tf
U4FEjEoN/g7Yy8lNKCiRE2U90PgTsTxw+AUjvESHl60KimZeGwE9d0yk8wMJ+uMYrMs8uqui+5J+
zowF+e22DL9LIheCsE+sGegil8COAb6MfQILLxmUoLLGcBrxbrudSK5Ct11Vh1pCL4ucmsw8eVJl
yvWVaFvdB7U81LgICpkDI9CKFfUy+v5il93zc6Daw2WxvXd83KTxGiu9D/Hfao6gZji9iYXQI4Mh
xP3PdJYBu2ij93B86YfucBiE43pz47QgPdwGr8yQmlJ3OA35Y54+Z65zUt+sSvqUwGH+9pa7YXj+
J8DBkAcNer2VDqySntd1F65nt3p6zIDNiRdsYrS8Fle2Jf67pSzyA/EMCb2OXSj2IF9gWcf/n9/0
VhytwRcc62T8OM+u2DfO/wL1+FU8c9LDlV3yBEnd3ixdN/+xfyN4pMSPflVzM4qfPGKM2lE+bp6A
coYjouK5z2F/pIxXV52ofbLx9eV8pVg0QW2nNgJehOX+ZOqdLEkdygWJkBb5ozL3UID44EUX493o
sAIc8ZKB7QPSMEIBxaaBgmFJMeg+4gsGNOAmty9+qiR5Fh0VfPZTHdMbCkVtJxQHv5MI6KbwS39s
oOz+Ro2YzgcoUi42Y4t33Xvm9g3j1JWHEgimDQCf5TRcbMGmsdKwDWG84e0fmk/dKnCmLFg4CbdX
xIw0aqCeLsw326FCzqFkLOOhaXXGDGns442pHwRN8crMVSokpi/AsdaoEQbdM/5gjzl0b8sV8CY+
/lYiv4n2LhQCDQqBnC2YtBmHpY1JpOh7huHXBqSAQ94KXkykrMRI3lqYyg4TAT/uHCE7hS4Jv/X6
HBdmngi0ite47Z3iITwopCziyz7QckRECVA3aP4ng2IdTzq6nlLjql7W8M9cDj1aT+hgr+DhFYIk
K9cWjUwmeyCLdreGNOKrFzxbsPGT/mRgyCmOZzWQ4D7k4pxkuvyOUJRzZgpnsM6v5GMQPO9SZ6o6
Uc1gR52WamyD5PAXOIkg9vXEDvU8KKl2m5lJkZwGfeAE/b4OeRmj7eMWmDwpQ0292+vufVx2Mi0W
DoClRJfMQnh77aL+ubbqFhgrnpp6d3y6NCAWv2swgywI/LqG8NzYUCKhvP9o7q60Zp9I0BmiEWoL
9DF2SmR4Kx/iQmcZbPwiruTkNhpWVN1f0AtyX2wHgRJmORkS6e3C9Yio/nPdNlj1/Bp/ofyi6eDO
Brhh0IZ88mMYLYHVCZW7bUmrX3suFTokxeutAOUT+D7yj7/be5GOfDYDL4vGHpssrHh9lnenCvKC
5KScPtOJEg0KD16fiQ9V4krzKjqaVPx3t/VM0m0TdESwcpg+S8h5zasFnJpmjffbB/6hM1ZV6TD4
qYlZnFOkW0mn/MnWEjG4ppuzrqqFHcMdaU0tbwM65zplTW9FfozS6SvEfy7AXV5xng3rqySp39C1
QVX+nw3XAVIMLnQzsBtmkomz2nibrIc0ox4ffmg+X0rhCzcFZw99k2iv4wfC/hF2vNVZuv0LcHf7
x16GROB8SrKD3NmID80jtQ7AKxSG8Z67SMAhCnLWYgHhSiZlL+DWVdRNsu178laCYcWWOdt20ZsJ
VgkkkF6zOA9ItTgB5E4u3egC3RETVyvA1u0KXKYA8mpFxxxUQC3FYyn5AAiIMpTXRvSj5owCKbRr
rJ476X4FOEW3rAMOJe3eJ64zXR8XDm4OGah17VdNHRetenn2weJlSS0O21jk9gO/IQThUQY2oMG3
g/SM8hLGgEhzZnyCSWCjAyK+rz3HImQvOQPSIMDmBkZEJneh+bWauaEttveN2saPNvg0kQSREs9H
3Zy1KmDFHZcye5OVC+nrlbWtk2KjOwtb5+thDAZdEoh1zCdfBYLZgYaRw9pPqLU3LkL8Kemt31V2
0jF3r+UV95IsHHjxjKTA6aoIvyzLefX9LibAlmQPLhs2awAm+Yp/rH39/MC/q+4mVnWRUtVSh3Qe
nA4KNoJA31ZBMt18JgJG2O8ZNUfe+TGWpgINTbCQhknyPPirDYApzQ4P3oM2IWWpm545qCL/qu6S
TNnHZ9oenD8SprJw80zKwjgNPdGe01JKntRD3/40QWN3Hsuej1MnHLgiLWMPZcvXvE9Q0dpq/DCY
Qm5sO0l3wod+p/oQLj4n8AKdlv+Y9MCliQgdnvBq5dzrhMWwChmlYsJnTtJIzO7b9yoLKjikH0DR
ZJWkkRNse1qX0hmxmy0lhg0MyC2USSTz1+U32sEPKm/gWOhEK8/MShmnZPcvx3cDXab9IhZ+ya0o
t/VMJgoPif6dmURhWFczz64zv6lWwox2izFK+R73kaALNxFJA+4p9BkBHI5CgmGhurkBZxA4w6nq
TeoUvTr+01aDl/vXG8s3RUkJWDBzgOY0cdMyMr5cEnVANuRLyq5hipHcziL30Cs2aRGSoNpEnF7+
22UP4iKgdTvz8jsPptH+vr0UZMgAoiITZXI6px7n5d0UeWSDjPAvhxR/Rax0coldsPpG9VP1W0ou
HwxiH0mgJGXXUSRCrdZWK7KCT4WqeBf4ADOghgcGEbDCZvEu9udsafIskuGSnWMERQ0Xm268kUMn
9PES69VdljoHQrP8sDKsQp9CPLP0uwNw4NaOblrjOCOmernFbHgGY4+tutMtKjcut9Zo3GfjTcWb
//WRPmGa5M2xjRVzNXj4os77NX3LWchR7Tm8/38ZUORyCxdi5nUnI5EsF++VJfLC+0Ej/tbfsk35
wC3meaWpE3n8pwEbgV+hsS8h4XYfyB++MB9w0gc6e0TvXFoMdGDFmi5IoN0f+SSKpRL5sMku33zJ
ODCn4//0knDoKWSrBey2E4IBYEuXxUixvxUBR/nY6lEnMFf3ikueTaxtDMZ8Xs6CtdV3Vtg8jtKc
7LLS1oBwyV6D3Jh/19DufuYA+dk6LOPYQMTDwV+MQjqyxAna57Q0yl5oF+IrNEW5FiqcDv0v4tme
89VbYCAGR+z7mcU+kR/1c1J6yyU8HYvYg5d7zRm7EoEtXfchcgDn1+aY6FPsmExPyx6uJQ+dyLRe
3Ofp+htGfeZ1Bzp0cMLDNfVpOfxRaV5qWYf7vBJQFgbqnUU7R697E4AyXoK6fnOrbGIGa3i1bF2R
U265WVTvsvE2/zEnG41C9R2OG7u5rlpH2CsjnlkNlO8yKwRmy1CNbgU+e9RvixzvNJL79OIFUgHl
ZVh5qlFlLTnxevathdLCD/z40dRgPnkIi/Lx90cYjgnqpUEvWkCRefMcy3uzk1sXsy50UjCZ+/Sl
2qAgJAj6d9exqdetsWF3gNbodeLZnhTqK6aGg0RmJ4zr4aquVTK2jXtix19DpAhij5qVIHhCI9F6
QEudqLZZosmGi0WjuSNq01CICREAkJ1wFdHTMAPUkyDkRTx5OmiXiDZPvwWkabSeDCvJ0x4Kdrhd
/66ZoPCKKZ914Bdv/96lntga1tzIdh+G3IISDoLU/kBidHo/Pi1o08vKo3oXhtYhuvUYuoJaTlyE
hA65BAZKGYuwkh5EOgNLQQEbc+nsvgu2bmECUH5EjuGkmYXe5Dlzt972uHuwpiy5UT7SHN9RLDJz
dQJQH9py0ZSZ5cSIKJDZuxr91OPPec++Nw0Y9JHyGQdYaj/GadVPXb/jUlx70UF0iYhg6bAtoxpN
i2M24WpyOvMPBJUi3DMGm8etC1wX0tCo05g+nmiaXeVvZtoBYCLuuXCvGfrgdr9C+KGOmMUhs4Al
jr4QuFZ/tCbUlmxpE9P5tM7+83xKFFj8v+m7/5ev39/8SwJYuqvG+evEmEYs02f2gmAiS7k1db/T
XxtHu+zqgkuJRO1TF3oNswMVyDazj+BUgp3uhNRByhtv6QHrnPYSU/xHj2ET/mY+A48LYR56RaJP
/xk4cGKBf0Rvb36dZYeYxE8ZRU/jB4qBFnQ/theTAWQQGQ2pF4ICvInRHkj4LVUiBO4lHxVz6qHL
OZl/DYwVayqQ1ZZQVZ/xvqfR5oLsLGNC8sf+FM9qCuIu3TQE1p0t5HbofMsI1YpP+7jfWmB7y0j+
q2D8orUEkkUR5VLyouHXYNvB+Ga1GB/LuWmRni9I+GLOtnbA6//j1kyYdy1f0hV7jc+zi0dVZcXo
+EFjj8KdJAPdyrvTEFM4+Frj1/R/Sa1cxESMI/UNm7tY6dczJqeFdGOfZd8m8jtPxCLxnVsrgq2D
QMdfJDhp3OQNb67VANCEub2njDb8cBwIfRmByMqoRw9l2JeMVr/bx4XNCuvmKqJ8H1oEtife+9a7
aNRAwBzsLstLNI03G5t/boEb4Ikz5cifyuNzS+L8ZfJSc0Wiq6rC2ZC3Vx/kV0XWywb7sFjneGN4
zdfRuWYmbJJAgDri1XNsoaCeg3gNIHa79sI+uXlbIjEOiV3U3LNthbiBp0b8J1w/7NwdecSQAYnv
fcCL4o/Pb4yTrsmPqAvN8IeT56AWxmC8qURAIw5K/f+z4Zee0SYTrqhxsh4Xvfb+JeCipn2yvgOH
OB+KX4yyFVa8vHdrrO/HPaXOsod+sdNXnJYfMPPlMOksQ5P8uQfAtgD9AWwyWhnyYEfN4NC8do50
sFi2L5kDzonF01qYcryMvAOO6XHVoyN/sHpkt7iK9vPGVUCYe+MIe0SPUPYZQ/msoNhPwxtgnX/n
NztWNinGZWj/7IMPQsJbAXCPtTMgMHS+fwJfSrYADIJ0ONai2qzY9H5DlyYVFj8F2hsDFT5gDpun
P4eEmVPFtwwy0Tyk69owBvnW68CGzrrYuhw6HomOK01D0yyPoTSvhfaTPzinW8zxnQJl5wC3kMQk
2+G70rqduKYxWa+sjH86pTnNKwWrNiFPmFLURyWjJOR2XTYf5R8W4OdpditmRijjfr8qpy0+EiNH
X2011BSdS0csbXcaPfBow+M7uH9okbqAYOo6nPRjTxWc5aYuoD/0xsBn/8f/Om3Ky3gA6vrR5P01
/0XXIseYgIAV97MtefveiABwjtVR1EnADEHsf/xEP+7Hxud+/bUF86n4p0GUIace/AqCjlwayhFN
Sst1NwQ3u9uea8qNMOaWAq+jQv+I47sOqaBBBr3TPiWysV+SXCTi6HwSzZ5GU8TMoq7gP/IgK35m
FRbW2CqohzIoCEXpmoEh7z4kmWiAkc07oViu7ocYG7LljDBZ4/y/GcHyWAK9N620iamegdsxQIbU
ubrX0BjOa24tvhS7FcapAq0y75vOitM/c6BmNlGsQ+UYcxEnqmOMUzOX4CKj5/3zPANJ7T2FLLz3
bp963bqJVQ0pSfZGAlVi2MKe9VNkF2sGg53rMonalZJVOOWA4fLZxSQE4805s8oNp5K0rqunpQbN
/qowkwhige76C1B5BoRED2iDFB5rO9qOdEbpVjEhRdzsfGlJ5Jx3JKBtauDrsuU1I+kN0ACzGYoO
0cmH0owxuwBzHteCC5ZOf0LXFcgXIb2s4AhSAhe1tNzw8f15M2n2wnCdjQOOu07K2YmW+jcUORZn
tTU/0+PNdAs8LVErZUq8mTppvX58DFLGK5wh7hj3QDHhPnvd6AVpz/Nkeq/rBwH07hi/Yw4SuzCM
Q2d3oxP5Fx804NTU8wcfCsJ9lzwrxqwG8/ct3dEAY9l0X1oVPycq2a90N8n5jkJzGfakZqmn2rTQ
GWAbhGPmHK8Nn2b+NYcVO1MJ8nF6JJ545NysZp/LhStj6A4Qa5WQohFHd0wslis6cDxeyZMfZvro
UckS6qhPEw/w5CZ96fD52uMwG7q5igEJHnPKYjB1AcX7oJiNoTUlB5wCN4Mm9rOFW0OCC7R4ogSV
0gm3YFUu4VFXhzjSTYPmrLVvPoe6kac5AUdGcy0+Dt4WzqR9RA7nCSF8t/cANQX0TLE9MaFiFef5
PnucAz+RJy3bCSXidWzZxZjLCjaTl6/ATn8AjR+doqn0+hEoTo5mZsHHasI1jp9mXmw71Zy6fokb
sYvU6uszv8iim3UBaZolY3WavykyOE1sSSMrySjbN8IKZzrvrwBrGBGLfp+hyRgSfCEX9L7Qg6yA
avCiH24O9R2PqLj7+LRGrv3bdTGQ3zlarFLMa9aKVHhjXokNl6UDv24pxpbMmghDLezDzlkJyJhd
kuy5TW6vGOs1nxKmrYec9Xr3PHuxfyrp+FtkAxrdEDfMdvvEU0Isrd1UyrMPX4ZdgK4qHneor1Ci
JN60HejlqkzIiRm3CKHpHrB0uqG8egBfY4Q/ywOqY4zDNKbdwEtzY9pTq8gmxUuJ6O5IudIjJzE7
NndrzLvkYZjFNOaObw3J+LOx99NBFu/PVu5biqAY6N4uMob/bJU6DmgjylgIjrLTnAnODXYksIeJ
6oMxjUVn3go8oOTE2+W6RtRkWyut97jezBNOi9HgpWN8X9YpaEivYyU2p7yuYuCIMC2m1Aaw4VqH
w1+HtRL0Bmfh2zhh9FYBo7BO+NUIIYqK8DeuU03Jk70gmGTzUlYbRqYLoynl30GoCVDtvSncduHd
NP7hBDIiXucC3Nr7scidSvQwHjg9hIHdC1xA3QFm22wakMh5+snlSzBMUADMUAUS9LSQGC06WcEd
ZiVFAExejK9dQpfRXvVFXlCNLDoWlAKEo7E8e9YozUJj5qqmvKA2ABTFFTwBOkxnOFmHDjnPhiK+
4KkK+c1jWrkTLVgfperH/AMnL1TZaH4FHmtvKV12dhZQklzoj8SYKxClIrIV/4sEdTzuEkzNmc+f
GfAGj7UwBjcqaS0pma8NMU0eUA5lHTplQKPv81VVGdrdSW5IIA9DEwTAJGIqc3OLIdRfF7UyCE71
AclmoUf5yDucnQdLQ8N7GyYcywuIW24F7Nf7LmJ1RZTk+vWnpQwM9XMcZuXvcPfvE1nRCRtIVx60
rMzy6BkJ+opHJhvN8/SFJuRjiyg2ZpfB1B/OdKzJ6WMYxq8atwneejjqMMhhG9bNhNBcwIrdbW2b
9NRIo4hKpAY7JwMFtkyDgmqDDwuLqVR1XShQK70eQMco6ngNjaJ9aRTRdcJt/9gyLe0UegRbTd9V
mh9ouAqJOn6rKAnoXnjlx/pnxwNQv7kFe6b91W5TWm9KZzGGiUYarvJdE2nbgCSbUJWpdqMdc3Ws
woXQrGq51deuMcCV1X6musKZV4i56rUum7QwS5saPlMOO/VzZFewXrg3Lgycxo/Pv2xnG1NsWXlw
FfjXGQrMh32VJivDjp2tX0FqRYxZILhx/iEw0OEvc4C/TkT8cuRIat3w3Zf9EZaGyPNo64q7JdZE
Cf4hqswnYTicne7Lg4khrPmecEaDQplAgBiocvB1iVtBc7WJaIcGFMJI2x5ZkMpQM7x2XJU6G6rK
MtCHjRQs43NTIXkeEAggVQbZH79813eH+b50vd3+Qxapot2KRR3Y4EwV7x/XpNRUCaueDLuvemrs
edaxRbIf6fAsaPkm6HLlE3OjKbTKRbZ4A9K4qsQxMxopV74bxL9Xcqd4Oa1s9p0eH+5nOKQ4w/dT
70xaE7a0SniUSuoqpXBm5Hi2RNbDCuGSxqPsJCR92ou3li3QumP62wIlWBzhzEnCxO9Xy87O7AwS
3HDmyvhKJ+QnAvHRzs2FndsKFwsqkPcK3bsurttQFu4Zo8CuHdIllEQefw3KFdg9ZpZct4Zulg2Z
rRSnCmwXbzuCXs6YYrG/e8BVH4OaQEkGfx/X0PETOOtcOjSKdjWYldgJYyDng0qYwn98Z2idNxTd
DdArxv08aUZb+uIIlkHHDb/Sw+BI7GxZjVnhBuUIpn5kthxXYZgaRo8zzPop/ar66eQGjZ/dybjA
IUpv+QuL9UUwz4uL7HXBR8J7r3QSWkW93h96gkimjHkxp1v65YaWOvnMQb6dd1Knt4361gYe+7JR
l++BW6X6qDObV5kdjTQozWiZilFpd5V15QYVVLs2FEc+5+fSlclIvgrS5N+Jl1cd0LsbQz3UhKOV
kp8YrRYwcl9JXVbtXVAcE9OEhKhSDoxgw1E8vbjH9+HQbY56AC0t3MnF6tYO4D+kfBLVaqseRuiA
JT0IdrQCz0IVq9alvONmsvj27cE0ppLThdgz80/uSB1MA2koSwUW9WmrbJtYAeYgRjAz6tFXmcWJ
g/3TXHvDi03vK5fi9hglsUHIrX+2NX5nflyBrfvRFw3xy2dNqdVj/n3vqp7RJCSIZNElcj7LJDut
gbJPS+2F7iuuADG91MEi/6/sxPuVZ7Bgqwmb8fn3xtncLip+hP0/rjHgq9SRh56YwEY+qIIlK7sG
OuBn7VEOh3lPlrUJiD8xNVh3LJzQrn1qHvRW++r0X8iKMkcv5iXPdK+QgocmG8q3frItfwnflxsI
2SLilFSbg14Mq5+MKg4zg7QQmGq6Rw8vk7V6DKgxixOmYwhJHArMm3+/DEhFVy9b+S4/tcpBfMQL
TW3tCqsOPc9hWS1XtfyFVIZrjQgqlmPQkQ2LdwpnV8jWwJi0aqrQoSKpR41REt/a42Rrjy43K8cL
IwtO2xjNH5QEwK550IN5XnbpjgTMVNLVsjAQpuqINSRgSJH6sYeOoovsyU03UAEirYtIHqWRiAmK
FJ1j+lMHV5APFjprnt5LF7JIfZ2ilGChe98cRPTItz7A2nigYF6eVIuynJXWInJYpX0Os6uoqeQR
C1TYPa4+0KsvDCRu+pfZHnD/f01thAbzJnsIBVqvf9FFbuNdQUE6+JDCbmon6LwOAEbGyYrEgCZ3
fqJ8b+qSgQ5wEuhgqq3sHn3crh8QIFM/cjQa9N0/BEqvj8ARqvbyv6pRmzRgTKVCdfhWuO3k/2rt
DDI+PYT+R7C6vTzNgkGqztGU2KxR1Pw01z6SWtsWoLhcgSufLe7riikR5dtxxfKZwhFW9vac7tU0
YH/w/Cp0dCYROfkg8z5zIZq6zlua3mM22Xl5nqJb0YJEhMLhpOXrVeg9hxDLRskfFwx87BYpkwJb
ZWtuhMSY6pecge7z/PXok7dhXvV629iRUEkeevizSbhgD23Y8xHJ0ZuffNLU+ffkReXRegZwOaFM
PfMn5Pc60lEfe/1sPq8i1iy5yoboPde9z/f8Be4hs6TkLXVBTQoGQynbyAyqSPONCO3mg8DUmWyx
JXygg/8Dpxjc+uLbl+LWm8RqTqY9ojH0d8yiyMyzz+nC6GYDI29kLuGZYLyhkEBpQyTH1o+lcdrj
ViqWPXklYN+sfShiiMb8oA9j7ZqVtbCsa19nVDeTHJwyZH9zoLBIAoo+bn8PBUCBbSnJzB0ubFzR
aBOV4IomgYJW++OXD5i0ZGrP8hByIjnx5c+Oa5Ax78P9Aea63JZbLiLGh0rjfGDhEok2BPep7Cfx
B5D/qVtFRf78+sn0lVBqUT1v2iy0lf69xqSMizO8SpRxKcw6lles0OgC2wQtyYx+r3vVJQAFUHUC
3ynluxgTtDtfWvSb1XJO2rrU7NZVpjbbjIhn5nbv0kx8qIHZdgXC3BzZ4BdtuS1ZubiaV5yJ2wkM
2ZaAHJiydrLQUmBf4SGrWWIJixDrGmj1c23dIGmPHooFXZEWSnLoJAPtAD4TbH/3oULZl3qITc8j
/edM8Ex6v3iKztEHJEkRI2yqYZ7DA26OeMflbVl6KLMefQXfw+QZ0ne6yQVJ5nNyWnUXimhZ8fnQ
KZ8/7CgTKT3kSpnxbdGCG2fEuRm4NlfEW9Bh1xQ4DTK+IdpjOedfRB9cuYO2FZSaUVc1uell193E
zODmtWGGCd5QAVc8dFVSCX8Ek4H8O33CLZkTK/yp4zE3ADoqE/85HJr2EVoL++tF6+S75uIhSjtI
7J6gzF5azlEWQ3Lik664daTBeyeJKztcnQSCD6iIUsDljAPF3sczbsFFLfxCt99Y0WuZ8SH+Ew/A
sppBaSk37PbHRLj3YAQQSxEuTiori9JATcSnFlJybXC3o4GdhgZBxJ7BZJfTe13b3f84ohA+Kjap
I6eOcrssUadLz9DifMn1iX7qZvrBSIpq+vo9Fk74guCIiwooE8dHKL/W3cXs0i17br/9jnU6LR7o
4BewMCjiKvQnAIAwjcroj/Fevy98m0jezRSU3qEcXC5YFnVku8lB86EXmBj6KbfN662btBjlhMdl
wk8s3obMFyCQfYF5/87yHoHSqmDD5E4qpQkTehZTHHCW1+rd3eJbpq39dWOtVkeTTEy9lst1LL7p
nj9PIPnLjxhZYLrmOwmQEeQmyxrokrHkJl6HmGVaNGjgC+hVh33aQwNvC5KJPN+VHNbsazwDAMJS
hMWPKTmGjMWjtdTesCqz4SxdQwkf/5Nff+tpETIDejPPBJws/9zhzQfQfvzLGMwG3n5wsUfCZpO9
RlmgJw+Y0M1RlcLMcnLbNNG5H1R9MZaby+IPLG+KUq6xnmoNsH03eSgIfhyzeqAdxNJc7i/G7LPe
Xesp4aUO2N3R04yrx5BtBdThQIw+aIveSnI1Je83DvoCbjFrqOQFdrSYrbhxIg403E4lh4Lq3NLv
lX4rHJMxMGXTK9Vw2PfjcIly0brFJ0oQHZYoKngEgakuBLiGVHYTXA+p4U/N3EdR89bbWcc5JT3h
mohS0HydTFViud+dxWoiHwF7uQAqP+44VmyARl69brL45fZo+BTsSoWXbTSsVJW5HkSt2OxuqbIB
djHxVm4Pf+lULNoHGP9q9HZ8av/hR0ECH6+iQEPlX2LhBmBuQFnYrkPBUWIkebPVWiqEM6ZoqxCE
yoqcquypR+449JyuG+ROAQP2dN5dZPeKNqXwM3709KNg7fhnXhfTCd8sSowQxekYK5/jesL7uUhf
sOtAPE2ehWfPHoJPnFPWQW09ySWD856UUcVKI7CPj57WSQmyvZq+lOoGVmDaJrEQ3XB7etiEs8B4
vcEN5QLhD8vuyh6zEtp2pZGHDLyBRZsnO7kyXxcn5RnHTGgF3kKiKhSFdI+iihN4H9EggMaziOqY
LxD8u5wTnVAOGqXkS3zF7wXVb/HW0rw+FgEoBFHoJFKtF/we0MJvE/+o0aJnpxP/s8Oyn3s5RSaa
J8MmU6sbnLULVWuDnGXyIzld6YyK46X1sPzrC3nTfJq4974LAl3AmjZP5PZtu1Z6WZFo8B3jE+64
AeqgmTqrpDY2c4xgQJ7UXTw5vic3p3UBusvn/PZFaa5ns9G4FBjPJBDL0VXgW4q5ENKi7BL5NJWp
QNYfzAFYZ0xWebzni6GFKVb8onSCI3vSSCVaYUHLewxD9peAK08TMpmH9FoBSGYZ9yId1XeB2fE7
Uxg/QdcRt1Sz8TNRH2vG8IltxPmlxDIStQ2TwR6oobh4nrzUd1xWklDgy4dfAT9jXQyalW9UryB/
+E/XkD48wlPTH6eH5w8gzxwcsRyzhsrVNi+WDDCCjVsUlHwCp5nOiretyyyTCutzE6TTqSfqNGVT
fX/PRXm23RcLTce5Mblby2dzrnjhnVBR4Ujv+QHINo3AaaTlLSgYC9YR+TL3eQrkl4v4+Euxfli7
4qQnjrJVzxWRzRYFvwtdKRyVgXQG7cwfAppZscdXqgAp/TxN96VX44xaTr6dGXvcIFgc+8MC/y4l
aOT0+bNT7nBMFpw186Lpklx6Ma0sDQpA+RJI7rqCDJ9LyzO7nc4gJkynSjyyxHfBYKebj5f/AU8+
fTvzsgje6hvyY47JFtkMhOkb8yoBvP/leY/c2PiFNC8Xtq0vIpNDwY9JkGn+ydrnowmAY+3Ci2+0
vZz4gqJ+tn23/9hVBQRCCsYsrhqjWq2MFEoO342zg2ULAg8E34t0+D8zzeiEchiPQrGgHE8XNhzU
eJ6bt2oplDhOxZsF+eQv+Y2orDx6Ig+kKO2gZyHJvd0efYHv+xfX2Vvs8OIQJImX+SCZN3ZhQGY2
+sVmM8WNUn80h+2WoIUA1YwabaqyZWwnap0Jhmm2y4b9bgenLmwygIbmHjD4pLc7cDqfiUQziyHZ
JfMkMOzr0EK2lis019aeSBDu3/0r8bvjmUn8rY4NWus/q7tS4Ny+fVGvgT/P2U1pHdXtcrlGY77W
J3O4Qj02two3HlblKuP2rnIm08MnRSJjRmz2MbcuAUgf5IsIe10fl4clNI51yUv3Ffqec09E+BfX
IvPzywlN2MHjP6fNAmv5crmrCusCwtS4L8klEEYdpYaGC2M/9+g1pO05mm5ilDKOeaDlWvjHY0WU
KKMDuu9RDXVe/0OX6n03AlEwAeZtPdIzs3L31PluIoISjg6O4gkJ5+ML83QvuBzHp6Jpq0l6Mod2
etOEJDpIeHfEhji3LLPzawfoAOOlMt2X2IpSmqxwK4JEX6/r28OfRS4NHMczZkuz2we0/8d3QNs7
j7oiE/IPWypg0WaGORPZNG+NGs0GlQLIQLIvIuwvpJGvhGTMJZLgQmZ801ZQ2ZLc9B63eYuGkUil
eFnOIcMCev8q315Zv+zIj9ZQ1I1Jifh+7ZTHqronGvUZodzCiwN/9yKtbZ/ZceauYketUxCWYybE
kEgfeVajcgxcYIoQOR/wdK3WR14B2iSvW4eW2e4HVTxcWt6wJbQmlONO9J1R0ESiIOQgtU8U+zfU
0rjPAEM9SloEU2YQnC2IxLx6tThi5Jplcxys3INP0tluFrsTxwkOPhA0CwFQAOeVKXjK1lRVFFJ5
eYi+9hvLB/vGQ6vHtp5nW8rt28+KFnfyNXX4z5vGY2druo95z3FMMZamN76+taAwHN/ukz9xnjiS
jCKJNMtBGbTKfU4EyIE8TghTud3s4TyYpXWm8DOVfvSjKYOxH/AkUjAxb71VpHNG44rX3YbD1MIj
idcZuEujxky2sjnyc2v9QQWvszeCBA2mr1HpYaDZ586O4AWeUVlH95+LaAN24e/YQ93lBcQLeYlW
a2hFvJwGgY83/CDF3oUE/4ddYAZFcGeRqBqVGWk4uESR/BG2wYYRLujxlczyxO+fSAYsazQijJXV
0O7u7JWLXzozorvUwKjylZrVV2ofvjByvAx75kfivkWGpH6alVt8cO+RFEYf/PKu3G37a+PNqNnL
lNqQhviS9O06/PyF5jh0jsUbffPqDJkNU/o/snQa0L5WK/52q7TVF1ZOffIbZTYZdCRnTlFCGEvO
pnbpM7mp06D5I+FtRD+KwHIECZw2kLFS3lZzgNqVcKre+trOJ6sUIZhD5xkPC7mvZmSSTeZxwyAs
eUcpX8b4qzr/5JOB4LE/LGxfjNgPXOpXmmDNzwwiQPEtieb3dPVn0KQ91Zgf6IqLjisksv32EBRy
8lm2YovBKWm3P6Lci92hKXZ7+tWVrz1eXeJzKEXHePjPZmufqHU8xiIDjSmDl1yairPaIdNMhaNp
VbtymIIlcceelUVXmUrLMp4XwDQ4y0xXciyHb6tPaZEwkJcYmrrtbRHv2ogf8CHUdJxOyq+4AbbZ
XgWUS08tb6KixBBGuVMzGSt4vFkE0CNiHAv3Z174A41A0gvuLEMfC0UcNqZCWy3R1k3byIJlWXDA
HldvD5VbtBn90UvR2lXiIGTLEPovLekHLO5+d7JQPSN1IhaRJFS3YBsvIE1Q2UVWIW1m5RvKctVE
e++6EgxvcqP9Rz6LBw0VOVolz+IC7Vz/MOFv9E24iuEo9/MdrQEBVvVeqwL4Rclm2ZSybBMaO+AX
DRweShcmRP2EOfyue06PDoZwcUQA0LAujE2KPTAB+Z+2bore/mWhhzSSRRVlNlFaggDFMU2VWCZN
0AYxHVROJ6KZlW2rNO7BCwgicEcfTnxfig4h8Wum00SamdpJ62Q1209MfDmex7DIFnci9ZKmUtRq
35HmXOb9BPTeP6SQvcVfluBWbla+1+168de3LOkbLwnG/tocTRkRBm6OQivv5BNgih9zMK+RlEEr
P+2u3lV303SGc2gfvOGJ3M637efGlb1LTwZqHv2v6y5j+43sSVSR61FoDKRK82Gdvl3CWMZ04ZxX
KmfVLVqpVcU4ucfcXqGSzkxs2Vxcp+T2H+CatZqMkme8TZ4yoByuW/DYmqf8QwkF4V9hZErqZKR4
N8IQ8A8KlYiPaEUQzd69cqi1Ckx4u1NPpmj73LQPCMoyenPG/Iz3bQAutwl9l4CRLw7ST4lTUtB/
D2PTNg77aLavojuQ63zJjZ6zj63ZgIPnCInI8lIKHpP3XOs+zI1EW/zcjGKSGPpWGCcpl9hUUlvg
YbnyKA6AiTgVGtJz/10tCUiucw9cu+bJXs9884Vkgw6z/OEJlyJTmlaHTHn9bu7pK9YA8Z2MICH9
i1zHyqMtRDho0L2Z2l89IUBRukB2bVfLFQultqzTw3/kthgAEgouXqKmB5skEPYcUe+HQw7wwrs4
W1UKgBfQAisM42CIew3t8MOy7ga3hEjrG1K0xhXHu7+wu1i89/8wcnPQWU0xzG8yfix4JiU0m/VR
9kb6tluvXzXcnkhfmw/mKw1PV1h6fE01nJLdAmFGMGzChY1FfgoC/fQ8Q724356gr1x1i1qVqWdA
XO6oNQOQWunnInF1EAPI3NXRkgAajkpuPFQ2PvQNutS+e7aF0fLYOSPQX340sJ5PW15rO7mx4idc
3qOf1kg+GS5SjukqhHSM0ytjODGzoR8qNjm0ujDhJeAYlqdISJGYagVyA0+pvm19OQUatXfStld2
oB6SBR4vPIafloKq0riM3h64vtLK1NJcQ5ts9jsJi8BoVxDMjZoDsVh2g2rs4q5yab5c7uT6laou
grR7j7+qSAlLb1l9dteo0cXd3LPeRpsebnpuDh5hVTtra7bfaCowjJTpw6THXtB7Vo0BS4Ju+o57
zJGCj6XOV+Ebh5myEUv96Y0ykr9CXoJLdx/U+LuO4d2rHRAvlhTWESSS3psABuAnR8HbFwN5DPzF
ob8TwdEaq+FfPZ+nc8i0L7AQ0iq7H2/FNGBmwGZ8Tppey67VnhVET+2IlzsSJgAoIxbHjbW3vrQS
H+1DCZrEylvhH1eI2IlXFyL8TT/c5boRopxbl7ZOEdZJZQdjAFIV79OyVAAZmUvN2d0bWpWhARxQ
zJ1wK8VVjkUOQpi9Ye/f5xcKF1LtsAIbj9vUZCcRrOmuSOaF6gySe2wEGC/H8OFzu8zk21yZqY0W
54qgLVYxZRAnpwWJ6bm7UUYuDiW9VpCmnMctRHTS4Hcm0Z219BvQWbQqTUCNI+xxSHi0eLcwFyMx
ltpAs0QZ/Bv/2h1MBQ8V7qU613Q3DLgyuIIwHChOG5mb7v6tHy0aL+CaVM3a7vvyNvPTH3DqtATP
sYB05tSwli+CIbu3YjLjDpqinrDhpHpDEUCbucLhOFp66bDRdvp7BuK57fXwBQJMSyEjEdFzHGCt
fXfjJbyiqtZUUIkLXIwZib2VaOmiy39qy0pO+zRpjATcuyzabt5TrE2TWvdDvrxxZvszx8YON4y/
5eagfHkp4lZ8nF/ubSKeyZ02RNDaxm5vyD15hWqE2UbWG9PnxzkankWvftB909atLUfbjsfqazRB
O0LAHvNFB7yh3tgRNwhhlpnlwNHj0597OT52+rGRP4EVk2SzXpzTn3lLgW36kBwrrebngHbEhg+p
B66Sa+WzwE7q15wcDPL70Q22SC6aRQHaRFgpIxmXB5q6ur66YR4eAHssER0kll6g66Zkt/59Ymqc
dKGcdZPR+f/ZjW6rfoOM5Klj+f1jUYdioeOrgMjFKrYJv7qU373ptENQz1s3hruZ+4qViz5vdgaE
HIcCwnhwINnDyCP7whMNJ76knHEyB/bRvei+2LtvRtW8/xR7YKmy6Ibbab2YMHKqX7qCAOsuZ3Fm
uASFxqiLIhq0SfwOvcI35yLPOlFsXA2MzZk33wkn7ruY5+dxIiofQxp3dURK1EzDtTYhvKQQ1I7X
YPEdR8r3oI5ls+dXtOWUP0cT0mwGgtdFRPzMrumEXUSzF7j9hZqvXXpsMR2oO5xKGsbSVMDLx2hx
6CGoCT5Nes45OFvw/xsOboh1A45bl7KL+bjDFymb6cOFAkN04ECFEOCGxEIKmo0TzbZbfPnWyxMq
ZeSe+xRTLgAuCH9yw7gpOIyWJItI7oy7wzjMcbO6W2EzPlNhC2uaCMFqcRD+7o+vKdSD8GRhebTu
hjJvaKpUV9c2mGnS2EVtk7aeTIuZbMZ4Pr2L5c0vkBB0PjUx9V8zNN9nG4aVAVR10b1zINFXcEzF
7HDQypWhWVBXdZzKr5NyZ05fUiUHpt5VWVEYfz7miP9M+Wu0VhtjsP+Zvw40+lLw7wKYQzypzs2x
8DLQ2sBfmnny3iWxKCo6o890fFKM8/G5BLNqt/xcr6nxi7Oa6WliCBwD/Uafg4QqjDiTsz2iwwve
M9YhTySUg+eoa0B1VEHM0nl3oi++SmS36qnaUmz9jXjQbEiPIrgaQ1AqyP6aast9W6Kz3u3xBoM+
vDbWd0i5/7FsvoCF8LKNiprigBS5hmCTjYQYCj9W0kGWjvuz/70eafJIT53MsIRwlV1zDXQD/uiu
YYnkcyLWF1+hTb4cXY2xPWa6wjof+8OykLN3YkSlS6y8HI4aMnEG7b2l/siqd+S03ordvQgbav6a
vrdqB33PIVzhkCG+96pE2+wnFLHM1t1gIoxv1dpzAgb82sXo3jioAp0s9g6LnyMo32MnrDnuxFvg
0XFtkv+Lr3FIpa1eTSLVMWoxur40sY7KG8czadP/wSbrrRzCtm1RlEpj7ibV6eVzW+K/TMfFgIzm
QihbZfefNuyjh4RHT3Cafr7b1JsV76mV+DZyzZDh4mylGhGE7sAkJmppu49Ew4duZ51Js7M/ZnUp
+qKtQONOQU7ud4qk9BbxaVBnHIPG9458lRuhl0XXvRR178cG/qkhhjIaOGVUZYl/dCgBD8ig9OQq
dXYuESPPAtNpMMKETtDLEVx3N86SxPfp4chUiOptt8eEvl99VcJdA5qDuL9oJU9L12NR4ItBGhYV
oqKTppxStbSYoFlpuzv966tGzmDeLE8GtfaBEVeJ7FnhMMurAiKWEOIqLEof3wLCKpaJtASoBFVp
1NYI4YkRlHVaoW42+rbO15ei7gy2oMcVgzvncD43Xvcc+nJduycLmLe3YqNbs7dx4O+Tnleea3ao
Xn0cLi5nroZtuwrrRaQSzSJlHv2Qj6cCETKAt5gfgA9/gKKJxHjLBnuHyVPSO27fKatAqiLQ4lXT
aZoLc7ve2xAPwdVnP4kBZSI33B6sb9ghxyootpe7+wul1y5MOKMb6UEcm/dC0CxiRQCXnKaBVysc
or1mkb38W6mYBrplHbKjIU66FSpm3zHg6Yklym41WUycrzc0n87D9fRSYLu3usCD2/9J/t9pI/Z4
7/j/siVnSOloXUuyhBd1is3/3VrgEUUWoWZAII5JBA60fS1jHwgMpkXctZFmf1VcryP8XO7EJRir
pHFGmg1Fy/POSt0RUlkHYiETvSXEfEMt7uDefsWetNj1/qHyZIpw11U2ssR6ZJXoQddFrJlSNVRn
70HkED1AvulyHFU/1Cn3h3kLfPujWNEGlztImgQ3jx7AgtpYYUYwyHhC9gICP342vLQ9GjZ61LVi
ekCYTbPlfjc5NsPkytJmzbrRCPQf+KZTgo9fjC80Ds8/FgZnI0r7T2qeCSIEuwsPM9+xiITYNz9m
mjcLIrqdOAPaCw6VbikrtwHYYBTY1/Ec8BL2Db0YsotFLdgEi6aM9imp9WZZFsMaNTPIbafajwcu
mQGtHqfo15kX4oQVT1axwfWnLHuXVF1fTQEmwqEDERx/GlYUiTCJodlclMAXCiyYA7Sx6VVn07/d
Z+23ga11UP+qmCxd1IeYPX2h9RLZW02UW8yCcGGxgIYSjDjgyXqRDT4bHYIkRDNRjBTn7n026fcN
phzjDrw18LaSLe6BM0eEnLntF1A2dULzksvlXE0vRwrHPDChklzdcphFhMCAztD2M/OQJz3WtuK0
qb6sls2Q9N9Z072+Cehzq3zF+44/ZLsRQHTdaQMAuSEL5Dlsr68IQI3QFbb/5DKl+uH8kZ1pVZtY
chK3uFc5raJ2Jr8Gsau+PXzsSJLsdQ4s21saXsE2nEAUGWwbgT6uk1CbhzKPYHLG1yBy8EBVBygX
evSu49YE8T79ziELYiisJTW+N2N/Tte0MCHtXlBqhxcODzSgNnfQcIMytrTWrqsU2L19XojyfFCx
d3YOco8cj26XIMIF/y34waxhO7sJ8hIFEwQddea/YzaEEygcqFn7DetC9x0hju+r3zKdi/iyBjNS
FslBty5VP59qiJZcGVTA2o/Us94amO7dxcroQiweVFEu+BicuRWj/vEuQlkYkHodhe/P2j1+lqwQ
z5LfwzpJ8XOOhXaieXBH0Iq0GA9F7dNxkyjAgBghNmFPrdNvhDAXcHia8pI//LJRhGx2V+4t8qp1
/CscNqtxId2Fk4N5lOWqXNUS3W1IN9xCuOAivslf+UqCVwHiaoOtNDnwYXKi08gQRPdCXEonuP8t
XdoIGhH/3k78ZkKeeHKmSro6VBmko7olMZA+8C7F5l0beQQjQ87uubXTsxrRNAz01HnwrgB+asAn
h0+lSrFzGDqf7Q6B7Ee5kIJlISEUjeffS4rHzOn89/+J+0EIpVKSO/tVyLzpbqRRn/zxuU150aEP
+HRkeCiqVBW5Frui3Wyy0gd34YEAF2Xvp9XYxa/doERwkP2tOdqmvCzRkSRH/+Ky1JlvGErap452
DOYU1AKYTGYGSSceCJZwvZpKCTG72LdACoJK/bzqkuDCA/ZxMA8sgkN60kREAhagcXtQXbWMPTO9
4W9E+rFcrf+bnHgXGC5QZiJnhejdtBp+WUiT6slSRbemGWoUAAz2Vv0ezDV53Q0lcVAYe+uSXdSz
6WIXXyy/m6zEG0q2u8K/tLFrysMASDFKBjYBno03svXH+Dyjpz7wUGYu+/8ooFbq6u64jV2vS3fO
nJ25j7OLUGhmOSs4tGofOPLVmexdCctgoTOy/IUdpE3d/sDLFz7WPKpmU8PfvZnEMDZ/5h1KF94g
RuTlRdNswTDJOeCoKaOs/yBu70Q392jdMn/1p34aSmkFWfyeNwPURdunrhPfydWvsbGkTCT96fe+
xvcVRbHIscFVcjjU54znPEWA+YaeNqxqwP+Leehoqy07DmuYTQLX6/jYf0hyMl8f8bKIzLFzLrLZ
7B2EMqSkgOBoXa216QJJgbTTQ+UK+uV9TPWdU6G/L77uBLyYpfzLWro1s7fVJ6hlTlRNU8qtplFf
bFMFINzf+PTS6FyIvvaoxcCI/juY0xmYPMynP/Hdtwc8SsqYnJfen9F6pTmEbxBrIqoOqC3fi1IQ
PWG40P71ZWH9D1w0BOoXOoIrHpH0/dKIj85pPjsKm82WHt7OD1gm+mYMBIpPEtSh0HG4I45bE6J4
nGT+HWxWNIUJEj/A+jKKhwMw+NssHgWMYQkPcNPAGtaJTdoshhaDk5eTmPRVl/kd5ki1+wvo5hgF
edcQLrY8yD2dLO13oSO//kGBq2/sw8IMCMn3BuiPGrhv38Pt44hkcv2I04YrfIFCqtwESMzt3yKU
7XXrcuL//nxY7tHZtgs/+iYlxBrAi9Fff0WsFC7csqhX4ppGDpfBdgx461a5R6GceQlnr9iBwZJ6
hHkFYSujXmqTbU/GEpCKv5oHhUFhlhe5YYSMkyEjKZtK62wygBDEpEUBGappWCEbafoC4gGhdcmF
HIDkbfohY3zd6oEwxArALZ+maIlmI2Hmb1V5zYklHVZoFaZgqKI2n/7dnIHPTAEcfI+cDeAmy/8z
8ECxWXLAurnfhDSe3hWAdIv5SFRIc+RAbAUi1jIYmL6GdN6hEgFTKZNQ4+sKj01YmzZyMc0RiIrQ
apfIA/V3F0GIvXPeHQfWhC38C37/8tAE8l/pGODTH4q8xcP4TnzQmb1nzElIP7h2nSHT732zV4d2
9a/d3E8JZKEdR9sgwK0vF7/mSF1fS4803gyWhrPfJuqqxBrEqgtvavMfxm4xRSjv7bgVgqKpyVAX
ZARF/+Kaeefl7wyqV3NmkKrGHhoVz0Th6oKimQeleyrYoQq5F3tpUyLxVoT1MZbd4bmGb1eAxjzk
ExM4KW19pDglYQwp/Eeh0BeC1iPXzgoSI3bvZDfUNB5yLvo3hgy7BwjZT5tugJSShevmsSFcGluS
hAH3zdxyg7ONOoW7AcDdn4JZdWOBgZL5scNcVeW4w320GNKpVEriHhXM0sggxTaHMz8/WC4h0aCg
zrONky0NspyqyG3MWM06UFjP75hwdbVqy1WXSc35Y8vO9cEe4kwVnRsoLk7eAFK6a1hU9T1Ugb5r
aIZ6PJAzGzJ0aMQGDAZ6WKUTrJozvV3aIWI50N5zBDzZaB/GMaqq2v1WRoKtOZmGhxT/5kF6Q/1w
38/VwuRsF98IeW9ksM6kOYh/ewS+WRNlImANSzk4h9jyQG1nqi3bzV2iRH01Wg5eq52oen6Fqawo
oN40crjMYVQ04NGyAZ9h4m0Cdf6pEmtNk/SoYwU74nUG/rV1AcsLaNxSolI3yj3WO4UxtkTZxYiA
2Fs6dAwZUKhcKkOmPVt9As2CebBuI5u6z8zoj0X64Rn0uzxioDYqRkHE0ijM4JddUaurmK6ZxWcT
kQaFcFE3Zmx6rTMFgb68zw/pic4OHxnPwVyqrV3EFS0q30cqK3D6YhF8rzWzV8NZyDpb2iYGYfXM
+PIWe3eAn/yAzgJbi2/MnwMQmJoE5CsU1hSExLINWtSw73otPJzPkAHcrhkuUUGSgS/RXPHhy7Z6
SAyuG4v19gaWbisEWlrydPG4OELRrtJoBE0jjxYHY8IqTBK0J0cUp63c4XpXd6QJ6DCUUrE71NJ0
Ln7Zc5qB+hDIMF537vVka6d3H7iZckQmJj+A7893jwGtr5fKn0i6DQ69khKe//0sQKOTnCd53W7+
HEdIfej48cCzDaTiMzKbipzee/YhieTe1HlB8xN6Y/+29873hyOLcd0+1HDifow+avPsQYPoH/Pm
Y0m1wXW5wKuul1oBAzr/cyilnvd+2cz60oEFyGCvhiZb4FoDo2hAqBlZRHw33f6g2w6BbV2F4XQy
9PWWkSxeXnPcg2cnolrto//DZBVxcTwJELbTLD8oQ0KEdGuYuAzAUTdID4yYHz4xZJV0XGLKhqxS
w79WE+zwxSCUNnQGXHRsC29ZLrgIqLBJQazlktupP6JXcYeieLbbqMOzNswS6SpVDkMFQVGVmefF
TVwWHe3RLpMiXjc9Rdn8ryNfr29tFwFpNMBYG7Yl6U+m+VqL+9DKLHiI+3njd0B2xprKIQLIiLWZ
LI9DnAf+/+J9CJEncMrwKRluMgdTixkM5hMBwkA3WWPLgkdfUAA1257+EY61z6wInFoutPpa+FdV
et/9DKpFmgVWJTZXcHMXj+CEpfe8tINEKfBDPJbgjPMybqjViIYhvD1u56OtvLX8o0eqslt9Icjp
4lkHIvw++JjCkbTrHE04OXEGcgtRYUSIIn3GoybG0DuJ5buYyiQETCUH7Q3iM/6KP9zWp3RdcB6/
WjqiX42FeNoOJc2joPD1n6CSYU2owwlRfk2/MVuSRLgwKYkiZJUouG2DsdBvRaWZKpTpDh7fAMDb
mcqpajRuFKcL9I/nPdPqMJe9yZ+kB7wNdStna9hstlK7Tp3eaxW+o89H9zk3h7vLXFHixVEhn+BO
oQLHPI7HH0C1yZr8pCEIR1SniKrdqayQFmYaiCN28uCeWImqlnOO96BVPC0To1U/iqrAZ9OqkS4i
JUYo0druClwt7vf/2rt/EA6H/agXHHl90TQUErQNUHb5EPmJLUb9frJ3FMtm31LyOK9byZAAX0y8
1KsczrHZvhnHGyAHXkXhWZtvWwv5VWIFCCr/R4wsP2r+yfmf8bxwgr1g/gsGsUqSw3MvNLRDjQdc
g+zl8cvPFDJIEf/8C6jObZiutCbwaYJ6s+lQAoOSV6OmsnZLGqLMmnpgwij2H4Yj6fFx4bPdmUnK
AM3Kay0EAyi/Z28iGTExOV0n5khz2P/bBKIi+qe29Z0VzypZ6PLayM0INGT6fovXdj+nfqgXnpLw
wJeUG4aB9T16SQeTYXssJxZfypA951ChX4f4/cpm45YfacDRbKUzoiiCuJROagvdvCOCHcWJatrj
K1mp3nrmdxoq+8RWiyx+d7YIfwsXIrEjKXBEM8ixai4s33YdrSvoae+qZZHAlYJ/qgkaz0CEBRPu
W67Ay0mMd/zk8WYKvrICUoa8HxgWp2RAZnfddeWmlpWnWkSarFkKGah0irt7PZN8uq8m5+9PDIbt
peSSNBmaBMp5VjHgn6IyuRuJcd+90tO7CaW3r68IcGomO+i2HhMQKxWWN47xwDlNigWEQPwGON1R
TykgjCakUupBnB+f4BxFq3H5POmmwkeco44ph0Yrb0E7wTO+UlSYH/jhfJUIJgRIKaCk0mjcAnt7
tX3I5JBkF7mqVCwdKnSFB+jlyBvkUnpKF3f0ljiB/GZ9trYF1j5tI0SWfBkg8vxF3qz/BmoJjVvV
88FHUwXWbg0S6INdx09AKdQki0BTt+LMc3CQHAwPVv5V+32WI0fYvwsKkjRYFecsvCVmrMvqkiE7
xZxJ5CqzKM2NhohwqlSq4lcCEJz7hkI55S3hzwnUANnG7aZJeIHkflsyQaS8+LRyEf1QfV1lpc9L
rHdLBkenShY/t33hTuHG+JGDzl/6VDp5KXLZz8Ju46RV8EahxHUD1W7j3FN/XL9ZEdHh6Kd5UOIF
jmtJpu9acUZzYtRyKwnk+nXMOh9+gUjucWxcMRKyO0pXYdeHcY8PqzZw7sMrlAdj4tYp0WHce0+R
SMwS1JRPzGZfH+jBSRSpk4ig0XAJu6TVJG8Ld6F5zJL7nkxuNHb128i3wmbdoDXF/MAidsZ4FYqF
GLz+nQEmMFcT/lTeutQZaK34869UBhlkxjiRE8lBSQxW2LbkxhyNzweujYNqsXi9zl5cFkiHCw2L
4pjQdXgBzgmu29SGYNaquR+PdaW9yUePCaioQgoR4NGXHzCDQ30pGLJGRKM/+iBrq1+tB6TGh/eg
HIr83kgQLPYUTBRTTkdk5597Qjc3peJ7xpcwI7J9W8sUbWXSRoJwKAyH86DH1tScXwUxndoFzEXz
cdVaA86CHtY7bJ+nKAwSc/BoIXOa5TnrMj1MrrcJrhenT+6AD0/EP2viRYHk8K/OzWZPn0sbINDY
J/UA8e7XH1uyeJemMj6fSFUkEDb9/UNy9KX5pegNoZbC36bw/mRBkIDrdCwKa9rT8tINb+kvwRaO
5ictzyXRfPkdjBCDlC2BEjVhOcQ0RJOjfCF+6ZNaPQfAQr2RNLSydmgNvvpRRiBNIXffomSj3RqW
71ArgWWmANMX6aD/HHjiLEann0acnOu0leyNrPnCQfEWzT94lyrT4A+7vnAeVpbG/0fHTrBYWX3k
a+h40T22Sa0YTJKhm4mP03zc+qwYpCWqZ/ZRI8OlTVPdJ1nqYSND7sCxKCEDiR4W5zcNoIpGF1ll
iaD5g85M50KtIc8EYzIWbLLd1tH7y6fQRRIP27MoR74DWAh61Q3WIEAymxIpImRUnA0ATa96oR7Y
bD0CfLKG/uq/+2JlSrNQGY6Hm1pFZBMTu0cQMQr9m1vjvj1tXNhCss4mLgkO/Jf1liW+7oFQm4O7
pI22yNVjMyEQtg3xSMOW/DoZIs+K2P4J80ETRu+cGNlsxnJRN+wadIsI5jxTW8V88P7G3kpKuTVX
FI2coDSagJl8qdPTDAJd9WdHgFWtzyKS982elGrwR0wXZdubZqwJMOhYk1glgpJZzYV2/U8d+Dyb
TWQimYnj9xWOgNMmFXfn2dPweinHJYjcicKCt5HCOBX+5L79B2LnRD2IqnYDaEpSdob5XUvjaYYK
xk0qCG6YWUolWjj1sKpXJdLC6NHdcP58S8J0swZ5+TaLcZGtMSNBOUmqI00XygLVUxyN0fH6bLbM
pZbOKboZ6TlwwpA9OS354df1uCcKkdAx6f0WS6Te7I81avhwomXqGUFYonLaq39SRVRA4wAXTD3h
ag7W8MJpssI7mB+mJMv7j2AgG9sk6aCDf1f1omcLM8XLtDEUi7gnavF8HomEMQKV9u6xrfeVvCVV
gr79Zta/1i+v1KEs2Uffe+c5JhDGeOR1I68maxn/N7W6YgYFCb/jWFtXcgkFRxK6+6UGE3Nbs4Fo
ZmbA/Ojf+SOxh3NBVmiuGcIylijVy7Wt0zEaGGysQRGDJCXiw1uce8NJfsicVruzqQwTNRYIEZrT
MstlgF3Phsba/1ReXl1vuncPI/9RY+kQ+mg9ld7OcqP9pUqTMpD2KFg6zzJQSDAEjaBYu2//pqfZ
cVbwh1Ezo5KHwNg047zQ1hVKIuNWcjcb1Siu+XAKCQpab6nvOv4gcclO9a+YP7VuhMgcaIeN+G49
OuQgGMivvcTDNdApX0hs3uQEIesm6r1vZo3HQkREv3duRpyHcUedbFvcUFcON09FuyuuNyB7dE4T
7fb4pAibPbymcy4lDvzRaEPWIu9MizF+qKXmsBDb+5L5O2qE8aJyEdeqZkWBHuQcJblAPd202Ze1
6zVHND9wptzcSJsv2p6dGC1qQjzTBXpWSgMo9ZqCMjA077YpbUhRdVuKX2ZLlR40U5gtsfDB84jn
E6krAK3gGlH+fCcOyiz5GMkU8u4igXpOeenWlxq37QhAl3Ni4+Du9ZXZ9pqRGmDWwkvoZI2U2V0p
4yYVs6ZiOBfy4A0lL7XhxOG5XRHc26khgc3bjGPznLr2uBNBdO7r/1ccMYfHYs1N8p1rNPcnBjj4
MOJxdyx/A5I/Vvy4mxa2QyB9qTA6f5K1yrTfrk97lJXN15y/ZN4UQdN27H2iq65y5CzSftMKgQUk
EkZkenfwdqdt1ETFq2mx2HXym20SKdbSvjOe1aK9u7an5NFvCInieiTtHOnumZwahAkS0CoFH0SB
SNkcxExRWm63/V8A1qXi1tMHd6pqZFa3eCbPRTm8GRidz6zxuI85jWtfWpnrADxsj6oUsYKxVgiP
zlWhFAZOXp9L5rkxzjlvyf4LAIBkXk4zGcN6U2sBXlMbe6UOgy2mSZWS5xtnxcy3tlidGQFuuRn9
yzBpgxoNtzSIS12jy0e3zVJYvpxCvZMyYX4Xef1z+/lsruoEIc2uqxIWZcoOCvBRZRnym/gTXM6e
Mpi7PG5xCQEwehyh9v9iW7fW9Kk8gOskEIZTUE+k13PgqlEyO1I/VUQGH1J8CQzC4irwzoXXsCXj
OLi/j9y4U/iRqBLQHpomwUJ0h4s6N1yXmObe1JN1JuaNKDgBYSOUPYMLuuMxzOcgPbODHCy/yxva
QmeHm0QLFj6U5nJ5JAO2wU0+LIfEZewpPJRcobXUK96NFU8c7oKuthEH/xgx02ARjKwLT6vkMkio
/CZ2Y7Sm6rE5FE2v9fiVgmYPGbsq0kaD5keCW0/N/Bt3BgQ2Y/m/UBN5QfvdNgyE5p+ea2n9y0kz
5ili4TAWzp33JW9MlEa/Rp94stE+eBs43Mv7Pl5HVk0NMBrP6Xh2uGbgtvVoc4IowLZhJeFI2Yj1
CRDXym7X8u6MNWD8chCIY4GXHk+dAklUy+UYu+5mlDqqQ3zRtkR0DuXTUAj43lTeYRdGH2GL8qP4
yHD1Gns5MZDezWOCz8YfhztzS6mo7dI33k5wFUv5zWlvSyFPEph+DSV4gwJpKAfK7f+SNxbTXme6
o1dTZGvCGzgk4nvZgYPTz7PTus5wq5GuKt33yUb0GFmozSHFkMFOWLWLqWyr70wFtonrrF3WoRh4
MnWvnrW6me81Hvv1BzW6xYYcQuAUAmmtTGKp92asp6izU21yiAsxxJe/cqUXq1aLaQy9C/Kx/H8V
wMafciG7Kzgv0TKSCygJvbzgv2fZ1JTq6ig+/Kok7ltIYtu7obGDWFvoT66xWluvYUPGKXiT5kzH
IWt00eR9FhQjcIA0SCnxrKj+7PqX7gx/LxDY+yRynG3iYQ3MjSLSIo/NYR07dGlyf9MgQYEodZg9
28/b1XopBD6Wv5/bIIv1SJ6lZS/6wjKjz+mOgxVoFXfTtbRtWWuMoSP58Ju8ejgTawQT03h3e+5f
HKn5y8ezV4UG954MF8jbw4mwnUTfXoAsBvu+KvGVBnd+eQmZW1S0Hz/vIQcDZhkpeXeKrfVTlmOA
AP3cdYFxF32vqY2XU34PcO18w4pIz0oU2mfQjFD2xqpZg/snluW1TNSt+4VK7W/Dk9oGByHRvksO
zqtTSuVjhT6ZUGVXHjR96JxGDUkXZ9Pfz10h2VzaxnEofAFQr+fDiXq7E9Ktn4hSOgmK3vZbJk8M
QwAt+6xbcpZcxuFsYMNeQrngC4DCHmMABI27VUSpcf6WBT01zs2i6nnFw8t8KnJC8LQSgjjZcDnI
b51JDcwQDVO1ayEiriOUaRYaBH+CAiqIUxzC/viItIvEsW9YebUhfCioLpraCXDi0YieRHIe0XUB
xJhrNKaGjvJ9Zh2iSM/4CMMBJIkla0gwvB7x8veClyIAEctIIXZdqv2DN8jweJVCJwVQ5FaDnHP+
2Gd56sbi+VOvtnh9tAWeU9Dp4KVYzbEOYRy2lQdIt/i4zqzvj36j9aNp0xFVWye16LycGUXK36OT
DTKbhLVX1jeV8OpIu+bOOENmp5+AGUnUtPdPpDa6uGsNVAqDLOgCT4J++9aVAcjDh49c1smnMA09
gBqPAaZ1JapooBsw9fVsB3wINtaKORHrjs4K1tL/QxaRE+1HjRSwY2YxjQUkX3UP+2mr1qBBiKQd
ZLfXgwjioSQ8J6dcMPLLqoZ6MPDLogFiBPgjTr9VI93k2ppopvJFhj4wGI2gFdApv/WKq3coSkIR
2pIaO2odki+FjzDl/7EomuUWPBt1yycACrtUXqkN8phHVeIluZX+kjGCkYf9624Hy4qPlPSuJ47D
Rgn76tPNNrOMGRupe3k1BXqNGMYU6pviN+HU31spgYCjguj7cx7uH2MNTqcHG1aU3Mz/+kYOLlm5
+c0EZ8acOBNJkFoO3D6yHr5AYbu8U4RbdaxySeCo2LaKgzpSSSmzFL4d3WfSKUknTH692sjlQH+S
ubxWBz1XHuywJFO4nEnCEpdd1GpNUiO/e7L3Rxycu1NZa5MUZHx0Of0iFVfRhXgsUQEj8D7lI0A4
vP1oUyS7LfiTyPB2gK7UnR+lyd2o1lrlVStsz1UeecEq5weovQfFhx3vNnBXEQKayvvB6+qgUPxx
FGKbCWTWQB2QjlxMoffCsmHcM4hANH1OjQNYN72TadGwoEknULXB+6YVgx2wwIIpk5P6QX2EU81H
R0B74IhPATtHVVxY4dXxF8GBrE8y8PK0Usw4YRXUb8pLRTnwwQbWet6xBTPjNfOq4nx/gJfOS+xb
e77DenTH673O+ovGA8PjuQpmmLPjye+yP3ejlLMyIPO5Znb8J4t33Q5EnYGaNOAa9hfeRUfdhJCG
kkGBy1ppxE0rvYvw7Hgl+UFWCf14swpgjALKhwk1fWtBiu5mW2a3Z4QCrKfxl7KKQ9qlxu+w9mxM
Kf3NN55yKT6Kii1Pio9rb9hXflirsTvwlcrWCTJnL4lwfFzdhK4NMttckAOX2esfsJPZdz00jI4V
pyi6W4WtsRnPq453ot6eBeutDTOhn9tvje4PWYXkuEfxFbYdM60LslXlajIT8f5F0vdBob373GI+
gUz9o6HaWK9/LUGLGKLfTLMTH84h09+UJBtQ42Oknj6Sw0dQ8qQE0cHVA8nO8WBhuPaTvHfNxDG9
5Zoc9CC6Dv6mhYBQrK/CKaOVrq6Flx7I26N+KnPtxI5RpXYt92qxiBcdc2lpf7SIb+h/VRHod2Cy
AQr/eVU13ecIveM4Cu3uFGAJuKMxE9GYhDYbY0XhSiF6SJ4rP+KI/BBrrRGIRMjG9/jTrLR/caq3
faKWgr6YCyMyQ27xSjt/+SpQrJDyObiSEnrtT2fMPJjU1EhAnEeieHF8ME25C7/CUrX1rL/azlUS
3irWwaus9lIhmERzeAR4pmTXlNl2awuHqYyIuTj5OrATAoKCPPX3jtN2JzoDBkjVb24ZhQIuxooh
0AzLMHA3l3pPo0Kopszf4f2lfVKvLE5Mp4cEQvlOoi0vSw1ekYiExH95rG3X1UVS/AUju9I5BYKn
n1ngeeTrBebV9A1bZTw6GW0AbKceUBX4D+/OUAOSzDMCyEK9+0AyX8x51nh6vsY70SItkJTd0utu
CjeIOl2ybBsL7ZtQoTdBNClxkkAOEw3TDl+yKfvrDC42hc2RwXcolO1nquKuOEvXX5qdAPihYWSH
mDLa+TAqxW5elfrLWOdSFj1Xeee1Pvl7SQcctK4ZvXBzBlyproWUGV3KY1+9Q3Spntu3wKEb+YQy
+A/99bnqm43QFh6wqfnOXLiCRFvhMXWOD3IZb2jIGT2qAtTLT7zS2ejQO3c3n/JrQT7Xq1eR7Gp+
JN2bhcWtlTJ3IA8AGe9p0FwU+BIxoDLXOJ6LR338RIPS16ccTRaRUwUljkDG8JqwTPzZmuaTrlGX
jXVnci7Zs+Oo5qYhKJETciBmEzfVr6xyUJpgTXiIEKrdEJnQoJpsBBVLQ/brL8BpGHkKcDveFAmP
YnSqlvZZYzxNz+26PIWPufIsbMCDcFV/AaYGfqXiEpkFYUEn28EK+oDgj6Y3J839hUh1bAMs+byH
wrH93/WuWfUVPZ1YWv8FVNAQEUVCtl2505GTfbtWSl9QZWn/LIKtmBlgOK2i2tvBoyrOTFi9gYek
1zOBLxxB0ofBWOFdAsLY2vrDErrImfMDMNOgrtngkWRxZbOKn1S5t87pszVN9iEH9IZ8s/NM0S90
Urtz1W5cS8uqU8BF50C+BMXk6OBAm2e54C1/FQ0lrUJTEIDSk+2XA5CvHaHkzcBK89tGsEKQnPSs
+RCatcKQSMtwKHfGwrUOCAK6vhcCjPU6kzrkqtG8Oa5Y28/gjWfAwhs+i2hvGZAVio7LlyeEiMb2
eCmnP+7ajpiOnWWuHGX77rdnZv+u9yuyahQ6vMJAUuzJC0VURXB96LhvDh718VVXgCom6SdVcs1+
bh9KoysSuzgaXxYpnRfCSHcnKP6VXWnJWYm4wUq+Sjk2+nChoqD2BuwjlvG+5IXNlvVSOoXIvnwU
ghP0nNAqQQBdMi5zuErbwM1R/lsxk+cEQs0L7gulX3yhIpYcsnXCpycuPUUTIFMxWqacC4DM9I1d
hrX/316gbzpnMGA0x1FZdCB1RDVquidQAmtNgWLmoDQ9h4fCWjW4UGGOfgJNjYKIRceuBNSxfa+2
rpkWS3noreffsnCAwNxcVC4r6S3PN+l8G73pB0rsVmsQ8RycwDzKHj0YkzmtAqA5r2GC9OjSQGtm
2WDoHgdxb3AAiZ5CXK7eJOpTBRrOT7UOhOz0wi+5rqaxM3YTOCb3NOBFpY98OqA8OoxS8l01lGLi
Fwew6HY5i83FH9QfDQg/wXH05gvjwHo6qruRpxSbIquNf1OGP5nB2eZguzogaqD/vnHSm4xYFpFI
vu6fPrEG7PGjCDtTkjJsM3kUAg8I09UkHOcK6pF4dM0McE4Y2h3lUo6qv0wBYCIJo6jJDuzKtYhr
RZAhiy3lb2Q7ZN1Oc9G1MBTuDCMmQgke/rwQEUV4WCrHpGU4n7GGdgQPxaPZyvPe7ETlTuGxoaPY
0EnNctiTL27t1pgzcPAHR1lvS9MmmxWw+HTPP4WWeYYnOh4EeCo2a6aOYR/yOv/8kgJjuLRQTUTc
oTF7AqMCpncaCQyNCwAf0qP1ub4llJTCm4j7egHFbaBP21WP0x3bp7WV99RH7EtnLbsUePXIlJTV
lYL0mwllllZqhxVTgN6dkbyAXUFReWO3nSfYm9V/gxfN6f1wpjjZvtwbToTJZXxG7qocfKrHVm31
ytnwML+BPhbN8VEdoHWM4yrpS+B/4yo5GpL+6VJoUdwhlzQSJV5rO3laBlvqsDl0qOYvNCfE/5Am
OWXIdkAWwWQ3tF/vVF3+5/DbUQc/W1rELrZcSF9b8bGfwH05x1zquqZtykS16iEpFmaLoMyYXkdM
oRU749qywjK0oep5UGnJGwdmtpTcLeYHoGzExC5fDxrCLX7TOsGFqfdLOvJ2mBOATeZE5vi6vWIq
9H1+yY/j8EYsPEkcvDSHqTGiubMUphgkKupQOMI9oJcT4Deu885wS9GY/esrpXjf4tuVGRaaZDgF
0LfP/1AY/9lroiHm2gviSLZCgZv06JhRvVsbFcsv/eA7DYOP3hdWnNYv0gNunCTSB/nKth0kzhQH
2gVeujyXo++DBQYrPIlLSirXpC1TzHoDKtzR7QT/i5Njeyhg86MFNtZydrenJigi3cXRsYzV6qCM
EO9LSdTzq51EMi+9rC7irEGUmvdHxewd7yR63RDKBs55AVRXxloLuiYyQFurXeZZ/E97UlkMfKjJ
hgvLOv6ebnJkyFIAqAtpw7bcaMdkqpQUqki790b/Fb6bumBhEU6vEoDXnFov7vi6xlf0ZJYrLE2l
jldMN0nowhoJX65nIseCDSd67RVncMee4YlU1OgLnz9ePX0h48hiNedb1RnZ7aKZK752b+2KpDgE
Tou/nI7z6+CuRWZBYnOu3pbO+h3hWPHTaU9Rpf6vzm7uqCB0AQmYgrZoHnwfX52Kvzek+spFg7Cm
FRJ+I78xmDvwWHy/+dIuGkaKTwu1ENE9mCW6JSSH+3wM/OAukA85rVxrJtszybeyOsl7Ui/OMIXW
7/Ell6AirTl8Gd9w3cMs31h23tAzqeMCXjq7kJ/9h37Ilf0iRXYZN/xoZexA4MB1R1t9J56AnCUI
PtZij/KJmCyEU1tPERgFuLHAlDJWTl2hbetspPlsux6HOS1IjddDbsHUGlgxtZg/sO491vagg+uN
NFnx7Mqe5BAsshXEiMgg6GeLx+LFjRAm3oSwl3aWZtK7GYqqsr3kVLZNBRsaiAddZ3ZHDSfhU6TM
L+RM3g2/U9ja1WAuall9qDIS8R4RYNG/GK3tGHnfA1m1hCw4deQdan9K0nYDYpAr73mF8THXEPni
xWreLZplDr0LtwcBySJwk5FzyB0yEv55KkGUTq0A+/l09IGh+9402EuxdUmZ/CykgKvNFv/SePVf
f4r1Q33wyDJJLPzVaAHHPOTo9E9NBK0NRgw5T5DjR8BA0O2LM8iULPEaUKboEzHK4GismNpHeMai
cKDPC0J54/8NnZ0H6qlQ4EDmEMSrwb+wXAvUAsL9mAhuscB7EkHtUaN0Lemfrse6cikeY7ADTgUN
LYyH/JrfWQqV/G3JGbIlK6OyskLt/ckEfwI2gYlAZFaB8ET1h3hRq9NbqVduLG82A/9l8QZjv9m/
WGDjQdLaq4BVL+riLHAM0/TSs6qYBgrCXpI1oX+Gmb6meEYXuL/f+xHjRsQcVI3sFUMUfnpmB/a1
n+oGfd6ClENqSoaKHlsqy/r2CiOmGhpOkW9TtRVbk7jNp5ht4wb9V2q4UNlbbbNXv+G68YsqejVI
kqoE4pxAQvrSxJp554pn3L1cHuodayVqdTG6xD9ppB7lVnhfgLwSHs1k0dBQqkqiCON2d7FySz6i
ZxMEzwpMDgbSlkW3Q0efSbxdJ9ZCj0bBaz1boDj2bvfw816JJ0ibBrcAdMw2YEmo8cSpVJRX6hTd
EkFUamgRs0plPK4wcGFnTbtQXoLov6ONbofRqXEyYwhnrd+ViglorlVr0v875XOxPl/6xmOvdYnq
JPoYrfSCiXTZp8kCzegrDDtgAQZXPWHg258kT/hF37ObuIvLwyYnTF3wNyVAk4V28rnrQQvqVD9p
fa6XG8CCVlsF+72KZqz0+K0ESt+N8rQuol7MNjB9dP6XpOjkQIFheEw2XB9LJf5md7Odnre+9uCv
vIVOPDkD7xzEhR5tol6WcA9kaspPXoqsMuocgKE40zs5BqzO3fqtRxCz1TS4SBJWF01UktcZiaZW
DH3vgcF0kdwu4awWMCMxTU1ofjPboT2iYXKV5JP+vs4y+TCDW7KtahOU35hpKDoySj78oJZr4AlE
kBnDmDHu3ISanK8K3bCkmWI3qoSQb6K2UkELbj877uzmlUvYjPXBkWq83Dfrr/2yVDO9NjNos8lw
XNh338p3w/Ta9tgI6d6pgR3aFBVPgjiZfcr2St8aEcmXA06Mh1Y1Tum/sPffu5W1+f4Wzqe+oxuq
+YG9Bx4IOPeTYVPDq02aneVCUkctp0l1trkUYiLclmT4DHG9nuyI6crh+jLYCn2wHWyNYjmITLdb
cguDz6zH1dJR2QjAwNf8X74UN0HvketcghVl138QJSOBHP9808uX7b3OZJO2Vv3OWtQWbBTJxWBJ
SR5V5leDEPUUg0/ih4GyOPXzYGz6xA8q+t6bWD1keGD0vnQUQOJOH524XZKXR/895veJbGHv7+9P
PnQzXfiSd2Tvww7rW8PWVYXWOweXeqMBxhGaMUAJ6ZlP7MES3qply04rAXAydzO/KB+LJ7jhgAaI
eiJYFe7fiOd6cPzTU26lecOfo6/ByiBc2hBrPVPst80bw0WSwPZyhMzSWYvLmq1YW8EeF08dAqFJ
Rt7VmWQRFO3BJcCio4+hvuInIfWc6N4dX/PmduZJOX2kubj2HLkuEBvr/WpEMzuiO7uRg7RRw/cH
EX/3j/y4qYo+7KIplFDh0ykkWUsU53aq3Q1pGbXAgsofw54WtXLZeps9WeeFn6ev9OFQCL7VC6iR
aw225+PraFcY9uLWa6NrGJbFFlzlL7JCTcJAl1h4lk+Aop9c3jaLGuJYUAEfqlyMfi+lp8fXWVKj
jdGlNvnzAAhzUBndR0ZGAN1PSLMEe5OvAhsL97S1Obx+GFAZZFViUme/r1CshH4cFPUT4coppTBx
Th4ZMd5jrfZEkmbxhxOwRQUcY0TH+aRTXAok4FD/diSsZZ5e+a2jpjhYBS+FPWV1kyR31Jd7e/cb
3GOsDyY+vk/slEhRE7QcGQK0sQ0TMfmL7MDSbLkVmFtFIB8ooQg+HMCoEy+hT85iE2sW0J2oKACB
hA9RwBB92WHA5JixG1AAf3uO0B1FjQp86Nn2+FWHdi6Da/LBYYpnOIRJ/gMNZeiKEWChkAiXOJuE
h4r8Oq8vVyFUimdbrZYIOUpbC3DabMWxvEIwPpNtCCug0DypjoYLT5H9CHjOhxIsrqryYRtt6C6z
8Svb0NRU25iLp7pVlEyxxtIXgF66oYfZpoDp67rPKAQ0iwvZKm2GWqcVO3VIaPX3o+gcW8g9IcAM
gmqapUeSvt4lyn865NE/juml0A+It9lVuvD+6iaoeuPCOdYRx4lpq9i3H2kqdhp+puudQ2cgRt4k
9gOfQ9svO6+9cIJwsXyN/e4Ovfj7XlNP61nQXuoQdRyKQajqB/NMt+1PYhpcxYNKL5CXkexsXdlw
WxwEEPa0o0Ddn6aBIHXiTbk/8VhMnNY0aNunwpXyOAiJlPMn41ontGmHKSFLQZjx3719gIfu8qTe
ZB3xOHLLhMFGaY/FIXO6EjuEE/PIKgmQcPxspvapkL6xKtVbNZ5nllJ72/cqQlqQfjBq3aN3aMaR
lSlOrA2xkJou2D68Iy9Bl7dywoqacqpCklEh2EBrsd4rR/Yvf2la3Q50+7d/0NFt7OsVUCftC5+P
6zXTRbyd8H2LTtvuvkJPoBowPrBI1gphAviCwZ4BDnl7NggoVBtfvqverN8u8I9YYjBtLCxnFYmq
l9p4bXeyknrfCZjEqvwNrEHgwQ6xuuKIl9PaVTCrgO0HeHUiKVpkq87+7LJbCVOPM15AG5hjgKmq
/AOs7H7GHlUGudp1K51B68pjqW9aLoHskvkfl0zfefRVIl/JBqnUFZhqgfkIB5veg4KvFEnSQrJy
m0k+hwliMn8IxejvFapUt4Dp/IqvCARufQHU4yzR0ofHLl7hQq4FrardfrvhOB35DKHQwGJF4r9O
Z4cdVbbBCadLL5K65/SFwxK0rnVtAHj9ZBAcDCqkOuw0fc31nysvcCDVaJ3SawXjc+MSs68JWJwI
QbaC0o09vFuFePGq4+aydUC9T8UoR04aow5i0N7qrAtynUIwxsxcfK1S2+kyYYAleoEtS5V/LFcI
FKmG6t39z2C5d89ijcE5Pt2Qczh5SBRkY+0jFkNaEewUrwBkLI0sIKAm4iX8TI47XMFrW0LGLueN
+CNZ6oxrU7SZoUDO1jKNAV1E+i8jKEbV1gcFhXGjxO/tRA7CbR+sxo+YumgvYyBgI78JZLsKwy1A
gasjxLA02o2rM7ecz6RsG4aote6Vxs+L9vgVFrE1unJO4CKl0Xua1I2lSypmZN2JlekWnTpZ+EDq
3rAFitUToIlmT4uTs64Id/tiMMYR9LHnPEX/Zjq6o01s1CcpjuKHZcLWQsWYvO9iGRB0RSC151up
MLdZnoDlq/gEQhzG2uTS0BmL7XQeS4RuVDWMZrot5qXlacAeuK5jcr+1Rq679ib5IfB2f63RbDyZ
nsONVfu9Qc0dNnenTcmApj4GQwS0Njw+hr6FQU93xxwH+b3usCSQL3qtPMrK2Bg7kwH7SfXHIzoP
ZDPaPcayTj1uiDrsENbNlBkWFjuk6H8RC4/IS2kgPT2V/k1xWrrLOOcVITBvy1tKK8QkikmR9s2k
06Qid2HaIifXra+1isap9sDMpwkBnETRYV2qM6Q5D5x7rngpqQLKTLIcvAwRZNqW6c8OQl3XXMQY
8EgLq7ar08Qr7PtwR62CguK90iifEpDdLrNtJuSAsH4fjFoo3WDhYgqTHVOdxWIdyAHy7ylECy+f
ig9LI7GNsV83UuqGl9y54qPPT8+YVyL3qkwODNMl0ibx9yicgWv5AsyeYoUAJYryv9E20Qy/7rhx
hJL9XY1Sc9/2mjTUY/eT5Srotf+YRR2hLtHKcBr6LQ1esoxkr3jLpw77heV+O5h9guNbW18x9Xfh
oUqnsqWLb3SAILIVFPO0HaHi+7W+86TSWP7HGvGGvqWRCAPO3cxQz8vkqguDFhfFX1M0bLQTYU42
yDCRppH+KxOoYaMcYF3dANurqjE3BvYBEJbc1OAu9gVgpq7URMAD38LwvGqtfrTiYtlv9zSfmy+3
Btf+IwoJHG2tieS5ckETPqj2ERkjP0naEkchq9ne9/h6FeIhC/JyXByp9kso9qcU9v2fluCayeIa
vQKzG9piMjr/58RXh28cdEv+pHE+tSTSXt8FSrugSAeKM07ra6tazLPr0c6NcXBl4IlLnQvGuRCg
ZPGG/LgmUF64WaOcnHu28H1TwB4VZ/v+pgg38MkAnGIsi4I//c4d0zIXbjjhE+YiEfrJh4/dp0O1
lVfgdVL3JNQaZMGq7EdvyKi+6SX/VMt4YI0kIOCgz+16ljBN152LIl1AJTkYdiDEs3lhXokpbYqT
N9snDGU1ETXlPMrSDXS3pD/tnYotrJI3cQ3sGDHd6fjKZwaVHQ5UiWVqKPKlBK3SOfZSHbc8kNMx
18HY4hWVEr+h3UjLB5cxLo5Ux7JRRIfOgg+B3uJY0CkBWbGgyfrsK5sEVERA0QvkSXhfLEtMkEBy
y3X1AVQUbmIrsQll2eRA4akUSWhpZCQOnT22ESRIMwmwIu9aq6D6RGwDYuxFx8VVUa2qTcBuqvQz
UIrVrzs+EG667ZimO8oobNkNm69takpU098x+d8yAs//4vOrj5AsW0KdG5Tu3bD7pBX9iAlzlyqt
Y23UCkgS+ZsQ9CLLYdRKTv552HfeRKGe/WKvmOsWX4Q+Xs9FZZO6l98f7WYlPX/LS6A5sInzbLh8
Ulwrf0BifDoMiWKPDS3d3tz+Qk//XsUdmHn55QVIclS4ZLbv4McewJLouvMw/g02xo752Yw/3OY/
pM7Tzb2goelh04Dwa0Ye6U5otDS+xCZ8d3DFalMahZsramlmOjrQY/2G3Jzsj0qHftGhum3aRDBF
ezV+fPu4FIsuGHffzn1e7QUmgj2UTMROWRdTFPBaeHtnCcjON88ou+NEc5ZrDLhe8QdvDwXTC7lA
iGyCmAsbhJyyi1MiMJLTXhtgP3kYrr7y6h3Ytu2nCAZbRmRgWlZQ0KGknfk5by1nNbAybFVnZ+A/
c2y09d4rTMeSmM1iuAinwDSEmPSbsjUCuVWNMtl3LSUVwQSFRp4JzcWxtSuv0NrBFGriwJQSKJQN
+K0F7Tb9pxg42rGIFkpcZ2tXfMshbGWQ5AES0RobdNKpt548hTcVYNl7b8YI5Mqixs35fCXfUUOr
3VleST7YHwdfxDCkYUKPxqwbNQDYVTuU78m0Gy7aXJRaoohMfhMDwy9MSyUzkmBz0itwfH4asOAH
irJQ0f7iBAR0DXhzt9yr3HlZw6l2JB1TXX0rYRKZwlce76dntE4I8VG1Rra51yObfVgWtd/HfBeU
vDiQMOFRdATL9q/HUL9wh29vUzvFyNd6HhXhydLRr5BpzLx0MCqh2wXVtoOiC7ApYjcr7jgd+JJZ
sLYdL0Uws7cARUnzo4aYsGWmNt8lxemswlGW6Q+bdSaERGWWMe8scaJdsYk5fe7m4JE0s51KsDLN
3CmkZH8XQNKYeG6FduIGbbKXJBktijmGTYeXHvPRzVecueiufO7rmSQ5Ft1Sb5/F+x8PwjFMp1Xl
mXc70nj7ansnhNumkm86u43OwBur+ZEw5jKvKxDiEfTyOMIfCfcKHCKgLDYBfgrrlRpYbjSE/W/p
hlYAW1y6pVJfMdXOxzrRjHq5IQ2EQU7/TtlNVShfLDQ1GXoA9/KKZTlGA5ewKLfuoEaJDzq00aF8
3QZxYlUwMjjPqPlJpAyltEUjW2YEZExgt9lvdERteW9iFQSfqfiWBE6eEApgrTFLhSIbdbD+gOpF
QMILVxbaQQbmykJEfhtMo8afrcAzLFpFZsEc443y5PikXE8q5tLEfFBQJknLXalGbpfLTusgUkwx
PsuQSPYtC6leAzKjCGJ/+97GR5HYiV1X/D0TjDG98khZKgd3eFKF2GKc+Y4mE0s7ksrAfOdWAo0p
GQu1BlySKDLKxWvlH2+Nv8dljkuA1U2KFLkw0bQkPNQ+EIeKWcWiYpfbdlsQWJoH98EaCsDKvZIb
HjdUvoxRLuHByEi6liY3EGBpeXltjtrwcbWgQfB09gS/c0CT1WBVahhoifJ9+mUJdLtxwbvg+Vjr
Dr3YN9g2FOkcfCmpPmFUBQXEhhjeHBaU5YWfkKu5PjkyZ9in8yNrzVDjGiPmovt0n+hWPfwE+cxW
iLXINnyWIftcauG7UyBODvp5gABTNQSfH3g72YaBfmPvZjcgO/pEe9jp7dcHfleEVF208ffPPBdr
umSUFiEoTL/mtv09U++37/Hv4cEP0ab+0qITus0yFMnCzooGD9iQtDWGrEaRchlJ1Ohb01GQ3iu5
hwPIrwCgEtaYahjXEuURvtoDGywfD8Jbn2SJxyX1aoaEI9DrreBsLj94/Jf09o10S0wo/yywEs+0
kIcmWFWJEK1Jn6nwFM7WSqlF1rBBKBClegyxzk42VG3lWjNxFD2rvFIXC/qZyA/jTYdhq7mWsRSA
Z8nt4uJupUVEpLUk1Zzl0uLGLsI8fFAiav5k08M2X8juOkAgze7WaqdKBiCUKiEDCesZOWj2jryi
WRQacbXgpXhqfu/1g3/0c056bghcVrwPaj2RDv86l56G/7xrTJT7HuU2ISkf2sJHqSEHZjjfjocy
fsuMzXBP6JRsvxK1FUWieqrfZ01fuA/KFTfCIvgSJNBtCWk0lZVoDzIILyGQVMFRE7xm0gf+5pC/
NdZyey3xj1hmozgQy1AKrIxsPKkQy4+TDVSTiMUBm0Z5NjfnDj75e/cfQibP1gzrFt/M8s9/i/Ch
uLGzws8yLw46oowuvLcU9mHqqOKQblhbSFDMTNazDOP3l7AOqN2uWLM09FpHBscFiHL8PiLxJurA
XYtszEjayo30RCHwXv/9GN2q0Bms4zceZD0lEN8R/IH6fsm7hhE90VqozYOApvkemOsGQ/dhi7Nc
lViIEI+G5fIZmixtsLwnUOFH2oSzJ9DWZ6hzlRMWYglTGw5hrEDOWKVbs2Dbsd8LnBKWZmJOFe3z
s1m94tA8uV3Wg62cv4OD4jGTBH/mj6T2j/weWTpsqopLM8JiYQy/8aUfizcesllo3XjJNEJ4en3J
+DPqD7gsxpXFNbeTs/8aMi8juiIQP5sQlnDmgPMiCJzFuk1KHw6MQZw5XTQ/jc52vBYvW7SbWVbc
4wjiOy5uJoRC6JM5gaDO5MBHAm5OfIW6+coGy9KTPbvofT1Ugk8M1AtzSJ9T2V0Zy1CCc8b3Ns5K
ekNw/1HpD2y8XKNdWh3YlqlAkzrpAAEn8kK8idiXTcsI6qI8hKrX8ch333xkpGdkTVufGjaDHoKg
QtI089oA5eakzQAkItIe/Ba5UT9yBKp7/3C6QdUJvf4oBa3BGs2jh+Nmc39b9KcmOA0436Dx52fm
cLMUQPb60OqCR5T4nNcZX2xnyeVJVYq7gD8S1XZnz7pKcQsNqd1/b4Qh3gIt5zUuqplCV+xzAcPX
ltc9KPDtNGFxcUxpzrRbG3clLrY+HA0Z0o5M2+d6SwqKWUkltw6sULGQqo49scUA4BEe++rTGjXP
THvI56vW8qAbO3YtK3QGPNDNWVw19FXvTjGDVoLczkoQdv/TKr4pWO41zSB5nVPR7Dkovl1gBbCD
OCIwfvpO8kCt87T83ILnUvn8jAe7MFSWsYqjsZ6c83ucopztj9+NCYg7XwXVt5EtzQ81a8oyzBY6
m6/30tB6t3lvBkNSQQkQIcGUhBsOP8M/Ksk+CIbr0Sgix2/kISQ8vFWJBBLuo8KLWFiKZ2m73O3w
3jTgvri+sk7GdbN+HEQ06cIggzlEjfZaxw68E6r7wIB2AvSEp6GTX0hQwv2dpAzBC5HZKBctLFdS
6xyEkku9slRdSH6UM/SdX09thOr2wCASuiGCcGFPW3i1InZ2fetc5E6PNW0bEihEw1CDsKLkIwMw
TZp82P/z56UpagSBJiWyiMc8TieZtWTvGkr6Ls423OgBEtpg1zl4coy5IYJRa3jflH3X2ffReHVR
ADGWKpRxWeTiV1lFrzSzr8jDf34fR2fWM0LL9LcgBPWxhq7Bg1kXgl7yNxG6ovliE5zqjQ0EgBrK
wSwAGtCq3wunUzBFipu5Vlhr9yaoyRPUNTZ82QFm0V3azHOQatl2pwMKejKpgU9iwc1TPjvplRWB
hy0WMZYhfkcjsoW75dALdRb+mV2D8KSSK+qZpcxw6u0wQ9jiivt+8OwBjeEnllGVVmr/kwg1d162
MR1+OYtoe9anBIKEagn4Qt/ebHyhfVCjgzdl/M0f96n27hBv2EGGXuveCx38jGPLcp9WNuUM0QTq
JXuLIKKS0zCYRKbr6QA6hLxC2JQraeyawC2pRzr9/wiaG18v+7WKw4oK/oeq9Xhc8QgxALmghgli
z1QsrHae3OJK8ZObGUqfK5EyO47j77cGwG7QuHAL2qLGQRvDwLvzmQGewp0fYgC9hjHJndADP2nD
QP5HOa9PoiZ1+hkwVDqgASuibcByzKroO1AxJvVOHqQk+jmFGAV7JopjYJzWHdbo0Ys9wmF0UYiw
QvVhCUWSq3QpEjRgS2EL71aH4q2mq3Fk00qoCJYDe6LMZPHNkHKCkJHb5LmUiTFrh+8IJ7zhreid
XVZc4/5esGdlPwmkoBzzvjGXb5sw5pC+di9r08TEpFknEGGCZsWrNF9H4vot//xG7dI7KF+wf4q+
s4tW6AH4zkQOQUJj1nzkRYw+fuT3JlPm8w9dggU9EIHr5mkUddWLcIG/rrQxYpum+HidGMfehYQ9
I0VmfF8QVvPxDfJ5GSfWVlUMy4NCFZrcNLxzS2LEuqHo/5tQR9YVBIekW5VUtvvPGfZoIvYcxn5v
mGno3jQdFeIqjH7aQFYcR+eIucOujpHQonGG9qpBGYQQwRE5q46nituQlq7qLYGmgO/CV9YLp4cW
VMfLzpwW9/hf+WOSKQtqAoKVFO930xk+rnZyA6vD5BIFyqOrRD0bN/+oKJsFwUsusqx+JrNibEiV
Cex2MTWUWENddR6thBO4CgmbAhXsSU3SLNUzujUT2qt2ORRPM4TSlpfrtDveDxXxZB3SzrPZGZPr
zh5qfBbv4+f30l6dTWrBFWtL5G3VvPv/6Rz8hCVYc6ZBOSoRwnW0s+BP/vMXI8hQP7lSCDCIALX5
wZG/VslugojHa+aoSYlTIgTDSAL+WQ2VZTST+t3Fhr9HDL5VEeyD03h9jks47wq6gPfhpe9PXswC
Vv4DeIg+KsJv3LU3ZJ3C9QpJ1XsWRlb1agPDls3vlj8Kg30OdgxfFrAZY1CBol5RK/NmzFtRl2xt
sWWQod1nrRhX6X/JMq9scodcAJpKYDtKZnFjKxZGLKbALGV/6a2IaJJYNkumOH61rignHm0vlh1G
GrEgjSNRQLxdFC1IyPUs6ktD8TghO64euZCK8Mu1BfNkS/0IzIpPz70FB9zcOd2agtuwtUAxcbmI
hhxemoBBsIb6oKw0J0zI5FgQVVQot7MOticyURZsxDomfvZWqovD0nw6H3cxyPz5ATJ2okzUMNyW
KbUcm7Yt1q8o/t2o/H9iDJB5GZS3yYDDkiQLbZLWbTrJnG6icBcyig05w0juc7u7bZ5tu4COwytp
BnN+w1AG+Gtffuupv4P92tI0F+iKyxbG3WxPUVNali8AmJyjzWVcnV22OkoJRBbdnaOFqWeG3UEm
PW6lk7vYBksUAvYBaOlLF5bbhaRbBMUdOOt+GHkz1Ubvcfhffa7nPhgWhXV5++VY6Z9RiTDHyKHN
FjRjprYc7MET1voQJkzGxLmtcBWlniciZZTB+tCWFxD2E9MqKxL4FCQrFhyI0A98jBbpM462yIya
/h5bQjR9EhXUizXMEEM8fOsoy0sjRWAMzTpEa9KIwyQSus4Y+HZs047qtp/qdB6FrLGzLoti9Czp
6n0dvDFA5DpDkzrCo+IXXckY6W9dSW3kfdGIUj+c77piYl6Kre+R6XNzb4p9Xy7wsPaMRzLh/YKc
lDpxoR6eP9aWqdpXCZA/CycCY8YbBrrbbSXE1DJBupW3yemuSvEvPkqGxncSoNzQI9ckM4uxOV3w
unf1iWjnJWVIe/iqsJbzFfgabUC7jcfXXIxRGUzBlkAKQYRkui3kmvstgWkh8VMpz0/KAlu4dibX
b3CIcYRQpu5y7Fs5h5jh3xuS1/gsnSORVxqZUtrgG6/Wx6xAtuuoz4ZA7C//BiNjIPGML9ABdtzG
pWC85jb2YL740CYgOeQ54zA1DyvrUSfHdu2E5fSU/by8TRsNhc/coAnWeyLehDCPCeVXJ3Bm1sJF
4rGle+z1FzyPun2e4dQMdiMaacYsKGYaoEHBnp71wLFZ5F9TpYfcNREJ+0kOaVvp5Px8BVVt0K2m
AkCWZ2Wozsh8hcPa06Gh6VRsrSxwBz9ukXXnb11BCSO0n0hwt/N05ZajukOwMpXzrMP5BrSDq8Bo
HCr32kpQPfpw4awe9xCtBv89kGm1q/ohyI9EFZl6Jbdf+MBk7SIM/d4zn6pudr86JuvTKjfLm2hG
BcT7OLlpv0dIcoK2qYE8v30vw+L6csmZLZULcF/5azb2ohBzmBLPr0caNXSPy5ZYUyLzP8lDHkLC
biunTkVKuJ4n6QIvxNqxEVYE6jBziXbZdmT17rRJkAfQwk2KyWKiFKHH+8y7uOid4q8rG7Jd8YPl
u6Kc68Inos4KlsYmCWuMx7UpuffZbZFqTMt4v5YFiwKXZ3huY3NpRKMxCxb76V/i6Dm7H1tS6+/+
ScuxtXXJ1ulMeuiU9WEWfLsvr5AzXhh5Ib+tnxvux51JLRIjSGCqfi8th0zzLmxvXidjiMub19Z0
a5WV0FAm5Qyb7s+P7NNFWvhKczUOqAE6p+jk/OnFVuohvLdM0B7sD5B7pTpWRotenlNq1kxSPEuo
tp7P9HtqTGFgdHbH1FI+xJSGz8fJ74FDutr77dnoCvjL3WwJyZwlRViPBuElC3zqWX8OMGTfwcKq
ftnPmsK7/vODaK1WctDGesI/S7lMVanTK/XTxxTD1uE6umeMWwu9Lmf0GuTfZiK8zauCXzZ9F+co
0ZBdDySTbdoMnlyzLlXUpsDniT3DgC6te5u0LZtDEnIOlsRW+v6pjAYeQwf2kyoxHKCc7mQo89/9
KYZ/Ope553YarPx7eqoWt5O+c72+FXW6i7gyvx3QBAW5M4Z5N/asLJFRyY4BnsBipfiJM8hgxD6O
VLte7mKnRQgW4GwNr1rJburb6Z49ob/vhPZIa1ytctepDFDRMZLyrL4UsASjZtqLW944Hndc49Q6
ykJ/02vHAkMEfgvCu+ZpgHo0jEYMQ9R6jtDuEeuXInMJrrdIAeygNb6/Wv4t0qphKyxMSjFBAmMp
DYALjiey58+EW8DLAmMLnDX60Zx/4zfxWn0Lk0ll5qxNMIcKp7G8UEyArrXrRCdW4hHQMZNTMprH
AXX9bxadPFVI9RRXEHrwzTdQnGrTuHEi6HijWPbceSi0WWZJR0jWo2ipiWPv90HVxFTDy/CMZTVz
D200IMDGmueI8nD5JrRICsFdmCmJKFABKp9eQrNVnXPi73Euw33H6317SmaKfE8S+19V9HKHeDSi
d8wlNeS23/N+5GXqx53NE4QT4BmYz6ueSg9c0CvFq4SeJdvPInss6kMdSy6TGVWH4YnsfJjc4153
M39Znux44mIIABtupCbqQGStKSRMjNxl79vjx7XYza0yfLubVIT/4/9VnqLNwA8bUlEPG1h73NAB
fjMfzUevKwIIvS0f6BqVuk1j3v+QZAOO3DcyFtl8lvvJJWj2W88pn/PknkJAwaenAhfn+y63Wvfs
gZC514IVjok7Ak3rRq2brV4uEKVllOas6MSXuYSSNU4XGzLga4FFGZ8/R7053LS0HsGQXiBnseJG
99wsFjBkb3kYyQy/yfUwgW/rc61lWEH+ZWFG2pglf9qX79h0kmDbNkgZBYCktc6LYnE6u4zSYoMc
ZTJV9cI0Tx42hYNUkzRmIKS6J/Xw+CEOt0pW9qOCg67XURxy5f2iLSbpPOmdJjpRu2FDrPiP2rMO
QlP4OHk6FrPaKT5Ojv8qxF4cqfUCDq9qc6HjqVFCxZQkoMPkbqOkw7eg8JK9tUrYRktNJOJ5f7S/
Fg0lTRqSaMzR7VtnkCXcNgdhRIpm01QSa9FqhLtEHwmAUeX42OQmNbSn0OCGu8O7AcUnpECJVfEA
u6YjG8Hdpky9DPc+T7PMQ3Hkby5u6DxT9OuTPoQuDBbPhrjyJXHBa1nKHX2uFCsJ6E7MFxXsV6EN
898oXT1yW76wLjCzyp1as06NuFAOpKZ02+ClZ+OZRNYZOIk4gox1dpiA3lDsfcNn714KaWw8UaHL
46VNF7lS8D8gXhwUEk5pqtYpiNbM1m3LPWz6VIIgV2cEGIzWWagrABG4nuEonJYoPNR3zyCSQeU/
zyrnhjeFGBdlnYo2MoE/14vKZC2sjyFM+iqx6OYSP/irnxqJ12XhFmzDaGuEg9Nlt3rqIRMTlG1E
JJSHIJZnAW+onj6UuuVheTthqRG/k6y3bvRYt/TtCTiiR1tNnOrSPy5kUkuICALS4u7rv9eJ4zUc
F4XVns7fBH+6KkOhY1mKqYC6Uq8fECupwOGXueyRvinEBD900Q7I7k43SY/LCHs7HR5lmckra8zp
5jzmyYJOJGqLCZjhxbi25jpXb+u6At9JohLZrnOwajeDgoalibE8mx77vYoNvXCH5efhNNM6RHN6
GChe4G5oOvLCOaeV/dVM03FELeeWAKmGYGlzaI3DeahSfr/iaaTCg7CW5RIRFqoo/bI2jBX6j1ni
7w3eQIX77IO6BRk+bTrhYB5UM6+9QVmA7EqgTMOIXwH1IxEqvRpy667v6RmynPPCobKd0y2pz2rk
wcmZupH2IZvham9qY9WjjKYn3RGglylXIV99fMULNTCpRuRn7WJ46LKqNs3EQrqQTKhIe7wQywl9
WxUEWK1s2NIso7GaSHnzsgbB79BDzRPFk0kztFcO5+tfrDyXoBe6ToBbBMDpGImtKQiByBp0ei3s
Eq6nnz1GXOA+bVSkNmf1kcA74PK5ZwsXqhbnk75BeJBRUF+nl6hO8Wo1w7kP9sUX4HSlC6xkxJjF
R1YRfrAHO85cnCXXF0diLsUONlUmPNIHehI/+S/YEi+WB7ynqnOmvuUNg5RGsXQsRobpktgjPFiS
6fSeo3sWK6iUDzgdLBhbnIbMwb9gV0HgWPLHC8aLY/cLhk9lqEKyqAbSIODX7q6Q1iS5hANlDcmw
/JPM8t6znmmFG1X8L2QVE5Aw5QlQNQkmM+y/SF2dGtkXDEvyZq+m7ZniAj9eJ7D5TEQRtgVyqoMA
X/HBFKAXgrdikQ8aV0a0bAZb9du/WQlRmqzOomWuzi40KkPfmN3jzTOWjolJ2ikNtwXLt/X7h0v5
yP0T+JysrtuTgTItJ8UYkON8Q4hK9YsBFqtKwxaY/snFztwlBb+J6cc9BnLp0BPuPpWXftcd1j6c
KCOnKrApL71fDlBkNkejKVgNnAbm8evFC0VnZ0KVBy9ywIOV/uKk1z7e6kC2vFqZPn4b6neQqFgY
X4dqVt9WbB3zmICaP0VSs3o8QAYyGack5pNXsGz9mMEveSILQMOIsoFnXr+rbRpz80QrtULfVdIT
ESSd+D0ZC48nfnfwF8ulT6BWJnBCvhZVP3eYg02MN/KoBG+FxPcb0o6LkhGg3sg3RPc0xIUYcP0C
+vo7WwRRlPKBC4/R8AAfUcFd8X0hG85KxVkajxMlpg+mZBDT7utXqu0v61CNCjdHWNIwyZL9BOIR
MLYzm13+TjA0s62aBsbqUe4tHRD7sN/XV1jSC+dvTAbMOmnCAq9kCjdABEyiS4kvL1PREdv/kEuc
VsIsD5I+PwZNF5ARpFe4N42FXzOJ/MtnzleVLvuZzyIIxxzDReknLQULnB2JBl8zhC7S9k+iJDH9
11G3vqM+Zhbl61X1XhIQ66cZrtq9GYGKObljmQ9nKT/Om8Ap3OHkonCYyGHZbfc+DbFk1/RSbq+s
7GgfS13u3zPBV6pHlF358XU+DTvu+sIG2Sl/AZf9cZfvDRLTQu3cPbvyBHrXx3Ftl2npPKjZPuic
EB13CKuv9MJ80Gh+x/xHUL5gc119j8pPGSxuPtaOvZc12mcNDb+Aj1gmbBeojiNQGlL+d+dOe8lY
LNEiVLGY4SRW++Gthl5JndSU2eiF2qdfc5emk7B2Y1CkCHHO05J5VPBhoayviUJ6aCdp7RAVWLPs
Pz3jOLMIKDS9exEMk/hwWRu28gf7xNGmGkkqzsRgyGxtNhwrFgDtzHQ4UPoqF8YQ7NmugVvEUiFz
DAF3v1c5Wo9K6Z9TgcQJTeqmYkOnJwEEi4bMHI7fzjkYHouwtJzNmBbmayaEcIwnIDvkbf15WF7c
Oa7eNskdQoOm5NhsmRFVrPKDZLsvJ28ekWT89/tu/Ax44Aau/ZonozNfCfx3ZoCnkQ6pHhyN4ZMk
bh359R5MSBKxtCiASXvnUquGgDJTMG37l8ROAnMXUtUTURvg3dGJZDaUFFXfxVu0EiNVg9HH6cxZ
j+L5ubIZ6i4osTuDk923iHJKqiVk8U0TfZshyE99MqDhPROuN2NX8aLFzqlA3wKrnnn7JugXxRlE
WYL7eKmhKtcPZYaGUAG8a7GC2e8sMZusNz50uTSemy4NxiqQ3DBrcGrDaEODHV/V6z0aQijaKVex
bAubchnfFIubCyonfIfoUK71tWCVGbHJePiWLS488SgHmlbKyv2GEcmPuU6N0JJidQ9CP2vuDOP7
w2vqSiwn8yGvPjSGqLzKstexsH9pHebtpqxnuCJVstYfzrrcJx/RIqeCz5JR4jPHvNSUZ74u0mP5
YxwNBo+tgMRj6h/9kufciJnvPl6t12FZgo2hDb0nkYDCArPba2cgZW3mk8yiCdCr5HOu6uuWVqta
MUukPkDGT55Z3ouLjgTgKtj+gyBYckTQRQpx8vQ8yYuMizhC8/QkahrhlTYKM1GvNMnutOoTCvZd
9mcydz01lZm7o0Ls1BmUYqF8nKbK4OT61PA642qZrLy+iDLO8JrZKcq5uBMvtGusOKqfBVe1mnww
os3feo+BfLWHAuEj3G2+zDjrSvypYUR/hBBY5ClpctUOZVNMZbly1P4KuqAYo6MZq+DBZ0bxQSsb
8H9vIXUsptOBq6ivL4XkZAK1OHrbOsn9E89lDtmys56WGnI2PGDjJ/v2AQqhQ2l2Ub5DNdNYXA8C
oCeoadkL8s6f1rYgm34OycrPowCtjJLkY/MHkF8WPxqlwANmZfwoAGo0FYszItpy9OIzHD2z6Uz7
2moQmms3tUudfYDi2HV74GBo2D5YaJYsZYx6RjLEVMzPH7n3gs38w1JUqEOA4BVg4cDRk0EXg5sL
GuilUyfsSWbaeviYEOcy1FCOJ3TiWPrzRntB6n9AI2cF/94JPAXPeUbO3XeX9DKEbwzxUkO2+mI8
9vDH1xdZzCmlNORbuDOUTFR6gcT/CNPaEaNu7A8rmc3vQlxFRex1M1WCGfa/FATAkafih2qhNvB5
IpbHB42/ESp0LNTB3HbJinZZjsmTVt5GMlYj3SzdRj2lGx2szgs2Af2s99mjwyvhEUqu8CgB1lvQ
xFlFyn97ZFfVLvHoxhgOcKNhWqP7T58W0pd9uwj+qA4V48xRWcOFokkNl7o/7lsGorL1KG3ip+aA
pKZJTxoXJjUNczwkIqMF+nvfhZkIqn6FyTzVybfZ4/B069UGssh76NY4eLEyAEFsBtZCeKT5bMta
USG7tz8RZi1SFKxUWsJD4K7hkk5Sl3Fxe3/O+rwv0twjcPc9HdNp3tdX9LjeYYIKQOA5rhAtjmyc
06J+7nwvQZN4JXTZChuLIzkOA3nwIlI7lfl2Kosc2l9nQLLx3E7UHrqXmw8MaJx1e53aToCwCI/K
8gKLaIDFh2HlnH/7cVeXJkYSP3jl6puGYOE9ZY5D+IhWc6y+b2mYHfI8r+lNV3NE1LU+xFLbCOVg
PyXXhVrbB8Eq4gKm1+mhf2xMg4CY/q1l7HfwCFafoYlchsUF0kYoSKrP1b3LXJoesKpXXZfhiaji
MXZVo6JnXca3uD9Zh13UFoOdZbev7mE1g6FQkZg/e9ABmPwfkSHVhFTFpT3xM2fnoCQh+7VvvYqc
P0FFyheogz/F5bFZqM8eTsuw1rjuWeyib2h4S6Irla64pmnl6HSpJFM+5JeABYf+XZgd6bXOB5Ik
Nsh4m0t5Pi9HRJagpsMKnQTeAhebLMAz1H2YN++nbGnQ2glXkjlbdfbWI81XyfOQi1i3OUcjHLpI
GZM4TfmZ77WcTjEAUXAw+pd/YiLh3C0yBnJxNeDcqbFLmUG8tcnrSjCSwzUkI8uPVP+rTJLf/3z6
xAN0PdWUhtjyQGNhxPz2H/iBRLrGKTqtWN7NwwnXWVo5fmiHm02PNGTfjGb7MDQRrp4MUtdqSHyG
QaISBB7WySlVZ8ZJLNKFnLKGMuJY3ZU9ASSQLoeU59VbsmKOLtmSgaQAJ/EJMEyp8WNgOBtO96hy
3DpwamLuofFiJVRnNmo2OgVasOYkzUyAR9QHw81l/I07gx4yGZhV8ZBBPmYVuchkiZUpHCLmGlBn
BqhP0GqsZe1x7h5hVFfThjXr3Cowqb1gBVE75eOpt0Vyc2zgEK8kr4D2GbucDqM+yXJtSC78LaKZ
jlYV7yOssQaAZCJHKGoFl9y7DAbnYPCtZbp7cokD+HCzgXMLSq1t/MIkJYREAVQChnWG7xvhT6fJ
YmFATENeNI5ciQZ+yHYV3YaJ8LStgadOLq4zHTgbRmIvPwsVow3v4s/vrs93p20z8mBGJvekF+Yj
GAPrhi0/IWEVUhhA/lOQB69bNUmlQyT3KTcALlRsqliu9h0Uu7lNa8QdA9NCX9a4aCgUCMAZoOAu
eHO86yuFv0q6prEpekCEgZeGVRlGlPoI6nqxOSkjRJUJ2nvMu3IIp9/8JOFKISpeF+qZygGxioB0
qYkQI2kcQQTsOlyv/w0DRU/8KboI9qKCPoJRB+76kJVmbP6hmktENCdxW8rcOkEJ1DZ0FfijuFDj
cZ+httEb/5urgMa+tLTV5GsM4ppxE7N/zzgD1b+5FBKOAKMj4kzrTVEbHbOTPOqpPXV5rvk/LPI9
khigu8s5N4wpoq7M/+RxVVF6b+JWECbVAzMPwFK/MeXlNr0rBfaBThQy/7RBIAqU1kKvp+tj6wXI
VSyXVbniibiZweXipVVASD04EuvoCW9e4uBbLKJK1jMVBw8QU7jNnZ/q83giY6am+t1Lw/0A+z/3
xEhXY1ZbULNY1FrbIsByBJ1fCVnbekWGLX187I24UOExVzNxO5PhKdecGXOUazmeIHC7bntK/Yo9
8BL4OXv3mSFQEWx3uMbKJyHx6kYE7SjYiTSYO3IlYWo4BJN6VWfE/SiBkMgLeI64Q0BvjUiQCB0N
epYkbGadWpSALxN1JNuyN+ASU9arswpp0g0iSiouLM7Hn720F1+iAcq4e0QLTOPogxpO+yHKEx/G
RJKAkoqMxmriXNt0yfw+WWDpWjSBaGspkBei03+sjiUdg4tMGKvG+m+npAmUJ+bKccA6X2D6O8Kr
iT0Y4iZ2d4QhlFgwgB/rndDt90kvpLZuTPBwsX4/DA3GZQcDR645wOXbc89u3Kj61ChXRoF3QLc9
8CeFuIEXIneBrMfKwYncDQuG+2d2LsdQcoXLQ6aAjLbs7bNQ8qlbL7UFmDdGFBrjtZbu/J0hOINV
DY4vzGATd8lb17X0cLmWGl4PxumL6CxRlrsABGNEQfLpZfkP98WkfDG7daxje2yGfROWYoM/XiRC
MfbtqGThMmEZEO2k+ZPb8OqWQ/oXU+L+IiMDlVDEhDmP9qKhARX4eUf19umMrhsUh5a2Bi/4Ywrs
0ffZLFzhkEJYbcQGnPQEn7MX+l9SJAh2FPkRuYW/cFM4NgFPERnOud2s45JoLruhPm2jxRwIkARm
8Q++8ZMwe9pjb6JD0iM6el+N12uRYs2FHAN90P8bZCR30cP+QvWhlg7FelR1+5ifBUFGHaXSH7yI
spsdixQVu4dDC85HcjZGDpo8usn4uCcLdtlNCHAX61nxSb31918GJwc4WLNwWZVFB4LdwyCT+IGk
71/P0EVbnOdcKfjrfHd+slUNDXYx8iLMsDr21GAodfmoexrkgQ/+ppIjOwYRcl4Ai8VmvbrT9PLQ
MdXzTG287Tbj+yC/Ck0ej4SWi5LfmvEoTTZ5GjASDdWiRl3uYHTfEFXEUVUeRErENMa02yqASVx/
NCofRNMPOTMoRBVpq8y+YSn0ydRlI6YeE1gVhlDuzUKM+0l2xi2fGJWxJIpxwRAT3GZ9IN77rAsv
bnC4SawoUwrZ0773sg/FBC+l+07FmTJfQHB9y+i96iUKstJuOtnKL05ki5XPh7fm/mQHo7QmMykP
fEKrHI+Yz6gQMFa9aoE58RCsrNBcbTE2J6rsqsIHCrw6IaZPjKZDajAWxddEIQ6YMUfe0/jAfKmw
LlbAagwaT2IAVSqD3xCd1RP2iWAHw4W3sZ8s47zkLH/L2JljjVOZfBrGoH0DYXZg/kOpPBssWUDM
QzNhlADIdZwgXXa/aHl9UBNmQ2frRmrJv/ZEZUSq/AS4aFx7Lg6HiUCFudMSTJfgkjfnG1Jkzx6f
2CkvRWoj8CGx2DOCXr3VUyLkIfq6vdDi9x1AjHXoAryOE83XRv9t7sYkvgDCC41FqeNVrhexhE/N
36WWSmJP47aVL33VQrmWnXoVay+CHz2aCYhJQ+DsdP/BzaKhmdeGmPZWZJlR+rrLrplyLPGxAGyi
S4MHXb9qiBdrZRmT0Dfd3/Bi1yewUvUGtelaRRJO7uMo4vPfkxlmg8EObZP8KPcXdT1sDDiF+RR2
mvwalqeUZkjjTYy7Wf71trQYpnOIrmObEqtwIW8co1Fj0S3qRNT/sT+5HUbaf1lH5yu114ZCkwAF
NU4yC+LI2ZD12MnKvuPrjL6NYJIHdDtpk7uWxUfG31tXMhYbEMUQ2cKjCqU2JkFkvpBzwEcwSPW6
fD+uEmmTqpaeWWJ+e/m9hAJco66r+N/k3FP04EvW0IY1x1Vr6+7vnUdpBu7VA7hsgkSQyhE2lyKg
/EnsP/QKcFfh8t0/2mIgVIFP8HbjdeLIXgtHs1lsHU+zojE6p+5321x9yRzOilvObVkL6VvLiQOQ
ROK1DfIheR4beIAUh2i8aO/x4wakGu4fI0jNvym9KE0zG44WcAFA6yjYiZ1dzKrlLw2R37ZAnpSx
2vD3iYGtELFJklgMtOItWj1Ut0d1iuTIRVv8ShZtQl98mKqXvyeCb3ZW1Od/3xn/EFEnd+kLJEXs
D1qyHbLHGCde5gRlZO84inJP/su1nZ8z9EPlYVjloyudQ18NX82wxDqNtFVGYJxWf4Qv/LJPbTRs
MJnBoPNrJm/Dm1l/jN1xq/EHnSe4sYfJ9lZgBVBWsLxF8k15HgW2g6bUQuHBoxItxL5h07zEAzxq
XwjaP24Te1e0/UNw+S/Jhrp2iN9cNHKW83M9lNkA81PTvI8KUJv1hisQbabZb4AiDb6Z3Uwhgeap
tHySgE7XBQmuvHUkPj9zuXU90KDFJFOemXltPqRi8pMf0zGq4j5mZdXE94ZAYiwGm1HIuRw9N197
c958UHZkAYz7txGaVcZKTykbDTW5/Nu0MHYgWau0hGDyfjNbp6orrr4cMtJyvuwhtnnSqdph40sC
0joeBB73LWNY1Z3XJSgCMdP0gzDwpK6XDyv6oD8eH/PLaAzFSPhXXezzEWLYkYENpYVEKGDKsJPx
FcapmSPv033AORxNpkZoI1M+Eg8pioUDt+kHmkAyMT2qxeLS/FoAekL8Yz0RXGJ7YKS29nVpPxBk
aV1QkohiNrUSac8sRbsgTNMD/15p+GdVipwnDYzdKn25OoJ2G28xBZ30glVVcNP+at0SVdVAKbSR
vIhRo6gxMnegRifNV6OyjQOGWcd1LGitNBUSS3/odG9Zjf5kem3K2X5mr9OTPj3fJmBs1teLmaUB
0bKwHmmRbSqR7KbQ05MSbP20aUoCTlGqA2Vem92grq20diA0c9GT+9IyoLT26Vjj4qos2xUHTrAJ
JCtZJxVwOBaLYEQmGwCqUfirFegCQDOBI3xqHp5y32Nw2gNb2enN5vmcEHfrcPz/OdKGWHNs6a+7
+apYGb7an/cf1UxCn27Lkg/bHsfGWWSX/uQs9+5P2bUlmuFg/TlbPkrTzSA4wBS0PBLaxig40liX
Zxx4d4Zcs1rDT7327O0DaiGcDkWrRb4EjQb/flwMf6aNt917/jlgQtL6+zrxZoTaXSI4id1X4Oz7
aHFKzQjbh1tBnNKljI0DZgTolnFFG3CLkjUbqqc8ocSPnKJoVl/Lpwe0Gyk15/nHMWbKbdtpi0SO
Ubc+2C1Ncr4/kVeoCZjOxxF15yOU9D75p00cvGztAWMfrEFBNnWw8tMm0LrTkXbju+lkUkl50es2
y0j57XmerpN18VOtX2VMZ8hm8RZb6Kc6rBKr7bZalnMlWNI0f1B6EINPdmKf5OJv8psPHpK0TMtf
MDtma8WtAAfDjZFcsb2VXNOY01dT7siLdDPpO2+g2WQlE3/ol7olhGXKsYfB/uCGcMEoC2Yrmy9K
Twi9fEt/NcVwrdGB8jCK19zSfxsq0M7JhqpMIZxLPWto16Ke9VS6NuixF1WjJaRgEWBcXwe1i3rb
2hsAgfDo4rwVcH8sVn1pXTTfmNNAw2JL/OiWZwEgW6K2/9P/eQX9ypUgak/WfLQMt+0SzUuiidyO
c5OLabCJewbYfpGFfV0e3TwiNMGkzcv6Wdr9IlDHr+VmoMBAbwqRYzQ1HFMpqUdMGguzzsLcnsno
cb4xerB3iAwOxw6nTJEDvBwL7+X4zPt+WwtfX8Ugu79wKsMqaAqRlViLg6xk2QbgG0hPUcG04+J1
o2ardlpRJwSwsVpHBkdAibIYBfDv5hNSC/9t4Mj5pm80NjAz4URRgIuG5vWQ+Q+jyub/J+d/wsD0
gKS7+cbrwabLiC19Oaen9zQTAL48em3xoLvdbDuARO8Ivkwk8qykF/XLZq5BiTHPh0ekRIF+x6lh
/aEqBxfRSjyDO/NiUHJkkikNZS+gJRJHNaaJcFgZxGMmHMzegzRB3xb4ElmJ2woY9baZW5N2RrbN
T0mIxLS9sfffoOlmiZRxmAf65dfhXBz6fcL+UBkeWksPlVhhlTGy5alEkd4ocUOKF6WrCZT5Aa8E
Bjd2vFhYY5Exzk0eASOD+/KEo2mqXj0PMcqXng065tUesOVgOO5uXL+2vATATbV/SA8pi1hL67kX
ebItEwHkojeyv0Jf8KTSKcseXQRifx3RSTOk6PK2OmGOA9nu4ULm+i5em/jnHxziG09S0zNXKG4b
pziQXugB8y4FagR0WpUWRMZ/0/L6MjbBlIa0lewx0zr3RTR9a9Zm/WIHL28URCVkFG8JMa9ENSaP
6iqnHZ4htQqd3mdVsUA2t5n3lM1/jnkzmpWzppuZOF/CRsoXFF4yhf5RJuwtNwT2ttNHBaDpwIOG
chYWlzSS/NBqykKw8MXIUQnd1qcv+lZySfRaTsEbV/nABdDJGog1Byu5iT83bxO7MhsFV0A20W08
eCdl+9NXHJD8WF6hvsfow+4rN0sJtnkciXjsIq+Lyt7kFMplKZPmubv4xZ/4PY9ruOtoJAiFjyNh
8Ypz/6Ma/F9BCPsduhgd/Dyeq6yB2wF1CRy4c33ltqYAUkkTIse6uWXqmS5tuVXqa3Ho0Q5DEVpl
I0QxkiCUxO2Q5v6jq4nThCU7cCPZb//o7Dq7WrtbAlLG/pHsQ/H4DzS//puMNfqPgRrD7Ii9TV+2
RkUibn9rxKzOi0oJbM5DddODTww0r0fLJi8c44Ee+ubL7UqD/MgOW4iH334aDti2kb67oM/ARJtm
+PeTLTdo35ZzG29gtJoh56F44t87bzYceOPi7+gu3z1YhwvrHx0xzPRIE50OffdpRHH958fCjfee
UQHLQa0mdNgRSehWZbHNrk+2Kvnvbs6Z8oZdquA2XoFTzTmyR0GVfTsO9B1orQXklqns8i/KSiDP
AcgygyJNgAtiZWSAkOD6/HcA9t/GcLkak8VqloODPvl4AvbkD69cFZ1FIS4v9ZgluX39IHDcFyEU
GsleUgjqsjMsr14R+olhDybV3oqEb2JIpydLN0zCRF51wB18tTODc5Fs1UP7M6otb9UR7P65j1kM
7js/RJzsP4g/MNEruym76Os/cb9dPj9Ps6aZ66r/xSlIbrB6VVKXHPH+0kcS9tgYn/3lxZsrsF3n
wxx11snlF0N1/5MCCUoBi5BOwP0hd8oTfcCLucNldI37oGugix56jQKOqhxn5770mR3Ivx3r8ZDw
geA8RVmcv3SEfzxxWBpOUKCB3FnjB9iEJI85iNWfOnaMeFuULHFxa5iN5ouE6EeENZgH3c1fPQOw
zXuYBXeDOjKdyVgABt8aWHGRhDY3EjyfMse82I1nSmg2Ymw9KqS6V+UyKBIzRhWg9j5e6icb//A5
bxOnSn8aoN+tocgyZkvydk0EVnpEauriqzgsJId0hnbEsITYrZfgoXAgRHV9yL01xipC1B2X77Kv
pYNC4MEyXURIt9ve5mUQ9JVfM9xdfMHxvBTAdZIRER7MvgVLvgWDo3aS0/gJz++L6Gtlfnwfth8/
8n/j7fWrKsi2ULqnB0Oys4E+ErjHabeAtFgj0xuYpARxfKlWwbl/VUThW4ADA5na4yqddGsCWFLk
At0Y4ZxXbmUgti2l1+I2bjbox8jW2yp13V0emgqwtUlmvj/ZvFrhpLsn51gmwgeIiAYtEecOTnnb
Ipvd48x+nMTPWs/+d0FnQknp0WQipHkojIZpbAm9Y7Q2wqJIABQtxJ8jxCzYBXajOk6dPooixRmB
fGV+DFptlOvDqCn2EJfHYG4AIHGGW2WSbvE+Pe5FFscO/WJpOsUM2c0B/jui/hmZgV4x/3UfwWJi
i63l3TcKdMCzJ2/R6qi+QGpG4jR38pmLEgJzd2Ikqtwmktds0fOA4bxFpajzytAKUxU6O/xRGycL
1VMc1xkQCrlBnfwFKMUgnfxaRx/yKAnAASNLek8Sw0i1VdLYSMdIRHcPKzuNfxbJQkk7FNMRrk2R
+2FgxFUueQTKdpRVUn5aQ0XbaxLrIEnTbPyxHIWIplRqtgqNC+MKU8p6Y9avOc9tyXYZrNp3hbTV
2gLfdZfgBcr/w4he0xzAaGTrOf51OtiYJ6QUJ+ZjB+odNTsc39bOtHQiJ/N8CqWNw+3i2h+iBKSb
V6+7SElIkxZdORobn6TE9DoQsIL2ItgtpdRK6Hztor69U2NAdl/8vYtUYBRIgg16uZjZszQgsR9+
Dcp7mTm/cXXW7KJqhv9Ox1sbl2vaQ7IHC1P075PDyFYGmhYX+J+uUCOTjXhii0HPfSBPZL8nJITH
0BLtYQ5uVpzsKBTiP2Vxytf+dX57qDsWGjbXyJ2YFSX85eu3GI1eWVl7Va7I0hBND00BlnvhT8BS
pV0Tml5RRG3AsBHoDdrzwDZGKmzY8ZNmKprzQW5JYTuRs53zLPKmbGJDqdxJgCkxd0wrC7M78xQI
irfE3FaFN+xpw1tAHJ8c7YFKdGKWPazt5e8qn8XPZk1F9NdoZt9Lwozg7083tSHVz5AD67OB2MUz
+JofrD3vo3KX0QlLM9/K1T0fETPefQ4NDVMyqmXGggcgyFXld/P6QnHAdjNOrMV7JHqL/l2QFCu1
uKYCsg76QLovYrZBtKDSCLZS9bB6j/Huj2vAwMLMBxRkaep/MA/CMXss4zPwzTKEpr75IN9unJbT
BdUBnX2ufj6Vjb9xXacaDe0v8WUIplqH17j9I7OY3V9pxt2Nn3qWTUjSnLwHtewXZC3mJzNL9J77
bdKoLbJGFSuExZCuJy1vC4EsZDDrjdbcQAvhrPN8W4O/FjM+iYdLP0Vi9Xy4r7gV3ILidiHVY0CN
BQkf6f/Xu1okz2297L/t/3Mna8kgGlMOjunjnqveGEkKXG4dZW7cn4QzvDBAnkcYEOVC/xXGjNQO
HJVxZLcZ8Dpwzz/WWtg4ZZdOG9koVXgDOav5/uxjR5giCvhXiLtyLY4C9ackqHV8Lfxk/yXwheof
rRTmLew+EI1+jS/WiC8IYiqzi9j7M6JnfeBaDrqZY0vJMqjfRw8dIUCE2PwVDU0BTxF2SxFcCTic
2/kdB2wP5DJbYwD8pvVj/i8iNq6K919tpEZJlqaLTw3kn8MvagbNuzoNlxdLqBuKG69vhn1Z1uPJ
96i89o3tMt4OOWGYAWRd6kfQgBZmz4Ef3lN/V3N3QwcnfwCm27t/i3k9Ks3r4sEwCl5W/i0O+1Y4
R+nGs6OXNLl6fzN8TBD/s65HpY2qS2x/8jCp1zFcyEX/Ulh0H3PiayTyyAcJm24NQh5LusTGCsPb
7a+qFfMJdwY8OUUUhE367wXaYsDELsxd+/ra1uqVBw7u+ufkpLnFTtdPCJSOb7xx7zq9AMhqw30q
bISkjwU8R0GkersGTWTB1AwyvuDDhzQnqMZKbV7zB3BTfeeNz4YFSo4ADzBkpId8tC4QmQIqbDwF
lhaV4JRcRme6eb70CdQVunSavYNWE4c/3DitqMjePowV21LcjTXAGsLdy7bNbcRchJkqMIXNrVBL
Hzgrl+xU4gkpgoaNmiF2+/2Cgm1WbgpjIcuWf7SswHF7QBomG8svdjaPfgzBDk522mqdZU6J6592
tSn2jyyjKQ8/dtuSuIOd7Mgx5vxgo6YTen6yDihApQqcuZ44HWNIMMjSqhHHlXOKbbqjUWch0Tao
F4pFHTJLA3kDs/ZJ0hIjqaURPOq2wgz0NC1rBhOAJFUKmxd2bPm8tl/lU/8afAQbDSCKIzG3LILi
74+fQhe47uS3aNpQxaEMm1QDCz0tKh93obhqsftNZgxYu5Ed4MHkQZbEXPiHORyFC5c/3u61GTR5
jXQPvl3NV6KmES2fKgofxV/5lgc5hAKptJ2ZMJKj++wQG5jTqgkKnxNz0GYFWY8KkW09cqnPFKPV
7tlQOQvSHgnryjnN95hcab5l6tVC6gGrL6h3WqNoY/DHKKOXAbPv4LMJu54rrxrkuqlm3fvyezkv
JnbWxFBqflPsvLFS8eKJ54+i4IrDS0B54kO8OlAA81mgwVmLC99JIOq0DT/L/Gk9Xm64A0YkBTux
nBxUfweR7GlPTKryBFum45LuW8CY8iPjpsI1ieopj+EYppCgdJSGMjE+AMOzsZb52UkAW51tx++0
fdXF2yM8gDR5kRm+iHeoswTKvDIzFsrSOH5ias2HbljxdDAoBx9P+ocRoatkhQ0afp/76e2YP2zh
lOtx2nyREGYNILtc2F4y0X0NmDlQ4FMrPpZnFy5uiC6340dVtFgycM2zN1OddhZHyypBBFqiQhoY
gKkOEovu6aiGySdVi/R0mWr4RwrYzNG6Wdqwhgz1H3vGqiNhNKkhW2L9E/ZjHcZTKMo7d11o4Z0l
fVjJNI2iiHbLIXkX8w9FMYMY3bgBHYRoYr3lwKKMAFc7XEd3prCDzQ9y2o0wKJAP6S3lQ02ncHd4
6fNtY3ca38TKDKPRU3z5wfv9F2IAEL4VnMrVUf22
`protect end_protected

