

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
MpZqUX7RHqqBov6r9sp19cCgAmwWMQKz/kilwg6KfQHVNd7thNhiMjNr9jWB5lhCnXS2Dmq96KWe
V2+V1FG8hw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
eHZEt9aF2k9bUkzJgCuA+q4yfEhMdqCEDNKyWFDaQseZ/ofqbFQAQc2uVVXTRkEXQs+GrviVm+j7
2wxr0JrS1Xw60RqMKKhLpfqRVe2BmFAKgU2BRL0PnA5WtTOSGCOmSJGfPa08juK1otVgwc2Gzis9
06D0/bVknfjjRpJI8Po=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
s0TU3tsqHiK9WgquIx4poaAXQ17I+2l5Vqn12DnbEwMyPpn0YeINJkDaKFxRf41aPK1Wkun6v9Z/
YYZDqYBgVO9Z0NMkbD4LC5C9cZSBdk4ezqdUWACnMS4IR+6qI0nvPM6pNZernzgmYtMGFsG0h7AO
2CLMNIzANr+bYhHkAqpdx/KPtV7Deh8xOAkQeNSD+8rjhU0z6Gg+2FjdPjkTgWwsP8xrTSENuxiw
xPh+QM3dvd2tDQbC1sSMu3CzeLQh9mMzJ/R1uFQDv4VC1TFFFPI7VMPMlrl3y0ondyZNERO3SeHy
Mn6aVbKjlR68QJuFwdsz80LSh3ZTJ+foTk16ug==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
uIfIqnJL93Nk48nDUNvQ46MGSw+0jZe8QEp6D5vC3ytHCm6yvGspxOPTR0O/6R1kGtbYGX5AVD6b
KvoAJRDP7Wr2E6PTOWfFxWtEHCKiApDz7UksHM1gqF0d7SCMfsYR0KKn9LnLJiQxmEJD5y64ve5y
9s0qEeMi9k4HxMVPc9k=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
XH+fS8ngHwfDFxF50DT7MdOHeXbY/uKmg7Eva1j7eQ+2X+a34Rn17d34wKLf1Z56AIT4ksXzo17E
WT5KT9rKAQNao71yUm+YQAunOwqKEPRyxOz3bb+3Zvx3y9p+F7xTeZFLan3KtqwByX5rGkNJtGjN
oI8H+T5FEpTIirQ9oxghooMSVVhKX8RsayssyrgajR3SSX0Q0ggoCOy3XtjsFKfrcDNlt7iEsMAt
+8vV+volJUxGGSYbt9ATDx7fk+pYKVnFR1jV5fEpxyqiZQoGjkjsnbN29jqgiZBfhyEe2uAb7sF2
RnfrEGY96pFoR0k3gse3XEc9radVftI75N7ROg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5808)
`protect data_block
jjXWy/yfHtsaqReBFgNyV5DW8vN8ln7yW6t1xIWYrhFSQ/9rHO7X5bsPrYfjE+c+FcXJBYAvyA9F
u+Ukn5x2Ha51gU3Opqw2MnL6n32IAP+Sh9Xdd55RqoHiRYSovDuucUXhiCPi33gksLVTmDDxhBc9
S8tHL5gqtqVXS2iKdc32X2P/6f4jr2NVzbTibCOHb+ZHy/7eD+cFvJGOVbp11ddW1OwpUuV0rlUj
TtsjYjaaSyr9cXyTTwyH/aUwdzPQh2UHdFQ8m62tJ7sX0psJ1b9715o2j66OVh5/dpOKqlbdwPCt
ocVUyOGpXJG5sNiNI/xPFbVxjssew9lW3l3bZwgQCBVk6v/jfC7y/PYshnYY/h4KH7sp/3YATz47
DQ/hBtOJ6BWa4Cd1aFumx+z2UHFqZte5wlOfMuXM4SGxdnjqmrv2Qolwn/kbjYqTVT30noffzBfe
0dN7y+K3OEC+6mmBou4SsXrKl00LV4PoQcdyDDUFAANHiIPFiNZiwo26Lidj3/AxmMGAzBg8U3LU
ZHHi4vlVohWLFWIIgF0CDBw9ZzcADCaqLKKbGWVaQZe+naos38ATeyqzUHRe8Rn6CRdV2EUXpjdN
t0QzL801KjxQyIPNRYberk9HsfCfsBEg+p1Th9dKgilFcpyiBFAlRZvETS6HrI3738zyTYhH+gxM
PzHXd8jrh2OCHXKLjw2HHv471c///i6lr0BQCTf070UfC1dhxgsymXS4XUVqou9lICgr1vwBq6WS
Nf7guHs2Fl3SiACyaA7EqAMHLfpL1fcNj+4ycmVb9f5He6g8h8ST/+GO0NI4/2IXnMORJXeCyVNJ
nZRj9uwspDPZG2+hq67FGvdgFhhfWPTS5Uc3FNld47xmxg5VyfYg0O7VkQPbohMI4ahnolRKOFmA
7qDuZqHdVu72BaBcgwkdgZdyk6oS2knbcVprXDeRn5TyfipYOgZkIrXQ2TNet/V1ftcjlEsCRlXM
fmZrSjpGjfV5gRS68KEK6tzuMc3FcW890q6bxe3c/Ou9kRSbwKZjDZJU0HJo4H5Z47wjur9Aj0hV
EH9J3zQ4rcVm28OfR0ltCamoOP7p7Qqc1fSfYBrKbCrg2CgUDKznbJzpdt9R+VpOQmBECLP/oooH
NWd71CQ7BCoGgvdPnpIGXYsgeeYgNIQertNF6xVbshV6PF+HCFQRhPDX3XansXFD40atz12elH0/
px2FaklhJxOxL+VpQ61Uj3ay3gS8eJ0uqrPMz6Tdpczs/eEkrxkHiuXz5mXDHsC0z77uHVd/ApXu
GHVWlB3CVELagzJc+fE3hMM49nYsTj+prdxxv1sGQ8II+Q2cFY6ceUcp8voLtFfmdvfki7EJFKXF
aw1UmAIDtHNU81JsFbQvmZy0uGOtYUNJICvDHgRdOVgrwlTY6OBQAsUMit1a1g28PQ7e3Qak25uQ
QIESfzgk+pCesNszsD76wpy+/3v6kZRSECa0xVRWRb5vJfapPC75NUrEAeSnCCVWZv/mWvs4FTyJ
LzLrGL2sN3duRmv3d7a2EEjp3kH+fdjvPrZlI7Zah0V7wW/+w/lySraX9xFjNIGhcsc+xQz5j11x
kL5XZBs5BHj7lhs7EbJUoPbgWtUuQdQweGXiuFARkKkz6/BKpMmA1/agktS6us+ZOlblPUNDWeuq
eLj2h6sNrxmkkr1KbS0BgIeo3EOeJrCVhzo/37P4XEe8lQ8N2J9OA5KgR8BT6QMbRgYxLJdtjVOW
F9ABz1fYlkUNTQGfg0cTrRmZXTwd1msUnrtLDNQ76nm6IOBE8hY8h7VWOhGQBaGnu2qPY3suMteL
MKtFLp1yWt0Fbjm0ffrEjcFNinRxd6GqtiK3ExPC7nfUnEbufbj5m40L4Ihjby3xcURsRlZAoXqN
Cw93lLdbNDwZdOWNPipD338WwHWldKfsPJsJYuZGY7SXYlkgf9c8XxXJNV91b/dwT6nsMUuLDP4E
fdTkEyMd+SvmZfW5VbC0vR9n0ZwMnBK8cqnDFRnEGBqzHm5Kyzv2rI7/co6q5oI2wqkT8XfdV6k3
mxqSzO1nkoWws9emLFoyigkdL9z1jyeAuh6rZEHU1d93+X6R4cHFYmW4z/JWxNwNKZJa3SkTzod5
4bk0iyQV9z6bLVPjaP8jeFX2ICi18X13Or5aZaknpQr4WECKQ5/5hC907tVzZKQXYXgSpTYQcuom
CADVxRn8j/MMRh6B/OGH/smDhItEATbE+t9Hx4kyzSZOqWNSK0nHdzmhPsomgpZmzHsGWP7hkdqP
+EqIfBo2mHt31v2VmeITpIW4Ev/N7PsRC7SYVoHq8eJL9toUXaWlpTO3b1kuvsi4h/1cnbGDxrsF
VCX5fKHxoL01YMfOkWcT4NnzFvyigzLtliSi90GfUSVwnVrcb6WIJN4GI2oXIgJZe22HDXuo6cu+
V1x8jRE6ZFck4DC0tzf0LOncFz+O4Z29LfGo1T/RgfoWiFJUxjH6NcdMdJv7aiIuAfmOPP+tq1S/
N7CeI94PJTwRwrBce3UuIG/otkMVtihB8VAdqxBp6na88geevFrVWKtPfvihpIuOo59886BJlK/H
HGyMR7U/0z+klXmmf5Lb6+qaSWuOfahUiaUHwmBuCE2yZq7JxY2F4QpG9uBXY7STIOOjXex6TSWT
6xcc6rQOQK5mRoq2LZDw1ZKnxbzG9cMTQ019XCuqnQrbPvDv/iQQAS78m+wh7j/MbqKXs4PTJqsS
u3iE9YDeEBSr43QDklLhDE8+sH8Z+kW4dueas80JXDkS9LctjnxrUJUv1vG2TfgZcD/HB80Dsy1j
5WC8DHJW/TPCd8+0M1ZqepFeHY6WWzmCcD6ENNoQxXbK6P9tKJXOXJw0pl1yBQoIYRw6dxb9FE2b
vqdfSgGnsWExSB0vv0dNh8cuEn+yLiMuJBIs6lF9EJB+pSdJePugH2j6QiAuriApQCC3NbkOYCIh
o5q7UJ0lNOss9bzhr7MExNQdAHSrvUnloH8vGaT7Oi9uIYpmY9Hw5VnlM0OlbWh10SyIyFHPNHiv
BZcBj4yjEPLVk9nKvgCK3bPTY/C/c+6uJ4nFoo79gU95JfrxgqYW9iq6JvNS78NvMdDxhLXL9kFH
ApFqKmkQhW1OUqp5rNP5fFIouc9FWNmfxsfYSwW9dpITlWQm8iw/Tl9RI+oJugJffTYiNY5zuMV3
XRraUIhg6e/SSy60trno7PVxCe4BUYEEtZnCXVM2IssSeBNx/NVH+OFo46OqmAgLlUjiQyi0TI0K
kD3EveUFXL+X591hi613l1xehkcgUoRIn3acD6bgfd5lhI0Kvm4YFkh2fgQMDo5D0Jz6vwFxe1ku
F8EoODUP3JMxMTaBOJajxpZU53NC72KpWlXVG46e2TniScVJoAYu280DsV3IhPy/rEUlgeGpkmMj
k2TFBTadBqUXHNkKJsu7oscxaY9K9IXir31KAnrIGzRtB0LQApQfr0xv1FRU0F91YNypNQiLCkdd
Vw87kKYmfJ3S+9PyKdtmfW63QN1IrxTfYD1oPpJZu7Icj5sQhkmYISJWvPEIQ4OmuAeTeytcGD5r
KMcmTAy3Dv0kWdjuMiI/THiEM/EZQqXFfR8Yu70119puceCP4F2bMze9fGJQudj8MGr3f6lEhFy7
wVe9vCguwrghoWWaGhVb6vm8G6RCS4XsF8P1HCXpfB5JhxhorH+HYGQJ8zjwQGpbEMIaE27ylF/t
o8Y5UyjExPi6mVtvIF4ltMLsdTmMUrb8+blDlwL4lKrkiZi3PgP0zp1ffHn08uQKCavO2VBdGtuP
M5gZRORv31ojxb69wpR5VOXCYoiAxZo3xCxCOiBOioktkdRq+ljKIscUjh+Qrn1Eb7K4LOocl3Ev
GEvLins/n7bsLSyG0QkqjKUXzanSPFxz5LMAAxJK6B6qnkyBu59zy2PyXW4uFY7hlRJJuAeq8+o2
XTdKYobv89FP0NnD6v861nWhCrHj6wmap4kg1JGdQ4ylsPkp86aVTyulEhz5G0UJuj0lqPBGR+Qx
e9dwpVmXifWQVn5AV2IzI/hZQxVlhTS6Jcwne3e3zlPUA2HDFlsmstpgFUsw4ycnNYRxTKey77Hz
oRIeNObhZv0zOmzsmgGjSJC4jlbNjP1gXtXBl6FcDBtQjyCpNn9vCu1S1xu+3u5Z5VrYQF3Iun+o
zniTSBG1ptPoSTQoIkFTUkdcDY81dnUT9/GhHUnE3/DmoNF9TWJzFZk/mUEIFv5rXJjnd5gRjL6Y
SCkF3NXUvcxSWQcm4cfCSOGZc78ie+WeOoanwx3iScDUCrP867UB3vCwC7Nhtl6IImCwWI+7TKat
jMocQ/ES1y021cE9/4gd2jp0DnVnaB+U7E5V/rJiSX5pQq52rmQHlXQs0jLOgiGX5XvsU5Cew5KN
L+ILh3a1I0clRdmJOcylE3Yupd+t6TyQuExfRm7KbDVZv94Gmy4qe7pQXjD8ZvZ77TRjzi0Am+DN
cIGlCah5CpqZWQfaBlYPfCeIfSSl2mt+z+ruaR4AgsBNEoCgnyF5RrcpWXtMc29GfWO/KrG0QOZz
m8z2dj6cNS+mBcuLnEeaBOwxylntWDTwckM4DUA21rwWBeAjKJugwNuvHl9Ce9mjSxDSoD3EXBQ3
oVL46kc9mTjLahdBo+jgI1w6l9ZhkhTqjOGpJTXr4SpFmYAKWKuzP6anhKXCnzZYaKeSUcEn8b9H
2BUaZCGLi9XWGhtEK+XaNxKXB90gR36o2yW3ydUAh+WHnMvDthJRogESeMX9svOGHWsLo7TnfFVs
N/G6qls9s5lQcPZyZDxkNkUtAFwkfTOeHxB4yWq+gLxjr0I+FCc8UPtmPXieo17ypmjxy9h2AogZ
4LrWlowJ61N5lqWtnKFVUyQd6gCOae4Sdr0DzyGfjFz5vMrjJChqhWpqmdPwo9YUN61tnIowKD3W
sxoqpUa4lT2NnuN5qg5YFyVNW4CUHERM8Z3CE6Si1/CGHDEs609sGfu57GSNAQUb+BVHFoxIJ0K0
g5aknAcFtUrWQFDKt5bWVXToHS7H9b2V4Kenq6KDQfPuNLr36M3sjsnKDNAWlH9sDenaKCWyqk35
Jc8D3NW+8Wed8BLZ1LXjZhWubanQS8UJg33mg/4WEINp1UAQi2sZEThq5v6E5bKxbZm0chobbSlT
NZEk+taNHRTkOXiLZyuVyLgkOf9djxA1ukni3MJOt9NY39BS3Y3RLQg2kigBRkZ2diMtD38DaVAb
Zhvzd+kihb4N9rQmkm1axPA07+2Ay9bM8GFYS/nBv02ttXwwmRwDD4vK0A8OgKQaSjyFIqQ4JOi9
SCmNLiUxcT2X4O2DgDZaC72V5Ziqux56uG44mIYSsGCY2pPHcu4Yer87+HX6c/OLsOGiRHWuLScw
16eAnTsC19/5EIQj2wlxTaTMJITxPk89wcpFL2nrNz87JLhVAkLMjLO/aZuMM1dkG/fSqT5oWnjr
fkxb2VIsCKxW0haPPUmk4tz9F3mTxkdYMP/ckkgrqr0hvCMyknHFBQOLzZa+M6+b58q8HOpSWh7a
tPPdfrzQlB+VE42B37iaCTmb/c9YnKPYlfLLcYNJ784L1IKWKlkdVkTvnQdK4V5iWYHkvRJVwKpX
aRWgyedPAKdQ5ZaW34u416F1B60/nWdAs1t2i2SNeJ1U9LGlQ3zbyVpCfbnaLm+4CWPJ2MikM8IJ
ngSMCvL74VnRavjbI0Db+b3ql/jiRsveO5BmnjdCm7MAtRFh2pO4P0t/th2PmPobZvsLpxJaVi7T
he4k/xwbn9fSfpeOS0FDMRJ6QtEoso8X4pso4gACCu7mzMda5hsQMq7/NoRkIK/WMlY7z0wbmk6r
R1KQnjHH1D53Sy/neBgbMV0sfF33ysgUbXashan4IgmneWwFPRwJlB3QxGoxJdQzZf4Jlmupt699
FG1uROuEzcAqY9Gk/X8GCpsrk3YaY1ZWFoTJ3jq56rJIaCqzLEMqml3s6opYWGbxhjRW/T3qiX6Z
TXTnp6XHbcP3RLWPgMX7egxawCPRCQSpaAJlTzc4LyObPKqLwTp2U1mzSRNvVaprl/Z8d/eH2TUW
tdrXNuIJE++pK2z1wJz/Q8dwFTAGcfQm3c814/7XiZsMrdeIh6NLoUmxNpbsQji1BOJ15CVlz1vf
NdYXUacmIBbP53y9kVW+v16nTBF33J+4lH5UOI3y8x+xVB7YA+YoR8rWF2nliSZACDoeOVNS9CVc
TDK6R3hpMhmFAyVd088NlTDenAG80ydM4MbL8UD5cdoU/wzugoKAAicTCMDVnV0qq3Nom8bvOD8k
0tuoYK9Eu5N2Jd1yqDRALtdUEY3a1lI5gg72QnShz+WNgq68gDLImvlpYz6252S3PyqdqT89U41m
hnkzuYo05+/zJwGZpdQM38V3jc94lti625QCeGgqcnUYDAWxLOhvMIMEd1BjPmlXQg/+PFZpYqRN
8HyzJo78gOoFenSV/0DhBPA1U22rh48bWU305wPnjPNVLXi1QtHLYULCdf3chGGe+70F0oWwOpQD
wAgKfqiMt4P8g1puTpHXr1ie4ZlhtoXdDYyiMzmNFMwuonJFwhS+6lcmCpNMGORKpd7sGPbK8n7q
/HoGjV6TRQZeYSzM1d78m9kQqNgi9pX6EbtwanW9J+MIeKrb44krkbKUFM6sfpWNwzl10d2SC6NR
rk0gG5RpyfbNvUrsNlMqzTGyR8XfEqKkOgudic5QfW1vaIT1TcaRnjBJ1TYstFKP4R+q6XqPVxzA
QiYTOO3xxkXOUQoI/Ntx4Uk69RgNcH5f6SBOjAlrtsj7UdKzYX+G0QG/MLvlGoYQxQL9BN5upf+o
qjkL2rmHR/4xbribYOdIa0CsPSs1WVYjyZt7eRMzsQOINASxbMggqh2IROvm4lZWBp/3AiTC6HN0
aBfUdV1H1GLmZjbqkhwH1Cw/LtBxTsqOfXgbjuZBVttSHaDx1gP4Xw8wxe98HIkyFfU6UyJiPbrS
DecK02gbOoiR8XgTaGMwYFYiZ7xs1z+9lnVcRW8MSklOkzBR2ZYjxHgg2uYhi61BdloVRmLCnKFQ
Fu+Jdx5yu6a8KyajFTMQRiaGcxUJQ1re6bM1VdHhs1MNJWXXoT0Z0K4V67KRhlgFu7gqCBRWku/7
lLitl8fa/TUCF0Wnnjzo642o25CXAr0wHxS5GH1zmmW2OqvrICuJZlb9pR27c0CN4VvEtss3CHuE
VYXVGskfhNoNis8DRCRIkZPLJU8nTgBAp+LCxE+X+Ioy0FdyQ4L181paD3WlO/TAcpnF4aayw+RN
+Y6XJ31YYpXvFgry92jeVYNZO+F5kvj5525ZiUlk3UcvrT/ywTvK+1stPsEx7oqUbc8ckCL+EIt4
7iOusbiN6QpIFmNe5fbQ0VwHBukYTb1fSppUChB0JFQtvoKRpi0tTM8Oo5xFtpH8Eujjxy0ZF6td
1g/HqnrGna/XXXdT7/2TismDdPTi/aHQB0PgXLecWTVj88LBAyoAFqCL5aoQ3ySkouKs2j1Ey50e
YfPlbfeWMXkJWQxCFWkkZmoVyLd6/zU74OLDGFRvPdbUqLIolqc+WHmkvneyjR0NJwRuOJtdHDhq
pH4ELlRvBBb9M3KJHhZXjVM6SXnE8R08CBzgpN4L3VJVbSlilkDpE/g2uuIwxG1gs+cPlQ1Vr6Ca
8fVQGfyoLt0lHwtWBK0+eb4NuTX30k3sgjFofg8fFs12vHAaeOKPqHO4wiyhSF2UgpIv
`protect end_protected

