

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
SQUyeNX8cyskpzvvW2T3ssUGj6xZX5vHX5fJU9Ms0M+rWpNjMO6za6Zgr1K2FMwHi+buwP0Gw29j
IKEYpdzZOw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
hoBaDPgZL0nmY18FE8yzpnxIEfx7SKisNM4FVo3Ao91EGtVywU0Wb7yA1enrW6Xd+oLWYcrMdoDX
JTxy8JdlM3o+jyjU7UKGIkB+vX642Q6fBAuo3SZKPKM/RE7lQknQIOi2Y5V60nbw/AM6mvYDKdTS
wiPRLcQIZpvU4dn9GkQ=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
o9OFQKQt0GaB68TjFqZyGwbFj1TRgCs2FzlOtaWTgxoDRMFT9IEssmRwHo9pwJ5Tn3OigUlzbBbd
XTy7vthduMEKESguEgGeFDAlZPJdvm6/cpwtG3omF99Y9vBxA2K/3YI0+jDh2eyUvsHMcDbQ/C2p
zFKW1hcipARgm3A9Ys4mkgzXMVKYnvnQiSsmezjrXPsPy8jbFYPXFd6vFSGi/ZwrKMMLLNZt/Boe
k/Pl01HBEt/KNoY9VFx6N+e2ufES+vAz0H+DJSGPch6YdjmhkZUj2llujVX2dT6EzXeB2X9+1Sar
qYaNJFQdqXN7nDqoQMCiwqUZBJaHNrPJdzAMcw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
gMFEdGC+ckR/NJmX/aszkYoB651qUCnYvXxq63Zrpc98jREIyboMJaogrhiyZ1kntx31alD51ug4
ZAed1vud+wZB4IN9oJ1STjbhb+Zj5u4I029j7Gy2lllPl+1O8Em+DnBFlaNak9VTW5oxld5AFJs/
EstFEKIMT8MSbegVIEQ=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
I2MWBDnGcReW7SMjRXdvt63Rjoo/gu+NQcstRp+eRPxV1cdY3BaChhCXefqNXs4HwrSwjy6eXoRH
K9pkdKW/MmeSQuCCGBXm3SZnri7VuXOoNwZoR7yYcuzRHYCe4OVzWrXYc7CJVdShI1TzYNVzTc69
N+748OjVGLm080Ri6+7tnRVNASpwPZfo8iBz5hClukZRieQCUQgdHIAZx2RjUyVQaoW7cJ/urtOZ
zr2GA2iDsweYcuo/xtEmVehzY9Jjyk+XsH/W+/8SFJEIN/wAiWoW84/gDLItkUU21xaixyhQCl/Y
sHoICo/iHc8aTOV1SPHo9yWYmV0UZ8KJqveuUA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 6304)
`protect data_block
SgfRp2A7gPMpxWIoKx+SDPtxb1I67d1kVO1fjMd4CiJkMRY/lZVtMQxW3agyWF+UKhAKIuNPTWlI
o/AHVl7QwvDd74ZQW4olvUVDt+FeVyiHtB7CwtEsh9HyKiDYNP5WuunHpMm0QkLv3pdfYzduGwcN
iKVhQN93ASife4XxC3B/Lwpnuwwv/T7SQs8OUilQLBMaYJoGm5EagHU7yXAvNtZeGybvIQf+/9No
K8ufx8b0KY3MBbkO8CzlLmB5x06H2Y6pmmOnn5k0DKQ+gskNuI7WXPSob3pIl+lVX/3cUiWsxVTz
0W6TAjbJ7ogDIc/qiVSKDWkcIIm2hcmwSi9kqKlxguO+u8l6slwAfickzT07EdrykLp47RhTbsAA
DvV0Zvjk01QRGjPh0I+7MvfMaCEy7CTOMZhAJO2RDhmEaJOoC6+disPdu1vGLDa3VIBG6Jnt+s2m
qJ1QbMrob4RIdrbklTZqP89k+5VvgGL4X/ncKU23YRmFqG7faErERsLB/fMfIQnhzt0st2Kyqb3H
//t2HOfO0u21opEka+AixPyqFoXeKolN023UJPxIvWKCdrEHKaD8eoSRMwNhuNCUc/xASEgmKLAn
lkMAu28GQVz/1P37IPqchJIzsk4X3GGu6SGJGRXE3xCy46K6b0w/VWXQEQVwJm4yX2bjfIOlbrhL
rG3EJj20yJqoxqLSQPjCimU88ip3F6C1FtJd9qyxnK1ktTaxZw5qBZNWbIb7YBzxVPwoZc6XRlpq
2ttIKgAMzBNkQvSSvqFGPoCH/NrVVocWxj74U9s8XzB+5B84YZOjzOCkZWaEAUoMiXPEoWvD3c+G
iEfPrfACWphbC1QNm7zzrsP6WCodl87ah6jtqKEEFV8A6+tnq1DbuP5KQuj8dGdRrm7durQFpNQw
Z5N5dSVmHof79105KF6o3wET62klJl3lQv05ECp+znX187RYtbp9+TAxdd8gTGNKb7MZjWheBAFK
+SVLt0jRAgRmxXoM91saZ+BfvbB400O6C0ewg9eHvyYGxtEFxSHAtv+AR5d1emUUsFU2bd+gay5o
CniMdDuwarEgIHEBTlMh7o47P2h606n9CTyO4t0JqPpI2wkU66d+vFOyJwHyZIY9HrPezaFJ3lWZ
IFB0N9uyDmVhqiPWFNBQHp1Os51hVn1cVWFXgNzQJc07UJmZBDyPtcpOaBG/XLThYNgOkEGWGK6L
MuZxDJBxp3QQws23lEQCC16+UtRhMa8tdC4hsplUP1L6QnmBMziMzl/XCQRQUvg5MO+DTGE7yPcx
6v6gWl4UxG1MxBzyQrMAJ6+8W64BGzSAfk6SmvLuGRCGzr7hGam0mKC0FSKBt8FgWSKcin+pzWqp
iOV9DTSA9RluAxLtTKM9FEu8D58HWy9OUZgMgq+71Vd45cY6ykU/kVtK86gy3HNoJOcmAau2bbIC
nieIjQLh8JnkBRLf1vcxmu9Dc9A+AXLTAd4MljdTTzhczTIw0DLbtEkmqsAO1HKjnRKle1GQ9WcO
pJsflXM/KHI1ZLQdXE4fPnql88BhVp+O0bTdBR0I9ogm5VNdK2yo5App8xaEBElnuUdRCN5O1I3m
mwzBK+id3fCz9htmXAAg7MVTt60ohjEXd9Gg61r0KKpL9TjlGcpBTrNr1Kp8f25aK3KW962vpdjG
hu9jLdGrZj3TnmvdC4ZhvPJqGZGhLwpX0yVw5pXxXyhc4gPpnjMZml9yhkd6C0G1knqUZzmEtrXg
W13h9CAB/YK0v2/D/aGJKa+k8DJQne7XhmMZWCTESZPTVXswXHsNiuyfT1HqtHY+K4YxAgkyrr0O
Sb5JPC/6cz5IZ2hBrk+ppuvf4+y2LnaW686KVhvJMQM7opiDQPffBVv1GJ1lkLcal69LyfUywALI
+ngqmwPniWs8dEQT3h9d7bbf9dac7YDBlYrtHWJ/Fb0EyWwXaTIMrZGLZlRZeQwcCyIumyZX8vVc
e115oebxIO0B47Tn6ATc+UOlNdHZWSSmvukXjk0l4dTTclTkFTdMZvdbyk607aoawCUUVugtxpWx
rBuT02oOkkL1nzBFYxqNjTbV5i+BcB30mEevNhBAWX7dfo+bfmkUXIT9pbjKkvNkMSNJB+io7rf3
cq3Dwe6Z8tyX4SSd/88d92gRboBDQlw+fTQRazvoIE7mbg2yZsZO5NLyRgGFAk7K+SrvBZwlWupU
LTEyY3Aljn/FTJMWJkP840kt7I7QEVUvquCCb0HFX/GAAIydj74W/cRxLrOrXxCGnQK1hVgnJodE
tjVumjEQ2QpOQcjufkKjlxCelbhCQKyCXDfWaZIR8LZFXcMj7ny68URUXUbw+wdoo6Ic0YQQDJYp
xvN0NWpJqU5RfimG53iBzy1PNNCELM3tGLUjcIbHNLpCHRWxRnfRsKu+W2SoegR1FA47I9lFhW0U
8YcNFRljWz94SIh/adixJAUnDlV6QCruVGhr149rSPoKvIK6rBsydh0SCwpA/qmiiKAdRiPqGpW0
tdMSTKL2AWCczFat17eGCIuDmElvmNlW14c2HB44uDNc0g0OlAIgsnrcaq1drBSCBy3f7YhsM1Kn
RC03XdIRMNAYuaRamnF2XAtGa4KeAmptnrX8cDSd20CuMysK4zB/iL3DLyniP9MjtHG6tEXOSP98
riQHdaL8RzG4uOxqsl/qf7ufrScvROT2Mxc9xP+kehoRG9AL5xsU6opzFOdqarQOCM8p8TTTdNu7
oqddbVSDbBZI2+zNlb5gVHQBwsa52uOyYDW5pWx0kt9SsJ6Cfo8MA2ufIC4VIKuwbYTp7WEQqlng
sp6GUfmVgAXpP8JV2Vol29ln48ZRLT53gyKGHrcCdTMlJwSvrZDJuFdblsuVOzEphGgqqfjbzReR
VvTffhkm8GhCsPPQPjV7e8kU7+NQ72P1e3R/HtFdW+mkP1i9TyDWuQE+9aOq2Z7/LxwmlvjwSa6V
W4FWrC2HQJFAxuwmewhile957It22M40OA/xr1tMpj1P3Y1HE+fXm2TITiyiN6DLlaWC+XL3v3pZ
nVlqZzgGEPjRUWxCKtcbWwYHA1H38sNLJIIt4hWe3ZfZs8WHL+z+gcltnfwClwfpTPOPMLMjeIkM
zyuvSPeK/5bqiSpexWETumPHxR5BZxkrFVA1/t1VCasDe//r7mN2gM41ufLK6tPFAFkDaVjman76
SWgHgcGLrxDDW/OoN4O33cPDSxmz13S8CPlfJEG9HuJK7sJ14dI1unxX01wX12X5GOsk8b519UWE
250TGkkoy2WQuZ6ylEa/3j7dEGxZDrXS+Z7uBck3J8rx0UatR+co0O9t7tLbujUQW7F+FeiyAI0s
NZXKAOt3Gs8QzqYH1VUbVO1X5hsrQMPQTSZ12LhcBuPXoAUy+pMmZnJkW2TL0gaU6Q4Osh8vT0H5
FzmdnYL+AaffqAouNwF5W8Su7hbp+LRmBGP+i+bvp7V0x+r7LlBUwu4kXUdn6Bwq+vPpa14hnFbv
5ClHtPt8Ok7caxq+Mr+dxyptTqq4rwOm013XSNj1i1Mla5k8OA/ZLNBNTT82ahp3oVnZvm58KpLV
OoBh/ZR3TQOyNIw06Fn5LkYblO4bEAkkPX2jZx3EOhkzEpj7Q/aIVLPkA3q6Hdv9pq9vGiNAWpzE
MJzWmaBcF4/p/4PCycFHTFYtxWInRJnCqIgkEdYApMWeQJ2j0+e5Y5WHgMwQtJZbjS+rQPpCb9N4
e11cm95gtXHOhxFzKQqLPj94wsAzoirEpfV28Ko6HtKbfk243S0acf9GoBAt5t6V9ZbQdmL7ulrL
7CdVuf1y8aQDCrFpbEZ5qh0cDOKzasRqUnaUK6DhCbMmP0A3rWTbJvqGKXjleLav/JFmU0JWtk1d
wZERpm8zc+w/MNku+yDWWEXyK8hCRB+a/tkB33F+NRjRb6A8CfoSZr+qNgRHz+L1Im2Q8PB0MoE8
x1kQEfdG3Tz1A8dBXT6CdF9HkwjSHf5FspBV8Kz5t9qH9Ocoetw6ZK+J271QWrxpPpFVBt/3/Y2y
r8QCWl+rverYGM4enu5un1yQMyZuKtQ6LUMBhvxgiahSF1AcfNCVPtQv4n6iWJK/Xwk6rnUftfWk
tJt7YAeluXQQHgtdfxnmBgetOXnsYW4uP59PW0aoDZOUcpS8PxuTFHSChJenIsGaFJrz7/+tfsjS
meIm4nawCR+RRC4kkfUrskSztUTiMFGUqOBZqdPoJilWhmidbUBBa7Pgb39LgGlTEjEAhSj7rgwP
AanA4lKlZLaHaoglkqf4YyCdS0UsZFxPjExvvKrJCVhwjlTnUoSsd6ZRMRMPUnw3t+SBNGm44Djm
FxJ8H8noyf3jOEWEDt0E1n7wPh605QudfB4r/o3xTOhd4kvdB8yr5sjuO76gdpadPC5zFS0NAeRJ
lyp6+uWy6u3GWKWvQ09KI4HsqKBHz2qCY5PRtoedL5OQrUPO36NhvYF9f1m0KKHJ7e+2yM27nTKM
5Wl/ku2X+gsYeKYoXNCSdr6cbPvfXcUr/51gxgB9rt/NeR27hXiQu0HJ0Xe0Ad16545aTRREEcZe
6bu4+rc29Qmr/HXcVo0yL+mRBercllxvTNl9TF2lhmK2+wtgxpQrxlOK8kXgLY3CRkrPub9kMMRI
SZmQezB7qNBh0/dHU/onECVFmhpXRnUGRLOcYcHRGxPaqO5akzCZenY5lbIV2hvL4ZP9DblQn9bO
2BzOOUc/vS1NK6OJCK1s5uNwAydfSah5YGTdRZVmT+BJunp1VvS+pPKtyDxkRWtHS7IqF/bR5XSt
uLMhK2EvZ0y+LH01kw74rq9hugzT4x+WNgJ4p+c0k36ooRMvTim0aPJy2vHei9sVlEB5Qkev1rm5
TGvAPXDmeG4s4rRJP6SIpbgycQZz9Be589qEVgC5+QZuBQ62g5hmWb/HxMd8K+B+r/M1KEGHh+qX
u+0VNzu3lYCmRSJY2yadLboNnF0v3A0P8/ylIp5/PzJs8C5VxbklrakwqWj38QZG1SAYZxnFl3EF
4it1aVkW5v6eKXMRul7tAkooFs1L3k4cZrqTICnmBs2zHMTZoinFvMBAI7s/e7ftvlMxxgZ3o68H
81UVPu0bQxfdML691xDr1wntJLebzpPy0u2waq1gTs2aCV06K1rLCZCu0sTGhF9L4CIHidywQGBd
Vr3m79cmujvBTSGEFaBvdestLDVeGINlJqpmZh+QQiGQpndLcMf6yv1qgQ+5A7ySHImExIKn9Boz
xDhMmdXnhg5G/pWBh5vDL+N86FB4ihp9FLSyBtRfCvRqMIVaC1mdbPlaiDhQNAh4BG5XT4LBBE14
2Vdt9GTXYdEsHNb8mNEN/JtG8LStFSyl+g9WAAkVCn7lHTx29YBuZ1MvaMglAaebHUzBRorPp00N
NVgvuJf4eleXhVhdY672FLH83MyvGFUbBf+Qn75TG8O8PMLY6Td7gdf0mygJfVodoPHpFQYY600w
MWB/mENzxN/cF+7DM+t82vKZCweo99mJ7cqcGfCFzYmDxUxDA/miTyekO95W+fzqB2T0q/oVx5Am
apHEhmq3zMQAtDRGjwYgtK1mKwmHBKAJyeAs1ME8OAW8n6ZldKc77I7xM2lt/IwMjScEeX1Dfd05
mrnaH2Z5u0v4rkEZh/w04vTExK3TNuDGYndzFYCrYuIPX4O69YobYBu6Cs7iMws+hzeGH8neO/X8
pOAdP5f8yJWWzS0+EhIQJSf127xEOH01Y10n/iuq8tEg5UZNE0OjFE/YuDsqOzV0lnvJ0xqV73Js
gBCAmDBe1qMf04ge2PyuxtPlnWl1q6K6LZnryE85Tty2PPsT57w6I3XOjyPAgaJedNfruCZPoCFa
6P02Sm09Dme0YMORymOvsGOy8hEyC3DrTciXfcB2AGOUFADBTLHjBLqFXfFd1yIx/CZ/htk+QlJ/
HN3wXCdWPJqA0t0n3LdH5XOEfZRuOH7H5IFVf8gKPIvEQj6lvzDUfWmb1z1g/9n8U/90mfe9l4lM
XSrhLETA9dJJHvEGy9E6JBKFyxvj5KiQgLtKhFUjD7oNyyROU4EZQZr6wvusC3dJPW/tzY+ZEhEG
HeID4jy9+2zZJtd3VYZRV7pIVCR1SkkCCsxjtX/JrQznXgKUfao84abU6+3qPshxlot/Nr8ttnfp
gsfCrFGl6AHqGbHu5XyI6Tzj45FSjJ9ik32t39aJO9RkfhQYXpWWWtLIcn3PvPwfFjdyS1m4aXhV
ezWfisaobB5ujwkNZdnenm6sgn49ATZgmP268HOr7ckdLSfAAIvGxm58QA/bxPQPWdJB2llBORh5
UJXxx4uQcMQF3ltW38eBzCkrnebEwZTWs2T2MJQ4MycVWlKIt2UMA21u6pqlpVeZCj3t+6g63Jtn
SwsbGh7aNs8uPG7S3d0kzZARr2USR/B8D0GVFAOtbhM8U/T2bX+u9/LieSnkViM57S3GqN2HxV+9
hH3E4LhJq0AuFdq92x1+Ueg+O1mABrjzUrKnEhy8nRs777oc8Yq/HvHEaDBe7pZ1kw00ZMmva53j
lZAW74GHX01x1rVvZoEPtHK+L0bPmQVtEqdxaMvHUhwP4ycbDRmkYKL4P5A9K2S4SvdKW92hJ/I5
hb+tv+AgVUbQEUZX71WdrFQjeiopa13fdK66swAgG8t1+ezcGItl12ZsOBaPry8dgashQPFBwg23
CvNnLQzheDLEdUKbnucC/tk63owpDa/K1JPKyhPgXoG6/gf9SDBDQqC1WWUZDCnSedIAleEuBUZi
RQ/uqaS4lCmC+zuae4uz6k67EC8rvGz2uq7IMk0MDpptXwAm0Gor6Fd0xHzWr3qYsIEJ8/bzFGnn
OO+7GQP+yqp6vwOKt5acyf18uzqkT2czP3c0BF0ghS6DNdwqIw4PtPhcIfA/LFBAkHxrsp8POMYk
Pe/QTe6/Nkx9n2hUesG6kP7O37bfiqzYLSkQ0K7jK2UUrq2rnGte2VpzkzVGPbBo759DHNS3brPe
cpyE8+woDAvxjoFBQTh0cYgH4JVmEaNxiNB300oK1AQtMJXfr5CrR1yMe6iFEOoZScwje3FbKxQ2
7py9eMlaAy5WHlcKQXOCstxdR7a0ZeFogPFBhKPtIv8elu8I0Fu44Ai1+epqjuHBSqkL39BcRREO
dmmTpsPmu+ANp/OIsukeGD4ia3lkmaXcZ+XNoi4akMXCVHFcb2JIqbXcHdOY3LlXOP7qESvU2PPE
jddjTEvqLotgwkZlm3+8tcIM8QK2LtG3UMiTRufDCXCRWQIngHc1K9gJiIdilL9BSAWWDKWCdxYp
1wHteOGA/qk5fIWQYPsi6IfLjJCHCNmaFwSqukwAeenZAwiDHZRj9R2qDoNjb8SXvJA0Jn+Qde4I
/exTK4pm/w6kesbvqS7MUJmqB9xjc5pPMjXUZRvIqRhgDqldDx9qoRX+fbqlYA3VpSDrTIwbbDhI
2LENF934kbrRKRX4K1XiqOl40nkVJB5YDiYl5j0D6YPUTAE8W4o3+t4o8sOr5k3BPJHETd6omHXj
7ZFAm1gAcy7FNnuM6c7evToZMLFIN++2iD9YHL5RLIx8OBsXJl01pa0cxkU0aoDZGqp7trjRvcFh
q6dTyVRsgJtNpBLi5E15TuYSfEWajfG8pQ7mYlArCjAc8Q33emD/90Fe9SjazKbBLlQ7CxMmfUc7
O57qfya/QhVZ/e8n2BGcSdhYqnVJ2vPjCtKZJvWO7j4ueOpwfUVMmy37iIn1FvZZViUhwcHydK8F
2gF3l6MVGs1nm+NibaBVwbWYe+lMAA2yKte3wLOjONxD/hED9kW9WeqZYuUJIRnaPuxCm14s4vIL
Vq05MUiWRRWV28+9y5aVvvSCg9FkcpM+m5iHz26JRStzG7x5DnDCwY7mCGUSOBbdIwRNpcKC6GVU
pIuhgbhzIeNKzK5DtP6LTFihMDYIGaOIbbABmEbOIzeqloxjdygBqV7CTtR6oiEhMQFL8YFaSMNv
jl09Nosb8/OxgsCwDPJwz1zCmWceLuGivqN0rwmzLOVoJmztDxyW/Kx0aN5lmDCOgF26ekPLqp30
Lviz/2ehT8Q1+20d8BuyUNy6KtOTV0QN70fDgft3osK8DbzyGSYBVYUSm9hnMs7J16yPDuJFg8xU
vhwsdDYT5gekuBzKfk3AmgRuFWYWTybzvEQUa1gHIA5i/E6ACTGVa5pBMyEjUhwjZFR+67UD+C7P
8LaLQNAMQBL+pGo0QJcEpUJzAttIv8YVKDwSB/K+cpgDAZ8ixmdhedZkiG7dUmCFnU7d1Ub+fcE4
USvQcBI+kXRgUL+Mj7pQ9r4Ebz9J3L+fzcnS3UTiAAKUhUYfrRuPtk56wTZbuZScwBZL4wzRyh7V
3uKpkXtaSNL7FJG0wcJ1He/nqFn6n7kdCOBgzwfwD8cWGg==
`protect end_protected

