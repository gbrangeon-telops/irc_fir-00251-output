

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
jPOKnt2dHOagW4dFov86UptHPGMdrE6d2ZgqMnfJehhzqeTiVLl89did3kf45SSrRMnQy9YGjxY6
jqpfslmzag==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
TbXlwhQ0d0UG8+CBDSNOnRgRBfh1oNNVi5QwoMGV3zJAlkTsnTywwNiy3IArHTxG6Niq+d59upyT
QOuldsHqtyc6KQBpxueCYJG7Fv1OIOGGq8mGjrkLmbJVhJEwBvPv4mlhsXKQ+/UhmQDpF2ZyKhkK
EbgpRIm7ap2EmEdPduA=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
iaTK7nKuH82rPJSrGYALVeHLyxEbb+9Rh0wJiyQuCqzY3/f+ne/dT7ytF39Hm0BXD9csWKwQp3QC
vOqzo1FyLi+w9Ik3lkb4njvMdZauHueYbVoku659dslyFGV84Aivwjcg0Y5de7FqsEonjWrVPTE4
0oo4m4QHuK8VN0pa+LmuzTIHDEzIPM6IMp8H0IstAk4VaGHg6wlCrG0u2kbbhcyaOKk2xzxiDfSu
gcUy11TT1zHFME/fHUU4VO3aHMSGacP3N+kgMah6x7bBUjBd2rfEXkVcl+/1g+qp0xW2BzItYrMY
Q1wtoE+N2GipiyxU+AmrXQ4zQNqO11zaj/N6Ig==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
QkbQ08NIPb90+bNjwXDlVNk6WbvhfydYhJZqryulAczmjZMBvdwitIPmanwzKj9BPStsPNHXyOKf
9PFA9l/uvQOwVNRTz3G2U0+6+YFy3j+qj97mRopffETTpncxm/BoroKpRNN1DrgSjygcTkfrt06N
1lOXW+551KWRUPA+fGE=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
LXGnS/C7HF/SjGcWlSWMUKmilNZr5UhJNWaaWr/ybus0u0ctzmNkXcydCyfmEQe8OngFPF/IKSaG
XMrlZODcxs6BdW6TBJGvkBlKfbvIYg7iCmAit8JvgZpuYsROJrZ/IapJ9XCUZT5PW0Y/S/PoGs0O
fXalNP4hoIYlP5OYjMaSowkFFmCMq49fHUdBBmi6thqlMFhrdpbAhfGoJVYkjStWry+O4YcFvpKw
Q8WXsOAh5J64eppUG0x86EZ8HpsK6EGAeT39tAy+jNSSIcnklat3mhXxMF+BE67OS/DRt5H346yK
YrLlKC5qbVgH7HjzWMBFYeVVtUec0iic45xLPw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 11232)
`protect data_block
aRroxph5zdgdlg3Xxz4Cr4s7rtzEKj0jHKFBZ5lRck2S1MwoTcATsR0/PRIiyJa7cpKaVt/dLvi8
aPLwl7YVOZCPrWG893itnNmKSNRAfhhomZl/OQYEsysNSMhuThSe+7xHJzaPO3atlSUY0uwIxZi3
+sN9BfgsQ8ijZ0Z5AIaNwlc7GWydhh44WL7lJsrloTz1bmvJLk5ld5ISht5TVSgt2odln4q+s7TX
H52zz2EbVuVwHLobheJ6ZkjVSNSXzP+pidLN4/1n6p7tKM7idwJJLHoVCQIYWtFrHQjqkzHqI/rk
4UHwFi5I0RTWlhrn+7tywyb6gq4EFDofDIih+BOY88uv35Ue2n6BqRfvBfg53BkaSqyZ1kWMQWDp
ssBQDvXhfoAj7DzmZf/sW0TT5AdT97DZQ9CzA1U4Bfq2ZBoz5szS6OveKOtWhmsnUo6SZ52crjxC
6mTWe6cVDk2Qlo0UnyYtv607Zv0R1Ly9AoovFPEPLNPtWvidChn2nWmc/ql2DXUIDLdYa6zlyr2u
vfi5WPpoXyuhnZduC0zPsIvkZX6PLFB0kCgxgBtOSJ1P+W1v/7MXMMiEMTf5j2/bBoYkokFQBFEd
MwwU/bbDrX3qRiiOO4dsOAjngAGA1RQrmEV5qkcEksVqGjLPsNgEhTSOoeuQaAq/WErlo6lr57wT
2joWFDVgi+ZLZoy7x0u9XsXFSommnYs2/J/vARELtLGNL5WvMy+GpsOTWRll/wwlWaBjqsjp5szq
LeCz4NNUl5Rc+Q0c8tPYnEoOk4MS+vwMgRRe6sQ+nPfafOgdO1WjWjEgvISgPTpIkfdB0zxkIkre
GQq2ZeBUx1Miz8TjCwvmGoznQ8z1IhrtSmfmzKG2z7DO+SwLG02P3biYSYwazuoaRzw8yZskcZ00
9EFXie8DWkL7QSJJtnurHL27Cq/nxNtz4+MKqFdYa4fkb7jZ52jXmvL1yxm/j2Yr6JdJ56vJpoEf
3uiqbo8ub6L+fISlMkxQiWDAv5vyUrnmQ6+ZXa50REwh11mqtWj9fhbuNt4SwWS9Ci5re0Hir7Sx
2jMlhf+QtZx+ZtEMsxBqeBP5ECNwkyvCCXdj9LKBmwbO5OYIgktuIL7/s066Ly4b/rqw0L+3YPDo
hQAAOY37MpbOWdpustPrAhH7uhcq6H8CMPFXYsuoPA0Y5/rdT7VHHzYjHEXf2iO2dqhC5daur4Y0
FH3gjU/xfwFuOfV4myu0nRKnH3e9hWjLoRLeKGQQW7drstfYGKO97IZQxtrN9XwQ9nGSSHKTAnh7
JVF1VQShvGWi4n3q4MCrVu9EVER+mnY0VZXHpOpj4dN3NaKIjHMaHDG/6igYvoC/70U/0mJNZWOT
HVaydLygIjz2g+vMOm63YZ0WEeoZBv7wDcjcnuwzJ9t7IXw2UM2pQpzSHAlLIEjYldYvmY7b7JMD
6k5+Im1tzHA6Z2f4p6B0gL7in8jn+/T83te20mxlzugvwIbLM0AJnzoCIeuEH0GUrI5U7dGaxVZA
pJcIQF3UNaSUziB07yeTmR/wBZQ+m89p7bhdO0qDYG3bXhpbR7xWi+kZ7JcbAK5/J7GnrlhC7RzS
5YpqMFNng3zsBBHSZlrcqnFZ3KGlbkMFa6bLUYwxjbPed6scl9iNHWBlwH7T2Yld1ri4Na/bGBgr
6DyDRtF0Zm1A1GsvuvxdmWUtnoP0FyAUCfa0eJrmBrxG/Mk1wbADkJq30kOZPxTjzJyLu/bUlo60
TFLty8ocl4MCQZETAM6PAe05/gXHOLWusohD8aeQMEBHEQ7SYFHLXXroZG8L94/lVhjcbuAu9Cui
5wVg3eT3RYJZWY1FUv1nmLsWqi41QbQl1TjGl8houYhjuKF5e2eMhavJXf/5+codc1AzHnKZKrr8
N9kW6h1Pn6qJMolZkTtSsisHVSMyyfrCqtaKKjFFP7XW4UioNCudNsKtG7NFi8E/+31dcAEKj0LM
GV6EYghkm4vXnrlUx/4oHa4TMj3Tj326z92PSVExcf7fJ5mgiZFSvoKNPDAa0Pt3OacEd6UGzh0a
+mYXUyJFVFETuenpnUhJ9kaTRai6wPl65BEqZrH1wgz1uRmy91PbuKQVVl/adKAA5OP24L+/9TjJ
GTuis0BAMGaGs6uvsZ3+/+1XtUxk2U7QdSi3UUKkfNI3tm7IEtm+XH5yELwGVONKqUyuwjdsuus7
oCX/cUbrxSes9WpL0WhXPNDYCHQ/M/l9meH4GvMzpPOUu45XGFqVYx/9uomMFPVbwm/QF0d8NDmm
8+nKptleBXMwVaaC7oXajvTJ19vGkk1TzMlvq7DUbCUtHm70fGdbi9Eh23klKklJSQXVnkTOtWKR
L4/UbspJMYfyqFiH2KjBTVkUtCB7CAdJq4M+HjOx4GLlg0lKldzegD0w9oZOlQIonjzJ78ZYlu0Q
QILC3HcbKkpGESaFWz+J31ZPlQtjlmOPYxcKupb6Tue2t2KODiMNcmAdrnHERcNRQerrwhLNZVDZ
9eEXffqRG8qxpa98AX1Aj07OBVnISaA5jhH9KIF81Dr8RVwjkbs9KA+OS6C2ZLPwrwNe468zDyTt
OTWV0hATg6whSmFXYC84tv1w+pPqQ56F4o2W1oWWVUIWjKb8Arl2V3+P86tvl1qHeNaeNhc44eeY
m8eWxa6ZMPbV/CyZYm8MvU2viT5WYWoevVplKLkBLUnrfkMO5DvaMYltVzjafB93WQTuEOAnJ0xv
1pzReHF3i/NFPgqOoGAWEi/cW3ZPWtneV+LB2TZV8kkyIg+S2Mqh4dbxCAbYC+6vbP6G96ckwIoC
yx+vlFEiTEuFOh13uLBEDYPHH7Gu8/csohG7ZC4PjowClWnWn4pLlvyDDle9wTpCtDwT+knJ+VHg
InLH3TudxIoCwYjSsuvukol77xNwfg0o75Fq3OhWQYl1JnlGOzvB3a+f8TFmSjCumet2bPCEdkWH
42p+Bf4Vb125DIoCQTH5IwqB/0ai1m4/Ru8dTBcIirO+Ql64sv8A87uYpbjln5iiPSa0/tQ7tIYF
RkNfXUkl9N1oby+ZokoDVzWIM+zqbU+BGdvY2Bs1CLmbVsCJG5kgqPR6/7D6daN8eG65MUwPYNkI
bxEtkyLy7PtxXODBNZwhhHBhdd5MaTk6PjJCqyga3I5KocqtP/v2gUi+77P/gqQfMxPdINlIdqno
VnWRtQK2IiDEpHPTAuYs8Oa9V7BVdVr/tvuGd8Jzq0Dgot7rn7QgTrb7HmrFGvnWBMVbPG7y5iEA
4axxdwMvI2ePyHts3IaliqE9IF9A5hfP/crOeVYUhGhby9DkJKNxKyx0GgsLc4d1oBgIsnK0teKV
y08Ky2JIMKgeXikVqXOtLgbQLqKuqoxDcjVpjZu01CbjoIPtZGF3SXhttqTTxq0jbgis8P1BQmTJ
26uSaL8NHhZLpEN2htYrr7vfbwd0Svu0GDCvzgbPp9/wIepGBM4CSYEzAKIGZQxv22ZXuYwPT+r9
lzIwhMu+yRD9sEtKh+ZnNcz3carBHBfVP0hjgohGmdF5DMurIMrtiyjJN63oxSmSUv5IAwPlKiY/
g2jZdG9dv3NyJczPkpx3qkaPi4nIywApKCtsBX1P6fT9FJpGv7ffBHNei5HNnhLNEYzvIUSQ1B26
zVQZxjZ7HYKOXbIOfzjK6KxSiFsynI76oiP9AXGAla5dRffmbdWaog2dLirTxZYqY/YBLwxfg5xr
9T5b/e7wYVOtY1WVEww5/A2lSKLKvp97+uyMQIm6lHYgmfCMKKCd7gJgliz0EgGQVcMRAGr+j6ge
/Vp3GQTqBSRjHE1xu9P9KbOTgKszC0rARSXaS5AjDxuOZrmmiqL9I7G8GdYTNLg0VAiDSrM4i0pv
1WbAw3mfaXAbOdbKAtMDlaPUPEC97Ew+JgXXw13yZvVBD9JAFVifOJ8CNI+vihbDeHz29EgDIsl6
mysbU3OrjoKa0gYX5oNskQ232k1SLBWWOkTZY3y9aDb55rF3zit5AK9ISQK21K6Yi2cT2knP81b2
36YDhblJ0QubZ3IxBstMDO56YkIMa/lR8TOPxg1ezsHyO2khc5Lx53meocS6wJJ0CvbJnwR14ZFW
mkG5Kzb3ycHk9FwWL2NXuBPgq4pVe0hBhwj24PFd8jrKunghg53Tq4M9lXarAAFCUbRp2BtH1Q2O
42ATeCNnCIfKq7LHpSgOWPP3Hdmh1i5IZNbjB/DdGYBosFAmRXAOymaHdkEGmjJhsXqd3e7uDxTE
XW6ok0BpqKPlCYsC0D6Ijo+XLjcd7WEgFsRCTKLD3adOIXpxEV242QL6H/vsMhOrXj/bDqmqJ1vO
fOGEwdaNBNEblzkEZGyTA6mx/vu8rEVAfO7NNZ8fBFhVD9pTiiEXhs3QAgYOD/b46meGu3lnf1JO
JrPXj9+lLTkkcFW3qmm0sE5Dyg72iS0pRzfROKzzLOioE7G95pZzdAmgwSVhl2WkTMNJJF1KCTFd
a/Zl7MShpAQak7p0llaV2BtIDQ5qKWdvz2Mg89+eupJ1jrMs+UTTfYE7sseIh5D0100l4S4AnpZM
Yfcbsjgaa23F7VCyYweIfDof2AMm1w/N1dkyxShfu9SMCRJIiWfP2nVqrUaZHvSP3pgBMWGKqnZX
mXHq4bMSP03LcPKirWQksfxyeDYRcsoZM2g5PYUHjY4PElwKKJ5vN9JbeYuMH+KCoBgk/hdXNq8I
OOaRlGEArGfYPKd9WFboxmBzfQ2nxT7meDLseLc9rI9F5eYEJKhwxSc0DlIM4FFFnmUHxpc7G4pt
1HWHpyIkEnkaftlUe3idp87nWQg/bZ5zHssIt/3LOrjNw2WJTDX9yEPEcEW0qjXWjs7LDql4gKTF
J2KHMtvK5oWF+tYXZXiBZITKPYi62eeJKf4fnAlZlPJcrJ6Fev9DXyIIn2DSf9RYkD/BYYL9beYT
Eub7/tQg7h4YdkGVQ6T0KmzEpKpq65djvy7PWjkA8ebO46mZBDhhMqZyKET5gqy9xOZx/Vcn8qCE
AowEUS3WLgr/csCI1cV4uSgfWhpQQURexewR28uSgrPr0qR/jfrOckZ07U5bCklKliYWDIzBUAgG
Cpy9dVOmxS7ijFkUT9qodCdrF/aCkL8BAQ74bHG3925Nj5Hu5edQaWbS1pRMjJKmFjjxUHZjZcBj
DH+91OdTWerxWc0QWJfLPMiWtH5FH9+guxMjpPia4UTGpcAGrrGUG1mc8yKABnl3+EHb8XXj17C7
ED8lPfa5k5DOkFDzWH4PWZCf8Sb80dHJBCeMwqTI76mnbWHAeC9pEheu+JHc16Wc7/mYDP5I0LNV
JpuIQIeTUpt41YlsIN9DuRXpfJlCRvSfgk8KbqmeKw5c90Y5phgTtowXJMv7a6qYeSB12WCfkWqk
5xTFn797VTL9FELBId+q0oIKVHVd+WJ4Et35BsgbYGn1ahdjqSUvrufEL6sZInIwvNB2z2tshrsY
x2ScAdfG2Ts4UGYxoTifr3eV6N2mvnZ+1L1tzh8j8Pm4uIfuCg3tmTaVJoRch8JtgrmTcKLkwkwF
pJSZkZD3XXN7+dEBXHJ5oMH3j6EOnCaiKCGSAlMyZ2gZhzsw30OqMp3djQq3SN9mhllCGznd/6yo
KscUNyrQVxlpQaAchNQNPMKaBaQr5QmlmwYW1OcRwfGY5bUJ0/pt1d/Rmj8EcVbubY5oUyf+mWQQ
l/DucBET5ihU49mf/YWGTZNJ7b1+i77KrphXqH+TwPAyGukwOLED4LxPOL9v96flWRQD2AsyKdsi
hNgr7kiPjrLUSx3YSNLr4geAvamM2OvjhcghOwI3U9Rck9umV7nVR6aErJ949dSxkKDALB2sgUFc
F8xF9zclWGHJeE8zL1KBq+cLrSbh+N7eJ/LBQqq7GZpgGhJ6aBNFmTU/FgHNSG4TTvWrjPZqPm78
P27arogGFwK1APmKi3Ahrzx3Q40GA6VXNJ0wx2TBhYFhnazBLuw0thWm9Tek1/WlrSNatODum4VB
tffkZQviQgTU6NUUzXd020dPLZcq+pT8w/U/g8a0CGEj5u/ZZmGC8drFKhuAsWECvv3o3ZvP1XLB
GAxn5NWaQrjJ1v1pTpw9smQS6RrHbffPgBvlXnr3OuhfDvT2Vn4gQQL6QEecbSR8aHDoHCSSWdPZ
W3XVwAAPAJHgs/yeaR8mcrc1IbrnZCSrxApXAaFCFwUCKbN4POVca/gR45Rh/k/pu3JgTSB0FWo4
bueU1zIVUknOIfkEX0UiJAUQRMP8Dh/48eLMQS2vzIF/stoRC+2wT+R6kjbcAjGE5pOv+isHNE/0
QolnCF9Op7YNDY6STj6AuPXmw6hLwb4kCpRcUQsxXCSrDeSft2RmfBN9Bmg3vevLhjPkKbo+Putv
QQYhUvH0dwncoz69mw3qhBt+gjikuipz+1eKksm46DGfpIdA9IPJLEyUEPVEbnxSMpm+/M+lRuQu
+xCqTl1l93YKMsHdRagQ0Q92If835KkUgkSL9/MSFKHuD7cE6Qa2yGpoKlYDPT1gfrxg5yb8fUGP
o8X/gmt2XqHrDRTmuTZEiN+eoNcqHDOAoCfL1gA7brW4uQ+vY8iF7lvSjCOdGY+LYclMl1tXW4d7
n6NgbDfVUXlUx3qcQyonvvcEoHWexs/hqPQ/OcxR+oRe4SpEgCsCci/TiitV25cS5yhV4RrF4nAv
tQ8+rSeg64hAUewVWvw/QiGkrAmrm1ggLp4a2+IdoQgg/vHTtApFGFbyTqEEr57EkPws4cC2sBgd
zyzXsVH2DnjlDg7jrJAs3rFeWbES4JWZjrcZTAI4eWT0eLSN6wCeUDLB+rTdvXvXzrumjTM7j0po
oK/ILuYOBKtqDEeyZh+uPT7t4lREdKCIwyKT0OMAacZIHkiJ5/7ADPitpN6ajnbB8On5sQljW8t9
g3j4QK4JDfU2EEwf3ZXGizCXbkSW+eW3rDbik9psoZ6LVMx1UVQ6h70XKS0Rc3MaOHXbWh39QioE
VarXk9tdRMekd5PjjmeVkYOxbcMTwTOcGrmTIyMoJdW4kUMZbeDp9unzuV0amLNbvc7sxmw+0qOC
BBL/CGIUnCc0udQvbQX3PuksyBBkWAN8NQdyreqk9oXN3qg9PU1+yl9LLbE13pn3dNiPNdtLXL6E
JxYIXnJ0exPrB3KhCxvV6u+Da+edD1uzj4ocfuGMowVHaOJAUDQBT33tmwsVD3ne3k2A5PSlQFyA
zCJ+1fxqarW9zGic5dhmV9MjtTRrJrgIWeFtgS8PDL42/xHEY2PNHcvkhjW5AL30J7RAkvi4qAQy
IvqS6gjiX2DVm2xVCsSPZAB4GnLWxsn0tPJR9zIipiKuv37WTm1npmXEh5UGiotyb1P413O8BjhM
+Z5qZcTWAk8kSqmz9yIlH77VBl98p4KO8uPdifjWND7ujNK1y1jp2joqqTwsrKSq+4GTEkUGC1UA
RVjqRdtsz1Umxmws3pJUnR0sBJMgXY8oT0R15yutbAsT9KjS9FlQOqF0AFBI8hL8qmut9G4cSfLt
ijHXGElFQH48ZddwW2+BnOLLDHweFsCslMK9zRTSVtYtnv/lcrkHYsFf5G1YncaDlAwHwyMklWE0
l3zxwtQdXgUmjhzxvgJfZAFKtUZSIHrV7K0NBy3TtwDn83rAaK9ErVnruUvrTRDjFVXln7FezOl5
ge/vMm3NO3CnkWCUGI+6y3dJFk3Nk+O4Nf8Uezd4SXjD46+2lAIoq7WZyzJFi0iBbxqSqcJIY6OO
G6DynOCtmHVx/tE/K3NzgxSPe1+mJF/7UlhuYSUvn1LuFqTn6M+x48uNRI/AWNIpumdkCbeN7Yuc
JcMUGgEjps2d6T6SeymwLUQNGJFlJVdtfRDFQJ40wn3KeVJW+dtSUFYHmB7jSD+afxl9i8ffzNTV
ibU/sYnoRf3/JtG+b/kVscO000SyAejWDvs7dwnfVMneC8h2wyaRuUy4POQdVBmHgiFIM5kHPtDT
c0VEY30mbK/KvUImelh2xEzeZq8kju1WaKNvoTpMpTcwdbk5MO1N23Ub+F1hBP6zfWldXc0nSbkw
mkpf3WtdExfZIhM1J6Aa1VJ19tjiebUjM023ag3i/WDwz7rcg4HIbURQcpqh20paMBGmimmKTWE1
hNmd5fpK/QzTWhG4TidOrEAdwUL3PkRMS0zGL3oeKojNjYYv8fnNLtYfBi7oswLwFp956NHcaxFP
eGMnMkx5zXITjYswvaj24pZ52Gf/5QUQq7CM9U/Lm85QVIxnZVuuJ3AvEZD6TxOqfAL62eFqWLl6
wL9jcqGJJ+Ih1Z3q3hQ1zUWOk91iBP4iEzVkLVXkoNHw2ax5fcbVCG0f/3D4dCyNlKfJSBW4TGff
UNYf/np9VW4TldoFTHZZZZAUnKEnIUYd7Zk1So7dRGgHgZ7JQGTtiG29QWlElylhTLNM+yaTeL0S
muTL4UnqdczYki+iCb+xAVf1esMa4zovk3Vc59GNsVY9oFoJx6lzExGAmv00ORc9mFVPe8IUflQG
eK0VpH4Y/P8Nhsn4RoQtrQ50Ca4P0axvqKsa0lotENe0Yux50xt7rgMYJFaIeAj+AObpaAgmP3b8
82KUKMfkiB9zaQuJuH1FeTi1Vm2wspTSB9DSz9FjG4IL/dj0ClIgJt4amMJrlnhuz1+Ac6tjwK06
6sMu1uymWArYx4iFM/QqkfOVOI+qK6TCozA+zylyADLTZK9uu5x83I7pG2q4v1koxT8DnK40EVm1
LbU4+G+CUbqtbynEqtSaQRBoLtq4p0TlldkZ4ro8SNpqJEHckiPYUl0BTCt391bWaq6mz2pCXckH
RN3e8Q4+KukeSbsYxDFREg0sqkNk22p3ICrwmK8fMjIuxOHZB9/aTZJJ8N4NsCU5XTMWXm6FIhSg
mAjswLyhr9WYRP44Tr2baY9KmZRNEZ/QPWvxotWzLmL8L0r22GiGpJX3nPqmVAwKV+5SKM4XlVaf
xA62YZRzE45GMQwPOEmJ+34KavDm5Z0pcobhjHbbra+4+JoPwS8hNK3TJo8T9DXxsR4aebcDg+Kq
LeY6fRQZHzugSeZ8ptej9zR6V5hmzcQoEKEyhGyxO6YvxZ5ap2s6pnF0tu1nkltluVA6i+hDMvET
lIWSduJRzM5S0ANp53rgoEI/+AVRV4569FOUIYaXA7LgVfABz/1UuZjCjjeNY5HU4PbgVZjzidyG
UzrlFjkBP/X1k3XKnxt3+is3ew2AePgDkBG/Fe/Ls+kJCQzgOE8JdLm7Jp5ZyG6xBk4VTbTcmIww
kFxW6ygv29B8dWojE/H832NQ8TleSLTHYJQY6oQTPvqKxSCD7Nj7GBgJ/fDyZIp+ifUKBEi3atrN
osLnWlb9+7DPB/X3BRdpZi56MYRMaWOe/ZRVImnUl0GEccCusAOWUQvyiVJaKG1LoHf+GaUZDYKj
ThOJFp6aD+UYtHhdgyuf/nSgGy780xtfI+ZeHEA6dsYcEgKAw2Rm7D+aAheQxbAcf0YAhXnSjq9A
fh36QGUbv3hXq++IfEZ9AV2SzqVT/pNOFf1tlzy2bzffVhATkxgdC9zSESiFpCgrd9/2JQ07oGjo
vXFSEfrAN+YhLh+5o29/460ICo8DAe1lHjWnCGuZBHFIvh29Xu0D2CrzlufFlS2Z4mSNWCT/SuKA
Xzihj2TqG+lXwOMi9kRyoImQLAXuFKC8vAtlR+LL4e6TKEtxTtV495hmY+Mp+A5ngoa6ZjjIbr+l
CBT/6vvrTCfQA9RaLMdrhHM8k4hH8mLLTQT5h3b+t1qLmgJibGIv3PatiyriD0SnQGqY9RKTUkNV
EIIv+qlqc/TA96M8sYag5AJj/GmKSYbMPtDp9H5SeE3Te5OyIhJvklAkkh/BPCOLpsSapIoGUAFU
mihObCD6r+BkIjAOv3GJ98fa3a8NXAG8guOD/Id6CCDtlSpe1jhie6ETBCCPdt/zc4GK/PIubVOQ
rAdQNpWF6NGpzBUYvVrQwI9qJAZz0pvEQWtriSlYpLElkmBHlLRg6S1CWVdKBmQGhxXZE5mzDTBB
oqdPKp64oH63GvJOdSITPd+wuUu4Wke1em3I4OEwSoVrIuu7PNELVghwuEbg6zb6ldVcMJiPgEkf
fL5Hg/oiLJM7BNp/iBjwZzxS6C6/TDmPiQSSQdfbCR7yXnbmLV09EOYlezRrDhwYqeqd9t9ebXeP
coeVWf62wrCGVNsPHlDrESmr+yD6tf90bPdY5xTBWdWl3Qr1AInKB5U/PnzqzTtz88JjAdyGKoc8
OBohs8kJ7es1zjqHP9081glL7Yqx39jdnSGQHK3GIhYfBNZ11vJe0M4g2m6QeDpLa/6HVeU+Mx21
UJyrb7y3NzBtSVjmkKC2h1bedSKt0Y1Uwx4pSCX0tmffDAcwYFIEsiq2sfaWjO7RVWUQSMPdzTBE
UD4xUNENKN4JLz+MqE25AIWHZwCni8TLG6PJOWtoLld2HwSEgSGQFvjQPq3GqjqAnD/QeyQQGH9X
5ZF22PKzisnQsXDA8IZmkX6foCV5u8LCnbSgADvgvp3YXyNpbLidp93Fijb4oyN52ptoFQ5yMD3q
IHUJowTsGuZWKzKacdyB/3v6csXlzl9HpJnZd2PgEKNCq+n+ywE2vyPnIlB+KnRc6NZGSn7vB/mY
ZCzaut0W7BacbrsO25Q9vyWC11b6vxKhSy3gT+/cI9cf4ZKRFG/lTBj/YPcUlYC8WJ/bu3YabV62
LKfuoi8ozqJtjzEHH/iVlqKqX/tzkl4h+1T6m+7SexQbK61Md3P+t0jkhloOxih4VJ+lw6k4B8ii
v26tXzZ59shn5XWJz+nY2jEQpbDgv5xcEbm8RcYzMNR7fUMZ8O/kbC1NcW+6LUr1SGPOREfJLctU
q2RcW/PRR0td3nj2/TQt5/nMMyjiyb+LN9e3p/e0pHHh8rTosdWKt9RGHF2SgADyWLqoVHJHXPw8
slaouUF9GknlE1xeP8vha5LX5BSwXyBobeeDOrpE0djPj54WsDzXA3ibkcqNPKLf0y1f5oj4rDE+
OvQDE2L42AWVmEAnf1NXtN//DsSU5lEx2uXkveXdqa1kycods6SogfUzSe0nEGd/JagJBcSuxxwi
oht45PQ98mdjP3f099UoW3fqp4uN/YAGS9yx1cWYE1VzSTVgERwZbcw7P/Jq+y5QbzJkIhyI48rt
+997z7YySeWF4VO5028RYL1b6PleG6biEmO8wI9Sad/n4JabZ8QUKQk4pbhyMFbOHnupbUEJgm6T
02IJrTA0i4LAooPVm1f+wj3J7jBZLvO7jWuolVfRflk7Sognpgxf1sl8PNbInU/9jDZwG+PbpJYz
wI33WR6N3DNG+/t5BaQtjXmsW9uwIc8UYMMqfD51zjpAuE5ISXXVOsLx1IxL9mCSc+KoRE5KWr60
adwyNNLFeqvKY7pkhQBhDK70YVmMJEzzXH3r6Bg7flnyraCXjOx+MIuqeeQDGBydILdCGkVHsXS0
LkDGOglSfS0Pao+NbyflJtK1bIUGDxC4bgf9ZtHoSb3yQCKOoJkuG0cm+YZfI65z8Glgyn2ogrJb
sGzfV2xvAgjnJ7SIPGX/WZ9klpLtc/1cmStn8lZXvrk1XlGh+YIvPEkJa0c1UE/3TZM8hjhzTwf6
J7bSTITFYOAelPnjlNwxV0I16y3E9vlzca6DGDw9tzqE3mXJj2U7B71ZckQIUw8t1+OAZKJu+Dhw
OXVrDmIQXJcNaoODfgdzdvYTPVt1Emd6Pb/+3cLTFAgHLxf/YdOAU8IeANUsdXJ8kkSkHzpNs5HY
1XmUjKCUThSM/Ep59jr5gWMUJcqe2t1gcKJbR2qSI9npTynMe/tYO+rCHvhmw4aTQQf52sDhKJEI
1mKYZevn14U4rdePJnQ3a1a28VW2r3xxBJdwYVi9SAry1kmAhq5x9OLkr0pDPhVXSez4fewXYPH1
b946qVhgaVBUXuym13R/6mtqg3E5QoReT2ggWDM3rHROkADswKkkejZhdaNBqbnVLPPrx0dl/IqM
BBiV1d33pLoCAmHv6tgu9mWYy8JlWO/j7gZwW2swZEP8qVz890wJYZVp9z30RxJLSUdKwlTfHpoh
txPCb8BjUWJrFLdCWilmXxCpUtW8jtembUEuWf7ynR91Kx3zdfzlR2rFLEUrWzNqPL6sKbEXyCQ6
k+VvftIuLiSfWbMk36pnipcUBnfvj7aReTHTviO8OycqT4aIHq6uUo91wdkKlqf8I+u+nJlzOHMK
okeIaRMJ8OTQtG/ducOazxdRKstuAHcN/DBApzcGlmlHJolzWqs1am0mUY8l4W6XgeoKf6B/h8I4
wndTV9ATTBj4qcv3OH95nuuVG6aJKWytrri4CcpHEcjnyvdTyRlUINx6jgJoAozUBL5SPUQ7U/59
ul5ruDMnh+A58P0UEDGCnWCHRKz+woqPD8YXHhrKYHpDv16FjAmWMO8LL8h6G370QzyiuYFeWfsY
NEuX98sJuDX3xO8YpE26C8ZoFWCAOWgybiTmFZQbs1z5LpV+PkC0GaTwfeuudFXKS17oktanwb3O
w5p65O0by6izvcgE/9F+vyEkMnTUzbxbwP24LuC5q9i4OsxtykMBNC93Mi9IHBOr5ruS+eXxgO+1
WNk+CF9++WKbO5gWd2gg0UoTZwc51EHs9Rl9DKOGWgnoiPLLFfPahaF8AFv9+qO7j4m98a2C9ADD
o0mpeE3Ar5QdtnoQb+ccEQxMPdfnvSJ2OJ8/zCQatAee3+tQirb8nGHjYhvS7VtCFxEe7yoKs9th
bEB3JaptOulJZkzgQZEQoHug6bUqqpBDv29TgTqSdQO/huoOc0v/01uMAIevEknLUijmtZmR5lv5
737uuNcqlHDFczD7ILGTpt+tyvooaFlmO9R8MUVEUITHl63PGjqXTEXzVcdP18MAeo03SzdkvvgC
/IXm9Pr8oYn9aDvsJO1qMp0gzaDNr9mLlmnVOy9X0nozcmnJaW+YixOy+rCkg70Nk7c8yCJMwh+s
arYfrAMRyybkUgHcB9+pmWjtcx/KWWUJ4x37+EqoxH/G5TJ1Xamw0JsoLPgZP1Jxh8iQgAQKErMR
KGNlB8RgKaAS5rJ7OPHpADnKWLE9n6fhqF8fPfU9sfOoaTmfKtvrrEdGcQhiT6mrs6AN0wiSoCci
8++raXZIpbUR5EnSq0OK5JH6Oj4h+71H2twRhJ5jcDZu3JOpPXVc6Azbxr19WVuUnNGIlLQuPtf1
UZGHqceu1NQXnEI+fSyc4t409qfZgd3F7m9pUlkgRMYOVx39xXVw2rSRd/HLTZgZ6EYQl/rV/5iw
WX9jK3a0hb9/h01k/IOFTsTI/NHupxt/u8y36GI4S0fA7G0m3wGeg1tVxrmEm2D0flwUcI/01F2g
J0+XUG0jElhiF9lDZ93PxPjhIgLVv8DCf+j4mqG2QATNdb+0lRojYGOPr+qhvs7vbWwP184vpuWn
IujmMwbMo6xb0G1FMcXEidVqX1lPs1hjGs2kv5VChkVf9tgC57KbFQ/m3jPbDpPdIdiFw71RHDGO
ofvZrnvLSYESfB0kpBu12Ry+VuimMAipU3FQ37T+xyzsoKzr3hlP9g7oLeGDXOQZtdEPfX8T1+VD
Vug3oKWcGzLC7kOQ6OK1odzlx23ueBTn5t9dM2ff0uvZ5nE6nrkWkoXiyYlBMVXyeMaQVG8wZosG
xHEYJZPmtupktZalPlRn2ZH5+REJG6GVCkaghOmyISbKG8HQQo9IZmkiGI3Ks+p7BD9pRM3j3+JW
Z44lcrSPHnMYqF3NK449kvhLE2+qEPTeFKgwbEkL7qKps6GrIVlgZLbeyNwFX++tKpAsuO9rzpdj
W5YNWecgKBtZSJOnJc2vRKK6KlTPAbuVuEQdWSh6C1faJG0+z4YYjq1mBLiiUFSeJBBDnMfiKfU6
W4jY63LPlmT4tLe+GcCgVfmLOWpyVQ7GZWPtaaNJytZhktDm6aymX3ZFcZrEy2Vx/J85vS5YzDhS
NIRTZlzvZ3ONfW5IqKopd7TIDZBEK7MfMrrGDZdWT2E0VVg3aJtdRQY9gWhWZdy06a8EG6dELVSR
t8kikH3DQ6Iv6YJQj60cU9mNyGCTMg7sUlEzt0R25yiv6Z90oaFH7nfIgj2xYFYQkaoIF1pWriIf
H4XP/xRaVEiqpgmMaGHMwWMaSRpYIRkCsqWUnmqGa4H+23DnHxwGhn/M6F5fmppdN8yRbzZ37POf
TnC/BJGm0jnqsiq8An3khs1sMYe2cF+nK2uJY8WPKD8/lHx9FKVRk6xyZpT9V8HSXaLJEkzvb6OL
yURLUUj+ZLjQH94vmlo5klJMWsCXxXiBmfZRehhmDJdxIplMNd1SmpJAApDwOgQoQVI7ALU8mEZ8
AVdZXRSXFi/otb3Hhh2HmNTFp/okGrBi+7euRgq2f0nd7v/XhG58KW9lxrxyeGoJxB9Fo//Pmu4T
cvj8Ep1TaVNeeXfhE6Fc85f61BlYWwZa1oNSrkPy8dNK3BB3/u+831Tj8nGnSTxMtq5I6FZO10wv
V8M6htY6J9utwUIIvpzhJEUbIwFTYlhRFcpn3e+7Bl/Nm1/WX9IJPQbAWpCgZXAI8kZRWOnAjLtl
WSjM8M/GVgzvuzILyl4UZ7RqyqWJXQqEL56SOoOIQjda3KtWlp0gk/gGzP8hsNSfC1/0xXCy77Z2
hGCOKWHJb2OwbEo/Rm2idSIv+KeOesgnBTiPl5eJWGvB7bqYH0aq48FyXonhoD3zw7ZNVm+BCJQE
cp9eYFUxfFPugOqIM/rm5w/brrilWq2XynazEi+JMRXYnP4tpIWNZCGTdXYnLbw5y3ZDjpcO1iM4
h0lVi+YvlDVhmMpqjw+jbxdDznRRXF4fwkFfEP90x+US2ZUmkfvlaOxd/EOcRi4fpj/BLBFZtC9C
gHjc2UzSUB7aVtTRyuKqMm+eP5zd75N5shjNEnKS8slEKY2NzEuPX/dTA++yrcBDiCdl3BKaXU9D
MljR
`protect end_protected

