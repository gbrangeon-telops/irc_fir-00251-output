

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
jAc2elpDF3eoKND1/3jp/zR+PqlylbAiYUxqPEeJkonmmMj0p4wWQxczZkP8HQmv7tuBnI5hb1Re
XvZ7MbtjgQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
NcCSQniKJvfmu7+yh3FyGy0Ym5XaJUypJ6Y0uQPsa1akcjYi0ta/33mMsV5QsYvu+JmAYVNroROq
Kz/qydAoj148DuSUxGpr/Dh6K6KFEJQ68T8sjkHECM7M9i1ksK/n3u+J02M+jecJiy0HOyxQBNjN
TYNC60RH/oHr8eLrkFk=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
bUAhd9meaxo49J9KB0t7maJQYPBZ/miilGsGpP50LlxHKsJESMzras37N6FY41fj0BrwI2d8gwNc
EAnUne+xYMqJWaUJpkx5tkU3/Cq7YHGk19i4FrTEgtDQCfuJmvvnxIjd1KLqJ+tz2Gc83+JpCcen
LoaQjHQoa/X/vrkqv+GBi5yvXYw3CmPRVPihw2cyPAHh/aKqVK9U2rN3QsJFh6K1GPjF0J0zEoGU
HwvENWUy5CJqY+RhFtoI4cFMx4zvZ9LvGAYIaSHNcjGEuPxJtjqEiRDoZaxAPs4fPiQgVWKDuDze
FLb5NkzGHVW3Pw1VKV9puYBInovkYfTC4nb12g==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
yj/twyTkVkmohkM4L+pOFWHFJL5INTv01+xvkfId4SWEcQdYpyZZSWwRohyHdzU487emKgHzTSTy
GFDvnAvaZMJxmURlvGRprcX/FxMbqrYJ/QXjtyclneLv8hDwZCLiXegIMxugiwW4gYlZjMaOoPQJ
gs8ya5IBC3x9kMPV5rU=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
tu3CqLR7y72d6lMu0BtbwhwW0WER0YZdVAODwj27MZbWzMWHxGpAy3KeDW2xQMQiri7N5lQ02ec0
GWpokUjyJkcJKOv6cAVA0bMYymP9zM81k2IaifDaYhtB5Ah8VbDj/ArIWXDmp920Nuuu8ntuPKBS
17ifrJikBEgCPNkkESl85/+YxK58m3UimCI0iHmw3WvHkIj/sAUsakbfIOXt9rbFyqcIak6vi6kx
Gi83B53duhddmOvXqbhgzW3SRCCdyG0CtC/tlZjBXsJNv2kpjQBMBZf4BiACBpRjP60jLswfeEZE
bWRI3cRILGIwfm5V+sLTGxa0jiUVbd3TzGM7gg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 14464)
`protect data_block
SDO/aK+Nng9r+1crUf+hg3ReK/XV7GzZ2DQ2/YV4Bx48HUrghLUODfrAw+bYldUF/XZfUkOFJTQt
pDA+hwCfKzDAfdEvbhz4ETonypGR8RyjEwngX6msZWQl9zppzxmcPNrQQyiOCxrjOtFeLpB6Sdaz
R5Q6DA2WJMxlxjUFYggUfrLYsu2uoKchdC7Bb7CKr5x4MErxjlUcu/mme60L75R1SxHNdJ0bcy5y
BPEPKCW92HakZBfRr5KWSgPinE7e5SgYQTNWY/jhrvMGLV6ptgg0ZGAb1TDc58aYfJMZupAlkB8U
mnP6Uj8UpdDcxj7KKElB5S2s8n1oV9tO0RvXv6ifswaVe/F8pfSqSnEsRzu1+rJw/AAocNgzyRDF
DQaiTrcfVodpxVdUCuUo7jhXz/T9P1q02GovbESBCa5qU3sXTsy8HTpAPzGjOWCUWhdteV8ZoYIH
sVWwpOjRFYLA05nEWECmnCCrOrjjh2L7czaCZQ/X92WtERiuXhsQxPqu50uXm01mAJiEQzV5DJKi
qeoqtVwfDVLjbWu4InkXEmNpRFYo9EVBBUk9ZnrXZACgLFhwrlJeBNv6fugSw+PXB0En53Pi3fPX
72APGCeaVfJLz4cKGp7J1qkj2RBle9yJZSRU+NveA7pFnUXCgQFJkK1RDWaAElow1ttqwbalR34e
nbnuwjYpfylTNciWc5+tBBjj/lYjxov71GW9aKuLUzdl69i1huD9qk4SRwhoIyoy3zCQhqY278TT
Qm2lV7MJ/GqgOX0wO1YCrMDCXNG8ixXr8I+ZONefH2MmYYYp/O7FKPzBG4tvusGVc0x+ruvN2PJB
I8CiqR7i62xApdAQuYl2XJRW7kHBlDDEJYJgK4CBciysAu4uahjWVZfsorttW1ugAkF39mV653Y9
jdTzNWkUvcuLMmwhnlDhIvMUYNUZnZ7Y39EFdftM+6cgfgr3yauPJHqafMGc3KHVJgnhiiOR/kF3
l9wx6XEKlVKfhyxJhcZt85q8ZEZm1/iD27PWXbb7hoV+dvPIzS4AABV2GFDDd8D7iGTlOVluLcb3
KkiEV2NxUW/RrCk/UmWp91YexbvsNDtKnkA6NIRJ4u0sbQiZmZbVsxfC8Ek2jonEICjUxL7RQjG4
cLeaVFb0wCQvOJX7RtwLeROm+6zGeBuAAVaORowkKH6TGjzTYDpsddFs+wszkbuoVOTQ8nwncu9V
iGIRf66wHCvBkHO8lHLLTYb/8wj5zF+RL/UzDjfLVxPBKJjsD1MEhe5F/OXiHcl+9jpuWePRrbcP
g9cbA9qUyPFr8Yba/8MUz/d0Scswre5oc2N5pnHPv+iRDdmL+3WHD3obk6P6CSwiCUcVbetur44i
wdWv1//8+oWckHadbzHw07QSFsDGnjgUjo3Hv1UauPtHWLOPnXcI9R77Auy7CafawSBKJLtcxjbH
YKZ43Qsv4BCx0jvUpuwffMScLHWZ3caeA1Nnrd6UGY9MIY3FPQ1oAaQd4Jg6bSolppTS/7TdgdLN
PQTtCgIxGmX7W/dni7OnacTjVTQ2FVkhWYN/EfKxYvXf4WRvXoXmgXU4iHH6M3N6SyWHsI4WEKV2
71l1vyN0ZckhmaYdSurA1sb1ZTufWzb+JUOmysCO8xPVN8RfFZewYBEmflnW5FGPWTBTcMxeuK9n
A7rwG1W0BUW+JkD7f0Z3jpNcO/t9HX08yJBMrbZRMq84x7FLD0ZpXjOXBER1oC+ZfeTRlsUx6rdz
2WDIPAq2qO1ETVFXp+d6jDbcQLxWuqqnHOqoDk1QCLbHAGq0IbQ/VddU8gosHzuDHfVP8DLTKwG8
qPip1lx4eoxcBdnYcoD717fMOGfGn/LFlLa3vQaKp44fbY6kLk7uaDCJ0zIW1rZXS0ZpbWS64/KH
j/DwscsIRa1eN/Zt35Oooab8RCww2YzRrAGKOlxD+IfD8P2H358JKGO/GXeLiZ+JRfNF12kMsCYf
1C/DVW+/n+WfzwlHKask3DVJJtXjJaD2ZcP7x1aD49dHOoLUDcHvM2hybHcUxWcHqjsz6Q1fyVGi
/qk+an+vE/KDOk69n3dJGXY6CdfqXHzM2HWom00NJIaM9/BfMvkNuYRwBtmZjXHyb+Gzgfk8O/qN
WpVqv6YRfmpusoi68uYbcMtv7p/Od0UcaOa71xkX/9/CoczYRgFbuYw/dxMyNi2fUCsLQGyWVtf+
mQ1bBeC8ZdLWOPL2XErYCXucPaiRTuYH73tj8qHJryhgpaLVgUd+qg3nmxXKNLZCt9nNoNuRSOSe
fsSRZkNrj5Hj/yI11xfy45kIYBTOZYmjpbdmT6UUCYyjfoTdFi1S5BHyUm8wVW4S9FCKHHilBVvt
l617DIeFcuCm/Fm/bc3wzgYnW9tULygDLWgpPWA968SL1KF5eL6HOW9TvAZpk7BF9p26yryeoVAL
MISTro+nl86b10wmkkFv3kFwfTHWsn3MvJ7M1fS1KU/1XEq6cjwFBlUxo0Lwpal4jdwI8CpAFEUH
D09J0lOZqKPzODFTSSreSvNLUx1TaNPs4AewEnWlIhUFaqTCHDQ9C7Pomo1sa9lsLiRaGUgb4Sal
sToHWDTP/U0mWvKxO2363Sj+JxZ7iSk5KYVsbPjz9iDza5N2ZIkecX68oDJ9APL3yYv6hSE6phLD
0++lHFK7DPa57S5S4PlUXiNAMf+Agi3gzIXvF/rb5RF1Hu8RzGunDMCUP/NWABcWbMYElpg2c/03
4H3ZPzkxheM2Zjh8CvMOSvjvNJOaBy6fZtmZRg+gvgtky8a5d8z87HKeJCKu0XroiPaQt4C9VRyh
QeFEdee7usn5dWVfdG+5u9f1C91z8hENBia14vlcIf/5Xvig7bynBRLAmAzIcA0SXOmtXdxPCKJi
YSKiREj6I40Is+NlVa9gMTIpUnezvpUziQoylvMJtyBriQ9JAGha7BAGuOFdJhl12MEerYijlrIc
dOBZQdWCqCRi9fJig1Y0pPwMIGhIEq/7e+UqG12xV5aty9uKeo3bI0qvlUbOA7stGHqRwXzoNveL
iW/G+HnnHmbZ5Y2Lw8e0sVKjgosAY2R97yhvI4viIjMKvU/oxKGf+nCl249FMJhu5nF67rwS4wss
j7GRUDItorZEF6c5qtO1WxDCURAhUQUpFGfuz2Dk/HPskpGWIvX6e5NbQ++QUcN4iiIOHi5bc9NH
Ti6oGoEnPsyC+VY30B0YgaI19+d4t/mka6ZXy718ZWFEK22+VN5oWwTZTMYue/64vsvq65kdDY8J
l6fDvx5FsZa3kffI66SeDI9FRuYs/IDOR9iXp2n0Vsx5rNGj9Vb2quNmftPxJwnJoCNLmI4ms374
CHwNp/aij7znVLHvZpnH9Rx51qdCy32/n2fRsRi8v7K1gi+5R2Vwma6Y6cjLe6o1LUbsKj0nLFsE
gZJhtkIKhzoP9vzuNbVYDCnrWW4CwSGpm6fvY7Ed9ZF3//d5HiDvszroVZDq/6q+Ivd0pAtOcTpB
fvGX3HYkh1B894Yis/RKup6Fv6wwam37mUNwq6Ow2bYsYO+FaI3Igva6tA9nReiZCWsJ/tl+RRUS
Mx80Nhwv7iRoIPyI2EZnNES2LU4LT9hLBGxqo5bYiAzEP1kIqUofkQYs2UHnPDt44mzCvWPTr1kS
trTiRhvZRbED7mlQhDlBkCbNcFAQ1Mrh4NJxr/EjLPcVxvAMgiH0NmuvYS+HR7IpGRwnStYjP6EP
H9pVJeWGlGxTJ0wycXVBuPngfSCAOTYOaZOYj1xVMcwGqr7ESm+w6YPoS28sOHIpBw8JOXqcKRmN
R/Wf7ijbrTu4gLb9jKdidpMKhO39q+QypFu/w8cHEP5db0YNngHIvRQpuumdRQlOtoDGk76JqKHR
TYsWJRS3bo0MuhBVyJp5SIa9JPU83kesxOWCCfCBVfdWS1fifoASIgTjnw8k8j2IaQ95Gk3ADZns
KqZ0FJkPHiDjfcDKlo2IOPTVRLVBuzT4w1+QJHF3ZHs+GJZma1Oh56AMFBKABkgMPiihyu/Et7Rj
cPDp5qbCl83dcv2hAkJ8zQomp6KFhdWSu9wwV8qbWjk19BswVZ3m8FFo3Ks1brQF630X9f7ETXjq
G5QOwoADWXtcfWhp3YPhEyKUMoNDJ5FYTBe92J+PTfklOIMBF7l5pzyfzbXbyVnALpBnaHQGvjQw
Pg5aSVuvSYIDJ+vPSHSeGxgBM3zK2YyClndkMU6QEIt6XRLXvOxj7w6TLNFweXxZiw95ydnJCZEB
SKhbgLIslGAw3u5uxMGMp3sWzJyNo4VbKK2NdOUF2KlrAmSgONFjHGu7n+G2EMHJmfPeUZ6CtQga
k79vedsYo0PuzDsC6TMF1uvufr3bAcgRE5MxvnXuhD8BOjOnLYFJ7VGaC9htr7v+x/K3pxoTyO78
kW8BRQyRBj+a6evHyyKSxFyKRlT4lf6kNaKroCBsHWNTP4+1ildE4V0eOInIW1TBkxZXwLRa1b79
SypNW90QAVIUaw2lqjPQL/z3MsPaVim0ZiEmydGr7WqGfkfksuKvrzwAtsznmD1qRk5hzWPlugW8
vFSh8SiiwAevugiD7JzWTP1i8Np2MTqS0cSt8Yhonli1i17Ma4Jdf1h6YVO0zyhB+FzmyvySaWWK
X94qdrCzQ6F3F1qqado8dqvBjJwUy1CasPsLC2qYrC2sLfQQxa+p4PZTcRWkCmM45GD4EngBiMbR
v3q4sLCeGiGhU4i7FsALEV6hlZ0/FOg9kyHMXrSVchIqMZzXVvbqZ5/znEy9voazOx1SoW2RXyXx
0lTgqIpB9GgQvsalOET9iFIaubSS9Z3UaiqKYfIx43CShf0GuKzllFrhnFcSAQvkeWduA23My0cy
MMLbJC4izTee07vePDbQP+jDi/u9oj92Lw+7pEAjToAZWz9NVGHOfNa/MjGi4mRwDML5nl0+s6Eb
Pz5sLbNBU5qvZJcdQMDLhTyDUnFOC7Dtz8d6OwsJgHtxTT7JUiLssZjKam0lPYpw+N4CLoatJZ4O
l6L2AI8f74PrYh64oimhWSGUL02oqQkVVbC11jYpdlImHNI+Lu/RZVLLEHATJzgpoIz1MuToxM2x
AjEBDp68XX9ux/7C87FO30X94HJoT6sDSlYikmjGOdRIU/xBCVWoQVLmKPOk7bWSD9d4vzIgVzMd
kgMAQIs5dFHJjCYTStsDypCs8wFpFC5KdJID1xXojb7RKTmNIgkCBmLkgvHAl0alNDo3DJz7PrD9
5LytSE2MpnS2kMsLnaO2kO75Qza0DRvzix4fAgALxAxwgJDsCVSVojG4/Sbicxu7CU5Kd3wBfC4B
VVjp43u9QYHny9M5y6K3tBKDsC6maj0XyICem6rxKhFVH9aPkoDECnoIbus2Ca/breegNvFhX3AD
7/o/zyhP8liWXOPclTv3BS/V5VJ6vLQoGtG9SmLEwUAsollGj4M7q3SKMiHNMq5nbvC2Yp73wv9x
LEZfx8PBMRurZI1rEP4TA4W7EzHLzTSKkIZ3DLFqwXy2pEUIh2ERmrpCzYpja7cmGGKdL3onVzQx
oeAOzhu+ukKWpeZCy6bj7Z+GavMLn+GV9ShCwIRBEAEJyR28SR+UjTKKcmns9rVXCqPSY6YVWtVD
JrC1f5L2wfkfSDukrjGpXy70vmC5LyiNHSOuVoPr/Lzg7xKcR5EYFCPtXQa2uSpcw3cssOrj7CwY
Qy2ZXu+/Xhj3AS+bB+IwP3XiyHGlXw3Kkl4t8+mUF0Vpvm+QiYFIkd+30QagKuhK8V8HJB+5cHuq
iednnEJLVJNo9dOyluQyWZiKDJpFwnHsr41rK8jI8kQpJ7/ztCEK6vAx375K0v9OsgYa8sIKLDD7
1orSa+FIe7kHliLfRWMFZgqh3KNQC7Kt6ryUXr+XhV2wmTlJsGvDTVskf5ENotdUIgOm4yUADzRo
rWrpAsvLkBlkcePoHbNaya/ost7SzE8pkzQYUZov5c/PwsAYgbntgjjmxpWBlouN7NzPzcYOzBaJ
CM5ktBX9OuCJANQzYlud9Dd/tzpbUO6kOcB9VDHJwOsg0cSx7go4KcNw6qIjmRbMDYIHPXd9pJY7
6SodCZ6feGwFco2QPDdfkXDsR6lfQXv1R5d8dzGX1bcQQlWNQOiyF4jKfvTn4n3Fvl/UUhIWnELz
povLePdfYQYnJsFU243MpHdIZc6LMVOSRLYMuVu2D/ts6IKD8wHznqVbOcIGRRPOybNLA5rr8MOq
w0rct8wXC6/tzBFBqErQGF/3QZ8n0NpIqln7Bm7MRYdjdeo6iB8xcfnBemMDSJjv0zTxn2CTQi64
Bvo9Rz5x8OJglTqfxlnWiSULWsGgYWU9oms3sgQ2a4UKnO8avxv7V1+xPGkydVE/kUi3Ed7EXSjS
nUGaH7+RyqzI+2vBVrpKruP9DYvKTS7zuOk1CCdrxWk7hjmk58qH6iZSxu1IeeGPFYnJxJqHifjj
6vAit5VVOGm9iqFwRtrxqdf99djD0g4FaFzqbC61kQLz7dXZlqL14288wIcd4FRrv/4k3A03+1rq
cWdPiKgMuuGDgUsbkTvrBl05s/Tb5Pox+XOsEEgARCCHpbbkXBMFpG5C9rI73nnpvJzuAqU/jHXq
ESKQ9om7SZlWXSZZB3LrrotO8B5O08iexmML45+YRhO7WW6zCqx1/+wa60kEwF9MabsWiW+QuQfv
T2QoKMv7C/BGd/LB/oRQicSTyOVpT63fnoLPwL8oRdMXQCakfi1hYdqOmRI8CLmMTYGqB/MPGiHD
Szdmqo85gG8cWrwIBFewh+nsPr2wmR4xD/zfz30sih5AUvgpnnUBisZ8v6WuWbnZjTrEEFWfCQ+m
R/bTiYu7O8tuwrzXQIX7MR9AV7vITeu0NXa0XPFgAC7724YFy0GJ+aAxHdRhthC2xXNB9ZkANj4o
bPP11u6R24OsosPQVu9/6kjSJ1eCGsymtXDjkuXg6YuUQrQsXfPEqeU/MB3RiE0WxZbEy0YolYi2
nQWpvnVG9j2vrn2Ikphbnfd9ZgojCZ+VSNV9YI52+MzI1MuYoZDOdIyWoh9M0LSKP+/2Dhg6fzgL
iWwGJVEtvLDbPKbDAf0m1eqMbGvTyv374STk6aLbCcStQWVCga7vcb5umgDeynTssTM3VfDw+rzg
DeT0Vcr99Et9bf9AJ/iTsQ7D8T7ruEDSqir0haVk1Ysr475FTfX/bmVg1miigAkqmb6G8mEGih2+
+cIBqgCeevIBMmvbKHpnrK9fj6k6ExvaheD7wXkIgRliEbZRFbzrn/6Ir8pvmHhDv+KdAZ+ohJ9f
owYw453t9M2tKSLAeDqu0UNoK/IpCkRgurugJXaDfod5tkQzCIpKiZGENvtN4iwi6+rTiyGAVLPS
xsQRLytmin8TXlu1yTPzoLjzIVJoWYDwKqRjqWKYhmF8HegG7aiA7xNZdCv5uH5pXmpvZL8bGnrN
OgPFB0ZzNlLQ3d6yMnfwl2E1GELWFdIaTw12GXYPxsePWjXjZ2L0fPboIn/RF88O6/UW2amhPG15
KeVs6zMtsw5AKKqTtOmIJ8pvOmxQcIijA/tByl3Qvz2Izo3zmSUYkXkQcJeP+XY0diubk4veeefH
zn/wex0m1HfTxCewMa2Z1/ClEys4Zygg/ZguLMoS864c22YC8ObF8rfC772kj62w6dM0VHqve4zf
+ny+sSie1e5dFLBaGxI4XJzAHxeO3N58SlDQwtR7eYSf7N2iA7GczI09JlqS5iDER/Nlx/iMwVbE
lMmdl2xgJZtB0ab6g6q/0ZNFRXqKy/gZeTxJItV+5suGLAG4yirOMtKJT1YlTFZu+HRq9ULyssS7
TnFws7qm5ImJo3UUfeVbhOvtJ9i2FvQtNxlCfUGGBZDhLNMT1gnsenJtJAYTUXFIOg9X5Hzk7KBV
T2lLU2N3KaOo5vtRnVo35YJDsGeB3S3zmNU5xsh+9874sCu20NKlW2NSiky9QGiHZS9KKt5u6gL0
hwd3tafmfIJtILC+IiXr9/32A61IS3LEu9oSFw0UYF4rYgzr5sqyKgtqJWKXyT0l34kbPVhLFojD
BrIa/AeuoTBSaV7auyyvlZGhH6VyIlZP61DgvyrYdOb9FVbf7iwYOMBDOmTyH1Tt4S8WDtpiAHZw
VZRgUSmxi3H3kfDPUhitmhq7dDRUoRJOR1YAVPgQ2dmW1f6kcJaO8prKseP2lrZePUfKtpJilg5h
zCecqgcOTTXE7rHzQRA/SHqiEcG+aoYYKYyyYObaz4iqMKU0F+A/LsuzTbz4UGn3IVxFzB2AwSHH
0wrJ2ZQABIjAN7aE5Pd9a+q1jOkX2IkdGGKPo7tFTl9yW6xO6b38J6qgdI4Bp6/QMfW+2NdcpFDi
wARZxfIpKensqgVW2g0uE6bF/xj6SA25Bkh4BFbQW4+qwz5IbWkOwBbzctjecxmWibITquNAPKrE
2UJzGCzSsRpUdUSB5EBzDKY91SCKxwev5YN/Lbmj8Na5bicvBd9vlJgLPZh0FJSvvxgq7Zm9nTl2
guUOsf2I8uZDHHJKpY4FoALyMAELQqXtOBRKxnWtyv0K0gdAQw8bCW/yQJGtwGbFvYSSn7FbDFFW
vp4VDD9WyHtUnWrmXdRK5R1WOP3HKVvgN8o9CP4Qa4jRABqT6cXu1mNU15BbmA7+4M0Z3buaB/N4
bw/quiGQELV+crfjLe4+8/zTgXUXMvAoyTkPzy5ZLBGU/UuzCwgpI/VsMI4PfGWoim3m5LY0vRo6
bD9cyPSg0A2uUN4JbRREQCaS4bro6/61oWBBjraQQ6oAqkYFaynI9yf49ghU2DfxyytOJL9iN0ZE
zQwkX/zTAAEbZIo9QXpSKxDRaX3rvHiAiJKvimzhOfHAQg8KAOKX73eJHY+Xeb3gzaWqSBtNIgoo
AXbg01XNsRD5zQBGBPebCV07pHKHd2D18O6EG0V+O4j/Xzq48QmAbbfbOmR9nzYZEo5Nn3aoPWHt
wLrlvE6eFCoRbsr7eB8jiXpfjtmQ1zGLsys7gbNmFZNSdySs+SlEm1ca1Cz0HnbVvkyqHw/R9LN4
Ze1itGfbHr4/n1Gg5pzjQtvQRc7D3VozeMLoEgGuh6n7qKa2sHmg7GGwVrCFU8CJmGNSvo5kI+lD
nidN8jqFolNJt1U1ePj0cWe4KuZDRXm5Ii3h6NIGyN/4JfPsf4/dF26u/PhLieE2RbDRNamx8oQI
tSVURd5/svKebUC9q9BbNT/mnJi77UtwbaKgrL5JbzJW31oj5pOrY3dtWZLaZ0ypSTayQXCxSBTK
zxWG3pcfKzz4bcvrOjm5oFkyO3iFeLf/Q+PUBTeyJa009NrgECyYyNPodSfI2NnCQokTkWvw8UCb
PYG+AqirOU/0NIm2K+CFHv8O1RNN8/9q+uv++05XRejrSeh9yujCcvuu5lhV5HG4Y/QxwIm/3ACy
rJ5sCGtuYvcNE7Et8EuCYkJiowX3AgCdhdOLVyR5wS5VGeJmEgSKsvUHRBbWz0+QekCqIOlIH+8x
YofwcNHKobawcWzl1r6K5x3LBTccOh2mLYm86WxlDKIzN3dLd134eD65/Fa4xX4IMUVucJgBBTT0
ct1gKASUVN1jpqIRWaKZxj6ZTBtBigJ80IIOPMT7bFRj92urXmSdefCOyz9caZ9a7dFcCE9ejTJc
kYweB4cIax2QU5X8aZc8D/jNxGOcD3yOfn2tPMD898sCk0eJs/qhMz67tmq5RYVgmSdqW5gg7sK0
h41a3E76fYsi1j/t6KtHzIuilfAtjmlRX0dmpMtgwyJMiXedzOOP47Rily0DzXT5qHz+WF6s4QIs
eEGATTFl4hsWVLls0rfKPorEEY4gdWef63ToAs27ek4QGN9Pfup3RZ/IWaCGjb7xAcDI4fdZBiMs
eRpNwv02e0BBbfT+zY2ngx0S9vtJQiNxDH+MUuFDuVn6G8izqsXygAb666UF2YaBUexMSEyw7+PX
0W0oPin4o+9CMM+siHSqYR1eb7r0F7bry7eQQeof54786EZxXbedhWO4V+p7if1dj7gR20nR2dSk
a4GMqhhJA551SBX4cq7aF5pJY/2fiBQK7PzPscih7ggWEgZh7RVTixJWxWoEbsnJquZ71Fu2vmq5
48R9bGG6kKdOfa9cpGHX1Nl2JgZfX4hD2hKksnlFS6otZ1xp/XzfJEWtdA+5E1BI+0ldHdkdFQQ1
PIiXS/+WhI8ti/hhxh0eGlUEkRx76X43bpFeZzRW1Hch13YWIQMmCVEXsgYspeMYu+KlhXF1WtLg
1Ro/tA9wPispypTTmXw7cVh13Xlyjwuq8JbjE1O1tEWR5S+lW/hHr10hFDq5vbEm9qRMHqUn0Wew
Qe0KO5PxSkmhBPp8DN3OGcq5dH5bfgL19WNqKKMTvr5McHRgLADzYIGmIpUlQld4NA1iSr3rVYgV
0excNP0VYBEVdj6/gWO2NrMNSe9GvXKso1vlqInoS1LtWP71C+1Dl0B/JJ1M3GxD6iKHy/U7LSsC
aP8oJzhHCWwXwUJ4Y7npUTEbaS8cW1lJvYU+qPZFYuQ0sF4sBQgneKHzgat5yrhV3zMQBr3hzo6Q
qYuNaGGPbCO+hEohsPc9IujIbj/L8P7gaqS6YXZb1i4MPi+zROI+dP/4lCX09iHYa8hwu9KnmNe3
kpuYAGtE1k27c3GwL38mvw6xcU4FJou1GRE5aDhFrtEJSzT7wKvagr3Vmn6HzmzCKKriLKsFLgAt
tsbWa26CUS0BPry+dCvnF8iZv+laJAOlCNvj8XvCAd0ZlYxloi2MKeccg9mnpL7OmF+P9O32tlCx
20ZKp/truUVIuoiulDqIcuUSHN3XQJ7WnvP5XNeN/BWDYJ5OSlA7x2PXiSKHI958vaD6Gr3xPavJ
0NIAMQEJAM9FTKftkzvbiTBs5rZfBEaLoIFXGJtmC7PiZGyiB8TKH77uUqScWnU0ZTljjHLOjbcU
VKzf83QVowNzdA7ugreIuVB2IAZrVNSjux+mSxdZbhqi3reV4+h6Nz++xZJX/4cxaAtDjQUQ+Ghy
Cf5qWkOGiAROYmy2y9H0KqC7JLVGeB1HUwZniDH/TBawq/ndBW6Oodl8mmzFuM7YrJlqLybS9Pab
NiEz6DIlZk7PvvDr5LEAVKlHhFOs4MSX9Oic7m05wPyDEQhTzlVjZ3d1BsfTn/p6nSicVkvwBc82
TVI1HKl2WW2IY81W4If8FPBRj2tFLTa/QVTFCp7x1meb5/MjaaTjofNVfA00Bwc2JTMgQar10llg
wNUz7H4ju9wG8Sl3WTVZ45+If2xh3jdPRXBUuJIMJHbBl8pK+p1UsR6S31/j3ykptFIjMqJ4M0i1
9yXZ9JD7CEM6vN6VF+jT2N7g+wfzKASpgioNqvMXqGMR58fe7pWy+A6+MqbUc0pLbjMmlMV7yVqW
xgjc04sIh0CTRWbdeMAqAVzR9nwJ54UKCqS11qjNcEKjeXx2K0E5XGmpU95WLoY6bD1jlP0ycf5f
Z5TyYDzsTSG9nO/Q+UychqpAkPTlEBK5N7s8li5YYhNnTEQ6mFjc/9866HyTMItVreB9NeCHE9HE
pcbXo11Trse0oFrLNvOmX+kttAKQuRgbDThIQLdsoOachGBE9xlKc2qfJZaMqPKD+xA/bFSHVbFM
xCU3f8DkLU2iUCNrm6LDV+1aCOms8pwyFNd9EjTsWz6ImGgCtTxeT3pfkmmOJjO0oYeCnhrmBkpW
SXqTXh26xqie7c+QzkjYm3SPWS+wAJQCmukWATypY+BYvkOExgOe9oyNSgFgqGYEF216GkM90L9M
QAa0XaNsNuz2RYgBLTqSvpZiod8miuYQFkFG/886t6V2Rjntpn2C/MTr35kQqSsXzncsCD9oKCLq
RKHGz2dXMaxaLLCUZbtwiucyWygRaae7zmEVR5o8zXkAduUttnoyBfBmfhzfvAOrFr9iw6fo1dpj
qFkyx7h5gjfDQHfZpnVrGGY/jFyk18GoGGG3fdFDcL2N+h79fUvRxeBxBB2uwhPX11C0olmtMxhI
4wcx55EMRfibykq/nJs9YNtd2IWD29hMFSV5tcbewsHVxaZ/ecwygnlTl8qR/WmBljgpYJi17ZlR
JX96kqMRBDdJGAQFUmHCIpFH9WhNwFGebaCMWpeUVc7sX7K64IIgi1Q43Vm3F+LzVolwP5xH7alp
jObnViCpJYi3d1RblrEBbNU9Ye5L7gKb8Az2tA4QGa7vrVjtuzDWNkL21Vl1/C/w75DG3uu3cL0P
8YevcGLCNHJMyYAqnkckx6ti2d2md5rKfv79USSlca3G2CgkCcq64WcrrbR4vap98CPmQpPcEi0s
MzxFYePpcTrRF4ZaQPuNNJ71KZIy4wIwnLtOKjyA789MrTA0y/NIzwBHqANixq+2XnzNWBWIFETb
6t4qmPrB/sxb/LhCDa7pSwdvpvvGLuE9vQTiMjVkKMO06VgbXTHB4jd2w6rb5oP/YoAaUg6oMDej
iWw3Deocpe5zApP5rQR8eGecuF/tmGCZSaaJW3jOPzo8sw+Z1vTAs8qUKlzry9pJlgpcz5aZ+k6a
N5Ltih1h4cMnG00ijxnW6exnO3ZfPJwipHXQ/ktw2+DNoqAPY3qAZgRjJTkPZezET5JD61JaDKsJ
JDYmXSxSI9q+UoIO8Mx6AwkYpx5chWS6DTbogcf0zLQtjtUR+M8bkwsLnFF8scAPFVch75jIJFWG
Bj6YcuWoeSrR4MQArl5I477DmUpMlTj3gHDzP7p7oBy58is+GS83HuEpSoFSpoCdpBARAa8jtVts
Q3hHByZzMnJ9FZdz2Xbjp5hOgJP8swU1UJxTV+3WTm29bVmp4Uskaro6WP4388ULlGzpXJff2X3z
3OKdHR5MypuVEiT7ipNZPHWxzd66t0cMrzbf2u7aBN11AOaT0cF21gnQLsCdcydtwz/KvLCfkhIi
L3U4/oVD+z82dv1qcAQ7MRaJydjYEnxGU9uejMvOfJTeE99qvp8/c28+MfOx1wd6WETKW8RCW4PU
b7reHFf8+fRlTVKApzSPHBn5Y38KHvk1csga1yMeDFTZeSJBr+B+csRMUTsC7uIE7vWYfW/RkJnJ
zQh6IsiqE8X4L4AB4DEnwKqRWOsyb0hQyOdh/MXNpAS5iN/ZF4psuJg0ojSmdfhp0KV0SXgYaAwi
CcjZDHJ2o7urET+zJlLY6oPXIqNGN4DRUcfna4BgF7k81IFvVmEOkeMcEXo8fNlFGWmQG4bIxpQQ
70K6T0NkM7H4i3gQQvCZC/fcbVPWCMJb9EJf2ROTFSOmY3m+RM/EkYu7QCe4lGJIyzs4j7BH5F+6
SHYhrX5uH0Grk7afnGCIHGXSotlDRd6pJMsserVuF4/xr+zlM36kNtOhzJMU0oXck/Djoa/Wmwjh
xmiFK1lNZu2HHjYEDYzMR3sPKPo0MpCDPgeSOKeEx5K23wWOwzjhtPeRp0O3LPbdcxVxV8Lud1kg
IvWo5Alw1tcO0oQONdx5To8TBN0Gq5OgLxjh048Igz3fIEbkFT972sq/34G6rTllTwVd6pzmxEhy
J/G8eVRLcfeGBCWAImeeomN66Coij3p+4XhsjQJWhbRFXtD96xn1YIb2zvWPMqTxPMhE9rpI1Gri
i4kF+ph9usryhwYw3NdoN33lKjfTdOfZruW2xEdZz2c90NP9D1EVB27RuXAs9BFgzdVTNacWesCd
PnBUx77RIzwAbFGbebBzRSH/u2itYJiq9yadGNh0fS3B4VBIv03eXklZ6JoH37DFPJ8wJAgGHL9o
1Vzs3NIO6Nwg9NpMhs9IyU1ygvCjIN30q8vRYzT+HOwSRki9uHSYQTuFxk4LuXuS6rB+fzF0AM1z
utG8EKs6ayndFN6dFF3rEWuNI9DwTDI8AFdXmXHjGQecYyrSS37ZApxXYDCvusWAzrb/xWSCiz8U
tg0ow3cpl48NobsrI51WzpUNvS6//H9qXoSvWnP2NPoQxcns18TblixquqgX2zZKXJpJRyFG1NSp
JF0zGY7G9EbgfRatfTlncuRSGBwaJAxlFMWHoBZL1D2T08NajiGcUo1izcu3zQCSDFJlJWMaxH3O
mXafJaiV5hinEt1Fn8kt6ug2xtj306rCBh0bfPV+MBFmfUUMX+htk/J90M7QVC2buWIWljo60mUd
35WptL32AvCI22HKEBfXUk5Tox9C54WR+N+z2DOydg113oUg+78CgpqCqXqcsMvHsjNlKkQQ63sO
TzZiNFr8mnydhhxCaZzGMdg2UPKGiu0L/jwzTM/5UaYMdQmdTXlQtWWP6M8htfN8xFWrirguP3mQ
umSa14m4t3WXIaD80hfAK03DeMT7KpD/dSz1B7jSG0u7gh5fkNDy325oUFf1oOYRUjjJD4+wsYKZ
s+2+KjcQLeo4+IGA6diotRkJlm8fZ2v3v4OfjOftnhlATsCAWE8sYYfiGXP0X5kpetRqqSEaep/a
3VFZ2c0S9eH/A8ra+GsawtWID6R59xk7M3wIhp8FCsYPrT7HsjIdo9CFQbLk9Rn5b2rbCvLoB4Ul
7tKvwKhThEk2y9S1d5lSlcuv5ny5LscXJk0C7fwIlT4a/0l/H0HaRAimmxJNVBaqYt4r2jRdLkT5
le3WNH+ccVi9Lm/EuOsSrmv39fzld+VCSYEXOuTt/FmbP0k9caQ2z6+n7BnFXI5MR18upfqOgiuU
o8i2Xj0upbLtKLzqa6FR7xyqFsJ1knFCs19Am02Zjxfj/XC2seNE81+AKWiE4EPHbV/wpzPcugEi
pkO+KnbUeUfX7bezbmJncXjzCQ2fGTUI/jf8sCZ/n7UkqLRHfjspujCZloCXMu9xHGM2QFCgGP6w
AJLF0HFE8WsBlvXaMpaa/WEo4y8lNIajmUxPRwPonk1NgHKZ+wmhZTk72mVSlM45P2oCALO4Q5PF
X9HmsWOkTs7bot5j3wWEj/2hqLS2OMIV8StIlshc2RvddkZTHBJr5tUpPR2isDDLHQ3WAoe3bqzn
jZp2Tg7DaCSOcsb1MVA8U69b6lU/2BVL1gxHsU4pL3tW7xYpDKdXIibiPoQPinCPjRqRGh3t3/GY
NlgbS2stXroHo+DTYuk89VViLeesMIn2fr+8y3sQAgiLxjvKMiMmre9gWAelwx4/ZZMwan73ZYhg
ioEYKcxg3MErELVWx8RTdxd1oDqdAc6AoQDv8PGbvqXe6Ggi17eLM+/Ew2T7ViXYArgmJysDrMl8
m1DoX1qh9Op0S1HJ77fC0FW3M2oBhyIhZHXFpjEYY0zQTRivdXs3r5nVW0x3k0s/LYxSWsaMhyth
4uRGT9tEZ4woi0BLK55YxTdAgX/tBMKY9tGz7I0VDKiQbi4Wg/IqaDuzfr5jpRUx1Et4Qz9iQVkM
mLLQOhrh52hv0jbFK+l21EOPoU/GioRm2Uibyy2ZHnk5ozfOMHwztwM9exNDbT4szl1hcPVHltcL
T16Wp5vHgrMmTYRwwIN6i8UYNox3V6tYeUL6s2naSvVowWQAM86HLpkGan4h0DJW7ihaBFDQtqBX
G+oXSx0xtmqEqGasQLIzgUBKIbJ+9zCKexCmkL9A4qix0JuT5XfJvEwpI4/jEGeXiVduyAXdaEZB
lmEiCL9Kn0u56zGa8X8UyxAttjXvRqAV8fVXtXPDmy+pmN96GC7rz5JzY+gCzlLBD8Pcxj9/vK4y
mJKFulaktWZPAkgUjq3hiSrycEi2aGjCEWXToDhiliiM32c9YQO32fo+anZBl+FtLS4JCzG/6NRl
Li62VtG4z2YAM802XGwLgNKWbMm6R7L+dFQ9KSmM17GcAqu8QguqSM+Psr1pH+XUc9NfTkkWTycA
7R13SCLLo/ZcpGueaWsexycUz9XsIffTOvfwE9IAMK6BM16r9xcKkJ576NljMRSssXk3ksWp4HVx
QiXO2gYH2dqmkxcEFVQKcKw8hAf9YCQbmXShs3YxOxiHn4U/e6hpfBySAVUecgpD2pkBtjdV4Q9k
oILNB/XQ6ZmPNVrn2tohviRDlmR4eOJ7Mvf/8nBLQ7n9SzxAvRCjQjUjKasG/b7zi58KmBH2/zHB
kdExaEjVHH27l+koXBCNX2gwKJzGz8u8p6lEXwoD6ZSlRMQZqoglzv0Sqwd5T8yOsylLp3jdEeXz
W7YtzXao6002Rdzl2s1u/w0wrUONoAc2QVULNJ66cdL+HYOFh00y+6k9StFHU/bnALNMXP4WIbx0
X+uI7AjN1baLh2LViEbMynMDEsztj4Kzjit+AipaMCMdbIVwNIRAgBS87ceoDUneH3WOuMJhnLsk
U+G035BIJzMz//w6kaVYBP8tTp6M5Nyb/EqnhJ/75i1Xp/CmvGLKFLWYHHXbzAGV0n+T516v+p9y
X8HnZiyohDsS+G2Ej6904ZNUxAhIwxtQ5u6CTsuv9g40046qqUYFX3Gk3KSEQtruI2ApCeTTkXEO
+RElFaT8DFrteuVvSOBJcz3ujNd8Z4uLpAnRsPoNUN665UaUyw4xPQSnpguX4Jw+ecfQoyrHBIOv
5L1VtarqPKldryCdxh/26NsZQ7hI+DxrshQmdfeJ8nqeGM4/pTffECji1zmZWE5r2ZQHZ5Fwj8Yq
eNzs1MUBJtTmB7OI/RhUrkEBz9Xmb4DotO8L4X7kiATDg05HTS7wdD8HaIGhJXYpbS1qjspT6aOs
gr808vfT5XdFFn9+uY1ZwwFubWInfnOUp69xYUQld3trghaWGPP9e+B8X28S+Gph4JRKYEFi1Jf6
QTJ/Ci8rOOTyFypIC8NABrhOhhftolQWdDY2LQDaCM7lWNGeBahsurV7a/UCNlMDcpVHDRp3FNPv
Yb/iEswEC8b16lFG47CEN8Xy7iKHWfHZ/I4eRMbjEhsB2AhXAEie1n4P7N6zyOpoLZ/jcvnWUW00
IaE7VeBP3YNu8mmEBQSkgF54MKZVub3i4YASrAk1qJ4YhAd6XKQlSPtszNo3R0Au88SSnfdo5miM
P0+WmzwRBolWlIJq2XdISCOZDfGYp03oWP7kMveO7u2unZhdZ2PxDRv4FKeHFuDy7HYUKloobsKP
YKUq9bu8331HF0+wAXXiN6+Moqisap2o2QuN8ueSE/Qr3SS4bvQ75RBxIX7Q8fuJJ7WDY+laih1t
aTfyDZWIBz7KcDN1LymTmqX3Sn9ESjhF1VJA9vRF8yw3vElpNuSMNw3tAZWxANimj6XS6c49SvlV
DnoYVv9pF/ISVD9EYWn3woJ+OuyTwbG1F8h9LRotmtoZqYhMZH8Kezgz49wbyBrtSiJvISr/ApLw
viQd6glUeysgVyXIAtJ+jaSJL896zqC9+uIR8fBZnL9/JUIE1UfkG/wYbP+X5+Gqqgdh8SCSV4P8
mXaGVMwWj5U3+jtJ0803+YqYst3eO6u7ekpsUcwKti7R+5eGck2ooFx49WCuijekzWPrQXhxy3vB
s1IWQgyU0xdEjk7pQUtsYY4Kx1lSrgr+aM9e4dvxJDXWqo2TmenNMzrkFtbcj1t7t9B61mwJlCv/
rWtYSbW1cX9siRoNb4i491UP+Jko+OmeXNLqG1ynGbw7B6GYAHwuOPV3nRZ2DLSzlw1Y6Olp4XK4
76/Irt2EmxLKlAHirzFp7Y04PLYmqHBibVPexwF2zKuJBzCbWvzc84ECMcfDZJchMEjiPM/E6tRa
axo4J5u6W7riUGKheiO8PdijkjMzJ6ld7cXNy3WPPsyMQWNG4x0bxMCmVkTGsW3EgJdBwKMvcdqm
y/T/DDHq7yRLUAIoC26Y5VBvNBwM8Xd5AnJ2ksaZe/t7Vqasb1B1CwOK8U4xGky+U3fHbbLs7iN+
Xk4rM57Itutb9+r0Efcod3cKn2ezO8YWk/ypx+HDTRCL7GbTko83gFU04XtF2Q/Nbu+qJq+fN1LT
q24PC3pq3V1J8VEzfaDWekl497rL28NjMD4EIlIrg/T509F+LqV50DsCt76DOn2ona8ZMG7a32G9
jA8NCJyjCQHpzMBX+cEW1h/e6dsVTdYU6pXwLjXenZEldS4tPbBQA4SHBZRABYbjU7iAU5cu/rwR
NZJPCRDBK8nT/QR6F2XI9dSRHfAG7bFJV2c+QLZiwFraDK76GFn1N/FiqaQUY985HVcHjaRiVsvC
nZcxKNyRYq585mIIybnlgOBSzNDJ3n7S9w1H9mnbuiAzqWcy6Ft+ZbLrN2R3qfZaEXyqHWmWGFZL
hNDciHHoAdAmD2JolktsmiDXNUO0JViThcaRZuUMKQKh8sNC7vKepRlZiyLcuFxQ5lDxLefk8Da/
mqguCEGCOqqLOD1EsyAGyffPxoQQlL0Nn68VlQVyvN4GabipKleTCcWIX0rhE4lhok6ea1bAIh9a
i+7v4PYR0g6KpU1ibQ81qH07/drZoRJQSGbj7x7XOJEdj8z9KkKu6mmd9xOU7a42JdvihpJvnbuz
xiNXJmn2uQAgqGXGYFjdYM23Q14Vk0sQ5WLpntw/GuPEWpOWX9Hy6RBCSCe29xMrEdHD9tjd4RIr
uAwekWSNat8E2BIi258wTmLCjapkgtbjQSm6ZfWZ/Yk7j89lmC33aECoQnQFO/ZGaozLuvfZenoH
KJKHUHcb4zdrXLX7/nO+Stmt7Y/yPRpnB0Qds4DP31zPkGtS9dYtz4UIbOtqTuCNDrfb9qXtBDJ2
9JBp8Zyog3AWdWcF7W3uctjdj0GXD89Lu8pydYGFfXoBKLoF1NHepew+Tn44esPFd4Rn2+zLX0eH
XGYE17NnR5E1lHTg14bqex9xEongEU2QGDj/vIzPtzR+sLJe1Sj7qlVO4ws28aXPqWvTHp21J9Db
2xOj8+42DbAksk5Icjhw1wZl6zqZB69Po1KW8xIw+bRArxcD7CDVDw0UQau0gYCONoL0eCZUFYZf
lNxfRS0AUd0Ut2tMtnR0Lx1hbArgawYpRB7fYuTTk02/6K008OvpGuS+FID+5T68kFqsW1yiKZ+s
wGs1WLhurE8NrANArWYVj3GkX3cME9faFlEwCHA+PgCoeTq5Z/8rl4TCAViASPLD9/9zkeL+cAWY
iaZp0BS96AZ0JEUeHroOHPeS3W9v+HuOlyeVLsev71Ay2kGrbMRhuKfMs0peGwYpwcS3sVc+3OWp
N7Y38aBwMFSZn/gqHsFAN20e033wUOnbzqLE/Cq0c6d9nima6jsxYbrp1lNxnzoObvbhByEoVKX9
CSRd51gZkKwpWLLe8bTGvOH4vMjmlMJXwKqbRkNXw/ZSvaxQm/VCLZWwttnrz+scz3dTVRo3p0Cq
0QDX1iKL4gqehpYQgmfb11t47KMNj5D7b388ETi/uqaw3oyuKxHgswFH6A==
`protect end_protected

