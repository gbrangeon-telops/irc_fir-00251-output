

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
AAcalZ8o/jQY7YVFFozBN2W4CJ7dtDMmc4qCXcw+X1HsQOWsjlnqJ0ExLq/9HwwPaBdBtHuX8sNt
9MbzT1NoZw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
eb9fumGdx5oOSTot8dVQVSjhrvPnjy5/uUjD/aIEqv1QEwLJo5EU+m6JllUu7ONkl4q2pMcv3yUD
DaaWMJ5SKNM9IQtYV21pAAxck+unqu58lsMHcSYeRXYcYP0huhB41kbacBO7fQsq8URHfGRa6NSF
6GxQzFgW9OWA+QBW/NU=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
EWQNTRM+yXYG4PYEP5SycD9fkQkTTfcM6sgjpG7m3z8pRk88pPYs5UwluFbB09hVSCMPYEKLENX1
JIPX6A6AjJm02cmQD/SZk/c9uIP6nVMvhv4HT2PqiJbMwRsRLnp0RV8WJNl5IwtzQhAltPQm5tcZ
c9/ABn7qb82RSMRxfzibhF2Uc1QWD8PnV1j6nVmyG5zwtPXyKG+iY84QCANIn7Soa/s6m+bpOho3
0pAI7CU0STIdsIAbeZ3h93cun/ow5TnTga8aw0A3DbHVrLc+5xM9M4rs1eiVbJSSdL5Fc7sYK0UO
cAQhBC40rZd53OFEkTfLRVfwRFeSU8VoPsBCag==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
EUZqFPEsLcyFBckZdNISKg5E9SpkAkJYhYdYkwRh/xgSz3PN8kMAAO+ttVMn672EPHPSTTeJWt1p
AvumrJCguaLVBM7NIXSVbD3Ckha5a0glBfzxCIJFFOPOOxZ1B+rxQ2W+YUfoLzcw9DE42G8bHsgh
CvpFN0Szn2edsSc6Ou8=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
OK0W/E9mRq/arn5PVxkw4+3w3BGYpl3KNYb/ZgKXRQbbZBHdfBtfu0H1VHCuj27qhD0QdkPpdnd6
gHcvGTEag6clv0PLJ5PHHHzcIl4hIp/MStOr0nGLUPNhqZtLAZRqiy0IB5ktSoIvGu4wUrWu3P7t
D9RQYPlFcbj3tpqdazX+5GhWSHnpe6FaCtaWmer4ZDmYZIG1oGk2h3p7ggKQ3amLtCrg9RLkGQQj
yEO/bz1jhZ65yzQA9tlLPbVh4inksrXMkvmJzspRm61mhZF1ey8gENJN2v1TzCuN2XD/gXtMbo1u
8igS7KocN9wbd7hsHdkLAK4mTBcgTG5pa81agg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 998320)
`protect data_block
F3ZPclJvoiBPosl2GhOGhbT7RuBUQInyxTBMJkZDUe3B+18+JN3G/r1/9wrq78pneO7usZEjNjFD
BvIz9iVVK1rytf3AGpgiBfW2WsRLAbl/yNJUu4W+NPT2lkpzSqGthcX7+hsiVo7UUTtmiwRitJkR
I5jhFRXLPq7Cw/mvtcSExxf6GEYbJfVLby1eXiXaOHVpJmp8P9Olc/OsIokNZUR8H/F5gV431Ils
w0azyn/1macO73Ysci0EeS4MyH9SDAuiR4jBEuJ8bWBSIlDmssvUiyG7s2F2O384ddmt1c8S6nXb
c7ppsHBTUbV8A8NCwZ58SsLMdRgEED/iWdhE5EuuSypVmzSoKD3l+1z3ToqxFAcGXyQrd48DRq3u
W3JPmRx3eumE8qvXTVb/Nn/97WQAr+nVlYiz/eDiQlTPZRKH1R13T4OCoIHHCfhJZJyqU03h5dY6
DrdwT7G1UtXnvp4mxz+XfRHFVC96Bn8cO7GNzRvP34A8PjwD2AtNgFiRnKj7oml1c5ohnkLKdwtT
utKWvmw8rfSZnLQ1duBOQNS0kHMHM4zTYIsmLE0XFPN5dlZdu2Uqa+GQjQls1feS6l3C/++Mz6gj
WPCq327n4iqfm7YKE1hCaviNEGWeM7wA0CV5a4LSD37BmDBHewurYGKjy7wEvNds1PiHthL4P9XE
zBKoKnq8JqXB+VKiKrlSQvz2h8mhvxsTAffVB4SWWu8NAid1r6pfuiMe7AqShrybe3fiLDBII0Ou
10jqeXX2IikvF4zKIy2gQlmKsHnamG/QyGY7hb7SEma3Hp+Xc80hTvLEK2jt9FBgDTuxEXOHATRp
SHVoxDU/dbJzyhSdVtBHSV3HEo4Hs5/3lHcMqN/1AioNJZlj/qQXB6StDcRIvHmkP86HQd5NiA6G
32bsbI7sn28YXmQxOToQ1+MqemUoBnKYKvTZ9oj+fRqcF8L3cdJfsb/4HWDM9xYMkOMCt1sv1ciA
dSYrjIcEplp77dpsoTu8ds6hiUChO61PAEWQ/ajjFFW5TbJGS8yXaZ8dLff/XHwf7k2LFTFrqeFT
VnveLN76mkQDokUYjdsQnILsDokrFh1v+TcaL+pNY/iw8VYaDNu1LWG8fyb6QppEQ0BxqYAN1J3f
4Hq8IfiyX+cQ3+JxIEiv5X3leyM1WX4CKSTZ/neqRgYgyY7+apTvdrEC+lLQY7iiSqN0FqV20G2o
ytSmND2B49cMhpRSG7o5v0btPKmrK2/Og2Xe2iGmg0PtiTawaqhvKMH7C5CvT8K4dPD1VQF3rVTp
r42mufnMaBsvQJvFjkQmzG91tSiKT+ugab0RBjLWki20ARnKlAhno1IdX6Co+Y/ea3YI8M5T5HYj
mVy74D9mfkQ3nMBAV2GmwX8QXqV1JYiDH81PGP28zcOjKTO1F/rruRACIX/oRNZK40xvyAsg/evJ
03HjISZHh3gknu0GfiaptSbHEOFMauWfsszHaDVi5wjbJgESVOU4c9n80WX6NCAa9q63EgVeO/E8
OR3TiX95DIoMYLpK0q25iQjaPVQURyMHJaVgx38L5gujreMppQDpEPirZiYMomCO+Ah3VO9MVhJO
rCsdmDdOSaVA6BdTW3lKEJbV6QSXHluaNGOryYGHk1dj3lxdRpjXu9nJYmf3z9YCzSWzOMpZTbWV
bj8YnuJzhKwBEq40J/09+Xeib8SxoTd6zTbYbWm2dtkZjW7IFldq9S3lPFEMXFPxY5Z7qF1h8IRv
1ZwfGuUiB6d4rDX1w8/62Vjzm6jj781xX6Rb/wX8wzkplt3Ot06icF36XOIaBuM1L97x5fQlUNyA
9VZLt72CaPvi252ra5AF6SmydchYzJxPVILPGAHHWNTvow4WpwFUCAV5901qMQHUon6qwIpyXWhM
vwEFslojhx9ThU2HZIzUYk0Ras2TzR97qRSnmHwGX8RWkBp4Lv+8hFVKibd4opIJvLjaZ/js71i7
raVSehiOktJd7fR5oyn2lIKCkam8Q0CQ4n21gDZjwnuNlPsCDg2J5hYA5l3WNYntlKLa2jnaOErd
RjZfX8qUm2tmt15+w9Ld872ZZSsAOCRL04vcxhc5GPiPYZ6c6oelsGJDE7uZDiNq2vzZie946Suc
kuiNkk8wu3egxSzYHXT9BOVbnigNDTrGztv3RT9ajc1UyxECuaPkbRokQa4Fvu1ahYgkjkQUP5wD
yhTIL5uIv57lrprkcsRgsUuriYwEysx8iEtyzpTDP/T7NIXIHX5vKYAS58vXN3eWDuV8I1dgJcOl
/QmnNOw1e1bsNk5RHqsE7cFgrWNHgHJfZV92Soq7J2xDs01xBSgBQtHZFQfW1KRch53xDtzrOeVI
uVDDE3/ftYcspaxvwXAbakqhmcbsS277ony/baNBUe+wWvXGuveuRZ+eKSFqxDA+vfYP9B6LkwGR
KCKBPWe/fmazcQ4ZDGMZNyNqmqTZe1CEQmHCpuD2v6t8Zf7bpcRjg4FxzxxPBDOJodqzLOAM4kSE
WI5yFEerfY+EuRQrBNZcm4CQIotZJj77f2a4WGcYsA5w7vDA3i+quVQo0Os8A/wWrnPAe/ggtWDg
TkfBekAurjyaoCrQOkOXPJBr9u1XO7yw+QV3dSla1xJnPIdUvEgwGLmmV19AZtUVyfDySnFzIy2n
4SX7vU/5ij1JLam8b96SOUqz0KvEHOjCQV/t6YqBP/t6kmkhXCr+zw9sBg/XZVGDqWCGIRBcwUji
gCBT9xFDM3gnCDw6vkDlp40qaFfiBvqYZAzQDF7KyB6JviFos7tqwvbpaurWum1fz7zwJIXphqmU
ssPp0o8LV3u5ZrPpnQ/47xf+VHIZMflN9NvQ1HERhaSvqWhPDNfZOAsiJFSebLFQ4eBZEKxPOzKx
fwUd91vIbXJKFlJb5RLBiIWi4LVfyKoI86z6Rjwofg7H2CzCRZZ6NFizxIX3mciFJTh5xLx3NpGk
Zf/9E/5XGVFRO1ZZjErp8N5CsyBHzdzdQ8XkNzDwzt2H6P68NyW4sFV2ShHDzaR1vPrYscp3ddHj
P1faQWpxGfZfyt8SgjaAJuoIn6w881ZO/y5gp5/agSqNHWthre2vxbBqz4sL41CQz8A6NUaBg5hs
3e5iw7UFm4HMAiQKEVmmciOPhGa1zYzLLGfEEPOu1RZr+vJs8kXRZsPYQ0JuC0ZNDFvBtpPgOXZX
1QIqtQ4owTpv5FddSweJKLUeyfLMnsagz+ADZhZdnC8ouyyGsprs8+HXqbtYThidVtSbH2sMgVAX
rHVf6VGKuVMTmkP2vau5GlyH9Io5yHk3m9VzxgMXz2TW7nFNK8affKGU6McELlJnzCZPwIMzdbGW
9bh6aeOJn1iWTVSnWJdzsC68HD3LMvcl2X9nzNPiJ8z5G5WW0pakVWH+wOPcs1uDuj7krL0DmdPS
NtJLDoUiOVq4uBK+de5UdbatvoeZbHNOX0+1j8/79NuPXHHi3BmqZLYXmFoTKST2l42ynQt+qT/E
4OJHAs7tImY587ygbbb06ReKhsYd1OohS73U5yysUhlPKUmQUaHUNRmfYrPT1Ntb5GNw3zbyPiMC
v6qpMCZZmfy22yM2wJWPVmILLbGwxIQe69R6t0jLmYZ0Rs1F/wWmZYZ5odHcuqmcpkLzMRw28+6T
i9ObXlMQ3bs1CEVPLR/3eXdRh/Mr23iZlwG/D5is5oZ7HgZ/jyUhIcCOR0sjZvU28H5nuLMZmI1l
4XxkcJXW0YARwxobCO5gSQgAotAVD6n9oHebWDUBvysqy1zSmmHY4Jlst6UBGTpIXlPJgnGHdIQo
OOkDZWIs2xafLa2q7JVHeoW7mL/POrlvoInKugc1t3bWpWxXSa1xVet7jfFEsIgKofsSX8qYZEVU
madkyOIn4vRG2MV+9C0WP43ZBt/epIr0gaWCXlCiauCrFSNFsVhirlGZW490mEheHgdQrHD8AwFJ
1Y8cNPpdYEIS5dlpB+ZofS8Fy3goittG5ZhXCYo6aOBKvAWFGduXkIEwDzmchk/wMp2F6yNRJGKZ
OgYNGXcp1JrpZleBdmzZMd8ojC5W7jfVlAdvqmZzTmojcUU1RwxhMf3nfPGrdHGqIJ0SQ5DqCDc9
tNdAZ6zjQ2lTrkSlZxOFEv1dvFM2Z6lFtSNeZs4YOzqFODjK9MNxSTN8zKPyvevcjcVGPWrk4maz
wQJI5EBwbpgdNrZeLR2uetdAYKG/+Bs+k2MX45ycPAk0av8CtezYEe6CPAtDeSpmW8/+Ie1sfdJ4
WWLIRxqD7MFLOl1KjjUebQSlAGXdauJ9bymU57hRaWNOU1A7nvtbfJkEC9WH2m9Ai076v2G4kDOi
mSetBELKVoJTLfyQ9C5clo/VzbzBceUvV/et8XupAJUYbH2yHqhruBcq1Yc56i8dzY/O97g8C5UW
DO1ot8uoB+2pAVnDRgOxNJuISzcoR5Lhdk1Fdm17rghgc5air37fou077+1ET1KFFPhpR+dd47bk
p0sdPWWx4tjTeIa0DdNA7CJ4HOpckanCGktIL1IEYMk5O22ZNPAlapVtzwLIGsaZMGb8stngObfl
U/CZNgCpYqq3g1RjjM+vVsd56yhimO2ZZjYxl/RaL/Ob5IirbmrNwqIiZT9kewJjVDdCpBoEpVt+
z6xoQ+/2xS3Jub8kLZBdZmemu7gb1T1DTXVuQD6w3qNq42EVEYi8Cc/nnAhv1xFjdohisiTT1T9U
iz7Hv7cQDPflw8e6wjhN+hZRBn/huIYSJMlXLPySuyZfK5kekOnGclFLlLQPbtaryIyeRlIP+Mnu
BPh90CvH4bg+GivvzYNxU3IgsWt+2dbM9U/N3Os/k/P1NR3Bv86EJEfz/XF8u5ggKjbgxnkIRJqV
PiE0xvApTIrlSTI0ejEaEHX1hxR478xdvFxOvuWL6UcKho1uINRsM/fN8eS2n55vdjrYcp21DpJ3
LXAuXxcgQbsn26bBtadu/aYkje8G7r2RMbGH90Dq0b6AJxaGjfoHXmARdZSq97m0Bu1CtFafE9iE
Qfh0+d0UBZEUId6ZPDaVIKLF2R3EU+C5jx5+4KWTIkay+c++XluRfgO6vsNt579xBTadq+/435ZI
4G2SlDI9Qxx1Oc2kB339sZUgTuJWnVqGHUeU/zGgWe98mIdL72O8SsGIWFTz7x4aW73dvTLeD8fR
msKkmrxoHboO+Q5vSKE2DuYhlynLGbUAEmEL9YtD2CilUUJVo1KnZueZ6YMOTi9ssW8qXXzFSeUC
okRM16kKo7KERK74x40xsTmLQNwsAFVcH74fS8zV1l/uB79jYGLqzSu94/0mVhLAL/LcLfLfvWCF
NCIi59xMHli1LM/5TS9fKJeM/f67hUqvquckRdQ5I0QqOEXNIqWZ2PDC6Iwuk2nGkjJYHwd637le
A3t+05Jktw7QBzPMPLd5njN7k/qPEtaLAPqOJ40zLa29rD3PNo1tnET+cFfBdITFErsZeEQuLO/y
hiLbkxR20N4XEZO2quYH8CkQB2FWTVBFSfwXIn8N57ucNt8UfWkGQvBrLhqKwjDBAmNlD060aSn7
Y9x2vHHlPfYxR5AT/tZn8vbNujyMhd5unaHfdjU50PJPXaKRnPp+Qei6W2wr61Obg/9Q/7SYPdXw
E1QbSc2aWUjHidH90VTigXo17P0d3lkfrp6EnngfUmg2hcZSvodF1ZjUAFXQF4Vpdsxev8Xa8Uxh
ievElosuJiULr9GWvaEXEIZG0NmWSroHy7GeRe2LrOtf2sb5TIupWd3FhaXQAi4uqRDjExJM3SHt
h7D5Yk1+HXR+/b0XZ0G+TNxk1DSUDBmcunxJrtBlJ6uIiYCWA3/WB/IKs0d6Qb5MS4CTbLUXLZ5r
v/XWgj+UHIT4UPJQLYykAs1/Ij8t3rENM3jm/LvSHIedLDxklCrN8EGeZ11uXjD756D+LskTnk3i
VsjDOS19BQMufNQ9QSFMzRfFNdYVvxFwKeeOsnOO56sRcoMWsMQkiuQl3GAwpE1jJP53Fzneqycu
Itqr0m79NhOVBY2brUVq4v7Pny4BLfUaZQw2rm1hM5aFYsGrec11Qc6mmeU78Iaj5+Ps0J6zECea
PdvUjRrTyWFqZH8JDw3EiGkqqY/G8lC46CnhbVFUeXEEs8eb6PPWQ9aUhiEcRte75fau0X9hIxOd
g5qSEoXTzYi6fAnbUXpB+33PCgaj4yMRESeKrFsMOJ3P0ms3CbhGxfB9W+bOBOr0ARtnqxCGIsBr
BFaryA19EGwU031NSt0/WX5Lbk4rRM6TYBCGxGufMW3Q+22tS2hHhS3pebKDms3ZNnt5gDGhf5nC
Y1EKK6zBvcOEdOnnMsamkbTUrdXaEfxBL66dpVwfM3KntLKaa1AaCo1PnxL1ujoAJpGsR7JJaa6G
9+U7wnOuubB3XAkCKWm4yFUBLIeBSAvYmEXUIzkJfT5dTMA1r8uxq+aP2rzFth+dFPVwpUNcp1ue
Dt2HG0ZAv+wIqNvffeJ3A78t2/VogR/MJJDAZKdJ0Nn/jE7aXfBDXruZ7+rQ5p2b9EK2pqqjOBqZ
71jfTZzdhO0kRh3UIzBLdjUBwP7HskTWTou0DuRm8i+VFScR4Z6e5HPU8JSC08PTNo3fJS3otVXu
u4KSuBMMPqLj6qrmXkwCmdr6gpUNEE6Pb4GtQnejO4hY0GMu7atGpqBMvPxqYA7LuENaQGPyL5+C
hy32eaL/F/e6EQ88Fcn+uRGqqPrXmB5VvKoE59/dmFLaBqnv8oarKnshKCBNcK+t9cK4aPDVZhBL
Zg6coJUf7rmx2p4ckA3wmaKEBuqu4apkb49l2u4rOTPBfesXC6e5gLwU2U57SWGph/nobCccEUBK
CF3L08UlJfFOja+bNdyg3vzUPziCcKj6p25p9Fh1hQ6USP5KVLKlwrrreMzf6J6OnGovQcq5YzXM
fpzPGNovW3hON6EtgwnjqHiTD202h7VzPKNwagQ3Qv2fL4DRl5TN5tFOe6GBdhjjsp+3cNkyrqaB
tpYcyJbqpnix5syKgSv1rhibiYR6czr5N5wq5YuhPMcAEfTpXzBgdRE70BGNBt3QlKOH9KH/Fq6y
Otiicbq2aNJlmGIGn85RvKUfnsNCMS1fQj2MCiPZPObljNjA3UqRH5fvAnclr6k8VOm+a/9kGjtJ
p39HwwqFCMlJAdCxVggnyW680Pk+XQujITkAOCu3LYUq/QMwym/NzKqMsBNmlbq72czrm+/J7KeG
+ov902vBjWzB5R6Z3tM2jiuYqg5zC3hlxK3UX8REDASVxzpvoPBkl7ak5WCtJXZwNkiPCPe0nbb2
FdEa1rXGoeP/NfvDlZxcacOQw6SeL36u/6Z3GRws2uklPTq+fAczrcxmv6dV+EdMFL+w0U1rKwO2
FSiLTZyLZzKIciKQkoUR5tUYMidjn3ybvOa0YloUtppZ4sCad1q8dljclmMasq65iIVl6I6GDPca
9tcNUDl+WFews1AfMxkC49jUu7mq/K3tShTifDEStVTdY8L3eJOkxCJYFIQ9GjRm/bk6kR6Vzemj
ICMIgbHqlht6C/QRj7wRHOaEOYWOFQs7BdMQC+tnzOj4xE3W7hMHCgk4w1VVri1rg5Wisk+t4hv9
JO7E7HIWcgR26XgHRIluGFZILhsm8kBQShs0rKeoYxdYDYU1MWGZ7kU1hYwcyNZQJJfjkQIuRTR6
dtNpWvRKirkmh0EGhrsYnmLS8+4FfvSTnLQFdShNJJJtyF5tazBdzGkDKicHu7sjLMd0UgR6M7dQ
Pe8tSLKKj/y9D0VODRBrL6w7JhGcEbr2AzoGFoBXWCAp/dcxPXKVl+oDX5vB5lUVkzmfaQW2fCJd
nIVtfBVm4yQPRkxWQEdb4iylBkorharP8JqR/b+4OJT3iLMjezUc9OYPWMu4qrSuQ2mr62ebx0eo
O/zI9pOj7spm1bwDi85Vlj/ltbiomE4TGbToJ+9qZ7hcukHGSa7UnSxzga2CZLzuW/OkVpINNZkb
y2WHEsAZpckgO07+9VxpJFtqihfGQpTFqQDcta/vADr3W+nsb31OKyEfP+H10I5/xIx3VWs71qQt
FfvBXkEj93Il2fFdCchk0dC6379cSCIXDmjQNlz+5lv+DiM2JNzS0eD+xmWLoDtIqQyC1bwjh9TN
3Xk48FgEVplFKRNlQPLdinrq3If/69HAScp4KGXudHnOBWsoEvuRep8Hm/oCIlv18kbnc+b+P5gB
003DS0R22VkrWQFdTj7IN2Q04mFKJe/Z+c3+Qe1eLQmoW5zcEd1FYq6dQZsPf3L8kZkTiXZh/TqB
Yq66R3pELmOtAh++jlnwP4f0FG/5+DXmeP5c1o6bRFIej39Whfoo8Bo3TbtiA0TeoMMNcPpJmNnU
HnhQtfvgVIaF6YJu2YbVSa8sH52TL7j2HOTmjkV/h2Y9YYJ5ZE5VGLVwBAgg0gUSIfWIAnUnZAgb
ABB3qiA5244JfcDj1ryONmqYNpHoSX7OPj/qRBitptGomj3Hw6sUDMiKvuwEbSVN7D8Cb3N8te9k
lqcJrEdLGQoKzDsuTKGvo9z1V1ewPWYyjJOr9YuqNykeG0nk7ZKTJgTCHFi9hcmTo9+tGM1QS++5
denNJt70nbe3nnW3ZVlUPom/KQdAv4C2CIdt9KQAumUquGqR9nuwt/tBqlzmNCe+uwb01FvXBLfY
8/2EsA3dUljgd8pxW6exXmlz7J+08kNMUpYq77BopOJvRfOVV9/JjxuwPaxnyhpqnpR7CWRCDKiZ
1gC97bDvdLEsVgUaKbm2Xt3u71tNj/Xa+UD/CSEnvTvNRnmQ18EaQ6nn5dvoSLTIFN/pUcVcF4Uv
rc+p+fY4upZdyEKb1TXUTRNjoKqUkboPWm9xTsBSk7WK3mFBl02sD+iuJ3xfh0RMOVSTMxWwx0h1
bsz7ld3BCfmXOT7fXjyfIztdVYfAYF5PvcWKvzuGbjouwjceQMMDVAazgAmhbHyNbQRkF/VMsWJh
f2d+jnD203F+XnnL2lioXmjeTzZFsTrgRpXKKo+0Db65Ytzea+K6Q91RYE9T3Utjl958cLFyID2I
p6oUg/NQpIKjnNsneP2sZPqC8nKDnnfaJ+15LY3DOcSmWYFXzDMolczmQhFy6QG1eBAGxzfqjNFK
F5x5E036VCXcNYfuAAfdEiSe0qRf0DS+gcCDTl2H+nUQvRAMHEY870NlE/KzcOVwLxNqR5IebYmN
5icPnfZy1cz3dXpQmHu6LFEj0bytckKIK4VpfA0uFkjQgT58AgfA8hCec2Z4NTqBnHwVOBRz56/F
xDMgVcJPytDsGvXjfVSPiE/gM6IxCw+PZgBxL2MTuRwBtYKLZlTBjV4E9p9dTzg9/xSXFkGhZPF9
r3AJsbbvzBpsIL4xaGf0c0CBrzSx3hJVh1QdOR6onshZFej8Zu44/3mwW+vsdU9bFxHD/cJgdZbU
E9uwCjDK5TUosVl0YLPDPvsWzzEm3hL46vnVI5pRxiADj4M7Og5IcNBFdZOqZu+Lsw8uJfseh1hM
yTUt/b/fTxMSJbyL6vPKQHUxG7etxNCuA4GKB+XRDSr83R8oXLm1QOSm2eA1j6qvP9YfDAmLMKBa
REvgVu82n5pccEa4dyGtMhdy0l06mROKferKn4HPb8qLodZxK/TAYJyX0Pbo/QFnB0UKAJy5JAa5
9yvk8obTTc57I8ljiKnduIgvX0MWhNsuKeAj4p/XIz4/82ATIAMas2fUWHZPbBePAURg0+0T7REe
n8ehgrPMFm8tLwN4OIwXT0ET9NdLhVduOmZHump88dzDWuPL9rdqO9nFkCVnXbgUd4qbzALUHWLO
H6dWy/btVhelrVK+1U05PYi6LWTemS8P7R/eZga5fBdqwjTwE4I1bY/lCqSVurr73QXazVY7wczt
+ZnIDCuGXWToTXlcEUaCsvXC9dcfuikIf2eoq0uqo03Qx/B7FSTe4D/oCJkk/BMAHeH1/L9gPaK1
wKFE0kVofLN2CCalBqWKACOtnh1R+Iq2VBWAJpRZDUy5JG4aNix5oI1kKYluggqXKkiReiicQ+HB
mUIIWHl/kVoddHokaEuZfgcvwJEhq357Fus3mnz/Ltt2la0MF4gmtd1rueRxtkAPOBxwvS2n2WMF
rlhuBBDUZkx8myODFgaRfe9l3MPT32l7Nm2G+WCE4DZxNdDI9ab3JyOnhbBb4YUbFqcNF7E1F1wk
vJt0tYiXTcCxXuwbsbtdiARQx8sU80gt2xpC1zvT0WV9upM2qJS+EK+VvaRwJC38GhIz7+qDuHtf
gMn0/C5uzDPes2vm8FhngmM+gcbOU6dV99kPhTmmRQSaoH5WQs8I8hFegSI+lvG+qolV/pyLffSv
eGMJpxYMLY7pjsyiiKsbvAHuu9JIi9HY3Kk1WSAa+IkQmZT0QvkgW3Ku1U7mtcpYHcAqtFABUCXT
Mb4FQxEAELE040Oj0mizCL0AkPK5iu5U4nKTJaVvmB510fnonqenMe/MBx5VEgJngegTu4IHWurZ
ujKfAo6FU2zjx0je2dns62vvgQwAThOFv23LCtCngPTgbrXmrKaOhP8hw3iicnHZ4qSYLidztiwj
OH5NDpN7dx7fkYKuNfGwk0+qlXIDoZNm+uxDmM7NCEJOJhdJPHLPsJlf23+T5zRqB/JO3QndOy5a
l5YFcval+Q3wsZkC224bJBAFYqP+VT662EIAfvaZtSciSFLJH2hPebWKyAcYLLq+wa10kw8Pbqv9
E+ursOgkI2nwmilMMs0O0Fy1qaCr2KVKLnF6k2QA2Y3UZHbh6HmXVf1uYyWp65B2Xe37hucP777C
OXMmJkfghHJgKMMwuH/BwlXdUKly24a+O7mQAyF9HQWOrPhHlTCLV+wT32z9s0CeLbEuJNN5lN9y
i+KGehalWhrMwPelM+Z2XZBWPUMSHqHGlVk4xfdRwdMkayrVcctY8CgzglRFBU2k031HnehBjMtX
Ug7rf1Z6rkbe4FDoQJQm1QG4SJT8Eq4kSw+u2bYVXQdBS+uTTdCiCwDU4bB4M2H0Dqp/+CsIMehM
XtpDkbi4nXGG6nD/BlQl30VHiuzMJ08PXHhSi+HRSmILHxcmksx6NLH0ynYbnHNNTnHj4soxPNBU
3bq88Sc7sepR/GgxxmaTtGDNM6oFhNm2BnEobJsKiUA53Hxa8DLHBHz9HVDwGN4p+5JwTAmSIyTN
h2bMdoa/Q4K/HeKSOMoNWodNGW3nbe97850XJn5J1Gwk2EOXCYAyj411HcFvqCd5XlY/P+uwIgSI
bnvbDuZC5Ovw8AZIWSATnZrVuXUnA31b4jMvPTeYfA9Kg0BkDZqIKUm2Lo7ys+969H1Y+5L9vNLg
qUYA/i5jT5jTGiSRCc64bi+ajA7cvKyhNcSl/vC1uqagHMD0ckoHRPgblfke4P8s9KWBW46YPrlP
wx06OEgqfGQ5uTGUItrGloOkVMAhrq8axkMyGITQp1FbwPHYBdxBcjsg65OQWtlU+Y+3jOnhpztj
4J6AyBP08hngpVV7QPIe3DY/2nA5tKSxK4ccHxtWl8hSjTU6QzLwaonyCWKfchZlfVSLkUnrSpJD
znRM3EG93eV4Txjt8jcXDOyopjck2zE97q+mjWomGkpDqx7P86lypQkNClJm9ANsf9gSbaJiR/tq
OU79Ol0nPScOtNlunS5dU0g8Y5IX5hKBGRqsPEGaYgSZxjuMZDtE1uOlGwxs4x86YvyX5Ymsx67/
QZh3acX+Ma7Mx/5J7PsEPcz6/RVYuxX96VXKV6aIQrtmzAuGZBe/4wzrayzAYv6uDfJVaSmznDUt
08sHWc3SfC4fQ/uLusjcMl2mFNR3REqFsFcs1iUyTp12wm/T5uD+YDLmJrsV/ql1dLzM27HZYy56
zyiMOWZiOr53px88n+T00oLyyFiFIHhm9QaO4sOJKTdOM3DV3LqcMytrqEVAN+MqHC4G+i49QsXH
/4YrJU26VtK7rCeWY0jRZzfaXTBopryTkZmbpDgAO05MWR7iSAeHP7gFCnVvGvFv6ifISSSuqYiK
C4NnHXufEO2A5XLo08KQ5C70TMSP2pVEqnC8iaKRj6LZjuwvmAmvvCL+Ah7WxLi4Cm94DZY2lCTZ
LxT5pVA4qs8c3PTCzE71HzNdLQLa3TX7r0k4P8oQZH/SugGqiKxdTfrdP7+5zGrLJkrjcjIzrnLY
uyKnHuoKZQyC9g+MW7bwgJL9aJibG0iSwjAaVxZr9KUkmOzp+mbptgBe07jl8HMj93ZfHQRrKZxm
cuAkCkr6D7YRwR6mDpvBlcpEiJEEZUp6rrFBwnrfqkzAklgaQWTr6wkDZ3tDdLZY66vVpRCprHRx
Ix389+7bNuh00WLQyAEOhQ6Pres2j+e12SeMVKN92lmPenh7isqwMie3mMTSdN3RCzELcDrcziMC
EdnstDDrk5ygtJM8UlEwlldvzrEqGzWz41Izntk1zAD2a0kWl3WAGxWTMMhWlhJllOVESMSx2VQ8
jrlSbMVEIdHM/sNI9+1lGbSpnrG2depWWP5ynPhryrkWP3Cw2kWb9LxnllxUg+stBZKIkBy0ztzp
iJVSwz/USsKalRGhHPtq/AGwXWDIy9ypEGQLVARbOC6cyovHOYSJuPUF1OvNdzKk/L03CSWCoRBi
vUM+wdAFyWmJf1HF4R8jGWriOqkBtGKPRbc/dnLC551zoSrQnTvV1K9hYFMAG3+SLMXqzWshprIz
oMhP9+xJ+NDE5bAXpr31F4WENbs/W+LGrI9z4g+n7eVTDe+y+BszTf1m/oOvv1bSFRCB2IkOu+Is
W4p4BB7g9IKzSVVu6dzJsDQB5n9gCvnv7b+RT5Ia8FBn/DhH+tvV3RyGK7/5uIJfDfdKIB8N2MuS
1yRjmInxoPO/swDdAF0LRgRKIX+pv4SXncOEGSKhSYnQ/m79Z5PvPx0whNocsZAY/vlm1Ofatn+F
HR17iM61AYXc0hqQoxpJtWbc7olM6DngogpFBy7rKdNUXV8S/qs0A0zPLmiCwk2U/VxTu9pkE3GC
j8Tr1bOyayndDAHc3dHbtj2+DtxhpbMMzv0j8+qOPXHijBPI2+5j1c1Zujb6cCftQYuseFv6UDVc
JtfF+EfBrvEWg/2gDpCN1NUaKBMmFbP3up7tKUd3XA3jvy85xgmc4hvPgxFo4jC3gNYNkoFScbUR
dpDJuNwahbHvqwMbbeU3C8EELBXrQyyhKDLtf6COXzd1UjO1BUIlKKHSsLJwhU4wIPlqDrz8BocU
I/b0H57hKYiZou4s0APES8zhm6ZP49mSfQCM9oG4zs6X69jPcAvXWLYoBqdGGJ2R8zJZngMITqmQ
my1DnQ6k9gQCReCCao91L7Om+ZP3RE9D0YX+cO69mFGI9oIpgIl9SCsL9AvbCsUZxrJFxtAFdIPc
Hn4nqnHG1CJbx1vLJ7vudV78qmo+IkgfVBig4fF3w/HROQ3XkNvOrVQsY1iFen1lEps9pso42AUL
VUpr4uHDo6BWB5mXgHMCY7IY0rniOy1y9is22XOY3QKYKZCPuTzGnv6jZ5UjfaoqWwZ6dqNfe2o7
EL2TuP1MeautdKjg2SvOL5vkm+S2zZYPA5HXTnZcWEvHeVmhDOXrgB3WdjPsrm6wCCI8bTCfed8F
i40zpZAT0157h5IgCGSYHzLARVPbuPmw/w/Zb2xE3Ra4Mi/x8yX8eSAMQy9PpV4Jg+PvTr4/0PEz
BpK4xb6gb2igd3QkXYUQnIsQS6ZBYcCIFQ0AazKpdI8avflyy7cfWNB8XOffHD6ewTBIYPbMX6R+
B6TSPCzFKB2Z7op24Ucqk2HqAq6voMMdEsLHjRH1Z35G5SI3+vIHloidHhcmq/UyiCM0F+keJyfR
q8rPPR/nL9R3X2dQJxbr0Bf/McpPzbv6resYu35MIjMVUA49DN1HCyQvCwUpmL0HsHJOmyiqLOEk
pdQhfUbw+UoqnJMorn3eDpPG2CwsPiSvW4EP9FrlwbwnF+ZGrOrD1IAIifgVcoEuY/4DkfRKxauD
35zz6O9uAIQNDVDCdFbPShbs3NsUHtYXBfi7AFN13u0ShnRxjCmAieAhzEOZo+TOkcyBRnD2083p
R/xRjb8Fp1SSB+Wf/VWo0tUqIhunDGQFuINZyqRJw6UG96jUjYVFVyBo3MtMVbZNo5DCwTVhVgaM
bSI3gHwTh6TgawSyN4QoQhDfaadWyKQSKoEFVdah6VfgWzHnyI3pjUfQvR2ng0ByBM6PsZ7pJ+w8
IcUCtaEzZGmB3/9/nbRHSGv35AhI4Da2x5iSLqzsSZ+STY6y5tezvFzEtaqyaxiFe1HwW1msVCIR
L4zcirDI0nWFnjlfvqblWpeoxh4LpPM7svYYBzpSe2yTkhc/O7wooeTV/oeu0tGIV9XPnVOj47/H
SsR+B2EC8Gx9sf6a++iPQNXhIrVdrb2k5QVw2plv8jJDlSQwitsW7LiysuWLeAthealdiUiFLo1Q
gK42Zwq6aCQK+fL5ljyzuds87ayeYwmQZE6IrGMv4OajUIX7Jecu9T70qWutjKhhWz1Ov9tgoYJd
gP6U1PncTbs/4sRfW7k+xCC2aTs7OzQT+4AHVWPZ16+i9enTA7LZeYXkEvYC+V9pDC+ukY7luQT+
o8iB+Cy43QDT9TMqj17aOfj3NqZxOdG18zDH6KNBnyzDHDCwTVwl/GFh8Str8ggbJ5nMlO0USO37
k+Gp+pXtLAKuwqI9gBQjKfOHABOuBTkKH+EtYm2/rIB9SjvlSQuGUfK8cobNdHS1tLL99vUr1t3m
KEUNAECb7FadnpILn7axiEht+sw/iclzcv8EFDr2qidL3rXMfXSPDgiYrH49i1ZL/GPUL5WPAMNX
ESWW+Ukjfjnu19+RlM9O7qFzrDx6nk1Fk9CrbLPu/kSVzOUjJxYX7tLInkN/7hXtlZMObh/f3L/x
kmOWfLKqzCtWCQyX7K7TofvxpzdCz0VpB1+Ta1gwmgl3CiscbOgl7Nq3wojmUvP2bXotbGhdnfNI
fejeP7eAgdgUC5XWIfITwA1nTIFK1jKIlx345tu0drrAt1XqCn3KV/d9iRYY49INw1tegzuhlMwo
mlmPOHoEOx1Rl0peqTwVXw5CyRHGZA0l/SabsUONbij1r9bU6a/LrrjzeNm/vI4aC+EFWkrBJY+t
N0pJNYOaKBxcd+iqwyClXiUxIFHUFL6zSXzH1I19h+taK/Gh4vyJlJJAz09CndGsVQDccVMabSZg
4BPiu/Hznecmf2jsy7U3B869fWIwesnmLlwASMVBuzit/Mz76S/1sdpx91zt7ynPpSS9KntbUkwK
9zYmAVDOEPFOlTERFGNabt8Ecw2S4+Lt9dgbIWrpTbMe4jq/EMTKdhfGX3311IZgVGBT+Ta5ECsR
BKnVZj8NZpVYmQUs4OZOVp6U5JizjaiRSmhzK4Om5rNrXqgOWoCdo3YDWwTfFW02t3w/J1ptwti2
Ij6kqJhEFSvSLeoM5hFUbi/lhEOekNGaRhWpPZKu0HnNLunPrQeo5zGGFPgr/dzkgH70d815WI67
CJOS23s7DrDdA/QXNkUBXxjwdj877PXiLS9kHRaMu43KGYKHtwnNIoi7Ib8QXz5OcI3ccCYMstX4
BzDXsvuXD+JjkwfauPcFuCnEPaYQRl/Cu8rahXde0QDA0m3DMo66dqPWzLlP2XQuW1Sw4gRRnVwt
GJAp0jWodw4CZ+TX0yW22jvDulE0RK+thSm4wJq7oYiR53MwOsU76l/Kc2/wyfK+KJ9jA/NOcZ2A
E/kxocw0HMT2gFqjDjaBEBg2hgrx0maKDlV/R8VJMqMMIKH7EXlsA7Ncgk7/VJn00GujeintK0qX
WdqaQWj4n4msV2pzqAAtSSPxz60hLghqXlN3nUBmD/g9uL1nDG7rVNZovY9vb5MIgPmFood2MpNR
HeZ/+3bTJ6dQ0+BNXszBSnWQKs3rn+S7AOkdkmJPWuixA+MTrzY5Z256DL9h/v9LwKdw+gWvYuKK
3wIySWUb9ZPoFm5Vn/QLMah/R+jCL/OpXaaiXT86hljtWicO5sPWGoKGddCkEJPwWAId2422fwZx
qZjujFrTi1btjo4CEo0wO2i4vaZgsPNzIQ2p3XOj3yp1/qjZYwWOgy3pRIo4et9sNYz48UEVGeFJ
THQUzdILpwU+8OJB0JkGQEA6m9NiCggJGFY39umxymb1rdv3W8nTyNjN1q7RQ9Q6IWCbJPjdsDuY
iI8XEs9I6AXE1igJJMW8LH9jGIeWQGbVKfstEmVTI88o1rV+WTaZR2+C+6otXjX8/l3GnJtg+s7/
MrVsFTkvoZqiTBB2X8kColdmXom1gnokVjBCWn7MoSfUqekK2+YDBklZvcwSfpZ88G301Lq/qneL
i9j6cV8Ci3ZTCT3SNHFyMedvBQk1S5brydGfGRRCPOOSAzOB1l8fPj6ut3ry6zOUOJAeG9f72J+q
3W5EYxj8n3MnWHkI6URIedpaWLKqve9Lvc18+Se15+ScK7Zm5LeakHNYA5vppCPlzS6EzQPoIPOl
wkZBKw75xLKxqGnkJKdVEJb+/4NUO+4ueTZOkhkfNR0qGHql8tSx5YSw8U+jZRNJFKlNvX/kqcmP
TdO3lOEBDWoWXfZWrlwKcty4v5PBpvN371Z5EfVlGguT5ezLq8gmfzLse/ImkkS3yZ23yWdfwrup
Z2W7QZeufKpPz9JqtkmPz3lnmShTHLHxcCmpkX2Zv4VGzB0Edf0DMVvTPBFC4HmOqBLCGWAvnZX+
98S1jprV036/cWpsB4W//iYPZMCsWs+e1cGCZtXonlmfijw/INiMpCE1TWORqP27U2uOJLF+p2BN
QguDkWU9qns4aHtIUCOJ3D5xiz33ioc7JqYOpjfAYmJeD98lv4eLcEOsD2rEKRNXr6OIzlsLYtzj
dRkCcUr9TWPLdBRJqMhjgoOLS1hWm6wk8+jLpUOwsQBzihf3iB4DRNlMWtQSQf6FxWrtaR+bDEsl
1cTYwv36x8oE79oC8Ixmx/7PfRbPKrGCQH22+efAWudUJQTSORuV9jNa5JAulIC7ui3aubInEfnp
133bszlAd7ZsHOr8LCl+ApLXHFWq9n6cgI9eolM3cok0gipvrRlFb5zjSNa4Y3SSZOWUq274337O
j1qBcwXMLArlen9eQLPi5zv3VvGzgrOUjibHy5P8xklFRqRc4FE4gpMBtEaciMRzbz7MfB4nEK9J
2AbfTMPvaxeR9Lzhj+b9F07mcJ9MbiZhDJuTmWu5RnWtHdqbCUiJZL7AIEKvf1MGY4Mj9yTMwW7f
PM59Kr1SAwyDIkskpe1HeHdFsAqYCjoWaB1b5DRrUx0/MnQAFVygCCKR6vobW7YVkAj0zNvrR+vy
MAx9iow9BP9tOX5AFJCfxArKUKeMFZtIeVKa7Ob8tV7Ta8FdYJep1FJTGeao5nnzZSyWZSk0Q1HX
nNg18o0/r4XJjvSpErtZxI3bXjStPARIofxhkIHshKs4jR8uraQvzgod9jkoY+TYNoQkiZLmktof
Sj/uYAoVapqP736HF4g++f2UJG0ZRWWVcQ0FGd+ToK8gcyk86vYVogIpbj7gbT4PZDXgNMpp3Vry
ns2HbkhkPe7+Rxme/I/YZ8Fzaegn+cmve730F5VX6LA+ppNB7DhDp9uWZM9+kt0FQazU2ngPS5F5
W+AJ+c899HbBddVBfDTXxbqMTIWQlYwZKwVU31k12I3xzu8IEaUSzz5AaZaY3YwtSyBgn2p+P7lu
OuyiMuhVWOuMBLjldp0O/nFTA3VTzWsOO5I9FaPniBrcpEZRVUzKQQkbm22d4aYbwXdLebYnPr0j
opPIxycxIkS0zZn2GbJ93z3DMs6g0sQyQeBzQXu9GFMfEx+bK+IPEwtullUMEDE2PElf0SJ6ytvI
Xx3nHwM6i6EZKr6W1SU50qyQqOe5lMbFHacQD3u+Gfuhp78Z9aFuqF56FCuhOzeD9jbZOi+r6slq
olHl3SOKdXjBpeLZH4Yf7vK14m6YV+Kfa/R2lGwHqGkYhfB2g/UCr4JP8arHtaiQArcJTZE2OJRs
vzsQclPv7nH4RmAbCCNX8lLmB/YryLbMrSIOqPTn2y6LAc4z3fG4enrIdxnkdSFzdcXEL+GXq9BK
TX9CtZsXxeUhKjAscAvbCSRMOa2qYcE2dpqbD8ofXgksuTjvNKz8gumyrpOROD5Wyvx8AQEhaA9w
hpMz6QhkCnYS3ZlDzEWfexLGA7k8pHQOwPsRsnwRTqiTNgVjhzu6+++rSc1sGaY0ufCZGeZmLdIi
K181rI0lQjfhfKZ3XVDlGhGXnKdolAbfNuW/jlbsQiLF5+W+KPpeywcBDmAIzrUlGs7051UFMZ4d
mPIsGFBVfdVkwebmaQ7x+rZoVd3kcLbZiocNja1K5ObaYWyuaLbm6pAsYNDt/0MUuQdNRcUPfCJD
jlz54YXZlqG4FkcwIwku6R+4jbVbXY3Eu4qFUn4ogKsd9boFxTjBXhS2AlYN3Bed2b80cGIniBdp
Ph+P61eVqAzAIa0NGJrNNnmmx11nNBcjhEcbivHVSXG+7rUMORuGfkKI/JHuEnbhN/scaOztRgkL
XgXgdsLlU1usmt+xo7rxpaLqgKrX1qISNX8eS42isSmbw5cfsLvwVLVS5AxKdlrym+YkKSc2lh7s
lvhjrZO7YDr/5WlB69CJ/q/5n/khqjgwXBWNDx2cS/3ni5YEtaMWUKSraLztuaGnfIvIdn7wuks7
FREsAldI5s16tyYDH096UU1gyPw8SfVTyUyZyuV/a1gzhAivm7ZT4YzL+W9PVhHstK1L1ct12Fkm
cBrdmoUJayq+y9X9JEYNgKJdV6SOjOCsLbrJH9rJeqo34GvOVNPCMr/YuZeVjl+lhsT+ONTZ2vgp
HVVhwr6gbgUbPWkE6m95fNsEdJbsCxcSiDYX+I9ZDA+JM7Au/GkoM1zsr0oXVy7ey5VKHxdpzQGs
oAV0/YWyw72cHxtIdz9yIUVFyaFn+GzEit9Vs7hKwHo4g9PdC/LkNWHP9Zq/bMVviBUwTBgY1K+p
VmJ57xU0NsYpzORVsEdqntZuOfuGwMVub6TM3WueFv6VyQtIFwBw7YwjTZT6oxx38xF2n1v99eHy
2zyvd57EQvIBmWxflJX/2NLdDFJ4GxcSuxycZdKSoB9stIkUm72oFAU4pfEhY7pP7kNiG0LNjZ+6
Vxd0+/lPdy/QwDhXkw6g3m7hFRetOb+SszUWHQTjLsoJFwG1yUiYvDvIzpcPKlsFKrAfSpGw4e2b
xQ45VkP46EmIIkA/E96p1ANN7MKdGrbm6+36eJ/Kx+SRV+SVnRuSwkI7sOHI0PRh8SBzgnUhpPBB
GtpNTf+qlf4XF6tvwcXNiZ8aJnq7FyQFl0hqa5mkLsHyBn63CjlU16RIG9Cp2owTNAbewyeE7y0p
rLQvlRLZ1SMWdRj/3ipi4JqC93wTRMB+kUNTXMloy1BYyb+34pDfCIC9JusDdtX0biwvhxvnvEnm
M/+1FTzJzR11EF5E2fVBXIVcyd53EB+w7LBLiIPPwr9VONg+1e8d8WghKet2yHzDqouDTlzzoVd2
U678g5ERlPw8hq9oPOWczU6W0SSEu4VIHeCS5Rp0oAsPF8B/SFNAMSA3E0WMpZlMvxLra8+BH+8q
sRkioH+8YAFXs9jGltFkMtyy+/ICI7KDGPya3sZt8WfyMz9CogoE7arKGhmKI71OJQWcQUOK4kAi
h0qRTc1VQlI/jjSb9gAja3CYNEPVFv+LD7zV3/7GFFpHgYTnpMXeGzwIMtbeZ16hWPR0GkZOqmnd
UZT/tkgCzxu6uHZQeQbTWLdVxIG0o9YnjNtuOHCyUhzmyCVFD1lSSIHoy6Ns1PO4wFQy//Gb95TG
XvVRD/A/dZUHpg/P8vDLV5JibjX4p7lpLjRcbaPN1ayF8B546JL4mvEDdPkTI9aRLKavuHik4R3X
abrMZIyBpuD/UWnpE3QcxzOXNnTRMdydzmXWjd1ibyf8YH3MPCbpmZ7VKR6lG84weqdi6zL9FTuQ
SgwrO95aB1SQAemuKDkopiqjjJEdL2J5REjA6ZjFDJjxlFtX+F17MuX84vaLa4stlgxm615rnIpZ
D950RdCBdRWr05wofuUJsuZPD18w4gmszzJ5EUyJepbZfpJarQhI2B210EBmB77ZVq8dcDI/2CBT
kLmpd/AbGTh+Pp02ePuQLKjEqSZC/keemtS88/AOWsW91LsGfi8IRScAQYp853yneaP6mN9AS3PX
gL4KLJQoQfNaJ+e5UlxxWne/oMTu8Z/EKiGfjDiaTD4sTHSAHRfbNEpVNIqd1InTaluTet7nfNx7
i2lTkYVxZ5/FmAk7ikn6nboADibEgIl++R4KUyVqgGh4yL9UJWaSU+H8hd/0F74vNrdjcV3l7XA/
ZNZ6g6cYrVE57y/xKL7nrqtEYG4dOrWtJwQtUhA40sqiX50g5NWVrh8fAMeZOPl4J4wgcL901pux
lomu6RLs5aJUubFFzXf0idgazER5DmisG42R63S7noe2WoZOf3Vb63PenuGikm1bl0DYoKeE5DvI
3EfCaD0U7qaouMMoERgy2iYIF+oakBpYxeamlQeqb2GsjoQgIz7Vs+4LrrUIbNgz7qAd4nzP78Z8
4b/Jq+afawRb8m00tJMFghaGi2MiUpr5I1ZiDrrzx9IqVNFIN9CYXN3GxKByzcYGEW7t89I5A6L1
GiWvQG4JD8H0auxtJmiTW/KdvxTwyGa5GnyBvzsAHwlUB3WRUB1WQaJ0//+2Zh7HYrXMh1wTZSNv
APgKpPfWr1YREg5NKs7v2vvHkhtgK8FNJPjPo0vROEgA4razw4WcUiWFdBJ1HwC98zd9P+JqQ16E
ySN7jAedxxImzfcxj4U4B/PF6z0n7nwPWPbg/2UWQ7IckHGl93mMenxE2JfJkUVAhuks8bBCQ3st
+GX7QtzooBXV7zyqm5PzWEqajuvJfFrPRtnVx2lIcXZgxF+wv0bIKprHPC/4l7EDdL4Sb4xngD72
Ynt0dxKpEyQuLHzDKkhK8I5caKA4SqQyBIJEobCD5WjwftQ2RNVJDG2DKu+Y8fd0+2T47sQzyOU4
/f1G5N/BtJxUhUs+gWiBxUgacftmTEy6CIKy96UDG/6XOn77+YJK5m1PiR3355Of4N6FNP1oYwBv
UF9HKA8jbQUdVUl7KViYGQBqUUW434nj0DvxL9Q2yLPkKQ52RRRiRJX56s3WQCqXKMg47l6Wms2X
wBA6DnN+Tcfq9JpMKZNGFat6Ce8vqR+ASM+cbI9dp/TIGS2j8dY7wkFSqW9ZUN0uJM8QhGexqZkK
AZgjqYNGJk2YZ1e7qRXEaMc2b20CRS75/36mFBJirEvtSlPfbaO++wITXP7Ndw13XMM9P/BcReiK
UGq4SHht2dYSvz3WO+YK0lYfnAXOZEz9VTQ1vIds/WIcKGRknXJiTxW29FzVXGRI6bkOuZc+sg5y
+5r7P+rCGyhGF8ymdBi86tQO/9fgvgglZ69WovKkKfyBfKTx9Qyrdd9nc6szcVFq/7sxmUl4WF8t
VbzJZ20LqUpILJoSo1VUvooAdJKvvJEkIQ6fkU/ESl1RVUVZcvuJmoaiCPtqXxQShy00dJFlbOTs
Ef+jCEA6aqQffa2fZ9s1UQJZoR30qMuinZ4IWO1l/a6yik8wSiuOwmSALX4SjTkpNjzp5nMOxjT9
dENjhdQ++lS2GpfBBcNtQaUZgZK+JfqaG90hunNozX/GPL+Z1H5dF/LsPJsqkH4b6EcabQFCeoRg
pJJY7k1+jh+GP0sgmmaPYgj2nIJvzl7sm5vIkOUrFYXU6gZVRY3I7ThFq608eCg571ZizKIuCAbl
bhXhwxlp/9oz2U/DkHT2jNGs7muINjddM9zlgqIvaXk9CM/dvqyVXn5SKqPvLR+Qpe62axEL33T5
JqNXbL/7fYia7WCO3LBJEYoTEZbAqqf8b1rFd1d1OnSQ50OxjD75grKDalcaRSa3RWZIwXtVJzPo
L4SPTkJVM2OF2V3Z4AR01n7spwylBBY3Xr+xFx5TAcoPTr5aK3DoqEY84HuRTxWueDuQ621st+PZ
lMjKc3sJ3p3vnVnDqlti1mxFhrf6p6dOD1YX21c5GlJh2eKQMpGIFnCh2xGvdq3Uj94oNeCYh72Q
Juv10ORX6O55IFjjHRJfvaadrSm6LLx9W6ZyanBak1qgl5szVWE47LMF8BYnF2PJq39EMWMlPNsE
LIMCXtAJkJEzrzCzriRGD4S2OUWXGloUvcZXFjF/qsPw2XDSnqMVAGZdF//K4FAqFv7k77U+xHcC
j2dwlS+CtW6HdSxu0PocfowQpt+0NxGa6EYBygIP/TaIeuNYLiZtIUsls3IXtPlZ7sJAx9VoJPeF
MUUpe8tJKBEFH4GU2TfVt7hO5CFtyOnu0vfUNhX2bgkaG9ObQ0yFw5Q/J8yLeL7a31N1Vu7jeMfb
jGmLdTprWbsufSMBQgrRgn2K1R6Bfu+oA7wC491jDO0NnDiUd2VsdKVp0KMYNTT7se2ajuI2DHWf
PmJXTrLtcQaRaJ1PJ82Uyincwh3llll7VbCxcwBaXa7iJB4sry1VorlEyteVoM/XQg/wqTakvGHx
xLbZbkUItCns6tbECcrGVW1DyY01IfkMHFEZOzUn5KeAKvu0QdkJz254IxlgVvNllHExF828DVmF
9p42Qn83H8YUsopr/3vUt+/XnifIetzS4S9hBSCPajGLM++ggt9je7uRWnTvFzx5NsGJ7rOPqpJa
RCBGq/BQQ0Yk11cWaNxvwyPG/fHwlkWgT2bJDPf7e5114mvGkEN/7XCAQV04nPOF2NVxeH59Svjd
JPD419njBXzfvCjZtMM8amUPf0LjdRViyOfuwvA7buiB+eL1XADsyG9s9Y0DT3AMI+SSMInPqZAw
FxxY5BYWYuGeF93UeSeEGGjUHrEQL4GR5gt9pr+yK0QqMvnOYNVc8N3IZ3gbcDYVph8gEvjrojqZ
qQGa5xeFSs4+QAXyewSejMATNeAIkTzr2WrhGPjBUDT3h1+OExSkMrQBaU0sWvCdSCf6m5gH/fWp
HsOrwXga8dRvQtxDQXiQyutv317m3mX/92EO1rCIkyRq2JXgy0sCmApFD8x6byPpAWHKB9RiyUny
A0+8hPgIk6X5m5rpl1g7aFe7CACxfpdGWdBuGumRgoO6MZa/PCT0kRu8iliP8pFqYkih5/0TbY08
kACvwoGrCxk9E0h3qBg3jjYgqSyGp2ec2leXi5dNSWIO2TSoTpj+xINZUlJ+/fYBJyfDg/pkbzWC
VY4giOdvaT50GaELumIA4EdSyCHeBwUAyM8fPW6oz8W3p1Ct6gj3QYKQPT2kV+0iIDhDGBNA7+Jd
xJprd948Qg4ke7WU38gpB6th61+k+wEYalIrxtZpWjCRdGR4fV+wL3RANfJS/fXnxBnRztAN4KJy
J89IVdf9A3NZHJglOwwwK2l1qVttVbwEoXDUf7x9+0yIY1oaxSNWZyfet0NwhrCTDBVTr1yqKncu
1ykiQWOGTZ5n8AIU6O6MZsf/kHfRYii0fZwtV06uQG3PgFxvYc621tnMUsovGexcuFAXvXDtwvAN
JSECar9BVtaSWoL/cGfkdc/zomkCOThSKGYfoG9GaiITtpNO92XM94VYNHGJZHG6+ppj6NI7K4J5
eDayJbIGYMzYUgh/iq2dYP9kiI6JmGWPkARdAlJ2HrTphlthXiJ61hKTDP0mSeDIdBBmzt3snX9Y
k3ALqkWSuzDdPxGK1uov/21peadIh2yfh6DGBhysmlafPUISMs5nO6LFjU2EmliFbayED1hH0mn/
0vF/n9i7hiUjpfQci92ofdTsEhfJq6vrEgL1PzF1R5rTGX1LCQE2IcZaVCHF/dHax7O6SY+b0Ztx
ZXu/awtJyTAQaRvwfksDvgBmEPlhljJJ6/8EkvQX3J7oG1vADNU56UWKOkHgVzSo3l18tVHnOg7M
dJaDkpEk7jb+WQKYmDnB9xGrFL4PVy0WRe3MRBr0PyAMWL3w4GE36bpRtki1J2sKQJ9gEDpuEIqd
i/kwpbPSDgprQTCO/29TcKpzC5ZyBlnHXPbLcyBPNUMtemCAeqj0HQvajBwQZGWuJMQKrB+jGc91
0oOmzcM/kz4vuA3om9Lwik4fDBRUMc6g++GNFFJGRHM5JbyC8m3JSdef6aPrVfNGkUEcMoetIXvE
cahsPEnPUpJMIhE6itM9/8kO9Kpu4QrN6Lb3mNQQlg2UF5MJKut4pCOQn5rwdtie+Qxr4XmvcUsX
A+JIHs6emC7omwjb5p6KPzO18bmcCCWx6YF8RABXjLaikBkhstbcsjBbtvxQt5y2OHdB8pk5ghQ5
FrpFGBhPjxAG5qdbIyywdhcPzwx+chxYYfmIJJ/7zsoZftwV8zwdUhwXvAux1xG9sgfejMs+JZrk
HKnx3+Aovb7pyqGsxdbjZ4npqpNOx3MmlM7fMT6fWxExAXG05PitZTVFODBvQ3Hb2TK9ZmnrBM/Q
Ey/FHDschyey/F9NUwdn4ejj1EGff+iPQRRQi+otdUBIGCeov5Og2LHmW9qrgFWDfocaBN92+Pa1
N12Mbq5SN4FPxFLrkFY5zmbsk0vTmg9ova7ar/NdTkNXbyQ3Z21WKnl2z9VD+vHsJOBM6G+4BXJT
Qyfm8VKVx+AKzRFwdqtacNw7LRmCGAXWmZRVg+GVQG4mIsyiulgDw3xORfUNeuj1v5rnl4vNZZHD
cQ1JR+FIDrIDMcy3s1VqEBFwkwR2vjaMfAZek5g9j1XHXdlpb/AFc2OEFE7M8P1Kqm3F+lrM8I3a
9W6L2w0C/HZdurS9f6jMcQCA9kaE3qtyOQoJOqVC5qPEqcv0PvEPcR9Bha5gm6xOb352YsssMKLR
St9BH5YapjjZr/vyqIJ2F+Ni/qCrjZZq1e2QaWmHisO/FD5+Z6/5Zapz6GDOFibLghe4Uwi2Sw9E
T2J1heW5eOsyufjO8JwftxoI2/+10rz1dbuRbRf7YVWX4svH9aSl5FEap+4WxtR8+NWt5dumsj/6
yjBOmPwRDh7zuaC4Ixn5k6Nu5L3LPnkmXr7/CDLDhUSLjNG9V2v+LgmzO4yQ3D8gZlXVD4co/kYN
9THpHP+Ja9yuyGeU54dOZH2JYjpKawfUzhWz1ynlzgbNz3OJ8jfFR0yv8nziEgNjLIEfhR+X6gjQ
OKGYQHWG7W5G0Osoy6ma/+PUltogmnx1XhCPNumOLENc5pJA3+M2zK2gBI1T8bo7MkbM3GN/Ocfw
cCXf3G8ajjmkYJyAxwrXSyj/rcnSPMOwxp8KFXvxOnOnD9oJB05w2UmFkzgAMq2DURewG1rdmXee
Cg4DK5P6E5TVGvcz0iKrrkO/i7+zgj4RaMymaliGEDjp45RSogVQCOVlXSkvcF9JAbjX8xshoa6R
LXblNpPi4dpLCuFq2VrYs0rlYV8+XfvpfslgpnFxJr7fq68rE+nUKBsOPHRxWwdK7vGGKfUFe7N8
OW/hJbuiJ4j4jTjJnBkcTXrgg+Piy3mXFLtpXUdQ3qRK+woei5hcuOworD27BSNswYwupAu3VuOK
3xTsMAotrowYBwiQCAxm9fjRIk9JzRz8BABnQ6GtKC+Bnvzj7SHjZClPHXG8FxSR0/sHmr6fnW0V
PiK+S8S22I32KqMFGvTHRKenue6QGGq/gwClfURMDvVGkdpBa8LhsCdTKrAvDx0rujwlLPtrM/iA
qNiI6mki7CAKiTgEdK9m9saDbuPdRYeZ6r+SHPX8SbCAQcMPJ2afEuTW8TyaEv2jqQtOcaTcAKZC
ufov6gvVV6QEaRCRZtR8iTd2FDq9NKPmlr8iw4SBMIBwnU2F9PZmDmaMZJD29/JdKTgO1qp/hlVp
0z2Jr1vCBkJTmcGApLEOC0d73KzcRPjbQA4s4FfIWuTURTYBZAhktbJntkGDk6VrQyXTWvbUATwV
K+vARdufC4Zh33MKarvXuLCqBkvV7g9je0Ui5HhOpzmLewMVAeEEOtTK4U0YurkIi+klkEzQcS/Y
ikW1ey0Fl0fr069P74qCP9gkq780s5rl2AiTI8NW68tCG6EqAfBL0ZsZ18aU/CWeZsXmJhj+yjAS
YhLguu4eVtHPr1tZHwoZmtdV/7TWaO7GPz81+OtQMCGOdjKisvNcMXQfIzBCDzzeH9t/ddLjhpqD
myndla/w4jLIowYCLHL7WT9zisdSy2NeCtAmfzQjYGY4BBQYjTGio6r82G1hQpRAmgntC/mTXgpQ
IoIGugLv7LoNGXGAa8TZyiZWGbte6rnIhhJyXYMkpKwe78BNb5V9bJIfhLlW8feMtareKTwvtOV/
boyeU+fOtTVB3oMGNtLNXCrG2QUhXg0zKaGWU6pTR71YraoGArkwye0qBVutFibVSJjQBFpD2j5e
M4vWcPL+71ucae8nf0oaBRGRLmDSu3ZxJrbSo/xSOK5W/NbcjNvuzkDyc+TCuFI/hCLlfESgQRym
8he54ezw1+ABfBRvGS/0XsMPBIFT3zenHBfAfTCUUSi+LJO/IWTpMyAY1X97Bajlayu4Ik++h10+
WhT/MupfGaKTJDHwYnrMnIUR8VWN9pO/VvO9rWaksv59ERQDMhp5JgP4jG0n8cSQBjTLqkSYpX9e
mCGaFkwL2KpCa3J0MM/ER5N7H3dIrrBigqgC5bEVmZJ+Lt00TZQHKRFToqigQT+FK6VvnYzrMwz5
FuIKdMq+g1XkhH6tZJ0v6aD9JUx/ybL0woutFpoX50tmfzhywmrnwSzi+/YFdIj3c9NWqzHz3aut
2elOmg+muulJsCc9nQh5XiV4ncZT2zJxtNcJrUjM32puauDzzZICKjJoR2aZoLuboLP31BI+uCff
G9Lp556LRkRhyzWYMivPwfG+mnwPVyi5reL5JIS1U5z0w6hN/ZmhJO2zsZ2wwKLuC63L2/iTHzW1
OilyQc9C4gbBdK9BZrp1+e0/NFwiNvm9EEQ7B4apr43c6yr4VKq6SfgBK4iPQkX5CW/LOCYAF3Yx
mzz6WPktRpVvbKKWMQraPkd7l124mN4VPv9kXDkHEwmx+xHYLNnwt8JJvZOmL28hthRaQVvBytaN
m3qYSbE1GO9aiki4orq+w/WD0QuBk55L/TWSxPU5e2OkV+8tMfU3RvPHHSjR2N9fAKoOUXOvcNIs
cHlzAFo1ukuXJMtfjb/Zdp+5zkHO+PUQEtsjnw9WRC1DotDk3PWYPgX1plFdM1RcqKAAE3Oa/E76
gLswclAu8JnBwNFHYgL0vRYy8sLW4Y0tFDUxR6vVrWauYuggcWmZez+LyG/HQAp7nFTWR1xj++2h
I3VYgRnxCIxv+/fkvS+UxxpvFvaiZNodQECm44IIwJFdUAKVVSRHaU80UQxfN0SkhXZAsV0djDJe
CIXOrvIo0rPi3BWCybAb0EqPH/CB89kw5YqpZDunHwMg+fb6iI1/9zrf/lZmvozv2Cf/ZpXztLSE
y8xVT3HnNN/+IZ5goNdVldUExwj8RVq9Zi7ADSbx3zcLJ+pq3ENtZHhd4iBr6+KxtbJeiJTQiolm
bH7aafZjMzS/rEywnR6hDNhSjnTHVfS0M/E2QyCTNwEWh7DuEkVtkFeKTBgAgtsRf7CGEAIo8s+l
ZUIJoRlzIcf/ScgIIAzaS/zlWTSUbTV50ytaeNA8W+EzYc/DCJSUbLt4vNXEJ+I7uAfrZFHlubaV
WI5wakRErpEQLq57FlgTuyrn13b0yIjjXjrzCjrZYdqFDrg7X45tLxGhmBehjeLYw9RkzebjeBxJ
8Vj/aY664sLfdn4nWkMZjzzarAyQveElTAzbbJVxpOUqymTpgikn+LgOS4Ayc3WbzWWK5EOeBkfL
Lv68wIIQS+LrAUy5oUncN40RTdDMB2Rczlcwo26PrDqAoX6D1b46JR0+y1bF2wkqfVdJr+2bW7pg
X7Ibe4+C+8JoP6fU7BLjuElDaurDwa6VCfPK/47TxvNoj0ta6em8v9fhhyEpA0gHetMrU+9tQYOz
GeihDYKmwVXKbB2UIm9cW4GSDF+QrhUYqU2A6tVBIN1SKXkD6iRdsk2CrqG+e3JyHGvk3suGhYZf
oRsT9t1Px/aBDx3LKRe5kWPR8F3YlWJrHRWdEbeszJt9OBv59VG++P/6y/K8K/UYENX37/zpUJn1
gRPSMF7CNwppJuwTLxfgfOS44N4x5kblAztYd1IXoj/Q4Do0/54bCUnyCafC4QsCsHD37cwZGu/y
yuuVMfyFAuvOz3+ZYYPx3KvbKs1xPLT/8MqF3PijGN3FSNxARBXCdzGY98s1wtexoWSmL4flEyed
Q7YcOFqB5zYS+gAN1MF5SAmdUn5teMXfqULGzIuP/5CzyBv9pDQKbsag3jPMBfvvY5coTsQU1rYj
YwA4MRrnA5g7tLhzJKJtErXL520BoDyXfvhSUJbi8ZWrRkySMsx900p0z0THEmlxgm/gr8HUFk18
0xYWJjMFMahoHRCjmTCUaxOKARQXd/A+ytYQ4zhRJ/DCEF3QxQsYiGQi3t+HfA+0RMg3py2LYnwR
y5Wl259zG6Q6X1TInNFgOmEmNqaq9M26TNKuFwAZLb8QuUI4ImbH6I0Aeh+wUVdYjx2yRDAMDJKH
IG3w8Ec8fdMISkdiSuUmqZtFsBZezgSfTGgd9NDMJNXtxXc92gyymR87WOoKecQNEdzaEkWdqCh0
a0NTzQeLJ27JB3KR9dwct+uNZf6PcF5zgg6kOfyCcKMBZz83h+JgJg8axQa8hVE5AzdRiUNgNcY1
YbvQ2RN8TJ7iis1MWtC0CHOVS+OhZ67oJ6wQxNXwaVx+q7NT07XLsn2jXM/vQeDy+ibzD9lyTfpD
ja0WZiFJGXB6Y1aoZMJcnS1+2WLyB/t8xMvvyP/upJzUvOa1haqjK9MC+QhWGjJz3asDrJXPHDZp
nxK4FrdPjxY9mqs15IaQs+Pt46GKSHk9Zks+PHnTiT8aVVu7EW7JC1A9wTRhSZ1ljbKniN4909hI
Sqx5SuG0IuqRGQoYSSPZ1TYPOVVKPzp4es+8V6uhaN3AZe5crLM+VByNvCOu2DP1FvFI0xsISTCy
ku+z4D6FJJfs5bgrKdDfywxSqWhXnduSMvyUOfFNnqSUT99D2dLIBmqR/uq6njntnSKD+7B9wyzW
tXhe2LxPO/CPdofnloYOoqalXQUJacTcL+adsbfTwGI20sk3nUiGAyYuD8bgeVAGSppR1coR9DBO
ATAfvzOvzfQnAi/iQQdQO/jgygFt5aiC8VhoWyPF0p2aRUyhjNiWlQQQIOZAqSot8shNTG5T5OPz
6TcFSSf35dssNLiIIllenllF87gPmWU8XeZE/PbaPZ8n0w7y/l55+Aoe6o1Iw99CV4soR5D12iFL
LS2SyOVhquzu/CVK9XFxlCv37N/5c1+qMUn5/eZChxd3mOgCCklSCA7PmamydeL3/+XKQwbJflOc
b6s9wRzrpSVjDPdCIA43+D+Lf1wBCbnhZtSrJ5YxRV/InN2yglKPnP7wNN9tcZyciacZamvFpif8
2YMBjNt6w0TDTKgEYfe7icesfPzx0VB3oUWcFyp0ftpXD6DDPPguvjmO+7X9NW2s8S+SLDihwMpE
nHhgkHMEHbWCOcTxj/hMv6SlVIE2mbQio9kBfEEq6sTHD5+vS5XY/08RbeZqWvrGzUISItQQDY4I
hCevFNtnUQvcdNiDwUCh8HGRPTsmZpoPSXn3jFr7iMPHelGZ4EraYbwd8Wh1h7geojqW4epQxrgt
UCWCXfQrsS6Vw8oTbIIqAvkteZ5KNrr+3DOBsO6Kh6IIb8DvQ4MZAdU8bYJfCFZUscbWMoT9BA0b
TZ/2dhXUjHq+3KNFB0OmY8KqPMUSfLAD9N2nrGfiiOi7Y8j73XWfkA8wAMoKyKcXAMu24sYnrGR9
1h4qRCn7RG/M6bFtIX5gzI2oysMC8xNbQBMHkQLMWLlofa7lQjGJeyhE8I55mYPdrZdJYY4j2YCr
KNe+jz0qBrozwNi8nI5JomOcffJv/ls2aTMf6/MbJwswOxRtF7M8cXPYY3LmyptA4AAoiI8nuWoX
CxelAaTKTQAHHgDPv0aIiwGGFw6CYlL0r9s8f8Z+8g8SJE1FQM271tzFHI5cGOqRHJklGMu55bl0
Y6TGmaWtlJG4KZBPQ2kTmlgGs6GYBKu1dmnYlK4dUNecJ7syonOlTrqoyp31fG7C8LvHfoguNAbf
Wglq6lFi9zI7lhtdlqeMAnyKNDBY64ZHBPpZGdd3jtR1453oNYd4wOcITgaR86FI4tCROPumK5Gh
0eyQg6VnYKUB3ZteAFCR4f7/0KXAXYnrTOnz/hPYzG78bD5w7KI8jk5eFxKesRp/qmGv8MtRHjTR
fqb7vUbHDye1twEaQHGnMh1HkNiMS7O+9fG7SKcL9YOtHt54sPpRHHjqlNjAdLM9e5ATq37Jg6ld
HwwykfW97VCr5rVx8jW7dekW1QJJmGV7wufChy+4kK6GatzMGZOMtJV7T6RStgOx6zj1zVbU2I0S
KQPQM2IDo3bULf/GjwJafOKJqU0cs4yEWQ5tWt9PsMrqU6Z8tGXTl+d/GdUCB+DdKeStbn18PzJm
vk5AtEgbQtmwo9TEOAFfluE7lmI4qB5n4d3iYxzrBhJVvVhgZo0mKFsqlNcmoIqZ7RDNnQBzOBAt
51HWvT8oc+752MoEGKJIawMhvO6JWFMmNSjsVPn3b8UIBzyLrFKSI9PCdxwHNgcLPROSzlyP0qIB
PtxafVjifBDXszjw4el0J9zFZfM18goQJXQGbdsT03a1X3s9I7n9k/REa7x/MYkldpuzy2Cd93Ax
hjElKplF46oKP9YCRmfh8x+pistoz2Uqb/i2/Z5BQA/bDeOA6BJqOb9/Uy05aYer5cEgLWLNasAe
e5oONobMPD7k69JT2P/vt1XLMOekqdCUO29nnnr8cC1JFTOUQKsRFJfkN2Hoq+iFrUhIlGbhNd4r
pfQUdoY4rOzrijZfmmPiQ/XxWw1AUd8A/XJw653wMl7067Qe9jjLiMVsKNKoy84IDGzxx7hLhBKp
bAscHxRHHh6WUhZE/fvi5vQcK9NM8Ysvy67xcM0jQSdnSn6SVlKuZN3J8JmdI4s+33K9SF/uz23s
cR18Nj/nBG49PdGunFZuWcAINBG5NmRu727UHl3fpPVsM7KGEXg5LIxWl8bupD0K8Vn82lcJZzUP
yXGnYvIDkLVk8BhC63X8smI4MKOGoZFLWrWS5qVbuDrGIYY0X/hYBVRRaX8axjSp0NTf972FgMX7
d2lUvOkMpsmbegt2fhqlWmDGmqOXpyRHwLy6gYFkkyNjYjVPIMFVfgW+ZpzPnMZMZ+8o2VK20b7V
XHt0azFOR+JTP+3M9aXpNwhYPudjthZlPHp2UKYBOPjHrsBUjosCRtCGTslhAPPLF4Nkn3MaHCId
fa6OWC026lbeKT8pCyT9ff1CVeX5Ns1ZLsFosaI2ZxQnXh62fS+eiFEir10j6bC8BXoYl4XOaQV1
fAJufDcrkh0mfcToaZTIouc2CwOjblDjuXKyIP4oHGxbjxuiK156r5jcf85gsU3QY9YJ1xufDeQt
DGpfh0G6N+FW0xjXsQ78xTdk2WGaSzn0MykY1nYA0jkQAALIplidwjVibQQNim/fwzCBhaQdjvc1
TFreKydlRS3DEyxFLm5zTcYWqYhMUIY3OROXl0+nI/0XUtHCFnZ/LPfPNqJ9WgNgqtlL5hgjwbOZ
APmBHQaSrhxb+Ni/5H98R+cTnxM6Hf8BN31XBTNoKaN4EXl/Xq/4IoSd+r2xCuk8n+9udZMcN8/T
kC0PJu8WOOlPzW6WhjKBxDGBJlRAm0y9Qapy/nXqEd1ABPzvAF8epof2Vo8q+r5BK4stZfjrXHVN
eaSyVln6a8FHd7VHbdUUOy2mnyFB9KCPXENhK/0zgXU63emNhDbgSxldbj3GF+zoZxXkwq8z0KxK
CFowI0UGhL9i30kfyWtZ3tdfAdPJjexUwdf2+pFzlZ3faAgJl7JXy/ml2QMztTHe8/ynIv+OCkc/
whPLsHaDhKQHIwJjlwMmZMOOMLLDjAmce4bIe5XTWeP2yubwmZmkaqIPkY9xAej0VimGpG/iXghh
iyLuCPHypxDVwszcaHg/Cm1h8aos2Gj10D+4PbPdnRIY9fdR7CgU+cZickf2zNx1i+/fQPJDt/mJ
UrkWRS5OoPDc+b2xbPR2vSa2u4hpvgUK17Jmk75OcmF5svwaaQAY1+or9K9Zq60Zbu1tkVMSnGCp
wl+060TSObEBCH8hPSW0C0rjSByol64FzfRPJTZDFzLZ+E06WG9pVImasvoytN9biH/b+uUmBaXV
i26WXeYx9KLFtM1aAqbllf3kWuY8xnuGoPR7xeUXNJkds9ZqLwX7aTPRDkw38H2NXQgqR0wx+qeO
krsVqQ8x0a32j7BiUMeAWHUrWWBtwkxifsMBM2HRCmuvps33Ulfxz7xw4yZOvYHAM925H7IXCdUY
9iU9n8eGeggDYBwCTx5hGdVkgqihvGDzQh6Nf3w0ff44gVIXGJX7G6vzo90AohgF269K620G1TTz
fdfIx5cHoqwCRWgMZLr2QJs5SyVvYo5ZveBEhEKLGfFumTJKQI9HRuD2RSQlAriYxpNAIRwvd448
C4L+WmS9tbDfRwOFhrlwguVIUHGHJY5s7bWh3ukEQRG2sQEjQ7bagqQg3i8wkx/6uSL6/zLik8y1
geSGFSBon2rR29HvqO/M0mzOyRTujYudrhpm6UIu+cXCK83GxsfQG1cvB08f7XztRjqUL5a5oR1O
2bj9Qekole+rBCDSATvmQbVuAux3EiotSrWbozm9Kw/ByG7dVWs9B+nIU44ws8YXhtsHeKY+ckfG
kenP9E/Fsv56mCeNilDpe1GyOMsbJiZ/RUcGr2A9wNbnWgeCmHD4YYYdCXioJ6jZ4rK1lm1hEntb
S01rbX5mqdapO+NszmrHNmdZbL6V1mTI96JiRTZQrpW1vyeY66JPICa5E7xP7/MxCGcM7n3Pmoob
k502wbxhAEnfJpQXHjwmAPCgXgInuUE7L05T7EGmzR6zyHfi6o2msdTUpetPK2wEepcn3T5pXx3H
ZffGpQpqFo5KeC7LtVXkXsa3Gfnf3iXUPPgOktgn/d8zZ/QTXFt7i7wqlesr1vNaNzeKNRGmnlf5
7WIS1/8NjP1wtSO2mCAiosm3jwYv0tscf9nhIzlEK9YTMEMMQX8USYS1mKEjLe/G0JxdvkFtD6nP
9qKmu50oU6d2GNMA0kgb2khKqRerzYvmh7xiPKAdigy77upAI3ui41Rybd6ZDJFf9hrFfddIAYHW
wbnouHU3LrOCJNvfVfCWiZCro9rSzRzhO0ZaEQaZ0yRpB4LL5NYgGnPRVOgNiE9FaLVK1HenHzQ+
RhX+8bfdCa0KcF8MMYcMEhOEDLbTRidyJ81iUyTXTEv7E43oxLHrzPL/9m5pkXTqe5XnHv9l7HZr
5TJLjvz9xGG349Fmc9tOXZMNgI8DayGOynVopKVcvJxzs5hls45j6c1etfw72ttB1UhtSqwcVLqc
/rqUvaAkQbe9XlPXns6cJnxCljf8QzgLUWig+xmeQcJTso3LZTz4eXLTAIAW4sMeCwQiozOVlnkU
YNug5CvqSCNXS/TWs71lf1ObmSukM+Aewyp2DdteJtxbWMp1c6zyW/XgZfFqOykS9knQtHNESCZa
fILSMej+ND2KseehLb1uHGPqiCM1Ms1G1cozqb+8f09562lhoYDrKW7hJb1Oo2hLhF9LzHp9vWwM
JUcTDaAAoWDWgHNLgabgnoKPLTKhsbElGXxukR1pOWzC0nQdOJ2X3RY1GTfjEJZ9dPXJJlbEAMln
bFiey7csTXJJJiCBpxWTfRfLbxC5XoOZw1u6pEl9SATk45u+UFWcpDBMQIVGpBUwLMC9bu78bSSY
3P+BB+VkuAr0wXE6Pso4z98hPrWASdwJXLnaswItIUeXT7fMkgzyuQFRQ2SG0saARxmMp4Kxhiju
Qq65IyoVwUeW6kIsOkeNfwntOVwAk5/7n2qkxORUXr6Pznz2oJw7u618DiczrOum+q2h3StFCE78
UgJ+62M6w9k9rf7uiRYB/m94MiJTEOtx5g8N8U22PoobxCcqvWUopqWEzHbLqQV4f4yozOAuD6SZ
HXuV88ee/nC/i3cQrJN/D77y6lePdKGbqTN+ruthAj0qIEOI+YwvtE/yv77H0FUsHH445EXIpql0
oOd3h1VRkYP9oR6qw4bYaG1HjS0KFIMWc4xeBxy8upRkgJZDhbdHoWK4VFhfw9sQbaF52oBBKlk5
nqTK1kLH2vkcY/+flir/1TXQHKnzVasBhulFMohuRlOeJrRhzH6jjWAzJ4LsaE4Y2M2A3S/U0wxU
B8jOXS9sfh+beqR4moWlzx4ak0sbNMpIMouaugL32wuM2j4GFmDoJ7B3Gt1C6VLXlCRPMgr1Jcn/
Xq4hDZPJZq6dMsFhaZo4M9suibh0ow0rRVXhbhqi4W5pBDr4LaYP3xs7szQkAXAKx8XEM2IxC608
U4aG6RRdw5hbdOHYaoWy+dHHF9Ldyx9LkUBdI05O/0MceAlH8EnZoXxH4ejIY+BWv4yFPxzKSsO4
BlVUx49VrNHjWc4COBYjD+qqmlfytBGvmkk1VaAvq7QczdKRplD5wkUEvfGCjWZV6lh8HXE7o1Pq
79pTy74TX0fxq/H67NsOXYIztrQrDlOTwlo1Fmmcl9pMaw46ifQSMIdCbWlY5oAx1aUS0yVsaX0w
lOzktqoIXQ8E105nScbBtd8PKQ+3Vpn2Rh9G41affqcD3hyH7scFh+Vivrwztc1rpDu7+9yYZ48f
JBh2oLBanLs7V45Yg+nYKWlP7C1o/i6JSFGruQ7LeE5ZrysLNeKPzjWe3VPl73Qj9OnXkMFumkGz
8BEQ7PPBO39aZXLSgOZ57RRd1Ed1fA15XK+F4gcFzH/n5nYjODprdBrGOF5XirZp03PARwFRbGCy
vhx2F/bPx5hnlJXj0UKPwzuqr1kAEWpnbkDG6Ey5gX4rK9dcpYQ8JdzQ24hG/1FtIZAFQzdc2cej
pS2JbulSIIjkfvbQsszX6L0ZH5IZJcMPlJgkRxN3hBYAQjV0ABMBSKcBdC9UvqOBeJokXea6Tj9t
TFa32ixV+pk86tE+V8U6Aqr7iGAqTlTszITj5xG2vCYfUwYKjT/3IvT5Z8c6aLZqRT45zDB44No9
EbeKVZ5/c/mDsxsmQjWni45z6dLIZlY/lK31GESKSxvWEQHvlo8sHxBFZr8NUnwlo69BeMnEp+Qv
Lo/bhG16z5vJqwNJHLK/Zqw0WPbvd2oTSWetIwhgZ4XGCOnXw6x8/oMxY1bdE5tdvaatcmkJqUPi
S9MpCFcZPj1Qp1m9i4byNqs9aOrC+ent+7i3yz38AwGhZIwWEQaLLpCRBlETR1dMZ+5oA1F89ce+
0n5jrsbVva2hOrc9cnVtGzd88hq+v6q0PxigYaYEbAaIwevx/1OpOPTMLNwGQrsddfz1L5bJyQoM
EwStYVYCcrMlrL0IvO0aesSorYu3IEQYYtZsaw3tqaC5jxxyfSC8K9cyXXDV0b7duViMSx8tFBKA
HigmwT5tiPM/g1aOQT24mXgHvZPMvn5TK0Jkf7Das8DTSpKgr8nvh5WpvnzDRt+5o+ffRbxRUFQq
KFtvb0+FIRrUJvRWJAXeBoNuWjOwJZB+wv3XtQjJ2K/rG/RyK1a6ownmYb0U1pc8zV7GuNaoBV95
nr/CQk9MfGLSwRK8/jZZLQpf7YBsMOGIJDfyF89L+HT8ie3OGPxJVgT0y+JmuvDMqZHvdOyFjdkU
MtRI+Rlh+9HYYD1RC4om7bjIOTmyiZmEghoXFq8hMPM1nAuLuBWyLYNdS2lq47dyGS6g0TLmtAB+
wM7ZNi5RkM8aYOsjL5JSCg2BAL66QbvGmcRfaOhCWIetklAEQbRX1gWYmDYsGvwA2P8NeN1wqjjR
4YkfnqLhOPc54oN/jRedxnpqnABJw0SbNEVMA0D+gaeaJzckjB8cVhA5BbSbCaWjvwnsrrQ3fZEy
ySs0s9PXaikXMyAtoBDpITxDjt11KoB9pqfYU8dM2mMV2drDwm3SSv/lFLnQX3s/8pSZcfKs3ENr
PIatGFD22v1H+4KKqGA+AY/GKoxgWT3ed/TwGa+xmrZ0thLSbT+TdaZ0W198UfnPFejdIEb42VOf
4pzQDrFPYwCVO1kpHlaxrKjRTF2tsEwNcg8UtlUZnsLNYPCPSc58pf9hoeymYlH++qL3S9DOUQQG
ClgEHb1yXRZcS2PmSDzJTc9sgprcfel376yqrwmBgBaIU3f5sAFcLutjJ9WvbTewJEYQpupQOfWF
oBQZn9EgbJcA3YW7ej6ldRoBA3/EEOa5m64uW4xB7hb7zBD1U8nfVPXwW9s6gxnOuYIs/pIkTAFq
CG+WUAUR9yUiiLlXW/aHoguPBZRcckpY9+tlj5uw19hXDBBeU4sqpa6nShtddr57jvAoDYttcY9b
zCwvhf34rTSPIC0O/E4OSqDXxQVDm3t3biBMZ4J9rJj4jIPVEnf491ch3qzWmRMokH9ZOX0j8rZE
DqNqc+qHsgcRbm7b3rtkRSOPTElzMGIi9chyXVavtllAuI9Yl2hnlfNhqZ+GPNeo695t+aDy6dms
RF8NfVVPtUIV5qgvReGwrUWkGaOm33pRIYPcNwqkh7tKE2ZMWcZ1rOKZdn9LrklL+63ywIzu4+5P
+wIZe37i0WqH35AzrD047mcnBjeeUvSVW8kZR+JPrmXPXemVj4wADwLdkqeRskVpBRTYk/puEeNp
S+xeOP+ME1Sod+icRpGdPf4FYjZAj5/IoKnce0R9P7Btn5ev+i1UWi1ABM7qs4gjivSbrMpat2Or
DtvHRCbaynKncgb7wwVRC2tEGEolbjJOp0WDVgNcO8zMqnMyROpv5dFScwvfL/sD3MnltRT0v60M
Adwwltrdx+RwgA1LRmrDj4GofFB8m8PtlA2VWz3geYcfgbl7qwci7W0jhHCK9gGeILDLm6t9T+lV
b0Cy0U9cOk11qGwm7GgUR8aYQVp3sFhxsoYxg0slqEg9GCTK7fFNoRqq3QeEEZz2PAT7ye93h4W0
v3ef246Lv3wC7I1gukf/cmTV4zN39E2Df8t5JVS+ficrB0UJvepHbUelZFNzxBIIDZ2c5U2p9kdu
WmJm2FhLQ1dM+Oh5Pech+9niMH5m7qFyMYb4l7RiTNMcaWI3n6BKxT5OLxZhwuPBkYHQ8NDB31vU
IENHkvx/ygjxYNtKP8P3czcIR1jtJuiGNtHAn1R6mG0GxWrPCCZexobn0P91hGVYjT3jTrSOVgTG
m87+pDPsTb7Yx6nm6IPKZT6hCIeuG+EJkaKjb1nTvmBbEFN6bG1rGgDZKg836vzQ8adlYLvokqhR
hA23vwRMUKPk6J6zDK3OP6IpoNb5aAFVJu/0eTsPMAaHHQbiJPMKEU15XvvpRyGDaJOOWYqt9ZPo
a8NiryoaNR0kswUTs7tYDbgV/6A+dIBQaUY9S6/OwV7jP2D09Vv1wbTBjfCCvVUTxhc7thXOG+jg
krgZLQSfbltyB/M1mCyqjmNmSexmDR2Aa0MEaMg15DGp8GZb+UJpKEjUrUPt4HPw/pm49Xz9DGA2
B9Ov2UKv5z4zmGYZlwGpEWsx3OHDNxhmCPxCZWIUVI3X3pSo5AF/Ij1l0mXwP5fu+T73SqHdZbg0
Tv6LJ8cBZq5laCjVIx05aNx947/H1JUTmzGRm8Y7oOdsgh4e9Y+/FvjYw2GaqXvP57zRWfQB0nvu
njpVKf1S85M/++Qd+pWPbImYaB3eXlvMeAU+2U4mDFGm1EGhecxnxjkilZabHZ1excNLHNKOFrMG
8UN0lY4QNvfMJ1QUaxo8VQRI/fYNJvENJswZnc+7r4BNF5mDcba43L2fxiSrwz/VVqFZ4NyvK8uK
7JtGWD7FcfQPgwGVx3+iJtTO+fsGEzDZNBzJgWPSNggJsoXh0PpLuF6XL/VMzG6Bi53DC7mj5IGq
OEF6RCPMPBY8r1QTR0yoGILZs4+BnJbi5WnDrOW6StzmzYMSScY8wiL1dQIY9lnz1N164Nb7Mx84
WjAuITfI+9WPCgkr0l/BBpLmSbjWAPR9sW9WFZ7VbWGOMkNMiam0SIyrjRSZfEamJqq4v+Mr1axp
jEx9/JQVhpK9USlxeHQITGQXQ0Rz0xfXVVkOR2M/pnsO/IJl2OR5RDF3ovou/PYQdNn6RudXTTPN
FUpeBDMq4ymSaWD3ifGgIhp8GND1azedClsThSX4O9hnixRid0Ri2WHqRnLhHUML5wlxeRoSafyM
WJ6le5rXsl2l8208YlaCEQDMj778u9qXAoMNhX2HJ7czOvQkTmu2F1W2DAtKdmfsj31OJgcRp1Fp
awMXgsTgmfcBmpKyalL1i9MUMMOMWqJncAC97U1q3fGWXaYPWmkXWqy7yii+N5VbfnLNTj2mQcpv
nJJ1Fu5HUEqoR3fPP2E+fvOagYIIugDKnnSwKaRU+Gz2NS1PefpI8UjDYhOUYyZ1FTvdLsrbqRdE
V77Del6WVCXt6NdhyAtvUfwcZfze1u5EdjjbMRQjBZBBAJp/dMQVt8V1R9YHieIBVaKC3IvG41O5
8AKnWwCiXHq4BI1PpXcwlMIEdnIjHyyBvRc64fiWAGr2u/2MAfW/DJ/yXPvwoG3aG2jh80tq2iGK
4VR9Q8FcqTsO/HTRGMt4VaQeotpo8OctBnNzBQcFFO0GXKGUgjrgzjSeYGlN8iFULNF3NYPkoqUs
sprP+sXN11qQNeqnpVxUxLxsPxUzhU2AW/q0+MdV1XUf0oFln25iNockMqemNRbEjIby2rQO47Mq
K1L+roBtgD8Ro1d05+g578LPgPhSQfF0WNJ3wZm0By+vL3Cn7CJ9TLciyG4GfK1F2mo8d9JQg3vf
JWhgk1aHow0Hs29r44armNzTSwN2x0cyp2YAtgc6omS4pZQuOGrVwFFxnbupq5YHicpf50WV65Cm
dJ3zJyP95RvLhgigHez1Iqx9N0chBAoOlQXIZX34SZoH6beqmvdu0MUbJrrFDqEpI5OuoR49xdRm
FuZBmUwi894Uv1RjZgvmp1Onkl6o25vWDPOApq36sZhdlxQlt9Yn9FBxcV8iSej92yL46pO1eRpv
AJKfcH3HtfiKOBWnF/WVv16DoC1vPcgbXvqBQthkwK3sx20xQGBchzX9BHkkEag8/s5UiWTPlGOA
jHvH/cghI2+i5nQ7MYvQPVyG8ncZw9g1QIUN2Pl/71ckTizgeokfp/xJ6EvvaYYoNghjggTlUKnZ
nRB00kt7uxyWjWRcR7mgp6XNXS2xyAiErz6ZuZ/KinxNmhVH9kPiXLCYBwCF0i4A7kReBJC+igpK
SNgNlQphQYnlXv4r/XgU5fy+zrZxuADDksUHO82lb4BZnal2tCr3VFH/lKpKj7Bk/VRQ+o/b3VX1
l0Rdc+cV6omdT0dqbO72rQNGqCLfdMy53X4E49LbvmaAL6lddDb/0QW2rDRSFDdvtGChYEus2/iR
4Csghi77JweGIzDDU33j+6Di5saFSJgFhIe5ySJTcZD6ORDUKY7BHbXG2FtKEiQBpdHbzteGpP3B
i8SE9mmle5lIWcGVEewE6xfV4WKm8KpSM7o8O45Gl/s474/O6oi9pTI0gTwlvv1j0jIjftdYOKMe
A8cW3Y9MKrRlzBd8vLPtjO0G8owAGtTN+W5AMbVqB6iumkyoy4GxseF/PgTNHdN8kmckfv2ZBG8s
d7WYt+43Wxg5YCOQ8bhXzwQMkm8fhU2QsOegkDfC+KLXxAAW+o4srb6VwHc8RPE2m4Utb5eNUfiL
fer0OhXzvzZpBL1ijNRyNSmS23Gps6NLuJaqmW0YNNENwFXJHWpzQRIvWCBKMJvFPX0WLehTQJrL
LOFasfx5HMgveeUwfHQZ718WeABfnMfH6vFXhV7Ijj/3aR4B6O36rsRDqexsfhl/sRmKgh3ZNvgS
2NUH4Sedvoty+RfLj3P/Clc46kuUz3YLTom4F+H9JmSoiKoebpq21Jgc/dZrrUerW2rjDyXVSNlR
R6scMLddL3UswFtlM5T1HYpjUyMKwaP5i20FFD3ghp9Af9htvhddK8PokIGiktFnB9FGElnE+NC6
/NT4u0IaeGJyOUuOEzq5DvEupQ74N244GXqQvFOF6vxYJO9Fp4k8DHNtXGOUP9K61tfMXm+QMjdM
rWcEEAdQ0U5xqhsDIgOmySBTaq83ie8P7bN6T3AHl5MoLkZgePw75tyThhGiaD2ydBQBPjb+nNgV
njIS7f+24FvcgDLvazzEtESJMAktVwcDNt8QMP0KNWqcNWqPkxkIh/P/VJnYb+ii+P7dUlcUFJqc
5iDFy21+5g+N7T4IPPP4blgod6TZmve4vStaRrsbK/CkPvWcroxEiRno71mR1NCYcNKu4idNfx1A
28HVv+nUtPRRQ5GugoIJy9qpy9ZNIe1beXU4XheGLykiG60rYOgU5Zc2dccGZilUUzjHiiWXpVHc
tqhzWpymMWitHKj3g7eKXXHauJXXoDPz5vk4UIv6ZoRWq/m837FvrWd3OXriUO5V4XFfm9oLs4WK
406qFsebXTgW/+RKGQNOtdNlb0mz5Ea5KxVZWNjg64DKP3Re9uYWcqnHLprpmK5R0LR5KHA1L235
c0yhnnczqeN0DuhYvSgQ2pREjVz0fyoleKuS2jD9HZS5/Lq+G8v/u4WlOxsYHXHVAJm1uO1UcvNs
9rAV5cn2gsrghXLOB4xuKvtXDaf8rJ3FEmRJd685iEiO6WGiA0m+Lfb1HdgbVoI2FTLrEmm4pSDn
+8aoymcJprGvfZIpRkimKOfS3vP2Cl0OK1/AiWZ/IzAmj9hivjL2+wsYBDbbjAfOdJJXuOQSbJkC
HA1MEKoFEnlKW1LtkbzfxI+EKP2WzEc7Jw5jdB5Gfn3qRlZvoGI27raNdDvsfFCRqfIJsAUYR9l4
6I7CWgmJkP4iNvxGG8+ui4/rPCZryNCgb64MowKNHs+JEyVXtWn93M9u1cBlWKLhFicLontKxpae
MC4/fLM6o8158h8mAgPN6HcXtXJ0EcfBabxEjO8CHnMCoNl8mxLXyNXM6aWve3oQADafOWLpIGn4
lcvRBCNBAS317uKbxqU2I5hERmWWHKTUl1llgXDjM4O+Tw/892EyyAnOsGZfj5ubclSEQzKW0vZi
3aL4hGy7jSAFoL2MhVLbD3iUD93OZVl/oz/pw3w11RSM9chnJyf2xVFd/KMApMbUKI0GyHjMcbn+
wjWBVEQunNgd96hFtzrocKYxhL6a2MK7+yQrjNwQAd3efbT1icoSpZKH/MCWLzrYDAj/UPNHvkBf
ISJLpn6akGSdAKQgeY9suCqAB1MJS8+YdslEhUYaj1w9ufzECZSjA/1rKHlSaUCDwXf0ceYLpdSr
oKcCw6PMldsKuZK05Lqlr0CcJTmv62bjEyqNcxJiWPvtXRyfDljyK8Bh28/k6jPvhAi5ZlHYAfs7
DnEizE1h+SdRKnQKhympJqx6AFTRPHIDRfdf9xuLCSz4ynsrvCXtwJV+Z6hBkf6OMsHc15VC4wLr
euCdKhKKH1ym7YFKgfcTnkUGoc48q6j/XJCsqvpUpdtHjmEiGn9stDp9C2GRhAo5oBE901kGyVJ/
eheND9uDpu1OsUDSzrXn2W0PTICXrZ7ggXgVyPMNSOerpYdu4nONLBBwq6KiOsn3M46B8uEry3Pc
L9lmO06VwS+4SWZPiLJCk2bSanvqipKZaJNUO35GwO2qxI0lz0d5Vk8d4KoEZ4pRssiVHuIlc8Wt
0QlSNqhqMpMCiHfU6rWXHfHQ69lhPIu7XchmPYBH1hDttaW/4FopuKOuuu2RiMJvE0oMdrEwsIPy
URy8J7UV81t7OcAXYx8/aaCuskGmxyEFIH1qd1SF7Nb/QWmEFQ+GkV2fPyqBh2ryA1QImviGZhPe
exWjAEbi6MyqK9mqryMrd3uw8Elxv5g0T5F+ajoUEy+LfptUT/C1N949ckwGyCLpMbOl5LYOIt2P
CGM4M2SJvmROcxHaLC9NGNd7OwMxhvotDbutLbEoTXJa96U31M69CwWDn0EdPIuem+J0fn/0gUeI
BUYIJxnhKEkA59kKljlzfLYGNX5cHD96kUZBciinjp8yY3YWIzoohZPGDHvwI6Y9GZ39lrjSxo3/
kx10qO1L+nqcynB0XAf9aMlroiMHkmllQeZWxhsdeJ/Vd9YimvMd3B3TMqPlYIg/XwStwV75vJM7
mgC0Gu06DV1wsEt3nMeg9cpf4bi/i5B276abnz2bbRmiFY5hqF/q6JOrrlqoMPU1n5K8Ii+VjcA8
AA04Uy6PfLOHKsBSYpp68cHXy2ixzEDL1JJVFrp+3reenIm22heeZw0tqvo94Y979An9Ub6FtKbw
tFohR6ow7mcwGE5XXQUD9VQhtwYRLZINBXzCRLLal9SCTD9kr4wau0YfPHoBkEkezulEcDzVs4Q/
6uDNcDs3Ho9BDXmcljmaLUCSI4f2M1vB+NeRS0x9YI1qzobuoBHVcEXtt/qwGRu0mMIXB6CQOOlt
Hy5sHzl6ko5F+kbZnhKa2zUoYcia1j6NJgdoCBVw0SUxf8y1b961dOUFjI6Sun3lHZqlhuHo3jCu
gfLzFLeIgmghacf3S1RMe/R608Pj85JnAElqu18RWeQiu8fds/fMiFXvcx2BKQmXT2As9NWZkd5J
iD2m6H/mBYQ5cH5NV0r/Q3qyqK12i7kVLWNf4Oa+E0vUaDzDaHiial1tqzb/AsiD7OtdcLZOEW4Z
N/JRlPey+jPM2VQgI60si5NbwLt7DLlhwt3Ii/bosnjXpLrY1jsU7h8vdtS/RI5AojSYwnW/9DoD
QY2ptsFi3VVM19WTPluA0ElU5n1bGHvRapEX+X+bTSuCUWBpcxtT+Hsy2cc9lAZgyNoJ30dxIZK1
Ah4sa2+wn6LnuLU2mC6UnkhtHekiucYZhpX3kE/ZhGheMtAxNtYotgygav36u1L6d4WaUHkDL4MU
4a+kbngvK2cF/1KwpvXjxmYBe5lWIxLo6aEqAKU/aVcxcaV+iduvoQsydJikII3BnRfb+gIByyhi
kx5gDK1ykINdWLfakH/40ffnq3g30qLgWbqAaUlowxXvx3PeRQ5f3frcmfIHvYfhz/6xfWSK49MW
UR6+Pde2sRgTrXB7tw0ke4kqZz51C4ZCa3O/3vUZP6e5eDFCTrgQNxs1MXByf3ibla92C9Q/muBi
kn37zS6VUeiaG99GAD+Dz+RHD855J5aO5xn4rFAgzhNBD8XgRGACxTi3gszHMFdM29pJQQ6hAW7S
YHY8GPgQmWyeyUg8ebpX3pBRAjNsr3KeGF33DsCZMiAAvoE6fHvJyDvS5bFE0vtpb5L8BohffI++
W9jB/zzCqBzYkqO3qUd534W4jcPxgCNO/gy5O0pRn0eRhTWmaIV0jagdsaACRbDPbgcosUbl2445
kjAAXjFfDRk1+NQIjCRTgjnH+XFeSlmphijRb4IA/Jv92eGv21I5HnmIKb/27krC65yA7jrix3kx
Eb+x18d8LV/OytJHWQW62MsDbQfPc8yxvaXZDZlZiuxmS3dRYnRuev22FEC989tg6RBm9EvyY6B6
dyk4PKIquO9onXJFaPuhQgKA6fZ/2hTydob76b1BMGk+vWJS0Z5mUTsD/MOv0kmhn42eyrBV1eZe
sfYDA5v86tYP3IQbBpPVOvaa3HOIAQROnFul5irm/pKUJLOrOfbvJIdC5TNDCD3Ay2dLck4A2fTM
p/K3bNj6AmzK2FrFyOAsbzmyHWec2b6UJtAnqxsc4bv/FwG4MwD4imToYbDyh8m8puQg3kL8nqu6
lu/V51DIhCwejD/t/pJ36/KKl7A+6UdRa9ZllwAAgV/+61CJaaT4mgtzmwcJsu0N9+tYtbVmHV+J
/ZoMEhtRZdoD6nOCuYc77uWU8uc1/ucbZdYwLesxqfH/Nk/Y7FXfyCUF5ykjQH1AzrTWpUArjkG/
qHJYMswbp0Ka9ZvCfP5g/2UedWPyI62Y1kYJ87NvfZP0DjRdGGxj1HcEkuacJgxNO28saSWeFxAG
osHn0Du1r3nd80U4LJ3LbFdMFkVWkJt4c2nePf6ZMJ9ibTM0+JDI1D5xrjrZ72LCCFIHkLVb7z9k
M3LnB8aZ4otl38rmqZdDgy8APIU7GhptyyCAeYZkfSPAy3KzfusVrRI7Mj6/SlQ2KDeNOWQHQ783
4pa2uuwM6nEExhti/2ugpTE89aA+wR0zIJmOutROmQ2v/8uVpmqKBecAYniQo7m9yeJrUp2OpnVt
vmpZCQ5rGgMnEB686JgJgShCiCPIormXyf2ur+5l54585LQ/9WGdHgSfi2ONhBjtMCi3fGd9PMxS
q+cVPWsxUc8FXaglFPGk8ZLcoLNUBOK9CusJEpVZwyHLNSGMfbcDT9zB3yBjyZ2wGfJP/PUqTHjz
wFcLV3Im/SyWi2nWYhuCmqa8uLc6xp9VyCT40FYL1n4lyrNdQhfDBUslL/7n7wYdGX/7l7EVD7QZ
EkY+35GNVZcGeHHuU/8Fs3jcmsuaLp2OC/OYr9Gt+clSgEJiGLarhet5f6FeW+WnIPQfzpvnxi4c
xClotlviGyKMMxPgyQv0LoaNDrKwD1yEL4BZ1WLaey9TK1HbVrU9kRvfQwq6i/zEs73UkCwN4QkE
F4B4cakLxXNCbIZNNo4/ibqXn4jP4y4nvgi8Vx53bqk6Eu8M5hKMWDkRWt2Ean+h1Dyh/dhA7EOf
41qk9DDH7i3c6uTNkKiF5VfF8iEOqZWsr5vUWKHVNTFZj9LwK5VxbZ+w0PRiwO4FZKXXtk/LYXcE
GOOZbhO+bKVMVtJxJh4edMGChFC6n8pQwlSF6vgK6K1+gujIydY5Sn9mwHeb0YUJq0Mo8usWkytk
tmYICojcdwbtqlLxdms6qfkop4DEarvEqMcDrpuw6tjYW8NYWSv4EjPutfrobw7Ehqj0EK/qDVn+
2LaFoWLyWsR6IXfauwsB+0dlB/bsToNLmatNNEbQsc867SCShbpquDiOHhw0fGO7zciY+KNN7gfG
Ad0bYy/j3o5RzIQmFOZ5wmKJAcLzLIPK7Jyju3n1qWkKS/SGVM5mbY46hDYEuDZdgkYwQtcnCu5M
kRmzT75PZ68oz3NvJpruddVbxrhNSjQpVOjTG91uMs+j46tIhcC0MenPGJiXEWfT/3BUZoBLDVHZ
yeNTcXSTLZxfqv0+VwLKgelb+jiFp4k/4NzB58zHt476rYOgICEGWCVYiqFm+ADHPx6PiJbZxKio
iif7CFq7TJAvU3oLZclRXDUAaIlR3QqRyvjT+EA8MMbHS8qukYKFLL878Uahlv+kVA+pCv/WrIiE
IPjPImp9dofL2xKuQreGdGztv4yaZuvKVmxJGTj0pwsxS6pKhb5ZJOd+ZeeDaK6eOyXpXqEGLsMs
MaB7/yhUdQMD7BsCmDAiD7HjleGyld+y5/7OfGl1YbQJxyEVtvU1frVtDeQBcUBRTfc5gF6iR6Mv
AfbrYKNSVHFYm6E6xH4Jv9uA2d20aDmZNIhmMlUaygrkZkkpFxvxibjNeTBnJHpTpeSEbQO/Csle
dlYe3bVGBv7dpo68rOmdpziU02BIEnF5lhjn0GPitd0/hQhypEZoUx+oE3ALrkVq72pDFE8KNFmx
z3x8Fa62nHqXnRNoXeHPUla/kKekjTAkAd8k/IO/ztpev5VNziLckdjLYaLh7esYjY64xL3BYm3v
6AdqYXueSl7p2WLBsVCMLJabriCs4bhYE8C+IchGoEAyk/bMO9mkoWWHZ1DbKXYfxhIFgJCLfmt4
US3IvgnjEdVOCRdL8d7bpxOiKkufomsO9YNE9ede/3ZHtz5ECekyOjKmtWZ36VFWI1Vz3Stpb1To
WkvgEHpoQQPo/I6cbfdpA1vSrkK7/lVTo0vzXLcHDz+4P/kqFyjF1s9JiMbWLHf0RH1AP/Dsjgt8
ADIWrOYL7rwNLtB40UXsf6omYD5d0qxeht355q68GnwuMe5nRObYPAuLwInPIiXIIcHvBWLp0+SD
G1X69/t5p+5bkQexaTozCGy16BWWfG8rWhVcV7iVS0Bmli5QF1IMSDWhRkTVvU5kDYqxHvNE/NEa
sTzwHfJHIPNgIlTmiCYP1NKX8utH76qmz0rj3zWAIoi/4bwXN1pqlKGeOTuwCSkypCYsTQDm/vfV
VxFYryV8yFiftMdRjCFAziVaAT7g472TeAY5/WqmbwOfXA2RY7+eEsLQHPb758hBIIRB0T7k5ze5
cPkA82r3i4e5T3y9rh5XFDNyCH8n1oks9GuGGwEoBRN9m3309iIR/LvYJ2J+K+JikxTKmVCGaIIu
BJGhvgaQTTrTVSKsFqO4JwfR1De0nFbdsCwx2jzimc1SyyYRJyq5rN6VJUTGeN/AiluEfGeYOynk
E3nE4HrO6R5QHuYaCZZDGpNFb7Mdx8KlG8xDh6kBcfgqD9ophDdp71at8ie8ftm0P+E8Ih/ZA9IL
Goyf/h9yDHAlkWisF/WlElz0jWuhse7nSxQBKKnTSxFs3XutHV0/uhkqS79USa4iMJAE4qi/mLmJ
vUSmZ5UubSFzbyrUCvC8VLdJNU0nPQQUFhs3ewHnsB32Kjz4aef9YUPx1ySaQPezrA3+S7vGxq/w
6eN8pQBTbJqt524DTYsQcGCIGgyiIL6gNwn1vxOhIVpk0HgNKVa9mpSEnrDe9XloLJAZ8ELt293m
1fg0ayGOn2m73qGe0O2ZYsAD4ZLwbQvWGWYwxLpSuin7eOmYeCarGHtBmKkMLNNyjaLJ5ZghHoFp
YAbXX0PsZP88lJbWk3obdO5kUu2o7oIVR2N5Gc3iG5wTZsTepNooM6Axslpemrh586tde+fDmqD+
oBnOIrzfBmuVf9Wnx+nSV1Hm6ZD2SjBax3/OnVwBmUVoqZ6ne6DhqW/JOAU6PRWWmdrgGPoBb9ZT
lnVLyV1qokMMU8/EnFtfV+JCwtEtsmdrpAbZAnST7uEG6TA2yMuRFjuNZHAyUg4GcSI9jEgtgvhc
h68lrhtzS9gKVqVoQsw2RkjgR44VGrQpg1vknRU/3D1MQe0BcDhZdFrIz8bITnDlxAvdDB17bcaq
kHSmPCFYMcPZ7/M/VleeHjsFlqMlqU6y/Tf+WynJJI3Q12B3RwSHpfQYNtYOwgkqMO/CfkEwJ6rp
rvlupj/7+ZAL4qJKio2d4lud2Foa2f/q2AcGSkMj3NBMOPt4YjVH8xja45sVOJj9vn4AvJXXZqAo
ocsOkdBNutmWh8Q7EPTqNoObTP/nRYN9Ej61tLBwN45b/R+DLmvliTmZauxgNnSGR10Dj3NrOv14
Okt/LiPNNXKjsn5Ob/JWh6Qy4y/KmNko8FwqelYIfXSQfN6sN2qPC2XFE9TzXkHyZXkL4Jk8ZLf/
Q7/J6I2tC+XzVmh96yZAxWfR8qDtlSTXILPDn7ao/A7IFVGjFZNSZa+GuCYfUaOGoPNuTcNSJBxt
N96bpoqR0pC2P4Acmn+PXEH2rxi42PvvTX/Z5CyYUccMHhokUtQgPSzjfiDShmKJSuM0QSdewDQC
jJPv0QL7YpN8fHRhsRMjd7weRQY0/GIBEKXVKAnEvGke80tXEUGStMdPKxmv7+t/CL5QP82XMpch
60SKdNkqIfCLteyKyWZ1UyFSC+DFLz1rQOG4/zVe4cr+EaMbPNKAppw4ql/Oi60PK6u9GB1jc9ez
A7clox/Nbnu0oliovuTHXlAj5WWsL/4rQQeTFlwvuyCDlpruH41LY8EJiKlCj9OSaUBKgks//phB
0Sf39ZCg1Ox+/qLMpCfyqydbvv/CfidLXSP4W4rgRb8rrkO5l7RdTEBwIYP9k69isZzqLC7AiwXZ
8iiqBEeariF0o4lmxLzRwRf9WV3dcunNZG42hd6yIcFOR/jOFs1/DeqSURI8Edn9f+QXv9aJNab5
kn8FHRjtVruPJ3St7UcAsobjoAQWD3mD5WzmbBcrOFyiayo0KKcVcqrgxlqT579pNU6MSONIHN6g
+mrixo7UBpV3bhoGMMnj6/n9R9cjT9yH8GJTEiDeMQ1wLWJKNNzUeXroT4MBj+3RMKB0kA91Jzix
fgLTmCCyTmf1DAeaOfLB//8Jc2VfnXJ3JJCsyS019o3KZ9PbnuelpKxWKmjNrhOywxDJ1I2+IGHB
RZ/KhKZ/pwkCro7OmhKOXfneT4iuVzF7Eq7SpuNr+TktKJFmTLa4ofju0XoRqEoEgGVWpqyxJuUw
UYBE5UrtEULXQHwygzGc17cmWLlH09+gdTqxEJ9z7tEmZ4jG1AWAwxwTUlnaGbr0AZmCSk1O1X8h
v9xqoImQs1C4YCCB/LYdqqvMlpwKIgf43e++lMpzUvOIcnwRRw0aWiJtoJbtK+TU7wGQKh/bpUbm
MEzUZQRw3w41FLLOkgvrFvLH8K0m7YPU9Zeuicy4ogY87rAAdgWH6d7zELVlu5cb6PrlHGzwVwHs
YzMd/93/N2P7kd5NEQfmZJqntndKsGxHIaMhIXPkgbnKCqLLGcVJ+Gx9y0e9MSrmpbDR9Qg+hlra
gjEVwjLlKGBCb01NVAFfhnk3DwhIw6IvAuzjuK7b0Lc3iN0EQyaElqNjZ97Ul3Q2X3OQCEtHqQbt
5vddZVmmwvYVLrUdLbXOq66AI9qNidu4Nn99oY5MLIwxF58QK/w1G2uzmsun7dEhiI+Hh4RqbLda
O3gzv4SJ2UmHAcDb8Gkgsum5O21X8IfKfl/jAUK1RGRq9Af/Mn6tNliWRP9+B5jneW8aJUSdUpf7
vHt8/9w3cA8H7fgrVzva4xI3DWwE+qg//nk37oiggcn+ggnHb9ewPejNIdF9yrSWw+P7S//PPXbD
IGd0WD0MKWxuXN9P/scDaYxJqFoTpulZR+oZxMHEAunn6EUF2lBV5v4ADsyNAPMkABtZfxSSRcHz
WSv/mz5SPzVtFxfsxaDIWebkLsgXGVRQtgnHTmdiJbH1SijjKF9vcW2obThtwgHAmKM75OaxEyFu
H6U9noC3fojozaushzutP6hRhbsmIAJ2qRucxPoyq+8+P9nxgZM3RBZGjqCPqcMxDOdwjv2+IObE
yYbrEktWyrmJTZbvW/nlWISUsmw784WFlcOjCG3fl0AJyUvSz3WHX2AmavbQ2AYwhb59XHT62SFs
EwJGuxxR0qRzqtjGLRw9WiwbBXa4/JJ5QKlNGgRFyvZCncZae/hpU3u7tCLCbqTIF07qypotVh0z
c9yiTzjrp40JReCtfp/3CiroW911WORoJekg/NPD/DWq5yDG6Ko5wUxAGhIGmZ2AFOx0CBikILP3
4imuxtL2DPwALWoK4lbVIxOmWRHtXHJy9WgrBZaLLh7pV5dO6iqttD9aTFLwWSBufHhkD02I6I5b
Nj2yXAbgW5I79kNf49ATFhYVyA+6KEsYjI/T93eZz2aSEeyLK3kNbCS47OdcrNn9KWXaliw8pv8I
aemIbqhuMxBkAP32BlUfpSvY1W5ih5I+f2Ue8+Zn+KXDNqADpxrrvc6JX+xOdL5XMo4P6mb3INa1
pFjszyE3ThudKec6U5O4+o+Fmwfs6ab3GkQA9ynh0k6SBRXtbmyw+1STiopbvEuAe+JvdN4HSf1O
FEot1yPL++NJb8XzpeLPARaQe1waTVJQ+tbLNdVLa9kdNJXVQo3kuDtAz4hbQzxqdS0uuQu4lOYo
VspLYP+l7YF/oQbMh9QD+TQy5gE4Pt17fGD1wRkjUMBmTneOJqLB4kp9yD0rqAyvifU0+g8fWxV2
75Vnvo3F8MfQ1XQuCnsPxt7S7nBQyjpCLq0VYLpugHAQ8NJWUAwOAD7djXo1lffvUYUGU/Ap5+qK
vIa/3DN10YnYjUACXg1W5d/YX8hcgBDa/ITpdxsZwbfjsT+ayxzEUcrJhPZ+QVhzwkByVWdb34+Z
eL7T+d9DU/Hl278l/qw2qTk/MdM+amZFg2JLYINXOMM8TFPWqoOxGl4XXMRYOlKbj/J6Cdp4Xl5P
M3dLgGtclMsiuthG88B4AkGVPfBiznY4Rz4/3VMrBZtwEVQfHRh8utcDe5n72sUj2rDsQZ1jjPRh
C2LbwbAAU31QvzHwEYr/Ud6wC4aqQw30dhL2/m5H9Jo+MnWacyLrM5eDBYSYb2PT/yCFq8vXodqH
qE6MJwYOzBvH4Qm29LIgJGy326rXeM6ArEXH6e4R5djMyhzm4d7Igs7bIU4cafHnwHsI37SMJW7f
A2L7kQBJmbub/TAH/JmJ64pSuF5z1x07aFw7F00Z9TNBR6jngyq42ffrGKdv3lgoWd6vNHxZZ7sf
UK+pl1dkhuk5IjbF2ru7+Z7zpQ3mf3440Jub3K3WorMCeowqhjT2i5XSm4Oc0lgwTtP5kxr7wV91
O1QacVR7MuQNaGnJ/CLqyD8VW9zQY8CPN9BZTrxqxaS8WdxAH+ivsR8pH1cHhIWNgiKjsArgEoXI
imqEAHsZDSfNasd4J4nAxKfVHQZMksfGlp/+Yzu81/+8zpnX8JpXhQ/UzzEIFn37H19AjFpQ6+4D
8ROBxcc/oRqi3vztrEOo+SHhH5UGbTX7cjmhWWWT+RkMJJFsN6wfwhwzhegJ7HwQ9mYaa3mkk7nT
BJ61i5CAqWtkpOTS4ug5fCKIJc1xo13Z9VQ6OoT9ShsH+Uszm7u9Vd8+RfbZTHQNbKdbQ3Poldoo
vtVQNaU1lykf8Mb6nGaq3n3mzbOVH3eEdT2Lx4tMtTbSeg7A75Pw8qf5U5d9og0cU+xnoCT5yfUm
wkDeXWyLnMTS9YqYEsvKC3WQN1UJZlhYhJsi47m5GBeTqSFjWlsZZ7OssbwN43JjAa7IpWJNXG4T
Ktg/bNtaL6EB7+iZISrthRIxGRwtPzKTfpRK2ctVggedlBtl8SxftMtSBsn3AKcWKJ3ViQ/GWb7y
EovdXv+EvXqFrBrtPVHElGEjJtawU+cdtzfM187Z0Hc61lHSgiMqVQ/kxVl6oZczUD1MBjrUA8b5
j4JckAjmBHylN0muzVcINimJ4rJ0Fbxc7RiydkVB95QhyiaHLxp3YudV4PdOKMT+KWCJHu92PKMM
pLwvemYRrHmMrGmj8mr4FG+qPqoAGd2vNKNVxwXXidnUbbZp4wEYLRcRbD7U6VylXZ7yObSpYCtB
Rvooh3MIZCGIf0YPUmk3HdHSxksAvgMrXEucpzUo/VgB9djRmlGTsjX9j4wyA9MCKdqJRSfx8QbF
TV2mD+5rcZtw9Y91Kha5TnA+JXFY97E9/DZJuiSdy+UdTKIM9d173DDZuoJw/hA9PZQ7nTz+E5h6
He7y4OALt1AMja5qSwPiIOWQ5ecNRW2cFSvyD7x1cbaEf54cXvIYwJFOmcsu7LYG+U3eArHyChn4
jREuLbjHdpiv9v/bOA2IVVVwYbu7hnMyFoxb3wBpdUvyinWyPm+qGtYKYVHIOAZ5nboLt5AJBKWe
xwvWm4UngK+iSxk18AWFpG7tFrmJRXX/sw1ZXxSfT2Mg0NkIpABvO50SkadYU6U3Rdd9BRPPRTMQ
5Fjx77F4XpCDJTxelSNo7mcCSW0lezNcE/G3oo92vljkoQd4CWwEsvWEEV22puf7bqfCfqzLCxld
AeeX7stcJOAHBE68hx7jB0ZbYyrVTOS2/ziHeYCJVAItBUR9dfKrgjIdI5l9IKqFO4PeLbunUsQc
qEvbr65Sc8GfjhYoncYBQ1uLld5xChkUhdGYiNXV4RqxrBFklNRRHugQmH+Sf9dqwMlHVLCwyZ2e
X6Kazo6ghF2kMd5Xdlw7vKdRNf+04TQiItIeK4dUF+0T6xwBDr8yZQeRazHGUxTp3mpP29/CP9XV
6riq4fP2nCCts4AQ6IitHcTFNMzDi0p/O3f7wdePpCijW0h33BypN9LR+ja+//Z7ruTQIGTX6/9a
lNbPRdAVnKd4rixCOeRMxY1BMsoJqK1Ns2vBIn3wvaFYH9qjpGpFj0yoYP01HEuy4bLeCGlhSl8Q
FFud+KdkQ2SK1JgMdYeBMF/CtA7QPcvCO6O8VUvOV0KPRUQfMy88mbAa3/7PotsjOPK8aOISvQ15
auhOQewsCTmdLFWNfSsd4cmYWF/iC/3e5butDbk5cyVuKnS/AHIjB7Uhf5bTUSWJmpyeiObnfQy/
8PB4RiKaMhyyFY3sAFkJGZhSANbmC51HaZrOfjM+jyVmlupdB88WEaWe+lnFpDMMM0hsf+Zx03jN
+BrDlh5sTwZr4gAslaOMrKGGA0x1OH4yItOL2ify2eL+3pQ0lZ7J3GOi27/1kthZIjOsMc7aiobS
vldYx8E379RFyc8pUapSFgCE9YKi4VqYZinod4nx9EG2ZvShLZgU0x3Z9284Q0n7Si3O6LeaXv3/
UduZ4sgVpJq9OQgPOF7VEy343NDRRd85tHtmcugYji8BaE+6Sf5ZdrKSJF3tQTw8ROs5FC0BqYdj
h/jOnoI8KEVJ08ukiGnKVd0tpV9PXsY1AR7FnMkcZmveWONliTWiRE9DtvpbjxRHSFiETGSzy5PH
xbSKbqj+g6pcpxNJi591nEjM9HOLYnWfE8CaQFaWHOk7V9TzUCRmE7FGKZGOtFGAr5YKlAWoL+J8
8onnTOU8W7XeUHbO81XPE62+kC9P3YF4CMQUosma170tOX6iK+sV9sNhM4NfAT7UJ5fwTS1xz7ry
CX/MiWcczXzpKHyDOTMtnHpbiCuAtd8eT2YS6S34Uv0iJrMJgXKYrKhmZB2V4hC/sCLExnUY9kig
x3leegEwih/bIkUt/HpQtD+U5OgAzShWQ6/dQdzPZM9CGw7XyKmujKZdPxxstxzaSuPumjhps3lI
wsxlx+MqE0J/u3OGEKUSAmC2dxGg0qUB2iGrTYpfWJHbSEgqz+2j+dQFiLSTSC9hXPorG139tcyW
X4xbRiuWuV0kwmhC3OHLBi2SYtYdfzlhnHccu3jAvYFaY0WhHKhI9QPBKHwXB7QT0BoUWNgVSRO1
4HbeUQZQ1Du4Yli6dRwQBHdQXC3DrR5vv2UpxIhtzLVsW4Lw5yktBDa0ERiCjGpdzXOhmXnQhRRa
IB2PdWwe+Wro0uq7q2IfSEnpCMXTRvBpiqiO0V9j640gDW/9swx+YIuIaBnKvvxwHJE3iJN7w18I
huDJ2ZH30LLhwo6E2FTzjxz7UqgJD7amkZdN02wcaHcvQP7oaV99XphAV9CGulZbfZMWwEU5zueL
dqD0c/Ek5/2DUqxrragqvogmBvqs9Hkna4oVtf6Oqfi/MbdUGnhS5j2z64hagVTucTECBNdhYWke
U8NAy7X5Lz9lRiYFjPexn66BHKbSHRksLkP5sPgZ0tR/P/VeqCYFKNIvb0jAOWRBvojNqWzM5V3k
ipCmP+f095BLEJFILlacc6pftrExlwYNNUvULVK2V0e33AYcRbOG0ZpCqqdKtpQMRfo8e7JHJvG1
MLTAW4yqtSopy9up2rqsJDNeS8aqf9o8t85yHey+H0oGVHNUuYVyCX/9i+5FsocnZILU6P8d9QiU
eNb0jM3rmuwk+xqhIHeqe3cB84YngwL4/s0uX8x68dtFIQIpiIcgIEledcVzc/6p9OWvspc+cZSW
4zPN5lkVjM6ztUYRS3Z6s34rkcbMROvjoxw5UzM76dbl/haERGiOdb/JtoUWgOBV39qgzDE4jG32
IPij4kbXg5tvLotP2rD2Hdf7H8VaZk3yd/l7m9xPRhq5aJJS7QOMgNVU5d/Zr6ccNBLqeuc+EXwf
PwUXQvuYiBQPc5oO9rszLW0GPnTpiXKFunsvcBPL9iZ8nJ/Qawk7gKDAlWGhPHpQpruje2qTKDUo
CkduJpL+GqRToGbgbEqLQCbsGgRjI26bt9gjYshcSsJSEnZ7GZju/egGRA/qvH7U8jtmqmtGeCFw
6Z7VgYdIZggRN0970mKQU8h+Cpi/UPeWHYJB5S6YpN39+KF18om8ayBw4/NCuYuV5mdnbjz6mXZ7
QaOWIPmZTdxqpslQM8bo2UmKBS9YYep0iY7V7e7NzC8OoerI8n+2ZO7RCnvpN6Xnbbgkvp1MVfq5
Qzm+sOXLTucDvV9/HlIBCIm8S5TOZBvzdn0HsKGDUVbTalfCS8HX5tL4k8kFQiWOoYzIivB+DBFl
ZvVZweeuU2kXUEZzCUlPCg3MlMuodc4OP9Idx/cbvKNy4zRIAXOgvbpyCjG8TARb2HR66IbmCpwT
+1t2kwXttadKYir9wMk8DGyucFxYQa8JnSsmUGUdFBuUh29csWeJ8/Qod37cibKsyV1fC1jOrTG6
oNBnvdPqr82cxsG38rfGLtx1aanLdO7PMP2sf355KPf4uBhiGsN6ZWijAsi/FQ38MtdiV60Bd0+Z
6WmcL/h5X9Zs9HF76x0gMzFoAqz48c2zVyjBu6UMfHJm6a6iNVb+kkECwt210ZIrCSH1wBgcq63I
27on0ngX3MszFxuNViDuxriYe8HgC4tuZ2RqmzKnLIKmAzga30gZv35ZN5dpscEaV0JkdBuxeywz
fwBty9Yzzwws7GrTkfJINknx5p1BkVgHfFrwyt8soL+EDzW5gS5OuC7Dq7BFcXhSZTG94roL8qUy
SXcUL9BjOWSlfEmJXqInhtvFPBVbRUVJMK8SY+soCq3AL7eB9Qi1rUtoGW1vE2WBlIfIhReLw9RS
a71dV8FzklAak3H0tYixzbtYSsBL510S4ZsqinnmeynR1Yae5DH4iGQL3jJdU7evhiBg6W5PdH0D
Xy+8oBSElln+vd1SSUEqElLpIngSO6hUNG0/qX9Hh6iS7be7VxxOVG6a/3z1Zmzs+XmBgD5V5aKU
ysVipGhy6u+YiqkhfZhJaaHBmhXfndfGDatu+MnUFkwBJZCPsqSsBUHitMUhV4zC7wpJoUdpajsg
eT77TETiWg8NHBWP66RcDvRBglA9BXGmmZH7wBU6E2Pt+UPosgZlOuCtsKdAZrK+FU/BMkXQleMC
zb6E7ILasur3z0JsmyExhWd/XSuEvoGNBkDX6CawD5M8+73tWXIOW/S7B3ZkFUoGELl0Yu5cbD5V
1w0mTmgrEAWmWih+U/WrjoVkCFTI/wu+8YhULRrGxy0bnF2At6g87VHjeLEFy01jF1AWHzzvZakI
6YQcN1cIIbxytA+VpP2QpkjMQ4ZSFU1RW2b657jD8NzMPsCqvfuzhhNw+K5hY1We1x8tKzmlNLc+
gfcJYbMqVusH/62Fp2ReaEOZ6uNv3XsoizznpT2vkrUnVsVMAfBMYuGE+gLf4DoWlhpplxnb9lV0
yE4T7CY/wuBGo2NUqx0G32B8E4h2Lp7AAR4lBODFByscF1TBSrpp1v0O6TzduengkBgSH5PQd7ol
l4ON+xBAswFN1uEZ4ulmWAfJLAK3W1fNCO2lqKBX2BmW5k0+iBmkhXuqUMBxeBMZsn9EtnhGpfBa
Xr3bEmKBl1nezMpK7cyGMaECN7FX8xfS/HFLSprMUCleQ/BCSTyg17TJkBiAD5hgRixMVwVCvLEd
p31T6WS/de0Jf+JKZ26P5+hAmQayCypvV+xEiNCrmFE7zYBZd2e/HS1d4KcVKezJhl/XOMrjJeL2
s6nPxee6+eVuvFsn0fcPPcIrcs2Zoo+VbWqeLBWgrVxDUZTNyTVr32eGTErNkaWQi35ZzGjNBcMk
G5hPnoPiUSAwa1Y7JkT58ZcU6GO51uThOHx0THlKjnTJpFM5PEOYT2LIO3Y84xpXo6tZu1b3cb2g
fcpeNbgTpC3naKzvTsurAbKN3kXj8lr03wZzk5xkZtZBhyB+b1zXtKSRGTlixjyo/D0+QK45B7Zm
UbVqKN9pXmq/RvtGOxb/oeO4HqdgTexpCciOvAIo3rhZq+QlBb6SxzWeFrKYUSt+faeVO7OS+/5X
c2fF7ArH9QGr74/EBJJzdqF4tXEXyY1Wx9/yqXMKJDOVwydGagNW+t4HPANiyHq9wpyS3O5FkQHW
Q5EtDEHSL+lANonCudVjOWlZfqqraepXN0oBHjVRi7jR4cukA/s4UquD9azM70UEhU+R6NjlDE+4
tyMm19vGD4UBIRHHkmGBiAZHbrftDU5g+G/oQWdvJbicD5fKVSGljP6T97t2dUH/BbzgDCKo9Kcg
2/M5PP4G0gRhz9OPP97061I7UaehKG++eqH0iVsXGtVaGtkcUY6CLjjRbV6K9jjZckkZN5xUyLEX
HrIlanOwUN8rVV4b1lIp8591F4IjEde7uARSXjuEpU1FQDJK1cD7y0p5o57ucCsN1r9EMyRvT341
4v5IO4/Tfx/2XhuHrz77X3XLQiZ/hqlzyfvPEVsMtfZSoTNA6U5N9KFaKTDwLVlelJCJOezQrfqg
iv1inneXXC3R67sRRwPSQTdmykzyW+A7ExmWAEIcIJMtQDwKw/kN3dxyLGEHPpp/CSNP8GzyQl31
2vuZksZcJZtVBFEPiFezR3+PRQGOOiX1TRUek/2Ld3YU0QQg1Pnglaq1Fylu+y53U3rGr3i4ccQ7
J84flpB3YE7H5b26O052h9zAYoX3xQwfy8+Y5AL2qqEegqR8rLFti3mCwvHCHOrZkPbtk0h6qDrO
ivk95qi4P8G4BoGxSr1/cliXEDQJkUaZtDpN1tALfTKiQOChL8cuYWhwX+EfxH5O6ZSVhKLuZ+Ye
s2yzRPb5iYc1DY8q3T3HrKUMUAbozHdYkeHkqRYVYxK1k4ciUiC02mMS4E8cI4I2RD6NTVWlO0iL
OF37ZoMv0wd1oovnc0qD5ePCaYbrLE8edypkw6PO9h73LcdN/Z9edkloNaabaBet0TYQOUQefzw6
/WpN8XvcLHviOtYFhxDEpSs8mk43LuAFVoaTTOQaq2IB9KhqgG6q/MXc1E6b0sUs2b98Tlo0mEhR
ZjLNiz9ZG8DBJwwTlniVHzZvOlT89/17Xa7SLo0a2wAT3nqkTT9dzXzToKjyZdtGttwvGaSoXnd2
sXhxcCIaJq9FtGJ3A/nScqRGEk/yzMAT6qmUmyKLlTXbx27QHS/Xgij+8qOqf+Teq982mjls6wS9
gz4a8XvOcof0J0LJzjwI/YixV07TLDEYsQBpK/IsP+At1unWL0+ug1tZhV4nRck8ufwoc4DCyImf
idRJNJevqd/zObBpSfXtc0IvdFCl27r9Ija4jxL1BLXZXz7jzoFzClY2CGJQOUark+2Jf0DPjHNa
rMxpQrpBSFvxRBlok7j7q2ZgvgjMOmZ//XypblJiR8oR91K3kx+3zt+5JMh0McSwCoDrYjaQWnGX
lzy1Fq67UOMWW5v/M8zM7Ww6EDaJ3z+JpHF7Mv/uw07ds9HIiggnWK/rvFrvHttkrIF2zvTwTmwM
gvqvw/kRnXEMXNug1GyxbNR9IennISEQYn8h/ojRxEIUIaFAX3osbOIaN9BQrmuHqekgDcvktWJj
42hQjFWfWzbkEOYOroNh9F3tKoyPLrNr5RiStD6L/2uL+0SbgxcVr0k1zA337m1xe+IG1cbtK267
pTOmmlirdUWVT+bTUvZ9kCuqUXMNY5FnOYXVlKCwr25dqezONB9FfajqqvUfshWusuAg9cggen5y
uN0EyY9cqc5eaKwg2WqRuRZFrbvo0+O7MB+dpx9KyZRBYZIWucBttVtcXab45sdlc99k6tIBIGEV
Nb0xx5xY3CKA6fgp5UA1LwNW7QgCtOSkcNsVv9e7p+NEEKeq659SSFGANtnaxPMLYM3ujfjs4Mmf
I+uvbNfu2y9CbKYcGukFE8eifbW+Q7FLvDhlBTUcjQr8mjEI0oZkGICrsK3MgFm0wwG/jbJ2umnK
G5GxenRl0mtuADYVBmLjUJBJ9pBFmB+KFz4pVKjKBySnQLcQmI1fwzsKgFu7xazVZQ5QDDt93ewb
xwaa5FxjhfMI2PwlZLdI3+YMOV2V9BTsZRvJTCzaY+JXWLD9LadmLIzbmRQP/miS+fDCgItf+cBz
2SgSMZ4J3mYPJIIaVjj6h8WtWyrsMBfEi9LbpmQby15V9gB/YrFgR1tBv3r8F8WSF3nhxhshVlnK
mDi1YrL5LMig4wNPD6Av0n0vNNFVfpNmeah4mU/VYLwK2BrHKnDeH2sF49zRNkkDtYjRABYBmYM1
oJESvEOvpxLB4NUYLT+bTzp7u0crtw7FzQsQoD70iBivO4x7al6zrM75MQ4g/E3zcDJRnGiDwWH+
Wp54TngDoGuGc8hO/m9EDVuNsog7S2H/2YNsxPAU8U/384JlkvG1OOBQ5GjPeozOt/mW4UM/nmbr
/2ZV3HLAPR9sK0m651myI8xScjI1m/vNT/GJAT4Dz68dxBIvM05026cyCcRi4biu/CnoOuG1EWq1
YwHMw/vY7eGGwEhhqfvIpKFhU2qoYB52m+WeOxTeo7X31YnvNdK44w2xl0CFGmFotYSc68N6nGwg
6voqZtRFGffeEL86g7aRB2YhfYBZFGmbKv+FhUyU2pDqCUkfOOnF//G3IVvHR4dIw8lzAylBQ61t
JX66uPJpQQjaV61qhhd8g33Mr4fY9THxdCAWhSNYfrixVz6IWUSqWCSTMjnbQ1sLX6evb3fm3ZsD
89Jd2KOIkjSe9A06I2s7B7LfjNq3BkKaCDBSVHIFNkFoVB5a5t9H4xH5GbYneh7Z9gSaW4kCnZW/
Q1ZDukbgqfjkW91PcDcNARhm7C17eicCm6RVS92qKVUC/VJYn6p7RGwc5RVuckZCCnCLLrfizDo+
0zlIoNvpp7GfoywTMYQ4A+td6LP2MpwadJoV9/j56WR7WH2KBdrl1Tgb+ZVk2CPgH7ZlHqWSetwX
VIHxrmtpI2BCdr0l2chzy5g0F6Hw5iCZLZ40sEHtKumgeRPGq/j6kqrxdIeOmfuokbUBnfpl+cxy
mbI2zPmi1NnsCm6lSTZMZohFDg4ZtlJg3ARpWdo6cDfjCxawB4nzZVvG++2HuUs6OsPAId6TbJ8Q
3CxOWpt9Fs6CHaYjom1sBUyNkw/ha4cBW7+e3Fki22ROe0yeck8bqYx25t8sMt+4HjA2GDfm1PkW
hNpkDSj6xfqYKSQgpxM+mxNKkFNtyl6ANN80pX5iVUYQ2klfoZhWGDP5MtdPfoweJAf3bn39iDIq
4N31YcBt0q1+7KyQGEvHIEAmpx27XirYX2w1ctaHtkFI3LLGCpGpwk+jCB7UDlD+JDKI1ZSi9Bfu
L5Tgvh3SYez5/R2+Af62ie0DxFDp3RfxdLhLLb4GyQMsV9cxBDhDVJnxqX4yimTiVOYAYabYFLPi
AknBMibAalH95BBOC7rLcIuysezt1oeh14YAajhYce/OroPc/v96M+5sPD3kvsSLFF6+ipOuyPza
BVm/UCvagz2xW/WAL8z211H0TqXw1sCsnbrHkAgUHeYQbKC3BwsSwyDglgtKLLyrndwzuuH+IGza
ZQSJP8L0n8xFjfSxj5vMUeWBVoEoNZrrwNZTi7we3xFeQGH0n4fpmfUeURCW18gMvXcNqJfPEpNr
Gv365LOK1MfbgUCVdSlmUWQe9J39u46mbbWphgUo9ArY/j2Ma8hqin99iRk6C5rnBwYVJhb6lUpJ
8Esj3ZszkxbUkXbVCncgxng8GvjSHDX56KMdDsReZQ6YG10v04OW+GdT7rw+lUSaKTZ2br0Ka2dX
/B+vcenkKodWscf3so8p3VLOhpIQhM78aA41GiNsq40NJ+hJlAAMY/ebs4d3dIckhesqiXqPRWn3
TXe6vG3GAf1358XDGWeZgm4SOmkjPNzsj+SGu7iiGWLmts4tKtBOLr6vLVKMUTRC3CXvbFo7S2Cm
ugCT7YgyQfUKIwMAhzULr91jdXw6nAB3vand5PH86GtV6W7ulmLK+3fzKcooWplGW6eJI6tulAWy
nAtaGfPJirs/IHYFrm99/YZSb7X30Ka+oyYDGb3p1vD6TJT/nkUcBUEToq3HLMQAt8A/cRaQL0fP
yIuwgyMNuDRgwtxJDI2mUqFqhkcd+4dnkXhq6JLhIOD8WWw/Y4Kk9sp/yVm2VR1ZtiPC6ImWUUSr
qdRdhenywKduXfGm/dMHyV6B/2nx3V/Y44GAwECKH6AcZnBmZl17qbXdyKx2UhBQJPxWWQWIz4bI
NxK6+d3t7Xaxgkhsn7kWDH287Uan279aP4fsbTe1QB+JrxhXXKM6HDpF//gToIXi4sQPsXE0NMI6
65pUG0Yulo1yw++FgNXYRin2yruzAVfaroBfQySWIxVR+PZu8TT+mXQsY8/1IEmfg0t680VOU+Lb
IHCLCnNx9MiF51Gs2hnsOTG/6NEywA1l2kCsysrXbsHbgnWpIJWF+gljK4MG8maM4hchZ2bMNNTB
63Wd0I+I5TFYO7INQ7mRNAL/xvszhc3UjVAbRtm9xzv2vyhkpswTmoCsE+ZknuKfikmq7TgxnjoH
FdMkzxA2Tr3oBeWI8arDGUHYRa+9gBGsiRqGyvF/SHu/uhryAt2+thiRNx7iiSW/4cTswTsfhUYO
TQK561/UnAaMrjAwhDCntVmfDAAHE2KtVDNN7TPgZic/2lNdR6xFBBQ67l3ib3xf/fXEoq2gNyiX
6U4jueZgbuAKgFfDLFzxp/oe/3i7i0A+AdVExgLjTjsYF8ZDPpmhzh8KDQLwayh15DkImLvAquGW
AYlVEicZQEHuqEYc5YfBt7tgUaznZfHxMFfeitZhBXGsCV+tCUfvLDl/rmUSgOb62BBqjcND84vq
w44Q/a5GwvlgkDTEsY9uveFQFK4B7eilNZxvbBuKfd5UbtUAIcvk75JCEdu6D0SeumzUk0ppDqb4
O5qoJq4np64h3zuEXXSNM3Fx1D4QtzCy+gubjClBP/k3+lNvFOaUv/hC/7Wc/w8LlBaj88rLUZWc
qRYTTmDQ1MHbvR2bxmZg/y1ZUzJ95EiuatcShwdIoNFx61wzVadYx/XeqtentrRasV+dtlWaysMw
ZB8mOW4Juv7PGqKmiKEnNLA7tOF1+M7PmGdDk/Vc19Gb4rQr0V1upgcKFGZIQCJXpXji0nv7kufk
gB97sF8uK7Md2oQa40Nt1wn8yU5OTyy01n5PC2Cp2vTIJ5N6A1kHmE32ln87mV38HhEV9sCyBOvT
Scn+3zQVU93kXsrXfFiOeNeVweVtOI+2LC4jmXk3gZziHN1zFqKhe+XadvuNgoxBjm9Z2+Yu9xq/
rNVkral4VVtfVnvEos7EV6pXWlIcZR+Q3DFMylT7KvLNxGILpT7BPJG6yd0yiThtSH9JDO0DQ0Yr
9X1zaPflfulcF6xNR/9lrerCGvRnSnkjZ38WwpR5snflpV9brIPm6Q1N5YuV5aMhfBZmDHwrpv5G
7b4QSINuYwVjf6bcbuAWEFIXximNi/i3jUiG4AyZpNBKOuwfnlYwfCNEaZoJEACvYbXBFQrXi00a
zSYyAs6qguYfEGtEjAJdKg9feNZBLe5YlycX1ZGwCxHGXFGcpEwgCSqMAh3B2efOmiMyAIafBv7T
k6IrGdIwjfuEAUjwEARdHTiAC+cfdsy7TiAhfJmzC2Q40t9JCIxzhn86J7MbNi3PMyWJkySE/HJZ
ABYG7iFzMO1Co6AuEd8pTJ+mOLrhZlH3uyDOicuZB/vJuxrIZiu5mH1eHBtm+mRfJCtwek9t+4Wp
wfza+MCDag6Nu7X71IQNA0Ayxq6IpfHM54V0DhEswnJbs2ylHWcWiK9c92gBc477gslB8XhYLjjZ
3Z9opffV5Kuf4do+hQBRW2c5spuN87t4a7Ml5AZQIfJq/q4n74SvLT4Bhs65K5ucPkDR3zQCQXbq
sSl2frJYHltN8U4VyhMt4ZVffZOp5fgvyQpuOE+7Dttpu2djMgRdEkj3JRHp4avV8px2KFztESdy
uTdbUXB9Z8ClcMZKaO/Qq5yYaYn/xb39WVcuRs/B9nyLr5EYnZeI7uxb8TWduvNhg7WcSf2pYjPz
ODmHH6IotUYd5KqbUQ2yMRiVo0mNL/cOekaHJyPvz1JSVuWHFG3/xJojTb9rwv42pFXyRFZdQIfT
B4+WoUx+vLdNpP3a7m+E/wQyA9sMMslYgO/nQfOhf7C5Mi3rhI3XxnUZMUvwz++Bw/H72gp+nBgL
evUYC2zL9pQ2bB1n662Ctcd03/uOaq0BZ/byXVR60/jeGpviI/pt8374qV0pXZrfFKwdDzpvpsQU
LHoDzqnPzQMGxYKjLIZkB236M3bimKgUwoGFlQI4BFrpqg4roPRtOwOjB/S1LGbOU1GDSXdloYZg
rxSXlOOI6PHDPoTCSohuaXramyfNR5VC8ukmPnQSIZfobjsu5dRHach4Cw8nfiomL/CJBv3Wmt/T
28MvveOsn5KkyzmcNuq+vm4mo7oD1TCxBAQG5WNzPoCFcjrjZZEpomgQOOlTxWreT4UncNC3Gh02
xwYDV6pQZzDnjB4svuDXTuewnhqXj0ikcEMtENmsgVfbK5PaUV7GU0LrHTIdj/bJzo01XDICFWxq
pjJ1h+fjMYYK5uV2IbnZN3hsnuE+xDUSWzsm3sQuSnU44w2t3aXElQxr8CT1WhLfIjgap4tLoxHB
g+ctblq1O1qnOjfprEC7qK1bCCACDT+0eGJ4u7nQWiveklw0hLGu67/rckTN1ZdwbJD8qUsemL/3
J5dPsoZo0EI9W1IsevXqVHW+t2Ffks8+EdBokTZKAemC4l8+R4qjypykOCbtsWaQCUs4QmyVkLc1
fWKy3EFNAxMld60L+EXkY0i3yrdyr4KiWkvdkGCPR8ZSxcHx4pT9/inpOov1l2UB13yo+EURmusN
qbRBwUB1S12LHvEaWwKqLlaQTZyvdOkQ5ZEU697yWl2K3TRtdApRsfycQDCfO80iqClbGAk06VhZ
Xn4Z9oXeuVZodhbYvIZ8AAvgOKbXpFy9XbapXUhPQ7zPIxEhnDQhlLnJF9JAQnZFfImiT8B1AzTa
mXf2Lgkh7vmsoUSf3xTWjQO2Q+iWzrdHsOV1jzy813G/Mukg0bBoGXDw9EYGeA/E+o2Xyco/CDVT
QjYlsvLVE58OaDZkTEJJckDXWmEuK3FOqbFzRgk842v+uNzEdZx7QVr95KZpRH51M4fUWbKltqF3
bvX59yTNLz0LaNeZySI35wmwgpTDo/OeXC1q+6PP9cGm6H2iNftCntwn6JkfuMWkSqSnTqNB3yoW
xtHKrk5lW1v7u28MAhtQIBXRYM6OAjkCT04S/1xWvcVoQfQ9RzyB6BjLxFGCf/jWDPjG+UlMFki0
4m+ZmszsZ+JyqIGxXuTg6j69ySOtW5x4mzyZlUYJ38aicENNYoWHtKsphNL0QVgB09+UhBXNaQ7l
TUyIgdOdkikv0/Comrq21KSfynnFWyNjdftd5ynsNG6ikqjSrXE7ZNYfTfOLFN77T4SR/kIXLUaW
71ZKts3gywFxehl7WsPKYnHnAFElRCjS56DLdCbzhRwEynsWh7+DOrxF7PHtQjKaU3Y16ocIUoCu
94Op8AwCYdQ1YBPl8qkH7+L0er5DP1mr9gOXgTXbWNGoCAcowgKLJcahWBI36iM5xh+8MVFHkTum
EFKYgTpJ14ILgMKDugsMODhxhXjhG2rHneGjLGHk45u41RhF6qZDMsZ/COkE0CdKMFKH+FICxLIL
99w9N3//dH7ZfVHgHaZ65a7XMKR1ys7UFTKjFMUy9Xa9PIAj/7876G2FYk5lD2EA3YByQG6pGyoX
tBT3qXhgRsyRAIlrQyojZVzjRSIW5KLBbf0twNzEfLBuMkIisZSpD0ZSVT+BT06GvbfMDlxhPGzE
q9mhEsaAQnZiM7phVGJf7j/fXbdv6BSEB4SptODsVVOLnvOkOimJ6kFfMJ//E5bGRnpxyqxEipvX
E4gFQ8rTcmcUEWVIj6iV+DIj9y/QAKoIV6I7dlYayOa10k6JNE17PkFBXSqPzDbsxlQItmGMSDPy
U4C96xp9RhJlNeboIQ5Vff4AGo+WxM2gtZFS/gtcSUL6v0zkb9bMFwht+elyGNoI0k4QuXTI1R3/
n5ipU5HzfDPMGWKt3HPPz99538+7qeYSUSNXXHkFinWSRrqrZ8kFswLoF0QYw/p5QyD2/sPGoSb3
rY1TWX+IiazRjWhC73MThboCrXpV2IXvfk27krEkGMrhIvdrSncc89/2hgAIrvQyrur6/EpMJ6cf
+RUMPe2XL4Noit5QqpDzUBt/QpxWXcnw496IMKkJAPrfWHVNvXrP9uVLfmJwRF3jnGLS5mxQi5PP
hhP+LCSoc4k6qIJ081QVcQSYxsHwoZ10K1wMD5sKHqe+Nm9866OI5jF2lWuiDpOXjlTy8HEodZfH
U1lP3Aglm1LBm5/6+bSdWrgxYfDrBod4d5NrLR0xXyL7rsQAeD0P2zGiH9PEuomZ2DJHZ3guJ4WV
rvpt8gbv8d/2lUgeEOxKM8qYp5dWMNQYRjAyf4E+GXT3NXjfgRHnFGpOPFmOFrHwqWavgwS9yvL8
gkJH4KVHI7XV7AFCwD3wHkwTi6Bs+GHsq6vHlbK/LTSkxZIwsqKf9dfwknpmqGf949/nWJ6zxHB6
gyE55k7/2rjkbESExZgsaf4VWMff3wf2Ya0crhDMLRU75p2n/GXy9JXK0Dz863nrf/h5pGpFbqYY
ZAVBJ/BFiRQ2vQUmNyADbPrSc9nmx+OfJaisBQc7TZCGuyWHPQyr8p+QgRX0k4S5RBPt/KB6UclF
2poAz05jrIVNzivH/avhidv4LfSV3ScUdh6IeUViaIvgCmPLqwYjURZ6A8IsdPi9KhGTI51FDgTP
xF+Xng/Q7vZaUjIP2e8KEswqjNRN+88/0+2YdVhq0fpDRJG+zhjt/FEupvthL7Dt+TqVzkO0+CDY
RMVZOJ6AMS7N13Dql9BdBUWMMWtIJGn9C3+KbcgDPJndSZc8PMKOeP5Ji1mjnjtcfBlCAvHZyi3Q
aVjoSYCsMc8QapA1fIqwyGaimcPpHR98F7erOmwsdEf4QuQoU8Zlr47df4hfA2UBJydWuKSEZv4q
VJGIaWpSB3jCkoExjPBO+KujZgdY1bgQP7ET+EkpaWZlvUzMp4lkWbthg9C6mfKGEwGfKfl3y6gD
1ZKSKhmWWm+WUoB53HfJWjgBEhWxHJo3rT4lC2MbjPtw7+4yW74Z8Dlpw6Z1mpG0p/4pp9Zh8MD0
8hc7pQ28HeYvMo44FnXFrgX7j9nz8uqZFy+koUrn5gyvuUougF0a3CgF1QHmBfifoW/712NYrb4R
Ik/tT9QOhI2rALFP38wuSmjC7B/M5RGZveTNp+8Pv5MaBdS1jw/ylaeRI6NEunE3ldnh1ieEOrOb
YnDsfz0qF/wQT+1T2p5XVbmb+xPgrF0bif7dzMkkIhILtEzFMHZFOYtY17LvuTiyuKVawmYSwOLl
KH7sKEyETON1XqPoD5hh7gmy3v1C+0XpnSTSGL3OkDY8Q3xMnOuKMurpQXVZgTf4rDA6g3ym7tTp
DaxhYHU7be482azY1dIguLMmTr7ugZOMHzzdqTMH/Pz3ImiEuazpS8cLQYN8uyRsS5HPqm9wMgoN
Z8q7efHVWGILIiT/9a/1qNtaD9E7TPaDjUa+f9KWt8YXeYm5Gq3+kIYoD29v69kKewGT9ib0b7Fs
tGsjYscNBZDnZ0RrCBibkD3bVDySZcXZX8TMBFqqc4pHhxX8ESzoY4KSNTzF0oX4IU/7Xlc1Swpc
pndYK9BJnqU/KNM5+khrDNBY52EPdzdShCimtGkIys30O/QU2Apls0cIsp488aaLe/k/gCSRQaP5
Tom5hi8WuOrkUG4VBk0StL3rQeJejTa5f7i2eqDUkM5gaP1NLo44K73oBUegBykV63UgKtP1lW0q
6uYBpsKCioHaq7kmkoXjXGzPSuKuzC+r7lOH0O5MZhSOGGF2Cj3keGLSXfuFeI0Ya511SA8vt79y
8ybF/eiWQHIorKyhLxtsQw5q2RvnzHLwsl0cwPKVapGv2SEWMu/nZ4yKrl9iCv4wY5w19Hyh3Awq
qKah2EFlK4RwuhLv7rEptcpBVJFwapYQjLcrJgaBjHgVBTILzJRggKx9GIEkDPcicFW7nGNCXWEJ
2kS7qLg+4JAfFQqGOzxJWZbC4A0hIwaSnKpJpJjoKfpMd2p8uT9IwS71+wPPISV6swporQNk4e/g
aGsFeju4EK7HXvqWh92XRs2sGbEEI+aSXcjYxTwH4sGC4ZMW1W6DVNL2rDeDZDUTxxophu6ym6tb
vLEscFaEc8wI0AY3J7iQBpBycIcth9Vd+MXaw9gQwKG4WnYUPKOCEzhEVibJz5vfAIAuHa5IR8wp
93i6uhgKP/DKkSlwaEXPmFq4o/mxHz8T3i+n72R1BYG40aM00fJWazvmzM0YauUCbJoVlkyIwK3k
wE6Lh9ENqzfEhpS0GFQboJqsheOLeuKsxdenQTGSfK3UmrPGBlNPq1njdrUyLgMq0bei30J7KVwu
9IxjfTi7mzeZhd+D9BKFEM3yb/NsD47E8Mj4GOTd8JLjs3nHUH4qSFoIRXCubnhJcCC0BauqDZr3
DQjaDKfAbVhJ8T/K2lo6yYQqQRYrXyS8+TUkFeJ+dyW9spyMRfjjcdGAMoG8IG3LrrwsGaz7Yc6b
RdlZxtGhWOfeWut6/4Fn80GXDSGU92phK55roFo1xx0eGbVJe7BJMaiD4EYL+Rboi4eT3IaoYdI+
VHcOhlJSiXB6mkdIxNOAOdfVEY4ZXplQ9xs81p84jJ8MqfeLlwIq1pzv1JqIAYbi99uXawIQ8vII
dBegue3xJVsno/6AJFmaULJg9eC+yND1d9EW/SryfDHWB2pCkq5VwTX5Ggm4AFdlL9sqs7Pu/tqk
6cf690JzkzpjT5b3+lNutM+CDrluHaDlm+84lVaHGgWlOH5ZLj0/XYl650Xnt7RO2MzF3IM4G4lR
2SV4HsqpIXstti9vAfhBR4/nRd9kxhLsIn79JSPAbACSabdYc0kbcnxgqxOjiSIElc/3mnceBvrj
WC+uuHmcB1FmJVxsb9Z7txWN7gsBfqknCtuKMJSsb1UeTgU+x4Dq2Aohfcg7iA8eda76XMq91pYo
ESA04pDYhCSg3B0qJ8cOlrbXwnttgiHd6mz7uSGv57XyNAbV9pQM9Lc320XI8ftHbcCix/s0Kzy8
y+RETe+JskIKSQ7zCK+gJKD6F7Q8ICQOdGJcgzctNE29RHiL437hA1DezE6y7GZ+zYeZHWcqNpRU
azfaX64LQWLWh8m5ro8YLzGvivMfjbcTTaCRNV0b+CGCR2yJ0dYAdncjUoRT7hZ5l5otG8KZ1G2W
kzfzTZuaOIhaKEhp7WZDljuKCULAEc44cPx6Wh91uoXaoH7cwCl9CMAn3D51meS9VrG6cZ/OId/z
jnLwVcpmFWIX4dSK3RiJpG8qB2kLk2gnyYUcNCzK5kvJVl2IHJE/cYdph7AUfnQIzi3SzyV0XaW/
rmXCTT3lshq6FLnWPnYMNbuSMQcrAh2OQNhQZXssFcAnlfwJVLVUNDLVuvHNIl9vRX1BsM5kax0W
AfTsAaA/ZAf2GI6+LTF//rdEN1Pc1JmB/7bpe0hP4uHnVPaOzTpMWRm+q8LvfxHYpI5U5G3+bL5N
lzdXU0YgPLGSIn4orHL1cZm9aTIpozLGFiK5G0IpRFIih11XnZw5qkatSg00ySW8qSfJXnsYIGxi
hF3dRAZIRkMjxmh8aahGpurde7Fdi+KWhgBJBAjQz2JqGGz4Fb8W+OK8uHaYfVCV12YPIMYh0eZ6
8VbP1T8mF8icBA2qq3AYjaRFgkOITYSZ5W6LjTk3PuUetI7J8QKlFO0bifbEIGhDG7U91T1dOIZ4
HC0DY27/llt0Q6RFN11pzjW7QFc8UcUwEQnNmrk4PPKS1jnI8Vz3CtTwS7KbnZMB5pkvFua8i6BA
dE6IpiMuVDMqN7lg8E85ZBDDLDVjXO5AtM/aR+TM1fyi3sgA7yAwFC28tNEvGViKo6D+1Xq60jJk
BaMzNFofC/weE8f1DBVQ8p2CX7KtUyNfZ1vBTXACQwmKIQwqrjm0nrP7pse9wDiawoi1KZ8D0JE0
jWa5gfTvL0lvXEuKh37jQyDjwvVKTvH6cg24EDw/91SoREyKQPsLMAeAMK0XkFvSSlAFQ46sYXxy
ZOPoa+gWSyIVxfegWWUFB3+rMco8qCmaKSuQP3Xv+G7Uc3zQ4jb0Z2CpiTxNjxPNf52HwEvLHuTo
1hCmYc9OvU7TG44nqNPzVbKz4/plb4L5XiiQJB5WNWfR6BdLFxmaZr1HS926moPerWBmIspAbXyy
/bRqJGtu4qB0EqEEOJDMh63GrEQDQIcP4dsEWEmCFAK3YtjVaVFDvA1ybuMjd22UywHOqNmKvKnV
gZSXHyMnGvoROKO7esBwE7zpOl6jd5YuzIHyMFnNavxsGwx6231sw+GRvgbjBXEKMFv/sruvIIJM
YqHl6pGkolWVm0B3SxkWpDfUBhy6uXhvKkxfwWTa1qGReVJpevcFeN7jK6Tk9jjZ8btOmNOjtKUS
Bz5v1U8GwaYbVgZXYlgvrY4g0KElBLJ8NX+U5sinnwucPFJKdLzjO0LdhV3LIuvW+Ki0cV+bhoQY
VskK0simJnVqsE2Ipu0dUK7AZOJvA3cg2nMW7XpfkV7nr61P0Rhy5FFjFW6Xo/C3GWKAOi9aMaG8
Z71+wWcBhrxKXSfOFcvwvmOMRL+Z8s+t1Dn4I471CmuAPN8gwVIzws83aTrKJNbOCl+50vg1MSLF
pOh0OEJuR9itgkQ+pcb7EYNexlcgMzkrpLGiBnm6peUmUCV6EAmAsXmZF1wO+heZxBZw4ZU2WOs9
zl8wIgoIXd1sRarI4Oyng8DaO0lVcvZAHqMsP77D0CJ0uGYXTOJVdGrEYMXrY3c50GH44AOKYqwP
63gw6cdt5ZxQlVGUx8pAT0eEA048aQNdT7XeBDAwcEUsZwlRZblZSdZfIS1bgqzY/tbS25qIONWD
beICITH1hdOvLhtWNlZjimNyBWBAsYhdjB1UXuxH0hqo2Uv24YVpwp06dRw+zwxoyRvZGRRLhsyM
6YV32eFRatdYRNWUfl0EttrGHK5swiJ9sjoix3FKp6BdM+UGKxTcMoU7WTWBy7ejbwCaaVvOOzlI
jxVcvMRbafDxuMR3ymrKWr/E+h1qoOXnb2Lo37NuHMB2yM1hTMPdf47zU8DzJ+XaKl94wObildN3
7tSQcabxV3K1ZpNviTAGPEhKNoriwCa42AG9yPnL+VR52vOOh0COkzIvMqouUxCYOXq7TlAFn/jN
Hyp4/hx/2bNB+VPRhsWQQykxLv3t50GiJl5Foun+G5+sd63gwbDgXYSS+0RWjHjuiEpJ+rcYu+zN
hc/S8FwI4XQt4xcSBIQvcH8LMly/pgVlVnFUXYnA3KjneNh5L49yKDHjky6mQdq4DbVMLc+46KsD
Z5mEC5aD7Wz5RZIDEXoa2Tvh4PpCnBzWrYNVRbqvb41tITGYWbR/mvTtn7Esu5qIUQkfIORCnqJf
YbpN007f+yCbvKNNbrRQKwzE8biMNnDEGtGMOuFWVOLEPP3ovWD4G9NAI9q0dcBGQajvgJcWXUiJ
0ruogrv5358JIhf4zYTibM7PdM8oIDxiapdObx+DATnV07b5nojnPYst75Hz7vsDDH8goWi/YEMh
lzwAUe081Ag3xMkUexRGRpY1GjdambMdj465auCBLBAArbJPcNbIwLUhKRYYl/Agjk8ZkmQH6Bsq
Lu4lTSuF93EeLZng8JRDxP4AWNbyJh9f1YIHHqZvKZHH5jED1JjkT16lIBWQ4e+3VMWild3TYug+
GeQAc7DHX7+bsQDfO9aDjqrMxrFgGE2rN712hgs5dJrJ1RS1lEqF0wpw6gnqGTWkMA+vYKLtcvQ6
XonjIf7AoxVj56Z43sd8NhAlSDXUOY9Y5mD6u1Bqfb7vmGufB7i0LJcDQHv9dHCbaWy5gvl3F1uH
FclQZE7nrQwq31tmmPKgK5wrL5GMUj7bA6kqNtEclHtmoljw/Rh2oAlkYS4yUORKFBV8tVwMnMSH
lN/8nIQw/Alm/9jMriUltvQOHohdIhbZgu4h00M5DsTU3jxXU6Z3tv2dBUTSZRprnkfRNbtnUri3
niT5wp99WwxRgKCEyd/jFtFArzHCRP4H1qQ1IAAh/5yAUtTxsnid2gHul3lrdnSKfbZFtU2geACr
uLXKljB+YA8xxcLxSEg+Qgj74Etb3FO0I+wSZ82uxdHBfBx6HmbNu5QlzuPUUmsTktOCOpLsJfd/
NGi7DusCv1IPh2YHI5mHiyniZi+QqLpL3Nt+2J8EpCqCSo9hPTV1NEk6NgJB1ATJwTmSnspgrqrV
tEfhJpzfNbOwU8x2q2kAQOi7ZuA4pj4FQ5f22O6PeA5lxcfKwmgKoc8/vFKwCb5ql2UUtYBXbvhG
cyuytKDxr4/35Bq+afbuK/DNjmPH4GMR4xwdYYmxjuzmMCxMVnnpKPSrLmkiti12eovmIHCW3T0+
nzJLicIkQXae4BsjJ4I/18iqzoHe7X9mGVp4VCZczhl0tqBSx4yp0d0/STu1IFmTDuugejtMxL/8
10nYkthwOg7oCnqRa4nWTzZAjn45au96yNVZhgsQB0h2DnBWg0MK28Lt1+IvqDECgtj/q//IS6TJ
quQ6dbszmKQVUQ+fJuF5vryWrZVvH35smWy2vr5s/p6lLmOz4Mp7fIrYUSNhHeRrBCCJrkqWV1bg
88yLURo7TJXOUTFCjc1iiSrufuV1EBECL3dgvM8InjQI4sfowOU32lMru7qqwL3+3/V9HgD8lMrZ
gpy0lCRZ7aGUXJhRTDrf1ZWaAHqYrayhMLQnhHyEMMlL3QgNWZlCPZGiMGME1F/hkt4qJUFcxCJN
d3/N6ExcqDGa/HUSBb7Oe7TTm+Wdwsg17e7H0jZcKspRjrEGOaIK/FuKjPgNCL4Lk9rSAj1VePMN
lUc8awcL/zc7135DaACGi4vRB37plDsnytYhnMpb3Rjnai6Vl22skaDaYoT2RYEkF+TcGlIUZ3/S
boPIXXLPT1Ap/jfGdvwIJwW6jOQQm2ee4IVj3Ur15StaMbKNEZIZ87VZ36eox5KWBNZQsVaxI8wb
qfrg3lvJvEzzK/K+oVyGRCQ6yGS2+DZOucjUxiuss7SvOMcU+B4o8n+Chyo3Hw+OsRztkgbuD4zC
HJYg6BmgMr1BUab61LHgU+M5Yh9gkZymvbL68z2jEQo0G04ZolLKQETS6h53GXhdQ8+EQRPs8Wwy
c3GdPg4dOsaPEJnHcVDr75FKRQk7Ky51L28utTkHdWnDJgrh22eYC3xLULWgq9H3dV5Mzlybs0AW
ghvqTMbn9JHAd9x/M/i9pBkPfP1qf8Bh9hY6+csrZwnk2tg3f1B4X4Em+7/Eannr7yoriMu7Y+Jx
gziMNd4aSxtEjWYBPMwjIVWFz6/KNOt+P5JkmJhpQzHKkUQjRbbwjdMs2/KRfpSceU3hd6hjvTGJ
2XDFqhad0HW9p/Zu6C9c53hxbSfa3YLnEMPiJWIkNf7wYcZp9R6JPqWP+oJSC9Pa84N2dDgBKIe4
Dkcfs64q2JT8Y0He70SM03E/mnI1I1FF3KQe9U/Lv8fElqi1xEvHK+HnMq8VoNx/SpVMe5lJTt4j
18ht14wCEjgew06qC/A3X73KxPZGAs5qwPK7/rohumaVZSm7R6/bkY0RB312y/oBFrWNpq46jlSz
U7t7j3yTaQdXmfO0QlaJn4CS93K0HA1L+2hVZB+FxOwkpjTc14O87Za8lVW9wHp3IClEE8Jb1Dvd
c5+XduirdvMWfCdL2rfq2/Ishc1LwAVvCdmb/b5wc4OHkpIqB2luSoVj2Vb7XEtU8m1/2nsUShmF
5moST+BGrq1uZvOy7Z1PYIxrOzc5IQAAuhGG4jEilMrY50d0zGYYz6rnUsqq24UqQMnwrTurvs08
CSkrN3b7tDMz01MnDH7+X8imGtLY95BGPC2YhIzr42hgrCpHHOpty/Eu2P4ALqAG1jz60wXRQGqR
dAJxb38HwQMjVv37n2JzoBzgcPkqcU43qDRbYz+TvYRhqw7cSTGmRqQPNW75P/rdS+8jtTOIMD6X
JvBfZ778RCBqjFgbeV7OpaG7LffcBbxzrLd44oKwKBx7hf6U4DtZNKrwl3e2v4qtPKcDuGocqvCk
wZ12fkzhr8XVq6cVrhBlhBI+IpBIwFaxUVlsvM4WrtY7JzecTZYP1ONbinMFhH261Yn/UsE5Vnhr
d8lKM4lOyVGuAxJUHM3OZHNxdTXmZ5Wy+s43FzqiDZ8emfa2u1ig3r10BMIvYksjMwFW0eErOisI
RZ3YFSbkE6QFysm0TiqhQxiuDPmqjhf53OzMaNIQBd3MgjDovtaGOtKaAgtJsU+DHHuIPSEAnP+j
xa5DTahVC/lrtKTvLuxIfcEHCJMHJUolXRtieLghQcAdxGGmgLDMnEOSdj2L6xgUzZSYfGvXznqg
sFQjj5AsBWvor3WnpR7e+ko4d26Xky0jPmJuudwF/V0UAAtys2O+4OCRi3lW8kY8I+ILK/H81lBd
yo5NbJebQZRK+uc4YYpAJzV7mHbKYC9ADIIMX5MJsGHCUzIoZwOydgQXWtydOiSorfc6RNpwpd0G
DOpASo35zI6AAVOGFs8D+sWZ5NonaLJPgb52clOLkTMBK3D9Uid4T+2E3EP6I5/96EYxHbHhWt5w
EBkWHw5i5sJjtB550G/0Gs1JimmAz2EDGKzUChYCPKiC3Lq2nMrE9Zb5gDSjbY7oGH+V5pnrGJBj
eSspX/xUG5LgHCESRrRRpcIVcVKHmh43Ovdq4vu1c+qitjZh7u2eJ/47kxBw5xfHIPTbLaB44Hzk
nohkJXhmETRY2oS0sBF8OSrTdvXjZE6K+DhwiGhdhP4IY8m9o1ltPSgjXtDreBtMvpZnEABMae/P
wevLyXYXE1bomZ+vDtGUib+cCRUA2vpq17NBt7LEhj4GMrlKBkYm5qSyXkTkBiU1Ao1PKOrMKX7+
z7on0/uol7nqfZ8t8WBV1gOxEMM5NL/Hfbp7TgPjhyV/oi3AuCU/IzOnIvsg0vstvCnauPJv9BXQ
qs7w/aHdUmsQYWRRxvQpaOt78g+DssqVFh3Othz0v+R/aSurhZ9e7MMPafGcJYXk63eGAuSpYIu6
TcJOzO6myxBBTwyil0NAc0NyvX5Mrha1UlfYwT4IpbXe0Ud3XAuA6hCnbjw9Hkq9oVlLb+igwgUK
wCm/Qoa/JW/OUMywmbavrEGtgTlcI+ySekMSwaVjQtn1VwnbH5Mg+tR17Ddy9LopbXojGFswuMsc
njnLKSkNjdCVn3jPG05iG/lEsz4ESUHNHKfy4Z/ulybi950mlrlP+Dl3TnsfFkL9tmVxkSr1EHwV
OVyeuwVxh5K2X3Ggemy+srAJwiX1hbhHX5XjnHvKVgevJoMoEA26E0snoAAxDNy7IaDx30tQgUyD
7bh/8RIedUbSaRUHvzsRK2JMRRDIZbrt6VTjOMe/E3PdfJqvUiiS3750K4gVJfg7W1FpUPxHK60n
qUU4CnO7T+D5igQYlmWFll0d2Zr9/j5c2flg4CvXBp/mf6aKVUs9uCvlq1sO1srGSGk19Jfw5haB
HO7tb/+t5TQZwf7Li89Dk0tEs1fAqfCXZSkDlgXMinHmY4nYacQN8KrOOYoRKuMZG0HC7kieVRaj
Yqogwge5ZHHFhNlDZUwPPwE/q04RTDPigApb9+dIE4n58CZRoraCJJI+FzXEFrFm2v23IIclorQV
QADeWUQphuvXXdQv+LyoijTiGqLGxQ4CWo6l8ls1vVPu0tG50c6M+KrOWLgIPjLCZRjeBXDJIsvt
RicaCNvi2/h82pqpmWZwgv3pH5sOV8ZUx4VnJJaqwcfAVKIZjwSneqrQGsFfpm91D6STQG6uPZfx
KEgDCoSpcP4tmB+4FNWPA2+CfspHvwZs0mCe+w2ZQJ5MQXoeb2t45/qcqaNlWO7CAigAoVzzAlHM
wp8cb6QfUov2D6VT3ou+VehcfXfNcFLdA5Il7NU4LNJpVeCjhbuJu0pB2ux9TQqssS3xr/Jt4HVp
Mqo/ycLeyU5MOgD5JPPgIKVDePATru5JNsleBOHZJoANXzQmv0Agz2ATA1cgb7aMTM4OgP4o8lmS
N28+gAS9ke9NrCapqK4Oa81IcUjwfoBTiLDX+vvCqBOICXzUhAlfevyZvxvZ37JnbrV2UH6FjNpZ
FmhkLQjpsAcCgGdHH215HuKw0FooswSoi80YCMcV+gWTxvATmmICaLX8tdUf0/FKrg2B7h7o9OHl
wmSVdqE6+mTgO/SZkJEmwgkQzWS5YDRfoDAU26fw/cLYAWtQqpQ6X+6v4jwWZklJJk72+W6RD0FH
ImJGOhxDo9CKSdrqq6ADApTvPyOQwElrkLEGlEyXAMivchk47envnepAIYYwcTTdxVeXyvegCiJV
+J1gm21sFm4ZwxnADUkftfq63Q/AOwJ+Og2mYOJRQ38VwSwZz7AJHidQmD02DDgo21Bc4nFNjer8
6gh79l/snGUd8YQqMBNKEi/cEsftX+3UZa8o1IQUUO1LLQNhFQK5lEqQyyr/zLUEeqGo+EvPC6Hl
fARoLFGAT6KMw6G63KxAi6RT1bp3VGX6MYwLGUKJCxGGvIM1sF+A/3dk7GmAxvwAnHawcx2j1i8F
yZ0pRmeHOQf3KLYVAQdms1W3YgsOrVwxAIFZEiNjuoaGWZHLVMSIHjWue3BxPhUlUwIKoU13Is+v
pEnTZWMBWVID+K4R0/V5GEZHZJ89sT5etaZOOK22oU3FdlV2Prc8f7qMbV5d8O2lZY2qlTGbyo7p
j4APyRjdU7LZZe8IlJDD95xMLhd3YEcVWnArV/tMlvl7y/an1ybA7eUIoWutGmXNQUFvOh/Mo++5
xbU9C+0masfOa68Hmsu3Knypx3fGI0fgs/USb8h22WHnO0wkg1qLxuPMaAf3ShJ7SxB+me2VyOPl
RzbQg6Bmw/pUPQfjj1Mo3GNs9IwxkLEjwZm9B+E+yFU6gCIAGXL/oBbl/aZp++W9lnrqS6cMcOIN
do6eR4yE+hLgZzJEinyQ1IEFAgfb0XgG8Ij4rsK5iE1kzw1nZiheLyxFwr2Xy3uoSGrpK6BywEW5
S3OhmCge3HyTR4Ki5D7OFMw8fG9zQbripMkiQDxiQYLSWQtFkWgwpOLh2V28Re77KQbT6n0gDGZ4
yELn6/Q9Mn3J5pgQzO+QNOhIUQ4Ku/9kyJCKw5Sf4cqHstfoiWEGQH1OFWpdRb3jZSf+SuNIJ8Z1
gx9cG2QPV6SJVBe1bIghLxzky8tQsduqsO1dJf+qfdocRBFY+CZRAEtnmmVOP5RN/SqjTQleU13E
5RKsfIoR6ueOJT1DaAaZcErnA2djwivVmL2zM1d+dRVdftjlSr/9aDYyIOAGEe7vmFirWWc/PwmX
ioc07fDzg292VL+8rP4hLjv74h76SaFZV85bTbSg9civ5eVePBhZesTmjSZg6nysItRHj1Lg7sxY
FwkauTXd3VYPfclYYwCVgHI+D/0TFcn0jPmM93IPJEboscHz1rqj/QEGIkF+vLuUQc61IAEJ0TGf
kyaG4CZ3OO7+ZqYhEUfL7W0jU/rm5qIlYlmbHLXw+gxENFh7oXV78JR6EUlMUvR3kU3cYPxGyn2J
ZlTjZaH+BHT/gDRuDQ+x9bEDRrXDPu2E7Skwpf1k7OLszT8mfrgNCE2uOleu1Mx1k0cbrL67CMKX
LHUls1jJdb5kbLcJuiFvnehHOSDm3dnqjHqyy2gO0M6/fEtxYammqv3Kioi8Em0Jn3QJuK8e6Tr7
Wk0xcM8GTv+wj/nA4UlrT6g6ZAy+jvQSnQbE7c8f4bg5QLgQwkP9lFRvkkZsdDmVKMszl6GnyRqY
n0eC61BtgV5cY7AnonMxJ0DMmTElLK2ZgVckCANvYo8O30aaA6peXI2rhfS/LgNbELL9YwFLnAiE
R7ra9OptfLb+bTvNFcdCur4ppRIX4uHiUpgJgM+bIQgFCAArtOJfcBFRPTRkPymW68+z0QbyLrKK
S7tRHONHkOlRqQtS9f6ud+s3XiaMHjFJ6pBzH/uxDh51c5YCPK4FS/tq0IyrnnvrkPlz3KVYap2L
EeSafHP94m0EXmsd0YCVVr57noYhVk+99Pz5Z1LpIqlLhSJ3AkV+HAMF+ro3DwhZFWp88CLdeybV
0YizbfT9UgxGYmzjserihIW0gouYidPRMyVTGO29AYdfR6lpnNchJ8uiScNxWyCtg4MR9GIIODCM
y5w7qwli/z/htr64T2FBthIM/ZcBSfMM8DDYb+dlntp3QPBdH8PnkvsY+cNv0CO4RneWGMC+Nb7J
90mIiB+hO6vMczp1wyczrgyOExcYrgyl1yZYXCAXrpUmvrRQOtsYDZ1lRTyo+LSU3LzbxocLcsUG
1dRBPfJt96nJiu8UvmThXMUmTx5WV+ZkLud4sRGX7XEAYTW89cX/QBPXCFBcy7gGb22M3XWKl1y/
KqERU2YoNh5p6z26Dtnvr3MIZn9mHhKjb3KWlQepzwQAczAj56KKi1Sg+9mZGMsH5QBMLzXsKpFg
4/uUL9u2G+FfNrbHXZUsX8VjzMs2hlrmDtSdUkOEXZW3lYsFTKvmMfyiapq0SWbVWqALiLamWdUA
d9mnnkp+bP7dG62vo6xrlH1YRdZR9fvm6FskIGP/igVe0BApbvbYKQReHy5IV6h38k6KLl0Uy5qw
WjaPv+xLYeWkbuuJWE9T1RoMNkUuic54DCA2qIjUMPmcU2ATWXKDwXDnAwo823BLn//69E0NffZu
JOCIHJPtojNy4YzeuoQCUF9Tp9uVFRTjxQQZVUmzUwBwz07mPzdchndXov1uCdpGzHTXeT6Lc3KH
RBycVEAz1waj9N3pqZN/XWQKnViqBH1WEtpSua+WisUdiNp+f876SpRqiplKvrPYkq01mNGmtS9t
NB1+2JTEse8WlUm1dbSvLTJmKpOnDhFGObsRh4TUIp+87J8dio12oNwLztBZxR36igppuaMVhjA0
s3i6JFSPOQ3sx0tuLLlDK6rfEQZ63B9KV9+BmQ3cVXSCFDzufKFbUf9rN/d+lueBM2Ky/F9DhoTn
DdUsx6zYhoq0nGHV7209T9KeRWJpqne8w9zREQJZqQBb/GrCFD3h9A4CJxyTx4wNphIindpd3eb+
VCPyvDT9lTk9Qm/U9NfpEn/GzX6BAAZMqYMive+WHuJjMX9sVttj9MHyluS2qVU75RDv7NQeWnPj
bNquSsJF4T9fBEM58lvbjlAlLPSKifXmPcoaoyLDjla8qlASu9Ko+mYWtNHX1TMMPoS6FRB1UsQ8
LEp4xyz+K/7TLu+uelRa/swcNztWQUmVrzR/HLK66A3nmF9SMbwDkXQbYRZq7l49SYKxhDe52BqK
CMRdNMhfcrQWyEEYCKznJGSqnsq4/ZTTIPIDniDVn7Saz+/yHydiR4/nOnhR8UFwK5G5qX1/BHeg
wz7eeIWa/1wBafmmIllHqFKOn3UxafPJx1L7IsgA9Qp/iVKchJ6X8+KlPX+dmEihydyGlvGeJ6Rt
wLUqX4XOiowjF/6Mutx8kv8Nkwek0BlHA9XAH2pa7BQTDy7DvFC65p4hZOuOTHHR5cUsiC0sfBkB
yv+5aVawuvM8swmJ6X/CGvpEPgmYx0Rw4LuY5whBMXZ4uMN2qRhmoSD9oYBOkNu0LBXQhNYMZGja
fE4epd0F9KcfNBQazKK3bBcztdwtowh03oaAgegd1yUyfiNAEdUKWc+g4Bqfo0fByKxvCLSBsFBj
erRjHtK8uAphuIM+kDnMzFjEabcP5a678jLdT2sXH7LMq+WhMHu/4uYyQQeice2EN/9SsbVi6Oex
FR7IkPiB7mmkRggyc1rBolbK5DcteAls/7uJ4+iZe1pxQ50oZQ9Y0MgmAK4RNtZZdT1VrJEHM4q/
CzvS/+UEjF5o5DCIO4L5UYd0g1MsqkMwcIeFsiuF/54/ZqO6jYvsga4MnV/GTxNFtC9M67mDzlw7
wVoglep50njqWMDeny5aQBQlx6YBFaoYbzZTefMPe9bSklPJIhykOzsC9bpBp3vqQkd+yq4AnXbw
hkjbNCdsgx8coBb5QUvp00PACx5gwHXmbOlHJ/c32gvqOlW15Zh9V877HRXHLLUCmcMihzl3LO62
RERd+W9rNJc2MT9i7l+t6aoEK2AA5kpieULK7PoDwTi94aHqIH9USSEAEm7bEerVvp13UqtNwthW
oiECcleN2tybAyBnEmhXtGMx1UgEylU48ecKRAYwvy++1uIzT5yiwfZCQWaEMb15biaVY3ddBfW7
W/hPSJYapPKI+aUEiKTGP6jIZf4pLELZt39qFcHKje1QgtxWhXSYae1r+2JCJMWMd/Qf6jKzVJjA
sj3IY+sELgWyz4XG6aLeZ62BzLst+Om7VU/BMnftcbvhI6nSRoHkXca71fSufV26OjDjH2ykMcp+
iJEsIFMcF5OPDJAYeqlmLVqudVndnJ6tVCREPKgKtYMwXWajiBRu6yw51zQk2Qq/jzphTE/vHnZC
YY7sLhTOoQi24F1d+ri0cKDdgeE59C12Peuha5L5FIKWgMT79gMHC8Tf9doPyJbHwGhNNMBQKVPH
3YvPT56tBT2ocUgZa8sygvWGpEHj6RG8bdqq3UfPAwRi0WmXGj3NbHHC2doZlyKIk6V9lNUWd4XE
5/Blu1z704pwUL43BFg+6IvMx/oIL3f+Gf6lAdDSy2IGOFOso9GDP3KO+D9ARVmRM2Rp359wttt4
q20RVT3W32WbOyd5qmh32tBIQI0m/7wva3f4/OKLKeO8pUpgHglLqn0Gz3MGeOiF8iuUWWOQF/6g
d/6NIgbcFSG6cI8xf0YjuC9FC5t0WcKstkMJIlAFtYRQKrlGNhkpfMEl/3cmFTUMyGKL1bZnrVg4
2JYNM3HHuj6BgBhdNqIEnN/9Hqv5TKhYaB1pFtJlUglWmi/KWC9sZg8ozE2CR6D9iwfVnsHBG41b
WnXpXlyp+c8pBiEGq0Y1X42378xz6FelPl2gkamUbb8I0o/FR9z/qxkjGlQWQrp3zbOCdtVKO/V1
OXr9xejL3mZKqQOffH3fZ4ovjUfVWosUX4lgR8wkOhZTgowKxtYenjvO5yqMmzb8Gt1ZZT+yh2FR
M1Y5yzVHcMNd0lQr+2rIBXQ5oUmvkQirj2+TMKcYQQgj663NK0PWyayQby4G2ii5UFisFoW20dGJ
b3KbNrAEbQ71Cyze5MXcRNVGy+tc7hv0IsO7BpIbDUGhafJSYl2tEz8uMCJ235Z2NoWS4ZyyjDKI
0+FqOpN9jOoP+3iXJvLAXckADMu3sBmhxruBVyty9M+xlEoYdWys9V2fUiB6ezIiQTsYLZXJ2cTx
ip3wpDoLuOhk6LH0IN/ROQ6o+4i7VB5MsPlfHgegc5iUINFo6EHS6KaaMlcLMHeuSfbJ3wuRZkF8
wL6Nu2nH3nIVBp7C6OakCZd7ot5Fj8DZvqlbcbVLBk01ecCWkAgU5i3q7Dyg63cUSQ8lL1vBmcoR
6J8HIJbFxTSbjjBOkt14Jo0uyaP1WbloGjNuHvDRC2fy6XmEwh9xo2YWOZa8/mFbUeizbLYmscXt
sHWvbuA8HwbSRKiF2gUq4d68bGMrb9MJGmN6WDYHNZa5Ps5eO6ioRqxUvZScbkyoOHquIGCuamT8
Kioe5dtqnGqXI2vdOsJnANuLKarEemZQdjDp1g4vQ4lagdW/l7dHgXHPWG7B81HDAxluC57+bq0K
u7Gp3kGEzScBb6Mwm0gd+bxPCwOfooTYKqiIaWYQFaYbhnAHy+9U72M+UXE3RdI/97q7zUXyog62
IVii7Q5Gu/COAuci6WryH8Er8qZivd9lwlVAFtmAWwRnl3fOSxwcK/eSJckGqGXjbebPobyUKv4F
L6mPScnTDunxfe22TqTpG8A3krItWqsZhAfclwFlizu3Nuo5toSSJ9M97CNoU5Nru7qbqaIQ896q
DhJ9zk6EOl4uGZLzUK2J+6FTUADiQCXzb+arcSZxF/LkCLeCA8DzrhlyObxfRG+/6ZDCXmSlml2F
w96K0V0nbL05KRVbYTYT8ugx+iML9J3oZ8KHrbXotbMuO5fJvgKAtIXLYYzoiK3peCDvvT9jE7ek
UjITrQlQHztnXxGLxzVJ26CDSGZf+fbepjNOyiLnE8OuUE6SM0f6EIMfN8vh6JbGF4ps62nPVVyP
TOGUqXTXk2wHO/vVfECNGD/mIUnEr6cXpvtU06sd3yo9/Eoy6Xh2RsiBstyjOTYKJcsLvqxSCO37
/3Z2ZKPLkYkK2xfhc+tAEpf5i3+OPjvQezP55BURNKCDjyIQsnxPA7Up9ZNhWoL26yru7jB7oyNR
NYw7uuO19a9lc2m1V+d9zA/NW14290lu4f1sQ256PH9ZMXlA+cQ1giMcUgyn+xJ9+a8UMpPG+PGv
/7WTiIHeDX3fCwziYo3YSCEcJfNR+ULIy6yZozRyVpVZooT+mcqeMRyOaqnrDZX9qzbCSAZUC8i0
NLan8/1NCMZHeLoMeOQSMjPZPONkZFsiAUyizvDT+lJ9+kR7u5gyQ7wV7PWk5JnUFHM4aI+aDhes
T3Cj3Hjn+Bxoy+R4nq2k9pov5QD0lZSV+fY+H2vIS36ESDPNfyh1bm5WIMUf6BxLOa3oaXadZ8fT
ecT0fUM48F48MNbgIT0sKu4i/SVem6A3GwOKwpkJGuV2tKK0MFqKznAqmNpPDxrBhINT37kCIIN6
O2F0wv10g1mpLeJ+hlF6sJK6T3QgC8E9v6XU1sSmM6MSxBQtAV8kX4b2bMh104xZxheU1Pv6/Iu+
vV+eM9c41Lf3tpQp+GxGopodl/Gy9UqZOKQ8sQk86xcFeRaPe5fPOnCoV8yI0IrEJmuqAOHUytrc
1/5yLCt7IsYgq8GIq8xQkHXFKrAIfJWKmKYuFhL/uGywldanawl122W4PT5bhs8fSsVE44qO5T5L
82vG445nUVvDKDb2/2H7cBmvQZ/2OH+W8HMf+fQ/cx00ulTeb0EzfCZCd0FHSGvIjbapjGxQRg2H
89n2c0T+X6hWY1ascQGLtJV/YPyEWH4eZ0W/MUBOyO89sNPa/QqifZGcmlXGvyeZ02emTSu/LliY
IGtaYoeviNGkomkvKL4akSuQ3vd8wCWUfAzMqsdTrIvHeVkoyDhMxVEBKeZEsa86l4a/nUX1MM1n
YPEM6YEhO3kY6jjeM1xXgJmXW9yKS79mLiUahbdMWLyTfxkdg6lB7SOs1GAWG4NB5MuKa6NRqeel
THv4a9ht9LuGe7WH9dUWysuTjCX7qUR763gmZX9SYeuJqQZAuYSe5SKNMH0UrUrtoA9DDTHc+voq
CvlL5hCM1h5HmlQu2HQNxgoMQ5V7IyFSVZMVqaA8VSkK26zjqwX17F3TAbnOuC5JBUBRe7E/iZTK
3rq0Iz7WVsHnl4gPKYPx8OqrGqIZq47hFQyH8U/7HlxpvmemATKzolG4kVTyJbIddcDo0uDFUDfV
6yFJsfU+Hm6B4YqhOJGKCfo1++HzGiFs0NgpFtIlNy1T7Juz/OfAqsHWmfHSSZR1qs1ZsJgYJpSR
k2h/a/o8zpkZ04P+cw7Xx0RpYAPbGpgib9NbOzly2MEfDsPm/21WTkyuSqpje8VZjKHu+u8kM9ng
Uivgvz4YrHEWfRamkkkz5pjcyJSm41GBN99mZJaQ49oIFyzn7UU8GJwHmDTuAXRLTNZhSVefY161
2xJbMYMWuBduNzEHfj4tZjqH7w6jPugBbiG2dU3J5P3yQ2dIjiKxeq6jKchydTJSe6G15JeMcxWS
W4ATKdWZ2rHtXkFeNdiIFqwi2rkL+zn2QX2VYSwXNg5+AKot+LDEAZnICMf7pL99F2EM+l7aztXG
CilfCdLo8IAu9o3FZ4F+iYpLVAXdf8l8Vrj/VZbrR/mR9MSvgm733+tE0FQiyZBPC/aJCfyhw9of
jZHowCLDwqZE5lYBDHPClt9YlmQzBUs9jC1Wu1PVwY4oZOBQpugqDgEJhIW+m33BVqZNTDLu9OQJ
CCUYwcuTqDDfJ5sFaLOBAaEqf688HU4mVpnl0cw4YYlV5A8yT4lwv3weKtz1O+myK/Ep/dh5rIYc
BC47aJ+Eji8JyLLG8ArFnilzKOSpofQ3VFtIDSvpaFOkr6a3pYc7wPvHKUmLVhLNsadNTPF9S9NQ
XqiexLIPaYqIt+J9DeJj/iFLxqM/y3UKReW1aoEYEpKxOi3/ZzFg77XWCYhYzpQAu1NZ9Ijk2BxJ
IUgPq9eOQ5bbu69y4ZYDa2cmDND4AP5MHJydnvWNaOOxTKSvNjdeqp4KIaBCnYifLWaEWaSBxcHg
EtlLRgE3u3f/3ZNNqrRQxnvh4a/SpjGGTDNsmBmba0W+CLHd2MBiUoLcUZeLtDBpxXVrhVD6MSYA
vltal5n+a2yo6qR3AUfYrwiZ1BBPEK7YyeWSOjm+VybrgjQOdHLg5GRM6zOlfAdh9ZJ7AuBHYdsJ
8kFzjdLzdR57H6KmNtiRk/1JDnRBOSru6ivnwy7uzQxVp62OSXZ/pZksatsVdxNaD2hyI/glBlGV
LLitHTbynLT/mT93PPmH1uVlDgElW9rWYvVD9HTjbs520LSOPdc+KYPF9ofK1Q6v57Cr74/DdIMu
r2yhT4g7KzIHl7+djdnecFo3ZlWpnc70ksHCt5+JaWL2yeDCT/Pq3ZDal79AU7WqcjZ87jWjklVk
JnHRxGgPIwybx46ZhA4xGfZf/4VsVwfq4JIxR4fVCSoOS7BZNdIRHqlBL/oqImXSqMumetuhJDWb
cGsiKKDjWcpbbM+ou/MOUZhlkA4BKOWI9K9/z+V1XaGaxI4RhvzKsjyBgVQHSu13xk731iHb+Bxw
9ZheIv0dzDWQBg7jLRvxPDyWEwh57oq2E/f9VG2H6fQzxu/4b7RlvXcJ4aQIG5xAz7KVRuV5EP8L
shEbf3I/PjH35uKhAX93Wv6F+BClPAimjx8N9kbCWyhj1YYI+9cMPfMRGGP9tNA1fmDGrzgkPozi
6y+nbE0gBPGRADRfCngkaRZhc+EeusyAfNp6ZGl9YTW6nmF1TRekHd14WrbQX9mLryt8BwqgQ6Bj
MHIbVPOqeUQ8Con+kxOwzTKP9uBkC+YxgIyLQvGR6YD9W/6zNnpCGFWdOkCGdhO4lstVY3rRumb9
d31pM2HfaHWKL42kVzaT2JSYFiWWRCGw8uRv6n6FQGtfMfK9iww0jzAyD9tJ2aQ3BYh7pY2ewYN7
QirH08W+gyvlSwOhPkoDOezbbU0FxxEGlR5NU68iKRGSZXQNPLBr5r4QYsCaOVH5ocSmgURkItvd
juRgPtb/MMb+qNNa1gEDU4v/plirUcigAZeSfe4qIbNT3SR7sFFONvuvAqfUgqw93Gf3fxgjyBvR
16hmru5vHtR83XbgidaIgxaLvj7NjnuK07fKoiLa9TjD9V0n2mQUr4x00bSpZup35fCBKAFy/jLY
jrco4FP56grth4/7tDzQAUwtyMnqCP+G+Nd5cwv26eztQi5Cm0O99fbXPuTxSoX2luOeiSzTtSh7
rz4GXKi0DtizYkyoIVAolYpswEMg4YQzCjPk7+hK3NkWGjU24uJROk38AIusqxJ+WMZNj5+VF1d0
97hnCPOOvQ5uE4tHrkhnx5DMWbACNkZ46W8PrJlKjiBq0cjNS0FP4zut4xMm5lDZel5fm9i3/2CO
AAu2xWx79nxw0or5ANpR6OlkZNs7lQpJYseKTbXdgRcCsF6TqLKi1a1rg+yd3DILUw0Qw0nD8M50
IXnkN0H5OoOK3SMlDNhbuymjsL0AUn9BlXg36ZVTbXLa8MnT/DhPLS9ZiUod8QG4Ud8HFo/giwYj
bQFs/zwEpZHUU0tQKCnBvn9D0MKO9dCKCRIvgZQZ3iAsIej7FkU/IQuLxvlMk3iBglrTNM+iVq9C
o+0KjpvDuDeYS4Tx4p6rSiQp+vlysvswTc/R0iQiR/Zn55AZ9zEpr3aJw8+YIpkTe/txGMn1Hb3X
CL0toCdmFqsz5zXA4Ud2hCj6O4rNxXnC2Oyp+TDIRcZAMy6cpAa3PL8tObMsi5093LX1PnOcwVAo
vRx+9n2B1Zug9SK0vQgrtjZr33C1dTWwFTeoluMq5pASOx2MlpDKuX1sUK0nTjcmcpKY8AC51Hew
gfPJAcuZX3Fhi06TctoLQlN3OqsC00U859mySbB4qsEgE73LQNyAmj2EbPWib5bl8WnHS1jV62q6
Dy0NBeggRm0agwgmDlfAnGMb+FE5s3ylqwf5Ut/QUs1/hqLWriaIzuaZr8+MRlzS7XTbadHcFJ5h
W7b6tywpIHtrdn2GvXSxu2eXM97EvdLjSeG+wJeubF+01MxD53Rw0xVAGTJWz9r2PtiZrsr5oRhA
lrOxi/4rh/X57fBz27vB8FluBITbe2iVhlkTE7FwxEQtg99KcI2b2v+4zT/p+qPOFY3rnZoieVtt
uDET68v6dWqheKBnVnWdSBmus0yXBjB9YzrBzjaTLs4gbQnS0wA4WydeWfVzaCGjU2GM1R6uAOlF
w6aPY9DfXx0ma+Ta0uS2dx/mJLwc/35yhRKGQHGlipokYJdTMuV90n8Qm0OU5hrBwvICkNATipf9
HhyRWKkwnaywsDE5oCIiPTl9xAlbyg3fbnBTtzmGIGhITq8TmySWX/gPmXsbbZMS3uh+17xPom2w
urTgJaBNZopnG0uyuC0tBkd0MiUsG1F0ulL4Phcb9gq1AeCnlNAPLh/E9m+9oU8OHNCeupTzRs2f
PRhDlgR5CNyT3iWDQ92yj1I2rwv32Om33r7ntS1edlXofDRmt5uakUcM16BZsaedeyu2P3MsEKIp
+GTG2JksqH7rLl1CwXdlbiwE9dgdel1WMd2Yxbrn5qyZZb/S6qfxZDFT4kGTfL/dtgCLClMetKZa
OzKV6vDuDqZVbQtQC4bc0PAxjwN/83JuTb5laEttdjYFxQSBpjl8az+EJisGW87Cl/NJfF9BugES
D5K6wzP9wlkLwHy9CawwNUy8swVDCwnvfeHnRuaCjPT2tRkjRqV8Vhr6Z4p3yAXffPCbhBBwYLnS
tThQBxc7ouPuCRu8s8rXgZ2tw8ihOycIz1Hb4oVmpSTYxr/16cszqkd26YF1Gf3l4Ttg3WnFTLQU
uPQlEZSc28pqOn1/grNj7643AvbHhbg6qRWEf3OsRRC4G6P5CyStuPuqq6dKEaYzZLw7nC3BwDAw
SdRFmdUDA+HDEdsxDSpClR6ZBk1ilm0yH3GcJ1FxCnI15IiESW/El2ArN5erVNY+c9EYXaQ/a6GL
EevAAkSd7wl3wGMA5sh2BPlijxLXPFtL0KOuem+GGjM3pfIg2lCIp/oD/ArBDDetpwomX3HMFA+x
QcA4KeP8+pAZAn/AkrBHaAq/evRZMMdMZGL6dJttgbicRu6ppUnRaTf+TE8yuFuyN4mX5TyoEZTW
ETrYugahh/bhlkfI/v4jBEa0Thjqbunub/MGPw252tdc5mQL0G7DLhniU0FrobYQ6zHeMkDKkg8Y
38kuAHsnDwJhncxQ34Gae5pJD5Y5C91BHd/eziMy1BK0TCcGCKukZEkKf6TomcBAkn1PQdAnjJ0Q
f4Os+eWs/Bo2Jb9CiROimKIBdXCU632eRNlNFNQeQg4K9xeMJvPeb7ToJbDonxAEROFjq0InGzzr
5XTF427QBAsdcgvOaFM3/bBqpdbvedqJUc3LIVhhrVjAcLoSJ3pLX/AyB/UrjGxXTNzn19665D6D
SvqQLasp6ZQpvx8lCbi9hZunUj9sVJ7FWgP4cA0rF7iMktQguCLBeB8ugzFRJhKrUYN95lqP5hNd
aDHDtDa9Bur8jFYi4pUK/cII6tAIU4goCnPGawKCbDZhqoJcNqHPT0ug3moHfPcxzOJa9bE6CMdo
kC8KSLzKZu1ymGR7dpEo1wVlZfa3BPW64nFD1LB5Nl4xRzcoj898swkxtYpZlEYQP5m8PblPnu0s
ErBfn8gERTkbXv3mZqw1qTM82JSiE9afZVVYBOt1RQfiEWJS0FqhCHStS6Q0i4hoa/KDDfqCyKju
+e+ci9z8Y+JUexSALS5V6EfH2GEDSdL118NxzXu3TrZAyfppbAXM49ZDxMznblzojtDrxv5/+2Pm
u8DAW9jBOBPI/ZjBDoEHahHnsBKzCCeTZs+r/SLU3d1gWeCzpXsLiloiVzuf9+zNLBUV93CpIp/p
ItJismW3JUdLkPIMtkbe2ZRu2X0p9+Mr2Ho1RBd+Yv1DRA7eChTFeRjIUSsnDyRB9HwlZgCqzB6Z
cvaXe/mcDy9JwCd/jQ2Wg/MAaRvNaIXpJGQbkvIig4NBkd4BJPSJAGbsky4fURP5Z6kmbOQ+F6wT
D9Sb8xROj7XC7Ba3gxRea2UE5nY4UmNMNwjO0c1m2gxxgltF8MV2iESZrSANGWh/WvOhLnPcga/u
cQBl4oBQpcDI0NzTs5CNGYFBqbEAfK1+1WdHa10z8CcPICv5NzvkpyFch3cU2DMkj88tMSlc4p0T
pcCfkbtIxw5maDN56nmSVc+0L6AU9SqhMtjCA3EkSe++O6gi+bpPlKMjrhw5fM5wGPBxa3JATgBC
UPW6Gg+y5TLVI6C07tXQp6i/HNdn+BslD73CyUh1C9WuAGIa8Pv3zDIAjdI1fXzXKKalXs9NCmG7
ruV6ufILUiNbTbWPSJ9Mso4y0EtiUQjHH7sj3bSQteEWDu2CizNTLr8srC9aVtemZwlZOwjG+bSg
HE8L5nD6lM5WkTF/ky5uYTbm9Fy70KrmOA4ezFG8SZ8JNa3/ze5GTkQvn+0MPz9ey57nWbMJf8wV
+j2Q1aIWodK0u1NpXAY8TiOFy3lQGZRVN2VQAMarNoWPb3WdP/L6awpNLbRRpwEqeVuPAgVnuAq/
RQkHe+gcxFHBhU3LoFgDRCI31aFf5+o4xPzwf9dBQC65EC8pyZUd1Z1iTUOscdl0rtCnkGalZhuf
r6fJKOKfqZzW2l/gybikHhTqiYCImDs0/QsKpyzvQZivG9CV9mYQZwMT56Ru6sRPh0YsGxMqIjAC
hngo0ywHRIiu9wvLkeKKFTRzkCPwnf1q0LtavSvkSG+dsqER9vxga4dF4CF0ZADoEgL3CH+9+91p
ZxFdNT3Sa7U2qraZvHK+lw9F79X0FnwSzXGDNyYyExImbZXkRL0VVEablYWZJFCx3kxCFgUWYZDI
TujE+AzSbHGbbpONuCigJn+AP57SGDkt6mXOeKfJkpijGWZyJKoZA1leu322PUGzY2BbEtTpNUbW
BsUdf2I9vwaEMY7+2HDOktLwEDigtf9+rFtAodEFWiQ9vEvT7EjK0cazyJF/05pahGNvTNSWoNv5
bN7RAX9IvwOdBCY6tcI1e7blgwr7qAb0SblPhejdGJifJ2lNXZ60DGPMsTqnZwCvfYkDJsTcBxcM
wJhgUBY42t0laK/hHMtkNEpwNS8lem/fzImfYFkI3Bvnc7aWaMhTju1A+vW2+yvG00f+c/fTYaGt
6F0YWOM+hYNqioZs6+XVuwQAmUh2Veh15Lh1UDlqgR261H/1TUMKnMwVPOKVEpX6b4aP/RVHJd6B
R2ZFetH0DjjusRXpNYxafzebNbqo6/smM/uphfTxtr6BMRKxIKZEch/Zuh8FQt/ZxMi3XlagZyEn
Jie8VTqstk6YXtFwfh6d0ejWuUAz2l3esELhEwE2+CMBGtMIq7u+YHrZcHxK6nPL0FhUFEx3QZ0l
JkIbWThzTfkbZwROiiDMVYzfpL2UoFvpv6Tuhw6xdCG2Pr1O9b/IVFcenfLeLvPYms6atlGleH/r
c/kRt7N1XbZVlFwxslyPDXzAeHdjIRuUji395Zo+XGZ44aIJH1hg1JmNVdTzLJL8yIuZbsOLA0nw
LkTWcaROXDE1iuN1lFL29K8KsEiN6j5JJ99SILqtOSzGrR+zwIhGpQFdH0Uu9nLx9ilNoSjkoI+L
MzY67hMJqWFczG0PrnOrtkTnHSyYGLJQsCsuRzS8uQabS1oe5rHWAltpzq1fa/YW+0dy8RfXam1i
dAveQlwUJCB41QgKjzf55ZbxGx/3jIvZ4q/vyGjrKT4GbZJX3iS2f0H4S3Qo++wzQEF0U7n0urKL
DSOpjuqNJcex3XiTcddS9kPW6ShnGlSoi3gDQXSUDiCnI7ChxZxbEDzbdjw0TsuJPxlB/73rPRu4
WOLYiHyrfDINPHNOCxlWYDxN40X0UcyyeenrBwnDz3Byo98fVDjO8zdKBhisn7PwsMoFe2lNklmX
OeV9rN1rjfYd2NEB6IFdvqcMWQIWSzaB9uRZa1ygiFGWpXnxRZrhU4A1qJvjBC/4er3FDlIMMYNm
hWsV2fdG4LQM497rBWP8zN5DLXDPJPjqo5fE5/NQ6GIvuj3HCioWnBv95J9PIEt/mYoSVFJptEIo
90NfMAxddpe2yhI+cadICmJyzJeDFhyfgbNANri6yebspkPvpbOmlST0vWfY8089KP2/2uq4fW9J
XDoEuVPusBKe0TxbKom8NnhQF246XfKsC/KAgOcJO6eYMiwivGJHlnjJYQhof1AsBeNAfqShOwmP
NsviFkPJCFuAZbowL5yZGFW/o//Ld/JtTtAcJbemOIFwQ1QbeZP3Ilfdue6f8qEgC70XpkENtAF5
jixGiHJG+0T4o7HGvkgDPTvd56VOMgIWpVbRWVON+vqSR/oEsO2Lorti3pKQgAkYtTd27KKxg/aO
CU8ObkcNzuaeysFHC1y+1wiOZ08Y1mzTA5T2Rake2GrUFwfw39qdHglbHSHZA3L8lp9GapdVV9GN
291hf2jiY5xthorQZsm7crjddBJ1amsCbOp7R7jLDt2PrDvukJs0dcBIaP+MYDZq2ZbHWI5LsEd2
M/VSkhvUswy8/zpEcC8oftSA6xhqc0irXu7FC6veMaVV41H68gySgr2XCBiXVTboC1dIiWfIQT2i
J6fWGJWvY0n2Ax/GaQevuK+jitq8JFXxJE8JazKvov5wpKNzUK1ag9lf17aTe8tbHTgMcx23aIyn
bvjbkxPDNZxFxBFzoiECjqCYsHQAS9gHOlhzwY5Ol3d0gW606Lr0faN7xxioX3i6YIXLozWSkC3X
yPwzLjhNS/QukNwZ0Lhj9b62XGTc+JCxIkjoEcWyGXnoM5PJnXD0eZZNxWo3caeWUj5j0FKBAsMs
Z1+oxHXlirde2twVeUD56XsqH1mGDNn0RghHQmik9r5OuBDUQXGqqUJUOsLXQBvpoKphWDak+fmh
kZvrTLHVLQ1s2wUOARUVgLRybLuAhOtW8reiAGo1nX+Hc3J0wN4Kt0HsZQG6hBGNOMX00RtQqtWu
NZKpN/b+m9ZjYDpU2/GlMABv/QMjP/wDy5QewwBvk+HH4+g2TO4Ui2v3kujVsb/3aaj51+coIreU
U2ZvFRip4/rXWzVlFED0qEYf2aQp/00mzjV8iyChdh7Bzr+9TqLCgoEnrftRtSWAKZnQraUt1lLj
/t/1z1Rgs+MV4jFhvupNN1ZvAwq2JwpLrsvv9DlAfOR+Au/2Io0n7THtVkYGPd2pGLWzNSt6/+IJ
649FMyi6/ATPmzHjgqCQDzNfr0Ke5rje6WcwC6EFScP2tNCLD7OwRtW10aA/DhYA/6kZTAdIYyXN
v4O4WvSn2z1RCIgTt3w5NWWSsmqwHNY0ie3Xs7m77z15PrHH1xp6X/jcTiiufyNuBbX1bbLYCrEY
VPbcM/tRNZ73gjTF2xr0DktIJjdnrDSU6OVzJ65fwEAUC/RJyVF4eafdJv+9dpH/kEFxKFxuC9Of
JjklwVGQnTDFy1MTuE0J0hXW1qdLANZh1/MOgd5B8E73AXTsXlz6OJjAfAUlxD/2x3tLglFxbZN5
Cc9lhzlZKF/pI4liQF6Ylpv4rjKM9Pf/PzAW+JgqWmO01I2+vXEUbiAIBJZqnkRqNHm1UEvkuHY4
KlUhkoj0YDDVFXWsmPTIBjevDyL0aHdFFwn+BLpMJcYJaIWixsBT9MbbHE3tAC9n7uTRMqp+VuPZ
oE0dujCaKv0xJIaJvdn5WfZzmFdOSD68ww9mX70aSXRWdGKsX2sdsuswC6Jta15K4Fvnw+Z9fuOz
vdj0etEs8tbKmc+KFEhBVX2AR8a1KtQw23OJPfPXGMMZLAmbsVMqkBqG301XoI9vmzWTcHOhEAxY
12WQDO84gw4VvBEBTK2Wpxlq7H00z47zUaayYNi7+Dct+02+xIO+mw25IT2mb7A75YMzswOD47oK
RascWzHVb082kGCEmQ1MHyM4xFfz52RyeTCcrS4KGH6FK69IEVi7WECoKwyljYA9ziJ/b/uQjIey
QAopuYEJM4otZ0W1JQBuHhzwZeuUybobHru1D+dg6/BXadd8QFDGhATrp/HOGx1jnqhwFGvuTXNA
VNwufMQorut1895YL66Tf3WEPXbTyPtZF+oPkf9QqSKRcGYt8e6M1hmmPFydqX0omh3x/UxXRndW
0f46qDUgwMOn7v+0/OjH8RN7ReELk5XYdAM9FDI0XDEBRbYO66hPvJjTRnNq6WPzeSQpalYikEU5
d74/sRLfy9FerAVj8ssxP8p7k3dmeOypJ+SJZsssmMCzjyOjAr0FB/dHNV9i2zbvdSFUmobev6Or
Lzs4YghKO4oPRtc0jxUk5dYj1MQKdSkQvbRwP/O0ofhSSbveYZkvuV4CinNTuVTTZIj0lzwhnlsU
X9NmaK1qcMAZQZSV8Ki0liDsRY7N2HvupYDPtxuxRtLlBpc1LICQwF+U17S16/TaTAyiafCqs6fo
aCpf1M5dlNqXOsY+0CB2iiR6W1GgXL2L3z+Q57a5XqAQ/nrFpNi1dBKl7pwwlgRU6fzNYxQVd/Wk
U7QQXJfjT6PbB9cBR32tEORhc4lynQ79oi3yL3eyBtHifBmWd2NoZIRUvJLr9p2sAi2SahHMjoHb
MDRry6YzkQynBPSJzmc0I07YGDISE03isU9QzogG7K3sALfxrZ4u7L0Mdh83FnENElrgnp74qCoC
XRUvIEbLjo9gWNPBGgP9oNWMR7cFlW5RoHYGfU+vmENEqhXMKAX7MVGGkVlGhW18VSTGa1g26yJ0
SV1fOn/km12a2XOFyULwvBFe77DsOjdYyo04YBf8WttDRmuICCgKPYkX44NITpUOczpVUVqh4dJH
due9eAZi/IF4Fq8lsK3Aoj1ys1zkX+D67+X1lMQ7iLPI/2uzamURTs5aDfiqE/OvacB0UUcBhyur
UOwSfyoIn3Sqi+WIF/HYBxcRFdMlA5Jx2lOApHF613IDd0FoGDei2T0EPzcmZc38BkZGNhNfnWad
7Z9HzEQ/l06XtWPtVAhsCmXLR0Ff3EedQzxJf6gSH8GfPRyoP0CGVfdyxfIzlLUrgMjT6NFBLCNr
gAGBIseV7PNIA9kaliR4pY4wBWtFwRIPBzNNRKn56Jb/LuZ7I0Tkc5p+5U9h6C+LGJLODwIC2eGQ
/AVGhLmeCtGVKzjJ8x5biAuhIUNsIIQdXug6Ssp+1GzI4Gxjs6qSEsE0upIvlc/v4MpeK7jFbZbK
WAdIJx4/FfFnr6P/Hcu+VJm5ClOK0/ELATQxMwcddTI7F5EDnkpYSPLhgL0LkN5ZVRoxXUMsujVE
3pfKb/BC9M81XT+deLkiChqj755rmecHKeDemZRK87tRDK6aVVeO5xorcQ9Ls/tlF8PXpqymI9v8
a8DV1TNlwXjDPG9/rVK/I7ymZpS+s69fLWUf1vd9MR/A1hrnuw8g7Nzw/1O3QQcXuGNU+2oXzBX+
LbsZZY9Ls2UljrNdGaleCCiWZCEKYgGUUDcR0E8+/9jgk/wZAY8eh8YakEDr2FxjHr5tGRm7120Y
tbN6+TdFFLiWbs05lKrD+OanGvPUW5KABkM1CklpScSxmRoWOcPA3Ap63aQXvZ/yEMQMj26LRDB6
aVCptUEB6RzA6/ytBQIusTgFY013jlhdvQrG+LdNWs63+CxA1w3rnm1La6CBOR5A7ql9jOOs6lYs
NOtRwBrvF3zR29I6Du//I0qjLsuj4h8J6WkO8L7LL9W/2YFBrgNmZWLOdnsGqi6LPFrKXWQQMTgm
Ll2fVggapUH1Lheit2nUIOaE/75lf7ooi9o1q7BPVCXZb+6Q5YUlh6amIL5gD+jTOxZQLEDVStU1
fBfqHBRsLQBc6Hx9h4o/CmobovDjxkbAXO/jplhbjjP7EW/L57eVS/dz+yduB12tahT4QIDBsHO1
NPQXnRVqC6bfvzOmUmAZXlSBL7tGPjfBIk/OqJIZl/Dad+jGRWJrwaZ662yqnmVQ5+soS45TOoZY
UxKNn0IHtqHYFQSH+sHKAAXd62O26KZZT2snx4ykalZmhr2j4m1UoUwZF/SIyR3m43JIF6eBC06h
40zxhX+yFbtNvj9lcpcOkySvi7YGB/1iQUJ4n9B9QQHuwzQgk4AT0sU2hhYwScroIz4vgKhMJ+Wj
r6zkk5L9itYvtfDXZAlOLDFD64V6m02uEOX/2XupxDqhu1qSLdfBeq2V9f/gezAvY9KOSWHuZ9IE
4aN8SLzl5Yb75GR2o/q5oOVMcOuWBI9E3QIF7jltCzz21BCZWqZC6yflGXgPBbjiPp96ktTtPATg
WlgEQBhXhP8DTpitNduo7j7ABuuoMGKKrGG5YjJVnuQ9Pq8ICJSpMxaDAyCHZYcmlFRjIsM6cKkQ
Ph5YfpZ6TWquplAACjJmDW5StTVL3W1bj/kXNE1qeE7Q8z1CJJe2fASQTj5CAOyGwd5eehxnLc9b
Q7TrrS1GA9GUWz2kMKAheRDDoT+E5HKEGkIBst+i6Gc/EtLuNvxX8wF9+dvEotuuidk4rHLuSsEi
sUPF5KAF1jPuDp+QeLjThjNvmMedqiWfECo38HN8WOwTYx4jStMNxsoK4ii/HLKFNn9R/tEEmPd5
0qlvR6PacLx1lLFmG8e3CLSkY4rgMkzkxStGyIWt5S9SY5ZvPrY7NWEd9Uu/OpRVahBZNA8Odhz+
nzFaUKdZdKLLPX4ZOBPdLvmNioMKTrPo2a5dJhhoJwTzRooIImU8aJu719fJW2QjztLSvwRzYs3P
zsOpF3qF2bqWSL6YfgUshytewexy9XehLlm/+oNoif77HQU0QhK1zKt8oRmDuqKXoM8GaehO9gwE
W2MZZ7g6542Pi/5aj8mSziAzzihpldva88us33O8SVTbORdo9Rdnbx3fdWqAPc0f4eD8ZWznFJq5
knj5TDjY6AcsPZpERObSlhJYR28v99LOJ8C92brDfj2mT2iQ7M922jFGWxyw4GAN/gGxpRggPxd9
TMuzoMfHKjySFgTgHkcPWbL0e6LwbbynqaBpiu+SxcbWewRIhmxv2mKDXWsF3jYKWodB1CqHqj1Z
u5xZfEZluQT89gRUKpAlF/U1isxkVvGSYR7ZtV7yAtSEnpn1IgfrwOYA75G1IGJkqr3Gi5Odjo9R
hJuIvV8fqPlTZaSy5jAQACaBinJ1G+q7j/tiwHMYCJ83VuPLYugU1QTLzGWYU7LLPKE0HQ+7Mx+8
mDCrVBTpLmuFmT4ohEBlA2Rt5Vnu8M/Pn72YPgJWzPqvsniacMK5lHO8cRQlT9ngOe/fM4KHumnu
MAZeVaD73DMcMh498Q+lJ4WltUy0XsajuMKoJnQK73OHs6CO5yks1m158A1cWFaUmbbdLGx9aY/v
doA/tOPxZIk53KIG8U2DhAprl+DFuUlQXNlD/Md97vrh5KT26XZS4fsdo3nw3P2WM2/KRQAysJEk
dNXWzTFF2qbSVyMJGqbnoG/DW5CJcNz4YvQBp+TvmbfsVrtwpTT7O/vf136Vu0aclHTGdPCj7awl
eVpqizC3Wm/4stwytQ7tKw43ZAS3BlGBMU1ilMLrOQRshb7g8GRHg1zBwwFV/PBRo+HlsfAgypXG
Ojaf0tVVqYNRDi6fPzQ3GputzT/kM3NWsf/NOH8P+FNtG2qBBYSFQMUT7+7fcPZ+uDVKQaYRglAw
Mm+uKwXMFx/fqu5ItvtOiieLQOx/2yrZOl5c3GTs6G7b5z8HaI718or1BM5f7F0NMIYnHBIVijEl
xkCS9VLX0WJMv7zXjrYCUJehf0kxwj1TqfZHv24Hl+kuGhOijpz+TTAYDvHKSvzCBG+IyN6L2uWK
o5xwoilHNkTG1tTWL6crLM7tUjgb1/IKHgTBV3/zbQkZ/KfE4Tbc+qfR1/GR6eopA4JWfMMMDUXi
+Odl2UTASdjygnygHJOwnK0LSw9Gn3lKB4Km6bTh67K3rTnOhTp7CZH6gzH/sVK9GGwxu7hd6jdp
J3b5sGSFyIsLTDZu5fHStbi+OPOgmxpV2zFoeWXRw8QrFJSgfoOAsAUaLrRQ/7EgtYt29fDciI5U
1dQx6rgveS4POmxlo8KIxA9MqeDwVDogf+PoyqJSCikPidjLTJ9Xqdju9pu0MuvHOFgvCFZd52rG
7ZnEp5qhts330S0eeG30gFYSvaIx/YfO8X0XEpSJsPbClYkYjXD0GSYXzQD3z5vC4cOrpoiiyCMn
DoKjufV0/PlC0/zBsjXJk+hgthnj1hsa2BuwBfOibdbDgQ3lHUeJqNwG2SMl4KNUiiggveqTN86N
Tuq5ue39EFw7erMtl8YPvG6qHiZW6taAz9JtuXIA+lJ5P0EezZNE4p6bWbepyUy86TSVUDIOUbg4
WV8iI1iCsb5XcelFa34fe/qlfA8Zw1fnL76ODVr8ljA6qmvihLOX1ANY/vrCvznDSreGPd3op5wi
LOw7ZMuno4SZN76G5UKMXhs9QpTs7XkZBYKugZ+AimrulmH6Lnx/yST6rLVAID1R3FfTs1TfBBhh
naiEQe9qVIzGS5XVDHBWmiDIvlsLzCUlTanygz4eojJdlOcGycZKYnnFchQmyAH7/CKzIEJ94GfY
z89DhQz3ip8FI6KmFWbdBjvxCSB+halnp691V3+Y2h7Xbl/uoMpShnbvZuW3RAPP64nb8gP/UL9j
fDMnsvQuSQGXRiRR2erFgExtqM1ufgdVp0LCpVniomE6rdPEoH+Xp6Wt0oTmdB3pN35ksbbX87+9
I3i23IpOO1hMS+6IBbdWbeAKenwfTEKAksKYhGlucZQ3a6UhYiyZGeakF48i0QmwKQ+sHWjPyAze
EyDxqLPyvkMf+68F7rOA5bZ3j4nQxAgFt0qdqpuZdhQKtTPBnV4lZmFEAi14gUu4wQc2apF+k1Nl
woaI74McaLiP0dl9JMufUB/bDiTdFYl0KhwIYukPeqgyHa9xv8Y5zdeK2tZkTJ9ieVlVBmtcSJc2
jyPfaSHgYC9P1YrWOtFvHoC0EVCRZI1/zHD2bv/amouh9DLTCnUgju3tgp3nvSQe6PMyYfFdsP7o
sV6+k+DJD9sCuWf6qtLVjUot3hV1P8WVPi/Z39FHrrRPbVkS8n1+pAMlFJtSvdQs0GzU2ScCiie4
NklJMB1b+6zllkM7GED95X/GI+BZAKC952iNSHWfAHoNv3V7TAAJXl/0Hs7m8rtBtdDL7wU4+EFY
zf/OapM/UvzEzPxiEdxn3dyOc0G4A/cwYqVMD5rd1ifjsBYn9XkQECxYBfV/uhkmTHlarTMpoOeN
2ec8Hga0ThmZKJvczk8Iki7gOld9eN1avTrC9kw1rSavIlPvqc+DrV4wmNXrwVr81O51y4A27dQt
IUruojkDohX8zoLdVyMEr36wvVVMdZe9FVNbBWqGbHaywYyHvY2liXnuYU3vkbM4FqJemmtW42r0
H8M19KG2BvTsN7osF807bYGrMCs3T5irWLgdSQdmGW0IRQ9Lce10kwCq0MgHky6ccguBs2mA6GSk
pMqATgDfZ9cIei5vRUx5Nm/xdMokxGTKEwWf3NwQcGzs1WjoguYkkYEJ7pL9qoHysSEsv1GYNN7K
xKZKKOCfeyw+dwPfuUXDcWml7BqGQq2awdMqZQ1A+BpWuvUo73yqReBLrDjQT/DYePgihyrlS4dr
dN5msMSryO4jJVVMjI6U51Md+k4G7CbtEDwJe3io0emRxrh726OspAiUnCgt1dI89GynsQjdu3ZZ
rro/uldYyRq+ZmSwyfagAYjpN7ss9hf61LfzzmSsVEC84O41LMpLx1pmVNAC6HFX2W8MVlwGlC78
mMq/7ioXujZWKrt8HJSLJ8iW85scwfW9FUiY2aShLHcw9yDTedYpYDqLEhfPL5fA4hRcyUCKR5Na
j0f/I2CcEHajIbL0fsmoRQXIOVvTk++EkWh12nB7GdeL2LhE+0qULPZW3kfi7iTPfMXGhhUpG/sO
cm40gD5PenzH0mhosXPU94z4CuCk1VkX2p3QfGtu7CKFFpoGL1R8uPVjjSpfaer6aSy1haemIoCU
BrdDQdx1/rKSjeGpxokOV0H7O7vqM3T5E33DJ/w1CepMdtrCbPfRys58avZ9I1v8+bEdqXRdsBRg
JDbnqEXNo+tJ8T1LCBsTFE4bUKZXgFWn2Ioyrrn/5zoTkTmeV02GOa9r7CBG5SjRu3thHolb1bhm
bydHJa+Mf6/c6o+Gaxsz7o+6DvnBSQWid2JLtEJpbipfcsOoOVdsB4s1UC7oTIsobUmAFwuZI3qA
rF40h6JQrMaNetMRlk9+vyGTgWv737yTnxfhRnVSNZI0mwJ8TtTHC1l/gaTxWcXHc5ZRuO+JX8v5
RbvVu/LCb4s1xHLuyERfcTZWu+rRT9xjSdu8YEzlwgt/MWx9YH3kOL4T+Bt4XhOJYpVHeAtIbxtT
eFRkw82p9t2A8r6rYl1UsMLclJXyfz5TYwDnPfZGKkFwq23tYT5NhCu6g5fndA2P97nlUtUK5uWY
hUbSi7jMptEEx97NHgkkn7WROHvmdf3z8LNqGPRrYLxSVzf0EwvqFKTDlrF/1sgnAMwDJfXwfqtG
5e9S1AlR7W6rN+aUG2IePq/j0P8Iv8WBlphIqVhbwQzbi7yTMftlbM6V6glxW0mtiUw5za9j2iiZ
wvNNNvpkaxyiaYlvwUQGO5oW5si4Vjxmelmn8WHbOEThyQJdaqowPt57KukhiR2NhOh5d3Fi3Dfq
qEf8tOgPJAiVQ2Q2FcOBe6SKyifMe76gEdo/h+PhKBMLPPv/qWkOjXPxduK06B2xOjAxUbpiDH4w
f2Y3l8iLe4d3r1sIfLCafrD/6jikr/Rwk5vxhmbMk6rXDYvAM1aB0W+rnT1hkYH9hQh5zokYr/Aa
Vj2rc3OMEqWER+IELadTc04chGuNvFNYUqLx1Z0zKmmhr6ksSysDzXEpgmpXhKdTDIBqJBIOYTH9
D+6h5C83G0gNwBqy4HbY47E2srbPXCyft9w8Tofk0H6sl3Kw+kEKz4XUPAXXfyOhYqb9kLcHNEz/
Qj1GRxjcHAUP/3ot7J46uQrhR+NOy04A509qTUrqg+b21/4EGt6YS4G7dDRXiOagUN3DVysAqWvG
bt5MEk2wl+yKK01x4zT7SKUClZ+Hj4/tNk6089dllonuWU5uH0bXvhZoZZbGwsKEdihIKlrgROTk
KG2mAoctOWGr6UwaUuJV7wF8msSTlrxNTVDg+f7kBTICvlYsPDlve4CvUBEdP5WS2iP6pYvv7KX+
83vqiA0uACNqwXzeXyKyfNY4xgZheGOkn2JKbdx5G+RQo+Y3ZuXSOBgLV3Bln/SVfn361HIjN+es
DIEwEpvN3k6QWUIxGZo9bMCN5hId9KiNmAtCPM1Mn5XvZNAmJKs9MHdCaCbjWuxCvokXnwJrYtDO
uS1j0RFb0aRFWplj2/1R4tqGMJsV4Z/o+XfExr5vamyJncuXVhIfFLF73tL4ip7bPS0lAWruFlY1
tKQItnJSyN9Pkv3l2P5T8IoN5nT0qOpaeSsp9yg4Yw9z2AVXvD+By/F4AiCB4eHfLf+O5wYrjHin
t1zuOD5ktxBxFreRIXFQgcqonCeTqHofWiBqWw4d6Nmn7tlBqdZe9FHwH1VEpT2+H8KcwVDHmJMH
YkhhltA2k33jNWBAfRCaX5tewGK4973sAf0vHLFGJUhAbyzGQVz8N5VOgV5eL5HGJtFOwTbpzbhg
4VfXcgbwRHLeyNs//WNrOAIDd+RXFJcLbg7OWX81XnSl9DfJ90JUIi6Prqv8W7NuhX9aK+5V04H4
Bji3RhOQDgapQIS9Uv/9LbGAetCBlO54b74no5o0+hBaxJSfekyFCAXzi6Ti27HVrqB6Qx6Lfagq
GoW+LoYdc20obPdLJjkdIAJO3+OdIzORsHyPBchmLl4/BIaIFwjyaVY0fDO+lwhwjCpdlEoDLHpK
C4LPs1xk1kZ6e247HnY3+guw9VYcYgBSvzTjZeAvPjgidV0SfxSwcvDmc3h/asldWt8oV6evy2dp
bnmLSulytsR03cHO6f5laGiPFk2lwG7cUc320ZV5d1xICqABWcR/32LA35DbEeU77dp3+yn1+8ad
xh9d5Z6T5oArUu6QZsLDKPm0OAHQxxBTxIoXV3BfCt2edtWZmTqwU1jSz8z1/arrW3HyI2Vt0QCs
Q66oljnI8TvuH93KfGP0eleptPETP/55QbggcrJHJ6zVRlbW7RwilFOh3looGUrRZieI9Em4SPFq
G3NCvMkOxR5lI4ovqauP4KoknTBBuHMvZ4G7v7MWtdajNOITZT2ixylKAdxc1s7osxNg/m7sKAL6
Vu0RZaSk3L6Buf9pk+q/kbtzxo80B4ePJniTDthdn0YJ+3oR/3rWs/uVzeds//t4nwbeYjfegBgJ
7sA1u5K4JMYR63Qoag0P6s3uZnMeaDLjd7z7Gm0d2V+njNcXP8NI3nVAaHqu6FP8Rz9EEKCfQiaO
F2mEwUSFNCftswyd73wA1BWgY7Hi2MKp0oBDlb4gUoH+C2NIXarK4q+/RXabacpBm9em4BWpNewj
snXMDddj0KOJtz4rdmidzNnxwnZyUOsfk7ptMVxxWezFZgyTM85tAUJXUSRJjqqmXgRYRdUJOl8X
7Yzbhsnb9/Pe5QYK/P4YtmuizLfh5sDIdT/dIl3pGs2o45RnBYhMdcsfDmk6KAQG0VVtjLKmthqE
934i/w/KnYOZoZmIPOVcSTB93hJn57V/JOvX/6TmEuORAdozd2YmqcSFU+v0nHFOOm6aRS7lsOsK
3jNH2qpfzy1Ky5+vMbja5XqR+QNpJr2jWOd32qQ6nWzc6PnBXIS6DbPFqAFlxhTnUNsz7qM+ouY5
yYc8lss4SYgZD4VSAywlXwow23P7hcH+6FZ/uyqV/silviel4nT0TLOFocncGS2WX9ZOHvanV7bf
7gaodQ/Ciel7HQPpzz569+4fex3kyl3TP+f6WDPiN5yJS8jN166uMfQ+k1E5aWDiSDkgdIzpgaAS
hyCwIC70Wubi2/gtqDgNzB8ZCrcJMNdrE2H0MUpMvtYcLWtNLG9qLyLwqbWCbQhuObwsGJXB8674
nWwfkpABjK7YMkoeXAB9+1Jcz1UuLH5JiHYalYVpiAs+pRjppnX+J5Dn2D68wzWXw8DsY9t5LI2t
n2RhP7ipr56Rmp59Ej9Mj9el+gxXJGDnUqL2l7lelDDIJ46xj88VW1uD1RmN8mpVJgNhKroV+3t7
3tbs7Upw/v08rY0C8aH+idAbwFoAoKHgUvTgQHEdUbrnRAX+Z+XC7uVCOXC/cXiRgkcb0q5RG4YH
DhbnzoEC2Z652z2e92gHrtx3Oi0w0NHUFqf6TtU5ZTsmMP6cG1JtafcOsmbdG3y34UNxDl8FStSV
CY4ellkmxBnkfb/8vXRxzrKiPN33UP4NDKiqYlA0BBeQDXx6E24n09QC1QUaul+xuqvXUSf+SLnP
1ziAux4N+801a4B6LVI73uHJqlGHpx93QKFh9RLxS4rM/piePWDHiQo/dLeIXT+tAixekwUKXXxV
AIagt2Z4JarEwBKrWN2lwvVsmhLwmNqbv0i2PYd7JlnRq7vJ4mqER0KIN4NtAeiTPi0tn5+QEB8m
UIFghY4aAqt6mBPDWdVjyFKhBMbMDhMF/F/YcTp5k7TfFKh8UwsED+jnSk92+3lsJwvUUeU4jBK1
diwDNTzt3JbBoQ2qLe2BIa6z5An2t7U7Aa5Nk5LXfJuHdDKBWxSXYxkMhk9qnm/WRihGsfTCkNQH
tR59hz9Ssp7iwCXDq2OJs2PcX6XIX1RDpDLuxMcuPC9FthbakFGK9Hs9+CvX1vuBvpwjBrkNaHvx
jVpdjindfUTvRMJCAO2KXQ+YetR7k1OnBU3WPQuM/HnB9+Aerq1u5yW6YFliQMbwlS3UniwLa+2m
8/A5yGNXcuhwQjV7wibC3+jGfgS1jJge+zjlkvkdUrJGVHbh+ofvdNLGCgEQHmT3vRTWoto5dREa
8vkDneb5y3Snhbr2bDAWUPz+dJM+Pb8qp9wmnbHg9SHU9ppKqnFXMShTuRlFbQxQb9H37X0YUlke
Xqobw3gPIGhsTlFv0lgd2i8ZsTCLYIAHmWsy5PBIiiUqr7h0z2AXe7Dp0L/ByxQdkRgrefib3GNx
Nco9PuhX/biadJDD2Wqtnnddk2kIuOt79pW1+YlSeMVqJVG+hFY2b+aeIs7FkMKqvEZVQ46hlQ3S
0uN4DS5Rof348Ebl+Hn6PRT/YD2ehRmo/u67ETxBvVmzlh3Oe6cSiviWdmxHmIG+BFDznMzl1+Ho
upXLqlAk6gCXXlq98l0TREjI3iMW1y/J3NSQgxCiYJ2M/CLz9lylCgG3IhzslU7LBTcsU1c4riXc
rFLLJd5Wy2AaFdhRgP6nProsjYjV0cLM5iIRM955mGARWZl/ia+XrXRXNXa+BN/kxVH+4zXLLLPZ
mPURmLOZ2MSWL3N/Fmg61Re1OutONlx5DcObAxWUWiKCtZTWSiBLj1aq+C33WJsLykJ1Zklllh46
DJO65laIn5fzXrh0yh2XDSOWj0pok25WPi0IeXnnBjPbaLLR7ZXDJCzaQLCgC1Qrr7Y9Jh/196H9
l7IThVFi7P3bKtS67lUSWCLuuVtgEpR3trFCEr5Lc3VPSU08Ju3iueQFugnIQg72spn1u1r3M6Pm
Pl6YXq8ivI48NaoKKhEybQl/ZZLrSeO3X9ut+KDEHPxfFdsb0fUeu+lVmzE0wfuQPNz9QNOiCU7f
c64Lp11gdGml7o7qSQuBZZu+Q1f+I54y0fgLpqhnf7ccM4MPux2U8gDzgaSjDdyBRF+CtC01Skgu
2faU/bmIC3OgQF59qEL1q87ZijEIfBE/TW8qinj8vLIVWtEJtS1TVxLxjOpkam5AQZeHGjFWMxaR
UJQ1pIv6fSbmsg2eLgd2laUUdpMGgcx3VEpkSZuAAEvB+NOTK4Tqp6l+ZZwqXg+WWcofuwwezw/y
iSJOKzm4XMDBvERxKDWDCeEK7pa3KdW2+M4COaWWJ78H5bLwz5gFlMS+UrISlDzlyJQdELZ2ZmP3
4eGI7kf4pEX8Pgji+nPrXmBHhT3T2iZHwtoVR1bC89rQ20TLpsUHS4dF8W+2nAlZgjOAltdlgUmB
FUguFUsUUR4Jz2+LGSpYzPqHaX9LkErAmJxM3aZRG62FSQiFBdzq/vNSHUa0wso2hmdTirDg4yu2
wj6VfKWHhCNpmGEGkXKEBre/TB/IUTq46z54l3JWJhgp+V4BVYkaUsFJKlmBST5i58/W7J+icSCF
nauVNxXdfEUf6m+Dwr69zObW2GSpOtGLvGIHmPRLZ56OCBVn4YK3Fodg1knnuwFclXqW21ZDoJ+N
gvdxTpjRh2xu88DvBWwU6fCnDRxeE7Jb9cVll2rnZRXKwnv4yvaV5/HUOKCQJvbqtyZM0oZ7Oi5E
w8fR6VYbUA3kXZ8yICvXPHCrcCyEvv/U7PLe4dmFW1bylLIgSuRSBkyLeUN8TP8rtDSRKX83Tufu
J20JUKxs4x5rzXbKKD4eKW/ohpu2RdG9+UynrbxMxFpXPT6+ik308GchkRyLt80ee3Rnvu4/zVXe
NISeBHQbPd6ZHHn1AdA9cqJJHLiQPIiQzdLqr1hDn/v3hCFe8a+oqvW1yhOW1DW+i5PUKLJ1FD9Z
YaO1Gjz4r18a6RdCgiYps4JVpkruo7nqwZyL7J4Wh2uG34ItlOncmalmARK4X/Q33lmDN61BZ7qe
uOiKon7yUVKwdaBL+FNnahQ134x2t2e6m8+3kL2ewHAxcgAj6CJ6moTwxUoJygoPcxXZikBmGO5V
Zn9MXf6YovPhqUrmbjvxDbPGq+RyncOEe7d5jCA8IW4W5Er+94KJltHFDX4ift44orO7ZtHR7XWT
f6NlEwIwxBdUqkjhrdg3U0H9haQfJUiw/TVAf+3+x80yYbFQFg6H8DXGC7XQPGd1KwHaEE0Jzi7V
+06HSH2I6eqWIcMC2z1wa6KZ3sUo+bZz/HD+SImT1tjVRkT2qRhLd84ld0w/tR5VYkyIjebIRtkM
oicjCw6SHRb9GrafSwdUYslZ3sFh66ur48AiJVl4qQlz6YLAf3sdT6t7GHwGwvdvC6Y4+3/Edc1Z
fz2367kp1TOnDRMeZIvMZQ3meeM7HvZRdsRthztn1uFY02zsa5wgSoRw9V3P7YsEGRzMOBnjATQs
II0uDWmiw7G5F68SE/VhUHcMwHH/C75VDhZHyyJXnU96jVDSCrxTqW6j07t1Uc0JaGOCZ4SZKXTp
FAubVOOFUVsEJcitz38hPv5iXR2Tmebluxajx7MyEAR5rOUjwRvELDD3L8Ng96PAqFVcX0UoLFIt
Y6fJbbjRAS8E/hOjwlvUlzsblCLek3au5NzBEyXETTpbyYXMKoGy9h0obX+vwfkukz/wIUIjFpuQ
1+4HP4VEof5E/rNx8e8/0+gem6niWeIqoomRk5bm3XILBeWZY9j8i+LQuAueA0Lko+bPyZLdGGw4
/WDyJZmp8xPCFYdZFhkWy/SmnHhb31EwwitqEQc9GCqIGlzM0hvLZJ/uXnKSSFJCa0+aTddT50qe
m0IkpBzS5Lsg6fWJiyeRTksTvVtEup/rTyB9QmbxyV8ptFS0JdBxxEUWBSBV63cqXmLiyoMYnkoj
zBt5EqA2xC8Qzuqb71jfMvuY2VX39Zsh9BNta5islwtxgk1aDXctovRHlm842Ek9YxPP4ymZW5x4
9dERuQREJv28ZGlBcWctsOQHLXD3xZ7kkDZ9paKF4B43fPtDEOQnmkMadDteLiSWCBfyCTwv8Qyp
m2gCyuVCyrIUqIrvTSMhzuRu386puUVo/nQgFBuW9FObN/zmDYVJT8NIpv+Ynu5ckSHwazfOjJNr
P9Qk4vr+9S6TlMlFamun8SNm3nmDlfX2deg7MBFvJpYqY5QAGrvb4AhRkUTcfCNscSZCcT8Z3R2h
zIcxx+YGyERASjf62Mq5e49y9N7iFzpmglcqyCGpR4osoR9Z7zB7h4WbkMjxMs3Bzw+6ys17lpm5
/QXlaYftv/FJO3OiEFHzIp78NodDccfDTI41/i5+md5BKDSNKUZ+TrAC4eGane23wiIHxdB1F2Bc
JQp9HiPVYoOs/gw8TxJoLYFU2ZwQSv5tC/1tWFTH1QVSV6OWZ+lCLHl9m25sdOD3qdCoHGSnX/Q9
GLSwxmXgpXQMVcO3RktSIgwkbFjJHnic+ISK9qtok5aoy8r5N1cMkF2xafvuQYSQ3+DITJabU4Hx
/w6aZ7cCmXd27y+xBOWKTB8wJOtSgwBMA7Jk+r1qm0Ek+7dnqLveojFrxswWOvb6XamPA3BfEG2s
9bO8FVZ3Yx4ppCiOVNL8PsDwmUPHyH9T9IM850HV5AvM9CYRmOK0c6KoiOWD5MaeTKofkxKj7V52
mxWmeh2rfeSGN+brYIL7e1cE+FFg0R1Xtata3XzPM753gHSDiCI+WxbTdNRGwxC9ys6dVK+BM/xK
tkpl/P5inVr8Fol6nhYjLMqMNIXfeundzzvPlsyr4wc4Z0OwVCCGQwzeX47P3jE++M440LsM9+Fh
dZtw43+alqRreDoWnWu/Y8XBskO9xELF7cttSwsAEet1gQgGLUDZR0TgJ9CUS75NkDNSkWqU7L4r
GqxqMl05V5/BOhPkBkZCeSDtnZ+PJgOmkzRhT+W/54BGbW717GzIcZJgbmP8WJot9Lkppz6CcAU/
6oBuxfmBghKa9hf0W7TemUdoGXRlGBhieJKPj4KEAQFlM9mJBjWVa7wW5RDGYCaMPwUEyHV41OFl
ZRH+c5soQVvEhlJDtYvUa2lOEMnoFIzPCplZRGw5/WXzLz91kUvy6Z8f9GKsssEPDHpCe71Q6DoB
du6tgVfpwiLASZtXUlvdic8R1lZVGbaLu+jufi+TrpsUeWvCrU+GvtcQBtA97aMLwo3VjRIaqakC
ZltmBJ5KfNkupNvEPDwJdUkFoZTssgKY3IaZhK6CG1oHPUbq+5aGnAPvtYDYrxNyk18X6vTbLKxT
+Rrz0zXPibxHSk5ACFnOq/XBystITblUk62QTEjGm5tAA821WgzJZXZse56R8o+4mtaG859XnMfq
bK7KXXEAS1USdvanwXf+bLAW1AXaLjp6d9IQ3vbsTdSLFdOfUJEMlcE4yF4IJ1HNhtjGt4gZ665P
YJjHJcnDrN6yP3D7J+ZJ2tfiyxz/XB14Y0hf4FmVmNchAeIVI1wjQPuRBu0aWsRVWNKNTA/eum58
80diJX4BTcBFJi8ug/MEcKMdWhI3uqyeENp2HBSTwvisSXg0PJdV8gkdwM38ay0oHPH1kQYyhAUa
oIEySOXuHr4YZuQnYDg9tLBf5yv4nW3lUGLSro3dds0vyFwQqhFQs9clPESNwJMpgWyiA2X7oPWH
FiZjCFnbXW1B6T3ajNq6GjxEIcy1KOoCLh1WdHQWGLiK34yBbjBBU0hgilWv3L/sYLPnRq6tjcP+
60yKWDziccKXwapsHHMtotoLY/N6tMd42g4hSuhtVY2GELFWcc/WjfNjLCe5cyW/QMA52wMbrkjz
GBZ5E21o0gkrzLePPm00rm/a+tVN6/3v8F/rL1NVDxyUF/gXocJ5ou44Vs0Sjg3CRHUh90IW0EBT
xSPhFu45mPXQNa02YRcVIkkPPOqxeidPcsBxoI7eQfdjvg4RgnLj9USMq8+leRL/sLSAUF9Ac91Q
1edtfC3Jq9TNbAbA4l8r7YKsUpY8/xu6rRC4pUFj+s5yqYvCfg4XaOmH9X0XtPQu/+64Z355HoW5
Z9mH/XZkRCIVsipapRaNMGgxvD2jz4CKMXo2A7/rrajYjWwgKNzQIyOU3hvIVga0lu7JjsOIATSi
BqPuuU0sKkYSg01iJA7T2km7MdekEgspDAFIykryecbp2YfrVbLMhUjDe38Glbsanh49er1kwunA
0M3W3hVE3oqRHXH/wbEBjdoMaCO58KxNr2I+EBzQEJjb3PlK9ExplIGgFAjEHKKvjM8AYhWMlKOK
2uxAysm8N+NM22/9ElFGP1OJMUu7/S8gcTubZ3oGKjU56oA8HAFjPHqYHazJEicUVGOHI5RALqs0
oty0JMnIUqQ1ZDxFqPt0TT7OCY1Me9EAZReRKoX4W1ZYGbQinEjyQXzrT31fei/kg0HOAv7P/sif
OkZMP8/TIAjPpGMD5vNBpxlDJUxTg1vWPnKRfJzjBR7UM2sMVgbCdfm7Y+4ZJwQ2eE1H3WbrxmKX
rg6wg4JsyckEGtlRb6DrrblnLw65EYhT8SeEBtSlLlWOkTz5ml4x8fo+cxcjDlN0L9hf/+SBq5dt
UqozV10G3BteGnU7SDOSwFInt+82zR4/41mXlKjAV2Hoyq1+IKVZYyDcjd1uYrgIJbvFlp+Zu1bU
ODDiU6zgs0JcvA7wjYsQBnk+ePkrIms+V7HkS7KjP2ZKWPO0bCtDuU5a3Z9hk5aYauS2Krgsgc/N
1H9VKv8HgZmMSP/uil1MRpsN1INukYPEZQXJhBq+D9FyXMaj3+eHfrxjqfLyMMFW5fbJTOOmw9qc
mVptIBkNrviN3RdMvVgv2e7NRuQGrcHjFk9CiUTGIAdIzaxu3WpGvJjnwtwxChBp9UOAgfCyd79/
DSTjYms/zg92U18CG/TG+RVNE2G9JgH/KHfolPJd+hDuXiyfTDSAWRmv1fPen1AifxOkxox1PvgM
N+11sdvU+D/l4LabZ7Neqe+P0F6fMT5HMA3T8OB/jJ3++jhf7YyGgM2WI1+z0Cjv3PertVC0Hwek
yuG9EnWlOxnCdGdGMjgV4E4mkMGpfWBODU+e4Fx9W8+THmFBD7WB55LSJZOwsYttyVtpFnR3s3z5
lhLgZx2RIUEw4fywidFM7WAiv4T2PoJRwWahvZgAiiHvkn+tXH42LHkRehUlJWPTsyll3LsQgIT/
91rW8p+l5Q9jXZy7KFKYXq4AHIWLfa12JGVCUIWDJp3sjC5jLnFvk8q9HFBPaVLmCkWpvRcQ6k42
EFHKu4QTjDv5QRggrFx75Ut6Z2oCn24HwOonY46vVXRSQZUh/QOfbg7I07srqbX1gzHLTrgCp74l
SbDXFd0CbNthdM0cYWwWxFYES8LuaJncVaRdmA5+e+u70WtJskJUkUeCw+8Y5VW0aMmVPTaYEn2w
on0Lq/AYLGF666kzNHIfarzCumCWuJbZ0vHrPDK3ZhU9FFSesikFrI+QBA0HslvmatUHQ8XQygUz
9Y2dBzNW4LFBIsBTMawjG/TSbZLuQXil6rS9OnJVTSeRgn3MAohu0OzVcy00X7OwvDwcNOeniv0B
a/Usdprbplyd5B1FrPGF6gpXLYK8Mp4HhW+OxbCCFrm+8kl+A6XqjbqyX/U8fNAcWleWS3zEQCrU
+da32qUd+8CBzQUXoZmWK9qDj5T3N6demu9h0g6OZU+o4n0SVmq12AwVKL9KsbRtkWxIq+zbDSoZ
u9JglpQj+uIS2SPy8OMY733bvgj7Sby2h0awZ2s9sekk64cXLEnCzgR7Kli6JDN6xXbfINwW4hxG
0IEpoDMHwl4f2rBcWvxBVk4+TBNn9uwyuwCmyJyIxlHg2XzOMYCqA0KlKNLrPvjfuv6Qwq8PsGwn
Y0x/6otCnv1O0m5qnWLaBY0BRwCFH/ted5lWgo2/3ZOpja8qHlG3/mR7VIV1fOwtkFeKdQQ0hWlN
AWtDKCIXk10odmOGVqeFafoDly/E8DO0oRbM4gc5dr5pdBITPJAkPwr66ZK9eQW8mGqvsq9ALrEt
3bb5+nuBws0c8d08KlObjwRcnryVeKKV1yU9FLlCqxu2w6So0GYOiCqMxiPc56du+BZ/N7/OpeU3
PXj3KOyoKfp2Bprfg/0jrPZLt/cAPRXvRgIugkBKTEZJ2pNLeGVdUG0GqgwUK7Kp8VLglcOVOzvV
cBbeUDhpyFnX+ma26F0+bsNn271h4Tf+Uk4SyPCRm9psNSlfmHt2khz+N6KDy50KRjzfxAFcTFCT
4PBo/usHB8RJP93m6H3qSM0LiB8HNloKH2dGuTRDRKCt76A3OnLlnepRc0eab/5x3E95BtU+l/2n
wsnrcbqXK2ADp+ibqp8eHd2xQzoBhA/tV78vaAqUhL2J8b2TjL77uE7r4Ro4ECtdzk800NQK9CRb
BxW7ydNDmMDUaUQPsC3oxlu/JxvKPRx9isgBPNC32pklhTgXR7TFV+b+ipxg7duBnvZFmYEibOAq
A86fczDc6FHYBjMxPGxLrKw0krssL3k3Jeys4GC2St7QoqBI5BUP6PBga3cCURCuHohXlPmYxEGP
nyhrWrAOD5yU2KQvN4apxC0sAAZ58kHn5+Lzn6kxuSRQtgxWn8IvkhD+cq3z3359/SgYagg4vxmN
IV9WmhLp1TdqMETcncPgrTmDm2y/4aFJ1qSE2KOEfeIqXlAGjac0qbC9OgKka2ge3s57zR/Dm8AI
R0jqEdYiZvdMKRhrvZBVUEjS5pL7Ce0EZpc1YPUmLJz6nO99p8mY2yKsTEoCZWkkMFtqvHYrWLrQ
zEzZsxVVqs4WcM94oFPzlwdAo5bziLxsjvUOYhpsip8vJ1vLQ15BYil/w15DPRZ0md+i+qPoX/rz
ugq2ColaMCKjZzPD/lHR5jVbEvUA8DsPxTBJ/LQTq16z+p/T524IYobNJoqYzSe06A6wshckZeUL
I6Ofopi5rfcwIyw6z17pchROdtLey8ZJA9fK204ESpDirMnaBdBkxYq8Vx9mbFhBbBQrNF3478aU
SqPkm9Z/Gi0l1OXyUiaSl2FLpM8pJFHuqKLDVoo4Wd/0juBCnyieifKEKyvnsb2vxDb17czLutbE
+94RBmsXIqjI2CWW9PbCEfugFpIHuvTbu8IyD+ZTjivnWaGn+3F3GR7V2H/iSfNkZK+SqbDVTj2l
6R9V4a4NQJb6M9xlheRqMu2KXdT7KdGSfMFE03jZgDnw83wS7YDcmONAyj9BpJ1aEWB3UX/B5Tmu
fI9NkKaOpdlM/iLmkn3XWg5q2fN4ITBskIIxLLllwsApEfd3zRW5vOERhtbqp4HW8wHIEShteVH8
tr7qWv0jjmkVHnvPYhlk7JxAgeq+RZuxI/t1/S2DvKHjN/byrdliCm3CMFF00nvorHoDEEwr/x94
m81uOZzVx0Rw3qQcPRsL3gUcMRT7IrjHr/+Nb3SO3r4e0h5uAhvEmn0PcZJXiSSgSWquoJFTbVAC
tNtps04erxedBH5V1y/ZyGmIwsuF29Rp6w54ENuyb1dZb8IguUtdtzU8qSXZ2kyXCE9aBeD5tGba
8u3I104P0Ez9ZDeuBKTbGLHii1EiLKOp4kqSccnv0vYEJGk8gSjt3CwyETXliKwA8JOH8UBkYesr
CTG0/iEhOhUNsRPSSvKCsF4066E6cDmgIwlgwnXB02j2gJYaNAiMDPnc46qTmJa4q2ENjCrf1v/R
aU0hhU6XWC/d2SaI65rI1B5nZQQcvjFbmsaWRwRLGrQaZFtKoZvtlxZVXz2PwEPO9gKrh+2+FgXY
mWzTEGymnXwYbhajwvvEz4o94tfTVbvDs9FolE87iiasRCDy4vhRvjWKLSkCS2t/KoJtVSxie/H/
jbeTK+JHnFG34pfYCDtTWlpCp1pe6nQZW55OSN6dC0Mi1Dj/MEJbEFm0Jnn6EqTpFM+JLJraX+6N
7U+cliscK3/2vAOizV5n+04O+zN07ZWRnVSJ9VShDyt7hvY8nCjwJvXIJyKsZHbsERknaN048WPz
+juXBzL+dGwZxJjS8nT94H7uPyHmP/pZ6CUlxVa7NxI6qm3R1cdp4h5DmqAXlIofq2CBuL2rhcac
ZZqlJVMfKdHE7rGvF9hduRvEkZK8nJO5DFNhDcTZoTuEnwHA9o6Y6mS+P1/CEM/iMroe2KLpCMiQ
BlXF2k2LrVicK/2I4cFhZbhBlpq1Pj5ziTkfOwGvFkiV+JAm3CTSnMj4BCH/4Uq6LEXxGrA9PmQj
+OCeTM7kD5fL+MEPe3rPf1piw4PpI2vXM/Tz0i9nslVgx5agXA9w0GAdVYG+RV+3sxxq58cdn2vI
yFv2+P3+TKe+pzh9wpgMzY4pBTamOuxTUtwcYLIijoYnVvzkpb26cs6bXU5mHg5IaxGKhVkBcuJ/
D9s0d1JZvQlJIna7zpzPgRMjMKFzvuJ26/LopDBx69W6nBkY0gbTAzrH7UO/HmycAxbxgGrLdyFv
ZhWSWv2ZOZqu4Hf3kTY7QwZ3n9tKFDGpKrZomTJDO3ZTQ1OX+yijdt1Xl0BT8EuAIGDidcO4qb9d
QM+ScoR5pX51jK42FcKGAfB1CjfVNJ8ZVYAciT5R6wCr1fWfxPmLhWFMBIPMHwCwJr+lQDoLXwBT
Y9zPZw/HWTaze1+G2q88zMHDimZIibUZ2AS1SjxvPbUMXv1F1DfcVT98zEmiT3OYbfhe9AezVaRC
JII+HQcKiRVojSI97VKc0X3ZxstFQS+eWS0lG/UoyvJGDtEAbOCN5s7MP0wQVBYzJk/DfTQRiWKS
TKNzdM/Tz0XcjAAsN58Yx+FG4AohLa+FNV0Jvgqck25GUkKI8UQWawAcGJvsuo5LHNRSSacCDuw5
6WjqJs8Nqc7BsDZiXY5EO02ucKIgZhyeLd08cymM4kqE0A+AbKJd2rf2X9JkvU9v1KcochM4iKVx
F3EMiRrYG8t0lZiBVy06WIhnEhqSGe25x3z8AzKo158EPa+NWy3FQ4Vk+SsZkVRqqTVzJr7Paq6J
VQIeXOtuvRf/jjfMsdZnso1xvuO6xbmIHZzgznRJzQItP9dQV9EODOt73oJvU8xk3UOcJqtMdJG7
S7SG2rvE6jxwEr6eDlQjejaDp1w7Qx5KSj1kC1BcJ841YL6pn3djD5m5fL34t2T9rTJyoSDREEWE
WA9Fy9HWSrRAm9cIbBeZYdQ6c4kIGbV0fGLV5u50UH1TEjkv5s5i5vBPj3GtrrfqXQxe8dYhMdiX
hx7PGA/GAOjp2XepsYyi59r6EI5JEuZOz2KRoZJadq3fuP4EGlrCRMsnV5s8luqT6nhbfqWj1EXt
j8EGWwVflTJEnjW2qgYASnR0FQrloElvd323AinaFKE/gK3i/9qKn6x1W7IdUDeyKAWTNP0kpFuh
3bF0y5hATgfmjfgMI2tJLXO4fhGy9tvjlxD4cnfTp7eWsfX9BApdb+2Vgv6bf9ihDM837pqyc7ir
bUlCKIs3djnq9RoddWXtedVRlU6PGW7ykh1N4NmBBei9sVv4fgFUn0QIRFk9hgxgkkZT9tYb0aJI
Cv9N7Ep2JWmvFIq0YMJewj6m9z/Y2lIf3kHkq34LTFUUZIKgFd00YSn//ZXdSqzze3ROvEVsD6dM
ad4x6Y6SkND7/zxJpF40KHF1viUGE28HXATFtZZFti9+WMrVSgJF5M3CjHVeu2I8lnLvPMVUAzle
/piTTmvek0Bvad+oDADQbw3szPVThsm9b+vSvUckx/iukvqXTHKHrNfrsUlplYmSnpELf8CfuDH4
sqphqtKrt8gkOxbWCly66nW9NjHUAOW+EskeGPkFgbtSoJ68v7pZ5ulDLPd6NYrPR9vK9YKXv8Uz
hEh63hPRxp0QSHG68pT+LjhO1ddg3zokLCgw5i2piQIAjIKq/aUVL6T1EbsLowXKd/t+xsscJW23
utmGLQe6a5JsTiG7+8kXVVm2ZRXKhm9BtAAjNYkSFJ8lNGW1xbcmX/LZtuGVbk+gK6nLnsOUNQx2
6DJ28Ux48R9QbeaIuxLdFYcUaENfOhpndk1+k6Ibz4L/bUkDHEvhEzFk0dk+iVKrFFMmE2JEyRcV
hJKr3Qj/VxkLkEYEatCiGpy2QG9ggIeckhBd13cbeIul8FmT1oqfJMXvaXndc1dhIED7Pum5ohvD
4giwfS1QAAMC7mnwEtFzIZ7UcsRLuDYtLkZJirJBzcq+2qcLFuj0AdbjmnnYhq/t2REUDm8ArXf/
C1lb4J4i5bupAwD5BeO4eeEW6+OdiY4VJOMU6GqZE0w24klFt/aHWT4IrJwgVrG0W/WS6TLuOneI
sPyd6qc4OlVFViXDxm4OrVM/2+hRFOQVn75JaoT+wBfcICP00kEUe4JEPymx/blyGrqm2w+3RK28
Vz4ncRrVgC3mMxUEr3K1Wxd4+iCj1dBjPc+3NxgdoYtXei0gyQvkXbiOAKiZVj6mAg1maHdBv61Z
TO0QugwsmLuJWD/AoLdC75QEhKl4QuIfwlQd8T1sBgYKiMU0doRI35fr0tER65EVpmnmk4aNYPpT
MvnzO2uNkIb8bmx4zb8bdATpb0syD09lAXRTZKzdLnyKf9XjMnKzMPBXmDoKzolZPn44bzSouF2n
7uv+eKQ4MZGM3PVvph/esfn6EK2ROrD6sZPZcjkyc4HEtdmSjIPcRek+WkVwNsA6iBxTglLGe8vl
cTVcFq1xxRh4pr/DujjDRkPrQdQBzZIgbxcz3yFY+sgcpdYYRHWHNuz2au+jA8fZnGM6kbDyyD82
0/PRM17LgCCc1w1IT/yMD1vHMsZoX5KpeOsyvnxsRYtozPYurF7jLowJyMijmSR7qZhVqUaKV6bv
dKSOtKVxACTNdWNQw969lonazefnVVkrK2kd1p3v7llqO/etaUAagKGgwp6rZfJXhpfPCsBzubuj
+FZOetOwHn3Gdnssc1I/UNDUbG7lyPgqIKjYFoB7lf9IFIpfhvuqI7JxZJJW0jRegsFjSlGPrV8c
FqSV/0GoW1Vs/HtIZDUyCdSoCsiZ2hLHaaK2KVzTgHm0YmbBbgMzsg541L0lsUsll/3IIex/FXBT
LouBdWy59z4WyTR3XL6LXEJUHvpzgovWG2jnnSTYNwaLKHxBwz8g++nsoD9dyf3nj+Gliq5tMI3Y
rfDvvb9J3gwUL7UJavN//wJ7pYhBTa4wG019wjmx+Zc7Wkzq5hfaYypxYWdqlo+DbSxrGKkCyBKT
6GmJTkPo2XKh+MWck5K4+ORSmXXbBQeLW3YgKbmaKRqCuOk9K+vpbt9ao926nP/8kVtxMF9fUhq+
w9z415m4YuKgz4VPxW0WBKFuHjnMM+xDAgfIXh9LpmvYFWFXzplx+NhPuqBM0MRqY+M6upb7+wqv
1xH9VHSewqLAfMHnn6COGy1efnMWI77W5cpCON5N3JlLmUmPg8AL7ABKCvXhqhBKlkT6q57eD5aD
CFeuzkdykly0/7UhD4l4i5OhfKolVPPZAMBApcQ/9/zoFeZY19GwEVnROM8t2rTgC6G1TJJAMujG
/3LC86OlfyR4QgCdMaeW3ZerAnFXMoSZhWFSkDBnnluSEmEqEqwVc1MZnu5RpkY/MM3RmclRh7Kk
2S7H0ygxMRg/D2h8YwdEgbcbWwZNT956xaKrE/J1ESYK2YKVUiGPevgnqRFkXNGmVUZbqGUcWta6
C2Ec5tEB3pYOTZ0K/9XKXIx09+wy87Jl5Li6ofTlbQV4lpsKFMSq++fApKZK4Bmuq9JT7Dv581Tg
FfjicBbg1uibi9PMEaW4bSje0pzwPTaVPJO+RXF+8pwCEOYE2OOC3LyvD9rfDHcU2M2oIxyK/yxV
cYngSe+a285jw5FMiJ7m0FRao9eiQN+pY9CLhCQH7qDb/+rKynSBdhgCkCSLPK/WejVD2hCCNrKW
xaldg5da46y64GqMhCHo7yPaznndG45+woM4LHOoBRYpxLOK9z6XWzysC+OJd7/IdFCJLYanKn7C
l0X0UHVA6zEGNetekB3o9J1yovmhqj4xx8J8hiEgJBycC9AAyYVRO+BZiBBbZH9JNBK4QSJpAPmI
vKUWicJ4MubGifpRGrtwv7hNSqn2TeOhRE+c/sY941nVuIzQz9qUPsTDYqqWwUoNaE5ADAM3aeNC
4NB+Dl/Xlac5bvNLPToh2lVCp/CrdXyn5LVr7KRr4nEb32kXGJYuHvvurF2dxq0NxV4QJ0y2eQIp
TdF2nJx+/JpFd7OrlBKn5iDHQYPXimbyrXrkofLAJR3OhbAfO4bV7lwJz+l8rgp+/woCBCbfQ1EF
jIY4v+wKCtY9gX97/+jAS+llbJY4TLd77GugjJoH1mFsgoMWKbLsn30tWRx4RkADL3P/zpqOUVs8
HhM6FqZU11uC86/KxvzhdMoCXootrYWgOrSDUZ+eMytpYamcZmiDDT15rYoVv/yEyKvRSlv2kQEz
yltd6pMpz4HMn3wNcclRpZNxJasYAToWhRZ21Wf07vp9VERmW5lZ1nTW7TXNFctc3z4wqEWM9MiN
RI6rDLZyZmjG6QsJSDibVUjkbuijdfje63YA5fwHN6+vz7chVrqOkwSLD2JDUz0InYrFQy7QfKmZ
IgNrO2R4rZFJl9TlU+0fxqZpQ0uniuAU7l9/Kk9cIxyLRkELGT2tR8SsLOLkJ11K4gJfTN5HcXbk
sBsomnJfj03orb6gA3m0uZTXXo8KoyxKG2gQX7GmwtVwPBfjQ4A+Vu2tPR8Tvpg1hx+GS4nHZae/
OON1aXh0H5eOvGoOQT71xZ30WNr18Kp6dfTRKqHJnbsf+tdEGkvjA35BxFclwkjQ4fpq27nE+BW2
ve6MwTu0apldnfxQ4P2WP+ao8B1ByoyMmImh8Z2/bFiDFFNt/bCuE7MPuFGfF36tENQ6gj2CDLw9
ksv+JGiC5JZ6Xhg/RI5YKmX6UPlq18hwT2K/HvJRRXjQNHEdB8PHitbROQO3jBWbLBuhyPXYcyQH
5SNE1HcYCcrgk5SkWwN7TXiMjsjDEs9J3/h2hMhEnRydVNFbRO1ltgQYb6BdJoG8pMF+eG/a43FT
+JXnLwWvpIIz25fwGKDFlgXTXOc9Oi78v6z3V4928m1lYgtJDYqEU06QxiNab/PzWdmBhI/38UU4
ZyOF0YDwOzJ+GrgJFIc4SqUiu/5zowJ+KzklnBLRd+6VmvCYV2rhZEFs3mIvb+38Ulv0y8xNhaVW
QMdABoeQLPdUxl4S3nzFEbgdWd0y5YQujDgX/VAF0kkoYrTBQPssxjLC31xyEFl1rTpPcytBSZBE
lDhDZQmG5R2c4zqVIyLZT1b3QUYD8mCeQ9MoN7nY4P3x26xFLpPdTsNWSCEyujf8ak5wOwP7+1VU
3rz/Veyoigbt5d1j+faGWZMwbgO9n/LR/ZHCFlHCaXVKLxeLR+P/VEyPXa1OcbpZUjpakfBmor4M
+4sOLUao/wy/k5T4aFEW3d5mhCGT9H/hlbs96ErmFQfFlU74V6KjEjlcWtapdCQIFyoVu9l9otjO
Uga/Rgalv9Z8pTThi6nwuBRKBY2X+z8GGIWvgsEEg4RZ1CLFMkjARbbjrpcuxcBlM5xOhzDNc+8Y
1g3l3N2wOwRb5Yigj6NDKjZnB94suAzK5ECu7Q5P4/wMndET00UB/Bw/tUL8pLMxytgbWZL1D8Rh
cUfQhElLmu+cYRzlEoNWiq7Z2oyUT+J8lPrx/HIdUIqxwU5s7itbc+edPbW95Mb+JzUQWyEd1Cn8
p/gHClb7BG7pIWKkjpieToC4pYZ0+158oV5U3ZmxRJVxiz+001xo5VhW5jtckRoLAe2dMyRbdBVp
LnmIiymkn3GHETOY1T0/OEBgyfNUchpAGcyh265MFg2uAAcTD3hC/OlxTSHlyxoNGETzzQXJiL6b
3klIkKV78F5dZX0z8Zr/bVSDg4udUepufR4OHHYt+XXUfjJu7CCARBfnnyfTWJcMvPNXoeNUV3G1
/st4el+4wl8HshWJ/JeYmLA/IjyhmQ264K9zjjZT9WV5eVxSOEkLALA7CUoYOsoeyYyK/dbSuf+j
i13hrW2ye1A40CbsY1TQOp5gPLZRcV5r85JGY58bQUAeqXwmv4VAbx8Op12KZXpwiXWb7e33bliy
xw1z5X91qIi1bN7DSzyjH4qfp5+7EBY10todDVjs0vRSKTwXyChHutHRFWaxqjtLlySY4Lm34El5
NJzYMbdiG2ol/U+/jJnorglBDDRdWSmb4TDo0NN2WKAgnvPlVJTf/CfY6+5P6LKf21DyT4SY20W+
rIBlL2TWQo18yqcdkvZUPSRKuaj18MDnzS3JHFzHte4V3JJrFTscbQVaQcHubG4oNRqVilPeQkZe
KADEXPFS7ucRqWtsCawkonFkwujgJfwXHJ31gqzta2l9csJnNIhdNUH+X5PUOFjdEzuYuKzN1wyn
WsXBSzkcKbGSFmXusstK0/kP//xtqPExZsuwvk3mxWqJzN4KJjtghOPmlvP32CGoLfqKfS4T9zZC
/ObbV3cJtT9h1bSC3/+O2OFXwh5qZ6i+fXJ9+CufCKJ2U/IdffuRGzkxhmUBp+WB4rVuZbXSufGf
KrTE158pql0mAMloKzTwkqDFVmLe440/ip8SH67FEjzQlRNAHM31lVcLdbQojBpp5mVlJkbrnRsQ
gOYYRrwPxuaaCjGJmMwPMKi7j82o59ANHc/F9GCIqD36BssAtWM+FqIWKPwsbNSKjP2691JJy4ct
86ntn8yb6nw3BmXgirgCxpB/kiqsCCIBytcJB0tWGXhVQuzOII5+8g0wCpyZVk/2X26E+0pyMgzI
EEBTk0ghcndW7GCgVwq+OPXPKyqs/LhSsQVGomss/lz/uBOsMC8K71sVCidfTcod8p0gawO0hprO
aOk7g0TZZ9HEu6MhXuoFDZNd+Vwt8Nd+4xCiFKTEkf6rE5h0sRVYla5ylHWKCit8syfqNxXJmxB0
uodVpVPMDCKvtZQSGy5FiweXmJrP7wcaAPmeQ2Ri6E7VNw7lnavPiZwp9kFJomHpk8Mfz8TlbTDn
YzTqmXZ4H9i4/zDZD1rSnfWYuyxdrheXZmAwEe14WLfKYeOxCFk+sNGMttvl1l7ewslHMpyWD12C
pHOBOjmiYASu/NJHbH2NPAaUPdCWv9oT/r8emEYvZnunBqfW6+pARKIiEMBIrto0INfOp9yeOlAj
+mguPCFphjERc1eSvB77xIljG6Fj8cCLAMukhUUrkNen68sJrxbAs5zjBNdMus1KPDBefENTt2eR
dQBi9sgESUU56N81q0MWaIcg3EYp79cmb+V9qDIa1VmE4swN8i2caN5VrBan73uJjV3zlt3mcDew
YUOX0jNHpEvDEdFVhofngf6A3eqkdjTk9oghxoaPCfV0fHOjYoFTiVyA2Nd3OCFetYV2JpFdKki5
AEqciPT2tXoqpXKaBDqKZMYGsuZILH1KMdz0/Kxz/6WuwYiAQO2YfwAdHD/9z8x0U23lj8C4qdtL
ghHXG3P1A59FbKUaVOBSNd+SVi8gp3oW0IQX1NtlE8llF/2PcITm9VdubtOp56bo4slcWZ/eoEDr
9Na5VtMjzCZAnoE6XqhszFqjelwRe5wkR5TkSy8UH44ke15NOnf4e6ykIY9MSm2ihqVjIytBeXaQ
7d4pjdR+2D7zFJm9IlZ8fiQMpGkj7TXgsF1GKgNVqU9UayqPRxf16OHGRL6Kw22Frt2fV1i/Hf0j
SK/0n6yBpMaa9HJj0fI/6zgaIu3WTh9p+4AjonQH1/cX5PS9gT1aeMImQeT3x6b4xmcvsL58xyLe
LtKbpZ+DZe51FSxONLiMYyxmPfAe+N3ufZSTGNq7Vz7wFwVDvk1LTXk+7YkZPPX8Nm02POiyVrG6
s/FpzZoNzbX0lAdYaM6wwN7U4zvHUM6wcqWuu9svLPJmcpBCuBUUCSdx+/X+42/5pcJQ2xNfhz9J
+1eCOLKYsh5ETXk0bJEG+RHUDFg8++acJdqN01E7XiugdYvQaYq6XwdKRnx/yMLlxfUQ6jtcS/Pe
SfGHf6Yyyndqp4Msd91zYb/Dudo5wiz7iXNtKbtlN0EkGFNWD65aUfFxbmzRrzTRctm/LqG3ZKhr
YyiqM1DjZ+ISSzpKM23UCoEj7Bqef8JEv3yD64+Cf7WAkqqjFWzedxQRV72t1Ov3aYWZsvLDmRTm
tKDUipsGlkHL0p+h4PeoAkpRaMSFWGiWCc/Hw/tdDwmrv4w2rcdchlb3s3pvFxewpyGUsJMyujwh
X0LPeLRCMvDl6NqaIFXOl7MmrSbGHf5KLQUNuY9M3upNeQ5EjaGdTbkIxNfVri6t4VzyjPvA109g
g5oimwwdqyhsD3MFtKgb6k8QIEbijOo2WPnA9w4vXZl6Ls+anW7F94ZLUILapvhH4xUJ8hJ5lq8b
TIZ0n1CcsTrD/GBPmcCAhIxrU+e6CpYOxOBjMGTPbwFJ9rfRQLk+DVq+zC0yR9NLqIF7oQsMCoUq
M4fxPs0CjQqsTzbThJxiIRqLoBeTM7AIp8AP+PC6AsDdu6NpEWaXhoyDcZVYOQD2pNmvxy7SnPeP
6jWZr65GuFDDroyEkHRB9fGFyG6A9ql9l3wVfDll1mbY+t2D6TNC/6BXLRXD3HMe6BdEJexyszJK
eDNijLLmp+rGvz/7sqjb5A1J2N2jxNRLfIB2Pq4BZ9JEeh2toAQ1HBQNtWU8LMagRrBTgAWeKKtq
25vQ3rboUbID3R9JKqA4Sco/m6sy/2zu+S26qbz+vE+5HyGJ2s2/G6clyuipzwXMTGPTIn8LobMX
GZtEIeAUHG+TXiWE8c/whFXdXkPOOY/ASkzz0CT2x1YahRw0wpGGcViSB91yERBk5FwUW9IC/hZO
2plIEanNeeDfZ8Q6VklmkZnOXO0phd0o7BSoiA6r7pcSwrytSpY1GkJ6eJ918Omd95zReh2zNdi3
k/4MpnR0Bsa/M3xMKQ3Aoj7ir5bXgrP+tPXTcsVeWWyv7E+ucSd0zIxaqPmwkfg1NglwHqW1BVr8
BhVH8f/3H/eiL+cCyxx6NyrYWP+oJNRBH+871Ja4zMeS9XUSQ5QvItiR2hiSyhcZq9ORrn8I6G28
/mVwDeTLbBXGePDLxQfnDaWuOyo4yjvY0a63MapcH6NNdm2rMICCof1zoORMO75SUpC9MGgAhAKk
qqyfgJ10gvC+5mJjumrelpkyyoMW/6FxYzUpWGbqqD5YEIubjPzovN5rjvS0kjs44W+/SxyRUOuO
WeE7q0dNNJLP5U2Sr8vkBshvebwWmUusxIO6UzKzZyspHFsi8XUMzHkzkQ75t9FtoRPmn3UgBtzh
+Cl6NNN2TK/Bf2p1M3BBLqGtnxesg7C27XsjH66iLP2zQY7fTtPkikKM3U+OdrW/fIX+GEE6QCCS
qWGyKqP51QUOwEYjGy8ns7TUfD43ERlbU2EhahtbyDfQFCijzq+FyW770tlniVeQ/878MmIwUBZa
9pBeTRnhlaSl1nKQja/HQktYArEm6kMpWxLtX4u7O7AluDL/uU5W0LjpvtKtMiYASM8s11zFl63x
Nc853oY7+y/sMGXlbxqjUVvOum2PcE8tKXnkRWrr+w6bmfw4dIj8dIBRuwgFDJ4X0otaYTiZqZ1h
83s+DUn3RI62lTIDv8Ml3pIU4AnzK1vVL+bkjP7QFmkotYXkcqYrbttdLLvDVIffAifzTSjDYr8j
xmX93jY0ASsPOcjhapQXKqBfalf9AXtVilzUXqExGUn+V/+rj9ztx5+cEyq8zY0dzTjj9OifvGoI
9K9prgmIp7+gohsW5yr+ijc+ROH/vaAy5KdlYQWoyPkflc3uEf4SqAUqJNuFsDNx2AF4cQQIlqxs
9oJGO/v98U6ZuH8YFubyUhcPHeD7+UUegXjS5YIxByUEsDl0O394Ga7gQ+bLkEySagG6I9yV/887
D4MuwerVS9eaC8GEiQtr48Z/TTt+ssM65B0Vex/JlaDqDgHdrEpBVRunWnQwZhmJ2gIk5iTFB980
i8o9YS/RGiykWxjTjTtJY8Et2mrdMtWrWZ8CWl7242yi8a0trtwDHRMnFASyKpN2ZMtEnFuR4uNo
UDomLMkjt5XwOkbgY/415ogxYTvcm/GQMhJ4CIqtKCKjUcn4cbRt521lNN32CxHV2Layz2TUN6wq
rknYe1JFHHWxjr57amwO9VhMwm2jX0dCWo4h4BUnELN8f6Z6JJP5nY4ZCUlkg0oq9lMl4Ac2usqF
CSVGc1nHyfIl6FUo/akOl6Xiv7hWy7YnouH6F99nO0w7u+9E411u3Vh/waN26co6io4U8XUEnQQQ
nNEInHTOYr+mxwjeHT9aas7gjTV3TB9ExLZbJOTGqI3qDB+4b2wkI3KzXQgp/SGLDYTcZHwHKwg2
B3anJRK3Dx9LxS3RBgIsWnvs+wgFOXmLTJ/BPYr8dS++5Ta5Ij8Ud94N6fWIfPFublI2bXsR1+RN
Et+HPqoenbqkG1AIKwGELqbuoMWm2IfnehAdRfUvxAiT169XgFbjEdqopvif6RlNzOl18D4YvH6D
kcL1OK+SyCwv84u8HjR4nt+mombMcYIm++IXfmf3LHYJjk1ZZvsSSgYPG9BIqy9M4WWA338LO+Yp
hiNvk1cFRJjeqUW1oZv9naBjQcMNK8adBiwhZLmvnTvKjqpiOl147Pw6U2fnBYunv719wD8Z2GaR
dehCHKm+mCdsVhqA+8YLCnlCKdGH04HAnNUffAGgszx0r4vXlAUgbU6SU4c5JWtiS/p0LMiyZ9G7
43sDjGwoKepw3dCiiJz19JdhzA5muwAvk4LZP7TgAC5fzAPYIKB3dZiw4lohW6o5Q/tBoByxrf1X
u+Y3pH6ivU3CkLMm5gxJKsw3j4iHk2T4jY0fhySr6NB1w8FdGvltILXkk+rAnZSun1DhQLg/zN68
r2edrbCIfZxhGPoY7JWLfBZDizD1bj4cuFecu14aM8IHVDFqOPcsN80JVW1F3ugQP+Vhvnw0GCRA
IIN96Y1sTtaN1FgeDo9CelNOy32OAy6xTa6b+ESVGJfiAG+A9VyiNU9GEX0d48cGcFhZHQBuW+Mv
KqJzSDzO+7+2P4f2iUWu8lhyPzfIvLrcWxPEpZRs4q3wPXhTIyFoeKvtK2jzsgr+3gBLeW5HwvLE
wL4gPN+detml9/MmthzH57R8Gr2KUDMS3QpQYsni2YKlPO2uHjN6ySZZMI/F/Z6FYunpBrh4c3/i
/N6g2fXIht6biwPyLvJyjqx1YON4Q2qmiZwm7hwlTJ7Y6mohNI8pTi8QIiTulvXRoy52rRbExPFl
NAz12lRV+gNAQ7WX4dlvyDA4P/3BYzhZDmFqfUZSxlplzFlBffzLoTG98iBuG2ovVNh3XYilmhza
2qtTkR0iWj9kQ+O/goy83FvrZIFho03BSA7Kt5/o1OsV1UFv+JDmWMmMePAcENt7OCrxLkgpq8Em
MzLivnr1wcA0rbKZQpf+HJTjH+hT9Ogky3NG5gDuPsy1mgCRxnDwrimfujBzYuR5UL6bIWlcoXz7
VfohZRAZYni2HJ1oOSjQWMlf6v2ih6VTZb8kV1PhFoy+e0pLkHL+uoLZr4hHIEh6u+L9So6Awsft
627o1UDvWLu5EYgYeLsXlmEJpZt/rSJRI7ve/vaG7UFzG5eSrCPCeDzZz77QzCUkA8K4lOmZw8b/
u424VNXWTg30sWn30ZbONyPFSpprpRBR845FNvO84iqzo3Tbbu03b3vWfhlANRl0cCoYZcd/4wIg
+MqNIjqVm64uvFh7At4hvH6NbyfetCj3bGPUUANp/LxtCCR5dExOLpenv7SXyVM38IRLIWMJEauh
gY+31YPLcruyhfsf3j3MVqsWub7ahbesOgAercg869HxZxHDDT9kSh7hxnM/NvI56X7LuZ6NA52a
Dyg+D1KHSi5g7OPh0NzULrh141kde5RdaNi3yF7RCnkJX3voc/lrYhVQz9czybDBNHfLi+muAMLd
auIHyToIaARQ8ajcQGbqsvgPWD2KRlFV9tP0kFStbj0KwRwCmyvCz8fdJ6nmamJqFMgP87Ma8E1a
wwhNdIcEdWjKGJeJm0bG21qpnRoYVCDBfuW3MlpKxZeLkVtqkha19tUVraYzyImv07IV3gt3Q3uz
B6jjngexReVqRgbLXpmKlFyC94Kidl2+0BZM0eEwFzRlDBYisX/vTYyqzoy6m/tRS8ZRjYloN2Xv
Kxs7GRpof99wIHcWAbao7uJ7IZ5PzIF8rG0aYSfo4wZjMf3vPCEq3prVCfjmobR6656GAf4C1kc6
ZfGZT6qThp3zl4FzcnfSa+CPy2TsH3tB1E5VilaOYEClhdqbtWju+3lBNPFPODg+fn3cSTb7Ul+W
1b9kI644BhsB4PZNkrtAdJB7sV0lvOpebwu3C6zHTroBol1UlN0hLJGJMpUY4TbLXIdAp27KOkxn
6G849MCri7DGaja1RFt2xzwcSLm8BAfSMO+deQtSuI/yGdj7i6wBqG0lkRKg9xY1e+pSU+auichY
d9Gpkhj3Fe76FtOvz72li9IkxAt47vjauUTKeYa8QMDKe5oN3gwfBJNPTl9ZZemjnWVP3WNVYi0P
NRo35ZRqW6cV3apbRipgqv0WC2kcX4m+z3HZTkgCIbPaple2PTcyE8VTgmDVGoY1MWuRSzq0ZZwY
ZQo6Ai37oY1QCFdrk1rKnPejQLPFAS3Ysg1A/Y5jBRyO9WRhC/okgrLWKen83Ooy0bBWttmhR0Hm
n30kiipGKcbu3+yMgS1CV+lVmxTYyTjDgT9Xsfqk3FgeYu1BML0TBrHnWjBBsPH96/lPE301WupU
kFLMIKKIXHs+H4ZoKa5wqdqcLoImZE8/3sgclT0LAdG/PXBj8bi78hkcVvckGSP2+397WTH5WqlG
Va7y220xE8Vloc4sgOd6f4KRJLxYzMCiVWfFx/gI7fU8lasXnkte3QYAF4xGe41Ix2bO+wUwfOcw
aULPxEmbafR8nj28rfSDe8cSvJdT68hku+bfT07ff7bjCVarljTFgHbnNnk1wKzERMEAoJnIb/uH
w5ZL+az9ySjnf4gw9ZIvWm0FINF3q7V0b968lbr+52OSKnvIV5ko7FtSqn3ujbMI2rQDVmetkxry
jXF3ud3ogWHH8ecRrU8Q+8y15amUxlfJm8ObyJHxADy/I6lT66/aoY1GodWJUxaemHmbv6xD5/bR
GCkO6u6QSO0KAmKdWsOL9/Hfo3ShrIQ1oQSrOH+pX3ZNm4RjVgOkFW5xPUb0erjKWSgk7jspGb3g
CTV2nPqFJEn7jV6JZLtBFieuETbMfJ7pnvgHXd+jIG1Pozecnea/dPy3E65ry34kNIBZYBcVtl0S
992G8i847NytvpwQ2KhSh9Oglsy7P1bAxNVZb9ojtQJnt2Z5kSdpmD3KIjRqPXO3oEGshjR6M7Ck
vevmN9xn/f8KeNSZHqAgIVlCuon0b2PWB7CbVZDzPkWm0gsA5kX8jWFEFqeuV2NBZhY+O8WWc41j
F8Eu3TUFdN1pZnk39XLDwjN5ZzJrRcKb0VfDgkrs9lO9247cTapUO4WApUbSrrvd5GzWgxjbCV7u
PqXsFo9+P+n/irfxW/lwYxKunGN6sX9rSSSJZJRsaZnL0w/KHj7pB7H6PV6YrAi+SKR6j2/GPYRf
tmzDLt8sL0m6K9sRsVxrQe3p5A9T0Fjl1w34ibMO9aD2wep4v+h4TlK41MwgxB1qwjTnTlFgkRkc
h9Yw0KZbxoC6IlmbEDhJ+apLfv3O5RrVNof+oya7b+bdyfuUYlKcWAcbwvd6w4zjKj37pg8hY3TA
FmjuvdWYcwaGL4QNb0mJnQWFdrRXRvnZPfNjlJkcyOvxGjg3JMlHbbcT3/Qh2CcE4dvEbVJmcil6
3mwqlIRYBM9t1PbDOh3tPxcenWVHJhca+J4rV4DJWjAwepwzNGRDTUJCAeT02/V6LjDsazKKky/B
PmXKHPVv5QEFzPs/e+kA6DAeCO29vQIl2SLY7z4hncc9j4+i0IVrl13PMMcxvFbtW5wybKQ84k/B
JOiLItyD1s39vPzxGNktMUpSFvrtj2LlWLC0NFLhR39nLzg3FYKrIW17aGLpQ84PV1H8CDiW4Xxu
R+q4w8MGA8X3Qcgf/9POwIxg+9BIHDbakelxZ/dH+V3l/kAdvg9YXtZ78a6AtqA3jhAFkLhvwqhQ
6jc8hA9Qr+hc9dyuiItU5E8Zl4ja/RWyXW9XUmlAnUE1+QbNU2mdCUZ2t4YEb21lTAa4h/zOt++G
X2mS8GBsh+tvkrt19jxCLGP0lh+w4deERtBAgrUYipmGwLH7KEW5+gtlJXZSryQJU6tDaqphEmum
jdmz4WZwvrYFjDNRCiDLLw8V0XKRprj7ASWc5znUw5lcOaBSnsTwkGePRvH5zygbsSDQTZdyFhuW
h+G3gPViShUk2C5UfzQPzf0XhE74sUvQFyRZBgdukDR4LPwf23OrMny5ohjsQGEMZA0HtFZgBTRT
YBRUXBduNRRMDm+k3awV7odSDK0h7SVfyp9+5Pw0OAJqoO6hb0YigGAbib2k5yKA0R4qvQ72jbU5
a8R6c1QzVmJDe7QMGCVa9XVrQrnjd+KLGmFAbR721iAnh1a8OjyMPAgqMMVyMDgNQMfLUWS9ZuWk
gv0tXi/sBzov9wfIytt5ZPOAMJD9Or2CK38lfWzWBAERfSjodFryg8SZUvvFFpmGNbbokNhq+bb6
Qi434dSUiPx/4sSBJoqfYKqxW99648yyPZGSekJji/F6BlWJZMSBJ1I2lrGCPAtPfylA6LIPmG7h
8C/DMHOp0h6LBgpYn8LUoJmEsbKc7UYlA0s4oEIvM3koUZbuG9luXWb6U34k7yVKQKlS6QYZi0qS
4iK0tauHipoPMnU9JMzYY82gcC1FcWJUs4p58DxfqdRPggLkGyFULP6xWkN3JVJN7vUKe1mtlFTp
OlbTGAE6/XQ0yUmtVv6eD/FO/zT9QrMhtPuB4WJSdvILyE2ft3AogeVP1KuWFNc9xBMxEHcE541j
BdsQimuRtx3l0MnxBpkaWgSR/9KawpRW32tVLnmQcTdhQF3V6FAxQR5Snb5jAlt6NqBJ1oYmNK6h
bGnRnwXqJJwcFa2Yeniu51zxSge7rDveA+Dgg3k9bbEY0X5Ua8lpUNUi2ctaCS5Xy2aFmS1Dut6r
elNZw+bZ0IFSxtLt8PKh3umUOL9wcdrUed0BVplqYvzAHYbvNMDXuf3UyOQYaygMQEireiL/8/cl
Cb4mv+MAHiDMoiHgwZwD999LcMeMED1QarhHSaa8D3oZw3tmveC7Cugs1SNAzbwYF99F1Y/ktwQy
fTpPDhy6JlvNd85CM7n786es0srwMXDB5+Ob9puTlUGKtczpcSrSo/5o8S/epWEl0361How/4tC5
cwqjyHdjzRnAIncnsMcPRBtBrf2vjvxvAg4K4Iluk3VhJNWOCrEnvXUG1PLgWrsn74FP8VclXJSJ
2thfZXpYOYLo0xDT/a+MDCVk+mtaXxttnr2osnI33WQafe41PhpfTvqbNE8w6YuVU7UBbre247YW
iSkm3EWuVe7imn0Wil1FexUaeYtCEoj7hFhyIiMQDtkgqu+rMJLhFXTJirx6Z1i22clWAzkuTtPI
EG2xJIf1OBKYUKAoCt+JN+LB0Wgl3Vgjv/wEGayRf1dhvCnyk74Xxp7xSH+b2Pvx1TC8k7qNEW8K
CwlVnwJlGNdAA4mobkdIr3aP6m1KJkrWk0MfRW6jFvy9i3CGehFawXNT2Llu0Sqwv/lRpoLKamh5
xXOKpfgjxG4Hz+0dMEBrxfqy/UeZNzdJzx+7hRUDr6mESOOG1reHSdjG14ReSbgWBqnTxDo/4WTz
WjFUr4Hz6kyxlZ4j9WP5M8DgJ1Zw3Auo3drb9BodfMDg0GxwrGW8p9xIAlfNB/k6we7Q343CVa54
VlZGtCFOFyD8gN8IVFP1tfJPxuWFH9CGf3LX32adRSrY+7giOtahnxX4RO4HY8+v1+VrBG6UGK7r
RhvqpV72YAkWe8OuQgopE/ZAm2g5Sp4jssu+0xErBI1zzFEGWwR/If0rqP/xZ+N4KICDecY8++ew
3o/cNpPW8slN+YrKh5foJs2K0baY8aoiq/U77lEEk1msSF3SbyAzSFp+8zAtJ9IWiSE+0G8bsQmV
7Lbbptfs4fRr/w2/A3YdBg+wj6LoNArFkzqHT8lD4ZH7On1JBxJe1tg7rHveJkbs9n2On3knvKJG
A5Pi2b5joWYCmFGbEVIm58lHcQsmV9iESsY6bc/2EGBCivvHGkveZmAKVmnGyKWieZAygE9PtMu6
hZreNXa5GqbE48Z16ONtKEZU5hxn2cHaR7MYlZ8+rRlN1NtbMMNBxtfb/FPdY+/g7xhuSpKF1may
5D50Auo7jbYoevIqCZ8MVxBkS4X4UOE9rjDqznalE8cuBbf3ASXpPy5MisGtdjmP6K55xjvYoHcX
06Ht8/TY8apguZf41IpIf0+AG890ksE4ZUgybcDylagg+BxQ8lmo6Je7vT3DIPsyEB+ULzUlN1+s
92iMR0o7qqSmYIRRi+YDJng13kVflT99P2hDHXQhbKekIRYetnmvQnS5qqBRSccEDctGcFnuDjc7
ZvFhtIrOpwxjVQxu7P+kTzwx6xTSmwT7EJgQDxfMnVR1QRk3tSlbomvqTBkPqPZQqIIrUao93rMq
UgjWZUwzGzzQ2CTd5F2+rd2LNp2Yc6W1jkoFkIKd2Mr1zwr0DsCIcxwKcUU+CiiIesvxgH6OElFG
4Tz5EeGGfzVLkbVAyDYG3jSaZ/dya7JsHwt0wp/5qI66vJZq3cEjqUnYrmIMy0y3cDoq9G0qXRyn
0bWvQi56vktquXY5wEDlSpoL5vzJ9k7gFHpsk3o7NSQXrZdJHw+SM816ntffaZ6i1aYdIrl2xqY7
Sr8Eg2fMvu3/H8PNa87h/HuGsWBpV9jsFFK4gVCdk3tRndwmhJcp8dssvtyI/T+ZXG5f4ylD3/GE
pFfXr3MhmcD6yECcheVgOa1ehdGYEzkJgj2rQ1462HyCDHVqJwVyHdVy/M8nsXNCx04DjPdyFxku
6FQqb2WkwbIy24YwzQ+u5ex5L5gXHRbCvOPweJv0KjjA5HUyAP7JCL1RTrt9Zm42LCeQZGIvD1FX
akVNqj1OiPYVHNrLc1SqYLV2Z5V4YhPmduEbHQMM3KKSHlabbiRUtn9aYBZzOMLn4h2lJrgY8juh
FibzIl1GXvf7Wi1UwY4J18UPb5OA079oduVwzX8Ihr0qLWFZkDf1+yMzqAnHd5IepO0UcFF6MNv7
w2V+X9oVyQ8eup6GazdY7pIVS7Kbe3q3MFLzs9U4o8Bj85rAtw/xLAwRx+2fQA1aTNEhkeGnmS3k
FZnxDLScNNg6pdavN94D+8FRSXUeZiBvhcmtpEVhnmZ/jVMWuVml9TEUkSQm2cCe3WZlgJUyfwqK
EIniJ89H+Rd2H0gPXeVOLMPHlDDDjHFcaoTP/ZrWtt3Rsm0Wn6mzG4fcW0Uxt/Mqs+TqpeVitjhd
YULoYCIL/WUmopUSPdm+zueWhkisJ3XH6eimJtDeK+1m0cqgmQzNeKD4EYhXlicTONfqgEhntlYe
qTP4Fl9o2l44zQsC9bnFb8gV/bXRugv3gBXWrhFKu5Y0uSuDJW8BITKZ5Qt3XbnNwtokTvx9QGjS
J1hFOA2EhdhXnYJFHM2TIrfO3r0xff+A9lRSI7cycsSPiYoFk63hZ+Sq4ITSzMtsZnKCeyo7bPqZ
uT4EqwNcU1C/IJ33wy8sa+jTFUpcQSNXuBfVLiSd9SN+XFsyKjKwBxsV+PrTrbIfmkDZjKJYQ2G/
stNfVr3HREmLk0tI3zcqGTp3d0gA936b2pZG2TftWnfPH5xujWqV6KdCh0VQxuRgoE8+d2y6jknM
SzliP4VrSb5mYc1ADFUPIrddy7KnNErlB3PlqRgxnddYyF69I5Dt4CRuRGory1MN4Twt/HZ6HC2X
va/rTm01bR22h3zJeaB7l00DJS/G7BE7r0q9r9nGHX/uxCI0LB8ukPV3HbAEjfAS2hzeKmta0BiC
tVDjhdJ3ZUA2Cd8GTb+5sToybiegkt83R+mV6qinRyQVRcg0ZQlynXquRZeOSHt+cChaG9F8KUlT
Wl4i4fB+wptsX+hFK8AxXIpsUqoUb235ogdqr4/J+aac0j4HYePTISJYmn0bQ9o5a2LD91tJWf+Y
+DvHkeYqURi1jB9l41bYYWx2jB5O0zIaGOg/sjdUwqGxpcPPkfup6yYaQlPmr8aUXgXRRnt6o7pp
c8JuvyoJYKp/UE3m53++EeFNhC1eUNz2yyT0jJvm7z/1oUvnu0+Y3w1rrbiy5OaRq9YVjvd3i1DT
e/sI7VUli/LQk+ktTkJZzJD9P0jq7Nz2MDAq5dxZC/qN09VxwvHvis6hBULEFJUBf65l6pS2k5gj
ZIRzS9co062cjUtIVif4hPgnMA7P5rLg8aqtMfCdAVERCIeIvNKNcUpdDoan+jyiP5GSgX3q1N7z
n7tjm6m5sP/EWvgwhLIk4vQLUi092c3fCPytYwwBn54nH3/spEF+sbShl8h2DYb3HT+L++u+zaso
g573MzaTR6bhr2bbPW2ysKH7GlWwdGw1HUB6npQl1foFwtbF8pzP2t6gQEGDSXM7ly0AVwt9ctV+
coMc7tqZnvYZ8lKfNFnyCaEjbJXmVlsShxz2XSyvis5n+155OZixZuMoXLg0MZK1Pg0ILo6LvEjz
ScpRorpSw0ECWo2YtHrS3i5ebDBqcYatWDX2VRCxnKSQ8XOSufDwA/KLl4hxR6+IvpIexQ70VwE5
Du1tFrL7j/t5+/4k0vRZOcj8QbquHrnsznCP0HJNRsMpiXzqobg7eQHaYS065wpoG8h52k+xGaIV
nItijKOBqrPXoYODrrpKaIasPRdkFS+j1K7yxTupDawTh+NBB4oehqsXf18oOf+ppA/+vfeNJDMg
bichrLRiTREURx5fdaOZBZADhU2d1Zw+idt61ZBshIk2FO61AKBEpTlFVpq1ExMzOzTWRLf/4927
m8cA3KLA1HcCBHoV30fWh7hcsoyY37Lofn4nZcTiOiglglmXegMt5eSohep03rMKqzZ57kVyDKPi
ZOVfBUbUwiHJnyQdRXAAATHhxNOAFe8UbjFxn6Wv3vEsoh5twIFGAVa5RfbeyiU5xOKxesJM/CfE
clBrWbYXFI2zgtRPDGwoANRbYeU3G2HQ35ewFXOR6E8K1Gf/96UiWK3W9Dgq/kIXtJxaT4MnRaXP
9Nv7NJrj4tTQbtcLjSEVKIK9mGqzvngR3PP55E4bXSGhr+xj91nbRGUZM/PJGUtWETpwwCkdKtmz
DWuv0Awi0fEG6qxoXcHJ5nnd7F9ZS3hE+eJnSRbmHCL5efFO/koi2URhbIkxju6CRORxp6nQhaRh
kkw8H+5RgLZTA2znObsN09XO2Hfv+qvD0c+30xV5m58Y1Crz4X8j6+kXtcQTC7nDXJW2WtvZcwyM
xWmvSnQIZ7Z/hBd8UWBoe+xmd+1KTDH5GD92mFFNIPyUAn9F/vqglvbgLf/4FQRzS4Zs3t457lQx
aRJiXl2LOHC03OcDfnEPug7wiMh4QTu86Fc0/g017wZyWCTEeASsPN2C0Z4+Rdjs+0arxJJ0C2K6
PdN11814SAX+NiByR6oLwXvIhKK2+xywV+qUe8XJjgUKpaBeZ0CNp21wSWpN4NKLXvSUmnXD5pFB
LjWAEYpdk/3fC5JgnmBz3m9StR6fjEo6NZ2QLMUwKBSEJR+HIdN1BMOrXRwNqr3+JechwIvQLvdQ
OGpKGySs0UR8x63utOLJJJESfyRQGDfchTxRtOLhb9PQhS9WDdG4LUWmWd+BL8gs3MtOry3pVEqY
mep/niIl+N+jRvmTU1qsOWcF3odqc+Ay5Nia2tpm0ExH/HDbDVLu3VG6hZfKbx/RAtnYaxnX5B5U
k2i3edeaPp5YU2n/9PpetOD/bDtj4DObl7U0NrE6TBPx+PriTSKmXm/9LMtpkpB19X9VBtfajJXD
zf5C0dxMxaXq4jEK+Ep8RCWhplwQPgD+e1wrv+bCiO7Au1IvMI1bzE7EV9D3CO/bdjP2Nk1hpy9c
2z3zvk4aUovvHnRXLVlqX+/Eekzjt2yCIpGXnqZzp6xzgJHIn+ShSC9V4F/LewnAo7Y62uBxgqDm
Iuc7yKPYZ6XRIzRjwhFkoYqdxM1Fx+P313D4YdsG4tGG76CfidK1oKsB3+bls1fTxLWbjPz3GVWK
xJoCYwNh5x19CGKvsBKTKkesQlvIr15EzlQtdjkNkU5UmGqniJd5wxez5H7jKYkGrt+3ZCh96UVk
gxUcCb/8z1/XoqulnSUaxT3eP8FTZ+GUT77sNUnN9WTW2UoEsGfeeuKwkXq4acXkFnsBXqsOwsG/
nly1mxnOxFN9n1U2KblYgeZgeAPE7Ymg5xRBE/seER8ST2guQdYSZ9xtjwwI6Qzc8F/w/i3Bzt/x
ZjdFEVnxv94jBwUwa+h/wRrydoIUrEmIUVqjaHy6MffjUmwuMFYnxJxWgYObgjEyfvHaeO+8BQSU
g90fJktzcpdf3bNL8C4mijwNHy8tasnGH+XHSbi0HRwCcEXegekf2wmAVphBWf5xn8QPWVf39Szj
WATeg4b8C8HCQm21x36wI3Hsc4OFUct372SDcT0yK3rGIYD7InZ1ocBR5BX/WdUzvRf4SJkPjC7P
0esfP+8oc8EmNln5uFZ+a+yiTGXks1YDY2VxCGFjubEgZjdxqJ21XRJyDexzQbZhvADc6gVlkbbX
2bFuBxVZc64nQY52tdjQWwlYNIguf27ra1gGXuZQlzVqpsIJxCXOOvj49sesAfElv+3UWM1aQzTO
3RIrUFEJzsQlAhWDAA3WhxM+sbPwh0emDyEqnR08fngB3scLuqTR+Vlr1o5kFhFa4AAXZs6TpoGE
sTJbTL7kfe9e0K53lHldMI4QikGG0BBZirrzIKPHv8S/irbFcJGZx1AmUDq29KyhVkZh7N+Bxv1m
OXw2HZ3vnyjkf6TRUxLT4Ny483a8AWFm7lIT3xxmzeimEMb9k6BwMkl4kPfNx/8Fl16PZHHp3D7S
tU7vC/wf9LAhFKFIJ9KVhUCuiHZu84ekgeIT9uT1nJCEPfU5cEf/PYZJL77YgrIxVu39T9bFmRUj
Mkm3zS7QOVCmazt/p3d2s0p5QCwetsrdYpktLqNqtgfKWuW5NUa6TBFVenVtE1JrTq0KVXGDkXvf
BbB8P1tEf5bnLfPmBIVOnKqQ+ivfgGDLYDcsvCgnKwoBqSDng614fGl2q8weRfAmxtxBpnhFpcMG
USK2SXvRVRJyIpGdot50dBhvdY0TXacov9yVtYCtk6AWYvEqhzpi6BcerX74lm5Or8tzGTmeVaom
VqlS2UWLXTwyXPqzgHAN+FTjx/BF6XtffdnawSpcJSclHME5ELCk3LxXnk7j3FqYhq0Vt0VEgZJY
+zi0Nj33+xf3sCF7lbtYFVdesbY/vSOb0ovpTTFxnQiW1XNltaO+z3OdhFQlu5XSkAhyaMqnpWG8
INLKSbHYQt4fykQib4iDg8Q+v/V8j30rSThzf1Uq5nphSMhCzbmCNyVrLXrzI2OJw3qCFq0yOqEU
gdq5kKr48Y35UEH3V6LT/8v3drxs5MZK6GOHRlBnsbwK2JMDmEMGxHQgwMMfLUYoDZXe31pNKVQY
Eyy0oJJ42roauDqc/+hglphyzMFpC3JHhuRIp3dqI/JvUF0WTKW8r8JKbIRWKXg40Bv2veorbPEm
SHRAgidMJ5QGRiLg/c6ubxtmFJH2eRStDAt1zPwwqa7tmT8fVM8gYRhDtWIYqYgk0zMKV72io0A7
iqU6r9GNFzfEJD+/3r2WIuTtl3rhitM14S0ur8/Xx9j8ROJXrJOOcuWGp2qttVpZEoREXYj1G8W0
HKDgadPBxpZmkYel+iAfxINzYuSdtoFaP1rWJsvVERmFbAe0g6gFZdf6u/TcUveyUS51RmF2AEJT
9pTM6EAntj2qt/PNuVU6G6xZWZTAYDCZ0PMSkEgBo0fITWfkh/kTVwsI/hYKzxPwQGX55+KGLjRC
VmO5t8DCjOlUNpEQZn5tu32Szyc4kGU0BlTV5MFOpQL1VDmDO+BmcZG+rNLcGAh2PZINcQXdQuSz
mu8C+yfpEgOQ9mXDCPwqPTII6bIOqC6B8cQFkFZeqNN2kaqwwg/58VodnbsfBAPRlJCusjQNFs2O
ppGT7yjpBu9xaeqPi8X/nZVIuUovcvHeGSanjlLypNwWq3zr1gWIaZrvjVaoNKgCM9bzPVvkYx+9
RWsTLkgJAXc61ZVupZMffef6kF3+jW/8HRSCCp468hZNUs6CgMgtf+tQQbmR9y5QsrwDAlp+WsTr
C7KPPdt29KZVV7KENw59wCBZafpbpWxRELpE2Iu2NfM75ACZPXkqii8wzSlGW+CyrSJkAkC0bRnf
ZnlEXZNZLIdDRaZ16fqg7oECpS6Bf9kYhvT0in4N51kPKDtwVw5kNX4TAa4NvWiqVjzSQ4XHBOnH
8d29Ch7z5Kl47xs1iE8gqTFynhmYlpBvdGtBVCTjxi8Lik2jrAuMRVGcDd+XZ4AXMLM9Em06mGRm
KKGbHZeE7pMe6zzG8g5rvXDpyzLyp+zOly7l2mtjU3GFRQ8PMhg9gKt70jWKNO5z8nB8hpzJ4K4S
B/8PdZMkxzY7jRiCPWLCyVRcjK5bMfNeDuRFGt3SL846sUSdZ3bgjcjjFgJjllb3zpCBJSajSPWD
SPIG7sW3cDj3NURu2sNCnRfXXmGt7v9489Qrtnnt520ioYmkDZV456XcwILtBsT+/QkWyCFMY33T
smm3ikRa7JAQssbwiCDWw6SwOoDEmA1qlK2dwVcT+etdVeyXT7ZVhGqgV1G6PaZzBK4QxlY6IAwv
8qoQ9TQqfkUZ8SUBmS8xWHFzLmEKYo3IzqNNHHG1HtEtZ8ic/3S/ON1Wcu6fiGUb7wFAR8IWqC9t
Xg93nAiAAoOhxO0H5Eyja1qjPOHd3WHx6einrUUlbrS32fjfQ/tfcDugV9ijnZ1ZcDHizNm9HHAE
1W2Me1oWAUfdEWTGtmqwu2yy6YBLa9LtIUL3eJSwq0jKG03pAI6qRscEWwYkGftZW+9CWMa6I9FU
235uFaHgkvpZ73XrS+PbUm/tL6bzbKVc4LD49Xqdscfpfmljml87oMJV3sB6jsyDXROa8XjwL2B+
MGF9Sk9ht8Zww+UkcAyM22c1Os2CLO6vXF5Ifavyqqzi7xbVlluNvo4YWprXLMLnTiB1ScF7agKK
ySiDiLqAtLTNtRGYcAeVzcB3MdwnuyjtEIaeosyUGJU0jsydX40OiN0qAReS/PqM9FXTm3/mu6xU
2f+CLTYLpC6OcYfYN1aZW0ZK/MigKhEjtS9FaOnUTR9Tz/a3zBxkfRqiHovEeSOSsCegawytfsq4
DPVhUdr0hM5AajHurlKxmSyuEsOCu6DIJvB0J0uDXBeQOaDw+mIWGZcBlzC3spweCl61OFa7bFC6
s5H0u6A9YusNA7gbGwzGPWOXECHXIrk7iwW53HJQ+ntGPDyJCZC9k8fL8ZwJ+S0gWZjk8sRsXUT/
pcIJp4QhXa6oFJAwky/MZs+6dHuV48XBtpaDSpxwXAhIWSu/PhNEwtD6lfmDrM6S4Wqij536Ca01
9p/Pi5wBWJ9xBuWF5cUWmZKbu+/ZMAGe/60Y5fsbRE+Wg+a59HiMfyeo5568xaTrI183S9+GOGzL
QfYCNHlZzBudzC04vEC7PWek/N3GvNcYaXuedhZVlR6rSLYymowtEQJ8o9LHbMBnA3CdGgxVdKpV
oAssDm+mZZLBdW8jpQGLBTij++PP8Drmg3mWR/wf8Q4fF/rqAm23b4uqurB7b4rnRyLd5JijVJKm
wnkt7lfoed1hoNnrgb9f+rFE6SEuyP8oxp2qVOBqymGsSMZCV1PQ20/hramCm8Lg4OfG7o9pO8PQ
fIZmpe7d3cZ37xNu84leQx3CxAYso894EywzqtliJN2qJbB51FXJc5OAoZKBU8oluuP92/eTt1aX
7PURYbayGASQaZdk8HvrsByW/nVlZL6xTxbnIxrS3QTIkQ4m2AQpUFALVafPmOEEwlY9iXEGQIZ1
Thdn7lxGLlISRpbtHMksZElJ9Xh9y2f7aESeHWQEPI1kzHMZoII+VLa8YuvAoh4jycHIVhIB10xG
fcDVJo8hbk6swKVyDHkNqvKd7HX0AoV4tlqfV87lfEZ0aQuNOceanQUG17OzU6BuDyxHIWysq1eF
jBwGFQszN49ZAs8YE8u/LHv2lXDwhLTwWNp2K6s0qtOUutMi6u3U5P+N/zLWC9CkiOjsGq9sA+Ez
x0iKTbSq6+kerf/fyRjBb4e2+v5Vtabo1Z7DcDLb2PmfU7QZOenuctlPeg/tY9Mf8HCUKJF/4Cll
G7gvgV7V1CQOvAq5J3z3iD9k7NL8q55ad3E/NFQeyfcsRsId78sZYiAHyNAWd5KRoHbMExeNf0kl
VCkTAhJsVOTGP5K1o/BRtxJ5bYbH0kv/dfjl6csewcAatuYZA/7VdOg4RGB+VotzKMH4LcanJzZ+
v031agJ/FquVLNtwbiaPxmXERpur/vuryHnkiEkZ73ziLiGd1WGY2/MMM3WwSZzhUS7Tc9h7q7ty
XsZeidgtLdgcWPA3WU6Y0Lo3qnBWa9alLXC+NLqpcjRWAfuBryCJ05/uRNw5Gfw/4W0tGXBcEiAx
DyJmMQFsrkq2oalnUlPrVHh1e8Wrzrlmd1JAloZOfUaiBSSTWf5l1Lrr0pReM1EE2i7VimzUB0PZ
fvmg/0ZYGeMdhh6g9hMRO3uSOAgf5aLAntxcXT/m36e9ONW4EduErSKEH0JqpIIpcOcsH5RVb265
br3ZvhMQ5AfbDrGhr/dBtWCV7hRA3pPD4wKqx/I/ZzN6NCyqF8FssO4BZC3nHljhmozW1OgepW6i
oYRrUzL2Zj6Dh1NYcJKYzIassD5a0L9Z4GVOMZglkWC4bUCQ+AAaxp6sMjn3GXcgbqzhsXH0l2wS
WZ+dGod2lwMD5Yui33nqH/sTK70nuPCplTAFNbVKIGJmPM89rh5b7JzU3WSfqkqtLN0cXZ/2lEl3
W/pA9rSkob90qMTfk9dkvhZD6+UJS3FlbMhYN2b2Q7Axpa2oq9JzCLCEgkM3fsMcf9VI60d1a6E/
FB1i7LIrW9izR2+2rVMPPBFOtFpH0FYd5muU4Q16uf/K1KN11GQbyNcT+fhMI5hVrhIwM55bNEp5
arC7Jw43UzI53PrD2u9dT9EE62b7SVAR4rHoWTwFdTpYnYyCSOXi7RlSIQZE8LCuLZUfBndzWhsM
FeC327NgE1O8qFiDvsX1iHEhLXLyuC9nqMHNUS90oho7oee9SYSjjXGXyRZBjOpYNKLW3vLTJyNr
TNX/wzvadhDBXCs0j6Jjbc8CpXe2wsSywCnNsw99OQrVPI2Lozfh8Wj40rB7j+DnDw/OIkFBp8WL
Akwfmxxi+76Y+tWQpC6XvIA2nQGQZq4Ikl9irE2w3kvVipP9QUtfM+2mT+c9eQ317EaeMuKC07pG
wOTZpB04C6BRbhz2XB0qQQ8gK6kvybtARd2gZsd9HcVuOdHGM7wL+iE+vb+zd8adSAt/9Wj25EZE
7ERKMVeXSLoo5Kcp7OwjuG1kzop+fJ408xgZbKf31DA7TmBDJ+wfGmkYqTivOKq6aqnF37vTG0UI
auo2bksI1yrLh0QNkc46QRggZoiD75/Mfx1UuWRYmlMuUPg3m2FHXcAmskyoUSje+SyMhBJRQWdb
xU9u8sv1pBmOmiuG+UI3dPLzFmvAk/sMchV6y/knTynpM8gMFzSl+RcxQHNgex6GvfGhcKKWgQ0O
zepXl40AjU8aA7T10xOn478LUB4coNIP8eDp7KAytTDbXmg1a5uoUs+zdyscpz21SgPJ3l6OlQa+
D2VMDp1oQ4yJ6qnGuRHD6LBkxrYF5dOYiFa3CH7sLcOW+54UhR2yZCO66NLomnE5jZ8MWyBAyDTm
4P/l0mtZV0jZOHg1ZvVpWws0x3SZb/gjM/AYKFv3GcHjZQ3yvXD1sF8BEnU/pHgyeEoR4yW9Cb8I
7TaqjNDNJUTcBn8JG3mP1h2LHoMw7rkclSVBvApWnmGYTmIBOTSdfV24DTdlKze2vk2VqgGtxE0d
ETyXK6Vo3BcmNhlJc68yqc20k4+cQpAEZcLA9xJClHlN2ZYm09igfIRJjhqKV3gfde1pGZlm0Bzj
5SdkpEHbnU3iDdT0Q8NIjomMqrDMQXGbpG/hsodw9bkviYb74Su2EegBQSrinID8cNG2hL/40gSC
zIeUFdNjGsklWgD3y8GId3z8oONAq9ayDmXOOvVCb8KwqP1uDpz7kPpZT/w6YPSI6Hpp9DVKj3xB
9WkvgP/QupxpUaJvsoDAEUeS8ggX9T5STVMVQsyAbQHN9IpyQQQr4wImAK3/VSQjGY6OAoFRJFv+
lXCaNEkcAChjrSKUB5AylHScNiVA2NBKJtN6gkk5e09sgYYckxf0VuTfWWmIgcrTsnvYysGDW0/J
KRAbJdSKzXDRpwvO1SS3atTIOnQH/WGzn4Xzpk7gHwlI/YAO4DjNt2LGwz+dase5Fpuxto2WeIdY
0RlXgNYK5hgpefo44hao2eUnOtr0yyShWG/rym9Xd9sptJyRsB4f3oSac0VOQGiK2iCG9UfSnZ2B
qUfWQ8hYAzygVHT3/NVAtGQ/fhJbzInYRL/zE310l8DB4/viDWK2p1ym0VBvCqlpMpxyBqOJ1cBj
alLIhS/an5uIsrSD9z2wpOmI0GftIwzPkNmDOdr+nCA2K3HkZjo/gWM8XfC2xRkWc+mxm1yCizjk
8U8Ss7YQuiVD/Cs98zkwliewUNqXhSNZz5fDAs6UJkt5/v2NsKwNUxqx9+0F1y1UDedUwl+SEzM1
sZNlh3B+LRWlxMEBdck4QWgLkAUcJzqAeTSXnu6/Pp/jSuoZgEzwRwpOSluEUxn6AQhuJgc8J7TQ
+JMWWo1O8bDqQvhuZp0gZRLljEeV6vcQOlLby2n7+tspUwwTzKvnO5cO0JqCYjMmHemKOQsigjbk
iYCenwDIaQGvksAD0kqLgQ86ef2mmHuVtWjRYJKVv4UuUWpYwEdhLeyj7EeQHvJmeMBK4A3BErAZ
mwrSW1FIX8L40fWU5YPab7Va+N5AjrPgYdvng4vL4lCOYdNqsTQq1lfVwd5iXwmJvx/BID65/1Og
OeQOYbas0BiDdaQ/kTGUtbJisqbFaocICuLqZuk99eu83yS8MwmivPEQQwQenEFu4b3hFC+TtmEa
UZzvXG4GmMYo7jQ1InNjaz5n+j6QxJfTARDUoVZ6yjgIfGwKypUCViHQS3Dw2zO9nNY0WH6pQg+6
YxXOFT/Nys+d6gwbaB+uqvs/dFunfbwBgdz6SVY65unFX4eREhaLnRiIRixcQigETKroJMD3sNVD
8i/xk+0GWEDIbjem5uqQzkrpffDgl4N//bEGEbpOZmLgfHnAJI0U5PH24peWvYh9u6OYDwUjGFfj
8K3/PSePXnac0+jrdQPMyEo9pJrrETJTShId2brgWk/Dq0clk+XjeRse2g+eWyJOoNtB3dRxsFNb
8WLUTwNCiGF03XJPU3ELXm2luGj+dOdwBIC2NY6LnujjSXQVPHom51deTHtXtNZzlaSCwicQWftm
9waS8i4D2w2rPX2YSePYEbHKKvl33GonOvZ7Ag0stavRtuftS2r7NRXXWyXR4RocgH0LKJg/G3Jf
YQeVhQBIpGM8Qt5SQolOzRKCNEJcT4C4p/fwgvzjBPNR7yPLl3NTfgUZFogyt30JV4va00ma5R3y
Md+2Mc9xDHoF9x+bBbrItTHNZSF/SKNwkvKNrZJosKRZntY1VeJsagwdOaG+oVyS8fu17zx61drF
JKic/4YH0A/qrF32SZYkS3f0fYEoAWDnasVKkJyYx6STXiTCQ61lPwJvAEW810uh649r15hm+iBl
4C6+tGtnzuXeDdtnuSkEESBXtiyOvOAYdC6DjwVPQ01COXvuMAm+rVVitMeaoPfkDvf0UrRReYDu
i/O0WVAnopLURNRuftkgtlTYQU4vwcKsHRx+fn7FFEK++VYo10d4bXp0B6RqSoc59AakDQqxZ63Y
QvR3I7jA3lmfxZVc8H7kruXEBKiOCQygM3jkeoOzTr9Tk0mP7GLYYiaKOFLsCuCHvt6tigXbADSF
VcMp8McyoHTD5LdQjSQEJmg1rKnYE6D1v5h3OLbok2k2q5dyPVdVvOgsaN4bnSKUQMHA3raf+63O
v0f4a4Ij4LbU7zJDfsp28Xo5P8+8AX0B2zbfagXksBOGKeAqGRjjjVh7eoOtaAwbUVIAtBs3ObDv
Vhi0EuFs73u2rzJY9qxNHJzgXVEmC4aI4DNIPeN5UNo7PB5KP0DLurW7aIGfOTkj4VWg47xklLam
5geLkykBnvAIwgIEG7ZAlAL01Ju/jEG2j+chuiAZmxIXyT3aAhBU2gHm2ODcJ5aEnPOWfnAgmnf5
8md884WDORRUpjhjeXOQwGg/iMYG+cwW+zbYCEV5ndZ+ForlAQE/v4cCYfQE/xDKI4RyOKz6RAy2
xKisMKhQW91zDbpZuTu4zLbI9tryZ7Lp1464P2f5GcnAB42CF3PpinYqcRgP6JlJA9E43jQIK2Xl
sle28+Elf09R/Gsze1fa8CqWBs4S3DEtlQn/4jcTTfGMDGwYvcHHPbxaZMyXyLTnwMoRmhnb4m37
mKUXVrzPz+geI7DE8OhqX49pS3ZUELW3kehHHtg5JfAXiroMv5Au8bHDuMJDb0pHQUSoxH4ounTm
2ndV2NVnCTseMQ24dEBa0CIBLjXg+E9Qq5ptRdFE3NqOnoN86MuHSN9bcN8nT24mjjSwzGdrhQKg
qTTRMhXtMVy5+0VVMmXM6tQBoBRUYxEOnQj5SxzlzEwFDSUQ+b9GAOQW5uOBRC+pxVrT6dD0L58k
+Iy3CGt7ee/mrci1gJyBJBs0QpY991j/l5jQqcXPKnxa45357I23VFmtO/oQVl7mMCSgrtTBk56v
YDJF6yR+Fb2N3fB1WGUdEg6tmhtwgmn8gJyfFwcUNxbS/gEGTrtxEHmyFuBcb4RfO9hnVWhYBxKU
oeNKG/x6SGogKx2Mu41QQqSYn3dmBXKk0RsuEI18/10R7c67GCXF6k4EBuq4WUz3/BzzOIPN3LZk
zyS+iT4olGCFYU+TcY2AbyqkEVfva3902iUBHrfpeJoa1vw1QZrwdDDEpHLWJqHVM5AuehxCzhW3
5FSOz2GXOYmGUgetpMJ+2FV4yaixdE51djxWQJlxLJmYAfeGajWk78aBufxLIZqom8iS6ExppabH
0DlEbfZo6rYW7xXMXsFQt+7XQbeclGfRwYMP6/KdEs47TYn0gGnzru+GM7nAU7pNnE8J22nDeP9G
Zngb/XdLI2hQGyjQUMJxmiAhcqcoLYycVjgMmXHVdPCzeoy+cQNJkkZpeBiefFi3B/DFUKfSaa7M
+2J1pkSlzQjKq+x9omWD+8fCEfc9DdfZGyVSpQFonjlpUlqw/mYu7YAcIg7EOEAvZKdBnjlU6ya1
iAHy1Ya/5Y7Fq8vWlBzx4IIn9nGIclwVom7+c+z9iur3/WXSQxPS4yEXXqixhn6iPijW5CmAJh/L
eRQMVhczfMtDuGsjcnr9KzwuTFViZ9kCAYxdCazhPEf1q5ypS3rKWtnnwjiGso5H2Rte5ssAaMSO
H1z4hjAcygBCfUAnZiquYoF+jVHlClHexwGFUjKGfnv0bUYuor5Of7ZQb1X7QGgSGD5difTS2gER
xTB/r4+yUs6EdRQL/glz55+rYDLj9HCqBpx/2YNqjYOIh2yaQ71ul8hjXCGTCxbpAP670nBpYjyF
q5bCyyDoAK9mwkluB9HbFjIkZoLkIIWwmLeogfxzcvVvm9qjBvDgJs4eIjZGe300BkgQO6CkLJIC
ObeBNdWiyhJDihk/d1Od/0Zzf4C/x+Mx24OKdBDRPdZJeSOtkWwuBRrYNklkU65p/aK0+Vy4MfMn
D35A+TxIrCHe1PsWlaNsEUzOvhdzjwi5R1m3vWN564P5gfyYu9wNvN55382hJQARnBt3Sc0EnvqC
+pQzg5FfpffMNs4cfBRkEh49Wh9CvoCkSE99l3vqacTiLG0YnUFMFp6rsDRZQsUxMf+fsPB+ap9N
sEdm/vnURgJFDubEL4ANgKPwgZNbQ1M5uQi4boc5lucgGnBZTkvRvPbhIJo24xc+LtqWybxrdYAz
WjDRrSKuxRTzqAjyfoSoRDpmzooXbDyUXT3WX/FFzrxnGUv1K31G7AHJvjkwgis/L/c4wnRzm0FC
2lRrLnKbORKSCFn1QsNS/bT9SKT5B10eAZEJuuFf7YBnZ0+31engHnagfkPAm65Kx2xduzeK/7um
zbsB5bkoB/8tBAWlBOHeD9dCYDNAC2138WKq3pU57t5jKpMCGHXasKvtTEYIwYvYG2KbPkv7M/3f
dNjKbT/01PhnNV91eJWn+ITEhsJxJEFPh+LJ6558ElEP9QRuFEAcBtn6Z2o7gqEfMWAGjvaqqghC
fxozWGlXuc7EVYIUgy/vokUYzf0b2P2l+9nnG7oLBvLZmNisyQ74+1/SuY1xAvl34RxqhQxdw7ki
ziRv30qI8hzLNd4zehd51kAsPSYENkYWCg9TpNHOmCCZwctCHMo/hoQGVUk076RYCslKGrM9M3SI
5qCzPHpeENJg0gkdnC4YNHrn0sGStEPk5ofydfBaqrrBRO5sLRhDNEPD9tQJBvrHjiCw4ZbB4JRN
xhsWZB7aXg+IEShB6xdWqFqmm56q1VNNNKYft8SKkqgtkDi2g++ae7BXe8Zho9krM5rGVm96XCvO
QuYVpmiRNSADHuR7EYv+KJAMASRU5uhN+u+f9fw7EXI8QFjs/V+ew7nrVmBznJh3QDJ0ExihoDuA
ymBsh3QReL9NLo/ldU9wWNCf9StHlfBZe6NRjyplW4ifeFgzbG1sk1qzyuNYneaBoCrRZZ5pHHTY
jHPg5ggKGf7YeIgOZJtJpOVHdJGck0hgvRAfDLyHti64S3v+wD0QbQKdZW3SeArb9m1yBIQjj6Wp
fijDPJ6Y39fq1qd5HQUVEFMquUKHUcE+DKtblH+sU19gyNJK6jxLQxkvI7C9Qclk5Gz4uVluOgBG
stJ4SKccqcBxlofV5UaFqYqQNfWaBWTKhiQBTispAngiiLSlJNlrI6oqK80g8XCI8dGl3YADs7IV
0t6tpCqKKf3XtsCZWqAowyXyDf8nOqUd+/fwMZniSVzU5MoPxEcXF1CzJzumNnBDKqqz3vYyD/el
yGQRaruEjYccTxitVQjgF06lWczZSNi4n19ybB/A3vspOLtCNu+5YEvkbLwrVM50nW238m7sV2Qe
QOSeT5GDTOOwbJxUetRgA5tOsTYrL+SxbBKTGAIf3m25AtpsVOY4e8VZmbRl/So3hWyASlWys7YY
yqByujpgBRdg/qIvWxzXgl0ynCzhtQhZ2wPd/i27rgZhzYgV2wr7ruvcIb6bpMDaHBc3/4AJNPIS
Zs2SDmvvD/XXWIrxpaka9xKysODhx/Utx2o/nnxOL2YDDS5qEMcA9nHM7LqcDMTsDIWclu1Bgz5p
sNTpQWduE5P0dwYFtyTa36plm9G0fATxcSj21Z78f6iQFdGSnYsoWRTM6btJJZ/oAzYEzXTLSdIY
cyJ5JFKTPo4ejPZOhrduqx+j1s+QkXhDzZdlZYGk66OidORaa5Cvby6A8IVixUdESKMz7q15v8+x
IXSDP9AyYuUM4i9m6F2zV7ScavbR9VLuONFQR5uGDDB4segLu9giEHeuGG7wfNGF0TqndISCWpFA
8nPHO8BEJJWryhE60I6igUaL2oc2QnUXZzrchN4wTLECsky+Ib2RHvOG7ZaeizFwFJtJm1+vDrFm
e8KxEo+JVDMaZnzechE0o6vWzHKOwoLbs0v6x9NqmmFDS6QgKLPyCjkjKFJ6TFwHh0NNL7sUkr8x
IosMZAyHZBdZdINKWxlV9F9h6NXxKrCrHs2Zf3grFavjDR2CDNTvMB5BtkMHnbFKXyYNtie7MxXe
JHcWBYUca2eIzrUnz/xgiH5FmhvSF3Ap/PrjpIg57yIvwce0isl2TXUF9RWE2/yItflprN/G5Amp
mmGQgbZVx1fxY95x7PVfj+Ugf7w97IVrkCV35vALTl69HQQzJf0nDaVWAxXwfqmV3PEfe9Uwa17z
4lLuEGpMkZN48nVIDp/nOcGtkACdlYS3UHv5urZRzRzFbcNO02UeQVADOyrHFKRAHWrzqS1QjOdd
JPIprFU/SXkRhejy59zlQtKTmPrFHKZE9PqMq6rqj7e3wq4x9KlD+fcwkkM9UKY40bfqHTOrM01i
37eS4KNj2ZhNBP+eKqXnZucxARjGQ/sWfM7BsF3vge1/8w4LEULPDcUqsAzlduWqy5u3jCRbH4Wc
eq13V0rvAyHaB1ssbG9jtnfu1wXFCP4ejVd+quQic4ZCxRe1BWGNCmx+sk3p5wz4q7d4PBxf/5fy
G8vjcOcv2vUYOfk3N8W/ctn1z++ySiYRh0ueZwqw3DWDCaYPG6orYXPBKkQyTzMt7e2vHQUu1YAN
aog+MLN7aK2rKS16mGUUcYdWZkzC2ShmEzenKjJYavriplxrbYBhbF+uM78gy69++lKOj36HU/EX
C81f9jlYDmqbIyD0x3sdy8ypFgVKic8+2IHlu6gD3oVLDnuk9IJpzKKEzlKNGhwBJEnRPamwSJ43
v4ufZzLfS1YT+xrj/8aY0N1kVCdUHlGmSVDZncWJ5j/znJaNla84yK0iFSL12UZYGRubqbOgTzs2
G4NIpxLW6jmFxcerIvm7MF6OKRMUnbzodzIS3rJc/RRiriSKghBvOzLskRAlrSB6KC9Y6WJ2omJJ
sSgelRJa9tEANrxzmjfusTtAy/6zr9lCQoo4XSxqDyz6X+7b/8G0Z4P3I94L2aPRe7Pj/me9VMCz
euC09AgzueWN5V02AJK+PuR5g0oZBBoG4cBtK7bB3FIUdCIyQXZxa9G78E9v+6L9QmZd1dkbE1XY
wMHXu8vRlnzamO3Bi91r44cxXcjEkkyIpdZNSihWilkzALewUxRzd0KIfAkfPHrFW2TiIrZdQAJm
rztheTi9s0cOti3fuMs7DH2RWzDs6RVJJZ/43wONLeH2xKSHm8gkiXXpEbFXviEeWnaUhnWTi8dj
ZwY+FdehyTAMYJ6EsBaYCm/IgwAytqv81nUcV257uxxh+Wj46XS8JkuxGNXKjeqHO4JNfZ8X0kq8
G3jQeSNjyfJl+8gx4eaThX4VZMXUnbBRXWlWjgg+U8OeMGDoEA0PrTwvQlW2stLbqhIlBpQCKrsk
9ZheYPn8IAZl2qUR0SzHY7jpzoavGbIHJs32CEer7pQXGGe/32RRYOzqiaNNaVjau0dJpYeafXsm
t8TrrPs0q/i8vTUf2AcR2uZno7VlqzeGkokQQBxtpMij3ixs5ItuB4LC1bGCZxmfk8ceBSjuYNt5
Y0dIpfCv/r+uWfM8gSslVGwPhV+AtwyqSM97nl4inQ5PJJAn4kQQm1RP6KtOl9Yh2Tx52TSg78N0
Tayg0jEPgjE0DzKPyZbw7c0GuADjo9iwLzZceWlGg9xR2aPEM8iwtydAdKYe6ZazLAFQP+MaNwuT
t1xGRkRUIEnV6ff5FuHO6jsy67mdbivD8u6RGtQPdrWAJ/bPUt40tzvogxvTjjnWuwicRqDZPLUu
2+O2qzINFIlbVqCVyiwaADMIzcgNbY4Tx6RSEH1GYpjFRFjBiXL0Y5ib0dgs27vygvzi8ZV5x6A2
7fs5d2gSIWULce4HsBAyYBZ8jm2N2lTaaHxKqgMBdQ/wE++tbx/Z4D5wYQOnM045Lu8ABixi9YvD
aDUM2DQ+ne5CnN4C0b8gx/Z/1aBYKHL9Poxv9n+pdmzt6bkF+EK1JcQ0BHE7B3AqtLVcSApmvX6E
qCMT6yxk6inwrPyN490DyHKjdkPbDethMzsLbp+nTOKXylzZZvKnACsCQfwZ+5nVwwdjhyDs8rTk
5vgrldIiQkZNfiM75vaCKqFfvlLKOfA2LKcxndBk4/9m5RnoG7KtrmGeU+xdVsxIbDAOqz5E4Amc
3uEOFRxjuaZN1fXb5dPG+eoLNA0WH+mYU/6k7W1rD3rvhuvC7u0eSwAfNvVIPNrV11vMafmfziZm
YSSJ3ktrniiiTRHqIV7ljqi4jniyYbTDzu8hv1FItV99BXKQ/5b7UmkV1qDlAEbZGfqbZSN6keXt
7fSex73MPeZTZmIaUwsiqGawtIWAEiow7fi8Ga8f05l9JBr++x7SUOJsGyXDtk5xHwwAbhUQzGts
F+m9VyPytuWlhm87ygKPjjqxT+Zku3z7AGyMMuaymVuI937QhOdJxh0F/Mn6v+m75PERxZGjDsVQ
8H/WfvS7F116xu65ihiiNwoou2bnwHCx7d4XjXFdmKquMTRLsK57R4CGw5Qtk94CKDPcyOoTP5uW
hkTbfiZ3gH1JkKWIDN3bU/NWvYBXmhe9qlNZCjrkTSiiB/c3vzyy7AtdHrTzSD5VK7ECy7D6RG5h
ijo5UXuMx9F9CuuGxcc3Wl9j2Gq5+wkekTOBoEIfawtGa5pYBjdwXX83f9YEn0GA0j+/XhzOMama
gl/ZGFXifUopIaFSOajIkFgUGQiVmT/x77SLntpJp/BZWBXgsp6HWzLhQbM++UPvJ3eLcAKNmeRk
HuzJAeJXCZcKKKFI5JsEgeSRVZJGuHxeL0f2g41C0bD/aer8JC5yPwWiDq0anFgiJ93qiER/zgAH
khPaJaasw3R4jAFWc0fJZSqO5RoxPXy5z1LI1OD0OET1dvTbL61Se8pnEuFI8jiHfNNlt4pwQdRx
r6PuJeG+P1ABLGEksR58f0xOaeJ8lmPiabAxPEyHxCO7w+n4lPd9ZCwQ/wInX/42JuSbMJISJ9gB
4cTup+YiMG1n0CrmbFT/S5I7KKA8bwnyK9nt9ZUzhwlnhXxx2P36HHObAV3G7KhzZ+nB8EmJTyYF
HVRNGgKEH4RTCSS9I/r9bdZneqqy7hD8BTcdG108qkI+FNZTWBI5tgJ9bspGDFc4aXIR3RdddOzy
d8SsR70fm/cy31flUZZXMf5y0UZ8wAP2cm9kzFej04t05AOawxHzCAisDljzakYJPX9lEABLn5Yr
UZ4t9QYOOdd0XhKGZfsnn5OK6V9SzUGmxxXUeSKW0PfbMt/73XmWkrs9+LL7wlFSTmoW3llBq9q6
EqZDG34DpzSxSh9BUgxoJF2codz+hzACrLsVlJHbjMT+faArOafP3MUPlHTzSHLCEdx6GQulxqfK
2gMyUabtonYYm3H6EBPdRTnTjSL4iEVfv+7qD1i6/V04tNsp22blwNtKdjAwivLt81MNmInkLo7J
W1wuk8Cq1uHzbFU7lpyb2VqN6LD3qydlqc4W6wH7GfMyq36ITM1oLxxq5qh2H9Z52m8l5mjA9ei5
uvmqlwkAqT8NjtNCvPHEtv2x6tCtMJjmLfPTQrrtJ7dnYAf75UjZa6habrnnF77TNL0VlMjTcc21
NKqIZCbaciodJKIFcGtJ6CYRRnj07ix1ea2EcxKJcMxQxd5C/V3gBR4VxCSlTkmTw/GnMM8UHAjj
MZfnTyH2LdxA1KMtOMvt1+tZLfi+54m/ccr6YBa79vUhrx7EACiq+qyQax26IQpvSA2VUmWgqy8k
RrHFiHih6vTL401d6pBTcqwnipMcCXkr8ikYzchpv8JFPe5/Q74JhK98aidX7T360MILkf3NWPEC
CexPT03XAEfLzhmTZ5IuEtumHXfN0CVUpAXHCDxC5TUdRN//RFyc70duEwPO/fiSCswFwwaK5ucB
QB+Zc+tcHrSyq5mUmet8VCy/lM8Y74kmCrRxvD8Th2Bl3iS/fGzSjnt7+s7MXESEgSGrOfodxNLI
OSVgAJ8oCOM+kywOo1P9pUnhboJxXqdbde50qkQf7Gq6kpP3NVzFh2Ah7YU4foCstAd4EHVI1QFb
jwRmdQnozfIVp7rprXoJkMFKWtdZbfJvUHl+kAGi8ah02mdCIVsgNPounsjSip8kNxP/mF+TPBGN
QY7P2Hed73F3bM0QO4oWveOfd7QDomuX1NtXMVyyUVdw3HarfcAq03xoYXNZbAg3rBJpafymEyHh
lN2Unp91QJDKwkt617VEqfHnkK4QyBGzT//uqPPA1EnldPaVLoQZhFlJmzzIpT4gV9lXkbGLRt2l
tHsVMJ6qk7TCBrBQeJz6n3VrEK5v+gvnOiyCUxbHEwgg/FbqMnJzDLLcbXUGUy9TQ761dMVGLuCv
G45U1rga4l8Hnxpvnz5Zj+VzIk831jeW/WakK1YCdD0DqfkS2LlpRirDRhcheRTcmHkipXcOCm4f
GT1hD73Na4n+8plkWmv3WB5NaKhvo91oFx69IfattDLzC/21Q3IJrfzzZ7wYXz6geprSAI7yoNOA
k05WoLX+FJY+zk85f3PRceM8/UNAbdbHuZ0V1HbyZMNlvJA7Vn+FuqFhbamTLXX5tvaThxn43AxM
3EF/k1+mVexDCnBhyl7R6DxaqxhSfQCA8yvkInL72OjG30lXJqMCvFN2Gj15UzRXAG7ILGWnW3CY
7ipzpEQcGr5pybKIq1/Q1Vkby8XrKSmuikaeKuUMkVzeLOhKZvZYHgLhaMBf5CodqqvtMV3+WiJR
8RtP9VXAf1alo1dnMwjpnwgeBu8/SUcXbBCPv2PqaUHHGUibPk86+WC4CmQkUJyMq9AspnJCor7q
4Y5Ohi6JNvR/YSqy6osqEq+DVx2nWfpSWjFIJKoWfKYT4X1tEo5iOpNaEF45n0g+EXVvVt+b8AVO
A5SYSNeaSzPt0tR31dfyhFnXR4iWJrGmmZIrIWg4KW+5qg/KhoiDl4bgjYIoW8sgUhffWvS1iMGY
Zyq5po4kZf+LVrUjXymC+2BfUVEmHJFlPQcsdZsELQnY0L9oixSF65qWDqS7vIS4fooKtpnFzNuO
csLMepevaJbph1AIoZzwrbEpjyULxZzBInTyJvzLryv3ktkoXIqR1UZ0nWME7XmXmy8nKBDrtzYb
Ep+d7TNtJSjFnvjGORMLQA+KtXyJA7L81Xdulf1yVy6o7sP05CS/IPMt/eY/tznXrSkEdujgjBAM
XAHOuJvwyNCvrp0fV16aYojv44BbTbxGmAzM11jVn3LAuzMg23qolBVG4nqenZ/Y5bAWrw80wynG
J9R84iZNjXGyWCaLLMWyBpeDF63c9PuIKPB3QV2pBM1L0epCltIY+b+URYXBeNzr6OvfegrWXE3i
scNpHCqhUkVHl3JZebRH19Lc5yCO8sXeL2s2r5e6B0ofBdsdjMpCGzrCuq+5wp/D3Ii4xf9A8H8S
1izVYJSuQzth+5XYRs7aa/3HWOFNdEl6cCzd0nof6Ahyh3yj8CPNRTUsPDq+MBy4cy5FgdfrqZvs
mASVQivN7YB9Ez07jZTvzRmQwJl0J2DKadKCqcuCooEzcLGpkz6XOD0mJi0L62dGUtah8g8WGisi
BzmMj91+4q7qxFJJYHwflb+jv5bEd7nGNnhyripgPlvOy8OoXiTnl9szeCYJYjDe1inwX2R6OPOH
7ewFUZ+IqP7yZ6vb5Sk++8G+B8+HueyuQlsdJfmrbuwrxR8VAujRj/9DzrTYmARjXLAAolcQAGaV
3vWJv/pSuDYwao6uI7YxKuX+n2RhxWUn3WlgtXAb4PKouLYa/tzEhZ3j20Jq4k0g9OZpKObhvOs+
tx8EUtkdMY4LA2zFESNsz4qvLkPk7/4NVOG9zB2a1i/AQL9SGD5etVh1slxaRSh3yuMTJeFqbXBl
pCBUcar/ri4FeuArZaQPyIOMYPffKsZOj1piKx48yi3tw6WdTPHjAfiZjbeG5HzP2I5Y2y+CFwJv
KLXFh9pOGaL6p4Z/KO6dvIHT7SgZ1yTiYnhTXJPBB0PFkd4u+47O1PPOclkB4ruWIZt30SBicXdW
eimDOeCvXZe5JyhPYqXh7qGQFrqYKep/YC21VfI9LmeMvhD1GjSIqr551aDWCYwyeq4f4FLHN2iS
I/Ts8ZSZyJrF7s+wB04jz82utZXT4v1Bfos+S8pABBC+DpW/iPpl7ujoa0cnLr1RVOIQiPP+9hjO
mb1nEnftxdMW2UYKKln7uFlA2kUetVGY6Hy+RDL1NEzZ0JZ8nSs1nOedUNgq+bgDgW+urSR+IsUE
QzdVlVpBIcvHlIW5/beKusfzyA31+4xbI7ifxiVPF8znmszMQFnvuL0vobhKLpA4t7LSrk9VsIol
weKhdflyzop077gKiQrNLRD6tSZ3UtQfB6wmTtZNnFoN+ZDB0LLmkU5arT4XOjJ6n4+6FXQ/KHXB
XRwrpb/qmK5lKzz6RGM2g0gwwppHkKfZkWLYrQBv3s+wvKzdBLAmGrLV1/Z9vaPLBOHsSfxqp5mv
lHqfTdpqAXFHMWMIX2vx57DsOB4r/fjfWkhRPg283/zQ3yeG5Hef6BKUy706gwlPhNbe1tcdXNrQ
LxCW4egkN/vDN0B38jQ7cWvSYZrraQttkdAaPe1FqQ870kV2cSCumhOQryV59ZbXzdCd6zStMmBd
AB5ieI0xojWZMD6ylMC1QR8Zu5Wu96HY9/heeSpGzwzozvH0j04Zxsh6pxzmoMORg8rUIP2E+NAy
72uoPdi/zO5n/ujWlfAFZPZZLEUDG09ZicnotX/cgc1/q/78wgl9ugOWTfRvXJNvrfiE3D18WmXL
630y54491xwxq8UkCS/x7946zRw5jtaeaSZ7BtXP3Bw/Rkx5RF7fGjDFDS1sDUXKHFAuam6GkIUB
BJbksc3Jf8XYIom0ti8ocE5SucPsrwPCGpHtD8j1LG4Q4bHIo0v0Ow2qXZTss+UIgMhvZHlgpads
EEfiikQrnGU2i/IAPxIgMIvZtzdkyoSOZkmlx3XoGL1/pj6ep5xM0FGFiNbIdCkHs9T4Jx2cX6tr
HlOlgi/amLvZsXDgpjFuKPfXALqJeRrVFZnkEPrKGlNIV9VxOMZyEv/SqsOFhlhEvrY1f8bkkrzj
iB/brgzA+8aZHTu4yXN3OnXHgk5tZbKNJjbHaqCB3ScDPrXEwpl/Nil2XoZeK7pHUUyTFUyA6XDV
cQVB0ReJuAzAUM7DijWaU2FJ4TJle4txevcm3HEG7RRfLsyABWz+uFrp7ImcCmERUtzMFk7woTTv
YH8y22QfXHJIniJh+j+9yUHAxHfU08bZyue8bcCAGSBO/VEghn+Xm/6c5VdFMle4BsdWLFUuBkln
XcsF+dCY/OX6X/s/kEPZ7Yi+9i/ZpOuxCaigyVGi+u97NO19m4kv+9LQMEZRTV+gFLk+aZzKiPA+
rN5iEy7ginkocqECBz7hI6h1b8K7k1QuhL9h6B1K/qPmMTrGRvIvKzMya/XyT0HANGbK1bCu91Ic
EfQkHdnGQMSLPpRUjF/xwY4VQ0Hv5XXSrFTuVFSnk29f4D5Lp8fKPL9XwHnjKQVjT6tL80G9IRaL
26ImBg0qDOdHHUDg3i3wB0KoJAaRJN8/KP5ybeAVvaQTq3Z44X/JmyZPUPvA/9O6Buv7X9xh73ws
scPwZRoYL3ABHCydaDzLaEO0dv+rj0MLQBpEY+A84Oet6nTwsYz3YEs8tAfs5Zx3U5TKobFhC7BJ
f76fsCn8XpCAXA3RqztNfYGanq/VtjXuF4oh+oxG/xE6mOWj/GdI7jhYhP0vN6c7NA1R8TYQVwsq
KJU6cU6gUCxcHIvs+rn4ROB1rDDANr8T4/o7SnrHb0/U93xS4VFhFPJKBwSCXa6yeN7qgnHtNJgZ
6F6EZbcIYz+kO/aAZ+mQ61y54HycJ20AxraF2QajubbguxwnX6dX1BHhbOQgHtF4ZqwqGBOzQV7e
FMVCveg7CoEUWj2Vw9nbSAZnO9AsHH8sidMwR6GBoE6Rpg2+zVYi6tiblcFWfAbJCTYI79PaIzsI
QW3EDuRIvKpXM+9r/CA80SsYThWGYFI4UXGN2Apm+ognR/7AtDCCI+SOLs/9t73CeZEUzVIwcUnx
MAEAFpRouCdAoEEkCc1Tab9O9c5QNm0apCVCfwVEPPGLKhOxORvjKsW218JiGQB00K2PtFIQO+Od
xk5V2uGsfkMqSxF2ST/9R8v2fZS/tL7wymxD2BzPxGWQk+wb8K8DiRfkdAL0RUMBcy3vxTvGPgP8
wGdZ6IInOwHtmFaJmK/RCM2MmYx70jPhJ4NUyiS/S/Sv7i25lBHauSEVQwt1F5WBv+bONlqRpJJw
lsizTj1sGVCihKNC2uLssogHHfPEOX3JKRMxmMeTouuzuMTWKOL7Y5mp/NIKygys+80381ADnm9D
Zd+aR+2ecV/Zey5kWx5sKSNd+oYvNW492SXAqP/EkT7bOWkFVpS9G9j/POR7Tw1tNpGc4MIYRIU0
NYIbWpDer6ONlQBWjSw1GYnm+R7K12YBPooAJFuftjCydxq+yXY7OFKM/C03oaLO1vVeo1GmT3/R
r1UU3QtCi1c7OuLytwvTk/43nzj07y7D1gV9ur7pkg9CqKOJAquWpuhE5J0lDaJEpwc/xk4W2I+2
o3PM2NBGLIb0QNn1M3owI5PmcYvL5C41KapUqNxBp/Si/HgDS9MyXVtr29ckrHnv+D91N0up2bQI
38/boOaMRhwS/q7tDGY4is9R+6ZRQ8f8QjW1gd/LhuiSFG/TQ0YIx28/cVokm9v/p0bcN3u4Ihi0
qIyN8iOgdAFRMNERM5OY0kTttdoY6Sr615fpV8QihfS/iNkjBNqlai105NrPpRALXzBzAQyoAdp1
39j1eMCTDmysgk/eb0E4bYwoU6aFMHL6oXedGQdS2th8v18/MXnKwjCrv7dEoAo1m8wCO/1tJStd
GPUOhtn/fWlu+QP3RfSqh2MT2OG2CLQJnZe0dbCQHCLo2hqmr442xEblj5B8CXSfjSkMaom0D5ij
YDsCZA18fIyJN85K5N2Qx81oPVuMlhz0hu0aVwWUhooHmBHSv8tgTNh8rakg7NxszfTwWHwooxvM
Woy+5A+Z4WOBKNVeN7TBSnHmrFRn+QvycMiOtlXhPcoiRO66xfsE9elOke3XktIvvZqSfl0yNPKW
p3sXhVqzBwVBCgXXXgkPj7eySS74evBlh+rmL3YXV+HT0HZnXbK3jZq+g2tLJK4WpE316ZEAvKeb
ieMt5G2oyxvXJzridmJrMeSE/P0SJCq5Wr4oj25rsaxHbMrF9epkgfM0JWx+UEhJN/0/PXPqNpYF
DtCY/f8q0vvgXfzKSShF+Qu/7D27tvj0Cb/pkPtikV0HURmIYPKvIrBw+wEK7QeByj79JVUdl6eX
U6IElDS6oUBw8yLxn2S5OftRDJ27Fq85PaKdZNsBwyDFT+bv3w67dINf+TmLV4MwPi3Gn01qT/NB
dWcjgJtXpaX6152it5NQ8djLcF2sp39Tom66rvNqtu1wXZuUx8dATAR+EZIGURY31Xqud/l6Jp7u
jUD/KQgymEg9FKqq2uH2hQVLSK0LCuLfZNf6ULicmZe13SAZVtGQR5FpbZoRHYsgr2rIvT8xvH6x
x9Ka2ahRWnttMHIkkhQUQl8ywtAlN5CEWdrhIgbqPNjl7GiFjXWsMVOCl69xS54nkVSUwvATdn22
/e4shenZhXGgZzvF9/bWCQpoXhQLlSu8upBVqUjMV9r/IY1A8oCJDoury9FQL+fAXYKeYyYuDzJg
/4LMURv9i6fPQe1PBYQwQDMirkc7o0RkiruxKTNkVUyfisAte7UdLUUd/5lkRZpAZAoAz0AMDZrw
Z3x2Z4fY3a2PHwOQf6Sws4fdXyw6hNkgCST0T3AaPjJN6+VvXIKu+e+Gka3FO96VnacDtWwS4ORF
YvaiZ9CMUpoYPT9ZdPb8gvFdiGRBGd2phne4sWPHHEme/NMVT1ZR56wulyrVAKwr4WFtPdlqp+hD
LaWnW+2dku79jqLQVDzx1bptN++UKXjzNNTNyhOYEf8BGe3S3q/0wUEghBUWiJZrMmtRuUWw8yfF
hyJziQPCENMC7tCkcSk/mn9f6x3KcN1hhqmiM2iExSeXD9rTP+gxjlYrdaR0soI1TGOGIqKa3fXX
eYKSoEgwhPiSIH3rK7FMgTSWWUk0hZ3PfW5DTXmMwGO+RmC2IbdKnILkW4m2F3PLx5ReHsEX+Rnt
7jQ28RDBTTsSbaAA+p/3ySZ0mb146D5zuFc66MZfAHhvIF6m40jFxPbCE8B91kRuGJJH6XI0R6h1
Tmu/Ma+1ZYQREzbqUgXKexIMAHTs6+y2mlPOywI0rdltTr6YvbqPf1Ty5DcP0yvesJQaRTCM+hz9
ZZ3iDsrcOTDbaf+nQVDF+S7a/5VxVSa76A+4MrDbEZUlEQmcw4lSE5cIlCDfj2Gr0KJjIWdP4Kgg
dK4+3QDP2DGWhdn+1mrocmKUy5TdMUzCqdocdpLv1q1cCNOp8nerI44HYz7Q4D9Gsr7LgFxaRPiF
sp5Rje9LxlPH0rHz1U0KuI/qUAjaC4YO7faQt0J22W4SmemW8jLLe8C9bsv3wq4K0MgTKg+Q7GIL
lfmwEsbah43uXWSWmqLwNc/1UKWkcyn/nvhIzPNJjcgBt92CrrIcqmb6wpLLMadWFKdXagFoL1Jj
CqGanSdtqvi43iRypAQxppbVheBZdWjksTprhsf80WJiwULoiNW2ivjZ464KnISNemHeeZv9fzSK
Rrcg+kZFAS7bXYQ9RInTQhwPTXqb0OtvQPqT51WEYvlDUBT1uGfcZp8VqssRPExYhzRrSyFVSwuq
HTGqArpHrUC0XOUjtJx+tuJVb+h+yFzX+i8Mdo40PSGib3bGTOqgOHr3Ncz/+FhpXaDgJyNPH0kl
84ZlKwvnNOPc2hDPirm9gQPwmBfPmS6qSCeadE5fLywNMpMj7GriT27C6Ol0k8oIWjDnYukg+68w
aF0D1k+zcfQdNdtdsW0+bFjr8bRrHA/Cw1mmWzNBbbhZHkLBmpUFRtu9BQQg/JfszNrHhZD5SZ5V
GfqUkcyoQxyhkfe7T7Faah0/9o/0VCwfP9s3K2iUVLq435MfVVB0Ol3FriEyu/g+JXafzI1DKssD
JkPri7GwAzCzXAsh5/dWf0OggWRvhazMbhoapc0QGInykuTkyOOOn6J/LWsmg4wve6MJvlo0NYjj
AQ5qn/GtMJ6t/F5vjPdBQdO+ZfR6UC1RghJ7l/oMGXOLnspZccmQy3nIXlvhLqlO3mDOEL8iFRM2
m8tKItOreULD553bR8tYsnj6CAiJOtvqKS2dU6V1/+6KnNY3IMW0GYrhUsFcPe+lCSmANL7idEu3
6LlXD+ApP2KkX3fggMJopVGjKNepHIgbbfrctI6iaDUzbfs/3HuPVMJZzllrgZUxTB7i1Wn07DrH
aJuwoqX+ZL6J6TY8A5Byd4qzkMvHLYWOsuuFrt7qKpUrQqQ3m0zIU8/B9LfAfy17f2rZaZsvqpqK
9IK5Nm3Jxvbb14VrEyxFwsmOjr5BfP09aOWF3b/3+0WxH97gglYLIDz+nYM+I1joZegxuuduYFZn
WFLGknEiyaQe5LYwVWOMn97F+UChvofuSjuM8Yo4K4W2CLMUZ3slrHhpHzjiNjw/T3qWw6eT9eK5
hA3rWwxziUI2KputUGmwXcGv8qDeY+RX1oz4MCoIvJI2B4yD3h1VuejbrwIsrhFByM6FJ3vOzS4l
nfz/AvzlsMjPgFG73T0MVYmzwrhT1II708UUKQCuO+kXHW5YjfEgrgBYCyikF6WSJjpSJYIefJZr
ZQsniOh/E4zanX9b7p5BQ1KIfKZqbogjuUFZDFyMfaRyHL7FHEac1AI0Zb8560J2c7cJMEmHqnTO
9k9oCK/ao0/RJzZhOVbpePw5ONkiI6jeFAWrRvcVLatey/n1Fqt3LTZyamNCsmOr0UjHoXagKxvk
urqVGUwkSij646X0WalnpVSuGb1cp11zMMHVFLoEyHh0TWqxUxXpI+oEdM0kE+fDfzLhKFuDg3wm
QyX/1UEj6HnaWNlfhoP1l2dxdAK/zR6CQYsaJ8q2n/jPi9QNwaEeTgYzeoxPdes8uslFyHaPEEkI
sCCodjOh/RYq78uwkMRXWp4agpSlHyI4xkJt+DEWRt0B3QL41wLUl8BxBNYATq0q6Ln4adw0o5i7
75weEJDJGdYUhDODOhEUIO23T3Y2ejg5vlBGyO7/UvfxQMhAL3x3iRMva9WMLrKpl1uTdLjxJjS/
TtZPIcRJWg5oIJ4z/CnQ9mZwI1q3LI/QW6efYebOiqnRA4KgzX1ymYK3Wzy+MvBHr5mB7PLjMenE
r9vRaIn4SE2zkx9Jga4cMtGOpM/bRXe04SW4UIRTaSxiSKIHFmCqG/k2AVPssbdQnh0CSA4RJyXP
iUm0WBlPH9TeKik1+/GCgSsoXlSx0RkxJqGs1rMc1oht51Wscv/ICPWe57FtyQXqLoG6XRgYTpIT
S8pfvTPZIYySIsL+dYzmVB/NTz/nq3HzpAdT/YvA2AVXxYVYG4pcoQQiHUzUFm3hKp2NTf5EVVeX
ZzyO9A7WpywuGeNbecDzELsocNpgmwA6fbXFuytPJRFKTRv/NUxF9uUltC05jMooJps9KJ8y2ldZ
YfG68BS2QCRewhgNWm4VmAruVsipbESTtlBFXUGWQPwvFtvLkKFRCeGc2AtlEJCCxD5LIqedsCKq
VD5UwpzauP0xY6jgZIColz0uweH/jLLEVDqWO/Os97itO4S+2qs9HkDzUqdLRtPnYjHAEwgRfQn4
xQ3N+0pAgP2SIoxt9IYhviC/fHsVL3L1elH/VEEO+7MPNW5pMrOz3s5D7aajUUToVrSVlIYn9D3/
7z1nUUbht/v9/G8BOum5licLUGYbcELpYYK6InVwHc2NpQ27viPHTV4HSCTJnAUcprnBXFee/2tr
WkCG+obRFLZ8ug2NYeJ03od1jzDoe9FgkI+LVJnLcxkZnaA2DfVwFasYlJkwETqr5FB4aBkyus3v
G22Aa0QGfUAiXQyQOHlfxnBywxJ+uT47YHAz9csr4e3Fb+g8J6PvsIYR91J6kXnZBc4nl1QFjm9L
bNhhizCnwpQ5kuBHlqVAwOsPaRyRavc7Vdj39hOl+RXPpKXusyLIiC48Y9UD3v21W0RHGElSUAv/
9mRaFDAaCJAijzOAXbPts/WLDquTEhFR2I5bujyFOzCysWWehQkOv1TVL9Om7mYl4G9ogd9tmnok
g4tBOW7W/pwLBV9cnKbpTIjJDI4zDdVDXtlU2TT4QPua12MbT6q/CWG0oV3ZqdXjIAQ6lsFLNpaB
qGCqGYCVjoj6ZARiH+tbW6YZrBRqQsYVlmJc8s7KKToOE0Am6BzSeF4tqRqnj5stH2bQxrv7b7in
wha6f//dXs14LnUh86B6Rnz3fQp3NwCp604WZe9yA227+YACQJnArSaSzkVJNLDib4GM/O+9JNRn
KdwL2PoybuJXwheeaO5b3oXNF8EeRlWXmOEbI0UesWMiODDX4/tDhHzevTXyLB2p7AcRt4KClvGa
VDEio2scoXzLmTXFEv7f5eglNfHyIn6xPRCZI7yg7VuVEYgMLHnjVa9hJ4GgV3ELI2FVNK8quv+9
kHN9gcO1mr1zGzm9AKfI2hGmArSCYikFyF79rtKGSOq7h5dT8GZNqcl3omfoerjA1zxOkZZtBBxK
AVCnJKS265qRV/IfQuPkRCay4gHTUDEDx8ZI7w3WrwYs8comPtQfx+ugFoYYu4YUsjeb++Kls3YE
SGYYJ+ADYScboeSHPbHnEbGnjGNtwD7eSP+LmjV/rrW0u2TinEyYUTfBHpycEbWiCCudBLfkFfg3
FQeX0I+moAxYyKRS5eytlICET3xPGYuKHd0LWMffbo4UXAoEnD8iJ7jm6m9pTS7zfzKxCYUnpvQg
UYIxJhJNavhZjTc85mc6RWIabdCtGu15AxhnghNP/s178Hp3zXtSK5CYnTma3PcF0+wyjLBn6WXZ
4eRlGtlEaBWku7/BcsZV00p17IOg0VCVqRrNJn8tIkgXI2ceu3g77phorpvfcjGyTkOZTHXbLZKY
bKCbbQdha5j1K7MxCe48h+bWSZwxqFcNjosT+z1H28E8WyiN88nd8Q/7ZcKDtmG/6TzrRC+5P8cI
Px3ReVJJ+L3wyfERovXtMcS3q7e2XI1cEV4pq35CLv/1U3BxUFlx4S8wWiq8UUSesF6VMtyqekTg
Rolx75V/tIwGTElo05T8E83tJHgtix8P5X/kmXmnWq4rxeu6ldNNMFGk1Vn+8/A96fDO3045f6lx
9CQUP5YmdOiNjfSCA5f3VERl9tGckNGLgGKut3UBtLiXP6VEjcx+fvGZ0/7kooj09BMZ8ZxjYAUp
uv5aUA4wLdGeULmpq/T8TsjnoqVuc2e21ISIEnq+oHzkwpD8IJRV174k0bGlPbq7w1OeBbUFhuwu
EWO7kYKVE/a3FjaskKpCRAlPLo+zEKK+H3CZsNheI9PDf1vwLQQf/+fYSIEveQ641jQRUWYtIAtr
io2yJUbdwfa78UCSgC8lkLu+jntQLXBQjXtiDidM6LI2aXqxnxPZIs2A4ytOZPAxIJgXp2BOSr8E
ynLoiZ9Ixs0hVzac3QiNzkGpsTcLzdv0/yPML77NTSBmJG4U/dIW6CU7c/umUFnUqpwSlNBSO68m
NclauQ/bCG54gw/ly87mdm8tIF7Tv6gh75eKM5lC/FPOZ1ONt6SkwXtXvvTlJqb/IcH8Gejqle/i
KwB8lYIBQRzls9mnFwmKFJB2UnhXXdizRkYJ9EGsLSol6diPbtoXIhD/iSuR+FL7UVhEPsA7NAiW
CNxCMjZSkPcug5ZS1c399udz8ANeIKNAG2eFKJVlGG7gnPBukUGpoaoKt4ndcVczIBjF6fRSLM0h
oYqmlMBjsdLt88zu34m7w3zMRE5h8iQr0Zf4nBvgnb5ezqVCaCSG3F4HGFOca45RKucm7xv77FIC
ms5i74qZMsNJXe0T1NJqmSyN9K0wsjbAGcmpKX0kSkPR7Yc5pR781s6xx2GPuQsnrCyDaX8ND8LB
3Sx+IJlScs8UT2z8kIrqL9BJYPllcIpfwoNm0z3lwLRNaBd0D+jZeUDVDmQR0epWjIOVh+x+njhN
/c11QW9OC96vUejOUiTS692qIKOdnOjb1b37mLDghAlptxG/y9kBIZF+iAEy1VoHC8+527mG/pmY
I8KNO5IzseWrzYoH/5gLQATA4FinCv/kWxIsNG7RCJHTP8OVRs5TkVQDd1GS0Tg2fxn7Cl5o8bvh
u0BRxlkkOFwdYKe9izWSd4KHqGyxx+1WoyUkvdZjn3isAq+LMhREgjtm1vuhFF1j6H9X335E5Tf1
o7MKLDr0fo2Cb60is3lmlTxJ+sP2dsWTJ+uhKYLOWY47RAjUNZM75hEODRSBgaQkAZbR8DJtyGFo
ImTBwlo/ZRHhwvlGq6zmAHGc4GbJvJDVBdnPRcqqPA5Npk+KgY5Wi13J811tQN04im3L6u5xFVvP
wFIXcfc3RWtT+oXVPaKtl9sA6JOc5HSxjeWe4Dngqyh1yZ/3lBNmrGFBzmTBnlskQI1DcI3atY2o
Kz6iRBmfwOS6yDeg1EXlpAKvQvDwcfXDcKE7mz42xuaIkzp7VkW3NQ68KaCs/LxhGmraj5DilThP
wxZJ7WeA5I7A93EbRKQJNqCaCfanCXKkOfHkKU2xe7OPyqRt7EDwykfz3Ik4Xb9g0AlaWrKNQqb0
aC+VP6mLUKJFWzqb36Cv7hsc1nlP7mC0vjwYEXqoAeSsnK7KqxI6s9lLG7i95dk3cNDlRKwCItja
KmVXoAXp1T8OM+zuVTGHNKKS2K4f17ID9J+p5Ma5g1HEebNrWt3cH4xYRajO6HAHWOYYNiBK23kG
S/u8EoKJu2QFCb+Pol8KjOVFUxvuo/4omhJ8Z3k4zppxQt8s3qfKjeaG3N65nmrKxgbmu7Qk9U1L
gNNU3/rVFDyjoVg2u191UarI3L1deIntTdsRTLQbXB0xjAUZE0AKZgUyBPAtnialCmXyM3m0/RkX
g/bE+ZYxs9//ERQS1i2aJgHpB35FTgkg+StIR6FdHgD7XGfM1DB6nMZCPNNAij28NebjYQ+b11fE
ulba80+Lp8BNvmiSJn2TxQeK0KeOCUxV79VNSqVCNHME8W4Zy91uzfCEt+rElvCm0m0ekLTjG/zd
iYYxMli+5Gfr2jG3MzS5VhNS1EUOcYVxgjsvG1kU3GJIpyUTR+Hja81U1Dj6vqT8hltVGv+iZrRK
AOJQK8csaXy5tJVEMRRMRmhj07/a0ncqdB8ywQpIIEHa+zJATvo4qECyYfdHKe/9MHO8kFfm3KaJ
U3aA7gLH4mHWFf+xu3cawQ5w1zRlWhX1kgphZY9Ey/MryAC9Z3xDoOupW3MnLl1x+uJ+34YokhgI
+JGhKiYtEllyX0Jlt/PRQp6ML4Pm0I6FL1x0/+fHz0DX0DJqiJalCfj5AXxRzPDwVI/QKcDOQfTx
4r0U4A4H0GRNhnJKqb2ev/YNWGgCjL0xepcZ405I0oQ0dze5ygzzsxdzRqXIaD9ve6+7mTes1rsB
DGTIJ0Te23S8hi3PKFTjWlie6pRrSmrbaZOaYQKLFk3H6ssvRZEzyThDAXeI5df2yS8zIMVW+94c
5tlY3qm1hq9dP07Q6/2MjNWhQ7wwVN0rggWTsk3DKxfntYCSf/sLwv688rMQTwkELN/pwMbyzR3x
BjX37vQDNeFFoPAsYE6MB+aXIjWYiq9lMRrN+kCspxJm3zjgBjQT5R4uxmz6BORYoV/iLcXFHHbJ
66uYFoF5eSzsZnsN/ZoZhHYZKdguhTVSqaH6VSjjytiKT504UwOjdgrIi6yuVZvfX2E0GJ6yqf2P
rdZE0SzpN+59fl9qi8WSXFK1XEGqGFrrNyG2cTx5uGeSTeTFYgZgAjmnIANXXC16s40oK1EwJUSJ
h2AJQs8byERc1N65wv+sTBe6QX1R/CBL88VJI1E8vSpuSzA2TUfP84f8fSfKmg4jHKkTS0++y22U
sjMujpVVjGPok5+aj23VXjcq4Fv58LjfzS1FHITkHdhEtI1+MXEd/OqwRQF9YKtIraf3/E4Gu6k/
fIef5iyt8CJ2wMT/+IHFoPujOUaBpgWYFGPazOq5Y1UwHp/RY9dtw+jqoXM+uAeP2tNgfFw8WXXf
ttvKyMXM2qtIFvzpxTzdldDia8rT0c6KhooP9mHp9ftw9FRZTVPbWWoRtRbrX3nAAb2NCFMAmQKg
JlSNI7c4y/WVp/ExewBWp7V/r1cxx3pngPepRUc03jNJp6SLNoF+B47oFrwjTqZySbF6eS+bCpN9
3fgimPp1N0cohv44NwCF0+or2OGQtrN71dE+EPLi5m8oP/W4qJkp5+XK8WdjuroGgYpp4hGOfLk9
eegUwGrDCKifVTG9QkxTyUfOuRJNqorZLE4T274Nf6rhKTNki5HrYRBx9+vESrmgfqKTU+QQbr26
6jl+kr4gGT9PSkIS+NUzlrPLTzGzKpP/xGKbemWdCECirKYN3Qr0T0kD6g2iW8dZDZM8eQIQrTBy
nzulvez9SeG8rqNQJr5/v7xQwOQB2mF59FdD4ciTVErCfEE2uPa+cIQWEYl4pu12qVVPuRb69tg0
5ry2bCxQpDlFDkgjOQctaNfQudpJ5ADWdFHrTHHPJsq/zejI871EnV2ZwnrJMuNnv2iTIyCN3IzK
PTb8l5ohQtab+l6b1xcGNMTDJw/aY0/WB3TG1ATPXEX9dvps9fSJX4OZIY84Qq3tvtmmdga25JWA
WcgnPZHr3E7RyLR0rHUMBapymSWC92GLeya17flsD6rX53jcPb8frmDcYk00OdAjO3r9UDvY4g97
UfmuvEXIPajvJHIMWClODzdO/TXNLEnK3Tn6vOE40mhXArET7/49+wYgoxNam2C69u/qp4L0dOuQ
wLWk1yH18cUItiOZoLZNtBHh+/ugBoh0kZNEeXeyB8SDMda2wCM7fobR7x2eOa39u82SL5Btp49E
1azkzR5GTawdfjHFLbAUT5nBULvwZShvXS61G6bOStNeL8qgmfxKHOMAp8AhIzGn2cg+3tSot71s
dWC3TpehXeUM+YAQYQ2q8ifFa43ZHaMSGwID46vaHbq1GX8OvlXOAjkYhR+auHFwTgtgHrYjdG+w
33TQsE/YyUaO+93OU7bAL2YBTQM4fEBVakJCW/+SAX2QBDQ7Fz5tJhOUqrXZKhklA9zBr0HXsLmj
OlTChy4h2VaIPkF4qZ2JJRZBsbgW75I5Ve0Pn4g9MJXFqlE6dlqlKQEqQhV0h37UZWuCMrroSStf
U8k9sBlgmSmd255PbgCVAHZux0Ld77RoQ2x2q5LELJoBko2V5GLmkU0gqsg4ZjcNew6JGapcsD+I
O9K0mnkt+99BtK+3rhjeSQ86AOEo6ZmUr1V2FVAhcMmMNNFMUPolnh8JgGaVAo/Mata8BGdIl+gu
BVQtDq7Duu4FPD1LWEYeL5nhKzqh/y4r7B0bC56WtFpWh55BOJfS40OsRDsWcZ2SDf2GMiLuvbKA
/bUuUTQ2Z2v33xrPV6558dR9qKKzePHb8iQoWnlF/+sWNi9fuyvR2JHem6ecUtgumve7a/sfwpJ+
OQqbNs8yJMRjS1qiIzJIo4omGWs7TtwXN7gksFQhYZ4BMlefg+zvBa83g7YBlAUeabb0tnDe3Ebz
Ht9t6GWHRdsprfxW5pYRZPfJbpYsTklR799HPs9eN52iKWhIIOQ6Puo9Ww+3diF1e7ZXrXQu2j/x
lIZWCBjP5UpdB6AL9ZMlOA2h5SyGS5/QmjC/aQr1ZgSbjJwc1Hbryx14Ry6Em+RX+k8T9vNE92Eh
r4P6S9dmOABo3PEPaKqpIK+H0h5cUTqmZq2A2lK0lEBYE8Na1Qned66gxBMIkxn05GD5Cscwnjsl
wfjRJkJKxAfInX4qyhUdl2KvVpcb+FHbDSoIlTFA93k3/3ol3uo6enh5nS3qG43OmDyOWqpuIYhD
loLaaa7nN1OXZ16ea0Uo7mnpU8DSYw/smaEzorpqZXs+Z80d1hdDd8dP06R2padIp9zdUK74ngzu
F6Hoof4/38hzcdre6kdhV9IctD1ewGYXTuEeiHRqk2KkXdIzuH6pXb7OPOg74erpyDktMlgixhSL
ZVZqyxBOMhPOSBqtJmdd4zT+JoP6XTXlzYHAKGVSIPv98PSKdgipK4BC6xuQG2vFPmN6YrNfdM4q
fGVnEl3T1NCvUB36qyTaoYLNHX47d+0CyYb0mARS92aTf7qtrrkg1d3wkigoSv2/7zkUVyh6vOoy
qQZktoHpDOO/Fog7fdYu4FYL5QEYFp2WtmSug9A+QJSogkj8uB+Yr8DIcmL/PM/dgUyVdLRfKxGC
9sAIAf3EWie4dFHp3O2KKozt6XY3nsKADJoc6abLvYr7GADJOjAMagEgUC9EegtCig9MtlFfNwsP
OjGzg32MLurSDcPdtdj2V1rVVI+9H/C8hVkAVtTbVHNkhk6JncjOQxmlMuQIrY1F57LYXNO3x4AB
TM0iL2TfLLlxP4YWaM++zCe/38PCvrGkgcSRGUi++qgjkf8PH2dMBsgRbwITc3uom3QCiDAWljIP
nx2fc8DORxGq0GoikSyYUVUZVeLVSAsw9G2ZAl6uCCNsa0mXDXGZtwm1h6K1mdKoM2uHgErShGqh
jHtW2fdQxtE30ECXmmVSP1M/nggUuRDsPc7h6T7kk3uywucxnRCBYeWQggqxJAE+ICASYxEHd+yX
tgMKuU9/aqswfpOzhv6c3KuvLQoR/ImAT3g0SyKjtNZsa2qq+tcy/NhX2wDgI1bGJfQkCy1NY+Lt
+3qbYPOHYWn1tDv8jmZAByAqgVlrNMKHQTx1eVQaxNTkisP54IyRby+rnHXlKNh8dT42/T0+upI9
K7tgyM9qWtWaBiLiQLKNYmICa7sKpu+k7cTmsFKl0ucheRk7PmrC5NNBex+W60XxsTZKN/qJ6d+1
MvCBr9tkkK65YF9IaCX9RG9+qTkyxeDiaLZTD77gg9RU1LGlPmO3MbfSOj4WPn0DRYoCQvWb2jhN
OFa06BG4eZMbpsYOBGXiGYCM6b7d4xR8fxAaSWDPGy398/z/7rvgRMcWnpD4804nph0OKGJCvgFX
qP367fgRXkmZ/ssTfSt/sv9jGY+tz4q2wfXYTrhE8sVkxAZLlI2DhimTSJWOjFRAcBQZC2NKvfaP
b4ywbchEEE8NwJ+l2zQFQTMkh/0o5Mt1Ph1P2+t4G2K+O7pIUiXERnBHzyJSxkIHge4g6YDnIqaK
evNTZ4vaG5CMfndY4wJWUu63oWCT/BWg7X/mgXlxpQtV4EvVjNSVsw435TdX4gJHL5XzCwCO4P4h
M8anwVIsPtac93940N/R8wT25wEcG1DnTbh8CwRshNPhIwVA0v5STyqu7XVBkyhPlyYh3+UQS57n
o8bEgKeldhafclmz78PWdWEabBmv6poJIjUc7swYRmbSDFiBhURq+EJyKsbHWyeSKw+VvfzhSTiT
cJ/yQ5t0/MFmAX+cEFJ8v0/nDpkHcFgYFJBav4UFm093lQao3IdD35TXYPsBDNl0QQJpp2kiZOjT
Bz4w07V5Ik29c9cXiQXxXW836hY28dm1qEcBnXLbr2casvlQQ7DSYNXCy1XNY3cFk8wvPFIxau33
ShnFjsUEv5PHDe5Ox/2/7K3axKIhbhXnyqfm9a+kOa+pRRptTKChJQ6Jzd9CZL4/rrbRGynuiuUr
e9im+tii/XtgshxACcPdTi17fqh39eWEjPLudTj+xCCdY+b1LZ/HgBoAlLJBbEsNB/0eDvv0rp94
dksdtXdrnryv20YAXRYhHKKJ2ETAiny2C5t0HKKeCY6oCcj4epn3EfBWLHoS1edemurX7D4dwt3E
zMMJTZ9ailHefd5jlAMNtKoElh0ymHc8wDXIUSFq3LY3OQQSDftqS6oYVlQluszowKmdChiNThNs
kfsft9L9Q6lrW5apKOIXstus5cK2Il7mzRJEA5gqjtamm4HbMlWEYai7nDA3fSNDYcN36ODKpFtk
WtGiC7CAskOvqqopJ90+2uO32GEUbUoweMePdcnL8pWvV7ZHpP6Cuf1IDX9eOzHRiVc7WlZ3OR7D
n3k9ebgFLuqmsW7auD0hpkICu+RVtq74GmkOxqgLXt3jKobMiyzs9DS6Y1W296AkdEZbKzJdwVJG
NIBEJquITC8BfRMjPpYzooJbhk1qlyd2EMamyrYu1KyP7TB07tvzVgCgw9vomq0MBFYUT45tkDT8
HeXG8wT6gSOkqILbePUS7DOs2OAYiClMzB4DRmx53ww7vHzmlYTpHSJbPkKkHlrB1DYEKxT73HAm
UTnJ8YGsMM9AZQrBoR2hEnHJIBxIfa+HgrA1YzQbznZHQQThpY0uEQwNeZwd/pHRjrqDVEIP6p+R
f3OC6IKel//v1xrH/enLR3j/xYSYuJO56tnqIBJK2XLdXgd8WmpyhVlBsqNFmgIihABb4k3x9XC5
1Id7jPtHx99ARtShLcG8mrwPqVp9GG9tNcnqgk8qQqbco9XF4YZF8sHVC8mdrIAVw1CQzX7U15lf
cocdsPebkx6QamXUl+Xtm2LmxcNAEJi0MR6CUasTjC/fF248iCX2C+bHCY6pc5QXYHVR48HqPgnF
IkafzrmvzkvG6E/IUxjaPdr1HZx2/jxPR4kwHn6GdpPDd5qGJwk0PFHSi7Me7wn/mSl7gIwxrLdL
CkrUYRPPPJyIYCL2oeKD+6YF6NCjuta/tYgUrdGj9A7zc2zlxoY2F4U4CfixAUJ8P764H2h2x4kx
i17jNrQ525hhW38VCEjp28mMXpr6+WaA1kkrqUjrfmTgtyngUd0cY62n3kjenoS315PVfrO/kmbD
Q60mlMYkeT4gJC2VDtaJ4DEWHjr4d9//rR3OvWbV6yOwWq8oOujV5HJSwJX6XQSc+oCS0rCvvCxu
FicmqW2bCjVcwZmhGQ1Lq9VdIrbLMn5NS05tIYdsRz1q0vyQkWl2j0ze3pjzUJWcfaFTzb4Af87U
bWMudwlDsibJIZvn4jmQGr4hoeKIgnKbyXTxqsgXDDgqkgzqNTXwtBIgpVevDMuFejOK9fKIIWuV
ZfKVACb6XZ9QcMz5gSsx9oqSqL0pX+MFrn4deO8s7gwz3P4GspQUVL2e3NI1YGnsvU15SD6D4YvE
fXcfPURX2slRtli+wwUbAge+T6UyG6AOXbvor0JTmu4OgwtMQ0kvHYFLLaJujbEzVx70MHPwmhTT
65A7q/jTD2AIXKRkZmHG5rj7WKYGM7gcZAxLATl2ys0MVG6cW5plbQfVP0/uWmv/WaMRCi9n6tus
JKYT77+Ilngau1oZvYkCcduqkkhxNZ1/+ghl7XRNoUd6MxruLhcFCqeDioyLjXYEUsM6zlaNzMBs
4Pi4C690QSEb3X3twxTw2yVsVmgQLsHahMejS5E3Qub23UPDw7jw1RFsOQ7i4xqhBhSseinmCI//
GDoK3fkPlNN3FwtvaBQAqLNjCVB6MaxTM81jq7jUbw9Xyk2ms81P3stRVqw/SHbOGggBl810v2NF
qqLY4jZ0xp3CUNQmBFU+U9SBf4b+2v5gKmvU7qAULd0gH8mVRPX0tlfTJstbVfSxZ0EYVE2CcvrA
9r98SKGhXEmBuPSLxkt95tTqRmAeP5+F109JLYYnWA2O98MgFZ7zgEPy6+N0rRE3B2ejlYhehTAZ
THitF0MfeK8UK/tPHFBc9/HAIn7lzRQPXd9NChyjaaMRKwJcqFm4aYrhksnN9xZOSbkzXYtxNWse
OLRksmdr7uA+uFmQObxJrIViJ2FOnh4Sk64JBYrI6chtL8v58jDc38CXN+JxldC/03XBux0msVZQ
dUif/PrrjZuAsEGBAzzomD20GGIxmQg4tPhkArXdj+V5IyOh7gy8mZgDPnthwZhtyw2JC0AcUodx
ODA0IfbDkd1XmzyxdlC4sF5ycGpgUwz2C9KLIrEJ5fSGBVvhfRyYePCeJE7vF8pBr8e2Rr+brrT3
R4khR4fpVY8wb2F7XVwrRGhUeFFurQev89EnVDmACfs0rJ67CBULiNUvHHpFAZoNBKSUjc81gLQ+
w9x8Rds6F743yaiqZ5T3fo9A2deU2+/fgOCH3W3U8Bu+Kt8bJALL477NrNnOL6mSiG34D24XSUOZ
288NOb+tkuDIDY/dx9WmAJQIroNwYryEKk51s6zvzUJ70GYvq1Rt8hmZaX7XtnkuYLRaraWFtdwk
kUYVRvbFG89RAcgwpYOkFbbb+z+/MqsA1BL/w4ZyGF/eveZMeTKPxmLedPTzrfRS3PyQOVv1xkJq
bwrEI5lt1gLr+BQ602GDuwJqF8tvhsj+gfZuF+lqs3cdR8XP5DTQrqbUNV6lOuBZTwhxEmbS5QhV
LSBHnOAGXjzDb1j77KZWb5j6OZFw7hfq0H+4RdOfQg3kQtudRP6Q1NWunEu0yk9Imo/9Dv3MTJNQ
3cPjZu/dkB7oWDBwRE9Jr38dE4me+xgk4jXKna2jgChagteK0z7utmf7c1mM/ytoq0BP7NeakrjN
YBpOlsrVFM6riOBmXw765JU3p5YJETQSbJqrJpg7F4d1qUMF4LOczdr0UgcJQw+UJUD9Cmsp6+eJ
YRpWYWHOVbzTjyEiG99/Kexdl7wezOfcF6s2eCDkDofhyvOceVSQFdo1OrFdTPoxd8XB67vuyrrO
4M2Q7SJjLJsub5Akj9MyBEgRiXLQexePomrXcOGYlzORPtL3la7bI9WgOFd2T1uXDclvVPV7DZ0x
i2yXrKxmT7hqxPUkbCNNGN0uPZ3i/TpR7aNVo8op2acEu4+g5x1OHsZyyWdcVdFeIUK03xFOebbm
zf+gD4x4obUPsYMfIwYzueU5/0PbF7GLqSjBlu3x/YoxXg+a9dHKb+IUYGnhxpdE55UvwLais9Ag
kKMX8aXmh2V/HAbhgzy40BsDDgoLqtBMmqJIfrTFkUtZM5dLzpSYjm/WlgLhZn+BXabLlCuHctnD
jBTdDM8AhL8xquwnkBXt3tIC4DSCrgWOcXIVVArdOLZxzBNVruMAYx/8FST/8M5s548mk8dK8Oml
Ag1LeSEnlFuUNkYzU8h+4KTdqEBYI81LwDwNtqA8YLdz0kGnbIpqXw/D0c3M3nvaqi7T5SqPjoqK
VQGGtgRiMJ0tgJKkP+drQ0hI+tUYkbiJbhrZJvCO+y7FUmVZXiHYpMbvJz+KNOKbffs0jnPARIrp
7u3DJHf5on/O23CF3ihLsER+asZVpnh33FhJr9xyvJ5piYamC6QYntWXh2GeeoDMLkjtdwjK4zxP
sP3pXzJFoliGylCahmzZSc9n3BYwLUBw4YqW1AoKv9T/euhmecf+3r4jQ0pKyeWe/ILrXa7pwlPV
Ef5YgbIc93IkTcA8/ywPQTZMa30FxW0gVClVAcn1yioA2znJwir4BIptVc4iTGc+fW/lbRL6UEVI
Jgb3o09iTEeBbRjdpna2d3Vh2lqyV+/36uTU3V6jKbFC3pFvFNRxboqPoLwu4h7u+n9FTlJ0waYU
Ff2p1F1zMaF9I86+81M+VKPo2chCdJbtE9+RNSEF29Bzi729gf/JAYcpfw0w2vbls/QRX+dXXC9g
HP8HcXr6MMpuBLfITvVySbq/fkK6Mx6jisKACJW8+IdTkNcD/jZow9mimLmiyC5N+xY/LipO9B1l
1S3wbdoilQnMhhPWrgv3it5HxCBjOWdl3B4jtDu2M+ekt78+lW6GutAwwNptm5G1P8zTy08qR80G
tzFLTY6ysHhByY4tpm99NN5mY0AtpD0eXeHQVcffq7ldjCYBy3fXqFcD2AEqn1vDF3CVg/J8vyOj
vOO+y5x7Uq06b3ATjo5B9S687fGzTDoPovNj8sXOCFCbvHiLBi1uRLo+lBa/v8A+EQbZcCwVGPSi
hqYpIe3/xsM3+tzBdIaAhr4g+oBqxlgr0CnvIrk4cp2H7qpwQCGY1Nuv88bWBD9vDcsL17+s3Ch4
K6TnK2ks0NQjwh53wE/jXyiBqOvn8ryyy3XAXMAPTb8fFb4MiHwOIspRoGthKzrXDdg19Fb51hhS
+ILLtyl8jcXAU5ywtT0FyPVpwLLmJvQfqf/MOJV8uh6Vh5mK2nRfObh+HhwHxxjbQc4l6Bg5w5t/
szJMOGwMLmDPQnwb8F1+5MriH0BkPPc0OQwE9Qdmmo8CcPDA0ggiSIUqwY/qtiQYU29ma/xWXKqo
tHlB6EGpv2T2RYi+fqYwjgof7Pl57m0O6eGd8NBh/cvZgPwblkIfY4mmIbAlyts3/AZTK/ZcixrE
llcKFK8+JhPabXP7TsbBNOq6njJG1TFPdpcZPKmAyCyQC07VQS8KoTrpe1+WdJIUsMg5GrkVnudj
bA8UmfGTCOU9F5DvXHHl1gcKKvsiGAXM14jtm/rnVxT9bLpWpMnNIjWc1S4jon+coz7qhn04IMKn
mBU4ODpqOcKJjMLJ6ShdgWBLyaopZl7+VcF3YfHOpn0qLEaFRCMvmzamB90HSntCgtVKNEfa/KSp
d6w8i0k2+a/KqIcHKpLu/T09JfRN5lDtPQOt9zEnHFWXJQaP+gERF9g5GzzSgb7w8hVQstkRk3M7
6a5jULK0Zs/sjOlqqkw1k/JgmozZDdSuq/NEzPp5VizmCGP41tagDeyn2MvxI8KvOv9w1IUeafeb
mRjheezIgvru4IAl/RLsaYqul1+oDulNvxOU1LnF5TfYGEocq2kV/QUfqhgE/8VcyKyRqrM/xj7H
pYo80p0lDF+vKgHisxwL8lT/MKFN2v/cLK8793xLGKygoxis1KGupFjZ2WnDvWZAVi6jBxbah7Fl
VzSsGugjpFsIe2HkOWh+r+5Fmf4cwnLd/OmPbH+b6jdPRqD13Q5HgvpQWEYC6bcX1OQy5f7wrx6u
NhiRGV/eqHrHjoQhk3v4GwYe4FqdlgnO471O8Hx25QrfkDNXZwr5qPHFW6S7Kc/46M11b79CnyxA
IrwOpqJ90ZJtz6ZFfOyrQfyYjDGp4shLDWg5BlP9la0oYOeI1TKEWEoEazvxEbDAlkWSpldr+Qgi
A23mkgfsm/xev1zaKQDRIGma/EUSvgO75pob0rMfpHWNA2bbsOtyBCUCLB6LdvCMUdPENvCDggNP
sQPbpA0fIkPdw54Ryy8M35fjdSIKuEPgP6m1JhYvwUSZBRwb4a2Ix0BF2IHtGlsewLV/TmaX3iVW
YJyk5k2vOFDSJwaSTQHEsI54Rt3tGofsfat5DvIlvNPW1ABX7/6IGU/sIYSUmZ7GCuO6r3grin3L
KulLDMh1FfT8L2KpvaZAcKTCe8Zd/0JdOuNFMaE3UJd2j01Suk27utgcJcIP8wtsiNeFN2KbhH56
yNFFHk+qO9k1iQRg3KmeergC8L5f7bkYS9Z1LYfvPL+XXjQflAjZpNa2rQX/vAQrFwqLocQe7e2Y
kINiT8KyMWEIDcVKT/mnqzYNVybf3oOdf3N2gzYLY8+/XUvolRGjH2KmBQzzoYyuJbR0egGiTVgO
aAmfuVuKJ9ws3W0tOk5D0qaah2axaEajIYo+UuWwx6aPagXc22splt4KsxuKdyqfhhLbqntKjcEm
vN5H9iFRfS1yj+vjkv+hNAvOpW26QQRk7vdnnfjbDmg7ZscdTHgh7Mp7fz6bQOvIekNwzI4uHTYp
RUpmmcX8DIq/HeXXCole1fMS1Wqn/yseDaWamswqvSHDkUm5fOWMIttGO6AUeYvFPxsOjDHuL7Wr
eP1ajyeWJZmr7MlgDtBy05DiLyuVFQrvRKQT8Ia8oDJAR1wFrq3ncl0oxOBdJT9SeO48mY0xDgNy
vNb6/s26yyiD4WE2Isd2cgSadl2jefvhGd4SeHi0dNLD9PsdaXwVnlr4LEV5HhCXHnGPQuNGzGIj
cICDyI7eKFtF74/ScTc8pOCFYr2q0dfxJmkHvslphrsxZNMwW2UIr41fBBUB8c9bSVj08osy3gRB
J1b/O7g7VLJQVN7RQaDKu2dWfN2r2EV7f43EVhkn/OhGFmljACe+BPVX8ifWwzf74M0R17SmRDzH
KR7Iqhj1fSYiLd1AFuw8IxZD8iCHDibkILHPmB+1Ym72WK0jMDhslmetQO5ND3FiyNJDvhSoSbcq
P1R1uDNlc3hMhZEBy/DiY5OIh1p+41QtV15QSSNnbcBt5sqaVHHk90e6fOAq9xUObV1zUOFgbWuj
Z52/0HmHIrO6z71tSSBt1a8DmxiHxPbNoUSbaQPbU+Fl3zi486G07BQihuGziQeQMfhPJ4UKsFcm
H7la3tKlEAA8uQoeXO1uzbqqttvWGVkGXvvcXI+ETI3m14rCdrD2ezMUei7bRU6io+i0A5Ih7J8P
xLJOgDgRodZaFqq9S3CMhL20WzSsVjKHi/T5piBifgLK9epb0IfZteOKXaeVB51ovZWEh1yN8Cer
/EPAvv3RH+puJ68a9+jYA0uEqLi8vv76ksxFLuJVqnivu7+VSk7RrwEz6nzuPgMCgXgOjNjPUIRx
EThpM+j9E1sbA/VTCqTeHpdx4+Y4uHW0C0feMStzseTCtG+KCqz+qc6M7R2PgpKT0vtmY9k4GCbJ
hsEzffR+/yawbmcY/kNeKZ71CuCpV4DrVAJmwym2tEQKUBCaq63H1KWmcnsxZXSTdyOpJw5l4rkk
hizEVX5DTvw0YfWHdJjzgIvFBS3XCqA2/U9UQOkvvcOvhmFNNs6Ytj3zai/D1C19nXOGFXjJWSwa
NybuoxdZyrkAaOLE/GFTknW1vNyQQkMRS9sZ+Fnzea0FUZNflPpo07aShNTsa7CMEYXmCjjLMOK/
3Ta5AXmVRPVDQfYgKmtYO1/K2rRZ6FG2qBhfAGM72u6C/pLWsNOMpKoaNjfTV8UK9o4/znXsGeKc
z4DjB6a3b+/iALd4V1OyHrsoe3Y6kZbagYmW1ebSBKRnhv+LvscsFm8LEPuiKbUTLB0r8GdROoHs
nhPXP91fJ3yyha/qawu5Hhgmyd76qo0ciMblM9LuA7b54ZbFOXcNSQqXBxvLbCN28F1ZpDEtkZMK
gDA3UtjfeBnIA466ci2zIjWX2Mq2HGkQ/zpjsZwQ5+PzoJjfa7TLInNpylttSumB1hIhWfhK0C7/
kU4vozRcC1swvJctnlYBhQhxzNUHoDnTdEjw7pRqf5ytDK6R+8InLmI8gcituM+gdZDurQp1NV6Y
JNo4Aggf9KruLUDM3d51pC7IGDYtdkustAUw4n0UF0xhMUsmSDgOAiEAxuhUHusmRgQTWGgoifIu
Em8bqdRxCnqPmR/8UKi01wsdEOE7Xsn1Dfqw+VBLbS7tsAxVQIXxpO5PELpmTACxFPc36y8793HN
2/hdlrzUUPsSMfNCX2DajLpYrbSTWraBm5C6FltNlVPzyfmTL/3cOGV8gfmTAHi+GabNIvecGFC7
VJZ6S1wsTvawIeN2h4R+aQ5UUVdD1YU03/lMawRgJpEljGFQapK8iE1aSvatfq9D3XkHrk0eJUnq
EEjxwyYfUzYejFjqjDx7/WISGu2Udl0lg6bPfuBgixD0C3Z6aviPd/T8Se4ON6nOJw9vJWcbnMBC
tJvBf5/JuCD+cf67NS5bheHjk+/mRurz/0twkFP5U97hFj6HFJezkUSNFK5GVkkSO9VCnYJ68e4B
YUVkSEybn6f4W78HSsbzyUKI+1XkDH09/qWuX+dD0iXLHt+f3yO9k1dDVdv6xfrSMgAhEzwwJqSz
k5qRsygP77EkUjhIfTWYCIL6PQ9jmWZnpUkWlbtrQGFGLZUbJ9tZMQM851gMcsg8omOBCKEi9JiR
RrhzHeBRrTQY2+YiWmO1/oOrco36E8h3ewinvrFWNiWd48cRgYoLPcoXVfGSzp3jNu6PMhG/UfBc
fnSiZS0AQF28SSgauhpeveI3qVqI8qen7MDG5pkcvIWy8rJIsJu54N6ezibHTjZN73EgKQaNMA5n
HhQWhje3t1LKgY/vwnsky/4HBibF92hdh8gGsmxXsVyP+a/oOr5kflOUDxccEI4+qF0V/0woa0uT
Cp3TxTZRKAV4mb3W5HPZu2MzRzm/863tvtluyYw4e3CFqyS3SRj99pVbSOJ2IyRhjeEIdDxmy4R+
rANE3dJigRV70a5iZiJa4dm5AQ0l86mM2oVyh+ucIvLENpAm0eQ9RRa7+AkcDKOVfxGo6uBnUyNm
uYgHtV1fzuDjM2LId2xgbpF0CyLywApNuPwQFojaYwr2BK7kHkTZF3xbj6p/iLXUw1R3X/wDrULT
8Hc+DnGmtIDqIU/bB4dS+4gtKA89xUTMWZGjzmC6iq3YEsdThK7M2DAZDLcQ7svsZOZOQu53vyrq
pDxi6AKouaJeoVI1j01DOuMAeQu7OqvSAByJACqzImD1jA20p3JEgYj97laEEoaTgQK9Est1nOb9
dmS1FiHv9o+tj0tl+HfjvgemV5cyiBtBWXureka1x8HM0hwkujB37f7n1y89NnunAZ2xuo70vX4d
ZSGnllLVzUngq+JVFq9OwRmAYmQF6Ii/moY3XebK9yo6eidZbeRlx9+WfJoNuNzZMctqObLAu+tr
uWuJEsL3KJjKPznEB+4o9mj4AURwUExEs5TunPikY8DZmR7W2QIdpyQR3hPUd8wrFQvpOm0UhOHz
uhXOD5V3NqtNpsLp05IL0jAAIcf+YlYeA/Vt+AjmIrqiYxPsANnGTaemnRQU7xlehH4xt/9fHn36
Oh2muyFurkewTorsHB9PHYkWjce/IFNyjSNyxSOGJzDByjmaHBeAZK0ouNZ4PwU3BHyA6feNmUrb
oHXLOxyt/bfmdbHhUH+iRPvZtkhAyUfA0O2M/E86V5Y4HjmNRtTCCw8/vO4ARzx3QhyqPFHqYJV1
9uDkY5VgPAxbNgSoo2HUeo7wADcWExkEsYnrjvtAG7rxfSIef5aRPUlWuBzbFetDVCZa5afUCBJz
mY0zc1GMffjCNK9iLSTpSrXx0Up7NExwNZ9+8x91F9p0AC3LBvXWqLVP8q2UDTa3mRS4xtfgQWvw
1rhaPVKf9Rt5PdM6tm1EQ72TJtcyWdhRCD5VTX7JMdPKCMu1GHgP6bV7lDqLdMV/BAc+qRsHTaYw
Ohbyv5ynjmZ8ZAJiv1oXZ12yo8pPZTkj3n54xq/2S8+7CcevCZZ02X+iRt/rdvDK1MHjlkt+DnTD
fwlJ9WLcZMwRd4Ce8cahsEr6DJqz8HUvLBYfwUk5D5GyjxN3wKkOnUrlsxmza3fAIi8Z78daVCc1
8/egiUVQoaCjOgKnSU7wxoyxtqXfVXVfraTyfMWKBK9ipBgDT6fkpBCnl9AwWdeTE6KtkrZElCrj
dPPymD5ByK0VkgNykhi9rTri2CCauSSqvI9qtajJSwy0fEncL6VjA67hzHXmBKvsqWr438obwWli
RiPmgqRFThE02M4KOGdkRJUmNeqoHH+8y80XjUAxlodnuQx2iQ6znny4dfpFHOCkCx6d+vEqzPJX
fmHTGcddAyMcmDey0KWoxhibrotPQUqoqS1y9ke7YxHf6336qKDLsp5Qm2dnq9f408Uv1gkT4Mnc
8g3sdp3ChB+nZq2vVRPhcWU0IjBPXbqxHYOD71Gm+NGTisaQvoItFV6X90hPWSfbOAdoBaCvXfiN
kkBywzJCULefjEbtWlNAJ+h2Ghws1cescmXEpTbYujcBEbrHNgYUXXdQKE9p3EPD4px+BqbN4QYf
1uqh1rzqv321E1qguXzuzvtMzvC4pA7UxF8QkOOAOyVWl6M9/6NEdF6tUWt0dyDBxOZnsvXszmoa
qMauQh9dkEahYj3FHlCOR29fT7DDWNl2VQSKlMmJH64WMmRRsaezMVnoi7srXn3GGYsWcgyxLTmK
W1OhXXxd8BK5Fh00JIi95VfTvC853Kzm1DJI6+exd2r2fTsTSaHqvJE+HmWU/g0HbL3X442ROdrs
mDa4UyZunNnRafW4op8qJJWIgis3lGZtwtnW9RfhZDs3cE8MsomhImeAJuiUaZbzbIowV67cKzMn
e7eZNiNwq8YiFXVSyiYjls8p8h74RkZIBoUdD3J0Bmr2VEwwAUIieeoocmgYMn/gr/6o0zlz2t/7
8jWWNMlszDOPJHNPp10B+Rz/oSlyWWfbxdH8UlxznHj5EyZDy5ghPOU9ipyiwi9SP53DPhHDa8Eg
r62XvlVmSN1sYZFoPT8tqyyebvGX4yA7dw3l6GQ6qpJYkpMivaURPabP/iMqAbg5085bFxJDDELV
ZiMKXdcKsd0gn1X3hk5HF7tQ1QxvNFrXFeaGAcGpV+OlhUb3gkFLbLPbhium2bX2Uc9OdRK/fLqn
dmZzmkerouGb1CQa4gF5gagY8oAVjvaCHy32/v0bASSO0zmAG+eeXqtm0TDkqOEcazHSkkvtI8D9
iHTaehYxkCFVf40CJtgjzSsc1jacLiAP/1RrECnHZ3kFKrMFvCFlcaN3udqIbW8O6u1j/CSPt0zU
bzD8oBwPOqA/exwRvw30E/pX8eSR1I//DkWb/aoAbbHcrSuuJV03q7QOA3jK6s661aQ8sAWxh81k
4cnZJDpsvIAWemGdIJNdm8EXSOkns2DhNis8zutQx/n/7WQ7LuMdiqeLxs9Xv9kRY3UNO484vLy/
LrAOQS6txXAW5mbWQKkhOXoCogDSbtDh3vhnNBiY/k4eEJpLuDFyPTH341RBkGrpZJnZyjgyBT35
nWbAX74IbBjW5jcIQaOZ37xj+UvhcCW48z4Ty/IbbQ2FLDocevJ4++KNJMxgE0pAWaNkA6adt6+F
8gyLbACFpO8eTgriPL03mfSvXqXtuURsLPv30dIkeEBcBDYa0vGpk57sKfrXD0MdY5Dz6tALDUSm
7V9VGcXwcZpDdSmwkACMSvGTQGqgfkU+GKfMyIVpRo5Ewf9Kur+uYG/7wFxZU4v9KSi/YqlzhN5G
g1w/GzQEEaSXnX6MaCz+gRXll+wjwHDaueJX1rIMRijyHhci4xyMB0qjDsDivfzOrIBKFGXjMD0W
sB0H+W9rvmO61o7xcw+guvnx0p0cKVu+REcH3fQdN//vn5lecFXKHQSFvW12xyE8DUoXL3qUtIuA
m2V9BuwPP8E5PhGLRJV/fIWZpk2F/l+RwnwKa4tl9Kt/U/mbQYabGgC3t5zvhLLMD0D3p6yE6uFT
/vNul6ztjI+4tTOZBShoWQ8a4wAhNGsrrU5O4/GRCQzpkY4pI0vcs+94iCc3+jfr7/BhPN7hLnb3
Ahf8GhtItd1wDGDoPt5D64xP8eHgyqQUY9AG5l+9kaP8R+yoq5nJv/oFlS9Y5P8j9gk/D6xWOa3a
pOdsXK+I5Ilbo0kaIvnHtsz8lAcWG+J5gbF1w9tvXV6QDXC7HHwPkRQMrVFsQsCXXoKCWCxZe2hr
Md5oLJZ+CM8ZcYW4sl0jpBkkjpvH7T2tWFuag6+Rv4j7y+uQZKd1ZofPkkTTW9dFDaVPkektQTf0
WaW/+VmqLc7P1Vx6hHso850OAF2G/a4KGJC5MhcIcTz7JFe5Rosl5xkdQuYW0YmFX6G1USA6K9l6
1mUX76jeSggg1ibnoV9/jZCM8+gJfQ4WvjJzQQUDEkME/H+ZaXd+/jn9L9YHAgbxlHzXzpXc3g+4
w9Q6gzOtvSkEvF84A/+FouWSiQflC9hAg+yoEERRwNvjdqwR/8Ys/938t+ZInb6jqgI45HxmF/Oz
+GgP3IagoObVaTPPt4QGhESDeSvwxsjXdhUH2uwUGH+S5ryVD4gaqRm+PcfLT3bC5AFS99wJzjNh
p1VQ1XympT0cZ9EqHHDYZJ13Rqy8nZkWaX0c8hLGzNaxJ1xKQhV1lEs2C0weNzumb2oz3wTfOT5/
aRAllg67Qs1BcEs+THzCUM1sWQqPfmF3aiSd/zNKfAMvjuzJO/jiIHuGuZwBW2qpjL4XSgEW1jvE
xdXT4WetssgKyO+eo581iUy9JxXqkIPVWOC6V28GvGUyFWYf5vdXUEjp0EEOnGoTSQZHo7f7wxVI
4vATDiId04o7KFhBc0ph03DYuBPE4XaulUqjh5DA9aaeaV+XQ1dqQyF5GgT2NM5eRG5sWZ043e9H
UpTpeQ4ntLRcODkORAG938O7WsLkMiMR4EhF7pjwzlOspKa2ObRV1gkECcfKtnGdLYfZ+RZJk3pE
sJiNZ3Mv46rS4B7PtaiKWg5ILpxVxO9NLU6a07NF2V1bvXqnJ9zpLuzX3M58DeeAeub3jVp/h+F7
qR11z4INs//2RAXBQj/Ja1Ksbd/6DReRQlZKKKC8dgzyaQrZZ5FRuamHdmIBc0ddRggbMynLFB2/
YRUBumsAztq+CSDGp+vNhWCmQYY4w/KtifVfWRx6eyLynUwui1m66X5LF+iz5PrYwov2VQf55lbD
cc8nXmst0U+32qnlq+cefknEZzJ6TEt9qsAaPW7J4mLZFRjKBK5DiX3eaamlZAVWXf9yop+VSU6f
psUo/eclVcwOyf/eZk8UXc+8VOGXOwTlUvAzfMs1XGRHsAPfn7Htg81X3iNAVLRfS30BYE/iZ+Np
succmo+OvW9+BlbzVknE4uRtb8h5i3uBHPVoFoOX7HZqqcVND3KVZlY4PYloCKckAyWlQbH8OigB
exDewwBEwxWGKYBhGPe52GpHTiUkfY4MM3fzHgYHNKNXIOdD8jQn5t/JHyk5qNbd6cOl+0R7spBO
srzIPb6/17pOF9k6vwl2X+CDTtbnCmlUVqC/2mHVSzxrZY2uuTBqUOGB1cquFZFwZyFQrUfRWhu5
Bn8i3AfTVc1/3bCE/M6LU6Ua7IzQ5/qgBAvhWXo5Voe4BZ0KqQvZxXHtfAaG/zh+i7znek++ocaN
jX4dBTgXkc6UtsGljfvytXURwVGT0iKvkZFmJGmo8RpuXNZjjWDNLk2ps2ILRQk1R7REbMdqkhZM
sLete5YY7pY4bAbk1ZXVJiSlwyF2eftYv/9JMnBqKFYr4HPzKUsV4To2cYLTY6c+cKtnUtVXHCSV
hwXMWKLQWPN7NrX2pj80ybA5TkNPY39uhBRxLHtIyQlZZkcZAGqVvaFtvfwUke3E1kZrLwKHtOFK
9hLsWFe2IPa5nTzVL9bTHhdUK2CQn/w6GptnpiZT43Dn4V8f15eZZUPkNnu/0EzXO1pF1TWU5luN
bUqLHOV1aGapg/PSnSOgZCV74hC+gf4fw7zgF6x+YZ5bdXYJySKA9Ktc3AYLcX7+xny4rJGrluOf
mcOup5L0XzeJs0y5ASgT0R/nZ4Iq9rqHLg3aBDd8AYW3l9D9SHthMEvcxkWas1k+UkE3Mxl60dWK
ILT8p0MauI4Q+6Vt5tX5hPmK9RrJKbzYJzFFlmbUWlH7vhszUrO5D3Rxf96Byrb3/Ufx57dIQmfc
Vx/6+Ji+dipGV6WdNC3iH7QmlBX+1UHnbCkikV+WJxueIywYt0sylzfnVfbenuw0Os3z5zqxSdwu
2X5gwfpcnIC2LaRq52ZrQbyghkqkneKpEE/AjUHo5k/yAgrBZ0APXaT0DjZHMdkfL5ezPc0nEqp4
IaZSjSJBNdTV+ERRX1tK6G1gohbxDRvE5Aa1FFrlcc0MIOsxSd+tDavEu2d5IvoXilVsMmB7MVdW
J/pYhRNtYqrPrB5pcgfFHwLvSmZ0SL0WT9aDkzunDmyxsBgC2o4vY0qOYrGBipQBoMpjc4JBHFmX
2ND5ReNPtM8VcbsHfmwm+uFGPCoHq/hBeMtQp6JtKI26MR0fWdYf6u0HAmZQ+cfc7apevHyDv0b4
eVD5MCReSB7dF3Pl759S1rFYx/E/7EwMKuyq1pSJUOLSGsUUjlo9wTVExAqW5Mzy24vPUrfRZBF+
j2NWBxHNNi+yhLUGTF/SMhHihteuPCFM+7TbU2Q9RP1O3GWUozudMjxz97Es1tThf+WNtlyzlSrs
EbpyIm1f5BJoyaGKavHw5yi0Hx5RIfKyVqoIsYD3YEa4/VMTfzRUfCzajSxJXLwT0B7z6l2HHS+r
mfj+3vFz7QgvJvXo2LMBrkuygL4PMBeRIbaZDVVMLxeBoGexXBv1yVsr1ZB+p7vaD7vAKfmyN7i0
Ag6fPc1KoZMlCi+DXuCCFWKME44nhrkYCEqL98b2fvpFAu4JmKK+5zWKmbVM3A+WwfH/47L5ulXS
OiSS1z1zFXpzmgUVMq3pgKwvM/Z/YViqKSkJdWsI0UVc629k0B0+FeN2cTEZ2lDtWB/Y4STZbq6W
5lvvmdFYw7oZ0vj3tH5/xlHDdtUDYrlCCyUotID/Tc5cEj4vTsgjXWyQaCwHVexuIByaSkRtOViz
BMldD0wD84Ks81yEUg+avlo63eEV22XxeL1ygwbA99kA1/k8GwIq/dSqOH5T4Rmwy09d82sD24lg
8HU+UChtCmYj8mk/TR75F+IaENk/KYjGXw7xcp7abIr8RO4uYoA8iMVK0EokxLNAhM2x2CyVEDyc
7GQ/LtibNnDU/uWUMMQJTe7cDuXQoVJtZB94EXOupHm0vFvXOaIUk46GlPn3VJR1tJ/a7qYdhCI7
7QwU/Lkc2XHS5I5puYgGACNFuMNnUYcMo6kc/oZWh/sJ8RBtO2BdQ43QWDr38rJYRaMRZFkJEtpQ
YdZgY1a5LFvkFpV73cNEuYftGVvvGi97fuZ9HNmlVfyIFoSs5sSf+9Lk4pkD6Y7HX46+gDM0faVQ
2GngbkeaAi9lXfk/EykYxWlHPjy+nbZHdEpYVQzLtGldbhnuzcQK2i++GpmmOWiiNfvw9VwLiruY
bVuG3KcgDfEndvkpj6CLKuVm3Wf/1KjPSREJ5C9Zt5s1Pbq/RCPAIZEkWpj7LFVbMKjnyYvyE0Se
C7Ktillr+wlhAaAplD1pdEypNheBRTprqca8fW9JzH9GF1OTNlJX3gLRPu03KGI1c6OoLrpARELJ
k9r5f8f7Znb149GzBJWS2EkQPV3d5pDKsYaxMREaiac5xlLSzo1D9wFLc1NgKlb+8SdKTOAWGXoc
rFMVB/oZJfAxreAdxDDZJnwNVCiHPO12SzUiLPNtCG6rtMmU19OdovJTRgDcgWGWp0Y81ywFzKvx
GipvaWnoOEF1zxeuYrUIp26+l6OASCF21mNCdMyoS/iwNO6PxkxTQ1VPzDcAnGd2444vpuanTn0z
AVmvg0RrV1Betp+Q7jSXXLFl7w8vnICwTBKQGYb15ZKVnC+1vDGd4r6mu70/ECXUiSZPD/gVCqoy
pkdZ6JQaMMA+8e6Eg6JWVhczmoAe5QBtSqegMthBD6m7RNVR3lles63m9eYZNqjC/XZ38jGZNVG8
EQMELWoCatS7tqEwEe60kVMLrh9HWWxOviAURKUmvyYigg30tnueoth4JtHDQ0DnrWW1DaGjUth0
v/VKA6BANuaAEWuTQjQ4gXutXnAJBpIHsSehXSNPgzCMyg9S2dVOQHp5N8ViqMvhvqegcRzesZyT
F5g8AG1GdiFOdqTsp8WxKniTy0SNwr/UgYKpWj2hzLmsNhdRNmL3OFHqhT0VnUX/6w4fz50NhiSq
BiHX4RPICEjIYzkNQzrXE8MyQH5zdoewq8tGQT2Aa0kXUXTXK+zo37mgl5bGNRNhmW7thSg6tacB
emV/9BapqpAhuDzLLKVlTA7PpVSgWlNI/9QkQrJJGWqU8Z/LbqCFGeNfHo2011pM+XgMlBPZEFHq
vwjgUs0rvS/Dtm+MocVDlKUEPP1Z04xeLTrvju4Yalbo4v6qqFMYzYSu1RtrzWRW9a46qVsgcz6K
3O0Vtd8EIFBU0JR2T4CSyMuL47nOb4QDna5BQl9pPYTkbdpBCEdONL7rgyM0C5eo17bDcvrpQq+T
TXzc+mtCqsnu6VBv5eGQzTYBpKor8vqg7PWTTkNEgpQk6Bx8MTTv/Ngvx+5Cb+THfU/52DTY2l/d
QGFtX1/VNlija4f668EWdLHze5Cbu735Z5FFE4k87Fdtb1hDu56uAcMf1vXvQHb9mWDJBjqeT6FB
2mYEpyKCTVsoG+p7BrZRX3B5Juql9ItBHR1LOwYt3G9f64p4q8/CcXjMQFiY/RCyEVh7JnlQpAUN
KfLGSOSEcr7yGeFfCmrmQBUW+gRQteIgwJzhiJXEN4lqyj9NOnOwMwxAqQUj2j/mmY4IPVKCrw7e
XDC43TNR5ZhrZms9cDd9M56lDaqy6OBF16siH/1e8I3PcQ4MpVYoqvXxD/+v81QXvhkxKOB7MoGY
0Lz7zuRY1ZxxvGNFijV0w/FyduaHbgdOTGVW9pGy6lf5hxdqmbOQdWjddbd1Ih6WyptiQagHVECh
RkY924dH4VHbp/nbrQiHsHoslQN8s9vpeIN2akcsMLTrkvmBMwDTtjdtWDNXWDWS/JzQiHTNryB9
PNfYk4C0beEP0tYERRnJn1LVzKQLjB044lf0VMADIojjNLOhDYwMsxtrzI+V5O+XDgwC8+AqqPt0
08LH7KMD4Cm2snvYMFhaf5P63R8fS+5zpSjT1QW8xSy3IIwPXutSNlsKJ+ig2UE8llrKPoQWlj2L
j4Hwr9+pl5CSjnX8xNsmaJX9hkhY7NF/lx0gnvpgtNxSK9zlfm920FHv1U/+Qw+V1Uadm4LrXdWb
6IAFl8MjIF2Q1lnvNJKYllDZXh4KFIUBnv35l8sOl0cYOenqfiyLUdRRDGr1Od0OijenY86xX+7B
BABrm8tVmIm7yJyW66UYRaVZombwg8b6kRsZktJ++3y+Dv2I0xpJaNxcahVoHN2qNvmpvFr64/49
44Qa3QJbE002kn3BbmjdJza2Cx/Z5t7XkkxwCo0SOtVCKQvZBIEwmcMCdpdbrdwP9xdNh+IHvcf0
G8DUW4Qi6Enoea8dEurSp3DUeNIrxQEGgoC0g9xsyCj6DprFxmQIQSizkm697ldTsVu9c1pDZ/Wq
Mu/Qx04abEFskh40zyxk157CwwwglkZHu6v0dXOUYl13pR6ZDBEmLyInBafENix4GtkKR0IdLfkN
GdHywpPvvgA50YCtdEmiK8MaGwEr5j7UJS+ggbxukV2uR9+1SVo9eM7Ux6Q0qsDctgaY2X3d/XFC
SoRlhrH3KMm3Mm1aLHWtbZSXpYIPLuztT2UBAZidEvBI9O61Jk3ggYGc+QQRzbrK5m1mgyCXsQ+p
V9b4+rxWaOj/UxnSyZT3spI/wTPYcBuw0xCP3rj7HclqKOmwXL/MMoV1N0RxZnfrxjjVd1+Vr9dW
GBru2gFZ81QsevPbi3+6Fq6KgM6zrCm7pl8G3qFPgeeThOMzHbWtOeNP+r9bUJVn3r+QgF+mgAcm
eTUuj3wmrXkyX87mJz5P7LR7jWXvzWnWfAfFWZn8SBv1PfFczy80Ja5i4XOtmF/U8VCQSC1fyy2n
uyEPfUINBueLjzvcHx2my/8E0O1ImC0DNemN/t5A18flZvl7/QYXiWo6d+r8ZIaigGH5/yTpvmmv
4l5QAx9zRAlnFBnaDUx+oyC7+KNNkH0BwfLNJ9Mw3KiR9p77Y3oNISWxtZkmucjSMEwZQKaFNquE
4Z7eA5HssUL8VWmWBRMeNZJL7k0+/7ocsvlQN6mCn2de3JkHO/BFhYkr5saJ0eQkD02q9bi/FFOm
j2k7J5SpXpNPSo9VNDVTBpSDbQ+gOSYXsm9ga7mZN0/20X8NCiAHKPgYGItGyQrOQNoVZY8Mwx2r
aDJuGGJKymuG1FMVSiwWXkOEo3cwY74bs92KBsDCYRM3C2KfXI8h6bsQiyX9I5pP+2iSpVeeWs8V
auxRZjuLKfEDWd5B5q3T9D7XgOf16nvRJRI0V5UWZyM8/RY0zAnmsbagFnt0LqlCWKzbJBb3aPqe
R6Inobx64FrYmcobF2FlcqgAnvYSJGXTFzS86mHXbTVPLvHlcGaUHCB7cbrxYfNitpY7jfiNS09e
YHqpqFZCT0YHVkqC0iaDiFORhGJs4wt9R5SPbJK6x8FgxtxofLTd3VhB/HsiOSimVyXv4FovjjEg
8VP8OeLiYa5nNyq8ZHhJt+ubivfwZ2o+7/Ejz3CXXE2aw/RPirbcjfkxE5jriaJzx+aDSQTNCkaB
fPMGxgywSFc/YB3tRK1smAceVBl4S4gPW6D37Z5ZyC6DiY/F8K/4lsE3A2npP9munX2GhEaB+8BX
A1mT2J+g7AWROJ4mH3ZgWTut0fNGF2xWDt4zUXBDXqYO9Sxm/EOhS+n8jge5eLs03b22vn/bsN1N
EmVdz+Uf3AeYixQcERGy9bEaEQJmMTczWfEQMO6G558pfnF60ePwoUovujW1v1h/yUzzekDDhbq5
aVbKnN01899faDjDvzWthj0KyMytg8tfxJEt/PvcLFz0ZnLxpi8olVFZwqblHcp5v+4oehFMfjWn
iCzXR+V+zUJ7YHZIlQyrBAv8EGwWWnkdpD7hZOMZC3p08cDM8HXEiETgtJBtulVt/lL1KxabclRY
T7EULUa4FkmrdWl6tMxoufv3UhjVp7liQLSy0jksQV36L5GqkMqvrMx7aHp9GHz6U8DNr6V2izU0
NuWd+gnHCKP7T/k/1N6pwmgBWAu081OZv1p3zVbWL11kSWt5o5ZF6tkPQzw+fawvctHXtdha/sAp
u2ZhPgY9bbR6jOBiLQSqm7wsZn+XvPf6dhXc1+jArV+mJhNFEQ9ie2StSHNXj/5/4BWWjiiAtfsM
QzPeQXUnIYtGAJpGE+bxdBUGLBaA+rDs7Xf85oOX3b7QCXJBtsJsX3oFL/JqZ86LYXiJIiuESY+y
eMRt0g9E0x0rBdEiHoEeG4KFNNV0OdqWN22qrF1A5a/82gCwNfmRojy+9ucsOjHQ1X9rcUMVfOYd
H3kG3uaxQV6PmW4V+o+1gbxJMIpxpv4qzzZT9YN7vcs1a/2xBNeHhbx7VFY2BUoRTTf7n/E7irDn
txdACIVnNVA3a+cI7idqkkVeNn98wl1Blplfqt9+9dM4K9LjsS/UYMvTh27zF5YDEgjNBiSsDgW2
5mNO/A+pHncvWH5DF4DxuN88JEIOFYyWO+SX+wTu/W3dx07hRsmtA+Uh/8kEyj1w9YArlkZ/y/R4
n8D6V6Qz8TKmyZfG30mxWV+44cuzMJf3v8SpP8d0e82bTBoWq6Z1fc7Sh85AlaZbZT7S6hMHzOat
IVDML+NVMCDVsKk/ivkAtJtA0W+ceUjERNyE0HhiUAvl6v3qvaHE9Iw+vUO1AlB7gsh+hxM5Il4v
imqBhSceHD9q501yg4XEBNONJ6uRdVFxkrZnU2egQ0NftLScGnfzSms89AiqyyC/WNyte+/q5iWi
vkrDtr9ghsG6zMYzgMDF3cwlxzncJ6xIbFIP63YKdRlru/mctGvOEpyoxk2IHKrdaZE5xOeVaw1f
rGThDyEO4GDkV2JudC9Oh8lukLPAKK4WaIEHnf45PZqIQJbB50vhetVtSKTWfg8mk30KJ13uca10
xrVsj0bZxkjJt6Ax4ktfcpjOiPcf00OZ3/V2HaQ4Xv/81YCy7kegymCiAnJqNAofL+ehtFbgO0i+
lYZrxBtXldeCWnjheh1U0Q/Wo8dz0KEC5fsDqH5XSAodir+qXzgVX4aJMa1anh//+S+FasVtMkOw
ctVG2LvYxo50EiAt2SLl13rKgPo+t3DTHR5zQ4lBgsFl9eW6jmCIWFAfuih/74aAasYVEfk8OiQd
nz1Nkdz9Q4grkiVZtnigmjlEteG454fYja4zMr/XBFZ+/TOKRKhphoGNUFqzyVDIZUWtjwXaLHR7
QjG2kQbnPqGdnBMqRmlMTJQVVDWSVIUpP3Z46UxnKeBYze+AojMav7aI2asuSALmw8Ft0dBz4ucb
THTe9/nrxlczhHMzXXcD59/keK6NPMiZUyEc2eLU2bZAkturzhs6RnNCr+tVkDH+3KrnjsNxRt0y
H2I61Se382UD7b5AuYHPNUTaqUPLEvEA7aR7egzlO0k+Lw61vhuVWV9BkDnK+ZGVQWdEiHwWnELr
vmroSrwCmpm+RYssQE00H2jLHUyYxHIC9IEHeZbi2Y0QrN2D/31mr98cH/77sEZk8QOotNkuVWTD
d7fVWVa56cXGujTjiEKTwiICjaGx2q4rutFMBaYCNSEFELWIUmeSSxznrIdOpVZZEExQ9v7bD3Ef
nbTJvreZpC5UsaWBRZ6wTeuwX5wMrHlto9lnkflK4xO6m4ySCnWybez+KjQf3bgwuYlwNA5RPj2J
EoyVt65TXw8PLvwFoWE3YpKAGiFLNq3o92xw4mCaG89gZXzJupiFV5d0lWf+B4RQi7btIQor6MEf
rlDcoYWNE5UekyoVLYassttsRYmTpCLAp5wEb5MDc/AkjZn7j2+gOGHKpRjjFDfRU6h0HQIdTylA
nrhoRhomPVl9oST27QamawQAwdQlfCTEO0igYeo30P5V5yQ09dqsF7LNDCYDe0uXXxE1QulYRCHu
l09uFkoUwQW9dWmsT3YGBiix/Ftc2OsbiFISXRxjDaHzlDRn1vJxra0G4d+fq2Ui8ByVzU9wfByx
W2HZhPyj+n8ZBlSfwhqusDzzgE7uS73rdPqiySiU7EZ6Pru4nf5dfLTxpXqbHpyAtJx5ok/10LJR
rqm4NJLI4GBPl7qOmWAjSw+rWhG5msLxsbG9xbOft2igLe8+lFUV3H73oaY+67tR0G9AKTu0qhKK
UDQtZ3mw2IbMJ3aQxxqY90EIXCNxZWy2o8MAAqtSYBHh9vdOJeQ/9an29fTew+xoH5HYARJQKyyw
e7WVmbDZmOrwnRtzePrvANOBDOUraiGHFE3UpaWhhpL5eyFbx61frgTuVsUhniu+4b3rgLPL7q48
kRJl/bAXJsEoiSzFuXfV+it3HeV1HQu/GyK3Tu14sxV46YpGwuKBBHH9h1F+dpN4EFpPTo4w9MKf
r2naGM6aXcjCp8sc9sMYafltYmSosYR2IAwpNcIUnSqEp5ElUhR4K3u+gUDnnZy6qe03jNHzUoxG
J/O8h7Kil0WvMO1NEA+B5UcBo3477Jv6uGpdknSlDZeXf1kQyf6CjKPosF1MrZOjdlw7VDTCtOLA
oL9l6lkrGe0xCXDp8aKhWP17p5zTFpm3EkzO2mT1Dz/FbialRIl2Y81OA/j35plGb4ib4ycSV14/
RvCrhVfCbobV6Ox+SKrOUB6+srqMhr/XXoKKbN++acNJC3ulJ49YqnnBgveSNSpze+y62BI4+Kmx
VPBfrqC8MujIWZQO5IAlJZ1z+T0+9chn2UvoI7JwVc+2ZzWo6RwhynoubGBVuRE5leT+anF/bPJD
nn/9ktz+gcu/sj0ieM3TdLz557BNBQGOUTCIUI0togS+n37k7BDZy9jDn6T2Ka6UH6NPP9RDnztU
IEgtlF2IWAMsCBK7pqo2ah9okX1CTuQ8WdquhcexMT+5btCX6bFqe9f/7rsOY0nwG1A6lwbkrc6o
1U2Jj8mkM5y5i/o651/5a8WFIhUbFcpXBCQRudkO9nHr6W62Wlrm5lAiLS35Zzvmw2Z5czjM55VR
qMwrcfbfljjVPUFch+m1wWY3fKALqJa3zyL7+LbmWWC2n1EooOucsmbTbXWzmEgFBsnEwqVT71mX
3SjO40bgMEsqKLw/3ASJgzmXPrXp41M/n/zAvbsqod1ivCgHXBPRKDNcSBbMrs0PdZ5Efpf3kOxD
3jUr0hsqWaLOSRfLMTrRsPvmB1Qpm7s0AVUG89uNUmRgfACMWtutcbO7v/01v6+vc5dZ9ayOPhjd
Y6RC1GKjiVJFrYk1EMWZTXxGgsI7YdBK7vE1uXw+11eQmxdmOZfAWrfgHlZqP1rX4n/tsNJ75sMb
y+pCRoErYQDYwx3Mq8uGnBbnRPf9AKoFuvW9yNNjOXARsjh29sbFtKvG808rw2OdbM8b0d8h8LGX
U6FTQy+eNjMRKJhBTh4A7Gg+LsXDEhW7uNDnujyK1tLMET3OHKqoQ3zu7IZagFnKJQxSdsvGCHAo
2ka8Z/5FfVy87Uy+5+CILXbPYYTDPmCO3Vhdpwj7XGJ9am0xilohFo23HMLPuEf1cvEsUfe+y3Az
QuGb6yujuIQGpXu+LM5W9qocu54YHkKdhXnKO93lZdvF8J4oUvBkhPVNDgg39SJ5fOoiy4QiZt3I
sURsrZRHwCNXtcl4CSpI6v16YaCvu6awlVzC/lPEhvYCGLJtyzGa2MqoTRe8X/1/Y0s0T0upVlOI
XOynANTX4GFR5LS7noR6NqfxxQDs7/M+m/9UUXHHq769Xf+aicW5iXodiXxZLxu4vMiGUWimXE1W
BLPbLZCBOPlD6LEUkUj+leiOBaKoiGYyYXzBj4GJ5dJXteZHVEHEpVDAu4/UDC5nCq8YddCcQLOx
aHfbvoR/dMwYqgey3mLXqhajshV9nP8NW5LBkI88/VT+hiqm9WEo+Qfz7IGs+rk9FBJvoTp8AiTe
bQKszK4rwXl/0Sg8Slv6yk0UjrZuRUtrx30dSUzJ5FTnlWLRCbQeubIB6X+ZYNYz5BDOWjD3FH8S
rCXpzE8hQOCoSb8cq7U2QixPalGcjD+FAclWR4Slx1uTdTwD7wyF3p48HXZcuccQHK0eAwVvzcnA
fc3yMkBIk6Lywt7GoMfKGOw6t3Myps0X6KKHQf7c1gtfrOF+WViDiGNp4F5v5Vy96CSqnOrlRqmN
v43skl90ap9UJ1fLmz5/7w/2CSCrOjY7ZORAIltlZPvrH8rYjoHOhT+6pD4+DXj8jYWdCk+7XmhQ
blHzB/sqU3gheqx95JraJyV5d1UnLbiPFaYONRE6xhyINuw40NQOgZj0ADjDq70fcmEoHnffvdX+
xYEHdnxCkncHyZ7VBby2XteMHhNfk71x9B5RZGdGecWwDZRocIRMnpL6+WSC9sWAsjVDW4LWlOSO
rgBXhm/jh7H3JnWgqcg8s+GlLEfczgrOauUfzf8ha7WUaXK+80sNYb6UmmctRQjAOSVE+QpF5Kv2
HatNoSjgQZa1nB3+w93E+TUHpjImcxkiyIPSJrWKRxEb4Bh70kab5oy6QpPuRB8buimPrlsWT59F
5sEaXLw9llBxK//2GA5hG3/gyuywqSSU15Me99c6h30lvz7qt+CONrPkiBzYr09nMDsB+4hx2NFg
S5Gsi73c2G4OmIUsDhNWAZn/gGSrBvrtH9LMyViD3E8FvFTQUFN0MWYAAmo6zJ1AoQCI19Mz/3tY
vVLYFi5bnIT8uy+PSlWjSzHgp9GZ+91s+0p4N+d3wtDBBCyGJJyqwDJxa3J3Wjh26HPIHhKyWJoi
WjwsAYUAbWwZ0wSy2wZ1HWVk9z0pjJeAe8CLg7kOEN2mZgA7Gfe6JfXgg4OvccLVej8IYhE5FsNE
ncztU96xf4PnqaktdnrARvYVZRsJKDmcDzZWZQK4bYONdIqfoEEFeuNw4+CxoNBZzh0DYYzZQ/AY
13lsEPgHZHmzi8AIK/indYkC0hy3wNkjOlu85qU7Z1NYbpjyojHkZgvy1bT/wHoRj7mi+Fp7h9a2
caIzqDVZ8ZqA2CTh3OCn9afosasjhiG21x6ynp+/BF2M5wIGJ5uAQ7WSblkRHDPUT2eOd4ACVd2O
qmKNzpJ7g3oeUUymYQKAh7Y82YKa+dbBZDJ7QRK+qTmv+6HCuDVwlxSs0wm/uzIB7ry3jrAja6zR
UOhXDhwwy0MD0xhG9WXaD/i9lXLWomSpOCnnrbhe7QQROMD9jIauJAKdfq7rccTuDROFXTNyPe1q
zu2GLuR6F1HG0xkibYiY5JGhEZMhPeviADwqAy8MkTPHpWPv7/vDy0TUpn6MHC7u+vyqRql6sVId
Xfs1QrPHQrvQJP8QEAIYgZddnj0Ef67IbyqnJ7l/0wHn5wEKV5TgeOPZGCjSvZkKv0WyZee0Us9C
tnlv5StWlVyEsNYJg2I4UdGuXyzdAQHErpxYK0zSOofv2nSrCLLND2BtrSN/K3FJCCZ+jxAeuDHl
2PThZbIWWO8OfqYPqOF8grVCj+qpYhr1yzN9Lwycs6i3PL2R81cwrwPMpTdfnJfjIxgGktUXCARe
XMWZZtk2vSTtsmFrVkR5uXq2S6UVwmvSG2w1w+yIXU7iIrTkyo5XnqZfJyqthY4RiRfTzLoLfLs3
XzZfucg64Iz34ddmQV/MM8eJ/n5tQejE+6E2nNtKF+UHuqoZkocF/uV1+Zey0cKIOcSB9pR1UR3k
3HGhbHdAgEPsCedmdPCl02N+gjOdGikQzNiLV1bUTmISMT7QlAze3HMpLx3nb4A3Iyl4/X1daaV4
ID+4QtP1g9Yj6Yd3XnD1nnZ6wo9WNhRoJaxHvFkWZiEFp/aXW8GJ0FXU94EWGTjppgt2XSaZE61E
1x/+TVljI9jeZsn9ZvHBNa/sFJbNUrNDgHeLozVCRlIRL/gOfmlaLhyyEWzeG6++36/SMVda/5gt
Q0zhKGtDGD/CAUG+mBpye4rvfW6MBTrX9psTIxCHzqJrJZVEIJmUo52kyLZW0UL8uUy/lvV253R3
eWn+Rkb17dDEALQgAS+be8r5B1NKvm7PPyLhFi4DQwNTiq5L2EWmG9jV/0Vo3fu4CRR9AZZNQPt0
3PsJAkHoNPV2pVVg80VoxKS3dOOSg1GEJIbhN5T5H9XVYNhpjCYIX7bzZ+zzQbax5KbM2NWjZjJq
ddzNRUkB+VGco/iEDn+GBXkMCloHJ0RHkQWye+rwlUUG8DFeYp/4tEQTzaEX0ocDDJwQKOC+AVfQ
Mdddt4PjT9OkyEp8Ma7HSFICcPqxQkqBq4uxltTP7rcvJzOxBKMV04IL39UTFTk7HcY1Gf7zQS6E
c3bM5K3+ajnTKwNCQFG9fo3DGVjQto1zJeQcDS9f1UL92JEELCk8RZzoNdYfJgtEUpocq0nAQgqw
hNQNKeLsYnasUOnIYPAZqYEc+vqR3vnvgLPNg0jGkBCNJEjPXVcdZeJpn9LLsgTld65h5+Pn+Jjs
S0d9ISTksjrxSH76L0BWUmaijVDLqf+MY3Dn3gJeXzQmNkP+wHlvi6m5lGI4FZVTEDAGERvEHNYi
OhLD0PMNuD9HGV+QK3OXXFC5LTSTYF3YyxLgoypPXBxrmhegMv8HMKPqe5NENf+zYtSuTLWHN143
koJmuF3giaPmDByRJrliY/lS45EGyWf2s0i0UwsJvibKBWxc5ylAEICs9fSvO+inm9oUqOhQ8gD9
+BF3kT4FjtYAoSpW/hN4e2RYrosolx+gnFFFfBejQgk2ktBsJYKlpQjafJZgJ6pxOb3d5FMvQRBq
33veO8NFhF/rKF7nGuDQDCT11QKF29xnuZi1nig4Hk/bD/RaJReY/9qYm8qF03iKbqS4uO810aSD
hnjtb217r0V8mC0c9sxb5J2n8u2YbiLDrS6PgAyYXUYMhQU5eM5ZrTbMGEHcAS3uk4Py1nryXeVb
BEEmApg8Ya90nphE5PKsw06ga7YfacykPWd7TJGb2fI/fDF4QhQcEPU+HYsiCrvK0f0xZ18NaeLO
PCorngrmohdmj3x+jXX9EvKCAmlAqEUBuEXeelsSmBh1KSxOG5brDyoG7jxfazIbTSHEktfiVQ+M
gH9Y9nz197bWgzzHL2i7JgBpg0r4z56yjMzCDiqwfAmnBYzPpim98A8eeO3uHY3Xup7mY61rbgcj
+FWW8vnPGVF3QUBOQ2PgZsQjhluxzsCo7EPc828gs0maZoDspiPtwIYj5JHPF+iyhufR681juUKS
d29+8cTKkrxj/ivzw1QTCmfLQ+QVwSirrfb+VjnvPnaiQ47cyZyIo/wfrFxaDOD2hl7bkK1IjAdr
XdWbIVtuRpADRFE5cjMhhrMkzWS9BFC7xytQKkv/+fJaC+AiNzpz/bxGZypGW+y3V62X8wKJDhnE
VuE5xIBTakENVae8bQieuorn384KVOKwEaFPpUC2pEaTxChoTtC8FgGqbF7n5CRhAz/oP72kHS3i
mC/TW1H5jf0m7DFCO0AKjIZVZMUyy6MDHGWyQ69wEZBRMlYce9K0Ey2UuFU7rJmK6tcq4N4Qvms8
OoHjVEggOTJK4cGmEqLbUkhFWDISnlOUFiPPwPdeqdgSdA0Wyo48RyowGcHCwHQN0fdhZebCTXzi
3KvazaxvkPBcLrkH7nzk5LGs9tZnajyV8UpN4V7PjC+HgRP9ZLB96DOA3U8ddR3303yLRCDQzUP3
gClUac+0XIRV9dTdwMiqbtkbIEBdr9SiBVMe0r6IHDBJfvatl0m5+tT+Xe8TwKHnPvUro/RbxwGK
wHFTAOenF4GDiUG8WvPbZ3okWf53Fl6/yewxqRr5WPPoKwccVYLTfvGkkOBuhkbYh7gYX9F3lMBb
0LyDaMJMuFGA0UCrnKAxReyISEsQ4YUHs6BcjEyA1SWEkpV7z2Cjfft5bFY3vZV8W75gtBkwlNSg
+ZnUxwcBT0vxvsgG3dt7n7OM2hLQbugQNoz18EKPRXm3CtTDXouM5eWUQxW/yDWTBkQ+Ur0gnZYi
C7sz6lT6DXfdLREEDSLoyJNItQijLiHoiLeWyu2CVzPBlsp4twIkkiBeuvNMj7KyUCHNtlZy4uzy
0YYPtD/UzqH23AoOCDJfomzazEt1pnw9UFVlg98BzTHA7YchL6aBL4LdNeeeDePVPTxtEDr8YQRw
VsKjU8A7YlxvKKCcGvLOocYoDg6ACxnr47Wpz0V4nFdRlMvG/aUDUZ8Km8yqk4c4h3R32wHlFGTO
eTn+hz68GYlcrEZT0Vsw5/RETyIksuRxsvytbBDogrUKqlh3bN7KjevyVkh7aPpY8OUD9Z8tTwBe
3V+PKWHSoC3YH2AFF9LjV9fOFFghNk/PTAv1ABrJgbyHnMPYKFNUpgVyZy+m6A5cfMYlpkbRh/5j
0DMRMyMs9MfgdbbzGAv+xCWngVWaUthKcRNjt233rsRbcNIrCEBlRRP5MI52jdLSKiS0Hf2QiySl
jYJPzx492GR/SROqedM/gChcIf0mohFNr3G6bcggUcxjkQ3CSKY06pPu9Aom/BZ6fq9AJL43Qb5o
/wJr5Mc6MmKgmK5m+ymL4JBo+WISmHpVg/73oo63xBmYaWvYa0v3+ikyJ/5KxGZWt9rdpmSjiXZE
JmygQlBYtOiVt8uesg3sXr8AGnikerzqz0UsWISDaV2VrHvw/Tx64QtcQ4kv6+e5RgQNWLWCWG+E
jHSI4xCHXcswuWNBvQ8gEDh6RkLb5/l2cINdN5T0z2X957BWT/1mE5+P/i4th00MozHPC1tih9/r
rGH5SyvNKpFifGk+sV+593pqN7aeQeg4U/HOLZfcXllHxhTOCHF9ai5TfExOpAh++j69hXVq8OkK
4U+d0A2jc4uSSP+zsupoK9cmCxVe9CWis26cIM+dzI4oXe6I51L0tdrR/cSFes4yaoOx3dlcUSnH
LR7eLOPEO/ZArTEioxVb07L7CJcndf+1nsddHQRH5veL6DGGgYS+NNQQFkkv8DR9oORCZ1W96woK
RaQ6YfbdjLp7fN4A9fi+TIes4yBkfM/uIp84cijLObIGBBSGT9KXjWSJjcMGGWsemt6DgrdQRIah
ysvtRuF+4hiFunx8Zphhf1t0GNAMyAqE3qITzVimri3qBj5pKi9XDum8moZDpo+UB7I1rwUpqkxY
HfJ6KNb3YqpUbPAtP40JG0UfxLVARSDMiwkR6EMBaoK970oKC6dpAANLhgPPmneHv2zBt12lkepW
oxNlCf+vjcJsawji0SIfgOmcdXwZLUzpp8bdY5zIkxtJe+y1fYuapLY9nqWIHiMTvfoHTN2QIpEk
Ke2zhh5+gH9kDXWJVNtw9jcr0hoUYk1B3L7xHp07yl/mxKNbnWN6HpXcD9h+MarNBZfGaBi+HfHq
Hz5EJKtkPe6q9di3AH+EBMQmqjcU5SnOYvDFL3PpCv1neBSG3H+tIpRtDXO8xmu5Eiiq19uh87Gi
7/1CdRd8vIMNMaHQIkiAfuNGuLfahVfCDj/03Gr68DR23K6VmtY+n7ffTWnacfF64PlcQQqt3V5Y
ICYWdmnFAg7XV4KjxAaB3pAE3yvN4i+VCU8D3Q/+o8FzVTSPDO5TAXVxUtjNRqLMrO8uzz3+lrAX
1xjy1CwkW6Ik06F57wKaR+nX/NZEvnXE6cncobu1X/+GURD4zEuA4Ku8vy0wYUFPmk5KmqSir2Qt
1k1w5m9ZDxcb3PhTTgA7ZKpvbnYSF9DA4tJsZI3F/zYWduTDIVV+q8h0yCybOO4xZjfJCJX+GmxA
rSe9FJzZGsyaxY2soyRtjU1L6NJqUFVqUNND/Hb7qUrF8S2miOmN0SM0HmhybdGOjZ28Ud6owFsZ
v1JoZQtnFjf0keWeznj+MVz+RhSuQhDU0Mms33nNpCue+bpDRmt4CSN/neKpNxN8LuNU6EbsQ3yn
KbSr1jYe7O/Zfb+foH10ZzWIfNVLrVoTYWC3QKq+i7ZW9kMhYdyY3s6RWnwq18DC36fp+FHGZERu
RXEq7xx09LwyBkA6DgRGnvRwsjKYZNa2H1aLoxGwe4AwKITtAnZsBQP4EBSqMD21qhEqCIZUPbiX
V1IgMXw7rKnwSIOrfb5ENLYj1huRGADJS1ijs2W+V9+Buq5j/ZeqkPgetc6EDlm7uCwTshD8Jsdx
SmwJyT6rIsCLpc9ZCGMrbNW/l/IPXIla0wkz6nlbKi87O+qqmrQfe+VDGQPIRUCvE89IZy2Iw9nM
lcc7CVM4nTVJ6NP585izyEuqFyreXo2wQZF7rpRTCcfaX6poNRspkO6R9rP3Li+SlOoFxV3ACT3H
7K7ooY6QkC3LLQgS/aEJ/lpohqJvzpCK1LakfwOt1fi5tZRadd6HnZUX2FqUKEnaTkrZFAFelETL
Lac7Sx7YmiC7juJ9+7hH9WDmci8bWWkfpluCMLQh8QioGUNFOGtKhSqp8l86z+654QChxItoJA3J
7VxOkRgL3KUeWXjjDYrRwN5eH2wsb/33aOrPWgm0upe8wyvzsKQiGMlfFpsnbrR/0F+kWfMC0bRH
AHFN2Vx41b+C0qpif442W2AkLamlZRCTbl3LI6P+x1tiwOCc8p+MUfHz2VRZS2uTZThYz8+rIiK/
9jLNSrju2S/zLYPy03hn+AB2lDz42jsBdGFSVbqva3sShrYPxTaxSsn8GGDBeFucL/9IyEpDOKko
bsrRklyyAhSfngczlySjyvxUb21KUpHn7OKx4VM4SOhahzwi4up/CRg00ncJyAFFGmB90YLZQa8v
95+6jjmTZ9uAhLB909PKR7dNiT6CkjR94BZ2dqDIP/G9pzun04FoJifQX+MVedJ1gs22w86TPFfh
tzGJFe42MCYqm+l9+8DKAe7dN+79cwJ5Fkl/Z2df/1f+/JJTjAIyDxvoFR8YAJ8hMsqd0iEftQ2E
tQb9YA+6PxWqWzfRWNhEdJHUp4ns+FSuMFFwPPHFUGLbRi0YfJge/q4tttoAu371Nf12pCWuSbnw
/EKFElFCuJwp+UL7u0vSBFK/0xOLFs9lkKRTKZuk3lO1WO00q8pLcXfi8JkZ4+x30GVGyoZaTYu0
VuS5GSc+oxKAU72J52Ww705cgHeoetD6+0K01HI9CsSNQ/5G3DKs7bz/sRfQr1zOmzlGR68zVAcb
KWtkdoyGAjDVTCzPotMy3HyBSePYb7zWWaVazXbnixsSXD/vjXBWgLulyoP4bWcu81fo+g7eWSfr
PWxXIAJ44T1HD9aDUFiENXXBnZ5OcEb0wemfong9S97zThTLfJ9LXjwMK2xzojQeqw4pOc4sMGrL
s8cuwjZLa0iGDzUGA5VgBn1SWCU4YDc+/2gO1Cd3l/QBW5YY4fTmPygRQ/dG8uxVfVWJBtcM3HKE
9TG/zjLZncNdt8Y0HJ9zQckTF8txDnxK3c4ZZE5L0MnOKJYW1+jpSaRXCSfZ294vArcjbghAL3EC
jCbksuOmBNzOYQquEK8yZFSowJ7CcH6ljvY/9g4wHwxna3M5vddAmRezmxamRjEmRhzEn5McE4eC
meN8pLdKmwoBT2Si0fvNq4yMXj7LqnahymnhTZpePvtHnmUL+CZdU2j8YzP/Y5ukXz1OQKLRydLy
8LseukvuyAY+UtwCVIM/FehhDSJ23AxoMU5acAvud2B5xc+JhQFpzo2R/rFyCCFI9wwrD/bfHsS6
j4fYqTxej2Xjkem9iwVLABtVjxGeZRk2ax3ZpoCH6pQIYYDw6NGd9QlLrHBq7e2UGiNB0CZpqxnW
cpaKnDnysxbr0FdttPT0cVwsL3UqUruyIRNfHAIAQf/hRa1L4QKqTyPSw4uvgdt87COYFtqoYBo8
Jd61vh9GsnOqKuZNeYFTbjtUcLsCTLUjDbTdkObDEMpXOUhECc4hGuF1zV9kEomjlrwJne75H7CY
KLo2/vAYbxLIiZiM4NoqtBNIwPnoG3I5pwILML6MpJi/pb2VD1y7RMMqx6n08sxhfzRYAg4kpLdS
C/KfCKKfudXcSQyDnQ5vuH/k2qWfTv+GIhQtqGTtYZueNJ6QQTLbCm4F/QE86eCOkaCHQA/y6zg6
ZA02ZCgvYIY5tU6Jgm1iaRReolamgSyYmFTMsqQ/sxOQeLF4l/PaCkchRLfHXezaIFVqmRxNGJhA
VqiiKslWJmeciyfGBZwuOHwOwXPdHfxJOPjZtM+lRUgKS8VkQO2t9VZ0WQBEpj2Y0Q/1V3EmiyTv
2Z2AfSnU/TC0brMzF13TGZ8NwCYlOCax9XBNJyX694Y9mYQpAleCyUK/JRJmQbZYI6Ov7HwdHMyw
TyduMQvpZAinVv7qvVEKx+8AQHFoqi2wo6oY2xQQIeebF8QxOJSRIDbF4xHGGS3Nu6IwC7TqRIFz
pGChHj/OYHYj1qIOA0W944n4RGXaOIVRv4NUGnU16wfZjXAZQFjPCiAPoFyy4uAsVCLvjKfLh2T2
fh1yFnnoat5rkwufkUnbqzEekQxZBesOU1gUH61FAMbpzQJ1dp/N7eMUdtJxUI+AJB9SJTY8Np0o
V72E2aFHgOCHBYNKt5o7UQG0Qq6+XfNR3ZwNEjLg7TxcD0ETsKFMp/ec7Mn7bdWzY5oQMKg0q8YC
P28DG183UI87OIK2fdiOB9M7nDCtGzrM8i2s+dYPCFBQsJhXwgcPI9PQVSFZDsZROlYuVsOMVuo/
tTvFHuVwNZawRXD7T1PYBZrCJ7C+SXJ+PXhZyoety2qiFh+J869wrQRntM2yRqSLR9YB5cXFxV8L
mX9SXHNPq3ByaaH2kG9RHY8U9xk1WePtuzyE+XEEw7g/DLh2wLpcPaET4KaeQmMvb5nxQA+ILIZE
mapaoWvwGQwJOSqnok4IP0WaD6Ze9C47+owPIi/dMVmG5Boxeh1lQVFw51OMyo5Ky2nO6CBPOovo
LezyaOLwxHTcl44v5noSIMJamuju8xcNiQob96mDECoLnKZjzQbQdJuAVZB2q1lvHLRVLbcNCYZ1
7IZ+NYrjXRTGOFS8krFgiBHZRbWqafbugx04FCibfF76TXanvhjbyoZ8X7aPo7LIJHE3AxXkB7e1
Cx8rIrcEeUHTxVqFkif4xM07kvI1gzEBiRAqMRFCBfotrRrVY1fAsI0n/+xTsh+iiqzaG3tAf2Rc
VZCHDBJ8i6axMJkvWcmoPnby9NIyJUzf3yC0NMizn6DQCOHl9uqMYcmSXEkujOd31YHaoky61MZR
YTDTHYlSn1h0xtKsWhjjnbuy9SXfR1p5VEQXPe7ZVqElJsgLupIV4p6Ps/HqaWMYUJgd6ZX66LJb
G24Q3anvONRXUpE7HzvTolSTvlB/t8gASfrt25pxjllQlUvV6yayo6lSursVKXAbNK6oYlxO2Tow
Wjqm8CyY7HLVXhA/4HuGW+84Yadq1drnz5tQg4f7of/q5TfuoM+RORK1IZzAdYt6KI9LmSeXpj0N
T2WRZjpbI7LJV8lzr8ZaIgc+N2zHzZiBwC5PLK4qMUeroI57KkX9sMvmHRDUmuMECmbys5Wzm7sj
IrUAX/5W6pgeRNNeVB3rigByN0QGpfE13YqB0BlaqcndB6v+R48fwuhCetFduhLAM98wwg/g6FUW
L0boDSSK8HPMckLOsQi4SaOW+8ET6J/BkMaTFMI+9ek3cMAORb90Ai1fM921DEsmD5V2qVg5Jk2E
2P2hZ9UNeMCe8jD38wbHa3+fsDV0azQ08wFhW4vMzmPuFDjy6d0h/RuHEMdVQ+3bl6ehUrxnCrt/
+Nu1k0I/6OBcRTGi9MLTJ+FwSQ2kzEEL0yeQjEVnSJoZ6DyUTVdRInaRCxYdJ7aKTHsA6RRExj1q
DDk5j6Yj9v/PKQMAcuEveVZM5yMR011LNDsWaqATcnwkSeXZ/JSHsugFVpeYDim6smn+PCFVSX34
DGdGVRCoeR0X/Uf/6/X59eTwjujS/5svFxyR3XbKOkOMc/Gu+TNS40N5zMtmNf9Ejg2UqRUwbU6N
jMITw6LTLkyE2RQW/9pHgL1+sxoEDeoCyKqxVLclLOSQnbpP1b9eT7iaXXDoYVDK2tw0DeYUFuDH
XzER5UZHWaSR7Qu16CFCfY0MEVkWWHreYhI/lENxWAVWEktE3IjM9MLCfQTej6EHFYpkl/nNkcoS
wR3xqIzGR6r+SSarIQXKXYXLpww6Src5SeZp5BbUqxnd3ITztx0Hc7zXYWJecfOdjl3O17kj28xl
0x9nEWwYUcmSZJ12JnBlew9PscxXckwHYHYT3Sc7ZCq5j0lCppIdaK0JKOotLuuELo5gSyyvs+QY
WMXpE27F+OnaWkTUeatCv7qDmdQ7/+jev3mEPUnfYQqzFUV5cHKEQo3Xh30Ph30ClWHzmaB+ssae
xB8UC6nr7dqJMxZRFFdPw+EuwHQIGHLLOVNlDRNhxz+19t8swpY0Zq0jd8bWESRsYlA76zg0CMRD
DUI3jdO+/phAPh6yaVL/vZdQn7zLFdLTkFxSYRiFycHhcQp5o/DT/hVfCMPeL460Lsbot8TXpVE1
S6bjMTluPqt3MHG9tZo7Qo55ugsNFzPgUdfGNXc5Be1VlSE7wplh53Adu3kFirXpt1sbMiiO4eZ8
ivSp7ev9B7SOvHIv0qzxD1VPNLZAqSR9pPziQKoKo+wFm3Ywz5qz/neUnYnYm+E64IhAbnLSeF32
OtIa2Z6gJgsm1Sg9u2qRGe7ZuugNhaF+sDfxxjGq3UyP8SxmyAFg75f/sEItHHEA5Jy6MuApnvMp
RaychUa8/auymbkylzderez+E8o8mMGlT4nmLonPp+F6jQYlxFQ2eazzZN9bskV5u821kJKAKZlX
QYn40qgTGkxI4m9gORhWzMNm/pqy+gdBWgdc+eCmNP34I84+hMZPtRH5AXp3N6rDz+D6h20dXcpR
zTM3B87rmhfgY7ZCJvFNtpiTccXob7NP1MFM8NUFuTkYoQxITAgf05USlahfYDblXDvpwHAlk8WV
mYpK0V45RI+xiAYo8FIaPqcOqRdpBSTmCgtT5JN2PR5jfmdQE57DtK8PIZ8U8MwAAekzdPU89zUm
9LaaOMIsJUec/WrIJhOtQyeb/8VXZKohmZN45r+XNwP5iETqWoilMQeu5Jy8FeDDYjv8/YmBMu6M
Oxu7YeZbSMQj7auHA9HVuFPVuzcD0kze7KS9XMHwyXltQ+XEX5kvgRlXFwbV9p1GkRSj0GTEprO+
E6r5rfv0pRpXdIHs7o29nMRjvOn7OL0orWsVAtN1dKCRuKzftY+xVbKTXSY+BHhnN/WP2pSsiDzZ
2H50Npu00r6P7bOjR1s6HxTtSUAUqJrVwNUaC9i3VJrWiM+EF/8eyL6Ha8KzlRJz8H8OZRX3KWEq
yz6FzJORfah33j++TNNcDTMjwi3klN70vOBQ1gUxeFnIO/iBohcwO6RkD7qakfN/edASfzvd1pqC
uJn7OZtxx3R17/Oybg8qWaOA29gspJCrxTIQUaQeFn8CGUrwy01I7Wrv/8Ko1cgk4GbIMfRae+8L
d/FXwnayzP8VZiUdZo3HfsaNZaxq5Bkwk6Xl+X+qE8HigqW7dvTAcMd4rGwstzOBCx7mY31S1qXA
Lyz1TnoBtWFqXpQnJRyIfzQtenSvSc1fK3+MDA9HqCBzq8vzQ2x37/lFac7+LsEBpe2NFuZIuJug
lkhzDh1wfHc3qTwbrscX2IMbRGK4DH6SPMDOfmyF+TGDutjT8XY2Lx2ho8Uh0LkLZDIALNq0lFRC
kv96erGqLDAheyyaP/D360zEQvNZP2qfpjSuOOvpc8/tHxRJOo6mwt9UclBInRrY9SwI6FJmQeY/
P9ANbhxnCxS1nSABlQR744J4frU27VbnE0INDPcud0ljnNI6fUSa74fmarGzjX5aQWB97LQegDHG
1g7dJxAugDPo+OqvlhdrEqEuo9weJdh3PwYgUzbn4arH7/i0RC5hLpA9vLWAaLdqRPkStQDSaTXJ
yKFgqAua6rUfJorpxwNvwxhkpKFncIvGcbhwU3xl4MCRM1u9DG4xw370QjfMWyJASJn3wfzkqgLp
uqNmb3IWgUWBHbvryZ/KZ8b/WTajMvG4yA4gln57W9lWTu15tPoLTDIzYTWMS6fC8yR17ygMVlCy
t66yq30P2kSFEN0rGv5dJelr5n+jZLxASOdhdxjsNxGvYXh6rDfwiYNCjip7evhPXZccFt5xR+oR
A9gYhIzu2ZJIWOLkVZFSuJ0kyRMKu9qLLijFvNO7nJGIUOFt1cEP5rd3KA0xlr1gHxZJJBgNAATA
c6bEeSaQM3cUHyCn5PJm+fYTzxPDVp07oEWFvGi48ynWA2NdlW4pvTD+fnzuXwnPDKcV0OTJLp0R
JG/eVleTuxxytugmotHPQOx4RgGgdLu8fe6DOGbdNrkfWh68UaNe8dB8GfABvk89S2nEmduCGTiR
OdFlQS1+u0NHh5erM92yo9W3DVhPgmBByfuXjcqcBx31rWKQgIwYp/gwQVJ3e02BcXbX20bQaY+9
XM2Zw+/VJtkz5rwO8+7Z3LtsyMvzLJdCoEiZvU/clXZec9PAalugy4TdExyvg6TvkascKOJQ53LH
7555NRdhm6DTWGo99VSYvGdpPz1RHtcYEpDgGy8R/+FYrNvldjNdpvyRQs4MTeaogsIpidH6qTOm
TuCLGFUGiBVe+o+9NIyZAJLfySJnFVc6vCkkTQNX0O7dJ/bBI+VABIsn8O85z7YABFJwLpm+eVlH
t+7mqGx8aT7H0yzc1dI15amq+ss5y3jhIvHaSlZUjekRalPe5OX2xwthd1aPZYlRz0Vnen/+8uEZ
6YK52CqBnP4bffbE/3iA9cZByPYKG2LIibjE+rZjhgpHx55+7rKvLTOG6BQqCPV3D+otn2dsfd3k
qOTZuaBdE0Nl29DD9uQ3RweqfE5GEhLpPZyXBqCwblBHhrcqRxJzeHf7TMBuQ/xYdj9Xi+rgqaOZ
BQHKfqmJKN7/yYQe8/MgDdoQ+chzH3LlpRLW5fgn+YNdlf/BJVoMCCxqBrsnkLYYpJmZsvplix8j
vti6qtMqesjFlZGyJWRvL1Z5z4DJfrAbHSCZPOixglM+ydtKptYZElftklv2Q723AyBPcYAntNn5
JxGx+Hi9sHB3wnLfzj6Qh+a1/+GnlpK5LnGwDyjkSCW8wDJUNGk2jZmdD5dghX+Vgok15DBAHGF+
4RyOjwUDM0MEeeaCk6025//a2N+mi5VagRv6JjBTRklffVg0PWjsRAe4t+X5EwIoyxp+zNYfsXsS
NNmc8cqCm4Rf+gH8pyaeIxrHd2Fz6aDA8FgkOnWEPUXY0sRrofTde774HZJ0xT0SJ/5UD3eSNNTV
+8D1dZ7OHcRl5XmtOsv5lbJvvzcADhEDvOS2I1n0bbPMJmSAvp59mx5YYym3r96Zu8LFQ7+X41M5
RulIa/ZP42c7cu51bay9JsLwBdKmtAumXHK5tQpt4WG3hQg+9MWpUZTYgtxgLK+qKWHmXo7yZNSe
2ktiSeFmQv9yPi3d4ygXlYj8B6KEBkPVJZsuO2hjO7zPpmzFwml3M6bqK986oFvNsZpPiWePzjzD
Hren37GiOdPlF14DZOZxZUMgQurSW8/thkaYvQl7r8xE+PSKCjPsx2v5soJ34H1Zf5TIRxbOATAA
Rey6yOeqFfRTaSiZ+rUqA4WzSfx5PeAzpAbLk08SO0ZqIV75I6pAcIohE+v+7hF85cFYhyPeEDQW
EMQm4n9rUHPoIcOZKCtBpejAqgTayHHM2ahUK5f8FNHJNxdvvDfDBmesUfnJvkoYSC6fY93tyIt4
WGRoIs+GXgzqJpPbKhvAIwMyaDekP5Wfrr6SaROysDd71hVvBJuiZK4GA5ThppEsAmZ9IZqu7m8u
CI9GlQmEbyJwmnnmS5isB3JT6XC8OEVgZo/19SZJ+uXnGUTFTHgPbrmJ5HqSOsdSJtsGh2KzW+zT
gOc1pRry3oN8cx/4e/fFzQpjI7xLG/5605itCk7hsiHAhY17jbLeeValwfvMAfX+vFCmBy225zgm
T0KIl6sgfVPTlXR4VjRz6c8FyHAwOVwEhgx01wj5+O6rvzaDKYNF2oVXbUGgcK++Db2GUHdU+2nU
5aNjD6tRp6RJ4IJaH8Ikxq7MREopRTEPm6WrbPPVn8l1AmpHSf2dRJ4QO6+QBL95gXD70FHD4uP2
I82u5sjuNJa+D76gyTvOa+05gcECHK0w3SebrXSSJQfaR0+EKUczJiuSiTQ3VCi/BAJFFDT5qgGz
k1U5IEoaw7vegMHoe/vIIjvWi//31stxCMeJOrEL5uLe6IUka4gYU3yBMSkJQI1MMcbPOjBRYim5
HedQrlpFVNUe+6vkvGOcgtVGfN18jZ2LGySIb8CLEuXQPAFrU3G44lCLyu0Nc0lfxjAfMBdjVCTc
qRUin5CC+CQurnkEtutNBKGgMj9V/bImGQe/iN06g/8oOR8Vupj2DR6dYO73nATQaSH8kOXJiRiU
eyFn7uqtgA5MiqfaiZw8p0qfbn6ccaTo0z1noJhCS4KRgx5KjHzHkRxlqE6dEEbeae81f7Ae2rnh
tMMCs/IrE9llA/rdRgWePlvJIdAT+vRSPdDgRIPp1sljYFoHQ58z7VB+GY8IBXX2iBfOduqlgGL/
PklFFhzzJsaPfsa7lY4iewXzcg2KW3plPh9l6uz0xLZyxXYAkt0xWalm6jOJUrnI4PFjkOf/Lgeo
nkGbbyBjnE5bF5VBA8E60NnjLJG78sVNvECYzyejnIOLHg4WsxsAE9nMCSI+nmzx1lpCX9nqi0Sx
NT2wqwtW/wTqFx59vtKnFzMpIaI3zUJuiSxSs6knlftMiyo5v5W6Y58vg5cEF/6/Iw93NkPhp5/Q
+rnmIYdgi24LYLfDbDhaHsso9KX8SOJ7dwe8xBEizcGLqzMP9SWgkQU0kiOOj2vjxuvbtuXh9Nhn
Hx4KIrHzt5rb41R4Z7TNzP4Yl0jleTErpLo02NszPmXsR3+b59YpoB8vwAuPNsQKHkIMHCAeqmKX
HcCTidepFl9YKhazfIoR4cEk0EHoQA6Nvgk/wjkXvkmoq5PhC/LfRm+FQOzUC+j2VIdRcU6B7HSw
y+qGcbeAOANvtFUgSHyqR7FNY/6J4ayqb8+lKAI/fn7b0JSdfJ9ADyeaLVPbBmO+hCATmTcHjo0x
rvaPUsDpRfrvV/AfEAND7fhr5s1bv8S+4bRaWILyOAWsoYgKcnyEUsMevy1Thmrg6OE+s1un0gaY
SM01omjceSxzyWYBSsNddRkwme3H/C1bIdfIDrGZG8xW4o5i6s6V07s08jdEdwKhv3r2F+pYJng5
qot1EpcOeDi65pnyVL0iZhygE5i+rfIlR3CGYB8gT/qfWvwowjuoCDDIAyXY3GpdlfnuBHqgxgDT
DO2ckmiE5XyT1gPO8J5x3HeZBqCLe3ULgIawv+LibHoXgf7bIKhuhD1ekrNTxUa5EYbx2BI8Uv8i
oAkRJFrw54jMUFcx2Y/8c2LbTuBfacJnqp8nJl0x2G2JMDa8YB+X40uU7vBqaLPhKJkX6pg6qt3o
cAfySpHnBlE6lsmCEtX7fioRjjbMDoUCPX29OECvqiBOiEqJ1gpMPEFTrcVOh8A/hku8/4Thz/3J
t4A9G13vYWWgOVdOhnE0EdPO5c4Fv9DciYmBGxbktLwXifRil3zVu4aa3uAheg3T8vudGyLocbNZ
czUU0IoFrG8tyqYt3tpDKyULRQjGWeHPGLMCXAT538OGRxQBr3SVNuhUe7LrVeSwDoiCTh/AnrJe
oorENifVoFiXAn2EZAc0Am4mNkqG4ajahXlYptxVaSCMsu336rRJaIvTdouglnEzn/0Bk6MyEGX6
VtxP0CXTj1wK88EilCKCwmrIfYcYqZpTb0aAnhRs58a65UF4ARgPNZSQhmFVpclk/xP/fzj8TF1S
4tW1V/Xfhk+OoLjiJSbWlF00Q29EV6+dt43WJftUXQTtxAzVvZA+47+riD90Ctnxw/rrzubqpKhr
yP4BzmLYGMK3XGHVSO5BtEs16J/FhUiPyzRz+Yyt48Utd+LGbhyZBt5L6/Bm+APDeVEPp/a5WcTV
EgWVQAJZUcvPo4r2iEgtQd+M5BguxTEiWbGhxNvxWInPdWrErAnop1v6RCHmCbBOCH5e4jStnJGH
PFQnJtgysD2eCJfHjgiKiyTQ83VaE6TadLgqErugs78ZAAREXI6LdM2cChs3kQj6RpOSVFOItg5G
iZOugGfAnNVfGz2cA7DVuAHFe3DiDuG+JbU9ZvFFxxny6xhdwPSLoHo1fm8uWwBvV7fr6GwKNqov
QR6/t77r9NHhPQbteMe0D0XchnaxBVVIeM3MfXztVBs4ahfdvXSDbz/YXwMS1Z52JoJM6Cru1I/Q
igNgOsOQhlELnJoe3Jz+YgXVK9T3zbvGUQqyCG+BZPHoWTb3jN3gWLG6dcsr17q87sx2jp3pRfs5
YbEMnL/vBRz7cvWQ8KyBr9mzSZxpAKxjraMRLdg+j1OaLIsCaqwsgsQTV+mFCEh+le1wh+tw3+xZ
aJyBr7nLI12A2Vjms8JMcJhURF7RaXdy7hNTQvabH2ER7wbgS6YIRZrQgWh0OpQGcnmuf4X7/TTc
NOdsux7RBdnfzoADVjAAlT4IcGgAdEymfDztdG+exVY5qa5jA6DUje708QxdMSsLM3qjy5t8VDjJ
xjVyNKyR/HZNryf0Z9BKFnY+kWBGJWhTSWNB9poxhWVRWzoka5UahGGisHxwM2DZZT+89AhUjuyM
JM+iI+HUdACx2UwITpgWhez4OLTcQ6w3wVmootYY7KHoK3jwqU4iXQvOd/vkEFmp3+jrK4W6m66D
v6mk4yGerncc0I+6om8QmgP1bvaMyLNz/p+uDoJ9Nll9ZAPxlWKBE7uwufeFPL5+rSVp/Kj6jYTQ
YHscE7NHV0nl2i+qAYWvqGrGwp6NVchOBwr/5/NS1uTOWGSE/DdCjUm+BUUAzcogyLLpj8p4aJN8
Ja1dYC7yS3Vsfbccut+YqeY1DDAQFCcZAqXxFE7kjyoO451Nud/bX9HJl13K0Q4ax8ki86YYOI4g
LXteo7cq2hmzMRUG3beH9EBTCaMlRwf0EGLUPAzsSEVdkm09wVShI+03h2R0Jf1+UKnlSj4YauZo
X4mADSSzowo0E7CuoBf4HYnp4K2GPhl8cou1jGBgaFvButsk+S+i2+VvX5jUshFf/S3907Tc3j+X
jX1p5SEuLp/eLz1cagpaOp+DAcn4Q+k/r/hoi8dbWTHOFW+/Lchf+3MQvNyi0esE004nZGrzlF0S
0kCV9/hZvFhIA5oCe6n+/4hzwMuSJh+F1n/jAWE9XyMkUuMfOSuZ/XX4w7kdwZDMHm1W3etGVC9G
hXeckTLkdzj//nrz79KhoGhYdLGaqHUCDTr2n60Ctz/t9wKQ8KkDWrV+7ryyKodAnw2mcuOcR8zC
dntHCA/kRaDPYvZ7t+yDxPc43DTmk0OsI9w9MH51gVhb9HBB/I1PHt42cX21K55SnpKlf1X4k001
OWh3umqpQ9i63T25fHBGLMAMw9gVgthdiGk+LyBYfEk9jtcvEudBCS7feWs1xzeNqFaECYxk2d52
MjlNWT4zEMqDKtPrwvhiTFnZdk45NZjU+Vc3uaiPKEur7Al4FSdo4OEbaRzTzlTt1msUHyy2WYKu
oaXlXoaMI7uIZ4EZUDsh8LG767owApBC0ONxooxydeKV3iyjW0XuRx7vBqcAfiNVwhbaDWvZ8MH9
prpbgyNCX/NSeqQAMP2M6N9f1ErBH3xfO+BMx8HbU7ae4p8GQEZRMzkzRjWYAOnqCnFKBxZclkaV
eWJ5VtwfFmcTBk23iIaa8TL6toq0CCYOCkRgx+XrAa69jgOO9ex7ru7s07NjHwfJaJTR/Gp/lbNB
GKiwz6kCvtptUUMkKRj7+/mxEQ4PV48k65eYUEpKu+WOL/Eeh+Daz6wO1ya9Y8h1cPiuEfG7WEky
aquSYZcTrFCdjhWJAJo8I94VP2MBn8VX9CNUGqi4EvVTEJY/4ilkIrEGczT69FRnvylxiU9fUkCR
K/RZsoWSnxa7DvXu0rRkYXfh7qeAGmKVHhTfQL2sjRipomr1z3tqxZf/B4ovT8DDbZu50mbcn8zW
rWsOLFXiz9h+J4dilW2+q4IU0s5M3v1d5drmod9Ag2a01GgnN/9KM49AfpxPGeZJALUSwf7xCokS
/l8Rr5lXqpocC1LxMxW/9ZMFBMz5p130/nDID/FOS3bY5PKterQhoyB5vr2Gt/DXtJbqfrF4fS59
k7iPRwJbaufQraHaNkdUJSGN4yQPiOVwPGvP1j8zCYK3yxBPcJ/UggxPRPm/WdBaNCGV2ex1mUSB
B7F6VYbhK3sy6mbeeej9aUZTv1DpxoDT8b3i9Ed6HfGPxT7FVDHFkNRpY5YC8wsaPEksnoR+PhN+
yV4k7L09pRF8UQBWgfWZnW1bdpk98V5StWR2NpcaNZ7RT6lVv6nDEu04vXm8SrsvdodiptkGZlsc
xhggtYLH5DBTm0PaO/0M+Lm8RnZr5nw5kW0X5ohb/4mC7l2LieUab3Ckk/pX1yW0NAUSd8GYB4Z/
A4wHBhFpMj/ZdrMBuvQyUigBJfFo0ve9SF3cjrwE/N+kxb49Urv15Yx3BGHEfSSq6kTunJWfSLA+
Xle2UOxfemSqPgT+8dcTnEOnNFQMtSR7bEKCWsONbMm83p8f7j8FGobRWiltcbVYkKoWmWSEbD7c
jDIaeWAay0qlsyoh/TSBoDagzvthp7a6zqtQ88oDa6S9oLcwj7TPsvIO+aH0YOAcaUsQfHnCm5of
MClR6iSai0rKGnJg1Gkf0rgt2kVvx7rCzp/Jgx5Up4eWjcQOYfXqGa62k+7eWGKwgF9muSlaKvrb
Ad5FNqzOL26WERWLFg0CHdEaeO5kHXH1218osLXu+qCmbVablEzwBQqkSLTk62ZUNfCskjeKrGtz
98d8gIe2oCnun7vut68KcHP+AbMnIm+m35F1uakBmE8/nIS9+QPOWmgAsptjp9XbS5q4q1N9ZUvz
ybwEZfZ4Vm6A2+soVhAzUexuLnc6WRNwhuWNA4PI3AgbeEUW+MQvDyL0dOn36adh0/BofR0bBGf6
09bFU4xd3B/omDssrk/PdRMbhFfqgOALBPc/CRTYt+M6y1qu0zlWnbML2dQR3G1hwWGsme4zE9mp
0fE59Fqn0wiile2Rj/8X+Bjnu6vLXD+y4sTq8khpsDeQ4/PELm/VUoQ5lNt2TI1jR66nZ0nB8rCJ
TxZh9FwP0raP5IaDr3p0UmvLPTELPvpxkl2UR7YYUsR+WEYtHokj/jw2VjgziPVaEeHKsmr0jENZ
I586FS0HBsT/IIwTl2RxtJ2tEaedNSV49RYJ+5XIvdbPG3CL4N1pAuCdM43s3Zv00yUuL/fCkqAI
cu6VsoNwMmhTqWSJZ2WAL6cnc5cz4i2lw4S9mtidKNfR6YJhodRIISUN7Q4mI/y8lgqbidYzow4R
SHgauQ2zM9jTYBW+eoAxiXWeSA2R12gKQWXRlgfbFUToN1VoI+8dLMslS42tawDrCiAOqFF4nBOX
l8rZ5B7k3n2T2jv6QPOo3j5JNi662gPA/m6/kdPeY5sqABTJnvHHy/Xr9Ofo4a+QA3nEN3wDtbrT
FujKfIAgQTN1/MwuE3ZQ5lVS52UnpNdl2KuxIdCuzonD7J/zUkamarW3xtViB1GQsLdBd4cRNk+i
EGfMdIrpWaTtfh7jwfZFNnZ1bVYuG/WI2suidClZElPdwStX19XymSuuhiGPKDbxWV51/NIpdrx9
txpxGa7Oz+VQh5x0YiNN73/cQ7IPjafPPpu9di80kBXgoF12lB7Z6HyBA3oM7d3hpBfmk9ksYE8D
/FhVgqZbipN5Mor7Me7Hsgd2vXtVgbvZkupoO9BZ0e5o3c9jeCmeUljUqsI5MphTU/2+lTs9iZXB
Dipsa1z+0ASKkDkqSbfsG1Khnu2yP62EgCudik/vpg6D35L/H779kyamxFWdQHIONpwoVhbL9dpQ
GdA8Bs2Ly4tmQiIQoTAVnxgFuUodqkOOO9E06zeDU4sU8hHYTzNgCYTdl8d7loemhbjW6QZPKxHS
jLf1iJx3+L/77kq3u7AsOMjklGadXgRxg+KUTzMss3y1fNwvxJcdh1S7GRzCQN38sXoedlWtI0sR
r8TeTB8luNH0LV1IX/rRIV8S6Tpvdd62VDZg8wuLI9xBHZCfb9fIxmV/HNxzb0NEIfsTOKUJDj1i
9hrblBC8bRP1ihJwGBJXWCElxiHBLoKGQDGVByqzlML+XBZnoqKwnmIxNa15f4TPRPzbP6K67W62
Z3IC74H/4OdQ1B2+7tiR0ZCZBVI+5dxxV/pljM4TnaK0LnkC9cVax0ycWfvFUnxa4mj6DMxUvFrz
vhN3Aj5/VbLjjeFmDYdW6kxxO990bGyTujEmZvVvkl8qJgRkaE8sU0Aq5nnOH3j3VEA9vrzoEA03
ct7L+PBCPSfrVH2Q+x9uReMX0+dFqrdQSv1ucA9s6U2+6cfLbml7ffAHXGImGMghB+Rv/N9NSrfw
9EDlI6nUqN4ez1zmwBNb1uY5QWUHGapVZt34nmdtkAaicwEiRmeZWenCmjscm9TL7Hkzgd1vx6GW
T0T2RszdGn++cx1hNzne19DD5386BEjF2pVlhoMW+04NM3Ozr762Hc5VcMkeAj9iYaBsdlvKvQ79
nm/5rs2zcLFX27kj8R6eeEdj+nuwEwmud0u7Vw8yQZaTKC9nS5QH1VoWmasr2PcuQl4Y3oQsr80H
D2iUzMVZjVrFxr7J7ukmzYIhUuP0Gk/kqWTIX6Z5hAQq61s22BjejRbQeeoHy8riMtxSKHZYynNP
/mOUCvWMaIsNvSm+VrNApCSqC7YEodpMB80br7Z3IvU3EGyjnEYAV1qiVJBgKMlmn+bb/kTAmjCl
qVNnFaSGtGqXIi1iSWO+khv0Ffuhv4N6d3iNK9dnWZOQ8hZHYxDyy0DevAObCbACRhCdC4idtEWI
N+YSwSHn1PsVpCEKnwIV6rQDd91jMDjiEa/bgiwIpbmT9nfE8c0NOPYHxDheIW+68aqWWjqgC4H3
V7lD8wKkZwpL8dmIEUeWYHhnnKuFFjBlDVgpLrnosrqvjbl1rwipa/VEbkTi77w5dQ3Nicg+yH3U
oqXX7gUEreyKmNfHCuD3QhMh8xoCAx1JMcTBRZvLNBW2Vu1JzgZrwi+QtjjF4a4gd+R5C50odXtf
h2kwJIdfOmB1PsCl/NpEiReFhL34FXuniS45s2HCGLZorbc/7wFKZgxbUz9Z5n/4zspQkaolxpdm
BfKW8b3aBKOnGnR/++SoAJhsSaRTXP6i5CSqDdTbNpuwcyqgQ4Cxy7WTw5x4gyNJhkqlt+5D6NSr
zdYcmXFZxeiwdZqLHk3eGBPHGeaWK2zil33GAGGB5vCK+0k75Ml96dSql1mo15dsOqCrdpoO8+Yu
EMyXPUyJ9KMWEW57JSLIrvrjtrVCvHOtKUGATzmlfNplyeucg0Y1OrD1z+nSJ1z7Vu1bPpfGw4bd
KEfQDGNoGvqqC82Y7yEE1In8f9/IQjFvWGWl6Ry2uIjIs6MWiWZotGJpPBg8kCoWlqIoJNTb4JFc
lARx9raDioNHlXSA3hcECaeO19q2aBKZSDDiHwpCp+Njm0ab6BHDvVOd+8awE8JUf2/1c4hRyvTv
f0hqIUGyPh5N0HNLMhMQ9yakXiHhcXKUTxcReKqIKAEYI9gUTGoB2f7xA2Tmxy1iECYgIgNIPiZN
DmdrVEdeL3zlo6b8AlWKqCHCnWOaAoeZ4K4/C1mvCBLCzgYJ1Hy2MrApG1g2cgzB4z/p2fbEpoD0
FVz0NXt/+BwSr18sZIKc2rVKv4V6QFSDqAFuvtEC1fZ/DL/1S1byZ8DJhv2++OjffZsauPb/ezYo
efHo9rcjcPBAh6RA4bcPyEeka31RRAvpoaw5a5Axl0HzSDKkhlUI4CRVBssltQ273rq6AYIml4J8
882Zni6hKrQ529x1vDul/o1vrIQYBRaCsHWWf3BryetSwgYCaetQFNcrZLKGwVIo7hhN0O3u5zQ8
B9NtTc5r5p6HeiKzCpKSFnRc0/4hIzBNNvFBAj55brurRUwYoYFfzxt4/0M6dbcX7qC70MVF5MGU
BFxcKNjr9tfVa+VdmOzFBTxaMpktaY12UoVt10Gc9k+98Mz6XNDPIgNQL2iMoSYXSdkB39P+k/Iw
TP1RaiAgCfQ1BRpBeuz1BErYvuLcsFpgRM/Ec2Vd97lB0EW3gMfoUxaA6plcyi6NEBBmBS5S+lWX
1QgiTm0T6SEq+PS4eGIoaFsWvhQVQFTR/R72H40PIRNg3K+AW8ltRApYCJbZR4qr8Xm51Ux+0VGE
Rl6/2aDa2nfoFFtMzqoyfKC/TA1y+H5Kum6Blx/TFqBjXM/FSv2Mj3GuuJPj27RlON4a2CWGfq21
bbKvr6YStIhGz6QPngQToDAat+zfHJGTkQRN/BWnKIU/lHCMvgrkZpjkKyJIAap9TZpVgxKoKq8Q
v3H/0aA7STZS4e9skG93zb4O8A89QAnVHHZqKWM8JXvXrG2VCza1GVuXkUaS/JYfWV7eVO0t6XSM
59nCMoI3UD+CxNr31FT8G2duh+xDX+SlOXnyjZhxuK6Oomln+NbsY/PVmHIriRku54lWmUu5vWhX
x4St8yJIVXiQQ2hncxlobvIEk5XcEhZlHqgfpXF9K5AXt88W5hAU+rYa5OiYNax6x4PF45AUT7Vy
RXcZwKY6iL0p9VXiqCx6QXpiGzO/YTsamkvIeFT+k7LFzZeb9OX4oaLSPi4ESt4yKPhhJWyoNLmo
iE22p5WssY3ZrE6OI6u6OwO8WZOcA0a+Szy9Q7QK3r/gAacz+zgTluCeWXDS8+OrtQf5TfmzfKUt
nGAl6bIOFXJukI4FXHPEo1Az3iSH9OaaqrI9iVgO8NCnNnK5UeXH6yZ+iYy9Fso8wY4rZuuTFSq2
S7sgtXcvKj8WAuwaOvEWQShJX8UeWJ0aPrQoZ9U4KJ20kN4iJUcMhvxY3hbVC6rRo5rUTKgaNQjS
0dF9X8XXO920BKx3KJ7mIVeblSNaSwI/+4sqP0cwXDeEP56OsT6KxwXpvlefUlw81oaoP8XgdHSa
wowgZ7CNU1LGLQt7+iFS/sp/WSw+CF8+1zL2yq9c3D3U4TmIpcVLzJNwZoFkHOUTIVxZAw+VNuY6
0x8NA+Ul7UjhQAOi8sFQVmWGu8kEb9dORHGiudIPWO0v/uwX3BIVoPUPnxLh+Aldi7iKMCM0Ap51
kLzDJQ3KvoqlV341qK2zyyPASIGLWIUD3NrPyVHLzKHFXAplTz8ZsjiutixvKbzeAe3B275Y63Wc
0kcpMrSR6dJxfUNBRPkayA2ZElAxweP+02DtoxTTjLfIr3bDQIjXrg0Togl4YfiPRANX7CaZCCqG
hD9MVqX4567bo7/Pk69QwjLNkJCJ0AP98kA5Q4IhCcOqSc66tWArhwBxiepSzgLoM0Ll8fX88POM
GQd/Aocg9AD6nf4OJFPoTbsbBZlU4Jsb9YIAK0Xnj2A+edo2gPjZKcnYXB9FLdGvcPB44lJqZpvd
MF/TUk+/ZVDER3Fl28fiuh3RtBwIkILXnAR4hvErpmIYW/SFHHTAKqVkN8rk7Ag2xHtfvZOW7Xo/
L7WVVhHJUSXzilQXWhEfmFKI+jOrb0oIy6NRQ4qul+MzQvMvz1riS+8ikNj6XFO9dgsG2LwrP2u3
WC/GfIVU7fBqoKqKIWWgDkqo9sKtaeX1Ed80E1v66RrB9RmbznDOYEraiwo6+76Kt9FNNc8JiiXR
nZoypDT4sm1D9a5HydXnlOxEtE8aeRwvbef4AaU0k4tD3N7VCsuiZbaymLAMpt57ju8IRYxWTBSh
KhqTJdVJXxwD0nHfpU16nrQF2iMeyyBgocZjwV4bRIeoK8LpxAqqSh6AJ3jN9SopuHnq77TWbZ1v
/SwS+/pYxf4xMhAi+qL3WGq43eVr0ZLiqGn4byDddftXDNB9HMOY/l2UbWGDVfkXB6IaE/yp3OVt
BSaYEoSwAqTFF6jVcl3kkr/OU+rPgynwSt6OUueBZC13qYU46Ksy9nqgdreh1qxSM9w8ZZvfu9NT
nGLgI1AjMz44vQlAM9NSY0ILKgy3QSCuOWZzgXxmIR120gAivxgkdHgRwGcS0ao4/nFJOkumeSTJ
MKP5Z5+LneQRDrtJ1sB+yFYB4hKWlFwtgcrnzAwSqsRhIEjuWO4xndvGdcYa/nLsA+P9LTSdr9AR
xMZLgIhrSV/i/ldldfW1a7XK9tqGuqkeXqfXKvM02ZW2DZuMQyYhEH8vFJ8E9wPcLzn3P/N4lf3J
D2g2dM4ziqpJhsSrjWR4nkk0xD0Bi3q+4OMaFSFOYBNbRU/VHv+ltBL+bB3//6i5chF/UGx6LzsL
JPNEcw6X8tzNQJLkZ48pf9/IE4H6lSsWKYhhKB3TeXE+fTr4ijBAq9TWKf3r8oKaAl11K9Xj7ijq
h/GDS0JZzRNEcslXEXwOGz9FZdp0yhA6fuM9TXdWQZriSqo7+bmeZsF3/9ePXDHLhPuXUb1bQgt0
nrv53oALxAL3fHUh7G05PZnRAhh/ignZF9bqIDflZA18PDRUVRJ7UcW1iX+EDLv1BaGYzl7p86us
JPR5HoAsq7MQBPBs5cCebuu4+TpDU+pBG4oJoIeNisUPYufqC9pgxk3cGv2yDPhK0IbLEWw7WA2g
UgcjFDf98VSiXbpskUudMGUnoCe8I9cvgwoV6PCVPiO2962YGXS3IkuIrGfE/8P3barlJtbfJzVe
u3sqN1ymOZ4R33dmXPEJAIR4I8H2RBhGsT5It2Nof7yXgfrSOJfDpQV3N5ZMtb/9yoEkRXb0sndJ
lcgpbU/jaikIOZdx38GmCDxcqfPA7OAdJ3KNLknOcRgQ5iENlvxNg1pTaTsqma6AWTPrVoh6C7oW
ZVNk6RvIUsexZ/Cn9h5/t7YTCrZjSWQVB1wd+V79hTE2yLWMpGxVp8vUvqq6kGM7Pzw7oMgmyH8v
kBSaQG8n0BzfU6BwB/Nq2EhuDlG+saNRpswuOslIybMUvQZs7gqpsFrP73p0uizHx3kXtd+MkMRV
Xzh9laTV+QVNO1BmHvbco8ly+7HJZUYundQo0FrW3wPdoqkbw1vslWUqOZe7c/8J9yzJihTADMat
nw2FPtBuq7uCSwaFfmYPNwaJ5WFz7hIUi1eC22Xk3Ui2jV9tUM8kf67xwPmcbUYwxBC8NpQI5hT3
NTfwGWROKz4LelQFVZkR+xZ3BZTfSBLas2kEsbZScZUeMit0ylHNpc5h78p9yYN8japguuBbZCxO
YirhPGXs2/F5PiSPYXCQ0wsUVmTzi8O5eXb1v2gNFAWANveLo90h+bQPbVDbBwRO0SIb6LIjTzqo
dRRpBn2/8D5jMZq2+EEvxBFbwTOtdIPZ6o34HWSsgr6VQPThzQajjGHTE13hEO0gFTEwTZvxcXLF
qZKnKwK20odLdiZYUNUw5TgFVRJlFygQwvbs2Nafv84zKjAlOeXQB5LXSbp1SnTncOS3mmbvV2dC
6Kh4hJnQxxPRrzzGw3/q7frPiE0wtWA/C065VwIKQVAILcv0A9KtjG2YiKPQjVdvdt7gtq8Soaew
CDARkC6N9eHOsZ6x7VT3tH+j79k4++M7+i2lpn/El2S2mhWTIWXdbK/cyS/n+U4e7uwRvlwsYdfU
nmlbLxAe+Zw4kEeqOk13nxltK9VFY7hao3cQk1JW1UyOQZmm9GM4pmLmxQngmfwxkcjDxDzjmGDg
Qn4gHSg2PNP3LHplZGRUNowJM7Yu23sGSx10UPBONdNAJZ860AVf/JpNXTbVnfzi1QD1bXenkn5m
nXsktrBXFYPLeAlUPRgQz6SxWCV8C+Le0C5S24KoZCpmOUElAOBUzZOP6vdAV7FpoL6dxsYkDJlV
/FSZIVnTWhjbwCJ+vBQU6Qz0E5RQj7sxtLepcKve/FzFEQ8NwoVlcmpvAVBjK4yWAFBqmWGZVXDj
uC2RaSXynk3XPnEU7wgxP7GH1Jdq0QRtRRZTijVEM2NhEG+RNIZ03R0dqNI5cshZpJPdtf87xnqP
T00v2qoRVDWBl50gSKtFFYLt56b6bDlq6lYAZVIvVl3lUyp1PFdNilKbENquyeRxxAVmuSGaoQ8q
MrujMAbDW9V51htBeeXUmfa8JS+FMKahr1Bk/++X9ZH9oIakXMrp8QZrVNpa6+Xp0zz3vASF4DTJ
39qadNCoIku/jsdd/THbZ3dXqWRnDN/r+/Mi0DGFdp8pYnkZUpGxehLzphmmCB6w0iNZlIn2P783
dUn9FctKcpALrEW2nbnfLUHsaAfeVTyO/VSMnEBXXwa40JYBeWpY4lmpjp4l/I1uJpQmGLGo2Ogq
dTVYnArtpfK7H3xhW2X/mzKqO11LuUR+JXJeT8zxWWKfPmpIih4w5SwfGHTlwlsKl5YnabT6AQ1s
Uq5xwz77KqlXH0oZUdT+IQ7BTxBmtW4m2+4nm9lyEOIOLxTfhDnAa8HRBcG1djlZR6mZ9ltGefmK
I4EEb9oCxG0Powhr5+bSC5kA0xHIqu3Fz+zPsRmkjHlZhhxuVehS+JVne7Na/ZLVQdrWcQmqRy2R
tr7q0j8LDW3/b4szlITyzrJe3Zx4gEr/lcvEr5Tx2krnSxrHPpiTb5C51DD0vKSZViA6VMs+W6ti
Vie0o4EsWk3dzGYM5YhiSsRL8yG+BkjhM2KJLOF2CFYdOso8wNM2xxDTZnanegsPdYOlSRFTNotC
sCowY3KS6OquTOT5XNE6Jh1tq4byBvzQk9D4egQxIsAUxNMTkUQVKhAKIMTGNZcLqBZSpf9HxhUV
B3dX19+ipJ12ETkzafG7smzKTmoHOHBNgCGTHW/9Shw3hPCkXz4+z/P24doeFjIMTrMAHmbHjbIH
NGygBlY8K8b6QYhR6LPKkBMcQXo49Bb4l2EVSBJxtHmOV2XTRVMwtjbS1I1PenzJh2MbNYGTfESU
QEOBoUrFOjENbAkveRjVuVVTbwpAd2DgOa54K95vAQ6on1OLI2kzDQIgGQDuJ7IyqZSy+5aiCJAN
FIdlxKlGWOz5wvwFDCINwmOR5r23lT/fW2W+QQU2kQH/w3BMX4IKaWggOVyrTDr9S+ENvhovmcrK
dZTHGmFTjngVJAwio7dclo9qbNVtiYLZdaX+2Jv4ImbSl+xVNq7vg2SnP6oS3/UMdciyGrvxGnPi
v06YdYpmyLKKSWslIzLu9OfA7uwed2PMAsItkvJ14aSYT3OESo36GhLHWBBozVP/vR/8Nx5xTLFh
Oiyf1fyzKKOYu6fplUEqABmtKQeOjLNiu4hGBWCST4wDOowv+datEb1XKNq9ESnNrRl1UtGBpHsq
5sE3XE7oHJwvz38jzm7PLx+4zQoNXQe8+HCcWpkQwRZBaE1Z+ohGe9/dSFFyPV5lA6XhwIMfRL3A
R34ee0RsSGE2Y65zQvgvvuf5pK4RuX8bVEVeu1/XIc2zxxeHMwsT1BsynWu6XVtiAFdtIULGipf8
Ask/aB7Id64CKAb1d+dcIo2kVGYH+QIM/NyUtFtN7gY3gvjduP7N4dL1tjjcpul27xGV/0eoYTll
S1nTLGBy/Ha/P53G+XYx36bz1IaiBRh1pba3ddp7rlPLECdVlxTfsN23yyKHcC6YIEU8K3HL39Ln
/Lb3skPhgh/EEygzSVaGSHqrJRxeUc1Fip9N2zxpKwH+2r9SYxwNN9Q7UizA12HoHUmPOQCzFaPA
miSPnLXjnGILjkFg9OoP5O+DJnG7oguXlGVLUlpNV8toXvhwat8AQNb0shC+8C6UEfR2/62zVVGI
NqhjIthnLZMNJiLA+Uiyq3LCBaowV0UxbV5P7Zro4i+5q+5OBeB62eHnSTN+89IGBMSO3e1bA2cA
AU8pHNGBNQ/J4t2ct3UHjtB4H4x4OWOQbv4re74vT8H6zcxS/5iNYlyXqYR01F62u44SLqT62WEZ
zJfQc+iz06z0k9ufaiAzET9sM5NiJP77zxqnuYpLWacuUZvPeSIrsJZJZAkFr6rrVQwbL8R4OrSe
8VRqQO4049rqGvRH7OA7CXepsfD1HeHUC/QqjlfGac6BPV7uNKBD7M34h0/pvq4TUcWQq99MgMCA
UubJ3xnzcV+2xDb2B/Vberhu3as7iZAEdN9HzINishGtwjQIKQOcTNWP9MsY+VCuNLWjNue/Abro
12zsJdeJ1GJ4hP1CMULJLLTjZdVGYzrgZYuUxxB5n1qDfH9KHf808LJM06VgH0wxXe+PQho/CMVK
RvXwuLl2fA7I/mHnwQ5noMfxjqMXJJ+qjAC2h9y38EDd+J410I/kZl/QmTLk4X/umt0j6En+rTK3
xxYYK4JU+PzsbAgseAFWzyHiigQNh/1ySsE2psqvuQeFFYfyB5f11CJHXCpyK3ScBy1RbaOzt5u0
P3gcBaEP10YrVzzxobNZdeQJxCn9sT/sIkxNzsLLuIdOkCBzJx90agNbZOTXEiNLmvtOwIbJLLW2
1Y5ibNYH4jnvZs+6ftn7D0Ewm//j3xTpjUqnVlNbUbWqZbyB1X7Qc2l2kRfbVzZN5LDuuPsY9pFH
/RlfZ6TUKC49aSvoweDZe7YuKMQN1cX+Ov1IEuhJWU19esoyPBpByXTzkvzY5ifIsr+u9WWhSzYH
ya9Uo84DxYDTYoExKX+4tumBNfeSg5OJ9CejWE81W2+LQbYZAy4ATRR8Q1GlwApBsJKCxgZne8Xl
FuvBnWXxjRSIt95vARLGNbfA5CuLSCwmy00hKDRA5It8DP/R0KKXil9uAtEKtgrQannXNKe2oqkG
Q1n2gVLLIOZBOi6zCQPNW7JJ4/G42unI8UsjyT4sbrnDZ0GrxLxn4p62ZDDQlXJHr6R1vVq75eE+
cisTeCZzVgFPz4n9VIM9X925wxQ+D006J5v5uzCBAhwfTsi17MsGVPHi2nm16mGXGOJDtzsWPyDo
IBf9MW+0fLAlFgWDdi6ZCEKQLL3hdz1SaMdO0k5EJHr+n8NM/QUAc7Ddpay6YYfFW4TBMA9Hzu7v
YlQJ8pSyeuLc7kqZDrHTBHlEWoqKDJQc3BSsLGAS+z2U0SZnsGZIlHl+2kiPgU7vHqsNfxFObcRx
iCIZan7BW2mTpFrr6HoJCPKbjqBJLeaKpxH1uvwwMsL8W4IsmJ3zjZ9lkasltTtFtQQGCa9KxaW6
VtddetoI/tyw1fuNR00EfanogClYuifJ3RlF/ZFjZ1OBFOaUC7UCfSA3X8FEv2G3EWgMRNrgUEX0
MmNxK48V/ubPCGGPNmqy0FDy4jM0EYU+y9zrkDvycRceYT/kvNSPc4S2FfE0sXq+FgWsesCpdvfD
b936gnCBLQFkRS1gmUL8h/dIdurLNB6FyKnKP8ajMSYT2d/FtSU4TpMjvh8zhcS2f0THOFWbsPuD
51WPNThbteYsytQq8Lv4yni2RVo4RIA/v1vF2At0s6cZ4v3gS1Y6clYL5RC0NP7FKoJ4J6zMRa/g
D24A2mdKmjSRdG8wy6c7yegNpb4hnv6eq/QpaZOEKNzsWO8FJOYxwFlLYaPOPPW3yrX3oNQ1sMva
TNVpZW0wUaFBI3bU2i9GRxA9OvvHH1MgwjIJRLpqq6Su/cXkB5smWN45wOz6mIUOfXolQsHogHuy
SpAjTBWK7UJOhrU2KVmBy8IHxuLhk91Jy/agT7wWaBWc6wK0EhedkNu9Zjn8xvsp+gN+I1SGZkB3
C2l3ZkKn0gidNVLaUTBdnXW50Gwbar0qJlyUU1XUC4ywR3m7MAgHOFmHCKWkY4/ctIzlIe0frXWE
nZq3Ung7kA0X08lahEgaisG/D5qiWaFQJE9TeuN9YefO7gFXhIyB3NNwyzeeuhanNHwwEpp8zhSG
FnsZmLr8bTLmxnUnIRlF6SQ++l4RyIvwFL0PBT2RAIedkIYark4hc3TVlPPoQLuM5BAqa+D9gVSD
/jgIlIKSgVa2wP2XAcnxIUowE8a2XPNEgoEjip+skz8Nz9XTIhH8YG6I8LQUrGCTTZrM7OKBOpCT
c3fHrEHLLRZAy8uqViX6bPM7bKCS/U41thFLUIDKBAx1oadqQgSGlc5bA7AzIl6Un8/kbSeEP4TK
pZgiTNGj1RANFTZSR0WewLukvlzX3Jn/NOEst1cC0oLFthyu30PrNolhwcpP/XIfdpJnhN4aAers
tqzMxjDWHPPlTO1fRBpRj+MsxuBdgRG1XcDAJXxcsdUSCRhNzD5sYwRlTf05V8LJh7/kPn7rJ3gN
iNpTd5XJFhSpuG3QADjocR26dI6JWYPPtRST51ZyUzaBNQIj8DhON+6DsONZC71R1VppAyQXZ7pm
9CdjWObXOi7cWWsBJb7EoDdzRffj0aLDDQLWINJtFJlUMubg6+VdPNAvPTF7dRIlsb879mhq59fc
I5KLdkjPJqxXnkEX2G4m1gYUXiGqarJYM+51lJ12URiUpUAgxz9ouTx4yFEGe5eCIdaDh0G5Ztem
DRjMlPZ8zTmQLcwVFoRL9eg4q1/U+ag2qHed52M1zIML/H37gI+3zYI19zLo7tpTvCuIeQ5kJ+gi
rY24UHxEpA4vkmOQycbgJymm6u/Wx5PRPSyt8jY9GRmIte1s0gjFb5CG83WIjKyt1xYXxtV5z/7b
HjR3jDmbQCstwcJud01FGeRZnKxWcOJ1Rtxojas2LWy7kvRasPYJu5rIbstGJZfxcr7uW6KSs+g0
ZEFfdPG0NgYMK57dFKKL4eKy2xVx1dL/ev9q3GhH6YvC7lGLR3+Mg4VlqyIKvysfwHPwkN6QHK5a
HsHUumeoVtmtutP+Q7KRy876myF9zyd4HN5kgvIe5Et8DkSyXXnI00IjA5irgg79J9ccySTYzrED
eBf18v6DKvnvgttZZ40aoQa8RrOvYk/jcfloFEqCqzvXdsM4085q4u2RT8u5yPyRgDg+Ew9Nm725
ZO4E9Gds7oauLNNnFHH2JFIrjWyJonr+MEG2PHxFxu8WNonSifLShBOxLlxpGpui/Ny+b0xbaG7U
j2ki1iFxNIf/58jVQKUrHnc8nTchgkYDrS4Uyq32Inpzvm9ZxJdndAkHXWo6jMmYLa80lBCcPOA4
hvURQ0A4xfunXzCx+BrnMiyr7lnaERiLxkmR9YWzuD35PRw7HaAVof1hY05qo02lhhYrCYcWtxKm
dCsDZz+2zbEX2ZmSthVOwjWd6cCGZ0+pIFbTIZOyQjOw+e30GfKBeQ5GDRfE+bVYudSMNG5PuW1v
0vuPsGMfRwNwvREll76beKqvhNogv8FWccYcrW3wiaLbY+upGrMHfwm0F2/xFn65Y2XzJ4Bg2AG+
PD94mOWmTuNd9s/RwvAsC6CW4JZTPCYn0/C+ammBOreKRpIramEC+j8d/BY2K05HhswDnxu1uQSE
MiMha/UaK+pYzc8/GSMlFMsFh6dMuaHEXQTaClGUppHDKdxCUXr+ShE1C0Zw1bR6HisGMHwv3dZS
LM1kEoMbQwY2pNCFpb5U3LxV3G4hEgI5N/6mDiBonGPC2y2Upyu1PkLHnAn2XKPPPHZWSUq7cOB1
tVdNENtBb93jFnC4vNGqg6sbXqLB5EzgSz2oQD/M02WGsB6choaRdRKxZqMp3LwNqax1E/rPpSzx
vdPdEytM8b1bf17NZv4h/5bQCUrfyFTKIWk3P2J/DY8acO8f2hjrr2A/EsrLsNiOZsO4SU19ddJp
64BiAGkqhOGOhfpze24vXksuNasVzCgve4iTVV3NaBqn1NuqhRl1ImagCHB2UOTCN2dxSZ/Wuf/j
Uo0Xm4FvhJjbP5H65/wc8xhxeyVmvue/+T5Q++vr5tPlQw/XIlBRtGOjExWuA6qSSYxxBGQAOlSf
xOET8FljP4AcOvRshA6uKQh/ak29a9D0EF3Yk21M4K4hTF29H6pD0tfD8zriA5NRMj+XNhuRVjHO
uxghkpUkB4+bk4l7ONtlcbUAGSLBNvQjF4cISzoPX2PrHWu2h29BgsTPhe+LdxqlGP09ARASnRA3
8QTwln9lnntkD3pchEk0duMGuoJkNA7fKJmQaJ5cfOHP8dG7IrwC4HpV8MIyTq9M/fJLhEGf6QVi
4/7Li+F5YacoZJLesnxyRgCM5QT9SNzbVaB++LBfR1Y/e+yA4ygDF7myKd8Ykvm2bMj6z9OlO40j
Ee8JmfNnxX48xsXwXMFY2nVGK9sfq2dvGc8sFLo1jwcs1ZP2f1ao9I/PWIvKXHiyUWeAdnuxVPLv
h0GB95sZArv2ewOJpabxJvJ4UwwbriASEVBO7bGCKD3+sXEc1jdem8ZBFsXcD8ztLNSNm3p9Ej7f
KEyhpD1w9u3iMekfL+w9wTUT9aXAV1lg9lmlIVD8CE+FWc1uzPUHtk0h+BpUWgtd8hm5Zjxd75Rq
xZNzqKa6jrGEY12zWBalMFZa+qDxijntUYvToMSVQJXVkXq5kl19PyumEvAntwRQPjg76tjx9Jod
A96wSLrWsBjOFwIXE8fv4HtQgsjzJ97kHMruUPCzuSC5YPONkDI5n1xOgNxmZMHCSPknozS3l3ns
knWjUaZG3Mg5S/gszwL/ZF0MoWooBQtSqx76sDhJeuOfhyzBPdRlH2aIvg+YqblrhlU9T9t+hN64
nM/UBd/772L8y14+7QAS66KH8oyYnljO/WXWxRaxePhLJT26vLOkrCjRFQPFL59Nr0sndjo9jxSC
jC5b0GmX4yfk88n3Lqho+bnH4DPOacgSQKiaMzc1AlktfazF8GVBn3xFhRJU5X94TkqzfXXpjHhl
bB0CmqRz9BZl86Jg28QStQQlN8ZQ0qAlirDnxQJTXoFpyh64ec9/VRLXtXMDzamsBzWRrD/K1rFG
6LSmuCfI3zexcs0ztf618tc2bdB89IsSncHVgv8AKgmHgup2JZpQUXGDhHpOv9eTXz/lHack7bbV
YX76k5715XdS/WJcII+xJcHxLayj+FzDsV8Kp9inW7LTPMRLgo7p5CePQPi7UEqwbYquEChOKM2F
AwezLvdpogBT6E882cp3mKXzQtOtyos/VAOhjy7z3NQB250iCYr2YFWFUcWfWGlL3JAfnp4yQQZu
rnamZzuKSStN8A8Iy+xlc5i2JVmGE7W5xSaa0ENpp1qLqP+Ok1eAqkA5LQbr4minrSfKkDn1xV92
6/CTnTc2Z1K6RgwwOSw1k3nnJyMNWrrVaqZGyyKQ8e5z2JjVH3uwAqPJ4BHY7bPr3Sqy+JAE+eyZ
+XjCd8DHsWxobakwSAMbdL2ZxUa8Oxs2xUui00K2FNZNmEUvYzZpehy2Jv2tHPjef2kYd4KuVBqI
KP1YSiMOz5AI67sekkj5msnRkPD9hMs9xORsHNoeMKXz75kFUkli/e2Drq08k6BSodVX9KEIZHKd
WBY12Gi8LZMPsvjqKrplRmz+ZxwyoOstRUNWLPI43qhOnSchYQo1vhkRP2Hk0VmeTM9nNUgzRcl4
LQBi1XHgrh9TAtmwlX/kOl+4HFTl/V6Iv4gk8kjQuoclwaBgd9XmOf5XXsklTG836I40NGC9kqlb
BN9TtUrf2N6K9Cb6iILCBfnXOuIzaoz/2kVzBGRIwzcZV3rLk30t5akyigzMi9qRhZDpMtewOwzf
1dJFXvltSWb5FPhYKUPD181vhxNxAmzKSoUro0ifQiaXTS+SrJWOC39T4ZUSbdSUl9UZ6LtyRq1k
Xd2ADtwqmn5sUw0G4yr8m9yn2+h3/KcAZEgtsle0p+2PpSmXYByn369xYBCLOqutjKsm1okCpd6E
BPJsojQvwVBLOZpcITc7Sz/Biy49n4YfPDfkknR1ZkbbcBbaD8kuK2I5coP61O0MJHdAaHJpVbe/
SECkASn4Z5161QhkvU4EkPECZjPnTjGNvtJrMnfOKdhI4XAIlGyzqVcLLi8DMRyzRKRxUEGB+Bz9
zcnbr1NAmkP+FtHXr6QzHIIBwwnOc8F+Z+BqZKzRpQktvj//OcntwRpDvOSAhKqKc5Frc8mhp7df
uMuWc/qF81X3BqJtb/DAACDCUsMdKXVT8mKQn4IWD3XWLUg2zqYLpLeN0Y51vlC0gBXTQaYjzk1+
hgYPpindIrJ8Q1FxEBm2fsbANK4MlP/C9lQlX06Ji0/rbTEND8Qp2N1s1GZWsk7yC415zYD5V8DN
w3q6zQNep9MTiKnjcsRpBy4b48uaVUJoG0cp8F9orWlt5Npfncsli0tRRvLjXz6fwHD66HVpt8I1
90EUkqzIw1Fow9i3HP/QFZD/RxYQBZA4roKvh/Fg2vwQBjbNMvEbuHx6z2WphDNbZvx+OC22F7vS
3j9ObmUPhbP+UAEVGYLwQGpOyT20AKLrH9oPX8LcTjMlVJdN1/PrHafs6Ih3lCoL6V+MA2Q98ovg
VIR47wok3MU9THPqp76Dy/rWeOu3aCRw3igbusIiW276k+XxHg7JwOADfW50kF9rngyaZUWdvxjy
UMEz2wke870NAT0L+Mamg+ZVIfd1451LsyvOL2mpF4bmzMojdloskbXPRr901N/GFw1j3SkXTOWA
s70yKcA2vu/NRB5MeP0jQ/9maErtxacrQb84csnMDc83ymZ71vbRz0Iw8p2SN0QhdoVJBX1+7eUx
aJoAXoP4LcMvxsaUEI9K5/GdySv1eGJeIQT7gI6LSHFWiUL+GgjfwF8kYWxedIEnRFaY2GF9fo7h
SE21U5falicDqohTakglU6OSxislTdWuJWJX/4YMHmyEBGyreyhl0ueq4jKYkorcddK5725AkRCn
I396lEAQ9aN3pJ7DnrEqcFrdg7oOwuT6UuOoZ81/K/QFpW7IeGBh2pG1mY9YJSUI2RyYadNweA91
IdfveX2N6QlKwx5qmriRnry2xHrVE2BweMITrhzxjOgsu1lxhxym3e78y7hC2bbs3ePxMHtvzULD
C2nUCwkxKU+m+o5JOEP6J3Vny1CTji6ia4joWbGPrSP0mHt3JB3BITN5p9qBskIkOUBq58eeGQhH
o8tlfkv3Ohlm2dbIX4ep+pt8Q/VXByRXezxee6ycrV4UzQnSSPSOMYPbkSypZx8vgvKNhmeu03Pq
yzimoAiDBuqH91KIMkUPStmkintBu7vPGoobJwf47xzH7aBvhZoZbrsfjyVchOS+0Nag/OgP26qf
jltsrMN29hhhmgbbhLrYwQdlpfgc5mz6q0wJAEjHoPl8j2s9QfKgWFci6EzEfSPRk0+LV6x3ynpx
+eQuNTKK+gjwflj+/PsvVJ5pCLwchn3bxkii13x9QGpk66Yvd8Xk/Vf+BqHw03Y7+K1SZeAvSY2A
sPOtHVfkMBE7pcTjQnP0gIf/R86WZ2dAbosZNmLD26I/8X4zXXlqEbJAljncHWaUvMq/ldoDCh6I
aBgxvo/M9+A3xjooLRnmzfzClxDjiXTk5yTlr/GWWKY1hB28LR2pDTQmiCq9WhYvU7Wl032ourbM
ObF03RiTYaGJfKP4MXKO1YDzcWh1TwaNDEYPTbL5jS4MMh/ssvd1AsZjI6E8+gxSHryFQLV55S4f
onKVXpncvp/Ge2CaejFjaZHJaoGp5bzWssr6U+/aUazk8tzI/hGm+s1qIwUGvsuyF2Qak49hFZek
SsKyaLZ6VeC2vBFkso6c/Ei5UjtKcGbzBEwIgHP3mrz63/juiJliBged+oKpLqgX+pb4aC74kCrr
X0KG3LXwL3wBuC0zV+SvRvkXlhovm0Z5zWhZu+IrWMHb1R4JsA2SK/4oXrOU4TIOSopC9KMIy8fq
hF5877kGDGK27wBCQtfnyypUBzy/ciqYvaB42h/ypqlAjFJ85H/18WlgKGPrZsE9+TAQnDWIPPPh
fp7a5z+LwUUKmUsBG58IJcgZ50GJRvtuHc+QgZb9bwWDtda2IWSUORiC4+v91RUL4Kn+D77VRow2
FCPzVEpuDwKTNKA2DwDPA9rkmcBcWqyUcHVTJDdY8d6rMfr6KTyIIycHJCaFzEOP0A+T0oSvZRuA
jAJPckTCvVUlypuDgI+ey/iUpfagrn+dPVaeaZdmbSJm3tdPCSqbp/gvNaPJ7mvOnHGUeBV0U+1J
GZbnDtpbDRYIVo7pkaig8DPAO4Zyky5ZPybrsWHJ1rGmisyDcLnksQe2ZDsqD9n1Ir0+TreTqXvT
Bs41hccPolYvdN46g0Kqd8ARR5+SsgBv7OWW9JPZG7WdtHhhDSkurSSQKDuWrl1sELXENq1H39nC
5HCowm8WIcIOZ4FtG9h3eh7RoVwujL3U/L/kDnB1dTyS1iTv5SZQB6NcN1fgHpoU4QxSwuPJEiwT
6zxBMwAACUHQkxuSf8nZcafF+DTebkNQFVXWdd5ziU9Q51UaLCYUbnTWjtDNcy2l+mkmnZQotGbL
Cq6QzVtN5DF6uFbVXYdOxHr4M3W4bsMnAwwtGqKJteqhr57irGL7lf1SMVH7Xicm59dNppmov8ok
SiepqOyUI5UfdIRDcHocDw03Y4YYUKO7ghu6IpYoFnLPLkSfBKsKhOpbNGw8ZBZ5gPcUca1fXeTA
UN7Afm7+nZc+K4BYLQYdXkhaUvxlzXSH+ePxolGbV7TP9wn4djBgdS8uQjX4ejjVEdavIS6mNH3h
BdPvh3+HdI62y0+QH75ujGEGilW4JlZiPN05Z+WB0cOX/UmzyN9v5L22i2gqGAcPHxrQV8Y9PC+M
NiXeYJRkwCIZggcnohpRufVDab3VBfqB0eOPlxoZZQsneGy5otHWQ4NH6FyNUUQdQU1W0IDGbyro
aaU9g5/R0CKdSxWo/DRIaT9Li31/AF18oIYd27uPofqbKFd6CyjBao0fRAfFHHuoS4kRhiWpw3YU
BiydkRiheasO3qMHslc1wRtag0jG8jeuqw6FRVoKgvZtOSBiOZmq3AXZsbKf3f9iCIyFoFKZ5yrJ
43SfWY4dbpl9iy6dephqqqNRZPP56jqWt0HkmOLRuRBobQoWa0/irli+e0ADl5qsMNkAkkle5g+7
ch6+ICmz1Fu5gmQDGhbB6O5JR4GcG+EhJcZ1kQMrcmm/hRh91Ks/bAVRKC+/HX38caD6ZkASGZKM
8BL+1z9oqf+9JEAl21+WtnBVBa85EboFsFf9ggKXUiZPnNsvmdeTG0VQyHFW0REtPX68OYA5NFj0
lunhOY5o+iXbEMowsfhS9fqhAf/uo32STBPykSX+/443QBgzsJ45KKkL1MT/w6M8mq5VyjJujQC7
E9DMzEySO5MfpHsA+K7rlYWoneOo1U1Xrh2h7U55udKpHeYmDIcCMHmO+9fFd38hPf3YPN5avHDI
Gms27D8z2hMakU9SoCH+AEyXo7GTf8f7xSTLgItjNr3oB3lL5FL9av4YxE2GJoYdbGfaeJq3vh8f
cHI0/dedVkmTGfzdaVSm6i2+cBvwxosK2ToPtgqIPPVu2mQQRNFxc4Sf7Wlu6q5RGDSXsC+mR1fD
B12SKfZL4adLJzEY+pIUhzMxquR6xGSaKi9HTCVBmOxey870OzKuSrPl0bRrz/VQF1LYmHEquVR+
HoYGW97MbL+viiWxk2NwYK8V6NsgyQCUSrkpp8h4L6hDVDh4PdBBKosQtoDgwbslN1JhBF8Kw6sU
M+qGzJNGzpwAPurhSmm7w0w5q8Xwv4zx0RgIzDImg4w8sPu5wk9fY6cIWu/avm2Muf69w0YmYUZ5
3J+EUSV0ic9NVbENeUiF6ILQQBLm3ZVVq5OpBRU86pwaYzpdppC9Wrypesc7EBiT9g/F199oYEfn
9gNtGeUoTdsn6c2pU14Zx3EHto8SlpTT0/GIf7kGlCSZB31/k1hyOSfsvwwDsOL3cAcTXVqlJ+Mi
YJde411kqTHbqrUxOj7gCO78RDWFhOvVZZpGRjF7JuvtzhjldPt5fiXBqNTRslXSqWWXVzxQUEM7
TvwciHFpuiafoD73eJwKZzn0kf2mG5SunhEwfT70glExb3eJOjpchd84FWJO+4ufwCL4ViTrwbJQ
W7r/FLIvn0knMEbsIArteBMtxU4zJHFj0RaahOxz/Y8Ykb0FQuBt4wGccdYzrjI7MqW52jcRgNJM
XC9AYD1Q4osZZHJ3dJHg8uU2QA9cKK/tfnIn4jYUVWnFylrBuxnFV+Ux70sz+JiRfC8V/x5GaNOT
2GBcUgWZaevGlVU+EFlvxXyr5NhJ63TPhOX/T0Mu3XH7PM60ekjHM4nTGNsTBO2BypdnY6CuMxee
2E5cybQSZ/y7h1L/FjwEC+QQZj9O9okmPC5+luCwX1RqxS86xaX3JDAi/lVs1tMIVtWhLtHfMjxF
QHlgZp30baJjAvQpmt+6UGGqOfoQ/NygpRXlokC2C1WIKG+frCdOdtnCvuHsl1dOFJjjGzZ165il
wiXNc53k6pbFEO3N1pcDInXsOKFYq/6KPTGq6SZVIy+OBC5dQrwn6yxVxigVfYGbu9u2ecPcFmgd
exYdwblmtWBq1acA5jLNV9pvewphEX0uMiQM2XLlu19MvREhnS+i8rzbs7qkPeUOHsVxTClJATQG
fp1R5sm7mCkaEzeF3CP1Lx3j8nuTY795YBtLkBQ3iw6VtKDMdvjkKSDaA67oUUy8MeVVK6oEmvC0
KDvPkpQ3tQF4IR4xCMZFmOQyevTDnbkKDgt8w4PrCcWM7FB0OyknixmwY8uIn9fjoTwFFCjqysf4
Yzwpt5ImEStAHfRxgU59zYVc3PROLY0T+Mmwiinqd3c/jgTTl4oyp3Iyt0E8g0R4IxGsb/SorwtW
22de1XdZEFIXElnr4QMGHESWkMDNNc+ieehWv21lobB6dvedYoKnMO6f5K7JArtfAnJsGcDixoCt
ImlsrY8qSD3mZrGFYCbES5PqnT/pLVOF9ydicVUl+FcaUFAWMU/iAmefE+ckuFq1HEcN+pmonAAy
LvdXzbQ3FRqpJH4tExrmWApAYFzEVCDN42YOdDQ2D5zn7EHsROR3/NtKkl+HUXnfd4vHZLl5t60k
UmMwLSLxgJDLGEgf2r/o/tH3GV9zldseNOw7rQGHwrKjhjEYIVv8Vl3Z9ttFOb/XLyMWHr4/QSK3
I9p20S+z/rwbS1S8fHjDt6GaQWnF4tUNeqGDIpTMYlESDklIMvE8+RHInNzKTuGtBdlXwSdghYfm
oGqdNMFRon5adGI8+7iyPUC2o38EKQ9JxKlq24WyltejG+WcXyfvu/DJvQIMvAQBpOBTMIXsYX0o
g5uHmfBF+LGsDCL6rcR6NjSVQIcDqG7QjUyiq3lZG5mJH7rFRpidUKhf+rTWIstP9qcK+hgJvs3A
2BbXyEQSeeyFxOTSKXn5BilPxoudCgV62XucH26vXK3rAN1wsE8zzXJ1YtHJ6hhMM4qbvRIqgElf
A8pFcMcjqXusF1peH/d+URgE57JnF0WWp15nUWHExXqVZuOQV9U83jcqxgi0qCLTB+EjmhKRgn8W
+ZeMKH75HztdWw3qcL5nqJfcyfDO5grO/uVJDGtbw8gaPMeAm52DyCML7wOuWYHBbqOQXdBk6Yzm
GbhXnIEm/E7qnaNSdGmdSEFrOWwpHWKhvHvjnUDLtvUXEH/Iog53NMCxrZ9JQIAjRLBxu9lJTTZ5
yTLiXIBzpMCuufzDZvIYfHswgyNWFCBsSut3GOGw2ecb4aqVhFL8+K/ua/46Zpv9l4b1hlqFkij2
EtaJgHsguBkoC0hesDiwcER07Aqv7xUpEHDJIdWorjpC1Px7rMEHPpoI1+9vRNVpnajFKNSuBp2T
rZUpe7vjLOcd2eqqLd6lv5Cmt+4Hm19WpmKxLSbYBuyeboVIrISn4IsuzLpvjtY65HXgDOYv7HTM
/2geTRp50yaohh7mPQ3FDYUamg0l0d2YYaUkP3tQ3VeePwfrQ3AjEqfGluEqbTtdEkk0JXYBoCW+
WKOeNAHUi094gmpbGp+oLmcKdN3m4kJZTLN4YklxMwrkwAAnNC7ARq/TPVLnfjRwN8Hv0T+eDcWB
8RUl4A/jgcFtNGcEOX4v1uGrCQ2HLMPxxF14iAvB/QUit3xRKW1UYdMKApO5rT7gTPphVmXbW9ML
N3XqoJBpYIVN2IB3QSsithiJzC6vpBTaysM5bM2i8jtzlZfaH8qTxr8gdzPBxcYm0FKhBpeKggMg
4s7KmEI+5K/E9T6cv6H40msXkzcA8D77aHJcDCjVoP6pOYMKuFe5sS00HPhumPvMnQytQXiNNewE
cc61W4VL3gKcfbfwcJKMudf7c4rDj2WBS/0SVTZY380C2tc+B9eQ+I7z3xXZiJZxx0N8TyWHtnFV
Q3ByC2DxCFRXXpb2B3o3VvCWsZzeiT32LVTjZzqmTARfVf/EjsccDTzAxYctpIZjd1v019Alk3Us
ZLzLWm5iW4sQsmBAwzMMIU0QRRJJRr3u1xOVBWBgumU4YM6O0bWBR3+BnTV9jFU3ssYpZ5tG5xUl
hYxl9MBXvppSoOj/r77SfwWEPcPKsNtuNcCiHPcyg7FTtn/VCgVedsVcR6gVN3h+9mWu5wNfMo/r
Y+MYSFV2zwberQ9Mu+qBhfTyhCdvq2NdOJ0NhQ4ar/RtBnY/8pQaG0h3JigogScctOo7U0ymu6ek
FYStlyr9RAAbi2xMUZjXnyQBYH1ZbvNETQ9+JxrP4mZpXyrs9bhoHKkokOgsuFM12CURG600OJ1n
ClHzNPHSuP+qPQzL7G2zdSMOPKiAwR9q+4zolGm3ojVaDmjYbITaSQR2Cnaot+oNMbcWSciq0JrJ
jkawxekgIZnua/BDXh8E0/sUfbydxSVRA3S2e/MU/ZmMrevqL8tLgXCsEc1WI06fJGmEeRqZ240w
JgF7bgJPhJIerSQPGyptN7CSKyTN57dGON5dZXf5Veh6HEV5wcjHv9CEn5GWxAs5jFO9abhojrj1
GrAKDrSS40W59VNqCUYhA4iuW3OTSTwnX9pQMyLkgZOqSCXtQQssq0jIniSQo6MlJPck6h0Qx3bG
fbnvWxZUGy+0F8QeTb87VgQAVokio2i3R5wqPAbxhby6PCmwf/JeGCmoWar2RsII1sSWLmGG41BH
hw96RDrUmdMmOswwUefBt6a3YafMVWyQi7Vsy+u+Y+N0A/JMjTG2G8eXZgOPt0up3jty0VLXRtkh
mVT/s6nAIjMaKF9CDsdwz1Xg20rwyY0lOuQkHYWK+fb3rH5ZyKVgglsgJsHrtVisY/KwP8DvdxHN
+oTpVI6HW26NeHvFvQ0GCCBKX7xD2O4Bgk5RPo38vXGBb/qFXHigJFiG9Xa3Od1U/vxIwO8IbBeE
eMlBsUZc6f9KLtSpW8dCSV8nPh9XhLg0k4mqFwzpzB4EVld5MIwQtks/n2G7c3l5AzwIN6+0eb0X
VsbGi8bQfHNKilVtu63anGriu2D9EA7Yd7TSISIXYeT562bifNwwpssWeknc/DUyq0yPoUr1rF9b
h0ykbJwcuIUgLFn/c5R2fKngpPwOOXFHU38o6baVsCSfQgwoqe/rpthRktqlRQNJgLkTLZotvAbK
Ln1cSJ/k6r3YFjqwO2x/3I4e6XZEiLxyShRKzoZVSBKKCKpe+Oh02n+o2jTtNlmc6ZUMtUj14/0r
4JNg/uqVHvExG92lz8FYYJdGuSjQa60udVezL6FRK02C0IOJyXlUpY+hrvjjIA7d6xfUu7xwDEKc
jFMf8UzvG0IHtql3vMeP5i3zJPSRgcjT92fdDTcxhqsf4+U5ZmefZSmPxWsf530xqWRAF6CgBpXx
TKAIbxxxS01nvNzSVVcVihk47UF36v6MG4AVlRcI1eMMUJWRGQBXqxWLCev8tydWOK8CSXKSINWO
BxKhgEH34LYzBlqoc24mlmfrnAbJ2aO2CSiPWsHwpUsuNmsu67yf8NoCpQXHbGNS/MZLcbG+rmZD
jDmAo/N6UldLOjN/i05hhM22yoQ6E5+g/RV30uXAruHthPBr0YXuLp38aywqI+UIY2DBfV03A09r
EFtavskKtOdyJDwp7vmELUit+K449hL3zUksBdKjrYg71mftDUVd5STReE2FztFIFYpDYz3bNwUH
8bNilfuhplaa3pPLDXJLYeno1IBaTfkxnLWDuoJsu6F3YZDuvzCdrnpA/UkysmzMc+GsDEBcoGbi
e5CfyLPGx3pcY9SybOaK61QqsQJ3orFveil5WwtPaQVnrx4xPp2q/W15JThgK28817FhI4VS2SsL
+NJiOJA8WvB1s1TI6PPk6uWZzC1ig7e7chUSa5KFJuS+DPXiWlpVs+AESnQp87eLS0EJYHnMDSEr
svFmYRCSwnn1+yfUpIz6zfumDp1BNo6ee2vnplj2diMgmwaQ0pOccVsRxnyi63uaOQtcRORPT12x
ANzRVokds+9mKNTsY1jqLKuCptRLzYI0xESmNa8yFxBwpiyzm/o6wD9GDjyM8Fnu9WHWQhZ3uZZF
BA1qd5U24l8ljKh+/4M05BvMBiPEqy2c/WQ22vEPxAwAT3mnm5sPBR8OiR8nHmJsMqjXgmrzKzwv
MDTEhRURNMfhwZmImQ/PuEst5vQmk9KoIfx7htfsU78pJQ4cLYhLEBJzW4v09lp0z7lnrbW7JCOB
uTpUlRkuU07t8IEtqb49J8jMHb10TOb6G9rNwNrMHH7BSu804AHu4GipO2cLo/E3PFunr+jWDrO4
xIl6Z4qRPSLIsRQ25+gNTIrWOBDcjYWDfwQVYxSTy4BsNFUWATxYKTAchZQB55tqJaNu7x7erFjy
4uwtmN8GDE/OEutFwm0A/E6NZxrMQGXZ9ma7ZclFUzPAKz763/kZszlz45d0Ksae1tczQakbFUY/
1o/DKyrkO057Kiz2bIRvGM5NDtjohwdjtcsFMe44Mje9bbrOThQcAfq490Q3HcCZhw4MdgOhY/ns
g1LbakZQq0MVsqehWTb6minsK3BoW5oFV2fIynb2f5vnkED/oITmdXlyFcV17fT3bZvixG/Kgaul
yyIInxAAn5+MjZJOM2I2JXMXI6mm2EHX7C2g/YkdqjYn0hqA2DOVAvw6/epatnAas18nYHh0VLBn
bFq82X/30KL4CusmbtW1+aN0DUNy10WxsV4IoYJ2X1ob5SQaJOFD+EhhZUG1GWFHGHZaMkEB8/QC
4QYeR45Tk2jbjlnv9IAldvPmAFKwl4CIZNORTKO5C4VPufcL4wff4nED+PKbXPhLgiomS1ZtnR+z
HoQkoYA/LlSlXJCZmlOyyR3M07kfyQWEj3mJvwgYT6nOPJGfv4QCsVTAbmiEOj9nfFCPt7bG2Vnx
ofFtxW1dvXjyj4r453isusj8pOrO0oRq46CoeRrJH7FaX7fvrG5kpVuUs0BT1P3gx45B2fj6q40x
90Io6ZrrRoROCW3rkClqGa2bPdkmh3cGCADOPfBRcuX6xZZ2Hv8I77dfD0HZxnARQ1SVPgmbyE4B
sZsCw89upNmmlys8VAh8qwsNXyn4uMT7EtX2UPieQZ+NEq1i2gzKBvnxYuQt30zOPWznzQBhijSd
5c7kGspTkSk+yj0VIxhBQOlb55j4foU+1MCHkdMuhKnOX700gewzPj33a8ncEvmHnnqITsTN5xXL
3J6czxGyAeo1fKygg153oo2Zuf3nTIsz/mYagB2UNxVDPJg9HTBKaRY7zLFK8KjUSoP6W2tGmuwx
sR0t//XD0/A/sWu3oS3VuzkUwYtY5A3gNz4N9rIvmTQPuUoF2gkjDw9sHaWK5haSiYso67fCjVgr
FrR+eZlzsUMKTMbxbVRh7aD1mykcnvRwd/+UG/OIxmMDph3k6uGtKuqyEHjQ/pBqgge9OvLtOSHx
3Ts6+8c06IA9A8Laz+59AlhgV5QyGfySpQOc5IKYkWZ7SgCmzOV/fNJCUKwF2sZBopnQUNI0FP99
6HTc/yicb/wzYJrcPPEKauXgbvtzvdxcs7cLiz6BqmfTEpBib2rgtYxHbcplNxrBl1UzL9VPH9GF
nNyjE8SS7Tm3veDAokg4camDpcPxENadimE+hjizFjI3uNty6Q/Pd5UbXg2bXgt17j5bKH8ZxiVU
b+/RRLivN8JGixajUEATJfTGCMAv/WDJyRPN0u0AsRPwsBM7f6bEe900HK/dCzuNdkCrinnUqtIG
rPPm+HnWRlmP7/Juq6FE3qwvlVFzT21JCgAnN0VtI4Cs2Gr1AfXmOFtq5wYHugcza0bNVSiMojJ7
dfbCjOACsaMjdIMz4ZRMYQhujbSneVMTvnwJ26MDOwAXKM4lcFaatl6ndA4DgZs5ny0Rqn3gbL6M
6YVdTlCyvqgSDy7jH4GMGM4tJ0Huz+LHjJ2j+SgjjmKi9gnfnssbcgj6xcP0OW2qbU7ReojBuuln
Dvjqlr6j8PskBprUk+Q1OV6yBmfR+f7vefZvqBS7MnoiDJADiP1nAvnWqGzMwbLvejff2bWTKGrx
xetIBEkuQGSWP2yuyt9vn61nUauNoAZTwXz7mN0xh9Kuqz/5muXnmWJu0TD01zE/kOKlvPnfhSfE
w9Shut9BmrXLW+ocmFk9R7RJwZ7HMJwmMOo5FYZDWld+0KyGhfu7/JLfi5YQywot+oaqXDuw/Eg6
L5GpQFqaz/JuWdISStjcCPFNSURxGkNoy6DjBgiGtIbG6xEH0McZwhFoL8MPIey6WqJ3MK3vQm+2
gqVE0UZsZlftZZ6+Aw2Ki4BzHg0AjRk7ikVJekIWVWtOjiBlurzMs/hePMK9qX8BjZwgfU+PhhSn
U75hZEpt245CoOnMOZVZ4BGFOpB/If6FURjxMNKgh90dC/0WihA81H/GJo6k1g0owruHQz2zh2BT
ZEFjZ+W/oLlHKRyN6aScp/o1LrKZB3bibqGooFIjsEUeQOekc/nzxsHRLlYawTlRcwKXI+3UJ8Sv
Fl7Y0ehgnYohc8mZPkdNoM6EbCwp9y+dFrw2B7Ba9f5esHknz1LSJ39RgpRenn8H1nnAt8BeCtx/
F1/l7aVlysY5YyXUqVTQe8M2GIz7mKJJu+K3kug7ijI7yPq1xAcGfv2rpztJGNCNf2b9L9a1M3PF
/xWupARjqMxG6W6RlTON3D9TkqWGeQh5zlwCOK5iccl8Ge45/K1fBBzVynxJMwpXeqkmGc+8B282
g/z0atxSG1pHvO6fzDiNdW9jm/cBUFhJqY/u+8cy+F8KvYbFeBZ4PD8bbzKIFcSmP7efsPam2IU8
mhk3np67KunLoeE9aUpMMtZ56XazUQ5DkSN1f8Mp4+cdBvKtxWQkaLFcT+FfRn3nKxRi/ufYR0c6
SUzjKOsrShN4TlbLrweSdJQCQA09RLF9ORlwQhBuLZY6BM80v34BLqN7CqWmQmWUUEUz3gQAEJAa
+vM11CQlVafq8h+4Gb0ewFWtNiJZZrCIVmZ23NH0C4Ywk0cKY/hLdbpdT8+90CX76cl6MbnpI95h
UF9Nsw2XGA+jXN5UjtwLiFAWUSrckndhWa7erpIXeIazdasLN2aghyaoyyGpPChC+9QDuX+f5/Pq
ZshJb3BCRehLXle5FHs85rKcX9Bp9OCWI1V/J/YYwHFBE8vVsmpUDYyzePTI6kjecb9a5iRoQQ0E
H2eksdJrbgCYBidNUBTVm4NY+o/1a+IiYz8NEKFprYnRIxEV1SdP1PzZOY82W4cKJads9K36JeTn
GAH73YjFCK3jzr3hi289z89L5OxMTupvTTi87cUfiK+5gujDdUSRuEwHKq/6FFHr/wYQndhYeFkv
HmuC+h8Oerfl9u4uyGUUYMbhM5ET3PrtFj/JwuV/n5l1j/Y1Q/fkO4jX4BPha4/3go78CPBYN/gq
LI1QAhpohAxsn6UaItLplVej4UA5XqP7+3jAMzDGDcpqjNGttXzzta4dAtBwsH3B0vsJS/DS64Ap
NzIrWdhk3CMnuAtg0aCeKZoYlpPtUV6k2kPKNQBmpxNdxU8+I56KuFVQQfi1HdDGRufUTAI6A1pH
dHQZi0Zso2u4AJT5sixL+sDMlhGbdibEhEqpkHYU9IzqCcdJyvM45YzBknlevo440muAcaNjDXvR
hySfz6OkZulghV3BBGSnmyw6zA1xqAc0b5OVCOk9fAnk2AF1UGKASWThO9S/aoz8qeRXRZxH8lyd
Y7DEF9959DfJ5eD0/j19izqJotAN7kHR14pGYkDkBO3lPP7uph44M+TxztV6mKh0D8Ef420Vyao9
g4nN/7tIGkO/4aL9LtqMgDMEyba14bD4Tfydwl2zBETw7eV5LOcq4BffpWf7/yZUrscogq1XPPkH
GnNMJaMh/TH6LUoIfkbRVVr0kP1QCq8vM5UXSeybIbTqW69Y57Ny3KbpWC8hZ2lG7UyPppqQFKiF
Yn3wu14GoqL+pC2WgXC7wqHxioDbiGvz30ay2DnToxOqHEw+8bqKuGCzoUhcQO2DAmzcNqg5x4Zu
VtYGW1HapL0GOQhRizqQ5/BK2WesEoZaQFLGR74ExU4F0c20YZJRF8e11N8s2zwk9wzPyVctKDXc
ToCuOQmp7eLaM7bmT61E7TLbuK2lIOByS7Qohg3DSxc9zmzjxlkZPCILgzSt4FoPoOk0yHwIqmL7
Vn92PsUD5J/3+x/iExQDbNFMV3xCj5iKPvpWUb5VjBmerT3z4rIRe/ZhMVHIwbgM1+XvqhkfIRTB
uS8MEN6usXAMc6dOMNC4kk10SeWJCb0HhydYmAay6s/ichoiuKHOy3O59WpNbRyUacURJqh2pDTW
yIGoahXXbccUeYfInC3YCTXo/XSkFvpeka0cRiVxtn6066vp2xkKVu0tHyNm1cdnzA0dco2kW/3L
E/3gk3JwHpYnAPaWITlEELE9K7sLUbOsDNiUkUXAbDJr6tVuq979/P0DWQJeUhhlhwub+R+vmbPF
3Dq2WcyxSfM3T6hBNXb2tdh6TzboEL0wAyaUqnGlB130OcbBujbZqVPSAEQElwFCU2xmh3ssNjIw
n3k/LaiFnkBDZDUwToQHfmcEa+aQXSPvD4sBsEMF7cc+v/jBiC9PAVcoKqJQDv+ULYu0edx2U6p6
NQ/8NlujrI+x/obL4pVfeerYGR/+psknK9ytVn595NDLwJHYJCtMnp9J10KRIXgMUCDS0rvEtli4
o8gzY0ngElpSP2/4+NABpo3if+xbm36MU2d+386T7C6KEbqWJl9xA7O2NyOpVR3efdSz+MTUN5Vr
JUJXIa+L3lfqgLLk1JKXzvB2lu1KI9Ov+/Dy6jln956d9SLQ5WP8I9BMIrPUMxvxHgOhyG1or8/k
Z320DcXFANmbZPu1ovOxxPb6U8anlGzLCdrkQ2zkd0yCKrmtBGKKGNtlaEFasWmCo4jAlsZ+cQbA
krjr+xLLc+IYSP9e3Z50cfvJPSrjp89WT8T9J1/6yMq+ESxhLpiDLmqLezBvLF5CYl83vEnyYCBr
VyLc0whzaBMXT7eL6ahbg73dlSv9kkyjACknn+ZvAIvAExdFv4AAhkbEdxvrz9ssbWsLbAKMRcep
UeNHJ/2/LxHXRWrqZ2rMMaUkalkVFPhWj/9yVZc+Y/GdST07H03RW8GAPyl8uuFT1hATqFoXmwQj
sUwm6oAvDeVFKSFXoDYnhlfsxPKQh4AdJRPwaEh+rzezepBalLyKd9bnu0lOknkGma7GR8gE/f8U
ZZ3QyEgz4a52sikHX+8Bi/iLVrOwZ1XcgX6L9EAQLw8I5Gp7yM1ddBVLMvDqK3LVZOJcUl9x3Ht/
8qh+QvuGMh1h64bWvH5WcYHJTvJPT7yu+0saW+coVKtq97ordlAM79MuB5h/Umy76UOLMtBigp4d
p1VLxNm69hnXpXO81YY7gChr816od5d4oTYK75zwR7hgbVYyxQo4zyUmVGOlYYw/h8umVt+bnfF6
IBOpOXx6xy1XO3c7Wc0z7aNrcrQPhgYLXzl2rbkxtsqqSqr9Mext1p5nIk5VKcq4grzaYNg82rua
10HE19WST/LjXxl0K50k02MP1IazvjBDh16B/RfQY9KEutseomnTU4DFDsazUeO0EmI7w2p6fr4f
wRY634FrA08IxnlOdy5/FI4GsRZwPlGLr4U662WoCgOrIFP9kBzxnwoV67DiQ9X0NZnggBgCy+lp
9u544wptZdYAzsWsaN8qZO19ZIRAjORVcYhMKaWVR1/BQKpi1uo8DAruX5riVhcL4yjq3xeUY8dM
Ug3nJAjO8j1+mCTOe3jVC9W4bOgFearVnNqfUhN7ltuTJ48N/0jpaZay1IXr6LBnEEFyhvIeRzqk
ZBTJQgpaVNE5NOlRwDOB1QyjT1bQNm1Vz2oyrb5d87e285SroQ+gunKGJeAMeL1A9L7l2J1WujGq
zjktvc8fz1PUJoWd308i7RHUA1Ic0eS9YMxoIcgiGlFcLU75WsQYMjj1T1W34SLlTg7/4lvJ2Urx
Oe10DQeDPWvJEehecaT6BGlFj606qsKVHalOJ1VOwHvLxufKPgFoFJDfHaSWeCVzRWuZE2lJrx0w
cgAhGgTfHiCuGB0pIWmR6WCAzEql+jY5wlPOpkmyRqJiShx8uYc/MxiI+yaBSxTbxJZLVfos3YzD
lbV3vl+iw2cbUDSf+KgRVaOm3pmnHN/BlQjPwTKoXpNBXgfqEarPObM//5No1vG68rpNfX9nJQ7Q
HFW/n9B9htaqe+CwlyMtIUZQ7qbQv58SSOSR6m6qX77SnXa3RR9EDJnpkXY1FOPmQHMVPIXOLBg6
dz+lGmAp1dIXGzqFfxQnKpUcdIfuZ2hhvOiJwW0j9arw9gaHvpY7BuE0FkjlHs0kh5bMFh4/tMSX
rb26TWN6rXo86KzPpEVpy3lfMniyA+crQbvjgZjGFrjSFWS2/gUUvhp7KdnZJkaIlWR+hurmXqTD
mEA3AEjq2ATJHRBajti2nQUM3z4VY1x2e261wHff4NUijJ6KMeFWUNv+oED5mg06E0j3z0QCEK16
mNZAnSXi770tSsFUmdOdWfpgDw/59y1/X4xrVf/H9PVgGzUFSJWw6cTUgg9mb8I/DIsuJP9D2hSx
9yd18ZA267KfJXVr4TErV4MJbalDqNsSxoqkCW5ciE1ddx8etCS9ri7vIDTbqF8fdRm7QPH2n+Pa
sdfM2VfxhwknOQ7SMRIAmqsIK6N7f7o0ovzdQqMVA1j5CUDtEKQASCV9sC48Hkcslt+wUXcQXe7F
vUr3YBQUPlOsuWhTMw0PF7C+xDhCIZoGQAkvAzZ98ifGlyRom0PKxedh+AMFYvhzurKPTmGynOkX
NPyAArq9jolMCQ9Ng9JBQax4KMPh0nreHGKqB/tTHocrfEOJokaHVS6B6jSIuzyJD7Wc2OAITrd4
oMipZhSukIDo8FGdgHEsNydhyr5yHZWF0JyRJFHNaC7DSqGqDEkyRjN9KH9qyBUpuEz6ku/gQbjg
J+UfuLnSzbXYF/+0LUFw4SHHpwKC9Ft2I39ihNLXq9duynEXCMQePtkQLSegg0E8QBteSsu3DjnE
xF9sEEeeXPp2sG4NH9Ky0mEI3DvRzlNBLX6UTj3K+DYcVsF+wjHyPblt/JBtJIeRn7l1XDY8Oawu
ngYiNoZ3tGxNMyBNjKzqHrBoooYzObvAARLUNzC7Mzg848juezSanxHCOFbfhuX2UsC7xTLWcPsS
9sCI9vdTMWg3f9ryBtzS6Ar1jToyJ+OEud1TYaGP9qxNX5JY0nEjeL+xiHWR07N8lervSXC7K5Hd
b6CoQXb2/hcu480XcF56uejIWqv+seZS9qUJAsuuYF6yHqTCSh2NCKa+AnWWCfBye3vN0dkb/Z80
hOyr9G9TZLTpQ0ygObmjAbui9KBwSIPUIA7H45saLVIzr0h8LDeBy4ZYC+euOok6zuI8AuysWQJ8
3L7uOT6DKU3joYXzj7ysuLOvkNAe0B6Z4gG0h6GiCNGRZaAqndw3XcSAvTj3+de03nbTuvp+q34v
qsmcvPGM2wqUmA/49WX2lmBYbeJoQqd2tsdZXagyBhqmmaKJ+zF1JF3R46rma2OUXzpk8AoZjJnn
+L2Pk589fhsUtJokWH1F/SQWF16mItl4et4cVbs+g/lDVx+4Jd0lzpFqbo10M0wS34O5GMuloCAA
cK9nq4tKzLiFQoA23dsN0jE/ffs3e85+r2MNMNt5D6grIAOMHk+RdS0K0cM7zKX1vlpOgGg9Qhbz
yCFBpw2ytTxqGvG39y4nJX+uOaX+k0b/s78gRXtRd5qfKNFUjuUiGKD+X5usQp0NCMiuqBuhIlYy
nrX8gdjPOeh2ZVJCg/d+xH6t+vnmYDcGVIZJMo5f+GQxuYTiAIOpPwwt+CAT79NMhQdWn3rWZaeL
a53oxPQ7YQClpRAHz/rYBy4OwOqDbg/AqJKk7xLR8f5I/jXKLMeMhmi1yT5JmN3/m57MmqeNporl
B+c19PbQqmY1pVqCxjS58mlXFA8U8JI9j834QeWS0Cg8lkwEUETV1MXRXTz5XphmHwPa3TJV7Bru
bybN6aBp+HVJxzaMifJpEBh9d0SMTNWQsRaRrh2lulMjTgrP7PksY1I8c6lEJl5Z8F6M8pVB0SgH
qFEyocmvCsF39+L/0nZGh1O22nNNi8KfGiKGAN8EMqCz7e9F6JzvG9ffnYBLR3oOFKryOTQUMxAo
YvbtKU1pihOpNn4P+Mv8HA9CkZleYOU0lwwAIzt5kYhoWqAUA85Bjah1mGYLVOy/yWkpqZwjhFGG
3KvtR0iGBGAKlDj5XQ09sUHxLPWFh5I/XLp+BnuMVs/Ujthh5hhAzXPp2cKMDFq7TfGwxtVJbAt6
GnogyvCk27YP7mcsFEmXd2UmaigT8bnrm4aXyLaQl7efU+eqUA5YPFQZE+uTrd42VKfOufpzZcLb
ykArX793yeeA0d74AoihJXsFUwy8kMnEXysiAKWcKXFaORsMU1ANKphZUMZntM+P+vUlWwLkX1+V
3zsYZ/6ncifMy0fy4e6DaAgzddfytA3HdOouHflYBxWrXwBI5peYQKF3cw4K1WiBEWVw9lTOWd7C
ENaPNSBpjn6d++91qbPg/ahPaSyfXc+jSIE/aSjqO9gwlo0XfcrSLs7U8F9h7Y9uvaTFkxF0mE/7
iIxHEgZaIT2tEnQwx/7bA0nhie/35Rrkb41AZq693IvpQ3gfERiKgaQhso8JTuWMyJV1dGsTxd8K
qSHN/afLasKFQ5si4hj5Rf8YPrKYQvR1aCsC7X3OJEdZGOGqFZheHM4RufH72lHNmq2rfJxMjLGQ
h4sp377XXr7Ogw0q1T+6xv65AUbmhAtv+P5Nm52XXCBC24XA9hD/LBiwwWVb0sWEu6WOXdU9i/Eg
tv0b2tuEOhVo46Q0iEdkEJ2YLgOGlsvxnib1f9ldN4cybq72+0ZhmKGP/cbRFP+LA4sFkqlFFGTt
HqBcvvY+IJt/Siv6a8rDtijqa1ziJOkOmdrQSWtYcrUUu+X7NRO5LeDAyz+JUlGdwJWbSNMvfHCl
jZ2mUVYYg1Cm4/Yo6t/dYAwW91/LMlnMHjfVEsa1wMUItZ6gJRZBqbc7Q4VoFhzyAyP9q+d6vbGH
rgaEoOehmC1RfJdkFkl6OK7Gp+xRM9onMv9Tn+G70e8FOmVyAzekzpEMSk+I7UyqrnExMZtM1cRK
LgSNj+RVKbMlMfLfVTku5eb0sVkBbqVxFNo9TnWkR45J9wMhleD/rlrOi2HsGuzXpAgim1UqKtRD
8mJOO6OxT6AY3piTgfr/9tHpqOr7CK+I8TZeIA6sS2VzUhKUIhtEspbKL0SAEUTNak5C9t4mzbGz
RDbblsfDsbMcCMZ3XvPykpQX30ASObS19Bz/VZVY0/diLLcIqXQNin1NBPlnlRA0r5LLuq6VdgzI
6MV+qScANX/RVz3rT8U5sK3LV8Qk18dhtCfWMJdVrNVh2GHhF69447Zy4+f1dK5XMcPs6FTGbfEl
JFwhoQmAY194bHT0mkUOYn+RJcSrWA2tXg3PRrct65UsI/4Usv4G1ZEa4uFlXKlQI9sHgxGY666o
36rfoASj4WWZE4oUAwSff2XwZPpKmUS1qTcDYozqHEqXRrd6jon3bUiOZj45KYx2jKeGkpE/p8GM
CIGx58qo/PFRE0p6HVCkEviGct6RiSmSQEYIwGcchru0UwkjZK2+xY+rERN8/xDsLtpZM3SqpsuC
JxSyHmug58BFA0Kh8wF062dPPjaZDP3fmMvH2b//jVuYozIbYFJGEN8tq8vulcfdYIYPYddx1KVE
cBv53fv5IhdsG6rGxipgrfXFB4ru1r6dBOI6CjT1rk2mhXXjYMulEiS5jtDUZHT6Sto7IKAe8MBm
cBu+pahK4/65Qe4jSWgAvi40bdVFMpbSkkQ0VUr70a6tlDEWo7lB/V32L6KvgNmfoWtj17ktw/37
BX893NeZzcpFFq1Gg7BwhF3g3BnTWJj/UISCZ+JUyvDoevTkV5Edruo6qaqcbN8md/QNDvjTEkr1
gdDeYK1pbmFtnBO00BY02/BEEjGvNkP5m3XH7qt95KieQcMUiT51FcNE0s4kSXyien9Qt4kwwDg4
7HqmuviUDEDl872ieVTuntLXJ3wSxRtjeRxJOwEJJnHTtAxFif3mv3Ry2iOTUP+f3CfIkH5FukO1
OWNoI9Yc0n4wAZdMFTtXcEtEL7pqInV53Bx+9l8+vftK1bNm2YWVB61R68LAalfdeSfTBp1Yy3mB
FVT/dklk5Uq58BvFVizuVS/c/45uI4U3V+ufE/yMSVOb4mZ9Ndi+ylFW/n2zvfLOKqNoKCcifgD0
nvQGxjU6pAQ/hkQrX1jqq1UQBPeyevFWrNhEJZy4OqEYFNxe7iZFn530j3/+TfAvzK8n1cjfao0g
/4tvz2I7kdfmNBtlfWc/vhg5i5bMVthkw2+YaIGI61u89s+4WR/9j7Rewbrrg2AjMQnhTXh4p+gS
1CyllnLGJcbFPxziXqz2UxbII1fZCe3IlGIg994n0Lt5mmgi9VgQ9m4n2SbDuwlMookxHifX8jdW
iVR0sLn8d9tYWy+Ae5Es2HPA1TtzbzznyaSiLGU4mwJXx2T/9twHmGA8QPnS4m+N0VZODFaRoHIQ
sfpcEMT/FkBtodJ+befNU1Za+ZFf+syXBwpgbz3tx8v/tJ9nmBYeNpj+m80OZZybZxjYnPNQ95j+
4gOc3ZW2FZ0K2vreb0fCrUhP/6pzoPPrIlTXg8srkXr5N+nEFbuxhodG7yZvJFU9SXxIjIdPeT+j
LHx9BPZzdIdsaE1zYFrhFxzsPKxo/uS08TGK9zp+0n3gg6Z8JG9sggnH0Vorevku0aUNFZlGpMI+
FoUDdD3RFMmy+BWtCKACmPu0aExsGff2Z8NurDWYQnyVeeKdENs4064MQayGCtwXrxdV1r1uVs3H
pBUoVxV1bFNI9unbEDiwSITSEgmnf4CkxeEWEZseNucjdSeBY9DUBZwR/ezhwvqacNJlTF5XVTxS
g2Z20MS66neeMN+VlElslX6stafDxD5DLvaiiciYFzK9Rr8jad4kPoa6NJRamYzgpUQvhCaNa+e6
zZJUqKeVYVa0YHYZjiKvBWevJwiwZgBI/ipg64X34eL/MB/rmrg4hGTiAy4OhidsTr5RI8v3bSXI
KFGwmwlqkGKJvh3qbAJiNkYwfkS/lcMoR3suwfAxEliEjIxHZG0WDae2Q3/5AJB49RBXJiBPye++
zWqjS8fAlXj/dd0JdxVWGsh/FFs0BMsVdP3tiC3roYdVhnZ+3MWsIPMHrkl4ww1X7ACtyFTneiMc
HXQpLNVQrHH5H1LKKIfWkh+kehKMxd6wmbURU/qt/khb8pn0NDTMkdst2HFz6xu1Kq21JVVBb4J/
wSsDnknje3q+/Ja1ZiFcXxMh0iQYWUAvmTBGlJZHKpVVnxLNPaAzRCFejPkbPJvumiN/OqgKtxWP
wnmYsJ1fWY8WnpkPPnqe7SalZYhKOkt3nG85IxjemT6KIzHaZGV9EtqoXQ6TARV4yKaovX3Csvvp
oCQlvR5WTYNq3Ivp8WVMxwC84bZrUZGZb6v4ORUiOxb9iyNAqK9wTOj4UvXrqA7RGDf3CkOlyIH+
22syYpn+BooLzhVdo4V9hSeBkN4SoT6N3+MOm7dM5Gazs1LzMzPh0kybVfkQi1RMMqMUAZD71VGZ
pOKAdc2kEk0jg0hS74Tgy3WUEWMMgZVDzCA7j8oZMHTdR7bioyx8ZxF+yAbjpEfvDwbhZlO2WmcB
klDJfhj8ZGX6lYx4hbNkfQyJthiO4UNYLtIA+pIaXEwpwlKPnmgSwvPnz7q+JmFv4eLxR842iCjj
183cxMvhLloF60KEHtLNYqVE8GSAJ6AQSsbQLdJN2bBF/OZvejDPleAnll6rXKazrdQHOcq5T9Oi
QchMl3qXMPBsjJPgT35PEc7ZCk3CS971yvyU7hRsvHENE/Ve87xLZwjQnXD8qUa7I1WKWTdvyFUp
VU4sXdDajxGfIFQmHd3VuGEsQAec25U7HzEDrZgC8Q/wX7scQKt+DS4I8T/9N5CKRi+yvX3AAhfT
GEb3zbMvHhZ88EseofNSvIF5AU3Kjnxf27g+Qqu6XgQbYysj6eZ3tuvMb1UZ8hqB9KFnQObj08Vs
k/isQOX/8xqRwB0fw62V00Jv42KiDbN3e0mTmXwbCdZR8xUmBJSdhtQq646xjgiEOENteY36YrYu
ScMFQ82C06+naVgzxpJhd1bmShbxrE0ldwVekTFFnpQoJ2mv2gtHurFmG0JOxs7OLbO1v4f2AP9e
IOXl/r4XonGY1wvDgiaYiHyTdZNwjUqPggsmb12Fkl4JyOkvRN/1Bjt9Y6pxotKu8zh0eu3xpycK
8fQoF2uKUdbJsvcgKKe5xh2VQx25KeO4jgxPeA2bcD/dRudaBGdlyUgIk5Gfo275Wglp46w8svUP
hX5MMUpDnlffjQpnsoM29y9Sk7ql1I6rtBxFeD9LJBF5PEdYQ7+2SzIRMBWO/PrngxdP03gGRzjp
GVaURl6/O6SAM7r+Pt8XfM6wjYFb0pWIlJlYT6uTqcVuwMmD8ueGI449J6CCkvHF24KiJCqiQIIv
g0lKu/H/KM4cU3s4yw+RmFMu6haa0HTxmq4u5kmjsgRXxTDz3LiJ7YRxXHBHEePM5oGloJCVb4nW
Nr9/Ameoou64RlVaVPwMMNXPUA8ON8Rbc2eLHZXQus6853Ca9yKZLOSe5bhUncRERb5gOVHFxwGT
Bmk5/Vb9TuzhwWymnKH+wIX5e4w8UXo7FRAXXrk8Y+bDOP6j7BS8AEYbCzt86iu9B6hCdLuMAXk9
VYTD5TxqGtyN4RJx7kBoSf3XdJVoKouD7EXPCsvO+4ZmTIislBRMjoNSyttHgA6cDnEzoX+u/soA
qpbfgfsLWNfAnE6k48CaC36HqFI90HQfclT3VoO0S5tXrbatNmZ235W5rfdwAmY/MM07R/gG5MwB
tBCCDi3MTvHOumhzllFbB3MyRZSn0O+mqAzWpKNYp3VKrqkMLkNi5+Xi+gBLi5x72iId0DMgMqFQ
v/k7Y/gCJ70F/Q1uvJa34d/8ozEdkWW9MVIqC6aMe4NA8jRwPBRH56q9p+TyfyVjlRIFHognu5bB
NerZRtgfxP0E5h/G+MSwEl2t0BWAX79oR7mJhZ+MmhpXkBHNyI/2k/8QxVyCw/oknUzPzQfEADvi
wvesM798+qGAvipKjIRb2WXy5MQqZ90OuBHAnkQVRdJ5Zd4PJIZSbwqhqUQQCscWFmRnj7vSiLPu
y77DyZP368ujMJylqKbw4rkFtvnHcxLTCOClj8fkapDj+fwGWC5x3PbadLzays89jVG/FV0/7G4H
PHFSO7Basfp/KsfeOwLmLXA3bWpERk9n8oFFZHB3wjwnopzyU5qRmUuqebu8MxSLKiIH3FLEu20k
aDz0KAqtic+MKnIMpsLG/of8UVd5C+ugrjzPaGyPxlBlZ4I3r/roMNaY0Uo846FvxAOHB+3SiufN
SFStXHxyNl2SC9eea8EmAJZ0/k5ZLz0CH8crDCQmfxIfIK0Tqkyu1Llrb811RXQxh3vbAZCvyZkn
tSH7gxfG6aHPZnC4PGVTOMo6Ts31pTn4Onvm2LLoRb1WRn2yPecGRD1aD5CZlHFyAVJEemb0RhL5
BOakxGCXk2Ci4da6i4e3LcpO+vETw/1R52g90M5YhCxLUdYVLga51EgdvxzumKUKjlUXB6CCnv1J
umMvssssXr6UTcLYkeXNhQ8PGXCvHQRADATYnb2YHxZk/+ilZo/StASOyGe+RQrKm3mECazgUqc8
Zs7WhbUsvcjitEw4VyNAKcxx+vtf0GqBSwfxKtJjhA/gmSrR83C8UoyMADSJamdoEr9o+SZGWVw9
bzQIu/crBV0XrWnLvoQlL7jF8bzLq+o6sEWSB6U/A8nyE8WiLBA7f7KJdz8h2CZj0wmUNsGulgEM
WbiB4B5NzDeVhENSDbqa66RL5rUQg720IhlZvFNmivX9j59RXNxuvVKWC9gDO1fFHwgwtPCFGM3F
NzROOYMD7b9XR5KA8K7GVnyzRqaO4Mfvr6laT+yaHcfrtqGc3nLGSSmOmjRD/FiCRV3JIxZRB7/r
vX/zHoJagycMctZDD7cpcN1lAGR+QucmK8RQASH+gr2Ny1/pNNsxkmE2lt+AXcW05ojzBS5S1SVQ
Ia/xAvQH/iultcDNVMVt+RUmt2FnsHISQd/cuSe/Hf1arVg3raPix145E0loccnNK0PszfE/kMhp
Umt3IdcJ6FVbZkMvVB+Re5uJT2AVWB9sdek4FwaBj4RPytRJQs+T3vUD5aiSsTwur3VqNI/OFe3J
8xAvv2P2Qhz5AF9s8NvIlL5mN2XOSjFR1Dd5X1aLEQdxdTlkO7AVZc9kh9k8ZlFWOMWg6QQxCD7r
Xz1Qo5anAIW0NrCbzNb2akQEjtptGQI+PD0DIfOcgEDqC2Wnj16OOMDz184OtNW3Xh2GEvjJnVXo
IjsQ2qEQwSfPDIe6UCMSQBnrBXkI5mFtrA19yk6TogUB9N0tOyBAaD79g+BhJ9X/nKGEFQlp4QBE
44DiGulH0KjTz0lvKaoofUywka1VVEi0zbQhtRFagamskhCyljakMKt6iMwiwYJmvFpieghcHRGZ
TH2QbXTaTPLW4eYcEJMY4m9L+bb2OIUVElEoQrperdKmTDWHeU3W1h96Jce5roO7U9KUs7VK0EZT
b78ZKC7xJIKlwFhMVuha7k4rJAO+6Z0GXRnmmesh16EufRAwmpZTTOks3Zjj8+KuKGrF9QRPkyO5
kEPsPJs/albT4dMu321UCtJn0jTv/2q/lVKHMT+dUJcXGoLqct8zpeGqRlLdq1VwQnz/SppCGpe6
TtbcQ5akfFiFGbEpPX66h4FdUw2YnFrNaZDxnDgcBXispBwrWwAd5ypFTgrgW7IHwrghXB0WxmMx
SZfwlfBWJWk3Aea8lFLlwMHBBAZhd8/V1uz49r3dZ9zpZqJ6I9vnnEzJ6Sd0u4BEcohkkp99yEJ0
uJUS8cC6h5NgYbC2QUxx7koPXf80KPz8pm0Hk36RQByBqqEBz2nK4wXfdXUMPEhkbk1xzDASxE9z
gamBf7pC2dBx6AtPw6Qsnxou3rSeORqEamjgP7Sa7iVVAfs1ykC5PFrQRashU9kBNW9nzGbVNsnN
dhnMbZiaoeMWEOPKkieexPJRWxlDz2zcyGmgIaNOqup/Z8WwBiqLu2e6QGv3cdWpXi+1m96R8AVa
HG/8+wu7vF98CDkmFM0Qemt5htJ/8H9JgxwjjIWgYVu/hhN9G10YS+bQfxxrDk0cKrRBVatPapZI
fp6B7Cp/wZ4CY2q97ek7k9z+xZYFYh78A51lKe1JooHC8VrNTkLrNS3syPGwesa1ZQku2gNCxlWB
eliP1BQVkAycxelklkU0RWeHQn2mlxCUa1HSdjksUdd1Am4Fz52Vz82v3XEJMAMCdirv9cBk18rx
8lRenEm5HQcMI+hqNxwdLHvNvmk0F8RDUWQBB2YQlC+bQsKMKB//tqELEJIqI03x3g/vlVPg34Xk
+f+/zh4f1qQzaVjWY/feD5Ht2nYPuVIAplfsB6sni5RVOR5KOGEIhRParkCnll5LD2NvvrYzAXuY
oCNWr6su1BWiIY9rI3DfYkb18tus9Cz+W/u/u4qDdhqZHXSUkz8EZF/q91TbDBw/FinJOLpnpmHB
x0167xz4XognowdGp+HUEI2lA2dGTXaGVOImShFik564wt/fY3cGDfxrAgOvyU1MSFnjzg4i3K3P
eCyUyIfLVNqX9boO/82Xbh4jFLzfOq9uTKzkO0k2WqAUVdRISZEjwUJEY2ucfyvShr9+flBhybk+
6MsZZ6fP+ghq7GGm80P7xRuOylvi0ZK0X+tXfc5M/PElZxJD1eyfLrIRHGwqMwE+njVNB0uvqby1
bXq0SgOpHW2D/cDujBh11y5XoPx1eqhQdQcmFHwKr69PtfrDFv5u4m2lMIcYpgd8xWfQepYhp/Pb
M5Uib2YZzCwa3l4uxrSSG6NtFPvAK6Vy4h36KJNlAywwIXm7Zwotms9ySuK6ntFwgn60MkLE/lDF
DiHs4yyvTzwylqIS85DJdcxpT2ijGbN2sp+ZKGQ6hWkTyKNS/34fxOrdwdMDPVYk94zza7SG3M+W
KZPp2RkKNAW4HYn9p6WAYGYJuzMjgQdvVPF6uRjKLZfDSAC1weJD80ZaSmfdJLUvcgZvJo5lzNfp
7F9mKD/GQsNjV75OWbdIpGE+yqYiWKjDwSpjHj/NvZnJkHA6/rYJ9IAGrEkjE8qPRw8R352JlGQP
mKNJFuiXs6g6zKOLPpcmQ0jHANAj5c5SMKCOHzq6MVxuOZIwtqwC22eXJm63Z38e6HwPtjCFbLG6
XwVfR2jd898qTmFx7j78hKL/DWmk7stbFt6D5pPTCm2vEh3YDLeSYwTcMTY5yfsdoRMNacB7U7kL
FBvC/8NwyO8voGDmncK93Quplyfg7bmsR67Lpwek+JHDunKI78HRkaOKbXdy8TKqS+HAh0skiVqi
BHbNojMI86fsEKZX2OxZHU9BNFFM4IC/6d7DhaXFc5oC9XDc9pGWV1IyHAORukL4bH/Zww0a4Rps
PKGFbIHGMiCHTsazmvB9GzdjHo1RThcqCXpYgwveZUANmic2zFcCel7MT7xa+QvL92BE+JgrWYv3
6P7EJO/ybV+SGgMheaN527VNRDiccFA+8HMhkz8lrvRigOcJyny0raTkFKnEMnGD/f+/0w/NgnRM
zbc6bDhHsib8oiHN/ZC+gtcqdCBecqW10dutmGw0wMh3iN/aDpgbcenzBdcu5gq2t5GVcbT9N+Km
pOeEOMNEj6cqGdvAII48RQqCJyT3bDIM2rOePqhi5t03aA7fBwX/MkQsqFKCtRoeKVQUaSW5ExeQ
AaHdvxnFv0CTyd+2BRwR0vhl9bbCu0P9424MlnC/GWUBAccNtlLiu63oT6v2QeWaUkNNWwDqwqCK
n8RYbMH+yRJNBtaGpy79VuXD9OjS/T4Be//0OibW7bn6HqafAvEcbfx2Zbx3s82fhUGgsh2onMj+
1DJ1UDrKOhBxuu0X74xHha9nAmP29et2LCyBytq9uorgf0nuhyBcdM4QE+tozYkNmMDQjrqY/CEG
Gck2iLlyO28e89ufE0zBxaz9AKyoSOBOpd9Fodjt0PlpjzeKSSOu7acGqJeNxc/JdCb1IrIwTuv2
UHPQqmuSr95cUTgT5r2wsVop/j/eBYRHXKrArKMM6KMjGGTJq4zwWEjuf5YDNtmd7HfGw9XJ9To4
WjVYy97khrYuzvswNH4+63kJto5SXFCWAs9fomvHrf27b6dsPKTLBaTKfYNPspKntsKho+UGS35M
nO3subTwxcoQ9iaXfMdMrGgyQ4Y/D3KgU9vqVK58Yl8wkap/xI+6t/kU9R1+7hojdhYIGx50Izia
Oeex9MNC4cqwphrILP27FZr+8WEKSR0nPIZDOB8VCLm/DeNTiailrfd0prqLZ5najX1sKQe8yT5O
AcfrkhmagaEbC38Lo5X7nca//7QVM9HSHUS0bCGQwG8CMN0aXxHr846brP4zIvBdLOaQwGBnV4aw
Nh2XVNfpntjOAmEv88H2l++li/NCudhumuG9kUVnMheyoCCmmlUA0Mu5DRfrv/2Rw6A7s7AxV+lr
6cnpygDVoU2aSaY4zzRMLcyfVdbdHv+/esULUg2CE95rtv3WAEYAmtpQouoGcrD1O/ndf7j2PLW8
zsZq0LuvbiYp4N6pZpZOri+h1z8z0FnTC+hbgCGEC+Gme+Ll2/B7LQmLU4oXE9zBlHDTx1Z/kBy5
uy9FGV4sUUnjFEdWdUkgk60xJqpyPdzQ78t8FkTGAtXrzKAHem8z1UVxRXR5/1137bVqVgC9lzal
YctKoFSnXMNkiW5MQREb+FWTvSCqKuoheasnukvTKl+OGk3VLeSHvSAjdA0s1caJAFWsBdXLFQ0g
rpF+4npDPP/tOAkCkV01lNbEoqi1eRQeK77nhXEA/yofOuGpKb0+P6cHOI+DpwlcWy/ImFtmqTRh
Iv1vAU9KMUOqdycEoaVtm8dTfzN2g6buGkOvXMo5NQIY2uclpGs8RbAC4Ft05+wT7LCoaA9v2zx2
X8/weXvledHnHHoSiu0g4z/0h/53qItmiodNpn0nrycjv/gimW758F1tok2pNHJhNQhtIB4uozWY
7kvR/n27u8xMk88YXUYb3Y1cQUQTITt6gqfyFRiT4ajJxv1dxGnZoPzcsr3pdWDHxmsBxYYmetGp
sS3yq5LAAmIYgizSMaMWgieLFkr73wpWUTMC2oj+tAIy86LwnXc0rfc/ERj35EE4suOphpiUUdzn
43dBa0W8kxwXdbMz5gveBgJmAl/j/Q8+CU2F0Iusx7xK1KyHX4cunY7+V4K2nvzqehKkYvZcAcoE
HDZZh0Lb6dsJIjccsJmgcmZcR3/oyZeewyNTAm9M0cCTnu7hPddmlZcT7nK3692lQSeKLm2sC9Td
CoDazGgUJqjmcqK9Sr15OxQzs2KAYvJ0X4B0RpfaSH5rwlHi5Hn0Ihivnixnp1TFuH/Fjtem1N3M
bp/kwifpKr5+n3fZTi+AH8YyUry/+IlvzNXiGv9NlwVD4L+pbKZRnxez7h+XhNi1ZyJaQLxu0zYH
iRg5J6zdBs+YdOMD24Rmvs8RVUSXcX1zNa+4saO2u5wJ5SaJayVo3Z2kLJXChOjPixrjIZ5DYjZG
ItwJ3Hn0pN13xq3xcBEoKJoHkzm0DpxJXj5BRLKLT4KW9hivThFAqQKyYtL1XZtc9VFJwtxyYjbT
2tDj1mK55rHTsQrQemh8oDvqBheIUZvc9zDWUnIuGiOHAOLtXnobOH71nvOW6RiSsBvVBDE16+9H
udhc9eIQ/2AGbNsLzfbzyFi5nFJF4IpdACF8ecbIOUG303fVFXNNp/vy5lhhktC+5ylYgBs3OxT2
fLTLi0Wc8vH6ndDnubFF8DZZW8CPmzZbH1fTRLQPCtnb9uNwPbc1JUUDRcMDnx2mZU7BhhNBbVtO
mWpDZqTSPDvNHQQTDnloM7pf2vhfIZ/Bq4tR1557InzR9GPmB4ODGshYdJap1KvoCXBXDlqtCUnh
BLCTXJY601zxtDEiGEph3jfc4cWuG50fq96UbggFYwsHAA2VifUFUbCepMVn4oImrE7U9+o1XNOl
AQemkA9q9pC0fuvDl4Tid3h7FORHvMumxNRXLNvCQ5KjATcC499XHFDKv5OPgxFt41IIFIyOuzNj
5mTEG0pAzLjrvt64/11Vf98ZYZXFK2xJuj9SXXTZW8vdf02SLtVY5besLiZAfmjvj5cmOD8BjUzZ
+6DU3pS3p0bfPC8lNOMJFkC+Pgs4C1usUjbsiNALCFgYUJhTDxvlM5MqeD5TVmZTMJmh3AJR0QXS
UtJSKzdG53I47XXPeMCSGv/82SkquF2mNr14cJhCx7rq3OYAm1WpssfuqQ+YT4RdxQPPNswS0pZE
07URvbdyJlJ5v3/FASK84BBT3Zfcac2FuQ1WuLBZeQZnlCIydk+WgAlJuuedXCuRxRWRDziBvVC/
lCjdZRfRlN8nVXKD79O2WHsF13iTyFAuuZr6bBBrpbratgUI0pT4MqWN4YFaWi627qSWU/mAAUNy
CnEWBqU0xKLPuWf3y8MB6TCiXJFMCKuYPFu+AZr3jfooCaoQX6UdrKc8SUBKadf+S2Vdi7k0+CDF
HG6lI1Sxb+/Ezx4Jk3ve3gGcTrPExhqhc8t+USxz+kobklMzWh2jrtY7cV+43rPiIHYAJ+JGyNvy
7uD6+kX0u5vpmFxELKzZZAwIZLIQPSiih6/a/G2Op2ZZ5SmTz6eR+vfhwzyUgjNbIcmxUaLaRq0b
ZLBP39KbDFJ/xGVJlkSxZI84z/5OoSqnd8MCkvjhwLRvvwENROBEIPScNAjwbWo9odT5PePq3qRB
BpogwzSRNVjX1tx57qgfcl+F4P7d0agkMhjGqJ3VZtAo8uAeTNwCuKq8IduIy6Uz5v7sn+kR5GS/
JNX7AFHFzY+upXoscydr1zJn9FiosJgwqvYgJ559Q6SvDZPEN+DuPpVooi6p5cUYJHA7Tj+0PRgR
KZrdiV6AJDcC9und6UkV9dM6eciOkJiCdKobF0WLnx8Q0raUGZjkvjzillklSrTxbp9ZbYiMeG17
XZHJuJtpb9VDKGkwqgBkUZCjCkyOt2leP3sY1JH8KwusM7QSUEmQafuLvXFcsM4YS8MTyW9jXGbG
ALIdM6yAzzIYS8UYCsKKdYeNZpkNcewFVR8/3qbwlVMtvH8FcNa/gKIJp+3D3A+3bBcVeeLJqMo3
V40w9C7LwX8qLdrbFz9Akn8PCMD0H5guYshB/JULyXUTjOujelU5ZOaOq0tNFxeFe4W6yYvz2GAI
SstuUvdYTUrpM26WyNJVchmWZAb9V3k1Fl3r4pjRtxWrbwcbh3feWEEO6Zfkjj8xwLTwTpiZgbD8
F8fLumfSaaNbNbV2fO9GQNOqstLCsGZafWojfIX66s1u58w4En2GlXbG2qzPe6RUqbgHkR0Lr2Ww
FOZDqf/Av2QgoFQPCdRDjd+2AL+/Fp13XqCAqxszzezKBN6BVM1NuamOKbB7uL21QBuLlo5SO2md
7Lwm7nFcXwFtatV12tX2hv2Gkp4lfIYHzurmVN5478GEChJL/8ubhHJuVox1XGvMf0KIYFj7Fxzd
XAGJc8rIoCiIfmythG2Zs4LFGUYl+DhPyrmeN4rgG1+mJQcEAV+/5KpdSnIfrjg70zP4cFY5Biiy
w4XAXeovjLB0VZ+YApIfVnWK+pR+jDWhB5AVxjHcW6NRwCUxYRKeOa2Az7vRPPAbZqgwZS7t/nYf
PWBSRcDc/X0H5VlVAHescKI2h7dcY566wlsL6Y80JtU4sSIF1IoQL4/BES/W5yOxaC4EGtGyIo0h
MrD3jfudQKYwQwwotsKYjMmqIEx64TeU3vZW+lE1zyL7A2HB53D9ILR868pAxPfUufp6iqvCKgas
2r+qSKFd1eXop10xAn/5Vm9y0MnxCObllBJKkoUAA0b7mvMXaLKd7P8F/IxD9l2Xj2aB8oiso/ha
qF7OK0QqpAoMzBOCk6hlgl2yoNq2arUXbEYQ9DdyA1v5QG8CFt/8CRJFQurGBWCrsjntdg4Ff7H9
OMTNybZXUHqoUWIPVUj+EYJ5InuYClEFWveFkXSW+iDhWdNxR/iAjyeifZCz+HynOasA4QTL12ns
ZUeR1/zJgO7ojvZFzudvvq1Qpz0G8EemQM0Fj1WMKWB2uWDETSFGKM7sRnOpyHlwGig4Nt6HZR0H
q/RoiThB+QmJvJbxiJpl2ENUTQqBCS5JCT/+npp05BdSBoF5MjPWQljWulyYM1UwGGJ6hPbbYRvq
FV1sG6GXK8kWiC1Ulku9UicrKBYzXgSYvBcQFgBM0reZrQPng7DfOYheZKlOqOTMVppyRkUVC8X+
wCNyLNNSTOl3rEnc+FNqA37Eyo5U4vc+K5ZoVXE8zL1yeHUIWfCqscN/QQu75RHKrLI/J155lLXj
JVyxSVhbWz+lKODwrLL2CsH9VqhQtIku7fLjSke/kszGJdyEryqYuuEcGZ+jmTgtTFFH/l3xl4Ba
EN+4Jjdtv2tgAX5nPxvTm7jgHy7PuSpPkdz2yBNDfla2wku2tzBo6ipCartaO6QR0tifU9Y+DLhf
o6zZSdGjPX5HECUM2gL7k3z3V0jOFZs++4FsRXtjyrf9lXFYumbWlf6ejBBut7sU8eC/IXcd0SWR
r270fM5cytffWdMbSf0660/q8a+inzduAyoFO7AKRsClyw9B7RQUZplZyrx/D6Hw4GE9kPmCAilK
t3du77lXYmnSw91PotQ9ehZYzKgBeo0/dTQ8bMezpFhT/CiXlxpS9mwCT/hAziAoljV6noPvEhDJ
7GDY8/lPZ0/nlVwJO1QDduK09XawAk4gXF/X+8keNH/zcMWfeHT//g+7S3SLC+urY4LzHswY7TMi
nvCv3tJddHCG7RPqP1xV7g4qQoZmijKR33SfXYkUnyaBws2zGzzBuxgHTUaACORqojbS3KatAJbW
70PbxxcmXGoI1PcWfDXd1udWJm0tjqTzcww983uaNtslNVbqOq4Tme6v9NoIqXDBv9BqXfM+bAdH
O+hXDBta158D8WTYfOTfP/w1Jlw98j5XzZXi+i5+mYckY1Exl6PBZLWDtctxcR+u0lu65OwQlFHs
lytVWO8keafduo7Hi2cWXJktFiv8Wlihg8D8lrUXhrGhQzpzl4fm5jhJen6rcZ2wK0CC8kCN4sB3
Riet+Pt3Te7FQbIgGaR1pGolojPjuzpEZeP9AvaHrraZYQ7LhEAwHtMhNKj4JfVyXkmkeJ3/clsQ
sMaEaOYIvfH/AzlfEDwJZNcWtrv6Pb56XxN5vqw213wnHPZhr9Ni1Um/08eCDo0JT7Afz2t73Mxv
ycVZMLHsg+dFVFa1RalawgC3naYkq1qBN9NHqIMS4E/cDyUTL+/4jsKm2vEapc1ykjUdBy8ClXSv
UdAyZK02hLXRdZ06ke9Pfj3XO5ZOzZ9YkExvj9kdOqIfrTO57lWuJpaBtKepnFTFQFK/PSvZ57pZ
TiOQwAVtpHcDKsnwdhglEN8h+7dOnqOf+3z0gZFcSQUBwL/nnv8EzeJoYz2NniIyol697D2SJ5po
O0IGuVc49uYv74wR05pfEthWAQjcVQ7n052N4NRWB8ZHgOMDY8DgJNlugSsg2WaIXHh1ouFG+3cs
ZcGhcKMjfj5kMjhTWQysbcZfCGmv1vZ0Yl0R8IOwlGPAjmHW2OkQQI6wmW8otFr/DORIkc75fiCK
xZsjhAls6b4bu3JmMsEfPjIwVM6hCALit2D/CPprCoi8jgGqyw/0PWlhQJmE1wCsepGllXgeWTin
0W34xSMsP8rUz5UYnPeqS2IAkrWYVM0WcfC+nUNrKy944PYDbdSrkdQ3aDepg/iPEZ5or0oSEy5D
Sol63668XBjU8g2O5uIMxEayTauDOrK6lbfQNNF9oH0t7xuIGYKlx7/mqXnE2tZnsW3nqQU9O/Aq
xfV2VdllfTceTEQnBEr20b24XBYDe7yeH/Y4y9CPjpeyW89s6WqV4kwfhkft3dbaLKfiqEb78KzQ
evYtCPAX7pE/iDRuAUknIoxxYkwUFHA3kWJqnehU8olzJXXXd+drCeVuNpKEBkMFabIR8DMHMb1Q
QyaGYxn00jSEi9cO68oWKGuezrLA0hRQsCrayVgJvgmcpFtlnVy17UF/vTrzZ8Vka/snovQ7HAys
HCv7L5QgGHR3nPOGelpNHFu+wRB3Ih3kmH+m07teL7UglZgZ3bl/ILkucbtzQTEg33nbui/aTbIw
OGXrqlqmkEbgx5Hb6502GteYWTmsYgIr5YH17MgNUngf3jb9TCLAFopyGUbxAaaa+HFHzPrTAMOF
3K416f4bC8irDziqzvlE0wL4wRLinD1HQacZd141kVE+MpLrhzvc01PbBnLrO8Bv2aIn7NV0q07O
wc+1KNmIV8YD1yN7l/w8eJho2Jw/PJrSng7S3s+miFZKBr2FiX0+uCPDYwrGoq+USvqJuzC3ANYn
SLlVO7/jceK7S7Aip36ZjPTNm0cwRi0/BJf7MOMlwgNYIbkJHaLViNosVS0A95vN5JN2+gxgta0E
Rtfusdep3vAg6fxTDtbiCLKEOBA0TC4578pDhqLCwRfjpa8qhcmWqNY0tHf5A42pDVn3tNBanWhM
ck+4eqTs4LVWgHFHVZKVGR2L8aufawcFv1KpNXvQeQIgGW3lsHx7vYv0+CBxQfdRC83NlessHNbM
xpeB5K84drmYSoBa5FnGoPuZyGpPxjKnvakghoLZsQS1eLVsi9fyy0+jCpFVU/jmdKVk8A1hOvUJ
FyqmQ5ERQ1ixztzMD8JV+SQe2tFCBaK3R4Ed75nBFDzqp6qdAPYsrlG7mTLMvdYH5NPWZrAkXiyv
a0f5bXPu29D8in4glsQ0/g1Kxsm9RHNhnFj1MMvGNfqCtDuggPSojYcLocml1O32lYeMgMCsjycJ
1IbccVSJIGBt9r/B2mJPqL79VLDfMHxLSD2FfLWe0E7/9ST8aQRRrcAAHQCHH+IcYulKjH0Mq3Id
72u8+E23JZYnvuTxHm5vQdclhfAvNteYVdyb3sIRc4ATNCGNz87ZuURJyd4GMgJXFMCracZcqw8O
vXSM7EE4z++C1LfP171J3y/45WYSnXffok+Jr6EAvCPEbDd80+L11cSmCncN7otfPUn3Rzz68e6I
IOBSeDvhMKvEFEDo+2gYJIBPJmm2oBGbl8s0JLvVUQGrjVh6mBsZ33hQiF21El9vfaVjjUZcVMfG
TB4FpdVjqu6n25Es1SjUfend+n/6hVrxihym+Vdvp3v6+zHIaIAc/k31R3v7TGV4AJfek2Wny+Nr
hQvXOn+SYy3FnVJo0e8+nxaE6VOomfnHGst4Z2LVcXzSQ9d3HX60KX6dcxFJ7lBTP72Xm6QIlquJ
hl4cRYMz6KJw5EYxgMUWpxdNR/rEXuV2DyHQYVdF0vihsXT0IMiGlq7ZRn1rC/NISlxz6sQBYa5f
CxBtE36a0+QsE5D65Gegq81cFsaOK6tbZLs2l7whND+pTWjbMhh/dPUNsBt0XmyIzbf8G/J7R8Ef
htTSu3q/Oz8sjbXKj/naeokiDWSsyE5JGhTdw+lS2/5ne1uSvUBnbHVlN4hk6yPJSXzk0eV7Au7f
N/JLNtna4v8W6+AlUvt/smTWyqInYi/wvgE9RJq+UB864mwS7RWX60nUvQ4VDUJUrWgRRWZ+9u0p
LBKzgKqwinRxgUjPr05gPNiVOCRqaYlDXVZMtQEIPw9Vspjv+GhWiCG9jEYx1TNE4Z5wY2AYDv8g
bHaBbt60fZyKIe58ZvEgyrNkrAkHtKbnyn9HLdX0CCvN9dZ+eNDzch9rRW6YCdYxi7aMvNJWk53Y
nWjJrBsiR9e5IIxouk6GxCo0jETftWXf465TmorCj+FIuguDYMaARTi3HKI9rvBwdLh6Q761Mm8y
RRykyZXa9L4FYzQ3Hs26HvOdnxUgb3g3fo5N1eyY5AGI5HSs4bjdfILWm1P5jJjUYF+F7rZP/qkK
rn4oqp9drlh0ATPLTNtA215lRTU4qkSqqU+uCYX2n1wLfW9pWwLYCUy7pJYLL00LKSvHU+AM22C3
9W+jr+irUwJm98yb6wDQ0d7NpOAhnCFzsdk3X9638uTj/+pwcnrqH91WGF+2oP7TvXKq/H8idDLF
9YamDzbF2HMFhPWT7Uqyxts2SXzGLcuhfu7h6khb3A9eS6GQTR08GAJ8x3lJbt8WakkImn9Rr3Mu
AVU4YeSW09UA9MxaG44bA5yBx38yNAT6D0MSc4Pu2QUFo1F++hhaxLgAHnKcZ6+h8ZSrjkEysHzU
L6zvUlGvNZ1h828NRt4uhVZuyXcyaswdqGpRpSUgqkhBZSBlnAVSuNa8TIMG1bhqndEG0VerDOfe
l5M/uUy84NbeKdJSK/IV6vYZkNGbMjj70pupRO2ukZdvbOyppzvRaV5IeWEckoCTUdEWVi+F5Dn7
9RI461UYYe8xZNx7Hwy/Y812X+baZO9aDo0WcGZT5ThI3yIf0YSSqrJaJVgmoHTLK/xI/nENHgA8
FTO8hQ+84z1IRlWkeexAWRg7ZQdr5ZOUGs3t+DMk4/MXQM1IrOPCRBp4k5ypr21IcoPQxbePdPvk
aM6FEkLHUgL6t13TrE/SYf7rb/wh7ORiJi8AofYu/B6S7rgvlNREiVYf1Wjl6vdH79aPEzeVAA8u
0EL2+lrTx216Jw1onytpRbWw1poDiH36so5gi0+qdx7y8Mc12Rbl/IZR5EpaBMBSm2ySmc9R34z0
jAnGa3pNds2fICdxWJ/5r7F5Ld8EMZjHKs91MIECzAoXusvt0/5l4QAsly2ru3XrNlgPKOb1703n
NMetKo/P5Zy8O1uEWwAahnjD2jfyLXnqyBOf6mYE2cf4+WUE0hDyE6ePbERezb/A+GXiEdLLiL74
mFK7uYR7Ktp6v60DhYaV9p8EIl6anDJXlPoQch9kYW8RGRgZeP/uPfYgI7D33fZ3ab6RQrt6nfRu
M8cN5+haj8VpKfS9LFeR0JUt6S6KqXigeiK7RwAcyj3EWUB/H7fHDaWYSUcc22pMuRDLYDRG2sx2
Wo1roPNjSKirXh4WJjCoACXCORYIlA1FKCWGJhl2iyFZSWMVHNryIJSlCZ7y8kJPK+eAw5XmLiz1
tE4XAFtMAlYJuXfQ6VGpba8iMX+2K+CGnH51YZNWVNifvIwhtd5L+1YRs1yKM8D/Y0gMtnCwB7lv
v33e8y0Chc05ppePGT6kFW7Za9ust4SyXpAZNRgazFh/FeXPyJSnrVag3j4EYBge1PSmroF2pxHc
VEHv5Hgrl28nSXWIF9oiZB0C81Esc64aAMepLgihnrNNtCFwr/t2/JekimUGylhb7933C46qVnl0
H9HCaTyc4rtx5qj+Uvuq1kvSRN+uReuLqvXbGWWhvhNY+D0clnr+FMXR13vTbk6d30IxP2OHJfwB
sRw2QMGHoqA26rdNJVOYGOAkcLv1Ln0B8l5JtqlQwL0OpTAD24oskznuKqqALPjnG+/Hfp/xg9BT
nEu4fhPm5qAxmDb1FuJriSdeyDLC7TpMFFx7AH4YO5ZETRPCaBbTR/J3Yo4C+6gjOk60HfxmWRq1
RyA7I2OkFHp/xaG/k3xllNo9d4+qCal+jaSD0Jui5yPYx2AEePC6bN8HxDhMVrqJU6uuy8NeTvmx
YpF/qsdieurxfAHYTTpekALFEDa9yOQjGKwlYui3OgtzHpezn8Xn/2WBChpBvrsgHHm+96QvK5N/
neOp3R6D+fia1e8sZSl5+MO5zrk4407NzF5s+pVwZdyRQ+/XNvbLVMkYH/Euo21gDiPC2OGMJXT4
LmwuC6iVBQlpmKsdHlq4J+8CI5iu6mJN93sGeJPdeGatZWJR3m11pvPMuUK+6x2NU2a2nyrXqGPM
Lc8TXzKe8NMgqxbjyJ5RGxrVNyjrzbBAo3WG3k6FBsa/IAr3SU8aMEVrGaKoNgdeSN7yxWmCzRdz
wz84sILacnelivEBb4zfRCLYwfrY9MeeAdvqjO+lCMDidkQeIcR6FVkkA1mHYM74VI9c+X0z1Wx5
LvxEghbOwlZWR/chy/TVbKVspLce+tGtgWzCK3Z92UZUdsjlIoi/5MLo7DX/gWFrZvVm25cMbSC1
BQrdB4+/ggfgnpRLodbg291FF2j+z4fG6ziTUBDRZZiAR33FEtB4ercyDaPtgR19grrRA6tGnJJA
Hbk5cMCAM4eBcV/3XA2M7zJd2dJY/qt5HfXSt0x59HH5NshnWSt81fYdAuwwtIs1ZYsVFFO3FdXV
I5AdYeaaaA2ib7MawS7WffgToSd+F+OT5xpVsB8trm4gYL61zPRO/BG+LerteshtA896WSiQNB9G
vSVVSxuaNK/kHWxJXArBu4ScI4S91wrHFW3aoSlT7K0OvC4+dwJ3eSdAnrp48lbwjEWpBSYzUhPP
3TFebTpj9QhYU4di+QEMHbJPj8rsL3c8Rywa66PMLoOz5NljQN6HqrIaWGXdBnEgEmwAlXhuHLVl
9YHBLMkYHlCxfno59uS59nSFTTZQXYNujZ4fmbPbnk4h2VjLfJXFu6Em8JmqV7wrsQXJmohsl6cN
YC3SfoJw6s/QYuFj/X82J2b88vPDglfBrsTcMRBTiGGRkAI81gBcB9DPiVEFC4N9/04X6wVYRCk/
jKZe3T4J4sN/rZb5DbS17tbHHrhdOnuru5PE4E9TZp4FN2zHkTSUYUiXMUnJKzV+zDHg6dStqp1x
+dFXAlsByP1pGU6o7ILRY3rYAD7R5749u1RkR65Horl/pmNBvGEksWeOTZiEU3oFlzXCHtSOvNeY
8n1Ti0LNRJFotlJuRH1nbqbd3UX1hbCuMn60gBy3nqSV5iDpiUw6Y5vffW1w71thX/mKbi7wa6st
dxIlIQRyiBZDHo1Igy+1qzDb2h6f6rBfTYziltuO+PRCTWPuMjOKBVLaqBuvFbiJzFGRbv58QUAJ
yMhmhSYSTLkuzc/AcqhEMVqmNJWm4zt3tGlBfV4N6Fonb2GmK6f8kLBVxE+o+C/SJBYdqqT+ANPk
SgodwVL35GKeJb1sQMH3ZIXRIWIdkxuBwsnZ0GwfRbIw6tBokaaeI8veP4m5WQZ2DCeFlWJyuaW4
mE0XvxodP/SoOoFFcc6ZNoaE6PHNXuBytp8dyfAbiCbEHzh7JLtGxn0/vRjV4kbsootSAcCINBhM
oD7kpW0UvFM0Q2qmZrTfx6Na5EQuMeHNh+V+mO13c0OLaHg+2DiLxKveKbLKPQpoXmeToeLRCPqr
Wjk5i8mlk4WirnoflVRDdsN+IEJDLwZ9JSFb7v+OmiHs+6HbFW4MsOebj09ckEAQ6GP3vJQMMMSv
7gL6auaKa2WN+akJVX26oM1mmVb0GoB3WeVfObF3+kBgnYI+ro0T9DnxMM3hvmruWy9Se5zKEaq4
ws3JIKqtWFBvekhkX5d7ukeoU8rsq8tJNt/0RaEyvlGUZ97oS7UvV7mavYfcA0tUIJjUlm5K/Oks
liFLKQdSrfpVDx2Dp6NlsozcLHeOOEzXFR1RwNFofxcsGx3Ui4HvyumfL9kXYI2Lj2IgZT6wBVE/
1K0AuYqX0euMxvqyy3GME1GkD8ntEg5wUaqPT+ZJRWneih8Wh4xOxc46tYS6CZupy+mW/nHWQo0S
P6iWePEBzqejHC043JV+JT024A6PFqey0F9NCBeFGyaR+cZQngIH8k7JR+0s1lguVKUt+1lqZo29
W8Me3y55GtQ5AtFrpB2xeHj9k09J/mlwqg7JXWILI0zQPzRV92ynAZP9y11H/h2dNHvKfO0NEbDC
kztH81XXA/DmGtAmSEQp/GQDO+zwruquGhYmTT+ipXxvX9vb0EPsRonh3D+SCMgwHoRtJ/AqRlZP
ysQLErXx5MvhtBg3M444aM7i3cIx/8oBJyuCy+NNuzsLeRPgYwcKwCuWmjNEa9J4V9cY/USZ1egs
nZMdcZDUqWqxKecVgwvpvi8EoysPctut/CFB1FEOzORSFEEVf35lom2mMHvHYSkU0w4sFTdAns4F
dsJBZ6qoledIo+hnRr6RSzdQc7dnnHlV10g+9IrL9IUdqLo/Qh4No1680xw28kE86Xwhq+ICMIES
xhne2IgQ9OCZ4+aaeIZQ3vobF3Dzb32HUO3Gp4wDuTEfWhMeQV0e1DonF8VzSAqcKgh5qSpHD7nq
RCfpaSnryywykagyMvqoCeW7lnSBEcFDe22TB7pq8F6fC2ssv3GRpSt/ork0drdBidh9177Twtt3
jac5/PJv093fMgnVIyn9NSesJm5L6SkV+DgcvuusNC13WMpnpOohpiA+FhjOgQ1qeVoxtW3jJNfz
00MNH9wAE5bDF+7+2tfy6e4nwronNndVNONnVKy8r5uEGiU1SoVvK1U9aG0TPNK7F2rb9OBLGYZ1
VcKHb144YkKDEd8DruEfAQkvqcJnr+Wn27fItMqkSccEa3Q/dCuJ+vyjxWuODGPUFBVVv0AD9dj5
PEtnQYq3L19AWOE8CkVamSWWIasiryl2OSN9bYcg49vjA1oUbN7s5TA/UQcHMlkIDLDNbxbXDbQL
AjRHsArWiFLguS9oXjY0E/Rt9HehGDIfa5aIT5SWvYivtosuQqnocLGJwCD3nyx3yDQDpgrapjbP
BCUyKXcg8DYJPB2B8TBENPCM4yNOgUJI4CEqTzc1DXo5n8nANS3FcXjA/H2sp+MGQokikrF6anzj
RKtjb1GnS+EbS98cD6fcRxux7nwlR0jbkQnzJ9AM48C7tdrHDf9atu0eJ+sYLKX2MumGBb8D5Nq5
06h/n846shtKtABeQmBfiFszU3bLfcW+ziTz4fBi2N8J8uaWEWtxs226r9denFd5Rjrk/pWH04hk
Qmo40jA1oDLJc6ffDOAkgn1xKrikSTxdUKtwXaEKuyDFFp7IwmgPERxw+46P+TLPDYRsYprQKMQy
AolLX7JL1Lvt9QGTaTMKgMWpEs3EqATBOR87m7vvemHq4uXF8KNK4FUmGxkNfaE3Fo4TmnZ+Q4LL
nAXxFt81MQUXLCuB/CFe6fFASU63LIe7Hd+5lD8pB+WUYkyMZF4O0aXcTWyiWsTe04UQS6XwSCDf
OSrzmWmhotbOrFEIWifpG0LBMpP6pd6xPda9FgZKgFDFurhN/BVsAdW4zHPl0JIqZwfwsbQHnAHu
OWe+sIig9sadfTRt054non1HhjAx8s66gCF+bbmMG/Uw61oXGOm/abrKYgrR2XZJ+SQlJL7Xb88j
DDrGca5E5bSMFm/emCBaW9i27xHGUNYyhfhPcrC2PE/oWmZpajwuvxKan++vfee2OIoMafSuy6dk
Oe4VVnlxMTzOAgEGjqqBJwH4Oy5glO5lTpyBIlGQdpcKnECILTH23G0CFfH59Jc7IdRFAz7honpY
uDIvITz+koW+W/vmOfdiHD1Zk2hK3QFcooOENGPK06OveIrz5h/kD4GzjeVPec6HZ9/YE9tGsWOT
VJBJkAboZptW4i6YyFeaFUL3CIT7+j25ZYop4lV/NnwyulPx9REEfbeT8/DhWRdltJ1xcKqWYvB8
/Lg7yc+Pe0gB4BiosVTJvrmnDJvZ8obHXIp4IpUuzULIOoiV0oRIyASAgLDzLmrbuM7qifpLrb3o
uo2JNeeK4hOaHA7aCrkMM0LoflJ0wDLslEqr06i0zQlPCnCdxckV+rkv4Xr0/MJF76I8SMyN0g5k
e+vukUdlK93ULwsw2+oGdFpqZKkjASSEBGIV+kK01/D0Ki9YN0QHvg8XnLRBFrm2xx3FH0oJFs37
qAWhdGbkttIx5TzQqD/D8IZQgMj0hDvpPZi39RBnYBBBoCvDKqktADgBqkVGKsYKBkhuol/UJpgm
1yZaRngA15zbYiKUjXncwZhOb+7VBGsGjnVtPOQ9rQpq0btlM0ykqQ+4kiOdQ/bTn6H5G7eMfdl/
zarix4pc9cOgAEjgKY2Km22ZCWvRMNM33amoY6vztpUXumSNChiOt+2+pFeJeM0h88sqqjlPP6dQ
AwVX1OMIWuPHUs6yaKK+JF0i/+oks4/baHHWwpgb4YlMx/QYuGNtuBOICH/JxCtyls6BqqrBQFLL
fyeSESIB3MvHPlnCc5rQe3F8O19VkJMNjkNrEFb7lirUS+LVTF0Abk5wL3BnRP1FRWoc5T2/Ulv2
sLHecEOnRmWBYTT4ySKOXyM5vJkVSGMKklgzhhmdKayQfWGk7wuBmxXfUvFRE8cOYMs9jOFl+G9D
y5Dk/Cm7bdQzcwhz2VtWOitngsNTqF4GGzBN8qgBrn17aNB5WOyBGkZ//a2Re35sIGb/iboCuox5
XnmU78UoOgcOmiaEdWSAJOTNZLY5lRa1ezEtcYUQIn4X5PuAKbvVJwT5CUeilEpAKK54hstAhkfK
USyHItnKxbeggqPsTShUHDUSi+X6bfb879lwm0r+fdbKwZb8BAh1bXLPrkhw7c8WnoHpI2pSd6DS
5HQiwUohHRBP4g0+ntmO6Qy3kca9eMAF4q5T8eSntY4+jp94LI89ocoKcMCicN7S8v+7fQNpcJG3
5vS9AldFG3dY05RlMpaE1Go+kuqGx414Vwl0G1yg4p601MtD2rBebmKA8v/nk1bCBC9kSeaRcpR3
ZKfUG08ab4om4cTB+bkSl09/s2zKzMvaSMok+W5bbK3lNo9Gkf6ctsDHY+0EByOEYMZKOc1iv90Y
EAB5WoNIpgAFzAtk8zEYtdp/DBzojyZ8oNeVqTtlH8i8Avye17DiX5tBuSLBCE3IV7tReLBFpAVy
cvxE4CXuG7G1j2xaGKGrmeh3Hd9bnV6skknNudpH2/lvqCAt3SqROHfmU9sF7SlBMp0U3l8drdGF
Xddx/MgUEtjY59dvDdFtGBR7MeqwVyftZWC54HJuj28+xR9gZjAgUgM5v0dMP43zr72NFQ6w6u9e
DbiwqFYLIjyWy8JzyHpJuTEYXo55tHb5VZPXCg2rcRckkpaoxSMBcI4P5jKCwld59GDGHCZ/G3BZ
DkdsqdD6O+cNs6s0nHg/43kLpxPsxJnfE5uWz0YjXiKzWLZZypr/JNR1WNVW7VftOPjOfq7PJLIK
ybX3F1x7m4rk+aka6Ug1q4obV1PoCO/17nCBporqyKMGM0pMjkduC+qmL+//uH8UO0Tjmw7N28F7
tFed8yAHOaYnMbVYUyhgPIj/VsQ7z46+/FivNbQQEFy3fo0vLaVm9sHoEt4ZWV8dvogmZWnHioUm
HPXSacp1jIB6v/l1NBQLwwVoXX45hk+LZUEg8kx9MQ/w/ujYGjGPWH+X6VFhXolbuVehyBFQdGF9
Eh7BfrdDknD6AIvu1CQu72tjCkZrwRD+Qjd2yGXV8yg2jS2rxU9d+lg2dBZOA1fhEZnZ45x/00bl
H/PxPYr2vcpRHBek9x5EPQAlAwvM0EdWQo43fT9imqkW/gvkeAzoUwi0d5f+lYMLzofjsb+7y9mX
6hzZ22TfSeteaimd/RWlZDZw0G2IJvOqQEYxDp0jWRMb8xQHyl54T2+W71AU3xOFFjTYQ9rQw1CI
d+UZUjSHU6G2dW1a0JKy8ZhJ9H7AE6/cr3M5ELiZr+VVR5OSklj1QlgtXfQl+BY2k/tavz7DABG8
e2Xk9fOnjMP1GCmPEyJYrdOJZHfkIOSndxwRZvATevzn5y15OGxjSWjkFVwnvpSHn7toQBPHImX2
+/2ftlcIIbDM9HsAFgu+KkS94qsxJU9lUdN5BeFuHOST2KomqI+0ztTa8EleBTiDPoHCCOmNJ/kF
fRMyof+vdiZdyDiAMzUL4QdrsWl+MyRnCUS5+VE/KT6vPFzr338GhHiSye2HyY7NsLf5APGRUWyd
e03l5VGKVqUeQgLo8yBJcdegxUuzkdNCO5ucpuwr5/l7w/Lp++bNKqNAD3yTzDYeuJrPrXaK8TeL
pYfyhYmbf059uHEYZsqe6S6arshRyVpA7R1Ej5BI2TEGSE073GrF3TnlRxZs/RlQimvjUWStRo/B
0YW7xOwfFo5EPs+aC5OoCJnf3E/2RpPE/GRwMxN2hCruASFNaTmBhGG7pGI6zT96ozCEU7t83tEb
vnhwV5yiv1GvJ0WKpBaT3pwm9pXchpwCiGRSa2zFDrV7/jEVaFkwHhgTslg4wHzuPzW2RBPkZvGQ
6FUgI4EX5jq6TUSFcV7e2jDPf+h82J5+th1bFMASF2Shh1hJZBWJSNKoUvhTlRn2JkuJokVQLzfZ
+n9hGIbxZNNWoDGWexj71IWIExpJ4pj5RYOISROQeh/tTPWLDds3Mmie08Qpy6zR/tTf5d4AGXb0
aJ+JNzIcrxfIKsGSeKQz9v3ZMj1/ssREszfqPPHQtjLjlBzUwWkr3rTGPZYLl95O9mYdoSnFHVb4
tajFSNSLax2+MYBuuVtTXFMTNgc6tRf9bTZq5jgvfDJFOE3ryUoBJXMVIezo0hcP9fTq+O8uhFtM
mfKUKa1CVmZZjXUGRQpkKO7Aw49WWUxCKSzGE5Ct7vKzTQplCxUZtsn8jFifZ1D/XMa+vlf/VC6M
3RQ1/KhbItDcHgMGkTalnKnwP2h7wk4WlLSxAbR14FU9gOq4v3aFO+44F/L3Wn6AB9i/6DjlzYzo
RX3J3HKso0u7zPlkgd07L5+q7A1b3NwqniwzZWtdI/QFl5ritP5qIllQFMPDs/T4DlqpXY3Ta4qn
PlwSTgqK6CTQopEQ8sctvyLL1Va6VNwkhy/5bQvC5KDTJY5M/NbMHuxrnBNCGbLwTQFbGueEC2Eb
ccXgjkl6SVpZRe70BAAiTqo0zL0ZZm5WxThEiG3hMVucWPoy8vKbm6eUBwQ+vaj02byqnwGnn9gI
w9UNAH8ijZvuLkKln0K3Wn9ThpOhZCF8272UHEgP6YZReEHtn5V6jMtNn+ii3ZnMuHm6tY3QZE2U
2/51grWmXAyp8gkCeAA/gcHTFNnXDOFgzTP3agjx1ASUfPmRCsVNHr54s4y5mVG5YwDeEXb6zgQM
Gcveiy2P77ooOuJ9z7F7CxWAxilTjqAof6wl9KIki/blem/9+/Md7uK852AI/uknt7FHfBs/6aUT
LrCMS+nRw39wgqz690BUzfOptlKFAva5rfRuy4jMidm6OrPXl+mX4lzDVFKoGQzWHHz9b48u5vf9
IvQKwRpIKYkbneVSN/7LGkL7X9y5Pb3UcK0nHmEGmm4kGgU9ocG5hESC03ca9FnUUDHOHNuo+pkT
n//24t/lWZCPKWMlDZ1KVf6SVBS3o/AhN19TAyHAut+Q5SYQydrK8K4P2o2BheBNAkX/DTpywFnZ
KoW3jrtA+G+79gqVv5ivGsl3e72n+FdOuanZQnqgVKZgcjOLSV8JhGJhGS4m4wdraAbUibYHsN5g
4zRUZ5v5V0POwdfncRrhXHmB5menSlLm9zoHl9xUi5HtkY4k2Wqq6fxJddNNiekiVpcQsTEnfI9x
Bu3YvjIIwgFNjmJObomvAwwIeVVKTB0MSwzlpXMuFkoogLlilhxmXeIgE99LGXdJ2JegbLgvuFRy
QChnVSS4HS+p+mIuiNt5hnUQVoRG6u0KW0WCSVMCL0AUzqj9GSjqNIhCs313VbQ+wE2Bpt2o8Bfd
972IxysI6tlMjW2bSHf48IZYB+/jGOyBL06drxtXCSL7iwxgoLbp7plNroz3jymz9ivr5n47R26T
PZNhm7dlDCNBZ+FrZzpAfdIYSE4xgJilHNWEf3YKLKG5YiGtIDDnBIoiiaRPNMuQL7JCsm+Ce5Go
nLZLE0H76dlsX6ZxY9Kb/gasqg5EP/EP658Ohid7hv7Plav/aOnKvGSvSfvO97jLS4/VLCKyolwn
Bd9+Ktd7NvUYzrO66ctsnS0BN5hR3RIViNhmQzzu6qEk5uSahZgnTAUWndZrnN677ARuVVWkgd75
2pMB/+Gs/NBnx0Q00dc6XlO5ZGxp5B+IlwWpIkKOYDrctnqdCP4G7OHPWfnLznVeCDjc+4+PGoAI
gNAdews11IS44T0OM26OWPnCdpzW++nhcsk1zwnSwJ/QhDtT7/O5rg7XYQcxLbkpEM67SJ+DW9qC
ABjQ0IPZlC+L3ZrP5HU+y5o3RiBG6eOuaZAnyx72ux3ugaNgDDOYjX56Umt/huY/cjbmqipjI9LN
xsNvZDII2mGSn7Y6tp5/Od3nRqnMa2igt+A4a/MMn95uz465Ze4Ilo5MF9RtMTdbolrGwBhTDtPG
9pKxO6wcDG5h/MhuXaEL2Ff588s+pQMR7ioDkMgC9zeueKY87djjP8T4QGtX7eZ+XTP0nBGxyvQL
ygNualFGHTbHuQRvW2feXsGPRJkbrk+LBPGghLF3aNxbT/LlniJEDi5INHbp7FdfxZ0uQSpr3Rb3
AK9Z/+QmxlPAydxMiZBndQDyXThou94aCYt6SuMoieCv1ibJ4dvIDrSlK5G1bVi+6r/P0XL2cDHS
eRhpfjwt+mTagRpF9oDdQK6gzz6QDuEkDOAAQslSJ4KFy02c9PUP518fWGx/tUQufUyat19+B0Wt
onvgjyk4YuuG5JKCsNSjKl1pYKOvD6zRsrNCXQKxoFDrXFK1u0FaLGutPT06nUqKHjF+uBShZCyC
LKutuC4JHOwOfA4QwHESZfAgzXPZjdzdD+bMt24/sUYIAIK7KlpTEU9aCAqbwf8w0CGzV+sRISTr
wzqGQkcRHR1S6mVo7J9A+z4GInghcApaaD331rIOkcuLrCIktufkiQBeS9McJL2MtibjYTyHoYyv
WntWzOMmmav+PDO+Qrd7MyniZMhhqRouuwwa7NdpGX36pCn5c9f07Cpobhf46b7FIHsxM/QllwQ8
oSd5ur4NBlWTeoLziV+xQPCvufLRl2YkJ7XpaXIt9QPlqKkFlgyy5CnqTIehcm83v+oNId8MGjvQ
m59RIo7hHq1vJpZn2DUbrcBn/VlgeceFDKzYH11I0rK5VQR9JMEV0AnvjYHvnsL6Ca0I5c/mdOyb
pwmre2+EeeIPIQ3HAoW0E6DAf8TUpwVmpBFS4BdvKmeIgq4FYURu+YbyAu2SIZynMbc/jVsHakI/
doEBfNT9ZyjbS1phr7Rf7WwxcWF2kNr6K3PwtbHjFSrQ24EhoXmLIoS1lADvwkY4hzQuyTAPjbEu
Gqc783+Aq/XqRBSdCQdI7Bj8HZd7PVJSb0gSoL2o2Pb86/UAKkWBofOhCGm3zPDJCGH42M1J6Reb
brtNIq+4dYcjsJULUU5QWJHhU3DvbLP0fCnldJg67iGeGASI0EpGDwBL5fFKvztXaVN476/KPwXd
L9g1of85sPYlme7npA+Jp6lssfOlUM+ISOrJVufgZ5ju/VhkFrgpK4Ir5PqKAGuE9FbEixAM5EmY
VhMp67UBsy+5aotMFRfVpfbc2wV93RYje0Fywhl7jwPPefKMk6mPfxw8XuUeyC+DpOTg/80U/0Tt
OQbAbUwJBESov33A0c/tFAMp1SL7ICoICnZmGzYzyDyLaDGo/YWAHu1WDGqQUJuOAehtyZFMIlMD
CVdqEdHRTb0kxLYfgwmPCUst8+gBNGwkJOCih8rKudSlfu4W/HppGGxNUeNEJYdDfWheSSkvQqkO
fYgoGlpLKGBOq9NRrzPK3PRruLPvF9x2h0diYLXMVwfwbPITZHsaLY1zhHAY+QcULRlMJtjyRsQs
7pg81kzHMUeIOHFtml9nNTDNLNDagBBlTS3nUzsk3LZ22OIBhRgjNGq58SR0RsXe/QYlWXhfRHnM
SKO3+XPucqIVhtGmkn3ca+RH8okllyfGJKpn2XDlS0nrMYMxrSZcm8h5SG444K824TDdOYH/8v0o
e4+D3m/2DY2BOfuTSGGF4K9wpvPhy2KCryeGJeMuG6UI5MC8t2AJILopads9C6KqQv5wWlbAHRZO
3SPO1WwcAsIHoSSGTbtSQVZ5NYcMT3zsTlJ3KB866zgrs+V0fP5x36Kl4Rzat9DE3LA0Z1ZXsG3W
4oTRAnbAgKRJIxWW5nlWLFKonsxQBEM1J+CrhXsw4/wQ82Mcw5PGc1sS+mXtRq4G6/6sr4w4peZl
SPL2HJPb8+B5jrmfN8WbrJ5klBuKiMMrEVNJ7HrkB0LU4u9hJFDUkxQdHqwr5KzGXKrU4F6m32lw
Fsx4icy5B/GuMEqDHhwkP0jWDOMtifoL0Ox/D9RjOM+YHeG/nTvgSTeIorGmro2TEDsViV5Hx+8C
SksgYOIUNXzQ7ZzxUi0xt5or1mSM0Eo4XjnfoA5cm+Kn1B/zcQseycBY7tB+cj9VMB8buaZ4Q8E9
zs68+q3mIMen7wdXbKM3UuLQwp2pm5wukHNPQgI5JEK+3wau9SH+TerTgLaqHA99LcEmN3xil43L
btCsobNiyrOdZgrqmtCAbpzl6bRQOPrX2uEr4RwyisoXPNfs+GdkenbRICn2QC77nHfsCA6L0XVE
QDDam0Wn8JXcsUkGCNvKokniBFXarpTWzHeBKohdzxVvDiQWDB71jgvtkOE8BNBq98uDUmpuegpb
6zf8lNKKK1RNGAGdHmI99no+pb6gE3KPCnfuh7Pu/qyctniS66+4myR31zEElieuFLveivLVnim9
0djbjGdLhedu53FbPLT/HjMZNCqYdQHJWb7bVw/Cb+vNw1atYZP4Y8OAj2DTo5GluG+0kpNjViht
TqNkfL2tdb7qHfIesZMlbycPZXM3kh9HM6p8P8UfbKhwcjHnhJ+6x6x57QPP1a5VqQEAj+EwaUCw
trufbz3QFuexTNCUS2Y0fOjbdD4/57RaSNhwXQk59IlEKD+1yilfxClYqpL27tRmM0XcwWQxtbnN
mbsMqGZUagf5GTYegulmcLjD3QNa04dwhirdF9vPtcUdLR1UNR6i9oSlvLUeb9yQyrQ+8ovIRf/w
jNsALzHEF8ZmxrBK2C8KFxXOwHS36VXMAS38u722XNila0pPU1D7XypkPiAmtSLJFyyebnPr9Lw7
yFm+nVO88ITUdTSNAFu9eXHquBmnWLzzswoYH8JUm/ruHl9dhYrnKDKTNvUu+/1NV4HRhLMnIr5m
+GwXecO7g+xuiPBOa70tj4JWMom6N48LejgS4OEUfS6UiJIOg0u9f74CjFgwFSIr2sO/5BBv5Nuc
n6SLym10kNIFbvtXWbOUkHlywlNMW+jqm6GOlmjLY3CtRjbMn3y8WtTO01nGcNyIVxL6HyWvyUnk
TiIsFsGrre51Z5Y+9bvpjUrbveCquj4bk3egL4GWcq7Ohf8gtAYxeSYt8Qm9sqgXbJbKg+VlsUxQ
Ham9p0cpoTFzTeXAh+9K9fa6Hnoc+52XYF6BhlUWoAbx0PH4I03+flBj6B/JoVXMtWYfCdY/u3PZ
B8s+vrnGfZ6A8PH7oDBIClswgI9DBzMJqKcGlzntuGPHO9xgVR+t+rdLqp+U9TDhfrzE8jtudgkg
0WVTlXVEzoNIHt4TB68gwmx5icYmH4mev8lM1Ni9tp5+/BD5m+iVBZOSvP/UKHa353cCTkl9CqUh
iuYFWMIb2InXoshte/qOHNrzbQvJgTMSCZuSk4n/tO3w94kVNIxUJHY1Uw7JNKMw0b3ICSJOGOBB
dDCM6VG4BEzVZuffYM7tewoE8L6bugVnpSYZXM3QoJDnNmZdJNdxVJdAuAhBlIHEt3b8CVTELUGS
QnFog5q3nonYKDTsbdAlCGZUoomhWiQ/OdiyczKBOcXCPVo+EIQYZNPBfYwGw1Jmo8vEcelabWbS
F50HF/GX3GXm7NWxYoP+8N+a9jCM+k/WJaK2JW96aYynalF3p8iDZbfCSP2OCpiHLrfZFH1A7tWr
hWQUqRUMY0g67b1TKqh/l+0o/5dTIA+vjxaADPmL+yrML4DmkLg09FhaCE5ITqgHQJT2bFlfeQnl
F8w0PlG1dWy66DMeq1gCF9rU7rfyid6zWQqjwaXNwtTWD9jYUYll4JIhGUqCRtIZ4dD3ZoUg2Pf8
Z7l35+auvGmQsjmFx714dvfNNBNJaXgYaHOJEV1eJ7l1OEocqw+bE9yFci5jEfhflF+Z1BegXcFK
u5AoXjLXBFh6Wj7oLM7/YQzRIwP8BHk7exRkRXLpCKgLZOe+E/Rktm/D41vEujPltDhpy2UnPSSP
/j3wNP8mk7P3kYaOvFpJlnLmUY2W5cyzNlRYVVHQlEq9n7Po89wMYL/O4ms4rtjErXQ5qT6aIWBf
IAHGRev/W2j/eQ1ocCqxUimTSnpJH5bRQTaF7DYuYmftk8GWktOjBrZaHLmshvPC6X9JhGVyXvHI
EJFgzjDEHj6OgMEQWdO7SBZjc7AuljbdH9DBxSBE9/11+9Kyy/qWR1JJMywebw4K59/3QLiVXrVI
N7xlWNsDgADdvDWvJac18fdS5DDAeQmsXBcoUbpwWDmsJ59k1ZmzyUkui+QWRGrVV+X9+zX5WzrQ
C9Gri0fq7Ugpvpile0DrcvVVewwKzhRxtcit/y4HzEI7rJravVSrGGQGrqRQs8G6cGMkXJummw+1
XaUuf1KLnFkW+CvbkcpPuTh51m7PL4er+GmLzahMX6xIXvmA2whLuWzZTXYQr0G1MQSrHMHHfLgB
0nJn0q1UrXB3yWFyxHGO1winu1h5WF/mAbzrGdqvNzWFATsU8VHJoRovWzu7Ekb6JnBeivh2brdC
Qho0VLGVTauKEtPDGo6mrfE7WPunD9y8LOawKXQ6CBzJyKxMXAd1W9/xp7deA3dgvNQAHr3zT7e4
/Owc9rIU/SSOZM78wxAWDPkX/2aase1ta1lgZgLGdYcCfuBoEW/I1EpJBUMyErc+sPIAxnXcgCHP
JBPm8T9FE9Q+MhdNnA6QLnmVEG8nRLQQekp99NTEPpQ8l7zgyF+CKdDvyUTDmVgltzSFl91gotY7
Ol/NlO0hoxa5O4u0YsnOnBJ8+Xwvzs+E7b3FUP+sJPmeWIe1AliFi3uVMQjT9yY36ssHAi4sXZQo
mre/sgFh+0yNVOfOz/+UHOHp5sJZVsiM7Se8g+THeDM/8uThxUH54UbOYpvn88ASfLJke3wxC02m
97gKqWss2mGLpFZWwt9RNoKi6RQnQH+blOUJS7ZXrvqT6tMZBfMpMYDz05Vpyh8LZ0X/7PSlRD/U
//xZomeyqeZ/KqGA7aCuLdMCUIXwl/DP7LCsb+TkLauMmXmgkXvyn15IsEo2ZRdgUZsgM+2z9EKQ
k/49ABRcWeXaC355Eb0q80Reh23WHWmpzOmiGMd8KYFpYVPRhILHNgwbIHgPFBhuzWw7uP8G+lje
LZgf5DXL+uja6I+CQA4rxamFLC4FhHvYAnKUmlStESKaMnOTiCELn84SF4pvMnqL7oLzMU9H08YM
9b842c7kqtytMQTRvh9Pu7iwLrUtjFzY/vMcc/VNlgLEDXqLJRblYu7tvONzhgSdoWJbjOH8uUvG
mD48dnLQ1w2eXJj+1FnO7H/EyiHz998U9yUd7EdKPXULq9ZtF0fjupM1u40lI4k6ji6K+p/ZGXRf
Wiz7KNKuMmo2QxmRsLphyFx33tymXuEzOrSkuJA19mORou2vJmLAk8OxWZMMfBAuM5VQN90heTFY
KST93CkVh82jYmxQaqL14KC31bkRpAjws1kRTRqjRt6LXHeGjuoNdd3fYTaQSf/UlAbfvZ9+LM8W
6bgAYBoP9EiH+kDtea6z7GzIsez9gHFs+/DOpyNmhKTxvvUSRU9C4DHER+xXrS4Eb4e1LYGnxvtp
OqdNWdGFKMqgfWuMXK9WyqKpF+OjQUc8jB2Qae8nK+TbZ3TqPyPi8eCajB2a9VGGD57j8Ufo2IkB
bO+emHki2JwBrNFddZwxWBI6GyglFy3Ypn1ufaCUkNLhsOgCJTfu26KzOWXFg47MnRchQWSv6+UW
Cn6EFJ2DgPuM+6Va9HMzVlhZtfXUF7V9RbsikcArIf6vzphAMdWwdWJY29dWCnWdnqar9sbApZwB
yemYlxklKso8I+ijreTqXiEKASgjBm811w1pODfIrHWg9G7g8PA2C+j9X5PInSnvWDnOz+Nst0RN
/SWUxLRIgH7EXWUOvPaY/cwhX/CbZMBn1aGbyO8pzhBZT/2P7MixnJ/yEhQB7ehE1vx2BXx9EiZd
yvfSGVyDteTTPxUgAj8eMto9uvQUmfJQF8Tfu9kG2u+EajW0LUPoBJPW1jatwErU0lNr7aQV5wsY
j8P8D8ZGH6hH+J4FQherzt3g6voK0FPzrleKykc+DqnvZ5J7LtUlcuyV0j819tReYOw4uK4JYopG
/ZxHyTCYxidpZqwmHCzU4T+u7tgrOwMDOba22RxLbvMU0PNZ43blLxAlSAVp6/jQxxEKI2Zf2bzc
J2rVaDnNZNgNNwUasICpPk/eJh2M2ieOqOa0PbHj/cTweeFX1DrQYxaIEv3rft06UuO25yqIFl++
lmzbUD+IQYe51xbWKuyUrXyQtZvPvo+iW1ZbQ6ZwooIbz97THKf63bgUKl1ZJ3FRyXZ6fQ/NXFrU
zhsbtnrRe2sefqUPIZmuH6tYupZwaIf8yZ7SkhlQkCq31Lsa5R0Ta/A5TM34AMl57JlpHHp3Nykg
pvovgt76jPBqFbNjFo0Gi3TXC77Qcfw7xsKCj2VJBRmKg7vYSZ9uclWBdNIb2HLBykiItMh0OTUm
1HdGeyvp/j70BF7TBq3Hy8ytwzkhvYq3Jq4ZTBl5AmFgjh6vSdK3letlbP05OKeZvD79Kgr2AgHQ
URns9TRFwUztPVPIWWxd9k55bGfK/RWHMi17idU+FhJjnC586OpBZrP/MlZho0F53CkoCjDDIs5B
j/zdiYZE6W+h8e8fyMoy54KaFt0xYxkomBUKoEhA98ycAxckSgNC1HNY3bGqU0sbdshAgBh8JME1
UXZZ7BU9HWxEsLTbsCJoyrauIXhwfuFZEOJC9bQlVvY+B3Adlinw9w3MLDelkhdxA2+may2oPA+N
9wBYr7k3dkwIaRbq0mf5HYXII5sm03VdVVCKq5IKuucbfVXbc5p6kfzPJskAj3NLUcqFpxcl3pXP
vx/92wqAXrO9KweuEOJKVmanToanpSPy6LkW7FpKj0jsoZ8/LkOjaNQG4xY2EHbzOn6cYW5+HCLo
mGsr+m4PcawlGAMl7U7HkjtvvjEEcBw2VDvt/wGCX5/UpJ/F83d6/56evmksCrU4bZTmUgFN3kJq
06BwqyWn7yLoBZrEcoc1EUenJEZZ/VQRGuBzQnzV76Au7T7EI5PFABXagO5TYIj6lZVFS1gpx/vL
xep8h7jNiEgIQttatOzstxC93goZMHuupADl8BLunXUjLNinPTePABRZoiyYMQg1F+iT7r4n3B9w
njO4wGROlRlO7aQKi0xCgYiJJgwaSBZV/A35Ybxu26bM0DfI2WDyrFPAhJHVb5tHPYd5omXWBKQC
LRu9Ncu1hK0kOJYotGxKQFmeQKPlO0R95ExOtBo+LZguBk5O5qNt8LZ9CXLaLV+B2mcsaglbM4A3
1XaIJLnRCrmtUTsOMlv3vRoLgB99WBpZCDnDkXIEJZUWQ4rOkyl4o/e1s/awAMfxkwK1ObWqGUME
A+0jojUHS4xJtThjoIusp66zajs3WkSpSrDvsLxU2R/IRkCUonXBZsNh5hU4K+ZGSr5CBnbOVkWi
7AEP2F3vkQMP+g2wiIBWTwGo/oTxWO44qt6UK2+dJqz0ql7TtbaFIQjGPRA1mlM3rLVDp2ekoEf4
6vB50J1fRrB+r8NHAz0fQNJ+aAyKGHfWqxGa4Y2oNOYQSFSl2KyXsznCjMBeJASwH/jeIvW9N3lx
tlDhfGWeF2BWZU2565VnNB0upjwGzM/uWCz/OAq7W8G5gP7+ZyoQ+QZHrJN81YEbeWXmaGH3kzdr
2t856z42Zy87WWceLifQpyBlU7Q6//MMpdbzRw3nEsrAk6ytNRz724h5Zqkc2Yd8YGilRzTWc6lB
atGL7D8C77+dnmaogANBzjPw+u2WUy9cmbZoGnxzORYy4luNL094GmXWEoq3d1ENYr9qWcTLpOiA
GMh5ZBPgLC6T5BMB30oSr+01SjybbE6EcRLGcaP+5CM6LGEPOdUVKSXhXM7vrIU9AazqaSymjDqI
mheYM7TVQRgtuDEjeOO+nnWG5HjAvOYkhWxKrsJRCopIOCamSfreN0ORLHuSi0KJPg99WNcLPcn5
8ty5hDdaanAh8PFUfOuxM72KS33xnvbqsz2FRafgAUmgo1Qd4jMO+fYwWFO4oG3wrHEhR8NYiGLf
H2iLOCXwQKJVqLnJbkk7V8Eq0FkF5coG+3cm0maMNl2mK/lUAtZZJMAVqWAoKvj8Ssj5WdHmlGSs
R2WIl5dW6FVCVcA4U5Jv5fgxUbcqOhBJCvgiCq7A+cfxCJGIw61uiB7aXzSVa7mQr70PynOMxkUi
dG+STMUiQyT4LMeRtD0k710YsNqJz+8UOckJDns6/gdoJp32WZnpGH856VO0WZME/xQueyTH6J1X
MmMDde9Fy4svJsqlsGNs15+M3BLDooSU+FsbkHXx1IxXVTxAhUht4qD0KBFpyoQLMX62IjBItG7w
u43TMjVlifna9CVrSC/JprWZA/I2F+NdV8J6aw3rvV4lZEHAEtnU9WUpjhWwJuBQ0cdcUAsLZxsK
yRN6BbBGhBuKNxiKZ3+IsRrDg97MMfmpBrIaJtYr5wZJTGEihjXwIPifC3s8BzlRBNuetqsGyBUL
ZlsIQCM76SYh9MfZRLfgxtU6eFRDFxXzl1lRLmWw+KtKBWZaHJXd56IYBAIaNo5dgyfLzrGx3g6M
Q6i6GqNgOeNKfO72tBw0799lFkjyFQbUNjIUze94vKU1hoEOihHWy404TXNVwGFRM66+71gznNhL
WXyAc5uqE8gZpgEG8WDxCGqB6Vc8HGFzF+3t3YePNijCeBYR7jWtCqDzsLce08OkXYoGlo6sgp9E
puBtj96pqWjnQKqBLiWCapG0L+mcWfdA9D3zs+dJk+6h7l5yhWac1n7LsqP5RqOV7edEujYrR6KM
VXjcEPsG9p2dBMWcyuR+9RmG3yVjVobnMGuDVsKinLQnDxXd6P1gQUaR5xYjpEsr5TOyLq5AZ10G
cJcM8z202w1irWNZ1s7/6k7sbVOgfnNAFLHHvLjuJ7RPdByAjmSld/Qyl6q6LVGOpG4Mn5VxgeXW
fanoLHJS/VQIV3cAxCYw/ctQQKAymTgl2lRTSsy5gT7uID52NJ06yrKrBb02pPlDnGDbFlE3mB9j
sT8NzDaEGcFPhlydfr/drDleTa9eB3nqSg6sspSxl2E1YB39ILoH4rPX2L3A95Gxv862EPoMhixh
mrsdilCYPkfUPnO4sxZ0qZe7A5QwOKyANFH30LOxlkI9zkXHGAiWzbCMDlCG+GswHROvaBV2AYH8
B5FUXGzIWQ8zLb+3Mptu/OI/BOkQdwnzEx71GCRdqpw0wTyKEuJqdgc+5jJbxC7Gdta+BpMEZxz4
yivVs+g8TjVyqhbANfLprfNwYPEWDi9RULG1zxKAEmWgy3A4BWRU78a2PDbWbzzif2uAy3saTJU3
+iw0zS6qPkCCccKFZgSsWNTjkVOU9fAk3R+0C8go/qHXQ1Uh/csDp8zsZ6wrNQ9NmrpbqdcwizDQ
0k9Fqu5Vg2N5bWWm1QwLOA6SuPkD/OG/lwB2QtRpWgt6YyNhHJXaCmMUTb/x2FFWhdIGvNPv90iS
popz8LOod1EEHF4Gnxp9605QJt9nVKCKRZQDqGxAPm5zgLvnRERUkfPkC2VzI1aKlgKRYUjYfbZc
kYZLisvnlVbfcK+oDIdusXIWY2tUtIvLAX/dGO7TGbPDd4IxYcQMTdLk7IPwx6zjJunm8m97JNLf
zQXSUoK1ozdur3gS2vqmwH9ulEWaRpoLaLPCuSj4Ke833tkHd1JR67wFmy1v7abBNSBj3wX3qjn4
C+W0A+qF4nUh4z7mWWG6GGYxdwOHM9QUXtwMmCZ/cORznUkiWni+I3+B3W0Av/YzfFG7yZRoizzQ
D3fJEa6R7Ervkri0XdwpfCgT8O+UsIEpWEL++UoHhITluLaeMy3M5AWrCu8ABxJyACkK+d1Y+tz3
CFCVvFoF8C1bpQNC7Vk1Tx/jYc0/C+ABUFiaSdF6DYpOe0YEzkVWySsuE+gHnq3dgD6V41lMWFbI
VQYdqE1PdEeXymbtAiVmG6MoKPZmsC1Nlt8DCy1SlghQnFJubDZjKP6CW/Rds2eJ6ml9hQl9A83O
h735g8FypkN0OixyPxHGK6OF2+tEJVqOFzkcDIufgT6uYJnuDm+ZXt/B410mWIoequJcAq5cGs/l
QxYVN6Q1FT7z2zIdCj/1aywgT0OG06p2dmBrMoUqMumuo3c4Kb1bGPIk0TCTjgXa1RTNCxaYcy/2
sp+Lu42s+y1bN2NvzuoCYf8zAqvWpm0aezFo+mLiDJvlpUwEfPt+SB8LWT61ZhOzRl+L0wtNOAWC
zXZoNlIkDwwOIlBxY4UR+cUdk92/e8DrWGjRtePCKoJC5+NDbzVIbjyFYrQmOTA17Cq5gjqH5iNj
HkPKoLdhJ+U8Oxs9Don7hRKSQATS5IyTfFmg8klpl8yUlmDF3sb3SapFsDzKNHi/x7zN6kav1Z1I
MOn2uf7K4LA9/3SkhTshmBxVPmDlWJxRHOK/iTNkb3SaIayy2ekdSgSOoyKr2exB+i/x2KNsXymK
ihRCkae1JkbzKkIREK3tsyvKHL1jZUrtudVUDIpLVPw1Jd/lqIOGG+8MnjsFxwB19gYpv6iqfVDf
FEEn40DjowBKGnphi+JFArGnq8EEkRJX7g0BR9TNYjNhqskixzbfPcVYxSxvzZGOuHo2K8iL8SR1
cJd90fleXksGgRLIEsFM6Ahjyj6ZobcFNwnZJb8AipYuFcH9g4SIbO/7W2czSsCWjzoSBGUNrRLx
BFYczuCePiVC/6C3sy8xz5giXZl1laN2vnUoNojL6GgaIvAyr9DrD7oRp+ZXGTDltZOd9apquxG4
kiP7mdF2oO1NxatB8tntpD4XmaTnLniSQv0eFpj9glRmzHmz+QJ4z+T0U9L4TcsZvg9AOQf8HfHp
QaDswX/n2vTiwx1nf+vpG+Lk6IYETgr8+d6GsMY19tgFJHRo2fJvyAn59vxnJnVDQcaGQsJ3bmTk
/ocUVRe4ZlOEcOdnhzTMe6jNbcTsAI3lWdwYFytCX1YtOmzftwKdiCzJW6EUnu9wgnU+Bv4xQFh3
QFTgvk/r9AS3TbE53cR/0/NEwMqG0HpL3igI0l3Cu9SzglJTb0SS6Of0A5bQKnl8rPicLw/3Jdsi
H/oCdk8qsvfJm9F60EigQsHDK3H4bhahJpyMrTpm3SQn0MS5w6DO01/J8JseFRDa7uQpBRIUB0f8
DD55eqBvVF6vgDkP9lOORLGGkYwm+U1H9UoQN0Si1YUOGxAaJcL5SClAH+wUucdjhl8EJNf5nAwj
+LUOHdPwgUQKv3HcojsqjkHgbAVCo+i0LPH70o0TuFS1ryd976CbEkQKo6FS+USAF00f+MOs7+4m
KoM52ig400Bz9SXsJGpFZy3iTe7Su1mRFXHDAo2h7p8xtFPszbNwTq19pjMdg37amlUyyHDnweSv
lR4cTg/eaGLA/y9MEwMfaOQm8T+jLOHssk3YJL4goys/hdiANZLPPuwC4lUigXezotDHXyd0cpkx
ibNYCkNVbwB8cMGpT5YhrrVCPlCx9i/yMgNWaSOkbqcUAQZHBp0svsiXX3Z6vjGQ/LcXMZ/tNhoD
bWK2Mvk3h1f87O+r1R1uPE5QUE/X+esX7aXMnc4Mp3HcYnU5fcgXqL0xcseLE1o9xR6siYcrut0E
0FpuGCOpg/IwaNDUk/0KmMqPemkk/UUqNpKcIuQ4mFyovqXOAJRGEDLCb9qGwAN34Lj2zPi/dQJS
keivjRcPOs5TBfCFBSPGTV9zO9nCq0NTjOljEvE6SaGttMcL69HxQL9nZSxDhs7ORimvD3JiXdb8
rgF4dcnmXDIzExPuxU3WeQs0up+/l8OGojRxgdGCPHJ9QJvgimvfAeerNwdmoxAnI7PhOAeqVrzl
RVvnc9YdmxDbWyKp89m30EbrEezgFwiZ6j6DqOdcmeoR9AN07p8Hba/Oq/SvDjruI3lOZJ5ZkMO/
8rYYrdDLy1r7QpmAzfjYzhS2lZyyJqkkw19b5RDpA/cESHcoS8YU21c+xhitA1aAGmrkSOdQMHzO
IyJp4awCFsnnXtISaYGr81jstTaxeTghb+PyMY7sOym0ZyGJrxYdHTFS0/7dMFYN1CuYvAA7TDM8
CgYq6LM3NMoih8Kvbm9bQCUf1QyNWl1NwMK+1Z0ykZCm3c2KQURTknlucvSQNsn0rAaWuHDOvyMn
b2QRdo4tGTQ75pyksMU5ik0T6JvBBrkt7XXO2NWqzD8t4pguDLySl+bbJwQERsqiwoznSOyaSpS3
OH8LwI837o6WxvPLZHXEvXreoN7h3BHeJLB3dpNvVCDSr6CM/JaP3KV/VirKHDXS4osIEK+XGBKF
TOzUZz2NUCulA5IrJvO+lwCIxGSkvSrXMxXwjfH5CR1iZeZLrcCWVcdWqHjj10f0WFnU1EquSkHQ
+LI8DXKTTN8GHvn/rZe9cXFybBv1b5CNgzURVvbjtVeqd8iFuseXejTi2snKT4u6Qs7oPOsqvjbR
06zCf/yunFfOS4bGDCJf8J/ahdbxQyEV4/DCg2Xr4GaLiDDT27cJk/wgw/2IUFOfFZ2OR8G6PNWv
X5Qgxt+xrUGO5xrH2R+yMPLojc27y3NBZi35tmxrPgprMkYuitzW9rcbqe72Qt55ga0hEETpXshF
Q4kmAgy1qiEj8zmnL3lKiNy5pDguvct9PdUOnxzquq8VRmGfuEcbV2sTBLkBXraDGEgjyb3QWXnk
uK91PZVOPd5aVuzhyQElJJiocnLTB48GVpvXsgigRbOmPNuvG5F4mcSJ6EkW9Swynb36dogbp2QD
ebhQWws6ViGYtQVJajkU5AopxtMbhjqOpNqoNFWTaaixExbwS/k5IEF+6PYEHGANgXD0+WzROW7y
1KNy5e0XJ2IvWA2SQkei7Ck5LnITCiIg+VK5F43AimiaDALXLb6Y5s9MEMt4uChhox7PwponnYrT
FfoO6IQXifF7EiLQsjrWrf1qK0urmc8iRsZmv4OmunMK8Nweu8TMZKOO4zTg2/+ITV0zxZFP4LoB
q+hc7ZJV0v4tOyopgNH1Io3MPu44vaUYdUUmcHP4eLj/8uZLBQ8SxUStLPje0aZYbYI+H/jzlsGh
7U2ElvB/960d2D9hUUlc2q1Tb3M26oFry3mDVroIBHApKmZKIDaPKBY+hLOppqcOcGYjZDfofzj9
tZEbeM0CzKM6ztRa+2j+j0QYf2KOHxJ3w4OCIrWXpzrM4F49bDpz5jBPdthvVh9bLv6Qufnu4XWy
TZZacGHyoYsy7XaIw3PUBdHFH/nWIM8VBnRwrB6K9EBCYFHyrsIRILQrEBhipkPQUiD7iOrWenH9
5/TLd3jXSLPmtTXgiPMLyaHcWZQaJtyjvZiW32uy1ZYIZqikm0TrmXv0bvmhqvT5HiTODS7BQLva
WrIG+etMM9/3J0VYQWjRyrxaIePSNpVna3Ye/iuK8wDizDIr1DbZFKOTvvqVw9OCV6kNz+ZRzYu/
tODk+BKVIqMlACOgvpnV3NrCqSBtC4x1T2Ksr6GNNTYopR8w5zH2+2dHhB5hH8TWyv2Xy0RZJDy7
wwHWXHAPpj+xTjsItUK6rnFe/rF5hQtgxAau99kzCWms5G3tsWvAHGcglMcmPQwmDDuNI7/DFhdv
HGPovVDKrnOhNsDchXBXW+3ysWvBCKnEzf68ghW3hV0IRKwD3rnAzFqD9UciCaAUSzPIz1S9XY3j
fYiElVhdT7vWPhWq40v8c3VN2Df7y5eTaH++cORgMa5DmtHopVWpCXm/DJ+W6z0+snub3zp5SvYg
uZt/n725POIpcl2Mkl8TMbNqWPR2ehSD72mfoQCIeCQPVMJbPxR9maixsm2DN9nb9SBXLkzBYFka
pOYyCNIDMVoBK6J2ZWTlpuDlhXOv+CZlw5P9bjYz9Tu1jvO17MIxvvWralkKgcdSctCBubntiHay
ipN/urA5RKMEdreNf3BwROnrg1GbMYu5vevfTNz8wFwRDENLeodZuZqy88tlZo9+vLeydephLNUe
CEs81bRD0PL2jVPQaZrAY7C8zRUIBMq7wPQbL8QfEUxRyrHY5s5ue5URxCnmXFwp1mWMvfNhSfMg
6usnUqNbZdswQ+09+3VocOzqOiOoTKdGvmC0sAEVkE+l6SkLWC5YeEE+iP7bKQ9fduaLV2NarCfj
ByL1H7ZiHOW5NNTaFo8CuyBFh8It1GUE9xf3NXuzcuBGJoFxPMaABFu/If86CtJs5O0oSmMrvdkI
jfm7ObIlfxYBGlRGrfBGqATF3TxotqsY7EFaTaEjyC0UEW0LxSHVjvkTHywy/0W0At8eX72xt883
vkEcNo90+v90yau3/vnXxFzxcBe2fICUWVAIRxHYsNE27D/Y86UeW0lhPJ943G6mwJWjNBJySovX
24oMvWN5t5vp5aeSE82E95ycjpiQ3CmbzTNtzrfY6kadABAQZ+m8z4gho46LuVMnHjysEUv3udhq
CMGdWM0wtDq3QmoFmR2xUJzz+KoHHSYO0wFOy/H+wbhjm5CBkyvMJ10cw9SHYmM10aLZuKB5RyQk
jmacVq9o5YcvuLJpLyVkfqJEYcaRnRobsi81BfUQkFKqTy9xoE/gBNrfc1Afzz2vw/c+Ks64wQTU
EPw+rnkox64J4o5qsutsebtr8lF+pAwoJkdiZiki+pmowX9oNoywyJUgSHbXDD7eDKTkTDqDxnci
euZH/vftQbmTbkW0yhElq1COnbk7V4P1eg4T0qErL5Hx6bInVjhpydoZH6caCdTEMDut9lhoEA0u
hT52apP0HEUhLUJVshEgryJw/FbupTFMLEtUSqpa8PdbMwspP8+LMQeon9h1c0fwmrx8sF1vBKnj
rqvD1Y62VD4+QA46MTBQQtuvPdu1qjQ/PumdqKQKHX5Wrh8H5kt4bj31sAK03Ko4eLuTdKEuxCVy
wUPjLelSwHzpcpANpLMZzYu+K3/p+87+XruLIgYOb7WHSqwq1kh08GacO9Ds7cZcXDcu7zsNMHxU
bAy3MzRTulAwSlbAOoJWVTJ/0ZQYdW4Eej0NZSMwPASwOI33BHyP4tc5UQIWKaAAqaYygt8ciVhz
DomLiZUmSYLMRqBupD7bKQwo+F4QylV5jDCFUiLk7K5Dtm6IerMEjSrjb4SPrqr40gw7azwtYHle
X/hDydIApOuLvGG9XegEHks7srRDK7YzFFZPcvO7R6USuY0/qchDxVinZegiwbKy4Bh31Z4HijX0
niSkR5WLKN3XgroAxWSZg9G+dlAMNIJ2jk5hqLt8lTSUQ0Gk8OMAlz+Wlq5KGEVq9t1YAwtoYL7o
aqvtntIrM2OSb+43qr44c7iLJacphgDjCB8hEDabXyEh+TY5xbX56saztzKNbfJzmQNE5Jgzj2y+
7E2DcuH2R5nhdjJUoYjvdHBgns5XdTp9MtENyTTOXTyvVdVAFmd09QfF+IQWRQEwmJzi6fyJwZcz
qsuVMnJHBcHC57R4ZsZ7relG86cwxNktar2Ju0AX9KZ6Gyu2s3fhjYODEa4Vk7/Q8yLEc1fcIyC4
bbBkKYUf5yrCsslorC5Mqo63YS2cl0hXKTRnEXVfdktRsy5FzXjbRpEjj5q5kslPLXtHV4No4VYX
NpczLNIs6hT+Es4vUehy3xOQWvuYf+vDZkpww/YnXfhlfT+0U++72fADimrmQr1fXD0vIkFUn1Uk
cXLYKmDY9JKdekM8lF0/xjYiIRYP3O3tKntyLRJ+qjfQkn4363Nal8sHOjkIdJwxUBWW5/x3IXLt
LdCbfwPIGdWeBmZ4g7L0VJI+elJYKyQwW6pEeLkz56/EXRiVHyr3DnQuq2X6O3wLDMWxsaegPDzX
VfvafyzQT2xzN5nq9yyNAWecyW8Rl/7GIYarasDYqfwvp1LG5bs4iapff0/TRS3T+hLdjXAMyioJ
/H7DND+vENqpU/BR9UOytIwnQzk1fD3PpSdJLBhyWEoUJdLzaYFhO89Wak0W1Ih4EEMtYYg9z/II
yhQfkHLjbTCJXFTUEQQzi5C1PYh3LkN+SLX/msetSb5djWuyeXib6FVAyRctSbd49TpYVWJK48Co
21szej7Tj+7wMBOBApJqfPhRDNi8QhMLTiVKqGQhQKwp1GC80UEJq6ikZUyUxaCemJcn/QicLKyb
KC35KOt4GLFQE8xOkxU2K4xJ2LftqFpZhG1ZWA5sR7Oei5/uamElLTo4CdFlLvppiKfVYuGBqY15
0DgBdo/SBy5N4MrbduIYgJMlPFivobDZegTVemqH+qRjdGklSWtIPqgxsZzo/msptVEAsXlhuOZk
/MZZaqe+cj3xp4ATMtQC/pJOSp57wh5sYtq3L2OtB+RCaU+gZXa5G1NxtGlJWakIKCibr6I9xkx/
iKITOpsYinDfUyuWKXxS2f2+alQqlegXqGcX8IpYKBynY588tIj05SzZGzk9dCNSo4x3KzJhXq0p
CIlvnraERPmue8yGWAc5KKoUp/KvkL4epGOQ2SzoZVms9SArkUQrtAaykA4MB77k9CO5OzN46APk
ZbVSpyB7yPeygN/NDpGtJ6CIkmpHEHB8mSCRVlj6MWvmCsiUMiBANvKyOHpUQdnAy+oBLUeNVwxx
999ZCS2hxIIzqJEGY5hRx1A+uT8RAEapdedZGibYkmj77AD3LrREdstw3C3O+2QDQsvdqTNJn0+p
NkkqJAvRUilcwFXA5mrUpq8IiA8zKqM/KftxH6tVCkd31BqFIW6g9V5jz/lfvv/9+4xKrG5wdDsk
WN7tUpWO6tUxwaUS4Of1hnHk8mJgVRcLbrXoidQtl5YPb0qAuyA35J0q2lHk39ga6aLKiotT0Lqi
111komqLtvTrN4X/MaWygLFposYI/Q3ijTGMZDng4Bm93ieQ15LT5MnS882p656XXqZiI0bWyG8y
eiP12rvma7AB04NaQAAZwtJKTbF/zKVkRfZsNkaumOWatShdqv/w1ixEDRAZuJUFXHOeeoTbvuNA
6Mv8C0CM3O8Bfa8AOS8u0AIkjyW0hIWonFdvZ1MHmClqbbjO4vwZSh+BPBVSbBS6ghpZcK+8KQTc
IDxh1q7A0xEtTr6uZ+Q6/jYE5mLmywDp0jJiRyuavjTFFtvz+Ka4XYD+c0HjRjaTZvGoY9OEXgAy
RkgicYkryuV2Zl88h5ALt2zljDDMiw+Twg4iJ64ILNY2ulXCaFGe3Bmf+Up8w3J/leg5Px2AC9cr
n9mZQxXyRZyCcyiqLDuFw/K2GmOFE2WKh7b2QzoY7ij6SSSZyZzrrkGfV0pTTjU38bN2sC0bYEvI
wV/gjUfkaRjkfB/oxNSX/AGnampT+qaKoIa+jmMjaasfBzz+4Ix4SKk++63B57Cu46q7rNI5U4lh
FeJ7waBF7+V4kpthRcWrGIfENF/L96tVhV4dv0H/EtWsJyH2/2GseV+flrgcRcAHLAq42qgJNDzx
E1+yvw3+9wHQOcHZxwebX6ojJ01YH2V5UMoRkAK4OTP1Y3oeKEkrm5owTzZU1QiYIKtYWmHJh9yK
4aA5M8S4ZQhCBfkmCsqdL6du0Rbyzi+bEJ1PJIckvpmqcKsYjSpRLr14ZF9gyRutNvaj2zq32b44
sI6n1cuo9u9o44ClRINBXUgYSe8Ke8dkCSl4Dv1h5tUEjKwAaj6HohoY1fsNJBRTBvYKCwJg9IKn
iThxohRTFCHp+BdGG2uWwndC5iLKzjZXjBsjtl0Sh9kiBG807Z9MskHqe/piuBJqNlXQRYEJ9o/R
9p4dx+ciS3aZzF4Ain8nrfOSIXScvm43gkzRzbjU1s76waseAMLGCErXGEoGdKGi/L2lj0WJCnfN
9SqaRBlnSgZQ122rWjz57jzbDKh7kr9aUp50xzmk1Fj6t9kysuD/Z84FTMolKGHc6Qzh26sQS/SW
/7n+ghw03oOYnMqLfplZ4gYoSqNdROPB1BNrs1f+swPsPDp6TyhOKfzhmws5+pUSEMC0OBCkLwAF
WIdOblUeUPF9iNHfuBZ+nUnshdDWdRboaVYehV/X8X65G+so7QALI6oQLDAcJ6wB3TgXyl4CnBtp
o0SuascX6GLI3bwO5Tg/mS4U6QdnnIpEbOmN20Yv9F9aX+K9HoSDWai7c7YszC7OZnbS7vQNsXYW
ztgbahpH+GLtRKnKRY1PeyRF2mOm0HtqL8IiB/wb1+I4+1czR9s6iltUzd8j6ZHjs6IBwSP84gEu
tAxrNb5a8KmpIXN/EH5B5d0+YykEsJRRC3GsLCLDhofFNpcFJ0+exGRxWQ9rgDH6Dpfq2fy4zv3B
/aUeEH2LHkoVDszOOpSY7PfIzoLZWwzQG1UaDk6PJNBZDOBA/hAOxhniph9Vb10HiKSechwPUjT8
nIygm0RJa3y/ivuVWMexpTct+SrYVgJPYIYxLabpDj2TBnzE9Ya50YijCTYGeDIDz3x6hGTukGyq
D5OtX7afiOxFQpha6o5rYfoSVKnSnGrnB41IDF9gWB8AfXRmda2pivft6kuC6Ypmc4oDdGem8oTp
33xEYOYXclk/W4zHIzDpZ8zIiG3xH/OOVp+bOyuRL4AGDZNwsK62p1E89bIj1nM10NtY6uzacpgK
eVg+d1sN5btzPS6DlzR5Wv+oUjyyS8JOkb6eVu1otuxphsD5CkZADb5rvXUlD78latTwkplWWg00
xuN1VGD+TnjryTR9NLzUBDLtqO23wwKEuVmOYDC0xbMj0NoEBh+veAQYpoLaWqqRaZqaxKsHFIrv
WxiqseLI6+TpsR36sgwqffduiV8NITi8PnIeQSRem8dfze9t8ZxlQuHmRLo4fNZ847svYtPJvwaT
WI+fK8Z8IXpA5EtgLydS0ltPwv5W6zEzYYxx6LLg18N5RoDZS/mCK2vAVEsjzlfveQ2vaQ5elGC6
ZkkMBRymdUywbr/myjNMPhF2txewsXZysPRAIgAZyItNZq53KOj9iuZSzO3Wg8NV12knwaF41Yix
c01Hf0FTJy/y/0eFXUfP/6TwHeTR+KZir9dgHjY1lPnLZtQE00viI+D3F3u/YN/MeGt5kr+3RzXF
J9u6rmUmTkyNieuxo4RbXILl14Gm0CHNFMz53kiUa4tlY2PJSnMKaWGJrMiVhz8QjR9Ev8swWhOj
xlrHcF4KgQPJnJsCWmN/w20Euw/zFE9UCRx/D1O+0hfkpg8tE2G3Wsb1fO/sIXz/cakt4vzIK0Oj
DjLYnUHikWSy0tjKrSYofDqz/EDXvWEaR5QX7OfAgadmII2RHugswul66kRNBCokagYENyNlmIwY
NWSJhKCesJJLQhk142QZqx06Weh4eM6zG+0KsB7005xmM6mkAcr6TAn4+I3xrsJ9+JO/YR7VPHA6
AdlPP52J2CuPtQ7MV0Gwi8m0esTKoNVA/ov3PNW/6MJDXC1f92r8AfoUeHji01gIrZv7WPN689q/
tkN1VZ+6eKMjbp9upeDAS01GBO1eQAIDAtpAWTHNl23efve8IGIyDaPScS3zQ1bfX0sGUfQzi5CV
6en/2k3g0bTaaiooZJqlFrZmg8s76btWC8SZ8nIhD+HZMAEMriwuT2tkgkuEcaVOgZhN3NWNa3Ha
J6Yyc6OO0plfwbSz1p3QkqVqBjIN3ZN7K5Hrfwvc0Y70Gn9VVSJ63Lnl36WVF0RO6c9BrDDFBozH
TsC2d5boZVY5iZwCh0aWDIHiL2JIkP+LDVBmCwbpH3Cott/XX1U/An/7nvsmOzGQoAE1V9s91fUe
Wk+bWgacb+///wkaSA73jsdPboRqdJoT5BimlNHhRENeqonaVYkMW+4tu/EMetSdWvJxiA0Welwc
AQKy3P6WqRxPRdv6dBjFR+CqU2Ar+XWlYqHban8YaegnYJIURtZn5ZoIx9yIg1CI2VFhm28BbMgf
neNzwYsZ4TojpQW5auF7sgaMjc2WpRDBMfR7zr5TU9fW6EkSB5gyNxX9Y5Hs/96hl9S3oJXtwLn8
cqOHO2ro5UUOzLHhGPCq4JNqHN6Kjfl4I/iF8yf6Jcwb6lcOJrqzrGYcQDQl5LMati4MKaiNi3Tp
PEo3Dc0VVQnt/uZLkjFbGyNC/JAFZq8p24cUWwrvMoXNHrGMZEKnKmZRfGlFEZA79+0rfx+cQaJh
+Am/XXXBMCU34g6+HD44uIUuQCBAUsUILq94Bv//H84v1Owt/4O2wmRTFQPhe3Py/LlqOA1DzdMq
DqTEh1aLXsadA0mX9f8FgeqoYAR/ujkJkAcK43Au1c0Fvdb0dtATigdHotNu56cKfa24f5xdBXcQ
O340oQsfuyGRUJ3PN1g0lijWoqWx+u2/HFwxmWrbbMdmPIFc5evTnW4go7hKEVv13Qf/jZiO9oYr
ug4Q/M5NyTqJWhdAgoWfAgxc4D7UvejPgbC51Itz3ReIplwTzqW+jm6rPc5xpRi45xo6U8LpT+UW
yZi53bu1j5FJTiv+zAO26IjwGZwaKTvsSKJMp89wgWe9Fec5X9l4kvkl7JeRccxYPSjuN8LMEK3a
RndCQAfd1YJc9yTW5MXNSVrNVFblW20axPaDPR0fQit7gNhyrG//pzPJEhwPu9rNkIj1Tz8sO4C4
lToDT+IoUOCsDRTCiy3AOMLm94NSY+VJpG+PlcvW8goWmal2ObWTFH3ljZi6uxc68YJQ4GW8QLxH
c28ZKg55NVejsTqUOYvk4XFdRkrfQBohGWwRdiiUwIVYD4ZUlawwdOPgpCPNtC8cTQH0AKpkbGPG
lJ/bTebluNOtrYC13aobH+LiWQ7rjhmEQgvOdgFzof8JzJCKhY/I7doGVBWkCOM5qkwqTozQREaN
NSM7I8c3CpJHQLvMxUdfWKQfkJIQaXHGeRT7RGSZDqzt9N/2JW8zJ/IblsRVKfXA0LPRr+/6Sah8
EByfVVx8WGgH3b/qV/RbyR8RPA/lwjxaB/Q3OJmqi2J7J1bd8HTpUQY2uNPHy6aKa1zSeVHsWKJx
d5Va8gxRvm6QZi/bWyweYCW630FyfhIvlepbZnXWCHOPkvqlfuctqt7S7wvYGqQO9BzQ/VxD4NMy
rd15Te2fu1X0VU31TOmQHdNX8M+Twznd9/bXx66NGpihlV8LGueol2KcYm1KpEHEl1CWjMHGzbjs
ts6cTg4C9tzUxbyoqveCBL4U99SJtt1znAAJOOxlK7mp3H4cxhWwKQQB8xPrhRI5x74RMpencz8I
5IwbRTevS+ityN4vt2HZ96FXQHZwIGJxr9iyHjsKNLBOuie/0V2Ne3Vi/oNG4Hz+0M0QNWdsg1z7
aIiKrX5Xnc8RGcKeOl8ZUQ5S4IlArG+AtrDuwGrHh331cgpWgErhKKgkQWQWx3+w2U9NPuK/wAQd
g8Gs5o3mjA+Lha4HiN8l3QK8ovDuSc6k1C8mKmE1Oi0MdoYjycDfknIVjvxw5J33h5EI3sNeGBhG
jScXh4SWd8qMq0es1bHRx8+BmKrAgJM3PK0xcB4C106nb79Pfq4c+jryRxVfKOPCpZ3pH+ul1nXD
XPTH4qREp8Fq8MoK+/Yhd7w764qyhZ+kjlNq6GlbI4Z80tl3ZeNRRwoAaloE2d3BHpSmeS8hiUI4
kuZEsXwVi+++tdylkd86ihwrLjK0mmdp46BS5EKqbAZJqOmigN30epGvibZ/obemHELCAu2TxCgk
/PhpiepDzm2g3OS7BTk55Rq8VB7oBo0+xTVzq0Lx+OCKZZPABfuR866A/Z6vSxtgZnRAXVfpiPc7
6+H8GpfALu+W8tcK4jj9rhWx+thBnj+o/64VVl4Q4vnQ3hixZj02ZJsMoS59Wh53tCCHU19AuYgD
8jMmyUdf4PsX1a97ThO7JrwP21Jppji2srSHqHlVO9D/doHS1TOXSM9k+dSH5MlpIkfS2PJ6+mzJ
anWa97uOv2QXPJJtQKAAW/CgBVDslFTmHimPR5EsxfeWL9L6kge09UCtNFQj7zw4UsKDq6YM5VM6
ATo1nLS8U4ppb7U4HPbeBM2f5BaufP4YSPeS790cDx5sckt2Ng4qFQ0E/VM8XNFLFwv9Y7loC2vO
xGSVqe257TUFCJPeFVE3Fti8A4nJm34+lQrguQrTyPUxMOaOI62mGRenPy9wHRTqT2Rc+1AiPtpH
HwAO035wWgzA4jZ9fE3f6lSbkFIaqH0K1HgQwEAhS+rg53O1Z+Evj7sY3YCp4wK6KjMUyjJRvSqh
NNSuwsBRh2oI5rI0p+8P0hCTC1ykhmKJohJfQamzNQGBIxMb/9QIXOJIIutUBq2fu23UXItOBBb3
A2PQose5EnDUDK8WtHyyVDyVDThO4mfHS/nR7wEsQwsCphZoaUyxwghBgGpEh/OqVnAXAvjd8zk8
fJg3VshAabjBuuRgfOuFNZb5OA0/W4gosQYmXsYfB9ubzpxPyNXTU+G+MWKy8zwg/ntan9rHakG/
+tM+LoOaMSwMzoukBxh98nfDOCUB5xYdni8en8z188MLHmwwX4ynk7eYX18hljV2Zw5ZOZjSC8kL
yOymNsgev5FbOwdh4cMCGwPSklkcg+BZGXybedM0hxDQiG1ltCXpbcPSHvTX+wjUN9hsaDJDxAtZ
cW++m9ZjgFyTXfockTSTZPhW0+4HdUm7Cz71RN0hTR/x1OywYOIi8tmC9HD3w1bpVb3IVlupqyH8
96ZPu1UiOKfVc9W0wIZhlcywEq5dfX4Qjez/EJ566e2M+TqQF5gYsyb1yxxMHmohLoGHTs74gap9
nJ6JtzA47mUZk0yOq6aUkxUR2XHm1luWFKxnGx1QA68OpSoMg5/skfrrF+UMDzOXpPQC4KgOk8S0
qyokxfdntlRyfVpdzgweGXb87FtyRDKs6CQzCovmPhjgm4K+Mo7QpHnwghkOfdGWmXmXWrKj6oMw
119u3zULqGgBwvQXa5V5f1a5x9NIdZV8AMmuxDpYa6RkK/eU6Ug2RC5mJnQoL65i+qG3YBBRRHSV
UBSwS2OKpwWrIT3XEPbzgq3DearRm70WcjFX88GKTQKBevAHjrAqx7UIS/S/WHSUKpWPt4kNyxIN
bQuYtt4JoRAenfjSFczUEXklv/ioki2UUFewT721ryrWAXZPfGUCRdWvrMHZf18V31R/kM1hvij5
+UCMdftsUi5w4VfUAJf/zw2O119PQXB3fYcPauVNVYvp0qMU+bRLbuIh1F2oKjwqo6Zb5t/I2ZuP
vAOofBkcPJuNzpxH8Bk66gZmHu6ij+Klxmyl+/dqVhP56ywq/WK9Lr18nSBj6uVwDTbd9bVUOG/j
mN2KMYIrPQ149KaGDbBjDEt5Lm851W3fqX5hHTBbQjqnc0nquo97AT5O3WAQBGb6ZoHP9CWuRC1i
Gnwt+qNxhFoCRVoITYtuMRiHC7Gjd1j9wq3r4cr2pR8KowCbaO0jk9M/yiWIXZXfLOJU/MJ2K6iP
9vvyZ59lvSWZERcppvf/0wJAWcqwCif3xNQ9MN/OTIX92VRG04w1CWlLNPde8Qo2ft3qX1Cl+KeD
Ed25vmvwWeDjrC8iafdeg6Av7k1NZ+VUwcZJcTg5QOAX86kapd7I1gZvGp63kHNSGB7yj6kpVCBf
ZXwGH//UsyT1S++IpJfRGWITD2ncpmcfG9W4H/2H1cT3oqyMOieVWGrVNUYAhcfBb8LI0W3G2tnO
cGx+8k/51c4olBJ7//9SepifFAIc4j0tIiQaYW7B7DbJjkc/vg4qf5kF2c72RkOaGxABe8YNBAd2
diKceBLacQegMemUBLsbEOJ6om0izob+ma29GN0iiI7cKZSqJRFgyu8+3WOtrEdm4UOGpsfofZjw
5ni90zzsV/nMaK6RxHBv4QJgC+6Z0wgcu/SpiHe/dZ1k66OisXTC0h8U+FoZPTYKCSJSpAUPq8MJ
d/8x3hB1Ps8FeYDlt3mJEv5obkbZ89nUY8JpjWzFXlDN2knCweC0hQ/Z8Qp1yEgubQtF3Fso/NL+
daYWj5rSvrjpW4c8HY9aCTiXBy3V5/G+gdjPRfrqzkPFeIrNwRtAIox3fADNzX+IYJVBRqN+YVfU
2sTerETeOWLQoT//988PF1/HRipZtWi3OKVTuqOGlnxetqaaJzU4urRN20paF5UPLpY3Kt8GvwfJ
rvYGv3M9nAIoXEtbREWdSN7g6W25XcLdDhRjvLLDHrV9nL3KWcXTLhjnqC51ZFDi/QCzr4X9pRrg
t3E38iF2RhqjRaKcRLuqDwNpWpV0n1aq9AxoTTTpGTKDcgWsn5rMsA5rM4t+evJOOj07hshJqXMj
BZ99s/+OlWA2qtKoQCf3fOnDACC/Cm2IrM1jYVKCec+uLX6GeKOPxCtZJ7t8zGuqCgbfuQXN4F7L
/o9z4gkPCOHJhESC+BbLHA1QoIRmACRtjY/+sJ9Bx5oktH0tILaSPC3kleImMliZaPUrYdecGAXn
yq8qQAdBvQklrXEhSTfKR0Xho1awb+2jmQykpFW60205M45wiyii0qiwRSwJ/7Y8hxMAVMC9bygN
TEcjVi91wmBk8xu6oz/JVmmTJ3KJwtLtkj3rGA0/uFwlL0MUxwWD2q0jt/8JBKJoq8/oX1bG+Yhe
O+nwOuJamQ7BETKQimvV4E4AetRp2eG264mAUYRNKLV0+zDr0jfNDChOMyk+4fK/4O6YadtKCeEf
2bZE5SaXp/GT7Zd43r1U3j0NDP8zPzRTXagx6Nm/U0fImYNP5F0RPSi9fic/74UezPkmiNaNn1wf
ScnCo/runkuWcolguwAwb6oluoVQ4DoWB3oUk8kRDgYi+IYbpskMXws72BdgvvJBqryPOJzYXaRj
Kr81cLDW42pPzgB6YqdfEz5FDe2Dn8SB5OVWslVWiaMIK4xClc0jnCC8mfw+D9Nod7mWybpJ++iD
E2rzpJjo33ZO8rkQQk5Frl7PtPziwOhxnKCJnNH+XRTokwVZVMVIYAVAbdp2FNktOSyQ+is2Ixtn
LhSxq6PdkDQyTNccYCtF/nMs9hBy/tCgAiDRtZEviTOPpERjOxtx/y2r9XgbS4g/dyh3k36DsDqT
R+R7X5cA7yubOcZ6X39aqr3gDqDhWmKhaeEWT1fKPukTdZ7Ns3ypnyE1xGU2d/dUrlkDrQGHvqcR
SkKxQRGpfPVchokonXsqZTZQ5ZjRoQ+UQBkCes0MhnSZcJtCUPTxHPfO0473kg4cfO6Gf6WxDtZB
JqVs6HIxSYjptC/ATUIpDiaZVBouHMEo2iA0XQY4g3KpckDM9RpcruR7CBr8dEppVOUhlDSFNCCY
JUsguEvFdF3x8kbtESSucYt9Jz71Nm4Mx0B1TxouiTXvtjYsfSdujikZXSVua527DI5zPQdvz7S+
2ZY0LLj+JImR0CAOK/SklS+1Q51xNxEaAvvNT/EXR6azLSEBEYfSXpc56uJU2MxthM5o4lzGelUS
JpUP8i8eS8Ub/VxgHXK/e+wTguybZy9CC6xjdWaGmR2JSdkszBmvIMe/jNSRM5iC6VXPEeDs/FhW
IlNniRuZ9pnuaLtgnN6XuwtNuiOzUVP28IYGeoVtVop/jYs2pdAErI6B+eTQhn4PGMkcvHMqY+bV
oIoDVBp9iG8OUaGK2CKuhnWu8+9z0AO0Qkcjyng1QpPlH6UWlCfJ2YG5RsyMmjSKdMqCVw2igW1m
YMd72FewWa/m5ivod6/Uj+pEayw7AOAFGKnKbojvM/MOBx7j5rAkhNftH46Ck3dRlNgOsnIDA1O+
yr8lM2V3hgXawx5IID/LoWMIcSE7SWnS0m0cQWzYukUJ92E+H+7wr3+wagbwr126MVixjiCb0MxD
DSWDQGUnS60lby5W0qm7fWW9Pk2t80GZSxkESKW9EyJ6pzFuhwiDaBufxvvLd1DhdBTojGTl3bVq
/G+NhuRgHqrUf4gOQA0sFMQnUBONGRO7Eq5AlxHUYi3qHo/bsX1HlQAtNSiLtufIaD5zFIr/Dxjg
XU7WccMnc6Ucxl/jftEc/xSBmLG25LhJQ/3MvuOoERcskZMNgVp/5Mn5O8pyd8ydqGaBu3eotcoH
9ibB8sasyCbOCmDhJeOVJ0uIVqY9uYTgN0vNM06czlPR7FTVOJq1Fr9HQOvGBCV86qpZVQ0ZIGpj
z0Im6268PRA+mQX5Umg4TL2arVl3SaG9atdLB5sV+9Xghg9hbSN/3+Tw/NTrIdRkBMlCRM883sIP
BAFyDKvrK8oCaNj7EVUEH2Y4qS3n8+ebE5b7FIcMDoc+mtWIPsBfSo/EiPqyL5ETSoJGDYtTz221
RWktuL4gGNbkAXqjtsVGFqCIFtaQ6O8Q/n7pRvXmw4LIgtbBwlPQxA9u0GtuITp7TemOuJn40Seo
ji0UBUoN9pElhT4v9ptVRWLAX/CmpcULB9Xas/6R+0Cl423Y1cIpYLGLtv43luDuBp3ZTWa8kVB+
trSH8eI1yjI/Z6Pf7JxKI2vs8IetD1t1W/JN8SSgVPhrvtnkf++3fSNN6p8Oj/Gq0jEIQb4SGnQG
/4RNRurLc99Pg96yNb06UHlK+xaFq5bDSU7Re9/qc3OoTKPfzAPK+vsA+Tb/9NUTBkhbddJl0uAR
5EzEz9p/zodINBU8+htTfTD8b22BANO2Hhs47+Me5GzFmFoOXGnW2SxhoRb2jpLVpDAmDdrN/gis
saTfDUy81W0xVVFHgxP/xTmCb7Z5NcySbJgy0v6CmVQBBQ4UouHxauVtrMZkOOGVVFKRfwT8i6D5
7rGg2dta/wgX/SAnQQba4cJLgUhKbojSW5rrOPE/EdIzxnLmPLwE+o9iYGXUIYFqxThMbphog6i4
EdT/AhRXl4xIn81yB4oRH/jgq1rtSdz5cXDcZqKktqcRvZO+xiOHwvsSBxssChvPCFABbLz+QYfu
5rbWt8HMsJ7NM5qemMDW/7UuyJuAcNZZAXFvUp3vKBxaK94XJSBI6qeJUnrc/v2ZtK+SHowxvJn3
NAtLjlFUXAQG6J1yw/aLArQsDwtAT4eJ2NYGxddbvMYKBVvtOWCjwQxcDyMr3gBaQicJBwkases3
DcTTksbzV/kaqYCoIlGnpx04pk9T9s2/XoPLXASPeJ8EwgA74UtqYN0gRRB84dW1q4Zxj/n7vWM0
CJws6L8jVxHnjnnqwaPHE/3zMMKIPlWJcVS8/Os+xFJrR4F9YixnnYlbjRxq2wsMt9fjuMOJE1jt
ihFsDUn6XtwhxZy7nYIf/OT8OuDN6CgSMx83xwDOnLah+MoKTx8nZ3skMnQllrBCcopCZCuoISc1
ch8u7rU3GCiP1iiB5TJXmJs4z9jeDUTSTQB00QHK9K9VFokvb3yFrXuZ3xmDTGYMWluZ1nSMEgto
wGUhMRfF5HjZbobBFAEIUXgW+UlOcrEHWEcx7DjZbgQUxujxxgSz/OB9juBEH08JJuTY1d4+RySy
y3INoJtKDWQS6JHnXTZB1WzG+WIy/5lb+wtshsscQZx2wfVWhhuPbBhL57CEZ6JjGbS6RRcGRQBU
uN2Ti1twJ+BTjxVy5z7oF9ezIcF7SGo8FYmpz1OMTmutJkDmZKh5U0fOWo3FlitSw8ymOdXZ1k3J
INbbNDThWfPcmyBB74HAdyBZFYPD+ZxSpF9/cOn0D0I+Sq3prAAkmUAQAkXLSUCmO2p/3K8Bi088
s+4oKj8pZeCB4HUjUxEfnB9vjq8jxQc9odg6XKGMcwufjf4PcUA9206kaGtld2fGWKAARfIsFWaa
qBPoA8HzZd5RAX06/B6QA7tVYXweNUXGfYcAwlV0GUYB2E6M37ykfQJQG1aexCaEYKyS1c/oI3st
K6bOiZBag+QZn/aew+7CU54WSJUHnn/SoSCcEv59Cz5yOSqrFsl5VDq5p8wP1vk/8pjlPia/qmv2
N/0aypvV1pvA7MQfJMaUhpQ3JMS/phC7/DCAeLIviMyajRvDJIk5zvcDE9dKagz3JsebOWJ0B2kd
PGOF4DhXTqVYtbEKHe7hRxmNMorSiEkMcjIFqqxzAKvWHZBCLS7KglixeOmM5m4Aw8vWVVbmgWH3
OCTV1DiGVI9SyUdNgzrIWmOQqDmPWn5u8b2pXp9fr+OWnQ8qqB26QJFe83wFyX2ZqbZ4RqDKyx1d
+M/E2kgsRN/PdbWPyhIp1u3GtGwVHxkLZwXjfMIfYSwFqo+cYYYbiNT0dwzwABhWG2Y36fGzav5/
EIm//Qdo7GyKwEYCN6OThAPL9QZozGS6G4mTLxGskl86W0S0Zq79hST7ktZL8UKP3a/2NMRxAXJi
wYCPRdKLIYY/m7aDKJrzFNJrGvr/CXK4dUyaxFcsbgRlxtahWGYmFDPUNZygdBeLP91XnYFJ+YWm
A0aPcI2Hu+c522rb32YX6yUDsTyeStvO6qxRVTn/qH2FE78kZLOqRliT2tmwy574GxfTc1VXVSFV
lKhqKfMMPcRO6BwTKQg1gq8hyd8uvgWpB5envLwdh3p5IamLtagg7Jf+tuLWuv5QqfucbydLBo3t
92Wa8EVrryi9UXuA/OpDYwZfFdozk9te0oZsExMzWi3VHrXlBSX3JJCYUuj8HOnFXnCTK+T6zsAu
HccdOwTXTyjXXqszZVdGsecmJsZgGXjjVLXgZkfJ5y7Y3gR1HikPwogBafErJ4foKBjFko34Pxzw
m5jMI0xQhLzcswCJZ2P7CFFlY05Yyb5vREi7CFSc5l97P0FR+0ET+w8NRE5jbyv9Y0TyaTnNX6Ok
oTzNRKXO08bRMPoomBIwo0RF47OaTvDm6Ljwofp21ZJPYnaYXEGh3o6IQdOwjqc6Js/yw4t1E9Ca
P1tg+9DyHUOHmKtQNhGeF79ccdQd9e8EXmyEgysRDoSX7sBu+9HjpHYtKTutzv2IbAwNvz1wHn4s
MvGJgsB0hhFFX31ZOUwSlGA0eO1/8TKnZDinTycq31C6+B6xcbA5JF7OUBoIumX0QS1OtBKIDIii
FKtMyKD+eE61tNUFxRsemKsbwMo0DCXTt451fhYuWMQ+wLQN5SAoFkVnAdNf02pRO+iPztiZRnPS
SeEN6Er40h1bXBWti43aZf7afioG4xRBlTiAKL1JW0nc1WwQIWdZ6MgMQdS9o20O09d13u3E1Wqv
3O0mjeORRJLBKEg4AwRfNRy0ltAgwtClPG9uG7ExS6ekT9wJgvLyIQQ7liWhC1OyAgYdSKsAdDV0
edEidmpqfemwPl218WFugU41v/qu/A44q+4TZKpCIcEXjxcXjjN6eI3Wnv2QsHjyvTsRwsGhk7AX
q9AOH7BNOvSoKhKOeKJsQ77BUNztcOJ0uq1zytXS3p3M493BH4h5Rmo4Xpj27f221QfKly2768P9
axuCKmSxTXXoI66fQ/fpxG/ejuuPvHQZYscf2sXzDhlWYahCf4gExSMGyNlXruUq69CWbfE+QzIM
xHDFLX5ojTMKl/L9XuiUK1i+7O472Fv8iGRUpiNUlmiw0R1I5zNrDgxQDNgBS5f6Kufr7+9nsXw3
Eo+5p++ZMIGOMd6kjQsVrMd4V2I7WCG+vAh6qFs9HLH4jAgVCvxCzlycAdrrIR8AsFxEKJz37SkG
gXhOj+vBbCrFjymrllLEkda/Unpq04MadjgnuAZ6qDOkwzq6GVnWYeHpWbhPfL7zcXpal8b0RNZI
Yt4iQGqaHvkUAsrSQFvLA6oYcs4DMA6Nbnd/hWYvN23vr00bemIxmWVdFK7FLQjGwasowIO0pNDj
c5dLmBydYbsQs9RqMI+LfXMyYbtBthZaDQbg8SzQxp5LTzqrQZtjPvJ0+rDH4QcGlC+C2Amo+okd
n5rKMerLPfNo/yylLF+gItFZocPrA15P6z4sldZp7E4tNe/nbAfV594o3c4jBBpLoOg3oIQCEFoB
tQg7JIpfet5GYO8VDT1PzpCbdP01KNj6vvz3YgGl3mA120yES+RpfPdwF0HG6dj43vGE+6Bmo8Sc
MyGW6eUJ0NKxO5DzgOYefxdEk+esypnsrBN2DHhV4BIoOBx0FwzX2XQ8Kd+JE7TpdUMpkVh1RLn5
4tvW8pHiYF1Yg3L0eDOGV9OqLCoIWnIIs6rUlv6iB1Prb7o9tN03WUcmvoasqBe8e3jI20tMwdjG
kh/Tpjcp+Te9e1ROd1vkCY1fh3OaH7I2qv4dSfzTSCNJpjtipsmLTNl4NQMtg4HAvwNdy6A0bazk
3qscPQFChYLuDALMjgSAb0XqfPDXoSI9RvKnt8dgZ8dEFZ47tBfujFqID/SUwvtv9ZM5OZXIsI0a
ZJhax4pMYAtBdwi6GsRGdI0k0F/6KRSdYC6Otvdjpte1GrBBbky+s273BXB08caufnx8pysb6EBu
SQaC5Afjmo4dDKJhw2WYKFhR8749E9bvTFOKwEJzgU6ss/TLxNMRRYUB8ENO6LXmD4eli9EirUqB
Ok/QXh1YcC3xf1K+rA1ek6+iZg5VCPgbCpo/HoT2mYjp6NHnioXBLFyDGx1+fl8KzXZJPAfMvFBv
HwF8um+eZpGmEzNJPKm9JiDEzndLEIEMwej5eQEeY+zHvfUI+HeosDQ7t0f0/ikUEzWbv6KGply+
jWXcgf1ifLPkZJM+YsahP9Cxu2rJiVEuvhTB/PYn/PAGaKTU+UrpnzGguJezCnw3ps/U/LRUAuW/
crdIU3MVtAw2R2vmi776ingD9MqW74MZWQUZiIhuP0uS4p2DmTHQACFku8jPHR3EyEIJMz8dG14k
1q/4PYbay5O6KGMJ5wB/XfPh0bjQh/fnR4DRXWiLpt2Bfjz6ym2xaQwIIdVhi1+5eATXmSyv/S0i
uvRQ9VRkKeoajVACOkyOcm+X7r4hv/VL9W485rWX/VbpYjPOIj67peG6cPxdmbm25jAnlZbTcs3V
GQkt81YXDg8JFZPcIyPtIH87G8P7PSgQxjxfweMUQvyDB87jqs4U6BEg7kRAuNlBBjx3QlsT9qPe
3EEtEbumFc2u4Rm+PXYsIfCJtyGajCEuhJcrEdA5sqzFaZad8pyTth8XRxcnZ9JNUNwFZJX5O6Q8
uvIokYdTIgjgQQSC70q1fVadrrOY4eRoJaqJz9JYmulj8E0ZH7I2njtk5S7oFe6WM0fEtSQf3CKw
Cpy9CLZZdKwybq8NGD/4ySFs+oNXFeMEhniBzDJPO1gBv2V0nGdPpt2qjqJ24icCR4y7NbDMs8vA
4VpnIfP1KpcN9NypvGso+k0TuniXCgLK2QNbEUYsEH3tQpUMZULz3Rc/0DYMi1y5dYKf9URY5HzW
EQFOWtWd2Zo3SYbEkrjyTF+Neidtb6dvBo7xLoXoM/+sz9KcKHE73LdW7SNC0eV3Z2Tl4LNOO9gP
0XqQtp4txhsDWw9weWtRnTq9nAnD7kcWboQO0T+5iHlXZnf2PEDh8GHGEyYw+R6Xx8JYi1Tjk00Z
yICmqr5LHl8Yc9tliIufag1muYpvWHMeNxAEVc/mMW6g/uTpOiAoEviHLbk32xmkuRWSzncEQmic
/Si4lWAto3tmC7ElWZwI14C6K6FSnlINwnU2szb6G26Gin5ggpI3NIQRG6b/8Zl7BrNi26TVn7Y0
bl9ym7JhO4YmioT/jHkzMSndgRdr9giTdYzePCYdYXNf/23z9p4EpW6xH8WsPtRzBraS2ghDWYll
xk3pJ1HzCfxGCdtMVgsIl9DU7+/0yuxa9Teg6rGuP98K7DYRbtQwvmUUsPIaFOb4RQVE+DlHcKQp
evbbd17Zzc/ZeCTi7zeSJfvqQZY8LCYSKoxpa2rJykc2kzit0bjT8Xb4+E1leO4ZMzXw/5g8VG5F
nGgDTIP95x+NgtTCnG82Q7hqRcvj9zQf7R20V2zaTs/I0V02Vu8qDGxKzrD5HQHgyKXFY0CqMswr
PDmkfpRGBMvJ2RmO50q/yhgSwHlE43zrClCrA+0haQYQe3O1yoFP6E1AAyMNRRv2fGwJ7fzRCT3J
5h8p7QHxiLEMnNh5hMEayVE2j95seBWvc7fsOfjAiWut5SpBLEgB3Ay1ZmOvDv1JFKb7TY6rPGUA
jUYGB+Dbcw98r9UsclbOdZi6Bf350zOQqXepA4PSF4dgBAhngLZ1pvntr2JWnRzm4KsT/MuKZF+3
DQUMxtAJHWu1y7qZ+u6cIgY1+LmIGqe2bZtfkiBD+HlwrXgHcbs+uzIa5CniWavLOkgzLnhAHsz+
cWOe1fPYDYR3UUDnLvmCWiv0DzLvZZx4QpUSjHsdaLihiRvZrOeloAnOHijTb/b71+UxoklsZv9/
3HJCjyoLw8LDHREChod2z+wnZohAMNRB5POAXWNKIfT+cLEJou/yuzPs6RmaTzFjGe6aue5xEyv3
DHZc2bICP+KeZq6hIOj7fcH66lR4lCOkAyXWok/OhFLz2O2uUVIAtd/5WV0Av/jQYowGY0hG4V4M
Lw2pEFXflxxce25/PuUYx+hleuDkhuQr4TqOmQjderkaktZfBKmx67tbAoSLTxS/Ch4R2SKB7tGr
GLciCP5lgXEI68uLe7yxYPqDk0Ox8EpjsYGWJWyzpPhj3wlGDaf0TxoqvgHHNmCH1ue10qnRRelG
3kPw12SJj6QJzKMpbBGSMJ6Aw7c9ljtZpJgPVVd1xVcgNQ5iFBdS09YwjsqOPZdZzTpqnZA1J+Vf
APiHypF51RkDHzuLboTwjcU6iapBH4b4aAE9f+v0F6yzA7ioNNQybgHqs4DDNgtOaL/VWFKm83qg
0/EKuVDZ4SGGhAxXxTCoNRMP2DrgF+Kd73ciDrlvHEl2hpTzjiS8XE14BCE5ekMxythEpi6ZRLlV
qg6DTIHaMtWkdee6EuMR5IkW+Mq7rzzCkYGJLJ7jKKpZVTcFu2fhE+UH+OETWRKU10fa4mzIlTsy
gBu1/XT6cl2rw4l48DxY6nylvH76q3UA+edim3iYoN5xIn7CgUPJm+aHyLMFCCtvvRzV58cfLhCB
PGcJFvKXXWIvw2ODVQxVbjJXRHE352dJf0fsHfgmvpHENq6UGLWo2nsimyONs68gpYsuVPHtk4aY
GRgYyQhfFwSqogyFf/KTtejytz/uDBn7s8Q21/fy9M91h1F3jK049ClzCix/H7zTgN8TqGK02Hdc
sOaBW/pkmj0ibYK6oDCJJqXrUYV63p6jlzbyccfLSsx06Bp74pOzVFrgz2NWDUiCFuj2G7fyi++f
NLaKFhxwSAJkWe8CJMo6+2ilTBbuOVQEPf2CmWmPbUSODTKkuoETkafDMWPwppu+qPtjtja1mD27
U+UrttCUY6LQFKzjdBul3xF2YgzS/DHydVcCFA5BWyLI1BocozT0YLuzeJ7sUPrT8vlLaFHE4odl
quDaH7M/kg1FFS5XiHd05gvHxrybPz5rza2Lw4MutGl3r43mCWdwVnW/uzEfEMPFXpsSy6za9Sx+
G32ZB9v3MoQ5wIa44EJYyD00QYwuMBpRDKT+j9R1FEH7jHYARB8Jiyu2a48iwA+NZAyq0zJFlvml
1Db+9ccqLalZuv4wYm2GpDpbAjnW4SO4wsxLUuASpSYglxeShYThC4J8CTh50HTZH5pgwDpZfv82
xu8pp/vRO3p71W4AznQ7Af39NHlgQG+2dTJs2jrLcr54/PwLUn690TtItxXYiqXaFQwnM/S5c+At
HPq+9kUF7Qp8l4xXRXD30+DhJ1jiN/9hKFf2KYqvyD7o4F3wupcEnbcebTr4yCnmCa+xmulrpLDM
+3QvYuSrM/7YlemCMVQZcuULn+z/5T2WhHjK08o1sJlnGaMncqbwH/w/0N+f8V1Qmohmu0b9zsAQ
r/m66p1QKb6CEOr1tXKsTrZTb9cJ4/o8xl/J4ZcMnpMwtgK9VvAIjrw9ob+si4cFzLiNaLUEF4Zf
xpKV2Je8y5WGll0y/1cEfHHNStqGtFSy2N4VrYHYr1f2tvcsr4v/cRHwqW+nYNSaRp/Lx+rF1dOs
S5TE5zh+Fri/4fHm+5WJ8aj0cge2/uK8CDviaj/QOfAnI9KPBbT4XTOCb2fKTk+gExEHVj2Iscry
/9Y6utCdKa+Ry2elB3ahQwoFeOZCR726taJZ9BgBuzFXjLs2J7Rzi+vXOQW9FaANVWBM9O3NwH2V
a3TrECDTV/hCiJjy6Pvi8OEy2GwaQEtFxurg3Ui+CC1lm+dhCyWbNZzpdXLE83GjG6QcdEeVzwiO
q3podzIwtOSMoRJsgo/wwTva3aNEKjLkasEXMBus2m2c+I7/TLYa/iJ+OFwjWmgikuRoS7ZBSHYI
FGP9GyOpg2OAkSs89LTRdK7lli9OrnlWvlajaSZq+unBhdH/465/HXPbNldVgtSWJSJn5nGidOeC
aN/CnVGVfcW9xnQWPjH1rAj7FPrlvCIVhWit/XnS9+nv5eF4y07hW5HMUqAzT+MF0LAo+R2oRKAt
KhPp01BP2zl43OjKHbjYO6dg+T3I2IJDBSJA8tRhkDUKPm/72IroN6/p7PufJT0Mc/STyvxjlc4v
v4dpi+5iCDnnfC9amKjiqfqzAeS99c2v4vbkxgZVS/qmghq9sui4t5ARWMT1uM8VfTiQUQGozI8R
onC3NO4phl6VQK1cCwb/3alB70c5FF9Xt5E8NaXR7NWlNJaApagJoukuwjyyPDXK3x8NcVm2L+I2
7UWaaLDnJoiDcPdtjRAdZ4PtOnQkXqTPzyt71QUUnSX0c9JlK9W79b82HYNj9hCBIkGsZvLNSOfl
DWgux22vW0au0+LFMPaHPaZuYV4kR1we2sNyJ3fW5kRddXnr8rQCJ8poddbFpj6TSXK3nuN5oUDf
CjEiXLVSB7LsBjOL/ycpyvC1g1I505FUy9QYqqGwjGvAkEFmbWcqbxJSFCBnHjsnJkgFSYqBW5+r
puBf/EMIJPjitqDVDO76VluSYH7hAY2VjTgJFN2qsK5MzhuwbAMrZq+N9thz2dlBHNd4+sZUlwXH
gfAzIKWOe0wEmGlA6S7JsQJ8ydnVrMiCLFkIzeabqPBVs4I70WSicGpTzYJexBxZxico5eaweRty
mdIeTeE7XWWxGOtFwjltd81QRFrF6cPeEP17izNpRWGWMY6FdUmN8np+A4jwLmuNMvcDSFbrrEoI
81v+BzFGd3fYD98iujUnvSjBUIJyfqhiZv44ntu8nKC+Y8tajcjuLLpDTJqMu0Nrs4leuZTp0ywf
SpAtAI8KiFurpBEknP7h35pMNc+pXkXJtswsk01VTGVhRtbHHTLA86Bx/5jZ7S/Yd67gyan8L6J5
1z3sqOclfNZ3JAjp2pjxGULkYoEKmKWXpcFDmDARHX0rECckkLWVGJvQXXTvkA7c0aH00B+FKVW3
Xugzr81XvwWzLpv75haW8coZnDhFtY4iucFS1cxuNzbltNFKK+86DKW6S3W0CkxsriWi5QJkNd2N
vxStRUnf7yCnciR4Wt/FUF/Mc7LKCtKVyCDau3h7n92AKYFDffFW9dtKB/WuxNwuNeUk7HSPxtNa
ZwcVkiXYmseIr/kH/zdhn8+I6p/ndtcHJrnEnBSLQavZVL45MFsC++amuBajHPLdbmtmBGc002NB
i47KV5gV1n5LJc1kvf1WG+NH4C9aWFm9Dav8ZHOPs1uIoOjltLtqFj1mme78WOhl4j2zqrIt/g8T
QO3UwZA1z2E2QvR9xHUcO6T1aXA/KjAWc6URtp1YEnEazUuU8i9sb1w/YtIIy3PKPevT0aMOtn2F
xMhj6c7AIuTL+q43O4JA2zDUHm0SY+b/kCRBJHM6JPe4tkucAKNavr9xLEgOsb6kjNje40p6pEl4
/m1OujqglfcLZuaF9kKI64LwcyxcNniyERvYL8FmTuPF7QNjYEs6rg1EeRMH/cMhNUXq5lZ0LFug
Clge5Wf1+7cG3xSwulDyXS0MAatZuq7VqKrEw0yhFDifvE9rWa4unMo2uL8Mu/TrBoShwBLXePyl
5k8IMMTp0OPDIEbeUipVYZhzMxSmEHE7tDdMdYsm12roYw+VjYNVVHBgO3/rkf5ojNwrS3P2MntC
LVzYIViLXhTw2VAE3DpTTod1qhS5dpLXG620tIVje//vk5kpOWMC89qxAlZswDUL++TuucqT5mNw
hLvxy/zcJXjuo1FxJbx+KUW6TnJ/so2PbzXUKnwrjSCWW0uDuxkeAd9KQw/ShRd8L9v1Yz1ny6cX
pGqrI6zNnILIMR2842jeh25IAOgEHAzOf2stznZftIeUOD3+vmiuOlQFsoBST6rVYepLafSjxNp+
iEz42FYTdRenBRZqbtMNIEbjP/BposzEPTiKc4LNM6IEw8zU0d+3o9zEKOs1qYCkJ3y2xh0/txiO
g86bVa0XhWcIuQCgqkzd5+VgNYLvORHJQx77qKoPt5Cy6JONMGja5j1b2eGSpteTXSI/MIpNk7wA
BocH1jBDf1ZOVhopFO6ZsY2nNHL3MEunN0KIyTM0jfvH+8HYv8bwdkEtWK6z3+drf6vhKb26fkOr
tzDsbDi1J+L/1d/zP4f2R/rMQgLu73t11aWT32GAJJOjjvp5xTSrfctkRa0RZv3SpJ5xm+khXhM6
C/NWNgM+NUeCBhugArP3IhysTE6qLdQ5SCi9R3oK8IOm8Au4c5aIx9oRhud5Jf37HQKRjH/+qk49
41QZDhSSvIK/GFZuseymS8Xf5Q84+CZtYoCtYzL9/2OIiyJlRMz8r43Xl2/nNkvMJDLlAuD6P9XS
/NAnjs/CErTisduJra5wjwpW8G4O1sdOVk2FPBQgR/XMZrg0BMiNhSIaP95VmI//nIByqh/JLMRE
aL6F02nmT9XVwuL50R+dYJ/jrCP/ub9yf/Q8Tw9z2Rs3y/+itowsnXNRtmQrq/hVvbiLtXzdUeJM
h16lB+H8V7QjdvYipfZ0RGj4j+Dzaf2c4NjFPQGVAaF43yKpJ6GhVxRfZWIf129S8c7zEz8gYwcw
Y1609TSntxJphiVbeizWqfyp+AtrWXlDHPJZ3tLzq5lLnLePjutGjYxsy67bDE/hEciLdbYgXgiR
fW6SJMN7IyMaTMiaxbIaEvWwijznTc5RTdJW0v87lGRStipIsBQcCxck7bdMz6J65Io0txTrfjeL
j+meTgvLt/bvUVoNTRuWe/oymaPysVqoqPGDxee8MRfv/ew152zzY8Y5BD4UGmdIpN2hghQ9Kd5G
kOr5JoGf1IW5AjyiqsYGeBD4jVazCCyo4QhUMC0w1iaEPF3uxhfNkAMUCbhwfI+adf8MgCZWZlx2
hYWZK/UURMbtTLRNpKio1ZJSJfkCrLHu2Z5XH2u0Bn8dbYFBRW26dcAIfU20dP1EJmhEfhMx9kCa
Lsc/a8iHHMywtY/7g/fvUWEl8HNdOOLPyur27gOHb2eqeY2ObwB7TxUrFqMwOD5NLG3fSa1Hxq7L
ybR+wxrXOfJRy7itwST8T01OJpBrTSJuiglOUY/afOpT56SSrS/K65Z+93m3+UDxoMoAYgEMUjfe
dOnu3H2jnAvmdgUEVY9Wt156kAti5AIBoR1mnA1CYvpb+oJVucW4f+RWg2lZJZKcVx+vtE5FrSPd
GD/hgw/A7OCsNh/pVZZSCMaU2EoeOtAVQqBGZQeCiwo2X9yRTpdRsp1GZ7cbES0F7d3FFQoEB40l
jErDy+TxlZX+zHqFt6YY+U1GnQMi04UTIcdfDqYStZ8ONeXdGSH/GzijMX8ubkgFKjXV+h6Z1kKy
n49BzeN9ATbVHLvysKyf+YpRnhtZ7yFPEd3hDje+8C8/FvU8LH20ugE4Kdf3VwrqaT+hkQndgY0P
21kfV8/9j3SOlsAGFngNaPquUPeCdL0Ezj1/bROwSflY0BvePtgPxGI86BxHiiJ9YlyPP/s6oQLQ
ET3cMc/zODMJimX4OK8UcwuXEfN3MHqTbHNyGWVauo8JTes/8Es27DeI5OGdminpTZtj+5nbFnKs
grCqcp9/VuYvkQ6hLG5sRQnl30I3JgNG9Bf25ggcyKzdYx7JJtcEUJYriTxhED2uziMKC/xY+2CN
6x236AKOSlQ1itW9zvDnyLG+IRSU7dT2V1Locp+AbQ1654fLFSJsXB0A14E4RIS7gwDjTEa0+MkJ
8aBtf9+iLZl+KNnyzHrtglLUtimgKfTTOjD9tVRNlKH9/eJAJ+94VwZarC9RNcKVymk8+Tnr61tV
TraCH2n9Gv03ipysymGgUuIIBJz3dbbkuErL+qc3SAWMTz5HSUJfJEMBz5JJWWBrYkKKM5paVrEm
SNsSD+TOP/TdGyzDVDlj7nQNqLJvgjV+T6QTWDlAJRZuvJqjyzYwrW/u3dsozcHkXPpDaV93Ipz3
rC78p1hidDP5HeH60Z6Blk67AMh3Hqe5BeIWN0c1l0qYyJLiElOVfE7IoMYt4nHTZ0kV7jcWXT6d
uMrgUIajS02/ninHeWjfTXOhoubE09nFshNCi4+SE+yOc4hpvsQpKCdQO9X7hZcdR4YSWzv1N2ek
4UDA2J47Q3h5HPJBMqV6ZQL3YGB92nR8b6tNRrwemXKp/bzSXko4oxL5dmrE5jmD2NEeTCsKTRDg
1C2fI7tqoR9NHzsNKk8z3forbfb7D5YHmuxkhRjHbd6pFnw2Z4E+UFkkUQgX7qumXVr9oZFhQ0w8
tW5/z1wQCKY00dphj/tbRVu6Ic6IHMJeT1kMCfh5f5XAfXzqnAJE9BtUAO0K2DYg//sBgF3RpaZj
7A7b6xz92QMgGGrl3fnPZb+GSHzmO0WSvAjoHA/L4hmDeOos0gEPF2UAHxYn5hlYKhE3OFL2KNia
usXeAk91DbjExzFHYiXWowlYnKIt1vZkSVaiNmh5U3EXQtzM0l+YhMkzzF5L0TV76w9f6Ow3BmNL
UNX0PiZndcN/VhS4Jem007wx7SWV1sZUHqjvNRWlC4MXIcnePt5sXnA2Qa7SOz+4gMQSpQ2npIgB
5jUgTNy/Ocdg6zzIURgiGffsTo9ZnvyqegokzaH0/K7rzhgmHBlglydWgCmcM3loR0XMdOcN56WU
5NdC8+CijOZdIoMK3E1RbkVCb6pYGUVzVwHUmHcn27Yrs4X714Yz/5P4E3ltnMr3UGqrIzdHZKXL
DetQIvD+Q/jFbz+Q6tEAvMMao1MwVU1JM6QnxG1M0Kku7SISztZmU8YsE02ZoKN9IPAowewSnZjM
xl07McDVzHHAcy3ls/POiAG8WMQNn/kTPjQN19Mo6GxGMNfWeMlXAdAD/U+dGJtqVIEjZRYqhSGD
AGoEVrIw8Qxrwh5KOWbvyERZoA5rLAnqI8NHi6gOu3JnE8hipzRbPkaUDaEFlZEKO1FfoiDummid
/A8xTd3w0VcZJfPFOXVDqCdJbi5n21SpaVJRJ0OpDYxHGukalPZSnVzNAHQag1jQLFhacGvsBuId
NTmZksLOBbc9XgxU52keoxt//CYcHNkn7TK+2zFUbWxkedIhZGk9RdviKWjULtZAPKPdD/RTvvse
VcMi1U2assshSZVeffOaeU0Pqekw5aqmnl9pwtYGBXdZhMsMnYjekHPa8YDGXcKAWutbSkZDFzvW
nKMCQLPLT/wJT3vQdeV1bBWz+PeHKgw9c8rrPyO6zH3heMvHIgecVgSgIuE7qqhiBCH+OJxxMu4S
hu3t5a/sO55Qy35os5r3Jo0ocQWY37xYNdtFI7Ea0hEcHNRDqG3l/AyN5L4zJCJV9jAtDL7LXP45
DRqQgchSkchfLT4xb57bXGxVU8VuKjEKx3QzJM1eyK453Elz5hzxKpV/TFcP8IcZjUATNi4px6A0
2D9VScwUhEffsN8u0gnV4+w4nIuAPag+SeHIA/3MQBrdlQjiHF63/ngk8ui14EmWhza9ys5jOss0
QM+K12llfda3hje+pMaM/C/WqA7Gs2FCVXGknZ1Wx+YcmbNXQ3qUvKXvCZ4gEN2VGiqfzWMuAKps
LuPIIytttSae+Blzw2qN9cIVXCCzCO+yvp2qagRZveitcttAFlPwp0MMoVBzigVM0sXadTUKzwb1
fV2iXMX5mdgDMBefnc0aHmzilejqyG2uI5MKtfaAfoi2WXlQUaKwBjIn4FqSTYmVVDesBCiDsyY0
7bQYjeMeLaxmQZfojMGTIlrGrRtYTn/srdbYf5+PReJTP9XmMr8QV+yF0t4uSCQdFA/B+ibSZVxd
uXLLMJVktqQeL6Qz4tsTNfFMCBRba+hLLJF1E8ASIzkLSGwfIIkrvASfudM0p2VL9zLUuBnO49OK
Wc/WfJn4YTuT3sgXqgWuSKSdz8d5ofh3phJRmVuuCTo5D2t1QgSfEFybQwRJ3ShDqAciuq65x7Ny
Z8YjF16VvwqhU3ArUeAG2SmZlYdV0pOyrUQcGB4kPaKJCEOxXiOkL0MeIEDSEHhTCa1jxN1qKG4p
gpvDQbHYLqceHgDW5IGtLtFQld+RrM8NfEKVH+p/HDQ8tVU55ux0qrlo1UZTmHl5Jeo9TQPzUYws
OL0HfI5q2dlRxqsCs8CWtQh8CwnGc3Rl80jABZdllgEhb9i7Ql2GzyNtFSm+xA8YeoP4/o7WfPZ/
1iGiKAovjJ7cBddZHBcwSKVRfHJ+ZYBHHkbyAoUNg9d1tqxrv2Fm5Uvt1XLzr1Z59Ber3cledKml
lAAsX860ViQDWO384zaB8bcrNCDDrLdUi4DGRPoO1VYjHiZ/hRLfaIZpbm5UTpwgPVLMddidFB2r
MGdSvwXQR8SfyXg3vhPPbLhj4XG7f7swWfx5gGCK9TZxqREntdReGaeK9Kq4iOpgQn0ScXF9xQzO
gjoM/08N3yDFQl43D7lJ0OT0c/sz1S0wa2eRevfrdw0CxQq+t5n5Jy53z/sh5unFOFvjIOeMvGE2
qcujlCCKiFqvF71x7S5CLS6YCmTaPXjWM1nfegJQB/A5zjfXxLog31FKp06YxIuAdt0fJiccYBXB
dIGM2lgj/AfW5neYcUqRMu7oYAty9SAjJJvEF99uH27X9BTX0fNZfZeGJkjmef8fkXj+l7IVkyc5
q/Rmm70Z0PJr+7/RNohmGV18KnknvDSl4l+51W95glT3KD/4w8SwgrMXUBm+4YBtyCq3RCb9NdNU
qu4S3wcbX6/D1yw5wzeXfiEaXF6JsqrtAFINaPW5WkrFAZcgZYjUw4wredmZPYGK1FkgL6yQx+l6
bdwd3Y+X0Q9PN1ooaNWYWwxVw5ceSyywXriXiO44UFG5jCJzTgF+asP4+WOuf/xR1Pjw779g6QTi
/sk9klxr6ZT58VfXJFKrRzuheIqRN2N7mrqbpFt7WqinAQ5nZTkRdghlezB5uBmOkWObCwOioPaD
wzNsFGay79lkAMrCDmsGFP/Ch/Y6C6IKsSvkYb03lqo/Pk8OWvt60C5Wq1T7aLMbRLpGem2GGYCB
hUOK/N5IYNhbfmAkLVap4aEug+uDyv1Z+yM2xJY+c48pfLmkoAs37hcDVQBiiZtJN/MlLl+PFpZT
VYR+5Wtj/VlgchAqj66bkve6+jcrrP4FNcihPK3SKQOLCLRLItE4qoW+ciMKNKmjFys+1OPRQM3c
U4h+D9Sm9weyLMFQDEWvnHqA9LkJ367LO7S6OzHI0nsaseqSbG0T8g7IPHsJn7Jd+YqxmcJddwhj
skW9bBGqh7NuCkeOXUQywNZvfbXU+9BW9P8OvM3A//jcROsA+HUMJ90usANzGErPNOhFiNmEJvFM
zvCJ4KDcV2QWIZ2pwQenFQRZhvWnFEw1vP7+begyTlU9hd8hkppe06bceL4iKVhPSDURoeOerZ/H
1pC1StIufKbQ++I6bPdPTqImY+OFo80F7AHGZwHZTNeChnThyJyBA3oE3bKvhvJ5NqK39XHcjWOP
aImsAvD44lHU5yd8K+IvKRcYK6m+5Upa11+3wGWBIM6X4rdFJTYO1bm4zpeq6S/33sefltwt6sUo
qVj1i2W90KQNL7y/g6NaaOT5D9XZnToc7FVtUEgJjsjEG8sTXk7Kre67pPiMO64okPIF/SaNsdm4
icmxEloN8uWp9lsjBLa5v0C/ay0F6oYwJGSoJChww5XzioLCzmBJz2E+Onc4/R4TOg73s+0KB9yl
yuHfmnToLOBMLDWbFyBSIXrknVKaEjBE/XW18THsx7SKRxdH4J4pqQwvQ34K/9/BtzFeeS4otWqD
lFnNiTtFq2h4WHUmAg2syEh/BFKcN3ZlHLUHyDqf/MTN2BJUJoqHMTvQeQk0MCp43eLQ6Ou9Bual
lv+QfBkhqFDrfhoWpht6O1LY7hihOuziKugfDyn/RWN+Z9wM2CVgYQ4KGRAIp48j6h/xzh59LgEj
EvdHbvIoX9yDlgFZEKLrqUj/CEchZhvkab0d1Ou/UXcpWZXlcmfU2l0lInjoF+k/tSWiYLIk0yJz
CaTsSC2094Z78JXIs2+beO9tKEQ40ejqytD0NfcIh+dmXkwPs+VrcDikCVtxUUQ8UztMoK8Ux8Kb
ZwA7O7Fl5S4f9B2JlGp8V9NbKAN4iBxpbqwNNzX2J83HBVAj311eYvxvK3+tVcA7Ox5QrimJleyO
nP9B+xHd2aWf33d7G/E4UMkea6dUh+n2DH/0Hjq2yFawT/iZ0QulABP/SvDXOnzj40xH/8XgGejD
ztImSiczMNl6n6hfF1d5wH5Axx6RJSe6llfSL696BRRxGIevaRLM2eWsjdHpCom6SHEq9XfS5M6+
VLGHb/kBSXZgFAjeT0kSd1jUoSnM34+o5zSbh2SJZU8KjAJTSOxpk6ym9u27pjhR6wRjW50IZ1uP
xLPiX8ihuEdwQMaOzs5ddFT7j9h+UZnrjXUbKrQ6WOe9A1Ade9o8HqvqtlLUoGD/gCynfhGDE0gB
DqyCPMggOfXtKp7r7xGxNChPIR0R3p01eB2xekNwK2YtAGGHYCHXUo4t06FW6/kvFff1EIue+ZZr
qH1mr7wsCJC3D7GLrg0YY96zRMqyzwwuMpwmY/JTgHzpllqJ/7mg+OoMkgPfBEnsAjshXj+0cvSL
jnplEXJ+JmNfOiXtgvqPDc/3E4ydBMXZ1a7XhWAxKTu1nSgIXCEIoeXgcv0d24a5W12jN395rVmD
KtdG7UEM++eNm41wI61OG/EfrgLXXJNYvVsm2EW0nJL9XAWzBk6advZJtT2AYfkh/KYagrIVrH+D
XR86lfIavxZ/u+Bkmb1r2XXtg21Hw9LVQdFK/cawDZoIBG13akjFMTirL1klJygsBqo7DAIIenJ4
JZy9z6e6p20qMVetD0xYqwKHoU+4kWjvoY+a3R7KvFFh+wSmnNepDYa4GdI3BLHdrPp4TaUh2vwc
Gpc9w8kLLwDSHNdlJR7h7v5/8KObmLg0W2wA6222FoFpJHfNIsXQ1zJUYCevyhb73PWLN2ESPhhk
prHXx7juX6+EPGHzCZvG6TPDJxbLen5/DBACdwZ7qEjq1WrGOUvye2qC6/664/IUp6C/vrTG9dRm
TyKXnOV+0hExgcTcMRta8kIa4XXAHzVDtoOiLskKp6zphIbct4gvtn4QjexmsQXG7aSVP52pvmx0
ECN/2G3alMjGVPAOH88SZRc1sMEIS6rikIO/L8aMAOBGPhsj/LUD7sEWLJmy2eCFGC9Dg4a/1TgE
oCkBkQhMZr5BlS5C9R1yoe59j0fOACN8pHBx7A5klVd1rUwy5WR/L/Z/bm+tQybU+lVC69QSex/S
WmtfxsH+X6HaMQ9mAA6mG7iA/ilyKKq9lrpELW7bAmEFahQ2ylUryFS/pDh9Ym6fXvLz7gy3sTkc
LtHtPTvNQbwo6EtBXK+JEL0t2GqUJdPfKhZpA59354ZQ8ag1Xhiqh4vcgtaBIlI/OhA2crGHYI0q
t7KNli0VLwj2QGIgTKqILqcX5NgOmotuqfmQcIxRBiKQvknIDSVva2hwTnf1gwtqCL4qTynFS6I6
EHzUfsrQ6yFze00nsMehbPUqtd82IKTLjZLh0UZH5H7oJ9iFKJYqQBRCzWkwJgL6RnaxIm00/gCy
QU4T0e1KYHurKQqbJa/KpnDSYrPgCnU3zq8ZXF3vL9TI3gukkVDXLUU5gXFhmR9jDM4KrA68w8wn
KZAIPwpTQiazibsBAdi/ZWWZYKbe5hDjF/AKHRFHK6CJzEQxSOyMgOnmkdYiV76HQy7SVKHCGvDR
pXJtrvTLoRv4wGBbdFdR4KZbQtLVWUzRPKrtpBRRLbFBthXFNLoAsFLkEGWt3L51Xhv+hJD6ShaD
pEu8GoqVSq0RCAEYL5TrrWbJ2Jlgtw3MF3kyYEtIl3npFtn4pbk0ylzdk3LXZN03bJ4rGnO3Wdzq
/R/EtFvBpniUXNNWLAdhnlV1KVBybqG6fR1Nb98DGDF00Dfz8oOP+Ih7sRLEX/xKu/7J0N7xQWBV
CmDMIdhLNK9AKjb85KZ1vUAsaBQZAlz9Jx8EMPsbggW1TtMquCAo0rfTYCxP0LNrB2btRE3vYJbC
dQDshpTbZQ24S4Sqhwo97JdDlmX4DwVjf/xw8hdaPxhuQZBy+r6OGRTZg/39RVOGB8x2Yap+tx4N
0Tw22r1SxkI4GCMmhT/XUm8z3R6bO6Vi5P6Hg31vh77MAusbuUTSQ4CNPgzhLctxmZxAvTSgpwcy
NGhIoNPWWQQ9HLTPAoq5f/w84g413QDDYPZKse4CPqha7o8BaewYbglq8iaGZbSE7HWtGbbvz2OI
G7BtT5FxZtI+nCm6oGz+zSGxDHomynq/L3X1Lt8GkW1w84h3rU7TMA4Dlhv6dMC8sYhfiZGfx+o1
7lkFk7RdvJCx7u3XjwaJGFseHmlG04nmcROtBzpGEPlQmG2hQYIMz2bXhlm+h96yX8kMvIki1oC8
TBHLR6A4XxutlYCc8BWSEDFNoLEzzaoDbM2JuGFRsVehYzuHXeLfhTPuNOdsPS+udgHk9G6c5IWV
+NtAR7DhsfW9FYOv5izCkWZcV+i1XfE35M0KslHnaoPTpaeXPhUOMMpfaZevnY2iHK/AJDkJUUDg
DVY8JkfYLC+JpRuQCyYCZB0fN67AEQ5HmCMuDHFZFGnhHQ4iKae05hjPOes729soElJXnn6Ptixc
/TNNQVcY0KTi3jQAsM31VvRl1KGyMthlPO3zc1TDg5nzz1tU1Qis0toxCMdKHYePu/NV3wDMMg7+
WMass+N9w/FfTHBBlrsEk+bGxtNvQzaBgjjbR8lOeCRMXP0NAMdhtRfh/Xl5giABnG4CXpZUrJHs
g1Z7lYdqed46lq7eP883xDZZvrNJGg7W2EFtWEMdSdOMBQZZCR7kdFibyt8Tth/8byXX4e2/RB6h
8rfeTJee1r7V1y2SGZ84YrK87zIe0lxqFLTmd6uAmHR1tg4ERqggdr6BQAzeDP3fx3TaYDmSwKqF
ggBMO8DK0zCgUOBqs4/hYj+rKaZhlpu0sbFwoLcO5P2dee0L2OnRymi+m7N66/z7Zk3PfqhyTkBa
OlaxOTu+0oXog3DvCKeVCVQSkCS6tn7IzAMkZEAcaBUp+szcRGggUq9yF8oCdRQA1n+3p+8O3rVg
BDh88Rfuw4fi8C2UeMzX8LKmE7iLYEAMyIRmCHBn3XFqr/KNL3ghY7+5QwShNVr6k4b5ZdinNntb
dxRrvjhMA/IhAsoSqp/JvEgpiEQKfvFJgF/0ooB/92WhuFTpe4GJebgoBxEITVfaa4iJalgQ2pT3
n27o5AGLNK89Ml9U6wLKvuimrALVsCZ06Bzi4OwNvwbVl8nUFGkxFbB34cbA9lC6zebBQvsMaKUv
Klhf9g/z4tmola38dbeUBrn8u/VTW9MbBfKt5olyGiN/9N6n+qcIwYRzHX/2374is86dLAAC4N75
wLt0kcM0JDjKfHaElDYfIJuyleGQ/1Xx4DEV1iV4uhyHDTmoA1RrELF9hocb75/bT62Ltp7YhEiA
N0ir8RZABbxO+Y77t6h0yTYbzCmNtOm6kNNYbtig6kqHAYsGmFc6liHNo8bPXzQeg0hNdo4GnVBM
iaUofyqXlEnYR+8+66Bpe6mob5+zuIKeBWYjqlDBOV2ZI/Vcn5RYNawDX6q0wPhL4cGY88ScO2K1
IIRuXXZS+JVkXD+uu17gJEyc/TOAS9+0j2o/GVui980LUpD1MQ6wQpoGbYx7dLEZDyMbWPDqSUtD
sCIMF05NdR36mWhtSieWFng6XmR3L5jBCPgEh79sQj/aXpOjEtjUz5aqp4RrIPfWk+xyqGUKRtOI
UYQoV90304wfDFh+gFZTqUBIJLPAXG9uauNVDirxqHCUlqsYP+6SHeQ14zWnD5RfqO6p7Dzw8b9D
OBaeEzexHxhPtNIc9YaN62CF8PCiTmdAkP1G8/oqyqUgIxG+q6RTyaD9BbmT4iOqASd6yp7z10wf
QzlGZYhUOHmFr32on7h09rRWdi6gw1NnsfLKTQ5W2FbVHVj5z7oyIceiqZwToAEd9LUg7+vv7kp5
YhSsP3AzDpnXz7n3xy9f9Anz1Ce5JflRwf3ZwLuY41QWS9Pm+SNqf3Ji4OX3L8nIBvvW335oSf/E
+Hpki8QPgluOTtSmSjUzpKw97pGtWfHye1Ye4BPHr0UsozVdzak1CoEUMocSES3qQBeSwHxfUdGw
UJQLBrcHFETCLXFrKKJF5gQqF3VV54Cp4tuzoxnBPhvhCRSKxSdald/AiLN9riK1TLUn8DDwt+se
u5iB6ujzC1IqT0OWPlPnA0K51QhLd+X72ncmC0VPg2WYVdg8cNc126fcFzeLFO/W1VaG+GvdPZUe
NwHf0GJ/SikVYOYjr/OysbXYLvxDcmfL2eSjKfJNbd2IM6wnBTEUvhYSsiT0OB0nV+x8wSeCDaBW
B1rSNW9fRf2HM7fuKn6d/IsxsEAGVuOguAKEuwEfL3Ix2CaG3PmycuET32WKsNOEQmUJnL4nQo/q
QOEHjeGhGsdCqXVvuM/DuWaYSWFv8oPxMONZ2ErUcxWWFu1y9rwjFTZHoKaAwBBjVIMJqKVlB0mE
1t1tXVXJH4HSUy+npNc+dCaWpTlKqaxaABS4vVsYZm9Txas1t6n/ds7ficWzXDxc43pZLjnZVCLL
6b4BR7LeRGB11BFfk2WE/MBOzEIbRRkWu9IkqfYMdS06PvzLr+zO6bz9vb9fps/7uRP3puoOy27k
GTl7KpvW2swLQ/RSWYMVcnMX3kwpQ3xo2m5d9bbgC+/N3vmagT/yWFuMJ1H7/s7W+ihN3B+LDenS
wN+ban4p2U+tlSOItH1X9ceyJOsJ6CM1VLEvzRWecnYVjbAtA21cnhBzFw5Pr1zBRGMnq5CJ2V76
yUoMraXuKgbNwJADHDBW8eZT28fqHQxq/lgbu87OwXrohLK98bfXjRZmhHESyJCOOEbi50DBAhOl
IRpplCYTEj624aoDY/odghCPJkiDUTvJOv6TF89z4yf0AJr9Eq6HJ4fhMTsj7+OHDwi1ZI6yJs37
eBgdcp2pu37I5zs9PakQQ4SCvAVxd0JpsmwCHBxQOA6reY67r/9H0JSgiiyi8HUHdl9Lo6nkrYIY
uNI8Y5wbL254Aq8LoqAnBTS1i22INRGg9IWBSiNoOaOMdKyeVhNRww9k6aL/senSBkikYU09Pze+
QzBwpDgndrLpEoHu982QTfDH8GlORau2KJtVtyfWlv5sBF95WAKjkBSK5rOLrWlv79pdTnsZZLME
us3Qlqd6/W/qV7Ad8CpmajIFQSQd78lFQ6ptVHdn7mrU1np2kCBAS1wPw+GfapqcwJSDyrlXcFf4
78ztlENwpv3n7Xsj9Da8MiBkTFNFfd+JDvxQ925dm2RtWUqdMSUwBUSXXauqKYp0PFtsUge04Ma1
MqXNx2fnQxlIkYMwgQtk7ZdOkW9VRrR+BZTvfVr+0wPUq/DrtbE5Sq2KvLKrbFGi/3E1nx5nkYji
2fyEHJm1e2ueaPPNi5WVLd/7m3pPw0H+ZzoESnCiJi1dR2ksAWwgYNXNyOZBVXcRiLsrqc0UtcDQ
83Su2TwNjsJ2srdjrRe7CM6BwSCoz4SdXf37Oi4f/XWm/J+m/8KepJziAhYNW9o+Vfs/oUARELBi
I6aaQ3MlSHRuER5S6PZhYeuFU5JdLGnt/MsGXAQYP7GvHWKAxKH/g2SoOSNbU3cVGnjkHhcsc3BC
sFG2/QDGfYGkLjOdgl4iFWvchcFjb0SmsRqPPzvGQR6gyJzDAkegoab4l9EZH6ONFvqcDVLjPYwu
+BDgHAXJlR46sEZmfuRfteNodSse28TQmIKnTCA94lwQJFeOQUyxwcdBlh9X1HLOf1AY/9YF71hY
T3bRXJ1MDTXuCMVzOqUQdPy9ueQJOt37L5bM4zSLhytbr7VcXNbnjEcaBmKa/syVhuLqDgf+tlhq
BhPleyUA8kgjp1r3iOrDWkUB2AvKTpz1xt/d0noHfMkkIL6DtDEpSYzGoy9U4e2Vf0JyAdjLzeR0
5nvJ2CDxL/t3ta2GYJlRqqrbvzWdt7w8UXibNcArBV8sHaSz/4EIdBPAbWGsv+NLl6BWjzYC56E0
eYW0JJ3Am3jQeJsDNDFLbIjVbKrXMNLbqSWVPdeo94qcEk/DDouBR9sMElIy1MrQvlX6qsG2Ck8g
5Q/OJPL2oXgXPC4uOsub/VcAflxLU1KYrPHiO5PmGmY1lnfeRZHABj48p0FTRsdawm2z+8VaqGxB
Ov9XNuaFoASxD5UyHlqLfpuRjRNwlanTHf7xX9GYBDwa8XsmFzi2QQJC/Hb7d0LKfZxkg18VrTrN
UcIZ7cyr+/NSbGghs2OuFtFa+FiyY/ofXj4q5GCTd7XWa5yuUj/BhWyqo0PG5LwuYahKQDvlH2bP
DV2pHv4qLsXhWQJHwMMtE2ITFxerjDeAaAd9wdo+B+3/GVEW4Q2P1mq7o3aTiZlBS9K1RCh7rzDK
3tbKRi93plDT/hjmNlhS5iU5kta/J/ckURiSkBDfCxWgS0CNs3NUJDAV9bDP57s4FgWEUoG+S5i4
JLJ0s3Ly9Df7GXjxJi8ELw0E6h9iVoz9444imkV35fLDK6iVufBn+NZUZn41hXmzO8udpti91EaB
QCTFpzfpJH3o5cRSJhu9TlVlVNSX1jYLbk791zm58iKB3kBm1u3JXvWOM07u5rBjNXF4k0cR68mk
hdvCMiRypZOizAtZqaij5ykj+DgUMejkgMjKYX+An8S2Y9bJRaR03JuvGbxgCamswBToPWDpU8+C
2jiztAwv+u0mK63ER/eiw/r4P9lmFE1bB2f+piDbhqq1+x8GJktoPN07sJU4UasHen/giCbPuZd5
e5QhzJPNeccYrOVXgbGYAwkgz46GVI7x39Q0kcILFi2ry50wsTytDdA96pMtT+oJSVHVQb7nZX5V
ajohqL2QfEXpznDaYrlwlDK5iZM4y9WceZjke5ejlZ5V2aoxtqyVDXRA7PHGy91fJafzthU24Hb8
mDVlqjWlxOLHWTvB3lvTkqJ5zA0YJf66J8ozBFHawEzzqiMFoXG3ugnOdWJO3Ki6gt5yA3RF77M9
F/sPBLUsPn5k4EcZxFzG1a1zVPAi8J/sV7Mk67FrcNGs2r2jjUdp+b3lICOtIWMtvZy1Ducioovw
68NujQWt6FeXfsHQfRwxItpuPYtkv8chPoWVBrSUV1IlnuTmAWqS37fwsc0fVUbRN3AgQIOCjBCH
P6J0jiV7oEoycSvuPuxqnKuewpnGKOWw0vW6AapV4ogrcGXGz3WqqWg+CTv5xWpzWqvRNqxWagi9
F/C5DmjwwMPm5xwk6NtC/o+pPHSQ2lvrr7RDJIKRfXSkMhtyGRKb/QeykFvShNDIgECbC/BUgV/Y
YQ19f/QVD+H8a1SbFWvEjG1zjTufITmu9OhaqVW8hExQE7bFjnHgaOlhgNgHY6cin5zzrs51g8vU
/O7lkjAyI7l0AausGbU/1dGjwwO7IlNA/89e4AU3cdP3zLwcNAdKgQ+zqXV498EGGGvpWJ4pIbyb
PHKVgZAbBHQzMoFbrjNVw8nPiTLuLqztX1WEpJdId5UtoxAuHKxIMW8FmrFXKWHNBqsmeEJEpWpR
B+7ShnPikuplBfcy/j8LSXrPYbOhfV3gaasPtQHY0e1SrY/2FiZXslfoPAfTgFv57ak6ZwEijRob
6nwc2L53jIeLnDB8oj6TyLL0FmspsxeYJxkGXdoepmm/KjPOLh1r5jTQMhRBUsG9QrSUxLKU5QGR
5Gn1Z+0+JwgkuUJbgxe0P4TxmLQPZOfrFGgD2NhdO5qfFaU6cnjf76HTebww+8eg7qvKRZJQs2uT
EAGq97whReTy97fwSwEDCZgAlTcF8HFWEIlhbJx5b6qsMKHg1ELLkjSZ9bRGDfSj39VDhMy1LLlV
lzBS684Tn7jiwZAlilHVPCZ9gbAcp+//5YjmCzzCUC7oRWxiksv5AEeDZ99Nspz9zTwCdO+GX34Q
OQZ8fxFqipHGT7X7tuioDAsK3s5GqOdRJONTsraZcZOTGWVVap/CfacSOHaFDXVyWujUdAqB80ZS
ARZEp+RLVmrnPFM96k/gS3p0cYWZsVxpPXQgebb3Lkg2F19/jvnjMsvWsHidyPXSvX3+LmOImdKe
gRKFyqb/QAYq5Sh91zJSsHVTMFob8b4nXNMbS5+a6iFj6wrr5LLw4mukkyNqVvhbBboV0rh600VB
4rb2QdFLop4pATVmwtR//MrbRdtNprjF4YBlSwZD1HEBUVqALsCQX21mRVl+nmIpPQ5ifoSAJwPw
d7SYft1ArLfx949LEqCRkaj5rs1SthpXlfkfcgBY0C/sdIvaRtmdJ+UZygNjYs2XZv4rOw+n5kJ2
p/ZbELGIiSpehLBOCAVEy6IyfnJ5R1vwfK5J4LCZ3IYKl7KoppaCY9MUNwJSTZrVOJsMohDwuu2y
HxeeaF0wcIni7chBMwsSI/UVeG8u6oPtlqzb3iqZd+Hukwmkod/Kiqowomw07a8IoY8uSeYWQPVO
71+zPopglqEuea794qGbYb5kQ+LSGv63r6xArrr5/cJyW/jiiU4gNO+DjdwFK3Ok1EevtjN7WDL0
ShYjfqgcle0pVoHq7cbdBDfkknItusiCWh61HrnEfogjxki8h+LnS+vWVw7asrjBz91R1MEgp9U4
+bMZt57TcoGDPq4yTmoJZJQPsF6LWbhxfa105TYeb780hPVXnvGsNw37TUvBQPrJlEQK1WBi2XqL
14J+mmvpQlcRgdw0h0qyi2rGG0QCWBxoY5cw64u9SlQDhtPPIYaxK1mcx10UAIVKtjIyCNuQpqfL
K56onWz9pWPtTaUzXCOWLCvaNBj4l/ohNenbGh42BlwASfNPcKRhsu1EPchvAK0zEl9TVSs4S180
tgVmCZbHPx53PEKY/aBzExT4yVOlf2Td+NivVOpX1v6gJuCehfgNKFCeELyN1+o640sEv6Yq7hRO
C2FafgxRkZKLWWRg/hDDuG4Vf/9cWMJ0w0pTa6ltHyvBoPwqeQSxOm+d7OHGrSs+nB2bKJhgxKvQ
Vmq/CnpNIvj7yrGnPYx4uJltixOCwdyAIREX9fvt/B9UjASFFG9Hld8aXAec5Q4baV2mxMY9UDXk
PFV99JoSY6IqeA6NFyGK060GAOori4DF8DVVlLjXIgnm7QDgWF/ML3/g2t601x365Pe/znuO1v0U
TK83EMuoL05PJz/lateDOMmDBaMX2O0OH0jxtYtUeYbzCx4zNMZRfnX5VYf5JTF+PbN/ylEj1We8
BZ2Vpd+TG6Q3coubV0JzsDJ+9PyShRRnkTRqQkT8dLpK/XFMiqs7U36Y+XsHghRNaGpbjH2N5k0p
9Lx4+HAMLQk5PCqonSpIl2wgJXQ9NzjpOBFIjC7A/eOO3FTi2BFbvZDKGoFiTX/hREyZ7Quj9iW/
WfwRGvFk/VwuGfC9cuA6m4JYT++ECywqP9DxnjpOc/K/rwy7kk97V/UTL/Nf5nf6F8+e78OoAFVW
V4UjeAOhUdjSVce0lk7bJZkRbmDBCSlpXxNySfT22KSgJQUc6zHiEIdOjwpCbp6fqrH0rI+dfw/k
MYSYCuydLtk4ARvraWS8JYlKnWgXdj/uftH0gzuLNvydbIMHYI1uOKgyhUQDyS/C9+XtE3qV3AqD
GeHZFNx4i3u5Z8EXExps43AQzVjB22eyxihpg3zJVtd0Xfw+zryPSv2l4GQQRgIcS4OmA8zpQN+H
FKPZqgEJwcHM8gbiT5ToxEGRw0nMHaKbFvNN1T1GsFelyalFErSR+dfBPfMpKo0rUV1w/EX+ykyV
dTebiUdyZmFPKFWrTfj6VQKXtTFyyx+x7iFu38aA3rWv1/2gyoorDCH8kMXrFNfqD44Bitns0sNd
Vlgc2WdxTu/u99odeb1+FJ2m26hki9CoAaNKQNZYd6Q/Pz4dRKzBuoNcU0sqHSpoNGZ/60Ivg53f
SMZyeTdtzsOyUi23PKePHN5l+sgwpZ9P5krqv8peMSxAdQXLBj0vR9YtFl3Q7JOJxO1/3Q3R6qLV
OoRo8VTcnqSsHSbv3KPjeY8J2thULhX7kWCCTyImDDfhT069RLi33P+fPeLBg4YewwthnWMsC9Vg
kXnhmvYJdzdKELoEaJ30do+M9WUOue4ENU7UqYOwcUN0PcTpwuykPjvN41BDSglIqFkZphbh8Dqt
pLLp3Yiu4vXJTd3a1SBMR1V6Ts39WUUze3vIs9ehJfZjdT1tbnODhkG1Jlzwn2YqyEt7Iu+TcOFB
bQYl2HNyjg/OsolcyMGzbNl7EKbc5b+k9Bm01+oDZMQYaqYBY2+nCVxaGjBJrsJP2Zd6jGZOP0s4
BvEKiuJryV7kMOyKBG/m1Cwc1cB4suCe5kE9b3y6TfYyAyhPnDhCSlwpSiXN7LwnoIY+x01fiB4V
OD1W8Wig1UtRgBOX3xSYw2IGd7Wb0NNvKbQIbGLqbX9Zfps1g86Ljn/dGsDrJJyArnAGSJ/E4H0h
QFcyYQ0jZea1wQTvdstrULtbhpdYMAtrkhWl8Uof6zK7aE7L8z/sL0PT4vgrdQD0t3ZTJ4YXjQEW
YSNRmZww6u+ue8JiPNjT6g/cWltj/XYUW+6XxBNTMjwyx/oXskHK7NJ/4ypFmCaiSFyIle9eiwaz
PxQWWTa5XHX8O9zRqg/46dRQDITQB8DnmDlMSW/bXMfMKMZTi2kRziD9JFwxoCHPEixWsctEE1lA
9DTFrVSEK+r2PthiqDSTqa1S2mLOGopG5+KLhr+isbn9azDt+MG+208djxoPKFvbqO6czdEZBKyn
bcOotYyW2pvmrjWpLV+KbGMDUYcppir6DFJ+hIG7xXq3zckM7MTWp2kFXQSM8Ve9y5zMAC9VTl6D
hFklmLa716K7s6NxTezqortb7SKT7S4TjMz2LTVCcc+nSChQIYdMvQoQQN52zCqhgSQ85KrkGZXE
3UbpzUr+ctJX5+Bv/SbpGsfAZiDLGxJD8Hpj4OVAB2ZXaK604hNUfdIEjU/07AwPUqlf3VJLECvK
QZbazVlTDF+fySNbO+rRZTg0kcyWzkbKGel1wuzlV+EIp2R01in/DATtmlFeCYhuhKpV00TcoY0M
E0C73uCRbbRqSyY/x7lMIpgT7+5KA9nLSutm3HTsvekjlu4Ihvi1ch9tO3jdLxBVNFt95y2p+o23
pEwtSa8V4Rf2V973RHBhOm96QJqpWNL3T7z8ixi+qSG5cYDlUOt49I3+CLyRhzrcxJjM8lqfz0Qq
69UX6OY7CZM4w9rEcwxKtQ5PX02bNMbok9cSkuXS8tetZCa7Ic95EZb7zNflpMXTYCHDIPU1i/Zl
D+BFSXzC4tIKRVR243nGMgmZ65yTq3mYpNTYibrhzlNJiZ/YgNuddG+uoZfslVpg08T3/kKQDIlv
6hTaj23HAO7o3efqnsC2J3llHj2TNjeAbIv28Vf01r+3p6RHhUTnae7n3TxA6JhYpF2did0cpOS4
k3vWv6LrjZxxXro9fvqvL2QjIptuDPmxgYmP6geXZe+CWvqSrHWi/2HzmGL88SylSi4tRtSw6Ct6
4xL9h108m8JEoA38dpKtmQylN/41Rjoe2h3YMX+o1WII2mVOGFJOx+eb4x+H4LXkn95uUrYaR9ny
1mRcsbh7U8Z3ie2t0EqjWoH4eHQLweM0HLbP23VdrLsFWhxmmCSvv56VwL9Qewykvh2zsu5DQ5o+
5e2RqWjcc4B045Ndh53sPAu6PmRWmP5JeTkockPTPwZEek8bU0lnCo5codorMkxQX4cvbkjXYoDZ
JOveXcWrg8X37PS/GllTkM5cwAkrsWVxqMmA+yHdMh7H59X97u1/sLymnk+8GadCGH7tadmGLTqC
o9RTeB9Fv325Mv4UJKUtxxQ9T7zQER/r2NAY9wpGIkJiav5bpBe58yM6ObReeAzmy32Uob0aHO1Z
Kdv7erihqa2v+1BwraKWI5lAKVCyiPj6MH5xbAEnzsZ5OKdsbPUfz4Tji40ykSBUujbx5czLvdY7
O0qmtMHIoWXVW4YWQ4sIbZKTZzY/ElCHUi7XbqIsw5O+KxS0BLHuWUY/WLWe/5YmHkzCyV0zi+Ra
K4Cg3OtyYuB5C8PMAT4gn/4t70LM+ANmENfboPbR3jhUk0RxEYEi+QZo4vJV7Tup/I0txd/7oWi9
x4jFVFSUV+5/fBKbnJph1wlN/fLYvGGmBUCdPw7oXYDdOc4UKSx+dfaeeNp0qyRMRiwyp+thKfAH
vwosNjwdBIDmODvK3pgTccXf7zc+ovgwyq40FfpwhDb+H8PUuYVtElFycIYPesed3HV8Opyw7dn1
URfI3/eqo8o4083OA5tkSVr65pHp57s8uK7nBHSxGSy9gApasnXO8UrbgfJa6OicOK0j2Qpa93M7
BzLF9AJNRZVxWtM5NbsTaEWGZZ0F1q+Kz7hLh4Ao+fj3covDSeE3Yq7KiBq9LYdXFCV6QRMr6p/Y
2MLzzEEXdMyzaIu7OCVfFRGavsMZqnHDWZDMZg4kCYeULkCCdzGNjTzB+26zXzl2CInkCNxAcbUm
cFgX5aDmulTtgvF5INEmYw9P8BEqOnRXKsJKKkHxnp3b5JY0kJCYOcbUgtg+Jof18jRi2hopYAvg
pDAitNvN8cDRmKRcmo3+Uy0mcIoewpyLShZU/m6XIJiEvuAxJmPZYjp++7T5dtaX1IdkG8fpsoRL
Kc7JOej4DoiCsbYVvn0cfEkq98CS4iv+6XOE+/fpk3ilzb62HTmokFiogrLuGrvnX6McjpUCJYqx
j0tS56AbVErLFrUQ5UbHPhpItmD0ULETGDy7RfEBMuoOupIyp8zlwyVAG2W3M4rNhK985AFqeMuU
4HgmuREh3OogjpIMMIEHXWhG18F8c1ehUvQ6xcO6W1JyyFxciwLIGlLK9KJ0ZgBvbKRhDcyzkiNI
S9BUvn8uQUj2ELT77f5B0dp84ztF6mHjyQT3Yu2sKW/7PB6hqcvlh1ue85RX83M7aYUGzevc+WwV
Z9nuwGKDhLI3rV2ApMPl/hFiSIvmG8Q3uQoltKxjenmPJxJGE8oIyN8btsa3nMLdgX8JMHJizcVG
wpoylfgBCBv5ymU7t/bQ/5Ve3fXaa/D5hqM5bG1bIyg80xydgrz0BVq/h47UvQYJrHj31VP6JTAT
3Fv1wJPu9ldvzqyFvWa3XPgl8LKy2PgpS3EEPZqk3XeeLaHP4sa+bIHqs56rD3cgnlq1FrgBeoPG
T+4UIExgosn/l/6UUu56JlKSGd3eYNereXZf2mGesEOtbR7w+SVf8MR5qzLBJxR/5SZbDJZuT5R6
TRkG3xQ+HMALKbs+O6ohPnjnXCFNziMET5ocv51owEYSiPPSKueLtOBDhUF4OsLRJZYdZh/OJ/zG
vuVxH3SgAWZoPupfaq7k/kcn+aniTevbpwkyDgcLS2CHVZEbsFED1HOqJD+co5Z9pCe9tIutoVzF
0DCEMqtd7HU4DVCCSKj4dTHGRr/n5jgRGiztwRXjIqqL2LK68BJLG9yahiRfO3KtlG+r02G53I4T
nzOE4to9DJmF66BofSYw4rHefrE4Ti9MIQH0kypkQTUtkC0IvCqKGlGWgUJrambSkTRUWk6j0AHc
qf+nCndqTvn0v/0iIes94zUAjJnK9B8NixIwILXZ/Z4Y6tF2GwQLwTheJ5bBFlI6qkphtESU8DIc
YtKWuZh504vQHAGjn5QN6craJFGCPwclZ8JukYzR1UgIF8zg+ud4UtieriBCljqdqC579Zjlj0X1
1j81qnYBjGEvz8ayhj1pJ24rRLPeomWVYAb+aRuuGg5tX3OkB5gBEbCH4dRidTKbc7poDok119EA
FKYioxXOn8MiNebHET/lPoSoirQvKL6tSUdTbbh45Lfl1gK3xFw1MG6y/Wffxax3J9wQobR9XZ7v
9qKubI1afBLDudlyHkeB8zPKRKlXccsnOdlUV9jO9q5JFuc9IPXntpI8YedDb2n8Yk3sZr54fOWZ
dmbtwfaf+pDhkQU3fy+mAarrC0cJaaorVjOYXATHykz/EQH0BwcuJgnNCmvy8XDOB5PlQZvPkley
jgI5a1Z+YKjMa5TfnjIsg9fKXoKUXizICU1uztdI+Q8tOwOr8QsQHiBDl8cH7if8AEopX3YeiZf4
acORvyHj6dMFlN9GBmP81UZVgFapry6v4pEo7689aqIqSlhZQEyH4gvUEAsvvrTQ/wJmt9/tUD8J
T1q31uMA63gN6Oq5ECtSH+KXlo0FRkhKCodX+Hta2PgfCJ6BXwNEq7ffZJBYnMP0FexfreHafyOa
YAvf/0DTWvVeCGN5IZRAMnjMawLEZUIjEQ367ZE8e4r3d4F9hCfFNHuKqwPRvAxWbr7JS5AogT9n
0x4X4InWyjV01ehPGosOKA+8epF/1I9QWlPouLGF3MBbNwRpMd2onPK+A1VLKZ/8JJh7VdqsAfer
+O27V77AveZ6X7EJM0QkuUQRvA2ze7D+rPnA0eh3cJlUkknnB2FpvFC0kwOLD9vpvJqZBRtZNuVx
F5aJlmfBOu/NYLv2bKfvA/zh6awlkHa4y0zZhSND+pGgyuBZ9DUXmzsucjaIPbP77TFVkvbvt4ca
468HNEb/LQHi4QdZe9CJZDyDOMFzOWEITBS6VbRMjzZneQPQjYEGcpSh3zX5ERR77gA08PsBsBE7
8vY8QEFB8cXLI+fwqoNQfmQlvj7mZffLCJLQ8MdiSwmPnH0z1JYSTyYbA26v5V9EXu5lPnY0hj3/
TC1X0NhRyGHQQw+6GNrpVGGvE+NNECwXNxSaLcKBr2pPDhg5aBwo+z54fmdFFUDlM53Yek3tBNc1
xFb+mLwTCJiWdjT/DUYaPy8iqW14p1zr+UXkV6DvgEi1Mkl3WQRyIPeD+lBEKY5ScvnhdoZt80Wa
bwbZHaXKYpvMTwdaqLQyPkeROORD5UjiBBokwnO56WW4Io6bug9h50dz9zN62CEozVt/4WDwFPY7
Z2j7wYCgDPw3hgKcHj3/h2U38ohTXu372OLjmkBtV2VY2AHDMGbsyJZP5/xJ0N2tvUBTwgZLu3N3
15/7hS7dF+MjQN5SUByrdVwXuS2Q6Rg6u5b5Zka77eOVQDAVl3kLQMSnRafJBBUEgfRJHiYBx8+D
c/VAAW4TYvf5y/lEh9HAQBKYgIH1XNPie/sGrnXL49uhrKwBSmh+ktfe19AtYr3dY1M8jYCcpKFs
FHgj4lxPl1c0W1KZMuyLGHzKj63PUmYVoNKjUBygAsRok3YSCAZlxx87e/Bfv9ANCII+68pX/hCx
uQCvadHSPQ4ZB5+C7OdOz/Jy2151d67i3ymtpgEthfxsHhXfAwv6+gmPhPj40LKb7N+LZ9+GXz0Y
kEY3ROzfPtfDF1jcXpExHNz+fcjlfFsp2AXfnu7xNOj0l0Bykb+Iu1L88bpBVToxd5Tx6jP9qz0n
vyIYG+Wd7rGSjHy6HxNlEhMSSw12ZvKqUj8NiU9qdkaAm3mJvP51zHmyhT6gsMdhPp7KsiXJySnD
abR6Aqd5gxG+u8B6v/ZPe0zkf5Umt8rzBMrwgMpiLCgSEYDYSWuGxuSKtWBOjQQQLcPoIyuCTbWP
epR7Gq1y+2MIkhynz42QnfSDVPqZy8kGRIjPiNXr8lyMUBwxWP18PJtNtFHpQOrDLN9TFC3c1hJ6
3HfHPi9FEVUXx0+1XtQjeDvNiKj893xXrX0K8E3j92LnBjji0Vc+IeHZ5nIxfT+t6X5NKChvMD+F
QIuj1/88/E9Sz6vmISnS3um1N/j3oEDKYMYXOhn9VaPTYfpIZu3sfPhmFDxVkoNtf/ySExy7c36x
9SSUBJMTbsAJ6faGLfJnM9amJxWRa9+20T+898PLy5Yw0W97vcckqvyxgg3fBJpJYSES6u/PelIt
IGFhowAGkBIx90y29YtQIOrjmH1GDCluCRSYTy+s6F+T1B85hYqyOAkVsPlSWuTG/9O8hsK36n3s
zwvTqA6fY5MPaOigkYuBTvEISLVUaWYVksLN3Ok8hTbmbp4Qkgs2TqXP3gpvMJ45eiPT3J/z/6b4
hZh/TM+zpX2brXRkauVHcQnyzAzHHeKFKm8fAOL6ld9dvyONwUN2YRuPkqT6BwNYBNDlWE9OyzCx
VHryEIBo7CGhWZnCR4I88DUDfEJXMGYFHGbgoRAtKZJ3e75XGc/kSEG0lsgJmwlAdLcJeX85Qb4f
ypX7DSmG0vSmFs4EcEfAXjrpKRIxDRqWeCZDIXn+XrbHvO67/6lGSREHP5XKqiRC2M/w+Qk/8rui
dwdKTGuJxGkFG7YJ1kTWBExQBE+9/gwheScg310l4mtL+D1V8n+hFeWt2MiRIZzJwLqcV6haeV3s
Bt5E/2ImNO7+xSA+d48q+xFxSyiiA59vV4XX8IN7cIDp6xZ0Rby5SZyPWYu4RxBTYj8C8pw/iruA
ink8Y04hF5/AJ7hES7V0K2GOHoDpcr72NXiFXzyIqMh4jkqwZ6PmRJg2F06N8qTauyFdfVUcyNkU
wAx5dNAryjEfPSvyQAhjd0v3tCsxs2KOFr89ypwY5yPvweUSominF+aPgbOGkozOMdKTqbYBhyDY
i+8DwCwP/iprQmTNboGwipTNgZIKUBW6Z9Qu6qBIqeME12LC7ulkFm87j+mzCsAji0AzXq2JKRku
0MCSRyGf7tFEXDeLIIgDTcoQ9ohBjx8YNXe0E71+wAou30Os5V7nAHTMsupsLtrN6ygq8NWUi6qe
Rya/8KATBuEGYU0w1vaTFh6PSCTSUHb7T7/hSQsOXceQXEq+uN61RQIUfh3wykdz9oT51HUGW/GA
8EWXomxZGhxa1N3E+3IEc5LXOfm3JQ0dyPeUmMmOEgWfJaqT539zijd5cSUubycmUoBJXi7M8Uay
Rab65o9I5mSYU1BkFlv7Arbhn6CghubjwHCNadTfIIpKJ15M/ArtkSYyMgCvDphmPaBMdNjgSZS7
EKz4qnGDETkD00RDuO82vLGvKP36sBSEdAKQKAk/Htydwdjnzow4q3ZVl8IEtdCZxwYPOW2OZNPR
SMFyWzmSf+rUhYahbMPnfAs7EuUn18UlDZ09/0zrG+qiAsbuDbtTLK5hxMpEBWgYFrrnjUMdZ4E4
7bBP6RShNoRfwK/7+ZimPzGXBi6oRLTiQ4fm39uOoP74Tj1SgZLaPNbu8Wkac8qgiRRGiee43kle
CeOp/YKbHrFrGR5B3NX8KL2rbtomWbYf0OA/CwtTSqydzRRPLzG6mcTvNA2DQqe4/aLZyfkSEw/b
FuktUGSZRIUkOKfrojX5e0BGOmVREvsBbLVsIn7XYkIrnW0HDv6LyDa84SDN/dPt8K6gMNpijJrS
YVVNA58hdwSYook84eSHoNlHUhgQRePF3MLgZIpvLX0MBc4imq30ws0jldPXt+cc52IuOfVlxEw8
lR5d7vbmm7QcbAiXBPkb6VnC9vVEMw/o5WI3dlrLGq7FgxPI3AgK+ZMmi15m9gJc4ezIU6ZcVWSH
3R3AYO4jFU3AOmQTofgzX1VsxVc/SVzJKqutBbZFgk5BCcbjQZ4J53OTISk8U5UJ2sLvearAuGJP
TP7ZgS/U+l0BEQkGqEpXjAq1q8mhsCk/dpM+q7m7pBV+ngAitcCSPuz/o1YIReOrmTG4vjAYpfIL
PWPFEEYabm3fVngs75v7UfMHQENEc03kpmNIiSd4ZJs/svciGmYnGbUCvhL7DgXrL4Omz9T6Eywv
nslln1cvZKHCPLeYGBqGcJoRAzELRpNBZ8jXm2r+ZOTb0WJkID3o12rsw6eiMw5lZB+i9At0EliB
wdXKnSGiD9OY9nUYvdQCRYZmMrzfez/VIZPYIUp6mUvIXdsmgtTuE9+srCxsQWDIsn3lZhNq/v7f
AmDjhav0EBOoaG9j5r4aDDa4qs9654Q7mvgUaSEXVmKN24hVLMW5IxEeBksn//q7Rq/aD21aWkM3
+oi0uRYift4Cpku0rE1C+vYSxYzosYtpn9iWGErssfNBVINh0aLG3lANC5R5mlCR5c946LjNXAjR
g4wBA+OhlpHfXoglP6CRxLaHF4mdLYBLZRIVpq8+Jwr0GE+jscJkOcN+CT08zJDC5u7ZPtfk0Mk7
nk38WKUDLHX2HM95Y96JMG5bF06VELnw++x8y0VyB8mWMdkApDyI2qlBsIXW+UTQrq4DEU1G92j0
O7r62pv6StbAcoyxbEZmt7bx6vOe7DzKTtoxjWU9Ut0o2yHeJjKOKRFvQCHs/b6DB8esgFFce9gT
dA2FdtZIrW7ULXtCOMeTwkfIyONm3D2hMyp21cS4aUfMBs45GVrJqUkkL6YGlSjPOpueO0hWxO8o
6OTW/Ftr0vyz9Z/Wjtkm+AnHJMdetQPhrW5nhgnc7HiJbajGJLxHUg0ITDnjD62D9/6gHa6yyoQ0
P5tDnsUGHNmol+2HGHoWpXaUMkj2ZwPyYI76YBHECJicdJeg2s8xO8zIaiImbSLCnFw0rQrAYJsh
xUoQJkkqQXnAgTSkHmpNqWZfR4bU9UETNIyeL0BFm6vL3La26d3qls+uSH4m8oUGHlNpyPj9dpf4
rL28FGgtqBzgi/XyUtzLLAAxX+C0Yzp0qZZ9slh7zNMjJiaQMArbszvARVVN7FK0E935p+7/Pb1H
MGy4cePsSGTkpq6cReLCRCRp8q0T43OVoxY/GCB3LnIKz32F9vS2dSyrnaB8YtlQ2CFNOSWUf7uB
YjLMOo/1WwDoiNF7ZRnXjUTYiqM7498EORpbCI/3UxLwGqYBnjngOp0R/kVx8PaFvwjptG9iFnbl
QuCtvSo4Glyh8KaBmTX7Ydms53cenMGLFRFhRFzSFSv7yGOQh1gNm9SUVsxcjh1vjm9XU2ixyC2n
Vc2ZslSS1vZyMjldSLHdmDaenRUpF3eJlhBn4ary/lMbb9w3baz6UG0mGtGmvVwhI0vjiV048wW+
kQnBJLQWU1q8pyDS6nca2aXn0kO2Hr67ProquZKJgQwBzx9eVAjYDF1pTTrkOFioVoXNGU2svmIC
DLAOUHCczpsx8aAZJsg0zedrWZMZiVUnC+QvwINp/DCb16p/nA8+n9hBTAvtpH2ziK3yuRMMoc+v
T7Dt9pLmN9T/LA+GoheedaLaWEDZz4Dd9IvBcRulDeZPMJixpFZbvfi6qTklWQrW/SL7pKeBen9l
t7Q+gNl5lA2hpbsJARHIg5AvugUPZZTIml3oMgA9YfaA7n9uptHVBSfsYERQM15foVUgsGHeBRbR
SPPQW8//bhz2WTYJXj/YMEwyTMQHjpg8GRyC9r1fOq6QbwY14sKa2Fz8ZzLVKiolVK4xLPLsNuIq
1KadaObQYDFTmf0hF8rcJEuWMHWwwYQy/wB6/+cc4Bt5ktECiIGJ9AmDubExJLQ8w+dE8rnzQI/u
c9s8giDUdslNL9d2VvM4pW85Ot0QNxAERvkKUHcuAC1Ju97IYejDW3IWMezxO1C1UxwMNTqAOvLA
Qef4moXl36EgoINMO2nkoV6FGDbF0Ike2eawjN4FI7Fd81VOjSupov6EPvGRhQmXNyUI3oErohJ+
zuk5Ai0Ytm9vWx0Glhl1+ueu4C/9mNI0BuMamxW50mbNeHwB7Vr4azoXETYhqkZwGoTRNYeeT6Me
f7mbzvSIoQiLuSAxkbtDQ8MxbKaqqHu+q1OqEK9OeYf5RDYzUQ1Kfx1zGTmBVdCSOJCEepnRJsLD
+lRDABUuJBAQcQE2DYcQsL+7rI+abHojwjT7M4a5RbwIbFjeX19ns4rUGBJyayb7Vxn59QtcZ5NZ
b5KwwcJZtU+iU/M7pT1EWzpVbqzzUQx3yfRUoPwqP6f8BdowXicB/IsFBSZXbXLkGaAyhpcsklWj
lGsX/64MGv4H0xBeXoyfda/1SO6RV211vis6CY5N5cxlLxtRrV7MjQHcAcWr6Y+RWq0icMVyOhUY
DGtGhkGDc6tXvt9X3D1OHTjQhOanQiUaaHXwR35zeK/rwJUt95Y8vkEZRuIMHZIoVt6c2Ad5Ocel
SEFMw4fsR5T7iAbv63LFZd2kC1XfKsIEPHKAWko5ed8vLujCUDyZ1s7FiqX/yUgqZl9YtnugDfTE
gRzEt6tx1TgzYlQG5/PTUi6nnkTcPUVCHFy2WISq1cy8PMQHztqJEM1fBo1Ad875/OzlTcH9pZAU
R1SVJByyegij8wONLNztHGT4nvxfIzxckBMycrZ5IU1TfiTO//rFfhvjAXLKjh/UDSLBD7plzwJi
Ts194sCcZ0/IDKkHgSRTU1cJhQESE+zEu/nVwRX+9RwsI7b/794Hvh9U6vvIRut+eQtb9pYCU3/5
BqKzQ5Zx+HztuOqS1wrBuJb/cPYRjIko2Jk8GtmzXSLzcUUbiPo3dA+HbCWnn1/nC9crhNJYvtxX
0O6truMLeq+r1Saxwyg3ge2JDU65EFxT82NbYWjjVr7hywAEXybXklsyonfCuOxaka4tXncBy5ng
0N8iHYcwWAnCDYrrKsHw9hNKYl8BwphB58M/I2Cy44y5YwRXM9Oc7k6RGVLyUcEHlbnm4PUiWoWs
Dwn2BUEHhOA2VFm6j6fcC5ayErdQbysues1eO4lEasFV9a1aDkyRBEWoGAzZaGRwXC3fYw88gwMz
tMEzLulMYuWZcMqsIi7Kgt6Y+VInJgugW9LHqTk9nr4Kw9TW710itbctVzQxbs7l72LgAb2Dlz4N
MEt/GlHIsCHVqBEH3QH0IjuSVgbBoe1K9G+zZQi82FPz/cLiQ1yHDP8cN47FnIzVn/kw1DSNMEx6
RhuY4phOH2QUFS+Ig9V7z5f0r4j7DGoQ77rUCERZjrGphsi2IM6hufjKAm2Z+pBorHXFrAK/NGub
UGGsz82MISNagfOT8sfUGXETcx7QhybYPInYyp4e8wWSoCgct8y2Vu8T27ZfevzaxgjkDpCuxK+t
x//xfgUABscKhXED/lNF5n9lV1+IdNE015ieoQpJMpohmzop9otZEbBDVcDY1cdkyVhuEO/i6LVx
6smqHQItMEv5JZ3a3ffCnU04wPm8qSgsWww0cCLu1osH0Mhd6fkH9XHPeUanCE1tTU5AnhN9j49c
vuSf9UipqfF4Gf3zhX+L2zK04tzsArAPR+5GAmb5iqPZq78EKFyO28K3I3PKCVgGPs60s9QFpVLH
XQelnE/mfPGilJ6/DLJ1BOrMPh7viawctuIORleUFa3ZhhnCY10yv30Ykba+PLIi+rX5VqNpgdra
InfKIsVNwCtmPyXOfEk3YX57hMDohu5kSoJh9VNCzxUPfWy7jj4xBi+IB3YJLxTW2K74NohElTpf
ShftEVoZX2w10EXjqaOaJ1Msx8K+9gGODUr+8cwPH+wzIyp1mWjK2bMHsuTy6Gx/jmngNlnLegJ+
JxwUP4UyasOxFLS0xUKkjVoDuCrGhNH6fTahrWtrZQ9LPvhmIZ6eXCpFpUlOKLHNh6SRzujhmHxf
nh1mKU8lyNshEFkbpiUYtgo9VrfdnniWlzQaNPq7yVXaER+/8hfHWuQE16Q3mAAuMYrQGD3uROuK
1ijbLFSXIDKUFO05fZCGO15EoRqUfqKp16LeT21BOGS47maGQDunfNnc7P/QEpy5dqXRnqg1WAar
/SyViWW55qGgh97TYCzh3P2JaFDWT2T2KXXFlXtyYtTgpF2nS4bVrA3M73GPlIkhXXjlPk1kfWMh
69jDLl5WW3YA8Kyhl+JcfHwh6eHRPSl5ksKMRiUs6S2HuO0n47mqi+/ofTMDj0+NxVT/RMcEe62s
lZC6SzfyOrEoyoqExGnVEpK7jZajpJoYcy1OOzTos1JT7x3ZoQJgi3B5mBXjAmD6T4JFItC463pH
EnrAwXKZJSBqTYzephiopNRw6QpD5oymqURKxvTiTD4KI7nqW0LyXG9jLmGEOCj/21lo1HP1hz4S
gtU/aFuUVHJA9eHlp1fGdSqrBHqCjCqLvNI3EfKMfuPBSCrCepwjfvK9+acjOFOdaJUNC0EGoO8r
PRvIyJGlH3GhEKFMB+yUCdiIpimekgT2OCdpf3q5MCkNX+Hm+s/YW/8bPJ7ev8Y4ZpJCkQUhsR6H
zytUPHMly03gurRwjdd6bufhrF9WPhCsVKcqFgkl8JeBT+6oIbIB54AuvalgtwEpfyFoYbq3QXxG
Z+2DxAWnJHm+Z95a+39XMl9BcA+AaMTFqZM4Ca7fremkBYulLdFoVwVLBWqoPS1qhec/9SJMKgcr
5zxbX4n4CDlHt3KT3datjja9ykI91rRmboCZ0FvFsjkH2e2R0cIVTb2V2OQsC/1RTFSLA6eo7A4p
yqq4jfmxOk0AY85C89SwrrA2nSNJo6P+6tWvk6TfVSM2UzIvD4g1f4DPY9Poo7woVyzciEWFAsTJ
xlzCrZQLQhKtt6DC4xAYGl2BmrETSpCRKLAast89kELBstHbaNDLsV8dUF7C/L6sEq0yRiuuwJ0k
Waav83lqBemvFn1pabKkqWWsdbZCmqXT43EDLiq/tCN2WPPiYuXg2FjD/HXXKbTXqXtqNdRm4aQI
BLc1n6HwqrUuRGDDlCEML0UmOWXYrC56cJMI/0ELAk/scBe5R5nnWqdggsmiC1y3f7BG2UYMJOD+
zlFusUBY5O/F64qIJHz93pv9gydQur67OO+xy6t0gBwPkomDxc6Qnl2ixrUaB8SjWV7G1jBFSt5B
oVMsdfAbmyQI0PzLONV/jU1Vd8ak5BJ4sbNipArKM+kv1qGah3ZXkN3xRni76+N0UlN7sOz767w7
arpmvyny7Egn4UCZmOz2QC7MtNDTGmwz5ZCnzT0+vIFG/TSTMA0XmuWIn+uMejPx/OrtaS9tRPec
cAg473XVZuLnbM9v62pUZ4wO9gWF0DE924i3QR5CnZsdnupCdCv+hAtMIqZ+KZ9CTxdlM5lOhUBO
9obbjc7xGMgpzTZZN1uVbRSf2Zb0FYvwLa0nnYzQiyh8Lb5xoFEy/nVLjeqTUwBl5stY5ZTOMQAW
FkMYHIWMUdBLNi96aCD3ndJLqQsnxEk75D7nL+M8/c/rC6l2/ChXv8lqIbTwWqVF/jJ1pJQbV5tb
VbZXPQDHc4Q+uEI4wcxtZDmvwiIP1GnFM87oOx3USjQESDOUgZ6jO4rS1SovKLkMLjQmCO2khRsy
P6YmWWKsvystse5MhfYLFWRgfrP6DPVzl+IUu+8vAq5SEbtftVlQEkzOmBDkE9tTVjZK01HD/iHY
StEqxXZ8XI+MKkbKlwjxow8BR3n5NGbKmKqaB0LZ/2/mxZ38mRfFU7Q5I6zkB2U12zlDKxEfSqby
QVdSiz6EKBN8fZZ6FlIBeh7R0oCVAS9/G3nBdK58ahAx1KOHvgyfXTeBC6hnv0vvnkxuxJyxvTFa
Okr+FBkpsWgE8WXNrIHJ9mWjcBG8hnkgF+JLGFDS3Ri/rjHUhyT/58vTfH26tw17aw7l1AFZd/+m
7gjkHUVxYmPV/ogRovnJlNAiM1L/O+3U6qs+Td7YatrJAMPHUvRcbaAKBK03RD3ezlXJnfD0tg3M
cC1EyN/S2S9anBbGyirkttHINojaMUxqURrHL6Q8PNTvrZDGl/z3c5yEkexoPhCFg43COFBM6Hfq
ztMqTt8l1AkGXUstWx1ns1/keEHhpOab132W3PUa9qpbhSU1yrfsemaBUf2MaZJSGpv/09sBOLcu
kDT8q+2DA4i6DEw6TYYrcu+AUVeghryV8DwTd6eDmysKhJZShY7CDYqmwJrs6g9jrN42mUQSnGNt
bZJYfKkrfFGSFmGXaWbwFTjfYLza0oFCSrlT6q6pE3AlzSyy/1zcboPIKISZ6EPcx82HzXeGXhRD
Fcc1kG+/piIPspEAQxISJUSmyFNyBOPRh3ZkFeFgJc0ocOXuNKsTpOGTdQYOMqJshEQNi1lk/mYp
pDQiQhML7QW9DVqyEndmGSjvvr1MatO/BfteDxfIj9SItA9vugTKpdA7MA+DOEr2oV4ND0SvOmZ1
J0sUVWT+bR1YiMyWcOtYwtTKTqdVicJtQtAEp6IvkqD3msVlgkF4Ahk+cn3b2s5IDhC8nuxa4IXA
Cscgwe7krpMZxXOVUvEiMRp78nDbbpZ3VrkqHDDXqrv52PTIi6r9JZIQNnhG5pwpTYmm3645vxzo
rdb8gnfbIaqSLpXDkAi7/zhjXYfirnz5DqPGRwlxo6uanzXNo6jj0inJiqerKZi31Yyn1BR9I7ju
/E5MnGksQvDZskA39uIIqHHx2lByIiC57NUepw9SYAKofqGbbMZXPtgbSIicq6zC32XLcZalJX55
RaSqOzjEVqrmWpWNnj/iVJNpUMMIBforFmIzJBCi6Ukipz6YH3wgf9+hibWTU6w5aR+1J/hQfFgk
p3PMF+UzVmksfsZDCgrReHN5cmVP8Opi+tZJyau/6osVh09x4B3ENSIC4feZVE32E9QBpbXO2nNm
iLQLBTxdsEi0+Sjz9RaUSg/NLvdeLEBTv6WBUuaejivAF+Ww1ezRj0m87fuUZfr6TfzchMSHir6v
eSxW1f/y50GCAac5mgsblnqSrLwDr4EjsFlP3dSA2WZOh8vIcve7bqGiCPofrC3rEF6clILZJs3o
gKQsj9JR9dN0PObPiYyWx8cl35I7bMvXNhKshj2VGy480A0o1ijrvYjnElPzA520OuoYl4h6Ejrt
pMWmxUgwNmplvxqpW29cvACDGTGQOh17+j6Gqoby/7keGbVAwgoWee1Ann2IIK1Lm7UVAWCZJ0A4
rbJbdW70KX9RYOf4C59G2oM/80yu9u6JuMjA9wxKFHcOyegApscsnT7XRjeHgAYdmxAvIrz8bEuW
PdidP4Yc4iI6xIx+wdop3jWvQ5tfM3NhkrIwlr2LQ9fX1HQhjfdOpfWkS5mK2te0sqDP7eMoWNq1
J6ZUDsXsVan7wlTvvfqQ6Dl5ZXCTekQRlhisRX69mkFhr4SsKSMjsS2+6q5UD4EOvLcAWikWC+OI
WTESinu+Lqm66z3gBgNtln54TPtt1kM5+kyV6O6ybiezRVWmrB89TfsB5D3emSbgfBEPEzd6+hhz
Ph6NnMfYj5CZiTKx+369IOikN2nuBOCX5sCJPeQEWNBLGmddqAIO0jKxtNIuRLu+4c4SVtcsiRgi
dkSJd6q6Wiy/NcDFBK+vlHYTOqDltOIvPCG8DbAHdVsYghqkHYYlrOMzmnWSIKrVHznYSQ5bnZgp
rFaLwq+iOD8t80Fh5vP8pQDHAzMYlyhNGCn2vLS22LZ6QcnQAI4bvT0/+FYU5JcHzFZK2j5kDFNU
rMWTnjrj6uUzZqlw1cIjYnGO/S+5ra7fXvSdg3idse2fO00OrNykSXVceWm0ElMDrulKf2s50b9V
oGgM0+pesi3YkmLVWl1ZwwyUmL7ettgjb8OIswYrJvmrwjzeKu+HJHBLGXHlf1ehPOVEvDRoV2+s
iBbp68HCe4vR73ZPA201Upgi4mEFO8RCCZ0EiRdKGLBuuQPpqOnGJTKK+oJfG3BvEaK0a/wgpnmc
Y8j33oa3lqFlnjChYhrqVAxDI7mE1yHEomijI3csi186ay8+iZXjrfGmcGFsBUYcgjuCcKp7jC/G
DWQUiBIn3rl3kaqyRiu1Eu+tdhTL9yfnFhlW9tJwAwQPTHPVi55H4SFuTyQ5BTnSJ29K7U/fZ2mK
IkwI87ZfQGvvJL4kJ+4DnrS+7dgs6mJMDamuvlX36/xMWwyKtZRwup4ioWIv6yr+pYlM1Jo5pjlM
z/sXZSoppa8CCiA3fAf5z+sDEJ7FL7VG7qDcNsG/6SUM6B+srVkwPeiE273BQSrzqVaZ3g5CMQOa
wzANU47d3dMNLNOiMgSBOS4CnZYAyrc/jxwJvOB5RQXvah6pHjCyW5c4vkqr4HC9sMzCa26tCfvO
3/HS1lr0euZqZX0ixSuz6OATaU4a31IIKpcDaim1JLL3EScOfaZkOm0fB4MjfOPzFB2i9M6+V2WW
lP1lWz1T4Vg2c3sxG0+fdjFw0bS7oUPWaWmi/zxDwC4fmL7Gb7SuOJ+qrq+edoA4EJQHB+NmSpzB
qap7enrysnxPiRSznz+XqYgkOVBAvAjj6k+cTzsOxvHf89CPLlRxn2Bz4CEs7bbU8g4I+rKVcoLi
q8O/5NoxATTp5+9hIEphqtgl8KiXlkyrnr9v+q/gEUsA0oP5zsX2XG1hnmBW3Zq+8g6pqdGSXEdO
y0R8N/W4tPaVwGerFwl1f+XX03vFKJwp4z8kH2tlLPskB0g2M810D3+j/yyDHXfmz3KsBSuNoXao
nYRTwrvAnG0z9YRZCyHX65aD2Dd6CA6j314BBUCsWXa9qtj/6UXF2AjrJHwfKWp7BZWvuOrvwx4C
JWFUWA1CwNWQpMLRRWkvuaw9zivJlVqkXir0VR0aeDEbLHBljQBzSvoYWns7IO6Yp09QnmX9Z1py
oaEMu7CDFztUzQ69GVELiXfp/7v9eUsbYnR+S6cgIFOVuwnW17hj1i7GG7I3si0s1s/EsGnQoG1B
HbL1+0iA7axRS5b0vnbu2XXukIJZ1G3TN3w5M8fC4Nu71sAL6/UDhi3htlMLOQ+gRtw4P2KStyMW
4+bWb9NC6SEBonuMZDfJ8fFrzGgq1usUzLwg7GS0Lx7nqqRV98O2nH0mrF8XC7y3Qyiro2zkAW2i
uowjAaqFPm8I6ruOOlk73mJ7bWfrmW48g+KWBCG2DKd9Yoq//TsJPB6d/4fLELqZ3tvcfbRdHa+z
E/rgKub/tQzILZCjF8qinPxti3mMQl1ZTIxnMh1s1CPVuOV+GC3PPAvkNbgqbwp7WMcqi60N0+H4
mVETnd0EYptDCahcSv30Q6kwnoKBReO3UJ4+FVG0xr3jkdRMrO9EbVJIzRKutkaRQKRFjEHHQcXQ
y88HrhN3F6Iv3X3afzjDbXl2bf55j8v+3Lfq2Fec3G6c9ioueRT9rZu9657Ig2eRaXpKRP/uR83b
oSj7uK9rAoXCAr98Eh4+YqdgT3j/OE3A10JRjCmhQ90JQxNjhXwHZK9tWE3XWGsKnv1Tu1KUVMkX
5OlhihxI6eVrLgjSyta8KXxe+lAPPKj3t0ysbOhSCzWV6RJoio55JtXekVEB9seiaBUONuSie3ck
Lua0CMaNrcPFqJkI7r+5mzjBuXhL3A+pTQAZ1Z8ti196LG6Ea7h1UoThR1uzAFGcVGewWv871jYg
xFNYy+sl/tNmcAZVa4sey7iZcxZPH9oNPLBqAJjuOiSbp3pofYOTMFPGZaHbBZwNtrBFtWj7B2oA
DRsUpoxZ1jXDDy02xntoz53Aj4WgJpmAK4PdRJXIaapxgTaFQgFCIUv+cC//xN3o+Is+vxCBwoBM
e3lLFTH1yg9rQ8C71y6aKAQepp1Dr87grT+1ibN67776q02JFZ8bcGE1D/sNzuGqkYm7tWQA/NGN
x9qXHfWq3A9j6X5Kr1DpOcl2sBABYsb9XRxY5G05I5ZdRVhavErJ3t7PcF+ptDLN3zhd8I+sj/t6
Sx+PKCO+v44ewKy4E2Oa1wCGjjsZfCcimu0Sw6mkS27qj5ItZxql8fktJoUNFOmPdc4MVbr17MjY
GwKoLakZQznKK2+Wy39yGeLXlDcAkr9tYvUotlJLakHj9bkFmeGjxyzDxdDOOm9HuNGQBNWvzeUB
Fpy5PCLTw+WwWTppjG+ta5f+KSPDH23f66pzVP8/Z/4qymgi7Z+Uf6M3m95eKJsWwWZm/J+enEOM
B8TqMAuw1g0zI0QX4LyllS/27bCKFPvBhoLeYgwUhuFlCtE0fOHGGZeCdJ0aDn0QONORuT7Wa4Xu
OCiEV4n+NMY4wXVmGyzq6YWTB13FPuCObn2GrLgiw2DpesD9q239KZyU93Von8tCv0wmGB/MvyuY
rlHR//RX37ORywdMOUCdZ2Tpq0wVtZmmPoLzuQsQIIXKB89eCJ//3AtOpN1PmhMKMqEupI/08Urw
FftJdSkg4wfywBLTgcHyl4y7RzRm34jdX6EeNZclDPkEu+Sx991CCr3W3I/IIdbSu85rb/DDfcpG
70moxRVYmKCrRfjeNtFWhYdOXzXSUnmqvUrenMPChgOwc+fZ9Pc3OxKgy1D5Gfg1g04i2YJlBS2Y
81dGSRZju9CPkZzhgufS0Gzk+lLtjOqkiYCJkthaS3qvw0T4wpBtaPzcQXetxfIow4CZ3w/jJ/JX
A4xF1odaTDSSQLzenwSuiLqdEW57YPEXRTJYHn+8qggjHeemUdJtKYR8/e4OQDE7MdM7S9Hqb7ZQ
P3EHmVKwr2QnAajRPJb+oum79RjKOuqcM9jZHUX5CA59KBi4sntzjx63+hfD0JK/6E7OjFgtopvb
UbQunRW8Ly4hLH6o8xUnXPIQSGOcU/NDV1HfB9VMNxAkxPA1aAqzevWIX0MgeKL/wBdEMUP+0Ju0
sQox7RpU1AaCWuTZLlqMVr3a6PEuLDG3XU4UKHjKVqH3tOQT8yDYA4RWxODcg9pU3rxp6L7PPeVD
fIu9fmMGvPgSRqjcMioJg+yJg34n03nt9+FHWgMC5kHAe+ZErlCh73yg+rpJYsruR+NNFE9L/FqS
Sh33aFpWY1Iokdg8FQzrKEiyU/NY3SNQbKggfUSmmSyQ5o94Lw3f7Vj71yLQ0srpanhCkjGDE+KR
skujI4kjefhXFab1CedOxVbvhIADNQxw/ROmKnMkKACJzsPxadpg0fys+idfBfLqCuL5LxHxHSCp
zOLTfYJdL3dlMVMCPiiY+1cPXdysPLhZ0w8d445WVSVeJeghsmMYYF/T8rFnU0fwdFM8DuFS8UVv
dij2XLIdMEG2NPXi0hJPsI8sZ2EakgqPqboZLWNiQif2cRLPasG58PjJg62gcL/Aq5N+EnRRuRuJ
WMJrFOXsDDHUb1TGHbSIliFQ8+0pvPFJ014yfPuv+6GNIcpHhqXtZAquGZLuz84rIes9GqVh0x1K
tHnGIsCEZJvT8mx1UdoOyLn5m02jq9E0NWS1SuiX7OEtgum2iKM861P3f2TKsj66U/K6PHExruBS
0ja9qMCQ2yJvV4UKYzGxREk3qyPbOS2+iUBxgvcJx2hYde05Zz+3uYjbGhIaZDc/r+x4NhVvd9ey
FQRoDmRtsVbC6hwbaiENSG/P0oOoxETVj735T5Whwjnee3yfkW6FyBs2J9k/VZ+Cxith3vQz5c3z
hT0saAQ8X+nVgNuA7zYxh/QwmthdbT3IZgi/BqT9KlgpVm1Vgplpd4m88GYvjViGh89YWKXQgxvF
6pW1IkhuqHEYnx2PtOdRfveLEs3j6+WdlS3jH8Sby0pGT25HvBB3ERskLS7lVIY+PaZA0UaD333+
HTA+qpONdp2+s3BxZjf67Q33Z8LWlb5TciaqV3m/FKXX1VVuMfHzvvs3dzU+ad43M4HTTyOEtztc
g/035nNiakwZ7IEcyAuPRmj/5ZTB31jK88eCIYaPZ2v8WFfqrEAc6OTRzcsLGjJkIwdmCuJRea+V
EapsHQcv3hl9SxAjcLkj03UcbtlQJ90bKN65fzCq7acdhKC+FkvUHKGcmaDbr8IJY1f3zFBxvfs0
HNxn0T8JO+OHlpyRzO0nhKVxCmO3lMxyQ4YCHie4rvRk3Rg39OLlE92rJCj0hqfG+lQhyoCj93dN
Y6WSbzFGATRtDrEhQ9hJ1bwi1TTuQjl54c7dY0EoUWH+wvIhGqnXgBFX//ual9GhHpT+4YzfTXYN
oZH2/kbc2uxenRsKTxX8qXM2P3cdBpj3kptpP0S5WACOQjIMAse6tsOcgd1lVi9HrTHHav5tpkGf
YIyR7MeBOHGy8mFNFyG/i67XKKxq/17F29nsaZ4KpKwji0YLZJiLUKKSOMiTzKbhiRtEbD9pEFWc
mNpAE7HSyxX1lGggWxmyqHp0H7DfaNJnvZKFfEMuDaWWHXuDYhHC36+iW4iot+OvaKkSF2BQpoTi
2ieUm43wBLRZu+sFBdP9eUZEZoeujPZee9GlAOokc6vLd7abaoKrY9jCceI7tdDE30NW4/YdGbNd
M1jBDLw46rgZ0ttuwQORXNKOWv+IRaAX8Qfc51c7wbPYpMtFipBBNe+lxoonKVttZ8EJjFAKWwtp
Fr+KJcxlpfptJFcM4Fneh9ogXBM6A+6UC5XRMSmrlQGGHFgKtmFXpzXEBfAE8flaik74aotTQicU
+PTZfieOFDPiPl+t8caUf9+eqgF07nOvJoL5+baV75g8LJPKtw+NZE/FjJHqUmWqdbt0s2stbF7K
YxQT6tLPq5rZbFA3YFBb6AV6i7sHqBt/Qa4Spt3TbC3KtOvbjDtzY5eiDygTxcxM6t58mmGkHbwA
WKKA+R+YZFaORyOjPKe8jMBqunOKB7xwn8OJ2MHzjAGLL6iVoEcyUZgD9TYO5buIPZTiRz3N4L1n
epCLzozH5qj5vkILl88M390bkQQcCZgFBYolID4LTADoqeoNdD/9kgpg7vjd9h5BbZF/8giHXdcR
3qfcZSJQagymfMTgwWm2BtTpECeXd/ExFiqcwP9Z+28KCCwahaiiNOV34ulqVs/xKDaM9mHVHLLk
npyMlCUdTmpojaYFUYs6oYcMWFlMI88Z9B7qHFgSbKuduMtC7QnJHQryU5iB7XCZQ9IzNAE6nZI0
vZeFVVKSoaVATUHyTZp4m87WbEDso7WZ0iRgyewcr5VeoaVcSfzFd3UUWJv6tSzNVNVoSpfYNbmD
yTaJP+R1sdsnAJXu+Az4ABUWY1YuQIJroKWn7U4htPVLWAgyueKc0+kGJUP21nuJbrJpNUcG9SVB
xDb16r98muqTrDyan85yl2mUqxHyZdV1e0vKvCQGA04WpcilQDbE9hUn/1d97hKottRetO5o7i4b
D4pV7XsK9eT8qu7HCzDLaSkopKPXSZO0monTV1o4BvVXLVSW9MDP4CA0QfjXRnVK4NoVM5E0nx5j
J6czewY4wqwRLux2NRtaHRYMjM4DYeYkbh5z9O+QELuCYkalYCt6eCiKLb3I8oJKlK58I9/Dkxx8
GBLZsEubUeEv0ZLju61BByhAxk/TQAXr9AWg0Ae4JqE9npbJ/W+Q9DYN071h25b2/o/g1Afg6OJ3
ZeQbXrG/2JV9mKWs+t1VAsvFN1Kn8zQz3q2Y/j8ZMjbyOWo5YtZ+KEr7CR8DiAmlpGXRA67XOXIi
jDUtIjWGPIv7tTcqXYwTSvlcfmaCAyjPkZLwAxLpmLfeUIQhAuWn/SuaBz4utWq0m+2KjDL/Gfvp
A80DlfO//yAjg5eQ54rQdOFh1fMHZm9vz9Uxq5QE/q+aVs6qKwhl30RgqjoSDEmwPtJGukn5VbOS
wepwZc1Pa2sJarYceh/QuVjSwNpnA5XkpwOgNQ/vqXPz8B0Mua45xtAyheoMS0gt9xYv/hpsWB58
5/lMYjRI6yGhYr1x5rCcXcLo40Q/cY/Uao+QGJO4HYz6lHcrMDLqt1ZdsH+Q9afB8J/OOMv29Q8G
HQhCxtUtVODv74g9xxeY8caC3ImVfM6eYTFmRC9tgVkP8ytPk+IP6k6Rstuk480bS2+4+HnMQ9ut
yz/jtlq/a7izuGVemHChfvB0d2wRnmEwafdrPVhag2GKs3uqr07HLxILYu41JBDyvo2zaCgXbIR6
q9zDnO1SYG6lWiQzjys2u/YNZxBw8mwjOg11if7EQJM9yFNfm0GkJi0t/aKV+JUYvwqM/LGP1gqL
xEO91u8S5WSyS3QfEA3+DfVD76KXywZWWyDy5kxNxVpSFdZoqGMigsw0NchXkvYgqdvsV8cii8vl
lPsEVdITInwHg7yfvCEuT5+UEZx1E2FiwyAgjueWnixPomSYnl//sj5CaV1Ikubmhne2n8XvoIze
cGFm0LLVul6Ll/LWlR6YpsmRuWegCMpLNgwzxyDt2FttxfgQEofEBELDSR48FI/lzQf9JTIu9zEW
GIA74N+yzBf6CF5dwej67eqaUFd9N9BAQ7OWBreV2GRZJz6a1/y3b0Qi8pgLPnMUq2YlWFPcxbSO
9uy5XhnXZbQ0gkw+sAhKtxMjRYXfAAN6tpn5IGcOIVR1eyRpUIcStyi9LAXj50y2EreMxgXDApH8
ULJfB6oNpdlpwI8Pbo0G5uh1JWKioMk0z1oTbMJ2FamURJwaaxosll7pNAjzOGn8d66PWd+UtaGn
Uu/RviPz1tBtMByMlGyqREb5Flzp09s+I5aMOOww8OilLldmO0cz77TGEsThh9KFFYxRdE66RzdF
O+F/xtHiFv/xL/ga6/5zzqK7EWHf8Dg734QzWxhTahrvmESBvgOeGMJiba0odNqf4jXPVtFGFJGS
pHwXOHflnEQopQLwnpC4TcAqimf9l7xdWAoe2eyCfIpDSFjIiFiCBzl1pLgqBm+tc++/VL0W4Ch9
BCube4dXbP3Md13eXSTEJIXbP2KnA+N7ZJRTtb1WsGhkW+lHT2XKGfv9yy1IEOa9t0czLta/tAfv
grSTOj/o/HbRvVRLQUkuvCOdwrd/Bgdw9mZUjMCO9ljuJ/IyaRBD23RnGi91H596Gdg5dIY55B9f
60axAZc0A7YmIJ4Y5Slu6f6JDD81kK9BVXJEYh5d7CPrcv4HrFgRjXr1j1XeJkMtTLoMyrlQbb5L
VX+WnUjDuivTkjQlXkbz4h1mPoeWTrv+njxcvDd5m1Bnd0P/frmo17OXPqSUFWxe8Af0qFbWP4IK
Vta64Cd6816doqPxLRXxwaFb7n38q1bCAHkfhBAs9E6nH3uCXIv04ect7HhxTBJukeJwlqZnlTzJ
KjeWTtGVEVI/OCPhnnG5brdrWj7LGx3p0b1xh2+Mf0jHvITul5fut51PsEqk6bxzIM42eHQ4+x0J
MFH0+0VN/GIGQCjVyivMbWrRAxVlqe2ukR3/oQOj/UHlaOf5ZpHE90I1xyOlDv5mgb8hhCvU2+AI
U1HFwQG5Aa9ioJJVoltdG03CHluRDjLuypw7n2dnIhOTFkmCO5TotHjVYjcANgparCR+eHYNAdQz
IqIAsoHfO8oKwLqLkDHHNZqz473IabzXCVtwcp5jSYK7u89cGTOX9qiwRkDmz0a5Q6hJ+iWJcdDE
4rB3lO44iOwYn5owTolXj7LHHXZX1gJT5LXIV/MaQ3Y3WngmrM1ptf58BvtJHJsaJ0XeDVvTsFPo
6Wg3x5TGvKqvurGubCONNcP2KyZxl06ELYm0bckDhZSUzVYMbjYyTrB6PrvPBbb22X/e2IWcqKee
BPLpUquhJ+noc5eidCaszUq1G1z8m/ut7QL3z7bqrcgLUlq315TQoUJQ39RwwebdEwryxVsxeySS
A6tLQV5PqSTUKGnCTyMajCJ4BF17BTD20QZWznCUv+8XuHvKQVvRH9ZWFjKLq7Yif/XovAgw5zD6
AuX8HNpVqJGjOwM7+8Olb2ja0oQzdvvtST4sOMxXWxn4+wKoj4AOXr/bJMJ0/YNaU6mC1QfmaejX
Tgt6jrZPP4z7YrC5B8G1pc5hsTTyt/2Q1kKj6zWM+BYmg/QosinCMsRjYCi9ZkStZ6V8z8yNcKVn
zOk4gBj+vA06U9muV6++mthvFSdDkVMusMb6+V/0iMjZLERDF8XQctj3lNI4jhyHvWsMgzwfJx8z
WRL8Zf9Kaiu1zQurJmRxVlSsv2CawMt1YpcpZKCclrQN+VvDGstkPZKTaH/FtDmFirsJ3XLIwdbv
rSVrezELoYD5OvhMFSpCfv8l+rXvPdrN0zpsNazZxAdgrwrkp9B1ByVRUcAMYhy0J17UU5tmAmIt
czZptIkSSNJD/9wU1WJ2wK+qBpLumhRaKap2r+VYlmVuO8Gtql5Hf3EsaMCFrB05kwdCuHSXU4B5
oYvEW5ZlWBd4jHA+HMDYIQge/pVmqw1Yypnww2a2sLQxFlm65UM1EcD0X03OTDR+k7iCnN2YOryk
blDB6SaBE+iLOHSLdAfOLafWZYTOJuJs5LIcs/ADYBVRgo22RaEWL9mRZrL1xFjBOwxAi7F7YmwU
8C8SjFQOzrcyiPbqgaCtj6YUZjXPTb4faysicM1jI0AzTtAKk6QJsR0XZ0TaRuOhZQnipocrbYPf
qh7JcWUS1MqR83e9HYkHb0iBKswP3d0Z7t/PNEd/vRbqEsfkpiA+NW108P7RFCeWKFX4Y3Rt5InQ
zs+Oz/1D1YWKwmsfPJaCmm6Ngs4vo6HvugtGuunDAU3K3r3/Qoh0cmjba7tUxrPD/VOiWnj9LtLw
xh/Mxq93maHoC3j4H0eriupjELwz7YUIiwkONTr90YVx/yeienqRmqgvZydrRP8ZB74wS2I6k+W3
2IIkSPIJIHyzPKwwPBRfqCSLIxDGPvaFqzxK+i5sax+KQGqHX8ccCpa/WpiGuZ/8TwzOGapd+SWP
WdUxVDSxTbjyRG5PaIHYdwZNGkpuMsj4mfOYHdDXp77Zd8dy9bSqpwip+GCuk94+k5XGFBQiaPXX
QTiIvmXAdsbGbgvExWQJlZxzdOYSgjcnLxu7kD1Pm7GA7D+d/1w0VWhoBNfUh9QA8yOvn7CHAEYS
DnTGbn05uf6cFEZ9v1O1Ow4ROoDjE+EfpNPYDjSk1Azck9VmiYhcyE8E1JCu7qJo8ZSTk0X0Hn4t
91MCMkZmTEyOaQDuTwRxylpev8o6nRP6unTRz8MmHRqrLF+3S7tVvJw313+s1qiM12UnUT/4FKMm
xMz6u9i/DVwyFq+Y8z/pNb3bKGO3EjohxHB+Mqx/x/1KS3rVs9MTUnuQ37Ovk8vMlPY/WUwJtcs/
iQ4LAsBePrLjDnEzv5NMNiONpdEXoaAfCjlHxjA8QvRVYPkMIm4oTHBswrUxb8e/37Q2GrJ8jcsV
3zY+ZmPrcMFVh6thQGmG8TSu7O4SQ4HQFJLECBEWsMVTO0xkwxdURSEq1ViTUSfhD5f1159Dewnd
y1qM9MWP4m6hFpPrdGXMci27JSGp/5lUo1Adc6qoAUNHjr0WwATpztSZ2ZJSNJsgM1yuh1F/H0rt
sR3U2K82eOwniVGxwcsRSzcTPnuQmnwgPwjhh6KPV9Jqo4cdQdcUfHm6YmSjX0S1MxqP0knNHqPe
VDzpaSMnIAxu/jOUCkI3/m0aJkALXO20yqDCVn7Y3ujByw0UbVxzu5FwnxKxO16SnIhAgstdfVC4
D3VMwZgqxs5ALvbdVFoUPvbnJvvNL2SRwU1F98z6LV8exsMg+rl1InwPrM/VyIsFTziLHq+Ewkdp
sFq5/kIFmEExzlX3mM07oI/RaaXxmt4Ndlndy/oZlOHlAnO4TKSSMoxhxiZEdtyT7SgWoVSF1MFP
J+W8TfooN8kyvDTIh9HJNNj5rNZUtd0pj4cpUXXy9FX2M/giDd27wPEaqxJyumGkEAPYYorLwgLM
f3oAakN8e9uMAYF7aXCy7L9YJYzqMULWvAAaKnjZqUQC3PaPIbkK40vK/nHvMK7yIiZ+QWAjhL4X
d4XxWJ6ic3VQfOWpRHsw4+FyQt1tWVNPoWgSBaTftPw0YxrrC9hTWNpsem556b3S59wgP+EEwPzp
pEQsivI9dh7P2AOnM97R+FaGbMiwk3VJEaaQR86uGmTMhYDc92AwNSgp1KAK8gpO43oXxBwpMBbZ
N64XzbKY+AYlpe3VrPASKNyiF7Kzg5+tENBC00IYN5oTnoy3C9hOd3R1gcybwSzZXsP8vCRuFMFU
xxG547R6mC7BYRrS0HJHqMjidJHmJMtTqbR6BDQ8sYrPqWo1Mbnl8igCqGhN58wv/8EpYu4mti2I
g5oYgl4nfQQbIQOyTRL3alv+GVAzlYckzvGiMTntuUotRiwtMO/Iu4zxsI8fLLQPAJZ6OeOQrw08
RtVeUK+iLok21l7QV+/46zSLVIRu20/o/r6vMfwbmGZh4rdM6hq/exAXxIy5HPDwHaglQKBN61aO
TbaSHNfebq9y0sERSwetYQ4Ym3ibLQqAGMhw9EDyCmb0c28jrCLuVn3VQ39L+ZewZOXbg+hwxUA6
V29NcbhTnVy8Mh4w1crsrhIkBJxqP1EWmFxgDyQbJdKv4uU/IJDLzDKHHNyQd69Drz8UmX6QlE51
ci5toUIvlClkgJwIH1/iaCVybTUbbe/tISB6OguPqAnFAF3qQFSmHah0WWZ+PQbNABOsb55TwiER
9XPxkxbz9tUmVph1HteN7PRepPTYJ7J103LZ6M44K9iAO4EL1BeAL552vvvD9ZWda96fVQrj0/ye
kHsZXwC+SMH3xxsOvu4EfboeuLGbDQb8qIGQwgj1tDlfYU0zVs9mrRzB3wOlrz4NEvjBcL1KI1CO
OC7udrNTYaRCEyzYbcmwKOt3MIX+XUgNkao0yy14mpKyg+kmdOzT+jE7eZdCRuQOuFeNkkAGPaz8
iOAwCRZ2zx2U/OVp1r6FtC8Q6DlOwJ8CdZ2VWjsVNjZu+/9av3r8Ys3t5WUbsOjHzvd9bO5aWTNy
i//Z5zm3FRNTARh3EiTUceWLwBkA1M4QXuUJERokXMXzm+a9hAhudmsY4czhSGeoMZluc6ShKX/z
5pd6X2OR9FRVaHZ9UV4N1v+oAX9nqkWtZPupAJsGGmWVS7oKrXTPKw7sSArvk3+B7my/ghk1wSmW
m72IKAxiP0RQxaZEOqubinpvFR4N7fiZKRtgrszApK36ZMzNllr93IywTa1bYFT4Fd4i5jGG1IdY
cv1VC7Bd8m/7fIT1xB+MfGGsRLJ6rtb+N9xYnZGDhKdZZnhuiVL/oIIIsSaBQeqtO0tyiLgnJoFO
Hekx0b0nW7H/Q2DuuL8zPto4vJauOAXmy0AVYJ9Ypwx6j3dRIS7ZWxnTJGzz1KZOzkyX+GP0qKRg
C7ohH5QbKwbPKc083XJ5kTUO9KYgqMWHEh/7NNcQARfk39VBmsg1HVlyqlioxceWMbzErCLiUBeR
7exabRcpBFiOg0MmGu4/FVxMf99XH40ubuKTeZ0Bup9/z7wPkabE1myKMMlpmjBQGEIaQhrOLCpo
9ed9KX1q1k8bgUElyde9ChxZ2uMAWhYzm5MRV9cCqgf9vCxQtSR71YI/Zg+1LW/P4k090pSkUnRy
dlM2uT95YoqBxBPar3eyfGFOvT5grYvETux10n+rmSutR1xivQDLSU4PUN2CZIdsyLFsBZIPk1df
uATs+vLJn2rVTN4RHQirs93W0CLGYSw18bvIeAMNrAcFWJMsXORmEpK8TdOdw1NtrDSHqLQAF/dA
ObFgv3DLA/h8vNgF9B+KiDf9PSwtcT3RovC4gyzO2lsTPeNI6yepsMx7GgzAz4H8jomrBLuc59DB
arPPDobsuPLRZ3hXiSN6xv0/dNC16kFnNyBseoaz3UcWebY1fEH0ep+wGqrfHjL3dgIxJRrYgg2e
h4k9YEzvJ5P1N7v3LV+ai8WwvmVA6Fl2PyNjl7ERZE0/nyCTg6ogz7wuu4qxpyMbh6v2eJN1CO1O
qBdVFBWXxA/PcKhLBIqNKiSrNn2S0HADpxcNcGtuHwOdhWmwo6Ix60Y/0aAPWRXwSo9Sj7X3ZYez
M3RAeaWzPMpeN4Ih6YmeUKa2F0m7vF/X4D3G8+5Yu8vuRFRI6UDiM/VcLCEuC8RxQlBEmVvU/k9s
P0RdkTwNxz6nJedPGt2etIllOyIIKddRsBm43epJQFI7FwhyBlA3/mECx77Nxqeb4Xg53q4P3Cbd
dx5M7oFwTsXqf4CCVj/mGmHTfVpY7vXFYAzHCNKfstvN6pwR4yAj9ztr/iOpc2KOE5EQ0WKVivFr
21ndqYir4/tXkan4yLSbkVmt/Aai/5z+c8TzCMLANIpQP681aIhuog/qw6Ma8Jk4Hr1KtSgmJRb4
ICrJj6Z6ZTTIDB3wkY1j/xZlXZfz5gxsyLA5GalsfV8qYw7MC5b9lLUaa2Ni/PXrl7+9lpVrETsS
16mrH8bZuwjOpry8SMZ0I0iGnrAgWShA+p0IiKs2cENoCK0l5hVd3xJ4/XtdwQ8OzXyKl29Y1qWL
vX2M7SUT12FZwNnN3e2IkPHuXC5B1LQ2Httx0GLwXVLx/7xmS4gvwAhsG1pYeSSoVHPJgjOvIruE
etyOgQuKky0l/sJsvf58t59tFHP/MLXfGJwIn9pCrDxkHovPRT3m6ajdOHnpYxG5Hsf1gagVFaAV
+cuLtNJdilXGS145nsGH3LXOcyIN/BczKe+KV3hH84PSFo8CiXW44gH+I5VcVLlODId9AiKwL8HU
Qi/E938DrxzlgU5mH+r4Vq7S7CFGrdNKYPolpZ0QeIyX93Tt8W763TORMxqlK1KU7cSnX857UbHq
p9gzh4SPNxcswaYVYzOYIjMonAYvKgxwmFh7GM63REaN4cZK9j4WPHRJqfEYtOqj7xb2PMGmwOsP
KMZtKW9ZhvFJbrsiU1VrnpeTSVa4TCDp2UEV5QAD+0sUaai4Syz7ndt7jVFfQNtooGtVIu1vPyq/
i6KqPHcIQeu7BfbEEP5bHW3dRldN+S85TaBHgvJW403do4H1FkWpBopEiEuukFDRrfPlXA1Nhpgm
3w/dL3+6YDbRTg9+yqLeffqXWiXXVHtw+dzn/oMtB8B5EicIHzoDJAeGYNoF9N59hDqqT1ygfnLB
m8JjKyYPtnzwMPd+W7nCZrUbU15qhOD8gmHmLZdAA04/NrSkQ8jBa1PYUkI79shME63nIyQY94s8
Ux7aCnUeOj4/L7VDa9J231ttiW0ZcMinhW35Ky6EnrriGsP938Ev79JOerGiIE4IfYhy8Hc0e6ih
Mem9HARa8kl4xPJq8C39e3m+qLTLddxTmyHSd2lbCr/Ovbl4UkMTDwjyrWSEJ917qc7ygCHCad2c
SBCALY2ipaXcvhtm/b9ZrVmztpYoAgi01Zj/IK2kWlsHRn4twYCUNY34zwc0QaJVL+zSGesqPmg+
Tyg83Thko5KS4MlAHbBAKHb+GpeVn8Te/U7/R/vhDas6rhtfJDMqLEoWk3e2Y+qEhLm1o4+KP29R
6T17N4R5iiEK5PRHWr/YuwWywUMU2RGcaMf2NA2UkwFLHK4Jp9gUwYcNAaNQ42OWzowp/LcmuknA
8kqxFz2rciXXhQnpGCtIW2KZbuCg7BVErEbTPcfd1gkxlaetqZXI9lW8FUEyt72kHC3cvNseO536
IKGXmtHlCmw9d177dCh6YLi2Z8ypRjqGDXQAj9bFVgB3GXzkPaMXo7M0jdtVVrf3qx17HcLaRp3P
VDt9wu04NHAjBqU8VhETuNg0BCsFSVzyimJlfzS3Dym3FRdWG1/uVoue5DR9Ls9386vlDLyCZJnG
Fm+Qt2iCH8NPhcJy2EF0S1qYeDGfn0qQJa8rt38QcRVKptOjzT88qnHKKTDFB5pWLpeIk8MoDX9L
eXwqILjmf6dEzZV5MnNXAknqwSV4uz6tYoyI9TJRF/+RhyU5YdIRoE1mGO0qhCwlpzu5nP0GXjZE
NmGBoAOno2V0oxrMaNpLvi7PnpSGyakmH7xJFFbxQj6GFvFnTDwcV6bAb5+zrn3AcZGlSJo4cVwF
11oqDqDH0FLdt8dqKvyXLd9wRv7xStMO+F5WEuPCSTzeRK+uzoQjwVHk3UIi/0ZfDlJAwPZa4iB4
Ilp5aYI+UWqCkWXLlcwO8dLAtGQpYvJeAkFJlDlxew+7pv/dRa2BJMJL6H8gGMmozKITftDhE5Gz
ho9Gbnj7cxElJnceVeQwJG5vK7DiDE+gkEPNvS7o/WRZHFSj8Ot1VW5VGJ1lsNHb9R7ADEqHFK5j
caPLhpAmLS2avw4rlu9v+zTUXph8FVgsIElW8OWimRpVGQP+E036qwXLC+YEHUnkQrBadTxQxa9+
g4/dYYvzrjAXkXOdNrYturuAkdfLQbjJwKhSwcUDIDyDgIe4A4Rqe1gU527AGaXqswquGKUaPkGa
Rmvwu6zBAluh6ZHQ5WEZO3l985AvXbinGyhBe5jUZYFxcNyteOCkLr82644c3n5b4pP8m2i5qYUo
61VDAOaSJ4bzqN0q+k22VPH8mmsm4cWODzp7acEKLEULLbeDLtwSAXe0koBruwwz5jh5YDfRkmGx
fuqit9Cd3nbE4hBVXTjWyCwiLUlC3f+92VJFP6MbjJxl9WCJuFM0KPiAffOkDffl5AVIBmuUcaXl
mTqCxhNQrvCHWGX0EoypmNSr0LA65VAoFBl1CDG4IDtp9WRz1d04EsDxiNMBra53fs0S7QJXHhLs
myg3BPKuTvhCQ5cB3KVzBNRbL8mNFUfAzXO8XLzvEZtNEfUD8U7Ir9fYISuPMSvTdX2fCvwa1+1h
Kf2PNyL2PNbm77mVgXO/jKIYNRz1QLKtGr4k+u/fJsAg1isGKrWrNvWatB6s8tj60X9NH6QY0c2Q
VfOAcuP85GCQbzxiPmyTSkRgZJROKjrDJhaHXaboO6W8zHkCYIISdKdPGY7OlwZIryR2z+8XPUvT
Vr2Sp9gDAs/nB+Vgec0tAQ/OSkqKOUGcqPRsUiShZHHho+1G1kkxxXK+zMkKfKpzfCPS+8lL3W4R
ky918gyYNYa4UpYj0SfJPUNfLqdjc/YmK3VpfKnZnQOiRYQDBawDqRTkdHZ17o5BSJNYlj9XVf2/
LblKBtCmu6foZEFTraL6BX9IgCeybymqdjZPna4p/GHQvkOvun0uaB/fvV5sGhOEvyQ3RhnpB3go
fOeHTcfAfdg82Jpnc8/q24Jjj5Qlhk1ikEZC/d3jlGSwcW7jviPs2f/UYf1CVypyblG6oAeTbneR
hgQPCPJHLYiVM0oj6s29cbsXuypdkLoj9+cVJEtbkSq239P38+oPCE0BnOa9kPvxB5RifiVxAVUy
UiQsUQcNBNtD1TxNprMw1iZcHGUBLUSD8RMPLCPmcz1Bh6FGgX9NwrvJ/wUlsQBZ0qDrqVj/k3OS
AonZsA6rXS06bKRxu3ypf6/T6DMW9HfYuQ7z3hy03b/QQYWUCZ3W4imk9bxibZ/Lp5kWRN8ex/9o
1H8L3COF2YrUbfnf60PCfO3NoSyMXPa97nWDdH8PPZeVrUewS//NFIGWV9qOUqQLMrteLNFOcEnh
S2d5HLsQ1fni622lIzMqGyxqpXBJBaALIqXcMqK2uLDmSvQXRwJQZv0gFu1Y8xByC4oX1mzOjz0R
D53sHOB0cA0B4uP+SO046DHK4h/7suId85LJOChzlmWqhmlgu7ozBMIhrF3NraTM/PoOETO3b6Hs
tFdt4Y3+HIcevsSbql/ezcURh0xyQljs282HuunJGuN224ImOmtpEDyG/rULPHOE8gvH82AcoAqb
hIn+cXhGT8iSUeXcICp4Y1odSJysh223GWCp7qbqZIEhU0lpnZX1HHyDZ8ZOvlWOEzHs95BBs1ki
Ax3cog8q1dlNNfLW/zW/ki01/4Jc2xN10UtmrU7hVJGtOmhHNVd0cCaOCvWrgTDmqwiinKCddEf0
Hna8au36s3yeqH7ijfMY5DGnXDYkhN8ggMctgPkZPMHhMRD8D8HWKPrxcoYTlLX+IyIQs1VbZ/Ma
/A/HjijqGxNqBRtUgAiJFHVPMZn4DsbLYtxgOHXIz+PG0MYDSTpFgQ+CJ4aeIbf9VwKqE3/7DZDL
seFDJeigco4aQgQSIGAqknRYUyh1wmn4juYII/p2uc3J58EOGj/NGkdI+H/0gI+P0DLKZTjClEiy
CgwuJ8vVzNfqmyTkfdmmimWKySGj5SqyvzGsOJS/B8ZT7EFvPk3U0oHbqcFgOpCbtF53wOCDQN9J
lnaE3uHdXnoIDsmAE9MC5fX0tY0FCncOUA0PnDFgwXsPbQepMuSAR3SRXSN05dmRq9zLj89YUVeN
NftqIB5dTYptxO1TkgghfpudRQi8OJMDf9PKsdzuiDcrV229rSOtlqaS6jvqo1yYYGgk2FLwfTB4
L0ThhgHsiTv8wI4APYI1JYnz6PIM3/qcKbUX92Xlw1c5xSJFSHaakZDf4TLKoIAISrcXUE93nt33
83TpRWmdRtYT5WczyrMRRsSzjKAOA0dbHYE/KNDiEOtuKpLGrvdb0YDzamjVIHHmtpDsWfzdXAcu
sVZOmvIcPDuEcQiwP3bzNpqWSdVUvcGHNYNuF0LAxR7Y9pigkhjmALvsnPJtgJRyQEtMR5PXvrMD
WcEGYlccdoQnIaauau1/DJ9ohhqMOaSCGgqOvsy4pW3oTThNnOTDHJyaTHllbWauTPbK7lqXmoK0
+KHB0SoEPXYFcjVuPGZqR2SSUR/dGPAn3FGuv/9U01mvrY29ORZPF/Vjx2VIEdYeL04PCxTuCGu7
N8z/2JRoDMj9n2k8bUnzUjtvqosoCNGDAAXJuSGD3/I1FTF+7xcwqThfqX0SjLNW/KYFONn1nDdE
tZyae0oqECNj6n8bmYQf4OlZzcw6OdzvY5f48YYK7CcQ5C4gNPCW241sNQj2R67NnbQjOBTD7NUy
+azypNntpHP55EMdY/31UEhVPZZp+f0iDlHiZ6c5oFs64DAY/xlqSBvUFD16JasvwlGuiOUNNcZF
2Z4jFODMhg1NtmMhhQhlOxqwnGAQFg1jRGk5WRrIEVurMUTPk9JyFE5YpoOTQO+sWvSaOK566l7e
M/u0bwf3M7qhxGFY3ybdkvhbc305kqEgHUHrNofVWAKzmkIcxAQTJkkZ730fHJMDFLobewR/z19O
RL3c03fSI2MfGwN+lV/Yd/7nRcjYMl3wNr0BPrhBvHgBTu44MthPdCzFRDVPuRaH/Un4550/O3CQ
LwFjaO0/UtQAMYg4JE9ZtzamjF4424itT6vSqsbx8FberUWEcZmPJDRrp5UZZIe0unle3kHPjRAz
xL0V5XlH/W3ccwhfaIgEMbgingfJGAGOyW2B+GVO2oIUK1mHNhe3IQUanopElne2KtqwbRIZZF5l
5D4mRs+XjyCkIz0QNXX9yevo3F/SKhrx1U1P6YtlPW6J7e/7vfsoow2SMzoKzi8J6vpIlOyE6jZj
hznzC7ogh4TNIvPcn1DWc7iStlu8hsXoAR6F8Rm0fXtkieGNw8hMVdDbPp/+1waF+I7zQp1cYkJZ
7wMjUa7XdG5zgroLYPF0Ywkpt6gV+RLZWC9vOQNEQQjfNVRr32B2y56AOjIKXUGByVex4lqGgkwV
tqYcxothBPXs/pr2WR4iDN6eZl/S1L9WuAJvcH1f2JL27T7OCn701U2owKhDso72IPYLbv5EuMBX
bm+1EtVYdPYCPHnfwjsuV+ckFKrWHemzqXMZJxWQJVb49kPEw5z9hGvmkkMdVQ7N0L9Pm+j38CIo
7/TTiXCV2jfh05EiWzvE/jZNwFi1nC/TfNi+frfxpWysbicErbq0BWCzPTRp3twImgyVqou8gmE0
xKQ1z/F7WgFF5Kl9ikYBEjfr/BQhVSxxu0Jav625ivGNcJEdLWdYLnHXCAkQOLGkyNR+oGqNieR4
ZVBb2qm6SuY+q0dnA8XuvUN8rHtPoBnlnVEHP3uyU47yhv7RvfAD/mHx5qRTPpWkB+mL0KWeE1iH
JvoBD0RCki1CAL+5lE3SeI66z+zqolSXbLtpeAlDwmJeG6cTqEfW+xtCGCEC5WWGyVAspuK5AffY
er6YyMq47dqzT82CEKxl6cSArTvaEcyK7KjWqEoHWHsfJ4ySON+FfbLREaT5jkNN/T9PJJTa+CuG
qXQBO2awE+7B8NWHzHn411ts6IUVf0zQUTfXe3EQaxQX7mWQAi5SR0pTCGzukwm3rG+HQ7RbBNYo
ffOqFu9muFAWtFklz0HOVXANQKWTG1CuLz8OgGuOKu7uxC9cyQNBdHOUuJZcXYwo6laYbSqujL1q
xWaLymlmLNWMR0q4SNYP+p1imsIbzSPUfx6UY3E0nGBLBmpXygk0g1Tf6zuNv7T7eOgx/oDuqnhR
Y7cGRCAFGE3assHPeouvyP4kLDgido4dZ/cSEF9kadXAd6oF521fOcIeKTHXjexPJVjZW+2yg697
EGHOjqZsDx2gERTwabj/mEn0Q7gVZxd6RPqOzxiR+HDivQvWBdodiW2Uumgce4hBOk/13icweAg+
H+nAI/NwtvPF67VbKH36N1yBUu3Sc6YcyMFLNYDjY2cDsMEp3lh0j1Kqx7MYhVHWDfgIDY20gsI2
24t7wvFGeZIclLY7D9iyUJTRzqKlM7cw8OQAie/oKpCm29F4tIptzh853lxa3YXp46zcghgMfZ/c
qB6j1eqpN9x4/casDr9DN7Y7vhUo22iT4HWNOHFrhQkwfUodp6s/eOrZb2fN6sSa3QS5h3OcYSJd
twAynC2+mfP/7e6A/nflbh5xPoibfA2lZ7SjF9/rMjO5BiXsMTborjAUrOI8SLbSgZyiudQgIPho
TZvcsvKioh7M8313I2JyB76UMUor8cX2XNT5q2Oey0zEZ6lk5MJtrMq+wYEehs+jVeDH5bqSwPvL
OFcTFqyPmC8GoG945Kg8Z4XHRT2ax4IXuhIiLKZDE8wDFKbu732nG63qz5JxRhmTUPUdYDPwgRm7
wWxRdRCg0phQbgZn/3gvBEl/0LeKB4XDxWmgJ1FqY6zQagu8LpTMya0f+NQ4NNQXvus2Q7C+xf/v
yoc4RwCl3v+wHG2aFROs+uI54knLKshEsONJ+mwNii7eGyCN2KSna9uo1M8eYpmWhfQLbOmG40Bl
x0ITj0XHk3uIL0KEnLAELes7rkFZrnfZkomPrwHQN5Uxd/fM7o6pDgOCPszW5DNXnaW7bu0I1GDY
axYm5AMZZImL4QNo/VBnjydCTGKPhVqPjI2++Guw2ttplp4OfQcB5nZAGs//Rs81c5vneWfu1+Yx
RptNohUbaPA59pDNlYX2Y3H01Y189qyM/GNc6r7nsR6PeuUa9sVcc/YZfMl4oWC6pxQ0GI0cqbJ6
G0gFFazZuy7zFcnw38pAMwIao0brA8IFnHNhPpz12gGJk3OwJi4l6km7ygrC4mhlCaLT+EzWuNKv
JuVGn82y3Cu37cX2JUP0fWoTy9hfknE+EkiaYPsUKuSpjHG8LXNljz77cu5/QBOC1FVMBOqkV8Gp
2VNS9bQyswtmJyCzsQYKAhByx0pa2Yb1+sZiGlvZyMAk4jPz3pgD5ky7BC5ruDKY6UGoouhC+gsG
kOVKAJuL8EiH4LHwkV1SszoWL/CuRL8s3Dt9jOhJhhK28r5n16S2mgNHpuGE4jWYS75gLONpGw5v
A26b461xMELxMTCbft3rZJMlgw/JBZ3l5Gga7jlF3nOVtQqGwuoyI02ao3DLbK+itkBC1Xq2p4Fc
Oksj8bRb0ZuXavqkO6W6iEAZ1yvf7+A5nmE9TbUilVgXTjqlXonqt/4SGMdB/C3al44vcLs4C1jH
/XnR6ahWxp5GHQ45TPuVCwI9pPAqHf787mxSy3BIQIx0WOIpewJn8Polfl4PnFpK6mrYtlICGRZI
ZDSEgwT9f4TNrY9vllEk/q9HK2ztFtc6v+Dl9q6WPEJqfUfyuAL5nAEM7MQtcgslr41tRm+MifOg
uyVuhenqZoBvwJd3PV7H0syPy6FRAfjeYgYHfQYDpTG3xjY7k0hDBr7asAwXC7Ps7qXCj1N8Rej4
3YJM7Bj7QjHf+2PO/+KHZBmWOg9+HgNH5gQ0hYH7ernlVAA4PdpfWQmZ2qE7BrdcVGN/BEP25kaC
iWGzf3U5amL1y08LRMkoc8v82gXkNTCeCXHbt/dUtfNCOM1VA7D46MhSPBQK7daNU4uXqd5itfNN
ScyeUCb8DkVbcUWqfqcNqP5gMNP/Mn9Tkkbjj0mxk+x50CiujEzlVxIB+ycjIoIuHgWjD5UJDmMN
sBBXnFy1SK8gWBRlT81p/1pR8hKKuUxleudEBZxeQ8v/OKVWFbNHrlbA5PIfhr/4+/H51FPEqk7T
CNKYrN9H+8Z2ICuzV8flCww/05gG4p2/VoRQHM+rQadSexsJG/ldp+Nw3tHRfhQmmk12rjIKGW67
ClE154VYEl3KYMYr0IFOApa0K8i3pxTg1/WaQ3g1O50fTdx4u64ovC6ujodNqTu0fImcB4SAOVh9
t2kYhkogzOZ9mD544sPjIltrjKYnE42CzedWnTAewGI0/iunv/6tCzLzB+NCZcwPYTURc7o8T8oG
WYVAzjTm6FB4Y7UzSKUeDQDFylRvCKRS6pk4lI9iUhqWOFwd+lN5Vawm8Aq9TGejEOWK/tbblBbL
YnbuFQyjlg5xVamfUxeor9zUKdiJvBeiT/1vxdYNxvecgljXbTgSaukq6nFc6ZOPo8nGGcqB/5hJ
yjGgWMdhedKoKkwSKhvJdoTJE++1hG10QkS7ZPdReFn62V8fTS10rOJwSqCez1Y4hj5KZXDGlOqX
cGxaHoYAHxXGkN+YJ31tRvBo40AFEsKuQ+d71SkycZG2w/ewJT1ZYaRw7aGfJOj9t79xkFweuK8L
wlcWkhS1F/FlA5BVi+hzGbxuY92CakZjE3s5v/H0gUYS1D7WowA+i+gwBhHJJg+c76cy6cdJGQQC
8cKqyl3nWXapYJA/0C8FVKzDHFNyCmeRze3/JQ+Etnv+Xxgq0p6Y5pScMa7DNqM+InuSIAUrOnJz
l6TuAW1aLPo8m+r83RNogkMGISwl5rIUvKMnuDH3CyAElXrm+CInFMVlELRwc4O3TUvCkuob3v4k
d7CsegDfzyOEMiu3n8Dp5eXgsrMCr2dEPCe0xTOGZKV2oAa+BKbxBqNtvosJRI9av5WUTdLuJqr3
JcfYFnNbxaM82TsUXUJUqxJWPDjuZCg4dR5kgq4QbmvW05a6/xfzUE1ZEGG3+UXUnkLHwUMWJnrA
PiEY8OsaNngq103GkxyI7TZqT58+7cClz9aj6uhG34ORXFLOTKA7s2MsyIXBtDZl6FcPPwseqE2T
b9mz2OnDN7w4bSlqQfqliL1EnIHuTKjpuTN5M9+22xqq7m+/u2AElO/hi72jBZtYdL3RZbwm8mKy
gmdnqLqqVPs9LJADnLNUI6vDfRDUhZ5aogV3/iiPoU21ttIpHGFeribi3ISPStlmuMIiyVPwuPSk
bgbkTQcyw3fyF+6iyv3a2/q2qeDXM9XdlvmudQEB0VdnGOR0nrvkF8deRKVppNqCRfPeEgyXNBrQ
FBzSd5QoiT9pw30MXReA8tvQDxiQROMSnHgRqlIJXulyq16qc04u0K1prFlcBWqt8S3s/PXjHmpa
h6pe4c24x4VJQUtRFXCQo3bB1h/d9o9fRvj66kSg7SwRp+EbU7veM4H+sWMsT6ow4WA7HpzJJHgr
RP8P4K7hkn+GRODNQ5R13cPRpcCPq4oFErtVjj/bvO90iFbdnxK1+irT5DMfqzGolyjC6Rhl72BY
Z/wmXq9iEeDLeH46ztGP0lZZQtTWJrRAPhLlF/ERG+jQYm0CpzwJ5BU4bkOVMN+k3P1m3xbv7Mt5
MFNSYiiN+AhDlfSCy4+m+2EEAegqzGVZFaRLzJMbvYsuzB+ixyWuY1r2JT4HoOdWwyp6xyWueje6
9kG1LwWiQ5OkKd32RKdsQaSPrv0MNjQJGpze1ednIxPhS3xtsZPME0QxiMaciw7sBknO28q9NKKf
3eTKjXddovMoNgMzIiiAV9fbB3oMsG0rEBB2wJCvaBhjERpwRYl9fABKWzzafsT47woubPAuS0Xs
m3UgDSijOvUcc8OCMxvm5En7lLpOAhL2dVpRRYj9fGSRM5Lmok3ZQDQqGWwroEIY+2AMj55ijjoe
5uoJbM31CSlXp8jdlCpZjDKhsmkzmKZWqYIP9TYS5EPRCrOGhGe9Thcw/6Ss45pqz/9CaUnVdlQ0
cLU7GHvxIdi0YdQdGmSMP/EYLxIcJ2v1rHX2J+9t+l6K9ZEKcev9jihq29lg+edHkpRmbxshmNY8
us+YllOum0KQUuleTmUVkZyP17dwmzRzT4CiiAQy4Rp6/7fGms/GRP34hMoTA9kMwjptT5IL4dGS
OAQVDlXvs9w/DGL9OqRAc2CQAXVp5nG/4wgu//yDOivSo9WrGDcLgu9uUmSc3pKIdcaf/huAF6i8
6jVyHsFnWto1BETPI/UcS0Tls0t8XA5Bsz3F8PvowGqwxUj/sCf9J8qzSPa3jRl3P2kO396TiykO
MPpfSXf4JSacwuBZ+9s8CKquCDpW+Egsi9kootTUb9WH2E6KuoPWl3y2qj8Yi8bMgEMGX8YGXouI
lL2oeI7e8Wh3jsKps//IGKTrEhp8okymID3rP1EYqlU0qt+E4EQfdaTW7U83z+2acJBparBO1HE8
ATmyQWY46Hgu7/aWttKuj5L5pgMloE7Zw3f4XMyovsSWvp5q20vz5lbImn1d3tSW/Z0vq6QdXxUM
2tVq1FWo9oRcyHejL969iFsOYwc+LpkpgjcXuKsDB74tXWAQyFnY3MR/n1iMgkIAjmHwuyGt3GsY
ugB/49+JHAkN8NcfpNB4+qup2XnQz2zkKDmm0+duusat7Sn6F5a3QAz9/bmAuebyOV85supbCi6B
NofveO+q2AHfASRLqCjuhl0LlzchVcdM6Jz+vWXvkM03GbnD62RZcZA5YxUhmld3o0W0KLJhQO5C
9CNJ/gmtSx0Xox8zSE8O664cvQZRq0haIKsLD+kzqSayVAysdjL43I/FtDaNxAs2W5zwp04H1DFv
i21cFrkKEJagpPXUEI2QCwvqvsliH68FNNJj8jQTaDQTS0vzOQOj2pGDG99TdkJS9D2CkjGDVy0l
rdl9+6gyLFTSEFw7RC6ts/8iy5CGfSJclbRxt1EFGIAyUxA/DqYNp+Iqw7Zbpu6cha0t8/D44Idm
Kc7xkHsjU1XD+FoYQRs48AG4kxo+QLpPRfcXcBDG/9SrTB/cKi1KmayF4urhsI6mvjmI7ryhDNKI
oyn48uvj97v++a3fHRp2Ng+dDe7Pt1S3DzIRTjkU1WzdSP44mDe9WpsooKOsHxqgjR+IFN1Mt1vz
tsoFpCaoKDvHI6YujRZ2zxPkVaXgQaBmsCBJHfqHPdrwDpkoqVzdurXwEoY8bEh0Pyhjc6tcwhEx
DRuFS2vkJF+c3r0ZIx219a/RzuXkWKtaMwvU9cRawwAPjXRHh/W7DKhdM4G7dbKtLZsJ8D2yhfJC
kzCWh/uKI8QRyHgBjncqRUPgqsoqFTNCT/EXjM9RaZ6lSuPgkR9leJ7KRV0M6Xmtg1yO9a41/vgE
AhPIueTTgC2nXp5Y8Az+4hP+L3i+eEpPfKPHBJIJl7k1nP7evDl4dw9OdIHNeavpQDOtG/ZtEYLT
n2nKNRw9RnLHp7PWxxYbtkQ2SnEFgF6xlKhm/Nx3HK5se69W/J5aOIE3N0pSbkYEDkozDg/tSIEh
BpuzIxfkxI/j4XySF6afNEzm5rkLpVFPkHGF6pjUXNAKDOaoYArh3AnokxHRhmX6JRnFG6vb3kME
4eItkqWhFlCjcQb3WJNsQPUD3eBj4UMxSZLeV7sIbbkVdHuUgwb1luU2BsrZQaKRNDVAPfORSFLC
6hHwDUku6LETO+2GyoSWRB8lJsuIe08V4gGR66pB/tHaufFUY31U1uD3GgDSukTFb/t04Yip+xhS
5OxUL6OUn74FsjV4IWts7VwSpKjQUF39NDYxD+PN5hc+SNnOqbiv0dWrgZqI0T+JQGadKqAqiClr
OWeuHYdYE8SaSjNvZbhK+lxVeqdSg52y3LADfbeezMsFd+k4X9ZPJ4C3bbGfxqfSkNaX8iGLgZ2U
6xRp/5i255xXyDn95n8XsbHA33Ro3VgywlDqPOU7D6LYH4hVr9c2AKuq0IXsDsg09d37mORBA8JK
vZLiKDyWpRFTnWbv2RnlCbMZiauL6+xQs53chulzEPz0UR6naCvmzBqT2GCe0wibAsMFuzUR3Rc7
gkX5JG0sxEujtZSwH/u1JAzOm6nYjrzQU8v1R1RIblKhxtnpsid9Q5szlefjOiScm7igv5xdTw/r
Isa7O4ggD25NSbiVd+WlO2S83HZ84jqIUnEiFF1lhv61P8hypXO+3dE1BZnq10S4NBL+g8hgZLTy
y2dHh0P5TxlzMS7jSWrF19tCXl9C5G+51h7mcjIHcYW3jNOp0eszwJx/sfAsqOLQDhnkbUq2opK/
cbOwaJ0feEC+K3GIKzBamPvrwFkylFkXCFSjnIdpd4SrMF9fRc8G4lGvKkBCUdv8ZLxs/sOg/OF8
nlXNqnePBvUAWUF/fLADsxoiJBaGU8a7iXianXiPHZalNJ5iefcwhIVveC+VSw1I54Vsyr0ucpKj
hB/+xQACg/JPG9UgG+/QSoe5YDtBdD7lgrGEkzbWKZqHy22PVJ6zXMRIeuhPNq4yDn0goOJ9J2qc
FvRtSBqgRcLtjlZXrTJN+aMXQCEchYzfHMCoJEMMhMJQYP0Ih9wkH619kkHlFx/e+hx5VMHCGY6+
5xR3ChmBFH4Z21+Zcobt7hQdL5Cp+GgjX6VabdPfedyYrIUHUqelHTpNWq0n+RIQ1qM2dJ0CspAM
mrBTJCIMi0Vqeh5gVKpRMh5yBUvOuQRwCnk4+vrL09CIoTH8/Ztr77o5r/9JZe6d/yXKuoK8WFUM
yUh1M2aVVgtu5NkRqxE3oH/hPN3wwOmqW6aaVn6Ac7eWp4IiBuvBrH5UEoxBTYIBLRIA1FgVeHhY
Zp9o8Lx+xbzbN4Fzkkcyi6XnqmolqAmBA1MOtEyluWqNRab8gQUtRE1UHC42qrRK0Vk4GFHC5xUG
TR84ufltOrBixx5Mo1LjSdEbyEss943tmdJ7JQE8jH43jY9d4d9hqivAarTYE408nkj2HDGVYosv
KjwghN9oczpxMlxnWy3NJ6H8Pg0GlQUFFIdifLqbdNjzF6xjT00YmIccl2SLIzABdjhKRQGZbBjv
u8rblJ7nnQYqH6MdiKLg+Nycl6dmLa+mI+AGutB8piijMgNskz0feqkkP3ShoDFr4PaI/RN/9ChA
Sya1PfdbXviOqhO8pmqYuOIL+wAbJK4hB3GuuR3wB3EEPye6BWGI7M65grtFeUmneRDnAtk6taVQ
GT94afl4hIbaOgcSkHM4NJ/wfKOiqHm9X9isef9B2PKwgL0nVhU1U3U1GY1tWf7TrIGigiYTCjgt
BCR+qPW2+0t17oO5X60zLgBWYbPx6mW035kM12H2so5Vj3Zm4sFsNHMVJbjwOPZDOm1QXn7kbgJ9
4wlsihMqFZeVLrXuBej0e3LNzZPfhaVh+SG/4HBduJNc8o2RQAv1ogWx3HTxfVtBiL+tfQbr/5km
T3dD67PqoI2B2NDfc1LVx8WTsMT4EAd17hqMaKYzxniNQD24G77GdbCyui2NMHkNfibSadtX4Kkv
Azf+RP1SdRpU1aSiHGxYyLhh+CmhHA8Nbtup76vQPJ8gunyNDQphXaLbBkg5I0R+lRFTOu5hAVnQ
VqP/iPao5/l4ykaTkinMojecZjPZIt9I1E3opydnN2n3SVXQ463x6UhBQc5rJjEuCho86IfFBZh0
G24sY1Op9jKhOSmgeWYGHKz07b0KpyKYowS/OO7maaeoK4AENfVZbbco42YxLhfOe+ITNhiyt+yw
8vA/DBgITLCyjYlu1mgE0jU46vJQht/K6CFIyaGgWuIc020vil64rJDL+emIwTHv9TH9tA2CTVvG
rKP7JgOlj3MRVQQEN79xjiEWkcrtWBhWiLOw+nBY9Cw8rGQ1dWevVO3i4W6LsfdSq0bGKcg2AhrQ
DnU+pA4LeJC83MLUVEa+8TTLCCVRJRvYNmJpyMs1PRliEDDc/GR9HYUSatny7jayTjoZqs2nO1kb
FrfJ79104dlzCJiayDPjfGO0cvKwvjbuntyUX15PIWpmIz+p65swpGOAQIDf6keKISpP5s/MPeAs
QS6VpHD5EzMzy+Ckq4JpJ7F9ip/rFwg2Gx4CHRYk5+W7p4zADF1DXFCk8g7sTYgAa0AH1BZsZOQS
3CWCqWFjQ7cOU26aOnjaIwTRGPIKxxhx8jBLY7TyyMmpYXz37nexCHkFTgRYbdmHgJZostrjPdxs
s+k8dHhJubh1YUbgMzL65loFcBlHLf/phCcm/fiFRZReBkXxk/hEjiuwL71OEQYTc675EZ/5wjJa
0B5nTVCzWxHRK5aCwfucOpnYfWcGKS6X2syUe+TMB/h2+p0kFU5uDDT71wqZV0mzs2WA4xoCvcyv
RiQKTyNx+RYVockYSWnH0x1Fnim6wAWExB0Zm7R8pwaO5hJdKvlELXzL2gB8DCzI3KW34IkjR1pU
whAcckfsmVNdxQ9yltqGRjMONickQKB4fBKFCJCaS3h4aQ7Y8hUXu8eks1o+awnvoB6s+VO1pR01
BJHP08+WyLo5NLVeUV4V7SdxbibiXT2USOlYU01l+TtjpjZc9iyPygNI+BYROBHwaHuD17a45JQY
b68RzSVr9hoSdfK0sc9tAha7N2fOxo9W8dvbXR6NDXsSWyNT5KV8ihyaJCDfna5cD6zbxZlJ1T2v
gWhTKyFfc3YsT3MMZ3psnm1walbRL7awVwXytrJP4Uo3lxzU8W2L5KEgBbfajGRX4Pd/tR/7nv/0
OmPl1ywH+0qyBY/7UoOUOJIeEur8SNWRTxXyCgdOUgtrMb55lqZfUvHbxGpYSfPQHKACb24h1cNx
81t9c1g6kRryHz5BvkfuoxKkbbegaVsPj93xh5nWzJiB/72frtyrHjhbX604PhrVAh39KEYkQBLr
FkKG/ZJIOE46WxEO30xZDQpzG8Wy9Oe6Kk7B9O0bwVW4UPaDclIvMvFVdfQpDB7drHkQtEQfG2ew
RhgUC/JcJi/L+2LKzp7ldo1CKztog6P8QtiY/BMMBR5P37LSX3OBgXtUXyBVARdMn2DTCrN38a6Y
Gtej4mMoYeykS7vX01Mshq7gdN5VXnm4jh1j38ydJyb0nmoXxGAMn0vRd5k7q23PKNmxghwZleKD
bmIECFXsskU+tjUiVNSY3nTZvgtuHB2bBFCbDtKCdLUJNMDar1UZ0f5k+qoVqqn8W7Eeae5ioI4x
/+jYYpENfmFUlJN87vgHQe5Azte7aD0E8GKZu7g16Ywm0oQpO8urZj+2aGlY23M1Y6y2O0tP+C8F
0QOvy6CoNTiVDw1KYNImSkW+YWodHM0PXn3E+sqyDB4jSLa5qjdN2JZhjWgG3KJsovOnEYQ8TRRH
iAsoOi1HrcI6Y+XFYcOXhnTMHlThPIwIr+uQuz5wgqe2e+lqP6skrma6tS1NlZOx/MZjoC+IbEOB
Gis67RwHaileQtak4lLV5yi7lENG6cTPNB/7PZvNvR0EWb1vKim5RLiess5Pd2ZECRCZBergptgr
Ad0ENLvZPXvMVAPzgox3HyZPiH0nR+VLhMdSVLBYVmBEdNWCnNqK0K/PPvxRrSWEoqXpwaaBolTz
xk0/0RO+BVLGNF+qHJsEfh4hbfcFyF7rTfsWz03rXFgyzq0Scw3b1FTfxx3jmnDDtkLKAfIOOnKJ
VDvrURik0uDmk9SDgRIP4aLaxKWPGKPHXOkBqRBJijf+WODTdfFaxJtTwPAuzUR0DwBW5w46C9Ff
ZlavuRnTfPMyI4yHdm17+wlSwjEiT190ZDX9cRykk5UvjZYoaLjzCfYVE7f4Vc+6Htg8U+Ct385p
yzIh7eg2UXw+DpTZOTHzca2RbNxmw6XgmA+GZnnuo65m8W+J9ig1XDCMy+ALXVZHH8hzz5QnWjrs
3nDveh5ifZ5W87HDbl8f+Fy9Q06i8V9UeVUVldAh+uUSeC6chWhEhs93CSbftYNww+7Rc8/hQNLp
1eHiTlVKc6zxCsDVjnZhC4pPeB6IC2vMHLHVJDE/0WgtH8psstgp1soN9IxJELvKZQL2MPtVmXu2
a3zP9p7iQGrxBldGgIc971ytZM1umC6emNKmUDz0WnoyxaLtdIXScaBcXMC9S8vhNCnDBdvLEYNP
z4eJddZp1tmh+IPCl0455lmzRvQSsBKYCvMry+PFdWW5b74PfhetOPUWH+qF5zQ+0vWALdYV0eND
KmEDvN+sMrKNUZp0M2/NQge76eUtEQOjS0BWkVvXvNn2+nESEbKeoFIKOshE57AY+RVACV2EDTbR
JzT4X98i/DVNcqdIG8wyj2wfWMDQkdY/TV3ufHxfY7ftEFPBWxvDQH4/zSlhkdD7M5HgUZJrLFVE
La6FpT63E94jI0l1deK9v3wNe/awOlAoexDINXgzy8AQp36vovjRCp/n1y5IAjNWKTCm13tXGFJ1
oK7YHCew1gGBA1stxvTo1oDxxiN/7RxSLwaF/gzUjz/OjAFLUrjPT1mghfUoVj08CuJ4Een79k23
oAz8qlk0nEgY8INIbbpRHzUky17QA9uPPHuuI6t5aKRSUYczq3oa3reoZqxwPQ3lPICEco+o/gZf
qQlIwuL/jlqABFsKYTWv2kZQrXXVyJlc/dnC+GKhb6PwCSX+E+oKgkc6jci2lC4qDBcUZTOf45UO
A2202MqnwMfCjWKKYkuqoEufEot4oYINw3oVakPiH/WSUjukGEuYEDfs1B1soWf8mkrxs4RvDxr0
Zt+QzgTds8hCpFHnobaVuRVSFdRqmpJaW59naJk4SN6pFaEbYln0NUoRus4koFAh70XOPpfgoZPn
05U2Kap2tGJRDVdoIx76pR+ee9u2t+sUpdmZviwzrrH5PSlQ6eIMLp5JISiwrq5WN/M+0wsK6xwH
swtaObodEOQhtdzl0Kxu9X0aF+i58DWfMxZ9I8QOBaJecl0qVly8/oSZYLtSDuw5ugsoOHosFMAA
nfYEN0erHPas3HWi0hN1E2qpjew77RXXAKpTR9KpEXAAPKYn4SY7nniWhvS5En+tZVGVShzuNAYq
Wx/9phw/QSjSPHPyRwOK8AYEg9Vk9HQLQIOYM2wtxsktXN7elpelFUK9RW8WsMK/wqFXWsdTbyxN
Fu0izOUDv81RZlEfD2YY9xkCM92TVI4M7pzfZHWogsv9AK8ftyGh6xJmh93XJ4kFlIleWy38oa36
jezKmh7Pj2UxPg8PvRoXTRNVzIEMgRSElw8fnSb89dro54AObsQqyr5ofOGil6+3P/pIvX5UWjKx
HWS7Vx4V0fk/AgRM6ohg9zzOd2NjcGXu9PaTspMF8t766vP1TULPdKGI1N+Ma+hxaDSl10I2cBEi
R1Mo9Jk6cd9EuY9weKO0WrdbzRN3rv1LbYE6JQABueIrbe8etiVV7FCxxVrOtPmeTQvBa5LsLMVS
ZLZI9O1h1yF6oDcswU3oQvry3118eiEex3KNHCKsy7QXU+U7Bt3zhURltfXMaLdGJSozlyjyXWZY
WMkQq2PA+oUrBS/5AGrUpvjDjVKwgkl2GEFpvDM04Tw7HETptSE2Ud4gi97ScLjotROPL0MiTXe1
QBHMJGXa9+uMOldzeGk5itlBi9UTcOgPgGkXtWMXwaYQdSs3FJTaqdPOI6l1cnd5epqI1EKx+oUq
gWQ1IoiLKfcsbVIzfsZNROCVysZlN1m1bRRVpwZM3mvw+VLRVV+0sMAzXjNuwggIuJ7evNKhnzyh
wPFJZiI6BVakKG4HS1Rwu7k21/h4OqwPA+a1ZLfgtzJA/zJkU+Pw6FQw3eqgkqeXKAw3wpVnQF6X
MgGbVhZ3KmFMa6o3LLwN/J4MDM4FoLZgQ251QG7Ic+UuF4Aieyg/ZIhXxi+5kprNfcKWYdLuHvty
0ApqGRhFpsq8t5hlc8czlj6TbxXgVwCjEEXf8qTOZX2sv7UQK6oIrr6wlBfB0leNzaVY9XG6+hw2
END9950ssXm62EgqYgNQXFYylvXLPHhcP/KJmPDZmGIlDVuoR7a+jmUagL/YpM+cauaBSWvwVIyb
FvcWRt4AWweh2EdgvIBYXMTxlksBWcSIxwPPXF7D/7/90PaiymMBPYdjBiWp7kuYbVpdFGx/vCyY
X3jBNFVaf2Y7aiQRjGuSEoHIAAyd0TukVuOfKXjyHq54jhcydEhR7MTQcDdCzxczl0Gxv0wgsi71
W7sd4ezQ+8ZtTajLxeJRMMgIKWxA8yRVPbvWYFf0BjGeXuedkZaJgfMlrLvZTH2G944DlE7HpcTV
hw5HhBqkGRPyl8hx5xLufBqh/yYkqz0kYpR1DA7vd+a1J81L5woWGVanXyJyKgDdCPhA6/yU1si4
x/fATSGZoC+qIx0gNnX0rIlY5gHX2D3h81Ix5gaFfsjAmd/hS8MI3YiOvu2RL8ViXRgE8Z/27nM3
n8hAXfhagY3aCiqfBTbpzJ4UkYfDA53XfzpAqjZU+e95hqShYx356FgDla5OLlMEbk0OFbCKCh24
NWZ07iY03stenKV3TO9q4x59pcI8iLPMrPlf8D9VdZgBhgw7pEixalSdqr5ZV5iyqCLYwEQAZf/a
HTLCKz87uQb+CZlpGu4Jn+5Iut/6t9SfOqYDuHl/jptKqxH5+pOnK0D25W8RKmdANpICdcGTPmBN
SYaviGgNEsZHPgquxMQwb94HY8ngOvIK0erVIBwl5V5ShAqioGZCoYyBs/vVBrgdKUDWhffr2Hb8
ahMgvXmF0glM0k/WRYw4RHu5YWOlLL16CdbF3x8kS56ellpZ6Z5/TpDEK2WqavBly6F/rgONVKTh
WZLA3ih4WWkIqetsQqiuBfAnoxN+4g0T3ai8aGj3rOCsR3Afey65WCeY04udTNe6i3iH4B6zmJC6
l7L0O8wNnL4gtaRhy3l/bpEWXMxA2pywoxcsUSjqQ0p6d493udWg4D3QbbdiJCsF1mrU8mjnjXup
NGjdfP/RCsHmxklKMN7ykCo3dewZg+B3AjhFz2LHnDBFd5sNSJrgpSUks5BQLwyMdoBsaCUXQhyh
gq23Z6N2IYLZ5YYMwKS1JWphb/fq0Rd8J3TdRFfoufDN1y4bbvy8zyFb1fKDeRuEdG0QxZpfeqe0
aBlFPdyRhnI9FyUm7Ulsu0vx6QWGZhcqkQ6N/LWMsEzMoR9E/Artf1D9caA3GtTTqphdTR6FxK4p
SaL/dp1sVD42jbQv7fnKQe6q/F4dvL4g8PFObb/rldH1bw3rR0azBJLNpRvM1esKQt4Rkqyrvql3
7lgeLm+1byWqSUAuT6aUhmgllLiE4nTr/INyuvQP4CPqizB4V87kPqKYamUzC2HZREg+pmyxU0xj
rIydpLtVEWABvbwqP/h+x/QPJMAe8ESGkI3d3EUWE+eVsXSdHOXzyJKLZVeg5q6jDd8UQIgeMt85
EFlUwEWJShxDhE8unNdR/MD2iObZ6u4dH5U4vUEz+kIVUcyHMKY3sZ+jOD6TGZy1Opes23EeTGp4
Q/HkHB6lG6C+SPz+Ec0iU0cBeQoe6JJxnYR/EjnpArh5StjHbQYPJ0zyRF2r0w3DmKbquQT0ALmu
W01Mg0p0thM8+nF5eE/jzrMyLx7qsqo+KLt97lmm52KLRyyWIqu1eqd9x39/+pzU2EA2J1I1Zo2G
QZhEjm09EDUtDBLC0XSzip3ecTjgmkNzm0kOm/4Mv5OzKZR+y7NHat+bc2Tj54uuPzZy+enFqdsK
MDlUU2i4n5+8cHp1CSsVgxnKstKk/lc6dy9GSjRlt9IkX55GPplX2+P2JRxGxcs5xu4S21ve8DpK
xHKsdtFI9kG/jJunnFwW5FES+NGmmbIksfI0IYLdA32Yj7IWerDzU6kMpqGBa9QrCCfhCrpu58If
ic5Smy/pOEnlBPFoGS9kUq9ZEDuUTO+BfV/+sTeRjSdWNz9rp0RqPT8iTNGy7CQS618nbC0jh8fA
J+4frhUp1ImnVpjBFs0vdkPxcfeWpx+X6Rh4bkYqm5zhGihQOKzxVtD0FFY++hHnxl6ykYCL6O7c
kAtjh0c0YypMWspByG5j9/05UaKW54jRVzu2u5JTW+/le/XxdHMd2Q3nvFqslqmnkmNcKBuo/FbB
513xJ5afqK1yY0Btrt1QACojLqgmbaWlu+HfRV8d4XcWIRpE8JngFNARp+8KvnfhsjsFSrKfcS5g
jnkqvm38nZo7xXAlUnJQxVo8WYp+E2QB952B3YUvRdHgzDu2Mr8ib5CPuZKDeqjxecyFMGDK4BK/
A/eJ+whj4uDYUlzVoHoeAGWnYZ2dmalqlPV5DqOgHckpzA0jFu4yo6sYbjSWsNsTKoP0PYGTs6xP
MldGrkuxSQnVDl8LvpbB4QB7qJ4oC+JfAooNJi2K7cnUw53xV/gkhG5o42ATDHTZjpT85q/NhzLQ
fb8UAdHZDZAy5SLL/ITphy1kiDrsFeP3yX7pj9nfjkLpj7jvKdjOKQv7FDSkpi2Ix5lzrj7pHHVt
F5ZRMhCe/VFH1iyF0GrMu0B3NZ5ChUjg0fmTDyI1T/3r+K7om2XoUKZBBic2soWc3XDn+SL4pDQ8
Kc5Nl8y+pydigHH0aoqf1C9uj+csSygVuCL9B/Z3xARzA2v64OTV0svPTSRsXLBLLIG3p9pEgUAB
LT70k8Q+69zfH73g1X7b1RqdNOlrsUmUnp02SVVyc4d8AYSWVL0ZLWkWKtwLkCSFM5QwcZmGZBtH
BUKbKQTAUaf5Sf2oUzYZY5vCyYw/dcZNoInR6w0I4FOrELtJNNYf72Mss5kfL4m8YkYaBVZ5uiS4
+zPqCLeYKPkqWXm3PGfBimui9NGH/QTghLYrHK+67wAT7nT5rcsZAmVDTskP1x+UVKvd7LBkwJBo
ccwhRO+EIabPq3plKZVjiAPNrD4HLFyx6VhpuqgsbDGtce7lDJwlmslYyuQcGlDnblbQzAfilQE8
eqoFBqta0vO52fI0PEFaCxCLGX77ELGGV84WRnp2Y/a67rW0fdjB6koHYJ0/oF0OU1TkrTDBMLRR
/CY6j00SIXpkznrloNiKlZQH6E19msRAN/ZroihEwtX7MlMVjwqg71TYJoJtDg7dxsPnGvd1D9Fn
i2j6iUx0lolAOde2T15P3VDcpaC2RtLQqzK4IltP1LriTscCZBjkWBaXSJYSQE2E8gXiMOqw9b1I
MjO23hivG2DPOuSID2NZFMNLDLS1JaeDQNvnd3chmHbtobb7P0T0bKhrAEPquis3DIdJLVS6SeUY
FJG5yOIb6L6qae7LnpzM6BZUBgZwFt+uaPsYnZfPxFgdqzhm/SSdU8geDgmsGtA30H3RtW6fFWsV
9Xw3O79V8pfSyE1qQXMfcFSVD+0Tl6hZUkj/HZs60MCzcYqV+vMELt9+kLmmqkfbN+CPNtLI0xrI
VpT58YSxvEZvc2LzBMfCJL9p3tcKQ7xaIQJ5DDDN0eKxJsdavpTOTtvg2IJ4Etyo3EWnzh6PYx4k
XX5+etdHM5hE2wZlF8WqIMGRkJCEgFnz/DySTu7n5xzpXpsY5Vyr/l8FLYUHgS0tmnX6aaAk/syz
Djhn0wjcIbIySHiI4aycEEfOWW+atEZzs7rX4jOs7qEb2gcbdwb71EW7XUQnIP861uAZx7dNWcxR
Xjm3Rkwl4tvFqXcddjdJpJXgUmq6YL+2sZ01fOFjO4J7KELF/+uyOokNAbQYncMlWm6imbTwvLtx
wlm7kgrJR+vViUMDWY46z/NPHkgncx3qjh5j95ZHEfscht/QBZT5u5cJhBuxl2DG9eyEFWrigh2d
F4l5MjGb0CLfM8sWnY2JmhsvP73iDQFDgoWf/3R62q47LIL4F87lGmvm+MPGxLpS+XmC8XT69csZ
5/2kpoNoGkuGILdHlANsuIzkq4y8ER9W8Pz1czl66+mXbscfVhavxFabBFtq5CPnvqhHyI5bTL5Y
5znHT2kTnXOky735I6rr7UZEA8+lxgbeVXiwONui7E1N7bsfLwtxNAji4PdkMY8fkR5X3zwhFaVW
SmcLIpsZLs1ZkaliPBEHHnsWdxelfrfdy2RjrQjqMAQTQLyZnKABlcf2vMupWrXEwQQ3Jh9tlvmB
IWiRUhUe0JtamPFk01CENI3D92jbvHM1vxjm2hNw4epYUfRtC5UNDCPbwHLWHN2xFYtb2N+sWUV6
eKn8maaTsbNIdLaTnTszJQ5ZFTyPB6Twl+jNrl5HJhaQ2mJmwp0fMPNyuolUCVRCIaYE5lcHAOnA
q6CeyHIp4G/UaUHQsH64tNEZQXQrJ3q1CNYgm/3vEnzhOJY69UDAdDSmOc9FWek5WbLMxuHnmol9
ekm7EY45h9/oDL8U5Xze7xoghzpIRdyIFNQOhS1QV4MOjBW5Ox0N7vj8mX8rOLOVEYYOwyQPDseq
Ybg35PX0DNbua+ox9nnbqnHeoQ+6XoedSpE19t6iAW3vMEuqJJsLGOwtXGBvPxmrnLAUqQLUfRoH
+Rljtj04EroE7ToS5jLdtEbuKaETLiPA+VdC1vhstelEw0mlLlgcPgjKuWrkjNrX7nvkgV8HQxHV
RPHeynOSqzx6kb/DiM9sJGuSaNNNz7iIZNFZVt6CthCEB4hfNyBp5FmjaMOBf5ad65VxjXISJ9e0
iHo7YD/ZV0XN6RPbhcrPTX7WF2NlshKCp4SM0v2UIDovdoIGF6M2qlSVtXFnhx/k2W3q/AwYBi1y
KfGWwMKroAgAp32jNhNZ+gE3iYvsXowmuwoua7zj0X2DmNjQK/y/9iaUXXDlZ+dOY1nUquP6D264
PNG855Z+Qj8D4PHOmeKOWAxSghSGhNR1Vfsj27fIetB1LYYBIDb1qpDWMHq/FOUbtXX4EG1w2u1n
xx0tBYPXta3ZKM4wB6Kb+7jpuHaIqdp7gdVTJzzuWdfPZpFyglZMflQngk4YsAUQ2DajlQmUbISu
9OXycggXWY7PWsLtPz32qB86+400q5m7eo3SpXheWN0K93SzChqsxp/d8LGkkoBk4tjKHgEPL4XE
gouFGzY5zRtZF8MIvP+T5wmM4Lg0YbaEfXIzBWye7zwt2Aorr/caAF75GdKjpw8Tm9UU5SEFSTWz
lK9t2YS4bpplmK4FwESBOnoarxYZFqhL0wC03W7EO6NclLmx4E2fzGnyRhXWl5bP1pCRyhb5PDEF
5el6lWtENOAz1u+ooFUickF3y0nl1d5h+HKzvTAuNXphaM3Ko9K3jkKxHZH8bbfACJpWT3FdMDxM
8ihISKfgD43/wYyGiaRIjJwMswjVaIdNGbKV4p7Yas6ED7RNXx8Fjbv3d8oJAqs6FCJCH7zBqaPZ
+ZTbI3v/KLDwIX7zbx6zSOw1bna/H9uqfd+mtv52WMOczKRPj48sDdzoRzVq6uJi8JkoAxirEe/T
xV4I48OFynfh4GeaQ+t1BhXwd4ZQFVvRe/s40TXsEkGea2pg/PFvC7C+DKjkA5XgMN4rzEYCrT6+
JOPAM4+7ajk/Uv2AvUTBFT4qdkmhBmxIkZa2SU08gbW8YSHB2QO25cIBPxEO3C9yqF3YtnGUPf/G
jR0DsZHqjAVFuv+8ZMCnBRkLh6rNjOtiYbQ7A1C3I0sqhAarXE3Y2vEmFpaGdja+q7iDw8igovfd
vYW3WfgEIPJxvmDL9eoy5yMgHbEu9aBA5cO1Wx39XVIgufr48mQIwpdrw2hhFQMD3w3GLr8LGbZh
xGeUgGQ6Z8Z5OVwI5qMvEy/lc85K6H1EtDvLzEO9ltG72Hw3CjXUUfHfbiPhH3pLkbK0GO/m1hwS
kiogBpeWPpO2F2Uaj8EB/4Q9BBGrWKykUneahMsFISDv8kLsfZ5bgX0ivpyfrjhNV7zbatYaZfd7
JR+92HvHffvcFwJnL3oOoTUlvIAKnDsNUdB+xASrK1+OmDTdwqA165ZYatVZPSuPJf0YkiNIINmu
WcXfFXUcXU3dgrXdxQTycyCIqgYG3JHhVI0r9d6ATOrIexUUrAFJlI1PXubifZ/Pz0X/XhdagOry
nONw02r8qmdqunZACPAyuufszeuxDtWg2n7bhxdG8jnW19WLW1IsuO8VBS/F3vKe1ffOTdN8o6ts
Z86gTGxuh9lAksc6R7XroATFXu2wqWOxdIqjpJ7P0gO494mDw5bKjTx3ISW1FY4kWFCMlRhljGkZ
4kdPhh5jMGLQ+ToiqVlaQpGAmsYVfJWJ5fbgz0Kfypo6uxpkqMYeN/Km1eNkINmHwFl//klyCfDF
RHaxl0vg8lbSrmbtYfNg+rh4ECrnec+KV670V3GDgmpmQE8LhgLy6b4XPIkRxM1dy/3KM6F9gZyU
g5ZVJpyWeINntq1O9B22MYSeNra+GvmRc0Bb2inDfIJu322OpFMvFwu1s5VPETIVCDFF7QO10WmH
VA+K7coiDnVjAkp1u82Jhi9//fQD08+M8E8+oTKYbVBAfwS8e/C6OD+6EaOlCoXqvbh6AeAs7cjO
uwAtavaDgLkRueMhYM0QyBohoeti/VaIWMtTLQmn6glmLU/40DtjwdvWTzDVpxW/UkwvhCukXIFI
7we4iHQ1xmaY1ArLEpA0JgGs2X806+VufRhaJivxpjQggdoBBvmiiur4NBA1FdP8BunzgUJCTLOb
x7pAP/NoVDo5XJd1crCQ86MNCusfRs/IMKUZCu/sxajQa4kDRGHVHWyM91X3oj4rADZuqYMveNfk
wGsaOrqGhHpdYPybeTslFFj7L1geuHYjSTcnk9tkKE6AY+OnEPI806cudRZOAkiFRbKL86Vo0WiK
ii0ZPjO8JhGsjCIdI8uQoebHCh0FkpwiQnmr5P2zk8NiI4wzTu8vCPXWYbc+HRW/upS6MT+6LGQV
CeEzcJVgAd9uL9bt402BECYiz3cTilQ9KFu8X3zeeMODC+VzJYm0F6q1/U4ghM5oL4BBd7OPIsHW
QXTC4pyZba9ry7EyEaaEeHURa8ENTvvx77Gf128KErAVVQpm+feguB4TGEoS7GsosoPCgxvuIR6h
cnHVOB3cKLf5chMhTGt4zce2d5m0XaC84vMb20DIvaxUA0qtZM5cnkyi1BouXxyqXRrOQjZ0KA6b
06AaxyZuCwNSJ+fi+26erroms32bXoLadXJM53CvKz9Ud5x3mxUC3lMMQyyOzVfFBICX9Xox2ouU
yCN78MyGMdMYACpYQX1HCgVasvDi1rvDpn0ON+EnBFjpYL5tEKbz257dbLJDph2vnAda7+naqz6K
f1K7M7mwCHPNkzOiBWW4GOB2sKxcFBsZQrfN9jllWLdZZ+jzeutO/06i23Fi/PzpHkZXFlJYKHE/
C9mBOaJZUiDIZInh1vQE6aFq4EA6ivV0E44XTS20nCr5IlfpgDy5S7NkclKTB6DHPU0DmDSKZ0sw
95YEFPWVV+s7cVYgT8Glpd6MD03qcMz9w1zqJj/D8MgZHw61nG/5d5stOBEvsQolyvPOmqGaO/gZ
AlhLT+WLUVj9B048t9+VT8ysOVm5fy5vSFSJ9gE1t+7E0ZtFPfAm2H6IU2MrPKORL0eAiAp7Z9DQ
LuRaloSv3nzsh7enr5HsOKxIMUxdLgwVUL8Ja8Ro7i7zYXDKXF/EgpsHVXGi2mZ6sVbOxlClKJiB
Bg2HvEJUV80X/CwxiKk3sHH3OdUiHR/b9RowFXAZIU0jgsUF4sWRTIBOQmhgEKVjAVqhrlknLX5s
ENzt6L1XYMpv6+omiv0asztBkIQXI0T2d5mjepphYw1HN4DeY1LjEhKzoqwzK+Sq2Uibg1o/XPn3
7+32Ffs0jPj5HPOhKrdPwg0QxufmqwBrww8iLYB6eHUQ7g4IaGYTNWBDaqxpeITVFmpMv+6RG0kJ
1CfDkeuS8EEA0WItvBDiTdnARvJvH69/s8v9ywaRFjc495p+PnZnKwnKbQKkuD5jyidpQbIq7zIg
fN+FnevdSDRTbZuo2l/hnilOdkXpDCKMoAh9jgjxXW5wrC6r3jJau2RrAmDpJNFRUTzyNxwkGUTm
OTndOOH8KufwSmpE9/by1RGa69cqf41nzq2SUFtlTO+Ti6xyufSDtq4Q9GHwMJn/UGbLCQwa8reP
eioYyi9c2HG046XHiHhgfsFBDU2mJynYQe9kbI9iHNYKqwdA7LabkPjEVHfD3aUxyP41WTCjo6HS
gIPz6+YanqZUdWyOad/vxrX/jprnUVPtRYvVxyXIK/lxW4eKAmOp8DE3RzX92KKi0w+J+6TOHdE5
UmrXjeQw6IJxAbXc0rhY0T8DafWF8gf5WsfsltgKtY/mtJyHkTlZZBFo0yuwkeJ54EhvU9dL9j9W
6kZEst50UaFpZ1BHnCUD6Ib3z4vg1NGbCzM63kNlbwcZ+HtGP/0PHZqr+UPK+0UB3xLlBmFI2CCo
KCF2e7FG4uwlwOVejNRlnBNmVxKKbydr9YLhE4PLU7n6OY5KCn0HGQRzRHXfi4GUICfjm8EDc+kh
61K3hA+2zx7TkhWkeaiiYp88sTyG744PuWDLz1f+qeR6YupDboAt8X/+RMyCMVCW1l+xbB0bY66C
eSVwV1lRVtzzG/brhMah5k0JytV0go4OO0aWIJM8H0nL+DI3MwdGJz0gTpQP1OXto96LHl8dg3cq
KH0jrtmT/eqCw06o9YfkwQPQtFH/Q42K0yfDYe5dJ4c5BjecLzRmeiq/kogmj6Qu3ArQSMlyCgvd
IpgOtgUvI0csiqp3rpLsDEnlfd7pxV8UDT6GSelJQQtl0XEwyWUpIj/WGU/ASwML6sUaajxYsaYy
QfuaGcG1vs48IPYkgmovywAtmU1CgW3QKe3JY1V21+P4xV2er7PJIuoLkThESkeoRjMWy8aA2iHA
3xHHiCJa41Nv2OMUVGjOgKpAKR02IIrfteFihjH1RJ7dWxXzj9ZBzGpotK4gIue80KZEfCONStSB
MEFeuRtQUdFlX7hsHUefVXcJs/qLB6vzS1zMd1cUMu1lgEj035FX2YDhKrItFKmqJmsFlmjZs57Z
Nc02kPvQB6zo5UcrNYVYpq5hIyt5L2yI0/ZC8FXYZKY1W60i5B4E4n8qFvQVXwgzDCj2aub+lRKm
wnnXBxggRofAuTfgZi6PZe3aJYDWG/hD93FruN4DKEECz/FD2l/KzO6wKYg99ad3Jz1MGXY8a9NC
DGRD4FRCm975kYzyYORWhE/1xzYmP/6KBuZX4KLZaxu1Ibpei0khI05BEkz5grEHqtPAjNAqX2GD
rRNnYGKjqdu8ARZgxAFRlcNr0pEva82FtO6MFpRZefT80pY6FHxqDnxbZRFqNWtqcXK4ao34yzSk
nBoSbmrk0vmVCbQmpi3Ll9hT3ZfqJv9sL+eGo2XC7uLi5WIukwagQqjadSlOH3Kqt0NKakRkdHxZ
Uv0pehGBw9b7aQhEzdK6T3uWQYmOYOhy624Z3xxFHPJyGgsk2KeyTYZPx5f77TqTUkSk04gEmPwz
tM1YZMn1ZQ1yVo6y9b2EMbm0Ab3fc+trU2lSMfO1VLJiL1aXumvSoKGb7JEU9owXDJJIstc722OS
pAvSTNyxjvG0Jfg2wgkBKNn56+xGDMizfoSSJ/k17xuBUcubC6KhGf/3UynX2QaGWXfp03UHUz81
EaZFae3ueYdqwF/KRopFIWsSmbEtt5rOgNWD/Ga62msOmhz4pPWWk7mIcSpxOXWfpbHze9rH+Y/v
xc94kYSV2+J+jwVrtWYP2leOwmW2BElu+f5m3Qe6ZAmIrHfXpdZcFCzlEgvnNOuGYy4eSm6YBysF
RvbrOxuyOw6vwkoPOUN4g79FYC3At+SM/+qbEp2CgXR9HGzSVXkUivzXavBQySOcM9C6ZgIV5JXc
FOSfcAU5jdwePkr88OSbqVqb29PmrvZUL6aVuHVpPC3T8N01AHoyiZat9ly1lnSEo9N+TEkHVDSu
4E5VD08OyPFFvutQSxNvM1ssknqXftZ2YsdEWB7EYYSFe82Va153BAzMfUxmTVA3+GeY01G4c0bN
7j/byI8IwoTgselBs37hKy1XHu+MjnfgeXh1eAScHoWGfY4pMcl7CYWxIhUzoKAgN0OZ8x0LmLfH
QACb2QrPp9M2hyB1/koUvou+N6qYu1NbM6apjAoBpTltOSzTGWV6V6ZZrwiavit1C4UregEYn4hN
FrCnrhQRfKzBI/2okRQcoz2mFOs3tZt8Qd5ov+z8hrGup5kxYF9VJegJq768fcPsmOQvAPYLkOQH
uwVCKvWxTby+t5/kLjhKIe3/1Q7PKszRUg/mbvZ45L6d4xDaxG5CUfOZAKXoDuiw/dfdRfhGBR38
BMfmkEhBRR02gkqRPyIAnllL/LEDhuUnzm/t1PWYsgQyBRvNQMziCoK/leiUw+d7Rp3nFTwR6uqH
h6t5ZPUVMaL4ZRXOFTRSFJVysizGLm2RN88zxMPRZm9DrjRH8og/fxneBGVg9ZJSAU57v4tufW81
2QkEQhPhSs0lA6Q+nJpRiHWWBxz4mrWfJ2l51aBxE9TU0DHtAmPUyA0Zgohgj/Zhul5bBMNKQXac
Wr39pt9+QWtmQA2x9wF6JfCFK3+osE8t2wQCd1FYWlkfAO2eFWd0c0lxp8erOC4Ln65pp/qr553R
egl750xuPRvu/kgzI779uqNQhJyBbqA5kUJHq5U5Ua4W2P/VRSEJ7GC/gSB4B8vH92TW9JqCJc5U
vLIG2oHCBEKwzFRK7RyTW5cHXd1/0FPCW7GCFSiTr3pxPkdzZVQqC2srbmGjfp00PgFulWf9rbj/
X/r3B3XoKmnO0/59xG698pUWNYHPM3AaSVLMTquM+OzFG7YFBtJeVgK+daLrlywagGDAf3h/0DrJ
XeSvps69alYNDEkJ9dw0nQBCrnwUNC065hnaDszgMJ0j7Hx0TZCWBTVZJXOzqQK0V6AuXd3flvNW
JtWztE00OPI40MM+TFyoMEcCL6yL49ABoUiSXed6urOnBuSPqzwIaTv8HPYoFUIgaulh/Ag2CS9U
KnAAXMnvYD/bElExzVfVg1NY/dylVzXkBsdv6PuAreQT0uPTAMqoPL0ESMpE7X404HiC65YCTT5Z
CRnyUv5MtxgbO2Edz6Z4u5LSZ9PUQ43Gp1HiCciv7SJrMhNwam+ya2sbzjRquwK1lkbOBVQnaqvH
4NXByrnsNs9sFcaN9fDT8E00aHEmpKWACtzO5vyJAj9dcJCLK3EWQYsaHcMQo2R/JK4RPVKDuuUQ
Z3zmv0DETc7n8aZI/1XgbtNaZLTYdSg/WhVgmZIpGsqq5GdAyQlwgA3Tj3Z4gHxaIJPlhLRmpFZ1
sGIknkq/p7jAugSxhJNf9lf3PGTkt8KvL8AG00EQCKpq8j5lBxYJa7cdcqR+3oLSoI8H1Er1+7v9
3cPd4/vh5SFmRrs8GABl/cmym8ZZfYxL9hWeWgePajpoWNfPT03Z3OlYzwdahkCzkZ56GlgZKUHL
2gAv0bW0u2WavSkyzZdNarBIFoLG7xqAvxoiGe0EirLY6kPdrEo6ye2uw2G8g9OhGxmGbQCN6/2m
wrDFlmOwY668A13v2Zrs+u1LSwa/SUyVmOdREc0/KXHr3qAYjhVDBUKSX6Kn+qjJVtT08aNH0yx1
MJpdAWkbJGzO+Eh/3Fd/f7lvy9Kt9mN6vHbLvKDY9T49TOIZB+niho19dxSYBL99lua1BETqdxYz
v7OdWa2eQVn18K1vf6IHdaBDSxFuJ261rILXQPInC+YplTai/3NkW47vxnfmnYOzSL+fphxGkHt1
0dfBROMb7Oj5XC8refYVun+FTBe/k8ur1OIERmJ8urTawliol8+NVFifiWKzFHxQj4++qKOHRuvU
1EQql2z/Q0D4csGmjwYTv4Q5PiFr3piDm5wijhxZ4280j3dvg6klZmf27JL4Y17EgoShGpCLsA0L
HYrLebwETAeJnyXPNy6PKl4s+X455CfobyzpvtqHPRoX5bFSipP2ILfkNfQXM21kvnlAs4BSDi7p
p75txoqRrtaSvK6ai1Vaze4a51zVpSRZpJy+HSxMwJLY0Zpy7JPLysn8dGiAGFqPSqTDSf3RjY2F
vBayiBPJPVq5VMWnJtdWLjWA40cdBq/xQgYvFsvB0Ni0zlE015fnmNp/n+mh571qWV9DNqiAm/b8
u94i/8LFgRtQFtC6jp2oCxijilhyQdaGb08rIpz1R2t27VacbJaprAab3d5v1UfAyjxKJTQW/VxD
h5rLsFbjSxAHEIgt4qS8ND091jt9J0evbtfATUHG6otHBQHoo/HbyDF87VFp73ytznm692Ouh+BA
kUiW3TnDtg3yq1EEK+rn7g/XpOBQnUqfpwpvzj9ugbprlzJ6SSuQmnaP1vfkzNtJhFBy+Jgw0Xj5
kzuq33sGmKeZ60D5scFnC0zFikDM4PMdEujvYpsPozdie2atRuV9nscsvFS1kIQVnmaxo4+Mwv7A
uATU21nfU9yEpO6QT6+g9FcHLN3TUqxbThQUlVz3ZHzp2Natnkak2sSzJt/6AcO2E4Ub49vtFh1R
zySoy2Wn2Xwtnu9K+i/hU8tkKprMZbAxzXmcoNYDJyyXMaKw7W4KIlS7fNvURn/VKXoahz/Ui6Lt
aENplPWcD5p82Pw8aCFnyqb5ZMYCfTToZ9lQPFQsaffcDVJwu2aD+RUwMh85L6FLUDPOHvKB8Ssk
/VHkuhonqjRykxaAjaPU4CP0GYbMElv8TTPEpGwO2/2VB4fAXWfXok6Jy4ZQwAwu7fFNHcwQyTnW
UGbNjrA0Kat0Q711OAQmCrm0HgwpEn6NKepVHAmA1cspDeFTWfJbq+IuGENLL/CZs6F1o/gpCmpA
W869fYAaUbMz76xE1Jrvc3QVipJZ2qNErCGejIgi/7FpTBjd9xmNodkmbuCH7yDc/eXY4KA3noxm
KJNaYsMt74JQdHXLTYTLPQ19WJ6i58bZUExw52tQLH/v+/A8t7FDZFpGrY+528E9q6vmKwqboI2y
uhmx87p5vO2Qry+DZBra4dHrrgH5AjbgrG78C5wqexRbYcI2NQhh/r6V5yqQ6N/eoxDn0kHSSJby
CYyqKT/cZziC68aL+EGgJw0hRwmaqBzqflrTWUHDk1dU71trJi7OV2BspeGmWRjCWARcfoRjEpdf
HuvkJSrZ/F84JWWZQMEnFHOzkX2HJ1NmWqB8zi22OueG3F6sbTzdqHtfC2og+SopCko+n6/PHMMo
G8FqIkS7yaZG7Gg3rl347opB+IS/hNK6ufTdowxXebbGWZLZrZtJSfGHTQbFWjoPz6bnrApHOeVr
iTY/d6e2Qc1KV3TTWatAt0tgcbgXwvGqreaNgB/Kwqrmj+BO/cjk5qhIMOmQYWOyLU5pMIHzYv9h
L94VWK1+oi7+Hrxay5syoQ6q6fUnVuKCXm0tiAWZH+8ksKTH0pXfq17mdIm5kBgvVKI+j5Mbm8sZ
dt1SP8FN7qWdIbKfbb2UzIYVe9Ungdr3pachHKhwHUivqCsGeDoeQjTDd9IZn1uW8KHNvGILDeK0
8aFeePwaHYSNHjo6RU4GzBlCmHxt16M4Ejbc7wUVYBaYROREbvgzcjDv6iXRR3+pMYaSt4IpvgVC
2uv4D2s76pFGh9i4Aa1Tsf3zMsP3TnMS8W80Bya+tZT05cjek66ZZ04UGZ+sdgnW9sxWeVGIhrTq
imze1gxnK6n8CRK8BeUuGtlLkma1TCE9+8NYlt4eNOtOSHj/mBVw4oLsPlJgY6CNZvpGrRsyBO77
m6qlgCwv5hvhH08SLtDYNPu2O7I+npar6gXWikw6zVMWdGaQH5Tq/22wo35at0zUl881NYgwCEwf
tuHTUJNXl6aDMJ+LNA+0b0UbaNd0PmCv7uogeqrVxYmum+JyqOrMc0bFnIr9hsHZtOiKApiCvtku
I6R7JNbExDprTUzPCwNQ9QPJRRyB/e/jNq4pxoVvtSARHVAu5ae7sReXBSXHHH4c8ChuXBvYR7rn
xwEjSZod2TZCAbLVdguKp8dPe0beVEc+73hd34398EAy1RLy5RuuKemk3sMHjT8zEeUfbwxOMmMe
cW0xnn/XOlVQMsprSdJMJb6yhGMgU+rK+D4EH23YThaUSTtfphkqWLr3mm/I/onyxSbFT4nhbci6
+4ZZkxQiTB+TdINrmWXE6uHAZ+7lgq5dB2A5miVpzPkVt2hZ/vLveS16SVg5KkOpsU7sAgS0LPHN
9PCqZ0k6aIAwAyNBaBUrZb68+1OhE6rbWtVQV/A9L4P3wtcxVlY0GPU7E02lLYdpWSbc21/0F2NX
tTalUN48Ut2Cyj7SROCnYxgsVfqLzgjOonxr9WP1pV9NIDTAfVEPT4Ft8dJNNDsMdRokONmLSXDf
lI3ek32ZySRdwmQsT7HttjJ7CmuZkFblsiynbPFgWi/MNk3xrEw+zv6peLb2yJWbcvtDfr4vZqb+
/7dlYIcrM3wmgwr5PFtpG+Ca3FpuQC5eTQR4RN8JxXf/ybQVe7dFYzK8yEdpwdWfUh2btsmD4QyQ
kRznLpsaYEOhUJ0Bl0WAfz3VVx50IAndgmrdKcUQq1prsxc91/Q3dZxVA54Iop+A3qjFDAlbovCN
soLF6zR7jLCODIbtejYLZTZMrjMv7o6d27iuKoxytid5YcfsLhospNZ5kx/ZssGocXTbwH5b5+HH
FcRObqEvGtsqRxmMIxBX2GJbHaYnaj7U46Hwwm34Rmeru3dB6TVxZi3c1rgBqbGAK+KmS/CMDDyA
RB5kgkLRbexL9m8rXlXM2f9+T5Gb/fFMnbBN32pbNDjOC02gcyjhDaZZN9DV/2A7I0QkZdQGyHMV
r9SMEHIMd2qg9kyefyB8ExXJ4/z4be/BPDp7A5DimhsR/UCgvDiZ+3fhSEe8j03Zjn/fcNWV7NY+
ydlbIxIDR77VIcIaHML/i+riNV579lfPX01OgdIasI252JwdKPl4wd48QGO7e/I0rGt0Z0aD0T85
SCy07WmRQ2iVcSnAuBuYVEGlUqlCC5n2QUw5FL/6fbMIUsRefXPIAiVK1D9jV/K2IzDs7tdtN43+
BR6RiG/6rXtNKLxyvdNfxyHnUJE4MtpEu/FU3cHDCoR7cr3AAhRsGobA5uqJT52HaphzvKgQbl4R
oVcKl/uXAwU5pKFFSFL2Ivf8sG1UyGxYIWpln/OhEvnJRlzYIY4j1wVs8CZ9oziqBMXeM99rUTww
RdTrRFpKV9wV5Ww8Uln5TQy9MTEiXqa1JEi8QA+ZYIqOWol0LV8shJuCnQsBT8nPwedOLRDhYpI5
618Ke7jDKvh/g5fI3aet7qkIGlWrNwCud7zfU1fOC1VrA095UFR6D5ffYEb0mKnBY8IFyp+8+eM0
4dATCIJ8negXpYtZ0PBwMtLokWbfcALMYc79fhrhAxycyI5shWMD4eDyGugn7xfVVOrSKVCbGK3s
BUKX4kEWEU2CdKFiNhsjGkjOrryIdFc57L9kdFej1C7Nf7Jz+qxTRv6KgniKDIlAips21rsHzGHe
ZHjxhMcZx5QcJMAxU769rtB4pa/fiaMqEGWlVx7YXsF8Og47TC+lJhvlktS5I3ZWgMST2IDg2rGl
wcsLVhsiCjHYMQxmL8noy5bir1YgJ80uvR5Q/RU9M2BO5v+BrzRgKuXNR4NGcrI2eQbTXPrknaXw
aRJWRhmYo8NLcPLcznsm0T6b0gawvSt8GCjYizVNxSk16GLq7uqv/QAj2HnbJK2JO/brgOIzgJOv
kDsTgZ3nVLIBbCmWkrOkUVqqb+Pxj7QGrAALyL0EGgA5tx5sIE9oz3OmNWgtnSiLc/gu2ul9wuYx
eDW7HEfZDoc/xY2adcrnBqxqeWUnk7cgVQC/aDmqdjdXDlpfKvdghcEfWccH6FVV+8yTUrvTBXK3
LS0nPFJ+SfMgdjcYCdM+AFeuycVJ8SjlVEzd9kv+zoBtSCMiiZBYHBY3rFjsbX5xYWnc1FyvKOrw
7YhuCDS4yM/cpfvyZPWTBUk5LwRwmA+/iJHXHIt+eko7l3Dk7TuvtaEyyIlegwLq65OwMJJNy+wF
nRtknnSHhIbAZurtx0OPrOOwYN2J8stqg9FpC66FiGz4RhW45SBnOMp7rFbvyk8Um2L/05P0ywWR
tbmcI7/Y9fUBQsA6wl6O/4FAMFfO/LfkNoFL7e7qevaspkYSSsJxL6nCuRN8myxWkmycRSGFhTEW
O98s93srSA/ltTeFXrn+QczsKF1DNeo/IYGQYwHdFgiVEscyMJqeWA4lPR5Q+cZk9IKmx4J0e52w
um1ih6TKCXaK0PNhlsRzxBJWMirCAujAjykrlw+nk5L0mgBp1z9hGVLNMpe8unSXkp2bFaWNER2T
/4Js+0q7v27JCcgCUrsdD3FaRSPid+zOrqRorDPB3tt/hYDoFIueIggB40VTec6SAEu3SJmGuxYL
20/nYyt+A1jm35+MDNY1fg+WxIrGcsb4EDHgMj3ByLY99H1tS4BR8Xr+yh9DA0T1zogGx5KLmmIn
DqOiwDLPqioSKLwKRVwtwiRyqvqx1g66FQK2jZ7fsWEX4YCTPqd59na4DYMxf7+/qeROPTBbsRZU
ApMQYVk9Dot2jDMtHaFqSMnMKVl1T0nYHAyJyiemm+FHVWTI6Bnr4VzvVDBSqrePDjO6Sbj0KZV+
bhj8h7VF5rFL0tFcKzGkZ5YgITPFfFgJDyOrd6jCGl/cQxW3pHqZP1DW8KyU76rdR4tYMbfoKNwu
h5yKC3/vbPkC5kHkvNlf4C3o/HOTBt84AN4xOKRgDv9ywPqycX3HNtgT0RItcvsSxFbuF9jkNIg7
dlGLJ5Usne51t7WVBm75JXkqxs6QQnFwFLIRtR2qrQirUeBbGnOCXUoR9e+VFJZyG7joU7k2xMzK
akzzTHvlBTqeI8pQARndnzdNUiZ/Zb7ic5kStesNAUR3FKM6eQAtnC3GXhpPhADa+mBDps1WCVPf
llsvnBKG6mYqz8XeuxpZ92VtsB3i4QjkWOXuJLJIm0JZlgaIfjboN2/MCnQ4lud0BW1Fn+TLSEuA
r2YafH/fUCSZdQ3viIW9llgOyIvDjYdxU+bQARY3lZiawjbqY9+eKF0O+3RGyFCAkRtsl832R5Yj
dTq1bcZRflyM+JiUUs6ITxacd26k3L5P8o3T9b7eS+hd4A0SESOdi6zQOn+3qF0clbsvfp0jI+3g
zn5NmqDZpNNv9CRlm2bLm+3ROTT06BCW5bmygtuCecNDBXvyE13hLE228ok0iJL+2VwDrT7/XUsx
dwc29KZVdD6MNuPJMHIYBwEdF5AigK10J2512Vrr4dMhNbN+DIxCbkZvG6WigmBH+LyDFQfpA4xW
TL3pOfBEsKYw41597na2y0GFC5Tr/z457JmaPI3wmBHROiPekRHqn4tn4avXHhs+ktUYUS9Zebyo
suDt6/9S5TiQN5z/cRsBuSpYvPhthp3Hv7qJky1yYTL1w73zOF01zCwL4ICXjMVCxEdb5wuULHrS
rrZifqvnZgqZ1K5i8RL4vpKGeZ2g9hIXvQNdr88tXo3Dv9YCCmNRGqNGYEmZUd7Jrm1Cb6ePAL8+
3RPsx40DnfwloHplUYFEZ1UCCVCi47Dr5HVeGF/MHJfdcTJ2KKOCW9qc+bshbr0wIsKGJ3HfNQtJ
/SAYUKFkkW0147xcBJsaOg11k+eyJ8B5TqnGmiXZzcaY/jkepk8aMgI74wxqOaATmSm6O5vpYaWr
4qCghbKVDxIXgllS/mO6RjIMkFeh8dgehGNQPvaLxucvjuzqHr7zBdBpzIm1Xw3AGsqfFyARxvVG
IsbAY+JvRyiB63vm/HR+VU0SYXQoitoM1yt1t9HFGVfs4AX3eELQ2thrnw3Lk1WCN3UyaDkkqMc4
JhL/v4n1cQU7eqCD1suYsCBEQL/WVBuY/DJNJXo9m0lQAYgKxiWvvXut+nnS/8wS1TFoDEzw+GAI
lM3SgxlZpCA+yaCt+pCxAXMzJr8BYwT32VxjafvkQWPRvclCNV1ydZpvYuZHKPHRa4xsVxHd3AEN
/yiOptfg60omSLhcSqSdPCUf3Fe+DenzymhX8Bk4aHTLVCmVGqR8VXIRGkmz78sckIrsy9X5Am69
mUihdstQlofCH3PdAVXuUF87pvgczStBM75KPkClSHI/ss6mlyt1ZBOnhcuPr3Q6n4jFn1Qv4KJw
UBR8ijSkAb5n9Y3OpiSG23u0mji9oeSKRdroKi3EcxsWa3k8GpXOEGbR3mNezRCzChcV48JJgbJ9
ajnxiXPrxkXcSwuTJi32liFHAAwnXnvzhWrnfaX/2SlithGZXpVQbBy+KagkcFnAONMPDqSY1Gel
y/M7KgzStdRmXTlPVBW/mB7iocjhm1f3YIhuCsLEJoWUaD4KS0TLBmbV5kBqUlXVoiG902dDNQ7k
IRoW2K1uTNcllEU9qGNAW8VqoUSztJp0Y9o72pByIxv67Op+SUbZmi8kCLXaUUeR/d5JrsNq7puH
F5e1pNWfbDlLjchTmzU1LYPEZbyRUJkDX1r01fE/e06wjP1EBZ7o+ChYxxehe0mxxNj4nUc6M2U9
TKe/8htgQGKvINGA7j3aTvLCAnyTUqWN2T9TUJ/PFnzmDB/4ehO+O/4tfSKTj+wFDp4/aIs0dU6G
3XaponWOQgsjc2Y1wOonCCUpZ6DPPD+3p66bvxbrVtUMj0+C1JyjxAvoEE8DELba012Ay76hJ6GC
MttD7/YRvtNaxt49RbWLXSIZJSnTFb8skCibSj0L5B9RE7wSovuipaKjm9QEncrkTX0QYkSfwGPf
Kv4s9gzqGlWX4WmsnBqz69Rz4bDAl8xxva9etAAir8L4WjCd+KDqxBsM+Hg1gKc7QVymPUBHTRrz
sLQIjZGJxvOIW+iu41NXQLfAO7+MFVM65FxkRxfoCmOWkVoTmZuCEepRcMyOz0WtjRLnhVc2Za5n
AiJl/exptSRDXBI8AQfEYPMQkXA6aLrbjqavXYBRo+G7pxAuMV5iDBeyCQxAXx499g67u/OJRaFB
dQJ5TBW5sRUk1w6Oapt924Fy4jurud6znS+X+yknBOlWdb2ldvxK9ARgqzOOgeT2JdTx2je/K+tX
JqpzH5egijCChV0tVpXhe1ZQJI3PJwTgX2V4E+nVyeup73BWlmWDbt82T3TALzEE9SS34PVUZQ3/
2Qf/r4uFc8ZyMZj1QqG4FtKXBtDpjw2hBONKVAAD0kAPRieiWV/oy5rl8NQuvQt37+QrVP1DHjal
Wje2eejyioJkwZ+eq6HAdKUcKJJc8NSj8FtEJTvGzmdekWOnXzJweOL/bSbgmdTGRi4ZAiMFGso2
GLgFHqNyQasvdrKZPeO4Ajz8rpHz9RSLQtX+0+XF0VCJYqOncyFRsMgwnmi3rEtFoeNGmFcrVNvP
u06S3YKLwkNbCTev/dQpZFEwyNS6lru9Y1dozNlFNoquXRE7hyhTI8h6UUbmp31+kWxxXsbiT+mN
Hlj9Mf/kMX1AOSxTFamIGMT2uC7OvjPJWqNcHiUR2ItAzHps3dNxlSSDCmYMbLIXARcrrUrei+6g
ZSQP8rogdnpEYl19Wu6OhZc2ISx6sV0AIl8J5BUyCvGazk3bIeNkqtUO5loaaTh1Pxf10wb8g+U6
4ahi1+yOPwJ1OB5HTNXaB4ttL1itCfhJB2Iwj8CQA28u1ba6ILNbntUQE8OrO3y40TbOH6J8nokk
6e16EBBfiXVgJ6hBXtiBYK/xLbpQH3sgYPvAMklI5/uzFoJoKUB73tRvNuAXvhCYSQkix5DeZ+J8
12wA0Tf+Rag3c2eSkivuUuw20vC52/XGspTM5wtH9pAyi3t46NeZL1vKIBU6AQrxld3GPfk3QyVQ
evyZKYMFSHtD/nk+H/TtX8h8aYRPbJkX5ylwyzHjuLDNwiRpMGd+xqT4SE6UIK4KApGRl8jfANeK
8EtCvimbg9Hr4wBq82oiQX6k3GDoN7WsGx3o9d5c2AX8AT4a6yyu1MNWc9wzi7Xb5hEOfkLrsSpU
NjsG1pedpiUy+aZP0rkGC2+6EUkFeDlpRD13zX8JHNHgpfWlMXv6KKxxRDBf2pK6YqzO/U/95AGg
DXkHlqxgu6t3+wB496WN7WsYiBXQ6+W9S5fVEqR0OOXExLl0gnIOKqc2fBNs601sbXZazfJtgH3V
YzPUb3cXVvh6XT77nZ3608cBVEOVy1ruu0F71PsZueFUjzHJPIl8qEV4ofJp7yL0UIOHQ9qleF49
KHu+XxAZWflI5quNLZtXHQuV2C2PW3Q7WWWXydL9EaLlMO4eblDNE2BcEbu0hI8gqoFGOtRAPoqW
CNVtAHzXhjzRx1h4bg+muloT8j+IcHE8mQ0NrLwN7BXMc20nrfthz7wrS8GNNXQ1Z/zKDcN6yEfR
7ozYvFeiFEG5XN+1YGVOXA4a7H6nbnM4UemVK7zf224EQg6Jtc0bTiqb/G5jjZb+wvggKOwEYYiI
SdjpAzJQ18y6Tty5KISZbighu3UabfioyAeFYyjrR5Td7JOKF2bhhT0IdriKPc4r6xc9oYuywYhM
w43ax2DrZ70hbnF5KLm9oCB2BxEhPCQXRkQ9x0F/A3UD607IY7Qnp6Ymg/hEj1nPk+73Sh4yNb4/
ScHB7ntLRoaI72xjw7/jrgk29j9PaZnlQRiGgn/KCgnlWx24Y3P+j51fcpBZaodv8Goz6LIhY0ap
OTsUiKNZxQjoWtDwVoEOD+ydjz/irMBeaevEc7UtFsCi0eRajSdK+Ftfu4ZAZ911Ah370DdmA9i8
Kh7div7eUCqtKyVpYTBUEvsNc1jUkUAWky9aKOyqLnBfR+8OpL/52ZbyA+JMi2nkLjSQn1jI66aJ
zEDpSTfxYcq8BvJwZnRVh86RGRuVvfwaDTcJMCp6sbAWVkdW2sX8s8+MCr7CPgRaeDTwBlJt/rAr
Xrypv1KU79OnVDl1SHS0mM9oDJyfy214JYG2DMXRgp7Y8okekcps0WMK1oXJDnfAEnj+mse7M047
qOP1gvoD7cD+Q6FEwCaoT3mDN1stjPgdLGHD/b4yJeSbVXKTbCnNX8jxHNVMifJMkPdKFHEvY2aH
p22nmwRoV+OO1LNG23Vv+bcNKgtSKbaLF6YuCb3MHlKTZwD/upY5tGrsxHFhsxoBHQ9HIKmBOgUf
wKe1S7Pi6yxun0tHsvSK9pB0zQMY9ALQUYr5NKmtN6XMP0JgosD4kgks3Dp7QDzpBskeGjV+5n4x
Y2xIVZqkFXpHfZ/c+I/EAaNeucwLr2K2jJIx9bp/QrKiN8+kkMieEwfBW/XBkUCiUjCPGVORJ4aM
RJQmHeRzoYaq5TtBx9UKc/kCn1q834ceskj4Z6zgGpiRQaWThN1lubnQCt7j7QXOgRJ4FoDBm7Wa
KxtslE4GfJWDwZ9xOB+CYLZ5piTJ4YTzyJksRKqx2d9uryoY4J8kBu9W3b3ajZIATjFraMnPOdi5
Arm9xyzCTdwnsHTf2f6UMZMSr9KZ7AXlM+yb4jrV5V87hYKQyD1DgK4/kUTtpKJNipk77i5t6R/3
riGY6KpxjI82kxMS48DZdRLogRYGdad039XSL1yBKfsj94K11WYjEtGv+n7EzxEdneDIJpc43OMc
h9blJ6scPAyTP6Fc3qO9NVtZEaTw2bVcZcl9W5E8nGkNKDDIXxUyMxkHPqv8A61CpnzAVgA4KRUV
4jEj/MFJ4Tl7/83ls0b957ts5I7C7tW6oKJGn/KXkecBKVjoLNxiTEG4m1etfadDUS62xBEU/yJc
xSCH569M5ISWhD6V7nnXr+nm9MfFlvZM3nOAEa4d57ATl8cjtEuyInlC+NJgMTl7WUPGPtyatZdB
rRGfwYlFqypIFCFcAymXErEoeop3pqkeO5BaNCjgwJBFFKBoFbK9iIPTegGs+eppjewQW3XDQsTE
6DAEJzpCkGYbZS3dnqIqEY6Lv3D0aRNe4FTEGDbEPzxTtpK4VGdV5qrsN4qnlMoPkrNH81dRILz2
iKvqCJjEg09XzOW+2aZOIv6picA47OHj/YoQIUJndWCYsqp7goU3AweWhqD+jvI9E1/vHTb/DFij
y5IoUsIG1uLnxBUaD16rOE5CmzVjuN+HTisoepcx+oABNc40LHV8NM+D6mrqPRcP9PDxQ4mIF+85
Q3KsVYZiEEk6TNIwlAMyyyHIOPz8Elsj8TMpDTbKiiK30vQYeFIctVszghRYjpCXQT1M80RY9hE0
aQTWd8q9aR4+Og0j+QQrzXVwPL89vZqsd0QvuEmHKDigxG0DqkBXQBoF/wncJPVeN5R0sLHSRjeY
lHBZQqOOlMjvth0OVO2JjrHtpUKhWUXKwHnhCPVJuOOAHWq/8QIsyHdc/F2ZCqjBGP2Q2PbX123Z
kRSg/uVo432XfRFb4zvvNjJY5F/DCOe4hfVJOid06iByErMzlmCCsNdLSnd3MJiQ7em5PK+mfoVv
8kg9hAgIxyV6sTreknM7HkXZQrpmv85CrHxUxqvNwtXKIp21FtHR2xaWvgjNOqQ/NU2jJSO9n90x
NXqIv6XVkdmsrfaWhCjAw2P2XjemhcT7/NmKLuQdaN41W7zBXFw1suyYw/i4brbKLhcV9D0UHU3j
n8ZsymusQ6B3EWPAhDbvbprLKbKed6qoMxUrskvAoiztxIJZh0RkO8E/IRnOZ4dV2U/8GBwt49vV
5EGSbVU9WpEaGK3CVTmc4N4DS2TK5guTqr2uROL0AB6PHuc3xhyjFoT+MxGqDHtpFpFTbHwnMa9v
OgN8hwtVhNPM3N96RR+Oc4Vy8jT0+kksLGE1G1HOIBaWkiREBY3R1H952HGrjZRp30ucN2aDO0aj
lWog7ZYy37q3oOfeLZZgkMz8bJJmgxewViQXWLlBA283GOK3NzgxJWt9D3elrzSVb13ox+Z0o2f8
NYrvmqHjln6d8kKKWPlSUKv9hNMfJ5m0yyvHt+s8GlkKb4mQ3+a+pzWHdGOy9BoKCGERrCAYGrta
wiroMZla6dn2nKdEpV7tyky1E/hGqbBk/8ghIVIfebiq9IdbLzbiww9T+aM4Ker7la+kRhqt+Z5t
OXhTtVFw7mhs4w/8pHerIao0r1hh/vU/BgoqLv1qDL6udQxnBbrPkDudbC6OVVPflANTdV1DU1gE
OR3nPnsQaFsjfqRWF2AJsTe2fsmXjPUNJ7GJAWwwZkfd9nhY4cBLKDYt3IChzKe9UohlK873nkiy
6wAFR2XOsdaDyEeLoJyNbzWjtB+qzxd+UzQ/jG2m3gBDTvEe9+w19rdJSkeCTkXTyBh2syaA0Ge3
ji4XBu5djBvYJLHVyx6Lt/0R6IpIm8RiN3gKyHAgpR13AxBLqtW8aPUKoIn+vQQDAn0Bw57s5Xbl
6O/RmSa95uZx0jGV7w8v8xjmbPcPErXo9kccaVPMeVJLOC7u3s3CSRXp/FsxVjpwgBRJtIqSggkM
YXFfptXluxyi3KyjA0nWV/xCPVeAQpQCNS4fpseSe970SzNrq89UjJ9SoIlUJvaHlas4vhZ1f1AV
aqVid13jUN2bpRzUoiKLpR3sZt4nJaHJi/QTPUVsseYbWC51HzW2EK9JGrRrmEwtDqxzXUTYC/0D
oBdZkXD6use08+33hgDoxzXTJ3gUfZBx5tsW3b0RqDmz8RlVtjlnvptPmbSxziwiimzZLfwBcH0r
252k4CtIu8hhIgze0xYCBTAdlBms/LehW6L5TrzF8klBDZ6G55cCgceWMxK+RFn2/L6tTAiU0Lbb
bMmMNRxS/c7pZJFanbu59kUEmYR+pcNiZmoXclTJi+NE4Lki2DWMvnhXYKrCXPooVc5fZnR1YSxx
vSBr1NLzBTQosOG4G0e4lixPDwvcLuegiTm1ZXzYkbYQNxTNajyrLtgEboeVcvd5nnZ4MYUCKVt2
pnBwO/44ybJEtre1/GW+lXP4Ef6r8MAxnxeFH+2an8oyo0FRh4HMFO7qQIgFVediklro+8hWso5R
rb+Vzr26XhU/T2ea+IHcGFvdyCmMOqsFmmQ5Vn1oBjQ/GST8dl6RQmgd2ZNzPFRsIy6S63JBd5fD
h7NfirQZs46uHMFtDL7PyPoPhd2UoKlnKMbl1cPl1s8WCwo9QWd+dUu/EPg2tvcJVxKKcpWKcno/
iopLe91/PIFM9DllMFO2KjzsCZ8YDzAaUES3b6kguGZcnyKqDJSlal5evOoOG7ZzRrYqAkgeoy80
QKJ3ICLcA4Mo0gwHm/gSBjI8egUqhYsJv0hppcLMQrAA3t9SFT50afDFjN/aSoYfkG8efvNPNEyp
V+i3M8pbL0LN1b2MInN3ds228+T2jRWkDTLNNCj4BOreFqZTxF8WVHcpfrn9aq4LZYPL3UeK9skl
NDpoDT0gqSVa9LKWAz7S5RXkbegE3GLmFbcDH+H0I7t5yA03f4ZSQdRKl75tGzNDo+7B2npRO+1X
tlbbG3Lvnj8GSUprC1DiHQcigwdt/3SDkQf6idR4ElRCtw/Z9vt5a717XuVkW2b4+OYAQCuAJWhT
d0hKkBqTc9sEo4FsjSL06TTh91yqHoUq0mGbcgUnpVal1IZvjjjhd0DSIhzbG7GMBJrxf4wCAPo0
HwSxUDoYbOuSZHchRexraFJZqwQNb597LOSgtyCH0ofq95fpB5s5/PM7DLeyTnWKGp4VZ/pEFHGK
wcP3/S/KYCa4Fcjzi9ERz4rnWL3X9y1dGsuTIl58bJHifJgNiWPCUkgy0kMDBBSAZ5fLaz6f/7Mn
7EtVmrV8DFvUSrv1U2YI/lHYLeUQpFXktxzKyZKUPiz7wudh5c+KIok7ZcJU2pC6aD67aTiVEb8N
My3IHlA882Q6yjP4Hw6vSfmCsNXMICJAdqy/UQLa6UW2Xr6jQis8CdNL0WxESkvTh2z9Bc10kFem
RnX7bmaAKZ4ghDMDj3MxdFh9SkBT1lbj6GZoNG0WpT8WN5RwInE7JU1nogkBJauZTRbFMpPKHist
LA4X9IA5rdDreygDZEVEm7pzJ2gq5v6i3paM1ozRSzp3mjWbMEUZxrmEgKu/DmnSWS8Ly8bAy1Cc
CuNTh1CnkOzXvkmbzNZdK1UWPON2gb7f5/f7qJCPywL5bTxrzbdtKXL1/iodvEQPOSkU5BvnT/V6
q8qBx/8Ud22M4veZvKr4fSKGlhUMNtSxMTtjGVp+4dymqT92OEQQ30mys8+BgJ0uj1Oje0ZwDNM0
UMvmcR4B23GSZ+309S7AWFrBly25G92ZSy707UFF5tIurg+u21K0Tx1Nd/BJvLeh8u+/O+KMN+YE
S42OJXTHUxsxk7CImSeE7IW5rQyAinR3Hs/T8Ipd+y89ggu1azdrHS8FYnmp8D71otSxY82Xw04I
EQdmnZDaWX3YvccZS+e/FINN9JF9RWB+3e1KT0u8lQAXnam0NCudhbthYImykbc5We6f44sD25kl
6WaT5eCMON8FcLdzg++IK3LiuG322N/WBtE67QTYAKtR5yHCS6KZlcSYDZ5W2IxmowJfzfpchtwH
2nkC9+JasxMVax5Ow8530cQ8tvOR+OutPLqy3y+6st03o1/bGjjOlMe3r5E6WJc+Lxfhwng7nrCS
9cRzMVMFAVqO1h3J3OPdzu8sBwt0BqxeRk4qdUC8W7wtfvH0MX5IH0HGKZfsMlnJJmlsLooBOyrS
91VAFV1adncNyHqC5QEkzKyVL12E5zHPE1toCOrqHfuqPKZNW8IKJ7S3COUJ+AJUqc3DavmWgumI
O8aVwOTMVsXTobgJbA/LJFPinUjVAcMsL6pDnu2pMXE9NBOe5YORVh5rG/z21ke4TbBqZUkCcQ8t
+1TyeEZjoYVL6FfrGQ/crOnnmsRiOtkWMbEtwjeDH+/atGhhCrIYLfYHCa1S/BY3Ebj2JjLDmlzR
4rRZQn9xi+LnWbpqN3qUF11APvARJABSP6FnXDHeSt2guczaerkGFiG9UMGfAlnGMsEbup0TEZrr
muBHmLWwztoQ4e5TOmFCKArojP6H/KToGYaYS+A7WFnTh/p0ZIekAGF3OTtWwwMHDQma0klcRovN
tMkr1PW5Mxmk7/gVwvpZSpqd0ytvKkUN5Kn9m9mBAnEWj+b12no1YwfnNAVKoQndr25RH1mRqd6E
RIXx9A/4FXD1LbAZO92vvaHf6rflS/WFv0bcyfCMeSS4//6qbqqfhU/3K/UTdtDHN01EYLwbiA/k
hkZAU6MRKO5u/eVTEqDMFik0XRW2X53FLDnM4ZyZGzDuVyzV+M7XpVD+36X9qlOnsNj1vJsJHCao
JhHBtJdDWinGkyF/BB8+HQYT4wyf8GcbBlMgNg/muPdJGaNypFE+jZOsVIqQqqoabBXrqXDKJZFZ
sk9K8VQMxuOPXTSciU72SI+kZKr0E7YXcPE21gAdUGBuQ44Ec3Y/f0cKsWKLFyjMU/RBWNv/uYFl
Eo4xs47uF4DniDIcRNIH4LtVJ6bdyA7aVYZRPNlQOlnlM3C9/JcbcPr4OiYJRxVY0xVtKw/Tafwp
N8UumK7L/MUrXrdC8nWbR1AIfVlex0uVEWzQ0+377+0VrO7m1dch5ErmZHgQYYuojyrfmSxWxo9S
JheCxnkKP87LuIk9PHciH48my3PkniOl+x5DWIaP3dlebferzhXNiTaStazgVc+Iv2B40EfRFr/A
XBUp37OP2abBP254Fmb+c/2EF6D2xNZyB8Q2jlVUJjaW0X4F2Ev8BaQeVEyEReomkfjKIxt9RVd8
3X3aFNhDeLldJJHX1fErnzouoZxiYNlEZ5Um+X1oq2wKMLL9zzQGc6pOtdNQ2JjumK+WGNMOP6/t
cAoO2ItZPQymSISZi2wnQ9Jlhn2esJ/geJP9rB5xznKeuwudTKUVUOfu24yg2mUmPFaytZrDIrPQ
YZm38jCyQdGhU42om5ltdEmY2goWRDU5apybiS4UvrGS+gC8FB35U3MGOCDRMBc8GIiBirZTyM8o
hxPo3tCbYwTDYzbo75SjD/RUYLcqeGjIIryWI7ww0EZazgbawOX5WrjBwzOHI4gCbvUQiIlz79AK
xbIrXvkgt3KpsUFsjtXaAdJIVRfdYj9EzReHXE6RgAAatBwXLTAHCIFAITZ3QSvgZG5lNDkAz0IY
Bqv8bqYR0j/YADx3YhGi3bDgncj0aPROEIFs4dUdzaSGzB0gNoTEttlWd6FporKjUGmXSBsULfYp
v8z56jevl2kRig3eD45Q+f/+EoRCP4ASQN9opNE75FU4DIsLSzQ5kpzpbOh0xAteTWJkasTNZ7pZ
Rr/6PmtcfOfAwEQPOma6j5WN/DEl3ATzi/9t18CsUdH9IuvM90//nLJnTnb/ySPI68K4mmVjHXhT
2czjCY9NZcoMux5E8VcO1PWVX0ILKst8qz9x5neM4Gr3XvqJaKEV3bo5U/HGYdO7tInmaZDb10e3
xubweqI/Q2mu6P+lNQptddWsoSkmQdRQItSTEwCVOw1pIiY452X6DxrXFmKtNNzu5qgRLjf5YHXM
PKQGSoTu6ciCdvMHx7jVkSg50hHgOW3yuNBXzsQYNuTnsa9iod7oOUTqNafidIsdgK+nWfHGV7A8
H/QoXdiiX/nGHLkuyHO0ZW7hsnINfvndgmc5OzL7RSgHwclF0ZkZhMvgyFAHVlIZVAgMkMFIfGW2
nCHvGQkmNZ4EObWRqOOF71Og/TevjTEHxgGjEaDe5CP0kBU1CLMCiYC/16EScMKA9RbnfUdlH8z7
b+Z7/J1mK4nNd9JLKPY7nMym2IX5uBAUmKTwCWtTsLwoczwmR2+GHfP0uSoQ8wB8fEEwaeLmVRoc
/mbv+9lbMOY3rYjQqhY4/cScqCYu0SruZFeVAoTnSyV8YXWcIlioVS7ajsXkkl2YV/EngI0Gfy6s
H23dtPMeyjbbXErh8fxrQtzlYuD80Y49uK1uQgWGnxNG/M6jB6NmCPnFrzgvtOmb4WM13kI6D1wk
x4zTeVaVnw5WhWtgx3xp65+SJMehkhJBbbtQkSvHxDpwmfkkbJeWF7DEK4BzgJwtDfwp8DBnCXaD
Oh1yZGrszyc2tcvfTBymK1QvZf0OhdB4lTXawD+YttxMnJvQYI7BvU6kVVlicB5uHOrPIUP95H+S
o9zLcpyXJX6rLZSeKXSh7Kv7RyFcLoXRJUaEowjPC7e4uHeKh1Ap/7FhJciuMny0PsvgOZbqzGb2
N/Sn7/IwiCu5A3olGJepRchD54GBiQ2bp3UCXHZvxonPOH0ljdQtdWJHV4e8/oNycP5gdhuTFrLu
OC9ScfFyhjEjl0rGjZb4V4OLRl2l5VycT71gFT6ent8nAd3xCEci87y/OCsq4bJnQK1VMcr335Cj
oAP3H4fXCPRzGN324+mHJ/w03LhJMA8oy8KS2C3Vf15wCv5CVwIbnWTjfB9phw6bt2o/4jSf1JVu
AlY2/LcbUU3EVqvCS191wRM7cIP9GT+VssASvGGqABIPMw57A2ETR6u5T44B9Zgyhd+4qRpOWrl1
fKqlUbZ/pY/hGOnG+qcUM0ENrr16p56Kld8Q9zvYz21pheBB2ZLMfATIj+ckb6j8DX8D8t4QvjgZ
Q+3xUyOOPobwwCrM5Afp5TKnsQZrEb0MTyddhtQRIJbqZmVmZNu90jXp9JWsHJsNN5BUGnZOCe8t
Vw1/kSXuaA/AzJFA6WMZ9NVii8nedKJqNjAhVYhIN6K2Xzb1BwXOKtYdW17St669/11wJhm66vR2
gv7LDCik3OCxVB9o+HlcTh9Nj5cweZ5RebjJFyKeFijPBu7l8wKx9pMNNetduPWdkj5U2TDFpwdD
fGjJmUw1m2Y2BR5+t2HkZA1jBIxs5qWep0jCEo85DFnR1sFX+3N7pHWqHtmpRPacdBSt6aAqeULb
0JMvJXfgC1rumVIPnolC04HvmqGcBtwqlCCWK1KCNHfdI0KmwhHUowy+CkfjRiBn+LMXEjN3RTpw
+SMZdLJWnXatPvPs4I5p+tJ4RSJ2pGxvG46OAXWc1fWJcYkcEU5Z8jp2sMKDrQWCq+xk3TrKwp2c
81MYuh8a4xSUmW3BaVDTaAOGWiPeJTnHvyQ3u1t/7ZmjTkNEgpRKNLWdmg/mH4PjaEd1sj2vvj45
pf+5Yv0+hMbgXkgR/tVcQ/ciMqDd6/GHcSKQT25gLbLX7+pRdUNUVwmtaZ3BGcp1TJ4ZZP3eR+j/
wPShgfGVgwPg9sBdpDUr1dl/b1sKRM+cPVFATL47MCgGMZNFkGP0GX1+1yuejSxtpZig6+Bi9C/l
Cz/LAUeQdr4aujmc3yEHsXuR6lIM4Gx1ei/AiHGHmUF165ppmeMIuKqT4nq96quFP8U3dl7BW6K8
Y1xpKYgkdTbMRq/GZO5gwkgsFFo7RoFMjm2AxaF9E+ol1AONo5daXOtn9se1WTfvabSD/WpWIJ8E
dSaIkvm9m23sxxcDdAm/Hs8PJu5BNvJOH/sjKkZ9e48Q9Cn5tN77C1N4A1wDebDITWbu0XecNiHr
ioZdZv2mlpwjvwueCgodXiPlFUQWVXL4TTMKepMw/T63PqyXLcBFVYI4xok6KAZ1cyfo1S1vzxNw
35P59r/cGPuCQe/XfbmO+u0sRvmlEchKCbws7+7TjieJlpUlL9p8qyAz7ws7oJzSMXLAs0xmSobl
WhTs4NCfJdmcjnIPoUEVvkBM6C6kaUU7BD6ntPBLu90+RzY9NFqtIoml5I0dlGcK14mRWB8M1jLv
MFu3/b7RFjRnsTMGdgMFAVU1VbFKm+P1tOQVsgDttJLNZh/e4tIU4dJColm61m+5POGpdors5kGz
p6nZZoyhjaZVl9/0VS4QDOlmliW2ZgIm+kUI7ZQNsE0FPmrz0JsoWQwmITpZjZtfOm5sEqkBgFi4
bEFJ/HPaYeabkb+6KxO6f13dLewboSQATatLiyrvtyB3uKq2O1MyEiytK2xcATGwKDaQ1ffSKvxg
wnr5VYa+3M7EEjZDsq/7tlKMYTXLBmb0SqSaQKu7wFJ75lapcj0nEWL9yN86Tyb07e8yVCpzcfiG
WAyZBlOqPHmfIgfxdC4rBM80uDn5qUoLECnoxC7tG0Z2nbgoGIMejhpXpIumAF/cmHjMEePavoRg
D0aihxetT3kAIEbBAyfc/Cxsu/egBh4Vm8WruaVhd00JQ49zeyfT/444iR7bD2NoQ1CCOY4y3d8j
jisXWvZ3DdYCKAr7uEoQQ7dhH1d70XE7dcUBSjItnCriLveQWK8IJf/7EPQ5XALUn4atgZabvN3Z
O/PLmvmkr+4Ob3VOKd/UdpZAhmXiJy//v50Ti7P69JHf3ihWqMoAJ4MOsh/FGOB7whtYq7psVxEK
qpEMZT1hZECmzVHjbGFYK2+dhNyvxEpL6AU3s9SQSTmOTq3Odaxnw17nj8L0wu9lQ7B18dICSZtA
mVX5SrhyiN55ZgwzhqD7Yc/jacHYpr+seRo1zYvRgsxesSU4o9NojW0PnhOzYxr75flbFHArfBw4
pfA/26gYhiCQqxJM4nEfA+fpRJqGSI1mYGpWsAEr/ljJ1zrGAdSrdlPUnRIRa7wX/IOA/8xikeJ9
hBTw7Ypckrlb/Ov5PFdgeZ/UC9txl3utzvxJEhGnf/0sGk2KxjaSP3qZXKf4u2w+UufMXVsoy477
owCVU5/fG2PfTRZZN5bVwmIOTtgJ+ugBPZtitcochrSzUYblCZtJW9k7hOyzbLaEKg8YyKTowlci
g/+LG2T4+h+AvYOF2R/xfwzH+AwL0P73t0h+JTROr/xVVbYvFxhnWMg7i2RQj52+8FlOzRQbqYd+
VYYFvAvMcbKqcyTR76de2GdILf9n5i/mKPJ1EaWcw2Yv3kSSKDo/xUUE3s1vql/UDdTK9293fIkq
BCLsKOwEQYW/B01j80OrMiUQREYZJ6uKxOY5HUNtpADMscEVhJb/jQdFX0VfwiN7q9J1VVRlZF0b
DSeUIArMnxhvqFUGGWJ9k3rKV/8bZ+t7qMIOqsiJU3ElDpeKnoYVSqazLwfKmFKXljDifasx6skM
iwzkvaAvSJCIBiNIMnXi/DmE2IUe5/UdzaNqRuxiW5MQ3xrOjvW4+iL3vZT7oD3KEqa1ok4MOqQq
oJOD4bzXJ7a0GDXZwiVRn8+qi1UjPAX/5bbmMGVkCYrrw6gBNyQFhJP2HGMGabCR4Vj/im/GUI+6
nbJSs5kqSzhS1ykyHAFFBcSnuMoFVj2vLluQVRZhMefgkoR6k6Z4+16GRWcV9+LR2dbxkIo5yfAP
wzePyfnlyadxB8gVhw0Jv0+pMBGlN+v0Jd5sm2P3VpdkmFHjFXIcWedzuueNliojzLawaAw7uOpQ
QMkSJn1c1nRtU1u8guxMVcsRigsrTfg4nOTjwqq2XTjbdtyHqNfUmCI8IqJDJGHbLpROC8aRjvw9
Qu4aBYIu3bfNRSCWwN24g8zPiz4xk5qR1/buZI6UBbc0ubuCxBT6FTjZLMoGDTPiXWqpyZdpGWq8
GK90FIPvBdvxG0FcajJSuHrB9z4q1Tsyxjsl6JVkTy1H4W6lWh8sodPiL1iQ4gkNlnK0IaYYQsvf
PWPn6JhHDdvK8CwGs+n8FPfMvovPFVQTbj5hfjMsc/BNbPB+q2Rqsn0RLvuQGiglSBlmgPDrHp0e
3PySw6IR0NAvMnq/aN4xP24PTHnbpokLoWPOHu0mF5w97hotg0go1Z9qSlCtMapHxPKjDAqS7A+1
EKZ/an9yLF9ayvY5Un3FWgZRHIy4nWBdinyGwKblnik3dgqhVGxK9hspstt06tMrRF9WP1bVx4Ji
BoSA3Z3OGc5H/oFeRcbNKRXZqN0bBeOeJkmRMkA1qPXXBosN5/htsss1bMRfpkf8PvY7V+GZI5gD
o6YVhso3ta5CTgtBuNB5Q0Khtl9xTNEexYaemJynu5wf5ecKCZmFgRMQmbqpK8ikS9D79AxSmtf6
ycTL/UulTay/7veKRe4D6hdB3ZAIBwRk0uaRhknIdxPybnjq+DPtkHEwWrQIzgJY6uFpfPLU4PtR
mhmiziCMVFwATJthCfYoLMqjxB6h1f+K4X+Rza1gnszDyEkwLlIK+/23sAWRwYWqWKmZHKUqEdu1
wBRCvvkgbeNg8trRHIwF14v+N9j4Eea+YEA6oDF9pxyMIVbCSqih8IAGuFPVMSlRzpBQpKbrx8/2
S/s1/XtuaYi3uj9t0ZB+210uDl75AeO2x5VlhoQz4fASTUjJCdZ3qqv5BAaqfLNZ0aqVJiFfB2qj
3DJY1FiH/rrr7b+Eh3p5Qr83luGvBVgEOhm/kvlsQVjo2Fewdr8AMQaf9f0MgcXkAFprn05pnP3g
pgqQWXA9aOEm7GDjexRhNSMDIIgIo+SZv7YzUZ8DyOWFiRffPmdMdJD5lFK6CEDRJBHLwQ0PYkDS
dLFj+Nu4vuBH4y2lrkkwl1Q8jBhzgB1M7/C66/OgztYXWDVlTKOPBtzbXlYtwHz1/Bre9dIuokZ8
4OR5rACkMjDiXazzOmkr+IeGMEC5qm2Z+420R+LOXJXSY9LA5YKGi+X5DonI+P1i70TgSovJhAuU
TtdItnRw+sTHrY5SFg3UkCI2quL33pgiZejZWgB3E7VVe6WRU7nIabsZPnQ1dWr9BEOBE5lcpzSq
I4gVf3hQfnSABWy+OYnwwPPTSMMHGEkEUT8WiXIharisc1uA4tCnAIpstbxXEQTrEncUdpfeBhIN
5lo3deIpkL6Uv4dXrXHU94ZDIbwPrMFcp0SnVJEmJk5eLGry56bipBp08cxNKuM9Hd7Tg7sETv0A
0ISYNFCbISyudvQwtBAIwPPTYlXl0k1AeOrJDBJZ0sdsz4U+Cf+UAkDuxGdjHH8BPP63aJ1lfCNS
qnl8S7tf3W+famcrKS9+WcnTyEJvmuKNjTPoBr0Wahd3qIkgNc//u2I1AmGgJVPUPpz+qq0qwmxs
Hw/qYEC5fXRwf0hQwCYmlbz2Nkrd6mXdJwnlnH0ruj0TSaTvvpr97MVDwfTmtiRi4AcNT8qJsClg
JcnuX0Ff1AdmJguUvOw+9rJbewSmoMgeZPIVbLQ/NQhqAJxWb24O7kmQfM3JGpeUbuORbPewStOW
rpfy9CGSJoOVf1G8lLZr95De0tqfQTGSC5VHJrOW88VFTHQUH2wGhlNkrgd11aAMZMAoVUpOooBo
di0DK9yHrJZ4JqiYKdf1EYI2zNLtWZKrFmtE4/SG08KBlzDL7SenATqzq1/tfyE11lBcwdpPV7cJ
nVsI0PDxWsqilkUnfr1XQQ6T9u8qZGJV7Dm9EindmDTfwxI4VkaqLcyIs1OasTufBHrdV0bdmWt8
RMG7h2THJK+U3sjJctmSL4KgSsD2aSPy1T1mgemSIlL3Fsk3RLCDKFTbOwyl1J3FNygeAYz13bOk
Ce4vtBrvv3WGdt20gIsf9pVq+ginVF+JeBJy5bVENmClT3fh4bAS7fqGln4PRtysmyYBsMIYlVPq
lLbJGpqEbZeKCkng3CC0Eg/X60O1DtQe9fEw9UMYJGQLTMVZj/UrzLxNq5QCWbZ5qmYUOkGohsVh
+KK/L++fDs5s9r7IsJmxjWwR8xpcQuefvlhqBKeRTeDs/jgwvET5A5c0z6gAvR+rmTIVo/r1CkSU
uMyiDi2y5NfcUAHnLi6kYjcCfcHeMLuTot3CdYURf+Es1XGPjJFuuZ9lQkNATg7K6+M7KwNb2Rtk
I3+zBJvMRjvj+OIqdlAeZXN3c+qGn29fA/WlXYGyKaL81RxhGIUZlwIODR4HC5AAvWsIE0YxW+RG
qCGWG3bAH4beql+nTh2iWBDoXpxrDBz6gvGf2xK9Si8E6GYoTM6b7rvRPaaINvb66HD3ms4e5v30
UOwQqyUnkPy060hc71zVK4MZPM8iseB2MJixcEz8oBcA08I0o338MtUelgtPP5P68BIqsY9vITD4
M6FroqYh/x0F8ozPSW9VPj6vZT1hBOe/p5AoziUCtVd70Jr3Inf+f1xYvUetf5CMuoV27fht/8of
0480MH6a7yvJ0bhgTIvyxhVjA53l7fE+vDJDpg+i2JjK91CieapJv5y2fP2ARZI6VJDIykfEwnCQ
EGzgoY0/HSezfuMVdeTP9cS0cBnBnmqCdnhAZtwDS5J1Sy2b1vi0twHIaNOaB4bipOTUgMeBb6K2
jv3fIwFJ/2XYNslc3tFv6tCb8XzS8AzrxCu2vQD5p5o3XwMQhwpQ76JEhfOzM8sTT4K7H5ZZ8Jzo
uXARQ14Jl8+SHmfH8pG1U/UtCsnRm0Ws61EZuGKPMfJsq1RaDXFdR4P3eGa+7q86d2ycbuzXVhlO
iJ6IgWuy4dKpjjWKTkHxEidKRP3B38cGs+3nlOT/6X6fzpugeUjIEgGv6m9DiLAloegpFSkEgxb4
JHhWYADJIKl5cg7hndm5emxtznfayy8S7nuitkx2xaEKi+bdvYJ0DCOgnKBjDSULowgWYQsHFOP4
hS7WDx75/EuZeQuyj/Er2o2Ifbp9dHM7KmioIMoB5iX9C3i1qflfhtJQnMe2O1hdNI+jrz9UmN6v
VtWMepWfRnW2f4XQ2t1FH+RL4/5Auder2kDFofhDdsRJ2B1M3qN7E/WUtqABVU3uPO7KoK7wvenR
UQ8U5XcsJTz23Ofh4LZ9T7iD/dzWGTCTsMm9A+lhL11B+EeI58851ajZeHDH80B2e0jzCi83hTzR
x7fWau4uidgVlQb/F1RbZPjoFJ2SVPPSi0Qy6qQKvXPFisgw1KS1aTE8SY6oPWNtwSrWdiNabArn
bAp7AgoYVtfHQHgg12DGAGiyf5jlMvmO7bYjfha22r6MNerIKLHjWcEO6ULTsGZQ26ZdagXkQGk7
ndEl9CgrqxcEBEpLuKrf1g+SgmFpVaGzEbQGmkvVk1x6ouoq48rpOvA7xkQnjfr38jIbg9oUKrux
4snozv+tayHjbfEHJfEH8STGG1pWCmkjmzeBzCQxjT2dfaDF1ixeZfsdZ54hNd6znKUBi7xzkmnV
Gw1Znv+oyamrZxX2lyp0kv6vB1m1NtbJnkmLNWvqgSWh6Ep37dxMTFf9d5jW33GPmEbi1QSy+UgM
+GdumigPsJdv92PjTsdBveUL08zB5gathRW+wR0Imr9t3HcIL4jr78/0LOEK7GbfOf4CeHEyIAkY
BunfKSLf13qSOuCb+Pu+ZpseGZUZmgYPpGcwc2AwX8Xxc1gi+htevYIJEYP0TcyyZ6AVywbpVYdb
/6881NNH3rlzR1RqlLi1lYuWtlf6jYFBF/zdq9DHuuP6DtXKy9BZ28MyjvJAHilo1UuMqP+HcTm+
/K6ZUv58ky03QTO76d7YzIZmojrKsjkd9kC5whOfhnYe+iydNoakWDbQXC6Fc1LHSNnITQzqTo28
KnhfGKQZTZlBCplPh7dDqEwD24L0nAovcGwyrMtpW0X+XhAbpS3JVItZmSYbTbFYHSR/5fIYNPFX
rHz0nOjCdqJFuxKjTMqYDxa7KU0xL850dPZ3RbACMEjOmBb4ZOaOM+maHOe+z/c99IDFR7KZc/jH
BFBzgig/C7cFbkC5mzpg/OgK46uxoXMl+FzidoMs3b0/PLbn/GmQWus2xx94mKikZRRBUykrK0AA
HbdcpNchUljbo9lbEJTma3EgGX9tDhn648rch019VOuvmpMLz0wY38xNfwqwC9GYZ9RasqTC0C6v
pcNylQJr+Oe31gONKKxe7NwjEKaX2235CsufcS3TafZlrwmW1nf4hUIaNC35WBHfjMAngxhIMW3k
jTJmRKZFelKviVkeBJQPwbGVRCxkpJGOf/JTlCBya/qHQkRCALKD936j0pYlJQEt4Ib6FRz7x43W
KFsD2vwKojn0+92EVSY9xm9zap7Vp+lSkx2kgmseoBssxAHnw1+0krCSgkZJnO502zg1EZvMsZ94
k11PP1wp5iyEDhCHwVG19B4Kr52VL/Mc5Lrb0fq9ApEkZRdTB0EoBNXU9+R0jyMRVKe+y4sKRCRw
gTgAXPgoWKPJkZkSh6NxyT9/mHw226Xo7J8hU01fnv9gMDxysXZyDgKrmI6FGmS/PNLEDJm+8FIw
K8XKRRfSZwnZ2VYC/+aVu6vZnkSKgRslfE+G/hsnsJMPGnSbO6nSjNUnW4yP/SWQrpZfWk0Kot/b
CCmZYPtEHAJhPk1PKxIOA3LSUexS3JIL9z7Oj5vG1lQDjX6VsIeqBh5ytwWW9hxXVK5PaPePkDO7
vBm3uQQauIoUNJfBQVPMgh+Dcwh+NKdBc9uWnFe26BNwQ1M+imM9hh7neIXzICLhb98wwM7uPCki
LyRRod0pn9Wm6F2rO8stGCMnb6QgvKWLWsLlDR2cRpp6dx5UzH4sbMNyDC+vrPJr/cSH4VsN/Uvq
bCOhGMLjL5E5kn/2hBiKbZCjlpyjeB8GgXKmKI52pdeZO8+vtFJ1voydJjapZMiPTQ5auRO/4yDe
8f63F0LDJRT2ddFtEQF8D3x4oMXH6neHB9m2xkYOty7bCxSL7Crn6YF8BoQrjuvieDOjRjCGJj9e
5n/K0moEYyoFPOegUNXp6y5PLUz9SAjq6ZVtw8rBahI/5eq9bbjy4zS0VSIM36rgo5Ij83cfxhCT
bHvo5R/Ck9TJmhWpC3m2cBsHAq5n8HVyzeScG+rIt4ajxO2WGTX4qcCJCIJKunMRKInq7lulDZgy
SNiG6T9TbfeZBGUQiYxPUc+HVi8VMboMgTSh2oNr6AeYvTEPj/l00uoVYByjLLjx5fRMs/rg/OZd
tI875SrVEhMsKOFp0jBliyNXSUog4O8gt82vrrTq5HLUDYpOfsYyEXxS11OfQ/59hBFWhyZnfFyW
hXPR9gMIPrIUc/IW1Tjkl6W//8SWSrNjdH05TSwPseBsCSXsk65GpU2fW/0CVxuT9Fpkv99X06ff
lAIzZavELiSvVxvdfJcMPAkw2zy7bYitI2HnJnPPDCDw+kOISNOJR3zbk7QlaMZS8q0+d7Q3bH3P
RdmbPFcuckH4LDDCec8gav6401gilm1Z47dy0YuEbykgnkgxZBZ5cFDkLmN51TBzCy1aj2Kx9VOo
UmUU11ohTGeM9Rr7+GLSzFH6/AMDnwlHQKBj9AmPOd6oYBjpI+VIAC9x8JWjt90Q7VPST5qQruev
8+fhb/OyR/g6ZE+Lym1RrhuDnUbrJDxN4ly8Oe3R9XqpqoVr0RUoizAv8sQ6kVZ1AMJ3pcNReT8n
ZnCMERRFUiKFyuPzBmA6f5R7FGdiKo+4xs+0meU4IH/WD2g32W5rDdEA33To6N8VhqKeobPOjaV9
3j47tagTC6URfPKLG2/s4KQpRbpFc9vvv16LIwC/qWR9WXY04/taN9t6I9uOyIJwlizH0kVc+WCB
BzsSALS/QlqleGhBiqxYWLtiO78SayqFjwt9V9YY965E8Uj2UK1GyS3VrY9hP0aL65Syu0YHj8E7
pM7hiE+yDszOgcoeItcz0mvi/cuvmQyOf4mjiaQIwfc2+hDLzIMTDLJ+DvWdeKGWv75qMD6vES02
nI7vY2zYGSCF8sWan3x7zTgdv6n5ClNu6JFbHkUCfE3omi93m4Q5NLTpUKbxkuuLikVRa12Q84wp
LsozAooVllnYx4/n9rIQULQ0zaIU3XzoIZDHUrPXA/UrBOJuWDomAMJEtOiKzglR44CljTrlzmUi
o8b2QWYUMdJpxbmP8S1OuNtbPkFGG+qAJnGyjt7sGbmaNC13u1qw/s6F9tIfhI+juZfqPr7UeyVj
ptpygoCeMo+GDvHFzeNzVYOF+fO558J/7xiLPmOXNDn0Y9m5t4jhmRu8YH/9tFZvBUwCxrYomtcI
YiMe2+bfsSenbv8SFEGXDU4uEt3jEhNx9zBz3+WATLuvMzGH4VGya60oJRS64NYVnZ6OA3wa1mz5
hB+QVNf6Fbhgx0U6/UTiqDtNQh8uv8Ob2dhHrxTOWW00KlbhfCt8zJFeBmH5jeuSZ4ziMXLuyIZR
ZIwTjk7tmQti67rpu5B3hBWfCGPei5QQQBJ9UQnkggNVSaUxCNJPxI8mxEgvsEJQXoYR4Dq5fy8O
UjY6YAV4SqV2q11Parwm8mq/Upx+w7dr7FRkzRSmknDRMT+aVRDgT8AS7ffRrcySOgjAShYyOJLN
7gK5eyLDogdmXnm9yoDF0jg6E84PwiXZNKEoSNAjn8d2krjgczS1LcIBWrP19fS9MKtuB672ZYl1
v0Z7tfQyM7pKNVtELbeAtGtfubyP5XyYsCJbAI66MwzEt5TG0aFe35e4IHJh5FhMGo646M/r625H
9522/5J1Wef9pUE7WFPc8o91ZUF9VFtE9oSoFICC/VLEiuRhkNCfBaZkassdy+Y/TuoLztn5egdR
TEIEdhzHf5+0JC3H4TWoTWtVagBh/J1BqV4BYSZNfZO4izz4XzklYhiWyDyKu/nXiOV4q+J++tkQ
9Gh0O4Mc2iQW15mBuYekASW32gpMWfspSLR4acqM7vg9xGhQUpoJPJJkD8rEPjJbaSWeHw4IfzeW
OJP1U6xNsuDDU02NIjMRe2kz1E9py5nJnCgPqm+ot5bqQ0aPrkx0oGCLNWJFrhBQSfNqeOi/YOVE
ceOe0PoTJ7IGts0OftSCLAbxHodb9ytLnlTJfgHy37wu6NktuE9tXv0WyYo0x67Yg0Uu4RLSTVq9
TlDyq2nlhtK9LWvFVd1hy3ptEkOrU4MVZOGOYdoAu8WAdoLZYdYreZSXLEkwre0Xpz5ltYjGiycG
6h50OIl0QeFj0B+GNO4ql+sEPARSRWW0NVA+Z8/6RQ47RsHPLX+bs+wRehAfezvvC3UQT5nHAAHC
Tr1keYyLgHfRBDOjyeVxkPUl7gWRSFZ/dp3K7NNkMererDJT7+m681jqVaaD2CzZQ6cxGoBHSFSa
vgY6tyQPfZt1Ghpb3ahRb5fwoncx7iKJsLCTPGgfatAArerOWMpYJ/ebmAQxUxQup5UYk2zTrLL8
ws/sdUAeOxYquFsFV0YbAC8s2EMJ4sZoCefH8a09V99qvECZvLfsl0dkWnOUeFwfiCG1jzBg9CLb
VvDvdvaSl31jT9Arr1UDCGNI5OCFEiW/HSEEak/AbFKvSH2UpAJeMZ1yVvYTOK3Tg/Exxqy2WimG
Er37WXCFnl1GYNKQ3f4jAYzkXwMDQD5Hj6EyZOsO+kE4ScjZDickjQ7+r/FqynoBvC9qWBh+4TK5
q6a/9teWFgLnQYcqyt39Y41sf0KPkxup7jdPpnXcSiU5MIovVZkMkeEDaRao7kZdKcFaKVFsJPjr
fcRlp+g9f69KJzAf1Ut0jqFTyrxbfoRjRBSas579CiK6OAWo0KERZ9j03TTlef8cruYK+n+bJjVl
0dxq93LuRBejHnE5z2eT46h1hEGgFZjJCkQqLEjwY0Am1+o3wNP4ScfFXAtFCsnoC582FA5JH5YN
5x5t7lKGkUi5JKN9N2jh92sdv7amDuvsYMRth1aud9h7lUk/XXB9xrp0fytVuDL4wGcFqYElCedl
pxUB5Bd6sXKCMnEPMEmYhtDFYeRDcdzoO2IUdtK0e//Unu04sot8aSEqO7Gk3UDvv/sSyM9moKxj
dHMb3v1z91r3DASqIaYe6+R9U9APTOloQ6kesIuDQFIJrivTjKrDUZVbrAC5GTtq0Zt4icgVwATd
GvhMFioFJZOTy+/eBrFBU93m6vgk+ZVAKviR4hGl0FlW2qKQncCNqYIkn0sTfFfe3wlsOsOJoLr/
DHPiXfveSqV+7d/qP5+ICc0zUlT9JqAHfdgYODxttCuvtXEc+VMFlv9TFzfejVH5NUKSupe6Q6IM
v7revwbGJse0WQrgv6hpyRXeLHUoi/EdZ8FCex01QCMU43GnXAVE3qkoUyeCT3mxYIZ/1VeWDqWZ
eUEUPwggl2Q4AsWA0sfL4I3iGEwMLNS0mosdYOCf7CmNtdO11VWxUN4W298Z/VQhw3PBFN0w/5LG
IuQV6QQkUo1ICTmlALPjSxKZjmfbrHR+8F8cLQfde9cwLcqQT918mVvgq8BbFrTtAGptSabzQWHe
7570eDU0thfvFc5NxZc40SgX0WO0699T8I0JE/TlI02TgLxb+WaTOUzK0qOuc0/EgdFw0IBWEWRG
++nx7x39VS7DKlF6AiNU+u83VtAtNGQm3wDFkl+SPkuvxau+e/s57MnqqfY/NxtiS2/PR19slSaD
DJdh4ozQGI6a3psMAReFp7OiSxx8MGVwdbwU4HojmzlrR2Pv70Jakw7KOuhK1Z6JnccjWbM3YhTy
cZneHpsR8ZjqF4HuuTKxASa7D/1m51KISe0P0H86KHFOp0lNt+Yz6hof0dQ1TkqthYaHwq0MB6mL
b81dk0ow9OO8jXhLkai47gf1Cz5pSZ3pxLGmvOFO7oxYZ1KvFHig5PGcFKeUwyBMKOzbpWa2DSeK
ib2TC43pH4OHsUiryecOlhWBCx/b1t6P+4XysWe7Rrg5LaUuex0/tIE0/qVDQxPEqFasczqQzxSH
+YfcYhRKx5ukB3Beuby8K3MhqWo93i4a4bpaQW0WcQulZRTy3gQ3LvzToPA23/71eloxGxcwtO4Y
/tOIIwJgEBE2+LEtEQAIz7wpUjxcYTmCratVbngB53bsUcaVr43nMQzDDiYIqJkeTU3mQJEVH6Hp
9ga4o+4+tpNZGndmWEqIaMJ6gz4vMXeLkQ0JD3bo1RgOeBrrsYXAtR+QiQvN3R9gSfPeValLt/08
+yGubMp36r1wcBoJlQ1PzPFjszGLcJ1mu459IzRfOUkygUoCPTb8aGoylhwltyQd9InBLm+hhi0g
uZiMiw0yR0zS761LUlkrkV6MxlVdljIY1HllkUBvddhwkz3qjtUaFF+OdtukzXkE1E84GScthzer
hPq+Jsmgmx/gNlvCh1sXKucJIpSd4Hq9qnfRHom7DqDu3GnJxvF2sjto6y/3tn6miMzcMijcdq+2
+w8XSLAN2Hw37aMFtzMXi7NJ+yCXypdu0gmS3g0T/GkCn11lH9bUjiJaxuzpcV6KOKkpAehUeyBK
yuXv4m3terfN1oitdtevHHbveTZmOpj6onaiEKa8ozgvJpDySIja/L1hafhkavF5S927pNFCsfnX
+3urAwjFMWVAfdbCX2bBMMsXWN8neivRHE1PfptVGOn2REKCG+U07kqP7NdCcCWtDuRGNTLNBrpV
UekM/vi1y6lNUhiNkYAX/7JV0pbLDpS02ucz1TUzRTG5MsZGsPBSEN7sRE0WraGy5f2Vvl7xB9+E
tnA9EXyRrK2LEjKX/igqA9wPUFm6jx1W7AN0/VKWjrCtLpGdPbMniCf6P9BeUD+DFJX1lCeBj7Cv
MUvUWQ/1aF6ciB8vSLvfSwklvuKe6lzeK3CoK4ScfgwEan+en5YJut/HCF1wNiH5nhanpMTthCTr
Foqqr7akmDhwh1RvK4KH2Xdq+3MatXSwuOkM4Jc4j/MsoGbHWH4Tdg3/k4/MEn/dDqNZwkt+gfAH
TiokaYnmp5P1Nt20U0OmVykYZXwqM+ePXmzRaDuYZt4i+zvO0i2eyB2SHS81f3Lv+7cUElRZvAZV
J1/2Zvi1ilLMbUhGo4JGD7bXpYOe21wJMPnN/ppy8bIELCmnAZbZqOHpOaRHM5QFjZw3yK/bX0io
oUPvHkzTQkeSUoZZnMU9mbW0z3JZCn9mtH5ZpfJf07AjyIqPAiy0+XrF/eHEO1DXonVdWgME4xV+
47igVIYCLgYzSXnnU394ivRuBZm0ngU03QXJHElgo+9A2GZiOGZZdjqcDvEGShKheSdrifcvKqhY
9/526Gj9haWO4VpLKP2k/sMcogp0tkbyTCVpMju2mpNaN3dgM/4bpxygF+zl+Uk0TVVHAWEYSG7l
i/CwogitwX8OL8hpRtaBfrsMKji5fdkD3QuNPq9NavhPZKeBagFipO/sOLi8Vcz2yyWk6mdGdyh0
S3sJEZeZt/NkCjXh3M2KhjfqNF8D2I+trLOYDik4A3t7DfLlIN3cocSBZwuyWNuKG9tjY+SugWjg
cilnJB6xIGWDijWafLRE26CjQGLNddUX5TRQzYZvzy5ZYKgayGDEHp/XZbfF8PT2fHJcz1KSTEhE
4wq4jEU9jDutfqWJNMyvY68XpFKMxy3TQP6MJl9793hWS2AZhn03i5ScFHpL/2iTksPYqny2Zh7f
gkZqPh4VQbYDEUOZJTfJI/NDvltOFNzP/KprSi72v68zUIN5ci3b1L3gr06FgoARy2e7ZIexeZX6
+MVCCmwKDb/WpeXCqgG1VMMTA2GhGi9CTtT6VfhLb+YVN8VjOs+QnOWGdUdgcFEBISR5YIr4AdqT
0KFtU/Kqkgv6LdA4+4MMR8BMV/YKjXqj5awkS8tuCZRMZthdGPg6ASCVHWYYoeWq8UBMI9p4DU0c
Xryu7nvSvVth/lQuDf7/WzM4N9hC301w5Qq9s5+TyOhaNbGvkU5fAPXKcDTUM1IqK+QoD61zpS1L
JSaqJS6Fg7WIrB/2RGP8bhsP30uzGXCPMcp+aQJuCmzIeShdVYIgpkTnHwa+nakRsraggU0K08Oc
r4pqc5+w1F0qJEvmIYFBxdq5jlT5peb08BGK57tUZiuyjcpcNb89W0iA8o7yDfP+YEehHXUbb/Th
scATd6V0EqVS/KIERDx6PMZeS9MlyOcGt6WCI9GZ12j/57wAJyouOl/ZbGXe5ZcjtPTv3bf9ZrbB
gLNGkFB/qkT3ZFCj9pUqlb7hfFuYzRrPHBQKy4o2bpwryjk+8Zwz0Jslo/QY5faSZMfchn/mb7gI
+WugHMKgHNtWyFuSKpeFbAHOnby4KgyXwrF7TxyhzcZ6zLe75xrDaw/0xz4w7bngycUi+Rw24M6O
vUt7PIABo0V5ZMIMJSIbpLxUqCUMFsKFWC7xi9RBGW7fzmJ6wbxb5WxMmKIEgS3F0fDdQMPpS6CX
QyAJ1Zo7z0IjU9G3uhbEGVPuUQUrySX7tKnzaYO779ZK8L/VRHyCDjCr4aSIPiiE8HZjR9/d/ZF3
VEtzbW6Z+/WE+/4VLI8Ri9qd5N/wdyfnv6QLUTcN2XuGnb52pn3c18JfFXkfwZhVcT2evZjTn0tb
8I697iH0tlmeum5RgNqwO5dr2S2mjBtOuYAynXR7gM7dvBBKnu7mbIpWT6OWdSvjxkV0fvM1Ph9a
s+6Wpel4v6xpBYWTIEWHSUr5ZL+Veb6W7CCNYXtqBfsgNvowf1IosuStUIoGFVwwzbpThTRJP/go
0Himxobh0Dl7I+dHK+owRx9sXv1Y3YdHYyjiJ5wcM+Q6VgQO53WM1/VPPVufXRFArV5dH22oI8i6
0FJAFGZzy+HZRXw2ilB7B8FenVOpBHRbqVjEs2sno6fSlyBmtJnzZCTlBalJFbWIrTsxYt8SNDUh
Oy4zvP9eF/VgOuB0i3c1LXePQ+FTgVqpRvzE/T23CZXMHJByQOR7T36JZ+P5tXI/mnJOI2sFlqcv
3cyPo/QLfeUHPVWI68J6f264ib8b6MveqmSvIxZkL6cDzN2YgDvWpFT2qlWivWPQy47tdrezm5O+
t+1ke/iRr/aaqIrf31G/HwhXtEFN8WM6qYtoK1gBIfFJ/ctfcArGyq4GQzlVtYyz0Lu0gyN3cabn
+UVhdeijoBs6Vw4X4b9mofymZuLkwaZM0P8l+LTrbQh4ympIlGqMGpHflLW/Cp+rtB6RqC0QbmXr
HszEN2GJQawsc7UP59mmwCACzLaDh19pMhU3LXtKUMcYWNgFiO7U61YXrwZezuYCZfnrQWji8XCy
ZkSIKPRS7BuSubP1D2b/75gGIMPf06K/5Vh4lCZ/SITN9DqwAynk9NAZKrJIjXjPgOOWf6TBBhF4
pBAH5JSypuUW0crq1QPeAlQo4W8ESgmFuCU1aWcTVbWjofqPPwLcGfK4N2rqGxolZ/ZZxc8BJRKv
n7zYNGlOcSSnit9KaZc50WUUIJNVK0fHnTyTVCDEsK91NKpBKoQeqoOYX/pWAmaobrAPBItnd5K8
4FNaOZgBTcghlHzR0LLqoLK44SSUfuFu1GxILMyvXs8za7iaDFUnyNrL4sSQsioChHlzgSXBRvnX
BFlkvrorwHYrcFJq4QB0Nkt0K6+W7rQMiazopItRQ5jxqnr6SXPI45ARp2C+lQbp7tl06vhFYzIk
JvMlThGF+7eY2fOf5p1e2wsuM/m9wreDBx7GLEVY2GmYMVd7lWJFUN7c7TcZx7DENXpUaIdAJoyW
DLm7q7URM76UskQ11YDRdmAGbNIpC/uTr6ODEuaJRcXAm72Y2h44emMb89lM8ZHyE4S0xiHussyq
c1t4BgZQzZlBuaR/0w62iBclUrQlnAY4WqhWo+F5MEg9wwWXgC+D6mIqSqrFZPK1LwRcEbD4tvtH
2NMZLHuhD+8B44PO5SI7Vs9NcG/nvvlynI39wACtIOzwNpUmzBdt3ULTscqE81b+Qz/HObzPHsyG
z6s9jIFEPCfkMI1I4DBEH/KAj+3ZYiZ1g9NJnzJv3lSfNWQF2OPKaHGdqVgl2FIQ2h/DGmDm7k4h
NGZ8TAiUNmRZlIRKZKzUGYeQ6/oV3763Xw5BcfJuJqxmAfTCFH2JRFLemNUHb/ncn0J+7n7Dwuje
5+Db1zDLtUvUaIf4A8l9GVXhljJwGaGjNo2hW00tMhtSdyR5i/SUWxCYJ375hUKnXCKgF30wuat2
IM5SpurFVrtIyTek7HHCr9tzWKALMmMT9WkJF/stW3eAh03hD7gKsglNmWZr5JmO1YLGqinqOknN
YcEFkJjK+MGedQYF6ePWT3XB/S8aFWoYPeshDqVqVBadyJZcqqZlHM4FrySa/IlsqLFHe7SiXI7l
zVRCbp6obS8+TblVYYbGN/cYRzxUikNHZ+aJKIVN8G05RKRNazTjYLPuUWZqQDmPQEpave5eP1yS
HC6eVd5htdm7aZ6FtEfEQMkqq54LMG1BtKjI5CvI9ByrQ6UCA9fljuRuwT2GHTkOQU0VuWJsZ5kL
h8SemhBrORuUrieWGxn8Qgrj+UROY8YvdnBtTemoHkg/Apmj+njcLdqDnAVoK97wX+1CUBIlbC6p
YpWiZNM3CWsBa+5bdhJsFpmi76pUfV7NZwFROw9Bp3YuKbQlj43du0zjQVl0o+wZAvEOFG6BbOP5
W0zlfOwrUQp1sSYXDZeMEhrqpHzagYX5pV7N+ZWdpZ+s3ClaO4Fnn4P3F9V8EwvLxAVc1eWeVHhH
eCiOT7ucyKrZ+vWUClpDyXHpyUTOI3hq+bTjzlNz5z2KHpyJ9EtOCmLhUkLNM8QfS7BLXxJvK4tt
8H/+sPjPC6mWQ/Y0n0Z2gGO3eZaKyE8jEa9SJmGhMB+IrXVqQiBDISVWd24QluRsmAmS/L1KqGw6
YAaqzEUGpd7S2yinX4jwWqubGTMfPxcsTzoazRySKI3xnQFcm+UOKL7qtCDz0U5LFwtRMad+C2jz
OECvIx/OnRcVGW+AaYdKznfyPggBbuDn1WNl7XeFqmnungPgsJmx2ZydUNri8qAcn8QCNWkqd2Di
+0Z+BsFOyXM5gCOfsoko+vvQVxfMM10NSp9mohGT6BaxTCWd4rT9CVJu/npFEVFrjU/Pv6vg/XiG
YZFTLAQIXwyOAVUuaj0RdcY6e34qYwb9WNSwmEazVj8jAB567ew1yok+gCc7j0RhLSX0Qh9/ivUw
fPn3zRDwi54afYF7VSD/tlzKum02Yf6VRkwso7xOpFjh1Q0npaXlZ4ZlIqpz40ajjHErT6gv/BQm
JAs8msM2IKK25jYUTxCSh2AQt3w8EP7rP5Z+UEv4Rw1o6noKSv4k59PhqP0AQGqVJ89N1ToOAHkq
UJaD/sAI1h+CJM+3Xeo7+6oVZb8E2oMTYIp+GQdWPjCyZtumIltpXcI0qw2ANZirpx11JApQwLID
2y1iB54A2d3zmECe7X5LG9ah0NGglYvkL1w0bSzYcAW/DP3vx5uMkel5YhW29mQxtTL3uMpq28gZ
DPkTtK+0tkpiPVMKyqBhaH6W5HBWisMzpRjousLRdxaQujQFK2OVayZz+CGZrG8fMvmN8gqVyYme
PZ4I7CbEo4uHhSr8wLaIMuacOqWi1YJ4kcAtf6LY0+zEsvcbpCZjfUBFoSIF11GIjAsAJEBjOdob
SqELQ4o5YtrSqDt9aXFKgAi10UagyQPkR2yhPKyeWnmOi6Ho5oNIteucUomqrLFP242Y4SsIgBIL
HjezJ+L6JbJrgpzmVyZcVSjKn5mX2uIXw4CV/LXExHJ/cf9awVYn1l+7SjNGVZggfmrmqVcaXql1
30VUVyNQ/JZF+MB+MRO1Efhrn0cX0gTE6xEOo8TPXD0EMhpdocE5956+D+d1wIBLSWmjvLwIfhde
f/pveYCSD88Ysk8ed17rn0W8qsQzvP0VbiaxVDu2oF/7BXiFAYW/367p5vbYsYERyV3rcm6ROeRX
KDNHXENIycixcq362YEdgK/54Fz9ptWrvr1zwjKt8i6dBOnblIuU0lnP14rxolr2iC9d/+WJ2T+1
vziRk3Jf4blIb+SqZh/XHPtamULtELUQmCKNHDCihdBuwhZiFC7pxixokVBoFt6hz8QdAShOyTKB
NEhtFsTDC0iAZSnP9A4XYtW9zfaGvB6B40r0ixebSVglSX+mUTIi5U+Y1w52H9/DKHz37R8NFLzm
hDT5T3lsW9Pl7QTL0pjTE0llDo+4qjYv3gUEvvQa6fFctHauTvLpgFi847QvCCPpVqq0bjWnbATE
DSTJetiVRBKmuyVN/9qgSUnmKX5zGDLDBbXbyDbzLjLjW1GTCnZUVXHfj7lKfdAM1H3yU9UN4kBA
NwophkIUMsMXAHscGRCT5R4IWAHXaabf4dbOobds/sUssBGwzP+aBHm9ASJAM/FJaFVn5zWVDlsz
gwUJex0yDGQ3Rnvctvy+bR+B0aUT1jdg9nfZS/r1zDpTe41BkmCZ957EyF/5VLoZh+fZ73MJqX66
0Mb/wDO/uCbzziE0wxNaJ1hZARCMF2KLNZNpEqFLLKA2TvgSlAOaA6vJi1EOww6QTAc5aQDtoEeX
bqFYu4+0P5QDJ7YDwznq+ZVP5CNx86riXqEc15f+10j8pX8tjJ9F0vnsA35c8bjDPZhcVe53WfQh
KOKB6mkj80BiqMBA5IFPrOLVIop68LtCFZSNa1l5qtY7VMenowzJAMyudf84TcLGTXNU7s+nVj3x
10E7El+Wyg0umumdKxzLhP7AHpbJrqtyDscC5UcDekfyZPYP8qV78QdRABmVJmUYHjw8MKQJ+tvw
PLxjBwoVXSqP81dBnt7MVnW7KPDf3h/sfy3d1h8Y7pre7gZ4KafOA8BSD1Ho5br31aZMnc3gxIMp
yKIKApJVshmAa5M5ldqEP8cq2i63V+vGXCsifYt+pJEEDhZupGYNhOE2Z+RHjkoMUxPaqRrqvCkK
NzuMQfySqEyw4b0e5A/myFHCqyTxA9Y1KwIcIYyhHVVfiLbDmh/4uDlrUD0Ay/v57C81IVsSvzyb
V/f5ilAxKI1YmxhoKWbVBklCjiY4fQmoqEHgIf4YuAnOWwIwohI/e5lgQbx8mTjJNaZpspIgKaA8
58cMZmbI/MKUwDnhDj4tuCNlBZRIYwWOL4m3meM/1AW/+vusw+Avot+YZdPCdyaoykyEXaDhWiEi
W+pZ60KKKQo7dm0s56paZLkzHwgD4cTOxQzylQxTJyAruVaRR15H0C3GayrxE7oFr6E1tiaxqFhB
WZQXh2VnGBroqjrP92cdgleRcrJcKT2wtOkAEnUkEqKiTAUGD+FinzKBcB87PYGpP+cRGy/G2Xrg
7K2xiT62OeCP+b1hEFSw/58zC9NkphuAbk7fYvYEC94wOkAHegOKjM5HRog0mmM8vY7dj/q/oXJ/
qq550sXgipHdHbgnJ91E+82Ejnw3y0MvvDAVdrTTbZADk1QpqCCtiugUx8xPhhuPs5rjuodJaLZ9
lpA6fjBkGZT8mtie394keRByGxZsX+xAtxxJF7P3Rc8KwJoFhFjqOOJj6qG52CoKQ/ju3uawOKWA
yYv8lPQ5un+s4ed4HkwTLPSrHDa1b+gdGOQJDfpiajpDKjsedIQ9HCXOqiblYzwzVpSFbB5yGzqk
t36xJtoclYzrjapN4XGppPxypY/iQodLDdyqxQOy0twQa/nezOkA2XplV42YQWcwqvxIha7A9LyI
AN64CXP1xjvvS7dRlhkS6vgotNLtr5pEqp75OnbMMNsmb1o0y5ZucX2t4muHLvNn8hoAw8rdLztt
3hd6a7YTRh0aOgGxMVLeepLd+3zZBz8aFYKZfHrLauvdYPyIRoBBmWVQZ/vHbFPw8uKKXFpPH/zn
5tM/yN4NbxPvrjtJXhj9541j9V18JTX83OHA83MeFkvJR3KKUq4sqpxjHQPZJz6tUFq0lGL8d9Y2
tVXu16h1yzaGYCBmmjcKJ3+FIWsFGT4AnW5wn2GOys7ryWB0p++iTrG7in/M2t1tBCPwov3cQ4fo
Fmqq4wYcdPfhZD19x679ev6AQlnSeei4im8hRe7sBvESvPWkWYRTl6f6a1Kiga4Cg4p1AvUSDSJ3
7FpNySakujuYObIGbXCRYc29Dhu5Z4NQfZQHNuqfbRkvUPocLxV6e5csYyME1LD6h4c2MPNC57kM
ZgItBKkTiibA0X/1WNYQZ6PrLTqlWz5PSSSsMP81NQdZpDHwzxj+s1hpSopmY8fgtuivH8pSowv/
85w8ylHf3XyFw6HBHc2NIFFdshALNkXdrYxVCKCg1OY/rfbiW7lAgDHpVjrrLDfPRDq55bfOAITs
wewqMv+CCvzxij+XZSBnHTRBRljMXWWKALtHWvcXj++5+ESg/yU83vo2wsEh0jUQpg9hHzsYfNBW
DWwrCIj/6Nhpyk7NlAe7RY4tYNGE4jRBAPAVWRua7MFuh31swaEGPx1RB+BsnnxnTtMSKtEvE9Pg
Ycj+BpZeHjt3KPOfm9abu0sgfR2suuB98fH0BE7F7NT96pllIeS0GMS4/gle2t3vnuX6fszhvjdT
tGBwpdBCZC2aqPzpAfDHsxKA47511S4irgkO4+cJHEVDJyvNOvEGRXFUr9wrfk8nA1DKckQd34Gr
13Q3NMtuJtVtXTl4OP8cOUOwK2h/OGNYsytaOv5192Z0JYPPVtHhje1P3ilBm4wh5Us26DfXK38+
JacBpWwK3FscrJDvgXIESWo0m2H3MvOzcuXQK7z3ior1JOllGNgLCwpkUXYFubCZ7wkWejdej1y2
nD158oUf4c5kxsHHyIE7e0ZmpouNKK7ns83p9c+QZTaneakzpKJ8HRVvLgkTQiwUAXgJ+HNXXfNC
lLZ67hXWO2jMRLacpxL3rJqk3zBIZrhwqb+tKEeVpQekUDFpunbQ5s1g5/DjRwMUQnYC2oZIfTo5
xjbQWZapnXzBlthWBOswEHjUmuJmIz8p6/aYLlbX71BKWBPLGpXQyO9B/hGVwAJjSVG9PgvqAMZd
ZCCSFINl2jjW5nyLEMgl6zr0nJmLILaRWnYoGOPyUX7TnahS9YWYQ1vcqifGEtezmFt+O7L23qyi
dh1b7baQtc+nmtyjnrqsNB+Ep03qR62o1bhzbNEyiV+gvVeDEySxpzU6qz3FBRL1nCz0E7hlgz23
pO+PZroLAKNR7LToZgF6TcU+FZR1Esj0NLsm/P1wvfEIvzGpCWr0AnozsouNOGz/8EiL5RQVpcxO
Y5vI9/ycyYruMXYXwpzYUYdJ9W8zdES1cS7WyJLvENRhl59MwRiZwZd+Aq5x4AYfU6+ixs6nG6uf
WPilSpnpqZDw58kTeOS7O4pWdcXNqlFRQ1ZqgspaEKXDF0zykJ3O+uilU5heaku0I3QDjShqPkk8
wwrijpu4f+dsUTGKAfR5/pMuFr+yFS2hHMgGsD4Eqcf9ZH5LMHq2H/el5xoHr+0I3sYfIwaDQeW5
4FhuOcCGg/G40Pc5uMsjOlROkAvm67bQtUBKwoUfAF5NwLqi4FeVhhqPuSPtWRpjqF8RSUSZquwB
H4sCMjKr7j9P2HkuVMrrlvwCoZaRhqna3+gTKKdj5nfF47gAsKfbiuggn/BSXuRPEB6G65/i2/25
GkgY19wrO3f2NlxAYcGy3A2TJ6fTA3oEs0Cjdm7Dt8kfHQQWky9xKTxdJZO/W92LqdgkXq8+wOOX
9HOBTDmc7W/cHJZ6hapIS8IWagjbuv6RQD2nsXST7LFnbQsljB9SIXa5898U2Fc8UBpoi6G2yvAL
/sfpufzG7iUEeqMvpvWWN7J4+JD2cGmwenxK8gzXs7yHSBG/O28wIKKH9351MQl2f+EIuzMefuoo
2asR+qs1qJUf25Lq8Lb6ewBM6dTpjO+KqziNU1zk6g+h5NRSDLZ2bgkgFTCNrU3UPPl48MFm2Nhv
hU14POunco6Ys9H+aOCQy3c4gOl0lI6ABfA4/xSp8FYhwda5Osp+pSnCL4pefSxwLaEHf4dceVTX
/PZ5yph8xQNwCJFDTcU2wVSyKkR750C0W2CDyEKXslnJa36T32i3b8HkjTb4WkUttnVilOFhwFHY
5aHeBOw8rystUZanxCdkcE+o3kbJDeBVAzuvpRt2/EqoBbS6+A5jZyS7xi33UP4Uj/UW2KXMJW5/
d7yoE391WeDuVJ6NcRldF8ZL3JIRoWAO9j1FcprHGDKPQqCBEHlCPO4MYdU2Oo/wStGRcCMm5CMH
7TZo4d3cyURdI7FCBYx4n55u8ugI9kKghRTwGTZkdf3YFlpGA9SuCfi5hDF8RhjIK7z00giT88hR
ARaQg/SE1eXe7xOcyhGmqyYHm6FXrQACu2vu7WeSMpoBM4rCM7LoyxDbAQh6iIzKo5LR+muhqZqK
mo/IXFosRriHMqMF6gZGuc3xD5NB+rhsJ49P5pdhefnQ4krw6g1/8eAQs9+UZbhj3J/qyKHQ85Sy
BIDtuHT6fBVwbTxR8Lew5VEyxOgS8QEg2Fke86KNna3yQQyxoqaVcFyvOQYmm0u2cRORjXz/TrJP
c7jWRMckz3CgtoL2XmL8USyKfCAnT7aZNNTInwp7u1Mq37CXevyOdvPENWkWt285knSUKQMs+piv
dJSQH64MeP3xACi1lZpu2ZwtlshVbw4fVA1p0C4FKq/9ILVak2p9F7TORQe49Plk9d2YSlhHfxWm
Pa/L+GsG/yBvG5K+FhHuocueG9ExkUUNg/cRjGaSUyJttJc0Ys8s96vx070LMFr1grVRDYh3LLnj
hCgqJHF0n+cE0zxo06jG3sQjqHqJ7vZnCyhQW8xD6J/XltbGkuu4SQ8k96j86ZrcxBxbh7zqUpoG
0H7k9ysdaT5XVjCT6PMS97VPHkLNzNm3guA7zuA2kQ1nbFCdRz1PWaxm3trnk5v8VY5qIR6Zp2xK
DYQB6ZdAXTM+LGa6HiRXqFukVLD0J9nluZMHZYwMVvhaBxJJaKqprw72ZGXrkU4PN10aGz8n7CMX
O0GGIlXLpLg3PGn3PND5PMTXvbSTrJJ4UsQdu3nZek8Fzrc2PQmFqKCx5SolJ+sQN8VjXxRuI4Vq
o7iSIVsdfLbmBAD/pLqyUSuoETMNLa6KpZFbfUGeRcZi16rbWEqjEj9zRm+iWJY5gLyDCe/M8vaF
zxGyPGyA+7X1/u/vFhxQ4LeVW6sMOO5NlGCsWllnRCSyKQxey5QS7AP/Alv7z89w6uZ/aoAc46gC
yB7yF+Almwk69Lsu+igGleuZGJ+hQ+oYkfAu1KqXmECZAq4ZU+rakPBgcl8jTD2r19mP7pTccSVX
2s/KfoyXFzWy99KICC13e5fAtyP/wzhF/ZFJXpLZIumbnfIYrLixO9poNXlNiBMX+TCiz/hhgSaX
uo7brAek30Ni5iAqiJL9nl5NT8WD7FY7qEIH+LJbJWmcjjevFAAtWhKa1wMzc7ZDvG++smeYjZLk
liZzeO0T5rbk7KpsBK0ohmj/naasPeoWCuc2GXeHFnaWco4xtaUta/QTPwjd7LioohfctDA8Crzi
wyDXzRlCA5pR1qje0VmjV5SDgEeAYzqGKucX1redDrHBb2KEAWdWlT6UsmUE1FEUVyqMkeZhTbj0
xx/6OYj69F3cGfHERQMwavCo2hCymidVGkjuXTZvn7b5aY04WXSxhAkIQ76EUa7Otb1Cp5Q2nB0k
o3diDa1MtvGBPiByPrIt5I/Jo1YfPws0Z2R/pxpZUhNpWvMgM/k9cKpWQuayQ8TFygFKneZUyF5+
Llsq6X9nGk0+T67w4XL4OyXIZap1vr46v4Rvr0uKUckXRWPG+hsLEUoRwI05Akb1Qi8YUFlDnOMJ
dK0JynuQUv2owooE8FcJDbBIZVsau9K/BrwfvUUj5to4VN6dLnfBmi7FJGHWT9kwaFNRkScWWN78
hyPYYZ7OfXMGfB7maA77Rquj73SV0PNYyHlZVuuEPbteh3ZpzfNNoOQhyuHcC1t/2Fik02OL0Erk
5KWqjctomQWs6D3sVfOY7uewiUqx58r0e91qBxZQyfjTx8ttTRavoUqcmJKcY1hfMRt1Ii7uS5cr
+ONBJGYukRt68aZGAnTcJbfcYsrcDAL2eSATjUz78AJWptTbnNwzYhMTHV8uz2SzuMMVrPQ3NIHO
wpUZds0Md88adTN9TvcP4t9BRuCj5XIFkfcS/Op50G2F3v/KNyknDV6uCpCbNx2rgPO5gwOLSKME
N4iG5tcQlMLat5nI/lg2ZYusFNmfFmvbHPPMITA8umYhDS32JQkr3dCnYHLGTxIFdRIPejKVw087
OD+sKDPFsFeTz30t3ucNUS552Qxfx9CHSV5PWsNl6YqLNL/ljgTEPi5zlBljV12xP4UtX0YiQQFF
yRZMWnE7inKIXzfqce7P6zt7o0boca5ISBR39I6jPfzdqchjkWJDxhGtDwoqLDXhoeu8aykQ2+OW
Gl9Bj/2DgVsRSNpLiDv0hPLE6Qr/VZaQW74DbUWIMDupJMZi84qnogi3JktT32XaLyNNDFuDWK60
CRz9VZ4uN9HFchYn4av2v+shAoUtIYmwx/YzGwKIG0M3Yx/+alwspGR7PHxROCvKH06QDEtvJDSX
VQ9QXx7m64SsrihcOoGaT38ovFSZNd0cSQ9ZjQOCZ6vIAKt/8Yb+G5t+kZGxQbijhA9aTcbd+4Qr
dojW4d9UWy+CpjxTsTUN+u+mJZD8BO2y9kG/uIEi5xQwIhRyTd+XDlmf/prLoWRe+9e9HEXj7bWz
dB7FrNpWueuSvEbM2MNTYgufJJHxSR8JKcJbMGjIX3b1uwbbkO3xXG/J/7Sf6Ve6ioevfilWZHQz
ebOlkZoGOcXXXaqAbHW9++fa+UTmSbue6Uo/WaGK2pBE2tck0RvbsHzsADbOOxgd9HAiAscuqHQJ
1kyUQ2kQ7SQocOtQnd8x0xxHnO5JPrNZyxuMiFTrmVAPu859vD4Tzm/grVV9HRC6oTFpvCtcVjzZ
Lf9nLTIy6onxwuwagD/xp6/qxwCo+aPsfSotr2Qk8DyA/b6zjLxXz0jqxAGLUqpmS8YWCu/ElkM8
OLW3x78wnxxz5J3InfnGtOI3bIGUJh0AHLVJFZNvgisGG8DREo76Di57DseMAJhNvHHMdnL1Ocx8
PIwPIpeoZJvewi3B+J9cZdxu9TmDexAkParjF5DglB6nXKTd/DimblMpXxFCMPL0V6kuAvquGtc0
dZzBzLe9Khc94F+CiJqzjGSXAapo06YCf+b81DtzHDXJ2lqspdlLuUJROIvc43YZB6UAx+1iTmM1
9oAoGU4+LrgJkNqejPc7gZlzJjCKWHmrIgwDkukQKYU2cSzDR0gOvWJ5W+7uoW7fTCG6PSPKCnIe
LKtUnd4XQXQkFp3Ool3uLhX0yQ3/Cnq9qUfOmXKi4VJiXVdSdYVc6Y8pbcJgCESv0xwhSNYVS6c4
6MRVtJrcz01iIbvLunQzkMFubrAQawVkopxlXT/+Hwd5PawMM7UnaFzLs8a5DaSzSSQPn/DQ7Jho
WQ/C9mN9xPT+lyI3pmTC8SrMY3pSOSP+7Z6ITCcm97J3+XBX/zer7Rv7sfYhb+nx03eKpM3m0Ndw
kEjUP+ZUZyOD6L4QrvDbY5goQIgBq51L4sXJLJNxvCvUMvqooK527lpKY0lLevnaHeSqQzknvbrm
6iPagcYPjz/CyIC4Jb1AKDe01W9Q165ulhrwo5GOkPBgGdQIvSIjjulbgVKm0VHGt/49N8EBGD7E
zUxPrXK5Dz9yG1nJg9NXWmFmPytvTKSlgG8Jo/wnNnL33v2wJ5DPaCQwEojxGPCrmyhzJ0xS4Wj+
jDQQgUFv/bJAakIUMckW8NoCUI/8hAV8G03121VAPFUqimBguc4d8RnKCbNyzlL919qfHh8cTpoh
R+powaFwKvglSC5WyY64mtPs5syPJQprq2jQkR6NKd76xxDEKRI+igYFsJa0fCm0EliHRDkLjjm/
YpUdE2gAG+F2NyBW2xg3P0Xww8H4dE7k/eo0lG7/vNAAdqcDNhEdrahIEzvQdBV/Uk5qpyOHfzJl
kXFFrygWvgHMXWG9NgG6pKiedAzVTn3lMvw8dhdbBTVsj3+GeFAofWbeQp8UYItuSgfi1wopPqq6
8BeDk21zzfwGb84emHWVYzptRiO7EEbI3rIsq6YN8Bd5UXWJiCrmMmm/P+4P07F3WzkttpmsEs4H
mlEb9ZJ9HlDDZijx8Rxw3hXzhremqFHnqTDlq78ytrqMeTEp3sFQA/WXAzSsGDXH0balnVrX83+n
hELK4JyJd6JenMgZIdrkhDn1/IWw7eFwIHScwPJ31bE6d+5ibnb9vVq++1E+w5S1oJwdR4O5pxK9
MrII5AsiDM1kdedcbYD1NLmpyLQRZH8P/QsmBuSozZD/n9N7tMWq3dahj3Tig+YTV7Oq5LShOQOG
vh609xvgZ7o79muMjkbMCSOqp4CGlIkABLoSLe4UbBuMDLyuSupF/Bs92t339JbjVlZoxEtzwbAl
eQCGgszNCudeqZeJk1CH8rcAGz5Q694CzduubogwB8wn3Z9SmRZb/M7wTTghVl06i+wWLoOn5tIV
DxkxKJfdBe/MI5MOV+IQxcwUbNhIQuB9+lWr/Wa0MdKlk2jNzJ9HR717LpZ5B7aIHMT0YJ16t6KX
T89h6t81pFaa4697URbrwyiYLD9diwOYXuYcrcFq2bTQPb9GHfiTSTqoWTDp/2C7VFHJ6bIA3cDF
93YrrdMyOHdBbGR6pVOOJJo2g2iEgcHwlHYGN3QBY/Mr1cGLxtD2j/68ijToF80RV8FOrkdo3fR1
Db66F1vmyEb7Q7lN+3xX5FmKdaJG1srMQddzOy8mCojL0rYyhZ77KKh+R9viVBPzWZ9PK8TRTYSn
JXhrxGBAIXmMYeyPephjiqf73HaIMeRQqDx1HcV53BkqaIOSlDJirHGoR9DHFIBLtPrJQxgZCEi4
O7pDj/Unf3/F5cHiaEmK71WPX5gvRaUrmNDpjcTxnv4DiNzfxetTTnQ8Jxue5XK8d6wXsLh0Q803
kiQx2LYtEFp8ZuIHZtEH95lvjrNNPcIHxX46Kzm/SJJGwAF5NWtFfqxow74h13E5mMJU+iBzsRw+
mdvT5wNMYvHDJ2zGgQWz3V98Y08ko3Y+Q4jTU5WRiD7GP08jEPAvZvMWw6v32iMSo1pTB/2Na+MJ
3wvo4DxumBiIFeeETLueDraOx9UXEuJvDlT9C4iVn2I3GGgBb8z88T8TjzsiTMsp9Z1QbwnridMK
YLkOEI9p8jvT7WZIUcWUfe/uK0/Wtfi9CFKgrqrd646PbwN7pmgplVFjhQSLoy+cEFIJPl2eC6gU
w3kGqcwMaWjocFECBwOSySygWiTrAZ2SgVTgl5w1o4JYdlBMSAJayQqjxAeQuodgnqmrm4kOgFzn
MZSxGMI9ilFt+P6eC+T28TOi913KWZjEjCpP6SROWJjLFlA0r2rXKOwOc4+xylTXjidxIgC+yS/o
1MFT/QPx7DtcwEjtVOUbYyhvK0lmCluV/8TvVe6lm5OCYgj9c7DPBLRrhekvZ/KlUaCWTyAG1UyN
7ei8hnZIxkffTAOXfdXAPyhnE6tc7VoX3QfG+8XAVSV/HifRH0HKSGib0p/mlx9gjp5f36kbVEG8
vuSXHKcMwQJ+CQFo1FQZs/OnU7dowWd2omRncHYfFXZcVdA9DrJJ+xOLXlaJ0ukYSWepUUv1lg3v
4U6Xg30InSusGVcSvAJLsaUulybh3vGys7YIqYu7SpTYDOlt8juqIbmGiwDthuwWUh8uTPN5dgf4
PFgo5ENrD7YJr8rTbiAwIfs+9ET8pVPShxSqdBS5FAids3RqxM8YODMyUt2b6tu8NpBnQgM6Ee1f
E4wT/9tLAy6JpmkK54pvQ//aFv5wzjrOrfZ6+iYo7pCyi8XMtfMrsIZSC5vcqQubvCTgTyTDDvaa
OnwVwX8yzzmJO9Udt1/wYwOdmEvsRY3WbnshBk+Yfo5uoETLmLNj5G1/qYKrd2xGcW2Rl8KKeLb7
yRp2wZEFpIutzK+NGNDejZWTXoWBvmEUE6JxQf/k6cwt68wFBs0ylC28bAMtELDUIt4E8XqLOt6Y
eF2UJC/Jsq2x4fwi56/RoZAaeLI78WbmqNkJuVD0O6lB69nuiqu/iBoq/PoETahcywKnO2yT6kdA
p5J3ebo3QxZv14X4NwkgBrtL64TZTOS1R1cD/Q9fqOt3WmCa61BNu+ZEannDPBvFIVTo48AXOD33
a8ldUkRcuoHWJ5H7EOGtAY/Nd6iozdPy2yme7Tmx08gdof+x//CVTPx0AcxJOdYmw/jSl0SCf013
Oz3E38noP21LKxVxoJXOhI1J5qH4AbP8LqC83PAGFbDEwKXKQmiliMUeuQTBztghnwz1p4NotDQX
bYqRboI+48qQ+tqIsMBCmLEWd8dmedGbKWt+pFRTMOsU9DzjaxpIAUWVdfpV1+krFZDK4pfEtzH7
LQO7muggGKyCIPUHLeInUIHTBjuwyoC8lW+3sd/VjcINUP5s3GfC6ZY2tRwWlL6N9uTZbpvlxsU0
38qGJ22fL/jdvX1Y7SF76zlU/PjJqetDwMvP57Jhth9TvM+rFLh0E0jxqyBr2TlW2EWkdEi4746k
pzL9Jl5GqL9fvdN4yiLuCNvhZHRqiPLx5VYyAqHbzsb5K3UFoidbLBf2x5QgZGgq33CmKlxuejaQ
QGpxOtdtJrDmkdqdbeBZoCfifjEtjs81PKQnNThf0UjLuthyFPKH5wmXpFu708/RB3YGBY59h+IE
a7xQ2cPxpfzyrcnVMbBRnacpBHQiMocquSy8DiNy6XjwcRj9zxTeqzjka819xFAjz4CJ1ssNxILN
VOyWAdAcg6W6AA31UF+5G2+VcM5fxkUQOERBF6eTTIzHNXVRRYQJ7iUDCWVauOCpy47FffORsfec
rC/1TAjzE+fGp6ADkJZ+o8C9oVi35IxLCuzEHb6iZMWLAx4+vNUnZwf7CoUSboSsB6WdK7romq77
nRlO/nfBlmrWMoCKfFzWctX4e8FAv0afWTT1+564S1EAWTAqliiS8mY/ZpSiHye9kBx/77fckw2y
8wFNrPcS+eMyhLcAAHL5O95ZViHmwqqZHAh/I6kzkxJtg+DAYL0MPuB9QRfHziHDeFXpry84GUfA
fc/6VdSphUimCfyzOuqb6TbqNT/eV/Bum66pJMDhqFg8Zy6qqjtwErlgO2/2c4DQcq+X7E3YrT4Z
cz6tVSt2sZ4unqZEXxuI0iyDZMZTBmBHq1Vn9q9MVDuyJ7aIyxjMN8NOhzi5Yaw0W7BN8gF0f1ld
L6zLcQP825PQaxmqzr2qd8bVDBkG1VSyIqxirKgulpVThPdKsgcapQcLpYwdAQ7OBw3hy95k9iv4
X2Eh61iOX3z40951Hp69oFQyK7Yak3JgfR6B38G5TNv501IJ6m0yRQkzxzueXhPEu2y2QHrvjxrh
R8KgPszPtFW6sZnP+V6HL/Iwzs2yjTo1ov+wTaqUiP1QB01zbDYj/GpuFcaaIP+fnYkinI4BC9gZ
oGJEZ+tt8rddyQ34vRh+s8Z4hVnFQUUA3PUJmF53YhX3noPqkx5ZfL0wMlAotjAdGgyf86KtJvcD
lAoiQFVQfRIN9O+qXnEFB1FnC9bEwlsvbNZ2FmiRq5y9xmYNIdWmmGMBo3jZ1P7FLmaf164ZSt8L
96yR5HGPYD4i+ut6RsKUqCEiQduJtuRqmRvw90+J+wY7pFXgyUMLq7y0LOOBcYg2j3uOj0jkZw9B
UhNMbfO0X6i4yNNRlGtatU5/hjgUWbG2Y+KCzQmoi7XmSWgSmQHQtV5VxbO94fsavZvVWisp7dGc
kZZWMW+rKatWE5Yo2kkXnky5/lZyss+QlzhcqHGUx1vwB2JE6rJndaiKCfQMrtm9pnsSsr95hYgY
jA0m9mGjmpiUrDlXPhNUAs6RTOVqP5wZTHpBpSiIiPmCB2N0Zx60qjn4l1fOC586M43QkgPlARln
qFAcLCqdbga3GELONhcNXw1VAQmtqTsIFhqhCKaKvHuWplfGEVGHZAmZlYI7UMS9Ig+r0oia/WIZ
2ywxaRGidDewRU7XvdbAchvrv8cj8pZgzjGJ4o3tNZUxlSmVTkoRDhA0pISC6gGEBB3nHMdaJSu5
Jo+BOe+3OT6L+5Gbh/G+62olXiseO56NOIXnCrGlXMRLg2c4DT/1cQPXg1gHh0e9eRAEWG+HIraI
4cPUKZDG0gxc3yyNOmTS4B+r3+4zObyb0/QF6ArA1sLzipHJVZmVrcX1UoR1lo4w6sZB/cGBUoII
d/FiYTMyh45VcS7Xb4wsHewAM0I9tYYyT7Ruu7Sjn3mdiZ5iLTEFm0H4Ak2JEVvUGUqv9UFQd7Oe
6ocjfDJKjbtGiWkJyc31raCpJM1opJhibrL6GvW4pmhGk73UJde8SBdk7ftoBL0Bc/D2GNp1VBUy
1kK2o7Brb3Qzehi1971CdIPnl/1pHI4FujxqVQatfBQ+m8s+qgodyt0eciBuTPAO6WigYHivvr6D
ck36WwncSqOhcjjXKTj0hKkI8p5jCInK2WQdMjANs1x2Dt/JOwlYHUANhyllWdzJIJYn6L9uBawT
mdftejHBNhgdZHV8K5CMmVUcvU08FDGdqUzDJt71J5ekAAIfIUCTMZEAE4xZuv8KRxzyhJFcdGQB
F+lnXkXEQXJfwvyVM/1uWhCjmzbigdCFW/Ut6o+KEEhT3hgAjoiPrCIU5cNahrfl49ijY0hSJN4g
hUxHSjAqDcYqwFGo93apXCrx3uZ1rR2qsUHYzqxnmvcmXd7OYzmJO66Ls2FiXm/ywjQ8h0dL3yU3
13fM4JziyUJPo5BCnzIoY+gfUaAdm/aKdc/E9Sp4raasgG9fJjbVBcmadkOBPl+1HHwsMOnHrGPk
Fa4XRXuOeIWpM7SrbEbudEvhk9k9AMLw2QDSg9GHg1pdMDX2ShFpqRARWt4hb7tMT3xVpE6YSet8
cl/Vlo7hQ5E5DlVuEAWzziDI6W/PWTu/HyENzABQSDrF25keqdyK3Y6IkTlF2pj2DIwcZcEslMea
UKwOSAJkQz+p6DnzePrzxZTOnjWdDOF0GvjP4o/9MojwVsWMCTFY40plFrQiTA9eaPoaSHf7AJ7z
tnOZ+zq9aocdYGCpIinxaiG2iLEpV+64fQ5kqtsZqkw17ArCF1b34v7yApG2OnsrGb/+eNiIAyvO
GIlAGwPTvsZwoJjew49jNG4bD+vS3pKgH+0pg6FvcL1Ns3LnUtXCaLXXZ5sOVO31M6LNH57NXS4V
zSzJBxFEAuvmncuXThZcTgsKcg20XmxSHs8DaEiMSw1sfq4DTAZLV3f5A5LOszfWGIFXM4fWQvm+
/qi7+rFRIyoAQCPrTJyW2QZZS7MwoaY03cV2Vd1GaDy/Stkg64swk41298bxfOGOh9UxK7+rWDbA
+cfKTpyaW518B6jDkVSs9iNpn1g5BS6GvCFud50InhIHlrqLYf3W2PY/P26WsUmQsbEs6UhJNOIU
XjqotV6f8FpCwDe0y3FJlKQ17UJPPsX2mxTnCooEJRf2QeZwEp73ZOpqvopWg1WmgSSQKs8BJS/y
ebx+/Ll2BnMcifYZoEhtzaMVUifY3ZCZp3FlrC1L9pwyR3Umquj5VuwWYI+6TMlh7Y6HoQe7hVvl
6AP1MKUY/7/SGQSBSWEHPKOFAkcmFrNt8zNPAIYP1y//7tluIa/1pa//jYTNIcuwbAIrQl90149B
r99DWZ2ATBm2PnsFM9maEnQtG2PPvXVno4InN/OJx9El4bUTZs+q9USODkvzORfqg/fZbxTqPUWq
ymV5PVGz31u9F7oIHHmyKaHRvTF/j+2IjpJ1PAeNfHfDvHbjWyjTPbHMyJm6XmJrt/h6DQrpurLf
SJ1Xm2zzMN5M7S2skpUITLBdZ2a8zlVuHi/haWFYWuQii5sE3k5dWV47+RYQEqXXcn9GgIOU4e5U
5xjZchYfiVTnB9Cjp7m3RAeYV05ckUYzR2R/aZVvBU9T5nwMaGYacaBwSVpZG9xWS7ZIh8Q0rhqO
gLIw0MvDprUMzOPaLavJwzFXRPu9GhmDZKRcLLjqh5fGtBZOUDa3kNUNo6gaZZ0Ent3WpbL1SAnc
/MZcbKykvIQfQHssKvCb3vcpgUFVvTVCRvMP8MP1Lcvu8f/oMVRRzh1hhptFvdociGdIEONMrWtY
tm/QLTbRX+qhRj3YKVok9BsDUjpWdWJkLCxoOqHjVpMLmzTe2kbXM+VPafeibNOoGLQIbLY1LLOl
IkyxOShkcK+nJEqUnRVTCTSMDxR2bxkQiZ09XH9JFVUTqU/wtieEgtB3awj10bvyQmhkmN79XME4
qnVDrGZdN9i5sgOBvJqNdBcF50+pfP5xT92rsPM0nqis6b/y2nln5I/u484rNhI4+kIW9tjCVus2
uDeUFA9vvMHRaIVwwSPFjxo188Thy+Eb58A16oOvI2/FdlqwCRDOis/OhFRz7FOBM4GQHP7uVfVQ
esYJtrXNInoyF5hduGRHf3nS/4FmGmrhB1h79nKQE0amcuTJN0h95WKy5gog2ajHPAqIdrkJfk0I
vzm2jWMhV2X4DNSXeBupMvkIXELDxkO1MOI4tu/cUxT/joT788h5Yq18/+4fDME7/jXRNCG2WFzD
RCLucyRNb0VaRpHefH2yxH5OpobFvRWt4oAkAqjXSy8EHks4sMWSzEfKvKyans/R2C8q6DI4IyFm
t7uzxb2u8geICWHl8m00AKCz3sjpWcAbqXt/i/K5paYMuXkzwyZFzoanBdzMc00j3qYwUf5vTsTc
KYTzBoba/HjjvOXHuZj+YE/tvoKdOdyK9wpcRPy+3CouLr8wX/1CL/5RpEdUpI++Far/+mOD/Nw+
Z6KlwhdRwDxIfFL3LK7q2T90jyUhqRa5rJdCKg36Ze96rnfuzWE9rqWXs4YK11NMnefYxx7io+7W
dikT5e6ZlgmOoVb4s1QrQFFm8jjCm8/rpR7pEwwrc91wl36vOdLO8nkhMb+TFz/GkTSTWv5aXqvU
a0sqVuO+/XGySQAD8hqM2Xjfr9AK0skY2IST96tuA72iS4CpBsXwyHMBv3KXHhQaIdpcPrTDKUH4
D/q0PsLvDiidKpDf2dUi+rWUq/PbLr1FV9mRG7KIn1tfDMz5QKeOUwuciCz5svFBfZNZUGEuKEIz
KUiZKDvxpnPksSm8KsKivtc813NI44EumZ9plr72B/fE64KV4l88EvO0RdHC9w02I7xjrXUO9n83
wURL4MTmGf6K586AXNbvrenvQPUIpekjXsfN/57ej2RpoI+AHi65qShCAx+Z923V1P7xPoMNnktJ
2zIYZIbRkk60/bq25AAQouwZixf1q8nQ9CkLzRugzQyyIWYunee0HUgxTeylczVtp9MagayjnqqC
eHCklRX21sJp9YFJv2ukhxg9txVFOhQCvc/x6RGisshy0fadukmiCP/1G5Yhp52CtVxp2QRm3pKj
cfaNy8m/zyasj/DwGL/Gs+doVVGIC1YFC0tioj+GTmGFZK0CA3wM9D4Ff8FUXGfCdFNzpe9i6Qlk
N8SCWtXqUyNr+5iWWKRzlokdLK7ogZ8D+St579VUfCpSNMCR/6xhy8NlUTRF28j62CcNv++35AzT
+BJAJ+xdo+iZ39wYpUQYv4vfcKARQHjdDeMJF7sVEezcyUyirSI7Qc1qrIHhNZsScglpnGmNvEXh
BVmFdAFkeaivuQXLp1We2EZExtlsBTIACA+1i8/sn0zxDw2K8TjopBoEwUkhadh5q0tSzVyN4ebA
NafEY9zX8+Tb5s0urfeA3gJnUEkCBqDukdJ7V1vTkygjpY3YDNTnRhnZp4Gg7LRwPlHsMC6VqGpO
MR/iUaaPrdshcgvothflpHiPOJ83Cy3T74B30RGTSjHR4uQfEoxxCjoKBgWOKuQ7TqHRo02bPtOf
9OubIbQj9587NPKeP9aDP1uT+gRBkYczwRUzjr2p3NesduanzyGIuvkZUryuyCWPDuvfUMjGry4G
44zgldzV4gTuEaiR3yRIKxVbMxj5sifQdMFhhJRQdypzuqPHCs1bEj8wxcCWxVtMboPEd92AEbdf
t9v1QdJhkxYDARKTTcriBerZ4A8SWklaGNvOcu+fCdI5QWpM2/Mhy3mIxC4kdsY66r8LCPMe0IpI
oiLtTn//3dhIUhlRjo3BecaSXV9KfL37MH0z1z/FTk8Emka7O/3Irr0wmBTX6tkODau1kX8itjAn
5mTfddhkd8e0Ney8O836Pz+Ghplhw8J8aQkTnpzbrtLSsmKHsMGxycmBT3pw/uUKUsISIdgQkLBc
a18VH4oAz52z2aEFz8yo7VXQWEzKwc3YGlTeIJN8Mur4iVe2tSY5NIMpIQ80gdsab2679w3fgN69
CLXhB60wKpWJaywv2pyrBcjr422Sjbx6jOHWb86Lpxr8I3evrfNEzBvbN/nD0kbb1q2SxDjT3Q3l
aUetW4+VBy1CAN9QtR1sMJxIsPZ02FTGKW/hIyl123YCiY2JQkVaJr1pEPm/u2fKPW5m57tEnm+k
aBjU7KeHNIEo1BbedsqhaPgSl53Do27/CVsZmrGqKL51gMLW/BbUEXEL5knEKPeKP6pq7sL5bpT+
U4pr/MZ1WaX3d4j+PKgUarOjvrCJ1lEzVOsWuZa2HCZHub2zH6wfoi4+YLMHzz0NXQDY3HGt1cBh
QspgLOYJQkrJ9RE1ctrvYk0scAvICJmAwrDfw6mBppzu0CuGCCR7w4r49q5Haf1CsH0B+Vie4itv
quxPqCyHC7+tuteUU88PM4JpvdCH3OtJEYWDt/R3QwotacsbJHQ30lrlIBbN/SZ3wBhoSGh4DUyR
osvIkIAKRH3ItV+Br6qayYIQQr9PjHNVZB9tf3+9dhbLMHSyVFApyZj1/Do1S+cmZHF8ohp0iNgG
gbO6aEyHV/cvgRBYTXky5blLgwzcNChe4P+W5AjkT7RcCneme7gFiwxLWeclyYMppQasDZKI5Ddn
pF+Qs9Y8Uu9lqYtJdmh1l/A/bkeqI1BXV5V904LWRXIX0LeepmqkNIIL9Xov5xItVl2HtQTgbFdS
LY8Q+8UvQ97Pi0D+bk/E5w1X5WG7gFXK4LQMIhsqSTyUoTYvJjfGY5ejpg0yxR8cnpcRKNdbvaQE
ONSBjPnyFaC+TqECN8yH/6mbx27byjcsFmqU0/jjrwrn1AStW9AQ6iQwgtBAGWbH5NQwxQM7oGEV
KUTA1fMZxcy0FTUPFRiuwsuoK1ut5j5n8RuY/VfCFrlpk2aAzymgheroICvrhRCmJrPgMURRs6ag
LhI04HpEwUJS45tVNrMnsr2KmxrpMqUG+joFMhlm9l24s4M5m2ocp4qgnPxhsD6yZ3PC4Os844Ga
TF+Ig0ScfH00KqXk4CoGawzzOIkOPHCCpAooGL8GTo8z/+Qlln/SNLkjDdvIjtX5E9z2wdYQnrpe
X5Y723eqw5DP4WV6fX5JeuYuhI9im7S2SkQdlulDPE2tO1u+F09ELtcsy5v5Joy9K8UQZnQ+gT0L
6QxDNXMKfO9A96pLwiJTe1KIaxpQ+T2DKKQP4+leu5/Bi3Ef0eeGmXxDNziWVMja/GYW8CSWSAtP
qRJOeLa3Qlj2KZYd5vbdNHEoZ2fYnN7fyommR/4j8bHHnUd4g3Dq0nnXv4AhZYa686898bajlCcb
KN1yHSog7FEe6rEAFkZUgOywZkM0weKRojkSZOuceIRADbSEphbpWFFdEGQItikaNHc9OvYWc/Ih
e8jY5qd1j0eRKqqIXTAFCXnkVN15NNgwv/BeHhhD8pFK62ACsShYwRHJJS5Rtm1XO3M7Yt7gmtIt
wXJIqmkr3GMZJzIp7ve8ymZZcLcw8Giv8MC68rHcWYLD6RvbBUWPUSxyG9pcswuComHaQ2xBiu3F
2C+S55SKcVJW+Qx+Z+AlsSru8KtQEA+b/VdtTdDR9H273EbKjsUU0V/jaWRq3KLLFU900u7RE9fC
i2ZWfKDjm/jWCeKjpLw3dfyQMUfvifmGHZQJnA9Wy0nX2Yzerx2Jffn7cf2YS4bodjIpWlknh48X
6a5RZ+t4xXvCkO7Mv4Xc/JFtB7wQLL+MDQy/Z3kk6TxVP3lE+eHGK6Y9/o2xIYHS2U8j1myf6bri
HqxK1vqeIfIEIJ6LunOn6N+PHRrClMM0QpB6zktomaU5dz/5sD+cQe8AXCksv2xbtHxU3y9jV7Wc
kAqv/dEGALI4shqh/Zl4YRu+RkDW/LvLQXOMGJR8GZDbbAlHgLImRMHgxg4JR/abv5+h+5SRKwKv
Jzb1syxJjEY9jkjnvIWQPe8ETcGwxYeibie1ufcY/AzdJtveEajGraxGV5M6lReSS9rxwpGBJbEn
cSVyLuvFTyAEuHym6DbNthjWc4XDQi//7H/e6KrjPqcFZ3cZEbQwCfIKAajwKz01/VFTcZNCMDLD
WTq0l69ktpT96OD8OPljI8t5EZSJUfX0fvsx9W/3WPvxESlRBT6xTvRQ6eSCk+zWZdbort4yOSHe
yvZWnhw5E6Svgq67AYM03DFjZxNJl7j1oess4jUHu8tx64xBzNZSoKjguUi3toANU3sLNGh2x3Kw
WZqH2Ufz/6yOzTwWnf7U1tYVbwcQWglGnGaaqeQvK6h7/Gl8u/UOlsvz3Y0azUNVVzUQsO1pDNBR
zg1NsTUnqi7ODijDjUOr9UfAQy/3Fw3EFd5UouBavSXcJYnpH1CkQg0n8pVFoMges1mocEuPHCcs
YIXx9p1i9j/Q24wQqzGI5CRi38C9eaOCIYhzc2XCOsPunAjiWtCsVshkDTYSfRWPqPak/Su9UNcn
7QXiIcttgyKJi/Dax9H0Jv506sfPp5D6n0i8LiQ3XZv2/nq6K/TgQ1Z7xZO8fHkAQPoGakOPc8V2
zVg5iFPJNCT/R5pt15JfEeWJtHQa1I1u1Szp2qTWIgCR+sQ9orqTTjSmOD/2BioCYSK6m0I5dd3S
clWaL5CN4DwPeJp2kHR8x6/oE4ofkgm9TrEBECxYG5RPE2K13NQJfsFa3ACWW8kEdeZuo2FU7u98
Avao88fRNeSnoXvUOnb7rSHeMjaxDnDdDtNyAPyJqDsOYjbfEvnWgZFxUb2VendNhnr8wmlenRb8
dcsZUMrheyqjPIdabYT1Vj2Ok/a28ZQx2Z6x/5Q5ta4+tZmTWdbedlyWBC1qRk7ZmhbovMqDA67d
mkw9P3b5+Egmg97e49vec+8Aa46hzAlwtgkm6GIBvx9YXxD2tDK9NmNNcpG1V4q7vlfTktCpHm7e
UFWUZuFhWXKGnuDVWi3/+Qy4k7mdAXDufI4BqdDNDWIT9ZDOW4V0CyK+3v5vgiSlnzX+LdbS+0iW
mHGmBuH7fFUY9k48RhyCotnHsBu3SULygpkFHfyCat1XNIPge9iiw5lv/PQ2NJu20Ttn/1e0eE/2
8DKf+OZB/FV+IhmZRS3e3wJ+2lGhllwOgTdI+8K6JEBDdUFYMoCJZP+gpxef48zfEHVBPpIq5g0Q
4uw1DxTOlUpw3XVZN49XP6iR1ZP1dYjHi5pPxpixuzlvnH+csHVnsfoQCWhUV183tTffJehlqdEX
n+EdytYyivwFCy1mhNZssCnCPXuq4LEbAyR1BsQzLruLqF6m2BOo1v83t9YtRfNw9DujdE02dOoK
TObDO2ZSLs83ly4yB+LRMGqv4bA6726RHrQflcchUaApYeJNaPx/imcvOOO2GJGuXP4vL6CDZlZi
XnImmNQxEHrwfi8AtjUcRrUCrlxvfx7zV22kuzFinSHt+IJGAOjkoSHMtmJsOuHR1CyOxkRsMY2z
WhTbiot9Cm0h7pXKxRTkCkAZHVfp81WVPl351UP2vzEOcYXdSftrIY7yHMJDeW4s6aaPXeAWtROk
zbBH6wbJ7XRbNO7iRrCvuj46ozXSanh1doP+41yMM6YiTMANK7B2YNchRC/v+UOlO57jMU8umqlw
JyikKGD0icJs7GhplyFpnHuZb0ZIahU9Gp4R1YmqT98EjzopL9r48LveBrEn2m0iBhAnP2zk64Wh
GN6Gg3289NKT/02F3ajmPbkh7Q/LUzhGLb0I9Y1qMZi9Ux+bStEqWpjFDDjtwxVDQpfOlgFXVk36
YZ0TbCuscwmn1F6YOZlnsqeLkW1vgSuihymgSRiUxpcpOopmknfKIH7Q6Cy+psRBQyfb1tv8IZ5a
qoO1jyBJvu4U0QNyvqCEjmAb92OKIEshpgFfgmIVYtc0sS85XsG7sgO/VxODQ/TSY4qXqdPZlWlC
+aZQX3xaV34imXrO4bPx29OU9hArf7fky0vkx+f9wcBOcjI0rB28unfip2CfQOpNmeoHqQ0+M/ME
Hr9U4X7ixVPjNLQqEPLwuhPg+sJpAJgkoXopLa624OlDx/H4wHH4Ga9Z99RYZdS+eerEwwwjL4l2
6gLwlwWsIeTLO4WRQ41sR5W3mcVJS+YRes+/G1GJyqhmrNfPg9qL3YTsI8uXWa2UXE9s4Yu/XiSr
k5N7KeFaSCgeynOxWLGQjnpGyFZRZHV0mEKslIlUdIbYfRkw/DFrqMvLSadvuWNblDfSWcO4Fsko
n5Xuv5/nvqib06BMX1jpUdqRSyYbUr0aqvTw1liNoJe1RvZz1xS6E8ZjGSIxVM1K5f3+dQErjzHl
rewopTyAHoMPwzseOi2xI//tfLEJBb56Kk2Bhvdf9j7UucRNcEgwSyXi0VgIMlQYgH6foBRIZNdz
8WzGKkWuv/fZin3OjCMJUMDBlb4P9adaRupp0qWbwkqVOZZDfPydDcSoiNnz37V4JB8mxFldT505
eSbBkV1str0HZxwybg2aOzR7zYXqb8W8WPGKDJ39yNta/w4tORzOiJZGzot2hRHHssJZt4S/XgR7
/Q5ZSyuhJ2xuIo6YMkdU3yHevZGhw7EgML7sbHZK4rs7AGtIGFa6Z4MIHa34Zw+ETt7HDP6Gqdq6
2fbunnRlN4QYTKiXuBC9ala1LLecIf8J7fwxwlFsksYtZ42pVR3kC+ji7jZy9M3/m2DpxvwErQzU
zmHc1nl3pz49jEiGLv4bjdXeb42iihq8KNQGYyHEQK8V3id7IyLgkDVSPKYqkJ5EWMnIo0g3PaaX
J4fydLQbicrkKxCP+U1UUQctpvG53EpdEHdidVKKLLCl5FZszGKqFw9wat1HoWzLteqd7pZqjrQ/
OWr/Jw8fxenCljZ/7OZHi//DspK8qsi0Y+F5Kg7i3IQZnkXfqyCZ2JTsilftqLIVoz4C/FoLMQih
q/Ry3VJermPF+Dq1GghEbufh3OtKXwR/y0Ys/zLPCHsG1R7L0VtY18Ik2SBVyj3oWDCSuu2EnZEl
nVDj7tSF7aiuZ8Ys6lYVavx9fhOS0E5YAVCH3Hih6/qOprDFZwnkwA764QJconGnFzplUuzhJRoY
2ZPbt5YnIV17g6G69Ly6BwFKa0ZBlGA21p33TTJJpXLBohu+vDi6uWz8IylzoBGwGtariag0eKPv
1lZAzh36U+mlhc8beRjlpaNeTk+ujoloqtXg6gDW0TOfLyb2tqPqc7PW8eFREmVT2hL6DTymI+N2
tu5yij+tHBVtkUAes0NK9+vHODuj8Q2/nOZl9MZpJyZSFzTzmGHjNB7j3LnHw7p+OJ5/IyeVgxTK
rM6XKeiWXSoy8snlk2UwDHysoS3Z9rM1TM1hCqzmqjtpDNstSjI6pyHqRnngccVwVFJPtEiK/GGR
JSaLzCxygmjEqiNppiOnjQaJxyjM+tXdggHrAolYHkapifzaCPpesM/ltu1O6LkO2v/BHfhiQQqY
rz7yFpsow9lei6E4+b02Iv8qeqA+gknc6TlH49zR+1h747OXD3Z3lW1vUmbujKcIsD4reB/dkYxp
eRkhx879rIQkp8CJ8OFLGHKjVgCrslrphDf3RlqDNjdSgpAp30NNFhZVDQjNoIF+Lq/wh09xkVuX
kEF5VRUjxfz48agBt0PPb6zlqLXx7KuGLXpeefX7Mozljf2iFtks8KuYgtKsyDkAuyNEsFUudksP
z3tVzpXe+zPFjO78h1w02nuBL4Rg/7CPjOX4T1EtGGR8M7H9aVjDK72PLccpX6RCla8cgo7aDXNJ
6mjG8iixffBblJjAcSfmGNKWnC9KkUeoNTVe72/Wm/Vd00W8IK78DFBk3/Efo87P7aOIiPZutO/3
J2HCRVFpYi6QQ11fOwQBPdpO9vJoPjmv0ArJF84reCvlFVJXoS3uIslc0Xy8/JcMGpI63mS9Ns71
+pkbyP8drGqzzpN4CEqxHvM/wGbYLDzwWtaBTi0saNiFBGcOJUnp1T483zTsa89VwHpj9UjrzJqi
YzpgNrah8pu4Ih74K8xNtySOxFJfU6CsPUFsK6cq5kTwVQLSfZUSM5lYZTAe9bHGiiZTK2WFmIHe
xayQgjqOvY+Zd6YmOz65Sji+rOMyaN0uY11nWaQe9vYDCj06hTivZYvyb/WesxO6uvxk596hfMNt
wqjfkM0e9NTmZq1fU9DMNVa+V3jY2HK6IBp5CVusJOOVuQZqMM8VakmPdg8LmqHS/sA3WHH04m9/
oBMbe2xGS8tL4IFK1wpFlcqmCnW3Gi7novToUrrpxDEcQk1UBaur0FuMBTiqYKvfSn8Ecyh8fOJd
SMX1y6uJJ3XugK3dlLjkXrZaXBmNq3/8vlsO1K5Dwtvy80GZQO5c99vxDQc7aqEoRjTlZr4Z0f6C
Zjbbf/PnwEioCDPPY8q52nqdXg4JPz9/ZT/DTL491e7PIMmzKqcJOILfYIIg1k9cN4ycu54rZHyV
AkTS35PJHclicyRUy1cAUk2bLI/1kX7vpapZBjQPTlUZn/1kjKpMVovJYd0b6XU6C3nGalrJ3UF2
BSsuAFT7AYszuVO8xyJL2ZUNe3DhGYUPuuY1NuXwbmHp4UjTs+nZzu0ava3RmeeBOarqFhmeggG5
3NJsqVV1X2+6KxpLjC9cRBt9Ig7UbQHwkPx/az70pOD12yw48g2h3URtf+MWmx31MPp46opzNQ6O
nnqPVxgufT3YRYdTrD1stCrwXyiA4jb60Y9gUtFn5GwY840UCc/cChmVdn80+dJsp7MbHuGUfjzx
XEtE99R9+mePLJhLrcI4eaxDDbulzVRnL3HKJWCMTSZ+lFFXslopEhLe117kHjvDfJ0XWGrgC7tL
m/3MGrrY8S5iY0JMmxJodpbAZvR4QE4ns0L3X+xpdfEsdwRmTa06D475rJqOZU7u++Y48ed9mp1W
dpixOP5mFK6tD/u6IhdIYHhUdh68K/wUmo+yPcyL+0GpanP54r8FIWnan14f2ampOUyCZSnGW841
Njmu/rDeWdLsT0xR2X5IO3YZNk567592oQyeYrmcNjEGBagToQ4OLvmm13KM6bSrrFfHv928DmTj
ygjeIgwkqsIxWEu4FELTayL5glRG0TVqauXHsWwltYCwUSOkp9+YxnuhzkbHp7vaG1v//O0ZWxaw
AGZtx/IwUPGVWa1SrsGvBybeZ6xfDgW/qFGl3zfwTyWkZYc0PFZRDKXj08foxdfzX5L8vHwpkSNN
YCGF2PLDKArA1eyhPnGj5ZucDTfORcDHIdYC6osnWl4WRCkwzTCortZkqWqBCoXzvjRBk5s0zcNq
65Pio+Q6TdzcmiCvk8mbv4k3he5iDjkKkvHMjy8vJencV2jaSDFxc5Yxm7vv3EULLnF128/FQUqn
jrA0tykeqg0etfaRbLTq6mnR1sY3aChGEDI0zmTINwLKqk6ucy5mJA32xEa0cnwOFHjpYX/D23vw
88RA/aYOuEbzv53iQwIJdpvAMuTBG95XKfnwxUr2YLVWFH5rt2YfBYnZbCKy75+uXjP141+PMF2t
SeF6bLeMAOBzjm1XwslC6NJqNUhRMrQvxpTJhJPq7d2yoo/sENsOceIT4s1s/SOQlNr+UCTrm3Zs
67XNpwdZDLBO7ZtQWGiqwnLAYnapdey8gu1K2H7SaNLVOFyOIqe34mB2BqkjSLl2fUcOpf92nQie
JZFU5gQT/FAAGb2N0Wlc1o/NfWa64Sa5wJTLoK8vu7v2RHSbqcGwxiw1Yeuvmi5igwO9CbBVDhBO
pf738bkkraJfI+/Ux+6UhwerPynrrs+WwiGc9+1OKjE5VO4gSVlyfMmKPhh0FgIBbZ+AG6BK0bNf
3yd84J5jnTX7umBzNQ4KPn8ajgIrXR4LZxT4BTj/nH9VfvZ84hxa6pNCRHdzXmwD5LtdjQ/hcc4b
Ym3ar8L5kucy6rqmuJ44k1zqk1tFAQ1LPMcorh9EGQxWXfP8+ia62gqS9AjQ2hTE8ZNyu+HhWIKA
d4eMHJ5wq5UduSMLRH1wj2JlDCGc0Tvn/ZP+ro29ZbiqNXH2nqI3ojp2JA5tComLsBrJg8kXm7he
UZxF63PmbGXuYm1Wm+frIbza5NUUf1T64dh0E0PuG6VSOEjU9w0V21AlFlxY7StzdOtFSXKBXUin
JDnMukhQ1l4cXZYSxFysa6SeSMOUfcRR8MSX6Rmzw7KIKozpwm76CRabpTyfxujPLh8dD0K0wAHt
aAPRbfuqmAvy5WxJE/Sf5oKQgyVSx8kohb1zb1taEtqYwxtIf7sR5WIqFj8p1h22dg6o4cPuDatA
SiWJDBuJLtGZNg820OhwDFu9sNloZB45BIaJ40OEiVF3D5/lijA/XvGpnNydRtrjcqF7HhcNUDwN
LA4BbODhevmesgWi6ahrPZRE1ON2F1jtlChbQCorkXJDukqI7twL4WOygVt4aAyvudv9U8SC6lPj
HedlyZ5xZHNDUcQ6qa68JNQa19wA9vTxlZbb9PPSxhKitMVjf53FwIfGT7DCvapRswqHZuq1skzS
Wws3Nx6R2SYTWB/W/MHSkp6Lxe2ZDWQ7vifAY8SRGod0EO5ZRWFVo+z6HMA1BDA/G1RjkaEeHzyh
+c+f6+jMl6n9Lpey88zAlA4+8M1MthB7uTZFVqBOf4+1DXseDZmWfWWUH/42QM2eiD0xrSbVnZnB
bPEsDJYhi7nFeuBS+jN976FILX9iCq2aH7snQ6lkguIFPcIzZpFqcHP9A1IPjxvlS0gTcPpDRB7V
Wqrbt0gXVg9ER5qsH03szIDTIwT2u1dChA0soHL4wRmnn9y/irfMEUfGCTs97CdwAwBSh95cXaxD
lcyOsfjbb63aYZ8B0ibpxVfHfMrZBya64qUvtzIB4KH5mlZ9D/md2tZVv+M8ljxqABcvvJpAuX0U
JwR9IQO9Tev6mvRTtkA8Oy+N9Xs5zOo6W1ReVh+W1iQcbxLILBlFvXlQxN8C2kYooHHXayz9+2zv
SrLwtCWeFaMQzjpYjYsb7d1Od0CeSU3FwwYwEWICnlkQylcAL7BNrcUkSzM8gfiE8OR4jm58y8mO
3/EDM3wwFODzMNJNLyw9WRseV4QPoOjW9XnUPbI6nQlVKhbzWzdK2Yz/xEUO6BVhxMDYx05vruBV
U6NyPd0V8OtBV3BwN5ON7Q9+tcdcZeUbdnI2zdhdsjAPZKpmB3RaUlHGzyig1o2qFwVR36lxClth
wb6MxhLc3G5J0I0R+L4/aVCL/ok4rjtotiazEN9yc0yr4PAm5luwyHIl93dsdiKdYRDbgo0KU/o1
pGhTx0Ho6U093ivSdPLr7YdNtsSak+plxPX8HSC7J1FLb9KDxjjkqBPrTSY7mLvFlgoCmQkpIHMX
I0iRkopdQv/nDSnXF0GrLyOj5NpuDMbok8w8EKHv8CftL+eKMoJiLQA1Y3muwR3rBrWVQSs6lHel
Y/r7A42EChxWBd+vuqGlbqQlV1nzGE0LCNoB7crhzaxVGzK5wUHp+Aj6grMdPnCDYe+Vr2fMab01
ODRkYofjFfhVR2Qo7wyGXIyLvCKfCvPNdlIqS74xc58L2zpY4ndBsZNXT8GqEw1SpTVSIdI+Ccbc
DGmAef2yIVJ8Tvlti+xN6zmMK/guM1q0oALLvLPBkNRUNhaIhCoJJy51L6GsstVzB0Mwfv5Q+LTW
Y2OA24BJzrTxc8GQ7b4NRDCGuyfM42f4M3ir+NZ61He84t3OnQtM01AyjOyQzoPMqCVMKVdX1gGg
vnG2g+0e9SK+GqR7Ji8/SF1uOzNlgBLhD+2dpMOasdj0znJzVXIFTv3u0QJiccEY6AA7OTAVi3BP
VZYMBmOHIIqI26lxNgW3f6BXqYTGF2y4ur3iSSw3BSzcVuf5bbTvDMdH5sBBSR61/XHPiuOOoMJ6
wlJDmreXtYf+OMRFFsScKhiK1rYxVPc/U3wKdPhhNU5uguu/3ArnO+QbQhDW+v0QK25UaYot/F3p
ETKrEZMwxkh12ZHkColcnxj3QJ7Pe3hF0rdk3dYSkQD8Y8B1ihkavAAklzO1TW1md7i/F7OqfX6G
3ggtBos+ZNP2VqcKk8utlPrOL74GX4t0BbojxBr/xMBMkrjCYBhpwDwW4hcJKZH+7+pnEg3uB1Zq
5/oKQa9J/gcd2oUvz6z6m1iVnL9cZOouEQwxluIPfzGmZuNNTpLM5c1fX6/agEg83YjgapLKHhVX
6k0SCdqdXUDSf17o6feIaJ7jl5PCZB8lpNXDCKWwdC/GeLQLs8sfqa8mCY8DTEVeoOrALHlkdvXa
wqwyRz5+IOINwEtX/WJjHyiovzHFwyvsK3oTpNTLyMa7ri7WAXW2AGmyp7/UC+6Bz4XNDWsIvueD
0cLH4GqLm9mHFmvYAUJVFYUJ5AO8gZozyYWp0tJyQM580Y19ZoDKPFCmWCmncWKukCrjxJ+l6Yk6
5b/fHq6LO4z6NNODCh+EjUnNW6CiYFNSBKE8q83jwrVBfoYm4rq9bKn7eC9IHjD6bvCWj/9/4q9V
gFLyTy5keSz+XXFq94N7AYsOcZvIMvN6veLuEMXB0K4+UcDxK1ZYgVLD+78cHEQRpwN2i9EEt8p/
burf/1Uy8MszIRNSkDjPmvWlS1zLev0tgcU9CEcz2XWKiLZ0B0eh/WhuQ+FTRN7TU7fTPQqV78L8
ncZVgx8PW6z9DhMiuBU9ZXN3CPZw/8aocyOty/6TA6+THKC7FteZq4S0ib6HoxOZrqfEDNmUQFOu
GUdrF2UlumMMBfFlVmE7CShG/vA9j81eVEDySMFeZrbC+GakAnM5VxAwWQ1jPaSuNoMc1BQi4C4j
Ib9YrvDE1w8IQCpxWcapw5GDFKwkoaIs73z9wYB4aUcEQpOlBb/tcGOYD3YuT1Kx3AzuCnZ3Xfg4
C8cWKPJn7B6jT/TtsxePyTxsd7jeChAlhjaHpiKJe+oRoy4m6UJhai2ovhJRdCkXg5pae9JbHcU0
8W03T/ftlDnz3octUc+5PJZrFzc0A/jmsYaZIdjW/g5HhWMu4qnLkMTSCutqdxLJpIuaQfTW6dQK
YCQRJlXB1m0BoMtM00V1m7+DqGooA3tfGr5nor99Bm/RSTs7TDWIrYsGTjSawaFAWTySKSINxbWH
UlQGBZ+vzUJna9uwta1K6eVagjYrH33L6jS/6dl1NZKWoiGeQ08/e1rEWmqhOVTMa/zL8oGLf2Df
hEWBvxAu7NgiL68asP0F68IEybtfZndRVFQYYHt4K9d+TS8f2gXORPRNikLKi3XGK3NVAF6h8N+/
VY9915EBK6XbLWn2+tFOilQk8R/4+LOq1z6WFN+gft0KHnoz8ya8Cb1rEIiYc+GYrZnPlkF+Dj0d
58IPpddgfll7fctKvyNsA/ORwv6IVH5C5mK8YIGoMrfuu6Ri991QBzjBsyIzqQOuRjRQs9fNJGQM
H1ITSoBHke6f+1zBx+gWQzdS9yzJfPommNANlPxx3X5xOL8DhOpqvjDfk3mN0bPNT2J7xsKC9QBG
kNqJz4ShEVCh/GeUIfJSexA0kXhiVv0sH5SYBjtrXkqrSEy7prdE1y19SyuuKFcOL9oemKk/iB6e
Lu0KAqdjJmtAK5FFe7MhM+FX9iHL4zV5BBdjS6GUlQLiQfJNbr3ZQmm/JMS5p0gOUEEbUm8siO2T
Rfdz1KLsZPvvTjjgsrREZX0Vu6Qgh+RYjfZTNf2cMjvYgLVgVYtNhWYYrkEbeEEY3u3MYjHEj1cl
TRD3PA6UN9Z5D6SlO0fUZVWi6rzor1bA1+TYBVg8H+4VrMA6F3O06jTK5xO0HwRF+k3982xmmdea
cYuCI9LECWJFixlSmqVMMaU5oMi5fGDVseqZkQUfrbyDYTMZnakradfux+72hd/NTWV0NozZDp8b
pUnHP5RKCKqaU/IuGWCDKUndv6yMHWDVarYCxd+zPuj7WEuKrLFPw2xWpkuhlJ+YY0rzdWtI6mDd
GOgTGx/1G0UaIGkKRXSczIDnCJ2lJxSB9DrADESW+yoMJLmMQtDBM6SEavVyrtSB7ZL1KIGj7tQ1
XddMMgEyO/m4DhIwAeE+M60dsjehd2RMZRUOQttmLvn6ZHUFGaIbtWESVQ/89wkiU4OwwdMXWDrH
qsGe0U9raTweqJZh6YzIAo1kZqmZMgqAsiZiUHx97tPzbaT1xJ96i3aiN3+E0ha6druRICY27l7/
ZdGg1zaiXPIIKaYKbcFncuW1ILDpVYa3Lr6WC/yvzxFaXzvN9ZvMtfVhpAifzAmQTpi/XtrNSw+l
Qkxs2bnELUB22bo3voSaWZKa2yXrQB5C8pU3qZieYzeVg7J0YR7cDlmZZ/Gkj3mgXLqE7l+KRM0E
h4l0kee9PcJaeQ9ZeAaS5OMeUBsr4bt20WR4kW8Z1tcqEuSqJ4h/QX1P5ZfOvuJRK17HX/Q9S3+7
q9cvfht+rYNlY8ob00Kk680oYXtw/fA/yaD0/8yQDAhJfqbe7VBr5/5EjNGmGPpXmFchYhrfUcWA
HxfCqpiVqW7LP0PLM/25Vt1dQdW/l9kf0F1z6Ur6NNSHcW55yIawKPIfC5PIoPMBglllBwIOxz3V
Gsb2/uNRspT/xpymxe/q8I0bG/LNoq6b/ywciBNy87eg4ZTUmsru01Z25baYmV80gl3lOuQi7R2v
7WbaDMYvw3YkxctkYkc6PJBPkPeB18Hw3DRT16QZbAZA+O+x7z2/kfj3PMYmZNivly7BRM0y626p
1K+d8l94chYVybdeyMXVHSMyBQb+K9ArQLCdnNF4QFesBce546FloopVSvtDWAyVA9V3G52SHPok
nnwPdOnPxi4HuJwRliJc6nbYANIVprHURkXAItIJXu8oah88LzVhgbK00Ll5rUFRpr4zVb7CC6b6
jgC3kPCEjioamVKW613iMxhj8vjAUwxQUBR80ewo7WLTtI5aTeDJuKIdZmUEfO1GKqfcQYIQlNxH
Tz3f1vW222o+f10jYXJ2/lrQOQ16VufoCe/zYkBrVh6f/FrCOhxUCzSIcoZjlUF541NYSmmZHRgy
Ci5StzPNdY+cDDrV6ne7qqM+usYiIaHM5LnDJW455D+9lxxmc85aq4pojbhebYh9V/Ht2SIXwzj7
Ws0rRLuv1HL4orc1relrWw6pdJOCirL8EhXl8+ewpeKxqB90KqCUmNLpdh8yDyEpAlmjVMUxnF2H
HEEJz0Zs3sYDtv/1AyEBbBWewghyi7yOuUbEa6m15cTxpjNZj9MRyRDyF/F5/c5veAeuErjjBiic
bVUS+0EjCrkyNNztEjjljJ38OlV0leCjblhWHZInRfffIifWr2u2jp15+0sDbyZ+kK4xi7VaV4BA
tfHqOlRe5x7Fo2j2Ubr1RhsHnegAvD6vD18S7kfvu/tWzpctTpMsrMgWSyk7aQT4AqpMjCgux0qo
nkHnQfQ8HVImRKzHJkP/KO/Xd5jlmXk6YMfXJ3NLW3VX28H6GKNjXXxJy41QdfE+8JqbYQqJcjun
w7ofEIfGgU+ivT3eMAkuqkbg6BTa35KQN7hrxXMIXnrhWzEaZCDIr2iDo/03uh7p/Y06B4yYXXMq
ex62pBM+mTRU4odm+MDSWpnQO/JRTbNwq5agFxmRosaetNeTLANJH6vXVh3+s+xGgkgCNRVelxoV
cArGFNEGThoAMneoT1b8TgJISir0qMxqPIu3ckZsTXalSE1s6hjGDaTZ0GxDng/m1AG9Fl5PHKW5
24BMr62A/0BHrYGV/o/hAhnIAS4OCJQCXA3SjaqfNfEZ3Wle6WHqXJ3KA1ETQU54MxHS0BMgF2D/
exQeXgCspz46Fz2K2bNi6CHzrqonO7XD0svFKofkpYhfEJOSSYi1BDB1UQPOoXFxsKl60Gxc105F
k3I6KcceimC1JKG4woaz1oXE0D81OmLBowJO304CW4G7w0mf9RvWZ2IZ3D12NiuPbZ7cSvjuSQYV
rePhaLaBFkc+5LAowGncwJoZR0TUqfV2pRgcCg2DHVg1mjgvhM9w3PgG9emO/hUODQrxZ0KNPXA7
XcVONeNjat8zgMFbymt1VhAmgzqiWGknlr1YiW2G9D3Xec1CQBbGECJBhUPZAXpi2Obp4NdOnLDT
XYb03gS4epu7hqVTWfs8TawfrbVZO/wCcH1YM7dGAwKIb7//tcAUhb1jpXZVyYimyGy0m1DkrWn4
LE/q4LbprwJdlvjFEShiRZmwtIFSkklW3Pu+uhWFedDS87Zm7LCsufAkbFj2TymyHHtvUv8YJLo7
OfLPvjSXXXqGy7fETfDMjJ6p++MI4JvHeDVRS6P3WO0DUSMlPgWpdo4uoz8jDCLcKUyCTQpCw7w1
0oC1BZISGE4dXjhJrGwYsHCli15OvgQnbS/t4hEW1ffB5ZKmyeI/Odjm4WOdYb2cz6ch4J26H726
0JVjbSF5TXR1Jtg/7gEESihrTqq1Ts+Uatontrii62J7dTIua/ZJdMIgyqfB3sp+ILM+d/dY7imn
texmT+U4Z1yP2R4oXdX+HuBsFdrP0f5jYMZ5By3DqgjlT9yCHfK7qDE2QTbcZUdGwnmIXJMNrqd3
y1bxNZ4t9QqyNzRAULg1pvBki30289JJqLlUpj0D0YGQfVzdAxr+WSeXuMPpLc35l3Ri/ZE8YXCo
pk0hX6npC2zrFPiDxSngKaw42Tp1EVANtTWXngBrROaHTCq7r4v0RwoxKKJWlIT64WUDLwKyIm7q
fF15qj38Vo+jO0kT/WzOxLjAQkVbZEFroY0tYf7PGhETzdSSxejys+Ls/uFCE9PpS2jr4pdIUBJR
voVCD1FjcBR57TRibTc2954TEDxO1gdcbmhng+0JYHTpn+ct192+47vLyRYSOfZoZXKlU/cq+S+t
2F5ZFJ9g41dg0jMSAinMpdYjRej8EBgW/8h3iGVCNIdJoVA19ASvCL4I1ZilgvPb8zgPsS5ntsyx
T97sHom+gaTImaY7TjY3/Cz4sMG2CdgGbFWql+ZrGrkL4RG1Xg7lX7fsm6wjE3j0fb2qZHTJYC8q
PjK7HfvyrZgSfxVx5Aceoha+WFXJ3egRtkdC07DoY4orzDxfxQwFaZxUu/fzGfbMvMAqXpeitjaa
rhlmxjOegTl0lcDdqXjTnRjSQ1c9PcsOHj3IeopuJyHmMe9BkJH/cXk8+uHcLH8YIlqdhUdLNdFy
nmahr/VolRTaZWOkh08a1mWHbYlWxaKcV22LnpVcsB2kws5U/XLUVQrMteFNmYEQey14x3hGOTYg
smJOABmI8vs0o0hPj0iEUcyKxcDT67tNCW5iUz4Nd4Da79C46AkMr55y02Qo2PPXZPl6jmKX193e
NMTjBvi/KmVwBxP07u5wNhKm4TaU9yeNpzFlR248D+vRhjIy9HABMdfngLHwPjH9zWmb9Fh4/NIS
Xh/GXixj4qOqodrumZQdUef0Vnzxcnr7G2et8knNX/VMImnR/Zo8fLrjm012S5m3/yVmj24c7SAU
gCaXsati5DVXnbT2a4VYAc3LFKRdOh9PsnUedqtp0aCchJ9wSW1ig4UQ/CmgTnFF+hPNT1ev1YOR
SeGSfKvB1qZOXk6La5sHAMnNoLUR2MjIQ0pKzNX5UEKa7qRGtC7j4+i8yevLIUOCwO0PL5OQ4C7C
1CagUj5HB2b/GvvLN5gftzPJ9u7qmtgILeBWe2zFCFbggaigEW4OSMKFWpPWC+wyzqtBiTJ+mc8/
Avwr0kTJLCW+5p47F1mbXP7dxadXiQXTxnfCqlwQWRPF6UTUDIjWW65VKu7jJ4atCs+yR8R16KbP
xxRtlhirNVhYjnZMsrjXBlcvqD5wle/ntaJ44yvNybpk9WVRlePYe8Eo5qPLfyxIigICQI21Xzr3
amhcX1F5TZGBPjCdHYbTDA8npek3SLH9SLqXFKP9Eg52PEcFpQFPeUui6GFtC0FNiAajauvHPvre
mvq8UXjQ2atheGPtja2ODPNrPUpG4rWQOGHW8z3XyebsoSUdM+c6Eqq5+GGoBY8It36nyxbtgW7u
x0qPjelh78N5SQnpEdnIsd6OxUlP9Z1je54/g2iUSyCBKQipt06bwQPjnm9uqtuhVthxarp5ylpN
XMXrfycI/oLNW1wzPDbXf5c10gGnFQIG4Q3Hoyhy0h+4PT8XFYem9eI/DkcSKLEf50uaaNOh7AOS
PFvtQPAilJ59t8fsmM3yjQTyL5RUeuk9/SoBWKQFalY14UODHKKznd8qrNm3wqA0zuV+PX1+tiy2
O9jRz92KOsOtyev8w8NUkR8In5XRnijrJHl4S1K6o6WWlIBrYn3sAnD1cAEwFcLI25wIMEOQ2x1c
8UmfCScYZWsCh0FTSa4HtGfX4zp/4NJbykKYaghmFxYWe+ux/XZWw6/W7SKiSoRWweE6BDiCX3F7
EqsYQBdsp3xA9Nxv/jw4UMcVGfSXQQYYNpCYa3OmNsjjsOVx6F399YzOZsfPF/rgLtiWdJwQo/eO
fThMVLwJ4JeGz6HLTjANMLKgW5nFzDGv/ebmoi2WViIgRGtcB2Xjgw5GdP25zSJ/LIkj6S9LInSM
GMnxejB7lmS9Zo82RVVu2NbqGBcvgQlFhBAK0QtJG4ekHcCYEP7dat+dYGXatOwFn6YR1pEHg8Gt
r2QM3icQHq7PKudBz1VMLZJazvoGvxK8cp3W2wuYb67j6cv9jedbBy9A1d4QE2MKzpbN6qwI0BBg
ZOWHUv7FMKvFzCcXsPcNllPJJEXTooDTk6hIT/+ULmXQIxQwslkz/p2y+FeK6nBvP23cSDQXOYor
bRrhlOFdKh1aU+EMxNbdO70Ui4L029cutXRDk+MvK15L7soHTI+9C4FveMgaTUsLvqTPweBEQ0L0
p2mhvxlvttlLekcAX/caSeN9zsH7R9TZpMAm+VLJ0yre8y0X3gDX18gutDhC2QPD3XN+iiV2aYB+
782BOv3sBQwHCs4N/7w/RU6n0pZffyo/8IH9dTfPy9M9aAOwhzzQPcd8s3a+db3H3aGT6MTKiaKg
ffKXdmMuPoNcae9zutRB9yw54kF1NrCCeVwVUjHgrH8Hnu8IEWxw6XXI0zEkebpPBHYIGmGxfkpL
EP1opXzMUnzNUlCcdkq8Pyr2xIASiJvm4sM4CTV0vNCIMGIlp0WWxE5oHbxZSeqkioikyVC5oCpL
VnhghJvCsc1HlqxceJmh19bPuXcfhelL+p5vhmdRlpbpqXDQAASdix06bLSjHy//kwPIe24QVm8Q
has5CudXziRigGSXXXYLWyOfXnsz/o2JQGUuErBr0Hn0WExj8naDWUKhqMa3T4yoKS+CJ+dxIKAK
QLLSIcKS2yCipiCOHhYCy5GrNnqQoiNo92lgWfFQSLXRPzHwWgrahmMJaM5Bu4ZWkUuHfGYzeP2S
FwD8ypLuHGqUlJgn6Mozt79uJtZrRCr93XFP9zZU/IA79kQKDw+m+0LrYsnaYNQV7SuGnuMdG8gD
9u8ywDyuhhLwPkfkKBN4lxQxxtq8LhNQymNw33c7xKZa+O/yzeX9dDLzsAi+qWCM28I116ZTXb7Q
p7fAk9fFXA1Xgua/z7n1ZEYh8yB5rRvwDsR3G3pzgHpYmlLmtpx6JlXw1cPR0Sgfvbc+1hU5rRc+
SHS34UH8hKnUk5rCVpE4/SrRNnTfOK0OWLw6UQ7COYgLgWhjhLb7wkeM8QNiknRsU6p4qIef6Fp3
ffIPcuZSXU62ruRpifiR7JmF9EU7ZBypd2YcOKRwWXN9ukGsrpj93OK+mvvmcbL8uRzqm2fot/ED
gINw+PfRT/iAKsDG8/yHAipTs2iWd1nYB8/6Yx7KW74lHbwVQXLnT1dgQiW2g2b9ci39l8OV2PAG
sXxH6kLGfMyx+RplNyraY86G/ndv5EmbJG/undEBW/J/ogp1+JyRyt5JmzuDuop8itatUk+2ljro
o4wiuzCt6Ucil+p/zGl9/mO5XTc0Zt6CIw3M87abtca1e3ysgxHk5lQgIwn9YRxY0QII0o5op0+k
Jycug/TXKeVUnmFM3WmQIIgIn2uU2lHlXe/jPCpkWezKbWoyLeW7VZGLM0EdqQwzsbNEIK0GkiAC
N0keH0lMdi4Gwztrrf0zH3TUkEUvDmw6UPOBH8pInX+JtAwz98/+Yd/zoVleBdtOpRQiIt1bP+Tj
4yzLpjOlp5ZRdWw9P1HdoaIWf9x2Is4CY26FgbY0cWLLXN51oT4mQIU0lAojEnLBYQMiYE+CVpR/
Jz741L6pfo1jUk+pMxvKBPg2r7avj8AYnWtIzA22nnx8+0u706WKn+LA9oMYBae3MDM2AN2AuojC
2MuYfotga02R26ahUbXhcamkqirxWjfYt7duoJIutWrpE8/VCS/7+f/2LfUIjJx6pwZ/1h/38+78
WfXeK1OkKf0cxOQdnz/emx/A5e/GL9lUnBVsglvxKDWzpnz91YAzigOqKR+9vlxdsCugeG1l4MZ+
cW2fv9XHLkFVpDi9KBL11NXC3uHzlJNVWT34lZrSLGJojbwr5G3jmIZJJhQz6NFpCteW1TBqc6wd
Z2o2fOWPi1OJlmjM1A/LaR3TMa8aOqf7zNGeRGU20qXXI9hKEkcHzD4cHWXE7VVsEsCRg8DpM71B
IyGSvijG1znzx3NIWK/Sly2QbE9deCYDWhPx+e9j0xEykZcEF94LQ6J5Rq1rB6fKo6id8+vHZEuq
9BVFGJmOr/lCgl6JTYlx6toQmRUhQJU2j9s7a4oelhmGS2Vl6XR/4ez56Rn+l+W0GuVyo5HgrcCD
7G9xaFkXKPFARvdKX/X6K+mhUcAkzuShytEEW8HE7YuyBKBOjX3RGBgJpHhgXGWZVadaouWI2+7m
bp/whRMc/mNn4EKK8RfnEG+mKiRVBExtF/iE2L+XB3wxVva4yBQNxCRYuq6wIdkOLI9UnPaVvTFm
FUtJL6Afmjz4fa4haRccuIKH7qzVksnFjgqwlvMFLqeZksWldKVLXSlgiuTaObADvKGyIQK800PM
p7mZtEF0DnwMZ+y6aZ8jYCm7gKApqwEcxCInUs6ACOWYoGqyB9hXAcckeUsRpNEoVHJOOhMStLdf
spK25NgDTcp5CaZND7AjypnWM00uLef2fhd9fhQnGlMRWP5cNvI1FYYfaRCPOCZwenVy7EGLmdpv
rWUzq5bpKdDGe/MB87RtArYr+bCRGaVg5lE9U24biCVBP5k7+z6CpEabZZ6UuFJly0iQ5tBS/OaH
UjGtZ35TvS0vQLXray76wYzkddT79ezCWyXtJLf4S9AxpNEhmK+9HN5WgfIu+JFkvFkGt+VUYgS9
e7Q1JIzoRKxNNIhaUJ3QSHtW8HlalyRSRhbJIDfjIJuBWIvpbJGKcNVNsAMrqgcKYZU1JThKAERa
IBbzBoKQ93INrOB1K2EAakuZu0D50pfOKMWK+6EZOEpxOxcH4mhQ2zLcGsZzruMBxd6sDaObonR/
SeCLd2d8HwnRq7OgqWqan3YAhw6AGuiVAzOMng8yQUxDtBIsKDv7nxzdxXJ1K5iQin7N6C1Gax74
phfwhUOYrLOAA3DjALH2+7F/X9cv4FtVadRtVtgFGcnklcxdga/fOMEB5ScjB2f7/4hed/s2nlEX
7KAX2Vsw9i+vzVJjnDamFDLAvzxzkJNqEDQMtbGyIFrCCye2dND6wvCQjWXD8yJOksaid49/pZ3T
Ztp+KrViJho0KhsPJMBX2D6KMjmit8E3iFJ/Jd2MYMcrO5YdcmodcdteDMoaYt1a9zyJbNjyD/bU
L3u+7ABQKuPTSp8GmcLtbC9BipzQeUuKGrIQ6TgqlmHBG7xHahEU9YQtJ9DkSoUhb3/hwqUMazLw
z4oGu0ukCWxZKiY5WkrA9CqyiKSRIia2osApt438to6V7RI4JXd/XFvaRZtyAS7EfwtS8j36OLJ5
2ZShyqRSZhMy0bORYwCQV9F2HVUaqKwAr5LOQUDrIJ25yk7yGO9k6VwqT0Di2iE+pEaPw2mklACN
69/AO9Koh9DHB6T064m6FOfHUXXilLDQnftxOHrMXH8yAmqafN6BKJaLng0PHxrFQhF737CEuhYA
MGZBV+X5emI56yE4m4ay3amSNz5CZW1RlYtHMNyRsgmVnPzG92WC6W8XD2NIa7Nd8tSzGFMbB4B8
DwqLjmeBT6SSKO1EvtM2qtY1xCVCn1YDx6oO2UG1cWrDN9GeWcZnEFx4LbJh3zIbCmz1Q3DbtF8P
iZXGI6IzBxYRRiPPZbPgrOs3YB8DL6XrMGyKoq5FPDyor3Ic4HyRATu4e6096vTDm5QlEwwxLj7v
AEYAUWEf9baPRRFnTd6T0lUS85uQ95dJO9lYRlLeUR9hLUh6rqFZ8I+9rUDSjAsLdHvrpnB3uDHh
Y5f4kphvMiNpOVkDZS06nylOFKN7mXUhyzh/n5VMtZDaiEE+kLVF9EAbmL36yoXYlsUcVN/5YdQP
MplHJJFTPw9ynr1t3CTpHW3jdwYx9ZOBw/j1L/Udl+qsxc/5/VBSKei73+94gHTX9rTmHDE3LVsh
Rf3GzOC2zVD2h7ENug8wm9lFwpCoM0eqhnSsHpQieiejERZLttpXBiMscfyasLHOODpl/aI3WhZW
7iXC1K53dcDtzbmW/bLiyYKNcUCzPWCWWRGstevEOMfLLP0EqyKamvjhRL59csOHV4WSGzosGdgq
A9ac4T+2niqTgZV5ri5Ejj5dDW0+pcyuDx1KqXUpVLiUYUt6bCKesixyIb/oaOvrt7ZvxN+Z79bZ
RESIWbt2x+OrSHxYuCfceuhnCEKW7UvpHtv7+C9hCNUFKDKc7EFvncCTsk1+obJqLel/DLqprOhH
IpOksGmRUNWe30dm+LNfkgVga6Q+cgnftyRZ4flNHHrykhHZ1KR6ujY1yMIe5AYhM9ZK8uej60kr
U3jsJDlZOEC3LpwqS9EQNLl5QJwJoQgHzFKd7ekHvia5BFeW4VJW2dxfMRWOrXz+QKgp4pA/ZNPE
gLC/t1vdfy+MqIifNmTMYaxd6dnfU9OVlXEOmqhO7KUW7N5G/wtndbId0A/3wbtQNvhX0yminC8y
PI+6iEU3n6W5AVwuvmLT1ne0IULJncamxxBgM3l4+VcEJKYD2rQDPKGKCXo8fcl97yss6eRnZRfq
Y8K266IMxKYn0dPhIxsKjDZJE/TdfP+QOxistndnvYj6sszSWhjrSxQLExbTuK19eXJahD94jm9T
9M4Z6/LNVt/0Ss+5HeZL03tqkbUvyrSZl/jH8JDDY1HpcpBOby1NCI+Ek6jGHYybuzBI3AWdfeQp
gjDieNxrNiqiEPma3rurdv1rupIMYQE+182MV1f5Zd19NthgcjXX7ncjo+mvBv4sQDEBIkRrvHos
76uhvdbonulmc2A18Yx/RqxhtwBx8SdKytc01SdBjTJbnQxhwDmyZ5OdqH2gc1STbq3yioTOtDfW
rtPvC4CDu6xstSCvdvsnpBcfRTSpKyePd/4tKyyZQU4PBm56ZVJCNy/i8kkRvE0VY9CwKajtnyrL
+E4gPZtXDuMxdexjpfNUPFbB/6J2+tQSu8/+u+lS/S/T5OZKeFcjR8X0oLNeOLQAD5r1NMyfUG4c
/LFxpMJ9ITOMASbKPzQm+Xy6wI+zgYJVMgw/2fKhmPUSMxoTKWPTBrZ8LWNYT4pDS0qq5Ps7Ng7Z
2hb5DwF5K5dg2qev/uV0oy41Y1qny6R/ox7o4jNjGtaSaDYwXClIuj6V5deIR5VJVwsq+Id3EKd9
le0QKyO1WSd0Fqbtc6YqvPc6bXmj4H3K027Ov60h/oQ07Zzjw+xZKtpYgDABATFM71hGxlvrQBM8
vY9G7qXorR9FmSmRfMQ+LNFftOTLbTa2gfmfpYvdIP1Fgd/AsVdTy4xXGfCXB9kOWjRCjeHedDuT
ztNaF0Mxhi9oDVMS/wOS4kmoEmCCAE6izWhltBWB5J/s93dGKmTS3KCngiJT4QQiKMmKKIX5Hai5
mr4B+gergDLyzgLUoE/wsUO6pE+FcQP1O0bYlK9iLPX2tfq8558RLtwiGM7EKYt45Ra2hi0n/+Q8
l6QRSgxEvA7BYmbgwnlU7A7jxb15Q9s4f73JuOL6YoPfLAoDrDOrHWxw5YoKCILFYAxxgouyTVOD
cE4F+5acDL+kfagzytXq97YuCb/rDdEYJrGhAheWncVDFLD1dQS/717pMtRZ0iP8x1BUGVEKtPsh
tzVXTrHh00YewauNV+WeNrjfvajQWr3dUGRNaiVAjV4IrEEfwto6quUO584NpjrctdBRTgKXD9Ul
BAX2K4CJZu8bJMdU5bN6ZW0NVcvePZ6X0TqyPewuveDnpDBIdgGDVcyoTFQ378onPtjPlov/tVgr
mstgir+8JhPT5Q3lI1QoqeDJ7yG2ygHLA2DRzvRj7Td6TPSzU5i4+fGJGwr2eqjZkVVX1eZsF4/0
yk5ITVCKrZcKn4SiYcfoY7bEZDAMJDZpEGPCddCUDRkNcS7iOfXuG70Dy1QcN3xQXVVI7QUAu3dP
3IqG0aR9Ae7XbmoYkxTqgXHdgX0NYkTz7m1f9b+8e2IPYjQz/iatiORAdPauPY01tnTgWzTr+VHv
zKGdp6Hp9uMgoFXHPOATYHgSjQ61iapi6T4EZuEpPO9qFgSt0YBXaD2cCtNFuRfJFiJVARvAJVsD
CKgN1GNv2Jq0KhEofMTXRg2QFODSBbcxNSHbn7M7kyMOiaQKXIh0+ESRY76iSSd6Epc4Z5KCg7vT
2vTZdXYhc5rQcmQAB91kDdffgNfy16EKtIRyrU9p2iNegRJhH/0c7VeyXFCWDY8A7QAU2u4Ku7RT
svD7iU4FCfHCS/KLtm7xBSgTWY/A1mjSo22SNyjdWsHCFOM6z2j4U0wdsOfMpYVYYc52Ij5DcGTw
L3rjB4xtZdSvY0y5R9W+AUXlPTyTk2W/Bd2q5EER2o1DFAZztu/kX3p3p7K5HBYGV5KXhZNpW1/G
/PdWcPYlsX8BCkILY6NMIVqnMXTYs7jGBbpubToncB5lGOgxLYd5K6Kd7SXlYJSTC5WO02z2NKCg
dlYKeQdJz7Ak8V1QmlZuu9InKAh3A5usZOv9iGhVSlXV8Om/7OPigOmO2uSp6OM+m2h6yBkLUHpu
Zk9PEMXgb6nqMWY58NwBhSfBiB8g7ZofvR8ja09rwdVd8KHYrNuj0D/PxZehqPYeUm9LCvzNK2e1
LIJ2acK5Up1M5gpXYhGaxYtFlj1XmlMjmWAw5Cs1vyt9bZSkjXp/OJfAGCjtANwKp064n0vyr+bE
kN9o5lOxRUShVL8A06dwOKVAjfthm+g48R/TSA9hsNkdtuUMjCBbooQQn141vO+EhQqGlB6wXdLQ
etcefx1gS6X0O1G4BMtGXTJvG87l+6fR+kYOl22HKzFxxtSZSZCb0yWTFmpjznFhi00830Sg2XqR
NoDUgV/VHPqfuRR7XmED4p3mJtAwQ4fYwQciNJ2XJt8nZL/GXoC425cMYeCIBSfh7NhF9EKAoD+d
58HJ+M8bgzKXQTFYFs0cWtEeCNPa/YIV4o3rvP7FKUh7D/0L0+m2lHpN5NeZU19LBz5qHcdY19u/
jpFUe85cNUWTWDCNtvi0V02rQpyTUmrlil9Ne0dhExVV58gVoSLpcYqHsVEKdoLklhuL6FKJhg9v
wnQkZMv7lSzUrZYXutoKT69aUMwT/I+e89KasFuByS77HoQJh4ZDmQEq+5dcPedjobwKHlCoJYAn
DmXkta0vKJCex7AH/Zi0cnvQ0ms5KBjbm8ZpR7+BUEBL3hqrrMtsuRc9Nq2TK+koK7YRdMV7R+nZ
UMWXU+WB1DAPm6I+zosGkzPTKFkAzA9Ti9w7ekxdO3S9AlWPtQAG9wDoM7IyLAN+f0gpmFE2rEKi
139xwz+zqXhAWnUUKUPDiIuVsh/5G7WDNic53Hg3sbujH9CNHjupXTJrmam911R80cqqNhNftzqF
t+2x1UN3UPCPNo/78qJ/Qt7AflHzbFxnKUKalAAKD2nRxNv9tD6FDEZbejMNpX4CcCnPzhog29e6
jUaIjJ9yIWFwdxmkeJn9idODFBSlDHyJaaUF5a1gDkHQdEdc+YVIHBL1ZRr+O/byaCO1xjC2fsAN
p8HTRCLi837Td+lRlPx/KK18M8Hrphs8fMC4rrm5R+v0LoHB3ACBTFe3z6J20kEvhLaCT6f+SWg+
h/7IoOPUt+3YmzwSQtrTGllPcF5kcYN64Q/6xbnsnlXHpmS9wisW54peqjytAGvRbsCW8NuG2cVZ
M3CtFnT9dYGUJFUYuKnW+QyY5pQbi7G+pw7C6LByLEvQ54qHeR42Mi0K3DYr9F4ZolBlt+i0I9ld
tWzW1JRo3XtpbQbc8yn4EzJCYhAFz+yhcmaOmKvdqsWzMEecFLbCouRK974dSQJQRJZjF42jc2hh
9GEop2rccbw89CJQcnjiksaC0709yrbRzUqQC6lFLssz5U3VB/aD7PhQg1P88b14apKtEXVusVyG
H7Yf6D1p1uxx91ikKbqEMtT9p3M5kQyaC8psRfTGs968gXBSOkn1T+/V179hwjL1jajxxVSErVee
5yz6S75MieaaAbnOZNbpNGdYFn/nDhlhKC/BL4ntp1QzjQItkmfXI9W65hzP+0Ame9VX903hzT5u
akL4C1jTNOXMvAoC08jb80bux7gb7k7S8En1LOFr4mtEwGSbN+l6EulwitOlqOVW5UJWwwyZXci9
Ldo3dt0fjD3VXwMWCAt30YCftx2pQUMSh52oU01ZhJWUkSxgsCgWA32Mu0djHvILidbgCzZQyv80
Kc/pCrnXy/grCymfXf+U+JKl5ksMEDn/CtHZQi12vQVrfV7AeMJ9DDj3ELKC/LiLPlEZvFCv/Vu8
W1GHnUap7kLMgbaAan/HO3JV3uX7uUPezNKw7cp3TA/2n5c6SL1GLZddUAHj2cVXsBuadBwOSRKZ
0w7wW2Uhy4v638lwWRbr7RBLIHhOoc0iYH04JydFP8+CWFezPqM7rZiyLCv6DYp+x3Gv7wggxt1U
aNO/7v/kNME86fNrQ7DLnYuUi4wGn6AigDDtptsxJMzN9WOwnSpoiRvYh+fUjOUm2oyWe/9GHu7N
rRpThi0EtKaX+ApXs8s4ltM7470UL6oTLyNDIc8AB8oWZF2PQ40WvOcjFdf4gQC0jrmobo3Q7T3p
BJmGA4KByzU9ohv1rM32F70XEVjhHcbvd4RJ1HvQfCv7ZszvxjYolnickTgsffnqmKk6EuQN0eGK
JGD3WSodjvtNYXCphl26UIx6PFumCEzdbxGyc0foIWNuCtyVqxUISO//DTy3K9hxkLJcv9EmK8ZB
3g+QmC7PDV2BCAt0zcIEx9VTGUN/U6LcOeOyWVHE/gLnl+grqOgGgHlIFYY/zxhGcKmB5nGdgg8i
HbuMFbkUeDsBTyihi06du3DvhmvjtkAAncSScEw34TwVkqs3C31zAyXVsIBFNwb/aE6JYG2ZFKIs
SByo36DQOwWchkWm4Ws17UT9VCRZ6WFZW/sZDemR2DvUyeIE4wlqrgj+af1Bt/1WwP0KgdUJbbHR
F/u5E/CMGCuxniPw+sdVCdGw8YnLbtuFxvTKOA1Q9alhBq8+tf8Sk7Lf0dx65xdxOVjHeAwFvLH2
h8WG6zC/CDe8bccMUFwJet9oXNuf+RpeaGSiQoN25nsA0r7RIoekCkzE8I4S7WYh5X2K1kNFOUv2
txmDe7TE8mbyzVvcC4O1q6V3sCQZNFn+7HF1RBeIRVcaZE5ye0/msu0azcr3BVdiDs4iLYhmsB9p
BGVPSbbO6QiKa4MTgayF44iioS8daRiNTEU1MMKIF584gVHQQMO99vEHtf+9YzNKLo0lJr7Rz4tS
TBHb81ZUNlc4PeEvkDM0vJTmQ4AY5KjYnFl01tEio6gpKHGSIeXGu+YzBTbhdKfkSdqP0Lt4c0Ae
IwkdzHgohBOCluQUcXf5nOk+O9sUcbIBJ6zpmXQQIhyOtcVzusR1x8Y7xVvc0Yx+vT6v2WM1dfIj
rkkb+zlEU0kQ66wip7wq6ANBM51Gz38e4sFImvNTf8UqmhtowwqVuyOlI6kc8Hnz3OSQtZC2K7jf
upBRFxAWj22Utg2pLdT2yXZvO2+ZyPG8Epzi2pLUDJgbSBxpWdgr3nXx0aCMScDea02VFosRQ4X3
r0LBkYqyulRHStxeCUp1EnXB+r5gJkhFPnbWRYnQsR4KoToJ171qVcBmnUpXPcldwMjaV1zB6YQM
5UUbzs+6nWhy5bs8iDsAaPM6wZ5Mn7F/wsLgVpGYVxMnnYvNJ75H2QCF3lp5ldnujqaRCs8vwFrS
QdKJ68NmjJN5CzDOmtMSsYumCksHGIZc7wR8sBX7k1Ventsp1zAxPHnq50nZBJ45EpeELLAvP+3E
jGt4GkXM1KAmUtIKKf56LkXN5pa+XmjKolF0JW4xbVWSEY5PFXGLQS7OZSy6mlh8VAq3Kw6sy4yq
Px3SXvF258bSTJXh8Nj24AXJDz53i7ZhLMVNBykFptqPv9V4oAJJ06V6BycaQAsWZvubtrcLRGqx
OhZ7oU2olWB+79EohXIddSm51mq3+BeDpB2hjrUNS/PwudLjk+MCGiem59Q/8/b3krKrg60MHvY5
w4FWocCNs6/9r8q9TEPMbltN7Eb4pR78HBY0WO/xQJPNWCXRXoaLsrX0tmh/6F/zqcZdoGENk2TJ
CzyoXONGAQQwcvB5UP2gZQeaGod4DQRUKV3/94qPz6y5d1X8QEF1qCcQefK3YdPlRJVWhRZfv8/q
TwAWHLObVaG/+add1qxbObRH0LCosW2KKrcbEg7zvGKxFHnqf5ZQLNlt9AiOygrWxWLjExlM46+X
ZsCjs18J9WgiJSqjqxzKRpiiqzc0CTihyTwClK/WpEshcsx2qlXs1cFbRFxpfvSM9qsixSMQY5Jb
2/mnk52V1WzS5W84lz4tRRRNU0e06R7aHQjDN0t91i5Yf/7NfozTWAxRueV4fBKSBXxwsmU+xGFm
COPqq8O7TdSKtipinLQfN/uj+8jqDQ5qsu82fQZD92hQuOorc26cszN+V0Blm4/kXmG93cfnlpQi
BP6UkQX71XN6nm85iCvLfqp9/kBsqmjsu8P3rN+M7NKzlad5hGOd2lJf54XwZ7uOSX/T3bLRw+Cg
wug0i9Z2Xo8rY8u745AUQKwiBEvwcKEvzj1GFnEdVv4CPHtxYlfWStFqRApTczKbcfyfpTbD5M8T
05ICTfXDmxwe2/IsAUwgAj5iHErUYOlEUq8iXVtBJdFxeUtjQgvmS92l4ofDH/JPOR4xo8N0/4Wx
VrVjjQxZc+akSIf4iXAoM7FAXXDT+Dll6EXUYkH1GuB7EKaJEvglj9ZFXujKERK6r1k8JtMCYaf6
ec/XS4QCqbjDChEe6XNegHzOUAXXOTaCg03y7DHQaF9FEu27APAIT9WWlAjhMoWBVym8JEyjkHIU
hOSVw9Hj9ukNoACWcitDSHDJdoyDWCovzDKzoZRDhGDggVY6sMNTamaFjsN+0pbVeuvCkXV6ZFEj
0EaN3ixRtcXBWphOzV77FBAocQjEzUp2CLKjDGjs1nCszZTGOHgzKerVoXUK9Td4N+oR50Qgt4nR
tBdE2AM1H6uFC1BBiwqmILKZvRMYoOskcV1b/epp/CVdIF5YMxV/WzMCI3GdyXqBSA5CutmfZtsN
WN89uMiNWD0ncwsBxeSMXvzPIKAvfQIgGq7YRFDDWoizhHuHM+TE6er57CgtTnUtpSplsQA9lOZk
kSz7ZJL+ynSc3aewFMtxbpPT/9TWt2Uo0rYUQiJZuSRI54H66FUAfn6TxDJQq/XsYTLGapgTajlT
IDCqndZTu3nPFVQYsGNVka6RzC4wn/KA/vo1ibRP42TSWAeh+4u7rsY5jG9Fp0p8lCb2YdRoeVA2
+gNd6O+Iqgc917HJ0YkSs7mftMu7GlL5npX+gnNGPiswclSrMBIyoNc/SYWzFgpMtMO1QtwhgS8r
UpOsprdlClgKTFgkEwJQOpDaJ+QMvnm3A2qMfW5HylyeJZgJ7q2fgnLIJU43JyYZOThAoog63GOc
YsgsFbsdPFAbh1XFWduZoqbc4E4xH3gqa3iaiuAlj/Xw5qc6yQRLmvdmq56uc4GmvNN/nMwHmNna
n5n7RL1O6itiTxXo7CJd44pUkk6wJRp3xPGz8V15mGptVjcbBvZ77COhhG9Yv16SBHmeeb4Iuk/z
JDlkCZAHxoaC9rP5MQzZ72++H61JzPD4VZHMRer3axDoVYgVKZvI5Z0djlT06ew9rojmNjVnx/vU
aDdrBB6z/b7bXEhPWKrLUCierLKvyiFriSyXLXmat0jwp/qN2dRiUSc1ZSku15Sg0jLgpHGn8UFP
Hkk4xpxgkWZg6bv02p/P6eTAexxyfOqWMUwQhqp2gHKsyznNV3NFcxHSHgKGvV7fLTe4U88cQ9fT
b+mL/l8YMVTfbyMj4bUxredBAfdf+jjX21lyRfSSdFL/g4ghqEps/6ZJ2SE7df053LZUUNLaUKw1
UIbLJnsOr6d6M4ojWrKrhQDu5QWjhDObJm0alrLtu1pQmQ+2fIejB8mjakTBvlOOXwlviQ44maiB
Cx8ih2Bw/yax7ihPgl411jJGzLYVVke3tXPiNp4knj3u6E5DRGUnv8nNYK5yqefGU93XmLlnfCw1
IC8hodLx2gQr4tMdwoGUIMDIDP9lLbFPkYLeeCumFLtObHlbdgioxWYuJObHVhPNqaDgzbgadad8
jzazLEzsiOAZmOcIjRr0GffCrGcncSOrs6Kn80ExTiukf6iiEstXGHcnlHnPHhyj3BPgPF9iGxpv
pH+abJaA7hyDS7/XnvTAl3Psw2ft0wqGIqdoE2jbR8QAVONgp0g0xaHhq5cBXxhEl0wESIJQKyBi
t6e9tiginFCLOk0TLVjx1KyYg3ygo3McPIqyWyU2NMjR+g4pUejKlLyGp1AiTCR6qkNejEmDUdc9
Pbn4cSY6B+jQjIrGdqsnot9KZRyaOOotc/7k0UXiYUDvb3s9zvjUtSWiMCBLbVrqe2K4Px+zQwtk
f9cbmAkijytVDJ9spW7UBEggUH7s3vMoSKtOf4wXDsIdaiyvK7tBgVORsILZPPoxTa9EXQqjoqkk
jnLpmZgjjTGdf8G5dQAK0U3q1XHYdDmNkY7TdNQ3wgAPSEP3LU48vuc26n1IPI6/MdKpVhkRzgeQ
xvI3Lr83XYoUlODSXZBtfM8HKyNLO8BOgUiHh0oUZ0CI6SJsxCik0LzU+sGBqMxLajy/CkTXY6Fm
YLg6A6bbhvWbHHve2LhcwA1/c3o901sUt4xwoyuAcaD7WDH+VM3LC1gz/1q8DdDbGQgkXJMBLNve
Gt6DIr/fQTprfY4I8k+Rt5NWoJjvfLa17bUJsEVMZHmaHVuvMzXSIfh85eKqCUDnRgNFsTvidFy8
Nt4f/Nx9Gu3dcPGi09woC6VraiRPv2nhfZ9kIhMGNfJmFt1N3t+Y78ZHIvMzuem/4t+N4oHLfiAV
opIfG12xUqEV1b3/dwDlv4UgCAh0lY8w5zJttjcNxLeqblpwAn0kYYEGEZPeXlN9lv/PSHbDr1oD
PbLICuEJg9aoM9Zd8wS0Z/YuArzng6yOF89dEsv2tnOs7I/9LvNxLyqyDv2XqqEG2njb26j8ds8n
PvLhpcZoiOtRX5FEsXSsTaMmAdUj0rYHfJMFywFlHfCCiU7208fyXyDHP/rhTAA1r6K8nLCfRinq
nxItxzpt4gHmCHFGNVoDtf4oMwtsbmjUB/L+taqTmCPcgYGWayPBeBCggxlXjjlHA8jcHLxNutef
X92Ed3f9m6ucV2AEzo2pYRk2EGBawfZh04FW2gxbPey4KrteGqxFbbavIcT6mQhGl7OntDFnHOcT
s6G1jncCvbvXqcnZRM4bWs7Ds6J6VwSrpmrkTP8aS3/tBi/gmco4LlPXULjtrUaWZnKWM/hJKN9G
MNtcuwtnMj7EBnDL//Mln24d+3hzhjt7ctUxAsg0FAmH6v4cgtnZWfGXFMSEV+b7IGWgHd+NOyaa
HszAreawMQ+KjWb3/wVHYeDVq07EDr7rCDtKS6y2JanPT1FpAKCjd6px5UPHxFDl3jnOQOOCqnT8
8dkjBIQXWsorhVCKpHxaSxvioLsEpMrg+nOt99XEcP9GTJXYKv4yoDUV9KZYckQInuPAuXlGEl46
+HZqkn4WQqxJFQghqmVSAspheY/KLzgVcP6k50bpCW/kNPQ03V6J9oq+4WTuIoHvh5ah8GXmGkHs
/gQSNLvlKVml3Ifcif6fDTlbS7grrZPUcwGJYQkC6h8153J7FABa+9CSOdI6U0IrI3fYP0op2aPB
j2Fd1VFng8drJAHhj4F/wOiNcnOjZ7voAH4iKXM5FhM4rdEH9Rt7WNWos/lMWygp2q3wOHBI1s3J
1UvKdA25hQl9SAqXoegsIVCksMCuIWBYRahiRW33tqNHdLuRsN9OBgx765jMbMtwx1FXYgADt7Y3
hNCUYpd9Q8m/xKS+Fbx0uPqwV/45TK0ifSP8ivoBPnLJvtWZsbC+7VB18QN/XUYxTurmSOwpsEZM
SzmTAlkLkO7s7hCcQYOvfMGhF+utwpwF+g8GB4vP1pFa6COX2Y/fLs0aMRBiDQIhulAXx3hVNWvb
pQQDqn9kdqDxJd4daJpDvfRAsQkk8v7Ll2cvdf1UezcXZGPvZg/2mQr+7gtO6X2DCGoME1ZcU28z
gcXAqMr5Vqf3FlolquTu4CR+KzWCp04rAYJRw4k1TxePSpotqdwxkojL7Zq4prcRafkiuFURK3uG
a4zwrHBBRcrg4JsC9xCtME6WMWLtKEzSLm+XZ4UdnPn2MTzbastkTi6fQW7GVe7BGmb+e2bka0o8
VwLkJA/LD07LzPUMkKmEIiApCnFGutGoMplfxy74BEpZ+obTGseVBEq8RMFZJXfCLDelx9eHEHg7
dQjhjn1N9Fc5dmwb/LrKcRQasSHaU0sdqKLBcipblsipfti+Tu4VXbw3V2CS5f80fPTYhD4WZWFF
hIZNn77SevHYS2spK2P8I+pyqGUQ/je3ORLa4kfuB1R43uJo8XnQVLx0tpII20UnOwUhz0fN7q9f
PcYjSaCiOdZvKKVpdGqNieXZx1Age0HVrqOiVdg2RR8ezOs0xYnZImzRmifMXEZdWesAnfoLqVAV
ZLdvM6pjsKLW+xWccRElH+gm1DDRu7JjomF8pE4EB++bl24T+ggWgOhn6IKmez3OkUNra/L/ve1o
lF2gLBagNWAVsuFDz+8QnOW6koxprlLsTCxRk8zl7ltw3RhJxHCDfE0UfXnPUc3uakRev19BS3nz
Pj9vLQQr/Fm6KyJjr5tjH1eZ2q+MRmr79NBW8v/1+0LAe5Jz6jGbsamskOh75viW5MdIKXlXkBFC
SjSEx0rig2eY+mQczMNPIyBzboBJOP3QBNLqFJRBMqgUqkH2dzuHTdwBqMMd18FPBJuLwSKKLiI7
y1YRTQEJ8Hvmi0jqzIfbY0m5shrqFgZsKbq0yluQSIfLzbnf5X4mKXZWNUZ7iq1/Ujo2S/bi8EAL
kusfjkFElBOCvVDumsYUXJzG8D+LYhx4ffVXDjGHzVgoO2aCX9nZd4k1Lf/xyvWoVOoFjZxyPLMC
w+VW4YA1BUqSePKvOKR4dM3Di8gJC+NPwadfRqizC/hPrUqX9IV+tc7vO7r1xqVe8Y1j63I9PPpL
fdUzchavTNtL6ouRtNB2pf7zte8NBZ3tCYjZ7sgG/w+sMOdZPLxSiQo1L3gawrxn+4yFpSE6Xkac
P6ZMa9qJsyX8C7223csd6y6k99VzzNGgdR/CGnd66njCbq4MY4iinN1QoDWOqinLyOYQ6gAmyUPg
O24y0oSaq6lU7lqXQJA3HX4LPgY5BuMFp4hpkLeROhnRY0rn1VWK5ZOi60tnH8KHHro1XEUOvkng
gNIVRyfV2yxNblZ9299EmluS914TOjw6m5vjojJTUENQ1AWjwLLceQIaXYGyEBJDqHGSwineTfMC
aG8oBH7yPhHQzy787mILxS/NFMB9oapQMBWk0Qez3eF4LAFl+s5oP4/raZrx6k/SYfCpAetxpzCo
5QJGFdO0wJe93bVmIkafbyr9i4EZhNxgxbfKXmmGKsO5wG59M/aPrlx3Vl+RKCM+sksR56kKRhkF
+4jTd9k/Gf4iFn67UjWRbMMKZjA1BE/rk+6S8gxpfSiu1qShDjKlKF+bkaxmi2Ag6ygJ8b4EwQ5X
wgpDSSVlohM7d4ArFRIU3OB4JoXIPfUYOmiysFgVQ4eWHsONG7h2dmUtohnvfw22bwIh6m2ZYrTX
rJ/Jcu5fBxReZhuR+PvmkHzSyZf9LprZwm2aMW7aFS3Fudsh/KlfbWm+tyHX2h7iY9defj8g5TOU
0y0HBl1nn2TYS66NdQKOv9UkIj1lLSOsHSZH5EsuG39ETCE2tAQjSxUHWYSS4hzn6F1AQGW4HDBn
t7VBIUJ0crNv8P5OEUWO5vN53QRhxhXtZAYkcM9GcDR5NdyLZUSVOiFIuc7bI+4jm/Y5DsJdVUea
QsEjRh9Wc0iJbQOrtYLoDol9zVRN0f8oXfYwNobYovt1Mb+eHSXIdSnJ5D8TH1NKUNKHKY/xktKs
JblYUVxAQW1pVkLWl5MID2x9Yd+3IGeuyFieqW6D/U5oDhgeeDiZIpVJ7UOb+eNMoRQWq+8gMkln
uMZClfA4/R+Wo8KjFk+itcuj8OxvIxffwHsp3J58wMaTnxecPAnZ6SDVRIv0Wgm4IeAX8Q7QKDFn
ZXs341LI4LGe0Eds4jPj+o2dq39OLDHzgGqX0HsQQ2Lph+Wqu+1GA5d8T/t/hdWMRm6GwPDF4Y64
sVWblz+tEpH9irkwm4eYJGEMePCWua9gG+BgR0hH1eY4LdvtL0DCXNz650G8rq6bW0F8jt7VzaeV
hOJpBjQmp0aauwwDPl8+fzNqrGmqdxllcCSdAvr/VEn6Vw3D+MiVk4mYMg7m/pH2ZNgcATmadGY5
qHiS2XxmTCOZTqsF1VMuV23XvTsrD+QoaPXFEU8iSVk8S2UN1DaQo+ebc+PKdk6Fc3UPDj035IYs
Cl4eqq2qpuuyWuTEMgbFI4TW/cPyRRfNbf1zoSnb7bZlPTgcZsEp+zDHSVBw0vXKufbJenFL9wJe
xsb6jfTwetSSlUxHP31vthxrcutq2z/BQhOYuWB9zTu3Noh52K73O46XaVvWviTX07zot3uYM9d2
UD+sw5mIgVmKBGwiHicfNluseGct4qChMU9vCii076I6sPRiAIQRGmwi450rYamf0eqcO8qOzHOH
mQyU5jwfyKZwTQB8OvsPIrBkJKAIC9slxGMxbzYe1x49iiC4IjLjY0thGP3u1eI3ZzBOW3pDX0Yn
W2d2hAKhI9dIFFb0xb/rRsqSSbw10l5wIYPDBuwPnXAL2/N5Ntq/3ajX8IhZ/NL65ADIQ2PqRs/r
4zdju8PZD+tNnO6rRARBC5sS/zmAp50HpRrmfi3A5+l4rJ3b/7ZjIPB2ud2UD0gbl7h7vwhgaW3+
dPWz0RrJ9VbAH0PIhffVX3W3twCSA7gueUh9hA5Ogdhh+KoyN8QrktgSXJKoqMp0CaVV9s6xxQFj
HxeVkavGengrZnyuKc0ZjEX3sOeNYH++FyFwuYpsXJyvrxAWkOVuFJnlMm1FDp5LUdkwi3U78+q1
rrCfEh3iRxuIK6m3BH5d2EtliB/9SNrG7bfYZKVGTmTBwpWrpfIxXVmVSONfBYJB6gkuZMvVz6S8
4rF661nQ4CS1PB7Z1dXv7bI9wjsyH3pJiUPvYx2bTptoMJN1rmXClj7AuBSd+zCnUr72YS1Pvn+P
/fiAMxok2GLIN4K6vhb0CePgPlVvmcFz3SHAHk3AUiIMd3HA/d3aygdxsjtwsDHE+tvQNlTwe8pj
zg6RuHRVxSW/RHTHq4NQlRojaUVSnperG+ohpj+lX8zkZjQocIIzRCQriQ+gNAEefewT1bh815V1
MD5/5BhEQuOpx2R1XxfFv7wKV5FYFUWUAF8GKXFSVOcHB6dBZivDu6evlAoHr5r2S8kP4Abj/3uX
sj02pr6if7s1jctlCHPc7g1cQmJUQPrP1oTHgduzikTeXoZUfrj8rlNZOslhdKE3xIX6dL2OtHbp
3spv2IECGa7iu7Zz6ZcILiBnokwAdIaEY2eyptd6ZSuD/qbyZBg92SrzNkE6yBtQlMQJfOwTrk0Z
bDBr9d+oXNAkUHLX0MZrmxB9KHtCIj2w1F1SPdNtZ1CQf09GDzYV5kCEAJhvDBpGl4jqPMpsIKxe
piFrUgiyc3EkHTYZzt6YCR0VtN69ONADiDFFr+2zTl3eRcMmReMc0xVmrX48hBOR+b8IWP+hD3s2
0WkLNABwP3x0vzEleC1PrDgq1lXa8msM5Uoeav5IBOgDo56uXp4R+cskYyN05CEVoD0u3NWXjpp5
C3zqRmV4KO6fIx5M02FIUH1ULONWtpTMcVHI17FINzTJE1/UrvHF/w00bRGCR5sPmWAO6lFSb18P
MiQcKOwxpphXV23cnsJSFDcmfkYAsAYvAbt24MwQBqu578l+C2ZNnMEgL/lV8uj18Jj9bSw+9N2m
lyJvU19YXWpYS6LwRs4iJtAEPfT7xBnx0hc6uM8linvb4kv/+mY4aPuZ2JiyiicSpm3QI+F23AT5
7WxKFoIeh80BlX+Y3vp5YozjxbcC9EA+o20a3nVeEwbRIIXxqt7685KQwq57WBW9th4VwpDO865a
rMP62Ck2cS+tC37qZ/weZkS1MG3dtPb85ZjAYvF9Z4i9X8NHU9RwUhhrJJKbvfzCEbdIZePxxTLl
mSV4RqwQ3EtiSTCZB++eOWbfLzsNpT46Js0NYD9iSlSwL300tAC2L6EI7uW71KVQ0bskrN69yNUJ
7ZjzjH+U3JFjqedjWIgmILDQpeCvKRgl8uOd+DxCN1n3HZHQC+YG98ubBQUFjbhbA/rJbwizQYJh
VLQBLGKhRsFab6i8OE8mXjz2ApT798xeYSlSgby+TseEWYU2Evt609t47WltLzMXSGkHlgodIYtT
eeYIigCxUboguEKfwCUuSWVuii4dObJKKr9gGzmSyVcoHOyjmxlZc8JR5O8qH5h1Ggm3ZjTMTVmf
0GU8FyDYURk2Sc/nilI523HkX16r6CvYrddS8UXjGBYC05U+AWKjE33kSuKXMEgxUqZPOd3+424c
fDObOzeFfSDieCplGufj9n2nLrxBB5LIxnHrkLQCtg33hV/BU6taiFBPW85vwJk+V3pp5YhIpFbN
Qg1BE/DJFwDmLkuoqxQVPnzCPMqhDgF4kwo9yEc5LeKU6eR/qplKjDGI3fzRChIEyA1JsUaj1hUW
VCtn35uznQ/h+spaXcj5DL2H9iChvfgx7EgQ22MPRSUswPmQmvAAK/oHNNZjp9EVwUEvs7BXu3lD
cf076G/QN0WGwOSQwpkLotp5tChAzDLwdOQKmMnFUgEZ27O7YKSZcacQaxWq3XLi/GnBnBIzGK7O
fywVhZhgNjXIG8SAK9O8pTr54ymt2BYRSAlgWUMgLMLi3a8CDH9+y/1sL3bzmyaQ4lqRoUNxrwIl
cOWX0onl1/mSQCEb96O3X60Z4XbjhrSKbpJbtKxfifNRjKvA4Tc+nQcivFJBymP2Pm69WQMGBdTu
MC63h8vFyJlQuQlTf2Ivi1a2oN6QEH9nLsTUs7YZTZITBuFaXo3PoEiEnZ5uEjYB0QUgfXc8TjTy
H+ULFCR//A3pQMrckp4Z8sZN5L5bRNARvYopzeiEKhqxUNjEVzDVMOe1mBUZK7bxwUG/tNoT4u+L
ovQ3bFim781POIODceWzwb5F3/NZScNyp73ZyK6hPgv8lrT4y/1a22kH1ky8DILZZU3rWT5pTwaS
4QAeuGBDjI4ssqUqBd5w/EtKsF2CQgTgMIWatIkh2luTXOT1/P+FlAggPHcTw2bMKH09jKVRgfZ6
kvZLXmuDyuxoUagVv2YKkrgo51bplHsVzPfWR9yqZ+g9IXnSVEo/EYYS/ynJsRuKPW1+3npJ3AcP
DzPgbimW9RKiOIbAR6ot7cOLZhZ/PslTvBxbllv4/pYmnMCnci1BFiAHjMVqpNLza+aO7oXtwsXY
MIzS0nTHezlybVgnsyThySsTcwyA4xj8CCR3SD5+sVmGgFZXbmuBtQJdMaTqph6MsiT9Ei1yHTHj
3aWKSxFUQR3oukK7zB/zz8Mc2gclEURENytMBkGU0WP4MKRXEnbjsmmeC/t9X3l2LDxJo5upB3gC
Y7yZO70SYKuCMWddCvEHT749PWDzRA1KqqiaDy/ivoQRJkOUsmdYHoTQZbuaVKDmv0468Wjty3By
kHLHemAVwrhwlIIbS+fBSHNaaPirhLXKKG3x6s/xT3Dxy2A9naZJrzL67GsfozFS50F4TPwLGfPs
WMPq08Reu3u3buBO02YQBpF6muQLaolKxs+xGsIngCsM9akff2W7VJ75XMl9CtqSP8StLRZh5nr0
aK7UR6TtGuN66+ViTonBFzeOM6ojOuMe+H/3hamnxBcpUz/LPUyhJgJnQeyHv5gEr86SM96s6z1D
AzKjlsG6ybsecHQWPo0KAt09iYQfyW1+E/IdTW9zW3SGtCX5M9N+twVHMEIC/tCcVtNXNa5Cd9Aj
eq07yikUiVKwcDoValgk4z6ZsTtSqmFqOF0MqRxxOXLg4PGHF0z4Hr73Wm1NYly4C0ejiYPNijgX
c2D9+xTNFN8g68JJ0NkDsqIcETBdyLgPnJvQebiaT3eXE5E3UWKqVULYZU6dwMDcPOq35+2efRXc
gkqz86fr9aK2c1vMSHVXXX2ctLK3E95G5Wx0Oiaouy3yTheK/8GVTUqxi5UkGuj05woqpSx9qKTE
F3090MSq9DNrfQlTpA0sH1tfK3imozO8/7KgLKtfzA1MAKnLfQvASM3Du9KHoWJddZ42DGF6FjeD
xrSgO5pPnfvAKpUByx8mZUIUT8qtyOwK7TX+UyJtkwvzkdCRCis9mk7INdmyptk0JZrtm0lGPVYX
S0JANxErgtyUNeGetax5FkQ8iJaIL+CTeUo1DdvkMjlAUR1/0w8CJrHL27y2MDOHcm5ZTuGfmw2H
IVvfg+QJ/MzIL9u3K8aIMLwMk2416LkR3lZDwWe1SwXNKAZT1bJugR5ggR5Rb9VAClYVXnebT9Ui
2HbAn+XYxJOX66JJFjlGtVbN2djkdlC9ut3g+G7MnUtcVEQwe/kOt92hSumRJnHDxCbrnrYjouYO
7/2AKlqqp4NmUHAfbXebyUpmrJVBx8Dv0hBYNqT0KDhXnFovapCE464iTr+i5ecgpxjG+uVUk5u0
aSn6cEnolS8k5YkG78AutaRiiHyScfMt0gQQmNhUup2clN1gGZQkeW+EBy6igrgl3gUMg0tA88ld
q2WE53xNnwT+i74mD01GFJTdnl4xs8mVVkV2e0hT+C1MbLBSfFIagv1LmUII2pdeFqmpkr18Ug8+
9hPx2G90RbzsETXdor5XSJsuP3JyT66bLNML7dAuRDiZBojCjzcdBTHs7AgIWnRjuRGpCUwl/T4Q
l0SOupUPaDWw2ruSF3ialQvzg5gnL76jTJIIr3fBn90Cbaw+eKqC63GTJNFqnrF9hBCDa3pS4fYM
pTVgU2mx9Uh1lscHvg1LDrJKjH2JpXiw7fSCEmZJDJXKfnzL9Dpt838MkHtNj8PomQ7KHbw5QSub
1xkqyt1pwSp+c9obMdKUJrn93ptUTVO9AAF6uh6l8ZWSE9aUJ71I25nPNiNoA4UTK3ALEsJdTEVl
U1qZzQC0hnJMOJt8fHUOARwHk9hShPskfpBh8AkAAJYFr4X7h9/nDb92qOdikfwxKgYyRp4SeSp4
O/ZCSKJ2sBFWL7xkuUdbLwwu2ftA2ChlbaK+0hR/+j/dtu7BaOGOocbCG/q0UfvZdcC2DuLenH7H
afGgjQ3mzOx6Ypkl7Qu5KVpMUdw7g09V0FTwPq9wPVP/J/7Ff7tEWdPuEqXcfvk5dttnIic+AENf
LN3bKkA8nvfK5C+PwEc3YxhN9mh4QbWJqor4ZsdgbgYO8WEZq+Ycn0EQho8KVha+iJu4JPKK4LE3
Yt9zPqZ+qTiZuO/UdPTCcw7A+9Ccxw56BxmLEFpgSpwfLxDKTmmg4jgVAJ7n94rGOQDL2HDaA0uG
r+lxbD+cypUcDOuJPvpaRXMtTIYpvOx1eXcrhhZ9ugWZZLHeYRysnYPRea6m6TYTuP78DLJmQAWP
OXYa5I+BprLsRPuNvdbr2sa6IkYxLMOTGPlAgY2d6FhhrDvgnf1fr6LJLYWFb8gPCpPd3n6B9kiO
BQFDspbMBehJiLvl0hccFi+B6WkuccXjgE90FrLStmtFQhQ9iJRO4BRwdjw/Uzg62KCt5UcP47+8
RPNsky61fY6a23aTJiEHGoj31rRyOgK+i2tii6nfKrCfZakspTOddpkhot1459sSt10aNBcBvX04
tDtiMmwQZi8oIzjfSYkanisBvrvPctAVBgk5C6xMCNEb5zuDfbJ9Eb9gh/ghO29p3rVIJjaRGMWU
a4/+ztlzPPWekkKJ8QLGXvcnNFFOx0kQds4dQWw+j2REDrU22nUHsGyulI8zjdmemQKTMgyAC9jo
Ie2yZyIDVjWdLDVLVt9SBjHCIObGtSwOHk60MgofVes81RnuAL5WM+YNZ29TfddzUa4IGTqXlIKP
g6FGzHugaeDeo9BpMlQiayVG73ETftKlTa7wRY9jh4FGRugKzeRVMHsT7MroMJrhOW93VPmD+pyR
YacdDRQUuPBZqiRWxy91uKs8bjWy9dWmyMUUZb6yPHgQfaqBBtFDUBalDO3ZzASkSlBxXrpXelUT
2jL65fEocJgal27x2Zbqi+W/8KU4Sx3NP+6hNIRHRwd3+zHLtHr+IF5bZ8GOIH9rwG7J0G3gV1+D
ypPi1z8b37WZmb42QGyBOKeMFkmmjeR9RMFAvVYggNbj8beaEs/kwgUzX8ysP3uwjTDTTfgMoHke
GiTKiVTnefIQsO46QKTaXb36S2iGCkgWAeKKJ2Rs1DftrSLN9a9uOoOpSqyMcopAO9lVKBoovuPJ
6E+F9Q8HORlLyvp0EouyyFzllEycWUddxb+2ZhdQMc8yzkVO3H0qUTrDTomHK/gK/aHjYcpOeDig
mcnawWdshrOyBD4jnCNUiN/oS0uEoqev4mWWnNEMapbr5ig391wdQiaU18vwKjxZMon33e6CBp2c
pcP9epGWstu1r3ORxcJX2zX50QWLDVV2fT2RgU1094t4ro+IZbGtOFREo/M2nwq3b+SlYUAr+u34
HT6STQ+9lLzaWX5ruJAxquq2qOJubhgR4/V40N+U6QHEot8dLOz2A1vnAeMXduR7wtpfOijklegi
Wxh3VDOMqqBceEs6y93vU8l6XLZlCxrDYBmV1qL+6iUkzk4CG7EeZdnp3Md17rbldIylwvmiah+N
kq9rFU2NAp5AR2K+GAdux2KQqCBp7aU+RG98QtRC/iDp5yp94Q9ppZ2tbIobAZcCjN/qH1W7AMkF
QOglxxG944MI1YhjwAy3Ui0x4nu1USVMZ/jdLPDj9XA540vaNuRVIJCIjL+Z2CfUquAPRcgclPDk
Xci3FVqYYusfMPOCfyExhOTE4Zon6AToyz9gDZGaHyrbFjD0DSqtJFsgAlkif1syHFYuT1bKdkqg
nUerZX9pOwiebjZaC58QkRupw/X2ojXgbITEi0bHd2H1Ij0THAZGCDVxCYS77ZS4bS+L9QPaiKlE
WnV0QcXolIDIpgh1Pc+/i4UPJrPcPFd2ksAlhrdKv0MPG4Vq0LIiEgK/QOlHuMosAquH0eaUYpbB
uWCOUlIvgSTlHEF0EgcPCbp5wn1hOc0+YlUAvKH6GPTgH+UY0wXFBzYjj9O/O/bGTQfbQXFHRDPt
TGIIBi5nCQABtnBbT9/XioXEa/D7tzToIlIXzynLE+KPCQ4BflTIW6LNCMyFlOofaR8Ya09aSnBH
Tm+zSyesnYZbJI4zHuvLuRT6ZTvG7K0U2KepENU1pVnvRfaejqEDZt1FiR1c4S1IjmtLwYfoeU7+
5inGcIWThp4VXTeCx1CZadlKL3NkdTMA4/AekZjszkJPZrTnDGIGfIMb3qlbw0Vm5FNtoBs8/9/Q
Wip7DEF+ghqybsx7WicjJwRQf1Y5/vSylaaB0O/wyFKgkhq4Vr/Ukyy1TI2MIzEpRTZfZ3Ci7oWD
HJo+ocfHAf1rHDJdtamPiouf3HajClOIJ8cSEo0Az+MfiIJwZJTeg7b4XxUmR5XTXl+d/ugBjI/N
lVn6Me3pbWEAFf+pIita7bKDeQJQ14DK2dsov++IDfh7KV5NnQwuHdOlpw9r6zP8Yqn93/5vNOCo
RLw3pDvXB9RRmBC3suSWTy0BT5qtsNv08aySyU026B4jiQDvtfnHdJ07svHW03fmOVHomfYBbv8E
Z0sEKqyBfCfGoATjIzaaH+yMxiqK+fzdLdvwCmRRAPiiyp3gVRpe2MlZkZ5t/T4lgY+UL+cb8d2S
wRzrzTH7QnQ1OtC1PpybwaADGEqrcUWLJItKgNHft2Mv6pg3pKa+Kdtt2hKEPIN3j5NE8WiXC3dA
7Wu4xwaWoeoejXPWKzHypMUr6mifr8NdUhqDuy0jirG1e8E3PoGUiK36tM89hIM4H2kUU1dU4AP0
y3gRxFQ8PGGXHs3W+smfBn52tCnhn2AIoudcmFtcRQHplT9rKZqPNBZ9Lgnek7wV+AX6W8tOGfqP
5s2fPc8ux3URZzg4blc/vxLECU7RpHO1Vnk69MgaSLMD188Lf54yEP98Q/N4ksF/GWAapwzWC2L6
JxaOvLYGIICH/MfLHNM5K2Zm0jboP3HW6QP1kcmsJjYb8DqxM1EWH02z6Ka4Use0QRFbGREVJrVn
Nhpje60lJEeJVQ/fL3CrXUM8B6IzAzuC6/1gIISK3GfpyRc7PD9WhXethFc8cFp5AYmzUYhEZpG7
zs7i87g9cbktDDRO6fZ/mGDIXT1YtjAijXCIUq+3NE8fnWM3fAapJgwKrzgNkaKFR6kATVbk1gf4
Rrtc5kLbCVK+Xo20Qr/a+lrpm8N11d6mJs8C70OPMQxrLSd7e+YAGmy0b3tHygrVb7hudL7Taa9I
Khl5i8dtZXzPU35HT4xascm15IAea2mZhdNzd5tX66bHbH5sX+fpaVtDddw/1zknbqQxasi2a5kh
3xiFx1rzbwjn5fbQ/4EVt/SYn+q7CTeQ/LO3/OQLZVb1haF5bcWrbOeD5c5R83C93pjW+A3K/Qqi
NXa005V9qLUzDpNEquD7wc4J1eUJCEKU/IZsMfklcIiWPs7ww2KM6C3d7zpCa3NpbHMVB4DehIYj
b1O7z4rlMPt17iIAIuidrVhPRqHmLQ326zhcPzgrSLFa6x9PYXmD0AJR7si3rLsLXUfM7mQ3Va+0
jChKouBQUQnSpA/9ij6XF88dil3B3QJshBruyHAjEXctgY8KRiOyLEdg7rYz0UCiAEfzXWh2n2sF
MUWMgRVCWKwp6y7mB7uGpQq6CDCW5E/XzWCi+w1gkeL0sB8olLZRrrnPFgsxexlO52PMNa1owsID
53CrYnXkBymC7Jl8IB6co6zxNtIWQ4RnVXVbL7OQnwko074NeDkNtblOZq1wJkcvSieqeamvIqCO
sdugTOj0fIpXzFEh4TTUk12eTrX+CiQhVMWqHIuDLpSgEQsNHgoHxQCL6hHEk1lM8nXXKj06IA5R
DcM6Hfa7MtyAu/Zw0F82MW8JUNkGWtvWMnTk0s4R1G8BN377dNKmvrhsQ+bAEFwn8/WEzAqRNtoR
Kc4CDUldm2mF/Yzox68mk72AMZP2dCpNhKHgtL1qAWaOUZfDlXpYNpGU0L6XwBbxRVu9e0av3m4n
Vw9eqaYPDmDnjZjIGzsNxhFTAAxmdgDwatXAiPUN9xXaA7ltY+FDgxZVyI/lN970/JD/V5rvV6sd
g/d4xBsW+e1ZbfIngTth4v3nnsQJo5yqyFWNKOGYSbE9DjilhWdlkjaffvg6TjG0zD47aZVfqkh0
NNn/8rHYrCiO3yDArk2WGXfwcSsYc0G4YwFK+/AuyAObZIyguALXh0I8e2sLJSpFlQnKf5Zru4cO
TztQPdqXQFd7c3m3VHYOZJV71gSDiem9ExKU0TNgpkQmbCXfbUF9hZqRvy7cVktSl/8poRCrmf1p
6MfxYMk0T7r/pgJ7LcSkeV+yzs6ODEorAMwvY7w6zmyWqT0wR2NU3SSqrgZ/BE5kV5vejZX+GsSA
QYo6CkKUXH0JjUeffMkV/CEI73KxmhogWVqo2OGvk7zriODPkjLQXVdx/lD4BXzfM/t7SnTMNS81
EinsAPFP8rYgE8kRvt03Cb+nYcgwWOikXOVOi9X9gRthvahNcdKyv6tYOFcFs0pAZrxPsMWstHjd
Fsq7zIXjBuMzM9TdO31KuFMc15eESELMS/ZRxBGuOOmJMxLrbunHe3B4i1YsYawxmMGOc4astXMC
/spXMbLffSae36y8mJRbsxj+MnxYlQ7Hkg41CkFuYH4/WHuTAmCSjgXQT5nQZdhQkd+exp2UFyPQ
7rxziMJ8Cc2/yeLioQiwZF6JvGOUZzU9FiLwTqrz5qZIYXesSCi95f2sXsQ2ntw0eJbPpFwwbS6B
dYFkn7LkJ8Opo/zLb9XMa+c0KWHr8nHJ9ht2rVGmGewLniSNBtzyJoLsMKcElfM0Tlrfn0U7pR+U
G+E4hCxNufmICH/JUBAbXz8CNQ1f6mftpHzirz5wjaU+TMNTWoSg4PZMgOdX62/oyxmGPQJJDCFm
VS5pw9bttn/rJ2ug9MvWM4BKN5spU7gilcJLrmJo/0LUw20FDVnOJ9VxbEq6GkEPtOEYAHaoPCF3
MfvGgKHtGGBzQs0+Ffvd3jMBTiN3Y9E6GJQHwY83t4zqmTz5MjQwmYXKBAzavNP9vFOai8P/h2Ih
NHjfh7MHFpLW/f3j40kao3T/9qyhHz595x/TfHlMiK4Y9uiLNNLDiXb+6TJqvqMiWTm2tG7NJ9AP
ix+HXvtIXPHN6K9D735XIeYDsNDsZVrNZOKPK9irK885gpaZuQrS36oAr6wBjIjZS2hTEzw7v+sY
hoa/tAcDSdFvWcwpcIAGCVnedkS11EQr3azCszuLZ/sfDjgN/3+kii1q/YYruQyp0j6ejcApN+SN
SVLa2NZIJUS7XJeqwXYhsgOwVoQi7LxupuP+2Pr7DYmL1KJkM+DsykQlbcQuPrdB0rfrGsqTM40t
euZp3hpQO0IB88FYdnn6WMq6igKU0Hu/3h/oXYoTNBs0Ilk425FHj17hFSUKKI8s4UUcUov3AWdQ
sfuwz63dT1HEb8JnkCDSFzaV3AamFljy3W8OBRVpjk56aUnd9E0D4gI+VhYgoFrkSNZl6JJCYoXU
FPPKeLhaRZUmKgi3XommPKBuBGVNXzbs+cG3L4ohRF6sl9QmV+HxFPvSX6XhlN5As3eS3NQ92QiV
DZJ61mYJRuhQtymAXk27xc+5bhrxLeTmS71UXyIItcHuWAn7HLfYnk/8ZcFV339xDsYOR26EqFuc
dhSRGCpiho3tDNXwN1YHLH62cry/GCz3nNSIlhoHMzL36KwzGjXPYjqdEV+6jnOIscB9FmvZFpGZ
o5Kbp/ANgFVo8q1bwp+H7Jh0vZ+7EUaEE6VuOjVtaUEIXa2npgHh/ajFcyhlJUuuCeBGcrfD4iLK
EL4FC2Nroj/8+h8pVFHx1gQlnPLHbaD47MBs8a19tjmTAKBFPnYpC/k1BkEQifjIdGvTmdkDInue
z6WqRuIFT5WZylmSGmp44y6PW4nwk1x8PE9GJBO098t+8d5ROwLtrQT4NmrpS45wGQrcxfhtNCEv
NEEB/gXUBH3cXez4aaHNOddQLxEIldF11l4E5PLXS26UBVaHAcjClSshxAHG4e94xgP9YX9AwgkA
BZp/QKQN2ZgFBI4jQAa4l8HBEtUZRQXfrbcgguBMfCYoBS82i1t1ONjxfuRamduz8llY82eOQoTw
GKrs3wgwCWOMM9LQYMi3sVbFg45ws1ANYjE5cItvworq60uesNs37Vjbg2jzw9u3DlMMNs3Gxy5F
6+eh/rZ5PPocqAOa7F9eo3Mjh7qdSxuwMVAohhoL3+0K4bd88D56GEDpcEw8Q+v5+DxY6myrcC3u
/XSBhmW4XHG4xPomk1Bb55mcQLKR0QFhRbL7IAKzfejZdqrpWH6db13FeVPOCyY+K9lcBLuZB7oR
NB6w0phaKYlDMnGRfsrzPJkUhHbj4auU0KI5QSWYUpsHz2Qf4yDNIHSBGRsIrsTM/5ctDZx4t/o5
1wn6N6ToBtG6UnBQnzUvNL8m/jMSxbU+fSnoYskskRRap/KRqdYUo4XaDJa8bGcvxQKKlBTV9Wu4
kD2YkQ6Z3x894l8mtj9SPLZ3UtAFfPs+43TbG1UFUDZyfhuj0LCLF7akBADqxPcMhiDxFVMf8xfz
pIYfiWlPk5Z1MdTZ3BY29sT6CsBlXDGVlqn7Pihky0IwVjx0em8g0bV4y4YTuh3Q+y6LkfOQ9Zto
3UH1a+I0CoOjZ9cSue2TYW7rnu6aR2rL9+3ZNwfQQU/LOBcl9CeoQ3ysEvxy7t9CDNtif83f5cSB
3zJPg9YMEbkwSrHqIl3iR/rOGmwhDNk+G1BAgOkXmyEHxf76xQDeBbYkEaL9r+ifRjcWfPbME4p6
tiyolTZpY5K9LfooZf0/W72e0gKWyGGLX2kRSN03A4hymp41jGvdCb3Kg0+oaXK2V3ZeXT4xtLHy
/C+NZ1QqhjC1mjNs9iKtTwCRhD5Nq9zjVdAw2ev3sAgfllh6hUsKh2SJOPVlwe1WhyD8dMrXdNpx
59fCP7mvLQeF2K8oTXSKay2V4WdYuoGUbahnFD8THh9O01gBYsV+3koZwZ97x4sCPIRcAmEhyR5J
FoQsH9dFa9rm5NGPaSt7H4+MUQGa7AnoI8rgyqa3hk4KUuMNjSLycd82WdWXbE3gGC3pl2APSwip
PyRV0sF8XJqKYgSzKoutMOQPlSirLtThNAhULNJWAHin0uuc7bLrzt5UhZSxFpITPnZv5ru8ybge
tQrtZjhcszwsRaoSQVA73BZQYoy8EUbhKRE4gJiKg5T7PbmdN0Djp8aeSi/kcQB2Laz2wfMBZYuu
exs1NaiEkUItwtqLhrIOFs2pfDCr7zlpEXlm8z5HiIkyigwJcvifdkYeoKU3DZRkuX7/cpbra77t
2vt0TyQxrisA4s7YGt2oZ5SAe7Rp029wx8UGeOtAgL++8ZENSmd82npL1DJ1dPGrdtbs1kyJEVKJ
S68nXufZkIf8NhwXqN6IflQgg0FBWdJ7yOtTRw9AxwAAEEwjxeFPaDrELvFkGPH0U2qvXY80YQWS
Hd+6ffcf27G6fKe8qI6+pwvqx51yxZE6IT0KPhs1oMZLu4zvq/uANEwpn4mvpEb4eXq129g84BVC
hXdb/rm+2EkTafdHUaC/ZezITDGKV6bnAs6NvMKj6EcDg5id0mcqoK90io+Bx3bk7kYWntdM/Yag
pV8RxoCtYwxG+SrvNHWQZ3n75N5O8amGRzPxPQI1cyADMsxUNScMgVPCKJTElBvOmva+jqHah1hF
6Q0UhOOOwWx+raftRQrtCXaOrU/IwSKrtu7xiBT8IMrU4QVxLygGY9l3gVwQ4nJcJSYhexc/ARe1
H5hX9ntvUOwtIZBFEeRHF7aksGOaYoXd2c+APcQ5zO4g9ITyz8vRjSVdpdMTpl6LnLD0QSo27yNo
EW2u/qdsLR1+cc7LhHG1evgUXGblCy7ZlH4953RbLHFirmEm1YR2keETSJUVCs6IPpogvbSJBDfj
EKr86V1tMalWVw24isleCIJJgT2flq1XeTrqT3t58lTEDYE1OKqKq5G5tQcCUN4tfWRev6c01C2W
ztwi/Rx3W/hkSouhCb/VeEAdLA7VkiQwZNoZcdFswVviBEPCNNaz+4Lz30ADbEGqSpJ8vfxYH1gP
SGJl965Hn34g1sWSdrs/SI09tMAB04TKVDLPTc4Zj/mBL96RuwQx1yvkP/OlY6S33wCDUaeCfbDK
bR7nQe+EEFWPUpOiO/1rCoGX7vtWa78VBb1Vy+DjpalsepZHjFjhO34JDCSyaEUgkx9iXh3Jl5FW
kk+t+plkIDd/KU4gdUrn5nbWRG0Ce5XQZH3kBLJmlgFvPX1ncIBFUDA3AaOEpTwxYKxN5jX+Ceij
E/iYCn8CCGFd2StbVAM1c6iVXk87cWe7eo5O3GT60EwNFlE2zfzjuXDo1NlGaQfDIO0NvRnQj+FK
37LMhX9CFl9NHszDrkbUqkeQ/bF0ApQP3BsWFITo04XnhI0AxG4ZpGtY9ERtWrL99Y1korUAdxZM
NqqvzKeU0/z5zFg+vlZILfxVMD5jqVXPPNogWctUXmiUiO7U08LDqZ4xBedrhQ8PlA3UY3jqzvR+
asjAa7LD19iKMG0uH1mOWJKr2IvuJuWSBRHRbqFHAVGZGPMuOZx6k2um0vPGBhsX/gozyNPzkhpw
meNz2FgQZYL4oZqKmLOZq68ugbDsofmxSfidaFyi0awDR/46s7wO8QYQ1CXMmrj5QcwRYzsyzku0
JNuS0u3heIDsOcTaCvYzTU9EFbyx5AMLBYPk3DQRjQNWo2Zk5sCX6w93Rvav7ChCpqcNZXDUXlKY
2nZ+GS5iIqjXQ44wnTltj29C3hEuH5elkZnpEbCRqtoJlqJ4DAZ+Oa6DQSffDIKZB68plZH/ERgU
vShyUB+PjZiju/6MKtcUZvOoyRKmjoZ9ShzMzilLSwG6LRxSa3zF+SevIc+eAa3Q3h5/kDd1Rz8w
c0iintQ5Aq+YF19YFPUvyQzycvlyuioc/B4WMTj549NU5/j1xP+HZS83vSVXLLy+/SaFMGi8aD/f
hD31R/RBO/NmKZdpenhC8FYefYXNijWTerdgMSo2K5sK2VT8m7HHSlSBkUvuajzDkC9uAhIybZIp
EBXpgYjk5NgmaGVGYqi89J9/BAreJzBahQzkxlPhEoTcEnzfmURsnNalA0f8XpxH9ub97ItG+yXn
neBNHFQGZYHnr0fj2K3QejJRp1i7MMa+SV9dtlTgJ8gJStRLnAqNngCehDHMq2LM0ETdDtajpvlR
PmGQdOCfRmiO+fLGsluRtMc0q3x+HzFR34dVew8g4ERIEn6xN6OdPVAn9+OKIMNMK92GTSuT6xaQ
Q2Uo183jhtiJg1jcXzWigEcxUKwgOnwK4qw8QwTWyXMp23pjWDK7ElNek3NMDD2Sy8EFXhGyFDov
dWuVDOGibxF95Tfuuzu+4L5Dr+k7nAzoJA/uBrxz8nGv/MlDKWb+IjL8gG6WAeumoa5Cam5kT7yH
wCXsCXsIcYsOohdCL3553GYWfGwhhhNF10651Z+7+S+MIaqFTs/rfaMDv9naUpK6JMdMT/+HSzsz
MqqH1u7bL+sUrajAd/O9Fbw/AX04qEY/j6Pa7sW1reMmftfHVNbmlmZPenFatL/NHKC3pLnrFyDA
EqLYS5O0f+BzWCsBO0YHEmrsVzPy9w6H9OX7aMTnWTxvnElNEfv263fmJsoR1YB+iw1SICF7FWeM
ct1C4YNCRWJLUIIoacYJhfq5rjOkGXcZOZOsQbIMhY6Mo8O1QzqipM1sJUDHaZoAqfq6EkVa2vjt
PrMsjmN4/jKE/5mFgk0hwhTN+RlboHnGlbZ9UJ986OjtUI4Dqn+s6Ee7la1EpKeOs2SVxYNWV949
SlPUoFOps0xjQbo6eqJymUXlv1+/j23JOEDQqPbu2ZBYGc3gkxptTdvup15QoVuSMp2AqO4hlOc6
pP4FL1MLnEsgWlDl/bJ2CbKpF6MfBDjtAaNnauora21qcEsUEGBf7i9DxkV4uzrrlWtLQtRzKr93
WGwoeeRFhwxSfRbM+THy9RPIJ6yJsPwViX+wZ1Qcelozy/7SWra/hly/d9ouPEsVVMyySX78fvIc
Y/qWxRNZU05cwZVYGQSliN7z8Vq9kywqdCKOhbDNjT6GhiBRTI7m2aKD6ww4+GD4arddFTcdFiFh
/XbJLQBCOiG6c/A/SG1P4p6KGcgb4thhl4UiLzxRQSW9/lsEZ+ySyyxwV2UXbO9DCmLqub2TH0FG
unPESGuhfXHWXBWqCeHo4zPPhQJ/AqsKf411MJ8iBEqIYUmeWD6wrdbf8qxIx2sEVqfJbVFzltBH
vdZODd+JxAK8GsZ4SSMdQG3287S9E2USVoa+JeL1U73OJSwny8hLJppA54V7SVZTzozZVQav/nVh
HWc9gVjmfr9kRBOWTUoyMH8d+s/M8E7B05k4tnRvEp5jn069V6pMYgNV9+kKCc1RsPZcjcYBbovt
pzCEGIQStXFk+6c1IL+8o0VcciyIf1BiDXV8diRstBYlO2cn9385AL0nakuo6YUOMuW2U8ftkf6Y
DtKL/lX3ENgy+iamfmCy8r8mN0x2DGUz8bEiv1MJovuQjcuNfLcnh1Pfykh67XM71N/TN93YHJ2l
MNLQqXbFgnK1OetvLwPR1IboNJa6NO9B0TOOuZ+eGK7A+kvHE6WYxQmVHbRxFuKMvlVZOkpgePdj
2AI1A0bdx4iNyX3C148LDXXD/phSM1D5OxSUU8rWulyc1krUNF/zRof5esl3oG7YW4ePUI6rGjIS
iB4poOq9jmSiv8vtJYHieQ9IwORagGEg4y8JvBUfTlUbIgjaesVpcB1E/Z8p45uXhAF+fc/sna9v
5ExdAiTRRENQKDVbgg3bDvC0B32IS8P/TW0wTv1FC+07S6kZHwhpaK08oQK94r8DBaLs0BLtp5Iz
UpMyrWa7PjthS44sfFJ0lz5fn3ppVsBA9skmHWDqv7LhorRP5Egm5sCn9qXqKb10wd+mc1JeWk9o
Na0W3OH/dJQfssi2pQRneULlPbZrgG6703SI+r/LfaOUdgLUE58Zo/NalxjK88nb0EWCc1q1xBQD
c3u9zaE/FOfmEuTaZYkfou7DMOr007urnyva8yxNZcBEwk9lK0j//qaHNyhOhfqGl+9UFsg372NV
unZcAuANWpejObe3fqx0vLTriOlxz/EpRM7DaZbIgT3oihPzzEaVsQ0y77dTbVWc7wchTWML5BmO
pJCba62jlNn6Y1tgao5iRz4oCiV6DRoe0JsEeZRZvq1cgcnuvDJJ/PGPHnXYwWEp6OmgY9HJr0Hp
tQgqEjMP/+ioorvdjO59PpjuXHuKhDlJNERPqmhkRMudNG9Pb3cr6Rz+qgOs+9ZBmKiljE0wQztM
Mv7ZBoYbP2m8KrBvyh7qwykek7/ARd5sAmVwvwm2xQmK5QyGzpZF6mhjAs9eAmMC8fXDjfGi2Gwd
iST+AfQx6owQGNoYV/7xHakzlsEgWYzIzFXzbV6R5ljwZrWHWtT58OkyJpyGfIraZotfqPM0Rgby
jxcbuiWgwL2nQ7oFmJ8U7B6b/687ii7S1+OvNZTy8X2girGp1HIxq3wnT0gaQi3MQ/WacLLEGaDl
DPkrI6jK70lI3n48jvSrrBfeb0XeYnNVdJjdxQz2+9rqCQyEvk2Munp5wTZZRTJFIYtXYDt1JIKh
8aeVBcsab7sD3SVnyDJvXBbFlickslh9j8A4U5ekWkm//gdrf/E4axsw/BXF0PPdCjb/TclC1caV
4jr3x1lAmEK8MuED0KVfd8c7whefd0fuDsrVs+0LAUqi4WWlpZvHZMIj6cmEEMPMEotoeZL+ZiTk
lzeWvajYdVkw54OyA/lQnz2HkRx+amCUBQVhIujue2bkv3Rr5DR1PpRer6v3occPNY8W7MlFHKvu
Pn3MW3iNORvuvPzlxqMWAB5zTkn4OQf/a4YMs3uucCD/An5/HMwjsPCJz2MGxZKVd1wBvERrLAvC
HYdMZte25OHpojPgKlD1+13ZM04wXCV6u9fRAwAUU8YKu3sDYvtz42pUKJ02Jfz8UQnQFuZZ6gNd
bUVRrBJUgroKYTXeEFRik0MVYqW2CwvOpgpvT7d7V4L6i/TXLJmZSrC9BiLGijgPR1Uy+7oM9Tm3
GFpIJ8CknGe9P2JprWXqwJngfceSOCZlBJXX7SpwiXPrCg/UUq/cOnouum2+PRSZSXLtrzTdJTKW
b7c1FXpfzKP8PhfWF6ytD5tIu5b7/o4Qf+BwS1eHhKmVJOC7ZIIJP6Y0S/9r9WQyUMHmabCzqykD
xTgOvm8dABLCWqviHGouQoE4EUw5oOxn6TEPqRZZU3o1kf8652Zz/kWGr+RT/5POQ34z0ALBbrdT
H217BvlKO+WGz0LzgC+c7Gt5E4rwptk2fjV3YXmgiZFsD4iNHiTXbbEtXD0658Oh0bNbghn0XaLe
xoe6v+kD3XLnKp35EsZZ15XsYgg5bLANjmeZu8n7bmRlAV1tlWon8B2yTgdMmihYDl78uZVQhBYe
z3dmZXg00RTyNQCAWSZ3WQFPgPuZeGL1boHZ2e2mBQMxsi1FgyDVhbhX6z92hSJAXiOA07aCALRS
JRbArc3VWJRufge9fiIYVTIH1V1yGmUkGWtY9E5QLUHkCF10BzI3/r798b0GCTM8ML6eCcZ0SnMM
IrLsRKYRvFUhTUqteh6PeWQAA3BEVrfanJclXG5J8rP+rrKvOJxr8D4ZH9ReMi6QN4409wBy4eTs
nTQQ7UlBC7uFcmg0izcPqK8gD6vmChSjie4YpVKmHykgawW8iNt4onRL3sdkDLpgoYyzZ4T0Ei9O
pw+wyy3hs2p9bfDBm1c/Wxur8SEaFyQd56XMAY52K89T8qiIJZM8s71dOQIA1/Q2fpAEfx+GQfUx
VR4FLM2JaqK8DXllveUcHXA56kaCo2dDNilgc2cUjuKfjkIjFoubPept39iw9NpgHVx+5tagFKlt
jK5OW8U5TY+VxOBzbSXal+8+bdoAwreRUAK9ETnxKQ30+i359gDxIO3NO4AtYy5OhveQ5H1pUbLl
3ISSWRc++EBVxP1IURzpoqQQQbpZ+fVHOkNjaQ28xX8pFLbKNefv8ygMkX4qrql4frIY0l6EyQ6K
1OWUgsqfN/Qy8YHeaNRwquSamFReI+/Va05Pm08Ad8N0HRU2QP2oWIWVhW66zBCTDV0ANHFh8EsE
K4ytUNLdNEU3NNgWOtx/6seVQAhDrE/q2mqFK1X/M7PfEZmVKgsXSCgMXxD4aC4KaNE98eDOQ1w7
HPocOlAFhy+qVI5qQhnUene7sFhqZyOB3qdcliKcCeEEy2L3cZwYzzWMNbmdVlcJed4UeIdcZnsI
7uEEjR5OR11xAiJ4lB9pR5Q2eSGutivi1dfxCWtqvhRX4O1tNWWshpYexg0XCdceJW9uvdybQFu8
98fpG+9xqfDSA16F3DgqVOgTP4eCruIONT+w+PVSdnQmzpzJzo0GUQeYBoWiz0iLb/Uzm6LOZw/j
sZg1DoPXmCVfYVVgWWt3KROuuxWfI+GnEG1TXEgs2oB5hrhJ40LGFy9BWKgUayZFh/96LbW1u4At
n3WmeEC7qQ7tlxNkrhfRdaTYT9JLTSdbZitT3wDeCUI6d9TEPysUoMOGox0oPH2BKDT5q9Ocla5B
cBBuntQvb0iDl5HS/QHmXN31A+dv+8rVxFtAqdDARoandPF0ba1JLjLTsRz90nrzFTH7ylxjURlf
rO6x3NM+dNl5389Bf0Gb1souWmd4Sr2SoPAay5+sMnISdv/A+OQo4qbhtoms3dZGPmiCKj+8AwxC
B8g0LwawnOK1uwNTmWsAnpkc8ZaVJA/Hc0/vQKYo9tk2fhhwokXqPXU+oQCparIHeWkySK7efGWm
5BoNadQ+TYjJpjt4YtOXQV0RlHQTfVOoEWqMbx8TT+PiOCZ8BdNDpJzgi12440ojbzP4uUF1+z8H
nVS24F8YNJ/V83ASUsVFQZdPx6DMoVME7qyc2iCNyYJEiVGFvHcf7PxVBy2XLaEbvbfSfzT4IeUL
Kf6uDU8iNx7vuBBNXNsZT99JEOwce/ABmDnZLjl1E00rLw5nVub8peuWAoo4um+kh2phKS2n80df
imrMQ8+Ad1qyqGbuBrrsAWNf4LNzeQyvU8pT9c3JpdE7S9PPYUl5GYzWwJeiuDuKtNC1QlKaPP6P
/nY65aHn5ebLU0FI+Q7A5AdxJI7MirCwZo6Yh6Et/QV37mMAOhEA2Id1SCdJQI1uLC+/wqsL7MtI
ywkriyD25CqQDrmMPYTD6N2U1TyABNh9ua/C+jgOYzGO8ywj2fK2lBNBMRjFrmJBmvwmd08PKzWI
mc1BcJG/7R8lVF+jYGnEhfmohcGvnwvWUHW6yH4z0Ie4sTxR63gy6kRugd6qSgz+h6l8B/ko7uwr
0jgkCq+QyFkF+PL9y7Ne2b2iWSXbmGlftgy1bkDGp+bbLuWRJWe9/NAiVmOvzMV4iN3PfNjvqUVO
AWWG2LjHqkegjCibNnip4H/d3QcD9CqhR3atdF9xoYGes+vmm1hOZ29Pl/I3EoMeWZ1Ru54HYDCM
DLPQ/W55tlaPUckDRQceYZwsHo2hLITG0W+iCfs7karPWQJvKW2B1TPdRi0fV0R5ZdTYjAJHZ+vd
MuPEwFRSGNB13YfN16mnKdoGBqYfuFNVjvkb50wE1lOdqgGVSpvfqQgWmiWG+GuIPTGvRovdso6g
EltUE7hfTnlm4vfPn2tcU2o/iBviP5faUUsqgPvxZZAEAD07HNqFfin2PHEhrloHNZqOil4JPNWn
EQfkNX0n/6wTsJH8DM3ku51qUWm+uszLUcQh/Uxs4Q8z/xlDvhbKqyfQyRJxDzqK6acfuiGMYgQo
CsXSP4SP9BceURNAX/ARq1w5kTzQ2wHpP52Owvw3ZWlYZK7O3DrAx1XqYHGIMZQvQXU7ekxdR2Il
OKolAt4r9jc8MyjgxRnJAPtWnC42yZ+7fwI+vfkovyOhSQ2cslxlOVwaJiHg1T1qSMJBlloSJN8K
tdoBOxaqIo70Dgvu2juefhgvToAIhv5dgR/45WjDChHE3nghR+dUR5ZTgjxjASbJSzfNI7v16IBO
ntwuNunm1wQCK3D0FKqf6TxCgU1rJDKSVzrfsG+QYYeTFlud3osQUcdS88D53FIWSFEnhSHyMq2v
tcdDHQg2dJtX7GeQQn5cjW9WOEu2KNNprqYDnyMTZ91Tk5MZKmamu8yXjG99WyCRuOBsfSSpgZaS
zhrqwB9abC8yHikQyVFD7NaTIfaY1CJ5Zo9/ef17AEiYkPg5z/Ayr2OWw7EWeEueW/86AEkwutXA
GtXuw9eqWUmy7cPrTsxZ9j4cQ6FdPlXPNHgtB8O9h7bjA1yNsqbAom0EZjddEr5EGqDM+sfA3oht
M8LmhdwM8USmokIJrYnGqj82wbz2G2e/+am0hTMXyMwRYUT/kF8HHls5zuYK1ymWJda8p9zh5yzx
r0l6NtN+ORDc9iV4H7lB/rluTU+YF73pDtt8xl+zGWwF2OuF9VxeCEO27MURetDTrafPEnL/IKcu
CguxsZ4lFJuvsgmj6meEelWoMIziBG0c0W+7/NXJJbrq6K/csH1JVjfUUIzVQCPWLhRZLd2+EUhk
fpAxvCQCLJc9ICJd33VPu7lQxbVXxlJSmrztA23m/mzUlduGJbhtawsPefkqHoamO3sSfxguZjWv
RfuXN3CaYcoNAPJ+YrJOKfoey1nCOnk72xJxqAbPBdZzKos1XDcA+6ZuzIQ0HqjtSwNP1BesTZHN
xE6Zpnn7Iob2VWqj1ajGQ9c+RBzcoLenZ2Y95MzTci+rVzDE0TLXEFXNL2NKHosYJZrWs9wPH60n
8Whz559/Uuw4NrdHbyKRIW8tgCaW0iyJf1qMtfoO4y1IurUAiqEWLP5eVTwjZk8lkiiW71SZElVy
rBR6ll+hXNRH1i0Txqv4mFgq6kgJVRlAslafzHJ3sCoNFz0fOKO96avIT8Offan7jrh96rcB8fc8
ziBDKXGYFrr9705o5dXw6EsUbcPWhGmGiCiGro/sn5KDpM2voiW/3PXKSPDXDPM1XRtGXK0mHjZu
J2j3mW2fqBewpuRx1tEJExcST+7/Vb50vwMNVskcoV8oIP2PyiY251OQwvs5YVZ+x3xEfV3z5NJL
bIwPxGGhQabBX1QCbllDYdFmukuShod4ml4W4SmO7pvBRo3a+QZuvJpIRKJsGQFliHnNb3+K9igg
8l6/kGgAxeUoYIZikaUrLtXyFgxyuDOL1ynib/Qqq0+JW+pV5kXR/A5vgJVawp36gUATKfl/ouQO
zdsgqnsdSguxbHIYp41pZFpFZYYlK146y1Ddwfuom7lVySF0TPxwPzW4s1+MH+64no6mV4PholMa
vau4uIzCrzRDhmS09GWzSeMQK9Nt498ZVEJUkVtkkPaQ3uDEMgJBNJPOx3Ih0jwcv5uuomVU1Xj4
YE1HcXROBTMBrxEUkeiKFxq5aDPAlCiBtPrQ/AYy4tF2kHSk9FqZJcz2rrlpaOoWwYLO1v9LrF32
QpaEBVpvarISu5GT4bYHTNAvjrpLm41BITt27P69nzg4/KC8FCkeupooD5YEWHzdAL+FBjiyhTHF
Obj/wlwVhkN2UPEYKfrajSbsGkXn7pW5Fz0pohMt4QPcxu1r4ce10Sx8SwQ72vUZOEMdUM0ncKnL
yUQ2ZWV7iB/kHChWhtRAErseHB27D/kX1ANFxVK5VtE+9dWfRSei2i8SaWddEtRNmYE25dFuJ9GL
z/4wJ1D6XnodUVYgeP0YdPRzkg9YC1Ky6ZP4hdQOjP2kO27JoYpBVKAW0NiVx2THc3e9M5M0Seqn
HhNWCEmQG0jmw34G2nTS6nEg3z9XG7fzSYGS4RDkG+kw6Nabh+cPIdDS6rT9EK3MATMM6A/rBzyg
tHJ+Fez0LiB+BEU1LeblJx7+6lgw5dOE51u1iI2wqiTGjMIB16xcLxMBgPdBlgKygBC35JVPfTbX
LPZZgmN1u+x4d8z4j6UfpJGT3GxtUSoIGMJ5LPkKsyNLi0rNoEe8TP1RQyyNvxp/HfxWjeqnj1kM
h5pJ9DDntr3eUNLPOocfatnbG4ujLxe//jVm1P2G1CCI1NpZbC6lOd3ebEPsSWhPHmosVeZDQR9i
BwHnME08w+z1/vRJRZcsYOAN+/hbqOykpl6U3MZmyajgl/I7ES7ZjJ9lCslYGH/eWgQv+qhn5QPX
HbshcWOjv1nrI7XGY/JH8qdVDAPhbG5c/1gKC8iF3/wXzZul9ecDkjYW6JjTU9lFfLUqsvMKvAxC
Lrnj8qKVmZO85Hforc7k+MrhyOIXW6fuui2/xlp9NpUW6V2gaFunhI7/eQYDSd5DWzRefG+on6xD
wVTbcERvvMeLRZElSfjbs7qe/HaeiU2kTpC+lYJkzgX64KpD4g2CoQJ9/CKCvwXm19arWQKAhMjZ
Zgq4pqCeN61JkVewG8jCuc820pi8hqw6VObz9vQXlDlbFi1WcdUYWoEYKvIX8clXk1y0l01nJ3pE
5HM5RejNlqxXJBes9pGSgGBvhsrBXhmOkyLKoB6BkJ9jNcRgEj3UkwEEao9LiFC0v/jGlFXPZ9XS
5JXAW6mupEHJFqCX4BNvfaR49l+4J7ls+5DOBujc/QGFCrWbVO+DK34AaNf4Tso9X+i/76ulSrU6
MBo+ysbu/hPxocEha+sg9zba6Dets4OyfB4M7qTrCat/4z/t6Aq9EccPWBLhiPFGEPRP9oB1epbm
CryBfjSQ1GmNt8JiEEWGBj0cxwOFYxfXpbeUrgHOv7f4Csv+YCqeAzoZoQk+EV8IlAgTR3kUwwMa
St7lLFNjmZOtag8/3U2n2+sOmkoMMNai3c9uXYhhxofxLWCweX1YbvNwPAD4kOIA6nmtKh8j5cTX
GH4NYgY+gYtVd9f/rBCOoka6EBAz7P6Z9enp1hTcS9CNCir2g81GMorrwUGdNfWM/jYIKxwgyNY6
ESXhHsiY2wvxnJ9bEoIGNwhtBVBA/uOb5ZjsgBkVXvnznEMXvfi8mQTOpXZmYn++lxthivMUm/qF
PG34SDLndP1vH1SgV2EimHzBhkBJn3ZmmCqVcPVUuhDK3zSRBwiz7J9Gz2FQtkDU3PzZWRD8u0wf
uVEC4oPQGcbLsb+GwguYbERo2JQ0crxk34XBdeP2EljjoL/tiaIXqDKHW28BMTLqxkGmBepetfNj
xXWdFNdiKwuUgCxXExFS4x+HdEk9kcljBVLHmyaCJ8GnRCAlNyVXx8N38L0Zy0/AqSlsnpShiXXR
VhiLdoDuy8zozICZPSEc+LjURgRAGqyCkgscexCTh3gPXw8OBFIaxdAK/HqOZGQfEI4XxS1oHCfD
gtNTLcTEsAfcdCW4y3xNYdrJLm2Az7FZUR8fP5X+o5kRynwIjK9GCSKK+i/cYMC9QEAy7aQ5KAyP
fqArJ7gDdWgyYd/2YU7VDydCcNxBVaKSpACKQbKMTrrdX1tMUHjg0L+1/1xJzUPjalYYKjk75Ck7
e3nY6TTZCsDFp0cs2DV9RKxnkMKiHlMdloLHpC7Day3jGy5ywLtsSzobFyB6MlVpO8+DZNYX3WlS
3C+8oRUc8EgeFtfZ3kVGqA8FTUnHEMs8xVE0FTrA+WUn3WGA0EH42hzrr9JR1NbU2UNmIDHPsXtY
92fyTTTQcIiSq1/64pZHuXj6/vPYqjqs3jQv9TardmG+ZK09KNzQjHMwrB0YVmYA3B78kYbSCivv
r+Sj1Pn2apk+vGFPeAsSj/OR422nLxc8xKoiuIbdaoqoL2UVIA5a2BiIPHVsqQ6bQvO9X8UWh97j
k/u/8MBva2n2phbiLWctf/dqMmIYiCas5a/9RFjQNPnO0R1DuWy3z5K7TBc58TFmcs9+yFiij/MH
DI+ieqoa9We+t1pCjLgRfLVYPPPRUAdNKKVQH403ISC1ZMQYbLxmocmwQgFKyUnh04CewiXIFG4c
q2b81QzMvDbttrBe1GIHNL/4uiedCcXMTH9SNMQaW/gO8WhmWgTrTt0qSfPjGmMAqYeO+NNvTopt
MQgOdUhC/DAJalCTjxEie44HfvkexC2DmBBmaag9b0lWxT5eAKBL90DM8XpsV9VOFKuuaStk4ZQa
nDoGeLup3BR6qpgmE/DNgUMwr5QhK2rB91WWqaIsNpr15XxuFwZ+IznOEvPIsPUhhGeOYpQfN9tD
8lrm0nSComkbbPBibBdjOpdy9/EMJBaP2j7HIq5HTdtI+2Pja93M6EJszhIvgwJXvVwErP5LcVFC
uyp6E7KRVD+L0qpnVYVcFXAYfxf6sSnvGL7GBqjlOamIXx+Rges4tRbNuneOFpTBSCagfYJA3LtV
jxk2M0dILmcfgIH+sJNpzUMJWgilq8F/IUHB3Y3Q5CyjFkXEbms3RYBOV7sGiVizEgVGU+SqaQ5L
B8W+/2t4YCObavdci227oRBw4MqNFJzEc0SN1CqaV3U8NFNiwHYdYW0Ld9wL5BQzVMTlLrHyBHBT
4lyWDYEJkcj0VSDcb3GCU3CZ2nE+PSb4YEUTwMu3NCpKgAGSX0szM3Wryz9u8EcUMygfcVJoulE7
5SRDcZdxD9bVgYS3NPOJ7jjb7HJMrTiCU7q5Q0MZbQxxaI0z3LQM3pr0uJkcEOFco9ZFpFdvkcSJ
5ephUqHtSaGHvWWvAaD0XcZRF9Rq3GFNvpZXE8D4De8TaCvaHBsDA6FTqf3thFKhGbqax394Bn4L
CDkqqNBte8iHtJp8rqOgEPO7Cm8srGf0grEuEk7KEfATnw3K3m5x0n/c7vbkxrt/2CBwyp3b4H4y
R8zCgDvWO4KCt/A5y09HZpxS1wDwoNvBOuyTn0F6yxS6c80Ej/iXLSvNpvL53qpo4xg59qzQQdI4
SCFa9nhjim5R/GcTmV7RbBw6dc7AHzkEG3SJiLz+jZmFZvL6e4XbwOiGC5VCGJYCylwIBUUVFU1C
+nM4joB4EPy1Wc+E7qv9Oxy51SVkKdnK8EjILgSV4dPWZxu/kpHN4E3apkiPcFCeZJVefaWVbAuQ
RfzA25C9VS9WYCCYeFdBp7tJlfGQhxbGL+joIvXXKIWD+aNcOX5hgqYl60hLx3Q+wQtFg5X7q5ab
gNvp49nbX0euQeEz3Q7TW7E6Pi05cUk+ZJQ7BDDGmRjpRAKE4a210v5zUi/CR+w60RJSQ36dT1NV
GsrWjNm7w6RDLqsvz8bb4WbNvFSukNos+5ep76F4/TKU+LCXR/NfCBnDk5Hi0bMn8Lql6PD6w2rV
uGrjoqXe6XCkaJ0jfGiNOMP4BitVmBaHr51DmaNlD/HL97FoylFotyrNKipZqvuy5KfPxGV9kpmj
fw0WlJoWyCTQRujsZfW9uK93hCOIiZT1aFS48sV6R6L4xjQtG25S0680VltYbqdz/LiXMpK9BvkU
mWV6bUZxjWGGqkhYXrRaH1mwnunSK5CYef8IWUupqDpO8eVqqjk3o94zZI56eCYfBrDO8VsYUFZq
Y6qXolEXdb6GmhoYcMly+vtdiMi0NfKmF7yiocDXygz9/Sep8qnkGpxb3MFO8Z67I9bKcVaj35nc
ljVb5DPcbXyRZv2teahp0g5j58dhFW6wTffylLrfc9oUNbN2i86I66k/EuaPsUm77ll8w3Az+0WH
0OyUoNd9kHLEEGvZRMlLYg59TvYTryo4ER+yIRrwL72giS2dHMp7DxmC/FI8n+vyU5cfFN1uR5xs
7JEqSl0XgoWtJnX/tsQn6j1nxxVBAqaUCbkKG/+TwBX1stHmtGSorZmf5jWZXynJYxGYwaIWsBIW
dUDfisWjGZDyXL+KLyEvOEyDQcQmWOMf5mKjAbUMLLau12Dgrg+4xjDmaOLZN4OUIgoaL/XPpfIP
yCcPimc3/+8MNY53grW6f05AilJgLTuBzGGPRLcQF4x/NAOBynpmgamtdHbkL1t/qYB5akq7oftz
z/tRwrVOCKFBYO8coz11dbhcB+nZoIX3924fREaZVXhfFpP9Nvn0V4G9tJy3k7YCOfTFInmczEPN
lcpaGu4/d1xlI6iAbIpn3ZFFpV2ixYl1jZ5dj6DBqvw1QjPnKHk8ip9PxGZFGWY1uBzcDqFXimZU
dxDnIYAdnLcR7zOZ6fbAjS6vVxYEOe5V0Hxwag1PQKIbov99obw0yF57VtYc0ZiVG6o2TOJikb+E
zP711d7mj9TyS25UqaTJGtovBZ+U+IJ8gPc/klnsmPC/A9wRtkxfGEGz80WmAupoRZVcP/kJgSqa
eMc79EZh3EXudSouslLQdWJAoWjGSYY/t4Eb/ZSUY8jc4lVK/aZ7kpPoklA04qBOMiCVtZIDJzPm
iBAg+JJmy1HPvZv+MTWCI9BqAx6k543B3oJHmCD9xb733cEeeFn6yNQbp5eN1tX52BQKV7S00Mvg
ML/JqSYiglUH/BKMkeZmeKMnmcibpoGyoQ4oUiA3qeGjw6oMmoqMpF9vP4q/COTE99qmdIIqs+1A
u2rz+lDY8pSA4sQTRhSd+ZYynI1E9O2vkVRWDk1/suawuG/+RVR0WwbDwVNvT5n1Pq4WnKk3+3oQ
euWvoXVVQh2WVSIgbm53IjotGssqE+8vXQsCArkVHgfFyZlKbJtaLkYBjRk4IFOUYWekS5xAaPha
uZSOalUEnONZUxhwaLfbAv9BkegS4RRn7+PqPpRWCIo6lGh4ds/mce4ueMtiIsoTLMUDWEDyjF6C
sapLuha3fQgvab346H6jeYZXZ1Rf7VqIY3GYXNCUc6iIJUFpJf4xhna/erY/cX+B83XNeFOgkTrh
vTLTuSJqLUjLrySB6UuPzMk1MLDv1jRbDvrul9JptqracGCSrdjYkJS2H4FVIr+xrQtRxO9N6Jka
6SfIUU6SQT3YoFtsXxh0nKbT+hkoELA2Cv6XO7E14Udk61wN95/iUafSaWxzRpYLbBUDkonVKVff
P7f7CZfHDkPmTwS34vRhD1iaMF3dkxEHFWiKcd+2VLdjX8DUvks191Ph6Nr2WaZmnLZope5IuyWR
//DRB7QZnHRfq0sQYZdUOw45QxwOvjNMq4vpWC9yPnnkPgkG1Afv4CklnZxfGE/mEaFjmlQqHjjF
A5yUAjFGtVsKUhS1RV34MUh0N1p4leAWGNK4XrXTz1EeCbrOx6wS+wbhRk+KXZMMnD7EFNNCpTRo
h5hP12kkkiOO063VCIuZxiw2N9cgxXLwondlbfDEGVRHS9A8wuYAQeFf0tX1wt4AaOajJ65Mn80Q
Z85qbLQfuFsK6vG7Xf2TZQbtXmvO4V9Bi/KtGgAB0uwsNa4llAh44qF0Xs3h+G6rjj1SzzlwIYy/
LvWZaVuzMAhPtpLzQd3emjNvdHCyihTQIf6oKxaGQtTmevHPaAHmVaXJm7qUdrbyv4c+4hp36+ha
w52xLrCCftbh1Q3rxKXkLfvKgW0CD8A5HfshhTDH3hTN77RBp4xoyCvAt3xeCczmGNX/Dtn3vlpA
MHoNn+1xiImkVCW1+ttYLRTG0g3lFZ/z64pRhogOp1CbHUA9fKTpqdYLB6OgjfqUCC7+D6GsFXQZ
eB7KUNqaPi15xOH/w6Bjqtk1Z7EGvvmlW2tcY6Lcl/eob2DOBy+h4ItF+6TGNvGKCRwD7FOY3LeZ
eRET6qzVSZXMAR19ttPNuDphHbo/zIhZ5ihQ9bFqpas4+Rk/NKJzES2AKDSMRYiC10+SQiwH6vTa
nir2dQ50Y0FdiJJ99IIguiWgSQQAh8fAEbyhWf+SAtuOSfSxt93rqKwpCRjaRAqNYkNo7VY62F07
20pBEd68zih3gBBE/aiPiMF0DWNxv0pl+geFFp14fKwRT2f/JwiqHz+zFLldOEV0c8jvtmeCR5it
0yAHgYu/LbIFwomY/8tHYaQjpS5cmZ4DteGazo3rrkGrsiICbFvbrdXEDrjgodzD86Vhm66vS44j
cjkz1iUyAymTvJfwwbQWzeYf8KCLzhrm7oZZtLZ6hWXCz7Xmwm4LmAcJtc0f9pXD1eVYEcYkhmaQ
mG9ROG7vZ3FrY3ugO92sdAUwDFNi4doauUfLs2jE1aoVuESge14XIk/N7Ha/zFVINRSCPTWWeToZ
LctZ1q+PrCswLZHIS8JJvK1U6YOpyVb/0ldI3rUNSUJtpixbav6MNv5szNQMUXu+ISUcsX7NLGJQ
nWAcLzcy8dpGXXuPfk/QU5gpJvtDXxyuQH0DpHBE7RdzR0zbb4m2PATka7Mgq89f0VnfPWgDB/X6
H/oqlk52NRcG93dXuY0lyBJ3uiKaily/xATMdUs8XuFGDfUj/R1iWbqiJZOS4xA1Bb6W+gvHDzcU
8zfQqRAdA8NGPKFrVWz2+5bbCTDh3l9FvT22xcLkXlzVdnbYJz4UH566aVi3cy+Uq9UiZCGz8gHB
Bpr2X1uIuwZ2i5o9GUBkP9E+ib9C3x2ORrlAQBKSSBZNPdLxn1psD45KpMQkC9SebILEOC973tQi
uV/NKB4bY4nZIeAhfFyawTzZ2DFioE27F7ekN4g+ZUSh+PPyJCamhJg4anZRViTWF6JBDCW5T6UK
OobhF5ydz8jUzaX94s6pQTgySDloW8Wd+XtSOAwVdAOHXNSVsotSkYaITA8pgXqwYIKJiX2t2OuH
s4jeh0JD7xFKRsf8cr7ves/DpZdEZmOU9CufkPEJSO4yfMVuRY2Up+JBkGNCTIUBXY+T7hUCEN4n
a/h6AHhY6iZwRjN2fB7G9fRJ/NIiONl0rGUbMjlQW1BIrB9fKmcTOZHhd13eJnaqrCUalrfSYDbB
cnDsKNsgeabve9Q4yx6X+07Y8+OTFwjGHkweWeYBHLu0S+Vjaaq7qIqJzw6NajxsqH4SK8f5Maf6
I8wgxKaDRR71q5Hzo+YNtWEWLfmJEE22hx24+no+0fTKiXQ0HZMdfk9l6jTzSIKuHln2T1PNNR8M
OkfUP+4pzM6I7PeAa6i4G/7gfokwWKbF2RnYoEi70QaQpvSXgYH6/AJf2WEJoXp+9OrRURZD+QQP
qz3hh3zAUFsYgZEKslIdYQEWfzpfptKM1GTzlPvZrE4CabcaWOFBZyfTAsn4EwrbgMEIEwWlxQ+/
YqutO4wc28D/SKZXR8c0IGWsKvhXHflTj9X/iwbH6aHshJPNu7IytBgUmHyEO7ECAroV+MguChNf
+Irof0VL1Xj7/n3QeUPwWkIXGKIops9HFbECWjtap69GzDjNFAOvrziT7oakKc3+q7uMpBFZckfm
YLhMZVlm6yN83Fzu36TIoYl7Lg8fUtdQQlmpcqNa9Et6VLZDY4DqL0B4vj/IrCYMXpm8naEbRBh8
PY3fZgBHjhh1NA6wgJbkAqACG4vPfp7Hp29QzlmD/aOM02kg7e7Kf+6cY6YMgKPplldfdBJXt3Au
jMbc3sVUpigyY6kndoVo1GI41UiLTMQxw5BBEG7/RveCW620nt6MdtPLt0/VUqEVMzlhgqf4yKNL
etVUzdZxThR7/5QVFt2Ht3tDtq+vOnoptwBXLApMN0LL5N+cALfySwjEjo1t3g/IW7zq2QlbWpzi
FNh62RIeA+dl22627oCdV36RHPbtGacPWw7V80Erfxjlj8LneWrYHkSAGR0VxRDrFm1zMMhA8gC+
koq6SUq7sP1d4VLv9MxpK1pM/kDJlrDDEbIVEhdUIrvtI3tlyIAuFfyJegl/xogLPfuzb55VY8SA
CYCAs6cgc8O5KS6REKwqxS/OH6yo8hMa4jg4++za5WEu0LE/BKelj3CX3uMTHHNSqHJIOquVRl8d
vI3TCFfTq+0USlhPYNjylZBmCsePshKXO2EAj/TlWpSiLYcvqUt1Qc93FT2rhVN8shtUmNNZSDP2
sshSZsQqOY1FC4rK+S4P90YD8lloSanbqW5Q/vADuc4KfJLWXQbMlnNdkI0M6fR6wzr9sVTFRiez
9wKeELctknJD6Ko6+GQYwxyuX15N9+vaJdK6Z0AJ4lsU+/cgRzTqvGhSq7vf1RNUU7zULNBz0I73
cOsbHrYFC+NFH6E6y1Gp7Y1/JadPY8k0QSquyf/HfWEj1IIC60SvpvycumEDz8Kny5Oj5dLzB8Ko
HxAb/msLAD0vQ3jNvnvAF5rmJQ8nNr2MTMMVSD3wLzHP9b1LBa4tZQ2sR2XVFLtY/VkUp5xiWx6A
Qn6nlB6qE1vlJUoQagi/KCUd8XnosM9VnWT27Cp54wnhayzUW4zyO9We0lPGwoZh8U+OI8wZN3BQ
Ka1cENYLRoTcRMO6KqYaxDXGWUa71c+oi9z2aiu2U6rTB/RqjwSKxnkINlJQ4Hvumt9OxgvTQj5v
PrjQV0yQuYydebNjVsk7GcMwbFgVViPjgsTk9+Aiay+e/PDKhxpdgiJX3j4CGfFRD4EM+pLKhUkd
p36Ybt6Q0QT5+4xDvHjxadBKOQ5Hg2Gbx3ELBavFFYwq1csGT/RiZxQnLoVO5QHrX9cHQUp2s/7G
hvuSJoHImhFzxk93/xViqhIyxTL48D+Btux3Zdoie12v/NX5yM11I/QQk7jhXPXcgPVbBX0iVj2H
Y+6yDa+S/FTwLbN5THfinwLdRvIgWAFtRRHO72s+u/FcmuamDp2G+lsKqoNvNbk5Dr45dOCaC2VC
kUq0L5VSm3EAkEXDzZ3WyJjNFk7bWiEf11ejGdhR9klADQZiOn2LVs3xPoOHf5ssXY0qfUYNtZmA
SpY1tsA4LVGAtsU7x9oWXF7pK1T++qa6rDQX3vAZ7XypjWsyC2Ldl78/shedGWsgNgBXfbhk/Rj6
Y0TPo+i9HHHs1cAxkyoRsKxoXR6Tl+KmGZn/SHsG74XnyjdnOqNmFGKgz0a3NMgKpPVCN3oeqjdD
uxH6HzRrthY4EJARyx+qai7Gc2C1qXewCHF96y6xNz7HoPuLsdCdIBBhnC6h9q4tuqrd2PLrNlu5
aJwjsIAavqsYWhnBk7rGqfStAxxFv0dpEKBwvqCIxu389IkypwXcBjfcwJwkaBh0QCs8u0P/Czw9
0x5fgsj4zOClXfaCOV3Yp/H8+2fdXIKkN1aN27VhchJhfCVrsqOJVpE7IQie8Nr/IVvD3Q9czO2J
JXroH6N3h6fnuZAhhvcuQecuzpBQWdqChdHfcl4vhxzch+oIMPHsrZ5lL8dhmoM5lIar4I1ekjVP
SUCSlESmswJm75T0cbJ38uYATwh+dNygMOPPVAnMp/VjtNZ1KcELNKQ5j9xzWifYR25FjIOViALJ
ddi+4SoAdIcuv1Ueov4Usns0Khiom+lfs4SMw/XczWs0z0o3hajXWTxtLCrqVoVr61gem4a8A59X
rmSs07YJPfZ70F5R1gqBUaY52h8+50lcEL6hSyXrGu3bRsAj0p1uITzGj/CIWPQpjmHzHlqUPgU9
6ophvoRpDnY4H8CPOs1fBbUtQVr5iiwuph7l8HDuCaxJ8bCLbDhsLCUG2w6s7CXaDuv3d1otiWBn
c8oekpSWOlTWbcqDCHfQFTNgc3AsEq2HYTnYTA64x0Rb7T2iNbNccLTHLBh0PIhvO+xwsG+cHCya
s/ahFgrdKKYpvs/rcL3tMZ1QKB9TaDrr9yjk8yauzOhILfbLMgw2wXOsIOHCUkIjZIA/bD34fSN0
a/4A8pIZzjCmD6REojo9DmmS0qQQw7MTpSBG9duA246NIpAcqzYAwCFkBlIzeUI11TmLKRbCm5Jr
tZJCixlbpFrkO3P/e2sji5fd623wqhoHH3Y3b3dO2BcA6KZC7se9PJPPaQ2PeGYbk7vwSHBpglt5
grornQUQV0gjd7INi2/HLNObI01SSlNOC2zcDBBy+6dItbLvtJWKTozWSY+T85b1RFPBTMruNFVd
WYLUn7R1Jz63FnDjpAzSbXxWZg6W7CELpjE4MuZoEJAiUghEJ8irCxLTVQgQG8hKuyEusP6rToVK
psubz7/+uKJ8f03KjV5rFKqUF2PM69M5MB6/WdbfWRRKDNv5OHm8Eu7YAMyUp731ljIjMM3ICrOu
kY6Ze0IlweTs/dgpW5c1vGTuGm+H8jCpyi8zi5CoH8Y+N9D6aW2V+qluDBvH8gQVhS6IMMJ5RoPv
Kn/zToNmpLPHVBIPaqFE3/0QNtGVGygBYFPZjtDcNlXaS5mOPmalY8bLMQaZepjS7agBjC0nCE0R
TYwLKz1DMpSHb7E3TzoiFxzxElesoet9YyAyYIrGJ94/eyz919KLWj6dpqnvsxok7t8fHOJaN0C3
7qcDFJZo5nwLWzE0re1Cxdjse2+eH+JFw/2/gdA0t/lYllCJhCW/8zR5Dj3dR21dFJOmCcMWr1Wn
lXASkHsi12uSmUBuAhS+rcfNYKuxfa6AwRz/IDM8wm4pCn+2ek4k7HyWqSTcJVJg5F+rxW+BY+EG
r9/ztWIqusm1Qap90+VIKxpU86LMJsyKHXRjd7sAGc54mGlN+u40zIbCP2/t/yAb9pLmSOEQQ9Rg
d6+UwI3eLfPoJjem8NSXvQnmQ2Jkp6rBGs5hVpzaEaL3H59ShMG4BUZai0ARe6ZsHoFFqubGD7sO
zLpyDSgrPKavE46281f6pyoSupBl04aBGiB4GnmLTBboolqvO5Nr301o/K/8DnoJqVtRL4aTOZTv
iNicF+1mgWPx6UE+r5jecuo8Xnan9XGfAHKB0KR1KIxGH7kF0Etaj7CrZX61gLaSHUs3jgTzi0ci
t5Z/YeFyViQX323O/z+KRmfq3YOKYF9lIAfPvLBaPiQnGv08fdkGmk+D//VApEKmXVOpXKgpXnee
+wR5Um6tEY/W/lsoC+YrKHj6tv5h6bPeUkrRONJohQgscJ2fxjz6NwHQMYmz5MrKBWt6KWFYkARh
eVCX8pEym0saApQCierw/VzI75qqbunbBYa+JgamX2R3l8zwGgbIE/AUt6WKtLH0wRAAJarvpCEc
Iqcyrg3sQIcr4CpL4KHI0X72yQ5Bs+SMYIJioAa9s6bQps1RUZxEyyiBrgMGnbcNPi/+tImJxk2/
QXt2t33R5wXTrZgbzzQFjeqhjtqWm/yvcSXfvSJKeeLxBvqNfLNiWbP9K2poJ7ddbChpAUjd0DsR
dNSel2FIPRMRXJ3tlyuLLTQCTzVC5fMXYF6Nc1JdzNvKAmKrl5MzNtswKsQsf7z2+jnvfEzrNnTX
LsKkgWR0L69Vh/XsXK4WfpgzcbQ63NmKFaArTywAGQvrjo12WpjpE+xL9RdDwa7XKvve1j1QRh0E
ZkPJBUlcg0jpitQeKBek4lHHS92cewk1bHkqj+lQFx6XS/hZcN3ZvE8HY4J+gcZmNfOztagU9VwA
UVp7KWfk7zZCQwMYsTYTNZneyQpryptzbGatBGQcd3HJnTyAoipiYcg5Ns2tr46QL0rPFXlrEebk
P0jCi6JnvNtXjIZ17/kNV/EsCG8XBw8zV1roH9uuFk+j/Yl46nDS6TYQd8vOQH7jgb4o43H9PYfq
5x4+/uY1VCdz4CvJSmqh78pkU3PCM3y692GCJEyzXABfVO6ly78xY5bAAtbSU3Zk/VhG+kxPfnZQ
ko2uiyXMadKeptJfLmhYcTNejH6qO9aS6TFFkMiDFIklD70QnVACk0gXefXUyKhx3yph2yLTHUcA
SsLZCmB1BW+EovHdo0MORN2nBxvdrohvAnlOYqtdXErph4zb5MxmzmbFxrMkWcxr5Hhbft325Ufh
YA/tzj1tVHGJeiawaXfRgGSVOLrbGNVjQ1a/aQZb6UtKR5L/iCtwh2lTOV1XGTJDnz1bdUgA6118
AnaxrGbeOBXH4g98Iwpk2SbYWWaF5mdcS/rgF8VnDkmqRH/I9/tdcPLWbRRlDIX2HDsScATNYgom
ITgVoWz9vhGJmOw6Ax5YoIuEsubhmCxY++eeyvqVorN2klUWSnp8Pb9ciUUk34q63w8r9TV9jBzq
1xl34PFL7HZt8uPhMDkSxmlZx5LMX42jaH34sDpBqZERsRMQYl9Xkll8uMvbW2lAscRFvc4pY/b5
U1VYTHPid6hATdEjJFgvjud87tMuwlncuyHgZTFExD5yZmck5+08InuRwq0JicF+QFohF2jQhsVZ
YUsWvm4nK6HcAWS1ih6UOnnhQvPKi1YVAtbO43MQnuKgu+ZitfxOgBLvk6QC+oYGt74JdINXJyFv
1/pDRh6g6Mb6HGW3v8y2d3wzLAFoKHzIWycEF0sOlZD7ML0Hp4C6J19IodwUO+moXhdV1swuSNLB
FxvyD8jfHAC1DLLn1d3SipSdpzGpzx0rlNWlHQMWuBtjOtWDLghJnstZL+CEe/31jWju1YmsiJrP
s8wG4nC5sd1RtQ34DfZ40K0CyCVvZGxU+kIbom3cdNbuGLHrVtJAFAYN6UdIZK/NKniLkwnsr7uZ
BWE6yoPi3ahQRvMiN4jy6aatVVtHSpWADcPVSapPHIt+3qbmkstLOLTrQ2Y0tfDNx6047DqX9SUm
jY7s8aYeDV4kd1TVmEzxX24QNt9TW87mAT6l+lSUdB9PmWP5XOr1kfhlQyROvefS/Vyon/A7/9Kd
SW9kAhX/Qg+TcAedH9/aoBEBPVgzKbStfH0mgfICdzWFWiJa0P9Ei0ZVyxLZecq6xsqyS9Fg4nIG
SvQ6BzduBuehaiUMFxuXL9gKooIRyBxQOMMq6WEYkqzOEz60ANDxq90cjwiAYsdIRe53Tz4565Oh
SddtGJP4xwkm/rGBmxw4Fb33TePdzb+w3i8c2Bmtuid+e2BGWIA67GY3zbjj+ga/rYaAxwyjvbMO
R1/nBdA2DqwoodlcffiC/bm4q3kZal//QrTXJ4u6hf2jvmOgL7AscOWxN5sQm+CWrQdZ3hpiepKW
e5OS4CBrtbzk+aSh261uvVIZj5fyn4MB2qMeHce0RMcz9+r0PEOrt2+fcs72ahtMBBS6ADgsWKgC
RVQiPf7zBsOqyH02opHCchkiIt4xC1YTKfRizt3B9UfJUVASq9NqzggmOtMmxIf+nC6eJMTU5iLX
kxD8snFo6lvGLG5Mc3tlVz3HoWa6cssUKOJK6mnSlE8D8z0ZRtqJPfJApOrBwsFTW4cS9IIQXNAA
tcCKqnnW4pCrynpLAizI/7mdI/L2bYASuS8mrRm/KuXpNrUquUilLUE0mxy7tPIKHv4eOLRrL0UK
FWrTeazKsGf6l3BwQvYD+chboT5bsm6kGQ3qf2xJUh1Dt7q3TLmb+9x4S8tclJTxr21CThTTLTA+
76Qh4qOzGvlo81HW1QNS7lM9JfMFTqnHU6GNEOGA87UgbUI2k0IEcUJTzr/0gFIQ+5lYGxDlUppk
Arcvda7XSS6Rw69VNetniWsuohlRQ+RXPAq7gd/6qyOCs30z4i0rsQOyYjvR9f0ntThGV7v+4VYp
IiulWZlibfpExUkzN4dEbvwB8UaHAIocvvGgtf44tttcaxU14UnP0aryl15kOj8lKZdSgQb80vv1
wDNv0O0W3mjLqWRnJuPo1dfN/j4uDil0xdIKy/btkSpFprTOAz18tFuNcqMAjbuNe4nKhFEFnB6N
pt0VcjRgyAIIrwu/BMjuNVErJLx0mrSHKb9yemRWOnT9NF0fVz3z9C/qfpFSQicyo+lehACqG3xv
/9EJ+HRJF677Z5Jnck5HYwTlMMMffkU3NtRN+tQlxkWodHXqhJeRA51QRkHYrjWrpB7WJqH2o40S
ENnKkfbl4EUZ/LYB63cPcgNjwcPb2lCAkLAZQ6/sdfRkvIQ21Zredb2PNeI9kPydHrWkiasuy8kx
FJ0Rhs0mbHw8NBDJw8m+Ns9K/1Bkwnh41Pcnlj2Yul3D1oS5kT9L+5AFCbyH4pXP1c2xTNmouO/1
d5ZUzZI3Ocpx3Def36ip1fav/5RsGvAIecDEPcJCB1/Qrp3VxH9q/c8yvh/PfJH4uVjUOy6ij6T2
hqx+mM62V0kzZPN8J24bZfEmY9i1BHjxc5Y6K8GfdrV+3r29jvJ7dZRky/1VtP83IbjomeLv595k
aoHrU4oFtqskClenk4mVNOQ6l578xZEdzZ1oF36tbf8yLRGgUPoZYgqJxkf0tktjWm1GW7EhXW0d
RqF8ldcNA6m1b9QGQH+Avq5F3s69PGAcwmtHHuQkxaOOiX/gh3FQttu29BLMxwnhbR3wEIccrf49
FQFA2lQb5sQTtHhikLhoJNu0nTfTN4P5fdrzP7TmEiZsRT+FOFPE6uaoaNmbTfKFXk9zurE8uNQ+
Nxp2uRsP/TPfEpaQFqsPdNpzAf1UgRdZQ+kmHW5uACcDKNhi4f/t1LeX+aF7z2/lyyqUgaV3sILM
89JqqE7c7UEIXZyO/WmfOfD2J/7WrommYdvfvfEwAGAmZZRChzCDaHqFvGaUKp1VJjEfJw2LK0y2
Zb+3CNz+zWHItFkVYVO8oeJh/+M3RwNFAU4Yw2idkpIEYBundY0kUCAFiNS8ubN8ZXELahKLFigM
u+xNiqZq39GubOCv9OAVw2n4cpy7v5FDWgCpvJOZMeENXgk44cYxylb1j8orfXUq2uNgk/D5+5qb
KMIpqH2qc2ccl5aRj9YnRPgOxyRef9vKX67mOC5KXwqaYtq809sYNUu4GV1QLd8R32wfz85mKvcw
ujVlizRhau1EkYqPgU/+cd3We4J05QppQvW29eZ29LzTYV1gVVIXovSXyMrSM+B7KfjA8f1xlRZc
drTmr77W+JqeTgRrPRbgnDWcUxw4sRgAFznMYC0q2GsZEfe38TxlQcnaS00+eijUDut1I5/SC3gc
ghIYcve15J+IUm6wnttGU/Cw0L4HvlgrfzVj9ckt1nefLdQkw1GZEQw+JMQUOTkLJSiQNQJe/U1F
jSdA5c4Tn5kN2VGC9GI3Zmt443GGgo7Xi61yJnXNSY8STBBGuQ7U13czxvhEsMnMKV11dYsXHrMb
2TBdMjYV06PqNGBKNHMR4iQ0ViSpU91FP0kQPjhS/dlx4qnLkJ7YWIoeLWyrCetYKt6PbhLIgR+P
1Y+HV9rckooJqGG5s5iZmGYcUi5ugVdMHCGyMrtE24MrnRFoN8wX/8Xj9bNSXGlS9IIud3L0yxoT
VBRriPwW/j1sxuVfoUrph6Vulnbi2b8qbwcKE4IaFJ+88NypoT+OhqPEsVVAk3GOsT99g5LyCETq
dT24kfhqB9+A9X8P3zRx38HsE3+qHkbrVAsWIonDv3usumvBopSwFYthFS+OJ5lD1+vhQKfe8muc
kIOCPHOxPKQJFvz8lFX7xBoPJ+UmZnTCs58AspzpVvtiH6DqTQA39BWw259L5Voo2QK2CGC55fYo
R0ygSDXpypgIAyLfw7wbOwYtJbKt3VzRVbUGQcOyTSTFkNgkiyjOI2dqMymD09lJ7jEtvodgHuHq
FeKlFGY1dEM6C322VJl6nvnaCKJZhHyxAvDgBjU8GWx1kSfXa7ihu3QO+FV19erPHRieRX4paQNl
wH8ll3r15CdUDpvnacIZzSQnWEJUTCEUQ1Y28nAMrRNsbm7l03Oc9UqONc+1Qp3O7Vi7Ft5lEoua
EtsLOg6Phaf+OIQKzoD8AGb5huSBlLzgAAoqzrPDHIXSKPG0htOSlSaDAa8qYsfovX3Zb0eH5LIS
dp3qldyegy//+Kw3n5XKcs++dunhWHjRayV6J6PosJPlTuVl/k/RA7zPV9s3p5dBva+Mn/qc6NxZ
VwludqqYW8RFVYFyx2RW2uPgMasnMesc1BeaxA9NQhIR0tul1VXsDRoDH1GyqA+du9gekpebwudL
MoNXYwlcPuUAMU4JipsUqfj4Hcop9Z075ryD5mYF+L60g3j6nflVyEjtlbEnJHm5Xls9B1f0Z6UQ
deIWh6OLiz0TZlzLmIr0zgL12vevY1bFlVzwTju5dte6XOw+ZgrUIVPLLN/z9+n/hh8s5geUvXge
jYEQyTmrCUjHx9cfChHy1N1FbP+T2hz43B6wPphYN62zO9Wd70kYdrGB6q6RGwq1Sz1BlqzFKiHb
loggpytbRt3uX3Sr69lmhqD2BRJA17X0u9Yt8Gua5qDvCQdwPqnuHlLNXI+Yq/8BEi6BN4fPvaJV
qA7uay67tsbVSUT0W1NJSFJkkoibv/1BiVKAS1CKJwEXq5BsH9bkng37hNn5QOGuqOggu0lPZkla
8ORFQtNsJKV9QmbGviPskTmlhz1pyB5uCX+Owh7Sc7NnJyd/ilAhFukttFtkWGlvXniMldBTcoKN
mdGoUdPRuxwBU2xvvBpAMvoX8kwObppfjkqy+fhK4YPa8Lf18SJaVgJTrn90iDE8EFvEJsxCBTVO
thVni+9JUXjHh72zyOg0UbYappm/3+5b7lZKKcc265d+LYQDrYC/6bsfF104S++pLkcTmp167J3z
65Ftb4smIGOd1Gycf0bKU1KGa41h12kuoKRagoHJgIcyUT2ENQ9CGyJ8hWnW432ivYjBgSnncFMr
8StlV0mSz05c8+E+AH/pzaYXc/9wd0sMfKiJ+IGmJKDGM0G4n136x+wdeGtK+QJHaSt5jam7OiyZ
LbppMY6+E491O8GS6NgfotryCo1onqr7ALSdBdhkIsAm/VT2wwh/cfyIxRP0tGtJ2AdOIrOTLray
9gpEgobolBjwwPAZlUHK7Ap5UQToH6d1Q5ACjT4loGZHv/qoMnqSTFb/p1xjrLbnBGHv0LMqw6Np
JuZGWK/A89DBXdWsS/KSVailysBK6eN48cD7MgB7Q0M+RmTArqB1pxePhFgPwK3QBEQePYNSSwZD
jdmmkc7rf8yjb/MBclRnQ8sBzLGR7CADDK0p6X/v55FLNv/Wnh1fxIf46rH10c5jd1XfPRWkNXd9
dxdFnrhtfzq8yGnjDxhPz2Q+90dzGn0O4j880aWIa15OmsGqcFshsm6K608nKPEWPaFc2R1L1YMH
pIGgbk8howOUuWbtdOeMvuvAvDIxNn38w7oqSJM8ZUVoIA8aeB7vSutNU9HTW+qymUy/jA6wUeNT
10hOphQZQOEUeDOxAdrUoZT00VErlUu/g/fshMdiejYCWwRX+QtGQ6fkvbVn7klnXb8icWIXwqef
AqUi9c8kG2QnzF3t9N8IfW0ECo41VDQvBGDHqrLuDIHlFIanb3anR+bTGRM4hdKQ+bbBPNnfYWgU
uJA/pyeAj1Ppvi7AkutCJAhS6IrSJ8ta0yXiighiJpOJbpahbCQ7wFc+wOKhddocrvdRaDE3BbMh
NgaVxqSot3x0LR920JV2flIx/NiL0CMm0A248foUTCvY5E+jOMzfyI0uu3IaUVxMU3PgsnjKQ5vy
+UlMMTm7nCQhHCZMEADT+/n/U3oXpFlj3nN1qy/FqP9dGZAbfSjdp8/+3rPMMHx6gjYG1fhoSnNq
tMzGKXBu1OMygGi0PpiZu3ves7ElAzB6KyLiuLkIPeiY1Wy3cy/rr68yiL8rFhDLMRufhPMlScOI
nTsHWjKf4Bcubum0USMLZ13lWoJyh6Xq4GN26npkETltFcHyJHNM7kyKCZ5E4zHswLux/ZvFLO/g
7UujwVZOD65msZ+FjnU6hIlyi2LhlrOG+4BNZVu7ghWYvohdCcltby11Ruud9IuSNR9GAQoK8ajX
qdKYYqq9+G5wlm6wwzDdzBqxDF/V84LkT6GW5Klu2widf+MPZgCusNG+L6g4Zo4QClilWpUZM9mO
rX7EchwQKPvIrtL+Yt6QGnbeyinQSCDjBhlEXJ3S6V7s20znDsiPIXksKlq+a+jIAMRIuu55NIAZ
ZYUIePjiLtq+xxO/4mVjRvSOcwbkUCyfl6G8QPxmt3SLleqtM7Gpv3uGLGNnnnhEt13MjpVdeVO7
WEGZKS6oxvfWmXvWABgSvoAvfbKxbFrvS7HZiHp/r/oUHdXsxbhz9XXAjVjql20QWMgw/Rxhhu9N
X5DYJ1v5lhEb5zzv5DncZ/dquZAzY+mjDwDgo8PRFeXQsCFTarp9+5VN8GsF823lInjwmweXLh8j
NrtZMGWEypUfV0cl7a5lyu95a7zGdi4739Tx1M9oIfNME0wVZx1aFt7478hqIVgmMfXoJJG1NIMb
sea8Aj9v89jaeFI4tNoA7KB0hhGWjxGU2+H+yyIyjBxaHkZyeBKswfNkyTjSrx4aQzqhvW2gBlC4
4Hz+yG2ZOi9Y3E3jd4Bg3kIp+DDwa1bEdR/hr1F9LaKvYLfq+c9G5rH31XqzX1daWileKNNbjWrn
4Xpy84bajmLVJR+aIqHHJYxVfyBhblt/z6CSHDuhPpsPYpRJ7dJwaPcs2M0nUkf1z4CIhXn+MAmY
6VjqiUC6WE+cQjDTe9NIf3jA7IoSkVMIHknbApIlWPtWZOvM2/hx763R/q9cvwDTkIObN7r6230K
cdvw3HLLSOpANjNErmPEpGXzbeDsTa6hvLcza9Id/g1VcQzYKWswSEGNfr4IB3igMFgPCbYC3MLQ
/WUrWxJ8WGJsOGsGKS6mBq2VLO6KBWt9s0XwG7cvhzXIHilXTD3bPxFyqQk/YP+X+9FUXRXQ24HR
Tlo0b7Adi/9mABxxHYo3bPEvJUDtsLS893JAEV5Lq0UqHuE1yr9y2ZySnYVO6QdKsiclQc24rJbY
iTFC+DA7ITd8tZKR6Ejzt+hm2xI/Ihxx9aYYTtevch1PGUeJwHLYoT9vLQ3lFhYevUnteRNkQCFT
xrhLAmJMdE4tJPlJqLSidYC8EkvmAtIrIQBzBGAVA+5OhJZnPfnBkOt0nqaDq76wvcncL3ehhwzj
pV63O7fxAmp2oAX4QwOjiHwRiuxbxJ3C7wMrYOznRoHV6QNEMB3tNMWHRddkGxMvostL0TTEuGY4
IQ4dGCLn5jwcZ9NfLDkaMM72QyGmqYKDuCB2VpKUdvuwFUWjSR+PXmo5tY0zBX7AMeHqxfSj9Qik
Z8fPGT5cZdIMpSidJybr5msUNkjZeeSaR79oPYRUjiyAkvfr1K3zUjrS5S9wOAPV6/PG/3lSv1nJ
HyGG1x+SmPJ69Qla5ORSh+YZAl/Hy/YMijFDmlBQtQfj4Si0bKUmkTeyZ+WixzQKaqeIcUW7fjCB
O1Rnvjsv4ZRRjOJPRcgWQuAA4rDRzjFb9n+KoCez6wqAPyyVNi5R527EJ3Nx5BlSVGoVxuU/kUkd
DzpJG4eUV9N20tqyY7rpnwyz+PWA0HE9k6YQzslEH/No9yb6nDJL8c+dXPEwXaXaYEdZtO/vx2qT
ZwBavEJ+3rrZRpxDaCsqAk4PBN6GE8WwPbSX2ewp86Pit2XbZPX0l7wKL3NLiF6thke61GifqS2/
BOHborr2VkbjXHsfNmtQUI0oa0Ti2d3siJCRdrLqpPY1ayU99SFKHPVGd1232weXaLXQdDyGS47q
iEXOgLB85IxVU/2W1iAvBFzpgZwmyMuqMe6aXDP8HVjXygjdKXRN62RhLJfZr0WPQo+gTNBVN34E
yN6PEYV5yf9Paaxcmvv0ZuLQkPn5mNbJWpHtAI78JnEaWwGRw1aohfMfmZy9vDDMVEfjiup2zE4F
gWPf1sp3kNGvhTJyx5TMg1NFAqLnfNiR+d073WzPQwOFw4dRZuJ1MfRIzy1otMxtpoD6HDMp1ZMG
Cxf/vzVy7wjofdOwz4yQChuCDR61Qo8dWbWJMUWgLJh88P42qa31Ohs0HJIad+nXbnODmeBWWCgl
2Emd8t6iBq5v6hutDNnKiZjZdDZIT0mD9WUo9kyWTvsoW8MqfiiVD05WuQaEp40XRdErzZV2p0OJ
5XRdRY1HYM0zw8ixTK6PxQ3p8X6iXYyxJr30TTGlLdlkLQxL+NSe8QskDWmW+6PEmDPFE7DmaeA4
UUpdobQSFE3dC9xBsGlCOyMrZMn5IhRP3xRs+BzgqCFCZ3hjk+9FJnaab3pH1VmA+aETzqpa3ifo
XTKNRVnHz/5BqI3HScf/yWKCER+yWb6FEkdovZuJlBdOJZ/La5//eYbue56DZkpyRjLOWBgrmsFJ
ouw0b5rv1ZiB2zcuVf61fC+JFDUFpGuGgE9uFRS7DQgtu1rZSNHD55GA81MD0T5agUIYW3Mf10sz
DIWPQOE8i+nbqjwQbogiIFQI9KoS7e1SWUEW/HSNePEkUkq9X4N3DhXr8YidW0ID+Qi9LqZVP8Fp
mTArvh8Dms+8zJldtPkWgUHPb7WqKpGCpgdrZjoOgmUEUXtUABBAUSeM+bgguik0ceCRDPcKC8Eq
qTuwQsLp8y8CajQjDbnaRJMWqcLqxfBQCUMilZu+hxLSyoUQ40wvV/7IHNYLfWPhUaEx2V8ZUZVd
x9qFgrt1VY7CJvIEt/MAOn6hmXHM7q3/JsZX1vefn0qfcoXMJRbrcZJYlHYLRNsPRWcjrF84lbFk
RRs0eznuO+41GBRlG4Xcl8zHgOr41bornDwqj4iHJRi5ZBZaONxgJrPEU70dMVA2QRpJiUHkKmnD
RJfCP3Jo35As+gwm7SGi6ndsxG0N2o2pNv6XS6yHLGCnkslWdWpLtzfFHzapXt7lJiF+k9LaAjUp
0fXUtz0S1fBe2x2EV4/OZRKnuBnt3N5C0TTJwlcqoxAGUTpf0sQbyrUkmKSzEz7r+vtPntzRDHjN
LAT5UbApUh6+5vLeDK4IYsBFIVeTFdJd9cC9F/sAiqEE5j/EsgKFWzEPKLE/2g7ikdZQCCwxFxCy
mRI0bdbGbiDnftE6XsgaiO0DZZT0OJCiHmr6pDQLSVyBhlptDceRTVaSDAWW/K7q3MW0RfQewZeX
ZShw+vsfb7qqFbdedw9laJG7FleI5ZwMT3lUQXxae8HjDHiGB0xENNXeWxNtY5b/5Gp//4jv7KXg
2+U+bgGe29VIjgTi2EW10uyuNOMGnKfpst3fQu6M+NazG5Hj8asI8hZb98kE//tdH3NONoxhABpb
ffyDymjKfQtaUqH3Ts8JLGGywT6w1NMP5IW3RfMLEut3qFxgu8qGR3LYdNJqe9iUpNq5sFTXGwMr
BKgmBCvv6GLianSsHgMIimUikXOrRk9b5C0M1QJNzRY7Y8CTikYkK5KxMb7RkudVc3dd/tmIqIB0
47DaWLFEIhRCoEMit1ji2glxE9Dpu3TLnXy2b1R9tXnMe+11kF1xZz7tT9OZB10+rLkU/cGi0ZdK
+jiudISY4SlOQQtXKuQynQANTeIOncs2VftXPKaVgpAmwm+4wPmieDHpH9Kyh7FX6vLW7UpmbKQI
aW6WO35cScfQi2+GoFFVU8kwdm4UG9BGV/2IRKtOZVRi5auN/E96ZSJahO436OC3iwA/hU5QfV0g
q6FsRraTelUxKbzGt2LLS6sV1V46IP6VvShNQiv3DTkynpGPcjyibZioAXAf2d6CrK9crgbPiLdF
7Vh+VMqKbSkXvPDMCrG/gWHLof0o2aEDAlptZi2rRr6QbOLgR8+jrlUZpsBg9Ymp/nLWJGd6yed3
HCuG81QpQQG+oRoiMhrZvGZTvjJmxp2nQIlnZyE8AHJ4jqGriPYnvo1eCRL2KJ/z3uLZwn88OBnX
EdGF1xfusvJSnOhmxgkQq1cLP197CF2Xb4N5t3BoLapWXFZFP8Huuld7lEeZgTW0/6f55MouLrT0
Tl0JLQkqknEEiqo/qTzLPIcpBClLD9H0zQXKiPE219CXauNu6w2235LtDAarUZQ3OZM0BN/6R33v
A2Kjz7iSMpijtwdwm4H7BGFDgVWgY2K9aTMEmBByZl+aKW29U/6AuJKc7JW1bAUKN1N/EDAVD1p9
KOKhr2Gx8StWFd5DS2fB/D13KcNrLwZ6wmVq9/uWY3b20D3rkkq41urcz+ra79UnIJDSZzeyMNUl
4ZKmTST+4Z3bnZBWZwda4jlSQMI/Vnap20g69/U3NUgfIXTqniTroc4ckTeZBFS0iAaqftPrs17U
SSzUty458l6mdk6ZU9aaXoZvIZSZHvq+Ut7rHZweDztSCKHvOm63AKvjkLo2qdhUo3iY6dAhRdpt
nZayx6T5tmYogFUMVA8Ye83LjpFsqfR8sfBHrekr5rfirpgpZZFh/wDo7Ors8euon3Km/5vp0TAp
kVji4amuHfN1Hw97ko/+UQcg5r1LjxLlGcGiJdV2pTdpCaEhMhLZyXDjeIGoHqMgSGaEyDzB05kL
qJZx3nr3yfY9ynE6ZXGF0lKOcdDSTRvUwAm0GP8qeFHIo3aioszXmmsiW1FRheodjGFv5EI0rHVD
1VSjpvDu2CqsjTjohmt1kFUUOs3c+cZMOj9aM2N1nP8TXztaaR4LFq6ISdkGw00M9rQIKaVmW4Gu
pdx/MWmmaxfG5o1B96s6xUymBJmqeRycnl2iAvO4mUP/lO1ESAQd209/MX6anq9KsBU3vdd2uPVA
mkXundONXMjEC19DmZA0qaUzcPDqGhPtajQv1pCAhfqL4SEeJ7BhZiT1pK9aPhsT/Iy6Wu+Eokl/
JGD7Wt5KRCyCOfb626bnyRZ9W+c8EjhRIlldVZ2LbvpyrgENR0rKps6k9J0MucMc52PfKUxm4KzT
TQJqiio/EXv5MW3xa3HRaj+HMSq0gn8PHi7+BrWrtuUjfx46f7fDk6qg38hgJhiGIYcbDPJnx+BL
BWQg15MScAVrMpcr/RUFbJ3J5Eykvrn10jqci9KBoG658FsIwH2FFGp9TRr6PdJV4xZffOepR6HD
DI4oyLBp8aYkahr2TxP3m/R0v+fA8nwM1hNvW6urUe2fbtRKvtAJnb5ICommOZyOfwFUuNYWBDAp
1u9wd06TnglpzwUmkt8NBoZaS6O595dbozqD4e6TtoMPqFrdURuOJVfua634vMWvih0h9A+CAd2C
KhNlBtU1P7LVga1b41ccC8vq+hRDELrBgy8YaewEC7l/g/v72mq1VjP4sJBk+Nq8do4q1KuvmlfN
m5yL6yf4+HBEb56H4SksirpEyLpJQBoNNxI1DxTjvK6M7c+WBwhVp492CCCtexQBA//up1plafjS
Qa7h+VHUQa2On0xFR3kqtDagmZP7xPprb2Xaz5b16o69qWLKgCkrYhO3emKfaQ0ErcDyrqk7lAqe
TlCPJlK1t+B5ixcWpOhkcmDHXyQosVtziNQ27ujHrD7NRvl6jDlo+Jh1YcuDQCzp91xXt5ZF5Tvf
SAV/aTyF8esJsl4aiXU0hVCdBzXybRpDPjCxpZKGOaCv1yg24RECgHDsh9iaEPNdf5FM5XokxSjQ
QgBPRHrBlPW6js5JbSdI32YKIVddZ9PvFO+i4HiA/bYi9Gs+MCI2GArCNj27vTeh2iiHkZNg5sfN
jUlxPHbQfPocYAhSyKSXobK4rXSNmZCyFKGi8QK21B2inoUwoEuYazdK6Lggs903K846stqKhYUV
3YR+zlCHijDNP2bEeqqJST77JHjpnSJRgqBeEo3l5msInqyK6M0G0neM+B+YQFhmmRwpNxBVoYy+
r7M9DhGeqDg/GQTrjKvvg5gWWrg+xRxN2I7U13o5o7q0DH0uTgeFCOPYahEnOA9pLyNba6iAwmvk
WwqewWyUUXbSrDcdsI1RnC9N57PHbSBOeEKWiUnGLsKYnbQWtGEZeiZqVXsVCxqrFgMH0pweV4MZ
VTxc9Q1NeGc7uJ9jwv7ATyue8EHcZO4QIOmQ5ix/aY4YAtM+chmKs3ip5hwYNlDYyIo+zgB4e+bd
7gx6ObQt4ptAFPgNrO3m9h1bfm+IVT40ZbnTO0PgEWBvlSkBxFMAon9cMDcZPyZg/yyN4pIVqq9G
99hJ0q/ZZ6IwNjjgxnp3jZiLISVTQPcR1clD5pm0owmaFy48c1HEZM3B5wbQeGdPV1C2seIsDl/g
zq+venuN9tH4UiuyKxyLoum8pceMt+nzlfvxLwryQ64ru/zatlWrSnk0I5ZXMuLrC6nkRnxZeNhh
16AEm7xCYqLSpnYwBskNH3FYiDM6WaRQlMkSNFukoaibzGR2iGl3LFJzzKyRnmLuSYS4CLopBT5Z
REKK+ohQJRFupNfE7wKklq2ireWkKA+NnssesefCwFHlA7y1mCNLqCn8JWiVDVyxnys/uy8Id/1W
cKZ27amraI2vS/LsMBtWOfQpL7TKAy8P+SokktDeu5LsjXWLmgXMgcLZ7EUG/LPZJBTe9Emd49+T
57QlXcKjNxvZSkSPkspzL6MbKB704OrYZEd9ycMA4nTSOeec78gswJWLTx64WF/RwdfofVy462v+
Dqmo26D1oSBGTTjNCW3VALDBcnfAE23+ggr4IRdseTQOqJmaTS808Znw97DA5y+TTFg5P6SP0fR8
mL2dwqiseXOv0OuBKt4vTZORNr9Q3Yk54V4p6HaMwWQ6haTip674JKtB3KmRRBPpPTn3s7SYH0Y8
q8e8CQctyWPzDl6FB8qsFqzCebOpeiwcw16geHYFUvJ5VZMRAoFA+j5ITIxrd9GcTfX7qJyOMggr
7L6+Gsoz19xYhWVXASLJ7jI7IXP/t+guYJYPLNtTV0VHqWvRBJ8/G8O4r1PudTxfb9leWszqdmVX
dyHOLhBo8NkhkVHQMbPqv17Q3JpR9mK1QQPh9OvMLR/8nA7TBiFrlKjdNzG99HsD7a8ORQgpywQD
WAU7m3BKf3BL9ySTrfqxHTIyWGRE5G4ZXbo0PJlXBPZ0iQS1YirMuHYcvDkGz7MP8AsPJDijLdOc
WmzIrMQAuEsxszTV+YcPMoxlHe8/JNrQmhX/gDr7GBwE1fMbJ5EEB2quGXXrZid36xJHPo3k2FOg
DyRyfUD5hZO2G/NnsWheogXRInu7+e5t+R6KMF9Zwp6NLOSeNDjG2xgfJUA86zL4fmRlyX9r9GIm
s+bIv2wrD1Vz0MTxWhCL1Wg69wHNrTUj7A/K5LcmwchRel/Zd3PH1+/6amMOAfPxJ7+zaR7My2w0
RrT7lQ9H0o135ra95nuKVo5haZNqWyJsxzXNbS/LHs5P7NsV8dfhroaUCOW39y1HONPCAcb5Zo7I
Ep+Ba9Tlm49dZWlfocyUQmXxa/eaWFvKhqtLy2EtwILDqsHY2+EBdpI8SDvhnf4ZjGXHHFJurawD
Qlhu8lL8JcH04V7o8+p+Lh+QgbHnC7fKnM/l8/xG9nPVDoIqLdYNg8vWo/R7Srx4kpeIyYtCzJTn
lJeItgE5/qn6SZu3w821x0bTNSjdn0ipi2op+M5PDvauZj/jD7xwQJi7TqZQcojdE1VDF+l3OitH
rINqba6V8x7mTozYbOLBx/8kiLQB2/uRACZ7Tm9mxGL9zVPbTVhIH5r4+V7oaSJZMFggKC+xfAKN
6UE8qwgsWbXgl1g8VkCW43ofTjqfkxlO6YUoW12YK4Uqfh2rsHh8YMSHamNVH6xEhw9xhvW5uhoX
qoULOPJ9bRHU3euucvR7CS51UnRznmO/xkmtTdsK0MAf8XC/5ZlIlomkIZbxownfhfg9FGePQ16e
sDgeQrkwkVwgRS8+WyX2/UNYEmllgrJ3ml3hNpKffaLGUWzHdocZL/1GVTSzmD6ob+qX08SB5j19
MS6v9ekIv+g1cmh8aRvQu7+lIWKlIoufqaWx7AUuVwdJMecm6a0JnckFAkP3iW3FL9/M4r18CJ07
JDU5i7iBs9h8iSFesDfrqPDR5TUnifyRyxUItsNFaXgVQsRx8BXlmpLpmr4dydpUxROtMYUD6NmN
9Ez2/UYU+IZ43gAtAD0Nym2iQbvaACKOS2wrS/3HJmcjJOC3P64SttEMTXTPhe2I5ZLafq7xfxmt
lzvKAz1d+K3X0jh+LaEuTTUJ2y1/9GdV0GKVTxduaml7ZjnWrpiNbl4STCwVMzzWi2paA4jUiqXI
+ikMk2c8aYflVIQ/B4qwWkb+vbUqBQjNw1mKS6DzXR/iFIoDAYnoN/Bg+BoizQJzkdGleIN9PRVQ
9r+PyrmigtgtAU+DJaXC5y1loE5PIRh/a/h724J04xBGob5tGvk+EFl7zG2h6I3Q1R1SEkUsw7BZ
KB9fy7Pi1BBtCknL7dPCDgdo1lfCmTa4mHbF/Cus4RCF1ukKUR/cteisQ4Z75eWE7lm06YuB+d+p
J++B3kj56WPlVRF7CwvBJj7CsZK18x2ZUzEljQ8GQiUkHBklQK+zxxWQExaL0iThInHv6qu8+tAU
nbYV9atmUaEZIv0wV2I3yjg7oJhWyQNDxQqewGx44V883eyigUMwWzAbE96SAXZq5crY5FkFyv0K
97LjqDUubN9HjdCkWIfDZRQw9MOh32+mFqlzqWxBFFLSG/nPMSx2x4RpSkdwd101HklnSXtqsPac
Mo39YR9TsgchCTh0QsLFLoa0xbS7wWZ+u4jKsQRBY1kRxtHhNS8fnWW0vmwS5p/vGfrvAxwlDJwf
JcOoPHNI+azs9SeXZ2ZTXbOLe6WK9iFZNrbK1IO8yhzy6we0LIxsJZBJmya5HCIK5u2/AnZOA1Q/
1PwZbTrvxWkHK3N56IMbOAhlTN7MsWLFUHpeb6AuEUV3eZOFTPNZUVWfIl5XAyF0K0tt+BJe1hTx
XTo9auRntW2QpJr+4y5YPvVCzD1hxlhu7sAxz3zumBQzH3XAS3q8FW+yTIwrUaavfKvO5dl3+aA4
H262yqbV79iJcslNN2ptfPWaCdpI7lBi2Ffs0JpXOb90KZhawPRRTeeJlnF0riXcEei6wpy9PNN4
3LsiqSz6TNsC2PTh0QYzIxOKTpBtVwnX7SYGyZHIJjg72HbD8/FTUvqxRPJVNE+rh4kO2Qp/1BEu
1hXQPAZVdOZD9iWFE+V7HgLgHpjsXDJcBBqtmpE6EAQ9wiNWbltXzHVIAV7b9tyekF+JNdQke54X
35lssWHzJHRMU5KEjjHAWhGjxVTBU5DdpDyZaaWOd4xXeCncnmQqp9rzgwrkWXTCKp2NOpf7ZC4/
DK8mvlwbHl2TLPIwyQjEB62GXN7K4npwk2nu0xtwjcpVoXIlc3LDBbEeGDO6iryVmvHxcADnybTc
9uDbJtFe7qheY2kxAt+3Fd9r8Eq3BMdhya+Gcvr1Y5KA5o6cPrlFTZCxhiBUos69+rfJI6GDMNrH
g9Ip93ezmqbZnGc+Xxn+YxSoC/DflTdJwlwkKlJObFFlraJT4BW5p4agXDdDucvVvdPququIus7v
nDybqMqIerbk/rKtJBJZvEpvIqLw7+9dsaadeq33WfBLa0pEOkLVUSIZaeWswzIeHngdfIaprZmW
QXqK8BxXy2tczcBcbPD5oDBLyToXtvrIgeQF0Hd/xTbUqG5Ot047fHzeNu4mV6u70Dw+e6vA0PAl
zGzDPWm9N15oKiYdZOubpftfCZUXqHEv1LEBfolzm3+ydNFRseMmXHWM3SbtXUFTQEW1wWkZci1T
5iiLnpD0P4NbXB7tPkWr/GzDZqaDzPrDY62csdkPnDbmk8uap87oRgH5ccOOnPptrNMrnyUCgC+3
SN1JcYLf73AM/3nKmmDFbQf99oWWaGFLAjkuIkPhUFh+Kd3QbjRz3Y4PsyBOzFFbhxt6xnQ8lSpt
XKWIw4E+N2c4PIgMRo0YwUy9ITDyj/p5D9KJt2EfNH5uWuQCO/LKxnYP+1JUwwp7joy7cvVqwrza
FyCYr/CJ3bgTf7AfC3HxovEpWppvnvbBoxLAsoChp8O2KNZqOLj++qfwVC+sql1EOVdy/QOd02lO
iRiKGW5gnB2/J3Uo1f7+pqv0u5q8ubIN5Fm7HFJnxdroHUb6Uwy5NFJhtrKTCtsChK7+vADa2fVS
8x+Jq8ZJV0+ioD2olS1aviv9NPhUVzLX9iv8bUKJtoU/Av3J9hXiBPjFDOyvtI0TvlMUHJGr6cVb
EDe0W4CTK3rv1LmPNd3JkjWoSP0aLzyRozkL3LJNyBYdyfu8cpUATi3J5qPyCcLNollPVXq4u4ND
taKyPdJGfDe9fg/utkJRLMB43jlS5T7P+fLQLZKf0ETfigSijyJZv9QeaR5wDpef5Oqhe7zJgIP5
DfTWqkXTyzHyvhDTgCQsghoI+TFvYviHJ6eEu4vAkglypFla1eYrM7UEanOuoXZl4dL9kaor0zBa
PAe8j1XQ37FTkUvu0kSI6NQ01qhvsbJQqu9hO//y1CdE+eAYtjqDZAKL0y4X5uVejsnkUnq85mQ2
uxVp393iw/JbL4InN5TIcBad13t5jt03S9w8KfFVhiMpETOtTiZXVqxTc/mW5h2tif09zeivRrkp
4To2LmogSZ6/f8OCcnaTSk2PSf7y5kB1z96oKSzCXLzu6PWDGJDmTnMHVUPIETYa/TBRwxiF/qj1
EnH4rZetwjhE+Sja8FrSDgCIqIUjMFyJ4O2633sfNEvAoiqMHqs6TUMkDVgOqv1CiP7zZrnxls8O
E7PDGKIXhIlbU8BAQZ/R8tBx6lnrzdb1oQUNWCP8cpamFVHwzL2UCc8W//xjS9//2YTcga0r9Qyc
SBwT5W5JMieF+EooxuZ2pH9HZagW6BmuFctQHGI6TG0sEl6Vr7xHjSK7EtBLox/h8lwPWRaZksHX
ArumPkv7xpY5lsBd6qMVvwNdvZL+75nvkDWjovYPKJ1b+Et8wP8vTfra2FDdng92BgFxTcW+gxL0
h/YNndG0wbsFmOstOUbTuVbeb4MuLRK7j81V4bQVg5p2sXUKOUZpTGbT+QevxsLLLsRwehxKy9dD
rJxxkviOYuJ7/iMtTgvaIKdqYYDhvucPT44PKVdRRNEs/s0lvCV5RnXQILVf5Dq8VhTI4zYWGi+K
m70N0T5n3/t4t9xZ8t11SodHzgvR/N5U2vjaWAP9xEyRY8NeK5fQYhNH6+4SuidfhKuUHMJhJbqR
6NKgz6D1f8viUiKouhtNDn8i5i8vGpRXapN2K+V2HUqRP9QsR3uBRb828C6uup7v6OX1z8DTFw4C
7e9F/gMTsIghYA9hnIaN72plzK+ufY+nFWDBYfk4f2+JfXMpmk7d57E8GeHb5gCL/xdwVVZXTOQD
egSiW2SkH7PnIeAwgXTQ/8lbzrJnGZZ55CSm5884pgiq1jMUjQmN4wSTgY3ne68+VDmjK1wRA9qB
wGmj6EGm3aTKaqvERhHa6VhrNDtL5i/dw9VG6bhBsipvpIyDTYNEjyD0J4fbt84WKhbU8px5clRP
IqwE1De+qSo7i0bOEKw+isVbdzeuvSn58GdqqqKlCkpwso3vOeLa2B2jLYLSaup1DhMZDLCV1soD
s+8RvpY+4L1Ckw7qZXMgyLZg6fGwK2xFei40mVLhZvwBqZrgGaHNPgNAzie/mhSCgtnynk0pR5IG
tZYDPf6rwScRwQi7ABtfPu+iO91vwrIcVL8VDYU3Qm7mfekIqnKRG4bdpaLlijLZ41YtUj1ynMh4
/G+4FTJTcZyQFctarRGmizW2ybcfWo3GlqBxl9Vl3T0H+4bZTQanwkF6zD11Ucdy5YpYV8YQySsE
DJe9729xpV1Mos8o6hlo2DawftVyZK9jRl7jGVywwsquSxHAE80kYdth7DVyrIbQeFBXZUXCyjQU
7IvJX2v04G94AoN5mKwXYFDzuKJLlnxoOGFiTLgbjoAG2tXf3nTYbqtDxLy8RHPmfjh8niGeUIxi
pOsJ0tdBK1nuTAsYlVApAYWNyYRSr32OAAeNY4bvn2f+ZSseGpyRO0bKFD/uxrEiU+gt1M53rv0U
AD/moRZseFV0CMUhnY8leFk3g/++1XuPedampZ8uZe7TP3tzVeXWmjwBQbih2A+2+3tCJvqWqoub
ubJk6piWQ1HMaLiEvQa8mvVIkNRrvsUzCHuqZqcOcjgN8md+ip5DHz+ttYQRenZeW+B2BLXtVz5E
QDqi2ol1ZzT6QG3NAbuinUgAJY97PfVyLVklf5b/AQEafMC5kK4aAy3wbrARuv5JOds6RYKdvO3e
WUUDZ7whd6VBh5iCQtdnn+oinwxRASYnVuU8NUi8ag+kr6nprLL933xmGCaVO+UqnvHOwQyuMN+R
Durp5EZmbYJg6nmNW2O/b3oM6CgshNhHmp1u42lnDQph8S0F8M6xRNiV4Ng6UAua6uQxWteD0++A
ODi8IG9SRqlxwR0kLRecVXC4m7/s8xxOOioRDYfW2xBhJstBJwY+Nr7BW8nQN/QBvkylsMMXSrUO
px3lWkxwm5YergoOKqZn1D0CX+yk21R/v48EolYgMmnRCK02EmJnLxQ24g+rJ41RHVzESOY3HSMu
B+03UJovr82XYHr2/XO5wi7BOAi/q5HLmiSB/dVqeRcCX8pu8ju0sCEktKOotlQLbbxw15nFpS7P
JEe31wcBH6DUi7QU/IiWKLBf65G7Z0CAqebwzwZ0BMjs4x6+BxX4O2Ui/Bbf1F/Y1eBjZ/JRRbg+
WqIcj8OecogoyD4Ogzz1Yvl5AtuyWwTpJjogZQ73zJesHBSNhKwxn2tF0qPH3R2f6h554PrAUJBb
1vPJUIcPQajJMJ6+Q+JyQCdfFteNPoypIJJK/k3i1P9TIYrsRs2EcxEegDHqneK9O6fbJ2cpx1qm
V19r7b31YN/us3juiX2o9ohirtjZc05dyJNrQ4KuqH6OaEm+Hc75vUEfAFStk7hIEQkhtoofVDdN
3PTg3ma2KywFjcdQtNVqibrhLV1K4yPhluR0ElFFUfDQN/6nWsZlGxTGGwZr1WPfBmGQzgtN//h5
6Sr/ieYMI11y5VzfIALVrj+uSdqrYvpB3Nmb2EARNvHoLTexTmvlccSS42wdZFnXJubMBURBrG2V
r/MdULeqxSS2soLygWo54rGkcOJkTUxGvmLwjb/nUnS0A77nO7lcHUPnJso3SkQwLwB1NMmJMEUc
5Nc90xS77RqwdmJj4gM9JkbyzxA9+soefktXk3BeoR0yQbj2DRJSKAviKKSPob/ctlmnzMyUEzmp
w+MV5fP9POWu3AyZOSb2i2XUBd1O7+W3dAG9PxDlI7DqXrhwIUpyl8coLLOt36a4layedcjLVSjS
lTG9D0BKp34dnwjL2QWvmxhzPutscovYYwkytYxr0JmdO5phvfazu0BOJdlfnEpalqyJPIYe+J0o
CgJZhPZHZd5yRyClQkgRseGHEja51UQl1pR3puUYo7TruHhOavFu+vwyKf/mm2WLutmre1ZPUzKF
vIoaVyt8Lns0FEL/yNjkLYqLkIH8JmGpKgYIyPPHFiLQiVIk7byXLK1b2D2ZYdv4ZuMui4px63Kr
oBobny5XLhAc2VHokVvsA7iCd46BFenmapRGQB6aUUdzm6THF1ydFhN5QxJqRbKkv9kLk80K5FL/
S/jJe1o9tBDs+8cDbSQGQO3MPl3vxtYLM69Y270LcsNVE7YxkwakmYoJxbsVOn9O12vJWlRoLMOE
mnVZr0Fl2ZgrYtVHyIkW/r97SPhio1ThrIVkoE8dJu9YSWyvqXuZoP+xcNSmR11Z6vVwNPKWnO/M
rVEM8SSjd6Wqg/JS25wdkGUbH66kS8moqQABdXaMpbfG1fFjzsP9JkXOy811XXCP67GUGOhJ4d5M
EcvY68KhWRCbZ7KLqr6dYjLvVsq5mNgow+0n6BLKPHF7rz6YpbbsWAvBBp1xsK9nhJoSLBx8GoDM
FroECl6uTE2kv1p2U6BTHLrzagMXa9GpG0qq2YdFaGPXhNAi2s1OsFElq7AWM1g31SnPi+U7996K
xFRZIzdgWGQcYkVvBER0MH3AGmIaz7XD2Yre+hWy80MUMNhCqn4w5CTc80f0gwcd0mgvGbWADBC4
xh+Y46/78pQptekmI0aduEc2sF/4J6hKfrbTisfIes79+S4IAhTFC8kigj8m+WEJZSpHkrdtynlk
Ke09KspMsdUg1Ue19hTL809gwoo9uuEYA+YvJUD9LLadElNjZuxyLpufbSzvHBv5ya7tfpu7bGh4
YQhNlDibDScUkSqCML/MjXFqm520NJZvBobUwmUQ0OlJkjrPnQUJQ4KvuUE/wnqujRqXHfyoJnLP
aQFxHZNwx3X5VklCMo8iu6nQyriWyn2dRTeAj3wPySh61nMTfwq9GQ7byoKCwkgvWvihnPAtLsd+
KO9QjAWS61jApmctwZXnsA+WCR+vKcOyqEcuXpB6F9Q6LlfzBpPdH01YA2MeNCoi1hV7f0kdk3mX
hXFuRHGXbzvlHDbTEMxmCsqTHgdw2WvtvSpJQvnDiTIuqG+ubmjkJLPJGs6u55iGLpaaaNYw8bVK
hEDtifUC4XcjpMz+FM2ZAgQj+F54Kuwixv73wDiSNSHTOzT5QKBGMv+IAE5zQ9JfQUYl1dlS4/Hy
vXVkJK5N1iUBEDjN4wBaYy9duPvwF7OO3PVrD8Vt0/Ax3ZNhsM8dtzAOlrsJHt9mgrBS7DLk9Xko
ZoLLvLgx95iMLGzxivuBQHeU4PLf53L+Jx0NPWVFNdLHU9NxfzdADDeJ8/e2mlKpik65DeG4pFOV
/idOxEkf5wZ0fDA+HjRz2CdIekD0V4mUrNbPZ/F+f1oJwiQplvm6NidtKUwSkwWuHhy+TihIBu7W
Ljifh9udhbUv4z/dSlZ2fSixJMudYu2fescQf9D7+2Ccd4tpi7tYTbRme2D9ZNwcWL9bX84TOhaP
8tvfsBgglbi6dtgTMoYNv61dNQsrpP4PnSafMaurCRoj3nvYgaRMXJnJZyfZLnsXMazyHnzVnfuk
DQlEArdPea5b9+Z1IdSxc0FIlpTEUZ1dPr5VHwBiyKC258RgypiIW6ys106hsaSGaiS6ACTIY/vD
L1wzytoHs5iKsNX76b+Z4/jnkzjg9GnYcU3cm5jwtdVdxw+aUB694auw/AkSjgQ37ZF66vXGkBFB
K2S3oFuaNzOXRfKCurPKPkiQF/vJ5jYXdgOe06+JULmlRefswnRRytLT9xPP7ANXmkpMMIREokcv
cPuA7kFmM8IktQVt4s0O7r8jAGs9xJmY+IfAuXgTy7tCcoHFBoulOLmaVB3gPM3OJtc0dL+Ei98T
D6+4CpoCcnWUnXUuLkCnpDH1I0vohEAWDMK3Jr+4qwrXCPKGY9/ja2RBe4mXEec6z9oEnPaEUVhq
Z1qN6ftzK9fC1pZufy9sxpm0vneXpu6ZdjQ0ydko/8JPakQF4PJyp78RGlGmPVI3nAY3xi6Dx4U3
1DGU59xsaAatL1nd436lVYdEChCfiVx3T63TrIZQ9Q9L2yhFBQ2nGeRA2GMWXEDH4PIhakVA+0+z
p2cRNR8UqHGhU3dXqbt3WMYDKE69Jdy4QZRAHZlq+C2m9kxEoTrth+EzY7+NIJYFf2lVSr4qhdoh
nKvPN2QbK8/gxBv55Fs7bbvaCPYwETHJQXnkpN+dAvJ3ZoWXwqKxy1mi5WLh53Eebu9fkekrvllR
Rle0kFuU17k3tpO33lVO9dbkdclRBw4U2o5CCbW3xjG1mvkSHQ6RkAZDuYU1XCyOH78Ku2zY6cGK
X4zW1dFj2PSUURwjM9VtRfj4rA9+zKO1UVh3SlXi+G9Z5R7IWmBI9YFARXfGxOH7jzBpFKORl2DP
J9YJD7Ho2QOrNqTeHxGKxNZ4v8bwcJFjGjI5Ly3QEEgNPSJQYDLMYI0BAbCmbMlvxidqgwwKuSgr
1NwEUatcOLeKUxcVWne3zWJY0ZyXEIBBMz1BOOIaABfWZfyMxs/Qqc9My+xz3SsGxS6x+vZTwvB2
GulU+B6gl8PCMRS2wGCBlj3JTT7PrmccJtxOuu0JFinw0pH7LtgUe3OSuX9OLaiLsjer6ZbyF5uT
N1vl3AzJOead5iYWIzo9No0/o4G2UlyQY4yroDedxcyOeUHQlqT7h/akIWCBR2mrHf0/33yS5zi/
uH+h3NkJkjsrXCyi19DAqKsQCNTOP3AYsMtjkMRrKsUQbWVSXBweL94fJZY46btoXKhSlIbGiQ6G
FO2jVY6Ts9o/8gOOPiRKWt1ZVTK3FWXkDOKUjTmjIvQOE46fY7Qr2iC3maSNHHzq5pC1cTYD0sIY
9rOFHhvVBbrkfYlZ4hcdy99tCkioL39xouHoszOGGw6btEm8h8alI7HcblUyAoDj45l+B1tbwvnP
xSO2jl2ywq9bNylnSdWL0nRVvXTUbKNIjz+IFYDeknu6av+i89N08DVceJHmlWDWpLBGE//JFcz+
jhftgpWIfTNsTBIhEohLKFFpeyFKsta5WcVMXf7xi4jdR6iaRHTGRWqyqJZPNPmI81Hx2K4yxwzm
dnKMgc7+KG4geo7lsVfmLfEugbyIWNQV7LD+v1yvHt1HpuBJsPHn+BNXHUdZP0rQyEPYACxn5UPm
66OMOugzZMp9FPdcpZFmSZU6OL1gV2xvjXpUYQPECq+wLqbceBoQlk6vbVC04tDApEj6D3DcfTK4
P7pyyUE0owXsOKDyCnLXAWiEzh/MUeKn8Z2qB6JOCCQluRKa+dColtT8Vv4kBAml1GVtdRT8dyEh
ir820QTAs3G2qepXhP/Kt0gzMqkCFWo4yWlnh3AEH0G01cSnCrrf3Y2p+veHpqW3CKqnQcQmOl8W
SlvnDLU/wbhjN4Si8aVgj7GIBYc/y5I0w7DJXyUAkquPEDHIccJzG5IvBoNRiV6QWsAozc4aR/eM
bQeE7/hkuJY5qxtkZtS2vsxGCo1Q8hpCq2KHJvaSzIrUFcPBV2eF3BbLaVhUnYspWHg8kdu0C2cs
8faDZV8cKG7wrjZvheIkvqarbZOoiflip+S6YpswiWQGZtt4Deltwvk6KjmXfM02dpE+d/Bk0on3
hBflmPclH948pg91nRYdiN6tv9sWJtpiSaaLf2uKax1AUc3we+dfefMD3lKr05yBFFL0BV4Ih4Ly
at4Rhalut1CtnLtS7kh7xmA2/RR+O4LZy70hoHkLWz9EOuz1rnq9+/uN/hBctgDJuYmIJppQ+H1I
//ZGHtqBfE5b9W/9s27kKGKcHJyXwhQ0DMXDTCj/1fiuZxDP7SA/OSbYwj7hFD7Frfx0RSheMskx
2PEzZivZLRVW3RqhFSbF7mHSUKqCb0sjSb3BDcG3sKbXX5pKIm/Qsil+FW4fEZSOzj0+YQdPQH1x
bwUq5SEm0C0oyfV48ouLKLvV7sxoYLSGGdg3ZoqMpIcZudkfviln4mXpiYAplW123QQqnCOT5dze
HS10O/wnkcyUwn8XhJtEJkniOiIzC+GShIU4qYbLrQJMfom02zWEXZLu/mGrKt/J1EPEOkqPcM7H
j21kMyG4i+Fp9cVczy8qwPjuXOgxb5iTyo2M8cewLkIEFwFqTJvIaGXIORqhf++uyaNdVVhR12IU
Aby/LYUnI1yh5i5DXgf4uW7ONhNZWqe/A7RtLLFPDV/kyYqvQY3rc052q5cyhJXoEUCuoqqiPsCP
V2FuQ9r3Lunv9MTYulhSw2y5ILDv8WP4tEDQJCDpyezgS+vSQ20vpxTE9Viw5q42xEkzlznCdCdl
5Jvj8f341CbHri065VCYQHABPe9cX+Hf3VvgYsTSnHh0mzJ+bCZaZcyJFjfWCWmL0hGjsq1UouJY
k5LJI9mlxvpnM6vjt2bgc+IYQha6vXJLG6p//nIn+VuRuckbPQObOQdlXJTMOLhyVcoHC58IO+dA
0NRpTS5YUs2YJTPHTh9qswhM7+claIxc8U3fH1v5KY+kEVLzjNEfq3m5B8Qt+RRudcpbLo6RwiXo
R6MRV1Ibmmzf5iB8t1MOPJOz1UlSH9W63vaVfSKXLOPOG+Jn9Q58crFPCNdnLO67GmttGY51ug6m
IkIg2MQQQ3LiDp16XmEBbQEz8TZT3DajJAahHiiD1APmK2N6yXs3+OMuKRcnieycGutoE5wJQe0B
J/xxygburR1gsul3EQoiHSltZOXRuU9TATU1qcSpQwPoMvBS6/4brA/uJMhuWIjwnCCsI4KLZ3uI
M+IftML8ArmMZwKMqZEgk02fTpNhjkRKA5o8TEmXDG6f5VAEYWliHb+B5wUgoVevjWj4/CGm+OcS
EQTFMWhG2M0C1EqLTqu7YSgbzyDB2StKIMNo/uDSwc9c3DcNq0PUhNNSetldvqsVbEz1fDJ7G35D
zcjww/DPyCKUhErq/0TSB+C+c9ffXPB5d/5oNU0OS8jMeDOQVg8Eq30vHZZtsYuFgF9+Ca+uqCHs
gUUsvO7VWPkmjOAr9SG45+Yl1Fy7wh+6R5mbxj6ifNrZaOrVqJ9Zuxk8f4S71WTIhelsoJ976fq/
ZRHni50zBtdSFN6U2EiFK4d14PAmyJJqCs5rQjMylz1VvPjUqchD5AOibbezBShMQPgEHKJxX2nw
yVt/BU3SIxno67qCFAAQaIPwwNl4zjM0+Ruo8O/q/sbWeRv7+rZKsXgRp+Hje18LU1I9x9Pr6qt6
+WiwzcDhKWe6XIfIWDmg/7Ie8fbXuFsbzsj/teh0dvf8jAl9M52vifXTPgq5yLsCbVjlAv8Lvw0z
qcGud158rXbLDZJnX1bAaPrEHTEaybi+bru9nTHMfJNitiDfG06IWgZNlh6rAChJEYaIw9T7sG/l
zwId0g+zpg1Tu2vE9JLGE+LrQz2FuI5YpuPEq17DFptWnpT1072zXbgfWFF1S8szuQyQRmPKeCLs
kCCblbQYGi3rGt9uBhHXN47EKXVowDxN/Ut1zf+PxMosxBYbYL/Rnfccw1nlZQ3op6i5BEAACEt9
uPnKWFEzfq5AnyhU3rT0ESZP0qnJT613ALlxE6JqJ9WgCYeqCdnqfLgkCFCejz40ZYw8ezQ+qFTm
0+HYqgX/Zr0aSLjIiK4gLcGWthVqhmB4kt07WJcfOdc81IKoTcYG8z02mInrGZMYUtL5z3gQ1d46
AZteb7W7Y1rikfeI3xGsAtyX7nSUIJDfOsIbb7h1wTSCfosVqAf/GEdT4cG/B2jGFl8JipMFYGub
H0fhhVnGxRKWbB9CQ9QdZSFAPVo4bPY2OSqC18/HUve+jdUJqJqUwEM8ZlT1xvXIeWloOwHJAEun
VttG1Ss2i6OUrQrNB31nSw0P4bndfFGbZumqoQgDr/dpteJx60GV/OfcnRx4eHTSdJBLfV/TdWIk
1G30W3DLeGJ4XppA/WVTO40W2PADy9Fs8ObAvK4CwjqNOOtyYnWsppZKZKm/Qhh+mLElwf3hmY+G
fq2PchETgPObdNpBW/D6EnFF6+gJsAaeUxaVcwmS8bpjao3tYfU7ra+EDaCNk2E5qBY2KP8Omx6W
3cSM91Pb5UxiBORMAwiw3/TTu8K8/C/MsvGAg4if+/k4Rv1xh0pX2Fiiw2VKwfUStWvccJkAnEwW
ZymqGVEaPwzVmxBb2DFDqGCUGQmekdWtgFFxmwHsRYTE9QQ+pt8bymjRX6WrllHBAQyonmASD/IL
D1sl22+tuGYPHZ2iT+ryWwMpHAq5e9DLhC5SpX59nojNSsFexpTGQ9m+x2sIyxFYWFHomONyskDO
bhpklo9yEMY3oqzwQ6tPi+P9IVJa1SakyhhoPsLdXZMzQexItjhvOm2eAnb0rIJcIUjo62rPl8Sz
iwfJhQdN1viBR/xXQhU/hMo7+6h5e6WM+w0mrsH7dIFquPUiwn0v2q9j1rYalKmnZAItHAu157TA
26u/XnnX5d/eCwC+zqZzhSmHVnkQ+S6ecyY92RjNUrS3ifLpHNFaDr9M0Y797RDqw7oPhu0E171K
Cuvo209hjyy6hdnbCNWlx5BoDmiL2PUeIe3SfWzGMzEO/Acz28+YngBNovbq3Y39IMsgkireaZEQ
a3H+vuevrna4ztuU2Ni4GDGm189GHDEWKwE8chebmpe4ZurEjpOq1lbzLtNiR72kNYtRwLeCoPS7
RP5fHxdHzJx0nawqeh6knekKNU+WuoVQWRT5SvFNWMrYDnH7F7fTALtWT6ntZBxY1Y2jcjqM2xNG
EUDnkKBTAMnYQmqNPtzbPCsf0x2bObjmcog5lIagPSx0skGxrVop5g7sTWsonYszi9cpD1JSb3LC
MOSC7PhxNd56o6BPJpxCy1VDGKNJYXR3xkKSpWbs9dnaGAdftSqHzBKltgC2yYpgsUPscJmCvt4b
Lh/lWlvnvd8wHvxMZjTMB3kx2IIKjfGHDPdZcqHjDMKn07tZvV1e0HHmk0PoUi4Ab1Yc5C3Nnw6J
h3qtS7YxBduIJvGOyzVLURmYdIk7kCWZrk52EwaL0MmFYg9A5OsvPVWpkvpMSX6Dl5+q5vLAvLuk
Tf/NDTdmGwybKGDSnvIl+yzADVadBu8GCHc+lp6HEL/sdCTlEB8PgDPSzinfLTSmndP3qCCrZL7a
hvzDrvqB3bh1QyAhQXvhKFiLEmmns8mUpGGUIDYPJj8xQ1ZO8ss/VdmB2Vvddem2SoVKIkzWg++p
VYmMQcg1KvEleFcUIlkoAeBF+Fy5EnsWkoPx8OK8Kt9qncmF5GSYu2sybRxpCV6rlogsZioXHXZ/
F1IttH4pq4/aDs1hcVJHsRKv/mXkeo/Hp+Me463A0VlTf+ap3+JUSS8CzZXP/d+UlDmD91qxqgLw
oUcm/V4UAd0lZCd7mg7RwKr28FZ80cg/RtK/1b4Z2xKqHMa5CUx2BAbtci7PqxuVZn3htQopC98C
Zrxrt+7KQ6OtVOIv7Zr6DzLRtPGoXeToDHsJgHdz5QaqeucwcjG4qXT0pzHAx65uCLW5nFWh0JrZ
y/pNCRVio+MUX1xsABQGvR+pNPnEVluLnOTLOpJiqfXuTTMoht1zX2/gFx4Dsm4b8qr8xktDyApl
Ire44GBHrrEHEJznyU6qTa7+jp94CuUK7bTsFKXbO0P5JFbjNw0EdkajdsndKOjJ3/8Pmt7eBiK8
/Zj6l8FQ6Jt6fU2Wtwtb8CbG3jNt41Z6TW0bHbwiuj+vsDDmRktI4APJs7xdNWrCmjy/py/Y94+V
UueraWZD9FZxSzBHQPONN1ds0zeZWXgLb3pR8EaAFD0Ebof3hYOWIg/AzFMtZyCCBB5woxULjPjn
eabjX2P1ECL4nvsKPa9fAkYvpClIBBp3vMScNgMw+g+Wc6pEcfitPPBu3ydD7GhfNa1JHKy/JP1C
Dfrjp6zfk7n4GLO5XsCMpO9vIlWfIVbn5iwjBJJLaycLnad5TQTLEoEP6QFTgNjLuZYf02CjqG43
VqeI63uUGjX8UUDlLAWHVZl8Q2XerVpF8G5Ibnpxu8AxNxhfDmRqynMKoKJS/uWyZ8+0REYHBej1
ArfztxjDfo/j7ba4sGMrTx0dwwKGxy/b86dVkS2iUviWCBjrpk7bTZAqAuzw/RSI/Og0JZ3j8+di
OWEiulRcIaI7YQxiNj7cVAtKOKh7uxeEUekSb/4F90RgYEPq+32t1roomJitlXE6fqqAinSj8E1h
Ym3xnOSfx9Uv7qYkmyDzalVmEfXzliEDbcZWomV2Q7ZlqUK4lRoMNSICBKT0ympfALweeq1JMFBZ
uft2iBjZ2M20XoVNwbjYJ40e6FjG5xjbDhl7tXzEIn6lZZP5yjMGwsVr8HPvxraVnmL+y/XddmJK
45wLTPQjnZZcWnE+ALGZhwB/bTKqumcPaRso6WS/xze5rs8jqt77b4s5bZ67QYfwzB3omrnQCEGr
4y8d3NnFXH8Pe+4V6sDmQ8QO0KePRa5Dy65s5tsxjKmxKWVi5U/aTTuuJarR10gxobdojwQV9IqN
uYpgMKmXgC70JSGjZrBa6eO5UIcrvhf3uxvEqJ5Zq27Ot3/Ph28c1bxcq1o+e5BJwOtZ/sjDxbr9
GlujVTl62Vzc85lmXj/IQUjzRyHVvC6l21qcdii2pikrWb5nZWcXaLtx8HmWg9sQKDqTiY1XnjI7
SVmKNTh8/Pe96f21r4GIPNy+K+A4MfopfK9g39cH0JdyfVqtMflfadfsHV/tiG8NG587ttyDMhfW
8VBpNZqGe78qLHaFoAJl+RtitVC/A3Ra7WOx1GVkSBqeg7gCVaP2qenTlUpVmcdks79f9CrjJdz+
BPGKgge7QiN9FimsI9U8GMkaoBmpAgP92appj9uACYxMmqpvxMaKxf1rd7/+M9DhdZRObdsrB965
XwEzFb71AsJQTdTmLiYJx4h8ifYMZHLgUVF85ZJW+L8TZXWorXXqtkfUvA+11RdguwfFLzszMOdZ
2pJDKh2etp6LeFx52NZ0ONvL0+WR04VkczMYsJaGVLk+ABv92W8uw2/OhSUCMH/G1RcA1ygHy5q5
zlVWI3d/Ncrud+8jRMLj1u2npzB0uEn7sI24U8oRi+e4PiI0lKoNHNcRWot01/4mGaffa0P86TCI
m7osWwbsf0gdnZMSo7rrJ84voI0lQFbvsG+km0YhR/8A4X9jTZ4Q4+Edc0THJfam/coBKcZuPYfR
1vricthPEgibRW2KlIIoENZlGdDH5GICgzUGvaJPiFi2A6tQdQ61J3ALCOjnEe4+v0d6WHPRp6fC
SjCsW385S0wLREiP95iDe5NFnW7CGmDM3NzRH2ImwxdoyY1cd7qeCoSZJhhPL23Leo5P1xDDQvkU
wBIfTUY5lArTFXUSGp1xQZjmR7K+2cGjft4h2wL+AiSfJukS2kyZd2xHrfXPmPqxc4hXglhZLL8S
rQbXspZjNfgJOPnujGaYlZcNGuoKN6cUyrMvnAj4RZsvMXcKaR2M0VUm8vlKpt8rjcHCiOmS08dz
MzDXM5PYn5HouVrhRFtK1Ug/yQmFO0ueIXfePNvfJJazqjlSXaHLCSjZnTE7eonVZY1hw+DUB5+J
Zbe8n3iwuTv67KTWS2h42BCsMZlQi4Tm311F69ifOHHS8jGNhCSeIPFO1/uexDxU2kjUad3CjsWY
OLQD0rm7IRZtloCcSbwEEKRFkl+ETFLIghUfoZonKlw7/re7nmTMfPeMPOwjdAPHDOCpuny0tOfM
6MoJ4BsWdl9NtYtAN3+pY8U3rfHkIE0war0B25efpSKuCG6R5CWbu+qhIIBy5HXkARNeyjuCiKxv
IKIkbKh63AZdQL32+C1VT2EjRT26izJrs86dRpK/Pbz88Abp2LlfNEw5lvJVmkuNtRy7u6yHdby4
v7Im6B8VH8bKunSsf/nV89glE2WIzIpUy8br/iLYX+SdoO7BpHw9B4SY2Sht05XPR2trGUi32xQh
818o0NcqUvlfYOT9cBJSOy8te1hPYX6NuoReVaGoa7NRCKGcqTUY4Tmz8GHJbgDU1clpX9/GZ3q7
/qu6FjaPet3hkDfIsm8nctN1Kf3JBMnR7GDSIt9TQq6t04Dcjrx1d96GcteSXK394zZsVlgXGekw
GOACdKL/jTxlMU+hTKyztq8yTFELzVWYyWszgUcKmyA+z8r7tjag7mfHIpbhvvV9fcQkuSXDxd9o
6SStJ8vxUheRYRVH7BTAKOxN16qGr5jPP+KUsDbUY4R4A49kPh+gUkxaQ9Umwzdq765PiE3RwPZS
WbFO97kRSPzC0ZBogNQ1PU69a1P7FMhfmXTiK5Up4Iwbw+FTD5ouGLZH20GgzNd+BirOvsesChdv
ElrU/XCTrr82iEPJUFVwvSOkw3klQks70nAlQFpekR8e+8aNvOztcGEpWdJEtbN7iLjTNWc8Jsja
xT2DINnRCfDaEGqT/KQ36wJnyYjwP8MZr5Y8h6Wj+8PM4xDmLl2Apw/CTWeF0N1TQmLfq/gOL8x+
FOvCZv/b1xn3TpaBT9U3pK96smc7cVXqyrMuPIY9FfTMSOe9OuXaUB+aYB9ii5uorR7yowFYOuRa
zuXNannv5iBA+9buY1W6C/Vv32UgFw0+Ffz/kc3+uLZbBDWfkIpmBANEFuk3i7guqodXY1WMyzhU
xDR/xX+v96JwuI9R6b2kgV5UZtIuHqu5W4ylEt1bh4jZFQ422ET5nkH4EP4hf2EBABaQt4Dtp2L0
1Ujjs7VkyOK23owOJAMr90qnEUG/JFKN/sGv4l4pAYXGsEjtqvFt60bliCoNju9Vfv8AzlNJAO3i
LDVHdh9JRUEhPwx1s7ENm2EyRmP4QGGh/qeFWyNTlla8LphX6j0CortUyonTdjTOj5bBao3h3gVP
qZjok8aEA7RkSUICKPvEa4nN3WF6pc/q3dZ4wAqZF7XG/CwiMBBlcNGvZQ1+EAv7FLECNguM2ZAG
vdUvM2Bqkk3BA7m38AFtO9rROlhjwZEv5bctOHrdFM6OU9O9FO2RVtvDcuehF5ie9vSxHL/h8nMe
PXCMhmYZ1PRFqZ8PVqPk3kKmd5u7o9vkse5ai7ZuCTu8VI3vIHEBBjXNLdQD/nvjU7f92rwCV6/Q
78d1hh8teiaADe/evU/82BWDxN6klS4EqzrcrNl6KO0NiEfbupAF8Dt6OWhyal23tjtqlJnpGhkx
LCP8b/6pntR2p5gSp6wk6YS262Sk/AOsNL5zS7uyN9Wuqj23YFGOdbHfuW8BbSu7hQ53CcoiOSMq
CWsLpeR/fMPwRJe/dDrwKrF2iY1S3hIlJv/x6HnLPvQGGKphbZYJ2uN9za2qAMELAQLUy/rGokzk
ZpVAXRHgcvZBOsqVYRx55jOQhCHCEnRcSa5BxTJbri5xcDVdqhx10POp4NK4s2nq8G/ANdu12Qbb
06MwVSe5zRiG993ubooXtGpJmU+d7zHgh5iaFvfFqArYKwO/pJNnsnJAKlURLuvvA+A2eOg4zSfZ
DkawJlJgYfAj7C5Oyi9dPBOd+e8+esdUIrZldsefzYTPiqxUSptXT3crTjrkbkoi/x73GnCsh080
kGpbR8MOHUHzSPpROf/73PLzBNPVi7iW48v5atK0mUBOWMfGvfLjmwYU5I/eVc31cVU+GXEkzzK0
t6+v/+eW+opW/eEzmCii7ju1kAEwQ/OTky3gBZhgEdR4ulNL3iq4SyqMJbLojzU0l6QifpXGjF/5
eqLsyT5bLRkdFBZX69ZzwW/qd3ZvoPGg+F/dk5pXcwfwZIEygfzE20H7N4fjzXhuBzjiTV+RGL8x
r5G5QX8s1ll1zpwxHuV1x+PFrk8xHsQZzpi+oerkmHktfvwVz9XEe1zfOjK2sk7ViyAxci3Ebx/K
seiZYFHHy4EsDGJpGfpl0aeedvw4GaX2lEuqq7lZ4Wrmw3DnGsuzC1XI6xX1xxMS22/eRXiGMj7j
xb6kEWID9oBFh6jwQIAb2tzZk4vUpXh/oJvmEU3nxL+ofh6xfaBwYYR+ZMzzfLrRQ90rqDI52cc3
ZyZe8AF8WoEZX0qu56ERgX0CQVylFcw4IYklJbMBs+y1KkoAiGdrN2fujzb+hXrGB5zmONuq31id
JkXIdidQkx/Zr1CSx8Q55dfqwOBDFljbN8jEH//JVEIRsovfFYC9nQNJqXL98U482yhT4B+Q1AFb
RxKtpY7VFe+qqMIZClbD8vckOZVcBJwn4XoDkQSu7w0uOXJHYlnHCECsaK39PU/z/+N108kBMyWG
5ljVZIlu6pA64uOqqN7zIgpd/rXvWElhGNFWoIB7XUuTgxIrTTC7RlUSwGOyW5KbjLT+e+7jt2ng
EylglVSRxNxceS54HrMtO6OgLdlwFRQNsgUFLo4v4QPfCvnupMF6OJ0o6wpT4V/WQo64tqXfA9mZ
vhtqPzEFM4std3qtXP/sr8EB/HuV9zT404KCGf9JPKG+VnNL9zOKCI75Y2UG6cI1ZGZDT9GxAxmF
zWcHp7Ng1XAhvqVB3V5cEd+oQiM8YDrWlhfojgoXH2SWum94KQvc7yy0wWCxrsBDKg0Jqy26M+5v
MEtb0dLjan8NMJ1lSZLBmhWTi0rhzMcFmQlqY0xXhMsrh5Phic3LATtJSpytD9/gwauSFoZLeL/o
i+lbJXw8YQ1U8iKYKZNl0c3B3sl4BRx63+6wVq0p46FHBJFV+WpC6MrDsbfISL8N6Z5izHX84BMc
gKN0BxLorQ7OlN1dXvtm8jVGZndZ0ij6GT3kf9Yb452Ri3GtJvWfWM14e+UTz89hAohXa2FVxjLK
uy8j+yXEw74dl88tnsvgjjYafpP6vUwgRVm1/T74UppKnmZ/2YFwedcWmRsBuQ7YBXxLu2G5lh/G
VvlEp2uWoHarn8m52nCi04SDZiq1Zpthblw3DwPvrYhy401Kmsq3VsgUC/mOVep5u7CMRzHCSihN
MX6faOEFpnoBOC9rymKpz9j3oDJorECwcAwvPNqrX/jmyPUBCOeOLom3OxyLH778y6a+OOQ4eLx3
BuOnC6YeMcHNWYmfCKHjWCEg7rN0atVIT9oZOyqJZv9z1ekBp1Y+cqg6CtckqUNIEdP7GSvTzSOp
G+AHG7oyzF6BWA3iimHT37i7HiAiFHkvllYxjd8hxkyfg6wcgxcwEaYq2RSnAplK+pcoqO84q2a2
K+mrhflO5PhuppLs0f9q0c6Yb4lA7k55cUWi1VXNl2zVVxfHlcN1U/6djy5Z8MTSTrbHD7vxfpid
pCyFuqMbCRpe9zteNF/sZTzJKa3gp5VQlLau4auVFgz36xkFhunjHuxKGsMeP9A92GcQB5MJTY3A
1t42WMYNHw+q/66TU8x5LrElR4vXoX6CJTpltufgJ4Kw14KGVwQcjSxHlnjrucKvgFWnTZksiL6o
GoNDQBwunLCll5Tz7/wVeTsiVBwStrxQHSXoh1uRLZcocei/xfGbxAIOunU+yjZv3q/SfDIJuhq7
tF4Of/TQAHjJylr+n2bjNnoLzX5Vc0aul4fq8V8Xd5PsRQoUXT813dnnt2ePb8DPALvOz4E1omQz
YHhE/KjbBYkWcA54+gBLK3Kl/W3ykmbQFFrD8mGYGJD9qvmhRC3rCCoO1Rr4QSFPWz10s4LG7sCx
Xav3Wteiw9Msf89qeLz+p+2v00DYZ4Ir05+HaWDAp3mCsUgAgq9lmXtTiG962iVtwK5vPPutSVF2
7Ch8Q51owdyfKXVQM9szLN38OINa4Wdrj/nHf86sU5Xi+gwfVRGmLOzUgwrCTGzTJIFcyRlkXbJu
1Qzv9azRpo2nJoBnmRv9SQJI0d/yQ/a4aUYfnvDhBj1xS/8ot6TDXs0VFoW7d1XTDRZx1jxIQf30
DPlBvSqLwcaD+a8a0AIkvBk6c6X3enWh9xaKSgCJbILSpLtLXG2pF6MweHhmC1hhhHgOSm6+WYsF
+glF6CtZTQgspin6FAOBQUVjGqvWjif0EeEtRhjn979tm89j3duyeMIqvQEca5FSSnaPKkluDG4k
TVeRLkBPDwbL+SrEoQ/SzeFVP6lkjIjP8vqSwwqw9KU30MEc46YNfVDam5djXFXqIHwt1iCxYTjA
vMKYDZ0H38/J7+js3OsX+DMgAo18MkJkIDBHq5DwYNjqalVwMI2xLfMtslnJ9R1hzul3WDizB+5u
3sCK9DA4h0PCNgjuYbEvTNQ2IgwF7a2ixXGc1HUajCZZa3fyjxC9oOQrTb6I6CwYeDlohubX6Gch
yJPi3h4CxF6LygnzRJ5iJNeLWwkKtB8mFLvhCQfcGBIadYe49biJOeTQUBxT8YGdBjgp7Qn2T60E
c/X5Tc9DjoQUQ2/tXw7h9AnQLyOlu+Hb/zGaw3OBfEslRc/y7NQHRueEF5QSB/v7VMtV2r76WxG0
prrINV8sGk1p8fDqrqQVD1G6PSasCCcUL2Uj34M7zL5PvPIm2quuPhSbzvCFgYPhYAvyqLswHUN2
MqiMrfGdsO2iayzyEejFdfZkm+NBZhM/VgBejQ9AmUzSFVIcgAg1XYLkuXhLSOpt7ZPid7X++Smf
QXSkFXY/8WBA0imoRPa4ocDrNsyRjp4/rneuNTfNui8BYJtpGydzrQdnh602TdD6OOObkWWlJPBi
+ogpcz0OKdRIFzH2Nst1g1uq+kzHbzdB5KUt6dAwjr3mmGoV6GkBM72YBVYrPeXHOOVV9i58d2Pl
oOPGlEnYudrQDW8y9iXDjvoOLgeP8pKptGec+MskAiIjmgq0taHMjhP8dBv24WMQsTq7z9Ng7g4x
F2a0tEMMRVd76XfDHUWqa9gV0xHvKHEMNa/sf+zXxIdwjn2npf8P5AhBtFBQabz//IsJkZh+wgj8
mxDCNlbFk248wspk4FcTLGEn9nsMksrOf3gdztxoX8m4hQzMJLBtzheGjaLNRgYDvnJW2z47TC2Z
0i3GwoxlBoOhcI5mGGcpEYEvMn+W5UmqFwuWBjfWw0h0O3g3L+eyVd1/dpPGKg+dgAibt3FyaQdQ
11HOPVbPII4WPJ4MmLpFUWTEg35SZRUb7Asnzl/3NtWYygTqXacYxMqlrFN11SaslKS1+j1hdYuL
lKuoTOaKLQIc7RI58AHM99CYCLzjaHn5neXkkX73CHz0a2s4OZvwmIKxE1KdJ2Y8Z2urjTRadpjb
AUTUFIrAZXRKAiIZ4XQlU99wFf7KbQe2p6MKy9nqD6vT07xsnPfiSYKBwOBKZPTEYOncUkNJmPIT
a1oFaVfOhPQ2s07Q5aj+cjcw0LorBayk12LglNp9RVK6AvnuwnuEjAvsfK8LWbV6os5XOYEbZyTg
YlW8b6rH3hs2GQsESSUq2karl/dLM91n0+3O/EqH2q5h8gnbYxM+E9n9mFR3MhE+qpaSL53xYS5i
/vsJNg5nKGyD8Dp9IsjIEq49E2rWnjN/hTC0F0vi1PVaDXwAcUAtrI/qIZ4FYP5jbTKrubUDeoT7
JhzHC5Q57WY0ODTvFxJ3M3XvVhUjGTH6UHnUwG19OVQLPS6nCz57ubyav6sjs7/bYWdct4gnS42B
QbY2lMjsLC+QN21d33otQ0hkDdsNXB0m6wbHPqkzUwMCv1AGcuH8z1xO2T4Db2eVT8yWgBegBvAG
Sm2XaNkqmxWKOZcaRO2LWfK8A8yxl+QeklM04sacOAUdfpEId6qjgHMoPtykXjtlBudblVDY4pGm
Gw5ynqA+l5F59tAwA5xLPknhHCxw6xqQwj4izk7pABgq8tS9JVuqUsKdKNsLHMArQWX5OhRxEyG5
HC2Jml6aMrFvkXi2U8t+XY3V9xeee2p943BjxsJlWI0NQTPlbQwnama5Ao4GwzzklS/83aLBSdDr
BtVLcihanusrJ4D9sR2G3W9n09b2QUEj9VOb03sOtM/7Bhwe1vJN8DeDRDHgsQm0y+Ean0XhABxY
oCHQHIinBwjWoZ+7y3AjDr64XRH1dVaTUpmLP6IxtEI+RjSh0aHGHpE8r3mYxy/bXKwt/nCgthWi
cMqvIGJzXih7tJ6o96PiioKatczoZC/XV0fj10gsC+UrMyr8Iw7BPWCyiOgfJdwlVAysPlIYUFeR
5EwCzt/zJqmMc7sVWtublgauvTkYMO0P1zMkbpkWeh7dRoVvewyB7YmYrJ/SaKC2H7MM3nDpFhSP
xfDwS5vSDCBGrzWlmIfFto/uHQ0+NICfIfHBA1otZEbluQVdrxzmDiIYHpKR4TJQYFjboCqgu4U4
m9BkN+Gy286SUR3G0z+kokW4QPy26U+0hHCzDznpd+6G0ja7rqhKtq1+Co38POerC+STbaoY5A+i
hr3dbfGDE0TVT9kF0KUy9uvbUsHhyNYb4WJdzhaKR9+xHSgS09eg62vwg6GmtUaJVr8JURDFUVGF
c5BFkBBrJYugXHIPiiKed8Ozwj0+Qj+YRvA/jnQPqOCoR3GcM6vfeuN3jz4DKyHeuA7+PwJt/szQ
PNLJdMrc7Hyq8ybMy5dZylKTQrQS9Zongr877MIDy5e2q8z2vqO6fq4olC01lDk+71GkqO8DRu0w
FeUxOo7g0sOf2rDzoEzHWi1F6mTI++11JwSfEaUEFXDG+3H3GHK/SiKGUmMxWnX+NjJERUFkiBXr
JZbRffOuYavYxE3RFfxz/ririRuD3vgTkRq32vEn5A1579AAvMY2kX7XhjTCWpc5WIDsiED0Sx/e
TJIA/PRmEYsebwxMGsL+X6Xz9H5O7nWbF8BiEvb3kSBH0J3csf0E4fytUd2t8XHhqq/8ys9BM+sT
0CSJlZttoGerCUwbiDHuDGqapX6TSNf8P7/pNP5DaRQ/uiMzMQfdrq75SnsuiHownYiK14pcJZw6
RNInpP4V/qNWN/azw+nB2R49tfv0GvXlCi0QyCnCNgG6aj85J+fGCbubYS4+ToPd0FNWFMXoURLs
FJiOhNJ8cLPjR8cLgylzHgJvZMIC1rLmSwpAL7Gpg4hduHcGuveL1K5Y3RBKld1k1PU0C3SnW0cI
O4ZHDn4CHmFODsw6ad+ic4SGXrb+FHBCjKdlWPJukIFRnNPSd8UstnRwqddUlspBii+59X96sPUi
xNl8f0pFhHO6SsvjPmy6mZuozRya+GNha4lMFpPni45fNCz6xyq7MSUl6IPDLNIdNxV/gxfZL1zu
HpeJMdJkuzlR/xRyi+0B2kO96xuQfYZl5TjVXqa5TJpNsffpgPpF20dmPKGdyVuKGaZh70nlEoee
q0FjO2mtxhtBsyxjtdFOuxrr5C8kOqaNHMLlyBw2Fsj8H8deomwcuGYdGB3xTHrc0/REjFobLd7P
NJzs+91Xaanunv+7S/80FeIwi7ZeWx8TfbwvRPy91cdhJl3Ytdx50j3xPPXCg1Y2pHFLIyKdnxPR
93ir9tnUTIKdntcC28uVziSnjAJWfeK7uorDsO/5ZYAgvS8Qh+tteD07rFzjGNvpptiV725Zu4J/
leVC3Wprc9+YU1N8coUfgdEv/fr6v+zvYWuxvt82/nFN2AZjSeUSbRnItXSQQTtBiHGYCvUys6HV
yVelPBVOBM16w4HukAtV+soPzGdIIbw9UyROaxzFIomA5pUAjNkUk+9/0qb33htDAWSNfAnfhFnq
hWHs90q4Wmzu7bZqWhJ8QHXyJefOI8nfosYb+npG+awrxzQFJDLfPSVagoX5Ghsu0+E8nj9XWl/S
JZI54b0L61GSEkZ3VoXVp3x7rRr0NnVEgbAFHJadwI5a4VuP6wTc9gJl67FNsPCzOO5WvFMEte7n
y/oCvf/B3pedz0TaQrwi5sby6BM8rNiVbdYxNRFPHozNJ+LOkUSqUP1CCbqSh22/4zS6KBeFafLx
0Ep4wV/w+3yxXejV9Bf4wE3fWsx/UeV1sqRKXVBW4orVPmtmpfCKJdZMxARLk7as2c+C/8WRwAFw
ks0OhZk0tWf7nr9i+GSTBUMAdC7zZQCOVPbl0NCbgDBrjQuQSURNBbrUqK/fTxForG84bzear52S
ALisOxC35Pc2HpDE5I6oSeOoZmKKKSRqK3/L5YEtMHH871/5Mei6I/a50nlEp+00t0WOr5alUfsN
t/DYkeTBy2+0mR/CKSRkl4hoJeoeezm0Kjy/hVN9A7AqGSTU3ufs3xbRHAtIQUEhuE9NVzJ7dVtl
bC9afTDAiUPJlAtLBKeHLyDFDVnuNhnKVxCt1wIQZw3azg1D97iXENnP78bN5WZqFIp+7jUMv0fQ
upDNL6XWTMEz2LJaTjNEIBiPF23Sspn9MTPPUayuDz/YyzpJqLK5A9VWX8721bEHdUe1ort70SEW
KXEpt8VooNy0vx87nd0xCjwdGFsiwOjFXXHQ1lvCNVczrVDL4HeYUexvpHq7ne7mvlGqM8TryVTe
Eo6AnuaR0aN5VXcgnh27PHrF3r+sk1pbr9S5u1oL76UWlHdhcaL1m2fSqghRcFQnzd3DVgu1yDZM
0SJDZhDu/jXBx29ReIV16f4u5hOrjpyY4U4sJvcZahzEzAE/rar5r1HL73/SuwNX4rEi82O4NTOc
jhdksFjZUQUfx5Yy5gaUol4y3FbWOjhXLwOSBB2OX1D4QNOObPpSHDTfBH8lUH6h5TwPEYkmUzxm
KvpK+A9Abrl2kIK/qbQ4xpjJ4k9wtEPrGgKY1uYiGSwT5LKIa47BQY8dZTB90l1QBYJ9obbg0K/J
3NeU6q9v+/cJUIlNx83Czt381knMM6C9sO1vVIVFj+FLIWNHWsNp9PsieheCa/3t0PCvF6P0vPmp
4BjBkNUo3ifQlKGkyoUBZdZSwt3UFN8t51eNmpI6lsac08RQmkJ7gIehAmh3r7Cgn0Febg1W7AYg
+JZskHHrfYOmLI6kcKZm82OCLzuhEnnOQo9qDi2vmvHgenbcKkGSfXQ+pJ3EudFxXm9g4O3D1Ik9
W75VZzZN/F/Dv5OBGdkhjYa7V2LFVn8zC+xOJhUj2FM9tzqY2J6KvPAjMQqpO5MngLnhMCkifswa
Mfh2iAfMif7q/+90OAIDVtc2SnPU9YmtFbRQZDwitgtftRxG2PoeoPPuvJ8JobKDQCt0rSHnrH2A
Lh9LnOg84ro3xaODb1Hdi00+5z+4g2zbdJzaKEAwUJ2acIQoLgg6/SYJJJC68TmtqFQY5gHrUHgl
KMs6lWC4cHpB7GCAAXhTKIu/wUuNDyXQerMnYrL7h6AGez5ng1Fw5JFGqta8YUmV90NMQDZqeoea
A3+OK8+kELm72GwUVTpza8goZrUClFTxGMjZyhhQz0mXj5opmo7E1bVE8feXRIKKELBGHbVOHCD5
GHbdYxe38Bm+7tyJ8E9C6nirFE89PXsfWXNFULDoDDFqlS/4b9XH+apJc78jxAGxvzXHiloM0AIq
Xk5Yr8wbCWfrGnH1uWGf3xVEh44Qbn6XV/IG2sQIy9i0LYrxGub7iWHdxbsPqAy6AogCwxUOxVeT
4EJ+UKPuOniOxd6o0oAdgVLDf5xCMW1A+/7PDx96RZ1efQwVOLk/CAkwjD8G/aa6WA4ALDYsfkXs
4P5eEC+caqWktlOrmgUTuxtaKyceBohds5+o3NVZNCnHnXps0Pqbm8W/9bN0pyZRO/nbxtPXbMQV
U7BlMMLPuvWss4KjtBnkHTiS2SD3UEd4P/DPVj9jO+oOovKwzuFgJui8tJ+Bz9ot7a1OQUslV/3/
QTKXmWPl6oFZfGDOf7VEXcvaWLjQYa3ergppY2mCCTGryNLzrzkr1qQkuG5UYAiCX1/tViqRTKvm
WsGlhtCfPlDzsBkCGzFXz6U4MgHmWnz37oeS4y5l2pDI3ufcsESEg622RBXfipepAX2etV5WITdt
xYTM9UOprhkGe7TEAgH1siSnBwifgejMUqACDkawr9t0kYlHpD+4PfgZnNSyI430679eFGamRHLA
gmG2WwCVhc6Df0cn2Gpb/lqwKuUwhPWjUwzvhuNIFwsvagJHtcK3E+WSH5mRLNzQwwa+nEcEzJIQ
Apzkff8I1erBw/CbJzX9/odmWCVrrN+Da+OpsQfQXGHCXwI7eibvBe8AXciGLsakQ5t36jt09SQG
xkFkJORsXnZ6JnaXAkejmcl4vJEdxFZQZWNMyju7CNNl9wRPxSu5Ej5+ur8xU5yvqWZGNt+iR2bl
v+maOe2bJhjddBMUSLQWqaXUdw/N/y98pSNJYMCxAozapuFxmnkxKvWddYfmsRdHnSKym97QjY+D
T/JeJ2CZY1oq17ynhXIfUoctgFvn6DOExkBwY6RxgYOuLckUH7e45fwCgFiDEJuA2pKuWHNwILNo
7AWdo+AZuocJKTsS17G6rqFVCenRnWpgrw0df58ldUJErzxlTykwPFr40ZqSk+ycsjxUucREPMOh
iHjcOs2R3BSAiXqKeRCelSoTJjVI02o7i1Dw463IjLLndoTy1EvDLo83j5vPdc79pfKTb3Iik5Kb
HCHnmPG1cz0NSKV7THAEsLAXAZFPv0lnCzEmA/LZHJ3CLzi5zdq+cwok+r/+x98Wo1K+ek4hWmwX
yuuqebh7KKqyQnfd09gEJDVSJV4nopG0uV5E7Yhb8Sy/WjKpF0/47f7Qf8FnHGMeeB9ZMXIxMs5O
S5VSN/1Ran3T0v2OjCv+xqqjaRYyfsxM8CG17H8c5+TkxySSI2NM4/8sHYPbEN6Zg6smHDoNsun6
bTVkU3EXwnYA28iENfPslk6NA12LBWam26X8DKkDHgTF/c4n4kWKD+PoCv6XuOFgyM96hu0W+gqR
Bjifjemt/pz++l4LeQHKoZJKM4yCD7/b6qZe1lhiMu7L2MicLZG4aPrmkY1CftLBrIgxSi56WDSh
FfNyMW6auGBAmA9AOhk+yB3YUjqWbMKUNnqVjYZ6t0xHIyZ9hVyGK6kuNXWv7UdBTK1aTfyTCTyk
gWhDoS4P2p7MW1h/aZsFIbGrr0t+5Xknf5RrubVNVuBM+lpOE+yCRZM9hxc/RGThBNwb0JepfR3n
AtFe8qir18ft79ot77QwBLnx8Ezk1fc1+AoXRn1F7Z2Mo8I1PsW6x1T9obj2snwe7cVaE+utkqdi
i5qHWquXAOUseCgH2akJRwzSn5eOtbro+KivVyj12w03DVyQMUqrVgG9QpZAuYhWSBi/7AOgJTAw
UZqSp+7gG/8iXn3rAWH5VpaYVofYJA8RcfgINMIZHf4JF/E2UF0VBHsGA9Y4kkCq/A0wl+hGsCaD
24TTONsmQdnrBVwOOGq+A0+0wy2wdnpMSCLmXN8GuQ2cJJjsdJrOLDaPMCx8+aT5a+Xlc30ksA0t
NKVT3sG0Kr9mCytm5gW7OYpLghCyzZgSODBBy31SyoMms2ZzGxnFy5bEdTWGehQdyuJotsAZodnU
UqjMQOqGhhkHsteo8g/AScu2tAUpQ65d4wE1bXyGR4P6MDgk9Jo6C2I8YqSTExVjfxKjH+7Nr2La
Epmtpnj1GKY5mznjmkBKD/lEujUE+zBFvOjvnKIAHxmASoOqzSC+UDfXrppjm0G439kxolW6cj9R
qJrhgoLRMsP921Ey2dCVzy7xydVzTEntyIUb9Bm1vhcJG2suQIZOKp+0nvDHjvnH4b81EV3FiB5z
SARs6PxKw7+/FDrdXgCxC9fmGJpJw4vTVBXWkiqWIUkrDPdJZzedkdcUxnz8s5E/h6CkBMLuIxgv
0r3GuBqHErrZLPzD/iYtLEAJhPVsB8ow5lzXo8U08GFv7NGEh7/2HVnS1msUqsqZtDcwwk1qdc4U
FOqwjlvfpC9dF9YUAWAGZz6chMatUMNkbQ0KI2mLFZ8LD2kaD/ehw6slE5UncJLg5Os0lQY8sRaB
3ztfrMVpYYSpyrIJegPf+JonEmePiIDSM/CcWoBOFu7CLCwn0GKyV+dp9mRe2Oodq+CuIM/4iz53
52S4xXqMTENXGCeRDtBbluKKd4m0heVhZUkRAoEzTQpIm0sgbyV8PtSiKHtryqW0MIxAvtVlrtD8
cMykTwsV8w5lCITEu2Q4g3l4kzXZRbHleC3pexliy/F86UiifSPmG/MMaC3can5nHnpvWkhQkk9X
fk+Og9PHJVjvossejjJXSqC4SoiLlp2WeSu+dnonEvoKg27aw4kWZeC49wbYGGIwCGej/KaOi0DR
RCro2IXuYR/tUw7VNqwx1x0nmzNMuOn/Abrozt/HoGBZ9TzFnP4Vh85GHR07ad/JxMUpCYNHXnnf
cKWOyAodeh8W/kU6OI0WXBWfkf5Jv7kUVO6jsz2eBtWak3HNYHEl/nt1XgUSpnWHaKwd7qccZO7L
H9fiC0JEPEH5j7ctwvNuMsE4ib1JoTLV0tnRuVDv/kDOCN3i7K9i3qSsGPos4DEO022lbgj1JfyU
uRNDiYCITkHpGcsO/tSfcFgRW8Ex4OwMAdIlTLuBbu60uYsOBOheKe8nEMasEqR86R4HGT7VU8TT
v7qt+SrEKRoUWHladsvPQ+EI6dzVji9+jTspTMygaDhv6hfQbpZ3hlV5rneL4D+3sW7qDH1uwCj+
QsgEKVbfOmefa6kIXLsH4bluueO5D5ayRg87iGdw6eEkfQfqH71YyCisP1wKOlGs/vPW+JTBUl/5
VEGlFIWqNTADWILs8c68GuZGE0lIA454zO8FEOkG+97eQcQ/n+InAJiIppIejBQ/9yVnMmMIDYxG
qYUGhEFKaEa2FXQ5BcjqUjkL1dLo+DshYe5b7ufD2bXsfO94I0XvQXrXcq2Lmk9WHwmlUoSHfXwp
Dy61m5dcal7TgKkAZgTt3g/tKTHO05G4xykGYbNIDffjZj+eouC6lA0wQ+asDPlkqo3J4fapK3HK
qVHSxveR2xgJosna9Rz/QGutJqmpCqSXJelwSYXy/cyWc+cCLVmtWTLYKk4DAubxE+mtlAYgTQkC
Tl72lgLzAqnnrs+H7xjayUdYRVtJEURXjmf9VIVncSe32BjBnOfn0C3vyNxGHEdWrU793c0Ad7fh
M8vNCQmmQhZhd27yt+9DfqD1P7lMQVq1+UDtyK9Aaz4XJo/oNROWzLTqWU5jHlKOYK/EtojrvcK/
CAhk/ieJfVqWG1PtyME1e8eyI718iHW4eCpvj/OChOyhJJ0aXj+IhEOeHs/14PM1L3B0j4GH3lF+
gS4FisiWjiHy9rNZTWuwv8UY9HRpR+UpghN4oZhROSAApDQMWdhtuzWgFGILh/zX3CUNvY4vMOE7
kdYX6bTTo9xk7wUrj1GYtyldRyjI2H6jubTW2ENFS6EgJ3TnmdOV29d9vrK5sx4QapEPzg1CPptZ
QYyzDAJPp7vkZk05YNWtQ2P9p9eAvv1Q+0YMAagTklYkrQhTjz+S+yfyXmbY1OtI0ybXBeaMD7lp
OVtzUrA6FmmTWqul7gMRl+EiqdcG9UqFsKt/iTzZgu0BuokKRFT73U46yP9p9sZJOcLsSfWchzHg
KPWYwNBM2Xd0xdmlW3aZIuH2onNPQVKSXsnZBhihnFsLm0dclxtROihRR95VPKkiE5Oozb+B1gLQ
Vm+Z8+HHUNZrtMs+jPDhBxNLQMR90ek2TeyK0wCNnBhYqnDc/FylSkV1y7oPuKs5rf2KYzRqkIiR
ct+pNhYoEUwKZ8Gsef0MxXepFXIePrEAYqEZGNby4T9C8H4Q6c3h/L4BJAWGstHDb+k5HSG0+R37
vduWkWAi3V7rbhWYDNs29J4vLakParwJqpmksa+X44Uozd2YJT73BFLqL/uWwXJ3LBProTiIrNbw
T3+bdH/su5x4QbYaKNvMnh887uYjyZlCStlBfC0XiH58btcVowFOVmRZDgCaOszut6Ba40obCSJD
j2zJdnSUX6llEOex3V+HMswcVPhzJ1I+7hBQR7jPP6k7kims9xNy6sSxvJRP5zkFbMdR8sVUNVPr
lwxjZLAfT7umh7zyfoEfTPflcWqOtMmk+wjW83gs5oxtnF7aMrmcM4MRXOO+uuelidbM4WPBUJF0
67p4Oq7RyaPbWC0GvUzim1U4UgVFGrNLWPfAqMnBQ4cJHnRJq5b1Qj6SIBG2/XujeIl3f2Llfg+L
fClum5I2k1rpDScyzs5PFDHIXGXZLaxiIlUPSwsoBKkOe3C8S2K1D+WNfyiFlwEo5miMBILlAoIV
kk4rFUixHNSnA2WRLvym0+JgNjlzzogLUbwv7AhtKtVBkMpe9hJ/NcxSfON48/X1pM6GJvHA3BT5
4sYD1W0+o3UOVBr+EYILEQLQmhLMhsAEI73+v3ui1c8hxB0HXY3APprvxTgRAQJGRXV9NopNQGYP
R4tkrMwuMMK8TQPCLMCofsXeRMalpk2kGpvB2HSlvGhUG3BrVGvS1Ll1jvSOYRTvihmd0Y6BKyD6
Kzx7sitOO1puO6l7W0VbthozKNwU4B0AG+6xwtXHAg2Aj/RaajcO4dtNZfQLo8hWVwstmTwNbhPR
WeIjlbniCvJYUxERj7PlMuzE/q1lcHNOBIbuEtTyByHMKLUonya0mWx1LgG8yZAop3BhHP7Ov+HD
l88Q65uwcIqRlyNIsiYV8bNVI21kxNN6ogueT2Xel+ndJDYlHcQTfE99pWS6METr/xtV0V+5ez3F
yxZ/TCq08qHhnzAJcuCGObTytUi+CjzaDRU93lTNJ+XlqcEI6/MTIcOf9LtTMcRGaLK9zmeA9M9l
KyYmJ5hRf/QUoj4mat1TE7cNwFG5Jvmcq+OXyInXN1hWm6osL65cmMvUZ6aKjwMjNeKKBtcUUKQn
Nlt1wRNBXavhHq82MM5Vr5kV/EBRfonzEWqhDTuLSOU57HRHrHBqVkc/noI4iFTdvBVMfVpvS8/b
iuWdjh1EaKLM2MrHGKyJ7UGpLDMhVmv7FydFZhc7ajQbqtivEEv6fDOdcTiHjN6wYQJvZZgMQLZU
5I7vTGbEfVVwlo86wqnV1nnWyC15FIbE6d4HFTx+/mNhBOp7kHFSCVKxKaU4rxw4eNjQEJoje9wY
exkXJPHtZdWd8ixm3UQ7q/RE9gz4kK2zTu/lVoucfGr3cVMA0qFYfdVKvCVMKMsipiAZ1bkM3j3z
5Xv+EbsuNZ4vyuExfAQBVc07w2b9rAQD180Nu01nGUfGBYiX01/8EL6wB98Zz21vGn0kdmVEmIeP
Mi0baXlHV5aZcFMfgri8B58IrivMPRFDmPyB6MPHKq65XnEDbAy+h/P4T52vnyVR4a8Rc1T4ipzs
eWnZTrL+WpMWGx94Gxh7a9GBEsuliPKHroRhx2/Z4R98mPnbWAUQAXrf5AxxoxCcsuCOliQ086dX
kmpM6jcboYgsIB+oInDB0e7aQmuC0dDaJZwMlTsma+OLI6LlvYfG72WJILwpsf+Gp+hyO+2i2i2X
/kTWlgIHBwf6NJ84XT42DciM9BEVfOa3bdv8b/Cjo1ue1ZQdOTMOyvvGzriTQuctVrSisyiUUBPS
bgqO+RwEBetHioTxziEYnUVnf8FdyuIB1jfEE/JjCpURcit2rIwlwLxcQL4ND1b4kCAOJBB/xX/p
q0QHvRzOsfvlT7M9or3o2VQsjitXTeilg00w7AbIBG861JUYsCWrAcFbCRkrbOHvVKAwVjXcSyYW
mtleS5WSMaxsBmn6Dzi3BTixXQrNQhnE3CR7H401XqiHvbYX+bjzpmL045HWL0bWqalkGBfJLzyC
mLMUc7PjdEiKkGr4k24pbcbQGoqwMCBLo9zebCSRwOQS+aSZQ0yLenWzot6RM+6g7AEIXqBB590y
d0eGY64AVkaKy9Uzrg8mZCdcGoPrYCHr7ztsvxE12z29pS2ChAXlOim1b89hMlWReAf92ZoG8Xz2
dgRndCMFAsRdGNEepaliWLcXaTnJzHEJ34hMWSSGOEqpKSsobPB4QS/od0kvbgE6dw3LwzP4IxpB
5p41BulVJzsO+5gQbV5sCFFBCoWQQBTE0EEIYeR5VoxthJHASrNgx8AYkTfe0rWRm2ij8rnnKV9D
loGxOdISLgyJE+m6el864OpSjHz4A3np8yoRWhMcMasNbm6Bs3SIipzxMkk6kabJDkja4QKuL7zn
71ARPKQMJCFZEERzc7qZ12l6scklLSK3xQDP4Xyuuw1VLyFLO/pLQq2jT8+xwdpIb1mJZd1yBPaw
xzdKh4SA2oSuMEgeUYkO5KgkcoX2gOFt2XzDQe7pXm+NqgrPqIpUcRca1CKdMNQSlV8VV7oeGQS5
VQtp65rYluThmNMyseNUdsQA+X8NigxcAHyx6NxJCTEpjjR8f9F8MTKVdhmumxvp02tsfUZJiTvd
bmucefBphIWzJtTKtHRdseJQ0l57q8Q9E/vFAgc17FzOcQiceVLjCgsp7b1fu9HSigaIquYtA8W6
gftMNvfoO21goNAanm7ZgpoGbROEJNCuc97b3YtEaLebo2+8ENtCq1fWmuGOal1CjzD7I0jDMJGN
kWLLjSVh1VQj3G2IFINVzaXlRdv6oFnNgmaIaKpaS3Kmm3QIQxi2wHjNaLmJ2JDmPSA1cy/ybtd2
5usKBhmAQNvbcyLc36Kqd/QJwiGPKUIHxWyj+vpw9Svi3iLFAl7sX6mVMNxJCMSCv/B6Ebmocav4
JUkp3GqnCoL4c59YXj1OyAJz+fKwe05+GSuwPpHr3SMmYWJgkzT+8isL99Cb8J/ClhD0JUgdIFAe
WT3rxDBc1P1ZH8tGkcz6lhV1hEjffQg8Ih45cjFRaueF7Fl9eiWbas+bFsdJIz29UOOJO05BOiI2
bNroY5iEM0c7VLNYtNhWl01GPcvjjwF9XWlCoeLASiaoMhL0V8+eHIBVe2JlNpzXw+B3hflfl7jZ
v8Eqf7Wzj8JjbTjN5DZc/8B4y5dz3xmm2jwF5TKC+x90pYss6WWLhqGT9P/d7gsZBBiIyRUAscD6
xeN1p8C6zhHayHHdCngjMCx262KYfBce6l7Ip6oYsRsSgymQy+j9OQDt1NB/mdVIflcBwwzwBLDN
BLjpM8bwynfrOaWt9+hKwAmVD4Y6BtExT8Cs1xIXIa4t15YqN6aQFYX9eIPoMsliMZvDJIWseSYC
d2vrUCZKD2uwqgaDUJKmB9Nr40sF+14kAxcA6jiNrXdnh1sbxcOiiu4GbpSLozgsPpxRlhMwjAoC
JvLiUlE/wCEozUqt1XQlhhX0CFRc4+3FFYQlow+ekwiQAPGkeqXwsSy9s9UPTMkWJgmoJqst45hP
q9/XksPFRwdz7jQ8D+LOaWIC7QOz12VIBSbEaNRVC4w7PIy/bHYopl3aNvrVLp1wlqr3mOibDUd8
49ghBkqqQ4yT8J+lB6U4KeTxsOvcjgqLWmE+oaZ7g77VOxytcJ1hMunH9F7rMt8A1ST6KWGGjoPL
QRPQsQdR2Sy9kWO2K6rpDFCVuAtQmhSyK7bZIFS9efCWXpIraOjKRt8irg02/SqdiycwrCLQUQhE
iVK5CAantVJSWhpB4SHQYFAA2/0MMEeR4HuXI82bju/H8XFXyqzZH0SAAhlXWzVlJ4O9e0Wx5Aex
/Rn1rMVhfakZhqcKmwBmynlIr/UwUrdd2dV9Hj2+fbHLfJG9RvUuUdv8+RgVGZHUJHdMr2922rPY
qen/n6xIMWCJ9w3zCvRMxhGUBIZ+fUax9+EgQQgpn33ewPB/ZH6aysk3oybEymOfistxo/cbgtJJ
nEhEQcVXAq3kyo97ISmescKkFWsUPD/FTk2FytLR57Jh7zaaCzSJ2sdw7faS9sYiIukli0AO2b9j
OyTanf3urYVWH2qcgmNhvK5mm1eAOPUy+zh0F742TeqDUWUFbU9sus92/tdQuGtzS3J939RRta3E
o3X5KwDP7OD3KaaRMKiw2OantK5711loi+VxzY1JYVbpZqDN0UH6+peShdIv1k99Uwyfa6uW7QHq
CcRtx7+1BX5CmfsBjH7yCeTELDUZz0XZWpr4nx4ErrPeMmI9l09RV8fFdUssJX/VU+MKdC3adxEp
swyMb8SQ4UfRNL90oe3BJN+Wy/pz4xlN1e90jLrGrZ1LijwVe75+cp4QP1nxgPffr9f2t3dWvysK
Udc44yoNhQMsnuuCsV4fkC62jFnBNc7dWYrGK2GWLTTyJN5xNJbFM/hdiccJcFUkIpXu9Tr/NtOB
o3cu9Hjj2R+h48kGk4mCHNcdmwElQYI+iod9voqmcTLmmLw7cZg+268q+7cl2OvV14nlKWccsEgT
Y8uVPvKLwF/s365Sqe9l6MbdOKa6B3a5+0wy6+BjFbe33E1Jhn2pJZ8ekBYqC+QSxJL9f4gqeMwe
A3BWQjk4HtElTQTwICah5mSGq8Q8cyWYFKlki6SIcru4zAxiVCqPXkjUHF7nRIazqxSiGO2+9Flx
0zF8zgFGLF2cH6Zmr5rWjQFB+QWIj+eLKy2ZsgF7+4KqCixJ92yiJdQV34ZqHxxmM4dPzcN+Xoux
MWhCZrUGYX4rKo+aHDSH5nR16uFue9cTaZibqHVD4IWskF+kqfdX/zwZWoNjk6iwU9/Ks7OiTMsk
7DBb40K/HEpfv1iAioPXK2VyI3tWTxCG+dbOjKZYXPsst+FC99VlkVxmy/k+6K07qjSHOQsoLgRp
mdgfF/KCNv7PgrKME+VEr+gG5l5auFy80cfgSS553FndMzrFK18rWhibQyA91q0VPiAi7i7J+UXq
xir40Dvswt+iY+JN6thfWOVFkRwl5ed55i6iApLaF4LTw+AkDU4neoiTEHnX5iugQK1X/XQBA+/q
KYU0rz7rNFlp4UhovtqqfA0jt23JPMa4jnTe5Dv74qcqWg1mzSwgZKVkc1vPn5XivR1tEFDRNbb7
CQ+l0MkpXIsdnqAnmhcmnPyj1LC9DjUSO992h0/54f4Hi3t6B9Pkk5uz2wtIkDwD+0iUluVHnGYX
HwUVVCu2NNqItJmgkbTjWAnzbM2+H/xxxn96rexaIiql9BFroDg/itbXWmcItQHgqmflVNvxI04p
4dG2O7hJYx5Hsx80izK4zVTg1J+g64xfsnN1ncqRxfU8xZ6o2DAfNrSZdtoQiW07JL4NwMxFnEQ7
hebX3H5dO1SMqYbQ1UiBpDkb0Kp78YgAGG5Ex46vHXZCYtYdMksTzo8wZbbEOL49lKldmLaeMm9v
mudDAIm8lJeaCLq393Nh8nTtlNOSniRnW4rQlmVKxLJdIWIk14W32kt0J1hePnjTJk5e7pxt6MbC
Y+XKW+4c01PdXjAv98WlXV/UQH+JOqzBNNJi/J/KNrAOUjL18QbRVexpE9jDUFVyugYZ4xx2CFXY
T6xH1PJ9cp/zRxMebPutL9yD8y1Qh8sOoOUAgHXcKxfXomCPbT9optvD0AYsbdw/So3eWlaplVoI
tiOAGFO0BQRr3K5cDpNxBuhOKVDz4QfuNG7qaqEQclDWaMUKWsm6O2Cvnjq10g/SnA/XDPLDmRjJ
aW/cC6XVtsI1xO8QsAjQuMlfr8uTSojzz67uAznMcStw78uneifAYzLTLjSsrh+Ewcl1IJMZ4lgK
XJPAr6Ta+p1k5SGfeExb29z/aoUZMYfVNS6RnqREsGR7ylqanGfdhOUMun/TP3SfobFNAUugfEaZ
uNbZsOebBVa0ZvKrCBuMOMlIzF26Nsi+O1tfoS4tOhwNkD8xbiWs2r8WkSjWgfIKsyHxXsuWK0jn
JhZuFzMj7T9pFz3ujnpiNe5qKKCV2BCkomwlzn23Rsq8GW31FLqzdCv8Gm3jFpLhVHAvPLZvhFik
3rce/EaIC9qm7U9sqFA8I1WWbJwKsIGwxqaqWhmPi3fUfEy5PpGfGvuTu+1u17uwB99v1Ti47OWT
FtTO8PFvT1GQWlxXZtnSPe/2lyr59GoqS7snSMpai7HUniG5N7U/0z7qcfwKEOY/Z6MUMRIBiUGy
AqXT27MZNqq3i0H9y7DO1l1WHtcTYqscyiKWIAp1VZb7Z1OzWn0ovWGYcMhfQkuovxtq0LOH+MAh
4OMKIya8REr71I+ES6+IL7E+R6dHjo27+xzZnPsIAE0GjDIzD27cI+0AQYCA4UYqwJqy3zSvtuMn
QpsOC7kX3+8eELe8At1wASO/A0L9D/4Ntdb0IkJsYgo99NgRyqjFC7nMAmeHVNHVSxDdB5ZzSr7D
Uk3luo40kXDU4jTW3L0qTXws92bnLTspo9XBy6lIa3d3hsXoIa5yRIeEIBxRbMPm1W5kAkAAU9xJ
OvdMo1BCGcFJFRvG1zBNmaeS3JKCUDjXIJsPC9SRvmZJRexMoq5V38Q3JLMbTXSO2n3NNaq9xaLU
kMkMp5LzNvmdNWhrc6ES59bzKdhrW/HjTm5CetB5uRJ+gdsERmPAEDhlMSXa0dTFGXNemYcHvqgO
m1AcmT3K9O4r1PhuQSOxgQ2+vu7m0Qjpxy6AJpkrP+m/rZNRFjvpsx4zUQrnousG23jBE9+NUCDx
/0oAPhYthVd+UungMLEduwv8dpPu7QdpjN0uySE0HRd+PyuPHleVKFPGlxPhhPMZXDV2gi4zp5r9
ODY1OiU5crrEyGUy5OS/KuDeybtz8HPlsBfljEj9H513DEzHVn6ODVuWyWaKmYAuG25uxxKV5gw3
XzQY24YDkkx3kIQcDE4WEQjnAvicgXLvZavKkbPSf2jHK4wjc7j/3ZASHB1E8fa6/NeNWbA9lCbo
lLEcZe/wOLmGresLMQmCe/sMksX8WcZN/Qz0uQOJluEa4CPBwvyCjThORPxhlQTunfoqzEP/ZSl5
fQy4P78Tuv3nOgY7zp+sWhLYEOUUno/4Gb5mZeO9PFzuhvpsgMHDqDARkRNyFIjoaqd1cH6MX0ze
260e5kClpFLmfjqVnmkHcgmX6k4cyNaVL41uX5d1vqQNwijEcRqZZTWwfsdFd4krL4J/bmBYZ/mt
zIDvg2nHiDXOeQ6CNrQ290LFihoE3uQXvuNYoGBbupLkqkn6J8EiL7B2MSwinUzqHfvqPNJbaVbS
SmYMqjZ78cLp9Ev/uqHCR+lYla7KjX6gWstad8fyWrup4c2TvVUBjV1h99u3eD4LXTfT33l9CVT5
+YDblr1P0hqMOgofNHxsHDveQ0NJwSVjuhE/46mxyQBT7HgmmW0AfAII2d9dQDjATgB3wudAkRA7
AJv5ZMEYkYdc1lo+Ooo4dogR3K0CvznaiFUByKyTQdlKDeMs18qgUvJE7LWdWrUo4LLCv7rbxPwM
ubs6mxBOBdBn7yQx4shfJTtbp9ndoxqkEfXkHc3LplmVWArQQR+KF6kLt+9IrTm1B2c9Oqq3bAtN
ikD4p7kYS2XsHnR27scZpdtrkLAfX6KStXESz54DFMZIfBi+2Rbooea6oIJ6afGcPajdk/xZXIr/
d3lcePgYU7N40n7r1mUll3n7UxYYaz6XigHMOHMXOObt94Lo7TbPyW28830fWOKyhRb35/DzeUO4
e9qStZxD9Nbo78LTeY/6M6IX7ihdb/cB5aUQqPsCSlSwJEJmLefw9jXwZceBPwc1i2UwpVJUmNmE
BUtVsBLeYc3GhtU9H7FZNPEn+WpXxzJo3wHZoSMRwC1UuTh/i31HXGrFsY3RZtl35E500KbSJ+jp
LCz3xK4AOM5qrBtIfVVc29NI9+Ab4GTMYl/+bFTNwbDHtzEeeo/9t2OOhKoqEw8+kLGv8wDwU5ak
lQzoCovIV8rIU2HKZmLp5ize9/mWl9ldf5ffwggLDvL7zvE5lvOwRBvZe7E1jD+9wCRB2dIsIky9
Y4LVC5GcL+gSMMxFl1IlrIxgBObqZRvjgaqCCeVi1aMlxdSfdCQuniYi6Hd3xZ573laH4AsRPFiK
s7rPWes3hKPzSh+LCg7fjBEqW/9eo7uhvRuywdu66D55mIcgqtWswvR08r0+07V/F232X5+R0SVa
jZx/QzxQClg2IBPSUJ1GKZIrsAGSdzH/LKaLiw+J9EMAc2YJZCjvBk0SLPXGd3JBkD7lex+uF1J0
B6N+JybdJtn1gxnOPjQ+8OoWMyh6ES8TQ/QQIWBCCz+gv1UTGU+L/Ekboryz3YSz9hAWji/ZDkx0
ZjUMmHXBlVxR25mMfyq/y5qRYcoy4ELqc38/3lucsrU1ZdZvQ1hpjIx0AGBhwiPmxWxR/JFOCMHT
0/F8VU+19Jvoh4W09WGhHdwaaVtsdzTWU3iiAa6uQKErI64ccWqCImfV2nCU5zpAMPlZRPXnADvS
vpDcp+Kzlfvy0vh5g1Ij2QgUXGP9busdIxVtRMyMrm89YvWgURXOwdnyvGXNyGfcNXf40zpR0rLy
GFwOqVy0R3WPgjoTx0W6ffv2ck+vHvgUAvoj9GBJXXVTYSKHUpSIf9iqiaydFEREThd+J/ajdsWx
GmC7NP1kr+52lgt0NNd6NEh5DUoHzq9VaI10cRCHZWJ7JKnPd04ufV8Kj96qOLhczn9mH2bzGklz
/WgyyIgC43DMTux+WqTV6mTrA6X7BbGJWwT1H+6WShZB7gc/6IBrtI6Tmjd6OAJbacAWwgr5u3Vi
q5VtYK4PTI979P7QpGXZ91+SRWuUDPue3ijRixxkTCYIIv/Xeg14XGi5SoIHSFJ9WMz7eekGmlk1
YxrfZBRYfEz5jo5ZWcO8Rh85mmoHrEyeySai+wrM9p8EDx/gqj4hLrKnzoQVGLLrqmN0SM1XrpLc
g27movuio8mi/lhWVBjTYEHe0wobuIKqvQVXVr9vVU/3hCgqDTdjnsAzcZ2O2j57gpjIMxBjuScN
v/hjDA+PMKe1JaR0zvOmwNwQb8z3IqloHDpB92jpGt0CegCYCt+zXaJwqHgkeeIHmMc9rNTeuMMo
OlXc9ldj413G3kysJCpO32fLyG30K2IVfKjCc0Hot47KPkOnMzSAC9TtJqZBSdXAuTf7JXEG2vu9
+jVKZPA6Wk+Bc+urpsjr3Z4nwejfO2rOdapzKRQUb9HwALOr6DQW+bRMiSO9pl+nZNjGe740Ksie
HhDI+lSs3CUieNwXco5AKWQ/SGOv23SdevZ3HdRneoK4iGoRMD55q4cQyUR8+InWD5B9KA863xl0
07IT6NhEW9pp4dS1+ju/rYypCM/nG/6Z9ezYRk+hGSGbUX/Tsbjy1+cN21/p87OdN2ocm4CDPTsK
CCjtPCVSZ4xwmC1GA+Wp1N8VyHb03BpIH7t4LLvoOR6t+eC8ekukm/KEZ4mmpUrZSLC2henvafzh
gd0MB+eFlcKcc+t3rBgMvpmmDup/vupUowIqaq5keng/6gSt/3syWZ/cTMjYMG0dsho969DL1831
TEjuriH6lxCDqkvX0/N2GzKX4y1N0p3aC06pJABGD38LfDMdLEA0SauJJXv2wMsJtDS1bqyxvfEi
3h3rxn/vQpvTPYuojzAURkWYMiA5hUVKiYGSC8skV1fzi9kQpB1fObPs3R29Up/MMyUndVI18PeQ
fcdetC9reDwJa27Xc+Lp/uyCVaiOVvmA2HLIOkQvRTgMs1HyR86i3l253uDuJpvSnrECch6Y7rfQ
lEgWMB5NuDFQbrBfIB5ivwOsoZQmZ172RjmnxrHAivRGDrHGM0NxVJCNokHDjxKx43RAELG16vpE
x0AxSGm1EkrGVamOe+jhSE/lXjJYNHxnlet0FbCFWyJgr4N2uzQl1gHxb1R3EwINqXAbR2DXUhJp
Bejd8gLINel5Rpd8YSIjbHMpPY8noYg2yIKKSxj+JM993+oYtVORU2vwSLR8xJxU7iIC7ec+69Yp
Je4uA8qYskwlUKpdmKvp+gm7JLSH6cJyfS6hdkqgGdZJJUYjzIcqH95JrCTZf+4vnc4aAYmvFexj
eAykJS8p4XkmcAlGP+pJKL4cH4nQoBLCtXr3q5CiZucsF73GRkJ5Q1R86L9algYyJUBwfitCz0dg
1Kkqh1oVLR4G7rM6hQL6x37XfOGxSz25ddMdkWH1Z+21BtDfjvOSeP3t+1KPHKSJyLVXCtlCICxx
0ab6/CWiun3uVo7OvDA7shlJYQxsZP2zI5kJfGwyMDpF591fHdYu2kVBa+LljFkRrYOnOCvLliCT
E+YBov13tm/lJ1kyALOGQFbzyNASUjCwzS1ypU9aohE94ZnPvgo+i9Q20/WXnVJ0MIM95SqspwZ1
xc2PPcHBfHmPJYT1aONVEXdi/ysBXJRUuscy7uaQWW986zGo2Zhb1RA99Z8VlZwnY0Gtj4H8Wumr
DykCcdX/FFBJUWgg+WYhEsFDEv7/F6Pqhe/9YorfALAS8JRZrJEOo/KHdOvcUhi6vH4lHjYYa5d7
CRVoZ8r6YlmDXBqTRl2K+Aq7J1K0nw+M3W+Xjkf8UmIdEtB0OusqGem6n/ESdin+iQtlvL1/EIEe
/X+BADAS/gLo50XEIjFFLE3k2GwwQXyS8g2pwsShzc8JaPN+DdEpTWf3Sdq/aJc8oY1acVPprg+I
ivmx2Ih+MO4rXqoa1RUOwXMhZtZrOG9mrNCvZ2NtT66rrRAOTFo4fn40foGgvvZyzmgLMJpKO1LX
tOMh/ZD8RdHsVL2ifhTS+v6hY/IY0sUrW5HFfYqcu8aTB3c1bohTg2Z6bg/q6SW2YBLb0spYl4cr
Ap8ZCFH7EAYh7PVB2f8aToo/ekHp0M8/EopJr/Is2NfmUZFbtlhH1rMN+JN761+MCL5KJDbLkEBe
mkzZ19IXA9lKcy/QTDiM/tfjZ8qjzfM3fg8TrQcQE7yqMHMYnP9hJLjFEQzKAWkddNdg5tsZqmAr
P3BkEEgh/X4Zey8GUXkWHi1hKZYGd5cZUY0ZvgJD1ZyiKo6U94OYbBYND83PasZ6LL2zb0lAcm8o
f45gZXjTCDwCuS3+YxnEm7EenjvQ18bu+r7LKRhH+J23GSJE7+A1fNCHKEv/hTiHjF9CXVzl1yf8
aFEukDobsWE/5hpXWin9T0RTSGk6UbBcLmHHTJboK2+3g2VUru1+YR8xwM2tbZ8XPK2Roh/xbexR
R6itfw1V6B77lgc9FQIB/McnFVpGUQGhb8AvcxV6rlcT7/cBXcO/+q2lF1D08jRYZd6upEVnc52j
W6Gqus0RpmvtkrhezCrQrwTKVRDb9fo88L/jG4kKVpALqlEIrbtBmVimmvybica+jOOGYhIXAga0
XNmQ8mitRkYr8Z+w4AQoCjlfLN6pIXy89xgo2j/RnUKXvA3QYrLo9o+Lg+guTKGmLXYLtNFoXb32
kWpp+scJMXce1J501DvYmrmhzyRaNVf/xX7rRIrCfpY5ca5+n/ELT968A+Lkcv01JLfEOa9kMgUh
vqRKP7jHF9BXVHPaM5opObghBmymisFZZPUqC+z/fWaioPFlkfPGSxdqG3dBmtblImT3WCCyDw83
LK9xosSk24igIHX08ErbJuxZcPw5NCICkS0F7XXDeZgL5Mc99AOYeWs7v7zSW0wZwnDWjwbbxqez
jkk3JM3rD/soR8f6lqz0DkOxQoASyjUULZCebjlydgdgvZxAVzV+FgHNk8bqyYAzLDJfjjqfVpyS
Phz77L8GHYTCB9ZQpD4P50Ycvno3eGJuNHEi5CfQdOXsZQEY4JOrUzEb6phrCIgTK76w9St1J9dF
ujc9M3HT7/xi3ypWjJYLtswhPbGNkHQufdP2WWgSMBDPfmcmVhenxBYvNN2g+ev0xI3DI/SZn8fM
f6jQmNwe9iVS1m29Q5TMwwhvLuSn4wnRYrq065RS5ZdR1PRfofzcaznlcXAF6Glt5N5UXZC6HXC0
bvMvZv2hkdleo22txZ168S/mhHNgVpwGPU9IxnmdSLtF8MwXtQLHrSYcyVmU7BPlmeeWXx5DOXem
AQKfaMPrptcEF5Cz830SjiEE9p7CDN8mM5boHgVCVWJmSLFA6ivKWFmfuhXrW6ttM78a6YYM68Lw
IwoMjJG8nkbppJ7r6yOWcSqW6tGywSP5z62CBpgI0jEmjUmk6fx0vd051NUNT3DHt6hZIiQJVMEJ
6erBuhdq8Z0jrQjtpqlnvpaJ0Pai7tSmpW2zepTQSiuJlapPj94vJAPCPpQPCsDg/Vra/aKY8455
AB8xWqWi8ayU2ABkBXWQMCq2oxzZa1MWDre9dwFrTB6B7xRhWkvTzP0dBu5aQdCB5ZWCkGHFpWrB
Sptx7+PdvLQXEa+bZZmp40teQEjQJ2RZNWsHp4mStBuSf4Rt4ZqKeyMrEyrIFcv9fLiYtMOTBBVQ
yBWijzBEqHZb5JEZuNOHfWxyasqI0nPxPSXPAVXcnmsBbwN0rYJabsDEjydVC9MCMtLWMFVJQWcj
5Y6A0QpijfkalXDH/plIEpvfxGWP0ZHNce8rCBvPGJBi5B0bLE4kPit754fucSSJaS+v9jA8L6QI
PUmc52NzbVGRsohQ/t62TcWUVuIMurcBMp17JlYwzzaQv5b9vEU7zCkHyl+Ep3lgoGRYvJzEkhLG
XZZ2AIrTz/0dJT1/6TAb4ZrampFRwd5y3OUKdKGJWjjeoklNgll0ddl/LCeWfSNahEGu3VCefjTt
YANZTCEc3G91dskq5cLiir4EkOnokMq499S/l3Mbj1pUP9KywWyvClJwYah99e9oCoq4vr3OxAXf
1+ebMpBKMIablQxLpHYjhgX712o/jzyD2szNFvBWNizvTG6IUlAPbQCJM9VQ/9KNa0jjpTLhbvET
C20FfvdfTrPNkwcE2nYp8TvfkXKNp2nNzNbQrtTeFKd35v/uUdCKcQ9wiiIHbOkD8ISz6gkZ6mN1
PlRVYIgl0e7jxR5MI8AP8BWJQQDexRfQONUxz97PAJjiDucaXj2NbDbaIiE7nOVUPA31nEUPa3LY
QteXkTnL6ZfGfrmVJEsePUoRRdIi0V9G2kguBdyAwj3tAKNVnCY51KZvOIyqFAswk9r4B8T298hm
eYZ0kwGDZLYlP4Y5AwxD9R4iUBFW8Nq/0rcsha0uEfD8BUPAwGMFeVBF4GV1Wrn0wLfmeWV8zzS6
CeCQHHMdsjoVJhVZKRzZq+IP9iBqDrolrFjeaKmMnQj7Ho/YSSopQX9cg2Q+AxhRkbX976fOohUb
GJbvlkrH+SJ/JNJILg6PpLSuTfpH16OleklABhF/s4edf+Bo6iL7A37Re+SpaYSK90qtkMbjNryF
Jx77g5EVS/M6WdGRgvgC3qtxKt3tfy0soVJIh5lCR8ZRc8OQhRS/kbzPyRL+UitcSQrjYedWDt5P
xfnN0eNUT3tmRoWaK7pMHTAeO08uBxLmJfv3OZw5/g4jjlBm4EojPHYE8BzJewL/Yv2h0WOxVja5
KARwQ7nihvgSsp8ZUY0/lC8ABbhOoLc0YVxJv6ulnDwxxoWH2MgnLeo0igHrXOVYhXe5Dr0xpXbB
HeQ51ohoz/eX6JBidea2cZdD5rFVpIoJ9SpIanHHi9YOrNs8ZfOlMZk30ucjIQQuwB34JYYMNLwQ
b4j7FnZkqEk5ndq0vAH14obji1Uby9D5CGqq48N+NVib7j/iVZTTGnH4y33ojLxKXSl1RbwGbfNC
ewr+KzrlZkoneTgnZyIzp0IVadLDmlSbkeGpV5W0lxu4N4UZ4ARuoASzbZCPsbAQhgPYAsvfdRAN
OSaQZv84sCPMukpYtoCme09XAXYH1y2GLNcknef+D/W/NhWkSF381li/lJBueQUXbxG+u3R9uyRG
Kl3AxL0im3j3ZyVkkQNgr5QhhaN2+Yr7ZeJ1kxlq0svAwNDNWMjPhZW2WVnBwxPAm9Swikv8YZ61
rNZhNycr9fQT1XWqsuMJWGpAan416AS+5pCCWYdtYFu66Zem5C2P72YEOACbEu1LH25tYQPNYz/g
fQUfrTgOpS/jceaT3+seJrqKcQhDRxNT47qBGy7DCF8iKO3urQl5rP4agc1rKTtoM1zzVYfNUUXG
RI6hv7N8kJvVJrk7CQcbNxrXU0CyrMMl536ccTemHpqWQnBCnY6rUTRSk4rKTUWsROfcMC6QVeGh
aNg2rGocrJ0ntSuuTuTJZ8q3Y/x2wUZFcIyr12b/D3fpXvKYPUEFXCmvpL15JG0ZFf0YglngXlgg
gKCgiKdHwfQu0q3HN2j9kE8w9kRjDUchmIl7KVTp7TrUr1likxVohezCIvJFxdmzAMV8/aHD+UjB
Yfl+X/XI8rAR8kt3u0BaeK49NtcS0sXdLKqT8XPX9IN46JcKo5TEicqB0E8HYNUbsB3y4WlWfDDO
hfTae8MEzc123z121v59q/uKE2KH71bdA7kcx/aOX0wh+bKkgIwJRzr0ug3+bN31savOHwOiEzGi
4YSRpMBt2asffO5a/GcaSEqsBJP0tXEUBbB+0BFBAE/QRtOtzH4a5h6tlJ5ExKcn3G6v4MAHSQ77
VxzoJESy2N/gP4jPhA2w6Zyg22cqng1sFY2Aixu5wYGB/Dgss5XkXWiBP4rqqRey9fKfapbeGueB
hSie8Q0PhbrtBIoHv5zFKXk4VMllVMfH3Vcc3DiuBHF+wh+mNw0VfzNZ7mVHP8X7J6zDWAhBS11H
mGN4DhJp7hYdVQuLht/9dnXGe2KxelswjULWXJ1mG6XSV2kdNAgN7IcmHZVdj2X6AKWGu6yezuIs
H4zZ8447Pa8QUXTvCq1Tf1+Gcn6v74IHP9MsX9Tfm01MK2ZSXLVzsD6M5ngQci60P/6Qv10mNq2Q
R6ir+CzXEcGv/ZwpfWUoas8lQKdiezkcpqe7ywCrQSLW+oRCnyAAqJsbszznjBzl6iNGiDPxdbj5
7O7bkv7Rj6+JRfqTHwSM7cfN9nzljlwvYevKj6m73phnThConFmx27qpUZExf/WgeVamsoL1zBKa
UYy+XkZMpLpWc5BO884T2C+drAnDa4LbWDFZMaC923IHiYNUK2rfXdwKuihWLwwQnvSyfvAHOCV1
4elRyzld5grp+hfOhbB79WtcK02WfzghmtKad4+7XPQag5ndVth0rMIh5W6GcXRqMm4NGBLTD1OO
hnuY++6xzF3tNFK+nWy8JFdu4r+LYsVTBLiElK/wu8PI50xRO1FtDX1dPLRz4GgSBguVD+1EcHLl
jniyfLSZK2q5E/Jz76smggkuUYBDkG3BFJdCysrgzO522NvGx7VE8Dpy73KUCm50+0HhjdYLZ7Ky
ls6XVnXCGXhnMVEKxDwWz5Aw/NUrjD9J2ptB6dXOthTZRfE9Gj68RzP7Kv9s/4yrm80a3MidMkU1
IsRl6Tei8Ii3+ElYZVLmHD9qYSMWFwu/67LAhYl5uvEtC4YGY56Kzpb9z+Q0fS69jzMukCTV1mkY
szH/jFzQzBb8AMYNLMMCfGbhmQUtR4trABkEGfSGXvhzZgxj0rfZrfD1s3YVKx40I4+oHrOWAGUw
3+zrc+l9v+C/2j1a7pOyybyLaLmzkdjzpX6v6OQb2J+EQy/MZQrmp9u7RqCjO8siWo7XcAEWI5l8
KfCMdhATEwX9Wm7pXnCkLiI8OjUe5wetsC1C/1hXVnq6JgUU54ZuYwUszzkYpX2oIjrvNFrdyK4B
2tm7ZR3uUgFbz7gTHncoxRMB+YYXvEm8BOsX3Uvfju7vUlImQwtdblnc86Fk/ShqlqcdSa5DBEWV
dyPLopGaEnHVCGS/FONM5A1yCt9/VvdvxhBogAf685NNZzXPEuBu1ckgL14oo62GEg+SET5LKrhj
9fvt/dt8ptknVn/3qf47IRGcGfqcNA97/I9Y93R7ym2F5X0+3dcs4t5CsApefgm0J1PtdDt69/b2
kuVKuCSx1VmkQSgjQFXgZ3gKtD4WwkSBI/QSWGJZjJ0T2fRtgIJMWYPnWMzsQuvu7AxNQpXuIZ3B
HR6mwsP5cTRcup7nl+/wbmJJPHPizwMXtve7QEQQ7HdfnSeUnFY3qKi2/vBi2NaDRJmQoJ7Er285
/xqT7nQ/6LheEAd8BHT+oVgUfuPdSDIgHMCoDO9oGfX1BRIk+yqdKjM4tjwxueYPLpASZbK85aRO
k0MdvZhftRqXKI+0BWIsNru8tsfRpAKdX5zUZPtHNDsUdVTKUPrHd5RtP539RE6EdNrUlaPMNHFO
5fIwT7doBZCUI9wGom0ys/U7WtN5Aq0l5YYf5Yg6bJelDIOpfwoBpNS/PQhs+I2s9Tw7f9Lx1n7T
fml9BiFTOhfmENH9UvHoFdzFEb/R7PFkbgClWr+xj530650X1vZJDUoOFY1fTKR6ytM1LJBAMTCg
Y5swTcAn2nP7oM4rqNDdruEzn/l7rATgFe7UNBFQvjZndjQnZO9GBRvTjjPKGlgECLwNH+b6Aj3e
KlL0RNsgf4wRmhv6IVuosWhHb5mnbNrvghIOwBLkWumMCJln+4X1fObXTp26k07R/RBKRFZZ8Pfk
rIfNUwquRp6iBJI9rclgyVuQ2sTHzQH93CLIWW9VEDroMAk7bl28+ru3A096UM1VbG2QSQpdqJnq
2ju9arKhBSeLyFYAiR1DlmLRyxq6W5mj9Ldnsg+KI3Yj8V/3PM/dX7flBjHyGTxZLHYAd9tv0RBU
eripec7sX4kYZG264If7Et5HeB7BMwPzJ1Iu8z2s91Uul6oBAdTwOVQYRab0M+1zzqF68AfcjPdH
ER35WaB0ewhcU6636OWXeqYf9PWKLmTkaiTk+XE8PtOkwfW78DOIFzVFt7f0oU677b+nb0CTSuNW
vkD8kfGUJyLKrFknk3xZ2CNUxE36VUsCnedCGCUcVTuPoREopLYGX8pdh1T39CMNmvfB0K9CCio6
UqEvqkbpKorlLTE7r+iD9Rsuysu+2NDxaiqGyKIHTgY7WdvG9asaECSKPqlCh+ZZLhOJYHfbjV/D
//ZpFNzA3E2PlyFHqtJncoLbtznJxo1lg2C5S344TcUO4hKyUTPqd1g/kjgQoi0JR3/AU04ZCT/Z
Kn7OHIQvp890n2LMGR/tytYSP5kDe0uKsq8naBNAbvPPOrZTGYdQ+TB5JKLB5o4spKVgbvGK+niL
zecAbf+YK5ki/wJXkOj7CNjLFDA1DKnf5+kPsyHUEIkYrzhoRYG9kPcH8RLB8Z8BzrQChZs15o2u
gVUUTkiSleJz0RAKWt1g3iKJgca7J5FIciKEm3PX6HU+uObn1kbZwWlDOYGS4fkhJ2jG5L99i18c
rM47oSLuNharOklGw6bZWK2fzd82FmVkIWPlha6Keyk4uF3dCfiKRfwuuBROjH81Un1CMxMQjC7F
qkMj14zEbEbq1RmQxA+7PjU3PLaA9m28yqUqPy5mWnj8wRAWos10+mIZURGbF1OXWBWDACAJHd2g
Dg7cilCsiG1iHLwhRsEMKaQuJ4g2tlr6lBQq1aN4Ic3tS4FiiIzivPfChLuMxWeVDlTh/ttH1fAv
VFBWCuMtgBR5GnmiRb/n/pvLjV1xy4pzLbofqY6UAwFHMtxKuuXFu8ZWwg0UeDf2fVcwNWt5xdVC
8w3mLNq2w2wljrVQ7thw6QredNyF9JfgGZhIBtUEpC70CC+8y/8F/LpAxyLG/MGyt6ko/sjTpIiw
s4MnkVEXOWYyg1GX7+irs0+gqiMX/fPLpKFgkECojwRiPZOb6nbL3CQ6pguP8InwzM+kiDyFIOd5
R2PuZ8XtU5KOu3W28ARUGYCS7vQXtwVNvLRdnmsS3YBSBSHeL3WilQW9qmKLap64P7iwVifGWb8g
RuGq3FqC0o73xKSqm4/9h/VPXtTthOVfW/h48y+M3gsJQ7kz1/HXF1insTKytZIoMkm6zxjX4UrZ
FNi3xoxXIop6oMixWhLqXCdj2ssyYIcoqFInSyOuZIHFjM9DEaUBE9r68Tp/ClCROzIkMlLNsQ5x
qroRmq82KUtbEbxDCZu+oqHthg0HUt3spyOtEoMizIn/6uFKGyyuOrCzmtTtgxdW5/MavhLhDgzt
MuWql6v7P90ll9peecPzP4kqUMMTDtYTIFzgqQ4FA5NvajyGw5Dkjen2keYpMQzchmHE/56iRPq2
ERDMNLpb8RHTjNJdmvNPMIluZx5Tyo7gsq3e+HATVdk2pyW6L83ZDo15cC44j4AZyo6kYmBmx15T
fdyJtg7xwF4m1pv44J7s8O5oP1tI/QtTcvG3wOIR25oJ8Vuf3LgWBrqEv/ZQxZzJfw3M01WbjV8j
1RRw3riV8QPW+3zRQ938xNL6sJX/H6/bxb4QP0vkCObedTMrwZ3yvkYCo0FoE9ZRSag6slv4yPzD
It04lcYwwcoUejqzE4A5kE6jTcMYAUdr+03/AJjBP/DuXmGgMAHWbEVK55pis805f755dy2njsTD
5eHV8Kaz44nN0oYHwl5voklx8etUYEGvU7amLRsXWKDrT//8ZHv1aj4It5P+hbeBMc74RJ1xFmgQ
mBUQQWYVfcWL7rU24PQqdklHhtYiCud4lF7uc9CciJqvBPDHze8IjC6qjNtSzof1BgLnipo6Cj0e
5XK2bjhK8eBLINn9ryPXUriypSFyJz4odl3zhAKqejV9aD9AaYIjJgWhPHEKuJQTQPTIni4gYh32
ifV5Hy+RoM8R1gJPhfkefdeF3fhwmuXXJNL6oc56kIo6LIewPBuLTafqDEgVMXCzMDj1lBDEWrXK
3mqed6PbdsRmRR9O/ZkhHFByn0c+up2aL9cOyGuJM61NEjlXNV5oxkpxAjpz8EBjY/wr/Vwntx7y
rGTIRpkOIyNiWvhzUMlBq7DRmvkjgKN4WnbuJlDcn/7RB4NZ8Arz8cN58j6VWtD650v1JIlrfP2z
QTgbYdIQonNkwmTv+X5/UaZ/TZSzDbA+cfFZEfD/vkkhMvmz3F9Ny6paNxh1GlhOIzBB55IVWGjZ
yXQDQUyCZf3mjufGQaUywntMqv0zECM4iztkn05HpnvpfYpItQ2k9FJqcvddbvlmtrl0LVbn0W7D
LzbCTgQj8DgJNVgP6jTfLJ4CPcDyd7mjN/hVYd2BtvlNqhgDd1pYSKHc7KGdhO6S8garQv2xap/S
7kA4PmiMlv9rs8yNYuonYdsQAwS+kBBbD0fLNcNpgSGjOccbf8hMGHtzqkiHUavimWEkk/TXZLnv
RERRmwh8A3OxIVeyEefx7Abh1T77pMxktbcYnFuTbfh2igJ1RPuVtuefvUTEGqqFHcfxeoOKtZzs
QATAZhVACl2ac3IFwjMAbBscD8f2hCckxlLT2xhhY3LQOyFyzTT9GcSPV91G2zKlNlqjIV6+TiGF
DE9cXKbEvyB6T2U2wpHZ2FbNNT81P0AC3dBwwAJx4ncQRDzVB1qVk0hsEE/rbSApBNDrzvM0VUca
wv1fJWwJlET8cNqMxhkXUoPPi93m0soMPi6sYdty1KwZP1WfoY+1gW2O8bBpf8cnTzB1Bx8VT3lk
dl3ix4P2YpJ83N8SQ251DrMoudJQxRtlSzo+Uso76z95TLuxPnJCsnf2TkcIbCXrO7+kop94umCU
Uuo6NpTGK5f3VKHJh9nUd+gJBFCNSiB4XnofEkuHuI6lBmBMKg5JkMeOUX/dKnrowbwbgfG/wD0x
O3X3x+vJX+cP6GCoENr1t0dVZUo469rZnix+6AGFqP5ztvNL+DoPqwc0KjQlCLGqs1SMKyBdcwnr
TFDaOKDbotv4burP8n58X2KSvcoqBF1G4FEUd/7ph7LUbyz+ZxCvbFIJ7wYMJO+mOWl3zo1836RF
OInMu267o3fYUoA3iljsNT9ci5Z+mEfW8KQarbVArCMbqz18BDyd4N+1BgcOEaUqARjJcTU3vJBY
Uxxr9sPSmodvSxj+pHcwoQabr5aGSYyrOEyiEab7aL64omeCKKtkzGNVJPVlcAfbj7eTqPWZnhHE
7+l7e6dIoZwxY/qMsyHC8lxK3ui/PDrjSeHqUy4mXv2N+7bhDbRIyCfxXo+cWcCOVKc/NKaZpfva
RJfsErZwgt5yeL4HdUOIehK9w6NQZbcAWZcEKBREaDE1+cH5fi22v0lqKFaVpAJx2t5TsC0cy26/
uEpfD0/dEg3/J5RloB1d0wV5zYBb/MZL+3tPq9OWLmJMwtlGxVGQUNe7mZDGE9DJhFcz0mr/YP1T
2svdlY7dMdcf6Gi4C+yK0hPV3ORy7EXSlmuupZ3dqc/FK6WwQvwx+uQAB7zd27GvLWugnsWBw3jR
RbWX0lQJS4mo4dHtLtOC6V8uxwPFXYAwTWQjIIcXFTQL7axYHSmGEwHlmiWagWB17ndjIA0LDvk2
WM/d3xWs93q7lHqkMI9h7aw3EBDeQGNvdxbaACAMYA/g0eZk7XoBXzD4FPiHQD/E4de51ubVPOlT
1qzSTkyi/saOMCODb6RbBGG7PU3i4vMGF514GXjomp+jzZnJ9psRSI6UHcTxFSn8Yloy4dt1fZWf
aGcWueD4+pxae7DdBjIKWsBGDsCQ/YrQGJWm0Ij4w2U3ewMxEweqYEXz56frxRt5BFAXqIbgWy7a
ilf7kguV0oArcCwsIBdpS7tDfmDJ+uM4Sw01E6PZdT/J9ijqxMeo6rn01yg0sXYjIXBV9Vfh/Bap
60YS2lyn88B8hcWz+ifSxtWviDyAOOFK9yyUFFfy9Q5IEU48hV33hGYyg8cBULHPIkynWEzOu3oY
K9Dqftf/DOzOxf6fH2x0PHzE5Sm1NSrU/YbW6JR3wTF0+5LYwcMB4WIYtHMGl4J0btofH12KGErt
EydAY7g8QAvahhIGMESCvoOuNDd4s36BU4myyXrdC6MsIr4TN+RrofjBFxxhwUW8jHjget+z2Ras
3VW4QUu1/9pAfzKy+dMI0K14mnIzAoZY3E2MaApTNDLLLQlGOqB26RaDTgTPnBz3cTh8RE97QfSx
dlEFr9iwzxx8pTJE4TN8wREBi/RCmY0RBA0in1/1BQ/YMpvGf7LsEys5GReEfmF3NX8w6j955rcP
aEi/vcn4Y1rJlsdOMS67w11prmLe3GRZCkSON2LJZgD6tecKHqAFDBVw9gd2U0c0OQNYgiiFW4+Y
4fQkcXEMLnou/od37/uzq7S2VwPGHORG8OuCBGqv64xhYb/f+I98TGvDAIIsLPMZOIU7SFvCtkGh
BUDJyF9EZXBg7Md4SdJoQk+4qimvfltgCklbra6zgMXKOSmEaQC9rG9WfMrcmcHHfQy9eP0aaTuJ
HfsG+akyiqM9H9aor1P+R7VCdWgOEKzep34raj5cJSYhB4XpnmHNtRVaD2YhY333s0vRdPriT670
rTVDXdQn9vThSkvTsT5XB80xXObpUViLHoYwRG8ITTbNtjfj0+cCOMVlbNWrJTG92IuJqvVmBuaO
erfVpUrTMSWLYhkJC/fG8LUuQH3VfSn+59ZFUNR1Ny1KwgklNnuECaBTlpBkRNE3n+a4D/3GEOD5
UxtxdsKLedSyZz7xVLx4+9rt1rCOq9JmnDtfpyVtXWc0z+vSH9RwaRrW+syg2B3e+oWE4TO4TWog
0Cpj/3VHGPBYBIVRBONwBhd3Ue4M2nF3iwJO2iUgYsf7GcjqtZceJ9OufFRwvB2AN/pU70FdeesK
GFip2RncoKNIm6zdDBBmzoWvEJlgehEhQ1omuHDMjlJnc4A0fWX9tJRC36lwezCFQQwqBMk9HAw3
QaQ0Jkj4fMlfy/nDzcJuleFJf/m5C7RbQTbB2jMwYeAQgp7OrZ6M06ZB7wVo4spMi5FIgFHuFave
vI3Y4s+ae0PayweihUuS5/Bvj8GXzediCFR/spSQWyvCZTmfTGzxHmZGJ7pvnzITjGtkEzRb8CAZ
mcRFudpgMwY6CmsyFiUF2qfm/Dotp08/COfgErfp+N96gxhAJcdLL6nY/bKmmdf7Z2NCSLHhmxY4
f8kF7HDNi2IAtt6Fqkcv+ZYYmuPFC/yqTSxleoq+rYRNHNLAuUO0nEuuwKyv8OUkErsXdGiiA2pZ
He3XB2qvRwGx58oyTS64KEmEZWYSw/k8UUpOKl0g1E42wt8zZ4ICGjd4h9JNKQJ2ngW65i9vNBHd
eOKbTtm/Daw4WgqZEwciUm7gQnpFRSg0mUEZypmOqYPQl5HVHJk0gcV82JQEeSNLjAe46wVc7vNK
X0lJH7/+0fNiGXLaXsczVftPG2oypHrn36kdz9lUzcSfEzBqGkZJLZsw4OnBjIHhTKK4e5FIu62h
9FR6scpsRWFNOAh2SFOW38XS6sxuNMJ+I5VMCfsOU1grM08M9Ypi36tifGwmcO88eYENvapEeufa
hsrGc2wp/XtDaYQu84nBybeFkLxF/6Ajp85YnIvFdoAEi7qXn5RIVpdZmBLs6pC265XtP1VELOdk
8xdN+8GsOiZV71VPe51BvdDkdSw31B6u5q5OZbkRb6mPSdLqtEWemHlURoVIE9OTq0zej/HCSTfC
6eboc8J6dQY5a+Tnyq1foHfXHKJb8jxo4rFokAqkg6k4ownA3S1eQzxkwwDRFXypum0OWWmw1CNU
TM5hrrNLwOD/LUH9Sng44S/pkbhNKgNCpeJPSmF0VbwMR41T04Ecy+/pBKJ0aJIMSsPsMrPAl/AZ
AiDvFRQEH4fhmNL71VWFgq1E8TS3pXt7SKEMlrzeEGSddYM7JwS1il3L15HR3vONOgOcWSKWRR7W
P9MBvED74SOAIeMafoZZ2uvdm5j9iAPXQiWaDXrqzJkh8gfDHLuYaKYeuIZoUCmEC0lB/2gThNUL
HkPQOIN+ZMVYYyaKXRVmVO4bfUnv8XOBV+gvU2STWyfO4KX+m1KFlvQA8L63Hco+B7KcXaGREUsh
ZL/fUac6lBS8POuD3zFNpsg6wKm72Sx5UanBTf0mj+brOiCh9Q4RlwfDsq+dVkxrEoKv0QIbILjE
JkR6jiSGz/BT9OMzQYu+dRQOvdlVahyEIsElC/2LogBxdypXyZ1D7vx/+Ms3GUJo6RGGDEcqvTzt
4AUyQCKEnvhzLgDcYVbUaf9DthiUmfLA9wFleOpCl4hiJPwmdSdCgvZr6fRSa3Cph+T6KeHD5W4X
56Gaql9YYWACn3uwbER43XHHHoYX7YJp6CsmD0A0Umh0cbaGj7+mXY0GeUSo2FPfyUbFFc4CLNFu
aol+2M1WqPNjLZPXfCRseXR40YDSMXfrITCcK8Fpy8FSzSIAHOJSEZRuGpAaknLNYO2+ygvLInmf
19Q1ceykmTXHjopdO8g+Opd/0vPrVXKvPeqZKjpY4NnVM9DsyR9cgWROTVKGLPpGxufBgr++Dgc/
OllkSAdRfsYICP8hqoYmB0laYC90TsMqEjIrFObMVqD5B8Nn5NyFYalRcmTBmACF8NwOOfhdIrgE
IRYb75B7ARMG7WNfphsXfR6SELc+gMlJY2z+V4xRjWFNKbryw9nAMM31NOdB6ST14U19sMtg5JJC
sRFeb+TmWdzkJ492s2Oo360jiNy9r/6rQJLWE+gJHDpKBnNzmGWjCgxh3cvUIxwYP2gNDrTptf/l
sytIKxIYxCDQgQZW/1D95K0lc5Bj4ONst1y9sAScJsOb2fikSrzN9atU/rDmLuvoyiF0eVN7X5kL
OBiDZKlv5Gz5y4grb1wJd3BQ/JflKfFL+t6XIVv/khnjEqkjAV8DqQPPWrZIKFv86le+viXWXxRj
YMvXaCRZ8rwP1Bnb7D6hqpDUluWfZ+l4ncx1LJEuLhA5/48wDSR26sTMFHAKH2cdBoibMXCepYbM
DS0xKxV+uQwmo0HFk4ozdHJhlcakfWO0KLnS/grkXvfjkvMCmDxWB2Ck2KMlL9yTfMq7LlMJXEU3
R4tAPCDcZzVTEnJifYyzc5px5qAsdigFyOVZGlxllWUbyNPmqszPlLwmz4Z1dlAuKadwbnEuFEIk
KtopUQmnRW1uec5gRfxN5ZVl3GlhK/Q58T//9dBh2GMbc6jTGbIdhFjUkwbdzVWYb8BFV10/QPBW
+rdMw70L7a8r873nkULRrEyLYy41vMDSeCgBiWItMjcK49CZ6GI7hVGiD4MK8pdb//3LfSe6dgXn
z7soFOfE2DL+xvLdjz6HPW475P6cFf6PjUUR0vClNiIZhMxE1icjP7REAMAk1rsZJtovpNUoduYr
ipDQ0XwKmyDu3/Bx4KmHcc8JjxM9LTm8a1zNqWI40WGXWENCf+BzGvIamsLa1qq/yQFIk9H6H/1Y
nQXbwQZ8g88HTgJZOLeQmCzrAB/YDlXDzkBoi+MktZ/1h2Gtrd9zn5GxfNc573vPrGOXS7L9X5d7
4NCxGuOLYyDhMXX4MrUiiLPjBWs5Hpto3Oa0cU4vz/UWFcQE3SLkdQHr9PlTo7rT9bLpUgv/q2AY
SyEzXMSWGVgZ99BB+KgUJWDf6DxLb3UkJEiFoF648+vnK8iqtCfCRSJtAa0HX4Nc+8AnXmPEVPg9
neQdf9FbXXvncRBCwsX7vAgl14pOiZSv0eJNlytAJe4AAtBBoTdbSnM3ggX1dJM1vNt+2RzZ6Aqd
mgfSN+Gd2d1OQhsJiWvm9jke3gOWyXPnINLFwsG2qWBVsBT6vKWbvaoNWuF4zoK4I6aWxygBdZ5t
mLQQdVg1+zdKOEggJmYN93/tnN0V8KWj+4O7XjwylvT3EgwvkaHHvrnRcVdJ0N+mEle7xxB3PHFN
/BJVrahISSf+Dq+JOcFr2KjENJV2DmxA6nqhbZ7Qfpy8V/Q3FPrQdxXc6W7hXGKlyZ1YMbbgqif7
j5qHIyoSacViErdahT5nCVOt4Sek+t5fzjo5DPS9uA6iSGd8sKgv8jDJ1/rOrtiTEKs0UcWOvs0p
KrAT4TxfDn8TzK9dCRo2DW04LV2Xfuw0wyK1SspTyi8i434+jZm2jzkuTZRJOqbT4KOqSChjTci9
5jG1G02gafrDXCYMt/3sZeLAcnYAUlH+jJjOnOoe07YR7J0bVPn/zF0I2uFof/AZaWiLfMMDzcsl
WAu2i02YGEMVHmXeJCxPwKOCoXHtrIxLp6NK5YtrNFRevgwkDXrxWOPNeCqcseZVPjaqjSnp3W55
gkibgofR5gMXENeO4tiZqhdyH1vPv3yVlWnsuSIOWtMoEGX21rAmUuEgEUsGtSkY/8PjPditYScO
tRI1ptxvq+6PkQnvFkaODIBSw8/WaVUC1+zP6Yl6ZhmI9GbXcoryIS3NGa3RgoqgscpSX1kNIoBy
zuNI1Ju+xCHRSxHHLcFqGgMd5tE15v2QxOdeoVn/WjPnmdm0D0q2X53DFUMDt0XQWNG3Nn+l/Tgz
39BmAuSU0aDdtRsmNdIAJ7iumh0AufzXAji+/TdzaBVIZGlUcXMEEpHuf0pVaCs0Ym9y+CVib3Fz
71WBaTflJoaVHyln7t0PzvYGRzrR36J8KoqZvvdewX/WWljCgAbu4e6Bxn84VGIsRwn5pmB1mDXo
4V+d95a9DAssWFCaPHJUmvyY166G8GZzVVdjAaZ4q71tAX+xPtWYBdQD39rCUpp/lEAx+Q4CzXQx
+U/HvNBADiWvi3e9jjFzE4vRRL2PGxJL2hAptAT47YgB3YYwAzb7LgVNsmYey7WjrU9ruAS9yFHz
3kfZWfeDO7gQ8zblxx4JSu+v4PSP6GFoIK3X7RpUH8rqST+wWDPwlVxmgUnW80CXrF6qgAAljmDO
8SLbfkr9PKVukJfY3u2m5ncXBoyQLKzCl3fyiuQBi3sAhm05yGpDghg3Uk1gLFPGPK5wm+imvDnY
PfrftWEWKgm/27D+fRycTG3Lpop9aKfMkLc+55ep9PiwBfcewfLH2bs0TDmAXrSoXbjr52yBlqX+
e8Ri/GmPJRVi+a5ch+VLvr8gqpCNneHDEXBs+kqm6tWax4IinXP8tX4VlMO8sRk+5Mt7Tdu4LTjD
cYP8jlJ7G4x+IEAq9qq6ghUprgpIL/NqDf3expYmiZWj/+ApZ4hC9QXnklVUieQUN/6/lvfMLzM6
E7LBkj0rOKiWrBs3E4quQEMrLO8QzavuSWEY59SkFmCdN6FYLj7bNxGY8D6V5yvFgWhWf+tSTxPq
DKvuMWqatUZGjA7oLViJLaX6HuucG+dE6eQkSCnE+1GXcYYoG06/M7DOHW+Vlc3CcAPMHUVd6fg9
zz9j3Kpjj1vg4+8mJ4PZiwUekNCfCauuVYVZSnKfsTcFK9QXziXC/kZ9fBEngGDiWxiXWituVbjJ
n0YYsGglHyJlozH/kBF3YToGpd7YC9Xf/Qd4P37KNYuxCecF5KzKMVzF/7t5afUZJC1LWIP33ixi
j4e6f3zEigDZqUS7yJdlJPKaELMWhtMSwcjsspXV+kMU1PaxiZIv6PZ7jKPkrVIXdfBx77eQYeb/
d1U3I0xBe15k61YT6cmFydQNAtdsWjvzz6wh2V3nLd4sj5Wpaw2tyQQ6hnkdz406Cf/JRPRPPHl8
NjJb3B0Ad76Zzb4L2AoCHT9ZMaLCaEyzUf08je5nUrmWNHrOr3BsZvMfPwPIpnepg6rdtJKX4GN5
MoilBnCsM/5a2dkQYJSyPmZ73cMsSFWFK2YYPRMg1jRgWKd5+T+5VfVbJN/vmTPQv2CWWzMVYctN
IIMURZ3d2ORA5FAVTGro47OFKgS37MCgcqAFYBlGZmMf6nTosksooHeLdC6v8A6/IYJhrrL3x5JZ
/+OuCRGbv7RdIy1ltF6NSEw3SNDm7TLoEWd35wd1DVONjIEkVV7Adw30hA8N0JdU2sQni95Pfkio
lbkOa0zfHMXyjD4nWk0tfSz3MerDFZ/cY7BWAq0gzOuGgv7t8t+1MimhS0YNIaqXpjKTwSAmxDsu
zQSJByIkdeGAxlthVE257v0BDryBJx0aRkdMDszIKRk4UfFDzIsreCGWn/ngBpDYYh/M5TlGYiZF
zKcD6Aqd6Ts1EZL3VqECcxnsn4JzsKkULSSJhTTfI/oPK/pyuP9cYcACPhSVSr5GjF+Q2Ob9Nf8O
xu0HDCQcVt4YKA7cESwgAQkwvpVPxue1IlXGAGFewMUxxoCym71qMUdAguZ3L9Y7L8UYtkEkDr6E
jNclxqLMmd3lzwf49RURI344gvXLrzrvz9r27j7A8HaRhz+QiErll2+9V5JzB+Jgs+yS5PmgDEyx
I2V6XIJzIwFo9BCjTVa3ZDhbJgyf1GJKd4LhLySCCoeQ8AWeBnwDKa9fNVuN2p4gyoqQeNs5UxIc
lNg5OHnRJUdSAwAapVs6CfeJdAGPPzKzEeXkOjZy5dP6+5HLuqXyRSfIQlRf8zkov2CqmL/OIq7j
hLmrtH7latRDjGroXyO42WTqDducW22rMVIm2ZSKAL/j10IAmSKVAozYCxW7o+VSRtXcr9Z1tbSg
1PE5+sYq3NxnQB/zw6848FzS9qeVm4LGmwsBGN07+1AnOvFOqSbMdEBNWTPuzRuTVTPf9BzDys/2
VZHAW+lQvAkObKPlrX2V5DYHXGHUl3bsxtPIjMRN3H2sRDfQcShwvRzSfBQAQ/2k2zWxY7JH7E/6
m7tqKDm7Wc+BuPW26yVr+HCnZO0UczFLQpU+9lemWNlrzsj8hXE+Mijw8JuJ4tMiIHU8gFH+Kxym
6PQtOAJDfYjwbcBp9yM3nTWpLun+rWLCwYi9ZhzgT1pR0Q8CeA8IOqRkytjHYYsIV6Mb4Zjw+Nzl
FY3wrKxPyYCyUBEwL/PAQMvVq1JLqrAm/aFad57kE374QKvdBJ67K7grFOYR2hQYEDgaTWdDgJC0
6jc++bYG0X1XjwYtLgsf2JR+uNBY9g3BeIX9ImgdJeix/+Zsigf21n8r7P511CxUMzokogXXPv/3
lUZWVbdzfM6UWMi4Xclam0Gb+yinSxjXdXTRSfnP3VlZd4NThwyk1ZZ8DNfETkx9+nIuR/qcZaDa
pUrvfO7sm72nTCdlv7vAQG8u5bDlvApyLfgJBmDvckBTt3Qwp/7P4NMQKvQlMihUjju2b4QSnEzw
VNRvOyJzfXSxTKcQLSrulzIPMLIIvy/62kP1jCscJr2t/L1T5vQQzP8zem8J2SpFCW42A+1lRabz
e4PtWANJUWEJL5odT7r6rhQzAU1CRgpZCm9TEwjO/aY4UF5SlxZpLIk45vBbFdekaHZ9jVfjbcl2
+qmckJ4ar/fGXzKbG58+A+GiYKx4NN3I0P8Z0yaIQv/ODK65NFn8y/p7q2ZezNm1aNyFLdbwJto2
dl+LIx0XiDzAXRfckm7QNeXIkDmxyGVg7hRTuaLvb/dYlRpUfIPFOXzFkFax3HIcPwKROPoecWnc
BfAAJezks32FtdYJk+oMsKuP2iOocXyWM/GKcWwUhDs9Jc+B9T2ICSg1X85/t5yklADPn+d3d5sv
G82mHwrAz6IRrsV3jz0ZTSBSs4oN49bJVe4OXxDJo8CDoMHwUANGZL/cXRgtzVaZyh6dMw+qEHMl
MFVJYUSr+/i/rorzn5jdDKSLQZTvDHLBKpazjAbVHGMRq069ukHSWh/RI44U2mlVR4xCekGk5KAJ
qEYcPd3cI8XTy6znPC36KruEkkTfeJjDeVyz7DGULxZF0Dy9wxy2tzJz2Et7uVIMcoI8tHJGso+g
wVopsvtDtcJp2RCX9pgroYPyFcLO5+xUkyDvNKhfdUsN0+F4HQqbYv0Yys2LR4KUIKuwnI7JSIYw
HNow9ZNn71k7yD/vn7Utx8ZOZ79oXID5mU4Va8U5MehRjdngw5zWdQDj5rO4uAfJ0E6FjOHg9UqS
AD5uWgsaJoUVAbnQEq2dL3FCg0SrJKJXir89F4Y5SHcRlUTl0i1tC46OhPwKpoHTzzYA1oCI08TG
3YhbtcJQ1qg8bjz6pwe7pp/b452TaTSLMsfPvpUwNlge2DhDQ3PGmu2nqyyFHEaAN8sr4B7T4ong
DSZIQVeMwzbePIMTIvNqUwHB7/ZGAlx9tO8we9O5wesl1ldou51tDfAN99LUvJ94mR1VCTI6/AyN
Exqo6/16gpiqSZkuqdZNhLEunAgZ+cCNy8ZW7yLrsuIBa0Um+Wjh4xpV1rwc85evuDxteLNrvydo
Kp3uj4D05Og+DQ7Gg55TWZWgns3fclsCvymu9TS3laXpJRu2inPHU5suQBhYi7Iase8XDFQqYfKN
9g7+bRWjTxpV/x9N7rLS82S42iIFHCYifpU99N/96qarF5gg8tAx8KyVtmFtfGd92KuIe7WTQlY/
jUsZu4WI/RSZ2E8CqPG+6le3Oq2uwCSa4RnyA14pyOTQtXPqwqMlfzKWdcgGeeGuow3avneTwCnK
OtdT5II51ESxbG2VZXEjvcd6ncJThr+Npodnvdz6uTsanDKHQBmrJQbUo5MS+15nduwp6tbs+Zkn
twqrfnW2sUNbtGN4stpV7U7z67rYE4WhLL1WhYpKgs1mZExo+yVpBQbPh2LuKPL6CCE73koEjax7
RbaB61d1YC/dhIQy3kqHEKElMXk9Qn16aTq5F4e0SYjYc4vncRbgPhCz46L9sVB654SoTbcLZfxn
xG6W/Dl4cpjhS7ugkvtYkORIbBb5yhTSway06iq+oj8edBl4aDd8BGmjar5kTp22wbILF4yVQU3X
t+/SROGMhdOGhFxuFeYS7QJsK1RWQpFfbXiv5cE6PQpEnrIHhOmbT05SG95sX4Djlmym30hTU9p4
4EAGrdrrg2GZvt55Cotc+M9HpsqxJrxs28mBGGXZcfVjPo8SXI0bi1LEuImZT4PH3E+zef7UDWaP
SO88CzUha7ClOirx2RJdtkoUyRUhI5UR8aVjy+1hyHq4PY8IeUmJfljMw0MApcYX9u9bm8cp/eb6
DIY47i+zymy8QpMQ7a0uNMiWTWQsUvOirzXJJMUUgA6Dgr/KEY5Ofm48zWE5HZuR52av8SOBZ26g
erf2vzlX6GedvuNxue7RM2WV0WiP5um1avhlembZpphl+H7tTUv+Z20ZNMS5bIlqNyXfUCj6l7zZ
BLQX38JIk0okD5vWob0TDQ51t3M7rY7bt3bD/8VHfQiTjFsS1XOR37Mo9Ud1RUgahg1QY42lCfW3
AaymVKMuNWT8PWQbtdiu4K2aylTV1hmohnc6S80mrvyjjcaKIEcDqSiQAz2WiX+UzPNQffCelCOj
QMPir6KoYSsJjUDkSb8iRvG5/tRENMvOMAjBXCwUb1lhghsfWkdojRl+en1rS0T6U5dSB7ccPzI8
/bIHPQNx/R8aORSuWLjZkSZvhi1VqkQcYQWiYZFXk2yZObxtLLbgtpRWOIiyEdVedLe00qBWMkQT
ixGFGaRjI2e3dtKxD78Z5Aa/Y6yZ7DlxQOUgbzUWjvnIc92zapqoVqAjyogjjNNO8Kttz6oZta52
ie9cGUbto5M5vpGy22lC2ebqk+a+y7v9Mf8kWzlz9m3LiOH01IA4Yag/mXfYxEWed0n6p/MDWvAb
L4MBIA7X23V/837Q/6DkoIBVVWjVgTQth2J/kq5d8XmMDvzh5JBVg7dG85tbCUGRd+mmxkwByaAK
jAk3nys1W1z9hDt1cWB4dwJ8S4mjsN3347sDA3hK2ITQ496VaZifS9FdZfkvdQ07ZwSEPzt8Omtg
WCrE1+QJZ6u5cq0u7KwED9RDgIRPUMxJKTBURy3pMS3hz37Ymgyx783l4EwzTX1iyS91v2mMVpPX
5/xEFvfdCm+ZiPCQJtiL3uiIscqBo807dziSltxgasKlrsPzNeDGWTcQvVl61E+r6E7O4UBwzMte
6kWGKs4UlJi/HBa4WiuuocqfnbAbxlKT0xD+wveXHDu9Gwmmo9DNwojoCNU7J/MdWTniqPKIEBpw
Zg6PPgoJtNveWCfBd+uqO+Yc5cNDyD/Fv+CFT60CRqESGmmmLhOzezuzNP9vMOwGzTbnucMkCAIo
EwkHiatNs4yXjXBrNk4xphrbtyotFEHCgFzeu+Ki4uI9Ui1PsbP7RIfA5jlsmYCqzLdpQ719gyeQ
EwMtAtqvCa4D4wYa01GdqlvLAo7NSkxI4f4UZiMtF59oezstToUvbORLhlRSUJ7FL13mrergbGbb
fHxjhIIkZcR2JG/ftwVbw8zaerk8lLlb0t0Djj/7/ZUkdWs72+0DZyq0nFKVWhElqs4jY9noPtzV
vUtuzimTnumR7owhj/9kCDmIHJxQl5QfEHbfyBwl6zENySQATemgODkpgbNlJIh/AY8jrqY6y2iN
pHNc3FOgcNHBs8/LXCQrtVQlEfB3F6GoewYR0RAsS9JORMtWrPDXG+263LFXjEv+PLjenW0Kn88b
qJyBEyagp5PUZFotcU4LNmmMRYqym8cIHs9jMoYJH7leHmTK0ITQJ++UJgvO0Oi6trormwhJeGJw
BwHL5UGyHZPjuwFWA8ciDQwyNpCo5dm340tAEXSfyygmuqu+0UkYiIbzY/WAs2u04UHastHO01tT
ldkjusD508E1yet8WcFH7iqpbImDpqSoXBDkUZjZQn6oylc9yvgFi4WgxHYWmxXo4pp0G2lpAz6H
vISibh/lvMEoZ8ipAfpM3hk2i4Z6pRBRBwdomnRA7mYtPpLaFcuNA9ScLsF2MRkI75QPcDVGq50j
DwkUA3n+d40d1c9ImXaz76tnjDLRqCzxFvG6kwey+GzjDOUM/8MJzhW2PuH3NdZMTZa3vbXI/ASb
YJbDflfYUBzKa49GEs2BiBQeLfnaJjp1gIJZ0hVaW2osnXPKZmGq027mogH8ljPwkGKjl+oRIBaa
Lm2wrfpUfvLpiRmfaWmTZAm5YIvuTeVfGru+8iZcf/0Z+p3z3sCP5cII1TQzgPKymEeCqpV1S5MU
P76t5gNWIV1N6VfdrvhyR7Op3b9WByO98KZcG2k8SK7h7j+3pRDQAJq6LvJEKSX4F05x4J04/oJ7
zTyVNnsn6WWGE9jsARWaSt+LyvpJokn6UxRjGVPS35uYAhCBKs4WG3FIJUNMoQooNGVZlPK28q2p
HEl6tB3Rw+IS/d5y/e31+3lX2BNKODp9OjFzT9RtEGh+QRIGp+pe9yBcuChrWsD3twuONi1LztFx
/66OkwKEhBr3jmnMBQcDjUaTTc0xmPxcPqgzSTchqSggT1rIc5IFWrxblztx8DBAF+H2S/dn7H1B
RDdg3c9Wcw1DS1IXFZS5e5FzjgRXO640Z85+EMlfN2yeMRhe8E998KvgPzidE+7RMsSUgXRxc1Eu
b9lvdNmsSv7XwEMCXo2j/2rF04vA6IvWX5Q/s+OM1OFRU8eN3j5zHOxmGflXJF4UPphFRnyCnMWi
VnOtUeNO16v8iBk2Xe/WHWqws1Uq674uN5odUDaEdoK/dCFeDy6g5e4X+rob240PV41fmt1MujJx
qglCj6Y6FQgd+1PtXXX4bkW66szGsJEYvPInabi1lq2ZorK0WCm51Mr+8XYGyEQ4slHI3u0jiW7D
IqZ4XqCVuRwYRYcnVhT1DKcFqKJGg0S5j3w5xXRrZckxZoWMYUtZ7MTv5jTitJCyo7lrTRMbuTPZ
RsFBmoQQSwBwiHAJrdprm+8U+pvztw/lTe9GfbI5xAoOAUTmXhUQVYxCX9nJoBtGl18Bwsuzbhb5
NyiuyiqBfPRDThdvxSUHGH35kCc0HhSj9vInGBxY35zwrFjoI3QWZGa1SeXmVEVWYGty/H4nKs/3
9aG7DCnr17NhwGYbBC4yDu9QNYzxtxa2i3FY9G12abrAvFsEUTMP7kcw9U3yMLX/odp1ECDusBPZ
6HrDwaB88eaeH06x8fOUyccQVBi4iAxtZWpCXSuNFL3oBGpsk4yIw90/wQBmp7S33HJagQrpJK9+
A/292lh+sk6VvCj+8ECmMSLFKAuFyZ/NkAP5jLpau1+zov1CHFd36bTxnmddFjxEj8XX5weulVAJ
7lcB4HhKIHv1BLueADq8l5REXpdFSqrk5UhyHk/46pKoOcrYbiGjYzvFX0sk4HJkXNI59mH8246s
UBmACr2alyuQdmOylSpAIOO52h47Va+eQ5iBfDlxNQwYh4OcVboMK9SvycmPmEBdJ66y1Mv62+X5
VYecqqi4dM0UKqXUkfVlWPy/TJsKPRwoAumPfIcylfWpeYd9rDIRY97a0ZDl0wj4whCEg4BbaNHW
ZT7jes+bLDgXz8Wz/VYWgmHR8lyggn2wBEpwfVDZSexiIZqalcuC/KiWVju+i1QqoytQl5vscDzI
TzD+p0m25Vgz8vGlJTtIs4Lr8m6rhwTz5VDotU8ga2T3FzYNPh4teH9LN79BPzGk6n4I5q/UD7GD
c5h+/7PbmGLI2eb652s6ai3d/dmxDrkmuiqfKVUZ14P9Z21qzCbTjKVBd3jCkgXRmmwdphB3QZhj
c1/9pbx7prSJsDpZlQ+T9MGVvlKTXtfAg6Ydd9G6o3cujkzasnZenPOlpaS8+i5o0vLtMoLu1t/e
ktlmfn5Ora/tcw26ysycb7927ULE6xQyyIaka/nP+kmv1dw+GPhQWFYToS4lRl1O+bn2PkcwnWzd
oD3jtt9TaeRjMJE86piY+5TI70ADz6dnP1dkN16enE6txgFS2CEQ4yPAH+7zmUEcT/KPIytr9VJd
BiuehkTsAQrYGVoykgtEwpBRZJpECHdEqnShIEUATFV7HlYyZsTZFPp6M70ad6o9ireD/5eSTHQ5
86bBNQmIlFsM7sZUcQ2HZ3+kGqjNol0/Dkg89g7DVwXB7Kve9cb/LtW/BbhvqkAIaAUkWL5cwEXV
Fw+Tf31AqZR67ichkee5ILaXyeAB65ayicXBlaXH8txbvEQVihjWAVz5/vS6midLUjMEjBxjKKnF
WuJ/S6mn/5DKKrmbm4fqYhlhtO5ISVY+WMORS8dLevWty7j9+RhqaWr9QTbdEkDywHqFcr6eroHY
lMINl48GhMQee6yMB+9pSyAt3OPb0S58/tdECJQiN41kZzHYcw+io1CohO89TEDpOltqKF1uOXEZ
L1HLT2bk65nDTsauj+APayTqW/z7uo26/I3Jw4G6P2MTIa3QwZc5QwqZx4QV8hzYPeZPBR50eiHT
QBEdjFZfjTlqb5y/OS6+ZM7LzkllipG6wpoGv3WoX7x0npOdOKLwL6OZ+pHegjPx3sVuSaKLtIuV
BWgATzTpDLZF4NPJ16Z2pBLJEWtZv5RQQ/MQsYEQhgiTzJt9DyK6NCtskgaj4U7Sk/H9Gb4+YUIF
md8/yVQNexMDUJdeuG9J4xRmR5LlWWY+gnpkOM0Y1EpmGI25Xzi/pLWu8Cu+Gq6TP5zvoYXFLNnR
MX0Q04cwA1Ytg/qch5kuO3SbVhARzdsVPxnRV54fabY61Wp4zSLSX7YHXE2FiZGILn2a0Gl/M1hi
6wWlYXsyK8hSskQ9HD+mRf39yMptFLcJalXVLOhBPydqnbT+9Rl7ZZ8sY5XJ5wlHLI68UZYCyZRd
/oPPnXypqhpKmnx6hjINSQ0BGsEjL4zwrnAWlI7TneolZ12waUHewqRk0geYyOeOwz3VJy1n33hV
8a44wYeUGdONmeEvDRDdGoCZwkjM//Oyvn5Z4jVhRGD1tXXyNZ3mqlybe0TGssHWMR3Vf4ATKv+B
nBF/XS4Tb1QPbGR6jjEGq1aAT1hNp9ZygnZKyGZyeU0cvmPkeOiXiXcNYQsEqLYakTeMudxojOYs
Xm5bRMpEz2V5Mnp6h/T6OJKTMZjMeO9Q/FbACEFIM0d5kv3ezUQ2ZiddpWbsGZtmQ8R8fcSJuWH7
WLAN5KjLmz10ocS81N0XuqGBgbNEbGoVLHQkczvMBt82BW59kpWjBtLdHcnaMOtXsTezFydpfwMw
AKz93QZntuaRurtH63j/y0CQ0sV6WRSjrcv5YRTX2g/VWVFOCeuXAmK5NvqUrvRGXRBGgNaHT6HP
avnVzblDEhOu+SxBf+CbrDUvXyfUvQALIwCuGthtH0mESW0x1KX+OYKQ5XT1kNGYQkwxwwl5otkc
vqSpYkGo0zWlAlRgr410kSksdTg6hHCu5S6bWXolea6Jk9LKQVx0gBYaKi6g1TkAOTb0FuB57Anp
AuL1gSxfRfUWGeNvwrPZttT/lzqq2WtccEyF0wHdIU5E/htelRW2x6/5s64265AIfJJ9P1NjveEb
k1vKINJy4QbprgwpWQyfp8d/khM21wSbBcHWsK8Dz6mNWPkHYR+JUsXDRbePxCNllOUdM64wk+7Q
Kdi+xvYVi9i4TRZqmFTaI/ZQYTa3uKUsK+ad+FRMa7/A2Jz8pvZnVvYpj+vprgTgL0sSEcg58z0G
yt6gHkgQvNAHeipsDtUgfWivNIvP6MuPuB3FJTU2j3duUC0ZW4w8DVGk42NrzppTx6n8TrnRSr2/
Nvv0Er02CUdYGkoMnIqMW35VS7Xrd2stezhs4V1E7+umDXHacOrjt2XkwXaEa3PhkTnuBTb76vdp
3jDljm8PUyOyfYQSqwQ7Vp8U87Dou1F9TpsSR3rra+FmuSX8S70rFUq2lB2bau1MT7wpX+jLF43h
K1cp9fLczjVVQsSEOETZr7BeqcIKBXlsiRlfKjPb1gph3lYdRCWLd+smXNGw3i/IMbOz5t1skBQV
RKi3t2uaD2c/idlSeSKMDaFzrdgNa/tQcJeSYHT703ZcObLIGWJbe0BuIdHSpVoMOTFe9wJLUNqJ
CYBQZEI5Ae+1unnUHm2mIastPTz5Fj9P/zGwx33FNX8U6soSe9O+xNujYwgaXnF6mjYMqBvcTU1s
DEBpo0L4G7qQLSg+FZvbXC4Q1HF02diw3dIiR4RQGP7X/HQHSE3tVds1oU9CK3CT4eTgxgatfkcd
4edvaOT1z5QhYd71vkzPJye44QQjeMHAL/XRWYOMmYQOldTTKa+jIjGY0QyeNaDd6nzM0PgIBhEG
iigT3l68yATCF0nSJVoZhUQLL6PORnKFI++aj7SphFeV3tNVPugyjHYBAc2t4ZySK5fj4oV1qyYP
SQZwOc6qAgp1wP0BOTN5Po1vnww1+1kVdeExp/rwQgSifxiAICi7IqHirn+Jt/tlVSvKtB5W1t12
JfNPXeeLhZVryLP51R2v3Fe3b2x0tFgXk9Ip9QvIAy2u2f2jeFiOyrWdEqBS8296vZJxTqfA7jT8
7qYhrC8OF6m7BTqZNaij2dy/K+UcfgaFaIFZOI68tyUDIdKzZIDP5tjIxcdtrGgAcyq8pxxQqJ82
Llw9KHdgaSPEn+4CN2DVnVMzt01ObQO1V6QaesFjINHNgiizsjHEDMRVb8YJG1ezNVsl6b6oB1N9
YoOrdkeTuv3ap81f5fDXozx1pIS8ul5UPJy1qa1oQl0/Jt8xO/zkztrMCyh6AExoiQKcJtyi1N8Q
UZHrKoqvWyX9SLgkl46M/9yRkQ0Gke6SSrknJzG96NSF+0TLkTd9EtdnSn8foFn/fXFM5wpmlLxX
/XjzImf6BvFEufFwhqhseHfLW7H3LLovjyW46cDjWslrjGNdWWlIBGMjpK3AHMT/Ugtsth6GSANc
A6Byl1+VsPZCrF2yCFyAX0c7hkP4nP2XeN/xMP1hb0AbCK2h6+Oq97sOLyNsz+TzzCKDbHSiDY5e
zwg85diD9bU6F56EddwxY9pFUiu8JdGgKilbp5xqyucBr1eamfKSEphcq7aXgNL/uTuRz7phCmR9
hb0pi882S9GlMOfI+F0UqxsBHYq5EUWcI1VpvNB+re/DDlmVmn1bDrPis2TwahhYo5RqhWzWP4Tp
IrP+D8b9KY6Ql3yQHHzr1qeno94xphzu7+JQNBDhbmZHKpu+VwzFP61kvfm0GqcwAbvy4QkVaE1w
XlzY2N/S9LJWjpSMppQ5lkyJ064juNc60sowLOwJoMDaOcrEP8P+YDm45hlW1KVzUvHKakcQnGWL
BvjY0dnxLRwVTQDfeXLYHSDruHIAwSjBsMPO3MxqCuk6ydwwOuNLJzPATQ6ZFZBKc4I4TX/G0fVW
LrXY/MdkJHc/J+Bf4vBYOwnjwuid3BdWcKzx8/Zdfbs+Rnqkx87o8utc47zGbdKjug3YdyuMeTYH
0Li+zJyX6J39bxEwzm7rrWnBHT84hJoTku+gHK0r6yvd9oxiuHty9g/7PnxpXIsJrb9SkqyWtyEc
Rw2Jv7sgHc9SxjLbymjMptJ4uw25uAMJ04q5FYDPY/MWI7KEz+ifbO9VSyn+ivKjAYWIoV6ycua3
pIAeqHu0d+tgzGDY8vlDRkQ3pezDNK/3tUOL9JBbCZzjnzmtWvqXG1ytiPKAO1LcVnz8g5YKKanL
wWUuS+EqmHb1c9oz7G9qFWQ22SuqsYcYk/JdrDKq8BbGJmBbswUtAP5slEN/mCoWbzvbbvjZnXHs
OtyR6GzEB9iDjYlyyiQ4stasW+escHY3MJ5qukYX57bcBTkoWadnj1sa9kw8i8gWOsF9g/il5oat
5EVyRieakycLGr8ol8cQx4Oiuvg0aJTr9kWbY9O0WNUU6ht+ldutpYWOYGi1It8eZAHfIPkB85st
xZRg93kHfTsn3xdpXBqb9xgLCzgwWDu7T+KMQ/PUywIMTLpnf4taP2a8cNWsMtp/l7vL/Km3ilwD
JVy+r0JpvaxuoiGUGBAnrWPXLaDQhFhuDvUM5unus6zdMbztE/WUqQXVBo3pWQ3wPQX99hqEeZpw
cd+WNOKKNwd0pkwa3pW2xOBYUcnYQoAaitmddl6jclOCSOGWMYjdL+/9/2HWExcW1PsKnNIRG7f6
eDSCznkDG++HXo5pj96tmBWP+OMws1c5Ke0cSs6Tv5NV7SwSVkWHapA/rsm4Q2WUzGhfQbbGxamH
Qy4k5k7TYooA10wurFobSC2IUtdSpOtnnP+c1lPV4TrA9Pkis85lQao2uYrLQSfAJ9BBReiel4/L
EB5V+yDqLDtsV1RgpQIQ8fOBrhDCxJLQA9WWW13iat/PddIwY7FMPYG5jXmkAmA7kL4SNVjKouDO
2PpFqnUtI9DVG9eY6XWFVIS7rdB9vFQ0xN1pkX438PaxIbXFXhOwC6qShXJ3R9ZV87r7IFVEvvet
4DO+sgyrsTq97he16Cgk6LnK4OFPnaFhlqwRZlE/ecaHVGSjyTb6tZZuk+oi6bAX2IoMHGGnX7NQ
7b6gf7HuCRJqKYKm2v/EaA9/g9IdFDLtVrdM5J/szW1G1CSCdGRDaVDAdxfwE87TAl+N5oxws6hs
+ZNoXE3TPAjfafGYIhJYc8joL7J3v5s+mpYvQXd5v6D0vN/643XCg1iDkrVN4l1WVUk6NIOd1Q+X
kQeXxkTj0YWX0fYhPXNut/l9uQTxXq9ZjbO5OywsMPTOR0NbjnuyywixgdR0G/jsjtZ+eXCkcEs6
ADZsJn3HeUotBQlmz+GALYj8IOgkXI+8H+Owmo+34ZrAng01JNuoQ74Ukh8R70sg+52YqKKJ9683
6BqRt4ZwBF9wdIsKyo+Q0ZiFePOQOmW3ixg9reKI4tmQPo50HQDkuM7cgaBP3eAx2DtQprUrIrX0
twfoDsKUQGOmkqAuUd98/Ze/ECPRcNkWCJ+0QU7OOe+TqkVvvmmzqpUVo5+P9+TFh+xfRJwVF6xs
sAgkyPGrYxj3VBtLApeLdv9t5oUJc6cjGeOfPeAeXbMih2iuZaA6XTqKT0yNJHPRinpPPQSPi92H
BHHFcCkkkrzACEFmeiE7TtzGkcH+DkYYdBZFFgImMvcmpCW2SWjcJryOPlcu0cS8iZhHAVm0kMIC
2Zah+UCMHFEKrqvFhRMU+Ad7EF3xMVgPJB/l97PX2L36istky2jgOJEEzzYP9fv2EfcC/TgbLdBs
zr2jCgztNYnCaoockzX3FFPV0MKiio1dv8q0FP5GIgVvJPPvgRqjKYDc3WRgzXi/6DXBBsED+dQw
kCPVFbPobtnBp0qENYrXHqxqSJxOvRWp1YDJFRLQsd4I8Is+UeyaRc0pSvDeO7TM3Ll4Npq6b/Ok
jkDAranHuYC+n8Djqsef7Ya0QmLF7RQZ19XOMI8HVGXjolOaNQgyHaO1bx/MENgs1hx3wDrSmfFl
L12itt1q2G3B764yeO9Uu2wXZYowIkuPxMEoaId4MHR3gnjB4eekI5Hla0JyghPGWgYradY65325
DjANaTa6G1Ka/v1F3kNMhph5RMcExhqp3To+DeCAVfAdK3wkFufTWJpWv5ogqsbwGy9DA3f9DcTg
RNw71ty5A3zXaqsL+JihzZfa5XhKAFAhomNwQs2HOploHrIe0l6ih3Yk1FskgdQMBXnflCJNdVac
1vvkBGPtlB44Lp8vM/2T4J7lqakEF0umgz5ydBmq2JYbdORBEmAZIaGZWjQhvkCoJC/HAYFJ7hyf
eu5ARfpbVFAbeYEJzmXwBogn7iOffCWh/N7ghh8IHE9iSF8LrFT6m6rOvZbqNEccAUT44JeOSog1
2ecANOFyMhpCv1ZjNk+NX2Maa7kvTyJcSDsTm78yjRRUihfqkw2bu+VomijexJWA8AGzyT6QB9+5
xF9ott7f4mTHJZ40rvzamVZzLdreBnYW4p63XxcQmToeBQ+MdKmuaj5rNmhrhXhvRVaE3NaWF3zM
RtIIDQaoLlbRSTszQ8UWUmBsBMW/Q1SIghp7PGoXRgwUlX54AwKzUBipms9Ys9jbPzgTo/BomYcS
Lk8nWHWCXvCqeu9ElKSgDQXc+Q0FfWaSPwtQ6bOVjP15bU2rHvg88keEEdXol7zuNPd9BNwm5ofu
PyvaJGiEP1UTFChTr3aKyoDmeEyCxL8L7A7unMR/xetb7i8v4XUVJn0Gy+TEP39ugRN9pfVykzMj
yall+qvfinzR0yHv+KbVfENvqE1YOQUxffFQlTPJVinq6YylyAZMoUgQRu6+b8GVu3tK1TK+DgXx
INMFdYcU+Evr3nzus5BSV6R+yWLVNzQXQ+IIFxiP3DQMJXvRgI7e3xgNbIp/Bx44fEHcMrvG5ijc
Dr6Nc/FaGOQuqnu8pMzwJ/Axjq4x/Lv+yQO5PEVPKp5fUn51T71R8zUnufbPEfT8+gHNZyCsATIc
oyZqjuZdEPiz9NU6W+BY2296AuuWRkwWFJgbc5qfN88bdbEOVHoP8jRunRk4s3I5axA6jgcW6U6Q
czlnJW6lkSxL2N02SaNenlu34VYzh8M35swAnheKRq0deEmKXeaaE+eoICMD9m5/d0GXrt8Siqof
4d0wDcUP2d2KeTNl55xxAfc+KHSK9uyTJHXmM6WPrmk3aprtXD6anjeuDR1C/gjj4r53lCPpIOkx
Etb6+v6sTxDHTYlpIHXrftfqvN2Gs2w0q+8lRg3fskfJR4AG7jf5K+e1uc9UPtlcekQUjvyjgkJX
9Mtt3DhC7PPc0ahm9i+TSGy5LrzFZ8p0/dklE8EUtHZFafDjigkV+tu7MMkQDwlfLt4G93YBM0tZ
JQSLaNu3zPmd+HjxkpUI43W5kuOgyEZR1qLrb8466z0DfF1vYtwWWpj6O7zaivvUUW8ofwrvWa5G
IDerNuJZ90Ctg95ewgpI6IzOqa7saU19U9+leuNS+d4MfjAm44vhyu5GZh+UruZn8wILP65BKda1
uM5lra/FKWXCy/uMhiZ8T/1Y84x+m3mqzgYjS+ISr2VSlQwv9I+wfA0tcJ+gznSDjhZLw+49L7q6
ImW/hcl//NfLRnFxuVG0zEWlBUMw8Tx5RRzj1N9IHs3aUxiY3qn9ZABcM71gMCtXFfJxwDDZAoI1
SaAWeTL3A/NAHnol06XQii4BB3xN5AfXbqgYEzjA+vLax92ts86lMYQIITZKN1LOPdEdhraRSO7C
XIb/5wQ05jj7e3LBTbHqIre6OHdcHXHCQzC3K+K8VBu4svk8oAxAA/3m2ME2je6ga2BtJnjJfxeb
PhYxzd062TouhHvUpsITWMa7GQ5NFL2Iq60x3LGURQZ6yRDbuLEwH7algtCGWHpnByM/Wzn7+9Wb
1Wr6KXulK4n0ZIcztpVDOQeRUG8SfpffFYLYJUVhRfA9WrdN6NxJEZmlxX2uq6QnqIDRXlLr4IEf
oF++BPtiO2uHdtmEIuMNuk/+liGLy9wiLw0TJftmZre1C0cQ3CcZwB3IK6ppq1GpgaaoeneE6B7g
vwf0XxdpN0yIm2560vJcuvEuBQfsn5LnSFLF7sg1dd2tjmAmbLaauBooxvMqPlqNlOOZF4GUPZf2
/owjDTJL8L6eyeXk0mhJWjwD4RwpYmjquwk1zbr1HCqbEdcWF8jkyvqhHUBIwtyy9GBs00r6CF3l
TsEnzgQhUxsiNcWTM2pXX4xsN3MJZspn23YN8EAgjomhhD/bKztN4A7vMRoOJkiSjUv9AXdcpxac
xFEiKRO/c95xvhT3s2JUrz7wr6Lt9/MzWe0AAlosj1FhWz6iS4hj0ONfW8vOyuBohQdH4IDW72Be
0VMu07md73ClUHFELnJjF0A0VE2/mMIgGkZGmGVu/eG2aXEQOSaaStdLESxwjK00rMnF8OSa53j4
miPh+nrx1UhLeK9yld52RFn+3aLZ3bZxbnJIekUYNSJoEGro6PnFcMtTxfRQvXoNIeL9GsSi6Rlp
IfhIl9Di0xw8F2Legz46Ff/6L3+8quh5kTwLyT5DrHANjqFt89Tum7kIp9TrpY6E8J9ftJ4LLA/7
585iJOcnzUaMZIs5azl6IA0ZPivdEzYKqsp6WiLKcBOL8Gr0BFjo3a8KrYhM3TrQQf35s631Clzv
WoPR6AZWFNw17/urUZSh4Zm0QXBW3MllEiX0F/Sj1oK6KhdPB1YQEHJL4FUUk4BeqpJu+Laut/Gd
QUy05rQX+hUgyANh2LHFLgScwIX4z40Jgf/WxyTNCGzuslTEBS6q8Pe2sn/y+0fEcroThV5VIHlV
zkb+9cuU7yxhbkcYe8BblN24Sn0S+7lbYLKTlPHOX355SGfVaEhU/v2kmZKsJaLqI4lcgj79FLsu
QRszyRcT5Mps3ENKB/RL505D5elAN2wncx3m/0Lz/DRp9q64S3vZSnU/sNTxUCi4Skryq5SbF6o5
S1qThE8zWkSW6jtzBKhwHqJWfpoMkZ6WDyaZ6D4OsDtQ7iBp/9pvPQDTCLjRwjB3b+40B5bIZOT+
s14+BoO2j+iD6PjZ0b2Oeh+Ynj7BmEakO72F+jABfY1OAQnlwWlMLYlswoOvovcVpK6hssVkq564
MsapBSs611wqNPYXn6mwzkwwLkq0So28xwjpsoZ9JxluVvy2yMYSRPxfwMFkODPTAQB9Hd05u1d8
O73NKWLPAQOk5926zevRUf5mswXvgXOYQrO3QvPYxgZJrG+lNkl7kH8ecPAIIr+kGOF/ACFoyDYC
CjaB3g8z87z9Y/TWK4Uo1p4IlzYOEOtvaMw95HqjCukatXjRY1RkEMRd7y0QlP9ilOhKO3N31Q6H
2brjPwUXFnRx5DNnk7PH4+sWHfKgof313C0spV9nbLgPbG8rKnd+ETf2oSWGFRFicMZXCRGjF58b
iebg6g3t7K272dj52uIwVCbxyxhRvR9pd1uVeV+BF3JRd5ijpq9HRCWgzTNSAp1h7XorIoRlpg/E
6WgNX6oxgzfrVSiUMwsLDWUZWw20hk8QSTzQW2S4EBXjV+IUkPtT7KvnDyOM2ZR7cCLpgaEa1cLT
f4aaBYBHRSjbUMkdJy3ugQPJKktD5WtXgth9i8LFitJRN/2scHysZ4jdo41wwEPciUvkQWxJ9HD/
8qtgFx7jSLdb/Onl8M+37cFA3phiIu2lTO+9m0PEkAtcImc1pEAQtEcN3A1W5cgDNEx+/UlA+1gq
qjUB/gIqzDDUMGW9FbaGIP+c5hw38xgn4Dm3HRklifqesxvif6OiG62XAgkws687puDt2Ur/4Rxw
vkLHyceriJNhqenyvYCR8pTOQfS6dZ3fsJDaPDCBQv0pM3Egcx1h2hC4XLEdmEPywoJ2AVF4wxmH
V984QCajzXmKb9ankh4bolJz4u8Zg7YMKSnzQu3reBphZd7z/yomZD7EQTOEISfoBmyrpzcv79aA
MDpo9a/YJsB9BkRVv0FanjLbrq82/JM88o77W6aSGNX9Io11md2rkNr83Ho34I8YgpBiVTuWzHIb
eETwAmJPqU/ETrzSSPKw5RgEvZ9Bvn7hcHmPKtxWuXsGkWe9ZuGW8uB/xjLbZIcSlGJQ3jStF4AF
BsBWQXjmXm5uCBUjHAh51RDGsDTNqHmTYWjQyO93hrtk73jfrAyzJGqoDMxjKSLYoRlHSi6aNnZw
Wz+M9JphXaQha3ooNGx3qGO78Yx9uBIIE49jVHlP8BA5/sNeun7+oPUCi4lGqSUNMw3TP2ZPO5IH
yYEqxX38rp3ed7MziYe9uQwYVoY4ieaGK764nzm337UobkvJPA/yNRQpuo4ey/rS7T7aD7mntCfc
3jKJFvxrDHxk5gSmCK45+o2kjOy2EPlbLB3iBqjCpw3iojN/Hy8is1gbLv3ciVRJnCmEUq/CizLD
+k9Sr0r0RuVpHodokF68H/L12XNXGqWl7AGorMVuHPgqLoFqIkpfALqr8Z1uTUm+kVKsM2WOC/Pd
bqkFSTI5Pr6p50vszY4xLjOld1cKOJNjafGfAQeQDKg7OFx8WCVVvq6WKMF3MKUYGhqwbqHNqgDy
G5Bf0NnLqYLiSIgkmKE3FB7kuciY+PYhNqpFzSZgYyiShbOnzxfe+Ab0vg0t3WrrzEatVlLW5Lhs
0YwVsN4oUpdmLswaHrwLeKBz0CxtC4owPZPw2pVz8mshs/5nqDBnfb29Zk2p9MsEI6MenFCEOuQ3
/9HDXHaVI68bESmfWJPbiybJ5lvQE6IQFAmFuoCLPNzKiGNIc8oidfM4/qmUz1Fqy0QbpfBom0ul
M+9oHVFipAHCsguwhenwB5veGOFxDNcTLn9sqFw4Kox1nOc6NIDQ5ePEZRCFhXCe3th323pgsHCS
DOiKCIvpgnEPZUBKhOzcjPZTVivXsS++6UcJf+bW5ox77Dwt+1YNmA77odMmSCUn9uBwcb1Vhb7G
UsVAffTwEHhUGd9y+nKrdklZtSrTB+KQsVDMxvQwcEoOEDjIpuoH7EOPkmP/76V3usAHVrof8UdX
vd+gGXlB+ObRztIpX1NlldfRz10fppoCla3SbWyPrrCphkNdI33LZl+9XksugrXwZgoiNfytmcT3
XCYQjop/Sy5Wk0B4EBf+moR5z6bpZm8Kj8+3Z1zuRs/Ci1zy9/Z/NxZGEoClS52K0cRG+EkhCgnX
DDimBbVgMKsV8zycuU4DJ06D0pINBRwrUByhBiOKSuTJXZoXA9sVhOiV2gOORRDSTtjJ+MYevN6S
KxOo9B1fR8heGO50Cei84zKMchvV4Gzk9YKz6PiVkT34bKUNgkIcIkziavbnGFa2WGeSOqvIWN3Y
SO+xadanRKGIDsVf41z8E7YmsDl35M8s77xTA7oO6M/jnEMuSZXmH8cltfuXmYBWR++b7X9ZpqbY
vq5e9gCWq1Tis22jafVFzsYPqS5yYEePOHQfruRy6v8yHrN9BMog7Rvwie8Nnq+lIdx/qeOn90kE
VTFn19uaRgr9C4UJyHKsSE7a12bMTx1fbrwMdJY2ebC6umgBHMAit87QJzx42pjys9+e9CEzZRSk
KPy/FPxmkxrScSDsXMWVi/NPcTwCHpEXDlfs+8vZZ9udDN9xeVGPUWFh9Oq/o9QoaoA/kIz0zkIp
7fobP59TX+PIiDgo2g7yHiK/B/gPWf1bjY8zLYQpPKQdSji8tUSdlIgyI/4kYXWqivAIlGBsThaR
ECFd75q9iuvY4i6ckGm20lEeW+X5US+U3egcIZJ4T2SjDLm7EBujtWR5h+SvwQ8rir6E16xNfVZr
7KBQJpdkhYjRrfT6wF/55c9e5H7yQyvklMo/308G/ne/VP7ckZJUhwHqIDO9/W7Gi+movRsW0G9e
2gWuGL65J7g4xBT7IAdgpC/jJAOgi5O6nnmhMMnUeqwuIYyHZDCBRXZs1slxEHU5uPi7TLi/htbt
NOxPXdouz6EuVCQf9oko5Gxwdk2abhrv+60498G0zpMY+EvRx3ftbEmoo+ISdRMUtWUtK8lQ4Cgt
FoppirEawMt9QP8nY2cMzCbvmOAVdhJzC2bgGzxCSRxutIg4qxR+Pa0JVpHXGcl/KTZTjXGooxCw
qeDynu8x9IGxTqLYkJ03tQPKmb+EDngP25/IitpGtE9tDfZWoaFdVx6FFd5chA62LlbIzu3u6SSJ
Kxmq57aMu56zIMozz02TibTImw9eSjLFSJ6GAScH96rqQF9wQ3D7DkaLThNXIuIcDVnUsxAGVV08
1Vxpi976yMp/ygtoNoEAnJSfCIeFKyh56nVEIxSVG7YlJy3MDfKe1bN5KdBD77sQiYmM6KaD/yYP
KFvlnBVHnr/qefSzfTAh9SFRcaGZxsvz+TE0lQ/+o1rVJumMSzFWwBufJ/Or3Zlfj2+CyTl3sr+r
mAzO5DHxKDX6e7cDS5s5puhUE3/2qF5wkvoCmcc2Xifb02VyPigb9ktlR51ZdmtyrT2OiuSQz+dk
usfsYsNpWtIxZusW+3vrrydn/WBJkLwqdJ5tSzT7jVBHBg7FW5Pa1F8/K/h7pLUXzjGakULpw/qU
y1ouklZyvQbS4N/BJYhwryxTjgwkoON43Ka8BCBolhOoZByrGJSithCwop+Bm0IC5SN0i5wbimQH
LKfoD1Q5oUzD2k9JkCn/LZ1ARHIPGKg0FoMXhJj1+CKI+A1/o4dbsnMdyh2DjMw5UTsJsrByB7Yo
wpfGferjEzag2C4PNRV+XnykC0LoCsamR5dTWYX+wzgdviLzwGewQmVKlyRzKjA//VNDXra2JitE
KYWWRft21ccQY9apj5J1K9ly8ICV9xP2tfSPFswojhCWw3uGsxXT0silLbOZEfdFicgJ2lxgcJcw
gsqd8EttGIAc98EwOc5n8wT7+4QCVb9w/TLXFVeZz3LAuvWSH4cTHhdL3/7PJMVgqMWTHaB61dES
8ikx73V+KBlhzHbNT4lvxJv00rpZH98PJcn1BDwwzXnn7zkFjBKxzTdNJ4kv9S6fBuOw9v/gd30p
v3GWyg+GIlVp6AwC6QrmDNXuoNXTxVKSgoz4GxiYfdztPkunWZQspFQIDt0UHyfA4G4u4xNndC+T
tzekCdkzf+AMPjEiO2em3/kCscquuC4JAL/0okj5PDss1fDMDjQBcXf7sk7SxtINobAOQcOJzs/E
yxKeBF9mRlE5CZpBbr0wtqua6ySogtJl8heGy4oaC1VH+fbjp5qz+yqnjLwTbqsrWUFS6nOoa3Iv
OUDdrwxSULm1U0kf1lOCGWHN0qNoj6aWWNdNn7ujpk4uRu68sd8m9Gxi2IWXGJxnIx2aX2AXw51M
R5jim5eFL+zp9W6WELv8QeXWWnE0QnTYS2oNAA/wwMeO/B1FxMVkaJUbT7tBDDsxjubajEXazUMa
fa4ruO2Bc01K1Ar4QhofsbC38EOlyDeLCKMruKAhj1ML+54LDyWWmCCsqRmIHVpYYmdIiz3r65r3
Bb2XuyBGBIMMokQ9fQ49SPyMKdZwZ9YZr1qSC+0BmSA6UjC05uGQAbBd/cLLr4Om+B3A3K8KRkKh
1rvzPjovbmh7INcFa1rV/Ix6Fw3jkNHGW7s7VAFK0YrhbyELXu8APGF+F6nAVPCRqXmK0+hqjSvQ
Mnfxc2W3Ho7G/ES2KGE4YGakg5jJMRCD3bvMtT7ML2SqVEI4bxLH/BnI+KJJyZksySgA2RQ816UB
WxCsNujg3+DbkQTUdVhKpVRhz0+2MFAMQv9mmVVcV4Frc5iLD32d7Ogxnlqj6CSWEtncl9NHAyvY
L4+0yyeYLkrucSY+pjinsRYBnLbx8/Nzlrmg1aJXvPcSOOseCqs4s7fhqmSy9AUqSdbsJZJSQT4N
TmQo4FxlO/hiXdvJ6R5WtvZxa+pXWop1cVpq1dIOjEO6uEnBaHdRMQA1tEa8q5wpAhKy7j7DC8ut
eSBEkh2eg2dJa4ODJIDEYLZgUTztT26QiXDTvsYYmeEorqw+o8JkiDHwMldthBxtZDMuSjCbEQKM
dvJT0zumiK5SsnBCvygHUYZ6+j/VGreAW/vAbubwlN6G0c3yr2gp2kt3KFxf/hzOj3MO3/l9ODOb
fJ3/Fb36cliB9D+54LLnJpNSH+fwPjXphYxWZpL4iHd9NTsX+lwa2zZ7IfrRYuWA1tCjueQ6DF0h
Bf8+xSWt45aUyVEeMCyAZ4XYx9Y7fetpPMqrUhGHJ/0aRAt+htw58Tl+HB0OGXpL5t3kP8wdlOlZ
rzlUM+q2JfCSk4ZXNcyzRT1GoTsm4M6fpQ/CBMAbKKsI2EgOuNJgCr+L8/SQLnqK7GLVGRBv+WYP
MN0w1M3Qa0EhmiLIRlidB5Zq/8FE8kzsf30F1nL0kHB1wfeuLiH15Go5x78F+Bd7tc4nKaMa4aU7
us13VNLpRfzaOoqxQc4cIlK4rgIQO0VrVJVEBWDM/RxrU1AR+wjqMmu144SXYJHy/1fqwqixBCk/
1yw7rq4sVa8WK4e5p0ewd+1JHT0ZnAzi0LwYZbfa/9uwTeUOHDGUnfKaRYpHWFCqBajaUzym4oeK
CugBCPQV/HjMCTXVEl59RH1QhNTradtG5+zfJQLb9sy6N/v3Nk6leIMxeMwdjmEuvmb0vAlbQqUB
92xoMkk7jAISFzdTt3dTeLFPdcSY++AIy09f8uU4W0dl+7WLiupMnq8kIg2V3njMm2dSQHhsnmZj
EzRgCeH4O5zIu+zfTaAHNYAwFrcYqD5sPLDxU3ANllFpmclsz5svGUWX/Me8sf30E/6f9CRHOlzL
oEt3S6vEv7zQbEm2Bv8oDjB56WFekNTYptBuUzZN3M7iCmz/HoQ1F54rfA0xkaeiCzXLI1LyxNfB
SR0UQILJoVvOpqHiLn8fPPwlyhTBsQSm8yFI4w+od2vgc0XPADDOp3sAAT5dQ7C2gYHEQlXkeagO
B6m5MQolS/OK7CUfFI9XEl5jeW0GOT+B+YKwsfQRPIfrG595lxAbm7x1y1+AZW9r4u80jXMagQHQ
L9z33rmSSYbJ8sOvgbNhG3q7EZQ2nAwtbalS5VXOLHho20wDlhld/1t/VBZ2X7cfhz/CkhxpnChD
5Is42gldfbsEEuZcmt9Dct0UCFe6oYuaOFOzIpQseilKPv/cZWv5PZfisu34SZtIbQgx8/kLOI2r
fwSIUSSe3JTnQ9Q9H+viWlKpxmg2pBBw81Ik+Z+5ztsGHiAU7m+ATnreRAhJabXwXK0QAytfs5eo
s+/ae66VALIFRegVTMciXQGoBGQBWV2Lfmi716J6sP95PD8sSYqAJ9wDA9z0OkVcZxfCz5oUbrPA
TpgSOFVowKuOEZop+96JKNBkssLCo3fzlFt3ZQKs9Z22PPMSfkf6FIfPr+O5M+Owr4CvZKq3lYtc
wFpA/tjqsR4wunDM0Q2bLJAMaiH2hjT0ExKNbMLYqUQVYsDCPFHoLQZShPpmw/Ye5pSR7ISNnqhZ
WFHUc9VHZLNbd7wzNQ/ADW+B0eOcC6Vv6BG99yu68nlpMXERPatQVls6KzkTmFGVUd/SnM6w++Lh
1y3isgtQxtw9e9AIDuPR/aAeawrQTorWm5HkEj96wKSHpQzJOkfur3uBnwTWw29bOQ/EWpUkjl9C
+lRghbbbAMPTwKXQ+FZu68A+T1KImM63J/1vb4+X81dacgb4swL+Bdjckg5glCWiXTtz6em505iN
+pmGbfhPsTR4y3wABB4pEnoPw21rDTPBrYxkaQdMBYPsicoWRKDoxqPmMELlznWXh/FgmmHF2WLW
yjZWUdsXfLQWLJFOC+oe6EODTlFlcv0ijh6e87ohQNLudmtoe3m4TxM25Kfr3TgOEVlT3KarypBc
LOJcvMQtCAqfLJtEOFT5N23j41NjwuqKiXHXI541MGtWUM9fyzsj/0e+ZWbV3ylD5XdsJGRyeVRK
mcj2R5eX7InRDKVej6dUIKg6JZswUqLo4c44B+mjudO/3w4IX87JI9fVxyRcLmnhQgUOgCUbl4HA
HRTaMKKjKjg4WwpbpJtyMLYNSLNddz4lwQhY4xXZsUzGhzIe5nyuJrATgx6nD14NZR50MPTUBCU3
1cZzVMmeMmweiWsrDcDWDzGeETD7KdJs4qMqLlo51UTZEot3LYXHWihEmF3cU8jSUUbFoWeid5eF
ghOaaE/DEyoHCG+a8VJH68CtqiTJa0CvECKTZEFp3pxYCpmqjlkHFRWVGH3dpJhwz8MBwKBBrYxl
gi0IEnSZpDgBmqM5cIVRFUGJapJtDtzjdW32ckCMrkGSCmAr29nemnuPqIFY2U7Z8UcN16CjDG+O
7zUkrhMYyE5JQ5eVkobybmlN58WqzbjzzUWZ7DyICkASf5XwCrWyl1o2+FzxeDeoCi+ZjFC+uEYM
PYsyXWvp0vyhj3LS8FkI1fS2o6/3Pbi9UsS5AtWUD6CfXxHM8FREh2a6mIiXf7u94FJMiwLdUbyL
CM87zDccYLX0Wvy2J7SZHX7DSP1NUWOkc+TIeAEQtep0QStquhzYU7/blJwRsm6gyZQlN65ymMhb
0GMo6I/D+8hYewH7QsjK+zEStKAlNlQO/u7BSRYSYJ53X6vtTKs0dERwj+3svdZ8AgsFLoAy8X1W
iVZf/pg6C4eysWJ77fGBGOkRW5A7xRZlvYU74ddsERUbyrLtVTlGVT//Fyz5IWQ5re564d4K3K5a
8holKlTv7IgOgeRCSyKCuIehJmYaczvHfmhFlB6JJId10RyNlNlCyUMli5C+2ZfPHg9TjodsgAFB
8yYwXy8KD/nPzVS6s+5Nf4qYaZKO36466xpXvOvFtkd7Il7lbFxgCRW8fBwwkjobOZmmlTeLRGk0
dys0s5Sa6pXdS1bIjFw1sn8pW2PZDUoR8fE4kBNcpjD9qAx+2d5bDWB5Fo3KqsyV1DNAiUB8NMn/
fi/FRMzQx6e/3Q2CrH+zktV5Rgv6Bcn+vyC20KHiM+YQDN7WSsBscmtokdUXGmVVGw5rbNvj1w7C
OvugfngPKO/nWIDch8MN7mWL3fm2kZalUPbeRNSwfZjWWRVKr7HL9SZ6aNiwpHs4KgZuhvzAtZqB
1/9NFtRs11rPttd0QsOl34wWWkW8eVw5FTSX8LQELqoXsyQroE8tr0B/IJURqnaW8Dd7/w/3sbQE
3xjdcpNQQq8u3+sMRZnyXAl02AEOCIImVJ1kK8AbW2/aklzmacX1qYyDkQq4OzzqR3VB0a+/Z7R2
elMtYLzSMOf5G5HOhudpS/PgizZCHy+fGhIydNznlBJbuDtMl10JslxX2enebtHYQgTVP1WE+8wd
OAYsFvTD6jAJ8P0ea+27Av3PSbNG47+XiLRTA+KVbbE16x7JdxCmzQSwr0n+eLy3ulgHu7gK5KEk
fBROPGgZXroXHZYZ4RNXqWEMgk6OVDtchu+EXIGz9M18L+/bOAOzDqH6ldn68lZ5ar0Kxlc8QbsS
xzzMZshHGj+mZ7o7eHZ4v9Bjo/ugOrbHtw6YjwhrBsoDQ9EuOKyfJzG0U83HnNdQ9ESzlAM0Ae9a
ZLQi4bLgBeX12cm4H/ZJQ0yLNhQs3fvifWq+8vUopMAGze40iqKz3Cd2Yea7U+eZG87LItU69ggi
qGk8Q8FoI0xjUODK+2wLMf0NvS23ib3fWCINmEU2JuhCztrEiiUgOqQcP802yejg87p3BLna/qev
f8M+N65oYgnT4tW9edZ433Ek2qQw8sLEIPaLCRiHRCmTtjs9k4YHoqKbg1i0ILCCXuIQVpJnU9lm
Wfdo4kV73VFPVGHluaUQWAKg8dPfq5uEmOh0hyjhzq5FYBTNZr/IZFaDKhP2A5fzT7LkI7JpXbY3
yivueJKNpNfl4JQ/NyK6+3qyhUlLpxQOSFi7T0bgQjP1gTE5DFIGAp5Fy6tqTi497wSj3VeupYGh
K0wxWeSuBpEQTrSaW+0ZLLcbvNqyBWpsO7ftyKLI7kXoF968k/62Ez34pkfm26JsfEg22dDVhZhP
1n/rKLtJsu+7WoKJwa/xNfGA2AP1wLe28bhOqggGMdLl17EHAXifNJSNvKQORQEIdnLv4hjAMQhs
z2oI85wh6gUShh23VbO0hiNUPVwg7H4/FAEc+96ObL9Hiym58dT44colCOejdIkTGLf0L5bR4cZP
gzRXRYP44lAEZYbTEwwiD+ajZ9tU4jsKpXDsZBojD+bBK63UciwwyI7baCbDKjb8YIFAmuxRQIus
SvwYXk8qXviKDVOoYXm8qe2DrYEAeQd3cFajItXp6jj6LVTsM/VVEvZI2eHjh7TTCU6L3ZTfYEkY
LBYD/LpxI8h4doXtOoOOQJN8V0tlPN00BgFtEdZ2BBFVIqVlhv74pcmKZupVsW+XHDJGItvckDjY
/dScK9CI2AZx7A8Hif6phe4Ke3+1s8twLVaUvMTRaSbMEcUwetbZjyNOqkUL80XVbb6fObvHTui4
QPiUYMtrBVzhsSrtpnYro6ckI8clwXqyD3KLsNMKPLLsMqLpMnXKHaNJOiUdjm1/QZmDqetZQafD
4GVvreQNa4p5ztad8oarhVNbUloaukPuhrLqlExG3rw5VccCJRN3gPVcwiL7jAxwuEeZyDOJTnCv
SjvRUQF12+3NOubefoPj/+lJP1zFnDJCFVJutQtHt7ZWxA5/8BauZ9csCoqFI2yDWzt+7olWgbN4
oOdtF5b7B8hxiIVMmyANNXzGwcmK/hlYRMztRPWb37zQWcUWF0I52dGybn7j62ElToGtOwXMMHeT
j9/n/craUzVJPwr1VUpDOavMPWFV5ZDVv0jSb3TocNQak3Cn1aho/TytHhyUgeXgCgsFlrpFqVHQ
OAfqXFeG5BrpwhKFA+1/a22U+dLFPyqtSY1sp/eBn+nKyRiVYB7Xu4ODDwaUti+PYqZ/ja2/YRSD
bZDhvlbCVEsB6geQ5YR/xkdV33YlaBc4Rw2e6C6KDQCyVU04KV1cpVSMG6na3/F6SWTAR/KygMW6
XBm/BW59pto0fXwOhoV3LV3qUvd3ltXx+UiWlllGLuitGfKfE5Tu5htMed3TYfPh3iEUZJ+ISx2M
14wQYbHxfbYyLf+vw0n/2HysYsh1V1p7gbc6Jx09DPhWIWS63Ctt37THG81hXmZL4Tl2LyKulHZ9
Ef+Zg8boZk4NHvFNXVDiRvaJVT/Dsffn6ifN8IbD7R4CjnWRTJEyq8LC99ElKmMJoh8J4MxiQcaq
AiONE3gRhMWV5KIB/fWtJrA/J4Xc4a/BjJ3MLRylZtE688jyLPm9DWaM+CssvpnuOj33ChPuhtJ4
fWvYuIRat4eaFBB15cxrjSeiFQCvMQ2ME3ucNJouBaUxrgUtVSXDQ24W3zS3g+URdObbiNsA5MQ2
CWgOvhEK11vlpj1BR/Q4VWztzD9vopm/mgE+Ttl5xnOhg6i3wQxDXKZzyHH094sPqauuGhiDlXv6
wjXg38/snC+T1i4kq7C6BLQ+x1WbShIFPSW0Lb8uny057N5SZyvjjJccpL+cxLd8Z/Lqs2BkprYd
kyhIvqqLh0SMzXp5VlGRiGn5JqMwlTqsWTBcJnXuRROoDUl4u/BCQL1FjSH/o0ec8NzoBWBFLA2Y
e8BMhmuC6QnfnNZcgIAe2xKYMxpvJJXqXQIcMURLCqwFl6G3zdCxdfWjPrXCMhasdzEMFq0oIACH
u+iNsXn0BFwqIUNOiffLHnQ9r13+EWVdE3KxY9guB3S6J0eNUe/4dBJJ0QLkwkSJjE528tyBCLQn
yKlVoi5Y6Dx6zt02imXfcLOISIZfyNEDMtLRgzSZVKoXrzGliO6UINfkj5wQYXlebSlgwueiz25n
6tMvS1oQ2TmDQAcXiI1U10q5GWrXOgY/7cQiv+MDDnlgko7sP/joaYM2P1YlfvVvlXEAXQDdF6EP
Iqr2xH9jsVeKAt9qB7AaLMgTwQ/t4NCEAtMGW6kxzKqKS8HNGe8J2JCV8pMQy/ZuYJvg5SlmeNut
mL3irIRPdaoOSeW/lBg4fyTDLlml6KiYlKa+V3q31+dBr6hCFbf3hxBhnrcoLMwYtSmclYvA/MS2
l1ISO0YDjw60/SucdoZJ/IiLV8sW4X31N3SyMYsXvlcMH8CcRAJ5bG6W6IyjMeCN/H7uxUiyfa7S
5UqalV1IalvVibxaqlR5z0HzHwvaJONNOHyL39ERknJ6VU4HfqnlYED3Fh2ufLWMffcZSV1/jo06
FRm+rCi6ujatUXmpdl2tGX3dFXaWhLUWGuvZWZetmjO5w3Fn8JepudVFlnrQG4p6BhD0mV32IxNO
HYeeDpcg3ImJSBXODUE7n84ZniAEqu/Su481Jg3iNzeSuPaSMp77PIarRqCyiB9+/FIMJbWWxWHr
+0Sq+OjyNbSqcsTNpzxZkyFylH563vYXffu46LvllE0WaCObUmJkxEtMfYb4p2E1WrMTZwtoKaGb
GLVWH0GIrZ816yiEp9oKQeEskFDWzBSWuFhLcCPFOLmh2lbpioU46OtKO2tc/or3g7Ag2b+1hpHK
Ebba0bpGrVt5Vou8+EJziw3ADp2xUBN/Ex4GvJeyW1aYt77owySwj3JGgZ5tidqkdfo2OKuAwnyI
HCaW5DlbfbWDtp+MkrijtWFSNNfdk1sTmncFlRdyFMjeo+9iQ4kGH9gYsNPpBJVU/0CrGasHKYxh
UHuFOccVr3b7qLN5+UPLpjZbGfiS13KlQMYR6obybC6IU/zhbAoqslRxiyHqAiOJVmOn0vtmspTB
j49bmIN/A1pJPHnv+IZCG+IQpql1Ls+Uxh9mABmwyxHreM34E1YYO2t7ddK8PfyFidA5KsNl6nAk
yr9Mhw68BjpxIW2SeU+4W2NeuGQc92qityjaUEcCeh6mBVs+FNRjdig4wN2PuSVaY9IDiOcPYjtv
Q6RsRSVP8rMhaiQ67UgmUjxekM0U2oIhiV+AUU6NJinPBE94Tk2LEh/RGuZBhfccYTy+tVR4gKZH
YrMzQMZXbQxSifY5TBkUPThLS4eAKaWGiIw8o4/nybGC8Ij4/0xgaYSyXEumrfBa78gXoqXi5+ib
Ep7cPZSSoGhmNLQ4N8ChNj/4zrdxgVKDpkQFzNVI51Ntcj8iYo+2xVjCpiQjJx+MJDdUoSj3Cas0
DEgIyT2mSRlL0xjWVA4GR+tcOj5Xyj+KliGxxibEoJ303LwfuOUqJAqfq3DiLVqHgpleOltGKLCb
56LZHBBJWl9DzBW7dnRtRH9NzNg9jW4ZnUTxyu6rDc8YCzABeQtFJcp2Ae7tZWelWOAor2kd0Gqw
zWYc/RzvqcohPIQwGCknPziYaBhJ/PHrOoFy0roR237VP8D71GtibM6ToQ2LW7+pxXkQDrFB1lPD
JQwUZW1jFURfx9LxQkLdCvz09A0ktjjpyeBWrS9iBLko4TH5q20pP5w/cDhmtr6GWi5Yk+wQLc+7
0Ls99jO6Go7x15s20CB16SglTHDtc/dNkCvad4ClkLkpG4V6sdpse6CBHMP9p0S4H48xDNVmO9sb
CrndX0gAszYoCBZTeJ1ii+ExbFO//FYAMQAvblIxRcCEw073AXCLCh1Qc2BpO6/JK1QvDPykBhre
07Wb1tCcobcx0S47542xty+MRgWYoQjZ3owzTtABQhe2LIinvATcEP1bB06GdRNa5nMJPdaefO3h
uurRob+3yldYoVGg2bpnwNUJgQnXj3KI8/SwdRxI70oU44al6MCObTuFF7c32PWZXrfSYY1JbSQL
RkPVFhFFItVzdP8osTTTubBToM26gJnMVA3MdbiNGTfJrJ3EnZ0rmUeznb+coGA/c/WKuHsZPddw
+5ItwppBUv5XXbw69UMU/64gLA7MIIsHX88RWq0vwvrh7wW+J3yhqi5BJTLdPVDPmlth0wF72o6i
1wr+BH8uJHWgf+f/NzJ5uWW8c+j0KEGBupAJlUZ6Y95ZiUPjRqO+t6X/7e/K1ffsl45Uhqeu8F1s
3Qs+dBdONDlmRYetY2TkizSeOSkEgoNLkAwmFO3HgMEJ1EEBtOOAZN+qW2XaozEha+QTgu+BVccf
Bs2Mg9uBNTYFnlkFvz4ZM1IEe9gPlEL8BHPv4jYZxIoQif12VgZSQ16ZcJ0IQCsiPdNzGHw34oF4
E9UnovU97ENnAMrn2ZDOk8Ibj5ytCXpZTEE1DuudK0eyl7hyer13FE6lJQUnyDL02NdY6sT3gvld
WfwwOXMOg68s4xpn13PWqp4DHiSW+UhIYANiWTZs98N8NsXIShnwzqeEvyo88of4KQb17mLZDPSx
UXcWFCUq+isKjX3oNXOkHE3IFV49utZmvAcPLIxOUAXuQ73NU2rikENxYzpM8VpmThMl0ZPqh43m
z4KhdDe0NfkYV1+T0fCFyaxsZmet/5oGNBxnV22DA576eX03X9NSqDH5NgKXBb8ImEISTGebt0rh
E/g4k3zussYKPKBrXYPHSaEsoyUomAgDMNXC4bLktCsFt2fI90GFoeLRyhclT5l40h4EP+gNTEiM
gCW/5/tgk82SFYt7QvS84SLaQdrzIhRV//EV74cOPHbOFfMWuj8vrHX+BCxULfoMqr/vEFegGRXo
7gDTdwNEAZJMsuV0ohtCPPjIOZpoiVW8eUCF+5ptko0u1NOQaij9b8ZKuUvxtx/hlissfw66SJVA
Dx+yyXX5oUYcGeKRS9Q3Is6llEmu9ofJ809LfppZshlEEdmqTuIZaghVGCvJFdS1+1Fyl0v2iBMz
CeLlwwdloCueYDNi2vCQ6SdP+00ulv6YYGdScuaa0ysdgebjhf2LNul3lvrpEDU1QCi4042hCjiC
Bm5yo6BcJf5cN4K1vUgigt7baBvdR5VGzHRuBCQB5MUN2oacuiof86OE4T/PlXDb14PM8uX5UBRY
zpn7r2dt4A0HtfWIGK3XeRpST39ODwLz2HtzgTUvxIgKNtxHwzgqU58/FEUXaMbviwv5Zqplcr5h
FBmx1JoOaTvsggeLcDviiiZKm/7UXf9Nf9KWuBpAejsvwXVYIzbGkXcaHBAuveNnlmc/pIpIdr4t
B87qLOzQatIQyzqNtUIJNHZKID9c78+7DHnsgJOGaKGPgpKqSniY8bxpDz3Fi1ST/BFJDyd+FDPs
RD6VWTKx1bqVH+jtIXZ4o5YVxPiGBf5paWMbiVSU5ZP71eT73FU48NE2KfkakonlDll/2WmNJ4Oq
vIjdJXLrPdpgwnIzw3Wgi8b8icv2hIc9Lgbdd4wsrAgFpekm4nKZX2UcpxsU1ZRxMkOWLWMpQa9r
tbC3KC2lVKjiO75PjSukjc/Tbh/l0Q0yLCyJC56rCaJLSZzmvyuwh5XW3/9uyLMcIZj5wIwMXzFf
xDdMoGYznIa6+iyet+dqeuXk8iupHsOlwLhwCAO6vP/MfI5o9B6KfmXjEabE8jsJnvhCCZeEUFT3
bdLha9VJB+PwWjjXoW2cR+TNvf7JpGbK/aXNuQcdZqZCPTWZELyIf1CrlR+VnMuu/U1i50763FYB
BWwIsIZTODIToXGCPqxb+4n0grnd/JI0RRjzBVb/Doa2aITVkhv9O8kT49AwdYDQw4+I4N2jaLoZ
K6r8pc7XeuQ0wzXJ279jwG6Qqi9G436ommrJGeYTGcL1oM7MC35EyPucyOXAbKJgYRKf5xq9d2jf
jsM46F4x2TjDbtvmKki4OKTpNGErqPT2SzcY3f2NVp5goeDCm5eznGpi10lJ11n56xnnouPGu07P
3N88WTeNLMkryL1X97m6yx/DR1lEgR9LYC2wwNhZ/0LuCfMKnYT3PSehwgboETKQ4y/0y+am8GwQ
BjrzXV4VY8qlYVEiLmlj1AfQ610Y/mS48l6PU5x29viU/IUtKFfElHD7fyt4swHoaC76kNPl0c96
rNmqKJXHjy64IrWCUQ+BHREuUlFK+guT7wsOHj52QB9JLgt345SKMHlogRjrGKG/9RbYQd7ss4Du
4f0AtGNocBkdnE2BaG+g6pDunfPskkRN7l1WEDW67Im/+21/iYTFGj7yItzkU7k6jwrsRHh+0Z2Y
YEQTL96DuFOIk+hrMASNLxsEUIlpACbe6wHM/RctVNZfE3bRNnSCEZK+I27/Pr1cIQ9cw6hoBjZm
EHU95fa0kjkg4xS2K7lNUS1zSi1GISm8XFyE+ZGeYtGd4lZZRQzJxiUPi63VN7RAo7kOaXgfig/o
Tk1VF4b9dUCdbvK12wrkeuu20hDn+YXCWB5bgkEfeqyZRU9dhZGoX4Op+jxjrDaljITHd2DKrms7
ly3xHZo+d72ERiuKmQYpON15oPmjDx9xmrk8AGca6WcufRzvyKqgxnMsgQ75cnvjf/MNeOL2ikv0
bCeLxEBxA5g27PbDy9rVOUR7dfdxPfqqWM6ueFRx5TiyQRbb6ddppoGarVLmh1/7bLO1idFKjN8x
c/nMVrdKahZHYUWG3Du/7dgferwUhhH7DfGIbcx05vFTJSCA/SrG+waR7EEdsPRmiRGvvHJOkokN
0KsgJCV0LjxyGaUYf/cQ8wIg5X9I8TNr4bVhHeDjXoShuAo8iTnyI3oFVODVqdW2jfUEVdakJpcX
5nImF43t4b+7NvF/nqqnmScFbz2sIMyID/ARux0HDoWJgCAJaJ8bzYkeyUvs5dnf9pm/GKYTrmXk
ZVNfbMgY5yyIoQmlkA7jfXUVxJUz2vVf8tVlpK0x/kjLWdZzoL25mKk+iXUVQjknt7LrlpRhzpRo
zscbHPC6xcrNekFRiR0+zovyExE0L/euKbkFGknMDrnHsKfzJ2+A1qBxco/H9CIwGK32E4powVcu
/pguZg2ZVewekV59d52Re4wOzJTVwErOoKPXFHtNx6X8VoDjWV/sRItFB/JrSqHmbqX9ry+oYAZZ
Xj/mzow6Bf5ls4kXZCjSS+Cd6B7lKLWMJoTL1L0uoo/qpEQiLM01dPEZ0QU2EG2ydbrCjz3K1SEE
EKkoZklUFNEVfKbt0eVuMJEIxyC0LqTHPGIjTCwwSCkzM+zg9xXR+k0MJcRw18er5T07e2eu0Qcm
N4WmqdeLHvTmARNWWvn8LM32hYIkHaMdkeXDdLq8JE/I8Kl4xrGMFqQ3RHfhRwvWswabfZoufuOa
GLZsK+lX2o1Uv0dsF6aSiRpAQTV/ezk8lhdxoLT6xOU1klyPeFgquVuuY1MXDAo8vU6ot3nGBf6J
RTZitIHM38uVNdE/Bs5tCidC4f3yArayf11GHiUAboupVA2+0GEInYf7rMVfh7wqfOY47v3i+6m9
IPaqYvgqH1OUla+oN400NOCk+xpGtdMXiv6MFDdDJAN7GKBxIHHLA13bpHy+C1aNbnQDurOmMNw3
OGpX5ege0ArhO10Q9jGlwUc+hmzSmlloKkdFrtuSEuRmUygROP4sl/Mrdm4LxaqcXLHdVrzMGhLN
doEGXHySUiUkUbuqZa8PnyAy4L+jum60+J+bFYqFl4jc34qFunXuGeo8afvlI0Pk9wROPmN7anTa
F6tLwEhe+k0bUccMjXX8iO5Apfti9SZNYab3ZM60mP9HZ4bW6o3Tbj/xzgxoAkCz/iryDt0KRkwz
4xP8tM8HNadDSRO1rD8FwF7ybaeprH3XYsYMXB7ucfpkQ9pllZWkxs0YY5Ly5VYrspj2zISm/i+1
LU9dbPZM4rN/8zGY3wQ/V5LBlKT+SldeQMkuSlx41uTqn7bIYJ/FT5XWUSm/YK+eFqzU6XD4AKli
KV42SWg8T+Yngcm6Y7itYGauin5E2d4tjLuc088e23ZOMB4gSza8mORs9I98NTnfJIP26RU3LOF5
+ybo2NHcITHbkogoChnDxRImTlew5jbzJeeNKy1xlzDU/NUI6f6fz+0yq+SjcSckwCTjfwpcCCLv
TM1fx6blOyXRJsRjqry6WLpJU225ear3gD2LWN+AHuUbW1cp+CTqJ9oC7lmsyBq/uxnPH9MptenR
v8J4WsL2avmPKjwgHfE1pyr0TJotKoOECMCquehNH/HRcBXsjuZONOISVz/Tm4bHmklBg7rOamxo
T7lFLIb3EWTIx/jKu4Rw6+dYxtWMNuQG9gB1Mc4zmxKuOEKdRiTBe0yJSv03z6cpawvnC+1KxYK4
mqnGPKOnOXjd5glvz1hUJF5p2vuuZ7ZOtpH+HxEWdI7oQoaddfP/zu9qFdlQ98jc0bYUwzvaLyAW
3NcLza2VTr8VMddW7tEYSIU2Zl5W/5msBOtngymv8MTYv9Yzao02RkprhSTQvKzgXbFpD06JAllf
Luw1FUmTl3xm34bwt9ZFiCz8Cv+P/goxtz9CIvBuSRhBpHHNjCDkgFRz7e572beWmiZttJWsHQFv
bD/mnbVUiBOa7/bETxne47fgB2ai/iaWxDwUYRH0ZB/ixFblya8M9u1KNVKfB0h3/aol2B2n76yk
BT91dRstqm/4wXAF07ONtkQZ3BescOR+hfPgxcUXEdURJTIugtraNd3hIDlELr1KIaoBUeg2KMuE
nGTkeW5BdHALEm+7fxeX+TrjR7hbKnudIzj9BUMjXnhccNrMcqD01183qPgg2Gmi3l1kV3JH3nED
C8XNCGozkF+RDgcxSo9eZz3FFmXSCk+bugSiGDntoDXVdfmJJ9YK+dAAAoimbNnTMGFUQOIKzoR3
J4vdtJfBksek4z6QU9KbEmFVf9iirGba2/mz6oGRmZcSzAWvTrzYMVak2ixziMkKs1vNg5XGqbvd
MNdLQgB40zSfoyWa8JQOo9UV5vm+2zdY7VjBstdhBI0npxFF3N7Dn41V2lTaRGga6tAlTdpyUT/G
hYuStSuT6QFEkktvgzO62NuYhAtYLB9kq6VGx7MG+y0zY+1cWZmmoul8war+T+IQTu+J9YogmRUl
/j3z+NmR6qNR137mZWhoNxiYGsp24AKzC/CnZZXaDAntvPZrXlqQBqYbKYmLfjFHf9maBc1E/+h5
giEojuX8cI09hJvm70cpJCtDKEgTIGJwc7+OFRY0+Kn7X5ejIvbynWDsPC2LhS0Odcpr316vM031
uvlpkw1dAFfVYcx+hhMzjlf1nfheg+rgNZjD+/ipdgcomR0BJLRw9wwyQkzzOvIxcacuc6OANTGo
mwBBfYfye4D1acARIqadYRUAMuViyw27kGUnDal+InugsQ1KrnoM6jTutgwrh+iUOehaP6+jZVxx
pTB3QSUAbeBG/iT0aN8xsYYWVAKLy/4Trxcbno1TW7vEh4FZ5qUDmlv2xiunncQ+7aO8VgslTN/d
2+7MC7UptEOyi4A/uJdwdvJFXxMdXrug8uqMDNhRAEAfDtpnIttRSQ5TmvRXER1RVa39TL1/ULJC
e/W7XB0r03/ZBJyGQC0d3ytn610sVqhvzDmD+tnxglMVruT62B4TZMAiOBK+v1ptWNoDSL7ZpxGs
d/cnAZuOWRanPjX64a7FAW0CPSwTvSkgjPdQ911IwHdUFvp0NZXg2PDpR1V+p23K1O0dCaeDs7Ze
eaq97I/CCJ71DvsH5JVhhqOk5Z/Lx12G//berjPIG2PXv+EiNqpB/5ujD7VxqrSAt4ByoCOGL9nq
hpdP3g7NN7Ox6qwlCfJUHkfgfXfF1DdyFlTh6hPR10y/0JRcixPA+OwAATN7U7fVsGJ3X2J04Mbn
V0Mmh5aVItWOpJ3rCxR7CeA5Q7dYVH3BxJnQSG1XEs8XJ/o7LMnnSbfjoWgC1IYtNdd/aIEf51hG
1GsqDGAHuBMkeD/OY3d4gP8yEPTZHwUrRE098gk3Xk7xCvgkt3HPlF+uN7gvguXFir81tfcUv2u0
4Lu5C7FYS0WNk9j1ap/H8ge1WdDrCHUWh9k9QKSJDtQMdxd4m1yz5GZeED9RJrdvyJzy0mcbGqV0
AXeSd7bgXqqs38LlvMZKsRND7bcajYf1/ihBm+/cQI7pdvNPaqYYyHiEcHAuFTAoGkadCW0lMV2v
qjJWwr+kzbx5vsRq04iRQgSqZOKy/9Hspvpd3g/yfLkCthqPwBIhi16MCkF7vyUD0JMPptTVqSbE
h573SnxC3DT2TYUunkOgzk1paVVsLO7L5mB/tJ84PsnsamKoElGPJJiQOeenWy2RHyuszb2CUKiz
Ai5TMrqDSWysNXrLSgVZkGdm1Ok+fWX9d8XLINs14ysTe/i7/PdCVrtnzC+lAHrdy+/QSZJRLOmJ
UH/IM7FuX70QwObIDarmXcJrEvl5JXLJC9rh/Az+4vX1UEL1qGRZVGc5Q9sfPoGJo70bW7kgqTun
4HwmrGF71ljmsOljJTYEEwm4W9K0PIyaFUcogmN/GQFyYNTz6oHcy13R2Ixf6VREppBxU8NGWSUW
sdPIN4JO46ykR9ybZA4GcTWWRAvvTqM9xxYrFbr2dg8EBfHN6IUPsUy+eawgyRdET1BC/P7eThPD
34Tf5+DJs2ZT7cxOtgiJt4Tz8UlOUalceVNCyO6cG36Hd0kf9SI5I86SfKSTFEcomGZ1OxB2EpnC
1gvhzh6rn0gQvjmLm63jEJY76BE5yIvxURDdQaxOvvOIOS9j0gFoZKRzWD3nB2iw7BUvZ99rBAB3
/CCE2Bc2umy7cWCgkzJlKjrh7JhyIH3G4DHWnYh4uI7LMBPiWLtLztDAE1JCaAbCDEB3aybROjh1
7zJUqzqJ28srCirKPYbtLBCP9qfyA0UYs6w0gQoF7a/MInHNDtbbnf/0nkEL+n3nVqXwbQW8rezM
HberIuhlqL9Ame7vWWds1hw0crZlOXJNLRtGDLXg8xv+vD2/a5YxcfeCOlCuTMu8Ia2IiXkk+/jf
5jQ+0TFQf8zF26JhOyHG7wFJm6imtvu5wzaxgQk9jnRfvA+NmXLQ7VEhDXjSVufnRv2zEwuIojw0
NPAe4XB48xHJEJCtvH1Zost942MzuKEZbGXVXX8EGFkMh9WzkGgh0aqUCtPIuMn7Pkjv3u5CnY+W
QAwJRyMPW1czel9KRY8tsA62yqkcpilkSUlAs/Sp5btNZYbvUJt7i2n1Rj0n0WJwvRjEF64Q/0I0
2qMiEsFV9KuF/0wkLk4Owb3i1P4rGwp8Rrlxb2e/0Axf9EJW6PhjgLIhY80Q2wro07Reb9EanIpd
BUN0maWwRaIYZ6NiqsSP8PIG+PXN0FreX8pKQwH2Sg1bFgeg5LgD5+xiSEVZ9ecxqh/LIdNCFm00
bP/ULwiLyMFQ2aZUw62a1uGa2WfihbjpioDvH6kd0h5tjwv0d2dNqOln2/fu4RLIYl+9GqdQZJbQ
E6TMdvlANI2JH+kazcjJLJDntZA9HL31XziAcPq7qLkHYl61jXQJIpq8yUxRARToO0x8I2Dnl7eQ
V/d+4q8tHeOq3gstpo6W0fKquzyctN0Wr4VeYI2eMWjbQGjCOSyaypa+BIS5W1zbjzTwg+D9HuaI
orx4cWOwrHgrHhz4cT1F35D5EhikTVLQfITxoyQAvvxI2R2J6sqmI9OrCG6P0QQArte+zXEMcyYq
02OEwdAdlb9LHXQvWM9S6L1JAkNp2Vn5G5qIX5N9uWOSsfOyH/TOfoCB5/exJYa3NcJV8MfbxDNH
9rB+5uNsTPsU1gUsyjfYho1p5cnRFdwRTNb9pER39VzzV+IxYDVX1rw0kXKENpjNT3kxsyqT1dWc
V76ahvLVSjyF8ThBSb/ooDSrxJhZyEFquHWq8RGe6OZwfR33XZOebjlWs5r/DlwburdTadx+reGO
qTKrNQzvFzzWbcqC23SVHZxrPjYXTaXeExbt5tw2k5F6+uvDMNGEwIyeCRh2iAlqT+IBnhR9xyQL
YseAF5c1freD5Ee51SQBle6porsGZSpVEIlnk8fLVfk2fDgG4hs12yG0OqPPSvAWMOdifLV5Qjml
ksnftubvNxkBTAiZdDJMT5RCOUYktZKEbqM7nQ7UMGY76a9sWF3+l+c6XeSVyOuNyMp6nKXhwUlU
aA4OtBYWg1b5S9a9o7wCx4sSx/hjMsa/Ww1iZ1P5tApYIc/h9FJvh3FG2xj/1hvhy2uihZ/1snQF
jQB6fRufkYYDOvQrnVRHYQqo3R9vnLg0ZPFCVUgWkfLPnmYsIuVmaJSIXFmjKuIXZ/NcH3MF/QbJ
NtygyjVxqpprCwWAjLPIJ4WI6PZd9NctaPuir311ZqBWndkSROFGVy1/mQWNKFKFSfWEYFn/F3mT
F3ErmRDdPMtIr98xPVmy0VnAkkJ+i4TUWB2KC08LWv4wdxUuX9sxQz6FA2FskUoMIGxgobpnnS1d
BSt4jv6hXtyW3SHcnMA+6plEguMnwUr79YrRLnrL+q5l81lrl73Xsu+3wpS/97VIWjGxySXd6dyb
30S7cq4F4KCarDhQeB3od/eGQ6y+v/RYFqKvoizTa3Gm6KUFLGrREnoznlx4QXU9LHtHSvnul4Ah
EzDehFhdtubtzFYm0xQfCAApmtoTAcZjAukXeDzJiT2hbY0dty4UEbFrKukaLvRxKHRa7pbUuHqL
XiDG4X5iAZJavZislkft1a5R6Hx8XiRnRZU75LA0ziERVx9cBbQWpQnu22nZC2aRdY8ZgHlwNGSD
pWXZhpRwHt9H3zrBbc+JdMVzmPgqv1Np0AjkmEgF16ulPt9WEJbx/2JtRhMmp8oq82yjrGU3CtQY
HZRhrd5EdyGRuKtIy8qoM6jUEitGbfTKi70CMGGRF2ME57IswJHq7XiEFylAqQrZrq/xmMomyrwJ
Y8hbDxQPUD2IeNa7fsHnUgh7RGjpo84ZFOk78LL/bYb9XxKcbPEw8CnlWJLt3BxpS5MLC0WgAvcL
SqxVGBv3z/gWDsSvbCcmSKsZmiNTdTfK5WY/vrddDBDsYPkhIIzO6XDu8WLZrnFs6j3ql291UrG5
+ok5Fg9AgrMNMm8NlQG15xuQkDZnxc9TCdXJH7Lt4U+ahSipd+0AKO3MDZoNQrNVciz8fOODQzWH
pAmiR3HwbfV6DhyI1wd/9brglhkWuX8B0lumIuAkH+0WcVH3ttILG2DoNKRApjw8wQz5l4K0IO3H
dJkymR9wdE4Sd5rcU5LSm2W1YG3LZKFwRvWBMwiC+QmJnUdoHVe/TmWkla3oBwWf0ImQwXFdzJrw
yc+sDGRjrrCnHmX6E8IFLbVwvVR1qk334kEeym+l69tr6QCsUC7AmrYbcjEjkAWRCJd4p39/DK3h
VwZikv3fmoGuhSA/4/wakOhEwZbzt/d8y+vaUuEEm16U57ERUctx8T9S38ku9zYfFlYrm3L53BEB
Kb/j09VpvqFpDP7agiosp0rLT9Rw6EuMtsTNV3nQ233I72r9zkU6r3KsEWtSCpUvLFh6t1GGH/C9
KymrfZ5gLIiAVBUoi3v9//wdSddbBrrGUyja5R6ej7dV07+Awl5Di6Rifn7z+abUEFlkdMpg1ulR
xs3Skn+uZNbBgM756LvngEiGipCQ7UgXbWSGSnm0G4w760INZRLCUjva4t92P38psSHi/65hjix1
FOLa37PVNkogPuBamqCFXPr0sb+oq9dFm6IgJZZaR+VVC1CJklEnJgoCBnyJ8uj4IfwDpEPje5Wd
RJJ0uqqh/u8y/dzTIEqOW9+Kf6B5hUEYjiTHbG1wkqMfMz7+r+SdS5VTjh49+jac2nKb32pssrio
RQYSaKIq4zhCPOQ+JehcjO/mSHO5lZBNt2XysXKMC2Aie/lmZfAezijizjOXV4VDmaY1wPlUwxKF
O3bR61MPTqw1acVdI+aUNSiFzBfdjRKYBA5utGJVUy1C+oAmoc1uxbxdzumldKvPaAy9O0a2l9B9
2nE6SAblqCZ8iCAJeAnClMbrYo5JRssHxqz6uCc++/cqRPTf4ci1p61qjrqSiC/gtPNrBtP3y5wl
j3iRdtvDuLYGqkb31zdn34jUINhyiff4pRki0lPXVSvQfGqnacKd9kRbkw304pMIWc7EBGFop1qq
31+GNwR8IM5JuXlL8Y9JCNlpNuIp2m3TYKGjIAa2ye7qkqk53j2ImVzeJKT0SyaJ592uUvYRgFFE
qsJYeq3WqD+XsTvFvF5Q2dnhF/eMB/k7aAiDQ81xkHqlM/xTNFTIxIXHrNA79+jxtNOuDTLQNz9H
u3A9XxGaQ6jmC5fA35Mh0lwyXY4soTP7+ODBxM1ZdDgTs9sFjR8qNhGMTHrw1WNXt0j4Hemx/Zkv
6jdSY6S32kMuRBKB4PBoK8pPMv2IhSw77m4eplAMt8B1tGoETizd7Pcetg0YBQi4mXnkhCnIwoj2
6Zk7d/zDxna1uYgzffkAg1HIYHYwRqi05qkWVW/ij1u7WQ7tas36SWWCx1qMWLkF/u86uNijP0Z+
16EMscOUj9QEfwblcVuL+atujWxbaba2csCGklgFJVWm9kBcLcBkVwGeQEzOpM8xBYCCqw+ugCFV
n3irRx5lCqrcAhK2nX/IdMFU1pA5ox31VKigERSLTZC9n6AdHJqcYCK9V/1MCXjr795zkoD5+yjh
Lbe70RknW0xvY4+vdddtKQm/MhrrRyFll9eLTdPpTbLgpCaWR/YV+h4pRodyqFMBn+zSLGJFypG+
Wj43vU3bzNXRWM07xNfx9PQ/y5zKk99uaHgVKFHrlu0tk4AlK8LSPoyPY1P1H5rtf8NDwn2+DKJz
QuEF4TQTRclCTIvyG6WisaMLSVGOiymzOMJyZNhWjE+stnZSCFnhNIU3Dud5laFDH8IpTtEkfx9K
CVczH5NspB8//brkJvv1Ntp1ynQEQ4lYzzeymAJ1IHhqQWEcumXGVA0ybyjmCOqJcFv1bL+5wGSK
z077I3b+5O//r/kB92xhcqwHRrBPumUzXrTmUsb7o0ervkpDnQm/tj2QbW23LATR7CosTa4U8NmB
b6c2t5Wxc2/rqF6a1PCyQ7hykRkJQbqzaEgha79k7HO284QplDQzWoZ1aIEHN+5AKCJUF9NoBvHq
m82CsPMBkfOr2go5pJ/z6fJ0qMhZKgY0QDvOIb12i4l1RnrXloGitQZW7DidvZjrTbKP6ZZRl/p+
09D7TOe0kFKMn3CPzsE94SHkB+QbOwwNrLNtlA6xg6OT2Sph16Nnjb3/C4Va/LKVR9hFQvdrgF8p
sSv/xMMP83vcC9224LN/ivwfHtxTysuy3puR7thlF/O7ogeps2xsKziZD19P5fSnjcgUVFxR41uJ
OYwcL6WTedHYJ1sOgXmaE4VChtChgtX6QMy4LxPW6EMzk81xKMe8UM0ERhsjS5V11Ytb/JJctq9t
LBUPW5soblPFP0LHzxdI5Pf3g4YdScsK21kXwvO/oOTVUMPpFDlEsE2lldBkDWD65nU/L/kkX0Jd
dlpncmTG6m7bPnrPLVwJOb+c5JIJstg0rojc4xfrt5i/oVxSeS8VCKcSDNBVvwhN9aGxoHr9Mg0g
Iozwx7o4UfJAL++Nm8YJJGoxqwkKOyxGMJYSuBLudD0oP+2/bmxT0JYnbIct7qz6fvS4J0w4tVEr
Bg29WxlyqFC09tdw+Lqw3MXAGrNA+SUV1lIYt4VFAh653/G0F7xNDHXi6cH6aBpXBCfhUuC5ohuV
JNDdRk9vkfMLBSJM9IUsba1MwBHxoG3Dxzn9JBxc3XNrajiAxHzFY9jvPAXLTkyMWJPLnxMfI7zY
yb7mK6mcK8JPmezwAwHq6B5Gqi7QaI9PNW7+9CvaFZ6Lc6I6hyIEMY6ryvwVK6MM5xReIKm6ZqpZ
98TAIMwtHTuAJLVfsw8iNYemxpZkEwVGQLPsXEzgEdn5RedwHXZW4kc+yrLIKWoVIghULVLsV5I6
MiDHgpONeHGqdygQCZrtuiiGA211SN+QUz8U3EAaq2nQoc6Wn3fjd3qqLMz00ppFui5/30vbG0Fm
kxDo5DdotBJJ2Mba/kuWHEVPQZAd4PLgwckyAL0duKAoZ94/xq3pFL9gcfyqaFXaOPStV2VSbeTF
uMrDXwRKDvGMJkeaUWw40NzlRQD5kaYn7ujOjwI5XoEoYMz0+WLYiT3T4VU6mOv5sj80dJ2wJEP4
at+dXA07cnXgGaIC/1HlQPLPndf7bLU4nEpjWKIDco5oUs9XacgPULGdv+rwodDHiIYwOO2qm4jg
i37RC8O2GNCvrYemKyIfestno/x9TdyL6MzZdoo3xNxdUGbFU7s3E4cARagHDCpjVoavpKyRmXB3
fZClbgEowNpg1N0ahUWw8fCNcVQlKKTytgU/AN3yC2LlYxglKHP1rSkaK5rZpMSOWnRn88EwE3HL
hVnd8hIAo/HDBc/PlEQGOvNXde0oOj99zd00IgUOp4Dbbo5bXrlfxjFC8Et0KBIFU/vhnpy87nIw
BAOUd3DLAe5FFcNpHVi2PANx7VQw4ldzVXLIck6wCZPfm5Od0WpwTv8HOmhIwe76cuW9t8jliJmz
XfCH7MnkrblnU048DZAz/lf9TTkYeW4jCLkpP+ErJwUkn1FZip8zMefnRFDBRSZJFh5VDIpreuAF
HW4qWGt1uuSCDiHEORMtaINZMKS12BH3IKdiIwFXqCXcl56m6qjP+ov7jpwf1QjFuvqTFbcyDi2O
2bfIr5Tgq1lDCOX41dqbnOI3lcHYO0HHXhg4opi9QgeZzajQTGDZ6xALS9fhHUgQziaUNIvNlwT6
rEOTfP3P9TcUd+EPZlbFxj23HavWpfcadnjGim50NhjdnpxCoAyh8OjFe2H7322F0okNnw3vKg58
1auGjg+Wu2jeOlbXEcmxVICzi03Tx+7iJqdnGfA+1dZBJQKa709jlIGaXAF/BZWhBn2JJ3KMAjwD
Q3YlYqdTgTYEo3zNXadkxVVUZzG19ym3a7XdcI/Q9kr1NYQx6hwYMDNsphMc/tMKkE64vQn5RfHU
l0aWn0K6Vm1Dzys0jg/XxXJzC7AG9OOlCX4Wgy57/LiDkVlla5HOjp04kyOGFI0SPAPKqz1WW04n
qOG6TxTRkEATp57kbtJF/axEg85wT5M2d+VlQBbaJh6+rMR81OcGZLzZ1+EhRNRv14K+nPwzguYg
wID4aOWudVmbQjaLin3/cO1HyELQ9B8zelXCpYoH8Q+OLrE+3BMdHv1/MQsvGU82irRIjFz8/KOX
azI5xEJ7ZWOVwLBjNmwU4c14nTtC9UUAq+1DVxjPz7IbWCXfLI7msX13o5jv8xle+u/IJywXVPT0
Mcms+as6OzPErA1MU7YN788gSlWbYo+9KJlcLAoD2fgiMDzc/EvSaGhdacScvC1MC6VqlFcO6ean
u31OO4RQIszYxGEodvECv4uDnV0eBrUASqo6DdTWi+QKM6wd2tLfzb3jLHMouIdFZ41k28vQEdSw
Wvj6qxUIoW16/gUeWbqpK4WljLCmWsHHyCPH7cLPRBDB9ZIgPQq1et4lzrWZOjeLQRY3YcF8qB+b
7SncaSrdwuPEN4BRMjWJ+kEfpcCDEvTAubuwW4cXeBJ9v80CV9uBp72FhpN41IiPdAXCktY0oINB
k4FDCr9Js7Y52ZrkRyyZsyxubd/gtYlfv7tMD862NDkENmOhNrdl0z9wzjxGfSY56XoFZ+Qhu19Z
fhysqad7KmD8Ix3le8lusFp2uZVmR+3WkVVxJDvrYoc5gT7MjhtzmdDdbXdyPjmnpqDAw3RPS01h
wP5ICoRVijEduUVnbuZSLKJZ/NoZwIfbzj6Wt9ojp9oU8vtk8KEw0h7LB263VhrjCjNnZS+TW3hy
eKGD0Vv4GC2pX7Ezv2t2TEirLEnY5mUrSst+CPzDNIxav7Xh5MXe2gowuyAKOjSRnBG7nUrW/gCt
zU8MTIXXe6sf8WP57VQWmPiC3GtlSlq6GiAuYNhtYN1l4pjnQY4XtJHsuSkB+b7C/Ogt6A+rOIfs
LAS++hh4GtKKjjArNig2dDpdiL1mUUsXYq8QzlmQUeBOy9OAjcjab/8/HL2EmSYz6SVExWhyu4i2
M/gdKUCTJaEnnOH9q01oTA675Gwh8/9gmjVRb7yKgaTxvVwBN53FZbcqEvNL/RysyDyJvwLPTYQv
n58ID954+x3kaJ93SXy8UBH5rOO59Y1Oe1LzkCIXc9gcacVrHxhegAVpgXk1hBaPMzsg/cpVR4Ch
lduZDy1O47sZKpiY2pmesIw6Lj8JuKSofwjcdYzFFd9o1HcSGm1Pww2r/HVfLzJfc2SJ4fvgmPaU
bW7JCDyulwqOVXPdM+RtiyqSkwqMjAXNWL4wxsBYOzIW4Uh6ppoe0NmCxrALH3/OoKMRtMyYEBxq
p2lrEmRLH/HCwLxVm8XLmozBnROqJgNekwQ0GEyFLV7JeH7joY68MA4Osv7RWR1SX5XK8oeNbG07
3cKw+V1HhUKWcdKnGaDWMOEJtrYYjgPj8B9rSqm/Ta+PJIwQ90NRFM6EXG769F4nKN/gt4zmjGXE
lBqt8I92FZo4yboHzNuKOQfOQxQ8inw+wcrMS6FeDr0j844X5bikEN036Nxc2j5gFY+ow4cycjhL
wHp5Ee0k630KCyBemkidKkQNfmmnZwmVdRA33N7c55990SvvslqP4bzMVixFjaRc3qGDlESyaVt5
ltdRhuc+TRPhmzWgaNgqTSsN5sGXHoNoYRGxKioDYNNaSsR2gBttrFVjx+LAURXddTlqrhqSF9JM
+W54BcdKWbA/6a4UWwg2+O0PQREp/l9vZBvHqzE/qPpqwYUAFcuzH+MJrJnKAm3PrhBdgkhux+VL
R74cFscxhjh0LBBPN1mbMcpBYYuzHE6P5iV3cR+ZCFQSFALXQrwQt4gFXEpNK/5z+qhXPdU0jhwG
1ThPmkr/VMF1UkSea7ZS73gcJYdZQv5mAtuR+wnomT7m49b2hT+wskX7KmWe1EHNzQtizkUzcKKV
QdoA6Hu+3ECBGkexH8GCL5Hmwa9k2b5pQOGLWr72vWxHGnt6dyshtDVK9ylK5cQlkagauJpPGpQc
81XcublR3P/UWZZct+Ke2VUZH3YJ/HmzZUx4K6S7iMu3MrocqDK0UnLl84GSCXTow0eNQZulcip6
YeMc/6w8k9gNRz2sRw3e7Mc9PN5b743BK17pyMYtzuNphkwdmjMy75GzUA1/5r7WykhGkjdmZBeU
JXdKgXDeOmFw2c1DokBk4vkiOVTZGbIulOWA2GtcL4vy8DKHDJHkjjpMFB0Tt3aITh6BNXqdgHuS
q+cP+DesARhFBv5+9ojIdDc856FQ0uMtuTAfonYY9aJSeMC0AR/wT08qierqMFAgyvFF6QcYvNum
igjflmBLrFbXC2t9M7CGolWxC+GR0YUgVFqqqYAhN4I215RPmKUMEZ+tL9jZgaPDKx3IuWpoAAju
iOST4YvBL+MP/mTaSDhYX8DtXG1/ggDZsUvLVdMNf293JWuFj10LuwGV5OrdYPM4iyzC5pFoCsTu
w+JwtEBk2/7ynA3WOXe1RvdGK5G6VV6chzV/2Qezs+s4/xQzU3H6jlqBxQWpGiWrEOgDSBKYiNMy
twhnUk//Cp018Jp0yIwX2M4xEPly7nJSDxFjxJ9YWMyRvUJWMD1HsIEpl1lt3cuRdtvpJsNuMtg3
YdMHNKOUf/MM16l58neogr151qXFJsFEEbYmZ858GqcqyQxx3v1kSFfcc+cdQqJjhfxhVTjnAkPj
2lO3YB6b3Lkt0fukCB6Of5Hml+kZ+pgqYJRMcMsUFoFFIGEI3AucRYxvuP6kkeDh1vyC/0JDdqh1
16CjPKMYp/d/3GKtRlQZaMXe/Vp6609DJ9VnF/Dw8qU9EGMzWdewNq6fErPr1dgJprEkuzi0rOyd
eFrP0FvG6qO0dp4IYlagaMRBXAO4ioedAQefGMR2u9Amx5/KpxJwvGqD4S4OwhVfPb3zUJSvtmRT
ksE3okHDqHsUrSETQUEtH2SlUvCsEp9UkF/0PuUUD3Trl+Al+u4wonO07uIYcPn7EKA70VKy1YR7
MwnpmQrUwq6inTWSvw7cwEmtFx6Il2IDEvhwuYk24ZPCQ7VNHshXWKr0VYlU5BgGqRueWWkziYnY
P2RRTg9EtKEFg8fiEsOguP9dCVwe12IrBytCT+/ZB9Hfn3jXVLkM06e1gUIJAE9IqSRffWygbmq/
37cEJ51H77SEcmqTvKtA7aJNbfmtSOpz6PYjfQVy41X01YY6h9uI1H4rwurztKaE5WR/E7IaWjSZ
brwRl+LP7/n6jNUeGDaJ9wzUsfVe7NKjsXUWS7ysqWvQ2XyFA5lk3HDHVp1NhU+LuLXKZ5RDPQdf
dDrjFMmvKOnoEmCVljgf2CCGhRbMEaYgO53nvAELdfvj1RMTlcgPBSHzCL2Jo/bkUpOi3wZGTv7e
3XfTvCjHAQ12p9pzh88GI0S43TejhWeE0cLsihUD4OiSs+MxkkVHGho4W18vhEZ7VCpoZCzJUtZl
JJTixJlSZeeQdjSDMatoR90x+G03NQwMIGcMFVJ5VMJb075Oh87MzPJZmI5hstkPnfqfeqsnHncN
HLPIYtISMSqi+3Y2sOs+B6nkVJlwfLEN0Rk3DuBOH5H+a4SH49sP/Vu+kM5K8zBHgJPXiGiHX+HV
1XWjZfSO7R5PyVcs2t+zcolr+PdG7RrST7dZZJ2zsuPQifhJhZhW5xHK786iyrtpZDO4IshFrZSG
GROx2FGatMzucDQ64UEjXAO2hAGWp0jz7vwU8iafb0l14iXgKWePn0zozT5/2ZZMCADyyTqPJGIi
CL3DDFxHsJF5fMNhFnYxrBs7sNKNe01EWwcBM9ym3wkCx3ZtnTp+RkCgrwliD7+zy1CJq176Bo8G
p75NVVBPrGZ2KoGkZnPjPiPdV0fesY39MrTJ+9C2cofPLiZEh4a4bRGglryla2XdFVo3VWdLiQ7q
TvUabZdbGHV0kN/fVf82/Vu+VlSiY5hw2cX9GFy/6Z6TAKo5yyYCgB2lsiA03vj4rJfmYvhN1Y0C
u0cx8FxYXIRH6aVomV/mImBJoJy8gr1HmR+qnUjSdc8BOh+uPM1yyfKy89mDMshO+bsthHDTuswm
y9+J75YpRRD4UxNYbgBTtMgm8xongq9CTPGR29lzcOZkthC1IhwT7sfdDqxNn6DF8UJVnYFrb73y
aqU70rwnwA/hJTByIxEfbFZWzqPsbMij1TqMlKpPCu9rH0wdZhDDm5AduD/JOMU0fHwO3FoKHOm8
MH23Hn1N94LV8fLPe8oSLIxDpOjijLWMqxHXczl3HrGUuQWN+U38UEmFFX5vucScm/48WZiJm55Z
ne7aALqPRa9FdAd9qJnattMGhqYUgzvOa7j7q+YEXnq+LjC4h3pVTUg6SyOp9o8/MFPw5oHqxoll
zhqCpGOpu6yy3i60y7XGrsDc78jJsBdAz0jKLhl47kvvUHA7UUrgAjqUg8dpzmq9ib4hF2r2ldvF
WkLotuY5Gj1Z+3mRzDGADPkC4U8bM0O9MvMk6tNMVKOu7Wkk+M9jBJZlOEIk6wVUVrLL9OcdX8+B
NQYvhgsl5DzsY3vqmYACs7rxi3EoZDAjnBl3N/47PtywTAZqF8JDpJAZdctE78TY43cSuGySi9zL
+7bh4lMy+g/cyV8fvpqi1WasRDJG8gOgTCUhFyEHwwFW4AM0aIB+xJHbTMZwORZ42drV9rWjXZ+U
TIdHfnl2AyRwhZsGZ44PpyoEihgpWLwsgud0Bzw0Wo2UreMVjjCThiwpHRC/t7Pns12xACqSeoKk
STWvglYm67HGom58VkhHNzpx/RrBFcCP7ddhycm/FniELu6c5rTXhnlfr7RZxZN70cyxtHt1+52I
gNKzqWr6bQRdQ0PcuJYxg6Aa2NOC0xOGnKTrsBjG8FS31SY2qavgZdT8ORlaFmCLXxCVGQCaUvOI
L3Ler/LSNEMhG48/+E7RqELEo9dqxi4TTDvs9NdvZnMSoYpXVwPfMgkhSBybBOcxJWI801JMsjUb
et/t4aEwkJg8uGnbsPjETw7XoyHNXwwokXJOLhqDvZezqg0Uuk0ynzhPy2Ht5XdLTbpt/zDMy9k6
LDQRrnHQVUI8YLWZUn750Nf6JJ155vZwCTGwR+hScHIGf/7dFZgO+fde1sgdyu0vPkEiKznK8yX8
NoxQj2CJErTnpX+04lUTmdlQwiEros6mToiDTlKt3DesesHvfv5QsECJ6sdYz/n4NPe/fpEgNr/S
yn2aHKr+8mT21Zr973jC+9IeFm7N+ypOPfNWM7herNOMTQCO8YP0NYBhMxOP0vtJ7ufBgGo+JOlR
Yi8qlTWsNGQyAsi1j9z6R8mUEzcYT+ztr8MiaHDaWFPToD5HXp8Pa/TizyOtGIkujCPr591vtWMm
pAh1Ox+itfpYrbAMAkDk4vXF2oSQ6lNsDRZMCjNPy02mc2v6+/x0HDXslyl1WiDM2CkxD0FomoyH
XzvcYuHA4DhCCbY7evMKIB3SrNbzDYwwXmW78v2eq9p0jw+El12m8aLEdQwg/XTstVwGRyWpLa5Q
Pu4BlrMBDE0i5BZ3x0E2PXMc/EDDr6cje9EmWcetVMo8WUoEM1EKXq36ZRqWdWuRQVfhQMbhIAzn
8+8qv6XGV4teY+frj2NBMhk+O+WEV3qohNlWuq6/HF4tG3cnCM5jMcujA/D4cpSwuZUZlhNi1Rgx
D+qZJIoWxO6XwXMXk1eNljl4sDZL6/SlDjS7NS8A9PQ88+sDtYlAb/bZn2gkrMhABA4rvpiT1P3y
Qinv9WdP+JJXU+KmSckq0Tt5JKMQGvA+FLv5+XDZRHmEOAcadjQe+dynZTrPtCLOdgd05J8yfGYb
weahxLDB/7qL6vQ2/Lu2881XCAxIb+YJAr2zAn0Mw9dAq9iqPCD8sc3FvrjDmYf3FAEWr/C2oZ2N
CltfwmY4iQkqUdKOy7F0f/L4C/lqDa9UEHywVRpo9fSVc6vNPHDFNMlHGmXh4KIx8tlxyNFARjL/
JzMyxUDcSPlLrGN/ZpEdNRYl6gdq1uYO8ccnTnmqdAyjQNWrn0WdeevRdIZQJmA3KW9mV8PzXf7s
e9Y+fqSvHYSsq37KfTRTDkMLzVcQVkKu3fE1tOJZr+O0bXA9SkSWUmxJBI9IzZsNQBZHCAu1rldQ
ZKBXHkgUEgBLQ01KRwRMkNAcFanr945NjnS6bI3jpFSbcN6tF0D1h3atIidxj5Z6JuxQamIq1aT0
iODUcLpNO5erSIY9BIAe9ebGycafAR3M+QzKd14JLveNLaGLN+gc8BzTNVlYMiWLa5leiRHNAaGK
hrFjF5CfYe1bkznGyzp9g5CLzfrwaE+Wst1EsmdnOO5LTDW8AgLP4jsbIQiLke1MI4JZ+DFClxBL
6iZpFY3SslN3VewO37sIeHZwl1fY/ght24MHY8EZArYEYfXzPu6VPExzM5u4CFiqWyq2DksfeKzy
8tdhwOBogwtPKRWO4g3SB9SqD91oyAigsx0UKk0cHhWe1v9ut27ln9xWBR/Fhx7lhwvbIRUPuXOm
cXwpi8dUHt3mju4UVu0or+PeXOzOkPMqZilnPd4OQ+BTH1f4ADZEgiv+PHDBpt75Hyk4ePSHIhUc
wBt0Wm7mAaboBWBjGiL61shL0q9wZUVTJkl0XroYRuQ6jsi7aRZug/lDpdCI67YGye+cKCwIUILS
eYajnSrTPeSYfJk+j6eijNxYgju610MTKLMHlA8MvH7AiF64V/TGremd7psHjJ7Q1Atn4zKFfQjp
TFRtbFmiGF/FP1zp+Q5l0wk6+PUkKDBKdh0U3nawZMHzuGjeA1oqrhPomfr73Mpu4RrC6ILsgoWN
sPBPfVoGIBGi7uR0h2XqZMJz4ByZiYEnhVFud26Fnh26yGtpa9XcAVUOcpD/0Dhg8end84k61Abf
VsZyyo8u1m2RmJTKDTtBbBkUmiLxPAfhbQat7I8Oy9gQP6PlzWkw5EJgnmwBwLZoNBMxMMrhidqC
BiRfTz+MyL1R6bWXiri7vwdp8a5buUlKYPURr+NmB1rxdRhFiH0YE2lKsTFetwMy1vGX2K8HOqYf
+8hQBZwM8nttv+UyZnLLKqlAkPl6QIF9mN3EA1V9b4D4Zaku/SPjw3HFxB/8jo3o4ADI/41U20d5
7VGtf8ZKEaqSt05yDDqsML+GDUoz3rjGv+9PQ1e73Oj3PEj3uc2sLqbzH7WVz/w/9VUQpNeHVwdt
QROtbMK3hicTnguDvXMYZqnkBAbLi6muHCp9Yj5o7Fupe15ybLkGNwyUNt5ITV6usl8pnQEEzaOT
zE8A73cMHZaufX3nbNAYo19MBL9Sh8rv9SHli2sQEwwUa6otbv8IqyiVhIc25U+7voOATgXDfRzH
u2JyFNUrh/kNH4RGvyI/Jg6wqx+illYHmPCWTJrgKSsLR87nCjrqQq+cpIRKuNlkabkzq4REsxZm
OzxS2i3vxXywWilAzKJMVsxPrUhL4g+o91Fd7JQ4k4lcDb6XdzkbaDjlTlmSUxoqQ6+E7e5t4aPu
Da1FhRML471FnToc+2nKNtsjwEv9gH28nkV5z0hksccxOnyiZIJKZ9ghTaG84CGYyrsPgVAwNjwE
ARbMiYn7JXwT8qFdpGQTGk/KGQfUURWbtbnjQmeqznChbqg5UqCyveiz9M8fMjT4IeRXA+YIrDw8
4hChlrkTFJK/EhqkYuKD8Lccw2MBRHeltAs2SvrthAeM+1lBhmWu14ZBRlucrQxoK7a6Li4XTA06
Aqumy8U0BVWyDUTuvSqhBdYO5qbuembJrhEhyQS9/VT9BtO4H0hu3k26fJax6eQW4gnWRAi7mfsr
uZsEUZAla7grDD98Z2C2wVHQdT2+F/3FWOc/IHhebyzQe2CtV3fprE+lPdo3LrU5k13brAKW74L4
OE+cJ9piev9CYE4i2DKv2dE7UiwdnXtg+EH5AGgFCZ1G0d3VNZI3Rfa5FisZI86PELERr0pbFXM7
Q8dqRS6zNCfWWnU4oZitYtNKRGzNuseHqkuYzShXZjthfrRXf7xwo8rwHhX+pz9U0Ha2+dcE/h63
jyLWCI+2PVKvfxDjEjfO2QM883OczDCHkI+SqZWMGBDTsIwgRfUWdlPvfHd1RgXHFsGWz8U8Cakn
jehSh8jPROkGCOk1sI/YVoXrL7tiX7fGAshrY00ZiQEGfK1B2fKgIhGnGvQQMhf4D+EHN7pQLlCG
P1vFomaUb6CqIzmhryCuh80HplDainzVkGfPc9o4EVgys1ejkxq1vE7sYyY55XBHWcUvIm1F9y4M
+pN8jLkQMPOt6SpqurynF9UhvCtQE0kIXRGG82X0BeY+B9mhfdKNs/nluswAZjU27AIzbrzQU4fW
plc55w5Lxe00F8aFc4f+7NrT6yBKfl/D+C6I2eRFpfMrSEVfXsQoao0dcRt57B+J3LvpLWzhIqm1
XrGlPpqCtWp5cc21REV0v/85FCUcSRcYsmLx0v2lJePzdCqepsYAx3xAasp//6cfyGU+XueZzIpB
c4+B8c+zgelraN/VkqTUNvdPOVltAY/Zp4Yue0i+Za/eol1ngFH69dj5GaQwRBDgc7zlFfsKKk5M
B7B0DEtry/wjIfcQoxG0bgBZ16/eyrmXRTcpnKUjqL4dv9r3vP7mnx8aqZzRgN87fEC8hZFfavpX
TsOsVgbEqeY6RkHKR6y8VHit7t56ZtXYMMdtK4jD2UEYxYvQypHwP/t8bhUpOuVpyMv/7oOIhMBM
TUEc7lYfqex4LTCvYfXhOJ6ZwQjl57LelDC0zvUm25VQurUsemMfpqrZc6hWEnTviCx3z3v+rT8l
Z1MLtyLdh7rNy5dObOR24z3JM6uvqk5ormra4R0xcUfMYft/iCMLnfmGs5KGO2axT9/tH42Pi46z
Meb35KiNEhgoYXWicUs7uRkGrLPdmdLvxdULnqw5WXeNRvLUDaw4z/iFIuPhqwk0Ud7GwV231NDj
kYhwUsIMJAe3Lu3cLt6iN1qTuSC+NHoiSWDJm6/ARMO75ij9UiukNe0J/paIPJz1OAJisv0FvUYK
AOEEWJsPa4cQxpFe5v3l/AItngPssg+I4I7XkuoBV1Q8rjIwcf3doSFwcGsr5v839ZoDF1VJP79O
DUVo+L32GvD19oOt5D1AGBZ8b8QRm4T39wk0ozP7+xM2Nwgi+Z3OmUDysR9dvQ3D4bl5kLptgUEp
EJswtw/Bf1vnT9DQmn7Pvl32w/Xh9PAPcydcMaRX9HmnII3qCyxvhVARA6H7SSxnS0dlcBxeya0l
xH/d4Yq0vb5ogJc96m1KsBcJH46Dsvv0ijfPSydZfvEMuXed9EatL3AXPRhLarkUergTuT02KQlP
/W2bejPm8Pzifhul91l70940kRxLAxz5triHEFVbhjreZ1HeoICwVrbahqvYBXeJXDA9uiv62bA1
kXmGw+6xfdkw8QRDcn+1TBspMxFv7agMQ6OYxvWk9/w7eEsPtSB9b+w8IOm6ERK/OtfZCgoTZnxt
DgmDuU1M8BtxT4oGQ98+NNLrqb201rpJQjyxDl/02Bq2MilTNId4J4T4/vuyuMH8kYJO7ALl+PDs
8UCDR3Y2T/g9Qh8f9a8OZKQHJGqSs6O4qLgT6agWwoRXakji56Sq9qG3XKo2vIDuEj1AzmZqyEIf
cmNjlbc7EbMob3z2m7GDFSaW8kmG0hiIR2HagBG3sILgTo9MYtOgwbeTEzJYkNxi3ZvoGa0zdI3R
jlM/VMMhJvrzQ931j4Y2jcWbT6mltw3X9uTJMzKRkchmYS8s5rwibpLVta/3G97waJVhlSpbQm2A
uDGoV07KiKrPv3xlGBxbBrJyVLYps2+TOOh2JVXphsrJQADUEn/tSsBOmSPrmd/vmkeh/ZUCIe73
+ILl/8xAYj7VaV7p0aBWt6zQC5Gib73bRZJfPUOUmsFaXF61PWrapkiKB5+UwIE9i6ukCxLZojPC
9zh0udY5GzfxnbaongDu43/MxENFuGZpJxEY7kPuNW8YDw4Q2hMgn4EYiLoNisrVxIh8aHfGA6BZ
43+akBku5Xp2Ti2DflZCtcmwCgxO3KC0UnxVYNROSk+xxp4EdQkJZ4FGzDSqXLeb+5urWN6TSvrq
InDBK8ioJbi7/vO1gbaxX+nCx3x8o3eKcELedI16RC2ZxCV+evyH+vUieOYPJjDqfE/Jwu8fI/Km
N2olmT2GdAZKc4jB+ibOcrs4qyjn7uTXPOoW5qsbw1Ypc0MDUn5S64pVUQQbDU+Z5qoLP5JQ37j/
nOa57gC88rjW9SnwX4/NTjFN8ed3djZB5RtIgQPyAWUDkBIp9qcmACGm74jXiae6rk3jqWWBP0sl
Z2f/fSdVY9URi2u0WtsAS3nSMsgs8fFFfijaTgSTVuOSlRuuDV9zkoKMCu7lu9AGZBrw7Ch+gDgp
dUqGgtfdgGt2ujiTODnkImjGZQpU174mSZpOMgSpCWC3LNIjmNTc31JKUBkaCYKJS8mX0Lu9wHN+
OnbT76Iocrn/WnQaKWWirBbYvXrWgQ6IPeaiU/CCEZmNCE8Ahi/I04wIRXwoI6oF866NT5ePhLcf
UYfWDQSjP9coNgsjQ31xtWmhs4Z5dKIm/abtMiWtLwevNli5kTr0TkNN86shXAJecZCiVObuS6zg
iaJkwkFtltaFsN09wDgIgyx82dSpBgXMzJEKowJHwnlIYARb2oWHvUw7nzH1KGir1+azAx1JBXcC
ITB4oo7+dzhl91sCL3XLHyJXXeemcLgtVfUVsPeihJSRSdTJxQDHRGqyBvIrz4M2rNfL77PEPynp
PeBokpvINwIS/zjvMsQ2+KbhG4vtQRw1DWSJtreAQpyN9SjZXYlBBfbDLLM+wZE2L/RVILwiADOa
V909+Rw7+20aGTJDbbaJhRsbpZAWnSD1dDOm8PpD7ok1wwnMLngYdNzXBGqWyoiCJozJbgJ/VNTH
hMRMgXvS/Trzr1QlO/jDV1o+1iar1ke3JCO7l5wwF/sXun8sC9QXgyncSKVzKEjdN0APbgQJ3jXK
nBd13bIWfQZNIVGefPSgSQ/1NmQBEX4EJV8xT1GnOFTLPsBqe0Drei48bqgp1VU7i3+miuGG8OS/
4OyeiyleKfCDU3FQ1wtsJvj2WsNgGfYRs43+8fwn3bAOt8UhJ8gT8dAkhKpaq8qCPtoXxTAd9086
Sq1H0qJJ1AEboQC1TJ/ECimVMXU3G/WrcZ1SPiiwwDHgRTN0DERljRQ42+pjG6+5L1fGrxkgOAEz
mJDFWB+YFXoax0t+0Sw+0N8XcNdzWvy+MbZ/DVKuuJFt20yDjflaYJVGLMLcvL+q1Vpy8CEUB3Oe
6CgH0gH8C28pjDolYygm+5ow/Ipn3rOuszYdALEBULv1lQtbafI35ex5V2wzL462jS9FwYrKr9Hq
NLjI9RI0f3oWnoO4XuhNaZofetaFeqjPS2gatHcv3g/D5rDxJRiKfRPTNJR8LlPanHJ4PNZmD3jP
ZNyIQ3RaU57b1KnWRtXbrJJlFwnicyLx0NBjHTMo8npUDVMYppdp28yJ9BCU2r7Xd4h69qrR4v+i
2LBi5FrJwW+u/slB64343vpP4TLPiz2mD4xke5CRHrGTfGHyfDV2/0b0171CvsUuIJvR7np3ejZv
xOYpmP5UPhHtCJgQ/AQ7pfLEcndM5AltB3dtImjuChcMLOcsjqqnK8Si5EGuNi84sjrUw8uCeN+y
klLCv4krtGGIxQ7XuSDn628NFzwtfvL3abt0LvTYt7PHGUENf9k6MTVX2WYuzcDCT6JLC+9DWiaK
MejrHK98FfhAnU1eXUgiJO1YZbOaG2g4uVa3vVSyRqhiLr+9AKx8gSNLYGg86PZr8DL82jDJRsnG
B0ASZnGSRJRaHr7WrwhOJZmrI9Cv6z/2L1QzGvLBFOH5sdv0PYcYtSSbamBki9ZrM8k0vv6EGSH1
whjvmILmTaBgZE+rqj/G86H2jVGsuqw0TxPOF0ILMCBOeoK792MvItsXvKh7G0M9QMnflJLbXz1l
Nt2o2NY67Y9nWZkK6MX6PMZoWA8tJ5tTmr8NftJfUeBCc9SSCtzNuTQ//of0zO0cPipxzHC6jcaC
pYIJNOE55I81AO0tEXIj+9vS5UwXScfpiwZwV939kwGEafD28iyf0uefvKeYsEDl0oF/moHW8qv5
qO5j61q3Tt7k6CuPpGsQhJTNYrey/PxjyvHCjbeYOtniC60qDdLJzTgnjdp61QC+uxzgkqRxll45
HCSxX/jKmAyn6UbrkNmD6yuw8LlNjEXh7qdh9U3h7NMQy5q5glVaPcbMyKAwqNy7UmZNpo0ihTAE
h4s4KJIzzuAaIsAiyQjuWIsRYOjgGLytcm2P/Is6a3WlI2XjQIABV3jYCMhxFeAZjv5Grmjpd693
Ek01SLlM3QHJrtdI7tinbWU1yOE76ITu9oJ8AnloGz+LbNKoJjAM6yhZTaaBPVxK/748Y4OLeQ+R
WhTN2VaktxcQkn1P/z9fBrQ4UUz4nFaZXuf4IvO/UiLNye1JavqB+tEYhLYcjsll8KBCRJtHjwuU
dCgtvXMmAJpDv3oYmfgkwHHlCATXBIhmfsbo7IQPgU1nxG3bZ/84Z79IiU4L9dAUcRR7Q85bivcO
xJi94k/Sr7pXkcFr3iDDz2u3MnkJVuwG0real1kX+g6k9TWToJFsWlkvYkf9q2oq9ROSdXuGaPHW
1Vhn5yVjtKnvTShr3RhGfp0KfKTtRiH5ouqKRgsv04YJZsSGaapS49kwpVAI07f9Fc48DIqGpfpt
ayJ+HO11wKRyXaqTOmMswcXMd+ulmHbzW9XLwoYdiDgMvwux0Ev84hJzp0KvVjRoD4R7ex/Bk0Mc
MoY2LfbAoekPd9iT1uxH8jfmOR5MQ9yJ7M2H9J2N6bWrVAxnUvwUNwloaz4UIQUhdU0Tj3NKqr6P
IIukoQgyt1xQuBBJvtzDx02CuLoqnFU044KMOgFCMso5HbExlUmIdvAhUdnjdC194Mi2P79lMQ0J
NZciup/gYzFtFMdBKFy7rOSkagiVIiEmEdwKoimhmzRTFpix9SWmtM4XEHtPAxDSbv6MQnAiNmQZ
TQkBQR9fOisgFnNOr+rBcJJjoHfvoUZxWIqBV5E5kx/3gPGnKfgAXDPOPGktAVa8JTq56FNt+aaJ
NCy4dqj3Gr+18S9xKVUqLYE0VM2j6K+c+oPVEtAlH0rCzj6dzZo8vOzxBaPl4kitWlPmqVEsVIBJ
IHYqpbRTxPrSU/lKa27nPZ88p7w+nJYdoxAUD5ubA2H6OHtZTDs5ZHOszYUknpC/q9UPgUHxDlU9
GMeFvEy9An2Sh7bPJPkdZCmFEP2SNc/8NtE57uP+Vz37ucZ/vH9GtSmhjgHFcdC5DVFR6YTKP/se
Bq/5N+I6YAjTpWJDqp0CwQC+z840Lr8qdGjCjbpDxG35yQFmqGOtC7LrjU0jxWmGKK5HfP0NLwCN
6s0i7GQqA8lPdyPXPWIQcAdqjF+R9QGPcgMaW/ahEvG8zFIasS+YfzIUXveN/Rm9qLjNc3iFMAqB
LuUML+pGvIUEGF6eTrA6/fgGOkevMlJVFscAHAyPXc/XgyFBL87IYXy69eZSpihybAraW+yWKpQK
5sIvRKCfxI56vBvAtXkHtF23RC5wOuWknAN3Y2f5DsZnWG7xIjBb4CP0a/JN2298Kql6uhVZ+h+J
o7747ozc0+0zIO2oFLX0ya0n+finGZO/dqD8Tr5yi0jL3qhCsH6rdjRl/fRzehWLAdM1za/Mbf8w
RmhUNACh0kcfkEJ5I9nwe5MDYAGkumI87TJHiIuLD6CSC4u1R3Z8Hlr+jNWNvPdYuS+EkjyoJNiw
iJkxyb7ZwJMbbgHKrXF4/xgGOc7q5YjFXh9/d5DsGM1quVisFyiGYFD6RAAkTz8KwKq19t4cKHWw
DEd353CKcz3mGU/wWBx+0JT0MXuv1Ze4hLyddEaPx3Nn2VhsNdOJ0IgqdafK1tvqImTX+L1GUBa9
RtcDsqra4ag+M+S5JT3w0lAvuV+YeT9kWZqrFy18I9i0IT4Eh54w3ePfSxSn28u5wHERFuptEeai
d6Lt0naneG2borDedGRapT/ZKVqxJutuNatZJV7n/0F8EXiqS3hZMGzeNp5EcPbuPOsLJSLri225
HwNMFeQiEx/u30gt1NC97YoF+I92NjOSW+CWqoB/18VYZuxykfTt6YDn7QauCW/l6FcCN1NmMSWS
fiRrvjZCd2ZX/he8rd6CBkHOdiwtQHJQUgh9tjuPgM7+W6WUG9PdGyKbt7Uri2Zdnw0xR3i2zJW4
r8zEDN1XsJScZYzPp+fc7FUE/1iTMl8mh4peA4hBcy9jG6BeVKlD8RW2dbMryoSO7yJyseBDVVvh
2BdV+IdO+OiC/vtyWBAZitIsdNsIzkT7GznRrkr92eLAxBrYtmeK4m9/pO7Sz3TvP1ZQ6+Z4Vt7o
U//pdV2SH95D5Ly11qsYAphEv8M9A/H422T9eRA2vvwE4g/Zx7yO07rqhhgR+fPVxOL9zBCblCRT
B1wLE0Vc51d/Vsh/RVNXatvfbf65vf33anwcQMJl8oKhk6+h0qPWZjGpxn7KkxETRde2zLERZ0aj
He6e5Uw9KB9VM0eLUTUDASoiVNloZBn2Q8VHmhFNq44TGaA65LcxdUfF1JRkHz0ZYu3KmkzhSvS4
SdkWkyOC0eD6mhKKL1hsf7kDz7Wsww4+ue0q1VkF0syvct6mXQKhhcCaesj8jnDqvvIkAP2mQYoR
GmKNdaHIo7ElrbhffAcxc2f+HkmLzd1NQe1lZbzlnIwu2nZnbZSkCruzob9aL0gfxmN+q5JS7Bmg
M+9m6JD74NVSj9AiG3NffeO585IwLgEim6WRYMATb8iAzGtH4OP0vNcwL7uwMpGM7IrvLEu2tj2g
73OauFp9bixgOegRex0DP02Wsgnl6rD/AtvPHLh3ML0z4tBV6ZOG1V6KptB38AGeFWMoWtgmmfX1
m2PQ/R99Wm1kMl13WpV7NpWQoWuCS9WXn8d6v3xzbyeBo7rcd40bQ6tXSrMqOrWrmB7nyGJNx2mO
TG7a/0/uwqhzcQ/tmJmQeFto7XZmok0eEk7VVT7P1WoQppwvLXn6G8AQZiCIfkox0ZIkP4yh0XHe
ybSNaUbeFlE4l7BAeaumYKjsW0moxYv+T8VWUeXFpb/eygsc4L7IS6KWhN9FaCR8G9vjOkRUiC96
7ZccX4FS9QWqOm6EN7//YUYwiJb6mLAGQHcABRBBLWKfKXCvibs9Fc8DN71WfMEk+mKPegd3Worb
aw8Gp3DiILQo2H4+uxlsaV2m4Ybng9ZaLlmKoqzLPcl1URHghaDD7krfVxL/wge0LZxd+ZDckUhh
oIHAa6OOb3MQO9C1jhCkli6T4vz2fWWzuomQYdpgb8c8hK4jdK581YNy3jlinCs1imh/YE2OXnEY
v0uxfKJjnjeQUl3fY/1qyxe6BZCjb7isl6XnS1u6H0pVPwQ2mVi7NRtzld2wVPyw3jYx1IwLOHbR
k8+TEapaxQGlXKDSddBLmRlp87egYBdY/iOFA5qNmBWvJp10SRdf1TkHFbbpAYGXnXk3Q7sI/CMP
6ERgInquUYTqTwemAdJf+H+Dl4LmpTtEt7cQrvu160dVgZma/1uQZfyNpu5kQ0AxtLREi/cUn3VY
gXHmLd1KFPr3HBUm742eH1ZLRT3amv7vV9ncdQLGBzqYb6vvZ8LFn24gLFQDsf6u3ND1Mww464sQ
8XT51JzyK5n2Haktof6ZtIK5nrZ909g9ix8hQ8sjYQyp7hS3kZkyZ2Q3UyzUdcp/XUNOa6aC/GJ1
/x2rKDrWNDeKHiD8vvOYopQcJvGbbvZDoOK062+WFv1VvBRlP/eROdaXK62fsGaMp/8rGFgtPUSm
BkEQniZwMEMg3ebQDSlqIxqYTiN3XTXH7YyC9uycPTN2bUa8qJJWcq5CDh6/psDjqij04f7+aNJD
+mXqZPy4C/5+b86qsR1gnDRoyH+wEmSchRM5N04+1heQokyuLsS13t2sMMwiN/QD6ewCl1gDGAvN
+TnIytiwX9OKuqgutA7ivMr5JRgPDZroM/agFxLYdkQAMva17aWI+DVcLWvSoUbf9G3X02mgLBg2
yfxy2Hd/WvirgcjafgQDSebcK8y1qksC7+keOWvu7Eijer4guNipw+iRyCdT00og5yHX3V+FkSad
12DfvhmaxKR/GTumS2NmJMXFRogiEWTym5Ppc+j2fMAt0kIjs+Jul9sHLxumZ918PdehAkFw077f
XR9Ms2l3EogeskJyFj02kPLAbwIFmENUAQd3QC0/DQJx6XLIuFly1N52EZeVFJtiWczmDCbngiX1
4aP//SLWLj8hv8iusgH7Epaoc4mPeuY/iywroZ4i+UOUpyBP2BB9Bf1odwXbId3xU8+q2gG+RdlG
8G7AYgT/wY9FYBok1wB4OzA6FbU/veXuFMeKfr3tlSrw6FMmGHGk7OQDkj41PGP2nJw/GGXWKQV9
GbxAWn2uSzGBMZiBwMf3C45AimA4EtyU63sSXRosxboV4G0FtB30R9KsphtXPicMgRbUtyXVezkO
WLjFhZeHG7timuZt5UrulrfFYQ6KET5P4CGLtlfd+E0Ta/XdIYNlFoSjPQv+dRQ/OoNgGpmwObob
4m4AzpJ5rpuc52VPFSik0sOXBcC+1SWRL9JxVEjKUXvBb/LlUXj6pP9fqmefk9Nv0LaQBSpzPkwB
ep52bqEfRfVmgYSGB2+VV6bBffzzomQ40yGQTOWtCyQeJ8LzRp38YIZw25EpkgSOnS8/VkXb/V92
VIs2VmYUUyBRJ79Pzvli6DUygHq+RcrgRu/k/SmWlT77l1dvJhGibhjNp3/kjnnxFsjhlcUx/vE/
EOcpW1tNkljs4IFk+E8BGojSN/nfrTvhRNv8fNwkZGXS9Yxh+qS67ytf2YRIYHhyYKYgCoM6ig0+
QJdRkGcJ4Li/VPzyL2RlMBdK0x5Hbwq3WboHjTmbs8hr0xv2iGzdYh8oqPrWjL5uE8IrtPyFHwiq
tAMSs4EGxbbSZRVoEKEGZFJP+ajmsDutaFeCDmwg39xlV4uvu4tEuNwO7DqOIcOQV+WZ91qaCosm
AfDOuGA7JYxMxFCnwiPNFLBpGGj1uHZMmHlYgOtMq/JUcYK8RwDShoegmPMy7ImtNj+A1aPn6E+P
W/TKR7jh5VgXKNs0gRnhytWdV/Ai5LtsYh8n4cNyiKef7TeId/x+A+1JJt1hs1nMTEEbv5e+RJ45
bWJQfh122YSZghpkG+pjN3DHQskxwGMYZwWQOVNYKywKItapkpeDl3YGZ1cdZNVSw20qEPzcgitD
XNORNbALQ8+/K0yA8PHLlkOcZxVzSxTIREMJANDGbNLpp75dP9zzj2L6r/0WpxtHhw8Z740D4MZv
QJjQ2DgY6HAXgk6BXZqWNpPGQMNZET7kSxvUdm7IyBTMLs3DoGiwxGLcHNwtOI9N1tVcNJ0mKlPW
6ASg5HVHZLRYEIDX5DXG42vVG2KOEPNn+L0x+hK6yAh+UJVJr4LXmR3+PUa9SiDs0bAbJENK+t5A
XKzI85o8Pb8vDAchok2IYlryrJ/ikaZX+oxEam9gx8cWCxB4fSC8RnGb5XV3OBvcHW9KmORlmqCe
jxZAibjRT879P9Xcb7iwFEgSKEKvZcOr42HhnD+INmv3ZC75+n6F2hz+tKM1FM0GNsA4M7+6lKCA
1fLxOB/TL0qg2umjC4sic7/GM/sAIjmwGP55P6BsRF/vXtB+MJVkECYRXO+rGyVtsRKlx96y55qd
fZyXSDT4ZNp/DyJp8UNaEIMQ00/ywkx7Zm93Kq/o5opsvbBd360E0nybNdUzREdBHJjUAK7y0YEn
ehvU92ANqHEimH521H2iL7IQwua3IPlcKNIMtd4Wr1Fvcl7A+N8+3GkEdmfJO8IC2/Y4bYZpek9Q
WRzFkRK2vFkVR4Ir3hwGk06IbDHddSO0mInQqpn6OYyGoXSFeuEYNXkyTFodtn6V2PYdSN5eoG69
IGukQc5rroaqcqiR1tVpu6rUdM5zDba/GiF+7asUrqIolBoo54bQUuP77+687as7j6Sznbahyp0w
Ona1EKxlvyDbn4T+DCvYz5vxmrHHYas/bgqZ6D8ZVRRke/+i/bd0wppZ0U8U9a0EvI+FwrgzdMht
SEyEEu8Iu7sNbSfZWAZ0o1p7tWkPUZSKTqIAKa2T5XJsEMfZUE82zovAxVj7Vyc4yBVPDZmikOO0
uCoEM3JCiBj457zXWBTxIjBXFjq38UfA2bLfy5ut0sZIKj9NtqWQtKjsFKXHLdj0d21IBObl8hew
egYirq8tOx0DN13DmPou7AAimZBcRoSpDw3O9Bq6utTjPWHmLOGvpVcULyoTEelT/0BD3+T3x+Te
TzWjGwKQYURekqRnSQAg1paE1z3Vj8P0a34QOEEh+biRljlD3E3L1AcD7J36nj6Pbqo+P9g1ZVR+
a8fPSZc8EKrU/yEwHao9Wk8OQx96HxbRfa0qwne/ZXmuVSmZUryMjBHJXv2cOsY2M0wR+LHPzYYC
vw5Ve3c9RmNLt/kaudIKTStvW/vJ5vH+4ZgeNu7y6fH99mwjamm/lPD9PcYM++6JqymhEy52rRmk
RvRxHKnKXqawPdBJcmMo9xcAem2RaBNuX2xSiSjSSXcA4rmmQB4OvnTpSOSg3KAUBIzAJqc5+k9B
q+NZA9/dofX6J5XSTs7C2s6Sowk1HbbS7r9QXCkO/EszGAQtsoDZN8e0qK89yxUC5I3Rg6MXV/Xp
qFNWYDsTWgYfDTW7dWj47fCUhXgP166lI6h88aftOEAtfYUJu9paKoJAa3IjpBKwOUlztLYH9FSW
UxrobWpN8fzI2Q62RQUNzEMkXnmQbKR0LOOTtzHPrIr/VunJg1BrNPAIfw0Pg7U+ztQYn/x/QP9W
e5xJK3SYk8UW7PWKiwjnfmHWoMpvui2iJ60nsgPfcoN/0w7KAxCtStunAuZlaSkOudF9GycgUwvN
xF4QsNeEL+/CVakTBvUiOuBZMpLbaw0XJ5glBPjqVOhbp0kY1g9LYJsTVGcYamt2cKgXlGvkM0Tx
mpxRxTjkxht/M+Ysi7h80hZy5tsQhb7E6HszahL7ntnjTptWnnllWiuYjCdCTJU4wclETFBtWARP
9TF69IZpuoyRz5tmPkpinpwPO4WVTxIKemNpqfa8I/M+gmVJItVH+LJfyN3bXVkaT333WuN9/xDB
smJj7aHJ+cETt0siYZF/bLq4VJ1R+ipSQRyV3fkYyZpX/10BmiwrtqmDsC5kEVQHznicxqtT52eB
6YzhydwLNndQrTLq32KBlhX+Uv66rVxw7P51CT8gxWXK+x4ZOCY+Rr6qEmoAt+H+mrxn58yfvMSr
I1BNhjFq2DiHfGlD00RjvFVeKgvi86Ws/AwjwiMdF3rI8s6V5SXpnZCQ2AlHVCPPDGNagR+YTnHs
sDs1xBuEzQREZv3YnAYwfIobDwqWVnNhutiJL3e24D5uV2lJ5gWo1EqyKHCdl5E6zRjcIe1dLkZ+
qFP9vHPYhZYt+hXD3bsYsDHEBO3DULFbwdAFGPGdONtaBtq/bBE5MYWUsFX2V0mVO05Ay3xsEG6h
hFb8SWV4hy0YPkNyyxkpzsSTFXW9zh6gzS4SJnnis4k/nq85UHrDwfJ6Etqn4I2ByrAHgtLpVuFR
Rob+DLc0fe7NZ/eAXUu7ezmnq5AEPChu4Uo2h1luiZ7ZfV9N7R9EmL1RWjpUeWnm84MBXY7i9Ap6
xeArPIk8syQc/BH0abLs//4tuGEkBaSNnRgx0iwtmZInbck0KhHkuoFeVxoaeATjnGcEYiRaSeIK
FrxTAI8F+nVg0Nm08H/3/rnyNW6qkCFnLTxXHankTXmbN+tVQTPEXuLPtoK3ytoZ8Pw7Cwh5VhQt
o3yYBAxDsfsXZjDpzhfpPiqjgFbguOHBG640esdRtg7bAuE4SYyWoK0bd5kXJUrZtCkwzUyb5tTx
6gs6RJOk3mCqYXBhV0DdvBOpNR3+MiTyDXpch1CUTFS8rgHGqROM89JKJTDNKQQHrma6ksHmwZX6
RpIzfBzZk3S22uDjV6yz3sqfvM+/iUWPtWXujRDRr9MhKAPq2L4WaeBdtuqEJS4M+8bWuV4T7vnr
LqS/dAJXQVp265AY42MYUz8qLMNLy42JX2i27dhmTB8VLQ8u/OROjWFPziThqZzhsfWkJ7eKfOca
bHs37vXFFWKmlbZsh/mvk4aiRNGZxhuzQ3AEfMmo/C+UxYCWCQmuSgM4tbwH7IKAj5pFqDOV1azu
6FZPXn0JZYcGDsVnB5rJHzkFmGJu/OvUBDJvAPqRmG2CPgW+ERH6yQM117mZ7NVjdrw9oOJBKA4Q
CbyexJSKpTGRquz8kejhkhV6VuCeQsXi0CEJ+1Qh5htM5ccbyu3ZFSneS+o1XRXrxIJpeRuEMCnl
o39+er1aJW3xFm44Fk2CjQym3PqiouYNokIfHWeCrH10WMGFkFVC//EX87dccwPozdfgofUbcm6R
snGOiPf1OMD0IYju5KIq2/86vJLmqFjU1szso5yrH6j7pQnhYMwMOMyTJARRv4Z/eGQsWI4fn/L6
MO0sDpzl1Ffqg4lgQuPN2ugT8lsXrx2NSjqbIjNJJ1aZ8f6VZFZoSznOe9SyHfNVEAXnfh58Xesf
qCPKKPxCswJrkhUVM9NMwdVeyMhm1tLp0r+SrN1cNqEyIczWrS73L3fV4HqkiXqvBdfkD/G55vo3
oEyrJOhzmDbQFT1gYRzdycPUyKRv11iJGs/zUEtStfbmvaOVv6Xc8QerTtjr1pJOsRaISSYhCl1A
9dsx3Xbxf01tkHJJTvRcfGTKQph9u4/pK4Txp60FX4oE+zu7ONWK4Mxzyc5+fH6wAsb5Mhote8wr
uMjR3J+EwdsLI6eXGV661/v7DmW4/7UgeQaPapB0o/+gPY+nPQk+Kh59WcfauA/ef79+bnMxsnNh
1VDEATGKMQ5ftQtxjPkOaHDJtNu7ME5Px/TubXbcHNOIGkb/TZYz5SIMlp9B3XKqxNmNiKmw3lip
ywrzfUqPLFIWFlkEIXxtY/MiuNOj/Mf19wUAPI+luBrylRwXvCC4n9iUUGluSvKnZGgtnDjbxObL
Tf/igHZWQCQ+xr50Jl86YHgCPj1ocDXmyzQCrgpil7JMXi/EYchx/SBcNpyDwtj3P8xYUwRUvBzI
oM+FOgS1AAXhQXiKCgp94vRVp2DmyGv+hTt9oWtFmtn54MOroGt3RIXLLVTq37C26VgRvatWyqcV
GKb4KypcJpGEVrdgEg/VvF8tj55e4yYCoUL0FH8A0lEV5J0HknXoNeBxikfSFO9mY87SOBZTcE9l
Borb3JvzLJ0W+Fe3mN+ZnI52t4G4gb5lE1PTe0X40t9R8CpRhmM6/LJ5d1gElselbzdGL42J+9F6
4d3/E2QcNFXCoUv7hEXhKQoza7UZQnCjBO0fUFNUhFy8lLasVVoWSP85jhdDqO4BWNuQfEUAQJvb
5NsEN+X6U94na51COqnpoqUpgMPEF5q1Pn2y9ClVq4KNbUFFxZT17+ea4EIx8QOHAJVVmIemGt+F
86cy2kb5w6G57TRr0P9Eowvfq7ONTnnLN6i3VCcrWxJjbTuDNtTxaLyo6ruTwiQ+oTvJ0dEGEHV8
JM9r/MBKjKwDyfXBZb7nMVscNeL3lohMFsPlwE/Ec2JsfBGE+9xDntWTQbXNbsVA6aH0rN8skjFG
fTOM/SMWyxj0V2C0/PJCGouhSIUB80B3RCAUvsCCL05HqjszDHEs26/xwvudwlhV0mLqj87kSkrk
KXczPW8drV1VoqcEscAtwe24IxoMssFxR+7GstdougoyHgCDcAlhPjRWqewyMmvimYvGe0MkGiFS
XUsBeFMdczPHD9UFHvtcGkVzuWuEzPfYUEZFCNSHjPAM7xd3XdIikPkKNIcE1saqL2oFTyzE4sdb
NSu3ZBZEpudza6MMwUBXqE7Y7v81fYBPlJ8I3bOhADqxhmJAJvVcS9y4hm8LPj3Vjhw7V133rQVK
zVMo+sC47UXIhbjbHeaMYVwcEW01HU9DzWWxwusGCRaypmZg2uUnzYj1lY2gGSyffH0EJiIQEcGl
uGeEjWOg5mEPLRv6mCBcy5vDoWBpzX+JGsI5YB6toQODm/NoHLcGukpndziL3DKqp8Uqck7nBSo1
ZWR71zTSkRtXSw4oAx6EW/WkFFPkU5I9zHAe3vG63462cloY3Jd1ZCsuCUOcrQq08aDzcI9j8mes
nVjraabjlCcVZSA7I6j99QB5jUsz+8dacpDA0vfMHpGE3/c6saxIG5xhTILMfehjOXN7LwWZy3zB
iVjvoYGQZXA3fvhb0vnT89Tj/8xFn7m14/7yhqpbhnWhbK94HaiShrzDM3wE8Xw5o86JGFx23+y9
EQes0bXWeEzmMuJGdytRW0XaF1020evK9GMhXJVelI85O4Ac6S3yCKO6py7ngTiZCyK5802bugkV
1Yof6yAkzftIDaonQ3nIaR6bJ+jko7LOEtXwu7MAxFpr+P4Z4YtR5zKWFfv5fMom2OBuvyproYYY
3VVMNeyYk/ruWDTN0/g6y4CGlmUac8l/61IIqd3BpChkAtqiJGN7qoj/O+VpCvoBTw4w/DYD3Kn9
DjdC+vWTqsWEEyylhlPF2lI5flN8NM2DLesroCZ4rDX4FfpCWgyn1KBKLOOki4LbbMXX7ibpgtBD
VtdfHg3LlVhFHjio+KfRF7vvs3YVeQxsRySAX+KzimdNmui0oNp8I5PJ9M3QlEP/vksCnt3kN97c
FZRGrcMgUEQ8EqLh2a7f6IJ6GFEMqOn5lpDWUx1XlxcCsvML71HttgBeGDZwQ9F+HwfYnQeZbM7Q
vJgaRSh9r2qah8rHY+THuDTFfyNpuKlQVh5kRXLBKKqwZtrI0INalkZ7EYY70pRgzBOeH1jsM8zQ
7xSklZqSPqDqPyW+SF2jUtY9f1RXyPBszln30oBvIXrnr0BCGm1plvElydpzmgt72EL5P60wabb3
cDuOUVf8jE3Dr9PxfiO1PXn6ejA7uZXMJp1Xrp4ssJQZ+Rm7JSjHRP0elQwvKgZKbtGEqSd+fMIM
0D92c45kepO/yc2RDmXZW7gw1YSz84EJZZbk+b9aS23Pjfqfy9i0kBygPyO8y8bsYNNCIwSSanQh
6A0anFSHlRCiXKt1XtvBuPKqUFYrEYuAGRT0PAuXSn95yP62Y/2zmKQz9A/2pepwp7jj9SGlw8bO
MDYIdGixBXxviArUys81fAgi9u6SEXnyVAGrw0bOXxuQPeunzXeUvtWqHJy1m/qCp+idWkCh36vf
D02cuD9IiWGi2UHTrqKrdpAmMomQXmC8Vt8+GUL0hU4gN/hnp4lNPKox8zkajjMY+6RcDVYoXVBO
W3j94x4Vd3qlteJSnRkMmabQYNmBU5ybCeBUCeMzi2bRQ+ySMCisxTT2YckgOzUFSZwCTzZPLqvv
VvowOa1ihjZbK5ho0yEetc0+JEA3OrhhJtRkp+VOF4V6ObFmL8lLdcaLN9RbZVKPAw0/MOj3JdPV
VJM8eM/F++9sIDqrsJwE8+Dvt0CCGpSsgR3uOsmOqmIXNxanPZbLCnCAYij2NlOR8CYpuq7Kcog3
7ef6jbx4qKvO/yqiw5p5Z+7eOm/AS16HcNDikjszzn3kiWp4TA5lclFuFYd/HhTiT/GnY72+Vlt2
II6FdS/8ogV/Uc7vK6nzBmxzA5VC6jgbGzrLpCA0zb2f1IYHucViM4J/QnSPDVV4Ms2PDsChP5AD
EXAl2JmA21xfVuBV046h0hzO7AowEntLXg97Gahh6LB8Fxf3RtPIezmI+9r3ci+sYrn4o9eybqHS
ENTQCiXbN5nQsYTkqX7BMlhwKNbP+aO32LPIUOFFfodJHoYn1rN1oe+8HkgZSMX/vT0bf1n2ITWi
faeWrDQVe+c4ArK2jWfXbwVCu5CbqBQjCEsbQcZFXQIb2MkEnU1E//o1/wRxzPmIJnf55T6QPgTE
o6lkfvmARu8pm+1AXxA8x6H67aYRYyELfq8tCxEL75DycNAH4otZT/gNTRrExQ3tX7AGRcNKWOuW
9ZZ6xbgfH0CMPBLGIwEmwVk6L030oogYNDn23R/0U9dHWq30aNdvzWsp0WRM/OswCBl1sPHFgdFr
y5A03vARdwzf9yCZledUqiHE6P6ybP9a+LEwuX0OLv6ms6Lf+fx7BWW23rqNFF+FtyrpGab+spQB
utmIyAC8ZJ53DdIzAsJaIKYWXSAXRrv471dWNR2C/ryz9lCt0xS+fyxTlCseWJPUbHVkfAaZHejl
XbeWBmFG7Psyr0i9fQuEPJneHwb8fEn9ACSDdJh2oI3q//r3RyRLJw1qACpt0jR31phsa+qe4kB9
seBJ8Nmy7oUeAeGd901FjQ0xqbcClJdi5y4VivBitVVso5B8lQ+hzF697g7ZlXaQSEy21WcLNDuO
4LTdc3wZVgPGKVBVYSp67yPYl2SO+zaaI7BsbkQYcB9MK3a5AFzrNjmv5FcD2B0tU+4tAVW8LMZW
p0ahhGUaTDEDf8ui/Maf4pNkImUQ3a+3NpbdCM31bdUF04OFZvxahnOaqFFDl26GJxDLcOi1B5gB
MOIaVO3SoTTKjw/68bS1pEWAm+YFD6C9EEbxiHkU+dPYm/2ePTRIifGDQK+iZOUfV9lC0ysaEP37
uTXk6PLwL1d6mBxPdj0BaDWDocqFt4qqJm++7WViGHL66N6eZsNwtlk0s0RrC0aWOQY2lGd/Ctp8
1fziBWZVTw52F/3IMh61ao3ajoTGv7xfvd0hUu4F0wR5tZyACAkk7brSSUj91lidRNoPyL1lepND
zSL12n/QUPenmmbo+qgENki47Zp3o/Lm03mF1OjD6VdDZgRX6FJA3ozE0LYAj8+Cxsa4aFu7SLOe
5ylsHpeV9pjyy5z47A3CK+UW1Z0M7zxxH3+f+B4cHLIPygN/2VPXqUlFqJyas3gwD029xO21W9Q8
DSXw6r9B8sygb8DMoYihTi734FKyIimHkX4vIvXBaMtuYCKJFsYVxv/pJZIjwMYjTwB0qn+2PwW4
CkvkUjYGizmL6rX5quXe8X05ksR1eQCzUUPb8hzMZgSacNUqlb6EjIhz1NP86VhUxk49luQ+b0Zx
zHYvThcE//zE64Jtf3eAnJVKxC4BXy836qX4JH2puhCVL2fo+QHelgzuB6gQDsMvFUsfHONnDXpT
hKtNzu/u6fhAjNwFnp/Qm9jDq/fDpxbpppmdbM5KlTj3ruVOq5eTq8NbqkJ7Ik4qm6kwplaKm5N8
69gtEKqPJambLkp/lXLxKyd0qVdksRWQZUfYtdi93VuLHNHMqa0GAIBoQL61gYWnlj4gHErMAQMt
ShUXillEarlZk1VLPp3XENNfQeSMVPzhKAgFbhjdA4R+sxQ/s4xkXDYU36+Suq6Y8Q7cRoWmPL3x
Z4Wssm1iW9+mNz1tBNOeX44xoLqJE40FAEhU+YReeyu3SXyDHoQu1Elvh7pWVrwsHamncEVjqhgp
Ib5YjMkXCY6OfHJHLL5eEmHQCBnUV0rCGtZ+UQpvQV2UZhnZIVa2IcuektWXNucpdJb142q2cFLL
caeik9j51k445SGfgkaMQDHR1PjO2PRKcOWI9G241o+0U2HfDJo0tExs032pXo3pVxGcBpMc9AU+
MohVfMjUJ1WYRLExFfWMfPkML7bzTjXRtSPmC/HCsj5YDmaTeort08ZO3es4VXyJr2ts4Av+ny1g
yQ809Ea4LaRCBggp/a//cxJyNjD5EsDmDgwUcukltrLvNLiMoW8Tbibssq0S7TSaN1A7mogxOIaj
agcB/wPlKrqI30sQ3ykDl8EpNG5JP8HfRZ5h5/ciaGsZganJpL88Y6uDW2tK6zr81m0YbkqYAB8Z
fGZKhDRMLScWrekJ+QWc+Q+9EvohmetIj2beDv6VbQr8+YxUgl9JMdFsOyt+5d1HG89hYd6+vDcT
yrh1N7LN0tCVoqmZvEbsREiDU9U/X6jk1Y02U0YExI3svkzsexfQ/4w1G66RRSl4Gyw7NrulDZPQ
PB+9f5B2g2hq8PbBvtdCyqeDjbwDDm92hk4l0+J1O70IIZatnQCJmGIymXh8jMuGdkbAsKaf+Q9K
Re84oBJWVXxeoLJiC0kzxiv6i95paLO1uPLg3X0319YfoDbWbjcDoj25pIXRwAbk+0uH8tV9qT1G
KkGGLZUtm/OBQboKs4o3fcaBqY+jkMTdXCIYNqosaf3yMC43dv7PlWtowemVTurpzsiGMOOpoJgn
Sbuxx1xNYBanAfNwK5339rhPv4oKBoHfZZGLwVxu9IejID+SmqS6IeNwYl1n8mPUzSGzkLqDzcDE
D9vq49JIzO8rY0gv+qygu8tHFVRLUEvl/h8IyqlzugjSR44YPK6pcSTIgo/fQ92LFR3u+2+XKNwd
4MAKH8JpXLnG8ZJaLTpe5pyZKXJAdT+xeoH5ywklMZPhq6xvLoJ/Za+lhJsryjhDRsFGvmIk4k32
lrDs8Io2z5E5jwRQBvrTbIf69RU6KXM/Oyk5d06XDZ24/1k40i9Lg6ec7xbw8Ocx6kl8yXo9Apqn
hOTbQNuxkoD0Mb1n8xadaiBEnsew3EE/KdC9UkYtInjRnQ4Hop1+EIXWP4Uj5RLaA0aU/CCPFo5j
Btwq4/4OcCg8fp3mUj+OTtVwmSXqzLQcUq+h2aE20qWdY5OK8QYjvdUzrGL70ktdJuAKwEjocVfO
cTD+do2tIMxB359rqKp7REkN40Gucv2+IPnEKeM6VRCZU4sGs5V73cVSB+OCpursTb4PiEDHLfGR
Jftx6XV+iGH/JMGib0Mvu9opJ9dgLxx9TQi7RxL80dHjYpyzGtyZ5dbwnMJwvSyJCE9xhZsTN2Uw
vo27/NIeaxyqKcVHCTWgj03grAt8BxGywAYXNR0ZoA6iMLdyoCLQi8VwlOz75EQUvIKd6yXHn/Sd
jDuRlVCRGSxWXzlyKtJiiJENvx/k8JVDMs4oQCVOJHBJ7N9LvWo4PlrAc4FwcRsHvvlbXFwPHTkr
1vzjkNJ62Hy4knW4DxouQSrspTwPyGgrhEjG+DQKedfVcpLuTiJMqxh0SL3Qg6eV9LauDc5XgVSG
AzZ4vAV8OiROc8Wv/TinnB6KyltR0dOb88puGrVyAyzT80a2r/UQ5t5lLtFuF+YnsjEV0BspFfGh
WGQWRZm5evl5tmRqhvmRfj3affdnqv6mWSPjjCebhnwKqgJyqJf+CiVc2jgfqcv+e1stZiQ/z1GO
zL0/oe7pdiIRiGJHhDOyCqkG8S4FFo9gJqEOSCZ0qsDL9doUSstj7XRRKpzvJvSNXqWoByzcaSWe
/6KLxAxbcAcnQxaOQz1CU6xKZJOZiNvi/GcSGALEVxvsWTSzzm6ukDvoTJx0mJFRRMAkg+hvX6fT
luc+VbAFH7Zv6H+w5FjfJC7hw8xCzDl9jJ4jBfaTFagzNVZsZfTBe+4Ub0RHzzFTndLT/Ysa2SWU
hgraTJNdTDcgrb9ToE6YkJTLw3W2rZSQ3d8hcuEmHVW3EvGjIL8PRbgECWDSq9jKkHNlY3qmh+GA
Wn/Y5XBMDMleLMnD50Uxo6xVmG6rtWJgqIddheOZIQpyh7tGnChvKsDAKHlp9nICeoivwfUqS5zP
KG89RLdU64io/z0s9MhskliNTo5q2unQDTOao+TyBIbBlRx8/Qcqm9yg7nRH3yyg8RgBTHhtqhKR
QNikpZpuIMWk+1Y2C05EHPs90BwZHPEAU/gncuTZgFl6B6mrPn/q8ScbBbiuMGZ1ccd02EWzOtKt
2p+6uZTnAB/48Kg7SKIfGisx4ZJR2OWcHti5kmNqBtnH1pPRhbCehsCshYoIaSLupyzm270hQUGH
DIJ0qgh6kM5oRO36Vf2fEFthqPaKO0C/MLUWShEISO5zqol4sg4K7LAR1nn0Kd9mTeD9eJG6uALQ
dqL//EgyCHCdPfSLhudit5etBcxChoHatxk+A7l8l4HTxZYPFhaHrWfnuA9woS7iB2AlNAxhf6JC
j6t2iArZc/zxzj1b+aewLLhc+Xij+WSRLrnd8FAQPcPIZYcP+ID2FuF3Y5pS9a/eBYTYSkec8dAX
XN04Gc2QmFehr7hBXHmsE/PtDccEqd33e4SDT1xvqd9eFbOctkcbm+sYOWkyGULXFtwlSV/LFk0x
oSNCETTmJ9C+tlDVNYlWth3e1I9FGKplL1ruqsM3su+ArM9ahfudrsN6WFeZ510Is0RdDOuqlkAn
/h03YG95p1tHE2zuhhl2/Ko7ylO588deSJP7RqI7TS2k1El/KRkWHM5UuaWWqFPTGyzHOYc0vczR
xyjhfUwCbRVPj0mv8XiT2XThv9RNGWNS8Mwv2+gMZ+hVIwAVI/un88mUp+21WjSpcIi2LDDVf1HN
H6tD51ysm8d1QTz1Yo3ItfjM/9DKj4OCtuKMbfu4v9E+Mz0YkqCP6HTXjLrvzzMiFdBMqohuFaY/
RsLtSXck81ALqmFKWzWFZiZcbLROkBAUo5jUJQa9K/XIUweIynHgpbAilcvsR4qEeOS+SKboPwOy
sc5yB5FuoHrjWXYeEMMOllpJ826rxNxpz4RSKM2SGRBoNgjJWDJJ3Tij69TpZAT9g754GE0j8QOk
ON4yEziIy9zu6ceN6uExi/G7l1nlyWC/YhRCyNFQIj094ldEcXsgUdATdcOQKYySMmM8mtLVIFbD
xq+HjbfAgA77TMu3ZpPcC0afqkdZIP+TGsMrpo+uBb7PQGpjSs/dFJL6UkWBP1mZTQMBClxsIoId
FXb5GW98BRdWPwJpwhVfMyNWdicoorov/cn75YT73gykjI8yh6hpVSho7TiWz5+ixITXs16DIZCM
kb2HumK4B8l9ChC7XBNPhc0yY+g2i4ASA6hYZIZ7lxqRqqR3WMp17V8egfrA4Obk87wgHMApBbrp
z6DwlAIYQgzmmbO6MqiFRx+uUZtwgxXvxheZt58oipmqVXLDKQJZWZKFmzxgcVr6vlaVZAEMR1jj
Ry5CIiPsaE/SWJ5cMMumUoC8Wqwp875yALoGDl2UTmeytRUts0kccs3TYpO5aEa1FxY9GEWNlbIt
imGyS39w9nhj6fPA6Ky6QNt1gEPvAMD7epxjxlMFJhtyN8M5G0i0pvr1hWoKg/NBDwgB3yCr5Z3x
BDYDWIwslOSG+atS9R3c3OY/arAw1hz2rXe0oAwsxwiP10espUlKOilqjegTBQFIFDMCysntstEe
azVRsMc7J3WH4lwle4N+XWNqTQBKGiMKJCBv9S7RQZuLnhVHF3PEJjwS/MfDdB4sZYM9cAjStmJ4
Gw5+Nv8Xc61DuyWxzZ+1ylzY/rFSyXyNJ9dLOJVi1xZqJKckCiSAzzKqKN647xDpHFrPCOYH2Wib
hiy98ECw3UNoncfNBZ7ztXbECDRBOiU8wbQxOnbcpt8DBA+JpS/Sbo80E4juJn3wICstxy1yBghk
pq7BThOowSXpbvqgmbyLykYuh7x/CP+3AqffXqmHjlfhYolIrl3c4KYwOv3uYjeBb8MuZbC/eXqm
/PBsUp4ehDXuj1xQKXO7sbB/v4XOnRSLhO4y2CKKPb+M1zMHN3YnOJ9M72i6DrrndIL2M3uRi0jX
OodMQQsqXiD4wtPHyAILKkgLYhOV3ZEQda8sdCvxlguPWJ1V9epCvLlW/MX9O0kdXpUR2SeQvjsJ
g20c1+5L047p1n/oWg2d7xCmqNcreJMB4wwmChPfhHI0MhOLs6DHoKBvw/Wc1r2Ta1/QwJ1OQ9jv
ROFawVfmMj6n5KnZpquR1WtCGTMP5LpZUNid0Uh3M/DBxRiToK02K6OdAm3XeJemxBSrsmbOedfs
UJK9vu/h3fq13fgQaIoDNe7k1dfqaFk50G8LU/d6lqDa785340Gt1AhLIg+FXSgC9di+x2JW1msQ
/yA74l22ZmtK1lNWdkT1akSqp7lyBiqMGkncrt42SiKEnksKbSJo9A6KAEchFB4D6lH+mI4PBhcf
4qwRKiTLMmxXLjHbkSS6kii+qyHtT8dxkLDlphqBT68Vb1y1p/U7lZk6l4y8oS6gWNTZMIhb/SED
7UAbG9BraSYhnipc6MR5P1gKPoRIy/5btmGoB/SvR3apwN+2yX4yw8OFGJe8f6JirxlKWBvXT2db
KA3bmd+V6phxRmjcntacIuLN9p+JZ4e4E2vVj+WSm1TlAsQUgMRRUMkjf4oW8EXmzaZaoyM0o7Fy
4FaSQznt9pgi0Qc3SBB3qBMWK3tT8ZBSSaJ1N0yk166r2EmGneT9kIVn09Vr5g5+4via8aO7q65H
LSHiKs/coz64BJTOx1z5T+L+qv5Jh3hkWcudzZfGOBDWCKYdKGGDp+q/2QU8ytFv1nMTJC1Z4smq
I4GvKvYo0jJXNUjX0zBSPwVxuVGFnPJE9eC6SgOTHv0fiWGIr/S4mGM48PL3r1UAcBGhTQYq1nco
mVU24Nf9ctdng+90juAXF8Q9FZK2o0cCmxgyesMExyJo7O6pHTkpThkYQHZlngHf40cEKoWS2OTI
MJe1i+gWXwhtz/bbAgpfoRfBpd2yQn++VFVB6/zIbzGYXbMNOhLVhe8FqJibYgb98ZOJJn52E9w4
AECo8CvsY4UqXAdZEAETObG6dkNtJ6bjRhKuwCdwZby3K3s1djiPa2s+cf3++1VITh/9v76GgAM8
UV/nl1//gLDuLiLTHEmLhk712FxgxAJLzirlFumro5cvwX9pXhPndYgMzA/bLG9yebi1+HqTcZSj
J80MLVRfMkuPXXic84bE/uFrsRLh9xs2HblZ6g0PxCwAqCMCrHIiW0+VBIlpYq6Q9ybpP4KuqVqt
FmNn+/cgSV2EdP9yLYaf06pHDE/Zo62hNtSZA2FTbnysWLIt4ckOblOFhXxAtArfQJxoHL+g9kuu
5yHtwsXxNnzL6KBIUFLNGqyqOmACz3j/r9FIUuM+lH6Q6YP4SuXkEqOwLxZtvHALPClcBWjr18C0
C1EIiQwTILDPxVteTq3f/Cu8nRgLQQA3vXgOd2FFO1qEiWvlQUtgnAtFzjS9wSMakHm3xmknPnxu
5ZRk1CauuUDqOhsGKV8Bqa3//OZS2M9xCZRwkMITR9AFUZP+0Cq7FFMSLra3JtaZIBFbTCyxRGj+
0iqRfY8opwn329h/Svnalju61zEWK68kQF5imHSbsVv1/9gcpSY7ZFmeen+po0fuShXY4VPmqkEz
iTSQoXmjgaqjhXIQJwULpGoluhhUAyKRXBjmanjk/53vjH9TmPiyd7Vs6YKSSM+WXul/03gUn2Uc
50xkD/01WgyfPpcIzeYU62yEpdRZWaz+CRMG0QJtfGoKhkeyDG1w92XM+5Ph3Wod5YNwaGycBJLi
nAv9RisHvlyG4sbAp9U+WEEKtNRRKaVWI0xwJ98jOg089W8luGpIFxyZjfbOw/5cNQH5V+hb8qnR
IlXXW6qMgvnd4tHWVTQS37BpJerGv6alBnyqHZsvdAN0OmiRdzq3c29NTzmmY7J9Otss7zuChktu
2FQlJdEAsv1YGhc1ZB3hBIW1vU/BXBJ3xbyVVPDizng4EbpOVIfj3w3KRsQYDtxw90W4ay4RAgF1
I9ak9xTRboxg8oNdu5VxLJO5/6nqgyzrSntFTQUG55Y+M6X2NBNL4EfPO1hn54f/QxVXUMYlFVhq
xx7+2D5rGVXCchvtTuKWcWiswWIx9rTj3ED6qb015M/MkLOvloaKcWXZFky0lh7pywWa2IcKAFYo
V3tmiCBnGubChQkteKHIpD9bg0lImJCS3utLF+XPiCxfEWzCoUS6JjTlF82Rh5mUTCX6ieRc+hiw
cYE5Qt8Q163eKv4chMe8jIZW9np51h3nS67aqxLpjTMANU9kVFOvbplxlkiZ0gIgCgEXvDh3sMiQ
8wICzh+J5lMFfGWqEWH1JfYacDX7EvzCN5nQCaSYZvnvdLLvXC94yd5cHymQ1OmfVH6gZW8Cy2A2
gVin2dj/4nkTdT011sU7IwnliKyy4RhidoPrJOb25zaW712Fl4hDnY/boFjN6LvwtqL0jDNqyEyC
zFJerYUTzDfju7D+OAXwHiQl5Fb1DIZM3lBJun1OO6iZMrxN+DazaLRWUOVkdq+i9eneWJFEDRl4
2MRwrZ/1PD3FKxhgLo/yKnqL6BIXBhgiztIz2VPI/GUYZh5+SXCBcgfWiVoN5S398/dhv+ghWg7w
P4WzJmPbbwPE7nY57hh577uto0K4y0DUbP3RYXbkgXO39Gwxg7AYN5cBujG4GIaPNwtKjXbQygyJ
donY3G15/xYOVeYhp2G9tYhp0FnOGUBP+LKCD8u9Adm8PTig8asXe/jMCVrtURncpJJ3E1Wc3w5h
M4XCthscP+EMay8I6lWeXnnFAA/OpuTXR/RGzsjbSGkCq/gWbDbhVCwvy/5ycS5+56oMjsmwtZvT
38HGvyA7/gh4RbSqBNssVUtVx9vV4syrQoSgQh1uZyMZKRcof5ua8n6mJpdUKkpo2oFCaPmPly/O
buihAhw8/kS8ILJTno5Kwb+VX2go6H2IqufOgYTlm7HyILTlNeyU3Szu2/eoY3+kmRzZNXrSRR/r
qz/2pTvbHXxxoTiZ46w291NS5NCruyDK3OHp/h3OWFX65ro2TfLmOjpWmEi2w2YKQhxfSfPHoT2W
uvuFGhRIb1OSfqK1p2czgijwIZhJjqmzx9qWeL97cpTv5TbdnYYQkWU5xmTiq1GycuWbN7s4EJ6F
g0fqbjKNV3rmS0HEWYYhE4h0nSfMzEfqeh7Mtzy3imGuhyUIpdhaSxumBOXrgzL+A0RVtgJ9ukv+
XoPsQWQIYS+TulWEJXXcwll5T57OWSDsfBvs7gMYrNZauCHh2NW7VTLWNSSFhCBNinggBEkFm4qV
RfC2GvF2lmSa+oOqiLMHiTOwQ5RiShmnLQ23R8vWqm9Z6nV89SwjSThPPbAkAU90ggOJ7m8hPvIg
yclpvpl2KfJdDkHliLKRTfcBJln71T8NSlGF/nU9wNnyKyl/2cJ5gJBlqbimcGwVO+QteYM/Rwp0
M9ogcV0gB4G+qW/ArEYcNofIDcC+5zGcgysyl9cchODQVpiLsVWbI8UzCzhDgEJinSEbmErXa7Gk
y7DkGoWsvG0E6OMueWxfgQT/TpGvZRoMPgd8HXT4KC5Lt/h/u5I36FSzo9wB4O3UMsvHp794Tuqb
TuBeUAlPqhW4j1hs71iru4idE+DxLmDI02cu3qRXMGa5w2b9TwHY6QFQQvmEFg/ttkS9bgrzkx6w
Vo2TEPtV0FG+pctyLeXE+bkcOnPVlfgEFERdklKLPQ4Gu/yZN9QfHUJCh+DA6Uap8mao5w0NqGDa
jhy07eYkTvNoLWB4PJAgAK2Pub6ULpf4B+idQWvnt/AhgIPhfrxZXX7EzJCgAMM6+C3zmexs40YE
tk1w5batNtCHRNaEq7s4ADzQ12pS0Qy3lMAwU8lnPff5R6vPbKj5i8toJBlLxXzpIJzp3SBcQOjF
Xnjj1jDZVatSolLdnpeoQ3E1xP+9/KtVvPkohz5EJNJJ8Pbmijfs+KYsB+AgZJjypc7uZF5jmQ2u
dciKey9tq7UIw7YrCWManswgP1nHVxyyjYliwb8WNe0uE+7mz4KdqdWpltmeECyVAHpkF6SiZ9iK
3kU8/Vqb2WPvKRDDeosPuUcR0l+zBFSXBQNb1dxvf3PgfDOLOoyGRZCkkjeR65b21CX0sCVQGEIi
q8utkzI3DLzYBrEvQ3JmGTkiuXPT7lI24ZILy8Xy7prZThDVptY/ndUzb0jBJR/dcZYuAyOqLuI3
XZJ+6vJbDy0g6mi2J2nUEYpwHmWSfNZXYwEX/BSfoolU668pjtou9SbkPgKaLzkb4RKELYgmH0lW
iSade9Wm6YokTxdJ/nD2M6ewndxPmrbg9ngYT1xUjAW1c/FDfLGLQKa98AXtGb3uLh4Nmh9hy+tc
WCVi87UANPcNCm1wzM2QSky2zr+3cH1zizHQQ6rqDYj0dTGaMe/TOcpMASCuU0mI6rCNCSU1RONz
vUajxsSfOT6Sh48G5oLp5Hj/17kYj1QouEH5V9ha+OPjpSJAWwTYrzsdAxQbMnUm8PdEoPyBWawW
MFKh83mAGpp0qsdStPwcksBL70vUDQDskRU5iSNZ66smFQTzYeI30kRZfUb/sb3xI0laHdRzBkTS
thvnW6X2t1O0XY1/HcYgBEvee9cz2kmr6BDvV5+6a1fW+n0kL9HbjAOMBexP1LslhlasNGg1Jsyl
huQNNU0E4BoN+NwY1bnmQYrDXBXP9ie98J4YOjUld8GS4G41w2HMNvqAYkpg6coLzXnIHjC5HYcv
wvQ4obX6EyfFFAMeulzjrmRhyUPpW4c/AriNfkEHXzun57eBcJkwvZkadxe+Gw8SJ8i5PUVC+ycP
E4+1NfZMI5up6niWPrWb5Mg3Rc/4oEGh0OlEDLLziePCACdadVga5N9ONIC4D/+XD27AuZ1DjJmn
9p56jf8vyx9vXnC4VrYcGzSeETxTazRqig1m0HI7o/J6qsjjGECLfWFhKRV83+5NKufEVXtLifwR
b/OyVAN9WDExcYshFtGeGtr1yKt06rZ/ZMOIX2eCwxU00D9EkM66jT0YbEJZ9m555QIIsCNgnrBq
f4FkOrwVJSJ8nAf6IssC5r4ABCkXv22PI1jVkjXJi1wBZ6XSwNi4spYTqpoTqg6aG/2bUeO/pyRR
cA3pe1pM3KF5VvOKVtXIsv48EQQg5UQOGWS3paF/iZ8dasXt7SXRQvdYNPWkMUjnLsaGg2diiBWa
iTay6FwJ+dW7/v5joieQDNR/CtYs9v6tgcradqSRKITVDNqz644RqJ4zSN80U1wUMEYF4ZUVOHq1
42yBDaGjx3cgJrxtndDWy6+xaNhxkMsl3Fk6Q4FV3wuqM/aya5NvlafhZXXyNnbIJ+cERfZJ384e
LOn480hS2ADfApllcX3P4YemVDuj0Elf4yzZ78adu4Et5H04CjBhiBUcA7OVQVriAp0RuzbEA5Zd
FRFJcu13KLFGHity+BhdHWGMemqMjIYKBc9e9N15xS5Pk9qKNevzzLmhXddKTltbMJEzqCJPpSPN
KZtdYYsR4+NOSO80gd8V1sUgpJUkkt2sU5RgtQsDajgSfxw0VjkAMlqnWp9GGK70xnS2Uo5y+pff
m87NVuNwQHWfU/Bc5TQ+SZDv+YOufsoPAoFnXAN+k7jjVCrDefsLsN2ddCb/jN8B/g/N3LX5Vn43
L3o8koHr5WMRhQURt6v962Wfu2E4oxZCahIeyftlF8+hqbrsQcAjAcKyo4SX0bqNVdNPucVVG0WM
8w+wwdJIm6Vw0jbuPn+h0gu2uU6lVeg1OmrqTfbZQsvfRQKox5fY1YCWBndyZYi8HIUQ+OWsUz4e
wG+b2OpphoJXJtho8sK8SJmKA8QmRSSyuN56G8vjsIgkuWxasL09xmBMQsnzgNPokKUBAcT7GxS1
1yCr8LqhrNOOEu9acvpr9/rV+7ZL+eJihufalJhrcGLcc5R5K6r0W0xRfxBGgIMRimPcFRA42kQw
Cf/FvnDDsuippMVVhyep2IGlALRQ7vwaRIvXQVVHrEGsqOwHSx31ouKWXohLLdIKBCEiIkmCian/
5qgn15he/KblmfTlni3VA+90l5O4wKbGwnt2nULFEFGBYPpMNuL06cfstw4b7YQEeh8h5qvURJ1H
5ortene4UfVHuVogmlM0Avtu4YjQNG1LuPxerxaiiDDdELGkFQMWM0uLBAMTuU/Zy6jB5DZFwL1u
F9wInzZZn/eVdf+/tXTTZ5aZz+rNgDJLdF5xPPVQfldbSssPv+gNPLDOdtEyRwoEpFn7OF/Oh8U4
DCpYTdCcEyqaEh5XVjy1Z1MMacBY6jS1a9Y/qNZ3dbs30Mc8EjEQ32oRvStHJw5hvQ4XSzCwh33w
SC7se0lTgfGGSnQ94TmBKHvsWRKgLi3BCG3MJ8SvCwRBbZpuQJx5pZc2DUmHqeI71awWpv9DKtB2
QKANv9dj2rgqogxqkY7SyA7uunSDjXoJPZ4Nn5vn3C+J/cZBK7TJqy0/Q03s32Qe//lw0OXoBnI+
NLLrfR/f+5fU4lmHrpYsndaAS1zltoasez/zwMS5JX31TSYKsCeA+fN7Gbpld0hdBBgnxrbJAoAG
+EET80yhFC1wnSV2SYODcAi210C3H30wnFn1EZLM1zWyX0uICWXsBA0D2z/2n2TW/mipssBtwZKi
bvFHLIWe6xHulTb549hPyrShPmy/ZNxBoNb8xoCJyDRBS9NDJ5reQ/hJHUtCLdjeNp8xE3KdnOKh
dRNaHOfJMf+ZZw+Q7NbrS57Bo0iGVIQxQFiTx6gsGfqvBO38SiNmIjyA1uHEWw6XUjxn8lbN+1Ru
f2ujt4OKE789A5FMA3YyAG3u6Vyg0xgLckqBC94mOs/Yh5L8qcT5gJd0QNxma4xKZ+CkA76N7WS7
wdUePpDGPBDkqY6RRC8+byS8yLrXFf8rzKumY2U51dutHeAtOdzweKvUsVUSVn+eKN1eTMT+v8cy
/2CMKuHGnBc9Xd0wJSKTp4l7A39GLWsHsyQxld3yrkt0ZlkVeePPm7Vczdu/v5friTGC73p9oaly
FxKUP/ySrUbn3Fqu5n3M6K25yb2gmpdjiA623qV3+X0jmnC+BO0W7Enw3BJ3SLPrRX/Y2LnqTPXn
MMZL+pCEKVSa/QqanhM+PIoKCm7+gysM2CCPPi1Nxk6z5wTgA403V9pr5PrzhPFKtTuw+ZdxmAwt
7N+UT6zY544nHRqaRmtrAcut75qp2D7IjpNmP7orNGRMh8uEoC3FO1rUgEY4JtsbHmXNE2fdm7E6
nMUzGF1c/Og0QG2MVQiHmVvJs2bQRhqEFAMeqptcwR7x9JN60jVm2PdDjsaG1sI/2R0vCFgG9ls5
ZOxRkq2aGbbsDQ+gOT69heIPfJGKGWfB6ZiThqd247UmQxsvVFXiy6+Gd1+aelRyKsV/rIjAUlKm
66A0JByX+Qczl6Gg06A4LkWcKG81C1Gy21tdsAcKuALf+HpBmVBoqtENLNX9Cb9JxUinR48Ssk+c
+lg86wT5CfPCe1HlMzkm9cpaFayYaKhgk7gjiHLxWqD0DCWdHMCDkUCf2WFw1iIRkMZiDv/SnuIe
r9WeRVUMWtqjIUWqa0wSVFUeYnd1IRe+ElZYv7y5hsSFNv/v7A718tcR/P2/hJiKYsFi4HwqnVYu
6weVwwWbsIb9XPa11TR6rh1EswdRj8Zz+r5j+2oyWeCUHPcq8QhdD+9THhY0g+W3TLtWKMLzw3yA
4BSZw1a4ydKs27nWlhSztDHYuuSTEujIuejC0OVNCeZNzBIFRkjW5/RjOC9mLOcE86R8zNBxq4+h
Mm/HB4iFh2V5VnA2jKNLDQRvvSvGcjq3DqX1HGE3btamGKl5CkbMY7HEFYdXyF1IFozs9NSciYlg
bnr+szHRHxjjTnt3BUbr4aLUNBoYq/2TSOSzq3klXLS3AGs3qsVm+uDO+n0gMUH6w41DPXM7hW5L
hVP9PsC69b4sV3JXPTlKtsr1KiCKCXg8fMfHPWlrAe3CxZVFDFnz2l9pF2Qs4pW/jEu5XKzfD5BI
HV/7kDK0xwtYOJQnL6DPWe87tSpwUneedrps9Cwu2KHQSD20PQDCacNfR/HSfgmUOJjHSaHLCW5e
PtSm8cnDAMp2Ly4kxAcxyVbCVwE1+GRIFxG1PqQdjSTrRmzWMBk1+WRZMzsZAyA6Chmy+MLoyeeD
qcH4K3c2s03v856Vn5M/LQADnk1LtpQtAmt2cRhx3AsaJkBAplQ0/y/MlMoHyvQygqjsekoIGyHy
NRGxxcs5XvcOXSSSOqwbSnm3yTsYghVAvIYtILhrHpEWfXhV1qK3luOR/2P9LP5YQtMF2/VJDF+r
0BXQR7LpE5QJOjtXyqpNbdyV1+2Q6nws0ibRZj6w2pXPckzRVdqlej7RiTRt4ABHU+LEmuCxp6FC
55/mX4wVdqsmAyxf+KDhsRXSMPpmj97Pn7EEmfDvdBndJmbQvZX5Ss6q7JsPkKyGe37tN5fBetBc
Dmdgn5WAl+A27RFGDgcoMD/khFJnhR5H8/U6b1CsWoTkQgjbv4Eiz/jn6FxyiZd7nO0r6Y6OdS2i
jdt/+VU3MB6URVMMljiCgmaKiGZnyOTC+2UmBaS1CUPnurrnUnwDDrEhKYJfKgzJOD8mscL2UKRt
rFMuW7riFTNnf/bQsCa4zEAxg1AfbMwDvcXfkkPyPGicr7SYd7neRZTTD3FtA/QMI6AsKMZtwwIp
cDZ4fDtL3doZFmPJVPdTdb0HcMCUA4wLwRlOcmPOEJ0WSzh1Ku3K08XfKdkg9yaPBIEuEYxRp+g3
uzfe3O2z+CBsJsTQUpk5NDaFtgNgdTqY1MTLH6kNSkSI9JQeLxVyM585uKWkcuYukOpYC0fuupUw
ikIpcoEgJ1FSKXFNlQa+b3yB0fyQZDOdC2gc7A7wMkdh8Xa/19qxhIeKxV1u4WzlQPUGevV7bgak
SHDpK9tb6smQjzZ6UGUqxPHjVTV59EumM4qIf7Pf/IjfwIJjak9cBmbBe3Gl4RgyfWLWp726I/qC
q0TxBWKe14xPqGzMM5Hw7u5Uuow04hqah/trLaSeHzM0FPrG9tIeTRlPxZJu7cz9UmSzCU/pXkgL
/7JZ09z8Sb+9PPRyVcAgIG1l3Nr4gVzdAsyN8X9dyq/69PKnnAXZMfyz6Jr+rMDkmAXqKqeaIEtp
DzyhHp5xZCyr3VQHCjLIK/7UwLgPpXUMFg/nd9ZY97LusWhqBeMXrp4fdckWXLJPr4eZabrpm3uf
OLt5UsgRu9FjLXoWlLYjWAtMIUdFcGMbfIry8vLK05yyEM8szc6nxW2ME3C2uYbwk0Y7/QXkVnNX
zhCie4KMAxOqdC/WJXjvJEMol8uxxnXPZoLr8r2i0/rcPzmHfQADN5qT2LMZVMM1kiyKjITVlhn7
H6Ig6BiAHyVIyJjV9k0DWrJA1C6xS7c7dS05uehOlkII8S3Rikmk2XfH3YLafyqqXq7yTdYFZCMH
8azMFi9tRGyVDIPGXFmHdu4p8XfH7Tzwpfam6IW0kCQZVJz+9Hd39XPTBqP2RxGgLK8HcvOGny06
MUeJ/A4lPBYVd6t3oOh159BQLDbI5d4B7J9plVdUrmzPyeTkS1SRRHKds5GsL1qpt0p3wIFoAkWj
YTb2XMiAga2koOQ+S0fpFZlayzaH6wyOIzJ6oZllOl6yBvD4KnBDQDPvu1OT2eZpPWcwVrJxRETk
D6Tm5YABzzShvkH39RqhxxC8XdsKq6IQjeknnR7Oy1ZftD3bzNTDOvjZ46whenkOC6M2Ie/ckWlm
/PkmjKLgStqzTRLV9nnHpxq1Y+3rqaoy1vT/WlUij1c2niV7U1Qz8CBTwEnffSYotLuY33grtmL4
z2vUX70HP+Gyx7kwN2J6wukQFDVKR5ucMRdcVOHj7qd9B+O5I4qN3UuAvlpMyxiw2mFynuwM5okM
gCZ9/0IMQAbwGyTKEDjURVr+DIPbQwKHzPT6vt8xLqutlmIOBBDDG4US064YxSNLw1TbkeT36/8U
rBo0wdBTmkBELzV/mWmZOoBSrFxDk2Lbbb2rUeSxUPUo6484YQLJzSsyL6hb7gQk+02dP4yML2u7
LxafM+KzzCEr+0rJcTp6UOzo33J9FpKlCpdKtD0Hwy6D7PN5dUN96/KOfoXjfgdPQjS0fvEi/GxY
e+aKa3K5pRACuFNt0hJYwCU5dvM2qYY0c5xYlwu4a7lkQcAYaWUzIIPi3OYy102GEJLQ3/8si9Qh
zSBrSxhOU+ee1B3uwBgrPl3mZSgFCsuILf846OymoQnSxNt+SmYuxRwLZqjB7MT7Yc6ZdlyciJyI
iDe87nBkZHn6u/LmT3w9WFUOuZg286pxEKqI5/FqhDxa1Jyt1Yz68xHXkL5dswXBgENlz60Ioo9K
d4QcUFxQXIeGUmxN23G6YkiurLPeEFfM2Xrm/t9JhkGJM3Urk8n3RgAKL0XrklbOfAnYzWxxXLOY
JcAeuak8nCtj/64zsc647JQFt1zw5PuEVG1J9WskkXqwm4JXfDmKV7hTJO5MBkfhvPzaIeVMlMzr
Ea5KOXGWesxi5SBXPu24Bq4qcTD4wYO0boPbACu4QNfcxf212oRpbPrMIG5Y/kdSesiGrw5EI3ma
9+jhPGyNbcMKzSNRlwop4ABZR2gKj9irVjxKZkA/DZsHF7kRuXKyGSOabxFVXqZXA7qMlBqGAkmT
w41RVHLopBWph/oY+oH/6GyaKQmgXo4bSOwiPSE8W/0bqB+Q6xkNv4W6k0XiQM/01khJ/1xLZuQ0
nKG9dE/AgSSr4OLWvUgGtKrSmHN1GxuRTWKv5BSALLjL2KUlKMMtDPHTkt1k6WPdy20qkSRpXDyL
qu/P/qX3vGe0+4hzzGhNlI3IY1UD95itMeh+N1EBTeDrXCA2Ty2OKQXdELzGBNbcfqqA/xByvAom
M54kSoQQ3T5NeIMSSxl3CSWQWAZFnBHhh5YB65nzs2ocw5y3PzegbrrGOJW8ZFGybL3k5aLi0ezL
UYXhTD2ptqjiLimOF9KiMI3gGFMiJqb1cz9YDztyeLXXIssNrQtI6kvl7qoE8nkQhlhdXT33YWDe
kcw6sFNiMdow89to8hE+JG+HLFPWryPjCud92WPMgCBk0CKuYZ6qrDHDcQJRRwDcL4AZQ3wgmOuQ
F8MSXvjZul8AvxFT5R5PyKEgmSKoUNQ0rGA+hyAfM4TThaRqDSAf3l1lx3dhI6jiL3wtLbtVv20L
drcEgjKac4JTGKkgGPQlZYfVIjlw6ZkgVNVIOWnciX5XUVXeRfG6obZtPlV4iO8FOuwViiJ9MSd6
me7dSaRYUN9bTIpdd6GL19+dlUkFWRr5PS/q76oCVRpl+GKK+TAjQqJr6Z06wQt1QjW1+z2ea5iT
nKAP+QNl15H8xogi1kMqKuCOu4T0GcsaUnz0GNMpwPVOCEzjAbghsMEK4ku0lCoomocTn8ieMrYL
CKqxEctSyWAcf6qTndW/+q9GXjsPf/ghEI/0tSAGVj4dYX676DKzYXF65OCMOlvDBEX/iG9/EjTy
7jC8OhvZMqUeE+hK1D/aYm+QP+BZT6qqIx1ZWizfyA5IowgqJI4AS1h/FChMtZE1CZlnvd7LFgbq
TuaVDdMoQX4KhH2ECyNE4GtT7R6YjE0n9R984awQcKJoqzkFE4E2kgOexC0dscMyzZJixNlvCRKu
113cZ0qmuuiHQmt0jWHSlRE6Hh12JVhlTmCm2+e755Gpmga6/aNVHMIPTVfrwcui2wkM4CflxnMZ
HfAidCfyLU0M9eJtLx4B7mYLIVap3wEChHGn5Dv3W7TbZqYGHMYD+R8vRXb6uWeuLjiS2mp/GI1E
63cxj9qY3tPW7QrfFlUR3MjKueg/GVuN85M4AZaZvGhvL/WIc6DZQM1VNQT3Oixo7Lmd+6khPufe
fYmkB2onb8mY4G4bY6dNySX2p5pvQ7WwOVIzv5Mfzt0tMBtSmGy1q/3g4zA5z3xrQZf934iU9W2B
5YzRjWwnKBs8yLDkP2bJqaCP/GOKZOfNZ/sm2vh/iQX+VU4dRG+ZP2PnRVJeSbkoSFmvwH6ruBBU
21qOpNEdydPCBwGk/0v454d3BLRj4uXN+N9DMjVOvJEp5tE5IiqZKTCiuNkjOzErFoNly5D0+17F
d28N9cjnvFDTrnWDrW2SrucRQ4/VihyUUNxvPccWUXln+XGUnr0QQ6dV9/f4z7kZLWqgFRwJaErB
k9K6hThTlfRO5CiSn215xlTfvQqHpIVnCUaQYFArRnFugeneZiWtj+9+5WOf2nOpj7Ycbx+5+13C
6V9bFFycG4nl861M2Wox2ii6J2JW3emuw75+FulF28BD+ts1WJLQbDciznIYuNFak02cDsN6reou
nbQoGuHX51MvnqdlOnokTKgcGoV9HGnJJZhzbAc/Rsb5zentvDCwq6VrMpoDWQj/B8WlDZLjPDFL
vI48skD0QLJeKQbKPdlJqAs/r+l8qatz3ImC0AR5BXtD2UWEpn/Kh6DOq1LFIX9q6ecMoV55GS51
37Dp/PJ7znTwkCXjFvpzbeukLrimxsqgekS3f/KcSqyhgVRQgDdBRl4UY95d0O/GUpfxap5hlPKk
zMwSSu6TNroFC0Sixl4Ucf/rdxOhsdByuyf1Xryuywb3l4hJSvYDpg4RpeQvsGrJCuMFWumJjS4r
p+YkvUcNUJ/yY+ZG7EGqr3Q68DcJcspQTtRKVtATY9L0rgLVYVi+cGt/D/hbUa6QZCvxMzZEvIlQ
pE5dXWMkxteDIpp8dTQ0R2D/6Hlnt+URp/X2O81agkvmiE6zB8iaAZZ0N/twxIkeZQ0nmFiDFFip
/e0He1N0sqwUWvQWktqGVFRgrDuXZzEABFbe2TQWQtve+auZZk87U5500QxdeVB6eWDZ1GGhWVNk
iDOjmhtnRWF93Zn5B/Xg/M5AsoaW67/9Hf8xQNA6vsqiXH70q76VeAR+hB4r9XH8nQfU6vkjXuvN
faSnXMmlvxtcu7z4qjuKlmxZ0A5ll/ioHqdlsypsAXwwMGF9BJd6DNRwSAwmyjbuu+UHRrDG0Lv3
wsjXqgl+x1pU6Jyfeb/zGkLfbDQ8nnqetxeiXIUDYqoVBgvDcLWPHhiWjcmV2YlLOqnLnP4Ha6Wz
XD7wD7MG/nZuFl/bMG/1y7ete+rAel3+5AGFPjgweAoVBzYgvRexQuJiUyY2UWO6+U8E4foDysDR
vsKky39lwvvXSJlq8QkHRTaxQfeBex9FAaTnjJlCPN2eixQkibzFyCjQn5f7KKBDV2gJirmpVjaV
Z5MYS9Nqe0qk9Wf3XY/tSiGoJl+XjpL6r1gNwfbMcHNFWLqM+BYOUREwsxPdM7OBxt9yCf7cAU40
WeTu51fQ3sYFxqBIUe0HxXRJuTVdOqOkED7IEOstp4mI7wX7XgC0osu8q4fKtBeL69B6mXxl/0mN
WO/CoZ4zb0Vfw+BNu3MmjRpRJIDAr4Equx0DUtwZnCxX3wOsP6HiybGYPmZ3JeaPAWcQv2KlWdro
883SQ0Pz1EzlKC8jLGpObOOyrCdvheZ7RZcgwxUTwDoEIetW/+pCzf+o3GtRdfFpuCx+elyBIaBX
SCd3BtpBJJp6Db+RF8UNR1m+vO2rUEJ3CDC2roDMfP5dzdjUcIG+5SEd+N0QAZLYlJHIWMX7zTCH
Hq1WZNm5PigQWJQyPgBzRoPcQ6K8hDibjBoeQchJuz5WMtkclUrscJz3aSQCyeYHUdWwVesIh9b4
MA1xbEtjROoRVUCNAlW/G+DXuccObt/c81cjf4PW48lZeZUmKU9UJ0/p9jiYVV9lBVZrbt2LpHWA
XHCb5usIYfmukJuXjS1wnO6nsq7sT2wglW9p/SGp5fz03Zeyq9Fn7K1i9/nIjZU1nRpPLH4yR0sN
zSe6YPwke8q/9YguM4FtvxtOq7+PonycPgCGyKz7KoGprTeRAuszKiL8czJWI13W3F/4DDvcHhf6
Z5GMLzAqunDmELB7lfibk/VS2JN5paGu6u43qCC65KLVur98uzN7yqoMuY7rNa0LUOLWaVuIFOVi
eF//lsB6RXaPEMEbYmKt9v21w3zq1V5DvtBfINVU4eM/dWSyeOyexCdBFxh4LA8TxieXXyPjoIDK
iZD+7Ta4lXF26x8aVjSixBQBYSXntAFKzD7N/0kUEs6sldXjVqz9C84VNbzh+3e93QtobGtYbtio
0xLiR6nSGofA+Wv72MDrgskGJHGVrOxc2xm1EpdHUVzG0voZG6IVc0KXs7sMSZx3MJhbjN5BBukB
EeABXscrbigsrMYo8L1QNVLiZdJa6zUNBG+YnDiTdAH+I7PbwPyVPlG+qKOb0cdegiAVkXQaO9LI
q7PQluBICkm8dnBe6ckSbp6e7crtfKIluCz7m1BlsHw8irIzmJxppiurTwgQAxmEzaUAIqev2rYW
WKz+h2yc2BkSHqrGbv06wLsrRaXRdAYKE8/qs/kor9O25BmWR8RItJj+Wxb/UDm3ZV4V18lks4wo
I86Y7oApKbyaew3Dt8PG0Wo9A7KqdRCp/HBR6QOvJBSZvYbfYKbL8DFgKSWduaq+IaZ+r+GFhQGr
SNn/kHHZ41VDcejumwNafryBNFckzW/ZwhLiz0Wr6qAXnC5njxjpYqviRrAmbocJUT6lqr4bVPXU
rYKpT5AnywBVW/DhyPJ5uA61j1DZccf6eP8YUdXSAPoukNxlizOjIapAs4PG/I6+t7sRFhL2xNBq
OlnuPfLQmptX8VDuCzZ8tOBUunAUH61ymeHDgxsm9wUT34SwE17V5CAYul8mWTGeXJXRTm2esZmj
0bjubzpcnqJUrrTMntmzsdqqb6fxkIxgltWYstYsZ1Dm+rY6hNquRfq5hnaTRs1/cw+VpoHENXQT
VxXqKpQhsEahTXKXY9iEv5O5sYEni6G0zHyY8654q1Ed9004OANaW1XLoIyzCWKQqsPAs8mBz7sm
0veRyRYW4StlDoQDhkAyCJXgk/MQKJA+spjGOdHtgQrNfOPauFeGiSKkMWEa0fHizcYZQAZDH97j
B07JONqyt1blk+cmmiqRrjJURhZ+LWnh15Rs0+1G7vVPWe4UpApiCw/OWLad6aMnZbABWQgXvjr1
Co5uMUb68ARlDYugygTbE8NNQhhGIuldk2AnmSxxi0vzlJd3AKuh76NygYKmrzIwQvWY5mRUN1B0
2AogX0zyhJ83YiZjAdFTFnapdJULugC06P1ysl7yMlxyDvB27rZaj6Fg+Htxa/Tf308xayqv0CST
XDfpGRpAo2mV7GAxNlzjL8xLbfeJw4NHWS8y0Hph1JnyDb2QXO0EUy4Vfk7ZxyHtxBESGCAsqaDO
3iKY1aURSJIJ92AGI44IOOwR6DXvUbGnV7WqMkDH7RLd5b2n6jyxOfj55h1ZzvLgmw9cP28IRLYs
5Nxd3vuzQvK/B1HP8Xp4+JPmSZHEZzneoEH/slKs6/Jcewes4WbBILT2ZD7zT9QDQmMA9dLfQRmm
R5OL13A+A2rP4A570LhrKXymU2KNDIR5c5gWmC1hG/W57M0l+o2U8XI591dv+xzG09a1fTcwYIQd
cEVBufFmF8IcXUjPIf620a9naBvNo9/igmto5jbf1gS/1Y+rYq88C5y0JNtg+5mz7CUHVP3mFIxk
9j/8brho8kv1A4f+8Tn81mwrY07nt5/SkzQ/hJHndrOSWJgfLf0BdPG5IvHrrPm3UqaVprh7KTVM
qgkIr339St9Qq9VZojDbQiKfZdaHOBAKLO/Ns+kii+RCXDfyDAyJ7MDp7e6vrPc5Vfj1BBBjO9eR
JFBiN6eusPJRgv69hzoVP8D1pkaxB08vPseTOg0Bpd5zBgv70SA7haoUpP7HqueiE2B6pMivz4/k
Iyd0am2dpMn3O3oWKBpJpTkyvQyIszpVDsfz43Nl/zrjqEdmHN09KmPJmKvoK2qDkj8dROXZMiUt
egcThqB1ogjI4OBmB4IMfgWaWNQ3/UtM49U0j0g0PhA5S+zc6O6QwEZDd4TgsKvT8QZ80u6Zodlr
XXmsczabYlzg9yLqQ1ZvL8RWBPToEc/ZaUTrKD4f+GdFnXZ0Vh4/j44zlMUDhuuZjtiIJpwd/9lG
qyFfAo4EMWY353YfJ0tGlAi+95eCvX66NRBzjGkbX5nOAMj1OTnFw9U14V0WHV9vi/KqJ8wDvkoI
91pys+N7Vkb4KFoY5b8/NOTFC2dgl48icOgkKcSLBiAznjH/lfU0qkr9FTWZtCrp4o9/FfJp734H
9cylXi/epSE3lTw51nrQbD4qEFyTSCt5cjN1tlZgEqu25fury7jDdK8LhenMZ3XMgxPkO60+ojXo
8MHIdZRsdayEEbp0NUHTAEjXIPZhq4KDQ5hvsBw7wDszjN9aVsd5/UdzyBiNlXaI5j7kn1qKm2K3
O6GFOtcFvH7tS+BAApxOp8mQ9otrASV2P3CZlvslhQV6rtbvTCCH1kw8q5+obpDIDzMoJMXcKffE
q0N7BJAtBxQrbwD1KUd37mJMv3ZmC2bzOcACj1+ubLmuZbFERuPlAQfCWjf3Qmn2Q6k6MK1u4Lbc
KNf0QCzvOonkqBGJIxChlf+6pAJ8tl3qsmeTYzo6Ba48E15Frmh9aqI61ERk79ajTyGcwy/jQSqD
0tjiALjApL0gk1I5M6FFgUMFNQ9bIu3l+VuJFoHuiL/BPaw14SEmE3GGHUlTEXWQ+06+QJdAtjxL
odub/jSDT2Vi4MY74Q3PvQ6FtQSs4noI9GCXcF2GRbMFciBF/aWQ8yfjti8tNQAXAAEytUeIMEAw
StNp61XVm1/D91e+ePPk3WCLHdHmZ+zHbu9QZLGB7iYSKiaDIs9S3Rqko896odF/dEq6jl4yKZAC
RtyjkeUH/Uz+8U+zMY2V0DvrL59y8xfQWoNlTs5pg8IZ8tTfOfH29zyEZV7Xk9K39J+2enACQBOT
M5LWY0P2UkpaQgBFuxp3J7y3mOhYU+YzgFdb6GR/jhneMhMVpHQsPj+XLJBXlCkY+onBQM2RhKz1
pj1+dV9xWwfacXKv9FBiLcZe8OUhJrHuF8ynj07bbbx8zY9uuTo0QvaDwSNnkPSzLbdxY7vFLFAc
4H3TWBw6u42rJ0d0Skp+hOyhbLN/4DPAwh/zaGRUK4hUvbZm0wupa8BTMkbR5MOPPAG/e6eIM9YY
cZQSkiJzskWDjbinct4xC6t46uhtYoqbLtuVtW2diahUSYOE/1gGYdFN/K2uAFVVtvQ3p35ND89i
Tb6YX1G3tQdBlpVk55NJUiiXzicvW4P0HqC1VC54+Nx6iF/xdl6tGS4h7ICvEdZI5GHIZfg5Zaz4
zyFa5sRdfz8Y7tAQE+NRJaK3CinpQYW9X0+NVE1JX+yhX8zR+I4ocLggE0NsS4ldBNBPlEebumg6
iV78OqtFzFFuDnQvTl0n/QgWDUnGjjS6/omdmS7nDSDKbMQPv9C6A440WzWxBwS0yXOZPUqVuiK+
EPT84whN4VAjGRFB9IFT4GKG95/MsU0Kxt5J7IHPQZPKIzi4PfhAZ2RViTzd4/hmKJRdwWKIU+9V
bo36s4jdEzqr7h0WOD4H1Sar/tiHNI7CtQ3AHB/Tl8XcT7FeG5Afo6UxXdIBOcvQxazoDvkfN/7F
7YN/KDocUE5u/VKYz/Dz8WFaEIur0ILSW4+q0lArnc/IyUpEk38bmt9IgdyP6BW/srmz4SPVtD7+
mP5UVlJ/Rw/mL5jmL9fjzPg3PyN+ovnBpADBrXLNxhbMYAIJCsXv1FWqk5zpqJBrQg0ihPEcASFy
vX8S/sOb6qQ3gJnc0g75eFtPc91WRurWRbqboc8kOUIGeRTQgxPAxzBMJFxSSBQ3YrqOCoqSYRMl
T4DUO2LED38dyD/okKTVfBeXp9OkGj9D9VB34pqYjF4rLgLXiZpbjR+ZS9ULDHd/oLDSkH4MmKm0
SOseowO8s5xHD3ks08HpKucfnF/Ib7KA5i4AEp616k9g34hgg8Iz9WoTWX40kymaCuWl2mXaNaew
hVEUF0E+LXgbLMZT5ZqYzV4Bh694xhJDvzh9VarIoTZZIEBFfD2FmmP9mTEt/6b8TnqMF38Fo6VW
TnONXCrCTnkYIlTSzl7asl6AW9LZvdNcnbbZjYuC7rU1ZuexaoehkmlAYKFEYwPBt7e79E7g21Kw
xdd1bW2QumZgTTQfDKFbyxsGwd9M0pmtuGESvt0P8crBtR6btQ/nL+uiUB/0ucF4KBnwxIzbGEqY
IPStLsqcBhhEfMj6PGQFh+4mlv7VkngFz6rYfnnV+ftsLCuX14am+p0Cekk+EcZ7ZJ4nJNeDG4Pe
fn4JqfzKOauQ6RCEet2pvLSJ0Fp05A93/dKExlD6ZJkuXpIpF+PwjHVYnyzAEF5r52/xtVRPGBxt
Q1B36qolApfq6ZlPHnoMsXl1NjcRWRtBaRpxSxhEEMtdjvHh/tdoI1p+ukMAcHxyWKZyQn6Ba3SZ
Xu6bgZyPF4qE2PmeWz0fUC6CrWWRG7eGIAJpORvJ01BK4Vdk363JUVAj82k2nL+M7GbrDVui0VeN
9NUDmt4IRdQQ55IEFlwOST5VaZmLd94wRt3nMakmWcqEzRqmJu2fsEgAZH4DIDWVEpg+8ac82j24
n8WDUOLga9pFX8IdY+Jwv8w+c2Pf/f3+deSX7vrUZ6Gmo5Jpj7NybVjZ4gAhpdrVWIA0MsNS88e3
MLo3yuWeBBoP3jPTFp0UKf+ZZ2WvBWlCLKFs8uK4nNM2LuSuBdRMfayRj6w3pDzAJBF124YxHY24
ApM1v+Qb+fi9Fl0Z8o4s9RnSUtHqE97OMFJqB93tTOI76l0ONnqAFfdNoWCjb6fl4gYFB7ltS2ZL
zsCp2K5GM2i78IgF8T5vERWS5/vuq2MJ0R2EKf/Hs/G5u1Qkc+rcaM1wK8L9EW1eXObHGD5JVh98
Z63qtRLQJsC40DVIW6Ln6y1tphPOBqJww2taXFbvBOFB9D9xFdmkK/UC34VO+/cM3CAU9f9Bucgz
A5icNoqlFJ/ag42UP3ad8+LWZAuyVsGgPFHLo47/GiTMiTYA7hqmoqbDXNjuPwEC5DuHXhLh5Yey
vmuslQBfke/BHcoWJUano9vBKVVVxAE1+nUnpxVwtjvPB6RH3+s4IWQHNUTiKaw+BZDKiQhX+dAb
Oqo114w+PVydFCG3rqu2DqMzfWiI/ChExi40AZy/mEwTNSMyPQtQuiP5BQ0QUrEYQ6UDNWXMqlFj
Ezzy4A0oea+meX8nxPWuKssVrk7YYPjKkFegpSCj2ZSDx82IvvmpLQM6oy0mgDFr4qQSmFeoiqBl
ZJ4B6MieUPIUBAGUZvGCsk4/x9Z5YzTGTGG9dvWvzz83xwd+ALgCEv5tiXq+8/hTuYw0n6mP5ZFZ
+GU1tkvW3pE1UgSWnbQ+kfv+jN86H2DloXscH2g7lqYeoG/cBUAUjCIa/CGtEsiaBU9FWn66Njaz
nFbHWkBcCco2TW2RxcsyVNa1+X34/TIMk/KmjQVZo3KNK4uvnSXQ4gf3bCrWr/hgAWnMJmmv2vxc
jgB4ODhQzkJ1gWdH2f/szBHLXRxcg7FolCh+dMd2gRpcRJfqaoTmDfI5LKvELqUnY5sBkBmkvYrp
lZjClN0zwoJRGWJjQd6gRaywhWdvHp+gQP3sG+IE1hvlZaJtDxQHp4h8NpnCjGhWIFoIwE/5L9hV
/YSocBKCvhzzVI9siqBoE907JaVfLfBrsgcH+1yTIe/c7S9x5K1PfJFnFTu3uOOqq1LcL4ahpwSm
x/px34InYMqTjRpXDnQquLNNGKGvir26/dT0EhGQEzFZWbVPv4iracUdrzOgEbj7dEZJXDhW/f90
X1tIkmQ5xa5F85pm6TUp6LdmM6bKvtdh05dF2IbUZ/EhuxZ9Lfwiiz63/ZrIJjRamexZTMHmkN72
rroXs8sufQfwPVVCZNBNilKt4H+ESZYasw3WyXv37d49aX7JwKFF7jHgan1jWlm/dQHRSy6wWwUH
xohJXe91N36NK0ZpRQR+grrgIRSSqJ/sYjXj+8rwZ1Zj2dUr1+iv/yqENzBQiEKBQSn1wDYYLFW+
h/U7DJgtGjMUK3zm0909eD0wOmTKrJDwYnwbLUO0cFLiJSwPbUV+k1t9JX7ZlORgB/hPOMk2gnZf
Mqt91S79buwvPKM6mf5b9rUfAniHDU7PSxzhshPkQcKmatXqi4uKI6pSG/nFV+g0HPByDg+IuL5x
+8imxDxOfQ9pDZHqHX010d7y4MlpLQ5XokEj21pQBNXFdJEw4Ke7xsLoJKNvA+VaPtuJ/u7ZDCUr
BY6hLDAC2APdFTUtdCmjEB5s5mX0jwluaYzXo7ehBNqhed2J2sCWTv+Lrd6/5wSnmlcFMkdig+zr
vUxglFt+BZ/0gVGvPKmBmqFfro3u9uhqNKeopramSSkWXHyfo4N4/FFDc3ibaTjBjsXXKkOnHmnf
LC9bDHOJdckv5LBbHAP9Do+S/3PidT3dyWwgKzHsZOaHqobL1Wr6yFIAGkIxh29PCFj9YW+MiH5R
Ftt3a2kWBjwR6bf2tUXRYkMige/mFNwka3ScEgJU6iyjrNyMrhugnvzmR3msVvjcI/B+GIBgS7eP
8tWM59QuRomObKht1CPwzmZKCap/9DdjpsZvsUlSGpqiaAC1Sh1svKTr6aDtUZa+/9yl17JomUTy
7eyLcbxSteutlEdnxo1tX7zX3DKtXt5u994sm9G3tLRolQ72+u4JNdl+ksMamKffoM8CJxqe8S0F
r5kPXtvpAwv+Ly+IPo/ybtx4VgQRpmnbnNv5BjjdLU+uZEc2mOX0v6Nqm3A5XKHVBQ4ww3M7RedM
eFRE+5LKhh2Y7wq1XUsOWThMebx5fXVycnaPkM6RM751DcH6ojp0aK/JPELY90pW0em0nyyj5vbU
EzcUrxi+wNR0mK4e6mfw9HrHkpIYyYIQqWqWEe4r0nYsXv8u4puJUiMeRh6jPBa7+bxKav73Oahn
yXK3x9bKjRHMYzDWZP+7JZysjwnFEKgTwa/ugMWgDKpBzu1krxJsrgzt0L8YZfwZxyji3Ht47tLo
sj7S0q2WoXdxuZXUyremfwhCd0DMGgIivKP8+RIVmguMctJYGDQY0ga5bsWksV5Fav5KXQQnuyvQ
6PEvW1noIVLFXnLg6w/pRLR6optSCzTgWt5GdWxXgIaLjvMmryNxSoLDBXB/UivwzgMVcLBCHz15
fd4a2bdOXmtIgZBokdgj1OnYM8kV6DfISuYXc0Mh9OpI+afNRN5kG7E6m8eRxEdB7fY/QrIkMnWo
WcMvgFha4cCrTX9cW1RApTWuNzErmq2kESGj09/l6JO70A931gdtVRqIBig9JumGYIXEihiAvw3H
wubGSa1QjpOGqNaCUv+eBKBvieaB8eOtewlnIk+Ds5Budh5Yf0h5NkK3ndyIaoHLFFCxzeOg7exx
nKD7CDHeucSrHbsswCTo0/Ay6DWULPyy9TCa6ZDLk6b33qRUPaV6q+esRwkN1L832EPvOISJlSoG
9fUoFQVD4CNworLYeZY4tW2a5zBgq3EwIPr+YErYE+kz+DKOftxbqzCjEBJwVHGs33aibsL8rMmB
YiB0btIuchhtSchjc1k4RWy0zDKSRJD/aEGXSNTKkM8zvuWq7dfD+qM9rpCWhG2uUZi/ncaxTsov
zC75Ey31v6dNsFwYdB2JojWx30EbApZVh+ZYhG1PpvbyRxDBIH+KKJYa3TeL1961yZTHnqE6/Fp1
46KgHEZ+ZE+u6s1cSOxGeJ1IQvyrR4TGRi0rfAqxxXthnJAvLPLWsmFbzgSm1jHJYmaIiu8rgkJf
ELV5/9b6EO+0HH0ZXzbi7sXB+FVteJ3r6pZSBltj1WUaNrY/dww3PYVB+7oMIto6V0pKrjsixCkB
E61HRpdqKGKuHgpdmzDpDh9xYz0sWmR9a4+x+SveJfT6u7fbN/cYSCAt2vQTMXsk1eBGTnic8Vz3
sgjTXXe+s3IoC/ODPQR7j5FOrqW9fY8wtzN53ihafaC3qc6r9Nxt4GAd4CDqKU1DjDF7WrJwF7Pj
pI2eGA/L8QGVk6zY5f6vhWcvH34aZoAMdPGwCtJs18GCOvEn9TyoQnJXFU2L/4H4P9jT6dZAnyJx
AsIqF8v3b3XMWowiBDZTxW2ynjxArChUW+EmF6SncNu09He9DHuJ+sop3XQjXjnnIO9ehucHw9X5
rLKXBWtvQgeT7paIi/a0PP8uuzZcniPEKa/ahbLcY1lbGN9L76wSn6ul+p137vGwGo8wVAcrkUPd
NSq80pQPf0rXRYwxlXzsMjtywxuvaTtw9JVqfMi4k14pgtJJCOpVTjXKxM34ED80MNK3N/QpKR4e
8xF+gruvEowA22MEf51srQIlj7ulp/X3AlAo+1vgxO2QB9W3bv7g9J5L002R9BUVadKSItTKZdQY
eim4YERclSPdL+rqFGeNN8NLudXH8EHZdhDDwFq2RnBcNw7sMFUje+7Y/P3xg2IFf8RFCCcF1kI7
SRiLm7IAFEtgMBY/Ypf25bQ4rwCQ0BSBqD9zVkKThWlN8F5CkRzn9PW35I2hSu0DBUUkeL6tL4+Z
sEGXo3ma/Ylr4t1e+0iM3Dle18C9vOf0U3XFnFPubfOFBcNaa7Bc152Z09NQpgPKxZqsR7rDSCBC
ttzZXVRYtg48C2GJsx4oQVXgNF/PxR/IVzz/k1xN+2YAHKGqd//0nY4KVoZeqvz6OCH6jS1yo7C+
SeckhuuZ+5jLYHCD0HE8cAWOcaDoeP4cYsAm0QYc36WwTTfetM9LAHXmPdZTRKNKrwHi5eHMuoLO
lqLOcxMu/vUah9o1hLUKhEtNZeKOJWlaMexxUaYMjvUderxJxgwoqi7d7t5J8CallYn9SzHfSz7G
UVSFmXPltBaJ230PvxkRqePTgv1fPgA6yn8P0Qrw5LefknsXyJ0bBAgr9NANb5OwB0yMDTBIVQtR
1QHVSf8nBx09Wouh5BWWPSQCHrwEQd3pwWmm69xPq+erpDoQmJ3beXygT8BxZrn0NK6saYgZvKcs
HZYWzuEU8tK9zphCX3AuuUe0UMVjZfHRqoe9YiAuH/4PW8ekHFzJwqtF48g3aiRRdf2F8/B8JCRs
Ql8cP1OFmLto8zISXzyW8Q331WMnx55z1oCgtO68FEFyDluc966JTII3uJQ7Gx6UMcspGSwVYJW8
/SVJFKYx35oWZwRQ34n2JQbUEMcsXY4JGJiSCXnbFvIhuNdAPpfdnVNjEmWLZwSKQSdr1Nzwp/9f
Pa1qy1WqV9DfarEE3oamLGCKzhPGCLKMDlv4EfCn9m9v1n2JCTbO860w720t9qkNMm7vaudWyEAs
a64sr4Mqdy7+uNM43B9HlI3DDOX2ow6uKKILO7eMABH3TVQcIoKMZaPj8cw0t1Ji6/GWThrFHQTq
BWigbAjlEgGGwSXbHU2dCLrWjU7g5qz18GlmGkfVhrClQF3lPM3SJQOACAP8vU8Dng2rkVDCPYqT
lBz4uwEXxWKs8xbUyOELPkwNFCeqhWpSfLDxS3Dorh+jgSH1+FAZvrAQqHjcLmbYUVitg5GtKUQZ
+YUMm5fANqFd9Zzzj7EoxaQy42WY2VczoiMBpbryvaPkFwIqjos2Uqd0BjHXg8bcR0noa9C5jcSR
J2mS/XCwnI+Crb+H7KvzDqf3xOx08lo94dEhSbiYHRAGxWtjwYAbZXKbgxD6gqzo6PjXGvcvaR+g
vV1Bm/6mrhvd+cxh/MEyFJtTMhk5la2yUCQbZyvsFSfV7KrBYQ/tPae0Ih8r3cwUT/JXuB6uPRXf
iy0gzACFTrDZrPq47v38Tt9wjyfsCPMQoN8LQbWbIqCpn5aF1zqjCcwZeoKqAxa24lNOSRxettts
QJLl4Otf+pOlWFD7cgXO95s9jnhijlN6HHgedUYgOkZt8jdHLCdFsf+VsPyk4CFMlppw6BfM3ha5
8pacxurI3JyM5asFt3647zgBv5Azktywhppie7Q7tcF+luEJWwyLgZ67I2HD+bi24zlbZmIkYvte
jrPX1D+jOXwV7m1kTkAdUJBBhn7APe0k+RKeqCy2t3JMEuDf2xlwvHKkKWfqmZ1JppR63qhc0s9+
rJ5IO/clZbypw+LidUA0uoFR+/MRdXxNdqmERvLrMXhgB7UNARtzEkZ0iPzBQJphnw/n0x8PUIGq
OOKDZFkvDNZhK+tAW/dTDxf0tmw27Pjf5bN0GVhFJxoFNuASQOhoA/nDx7PNcduY3TH8welYwPwZ
D+7vwGMy8A4A//C+K72L2MOM4KYHTuDLuhaTypTi9xOOTn4tAN7j+aJ93AP96pUT99FwxD1VZoYU
oyjkEZFtVMmOSS9UU/hBitxhaTEti0lbx6BayA3aNI+QOMGno4lK1mcS7F7mto+t4hIL20YHwQVn
NLK+Oadl9efCA0ACFbEoBHjjHARUWKUroigZgTQeMF3VWs5CkGwu8SsqTUjdVpaQ6nar3W5N+LmS
WbT0ph19N/bggWp/Hbt5OQCChJdSDta8lOqqT4ES9jCGnk7jJkoN13qU1qNvINBL4PebVSvqbdIX
YFaNpcRWKqZxCWrlR6V4lT3d2RLXSEogbOnk4BRavHCOm5QI4GebH3pBlSpEna8tIo4ZRZHR4EEm
WS9HYrBPirp/tLtnVMp1CpWgO6z5w84EfswmSQBSyHJwl41py3/ps/KCczpts2zpdikqHg92cxw7
dyKta19SaYFgt6qa2X4u6pKxQCCmYE8yVhny2lmtRoejG3t+zp4naAnVihfOSI26agj694RAcwx4
tbqdo9aGMymqY9l4bwFIJGBilvfdKJCgtaxCZbnIJ1Bo/68d+wPrX68z73Fmn+WP+mzIhNdRMW4f
VsjKfiBAeM4DOwfkzViLm8Lixo9ONO2N2zcKJEDDk3bOzjih8RPdXe2lgHH5qKt9ioyCQNU9vlI7
VHi1oMMjPdKnDJVyqdKTbPUN9HBqADsDmVitMj4LAovJZE5j1/F9k4PlbZmfG/ywLdWx2jJO0q5j
y4Ffq0/eFfJ/CWjMOSggbHJNgxyACqQjk3fYLD3Rg9JdnkdxVRc2lXDB2VwA4smcg6HqSaStft2D
0RYC8JMzCI/GvunxKWMtVonw5m/TIeTrtCLOAcdKVPSJowUtN0eD595RLJXWNkNWJS+CfXgEYVN+
DvdVER5/sxDJRL2m4PZ7LhKNDGGaxtRPcZlS4houi+oqtzAncZ6b1DVkbPABm4aDpKdlldMXqf4n
bC1zoHa54JF8cFtqbkupvRWwZH8K5+z0xrgWmXzVabno90qXeXY+3BF4XyGD8pGTNcvzZk0fd5wj
mWENiq8p+S41VWFFcXFnh1ahZBruEKPV7uwX3rhrUbbIl8+/SPRfd3U9m6BoP4ZLL0n9kIiGIokl
0WquS36JhR/ck5QeNlp9PBv+2uOQ3R3Qedg1+HroTBf+230Oz7XEdhy6v3liBNqzuMlZUWkjxCmJ
VOu00CJS3FcqBvhlcUto3QTnBD9rdwFQ4a/YDHcXoU1A2MF0Re1Sg/pbdkQETU9xkw65JeCTlV3c
nHFAjXeKWdd7VLs/BGV8Mp+nPWeb6FSyr5yjEbOaRsdb371pRG8nhkkU4oJ3qcO3NNcwyzWFF791
GTbn+I7mTntyHD/7GgkxzoGxzNXy6xFIMmigHyQCGF4JkbAERUprl0zBzXBfk+9V8nqRWb2pVmAt
9ETJSIgoyUdepzHYmWL86R9LsHipMau8nNzuGZiP3GOilXS8Egx4kPXW15zAtn0oil40sgYWBK6D
0pMNG+woU0U/kMVtL8l9UbjI+y1sp0SCaFTYF0eznLJCMY0Xb/8kYYPAwDdNYQ/vzzqCdqXl4MM0
ryzAhpTtUZJVx9VQkST0BXzDLb6BnJlVZytUrD+G7JerXltDBxV74sVlooxMYirBpdUHEzdvuzCc
ttSfb2ywdv6kZtIuzlNhzzYj9J/CuLsGMvkM4wc1rtlwQJcNPmnAyZprNtbd/b/D1Cq9U7f7XBj+
MVjuLSBNB7UfXrAy5nBUxcSW++FgKd9vIdz/aWtpJKTBOeO/M7QJ6a9RGcDhloaWktQkN9Y4WEjD
XyjAfJWIKVx5Di1PpwFS6WOYVXzrqT+8zauc98Sr/woT9JqNlJOYoNeDcE90D8tZ0RD0d1WU/Oao
06xRQdL8ka2poBXReRkstjqr2VEHIanmRN5KAv2rBus2b7C6GUy+h0oHd7ywDKxYZ5ok8n/WngMY
YI39JgjlfCbWv4HJhZ9TLyJSuzor7HstVEw99aABpZNWgQjO/2diweg0g9BttjV0HH4SSWDZYviI
aokuNRajFeTXtDaSH7WvANKqoM54yHdhYV3c/6Zla2ITg8ZhB6g6feuCMHwqOX4vj3wjpaFg+8TS
5imEgRU1odwWucFOWK/RI3f13cJsQWfCujNmTU3hyNlZXe7Fw0g3yTH1vme1QooZBIXEeFTrnJ4b
6CGu5Fu0KpCV4kWtadZoF2JOJ5Hm6r89pzJLxrttSF/2VMBAsHsOR7Uhye1nv0BVT9mGo/dGu0em
Ffs1T94JkMsdtypDPZIp79pG+srgZNFkS1JeRYncfaYpfNmBePzn0Pp0ykM3W4iizVxdfOReEV6P
0l/zFa1D2ew899XG7k7LxvGcWSsqIMYVGMPuo/GdI22u18dHuJDXRGd7/uQAqvTXDTAh7Ip5Hx9p
ypf6iE5oFEXzhC9XdtiSN70qFf2nPIb0Qwxra4B8jqTcE5jv3bkhIm6CTnjDSwPJLMW4i0B7ApXL
wZh1jZXQs54t7heCfV3IaWTJbDhgiJSvypV/rf6UG8HaGbLBTLXT8yZxqhGKXwvw7YP+NYO8WT0j
48MQ7zJoWEicFxVEHs3I2c4FYKQPXzslEAQHe0RtoXNipsRMsyXKvqilNIhC+/ZbcXdVy5WX8iqN
Z5cDXHXl/NxbZsJximoyhLmAWp5DhzC5o07z4P3hm7n0fzM7fNs7jUOk9dUyrMAdvn1a7VCPLSgt
Dl6u+DJoYnUTSZMykHBLp2lDpwpnzR2R3gohPtf6sISrdSDgi1P+0hCvYVDOjY6CB+vUs/SFONlQ
h+ntUcxuJ7p143lVUJTCSt1ANedG19UyjdVZTgNBbM7yrnwvah4vXXBxdlfHgBwTHNBZk81HeGxu
sVHmumQBjvMITkcnz7Je4pyNAMBEk+RcHvCkRhQCNFtMcIVVIJ1iKTVECUhon9u9/qjF7wWlfZyd
BnWuwJn7akVS5xXWgPSIjnM83L8I+LYbtI8PCz/xZUUQBc3A5onG/VeRAcEK2KwLUOctXh0oSOzT
Ba2Uq4ilYzFafYAEP2QC2QjkijdEGpUkPZmjrPNNKoTF41pVijY9DFTF/HNs89DJKUjMEOYK5Aw3
jrn1VBofzfcTowlH6hsEJ88+vIgrPbQs85+Y61KYQP0F0k2xXw20GOB16m3wi5/WtipS6d8YDZHO
Utn2T1wIiN+qe0jCvB+xN4b9CKDcSruNsqtaIcEgWMvSPMce7WmmzX9je89f3ijVPxQfwgFtyY1g
zmJ2Yoen4DVhyqZnsVqkvZ/t4lf9IyA0i8UEl02NGFI29B715ezh1xeyHQDN+HnjcK996fB//2Qd
iTvnEzvi6j9f/eJ7uBz71YyLXrxPN0Ts0CJy6wIA+RkCDdX6CQtEwOg65Y3+PLSYoSbyMr0LFR33
BroHooL5h3et/EtzTximFFoAhfQ6rHZhsnrs98UnZWrhlUfa1vO6N/SgTZG3P2AJPXhCcIiP3DVp
KNanLRl8b1QSX0BpzwmD099pGcH9l0JcfyF3FDcmBxMyVjrf+Zgrjorhk2WmWR1MyvDADghpXJZB
kJnRHX1ID3c2iO+GhWmRswNiyvhUS+SIjcbrvydbiyWpwCVbpxc7bxyRqJD/RRn8JaKuLNU6ak/B
X2UuTNWi89IOXKnuAqRD2K/JoXBmhWfJ/dt1cWr2luFxOJ/x4UjYSi7abeG405ljKayZtihbnOpg
y0DUG2sy3N0+UWeOcButDBdAXGdjSIEKwTJ48GqTYlp63e8l2E1vq/grgzH3ZkRqO8eQRFZrth76
Df+AlPzCfdDXVQ2OkFj+Weh8DmawQIX4D0kY3MZQWiGMLyrTnSxeJsjFJHu7N/TZtpC8NoCyWZrJ
0Qc97mNegrzDkG5REkvelI4PzlFqWnK+EeEwGL+Tm+sLPXf/mFVe7MDJlTJCpCwQC+iJm8qAgf0h
sMZKIBV9fgbdMD9ciuAwPdtRpQR+CePQHcpC0aq8Rz495CZ1oiiwxgF/rcSsWFWBi41a3G3RKy/z
nTnF9rMpdSmCLEWn5g1F2CdR+lg5rqSKvJgAh9Da9sa9iDzEU96zidvu2ldScpA82Fn8N3oITpwX
Su9C2hvt/qCHvmqt2QzDcmDuG7HqSRMCrU2OYFSErPreQJST9s6easH0XwOme2cX0fyqfMBV+UaN
da66wiNd8X1YK248KQOCdfrY3BEiprd4oWcUXmfuLDdEgMwuX1PYgehYRJwbaggnQqt5aADrXSWE
zSkcXut1y5xEmrc4psYmWx0JFWEp6du2vQNiCpEVejVeKrIy5A+jG3S+OKBR3esck3T7rxGUcp2G
QYFTWlWkcKbdGQBQqW8XXayzy5fQdCqO+ni0XZuTwBqWQwmptuCyy4HXgXdtrQLj7cg//qJanDfn
mplTOT1fgJlFvAogXRQDOA6zlMzRef/1mDGFwBLVNBVwcZuYivuqcJfJvxuN/clOkIluX9aeCeA6
LEyGBixVhGvFr4bjZnFwSMAJW/TmyRxvBHZNeCWtfk+pkReEIeatYgKLUoSyrETEMdOQJoBePiFx
5R/Ksfoky823f8iK9ccuP1pRRcn/xPdqfYUOtUv2SIzAiKKvhg4U5BfRMGApDAaKr/gYw8ZWMgqB
oskBtvWjDNaJTeLsxYlBJN3nbfdO/GSsKz1ZL8fM87rrlglyHMq5Wj5adv1WyuVe5hqq1t2xdZh+
e0uBQvJFu9zexyY3mkHkLSNvxh3m3f1EGYC8XBgfLNGMvNL3BoNj6FAgkqkCtf9V0kGVnA+EY4eG
Fyl7JOgyABj5ahW6/1WM8Q4haqNFdeUQAILoSeuVBaqaNY49jTphJqzhImNr2WF5lAOwyMMvFTvH
tYJkj7j/k4X55n9c9flpLm09x+EK5RHtKlSLFSHRO1oLjZPWcXHfHGT3jEH7ap0kQBirO6uRbdME
N5Ojs68pEHNA7x9XZwHFPDQOLa1Am87I6N6wdUeMr2YtHrxvn6UQUGFk5b15tOJewTT4YMKPDqxs
MvHvr7XWfforxXtGUO40CFaD7NBzpiJVWmfyyLYlAuoYMaiyNdu4muL2KUvKy8Aih1bDgnQ8D3Rz
NL/kGlQBMFupmvpn1nsXDisSkrI/8ZrVTmMsNMt7VU5pqTDSUeoiZq4yyeyzxhSLSWFroQAcUiiu
YZKv9tCkOp1Eu87RDkjk1DUp9vKUC8Q3YlEl70S+Zz4hqdgl6IoOk1+izL10dBECf++EGbEDwdGG
+F4JBTRfSZ+ddP6Ae26De1izAwqrZW5ux/bGP46UN8ovRRCHw5c4S/a0Emhu89DIEef5pQr9s4rJ
SgjcPZgRcYVEY+T5LFZ69LFLpG9Zja2ROekjKizmgUcMG5wqX11x0xDxUEtEJtutcH9WCw2G/vtm
bSNDKOojZKPOXVgLldfP0gnnbTbsNT0jW6PvCjbIkEcLo8WTbksCAKiQ0AXNg8vomiJl+to5opA5
93a5/PCrmDNPpKnhDrnnI11KePz9/odSSkUXT0WxXOnfG0cVtYgGqWmSWA5xLKCKN9+RO0xyG3RC
JxllmHHI5FLqndrxCwoAVLACfEAMD3UosBbieECBfqbTBxmW0dfwE8meLIRtui60ZEcjUROiYu2z
peIXv/SUv7RVfoKr2AmfqlnVtxMujb9okJegk9mg3Ds+WqmuHcqUqfs2h79XR3de+XVtm1Ngeok0
VGLfBI/gKn2DXL3w6VakpQQP4N4Zga6frNrkV+cr1uoqKAairp4GnntuB7/HZIdzU0aniP9/fnkD
deMPJhoMerJNYyZY4/d2JT/Ws4WJGzDVZyM8poVZqnYNI2MsnGLnSMCZVghcPnUWzxapiEJ0upTi
5h+NPc/YvXaTBMBcCGCUZVEPeSpK6rEf3/ElgBfwJvIOaWCXBrKJUiYtNMaOZ7OMcp9eZmnlRTLF
arRSS0eOhJ/e/8n/dNPOKtsAxClOKbxGDI+e+MieIP80jgrd5rG/va5k06AHiIscXE5fi5ZrEyFw
OGKoGBcYp14ij+DgK6sO8oWtBKVP3xxZHYtGthrESzE09Ls3ziNGnyrjbsRAd+zJdlqFN3zyaLsk
Qw7rwXuvqY19lcvgrGDeaADcxjOBa6kFUtOjnPvW3nIuUuMNlMLS8WVW4vWkohkMvHSQ0c1nmPGF
eTgFzSkLoT8ovlXPB6TvDHEqsCCvCqUz0wc1mLMbz5XAW2NfcUO31Ena6oomHMYnFXS9igftazkv
rkhYVD2/tiKnMyTelnNqyDY56/ut+J63K0zJBbFWkDriI+ZoM2bt4ewt5mFLzVRSfYd6/xP5Lbzs
hZheVuTTV3fonGki78Pu9lAiWyhnKnMJUuyo2z4rzhdhlPWbuqT43ue+jAjLmwCYOwCscDGGUlyO
TQEvMZp4d0YnycTZGZ/EUfwd1+VkAcs/PlUGjdggSSK9J7skwUGBYvMqnmT2seMriJpblpQk1SQe
PVLr9CEOgXhbk1fA5M4z2SDLhmHtTnYM4CVtO3wdF0k2Wl/YFKJe0V6YsImqxP8N4Ep3Gvq3NRNr
OTPHKajTZ+MVPfem6YcAPGBEZwxcC7iEaBtND6VU8I2Y8IGn+WYAIhZU5pNzOJGKGwxZrgpQur8i
jerbSQkmj9h+/HkA7qsSPaC8LanCUrxJU4NOBlqYgfH4U+UskEoaPq4umFNNx8UE6Jxjs2eu7am4
/sB4sY6Nc26zOOlrdrvK2egARCOaiDCKQ9JFsQaVnpDadQXhTrhP78rTSeKr69dLiw1F95iYoYDR
gzd8pfOgFrHUY4f+ZX57ujbiANcRB5Fxb2FQ9BUseXMWLoSxETeSebXH7xI+sbtJClJj14srvKWB
4as3RIzpk5ilfLJQ+MWS13fmWAC8f5lbCJsWh5sQwp6dSepGgazwiQX+AnMq/hvN10tqjy1Pdsmk
GZzZxlvG0jGN9pZcfWdhAPR1niQhDKa3qcvjCGyvDWWiw7yBCrC5EhHjdB237rcJnpaLrGSMReB6
R+Ita2XVZMRgCcD/1uToxlpKfvyYmNb+xVXx0G3Mi/F77z6/5rqiP/cy7D/Ize238mtNTz5XBafT
bSIPhAywysqVXo2UAsFU6/nJnS6cYzMk1CtCfPbSVvcoh6Hr5gW0qDeq1Gs65vcu6JremkhMKke6
ismtTQJWuMoDu0fkuvRQgJA8wpWcZlKj4QV05ygwQecUJHu2uCO6O1f5jAn/9LTilWBYDbg+oN97
fHKwH8U2Q3yzUCwGV1O+yHpL7OgLsCmaJD+hZ0vz4jCPCk2EePOJkji2VuzKgo3xtGJv1qcpo4SA
suK8mMzAbBu9nLsGOc1NUDxg9lRlvcYCB7HUj/ovlFrvXHIWTqncwAs5SYhhv62kGAKmZZw6qa0a
CYfK4o+wIlfpcNs0Cgh1RFM0uoWaQTBdp0ioc33XCQnlN8JwGMjNRxkVbdmxq23/+nXxxQa6+gWb
NEufyb81tPbUTNSteY8eDjqhIKWAlltdG2P7T5CnJVVxtuHaBxqWfBY19gHNH9o3Wc0lsbbq2RrA
TXn21e78EmI97ZHUj/92AxYa83y8GSd62IhGcktV+m3L9Q3FXG3c+WZ5RK9lBmpXy3JyinhcHJSw
sGehM7jbz96RkrR858aG/nBirmI5Cdhm9vsoFQ5yA2V6zf7Y3Vf2xr7rULtvV/laEaHSKAndaQrl
q8UybbCNvgY8ydLYoiMNIkWRnqwrkI6v5g2KwAu5es70HD5IUjqNAjnmzWY2zPkIMVoaQ3VQoftj
M5XmzWhZfsYCWra4roie6JfIEScdngt5HbmNkAXnuvqizs8jNP1lyvgnfdsaJUPFRTh9mjue0cAq
QCxvjVsgoA3B6GFF9d4/YljYmOx+29Zb8MSp4CXxTHFybQC1hNTw+phnX8iqkldUk9ngfebUBG8e
Gzz9JFaRsjZp520zcNqM2vbZBfkh32UfTY3Ht8fnlhV+d1p40dKHPKwhXGyiMSL9FRUQUl82HMJS
ucFkFj7Njwrt+tdqX9I7kvmDwaAwtpPTgi9ff0OMKhaZgK2AwuO15PxVzl/jGb06nmvvWBnxeRHn
sTW3Z2Ga0oscLkimSezYJrLtWy5fjUVhBmS6KuHarav6Zf4zzNQbSCZsVkZouSSoPpm/M16A/Lqy
XegiVnaBDyFA7mo+MnkX8gop/a/cQTVZvL1egA1jBDCo0lQ9xVAGgoSo5KPgVnPBhM+GVzI2DSlU
oCGDkZPoHkvoTQRJNLIuZIHCQDGEm8Bcx6cYpoIfWFmRuIrUIxvMG0+Q9LJDnyb4TFh/n0N3JyVT
xt1d2Erljuk331ENt924yvVqjMCiyEyQjNE6poXM8I/DwD2fIfdYoJ/4GJCYuSPNrJBxaRvyKNCZ
wt9x3Dt3ThXUN4GFS/wXUNFK9LwT3jwku6Zk7/vSVDSDKQbSdacdo5LdYtz2S3bJyr0YwSkQQYms
sNgjBXSKe9257iRPV85bulhlZcGo/eLzj2PRy6YWZYXpysTQK4hP9PMiM7H1nVIKc66qgpueop3K
7OTnq6KWmdH9iFu//+vqhhRFViv+kKVfn0BnupwEtJX218UVPdaBofyXtIZ3PCioHhH/TkTX2p1+
JdMCRMOzj2GrysAeERJJf/ce6J7vXaIlSkMcjsz4XcUEC+4rxYDy69zwz/yifwMAdWOwKiqkJSsv
KnzxWySHocIX6bOhCwxU7JsEvdO+nkdqGffqoYZt2RBHF3ddqnyHmRB0UOz4FcT/poEy3h+gI4Bv
Z9sHTas0dgHbiYM2iVof7kprQBjNnKMzqmBVZjEzAzXKLUT7fhTy5lWR0+k1Wik3ouckdkw2yFhL
Prx8KmN25Z12vVWMtWZwpaLLOBAMC9CGHIbEmj2b0VGhBYOYCDWitstcQo78WaW+YGWAchg+cLVk
swPg/Y0zDO/UfMjtGFxKqp8hqF9ccslJw8o6/AV36Kuj1OhzFXluKh/PhBtCQ41RcjmYwDzSVdOB
sWXA7/Zwvc45ZsE6COgL2Ty2LuXLoyiLZOMFAVKiCfHeGOKpa22IWNbSeRnRt+j9xE7bQgR4U9/W
jDroQL7mjBie+g1ymuM6EZhkMb5E+gicSqfomV+EESHKXAIPZvJIqQyNtc4yag6N7syiy59VKs02
hEoTCeIraKeDsWcVlY1kVltLge+R5InSOq7d9PTj27h7l/JT3OCx2UtSD2yfd8Jp6sXf6UNoHpB7
Jbdf96idSOMANXFdS4vafBQbOfPrvndoP1XIPLzFnqWxIvSJ0VKhGxB9Xwh7wKrxfwX+1TuO8HKW
crWvZ+aU2RVfu6/Q1xJek0VkZtCW7QBRr1kZyNlsRigUKPoMnsV7Ynz6/Al7iX2i/x/nIQOkICGw
E7QvrF6tEW1DXzwfRS5vSpZ3N30xw8QL0SbMRguRdM18dai02AJ4PUhPoSyUPzdTbdjaw9IDDN6s
ffmDHLehdkE9l516m9dNmxEfSxaWFeLALbr8gSszG70X941leiXRoZNQ+XEySKB/1UuFQRh34pPr
UOHpLuHJKawpyXOZM8Vbkhq5jFuEklEDYmNNQXqVGSw4lJgjRqTKi3qprBjacSM9IeDdDHO5lZ2M
kY3HYl7wnxvDMBw1DUymewkKcdjs9IGnm2QjNXSUO0C7L7CV9JSDHsu8FaQOQ9Bdum4biI6lXLfc
yrkrwfd77huUPyDH/Or/43vGbrhsUs/hqfhREQuOXpQKKB1NXlLd1ZpJwTlqOMF6xP8u29ehlhwl
q8axzMo3h9PtPtalvhSxzDFGLD5YmYWwFuytdL2+aFSZf7RY2gwGoOiUOSo7hyGFlZ6Vp3rKMpN2
9fWhSH1V7jp5WPQU676Y5BjHBujQ6WSloM306TrOqiF4cVwLxfys5MUhYzHYz8IlxAmQc4elBd7g
kIUe2eBbxFBmF+GyT7DXech4qsKz01iSzHT9XSwRaOVeMRhv9/P8cnyvkQRn/RQvfjhFqbMs6bEI
iYkXYtULMyENNzMjJSPL6q0xjqJf5b3h5CpOw7Juz0RAvpna/K4P8Vl0nrJS15SQ+9A6Q98Pc6Fr
hNI0XGVnibn9J2zbqMmIBXYXllzfchrL0j5H32u8rWhwN8cYnBDc9Z+MOWAiYxCw8TuqCQaYwHzt
T8U78qHuWRgVR/sn4TYfWrG/Wsf1NPCDyMSLOIIgK7HG/V1gJsK+qSTHky5qyB/EPAJ0+0I4mESK
m/jstXazEB3BtQJK9p5RlTlG5irPauJSbF+ebpWILkD0wFELKYUYUCk9J3d3cU/OFKBLnriRty25
gU0wsaTnGgVOVBitDwc+KX8NHyJs/fjZmOb9I1hFVu9b5j+DAFocOc6H0jVrWVqT3k6sXvO9laFn
6pAxFDynS4QUAcA+gsCt2HGtQMrw4Y6l2ITqiZLRgBDPlxohBG9hJ6tiiW6KflHe5t0kOOhu8cwH
T/nhunT5tyeZVZJvZ2M3DodpRUcCKFjzh8s8bOttLjqElV7/t0GZfAK1Q2hmc7b4Czx2n+mAgIxq
hx68C6pGoEQx5Egse4gFhx21x+4yZF3jTTo+BFIms/k+wcyWdIX0K6d56z02gBa+60XpQHlAt1lq
YzY+8v2V60VMIH9o7UIqfpu67WXEOaWMDgJHpzXnmOg5hTW/UzwPEPKsjDypVkG6T7ApJuCvJn4D
hPhXb+r/5jTpEtE/1BzXRh7WLaigJdKWM0MVOJEiMzoUEZWMTJ/oWjG5SWqxmdnMjTMmGyH2b0Om
47n7LN5bUS5LHdLn61kC6PZMRSVnSKwm9f4WWeBM0SdsdrMY7YFuwypAafYuiAQLWgjtGXF9ZDii
Km2+3mB22mHWLJhbgQElF+A7saj6ER/3uKtPYtFbwYovwV25oY3nV0g6kacYlKTNNT7hKbomLQS8
VPBhv4MgJQGxjrTinXALBebshKrFqOSa+bBMgY+4IsNJ8DNncANnPOOgBe5dSuzcVrqT+W/O/DGi
27n1L6dmvslBZljSdG2qY6v9p2EfjrC9q0DKKyDIhdujCVB4VW4D+2XddqagCGBRrqV7m1aAnqSX
SI67N8Y6YuzcuKJqhYXY+sS88gBr/fwWjHUThGEiejMTCgtrcBjh7bnUqy0y2yYO60scz2FbjXAf
Uh8T5GH0aIFfRSB8E057wfELqsSLBM0QlcBbk2P4LMj+pFi2d52fL+W5U5ceYnz4Qd7Fnoz+Z69v
g6MBhAh6HREcgO/MkluqFJbphgUz2ujOnETXLJaaxQvoWwV7ZSc37Yf77bipIjSX/UZLCUEnHybE
cOhrHHQATM2V6rUBlE1uVmPdJsak/QN+1FOfaDUgm5V8vB4jv6DAG850rDQwdbYDXw1w8hL5Dvxs
x89uHreEVI4QbXIJpYH8E1tnOHbxnwL1WIRVhFIY7mDWf63Bjx6uO9QLm4eiqZkbFPUo1y3O03pJ
L55Vv1AxKEB2ILUVNVnc33SoEwJnBfc3+NEaxsuN4Khe0YcGbPJQTAxd1+DJ6pvrYO4uDOFzg70K
wisKLaGfsE599BmWherrGjw4EWZXGnsqSBcvFTAAIFs6yggEY5bUFnlNWUEyOK3yJGU16htjmClG
5nZK1aRADI5MJNpezoeyH2prPUN0jnmrrnq5OuHRnfOdMIedqWuT8D5xBESLZ+KWEoTRN5dLS0fu
MK4eWuRxcVeZAIdhLuQ0gj3Z3I8COIGfC8bLA9f87WIhygQPFknmkwNaTQe53/H8x+Y5zmZIOHDN
58Q4nJqKIYEvZK0e87KBWYRPRSRCFyYNuZR2aDVwxlHpyWFGrTECs8X42cVC/+QoCW7WtIHcKjm7
CVTCNppPSSViGnwVR5Uz+XKwQXmpJEGKua+dZY39FiPQAT4cFSkxn1GILWcgo0e/ve4KHoFytNCr
RnBIDdwP6g5Vaccy31H3ROzGJCvuWUp2dOSCdZJqUS7/JH6Vsc224dC6luEnvWCwOeIpCuvPebmt
rfhi0bKQlfqYRQJydh3qojju5e9oxzfM4qF9Q5yefxO/VWjoZp6YhwsL8mGKXF1HCiTwjt3uiyVH
fA7Z4laM5Lm5Q0CqwBfQb71DkXrTgQtyA24TENDMTvZWlkiJen6nzzqTX7vrfN+l81s6jVQGlG/9
EoZd97ZALvSVT6/SRziDXuzpme4Nyw1BmQnGAqFG3pfFpZnEr48WXxUuWtbVA/XYeiL20yF0xiN9
k7BxuAPeDOKEfLv6OC0qdY6vbMw36OW8YgET1rbQDWxiW+m8xFP/3TNyQqVE1Hz0gAe3esNFGRCy
2p77jY/bynGewsgh63ryQVTNLM3o4HljMznJdygxqprjx/xNnSp2zauOHG73Muvgsqj+r/laL5A+
ffAV/QfPHk5AID63QoLkZu0QQQSilLUrIm0H6Rmsiwt1IwXi9q8zeJdclASdh/S2E4ZHnPEwMPOk
qK/hh51aeP2+0oXWII3Zdh8LwDY2t5njs7SgphwOVggP79gFaYjcw/07iCuTHf+V+qXWfyIcQZi1
S2CWRfZoa3NMc9BT3tgEgaVAtlZNoM5/rX2RmgL65vqKrF69yBhnubYHWRO7z68jZWld1QD0yeGp
XgfWVKLQgyCqXtsBxNqYzOUvslVAo2h3dkTvPfg98AgSBVApu5Bv5DxwjplPUSsHcBR46bMO0ymA
OfHTwBGjVTRl7ltQqzAMEN2E0l5L2YyI67CUxLzjZu8aFaISlxC883t8rP81tWo0ntpwZ778BVQC
+buyeF+sWBK1bgqbr9LiGwsJd/Zs4+yQXhiscnLYoK8LJFZWUSJxmnWkmnI6FK09Aj/9f9YW2bSF
bd/sv8fh4U4Fonix0pDKO7fwJK0QNjT2ZqD/BP8Ucb1USgkdyMqgaWbpiN3Q+z5uk67VIxyr0XSy
MpuFnEx/7kyrGM5BrdJFtYYviBis7NuteeDbl9QMdv88Oz1W5CgQjIpt/WCu9p0kiORnKZOxnot4
tvpG7U0/iCC/2MJEZ1jmFCpkXi4HZuI9xEy7HsMhNSDHYyC3anLtCuGJwaCg+3VmQpeYIDggJEll
0X8kegKuU3GRPpDTm8uDXGp+4JVlLVTj2+krUMKuppr7hZ8ThcVdbE2ep4XfAs7VVtH1HtY8GhMe
L8RZCHjCJ5vwVU/mP4XfWMiHbyUAztCsmcqWIRn4dRxCDD3FFGaTRG9LMTdY6VFr7XZE3PV+if/N
M8eSC7bJRmyTxgfJKUDyGyYYgTLYcQbgr+B1adAlUbX0RbA2AgKs5Ci8wn8/jOPVi8JfBG4j+qiP
BAxfpwLwke8T/cGzleCD89L7AFFVPE5RL+e857a6RW1OH/N3ZMdXbyTNnDdGYnXFF91SvWEmDb2d
eR2TGLOHU68b6O1UuBqui9hqlrschlwlg+/UZntWkBecaNUV62ER5Ye60bgOyKoWxiRSLK5Whz7b
7Jr6gxOjDxCwJZAUZbIXIakQj6F7GBrwc6Ptrf1qP459YkpN1stZmkqbzkJVUOB/6H/+o7DK7hwR
Stc1nV6X5xnV8a6aaE6otrS+wj/PiD4TpGY/8juGivs1PfQXclArJyGtCpkAJXT+4aUBChMnZ7eG
9fX/tpRHLwhMEDKV+lsLNkQMs6oCoi0sLEitn6ibpdA2LdtQEEB9OzrRjh+unCXms4eMTSupatx1
zWso418E/p1iHS4oLm59lgmqff9GH682m3bkxyYuwKk+ruIv6asqkkpUQAkEQw7K55Ky0dqtspz4
MDAD9cBTigT5+XaZqdudjQOQWmRVWWp+pgGx4CwnzrjchBdlAvdrtDJ5UgsjoDIn/rAQCp+02mMR
dV1veucmmiVJi1G+x3aSXFD8N8jGIt3tbdrODkyVaLnrqkU+1b2FNAszxPNirj9AA5FzMN4GOEEF
vH5lgGEhPpLdHBKg+Qf8x3G7jxiABCAGGUIVqlbFPpOzNz6MTRr5V9/hAVKlrn0wBKVVF1mdExsZ
NuN3cxp5DbrRUF3XhMPN7+ZWXzTymv7X+60uqFp+UHhLsf3i48TQMOgYBQsVk+gOWKhzlzfDNtew
bafPin19TTXnj+B5OG2JnFNCUlsDCugHGYEolMDFjKvVGogRllSv8tlvd2Bj4VfXB8YhfMNhYkIj
Bkc8nBiOSbitF/LpwtXtf+ODL5kZjlmXgZPZ1lPYZCVMp9yorQUJv6tzJ+F8XIrUMbThrTZkidPs
na8KbrgQxJGfbfiXZX1qrgZDOjvLUYdRavR1Y9BGm/ZrjdGnveO7454jTf0F4rmDQdfpDxICOMjs
kdkr/yWkoGhW4kEjg+TbE1ZSk4IveOZVp+bRgsmUvJ3aH0AWFP7wT2v4BV6kjhq75du7PbX4tJq9
IRIzCKP0Pm8t+uBVZHXKcWEpvD7ZnO7GKC/ej+4z17tGzL4xhkiwaSw1aH9v4oMXY5o2bbD4Oele
h5ooUXIHnCnsTvroMXMGV6rzK+WL/lFatJN4YBJgJeSJxVIQTxGsRJUxpwy3bk7XWPP+ChslkTSz
lnFBtUr/lRxIERvzRRK+YjWFW2Hlqu1L7/SVwPWCLb6AtgWXbp3KYiqrrbxepC3TDcMrzMi3B00H
hCGb0IogDGBndC56kOgzIh8jm+ONjWagpysOg3a25rzAfSh7ms/km/gQBPz2r+mUxxkl5iy0fRAs
IOMfEq2iMMmTS1xsN36esWlHw32qF5WoBSKcw3hapWMiWo4gf8qw45MR3lvCiwRIozOXWDDaFis4
c/g6S2Iv/6sgbXOSTa0TKtHq0Qoxguw2qkuuJAIsZN+02J5wA6xBHqdOawnkt1cFcdWh2oOa0iXC
9UF3chVFQLwDpHxdseYtcLM2KKSqCDBOnM48GkKsYGibQCO6iuyPjh6sd3/n41JeacEqNhPU1xGA
I18vAH55MuF25Gybx7PlMkUhRGLGNxNLT7eQRS4+T92gkkQ3Fwg6VpTilOsJV/ZHY5CVRiXYS+u1
RXdtoR+2YM7A/lZgNmQD0gz3rh/tgBpXdWFJflAzjYgRgDajSkgYKVZhkxLpr7r4rlFdOuNqZKVQ
lp+GeYXQyCnxl2K/2AztOndBb5R5BqKF6GioFTlaST+i1dXW+Q1kveEgjlGwLzbEgRHboItMx6mQ
HqRE+km/E537icKmNGR9lKFtZYGcgj1Uqm3EDyOAPuZ84a7fNzOj34A2oiJeHdCMqtqhH2NqbSZK
mnJgxAqe5KvFsfzqbcf/Ah6Ot/MU1ilC+j2ce4+7h8g4vfVeO0bQsLVraUX2JaFvSDvVnqVoD76N
kli1HJEOwLCpBb7hUDpasKjaZFsORO1QnCkYFSOqM2aa30+HAVFiFeDaUITUFam8OJTZ1fad7HiF
1QomWPnHVVqV9nWf/CmFKiMrWEdrYPGwM0BkqICUAoqM9vsDhJsFgUzpzjoNYSliUDKOfpNu03pR
/i9r+GbSTHxIqDU43iQ2jEYbStlZZy9czmMFIFZsKn37KkmBOvooYRNYhZmfN3adNnYRBU4I1YHT
PX2vlkTtEmpB2jWq6js411t834JV810KUfpUIhAAXgRR9uvKPjlHQ/G2DiESe5bP3Nghu/toE1i1
FQ35YHEV4FAq3xgMz5J+Jz199UVYJQMtdEr84JHWgHya2JaZtG3NGXjCcwLyrKqzRwxoIqsHvUWf
nUh3WO3eod6JpkHfW53pXbXR8px7MBPZkichoPyKC9yhWcYnmTxNMuMuXM+LeaEhZLd4jcP4Tnwe
OdUS8XzPHFo80pkuKN3FtFo7T2vRPjhbFI0kBODylmKVGfDwW3uf43MWpsjWNocGWc3APueqZlAA
FUB8jrVELvvgG1tIn/NV7qyH/+GiQ7ozLHjExwJyAfCHn6ashUFOtzt2jrf8xOI74MAjCT9OqUEl
idH12tT2GZX08+kTUHo9LyVPxyBDO5VZaJevNNfijl9wcT65mIP6CAj91XFtiIjTyBCb3xlVlxdH
PpS7lm1lMUsVqR3be0rdfa/vDgOEtjFvCveCGCRhLzp3kHRylei5Iis1Y6QM524HssG6oaLzSr3x
2FzFWoTTZcW0/5369nnAU0Edo42u99GjXMQQI+23bf3wpsBoE6s92zscCyD+nCvYEf4YKXT51CgE
5Cjyez40TGu/3vKHE9jaBNyfotMI8h/7Y7/RzNDUmTlHpc6EnX0vx1Xvmq0CjxCYSiUk3yVMROiq
YZ7LMIBEOPSbPV/mEOSwccGf84njhdWsRo1SDsTVksPZbdDIiizHkejoQxged4nwI2XvzONitiQ2
6uIiHPOUdHWVXYFpgmR01G7iKUGSOg2uN6XO1qkupecC/c7vxzN2H8NLrM27M7JBcLtbG0UVqsrt
V2Q5s3aLUewwxGd9Ov87Vdf/BaRj/xyDq/+p34TSkmxfHZ1ojPkhSjpIxp7LCH6H70zYjIfi1hDM
eX5xDfeuO+VfUrLOzwbg4f2IRLmGAOP89S4ZBOrlnO5t0FDqNIPk9Rwmwf74cM912bApT72CJp7o
Jw0F/vlZLnPW+yu2lHzQKfrkhv2Iai7Df8Kvi6UnNUV7AqWY0Q8tVWJpztubDjYZ7L20NoeAp+ET
7cqO2+sytvAqo8o9tohk7DKdrwKsNqk9+Lih5yK406IryV6S6pA1FD36A3A0sIrKlRL3/YnyYnUi
qHUvkxDnrcPEuhBfeotlhznVjw6eeqc3qU/ocPc87zxu7VzOOvcCInHPi1q4Pv4/9/fOpynZHXIf
eon1JrpC5avQ0pdTnSAqAe7+QIuPIr3kyJhANKenCKAbU1DmOXvDjSzVPyowunKZ70whY9NNt9AG
Gv5hJqcspTPRMIA5uawwPEdaOgxZkfOQG+pLhNU33w68r6yd6j8WToM3KxtDspCnccnbRjGvrv0H
2dkJgwnoxe/SXLG+cM3AGFcpxATrxymT+OPrVYQW3cJNLNo1BCuvKNUgd20pYNGUomfftVYvetd5
2qwlMHXPojWpaK2lokQjpGigAjfjpyaR8I9GJhZhl4WNH3x6JHhnGQOnx4UEy+ibgwxTf8rD9euY
cDG+38+WLJSUYvzODVczqIUEf53isDdr4zrhTWhOLnBSEvTwG8LEQ9mCrqanXKFEiv83o7XZUsbA
8HRD925VvdWyJTQGErueFYnIjmoDIVMmRYvpVUhFB6IqVgKPHjzk4emjmxOvqjXZsYrGCYbb+Yde
j1BIA1ZuAuIv2fgH2gcVQZ9/0KxzXD2PNHlxLecdNi7/J5WfMmYHlsEl3ZFJ1qt5RrlNq+aONqyN
GMswYuiNBYsBXXtyzEttHJHCJTvFog6vqm8ypMYNUokcQfMFoURB5f/mg2G3ZsDaD5CFlleszjco
+nHGGDDoUUU3ewaVpYYi40JFJ7KFNTudS15T3Mu9KlQxm+H8xVLvoVA+/XVW+yTFiRhbyrqpRfeS
Kpm2vMtTw0uGwQZ5AAORuMS4o5O+DPf1C2h3QtIKBRAJymXQ6gy3Z9sefVgaZh1bAVbvjjsRSo/f
mmDLqwgS21HU2CQMqmRwmAt+Qp7QYoFgLjlCUpTlTwkrfnGRBwK6IcpzHNFy7uSoxYFVq+CCMNlo
4yEaLgRAf5rY0Ta+LG9TQwGAE7apTbCFED2eFNljiLugnxY5Zh/7LN+jXzo4NLoe2Suow8iojbcU
LU53Tel++Fjt+w7w8ulmqJdzF4foxiYrZBsSi+NeK/eUv6t69j9EzeMI0ylCp9X/dBKNErCGEnIW
c/JdQFy63DDtS4p7qCASO0FC4spu4nGjfYWVB/12A+uo4yYxrxUQ5RO1+PsCPz/j+BASPJVeJx7t
9xI9kk0S4ii8yMR0RPsPohc4+C+tthaq8g0b5YiXfjWPXWtiF9zEV+msbjyKSIAmz49jRPoo39lg
LforvixMCCFGpDF/+PhWjzt5ziTtB3goKllzY5FiothNxFci0xnTM/sDUpyqU/tvGe2QFCiZV+ma
/j27vCNwIzDKoiPWBzD+etoG0hKJxYAtV+cuEOTU0U0q3FdauSiGyYbcj9oFXHs51DNMeTljeWdo
3bMJEn8q9sPdVkTGSE7sEFgMqNku3nyBv8siQE1oziuWg6QHYWUFJr+XXLFinSmKGg/p3L3i6REm
UrcWiVlpV0D1ktaemaWzp/nAL+DyORHklFP9ia2vntGjy2hxyLoMH2AbBIlJANIvPanP3xXIIA0h
V7W1S3zQOilRZL17t5s5oZIDjaxhmpnuZlHt2U990mJnX/oxVoZ+ZkPl1X5VEvQx/xUo1LEczvfj
OFORjAqy+69SqTu5+2MjHh5zz0gLxHFB5GkTZhMIrbtmRkyUoc+HUJ0K2nxgmHxxFpGkvsD/b/Rb
Gyrb/zfluFKtwBGPckKwH8NL/dV3P/2+XxJQTGIq2TaPunEix+I9BqLgYDHmmntztifNDDGYYO1e
ZaEyjRvaWp5CofOm8fyY/OYbzQ2L18YX5xK7Q+sjJ1ELlYgaWkeqsm+GQ4aQ4H9kf30coY/DuQz8
aM2LcBT6f02vBLK90/1+tLcF25YeOYBBaM3XXZ2GOkO13C2LWkOE11yTQAGIKm+SRhbn5UarfCdr
JcVMSz/jUoKXyDjrQzuRqEbgIUh1Ujd0KCktIFs7Ree20xvJEL3aQEoke/lOtyvQ5EyjZp92Lo9K
MfMbqyWJjiwZ991JwD0WQHM+lLltZulDXE7BEz/0UUzy25pA1w5AreyJCpht2KNoLSUScs69lPJr
/yTURvNn1SIbyGFbP4ri1HMtxicmlzl3tWub+XFFnHK5QIMu6cbWXsPNPQm0FENwPHhwoLXw172y
XWpEdQ+EV8roCxGmUL83+5jTyRsrE2jngc1oywWZEoksrBCRGffjvuY+1qni3kFpK2JtTDtmVTzJ
FOKdzxSbfJLr0cYdU0IF1laYgBk4au6nFvNSCR3xNhOMWD4ReYrc4eETmd/a6xuWHyy0lxaT6WrY
qDBRC2dr7x7wc169C9IQvwWuNse6b3fQUzlocZ9aRQa/T22lHxYmlb+rQ5T+0zKoKW6jDuLgyvgC
p8ZdkA7QkR8CeTgS0Lc08/YgVe4PVm/BVVvxPEX/i7IyslDKN7MCDhfHC4W+g/BWRfxfQkOPWVUh
/rOAiwdAGl8ChwEzYtY2YQ4iXvb6XNWDDO0pX01AEbs4jFvjwIYj9mifGGkfQstkgDJ07t7GRMpB
gUv6HXARpIYuGFJPA4lZpuSLO7UAk+gbSz2OjNuM/jVGsrz9IPK0Kps2v5pBPo48iKfbHYs9Y0r/
nwfkf1IL2hWOtLhr08k9FvbEyjKGlwLGkwRbsnX34oSGZfy0J1TaZ7L9EnKM6+orqRhpKTiWploD
v42u7e3XsZiDd1uTkvN7Lb8kmTkgDC6ZP5EVUrl5ZScJY0IwAsJPw6jxEQYKqc0U3uLwyW1X+Ncr
WCrqJlVm5/NdcqtUrRK5ShMEkGCci2mJfp2psIjALCe0bstq9qFGrkURTfwzpVhBqwrrOysusrOr
iAU8SwePD0m2HWNzzEWnkD+eTBOygDf624th+ue2V5G+GiSOjux7jQCfMFm1EEtm1vDhSUxW2kUQ
L5YpcldzUGVb2SImZ7I97cDFJPR4fkuoVMOfqzsIogazRvRRpCwvDY4xmFd1CL8JYd+joXgdF9c9
o4Zc5wvB+f44tuUcMYV8BGby+XMOXC0Ryj2LTGNXBSgTPI6jWhJ3iQCcgYME5omEeSqFS5YSdCnn
BbtO6/VBXDJUR6KtOOvMj3lu7R7lZNz8mBLb16J7HQbt/FI/BmqU/OoD4P7fBsejj5/B6+2F1FQm
/BZctQ1wSsCSOT4KAd5Tn8KkOqRcssGXPpDRuWyl7XcxuzLh8p9WBwu9CVAEik7849O2DIAFDiTY
q8oIC4BfjnGRi9NQfBHFgzBg83SgrNVj+YvcJ6V465CcvbGrY94fUfQrFHB9wX2cTP2fIR+XG8yF
ZHtUxChcIQLWdxuRMIn3XPe5Y48gsqnJ5Gr6lBD/yLW6CjhUrgZcOJv13eAO/0FRjg2pLKyuQYpN
CFzpeCRK3lPO/VtCndsiAh7Y35I4uKNfDhUwIsKsJmngTdr4gGankknf+1l9iFsyr6R126D3swPd
XLWexY4ED2Lclj5ISW6swlysfa268kroJaw6/6zzwI0maLLXRvi5BHrk0EuKoHUMD24VOCfei9mP
+KVa4yXodqmTxapUEgVlOlHs3CASACcwu59GaSXFca+6IwtETm/m8Wiiy6Q2usxQppYqoLMRtLcw
zlbodqCGgDAtePQlQzT93HA2CkKt9uVQJK7V4KumsJMML2Bx0vwX4qrFGqTI7H7fzYLZuXToRwdD
2wDEkpBSF4JgVtE3W/RthQff6dL2N6g3T9oml+sdfg/Y8PEtH8WRiVLuG4XPXx8aZ8SsObdrBKkJ
nZbHR7Uv1Op0I3LkzAlNzaPWeMXdquzybbBrCJ9iRppPVtOUB6dZgXJGhlI6ApcSDsfavMvEHV1S
sql9672lFm7w//juUfDPiCpPWIvKoe/ccwHbO7DuoHUtrt7ViWzZ2ayIa0YeyEfPxLI8mkpwmMPH
dRGJdFxeWoLPYlxZcj4Qq8lnU0ghk8eXafO4YnWt+ax83XQwJW/xTLT16ZfDLyT3BdI7Anj1S/OY
rf1sMewu1U9OekCAzNRqZTv62talhew+HnylSwhCAKTFutCGFVc/0l/LZBQ1045Spwxa9laKJTH4
KAqVBcDy6NU8cWnxfBGCoYMl+AvbDjAhDhRmCuXQo0qyUyW0xG69u9jeT4j4iZAVWNCgUBLVCXFT
M0KBdnzom+nH7+BIJ6Y+gRboc2N1U69hsdAO0thiv2/xOhXtAF8EM88u8hcMFMQ9aVVRyfsnFcIY
/Q+3M7K0H3WMHkQDE8hczq2pis4wDafCuf2L1tY/u+2YjJbeUigYZ84bmScQnCYfW41mr8bNeRld
GeEtny0oCpQed/NjHGLh9v+PxhIkvi3TmgD4Dvq0r0pqpPFo0hN8E+Y3VsTOrBsqFo464pN+4AAb
T0GEhTacQVopSqyWpRkRhgtrJz6A8UqvxfHpahQVd+24dRwcrb31YDF/zrWxmJvtl8I7gas6YADs
mmD++U+7xVdwNQzNapLNmMQYoPHGYEOgVf+wRLp6A87je/+UcSAYwETwYW/djBTe/OuNDK7bw6NL
xCImbmHmQnfZYOc5C1zbcBJiBADztNt0ZO3kNEuPBDnYjz7S1miFu3ltHzTLIjYtD3bDet9Tz9xU
i6JSsr+y0u01IbIgDLt2sS41XdofnSJLMDdHeK+RxS7WeLRS3Cflv7tUERx0JF9rvKLpMmGG/p9A
WmnxqISs+PeHxyO4zeWFoItXzGG0bU2XVY0Hm7H2SJzl707+vu2zqNUzcg7SgJnS7qNEwXebweEz
aRvWmWNuUu/jx0Jrx50i80xDCs8AvKjo36hKp4Yb/5HJO1v6S8MXpQzTWGV8k+SyZWLCfdBASTS8
KvZ8Llcvj47Y345e59Sm7PUJD8P3B/IfuaaTcR+JtP+3wH4utD0r3+12xm/LPCsoEUpH+NIxaPVC
Vl5BU5mKLc7OCJMCusbo2WKfF7RDBsEORi483/qTD5BXHKEKG7BQW66qL8AjUx71ARrAexAAm6df
jV3WkWWSzcKk1euEuAs3xOPXSbRUzZWgVupcVlWKlAGwT/F/+DCpfOvjsaUCIbbra0iY+oSB1cJ6
HPj0kTnnUw+hb50M5w2/QX01WmkOU5gSCCY7bdbUUYbmDKvans1+DkIFOYRdvPWyYiYn5zxwe29E
36tO/43OMryiaIJn1g3YmMKsmfUZ3ilkE4UU2+zakLeGOiRiOvxGpJu/8bkp0I37xR8079SBl71s
qEnYX7PY8meRpc+1iZI/TWaT8B6GxiUDtdUtVPugxuuDAoJRHPsYLpUh18jvfu3ocqDPeKFj6LJB
y1ppwr1QFH6YsYTM0xsZ4X5DJyPwZCuk+p+vAqlJBR3smRmlZe7JGgpyZoJWfvWxMT3RZYgr6OxW
Yiz/ui67c2wRqwGSXREQn+P08tOc5iEOhcJKZ/6+DZXqmedpmEY77E07LHHnDGJM2YnqK20MM3C5
RIDnBSbkqVK3mFh0nlwAwopRamvMB9tGzwU4nTqa0AjUZEIgbQIGoFOq2nsm9KgmENGfFwC+gVRo
LTOryaVnPmWd1UxGayqAlgKEJxNAALutjEEYZS2XMkMjx2JvRidLJnj6XTHiIcZ+OWA740/34iPl
jxnuUVJNXtlcv3UNH3ldh9jFMv4KTdA2mCQozZX12r29zn8tfqfB/6QU56FhP7kdB0/6rH1JdjQj
du6vzkk3t/a/121A78JN0SlFfLEce+mtuNcHahPqd1vnyDm1elmbTnv5TNtmmVXM+22PIvttyor0
rg5Y3YOJUuV2LlT+Ec+sZ+6evkDIKund4HpXtRwh5tGrhpeMEZO5/ByNg/c3E2qUhs8Kvf1wo/S7
PI691SeG7NUSdeNR0RAO+wvPwiacUPCBx7M6wc7fJm/ANHXK9Z7Ner44VBAzXQD532zfxQvvo4W8
gRQtAynUF1PIRKyjskGHvjnR19qs868z2EP9hWl2GaXG6J45RbsOH3B5kyX0v30QvxdUGkU4cc/N
ZUGiKJUc3F8I1nNcDTH4RxFGWxQZ8UIPBi49hyfg1yjTyLLbWxQbTb9PlT7vnse2JXv0ZtgtBEMS
U42gveHqfj2KzYtWXQ6r1JymPQX4MQoY6QmaPYIof+JKR5FwdacnKl9La61yAGsOat3Ypx/xOUWs
9LRHZQduifdtNqtBV59UBl9FqI9zHUM27cISeyCki21wm5rxs7wkorSAvVB7JS200G/TH0YAIS0A
S9v/d6C31UH9u86DZBZ4UCKQ9/ggYO+zjNBbvs4MyjMDU3kLCk5S0esq/3xS8WJsneQuKFTf4p8w
81c9wPb2Fs6DU8p8uOxRhDJwW9VlbaCptsswaoSvcUp3SsrsxPZ6knmrDIGscIOzbCiv24Abhl6x
ms/Jq9sOEWxaK7+IgA4VYHhsbBSx7T0YsCXYRsilywITs64WYc/WV1ZDVRm5a79+7EqsajRjcRwO
/3r3NUvi24Kji6ThbPkoHKK1FJU4xDo4zEPR0pjQqDWsYBDUfOjZ2p8pz/ZvI5VB+ydpFKtAN8sf
VHRNVTPhMzkpEs3eiAkzz7KanKIHjNNXTNZGSW2LI87jIJoNgSsAIUSVYnpSq59fTqIzOZfJ7HYe
ByWbrjEO5ysUJH/MjVMRwrkFXDp9sV4d+WjjRs0YqFaMYXhLqYe/+OhtHsO7qXV4zWN5KfZxH2k2
Vt9LFCcejOcAY6wNMqBS7EC4i9t9111uAzvCg4C92dViGNeQYDqgdvCN6jHd3+Ts7L4wcCkW4Vgk
jFBj599KUq3d01HjX3HzN/VLfLaPDDyrENhuVhUHGEXZhhhpIqtD2k3ridS6F9zhcHQZf4AQxlrq
5NM62s2SQsGzexdekxEuqEoKLu8TO9+/h8MqmVu6gTtTwVy1jNYE2FkgtRYNa2sX2AFv/8XPX+LM
6i66qvz6sfmmtZKcYbrh5BmzOrxQRHKaqwSf7FeL/5MsEe97vRT+4Jimfns7SXoDX7jBnLgFfosr
dsrt0JGKV8iWHS166KFPFsofo6we65QURB75Jxjam/hrzh1Un8PtB+AB4co6HyTDNm6CeHAL5YTT
aJHXxd4/IUT8x4QcG+A1hdp8V4F9AaqrYPuR+NMw8jpN47cET6ooQGv/BFvjWK2dthta3IrEglfA
pJnkeptj6G4A8HT9TKljTcX6atwPLKyqf9DS789O6s0y4lwpHpIMFfYTUGHju9Dn8QJxL+BuUw0l
Qvhyi30y5OJ+lmtoPh98X3gAAmITKG6moaixjbU/4Q1SGrmMjuXhzFkByofVPmCTRj6qy94s0Ns5
yfZSRhAQSYe2tMMFOqgvpWtSs/kn/tub+2bwMnzNVaNEmoyNVFzBFnRr3ToowMx+3LUksfr2Rzky
R7jqB+LYjRcbMGchK7Wq2OqDmsQZlKywdZzKHfYVV89uOec1kPRF26THUY0Y6XmWiPCr1Jwll8oc
vfjUaBKQkhv/prFvgqkPhbnwXPv9dR51wIDqE9AVzyvC/D8eHpSDljAI7UNJqj5XnsvatQtfot+d
bPlrsHevCAl5boWW2K3aY9NsNRZOCIJLTI5DPx5Oh4U5qX4rQfKgj3YmVs2w7Tq9rlVtQlUQ5bnl
Ci84wjK74YO+Tmdu+bdyV6WPlrutl5y9vaGSEu5+ZBmhYkVbnXq2mmhrpXDMBH2kKleEN2yTAcop
JPJ6PedT7zWp49nRtsKGd+bhGY3lAmHveyJ0mKjJA+kaP3OarDrKbEOLgh+1MObQTCUXSeRkFG0Z
00f6z6SOny32wkt57yXJd0bUpX2VcW9eDg4Ewz1o3dSrBWtIidYhQaLsWOBJh1MiLtLFpaVP1AEp
u2hsPpeplICo4xOx06azPjBwRHh8dhODMObQhBt1FMqOx1F7xGStBlTwwnm+CPUFOCYUXp/YI7s3
yNqAw47WYN6I3nHsGI8P4BpF+PZZAKLgqfV5g/hjKrHJTfDHizOQ2b9RRRzofFmZ9aT7y6L+dA8x
PZ8L9C9q3VnOJlEaanUikZ9HyrWrhNHxFWrSX7Soj9alOPSbhA+gqsZcJuqgXAsGyQIGlTyyLEqK
dECd94mUM5g/bgdriC1KwwORxgutZoE9/FKThYbhFMwiDEZK+AxrfEaiEleHrv9JkSd89BGJXWHC
onXmGILuY5GzdiGS4TBGFWwEFF6qmJhAa3HleV+V6CLDFT7+hT5HCNweKr7V+Kh2o1dQ3ZNWV2bB
+bUAwNamBhBN+io9xkWVZnA6Z+IQaFISrljlrwO9xqC2Q/dKZisWTGSL29xZz/I7AdgNMTKl3glP
oK2zb5g98OHkSjCu0aoui2WWpHnJjMEXkJvHqorhylhQs/BHYgOLqkxP6oiItCHAoT0wtinA34gT
rLx2NpLo1C8dzazC3+6GEXamcEbQHOA+qwcEfqF9JtpgaPTHdVqIsUFf6iae5rwKaQNSjyUnf6QN
LW+xqZhuCObo6QKXtVxKWN4T0GKcqE3XxIcIhY8Q/NX55q8YFUuXT8Bl3NHQ/RwIAftm+ndT9oUl
KaGufpGmLotqKH2Z2yzxIz0GVgnPTWrcussgvo3SHBjjCnQQ725Yn6upfOOr/dVhkg2crxXFLb9L
8r1JC9dW0m3nQPkEvJ2xm/C8AdSl6B1kqekHhjy72P9X8oOFTUpaQy3q2CQ8Cvqof5WLCg5dSoo8
uqAXZbLiY/MmfLfManUbmn4utyaG6pK7yPDMpm/55jkhohDb7kLE3GGJgT6jOSEGhkKehBvojdDk
j84lsV0wEsdJULL1AWl2wriYXp0+UKpVgrZCME57xaB1zlhfs2uPQuEs/YfwxdwQkuW41l1vAPn6
SZ5Sacrd0kRuk4tKcdtdrQDC76TOFKwO4XjFvbf22cbSs2GMmGUPvfy7A/ScCPizzn1iQN/c9C5J
z9CrlEs87HlXcpG0+1q2Y4dog7gY/fQ8xEAEEW2FNeL73smZ0ePj1TO/yLThtllNslhpJbp8jRR6
melD7zrTD9Pp0oxH6cZwFB5yY0zEsaclRw+c2oGWjPaZb2SRo9nk0Wk71hj6IYbw2eMgfCwvBGYI
k3y5v46oU4t0VQkolEa1TgscIkJ/FpMCXjtEkmj5jMeGKd0Sq/JuUa/tu4QNSeqjbRUa7d32/ITo
S24EpZwMVUBjh3/5kkyLFGYCCnwmOBSDZlyos8QwxQhdqj/mwuVOfm91LKpG3A6hjox08qp4zaai
wzbAXOw74WoahgkekX2YGT75KmDj6MBpKlzUl+YogEvTJaal72hS2Pr9c/ws6OrvB+PgayCeMb0S
MLOhIgUODQ3uubgpckbUymug2CN2qFRnNBkNf3J8G4v+erB+hsBxx1o4yP4F7QguW8lg0s9d5E3/
T/lBptApCpGFt5MksW5XqOywXenDGhcL1fpcPtdeoqBevuh3oIOk1+5q3mwvKJWWu3nck7p5Vj5W
8KU2jWBD+ivaqIHFr6FlM3nS+d3P+YKf4kztoIa93tva6BSfFjvUmzk8RcUuUs/5n/puby88tNjj
Pr3zb73ukZJr2i7nI6nnm1lFNbC+ulgxxw2O/1gT+UGiHsgznCuVpaneR6WpU2D+mCAIOXieh10x
BrnJJkcJKhO9b5YUOV1Np8vQe9HI9xjK9Lp1pNS4yqnItlAg2xQduDO6itKExkPcTugtv7JgP8Dx
F66Z2OawsKCTDJyA1d8MOU4o05K/SE6ZOfUzYzw9KulOJmlFYpD9BnjTH+NLQcWXjYdX45D72n7s
gq40jukEmeM7kXh7tJpr1toIumythkuka8INZfjmTeng7F0YeBb7TDThWQAol/APIqY6+fVnTEnv
Oc5eecawwxmlIyEG5wZg0rUa1m0hxKW//qWnWCxYLFvSmuo+ZwG6CVCdqiNTeThxC6k8Wq6RbYq+
jHuxUU1DEUDREOsY1uW6uVlt5AAarZWbGxnn5UXWeEVnEwhxjbCL/Qhjts/Qnwcwp4R0qvuVddIG
LSiJ81Hi1w07s/71txfv3hhJLeXFT4Y3ePrdZ/BiP3IkYLJw4DwvBTF1LztH0mB2XEZ4Gz8HwNQa
yPrgAvZvpTbXgGyEslWCJdWdgq4JCS3Q+aA14IojhmaEVtcEB4DFNqzh2pMW8G7AjqTSTBHxOwPj
dD2/LPTE2WZ9O3WblKXZjvbJrq69+CKMHVQNwX+gY/frlgbQDqhtb4+xtqEFwKPXhjNJK6r0iLII
DjEScVF3ZpJAuhpp8cjlDYAJQn9qCAM/sOl6HkPvW+ZxW6wMk2RvFJlhdWTPxT4L9iD9kk7FQsCZ
DO45d1kT+KTtAqX8exV0HL78G9GAnRtFa3xjG2X6gRHb3ebUa3zN3/5CJbfHoFj+2TDrJn8pG7LP
Xi1owCKZzqHistoRsF+NQcG5vie+SOn50IHDGVBxv5UEEKmK2UC3DzZcFniHXA0mOa/SSHPmNl5q
p6PX5LdnSqDrRxheRZZBqxDf5buGpn9siuD3BSBos+0gcumZPrwm+A+mNsWVYiha4tSvjTKLLOSK
cvnlY/jHGfxJTrfsdTLtrQwLTCTZGj5zTOvR8b/RiTacNUHe21rxTB9+iVZoN1JOCrPwPVsOoQOv
s1Zo/E4/xa/veWl7260m90afEKRqX/aLBhrrNDdXwbxHSIcHjCAwwcflHSLqpluCzASLLdpxv8ls
14k1bXj1DkZuCguasnox4OGFGyK7TB1aREDyqXU/7yzPhXVbLDyJioGA3lSOZ496nrJBrvsfeJps
VLSVmF3MvlL7GrBtmoQ2fscfpCIi1Z0vfIcnO/g44ynOG7SGD87iXoA8vRs3gp5uNGM2uJ8HTbsw
i/S7OrXv4ep0nlqegL1AmkI/tol3v/Pc3alAbWBKHH11p2seWmScAiKqKm8vvMRALvolI68+dZJY
nAHUqCppnmNQNpGpM+Aa4RkBlmO8m2ft5M5ExdEqlJzK4gPji0Evq7Gj03LK4AGVKq2OKwOGgokb
uoMvYoAa+1+jS1mXmWdzfjkkGEc8BRkzoRZhySrkUKA4/NYAt2AEjZVGw5RHwdpziexkvyIxHmKL
x9uy4vPkkopef3eGUEoXAp++1+lyOumZneojI20cCdD2dGHccYQpMCMep6fd7AqA/NbWL4O1IdVm
0yT82U+kytIBhumj90blNrrl6cJ5z2nYkdA1V90KXl30usc1qAWQWs+Ujk8i1zVHj9Fm1oVzEmJk
R0DWoHjMmZCoqU6eWu5aQa1piQSjBKIhlDY19tLpCOtjpkNbEbow3gZS8eCST1JT+hgTwSuhN9ci
TfBz2SyJ7NwovFKYHHPILQvQTT9s6IHTYh8xjE6WeIqe/uMLSMzhBe1jJltHraZO7CJYwjpnvwMT
jSUcA0qcz3bMwrV5XFmpjLqCJO0vLMjWv4YGPTwJ/QL1FdICV/8PsB0kO1NP05WG/1SBNz5d4fUp
krIfy+xUQt7xP7D8Muvfv6g1PyED7cq1wE7VmqEin1xEG9u1DAjjLyO+d+ywbmGYOFi/lK9VrRmG
4X9eZ6ZqdZWNy70F+/MVSTHirowutF3Pq8Bwe2IwwZ9fb0CztkjUIviSOIC/eAY+Gm11lr6fNCoc
GdseEQq4KvhzGbzVaQcLzPdyKX6tKW7Mek1ptL0qTuWo18ppnBWM4j62+m/95REXfU7V0z8on93L
mOBJrfjFA0B61f40zZNlJ32v53wN9vKD26j8apIBdOTEpb/Rgwcyhljw5k8fZ/ADEsLe4OywtlWZ
P1fBsD6zM4KWhC8/vIV70CJwNHtKgv8ApJC0Xog+7/5AhuwKE79x+26MsjGeHQm7p7J3HX308rCx
beSV4DOY3ZzPNBHJ0AGerOj0JfCz9XR6OaD/lai3VVD9DjIgYAtdsgOc+kdJrVS++PlAOkKVJvD2
jQQBwAxeoXF51n2pMZVZNiO7WLKqUiYphqOufW2FJLDBz1Ktu5daGvOh+MXE+PneZ0mdEvbW5UVz
Av/A+Ckiam7ehV6iktP2CXbHxPQEMeOEZ+ssql/Re4ntPtYAzslFKXgNBp13iiMplk2NLiUVlq/E
S+fQYdva4god0GJuEt6SX4dO5V2VrDaJlrtIi4f4gD7LETFzympH5wHAgQoWQABvR7GxI8wbcA1o
7aauOk09IwYJiXUAJDrzGXrHI2g55GKMmyvRuUPqoo01UGSpH9Z5VpV22qk1VeKWzfuK8MZf8M6s
Pnbr7a4pSYMpjDsZNxcVyaNQxx2QW/+p5uqhclT6A/I3wpjoXsoH6l1QT2EZP++plxGR3+t6aOzX
fMdSuOjaHqQiPPP47IEpFQqzgZWiZJPuhX21dgCR0yNIdZ/jnuksDQvGkyQiMKGR24hDun7KSmQu
ngYP3RpSijCnpO62Ws95c8jM5NLNAwouwCRswGvrLijOACP+GvQBXqZbbBHY2IY0TPnoOaFbn6tt
w4Ubr/zqZoQtM3nU+WdCnQ18qf3lvQGk8eidD3s6csk9+bKWk19r4JAx4ZG86mgafHpHtXRAwdKM
5BHt2/u5ED+TIATxg2gIloJXG99ZuduPBSpnqP5aPSTT05sNwNOsWjZ/LJ5tYrg4Dav6q1EDvNCY
oo3nsnce9phIuHDSnYsWivj2K+EUlemdPlqhaUq5ZPXFUmqUxBmbL1C4icdnbdp+Da9ILbAuXApr
vo9q12VMlMnRJDAa1KSvXON/12o25dh4TPgQeyoe6IinX/BAbSD9KtlZwGmTxJZFm+F5w4dB8FUH
UaWKJfze7msd8cD0nXPMuyIJAt5Q25PZCw129dAdWCOK56+lUcqr7pECbfyLMqtmWp78EEPeoiAs
LlQ4oRJ5vwGTO30GnOGeoHJiA4IFU88/+7gsGuHVZkHabjfJ0+vRjIyYKPddSr1iPbR/I8xUYmuA
taljYuXEKDULjiay5tl3sgzirvDp5RLj0lcmXkyc3Pu+iZ5YulL/+FGx4T17C9207ueYFh0B8QPO
As4C1f2tw6JZegAkGSt1pSeYUJLs8GrZ3wKClO1s5WsJUKvurW1Oi2ukrndg0RW4TvQSn9FlecT0
31VvYoO3c2N/kQ0BCGhlFVO5x7nzshl88Q5FdmWMF+JcNNdK7wyUnWnqK2ytuZM3r4nXjSHQ/1C9
GcSoS0pwhiXpPzl/N81iCEkM4gBxu6Wi+sCy3dRz66o26ZIvrsRTt66HgURTKCCMMf7jBhxucv7L
YfVfnVkSHa3l2M5L6oBCcbFuYNdpPz0QL1qizU+w/nm2bAvQZmKWPtTc6EgT1QNL57UJvMQB1J9r
uYz4HwEdiVYFX2LCJUh/QARvuF1W46vrhd+j8arcQgAkO+A4kVUfYC1YTydCZVbjLcin4aSGVNEk
AGPutQvuxFUIUgT4ryTF38gylaJxtTU3RnBGLitNkT5gnh9XYWCAusF9mD8gf9+yPg+1eBddg2FV
9WG7M2TUeK0G+uvHb1r7qXfOTSJoUBAfU01zDHwTyIxlnI4mw6LExC/B+ijvOB5A4CzLwNnvWh5x
+ccSKI8d26MkzvhxE8QGvUzshKGSt9+QmQakDX+x3D+zG+EHh4vn/ZaTqQ1GaegpYEmFGkt9VyKl
ZyuwNYqEd95N4lPnFNxt4kAPlz0135IYrN0CgE2JJSA1HnVuwhaCXtCzukfIK5fWL1dBomacEfIc
wKw5UKRjvg6GrL32Ul2aJ5wgQAR5NY7aRdghQtgULTA3NxdRQiJHjwpFQO3X09PKACEw5+sGV0wE
YHOFcTaRTRWxvzVAXUycgmnjS7UDilvlvu/pI+SwgoW3If9dxYVA35+8r4soT4grIkCeysgjqoFd
bNSYjbwpnv9DMhby+Lv23JEK4FqksoVP66jJi4RBNlrKlfOUYx9QsaAGHrBTVyRs6Baepbu097Gp
62qpJrXSE22cogD0Qrv+llUQurN07T+IwP6pHsrJG9FC2jZZouSj0JQmMmXhsUzMht+unQVNMPoi
PXXiyIzcjuoSWUGnaJ/3c6pBSaYniQFleSmB0MR8yYJCJyOqBgL4gHv6h1f63P4gXN8RKLTJ55Qc
ecYac8dgboL44s41CeZgCNhVfepPp0BFpVW50oGXdEMXBa5QT+FX6XAMjd0GjDUr6OXMQhNj9tZd
8vBpnAUS56fTg4wcngnjF/Fg88Ain6GosvnzQdfDJFDHSea67RZ9dVGmzaXzAvH/n9UXC1ShiRFx
50Sf45iLNQzg3kgeCJmQlXXmsm8UOW++zsvueuqhCXexlgzWWLohj8av91/b+ns1wSC69LernQ+2
H/lYJn7A7tCLC++vqe92rH8EzDvwdaUnup81fRdaPaPWz98JvwunJiwCWw6WYphsUUUQ8vYidmoT
RHrq/MYzHuSmT/dhs9rKy2Cn2TiIBsSR2XTou8OW1B1kEOhp7SVkRoZrbbnyRH3564OkRtGKxrHk
/w+K8qgs8tckRUOjPPmdeigRVGRxlsk92ONz/Q9C/wcK2vBcY442AyQV26yBgRtZ8GvZpNfkoO7D
H18g+C7nSopa5cNMtszoVZOZytnZmLrxKVjEZeNbhtyITimVxZijiUQmRAKuzNIZIhVWL/Ow1izU
jiOpABRcNr94/wMFE/0Uw/ua662+aUXFa3uMEWv7c950NVebfGDu2NJSpzWucO74I3RRq1DSy7Se
yb+KgCUz9JebmrVNIvwgs0Su0QQmRwES49ECaryMISu6GTy5hU07VznOlFi/ZU6p4xEpkZH2V8XN
sTDRAAyFqTsZIg3z598Fp0Cjb+BmiMwTMy7KbyFFaB4YaRsJovV4H5h05a5H+9n5yo1U4TBIYbkt
Jtbn3HUhDA+wSGfwIHRkKY9wfEtXygJ09Zdx9JpcH0DODfZhtqQs51rEfSxU7XyTJ9ljNR9V9JeE
BJXU6RPWPOfwaIa4ZQB1E4esd51QtwnayhPmDYQAE2seP5HokCtRziBSsH3lAcyXJmGWtfRJZH7f
lF9I0RDUPhgwfnK3n/ig4uNn5/LJ0zefx5XU8htYFIbUOicCA9rfn8LbBd8QgUMGsz7e4dZMv+M5
4FcY+hakU5OZwJNhEi3b9HFOTfwP/9QndD3m0Di/3LM5AbjTNJ+scO/cN2I2ROQ5bKsikb7HUyRl
SjCOJTLji3YhDTbJWq1Bq/2OsYkFJxYBSRG80a9AtgauIZjTmNhqF+NcPo5bhnbczbXlmXjCQ7y9
bNBSAuqn9kWW4NY3Ze/LZhCcAvP/HqPgXa86NauS5/hb3hwgkSetbh0FbZmnX3XSNR6/fwg35Qxn
nevCGByiDzZtdkdiOxMWYO+EY0ME64Gm1XhfFckhoHM4wLotowX06nZYcJ1QNH0cZwLoJC+OH8yC
ALA4dcE4sgI5xyPccK3WtrHg01JC8C1lEjy+HyP2rRR9APODWjH5pJnD8YYeAzvMfyaAD9T9JSq9
/mBweC+/uvQCn0wMWCeT2I8Li04hO7KPiIX8PBAkCGOuTXnb+c0ZxS0yTXc9dsVtuXVaFcthTsyd
Dibn512D3Ewg7RHcHdczSt2AGK64VXr7dXEgtEj8Mh2qktuSCdhvvdy/cEnb4lmtR3bMi1pMnz1X
8Oe+ezq3teI7x8Vq/x3ZFWdTWTJ2ide6Gnp2SVSq9EEhl8RcxzSBcfkBrlUszhvfO/QkLdBC9Rq8
wwx8mAwzGlJn8I8Tmrtmj12LYOhgKtDpAKZDf3tr0B6YCxPRrg7b7glpGuBtBKxYEPYkwWC2E/dJ
DJKv83dCbz7f9C7KIoCzKAdhDTuFmgoGxdswSi11yRJXGFCJt2VZ662HDP7ZeuqpnuRNHBIvRLP5
aMTT/zpBPR13hsM/CmQ+FQCg3Jv4JUmpDjXC/ta/Jr7ZPTaa2NlrDyckwHzbdLoP6hsPnjwfok0r
+t22cLx2bQYluYa6mvsqstoqcsFzYKPFSRdTYH3jjEIwisKSN2XmZp8Ac3uFrH1H8d4RUtAzxgZ6
hMdhI0eCn1VDHOapSsj5z1H3uv+F14EF1ye6Lr5tNFvJsX6WczSHszkJIB1zqpskcWQ8CxoKgW/z
31hHy/+jXTeI9U3T9glXvNiV47QRzdb/dQkPOnSKzvB2sN2igEAUxlKbwNwOxq15KlFzvnlxlMqz
fuOWSPjmVhA5kP7VL3+RbeZeiTfSS8+INwbE3pRHOjBF3+t4IsRmWPPvebdGrnoqu8UreClINVqO
D53V8BPHVzmMikW4ZB9R9JWgHE4SVG35c4lCAm9QhrEer6YZS5dZFtdeNsDAAalr9BXr5KsBg7Qw
04A+jiJoXLP45TU0iTe30HdYjB01qszrvMe9rY92qMXVjEPbsjfaKlK3vtMihWw9JbW+H4hk2uiQ
cbS5WP8y/ADwGdFALs51dogdGpzWlposGgXjjl89vef2z56jSLJJOBRa3YLv1sR6mz19EP1AAZg4
8kTc/AcvtM/n971LtOtqeMlemuK7G86ge2a3LGfbWMD+scl6obja2kx9+MPaCfa1rWJk1n3zWPNP
44h/O93hHIUx3TOajXE88Bbzfh0+Loc0vionKAS7G+Fsyo5p0M6qvVUl60So3LKYesy3AWQ0NKNm
gDuHcilsg+YYodyTsexr808tbP7mhjwFcS7GGctmzgzQOdGzP+Gbc4QHXgjlEFLIyhXkGrdiCn1X
T6sr+khQcqlk6lCeCPH2Osev8mWrHBlOgUJ+XhJz7SArw/nshDIq6OP+TrpsX6HuzfLULv7r2Lpu
wLWA8jV6MF2DrAOhsyl/+1ipSHoDe2INZ1aWUgqWvcNfl06CaTfuSNojo9UAOK8NVHuqqav+PxiZ
CNKcdAY/X54/iy10+e8dRkYZH3w6UuSCk9ynOAjGrPHPzv+Ath2mHaBM50JRWdqzWZF87CbdkFfC
eblmm7tMMDH+dLjtgMC3wMcNlAN1/S2CaFvZ1wloWxnqOiwMy2rr9exaLAPwRihnurw1RVDR5OxY
koY0NPbZ0BSb14Xyda8mypa58URCzPbp2uud5bFCpZ8t4/slwlDEWooWCr0WGf71k3EQPjuAXgBv
mu1eE86xamSE4ALmB5LsNAXiJJIj3rqXOD2vIiY5Gk9zsiXWTQiVwE1tykWR/2aLixMxT1pNFimj
yxUtPw4jLLsO0vsncuoWy7w6CkJ4I5S8neETB21HVVm7ymq5fjeTG6zkNHmqt0rvOXKNCV4xQyJd
8tEtneuT5TyocXh10a/bxyEhVqBVEerkgMIuRdDt+y8Pjcfrp2cA5QM66F0EcEca7DSwQjfFepuN
mqzcurIbtW3LAf8xTFD3galjh0aZu8YvDWTB8sj+5VfjrUqSBhhCiT+TNUa2k+7bgw98eW8Y2BXk
EdiX4zYYjnhJqyoMpHJgANFdy8FpWhyJ57REFqzHa6/cs4m3anNevJyc7twVT73IVehbttB00/Ky
P+IczTdcd2fLqJS2f7WCkDheTBMNSob321YLWRyzLVA5LXKw4MmLIea3ioaS4XKGUIvG0iUXyrcW
l+XVTwd4ERrgot1/0g9fWytyX3DKM3eHYXRGlRCVyxpJNinD2qEmJrccZ5sEVjvBcmjHKYc894Nt
Gmsdm0jO2nO84mSUrEdnuNSyii6AhobccXIaEQoBZJwweLslhKVreiFzpasEDKjrTK0GEYDRC45e
8aKu+a1IVg8+/qRvUvnF5H61YLRxPdYv+hhv+WpMryWtpWgaLm+UTgLS8eI8bIZbeU2nigNUTc4i
LO7xCwvxhlTZRd0XgWAMw394ut3XxFn15Zz1d8+ci3nhsPt953WsdIliPJgihlZwbTnPTyLq/h/i
QAw/mQNRiJAxpdUNWPnHZH8yCriGXn9tWGW4vrapIsIsVb/lC65hgbpP1283e0a57G4cZopw8wME
rD5p1jN5UywmVKbARsWRrmiEnGdcMNzUXz2JqzGa953NZGMtI19bfMg7LXaHl2eJRpI4+e9A2sj4
zaJZ4XdYpBX1wqh9q9JgjQY2oLqAw5Z1xC2G8L+99BgYdqRQA7lNGxVnfpRxRfZTxVefPAWCLVwy
LnybepuheJhqbojoJdQjUN2zdQqkq3wV9clzTKRNkknMNOY35bOyEp0JK5Gi1DVx0pMKwadXHPLM
ApT4VVMGnq2EvCpOBtOe2zDtL82amuFGM6Kej7hMuE5+XPhQBVS+17pqZfhtYDbcM4lbaX9BMGmD
JPzk3UYO4hw568alQkBKce2cywxnn65G6hoCdb3+jraHz8PRtg9Qd2BgutSO50lP1qate3cqugbd
+3kHt0Fd4J5zaAK01ooJAnjFNcuYQkDP8CR490phFyXAmiR4oAc35w/BYxNLYZHWvOKerYw9Xswr
6YVL5nYo9xl0CcEjHSOmS7k5Yrb/P4mt6QTjJRoLaY15B3LA/I+ti5vYIQfWgdlzLiH0XSUr12/l
Wmfq41pvsnXbTSQBUv8kJgELa+LXmScvo/hk5hHRMSUDbMvPywiWIn+TqAojkxr4+A6PmWT+d+5L
/67pPTrQNK8Y1ZVamc3cIb/lhA7YuhR6U7PmNhRNUdp3P1HFCNr4XWrweAMjCm2KyRvrWbBuGrU4
bYce6/VObrjDYqr3FFvUmlCbVqBzvysfBh8ve4+FndQpr04FcnOne11/2FhGl5W8qV7eWImLEopE
UnSlbmnNVByT+WHgcb+yGH2sxzd8kvSJR00IQBv0PIkt3MfB91kSuqCaasb9DeZDnHMiNaOvFX5H
Nem6KKmiDX/1uJdPkadeeVqumQSGI8XUqNtId1djUWmrbTroZwmG1jdEAx2yz2nGnLcCh7cRFMUb
LHsLunFdn6pjNnVBdv1abhF+8HLvDfzIjx+Vi6i6X30u1BRHTT7G7o2kLqywU0aQ4Gymb+Zimopn
EVtR2jX1hj60N0fgEHVZfqidNX/E+d7XqXukKKewkJ6vboHciHYsvaxxVUUiZAPJNW8ry2zajlRT
bNOam38uLM/w0BzTTiC2THpQIiq/6vyI/IEgLPahd8n+Fr+XvJjojAybbneciRt2ezYM8mktb7G+
Lqd/ljK55Akxw0DYju1Hiee0kI+c65eo3ts19DqWEPNPxMl5kpgkU1Fe8YAUUX8V9k5G7DWNN5JO
GHw5ZYO40vRxwKnKV2Q89M55pu8O5gWR1O7FaCp+VAnKOoWFUDj8dL+KZdtb96q0PJ3fSxlieZqF
mDj5+c4CybTeGyrh41bZFfvZGxsiBCZi7oLgb/sINNHKKG27FEhro5yc8VXiqhtUbpiGhHHcvIhR
y/T1cCYaC3FYojq/JxNmaEIsKNcbO60WocvipoNYmWCKVWd9w1MctzoFiveahs9ns1vXOLq1wJRC
iV/famI3NyyOd0Y4tQoqVUfGtwvITCVn8dfdL7iJ95i6O3SDHDUqi9cnYLPoyrA+P23SjRCivCoD
F+7o9ffhV5mXA4n5pTFTiM+k8p/eVrFZ68xedRToeZ8F/maFD+ulM2R3/KpxWIOcz7JlgKIc/I9b
u03kJJ/MBO8l0q2O4J4sIpSy5Eql1vlNsw8CKkLEVEipAbjfjCUm93Bk57IuROf4vxe0klai9i4r
EQTAR7ACcAx71RA5oNKl/bcncXIqvlK7t3QpgiK2yOdyLCn6ucporysO4NXJ1k2FCdS/em9MTYtR
i2t7V4wHphd+kfUX4c+UJvbIc83n1CK52g4rRwdbKAtoD8zYLDufKAErESXbUlaa6GScpA5TvhnH
cuUh5/uaWDUokmTsd03qln6z83FPtcXBExkVlHAsLxr5Q4Lfco5WGAkK5t+dO/Mi9LADc4N1dr4e
1msvzhcWdKQWdHtX31l5i7e+8u0oPZBu+FpGKgG8QbWOjbOyO8/L3sVn/V2nHwcdsXFr+L/AbuOo
slnqZ9vweBbSTsuECUqruWdscpqd8F9kJSjrPg7RaKME4F78U+lXQa8UTdHrA9D/U0ZWzg8bvcCS
C4VL5Tsc77KmIf4chmkxe7YshoMxEvKvr1Sok+hwFe7d4w/1i9APBUM2EzmQsDE5Au3l/bp1jnUU
TRF5KBxhnVJV5oLter4Hxq/BV0H5mpQctVB2x69z+ZRMUHUoj2s/NDrOIxN6GFjsK7y46NqcYpZT
jREAghuZk2nxHsTysZnudrOZ6Hvd9f8yKtZqXh9jHy45TyX1RMKv8919sNQ/w20seLZxWhCRVLiE
SOr657/BhAv6moxP3usWff2LxHDHGaNmzbS/B8GkM/xgfIeb7gb5iEuQKKk4+XuUAq4TaDycdWi3
sbYpgELTxYps6Ox0SqYOHK+Rb0PeSDTDOZ0i10o495IQqziQLrDFnSlJohqHemE6+xjkTIsOjW7G
q0pQOjPtfej4LO4x5bHQTbAVYOkS5pe5sfKIInqXKdUlr0nFr5bSy8Mt1G0oa4fRYM3bGDWZwiat
8r3giTizL9pFBZqmEP5joyK/3XQjG0Omt7J+5b3GgYSu4I4SjPoNMPJ5vA5+IzMN+UKmTyc64LRK
p+k39i5lGmt+dP5tz+yJU8gxQmRW2UngKvIjg3NZkSC3Q/2TegvfPkQLs6HHw5Q3xvPtsrCjLr5y
usqnI63ptNaztNi5svaCGcChIiQ6QRIE497+oTYbKsNSI0UmvEZfspWFti+MlnUQEZ0ORGasJdNy
LzceVTKyJH3/4jWX/mvUPGHjlwCjf51Dgtr6NrrlvZ5UUlVMQv5WSg0LFmQCGywWrRHFLJvHEe8/
2D4BhL8kihGefZFR1pJMBM1gBEuiu9zJPTQ8sbxqMJrf61aUZw6Uc+BvGC2StNsqfozpV4CxH0L2
11uynoTzb9D2ecYLXXay+Gtf8vztgJpFnIBRj68iTFM/AzKxUsWkh53gYx3rJzII/cH7vdoeqCFM
h6y6RqMJWdYCGro8E4c1oi4Fh08VCwDSAFVBUdp4oFZuoW4L6loBTSZnNQVk55uZXgD0gONIWXpk
M6ZDQeHSrdCWSOy0K37VOE9tLA2vsYt3S+mEURaSb8bHxKcR/pbGguRw8MI46pCshDFeKz2mFdhe
JoisZ0rcY/BOMxAbpl+34+5WjVdRMu4E0jdauZXt+TH9a2vHO7brq44s+nio56f5/xzZj1JQbDph
Slcb3Wi1Vv+DOcTxR591Fz18SYaXnieKsXlFfJpsHFlViapcUj7jcbD1H70I1tHmnCmC1ojRBmq3
UFrQd64wbGiGQnLd0XVmCrzenaoOFHnrJ9o86OF4CD+gD2xo6pmoZpY3qEAw7Ko+RcA17yQdA7kW
+UmNIKOYIK/MSlzsVfQq2i+CJPFZMVrabnjPm/Zr/KM0Ys+BUm3IGOgDC2w/2JdkL7U+duu2mY8h
13fevo4O1T6WkpVMmHOPcYu8UvfmQrBxEuKkIrv1Ein9tQ7f0w7JjKna3V5Q/jAaZRdOJHtaQs5I
kAO9Q4/EPgRlCZVS29qRO79VRXHW5dzXHeV0nJv335J5Z8i1uEQ1keWhnVKP3VCtzxaRDizmGvVS
W1momhFNHwdndd1sdl3ompAAzf6UC3pA8lyhRWyzsnA5JoiKMZkbHWaOd/9jky8Mrm5b+mbJ7fBb
rsciSH2fkPzYoZPGjW/7hTwjh9SBCKHxP7xdqb95laU2dVHV10lRM1d0Q1371+1qLRRv/xEmlcLr
lOJq5iRwXdFDW0QuhKE6iiEUBnsYLfZDGCHMC4yukUEVAl+nhOhgyTL7hnG+H8Jt/xAjMiGcSdta
zHX4GKIYC7QTFQzvASUB+2e+7Apqb7ugOs5fDy0hbDe0u1M+POrc79FZNgovKsPrMAkxfz2wEZcR
bp5rgQLv3maHFPhFifGIScNiHWBlA+IaYps8VB3Bi7fN2rtu1GGKJkRZsBA3Qw+k90BJuSzsjBDj
MtcmzLP+vsZa0+OwECkyeFDEaaz34+Qo335Cj8qaMwfhUyCb4E/ZRYUr/n87l9I8vbc+XJETGbLl
KntQJNQPXVTCXYlYKst/Xd43CVeSQv3ZpN0c0+Vfzs5lS6NYNyci2MSaOp9mo1MJPzT4j8PN8iD+
dyQSK4fsDPbtqLdfUDUc04yjg7BTrFH4Vj0HTFW7m93Wlfltz6qQ7BdQJhMXJzH4KkjUQRljNOXT
lODeyJr1tj8ZJzL/uTKInsvysSzlwU7TgtAGMGwWJd9jcD2kfkb/N4Mq5XCwGAKFEFE2WrRmjnK2
oKT1tK/bURv6ejInm2jEun7bcL+oazpJz6LSvkAkTO5EHuUFCF1+5b3vUzQyvxxNojVbc1H0kFxr
HcxNneGtJPhQeQkqw1ICCzV8epu+epbGwk+fNQC5hJLQX0NpD6uYyRAUmwyurNAKsVd1Unx4lqZ9
BNmZhrxOB+tHQEbHqKjw3R3gie3ygFBgAC78shS9kOJwOyUd1WYNisvjxncOUdjmgTyRJjv+AIFC
YAmzg+7K4V8B93TB5aZPb9SWShy9yOz2/eZ9Iy+RZZI7eCABFe9Tf34YT2Dekq7YWAXYgUwcDN8Z
/sdn/ENr6m7ab/Z+xcCxU0aU9CDziFw3oenptfC5xEZmDtYQgfjphTFOIeUIWlVcdZop/dpMA0K/
SQBngdDsrmbZr3fqrlAvGxXW0n/ZRYZKVjwprIAekOMYROSbaLstVCGSGYqlShnoHIUG6gaTR+up
MLdqaTs3nzCkWWAN2Ly+YPTPjBt1e/WhjclMBl+mGwt6CGk4MHnDo/MFAgR7PuLuqRVfe+VkDkqG
TyVQboPjtVy8JLnpKEkNG7UMS2GfH6Mh7zp2P2TY+7UMWaDpgyYRd2d8kaq4ukuJDNZ1DbikUlfP
56dUGbz8uURipUL/Y2seC/DRfG1gyQUjvkEVRZD39owpg3liZCJ/feCC/YWUYJIR1IQLEQdEhFrs
2rGSYceG0zw+Pf2x1EN17SrLBL1hwX0Tt5BovtVXE4kjVq8MCsFZ5GOlnBUpTQjMztBe323Ok7k0
OulgNpCFx8vqR8LRZpNoOA9SFeE2lFNaWrZHzpyrjFCWhBJex6i7fRhNhJ54isQtN3Bd0hWKyJr+
7D13Njs2yWIsadJCxxq/OwjO9BLCSBPQPMAOhYSUNCIBynvHvoFQsDpZrucSygZwmckibBJ9Bs1/
kEd9a6iNB4WIo+CSpB9hbsP/v/pvxGOSj3pdPN1srfIT6h0draXf3ndy8jL8T7ds4fuCPTEkmm3e
Jz85kYy20igZ/8Wn0ArliiyWO3qF6wAO4ROZZ4WWoRm7grB2Z3Q0TfoiepOd5LRITNiimz9n4CdM
a245tGwx4tFrYsye0Ny6eQ0Rd9jqUJ7N4LcUs6sKCtP3dpjhk11HVJv2zzrwdwmZptoiZqur96AU
oZVb2GzuaQMG8a9GhE73hINcZgBbiJe8IXdkn2UxGVl7yMPjpAh+ZID9DSuvBXYM6m5w8LCfLili
UcLIpM8ea0KaB31kwbj0rbngCWQPHCzdujlgASf/ZmWjsY8XIHT3rXaIjAmDQ+BBZiryRcTxZFA5
koQ5FGMYHIaEChLeKv+V2LYu0Id4+838vNHaGrB6DBjq8bIvyq/rJlXi5IyLzGO/zhc/iDCCEDPh
6tHNMDZcasnEgf2gXVdVi0uQWibAk17e/+Jdw+sbScHRWzPLKR1wxzKf22u7TXO4eWgXlNu08jFr
+U34Uyr6mV3fScs9udkrEkpIM+1l7JbbKT9LmL8LIE4MwLfAObTVtn9Mexxty3I/gZVG5cWT1cYi
1TS+6k1NBulIbdSKcK2eSv3nvep4RPDLSmAWxOoHVQNjmz2suEIyJuiCHKhIHysrNOymrFn6FfoC
woIz7m8fjoy624RlFDwSy/pG1iQ/loWm95oJgfiOX16HPm/AuVC5wemXhXzcr4FC0p4ZuaFLldMA
A0s+d64scBDZeVHwSqHwGomtzPYCbYoqZuruBot+qXP3cIRLgCd8z3hZCmNnS/EwtFVGmpH55BFj
2y6Rs+6Qh+QdP/Dhzy4uu8+o0Maja76FWp7y+sWT6sD1gT5EPcSmuZnXxO3NIx9YexWWtZiamRMo
msezYeXTsRFfQIu0UPKmfvOprMSKeb1chYzWqX3J193QcvjsAwizjdnN+dg/NSAqnZBl2cjxiylV
77F0djJ89WmmuzknTrjaAmmvX0i6ZtWnOrgnBs+qvU0IDAGDdiIcINnYzv1FzYazp0JdchbWlszw
PbaEVHbaIE2cNH/e9mm2SbV+1suROH2c9GwOlj3wlM0UzJ5CHj43qyjORX1GxzABIz7cHZfrtqEs
XkWo1EeNkOi82Gc80zzL4wj0GsfFz282piwTMiCoGbUBgj9eJ9Q/xVCz4e1OY3B3HJljMkYnAztQ
T+ht91zDmdAhpdUHlpTT8HWyXmFH/sSN2bwQs4S/QQ8DrbsBoTROHOWuG9n493al2OjaXWDPrcaK
OU79qzYkSwPG5ID86x1JB1mhGMI8NskgsysL+j1vhdhAU9xpTLE1RCSDfw0JxPiA5KC2JL+fpfEq
MkWRYY2LqH8Bfxli85DnK192UEHjJDqAaR7Cb6UxhcZAXQS3cYQ6P0VUWd/VHikXiuVPGBbNI0Rp
oSFYX99ZrYWVrx03XaCKIoJy5Xpu+wap58pkKhRgA/XumpAX3lCNRZK6/hMFJcxXypLU3oUEl4M0
R9AgSXcN3pzy6nehBlCitEe8DHBZtPd0ez2KYR2BumuGLxrT3DcBR3GcLQgknk7ZEgHyM7v6x6mH
uj43CznOaLpwtghZ48rOSbUiLoqGoLLfYAyr+n1IQ7O8UwvO4gUXP0ruJ7H8ytZeCqZAREDCxpcP
o77D7s6Q69/NjZPVDU0mFcza+Ag7E56wMehny+pCoY6oQBwJ8n2b6FdZ8SWUxAkJreWwGapZcO73
Zc6XCe8AmsjrZfyuw7u0Ex3Y3Ok6gy6kJPR7U63OjAbN3eE+jBPXFQbVXdXO+zRZzfpoBsEVsRA3
BG5KtWU21rSLpvROAGQUbOl3CCj3m2O7BwrUqp3fPESkCHhUpTjNR/PQyjpsfwtxGjau2E9PwSGk
QngY995h36a0S6AZqyW9t2hf5IHj22ZR+AVVublCpSIA8J3I7E3C5qGJczanoKt/OqtJ6/3wQD08
NLMNBs5XGfgnedhmP/GpCXUXKamQNRcex4yRC+j7nlbRdNBfG3TVk5hpl4hov1y75mp+p2PUHgki
DvsHyph25Ygum1CtH+EkcbqszksVKHgubgv5QWOMbXTXlouX6EM0yS9GvkZ2dyEr94YSj+Gr618P
4lcGVEIl65r96loVBatQUYk6Sb7wTZb/sIiFoBXvYQhzkFJe1v9DMZ8OEerGtpbTTGKbWovs4Sj/
/hTVJg69nnQVRyNSZIPiQ/l1P2ZbBeiyJ9JmYBpr+QRcSxfyScdfKrmdw9pNtM+XDu0Szxvow/Mp
1H3qEzeZB5mnoFrjV702y8ZYOdCkzPldCNzYrIc11wKR0Jb2AxEhvuko/eA1+acV4E9sHwwH1KH5
dCOpb4wekz16ORb3vza3/0SlcdVj0w/IohoB0aDNTaT3dUbUI383b2cGm7v8Kn+c1xBEKnI7ypkb
dXt9ntUiXwpHvVJHTWPz2JOOG899RawaXbgNJe5JM2sxFjX1LI/9om7djnt+nCnUI1Rb/dk64bOG
otezU4EZeEnytigfQ//bUeh1MxFp7k38MCU9nbwSVGEcwXvWBrTx4c1JMEZ/cnVSgcb1K5sT9mUk
damIbz+z/f9DP2EzJMm+DENp4mQDvIK/lIJu/8Uc0TuyWGy7UxMtwiUpl67sPw2vTiyYrKGSogVN
ZVvFqk/EiykJGI/IcPa5my8EpIi+ervXGcKExymTyyfaLHbcKsQNp2Dk+3z/iBlDK3NENdjLrVYy
251CSo5SWYeV8wuEhwsj41mSqumt4hIR2EQyUd/8s55MIVMNjOwyqurwTdjFV3jCX1x+iyteAWvR
fUOuwM+7BYxO+w5r5Q8ll6cALVJCDskrYByDHsJSm47hlsY0Rf+I+YYcrLpKhBzs5E9agd2d+fkg
EdiUdHJBqQK+b7+xioTBIPpUtenfbnBoLpRu1v5gqXbMPXBLHfZgXNX0CLwo862t1a4V3exxA9B9
QuLZNmGNU4xOFzecYUVvo16VDxHNpBHUmb7uwlr6ZUOQICXlg6UomjanRyqqRd9QMonUGuzzCg6W
bZ0QNgs3ECXk/w405UJYPxN7Cnz1srJjtxiP9xA6rLKcmHFVR7kt28Ao1TtHYbqxY/kxckfUw8bt
LpkgUh7qTKP8VevzXwtothW3RVf5B05VkvyhCl71vTyxNqEEk4Llk0/uNgGJO7+nbb/fhpE++E/7
PtCma3OW48+46j3hd9vOnMgr8C1lyQ35lOdCzXufqzPHRud72a1UorSnQML07qDGSk3QY42vJ1o+
ZMyLU96hmGlSVvBxMtdjC2R0qR2TAndaBOElIQeEt5irknL7jK+QShlhlVZIVFwpN/tcQ7BvR2oT
VXtKmucacd7mX5M25ooHzOfZveJMmvxxW0JsffLrww6tlom2hlQMSIyJlQ9C3AMMVlyABUHIrWda
UO0pnCjIczLqbTub+kydb6Rfk5IOrb5ZEycWcptATvOeIs4mYXCiWRzirckR90JCaxPtd3ymBncu
pzlxlAOehRpF5QPLPOiLAyIWe9eWbBxkCnitZoEMsvqmLPQyelten/royfZrobk+DUWsaTby+o6A
cE9ZSubCI0qlhxCSJFLt+dqTC7x0pvxFEHFx1bRJsRSzVEIyjaLGryiTos6Yk/HqgZawHLpYtR/V
shHqO6JpFI3rtlIPavse3IllMKRjIhfEIqq0RqgpzTPnz44NMzfPtCkH1xO4JyIIRFl39eXpYM3n
HVvnwm2d7/Ye9nyU2vWoHfiFTm615ULsRhdAih7UVnCcoaMTlxcS53zRdwumw/CoNUtW1bPsW/n5
MV/Wy7ND5KEzNebO8zdtIFLlFnb8X6D7qmeVfkpF55EWigS7qcOFuYFMVwza8VTleBTxngnfhZzP
sspMWjcMlV+CagVkK49yZ/DpvPvUM/tUDNBdeVa8J7Fd7BaiT9jKntMyg5rbLBKXnaWyYJKVRfbo
qJVH2+ysONJKl6mWpLULP+UUfJ239DjRcFAY4+Ixtq7jE37JcPs4nFoZCkjzZ8S1otnjUEWnxgmA
d566aMQ0kMrgFW/J+A4aKBFOo0UJQIoT3lcOpG6oBqAZNf2B2VPPL1UxriZFYvUYo6YL9zBV7hd8
0HldYzHxmS53mtl18jUnUBEzKj7r2DVW/sBrGQWgoKRM6hbD68jt4Qru7VVwrCISmOfw3MP9uhVq
ExZfNhdBqzc7Ve65g7PS3GqwDCHr04MRMbY/T8kNv/p9LmCzqHiMMGO40swj4pik/xXeZsknkpQj
zwDPM+PAcWZJTp1LACkOpRykWYPEzSOloFEb3/lS0bKHJQrAz34NzcSbm+0zvbEhFxPxU6kl2qgX
YYePk9tfAnK4UTU0UEjQaxfBkyzFtKmtI5keEW5x7RX17zv8WB19ekPTH6C6ZJ2nR0GY/EY+PwqS
qGCo+u4ZSk9IzH29NrwQ9mPrAy6FiCElUSrXmrCVeNZoXwaTJ06zR0UVQ7nLjsjGpD+dTCfgw+1E
2bkNYoPTjtLBX7n2SmBV/1maKgzwqK3aPKIjq6Wit1ISBRSyN9jeYx5DOGNzzlofxxBgScHX4G8/
DKFvLIg+WrvpxfWqqOqf0jy1O33BDOtZ+prnDtXRfGz5XF93oRfAWV3wiDjNXHV6vXqQKO89W+F2
/TDEVs+XlBT/A1qNJ+qH/yKuIabMqD/MsJW7R3QFgrHKcybT72pIVUtVCJqsnD9CzttlXdcH9uID
GMNxyOEjlr6mQhJncszZgDKMDzLHz98eFnW8HKILyghtlJZ61AoQz6JVQLWBrf6SFXo6XYpg783p
S4K0rdrgNmYcn7u4hJJ9kGyHXyUX1dTfOvYL3/L8v8JsHNqsCz8GYxev7Vnx3G6YnXb/Lr926yVO
yL72G6UYNP/VKIFBro2kdLmfKRfjyoZAMymW7heCQ9rh9Xi3mCqMxtVuc0VQ8iGs5zxtDXRZrygU
+XmjDMrnSoGA0Fiaj3XETH6y4yA+92DemifpVzhNRIlI42dCy0Kyor7xrd/AN1Wn79wi/nXRZkp/
uOMwDBW8olWS720TD9rd1I/WPI5Yx+zE1VekqrkviiRmSpsK7QmfuTdryHy7tNLj27LO/9T3D3NP
RWoBVjtL6UKlFuqAIV3FBoR72g3NGdPMDpaC9/ziO5rmTr2zwty+UZi5tXtkaBpw1aWMfX2nfQK7
OO0iS1GX8lLeXAIXDsxk+nN3LIV0gu7ox+s1hHXB8+cKMaoXOla56oz6V4rrf7fL5pL9tjQ2gUew
AVcQJl6Pqhl/U4j4M6XZbHGGmrewhCnkH8RGTTsR+vvGYBPMG2yoo8hRVS3VCQ/XyfQMCKNT1jXP
XRul78ZIp/31O8UFJnFj9A/GqpVh7oIgGM8ipsp0yyEy64L5ZVsoT3hwETJzgr4/wa1CBGFnVMkb
OSULCdP86TntUSA2fwFWAACaROcedKkrHWStJe953WbO6ai2TlDUclrWzeL16vwhDG6dyB3zdUtx
mqTUriv/vxi73/TS29bd5SXQlTEE2geLEQxJcIgwJLip/q1SnrU6mIFFHnM3M1LhAOzDP0Pszq+n
92QoA+j5biyM6pwo5DsPlIpL24S3JAXx0a5ikkX2S2FK1ZPg/QLwHn6upYRTvCleZP/IrWV4+9/G
koiNDMLdDpmW+2na+seasdqdEBKowQuEG4YNfCZKyiLsIlpqqTJAOEIuQRvAXjNGhMwJ3sWeAWbi
BOuynblINuU4+LYtkD5TfmIxt7ELosiTzCELQN+udkyO+NSboPtz6oK+Ki2eMjhWy2V4uPITHUcT
sSvFjINvXlIstCrnMIkv5MO1R6IfBuCGaXrFW59JYRjQyZ+hzO4JkAlohr/l5NpFPtBeUBb4gc56
V8Ir83c7xyqM1VYZvmclM/D+Phz6DYn1rTcu670WrDlB9mSlHGNSV0mBSSWbwdMQrqQQWPj5W4Sl
7PpnaceUKhMyNj31XYNZlUZv2xPzzWQDAfphnBExI+Nc4bIA7Sa8EBB2qvcFOokuOnFTLddWLLG3
zWe0iH5J3Yw2ZpFuffk46cBHCjwMT9Kq+GK8NgXU/p0eqxPn2zXo4PowgSRKLvLdwaxwoEJKIOSc
njH6TgzNHDij2EU+lkzk8lZWnV6Qm3FhP+z/1OEjU2l0wsIR2YjnjRG0NxSXoCuYE+1Uax1Qr9Ec
FR+KQoC70W2I6SS7+g+Sji/6FHpe0DDaMcQ7F3tKKUwJVgEoW4LKy0DcG9pRbpDXNvpvhZ/qwqpj
mRl69Y6ccO6lihdPYCXhh+JRGC95jTf+j3Xgnocz6RFGes18QfTQQbtURoFNX/uI34z3PxfsF81R
CvB6yOr5qRB8CobNPUJIW5MBYl3D1sFDMn7Gsc4bz2dKciqlpudYmzzx9VeHntVAAl9EbdUtnite
VzX8oX0SjKidHOXtuBc/jX7tcmqMYFHtO+qUDgmXx21kX23rUMqLMKNsmjgc3MZoSKaOdsDoJdu/
dcn7LvCHh03qADdjCoym7ZI17fmNgK8WBmrVwEQ5ve31NEtscGt3UZDOFIkBOHdK0kMkqE4fKper
9EKJU+FNOeQtJotRd5c8viKfXAprP0jce3cbIj6/10l9Yelj93oXqxXcOAoaEvc/Njq5Qul1iPah
lxNHU+CC3c41ElsdBSGkmcVui1HcXjPBe+kRvqYPQ/UTdaCYeyZ6pLMpMJQS+pt5+BIwUUge4r3H
uRNGagcnIl9RE7KzDj47iA6O4krzvjC2GC2LfuHYGQWTr8O/kHokg4TipB4nRhta9PHX1ThKt2ZU
ZUiAOLYGzD9VKOrSs0ZqZWT4YQsyiSxrrfTUOYJ9t+LGIctEQUpiq+kSiMZvX5mhrkXf7uq6ewzA
5mv1DoBRm/XQVPxVX6/o5Lsvxjm26UDIhuntDNUkl1CpGN4yMMz2Vf18LcCIvglfWuJuAOxXvYYM
Pp0EEPG0uRZCswVf/j5/+OcwsdsLp1FEe2YksVwkMoiIkflHwqeco4c5PU4YLH8ZDcwG56s0TBYG
QPPTMV7ndbeJ4DCi7DffNaxpACLpo34Xv2Xdc2z3wd0anAD4TmqB5UIXg+pvsroLXDp4J9cVw9Qo
20YherSWjmrKLiNJUfEgZhsZ7ikQ0A8Ayk1r6Ca3Xgylfy0f9TwBnR531TB+AQ77td5xbr8zcRI3
8hf2ryruEmym/cAWxgHwgNLYysw/T5/VzAqt6QR7xpMg/CldvoM+rZELNwLZHjNry1ALcxat7oRl
FiP1P104u5HSCUSf3SsH2KItDkgcFMQcZOv1kQR1t6A8JXAFdi/X9gDqlfT0ZT3XqMZQ+HC1H+Ba
Onh8JO+UP1gQpNj+smyUJJgWDjVv2ghkW1SXJ9126Hgq62JqkZTN6axoOF59+3WMKbwVQNPJ5iXo
kJrfLrRUTC7UcoH7tTmSUAuN5gdC1YjHaFZw0nQV1X0eFVgsuD4KdgBGfAk4Uwoxi4vojLkL9505
/zpS1afsaC3IQD4c+B2k7Mer2euZRl6pESI0PN32UB88DegYTUjTmTDD8hIid9ftQBeS171G3bEv
FaWiTKXRZEbmS3avjDy1QM+FoKBmATk8C6BnFDTGcOgPV21DRzxu5sqid1vPaWdttoFECW0hPfH9
5igHaBFCq2cYGg9PgWuuT+J5GDpZm2g59qMNHdPAZdBeQs+BmIDfC2GTfz4rk65bVFgGkJGFBUxs
EllLoUiKQmXMAnMSOfANeL69uZ67DOBb50GmKryp9dcmuEjXRb2DGP3Y+iz3NKhck563/LjZ7lk2
MBUVI3FB0tJt1f2AQtZECcP3ImdYnpr7ZIVusQRsoTGo7D58mvhHBMeRZiLWl/pVr/KMbEmyfLN0
CUrwtMfr64fVzcSTMNStLZneH0SaFmP34p06XUOJMoNZvoCP8WtBK1lIdbpdnm1Z+NE2k3amnJLh
wRsZD46EfTt/g0Io17XnTlscZ5xKIFDOvxROPGgN76pgKevy0DtXSMA62Ji/KRT3XDWlQRB2LvBX
I2U6MwLGAfPsPn98c95+9IR0baz14vaGOjRrnVHucOgOwvjMZFplisjY2y7OPlSIa/EWQUC1QKTk
ZE/pL8QElQOanZXuV4wm8L1gQXyvklkbZicyHEG3z6BJ7QLdaxV9BQSKQ8m3DDX7lI59moUwgssR
uujls/vignjPdiPN/IFfhevdV2Vh8Kt8qzLreSrIkfNjXP3z5IAa6A+PMizkmB5XtQejHjj4clET
W069o3RYdTr82ZTqNsg8vgaHF6wABqwIvBizMOaxNC3fZguyHNUY5H3WNi2tpheynRQ69/WpHlGU
+rQOQfjAVayRf9R3Du0JAJpRh8g1x2Md/2lUkkgd67iqDdB3Vvws7VnkwKh06K+cn5Jmb4mUWUgw
keuT1iQg8YNLli7s2J8aFJlC9swXPh+FDakn9QaAB1umFh/3k38rAzD7+UWAxz0e6k0T9DmLIq8Y
zaA0nN9/azwejNiqZC3dRl7T/v81Umlq126ghrsxFD8VH1zDYR6tcONfUK1WQGBIzXZNLlUbUyw/
xehIt540abRdjnYo1d75KLgfYnKXdvKJugMRYA1vlGc1WMUzPJJxqq17I7V5hofPFJs9PRo7w6Vp
r1TTiIoDMUBZFulB+Bmij0R8RDQ6/mbxLw5wP+dt0bRXYZRJWrbW7afapoT/LlNzvX9VxLWd3WXX
VPDmTbOOTO2lQ3Ckt4lrRbfo4BuBdY4wZKTiGlqGo0xrnm+QrhAEjthNe6SLv7xsWpIC24GqAIBa
QlHNV4dYkShlO3BeiL7bOXyeaXNCp6c78enrdnbB28oZriZbmSuXYHeZoo4DpaXilxIW1/qmw0gh
hCP+VYKRy2PzSXe2sW2z0t9fbUdn7zl5+AU5cOYgI3A9xDu+BHKL3kCenhhlAvKnDBxy0tYkBIfQ
drbSZmpKUcU1w9QdR+/6+iKfTsJR8DkW63phfNp2jfRDGkA3kvWa2uYmnzn5CCS4E9g9VydcZ4hb
bjZNZN+EokWB3WH6C8JFmgVm5dOTKyukFJ/imoinalRFhL3lSVH0VbvVrBH/xHjNG7LMeiQy8tL+
h+q5qCN/ukwkRatvW3nX7gy12POI+JuVEBCQnilT8BX8xmxJm2Jr1cfi7mutO8cpY0dA7xeWovqc
jfdgKV8KYT9WR7WbDT1wRNPTpt853BqFkz0jrn4jvBp+pmidzDus26PV3NoYLQD/p3TZGb7HouYy
RVUTBsLjKq2vaKlQX7/zWeOGyftR3/R2ZU5g2mNFuYM3OPSPP3TJ6hXm7BMdqSoVYQKEucwDyc/3
2e0/HWzZCcy20MfpM9JexK4Ogi0tlatgZEAmk+uJ7e1VS3rWvbYqDZo2m5guUrvrVvgUv5XH69HT
UtFsxR5QJudK1t0rLse/gJ8V+0kQiOvRsXSwJRzFkFng9RUyJmKFkJbuyMfTaYX5dpEiOKX0v2Xu
n8BCfhsmh38I9ipY/ViL8kvlgpxDRNhxPZpNw2KcmX/jcDJyvaQFLKrvBggXKkcnm01CMdfAzub1
kj7RzBAePUoUve0ujpf1GT1W1hGSu/ESdZU+hh18DvE8nZTR5GtgLVf5BeusG6iSPegPZAxOpyIH
qGYHvmpxm2t++Q8TsLjkufdTOm9CL1Kgvj4MtvCyHzlVkD9hCzLauIS1Mnvd7fy1L4fKdHSvagNg
i1lFsJ0w6PaqYcl7QJTgj9IDz0uMnsS3+TF0Rgyu2mGYUTZSRV3tARlv0nmNmjaxTVvqC2cl98YD
AdbCI8PqHaVxFaThWxnBw3QsGqOf03If992cTYa+GLXvV6jS54eE+NJ+MEehsGfd3/dM3QUMYB9k
E99qbs45A9XWux8/s8f+35ONM69bmBQL7oP9yaQ5Pdi5Cump4mV42nT//YWbX8jBPzeHkGhI32HR
gHLni0+X+cx2QdY9JzaJVim+V06ZvpeV+KguVGFokmZo1k5PsKrisiCZntEdZzNiVsKX9pjSYOmt
3vxywKxqaXvWtiBD+8wWnvYYKXe42u6G0sOv+OTkehnFLPyTmu0mZv4Bl/+BVdXzDcxYf4ypZz3t
NNdKhA3cNvCP1biNQehn+JnRC8PMSvCk6ECL1X7ItAX7XUKXtdceMWfsRRMX8ip36y2rYHloIQIo
O7fS92vo4gZyo/Qmv75KS6eXcSiJf/NLAeKguyC5x8f5HhJG9s5+UP9y0jRFAvenivLPPDQaucEU
ycGG8N3xRuCm9v7pfp/0ILAZBMvr/5FNkgkKySu/3bsZcQSF5TIBjTxWJBW08rcg5rtTxFw2948J
gOtjXFNFl0TlW6RLFnzWOqLtQ41nY4SQplWzfTn4C0QzYZsC6jbP8yHgh9K8BFrZxxFfXq+ZXN6N
7IrFyRR88cHt+AWN0o2uzEvY93fz0dsSo57dHXy9QkCDjjCuW96k5mzaFJafacdmZAprNEsDnt4u
sXkLYQBVeNBIez4OCUUHwGqyyOLT0ubj3qRMKgKtVgw5ACQt2AlmabtElXxvR40sN4Nold4pFtm5
Y7pOJL4f84B5zWae7FI5Rk1tQsc7FW2dtBTTOjQs4vmDWQlqR4ssrHt66XH2bY1laN1S5N8Es4ZA
nUn0HTj592Gzq1/KaAMedn7lc+H2LoK9Ev+UXE0eQ1iJAXYA86rYQPO3aCcYPtZEyXhFyx25NvFs
+vpFjkjgl4oVZP0feQoS0Vm/RbWcRmdORHk74bkWrA+edjFXtf4GB3In+7QjGS5JUfnn6CFEyym5
zy/Vc/GK+GspIWaedREtLxK0nWnOHgkJn9+MdHlc4H6O/Uk0E0NISvvqPuXibu1gXovav2XsP0w7
aDEgLde0V8nRaFzS2AqYjuRAr46TLQq4RtM0nkwTbMobsgRgqh+YKy0Eemj11wtxfGhywTU6pDwL
Dxounh5Iql6AD13fhPZFHHE7oB4B0N+ZYyV44n1+YtMUBewwQ/MXyl3EOEhgKJlfIS+7k5K9SorF
LR1JvuJQY4olNhtgCSKQGJpHUyr59cEWyz8xhmSi6jk7KqYgAZIjOzUQrpH692SiCdCskrQisEW9
MPNvSjwTunHUd4PwTsr9BqaSPG1ctQfOw5+u2N8lUZpWyCUfCnvRh14IethzSWG6CJ9YZ2Y0paU2
ARRmS2YbPTM+yk4CLMRq0E15vxuJMsnEfopujMaTZMZJN/T5wLjXyRc/Z/f9s9PQIj+1veb7htRh
wMgCbVBzmUutwsKisYgFBdvhXXlOagT62i1IcbHMb28oVjdxmIgVMRAnB/5S+4UbG0363pt1JU5F
gL8tf3AsmGlWTRYA4VKxIZjTN6vRkz4I077R/BLuAK/J58JB+NhrzJEjM4DaC4Le1dJHEyOWKATq
jHYjTPHo9/tez1bHgeU8P9lo2uLEDf/2J/hgR1vVLkfJI8ZEjDkcWlL8fY0Z0XseUtls0rBYos78
UC25J/vKmD0SXQm1INjoJ47y4AbEVPXsmIqVhv/YPWqUm9ngD04GAMsxXfNe1fWTVjTFHHqz3VcN
3OAmAImuvYxnxTIBI3gziXHFdyTXO97FSeMT5F9BjILPUtrJdFsMezNc3J5/CKf5qznY7+L5DXcW
GjV7XqMGCyqFG8o5fiCz9tSus8vgnQ4iUJrYbsQMZlCfcJA7aWRy61EtKU8lffdkj1pLXeUeTRs6
p6nQo9DyGxN7NHJBvQ5rKHBQ7NueD0881L8fYLK7NL2kHKwGojdBwAvpS58U/yOc0tkOdyUbgmej
JFZYUDRqiKteltJVgKSYBD6yaz0Jv/YjmSaBlenxEeeZCHN9U1NJ1FBjV64gBU5r2u7pOCPnolZA
sUoWawSOR0qWGHPK2ezpX5FSzjWRZmpHSClrMY2pU7Mgfv3Nyj8EliRaR147Zr+F+3a0ZZLmTOOB
ox9g2Z1Z38TibxJS6WdNg45rHvnHDkSCWxvepF8VX9Ns+FCWNiPTtdmg2+5B4xyzTHiaQ0mBgBXu
eqHblkSUuAXEqrVDiPN98J75QEslh4O5TYIkqCidIjIFn//50bj42/dekBr+qMFV+7ahVtbNomv+
MkxVlrIj9q1WXALakAsgtSaE3cS6M8lgDB1nzADXWvEGJKRSTpIMrQz4Yhiinh0wx8L9+TmM/+9Q
b2QemwVLRj2SIGZCw9ZLLQXvSDwnnAaB5UsaT+XxwkZrHYPX6LC0I9PpqatxUijNGyRriKcg0A4c
o+F63GSVnj7snLssf78uQM/O/CQZrbQrqUtpgcuMTC8W2mHVwltnwE8bMP5R//Enbvj4U4CvzHqI
Tgq8HaldemQYLmVJgSMiJI4U6j4LMyekAMJ3rKfkz4OV1p5X/FubALmFGrPL4yOefirKHwp5ENv7
+F7eWVtPyHeeNYkJ3R12ezDM+eRoflPy7uBZ9bISuQA7ecPteH7+YWkTEuIH9zza3Dgz5DNmCTA0
7VxJaPtr3/cIDwR7jFqTsGBBWIKKNMZD65nKgazUeuftGr1g1noNx+pjfOUGOv2AUZWpCrq4nD32
Npe69YbI5HI0Deu8fF/OCIw2H3gBxkeF4MKIgkjyEcGEyeH9eJ1DyMvVz7M/lVHhAxC+vxmLOENE
yI3m/ePhzjaRSgiGl6sfvUA89sQrZ+kBkrVnA9KrxRo4W5LgwbvUydLW6/W9jlmVGVtpQLCdc8Tr
mPR82jFIj+hJdn3YZho5dSD+TVNV6NKVQxSrapcedeTS/ooUwtaJTSQQR0YhfoUGNJo/KW9yM4nY
8jPde+mZCtn17f+4JleOlQelqNXJ+GkQXHoELuQrCqMW1UQ3O8EBEcxMO/Yk4Lq5ni2F953LwGh3
BZePZUShbevJIvUjRLrkjJ4uUhGF6NDTWhkOBTbirSMTkO0PqFJXnC0g3h3PnLB0uBosMh/qYZpN
YzFFdMJs+aM3lKxdV/sxn/rb0THb0FRo6KM0KBaQqDUU7trgXeGqyPPb3eUxcWA42GMlHtDijMBT
jnwm0T0hoyXwf+D/14srcIb+Mg9gTkffzuMYT+4GxFKnjW7r0HX7ZKgKYj03qQW3XCJrBJf2fi6X
DZqtMPn3lBcnQWf4WJ7I/Fa885r0LTbq0Z13naGJ5t00Qu8eqRz75U6f47x4HmP6K6eucu63Wqkv
OklKn+2zzbNEKUXi5JjXvgqagHtvINf288que8U/HtR+kclmW44QNLXhlZQtvRfFWLeBMimop0pn
POuK47T/m6JM3ZmqXLojmH3pj5+ZBqmP3pOIgNFt8AA0tN4W+qYXq6kXTyYClCPWqndCkdgsfXQK
NmlqY7w/GW7mabV9+jXid57Bhk9Wv//2NsDC8nrTMeooW43Y1hs7NswGYr/GVrK5wUgATyp+OlWt
7yIsdetMMrPcA6ZO8XMmVXwqeCzDtmQJKDdkgOwZr9SPaCdsybTHArm7ymP568gCci5tzdXoXJbr
B/z71rNqnA+uRNeYYbFrrQFgg6743QMt/rdAw94EoRS9JOnssIe1Vk9NI1lZGp2pQ4qZD9UIAua3
rccclrf4fn1Wq9IAFTzcItGqAfLiUrEEDhTlqrai7LHYQofrZOBRKzf9VHh1wbTkN4Jyh8m74xGG
Izc5xp64H1pqEVMIQMdgw09PfzVkbCisnUafc8woZ2ZOOmMWG37yBqnjoLKdmSdU11FwnUihupJg
om1rwzf8WxhPXq7fqFbVES4BW+aW1c2rEhaDAkiSUp3UvUQ/d2L/xCTwwdCq199aotSbtDHyV7bi
FnLpymRLXj5NdlaPidJuYi0uRoOy90CYG7d5+LMm5rr4tm7Dv1TyHBffcmHQOnrQC3HfSo5ny6j+
/HNQVJ5iFeQ6du44JWpYPTHADQA92Jo5W+TXXJx87iBmDtwPur1IgLQ7Ic/yjoY+tqCwtjom7mjt
43hoJlF7gKwooIRbaIq6Rj1tvd2hNAqOnNbT/Ygfsh9Lu7TkaNO96r1oq5fWkYVYLeOTXJawyPk0
OcSTFm1sL2fruBOEV3LL/r4Qo7KsEoOZQzHriSyWNhnxAtYqRmp7SQrEYAb98iLOu0qHbSiDrzH2
8oWHG2VEcrZx55fXzjDavvAFGIUZs3p1OM0StjJexrj2BPY/BdEqOeKYZB+n297ElabWWff+Swiv
hJnVhc0m+ZVkp4EnPXretEgIf+t1U6QdRxgPmtA2foEIIQyNeJFJjqDR51HsJj+KvZr3MnKJj73s
BIlKzlCNkwEkhG3nHh8CvtwOTPfgxWkg3EPHannS1v4sXXe/hqMUkF+b3M1YNgzB487tFi9/G1dF
XzanSPw9VU7Xfj1JNdgrLLipoF2Hg16GaGCGEpXVrQ8q8CB+rekTXYh2G1IXxJ6aChbpucwV0Woi
KS0J9Kj2KK5k6fUgkbnFo+CgZQWi6adktw9cUDz99GIrEFTev3+OKhprv/9B2dKQA7//CKPCiWca
nUV19hNO22bD6KHUVNOSy3JSKiInM16g6R0f3NVVV1h/7n4jTpU89PgRu4ZUO9EKNubflQuWkqgj
k18lYIJa2wlTlJ9EaHCd6pTd4uxnR08Yd/tsuNEFG9EAd1sdU59hoeJoGv/V5NMotXcFhzlQULQk
tdOmPdGPlg1cMGF0lk0vYPa/r/3DWv4dfochLEvUHscyed5JD74l0LWVshazofVf23wJZn8EeBLV
cDwx4W4op2iExwWgjiQXNVnQTshj8FFCITNR2VD5INBznISa5sZhWFrK4h3Xeq8a+ppTwIuW7Ibz
qmqVjXBhASx641Z0VNoQooKkQT0Qe1nHUSBXDtKuS+Bmfw8i1Qx2Z7DEKDVwsBgjhzr9naV0t1R+
A5hKpt3Hp+xwZ+KkoFU0JWTNKMuhwFTRd4waOzs1FSWu9E1LdmLPAl1H6yoxyLRdWK6wPNQv23z+
t129gjcRz8HZ/PdfQsK9WgA7hA6BSVQBMoI8aWo42EFZD0BFX+0s79y3RT4h72N7wZaU7+t0JNLu
rtbazvgS3yve0yiHKHlrUtfQ+UCQEgKeVr0R8ugVhFNm3VMabnFeLyHDchHMKlwaXlHgJ24RKVw1
GTEdQshkdobnJgrjLZSLj16K58CNO8nXkC1dbzTjKrr4KMUDRBw6yadpMDlFluvrXEwtSkajLvfx
cOnrxv4RRcnuBiGxX1fSExmaZ8aQJnwlwt93AhZ5pDe7O0A/rS8atwljSqBIP9e48uSNxLZ6l9H+
d2vc99agMyr1omIbmAsxYHhbByvhFPE9SufZgEoedjuG8dzig6bn0XDQ4jGo7Bnqf8AUBtYmaC8S
uKoT/8DVXntg+wRPSdwHa2W+0hs0MX6a+QwoAG0tTTKrptsHu7ezfHqm7lmvRWVRG7FzCyMBBQz8
AU7YPBgjB0Rfbj63m9hDOEtF1LuaCQJnIc2OEs/b4YBxzoEfgo4ZWBPkIrAYSYV9aSgbSE9PCMz3
MzxSycI2PJSNtK9iBiooaQcb0PajCP5ycDRlHZ3LaJ5c3DFh0EdxQke/oj8IdlLvfbhCct4VcLQ7
oThvuQQHDoAZeUsSBtHaWRcQgWI1rH6NAgFHHQ2QjH29lPeu5b8vboASejE/TtWUJ3fXTfW09AQz
usUkc/SpliC6GUDcP3Iv8JwsDT6bcpRMp9fL51i8QLp2NuQpNFlOJrJEI4cBrIOAQfJnSk6+dHgH
5R91j5efNjXUUrorOK76tv7ar2H03gXlbQAp7UKwl554Kh4rCNtIibfU/bXAHF7a/DqJDH1A3PWP
EBDch44XhaVIigdASLq6p8AuLltYfg6XVXwSXC7WmmWeRjpkk3Nidjb5waxcfnFBGuPB9+RrtNWX
UIldhWY7zGySyvyW0dHqDCE7YcFrLknsV9enMQsR6pGLAmiKLNFr361c7yiHB/H9QbiJ0+x97yJL
AgxA95TY8mbNKiMzag3eBUGtKaxfDANsoWORukOq/QToOy3epWnsqRbFjWUyJndf2zP+vuQgx5mB
LsV7fE88RvyRcE87+AdygaWIlq1NNIxcE15t4mOfCCrUIW9g5bM1KoRgKqMnpcQuTWoYVV7ljG9Y
vl/aGPwWZ1+XUydyKKqtSsdYZbSS1nbNnsXWWJMnZwf6YvHZIPexslxxetAv2kknVRKeaOk8iHqC
fWReet3ZGzqW880PabmYGZ1aHDZqn5TlEe+1B6Wz5aiv/zOvhvwgdv8KfOtUboU72ZK/C5gAtScP
1nP2EiaXD4JrBdjjGxhqYiL916j1f5akrXtj6XwzdnxiMNaQxxaUKzIovAGFgIuFWdSXSUHSPL0I
Mt1QunWrpIVWay3rdUhWYRgPNnyJ5cBf660sYfgPDjG8bjyNm49Zn2VuXH//bWdneQRwioOezTD6
/tbLGHpM2do0zUomjnS0OnMYWp0X2yWbg8vZnmKpb4lexq7pZT/OUAcyfHMA8FrWsFjGfmRRXOkt
T+uM8YXwM1JH6EVO9XiDWSPRC2gVURBRHiUqKbd1PP3DvpchNTvwXRutzkHnSbhdgd7r7yxm0lRU
89znuLzTue1UgJf0KKFockveDuDBFDb0X6uU1azIV96jLSw7oYDQRoagkleB8XQzZ1Y5PyZbGZms
aQfI41gPoH0n0U6m9oW4Jbbs33IxkkcwBArx2N0fqCtASU408fMx3ISnGy62oUrWjJM9d0nWkJNm
cF7BaTEnGOkjrIwif7ZD9fjhHUWwOYqmNnCbMFlrXwPUF9XChU6fblHndIKLUYZrOkbn5PIWywe7
pj/JCOLDzFqc+QQaF+mnPQ8wYn3sxFw7qC4SgwhBJETgmbcVTJ4zRJC6ziMOwlQ46w3//HH9roOz
opNcoHPp9nfNhV4A7v3npoBdy3dMclLMlvEkIwSq92DJL7HlYjL0Ul9nNdawCyh/JyoVbCyLg6M5
5ls3pycB4Xu7qwUSuuNXP7MoeKkEB/mLIQWa82M0zC9uqZYCY3watWwTuqyPtSaoevzsMKDEm4LL
WoFDjGSRTyNnpN+3NvSR96ti+1jcVz6cwOAZsxbepFYHvmnjCrlhwOftH37GYJQHnKFITNh6qTWR
ZpnZvMJOS36TyaC8UAwcCkqJYMrWSR4oo5HohAX4EjtyobwYqGiJ25lVm6HQyBqv42xTkRjmByaE
iexoOx5wgdNLtWP1OfhSrMQOhN9lQZSOaJn4BNr6DtrCRIJ2veTR8VD51hdeGMREL3+TglaYoek7
vWTTPgpHbXD6dm/QUZ8sYpMK7G443zJBLxZBaQZx8+XAdhA8ZctXFmH6Jkdg2VU57R9Vk3Dejx+Z
+TBSzgtBlrjtBA+9YFvgFxrHBp2emSYAoBnqI3ZpVhtj3+m7zu82v3WTK3rxGHjtGyNqDvcuHo/D
X8Y7+9pJllfal8nsWlRrU/b2h0/YgfAkzHxaI/TEmz0p20YUd+TJQk3gU9e6ojBthtnyIREiZfkh
RE/sqsR2J82PiDrYTL8rfZBliAxN3OLiAdyTdjXXcxAQY+m4v0IVBDdXbD3mLxC8V9upGGC9ymXJ
ywi0Gky1Wi6iubTWyG2gDiReSYXPyhoIIFUn4GDE32L0+OAVM/RrDLL1iUG47XoNk5St2altPU7I
Wpmr9UJR8LbufW51BmXyV+otdenS09X5OXNRQayrDeCvrDWTt+LYL/+D4kT1TeZTL0jpB5oD7KV7
+iTdv5eW1V+5fHGskaSKpDzjIDOh20wlONwt+6mrc/AODQpOufFRLTZBBrCSjtSkGWy42C5Kthp2
HSHsJCrH2YWkEBjIii61U2Tf2DxfPrMruw6eLrHbbiFAb0mq9XeXRZ8Z9J7TqmENaAC5Ck1seObY
u1KgNtzOVPbmG7UM47ZlWfrfnFcGMUMhSH0BwUVR2dit4ljE8wB7YZt9OJTzZxXc20eTGomPs1oR
8nlbEdRgv5zb9+KFDTx7AHS7THyFdoxYPV+VKMJaA9+qrmKJgh3AW/OqXKWoSpLVfumlnAjj0Y8Z
iV6bdU36trs6Guyyp7YldPMcbQnWWQTRdPyDFrYYosV7K/tSlIrB0w4Y37ae0WjmWiRFYCDvuaaC
qZP0WVns8Sc93ed0x2LZrT1rv/rmyMm1gm3iXN8ojqxsTqLqd8MGM0CROioq08yFK1cSfLsOtQ7u
wAPsQ1UBuEBD/nu82rALc0wX3ig69A3S83ocmMhXnjjrphon65OeBxw5SjVheDCAoB/5z85EZPNO
vBTb5HKHr3bqwd/EzRtQlLS+HEgXJvNd0TaFcMYiuTZPfqIbHGLzIQRjz0uhCao/CO+gguHIwwXF
4d2mcrnhBCy638oRIuEGMUZnN3Yqynu8Q43ntQUf9EHQ72RTzj870HuB/F5T9Wt7bwMpYuutAM9T
1Olm+z7tLM7hcNrGSchIk3bOAgh/LuVX4FYQ7DjqrQVvPjJnSnrsQ9t+rnHA0VQ7wuNPBnOI7dIg
7Kh5QnxQvqMOlxv1EW1cDPTOf/JKdwy6L3JLxpL0JAJ8h0OGYgBMrahuOgwNnNpmDefIWb0Yi53Z
tQThMs3B9NdUI51MWi61WZHPkXL6q1kWJKrgW5Eu+M1TqgihiU7fBhE2CgB3w/dfLVrok7lvlSe3
LkRcODIyc9ISyIB8Clv7OoRGShfflrSQ2nVvQgfKtmo8CVwQdVG05vOWwm2qSd3Z4dR2MV5lJmVt
66csEO1bX35bxEM1ph4OkKWXAYTO9KnE7v0gwsG7bjnrxjBQ5pDrkEaTQSCUSTxKF7SQA4UNw4R2
nBY3R+zxyv4DW//4Vp1woGvFLh1iBFizob4zwPhDoQs9ESH2yYp1ERJ0StJe8+RSkTFz6ad+WnjR
esEGabOsegdPy5mwIaEAdBi5uNRwH3PICemjDH9n9LTQ2qkRl6/RvMtB1CloH85g38jg9nu2jSPp
cpnUMtAhHFCbjBCeu8FlYcB5/ttX76NItSIdUVt4xp/23jPvmiAc/ftlHK51vesO/xiVSUAVoE+A
OrjPTH11TbZm1qTd3lVPd64H4e7nKP8ozeNlssRCzTvaKVcAAx+ZvnA0/obLpzo8xD4+SzSoEUTb
Y3iLPexgLkz8b2vKPF/BlWcPgChadRLGfwEw8L9wumiOLYMO/f0X6rxlYwBXYATOzTqympBSH3Lx
aUyd+LRjRA5IPmGCx9QU+FAYcOCQLhRt2+aLFyXcRBk7E3JcCHrqcViIjwhif1ioel4Dotlaggnq
2zCuyKPJBQ9qt2FLz8tQLjchptcPfXRUGy9rWOMKw5saBtRDxdUOTwZXrV+2Ppka+eGmw+gREWWi
2ulUYXvoL/U4Os+4AgQNV7R37bkydurj9OewQiBSPYzz4UJ3T+xck3HYO4GaNA7/lYBXJXa5Ji4s
NxmzYjzAoKR1jELLGAn6yY7QhAuf+SyXf5M93ZnM8js5WMG5J5QG4jU1OhRik1xzX5PFgikO7FJI
7KvNez34iH7qDRjRdSRbGdYZyWOuqcECzW6YzOBGDYIXE3PQ8/PwfZWRZh09OSSuPjPGMkx1QMe1
0gCVDBtQfIiaVSf1xGS/k5iFJArLfIT4iC3OEYBg9r5udqYqnftfF5KH1ESrzIfWoqQ4xiTbJ6iS
GQLidqPBR8KKhGrBM+XkC4B+HCuS0zMViSizJO1vm75tR76McUrh4jJ4E7DxTZhXlctJilkw/KXf
XpwQbuT4giuOfSlsypF3m+83yeYaW+yE8liQCaAXkDVGAa37GcSzzL34hGFnTtJnhsboW+aBJC/e
1r9hk63dfK8e4SG+scNOt2aO86ECR0DcJKdeWQQxIoEXPv8m/hCiE3yGEy2qA9x44DgJJ0hOBOJE
apDFAZVDeQjEET1FbRfiVNmXdxhlsxc3eb0gtoMh0n9mLrq2CD+Q3xdaAJBZBGqmeXh/MMrVVxqV
LFTmIFVLOGShG/B/a25YtKogCZ0LpA3XoHsMXK2Q5gF0NDAog2e9kqZKYIOktRn1vgEKaCqVBdKJ
Den6o4Z21AoLfYqIOSxkHTZdQP1z1II7ZrwJ2EzjPs3w3x5NaTd5ATffw4N1h6S/og8bogK5LHne
OzKKMwR+PwsNC/myHdOCWzjHUVJGm+fbj5EB/wgukY0UXQ0Thu39FT4cnSAkD0xNusBZztVBwa+/
3ZmsPfOiZwWm0yW4O9fS5OwSrtPRdoAO+TSo8tEUXcO/ZW4+/sXHhW18qpVpaDFqbVpLwBMF9Hyu
CaAstXybSP0ruxGZ1uyZ1s1BcyPAmJ2wzk0a3z5sDy0tCH5lvDSJ4XYuorBNKZKxnL4xX7oP/fRU
ZH9MUrTwuYJoP5/dQo1/p9uzY6QwFJpyiM/GOh3E8xn0e4amI2Caq3SYjPxsLnBl9A61rfgT1ZvB
L1XOP0Fd8kgBy0V4ZP/tJ9Da/ZfgN7Tq1BjGWPuaM1liMqntQ4sP+a7L5w3kck5Y88NtphGvnEet
O9b+e+iTmA2+tC7Tuhdh6du8FaCXyFerPAn1PX8XGC2v5qm+9pzbrnmOx3WB53gGVruibSd2q2il
s2Dldvp6c+om/pGCd1qYG4QDOWpw8ZqyzRK1lu/6cH4gyo4DBQb4YbfN0pjnauirXMAq5zny5LUM
CVPDrl3BcojsqLydpd4ICLX0dCvcugY2hGgQuhPObEWsLD83M7wMVk25kcpwWG/hbQd9EJx5OFVh
vPEN1GrzXeZCX6d/ibfuDC36lwUPzpPvIKAd34UaLbem2vtFQ7Ot1lgw1vSEFUZHOynCrKuw6qzy
T9zFotu0o2UfUpJ7AXIbknJHBfeHY5zneL1PP6DnS4f3MeXf7CTVDzwy554WBcECz2yR5epwQeYJ
NtPobraiHkDn5mpm3RaTKKbH11gsDr7KxnrVQbnlUQN4ADR6UiQz5V27fvaYVMJAWbTqwXBIotLo
8FoYO6/CETjBd5ELNIXjLZLNUc2bIiMm73LK/gEJqKh6Ip/PYUf0Arx4yc3HcWwWy4uTSLlkv6B1
EbCcvNL6IcY+1bgPqg1K5Bp43f/EKJKwAQaQnq4R9U8jUey9CwvMG2EVykjiwCYVUUmgRzXWdqum
u0UEaHodCxzIUa3Eis5H6rhXm3Grg9aQmq/B3E2JJCp63ulgI25QKcUfAQWjOYz71F3LfLlATajM
B2D1FWMXoguvtIbitIFqt6rMEI8frW9yvP2Tdtb3GWppS0AbdXkQ2BpeCrE0fpc2315rJGM8jhKF
1rCJZF056kz5ErgBz1LPrxGdP7xNfCovRJ3KSiUoKI4wD5uyrl0/hjHYGmkoZsMmu+zGcR1FBp4Q
xIfvCC2fTSwA0quMyfuG7ZYP6Dy3PPEp42vVKS1nKLA86c9Hyjz9VK7qPM1fxz71fzKpbC1psFWu
Jt9tOl1I5TDqKPwD7Q2JNWRjUWnfNLniIhYd3ImMIgdtyu8v2lZ+M/kOsmv4qoQkZozFKhu2YDmu
qbjsJqmpK4+AmRKqMh8wj6TMAuSMx8Oidfb1Pb9eUdqrEXO9D9qKx60MQ93v47jwV3dvOVGYqBz5
cSa+yD63bpR1ZaczW+u+hqs4NvlE5RA3qibo/SPhtfxhRBnjZzuYi3kJQT6+o9M2rjZPt0BDPR4K
uU+o8+j1eKntiX4X5rrQsQdzHcYTAFA0aCYvJVBNbhYCmWiNQD5y6GSDTka6e4uX3KTLJRU3exmT
7g4kw/Yy+rG9NzQ8nFBZKq0STY3krihpgPQdk5KGQeLoO0M+sXDb5j1mZhZEHke6Mywf1NFXuTlK
OpMcOQ5qFfL5q/yLqE5r9BtNxcFC3EqhPpYKzLduQuJRMA/RgOvj0UVPe9iUqyr2wUj2Vhjjfm12
gZrYS/dIGevPIeZ8EVLjGBImytH9+hFyhL4TAPxenl2Jongutrntg9nIyKGhb7ru5tnqy0XXSrHZ
dyvbqgywQI9yvnAZG+NwNeYd94XcXvDFQdnTFmyZF4uUYNVUCZAfO8OuM3oDD0eKOU2oaOQ2uvJ6
lNIeZ2XWMyHVm21CNkjw04E6X5AOoO4/+QboVu4cUxLnLapIuxp76WMp6KJEj8M7fSV0qK6nbAMO
sXkp0NyZwcohfEPIpkqVVNd/KnfY1SNBfxHfBP/5HBTi/74ULjxFNq+bt37q1yvep23znd1j0mFa
P7qGpOtNSCv05p/9FcYkglMSqy4HkRvQJM7NybvUQHehOKQ94p38X1X1nnTJG5xG94+7PmYFPUpL
fjMfj/STzVvNdTc8K3j2ivkcBuvZwgu+tJt6ajrxWZnQ1cfy3e+7MFAzguJ4V9lU4HtnR5EWPTjs
ErSgu2MT6+TKX2GdYmqqGTsGGiOceAVLLEyx58TWVZ52GpD+Hm/18LPqUJQZKmWFDvhZCCklOWEO
o2PxNyd6Ie1n9zE196w+UVxXrrQaqPOiqLt5knaJDP5nA6jIz13EGFETsSL2/wU30srQLI2nbXrn
z6XYHsIhnVXioS4jw3Oh+FWJZ02j93IPGa7K2Ktz5MD2f54oqFJ/2QDAmSIuy9OWY8yNB08YKR5I
ALKaArYv5MjUyj3l9uVguvU5wA8PhgmhRQTiV9zCsnNTQI/9WTNpsZd/FIdRDShxkg9EFawuAmwE
oeMBHy56o/I/zRj2szHuEWfFGXJvb8TCtsV7t71XExcaJ2Epik5dFE/gH5aFEcQHvkG2qRQ8ZvX2
Qy7ycMj6nQzPVrIOZlkEK8I3rTbjoYEEzkOlisRqTTKPj8L52UC/NA6DmbpPB4F4DZN6+H8uduYl
tDINDaJjrdWYKREfRiVdiHsg/7WgblWJxM8xVPOFOQQeiu4JRbWVjow/s3IqmnyE0G9rh//GvBha
jRoqYNzG1HtS4NcgZWW5Vl3Sc9egmm6myto+3SKvLsErWozAWVFsAaVCPvAi6jk+eyaeAVZpKmnU
egwNX1zw3Z3x0LMl6AXvG+JQ4xR4u/mIPWsWkDmBuU8EjmZuekvtIeKIkgaM96Zw8Ax+Ds/tZyFi
zqawQXyI63wO4FWwiFUApJ9s7o5IXsIn+Wh+KOk4cXtZB2Lg6M86xmaha34MQoNl8WlVFoBepHlq
TX1pVA5jzYfXMf6LnnYfIIqdXp8UdBpSn3Q6CvSLDw9wUrBjXtqtRKbnaLICdixGYvmQxWLIUCdR
IH7YNPGQibfjAoiiiPY38F5JewPpStLxOL9vL5BLVeOG8q8mJEIViH/VbEjT6JPOiNmH9wLW2+9c
avEEdXnk8w1GS2vI2YAzwf751M006evwH/wVvRZBQGQ0iRst/RfNWKKZH718Bgscolz7f3HMwCMs
vlqoK2zq8GOltP/sXfjUMej6SgD8OT6Spq1oOTYA8g6rA3dZd18c9hzDFVgiA5+86VwFXTkBGsGL
XsigeSaNAYLyfAovucZYeLZvsyiqIKUxg1hUtHtKfzd3Kq2OHXHK/SPDsKEUk1iT+exX83KD23pt
LnVDGXfcvezpO79udawojfTUF9PlCePJmzuAukvu7FWGaUsSaMQZpmKK4XIkJLC75bYDHk0DskX1
KX2JvbxhpTXq0LQyY9q7Islv6oX69SM50vqJg+A0ph1UvL4iCBiGAw0dSHYCcZ4JNQTiU/ReUOEX
KeBlAkt9CRoY6zz+DYVYuyqI1Sf8QsxPcuWQ6AdKCfBsLuH5fTkX6Zi441Cjusd0fD+e6RDONzEw
ssoVOKKksO9FmU8y2w320jqr2SjKOGT8GQNr168ycwDz7OAYaKRAuMd2L/RcMy493Hp3InXBoAGh
/tu9aQMIonT/5AE6Mk3SFSrlO67jvnYgfsqIWyFst6vqYxADla/PnYhjfK8iUVvu+QdmLDdsc5ke
UTD6zNYNlQGxtCvtRFf9C1OsZBtIuBX8ehjU1qW6X7by0ugrVofjNnUSAcQS8OMTyIt8xjYHmDxo
pU9Q5mejMySGXkY/n98HcQnt0+TiEUcCMc6Gw6HTDczrUwIFpY+6gh7eA760X744UwgLMiK/hKk9
Q5ApvCkOfI2ljaiVbLs84deuf0Ugp9jkm5DT023ezL/ekXz0ngwmYmGhWJ25EHatNMr04t1HQ8rt
ObcEn63gSIDMJwhqEvr0H2Lu192ZzlpJQxIqxhNL3Z8Ju0kJIKkR6RwXuuyXvrOtwpXz7JnYbxAk
2IbCPMgEL3DwFlKCSrnKix0tyY6pm0clMylBX6b2CBumn3IUyIr1l01u4vixQhSCSvrDWDbzrott
DywTmCn/a5RlhEfZ+xl4GpzAIgYdRFscDPHw4+D0tY/l3TZ+o9nrbAVBtQMzZdc/VEJP9f8AmKFN
0WNvexS9JGJggSIAHdzu2uR87GCUqj90Wa/orr+Y0lMXt4NUjQO8ivR6Qi/jBk9L3JIr2d3z4BbD
x7kP0dl9UM+j8pOhzeF6s9g2Jt71EtHtyACbuF8KdbGNeWAukUYhyOphcyi+QVwXVbS6cSufpM30
eFZwzzkKMbhhb6V0e1RIj6vd6l6pVvLz3dfIvMf0MsUI2KPdM+UUmgL43pu6KeXB8Z07FwwmquqD
DRhuDGC2uG4N6X+9NlnEv89X9JLSdi6M/cdWYFhntfhq6SVCDIyds7ng3I63BQxR0X2DIdeUrB35
pEXZ661tlUw5j2AdeblzwpOWTdNfZJTZuFTQnAyRV0YV8nXAF0jLutoWqntoqc9w9XreXO4u5mpY
ka2xbpRBN+rjwBTVHFF2nlqOO8BZXRorjStMcqkN09drNBQTlFbistyhZwdyzDpOjmEwC/2V4E3e
z9GxVE7DOLTqjL0p0txIKUFo8Fa6k0TvGGm2Yu+YSmFPyM4PnwYAf04zp79f5h6KngAw6oWlyMXL
xwtqjrtkHFXJIStobuPGnp1rLZvN8dwQS10ScKIiqwwYZzEomL9PRAy2h02re2Av4pB1xdrKk+zm
UDGXE2/dN9z8QIu+pq+bqab6eCT5EW/ttNNHdY/M/PEUFSx8V8QbYXKezhW42FDfmiSIfogtljf5
0v/zQJ1Y6BhLt5r2rUv6n7SGc8bDYGjQACaYr4FqbvHRnVjIShmZ/jte2JJ0rYcvp+tu4VIwCUni
itMusbYT+pkLSr8fPM7K1x3cUyGUnKdj0q/JC2G59Su88tuef1wK2jd3BW9KA/dW21qcei6DS3eB
FobhYLUR0LAz3J7OSPgc4vKPtw83MUMNU8hPTv85N7rzkKRxoMQqwPVNxWp8Ma0FWTHQXDWk6oO1
cNzn1SjdkF7hfJYueR/jiIGX9Ka4n0TdGdOtJBerRiNTcQzBFLlRcBf9pob7lWL5CRcPDhU6bsKe
pIUk5ZshkJjujH8NMsPxHzF2awVV38GAnLMpypgW1nrDFZzDNJtwPP7KlzrYOVpMlficzITJU0KU
4G+6EqiD8kuUWoir/nvNhpPXrJbyoke86qDrw95afqejTNJ5sKmDzqyJ5s2yyTC2NlD2APuF+AOF
vtKzgma9v30RTafXByXEnky9gXxNrU6wzqqhvoebQaDd3v9siXry5+2eP73alFEif1SKBYClVyQ2
F22fZyVC5fMmVisru8GkVSsrRp3vZ8AkoC2CWXNtG0/BLaJIyhy2TcAt/V32NAa3PJskGipMRvEh
eDxhWacysdnBQ6/VSJTGEbJJhrwlytfTQO1mZdd7inzAhf1TF/oNUSveIDOUpOL8LcKsIZ5Xv4zb
HJIUg/cTuYNcKbd1C9QcODQGMNtY4TtvNDn+9rLM5VqInY+2CMtPq7V+16sTZ2XK7YEezCBIrskE
V8/CdIhYi6LDr/IYgBkRbsxnVn4jwlDZQN8E57FF6Q9c5OBxUQ7On/BepwkI/HKYqPF2WoxMxucx
hB/AHlW0Be/GJgDpjcAn+8kk0RrQZwYNcbZ6XqzYMTRWYKb8BF77NR503wfrRgw9dwzdMsHiJ7NS
8Gmdv/6BEFNoeJG5YmCP8GfjE6kl851fVTTMl1KBlbIqREnZD0vVUFLq2/MexKkfTaEVkg5me8IM
sJ2kmSM28gpHnb02M1BCne6wt/bL7t8+5wRtixeeInZ9RhXq8uNuEdUuPhqiSar+uMJ8TpSv0cYZ
u/0w6Ogi+j56FtclLHRZhLYJwJ2pB3wJybN4ZTyMue7MhQl3CWRvTjwbqf/PWKqyyqiCRTaybivh
0fhcyQJRlf3xIjHMh/k+TvrT3m+qoadvdoxi81vEz9KuQ3et44qxK6m1WeHz9j4/l6EzHibH8New
Fs+3J/xKjHonbmTTOnWfFn3F86Xx8z0zDiiG4OPNUIanNg8sVfJNIdfkWEkm1/4RVBZjjl67ngYR
J6FK8cGgmegtTE5o/j89YMvLMg+cdwYDIStH5NfdDCMSin8px9WOAs5plvks/pzoMfegfuuNexU4
IPOaR0n4OtRDvsgfT5F2Kpw4KEe7w4BCuemcBsJ8gM7dpB9UQHAHTShJqUjATulk0mj7vOIxckQ8
8WVaqAkuPdsaAwY+zr1ZFjchD60b5W+a8NvobHRhhpsw7SYduEkPg9M27CPLyrk2t8oZM5JA0rqy
GtV/O/tOVIzeVI1KMOIcDi61Tdrtitg3RBC4OT8GAT4M1ex5n3zonsupnGpc1+d/ZPq2rAFGyDLh
qOCppTRR8QuH5a7DBuRM2T5cw15XJJstWVbFmskm9UPyVD7hCf/7yN+tJY/AnMaREVLY7ACQqT2S
I9xfeXKDWN54l8LgYBHdg0+EcdvMNXtyiLlKFA06j0veeSo+XaFglg2iHcNujkcAX+L7g7g8GMPh
0p2XjiIJdSWMnSYdtEAu6mLpNGwYwqmnAzzkzBZ0OSZrDpRKbhyBMrsxU43tU2ftLg/JlJfAnn1y
kV6osARFRTiacV5dzC18m7wuZ4uGR9xVJmbcDhfThSAN7nDhbswMNMqjVJUfitPHmy3OJ+bwzKrQ
0iomCDeVcoO/c6Ieb0pbwYjFmDL8Wl3EAaodLmzDjgcwcLDjmERkEsJOzLL1bOIe8Bl+BnYz7czb
7PBtfI70FMkhG0MH+aYHHkF215KpC5gwj+lZg3hq7HLLIUzjv0136O/G6ukmtK76gu3fjCu0pMWY
NFmRYMjd18Ig13h3AuiN3ZxFhSBErGJxaiEytSkvcV1Y0xPGekM0Hv66gNjINz/hhwzzL9L8aPnU
OLk1bdOejzCrB3px/zAeIP7aKTEkHqNeVw4lYqxrpBtImkXRFRA7mNL9Ivs3dQe3JmcZ+kY7BPqd
BXl+34yQV9F3DP+pzZ8DVrQMBFXCEHqDMIfMnBk1mVmt+JSKveIbKITk7K176OAE29pqP/xFwFab
LVf49o+Id0GB4vbflHYXx+/8tRJVrsig3gdfvb5lSGghSsMd9X7Rt50kw3kgnlOIJtyApsdgKzIE
IgvpeW8JlROD/PSwsZBTp2V0E9NpPoVwtfPUxw3gts9u7/VtnSsnANJF5UuC7QClcWJQ/h6nC0FD
OYoOuyTkubGC7VBx11PAc4sVFaR+hJurdbyuX+xJ/+JcJHq2Db4SowesSJ5fh1scDOEgxLdMYgw0
35CbSNiwY7bQH/p2fQSCNc6yos/eG/NpTfmB41K0wQnf7RfB+Gydf16BB7HpN55FmqjM19uFAiL9
IPXQY3V+LwTSYgTgVmTqHjAUfi6GwhcW9uTkuhDeGQMnaWSeUrm4EBqiZIyBWBNomMzgSdRVFZgz
c8vEcarEGbR5b9B39LJh6SbcpEDsbALErDoMi+HaeabiPcVwOTU1Yz3Htr7Sv66C/NuzAJe/bnNS
B1Exc9DU7BwTUeBYfwPOO/PBbJGuTHBaAFt4owCTxGnpfwRNzyItZViLga9Qo1NAiQtDBAB5r9vb
R4KB9xr43+Z5QUbOWUcJEM0V8ZjZCLQnCe8JzzgykjhAK+78f/Q2+6hHx8YFQa4mxpdozUnlnvAX
LhCXio2OBxN9+cFi0SspFCKuduwbpc4EUZKsV8HJCI0zCZyCOtgJUm848PqMAjQbLdCt00USwDzW
y+wLy7dNejpCV+xLCZ19i+TjSkjD1hSFhFy5frroLzlRM/YjlLRQQw6np1VC6YIyrnxK8lbhWwaF
o6b59o82ozQoUD/Aa1Mixle8F2A0vggUhdr64dsFQHwWwb5VZN+8jKYy87qrqo70iDXa68Wh5YeV
rTaV1jS3Z/EjajPsDP2SYrrmJa60wgGaA21s21y+T3J8/NJpEaeRcOu6ZhwmwjwsByZqTbg0TCvm
yyof8Q23HfNlpIk8MwRAIce5Pk6hTH+syPYbPIDpiEnCs1YF1YpKojVpvBTX1NSItxGCMTVprzQu
W9yn9QTj7B4kHenkkCbrbN3VfLf1o9a7wBtrnU+ktWwjEmqgDDzhF9QzGwmkCZ4MsBm93mzSpd3N
/BiK0/OX980LUwHFtyMC3XgvXx8AljrP0Zk1nPpn0bauriMgJlu4Rm4gTrxFrGp9+Pt3bqn9Eiuf
S3vq3e8iKt7lKveWRe17opF7m4LvFp0+Boq6ZKU8bUsd6/I/BmjrnIHyJmb2GzhhbLkzmdBsz0uF
Tm2mnmcxDgiYYtVS5tcLb3qapQ9etmg0cqyEERKShiscMXiMhryFB2p92o4K26sSoiFi0Pd8BVu0
ZyDGzlqSx+aXPyP9rceEn9nOo5b7Qocym/3tNSnm7m4mKofxAh7Zq9XZc6uSbQT/rKzA+MIuJqI/
DWNnuayijwnnjrPYQiJot2n18+cONp14bhf1EZjEYCGHPs+sdQm3sPAKAv334ZvmJCcKTXo2v/ht
OB1doHAmO0goUFal521TsCfgCq+d/5w1wMfU7WZnAcy/W1CEloT9dY3/O7p1hOncYc5H05u9LY+i
1bqnaR8ODPZxFkAFfLp2HTB9s/CnXf4+jbL6EXkOiQXii3D6lpGf7Ssk1W1Tp8jPU3MFD0CBuqQw
QGBO9h6sQwxRgPS7NL/9GCbEJAckkWF4Mu2ZrNb1RU4qN3KP5E47GZxjJaM785iF07+3VrqhD9GC
ZRGOduX+Hip7EGlI7QbFq7E5+KGiC+Dez41Sbd1y0U1yckPhNQwIpRoRhtdInhwMUwzINnljGwn7
sGFpcxWAO9gxeA6y40tttvyGbzTkZQAEuV9qlXH6uVzHJv4RKZstYsXEfakCPaNQctlBuxsUuyDR
VY6TJKVYbMq4GcO6e2Zwy8fY6AWdeFDTnUtaOYyibSdNTgeOLKpntP2jScJ0SremI2AvG1XMzRTr
SI7mL1DSbF8l9I31Cm2uARK8mspqAussxTqfVArxFKTMl3Avnihx0w3fZu0Kljl9npSpTl7xO5V/
m9ITuArjw2haPNH7o7qlcHdzGI10yWaSLTJpm7VzKHzgbb/yHVczfP+Jdgzpbp9NARmjaMZvEmtd
Or+V/8MmTxCej9Q9pnfQoXktMFGYquOkg8sOUTL7WiasZx4s0tit/d+6YSp2cV8Z/wwN/7q6Qjwu
Kq3W920tEPOAD91BJctELXFo90HJlNnpks4ZGq9zgo75dKZ2uLn4gP7CZwuSEHChdNi/eSpOf1FJ
L+FvXv0oWvyySlonLaaz6l3W/oAuX++tDtD00m7Gt8D5on55iDFM5cyewJ8ZJcRTHj0iRuGrDfC9
WWNL4/UP8sfuD+MKcYLiulXjCphS7Cw6aVC5hL6PePk2QeXS4YApARHXDN4oIUMc2B1loR2A1+Qg
mDuYXIKaK781QZR6h0HSyUhNMpdH2TJz5LiIA7CBBUzCFv7+yzP2aJRplTNBDD9r9jFUuHDa70X5
2Gzpky1aqSrhhkx4c9yxSywvbbEDUc7D00XQ/yOjOq1kq6mhNnw5mgvgOEeg4eGe5TLiuXWb2mFm
9BxTd8UZ3qP2iSJfmuHYqa29IC89Zbvdl20OrS8zDT7yp9ox+LKUX24m7VfNxCnlf2OhDaqNdGaZ
Rr/E8vUWPWAf+pkXnaHp/MrZgjuQvszyFswthsr1sfkFcICpeKtY0DIoLJ5mE3N0f78CNONePj3y
WQBqGgksqjmzx0LFvueisyeO9fIfrpHNFJhG59E6Yyy7MGO5g32nluHAzqtKM5zRbDxbl2KgtFYQ
yUtll5VpEOUsIE/c24ctVm47ybkIPI6o4A+XrO8mLW00VcpQouOcRd0mWPdvfWYVmjJEOCFmQl2E
V45Fca+OGyh9mpp7dX2tD14UUnJmkUSRc5Hbahagugaj7nHtBb6cv2UeSnFWeykVMCBEGRBCDCMR
BgxVh43zc3nkddNmZ71w+1LJUYytrcrhEI+eL15vbi1G17c1i6Q4N4kRPjWL8XLppy70OiYnXDKw
LAC5G8QNf01vn7fIuXuJ51W7jP30aOnHvPY53zae7qH0/p1qYNgC35iVHDY3sXLnb7b0auPidd7k
4o9No+wiJZviHyvvNukXmmJRGjeESIj+rlg9FKkfLXv8/49Hxs5FToylnSBsD6uzm1rcj6Ov80YN
sTe1WKzfp9DVo8uPVTrqf5K5idGgzWp5xgRAowcWt8lQ3cZM3qm4FwAb3sxRvMIZsaAsbHou2LNo
6w/X/jbER45MeT7TGWH5OgKU1LaZmRad5t9B+7HpbgYarWJLORMwlr/v+XkqXTtqz35aqOlmGp5X
M0Jb1RCjrZFB3HdrDg/pITXN/+MjuGBKPKN4SLg3RrI155BBCwipTrrpeEp1vWoUlSXbdXRuSbDB
neTVe40gKjfjkD9wa8DIPR0y7lR7EvRcpugRQywCKrDuVlJJ8s2iWIBlFmP8IxZuc8HBdf+pkumB
jKfhhLmRsEvJQfts8DVIU2waSJBiwKUytVmSUjaQkHEA6PFQg9GOi7ABISviBYeFEaDdWssaPZGb
x5q92tFXYrWbXdPIeGoz35fWsp40eOrKlWoN1h631E3oHl8hlFqWQ9h0ZqLs3YZt3jAVBYvZft1W
FZsqABK5hO5/qmX3vcT3B2Jvgm7gjYkyg3tko7z3F/lcI5ClGO6P11UHuYvPQujwnwdlr3YxblyQ
jLQgpik13Am4IGtibxixLg8WgjG8uQ3k7ZtraVkJscc+JUlKuy6x3EmSYjTlivQCt7FP8HbGmyXc
cny0NCzGMrldgXKUqy7FY8hQiEA5JXgv0JUF05qC2ANcZbdzW/fWmXnB5pt5MbuiOoTinMjfds9Y
vHnvBYIkhF09H68Y35PHorH+xFdbRw+MDON9kNIzKaI5vl5999029qJTWuXpecSjL4Ztbj39e3lV
1eS1Xp8ZwtpyVcSctnHgu+5FtKoXML2JKCt6D0TlDax9UnyAu/Bm6NXCNKHITSXLYoCLkMKZYqhy
VoChReIFemxwawTntYRGkq8LUQcU7yq57oFW7qhoLUfWZjZ6BEyf26xvJZJo+k9zYDsfBxTVE7I1
QWpRYuEUUfSouWy702DDy61+0qkX9Z2N1NloiBtA8wDksD+Of0pbypPBw5Yya148GPHPQmxGPVtI
WaMNUV2b2q6P9/l1nHs7VFLla9HQpuQBilPMhXS2UkKE3VVObJw07wWvEZxqJCv78LQg8c5vdOID
NUaZ08qmJ9cmSx8kuuzYy3QpME56EHnt/wmogLzgwf8bZ5E0byGwM2d6562xhuZ3Dg2J6rAviCGH
5GAfI8fwsACbchOV7tj1ZhF8DbNynE1qjtARqNhRui/VqpK/eCxexj81+gGRcLbgu73No4T4whaJ
AibZccBAP67eMQuEri7Rj0OYS3Wg5Q+urytmYDgAIhr6r/1+9asGAxxDMDPzAK3Ei9fjXYa62uJB
dE5cg+WhSRSmcVF+AAzJ1pCaN+OKhoOOTk7BodD4PPmUR6mzs0+eC3pIz9focY/IlO0ajAX3WFTB
MlMg//wZ3YC0eWqnMGkHYHoq+MPSxISwGErhG8u44AJ9OK4epj3AXsROTCCJS/U6PKUNJatb+s8f
fKzl6aQhYLuKA70Q2jIDrYaqLHnu3WZW59Fl5CBs9k/l2ZlkTR54rXewxUYj4jz4LWQawEVInPL0
5y1+mFUDPsXgzmW8nEc9SjLPWJXlE3QobUtG3KTYgqsggptXiEqrSK/yiC9DNVg0CoRAjerRPq/b
vTOlVi/RinIlR/z7cr+/yZyeax+5o7IG3qcOjIeNHatDgoc+flrbeDrFTkwKsCUed+S+qlY+YXi6
Gp2Eu40Q7WTxNFVVSYfINwq3qeHRz4NJVjlx6snWqbIL99M92Bp9gk5XY1kHEmeNYFDKjyYGgu+I
DetojbJVKyc0ZXNXohH+cnP/utGSp3IOjg87k965sQyGNyyoYjjKE0iW1VSOo/xlP76ieTvSjKHE
YiXXQH5cZwgbBJPL4tpsoN1B+b2QELT3jeOFtSY4PV444GSFhkvih0MMfjygPTs2odZnaDcX39E7
po7fhj4lVmaD/S7xMrTgT0AknaG9Ve5f0CuZ63M+WpC7XEYbEa2MZw1WlEL0T6M6zN/klXT5kQMl
AT9TxiwUv4fra9fNgdeXkjJ0o3scKdz4YprhFbnfqo6lX/6mlKEDhXmLga0dh/1ujyn8zRmud5eD
BgseKDwCjmgGRSUFK9gzLaaqc+G3CSzt1pDtxLs4PRuyYfa1b4JC32boVXS27fU0cY80EY1u8Qy2
Ov7ER01E9dayn6tXLdF58QxnNKo0A9xbSjROBQ/3bRfMVBpxuJtiDDN0+sYd9IvyJlDNM26efw9u
s8gEiXEm8SsOULrOEyd2uLoT1FQy2hnmsshH11iWRrHQyHch+rakuq23tBNz8ac2cITpLs1C7G2G
NV5/3allYQjLMVX3adeMmuFDrSZWMi8w1Z7S4JVlv3NEjlstLrYt8ENxxA3+K/G2nYvq4DkukfVZ
ohV9fyNCNaL2wByHvy56yeg15VeyuHkGoCdDZeMZ2scBpgf/uX8qUDOdK8Ozu8RWSV4YocdArpvN
KD/5Gxj4dsU1jaTHW6UKnPxl4rQ7KNzuPzzO0cPhMiLnVCUtF5tIimKnlE8Gx33MQqPcGTH3TK4H
lVK9/yfg+MOtHr4dY6FpY08aNU0ENZ6Nk0jRvsCpRcWVrImu+gGaSokEi9s34uaodoils+oirvFd
zMEGFX5hvlkE4GGzeGuZ58maqcf0DsLl/Xt1/k0CG7FWatAeQbLnwnj+KAXbswQVIms/3jNZZtUP
EYAJA06+8aaAZCEpRj53yisroxI1Q9FosuoswcuXgKmBbzMWxUj/+VV2iCwcyuafUqYQFbhbPXMn
+PmbdKhggftTMo95yAE9fvbUtDvcR2PH9s8nfdELdSHZT8p1AV18Lno8oizQq116aNuRx+HLz/Xr
9J0uCF6sKq6GoMC2WHA5UCvRMExqCvGPSYLeg+RQLxXhirT6zN/5YswzVNOHmXtbYvQ9KboBZnzy
eQYo7LLclNBgGGaT6jQt9YWmbrVLx4CRffe9BQF3Fg9TzZV33Y5nqm8JPxZF4Ck2nescF80Tz0w0
YMLz0wgNieemeW+Jtk6AUYZDZ7NsUWtuMRsN8qGeu88HUbM7bR8dEtVOzDk1dbGbhClZlalMRgrA
FIGzxoLrn88sdJzT3hORgvpMXdIaMtPmgTejPcmjnhEyZNHe+0qXH6hsE5uQszR/iRItR90RAWC5
vL+vFhIAq4TAbaRf/7BErRI24nVCqgUplqXWnv5qkaBiHVkcv0I7UkpZ/m/KGpv5rSzR3xxHaTHG
wT3Q/eA2U4crEtU1MQBQ9UAo943LACiMbOoHEMouKBEgPOzqQ1aCROKCDd8MdDoGk3OfyW6lur5p
ltZTap9f0ifuAGebBBCLNXnHOrBjiHH6o6vJxncUsaRF+IEs1XXnchL9l/MhCCHbRARDWcYfQ5zf
5GbQtdp2US3ckqP1DzWU4Zz5zRkAwAnLfMJu2pR0TXr+u9GX+tVWUaSzpshvMHdqgYvPD6/EKZcd
Bok54z8PGHULJMJ7Z+Hv+Lt5gAe6vrfGBJ648G8wbrXDyOZxW5J8dXSe+U+kejjnSqDMvXiDeviT
Kcc4Fh9njlUjFzam+VWV7JiIhrVwRIEScPxQ2lWuwscjKW/rkbybeKu7AdNozm7NmgOEHfWPcRJt
VMe7ehFGL9A8631O9siA1fqVGPqMaLr+VGC9SmrGuwYa5pz7+uwgsUJCYW93mKjTuk5pG0GVexTm
aPX7OuSXCNxuoJAm5ycjCjGzhK1AD6OlD8jGDDSyQ9ttFW0GVvkCInGJJ+iY0EGHCu49d5yrnio+
x8yblrZbMs2xCs3aL7DZZl91LDCJx6wpQvlfaR9SDaT6/6w8jJvEXedXQQHMP5obzXrQZbi0xaz1
1qwhSrMtzAoWtCAkP8XOFofIuV+40rCfUImRhHRbJPvyro5n83FxTiXpCPF7WS5I0GQ7BjhnU5m5
bHerQnbmrMvACeloWpEtgjkMre+G6FLPz9B3jIAt16XH0xZKeBqr9ToV56L6Hc2lRs6vITTNQ4MV
d+hlWobHJ/e0FEpbOsQHdf9UtFu0aGMVhzXXoXoLTMntu/NDbcnBEL30+za/UwxRfITnAKte+InH
jFrh2jzy70uwSvLRHT3o+YazqWW24c9GzFup35zmV1aIOlzE6SQmGYDY/KI4hkVydPsJ+eanS1Z+
Cmp7K1IHwzQLUGvrJxTAJuaNx2qYQt5ITigmOi+kp1VkluMa/acq51to39MhguDUkZgV8oK6ZGu3
4uYeXfvhaJQ8lgm7vTK5lPTtsuGyd0buFssmd8xm5WJxiDYgiRya4azaG/mj3LhYjfUdioPw7vyH
IkiBIeti6Q+6OKsBjCAS1d8kl2hsWeTolGcvQP79V5JBiTUCqTgAcAeUJChnQETcRun5ouGlboMi
kpCXqBgGSM414aOK85xoJfXLUu4KsiB0yknjZK+T0VRa7EeqMvfYhVCha+isr6uy5y10muqlQDHt
NFrejjEUIeS3xTjeHTV01zio9EvChi4ZxyEjFG3kw59rBn3a4ATHuSPM+nVXwAQBTYVxa02afVBZ
rcAFj3jXztlqUynVwDou+yPQZDFDr3dk/ziCViiBPBQcex8ZYZqkcK+AMMmB/Pkmc2Q9XWetQZna
UFbTJPpHW9h635oEoeSypYO+TaGJokv10vG7JY8LmvrvfuzS2h2j0mez/hwS56Ib7g/vKbnxOrul
PSwB5pVkX5+6sbcnCPieY9dX29pBRWX2R4QrE6TXekF5AVwE+7l6chvxNzcn49C3Jebr+vaYsDpH
wwyJK7o/UbRkeic9GoplwTmQBFXG68HHpI5RN+X34+qjMV4Cj/k5yj6S0Ypt4r2JWL1P6mR79OR8
AYp6XrWKG2AOd2piQKQUcaU3weYusK3qCf32dZoFxtPwn9A1iSVgFMiXGY1jvbqeUGqdA6LPboDn
wa5Ila9svKHIBnNw27MwseTBoO6HEEt/nCPTyDLJRz6wjL8dcX9L+yQz/ceqqV9b5HLXOrb7joxa
bI2lXQMV2RTKdOl9y2fm7WWdMDYEI5Rpq8rr9POeQ2kcSXbf+V09ccB3pNMdOHstiJ9PgfdJ/rMQ
RRTZ2A/fIaYPinZ3m5OGQQSBUGocX2TyNmsnCeEQscYkqq9o5cmfQg0JAnYGiLe9rLrjn6I6pUjs
i3gbHomaDej2Fzc9D1uJEkftmVmo4Vek9SQ7UzwbfqJlL9oRyzoQl4eXK1oBlBgAHSSExbisJIJb
FDnookGQxQwt/Z4Hi8Y7b8x+qHv3iSXrnR684xhaW3k0kIE4ME3Jnx2ksl7FwMbpXKOq/W2Tiuo0
GKdjXOPQHuspSKuxGaLUE7UTjsVe655pJ9wwMLluEKNzA4RyI+lgXnS/q+XPRL8YYTjc9MfwyQkm
NG8XFAVqyxBgl/+0t8PFf8xDFbyQE+OLKB2J/9jjUvODN7gBDjdbtUQqrW0pw2e6B0LkmEbyYerl
8YU+0CTVbVpUaN+AR+PXr9b2mrwsxLd7Ehu2Axe/bOMsmvY2JuvfcYKzWPtgz+AJAysKmIUGlMru
tZ3Ufr1jljZf/W01fXcYwdLXjHso0Ywyk3Czs4sPHxgUPBSMSx0+KcX7HcyMntTsvQ6sNBiDbgEu
bNVlz2ENUlNcV0Xd3VbPekC6898OGeI/6V+pyitVDwj8IuA2G+RQZxBPoD1YKH2zGmR/ktzPXqAS
HlGXAHtA/ruc4IHZW3U5M59lp5O2t2lxPM8cDKPYKW9fYotiGppGfld7h+P3R0HVHgFEgLBcI4EI
ApcJXOqgxlLK2Stdl+1KsQzjzh+dv1MuFI/qk6RaPXgUp49JhRNKgvutBDX68/wlvyev44ZNY2v0
RMUIu+/6a59eWZoGa4NvTwvmvJMtXi5quK6q1VADVUikSUnHFeCQkHdl1NQ0RPF5ARYxZ26/ughW
jtGFGMEWSoDWFTIPboy0+iqtPrsOdasOArMN6tRWdJ/0kMYs/Qe6uC2uiOgtA3kqdJaLPxQiSb+5
TZKwbydSJKUTLa/T+54gxjDPFq7v4Pocx47KRW5xQ5Gi1feIdV0gs+nR5kk3FUlLXxkMo4gnpVp9
c4mlOBST2UTpOATUvKQaE1e9blzNaZhTwRX3y68YWd2TRev5NW3m3YQWI1sxZqqBbQJD7AgsXAuB
xop9iBSjQAC70IhtOtc97x9qs70D20cANJFVHF0+/7vfx0J4WtJuiBUY1hKUhIQ82GEsZ3xdYeeW
GZ0DgBl6uEwGx5zaTSBw+FZXvU67X258VhKw3USCpmwIuoFX6QSu7mN8by5L+77DoJriCSg+StMc
VOVJXIy1U5gzz955borZmT8RpgnZiFaZr+fxZgLwCWI6KvbuPq58u7qnYeaBHQP+bH/K/yQ9utyp
swt8wiZzt1ECPQCp1Zyk2E5i7+DsMxY12ugBx+5l2ZS8L5c5zji/rZmAvAHdWSEIQ+TcjNUuVBLK
DkuUSZOAnskq0hSNFCFZkEsNPvqkEeNmlueV3/0Y190a98AUTMyolpsJdcauqnZltjJDkWIq1//6
RM7E2mOdKkJPF4PU9QVy7YaFSNDfkuOxa1zLT5vUno58AvsE2BpdIl43Y9JjuwHS9m4u3DPrOQE1
Uzbrx2/RHcJ2DFfsDnYOfBZ8aJififrk1W4bBH+3t+CY++DDU/+yGq1/LFujElI6uVyOxDNl6UW6
W6UoCkPgwqbW+Wprmvsdxii5/pnOuu65WUv9E1Eto8jiYT5o+xvzzXm9RrDyv7xyt/9y4cEh4GVa
CM0M2E7XNx6qcdVTEN3FPjbzItDfgOrYBP3Mf8XjAEkuPJZSH5nFofBt9LjjsnqRTc/hG+a9DhTC
6WNMdFJBqRPxJ/fiJZMB7VxUpS8h+qmlzlK14iZhys5IwLvJ8LGTMgdhLN+BT0A9fY6GUvKdmX13
z0+e48dQ4XWs89Hk4etCtpQpPMvH03YDansu/KmireTsR7uUv+RGIa3uVvYPbTmGLrPQLrEFInEk
vFjWNO4YHQKZIY4YACmq966UEJiGxLCeWvmLVXlQl7o3c4ooyZtyW7MrG8focwbIyAMyTWabc9oy
6d+7zVrZb2Xw3BkWgli6swnhtqojjcPuW1VufZXewq9PfOQ3RO49i1/NkBtInXCf1sXqc8A2FxFB
HJB8of3+2E/asQHJO8mTiriGq62LnbT1M2kFeui6xa/fXfWo9p3OUFsh+kYltCxPNHxQkpWxKSkT
Z46QNJ37cfzUXHCs0eVeMGYPOWMlPWSvlmGC2m0V8zH+jOqCUd3GFub6cBMsB2CevlUEvytEM7SV
mavtsoHsICG4L43hYb9uN+7POXeDHNpbtOZwHNuCIqdbhgDZkHpyj49WMHgL5c8z0oDQccTfsGFA
kqILzwBFuH6GIL0c2CHrjQjw68EmGuOH9OIi+Wj0tiyY4+ohECcYP5XG+OWjlLqQg1576eldvcHQ
q6XFF9oYrAZfsLHWhEgw5k2fQhWCgFTMGkJyMiEJMhCzMQqjFftEHGSUARqxzNQX7hnIx12ncJVd
CnXhDkJUZA0JlwCgbkdhaWrGWXOjGTkP/km1CKkDQPNQyVyBiLXMksY2JIF/kuXwQUYzUQH+yopX
OQfitB/uG12NStcueiLZ7THJAGsqZiCizCJ7x9d90x7nQRuXkoOtCfSLk7NyYw16/yJHbdMIrHQD
8wtq8a6Ggp1lvPNP7H/DjW9eqAALJgnc1TE+CAIZ3wzhvw/scHIXG/jP+wDc8geYHfxDVW1wvMNF
zsIUlPLgvNpado9metykvH1au7NWPGSjS7rDXr9+2qY1zVXjtD/54CjNy1mZmAJWZ17YwimIm6CG
wF7OqHVBo6RiiRng5lTklCNAwpXH4sPyXVint1zdcS2ArCOs+tPPEF0zugGVuCmGUAnDNX26mL2f
a9OkRSzuVRvXv/qY6TR8P7n8QruG6/76nRkcaIlyPMKfyyu2J1z7gCi1Ze+uRJ7Z+zU9hpuHHi9l
BHtvrA1IKWjvlSLgeXId0E7gc6CMaTVYWSBF2l15VbXw2wtTnKleakwfr3N1VTUpJyyQPZSY49V1
goOR7du2Qaj79catoNxnFMYA5oyIraD5TA7iWkbS0mxrJy0QGeTRyeqd92RCDbFwZK1CwYGQd0IC
w/JrMArl/0jnw+I/oSgpasoX37VUi9n3q+Wr59EgMc1cNmAzXbjX6a7Gza6ScC4xVS0QQHB3Pv3E
Gavxluco0whqZ3/Oa1AknMIiOq8T9K3tJkdGgLL1R4vg4j1pt1Lq6CWRMoky88TASx12dw2t7o1Z
bDrJfBT665fxkOfwaUW6JUuzvSpdY9etcg+or2eFtMOxt3xIZokqIaD3tRa5N7g1+FSq4ScKWbhz
r1J50e6ZpLRH08qMfZSZKA5y73RO7A6jWTWQh0039FxDvTr0nGu+LJB21Wh2c98f4ZDIiIH+UpeU
vMajtBu1kMjtZlCA9QK77QHusiif2mHaGe8z/SFwErMo+tpxrpZNvaQ1XtaD1MrNHfeXKZQsBsGU
qN2u3kMCPjrsAl4YuXU9x+VqzGRSjQaVqGKcAhHFTUAmw5a7qRrGqTHbGW4w/xNGWb2kZBQipaQk
zlbwnIDCf/EbmNMTErHUf8lyNjgf0yvl/09swpheeyTuyXFW2POKO4jb1yJ25m30nbEe7VxrZWvb
5NyGJyMP61zYUqh7OlgXlQNedCAhLxC8CVlBv90UXTcEARXPeccVPbQz/67ZpJl6pqc+MbTaVjls
FoDYdjOwMYnvOsWg+xBWgM9dp6w2HWbzhdYj7z68xMZLN/dU0QC1dLDE0lBoHiMfBhu3f9owPpmT
POIj5W4+zoNZhvt3OM4OiviLqNrlSBv7jObPHPAyBDc7Veb68rHK6Fr0S6HCVFuQmEGmP2Wmnz/Q
3L2skypDxIfltkgg88XJNjLSDL01+RQrvdL6pzba1IUbk8CTzmblirNjN85UdEi3OTsxpezewG3X
uW6DtnimIDsxmD4Qyjyxs08LwOfJPvgNj/nIjLYCTPuKJNB90xl1RIEOMrREwO5RcJH/BMgLb0bU
ouCaI/y7thM9K088qdKnSsO3floyfs/164+fFWUsV3/J+5ZBxFQIKpTtXnToZ98WJtyMCe0l1U6v
sPZwWxODq7DipcSh2NAjGUjxwIg7bN292rPveFeuvXvIPqjLkiI+9Ta6TMj3zpJNMbHfiMBl8m3l
+J7FBSU+dTxBgqBpuQ/mJZ7ziMlQsueM6brG5XaQDnxGd3mpK9rGY7grWO7Y+9hYvlf9wlBRyO5i
OheemlRDWad/D0rK765UgHQxbD9H5bIIkbjOoh4oKHh2bXOKkn+oX+lMAnAiL8Wsz7SejubJjz2B
WqH5xUrft1amX+T4PYi4mLH/zmHztbA+Svd+FmY/v4cEPNIYoPW0hlOTGe4+Pe2CBeVbwwale5d3
DzYzqj9fTbfFTq2rb13fhqBduQ9y76jZL/qc/52jrGTfn5ZxPMMkd5q5hyEM35505Jc7Op7OMIQu
jifBpY5SQjUNrYRxKXUHLKwLbFA3oTsHw82mPUkLUu8Bcgnmz//rGqZuqwnMMi3MFLbBWogiLms2
kZkcX6knTfC8ZhB3S9ORHsBNWafXrpK0nFzBiiM0zOpvE9Ra4Ggor85XR5Nj/Z7jvjQaSVQbinPA
Oqa5UFyEEMx8RjUPgRx8FIVmxPHHcqNkVQq7EaqWQG7rE7pFUzo50gZNK2WOB0/u+4RE2mGBYwDs
YqspnF3X9kMatz11c4M4KokJUhFcv9YOL+nZ9JMTCXJZlpuTBfh2jEpnYqy3Slv7NnjnrjusZ5yf
tM1T1CuXfLg15jiwoGtcoSLIvyaifFKLFVoHjT4HufMUk8+KlXEuEHk1t2tkcyRoK10NNTsFQls3
KIy0Bcgo7Iw7aLQjgdW5JxN0JqMJxFcbU95GkEBgk/9JxrL7rGEmU9R8mKcvTZBq5VIOgB5ZQUYR
tti9EoiI4lWdeGnUYr9qLy6PtrvUj8FaZvrz4YMqwJTnXPt9px27gukO2u7EpOyNS1JJLWoJxN7f
3Qyp6x2EzSLCJ7JFi3tMtTE2tNKLsOQ/v1bjMDqHYI54sPI+d1RNmHZ+A3PBdgrRM1C2nbYqxaeR
gFaytBZ2gxJlkXgxjbzkVP+j2zbSlDFCSx0jwFGI4xNzV7BeqoTrTaL/ew4CWxO2k1UBl/GT/R+D
sM3+tTZdP2TcNpuBshr4l5bPGcc3jkNCoFzfM12FbgUMt/nqgDqaIhc0vEMLcwRO3RKO7f4G7Nwq
PvckMgWt8vmy4CofEtKCDHwOeXm7VHrr6ETBDhgrapbmOMc6JEseeZgm7UZmpNRaErp05GaFy6Q/
M7pyw35XpinQZ/4CeDw4UGGJjNPNuvzd4AHjatB1uGDgelmLv+B4JwkyCJGx8M51CqnNMEOD8e7z
OSEiRaUCL2SAziNYQkAQMm2x07IlD9AGWT2LOHBKLKLHB2uMxgQfFUiCBDO4xiRG1NhC+wa3qG4q
L4QKeGz0vRdodTwqKIm8XQbEZqosOnbNRqumFr3F+AcuBiVCLVCNKcH/TvJIxFVT/bm+PBF/UXxi
tDzbntJy87sAX6YjkXo/1Fk1ybwWOFCIKdFrpSf47ak3uL0El/VJ/eRcKuvvvtaDq4UTsZiZZT8/
fzeisyLFC7j+x9dLiRs75y1Jh9pAC5/AxLuvONhzfrp5MhEBLmobxXeOn3I49eTFHlFsaEqgi+Ci
s0wSbJE+H3hFzMONmblG1gONV1cAka4LY5e3gGcbTzcu+sXrn9EmSsKV9Up62CBvaA+1tAwoHB4s
dr1U3CDmlBhXqF9Fnoiinupn/ermii26/sSj/RFCa2GUgHwgMklbJSVWbfD9t1gw2wHwG1EScCaG
5WslsLDhkf9iKbccCbekZzSIzoB/vqfWQatQMnHJG7M7Y4qOOqmr0WY+yRc6jdyubgzOinOeJjUw
SQjbyi92bXvMkrObikHJzLfa9OVcVzFJbfbBKXGiA4IO9eXxiGjCYFsh6rSF74D/bx844r+GQif9
tBA4UofsB+qW30wo0B8gWzhUMGUNFW0T2+ZZ3bSi2sI3xFwHVlWiSSEpfHq89phW44S+2Z6beMki
KSLbx/7FbaGgpGNjisE+iGR6ilQm30qEBDX/8fusAJuQd/5UZAzhs8elBLSbEYxgu8JCHh43P5O8
RqCOPmwO0+Cv3jup+dU8mAz9sxlG16GivawToJU/XZqAKDwAGlAr69AaNjG2eMmzG5FVk5iXzuni
R0th2ar/70UYQZnOdrDfGByAxlDyjSManzlvBzCVj3sGhA01+PmWQZ3ogKuOYacKOnegYxyVJuCv
lA+3aHObFQ3UK74Nq/0w6PN8dy0xwv3bKwhWDSqjxI7lBdDRSYp+tPW0bSeEF5VmtMn2uM1iPzWs
gqpVFJl1Nwjs1LXY86JNxp9jxCduTmbMmOQwvdt5lS8Fft8IQr584+7kPVl5xtjUJVY27SsazFrS
ppU3TnmcYUa10IQjmyVDEA0vuLYDJpQTnx6TqbhsoeBzPR0sYw8+pxYbir8rbHDKW9poV5u3FBTO
eXoFye5S05mos3ld57SdtpAZsYKHcqMhNAYeDSnFIJLoqHBt35zjELdcEKLA4w+5QVB13HvDXGl+
CvPEKcoLURA4KxZSICgpBQs79J42d665snaDfvQh/POJ0go07BjuwwcWqTBjt4u801B2hOnOgKK9
wj/7OnjvFwg3xHTMh8wq7GC1U616zynTkp1lf1HercHuQeCCjm0NvgkWMCWOVDB2eyeIgU/ovq5H
c9UodqLSDURGeiPgPyVgdwBb9eu5DCALSZzOQU76Hy0BMx6SqnjazSdiey/VKc5PCdYzDPVUxoU5
yY94f3U7X9z+CxfgSy2hcb9FHngNlbrRxBTEDCmXRmcm4xPs0e6fqsBgJcwpRKeXbhfUjcuru6rx
YFjUfUhnw2hhqobjDEqGySQgT3KejPEpvdqz95k0rL5ZtLrUdTOXvBB/YeRQ8S5yYusPejL6eURJ
klyAnnczi/2/RwARcpoNWmT0WYZ9aQ7TwP54rqnxEFjmt2jtY1Ees7jd1Y2oKXh8Z6OSWTEpb2+7
emHswjkEc9Lt3VpSDyE3qdfXbdF5R1qqVp2u85sQ7FEYXJrBEgWtKc31t/D9DMKaEbaVBgPbh8dm
LTv2KdPFc2QQ6V3IbrNZbgjBuXqJ5RCa36wO7rzi/YpkxUMGqMgf3GEAoLpUfF6eYpiD46vVdDSK
z0HRQdWmi5IfNze2MZvQz5bkDcQ0ST5+VvFdONXXVR5bPgN/NnERngc95dbrJ4Oj2fRcX0Z7X6xN
Z51Z+I0QY2vGNgFiKhGjKnPLL0r+Nho2S580eJNptTxXQjNJREuIgbSjKX8++oS4gL/D0WGhP4Ga
DlVZMMrf5cNAgYFnvDcnEE/Bq/d6PSaxH/im4rjOZsQtlEXOftELvZTZcbDIRbklLq6t8oa4PRsl
ApI1LFGi15a0pOlSQktNAfBOnoXvMscgybGbHwqTDLf6urW2O9sVri3LjBnU0CzqdMPAZGwog44U
d1G8e2tKXOsAQzslmYJh0hEpaGFq5G3HYxbyPk9KeAyg1R2Ca+TYY59qGTxPDKzxLD1pzcjcQ3xU
2sRxgOF6AjVy9+hWdGCCPxkzNeG1UJ1TrvU2KcsONzTNAp3aSx3leG9SGZrdr7Ke9cGydKHYfwhk
fXkOewIxn5CMG2PinxEKqkywzSfoqxIfsBRLfoJ5aW9nlVfZVoHA8vZLA2rx/y7M9gOaA5aJ1rjz
RNHXYiDKF9ahVK2cy72xOHt5DIcHJAtom4EkK8xASwqH2EEPrGQAk7KvuOqdSs5zJIrRoN5W9xiL
YpC2bWqyl5gPyvSB2CzgbcihdAPpJHIN6eDNEBxxrIkDbAzBGMmsEztQlYVXHTlifGe+Z91gZFM8
irRJvTCKca22QdpZlZheIHfVHWLK+UyfTl/yIWz8DZcORetfxUbtwsD+tC4pfVW3EqHSgOR0XPGO
JIOvdmOVYLg9pVSdLzgXdGTPlFAbPd3Q+hMEQhbRW06gh+bmGiOclUqSpnQpLTxSpzH8ArQp2byD
9U3LPR/7TBalnXomfxRVZqKQ4Vs0WnvDc3AEj2W9H+Bq3qvpQGJapQ5Dv3rQaxNcJA9UrySDkIo9
g/f+c8q1gf46hqOKomzL7ETqvhw33xTnQoW4H/1x8fSeqWIXJe6RgkOZe/JWmD1yHMOCMbRNTTOn
fDMEfMn5u/ejk11TfYg8Uq+8nhvH6tByah4wRxrzq6QUIsU7wav44mO5TahrrhpT0vKfueIFS8VW
p5Fku2E4z1wmjnwPIJwQGrMoIseHct6TP5Vb5bFeIpRDqaI1e2bl/Bu/qL0FZcTmGUD3M00xZbWF
2ZrZTC7e3ohdSEF+W76566k/ivI+VDNRAMqPqyBKmKCMMoXyTmiYO/lTs2qNZUHxYoBKrocLJztP
BD1vDKtVLzxdDh2zIUlXte0caxdxlzyR+kYJx+X1TZ2tA+LOQzDr1JbsO4n8fvN5GV71mAHJuMCS
jj/u5+lhZQ86SvfaqRE+/bfz9Hqr1XjGbMgtRdnwzKmt/mtwFeHRcqdUFuom3gIjSvNHQYn4JlcK
faRg+Nxlo2H1RsfW5rSHSoD+5Uxm5zhFrc8n4s49xdXSa5+WBb+MUP8RH55vML2hTnVkSU/CJRg/
4+IE4uKTWcWWacbM4w3GYqI25gvl6h3huBNqt1q7n+nJ1N9I7tUJ524oFonfm/8jsYVzVrJ7lyLI
deI5hx2h2IUJvwUUlfSeGWXajHfGQgTW2EktM3yEx46O98qIpmz5viSbRZtkIyKtGYJZBfxERP6h
abpaZSa6v19hWkF+osn8bqv9MAqjqoLMVDJXy7EdpESmscBOw2d4nE7mWsxkIL5uVhMHfIQxd+xb
bfPOOhtNxapZ0GYCW8PfhSn0tLo+UIeVXm1xP22HvEZg8wSvI4Kxsq3FCmP0SVcF3bfQ3gckWzwr
eYKdwmNP+hPFA8xTnvnvaINdI6lUbOVUUZGd8cpzUgQUInb+oWprYH6kDRFBrvsZvwoytgCXo+8F
njIjxPXEoez7I4RTAdFR6ivreuuJsJ/9q4mLWa7bSvhXbhnnyRvq4p9FugXLfT82pPKmQMRNuY34
kuUxgN1zzjhcNtt0v8cV+GKGikRXD7QXm77r0bF12y3z/ir1u48A0e5gkzk/9EJh+remr0ggeYxK
Jfjug/La8IF/oFJmmwMiPKMJsWLcJjbTfg+pY338SYSF1rFIYOa9yWk6o/xLl2eFH62m/7F8xYWP
JAXrh8Lu4IkuivJR5yKxq8LeSccdDJBHOFSWnyr+GoA07TqruVOledjKGZ8pm3yxfIV+t16bakEU
q1osTZYKawu8g6IoyV/nAZ0IRjwl4XumeUTqAmsVZmUuDJRPm7irtdxcY7WW/O8gSjVXhukR8pBF
ZhyeoIgCLgMTH6O2w1GWflXF79U8LAmON5f7NoNbF5OW7rIbG6zwNatQnanmCYbyabAv56/G5+YF
m7Q7lr53kX8S/KtKWBNaUkvTSVlFVC9d5PFXBzmZ+h6y3pzrvCmOj7hJw7NMo7p4bwYET8lE668x
DIrhoO3S5hoHo7WD8HkPnA23K+ucgELN8LAF6yQQujvsYkt3KC+10QVRuEFW7unBToxPOnI5C96B
ZZBQ5LkFOJU1qKRE218iuAjBSSeogdEZn4b7+tv0bCYNTM9bDUvPvmAPaY8TK943EJOc4MCp5su0
wqpgy8l8Z6jVFdqu37/nj3GCYuNr89DQUJkK3WzIKbOuRG+JCFIIOHNLUHokjosqvrk4XYCybaSE
f5mE/q8tdYVyqqKx7kRmLUx+HLsmyQoF1gbBFe+VjU6PFBeqTQXINSdLW7wk39GQ7PKaC1Mnn7jZ
/sfxWg0oZItMJoo0QFbjH4zytCnrvrbPHhVOzP9ZqCX75bV7bvP5UxQN3WVNcLgpTwqpIuLnar87
YxK0ji3OoI2omIpRmDvFGPwCZAR48Tt1lTLwFlJ5LoWJvK8p2ZnQ4u6rjKBU+OAcmF/6ozrnzl5S
a/b6ySPeqSnW+YeoWiGk0QCyL2EqNurYdIjc1KsFWI3T+I8c84HUhkZd5gwreYZLjsc3kM/jmRA5
lHOLeIxt47EyjE6A7tPJfrFixEoTAfzA6JPIP8dkW1Dwa2a2n3AkijqMZjAUTjCD5U29dwi6UPcv
9vIV3PAMwgSbsaiCgA1vTvcXI4ereuKZXpYcV4dJ0okeSNWan5W4YFdEUZS/n0iC3J4tN7MDdMbh
TLfLZTq9GVP4RdFZLqeDJ80QsrOx9J3aYr/2E718rpNl5t88VVRu44UKzYElx+AdNfbHGdcRVGtZ
mslNwKssR+cIb8jLwYJq+Jq2rpIrtP+j7eiGZORlr2u7w+ZMaDstDan8H2EJbftxbqvv0M8e+vMn
dlrhWzt6Zs8CC6etcYYMejgMG8P73IoLjKOkABpF+5w3ojiy7Dye2cRqbKncqcWhQj4oiarlm83M
1xjReE5PULwwK9gITosPrgAFf9kPKJe2twLnryqtVKtkyBRIImtnT232TPYr9ywKd+GMiwBui/ut
XmsbAqTYv8Lxrt2j9jhAqEVe+8xEhlufJhcpgU5ErwKUPuv66t0M1nQNZZ2PCtTeNc+OogVn6vtY
tdmqs2SgKnApAaC64sa6OIS5qlMlhxgUJ+sES3UWbY4lPTTjw6rNXJ961G9G8n1ghiATQeiYIidQ
1OW2ElXg+ZUNcR5SD6B0KM30yesr36QVGZtRTT82aW05uu/GXu7Sk2EcifxfAysbh7iR8VfRyTj8
QH3hlyciO3SLQ6Pv1vSmhg5aZxLAQcs+2+1yPso34BRLRRO8g7sLIrKcALsb9ZIj9kx327BrJNoB
E2v8c0Zd8m/C19JSBfbXSU+bLRylcs05ty5nxh1naIJWze99ocUzBhVNAOunsViTh56z9bTeLVnp
o03JiitmZtlhKnnDC7aWvhJc5W/uN25piRxJscA/5JGD4SpRjWipwHPDN1RHFCOtsPj6JekXNl+2
OZE9iJSmDillUePNJH6d/R4zqzgopWeGrfrfyPHY+P2E1aK+oJSDtLTlW4WPCdLinwPfjxB2V9hD
MICNHqEUNZlVfEyCJ0vZUDNNRSgwLF3fBythDxw0rF7rPUmtITpSpOBDu9UDKFD+BonnXeSFOU1f
HzMBaFk0aqXTBTmtwgpQJ3VYlYNsw01PEjhUentSNYb/1zGkw6gP625g7Xa14vjE88sSgjpYssIa
Fb9OwGTMZ8HJ6A/BnmuKLdw6IX+94JK4fmXknZaH2UQpe1AL7CZ5cuY3T5ArDQWmg9CdAbMEAQc+
1o4dcD3cDSYMa1T82lumBXUzv8nsdp+Dd0BZk0uMCNOSO3gWrrQdeFNIDBRfVloD7XU6Fy+z3ZDO
gWYRKzM3P5Scleq0J+KUFzu/8hLw0YYedANHIKVa/cOHxeDSJmM4HlC5LhX0kqz48BUS0yYQSgD7
UiYazlqWCEKZVlAw+jclPpoG4fgHBN5ICYXgdSXVpON53LNj+BH5NCiwrecFAUSyvDlQIoHrV1fe
4/M61hDYT85eLfIQOiG062rYFV2hChFDT+Cr4WQ9HtQVFpI1cSS4abSTkMas33iA0W3OglDKmBsy
JMM4B7/8n8bSSwxo0AngKAWj1WM9phNazd8WrWQDMLzga+o6zJPeQhJufjEnK3psisoMWMn/4J6j
7gFSqBL1R9KaCwrDyWPVYunY2J2uEXT4JgId1/kP2d87L5GVK8sAlGDEwAlyW1sWHjFQViwimTyj
EL5B4fz12KQW4/B0boEYBlwCAEiEE5UtkXaTy28witcDuwgMVH7LvL6e4gcv6URrxCRFAEvF3Qff
J+mtbcGt7h2YyNzNMhmZ1H64XFhYNDU5clYCOHqCacSy/KYJXAYUmVKMq2rYWsWgnGX4WxKNTIyy
3r7VaW7MVgsh3muVy4AxMKCJVS07AfMMflMQvLY5FDKqSHsCgKTy4r4ysaoXb/6qr6TU5rMwtl7E
TVDJyxKp26oifCmNrbO1wdqY8VLth+DbIh7eOTqC5rc/MDrhc2ySkW7sQi9izz+vEZ0tRdQeaGyN
pPE2t9WFh74NZNgg0vci6B2LjNUssiiUcHzcrl69L150jpSlKs7oFxiri0jWAd6+GlTwPYs3FgF4
fWq/8iZXEW4i6vijVhgDBKBvWCfvN8N8iQkE/FtuQihrx55ZQvCEpDh+5YVfdZSBSe6pc+eXZrWH
/3YWK3SxzgCF7fmS34qN9VQdqqAsGj9AgsDngYxwm5b8kY6xvkhzHuvqebjpwMUhG03A1FX5XPnB
ZX/gTxmzgN4PBuiLK2EcWjh8B+m3HDlhNQmmHo25UMsc36R9xyiPu0i/VcoTkCiSt6qZoQslVQRi
8ViGP4ldrYtpF8lbUPegmHaqJiOVUIM3bV3c9K0gXc10+dAireiNbfSmU0H1/rz0IhXisjmtMCYC
/ni0/PZNXNNjYUHNvCp5uipo/85iVrQjqcLq+Qmz/5cfxFsxnXnVhh8hmapea13ApfPqlsVHchj4
hVO+wSPunwPsJuc27E9/NSYZWABbKpHUmVICEGv1pHpLSlFXvoQixbI7KFxM7e6QxG0Zj1gC0Nzn
5khn32NTGZAcMpbR7EdDEiXAGy9QAuny0fn6PsYfDYI9C/RTHBNOaJ0xtkYu/Uc5P/0AnFmWRn85
+gCe4uhC37CcXPmPyUxvW3vdyLi5Kmx5xB9jXgjN5RYkRwUnR7uUbD0FXd0FisDUBK2pw4krrMBN
RBMtM0VnQ0pSkphaGqmJ1/HojzMT9y4XKT9ySOlzdP3szmfxrUVBNg0Cd4rcMEcjZWGDz030jlvr
axswlLet+BsjfCJBUoZTkeaX5Zx5+fEGfC11KIXD+P3LtPPC0BWSsXVsFAfCjm7Tb25oRBlf8MLc
vqF80u6PTwLMqDOwWbF+/kDNtQfxacY8HEixhkcHEunN23o72xm17PWSycp4ru9wfGnRYcL9kaOn
UZcGiKcY8BHA0aPewdhtR0JNonlIPATm7VQQLxu3di0RrPzO/LylZAdHQs67Dinp8jeJAxceG/AE
JRl3UXcsS3RMCZu7J0FoMeDJ9VkxwW9aVyJgWn+RBiB2NhtWXzebvxQmNnqFD/T2AzfxUxcwl8qX
xTFEt8RSkpCxV4tu03n3yUTh3OtHzQrkUJMgbucZk5rVVuiv1XZzsUW95QhWVpEI0I4HcDpHMu90
/2COQpYmmnM/4o8EpXc0aaZ26ByyUTS52H7gQrBM5afXfuBlM5FwC1jiX1R13qNJdayKjTa5Zq/w
W7zpyhKWijT7KCCohSYn0GT816CDGEWGD3yFMOB00Tt5eGGUrt9g2opc90MqjKQAe6LblgvpBuxc
Mbgc4n4KzfqPvcNWs87D4ECTZL+ZgrSt+zsJwGcK76h7Z5yaGP5MMu76htrH5c2feEgFSk42F+4z
hSKCkelrRYQWWynoSM+CriEk+7BZgvfwQxsvh5qYO28J/wW/k8fKdU7rS1dXBzHK8ArVl3v1kaIA
XpZr+hs9uqroZwAy5w5Nxor6hyKt/pEYD5+IxPdKjWnsfHYSQgBb5NhyJ3fKgtWvEUNAnDhv838T
jHisD3QpnarHHXrYILfYn1PZYeZHFpQsE1/sYyu50PK3czZ0d/ghGYaHGTxmSBGQkJwKpIAmWjFd
Kdrc2VuySpSXlT68fADRr+ksxYPoZdzRF6n6igxvwjfl2ui3BNcCLpFr9aV7wNCBtjYk/MQh3VIM
b2ViZ5lXcen3N3aatMN52PLe1oHlkznruquOQMAU+AsQu3wk2OM92IYGhHhvNsHnDFw6rAI03XiQ
t8l97C4pb3ZGfOQRmlS1EOOYrx2dR5CRNgAFwcAbNXTqBCdN2WP+aFaUF7Q6FuV7muKyJPactQXx
L2w+olJntR4y7R3l/v0T/QDkDiFdYm+LOi+lFZSgJH1C/3gzJqiALIrEZQaJ7zBa5OiWa34D7l3q
8JNTgy0qxWIhOWYVHHquqSytiaqafCE65GXwKOilvzSb3S4C5YIQAaHI5rvI1M2BJFLXomVx28yX
QGDtVOOSu1eP4/EShy8rTjhSjzUCoqcaPN4f/ywt57R3mH6H/VU5JMFHtqXVyg7Shh+oNFeQu/vs
h54fm/ngiKU/pc1Bm4hEUD6VgFVgSDRi3AH8OwZQmUtfHPSMEu2DqlEPh+ZIakh4Nblv13umYZeO
nK9T/dBQ2RNZ7crTmtOb+/XCSHqbudymm7R2mSpq3r9QVimELia5LHEm5d90xNZLWnOjmQYs56J2
qy9Es575rJ7Xrf5nNG2XDZw65QJErwisND8B0xjRepN6lQe36YuIc3WqwJheDBv81Tg03b6rHPN0
10HQK8h4j+VA4oIro9VD2gqIxLXNA4yGCUs5gwZ8TQExZ5YJ+qTexFyaBVzeHtJXrNK/CM2tKb/N
WM1XxPKCjgNSLp/uaLd/kITXLLDo75LH3FZyzrRL523ckRukHcZXykgbZ8Br0hOKE5k57BUOEN6F
BR8BdGgK/7x88VyxFUs7kT8mjy3BAJjg/rt/gqHDpyrzsrSgRgUzUQBQ6FqrYWBnEtXR/3h2IIyQ
p13Uk1Qp3zo2wtnan35GmYNKxdfnK1GK/esoBRE2RXD7E2SPIJ4RqSA0C+nstrDjsvSS0avlV1Fz
vaVNIb4xhrl9Rw+bYa9vqZP7qLccGAoNOp+x69JOHsMWA+IaIThwIbHMFnK8sKHyPirUl5182nw5
2tjlaMgfXD1GsmkYsABkChCBSJcQUvrm0M08nSo28xcnWWACqelA9MainPKU4gGMoT9IIl6doA0X
wB+S5j1jM8au2xn/xKrzenrN8Fqlv42j1rVMV7x6wsP+wOzK7HV8McLrLJn1C74FLKLEF6vTGbdV
77CqcJ1Z8zl+mZ+TVdmDyUM9rAzcxVxeFmyZx/4+fkz5pNjeRuG+Mk01ADIyNzbHP5n3CBvR3b4U
Fc1yomHcHS12/5BEAvThR09loqP/ajvvhgnQ7kv1b4cMSvqNXkhUTh5N1j/W5ElWogvOSLTa0e52
iwvcCzjnIfkMVNtciOlwOR6YyoB7TQ9k00gU+2VrdwM0AjIyMxcd2FQLsImfGrHxEp9jLCtYPOe+
iojeHet5TTl6OK21Ik/LzNLLzWrEblFi/6/S70ZBP3ITuudZeWmCsDwh6tPrn3RQHrYz+X2bGdC6
fJD19oOCh9UcMSNdCg4dHCVJhZUSKgB9Vp2rtLUKmmWzGheJzJGQcZRw6ZcPnxj9c+7YxutMulLj
CK9zoDqb+Jyq2Q5bTr+Tu6NYKwSec+xK9pe89EIQKPWq4xndHBSBu1HulfxG1FGIH+1E8NoXhdC9
B5rd2ff89W/En7Q8k8MVuS1cak8oamwKavL2kg8qxoORDsbDrqWtjJWIGxA8Cjzrp2FinuTb5k+G
dWheDKyUcEKmkiWXqssJ201eI/KGjGnRW42QAmKTKa+gnZwYejfDsh0CSAEzRXuas0f+vQqXSHZE
fWA+I/X0hCLdfW4U7pJc7dcY90lDEINhjasaHiUVlBYv0TJ6wxZZzlZ50yXa+oMdqkUYnVRdLpWP
f964ke8C55dYLK3FoiQQPVGwt6l2Dj8DkyYF76xzwCqgvQemyoaeWrnYrlfJwVAL4aBaLbyE32bC
18Qv7qqk65+w339XUxmSHFdH5O/g1xbp7mgbkw4/y/BDpIeddYxIC5tJ4OqqALUI3Ugum7p+/1Lm
V9vBr0GX/wzx6cJWyKlr2i7VnN3yAODLpEyCWZTqQ7ne85H7Z7YPnKRyyJtkE22hAPVmfDUB9+TC
N5fqtEUUBK4i6gjHQ2Qk4KnV6vTnnu0+80P6cxhDOI6uqIMEHFEJW2Zv5MJTlr7IMvnxXjKEXz+l
VkaQr+2wnKoPAm+W+B2bWZ7JccxC3Sc2FjO7R4shLGeVdFOUgOrOTVEWBFk4Wj49sG1mNBB5+Qjo
UTVylk2kT90zbBA5/wLsywQ/cuF/EJhEYCpTjaSpSuvvhotcm0FfKvBv+D42rAhCXK1zxN5HikrA
MvLl+5wrcKGBSeL9iNzahwXxXJ8h6S/1gyjnsIYWmn3QazXIYPbbmPrmfC37jmqp1h3UtpJFlp0n
EEINiX5ZAJshArsMXab+OISk5Ch6xQ1uRU3pfg8e8CN4nzEFZeeJZwfbw6rEgD6lW3c44ynZGtl/
iIWMGaul3/X3WzSvdjCkVq+/mOb/SQWH2MZCIWayKeX7F6KtuXTbk45sJs4Ttd2lbajoaWJUKjFf
LwTrXxaYXPuHYri1xS462xLk4YuHIf8gBZ0rP/9in0JUpp/xsw06js0/CRBmNRVC77MXqBFuspDX
RlosNeCLzVJ4i+P07rxU/BLKutAdTPGVnz3nVHyvQ5jgerHMA9v9HiEYrlkODIeAIxhrr/if0yUD
94gbUx4CyNxgdoMkRaPeiLfdeutiwlNkG41LCpzAAQP/ewsY22ExzKv3zjOpPvKK8t6Xa/t3QT3U
GXptD2FwzlAWAtUw80iYoGiBXi63LntBK/S96n8RXyVO7XEUdgESAwE2mlmWd3H4HFOdiXHtbvla
AXntJrxSW3aQdsNTtBLxASYlO15yn17RjY6Ju134PwI15MCfYJy1Z8R0U9dGy9q/2OxseD74yHEa
vhZ21Z3BL9LQYlrEP8ZqVfJ3zZcHRH/q62/e4aTLJku0fRuDYEiMavwDUqRUecT+Jsvv36xbrBnk
XVZsu6+n5INMQJHoF5lCSjiwqxCPqEkWmcuZbMsoxYJ5joYIlkIgj8gyLpDCEC94RvFMu+CJZv+3
kz96UYUcTIpoaXZGutJdBPm6nQzQPBQEUWxOIT10t/QKU1ktnva34hB2o68M4HKggNa/ufIL89mw
o9ouKtCG4erPfHYXb3gSs2vUxASyfVp1jYjfWohjqiakCS0OwYVkjzz5TQsw6Ylep3E+kmTNf4i2
C9CAgD6YFZGUHjHNIIUxMuQUleDgCMAwOpz57qb/XxwdfAx9VZYc8vOgj4eyTHlKxHOZebz7XYYS
tUdxJnYdFpCY/jNLikIFsBgSFtgnsf/hWwwy4i3es3RBQCYm5gVVcmrpgvajGvDtIDDYqfdM839S
sOvGc00mmIbffCMryipzUMBZMSkobhZyLDoVxohRkmDDEAGy2gyq2Updw+yOBLaMl1kEhOUKgvCV
hmMMgY73RfeVHDWXZ0M/VTBOVhpS4vIeQgpTldctQQdtvONB5GLHYxeOSKBHfOTUWoi+p0Fp4EdG
tLnJBxDSqE0PG0CQlg3Nt7omfpuSRnO7AKFfcWbmligho8o/NTYAlUJ7wPqUJ3rSkCoVoYC3impA
VZsX9drUGLx1Vdo4fN2KsWdd4h2Pjpbsn3Ij2/JjXS/FIiRdGyQX5b+1tsCho1BShZRKwGkugcxy
11zWzTrWluIB53Psu+dZgS9sSeuXwbzgGqsUmk9Q0CX3SVuedfU/tjPEToqDyECglTWot9Now7w/
7Lh5c+TV+WH+F5v57XTPtPR/nttr+MvEkDOiiV6P7FEcGoeSykZPEwujTJ6nj17f5sJGNaOwVvdv
mOJcMmYMsgVVsA1NiAUl4Lisdr0MVhE0nXJaudQw+FnMDqFguGe8ayXfg4K1SW8T/+qr6UfmEX49
6TI38w+8wtk1gOthiZBdyqU6upCeli/RZYlj0F0pvor5deJlk9Pm73eWC6SEs9+UlgCW5M+ATg29
+TZ3MiVn42PS/Bc07LHokSyOOj8UYqjdjXMYL6KLTf7MXbexOZqbhqqckIvsSjC/TJGckpT0F9Fr
LvbiEkwuQVeFsyCZ6J8Qmzbjzxpv0g31ewgqTQb2J9Wv3QEj+WldVbo1sLqtQ1T6xo05ONPWik7/
3oyO1oRCDyXTcqjsus1cZrriLmlCVFTRzl/zwmIW3T5B33JG81e8jY1I1gOx90hjxPC852p2w6da
prGKQ/BR3iyhPQTALYjf8r/wfWddc6m8fzj9SrRgpGPE3vHWhElqto43oc/JVICpV8pp9PCJqZNa
8PX6DJVnwMxppoqSbY+kGvcOODu4eRglW6RiH19sZH+15xEzuDt++SakToTaoP50CjsPsULR/Mm2
EaAME0vffmj1+haHHib9bdFvpdMx0VcxR/Bp1DT44jYx20YqftyJI/4+jRz/9R2oDQpbwN1yjsgE
KaBLK6ekuE9ECEygjfOj/0RvPPo/GKyHGTTPlEipJs7lQL2mP0ytN0TSm0oy6eKZF81Zcj+hT8mI
/p8gCCz6lJcFsvP8HGT8ZefqyYf9hXLgqo1NX1/TO6iFALd5z5JhpOSmkmy/lJxjUk8JIHiQ01T0
xZm///oQ0xLbUNjN6NvTq7+gfKY4bawr/SztxXsEl2jmVCIKJ5j77QhjWnPz6EeuWDhbv3vAWDfu
05k3YKoGyoRd77B52+drz+A5WIgX58uECosahEprqwVAW6X0ezg1Dbuf71h2VNPDDFgeOifHcY1H
2JTuv7iI7XaRi0iF1pTGdP0INuCz4nBna3tNBvPGp30BTu8/5n51Aw2ShBdsNBDDzb6zV8cM/64U
zxuT1bHjuFJFVD/bnT7DRErKNsnnoCK45X3/ajWEleElHkU5YFRzcGu7xgCb/nKp6BqkyHJLMjID
imrKK8Bvl9Y9CMIuDhXNGF+si6mK0DsGJ1nwJf2zwtqYA4+YB7wipQVKwIa8Kv45tcdiDLn499H5
Of2yjt2NUbaVCPaZY4zHnbUMlpWYWViXJRI18R5KGXz1eK69gYTTa15zqTrn4YRbtxFJg41v3mGi
NlS6TsloCoiKgrHYLHMy+2ay4dCFEFXr+B12itlu+9cAZEyUblJ+FkqE9aKe8NG0g3POCvNQxJmX
6LaWfPRvKNSys9l2OMNcja/W4Dq7976+i3AZubIGQtmM+4lUK2o5MZ+afbfCxz6EWLhuW1lvKTrR
qzlN3ncY0DEG8NhYr200s1iZTxbqwNDFa5lW4RLsbi3WkkJ0khjM3KAKVcewTmOfYZimybAg1rs/
M6LzivQ2hgAH49jlXWs2CRZ8kKvmIAjtNbm/KodYgldt8KBe7oElm9STCbu/BjTQlt8qQQ0JxqVK
HyyuvtrjYu8MlYiU0QUz7x8b4aq4NDihzkFBdfHEHLVc6EVoLi+T4PZCOC06LjSkMeGzvY5p0/i1
ZOPHQYGGRtczwr5lW2uV2HQK8Fn+Jc3iEz58WVUH4DQQ10RqkUmLwovGb1UykwnZ0l/EdWZQpyWT
hNQs9BRlTaGNNZXPHWMTgSJdm0Rf+5Pbhy1my9HYc8w9SRiAjjzwMXxsgqkTnNqcDASxa2xoPMev
aesAqH3Uvh1Z0W9+1qXAIN9zrCmjhFfINDf3JEPScsCMc1eRMPwbdUGBZAZQ8ObOx3imUurau+br
bpLSRn3/X6ES2Ymjy0yQpK98SCMqOJyFNx8+bRepyfwtWvQ7rh8Qvs/sllQD/WfWpz/fWtCaA7/y
fKr2AtqwkSrqR8Nbp6J5CaWTyEXEI43fU7SZf1wJ5DJuAUv8c39vlY7ei9CUCM8A2N8cNlfpcH7f
ju6r+Tdfog0S2MIZz6HeyVW0RcFLyJTnXNLLrLB10elyoRCtY7WqkiBJj9G5X0RVjHDbhkH0BNt8
BdOvmmL7WxFEDO29YYKlXdby7E5T5zYrJZ+d2UHe+mNG66h+wFBtAZhioD6SFK61ek/uXod7OM5m
mPK/TwoLB2lNuwZCgLXFi9I3nmCMuq/w3SV+iFPwbhQHuGxB9SVCZ+82bUHoOssnDK9A932+TxGJ
EpdxZMRHB8sCmxr0jBemRdq/ew8SYbwtNoBrdqv0EFD8Pcfxe4LH+0wcFg5SpgR477isGtMV6C7j
lvjD5DfWGnQKBez9FgDmAv3FGKW2IN+E8yWOMmmdQRRuDIGzgS/2mPNvm9sSRRuPz/NuOBmVv+xv
fgdZekUAYi7Gd1bC2AdFO+c2NzvLO550Fv10J7oV1sSKAIAJKDpYOWtpzz8QTsRjEWkkZFoSd3zE
MEG5R2OXrJpmMr2t5LOjzuSlceNSSzRO2gwgnbQht3Df04+DqKw3fXsnC8uWQZGjZfM6K43prWQ8
M0VEGqz+i5toEIL5xYTosxH2nuklYhchtCTX7J+BhTrLz3jL9AvYT0hGAa5GsMEBWkce/SjvnssB
55s3wOyOURR950BxvRRKnKQ8Swgafyc6rlgi8PyWwRY6pPZt/4kzrnePLGxVUU/HU/ZKw2m/5EuK
qYrRfcpd1c5vfpuxAn0Wn7fDKpk7EVpSzWtkxH2cbfy44BfyLwi+VvIP4XsC5OzWWKeSrBzXzIm8
6pEeEsK1d9UFpcAcaDa1dPUWA6DK3t8x7lNmW2m4tWXBEqESLur1xip0VrI+4Nr2kCy0bDM1wRaI
By1azsRWnklySavUI3q+cRFbBKGBTLcNeh/MP5b7aK2Q6IiEi39x2U7sqvts3pVKBDoaTbhuRpaY
3ePP3a7W7DoFMRE8eLaSXOiHFY0sdRngv6UAfB4XX9TFm6xEtAvZ4nYrhFAgl5jsoPBcH15CYsCA
NOxctAL+ZWyq6vvG98CQF1oky3MWfdrjzVy2s9i2IHP1L5mG6GUzLp//qIktgE6uogS1tEjSNBMe
Bbb5c5jO9LKwCOrdxR5FRaRe+wTaXqe0FTTrOsiSwITNMTdQuZRxc9gaSKfq6XBn/a1kdBswe7c0
M06fOc3oOp5ziy/oy2np0hbO6vHddLwkyVfsaQNGw6gZm1GGCajjfKP4iBYxFD8WjM2Fu9JVYgx2
Qg51oom8gOSXdjNiuxRHyytwOe896wv++JUT0VK8adF3EQyy/pR07BEIJr+FzFQdHiM11BYFnrO1
+rn+oLZO+sq/RlD5UxsDTb9xLwZKGUD1/HvDwSCHiGIDOfEEq+5dstzy5J47zCKoy8u0rfUf6lc0
1g49XETAtA7wK0x9WtPcP88tDANsPJczCp3AYEE6Ku9Z0HVlmqu1fJUiOKwRk0UO8aTIVHAbxsLl
Dl1+Z6+MlceK3wkc++boybgJrM0JoEB/p6Gg3dMIEGx6OsPooxjC/U4xHjddScMyyGRvyY3vGiR1
KqWrBtLKTD7awsMQH5XlijtLaKPYMEgSdBeaJrtqFmjEbNVUTj3D91DjuwQL+uvfsyn3DEP2K2ny
N4Pq31Jq4QFt8pt/nEuFmNnfs+fZqv/P1IBL5P7hrwNpQwsze7X14hjDiKbIB5h0JOGO4ShzWewe
zAqky+0BmJEjctyJ58aJOHfgLp1QlwqD5g5SE25SnXfep4ku008miQNuFu4OCkpvcziE6jW1YhCc
YyJihVD41SmOvAAVKX7dzvQSm6xf1ajbkEkafKB3imTtCf/vPH4Jvk/qtSx7E9LmB8NrjX/LfIHn
cSrysUkXFeovX7bKU5I3thdpHQZvJyublRSdabtwTNMiOtkk0wldbQP8+aCvi0xcNxex5MF+uVb1
cRvrqtA9fU45obzCrHCCqlYgz8Khme4kPI2h1vWyaCwAq3Pm30qDEpoAhYkopGFfAmA12OTsSn8C
wPRqS4aCZhmVEWXaZQAFmjIXPo7PdqbHzY2UWV3b6hmQ6a1ciEfg9GUMYlsv2+A/AKdrALtvR94z
3CJyvlkHYGETiqlPkZaHZa3RUl/BNlk3d6ULzjeN+XfHljcLKd+QIQ2nI7KwyBS84Z3AILEwTRRc
IGzZYtaTpQnOEykvJoBrOLBia73jOZph0/dnqnQLL6MYyetfXK4CJVsInjh1LIU+j0iNpx7OiXBW
anznGAzynJ73nRsnzcMzdtztPXVmAPS2QrMsPR7DGy1gm5s9UTI2iRRod/S7HI5edOKhtNHg1rS+
xQKA1ZvgRmUzmxfRBCqdnb59q2HeO3gNeo6zUk2Dgkwgmyakvz8fQhqO/VlQbW6VL0iU8xT9U9c0
sA0//40cBe9WJJpDCbHKzYU4qrrbGMmagNZiwH+KN9gCgbNHhCcDIc16EZA8feruCFkFS9ytk7Zv
2XoJ/tlyt4OwJ88oLvI89qm6Vhz0505K41huQcc49XLKPyNaIxQz/JllzU3gTyC2k76FLZ9q9bfY
vbr/2M94YqamZ4SNacvHV3jxojwAx0PUPT2R/oSTs4nlKGVcAwz/vVV0EHI7oaIc+42xKq7nGATK
QAsj/iaNk5r0cW5Di8GzO9CXBAUEHlU8GOe2AmWpccY27hNeAFtMEMMSzxC9RAOHubZAR1GMxAxE
jgJ0ZAmODcI3KvK66gVg/3vlWZOhKFwoIatt+HllN8bOqAz8fBvl8DdEOsGUDpDWJc19FI+Rrjxq
7tgPF8vcdhS4FiqpSZKFVleyPUm8XmXSvM27OqeFW9BIDVpqFooI85d/Qo24v4Dk2wKVv3IjGqfF
kn1RtyXwU17iiYONh9AA1h5gIPMgyUCQBQBre16txBTrNxLdPZnzaStO/+40vuxk121J08nlPYX/
XBzacpkT/uikZT4ShxLHI4lpRX+OGGot6Ia9I4X/5uYmtFuY4Cfya29ztZDrxwdzOmJfsHxap5BO
wYZeJpaw+Xw1KVUwYy9JZ3N0JtiaKoOsAaKeqZHnk4wL+pVALi5cPlt+JSYWJxWiPG7nEg0my5Zy
sfH8UVR2MykjWEl9c5N2dRZbkh7sg60zw6S6ioP8sSOV+h8WbvTC4SVohL3WMVajum2K5srov/Vl
JW/fNLqJQ0nZH88S5FHH1bboVM471QyvPDEcQqjW/GObSWDCFcVM3YiDwnxDnkiOVbuaVgtMqQWp
tTjqMrJCWAZ2b98FA8KhHlZCqpEQtKoOU/UUWvgDekkbQZEgO+QR/iOgVNme1xhchE++2KOv4prg
wGN/AB6OaHstReNud8Q9yp6jvgb/O/wg7gQ6H2qVi+hu8EetNzSp+4Em9uv+MDJSSByQ1nq5+v8u
KhB4DCazVs/vf8eXCIpTyuU0G6UdOP8lR2tMeKq9DUuqPwg6cixD6KS/Q9juUdFbiHt7mM7V4HvV
7zvK8iel8YIzi3VhT222DLzPWwDNXjwc7s6WQ9xgUNf2e4WJuUolmcFzmo+BS9WGjKrC8cftk93z
lQzr3OGciZ4TAVMTgbC2kyZDOGhRgzeZ/F261X+9s9h/nocRslN+QWlR44LtwjSLLjFWpU1o12x4
3ROggkEpf2NNGdGdF87esdeNu4ZPKDxgHKkVji4+mMvOtiFP8Ci95UAu7PnI7ONTSYXyfNK30Vj/
DCo6sSrrJ37qXOomF5VtodeV01kCh34zIZMbVmqbL8u5nhy3eTF012TIW3PP5td5xRcKYQVYgyzF
O5aWt7FwzC2z+UPxxrYA0h3dv8lznka7YSwE5nbrYukM/fsWU0pCyauhlk82tym2ziI+CF6M2J3i
8kkybgs8WJ7tcqiVm3SjxmePcwzY3h/51oGd3pL3MRvHZJqGpvX0HyN2GiMPs9CZykC4fwafZNDL
bi1LNdpCxegQqr7x8TB9GVWYGQCneKEfXCPadP9nUquwyREeMjeu6A6z9B+MMSTL2+rta6sm4bnL
yMqdgfuM6lIVMvtNJ9avKBN2Wd2UAbSfCEj4LZnxFqxo40Di6pcTuf0sagMc/f6OgEJc4Gt1snLw
bd5EDto9i359StEHtFcGNQyHNmE6fnybxtfHfqMt/Krdp1VbepVwAI9K3OFQkd26Td9yDVXmKqoK
A/zhn5Okn7AGxg5W3r2RGK96PcafoSKSkVTtMU4au97mnvza3QTmuHL4ZhKfIpOeehaYSwkiwt/j
PpabB+mI4GQk6fvHZ8XawJ4KVI9e456gMsyZXJvIAKus8pnKHJZVtXxmQi3a0nZuz9Rl376VInK3
FdBAI7tGRjtcmOpziieDgGb9x3UqR1u0n4E5k24RuHL8ZXSWF3gvQHr2qfzm4I9JnR+guno+ACWv
vb9azDpfxLueiBHr4qgNoTe5VF1djoMIQayZkInvxM6VZtCns+bK3aKvpN39Ic2pEPluwopmYudl
BqgEEvXNRrz/YlnrqtnFE1r30LQ1k5k60n+pMGHt6QJNQgJa7U1UUnDxhe2ajItEQKRfiPT2CF0V
+LS8K0VpelQhFrBgWK5ZHm3dRqGJN13jIdNmtxppAUR28ZFlL5sEkOF3IdqdTW/72iGVgC/B5Re2
VGx5B8ACfZ1ltXPYYxtCJcrqW+gu0rVzXWffNS3/xiF2XXfjVEn6jVRq+sgEs3Vt0WDIeeUc1TEB
o80xUYvwwUUVmtzf9ZLSV1GbGKJRlxtVnceX29oeGNRVlx+5bfJJNobpPhYQbQibTyj4wU+92zIo
ro5u9hvA67LhHpg2LFWG3v2d7tufgY9GLEeUwcvALkR2/QAB74lr/4DNiQDxxavzbVsjLGuJ/oZf
dLgYlGIeB0EEUL0szR44P6JeA/5C0I9+kjXrk7jSZ3VEw6bHFeK+AHEm7EoTjuEkovytt8Jq6QqF
8L8T3k4Qoxg4y86usYnsaNkIUpbcnIC2rEQKOfY2758/C+kJfe1O6V91b/cDVuxIJL79xqc7xv2i
FCNkVS24W7WUOmHhXEgVLqZ2y/reipng2F8pD6TyImu+SC7J90TOiuDEUOL9Ah2ARPFziy+K6qeN
fLSu3tL5gMndAiC/TsdNsvl/Yd1B2fhCcvkg4dF4Tm+bSQBQkgtrju0zGXoGURTyb0xN6v5yl/hF
GRWAi+5cfjOIq9T/OZrMqeMB3avA9CF656hk4gqkRVTzZW8Ml743W9QFWMRqOZPr5Kv995IxM/j+
WlXjBt26DHe3LJHazXF1nWe8Awij7QMaTGS/Ckub3OoAJtIQG+PaLchtPyP+fgpVmaqshobg/JMV
RR5mZ9e5sLTE0MXivgs7ZgAyjj85IeEVcUS5vnxP5Ty/GMmxalnftrOp3pHpBGf/a22J0dj/Qf7T
b8I9IcwQj/XnTxPNXnWg5Sh/R60wyDzvKz3BErLmOV7sttw4bMCjz2aX7+Y6jIkYMkIob1q7H+DP
2UKt9ThBNIrRfdRnOBVUxRpkznJZatCN/ZxZcfl4oLJfawW88Lw3u5k3ExqTX9jrOqez2kdIMACn
PZUMQXKJQTVfC3QgLiZ0xY3wbeVOBP2fhmK4nON4gATfTy0UsBEDTdJCU+Nzk08eBLSEZ8MZ1+b9
S7qAknvXXulTRKYlAPFnKkDgucY46SCg3BhzHnoZobIqTLpFslAR1qVYz0hu1QUGXPKDshC5fLx7
aDZ6GGJ2teG/ZPxpytfRi6RN/N1TA5o1UM0wXES2okwsUa2nITYBNfUaE/f9+Ny2ymreicxZK2eG
0u2bvyqW121DlFIUX20C+JBkfmEh5e25MmAsGj+EHwpZ9Tq1h8I7uEIkVrLGQd6qO4cQtovfo6VR
L6PNw0iNLUvsyt+/9ADhnlW9jE/fASN56/f6qsjjAXKE96+/lWPKIS7Lw92NBsXP3C5pnnGlDwPj
j3dY7eb7crEZKu6QYQPh+9BkY4jAzVVHv+qSayfhO1LuQv3L3f8CeK5Dbbba/Jyav0KpaEi65w2i
Oh6VbENn9C1fkBlWUDt8ZUGuR9qX9Wi+fNsOvmCvF58RRT6gQIvVnKF6NdbCuyIlnDE8R235xhZN
Qsz1a+/lMmUKVclGw6dJHSj7CBLTboK2PKy6ofb0ZvrEvGR4j59iJZBKTSfVEwUjY+lr0Cg1FU2y
pt44G34ifdNCatqemb4cVfOYj+JJwbDwwB7bZAyZGlWNq7NjWzpoS19Abw6SFf0S3KTxRpl2e/TT
xsP/zs1DxoYOEELCn09TIpJON5ZoIuGlG2N/Ayw7Nlmv9nciPeRfd9D01S+uYi9+Ci1KOwa7mu2A
HMfw3Rinim86I7g7WCbT1Y5QgiptwyvLO4066TMwbt6J6WsgJ0a5T6bsaHQSxMgWpuhZTEsIc/hF
vsUxPP4j7hAHnTfMx9Xgvy8aCqJhQUoooM7pl/hJvQ/dBnzil0OV3Ti0WnHOmhqdodNv6o0PDmUt
DPaP4X/0grAemZh4oMyBn6CTnqDv9BDgRJm8APGAY7f+r497ZF2lCTHFpLYoqZLbf9L6TvyK7ntF
LjWfWSK0puqpIwrmV/SuKj4llvY1tPxpQB6L/8MI1EXYUwd75AG/E0N6sPS9aQLGLZKrEGlETkFP
XR2lFm1zZFUb3X43Ll4u5+P6DSOP3jSS5kjzlMS/+D99cQ97QdgmsRYUst6KkDaHXumne0Uc6+x2
+imCNzR7djI6Y/3MKYXNnDY7aKkBrK1jW5gdC1UWddTw9N+EV1uI8VrAy+TrOFv6Uz7MbjQ8MB9l
MHKoiyQYYtKKCZkZTc6z4enaAR6VGDEiVhlGlFeHaQueL6W5AgvDwIqImlfcO6AMAwFcEzd61gaY
Nm2nPQq9h+7kFo9aKjp9E1HEx6kdHhx/m2OphsvxTrZ8IjHs4o7/b7dm5GeIltzbL3x4IFMqng3h
WOnjiN4zUdqi5fZV5BVhe2nVXDyGdKkhPSEe8bc7c0v228GeOKSeAruE2nCJK+OwJYMF3SLbNuZ1
GT1qEYeWblIbHiVDmsFUy+C9iGL+xfKKLu2H55ZZW04X4+HXhILU9wGBh25Evo2aH4zM+p3lGmAW
3TKapDNjirJ0ZDoh5mrUtxGoDhNaxfUeIRWSKGe4yK0TAtZx3ESXKZ1zj7+m2t8PC1FcHRQmq002
fdMXeb3beHPZ8JJVWm5VYXNXovTZOFVaMxuIlaTw0ELog+f6KgFDwkerDwiiLU2yYECkL/HB67xE
QP2ETc1pFc1bcET3dnHi0+8LndYcnayxJRunUg/2KnDC/hF4FCHTf0z+Mm7PjyIWHIkEfdyhqvvb
ZbyDpUBR98Su3/C/PPx50q6i9aXaAOo206vL4tJPG0b+8ZKrsKLKfXg1VmBp8qmXPmW/oY0jERaJ
/hw3tTkSstZwNxIGErjP+ZRgruGU+nnVfxQOYL7BeGptsfOYJqMTVnPdl4E+vVYOPCVNyAdIWvx8
t0LmiXJZ27/cW/UrTdy9jkPGW9NicmSrsbUoFhOY7a47CiNlvhW8H1t7c/urpVW978Gxh8ywdxhm
19mN7s/1gkzs/0hRkC40DZMcAMPl9KisbO+lYxLc6NirkyOUBuJNYFF32u5JG0SYMebc3sqF4+ZR
GmQcMvyib/2HzvH0TqR9R3KeSifRzNUhWgaX+xVglpa9EunGJCXITZ7MVumMfpnhRooCFRdHOy0W
0WfJFrJCoFg31dzYCrr+cXSQ/ztXNjbJJFT17wCzhususGUbdUPGAR6LovTGbKPwcR1PryTc21az
hxRrQo6+32UL9gWoKbSm1XElgiYHeOxLsZeUoctfHNb0rcJwoLabrKhcEigctTv3BTXJYMcV6yfo
csV29j/KtSGV+sNEO9tvKaRv+BSRNuYoWn8xfIMITDgATBTKZJwEUYFGnKm1bU0gwcwoLhLBLZ8k
yYkPNgrgd1sjz8KC4ceZcMwhmIT/zOHfhwyYCyvgWiUjIM0O7u3/SbThz2rQRQmetClu3PefFwrv
9gFU66m3NegB1DqIooBI+WnIAkVOIKe6HuM5n/SmrIy7jY4iQ7nCR3pDSzLV9UCsiJCPMYdWu5yt
JQOuruxO75Wj8M9DYCQSlQ+/WkmtQD22dEF3Rdw1a2LPiOVCgQ3dHyB9Z77zxFXkuyjQnoVMngQI
PnnSVnIgG3c5OUKY3SI5DbHmPXfjikljbjJX5KNbitZSu+hmgPlSgKHs+OO1EPO1/kWkU77l75mZ
obgECey4rjDBjqM5XLJhe2pP4fErII0y97plD1dOVcxTiTSYI7GP9pAmSGz+kr58kaPReOAR+CiL
be0BhP5rLhHjRVQTVbGJSEEVu6uJIuFSULT7wKPSt5lQALwan03vXNu2nYJcjq3gw2nVtcvGuB6F
LwevFOqZ0CI36ZQoia10Htn8Uy/pISF7zFTOv4FbqXZR9Gj7pvRHYwKoxGKtcpjPIOGVNPeykk5p
AwTgq0S9aSncZXnqKcbxUKlHeg3ZhJxZxDnZOEA0m0Fiu/VSzF19C02u9cpHMG6S6qviHieem40Q
3jIQQ1Z0FYFr45DdVwU3Yv+Ukakud2ms9pesYJ9W5WoIustHnRUfD36Hch0rRh0cA4kOATm9upee
PnSiSWioQbZmxeZjIbjygmwaqDk5tpXnmwryCWZT0RbITRx4lm/Of9t1QkOvQpY0peUqK/oW2DpV
VGKLWCMCr1x4wqounACKczWr2wzAZkyRqvEooABNThowjTr3gPrsDsFrgZVv2iyA9zWi0WjXHq5o
CcB3cn0BHaCEcYGpyC8fcnLZGzJEwOC78fa60uPKMEJaf5KLJHMPQZOxyuHs/KkMjXpt1CSPWbo4
vnwxyickGZuzqs0P+te8lZ0iADYw4TFosPRQTrZg/lmEVlBcxKULhCG107N6Ma0F4vxVhCb+v6ue
0CNCH63psuhXVg9RR6dt+2gx2PRlY8uY3eTpQLLtqWGUweaF/w7l5XLAeBmnk5CX1jnmAOVYZXs/
rHV0tXVoeGLuH8P/1t0IKChEU2LWxFE/RstsLV6qMubreKOVAazhgt4CbT3idO+u0w2/FfamOZOZ
XIfJzMZ7wVSU7gyxlnvoVZ/1huMHT7QkPQLOJvyMhttzr5m8nZIXNUHwlRq5clh2f5uhyPAbdywd
8gGdTgfi3xNBz266gkiOebKH9r/6fHJ5K6b3gCyqw2xtvn7w7vcPxRxN7PIC/K2HZSWcZCoghrj4
KY90fQ7pCy+fQzY91MYSYzEM1A+SUT0k+veMJYGe5ezZrt50s1eseSCfdD21VTvXPKkegjUheMZ0
46EIvsdFRk2iVu8fA3egc2bWeEfy5FF8tdmjnvjyrjTUf9UkhXuW361eKm+OyXOj3s3o0OnB/3pT
RIoX3bbustBNSma8iY+ZxGqNd9nKOh+aTY42VEA6qgdpUkkkL4Ik/05HByl/grS3L/QTQ/+S+2Hy
eylV7FO9CvYt/I57RoNVRj5gBy9x5CyAa/MIzxKR8RYK0YO5zc5Lm2Yx58klDZylaa6wj2Arc4tm
yV0NLfFBkuBJht0bZoCDvZegPxAm7o+5qZLPJra+SjEuPvejlvquN37QssL0reT4o6w38ah/edhh
Od0CuRbCro0JiKemj47LNakT+VaupKhuv6tO+QkMlx0tDKa7SE4itM7a1c0K9vhj54zwXbnPpFie
Dgf3hY0AbZuuqvbzqIc721BgftGlAyP8ZuHr+s4y4QXYnPR2DnVxI3nlEg3/6zrkv8dMNayXLHsg
F2HlKPIrXl2FoSBey6gzWvrbKOW3EQfU9UndQBHjlXOGwUGDbGkjWFbl9EYFB0YWr1JBcBBKeEM4
ZG19PRbGL/s4d3YMaWg+Cpsu3+3pbuG0WI2EZYW4U/tbuWvNh/LmMdLzZqbM34hKwII4l4YARRaX
WinaK5NDFDlL9jkG4PYr3yfB03K8rGDutHs5YDhBKISvKmC5IAq3WCeysfKci2Dcs88Pe8ArAaYr
5Q7A7uhOTHtUZCZA1ey/Ab/wtrViRmFxA6bBP1ZGYblYsKxbW7f4L1AxdlfweEnu4iAtUr8FsuGt
mfjZ5DTNNwKvwVxzenSo7a636B2ZNvNcPWBd65uevwaB0TVvs3MuN7GCdjylSgGjDdF/ZI+J1X/d
tRcOYZ41lTiisMN5dw8QgyhOLTkFwnpwZYNQWnwPA68bQFM5mnDbXMGCXe1H3TMhcNUlwabPNKHR
2BP2+qYWTHA3aRD1pw842kOQvN96KwDy5BdzLPEEgzbSvBFZn/HFtu7W9U/oc+wlO4WLRa5dyWpn
1mbKE2Kik3Yq43JXGif+0fu+B8SYAa/Zke2+9JjA9hHODiPvmDSb3bd0cZJ7IY6pqRkrAICNXxEs
dljP3K4v9ab0CQLBvUbLH1gMVNd0rm2ypgLBUbfAtxSn0w1Bt70bssW8QkzF42JIIwzpkh7+Uwd1
+AEAwiliLoopAALxmqRvY0rZZSxXi6nQEKQ3HgJQDlnG8RsJb20bWMTxyMw3Bwp6PB3ZUpHewUWx
cNAkKpGapUh3/YTQvV8RCY/pBWAX6pd+em+jugnYudRWgG/iVww6rK44cIUuZQO6eYpI9K5EuBec
TrFUZrVMxLLEJENh+FfplZz40KkO76Hth10vJfjcqlAFlrbGq40PrFGYgGA47GCBQBSzCVHjsqmR
a6WNTIHcwTltzG2Ih6o2jqKaY0EbsYD+QrXuaAF85IUXsxT7Z4xO+leCpwZeTDvgWbfU9KwlR8Da
SOKChnWFT5u5i3X+No/uAEtvUhnGCmFJv0JluBA/b184WvKx9zoB4grA+E+sNJ4mFqqGt0I0Pfxi
1hj3kRY252wb9V4idPpgnl5/P/GPU7M9hHq3PMUPJ8BsbLzwso1wNP6yf39lg4dqj5505s8iCqQF
ke/78ItnI7Ma87vKyQPx7lFxdGUJ/2/snibM7WhUOSusTdC7Z6dW8skfSI5PsKU2Asig5nJ3GbnX
CdJ8mTJ3LnMwcHJHojtw1dGNfPOERtkzi7B1NTg4/az5e12m5WRQYCmo5zX96eH2cVSNoLDGsjBf
hITG9k+HPn8Rs4mPiq4VklUXC/0hZO4TDN0tkoW00uqQYtzV/Fe6vSb9Ih0hd0OJHbDj+tQSJZ2n
TWt85i5Okp89jkY9IysSetyolTIZNEg18IEW+rEJz1iw5JEp3nvu3EoSND+vgIjfTvJHceyPIfQE
19TBdLJCkmP62KMGYq2+jvMt7OQrUsdbtDrJVipgQEp0tgmr4Hcrkdlg2bIc3CeXlMboZoNimwH1
mXoB4oGoXG1lupmg4W2mJJ10Fwfh8wSRggLLX8h9psVSG7xIz/BysDZZC86M2xk67qyzkR/I8mht
UKI5Nf1fYaALMwUvoF6XVWMEaHsjgU94mkkp8nZE3lFADimbc1AWjJ8oz3GrSZWZf0c//4DzRoo9
jc05+xCsvYjm7EH7CesbxtWvg1ZR0iaiu0tmyKvHLvX5RgMTUm4c1wA9muP3RA8loFnYV7d904Fv
fLvRbIpq0c565PfOXCEa4e4JOk+mz8Co/tWP1DDDf2UnvCgE5PiI3718js3WBDPm2U67ejdL4tNR
cMWLYA7LCm7ccuu5RU9emMYaQ3mR2XY5TLL8QURsWVqaZ/+ZWVhQ0zB8mqkQwarSshUTStPDKthf
YeAzx+vpyZjTm2WDd4wacaSUp4ZsaxuLVRCL30Pwr/4U0fXCBaqJroHT4sy2gjLpFXkfW+baGAC3
3nsy8EG8ebAwXE53MyVfiGwfzZHNyeHImA4/RnY0UIbtf/aUm/mzyYFrahp55pTXOewnHwIntjwA
zFlCzFz3Nv/v/GXAyfHMNIhh+yMbjAYrCTzecVv//2/2JvfNcITDu+nejmHhFsnwhSL265vR6VxB
x4/KxHucuQRonITgM3uqxDLsu/dNETK+Yz186GIsA1WHCMHrCVJIz6c+DHTzFmOe9uzw3+dwP+yi
s1QTd4xjtceP1w0aNZpPIHm3aJBO+bY3yflAef3+seDzlYaU26+IGMBcCqnHpkbAmiNdVanM/TkS
TB4zy+uZzdYrkKFVfAzaAjc3MZvRLjy8XrpZ6u9JJfOfbAvFUdPB7gQmk8MRhUVNjD99eQwmtIpO
I2GUsC8+iJYxHH4L0l7PrZL7O1MuhNOit56fGz+3a75IrH9Z8J7SQP3eGuieTy0VE0Zdn/N8oNLt
DLOCAWHdqU46EG17NM6P0CHd4XRHrQhjzzBFiz1uYR7Pf2iAN4kJ8Jz2syKSow8nvy7NDYD6OHyu
Q6hWqs1PIjIt+7rTfpb0dyLxEq42LG3Lu7skUva0YBrvJGxPIJR9jR0cQQnTpRYTYP9u4rD5xof6
jkUBop0bB08YGpAc3mfkp6sJb7jUcmZxhRbNXSYNi6EIylblDw1rsn8dYOd9nx5wSKZPd37mNxLq
o0oH8MbaYCYhewGb2LV7q0Ht1CXPkBhAQSahlTABooY27I68fQSt96CvBnDMFdaEATZ6HlxzoDuB
2TcvGKM/PafPHdmCB6NT5bXungxAxFP++EbYamddTVp1iD17oeiTyF1NOg53hsvOvbfFwdKjnC0h
uNnUYsZ/l5m7BMFWa6ISvLfQAgvfgm2rmZ2uyfxTcu7N1vUtH9SZvgbgElppY0hp2d8pZp/qGxkd
lyc5M9R2GWwnXqR5PkM0HN/bXklA/124p4/uNyht+FOwdjp9D5K+jm9HH321cBgeBRXhyRD86QlW
zhyfznB/0W5KgfSUB0U4JRcr6Wk6TConOXqXaK2jopqsPb5fw7vEWi0WMxEPEpK0zRnj4/CMJSoI
pFTuX+WoPQzZLq2d0SMJe2Fh+ZVMuQ+WOVFA+x/2WM8iKoXxKgMttQMcPbFXLl6gXIFF6yAyu0tc
I6FdfwGsZqOmxRSiYZ4HSkuHlJsJljlzjKG0rXpUA0Y+abBqwi7hMgrajQCcSKnmFRpsgupMY4Ht
gajcpl8eDKzCalBAFmEr8piNDm4RuV6HFkSZSAC3epKJvM/lf73abQYdLxzZXkjYDGgvl5cVD9lc
syZP0vT70Ywafyja5WPMs8eFRdcHAc8C5a4Ssv7x0EGdnqlE00Wchm3bQfDGBUlShfsrSe25fPzP
RiERPPMjkyQcxnD3pE5A+qvUnIvz4FYRJi7WrYZfWjyBX7Ff4BNxzH+4XcncB6yjTC/tgBGFg1tI
lpl65qfRXjeBma7az8URdLpK/x6SJwLwRBHVB2C1R3V14R658rm5pSOLXofpA2k0l3KIIXquAHIf
3d6t6dJ01CutgTeBcxgNqrbnnq1GWxvwxVkIMuY0jQSGlpnmU74VIghagqaLx6/BW+t3uWRp+OKG
GeB6jc57nUi4QiNx9xiFY0xMRplfCZNtn8wvHey+gzjZQ9PpE+Oa72UckvtmUGr3La5hxsRiOEVQ
Y9lnE74OuVGCO+1t7ZVFEQM4NVe/DLbqzN4TS77n3vg1n48iYvaaNk/WNSf87jKbO06YQRWmCmmT
CD+jEHZFRLNJCEbSHsfXDVF9gP9mCHGO4B9Vr2wix6h+F2kaE2nQGxgTNgZqkFYi9i26OWIrE8rZ
tSlxBOT6QnDnVpZd23TqmdM7BiwD9NHhdEQXd9RcEQ8gOB10KThKI6F1hcVqw+/9WX5fhLlHgR4Z
m+Kh7GsywnxUifHA1pOTcEGEl/Ie2WdFViV1To81/VHqeyF+94B88DAgNyyyX4bUp/ZWbDLWDAUn
+sUM4ZNALrzFd1LXCO5usYVP0Ky0JeiTYEGufyIVDLamAJ3W92aMdfu3XEhaVBs2+aXcmZ1TvZ3B
0TS6CNLSFYFCnaU5/7yO6PmYjBJ0uNb45PPAJDgfiLHs0glRjj0EEbd/ikkaU6gyXpALYwrECIr7
zRqXBxj8cA76T8cxemYbPmIM52VEcC5GyIK+yyj3ClHJ1DYp9w1UfYr77zOWyzhLDerLlYBXtCrM
O4KkoUu/Ek+2wkZ1CrcjfGJPQy8n8FtG0cWwTkYLKCM30kfm7bNcouPJGG5zvXZ8ehEthJtIJv0B
EO2ihskQqDpTr+0wwlDZjhqD9HgsMTGCPI9Pd+0wzJEJmBRw2VoRf9T7yAdCkDR0xmqse3WXA+jF
p0dFAlTe9MyF745yLfxPDw4Enmj8b0Ja13C+N5PUFTo7AariFB3IXLwxlaLwA4ii0bAF7c5/UBBS
/Scag0wXE46sdSmSNUH1rKly5OjnA1CcUQ5BL+OPN00ta0pnNCHhHhaEwpAvj6zMHMJHDNdOchME
JKVQ37kPHyMUqlLI9ZoIBddWPSPeKkwDCCt8lX6u8YMQat/4z+p1wUk8Lw5JCfYaB2HWJQDfVgyg
rBxiUqkPlGtGM0upyt0uHO+OBl6mxkmCyNXwxea1blLFonETEZSrOwM+8Tml2Ol8jIdWDlHSN1ed
MAnhpPhLFXkbq/pvoU7wkPNhRetEsevb6iaWkh0OQNYr4k7CINp7zwRvaCMvNinh886JuAy5nhIt
G8UW7XCOl6UPqxYHrOlomI+wwwJB70VM9lw4RguQo1rSlyg1Ew8hWTRs7cQKKIdLf3mrpWFGbY6Z
eVtG0tuq5c3sjnEAl58wuZ9ksV+aXnnR3ww15FbaPZRAThCSToBUUKK4OEn3pnbkp7aVcO3lplYp
MWgcHYkmRmSNRYsfJVnxb0Ie8MqUHEX1seFdI6KMATREmQd/NS8UiWVkGqz1Znuz6UVw37SWOuQ9
H6H/67xDGOa/H5YlfUrrETh1Kb15b7QOl9JC70yyVxlCehBiqy4Yui1yxOKYNcFuOyyrTkD6WdF9
JIW0QM5KOQg01f4j4Ib2qnSAhh8opf/+FB5/t3hq7e0sPkquoap/TbfYDoyKBkJDlqjsHwlhX9aV
3eBodRiRgX1v5HRKwKzPz9yvU2OVs3rPP8ZjJ0DtzWTy73v87rXUDaP/lRsnRLPp//uGSBKBXadx
Lcz6MNljT/008qQ9YdpCx6P2rmBQVwGEN1XN2j9QzqnZqWUtRyBi/mM45bhYOsPu3GbuOIRhoVPh
J6nZnwdPDoU/G2jmEJlrh6CgLPZOigxKcrVdycM2dpD0lk03dDCy20S/I1k+sLN9LoIAmVacH/F1
4I5kUV8vjmsYxhYQAYTrPYip+rdnWo0F/kzbb6UGv9ivOJKfhz5nGlRd3F/u2bG+SahWBRna4isd
9JYw0vF/WjtOLnvyE4+RBlK5oYsD/Q81USSpfPVRbVqjmgNzIBbLznpOIOW7GC5yxGaKR/Yj5DK3
cCwfS7lc7vK/OV7Cyzev0CmA5VEGJTYp8ZALusLzSI4oce6LkfpHoTUHOoBAdUJfHwLBdGlEUp+h
cmqRuuYWqGQd2z/eZ2IXRHGcoWSRWV0wJlF9lNAAdIMK2FdDqjeu+hqXMysSBND3ZHL6iWGEviUL
vzAy84A7T89f9lcAYZehs2oBwEAA1Ac3vDSdA1eu67FduBKhOnC21kPGjQgoIa60AkIOCF5RCQub
Ya9aLvT5nUSdropdI1XTiwRR556pXvJ5J2WND1sqMs9Bpt5efN6bZ2mnBcYqVnrAONEatPp58PdN
5iWFpOsMQPFc/awXqGf6UaBc4jLrAoPUuCI3cmg0anxRKGFUnIaA+Zrq0r2vZjE1Kqi5TEX2zVjD
JXJDPwrCKOzhbvMXh6yKBryKyM3+u6dDcjS73oVVhPWV1qaQTBYP7EqkBBX9jmEO6dWKQdb0orgp
oEUBOofNJ7oVqeSk1n7vWK9iRLJ1hGBxGOvu2puOEM4eWGQ9J9Z18nSMV98ePC0WhtiIyQnrvmJT
4VbKGY6/WRDNe+7gKWGanEEpluyAnXx/xMeYRP3+/pzhHGSD+g4aoZpzO+DgErX5wrgkZlQ2eGly
AHeeJb/WmU5LHon8v2eu++3totNEwUrIBza/skNlSCeT28efzE7AWKTNn+euaSOhzQmtFheP9H05
mZ4xtfNDSUm4s21HnhFajkt23WRAWI3cgpN4+xt0HDpVDvdzmheq1oM7LftrPtb8xc2ymVylKBRy
RnBykQGyfvMA1ha6vIU8Ipbm7NdDCNvuK/zkMNx+Z3BlxWzBYlp5z9nHOLr/R24lKgwWsYx20l/e
5wT2iRyMpEbpAiAHrBjYzJ9DRVrlCr1dGHqQf+G19KyA03u0CaFdvVyfDpfCmH7YyP9K3//g85QT
1zD1pem5tNUzXlR/ngdXWmk7jb7qLSF0XX7zWF403Ene0Ponn/VY14cPezZg1aP17qG23Jw6YU10
8PC8hSBDDutRLTus+7GcLiipBXxNjdAgttNxHzNL1m3B3C1t0vLmfHlBIIWDTaxPzhTVPxQH65nD
+Yd4abWgAqWPlSzF4hTzyjJQgqo3mR6xZmCEUbwl72Y+BwxGNC+WJR5eKOEZrZN0qiEDTdnkEQYM
6sFqnFcqFyUk4xact0vnt8xadZi3vmUeOiMBuEjjGmkVez7tQwaL1YdUxEf/sbtZ6ix026RmHnE0
96DK+8qsP61Pso4fl9K10MQPS8NFbqB8cPNsBNGOyKn3UrGtlubkNZ4xXw7XrQUJArtQd8ndk8Zb
+IiuP/0YTZy2mobcEvSyqxsuM3ueQe862wFI0kCvar4uMzpDW99Ak7u2SOiediQWpb47LGUStDYt
ICiVcgK46YaKwLKSogTtz+25n68RKrBtR+vs+SiW6ARyadirxxp/aXULVttk/aPiTVidVpnPWxUd
xsKKg/PBSNdier23Yf9dBLxXPUCX0IWdN5SfwNoKJlzoa+RPz9MRncZDvUtwyBqGF9AaGmbQMaHe
iWB1RjGXJ5EXINWzFnOtQQ+E4schPZvf9Gm+uFg1qp1GzslanJJ/3ByK8MLfHUajFde58qaTvY25
rJpyv//DO07FBJ6a8caakuZfCJVE4lEGBv1tStMUT2h4T8avW5BaBjR9diC5O6qtxdAQUKka8ODp
O5LgvtpdUzfqyP/v0FZiHhmNdCuVnZ54vuZohjaphMQa/aPdNPpePmhgaSs1Z9zws95PCbJ6vyiy
LeZlriq4tcbJyA40vQahvajbiltcUILWe7ZVPpW20JtFBeIpT1qLnPcQfEO3NBJApovJKpz9pkBY
SMyOEukQF+6ARIfByzZt0qyfSm1IhZ93qMLbFdeHU7i8SYPx65Lvfl3FqeQ4IUzXSuCCQfOrp/EF
+eFS7GDj28ZlX2LhXDoK3yrN02LWEaAsRfuNUVEWkLjcL2g46gJnqHuh1Q7t9bLQUNewo87RlcfE
A+Ja+k17qFHxr92xnpg3WtTxv90JZBrwApYpaSfWTqZmJqeKNSwt8SLfarkqItxyAQpViwhG04r/
2LfWxrEUu9wbdHnZzVXXu4LYlsFnnfLw/ueyizWBlCRR55Z2LRc9M6x5rdHW174WaQCWzEddj/GJ
HqIUJc9V5q+kLQEcrbBpUlq1aR8f6ZpRWzbJPwEdy95APsmgNQzcn5xBS3UU9pJPL9yE2WJSlBeR
ZcXyPcDKtZkICLhjJjTLa/2uXJWVVnKLylIXBA/jfxfn8VzeKXXR5nTjOiGRq9iHuIfHGzmBnPtR
zDzZ3MFA1bmVudL/nu2Aj06BxLSCAZIEH82cPT43EZZamd7GckHtWKHunIwdDUzAc1rSLOnM3OIc
9eQwLDO+pMfJYitEZCY1J2vdpsOl5Fzy9gr2chZUGofIE9xNWexY9Dqy47vl00GYMmElpRLUahHo
L/DXrkTOlrHsv3mTmSG+f9C2HugYSMksiSvDNR3Fyf4feYX0BNoSjz+NUocddXxN84OQiClEFQ+t
pqou6lub/8LWliLGgWUZE8J7TWal2h1h5gVmW4OonSH4WDGj6lM4p4FfcHXl9GNaxCKw8ElP8Q2+
UMnlatrtbjej2fgvGO4BGOyqQFPEzpBgKxO2FIm73yeRhzDCBV95PIS9h7fnBcWJy4wvbeWujS4g
N2ScfVQfY4Qwu3sPuTx4GKoNpM65yfrluINfqBjwg7vbaGc2L/lXrxlg86bdU9Uvgq92/qIhqVXe
QnJnBql2sP52Fnq533BQdZ7zMC+bF3W3GLa1+6AAiA1l7p/KT15hoH5B40TSupsrEhoHnuVfo2Nd
MKwwFvMwr6XgFva0UwpMsQXxIwPopLPj4XDoZAwxT1ww1bFPyRi0j425L8q7lYjliZiol0labLJz
SQcby8zstSCA3Aw4NWv97Kn+VwC+iFQg0/NV1pQyV+Z4ZQ8enFFVGjNQ6FNLFL/oNOWepFZFp3BC
gL6hyBsoPAE12FQdy1ZqY6oq7HCId17KCFCZ20blX0ykiFTDY8SChGMyI2+rmvxlzI9uFOwGyNfv
jJDsq5GviCNL4ZZayjzSjBPvS2ZUi1yOmfOC7sh+0XIPG8cl24ZlHrr7lfxs8HlwNSgkSfqMaf6I
FzgOvUkGw1tgT67ezwjSIixTZJtsha+Wx1VfEQXjxJoKLhqYo5PUYC41Qfrka2YaTHFMCLISlgJ1
yna9srAGuOcjg+P1Gi04/uMCqJ32Nf0ITCoz86SxBYCTv7j01RdIwZZtGCiBXasMlvCJ88O/nf99
0OHoIH7+nKkbf1G1ciBTf69dU20g4W4wy/SGBCmb+0uM0Fk/Jx5yLp1C4nCO0B3EkQgrAaZBJ1PE
3tHSc2BTTwCrPonpoCBt+YX/vf2q34vKsfKb2QWzIk/ODyHg0Vfsim/jDehfNm6SCRAGEzScQ7P7
rasoMEn2lF8yEZvBuNVx86iDqJc2Qb1K5Nn0BVVAxDFhoC4A9+uHfnVpPWucG4QvTx/CjsCSNDyi
WHmDcIsd+Pr7cneClFWcIwbqpgC6dxcRSRlhYZbeBWmPt//sTmXqap8WttRLyeEXe/vmfkNYbJt5
/oob5/tRLF1PxS/tJtr+aPSKpHL2J1F8TWTY4vtAPoHsyDHXRshnSMiTxRETLugTIq1h4klZT96D
gph/ESqq9Jg0CJKEJ8g/QcOmkkTTnkHew7xKGug5Hkx7mqYN0hfDiedK5+zMvyopv+rCom1TTEX1
HfGXPIU+GaaMUU5qAs3UayGT1SjFc+XswxVmTHCaDTLQUvh9n89XiIznvABOSDqy0+tnf04E7XEM
EJwz8tJUleBPBxou4p5fi4Dw6SuTVs0I4wbesGwZtGkZ+qd9UtqEgRTZTjGv13LQBOE8OGmCFt07
l8bD/wSZZRrxNjAJ6MzVq/0TDxKUm5gIVYjMHmwesywUTR20v6ACVuSToQjAe8X7WnniMwZtK4xQ
5XiG87ELBTGDhoQpAQBtcmDyngOmb0pyELtCfM6cDDlJKfU7MXm6tJ3IassTSY7uoeVwogFHspLN
pRw2Xh5khhf4z+4JfJZwI3uIzNknUXOOPsGY0DC3zXyClUT+EDBjznI11nndjv9RC0eFHfJo2dEw
mZFEO310cBgyIM0P4lRLSe3g/egFeQ0KWG43PkhkrVwbaQ8p2bCpM6TLqOWXsaBAxI0o5KijCuQ5
h6UhrMIRzs2TC04b5T0U4VFxhJKpJ95R6pRu7uKX1IvekaJjeK+xVzykythO2AYCMsF+uvdw+UBs
wn7zmYgYJ8F3wGEcBiwXRHPpVezf+UqaLlz10CRkTOu8iB0d6SnBxynDYzYcY0ZGzsQ28/UpX6zu
U1HMFl7I7s0XyI+55WETQNDkoqzht4GtoX31rFa8p7TPBeGZ+3XbecAq8GmFjGS9I5gJ6vz7dKia
jDUy0l7oahj3JcCLbkCdzSlf4xmiz1gDOrlKMF5ahLNNA3i4QX2svWvvHeZvK3DtpkD26yQiX3e/
ib7AlQ+YZllnMiHf98un2Klz/qivHf2bxV2jrRp44s7zqURQ48dOIjbhozr87r8c7iyEQW2Jf3Qg
tUNVpvSIqN8yIEExBfuCzSZa75jhO/1rG29l1liRUtSU2rq8ZpPjk3YBVALG0LBecjupFtcviNPP
KREFEzfcIlQZxHup3mLILlCf8+fKLIZPHWlttuG/aGb1dnKZN3Yf+P+A7J5OKVCXtzBBBHKcj5ZA
YbnMJXczpiDH7wic5HBFgGz8KfiqQI9sblmWBCFQVI0B/ClDFG2Y9yHNoEGrguAmct1gNhLj6F3q
7PW6ClGJoC2WC7t5v3WrDQgpJGFbm0zyobuBQONxXoudXmqD0OiVQlcE0WLoQ6YjLqy9v/YObdeJ
Zg6WLPhVkfzxMG7F7Xgi+yd4HBJWu1TgW/cfzJW4LLwmiD4/Fek2ajFiJs5J2mWU7/05YPKimlnJ
LYwYrWsX1dCG2M8iMQtPwWx1T4BIGO0ACkKOXRPTGY+vg0ALBz/zs+YuaRlygovx5SyTi+gP+UaW
NlinV8x5CQjBJuCYIFp2FAeMg8JdcchUubB/f/dGH+sOgSkgVh0rdc5whAs2sLuBsEJE7FkW/lqp
yyFjF9cHlILmQH8bBCPItjhqAL0sv+zRoJsKKKu94UWTIiywWFZL9ANX1qY8cLZa2pNIUsu7HtGp
TkCQYRfzBXSrce0KarLVCvS9CAJL7AxA1dxxHW1n5mQi4+eExyg+5MEeYJHgZQoAX3oV399VfdfT
YzKAOUAVPT/YhdXhcWPuxBwvBOyWaojqlVqKfj6eQzP8QCyBMGPrE8l6Mnn0xkCRBq6twRsTDmtw
OCn0sgkqnpS4HgYW8AP2rOlNY8Ej85Fjq5hOlqCbzBDTYZ6ALBciXZuPRNrCvdY3+p0q0KtKdgvQ
9LH3oGoadgqO4r9FGkHtKoL+sZjnM4BhgUhyZoqF/M2Lnam5QvW1Eg4yDShmzsdT/Juo1JzAQH2n
Vwk6rYhjob7a4a7DxerxP+gUC5adubCV/Vo+QsvL2Mpn6GuI6DfToXB1Bux8P03JKLsNwyrmeQEe
K/zEUYF92aqEibDOrIC+MCTuiWJaGEZpXsJ/dxc8LbWw3pfYpiqoNgITlgP8fznWyGosYj5EWG9M
aMysNSXTh1SW/O5bZFGvEBJWggzvVApAumrfBO1QHRGEbG6jyfnDrNMhUVjqL1KGee0Y4ieJSltb
x3NvwFLM9EUlqXww1BTSvf937qz0BGiGYqXJxwk9d4GwWwFWl3be+gvnPWvbkMGFWbM0U1/quV2U
TawVZYJuOhVyhdPZvxYnKQE69U1zn9QvJRoKCJIdbZujQDinfsTisA274PTdIEr+Y8AfZAac7h+S
IPi8YnhwhA7StUFFqQ8twFiYEDweG+rn+xZAr8jaBTbJMOlW6vMRARUjghFPYBbU3Up5T0agyT9D
NWCdZmF1XjoFw6IKm5OXbg1W5HPj6nPlfTx8Qgc3I2h7bNw1WaGp5kQX0RZq3eEvOym6Dj18t0gM
l6X42drz6JrtZ5+OVa498281hCx8r7ngmZZ6ppJ1ujQIflyaXx1N2WRIN63hekiLAWuzR9Osb9/J
AJNJ+pXnLdXdSx1T5kxs7pqCBPSU5nWqFTkmLLJik0eq2NnvA8jH5504HdD8CNTyWuG9Ec68oJFf
o9qZHbFntVcdHZ3mgYoN+DrTjvOAiv8NMvWNxnvoiCS8m9mx1hAbHK6gl3pSgYgAb3xEcmlCHQ+Y
Jsx/kgVzwQ56k96F1tzhzPusOaYr959yhGUFhXHyW86Ga/iHQo5JMW8OXcNc9N6Hy0xqzyjrZbVd
sufXi30XrR1otmD6+mXnYTgbswNIDUvKB6l+C9mAC37ZlQdM9EHDRCBFO4TykWektPycZmx9BRaO
N33zvphAXJljzvRqwTd2UhIEfo0nauvA7Dix2gcmExqz8npuSzbDd5+Ty3K19KJj8zT4pZVtwLxd
4gYQQg0xrjLwF64tlHHnIkewoB8Ia3e8+Ub7/gMJyPva2BiDt4FTXxbESWZrzqwDSh8NHxH0XoRR
Zg7BE8ueYziFeakk1RpPvDce9x+tnu3sPrhb15Sf2WPp+A+IZYKXJltd+YgYkYii8EBmnlWK+VCM
zxYfPn7eKqBFV46AsVTkC0cc0CILWkjcARL+nh+FWhXOh0+4d2v1QvNxAt79YN0rxQwHB3nS+vG9
FHh07zXUCf5yFSkZkjjBUVNoyXFBi4btLMo2Al4QzaXxp7aW6zZkeHOMRDwdMHV66KuVIPIBTPl5
D8oZqHIcQ1jBvlR1Q0yG4Sg6PkABX4pzFWIgosdMhvKjf/x5KWU43UmdIrdqitAMBTYBIs+QuJGv
X1aZ/y0LpynAgsouYyoLdTcMxpBe29c8J7fl6pNhRl4P8rWL32P9+RZiQpXBKZawDCIG7u7LYrNM
hB/njgUqiCXz9oKHZc8Ce/iBv/HsiLsiVDMXDRRK/2POtUWirxyRlWc5Kl0WT9YVh4qn7TxXvlaP
H++fIBTXJJwjB6YaJA9MupJzoDaDyoeTqKt54Qpv3VgDDxw40N6Bde0rq5z2GOfQ9BIwtkd81xcq
yv8GCjEL7GIme92HO5425Ya/qi7FV9jQqbJSPPuyTr5O4VYr/8TaZ1HAXbcRewPMSgNLbcuUUZzl
OzkRKbAjVzwuoOjdvVmjXF9+kIzdQx3+bOoP0DwL/2ClEkYNIKbrQyye3ZWiAknJdBWyHGn0I5Jd
MsY3rniytE8evg5NSiQCRC+G7ftnffHMxp5eRD7RAOoac21d9kqmIel7Es60jp5UVb8wMJAkuF3R
wfdC4fw3cvWNLH/UozHLyjfbTpmhsvUonf/6GLEU7OPFZcv1I3ZH5IR5Fs8CcfOJg8OXVqt+Jud+
8PBa5LrxZC4BHD77fgdmAnqjmx5KQyuk1UFfi8Qs8ZD5g/lY+8+G09Q4ZNNx/OftsUZzfOIvTFhY
6L8esfx/ZnGi0QfFoJXvut8jCLYW8oQG+vZ/TAwCkSEedGAFVF1VFe8ad4nkTPVu8iPsNSkR4mVv
BxEv9Y3EH+tLHD4cZyVNN/D7W2sR2P+lZZ9xbg7MFzWUmxNxQ9SEDVySkGX98CtG/+ECypPr/jrP
QtXbqG+RpuaYhJTkP0/NyvL4pRxU0hmrvQtgyeycuSJP2wAJIwZx1v7zHCDDC+P2KN+uB+TOzo+c
f3JA7ywIsCDVwSJAHDM6G8KVbjstP3x3Tl4leKdiJBhfjbk9W7C7fwKrhnX5X1gXbZ6LAjJcy84x
JWwG0j+0VchWcD6jotlw6GokcWtjMwYcNCBrDOQRmVXlD//GtSiaEsJ9kiFHGmoeAtSAt4Yx/QI3
KsHSeIUS5V5VSKWluoo7xVPD3WPwfJsSUZEjgtiHY5SZoBEs/lOlw0k5X4rqfnCuLSNK6wUWCU2I
rp/8AmGvqDzDVJsbMG+mMNc0P5UhjVVCMV6k/lvJoltDu5gPvDr8LXdhGJYigSb9AcmK530FQpZL
W6hCst5ClxruaWwNACqhcc9uEgFCA1PFQ8V4FmbK7TjMX0pAs8y+Xn0zGI+0Icv3IkEH0YtpXCti
e6j11PfAktZ4n4179kc2PYYQu0VHM6QNojsCUEQ/v1msDPlxp1noetu8DlL/dkfubEYoEbMGmPAI
yggPqnUgDisdooxavZAXbW2I2WPUYgvfhdtuPJMAK+MJAV5RqxSx9L1Fml9nQ6QQS0f+1EjDxus7
pdjDCbIEhWYLX9iAwZNjB9codCIF6xXWEqc6nLLaK91UW+VAwg/uax0hotqRYhrCQlAL4xvfESQ8
xwdlv+TIN8LN0H23PU1Hfm5JAZhpaSR9U2PiSPavSDK9DMOhWhGTk4RC79inWRe97rZ1Sg47u20t
treMCAsCKG/a1SHAa0VTD5cJiBxpX5NcfMmvNzNFwvOUO4Eol7stKnezgHPPEbQnfm/JhEHC6Wl4
kkJU+0oyzRb0i8E4heFPd8egOiNj7eHlwqJvsbvh5pjHzIGVOr3IEvZjfu7E0VHObUAIc2j6LJFG
FvH/YxHCGYFTJBriPcEiwUp9fXjhTYDkSiJnNaTWnfNSsex9CIf4RGss/nKjhC3wnVYgz2krc0Tq
Uv88mwnawJos6/b64dax8A9EowConucNtTApNKjn4XwoMewHv9kpfDrOtGu408CfwM/Br9STtTP1
0fhXNCoU9OC2AG9zHUjNvb1xa7NvxorKz6kx5PWgNk5Bmgpz4uObwky2z6uWE7kFKv0fzzrdyw3Z
EcUzgJ2x2fVEX9o8MCvqf7twQ2dMSfYHrw1jrbDDc/1IT6nwsXINKzNvHuzb4htlNQDi8x1BJXEv
6O7wTUOe5MV7AdKAOpbOEs3fxfy/quXPNP+3dGADoXiemKLJjswwPUqI96y9yGXHxzzJvGsFDt4Y
rEL1rsC0NfAG7io8pqpDJl9W4jZ0LpxF1+9FWHNFaDGPj9n1l1nXVuDvjNAbIwI/115yZAPUyOMX
a1P5oGuEbj90hyrSs2hbecmepK7j25Xh8g9T8C25MDRzTXXlWjdG8IUGsQ8fLBVfd5T9u6vff7b5
CCGBGfZQ1evKmwbzXuB1Fuw1FKQDgMzlowOCjTeiqvGvz3GP3Ec67j2jXLOzgVAloXI3GyN9+JM7
Q9RYeyPuga/ppuowpTyesh7Aj7daqCmHrU+sESDxCF8JGa8HGZPUBnCRFiF0RyDyUS8e41NT2eAV
swAhiT1ngoqml/kC2yK4Y12/VaE1CYo13Czx+Pi8xpqsq3OtkVbu8gRPdOvY84cM1+58RRedpeir
KL0UO70nqOxxmFnIb3pqYZLu1XWWq9tWwcPxmSondMO10UNVZ7ds+uAvdkyPg53os4CFMrR50ITx
uvkZlWnVAf82mCutdPEo8Jl52qLQLDhQRNeRfaaTRHhHfd+MDLXVtOwTT4Xwi+uJJ9cPxf9JIhOu
fQatOk20LdfrzhOpnhF/sSyrxxAU/sRIenTUVt1Vbkp9QvCrZv7fqyLdd6Osc/yqSROq/U/UfwGv
pGr6Nb02wtM6Lk+ExvCAd2BulFhUHxdmLJizlut4Ed0QRYPGS3k0l3kFDHxrPcS007HU8P9Mp4F+
sBCcM61pdbKduRhZ7ZWM/3X4RxBOzguzMD5glj7ER1zg9st4Hyl7e+9Wd2pcM0qgv97qGwnBRObR
z2dj9OLGX6EPCGgsBgtrrE2RuvYki3C8f4NPEhmIpfgV9N0sAZPmrRCQGQSCvAyVJeNzINeZ+8go
NKCkDiEVhpFT3k8UTUOU7Stp+gUWM0QkL7erG0h0CqDoJcAppBDi7jHZoWM9YmTOFS7B2AFQRkZB
RHS89wqTZrySAObU4uvRYGUeV7Y6yK6NEjaRSm1WTqNjj7EU0brqVNT05oinOH1B96DCtbm+mjly
sbnZMMOPytx2oPonj+K27mC9mqXWYPUw8PwkJAjSDF8Ar9cC1GBuZ1YWoVrWAuDXs8Jv6mMwDxbH
uZXHLCKz50HLMc+MpiiLLrgmdqxXRj5BPI3K+LOvEHNa0asjQ4KGii548DXKNL3UCdFJye/WLdL/
LffvQ/ANcSTWudcwJ7Z4VIRPyC9ZOYRaKcwb7cxN+NocQyCEZ3+BSkum64UfRICiYOzofVrdhx7b
NW7OyZA30VLB0YIAkntCnQRaRdjBeWMBNJx0KQFD7JNha7q0Zj9DeYMQmhfR/TUTMmDKIqeiDLSj
dwyH8dwwx23r0agva0iCGyZ8QemCilwwu/qB5RwzobwppWwavipXJODvB3OA8es4SHtA1YzIpf0C
MJfWOFXPzKX25Ifp+JWvw6PI12u/1mKPHk43qIjNW0m3wIf/8HRDlkltjpb9zkppn5NjEZETlHNb
bp1T/UPMwNSxD9L/UU3ruvJKFyCnmXnA4Dqq2zmQ9kRxFNljH06iGTJBSDDCHTwoboCsu3izDgMO
kwPPHLRaWtfG+QT+yTlauuA/qJQfQxIHwdu39FlUqGpc3rNjvTQwXitm6AiN6h0KrdqfYXcYy66M
uh0lxilIxF+pM7zZ9PDeb7YWPRdO6TOXLEDliONLP1hDAOs7vsjneTIHEf4JOAHCKea0ak5ZmdgX
QL3toGIpu6aDA7Urz5NboGKLVmvv3NgYtLYMCneYRFQTQn1oOAZNJ5t98/MfLDFdSYu5VKMpRg3i
mDKIzY/2i0auxCxUHoBwQszUhm5EF+ut4WAvqvB4gpUj13hlFRa8rf5hvGPJVwayccy/opK+HroW
f5R7N+rByHnGvHveU0jBGEDYRvCfl3XfK5SnfDXQHT/hvKvsyz/oUfK6y80OdQpeVLfMh5IFK/xm
ntEosl47cVLRNNzzHEWyPHIxkbyWWZe0QnIbekyEUkFR5U7Tc2vD4eH1aKnU8Rs1R94Agy6Orzpx
kESJ8Lr3ZcO57YqmyxkC7SeYujZLHAO4DxAa1nGWJFLtphYZrJNaBmzJ3O78Wj9+p4cyhyUfGXlh
JFlUN2Dh0OMj2OvVdlSBqmSEMDeU7lfO6fOmRqRTGHBXhZI6sssK0qtxyN583quA4t2kSH2Q7/uP
2wJljmFRdbNGk+Vy4XAuycNL+JTc2V5LVSQsNs582WUWVMHS+SQer6/e+bocSzOyUwr+e3A28Rae
xGsNe+LyJY4p/qgAK2qsjUFjVuOoe2sX6SibaTXrC37DcpbyL/cPuT1/+0sGdNfrna4rVKAX9Jzf
bzLnB/BsfLjjSwCl7IcoRtuBHjSwoHpy1tmqzeNv+NOl5KDibqy9IJ9T7Lvbj403eGkjB7dn2OrA
EeCoht5GlKcupEPEVbItdeXc/NDzWNdyTEv0vld6raW90KyX8CHeUAn/qo7Oag1tevHnB3WOVxv9
jEyZquG4rBr3duLqkl63iMRxKb57vhM0D+Vgss5l+NFxV0QZI/XGaidiGQJA/iEXDinVo+a/ivpu
YbIH3zQxf6oahDjsYCOt3NV1lpo0iLSR3HNzPn+dpkYsBuyIQd1TwyZoivZiWTgaZXJHG3+jz8tz
iIM10nDVJiw1BvBYZRUrvQ0Xc1+lv+FlMU5P062Rrxkp1pF03CpINcptjpoQKwhAvKeRnog+F2rk
fsWTA+v0hDlKzf8D1Xcd4XqkA+DUwAiPcuuMrfzPAsamuMnTeuGeF0rbfAg0AcbzZdjlzLwmA2bh
imJONC6sMBGDCdEyAG6cI+mxBqR9aOYeYnH8RAGxFh0tpPYpRHQKeCv4aQ7KHTsVDSshfGea/aSZ
r1Rn23LDyCUZHmOHbgKIsxY3Lpe9WKsUyzTXOFxbrvaa69aL+OSBoNi+dEBbrjhKMRua5rk9L0JD
J/tlkj5ITpKy9jTOq+4pVuGfLtEBrEKXURkzwl/QpNiJ6uB9hYN3eLk14zDa/jhiojaAEMx+nrTQ
9UzojKzRP/5usw41W7OJ0CB8lHK08fRDENqea//Riw3N6t1giO7W/IfxUAkKHt+MVw75DjL8pZvc
Mcb4/pJ+QMxLSS70Rcq3s1GhFQFRu+zASyI+PXKDE2AOFzc6H1Q9pAGux12msqcQVH2L55IDffbK
u4MI9OY9zPoXFzjHzaU1I5GTzKgL4UuIEnXeVbQlN7LdxgFbD/aR7XCkbyg1Q7Ocb+Ae7t9o05P/
cMqtXQJENKNdVMQlMDnuYmPsyNmB7+hc/As4H7i650cC9GWRjqoBwdbEHIMn60oTT43b5xLDmXCd
v07Cuduc4t+FyfuFCd/ODZnK5/4gQJGVzimbUGRbLopKX04TyMVZyGU1P1EgSdDB+YSXVKNc3ivD
TIEqWS4kSna0xNvG8wweTsUweO3NPKD1stB7VdFix14kpApPfGKcg1X4alGxU9E4bRxy3BrJq+bE
EDz8Nj1vznNrGtc1HpJqU4cLRYAPAHI6X63c9jd6wBa2C/FkG2feModniFV3XfDtOhfH8qnazura
8WlRXfldxTD6wRv7Mf4Q/+Eyjui5z9ljWAoGJy5GvinEUWid71pcwSo6kcxRDUrb04pOGpwG5ImO
+pcPXCxbeNYnNvrRdsxHDRAT4EDk2I92Rng/xpFNq25MeErBkVP3CzWCJ8NiPzzxHQqykn8B7QhF
HGMz4yru116hiOLFE4ybibZwlIHqpPTeWpcmLinnQxIEezi41o5/XGa5xKU40CDqdzS1nJ+gUP7n
l0WzFDQs+SDZdc2NrEPI0pNgPolfjBKGvpe2Q8UR3F7H+pjhJGtt5LnOc1eN7dSIcbRIZzVtAc+F
4YsqKSqHxs2bXhwIYjjyx9JuEMDIn3sE8cyfTiT6Zd2MZEOslMDmaXW8OXB3f88v/1/TeUerAjyD
GVtqcjQa3Fo+GRCJ6Ba3I3Nmhx1K7+pqwhvxMoBt8LRr3OHdBNm5j5KMOWYjCK9e5yb72v3X9Sdr
53Eh4wliF9SmrUB6ovS06T14yY5V+htIgIaX3GTvLQGWeyZ6vY8EvULAY3juXaIR26+h8Odb25C6
ebSFyMzPmR+ock3l3l4bFHncCe9OWtEHVQJrs3xkFsySeFH2u9onhghC0J89YgAd4wjRECKgBah3
DG06QtRjiNfF9c/9oaCA/3rpT37V9foYoZZct6zIMWTvB0s/9wtbHGRUuXOsuIBKnYXDGiVW4VjB
RrAX99D11qaGvKukCkbzY1nGQ0w9rTOrR4m/2hSDSu8pDGHx3eWroFsdI5ShudZNFSmupb0QNVAE
4/buE25dFCtR8Q8yCOyvfieW2bmRpz4FCobbvt7wYM5sn2WpUqnrXL+6PcCI2axD/I4Qc1r0lu9d
E1AZExZtdbal33k15QVxF02zlvsPTKiHqWvkqamuyW/8qBb1JYj6bBbG9mrCLMJrRpc9JoN25/HK
x9YP0DVcZYoQ+CP/toeqF3hF1TAmEQ65BLvXogE9yVf7QMHDjdpjEaEwiEJYsDPrE227Baz4Zi9U
tViR6BIzYURhm32Y80RnGVjOMh9ATDA+LgcKLToZuUw78glZORJL3jl2bpZuCo+wLQMUtLFWZ0em
xn6Edi2lcLp2P3XlteQfwe2HVeh7EkAUXkCwrgYw7N3xgAy4yc8zwhkQeL7G/86IJIhxifB7+GsN
Su3/KmjarVhsI+Kzhf58B5HNLNsWP4KFpRsjtL6HWH3Cze5iAdi2RzlXlXO3ddu9bBGb8vOLm0N/
6wuSIhlea/5+mkBO0YYYKDwtLyuIfhYIOS2NwEusxL7IbFpDoyfL7yitR0++tUipOJZitVkDmhpr
A8nFYgsLvpjOrND+b/Bf9GE5+rsn09v4rbrnpDrZGpwbe34OLIuNBREFepCM0jYil8HqQzDo/cB+
saA8j7LIiaZ3Cg8Xj+MgGe9yO0p29fjoxdqR785YLiGH3IN9SSjcnVKFizUBS4Rz4JdLA4OssPRf
8j1k5f3R8jCVgGZ8dwcDQ5qIDby+5UFrLu/79dE5QuJxkjgkWrY9FEDCG4u4p/IhSB0Hi8I46US2
PHRm0J0Z0o5UrA6+xwqxpCUpGZs+bxF2kliZNrOLIuMeBfhH47wsW3CWybcPfZyLmRYT5QiXH6Qb
WEIlQw333KyaKZwNR7lNlrsoZv4qbRqR1I1JxyJnN+dL3u3RMVe9JCKC7Hy8cE6MmpLzys3jZY4L
6iJaEtPkZ5Br0/VGRqaM+PfffzK/JyW7yoBvLCAsqocrH3HrVzWdSpEMCE9IXLHydeQ0l5sunn+S
tPsPHngAUn7s6jqH45j50we3I2IUQ0bkRSnAeUjKATt/beeH21EIBh0yIwGT/fYfJGdcHPbwnDCB
Knc8Uxctr/DjQaZ7PnlHho4zWYigyuRbE4A2wjp31NC92Z+wl7t94YfsiehH7i3AK1zldKTHUVVv
SG0V1My+zyj+STHu5TnxHBvl685V7Kl8rYmcFRh64iPb5+mdYL0VeThDGmZQMNI9ztSnEZ8vgk5p
OreVLZXEiZcB5cL291YT6Q4v7Qo+Ekb117X6xyeMzrShpBUesV6ZBnVFpVT4G7nU3UGDVm8Q49eT
uiwPK5jlVVW5dsiWdQuQ+ztUtERkOtdxHxoHoc/W3vE9apB94HIUZIYCushPqAJSVqYNnluhu1vh
k/8WbvlOK850Tij2akS434XQjsSa1dziSSilnkpLFgJ/0gxANrdvzd0es+6xgmrvhaoPy7nmf+4L
cAFJajT4zBi7el27VVTftf25bluD3BaYvD9rNZs5wJh6/lGyrXhGRdzwM2U1JRH8w3pi2NMMBBeD
KZpnVf5+q8wJrEEDnsN2bJ4RrgCB5isFEnK6N9xtmaFqlexpIsVHBkBQ9gvBB/zE9YTNoIkHTPW4
SwycBS6YeZ+3dlTYtDG5BKbiTMoDReVKR7pcPJCaJT9dY/b4C6C/RN4AJIQB1YRDHBXmytCs+d+N
K9UI7nw+LMUzZFLphzG83wotcXoxYiXbB+auQ6IBJ48NPybmkU8N6tcLTIYjyvbDn66iZijk8URP
+0BxDADQimnzeAWydRtM3FnG1JYpkH26XIUwKZz9GBIo0cKZ4uZQVxSVTCRhjRvAtBpmN1tcTWtZ
TD+fqgeuWxFT3KFHProeh+BFyjjQ/A2Ry557sXRYmm2+7wB/Gp77ZOhyLoUpvD0rgAHVZVkusoet
KIl0MtMx+ponzYEmwmgMKn66wkngA1IwvQ+moIfLyc/cPQG5LOpe9/Q7Hpxq3mUbEEyk2JutV09U
FgCtSVpNNIDMU7vhpjDKxOl4YQ27cJkVGv65lke8txf0xJlxextY9PDSWObVfC8L4i+wsIRc3xwy
Of3mjFhTCX2NUREOIZI1iB54gaMEwvKszpsqF/VGK5/GKa2zkspyeHN/h/zb/hKT0xlX3BXCAsca
Ei1ye7igPQQOQ7t25sOBV3t8mROLgsgZUSbzBxfD6vLnfKF/Afck1RPQg90bSrSqKRwzRL1T+UYP
k32F1M6ndLKYaLBCQDpUDrGu1I7zXU7VezN+pIfgMBVilAL9UHYLnqddFQ5LC6dI1dS+7rwah/JN
c4yOC+ShanSFcDoqFeE/v9MJ39oE7zrWdbbBvwplksE/9T+eSP+b9LeJsGIXAjVH2AuNAQQpIw8t
fXD9AIH/SlzsCP7cw2BvAAL1sG0wKY7r4dZ7lEz5bYKpINS4MhqsN1vYY64nKYkxsXP/cUbe4hcA
8cIl6ZFLHyrejvdfpR87mScGyhnDCNW6GtfwiN53GjLtDSKia72/XyeKrHTidKpM6C4iRa1+lkAR
FD3UtMnJw8kVchGLkh3a2R4UEkgFvbxjleCppVUiNQJ/g5lhwIZSfhRdVk0sTIW87NInh8KrjDcA
CHA1/46/SYGZnowt4T2OohXz5/F9Q5/TV3V9DLdSqghu6Fje6Uv/y9nDFjuyL+B16cfOoO9E8jpN
mfLAQDRuDrVaBj4q5y0p1cWHA3tmhvscVrMMztkzF/VAjdNJnMFvFmrhTfl9tCkpbVghGLvPTSFA
dnU+eiW17ZGucs77Kfyp0uOjUcZsPw/bMAnHThpoFRuHQp6ZWrJeKvJIJDZEe9nMpbFIWN2Qdyg7
V+5/PjfrdNPnpdrQKmv933kTzmXGUhuRjLsQQ+gLojwSQGtm/Lt4Sr60fxbu0vLemSC+8evvDhNn
wH++SEHNujRtIwTIKo32AzhfRCAZlVAW14uW+iWhZK6uYLf+sNFKb8tFLSKHgozI6ycR6T8RmCQi
NdMQiWMJTXvSdU1I8E7CHk7Odw8xlircM7xVaE0rOqoo6BVCtBI3froqPzXp/8ZMnCoG2XD6UopO
MPW0/obNXYuGFvTNN8ej2MG3+jM+EjUfbH49dV7rEMUEdWx5eJVb0N2Yb5Tly4jMoUNx7w+iC5es
rhebOJvlJrt6LXxUhyigj4bwvyXPoQztXu5ifOyWJ19xiwxxNQXcxIdfcbFTYHJYONG3yTA4KGAn
y8hpIjnNvdgS3guYO01BuMYB7RWU92++x8fHgEMIrWoE7SiObAEggr1TdhUjdKKavTfaFC80sw+n
kCBlMqYhdIy1nxLH/IGaltdrmiOiQNpSdg7V0YHif1F9tAAMRtwwzLJ+/o4r4WLVC8fVzhoJl9Co
FX+WgijX2M49inOqJZ0t5UMWcKwz4DS7h46wSP9tX6/Bg4AETzUTlFgEe3u5EEC3qKiXOflB5krX
GPZCR4CGNWnvCx2fTorv/JVzbriIfDexW/Pz7OBfcM1aq4N+lIloA6NIkW1R+sqyKDEArUUb9tsQ
K+wixdJghfM3osz5ecsPazEHJ7zelsMJBIBJ/wBo/bTFFtZS86MrVTwV9+MoWamG2hpHQiSobpat
T9tCK217mqZmKz8HlLbJ3rQBN/1ZbK7JxnOvatpSmYeXlxtVKX9FCg2jwpaX8t6yrC7O6KS0RWCa
2C40Qvxc0TKW1v5W7YpvAW20Jg1s+LldEqhk7pAuBQi44gpudnDJHKG7gFqBKEU/na0ysVtFK3jC
ZPtZXXITWBqAa+aDhOG8lE24UhXPAA59gpJgNwZ59W1RtWccQy2jNp6o0D8GDK4mqq8zoXFL+jo6
5ACPc/C+CMSWpts1UeroxaPGCIecprgAm5Vij3gFIceZvotLR0Eu9+G8DUgijZoknVWXCCLbmUM8
ENsOE3sou25lCLO/YvObOQUU0Gj58RqgPWU3KRaDcQLNjE6DJndib77EskoNurXci/ECQu8u5s8S
IVDvahMeNRRtvFUtxuxz2gmwyDCJTiQSrDpC1BscsFox+1fEDkMSa3z8iATHHnQDhbClfbuiLrlZ
EN9DiFYV66NvjpOAVtPBOriGujhHQRATkptKgjSGVreMH/JCN6ZyJF+hb3YY+raLIwNE+AuAUJiG
9kdacG1dsoDl/0ha/GhEW59IXG1Vhz/9hefZNyOJ0HZ+qGP31aVAlP8JEiavscnbmteAzlupe06W
FQ66FSUw1fVO4jUwrdK84Bqr2FOhov9Be5tw9PRYV7PS2TlJGaF3uZFBX/jXpjeKyyuc86g32iFU
GDfBewUng5HlBf9Z2K2LofjIXn8cP1g3WQtf2LqsgRM63ldA5iAoIelbOz8sP+crqvP2uBHIh6vX
F4nfi0qdV7LCiSwSk7Z2Wm5gillNRp6GKEMf2LOgsz8mjNI59Ip9IE5P7U00Ju/JCBgAnkJN5SJc
Wrox05gwbKupx7XuKkFobroniE+31fg+2RwAzToNMUcqXEBBacDC374Dx49wI1Egu+XdwJ0gI3ay
lO8arzc6j1Irb3nfaNHGUIx116eH/mELLFrOksfXdyCr48HbF6zGuWYZ+WseS/9Q10cKCLq3ADI1
Hw5jW+WAr3XuGDSum5GVWEVBpc4OBdLsSJ21LH6f0sbN5P48TcsW8TjhZ0e40OiRNCDwfZRpW89o
oJ79AbIMn+tC+EiQbc/u+g9SRlF9qToOY/kPRbvqrsvtb1AaWl5fnG+tqeMYg5TY+i6wrOeiTyK+
6VqiIUYTZGdXpnusPP5auBqLBiUsO4lz+VYYL+eES9rq5LY4WGCRydj6BqfyUm1alfuengLD1sQr
L2y8ftYQ65bp5QILWhe9bzbqzP6ghY3fdXDEkTJb9I7unajPtPstP9fxkHwB8luZI8qomEcs/lk1
VLjGppShfCEyK2HWJgHrprV4vMeOO4j2XHuHArNgdjns/ADEh5V2TmeYvcRIDMfPoverCTy1LtLf
G4CoTzMTH47zBIik5N1mvOjLATzqkv4TsyfSilmhRJUD+Kn5A+D+qPvKx25gefSjd1JUyvt0XWq5
LU3EyABW0zLCibrZAcHmdL+Ne+2bDvyKIpHYyLRSkbaPkRLs62Na1uhi2rErHu1LRxjjswH7ABOE
3SqhuSuvQKfFhAQVGbPuvUtgILM/YdVKyKSvSdyyJM8sq38OyAtL7sjsMRdbAnBCCHcHmjYAEc98
DvVR+ZDE6Ud7E5098kn4vO/DTZe+s58fClpGOinTZd6O91LoCO1eiDVd4Qv1RFHuwqIj8AGm1cym
AcO5+WIPQAmGHSaHkZBxdgbOsI7TMj/VG4agF7pdQTpboYwzIfpW8Ppq4qRw42ucsuQLXIvyGXxR
WDblIHYSKcmsoUVbEO8nChlCqemc/RlRND7CAhybncesJGjv6D8BB+XBPtjUBiFjkz5XjkkB4ctb
fy3OeKkoCZq+nbZ6kIFN+CfLh2VTc8i5DWz/iej0cC7GV8Mli/tof+6e9Dg1jzU0c93DxHqupTDt
nZeXzDdW+HUNbnmsJLUQkxSNEg6Tqamc3hqkJyt+QNbN8R7SSs4zj6vum0AAT3RwZ6AmH32of+vW
CV7vnxT+h2IrVRKcix95Eh7xXLXxmtS8KlmY+dfQ4Wb43v9Sd2fPbuKv1dI4SU/r7plM6oWLXJjs
y/+BbPTcefZUFGNZFcUJxEuGAWLBjjNw+1VKRf1Y7589SZkPjsddtuvprhA+GG2n169lZGWWcuzo
4qbgmjSRJREn6LKl43AU8RYB29PoExp5MW+L+0sxEfM41gYcErGA7zo86Fo/gqzqmi7EnD8B2XUK
7Ykkqah6OJmqH6k9sFakEU79kP7RPnyGMQnI61v45xoDbou9cYQs0jbAOEOzC6h36L7Hjraag/h1
LiJ1GNV0/Vyp/hEik1D7FbXM1eyE8LjoVfkKM/2SObsHEsIzG8Wk/lMs995boYku6ws5uwGs1Arx
eLYEb/iyErb6ZeZFfST0wOUBovhZNLr3OAFHz2dHdhOeD/s/cLh8yBDlbDSpek3jr1I0wc5kq1Ah
vZ7QrXJqyG02ZllBK6ehDlS1hxHf4C+8iopOFodqFEDXaUqXmNQ8DXesXwK8luTCxb/D8hmcczXM
1ZxX28HDxkOliEPllOjvfekbbOfGMFHDVh/ti8ywZzdO1WAwjqg+fj+4FsijmWdNs3q4Ik+FSQyp
DVxZS+Jsfadh3c8be1Z1S8GPBxT330QN8611x1syhTgyOqe1tLCRkU4D/WkGDdRK+eRiNk3xz7iO
UOc4c8v4CsfJ01lEhkUoU+eKKdue3RBN0N9Pp/PA2pbwE62Ub9TxlXSRB5+WmmhTce0ZW5us9J/c
voa7ZvzWnVY7So5EHE9bVK/TCG68Nh59jNbM5W/r163twKK4a1wE05eGe4HWF48oUXXzFvIdY+Fo
l3NVReK10G0s1v2+RE41GmAkolCUWAWPM2ROgkX9xc9ja6gfJD7lehQheI/G5jnb6Ddwe4RdS93W
w8l0RybtPA2IgpaYe6+nZHmC5O/YC0+0MbLO+57MSOb30LmDsAQVa9PoxdswaXPcaA0M0FymrEDk
KA29Ul0N3XQLzZzpPdpwomYEikS69ud7tkGIVa/MN6r0p/qjak/dp2ZSMjcB1csqmN02jKhFjI57
P8VUE2CeZR2ksXkQifmm/2b9aNK85Y6Ejhb5BpwyyqUtkMWkI0ZLkp41wklb5C6q+l3/vmFhywyL
XJd2p/Nl9xyaD1QtGBJ58hSqAtstHx0icWOTE8lZnmkwjrWhsdQnpq6Vpu8jx80fxol+8JmTp/ce
Gr1VIJGPFt2womNiJu3lK++YW35qEDT/nmTZi4EeB2/AH646ej2ecTxrWyUlwkn04Ne5Jt7rgPia
WWOsOeGz/ZxI4YtBi+FdNX3OcyRyre2u2vtSalxu6mmHxwE5f3LrtkHtMVw27aa7raBGaGsSFBOQ
GwWDvDmGzalXNKhm3etwgGXNdIM8/yL7MDbDJvyMewc/z1Jp/RBjOAZXdOgJg+ts1uLJc4UT2vAl
uyMdgqOTO6RxMwt8OPoVzxajfU5lzc5gkFOaZkGlvs9J3f4dlMH9WycWVPTeZWUrhkiC8C2tXf7h
a0V2W6ZBPmlb/Ue66jM1AkyN8Ns3ZEoxSqxJuc+yhr3/uiMoyuQF0RWymbGqhztT26T9zCx7+noP
+NupSS5I/HZTo/aayGh0UzJDcwXpZSiYywM1ebledX9Ojn7Bt07B8cdq49nSNjhuB7NCGb8xNPSI
cXYlacKc6G9UlGHd20OzHahgA1fR59CTqc6JaIthc33VBI8ZPXk6IKGABnN1+8sXgI2Ioab1J3gk
BMxmlJx0TU9AJyCKiWnI//CJcMahz2vnNqc9JmNXF4+VJAjKwdxgQ3gViyNM95uU42pS538nagsn
ydveWpDlU2UWhV4Eb+zEprMnIzt63nBT/qWEVg8I5USqguhMGp4mHWa2jXN/rMFF9Z2CjfcczxZK
qSGrqu9UhXoPk0an+E+pRjbkbag37myAd31l4G+flqcc/t+EjXvS4iZ1O40judSCEux8YMazrVR/
2rUIeFoKhKt4ZCdZ6LeRS6J8Bhc7uFx6e7qK9Fe0dZPx41MK4TcDIEEonBiH773fm2FMijyuaTuV
1BAo4mucy+qVW/JAl1fS3wHX1qk5hM2MMkTxSEgEbmsnYqIRBt0ilKfWNtIaarlxoa4jRqW1PvyT
GzHhkbb6DkmAf019bfWsETdnkZjMvbWDQMsIa+OGlaeV/RUe5bzLdO+R+JSybkMUtJS7HRWgkaA6
sDSRHekDZ/6k6WDOC1xBEZDX4Raq+s0oopz+QxGFdsJYDIEERyiBspT8mcgVYCzMrnY/EVIjRFZZ
kiAqyUhnvGjcvuT9VJGHnZ4kSLviWBaSx92uuSaiDDe6k41oblVi6awkcPLASyXqrNGrHefouNXq
FB/KE5CH7OjJuqLfvpdN3QoNA1vI8QTCsxI4lI4IRtvwW5KGadtRJzFVZwzPNZV7TUmSdRm73StU
EXOZDgN4FwFJhyco1jlDSB5YsISjBFGEawIgQ6WSAY2C7NzTZywYJwy1w5tL9Sp6LN8/bdQ66ICm
WGLNU1MzNQeGOoTi2jftXhVkzAf3VM2vqTtHUlae2M3VekwzlMFsnp0TAzIDCZpAGcZ5tXlojyab
CBLybjHwJa4OfHrvF7Cdgnyt2QlWVB4BWvDooGOkmUhlFPmGzbIX9Mq78OXvVKPdoCbbX2QPi/lS
IYevEJcqi3COYKN4C1z7K4jb8VKnzyWKw57wVjY7QXQt32aCqskBwVKJ7jg6WzO+LMx2Nz/OK8Zb
iX6E3ijPs1Z527KNoWxGOvS9w8HSnmaocEE6QwwqprSvB0cYU7+2JzbHIq9+C28k+F0+HvoFuCzo
6oUXGtvgtqRkqKcsapZ0IbKkb3GJMpO8FxJYwc1Gqke4MislA/DqH3XB/7ZkKSjIfjdtOxwP98Ut
mUKhX/l/ukRI6IBDl9NpYL+0JJymS1ksVX6T+vY9WbAOV3A8FBb9Rrp/3fDmlJGtDOwuOk7XhrQq
HBTtv9piOR+RHF+owUShNa8b3PDoeEUeqX8zK6jpPP6V4ZUq62OvGuHnYtpHYvV1vTmPgTpD1Dpd
AssZBSnaobqHyaSymyoRH/TTcTJ3PjrJgAkSJg7EyAwwCq5uGe3spWGg58hyKi2uBgkuBbmjWTQv
85xOu9t+STYdUkUQjZql/MyY2Hztq1/8gRGRu+thcOUUDVhmE8JDhhlAxda5LktY+IYH5JmiliSM
Au/ECWrpSUTbPS3Yw0FwbSI3i6qTYImHARaPxXKL3G9x7t3U8snMBT5kBf8TOWS33sfQenkcA83+
Q3C1E5Fk/m05oMV+cihdgGbnGNQsTIzETNhxfR9Ud4KWZsBNnqwVtqc8Y2oE8MdQUvbr1NThP+ok
furoPRac9f0zleh2Um5n0i6ilsbl9ni3DRR4IUKrXlgYOe6Dzt8yaBiHD0i7DwM3E2siE/7UDnhr
8nEaV+6kzLrSpBh+ZYMgUIzsXyH2SbiiDTmMaSXXkqEbNF7h0twoEUOo3Yhzkof8AOJd6gn4SuNe
ZHICDcIzDUAqnDzzfPKYtFoqaSnOUOpdGT356OttwjUUdPGbnJQ5t7PT40clVg5hYnP3un8VsMlm
WB054Q9sFVSg5L/bXVJX2/XgWdxXTXM4VneJgxq6fvvpEWkppK4UliXNPfersW7XgDWo9awObGZb
ipFnCPl+7LOIT1gpy6jI4aeZNUWh2f2ZPcr6b1eQPoghZBYq6gnjzoJ64OKDJFRorl/kRxM7DwYH
MclCqIRFwJF7t/r5i/f/L/78WpGYPLm+tO2lif2T4smTnWdyuvBRR1YYHd/pzBJwtuO/du82Mp/R
o4GOOXUi4/mEuoZNpOyxCsr+cCR/wq7uEJLYahc6YdNWA+3KIzY7qpYKFkExiAk80f7u6xv/ztTs
yHNuNbOjRMOvTkaRJ9U/Eu1qq7kxsQnAZ3kMXGfVQXxxEcMJRuN2mtl56tuKXbx6+yZx07NCXLrd
P/haPP3pnD0asDwZAI49xs9JwDEkf4LS60iI1E0Sa4Ynw5DBEqT631692aNEHmldk3RZIVCd5vxL
F9eRmpf6I/xrb31Ut2w3X8uaRQ6ohVMPdzoTxCMGjZo5JXcuuLrqjce6AMf6riQbUHcD/srvjjwb
BACHMFXG9/LtKI9OTlRWlRuPIoH/siO5HVpE7UdhgthxaNf3VvzDFYtlyHf2Qx2WLn7G2GjOxJPz
38daMsIUH5e+plQL0ZlB0DqduhF60CO/0f7O7QVrfBj4fgla93eN4JrOiYKC4kghlnu7yCp+9UlF
sNSyNxcWM4Z+7SsEfHLvw8De6GjAXcjHr434GnLCIGv/aOyC5NM0/uO2tasH5Q6lr0MpT7PouqFs
9ncwylmfqojz/ro+Lg71tMx+qucYwbFlSu7N2pnqyi4UvC1QNIO5w9AAxHlNgHTmftKh4abTyC/A
70k7bMErT/Pgyv/dv/tAb1pzrmRPRlEMtrCNICIqV5vVGWsjaSItThCJE+/tVPU2OmypxB0P4839
XtqJMBBccimiIcTHIBRPB8uyl2Qh8jW20BkWwS0qR4qfz6DVoAef91HpNhUiT6AH9KRicGBpCz+A
2yaRXdSwrCZxGa8FnDvlbC1Oqe4YBNe/bt0x2rxitSJ83TIBeLNfg4eZccs9k5tZVNMGh0+RydFd
+oXOoeEQLYysAMiEnFuE1K3F1Lgt7+9HdaN+Wq2uPBuZACmaJ6iqLhOsIP9YMgCXOuaHljlEDbet
VNUhbub7Mq+fZtxtki/rfQQwG0ItqnpkKnSA3jezu27PyyCehp1bsgCOxaYmj46T3OZUDj8rF67f
i5Bh1ydCYmax+lwLZEofn0mX/r+nS3/HRdG/A/i3QB9ktJwwBertw0hp9nD9HZ9SVS6pXOs0z803
Ok5fpyxgAx7R8aAH6vdjsVIqE4OT0KvsetoRcPjvyoS/Fxq3h3LaTe2bKBk0+MbJOYIjzpZgHQtV
oZw/X1EOVr8Qy6vhVxLcqmkLA03MY+qmT26G2SVfrPRp4Ob4qjsbs/jjRITuOdkgLaRFh72m7yCN
Zqc8v0yA0paEuauDws/xyzylJBOVEQu726ipdd54oYK0uqsBnO9FytloXcFJ60EHhknoOm4T4S0m
JWvGWaSxKtxechxRxdlsQ7vRu0OITn56kT30FXxrJ9zh94iEltG6dP7meoVGaNg8wBDJrVJ/l+/N
LkcsJcNAE7QazOeB9XTBTS6jnY3KVxipr7AGHPYAUiduoGwwrKgIptQ2kYJbfZKbyNt4wnWMqrAN
l7Ku3HDQBIhKP9CppOKGxfEoO4q+Y2tUzx36OMUpYg11iL1ktfWzLL4LOohi2dWkliJd8uO/R+J+
vsgVFL14pOIQ7UNq4XS2IXVZ438weES9qc14ijtyrJ/6ExYZlcJ99qxkxUVG4/BY3hMBR9QozHqY
Rbwpmlcz04pPiWxu9MpnXtdrvKJMCsgSLSxsL08aynC/K2fWl9vdNxzKIpMrGSN43lp9FDyZy1+M
bwtvUWINkWf04aVMt6cHArqWVAndckDJyYXTZ3eNJmXjbGV6x5kilrZvXmKKdbztRbr3LiBdhmmA
BMmnMdDBAg9uKx8NaGsq8rt3R2Lr1HBxbty7U/rxJFSnZ+4WVaQMftA0zKlPkQ630ylnMvwP1bzC
3q5z/LjQ4sSDsyuZNkQyUyiIFkz1AFk2mTY3e3RJLLZC8mRuexd8scA2EYF1ytKAbzmSGhbk7fPU
y73kSj1oiJgbhEyZ2mkQBVLQKdy2C6IiRAHACynTPSglrWc97H0VYWFcp8659ZzDP8/39QCo02wK
Ge+aChc4qu5sB2zgojQCR7AD6rHO6W20ZM/VM3fWfcDnfHL+YJMAa7XCrv6XnPUtwVLtV2XEbxGm
ualmMITlr3lihb6og1gJ2gnJIxZKGXxdeYLVIng2zUOC4/H2zN9RX2UF7jteu6aDI1MK3SWov22R
zLCbemo3RVk7cusvQvOnn78xmqOZjXOZ4Ap6sCAFhtxgucz2F9VRhkKQR4Tb0Vx0Sv4oVf9buLmy
CdlSo3H7YRMOcce8mSLKOseSK8g4gvCp4oTijBZxxhe9Ley96nTKS9S3SqvqkqjhVsN878Bb60H3
Senz3WHogaet7f2ANww+SRSQd1JRPPZM0Ev27pCpwzUl9zsK4abCrvjk0v4PByV6a3BPXMjEyBnQ
nh6KnygGMo7jPKoPmNpZRu96Fbixd6EXBS2lJ2qZWJTDTlVm8kAgZDZrUoBvEdAEeqvVyvjwOyrm
aSk8OyntHpZf8LCzSm983gG606jlB+bmx2Qv4305VtWKJL7VmTYAt3XDCccCf1jHIpE2AnAGA4Z5
9Y/f8lr/PU1r6Jew4o3uR1xFXhBE1JD4IR/RcqZpnW303G8pf9haZAgsxldDircjg2+ZT5PGUEAc
dhXLixVQp7lpSyN0Wu3kHO1AXeFpxteZnPfx80ArVsWsey4KD9bQ0Xlh+E2JoHuPqXZ7lB6g3ZY+
9hFpsb6tTOgBazcWAMVoAgYC3mrM7iBUeb4UBKCv5WRmXOhYsgngbrgD5L0NudMfG1aCoeqCUoDe
NPGCc3TZyI86Rxlt/3JPiuxsdmZh/siyNSCI6Cff73GGMsec97NDYxKN5WW3Ye3ZlMUp3j06NTui
j+kvlDNLOzuF4l+Fy8mRc12aa8InsYMgbaXWUubik+ypTAJ9q5OT2FClvh+o4PvVKmmL6zLrFBSv
MbvenKXJkJU13ua1c5RqgXMxbcKo6iNJgeVEgnJXeTWET3o5kwlM3l1PZkH4BG1pBQH7v09eoiCx
KxCM2OKpXqKfPylnJJwfF1ZzRDq8FjxnlFxfyavE9xTXq5jaTZpMgKt/YRX5wznkKvHInVS0I2ku
57d1zITBbHHDIn7xt81pow9FRdaO8vrwW8JFudysXiFlijtxE/erx/P9GLLM3u3DB/YfjrL4Cmps
LpsvbVDJi12NHAzYB81SH452lAuE0U7woq4kmRU5SEJmLZ9FyuPFo4Aig0aG7dY9z7NLNRDP2PEn
3JKFWnBpnGTvC9C2+aRzBHVf9hThwVEyOoTn4YK+fQETr7znjoHL5RTJGlx12vSmm6BQTSwOlF3k
cmDfxLP9unExNJOJKHRRsKUGeBY80WqUkcf9dLgg5/cvlkDscczxPiwpX3c9SPMkcvme80PZXHhT
10eHbWQ4ob81XnNXzjnWR7Th6TmAMkK7hzYPVY5SF3PipPUo2O/9JnlUUl5k+th1Nuv2exA/hAFl
pVt2pWmTuK3IX5tNtMpt2KjoXkBP+2UN0idSOjI6b8CMRqeevKB1KMLQ7+btQBN20BdFtGBd1M3E
IL8OwHK0sfJfzKCGRpa3S2v6q17H6j56x5+Q1FMaiYYfdSL61C+9/4zh/krRCghNz5ewZnkIy2EM
Tu2uerVvcBL10HVfcIU6ufe/EfJ1xf+QG/mC/lUOGsBIek2Ek2c0Y81swAYDTPrQeVxf1rIUrdht
sxKD/Az7BKw2SM6Ce8uSOcIfVJrW4tMnBI7MWmysDHKocE5choL53eI01fgpqExp0yW/1zo1+o8T
v7AomDrPGLgUwZw++n4Njr4yY7mnvevBdDh7u6qVa+vmMrLcrY4yoe8InPJc2Oxyt+A9uzUhZU/6
SjPQ1vfxNzmQls91pbGzLV7wx+4ZyMdKdNGe79CQgOYqLVQQl9pZzrI+mLPxF+68WYDSESmN42Ze
6mh+GUVtJ4EL5M/6ve9LBsLsYiSljDXcbeqxu/jA3rJGnzu0hCSmMlu3TMoMnMnWqu7OvU99xVdB
PMY4SVpUxgSjcnOyPe5vQCEGREylM23l8rKCuZkfp3cODEjhx1w02wHM2GQ0njmOL8MpjsEJugIw
w7S1EJZ2ozUUB0WovZdiqxWCFhxXRcmVRb0JzA8GG8Ui5w3bAkmDVGmC9RaicAujBnrL/mBZPPmR
J7TSwZamvyQ0thRdb5UEYNezEnFQJBdOkxEt3Zgy8gmbUVA/hGfIntF+yb3qcK8reTtZ5OJc7mvC
2M2TdE5+PVhpossFPYcz1RNuxTcj9U4aQT2V0zg4jxHjKNGW3XcD+NSiF1xRXUA99fr88G3AJI7i
d/fDwMMc8JueT0lN/rbuV/DIUdkycPOOLUdzY3yXQDI9gwnxcLr5C/AOBXcuQw8wtBKz7eeicjYW
8Hvyp2xMTTVnLRKJZoc8Rb5zPP66/w5Ciw5Uepwq32u1Pb6oqeEuE8Htr3lCyWUhQ7baSlm3BDpM
qmxNbCLr7QCm6YfnNIgAqbs6efetFVIynEirSSjWjpX9bahOLmw/dhbz8tY1tBlAAolLFjQ3CMNa
rQIm44i1GIEuBaeqrqpjmebmg5tGHbHZ/kCpfhmyDztpau676F7zaqsvaJWW7IEvRhF6BN6ciM14
MTRgAepPR04pj7fiym6U1V+zlrsIJiOUmQWU/aDtO+re6L32gFoQYxDmWfh1xTI78JTs1m4zQi+2
GsPDmophmW1DbKYjQovQ9M0/oqkxDaXbWjj0UMeWPqO8Y9VRLI9CZxGxQZDug8YFGtm0yXL9m7pW
9fU6XKem4EudP/nOt9ahN4U2X5lTxCjpJU2qkP3P2PxV8aQkfywunjJWiKs6zsGXoV1fTKcf/Mxb
JtX2SeMq3nQVpYRjxtROgaGMwK6A3XXZmKZtWUKsLhFyrzp74dzq26xMFRD2X7FP4A+xFht3Ueyh
baxNM9Ec403rNDHqT4RVKdHCOJqabkGMcug/6p1dtvujwhdH4rwgmJ7ECaLGGH4tDyD0BHZphElm
5XAhh7/PW0H8lYrgr9QDj7Zn8zXa5fd5r0J963j5+nhKGCc9dnORh+SxCr+xIWJKdE1DdYW6PnJJ
SQT4xiLpaVpJm5M/q4c+MH5bZl9PL0XQdkZ9iGO/KB3GOZLDwqx8qa6XKZIeQh9MxdHYnOL/mNW/
hFCJO0Vf4e5qwyqEEYXzUGufmeFiwtnX6GTbZJqC+HgU8rQKXkjkShR9CbJqHaCa7A2CgQVjntEj
6iFLqKbz4QwejkgqjAR2eyWhh5z86fC1JY43FcG3huUP4Y0X7xYGd9sJGr/+uDcDs7GIufBx2dtk
TxAqaPU2h6CKkQ4TI1mtDceIklvueBNhJfZb0LNIn4Manqu7bqUw6G8hx2VqS7b/tjjJyodxi9T2
JAXtxQy6NrJtgrcSJymMkY+reFuNpA7/IX3e9l9lldWwJ8sd2iJEL/f+NMcMUKNneOvdXCGXB45Z
HQe/TZ7v/bfa4IxHK7UJxF6FuPOYRT4eFW7km0Te4nP6cDIbfTsq0wtH/LM8Cps2kDJ+voKBSord
YDqe9ryOyjbXcI1imQR92LoHtCTAT9crGVfbOx90WXWaBPFWJyTKR6vqhleD2o11eOhVYGye1jkj
jVK97HV+F/oxyYoUkr3QvcYFTyZK2PrWlH0bjCNumhHbRKsHYpDmeN+tNJFdEcAa1ZtXsFp+qP4S
zz8G6qNxkvjqq3sNn27KhhQ0md+a6LPQsPPGyQoSeYes1qs+17TC8C1+o8vl11nhKTcHNm79hz67
49TszTA8bwTys/qa156hzT2W6qIIX4ZhissykR3psuXTqFu6WmXoR/6U56r6v+q9R50E7QoJj6FW
z4cdV04dSCqtSApXyFx1m3TbfYoYaNwx8i0xYZCvsDC0lAJY2488SfelSecUomX4nCdS+hw4IwZr
e2WCCrwqZOxqdSSUtUvfMt26LE79n0w1qIH4MRu4aGGgmHECfssOyqi2R/twDgp0ZpzmAIB607Kf
KDhBskslL6DnGE9AIH2JkHh/UtTPlm3LmJgZGDCBccpZmWiZiOswxXhUKWjcFSwGsH49WTl8Ub1P
HZuH4zX675kYVi1KCsG/zDcQaAW5XvRHoMpmeihXqC80d8UJ/Jo0MzXsWhZYTvzhCgRKv1gGIQxt
4NstQ4iWbu8VeEa284D+oCmAnO5xD8kShEZG5W+JEO7P1UQnt/PljatTfzxYgtd8WoRVAI5gAPe4
aGemoDQYfGhVPNFaCcMXWQ1omzFWF22syE6lQsA09G6WRbCXgjQauMWiGG4+4FXIP8n9L4Z8yBqL
buEXeorrWdwEc1TmHtIZzTnAI9STrWVAUeTq029gDeJujFqnLvGN6RQZWfeD1t2SutWbsSvrQkgI
e+WMKFkON/2pSulbFkWy+v/5jo+/buRArzi6QSSdItG4wZ2sxnyOTnG/SkdWvHftgb5e1hrhFd+R
rTZnXp1OpUu84ll02GW5CzOEKAScGtOiG6uBPZIQn1f943RjWdztwvTgFiQku5XiFIj8xtm9PAE/
MqaGOAp+M1yDGTPvTNJ9nSBB5kIwG/5923cdUwdH1bS87gfLYx9sQ007r4GY9HYhIhrIuZVMlxLf
9wiDzfeu7n6fj3C9opKTCP+UVuVRg3r8Oj0O0mQiy3Bm+59jpq24DvdZvMyhqpSyQCJZUf6HlWeP
xjFPnxub2829fBcA1WHzz/tR0NilU25qwAQaMk260nRF3tUeyNbJf+9l22sYn+z4pE4QnHeZgw2j
WQBX3XRQZvMKoU6+iDT7zF8e/uelaGsO5ywwjSX9GM/9/pc+vsEtC4x4/E7S26mf18ba8yZmA/2G
docGRRwNb0O1owJb4aSHPOI+eXY7JQNAg+rJ0zYGayeZGm10t1M/gV735yqQj4SNptgb47gEdGhk
4RusqjimrwUl/GAzAweMzwTyZ+syUUPrDL4qP4W/njFFblPvfP7RUo/XtUJNZQkm2l/wFSWpeBDg
e7C35ngMUWTUrjYlebMoIHYa4WloYgU0vg4bX96tJAUJAvAEl1xtaDnr+W+QJ7znFW2Uwswcn8tI
IGDCkYMgDAjTGbFQmyFkwZLOh0jUuQrtK4h4+ssVjFhsAlE7f8ficF6MnSfP7dH0ojUXmeZKkDgB
/i2zMyHOEChuoJvKcr7a7r+A90OOQRSO2gx2GtaxrpSv4nw7PCTXcvftqfKlVgMlE29Ei5IW0Ccp
v644pURVD5VZcXJ2KfaRXfG0sqDSBNvv0oFzgPERW+VeLQG835WplkDwZ1ldto2eQWDrttgPjWYC
V7DLGaKZf9DBkSBTZJ9kN1lISfYmJrIvRpWpvIYLqKGggMjrvz53/JjvTud1ISnqMwbWDTR4GX9T
KDwTDGtRujHdOGGt76DIgms+km9isjEBRDwJL9bPgTlGqhx0Pg2wnhDlVc4+Nm1J/trDef+a66Qm
LLOzwVXE0FaYfEJL5jMk71cdIWk8Cmta/WVYQR7hr5RrcH9dB6DTlIYuOEsIoZXtLNBo6UkTc27A
NhQDI4Bbe+90nN3+ec0xRsoOb81xKVADsh+pVysuu55Qkssoskqet9m5D2c9bOsEIWVKBDIvY72n
VgDjVQIOlaF2LEeaOiSWSeSSG5KKsyB91uAFpcJiQq5gbDTpdzFTh91yiWazPvzyHhpHiHNYlYxy
3vtyitWXwGPxs7H9uhKQoNGPgwrxfBbpSGApPIvIVxuBPNo7yLWKf0Nz5gRSHZ+0TE4EYdw/zmOr
ME3zc6MU0+yFGg0pFkfTxx+JBP9tYCen4FLXSjm5kbsjXCL+zFqfgKBOgDt/ixx+kGRXb9xGNUY6
Imn2OkXlDIZWh+vjXhoi6sl/C63XBVNerEZXPCxrsm8fGDwxldszeWgjKGraBdunc0cVSKTXtv/7
u3dI8lxgdbjFdYxJUXji5aLB+1UIGLo09XoZUWLW/zio9JuruH5pSrjouwHnQaE+P0mEFSvWRRyN
eYR3CwA9+8F2ZZE+CYG5eDhkXgWqVaQWrYlhJvzZ7+ZduXOrRCstXKytj9g77NR6rlS+CIvdqINQ
Zs3OTAsZHmiJfelrHws1KTA2aUfZTRjxHS61RXi3a87ftOTq3QoC4EFeCJ4iqso76Zmp12I5j6BA
iKfrw5o96We34hevvCA9PppgCSPfW0fzjWaTeqBb3kuHTFs70hGeEMz5wwOzP5OXQxOcafIPRZBL
Dy38srRvBBXRYYSyDkdlUS6NdwBznVx0dQ0rGZra3kOEmsbzFNDFC+FuemvE6g2jEqemy9kJ/LsW
ORBb+lKSmxXyqxDNwbWSLaceGRKTzwIDk+qqlTAwN7dQswbj2lAYs8GhN6Tc7VBVwGYc5Fjzw5TG
bwgyTq6fGUR+U2GqkMXlwj/H1jlCgd8mScp0YjmqW62nSZ1DBZhJJqv7lnGiJfPsXoEanLA1BGbz
DFNwpUf9f6263rBF+eoL67p7FHTQ/mkF83bVtHhqmat7CUepcIA8UPPr19VtaV6yqI6CMYi5oMJm
Q3/OUcCyCAwn8/I49IvTXrdUhLbX6+lR79JNYRnTvDEHZFhwB1nedabUx3xECmINP8yiNO//B+7N
PZjOGW8A7smGoVy13J9AGZlrus7JsQ0YD0DbJYEdc46AHeh77LVpm33YRazd38PWllP0e76eaYjI
zMaipqmecFuAyKUyCvL61Qg8wbqTNg+WTpnKbAncHOqGpsuhEXlJz94aYSZckdTC4L0fZ6fsQdi6
GuHkKHjP7V38FIVVFWcHekGmGhGaDEmPTvuwz60bpAuV3NiQ2Aitnebpzf/yqFpqXt0cmQwEKWad
Ua8FLmY7/GGzigsJZkvyPyW6bSuWUa89s1SppOR6csTsC5mrEGLDy+K4IUlraRsU5NJ9B2F+vNRY
2k7BoBasQrOK1z3+Ij/EQEUaTS21j2h5r6njy0BFcCC83YY8lPmZovh7d01Nv+EvclhXydy+Rz1v
zVsvpRslgdqmBsPZWvzLPDjco6/8cELcrAWMcH+6njEwcCq6fzsAlyQmbxfw9efDDiTMPPSWeNOu
KoVv7baM8M+8kgPR3izfdirwmxsWMxOGQCeWNkP2KlXrdstotTJ0gQ6WCShxgvgIwNqwOuIadoPe
p/JxTY+dAy9cl5x5ZNUX0by/zM39IBpskaKgPvflXT8pCF2qrrcbB9TPQOuc+nEFAlKUcYuAXL9A
B7KPO7UwxbZjl9YEIjGt6MraNFpJYHv7eKUxBTc7wuqjjoLC2V60QjLS08Z2ZhUxK83TRrc7DgOY
kfBbO01BLOCJoZOCsKiUXpn/LloxDKi29gnQfu/aTZOldgH7UKFLOr0Xc2ZlFKdXibvfYS8jYRxV
5A5sT2YWxS0BnidFE7WbUEbccLTgtvDM6HhZvD89PJ34uhNRB2RXO5J1FUG91aKaorDV8dkJy7G+
Y9dxMM5FsW/7+3v86A6qklIcIaZ920lEjHlqZ1Ht1yRYjosZfMzMdhYGnlUxZo/0jRbvGc0OFfjH
uSvfl10fMPfasr2rocwmf8wXoL8jqdzM+xLBvwuAmxFEmgnzMnSdjc/ere/at35/0xzzqaankGdQ
X38uwztNcd7xTTDktCwv3ociyxJF6/EFJ6rR9d1lTB1/fr967LLKq/zU710Gd6zcKNxrYdbbB8hT
kTT0gaPdVU4Nb9vzsvke0fLq36DiSX3BngxWmrCV5nfzQnFZ28qhCUPv6Ggtwm8vita7Vpyqa7N6
zAom982L/WVUtLQPWpAgzmrNcSj43f+kqp/lBsAO+4wNqubMlKm325PRCK2ey1uYPaIPP0e03GYv
7SMcOWK4DJ/yMzemKH9hzeAKasi/8botSft4FxP5Kltw8kPvaFQPyAQynC6PnKNqJZC9rViDez8H
MR+ZpIGctdBBUtqTgLuolxTDgR6DBv3wg7RyT03TVqQGczD2gK6JBtGCA9g57Wq/ZKw3YCub6q/K
XgAVhiQKmuuJ7OiSFHDflpcgY3VoRxdKuw4SAmClpitJJAOJPNF13vvUIjHYO10EffwWMGvzRcHy
0Q6S6nYX9BPTYyS4jfasSYbL8TPiL9/S2KWHv/tf47hBq/rGwWYtcfHKcQ8j1ZGUniXmyAFAfoTD
K+a5zkJDznNJjtAOy4IQmzY1x5gEW0OcvaWfpKYY48rRm+6AnIXkEet0JRfDoQJCLACJFA3w1jkS
a6a1t8bC6uuPIVc14a2/X2mpZcFW9ED+cG809m9VhFU/ymL5GcCSHHSc1rAvCyB0TBDRyxKfBo0S
bKYzyBjsY9MEN7gn3dUTMaZf3VdLVnweUONIu7Yl9yTRurZl/kjcQmMjioYzXX3uYb79Oaz91u65
0zOI/88nQ0BrJD43PqQmIu9I2qwkPdiALk+yqZliXiYj/Ewa92n3kOZAtlhztRHYsXncm6LqyzRh
itAz4yz3HH9TIIPTH+1u/C4q9wxVAQZGr8G0g7BP2A+AcRU7Dkr6QiW8UYAUFVSmpS5u5FpSN8Nt
5NXTQuZWddrHmfQPkCOenxuluu7y4B9j69Ik49Ai+ZzuC7y4iFSw5glRhA6HqhnOzJqfUOumplhm
/41HrSlB+ZU23R5AIWX2TwjKs075wtM/mE5YsvYL3qfxTXx8t1MYGNp6KUD9/mA5YAXvADXiERyj
REkw1abtyhjJ7waC5RwSm5EwSRhI3+Fk1p5wtSm5T2k5tYIz7vfadd4FghvIAOWKE7WsJBWV2GAG
3sJspc3g5ne89QrwnQuoy62k7cOSE+NygSqJ9ubosYp0+CFPqKr0qSPFBn0FV+JEZcZFwFPWLQKJ
FodPhP/W84rbBy3mv2FIOrWsBr8XVR4+o87w4n7MADhYEC2uoHVREo/u0aSqEoW8UlvjMSffOm07
HUTNr2KeKhTyK/2LA8ZdA8uwx+7nKii3uWpVbI1zablCoj5gn4RBtJp0lFVKl9CDbBgPLm7AEWxi
VKuOVrgUJcHnUvWCA8ivWZl3rAMkBcbhXN5jPEQCo1Rio46HbCW3zfZO4bg36gDaxBLc0POKRXlL
rbXfAfg4P272ss2bfTZj107IyFUnx23A2fV9lKu+k99NQEryJ/3lUjgUWhwdJmDVsnaSMjWS4Xi+
rSpjSZmI8R6AQ5VVvut7WC7qm1pW7MHgEZ7sV+SANAozQI4pXOgPyRPaL2hHyv/myNtmR+W7Sdjj
N4SI5iZPixu9wxWnYoWf0FbxKHp9I/a8oMYbyw5Ta1sCZBXKk/djeUj7XSUiE6uQ02JLiM/finI2
lJNz1G3X7ppMtdQbKrwJb+dxbkxGx8aF1XKc303nPBp+sXxhJsN3kYHHQ+3P5gXZc+25r5myYmBH
Xqh1jNwpw4lHhHXKq0hFKs+iB9LgbsCaWY4SzvD6SFHupe8M2UIv8LaNOnLjWdcZFl6B6u+eblFZ
lXrI+zhbRMmn4LAkuYCDTFrjE2mBE/NHjKpvmV2h+ZPoDLr2RMS10ral3LLKBCm3s6imdxFckNwj
Kk/8fYkv1kxYBX3tUaQOH0WAvs38UyZYv9no3i/aeTBpc6SQ7bdcz93RLTNevxgNS+lhL/EqjV2x
cWckLgOfCiSd4CUzJDLt4ioZwzYUr8fuo3OhGY8oZk5qHPz2P9Sr8z9p2+n/JOl5n0RGPQlK1Ojp
Q2rCjxccwwuyHBlg6UxxP9gcUaj+bO0v/C5RRZkTu6j+efgOZz5GgKsIiFS1QCxHdJbfC7T8H3O2
WH95BOl/hP4e81av610A6tSIqU6VBd5f4EPxhZpqPOh+Ls4/1J7R/BkhWhb/mFMHBXAeDWEDMCr6
SDMViwdzMvL6hHIsnuOoNgGXQGm5II+ymBgTL15WV66zrqd68xZCY6M1ATuiGLlFQZu+NQtTT4WC
3IBRP5Fpq7jtWDapFF3B5gb4cbEtuWNTEGOKeipv9qgdvAzEF5G8x4ZKQPhQTSBH8JznNssoSTfx
ICsdtAd88+PHci2HTD5nM4/D2s9HtY9OUlhrsGFjb96tVm6VoLmtyqUNvsvdV2kODjSa7A0Vd3Lv
b88EiZJ/8RTbATyuUAfCnCL+gibajOcz34uuPl2nwKWl0SqROMEscxweR8lmzTigd2B1ToeS924v
mirEgbDlJzZbUdqwt4wcuk4jzoXXmM6S4VELviUmyM0XwLGNRIf5Gq4Im8VESEyrE8EC5CWrxY0u
U+/FztelOBWG2WHq/VxGqIFu4b3wDNwP31O0nZhWbZwzXqAvG2KHeT2hXOltvDZD31LJtT5ccHDl
H9TeDTiq2uiO8u1WTTKW5vWzjmAn8P87viSaLX5zA3ndwhuB2SMDsVzDyZXR8QQjmuI3ijvIqakk
zrc4jX1OiYwLWJ4z+ljuaursFD41+UkZ1R50kHeo+ehYgdfI/HM8k3ZPi1bb38sh72REgEsigTMa
epIwnbAZh24FJwZIT0r61KSGDF6PGhc5NfKJJGjtGEcKMbFS5x6STQ/F235nWOfdqvf7dMEjETp1
/uQMmm+Vvs57+9DXP0glFvsHyErEUfqXCO//hAGhDw9xO2WeJOflVK5Ruql5p44SSS6a/dk2TLVI
4lQ1HrDykZKvqPGEnjsuWuE4YTX3q6ELwoqSjH7ylMxR2ILYwgqtO+ajgq9ht5Gyx83QNGO6iV7p
be04hmoHDppzEzuDaYLBWn53chG04WDgFddHYCvAv4DSSAcvoRTDpwaBwURVnAGX7vRX+qEJjIsJ
dJ9F4JiWtBUJ9T7sq7Ne5HbFjwhc7BPiYpGF5+NNda0Ru8qZIQJPmRHz972jrjyhNphOTptRfoaa
5FRZfRhK5+7xITbsiijU7iuYURgCc0yZqx4hd+F2SLcr9coNwaSQnrhY6ZG/Bm33HGiJ/KuFGXeS
ww8ZSmRudZUXoVyJs6WOYU/XV0FB1/8QiD9hjtIFZtI5RM1uXZlrqhX3zzhBiKS5TCjpWQGsGObT
kJgoG/mm742pyGUaXDRh/KZ5DewUHdva6ahdOGscGyFuDkrcHm1uA8WyxlNpnCatP/CAhHigzQ/u
BWCcBAhYzE9E/qQTIK66JNQPv+0nHNhiFmKBLmf6BXDKYzQVNT3G5yvojzDSyFp2ZysIBUpdGMQQ
9sj6topXuvK4zvArmhmqqjok8wA6hF0J3SlKNYAPaoPcQlVbNUzoYuDpiSuJpEntymQGsWA//kH4
vN7YVGrrtulYI5jFH+nev1j3loW73sBFH01GQMaARq30VRgeOG89b4rPTIDywWwBry4uVU/F7VJp
f420mVo37g7RwqIfuqvuhdA7fZwd4FR9j+H61RG20yMvFMia0JWnUGC9LM8uMbdixEbehVqxlcLD
fGDjbnW9b6yp69kOsfT0Lu7heYys472VJQMwFHmb/DRWOuf4gvrXaR5xemiOZ6vWirtov8WHO8dS
+0NNAGLqwQikouVJw5UCNrqj4ghjbiRve03ILToS7a9UjUDi89f+as9yakp8FE1/X2J5jq/mWlqh
Ua21JrP6CX5XbcuEC1SbBY6GY0I17NklVvRdU8EO2BQR2PoooSCQY1XJ6jVx7QO8xg1S6f/+f38A
CfezjhN+oqhR9uRrojolNy8OguXOaBi1BfbeU7Yqf4vIO4Ip49yOhr4dmmnSeGJiDSzbqBVtQE+Y
W/jUu4e3BA8JHzNYkG2cYU4kH+V9q6mTDRv8UmbrHc/8n/ow7GMHnDZgxAkNeIW0wCLQ5bmxAUFh
MuwziNI9OY9AKWF9E4kDZ/VurnQma30kX1cLZQQLDvVODlQPcBgDAXNBr+4aC9BiE7kBftMi2f7p
3g9GVdSUIzwTAza8pmA/F8aD8eMLr0OdYXLFWkO40Uk+HFRxmiEbMbW9jIuUQ3Ih9FYi58UP+wTG
OBm0RIehvxVHHEE4JmKlbgr3o3JbrsGe2Womp767wlv6MhsIvglkgJ5Fb9CYmPZTsfvFIWipfezR
FGoSfCrdkMBRJm+FJLt8QUyFrIu5bO5FAGxxze2f3gNdTaOWhsldDZSwINmAaFLO1ehbBnVrytgh
gAeLD1Z1L5eoPIWpcUxt8cYsakRcFqPcNLwoiWOmawYj3lnHAZwHrI5LG3kRj+gBl2vrMcDewNUA
YQNrgviUkSjcDTww4v80slNeKyBx1u0Zod6IKaZheRfDuxvktKhzniRmCLUXCOuKbRrMt1wkWkQa
XkqMzhzxGysHVJt0YWau3m7Nj6JqC5x1vExhXZ9NJ503dI64W3GWDY7axKMNS4SpukvfisYmLx9R
Z8lFQ3+zVHrdE8U3Iweop5GeDA+UjW/dqTPp//t6sE/dEfypce6nAsstNs/EKq/kcafhkaNTL06o
nqxg555LMw9Jzgb2VvEEDnyc+WwxMtmLx5awYX4FnpB2QF9KH9HhCCI1x5GaL0a5u+XsvqsOihAa
BjQwDZfCQrbZDtrB8IfTxQGIYvSYbcX8CCWL+UVGRLYlypQeB3ZSFxdMUUiFIC1xFliV6L3bkAaT
Bd+kaxasjotGxHzjWEqhIH2AwTi+PA0AXpGgZnfidRYZ3Sl7kkip8QLqEh8OgBK0ZAvV3mQMFJA+
7LXSuGQEwGnHzGIjvjyljXsGHOx6zUYc+0rEnMbqHPH9LykobnG1XjqCliB6YchkyoKl28aIDrUP
rRdeEY2G/qd99tlHexfhM9ZphVUJQ3V95hapzWDu7BepFlHW9TfY69uE37GJv7f2d/2/SNUA8aYC
ssPSuNLEuPvdYW9hY6IIe5iV3vEIdyHZZoOKqZx91ScCuOkff+G7XCo6eNNUY0CsVcoQ2UvGCMGa
QLsed3+X2DPS6rW9CqFFpScmRvtR2nXeA14+um2cPmDFkvdr4RXZU5mA+HJyHnpVSzcPLhwEFw1C
R3HVJVnJapBmhOrxwzEe397jkTKeUEA4mzXwUeS8TyroM2i8MpC60ipW8evpqdW5C5IH9Rcm68Un
mBcd15bOmHAKOcBZN7hti0UW8vZhVPZXCdOlEE5RSqVD3zHc3FXNU4Gb/oKmt/8vSX3NkNzwzHj+
SUEYMJ0blA7Az2q3icvfKV9Xo5yFtQqwwwc7nXV6F+PYVM4y0Bdm3bx8PlDiESjzOXtx66//4/3D
Zsq/JW5EUlZnJy9stIfgL0LE6MHJiy4gJMyWrnquqtoS510ryU0u+fQYue6PhDFhe+K8Nr9yxzxH
Xbg2g4kcnMzRr2mtMXnWq3EuCJwtIfbyU+3poTkEg3HtBwxmkU5cFV41VCwn2lwp9eQT3nD7WYM4
YE5jPIdI6ianqvD+2cvWLb+dKXXg7XtU93bQZUf5ynootvPdKCKPrtcPnsdn2qxtL8duWJki6rlk
3e1uvlLYouEz2s+7jbvljzq5JXKn6fJLXyCm3YSVRG8m+JfQFoVyYDTPseHCHp7M660aNKb4M6Nr
p0kXp/yVLWIOCo7vD5WTyOrz3egdMhBF67HMtmtFd2ApeW3zNgdRMYHsUc0ReuzFcBfPbHW4LzWz
OkHCKBUmCZd2d/pW6nq88uq55qPE7D7YtTA3YvsfaMYBiAJTzOAGAldzJj9vIsA0rWz5D0YO/+R7
/kIdGtpF4zKBH1nZ1poTZOcRHi51VLaMAWPC9tvetZxHBibQbyMFfzjwMF6nDojbq64SItOW3aIj
VSh4CVpp/W/txoMlGV4rTZG/CxYWTQRD+LXmauIdYG5OwWuVNlZygkhC5jOxVg14V5oBuqW/m/iC
8vadaKbO/VscHztv4Rf4kLLcmAB+2oG/5bNGJSxEvI3EmIFJvGsnU8D4Q1kXBshwX6AwxSjXYl0M
0nTrPGdlXeOlE7PhUHu0wI2fYDrRkYzg3m94/UUi29iVo7C4WsLstiv6E53YumaaR035Mph6f8ab
Fw2cGDntbwE01E0DlAyF3nnyiUUer02F89ZUFk6BO7o0UTk4MOKZzH1rkShzmcDiWdDq0PJJlCNr
YhbTPpLhMNAKd+vIJ0URhUZ6JpBatrLgv9kcylYlySr/uAmuKpnMh2dh92K18+gVWiZjZN5gxBa/
Lr3TLXIetO8ta7N56lgfbkdFcjYftFoKjYwNfDUIXTzCIVk8hMmKPIo9SFAawfbk2T8BwIfaSq49
W9G1ddmL9W0OXcBsK1ry7UT67dbZI9D2pwarpDzyr1nJeZhPLyAMEJumhtrlFlI05MnfPvZ2T7Z7
WQf74W01vlh23syrO7VmKgVCSd1bOeuQ3XOgv1I2UmYK1avGCBe+LrhKj5h0ujr3J4cL4ar2YNiv
i3ycUo305OQ+AfFyz8NgnN6jgMU4j+qelvH4y9qAn6av3FVc5rDonYOQO5f9TzEmO2Du1m+CS4AX
fQxwRMrERfQQTBZFcINrmrAb2gychQIraC79LBcZ4U2l4M05R4/aesKVrYTU51CGaE4FgxQsvk/U
m+hQnJH9f8bx+TpHmTbmT1hVryLJULTGKr8PwYSbCqNnewElNB7qB9cDr9bYaAdwP53Ln7yqWZz8
uSD3jlxnJHVljTUv/Wi6hIzk9BD2TlVjdKNn86ty/XmdpS+lZO3/zBmdnY/FIc2j7JbvGACC+UIZ
ZgYtySXGrRE7iOpSmQW/8bznDTjJ+aOmvk79/DdEPnGptqwfwCnIlzC9YF7yy+3S1Vsi7IjkSWlK
RIkYwbEJGNkZQnlA0hNoblDxZUm+94WuXZURCX7sowDv7QYsAjsTNQesiFXh+Md/dJrbc1ul23OT
cAkcYISmi7mRJr4SlRNa5gNKwHQP+xWgSieBK/wD1wVOMD7p1AiiQAO7MyLlHIyHlyMEdqHfGNTi
xoXoEwGE/qi61eYFXqB4cy/umthP6CxRCXev0XMMG//v4jb/zXHqDbEp4RqQ/YCZBroBzLBq08YT
lAYxP5ltgUSW04V42qLdPEeF0tj5PJTf6u+Yj8ypo1jXpgoO45fDl7A2eVRXd1uoOtyTxL2DKIig
2xfd9A5/rey5S0lukRPqjqjZlRK7uJ0KYVfGSwosyrQta7BI48tjKE9HEifjtdWOeN0FkQT8bBjH
gdR49D7eZJXzVBga360pKV8096SpwdPF0tCbz8VZG2efV192oZKcVLl6JV1HlXzCJ0c0QJ2JUU9F
h7GzsXOPCWrbNiywfNdfHsGfTpbgo9dFDYmEbrOQbtYjC1hhkQ9ATZu/BKU0ai5XJuJ5R4YELp5z
8XcRtH5BfgO9nq381xwbeE5Cvs9G5ruJy75AmxHdoHOxKKFE97/1O3NzDiRq6NOnvOKscBVtBa6J
G+qSPGi/AfGTVkJKd2jNHsteU1HTEhviltefm3Jd92xaJfKMjXMMEikR0JkmN0Pl0JMyt9xHjg43
gttDsUtQAYla/FjQw1gRL2RPB0+SUFOrpqoiElZ6WZ4imuLoxwls5loeAJInm7Vt9zYVl9aGF5GV
Hu4wDFA1BHucdAA+d5c0wNJ+YTEy3+lR29EmKty0Io69wJWxy79n1sTDv7f7fC19UcWxHoZE02GI
5og54ATSdBUOHSIrSlOZ+fTSXOxQYMW/SZkf0yjqExdMxgawbyAEmfYcMZgjaTkgi/3kF2KVA/0p
f2sdDai9D55qZa4BUulpqgGm+MoynWov7IKQ5ulikSb3PHfh0D4lPx5W2MYbRuu5ekMZQ4QFk2OA
MdCbdGse9IWQ4h2MspCdbJesVUR0BoVY8+RoI8yyOORtThivYXwKDZPnM2rjeIk1mTqk6MEx6gVE
ld74T0XWKlaxbkPTdX1CauNF31Rk52yukkR7iOii6ZnkeXp8LfdGIPcLTLdRjyyPdpSzQ1VZtn1p
VphSSroNp9mD/X+DAXkd7OqhEBRcFFKDgb2UQ5pMrJT+uRdkMPkNKtslOCZCHVtmuVpWnG0LEcHj
nkZR8MDMwzAwUP0+DO28FGShnUv4oH7lZJ8jgKwmSRiykGNx8t0n4vdehLwWzVZF0WCSxBtrTUAx
usjT7yLA8ccuWV9zFhBKwDHhASZYxI5PwlsYi6LIVoT43U4Q7iJ/D3rCTvu0FjunUJ6jerx/t5KY
Yv/yZy+xclBvEPhoIKfGSceDM1mBgAuEo6vtmVY/FLtaYidt2e0Q4krcwVpyXKI6SBWJ5RbHjBV0
byUpSxmGOFSlM4Jt8nl7uFFnb+WFFvzYwZUfIlfCxVbUUNtidBhcx/S/Kw8bTzaL9XiBJCIZyqLQ
s4UxHsFTitbwmRKhfu4kwyIbNWZ+UeCedcwIw6x0PXhEvKjZT9tvDf1YQj0zPfXRHFQgzrYpQjB8
qr5lBqvirCJaOE/WYrWKBFt23a67swCZcy97Yu1OAXCe8wCtGVMnZbROc6jN9ixXlXDw19tTtXj9
lTwYUnuArk8YvLyBlx3FHaKn8VCJHpelalbmK+wELn1kTtTwESaO/gFEd14xEDvV/VFe2ulZIoR3
yuAMtOxCIRTEdunnVQNTxqkmVaaO2FumdHFRHS6/uE69E3lfsQR0fxd3SF1Z9AofFqSi8XnM++jh
A+iz/zGZo3cy9FGSylgJmyigkYNsJdE1oZlaizKSUZa6kmPXr9GFBZEKw8gvOYK5R0ebYlk3VZyk
4AxysU+dx1uy02+M2gkTrp9sCED713iyNEmKnbe413YB1y66YIFMbEmMdEjS/8srj2gIrwkPADo1
ZqgYv+1u60eM6GtJv0YN4cvD5ZBOrDvcFwYWg/ESLEbIRWwbmaW53Umb/1RZyHSoNx7rZ9ejI6aO
C+cnLxIQ1kDO38g1weSpcd68hJ/Q+f7wv3TaSupizvxBH+09NFOCiB6BQQH1JWh/jg2KLq/NS5cw
jYDoScYIdRraEO3Q71vqnQfaEb1jJgBjTF6CO5Nj3IS9OkEkDOf+7o8gsBvbNY+XOHiCJ165gh3K
whLsxUVpjcdMBm9oUvLzDg9CHbN9F9n+Q2jereWs9/hl/ZvGhFCzsHwx7a8bK5jG8Y0QXAIqc0jj
2dbdQVVMJ1q3qqB8Le5B5wThaCPcynjE6Ji2GSmNWrYFTNiHlwuD0AGFxWg+u24xRO7qMDDZrUuM
iKJUrBbnwmS8N9terbIN11QkYVph1ZDQ8Mc2qKAs8rkkrvd5e4QGlGU+6tO7CaD60JxXSD94VfAS
FThk91ZIaR3I1DhsG8C7qLjfVZuvLGhy/WDO3OASqUDkCQzowJBLZ9d/fGGEepGTWF8iYCppn3qg
lBfzWB68osMiykcmAQ0KNqQiQ0F685s0eP9iepn9S8pKCObMxvK8P9HqczfcS4JpAlSLcDXz1vrA
N+5kLPPfPWFTQgE77SPufhz/EMaA8TgMpQCr59gA16tv4F+pOiZ6WkQ2IunY49ySf9FwCRLmpSdL
NqucYH3Y8EWXxXnniIIE0HVpCz50TaoR0xAuPIKvkmCsf6pAKOy5n3861v2dzW24IBa7pb3Qpg/8
mgsZ3DoBlIkRnuQO3XdMmUeb4M3WenS7nxyVeZbMBvxkmrfTT43/Lo/oEPDGsGg1OJhJzXHgdISO
o6kY268FvhxtAP3H7te+dp33oH/yygeM9mUsDewarQXZhB7DPVmFz+pXcsMZggMKQAzWTPtiu/Ee
MzxiBARyXn8mx9v2rccVQbmUqQhfmjCg0bADS+4yNbuxxFQfKV3TJp0jdUSUglRMMYiWUTl7cTXG
fqxFQHCE4jhXRxtfp16ULFx95QPVBiHbLnhA7htYJ4r2gg1vuu41FM9eO2mioBxrMi9G1AJxq090
yYmhse96uGcS+qt7SDFFkjGlDl+phuBAHFwJIIstdhnJvwDZ7UYW/NkcSUpN3y2v2JADt6Xrvt1B
JWLzZuleuyzKkCBRf37ChLglCiDGX/Jkq+4G3CYFaomJ1h3BW8bv5U+QWq/ajDoVgEJ6JdBCP4BV
7xaYJmi5nsMXUUgyjyoWwpRfeuES++vL30TgAd1xiPriVp7jv+GVpX6QUMtH4k6Uf9wsbewfNc1r
r9gBPQ0duLvXbmd1PoS3bbKfRcJhSCxoyu+z3NZWC9rfrXH87IFvGLVpIIZwofou5CU7oa/qYYqe
Upi0ERi0W1drHFdxaSm13TyHV80pyEGveqcnYVEx2xuI49kZdjfkWZdyG//AgbxngJPS4nh5zMQS
Oh0uf8CSrcUDaEDwUBT/UIchI4xzu/EdbwigRjzYSkA2XWKm14fIMN3jMn4GXNabYF2V7sJYmViX
V+Mnl/gwVCdFQqzuPsiDknaBizqlNILb16EIkBk7QS021nU0fT33rDHLmVK0Z/XQE/GzUbjEyMVb
YudWMp7DeusP41natKTomwctTueonDVevo+4caqDZuwf5Se8e1IrwNvqpjOCBmf70MIxNX0pJ2BY
MlQ+FY4t1hpQXSHNg1zsLPIx/6BQcIrVb5yHe7QZJhI9cGixZ3W9sLhc45KSfaVorYuJImxMpWts
0OWmXAG3wsNLunQBj829+eCdbKGcy1UzhZmckd20fwLPbvVn8ZCi0ERUTltByLjdL7JJQm9t0cDR
HzT1gHdJJdaJHI//3fD/djx15FeaT7sLs3Qnf6FE2JR0BoTBjfFafjBmLp3xhekFm/EHKEocQIpv
LWAjL0WaGdsdikzaAbyMIyak2KybFKT4e7AUGjQ2OPFg5kMu46Gd+tbmbtjp2WibUGLBeRnRwuso
UC9RcLhBEB++isGbsamhuOphTMLbAuSGU7ypad/9eYt0lK0+iX024PTrr0QYR4iXuIcxposoVr5R
f/NzzjYxqFG/dr9aDqbZoatZsxWDROBGoAq/VKnMxlOUwUhItMDi7KErd1c1usX1L9VUnnXm82pX
SSDgkPHSKtBlM4OTNqo5ZDKwqxtL7fni5VQM3kbXuxvI5g0NrZYtf/5sMtt0KmpG4N92XAfjsAu/
yDTjiuvi654TydWCFRUWU1djkg8qbQ9Qy98F0b+AxAzyJPnq40yn/14+xHzodtPlxKbLYyEmoLJl
NO40z7zgblTwOAEZWtFkQ+FNL0rIrsL2tIPyPbBP/zza5+HZvUjAvb6Z7cW1ZecNrtlGobSO8wDd
ZhEa97bCMWqnQ2D1yWCimX22oVx9bK/ks0exHnnl6z+NzUV0EIlr482/8Pochv+6m0KO8OIr7PgS
YvNQPBwskTb9gz1hZ9Y6GKQiFEPmffXPSZk7gCHcfWq1QvFC6lCx7BNgv1gCSIDZFTQp41IKnaw/
ZH90YEYABbBXLSAeZeLaPiE1BkEBNlOuphBAu5tnkYCcYSr6e0t1bIeip6Mgae5r1xYZt3tlxmtP
kym0gX+hf1juOf8GqPOg1L+PRSBQ77gRVvGUM7Lm0LP5Ry4DENsG7o7QStT4xY4yYFsK/vnIKSsr
FcWGfdw/LpTRX0wGvr7c3/T91y6FUsndTJrNxG+2D2U+FALcFD9er24nSPJsas3MgFjwOWFgnj24
Ry+bdi4+RMdohUpXYPzLMSSaaaGX3aRj4CL1zLZN4+oi1EiCeEDprUbajgNf1jQm1NaYP1AvvRpJ
R/S7AByOuO7SOdiQ9GnCO1pz61zMCd4Qj3e+J4tgzrnmu7tXAknGLiJSnzUbyaTg7XEMVF8UTZqU
wpEZhLgynkt2qskX1/wAQrOCio4BHIEdfwXz3Fnc/KiSi13BNvg8s4mXC4YFV3KeC/k9QBCDly0q
MlNzxv+ytU2DzKFzq4aaQts8RisQ1ieisBIj6CsCVYfwaXmKf9yX6uMmQLL6C3s7JzZvXWCw6ZNF
GFDjVn9bFpVeVZKPnp04GMFdZliVJgbgdZs3qHVMrKCxIoKk5bDFMcIahDEC6pCNNwU4r1CuhtSl
HzbRQ1523Qdq5zTQC4I1MevoeQaGlbz4vvjYCDu1qMtDua3xQ6ssj396doeUGAv/vbYD4DAxwr/c
FB7tiYeqYRP+8XN2lVOQShmin3GYSMngfwM1FpwcdheOUni5C9on6d9I+9EhzF4x9YrCzorWZQaI
Za4+e1jDDVUEUogLcfFJfWzJWe7BelL7w4t3bOMIJR26MnXEYrHKWS8S8EgI3H8d3kCihMbPJpVi
m2wyHVlnnge3ADEtcrLIbG3L6vnG9pYuG27ois+tgqWVbmBNPGduTBJyGMf+FEuvzy3b9Q4+VrHl
vvU6m1oH8a9FIdk3zYKgmPXLTgE7GWuGdGkKVW+ARtPDF1L4EL5jfIPtBDPE96WIoVVUt81uC23k
MWPHHhtDcM1m0npXn/a7rk50Jh4g7se6J/HhSbdumpoN7cFvzW+j9pT2Vk5AqVvD6pZb6NfOkpUP
A2iZbk34kcH/c6DluM8kvju7b7EInhwnKR+T4ADoe0HjlTlkvHGPm4tjZ3lRSJ4L7tYziBSyxCmA
yuvISWAnFXvbTlbF+8yl5fm0QdgsO40qKNXdLaZnWe/iowYQgJl03VUpLVgcPnT/yYNM1Pxbc9i4
kPOv7dfd3BrL8kmMsVM91k/jw3VN6zujKYDDsfJm8R/LJ9iUbXSwcGybPeph4hh2bVCDTNSiilzt
J1MpXczB9WQWEhJPi+NuMd8Ws+Zk51IyOD1RXO9Nva4R/djuYYZzo1LdlEIN0jUwSNUsj1EWcz4H
WgEp2BJpTbonkqQohFJdB1F2lGRYJBfvNGif3+bZsC+EVHS8nHMNTP83FY5IEkz7kKHq97qN0NFT
E84V/N6raO9ME9vx7Co6RisxeAsutjxxzIkIK3x0q/5LAYFmm4dmrKASQh8tV1eA9+3TQWGieEx6
Hrwky2TGnsXQXrHOMdQbEHezeL+os5vm1IgrV4YKkNuQDfg+9vDNw73ZcOfb40X9XdIhMzNwB+qL
pSzH99/mK0pZfdLm/n0uHlp/V4V3W1Vi/txBwgsuT4UbhslPeVBmteheRK5vBltiIQ7nJbtrZfoN
4h7WcSWjvfkig73rJM5i4mngLhvpFCvYW3+KnZtiVcqgDr0+f7NTm0ZkJMVm81flGE5B1ybndZbo
nfddU/tU49H9pgeNh0RABkn7rdu+DV9g/3x2wBKk1MdzWLaVSjkSQgnsKcRYMk9kHkhO32ESk0ZQ
Qx1BHfOj47LtlRsLX0kI6IjHJlBGol71EcjNUCqs1cw5W+hZLkADIDD8aroAHDFzsjhFBAp9umhE
HYqcDbCs/K07Yy7zexYuiVQ3pm3hprKbhbWllD9R3ct/2RzRARAX9jCAajizAcT7yRQRMr6sA7jl
JK5AbWZOWtKwkii4iLJ67uhwhx/VGw+CId43Z8YsR2YXBkBUSSl/A8Ym9c8eKLtrzGG2xeYlGq8B
YAeSeZIfxY0wQ6JzdZWXYEhmFz3Bsipju4ztpkbjvYAn7A47G+AFhqIixxLOQ2biKJBl3ZzEbf0H
fQvb0aej7KyMYBXdZIG6C45fgcEJS1CxLblSiPKL0gSVBOWYjheJmOb9Aw0g/xKbwo4dE4NXcz8n
hgpxrH20zTdbJeRDaIA/JDP8S2mAkGhftPQ9xy8yxlJnfFR7+XEsrUnCTtzdWt+aULE+RpoWivkq
UDxNF4xJ86CobImhCsSq92/OJ/U5K+pCDooq1rg6p/uXlc5hJj5//c3iNIG8Wvu0/gb9RtC19tqJ
Q91o1ZEJgowGD10pUqdm1exIqdkyu+7//mDVzq8/KqWvqToWn2Ku5r4BsvsrkbpJ4XFe7OkiwKAd
wDpEMxrw24zRro7kbAFtnPKeFiBDshumemjw6o4Tfp0wUhGksT/E5srBda15/pzI8b82JExQlYRT
cjk4lVrRAraWH2k9X20XDgyslqwYVwXOv7WpukK1+KUTwnShOI1oec0mChSlkz0nNj2lPi06DyZ4
T+6wT7M2yUdQ7qxQTx4q+b7IuwunSa8r5NFox08evklytDYT9n21XvAc0FwfsbrrT4VljTQbJ89R
88tDHLnLLanTC4ILjWkEACGAeHtU6czVCwhqkx2jEaw4XwE5Ey5K5OMbRAgNn+5UTaV9vp95AwSm
HgwibLT/3ge0JJ/z0ylG9jAxK/E5NoucOFWg1QrpBPMrudCGoqjqamPgF5Eg8jjYH4YltL06RWH3
kEay7Jtsagatlr59TlRb2y2RfOElXAs5m196+3C3pGTG1AlAA02W6N8UO7aRksiGeHaMCjNiQsz+
LgRjss/jWwiIBc/ipWRCYc4dp6OyL1yvewHJMnpSBiwfHTBL3fAILGUTnNXXd6xhdXLEs1CFVIl9
HSO9QG4hfT/ITlysD2Ft5ucBnFxd+wEbc8GNzjeE2DL2xv3M8AOmi5ol9z73RwTpbJk0V13DD5oF
w4yBD3fq6IhSRej+stIx6yyHeanI26I2YDaHNpv0DWTt0eMpLNNnPbm/e2U2Q4OLtFT9+3WZ3IKe
avpk7/Qy2jo6F3A76brdK7VS+QBCGbn+lcj6jleuqBBA/KfOtF60KsPSf5dpnk5Hc/DhZmiHcX2Q
tci/yKMinK4uN9kZxZvjFlcKWxmp1ZJvlcFLo7y4EcMhuxa614WnQNDiSBNoIQMNkK16kW86vaUI
NJrlOYfdd+9QTBtY8JE/b6Czw+3pPH1JEqptHTW5IbKvJhoidgBuX0twv+gyybA74Dbj1LFdLcJY
jTy/NcqQb7RiVk6ilNS/v3Veam3VXQ/czjgnaQD4QxiKZ2ed0EbJUV4oZx3b/WdR+VOf9hFvi7ZH
demAIGu9Wgk2IXvYhY0Jwz+6NsyloqOav6dDEUbSXeHe/i/4xdR9wtMNPag5/O4xTEKUfquzbdGn
TS43sY47e8WPn2u2dhvtCnEHD0cG0emkd6BSdKGDt0z5n0wpbNy64KoPdotw5JLD/pBxhaQkk/lx
ElOlICx+Qf3M9CnEcHE/X0thhopSJsm6YtBP/gnnqFpTfL9b6nlExIuDU8Gf9J2ar/mXuZQcz803
g5KznYGnPBgujPqcVqkB9yNDiZDpzqqcsx6ba3LXY6ghUK+ysWtbf993SulhICNEeqcDAfLQOEb9
INGM/Wwu87QoP5gUQTUUrBmCI6lzNmKeqIHT6/9zfeERobder/GVAFquWU796zE5iFoGMXHcPxjo
brEgybTEzlfkrjMgYxpvdTJCwmbvHyAqBuyqF/jWT6MUOpgRlmIwV5bPdBIds8xbBwB7TC5xpc6/
YUFmzMdNC48htldVPmgqAZY60pw8nHf1zoEvwC3iZYTpbZyodHEtXO/V3qjxxEE9AMhG8dmK8+AS
HUhGdC0fSl2/wqkDT9LgrglB+M0xoyI4+d19PWt/gKEx674ebX2CkEsNElzB/LeVq/JP3BzmdUTp
hPvOqaeDiWlSSNZeJ3BrOtHEB4C34svaVhJe0ZLca35kJpJsZN3V2hftoBqb9CAHduFWRUY6VhIf
evGnnO6IBvuBrjYzx3dbtksQ0UT7bC5KvcfX9Pgk05Jy3L/wESqTMCGAV9AdPH0TyuE/Wxekwyu1
Ye0V+sYNZiaaLvmu5G8PGyVOzIDoKLNhw5c+VJmqrqu6ak6sTsmmyHqchVo0L72cemvYR/KBTuc6
AUyR/Yyip+eqenTmTQ3u+lrLoxHY00vvKVtPG/eIO8ytbuMIhUnL7Qg7gpfdxeRhswHEUzUSrmdO
uk15gnFRlQmXub/jq91h8bRHDWm98U7eTIi4QG+utAFqOrmDRf6ru3F+3p4NlxIbCvQfhE9yctod
g80GTiE0JWD7VYdacb8wnp+tsZkezQ3FsQhgM9Pd5vu513WRHZ04MydCR9fSq6J4rAAkg2+nT5k6
ZZl4AHeuM4qDtYXw5zAih4ATDZ3PweE7/2YiQH+0nYg7ZuxJqxZK224JirfcUTfOLIy5MHLFbYKU
V+A9bzPs0GNxKYP8/cjE3NZ5mDyBj62rWgfnULLMlJQ4mQbr7CkbLGo0LHdAk4KzkYGppZDH5UJH
FEiwJR62r/VBjRXYBZlsixqgv3jG0WtdHvkEIV9ae7BqzT2elI/YBKMpjSP0Qe8t+78M7oYKIQHv
fON8ajN5hSJPyONVTbt+CTT4WgCprnhvZbhCIRCLTN/jWhU27wudyQX2P5N2yLFQ9/Jp+7F+vMaL
nxyNkfEfF6l5SUCssPtlooKxfBKVenRskIktTfeaNSQzl7tj7bgxjwEs4mCKO5723hOh0TwnMKb9
wa4SUpCDkfmQF+BekssoyslYhllbvPDIymnQJeeQwQie2Km9GX/R2bUun8iICmnGP9jDgCj2pde0
ZyG04L2Ou6kyOGkeauLU3yYt253NJ1uutjEK2vemGzLZqPgecOyNuC9Qr+gzYZi2d5mUesFEGa6P
eILxF+u/U7Bh/LgO38hYTlueZJBb3OywZsIyOtiC2NsEV2kYfjKE5CRZ7erV0XnlelsLWBG/c0NB
ffavBBWMbHrK4gm0yzpNsEXrmugQhIm5OW9sQG3bj+f1PLN9eacQjIak6XthrqoE+SPSrOfwdpaD
90JWUGSYzOeQaMUwfjt3uVfY76O5Lh0+PGKjC/84uUMy5SaH+tBmtp2q9gqcyZg84uB+lgw3jbUK
8v4J9MLmor7yb/NkVogWAMJF3NI8crfyC/dm9W8ZzoYjrPJm66BF8eYKzLRWtH40o9WjTRRFGd+c
ozn2i6XZKC0nGyKzE3ScefjGhviYRu2iHMjRhDjYP6wytrFxW/VgTkgUDoZD+UkDQx4+1SrkCWVY
1auclPGTX5btgEjReC3QhwRGQy6sRBF2unE49eFtlC6eVNI8jYLajFYqNhaBYQpW6yuzi2T48f2z
2jxXzmwN0VggXImezN5faMwTyEhZMEEGbJJuoBVVEU+83YFCefM6V/7zM/B+Q6FpH2xVblH0q1PI
VsbyY6LCdDcpmtmIATdLNTnwabopnH0ZEsfxBrRjGWhmMd5DGf5/lV0L+kjgW9Jil+AYJnajOYQy
utH0n2+bOmGL0QKeGtm6UBc0RTKszB0JvvSiQ1wmpEODzxKamBDX93bPfffN6sHniCerwnEUqbqV
bebyjdghKk9OvEudL0kQ4UZ6fbT6Iw/MAcai6wPebzFTBRktrc5NhoGcs40adEIqit5Vju3BsGIf
a/owZr/pYrJC9cJxPoY5X4XZylsruQwiO9W0jlY74+Lx0ET6uGqDi7e1uo1NLnoq17aEu0kzRbLL
FDXCPr/ZgIK0JioY21flkWh5EIPhPNifK/ejzlXGvPpWCfiMrWcjJLCHSOy8D2lnq8aPV/cI0cLY
PzDG8D0FHKPBbSjPGgx8TyMCGxdP2eK+2+3osT3iQ4TM1IU6eci0x+LKwMbIr8N5WcnMaQqVMQFf
TqYo2EeKf9Zu9M0pgpJmYs+6iV6Ee4zJDN3FU9oEJ2Atgm3ZgoXvRUziB9lcPUw95UUmCzb6iw7i
Xkp0vZhPKoXSTM2u32PWhJn+lTl3xFL9KP0OmgR9oQ7weCHRWkY0fb+FDhKY2VUUmKy44SQqu+/Z
cr2l/W2NUwP/WgFrWqaKa8LvInZHLeSCTGlSRFWImICMKwTeYWfavDT2aEnmx6zmECWoobmpHh8O
ozmCG/dsORIifH87wtErXiw4CEBnzpeUB+01vgTNte/lZCOD01IExE8IM9CyKtL9zo1S2Tb3dT9t
q1LajIMwkM+G99kz05Z0qyr5cGRfDJ4IHjSz580cTlU6UfkF3xNaCirJHP7ENSNKITh4nJ0q3W+3
R3R0T2I21uf7jAeMIu/LSFV0RTlTGCPY9ctMvYQg2HSK+RprkdGDTdwjD63DqW7GaL8w1jxp2UG4
g6s2i8A5SUWDUQajM8baMz8MCq3A9gq+XFUNcGnfm9uCvipP/RjssneYcgB9+R3qQ/1agRGKczE0
/w95Xiq1ZO3/72JWFmXkKpYz+t/WTHdd7ccb3csQE3tPfo9dlj8PxscYEU3p3d4aOhvlxbIXmq5Z
BUpsK7wPod4hu+Hz4v50bwE3Q84QxoYuoIRn5YffqRgXQZ/uX14RI3+8xjzdQFb/W46MUTwCkQND
6YvUW2Yqk2areuMr7xUisntuolKbJ0f544meRhr5JNpwhMRdYWLtKHf63ctAR6IMORH2J/sw+6QF
JImUr+6vagcTij/pmPErn21wd/29vXmFaZlNRerahsde/dMQP7SDmMs0rYZ9ZViwLYe8hcV74fg2
TD3Eejx3SH/xvxqd8WP0qyHgw/EEvuLIngAdci+82sE/mGLFAQZFgPM9ErbUoQUPpeMIVloNEOHD
ZQYzXA9A2oynfmxGQMlTOZe2n4kpncpPhcNflkm/NOPaIkR6uiNhcRh1KtXG4LoKAP32dv5lkQ1o
1X8JM0H+czAdT1LnFL57NIeNVAKuML/pOzstnSMzsY5Yt8Ap2XJwhHJWqfeUCMm+JF0od/XrrX4U
ICNNqAclBWuO/XbUN3rAPctvc4BVkMWMnfc5zXThWbN2TNiY9d0aCmNFsViA8L1qAHkLZVRz1mjj
3QY4UpYB2ASbTpsvUkfKzFclKf9gLiNccdt45dlp4BDuJdTF4D936skcU6fVG5QtO5KQ/PpnbMa4
AF0AhzHaixeHQvwgvkouJHgTy613TSViNVE8r9Cmo0S0NDTI9ouiJOtcZHoG0RlMJ5U3n7y1f3Pt
QmqGSyKyBkuIaU7IStPi/A5Ciwqq+IwBjsNgITVWPMusCM9BAP/pNTLuWRG8wpceHINT6W1G3L7f
yLKj48u76I1QSsZWD5IYaBocvEUd9qBiVoqjWoBrpdtlErVOcIbCn4MadHu2PR7CB9JAaxzP8Bbi
YvrZOPkiJ74RhdI6sJ07pbS0CB+VCP1SquY0nqHtGDc6gFdKoh3HbPJJmBMcgRkG5mwyIgp7Wg/8
J4VHGpU3it4MV8Na2pwCCiQ41kR2VucxAf9ICd1TxpJfKLgX8Py7J1XVp76ai+PIDYcfVJ9GIxz2
uu9hSEjybNleHJBPkE7MShnumbwsMf0xy7QHCNcjaUttOm1+GiGVgsSIb5cH0PB/yP0wO2eVgDwA
mj16S2qEGn7aBkAiMvCz1L4gNJtO+kxu3QiL8yaE+CTmd+kWDO7GiwbR0rXZ/EzhH/lfdDvWXIX6
rK8vjIkplA+Sascwm60Bma2y7F0Fv3QZCsmI1Fj/ASPK2OREPNrDhuRpgieNYCTrpBNcnVs6RMa5
4aMhi8Fc713EX+FQguTwV4IGGQRqnRTzZoYx3vZYfSRVmO+t4lCxSC7eZtc5H5o7cAEMczsVHH2I
ECwQ6rTqQNoPw/8giVGW/YPPQr4yTm01JEOQVT3mg7jRY1cUrdBYikgLlctYahEk4uxNRk8C65vf
BsYtjBhWn3znYKl1rcpUcATIxX/I/BkEsa5duSigk3PFJSAZYqkODaQUxCnz5OZVdxi7NAyHJ5I1
cMoYkXkg0bF98cBVtn4bRWTpWGU51FIE0iDdA1kjrC6MxKQ/N/FBpukH42Moj8u6j+mH6fvafr14
ggjEMQWmFA/l1jxH5P4CgtkHZIyvcAWA/lotytpKX096PUU9xkF40KLG4PziDAJQNqrLKB+vEB21
yI0faRFPxzHAUtnXAz+hX+76pFM9puOZPsFuqLM79oLMa9aFmOk8nWlBUTZ6lqGrA3tfEXyKzaK4
NjGI6w31DILGLqpbSP8kV5Jy9vUY8MyFd8/6jK9kPWie/cBKAiFNyZg4CA9oTmc01gsurTE+3uwd
jVD7EkggPBnIkEmuM/Ek2R0qOCzm8lu32RsfTmBylao6y3g62kPsLbYO6ojv39MThFBisy5r0+Jl
PM6cic4ERuFxJNefxotqruVzDH/fAT4RC2zhn90PvYSyvvUn7/HU58PB6zmPs2XSuZ8OYTg9ZkGx
xZvM/1tYc/4VdvAJmE8r1Esnqc1l+oNZn8dPO5mjT/3iOjROqjpQyLPr7fetL5RToqoPJR+XOnT7
cUieFbt8S4Iyut/0E8AKUPe+aftAMlfTqHXeE+2kZn86VrTygVdcwI/FVMfu7FFD3G8J2oNWP/MY
tSosG7bQObIbS6e9t90c9Ny2XlHrlTLDKK02nsiqYIb8yLqiL54tg+uK6KNdUxk52dp5suIQpB25
4Ko6yR6ZeLA6we3tBZHlRJpCWECEAE9FewgQipT02k1QXvT0bAe++nMnUsXPFbh1oW0q/z6Au2NI
MZ9uzQFOEV1QMpDAxbS8sy9bd/8/XxsvEq6XsDMwWmEgjc8qIjaBsbSU5IPF8L1oFPdEptsFSb55
snh6l34QGbF7oJjqbYiuDDMMgzjQ196hn8LFaO1LI/k9vhJaqNBfzHS1hHHVAPmiTzffhoDB46ll
PhC9IVTpDNwTh8J0eD4GFTfkY6wUePYAenZjXNDhIO7fuLxkRYxjvyUA6CoORVgtqI3c6ReBCGgi
yO9XKAamFKztr2EgP1oEDd1zBWuksixbajV3vAR3T4BcpSo5YGx4QJRpV4umotWk2KMSYY95Kp5n
rUsV49LDJo5NGnzaP7qZYEK9A3qYbV5bESuMZdTTw2IS4VNDK6AxyGhNBTQOu2z68R8tLBqiZzXU
743nWTR/khTKJjZoyOQo/BzgweO1wXi/rQrpgpJ0tC9IQ1gyZ/cLReqZdJ0qgWk3du69eTK8V6mt
Jyz1aBWO/mljfQ0s0Holyv8gCXsCaOPtFiobkmYH5EbCZYIGOcMJKk9zw8yvWxRx7ptYiZs+RsS3
P/tAg6lhj2xwKV1gCRdTPTY/GnDVCDExBawtUS+d6xiILztkJBibS7woUZHGAlmVx4Sghp3XGM2b
mh7e5d9oQrHVWmjrB+xbPyB0T5wrzFgymtVXxSWBfpjzcHG/KHV8qNeKJgiSruk9kR+Z8dUlsJqL
jDGBwMBxY8c5Wpvj4IAn/TKpndl0c6DelrS1sc2Ip86CYss3ORw0f3U11VpR+0X1pFPoyzwuxf0/
h1HE9AumeF2MSZRLAgituAKByP4w4GICBFgV12G+WX61yt0UHlvugmff20EQKddwa3VjaGTNY113
v7wCfLbefpOY9lvGPsyzvRhjvn+y4yFbX5DQoV0VQlgCksU/HlYuu566HE6ES6nutRWDVFmqe3MT
e/T8BqNRMlUFPkjuWqdusU/oisblvtEm7ZWUEmKYG0cvQBr//G2MSiI3ozkmQ+I1/ge7Oft2LFqx
00tQ6V7Lqva0CjY7WJZ9L0lYde/8dFR605pCrU8nnjR99clclzEj3zCWCWssneQP+x2nUx/lfJ+r
XjZSjFjhRLfC0/qe0/nfIjtlPBx+qWv+duIS0IaQVZ42IKGuAezSgQ+XBxUZxNcWvB8X2QVLS560
vdW9vKuAFGUMARmdszSa41StSSt8pP3rytucOS917vsNH6TUVvpsExNMCFUeCrOyVug/ol/2c5LL
SCwGo1sbmj8FQnIhmwttpVDrajr0cTipDjIt0wh6Pa9xnUQGf71OExntogYq/XiSqKzKM+YkPeGq
Fa3Mltnho5gVU8N8vhrpOnvJg8xaFLvSMiyFH8ZovYHXUjxGGDzMwbT+qaag4VBVaR8ttmpvmUod
foMKWi3kE0ArU5lUkpiYALPppqz7GHEikoAkUAd1E/05f8b7lNQ7QfdGyi1Ujz4Objt5BezJvKSF
fdY7bWHBeo2+0v5zxhBwgFze96nWgK3JI5HZ3IXJA6oiH0COOoR9Dw4lkp+nPXPTIf6BC6y/zwcm
CYcOwPi+PQqqkHxpliSP1iJW87/wymCAA1+8X69rZsRxfUzNqV0jZFQ61IYlmj0SXvQRS2KMkMOy
G2iwjV7Nau5iY3ru6TiDAW4kXnsLwpsvGTvomt49vwcy7W06MiJMz6fwHGQGIp6MkLwbpHJ/Ruv3
QNjSOzRVLchMeGvPI5Kd/hfxotWXw/UHrEgcK0qncfRnplWJ0G9Ucmqkm1SozjrWjk2u4CpF81AT
Yc5dgOyTsJcjx9wrdYmCDM6ueqlIqk4CHJIZOWww/seatJeNkDtF5r3e9PN7AOB23lYCvwSEPSm7
ShaoEvgo0/HJPsxP3DdZlzARpyQjesf7hkfB4yQMeUDiqORkLTGaAXiIIVCtEyaEZD1VoHAV3+Rt
leaJQ3T0wnHHZTaPJmqp8X75knM40VlnWa2Y6P3hmRytqvBetIVPnEeo8KlXNY49AKkoa5DlF+Bf
5TI+xF5q7Btunqf2UoY4V7jz5FR/G2kcYIS9fJh2GQGPLwYz9fajkKWpnWhJiN1iGsbXXu2lwW3L
CaY18kWUN3InkGayuWNQy0f+wsMZRRWhqBdLs5DUIFB8lAgYWMK9loOLif29LgdTTYU2vFN2o5We
OKTjLU/ROIunIb7SZYOxSkpPr4+yjH/EXp4nLBALkzKI9dyMXFoBlHFuy9zzQ7KmeLmocaUBHPWn
mBj2wxCOZgQcKQeMkm7bmwSr63tKOTLfETGtr5wYIt3jag+fxhncJwIHsuOrDwNb9pP5hRqP02I4
T66ebck5s7Zk60iI0pWAkxi7G+n0obkRtEm8DhD4FIIb9ETcPHY4bQx+xR2BOcrLIWmRGJCajPdp
jUKAm8+qvq7fN6Pj0xlAgyckx0jbQrp3TGgsYHHsS7A/QfnUP0OuRQsBGTRRpSeB3dddyz49Ic+k
4KC4uDYX05hNJULnySSakXVFLQEahKG68+1KjFwZdVK6nr7s/BPn3H5DlFnEJeeVpzjZr0+4sWcv
mBQhf4HD5For9+h6IY9DxKIhLVYrtDolU0a2Y3zVBfOueJLuley56e8c0j2zPNZTtMc6DiuJG76M
TDE3OL/xkmjz5uMv3iJgE0bJFxAB7PhRjj7R+cXiT/KcMTXWPtb1h5lMie5Dqne7Ij1jOvMCxHjG
AfUfRVJbSEwx/GQ6l7nyJzBnTtYVR6yco4wCfCDQgNEpjK5O5Hget7ttxXIyEdiYcAGYmb+TRz8H
vv7lhrHEcFT56DYqgoZiuD4EQA4KpBUHCgM4fSy1h44MKKdN2xvXYjcVbcE06ESPYmjBtw/46xqc
armb7ESso3+PXbfjgLpDht45g7Vwjmzx5ZMMmCbn7AD4GUR5awSjqFehkp4xqCeHVruNXCp8eb4k
M1oSWt/PChOc9RHlR9sZWfy4Y+6CIADO9LDVat7vjR5OXk6QkovED2gTFRjQlLvVRZwuwNGA7x74
YyOeRen7QFiJ5mrnW3JFNPGevrTXUK1zDp6qpPptT9GxuGKuvjPN+Gy521NlETteNyN/+H5pRTKT
90xmdggA98ppbjin5Gs7unD2tk8etGixdJnb74XcHbtq3TFYEA+EUEy11hBQjvho3+AYL1NtWR8p
ZgEd+ltPM0yKleyje6utSGkL75HQVoZtxulPkufkg+W9i9GlJRnuoZ+A+DCy3LLZU1Y836UuwhfX
KRk5rByAdQ0gk25hmD+7pQXIv05Nuhur0hv+kKGBvXWQE1/CI9UAfgO90OCQjMaKVUjQqwRginMk
FDsBPVYC4wiZtbexmbVttq+re+Y65Uz2lXPESWU/xZYwRWu5FkyDPx/spqSxaDEXBn0LcMBRvVAy
9R4udKILzjqwhzwb3Tc5LxFDoKn1mFcGTjkMwIb2ldseIezP9BC1nqTxX3N13CPBh4iffJE6Ev7+
n+/87xEKWFFV5OD1Tc/+KzPTstxjUQ+3JKtjbOVe5JA81Nb2uW7bfk3wLtNWuOvgnuiu9dqpXmPv
apBY506oNIYX49swDzBEc6f5hzb9708zzeQgg4sshfLU2mnL95QtcppIjzSpb8pcCwZ0FzaENntP
gjGzCnA0z/X6QAZSXtmq7R1z2uRISMAJlAPFQ6FnFJ9UXAD4gN1GVNRx1Pfp7vUDZTcG9VzSUGSt
TOT5iTaTEYB/aE8hLK0m9ksrkMi0c13p/+rGis8oJx2hOFxLHX9FSgNj5ojKBvYbShI74IvBLYVN
lyr/J7HtHgL+MabwKOC11JednjYax/fLryCvgkygUVs+5sbh8Q2EkuigK/M5pKS3t7zoiBe4mXMR
I8HDIYN9vSwJ2MtCODZaGqh0xA+I/QsDh6UMdw6SDdG3SwxO5zM6ZZBpel+D0/CIkBQvMzESzTXJ
ETppOh+7gob+9ATkfvJPc54beXh+P/ZzziECYxdzeAjuzll59xO/ubCIWAiQRKmZhRI13suI9LW6
S/HsXBjnP6b2baHAWJPtGJKe6cp2h/QX+IbV3hA9vOcA5nLQb21Vlt3IY7/o07bqRXg8tA1uMFvA
qqvolKl8pUjJkfM436EzagZzQwYJh6S01n43E7Q0eXulFcCtmXqHoh6Mj/xfWJO5nUw/9+xzalAe
XHzvxrsiY01vr4We30rfMylkPSmeMuy7xUlGr6gsdvde0DX9NPXC5Q1AzwUWqFIXDc6JgpZG0b5p
nUNXAEl8Qk8Ezk0ZYFZs9QbVO/17kWNjYVYS5EDKQUTbqiuDJ4CDAO/xuYIF6wwQXgMq6e1Yf6hO
tfy5DrxBZaysIq6Oh048wPnKLnbpKolBxR6QE4D9gDsNChTNyzQRDJZQxJ3dtln3kVFtktbKHzPt
wJ/ET5vg+sPnGLfH7RNmXbGOpqBYx5GY1AUo/XK+Skd31j2eFGjux7DTEkbuTbxdwnk3dntq+a5G
Zlq8JIgYh8oDrcKOO4n1UqF2O8w+VKLrSV+1uRB0kiAGXtVUBfrMPr1kRd/2Ze0HfM/8eVR4hgFC
6Pnys4yqszQirNWi3w2m//uDUlD1DJHICTen0Fw9LIx/8xbkzZuOPA3pKteaHc95gvLPmc89ZpCW
aTRT/PAPR5VdiVnZL+0q0+k56w1aI94BtNbx9dJXNFPVCPEl1j3T4cvrdwg31b+K6jBdyGNbN378
mprN/jNMwZmkJ6KcPLbo0yDpURZnwF9IKGuyB/ujCx8X4XxflKABEa0eNK/8aa5TjyF/n8UQK4p8
CcoCkfdVmdX8UJeS1JUMLlrCVgYW7YHnVOPKCoq0o54VD04EwtQSnuNQKhZa0F3OfT18uURAod4T
Jnhkh9o18EG03ly9T0sJsQFzgy0iJDqO27srxQNq95Vyr6Hqm2Xc0p02kktxG0Xl8g3GgYuFf/bv
T3E/6MGAkRi+/UT1ENAy8/qmEuv/fHY8yjr8HLa/8mbPtQ4fB+Qmy8wqDcB+NU/9gmKk9fzDTDMr
+/vLNZq4xsIcRZ0v7Nn032TGzO3hir00igFmtDBp4KN+jVPmR3DnwpWRdy3Bo370q6HN79RERsUy
2UCFN1BTG7BV6QsSheubHxk9dlJkjTZ5vxi2/KAW0Oo7iVRKNELm4Z0MLPdTMjKAekW+acdydOK3
f6F5EODeprFD2h7zjWZtuvrjOXS5muCQZEFxrU8waPd4YJFCha/yvO0+V/SULuWGjWfrUVhx8a0+
ILzCVUno3HDAFgDINH73g8RjtA3QnVWR7vfPhPvvxRlUHIov3hssI7sqK9O89HSRuz3jO15selZ8
V3nYyfRl27kdJWfW8LQxbdoHXWpkDlpzT9E4Pdh5ctAIwEaBwjxcMj2ptB9rVSssXGrmqRv+02Ne
5T5GFG4lzow7xIfJeXCH/yFrarA3vT9RdQyK4DELwamiAbtr0klWSddGBMWPHYpe3PXxxzetp33t
F8TFUB83r2x+nzAPYyo2vzRjhirHY7Sm4C3lWxg24tDdJ0XDhe6woxq7yDR0WUtBrxrehXtNrDaD
pK/qf//PGzgaHJBQYlYsavLq93DUNlQ+Eod/HcYswCdmqf3SRrvPrp7uRVEyK6sq54uPILKReq4s
k+yIVaEqBhYkRZILlfiqyu5522t8mXE5yLubp4QCoxF/8d8LB2PznI8/HxCtRu5YzM762Q7calDJ
bzpKFkG/QUs4CS9aajOzl0YTsy81bS+VxibQJydQrbGOTf3h3VbySXC/R7Scz7gcTIW0mHkI+XId
Y9GCXxDMyqLBEi5XFyiw5OTobea6T7prf0dttW9fSMba94dtiE5JXa00Z8VvtRDam6KTVE0kW6E7
mTWAMGNsdxVGT3Omqzod2npTOTjhcrsXm7DiQ7AHX+URLWAZDXXqfxXwWCzijCW78SKWGqAf5UwW
QklkvYgV6mdrdT5vhG65RZoC1Xgi0BO/DIMaNb9+VbI7ZSWtY0GhmEysTgUNBr/aLZMiNn1eNd3F
diQWWyriYElvPjnpcsLEk02dPUdqmoocSgsfZW9sPoeZQZpJm6zvLeNeX8LX6HNDNvJS8TYuguRP
gUwJ3iTFs7hLXdeCCnvYZEdGW7Y9Go0EPWGBhAfwJtTtNsXHDKkQTWL+sCRfBF8vsjvBqRLJwD81
sxLHuc4tFzLS3J+0XHDO6YhDXZusJN/FfyYDAmxGcgIKTbBbnD7BHAdSHAFS1xe8VM/mPLQtPrl+
5QJVrsBbR9pL5tygoFvqpVzYeBm+4SnLucaizkLOzjFjYk6cuTXzERG68joSYPa/pA9VReVaRgN8
6UQySdj1dV9Tq91Lv6BN9BsD0FHbVXRt87B1k7NvYp0waG88OmrE9j/qD1Xa+drb8X+H/MXHCypv
ClfcYC1aSuXlxf3iNfmmmkGNsdnJgBlKDQs6W5YcFj9CzZQqUKwCYkXRjZnrxJJKM2UWDpi5z9dL
NKBRbYAgwNW7E7KHUD8lFTIsxGxOST3KRK9dZa7LF6QJx+Sz2akOGa7kMdoQpMZHCK8cZhhcpUbY
SY7AhSqi8xqcSNzx6wzVudtxx2/bfUizCHDjKNOLom3uKaemBDqzHNPhCJO525iZHOK1UHrIWWG6
SoYZdCFz+pknGo10nn1Rg4LHWu8sSV0wq6plFJ1HgJnaFMXtGFxNL7pEwjM3V4kjTlpBTNjhh/Qh
RTP9ar/4qQ6EAPHgE6GxlugJV0+98Vgu5TvYpqKEQNgDwrd5qa3VIoCXTs54ipYAv0nVaA+1m+Gm
d2UaB8XWeWKCtFTxT5VYZJHh2L/ejO/aJ9YZI8vCVBZwD4n7KhVMlJMCdG0xpN+FELVPHQ3P+VQh
YdUkDttJIEhcaA1nyuDOPu6iNcaFr+knAK811ldE5cJNfOSYfu8rGOnBRaZ7QFWkWoaD8NkOH4nS
g1QlAFb7A+SpghA1Ry2Iv99Y8d+ejjzjlFaU935e9pHcOW8jMLNKbxFk+HvOidinYBtPdMFnz8jW
TNPiGHbf5al6JImNonzkEjHOvPJQSNKtu+hQfFwnGF33K0NEYFfPCtr0op7HskAgsZm0IrRmgBQu
X3HExr7H+Th1lJ87na8QS5EodiM1eK78JKPzQhB37kWL52KYo3ESIKXp2/vYTjjPSo8bXxZwuwCf
fQg6WPeb16UiwiQvcmYOmjQZfpLhxaKWxlcONV8v9SR2r0hzkWBnBOEkTn+tw3i4++fdCZfxlg0G
fL+dOr/jtHEFcl40xSbq68GvMfQLSFxrNDiRjKX0WycMY82mCZtAfoO19CJdjVgmbGK99prNmICo
5OPn8cboW94eiQ45bjeFSt7GxrIbco49HGnRCOe9fvnEwe8ZhDu9LkX6+hGFenGhruDoZ89t5POD
mFAsqNqeoZA0J/FjrWm97IfYPreUUSYHSJgbqB6ISg5/BOpXUy1dNfa2z8CfsJi9MgqUjYJbMRCc
2NLOV53AKLBpvdVmizGBB8dneM4rmEYHn7IJa4idsJWuch+XYqRyZM+cywSP9zWydY+/m7nw8hlg
oFrxW9EsKXHYeU/tVQ78R37foXyJCvTZjo5JyASZPbU5je0pwvIZGxPg4n61cM+GiXpThvSYFDu2
xI1BP0j5Ff35nhxT2Boi4yz5GrTcPjFDLB4fX3SISar+z4qYsJs6ngKm7vAOEGeZyjcq5xQ9HxTw
HakW+jUbpydtsh+yOgL+vkFwyrUwWdyRWDHWM5focMiPp+TULkWzC8TwAm9cKjqApv64HZVbY10k
ZpRHC6XzNBS7Hmu4NRJhmirDzbkPj2mNIxDLiN7xoJu/2BQxXlq15Su8MhNTOeyID+n2CKC520DX
f5z97HsNhFFPHvd/MtL+P6btXzv4s5087N/hBpnCc/eoL47sxRKGOg2p7romUouP1+UpXkPKxuel
opvj9xQwJdctQVRaTdEdqycYFBz8BtLhE2sMMNk3SwUfNor+8layPeMAcbrIsED+hw4FSYGiWsyp
IP/r+XDZz9QHnCY68F0joUWfUg2ecbFaa/ghHnqugJ3DcfNp4hCpowH850r3WWOaC9/63gtTqW+0
FsYrf0TNhoOBpyA5xuq5IA4zgeGAW/OvaJHHlIcnG/cTizidA04PLXENE23cSA/iczZJeuF5sK3k
YeIDqIcAVCDcIMPgMxoK1b94LK5h2eze5BlWQdTuezGqW7b5HN5KN8MVUQ7pER3eE6nX+IzaIFef
Jhn9PRUc/zSKyq9pzVTbqOplFmJV48VRshRwJc0bQaO9Cyaj55I3aMg5FL+MEVyiS948xyi7hDAg
ai2BV/saLykYH6NuTDHlQHoiVGfHJU5Vqd0tcz/iw6vObpwmLT0V3Aee7ms/6jIgUAyvcgyb2DJP
wC38fzCvjvzVreYXq9GWt080w5Z5nXRobml4LIVPFGDrF+Z7q5vEWcqha1aJah+2/CymweCjAw9+
AYFDo7fEDW5uc2Q9ymGBI6QeO7/w+MCOQsqhVUmHWFIGVIyHCqlLVvErUE5J2uZUDYskDDPINvRG
U/0EkfvYydMV32MDiXyGnNtr/DbZhqnzk2NZsEwsUHm+LEXN6Ohp0wegZpJ9/X36h+66nPtp4sMB
Tcq0y0mlPQEkV059BKPcuXxcypZLiopqHxgBp0M/0yBTRev1fKfrQCtc7gYaxVczZcTspFY1G7E/
jeMC5jpR0SMLfMgOubkSpvP4t7SPQ9LfU+vufrzXoUZjnZuGIkW4yDAhzwgJQCWsbaIuZjWlLKac
NeNyBPGkGEDEbi6a08yhK8D/45ga3+g8eBfjL0gpmjSLqVGab24BwSUXYuHh12o25VyxEdFAf7QT
318jBnkWPovjtD7UuUlea0oA4r6KmQV2nTBP/b9ncqB/b+1tgVZaJ1UzUb66rlDnBf91L18cGmo6
mTr0ZXVnnZUgWqPxhTrgJj/YB0DrQRUXq7iT19EfFojZud/rSyU/vyBnHD76PNp3FV13imfpsy+8
Q7S3pC9fXbbELRoClHZ9HDgMdfVmvoPtbqCIxy54JMBlK1E4Bd1SkAGpLcODbEv5k2g98u4LmkDR
fYHLhn27l/ThdH8Gb/5WZewyoCLYhYIxdVGI5+rN402XoTenLYJxWJ3WIPiFE3mDs0EFpheYojDE
igEEvPh93/Co1cyuOrlbXj2AFJ3ACqRbT+4+/m2dqZpg509V8UGL2hX4rnmhoVPG0i/XirU76Q7X
wHE+VXGf+a3DQnRueH07ehbhrUggGw8cmUlmyL4FqOvuEPx+LWr2b4yLEQp9/RsV+Vuil90+rtOB
K5cCKXoc5HhH4OaiW5iksVgmWk8z9BdAYY5NnmSyantNM8ViI5j8J7XWN8B73RYC/EELio8nwNh7
9wZyfUE+AcCU14g4tKVjMptTJ/ZHCgkGOHwb0LXMvhQSsf00uTTZ1Elx5WL32C9mTOGjxLtGqZui
0Yv1sxpSSMPMTMo0X11rsv8JFpRSYySBh1iXExmjMb91bNFKu77WTSETKUWLlweUjvdBeOgjOeTx
iK+LI2dwuCex+/0mCa4JcXm4mhDG0rV/EgA7ScpzjPazcDehL0oP0Tlxd0I1/oIky8992btWeFFy
IpZ84LNyKQh11HTs88UPZQq3A8F6hjbLUP/I/At3MfdqtnYSUhRg0XZKRlMCnxuAiCZVmswqxzZ+
oco2M0nre1eJ6E7uYeRFj75rfIAJ1iP6/n4wRHazKWjq8gwjO7n30avAxNpBycm5HYVdVZOctv1t
mMBLAZ/74wA4Kg2pw8Nc8xP9QxNUtnaGNYQHyHgALBhcjV2x7tNA1r2noN9AqpIJO2ffaAvMmwOP
0KeR+ArRK2wbkDqmw9m6vcSLxA7S71VnG0KXhB4pc7cxY8oN/wRrYuiYgwSxK7HaP4v86Pbs8L5j
GOesv5ql2vccBAlY4EAhmQ0hSx41tYn6UfTwNYOoKKdPne64avXFIiO9los7rGld2Ga8cfBDlao6
Sz45fbqzN4UpaDd2N1oLQ0P3KtDYysIcC0Drg7qwnZ8l668NZUHhTpSUeMsQ7mbauRSpqHtwLBbx
/+ghxdLc6IETTJsGC2c51TqILXxNhVjJkrNg6AZMpCWtQTYTwgCaaS1DhqCPASdxleO12zF/OMte
33YNJlPlw7fBpGFrmkNwg7FUaS0vTcmpApTmBpzFJdjBjcyy5Yfy6N65h2Kba8ECrdbIom4a2rZr
h6Mpz3W7iB/Ytxch7ovm2lElP28nQiVVCU6lR2YX39i3mWAAB7oQX8xLhChEZZNLrciti7EtdS/W
R3jOYUcnG82JDucRYy0DpZo3BqzYad0wXISuelPxKStCp8EeXbf0Wr5nhArZVQGSBwSssTXpjFE+
Ow62Uy8xWacAYMenBQjx+BNCzm6MspFPjOxmKI7+OKiW6ODIQEcaqBVKYhxB/PEX4zHsyjL6oEqw
qul/if1HU9xDViuL1Xjeve+umv6uJNdY+Bch95ThHmq2HggvRmYvhW8vR4YF4x+UwDrHnqM+k2JH
dTbPcgLAG8EyNF/NlsbWplg3PJqnSywsD3vpgtPUEiOqsK0aDxVSQL9x3XKTt09CWyxJpRf3zVMY
vlWtED27jAkEB6mVaQ9UII17xchF2f0jlrIQLdp7m4s0ibZPIpMVKQF/EMQBRC66DYHHGJnJmy4u
uGgtKTwwnscRA6Xah66tl2+ufsKFy7R15Tt2Ha/bEeSv3jVkgstO+GL2dPshsso4TaGyFP9/NoW+
u8nWDC8JiDQR8EibZ0c4kqE+3Z4tH9OStygD+yuMetMLnq3nfEosvPUOcAL8sBxPip9FXokoJoDH
Qwse6Pbj13TP885uiQYtuR8XNEUp+PBY+hYi4ATnv1PLVSdpxL1fHWzVmKpGNDD8FSTB25iISpmz
UWobwmkrAnxMdN/IwKzaOHjGXQ1KAhRX9Fd1SKVsAZXQZXrDQIbv33jH9N4fW3yvLwAQi7BdslGL
Eeq7yMK2KlkwlRbXlZk4nkI9IGgnQKpIuOMRm0wlKeC7Vc0M45dNPUkxKdcxl9hNBySopb740kRE
QLLgoD9S+xv6O9ZSqGgnDubFdFO91ldfLODtW6ppASl14EAxmgBYjoxS87yjy9Oieq+KXEplaeTq
ITX3V+2ycl7b2ZeBIS/FeVmEHuLsvSattHUfCH8qckihbpgFDPXBnZ2eSbw+sOScRHeEsKv13q95
8ZnLrp+0LEihPN5hjSR6Isva7esYvO1Xoh6NHCVp8SVIVdYMxj5gSVYUiojvlL7AS2UZ3d6EuLn8
OmQQcker97w0cWVmY9GnaL4hRVsybovrBuli+na7/tgM5cexIz3d6CFGyGfpAvPfaess2CH2D3O0
I3IdxulvuQ0W9dKiSJD7iSY27TtJkvEM5Y9YzrRxNTSLfcJY4ExwOo1uwtYKMz0DnANPbVMy1Y/P
pLOtCgF0Q6ZUr0r7f9RIf02EECIXytILWeLMOYgUaiP0Hfr2KIlPsfNYb04aUCN6gVmWwL0Dz0Bl
02G0iE/8WbXFUDRtgJnG9gP80mTieTAv46IQUDhJAiYPxS2Hjr4nDNbJdMXY+BABR4P96FvkMZPZ
2PrciAOZrjtw24G+dTKgTC60tFh08flol+tBTEJiZloj9Ne91ydcYpIVJjn43F0xjFzqA9h5u3lB
vZwaLAl/y3lkSsjthai8nt9JLqmaFMQaMKHkH0w2qu0NBFBCJHvyzNjwkW5ymh+YA1TbuDfehryQ
fbPhnlzrAsQS4qOg9jah9x7R48WhJgAA2p37rK44kY8WP8jSOXeT1kbhWYBpBMM8kJdSdvOD8MeY
ucpFjkfg2c5f5f2oeaIbu8vMeD8/S26XhM5vFANjMpIHVjzYMvtMwG0KyrN9Dg0OnzokHcy8Yb/o
yU6Axx/o8Be3JQDjAfHkE1eLKOaZNAaMMDYiiJ7I6Wla/yn5DR5tI4OjJoSmbX8GzrsYtfKCo9dO
7f6tlio2omgVr1zd6eLzVm9RA6rJ8iUQv6aMJBOMtyB9/AaIbdpGwxUxUcVKHgxYwFSTx5b/kkDx
5yajdy1BmE0rY4XpWBtwFAQdra50DLWDdkQahFvBNAHU/iNb/HV3J+Wo7dG6ZakYkcmvPXt7giCU
jcbx2XLBeGJ8gzYZryTvxRRUtQ20a/oh0CsuZ4y6DdevCjlDlB3g8QJHbkmHKB115TCGBiuZ2Dn7
qsq6TCMMwlRY7cn8zkUZ1ZPfLS/ZD/m/miqPfoPZmXki24aiTHvE0SNVKxBXeF6QispjW+zJZVxr
v7oDxTgv2i2msEYAgp0aEPOeFrVEOdScorOrIUTdlMSjPHmxPhgIDRsdvaLyRceZxY1UiIzhMsNE
uEC3QRchUXYfQizT4EMLqs4aevTikDlOISQLU0gbsSgbvrFxJCg+mxHVJAsgj7ta99vuqLopQmJQ
kO4fxsiZGddiKEqFlUvFXJjgjU0xU4MpjXYzQUJ2hIVLSjGZTohR6TQh1Ke1kExeR6rdHpNJB8VB
o4KUtc9Y57c+jbzoWlQj6I+dH+k89jvOkqXdVpShcJX8j+vSwZCdY7f3jw0B9Os8gsHK9Y75+ZBd
uPTP/4t7AZQhk/woyxjhGqhrf7aktdG9YOS9KKYbzj7rAJ6kyo7XEbQSDA9LRdz84+yTYKZkaMXA
0jspVvdEPrk4tDH3+07VwKER6kG1JaioEj5qEYJd+p0WwLPvpCnHI4yZF5B0OglGrc2FttTe2J7s
pYq6Qap4EICqMdK3bv5nbQNWv0eW+HpSFB45uJe/Tj2mlp61a5XWYzbnLuKLamc7YoC/tQXEhyYX
2kuHmxDfqXYrwFCnNoHTdZRs3kABvGuw6a+Yz16hPqaxk0TBLtJTFEG6/JBxWBT+O2PL8CkdRG+o
yiIPOw+dxMe9nQwm9zJjgLRYUH/x10SlGvIXceUPLAg5bT0ZsppT4m68U6oJ6Fiem15zLiT4hRxY
TCJcWEics+2UMax58V45n94RRvanwQ466IOWwUGc4chNPkcKBa/qVaBOeUjVwLA39x903JEe0nDj
y+u2180xMLYRO9zlV8/1yXkp1HFR+4NFJt5yXknA9DPXyQCvkKz6zNTi/smSxOXCy+GNXBhvGtO6
AREczmjibXqglgyRPlNMOoNZ2BxH5QMrPExvw2aF6muw8zX6sUUa7W6tryvm0yLIllZtxAhdmlhj
3dqvGyRz4IinqTAdRMhjSjx1BV23qdrmxrcukzGCK53yay81V6QkC+lbn0wOZg5X8uVlKPDEXmhN
CLqunSc3OUGM0++wLxpsF2u9loUOrQBvChoBB84DMFBuPAITAUjKpcK1d8/Ga0YTloT4ame7+BFv
p7rmSxNKGl37B9XzWozObBh+IbnWh59BAiuaOiPgMZ22Hqw+ANKVCr/YDKNJ5kPaB6SyUt8dxEXE
yuLXn4b6N9R6wahYTffz+ywv3qYe6cKgHTZ9VLxTuEwQX8UI4ql8wmE4feACDeZVtQKzEACtwfi2
m+CELisl6ZJ3TIiSkJtDeCFFT2MZduibMwrih4h3tjFuGMS25nPN+477QoWLrxhmWipx8Rcxki+/
b78/fvD1u7B33iaUFjf15/qLiIci+BHrc4IE6MikfAGe9DJVrwuoAt3CBe9gPFEFKFeYKJcWTvCD
a8hDRqsqJffkcsznu0DH4L1Slh3M5QPGjnkN2YeErFVeDLg6rh0MA6Cx7AgU2I3Uajjq6boKPlCz
0fYUggLTZRsEQDF14xf8KbWq/SqB4JB8WLn+74MYT8VL/bkBXP3oIIDlvZmg31X6Lv+U23ls4mE0
paFD2SYxmNhJf7C9WOU/XS/+d9UNQOsGCuHwzOfMQDzvWYkRu0RxNEZhKgiZh1NdBd1zhQ10xe9e
RvC1kYHIino8LlZzMbwOx7RFXnHjtZquSFVdtnQhs3AXp2eEgM2z7CD5F9QhLGoasR9w03reaIg9
CiL7xsnvEKnpiRpmAYe1owRx0q+dxlB4tiKex4P9DHPhfvfMVrSWqvsHgP0cUIsuMZEJJoQDDcya
/tkdQa9E0WKQqA8CnFrmMlLGcP0qfKHnJFC+wNtz0A7kO/K4EjXc3ShlV6W0truntBptCaKnv0I3
59K/FnAdsfYHDbfPZAsz3+RLIvQFfeXS7pfkurqjYRMHz5M81zlfaw/UyyZxRB4vk1seCuKsQPyF
fHKqGJXXMcpWHveraGYrDnjYr3CeCmozzUpayeSRUwmP45gJMqVesFBDxxepuOzdtIzXPxvWFrb+
3hziMrbIqrrs17kARfuxiTD5IuU+FZ826TNjvtp/ehtC6Hq3VLm5YzW7K2LQ343QI+EyysANTfKT
+mAq18vKnCf13PV2dCOwdnQ/u7vCQkvaWqwRF7Y29iOVkq+Wx185JXp0jkFUIawvvxygS/vQGZEh
Uzzf5TpPqEcouPn25d0dk7a14NCDiJz/TJYxhBHb0exY1uJnb/fsvQMvc2ebSeyx39ETHmwgJJx7
0v045WK/LzKaoigf3OvkWiKcV12a+TBxJT+HCw5mclWaOgpua33sBOZzrxweY9Bj5rsV5UeDIAea
GSjg66rP7JbMvzle+27i82YuG5XM9/JhUq0xla+Y720P0ymt59U67DBT0Wdd/u7GkiVlDBC6JePe
Q0TtcFwHQaiL+XVskTE0cly4bqfH8YMAzRwJPf/79e7/FBPgNhLcRVj0A4+k85F3U79AdI8ItSQA
ItIlecW/ObtcS57VTtOPr3vBphWIDRZgGWuDqVG3/Z26Xdt+eify57nA4JZRqHqB7U1hyZGzZZ0b
g2dJNHFd2JcO0fUwTk/fDsERJdsfOx6T4qiX2VegDilEGhewr22RsMe63tg8qYnPxAqCS978BuRa
kVSTHmfWutolOHP6S5Heo0DwN/zvvQbgK1pghbY9rIngU8q/+s2+F6zsnyyPHv7gQYdX5NtlfRDS
vq/A9dUqqDHkPs0O/cZJ+4xpF0YdJlaGLIGHD1F4wTo+gb6Uz+/qBNv9Vo+CWTxLpEHMa+QBN7gm
+NecF+XDfmljjjTvk7W4IG97t/N0pzGxN7PnUlZQRaau4n5ewTECsgkMCVf8ObPlnnlg2uecS0c9
e5A0Wxnn2oTQp0YUIN914Ie2BOqI5e5Z6yXi5wL7paSjdyZp4BAglCBnmkCCjXcTwMUm6bjOzJ26
JJ54fm0WLcHmGndKF6T5vysE+pyCiPeXfuvmqcuqSQmm3mElqaclnHOGeIpAlday/WMoqfsubE/o
2rWk9cPBS1NYWg6HarUzPRM0QPVS6IH7cvjfLLeTBEDeXaLSF5N7VCws+j1R9K9ZJEQGTUGQPzwr
vI0CsHyDLSBtddFXO44qo6X+vc0MjLizA3e7xv4cz/O/cR+A5XgGUKG5xYuqRM3rWtYaBSiWuQhk
E2hq9Hqvd0Bi+Z+tkmBdULJOzYjf0DNRPNxaNbuhZHxGdJr3jLkiGoQM/1qBo0cnTVTDDR08mT8y
pGCgCj5TP/a1XmIkhdVtGXwiAc8477LbVh2eC5CN6oNvqAVG0NU1bPBVLqZcQwWIdbA8puOfzhxW
PtmzNF4XGnXRNJDZv9tl1br066qJuHL4kw8ruVwOwoN7kG/Cjo0+ToF6g+9RxCY0thVVvCMlniOm
n2omzD5NrDBKIxSTT4OLRU9QIX5q6t0KrdfQYJJGiKl7gj54H0l7PYmWN+0wHg0kVb6Q5KhhkYnt
d9W7AEh9ZLwgE7jwsTWwyuOJxwhCcnmXDMc6CmsQ82VA1OkMhHgkgenCAntYUCHtpj3zbKueNL48
BwpB4fugujRA48LT4RBDRPpsNUMulZ/yA9tyNaMCh4ZcXMfU09Cu8cNweDqI/FSdXMjJwJx8SpfO
UUhHGrtPF3UJaexpQ9wOUUQwn4b9nMd2Cm5QXKA2JaS1iZ8WnX17V/31BKFlr7G7IrZY9S+PBknZ
+7HlUorkgIobNk3AVPCDJHC3jwOcWHavjylpEBRJCCIMknM+JwjStbLllNFpZOJdD+tFn0lZm+54
+e18IxFAPXOp1Ut7b51L+kUslP/OUSOkjLC6bwRyUGKas2R0s2F8RqmYG8b0uquRr/g9k40iX7O2
fh6mRzYm1VxH+/VdhIGW1KKr3mixndimlM5c1YItOI6BD2nLem4ip6rP1IEuOMaJYhAB+Xobo+29
+TQT+RHcip0E3/+QrczQ26chrWETzxU9Gm9cgvAYLqyARL3BRQDPKTQWy1sUccoxASxPFuQ7DVKk
wiQOz2pl/Sd5z7CQd3ikcjDCj05GwOA/rP3WQzKyPHGdlQ3qXWZZCm+NmuIsi2nV+pYW82P+0E8T
R2HyvphpnVITM4ctlHWncTxX3mdNhLOSr6sGNpSpKOIB5WO4PA/HJ94z9jzpqXXM6I5+pzrekA9X
QLoVN5hoEEFi7+lhiwY1k/YI89RkSXlwLeSloapAJPu7U4RFo6/7SyzgV+/vG50CrBpklx2M+JZ9
bMmcgodvzChPshzN2OXbCWMRgeJnFwXEhqOND3wGkrHXXmVLQBqRKoOgGwoZ4+yDBt/l1v9nbsni
QaLKUweVxSAYwJFMB4OfFFhD+L9Zu2K3UHanPt0k5S197C+4A4EMibQPPLxEnP+AEvfl6pnzxvtW
OZZLeWF9qFeNfU1LFAF+ZRIAsgPbW8/6F3YcBqpID6ZizW/QwcF/9CiHcDgQF8Q5+8c6zWbUG1H0
BInD0+KcZMjlp3CwA4HzxD4T/u/dtUJTo49Fy1GvhU20ilYFlmK+MAIOzzUcuWjzj1Ku/q/pBvY1
ZJ88MOEeslDsp7MBDZvX1OctXw1CnMKylzAOX2zfzINTlDSMToe7CcWHoZ4n9KER0I+WkOTl4Ch6
SRPyUK9l7lBA5UIx/GIsgZ01J6ogfdhL4XSZaDjYIY6dJ4C3UlwJNMQggtJK2hBfzo/HHzyaOIWL
fBD1e7WDKeCsoYynBD3gWgu+gJZkSKkgIKBMe9cRZLP2DFAU/tApeiNfQPa9NB+ltj4N3DENvWBr
yeKfhN0M1bnuomIZ2kNDNBWcEvm8ZalOnzfC6k8ULzMyjrIctChMSCrQvIUeA76yNqjd3r+MkPCn
/xvYAiw4ctO/yM5DbB2fSlkc2vJahFGqXm7CDLHaKPk8hdcpfeFdqoLYsAqcxdkFdb8Jsj096N0Z
RaOMapC59RrXQlD8HoGuz08ZOxJxB0t6Y7c4gmftkYM0ZfSd1l3h/f80dVlX1nHoXo6MAiwsVuIM
Oth9VqAbTDAnBEET7YchF7kFB1cHXqnjQdMhycHIoJSyiyO0+zGpF7rMTuEY2shIGpFMgjnY/L/l
IZoh1ZJ2zlqqZjNjnO/VMVnx6Kpdorknao8LRhwo2boRsQYuY443g6hkkOupnr++fLdi77lT3Xd8
7jhGhIasgiRENH+ShHhEJPHVFmCz06psoITbdWQxoWDOKVmFBAXoYz50EH5LAyhgNCe8w7aIWwLq
URU7Dxl6KRWhqd/xKJw2Sh8m+mPbxLds/0+QiV5tnW9voFjEW5xTWGWkpBRKC+0hUB9TJTcdFmmX
JCM+2qYbRaFcICbA68z26PKTGbzTVn3s9HFDimHJrrzhVlBEaGnV6Ts/ebFMF0iM8OJR2GB4UkH6
w+XUR14b4SEDP2jyhGAH/L8lv/n5PKkpIHebo4slDv4cZ/w4gL2z94rsxVMCXT/9N5erWxIt1zau
uxTcaMkgbObYp/87YgDIMsN3doVU635q1joxE/AL+Wz7fWZtVT+a8eKlfnfKIEtxVGqo3rfSZCmW
9Lifg9VWMmyjYi9z1lJLePDUcHu2X7GadKH887IMpRJ+mMpl2xgux7M0M3OjVq7XcexgOYXa16OF
IuhA2n7CUmKtW+XZptFT+7ONrY2Xf9GUr3s3pfr4/IydxjWuMzo5G4WsbG7PyxA8ZlUhxpAyQRW6
BRRDJGR834rGLEECX7a4AUjH7RdA8y48oS1tg/vjkfyV+/Mk8wpoFkP9VKDW8iq0HhmSgJnGVuoN
bEy8plcCmazLBKQTepy7mRMvVE1iNZDMQ0RINDeUqa2BJCrG+U9ohjxxcCn1VuuPhxG0YbcDysIU
7swJCz2nZhfXoiq93/36ABkcpYx3cscSuHxmwh272IKVWwRyRsq1s6CKeyl7oKMbNrqAKpseIVpK
azdnvzBWG0697MEaOku7jpEEMm9ZolIl64G2MHeK11YlXALhlPH/tlHlGUTQ1LmMheFWZt7of27W
2y31EjIjjhcbi8IxxjO2WWf2rp9GW1XjoWwlMRVNRksaf2CqprXxn0gqhkmDRebYSMKSuGXqfWrm
MlYjgAVEpFJSFDwHKX4kazvV5DwPW3/WKNPB/qUzks9OW7Or9MMpYaW5k6Tk0BuDin0dsgPb4WkB
sueqGg6k/2XNH+dVuIMNbqJCUpK4MbpN83g0QbcwbOAflsCeye0779BqI5QDAzEU/09gay0SH1al
MXO91Dazj6WqUCtZ7i2s1bpLcW3bbLHxOMEszELHpzSXhSzR4Pyr3egsx8WBNTBXYWIlAp8DW1Ut
OmWYZGydW+Iwu7Tt/T7E4mrMeWpjrYUgjn7akkj/ctyvy4McFipzGykmWtTkDYtlxIcIbSoAQntZ
YQ1bUAElTwLyuwWvUV3iwMYoB5QnlRRdWEv/8v6RTxfizyfuIwDR9nJx6KnrbBSpNAdBeFQOCUBe
gmSTlEZWg/KWVq/hUAPwsHSbLWvCB4pKEf+NyrR/QDpoj5sl/OlwxfUtnNhgKLm+9xPx5lQ/4Pfh
5kwJJiUGnxA61acndyKCAWNTDGiW/sxUzjYWPTIjwWgRW37xQe1CsnZmKffBsGF4wHGNkE+Icf5I
f/FWLc5YYx9Qf3W/TlNCW/H3xSxVC8m+/oU80FglCoPZNqXkTtwcaz9CZQwuLxlqF3m/ifEJ5ydR
I0kn/Y8tNAmdEcatSIhU6MArWvEpDx+dzhNTyqHc64amJtmLxHMDpOYkzHMj1khxvtBKNlHx/1gB
jZdyQ+vmT8duWAX1Q/JW5brtbOunic8oX0E3s9RYAtqMc4hl8K8RrgVn0kqVX/9KZexaONdm1vAO
hWXBNNSOJzubzt0iX9iiA2oMqAf1zzhgb4AZ2+a+cuMl0z/GEj2DQI1w0zjv2Pwl/dG18LOdyXSi
K148XoMW/JTZdpsxPt1uGqoEKkrenLm33tPWgTQHnqt5BU0ToKUT0QV/Fxh43vkCJYZjlZaFAKpy
HUNHgTjHLWgmxZzLmxFw7uYM0bh6C6KZD7bS0WFmAmajXcNehCEShEEst5czfYHOSy+OQ7N01Wum
SI1/tQ4yWpTfO155W0GbqeVX91/n6HDSw0YuYIHZCNdAAAYciOSTUv5trmvNmc76gSTS0pNSTHH9
UvxchSENKS7mmP5tOnZe0cEMjeX2I1fPdRoSsLHczJEN6oy2Yn8QDhyCrqlLDwHhoUN67UmhhWcv
6YuHtgJEdFbkkgM8iosIbJq+QHzgMnng0Try7yw2siUVL5yqVrm2Jxq2JTLO05UACtneEhX0ZH+a
GrtYB2siigcNEGEO6GmjQHbtv0Nibehqs//ZkSEjDJsBXDQCECKeuqmfhTUkPqmPvRh8S0nKsDpb
FvL8Ka99NVIopYGPeXY9dlrMbE6XHrFCPLgguI/BhKgsA++cmViLz6AFdJHJg893mSd6rhnZMleP
jSkSMHz5mTCBPVnkF1ErA9ckndztl0ZGsmQ8ytAehLgPWrDnoXzRevP/sy6NSY2pQ/CJ7s8vzwfd
r888mNSgEi8IUuztTttoGsRYfDBlYqUXCYEHrAVB1e9Pdd7WtCY/7Q/GGXLngUGBkLg5/jAlvkot
knMW5y62KISuT6M/47/ynPVWElYtfpPcOttNexlf/08Gb0UAQBle+sDhyZmqO3exQRMZL0gOe7gK
0BeYk7j1yGlAWfeYCjbmNTZRWZ4FLwNJbW42dEXbeNWminuHZuu+QDiZtiVJGECx41qK8zCLnctX
RvjP7gB6tRmwj/Pwies00b+lNEeBUAa/NiCTzCMpjMltteauTXL1SA01V/dDKfaxexns70DuWewh
4zAkS9QOv0ur0/dTWUu+aYL2XdX9XpYwbeohEYARG6qeqw4eAeEUUrEtKOAk0fHHk/ufumfhAuCU
f0C6p3N3Z8VR7Lan9bdB0W1551TdaQmKix7tBsqNDvLNXSebYFcY4aQIOOWY9z1tQyc8W3cBPGQq
AG9eIbUpzoNH1AnFU1tFQwPWvPxiDRqIMowoWQgDoEtkBO1CqocFYD30f4+TOdvUK5NG69f/RANO
AlwDx4jlHpxfehxNZdi5EO8ShNI27aE4q9LAM4iVx5jc3NdOT07z6OmjuoB2+XBoai8tP+ZoVEY2
OMFzezfa2jI0ZpartgC6FulsDDYpmJBf5HMe6LlPoNvtH50nGr1KPDneIiMmtK8gsvZ6Bo0L0mxk
az+w58tl2TgAKgG/6nxQxRCfKVnLIiQM2TrnHTGbW4ho/nkaIS4pZifV4MAs99ddOOBiNf7Zhp1C
hi/ixv3dbGk6cj4XeN3ls2StQoKjwHR7ZnRVkM+KUgxVqTp/K4QPcdXlsJT6DF6m7O6/bZUacWdp
EFBsNPJwY6dCxwYkrO+oDvaXbAoES+hwZ3Ex9eWpDEuEmxCW9DAtPg5rO8WMaJJeldcl9Ew8BgOo
qx1h+1xvSD9GTpgOiX1Sj61BIrgwyZQN3+q5O0rfvC2Dxuyae7S0Sl2U0UtWGTo8IHGxWo98O2AB
n52eZLpFxD9k96pWcqUNZGPgb3gW2NMUMYLRzCJiOrNL2MRrB7YlPVKmyho4JHBQS/rorYIHvLu3
qOzRrJMq2op69zvZJBnVjZ0DlH+p3AnKFV/qIHDskEf+ebnXdiIPMw9GFEFk/rehi6AiWfVyokrS
C5XhEoAZet7t7Iou8kVT/RF+gpvxrmcbtYG7fNhZIHWaidRIpPTQVceYfzggrV3z12TbUMVbeCP6
to9NYRt3BtttotrFNhLxnKy/SzEfrO0SMjgzJbEIgqLQVm3cj5CTn9FMKXHTRoNSPzahQ5CG8I0a
rLxQ6lxrtu5NZB7muqjjFswRhllo1sxwYxCjQAnLj0CftLRNMTsvaJO3bubgt3o9ybOUrqdD+QV+
00rgGGc05fDY81IhZfFc+zuvsx9bFdiiiP1XUs4mK0MFzbiFpET+rgWtoftpreWT7U2fm6h7vPLI
sjJvxs3gSWnj5ncfONmG9o4TgoNqPFG1PPgQkD0IRsWfBcuno7fpjCW+CLCztA22BurvgsSvPfo9
yfUQJlMAfoZwda25Jnz49w7DkA2SLSdrtbYiC0tN5yXoHE3iO4VAABh5O73s8m+jZhW1sVri2ZoP
Q2D5Sp7DtP7XzWeLkZIXlnxK5w3Phi3AaSOZ2esGLbVo2xNK3RHTvB6GPMZYjNJHO8fo+9UwbIGN
Za0j++3380vx5HMsmRMRv9/V4lOcIcE4MnP41Z2eejFv4iQcz24wSI/mbhXgMDFi06qsHKkGdBnH
ZPoyQVsZPkeDgZ8sAvPy7g87lQXTxjiaCppD8/f9+YgxbPC8yNpLANYPEGzyYVVFp6RG8lxg2T/t
6rYTdDTrgrIWtyBLke9cmvovZiEv7cZJfdteXtlS6rZ6N3Cnjlc4YYgRraFV2U7zaNdiEQ2v11aq
vKPUL4YWPscFO3Ys/6fvX5aTnEig/vluQegPfuEN8S1eVE2/YxJEkCCqKXTxSz+rIlmNWWY75ukc
hQjU3wv9b61EMu/C2k+FidoY1o9sCO4ZU8u6XC8T07TqXAiaezqK/+qE4fXYRkEBgWBq3W+5SwJ6
j+/T0F5fdUPieqPKqvDyJJVTmMKA//zVu8Ty6pU7TjfSj3KVSsqvBBv6b4d74+3H/yXL0Q6OPzuE
PSaYw4hQANDdNtk/8BNRxeS7hziRx/hnNjMaOzn7rKXvDqug0yhAxlv3bXApQwETbkLQIxIkUwO9
9gOq/eHqM3i2yuPJyJYCNk8cNA4eTzIP/+ERzf0y6jxsNc0I2YRuESaxHqTuDIod5uxOaGESh48F
pb8wNj0ngoOwCwxUofsj2UTMie4TRYVWulRNu36oAJdYzmZmtpG4OPvpUqLQ7vDb42Mx5iGjnBxv
dEujrD4ESlVNn0Qzhyh1RUmP4iUIvm/fHqhBzxZ1hpgCI+P77bRWWc4QYF6j5Y4lVERXPX46aTRe
smRYkYTm2fjDXx+OARgbKFP6ANyu1Nyz36ToYCmOjKWEeDMwf0rrTl86T8uhhdTk6c7tWBz1MbWS
4DJcOhMxPw5ZCV5y1ES1w1Curz/x+ygofeGMRSe5v1qtJMN23TeJU7neLFnMKJ31oKBkgo2tBupV
/tR0ecsyq1xAmp7iBB7AZUhSK42TErMW6+2nqdMROFAsrqIJulR+5culUAVX1RqX6dFq6Hqp9qXr
LxeLecttamWprQCImo3tzT/lzRA+PN0DNxlF+hOL3xprTWtw4oYuc8TUvXzyAbbSQL6M8hZxESc9
3wwAOiD5Rtxb7JWyYn8XeC6eWiFbfH55s1s7mUFTz7qRADe56uDUD0nKxbHZp4hkAY3iFuJ5NJCH
VmOeOGrSAOQL+9xEWovpiE34vVGf43Sohx3qQBI2d8cBHSAZ/VX6YHxDqpRFTOC8qp7tbeFXh/Vi
0XFTW6pvTsA7BHn3loqwXRRlT3YNcF4NzDzeMcYwv01OI5TulMWc282VPHvbbdwBhEQ1INCBIdPh
W070MPQ0vHGMisYZnAG/yZsHme5yIGZ9b8Subz2jzymMJWzfH468bJZC/D3+w7AUQfXB+hFs+M9I
PsCPFns9Ub3jVLQGb4Fc1X/wNMfGspL3ydMGaIaFVUGSrJPT0aEo76xerVTX2EvG27rwX9YOt0ZL
8wouPYXII4L9M1BLcapL8zLQwTS6Y/p3/q2bMAwjOUVfvfPLvTZjE4h25HhiaTdzm2O605vLTFie
mBM0aOl+gIaB2fxdUTch0zknPVviqXXK0cFcHdOgIHMg+x1EzQeg0o+twx11MYJx4h0CI7n1xwJ1
KXl07ZNVpNcYWROMK0KloO6MKfkd9Ksp6j9UlLJgB9SNJUsqGcvbrwlm6ykXUr4ABw4BasCGVi3R
yV1XXcN53nhOPTKdI14mwTWcektAp6726f4ECJKR2PJAu1gwRN6yJxM6n5FFwig3HJfMawpe0rg/
B/MnwFD37x6f3Y12lYCyrwc1FJuVjLKSRhzn7XB9JqWIQ5hoaozP56OLyHPf3g042Xt3kRIxDUYI
8/7WYslP+iapz1K5wV1da2qc8fODuB9YZ7BN76nMr2ZtYIN/rB5BY84Ym6wObEZvIo4iIxFoWVvO
XNLCftffxap14hBhTgm6GSzc4K17EZyQ/teiCRlUveM1eN4B+kH6QmLEldGTz9KW19GEy82qLKiI
R+OzNGs15DNqQt4ng2FvsNEMrLGJBOlrXJgcVdHHahzJuJNcXNfTz8x+puEtsMB86ZvNR8/ai9dV
EZfdI0gD9PBiyqbVrao5Sw0nm43LwPxrPJeiaVDBotAmtO5Vkq2UwaoeKY9qxDT+eqHjv+qpRcV7
l4KmmMnBPmq2NPto1UltAL3QhjXlCVIsVfSQQqFSQGI3E6VvHSxROoRSMIVgF+xmYmhK4ZzpELT6
NIAYgtNtM5S2J4bMta1rOtyXtt1cJO1YVzcqj2VroM1CFrJEw3xYf8ZPZVcvfgQlQS0/umkxlB5C
1b1nceFQoMnxBtzquGavRtwKma62T+y2ZhDGgY9gFzyu6KNE4h3aY/FLFvkOA5dM5TbsM75moVn/
OtIxDZ2vKeYsgU4X8RbOz/x3spdl9Uo3JOUTjQtitgc7Z6azJ9XRyrjjEV/oSBHan9bNPNM81qKc
/mUjhI1aiWvFa6J1t84MjsL1g9qehU9/TSRarROdMnmfh9DoXppfRlXgfEASVjH8I3PSPkJ1lUGH
lDu0uYpdK5TfJUj9VSuP+NEVfd48fwoEOucRCXhRki0Jt6iibg1PJy1Mku2u2Cg/5HvlAo8qF4R9
Mj5Xe9tmIAaF2pEtdOPODB3RelzhJU0IbM3TVhkUQdjSTfRaWy6H5APC9/F7pGwho68S9iSv8vDc
x/TxvfEj+xZjSXk5RKSYW+mNRgxKyv5VTVzRQEnMSQ0vPZl3s4jnu2VnQ4JlFJi8Q8lNlehQHfXk
8mt4+YOjxK+GQbW27z0HQkMquNAS2MM8hVFph/jqi3/5XBECBIBHsm5kQA97S+kW9Z4zqFfYTzr5
jrLP4xQruXHG2cecOC6QFe8IKHsf0hG7SPhJk/eF1+ZoXZvlxCFAuXwMFO/IIreh25nTUfXYCmwg
10+kABPBSobI/4VzolpF4NFcfQdllz8eDoQP6g2TMCx75o8xfY5xl/BpqgSr5xnufCxZazfWxA96
nEDz3WmZlVmdmL/79UoGfLKBH+pvlrx/tzFo6OmT911ivSJ458zTF6IcDo7cFk+DsW/YHRDxhbiP
cb7xUEmaemYHrg9bGqDtDcLppzqtOISccFfrZjv27+ikQ6sVMySWlO6OnHR6vgk6JoSq6E3QnWgw
/+ThQ2K8nmTS97Pt5uKjIGD41ZZVyeCKVpME/J38PqoFEevC+2Cdh+RUpK/y61csnVOkrBYJesE9
s4LxNnZSFK+W/sS1oUtf5/liwBimUpd64VucKY5fJXhJJ/MT8Nihra8CifdNLZl0ildhbYW3kCr0
+USAkzy3iJtoS6x16pcMsHcjO9kYOXAFd0HMq8wUCGH5g1RUpoXuQk5ahh5Zur6IHYvvhpk082oP
+XTS2cxDOKBgyk2nx8RTkI6INfOhPLKEipalIFL5sq7urNjyr1e6lRUomMntFeXkvCYg+vxi9p4z
g1Ki1nKU00PulpP9f+/JJQUck9LAg45gNXqz2FZtyfrPFurq7s+7m9jpb8LdWWPXbEnXkqUyb5rw
lpUHeoCEfD240+IPCyf+181doGdZY6EGxLUEuARUepY2NeaELPc5xaQBNmcVJFV75JuKP3VBRuOR
KUyaNUMHpCk5yHKsJI6LsBKgv0JwfpoLVMgcgkTudXArOFfdWu3RYqIS6X7M4co4v+J8RoK/RHvg
1IPcWlmLS2CDCRT0UFWZ2eRTEE5qDryRHDUk9ClLkg2IjXkXNE9881uAcRwufLH/7FHCLVtaDKgZ
SnxxwFucLtRAkJDnF7poL9I0LZp4BIrnP2e0pU5tg1TpnpQeX7Y9RChAyj+jgxsqsgnQbe8bampq
MS8nIGqQkt3ehgDJT14qooMwL7FFH0rh/BNCoQyvsYfShrBlkGu4KPm1Zu1adrv8nzXDrHEc/F5h
tx30tLZ/AxM16wV430wVZeiRV5yES+uBOLRQ83yvN36uyRd0TqjS3nx/HDmFpgeh//1S+wl4YCkL
oRLPGrag1NZYdv1am8pZFuk6m5LcXfmqha+so1Rtv5+Ez43K9SnP9g3S6lUqAaSH8HlRWJsVbSu2
d+QhS9e/KcxkKA3SgWNupfhmCiVZvYLaWoxDZyg1RFsD3l58j+8vlkYrFN3B1LN5SGy7Xd2aHhjs
c555XQnXpmHZbpjLJi6NQdhODg5talvJOIMMtpccHEIDk1r8DeXNka06AQq3bNUt+yxtSRo3gZO9
L3cOABlWVpcGAAj06rkcMhhjTuq/BX+REINfL0/c7aFPdKir8Pg2mbHemaF/Yi7bjrMG8Fqa8RfZ
MsgiN40wdgjg/1uihGetK5WFYcSUCZeUpwPVYakLRKxMKXgI45QQ6J7zJaIg7YcdUug/+Z/PPK9b
+Ih5zmlN9w81ymKEgJTrYP2PmWYjFk4uZNN2lpJDAEFFFv14UrEWSTKozFsVtEh9IGNjI0Q2JpDl
loGw4cNb1BMvE5M9f4bhb8gzMrQXQe1bPfwcBI53CVxbXS8bbtVvc5IleemfucsYyNxVVh91reXB
vxhKUvwTK4bSZtGKahw/f+HCIj5N1bLWSmZfdRghPSccT1LHiBkIvaMtPBfLkPHh2kCVFIXtN6CW
vDYUugLPOntz8IIQfQnnpo8UpHixUSwaPsCcQXQlbA83QK3I3utY8/RQJ2V8O4eZ4uXIRTwP6AmH
bxzrJeyFgkyl5t/rq61aVACeOGY7autsezPu8X1jjDhzihYI3iVLHYwJkAthg7nIS4rXHIrVv5TH
pm92gVpNwhc3QxnRVjehCcT8Sn0RvzLwZHYobaE9y2gHtfEVKYe2rDl8Z+ixJYkX76Y/TNtfEDcl
CrEJYNunW33ZzXXCCsLkPYFjZvgsAiDZge/KGL4NgWeOCkfS/XPYU8bLP3s+F+WLQwmzrD+jgsVG
DYYSoD9gZate/+uTHcNTHpWB5jGkZD6tKDxuO886aLria1gf4T0Znfwm0EqcUl9y9NT3pw20+WPL
MiPPor9hwWdCSKqSnOfLVtB19IEkvz3LmdWKjBYuhLVOwwCOL7p5q2WLjUgna36t+l90lBBlLkxq
GLA0v6s+UbHhfl4GI+nIyeT4691/v5TplPaMUpa7+YI2cK3N2qdLATv18Uu3xlRcCeQVs8LTJ1Y5
KCZWHYvblWq75aCxCWxs9OG6Ky+/gpFrgO8dUs2WHxvR9MuekDWEVtMVfDHIS0VEVKAJDqUMfkFd
gNmBWKJydrbNncBTsr0bulAz5w4nswte6RQq2oC9bfl5BaoP2B3w28+sk7Vu6SqY8/KOA4IUy9Tb
WHVg13Jl5lPgH18rSTA4gGJbUv0Y62WhQ42Fr6hwJofYeCEg8yTTpgJFnVD6D5QTHwy4OqNDX4Ki
m6AuDDXevv/Weyrk0AK2yUdHxmNWSKZqXx30KxI/n27dvnKcRWoH8sTLixSoafZ9X8xP8IjFC/w6
TgA+DbuurJaDCLd4hsQpqugueM1BPFt9Ai01bTKfV/40OOyw9SV7z0gU7Wwl3lHffhSXPVz2CGn/
dY4FalLsSlxonAIXi2hXTVNTr8CmnVaOX7FpFHbDfB3xCdOvLkhaun93OQs+TacCGNsPABNcYQhA
toWOFu7DqUshSyHWm3qHFLiGNkZ4JglF0dvJcsEg6G1gcg8czu60tdj6FQBI1kIE0RwtO/fYWDlc
eQ+jpzkG7X2Hc5rKOXudqHXTl5Ki5UuIiSrb0siW5+cSfY1PVUJHx6r9EQLj5QE6KrsSems3za9k
EJHvKf1kyEshwQTGbqP/dJze37qNx//pa1Lt91KC6x9H+JiRWZU8K2ROHngLI6w8XcvsAaGyT1yd
raYlhGYwAAqfCaA8oGzcSosUGBt4uVZU2lFESJOiSCsH9dFyKcJfChw/aj29Lpc1aoEnK5ugemoQ
ZXNkQDVLlFKGsa2q+F63hojpbMug474CWxDypQnh0J3mEMoAakM81poJgtIoR1idMkR8hQPQv6HV
/UEV85HHLcSlEOlFfGETQUn4gLvGCfhHp1jBj8P3K3Ok7tvsrRTHi7W+8bLh2kzTPU3mgZFEvfjL
FVSoX9X30SUx0XvtD9ZvPHMARI453eP6H+316UPdw8NS7milTrk2hAD0eHkPfSsyMMjLnSZWAGCG
iRqlsZXIuj+GS0Wsxm54P2ly5S/Xf6OtsmASmvuywUCfcP5yd+mnjADONlVNyqJkuQxj3gRJ0dqV
ZuwJx4B0F63NuvTJ/MsTYAa/OJibG6lrVzxHg9CrqmUBPGkh5308w1m7JNTkUpXJNPmFTWp5+Fl7
wIUl+bs9/E6q/Nr/AsFIznHkC2c0o6NsropOmUWwI71aeeuzqD3SkEUiKYf1Qi2nUwN3fORY1eG0
vYYzl5FzMdotgKJUfEBpC6wpThs6gl6ANyscGiIVMcR9GoisoTX62jg9CUdz8vQkcNZ3ACqy6sXY
OswTduHOtA5vOGrziquTK5JwRkc9cJ6Hvsgcfs+uKlWFG4b7Xx4WAVPyef1HbtvoSLLn8y3wwumN
SOuQL9YsDdJYndYB1dBcjE9vzfnUkn+qlHfb/SNMI6wFNQLHlkjvGlQG0SA9Q9X2kGkJUS+S+UnX
qYBY9Me5EDV0rJAwJYXW0ir7syKGBqcAQ4QmJA5mhltXalsFHSeoppVxqOyyI4X5Pf08/fpPakid
K1ZuOjoZX+w/QbwQqguP5u4Tqi2WLPxhybChnsjKFWIfuz6FCAeiW9o9oM1LDxOXXR5m3AQuD/p7
SsunqhrTtRHXMXQ5eNkeNFDD1Kmwmr/U6VzPWhmpksSkzS7pY0Y3DvH8UBGp+k0R2RmM3RfSY/Ty
QHzVhfMWlRJASKdRD4iyXxnE3c7jN+YL+8KuFAH7eeGB/4vT82KcteZKiO5g+A2v4Yf6E876SPga
9g7iosJb32Id5jYpdy42svLb438rilsDMNzfP6S+b5OqQaWscsUPjP62jFvTRG5mDANr4ISFyLQJ
J2PdSGaZSJcCUnm5gfv+OOoaWr0EIGm07qd2I1KAQt+ovBca0WB/YVoiXCgLG8KRpMfxL6WytPMk
xwO2yPFfaLh5fgds0mEfXvuQzCcWL5fUVZvIg8ZUPwGbCfm8zscgC67QvIfEpa0diZAP1v83CNP8
Kd1wyu5Y1xBR+jxsWderWkwpcfaiwIIa1zUVnwVZvNC4QxOSWe8zdgQYNAZomWeBE4mTjnL1KAHM
9SeRnHtQTvROqlaKWj4nWGSbib/R699zZxHwZ28bOFQ6cv4a29fPEIueTe8CvlB7lSY3fBwTTRCX
WbpoidwGSx9H8GQ5CBJw04sThPCw98nEVVY0DGmFe94Mc5+cTOcUm2LYiikzOs0Gi8wtuaFAlVPb
QroBUyGPnlKWYQ5jSYHoACC/qB2nClFOt7pDA3qlqoqBJzoDrK4kcIwFRj4o3mE9vxLoWOam7Gfk
fbEvGAH337WTP+UKEuTAjWlDnh1gL1+7B4AquolJDHiuCj3eCOPkoniahhpN/K3UNgmxetCUCTSM
HGt67PO5ieDlMRP8zwwG7ZwKNNwb/rg/wgdluX8ukGe46PUGOoFhN7cYsOxix+moqAAoAml7UBpf
RAtLThzuUdHVLyz0mYiLr9kjnIbtaSL8gJVkqKLL03EmJ2vPzXxK2DnUeKmmPnDwA6Y4atwzpe6w
556ESlfjPW9hALoCiBb3gnrsq0Ey1SNxV1c1ooVOMzH2MuqW18O1qK6/2t1uHCsUjZAmrhUjAMyv
6IzYFXC+oETOLRbkYbDcixn1dVl0D9LnbEIySM8s0iAmZ7MDypMXOWSvF0NscZlEGswyFYUJ+TO0
n+wt96QR9Roi8Bg0FDjUzWf/B1dgoiBmmkml9bc7mHgFMhembhMYZP1B94vcX5RHoprtkwA6n9UM
nNR3e7braLgrsi+ajRNkHH2XNNhn4ZOFDl7rBigNkaFxD2c7cRX33JVN4nomNbigtWBQoQrCFmyB
t35UlzSzAtlf6apCx8exV3F7ElfZAFpNyQItKmahUEugqNLID8bvJZtffx/OpTkFyDRotSGdvQEJ
zaymyglJ7h+Na8QQht5GN9iqoD5gXyrodJ0BFAiKbw9OzFnu+hyRUbvnhRTFUw98JEc/9xYub8ON
hBXCLZ8dpb+xoFG50UgljP6u2KFV24OCzvbK9Onu8P/Isxq1ZvKI2go7PIm9/VJg/LTRuFt9jxiZ
wKU6IVrQM9rlXoq7Hc9E7gzFFkN9NAjCo0Y7YdKWkCHNuyB287iNinVx1DbESt63RdeAkYEG34i4
Y1vOEt3u3T6ZU99VpiMLYXFohBaMj6+UXkh+v+pCZurKehamA1yUnlvqhRDldL1W5cWM7wUSvjOS
ZjcfIYRWXCj/BDm69GASp4//hY/nwSSd0y6JPWAmW3dKH+eMKAgJin3d2hNTGagCvafDrmC0tJ8T
8CeheG0vgKz6cp8DahHpXfXsKJyKKGRwg2iQQ0C9ljdevfivef1n/uTm2YKKHl6ATgUjGx5F063n
cB/zjFubnvtAG7Oa5AYlsPZ59z+bhQEEMzHYXgEhR3pzBwObnOCa5gojBYT37ooptYf2oqQaeS2W
1CJNMxqDoNNMm1hRpaN8Qim28UehOQOO6PF368urL/4K3ptcMaJSJ2fpMrL2ZPZdVDrFraTIxkqj
lhSwPikOhfL9FWVEVh/RvLrHktmRmr7GjWZKma2tmC+3hLcZjmKW7ZjPrb/Lnjq+R7RX6AFx6pFX
QirykerS/LQ71ZgNTwcgSeEfLypn/pgN0sn/JPbZEjMAkiRWGpIRzck1uDtH3fkf8C16kY0g0jyv
kaTGEtkYCbufkCdJ5bEmuCaaJs1iFZI+oPNI8/O2YvJ9nijNmPWsiHmhszxrhn7Man6EGGrjXCy5
lk9hzdB1nLf0DP48ZpNxWgpZMqsYCPXa1bYoi13gAu68Nf3e8wnuyMNhi9WbRTVKMwcHO9z761dA
UWkDjVCjqQEOtVH5SM5+RrS87ML91BNbe8hSu7XAamqj6oSoCjx5aV8x9+ZUMPrT2t/SvFuoZYxA
N3misDjZDS9VcD5vrqtivvZVBBBS8l2IzCARVMP5PnU90c5D5GKd5k1Smna/Zp7siw2sKQciuqSk
QyRPdTue8SuX4yVnKWdV7S6s/VIUAVFVbA2+afLVqV5HVOXZaqH0b4ytiw2AVRBQ5+tGXgV2iRKw
qkPDnuaIFQg/hRmrpptiwLTCSaafxqo2kyZ3skBraYZiM/kKy+WbnpEF1KinOLaQwFsrXg41Az8J
4vaKRiw8xz1pK5K1NZEiIV2r8DWTxxAwEbtuoNotV0qivGodU8fvh1GMZONrwLvOioqSBIIcwcdT
o85Dp7MLjRHSg0oT/tW1CoDjlasdK7m0RQsIfkO6zx7u1Q+SNhDSzTwyzdgHdgmospcObRFqgkx+
XoNh7WpjW7rp3JGPK/duOoJ1RoL0DnjbCB23mUQmGYkdbITaH4piByRWWZBnUwG5tthVgwRXmywf
WK5bebr+xIFpR1z1WUvulPPH7I89ih3nN4PXuAR7owyFmFRijunPuC/g+r6EL6avn8B8Ny87C0gK
U5b5+aSKE4cwzf0vOn4x4hicqMSJNlgcgt0rXb5hfqTBb0zvJSwQTW51PEaoPfpki1ss8vfjS6rL
Ul5Pi1FmdSuS58lYvCNLNhn/LG2EPhL5XyGfRIqO6r+EanfOsnngU4CR8jjQYbJJSo+uemnornpG
jSnHolSxjEAZqdEdeu2OZIDB1TkSGD6B02R8V5juv4sURu5+Bmyv0K72r7DXx3xdGsisTX4OEmHS
9rYyaPWhJQwVSn6Q7E0pMcauj7PuT4arkx3vgqebhCwrMc5HRgI+FySlGsjKl5lEOPlpjkZajKZX
Y1VZN/p6o9niTNITH48hwASs2zvKYhp2OxxkDxD3LJTNG75FBcQaoCI0Di0w8nViRIKdNbYn1p/v
bDZw/9lBNk70WmcpG/MQLtyB87juRZ8jNXwBXGlBfEYRHBnjpPuLF1B1ayUbtqv8dDThPH0AFCaH
eoxz0K+Pwrn42RlYqIzbFFQsjhgmlJuCC610L6gAEQ4P5sAHer67cFOk1jGs6s3QRKAOOwh7+fU/
6IzyTPaFmmPFKxz7vdOjA4Qzu1tNKdzZ5sQqbi+5YyOFObdzGUxPvA85h1Ql7d7g5iAd69J7+8O8
hoNdCvGqvaqxfPvim/CqVhBokjmDMUfIj54AR1y73BDvpBf1sqGLPBFeRH2b07izpFnJSOcixtmD
ZGVu572SzZICdUXaoxWe0PZ7X75Ec/YEIIuZJffN9KAAFEDSiJD/cFpX3CqeBnjHBIB8JQLuhoGT
BhTncksCzw0MJkV6unMNtyLi/iacgt8fuPN8ebiorXRS7+gq/1eEbVLbS4r6f6XbLhkL0HMlH3Ud
/bT0TyodNwKRUyWL1snPgAHgNcl7W6llpLB5erE9UWja+dnBxtH+4FhxPSe0efTUYAHZSHhtXmFD
5f6zdZ5QvkxPnfc/tlq4CffLTnjnHZR0c1FdNI77mP1vu71U5nLAvDHunVf0vim7urov0hQcI7//
xpT9VwQM+Jw67K9DB6AY2bzxWCwkktwdBbgETcJyi47iWwI2UOE3t8xiZxdxqPxhCgoXJyke8o5p
EO2f0K65x7T70eOuHNCSgQH8BhcRZMdSH6t3YYJEQ5XhT/Of+2XwiJpCE1lUippCATYVP1EUcMDC
/vttMtW0zZOceUsfpmfrEG1Z4TLmn2lLkK4nddYRWQD6S/10IJYwemr6CyTK+O2KspHPHEfT6Mnv
a10iXRRBkyYAMqGBMyyReFccl6aq0PW9LiTsZKq/CJUGB70OyHhRbITz33sXPID6q8N5MGJQ8jRx
ZgSgDzhKACCyCOXWIZbEDx0vHsip66XwMbM9pc7qcfT4trQHDpbMzDkrlW3FhWRfYRvpCaUVOeWE
s30RxAZ0jiDgQEO4zDu3J6rE+cEIe3sl6SdGD8tk0WEnADHym3U5OQ98uenNUztgn0WQKt2XgwRL
mfpZgN9sRyI1HKjv2DqpGZ6HLDCnfGh/En0wUaA6cVFhZHecfYl+d/IJUDnNGSgbUaiP4cyCwiK/
miW0DPuV9wDQ63atvtOtHRHKlieXUhtptkf2CxbzimWHa7+yNLD0MIyg6ZlLytw87gXCl+A/gYVE
9UxyzcBeCFiDZU04XmY/g+3Lvq5baRRzXhBhLpFe1s/RvSlvtBfyG++aIzIHPTeBE10GyiChparD
pCpIz37f7jr1tkom5UTNLTxjk1UVOaferKoPPBDqUYMFzIexuj/iPTdjRMXrPNGEA7S80rrBSUdy
TO75JiU4pwZDECUciuuH6vO0A/VvFC790SLEIVSClXA+Qe1q8kJ36xlZYq1Vn+Bh2Z3Jo4pJsEYL
ZsrV92negeZOiQSOIL7F6vJ8IzUTskNTXEIMsxlL7OSzmRyO0+PUWzmntftCgxtLKkexW3CijVBo
QWcynx9pUdxQVA0XvED94oo+vO/sNe82GsMPCoZdxsRH1E3fXmBINdyvVRqTbqqQ7ykTwoi/6z4/
yBmbOYkhIgt/3En5SbJO9QhV0HkvNJDi4NeLNjuKN7AChYl4he1WnLj2rMfCqo7sriWt48I71m3l
VCpGuvasggtfrU4s5b0kdVsXcp8ISl6/DRtkUwdloD7Grt6vpi74Pv53TYtec5HmwZJWxznTHOSx
8SziQAugAwESVGBfNOSeX+bOr0K7+VHG/ZZdxFV2QU7am0g7ITD1PRJMPn9QBP7r6NbnJef3ZYCd
aAiAMBowV2/4aHGKUGwKtTs9Z82AaFeoBT0xUOOuD7gt/1Jaenq6YEv3z/UvTn6e+JPWvd0gqwbi
MCvjGxDBqUdBsi3hSKli+S1kS0iz0Wnng5tUsU/CixQrU2+mdaurMozT5KVtoKwLki0UR99aKetj
YmPRZ5PR8wK3mbnG/Vvj73uOIMECiSVArpnVvzvXyyMQx2UsIire10nOnHLdKnqm4hpYqC92EM8s
ecChhAAd6mluqnduPrLc6C1wtGgwdPTpOdDMWU4ffsHr6JTSNbOWkmQNbTUO5thhWGLs6J5b98RG
Ne5+8Wd6rgW333RTedbDy8XXQB55jbOqnPkS8o1eSj0inCnG1CLbeDIrUNNMl7gCXYo2z8x6Q9hn
IkdbnsgEynAE9WIe93QFdmMzBh3mzQhSyUdbYYsMZtB3yl+U4KmvMmqM3VwBk/ArmcFCxEsMdRzN
9doc96SdJUoAehcqJq4/OVImyZck2aaFQNdg9DGhIjxwVZ4E7U9fnBNV+IXZVddChYJGnvJLDr2f
PyfDWcfrwWGsdS5HPt8x8uI7KYGTDl6vnG0imZArTNGbtQCS9emk9HLgLaQlBonJO4jnGEC9TYWS
/vm3Nbb2pJnGEos8H/oppZP5EN/sJPU9iLqQU7OAsdrNlLTCJewTyCvFMCmVQGat3eqTJCA7awjG
lpY7YWkiVzvYHI5F6RjR2xp26SFFksTpcOFC4VmbfbeRBNxgtMM+O0cy7LuOriySluPgnmYMxtU1
E0GXDW2wF03fErP88drNsh1KfS/+IXXq7+TrgFzr/saROGYFC8oX+4iJv8qR4KMVFiZwJ3U/NETc
z11EcnyQYahw9otbYoOV5djFfqXNNAPqQ1P8EYVmIuelrlzCujGCxTbT1TOTpLdMxz4c+O+jz9nE
iOemVS/og8nvrE+LkXYvW9N1T2ErkjSBM2QvHMjFFdyr/2I7h5jpbr3t+0djUw1juPyfX+ZStbAh
A8q+GAj9L0hWfTcGZxoPovcRB/Yen1QKN7o8o3+qFeemQ15B13OGIV/dByFng5hKTiuWdiPA5Mw9
/POaS0pNZNaHIa/FkeN11WHkdiNVw+BIE46VUGwy80inpaUWy2DP3t/W1r8uskh53LLLeOqkK2wq
cq0GRMPnKj5EWZRcbbmqi1Hl2rdSnFttbCygstrJe0o2rCKe3rbIOEFNK0OqLpM5jwt+niMAfiQi
3tXwXYWR0QqpplyjOdATn8WTyKTsLojSDik1auYAfr6h1YDfg3FdxC5fzdlhOIUlkQAx8O8vXJOd
5QEr78qJd281QedIXXyhUOKvIyqAp4blcLJQQwTriwflN/Bl2UII81SZ1jJVTUx4IaIZAGSIYJjG
uBgY8zoJ466frBgsah2SjmIg7H0XcznLS8G6tfFfdoLDPUa6pRjuM1uCbZLozWzmI52S7Zp+YvZy
E2dbViAef5MlSwe5q/uR6G1EIwXCpIMxjQJDsAq3u95p2kbYAgD1qkF4Q3qN+iBaY2X24pIY4lxJ
+UrSdnrpoBbpIfjhEmKZQPM/9pdCcWZFKTXOXVHo4OLhWJ8ao/GId0OrBe15YRl9zQE+ngbKzBBQ
rzSmPP1JMxl57+ouN9l3t6NyQIX1nyCV+qrwFFqNXmddtYyzi+sU+FAvJpo5I+AP5FUUROMgemvM
PZPfRNfw8Au0d4A+6wP3lEycoS9pWPL6I8MAaVuZ7b0wSc/1H8VfiQRjg0/8103kUx0BH9h0KgLc
PwYa2Vf0dofnuHjCfdLY2d5F6rh0b+0zYlWyGbSM8o8lFKuXpD5cWxTZgKB9S5dOa05ZCs2og5Jv
wD40tu+7lI6r10DoIRmoXha2xBNQtYfkQh6iqLLtKIFJxaLcgW1jLtOQKr66hnpIklJ3eGIyuA6Y
aoVd2G1IY49eenjbQLbxzgRAMmXc0LqaCSjr2WU7dlJbixH/hSZVQXiM/PViIHM1kHCMF6CPL6JO
4i0QhMP1hA3h75Kfakz3WZz0NC4a+i2JIaOTTXAjqF2Rw3RGQRnRTUlCqaI7ITcAdGYcAKQICk/K
ptM5s+OOq3mYfRsy568/OSGXovkONyPC7IJzLaSBuA5UJxj5F8RMWoiN7qgF/V8ySmIKybYFGOo4
QXqjF1lw0aCwSBbiauDECiWJWc4k15fXLLZ4CH/z7kTXOh992KzlHdl0YaA9uFkZHI3dcZmAwb4z
GPJVTArdonv+Ra05vVDKbUK++0IhcMbvr7WCOvClN8QOJ79BeFKETC+mnlsqM0fLhh0bzzDP0DYE
kUhqnNa2DYJl5gCyCsLq2rtxHr+/fYs4QIL7Z9DHUS0fps1NxeflMAHY/bXXA+Lcw0fdgbRSAC+k
U+9f7lWFvGl3cq2EEC04DpPeFnSFI6pZ9Ms0KStbyrthPE9fbcdUrOMzQSu8XvbQukcr1SEW0aNq
XRl1r2P6+0e3kG1XTx9MUa5qRCyD6PqCmjY/6wWiGHBj691anJ1Ku8xiEyAhCbUP6CF6nMAsv73B
NeHQpch5Vs8ZLEQwIAruBI94OVfh8C8oBiqq4OXo4XjL8r7t0bS6Gd2vyWUMiv6/6dpYtan2rg/n
U+xYLqDAkhlMIQgRWqgE6KaW7wqg1JTgok6i0uXHdtBjQKHstnaQwJdxEBLJMaMXWQhEqicw5GVO
UeP6GigaWbZF9dRl5pMOV972RotdWdZoW0d2z6Bt+8jC/ufSAWhAVmscfBdppEsbHECXIg9fjzj7
524xNNdodF7jwLb47cndouzQYovy4LFpzUHqE7H8a0QKkDbqYgZzqhv8mGZ8lmMC0JBwHPtb3vwo
7fWRu3AXk6iVvKNggDZDLD9tHaxncqwkeDG7cDOON2Koe+oLHR8YJnOwfyUwc1GJ+lpvel+RKRht
wm2GfjFuppJUR7IRpJ9n7k5TKGcQet9BLFvCpUIOrfkzwSLdKTuHBCNrx9Z0O7DmaDYUn7D7HKbZ
h9tbSToxgKVJmQkuJlOm2HewK4dfI6kUK0T21yS8jrwQIik6M+l9K15DjtQic/Ta4ES+9mD2TJVM
41dSK2oeQSH3qjhDl+7hvY2jTO3dmaCUAzr5owt0avqPwBDZ3/yJlQCaBKNesJnO77WT/S7UFwri
NG5JTP8/+WkIgq3hKMQUqC6SU54Lt4uur6flO76zVZr4DRTYdw7CimuFOPZTiAVoZ5uVPQSTtMRh
CnLKLbaDM41UFExFfrT3s4cpNMAzM4DPHtTTsMMilnA6U4zKtwrzGxc703MWj+gY73fM0BIelCwt
JA6aRXxiFKisI3q0hREtXb6sNRR/FXw3qC8wuV7VWoAsqkT3PNqV91fSn9yIzibW8ejkGfNDTp0y
juIV3woeamIngXVMhanJHdDMEEjy+oPo5EkptDOPJMeDov/zSHyoZaIoY6T7fImG/QrxJqbSMIvn
JMQRr+jS6D6nfzFZT+pp/6TNwkxNy1som9nGNdFeMO5AYBBcOqs1jjn3vBIy5cQfYAsZfkiYmDG2
0/r9tl2Ppd+zWefwA8ELfhkOThlIizhGMaFrl+oqYzZeeSCfdXDnjESSF+dQHP30QDJEr5du1D25
2naTDCkOpnqhpdsC5sxXBPzckkL8NVQfz/Xm+ITWOFQXmHQesT0t10ppDGCGymE/ywdSa/BZfSXf
/NOVaJXO3Pq6Om2e2+haRMhGf8Ua4WujIMiwPBuqQQsD8d7cSD/bHcJkI/RIfTwN/5WXdLBuOxnW
UklFZ42aH+GUJiS5IwWGCwFkNEuVmJRqVyZa8yF4t+D/pkwOmWB8D/LkUky+UnJNr28mKuSN+Ygd
xH4vtOA8MBESfN32Hkg1WaiAaOKZiUfOlCon8biXPduSS2JbNHR5DUixfGd2i1VI8fjI2V1aUd98
m5Hy5XuhtxSprGdwp2zWeySrUoenTXNw2D3xEDGRfDObTBd8RCYvRdllYiww35/F1Oim9+FjzSK6
LmdmAd7tGinTfTZcoeqioG/YfsZwVZW8KxMVdllCU0zDOLljuVzytDCrFYcbtMa9xKc8b3PCp6NT
kab5Oq/I3RriswQ9gxqLqAVCLSht4xoStADvLsDpsBFz6OPb6mPyYVUiblsx35McCwLyfQNEcKMm
j4eHppzkfNgwskLBS+J75q8rSe6LTM9cwoqeJTwmkvFESVUDI0BypJB4YSDAnQQs0sp8NhW6Jrxx
ap5J8huIN8teDtO3SldDxN+RCLtJj0FRJdNaD6XazTfeJA8DWpMMw6oJIevGipe1crmwqHjmPagP
f2uiVIL1HtV9EhRf9WHnpEuNj6k/rWFmBr7HBS0zh/WjlgsUViPq4W6WBHRY8dHsNswkvAV+U4Fp
BNG1pbGNPCqnN3eRD7UyeYVVp+9PonCbHF3h9eun4IHH64GsSqaItN2iqNahyLfTOqb29KgaBQpB
JaCcDJ81WoUrclEp2IxsiqKcd23ZeyWWbR/Qs3KvdQwtKVrxVhikNJEDDUw/jdjM/wud89q55AM8
Eb51TiAZKy3D3i2g3qFaDJnnrwOQVTaJ6UVSoBzCiM663/3jXmtVfnjmjh2ox1w9uX4zAmDu4Yqb
5/1Tc0rJ70wd3mbgNWyyI6ntkD2Iibu66pwolYHePtQ67BCNzXtwOadZTcyXsqVDDA5YYJZ/DUof
68EZsnfBX0ex9Xdu6mbGmh51SF/phWB3+9AAek3JGnc6kGEPK4g7xp8jzIkfRrAqRFuA7Fz23WyP
aZ4KYBrJ7SC22onapSFA2d1trGvnzr9kEmMr8r/czj3GI+nE47yt6SEhZprKgQIxE+e7ZX3ct4DO
7FtgjwSb0cU8NF2k7Lnckiiv38wiWhL8xXOGGPWZp7jS4NoVDJT5ui6ElUw28kL2Y5pS9gDQS80o
/2vI81rhi25E+s61ZZxI6YK+l6JBzUIJHh0f2RJYEXMDKDL2rl0/0RJMp4h04Cjie0Vi6Dxh6ZWn
QncInMih5clfmptBNYvTH6R/hLGLFy3Q9ubmI4K+Cz8JjQmv4ipqvTKKXfTqW8BrlWuGqt7+MOr0
+NSnEEYU4YtjRVrSimoUdIVSx6+ml5xRbXpiDRLM3FGEzDuZb5khM2s0pnBhrETvVXjDBjJxlWRG
yxNOphPYrbkFdT04f2EBcwbQtkecM5ebG7z7c4FQFd5E6h4UmwZ8rK74LkiAXpseD+W6eezZ1nKb
DoHIEXrKfaV/5Npg12o4xxnetOTSO/zUhPGK88VmGW4zNOYbAO/TI2bxYwqAwgDDWASk8MROqs04
JMpmkpSzQbZVEWL9+wYifOOcammJVg4AIXnVHtVUe6dAcBm1SsjmbXgWwCNE1KqsKPN9etvxeEpc
rhcbK/T83W71Q6BFwk/mcDAQdGi5KW5mR4rAthmpj07HRGNJQ+lpQprAWaB0WF8nYbO1es7HiV/y
IryNbbmd29YgVNafPv9yFaHVy01VTTbLWR7esmrXnRYWrlr/zDucegAh/c898o6dRcK3SQ87IaKj
2J4ANojj0/S/O8ScpbSonWf1/V53r1EV93u+HL330Lh7nuXN4QRIHGJJNASBlg+gNWZI67FkmeyM
oGAmoaW5HTqSY4rVzMQZaKwE4JMRVqtEhD12J/NLQ7fWHfKp6HOsIFJgmpdNlxv2sgcBmNLzBlt9
EUpqdRerfx2jvezXUgr8/Bg0lzMCytf6DkFwboTA4d2Cukn28WpAFHoZKvvxevlH27x4hXal42ZP
uz0o9p2ZuCUtc1dPxIzGC38F9FhvuySMhAnRTI/PuWGlhJOx+uqrETUp5Pquf5eInYXEX1rbFZ2o
JOdVBAHsZT/8/ZWNBRvx/mn8mNxBikjLsN5EjxurUdFsLM5/O0DeBILKoTx5U9wBQz6Dw7TQp89I
lsiU3olyHYqAmZVc6456xIIkr7M0KsAXVY+1mriWSQQpL5XbSxwV+I/FodNQBP2e/LfdkhZUMgvu
WbGh7rVWsMsH/vpI/ViHewrqinKVKCM5V246s+xcwUWc6qI1l4hD15rsCHKB2YOPo+xz8g4r3jg4
/xls2J4DDG2F578oel9hGWMkOkMC6DvbejKDRL6kCryPqoiyqTP43xcg8id/mPxNeP+TksQnSHxT
XJ+0E1CcmQk+kX+BP0j2ZNTHJt+aHCrc784cElJCYwJOlXMAz1GPmJkOzlUq7YHdfaMUegLkIbgk
W4Dc/4XW8LAU9Vwv3CinP1uJyiruluudnPHPr3Dt5PUfB1Ce2H8bwc6exZFsWoKjon1wXLPWxQ4c
mscBLh8kjwYL6myYko6DHhwWTqXYeZ7uoZSwOunk3eRu0Fx0Byd+UTN7lKKBeFou5ytsmyYIvjgW
dgtVZ4K1XdPHgrPzQKKN+rjrgd4b7E2/i917JfoLb/ch/MXq1MereuEPgRr9pPi6y37iTDOgNleq
fyqLFHNASEA1PpaFD4fyDjQ5u+cQvu8I4HuHiSCsWlji0kjGVOcs7Eg8Ln5gWLf0oVqvdt7tOcQH
fZTP5+4QMHMRQfRov30mrub7hHZUpV4kAAX8u8LKdro9VLASRkpQum/NvDG1rDgrPBE/FWQ2WT/w
nEAKFWrI3k/o8JeRQUfTN9IxzZLp+lCC2CJYYBCCGEiWlIQKsdiDRIslzZpaqIt93Asp7TOQNJdl
MKUXwtCrhE54AHT1ZZ4Y2g6Fx5CpuMgflwdNe8UVE2KO14yF0TO0zxhJXnpc05CLNBg8u70UkfHG
S0fpxfS0NbheHV/XkxRq7RWvFU7+lTJO+9hCJ0VD5TamJOXO1TK+mRNN9QZVQLbfO8p/Tx4deeDS
EKaOi653fX5onE+E81xrKcOWV0CnJB0P9SmrLdMJ4WxsxEXxzS7pEo/580EDrpGEUM6rHddRsc+Y
+tqCFZ9BkO56ZY7eAVJTok/X2pbGSofYsTPYsOsVSZNKOJwG4BHZAGfTWyS1Jx96hN1iyxk2JCJT
I/8ZuQpAO5wGkYgowwlTt4uXm2PdOW5MVnQ2WunDi70Be9uzP/lt6uVJMUNr5ty0wudtcE8YZ5eT
zSBXp9BZK/fbDWfHVTYWuiBUf7OxvD1epTI+Ddp5gUJshPLB97fExW7LVfo7+1oMJO8Qvz1t6rtI
ZSaVM6n1b+s6oY99X7pqeinZ7fhnY7tZnxBKtAeFHvzGjqdUB4qmZHdejwc3dSunPaj9RXh4Ie+h
Hm/rkI4HTo6Hyyr8Z4PcWnBRHQfu2/TuDpxGFvzOeqTA+g4d/QpBgRvkf0ViXSUt5bHNuY63Xi6K
35pC2sYNcAMSKOY8y2zWPPoc1cPE5r4XY+ztpYBVPhBrue0K1jkLj8qD+4FyQg9np+Q0H32Uetjl
cI+G/g6euttkKmF89OOZ1yNCMsLQeWSyH97MmoXjxtcEJdyeMADJK9JeK/Vz3h+dbzwMQdCaBU9t
XGG80kCIeLYusGlKfzYLI/WSuT9RNbRsVXC3dGarwUpVK8lT6KfaSY2Efwr2EHc4Nwl0o2cxjeCV
V/4LKj7B06KmSAFkCfMqwqkuNvJh1yGX696pK3WyEWfj10VsyO4Zfmg1f33XmpWMGw0ELGj70a8e
tk9vr37KF4hwu8ZmRtkfly3Xy/yoP31vFE8UuS4cd4dRxYOPeeRPQQ66maqnwhnkr9fB2kkM1BYB
/tKg7xeVW1b6blKqc5cR2+2MUXn5LAC8SLFkLXqL6UsfGxchB6YFKMWYZw6PUfUWf8PHY3LCLvQr
qmXF97k1hhSsr+1R/xsZis+3uPO6W5KPPAq5zaxrOHrsCF88vYMjocssmoDvufGEJToGGe6NVNyO
kYMjklwyMai3aLY7F3xPKRyA8Sk77c0g9DYY8vUSe7CD0iCtumO4JhSFW8BS9mzdnDsFgyQi3gga
wFS4Wrj7AGalU7Bet0izAvWyrRs1SbCfTRuid+giJoiCQKb4GeByntayNcVYmgA8HsVXRlfDmeWH
yWTJ+LxHdRqZlpCfQI9rIOFtM/xRrkUo+9PExaAMD/ZTpTxL7qbPWVrey/1TfCg9ViDZHw6jAbqs
fv/k8GdY93yW+dZBfsmCIYwfBQo+5wKIPLq1NjYEAW1NPUjHoY6N/B5HxOwiptfcjq1N81dgUMJD
gZG8qiutj0RlEblA4V42ZoUFW+ihfaYaL8IU1rpV/I1zMNxaMntTqB4rQlHdlk2h9gTIrUyWzQlZ
c9jvwmHD5npva7fTOL/iQG4uh1l6oXEypZBkEpPsMJKJ9oEskp1bEP7iiWoiAimLdaja8mPFtwnq
xUgkDYqvajfQ/slGEb2fqS+GdKEB1Dzk7zuVgdftG4IBCsgybb0JIryMfpplr11T1VN/IcNMIkQf
vfKw4Zcz0Q3YedgCrfF4RdbTY0zzboxUiHApq9EA0rAqGpFCdF9fGg0BqoRGO6jQ5OjKPMHGXZJy
/WPDSCa0l1+wFVBwRmuiaAhmf2a++1FiA5BXGzKpxPkrV6VrH7xKbTI6nim2Oz+BHTvdKrdm7MTl
R42uBSoxUWu9k/0PLsaJKauQDqOB7kuLN8+Y17Nfz0lbWzAQ1WiWorDE4ZYuS3eE+akrcgCt2s1B
SENAANFrYNR9Z8esOWXuiv406c1Qgrl6wPLOQxXTmhunsa6NcniCx6T+CI1RicoLP/v46eFXNJ4R
f2wUljF9RFebYXPApsAmpMPdEFdWf1AjBrjEl55dHi5+KbqyPtfA3ZE9cxJDoshGp0Dxm6vKpOlW
vPBcZGrlb1QnuaYxLHm6MfI0dMbO0SSxyTA/i8n9MdgyPyOjtQj+mJOKJAALPX+d0e5VNs6xEx/g
oXP3M1olgaYSpipkfTPFg7cit8N7Y1GNHnw5s9X2r/i7FFQ9WEmnIDBrgf9G0y0HaW7EYws5dJd/
rnx8OFS+uRcWmyytOkDrpPPFcbhIBbZxwja/Ogzg4CYY5hVxBcnxERvOmsnuC1SibtydxtDZb8AC
d4aT8gdOqRNKd6E/fC3VDKyU14r6EdBaV6e7L4PgIJLxaDOvkiut0V9hGyXtQB8Tae2oxoYBso1q
GIk2u3m/m8OCyR/+LT/K5xrTqbziNHLgQJ03XPu7EMu5Vk4n8zgvBjvpo0O4yQV+1tkrZUtovFba
ybqLCfKyAneEO0dYip9ifpmjRJbzrQtr2U7RjwJ4cYMgaO7rhVrO1dNe49HTZvyE+K6UmUhFxTB1
M5ggcHtPJZ6uFv1yNhENbPkeEKUKpkrb6krVYKvOlJ965TQWh5tqqvsyHOUUzet8tUWR4OW5RtlJ
PktBz3KEfxbm13bNdtdzIb15ROR0iUCo+1NBD6or9RjLc2+M2dbYcQg5E0WV5hwXhnGDxluioYwg
T6l60LWxv41+l16EtZj0zkwkSKI2jgkdbB/F3+iy75RkkMv3/qTH74MpECi2l6oheh8apza2gUgy
T/hfVK9I2IYSikIkIct7qP3OzKCUP6f2GJTQgEPb4KPMVlz+opcB6MexZ4UAh2TKru9gHac9LLdv
dXajVDEVRkzZy4q/+If2hAqsc6Qp0LF2vOOhWPcyTT5eaJ2kfNKDovNUrTen7feG0k07H6QOIHUB
rVhIxbVZzdbp9V7x3HyOK1Ll9gFr7rBrT9FwyYi0Pj1cZAcHxaNyRBcvws2A30t2xNkF8gbG+2zR
Fsv8iyM/90AUVHUdKer/gqnLAJOlmX+2xESBz2J0wfBbOhZGyk1NGR1VStwmpVHMDOsK+STTvMhM
2bLC4c3Q/i19DBzH4jq9jXfpVqH5oN9hOf3fMYpgyTHq7ZZ066x6W7Y875WNckUIyYUuHr8IMO7O
XJD6jKRFLO3D4+hh38GYlQ2LTGZQaoG8VO7znpTJ5vnKE1yB+QS3gc96UbSQ6s5hC99KuYjZHnQ6
hsvO+YP6hASwC1+Ba8Iaj8OucAm8KEIz7Rtny8nH8+cwsd8rtK+Cq0xJaNyGbjFzFlR+ysQpHZxS
GZDyDDRlEcECQHdyseO2DyYKtUcToU/boGxzLr1xNte2m34r/31Y+/epntqtC8OLAiHc2QbktLFf
gV9MKC8i7KGKYYz+cD9xJD73QUeMDqtnPwPL3maPi5l+9gFa+9V9/z1RzHn/CXiWQNiHMQcvV4HQ
3FKMZ2sfpy7Tp3MH09/XKTjRXUd53q4Hm9yL7R9pGWgZpYUYwk1ey79cRY9SXYlCfKtrjKelyF1R
dVGtWRtCMB3jD40cjGNILgoQUwf+9pdwZag1rDgcEQUCRuIE+9annC/2F2qMuNbgO9ATSnh4GDw/
Q7VqdUlBQmpx7Ysvqfl7ZgkX7dD3soKDigRUXE4Im5LtfgAYijTmKXVXW+D1OofDLNVD5lh6cbJx
lwv6+ptfneNL7vyfmb4HW8ZFu7/Kwq4vlI79nQw5Im6J2bCCF4GMFoyvUtypNZgLQaJnHQ3fCU7j
J/hiQ/STf2XLaM5Abukhs1njrqyRSNphqjoMlZNXKzmfhQSl0TGoy5KzlaYU1Rd9CvFdoGkaJjxc
Tapdj3YKOBnVJjlSOc4esBFIzFzJbNQcD3hDGj8VVafVomZ7/4Ro08E74jKjigvzcigNz09BqIvd
nyp6rrJfT/nK9E08IBVk9MkxjnEZoMoEsn9oAtD39Oyo5SQaSSxr1vWuW9SeRzGD9bELdwaAAI0Z
L4UhcT/fMPGpA1bbM5IBemfB5UFgWo4SyvBUa462QedNnbKyZjh6yW4cEnYML2G/DSpgDvgdL1EL
bt0LVcHUJFHGsczyRSDrETTljJIWiU2wdQqBv29uX2VHwBhbVxUYOk+2hubTW1bDJo8YaACY6fZe
DoP1XiDOVYWN+A2arDfKJrtflb4B4buRPfHUUnZrdHLsfVkFCkKuhZqKLjdo1mYPcxGBVioGxoh4
oPmVHpyUqvmtuvvgrZOMpU8R42GxX8l8AzhzW8y+PFSypTA+G+Dvwcz/8OjgNR7jTBjPKruJxnaf
bwjhlC05q6ap7KlMj0StC5Jg0GG/9xrETsizmk5E2Bj81wh2zNPmVSLOzmuQxkMC55/ejehvVSKe
vFdnonTc7vjWArdl8yHWVIa45vy+YCvSjsIKdHRU4t8b2PSlc/3ipR++E2oaoEPP14ciLBkTTw2D
O3Nav0bdwd05Pn5w8w6+YpWMvWlOy6Cx357iQWPLtI6rI2MIn1JucAIxQYw1zbvAQbNHZLVQhe7y
gE1n66FQyJwCwj0935+a/x932DUtAWEW5qxv7Q+APCNrxUQGitgdEBq3/A5neaMk8zepsyRkggAP
2tSunuKanhLIdDJTM37N+hFd/y5UnXeekU80Okv0lQLB04yHVvty7TObpVRYbHiPsPvNKeHpOWTZ
k85ZwvD5oU33cgTrPMWv9Z9ti52aRDiBsJgj+AoAwrpFE6T0xFRoFzyOsxkiwCht2zDHj1A8c4Qg
CAzMR5keu049mcHAhWOzt3N4JgUnRK3ajhJ+0Q8pyN2DPFzEfE4AHqNXRmzwmHOxOqN/SN/i2i4k
kka+mvCgxiAWZ1+CTPsv274fdixwyiEhWJMIAI3DbDWCSsAv7YVuw3HBjDkBRUljUpGqQGxQk3f/
Kf9pT7TMzyKeQKU8DtIrZFHla1yku11UjaXedCYT1Apbx1Dn7fdbVNesNCsABf49OIhYIysQkz66
Xr00f0/cXh98psNyOVQUIGaIY0u0+t8TlRO6I/3kvRA4ynJ4fVrZMqBWFWSd23Dq+OyFI9rFDyEU
f0JQ8l+srOBDO240TJn1c2nmhP4/8/wNqKN5f4EYScuKM52AA1I1KIJlh7WJD7D/+t5C3WdSEJu+
qjdZ8F+xuea5rvccsVbo/MinsrWd6RMM544MUIZjoQ1tj6TwGKDlYaHTIOhjZ4uh50kFMTahaL/E
0X480w0KVEgnoKXAsUTCK5cltdcAcJf/CUPrtFDSwBW5yO2pa4PhqwLkAPb9vvH4LHyVRWIjdIh/
tWnFrAZTPLWEipuQJz00JTeFfRq3UhtJBmyQVy5XxxVZHBuvbGbpkZSiyFaC/NyX8mNrcyFAQy8+
TiR5BQNydXDWdVbzOTsY13gUtBmn4ltJlso89H+vNibmeKo7YCvRXYBpH1J7Fln/iRWOBMiQ/1Jz
0pcp05nwpeNCL9dbZINgOuxs1IvNf9HbHS/BQDERJucabNitpwyrBc/GX/AoEyrcHvJZnpRMFfX5
lMbYieij9HNN0svOdIgQuCjuUPBCd2FQVlpDMk+jJkhHFakED/CSwbh8wtI7Uj/b83aLNWNL7U3v
xr877m85kuelk3ois0NqiwzP1gPnjx3nuNx1fE/BzFs/oERBL5ys7rFMNyJFLiDNAVzeHVnCBRbp
saR2vvfm79GidC1WL/Yas0Oz6cjcZLN1cpyYwDNI2VFFzIJipLsZLlXTqE1Wy98i50BhCmZ5p+GR
z9QpmxcsCzNhaBwXGRIu2mO8uI5Xl/GXxrayCo1zpHlpESbYkNkfjeS+kH+DUk6yUPjxJunR4nxQ
RwCIW291RIftlPWx5q1RE1p0Ab/lgj8ysXa44NNnBdnHc8iH8xSQVkYhH9n9aook57aGqPChtjvl
M/85H6lfFFlREdACEdDRk72YbBlmU/WvuYErGpVEDz35seCsxGk+/j8TyEtXTtI8ql0Q0H2qlIUd
u0YYRpZ6/+fbSlUXuHnEvRay5k77XhMk4MHbG4OtLLHS9Y0zPhfxCqVf97vrnI2MOUDh2o9wKX+1
/s4itrC3N38K5XhIlh7U2ALZRyBfPftNV2P+oOl71EAsK/VlFq3jc7rpUZsE8mvZj1+z1L7B8VPT
T4XjJaU59E3Mo6o2MHbevyk12ZHdoOhmBK4fM7rC5rlvjZJR/nz86em8cb0Q6Has0VVCB4ROUZXi
77FnYiqgZ5jv+0i3dC9Ougm7MZ/X7OX6OlBoeBCkAL4/riVQ/GIgdVcC1z1eY4VNSGIijnk5+718
eddPlRRuxxOqDDGRLmV317uvCzfpVQtLzsIMnAosCr+1nvvJ0w27uTUPFf1wapjEkN+gWexlXK+a
VXnMJrG/Ri6O7d3uucfMHElagNtKysQ7oTgzvExeM8uY7vs6GsU30+wZBYyBopS3ZWI13xq7Et9z
mG/8VQ2jHym1Vukcndn50W0hAIhHeUyJkmZHJXoPSAbPapFThGCLl/7R89HzW3bSqyhzS+r+CpGW
iB+Kf/lJ0Y8ux6mIc7yV6asogKIBo/CxRoSprUKJ15kjXGNGy0mBuyO+FRhfdSbRvAb7W3yoZXMA
kuzjTIp+IKBSXuLRRXQglsTnyHeDHdvIQks+fXlxw0PIi6qghGgXj7Sys72JTQIInOUcT147MyLj
zlKA8f+CCyDRFkDMRIo4BXABuqf5hR8bHLfZvvL6GS6CHPndxXiAkTAphSjI8b7+Ab7SgHta4sT7
nPMOkyHbpFT+SBiO9bK7RLA335ZJwKdyQ8FmZ/hIAxEdAWmvP7Q0FzbpkYz3E1yf9o3S8bzBFXCv
MbDmLLxUduL1uNSXOUcc8YR2HHPQdbTL7nxTY7CfKPLsZq9Ttt98qTIURwTlpLFlTnLQjOPqbCoc
6Ha1ojUpQH7UCwSlPGu+7zpLdAKwUls8Az2h9kEO77dZvfjlZpIslkEyk6PePz9IXUaY06gc28Jz
buq/1i2A3gUNWqPgvrYNX0oUu2/UgDN3eIH+FCzxIcAF0xnfSRin0YlehUDpBKJTeVXDvbRP93Ut
tiOUjbGzfcp5hv1iMv7QHgn3B2LTo6A3AcjX8N8+nwHTSmOj9s3qma8NQqXnGNSTtqIE0wNzCbC6
YeIOeBBsYXnxWBa4rSZuEmRwisLmlEI68n2ZGHbsC8Zk0V7rX7T2CwwdNrQYe5fp1H2yN4b+4fKh
kcsBus7V4wwkA5mMJMzsXkCde59k2dG8D8CVdwZVXaMskLh17g6ef8eMh1A2C4WqVrL2XvJqUTfr
woVtAbWAPvDInQQ1EcyXLY6GtfC/qvqq9B85JriM8EDjWLdqEQpIcnWZBmd5BPXaZqT3peo2E5+K
nAjxDdK2bnZ+o7R0fqO8Kvx8BL2mrJxmN8MCsS+4pnUAg2p6puBpZyQj3xJa7DJq4552oC2Px1hz
clFLnsMIRWpDwtR203vZXPcqOCVhrk+UwYDA/UEfY9EYtgHNZ8wTYamxPGD8pEiIdOAjWMjE/A/L
mHOpD2hNz86L4o50MI4MzEkwBxaXtz3D+9jxRA6JILn0VfeYo11WQciQ3+sauH0K4iPk2RUpVlFU
K+xNs8Rmw625fi6tFFDig1hDrax+fX7kFvZeq0FgvsR5jo9dtMPvu3WbqGCQ3mUGoltaJHFN8RmZ
iwWJptYlXMSLxBaPY4raYL7LWmz1CPLg+f+l+nuH680uzAw8bcDv6F35DvDgdkUmDRiOrQoWGYPs
N51sGcwcvZtmP9tgwYD7Oqh11NyAN7ODCIsOgVUJzbnCbe0wE6x0ElHwljQaxALX6DAgGbuSq31P
W1+kYIg1obRuDTW4RE0ZsKA/y/j27frWTepp37RSAYZoAPLd/MMV7GvRDA7gHUWe2W9urykaLkr2
XoRmRCYxixQIAEq4mP2M3n6DLkTdlkakFsF5Fk2NF+C8dtN0pHJYgNaJK8juoprmofZQBH1/PPiD
rkb9T69AAFIhOb1IiFEiISETlcPFL9qBg1I/PBsYd7HZTc6ogUz4LE6RogZWl5+FFO1s7olG9Q4V
WMAxJlYV3XRpnddyqO5ZQsfN0g2A4Pd9hMJxxcWDMCSK2wuJsjHGx31b2Ok9oBJymZiRD5FnFE7S
KlFYxjKOYgnVip580LNz1TaOyfK1IbT6ScoNcbX3hXSVqqG2D7TappCV1tyKdtjMCOeK5a+mJgRo
rT6eX3smAOQRIWo5XWPPd1VpeH0ziO/7JTGl6ANURelkr8PXMUsLHEWPgK0JXGBXuh5zsiyHPxNB
VhHZ6P5qpsG2ZwtmjOuONwNimK05e5uufFm63y43ESfKm/0WTvn4esGFsVH4om8zmmnYNkXG179C
wfsnPOS3BS13Ch6fBX0qhWIG0fhiR5zi5WDIjgZ3oy+cxzouXTybBxqP1MhofdyutJqYw/MZmjOm
WMoU2pVYBoZEoS3FHz2N6X9FzYF0Y5JHKZeF8YGB/DWMZrLpewvhAE9nR7h6IoElBqDrZCKC1d46
gEkzsfuHPGNTcu3EyoMxEHMu6453vP7xPzAooWGhpD4UUapstPTs1Syca1PNRujoOmX/ts0EO6e9
/IXJoUk4p/6hjlh2Bvo6ri/d7wW9zYjSghdM7EwP+SM1G1SkQKlcxAOqvF3RHQ3MM0Ufb5h4Xa+X
Rx+sRvi9XPyiz44RjjXiKd+QNEPQZ6zrjQEZmluJ8wbp7wych8trW4FAdau/uY/la184J214kJ6R
6Ywwmu+ysvRSYtu5XPReQg9T3dVxryUu5PSTB5XZEelup36GTro3KHY7yreoj0yHC8FjP+/WFl7O
hCSCQUJJYiNtdBYaN8FmY4E7yBMZm5XpGSr4me2o7EhfOKAgPckG6hU50u3rDvk31EoZ2e2Dd/iN
lhOzX0XjlftcPPtT1OkS15aGVF8JTl94C2Q8xmYCPMudF0VbyLgQVxlvzPbKNk+/5bgaZapyvH2R
xRimZw4Q6DIu7dMWyne+4jRkYCvVrbx82fD1/iZTC7NitROBEEd7kdgmt4LzYOGG9sgPrrThcFg3
PdS+CW5aeynkJPn+TqZtof2UoP88zHfOhf+SlOOejlhB8MWBabiurhU4B+An4NQuxyUw8urY2bPu
cXCQVTzjx+Fo5tCCSQU3vgJvJB+GYIy2Uc/dhHTpOe5wmTLGse5KxpNS8z5U/+kHtvKFGSLf0uWW
j3dzVo0Qn1VCuLzYrsaJTbWUxiGvh7XDeA3FdcWHSHOHxHzHmbnnalAqV0CWKg9lbKitUE7FvHrA
kAGptlgHHYFYwhIfljNVS/LeXVOaHZV6FrcKwgKxMfWr2e91E+4DCip3U4p3k9eSbudmj/MIj1V8
iyIZz67NSCLHMKJ7MPvDSXcWw0e2OQs+zvx/Xj5H8FdfjIfFNVwU4173ok+0TOYGjCmO2Ex/XmlQ
/MQ/MBHQ+pkgs2Nw1K7qhI+FlbLjq3xUVj5uEte5snY0t+gV+5pxc4YItrNP46ddzz4pvfkGI28q
xOOR81BVIVx/dEOjJVfGIdAKLf76nUtte86ysMKzqdXsD7zJfP6N3IEosyqFmNNq3K47jBiwAFMS
44ic+YLsZvpsUd7CZQpbC0/s183KdpMXuimfO6tzzZ3Oyj+uGBoGYh8p+1DuOOZlFSHZ4OU5KBPK
C8nqUPn403i1rMbDa3i8ygpWmnxPnMO1QVl9YV4ppC5wIc1eQhdltehXA7gFp7LewG1A4Y2NbwVs
b2RIRFUBtZ12cgjOh/yrlPO5MAjl56xdTvYtWAVwMT8n4SrAl7gbVUY+Th1WS5Us/8kx2pCNPw4p
iz4515hXY/cZNJVVzjVXI9OCb/6zuDk8WmQVdK4+sfTV9XC+yiTOiIvgThaHdzOHgJdG0rM8LJs1
24KtiTXFRlwf1D8EhtcB1vU4yZ1j5/J8h4O+vine4mz1PHutYH7WWB8cYUZositMkUJZbgvi4ea4
NeFH+6UxVDpj4U21ZBQA6XURF0d05cDXK8sLVUCSX49Gxokk76nf+XPZpa9/eJ2/2wm+DLX+2OJ+
P8t/Uzb+9A9ruJQDyBFFILPjZPIJz4//Zv3AerzeDcJphjuHS3TDQ/+9L4EJ5tX8w1FDtt6Vnj18
ZNTnc7nHxRdpYYtKwPzkBjSLECwm1aXi0qkrx5JYYP8rREqSPHx17G9dlmuE2VMjbY070ArNi2om
XN0PnlV5l4l+BN665Iuq4yS7+BBnczqIHjzHWljgfvfE1PtO5g5k9gvqgNs6mOkkbx/dOFwe1/M7
YHXRYOmxzvgFcLfmlfAb99009AWbZ1j3slMa5LoNW15iXOF+3Minq0k2rOHW2BcMd3qzVx2sKcMh
VowTvwBGLwMsMajAm7V7U9cZUPfIU/gXM3PZEMyPOhJvT+RRGuhBjgtU0KSvSxhe0ZQjxQ5wN8bm
pMvBOekDXyS+SKxO2VSVc2cdY6k4Si4pb/W2QnhaTeJAMfSFCnwFqRqEFgGOD7ZP5kva157cdyMq
BCsuNU3zeHDy42+7No+La6KZBS8ZsDaBwjj9WLpCp8Wetv3BER8xav9Qfj8CjaIPZtYrdDtvpKj2
vy0+DKwAsfyJqs9ZrbA7Djh5RnXv/c23pCLz6yaUSeEUnSuxCgUNB50JQJrb0eb/juzc/TggOH9K
UIMQYU/OJTBi8jHj1vVFTIaC0InidHnBLjmyvKXxV9TFjetLhZf6olJFy3d+CBlsZiUNwnarBlcx
tFNjVZ4lScrPGyV4K4CoCxRMedrRsXKaUfABXHg51MBaxl7NGyHnhHqg2k5OrAg+8cIFD/+C8zn+
WkASw9gmO8rSg5rGExTwR/8SMuegx0Dcm0dlFR6XvI3NSrDu2bQ9EpXQSgjnZkU0A/wcHHDfrs7N
4c81Udg9nOCIEay0Cr2HUNdenNqia8lksMBQJaaYkZC52yp+SCDFerRaIMInKLqh0vFh6XCwf8rh
SZgR9k6UmAL+MgN27UV6v9OXbVPKOWWIdtprR55G53sHwaUZNNRYcjC1gNLf2Ld3seSjNdciy4tD
PZ+VhJZ7c/iMCtGd8skfu6gzU52d/kt0GF3SCHKa9AGJ7D96rIJYq3AYR62YpsOHOg/y/ZK1RVhI
6xFwrsIJGcGhJvFjcdAuYOYAFcYyExbsQhOA0SnKz5CuPP0DBv5GhN4v42tkxXh6l18XlAzavOPN
hz+jOWmtjqAqcxE6ppf1t+Cr7nd8fvinewvheYhWWGpSVrku/WDQhDwOPPLc/X9mBeK7tFu9qn4U
CCLaCixDA0N2PTBbhHLE/tlHot+Xq9BTeUjINYB9XZHxvcMcrP2ptK+liLV1lii6BJGxKR0/DoTn
BU1OifVq8/bVTTaZ99sDfugHzFsnqCclB6OPmNj5NWwhL2m3B2Yj0NnOMuZ8sAM75wtceprlmkrV
i42T7LkjYPdagDE7wHuqUfT93YPiavtbFPWz4KXGaV6/ysmm0P+0pX6Z2wITGz+k7HGZFyK2ln4s
47b8bQHgwBSIoPVe3HFWtZtTC2GY573AeHXfkH9Q+TLkjkm6tOFXFUyF7DoLV3xXQi7QeFd1tLbI
lC7AcbkR3Gu3DeBbxkY2umoZVbDoNB4ZOcSQdyWjU/VluC9dph8jilwNfUoY8gF3LUxm3J/aBT6G
CRp2Vy0VsVnrD9egaITAXo4bQ6Jkcu07pog8i/5mEXviMwzCljvCQdZzOTAWbTpTctjvDigRi6re
rEvfAHr8MAU1yLMdMGC4X3EFl1a+EsxPsKNBtrBWZtkmwllNOpjLHnbAkhDk3PhuxbXz4+vosqNM
rcy78MzsfLe7SiTifRoUttavbEuIXy5CDqPEG9l+7qh8Iu1zV9sVB2OlPB1rhTuOrEHCims+4nLO
fPdNHpbxszXvN4rhPoavbFAHTOSquLeNtEmk1Zq+JUZXOW4D2zTxnGWRMZOI5K99v/TMUfXZCYzl
qZBPLnP3QvV3TlMLxp0bSB07YQnahYD4e0fCBU2FJ3SxGyIYnkJk4GMrW2K6tleSZMWqNEQ6h9lO
i4e3YVQxPtgzVsdTB0E58Xmhin3l5If2nVezYK6659PiqJVU+A/mvjRu4DQhoPw7J+tpWnvrhSpL
UMJ7U+YWfIBL3lq5ZTaFmurEWWH8pGEu1fTBhQ3Ma4f4NR8I7oouv9QydRUdUMp57En2cw7iP/rf
DWJ4UucrrBrgbFzhe7m+98MQEsjSc8/PCzyu5w9D40ljnI7kEuV1jzpLcdkLEzytI+p619pVtUkJ
m2lXvNW1bHqflOIXO3/bpGSR2M4Q8HgLIfNTilASAnoGTuYSnpCe3kduZZYI9jkos0R/n5IasLYB
yNidUnwkBMKTn1vj2zv3YapbmPAwe1K0dYD35amlLuoaFcyPEGRINTZH/kLL9V3LYbjzvoZWsnq8
saGSoAZ7/7jEyKF9HQiIwITBRBgbbwRvsB8OPcYLFhYLTz7aJqr9hhfwZ40zNPQwt30o0UOaxdxp
JAmfhgpekTP5bjXVPCSs9o0x+RGtzkClye2ooeM0Mv4KPIu0UoHpkS/cySDcf023JlKKcV922zp3
KpPYQ4YBflZy7ubdOJy23PqvRPYoaEV7Er7zv5yvL82JTRotm35ztC0gOUR1dyVGkn2wW5WCRjIw
4VuCtMeXr+hQA7XLg+hfM4LrnqRiQOLC8b+KQtaYskEtPRTB71pngmABgK5E0+CYc6qme0TgYQtP
5ukfyFnNPPLfBWsuVi9tzhwEVUyHtDBGbPs3Vx0Zz1pb59eLAi4TEcYujPgHjVCfepGZ5JCEDbmN
8LWhtTYcVdlXlkopX3VkS+R2RMXMwgs/v5XRVGZZaiYslozgsXUlvc2fiaC1VOnNtCAapbZmX+KT
n6bDGOsxsXySuchuUxKZBGH9xrSz4546sByFRdQ++cbZxoyVEMU4nKo69D3PyQLE1qLNpO9JIxhk
IiC0vHrJyMmgxUWlSWnq1amFbdhywgSrkj6RoNM/BlMABR46CBv9K7OhIDi+ygYE/2DxFg6i8VF4
R9+IjkHauoyK4ryXceyU98IJdp2F26v1zf6ek8uGgOvQeVfC06eowVmtW8dQYIPlIsTUNBKFHjeV
/TcP2auPPjs3b7Fiw4JGwDwC1dXrIgPB9OLIQxl6j2gN1jULEjVueLgTwpDmx8MqagUubEVQdjmv
NnKZkGbT+8C+cmXg1wLA/FHwUNO3kQKIfK9C27d3o2IM9bqYDMLquqSLD9p5R9kDlv5qj1vS//IS
2rLabrfEPZw9BdfhAMncZ+NI12l2lfHVdiSrKIGkQXsxYDmJC28KRwqWNXrJNZ91xI2ylj0bFzP6
n65xoT7JGSSHGrSd1vKCKYZA9NipjPdn7xWUuiaTrJsx5CgHW8aFUaJiYb0bXz7WiUOUVdJz5gmr
FuZAg7psNtMhpC7TpeV/kkMzHizfCUfRap7d7ESfv5R3pPHMcym2jnnykL+lFP5m8dsU6xrsr3ij
s6gYRlRKklPmRSkawXc588zgVLjaJqXyVJdAcAZUe8yUpamh8xVWMWRYtHcNbO9WCR370JhLiQvU
WmcySs2sC+L7Ft9Asx0IPWlIrf87T4NO4zKS/MtiEIbbrEMXDkcyTTUk2ahNaVMe42EKZ+KqK64y
dRA2cHUUIHANqAs7HJ3umtoLLVOZgI8g4uOu/qZDA7sjbrt4sIWxbdO6H+NPB5YPrXTOwODgVZHn
FdPZOUBspzMPJFgPLz4fbvn70mzSlT0YQUYCYTYudSm8yOe2T+qRVXWY8WO1DwHOOd0BKiGrYsNb
FUHY6g9NTkN/1FkYaQarENaXcV2Qpe9oUSKzFcq1grTkz1EwRl6jhIsPDiz2A+g/YSWetjs3vCDT
JzBahblaMQIGGt4G1YyR8dLai94OujbrSbq5u0Q34P0ZkbaCOdhxCxHAyXN3mvbVSPVuUAJuYQ0v
h7sV6Sgz1FMGE/JtGrZGSEacd8MIBblHfu37W58XDxZBu6MMdlEyYo8qtDIVeCwzJzYjBWX8DcUE
2ZB2aF/8zg2t+vyTgW147u21iS/BF9pcue2swckzqLrpJOnEQaY057Sp646PdOI3BvOXR3mkBUjy
Mu6I5YwRmh880TNN7EZdvjZ+6/0xLpw8HQ11f25utEnymjdrxwj4nbxtqQxv4lbouiNp0bPcqL2k
eq0uRdMK/E5c++eG2TY7xzrnlTD/0xNhay5ATf0PC9O1faVm/pIB0vA6fAGhLnKlsQRe8z4/YUmM
1k0/VINm9vplt/ml4szZ4lrcnjSRyph7P3dLSpTOqNrU4/0WYtofhSalPOCjrgNCyLv15Ti5WSwU
pKtrm0gWpYBiCW7jzCVQAdBMQKhwFpS66MWdMwMuKg+yXsSMCwFZ/MFiYHJK3+hPCcVSPFeTmY1/
9N/qLnO3oVMCxeX94Q4xTYi7+/glihQszEu2/kj/XsgRjjcju6HF6wRjhglhy0kuhJ7UI7jJdPDr
4Uir4mGEFGOpZahgZ1kbXO5fKLRnbh8fhOs13pLx6UmJsj+TV/WIOiFq4nnLWRsXn0k9yts9024q
xoaE9qGRj9LRC7MVtISLku+/ZIVEyCtW2l3ja4NKAQriTomVCXXCjG5XW9nB1G2R9dCLKScWxAhe
geNhqmfpzixGghjK+bhe+MppvkqESi+NVIgj2E/Aov/lmT1M1TPnJtQm29LYfP23p5O9yPpCtgEF
Y/eIocsDQ+t4VnCeco8zeJ9EptnIJkP0/Yof4cG+o4pbSGbjStp22199PI0ZMEajMZDZpRt8ehiA
FsM+/9g5KiRYKYhB2Rqm/M27B0Loq9TPPdsDSeSgosKxVnH1ra+T+st3/mDDi8RBKLZe1qE5R5UK
RgVo/8AMCQ+BsL2LK4WoJLlI2XL/UDsFgtouOhqRtoBmjbb4f5Z/5byOB0+BdQBTKgztwJPyAC8S
p+dhqUGsNuglYik8LRHagS2gMMpzrGwP2eetBb4VtEwy7JoCoi3bbj/Cf2BtIdf2l6xAQsvT62Wg
q5Xomve/Cvydo7T9B16zXS2eSI5+mXoaMMGWyk0rw2W+i6k/sRewG7EvdOqBXcle0ydN8sLV8Wi6
JCtKiMyIboNPetzqN5FZhmVUl0zLrWSg/XvN0hf1yDsR1BI/SHuKp1LwbQHjpJ71Jfp4T0Yq+xAP
9d0UxWfvZf1pMbfNIQYgnECUzjy9lVtWOXPrXoiw43OIGrkTHB5F7YviI1ZKfQsVMBegNdBNOqbe
okOSHm1PltgA/IwyXsdKDparUR8pE0kf8BcJCgQKIYR9OJiz+1VQJmSRVmOZIfqrpmZf2xmC2yS9
l3fqW4e6rV4fi7hSr4JGH2AhKY7WbKCk45do3/wnY9XMnbSRzJ+mJ92A/14GDZgx+qSC14zzQJ4a
MnBw8zp+qM42eH4P3ujt7o/hU0Uu+rwD6SxyZTNSJ8kNB2Ypar/QZyCt4zQvmrlJtRU8OvFlwFHO
ArjcxXx6+a5oPcUQnv16MKx9G+Aymu6kx3F70htCmV+HfxRHK1vrwRcPguq2gk22h+4laLx3pLNH
wR3X7uf5uO5rnWGjOp8u2RHnO5xYhe7gzOGyItCbMTE4+SGWY/Kbhtc5xaSdXXq24WJU+vx2Idw8
RnwNTUSYUn/jwfb2rbGflGz5zwUow6mwyxf3ElXZsSd9r4nZJwG9p+PjfxaT7CsF9trYCAylKgAN
YtI4VAQ0BJsb83QmJHuv5Eb7fYjv0ItMhYVD0WV1XsU2+jE562sn/u/H2GdNPilmKzZAXetV7aQf
hvjewPLLNGbk7TaQ+FjN0JbJ5eO4k0oOJAe2YAUNBaoPjXzK5ljeKytNMfDfncfZq3zmUCfsVA4E
2wdwIizah9me+Xi5SPJ0XY4S10++88CbvpGk7PaGE0o1KQQXdK3R/oMcz3oZ455umz62rsr6eu7S
H2j6a7p1rEV2RI9RiV0PkxnZYqUcwBA2xcWBVuWqT758ZHQsq9N3AMbSYgcbwvBUZ7bK1Duc/0Sn
gcR++yvwvDRblF6D9qRMORWQ/hypKxRg685iVDr6gLAXiDC8CSyRh5+YwOuXWA9HzRHubuIPqv4j
q5O0wUlnzIj8USVXXWHEHFMe4kjaRHd4DrJDJmwVZcfs6EIW3bBMevov37VkW2CPTQlV8GIxwpad
Jv9DPt/Xv8+pB/eVL8czuj+9jF63JNZxIGLifrASAZpgBjcUXt5wcMtW2XYvyBSdIEsJ/8h3XThi
L9qF96/H56NAXF/Z0fkr8r6zyihIGAPUf3fpXV737AW6kMsTvnIz5OK2o3Zr3RmAIhn7KPA8h39Q
LgmAaksR1A5EieL6JapC/Xhcizl2cQTZvBRA5hHcuqm0HJrWvWtAfTgHyE3jGyJ6Oz0PVl6A1OmY
ca6QZJy6mng2GiDK13yb9aHYVDl8ExwlDTiHdalu8trKYBthMXbDQlF1tiNGf7fSw4x7gbmMfpK2
FeHkIncgMoU7wCI5OXQgPr56ljkM+0qMVRdTKMQpREuR1q3bCHDDHclgR5gX60p+0rRTPwvkuNoG
t2cCN9MmreC+cjEZEbn8iH4L1oK2wSZDAZt9mugbfyKJBnj60nnkLbHbCHIPvXY0+uQEERyTEf1Y
DJUqMTOXbinOerRKbU3XAdxgoPpq8dKixOg6OUSlKV5CbKmYWh1zD6CqV2umezsw6xAXsQDL+Hiw
aN7ewt4dVrjcdJ66p7u9wTsv5t60lso/R/L16Po3pqsvL6FofqZHCzmA5fMPmt6QmQL5S8kwLnD5
ab0UjJvpdmjPNCOIrY1kmmHht05GO72W56tjrcw6xnrY2GvIVELbWadSUEVsFMX1Y1bPCxZBySDC
P8vCV8jcZ+UbdZPqGDwOoZwUxw7Gdq/c/2gVgFbT292NsprfNut1BdeUOfHjEBe2pBA1q2DjphUR
a/AT+AOuaiZljoaE+7A9ODq1ARX5Zpp6aBZOI87fBDOFBAm2LzrSD18PKj4BMGdPJkpq+vpC8q/z
CcNv9ZN62bMOs4d/CgjLIsECP7akVCQ0cFXtqYQW8L/FHn8AA8LIquCpNDe8lMpzQIbNJJPFlL5/
R9GrCJT7dI1xX0jVntj6+0tAzLQkovkpD+rT3LUwmDBSd77IETI02cwwedWWVJfF9G5ueBf1Qysm
818hW0M7siMLgoFhlkuoInr/xRRq4ytLcNP5mw20Gmp9rfVMdWZTC5hnKGZEog1mZJ9Gip8C9wzu
cF3g+YUsKJua+gncvBsPfrO/ip66nbcwil21YbuG5oOccNPQhLQMywknqQv4t+uWSSSR4i3NyUx/
t9Q3n+y7gvS97c2BMSWuxxwpuKJySBtQR1rFYjwkCvo4dllbGMXtdBjGiUsJEuQgCO/7QdUB4+HQ
rXB4blYJzqiDKS3y3xk5l1MrdqhKelxPyQ0gL1ffYrg3fdSHeedv0aebdu1zhoIJuFpKzoMAC3It
FPPAjEuktSE09C1VN21BkH3Q3qgJtFNcm93wkR1OfSBrUScyhLY+yENfx7BOxmfS9WSdLjUj3ABq
bUeo2DoAFBWfgnHK1aIiiZ4ASrocsd9dyuc+mRWrRWqinJytpgUF2oi2bpil/hkxM3XKKOT0cuzJ
vrgGR5Di3GUN4vjdNJoxCIJ4s3I6rSE/RPGVxv/oMu1r7Yy+6xJNUtWHhfdpPcFb9bBVCSMgGJjP
q70NtjYzo0WFRO1TBbe/FqyrAxZvadKM25jSnFkmKEQagL7w+hpGhrD3LsxJO9xPgiZT8GvPoUII
/WL/eZUEJzR67vBT86fJTfgYCfPF+U7E/GDLYCZN3OPDuThX07nwVLzlrQbBPaKBMnn4/mERor+I
LxgK02Gjy+YEDjIBKilv+/LFUo+Al+CrDDe32XNCX0QJ4gGkxe7utaK86VhzBCQqTW/mchMD8VIN
KWN9CX8yXe67P9SgoLtI7U1HmXQeSwMAU0yNyKEJU4xglyXh982fRetI+RjZ0YDNggeTPbCVGjk0
DIK6RTw+YjyiJ8UJm2jeRcFojXq+/X2KIDTHK3hkHPvALlW/bZyzrMPJIJGXznLY89N2Uyu5Bq/u
rPJdOCMp3gDqWLXji+hQNWDROUjSGvU4b0gw5cGaZZ35VPorKMcNoPqCTL22HV0XI+dqH5FZ6aOp
VEM199GTAVshNQhkeDo/Si812ugR8JgDS3rO5T+wRo1Az+EDIbjhfkL/WRkxaT30Ta5/sCjLNT6B
X8cOAz/P8+5w+i70/7QzQeZJPl8RdNy7i2l2e0qzCRCTS8NAVDvlJe4WuDqymxhF1GzsAzEFJK32
wSdSiiNV49+b7sAd+iQ4uQNoW/L4DMOP4FyGbktbkNJu2g2VNAhPMbzKiuSkgYasf0OQzn58WbY7
fo6u18p4o7NGop4f3XO6m5iHd+A3niT5berm4E/MemakWXOPBMJpIwdyOsTTduaX3I300hQbp+hD
GtX31DDdJGckU1S1teOdi0kWymZEzKzBuMWjs+wK8f7QwTNqErlEgzFyH+HMz+5/08vg1ocgXjTH
fkkDweRtrkW06NscwWhWyRYemK/nUtmEu4WL3RiPL08c+Lts6DmFhlGk/V9n39RHC0xEdCiRa0BF
E8yJPT8Q5qYAopMd+CLJbjAw8WRQ4PC3dYkycsKxQ1DCi8kZrBpuSkP+mEPauhTmgKFX+zKMwQH9
bAGFNzK8uzVlqLTjA3UoNn3cxOXfuJfC1gsdskFEkgZgjot7ZEv3RZZUT/G800yKgrYbFBbXAd7h
MxRTKhHggCXUgXvHvYFo+qchSavNXTCj5Ttc77Sl1jJuVaWM09wgxlKox5hBDGC0T0V7+lAiYWvZ
+kzfgrUVRY6j6I5/4Xabifm8DSqRTlFmrjiFaz7anyJCWLMo/VROsT8YKR6zXtmHMeDevZBpY6jg
EWkP0UwsfOYOHx98ndbD0QjWJSQLiLMI4y+r9huhQFZ8fbKlpU23vS5l6olrFn3QCjuBdtxFGx4a
sp5VqBhIgyldGbPWRSkGAkNGk14qGnM6TuuFNmckq6MMhI+RY3vQDoluJUgdqeDbEQpm+AJUmPZk
qEEMMF/tH/grJyvcyKFcsHVk6ho8Q+rmhs4/hI8c2vN5XbnyNbF2RJD8AWSIn0QIc/a7odFSf0gw
JdtNtGxtdBiQQU64BDrCMUKQ/MyxyPo6BFlXzwvhP8tzHAfB/P0UMz/V/+68H+WXSvziVVgQZEoX
0J3tmYSa7w8c2fYVB8j1QOAXyFW5dlk1EGJlxtiO6FCIIuM/L2yW5unsQepFi1ujMyniIzwBqkJA
c7NVYi5QAq60W1nTmKGB61XZO3WzYwajp7IS2WcRtehUHdQ1PZ2N3o5+MKMnPNFVUi7ruUXgy7dM
ikpwAyiYQCS990hQ8CyhThEHK1eTiWRZhrJqdSIGCzg/TZkExM+CIeQ2AWu1xJEVCG82lynDRGw0
LmsvD3+g1UN6XPP7yTr4s4kVLbJnm4N1ecZJSzp19ewOOs48J1hAB3QvTEFsE0Oqcmx3oVigH1JR
iSTO+rbD9bktnhY59KURjffNySBA3vLsPWktaEY4/TPgR2n9hvVyiQho775SUOrvdzHzph7Y21P2
+/0WYmUwVpBcTzDkjzVdBF/ylJp79yabnkO1WiCUb4n7z2hTPjnvmvHlrp1NGIaiakOxiJwxxz+8
9LLQTygOtZN4AbvtEr/6apE4FUpPwwv1xFbK8nnxdh8i5U9eC3TX6Ynq4bFeoQPsn2IHbRMqzAAO
fEf/MIV4zJCy71FQSTVYevP+4vE9NU7oXEEGgQ7vpnOpqObLmYHjAcPUP/bL0oMdK4TEEfg46DaM
5x2LeimVjSrO4ka7F0YLNgkJjzsuijJgfHMv/d+9tYz2xOTetKS2b1iR9+8Dqq9tBWVQ9lMenDn3
+zlCgiDV54XQLymRaeVxURUVOVUK2b0Gw6q1IBmZI1SPcL+BHJtBMiBhJp7huDAvKYoy3kKOxgle
AMqDh8lCviQXE9LIlZC/z55VzLv7iJiNxHtXR3VRVw/Q36BXBt52vh1BZRZPCKsZbZOCpdO4mqdH
ZHeNcx7gg0SbDexIjnhQUmExeofVorvpI/xwAsoqo/3uMweJ81lnRD3q+8ETqzxOXT3/Zscg/C/O
iiUv/ToMyfUiPfZZwvnaRQsMj8NscvKpQYz89k444F/kt6HnZlpkA5atdQerr2LSZmYYvcxG4/uk
/5UDfprSdrpCmWs/i/Li8cdMOBdIBLiEdhzHHmHVjkT0etP1wjOT3Z8qPknsuYw2Arwl9zYs+Ew2
ewutPytrRUOeM8AEZPIZMQWoGJxSENe4sDt1yeyKQTnre9JODzf45jwtVklFAHhvPxlhR77+mhr6
ykqNsDELlmbg2wPC1XlZZ4bJhvLQxDBPkiLlk7a1opcS7477TBm6dRHbnkBEOeoVRDNrmcCzR9Q5
ta+5vh+3hdstfAqE5msoM0Pq9om8M3aYBEj1jJHyZVVQnvkRMnKLKQzuTVeTpkQE0Cb3ojlLuZi5
v7pojDRWHhXhg+POn1/8Zc8w8WMXMU/0XE6IIHWYAG7HwSTafoquxcKMDf97NS7hhkJvzRoGH1es
cWKDEItSxUN8awJtGmncEmiUdf9ryP5ln8IS5IBR006ITi3fOhuhMmzcuJ/ES6SF7ge68JCR2hXX
BGaJEjDGNz5JTcFp2y4mToEmbIJdZbTwp8Soe2IaZrPtZ0YRE8yVatIb+/J+kj0U+6uPfyBHsF7a
vjYuGWtqUBfZPrvLI7/uDCzNnNZnWhBnhoGWTjPhKPOMt0aGH0RDzaV5Ft6LnxC65rgfbkfscxbY
2nYJWGD8obajuBYe1YvcyLZ8wWiPGEcDnhHcIYW2pMKGaixHOL9Sh0+dLRzSRDK45XjRT0GuDFLV
00bKlgx8Qy0m/kGR1x0w1ZHhf0k85kvTHPOcZVDK+eAzYfEoIZczfQDZakpnqzDL2MqK91ELEen4
v7FYW8iAU0T4T3jmAZ9dPKJ8bSUX7dAXQnFq9Kk5I3S2HqTcNTAZ6S/UYUMZVA/OyDrQP+MLLs4X
BkrAU6o5vAr2f+XbJePf3wEodsxyMbOlDW6+SUQFYemNaVw5IycaR7C/UNKEnHstZ5Wpz86ibP4j
sfFpljuLZoXZVqHjfvcZSiEFdN6YINkPv1Q5YiVpnRBA0k3EepBLgnrkylxtl3xFm4NTsWdx+dHX
+1XSts7Z171tsQhy0H+DD+eXd50/JSNMtWvYDt1irSqiexR50WgBrkKHxNHlrQTM7d37YMog62q9
zTioKOCVwCakaqUh2RROib8CfWj1gotap9KqdVyQNawWleeD8xJRm2MV5VdBrCTl/5vLkj6R/TVo
d0j2sQgDQN034DqZAIDsH+8IJzAgZtG2BSj/yBW+0smhZmJOMCCH4ORekhsItWpHaI2Ch3DbwqyQ
oyuowCxcugLxwA/wcyRIcuAFY2iTlpl6FIobzfrPENfiKZa4sP6ae6//o1Xl3ceH1JOpq3T1pBe+
nqvbEvh4FdOJWllkh22gFh5f4gVnuXNF4fpxJt/hnyT+yRpE/iD2Kze4xbJn4F4DnRQi+hopmquC
WMKvweyEwDmeVqE9Vw5FxHo7ag2O5j/c8gxFDzxuuwh9HLS1yOe0ZcDeruYwVZTxD8DmLAID2ZTD
Xp56Skbja4ySLaJ2i/cmgH2oebEf/v7x7zWdR77VKQ1QtoWOxsO1caAB7XGmuWT2z/CvGKPh30DT
9jeSnnTWwSa8bYQp1dZzu11GZcQ7oaG8z1Ai6XhnDj5o4gLm1Ikl+uJuyIHs6WIl4B8SxRlqo4zT
sGUszeEnyQvQ9B8TaIfXJ9Avbp5Hm/NYww2IWEwSc3StI2YkjKe2VSk9pzBmCTeX/G0WMd/l+us8
y8OQTpN+0GBGmJghTbJ2uDEvgIpJp5tqLtpBIi+00G48s8djIp2NsJo67TqhoKWRCt5E7K77uRBK
+9xap26b8yFPr2TNh3U+JozluiJ1f2R4qC2CuHyAsoNHaheuxBiFtpBIsJNAusScZCArzO2eUKlZ
czQ9QTl6P84gYILX8zpkMj4bXzbDGXJB6fchkiIPuNGMiQTI8mT5yzn7ssSjQ3eHqCVqtDr3qsR2
jweu5BwPSJx2awdqE4PTT1qZoi6AKmrU08IqzXRedX8S5eYrlh8N2XBmB2XNhLeivJoHzXxvxLf+
EKY2AxvQGsN3g9DojPx7naZ2ocH4p0jqwjMUSyD72p1ZTmRQOhK1wIbh+j3CH+4lKnAoDtXaJyPu
2RlEtaIMan6glKdoQO0ptJu89lxpIWQIyD96qXxMKR96BXyYelltqaLmX1bLthVhC668JyWkzdYy
VD1QalH2POOPKnVvNnkmr+HExk/y52oPHbv/2bnW09Ooceen7lvnAnYBJckC56FVKjf/1PiTxjix
MbiXAjEuowLyDSvTn1c2QbJ1PWfAmzhBgzV6X13LArSoTS67TSJeZRTwn/MznRvy1NjTGRFupDdj
EE02N4c2LH0AZ3NMO4+rcn5yjABUws0cRmrsTUUuZ6u/5acZZjohCMuARIhCpYwf5v0BFM7rGdho
1L6RQy5UjLm7cYM0A/nUvCVOqBkSldyeMFL2yFSIUB1U8XYFoTUu4Bytl0kZGwEhaVuRvPCrCwIQ
lCzFSg6CIL3GV/sYNSHfNZeisdEE0i3cfo0W151qXWvkRqmejzlvhtQYXGxw4SO+W6Bhh8jdZ+LV
zH5/ekTjIYocg5L0INeyig2KU6NDSmNZDDgs/A9wdn1AhrMxLtAXKsRhV8mgTPJWSL65ffdUWMPC
uIAZYr8J1csChqCgTe2UDxZ2gzJH2SVyvBbg5ilGHV0FCXPajP1MwzfmIH5XyMgameePa6nKoaVf
QlPXDcAmvSjsN9/2za2X4A1gf95TpwHW90BhZVngRy/Cy9B8dKH+q6ERDpK5v45s6v98KbOprY6V
84oyhht88vrUgOmJL/RzsxUSLckoRVkz5i4xYU0bqDSTNCDCga/0zFjJDsfvvtEKEnCWF9O0JuVh
6PxGwKz4L+w/Vp98WdC/mpEmI4qVfIlvx6jjA/Wk6feSg1mybh16S+Co/73hhjPPV4BjB44rCDi/
rBh4WZSfKHP1wj0uA0ylAUYC3efJ8bb47JUEyHpUjBKMNRJa37hCg7c73vL3vLna4zib21x+o8fi
h9M1NGLTmY5pQZ9HFU0rRifY8ccYcYmL83e/tDjqAo2suVLzlMhEfrG+rN/3/Ec6AASe7lPT19u/
QYhAdu5z3TabauZfdrIj8ql7JHyXYTuWyc7WemUcaeUWESX0j/iLW8gzr2+Do8g+uJNp86spKWuM
nwe0vC3ABsMU+cxnRWP/ev1J2CQUhAYUb4Yy0lEkOa7JJ/QYmFYXW4q3zCS6ZBRECkIIwxPbyjLy
tA2g2PumWc/upoZiRP9SS41Y74EUJ5bHaq+mkd/Q33doH/OXUIto/50pdq+n6VRLEH11EuAjrg6/
YEFk9RLBbdrV4yWk4dnhgcTNRsI/qyjQbHSqxmn+bBwoIvJS/9ogec5KdWTn918IUayDu46uQIrQ
gJi8DoKklzMIlDatM5r/2rCV2JlNpreHWxtrpyfn+EJGQ3Ag3NlJ9UBkwx2KAF/dyozrM8uaxNJY
wN8woRKUsonBmgURrzN4toE53L3M2khEvXYFQAB82/CBjYs2QLdRcbNYwc6kO9bEwrajpqQ+Jjqn
MQerVFuak1qD6T600OZ6u9UMTerfkL9p3bqns7i+f1Mry4SgM6RGfIzs8fmd9jjm/Q63C53r+lfI
yPB4AR8ayXEvJ+FXjuSbnjB3n4xBn+t9NOSO8r5WOyseq+dXEpt0tpd6VN0iIBsXCXYMwY7vgQcn
cp4cuKkXeMpHAhQ/8J94nm7R5f1q2vOOGBuSsQz3/1jbf3yXtxHjNmsU3QBLQssk4Lc+niSlVFHL
jpWKQJxbYNN7S06p5K8MZlItzD2xClDI82zSR9/WsbngvpDmWKOL3fPLX4UR8Mhd+r26dXiRsN0e
DRobURl71R6F4hp7O64Uzl/BaXEk0pM1lWnW/gSdnmw7EDiMzsaw2rg+N+JP0aiOtEtCG7vYQzzV
xU8GgndV3BwM+kGf0vkC29k4P0uutIz93eOIiERiF0PAW5SW9RIOuZQZAEDAlthLPrLWbCzSVtVG
orsItPoqwcd0Kx52xGO5N6cMvwmku6zSXHIyUda5jI7nLkv1FtrT+UScT7ufn6w+yZcwyWMuv54r
71bCF5U2eJsmm92gBgPgPKKN70/Ak7YP8W10trsVl/W7hUQKmVlArkUkOFKqAEYrxMLIE8lTBU4A
Jr3KrGyDaeunBy9JrcjxbtvwRrm+XUqOyiv8pHzxmOR0UxM4aEXOqx8vQa07wD+Suc3uzlZRbV1H
sRtrIYl60K/8K6orcxLkFlpqWImLwsfezNqdsC+CWP6iKsaqJEWJSIR6pH5oUBQ0IpXOcDMUUhCo
mexkB10CeyUdR3eOpKzvdqNXEdp6CYeNaCq2jIsWyibfVHpZ5SiRzzZ/JwLcP8d7GxrVfu72Cky7
qW2k/CBaszn5D6BvElpi4/+nxfgCybBA6DVNhR9dSQbJctuhIBMhU5E7nSMpVgEhFu0y/8ZJshQY
IJpXIScADIicPuaKQefK4HUm0IkNyYA5D3i6XtNh/+eqqUNOtFHeN01YDN3NtTT6lQlaLsteFL8x
YTjDPQRfuuSG7i9+H4K3n8OJUgVTUG3aHSTHpFpXIGr38jw6qLxUwthScg8ysgoR8VCTXGKe3jmp
SopmF/pEDLlUfkWOkXMBcyLr6ytshLqrtPBw0c0uautRYPQp6xGVfm4NsO1d3PzWpXuaNsguIDpL
xbSoWXEU2UDT1wHBdbxQb4WIBxj0FqL/+K29go2lJulVFHQVTK5QEAU8qMz5BW34xmTKJwBJWazz
eZWom9TmdGH2H25vryBFJ32+h0FveIkoH1uUaTEtU4E8SzeF6oZXy8QVZeSYq29GOxllanoWMqLu
eKWspnRvhWLdjWA9cykwBNlX3y1OJMIwa3Z2Kk668UtlNe4MH+tyCh6dalePkcykJJb000E4lyN0
5zx/N63qFqus8QNRhvWPYyLHXz0ahPxFvinSQdTaLGJuNL+KFuMnG53JWYY/D+7wJKaqKOtO3MFE
0/Xfa3VvTWmhf0xEtWL060AVFPuGluTEiKPsdJgHzQ5mLgrY2BDxCY0DYX6IyEY/coJd60zc/SkB
s3VTrfFqsEzKrs1WCk707ajugPfmEsIZqVt5acVsAcn37eOkKKsSg+teXA+H7AwtGbalZbucGsZH
LAkZX/bp1lbDN3QYfCOvS3x+6MARpEN1iNw8xxALlRceuPc/vsLtbahZrYjpU6y+vq2wU6fn8rev
Cp46W2VxtoOxLO1Oc6lVStm5CTcITLIb2epzFaZkqzW3YsBqxsFga0XDolFzeanRjunPeoKbOUHZ
glTmCUC6TbiWJTf9D/NDJ95UWorEOr/9knsiGdHdtcz6yd11iYJ8ZpaMROt7FrX8do8keJPHl48j
t6aS8usWUd5SiFhn52PpMXqNagWIA8kAlJah/aCLGo5B+me1XVDaJUPlTjt6BpZ22Br/t0GlIl+S
zocEr/BjLNFvW+vNhXZBmtldB6+RSeUocHy1RrlwSYpqLEjoioTmzIuLOda0RzAbRe0256Kmh6Tv
rsY2NuDcJOsSuSigSZ708nOR+l+7faPDvGDMhq3PxUVPEvw2mURCEMSHZJow6v0U9OA12KeE1Vji
cRrANzGFUd7AoedwgB4Hz+xm/drJ2Bf9oR8hzsEw5KepG1Mph/jZGSutJMVgxVbAxJFEp9OSS4lJ
gtLbBJtXe9FOguieI2KftSr7KoXvgFmTA1+BWEquo/yWbkcXX68d/JRAeuHOLjsWNO5KMNmhGJ9s
AW6bzyb9sGBYWx+vbShtqi5cuyzkkWjVKsi7x+ZvB3PKTN6CfVqHqAOhBWyeaddVQbGL4kwwbsrR
ZPzJHQIKIxq1LJEVoOT1b7a0eyUkmmKRelaw1quITQWaG4KgXHt15Yr/9zpH2B5GdOFkWXPVorIN
Y1WOVmsV8/832lui2Kkxu2Gt6ROv0rbpxm0rUI5sIxio+yqvGxRTCjAYWc2aBCKcg6rm5O4wh6oA
XnZ7CYgpWdxo+HV6HzCTjknccVu4SXZL+BDAj0O/kcg1nBq0sm/JWScyV8Qpvtsjk8uHyeKMt099
nAsl0c4cPL5KqEk+0NzpPKfSiJ8kPQHNIJRuJImYDeS/wLo9SACiFBsBqkTiSfNXMtv93RIFiKTU
MAWQoNOFJ1m64jt0IuuJDQ8stc/PhxdA6igKDj9t4bn+p6IEDkF4D1Yq+H59DyYcLJsCUWDf8eVS
7JnIfZXFl9TiDolpUocWcFhK03rDZJ/ej/bOprFeYtuBKwo6KZWAL3gY/1XNjGJok/eZEjHfgJLB
PqzM73BC5lOfa5d5HMwYxYs5ye86SGK0E/xzBi1epYFqykryCqSahVc5DezvXvVPUwn7HiUWSRPX
kn9hSmnTKkFx56cvSgzfNPUDlPauRfSr6qZNmgKyogbgmPdcNEDz1O18par2mZxjXnUzHNJ2d2lz
Ipv/6C4TiYPoVVGkpnbCYVXtKi+iA2EgOo8OZNgu6MQHLml57AsypIHxO15sPh/6jPnR5BBHyIvX
3wJSVSyQ4v/njARNw/b4GPn2G2SetgYlNHTYOXl+EBeziyFW91U+oZqZ1kyOlSSetxo4kDntfVjW
T+WI4p1RxhpVzPusTNduquSiKhEdxfkXTOKDLXe5ecQG938BuxVP1BVdlnOqUZDu29nEteAg+LFu
ZD8Xe0+y0EWH1PQ43bL9CRrXsGO5kcb9iSc0aqdV4HuFbZ3ZCzXeq+paF9KPWoDZUexoU5hiZtJC
+Q1FoKRrS9RzhajNW+7YLgBnPKSxm7ibVFPvM79SrdcDKQrmMwTXdCGXtF4dShe4jzY/gxGc2PCs
KXapDRVHlhfzRnrU3yXmkKOmfUQPHPvbMF6K9HbwtMflyoJa113NMOzEXFTs5AKfQS9wk5zzyMVe
6wZseGG2GCbWeoGD47heVnAMij4+x8X26BrFvTNV2JiINijTz7uNpqpkoyGICgCKsOie2NfwaxOh
MVBJ0xLKB4vPzIQT4x68Sqks41LWA1icxh9EK9bfGWQDbNooASEa+1GoiHssqAIkHwWYRbhYJba/
ssInx3I5pBRUa5SRcmKYdv4SWUwXLj5J1+IqFq7sLekFxQCVOYPJaHSEystwr+ZAN8D6qKGIQ+W0
fJxUrL3hgLKML2wpIM94iqkDHFHxgmHDJg/GT/H9bjh2FNasmRrQaBWmwd+dRopuEulevWCcl7nj
bWWkWmA4ri1RZPrJtZCwYPYZyiEYiOJlMHPMQsuFLX+e1AgNXoWcU0HoPH1IQQAUyTVxVUukeLO5
Z0QgmzozjjC0PoLCjiT26kyD1vYHC3LO6QM39CQDgK2opEqVNdPEHPZ0Bg/J5gewW0/G1bDvv46g
wCh7c6EyomOh+O88bza7DQLX1Jp/PDI/nnXKF7mPwtkZVz4mIgebbfbHYhgGe3LF31DIJlQ5dvwP
T9tZg9DRZ7joQTjQNawCe99vO3OEa1cXIoeivqo8hIRuChH7P6jLilUMHg2S8ESX5i1Q2thdKJz+
UHQ0TyCXlKaA8QgULplmxDXZ0kqbNAkFbZq8JPAcKTdWKC+ISqiWIbRS0Ozkqwxj7TmC9ISWBINR
fxnJOwp1qt/GAt7Laq0mTIQOsXV4AdM+c9tszr/6cDY/ZJnQNnOL8e8VUnyo+p6pwuS7RMw6XjzC
UGBDJFn+XUmVDCiIObq4ZbRXmlQXF73L5Acp2pWfl/1U5X8FkJIhBKmPaQhpS2kR/dfeA8SNpsUN
NBgAq4l3pAorhfEACqPEc4+yxxyI1vhdJD/OMC4tVwrl/cravAbYXSs20R2f0sg2uZ6Ido3+aFBF
sELYq5cQ9DG/VDhT6yGthH/JSvSM3Dx3j7quLa0ZGzF76vIl/g1q2EnS2876f4IdUSCuEhZJc3IB
k+ZE88GDNPes3FXDfg2BWBmryjXOIjTT8J7wFxIRqBjH+dx0ZiXL85hYZ2YHD1434NCL4sY4LivY
RqWJvD4f6kD5qSNl+t1CozzPexpnZmqSg0eG81PcxZC3jqGdHPq7pVkq5JXRUy0eHcY0c/KdLrRW
PtHaOHFIsc08FmaeLSlo7nDmxImB+fZrIwQQk8YGKycdn5535osaXDgioclAFH4BwtYNEbUwTJlg
hXICW24WJHQeF3j9cQCXJNlSpHH/wU+QlldTaFdgPva6nt3yy4ZGwHicCP1v36aPrR8a/HU0S7Te
EhtCO/P/IRPtRyGPgabf9OIZOaAKVkjg9y/MATjKmqqfXJCVjkiKyNEvsMt2sMH9lzKndJ06t0rg
lXf1Z+0Rs9WGEPUbbAC1LQFFn3Uv0RrbNvTZREaS6+NTfuUMypDYetcBbJqp8htNIIKxvLtgPCJg
4MHZpuY0aosg6i7Q2PA0+ggC+jKiXdKwSe1sE3kmZwCamh32yryplkykDbMsNjcNqxoWfR6X9HeP
dYJ1ZLYcnLxQrEA7w747u3pPJj0BqlFfquz9itdHH4e4aJnGoL/JpaujG49ffrTngwKd49jREk6U
pN3pxVVcp8iMPNACx36acTmZ2RgojDnXn5MqFkV+sdrurvpYrfErwTvosj6CR0FZNpMzdahKt+Aw
2zAfooFkCDPDbWokBeAIeuRZpTVRyNvKhZyfAJecKBSyL0kkBWx8Z5y8Svt2qGeT9KOqCMrW0Jg8
6KGjV0aiEmCKbf8MS/SWQiM1SP7J3/KmiPo5FH6nLUd3YUXpIXEzYub8DF98OtasN3W9TrLu8r7u
M5BVC3poo+hpgfwE4BdBhLOptPk5V2Yu2Q51mA84kgugRWpGBcfByFfJFg48KXmQogn1KDcLlBg2
bwwg56H/c3hhq71O3zqKy7OHUsCsUIb9/4J96HStuW5v1hx0DY41MMktdnkd3Kx7uq73xAwk4wMK
PLtMtPLbnbnjJFVrvW+9sxdcSRKd2z9ZN3JhNmc/yqeV6qLWlXI+d05WuQvTqqFEv6C19PS3OVEG
7Yucky/ELFWmfVE1twb7UaMPrfpu9D+XuDb4YGI4C2aoKzATXRCCh6DfvCMWH0pb5YpsHIHtF7KP
lJyQ5xEwSNzp6Oyi1nqxqc0s7uxGGf84dur8kicezPNDBrMAKvhq2I+zX/GU7nbwtZatZj4+lvG6
1jDvYDT2G3upTzxINLt9mkZ/6wWs4EobgHQr8O8pk+66lg9I8DbF76bPHtByXBmEozKgZUTImQAo
WaX9xAxvLUwHYeQGk2zY8CSCVX4NrouePmPB+z0rmI+bGVJahuSR8T3naZJ5X6TbUe8GCwVh5SKd
Xx+DUdF2xSjzvg+n0exjwhiEdUJv0dSAmvRYhEhh4De95j/329QOydQZ1sZn4bd20lJ2JxgOXuxG
0V4A1nk5jYiYndcnbvCFYJj0Vytm55oYmf4GBFfUWIQFNQkkt+7ryZ1e37W8k/JYB8IKx/oHpl5n
yH8H0wkjsYmtJkGDYOxfcMNwkIDywj/Jhksxaci+ZV7wmtZaoCBvDfq1clEGw4Ke45B6BW8GFs1T
1j3KqtgrSwZd6o54ZawhonqYNtxU5C1ZoH+Na2HWSv4Kh9Om1fSh3VvwHKXFv2XNaQ6Kp06XJF6K
QZpevjIb5VAV25dOtHvDUbZmtCQZAUanjpJOTubYA9F7KPDbMRSP3Ug+c42zjmr5pw0kY3gmaplB
JEPS2VR4+JCBWzb2J5W9iutGwq9NwNICAyttOvt4dczgtVrVNHGPVcYdggxOHCBMzYB/THNkQ/H7
5WtmBrz0vSCA7lhL14ps3ByrHjkOL7GceEtwg4rGmT6JLbYwbaE7uRnTaPPsi8aVezPLnNIio2Z9
fhiDXFm1smmet7LSgOhbU9l8Qi+cBa6CwzGL0OXXtNGYlI9PdjOMqhiRtfWgKx9Ite9IGXuWYDzc
iWvv88qFS0nC97KmpQ+LtGtikTeyENtHUURViQUXjhQESTF+FoydC35S3to5liD+A1q38LWyUM9Z
NdX3IqY0/h7o986CX1nvV/f3FFT+BwPDnQ5CQztP1wmABNHj/NsOVfNq4+TDXk5cBJtunk0dZKE8
53DVx0NxXFA/DBRTiLnDmXWW7KvyM6sASiOfdKRYldhwmTcuGyg8NeoZIGdHRjtwKdgFWX022NVq
20uoaRT8t2RyG2OmdiKFzpayxPxjiAg2gbfOMP5hBzUAqMuOxr4o0n0jGUxreeNU6276YmTHivZw
J/vgkGa5fvnbTOYuaBG9qOlOKZwtnQzXUC5eum8ZHJiSeJuforrk8F+VzggLDLMO1aItP3gR4sH1
xs6+Ndqhcl6nJxkZzpTfXFmm8/Urd8HqQNw9cyTv4GOqKyDUinBIFRqNgM7QdF3WiBZqWE0Y7/Ia
SlFy9BdnRHIjjUrYjhUGmrb1t+zWmiOkpk6LsbmDDbrTevaNW1V+bTOEh9O0YyRzohjqexS9NQ4u
E8Oaxcs49at8a5gUEXgt+XoWP/yM8df5FQC3iQ7FChTprEdd6huypDdv1kE2LTlj1L2uLHYQx/cV
P10mT2NpOswJl9s94rGQLxRfTAdjDBER4n2Bh4/bHbqBX4OnpmxyZEr5j3EZZPEO76OlsG5+E4ex
S3rVomPfkDfC6cC34nGbk45h0/PTICAk9ID0yT8LN8aL2c+ChS+6FOauoHVSQCsukXC2LHi3IrHK
W2TPzBCjBkZQAaUFsM8ZopX7fFsZNQp0OSd5MT58DaULQPw1F7j5JcRHltqBCyyn5YJsA/kkPi5w
op9cDbOONt05EFCNq4d/h2Po6g92n4gLaoJTHOXLcK4VJvLSK4jqyyxvTfTeC20dxA860/ZXJUcr
0W+7oDW/5S05G0T+BYlz/mgNrfKB4N+XVhvvm/J20WaOrV4FGYorxRVOvOKvmwV4Uyo6WW4jwAY5
cFf5EGW2D+uMcJl3eQQLZwz/Mp1gCodf3uaaRQU1c9XqjYAjfXSf+60+NYQeHe3F/HT8fIccu5a3
pwqrTYiMLVahjzbJEhiNdgRhQK/yw7gBKyuKaCMo+HBhANCmVIUEiQC3F/qzrBKbyb7xUmMdD2tT
m162RZ4sfOu/8I6YwoCglYGBfWbDdJ6yMBLgQlml5J3Fmi3885V0ezIvxPhSnbqIttP/MQRhSRTt
EpJNGzPK1LiYmtBysHVWGxWnhfIeYK1BDFlEpgo4PP+3etbNqU78LWo9q7fPDzKEGVq+R42My8uA
4+EtW5Q1cnDK78ok4abZg6CzbuOtfuh5LzgQUj0ECk2uuQDwsrXE/TzXLcHM+cavNizExTPB2+Io
Y+ZTw7/ijQWUo7G/ngliAOiXiCZTt8Jtft7aR7TJfwbxQvUlQ4BwIsLUcMgfBOEK8bYT6WTi0ToT
LGidBbo+Q+TRy1M92uETC8fV2LQpNxR+qYs+uatY2MienmciF/g3ALtd/cQ8DqGKK3tjxcKmAoTg
08xUilj1Zal7QZ+b2/9hz1XFM8kIZy5q3x7YKwvjbN84FxT3SkoOx1qanfoLxo+OtOoPGYhCL18X
Amfb55+GxaoJ81lJkxrClBmgNiYR42ARVsfNKXp69/Uh2MrXZ0MQm6XTWyGk16yBqB+KZ7I3bYpz
GuqEdeIFr4VllHvmbOELqxdCSwoPtVRqxoCH9vPnivJmViBTc89VfSqJQy87wg1A5qRuS+yigh6T
TQM/d9FnbMVUGJBaT7tfNRbA4npf2E13ehUv0SW4DuDfq+pF67TuspemsGAMKNdOvSC9SBaJIQyY
th4EFWeICV5eiX1f73HkpSFXjq6FP5LQkbTbblqGqHsW+jQZQbOKCqkRZ4aXseBkOSgfGIfd29oe
qgYrJQcsAMv+PN89qfzrr3gRFRYPqnx/v+3xIcN9FkfpgULdVBodoNvAYDLIoXq8VzS3hqxDcDP7
yxpErWXeWSEoXlBExU+aMYcRLsFp6Frc7EnVkQpu2Uz2C/L96WktdtBdSD+fbgmAN9VejsTi+fxM
Gb5FFBR7O5zD1bAFqmpcyNCGANvKEcaGdSQCk2OIBUpLtV53SbD7SufmVzAPi9kjmvcf5v+d16HY
Gs3Ec2of/GwrJLBLQH1RnntH8unTg9RrE/vpKqivH3wAMbWJwWVI00r7tKwYN54xZVFrniJsFG3T
Q8ksSQi7GDZn9db5go9sGWc1mMTBjJmp67ZYi6Dy2Ms3/juyf5PKkuA3YB8bOfghhLzSQDzamqLU
RVrt9QvYWbXdRC7tyvu6NkUrhlfjpGxLUNo7ofMy4RhM3qkMBK8JW5hix039346ydAk8yQiUH2a+
LPZC/y2v46Q4cDs1Tn0QH+O93iN15IXHUkgu90Eu8/auFbRHR9ZLuMFxjmy9Wo3C9WeI1rRX+BL6
+kVBLRhzf290k790K01I9bDIyen28LJl6256bKqK17psR3leD/i7vlukJEe1f1px9QUaJZJJshi8
zDN7ZUxHPAXNAYYCXqP7mAIPnfu4k3uC0CM04/JZuBdqdkSVcH0X7tMWYm3juCdLgL8smo7rQ7lK
SbPsjtiphxm++JItwBaC4qNvBe6NmHub97YBZXK65Ty142PDwC29Y9XLxYSJ77Y2XIdIzSjiXz8t
Rklk69QdYtZ8ESidGHDczXhkgtkNfEKmSqiDCEYp62stUpisoWvv1Ui/K0reCCHPMHGL83JXCiKU
0OoMg3rcNWe6pK/91po5d6T8tU6ck5R6rF/HeIbsqCbNZjve6jCTu/x1xMErYSuRKxfvd9DanFlP
MIntocoAULLrK2j3f4itWCBA4OoKnvePMPZnuzNXUDnjAeCrR5UzgW9fsA1ENR0yNUL2pg9XIBH5
vTiBa2ZHLF9LR77FckC2gbmLRBqErgj3wYFF1yKX1bhhQ7ISg0QfYBcxvRHfum/rKgQ5yoYomFeR
UjK4gcKbuhBjIRspjXJrOgSp0lEfOSDbt5OYdUUdW8mPgtFFfZJuoFR11tAFPAFyFbMpBh+7Bpid
ejjz3OJCicP6QbApQYWL6yzEqV83LOzlGJRu+tn8lzeayDTY+x+HGHHkAEwnB55kFtUccLRvhuW7
uMr2FMLzijv0cH/6aTdDcGucIpV+Df9Ne28RSiw/USkx2Pffkl+g1bkCGJsjywy8g58lhp0wxr6R
9hlEc9JoS5IR9gkFyqpAauC41TeCklOKZeBe3HFMJaqb6Gg//k28BruQCOKflvcSMYzsJEt82qTA
Y++7EWZBj6EovP1FXmbtleTw5uBiCYwdJeBW7ja+68K2iFBlNojeo3Wz95Cb9wu5Wlpc4jes6Ban
awINPkdi0SYyymI4LkjHxzhM4AUThmbPtS50+BFBHw+9PQ+LFzJdIXDjfno63IYR7dK7bLGQ3k2V
Z7y66haaQj96bjIq8oARyq9SP1S4uoXVHMD7oqZD4G7jSMwaqIX7Wyz0vRLbM1HKDlLSim9Iksdo
kwWrMC432SBo/Omgk0qSjQjIrAz2XnOW2stj8jmsvlRwqUiYyWXIk3c9dw3+tcWfkYOfvVTfcXGE
SBHEVCERJxcBD+E22eR52xzwQ7YdmBwgVt9+IWYqKi4NMyURP6oZTmophBQX1fBq5931Ccu59rJ/
0ferOWPNbXIEoWg4jdn4BzDcMFLSRyPtL2ozK9f6BuHpt4umt9DjsSDvk3boLZVyNHcIqGzZ4bEH
1FtGwdoxhGZwhiZ11w2iE2notSChLHGfm3c5P3zmNowI6e4ScoOdf3v7tz0w4Fvw85CosIEB7U2K
gTOTRohTjnRA9VdcWf8w/wkWpKy3fPQr+IQdtgqmM68rf0c4Dw77aZmo1c+HHyb8tyU3Gj2J6a7P
Md2zRUXwCgtpxwbVYduDypB8yFjmo/kqoW8PYkwp3qyyCYdDOnAOHRiva/xL18tfTg4UdA2KpdUG
CgDIUkg3/UfylDR3mqpkXGspPa2Dz7BXt0kiBqFZE/3RjNF9sZgY02iFlvog5O/e0qVLrJ5iCIyH
wUbaCYiAxm9c7QyC9XT5vidstc30FcHR410P8+k9e88akdZaRf9wy52xozMqbe67dr2CtMVQsJ12
KOZIoSSEBXtbLVt4C2XyQnbUh+MtqiMznJvQ7LA3vXjHTk0JUY5og/G+SvcXL952g+5hcgvNbHPu
8ooxRFXgRdlF4yMTPh9gZ8HRx5Bmij56mQdxwTWFueBHIiL+oa/tmW2QvebDzkfauvvpWkGi18ne
D+jqz/qVOmpxANJAoHaFncdKD0tmOaN72s9/O3LRw04Slrw/yM8VPnoTk96JRcbqZnD+d0QiCvt+
fAGAMJWY1k0pCVDil2MAc28lwYsfCn0UbnT9AEtOHzM2nw90mnEnx5nGYLFtx0v3PvL9OguWn94q
JJLXZ3CeJwaY9TbLVV7QF0A4V/vH93v18dkE4Wishm/oJVHTdSWm9gvofqocnJBcosB2QOvVWnlt
bdErBjmAcyfDNjHGy8EV/mZtcDhVjdvUeGWIGrNSqPBAvteEYxUzr+sNygxz8qEumba3/eoSgn/n
Mq9UaLogO+XHJ/kVYnfagTSsOQQUDknX0tb6kkRjoVzp1W4QjCmywfd5t8l6fsHDKfOxTyiysAm+
39ZD9W+ICQIQaWUHZ9lj+DVThmyZKvAE/JZ+c20LK7bUN6kf4nhJYvxu1ScoyAD/GKLBiZSdq1Sy
xKKnQJ9Z2dzcLIhJab0tGOionW6XL1JUOEkoPjwEKIDHbXwAeG9IlF8xW8ArqRsVnYxl97eqT7N4
vUlsi/uNnStH0Qi3MdMNI1fymQhym8U3+aV/VspdkYtKV94e+mhZgGq2x5Lj/1we3KeZ9LVSoM+N
YfZpbMLZokvVfSo4aczOVAVSdSsWO7ShFskg4d7luaT9tv7UkmghYGUu8z23QB9ODoPY01k+N8VE
aD5dMtJ/hoZ8EK3egMaDUZm3EM5cghZzEx3olEVQJdWctlrxuM1qQkqKDlSQ2FHtQ6qYQkbwJRkn
gn/9re7mlRGNjWx0ZaNXXVvF9uVxbY2t/+3bKPNK9aC0+kEHc5SdNO63xZlJJa73z1AK/siafUgj
ApstrKprTSBeUVXf2vOxYlvWebBwWKyM/wl1+w882EN7k81FiVe8RMJbyeXrjibVti2GMfpmIAcR
9NKcHlaPICuXUcd2byZ0k2wMQFFv0D+FawV4z6fDTx5WJses9iNBm81W9Km5H61VJTwfUmZBdJ9E
VVe+4APWBQ8wDdzjXw3rtruzmKNOf9+GKcp3luV71aAMKMKeKiGkV8YefcBhrwv//de0zVXJNFak
FRIm8oRxyL4IIBTtF+n/Z1ZD7lt/H6lrIKwJOfp58UdwfaqJg8W02mAzECkbKfg15WxXmmUNPH3V
e4i4bYQk8OtoBxo9PvTY2bBIwQLHI8Cd6DMrOa0YixMLCFwgl6IrlA+etVMEDtMXbzDCtsS2cP2N
PvcKz9SW0yK6D3FH019FG5xioI5+go1aMl7Z17YvP8T0nKKO1X30CnobThwZXHfFJNWwL24d6pfJ
2e16b3kOrd1svN1WuAgpfrZuze9TVI+0SPgom4CgE+/np1NrwjEeQNC4Hj8sCUopQC+ODgXMRhJX
A3Awi00ORUjXLxC5uyU9WDYbEBSEkQ/5iXpE8LU9AXUWBXUBkR2gMlRIDzTz8OlWyEJx+NwvQ9AS
QnYN/sY7W7wV1McvyhohKrpvNmmTr1nr7C5ZUtFqyuLSHh5lky0NvdkOy0gpq3mPYPZH0PnDlb8N
B0MPkmXR0JBnFFphmB8NT1iPAZJpys6hdS0qWrTCLsNnKUScN7hZTDgtAehcNkFbF0p13S0KW9bn
CuN3aadgY9pdJ3v0ecc38DcBWqiwcA1ioN123OY1LigdvQhTUtRZ9XH3vXoKkPNOAWdsMW2SEC8h
1Rqe/6Nczr5Z/hkahEnm8Ej9fgbLq7RFdj+COh2nf0PPUsCWsNheI7o3Kf66DpbRzAW2dFvVpDC0
U5W0YS6jmOVjSnLEfwNiLs12hqQvABY3hjWWWdkmFYVy9i1OZL5v/Vn9sNDtj4rylI/j/Z7ytPTj
uPv5Wa2dmvWybeQFRrcMbsEL1iISLc8Vle9cCGQO3FsA7cZEKEdLGHm3+dwXyTCRv95aSJuabow3
u5W20Hs76MnB+xRYx22pW1OYOHeQ22CbIn6t3CPJ/uF3eEV4Qft+0uVA+v1N7u9/i57gBm5HbrfV
XLT+Fgs6VLVcrcPO2yotgLCjIPcelNGwFkyKw/SqA2PhpZ0+apzeBy+nXGU92Dp1TcPr9PzhIrHB
w71YhxhqaP7uP02PgKkIakXyulKP+wtg0Bpx+y7KRPS4Gw8UrlHOG8U21cpZjuyTKn3rmnRm7eWE
bJnoPslVno0FPr4jhNoseON2clUXwOPMCAKVjgTSxmIf7/IU9rv/Xjg0pHSDdy6xNlnxMIzuMRxa
nf1Afg14oIOaAJje0fybfdxBQksOpJQiLda8GCXud9smyopmT13X7jKhs3mXOi+uXHrz+pUsIK06
GcRbpwFbBo+rc3pr3GhwVLCnaXQ+UQ1ynDSJwjISFNXjMq1ole20Av1VwkXEHW/hnnNNratk4y+i
LmMXOdpvN4HwPYC9zQHbXnZmwN2zN6z8gMmsK96hppIlQNzbnxO3i1wkEKs1vmwJI4sKq947w6xg
js7ygXHztwsDy0h1Fay+MNugj7t3R5EIPbdwmB7A2q7PpVGBfybZHtZegs5lFjO+eZjvoO7aO9B4
5fFlrgRR2Zih1ALn/jSpg7qO7ns7NUL8oDEGFYDcpzwVs8ig81ghj1Jic6VpOXXgbrvbOj7nPxyC
3ZFWaOpKb6zpiQ6osFB2X0rS7vQe/1Jq6eE7804vVXRRL+bo6AMpzMJ81v6Paeg0S9eyVQtc9feA
poSg1vuP1V3Dw512cuuN3s017k6YSc1fhMwwUgX2dXzR7S26n+PWoDxfpAIGZ0/fJBEZ/RGRn3Ie
MXQcU0un4s7LtCFoB2p4Hx71TvsT6InP58f5t3m3B1QUX7gV2jUW90uqkydsNWOoZvdpCtz7r3tj
zMXiySRZjfz3VTY4Qr1BBUnApOc75Za5YkK1OeQCG/lM6ijgu+R653+UNrEXXggVLxW/vgAvWs7G
WXuYxFV/ozkNydjlSO1/Fw7UP4NJBV52Tkcv0+yIll2KFyXxdaNuUOgvvzmEiWKk70cX6a4L4AXD
LnoPI0g0KaKvZa4ezxDIotnm0uO87SiuJjLsbMPYERw//IT+5jQfyWRk46wwz8E7oG9a2Vd7w5l+
TW7tg9ZTJ4f3xtmZM5jx/sNnpUxwbCbmH8GOCu2qFSlYUoM/JcIMQrfpGXizwKDwqTI7t5GCf+Mj
uys2/tT6G1A/HsgQOYUSwKju/oQFTePcjTClYWd4/AUOycy77yN7OlCn6gG16b/SxHb3mMylzWRJ
DZY+bSUkzUt8YuIA27SuTpA6b4AS5oELdkmzNfxmD+s/97gcXB5YEtMETR0tdpVB9jx3h2TOHACI
qm4Fgk0S22tp0F+pGqUqjn23WFDl1rYSZq7Xs5lqMGmS2iJd8aLj0CktvJAsQVgn1XoDeE7OKAXg
pQ6v+VqwzRIiVFfP7r6p0grhHSXcEeFOflqprxICHL71Myh9eMkNSYtzG+dm1AMzfAcz5XbudMMd
tF60vERyUC28vy/w4BhN6791tEx1+Vm6yLj54EHx/8wqtrNPq4RYditxl0PkwJbc+E+ihMWKqWKd
IbAU0VQZUqKucchd+Pwiyea6A8DkzA0VXtO2dg3A1jb3BSyHL13ROG3bhwrZPJ/H5nYhzJ1cdwWo
5ZJ2cqS2F384Sl3NGs6lQjFiegyNFMlSFoLSKnEOrar7QHiYI11YvW5yaORl9tywubfGsc4rMSNL
UUi7/Pd5WKzhqL/FkLIxalvQqaWmue+nNONpAIx2YO9ssID5Gncz43lOD+WS8zJh3dVXGHb3FhsK
xRGlrsK3cGqqtn7nkKOF3qp6E06CkM3uf4rudD8E94l23MDuO9/lOY/O5KP2ddDf4tC9oXzn3qqV
aOeyXoqTIwMs+IrCUn2VUwF7nLa7uCXvpbRh4s6Z1UyRZ8c0RbBThT7seH3LRP15GIYfkzcn8r89
rq/x3Jukld0+EUlmF0nNX67YSMgCtGT0xtt7geiqnh5utkztkWtCv7oDWWVRziW7K7Cyz21V9u5G
KQTTEn9YGv01ImTOj7yTepvFLzh0NoNK49tflYoXkpnmyF/siWhNfL1PE6+63IPPfpai+/NV/Vnj
bHMLYpKpJPMm1fKEAIEwlwsE/YnhBckEHHXB3/WlvrqRlVEDf7HUdNcy9OBY8+4ZPJrdkTzcESoP
nwrg4403GRr4gkD6LNZSS/OWewfe+elLXfvx+f+mBaAhvweNYK0CMjjn1hyfu5ejblDYGOJP5/qz
tqXNmYCawxBGdMKaETYb3yR6kTJSrbA3ehJU2oYCIausRV2Ts23k7eKvHIkBNrNsbGAq0A88B+bA
JYJf5jyBKHXglvmo2F+6NEe5DRuw8s09JlluNYeY17Vrrm6W+HSI/oC5lvF+q7BPgVYmJuAg9pCS
JE2j2/GysDbJn3MBMVqcbNmY3dGZvKKZYZMp0QtGDBFUoRpsd7s0/DyCXoD/LgzvI17xcZe/gIAi
XsLJY77e/VGZDCdxrOXi2anQSpvTvhF0wcDqdeDqx4WcmDPPaiqYs3lILghgVY6uqIvHMWr/qZBw
Oddk0Wn/63aU1sS+AhqTlpbYWca2lbH7UdZclgeofjIMgvMIwKkBFCxuuZ7nW4HPuPRxQkFkJ+g+
9tShWW6e75By0D2PI5eh2FIc+eQ3ujoDLjWvUFFJyUSZNPYY5+pujQIyA1u1lnjcT55dmTUvwdwl
8mNhl/QQj7oeyb0MnzABNNe7sgENC71H0F2Xvl+6CQqxUrWfMk+zwA2H2f3T6CM3Ot+z7o7vKrkN
UoNtXi7vFUWso7JhdHT8AYoZ9CO7d2fS5FziBvx+8UDIaVxNqaSP3x2we7EszMhd8mCaFU++EXrh
108Biq6vwkoGt4VBOcvPG44FI+5AFIWZyI+n+1d4b7cc8sKbbWtsir8nuYjIC04yt3QpEficzap3
bk7upRIDtIvUQDwB2T7q2UdwhAI1KPdBTSYkiN/J9Pd2sgBb0gSFyUl7Zuv8vMJRnRXSLCtt1DEc
L3HkHiUNkiJB6GMeuIGWNEQY0QfYHnsCeehD3I8ss8kh8CuFaOahD70P8gt+ezMN8bSmh1XW4AVu
Ty15vvQDn9kI4APtr9epebih9r4+mONQrC+MEAVBZdkCckqsJEg3Tq3uEYqccFZ5snIHwR3FCJUp
0R3wzVS5rmrefih3Q8vm3J8dBhns1u9yh9ghKvKSJqZkEDvgloLS+JN7z6dY/g+TcZ5uO59mhRcr
EGpZn5K9Esnky47ODhACzG+65m89PuXCyXnikghzNQG4UffF3JLu1YdEW5lFbMyJ7o0NgE1ODk5b
WoqdBhukqZkB0EmULD+dFhIr0KOfQSqvxc/7Jh8udbdqu5XTxdeR0GJ3/RzcAx4XL8JegtMt8ZQ2
t31tHyVoIxQSPfr4Ex4aKtTh03Tln48VExzvWNfTKXdac56xMVs7V55N0AZj4LiqJSoCCN4Y22g/
Vv1zmGYjSN3vgP7tFzcd0RItlLYevNogevWeps/w43HIYOLQFCvqjWAenLjv6eWY/JixGSVbo9A6
mvakKbBKEyIITTMumRhtRJ4dMuc8wg1C51WCvLmsiofCFcF/8vZtjalFNDE5wlZB4lU+P5ga7vjh
3qSsVDbDydxoAzvhCj4FAu0U2qqq3y7mlI/ur636zu/V7OwMXazAeNpkaIzBYVhJ0FdxSOIccQp/
G+eCf+bCKodTfoCfwNzkvVf+HIIblMkobtz1U0SvLd23DO7mUy60T5D5lpdPHR2nAkUnMYkl7c6d
PzOvb+5wvZHgKSlUM/omYOigJF2Vh7TkAxGkudCUX5bU7Mp3NkWIsGobq5zQX/0FXdCenL4P5VdE
GLWxFdqTe0CvxgMjNF2+6ZaaX4h3toBL10dRKOa+q2WmwsANl2581PSw7WlHxdKnVH9dn8bGRzGV
pBKFVxvwU9YY4d0RIdHr88EnWvdNuUKMPd5MHfWATy1NEiUvRcRo2A4ICCHuQaEbTUF5C3CmbFst
Bz9X5a1wZ9U+Z2qPwmDsDL9/+yG8XsUWNCdW78OE/M2O0nXoJovdLqg9sKwdSXMnKTUnWCBkzQjb
n/qTqB2kpkm8pbsXwFaKNza0eI4RjbYfzOpqLnNISG6ztDLFe7xyTe8w7YPSWtxrvXgUXiluai+H
Sk5MHahPehBHpEH4x04DMryYrbY2crzfVG80Ezi4ROVWEqrOQ8/EdH8MpBcTo3E2MV1ysbhv3cH4
Xut5CQHXu6k5Bm9k9VSyv7OyMoGqq7VZKouO7VN4w2ojC/hKDCE2upAruqVUF87M2saphiKBw5E0
MKMUgedzsVJoJy4pXD6ZY2AbSDCdC/UARBD/mODohIj5W8OWwLYHBSRCnIBd96LDfNUYVH56wzDJ
pOP4bQ1F3eKKyl4OPEdxSAOh7GhKF3plf/5f4sKqqcRMecJZ4x4a6vt6XQtH/7uuG9uO2sne8UzT
S+50FEeBcSkn8XWME+ITcC0lAeEcSZJEdGQOabs1YYc6filV8Ye0JV16gBXzgmBDdMYjh3+HQN6F
d1PTxYZCIeZ92KiDCKyc9k9TiGB0zIDJqaaoEl8sqZUVj1aVUfAbB+gEYT+CFHivY1l37yvrGINv
T6kBpj3XahNKsWg30IFRC7Qi0pVwwEPO9Qxbgi+oF5Zk5FWVDqxsdxF3v59I56bLgKmU9rLsBgFp
cah5Q4SmoFtR6vLt0gIs2DZ03iwV8GVbKEZ10riE2e7A6lb7bLCQ1PcbGD15GakbUcOg1UUXXuOY
OOsfGU2lGEhwLJZmb06n/Q4IeQ6Cg9d4/RR8kqJErdulkOI3tvz5E2ZR6MpswyJpwYhZ9GObEN+d
Q3yAJU7w03r8UnuyGUL2PtpOGIGwnI5Xs4vAdDdd+HwdyDzEqPT8WOm1CfpXOha16A26K6cRW0mm
cBdT8q+746qbXWu9/7kM1mSGTke43cB7d/lcpQkmGmXuFi1bwXxy+R4edP7d/rLC0JfG4W+0NSca
pc2gHO43TDfXNZzreCVmmPPiRiXt216D1unA5IaJL3mpRIs1fZrLtNwxHFbqRfEQEWVqSC8oRr/H
56nDgHyMWI4zzDVUNeUjWOd/lmalu4npcqrOuPOcPD/hzeIZKWnxXhRdv1hp8yYFmmBSRHZNEoho
Ah3cgU5JWSuLMDZ0JZkIgjyapaw5vDtjv1dDbKhyYOBB7Bevk++AMLuMlHOBbx24pCYy01r1IxY+
qiuAAofm3uMyiCkrnY6zptgNsADNR7EBomP2NEs3JLSMtjaqUVEhDhlDrvnGDnSvwknn3kQckYJ1
EO0p8b5a7eXbrn5waY3jr7sZjPnRdcPZ5jG/91N+6rRkYDWRQlBjUOlFWUd1Y6YcRk2CG5YyVTPq
7H40Uu1mRjCHZjJJNSXf9ykEBYsqRTnvAd3Bvi8rV/zcOYST7bXocp5lLXt9csi+SjRXAebkr8mC
cRMHlHkFbJxTNUi91JYRHlgBQBvX0cCBZXRnsdqfrpWjQ7rFag92k8HltmADvADjv3ZRQW94t48P
bf/u+ArTEtXMzDH0vwGy+HPFw9ypTF3IxBg3drkVi6I/hUvtAwwEUIcCWUOZLh8cQh3pO5M7qFk5
/sICVY0PJvSI+X0w7inBpeDBnXJGW5OMVqLhPlTGB9Lhgaoh30Y0sZ1mxcb1cxz8z+j8fjND+DWp
MuqFvvlEGVmwnNMsAn19dvqisNWKXw5qyRG4Odp+FNepbyc87O/tVvyf+xSyG1yiARy0hQUPRQUs
ZdRb2GUBoRyQPsXm37nwM2+Sf2eL4MM+AUSzwr43A0echPYOBimUyp49Kfh5QowUmykOzfLGbaZ7
EIZiI7vaF/+TNWdCGKHdHSmrNFgHFW4GBWY5gquMhD7yUi8hM0iCBUj5chaAdqpKw+tl72ICf907
2+MdTCTcz9L+7QlKBSvrs/gPMW2gE677pKfLuWWkr5YnOtyvX+luyosvA0x88+mDCgO2sioL14kQ
O+yu8fi/XmmNSCTaHmtn5ji9MIS8c9F6SHE/dWjb3qXhiL518oqk7GQp08FWlpiHr2vFzawGDzSv
Sn22zT/5sSGxPgA+1KRIebjUjxq2owfXl5vftl0FptLQxTco1dd7COHY5zOAGAeekpgRF262Jgtt
/3a6t0Sasa0mn554uyMb0M/802eNKXcHIiAUCS0v3JKH/KRR8TAQmlfbkFt18NPkCUFq4i0AlAOW
KoLQwI51YHOIMpHp8D9gDzE+zhIrs1yBfQGAyPlS1+13a51/iYPGqaYswbwXl43ECyvm20q0AGFV
Yg7JPMIsHc//cea3I8cbhA/ygdUrExlGUJ3TInKwhOLILAkSRpcSw3CHjjLP619noZwSK1Vq1n6o
/GAMf7ZagzQejCWOCei/CZX4GjNizR2yKOPeCqpOLhHP83XOqFvwXrCLxAmEqRWuvbzWddwOb/ir
E+ecX++7Vyujj6hY+KaSc6HzRD8HEiWng3rCDUADUdXYPuklURPMZpYTxyBncWcW444fXVHYE5Lm
3jFzmnV4TVGH9oyjurQiyqvlkH3MY7PM2L1GZ+7/i2vfsxOw5yaszjwsA5UTfpo7+pt8IOc7zxUN
ZjLSOy0Uc1Oi7XmrxKz22L+48ztFe4VAKFaYjVfyiFtF8ydmfMAK+hgVfLw95RGPhTbFamt4I9Pc
ZGn5L6uAPk24q/CvNnOHmqMFZ+0KYHVEChv+m/+GBQNX5qqBFE3yC0gXbwXd1Rh+Sull5y0hgstq
HkjwOcy87kn3SoEMFzy6viRJG9CSJfmNCHLrCaRDsS4joiz1kfurTC/7l5ahFAT9MUlS5g6JDBVl
0vNKRs9yOA5NhgiDgymq2G2sdsuNS1aUnzq4e48GTbg9lvj3TQIW8F2fVlwm+AEUDcMPbhKk4M4w
bDIfN9YRGi5rhS9OZWLG6J8tiIC8W+FAUr7HIAKs7n+Fl6mPcOFRnFwp4AYHIQqrPKHADOyf8PL3
9XG+GEvPFQjQYGyg4hJc/4QUFCcFewrHOp/dWu3DTubsUy98ux6N7zaa3K7dhFYmwaX+KYOMZfRS
TbWbJth407hWDzRIl7UmXKTA3XWP3QiuW52QBYQt7gx0RfHQLbY67DMDpt2bl2hCYzjG9rGcHQB8
A0YvV9OJKWrmrLgaqmn1TEJto8Hpr8tPNEjLvFY19+CTmc3Lmf61A/5llQGk0BLhob+w6mutZe0A
K8u/6vytX+Od4sQfboB7uBRv14heSlRDytwu5s0MvysBXPpCrM3MkDLArsBBw66mUvZwn4CF7NXE
b+Q2D9sTQNueKkqOPVJj6TkwWw80NxZ9leXSIrSkGn2Y+ZqOsuTTb0NHG+E/0OSSjcV+AnwXPjtw
TBWFYVCn1649b8Jz9qnExgWAIWaNg7C38KkaK3diCVSpiZXehQpZPiRBC9uQK79qN3eKq2nFpt4o
SdGx8p+0fXzAoBH8XocYJLCCdSAc9tTnqNq4W19UJjykJ32+a38zwG+YXyEhmixmoLZK030N/CyC
yQx5FrJy62/a4wkkwILP097KTL+2ufXuta8gvPJgBvDyHuUV8/9BAzJahGnWsOzV2K9oBQZ52vpT
t8oNifnFQ10ZfmrUWuHYf1/oUj5wa48k2cZy/lWnE5Twgn4lxRBpxUN55dmL4+ky1r9ZcqMkJZKz
Peww4wK2lN1hVDhTozpwDQ/++VQot3a5GI476OzHiXejIHdP3WYYreYvlye+C2MGJ5ywHeSafXhD
fVJxDtasDegV/Ki6ciHypA/U5+v6Aiof5FVbcvugbu7IJYWqs3t/pP+aP8OCtMc4Bw8RQ6+uBg2x
NBWUqyuXVONAwzBr+5lrg7SpghKti89D/c4/TKSHkGotC6ZVP2N92vPdzMAjXfOjxTd2WUUiZsng
qqPJug8/wrluVxBmLcPJjiHmpbDi88xMRKNFfzhYDDA2631CU3uvThjr7jVnVDY1/Pn6huQLpwco
2XY/Yfw8djJ5gSiGrWcIOrV7G8UxFdcTn+2Nyuxq0xidWw3KS09NA1oJhLAWpSn2vZR4GzV4azJv
zdXMlWBYOvYeVIOOef2LGX6edmWylAEje7foJ++RBeNGRzNa561X3bQDyHm8O5wIk+jlrKZwR6zO
5yk3gialGM6ClvfgtpHZ1sAU0ItvIDieRn85rrlwB/DDBM8lKrYVzobsjyjVPjqrJMo6Z4jxIynV
JUIXf51Rj4WMvYyOx6GIGUDRptyFHIXEH9cdINHlhzvoxq57qdUy2JeI6d/L8esmcFMd3pKKwMf5
PykdNVD4FGT5WhuRV2rrhGKT7bVKeWAHBnNdR9UxGJeM1VcekBw5+taSjOfVwL7bQ3MJ5l7PfQZJ
viO9QfQIV80bZmFyayDPvE1h6ZKKLl3Wo9Kb3RD6tebEZP+3F3YvYFh5wrvv03EpPF/FjGC+dybR
lbwlEBJHQua2swn+YefKpQNo8KObV6eg5GsEhnJiZdTo4M7+aSnc6+oEDzoffPUvIvNs35x6yeUe
qNNNxvxp+2psr7vc1JSzH0sSQgq4ejEZMOQDRCGpuykYQqLDl2zsYgNbbpkF5xz6nZp29AYVDiNv
mcAyPYfZKvLkcGaVyITUw2+ukVvE+vHo0kWyHNAdRBuM4YUyZv4ywOhB9LSgQmEtaHyYGCpl/rpm
3S4GnNY6hl4vLEpX2a3R2htqrXcnL6342Yb3HqVXTmlHYjK1lqMAZOqnEcY8IMpzsnh7lePYhL7c
yaKNNh4w/CYklBLJ5BOfTHL71LGlj7kvgp2GCJpNBQuXLi5D9xq2dsiKKNIav+IlyKuoobiO2UA7
LpA38kFkQC7+18DWQzHJUNS52nbA05UGcCmRF+0MByLmDgC4jc6DHmIS5vhnnYVjG5uyQSAMSxkc
cn1NvqlwtWplnl3m3Z50YMdIL0kURDr0LhSj8EFB2ePQl6m+RpX59IlmRHJ2HdT38svSoiRHf2sY
juG7WKWu35iXA4VNSwlk4ywg30h1hUeGvTkj9NTyipjBoKkCYh7DK+8hkFDKb7LR8dBPc96c/zBu
pkG9GnY3SZzhj38XAU8VQFoJrPrXloML9vU21Oy1zmjQ9c1ewOvT/E9r8XY4zGMWNHwfdQzRr+xg
vkpF7ewk/mHVnMbhMZZSx96QIs1MN0Go5XZyp857KTFIA4fLJ9I5xSae+NDIIPzKcIszbdJSwhir
9HhcLJGaZcGaoZUikQp6s4LjtK4pDJdYakCC0hXbnyP5ZpAxuwxvOTTvPXXuPqh1IXMHP+eN/ARo
TwHOdTuHnJ1gTLMrA1A75ujzp8K1D0TuVcFet/9lZflG3yhBLlFkCrpMkZpnwghiRZJKMorGWt6H
Lz3iRyy0o0feM0NLEMPbzLqANfxRaY1XzcJ89IMrYyNFUI0oNRA7ccO4xNnuHXsZsZnbwWm+7+mh
6mQJ0TDEZEPPX8HCRZVvOuxDWjm/wu6ffHXIbJptEAbHBVbywpmTM5wqaVrlUH/Cd81OkhzBSPD0
6fDPSihq70QFvY6HiGrfksvD9zf/top/L67OnZRzC52o228y3cVlo71atmp/fWZ2SBDOHwlNQMWE
gLFwCMGQaqLMHCHXLnkGa//4wvepzoBFE4Z4skhkkK0Rf5UwS/Reg1iu8oQYpLaezcDWvGMG0sHb
CRNLUCjMW74pOeVrBMWar+PTDgs1abNf0RleMuwNxNmMxs5hdGxABucL3BjLHxxr3lYLvOFdVq9w
MT4cBC2QFz8rqcLvqz4ZXVTOksGQZ4SNRh/RWfDLGXq7FyUfA2NMi1YKezKTWgJqqRZofpPEGTiK
Su3dsq1UleNhIfRURFsBVpNP6oFGxJIL7DSc9wXCL2BldIDaIcDFhAGm8+K1T7NxIHtP8tI3Kw+/
ESZVjWkCozkGDRitzc0NQPXCEjesrvWL5ESc1DGNa8oUn9ZSp7LDeAQzaYsYrI39PLkl95PQMRLc
dZ1dV7OBpnYiMuuTqF3Ru0DgtbZVKaTBSIEPD3B7X3dF5AQ+ELViVrh9blv7XSGZacVxC5V+SDxk
pGevmxz6g5uieLjAs2UwGfQ5wsWPMw7ULTAEfwzWfHthf2mJXzYzGvEtJUyfRpjORVWOOIhM/YIS
XnTORTIrYE1JM35/H4s2FfxPI7yr5dTgROIk5CgV7ArNcgmDqhV89khcSm1oinnQB/8m0agAmmu5
SqEJsWnMIVRIHL/fmDcZeK4AVl6cjzGXpnlg5yWC6H9JIImzprAh31gDe8AQ4ez1DKNb0NqLLHqK
vPWLnXoClMWMmdN6C1W5vIuh3Y56+N21N0riiP7KjlMfLCVbHaL75Tcgp3x/WlQEGx0MFgH7NzZ6
8LbOYE6P0Ev06htbhjQCa9hbpnYKkKonNrc0VUV3d+dsK3dyNuUZglSTC40M9aTsffETEZeaMuay
k4qBRLlgmgtJnsI/CC4rJRGfSjYzP76GsEmxNFfdDC/e4mb67EdpQwUWLlwcGpuVoUouFWcndtmr
7z1JxEScJLYxGQH1VJC7VtUybXGUfJKLJB0H6zH3okH8jltK5C4xJRuID0Cy6BnbHcYwHFd93vby
rYM1pMVlS3PQIHqj6zVkPDLUGFDZTEm0EzAWGTJ9y8neElVYR9haQ2V8hA4KkO7CgRAdmE4DLLvW
JntSHLEEWUxCHfhDvqLCjA7iKwBcVO/Tw9333rshP/CpJM30Qvknw1t2xjut3xG7oHBOacPCjuDa
5zLjes9ZeP1x7KjtQiPubnQbZYZZzssShnryA1BFvYAMWqm5RC0smtj6SRRhQOWZa8XD4YNsc83a
8BSna5IMdICPHk3VNu6moLhFNh8avo0sZ+9zakE+N+0Prd7rHX3O0/vSUxfGzsEqEJ6F9eLnzsMP
bb1TPuCq/wnHREHdUAK80CRZi6Pf66uWP8S3tIZ/CRZsh9POwbzldt8T9Dn0oA0C9nIsCNadVDVp
LW/GmMzcMjHTxuTrgMMCKZ2In6qzQq/MeqPRpUzD49F4cr6wSTgsHvF/zZ9KZtIIfta2MQp/Kzb6
53d6quS3+BRjYyV0vU8baalPbEy1dQELZZlw8ODEYuMZUtDaaallfOBFKhDHpeizmYSUdN3plCp1
Yr98E/Y19MN0EbP/b6zbiPAoCy+3lq8HiKJUoWLM1Jf+o7qDz8g9vljdgtkPNwsoRJpyXFyCNeYt
SVtR4bTyLQZ3ntysmhCmJC7/r6+VHhuIIxKa8YlipM7pWAZBfy8gGXAQdaA9vzEkvQWxlDWeFy28
MsFARWTBg/EKeWfJ84FAOoWrCq+W2upcYtERJbdrO+BNjlug5qnbIEkltnUtbJTB7OgUDWGnm1ZC
mX6h+wEBSE6QyyinLLTK3f3lElLEKPE+QAa08LBXygZ7PndBvMo9g/kl6BnLPZLbYQ++a2lhv11/
hCSKyyjwrtnhgUo2qETjgguDcWCOza1Hg8Ay7/AYiBhcxKjRW0Ysdo1fuMmV1ygvj+9owln/G9mI
/1QgAzsNwYQzYOM631fyvlZx9FJpTIE2SnNw8GywmV6sxdVeezop+duAj/LI/MDQq+UtuTNcfr9k
92rAJuZmcODWf2GKrSQdFRsh/qQb23wpvqNZB5ou7rzrI0UrlsZVqrRcFDGgzag9crI/hVYX1SDI
3/H0hNaPX1SKQZzvfuXbgwdqbF5v/IIKj9FyHZfTD9VW6Iko7PMTJy5h/cvy+Xt+sJDgrdjJkHsb
e2uJDMd3J06xQlHavpGCscklSXx5Mim3Rivcm8ChFoy9v7RynWpT8NCK0cfk4xRj180qxWOUMcd9
VHZGGJ2xrkFumx2MAmzHnJ5VcasJbL/yYAt4EDA1NON2cPrx71VpD+4C7Yu9S6loEwSPEhwy5ax7
2yXvfL2JKXZ5A8BbDMrs7QMigLvun3S8pgTEvfXxrA6XsDvoHflzTcxelC6xKJbzjYG/62LFR07X
hUPO0uzWtnvWzUiBSrSCDG4c0fJqGBZ2SOg7N3ws3YTLmOxPnBXp9XKF9elLAaJixojL4hlxOaDq
xeeQ40ITrSDWAT9vpEb47L107q/QMvT+rrFmebSqvwNLFN6qRxHR7LdnptncbFUR2Qy13UmosZBH
iKYxJK7FUqLsQW786xMqjtLd0iQST2476fYIKEuLAAhjtWg+YjSWGG4R1CXYL2PTSxCp8gYvotL9
HV4irmeQ9IwhksSE3w+hhrKyzLghPAaZFdCMGfrLhjDYabS0ug9jsU7wNrvxDyU97t8iVKQKEXjc
sQj0aZiPfz2V/bVxofw1aBniiMPxjxu8s73G+FpT0S2zLUV/hCbbhkPfi17Ao8VPiCD81gli4jg4
01bej9O0qaN8gGkOVXVfZJPi2tG8xAv8CfUWogTaQnwZQOKEjnvWkNktClMHWZWE/NUshpjI4VkB
QniRD37f6BpzsPMrYQWGTxyekOa8PZjcr3O3f0mKfuZOztunzFgUPQWTXiIIPrBQoXwxzxW1f1V7
T6cL6PJuI3cn5Y/7JjVvZy5xTJYHAPZs8wMDss63RaqCvwN1r9JBEaDdpqMp3yTdUf01YmwnVMyB
iesYZ2Qq+LyeIBa7CLIu33MXPAJwDQgLhVhNAOM4saseKXQmdacp23/8/TU/Nzyz1cusJ0p2RksX
twyYU7lHFOEDLsyljFCParFlukceVe1kF1BqV9NtiM8UAhU9Fj5EkFu5BTWAfSoNDbY1G7zqljcr
8AtTsRNQtjrGBgd6gzDHI3esIxRepKWOJCUS0XPS5oaQ4SC29VZOOvpQEocsWGgGNQjjAhzP004R
kXKX1UCyxuGlgd+DLDmCO5HI9UtCff+Ukby9+tCUZSBTBN4a2Tn8WJLkNo+/eWcj9cpmQ6cLyt3y
OCZV+KXnY8mDOOCKaZeLY3LLwNvLRVJjJzOS+YjVTipV1T5xya0/DrQsN9xQ1BSuh5TBi3t1gFa6
88LI8naFFudlf14gghdybfvmP/ZykycZXU1N8r5xU4Q1zW7SlWYk9DLji9q0oNX1YGjY9q0p23rH
tErnw4GMq6S8UiE2fsT+LNeJ50U6p6dxf8eAspKcon7jd0CRDqohb9wqAEuyrFsCyxY8d1tYBS91
Vjkdy72rD2nAYjTfgDQdq3hYUVca9/B/8h1z2XHjX9Op+Oek2vkSfPlaoAZmJb/OkUTDsULPgkr2
4fmpJrONzKwHdgjXU/i4yYEA5d4afRizcvjRpdlkJcppd/j7FWFS/eOa6mer63L31bu6xs4GWJ2s
dpoZLqTj1+cuKe58IALeG+DFUlwogJd+ljpDsPrx0okwWj68Trf+hTdd0gM8Cv0XZoHZtqIZKmkC
izeOgAXmgNot7P1Aiw4dzdsup1D5Y8eXdu5ReqnQwoUZY4cVtzVg2+dRx8sabgjv7HNlPdOJ4zRD
4ChPLlfKeNlh0jKWNnHd5QyEooccfysStFQ12eYsfFEZ9SZBEBZgkCczMesjcOguApjfK1QrZTTN
h0ux+or89Ftl6/5kU17mjgQeUDwgwB2uZBfOvfJ4kCZMSAlJ1XdzP4SD3C/PhK2JNmmoXFSj31+z
zYY/XMzbYBw1JvkUN/PW4zz8KE5swAuGgC09YTABuA+utjMUjQw928nXpXcLi76pxN3UMZoqlQPO
+1FW+PYfiFhA6FOx2NVdV8FaOGVTNtL1WMZSs7hEb2ujBAAAD/xsMNJY1+uRWLCsnS/zU2zm3q22
ubT16ATQqca1tJuhTtCccRyJeDqePH1D4yMK66rx60ZmT9GJD8lGay6133UEXYDh33DZuU59+nbI
zJwFxp6Lbp5R1Te//fcgS3WfGuWr82zxrGmJeWhw9s3EAAMGJoqABg+rbNCtCoFeLW7tDnwkcGbn
29IbwDzRmL606FmRtxRSM2V1B8W2NNzJAJQLnIToFgDLjW97gHnE8VO6FqMeVUD5ZuGPOE5hRUl+
30D1aEaDjoS8vIZio1G+dTkHfNT1CE0ryn6EP7+lw92XtHh7R1AfL3FN+qucjDIjLhhSeQveL3xR
r4VLnkQUBhhz8d1o+cCuEnJxdxcizgMew9kA72rPfhxx0Al8ysSFKNnXulI8tiTiKe7qyJkVAzIa
nNIpW4Mrul3s49WRVYu/jxpeiRgU2gVO5jiH+fZNTbAQmacNwLNHTlvkTH58B7voassGMzhyVysA
2YQ6xVhgnhenHm4rg0L/ETvo2bu/5tWshciKsGrS15PbGjky5+Akv47hwmVSebFwI46Mae/dKmg3
sZI2dyBkYiTyWCrdiI8eJiEe+F3TyaoH8c2AF8VB7KRbiyB2pTxMIWxvlSxmy3phABmOMAJQfRmH
s8Fjdxupsl713v8bRyiFJRdMyEn1FFemWQi/m8tNH/CRJ/+GFnQCgY0wH1dOPlsd7A8p51K4ckph
29ET4oF/QQryGplDKlu+lKodWU2lXUvMJVzIf/F7OW54IODGQdvyF7xKM2yC9b5Vl5Iv7yc/8ILm
2PWfOXF0GBiN1oSH9205tdVFYa7UQ8K+zijseZ7n92lEgrDKjF8nrvKoLFMd7e27R9mNMBqC/B9Z
36F3hZz3/EnY1MNi+XtM0stukMe5+1lOm0rUA9odg4gtygdlt7AW0Vrl3eAPMQjKxB5Sg/4nbU9r
8MeWip6b37ft9soVisBJbYzEqN8qThKizhnk8JpbtchFfAI9V9kAI+gy5LZwGPlQz8geF9gsN4ll
qLrUoqU+I6/cOL8SEJ/B4rT16sd71TaOv88FCGF1IyejBIsIgUbKiGq/0aPJCqNJxuXlsptk4RJ8
iTNGvCbX80vty0sishE01G6eqXfSlEdQ2axkzi4pb3iIBiQMK1SkN9FLKJSIM+ps3jtWDs7tDCSc
TdXtd6bNEeJ+X5OXJvVNIBDDrxjRYR/VZBmXE3XHJjwF9go6ZZMtcr0qsyf1QmdJMy3ZXpkNAWVp
qaWQN4K6NzfHfQ+4b4PCfy82vbkO+pnIFA5mVDRzDXdnqzhc9EnsXTIK81HRhjzYh++dspLtDmEC
C41AWgXy2zbhP8JhoBjUKdGb4wo08RhKIT7N6GqV7pPPziPUtaaCJ4YvB6+DLg9/61NAQTn/RfMT
1yp7U9M0V7R08oq2akXbOiRzAr7tI3WslWEoWx3hsZ/n4z/7wd6IMVi4q1eU165cUFVsqjJjGtBp
zitF90+Rc8fsJSKHbwCuO9UvC7zf5L+rxBl6cEE6QuJQb3adKlBhU2EbXIl1HZV1taS0QmUTVrgf
ymoRzdPPeA+D6OulLiZmyDTZXErQIX9sZHfpT/ZDstP81k7wBHAuqU85h9insP3ZSdsCbaRc8SHh
711RZmiVSJJGv9I+nb0CEleaSUDUkVEuoyWU3dpN5uwI75t6uIuAOf6hlRMzAJpen9lJVmePFZMc
jEt/t5Gm2K26MxtZLCxydEfkVluY7K84Al6IuNKFKWkbEWyDksnH0vTJkBKoB7O1fBjQipCto0Ej
texQAgUuGTc5yYjfN/SdahzswlKZNvZGngb7jhL+0EAjlVUo23mAkFYQSjoRyBO0Qfm/1uMk+bUD
1jfjDD9btEn7dvgS+HGNC+saemNHrLYSBTtUySoYWDNguZKYevV7QaVUWp8y64aKDdbvQaf4YJJb
15ZuRxO6qarKqYPHrWbsc6kH3vkVEdnDeDjL+/9pV9mxLUPUGCjROXyYHdj+8GHkfBJMzUUA7pIo
o6vF5oadrs8vVOfhkboc3HRmgeCH6QhrUNoNGLKDTH+yIq/udw7rhy+NikDkPosyO/Q2MKJtRrXv
X14MJH4a/zAJImL8nc81DxMTAUHmnVGZsuKNV+6ZNLJZJOCakg1Dj70YPE3wH5AyYBasdiG7XCHr
R5lakKI3/Yqbadoe/N9SCjlsdv9RloJXd1F0W1Zxe1NOoAg32+yuse0xbAYiz9KRfYow4A+W/zCX
jVGZqSozlMabc9RJWQERG3X0y+7h8ExWoGreKxh1q2v67+LgPdt+lw1vO4bz/oV5IESSFwP6l9WI
gnBGeqbngFHoFk7pcn5LNRFMTSqcOmRuNz2QvWp06Pu2FoYiqNjM5O3cuV6RKZNxxwSzN2wUuzh6
PLZoKhth0qd++DrwiJk0o8Ef3Wwkmsi4iAtCtJvDvfLpczXq1srE90Di6r4rIAeNqd8hP4BYhW+5
gl/h4lOmdNgFWTq+61E0/v0svHxnZs4FrJ9di+C+CVnEXZgqucEbDEf+Lff8LtGxSJw9HFhvgExQ
0+8aVFr9GvAKW7201R/O3kI/2xrDWwGEhfd9M5h+vjQ7Ai0fgo8irHhGOy7hvJJpOH4+odn9NMcd
7mEsYqVPp1fceXzly+cEmdDkOJPxzwTZR+xv1Da+6FxrNM8WCIZ4hak1y/VCvnmDr764ETWDt9x5
s6qtCQaVMqpxehZTSKj5wnY/mYU5WAWMGHRgAJFkhhAuNSjkDtils6ApC/vo43UL6Kar4LKrj9eB
/HoS8k98ak43rSIS4qw86nMeQXTMXJUgI5xOU3TLqgTu0VSYykffG3wJg0CYf0dw4RylB1zSLkQN
p49UVxNv+4+44R3hSRZ3b/IxqfsAK+LOmG7D2HjVw8cqqjFRQ8DsZLu+x770cw2WpFbVZwtO3YIn
u4j63dFCkTcMpLO5KGULG9R8UcYpSziUHG8NyFwSaKR7PoybOEy3nGvfXckHrSkJhBbIjx9C62ws
tCmVJdX0mfVHEUHcXk2tKFCuW0q3U7/rZaqSfiUuaBdphbYD+qpmHc1dJPtIVoyR7+sZCfeFy8Oa
TTG6UDbpQxmVT4B2Mp+6Q/UzFbon93AmlTbMr5bqrrZEerDAQXN/sOXfuCj7cTz9agy6ljbIlxeU
LJyz/s2BmWAjc/+/6cZkRJYZeTjKdnaYn9Skx+ryn35+n4FB25xzbj7R0ddBAsD8vKd+zb5uqPub
Ji4qXXODLmiDFmNZ9xV5E8OczC8ednIZ7FqlupDZjP0wjC3AG75K0Mmi/DgqMpxi/WBZ2WNXO7ds
xpT5yML0kqqS08uBIMr2m5WA/s8bxsnIRpe41Vz8eZH8gg93IIR1wuOENSSB0G6VCD0C94Pe9Xhm
B9YF2SmNSj5P1YLTGpQ/x0vWDfArR1SHn3I2iSY1Z0PbtgS/dKAKoJS7yA3SJGcsBcO5GbYq7H3M
JuW0OhdbWj7JvefLRSnx6+KUlIv0T59MHyCCJ5rObuWgGvTWhyHrOTbIpjYEeI1nYaByFb9ePe+P
DjOCq0vvdljZcCGE2B6W0ffVF9lbZ6PzPg6c2sfUo/RB1pqD7pUA/JNoOS+3jhYIrMtPz3NGZUch
pC+7Qh2m6yNmSt85Mr58B3FKXmeBqdLj9l2T695JOiQXpG0N3VskIO11KAg4e/+WUm56+vYydJy/
bMkF8vh1wDHquG6cZzSYsp80f56XutVVqX/Wun/zs+Zq4G0YhuuhZdelVqw3a/C5fs+25oWjD00J
bQtM3hPlR+md6ed+PzwkvotZIlDRZCWU8RMv1n0/mrEF1JJStcX5uSet0jg/XNVF5JYjCjywpt7v
UYeKsfNlS8EEefWVS0Mp+gjBpIHJaMSDqwZQpzwIwAVGgH9vF88GKt4MJJlwBG1B4SkSYhU+5Q7k
6qK+HNpq93pR60NiwtyqcwZAFoYjix4uNS7QJxxhkkybfB9C6yFqmFIU8NVsnGkfXgZof1pjgiQc
+0Xvwbm/UXxb0r6n+hntkuDhB37y0FrRgyjTTRvt5ng/Ouw0IPXLwikQ458g/RLxQR3IYT6ZU3Id
j+GgB8bXjKiIOqxm3tLWnrm+0mlcCPNlC7Wfj5tQogQ9ulLhU87NFOv4lHBVdlo7q0/9GWAQ+jYc
CgNttKshU0tT2C9GsrJ+hrD5BiJC/ayx0LkpwnrQVRW4fbKwHtH/JLD7qRnV0wrXqIDPxLz99JXO
43o/zqczpbBv7oJy8fywubPlmkWZwVNhyAztFDxorsNQ27KhNMNou/UIhibWAhm6f3u7pY1dUxNS
06tU/HLzhSycksMPoh4JpTjUIdU8dx39j++/MeIAJoT9+XSUCtZip6/iD4RBPhbW2NSN2f81S47R
y8owunNqwosxn6ZzNQKZcmmcFZlLKcKVQu2VVrcTKyTR44r+SUbsYyj/TAgMsjL9hkpjVSUC7rgY
5tppMGKFNviHf7dtBsSMtwzMNTqC/G+D05meCW4RDCnrB2aPv9NqqSuL2xhy/EtpfHaS4NCCHl8Y
VyrzzL6qJrL/Iyz9mJowlTbomyC1XBr6rzJdPwDnEdpWoRdSdQvgotqLX4/H371PKn0/ahEhUFX+
N1c0kSL/fpuiDXYhb2fIBOWbpZX5mdVNSCgn6j38vq1eFpfayHulQV20dPkeKqTJDfzbEiH/gcnE
Gs8sbEcMLhxb8qkFYvlPzTiKCZV/mgtYDkHR2btDekxnqxcKyxS5Bjl/LSwRr1UroHD09PQaU2Td
1gvUYYAotkcldF0U9bDudrns8Qo2M8I2vEnw59zstsjz9mJ4K740QjYqCic8oBGLJZhMVtDR4jjb
conivcRxF/pjpdIM0YwTVXd8wBKCAuErM0xux/MhQRfQpHlBqT0aaLW3ovgn5470Xbq7dCKKeqWu
+Y7rDjaH5+lqu/X8Or+nsqOvkGKGq3snOGe/0SQuzzrh2C+7tGQ988gxUxsJopxtw5PHy10lrpeS
yjzlLrPXDuNBZhlb3lYWqTyghtUhB6aFupRen6qiY05Iw6m62E/UPewAV3mtSzLx1uKO3QGvhy0T
s2CSxIaP26cR6ccULoxYUe1bVbwL/aMwedh46BLvbUiS79weD2ZZwbovoepVYMHp+w5/J2f3qrrl
ySrW8D0Nhd2l1+iCu+ZulnQMdsIN56vGg0zZMjetVgmCmKEUYu1H+dOETP4BNkI2alsQM391I+q5
/zcEeLrvd/00w3Jylo2f+2lnWBb8f0i+TEBCY2zr4QR6ZJEvR6gYHCFll6oD0rUFiGIdDC/6LB8c
9JuQPWFXRMmrtkOYyTRHND9k2UjswymaiJpn9fsqrtup6AzWA0ZL3niIUwlcmTWTYqChddHpiJLm
GsjVuJiDqHZS2wfdEUVmD2kpKKpjWqmcIInL1E794qxtcwNHWWIHqL6oDYHIU7JR/7ei3YOTybkE
mummPfm+V5wBktEV0NGawBDBcqvcY9t6qs1yNwuKXD6MqV2n19Ohe8LXmPFSJ92JH8W5huE4am9k
qT5bmdu6cVzYfy9GNNFCvZSMyfziHN491pW9YiGS+89ka9fWJ7YHYF5sHr47MECG65oMtkFDCY1x
fal5vHBe1CJz79YpNcxfHrPEtuHAPOubQoO/hD2qXR5KC1W+4s1Q6z078AZqpZaO6zuPNtpLcMRU
KZ0gIouGlcTyrYhg4K0+e+M+l2y38ywwKClVOHVrkMdJ1uW/OTPKmvwnM9tMcyIpluHWTP8CFYdd
/+7o/Fc8aebCFPCjTqCQj+/DO5RJKeFBcCWHPY3SqalAw3KFX9BMbk9uJiwtZrb04MXMn5myPMYK
KoV0cP+6n78GR9ksw6cYDVmOirJgBdl+26B+5srCy8i5sx+do4DEihYSZXEd4qwl2icRieHp39RM
ENmptiQ0EMV75xqXQCxwlVGcplP0hM4KVbJEm8WPzYTE5+8mefN5vMek0OTDPVHKEII3M5H1CDWE
Wy4LFi2IyXIdCMK6hSvkMUMpXI6XOt2c+NqBU5menLwGIsIInwr/sx06V77O/tMb2g7fJI5U+UJe
ycz3MK3vaTMfBLJtAasSqm6iSNVWAGhnOTFLuyAjMX6xix+DS+BcEQotucvHasxtTWJ2RAL/Rtdc
1DZRFbB/rqi2a3KG33WX73UDZAVLVHXB+jANMlmJXG3QDoLVZs/RQzAOGVSgYGduEv+VGYAQjMIG
CTpkpWarhmofaX2FeprVy/XQC1/juvkuraf1Bdx4XpMLcO770NVRF56DVNDtaG2teAEkZLJaO50h
a/SBGiqa4cWhhsZtAAb7YUGg/GE314fyL/QzKLNHQC0UpAe30pNyOgnKQ7voeUbYB0cCuZ0O6FXu
pfhUP4Cq9dHEYI/sauEJ9qXdar2ljjVmnHe00922ZXy2/uxCEqLw0hJLIrQYz6Y6JxdkFC59Q0bG
z2A6aIscCHmGou4gpPdB0riKDriFv2dLfR5UskrkxWI4vLa33WdWEnrYSUribvx70bw9fvQbaHm3
TUsrXFaiP+FA8li8JcW7rTNZqAWJkp82nDh1qkvQcMmZQZeuP5iyNj8nRXF7ZVhJNkU3PFDn4Axj
Pzn4C3yHyBaYa2sRatk2cIkYcVff1+D4pb+YIf4FQwyyVz8qbu3OczHOvFUbtMZMbdKRW5d/G0sn
c/sEw0ke5svb1/cWGNucFSh5SAEdmJeCCXjgfB10O2te4sPUzi7b/PpWrnD5tR3sy7ZE0FFOdcvM
oKIcksmv4ZzmT+7WTCH0oSeLAIqXn0GFI7FWiS7Ypo8U+Mv4CbjSXjvF3tzfMOJHVv6bFOlBmcO8
OIjEmUJrx9DZXT+qqm4K6rbUEmh6436plqhi7ZH/5aCgtCZ0puzpb24tgWlsoMdEPp6ro+ahf5gP
iRbMc7LG56qBzOiD3WxoiTJs2sPC/3fwtPjuxiGn397oYxAXIBW0L9fdWDJ3Bg2+ncLHz/1sknNB
dw/hVpjwipex1XLZ8/rP/JCondk4kmS/1OB++jBrs0e327nzdg0rJ1FRsud/NfpiI0GEmTFkRLiR
Uq1DDTLxqfNj6Ubt2nhN+ufLnCpa0ZJDLS3gf1jI1FO6WxRNbCeH/mKZvGFvaop3Evz7w7LeFhAH
4JCfPr6ukdQvfDaMT9DsGJHT8MOHV8cFAj7YpSUvMqftx1TdtCRo12FzrdBPQNjz/QRc+ia846xp
5d2Ii/wrRnAoFfI41RsYEROd21ObT3t+qnXNVo1PiXgO8BIsTXXo4Y4xcpyKPqCqFLr955Jrnv3Y
Pbnu8oKIflnOrS+Q1U14xtU1I8x/+9lPQKmQftL57aFONEbsNuLOC/S/XmtDacpXtablLvOlQVdT
AV4qw0wVYjo7rL93aspILO1e7jc+1bhcjH5S4E6z+qyYrOel2FIyUMgHaATpioShSvQKVVpt+oOI
uFDS96RNQTRx+KkcxE6Q2jubq5ANtfDbsXVc2lufAo55ud/IyIPFFz6J3KH+guDRJzZJixqzX0xq
Ey+Wz0ok+X2VBIsYjeHza1e11OAGokrml9WGcZuFI4j1GAjk/uCpMwvjlYAlG8oBrdaNJC/iGHR4
+a7+pZO7WTpKZL/DfbosoKKL8C0ST661zYzD5G2LaiI7jH9Bg+3H7AclFsMpuWn12szsogGmNuYs
RlPCI6iwEstYORbmc7v0F/TCug5wTUSan9lWX7NFh3c0I7kxlehHyg7YzUHp0xl7SAuImPsmto22
17mJhAChPIaO0lPEgYeu/Gx1GuEReixG1oa20Hblk1tXCYm0/C8h9AvMxZLj4L9FJXmpTKeGUMe6
LEaSCzWUr2Xqtwyq1AL5lniGLW80asPnrqBA3N+lay/T++noRy3w0aHn9g7onpZa8LeA9lrOJRaN
/asJz8WVXWjTs+eWmwaaQgyu628kOi6+K+kWULLlSawC/v/xag4AQw0Emr7WDUeEawObeaewnoiz
8bUpbs8Hgns70j9OhwTLDoU+mSiYBZNWtk7lUgebYlrILCyA1s8UVti3laeQ6D4b/8MPED41hdiF
xZBUYILwnDjuQHsqoO91tWV8oCWO1NGRZhzhzFg85KoEnRNpmJ6efdNrTqA5Fw9pUI7Tdt760Acz
ofsHpK3gvkd2W8ObXCO+fZmeMZCRKK49/YdIecqW8oH9Kf/L9QhsU4107ud7I9bNOr7PzvDLTyrI
hPFWCla3AfxOzPJm85gf4lG2JMWJFb5tWMK8gyx8HRCjbzALVm/CPN/OjsheWsVipu4C2+jHnXY+
8QJz1QPQgTBY7HJUoRr2/THQhvAOCtrie16ZrwsKqza7+tVd2PaGT+98bhw2Muui+G6fXxgVxEhq
yNwyRifuCfZz7mmAljOOg8XK+LSI78HANUjhHmO+lKXAtkcOlM6+urF5Q/6DH5/nX6lMOcQLqSzI
/anNxVull8yVQF+LDHVyriMl4bXq+9SyqyS/Az9z3CwGz5axMS73busIBnBNFInpNUk73TQkp+SM
U8ORQgM0mZuHCNNMwlxQXk8tdTRkXbv66otlsDhwLffMQmmOZKTmOtv55NQC+mtWco5B6EUOS0cQ
47x4ElRdq286ju3dKoZLI5Vdqpck7mhyq6mD3ZHw/wPgQgZ2b9t3da6o3f5W6qetdxe9Q+9CfPxt
9/1qMwt1BcGj5rZhR2xtf4zNXI8Y+rK7kmHtrJcceNKUrkHKAPHgyA6e9lf4cwJsvStiAe+LuPR4
kg/QcUpGhJM/VGSWkbrmsuzsVKtxxCaQgX9j+BjjWhc08ICwbVCIy9Au6wKI8aMgeyovkue5h29e
XYHN9pUVugYmVF2ARsie+BlhXa/a/w3AOhhwjQaSON74MkHBM2aizhczMiyzQjEbBlMRe8ZfKqMy
xTX/C+TuyBQ+u2/iSP3IF9ZvK7TON3/e7KmfO5+3pEReVJ5P3wfVwDCgmuvC5O0zdi5xV+6gulaV
d8bFHVl1N1vEbe94ExxPy0SRWUV7vP9s63K9UNCDm20qLRzVw6mFQDjpZKg3U/AG/ub7DoQ0dI6s
CUAv8aduWRh9/Zpclxf2QKZwYWHsD3IxoC+1i7MSyYCxZiGnncxHyTp/gG71wz1W7x31qT6DftQ2
7C95T9HtbJ4zhnlnmAdmy68dzmkMauGuuRC6hsdB0IPXA7IQrSuAsOHTumOPkKC0VmE/ThIJoBeh
BlKsmBZHcI5pH+00d43P/Ob3QBhf/Df4ya+TIZzhCVR5hVWR4NWiNiuiUS6bG2A8h5vBsHeYIQIR
Ld3O/yC0Oksh9oXjHSIvlDfgv9Ko1VDtWB1S0V3HB5FKzZ45zFB58WYGXLJsZ7jMvOYca6WODs+i
iCUvoWt8gSXdT0QpMTugRMXDBcvcRQWwR/TlGSdABDcvvvr97/IElRzT7b6WpKl2dLATIYnVHNSn
WALK4kMWpeK7N+GaKEnIReopPASPbQ/II3jXtlUxwKtt2aJAqhWnQzt9QmDGGRAwWTsSXKICcWE5
xH89bMJhpQ4qs/6VJ9Tw52QgWAvUZoItuXyreLeG2PCNHF7FbSysrLFad2mSnRaKK+18U/7UmnNF
1m8txtufRAGs647pqD5hItx2COeSrftbcJk3dlGmS3IInpj5zNdbY8cP+gLvprhBW+U5nNeZyvnn
5x4Nz03poz8dRIr69Z9Mbyt84jHgoB653ZksQio3r+VD+xkJfirH07GjmhvXKq1AZ0ieahBW1BHz
x4NXSjMJEVFONGcuLwP+9SfFlACNbCXMQPnIXgAMI3mDvgaLT3ftxbYmjMjCzeYB8KMBTPw7iCSw
yuEckKDzUVq0sCVX92VMG4DDPx4sG0ei1rMqquOnuITs33NMdWl4qZ+h2JsPRVETWit0fXDqGv7p
Z0geVquQ4pwfA+WwCcNOiCX2G80zpjvEzN30eFoVi40EpDctrNHcpFEkd1YDNg/IFwPgUzRDvUfB
9Vm9LTZJdzkM52EULVeshw2CVzy9dRSCmn/FjBdtFMbPYKW8Wu0B9g2842U18X40IHw1ATcbOHKx
PfL3nPFTrsZp66DL5w2nHfXAzigFZZqUyNHvO5zBamQUEtheTtV6F2bb2vbAdN961nqgX5yWxiM4
jJ9YTIvzUaG6B2FL1snGtZVr7tYBHsAyKd6OwrFlycyxJjGjdvys4oOt8uXl5vqRF5jZ6xXGIt8C
5MzMkEBGF0ZIpPe9xFml2AJyuCMW9yay3Ba2wEwFw4iU7+YdguM4ZS+A7XsmYiKcyDruiTHn45U3
ctZAxdf1yrKW7QE0qrU8Dn+ZmHDD99eEugnZ+2zmi9f2iQelzTLzvRGZ9BQtWsuKo+QDBKDg2DEf
EFy2qy3lNfM3VMwW7nsSpLHEIf3rnRJHD5AChEN5z5R+u72HjStUh9und4kFic5R7+sSXbjUQLf3
1tDlpGoFiG6OFAywIoP0QEHEIanFvXSOfFnPx5Pyr71shx4QsNFiAmfM4+pyQk2BohpwQM1TXs9n
Jx349TKhPsBXwzfnMEFrmXUImaW27DAIgERGmr2NWbh/DI6GiUvEFLJbGehUbwons4kh9oe74mhZ
bNa3R/QfPp51nuHIysvtadEYx9Sqoi0+jdA7WpiJOZSIWg7oR8dfL2LbocSgvOE6uZtL2WGq2sPl
DULT5XjdpcCoYArSSDqEcrbyoKa8iPxSA29NEfc/D0gSpA1Rd+AvAZlrHsycFa+M2zb0ZQGorjRC
Odn+KzFFmS7/eR+IXu7ixk/xvUJaUybeYTLfc2L7i68zK2NamQ04PYnK1itzUo/3RdeSfA1V8iV+
fIWkkapKvewSjA79QPLiZXux27mSagdTTokInp8Zxip/2Hfjkl+WFu1LNuqepQFr5MWVIPvwF5Bz
j7x/3i1U1LjAs97IJg3482wLS2+daZEOzSLOmN9KtK+Eb1VXLJXGVKYV611OOt+3tJjoFQsph9Q1
jxyF+0/iGruRfr1bteXeGa4NS8F1yNAiyxRpRt8ZMzxXZF4FOjAERT5s5+EHhZ/+8zhTWLujrrlO
feYjMwjhF1toS+lQeqc7RKzGNs7Drkf7jN37kZVsuFcQvsdAuRFeJpnEdyoF6U4b8ibk6eVWcp/Y
GI8gmFelb4VCLpkXTc4Ef/YYpqJY5zYqAeMLzBIH7DUer3+kIUFjU6Gb/XfxWFS8BEOQMRb4F8ct
XbMpwqxOGzc0d8zbABmZZN3rnGHhvletm44eeZRf5EEc2+dN4dtawlOuBEZ78DyCgFMcrU1/7XGS
4JPs15clJjFFvoWro+5FLgAqSq9w89KNir+ZVzY8v5xJ51q8FfdYM6oBKp058t1iDA6EVaYphwjr
8hzJznmqwq5btg9BAD1Q85Z7naFM+4FLZLuf3apgIHbi7pbQ7WsbtuNmXdOirjnaz6LXsdnoNuW5
f4xL49QiLflnUU1RJ3RKC0bAYVIUKRmKDGA1z56JTPvcb1y2XslG0XAKn4pIoB+W6+LrrbJa/asZ
Wh41Ufml8say2VutKnTITITif6nb80r+OkWZxirUQGHcfzyLj/AXiHqayDMlUKEG2m7Ob2362swo
ZTpzQmZy8b8L3VRqXY99M8zvVckmrK10hdsDVibCpXHvLQvbQ7XNSI6GOhBpjeuNZG3Uj0pPlhZU
F016vf9p14V+f7qxZwaBs6xOBfUVUrTkDSCgPAG8i3ol1X87OBFhNokXJQWD4xmvcy3dM4JXTcuD
DOTu3y/QPp+sLX5+aUj2aKiYilBryNWSEeJZdJRNyZ0etHMu5wK6M85NLc9hE05vBpCceL1XBi3p
TaO8T4bY4JEVIyHA7ZWiOBH94xrY26O9pBE7VgkR03/oQ/uX542t7cNAX3j1uExt0XXD+tVH+AcJ
yeErjfvjS6AfC6rm7UDZIqGxBD56Q2MR/sIVJRzOKrKFlVa/gWSCroN0doHRnsF7ukUFNrBuq9JM
3n6sxvciuR4tLWTzUBWdvIZixyRMC5/ehKp3vS8eZG1/PKIyE5f4aW/ip3srCdtV2LjUdmTYvZz3
Q4qX5TK2m3GTqtSlDL8YxXC1ZDyksxbcpkA3blTaIteZ7LJCX5n+WEFNNkY71Dhx3raepv1KOIEd
j81g2mp+I2kAOkvKZXt4zer4zwMEAR69Xa2tBA7/CMLtc/2AdTQb/XAxpZWjUO2YYOQANnsm2kDB
ixkaln8p8Mo/HK6dp9Ivn3ZH1298J2w+7kT9VWFTOs/VxzMv9sFadbw8WurR95C3OB4Cq0SnyRGB
bp8MWQtcZ66VofCp83fyp5TIiYUlKDG1hvymmNJKEKNJU2zhkmBcVFkYbv6B9uwbJs1mkVwFMvry
zAidBehHlJCDlDTGVfpo829ziKvLyCNaJu7C4Qox9V/tOo+XMDUjPrqfpJD7jzy5YabFl/dBZIyn
b0w5c29hOn7Oq2tsfAoSzVMNXolBFTLC8RKT5Mv7urgSIOOelaIqK2D9ody4eoLdN9jdI0hmx/KN
m8xcFnwohZ2PBysTYWIldbM2s8YJgP9ItjZ1bcj8CZPPJVBkJxlTwMYKPz8AdeJbyC3tSCuNCkC6
VqG3KkDbPp2gDZp/qZzMvJSshebgKGgFz4zTSjCC2LG7wBL2JwkzUxM7Av6VRP5NZ+pkri/MaR2d
X97ddsbu9wTC+bNpBlRhEQ40O8K+ar2fYF3jAAjIAITMQpakUKgfgRJSY4y5yRt+mp52ogXpSJal
M+i+devGLNzQFaOGyl6YN0sdeKL5n3/X33HCQDXcSlTFgnruGK8hQmIxY/wuy6NAPrpzU8NGVhlO
fGF1Q7JknEKps8MPPbzP6L/Hdqi1JKfS7eXZkM31cEvn+BreCw9K6Oa1eLt1tkwe1NFJFpgbticm
wWem5aif5WCE9LBGAvL1RNUtd6G3ywIDK94jO7cqqrwglUDwdyqMZpGhpVJB80LyWZQ7vqZikzir
U3aFDh6tooJnXcUqA4BJ0iiwWXKBYFnJIQRVWseawaI72Ubvx9dDs1DiYTHdOmqFWWwMCQsIUDWn
jnE4B3QCRd6WAaxkSueVYsXvBk/JdA59NPCRhH3Nj7/8kC+a7/tRAMIRYFmtBEItQsE5qx+a6YoT
aDvcZDw4WZPw6sa1RCxBuhuMfG52tUTFHe8HZaIS1+PsZoVLD3nBNM98vMGg3mLL6LetknHzU9vg
BrCALvfDoHlXDwF3gyuA6T0HNUL8OninODAqHEEJAhBjlgGl9OYaLp/3U16cr3LZwn3oAuHm2lqi
mIzqSlUz3AaOeKyOAi2wm1rqTENoPdlRsM4XbOsiBmBzQmJ9ulV6ui0PyEVoSxrSL6+T/Rmh1ZIp
xHvoS3aQxEtGKjflNyvIn2AZ0igntgVfpI8yVxEdOslBEGSAco5lq6miO8dqZrfAVL+3uhmrYTg/
qb5HduEmd9wG5ySVf5mzXHREWHxbUAaVkdQ7t5Ka21kr5sjGEiIRKuOFIVLjsSTZ2x8HQHcon/pk
D9tY1mk3PXB8NxdcQ1xCH49s8sQpYh7jNLUYywYHsf2PjlBXrck2bs3GfcWvyIpvPc+3NXEF/SQK
a8PRorYpbMxT4pvdVZAGRzJ8PTDh5meAFgtirIuwDkxzPKIBNPRBwDjjMKXc/GnyFtQN4kjBboxT
6BUHWseHOx8mPDIeMCYHKhOTePIwkjqt2v0Nshr+0BEYwfEihA8jthMDGlGEViiD+XsOyUjxsEWK
9MMixifDg9IyJxS7lU3fHSg9MQ/Xt5ZX54t5AVWJ/8kW3KKZ8b+Zh8ZE7g/PN4xtAumNKUOdm3Id
L9XPUXEJZRnJmqJhbpf3YL9vku0xtV7r05ZRDJbvz1fyvH1gZr4jVMX8uclIoVPHnBKmOH8ofH7I
C3UH/7rdeCa5FQVx2RZF2ChTnz6sQdTaTrrs+nLXZLTOx2m4lk9CSPty0a/bhkhHUB2WmwI2vCgY
2uJHWc0v34AtT61103aRcMane0aP+N5XAB/cLxklwWzj9Tb8Bh8e7RayB70zeKS8xZhxjoTB1lLz
oOCdvAcsp4SRY1p+0HUvFmVcQIhSBCDf241cXNYu+5RL2r3H21cAMXSLg8hMr6+6BO8BpR73uCg5
hrdNjg7T21R5PI/dVdAu+by0J2rGdU11I57Lw2pPsiRAME3hx6UbfCX9Qf19CZDz9o+S1rjSY2V9
bEeX7/SS0laPavLHYgYOvgB2KmHTwUoLogyrX191WaqumRBFifBlqBynvRzCZSrqHinzaDVTxkAm
CovCxvgylTL5dBSfpgSxTKIB2SNprlnr0FOecWCce++5YzXCmuYkISjAB+mu7QERg/MjhwD7zwtl
aLHu+1kOk3IByQG5HiAYPnxDg9tKcxW6824wyzwRSpyBxa0vw8Bc/iHZdGnHyyFXcQi0TIvy2nj4
jF9i98M1/PEJDkquBew2+r/5Q/BWY1IB/JpDV7FIRYoiC5fVilQvX7qY7rWKPgcOAzDgBGH/Me+v
zYNVa6HUIgrPOoDs7rnp5tuf4vwrMzsijcokg40a7FRmIbsDj5f0mLf0nSQU/1K5umc0389CTgPg
wLkXu8e4vhMEJ1WxbBPT9Kcl+fA5r+dKPuX+6nSmhM9y0uVltqcOVg0LS0ypJizR5URP7T/Oj7O1
zrnwxbMSzjAZG8oates4LWt7PkdC8pg5wu43Yria/hziGDYbdCL3dwhJ30FNSYbWAb4UlicK3jzH
w1gLBdCAnM3qyuFSeZT0ySRRFyRyOTUPi1a0Y+pS/ZzocPN1Yiywjsrdgf5BMYByWaTKJKOwQbpw
0fbaSxbCn04ggqvfxGWxBb441YLGLkP8Uh1IkxAR2iQ0MKqbpXE5vYCYm7RaIMQs1XQe5mWHCb1n
7Hmyk9SHPejy130lpRRyYuzh/SCr7yTFxWYt8i/nQTLlkyEW9LLlXvMUCzQFXZl3iuSch0/Fg75a
rcIYpbJsi7hE2IzZd3XJUTSwiFJNFDYNdgi29EtyRQywbhrOs6LCvpLTp0tn/B2Ww+g5jLOh+v1h
UOpvD2OfGQI9l/hL2VFo2WKPIL095bwE+c09eHgOy+Sg7pDh73YHHVYxcj4gHQWy32fL2a4VSaWy
jbuTHSzSusE3L+zibIHuo33WA4LiLSjFDfl7lFppwA4kENR/6TtPEjAttF9h4rGII/fCFb/htjJD
pFbgDWcCaVwfcEQz/4Y6OTCKfMv0Bi0OGbZmO4YpDGmrL+sxmWmOdVQ34Vpz0Q/hfsgZVzwihT8p
ddzA6Wo+2RB79VieYvrvZlv/bPfaX97dKXJudy1ODO+4bTAzEQRWFEgrOQ4IoIALbG1c6GnTmzYi
CmgTK8K82KLeFezUtjt0Dm6J3/prbkktOT0QYI2lapM69RPvh6eUddctZ98ATIEWnycVim9BR54Q
M184n5yZ9gtE6+xH+gsLb7DPH5FFPnOdhbUM6D7RG02wDQfO5ZZ3P232hs8sMNOJLPz/zO/Nokhs
RE5oDBVz3HRSixHc5w5Ajpc+KCZn1FD2RjXBxdZMsa740AW6bqBZ/M9qP+LGQNiUzVKCSVzu4/EH
rM9hbSShk89/1AvY+ht/ecGcpOobWA5idAkTGkzVtNJjrciLEOfO++qEpguP31lwsDCgo5YZ3QUv
8GrPolu7nifSzXnPEAP9clpGwKROW+OUjsjoAzohlq+TuBzzAvr8bWnolCXTmPy3rOlmDWYV9UUV
+fycyxQkF+dD4kcqAgOlTnBUS+PkpU+jIDJSfpu35EFlmMMLL0m05LiHzUyncv4HdYV2sDbEsQed
jFA7TVq9DlaLsxeGArmHZf1s4lPjewCtPh5s4KVYiX3y8Ks8wuVbYyaslf4AfgFdPd9dHor7c+vZ
5VyAsUTxhnLK+f2Z0iTuIKi7hCfgK/85SMB4qfM/keZGI9waMCiZ8T8QLaj8xwiQ+j4VI0qfM/W5
itGQjinHdSJXJ1JogXTflznj5IHVtfYOPWExV1C8VjS8aDCHodEQ4G0dbn3rATPQMf5yxn8LK5L/
KozeKjGPdQxjtkKXslNDYVoStobZVRfsNd6AirvYKl2GdUaB2oBv1W21RcZk1xXsRSjoqlndKFVw
1u3soxB7n1JwkJTcK22e9dmASBYS1yXZMZFU6ucWBKaDYPlBDdDIGWK2e1aA0E34BTD1bmgojyxi
lS4g0gzTolKD50gKIouhprGfxBHrUmMBU0X+dZ+w6faQV+3NleY/L0ATYlLGqeEMv5wDyiSoa+Uv
ne2UrAkqlB0HJ5M2bQRQ5zUaIo/yd3v9famH/OzCBpljdP2rzx3PlyAtuI3brGIQ5aVYYCbjjBcx
fyi9ok3yNZNh2UfIG7xWZsxenoNUog2KOKg0Vcyz2Fc3m0woWa4gg66Jnbxd7AqCQsBF4Bkej2pj
3sHniRbdyLhFEV5U0GslY1RPieF4raN+jQ7rCDvLiA39wwB1Q6kOic2yTqBsAet43rAVB7Jpkl4v
lnc+uz/3u+3nxplGIy3JRo1p4Bo9fh7WbRbYI2xBCMXwFqVODRCmWWgRcj+2IC3IcxIcHrvaXn4X
Z89PL9pG4b3r+eprdGuYj909OJytXN5zPJWk7d4tzCnt7fI3nwy4D5edCbUuvOdk+SpHr+0AfQPX
8w9vMOqkxrX7cLKoh7Tbv3VIwtwBZ7J41itTWnXpZoQPv032fUdqcvvy47A4vswOwshK7mA1yq24
uuFRkCvePVC3yhwysr5DlDPC0TPtQJf6LzdpHEFDHO9FJidhsgnl7nApoTcs7RpnnpPPwHI5DAum
eWv7JG4rTvb8nk8bZnlkXhv6bM46qWT6CZp22lt2fE/GuuiOAUChlgOQ8uCOpZIWqDDzXRNap8g8
yBW0iZC68gZDj24f73O96J8ky4bFAWL7vLcWZ/WBuJQB67oo+EhHGQbm7liz7c+CH8L4vjYHIiCF
EzzwBoEwHxpCCdsLDcV7lusYxXUd6aOPsmbLHiyIx7hQ7UEYEPUYrZ34UefumfA93e9i1qI/zs5p
RQQp2etB9u97iy6o3C+TZ+cTDTKEzgKok6N4u9jgTx4hn4ptI0tJVSUYWhidcENI4OKAgcS2+xbx
s6yyLjMCdTmCsF4fnWmD6jncRQIlUIMgFcgPZx0ByxxcwgncI1rd6rXCohDRqgMLIO6OLY3EQTei
4y7BV+I23fB7WSgy8aRqIUdfz5o8xLlaGFGKSAc1Qiy+bdXJ0rMYQ6/LOQF1vOLToJUrGa1Z86Vi
OJReH/vIQGYm53pXDrEdtIiCBo+cYQm7KIyHT9tLsscR2i5/fVdhYVyFQBvwI3JWmPyEg/FfI5LS
SlfTgdhb0NOHRx2C5nxMxeDtVdnKi2oIo7lYrf7xFOFmWT12xdSDFSm2MxAqzY9MmgawZ2GfH8+d
52Lr8xY9Gkpd6Ev/X+cT4kX8m899AF1ZPOnhCq6VeZRx79PRkkFl39yOwUy2o5Hhk7i37yx6Z98R
CuwvL8/BlUPn/yvQk2afVt+0NCj603T5u0rdYvnLq6I5baKK1fV7DTx8d0cTwQDbYAeCriMyC4BI
AIkZ2J13Nppk5dBNLqewtqxW090+8LgdBqAHtV6lQfpSwhJjg156fKMl2tF7gUjaUMYDEKjYB6bV
OLQl3yrWNLRLhy+2PZ3yXPABJEduxbQ8cmEecGctU1/0n/c68MPgRjt/BfKqkyqSch3bM4jt0xB/
ACtnTQJhEwwdnRslnsATe6OOX5RQ7P2fJ+yCyBP6d4MKBQB2x7zd2HhA31k7n77PNl2LUb8ms7vL
onlnsjxqEgf2jki73w7bVgqEz7h2Gp9UYDqrpOXSjzHwFQcpKGgQiuKUfZFFF/GfNmLvmFIyhboT
DFh2WdpN0fYD602+u8m95MVLS2Q8w2ni6bMO3IXfqYtvYcAnHhp7l9T8bS5NW//mqQXWfRsQ5eoS
ZUzbjN1fhPgji+8gRpTxUYiZNUY72QjVSs0FIMQql/IVSx/QNihnfasVP7F5CMtuxo8t6rzxK3Gx
o5qw6tzJDHbkN0UV/Cu+1gCW5bnbXRDYeHSFm/5wFMie9j2ZjWU+4xlMmDJnvrikgzBn1Lu/K8/B
NWFKVD1lrkVRJ5jEKNjo2KGHkwsPLF/XSsX15Eq8JB3XP35DXXeCHsipUWG11EVYgG5guwRWRh6r
ChWN+DNfajvv2PVBjK6Ht1qB2f79LTmT6a+5UUZXn60MOPrjJvGggx45DP4NRXJ+VRpV5QtQ681b
6n1/dMK5MXgT16vZBLJkiwEcuv0hMh8hUMudeUmYycEKMCyRniDD18/46f2ATUrurKUfcarw2+Qv
4C8GcqmIK1qfZF9bm3K38LCUCk4eKb/De//l+8FvwyDLIyCnrWLEUWTK5eoLQ6vwDfmvlr7h/j2+
FkhVKop4+q5VxhJFGyJru9xfRRdlm5uzBTS6fn5cmlUgI489zcXKxAPv4+zi+xD6Q+Z7O1yXFteC
hzIY/ob/hKt5r1WQBd6x+AW0vf8uuvExJz2H4B/TJgAfZpaDvM9ngPpfEwXApvJLRz5bHRvp2akS
gy0jgdbZgyRajxJaWFaCMEEjzQ67/HRCDmtrFfuiCbVOfjm6F5MZlS4GVtse+HOixv3z+Jm4a8l4
Llfow0n8V/QnAz+4MyV/kcdfg5NZWpWGvhzfk28YkM6dpJ2NNKbJkNbGRrS/gPlA4TzuCFT+6+/E
KqfzALW6s3l7gkJlhhEbiGmkjjsy6aPq1jjwewR6Fi+wLP+rPRm7zB+GQh217L2IxjeeyCsOIKi6
pu0HImPC/vjJ1q7tt6KSZcaNsviZoiXkQhgsHrFtZaYrxrBmO4hrfLFxM7pumeX0gMJhFN4nsMqr
TzsKgOIYm1TRWEzO8P1LdKbTmmxN9USmX+1mfAD2VvrI5s1PciRgBx++7s5wFeMrRXJdO+W9QgMs
5nPfgpv3ZeSB1vkmCS1oVppBjpv2hlBAmN6m8dftqxFSRFNzVi/dxaBHvXfvLdzsn3YyqPiz3/c3
+oEGWz0XsYTVAObKCFqy1aCcLwKm0FHwgifcvmBqEYiNG2bILwq+KQ4G9G9qhv3D/7fkOkMfol9n
Hy3MFQOsay4OxBf/EOWLRVcmbKKctpHBFl0KFqO4J62Zve2OH34radVstPIs5czjl2PShWxUT2wU
VpM2XFZTWtjuYeFuFy5fg4G8MRVexEneDHkXc5tbw/4kHrgAidwr317lyqi4HCG4hg5dQxA4KlR6
ThKB343BKdB4Q2dOGKHwEnf9Y6eU9StyLw5xDNoAk19cgXR5aP6L8kmrhVRkVnoi8kIz66Tdvs6A
qx/E6Q+G8zOEdFVVj1RWki1bCXQGu9yp61S49HN/ttUa5I4XQ8vm71KQt9tHpHdE0yiENIAJ0c3j
gvNRKJqpIwhXprcYJP4/i9AYXj4QlK6rH+s0oGdXnI+BlkZjIcJOjMsDcAJCKkbv14zCfNPibXxK
fkwe9E02p6B/L6/GPeeAfXQ3mqA9kqcNneZm1kPSXfhr0bWBxiLQn94X2B3lUD1cGcE01SbCsmOk
rjQEno4OzsmC73+lBYkImuFvTA7Ph98gX22RwzzohLzF1wHMnPyePLEacwltGdnJmz96ssLrVkJo
Laa4bc3HYlWNIpq/ogL268Vb8gpLq92wcShpokiwN5lpM7gQzqWfcl/pg9XwYdjAFYprn3i3t2aV
ggdnOrAIZneSO3wxiA//NkhfBHZIiaI7D9vGf/uCy1Alt/JrGwLKZ2ri+kJ2D1vFGj9iAurqSKv/
lfb7a2M4FFu7mN27MlcYPb9QF0MzC/d+MxeGOJGuSz3dOn+cwHFMUJzlT5CkNEBGXf5TFigxyDk9
K4D0lNCDGViwCAezUVXJf106HTfiyCkYM8zY+1zAwo+SIv6xOBYEcozgt8KrsOZXdb7nmXwkYiL6
THywEN1nBLPBe70GWDnMtoIVDV6Cx13wEJUt6JWaZGGV3wJrqu6oML+4SA0tgkJtx6kjjV/hwDPx
+MhAeK3PQSEN53iFy/NGrHeger8LhjZJDaGVyyFsTkA/aDckjIOFB3oQ5rZI1FrrvhQOaDRjitBi
oONLn7n/47tsLDCy7mHEZ4bX3DRYVZfzTCYDBSsC/jQ8GhiJETJiC+7wzDl1m/EQQsSd7FGz9ySJ
gRTQFypDJBdeQRwr0Dq7uXK8AV5hQvdnhyDnETNb3T3XOiQd3SWsCPzoHq+7Frdc/3tVRaYks+n+
djgFZZp3/G0G/j9tXZwQOt7iJq/EhNVmO6wVIwQvqJpKmBfRTiDN+i6yaAGX4uOW4d1wHcSdDjOF
xGfRnvI0ZhzvzwdprCIug2oa0LQKMYFgWNmS4TQ3TtzvonfRTRg/nzmr6sJ8ZclMwgZDDvDW7NqB
1f4Z/SLTNuVRIVEpiFggeMEbOU4lwfVtbGFfHExrPcl16h6ylA4ss7WFoHHKHCxb8Up+QVYa4iXd
WVgdbuh8nuUrfAWEza/EADAA/u60TLJpxEtdXkTfeX2L0BCklzkXe0vCu7GgnSzs0WC2VablHkwc
SX44rGiLzINZ7kv6Ahf4S3AbeWfNjBJtKZLCwu/FP6r2SznYsI9JfYN1zLgRriOgKWvKbFmV6XvA
hzbrN+hhMjn5RU5HxgiAFTF6oMIhyEMs4epvoB1P3gVxNSp9aRYHNvPKY9TLck9fW45kzHJJofwY
HaFBltuCE/R6RZu6bhQXxkJCMsqLNorHwiqGYTu9L2+qE/ZMzgr9NATpa4G81+3Dta1VVqdz5Tgk
MnLarLiJHOp3magrXTwHApCMlx0+y4eRr4pDQGa8RrLyc3dEwn7BMYN2T5NAGkuyfZNMe/hc23xS
2x8uOcV4Lh8GMbYlw4GmBYStWVZGN+DlvHKfghAJi2S+5QUX7+gGrVY9kP5OmqiiAjnjYVO/efBy
6uPDT/gfd2n4mkcxlyLRpgzGbe2SnZ6kNcFoRn/BFqQ+TaXlnMis6fELldrARcLRgStcIXMfLyso
A6cPofEdmyda4pABcwQz166fiHHdCSN7m0S3xGUU4517vfiuT34BRFGpRihacGUe3552Kmbyfd7X
Q1a6wVqRbwdAsT8M8/U7g1nIOixjr5a7DEpRfAjTeZ2ETsgtbpzulxIEMDheoiyyk2oDnJdFZvpV
0XCTw0V8UfzKLYsWSbxOP3FdRj9m6DS3g0we0a5mrnC1Q+ZWo1SRgjkDZzVsLbXvTRVmAEO9Bqv5
iNir7bRvdFBLQ9aspqvtzYRrY0UGg08TW3zn4pLXRbFPJTiOpMvXuYJIwp5/ye9cM1b9b5sNsNaj
koRIsIdYRAr146ZrZxSYslvW7amG1Ce4yyydj2Yz+7UQ4uu57bUERFJ9iOFNDjsgf63vA4WXGlGP
v9oN9sKcoYjt3q266uuoxrDC2lptZHyToMZ2Q3pzMAUrP2YhyURG7FWuxXV4v6wjjb+s5WQ12ISt
hVZN4FB25QbrhmaydpRIYARVeoP3TIT6CHmPaOgNW5g5ZdYi2tOKA/BFXsAuSUJZ9271QWm/E5lz
Asy+Ne0Jt6Pp73T/k4f9g0Loblrdv10/qQsJ7xWpv0z7zPkoeFPOSM7J+48+lC4+D0hY2VJpA02H
OMjDayXgtm9kApWlDULpDAosYtq19xETrJAcLZBx87dpRM59HUBW+MqWBWwzi1XngqN9mMlMJy0F
ORezijBuoKucoVI+cpS88BR+gt3m5gnzRu6KY1xZ2JnMxIbw28yGGgpDZ+MCKQmJhut/3y1/EIBh
UPf/IA5hnj6ICDdepPfZlS4CnDEizD6a1KO6KaXd3C1Eg75fCieS/JFJNLMV2SPdSgzJ3mC8hTnn
5QrjSCbdDRF8MJ1G/BUe7dxNoVpRinmK39rc06BB7znnh4rgbJu45/K1nl3OafkJzryVjh/TMN7/
uOYrZI2T+fdfWWyqfuoQjiQmsycdZiXwk8LEgURJDSOpJWiyJEzaFlni6Y8wki1KJJcFWS9ysmOG
ibaQBQD7Cn0Btqf1HxfTGIDDgvUtrFE6G0UbPhsd8MhrYC1r5vZnDCwkWwIhQum/QnYBP7YMY40K
8wxA6RlVmz/o9USWGTQO8dAUMtIbKzfgWVl80n+ec90qx3KlTQTahzb+kslEvK/hwPF/MnAFhEPb
5B0Tc/0a+8PRBXNTt5MGWh+yTLQ3hwa2/kPeAL4kbGgI0O4FYHs4FnD7QfXx+GU8gLZMeNRtfM1K
BjAdqBJ1XxrIc3Y5uOBmj3EC+2mfeKfYnORdzC8iy++2L4cfQrUjcEVIsI8XLLdISG4bZ7vNm0Go
OmVw18EN36iLGb/Zp0G2FdCFUQrY4NXm+Nk0C/lSR6htajXyC4sejKjXjAVQhST4Cb5iDW+LcU9b
cz3j4G7/93gypOzClDtoOi0RrFKQ5f/iiTE+VfZWgP+Um1Jq+dG7IExkZUy8dQEJL5lwG813OJc6
mtg4Zog+IdHTzpCLbPYDVLH2H4EfX5pJAmXgviaRLqnKpGlHXFN25cSyelH19R3A60qD8/GZYJjp
dV8bMsHbDef5stiKP7woiTG0avAWorEm8DF6Y61haqbBmvM3yz03TDeArXg9OGKckQhyA864a9sc
ltJm6RbHb2DQKME7AFLt0IjLBe5hxTP6lqv+ESsyiNSDxqTO2++uLP3/kq6nkDfONQJTD7SYlN1s
HKDqxbHxjrGwBA8DfMBOlYnmtyeKMKrhZoBBbcPnB0p/tDRSTrOslG9DnrJD0I4278vUdfj+oXKo
GIXeAjLWhFCPp5ZpYgN63Izp6D2p8QaJy/9rg/TfuWiJJQFEqWdJrO+5AnnaBv2vxdUDKqa+7JQw
YHtSxXm869spZOhAfgYWP8ywyk9whbHHGpxL9Izash0+1pGJIafmAlC5Q6CBSkXWZdElwXWrAjIb
hABmx+dGrXG6KA+xcc5Uzv4aQlgHW5pbmd5biPKuxEt/bY/gKIWzQDd6FYk7ug3w5OE/A/DUJ/VG
lRy70/XEw3OKle5fudkvfujkx8hJGKrh+yAddw0fXTtnsnevJeQobzBvdDl0do2a0baLM0JZnyTW
r66sng1tazO7weJiJhRuKgc4YZKcNjHqSFv+vdtCSW465YIYwb/eFEzSTK41aUePUR1QysRcqOc0
mvlaIBRUS3MxTH1XTvXAMqvWuGnCesVu90BmncJgw3nPvKzI4K2B2EyvSms5H3THzzlqx3W4jnCG
OZc1NTpwOXFAcqKBe8WTs5HVoLi2iEa2oQPMz7X6z+3Z1OwNt5rw+IshT1rAvHWb91pGTgdb4FS8
PZCgU7Nbysqialq2YOmVDjugoRcG8y+FjABkkzMMa7bRuybC27jeniOKuDVx0V1eMUkk5DmkEUcu
DwfsxN9RN0Ql7ngO4c6l/610GOXEprhh5qnfg59mMKDstPOf3tOaBl89SeeI9xtczv8e76gmRGMu
JWSIbDo3OJChxB7XePw15ztn2Z0NcYiMBklmyhD3YwIh41ym/WKplIx7Od776UX7GSUOqsLX7SG+
nuiwlRCV2lk7jmrnq5cyQjNiFBfDuFqzrFlkbXjQ9z41+oETvmw1mKw/FuVzEBcX/OPsetK+hYB/
j8ZH57PC+RN6EGnNmhoV/Sm7gJHwKc8z5vun1VLFNPMViHQ6h0iviUB6RuocawZXsZSkof8ig8ku
FUz3Bon9cdiP3Yw/5XjdqmBlu5VoygZXKOAudWXQBAdl+wX+W3EaCRb9Kt7rbWmmbyncaXhzT+EH
XZNqvHC95OYooE3VRdu8RSMa/HEtiTyLLGCijwEtSRSy9L1yc/fAibk28AregSPtGXhXBl1Vqqwf
AhEZRxTzr4tEA6EQ55Pw/0mZytEK1aXH0xZW+oefotpyxV8DTZlcDNJurOejSDT+Aybz6nroXYPW
pkxBbzT+U5XLTpKBkk2v+A1kob+lyaX0QlqA/X2GyZirzpCRpK9Ah5Duy+JZzq4/8fFDFW+8kNbQ
gacgqOvs0xD/ZiuG2fYTaYnJG5e/hOpC/jM9sATIopNo/9HCbPd1wIrpKH5PfyUDhvPBlgqcPvQ1
XPfWwXaDuVF800oyoEjJDSqQHpN73jCT6+MARMhQWrC5sNghdsth4QVljYOdDC+QUZhmc7w3Jlj2
4BWwEhNmLj9VbqcxFPDE5uek/7CLP90WO+cJFUdRY30fDohplYnanBB43tVT/cEI5Y/86hp+iYOs
ywVYTEkzdof5fpPRcJEmiyXk1nCreXYH/JIBWs9+3C88mqOFKVAplQkXJDghN2oykf8h0cW8Rxj5
c3xTCGaRZaaAOrj2OCZxB3fvnKQWQ9aWJEjEAYO6SzQD3uiSQJvka9+zDvYzdlrsbqbuESAKtAex
8Mq5NNMTYWMzJ653sCtrn422XsnfuUyz13lb9jqz6ZaRBDKOYZQfSLjUZO67mw+w+px22vMXy7hA
fBI/njmLsk0yxsGnJ175rt0+mdHXAfxcf7W5+twD9nn9KIioNCdIhtCTz7CGmjpxOYqNvwD1P7aX
U+hTnTtmDxLxaorlkmScxYwKTaB5mNNICeuQKXV/emVXg2eMtuicmrL7Nf25n3TqQJw3rzN+OdVd
uClSCjbHoY6pWI5jcRRAJuR/vxAjT/i5it18tboqclJ9mDCj60DPZ5QaefyvnD49w/3P8elLiBAu
nKphjPQ9r2ChMejLu+kHz9vTN27K/0ysyqMH16nH9G3zhwc38l3ujO2ZfazEkLSu88lbk5iwYDfJ
gc+OyKTBXYE0G03B6mJBKI9gSYPe8TwLgcHysQ165pbIzfaoqesTPa8khQlanRzF5kPiw2wsIif4
uJm1eogdB8tiW+i4ND+ny/OPNyXcsoR+8qVy44NFpjzk3Vveb3R4JbMmOMojzx88rNO8C4tU8aMu
9PxTx+4pIiO2sSMFe4w4OI7AcmCOCdvpMJ0J+Hvy+8hDaf4h5XEWbHb9r6wehZ48ZuXfaGyx/7Mm
kioGOwSlykQ8/ahy4A6Ng8OlAa8X3F9QQZQlrhE12dPCOFjJFXqR3932qLD5acaceQvs8y6nE0g2
n4dioY3SsA4iz0A4CP5sldi5wdmuEmUIR/L3jQllk3jONvTWQ54rrnFfxjUqbYuRI95JEnjOlhe6
Ml2NzRQ/wEVL0085tODvCXuzlof5Ydu1OnQKz9vnFRf7PlHZXU2j6Vlb6x1kJOoP75F9ePOr87UI
CxKvx7S1c+/UP6S6GPdgzE/B2LXWu+FHJNpWCkKP6UmSNk041WPw0CVqLtkSN7I02SXXZeVVdzpH
6pXWYV2RMwVeMiH8gkBDqrarDN5Nj0VeAulu83vfAVANTPV+8DtDaxDkwxfbVmhr+g2ExddbwTzL
zWIT4Ky9jRj+V2l9MuUkcDehdDGOY3HXF861vCO3bETOlQ2uHrfR0vPuVXMo0DwGqa7OyOp5cHKP
npmaUBrKV3OQD2IboWn/KmII2k6zfZjmjUrIgpSZhYDB3cKQb38UlU85oeMtR8g9F8Q1iE2+RajR
LndBHFLij6qb51rucU2qFrWOL3HOrBzU8XruB86iwvoh8tS3oeHI6XFgvBAgRegS0XcrI58bxjKY
uU+waGvuUx97qcwyydMMeMVWzTZ5GjHuHkA47vycwIdJ/ywpBLyYw8O6XiI4q4CrEGLVWx5pfYVl
x/mhh1A4ZmWyPXMlfuCk9bZaofDN4BJ7eeyddb0gfwNbrDvco1kh2rBrN8vAvpRtS0G/oHSmUJ+q
dsdpH4doPtvJDVPYx1hDXxmH/HayxF/Cy3BW7vJPa3u1e+mYin2twzFz52KbIc++6nwC3qYZpOqG
j9eDmHER5OZwo4HW4HA2k6MIxZAhB60LFUMDrjo1/4riaJnEs+BCOZl/RXsp7JmiyKlmqZhALJaw
KKtQQD8I7EPRepW63mT6AHWUkGZEQqvAK6RZKPG/t9zzeU6UwG69HCdNG0jYI9tbb7ppzUfROIEH
47OL+ba7QzoUFGfz/vsvnn3Bl1ME3DejcpWaGFRx7jmQrJOaG0KIfLqDnG24KmQkMJ9rS9QpN47D
yJTKZOJhslg9Hg52sDgCa83UUSkQoyUz0QrhpJy55ygXTK2kxyRp7ybXJJRTE1N0zX1Cu5Wdup/z
wfSPnE7ntyR2cqqQ8WIdNkXQPIWiSFyAxc4apadl1B3WZNttm2zENP/CUuAxfzbLpFflmp7O2wIU
eKc2SjzFlW4msYUfAIQTLQMZdEj3E8c7Hb8kTcd+JqbbiJmtV3djAgD0DIIQyKwUcnkmx0/3bmIw
9sI3N7EzbrF/IaPYzqssyiX6cE5nww8Ftu0GAPs8LAdaw+BJYLTLdNpY+LFmS33PeeWYTLiFyvOe
Id+ojydttH2xpacERzsatiWCjFRNkR7HgvEmJg62eu7AD/2/5J7f3ZtJACuoIDoe1hn1GaRHYQjn
Xt+9Re/ZG6o38zoEs2YOAQJAcr5gqO05/pWCdC6wF7GvYCYzFyX4NvuggJNn+YMXwYF+mAVYOehR
K6GOST4BE9ook6WoH04vU3QzaDU/I17FkOybwOyP2gYr9SsQlxwSZ+EVfINpGvEq5HelV3NU6UMo
mPjPw2Y5B5DSSWF7pqD/+pjmKWZJyEGBfW84pX8TKAedAvt22bJiQRlq4vRAUWUL/pk1sSgYm6OL
Lv3MoR78NQGStlwsPaXK0e8OTAqUGze854+DFfjxSRu96cPEUFj2dNvLyPIJW/IHpcUQNU7gduPV
/wsTZ1Yc2ibqydzTpBxeoJzuRwPgpVTlV+ADo030lYUFedncxsRXdj1kyIrs9u9az1herI7skaY/
KvDDk7G5kVDyH/O7d3zgoV97ajHEeFlAZDShq5T/xKbyCXf47VblRCjrA7i9BFTITzxIhZRZuzmC
92egC9GcSmIxElqN7LJF3jZFbrXY89SbwoW82k+9pD5c/RVPuVhla5qfTjd7n7E+VDkeoli1W1g6
A8c28Ih+HOT2GGqZb8t1+ixpsPfYXNGYSje4Tijpfverb4wloKCjn/GLg+HTjq2WgHU8Z42yOcZ7
gYESVNWlsomBWgTk5rmNheujEJB94SI12fQnNK6PBojDDewq2cE8LSglIbxvGZbabLxox8DbkIxa
iPth34R3Zky2nIv6/p9J7Clt8Wbpk28+FOLRI+0fRssrdytRQSH8WvAqK4NCBqIlLQ26XMXwqQZq
EbJzEqs8/RMLpSyefhuJyHNRuYAbOO2IFCyLKcZKb0cV1a0dprG0E/5FjtLtZaMWBs2M3y3bAcYK
DTEULLHuESRP8ObUWIPgF55yPBZAQEeymd2Y9PNA9S1ajcNUpoHTJIi2SjTQbivTLF9JwaQxpLc8
K8GPt7sL0nF3OVRRry+Uk1/wddydRuQTDaszo4JIJjiyfXce0ub9eJYQkiXemWL6ej+HTOJGmJoC
vnED9v/E9yvpqLNDjRyo6NlSSQqPhydYrQrYJtv6pHpsfBfY0G0ZgSvF2gTTM5StY51xIN6Qyibf
2wxVb/5VXWjFliilHs6njVGP/WE9JzrwRaVwyCilPTcBKc/FvrkZK8ZcsjkcYoHGVS+nQ7oLeANp
DC9CszLRbXyt4DfeFTXvXu42VrQkol2UlZqjOJBpP1WNsyCV+9OZSXk11G2OaxkRb3bTvPSJSrOG
MwJUy30+jN2vVm3EGwBXk4s+kRakmR8ERf5x7+xCwQKrHsbrt5IRI6WQgK6qKQVazPfEczdSSjPJ
LV8RAnl27vNEJCHOY0g2ZelHuxNtmIveinPOV7rNurBzKiBdmQ4sfjUl595hI4ghl9q94oKOcwc5
15Iz3x7IKV6xUTENTWUhkpdHWsDBKJAl1lpfLQr3HJ1kljT9ygHutl0HNPLL324e/BuaNll/IPQn
fUxMTnMYfGQdfevlcOoNuTH+OGRW89GWQVVRjuJeo1rHzIkbVpBvONy0J7QNftwXU316GVAojI6u
9/NQmTxfSL6b6lFm/GU+gZJSMrMq24LIrUwlPjSi/S2Mxt67YkVBBEfbLXVXDViLmAc7+Kn8IlqR
oUUhCgIkO9H+w9us+xhrTSGW0McJhbak1Hpqt3FF9ovqGdDb6YQSE2vSGkf9+JTwoJXu9+/08Yz7
MDWDRVugcQP5Jbkm4yo3kPUS2zSFK4uFqsN6c28zIjEF5JpyqsMjuvc/4T83sk960/+ouUefaz9f
0WvcaGYIgt7ekFdiwCTMY7SQYzbQoQoemmOnUQsNDkiMJUfHMe2T/WqaCHNvVYRQJMSHJYVe8080
j3rSRsuP80eX0EtLh5R2/LnNGKuM1ApY40lhTk88LE9wE5ZsiZ0nrxOz0ullqYAQY2g+KurV+3i/
M012VMu3e6i0HEaXBGKkPY/7SRGFEcdQTHBVJhvxKf5okM4aXyJgjCbfpYUkuQv2Q5J/FJKDVwi3
9tqI3Lx+VLwdNYTJCCRk6gJ1vNvzx9ZqttJ9/WTQh+ZTFqCszIHjd1iB6bpGpaogXEUjMhlRYTp7
qIxVnrlx4DAAl7ZZmmbK8iOWXw57jjGZsLDHYE9lcRjpkJeWGxKNa40ZFeTeHbI4oQvX+CfhM6+h
2TWQl/Q18uYLcA238McmX1zj31z4QaenAJo1AcK45vB5wmrW2xScuG4bt0u99reBBtioMR2Ibs7A
4f4EA249YjscfxHDASZUsF10UheLmek5iFT4eDTGGTYehkhNtvZvisfhAG/sxgVM36FzpFGAvknm
QqHnAB2HxSrtgeSjOGCL19hriY5Gr8y54heu7QpWbP5EuAuSURX/ot8pehm4bewyO5odXlwJrRnq
aYMQW89KVGAThk8OiUX7KVlqW/50hV6Vg3aC+KDwcJGrIxBCTkVDh1zQFPpLiRZNzPg8oTJf6/vI
L1RTdX39GCv5EvLKEflMcO0k1UI1P3QXK+jc3SguHhzla4eO7zSb6O+YxE0oaQ+im9SB403W+FJt
yZGH8ue9KqH4tRUqoBNs0Y4TtLrBEcSISOSsKjAMeUH5viaHK1+ZgCufmnV29PMBpl4vc/1bIXD9
c7fEupAGT4cXxEBgf3LnJkkjzb1mtpZQBf0lFMl8obSvHZNUVZ93B4QcUwdWUR0Ktf0NmOCz7Uuq
YyJPYGGqvoTnmWRlDj/7HpBpEw4w7mzpobQFDOzB5tfrpKx9G42zd0TKIMAbnCiVaB882pJdrEu8
JAUr6QLl12BZ1n3usdMoceDz6Y7FCWzRPstoRH9SHm47iaDYewloc3b1w6mbktUVtGFMyek3/Z/I
hAv2ogy04Esw5azWqvv38dg3alCpa025sl9Rsz4PgVZRW6ahfE2XWUg9+IqyW/2zErCl9rWJrBa4
X5a9/dWJSGBUIld/z+SCv3lR2/++4TyE1lHJNf0SmigWnVMfgfsUZb/QftK5BxQaAsQg0zRI6Kmf
JpDLcfaXBGkiaGJIAhmqGiYYb4relPFyfWVnOkFNH9vk9NnzyzLWv0JnOxlpWp14jqAeUVlz6Wvb
VGEJQifkEJoTd+z5OKH74zLBt+lUVDC4grTbbr4qePJFHmirCzeBqk+aAKERlmWr4KWkEFvdh3cy
lFq/zXBbeoV00lZyWD/N/Kn5bp1Y1TdxLAS8EB2SLYtynvHskRjmtbxSXhqPwgSx0RWl2lR4l+qT
0LBR6wK1o8ZIeyNHO+8JBgk4a3TxXC/MJf9X8JWHlZj/N+nsfeP0LqjLHom1VuiCzho//4EuW1oy
QPC5w84w5JhXZnVLK/73gtxYzx2sxocVuF6ts/Hfc4N4ud9pvb2GtRTSEm+U5W9mQtunF/udH2a0
/wnrm300Kv1lCwkfR/CDv7Zp9PKxZFmRAcgyfNXrC+jXKMD12TqciFBw1l1XOmKSNzK34XahKhCy
aAtXrYigkdk1OM1QlvGz2W332dJn+BHiEWKNFR9TcpQqr6+Crv7RNrfTTiugeb1+QBqCGj54QEXV
4DQFiibS/wAvimtLWOKAE8lkEeJMSuNz+cV0uJf78eKdNiyzrTqqOC7s5aGNVzjDoSOzMjEdvKsa
SshOYL1zABzbjG4cwvfp+iHWuXddHXKfk9nVnoNIn1OQHjskBL31rxpnjzMnKYbI5HM0UvtitpSS
4KBZbzwykiylUDbQGuco2LgvbFH/pAGNwL+Hhbmb06uYxbP6P5kNYh47XQ/zVIcLpb5mPSLCTYqO
X0fBK0C0w1mMY+QSem0GzddaTgQ4vXCLZGlT9Z9FuLfK9+0iWVCYsDL90ySW914n27lQ8/MJvflq
y+yeQSwr4/xx+O98YlZ++epQ1ImOmW4c9Ruuw7CPT6kmiXS84bkiDwtq+hTPcPdR/fjQWUdAP/DY
/EDkaNtPx4+nzPeZ7wieSO+w+KJwAlxX/QwcojKysRXGhAaee3O9xklvsGvK1/HHMDL6ltg/e8lV
rtytHB9MB3a/Rjw5yTBF+oTDPj26+e8TTSVue50Twu+HX/I+orI+RtE3HctbccnhEG0GUwJnssp4
zQK+iwlGDvtvBbQu/us6ry/RyB/rBkzaoiCm+YGq03+Fl/CW1WEMaJFJZnuSdSh8m747m3O+/IWc
iaYczS66MSQYVytTxFcuGUlMFx0f0NyjcFUR1YTkigtvJcLY9ldk6KSKVRBs2rXkWDcLmuZsJAQR
ldvlR+nYOhVSl2HiLNXI047e3yCcT9ciTq3jjv+25TnwkaTGOUhdGIzKQRTiYsj/MC+qtCTECEA7
wopTYEgQfVvjU3HG8bj40CAa8tjr2tmPaFefJgxADMRzJ4PlN7gAT2PjjOVAMV1I58D1xOxhp9SJ
CCiF8K1FOrS2dIBc1dQsaFpbGTfkWwQSrGm0JcsC0jWaSoEXeQ2ktOcfFYqNQHJRtBnZ2WNk23Gy
RuyZgAAQFY6LMV1zxELpxy3dhoMwxS/LoVRdOlac4XbK3VmJ3NBV2zEoSlPURJnTX4xT34oGIGwQ
vONkEamflPerMW5Jd4rWdzrZwrT9fu2n8JD5Ri2SZOJtoSkV1KHavJiUFm+aXu9Uxn46cuNxXtMB
qG/I71QDxWPjFsO+7zt3b7OgVquW37KWayiG8IAzmasxVi3xjRovlR+6iEhy9x5uE8cQPmrRDjgw
ixshpsqcV0tQF2SPz61C87fu0PbUpCWq/6QEnC/d3cH5Vc+URtBE53t3BZrXUxj8nfufwUtw/lp0
mKN2ajGI7EiMK3N+ATNSN1a8+oJa+xI6Hbtouj/lABSKhD02O3DYfQMBeXlmDaF15Vn7h8HXu+wh
qPn/AnPdCh2QZhSOmrdnGNzhrPNY2OViSqo0knRNMumUqey20d4q22GfjoCa2C1zT5X9Nkqp3is2
Rm7t7TuJbjc0a6dULMpp8CN1Udu4lNNfjGPLZr1IF1R1deEaSHpsR8UsNmc+n8jKRsuLmS6SPgqH
/5abIic1TtC8Q/VOYHp2834HAzVJaxAtZt2asglHWpCA2if4mT6NI/NzR43/MPhXyTbN5ymE6qM+
uiMzqdDnWtknYnhIgyEOxkyBj4IdcFhGOKuJONykxphOLiwQAUVN1E8fMGjlH/PwJqt+KE3qHHnH
YgTvm9I644phC0kvVWHR8vMr7eARjvIc4PTqsSucIS37Gbbs/7cVmAcfR9li+7qc1n0CFN9KuqTI
d3SSpV7oX74yI6v1+tpgfT/7AvX5dp84nJEbL8PW0I3eFAL9OqVcBwE2kMj/O4/uEZZuFXURv3db
OC5qxOINK9Eq2kGF2t0rz9Dl0BnKpaNQcAExNQhsIDkBPCFklQAfE8bop9/ZJ1/FCI1Ox6xMG7It
tT9C3BFUXaC6BXtwKhgMyycisAAvAqrZGXQDuGH3tLH6y/ddkP/n+vAM+DUkApKLW8r4ulYgWEd0
j2RTSvJJ/Nw6V9+PfvXrfooWkFm55F+fpy0flEcnv1GPmnMSVAgVT/HcFghpbSpWC8GQMTjQGm4b
5pDbVGKPEsLA8KSfwxJr1DF9rtV0IOuBLSmIw9Mg9Of/ay33LfVGuU5CqkQZOETqL+lZvdA2iqeV
hnh0YtIPkR7MJ+2DlguxwiTNlltC6CXqRjLU71hZkPNPRCobNibtvOY3SGZj3ggtLHy5SAvbaV3V
VAThlKD2hxF0tMy9wv8hupV2YA0UqOh2KmNlwJmOI1JGR7sBgwlwbN8+BXmpBqvty1E1Nz1yEVX0
HkGoaBGlnIC1QUGIG/0zd7iDOpMW6u6tHPVtL0pxZ1j8BjeTnsWAtmBGLtvdtXZ3cPV6maWp3Wbx
QvlrWKrkOKeY2/INqM/7od9bEh2Twzr4Cs/6X9cE76J795h0pYcPfQqMGwWNaiiyookBs6Nw8HkV
TVUz7urUpu7XDZLNU5NTXVCvz//7IwVM9rttWfhdfM3aE1En7N8117zDjZ6TBKOzTXTwmu70rqUn
wZSaO8pJbtBQbY12QSyLz54vgufjmSdlrB+I0oneGx7TYbHal9F8ny3fTUfoyFcjYfmA6AKqXloQ
ivB+gb/DNf0WGjQEh92x13IrimPJkl8TOEMitvg3Qsylxi5O4oUXQrOvlCY6INCA5QevXWfaD5nw
FiEbKvngg+WqVliGgQQNWwhg9DUKWwfkvpTjo8vUg/vR6oMimSVQqBXUpulVkzaROP6nv2f1ZNr0
4QurKrQQUPJmdiiv2RRqBrMlGWHDazXzbGXennJeLVX4/rN7s/I4jR2hYBBsRGkhXPS1vJAWcdFw
OABQHgVK34bFxIO5dy86lYSCzmzYrrHo79DOCk/T28yqSjhr54Hg14z7RZp+Wexao/8np+FIDbcQ
M2iCGR33EiwwgFmif2UsSCoqIVzccRSf2b8dq2/PnikjZfVfoMNIcqvGbfgmLsBZsDsYHTWaJxFf
BHA9sxFkIltca5cUQ/LH1K+g0AeAdJ9TcJE9+cgcn84QJLh7IxVpAQtwyf216yX8kWqBmy+5xXGE
m0ZfZPE8BQCp7xZnmBKPe7tJMs5oy9Sgewlg+KyJaGHjBKMicIoPPXxC91hC8wJigYLpl2UZDTlJ
rXd46tPE1oG4wDEkSwwtWegJds3CliiXFDlpREggwBgq0pHkMhjVQh2oFczd+IC4S7TOwh+uGmhr
UMlGB+zB1fcwaq/CDvf4338GlacRa6C2BEMs9gj5IcMtE2AdbC4kf18qSL7WI2JY7cUStgBXWgRE
GLOnlnGuMO9ZcFTTRQAqI7MTbiFXEF0/DNSCDmIVcT42Ql4Sl9UluiJEvI2g6VMhKbkWPI0MB5os
sn469Ms2TK44GgLF3tQA4kmHt4wpY7SHOGvrkReI1XNAz5Ry7A9RBu2YSm1PSMbhyMY6KFwb51xr
YuupnWLF9FnqNWkyeS2vtBpdFWFQZ2kVaZNT651M+C4nJpFwpv3pu91rr+DLo9Wsnqg1H1Ozo0UI
bv6QvwPB/omcI0N5xriNiMQAw8c95yT/oleZY0NGBAazVuNS62JbemqB2RxYy+UlH7MJti9AtgR0
IKVkxj1+4e/NaAlIhQ8nBcvDbq4Fag3v99eEWcdTH02PKh9pa6Q/fTzkC59cHeww6JinKhS4TpCU
3N1UGW9RVAJYYNEKQngULZ+KBfTkZnFAYVI47NHK2srpq356At0hvkAvne/jYAs5Kp+Yjc7ZRgHF
Xe4x9mkJzUCfX/jfUTb+0OH2DUW/FPPaM6Pja6MluGhZyf6X//ZvtzgeB7jiR199wQpeWcKLXPft
Q2ELw/nNayMmHt+tDqHPUVgIDrAj9aG4DkoQWycQ8vOmWEY9L9HZoSUfn6xwYIrSalj7Dd/HVLfn
neJEMqqRmgBDWjRhVfXYoOPpuM6lVlS4j8BcMCQkNGJDUx/ACJ1vggHgMx/x58FNvqmMHoIw/hou
crUeIfIxkvIAhr3Kj44D4/dL/g8/PBqZdGmbIBJyBCSrae6KuJi4l6ziFc/ymCf9yoXIECEmzq7q
0iJzCMyjLOJ6Mp1xpY74sddakmzHOFkdbaH1qPg1yRUQQ5GwMkg92s1A/1dDLZGgCIxBbXqJiypG
XDI+gN7/7S0uA1+r7ASx06uHHO1ZhKAoNK4B7CXxDj4Ys8L2yiDo3ItOOg0l7y7mYxGSEEJz3KiV
Fxk7FuMKW0Zlv9Cs0G5ibwo4szjClWxek42bP45xWRtBuzL/RTKjOJayDaS7RlGCis2HZ3dIJb2l
KETlol/fCStiLVpbTDwylMPntP5FUkcHrbqjFck1wDEDiYe8lxTLqZ/Lxf6VMmDdlIaeFqlXOVUo
PUn6Ptq1YmD1MoA0O1ycek2FmnVeqkRLsMo0oNHpMSo20yUpcUuY0cgV72BavJ8b1wt26n8AiCLB
IuAmR0EFYXqOtTEgNiWB2W8pyhzU/B30mAgUU4rsSvoYNaYhagv9wViBHzGDHg9zML3Y4myNeImq
rMOOd1YXLkBYE0WoCvcxu7PD7v+rxDE3+RXjmeb+sZfbHj+9DqHu/6CdS9IpRwI735Y3HImPw0lE
UmK7p40xz5eHNdpw+1KoHV0D2puwvUUg65ber6CLPRiJ285JKThfAh5D6ZPBE320J06k8v8lY/iu
yTa5RBTHP7s/yUod4GG7YW/qadrDBGTO8QPwFdfKHdogkHpc2HDH91UfwVv6nbHWi+xjf7ICSJCv
jfjcl7mne+aFGrs1S6QuTPimtIv2GeXPIHwjXVb3XlDA0rsIikoCHF6RF727J83tevIlkXAy+BJk
EGS5WVr+skpzLuzvv0t/0RSnhEY5N3sg+KyV8CBaUwE1FkP0CMTPMxacK+NWlowZtcrXZRzczKK6
PJP0+XZ6pNsLm+2OPbQ6s7htE3tvthb1+GJ7zS9DfFBS94axPSiZ8qe302ND3vT+zLM1/gwf5GF1
u0t1S4rwyMjlmr26qMMp/QdkkRUydX0P349xtHDBlRnFJNHIOBfVT84lu1AcfcsKc9WpliuLcg4e
OrAZe6QI2cY8sHPgK3wcdrzWdtfdNu/k0t1lwUDEwyTp4uRZ8uZBjIxtqLpzw7yGhgYZJKp2BGtp
E6ZDMFOZcyYlz2MF1M3yUrEJfBgQbNS6Xm2W0+b0GA6YwX5Kyw2Qo+PvJaCgMg5ZEjMibWTGFRxU
UeHcERAxduLYZnO8zvOOC0LTI8zvqMtVLDLPon4gWg6mSjrIlrtSW/4xDmKn9gllCSudn0keCh6w
NU8YncNx3+45lXtHl521zWWoHZUIWS91+OIUn5Qaj5gZS6FG1yp9Jv3+z2a/xpIT6zITD4uPIBs5
W6W/s/OfCPHygmmnztNlOFljgedB87Dxj11s+dvAD3EaMrP2TOGJLg7qmHJcK7Dd/rvX3cY7xUQg
/firZ2bmTyyMqPKtXZURCvkCJpepO1ZSCwpA33PdylRXo/LhWf4fq/lO0NXwlFujsmOnm9BoGtG5
ptW3y7X2PFlkt4D6oJPZ3AWuKJT/+urTx0+yXRQy2AsEk8ku61Ax6shPUIK20FqCI8saBIPghAQx
rvRw02onDW01UvOndrz9sv5L+wesXYqvSSoqrPIshA16tZMrrtXEQWlTosYyc5C4BC1sdiyXKB3X
apWRvwoswWtTwISmvjTm2q9Wogmn+UstJ8zpybBkES43GAeUvdWiLWkuFQwGzOsQQM2v7WF5jqRG
4zeQAn1sItkGyZB2ZzojZeXSpMfNhgW0M08ZXG13hzWb3m79ezAsHmd21HWFI/gTmc98gLJMv21v
LuePG1mIxyP4DnXsHJLA1ToGj0nA1hNbI/Cszrln8tKE9ymI8kZhbfPPqY1I4eeq9yEjg2K7Tnsf
jG58htaCVwGMlHe0YxobBCIS9mSU9ybvRmoqRdM6oRFC/ezvYqTehnKSUQNIQLakIZlWWDuw7Zbn
iTBqZdjuNCxZzN59a/Gfl2ORGXYcxiZi4p85p3v4fMCVlHE2x56/m3vzXBbmWTzucRb3hX/tgCd9
AATB0oLgolGA91Abe4nOicH3G45owP/2/UTCD5WBjk3xxTYEdtWOiwu63Mr+cysRNtLN9TuvFerQ
6I/8emTYmitEAJS38vPneNj6dVJt5GGDodSxk64jsgwgFRxZeUgUhic1MZ3KfSjUetg+92bhwhH5
j8m+vOv0OYrFxUig3OTvgBWlxF8K8DiVuRzQiSnAWleen4iAzzkPSGEK1wF1wx5drrNgJobK9cao
PTjuz0X9qYvIQB04CXChjp2LDzYTVCNhoyQXWrqPsegJRNel27SGKOzt2M+OB0GyWWwEFBBhwQPz
JFnxQqWlXHM3CpSYNbRbdacetI10O3JzZECdwSE8neE79jIo21zFbSuqXdLGAaU5SVLAvrL46+23
MTvdkzYukFRlC2T/0MF5cBC6uCH/Ftgf3znZQ/buycxULyt0zSvQJZ7UeUWlH5e5Mjd5GrGSlmHr
Llbi44EuuG/YhA/IrZcbystPlDLAFCfbTYxuA6wfvvxAzI1X/H+HQpNjubog39M9W+vRDI/E9Lhl
cKOmwFk52iGbBDSmik45Wy6jPHIiCd6zWSqV28pKBJ3sM0rt3PcVH8oZ0M3MRK7VG01lQ41A+QZv
a72aYu+EJHIFZpSHpZ0XuWhxVYtOD/ccqprD6Qcl/dxldEfX3KeC78hwLjXML5CL/aVqBiK7t2h2
ieZeZO1eP2Xiu9B3xe+lyLvweqTkELdZdLIHLjW2pN9BSC5fxg7MClBGaFezCLgY2bKVteM98V2G
LWUn85OpPBxONmca2gSk9bI9PWYXFBR4re0VALanTDmzOZEEPNnDeblccdN6ykKDHEfT6P4MNIhH
aLw2SgZ7aZP/Aof297VGVqfK6ZBC25YiySCYeAL4kBy3wePREKhhBYEIqI9s3R3P9p/so524ffsZ
gPrPAgTFl8/jvpQKnrGqdT8bpXUXRHrMICQ4vbBbg8VBFHBOdTj960cB+OgctjnkiyDRdrzXP1mD
rrkImm0aoa/OdBIuU9OvMzwaOAY+KyxmRs42EfCEwmmvTZFB0VFV6MBdf1gnu5h1CJIYve2sMYMD
+bjfPIHgeEKzv7K+CjzRWnGoXWdn+6eaops0Ma62zMK2IawK15KwbOZIM5sYJK7K3g88HlqKUp8F
SbHsA6SKHHT4Kk7cYw3pcWfRpg+g3TIQsIk/jZvn/vlIXO3Uhs8RVgXq+1RH24Jt3t8mIi93it/w
TW3jpHDsuWEljIMQ1ZKv/V7wh3Vijfus8a/MrhbaTYBXkBKCYCyizvF5hNVw92+8HILPN6Luxmei
nOjyB6PdBLgJuU+8lKMkrQ+ZTiFv+ZVP2RvpmHw8wm0BBp86ac0dCKCrhObV5hVyho1eaFkxzSE2
DHrBNaupc4/XP3vRLQvvFiYYgY9oOF/5CQawRRMiyVE3GCkFuS6coeGdO3PZkmMystpee6caQyv2
rVaSH2lmBZT/aUZNUNFvPRI9ZJenb2H0fT04SoCRyVGE52FYuw/GAVAzZEyVDMercSJsLrXJGCn3
jNe+SeVxxlkGU/YU/1k5rr7ClJnIAJ9pNPQV1XQvIgx6Rjt2Crqff3HeZ7IxNaT6m/7vGfO4ErJX
aMpIvYS3FxGa9H9y1LKf0koGL4yFVD9igIIoeX0Laays1SLFwHphzXHCGULrnmDZ1kUFUuSotVAQ
8uifOzZ4yJ0uSHLjzBGeUnWMqi9M/ddDkwNVOarvWCkwIVx4ve729XKOWRnRI0T7IzZe2gQEaWCl
LgcZiBOgIlbnHWRIvIKlO40dFWWV0jXojQ2wE0v2glWw5zrC5r9ckEBOFZrPDDyCejThNh5Xi7lT
3Nx4jy32SzCr8vuaphzHBQUUmgw1Vsm7lGta0W6JoLmoGnMSECdVHxFMBKWE0jCY50wQgrGLbugC
/G6c+2EdUB4FJ/1tSSoST4PRBu3RvDh9l5SQ1a9FEjynFtoLMVNA1LGEn9pQJrnYV+O7mN5pibed
32T1GA8pw6imqiPCtIXRuilKVDkJg9DdtECH3F7p1nBGbvqcUHasFJSEj6Ye/KTjdgEJLIYGW2Ax
/oBlrfq7ZU0AYtvmhvJdvieDBlQZjv+qApbpMj5JjwMO47Y3LjfJUZ41eUy3pTydxulEuvWXBptT
1MPMOaz7gfpSC+TQMDoF6DrfDV+4BSd1vFRAnz9m9OGqFjyPWP4NR+h3Z2Ea+ullV/fQ5yNgFc3r
vfhZaeoj2udrraZRktBChaatUUTwz6LgQkvUUWSCOl2UL3T+PR+4gjCvCRWNWflpIuApCR+9mRQk
60tHnRgTM0Bh127dWedngfY5hwtiqggpF0vWBhou8Hbj9RtEd/+tqrV9hKXBoCY8HRbWR/bDyOiI
3LXY7q9JsnKfxdPed49aDJ14wZchHBYJiuqdTkOiqQBlnTtR/+qTAvoDsPP/jKDp00YGmh8qRPN9
foeoLrM6RMssHwSSqMfAHGVhNkE7e2+B9l7fYSSpHTOO4unbAqB3d3QSWiltT7ePqbKlA2v561NV
2IZsiKS/4pyRbbFvz2Z5FOS6D45AdcQlN2g23AKmWPxVECn9uoaEk/1Kwab74fW4q8OnhHjJdqKF
LrnFc0RyQ1W7YU/qp9kHgw6M7l4HzKFV0b9Lqh2fpBDsUV7q4OsykIb5VPgTVrcX1v+vL8nnv7Lb
pT7NyOuFSl6G4jCvGTdb0KHHFBT6l3PGNiZkjEog2m0Tg3e3BO8zLOKXfcIUf4f1+qnOoyQMWvRt
m3sMzJl57bOj0W8AX27FOfiPv3AJSI43/ZU2ha8dstjJ31qhfiawMbirmrC8DOvZmY6GIvn6FMit
QhV7BhE5BdJDUI50WGT7gfGrFP2o7Ha3O+W/nd1m8axZn4T/VTOVF1138guFluFWyn+8n9FpJI1A
0YOuINHl5VM1DmhfSJnJuc/nYk5ChhC6aKEGy+Ld1upGZhjJO+HUqD4nGrLBuZzV1ofCUWoymejO
lMzhzOuMYh9Kn2oiCOdGgFPiFnGIzQ0Nog+JUyOiong/9MfL8BuzTdUnlaq5bg3bmKUOmXZiKBnd
l2qpz2BnnDDw8+DX61dj93d166a3L7lE3Qw41sm5Jf9Jhf3IiRO0ZhmSIPkjbE+5K2klGuFvGd9/
rmHGXjF06fCGnFkaa4kDLljSz/DXp20IQ96jKhp8vvDryA9qa2cHbMucQHyahuSWx/df0Btglibu
R5AkKsOZhTeN8wZYLbx4uAYW5CnQ44+l2/R/zchnzFy/1ilYmhiThJDuyCd0nMN7jOJ91NCAa2mn
Y9Qn4gJrQsegODo+/o1oc44/ZHmGL8fOXGN+eeZMv5yym5th/KpvBamGkEYJ5lZAD4IHGIUjr1IB
YUgI7IvNQ51hGVzV9LBTI7J894pT8sqB2pO0YG9h4gpaYScJMbkHN9BosEOL1OnuJf2fy257Q2h7
BkND42/zBkU/3Gx+4WK21XF9c6mMMXwSlotORj6RE8XF2EQCa8OEgNzE3oLXyIuv7URhIZ0ZGtiV
Zc6OCmF0WnjhQWscHP4WL4D7jP+iRoI65o0cZxZCPh4kuFsjVMVJFuKmPdYnvLScnZuh7orFyjfg
d4+5Al2gnQfp3Bp/iT+LPKbZR7eyOcmjBdGNYG1XexSBodKuQmFElONnnkzspzq8M+HEFC0QCwTl
AGWbJ1QjFjviQCcY9lfwmuUDAkI62SES+TvWCptDeznKeVFl80gHBoIIGhqwlU6zgUuAHUeqAhcD
kqXPrbmKMbYJ0Pedhj+N7rF5qE63AZsKCG65HML0sNg3OOFt6qnKzfjf60X+CkTZl75SA+ooFUdS
pd8K3xRbVIFi5fbQkB95xbY877WFKrBUpomt6F3NIG+g6UzpjSI8r7CoVkeDjTvvLThgCL+jksyx
89WqX+g8R0VD4Ts6rigJFjQJTILTSo0FLLSXdu036/Ql98LRsvcELbTNjAMBQ18KCaCYCSY6jUWg
S6nNCSRbDtfUHux5jQWcxiTZRgQXD2U3u277Yangblp5TYFbccXF2Ii2VkKoQ6JyvxOYiqq6pQlM
iNgkGGsYWk0T4EpqDcIBh16mlwnjbFCrDlqnT1zJYq8N9q1HAKRFm0mWchoxmZv6hz5PccSVMEsJ
mZ/ZxeXYvoszPdP/Xz/osu7P4dgwdJM32/8yuVP9Vbi3KMDJsD4wYIhJONbbhGZdZCHjtzblj+dw
PMt3QsCb8+5DKoqD7BQmfnlVhivaoPb8zGX6TCvPQW36nQ7Jlt1z7jUr6vJtJ/KgWnH3xS4i0dj5
Fv1ojoyMGOCH7GzMGSYPJ7Gzx6l+l7Fw7hQn1jRj0PsnBEq+QEwzYUfxkR6BrWkiW5l1hvMnSNF+
BUTpdiTfEFwZ2IZwk0wOVdR2oNKOd3cGtxayNBVJHUyG7Y9AUzvdlAD9C6E5MgYPkmx/bH5D+0AZ
IcIP4uYfTbE4V/1MPXIugkLP3jB/hhIP6DMIjnUuNDUkb59PP+QFOGtEFB0BtIeKq2/XnpBscmgw
c+qE0j89Tv9qg/Ppn7oTJlZzNHxMaUtHsDJuHbBtKYh5TSHU4B0K4LBGYJbiAjrIoNuQd8iRxoxh
ocKaOvosVBInAelidxhN45Xu5FWCDrZC2C03fYAZ+xfit9/r9pHOWU3w0VzTpbVGESX5pCmHQa+i
pUeaocsyFNowDJ0hHWb1o9KHOsdmaCYHgwRRyhPgA2yBO+X/RefmK6Y7zlIWZgUGmzC7Xb9HKsN9
3WO500CI8cTCVfx//OR4urVdW8aiKcSZAqw7krIY1jSzZPDjbcLaUT34txn6lvW2pWj4a5mj95zK
gSpmmRV/SfZ3CSqELIXjTMlEv3neBTzN2Dz0g80nB0/aoCVzFaP3vdQCTF3rttE2VPICwe5I69Zw
n7qhvnQmBnnhLsCXqE2E5poCFQ/LPYqVZdUrRWcclreE1AodWjhc0tHnE6c+Fc3cKW1ue/1k/rqo
J7PhEq726G+p8TVcPheayWTj86Z+ryvOVUzXCOVgtI/+xsNUJ8+Rec5DCylZBZkuLVd7JL66znuR
oskynmLq8a5l7mgLPdiFRKoxvJW10uYJq2OU3OGadOdUQ0Idd4DpUa2qzuepUDpxk6AG38gPCt4b
ZXMNIeNBUMuhAsS6ytZ+7Bzc6zJb365qtiSgXQPMsjwkkhTJ8aH8OFyyBtXkASTz0RYiSO2ZbW6w
whxL8RwHzqssYJ/2mqwmFK6pBERm04rC3aIdmvuiRM6rdiXU4zhe10Mw+/nt9DTnAo3ZDWB8+NI4
vUhNRLENLPNC8AQEp2NGtA3zjRCND9aSir9F2F+Iv0nkYtj6V0FpUYsrX/lNKIttIfb4dLFDGaSM
zSHR97Pr0MkqmiwLVF9vag8G1bfgDB4cUGQX/wNOp0MfLnrS5JWYUZhte6gPDnRRRWBLU3NpBEOD
NreLBBwvxN9HKkSuIqDIogQ3C6ac2UuoU8WMkQW//7aVG9Nu0dT9DsPdZnwOIN1oCZAfqmSinl9N
sHMF0/3tjMOgX099dk2Ioh6oQVNBI6rKqaLeJAspFdeBhT6nT7BTTzm6QSWxRQYzTxlYDSfACylQ
DSVQCLN2Et8riWnOItzDY91EkZyRPlpmVsQ2G4kNMV+5gAlANibW6tYa0EjIp3lsgiGitwWGqZug
H+didkNpF1UR/6/Wfawl7VBgScyxd1K3TBJM1K1qSN8TADugtsMJRMhFHY9uo9DjAm3zFCTPkvsi
askZcxD/Q1xmb5Atr5TLoDNJmj0js9FxjO/8rA93D/KR4qG3H1565HPa5XwFYyjOm7t0c1dsuqVB
IY1KYf02hvC6vD49+rwcLStiGp8XGVkvWlbdTaF4ea5lPUQCCfbqQJLm1MgrJLv8DaHO6WqPElq5
1edoEi2f5ZFSq8FbT3DwOzB6HJOOQI6PR1TUoXDWrwxh7A7Psrn1SS5Qd1CLBrETkXFy8oEMTgMU
NTjeb2ysXpdP/pBF20o7c1OjccVxrHWGAERsr6HzUKwyZmZlw0jignfTU4EeY31xrVMLwxK+ICbI
bZ4dMXDSlGJYxfP/ur4fTvTssK3V8SfOOl+bcORqhu3ahNPJCetk21xvFXWL7c7mOuFK3+bhc5at
HyvUZ9uN6O7aqBLGkS106zMsSgBYoJy17mXbb+iCXV27L4I6A2KUoauxmrFfDnxpBddZrl1XUh5V
PybH4D2H5vikaggKABnZolAPYlrlAJtDeY9rti1J/NrmzjNdmcKX/C7z0a1aqwuPZ7gItCSHE8+I
AOG74GxkazgptWvQspH53VsyhLYD/AQK9gQfwUvj8F3jEW4kQkvX98JwWcgvORjug9RhqS1ArGJ2
pi0A53WqgEHtyqxN53CzD150HWvH7mXF/YPz6p5aiCLWn7jhXUN8Z4fn1TmuBjfTXvoT18cDeJAp
zfcsQUconN+geTflJdmQ2TI6Vt8wT+LVd+ADQ/Rv4kNzBtItH+fmHoCL6yVM6ctMCSBnGbLPgFhC
E3wD3syW63/UVNeJCdzhnA3l8bFL8OeHRNu92LgdbPMU2xMpTRgfFzAx+UyhYRcW8tZTjiE2e+CZ
MyJ9QOjRfmCM3g/SRMCEl1+7LWnshlLZzosMIz/xhh25KJiXAey+ErCDMHAcE/bOYuaDMszc9MES
zzvN6qJsekBrlo+csr0W2YCy0dkfZXMl3DOfrSHSyAxMoPgipJ+Gnq4IXkuBzGyNa5e8Ai+bQ7B1
INICx0rRAcEtJnRJAlnGfeY/BQYmggQt8SIEj4HDzN7yqamDSSKaGjOXWwEap7KwuJup2720y7pj
yCYa2qnVwCvgnnywApWXqR9D7LZesYxelj2TZoXeMUWgVRtWeJbDkBuEjQOpiut5avsAYZKE9jfU
yzwnDHcRViEoDyg3C7iRFD4pdQvuPCkfi6c8u3l9j8c9cEsibyKuuDu4dDYwHYjAR93+5iUIK8C4
YLIC5LskMSgj8q26LO1WU8hC38SdF/S9TJpn8STjLT0n6bW7PJkHeJ+dTJDCjSqfCB32WBXueObk
JmYge8Eb0iq1/UCLSAEAdnU5t+lPrXIe8bauDoR9PHnOsgC9HIYI+8vbTSPkXSgwAjDuBM6cIR1R
m+Qgmbl51e84gutU0Q7UryBhRrSu2j/fdBbe2RWFR60+HCClKlBIYrxTVx4a5e91nehnNxVvzrqO
1js7lr2hR//XgZGNDJqG1wsRr/bEGUuBMIK2kDthEiZkTdckxBwwi5McSphZVSo8Rao1q8RKih6Y
apoR1GJlW4sluxWfpbOBWCua8Mh0YMnHAF9lLrnYutuPHLEpxd0ZCrBhKMA+bw9/vUX9DY+V9DYO
UX1rFfh30xsBSA23HiC8KGYXfTFm6j8vYilBkiLxJwwSKK6GWIS5Mf02acmLpBNFY+j+4K//9swx
eC5HTwsTTGQc1Ea8BYpIWrWOqhfRSQrN0bweaZDFA7Jbtyq7kUg4ExgSnP+IIKzi2S9TKy7ol6qe
9A95GBHfwO1hxcT9de9HCFurAbNTbc8B3gYmcOAMhk9NXJVCN/MmwgleQspT/1yD593LiGK9cEAr
qsibPgFri5RH9GkMyv1Pp9i6CVSy2NR9sVS72tGdNhE5L0nRdra1XrmRGKGzLbSXpZYq2MegU1J9
mI5VVxQjTW1GI4N4YOR1X18IZV7DSFD8w7LGG9nl+yhjQJn9Pfv6vZLLDtsrs0M2nspJ0DBVUCxr
Bo4H8ywW/33tlBD2d4+2BBswvw1hrL3NETReLH8NN5WniLi0iU3UjoBFnAh7tyPpbULZG6vOLUZZ
rSw1VGzzZEMeIbsfZv7HvhXNNvthB1cUydPzrTCNabcAUgeXghp5wHKtZf/PK6wdvydZh55i2ULI
qaEtCpUNSa1rf86W8QEndzuqg8pZl0eb2eCDGMhY4P0UouqTjZ36J53K+ObHyVAxzyrnX4S2qcol
3fjOPGEGzm5ZpaIOdphtyhplPz8fhfgS2/bWW20ocjymZ82RWoWtmbUuqn/aRt7EaWNa/H5tT4g3
tHxs2lzUjL+STwT2Zcw/1mxZ7ML9z2IEKBgecrriJWq0QIEus0J1S7P2vMUOf2ueb3CagDiU9Ykz
qgRX4HnM5xl6h5Alm6gaERtgv1Aq4ihqTeIYImkn3SmQWUSlXa69/HdcKbemUbSzVzfcK1fjTNFq
gHi7P1DTY5BT5wtK+q1Qw7ymNVl1p9cGOzy+uGJY/o6wdPbmjJI875cwyRX/1/Anpug/sTT+inkQ
nV+jpZqPt2B2O374OYzlQfcjnlnqsax2G1iMxMfVuuyW1LM44ETsHGd+cnA5mGA3G5C72A4CYaE9
VvkLI6yz6v38TIbpD92Yipwr7S63Kmt6ujy6pGo9qnkIIwZctGrYnlAJVBRU4v8F62RsP4Lx6rLr
3xy6P1EkFoR9VAOAXjAAREm3NUGz6WbvLpsYsd9m8AzhfksmwZ2CdJTUJRaOxYEsd8+82ez46wsy
tEd84QdZ9kV5XqPx31zSM7Zpee0fCOQyEMxU9GtAsY4FOD6E0RV74zPQGVz85SpTC3JPBPmYxneJ
mR4YYnvCFmmWgAm2aAVfm07KH5TvqJcW/vZM9taBjrD5MGCkgyK4cRS8uI7g/tQtqk6kl3hHLUPD
ALZwFoORFiUpd/Y9e0jszhr/IW28QC7KyS+cJ7xIduQBtROPTi7XTg7NbKKOEEpnxHypC8mnDVUZ
JIMAYy8wEzmYu1SkLnU9+NlBGbERz3XQtzA/vCL37Q8YGdx348sU2LTLoqx2EsouJlBk9gCZR1ns
9cp3oxq77TfS+NF7hybKVnb82UU4lalXNwxdXzzXS9+boI9M3GC/GpLIx2UbCgIYc3v9MyiDSFUQ
Kq/c/8p18pUL92x9Vy2GzQzgCous4Lm7FRuA9yYiJt+hm9ZnqIvEb3knvit7YC40JynFk7Ib0NLw
0v2885g5/mS58FbKpillHVr6ynw0kY9HINTlZ45gIGnjhb6kvg08g1GFQ+OnHOO6r5EV2vOYLN4i
quvRMadDnynudcbSK22ijf1PhAcqaKCclQZp/u1tjNmR5xmkpgyXqxRyN1JL53raVbu8GWARnyH9
3vW3e5PWtDflSFj7Wm+QsdAbSnFtXMURwhBu5PYtVng74OLC9E2ylgVoIuDodbZSzklVVa6aREdS
vYt12RKCgofxCjcLdK8HmZmIBhITQDaaBuZ7dFKG5zPqgHxpbRWC8wpFTJrxp3GD40dehVcbgraX
AcQYdnqwj1FoayQk0sBV0sfjAqaG65Og8xDIReadlPNRS3wlHL2ITqSCqz/BYEXKvRiD3MWi1LWq
ZteLW8Z5UO7Bj8Ih9BjEeigcTZr01D5NLsLx5psNbGWvQA0z8g1XzDamTrqMhbwYXTmvOfCEOBfA
DwjtxNXRxj2s3AIahrIan1nWqA/61zpUc2ie8wAEryLRgS4kfspPUMD0Yab1b/U1A9VB2R2On84c
VXJzJITq5HA0V/DaOIlzlOweUEBmlxSGmG6kzfNzUdHncwEnVmo8BeOoIdXlnNIF5dc0JGIYG4WD
7E6TzB1LMCxcxGvwCJCtv+eTsbrZvTbKUFBtT9iWjashxhQba90i/DE1UOpjWtTgywVoKr7hq+2l
oCrcpwaZs7LyixO/Ov9c5T/M4dBkuryWLvr4+61KgqfHcT+hHxLjSxcuf9WLVvfXNWsoaS/EWNWl
L4IfMf8T+ILyLLldpxCbhOfIlzNpnlo8gQdqp2vvz17eDIa9jca/F3+U7jCFW/0lC/thacAyqz+D
8z7xr8xRkDJJna7hEGwQe9TzwbEeZsZTyy/ZTK+/0cfkA1svvjQfyvkNpCp/LT0gP1YF2ZGC3MTa
4qy+Y8ZSNcLJGtHLpQoXgZ+cjM8/acfhsL5BYez+o7FSNJZxXx/IFdpSwcX1cIgit1E51HT+FHyP
HXupOulnIYqHqf8IaXyj5gssNWkjEPbiLr9TLIQzsDZiIJIFU+Rjpio3SXzCtInY4lmv9W0MJvj6
w/2VCn9BPLj5JtQBrKd4JrDtle728ZPdFGHjlw1VrJb4JvyOnKdxbfX60xGnUcZxuGXD0ostr2ts
DMh9I2PSHLwO6IE4lVXhHpp3+enXkDWQRZnM31wUp8olZNX+RnlJexZ4uSJ8iVl+UidRsKbHzYuX
tQCCQyrQJNH1rwIYtXdwq12TKVEqExoweq1gJnPK4mnYT3QydQrw4WwGdMP+LQ7pyJas1b9Gs1fD
eY5gz3tWNNe9M04amAvO0b9miUkZ2LT0ClANUUXr6Sp8m+9NIMa049ttlT+kyMr4xWwlGkVY1eVv
eiODoTnSETDbzaGVijmwKd8P4RflMOl+ThDhUPqUJ0+U+t0yTFNgpGU9DpuuvaZJbMhv3b9uQqvX
T99DZd6kkQZ0xaUENDb9jAb/RVmE5LYwuU0Fkx9a9rF365Pm0kq4rOU+3SomK9xxmZWx1MIh+yIP
x2ZOe09IyH9e0Ee7GeczBc0CjjPly0vFMeqkv3Xi5sQp7fUnFHE+vurKYOpkrZqVvyPaKReq3wCA
9o6Yvn1sgm0+HrAPwgtjozidZAtJAgjJV06rP/xKTRZlJrbGeBWrZl/7mFxfCTLvBMSTjVhjw57V
nL214ygogDWPVxejoSiSk6+5xnXLeloLdFtrAN2DcI3D6EJ8/atvk/PevXtdmvsYLpkA2ZLPl1tE
2S/u8DAJieHyQeE4Q29VYFIbrNivzxd2e5JlABj0QXeNsMiorI/HlMnrR+Cj02XWIKhZbG15+RTi
ybCZvemzcE1Hfqa5/ZFw2GPDwBod4Wk1GSCKvRChyDjsslbn4CjG3UfNnQWav5I3P9kIKhmqUB22
ZSMYCR6xMfnrSdJOwpZL6gJrnGleyzAgEJwiWZlRy4QO3Af71e0wEylhxFsv5BCTItxkfT1GL+EX
QY6137608YAUicyQpwNCkX1+8QId0iesUAe3vhWrjfTlUl6zu3PMc24kku+Ux74SGjcZGUEsHvAY
DPtuc44NqSP0oS9TYe52au8CjXLs6o+HtUj3zUgfSaX4BmpzzDYJqyG7ZCk7muBFZ/Zjk+tuOpmx
IRjN2s4DVpxq8ixfI+eOTuy1JsRNHYK99sj8pLMeJ8qRjsKq1vajVX7o5fgKB4Z1Y9QmIgouu44I
YWcMnf9kBqtutO6CjfZPBfxECNJYBPqsE27nA2Algl9ZdkYlWQ/nkV1jkH/je7OMsp0nGpexyy/B
aht3grxJigx8gXyyxE5dZGY184vitPLtnOgwgtrIRsvnNQVe7UKpOUgQRylf8TYqIa874aT0wheO
R2MPTPDaihnDQ9y2yT3HTEyQFUUXgLPaTgnObxO/qw+1/qS1tuHeCkTWtZt0XQaj3kfN1c5jUjJA
i5dRReYSPy266n98rvA+GBi1UvYONyJlwpZhqWTHlq7f+jpU31WrXZwBh+7PoXjRc7w2oplDv6Hc
CfmWkXhc+9kGmdik2s9jKv6MnkwQ/8Fca/sbo80XBs9qdqtUbXNqV7tiHZQrOjVcgtgAOqw1WVeF
8x7flqV5PlMLxad/0uboihZXxvRm6D9R0C4yzegvt1vZgqOdM3izbOVhqsBNObT5FqEinI3YUWxk
7eAWuSaZL5CQumaUNFMbT3qv5D7DpsxFkf7arAXXp3u4OES7EB7qLXgqwXhQyOeSN71EdOc8dLWe
o7qkpsG6oWz+eV9HOt7h6J0SB6CFVCZslZZweyk4xC1xTbwMEO3YDylj0DkWHMKofP/J6REauitW
QwQZy7sp9mnDi3LfGKRSNgO1GjAxI9r8XQXcdqwCpfRxHN7wJIBf67xv/4dnLCcGZ+IY130mWi8f
mlPcwDgMFbOE8pyg6PrAwWDyIGVv7Ogpq3LNje4fM50qfKEPN//V15SIetMabYkpt2aEg1Q0xAjJ
Khsers0k80dVEozVFhkmr8PHsaEQ6aLb3BuT4b/w37N8AuAU21NdLqLuDk1VFCcnjllU1iMVJGOT
MEasH+bdzRajGA7rITQFUkuuXjpaunbzDSbCYqguSQFqy7nCDNZeHOBN5YFEEZtr1dkgTmBLDI5E
ug7q0alsf0s8VPqMEIlpZBgU4qdtI/HtTmbdQkqx1hYrnbfye94o4T5qFgBgw8r3vxCz+VbJ+vUv
NMV8QpaZuysq6f8mOTlUvuiRRMIBmBu2FHQDc3WRa8/JkdjQ92JqJtTDF54mdc6Knsvv3oRlFCVX
3JTqASos3BcGmnJPc73Tbn3vbac/B/4VzBLyu5nEUs2oXka01XoLIBFd6xwyM99eLSOpJ1d8oLl7
pt0KCZarIgpKQotq1o5DKUmP6VtlYOKKeip2rvjrkXn7ssQMNH5VkqZUO1+UKlPSsH6QnaCO8JfY
OPkwRTiGwojd76lhLW+lJPO7tc89ws/qHbwgr1H0CGkLkSQj1e6nWxfiE0DwzLKCaaPRijDpW1Hn
QE8mikmoWarGVYb+NhrGLoDm6274OXGWe1yoXlU9a6ZHWu53RCNTZ52thUl5cIcyGHMKq5/uHhdH
3NFnS6Ta++7EsQm4cG9pw2oY3+gkBH5y0SmpVuR0CTnHpnGjrJgN3mrpv5LwKTtgdnZljEC3QIzz
8fBLIsHEMS/Ma2eUVpEeoXV5r1UbEw3/hzeGxeXO4yxWjebPwtFDmM5/OG8iG8tqjv2yff0yXwc3
SqM46UxHaQ6nHznJ1C+7/DkA61QlfAp3YEJvShbXPmMYbrClyFyjrlondu13g6FFS/SeKI9uHG5i
cKWgRXhggjRP38sIJM7g7eKLlceoK7lu/4LXS/b4FdCWUElKJavAOcSLfwxw/YdAjhPCX5FmnC/B
b8mTJUqEO5KA+6KXa8lkNjaBVtMHN+gXyQxVWQMUgMf0kgD1wB7yiKi1wz+2UVVrjnOB3QnkyC/v
fwf0ddW5bf37xZcBbBJM2IAcrhj5A5xulMPmfrI+kzfQuOuRm2smX/nrXuxN1m7yKcJuNWoqRZz4
410e3mvnXc8NOhwHixrbQUATGK8Li8gwahU5BwRvpMUMAG8VFSKL2UGNAzWl1A2gmVHTtz2SJ9Ct
anWzS6W6+gG/YQ7ArP5xGz5ska33UY6yBA+BRpxRtMiubOW/P6/l7eBDllVayl+mPOedLd2q6TUQ
L5cQaQctxDv9bAq7py8+m89Ophr31teF620YOqhknudDgg2vtB1Mp9kBs5+SFls0jJwMrhYcx5lb
bYRy9ZNl2i99mKO/w6JVBwRSYLs+hG2ONj5LIQ3Vy0I8KqbFqafUBkeDJVoYtarwAbzU29yCdAOg
euJml+3uSca5n61Nd6vvaRZG1S9lHyhRvC/RS4khOEQLWSTPDmyvFLgkQdqINuZhxqr6WML9GEZo
B9AHMTUvR2j8NjNMAIYjJ4Q0O7dZxd6ttE8+Jyn6U0F9vdX+Ct6NQrnEyxzn8ZBOB8Y6trwLLcZA
lT7eh3Y1hxGvhNW2sXovsDEsF9dM6FhvIUKIdYZAouIGZ4sPrC1MEq7nnIizwhlH7YNv87M7xtgs
2sgpklNHPauln8mR4if2mtc104FR1N2omwYmKNhLmB5vmqGSdI1phGipG52g7o6gDx/IMj7d1bac
A1yAJx3j5cPB3Tye/RpEJI6BVF2w5+ovzqAkYw6q4XXpeXk1gXmZYePJWlkQpeHfIovXtULz1cgl
0g3OYd6fpTOroDHDcQU0p9pSI6tr1Y5gCmE6/qi0FXI2P4IDvv1yvkwzsYTvUGb+shkjLBfQbNa9
tdJrV4PHrvMELrHbFgrt69qjn/0m3EOuU9mZAbOGzn9811Rs5/xMP8GnO8QkiNJUseuu/szxbqo2
yXXAq4Hu/MjGvtSC11tgexis4TE65VceyL1w8hmBuNgzYNZMMAZTB0yt1jn2+vk0lumjP2D4/7/L
m11NNEWTNu2eRYrs9yl05ULh7m0DliLsfC+LNIYGR5nT99HeNeC1ShIDgUTNLueWkfC+5UeTH0l0
0KsqGyK99kgBScalylLPEhZ8xQAMRTJm/1klhXkYwa4oy2tozjRY7eoIeWYN0X+9PHufX7Mkc+3J
OxIehB6IwZgW86u3qCYCoWcdtGIhN1pQodQRq/5ydWUmiQVxWRMeUO3vCt4zppRZJRKP3fh9obix
mCR0HCLn5mHhTMoXWryRYosuz07JjTDl6obO6zibo2DBi8MWQTVpPvCx+XSEcPTQV+R8HXFzaszR
+rhdHQZhmOzy768waZJ6hnSu3SSQ78Q4YkC4k5qkAnKmDzQTjt/50TGGFUXTDb6Rb8G6M0lfICLi
mgmqhh8wvnhncYCS9dpuSdo0JarFUsZk2oDIDP6aDFx+86FlyU58mH1oqr+ijQIGQSaXKfWhpQy6
ShHmpowV4uBqbsTwktHRJw8/8UX2D8IO99ZyQSqw5L9cSrPV+cEraLE3eIPePFikw6w0DOLJVzll
8fU+JbxsZ8OoMZlmPKNIlxuSFavPp9a2ShCQs+E7upUKz5Ch0DOIhiY2wDMgV7mpf1icdOVOa3ks
jbrqgUkV3jR5EK4oVdsqed3pfjeYhFUSQxRi/DVA85oGW38zMFhn6OR08ohuebBDQV0AvkHKDoyP
Y1R0rILQQBr+ODi1dmBtYvYoIdaZHQISPmXW2LoxguivT8Q2VqJJtitGKTyrxyCzwfTN53/RGD6S
NH/YAAJW9MnpMzWPCZnzDeYUuVLgfgdrE0c2UKTVnZMdIK3PlHXBxSBIrzDwNc2mWMRvjmIUzrXi
jxD6P1zet23CE3PJJx+CgDuAYo1doqEHxm/WNqGGKmv2FVyB16HMwhpnlFkUrZXiEO0vlKu6Q2Xi
/may++Bbm8VBr4RQhsCUNWAPFrLl4i645HiVfGqzp90T6xEUhg41u/x18rgKiMX2tcpgZ11IHvds
uZN8M5+dH7Se9vAIrJmbHUFffvEnbvy8nMG7V6q0WQf2TV61aY1UwMMWuuW0KEuZc9T8JwLMSEzZ
LeokYLcowQ1HGpNHHHcoKYbbp6HIL7rloi2VOOzloxw6t4uMwpZZ2ZxQcd3YmqZt58dmnJIFlvXu
VYXjIsuT8EmXDnlg1CrBPf6GsDDu9yxa0R8467fTf7ctsNsrSWnkZeSmvRwD8sVEEU6IzzM0Gzhb
7jt6O46Mx09iqEn9fN4t91odpZLH8t2b3qcq+KcEtAd9baR3vVtRrEEncO9znRfHTGXHwT7xq4WY
W5k5TpwLvvXH4yTDuBsZzb4gLWMXOMz5kxOX02jI0eRpsUNew1Pjr9XLk+lGZkF4vxOPLOf2F0nb
PY83Vi0htT40spuw3WN6NMPh6+2mdhL95POxAow+WnZFp7+6nXWSmQUtRbezuZ+H2N7zJAT/YpZT
/KQbjGznvB+sEXBarS2Hm06BpPaB+PRDaf0uPhSu/VeRqFXl9yUx6pSoYKXTjQsYiZtcQBWE/rNC
KBLuS/NmC/VGRkKUyzTcZxvocEfEZpupYr66JzXbHpaVhIZqFFT61Xe0Kr/dIWi7+cox9oO7ckv4
y9sz9NYNcrDoUN2Tl2zIWpBd9GAX1dEYylTeGsttnImQWNDDIU+H/wxQ/upro3aXZESalWgmRu9w
iC7m/jMihcUVRWJN3zy/TzrT4AoHuAhrStOD+fsH8Sc2OJ8fzIoAnn19FNLHObMrXZZ276s/ckQc
NYu3SHyoSrebFA+6+qhoibMA+Aliqpt1cHq1Yox3jeOYFlEfVE/JEAVTg0SUUB0A8bLhI009A4Zh
GlQ2j3gaE2/5lPkqib/U7iOj9cKRFevNtEotQnWQaS8ifRPBUR00A+NxXCVp4lFfntNAYsuK66gG
H/LSTmHHjZtw537T1TVLLfWn3xe+s3UiuFcvngdCxRGaEGKMy3xrIXPv4bUSGlO/nr14WGAzmZZb
+UctL1e5IE6PyViDZRARfTpeXqE4ni83QQPnvHZphSyFdypLP6/NqFUSs5YFjGVSxyW/fZSLYDjH
/Im2pkKcMRUAX0Ei8hNcMa01O8ZZaj7taFElxUXOKOrJ7VoDVUhVQsD+T/Mma9aT444z0uis90LX
aG26fMJYqMTVrLXZg0vcQzGencEae9b+xNCbGTNtXAWPMTpyKjIUuLUGUNhGm1ccCp4EJkPy3Shj
+LVxdlV618M27kYys5XLm3ckOc59AsXCYTFXeDrzcw54Blhpj5S8gNyXiv6loTyE7f1S04Ynkoi6
qNBCEPO4QIabghaTvPXKyzQ04aAuG75S99bdnW12B5ItuSnrU/9wKcleMbaUQd0SNsZk6u/8j1EU
pXyfPxCh6n7sTYnbf3l5EGVAlHVD1ykn1FmO4JiGUmliZGSQ7WJwDUilnWyf+Ev2T5Vw8EaZ9Vk4
sCmC2IejyJGOG4e3O3j1sbp+I//dB07vkbUdXZjcYzVwjW66Un5vxfRW2wrUCVP8vRyQIbu8U5S7
Ldn+/KPYO0SviNbU/RuxnN+Ajnepsr0J20+As8r9Ixloyfwi1SEyLJ9jba9K0PPE/pI6BwAULV8v
JMuWEnqLdCSF0VxPeiv5wW4RIVypJrL69Pa2C1Jmw5e8gq9xHHwyCKJn8POqmLAjqeA0AypWj8x7
mi4+SQ70yPzisXsD5QDRqen8ILVN8Y09lAA5uFZD7lVr5s2fakzrCo2umNv07YyZUngJZ/3vNq4R
9l7rWYJ2z4nUUsB273yOJhmmfXl8gaHuDKojFq+7P2OdTVLVziABFumca4LXMW5QRKI8GfWJRFrn
h+DtUpvGyuqzS+AhCThd2HCFONIdtxmMDaGcJEcFuvRanPdsARIPHZr0i8RaeWUNMwsAhPKA6QmF
PW9R23KV5ORlRkm6/lwrmMB5jd/P0pqLVzGPClrXOMm1RAHQ1y5f8oeJvF+P0NtXNt0DiOWl924B
TWCoqTWqfFaaC2vZr09stqYttSUGNJo4yBGSgiBU246Spd0giCYVzq2TzSxyLu87ngjIPU832oIQ
pg9lbAPo3dzvus5hnl10tqx8DLOKYOBa3Ksolqlbxaukl7FCn879P1HmiE3BLNlWbj9Ym3osX6xI
pdLfgj6ZBe6JDgXFQmjbU9viLjpW7D4VCPQyZid+C4+LUTKDUZz9IKo3EJYFbBUTkOoGvcX8SlMt
z0JqQRBsOXbZPmj18mW0nKqEB09tk2jWHCQIADOcpYyDuJg9Iza+FMPOL2aUZ5zS7f43sSZn/ZPo
RnSJT1VTPKS38lMjbAD30PDhuCbqBDN6S5knVQfcrPMvRazXgFtx91WEmDIggey8qeAJD6JJZpRR
bCPNMNEtAeVMPcjRFW1wbFfkoSfVx21cP6/eh1aalW/iU4VWW2eQ1DxZ+eL4o2xfVuimAta6voaI
VODmpKr8Lnyw3shJ1K9j8h+Gxp3tOBvL7hBoJgxQvRYGFcNJ6holYDHSQM5WPM54vIuydiweAzn0
iOAEcTErWTXhRPpi2tO9LUyR/GTgU8Ob0gLOY6i0W2HFSHEbsecj/lvBAqB9iLD+jbo3RBq+vFFq
OYmvKH1r9TSQ9EiKTmDHVhQvsZOY89aTPNB6usXGZ9ZDfaj2c7PVxOnlizxqpJiE2eSQ4DO308jt
/Rpj56Y7rWCED1ef/KXye3eTIBzRRZgVz3upzhF3ThSKTfLR0QKgyTaHhJosqJTvHLf0Lx1/IBJ4
kFmvg7f05ADRtPuYCv6DjOq/gHWD7EKG45jrgezeft7QkoN9J4ifAKidZ+5Omt+GLDVzZvMq65Df
RrDu6p5GmwTTK9INzT6Le+E/hLKujuMUYJvz/pTuOhKuSly0g8GE6+h/PZiQ7IGiGjUcXFHvB1w1
A+YwQzikLPf6YhaakszUFyk+PDOSoJ+I1eBMCxYNKkfHVYzbmBGLyBhDVviV+QIyowcq276cmVwU
OEGKI0/2ZLMZ/TqHvyGA/g1vVfwIAxUZS/Win1Dr4m5uAtpwE9F1TDkzXRQU3OePQMhm6xFzTNXE
xE0wbmEr7wHbwB+b343hmVmcxdgIz2kCF6KA0XSGzUeXH6XTqecN6lXzNR5GIDjm/skfVfbPz5pZ
6iNxEqRwLqWUq3nH96bNAhb7RAo0fJDyc89pClwA84PbIwsel3WE1VgOugMOz8XX64rUQpyYU+ce
hqeD+necOwzbT61rcB3jvQMIncDvrGeK4nuZhR65EOFOMQyy6Ymb5LIs4yNd0457Ty2AmQlTnq9A
G5OIEYfIRJD+ZASpCg1rcqjy3dTR4qKgXoCXlq9T9tepG3K2XjZSZfLYevSUof0sD/wzcT/HKhrZ
7TZwlSX0e9EDZwM4lCr6X6vlzDX9gPw39Cracmbve5RwZGGb1MkDAi6Y2fcfbt1ukRjiNdlUzyTK
nGecx+EJzqdo9BOoJbVIo3XdeLddSVcuwNMX7rCVeDpmvbiPn9zAqgNXzfrAUQ5gHSVUG/AU1j6G
1OJRojPeITqSwntg+1B6dA8ALBQ9vub029lHrNFFcbEUJLb7nZgMqPTlfDc31M3ac2RKV+tAetje
yazMW6fXDX+JWF3kgtOYQMh2RSn6Tn5yox6t2hzgTqY2nuSdmUiynKgmSzxmCfkA77aj/mGZ2YVL
woXlSXLpGhdpx7AjuHjsqS7Q/Co5Ma0kFtKwQb3lSgsJGAtDwUPwormYqU7ardtZkHhuboCJHWdl
7Za4bKB0X3ObJI7ASgrdTwG8kYzrjS8+sfE6DpHOOnBMz1IWYzujQ6w5NNcRhtEdw4+UCGwR23go
ARYGDsRvv5yqgZqOtVVRFF2M60CcAN327vFeRKQ0/ldDiE6lSTPiSerSZDoYG1gISSCTHQdh73ut
MC/5Qt5Xy4PF8nwXbhnrHsQ9NaPRXzbW/89ml/G8fIRPSVKP9x/YfG4P6eBbstPfZ/6g+sAPx2+c
bGShAvlf8HJRaOQ1FPrWhpIcnuBWkzP+CDeNmadGpXnSTMISYPfukd7w3T14p+QaRRFVe3/a9n1n
8mb0V7rJqA/FZRp+irY0HkYa9WXy1bRQaRRde8d35Q94rlAnoZSahKsaGeHFxlhSslHpp/g+2yX5
0w6Y53/GtgogsMb/0xnx3p2V2IfeedZdBxSdAzoooQh7UfsOvzy3hJGHisMP/XCY3xNOg52jEilr
egmYdlF7TH4YEcM5m7845+Qe2QMPzdsslNGOtISKHDyEyXXDF2k88N8fpKW02Io84435m6UrqXJn
ccUWiBqdyrHvXWHn+lthVR/jo+IX95qurJJnS2R3QM267vDtPMapS9ldVV25WHyiF6Qcz40QXCiy
1QnugRLzMeacUNJ79hWZtqGr+OLR5iVx+K8BYry4FnP3DVlwKcFYL2JXz6yTJit7qa7qatceFSCv
r+NhWWeoTHzVJioCV0s42XGHwC7FodPGcE1PV2TR4TVM391OolLI8ej2XXbwdTTv4KV2+Mw1htzH
GRe/dJmfXgOdvn6zEp4lRH218apUwSu1leUk+rUVczXsPEvwpoDwWCRd21NlPoE40xqIOelqo5W5
8itHTTrnZ81NyIX1YwrTgCuaJKLEpV7Xn+X3XLgwf+lf49/GZEpxrj9RJxkmMkYdRGTEC1pjuo5B
cEMg54M/3zew7BEg1f4hqvJrLwX+f9V1jrj3spykyg8PmWr9NFIkoW4ShIXMKPWIfRwLKMC68mmu
4W1QO1Eon5Ttg44juC1l5HZhL4bTSXpgrLah8PYZ+sJ+hotR43t2/rlILqq9xFtgWvcIXwRRxUrt
jMlADCD9gxdNd4VrDSfhJVcS5pq79deE9Zv5Kwng4CjHNsaKEZk5biA5226r0wOffyrXblVY33e1
FOYrfEXHFlIQaO5LoerizGZ2383WR01exE62qL3alwVHKLkUArAosadPpxpHDIJf7AUjTm/2FWsd
jpL2n6OKPO8KExKtNy56NHAdH0p4nj9+1vUEDVAgHoCexewzJV2rgio4gm6yXmUIb1qs6murrSs7
mlzLd2wpJBE0RxJvBMeBQceXpfXmGQd9ylDVhLuGAppODFR6djOev0Rt+ZOR9eLpF2I25NrTGN9q
cABuCBp9csF50gQSyNrG0qUNDqeHoNN3F27/gKtg17Q4mdYGiXYfZ3GXwlKnFeZI+hzDfvf+lPlt
I+Pb5TS3uYJK9yZXI8QIQu+OII3E2sjmFJnsEr8Gb8KDO1QzxDHQbgclLk5phFgwgQuTgbk42Nwh
tNkZ82cPGM1cpUYkbBl1ZwAhoi9YJx8EzCfqeEasXncRs9pbcxtuwIZTtg4DkufFlNMlIwVAbgbg
KvXiJMlZFYsnVNoMeVel0RJqOPEIwiVaRXd2v+PDZkqeBkoSAkWB+3Li8TaVlRU8ho722B5/VbUH
LTTuvHiwjzPhfyHL8lwSqPqeBsSNwUWqa8brqc3JFK/OMBguceOLJdZo8xkxL2WZLXf7UXBpi7mn
MAeSATNym7HqJ/lbIrxzMXfXQsWUDg3NYDsmITVty7ldsyxLgR15HOTB9EwwfBx/hIYTgKk+HwAP
6tfSC4FmZJyoZAkGOFnMeoN9Dc0fWjSsj1QWjI+pM8xPJjZkjKW27C1ipg5+KShvA8euZ928cE1P
XZ6CmR7Ig8QdXqVi9RBiBj1J1N4LXVnLaHPpuC+LIZPdj5mz5Z6GEWwWoVqDxRLX9/nEoIalRVGX
YhePv+wzjSw7hgu7uosp6hgkubo367UMMFXS361MwLrCPpmrJoAjdP0V4b/JG5ZgMRQ+mHwOVXNj
2iYynVMPIl3mDTbI+dOHhSMGTMgbgYx0zPI41yC+4cqiLzjIcJPcPAqQdy+v/v4k5E8mCEUmMfxM
2G8Onb4jY0KfzOJJH09XgMLtm2Ji3T2SZ7Ms+kk9rVdo0hy/3odWy+JpU8P9375mxFich8Ytzkq+
NncrIxvqDss6TIXFwpU/Hgp+lZuf8X0rauxOAJ2cPb7nuSQbvZepI3WrEzPAJnUgFy0lgWLS+p6y
ik8lR8fDnx4mr9Gqr/UvEIyt32J6mrPMdjJ7axkoHqE9KSGWWE8CP5S5YNdcY7lsU4rLD/wOISnS
cf4rMeWomN4POh5PsBvkRJ4xrnG8Bi2W6JmL4vSDRE3I4SxpCIGQ8jomtB9lTt8nX1JfXWQVVOnc
jhJZI6e9dWp1CrDxR0cCpMYWT3iViksTIC+U2lXqpwiEEagzrEuez4w1VmBykzJh2ZF/LlyPjegd
RRtx1836x4rMTZos9J8s6W22h0i22MuFPS/a4GiH1VXTCZfJnLmbujBDCdsXR6elpe47Mf9YA9Jp
V7MbzzG/69BcE2fMfvHYLj15U8qQte/oP0ixa6eW7D7OLgVJhuYdhzpoAS90H841jo2Si1ataKrY
yt4CobCv8Rg7YJsRQfJkHLrpAXHnc/29Kkt7CrDFOTl1xtXa5aUx81Wi7hXxruNWX74cW/J1vZg0
CYiYRz6rnYZF/gHllaSqy2u6yob+4FoH70d95szHB8yYotFPGySzyO/BJa/lIX073s+TiuUlDOeq
Qti/pfLq4SPzE/dTG93hAXL3ak0HNTJBDchHruQVbL8dvbLwR86rzCXph2JbpNFKXI1cukanbfyg
4tUk2Pd/uogLbS3nVapfACY1SBdr7Fyvvx5/KTptA7ljl7v7Vsy5c/jc2yxlSIM5zkZ2aIpCP+Dt
KR22WhSLb9Tct6qAxnNOb+z2O+GN5gyyMHHRoQXpnTYYJwi55+SBiGxuG/ImFtOAM4niyB85nwEq
eXBQOK9qwXWFJvPrhyA1FjGF50U6eOIunhHg8dVi0S3WchuvX1HUg/mOmVC7TBtMq2hUbM57xBtY
cA38r+k8s7REYFn4fiuhWh2iKgDT2xHvcfGrAKCCUKgmLAgd6oesV+sybGkQ7+sBAUCfyTJ+SzqZ
dqVKQFWsZhRidqZfmIhHZrsGVED9eBBKDavclIVpYYcAV3oROIei7en62nSKxn7FO1eE9CBR9vAq
rkM+YOr/ux7Y9sIkw69ZkbYhWPOfCeRzQWkZeJMtQ9qD+M3ITcLpIZUVM9+xmTHlJTGEXb51KN69
JHV45OeWuhjnLBass57ixpToBfC1h6TJgZ94trs68zDII1wilkXwgWG8jS0flxiZeb95e9iPIMY7
yKWletUBSwifz0Nf9qC47aEK7GtvEuBmE2PP/9zOxkibep/66/mIhwLcvwNJTLcE6RJwkvZfQ2te
OwIV8n2eMxFp/wTSfywffv7ueIvpWhHxHS0ujcLslm0KDk3w1mIqt4Pci7Sn5d0vpfOR5AjdIfxQ
ha9UO6R6uORf0PhY0Gb//G8UTEorVPdHT1cvUwKLB6E98/OQE7TFceOQNifb74n+ijVSzjLp8Cv8
E84e0J4JecqNjUV0z0ZVzQDRoMsXMVy350RrWFxpaUlvFitwBZfUTAQmmJXy2IJBxZ+4/zY+Nvh7
4PHAQxVOw5lQItdJeNl2k+C5PKzibCYzZV2JAQ1MMCIoVUTrjuD8NbjRgt+uAiTq050lNpfRJnVP
1aQ+jy0O7NxsLF9RXlyhrVyoJ4gcqsOY7WR89K4aCZEFfwhSSC+Ghq2evWy0cRYUK+Siez9Bnap1
VAGSJHPFf5ax31LeypUCBZMKTRV5SlgNZjVzmbFcIUH9Fldy0CN5Wx7O8k3xVSnBqKmWCwM2vD0b
ZLXACAOFXqlhoPtX+V0hfeYrehn+MqXzZKJbgAZm5y3A3vQgThi1acD2Q83LVb/FK8yi/1EjU6Mo
prpSkE+Ru6NeCd2IEBKP1jZO/NrwK03mHZ9qoxfxGNzbc6pzQ86MQCBKR55H2JHd2QL2itJmVmSP
gKkl70KyZRKW9LMiQd2MbdHAPISKaajo70so5GAfry6H21PN3nzu+kSIZGppJmYsy6SSTogUnI1Q
5mibn2009obvox22DUe1vyfJd0lr0UtYh+Evpoh1aAMEDIMc4w92bvbQEqavVUhjMyOw7SSwpAoH
7BbUZ+onkDmiH4CEEVkNE4n6PAHv1dQuJM8ntC/IjKXFHBrYyDqCSuSYVY0JPXp2vbiSQlLWrt84
PEqsEMWKtDNbuQKAMalZV9qAppmL1izOQJfRbdm62UoLzJL8ngkDJxKYEsB81Y8wRbwgG9CRvzr2
BXQOSyOSlPB29m3M6TD4+Eunvq2HqQxLsH6xj7J05tDpdF3Lvw/ElSNOgluaRNyYEuRCEkcJNYMg
3AitUKKapc7OVLFtZr8MwQDmm8rD4o8fXgVWWe5YnBF1J7+3/uhpG0gDVgHefBvxCKPp22ogv+Vj
2MOKwy2ypxe3H3jVGlCy6K9kAObITOt3TbGeLGPmyIGRL/3IdzCaI4MN1RqPakMRz75FdbVmftln
0/RPhp6L4BsQZSr7XwAMTxQgyFqh3avCacpSIq3NBkP8PekwGXTVV1vzOnU8CD0xqbh0psMzkmls
LDcyw1hZ1xlkdnyWWQKmNiKym21l0e+V5sXUoaaYkHjAsjMhD4gkrLLMxhOzDGBfA1CnY7cYUaVh
bArShwBZgNxoSi2iPm85G5PyGJCx3MBn3tT0TAjWkvNFX5Zgn0Gxyt7Q0AJvtoY7IgDUbmFYIL2u
mYKmYxxeYoh1/dccqHKrDtnn9WESK0X2DaA72kBBFBJMrPCl4XGCbi8ob5TabwTstq+p4yEWW77+
eYGn8eOo/XhrNXuYQkbLtW8QwT0ilZYkFK6ElbUUDUOls1KXlvwpD37JgkOzRPcN2ceLSmxUFMdE
jH6Sn1k6oXLqAnVYcVXxp+B8NNzaUaSWN6//ZiFSSaymhnFKdQ+K8ZR8pK3mEpOPUKFpHSY/bv5s
0xxTpPsaLmncKY/c0wYvSY4BaSBBtCaCM+PsGAJcDTYNExLZWjSVQMApx8pCtCQ9g9ecL/No5f9A
bOAVy4ylDmaOlD77I9LLh7q1ZgQAecORwIxK/w6u8NOxJT9rxAXrqKbF0oI06Ep7V+6ugWicrpgs
K6jd+t26iY2lQ+7HwHNFpFgLcnDtCNHzKnLxrwHhkAci3gB4a5Cfy+oU6/jQJUFKbrO36TmR3uv0
dot5hLpkBsX5S2kmt08VDsKXGhvqIJgeDjD4V3RaE9ivrOi1FYrnpw0x7A/lt+yVmKkDBNLmgHUm
OLmVoK9LCpI1q6p25nPTExc2Z8QUT2Gw6TjgEIg0s9VTWtD8Z0TtHmjr4iDhUEPGjwypOWKPgw1z
85vGZDppQwglFy5oklOR6tcvLSifw1Nfz10idSaQUkwqB6jAJCaZ4x2ZeghBsff7Oani5N8KxF5G
LLP8gYUkgQEDi4LRYpNPA3djyxLEQe5GELCq50uESUNHMIJf3Iwr0FzmsQH6nSxoYi2tpMw11SB0
/g/PnvD8wO3txgKSKOplG8Ccya+4VT2fHWuMnYdUxS7AXcsp+ZG4IxTWl1M6WWtA5DtV73PQt3O4
sYURP6lyATKOsO6QQ5vpBhKP1Kor3Z7bREtyx6mc57K3jkK4e0RRqzptpkAj1si2ApEzlMLTkmWG
z8HUBPLw6ZgYxYiS3K81XvEjELNjaqE5ppQp763x3cYU84GZMCr+JF5qYCP7s1IAY7BKuFHG5ycO
zLEzm25wTUdtefhJ5HSz028xJmznCKO87gzVk9E117wYEMAe00GB8hsSyq9mc9WX6Gv7P2zPLWOc
4l4yHce7DlXDfZYfzjLtRzXdoJJiPKUVtid4Tcl3hm0j8O+19EicSfUwQC0z6iF2leGuSCIlR/Sz
yoXAthXQqTeCWcE+GhABnNIOib8GA6zFY1OFFl15hj18t+1KdYCJxi3L+593wQndigAqs5FqImhF
Exw+HkIYIgbMFzvP8zolQzs2v1n6ZFEwoJL2q2498XJg2dDdJfLopMztdPM97eKj6w9yBelG1Tag
NciSsAMrewCaX+NR/KF7BhhGaFrZ+DUkYktfc87YI03Uayu3dsHyX+Of7xfcqzAqT91C/bZE9/lp
vhJvHB+RJm3dfM+iLJpp+l4FHUi8xzIomn2ujcaeMSFqfGE34yPpEBJDHF/Z2x0xwMdF21CUqf+o
Xsdka9ExXjUfiDYB3ko+t8MTkVe+I+vVUHoXb8evBsEhXtg/7kuCsZzlI2g3RdyfHawW6TSCMX2k
OPew9aWuR4l55GrDuS+/yEeme9cRkx+8i/76DDZg7ep/6q3o6orhSST9g5ys+tCexKtbBDReEP4y
2QoSnQyrJ2kBGlaP7Nsx4K4WfEFbO8VvjEXtWWRva/x417s4lYa+Swdw8cxoPLMkRBsUnKQ6Cpi3
vQxmaYpJGfzcNCEDERRmeS5Z4hAZC9T5MQOqxIjxkTtiRVVknqWHgkiW7zYNp3O/Mi4S/5M5fZoX
/oRKlTc8a4721S3Cn4JtImrpTbXDnJ6hWyBhp0llHel5A4vFDCxzBBk55VmTO0KlNFoWzKwcBbWL
ZuEodYYjqpW0zUpWcXYVp0LjQzsukdVHdwZFHDR8S2iVtjX6189UxsVanYHqQUTrlwhwDqO7to+p
cHoQu5E9UHEv/avs5bW0ADWHTKpiV8seBiHUOWVlGpJC/fUpy9W9ZMC2rTs7v5lOGMU0cWHId3a5
sJ6Ko/UZPdX/k6uy86FJEk59+GzL47fu2rboXjVqvws4rUx8CsIbQ/uYo3wvj1FT9JRLMCZ+W+ew
ibTWdlsz69zuFOxDlklqE/cO4m9TUkAo66gIlJUGYIj5HqbPqO1DYB1caA5qBW8xNQNwp/WrqqBx
doKE5UVKoclYhxQ0toc9DOt50fJs3PaInyN3losScr/BP9svYdjpcmBzxlFIOQ+BwBG7la5MrJBI
3ITn6SIC/Dbn2e9NtGcnjntmDxRww7eBXNTRaPGa03gfsvI8ZSDYENfoVmkdBcJ9+GKfjNEZOApq
tTg1OCO0AHBrpD4+u1jo0mX6x7YEOzzKU5GX81wISF1nuMLXiu8YeO4Iqmm+VeAHAuQgPkZuMq1w
cqkFcrRJs3x+0p24NkpqWHalvzGReaAZaMDj8Pb4SVQ4E6XD7RriCMr83glOVDpCPdW5NyJLTEAv
evoSSCSGnkfCkHkOweIgGjYhNcna6YyzbOLWFe5utfo+XOPxnHrrY7dvt1auM87F7X7MHs6D5rT+
GuZSyx68ilRh/LwhyOPxE0XWiWDZCQ4xUiHpNtvTxGp5AnkUAdrnkbDbxFJwuV1/CdBOTlCPOwle
PpVOk2U5ZZ0CTUIvZEJteWzukhxk0KxRMQ1kLAPhKQsOEh3X5zGlo5oQAWyFNKtw+n2CV1KejOqw
7m1319Xo1GRm2f9vBN6Q3Ll7q+Nl1jqWXzLAl/XBQgVlt/J4VLJoqjEZtkglolWC7Q9EGSWOHaFi
E4idCqiIsa+PGRao0XAEJsm8LFKQepK4HkEF7ut9H5qQV8Yzo/veJAM6kXTdI++MvOatWt1hfpZb
3jUR1ysb8Dl2cnCqIDZnHReLGft04dmlpVA7a7p+41weRT++hWDoMt59rrwgR+d34uQuN9EBh13t
KBeiV+gDhbzt4l38ppU8CYZHVEu5mefHsEzGKP+neFnYqkJsf5ucuHvkAWe75iznP3a2StqcAgom
BS+Got+bavL1EXU+btrb34MzHye7PUBoeU3BzZD/9PEVf/1e6Xa2j0KAQi9FDm2FVbsBovAZ3DUg
Z0pPmcc+RaAhBdhzpIxi/aukajVvi4GLHvhH7i2w3fOgNCbhsuyFEgE6xsBLBbQRKaNmaVdCGIn7
reV4PabfDOMKbPm7ZruEGXE+a9xsWL/nwneQyQ0LjIUyBHvgLLpnnEVxR+nuin0oc49XU1kMxbI8
1d+RILsauxc7SFCQT6IjabtmHoXrn+nUYVp3ObNX4tfWupQ8qVd7Y55pwlk2kF77VqBusG4m2fhF
Byd4lUwus3xStGB7Am8/Y9yATFtoAfED0JJdPMAo7b1gVAXMMuKz/qbw5Jdd4rc1FP2bMY0G2ChA
rGYkbzp+4LLEJLOeOnX8fP/qJpBZ2fvddiZouRmJJ50gYbh8K9w4Wv71RswIVjuPxeAAkixWBpn5
lDH8iyq7kS6t5TYHqwMe4JH/XhDUK2SD/tLTBOiJ9diPcX2mzUOtde9EQ5IcqzL4sIdqxoRgnwMl
amFVHXrKFSAy7z2fI6X/tLQbuijyzp3mM4U5509R/Dom2fI0ft+g4atdmUyLo3o37rXrSMeJaN2N
fg7a4m2Ze7FYzbGLxyaBcaQmmwczPiiCNpbT+T0oJfFG2Aa3ZtHB05jSRVmNTwcnfMmSry+QR7Fy
ISFqKQ2Yir+Wgjicn2ZBYlz9z4PoSDr/C6FGwSrKMk+50ACVeabJUj6H3n3PHsZaMAEjFkNQds2j
jAZKQ9ZAcwwENro4qQXiLyhOxo1UFWw5aATAMU6uf8EYujkhZoRNMIetke1EE2VC4HkUMvSgXIof
Z8TkzxEjIS36rKh+sBEGzE9hVZFHLBAxCyXpEWOyYM1jmvPBcS/+gOLKpzZDUqXhOP7dCAYdzsOG
3W0mLQo8K/yG/Y4kyvuTzdeJ7pSDyC4rt8hVF4klIneYq+e2ahmPTZBQ2TFFfHnvwUJKw6XSuPw7
zJtIpp3Ki/kD/qypM7Y3xEzt5AoqytFrATEZoneigK7Tu7LSGE+EwI97joaWYx32AGVDLQJSNg7m
lKg026a/9JIJ0FXijNwdVacDtrenrMSG9eB35VW3KAdQppIGolYkvmQUP5nNlxdaNQOalR9XUdbK
4mPAjnbeLTRuGSvEcWMJLS9YbfF9b39KuvlAkcxs2pMEMavI0kD27WCMxntU+sXB55v0UUWQBXgy
Gj88M0V+ax/ZC02VbjnbCbemskXoBxmRdIJdb/C00LHBFodPvQ2eudyi07q70WxCO5+FwJMFubcu
xyVSGpo8ivaKSYcaWZ6oHEoIbXWZY49/hNlk8vTmkzxCGA8sBiHTJVUkBrCh86j+7WeSJmDgHDH1
SjMAFnr1oFddwqelRL89D+KNaQClrVzRtuE54rdwQl2Hc+Zyl+joDKXFCidVFgav7Y6pn6YVxWMr
N1ZfoWnhfy0sz2w50ZdUfPEWTrDmn+JPdrUBJwJ84+nVMlupvwdvXHtXM4VOW2WWAmR9Mz+kRDN7
1ORCz55smNaBdNzNLSx+SqBLTU0qfekmFwHF3dWsynfbONPNgvLBb5DY619guzcBK9sr6useCTku
vywovFFvB8dQgcnWymGQWJXcJ6dQKZ075wvjBKDO/spnMUJJdoLG2VBN7o5p6xEbGArO9vwtnvTn
3NSwldIlJo4zed9yudnJr3AJ/3r7Lx3KIu7Aw3DNnvQ7p0eL5Nn0K43EXTBSyXF/fFOn7N5MyoWW
tjfzYSftqLdsBRKvPHinsgTFgsx0bkPAA/S3eTXMwC244RHnbx8K7ZYUJ1JPovUWXvhpNC746xQx
xFg9CeBbqX5CnrwMIOHsCtqeVU52u5SZ547D5RPGxwhLXPljoL7VdWHzm4yFI9ieIYPCegThABKl
uRNjtTNJFCczbVEkTJt2GhMVKqMoqdk4PfXYTRN1DApnTq8rXW8mW9vTs9LkCQOqAj+2pNgAfqGC
u8lbi0Pe5UpLKJXas84kT3siMOFsa8t+pwvABu/Bqbzqa3C/VCR7aYeDy0E3QMYy598JwhabRMzt
Q2SvtY7dpQDl651NDCVYpn/IsemofpjnHS/70KVHIo8/WHvrGwdMwmpCD3KBi+UU8BOvPJSGDvoY
jNM8x8169ym8XUqC/K0Sdood3kzyl+IKQlgr0vWJYarFePy3NZJr+EpxiqD7h2y1j0mYPE2Z9rlt
KT7srtp7cTmG5iLsPTcufrsAU+HdNMgbmr7VwCRHzAqVihRD7k3Ap3aYBU6j0vpYZHK4SDjTgBxp
M9Qzh+Nnq+vhb6U0UYIQg7+PVTaGYkD7UedkjXrRtogYNDpGxdkSBEysam4ipDqLWZnmMFNq0jgj
pGBfipnUGUcnc5L4HvnuyO2cx+jpJQSxyqjP9Eeu25Z25wwdaSMDLCpPOV2Za5YzW7cgpZbpJuDS
mwJEl9SZzCr02A00NFnm2Q/2LoSVLxifo73oXJDF01WqvdaA2fDwSrGau6A+nngOjSSswYpmv5Em
7SnMRkM7KAviKsdfAiQvgE5DXsnki8FP3wj6I86wH1YTV29nvzbM9xKM4EpjbXnpNXVef+JOMZuA
eg3Vgq+8PIuU8D6gfLHpoHPQsxsC6dDlfxlh9eP/zogx37aHtEVAzzRiKK4NyvRjLcq5R/jfFbwi
fh5do9tUUWw/2ZrvV6bD3Pf6kxJql5K6SxQE/L9kQ507X98v4fsZsDyewDE53wQid3dRD8SOPToR
emH37LZ+tpY6/6TYCIGcOLbSaTbBtX/ZvKfxz67WN8az0kdLCeWpnwnQcohBfqVoDc2EWrexhfqq
qxNmMqyWXTnTQqk/W2AmSRFW2wD4+J6wMBs/pvHNMGAC6Qzo/eFGunhuo4YibqpqfXZDpPpm/Mzw
MfPjT/bufkcN98PZinJDNidTXHkRgzOGA/sbOJNaI5Nk8AAnhh75Ymx0pEdknUkAORfRgbL+gVH5
vJqGxfyjd6rL0fvhgjdjXGm8gComniRfz6RP+Lm7OpMqz4+kLdJ9dd2aUjCc5j2Lxi7VFI2bpus6
C6zFjS7pPwpcyNWRRh7bDo/UzswCe27WaHPZFRb9BVFpjfRjsxOyIJ3jxeaGgXJ/MniYzGVKYQkx
ry4kwtT/bPJLPt917isWO5/V9PySSve5cPywe8SAW5lX6MIEAiPvw+cnBqYz+Pok6waQGkH3nO5a
UmDfwNRGYGe/uH4+nCcNvN0i58PkUativOpOZtPoV4ASUBqxuEggpqELtnXQ1sxUURKrjgmHLywp
kRSczfJcdingig4kZg5K7JslDj3XCty0sWIAGhzSg+/WvP1GA96oDl1jY1nSXFXJYdTqkCurEXvl
QHk3xhOucOM13mql0q4paxJo3eRE/BPJ3prHf1JBuYzfIlsWeyIkSdsblBHAnzmtrMX0lF90xw/w
Gqno1ahIRLLUHUsD4N3dJP+Lvx66II6QR/S512xmjCS5fNWjDk8jtYKAnT3ictuUv1MNfohT9ULY
xhtU/VZgbmb+x2VO7L19Ui2Ls021JFP0Ua/QUGqx3cYhJcHuaQ2sSn/cVYAhbuxpLpcGIFAKuY5b
9NuYuMkIX02sbLimmiwgUt6YR4iVtwCMiiOw91kNQ0TlpB+pfZ52SxV1ogql2Pxv7BNqsoE5fXTR
LLjRFJbeBc4OZMSvG10hu3B23LAt8LmiflzmQoYDGJo//EzhYehCaDoxCSyHit9ioZW0kRaWKhq2
lmuEMyTPcKMajw2CoVx69F6fXaxJ8SnJqHdvCb0oBuYfkBpfQn2j/QkYYQJe+Lc2tFuww+BcD6Dt
AJemo2/lTk8ycHGwuMov9QYENgaX4/rsjBh9pwtKHKgLBQkLVTG2LOneXuI/kYcInn3MlN+h8gPR
JJ3fVYwW4fqKPzPJCzxq8pWOyhQ130gENeaSeP+ONEi0RnHl8s5rXU5fr+eY1Rz7hmS094FjnvHQ
cdIy8JUtGXgp7UZwHECP7WJDdYNDy69WzlNBzYawrBdXaerHHGfXuD1IzPR91ve5IPXJoKn9OptG
RqLBErCR/7mC3UWfLOVTNYDhG+VrXPAHMdveDtKjMJteQcjsmfBiew5r5itJq8RK1lod1ztMLesK
MP0wGWRxtrEtjgKhwceoT9iKTGA/9uh1B1mcMBcxSOdsTJQNNyAeNDSSlxmhccwRkO5TGqY6XcpS
wgec0+lXDMGeeOkuMXyYpsQm3mfkr6UvgJQRVndUzHK/dam0Kz1OmCVU0zzHcUI7JR/uDxz4Iiy9
m+zs9BX86FPiJTm+QsmFO0gFc+B6E5RBfn0s/TXSqz85n/zS/SKNDVLgfRb1yH7xRzRsoloSugXw
J/RYF5rdEXt8v5eETNXrVIvtpgFYWvC84xIHAQcBsx4lylVUNQQ5dzsXrsYPjFtMQcsuj7SavM8n
xB7Zoyh71Z8Oi931yE/Tlej/Qxdm7XQp37qQK4JFQjotIO9mHhRckp776qQLsmDHF2LEA/6Ux21R
pFRTK49eM9pEVIUBFHXMzOZw9Rvo/myltFvA1kYxXP3ZEF4MpsGcBpUTFvtJaOj79TRfvQxvkagT
EV38S7BA5dOYUghjA5xSW63fQyM8lFESTIccBsDWhqJzaZcFfw96XMHO9qvVWFPrKNKDafo6hi7M
eEcEF/iKC2tHdjUHLCZQZj7Fkacf2bs39iM/EOKUKuxOdZJJ8XIfs6LuKSvy/IHnKLDRllqBwTHm
Fayc2uWM/6Qi+yVDcB8KgglxveyPTqiQVPuzhaMDN3/YtcYdX5RiKSR9P9sJjoAnJqFzZwvDhMGK
8OVRB/eiWiAwfXBoYRI6z1IGe6mliWyBzf5TtJttbA56hm7NL48emkAPwrxrfn7BGJwzf47Geaxl
rsSwCEJyeue3i7C5+pSlb2yMNiUJg7lJBjIhYnxOTbEuvHGkj6cjeLelCAjkTjXNBJZOtf1ZBx0T
mAY3E/pUP4WAIsCcqiP+4RNE1SToS5/VvVm/jMlVmhXDa4PITHVYDFalkvELirSJE0ZMsqdfRz1z
4Y8XRxd/YFH/OiaelvHb8yZR2FpS+/lV1xsD7bJGapB8sSISEVfLNb2MVP/z+ytW71ZUixjVy9kP
NerxoYZwh5hzgnWERlxrKFrLxsa/kd9X3S59vF0fwWD48k5vGDZfSlmejTdMJ7KkNUAiBqGumPIf
zsm7i6ctDec+mo2UESE66ukhoYLR2W/o6f0P5co5pir+Sv3osqjIOtqGoM1DgYqjmbUAs64btLTu
uWfUbtlmvzt0iWptw+fR/xlRcp+Umbsh6xn+hv8bJfU/zBwL3/9QnyVsZFsHrL8Q5CfCXmnbJC/P
l1Nj3RqAkYzlUVznIH5+vZKObStfLM/O4MkLZ6zENiLofp/VtjNYRwuYesaxX95T7WEo0SFPlsIa
OejtvyeGlawH8DtUQHziEqVbI1A1FsFzOXxI4qTrU5hZHwiEmOq3FKK/1540milKo0JshhzVcDvB
ENSlDExBHixlw+9H7+AxYXhPAce8J32rp9tSdoSwGcercnpPoHUuSQP7QQkWIv5LsExKsk80KaVB
/3S46d7CPm96Nud19z4TmahP+XX7AiXZEPiCvHTp4ea6Z942qqOgr1vPzObH8C+sLRJ4VP6YFEwX
cL/LyciupW3p5yFjnu1RQnjMYgNaVkhg6yuFaBTAXaddo7skze+f1gxsGJV+s/5+wTpSzB1F95lR
HgnL9y4Ti4AlbK82E2fxB7lHjkz31btrwovufNtAKWoeUU2NrjcFLWpR2wnkYN34XnU7vZBP7duR
xHTmAhLixpjhFZP5+Cot6CRDIq+qFbwlqUsyW7ELWlNG7kEtC5RrqjVs71KniWfxoJffmdmXhctt
wNCGo+0A79SDQwM7JfL55mizt8vgzgEkoydmZtvRS+lK/2s2ugetscgsF6DP9YSgDnQ1Bdak+cRD
NmdRb16UMkcfTr3EBJ85OKTuwyCiokozuYJ3hO36ZO6pAZAoK3Iz6s9ip9CCTmDfL76fUT+adaNm
XyyVblihzDhUHKR5QgmGugJlywNR5dWH0P3GZcU38KnCN2mdnzZhol7yuUz5DlDdkLAkVxnZpJs/
QTPOhgN38wTpA/svJ4mAhDfQ+0gyrqINnpiP389oJ6OCX9JiZbbl1Lu+ZNBEmi6k0uJ7n7Apmjd/
XXInsIwXA5LneV1rhVuWCRH3uUPTdYzt6yDZCo8/1w27HeaNpRHbp3eu46xW5fmCIBOqBH10RFVr
38zEPwv3uaGWDivULZwCaC2AXxVr+h7Kk1KbTZsMgVt1UB9ngaaMoHDyhbaKhT1al78DfISez7fV
YADtxuDNUKgolyzzga6paZ8Yo+hPjtnSoObwHmSHTEPYN3WaeJ75pg32wEaBOMq5Vo1wgQ/XEh7G
GPq3YO67TYLOFMjdi0wCtBPmNKW2yvx4JQ0+/9uAIoeoe6qmLHc2YmOabl3YbgENsAk+Tr8o8U2h
TFcmSK0Godg91D24qW3ZHcrQpqqJntVmIu47Nk9iHttCfUI2Xrw/emnLW0lVKkWBBYd2aONH0cQi
rYFBXTtoTVDZ0Zxziaihp6jejlb48wxMoHsuk3LGbxMk0UcMO3gtjZqgRUw8VKnHnEjp3Rj3fSBI
GHaeVx9yVQBCQj7JKZ+RvRlpBZ7fCYRUranzzaPGDa86iKSN9WKG3aWybxOXUuWVfXOk94TK5CaF
eUpmv7QDuZuABS5rHWkRzkyV89caIWWUGGh1usgXLdxmiUxdj8zm/sdFGOQL4757GlvyMpqB4FVp
nL8C3O6prPJD1g/WWawO+0n5yCWyJHLQNl/VWIkqh8Tt9cBxhpxAjHPdpKfN8jj6f2UMu3SmmEcr
ANfjgAhALzFr+emsB/stt0Sx9MEc76FVdwz0CS7M8OO/03Wnt/zVGfHZsxqWZG+jIx2dn23Xp0k0
hPRsjFf4qqJfJFe08Ou/UMdJoFn2vgnLcgGSDV7oHI5RxAx1ApTfARDHHndtp85WzF0Mfgi7iwjZ
wmnscP0y9db/nyvW08bq/pmBXp12oFWrvvLAk53k+uJy2QDLrU227kvUJ3Q98t4DotEyOXzJ1PXA
AZiTdTDwpRA1DfKZ5+cPoKSFhEoqqJHT5YcD1uKIsJS74e4vtlnKpsENrtP1LvDFHpCl2qiQ8PTB
f5YDWs2rRYWmstzMCGDOw3MMH86bSDv/Axxpa2PjOS/4UAMbsUmB0vVEiDCPdI8UNYQUzoXfrXPp
phXYEefNl7qtsEkNCETX+9BVkGYRC9zGHvA9Uv74l+aONhAWtjuUGJrliKvVsBQ65fBUa12nGLtu
JxToQt4JQPxDngK9eFVflr5TOpkFAKl6jGtPA+IK/jUzetVf765ZVMYmfwzsNMdd0PGkvasvFEbC
F+/GXlSuRs9vsiGaFea56YbFcAGbQGghtGIsqalPj81Nod19oRfKJdhy9KnDD8ZeHxGW832eLjHq
+KTAn6+XSkdzpk8yaNz3XqVVuDKKCBSH5rDF7vKj7SaJINP7AngRvjkol5v1MoLehYQyzSTawh+/
/HhmnPzZL6CnRwUFr+CzoXtDsQ6HEIhkWLA82pn95VHaTnWRLfVEHBnEOjNccXvuJxaVfAnJYdzi
fzQEhETq9Kg/tK3X89ugpCjyfppkuGPcO0xJAjpKlJr5JQLLsrTdoA6wIlEtGNeM2yvKpBom5/JX
Zqru12aDggW4b0jpobSlvnKm4v8oaVmwTGIDaO9u/Hbps8lswtLseg4mW+k+uCagA6+Ydwib3r2g
/7WjwOt5yeVySmEVzLfgEreSnXeE3Nrd04cfauxl/Mduk6efEazU+/VYf3oFEuiGfrM5RNxET+Ub
g9PPsGvoCvWbqJTekFxjrjjlxBvje6FLof9gCbHCDT9G9aaeqV/nFHABkLdeYsw7U86nMmTmv2aI
KbRtoRYT4ZBNaykibXff73WIqIDoIemElf/O7ovWm24yP7jU2Te9ZFeDoBoNhg3uVf1jP/tcwVEX
HtMaawvTgmd4LfhJdtJozk6SOjFr1CcCdd/G+KhpegYxPIraJGeixXfLTCwl1zc/xhPPfWNXCJwC
MengCzSSMXaadktN6uC+7uqDOukjPkWCQzjmYzUgwi0epRb2h8ggb8gLubYrmcHWZxm7FlqsJrg2
7VLs+lfRb3fBuwWUAijLlaKNqjaFORJVFspZeCKHA/IvHBYIlh3/S5IGbD8T5Y1YxUBsEDcY+5OA
FHHGpbe/zLL2T75NwkQESqIe4fDUCpSa1l9Bev2mwmUSdPveJ7LekACikXbQpk125kkQy8D6Ha1d
Xwm7DXsjJGLNtJNCiNpcvNUoyQYRvh1LRZKSYQE8rgYyf4j6iUEp4ZHQvoMh9w/W47CO/+AUfu2k
zlPWsJZUmYQLZHyCcDQX+RT3vVSCqIcAvlLqy7WYJSEEhVJu4HCQhxEftg6lx1S54p31TNUBtEzz
L8ZbJWBHI3bMzB5RKgHdGg9H6weo+o7w773tzJoe7R921hHMM5LVLSXOEIBRzSgDr+YucPyge/XB
p/nhIKwym0s2Jw/pBApkrAR0rVQIb7aXD5Tg44eGZO1CX93rU+cFG46nz335n8jwH162XDHLqlAI
YWbX+eTdkMwgKK6SzJVSQ328Ph2cC6azLUJkmd/iY+SCdss8rXzoA2cKfT7hInfE99pKN5NXPpH1
c9cSaCgOKGi9nxhigo5qd9Pdsqa5bh+QkrmwiTh5gn9RWKWkePHlKBdgAbLXiegYj6mv0NB9ctm0
72GaWDvowsXkaI7TFIRXHwG3LCv4y3CUkK2FyP569TjajfObixA2qDPcJ/6EyhIuh0Md67dDZsfq
il0oMEwJ7zwEdjWBPUZ39ps5r7L/i8xqyLkuushN2dN684jM1SjkRkLX3+HRPdBfGmgWtqMw+MDK
pJCmCIi0jm9YCxuzH0jxopQKp2/9EI+D2pRfdw+v3umJFsBp5l5Z9AunYtIc43IhpxPISvEOMihe
tl282tT+Og/y6uyvkDOi6vc9Wad062USOGDuDCm+5qRWiMq/DuJW9fKjsoyC9ngvyHFDV7F3FJ4Z
jkKmAs3EyHTmj3GA6qzR7ak8fb6cH5YaL1aboWX9GCo47UvFnKMYpIB3ZZ720VAD1RI0CMgv2uEG
yUWl/SakX6OSSSwukvxWUhfe/5ZH7d6twKk2uouXRwhoicES5dYlJSmrEUTPmOj/s3vgp+JeQtDJ
4eATJ8wb87RFbVq1+6dXov0jXWdvDWoof6bgvJL9b21gOrwDGf1q5NjP+s7J/HnH0nPq3KEWVjah
JeV7F69Ce4rAN89XUs1yKtp0Ek8Trv5OMbrK5b5ARf04iWo8XiUcDI3OQzFSPO0sjnO2EAowLR1W
d2xyZQ2m6npDmmCLE1xMmE7R+her5H1+9At1sbWcN+APY/kcAXrs+nJCAyJckCbfVi+RRZxo9I6p
ZzTXDVhN25YGYby0Kr1NHYhXUR1huiYNEczDG7upXc4dObj2F5N6FbIhmKxhWZszH9t2IpHfjay8
QhuJdML6NNy5yBGLvwM4WrTWhhoaRYB3ol/BxVtoZpimcy2RnnldB7EwhwGqUTOd7Cljiw9NxiPy
IAurTKagntTHJpvadOeicBcOJKTgHdzRyobdCpASVwnpH0uNkcu8j8Ky8GZlEvgjlgjUWVTUIpSr
CHXhbj38xiGE18PZIsa78eElsWQGs3ScpaeWpnRrfZyxwRN/EhmHrKGFw/g7erbH6TM2yjGR2brR
tMVWIHz8mK/WdcZHp1ISLfyrMKohlKSde5OPQK+7JsfEnb3ZRpzDZeI4DMWY4unh2ytHf9B3Nhcs
X4rehuiLdtMlbspz9tp3x/MTwcHnMfvZpxY9/D3N5h7KN05XAv0C3ZqQhMlardjBxyRA44gOnl0H
rquiQMaXMAC2T3Sdh6aOipe/+aZb9YNqHRs62Qs8u3EtpCrS1h6xYkRdKQGFgOOtr9U4i/HBLS0C
S4RR2d04TmEAEsii3zzojX1S5u+zrrRzbWlzFp+BJEF+DS6DuWtyfqddU4jgqIX9n3/7zAE8cGVU
L92rrhvC9sKSLGakFRnqNjGjh7DLg2tn6cNCFhmPMKzSP+1UWWpxizXjcVC894Z16i1u3FFASp3a
3dgD27UNEvwiC6yr9wP99UAdDfI5vhgulPHIw/VbOaaOe9lmTIjNWPhGz1EUfYCIExeqFI6i/n9m
mEWey7uPpTfveTOXNir19t/ZXk16zlFOUeoGRqcp6D2z/Vulrl0neDUH9AW9/UTc/05fHfrxijxx
bl2dN6+mxZ2PQahWlvFNlpkKfpug6aRnCSH/tytTZVrD0TFZ2ZCmLTd7X10tOkEfnJMjtWS/9eOr
Bdthd3LCaAhkKudCsWGRC9jq4FFDwVZCt7mM/RsmaE+tXW1DMhXyd8sWuyPZFcuqMWI4Q+mseXoQ
2YjUMnudlWn6p8Th62SE8aSvch9S7tlGmdTGM4yY8cAGTtDGEN58mhyEs4LVv44gpikXShRkudrA
yP95oFp/EKSYPf7YYOo/2E6hgzTFvBAgo74sV59mFjYQZF/fMJXLhsAxpoFp4oc7REge9Gf9EbIC
cuAukRipPGfpzY78PoOECEdAqaa+ltpyPXemWa1I5q7AujqjqZ+IvGFV5crPfHx/8lejMXgVjb7Y
4pBlA0Cu5eIlJ3DiMbKsf8J8Wro24V4E7+eA2CcbD3Suikz0aqHPdU1bBJ5XZud8FBkppkR37cT/
HioiSdolbiT1k9xy3yMVyqEPV3iQiAKWcSTOCmHYRHMSbrprEoHhCrHw5C4PiL9FChJnpZhwOygu
CUNhfK7078qe+iso/7LtgcI8cBLklnQXpdwBxr5CSWe8bVH2LYPuRVWUuW/qzZAMCtrhudurcPhg
CUKrRnbY6HB70MI9KsHDZCHEJDxi/b7VjyfqDOVj8RnjTpgh0u8X+FuyR4mYF6Ose1vY7+uaxPXD
QIpBugfnwC6IuM2gedUHKgwsNtnW2HaqYPH+2TH+j4GvpXrioX3GC784X+1x1kwdOoSF/2mKI+kX
a/quD1J0TcUgF5jG2wR3GAjukhiw60VD3yvvKTmWhYyEXLlIfQ+5sMCiiQygu64+yaRskbJVg6cK
m9D87cAF9JKMB7T/wpI6tha7wHJb3xgR6E1WBYkfRcW5rluk6Q+KR/ckMFdjpmBRipUbKw5YdKcm
lyMse9qZFg0clH7AcGL3p3eZzA65WjE4AHx+rMERqGlOdITSC3a/ce6kwnvmECBx+lkSwqsf/jQI
yTzcowpPfwAtS++O8K75s4R6v1SmogoY5ToR1yXaNjv34d1DACoM6PUuEWPMYdiJmTIRFADAj3WP
w4DIySP9ZpYURgcYTiNSKR4VOz0V9SKAuAC3ABrCHynU7rDDH6B4SQK7G6iS5KDYD2j/pnSYM0gc
vO5/EXWNvIo+tA68gvXuw9PlgA/F1gIfy2xOQKJyN/J2nbCHejtVkDKCu0h9gLyxMm64ReHvGz+k
9szZMGF/WedSi0V6iQqF8qWmUo0B1xdael+DUhSTcNPi6GULwh08pa0t9+H25tDvI38Cdqegiehu
qSYJsKZ4B4WgI0v9xuR8KutpUXnTJvk/5pCF/txD5a0T5xYQakMkvXmIvly5AAexHsTr0vk6M59Q
i12AVQq1auOJWh3iiY20MEG1s1tnaiOsNplOzDJ8wlna3frlZj1f38R+tt6Vtxjc+I0/4Th9bVpn
AS5S4wrH9tUtf+KDFfR9N5Z9jY6kH9UOSXoHrh3OmHrDFQGQe2OdDFZo5MIjlavRHlnar9PtBFVn
vKGDkMCiVozEDWJh5ojrqBX9NqKi2MOMXqeYkqXS4hP6YVXr0SQ1uUfj3AxUQFTgOW1GG+qkNjsl
bSJXei8dxBhQAMiGL2OnyYvGWnuD3YvMnykQUyvtkgvRKltUZHs5Bwg+d+839uDxByNCpvfWv5Mh
hH30PZZxxb2CJinRKDFIaUETY7fp01jCqLOkTrvjAGoXWG9KehfgCaV4/9xZ+xZb0F9Dap6zAGkE
AuFOCNPbeGgZoV0JDiomZhXner6rjs4Dzj8kxhiAyUTdIuAXdR5Q0vDeryD9MZrm8RX2klFiw8df
MfNf2dBCC0kWyyukCim8vROFKlna8pWsDOi6pICb6+gXWB4slxYr2udpJADzltcCUm6JnVxTyNDY
6tVNo3USzvKYgA04KcGA4YJg8fOIPBJ62hGVWd62bYtJI9xoGFY+f0SIJ3ynpfqQ9RdYsPBxCudx
CvbkcENEfpVAgIwqi/Hg5+msoDI0gtwUKJUei4DsxUXdNoyTX7hXtear98TpD9UWyXgNmEvE1EvF
tUbZd+VtiHY8tgdhrYqQXS9Z8CXletV7VEtJHBsuMgeNnDxWt0jfUOTtDewIpqIg3YMa1o0PuwlP
B1dUtS0E8g5S/OFFDyTda4PzwAPX+R43oqII7UlQqqzTNleOFuzK2hCqedOc/Ixrzytt3pmvQ7Cj
dptR0pvVnea1thD8J9m1Jzi6TvOGJsLUaRLsRMl90DSQKcv4m6fz8p0cFaD7/Zdn02SFkFZqVITl
cDYAr6O0KFaTIheCJWSbee9LG+l9UI6qpryZmBH0va0oqG8APG/4nBMvWWgv8iUX3HujwC3xQosx
yCtv6FawPzaZVvEhsDWguC3IZWhDQC/i+nDVSn8cMX00ggnFroaeoC00RyoQMLkA3dlCBAWPSGCp
6/n35mE62z5DnNhzM0jEbiiBsec3jiVrRx/5xRXRfqknXMnqJpScpWSjEQ9qtqOp4esQtOi8Pn3t
LlOfe1eydD1rHzEbmgRGYDRTHdAFg5r/LB8z2puPm5asTM3I/RI3WM8apSmaCjak0AFIKzg5CilE
Wa41tepTkWG8LR/Q279fTWZufdYJHD9OYun4z6SL77FTUK2GtIkteZ0s1/Bxtp4tJkJwWj4x41ol
MhPW57WQyaK9HPL9VSkLuHM+C3u44WKg36zL0BSy9GQAfCOZSvQ+9JhAOOeMHfG+TJ8ceMB/wNH/
4VmnD8ltr10siA5EAiv2wkG7i6OcCK/EUEIjrLLMwSocKbNK5eBpLGlM9wViiBAPDh9p/O4d1KVc
UJBJRPFrSN/E53lwJ6eeX8H3QfRdnQQmq2FD2kqveFyMafwMN1rvRciK8l8J5on1Cavu6K+JI3Ks
6V3BJzbXd3aMsFa0c0nIkWbHM1yhd8FzaHwu6xcp65An8LX3eNX2WulT8h/tNGp/RWPymWDjqGwB
fZBsW2O4YVE/dIFkuxO9sxHNQlOJ8h4ZqpsINNwN82vmmeGCYZYUvMMTgyb3gNSrsEzwnpPfUa9b
r/3CMEr+hsH6KUhR3kdtund5wr+kHkDKvpvdlu01r3BwtpXgG5aDJGGRibS7VLDzouvTYwmddimW
a0iyQZID99RJouzxw7X00K0z0onLx328k3NgZ1vdPesCFADex2ZrP4hmg8r/yNlrESyc4eTGqVKu
/J9TmUZB1JIPxTso52FFLWgZUYuxm3W4T6OJmjzfSZxHm55z1p1cQh3i1U7U/Je2iX4bmuiNViTU
PyfojiIKSojamY5/oHEZGQx9w9T7MmwXHIzb7cqXZDBE9JkPe7EhGeBZn5zjdcfCWNK9AYl9B8UQ
wkms0tdw73r6bmnRxoeX7UhYUiBvieyMgz4QluiJNeZRdUlweypk9/lOmDikYvFDey+R57zy39Lo
dSoX9ExBlGAOoD7g1QZjTwe2OnmYlz/LTQ9+lZ699oHn8YmlLk38/0iTJk014tO/h+OBfNnqgIJE
SGdWuuB7kl/9VWSuUQR1wvWDW0lJ1APodCOe7NNFaIaZyo3KWcvcEpP5peJr1fPE+eYLSrfisnow
j2ff/GLdefYN9u7xWMGx2HuFEmu+ct3DrIdxOZbFlg2kxPZCxsiH6tA4hHjAvtLF26AugOBilBUN
zgAVZwzcJsHk3Ml7owRsoK0Aw72VFoS586tfi35QVX8x3HtI0Lzx1UBwhrcWe1ElAVcfabjCp51n
heMASl9ztEEXR8DXiRO+3Edz+G7zQ9jQpOqqutB3DXqFwY1Y9UcvLP3iIGjtjCIkIoSBqeXncXwl
rfk+UU9C0CCfEOb1klRNsZpA/2Y3ogHj921TO5Dys+QtWE6sa+bIfA0V3NQo9TN9uyfQ96Hzg92e
dHXSEJPICJu+RBMGzoWtbah1nvMBPMQpMCuNwc+IRYxsySiB8/cVy7PJOgsliO9uMnwEjITWrYtE
098NbEvAJdHM8fGkh8HbGp0GkGjDpXKtZa9UpOuIsT5ZXE39G6zdNNpwbwLhVY/y7jWk1bJk04EH
1GcXs8RK3iNYqRWb2Zem0I9c6Jg2Le2FmtKGsyWou27GnhMCjOVmWFt/4Ui++bwXTrU5+Ong6F/1
ajiDgf2qmcZpYEYxUMWXbF43N3f2W1KBWzG7ZpejnzquRaqrjVnKs7ajHkGhE/8ioikj+hjiB/xC
LofCrZ74ZC6OaFSIHobN9VhR9uF7uvyS5Pm169x6cX1FhPPaCQyurVYjDurHHvth13cUPLX+4P+Z
WzXG0L7ScRYMShqfTRCWPauyYG5dHWBrB+cRybxVt+MoPWcq9JE1nx7alYz1SoGOS+JaxVP1/YpM
rp5pCKzb1cfccK+loMZ39KtyeP2tBpjeGyVYkQVQoLKG5ny3tc8S0MplMDeM9T6vYaIW6s0p9nKS
Tx9qL3iZ171484YL4z8pii0n3w1i9heoLTZsAt8PIftkfjavpt0+PuN2+Ng7OvqqjGPDngkGNQk0
m14iRwtpKyp8r6WwMAJee+qI3ZUCXqrg/+33ENjx7fmATgW4qOMaNS141H/KHCKtvQJy1DpzDR/8
hqVbUUGPfWws/USvCiFSzJ9CvU3+sUNYClvneEik5F3jnYQguu0Yor/Z+GIVfJs4LfftCJ1Xs637
IoRx+1vHIoH5Kr2373mPGEy+DCPwrkq8Sw/7u0Iad7BziCXeZKCYYugsev9toYg0Ol9/9Mp5ab7+
fY7rkSfqLOuWQGObR4GNX84fmU/lEwuopoPFbR15Ry66jqp6UIR+kOi2n+QHRlHhdnVdrorgAkKy
hM0LWvL+qvpLrOyGG8x5OuO5v1lgSTWV4Up0NQK8oydEW66Bb0qg3i/3+sgwm/WUl7Gd8LSdRuT7
xWCopqNai5UpeZ0N9PuuR04jbMKkRUZql2PQTdjpzlRFmIJ37tqbwLfMnvn/DzuBKBaXb8wo6drD
JdsxozuO1MwxOLS+3ypofK43CbG/TAaULpr17yMu0G8HQzlCYsgcYT/OqTX4ZvWIDiYxXgszDdfW
KASI1BdqMU75rNakvnfZ/RFAPJP2vgj8WdXyGjgdygFILmo7V+DM3vrKNxWelwBtFet1DutPWS2G
q6MtMI5UUQHITCkP4GqEVowW3nIwl483IzfDLRoUFEnikfdVzN5WV1dKcoSv9ylZe6myqPmB1x07
amJZ+yUiPkyNswdCW8u2gCtbV1PU7XSRVRA+mzGhN/KTSzChx58jsJ5kPKE/BJUA8Wghb+/r83br
iA/okr0o2YHnfMT4wmbaGsdlOPSUgnntlMD5lNCCu3Jl88mJYXH6iPGEGZqtMg3oLC0ZjhsW+lcA
9ER4DJ3/ab/9rZ5U96Bs1MC1pFLim/Z9Cz7HAjlv7QvaSm118WsScIVfKT9KpfobRXytv9L2bCvH
tpma37z9uiGr1u9IaMovE+BbgN28MwXjR0hMECRBrnsojUxqfH2rNIOv1lRGGJFLnvodjJmExTSN
DDREm1A5WfuyHS2VB43ChRSS43DkEGJ0NjD9PB5hAudfeOkwVKEfyp2b/aSgBpLBgVmofk0tprf1
X+qGkP2r7oAWSiNQQ+btgMpai78qQk0IjLnnS2Gy/TC1X/MGD2YUhftjHZU5XNIyY9L0m6Sqo/AU
oQLBat3QCsr0aJFb+g+xvXvAWoLWtCkxc4FzkzzeLwCVzBBCjxGgh0PmQzffaCGUlOOB2YGl9RgM
vZLPo+SpgTV25/irb6SOs6qu7NUGl8MgTCTZrkovnb9LHDsJGa6nZbSFPGQkuzW2fiIdqIDK9KSr
dHt+kVt61p5GfieyYqp8vGVIHB0lj4yK9c3dljK6SYLxhP7yzCCtA3Bdbw/KojtOhpbWxf9NfsMK
ZVmg6eZj0Z6FuCyOJgl7IRBbzhGAjgyTe4qlZanTE5cVWq7aVgfa9ycu5IJ36TreVBmxYEdxmk31
ghJrdVzROYAOPv5LWW56CB0mdumDv2xRZ862CMjFKIu9XUkPTrY6C4+zSOg5ISb1D3ZX9aIEHpt4
l7pGm7LHc+OPOm7LYYVE4D3ZVkiLPC1h4AdESpIazfWntkZaM6ikCG0vMh2Oz5XLcjx0UHnOkKPs
EhYoVfTwxahZbZ96A7JASngemGoHPsxjz7wSXddi+1Rwy0zV9f2wI9kS2/8XWmcpVMGTnvFc2Y9g
65KWDb/+Os5psXP3Q9an+MXcsvwXxso9zpE7v4HMv3rOfgIYHiFcDvbcnAdWB1uBTVAx3m5lgLAJ
kwB67IlNn2XwhsunafbwHKaZYxNGd+g7SBcK4g1XwQt6Ayo6PjJG1W10PA6IAXQyFP0ALJcs3StC
wuWV7NhErOQTgXFli/iLrsBUO2NMuGAlqbtdTYeOBN+dFk83C/nIXOueKva+Gy6iSXJ97ffXfEXy
Ol+fidBVnpnoWSSFS30xHVkkwrwXtW+k9U3erXi0kHtJrIJRGx/g0eKARtPDX8DlOopbL8GbQyrl
Bq5psckJppts2ZbZb8D30o1gLBA+eIlh2T7Cso8FgGAskFs1nLqIPGA1ZJ32XPQrNmE63VmEbotO
05MD5GpVM9jyMxEc0quf8eAPGj66A9jXyMngmXPy3YpN1BU3LZmmif+eX3cEXaAihoC5GA2sVzlC
xMmx12M6yC909Xd7+mn8jMBComJh/wiDcUZod/KpmTb/vm4xPlio08I4WKeuU1hOz3UCYPbbQSqj
pKIm4aiAOqN4A9NftCHzl1zTQXREJy/TtoNQ8LGmi+DdFE7Qy7d/fl/6n0A0WWPBEAD45BhRU2Zu
6Sdy81lXSnG2EpF4SSHzG7gufxNeTbE9sQ9yO0TOdjArY/Y4WTWXwgqQjiM3eBdOaFTVErdg4K0p
+lNX5v5HOfDRWdxoGA+h9YB/4WgXnd4ll0F3uUnp4oYrQvfRCzs7OvfD6BApwIE+r5FeytfeEG1+
AgD2lPFYpE9UqDPid0rHdLz2vnGrZbV/Xs9egPZD0ye5ZoB88R+4Ac353946Gu6Oo7qjRIKbTD9N
O3pnLCmcLZMUpLiizo1kmoyTfYudw/ePsn7f+gg23O/ZYzUS0OiYCKvEnhiFWJM8JywDZavOE/Pu
8QGtL3a8qdNe+ScGYk0brmlVZljKNLtIbRcJpIy6U5diCH6I5cLVH2nJwffdNn5GR5MM2tpJxyYK
9aVJlbnyd5Q/EiL2hEbFE4NSlqHD8bVUHzdm29yLNtYGNbo9qfetSHYd9Mh2rNfsc59Fi2L/Zswn
7IXNgS7nImzmWhb7PXh2lebdjKiFcZe9h0OlZwW6Cgn3NxUqkkVGKUr4lyc6gq7SItMH6kVnQS5W
EqdfaBaNk5i6JS5L06bSSMl9tuLOtVGQ6JI+gM4pc8ZlfscYOcOA8ll79F0cJCDcePoSKaelb7Uz
+xD0/DcObFuyW4lmOIBhSgwVe3BGlnnjt1uDFbQP9ssB/g9qgKXrkNqGWzHiAim+P2bB1GdSsbA8
w0C8WPQmjy7WLJ0eufE0LaFgjlWRdvtMciEv/9UQbLpY8P4ILgeiw4wym77voDAm0y4BPE46qOjA
XJae20xgCtts8NFRSF/NPgXZ90aqdu+IiuorgTIkg1XulX7FfXVCzstB37TnI1DJ79NTE+s6m1k6
sp1QmW/09fqSTpQMVcyX5h5oKOl7kRGR0hSIVIzTv7ykmWozD6TMdDlHjphf6xqovQoqY77w4/N6
B7jsSIbq4PKkrWRgREw36cjbB0Ok69V6fk9/3XzQ5iQbbZh+WHQmCWJdero8qy268a6YF0oDylTJ
WkXmz4UBEQesWjlbFjyTSLbGafXdvxXzLwPvfjUcKYUWw6X8jELqESP9KzsNpicujN132SvOFvOe
047Exls8AIgRjHl+xsxWn0QOvj7sIidAGFuDckT9TGoqhg+K4yHTsI77mBLTSg2EayVcxT8Auwdy
Hb+xMrNfzJyskf1MTVy3Oe/Urogq44AYKQtsQCFuIRC65ag9JmJFUHDzUi/JYit5DKPIUFPw8bJr
5jG1cgGmWBm50xOS7XoZ/xNi9FJUT/zmOTUZai76Mg+dvyP8WbKGiGj6JGMwcDGXIPNUM8f40cqG
dXoe6TFRAJ/ey2OsrXO/93tYwWfs6n9mypGELcw25EEAx7Y9vjotitVHdhX2vJWjsKbmgLcyndDk
MeqtdayHNEVqqKZtw8CYv1r4GpR9fnVZ+avkw4f8vdc983us01AJOJXA9LqDcsELNXWdrwwb1LYR
J6Dwa36rFypHlfnc7V53Nujk5tu+La6iDojaYuLDD2u9hEIW9NwH+HozEI/6YPgmmAgmvRu0d4oM
w56QO8HtvSCTPpos5Nar1xmbViD3QJKf7iIMFBGd9Pou0aCtLKX1y9PNqAb4YrsakDvC9f9qf4yD
j3rhc/WydJP+V39S/EOXgf4JGFdZwNYF2/kQwW9l+YCwvmJ2cPKqQ1El0FWbE/mTRI8WRRccYcqu
PncdfkQvQD4841/lkE4ibbh3mVW+M/7me5QEnC4OU6fQjTUxWwFeCB0vyvHeuYj2mt3gg2z/qfIz
1Mz2++TJsrEXI11E+64PsjavAs2CSww0WqZPubMni/cap0zOE5kd3yhGusBnaKsLM4YSlj3sjS2+
oCbvW4K9/ZzIC0gBdtqhnS3Rcdq+I1CFKbaWt8LucJMY/HyWaPKyvG94Y6BtOZ5fF/u1BR4fN8rc
Ac91F4uEFjvBEM9rg1lPzpv4yg9cMBDMcAw8NsxRVJWMbtSAnpVa+0sGTHNEavGd9qaAoh5yHkob
BCfDFhZ78OmWLQv/UuBnixjs3MgLNJqzLaxnQbA7eqMcacd8z+fEWOiVoQDaToX8ApSATYMTxu1w
d4tGZWONI+R9NqeK8wFIEwfMmsJonBPeNYC6SDhiIOn6BzbC/274tLaB0gXdHzTm+UvoeS7G440p
/5+RDtR04y64xXF/9RQGjhDDHoJ+o52gblQP6UJqTapm2xINh2uE+GNV4DhiUXLdeI37pyqZgrt/
a0GofOeSAcaj5KhY6QlswzXeAOLxKCVvTr/MmL3zujkg/NVEhXTqKg8paSiJhsD5e6rP3dVp1mcG
ewYNMEQfKSjqYvg1+MxDWHKEGdYdCA3Za1/Mslai7payuEEpBxW61w/wM/ptnY6VcGy6/ylLCPCy
WoUNCdLnyGAUiTQjeiJcd1jbmcCY5S4kuo7OdYkcrvwymNaUfXAgieBWDZrpfKWGBJt2ZXgb1OQm
mSXmKl3pXWXUqEdFDF2Nfh1/Qd0pHUAlYuBukuei6abjgZna8HYZLrwmMm0QukMCcaHLxFRi7+bU
z7126RFDZwIkiIuS9hEPU1pk3OM5iI+spp+ki8nSm0CULMyFwrxVS05GfWoOGfrelv0bVE5nXIhh
Qbi6tpdDUqzenABS2yq8pMhHixlFgWB2Jtu0Lge03bHGPBtn/9QVg/RuPp363bvvahpgnYGa+U4l
8KrCOiX4BTIilS3gpShXjv9bAzEDkK554EcGA9N66e6QvqwL7wDJEeCCsWNgtfP4A7xNWfBEJY7d
Ssu3U/a9DcTc0xN6DRvv8g7ru22iXq6YBdKuYezygB8l6EbeofAif9NQ+HuzqjPh8NmlO1/2j0zS
zVhMDFO8f1F4vJ0gnyBBfRR0CFOezY19EHKlQt1CVXyG0y606ZQDIM7DvFiWlFteIvcggyqom/J4
lAm5EYgq4/b2NanY7wym53Jv+nr2T/jyCitL+5pxIrBUCnOdovInyUe4ZdrkAyIylVN/hJA0ZMjE
IXRkZo9ze6HwI0ApDfrZ42WyA+yipRtf0UrMa8REwWowCRuhGgPWpFCmgd88h97WDe98itPhdp+I
8k+Nx+wCC/SQuMlX4Z9EC5kiuheK0GFC7Swllfy/WJ7oC4VR6gNfMDtKRzojusSIZhL2Ee89xqy1
8+4rQeXeRok5Mgtbba/BS60jLyzlQzA0laoipv0J/gMUnBuCh/ST+qjaQNW4dayqF3i5uUEIeAkd
DphTjcusyyDvwgi7Yiw2VCSNrejyps0fOKHQdbxG/VU6fONDUF2hO3Bd7iZ3G76FB6fkO4+fCH3u
CiNbJJOAOEsSijQQSctBGrSrBxmwGzGqEyFXpv2ac2Gm8BiJ4vwERPK7r6zY+BeObsQZkayhHuDW
B0wV+GDsxrmhxWGg5b3YZhTpyN6sQsxORpSI2HcnzfDjgpAM4vqNyWtuD93u96SMJwcM07gjGayW
iIzKw635U0/gkHG7zL1rj1woI/Yd1O5P3QBxi9C8/8/OrPGTDzwrSsCK2CnFMSeHPprVJFEbLJQr
OSohZmlroSX53mDe5OiFVGVBrFEVjJ4/RuaRPKKGlTd5h3rw8UfzRFBIf/Du8JvWg/yPFsUe51I/
9aap7A1zAbdNQlIkc8r3XN5rtNeZLULUiFD6qe04/sMHTC+wiXE19f2b4up9nsvjhM5oSj92L7++
ZR7to1yR/yt809sg82xt8/xcxjmmEaJvmN1Erepa0JOItiiecJXYxjT4DckVrXtlu8jIX4pHjfJ5
dtQQ5uYKgaNG8tMFqhOJa2YXxoIJZB5xGzcjvjRMtDkvLYOc82jn66W0iTHN0a1ezEEEV/BqFh1q
TRg1Ar8/PUGnHvdFT4H/QWmzlxpBuupXCz8JkI3bvU6X6TdftJHyr3HcUc5R/qx3hzHelwZBY8l7
4FlsjdoOIKpYQMT+vmPUaphSzds+nf7XKZ6r+q2X4oUJqlL9+oo2Qwl4L48Si9b28G2Wmm5giJPh
Nnn+C72WK1bA48wSkELyTcoOQQKZp3dNOlDFpMj96cjNDm1J9qSXe4rd8K9Jf0dW78Dub0G37mXo
8qISZ4NVfpyT8Xl9JCps1vBQwrJ4zS8YF8Kgse3EnJd/D2vw+4VZswDookohChTOssDe4RIJTgbt
p9sqq1TtDp7fgL8CZKvnfaBvek4on5E+F8eyoCTlokG3cVHp24eEiIlK8XQJ50cNXwI2vcnmc2X9
YtrPrlBUitEP5XZ0GS07OHNSoSJdpo7yj7XOZXjdU3bvbX3lrCRAr9lDgv3UQSSeGGX+pPfNeiaA
/kA03+tA8AL3VLthLo8UxuthI1Lr2y1V6PNth6y59uDaHGYN7XeIvVbmQjmxpgRDDMven5sYepto
IQDdTuT3FyTG3oID0wo2hPELcSBkbHnXjfV0rTlMaLhZpsV3MM0KNIHVv2dok6Q8kRLJImBhwlBn
4VWBawBat7ZldeihZ52KYNaHZn9VEmN1RhVFrVflUmJXGqQskKANpQbMRcotLRrdZjIpd7uU7VpE
JaSL6yvWOha7tpXEftByJjx1EXxrAARjuPShGY9axSWgPJVNZW0n4pO5NXHNJ1fCP+5rxcutRm8+
y+73lfLe8jIA5t0U21MstxNPb5hNqDELGzJfjGvUKhYYBKVvIEVS64BJizmuKSEx3oS5GO4RcuZQ
tZVVTS1cpFVrB3/thvIjuDST76Ly34LpiucDztMCzKO5MhhsaQD4vhh7JhPAYvhZoA0r4YXlqh7K
Lfl2Vs0tgppfzywKVlo7V2rbBBleawOgQcu0qNa9BdktGGMKKKDoZqhMo0PycXLoUU63I9u6SH4A
YdcOXqU3NZZ1QCcr9oLjNTk2ZCL25NiVL0GPyPNEujQrnuqDvCQ5DYCeppZhPYaC24J+olP5oz7Q
ObNGzn3oXSwT3XLXXPtpSPRuazTscGnLRFbLkB8lUSCoRC6gXWV8otlkM+iDuFQvnynEZMWLjYfr
GbYRSduOOOz/yopGXSePOR+nKxA+aHppenDHS2qigwJfs+DubPkV5ZbUooWw/pyd/mMD0bY3V5DE
XbSP9gQZxEYAot6sMVPwGf0JVFdQ7w11LQ0vbwdmz/5BObLwMNcd9T8Ct7RCSzozm/ygbZ8fLOHX
9znvrWAOjv1i5K0J6TqZJyuEDCIxIR8quIapDdbs2d7zekR5FMSFQ2TYBzdy6/KpHHmIz6g7GqDv
TdGkvEtAYnktBuax+28MxoPOwYBIye4ahIea5VbzPH+UNnukRBxY63cZXHLYTEZ1pnddwM7Y1B+F
Pnw1ANSRCVa4yGX6g84AEidZLzsgH9ZMnjhY5wRWvRT95WRPTZ+xuX1x/Y4aJBjyL8sxtNDQv9m2
Kz9gChqt3Y/7JVeEpiXK/yCxrqwImdkSei0SqLx70goQcuwSCRxdDRqbYjmIAAZCgt/RFoCetIe7
pfireruMAFkoKrSSpQz2dSnXf/mi/5IBNOQK2dgRAj44YxrGsdsuc8Tar4hhb6nycGVwYkzwrXSi
pQL6zcmIbz8mW6WsFmuXzLDuoZiLpAwOuc5UzoPCoduSl9YuD44xCVpHBIohPV7P5wvm4yN6QMEG
ms9Vh463Ol9EjsNYsL4hPy+cZmO2UJroi/+2/ASo/E11HQW9NVkuvrN8M8Ku0sTYCOn6UPmJ5s2/
xXqYtn5MyQ8TBVN8AcfIozXEsyjG2FVpiujHYp1i0RfB3nOyqEzZdIqL+CVyTuKAe/GYJYULM+5f
PDPhPSq7+NxAEA1jEyHMSEgSAVsVP9wNdP21/l510MCetzHWtYrdywjT0HTUN3N+J20XggUS1vpm
L1kQB2plZsA7IisyMTZr3NcS2iQUTUv82jYJbZz7Ef3pmePAHz43rpVKK3Wcm7T4Kwk6Okcwn5c7
Ky9bgc/p5fnTDU0tCdLIURXvzJLdD+MCY1gjihs6py99ntmm+4QtD2xET9XyM0sXv5JB8Ggnkg+g
EeK0/sLZthXeN4pXZC9wqxbIyhbqxoWBOnvgcdLe8UOf7zn4FaHUlZnCh79qSOJxQJgyRaSt2Jl5
DEGREG8xLb4Cq7FRvBL08ZGwo7gKfR/a6ttLKdIR+BC1qoYFZ5J4HgiU2Cy1TcoMQrZ7QcFRROU/
dcZAoPG9O9huvSXjRqF2MxwvUKLvCCJ+3SlOXSKL9jhiEfqGKf2Cwrnv8L7KHSFl4Mue3TWkgpr/
L9AHZb383pOirL1iJHr4iq49vReVcC+Bjz2vA68Y7ZnEpwJU2ZAw8cn8Wt8hGYsfIeQoncG/9BVa
nXz6+CDJY/Mu8JkiDnbh6f8GEbL12j9psEWJ5EmUOIPqegu1IopYSx55sgyvzfrh1ApiXkKQq10w
/6lJ44lFs/wV+rQYYRIbNwQVPP5HHBiAom71HINvAroSd/AH0/1q7eu7vHPy7odu0R1DfufXCdaz
rTZCaK4ny6sn/Ch+T/apQHd3Xw/XO8nU0Jm7058JZKtWjH4DTQ+D7QdVRQQnYQmm9UvFDndvs45D
lZcIpOGcMCKU7RSlgDXCN4YcP/Kc9nvUiu1slgNzhzHjEClu7rrAabNdsijYu57GCWSKdWVwFNBL
/0nAgaihpMeuED5bHrdQJR0O2jopfCNCopsL5vwM8KHWLZxmEo3IP0otnV7GtYn1tpzbYau5GzCu
oU7q73s9/JhG+skslh4v1LcHHuzLxo9EQ7BJppFlgfzStgDqbimhN9HZJOjrvemAPtzKelWmvdUi
WV7aFLDmA6r1l9JFht9PeMaAebNV92piBR7xKDaaYnGSCAVx97dwOy0Rt8KQdW2zWYYwAuNoENTT
FHL8HTXcIu7focslVff3xeQTypLw52QiDFD4rokqCAz5MkI8LBv2s8d2tLD/uGBXxHG/dWFipnpv
V0TVIdIpaWA7cU8To3ZYgxw1mhNGdSu3dqgP9iFmlxosIhcKrkAJDJi8Zbir7Eg6X17FzZUH/t1q
QhoNT8Uyr/9hXREVEXtAlpguCefrrnpoAwVdkfVr2gpIRgC6pGO2gr3j2f/Gu8IRO6o8ouW2VMeM
cbuvwJ1Jyf8pfGRLo/ryLcgNN1dexCb0lRD6RXAm9d7lsmpRa0TuVFsyaiPnyWxClsCP0qCDcFxm
GWyDVuuB/0CerHbTmeSlc2g29VMTO3be3qYHMJp/z3+wYO/5ZYxELPUT35blyTaOZn8ijBN3wjJu
oJybeaJsOlKKUchcyT8YsefQiO9BOhAg8olDYAhy/Ajx+tkNXBjLGkuInhmrsstPc+Xu9vSDY2bW
WKt2bxaxKU9wfXCtlGQdLhwyDGrYKCfP/3sRV4ociywwuulCLzfa6pLSTUazTc2699eABPtuEG+P
xg25WsGZ6yI41BMQ0GqNup+8dscRtFfiND/bn9H1i+vFuDz6ZkM4s45UZcu6Q+leZ44fS6JEZGQg
zfRW7d91PA/0EReK1yJAskaD4NFkahdStKqsc9pn918y7FgZm82+purqbUOmnPdsgliY0fomHgKW
JlW6+sf7vUhpv5hlsxwmtdEO8sQ7YlCNctnqebzb6zL2VWvTsnnc+d3nIwyL0zDVzI5DhxoxuKm0
Q9nOXa2GIaodO8CrUtNMMH8TAtDRquPJekIGmQd6EOHcDq8CJabQ/R/WXhxGkb+sU4MHroxfm0h7
jBJZP8coDwqaH2LsxF6Wq3jv1oee+g1soCJgGzQdiBResP9ynHym5unSgpLiFF+c0kMMD3X7DVbL
F3CZVyZ65Ihg8U1X2mjQ0wEW+G5CcdoG1R0PgdXW5iaO0QRCStOEdJgZYP2tVZtLMzFtLmP7SAl/
WWpi18VgTAcUWMjtFs3Of64IXhisbfksYM32BZ7uYrUpZxdSQ39eC1xiP9sFZgi0bwV6MQNY2CSu
TYTDJZqZlZIP+Yj9JpMkllSit6wcxwitUgCIQK967Kcd98K380Z5fCAd5gu+56EBY9ITggebuU0h
Qk6xc0Wx0BtQuNZLn+5sqeHQNX8yKB3bhEJZ4QD3k6qQc5g15oRc+LikmEgNevlx1IwLIJxuKxcM
cw+4co1vY0vnY6wok0T0G2zgETANyBdDbSD1GxGX6fIrBbNtmpD6xOWvzB6B+krWbI3hVi4Lenjw
O2oSL6bohP434FGzWXOWu6MG6O5qQwBJ6PeuPRsxBUBWgEDA/XZ69I7Ak8T2KBJaRAYAcjpPbbW4
F47jjwHAsO8bGo79Hn38A81Fn0fb8yTSETTFNgL2mzT4RI4272860iYC/2hO935cfySc9wdhN8q7
etmoIPPY+zsCDDAkN++oAeYxPR9HEgsEbBDNtW8lonaX8Np9g7h1N4wfsFA8NRUBjFb98kpRn/dD
B9JlkEKuPRmrldK6f775ce777m/K+8MNwSb+U8SEUfuXocYZ1R7qI9KVLCvFU1Ka+si7UCvGth5q
YgoM3gU246J2SKPjrSR0OYTtmUA+ripsZxd5hORdlraMv03gGCAFIkzJ9Q0m4gmUIexfDDAWYHt3
WAYm+qKtWhTdO26q6qghxptZE1UNnkIGH/T+ExOv6IUN7mVAOoQ+0iG0lF5JEF+21G2BNZ8iIGpu
7UrXPAU/dY6vBgdMJlW0krJrtddlPnlemhobGfAH4jYmKr1Rj3bVfyuVMVlpDsPpsbfun6/UsNdD
TDfB39sPNigK1fIrH2YEncUPycdiWpfzu75sQYDV90rwNn+1NrpnvA5DCiiYoryBdH1SwL8F/ZbY
Z23KXzZxqJHmkol57fI59AAOMxeQfiwQI9oNUoCvWMB9Y9pgKkZwy0xKsssXh4ypEv35jlPMhpV+
L6HcaATSiTFso5jv6nK9X7AkURS9hpzXJgjb1XW1VjE0FrhvuIeoSOlYat0ar46k/gYmHwQVBNPB
6JU+fYe7cwvJ40ME/+Hfnb1DpaVDOb2VVEB1ivgtfv/wpvDMhPFWGHgtGttLWOHXZ9OYzQWdMx4a
RsGuPfDLZ60eypMKFHFxiSqZp0rfI1/nBjvBkLPezaRCQUdB6fCt7Wv2WKFNtyY3YcLvamQq54vg
saZd0t+9a2Ax5qEH846LKAi0kKjV1eUuHP6ZFgB+T7bqjKQfD+b0bGxj6XC+9xkJekQ3m59lJcAf
eHRR6om3Gz3Qo+OqWnKJZiuMKRDbTBSPahWUZ9yZVv0AfEoTG4I1Ix1Z0jNw1imEsAbmvo6VISHa
owFH0BG93bfCgbmsEv/hJL2SjnL/rXmqHVf0NbT5R3bvA51dsf3gZyDs7Z+sZn4WzyBgdyUWQvM/
hPuMOITNes8GsvTc6ZWutMGMNie8xJ9vYoYTmPgyo1JuxEIw83wk1AUBSjjOexHF8lc6zi5NWlm7
oFaj+XHhjdMrCeUhO2ciFwN1hUqXYDJnd6JpX96PlAo9QhxL8fIXpeA8ONFivrFKF1XhI3O3awp9
yucM5tWF+HbVv3tR32yELoVHwzihNsmOIvVnGedI7VVgr14c8yw0rhHITOPiq8nZreSYj0L3G3iK
QIBr1b5OFHpCEuKdS6AMy8lNoNia7tvyUHHdIohPWPWYdOYVH89sq0eHv6LJvlyuNpYRzNWFXieD
JMgb/i5IjflUHzCojFYyTJWRijhsIXWATHffwcAeG9QQinLI7E5TvHwknBUtU+hiuecEG3QnvPiW
bM6l80G7Q1OF+su0EPqHKf95k8LNhssFJ2Ed2+45M/9Q1+Ov8Id8Tgd1DJJ2DR0DAaKPzdkM7k3H
u5OM8vqCsmKdbM6fBoOjKcBLwaqL13u0E9U3avTjP68qqeYZJCSmvbUlWbP8Z6an0CqfEhA0Aab0
DlT2cnY1VxnMpOsfH/Y31XZSLelcOl6z9PP8p+voaCA48birFgv8pXBRv91F10qkS8cN3gOrdMy5
/KweoMwb/fBMNUfb0n1/XAmBA30iF5EPUhnosHk4SPMiSlVo+lzYU+9tjHnPozbsXcb8T9tXXVVG
xWzKqdaIM2NJbZMGqLEesfvDRHG7/YBMBE5VcqaRSHAn8/8mRJImmUG5IalSJCZukPmAcqsDHZXI
0xzoEV/9rxUqqhdbTV2QaNE9YCmFP7n5+PCJ7QmF+bIql41AcYxCF8KoZ/JMO8RqOww4ktuwGTAI
pighejBEGIm6Hx5bj6Ss77XS0G/poH/E1y38Ml8V5mAXqXt7aRVwCvUDvP0CEkfCuwCNlGPZjTCh
xkJwOWEJKqwJO7CjvpPLsUUSPqtNtWcCQHob98YdbfnUi5dhipRvU+Ljb6QoKuTSwYjEnUVdldru
8+s3CfnlYbcRgbP868lr/FYpYGYymfRr4TfKEjkUqccAjZ77Ft9ZUv+lISvWMUdWlf4wUy4HuDga
TEpASx3WaeRSBE/Bo4YpOHYsnI59YzZs1Ye3rjKEp6TI8CwJjgbxCrcua2pmcOBx0B+SQv55mO+H
3IdabVvvVRRsm4TprNLyHUG3GSJGBDqlJMxQWS+qKg04iMvQNjsWVJMZOcf/XJWHjK+JEMoZM4Hw
/XEXgyeaaKrq7dD6qeYts+u4dQWplAE51SIum7GpEAn8kNns29Hy109rnrSPPRf8bBoI4ogWH9p/
iud+337LuSmN0eOmj7DOSCXXrFMhpQt69sRdHf7VMj4GogmVn0XYTGuF8pm9IsCqk9llErP6B7i0
g/iRwcSFhzNaYX9v0z0zriQHDJ/RHJQiq0ERRHJUaVRpjEFGFZKLLZq/VKyOPtJJGpQxzDBau1qu
8tWasgzzRSAp2dmddqA0njJGHYX/CdzJ0Da4tSFp32qlhaZ7fSjVIPSQxhn0CXCPryxxv8N5yN1z
rsJq6EbV1jDVK7amezlRzxRrA3m057sWj4kl9+y5rrNRPgsFvUdBaR96bbH4XH4cCW/OjdgKPwPI
iOJQHbkqXsM1LPC6K61kS6WEJdWxEuc7vYWsiinzlIO/7RDoTrNTEPXxJKdxsmTTbPGST5c4O8UV
LST1O2eY1LqOguycZMgi85myO+zNcCJx8egQRpU7jbFxgI2icqdqJtabg/o8MXzTg05FYezRaLQZ
n382P3aNG11LElrLuyO/g92mdHGQuYs0L/J1SD+qwpqCv0pmi3zKFPChDdDZluxZlAejjjxIwf5A
5ZqZD84smECVmtpv5YhGcGlQhoCOgkP4uO/WgLHMARwTC7gJZj7N23ljumY5/WmohLsyICbOcYNQ
7+oWY9Xj1iBHO16HIE20Rv6Wt9+Lo+FglONbOtIT/GIR1gF4gu9W5ObkTYV57ysedCq6anFxXR/H
ttRIiu/6iPhxe592TqR+GV7SJy3GxqFBcxhKWtjBzZ5NZW0MbXSfVR/ZsBknVTe+jGSZwKbsbpzq
H2JEb0dt++5Su9Ec8StLPPmmeaRdhU3Y91ac0Lt9TIVM3tOIuCgKR1p7YUQMgug4S090yu6k4Bp8
KW6PHp+IWIuo53fUOTQK6Ey7F6Tq4Yvv2WVJo1uj9Xo4Wl7qH+HpxBPdbMjBavCBrHRtFfgaFNw4
7TYQqXilcHAj9WWko8gdcdiGe5ma9djISf2cjKvVhDcWyP2Oj+IgiB99kYM5rLBh1brVW000aKgj
pUGgTIU2pwDGOjBi9FjXyfv+HRkIMc/BMMRhjH5N67PFAOqSAyDKJSsAR0Mtez7Pj+BJmYakOvgF
Kf5jP1lbyltb9JW4fGy6TzNP2LS4lbMa6NUwp4XBXlCtwkJ7NTfXO0UUktaWVNLS5wSpIv4vwGeb
r48bEdQXZ2hGIx6q1EKE0nZ7Od0K+w8JpI3fjP1E/595JsYLnjOq7tr7vH/sJZ8H5H6CVIqGDRcb
1DNbVDOipu1duP4xhP/Cy4LRq4aAQSwLZOuSfjrKLqGzsbD93lxAppt2/62UQtzWEELuuLcRbm0r
LOodhfgWWKVtPyuYBRRTUnBvbI41XlnNqNGV+nPIUUEbn2kPGpMXZ+YKYyDHhnXzGojRYgyziFw4
xiKOoisCA6ojPWk+nuwNbSEVpg9gMnEayIl09XGM3sAmTRgcI9gVbvt1JbLx5oRnTBrgEDtbIKEH
afWzykrFCuVfJDiVYW1R1zmZavyR88ByLh417rna3uw67Ph96NkVkkq8BKLPVjwuXuNiKRruktBE
Re1shqqFTbaeNNqh//pI/xDHCLk5SjwboRUnqEqQl+Hc+RNQMaLsYo5yxXqtB/MIrRMREPg0e/Jv
UJqvjVhmTtO38vTUJOpgdhvjhGraNNGL80f5GQRSzCjdmLP7LjYd63EWIBChZ+7I8gGQAHmLSIe0
5om7iR0Rj3xSX7Rp8P7t49JLQGBRjA8gQjW8hQWLf/R+8FMjUf1iX8UU0M6jxeqMuBc3JMvL7nce
Q2fFzcD/sEb1kQjRDRpLBnvwTaIwKRlEYn786wEe6MHh8bj7RSRlSyUf0hayx8wQZhXtJlT6QH8R
SwTINyzExm+JR+G4Fvcaohem/kC4NievFHIdFt96KgusxgYXAWTL7eiKOtpNHlMa391yNz8Sn4AS
6vpmEnD7ZO/Mb/KAHjoi2OTzzRHrM9arWaMaYjCq+WNAZXKvDXIlLo3AsQemD8u7O9bQrDRwFsSg
mDBWG7QL8JYlLUlT/1Pm/w2fbGhpfmhHPyk2RXKv4DMDHpF7fT7wPWz9ir1Bc6bHbmOIV+f9U2k8
r42DCfeZD9DVrHENm/UXbBCzh6pn9+Cw+AHIctzjALkkz4YaL3+ae32hA0N8HFF7FwIkilWlD+l/
J05Q+OLlnwZpELhp1ZBMle2vfZvidqIO08p9ZWVeBtK/ifegJL/ntVQ6mlqhVclG2D0lQY1vX5kk
vz0Hsy3qKGEGWpG/1kDz5ycHBtNGK8LWsNHdRJBsykAeyTUhvzWViG+14M9lVzoQU3I3p/XwU2cb
/NanXHXcWDRUSG9XtybSE6PQyPQ50fqo35G0usFXGnXUoR3AIdsMRW5Pj4Ucga0II1rgtUQQ+HpX
9fdunliTPRvmogUUAPhCRoKMy+TlvjpZPqU//c0l4vAzE9mDEgSIXhD40jchtgLiTimWlMGzQvcy
U3EV9marnytW5jpyzgpEfWI14Ynu6tKFmOvMDulCaTmko5suVAbL3XooAL/LQ9Z+IfK7bhqFTNZ8
vKeGNgoqNuimy+RMECyhfllDSWT+/Bz2k13o5mKNtGwHaubQt9j0cvbxDzN4eq1j7iPnR9hhW1Lv
ajz636WCuaV+wCKl467wbhCDZDiEWQVyjyI0sTZV3ahlC8DUABNzsQL0uDgrQEASNTtRgbmmJprj
l93rI9v9YRC1cwR/wCyqunqT3jxhIMLCunMMi6BWHCM+AnDPkYrsCmAvpQAS5oA/cTdKOZYA5OxG
8K67rhvTwedZYf86C0bDdDox89VBvdYgZ2O/GKxagl0yORPzDcc1R0n6UZ+AgPGjxH5HYoFSS+s6
Kehob/ziHcUge1pbGJtVB5TnkDBdtjrD69NwKG2M9f+wWPpIOwqtafgw0pwDS7rtW5lQ7Xx9LFgw
tRGgEBLemYL0/CRbFfywDio0WnsxZaiM81T6T2Cs0+o90l7bGlBUmu2EkvAcJLjTi8QGpyI++efE
VM9ePXXaJ3gJNpQdaMN16ghzuOUElWm2A4zm/H1uDW7Zi/Qe2JV5Vmg33Gltvo3c2GTPaeRXCBrV
PjQPbz7AAuMqMmBQMji/VSCdB5sHhPyN6V4r9OrBVDDCJk3KOpL66DNqBIr78ccwW7UXJvtyBMAQ
vfmC/+8jIvJyyqzy/BVmsYauO+aCNm1gBNtdD7imbI4wkdpr852JUKahAIcdKRbF7u64fkRJGKwH
8LUPy53rFDNMHqNOIEFCewB+xAo7r50i3RmZjkVMtDk18IYwoaZCAOwMCAAet+umjXvitHPkVVLb
Tt5XDtae/SrbnYACFbJGRYw+IpmfB9EBlxospUzS+fm0MWQMJmGl3NtG+wl5packzA4cLvNRauRv
CUQIGcjhK5UbJYb7CG8ph7MpTm3dl15Yd5YLgXcuYlei5Dm9TnNob0han039HfklW/7qYtFS8GlA
RLq657E69UanjoLCuaZX4GY+4JBEMLKWFqQkHTeh/kYxDEpkNLxrJh6bHpS41R3uegsKtZ2DOabL
CgpuBi6oi0qesa6CFTHjp53zY8e8hePNcKYbDiBXbgPru4TNxQNEICA2NhntTFE/XIzBUTa5X5tW
4vliUvSarlios7t422/Fi0KVBLITw10m+ANHnF8WnIvMOH20ykrmAfx3LPyw0Xk1Mt1ymyEXSopi
i7a7fI1xuFELC0/KQ06h1LN3GlB742zQvL42T4RLb7Gvtfgci7qIPuFOqLNE58V3AzMp3y2fe+Ht
fTJPiqDJdXn56fIWg0AS1ifeTGvqdJYkruoV34DDLAynlAmx5WPuVr7/a3dHXJJ3SFW1iPL64W4q
zzpH6P81SZnTYRuMXhMNa55epcrwZ/+kIX1VqvS1SP3+/0As1L4cD5U4uqDhfABIKbo3y4BeKKkm
IEBDXUSPb5aeHUQvtQWa0TDbC4DO3RzshGE87m7pDzhiYDh6UnV11NdmBPEq5Ncz2kHRg48/5fcv
oIDqkNXUTCNc2kWeNu82Qa5dCSivVk98vGdyE0COyLpkjydSBS5Rlztk4bFntBQDJu3sJ5MxOz+U
fxqfyw6W0lvfz+6lfa1H669iXLfFuGB2aQVxPkx3zclP9/dXnXXtAcc3Z1vwgBUWmD+CbwY/XpjG
y/WPLHKJL4bkD/3kgUS0uOx9tSTnusRGQjV1wznejvRdcToKCfOwVJpWr6KvymMMqgtcM3ps267U
OHBOGjdJ1NnTJ6uITPZ5wWYPwRN35SMJU4AyKd4sP5MZQYWAKn52JFxoomtdXtXKPQ4DuDaIInWI
lA2NNhW0xxkgNuXfazqaBclB5bigtYbBBvWeH32HOZckNb4Hoe1w51G5iFG56dn8224QMNfIkrYF
UW197XXZblKNt6M31uBS68XJp8aufUhlNUyKry+qeaSlnMJswf1oZ00ks9Y6PbAHNpV1uS7QeFPi
Y9IaTr7uNEAbhHWP2s0+GFbki3cQkDj6MsAPVNhTdEnzVUwjtpRCQ0XsmpqXbxnAdxDU2mVX0wHn
zMJHuSopNRTiQ3ardDDc3ZrWayN9ixcUF1nVjMkwuKSQWwBhs8FUORavnb0t7YnP/+qmAFpZuKt5
YOIS4sAa/XM0VjUkI/eH8FP+ZhzhLHYIQ4qrdGfc/K0UJseZBeaJ7f6Y0RE2XTumk6pYw4DQvWgo
bLY4FJcUf1atOsHK2yDiu3j2Ru4fyupIovNajNnAD3Pq2xj0feNhPzkjlL52Pkf3n+4Job0SswTC
n+ambJHQzqmoSVBh6PmFrsJZaYxCWdpdehv3lnbWfyGXaMX8+XzMR80vRbZxt+kTqChnwRDc7v5O
58vf2YxRCh4Q6apeLPXwQA77Ul43yTF371cKl5DtAWoQMzV4oPK/CB4xDW6jzEUT8xGCStCM1Ypy
kzY253L2XXkGnCSdq9rQMSTWNQ/UtWgSW1htob+U8lZ1xhWnYTqOAVB+Gmnpu+Tu/mOrXM1/7B+k
rl4sdtJPBnNhsK132upcLRduJlA2YmvatuNqbpZo3XWe0M9hetOFf2CZNf13LhQBvsaWVektb9st
4lhFpGSNLWDaMWpxKKBL8Uxla2UWCjzGxlbGoe95JD3QYQTaTVlexXY2x3SaVCHAWRHQXbTaYAld
Ditj8k+eVdYV5GvNPuTXsQQZ8PmAiQstMexVwIJiyasrZ5xQZgIZ/fJgP2INW7cTTw79WE+xyOi5
1xNGzsqADOfgvPWWvFolSi3T05RKvQf8/Z6laXa4GNNhfkxsdnyW5CdC8M1GWVw95eU6VOQTAAse
ev7/djarOpJTDcRjDZ4IhWqZ7C/XEvjQmTVflfhOoqQMDfFbZ9Jj7I9RZrN0+9KO+K6WxDdz1dFy
8cdpRDc765M4f4ceFgBC6fEbAVtVzb/z+gmvdBjA8FolJbrp/Matk2/NuZOOqUfMEXl+rvlEHvgQ
WE6/7jbB4rLV+eGwJwtahrTmyjNK2Xi7Q3OZY8YuPKdSDMoxDPKCBUwR8lHDHwz4ONwZXm4RywdK
qHoktv80sDdpt9DLARV3UUXInA0cvgKK4Tv9+lN9f8MG8dNmetsgueOcl9wkpi0/3AdmNVeEjRFu
yUXNQX2nhnHjeWgILDFeMj/sOS9VlvtoZhjEYvZ2f9pXl8E2+L4o8WoLbdNbt4Avxs/Np/gRzlRT
+KFe5eavuh4ylho1oqgrDGk57nJbc0V4cj1csvAmVMZTxtI417+U5JCspCxNxlQHUINmR6ZOkcUo
C01R69705Jfi7ajas0L5Nmyg2OWkQA2UA1IJ+qGp97q3M0m2QfdWIBso/Zo+IxEPpR8GoDMfp3tw
Wg4h/PalUt3EvwRu429UB9MCKytTM2Ki6UwYyDjCgNwLHk649aej7BjemHNa2ZICKUR4Y4G9iyqm
S223aP44WVr2FEYutOkaQwUDtGx+0irFfhtbw9xW1lxqSqHhflszBNEN7wxTGtR4byyc08gV6q8v
E+4wleiq3jNEtL3MUWUv9xj1xBQ4VmZH+PEyFWNxnmalfP399xfu+qPoftY+DanjkuK2uXl1JzV0
ReGuZ6Ggn9nrdUH8XLxniW66DM64EWx+3DYmeMMRBL4KZaemSx3hCzIA7EuUldnvBdjHOZe16Ske
Zp3o15lvWWk83o27f9trdK0AekDSqqIanw4sagwKXQu6ZQ8hpqOtDLXtWiv/zQ2L0blZ2rNmfMbY
QQ515aeRt+RYj8kO1n26VgRzocPzx15v7B/mQ9fX8+nzU0fzF2o9VPvUkfAPraVKW7nkmldBqS5m
T9HGyaA94JzX8PfDm2Eh+xw8ubME+TMh8H+aX4eDUvWTmH9pZyJHkBRUZ37+4enUiZp/sL242B+q
3vXUyw2R/tfge9eIksK15+ytzSHo3ncrwBlpAyMW8oOLlMe4rt4cyyxhHEMXbpIV5AWr3SOwwso9
fksyMU6fDhWFvooA9Of2lZ+r+6vpXzWweAqeAkOk8dwNHB/bUOSf8D9ZtMDLeBip3BLAkEaOxt9c
L2pkNh+OR1j1s3f9CRjJUQAYeU6B9ifk+tRreIHwFEJPemJdoaSO+Fn36JRAKaQP8xsmgimr4QW3
zNroKoF16dRfVrLPMBmV2lSUMgHxlhgToSr0qPlNV2Z14g/bXPExDWAX8tZTVp1z2BVGmTa0J+VE
qwO2vBgcmxPrA5jnVXibT+N7vwfBq6+8jPC5ojPmY2A9B0Y3UO4Avq3f+t+NURriZgADO1EYH2+k
k9aTl2hFZlvL6XWb6UTIFQ7SwYqB32JK74n8++PW851HUL0LoGNnd9WIiHWOker4iBGcqsDGaoVy
dXJBecogflhhzKKxPLLmyRxz8esvpIylDIDuH8uW8zBdLj4IQjBL1FAF7JJl4hbolxLdzu2J7fPi
0aUjSkRqrgT5yc2cgK4noS0sb3EbLVIe6S4i/xNhoWIIICmXGO7uQVYqJmXiEOsUKwkLSp6RRuCJ
6f7gV1fMX4d5cQUYd0gooFqlpui6TTHAu+ncmMhehMf6AmRvZ6z6um2od/n5156GrBUHYJVV/J97
K7rTP0cVy4Kam3Vh9OW0RzGAJ8nOu+WIjwLgVWHyozLIs52tzgfTRuOl6k01kwVTWRt7Bl++Trmg
EEcYvDRb44iXQmZbARTTxEZhrptXq3Rg7FvYnSj7V92HUfyymEH4NuznbJy+3qzDYGdUwf9LIvAs
lZ9KDzR7jcbmjmPHk3JydFWL9JzdNe8NV8c11SOZyDq5K7HvrsnK0DBYT+2ZsECgdEJhQMYay2B4
d/zuncNAtZyUp5mvoGmvcPqPFq5GNKMB8L+SxlP7M3DFW6uWPznw7QyG9vVP/SB4DzFaWLSOUZFu
bXk3sACCJd9UKOPsdi31BU5wxXgXOae9M4SnmJXKcl3lV/vpamjl49V6SpJF0h7gOZaOsqcS+nnp
kC8WXrkY6fpRsvLb5IX8pUCdkDg4I6vnmwgPPL4yjyAc9Hq8CIlmTTI3F/2A1s1oeMBZNUE091MG
Z8mAK+woJw9HgS+qw6rhr5p39iy3GZB0dS2Kr3Qw4yjttYgqlnyKYtJwKKLMZ9535wbfls73J6NI
EdFuPxteuQXdaYR/ivSLrBhQ93VYL4XvQUQtFUqrQCV0g2V+CwAwoB34PV9+1Sz5nWr3tMXgbaO9
g2fSysE6/sw9ULOsV3tlfh5Hk00ZBwrnxUC6i/Sv9wd5wlq6Y6z8T5s78e8aIVKj2EI0qQZqdiO2
IWM2rxOQSrM2YpPGhcfaVFM3HRpROjZUW6Y2wuVf6KOQushXZgDa9Mj1M7c91ziusOTE6TM5Kvtw
/jUpZOshVNEe7sYcZCXQ4D7oFsdrJ/5Lh2KxUMdjk7VAgtFswlr2ae64ZXtQrNsHX6LHAL0wI6nw
//8eMm+WOrCUdo0JEVkplV9eHFdKz28jrp6mndJ0Qh6qhszzT5BbEEbHglp5yitDKTrujruqyeyM
u2VWL7h8I47HSOZjoVrbfskOGH/cokbM+P0gvQu706Sq1SQrLe1l12bT3EoHCerRyqh7+Jvi0QFT
GVrBjMUApWDpqlTwzPEe617wxb9ClaibiDhUHyYma62bnKNaxXmb3BNcD691AmXWr1KoF/t8z641
jf3+N6lXWJpG5iTQtP07idfDV/+DX4lJisSUgttZybUlV90KUkonvIGZbigB3JUc9jB9NGL2Ee3i
DpHGNzsqeNB3Pj4+KuIy0WjQk9g3Am5Qq72f0EYprAi7KK/VRZobfR7DWDmoKFfYF92sSJwqvrqB
k0ysOTtsdz9xFx8zckZ378rX9xvlXU+/Wspb6AWiE6NYIBLBf4mh/aXcX9Gx4AltWhFy9P/I9KNB
D4uI7n0yIWGhzKzZsT1MTA+zOlit8xlFdZ/kY7aGm9jCY/ldCYsnMm2028S/XE+rupHRjywQRZ3h
Lpa1ZUD0Ul+9NiwjBUxbySdMDl1jMdioRL5TDYlJ3A751fD8ZcZyzTaDrRD948vof+FCcVPuIuRn
qRqJn8La9EkWaCaLwK8OYybf6JAhtcDmVmvGeaFAR76e/11fj0FPau5iT34LM6QogbBygCvJw0pu
FcKXb+JyMBo5B2FQX0C5iXGLCrV1GDy9Fu/xwF1W46C+0KEA8QUuVcXKbv/6Mv0kLKktE33qmLQR
pTMkeTG2grnFhfiDgZS2v65i7QzVtaCu1jzITUHRoRIYpA0pyRrIbqvIiGrA5WUdR58psYeLB1MD
G7HfaU7+EYiuNoeyLIpGjHVwXdphSH1+uGRQTK86IhliFxZaX361xKZztvu244iSAKW/fskg0AJv
au4fydF/E995DYQocvQYr2AUWHLXP6+QNKQo1WiA500p1lavoE8o4dHxmhBL+0yXMSioTjcyRpX+
EI98VoGFXykl4hKFz30zOmkghobgx2XohJNAwrtYB8S5P9Kz2n7ZiunOGp4+bIpToIC+1CZ5IOts
AviRYWKquJHNtwtB0Imgrd7CcdWAviEGgsx74fIThPQZEZyv3vDXeASmDxsliXH1JCMemV5KzFas
VHjA+XTXA54/3a3WB0TNV9TfN4vQoLElaks57M1HmiziEFHJHp+wcgVxXFawnYwJXTLj5lcELzCO
kquRIN/uIAq3HjEoNRrZe+XoOU5yp6nusGcxOvJleRj2vSaln1sLgWh1+c9nGKZ1AEn4T4D2rHrW
WzW00l3U6WM6NOX86IdLztYwwXSfaPt2SB+6JP/M6S61WjBSF9BJxYP8bMDkQ29mzz5vJZOLS2D/
F819FRsHhJPxEiFptZ8C85HG/Par12Bvl2XEFoPEeAaSC7mC4spcVIVzxsIFw61A1/yAfYM+5gHJ
r0Ft3d3uvFdk/TsgvEP0a9ogdtPVf/tgR5VCidLwyr7bMygZGz3Qt5+VnLGcxHqqNnUdR4RJgyVY
qAVdZIUDFXcw+FFCwZtNOMdQ/itfxFT/CN6YCZ/RzTkwQTk/S00Gj9KHsyUfcM67wGAoWyzbq7IQ
LzUzczVtLxMRR9DnD2XmsKorwMJpxwpBQjOvPruNKYW8+Rc6AGyHnTBDw1QoIFwb6EZ9V0v9I9Dv
tiIeAQDkKlYqUOtJAAysVuv5VPAYp84okwU24cfZq5Z9MoUrcep3IVIaWqOlWCY7u9SMzYeZOHHG
maVPSakNqk/h7KioQ4hPmb+9r+qfwEfScTQpemA6gbjPVsQWrq9adCfGLmSVDMWzGJ/UyFdil2FE
gYYN2bkXQEU8uXhgIzUh5vlW1J+wMG7+lAHaqw6faErrPfSiR/s+ZOHrYTV2OWiK1kcLTOd7GKb+
6oMAVQLw3ulb9/sUCgmsFZDmvo9/SN0oEf6onZKtNOi+PuWNhy91GLXo7MbAoblm0/PEredA9FN8
wdiPyWUrgOk0WtpiUXJGn3cvMQRG/vlpyn+n+zXsH/vBhti92s0KfoHltP6DvZgPEhAIBbHo/n4R
EntpugeP/OJspvtZGjSLpVOOg0e6SznLNFlXAGfL59zj0sptJBXvfRAqSJnTN9Cp0LnZ8GwFdgJp
5yH1R5RNwQylAaYI0z1zKj8OKY8upC+C1SvTK7TT/zQ4QfqVk5n7yynLsa95A7ljWO7T40KwCdy/
qS/p/wCEHbarIiOKMp2cg1h63RJ25m3saYhIgYhtwG8xF5esYXwJZOYbS0vqH7FokxMpYMSrOAK4
GfWsTnKXkMdSjSpT8+vHq1CG6g4dEiHRwF0bWonRaEXmTZExNW3Mneqxuf4GVea2JfBMSPmjezpQ
UhoHPg3IgtpNzrO7LIzc+U84lD8boEwbkv3kHiunvjRI8xhWvXdc03SkmPPHRl4r6Apu3L/PrHZN
VUHQKF2wy9XMP1IVbxtpRmg2FBz+Hf1lz1KL11Poj2fuinUv8Bo/B8TanF9Z/eIywua+4vlXPYSb
n5DLw8ycv27qIJt27/iraTGvHGzjyqzE0tEkH2/3MYGEzybQzUraOK0KyHwP3uEHrU9JkuwvbcVs
aD2DvI0XLBNFYTW08FlAKJKqw7hPhPgjT8vavCSBTt625SFAlgZ/q2+ouTnfqt/nJFRj4XLmVMbj
GcBR969ZBgHaD4Au1rQtsa5hulfOsiEvvIuz4w7fGTM1e+oEMWtRZmiPWfLobaXDlKc8qzI79njA
KZElBIU2LVlZdg+6qGVZipj7IDUZjjbSuvnNGIlhhq+BgT9fYag4ZOfLxqXWN0c1fhn2hBH7FPJb
OwQEKEm37pD4IrkLTwV66DBuHf7LIiCjDL/lL2akgc+ATLAKtLkKlkX62oAnEAjAm0Ck/0K/LRdg
urMumCV/PLrLM2M6pIilA0Dp7ya02mSehRNaZ5WstnlsbkKpKXulWWBPelxtrnD4IZc6TTvfACZ9
j4tO6fAVa2uuskq/HOmA5ko53fUL4h95NH5UgnLiv5nTCgL9xkG3Z2VrdRCytOWRK9Gw80ym6J5O
oUsXlAQNm2ynrCE0fNB/ZEwQwp7+mcx/hponNlq3dErp65wdPRx9eX1r9xgDfAHTNGyz7inyAFKA
N3PvOEQq1RHIGwanfOoplLniZDdIYvkm7EYJf8Wrl2cuqvnlccXE0cYUJlhEsvV7QMZ+goEo6Xmc
yhVTFsqnueH6bbH+JLi0cbngOHICieMqu3o/4l9h8UpgMrKkQfBtXcJfvryUFNngwEhWCece0GVr
0trPniCPy5iQj9d0PaQLG9TfyAK/7AbfwKzKyrRKbMy1gs4LiygcuYdZKvTGvwhnWRz4luScNn2u
71tMRLHmmWJ2025jLFX5m7dDGElf5yT93Z5OgjApF9F9VmEyRF4gm64qYHkLgqj1mAPf3vaYhLHS
93gaS19ae7wlfkA+x/hq/Q72P8q+lJaLZmEMhR5hYi07C9fKylxZfMP7fJDylqrX7wzwkptPpVqn
WXSZER6lgpKFoBDAqHy6HZgOKj6RNiPhBvP8exgv+8MCq2JcsNGjZDjyIf9/qGSQR4TNnQ9/D4nj
s84p2FInd/v68pKD41O9KihD0m/2fChulJmUrB//WkLT+ornSpekH0jEIukxlor9GupQ7BsSEoOx
EzUpGEjtbsnCbKfXhUrVY3Yy9NoE3eOPYJXQsVcy4xWvRQ9XJ35rQnJTT+vVFBRNx3wZppY+V4IU
1fMNXmW6dmRLMMHKMjCgp8deTFv4+448RKKhApfUH2vcWGp1PJYGZiSYuiLNJ/tTOXyj9sRKe1dy
HxqQvktnvY8vo0Iw2LC/LzYntkJki3v9mPY1UPs/1By3Up91IZF2qnn3yjs2Oy8uL+vCL1aKmz6k
xuw/7CyITgw/Fws+bHCm4o7b08bNx9ZHVTocQBtATA1+JI7e83z5vLiziTZ/ddyZOaiqTaS5NDH9
4lj3KN/iFUrX4qhRZ8MghhXFoPvFSso8eQ7wsyH0fQVqxXGO6BmfiOAouHKbgswwsNxLchUat6bE
56UFEovkZnZk8Su4+nT8mb2KsreghGzyROHe/Cvu4kS+yf7vKVqtQPEqIyBz7z726kct1KcCZ/4w
rLUBXN7jd6ocyTrARBtH3LbbfIvcTUkiT2McBG+3x2XafkkcWg0M7Cgv4k8UnHXETojySTQaCfXG
+spvnfLHzsgf97TtwtJ7HHikE0rQBQvNx0HkROG98RMWWzmiAsMPpHX6QGc/VoRWfuZNc/xw7jhg
aBjGsNboHBcnsmcGw5D5EL6Ea0iSCeX6gBtA95lMHvZpzw2tL8m5lp+kUv/u0PQMsnVXKTEHZOG8
r3lwgBP7Dw7Y7Hl46GEzeYOFV+uSM80cGHatPZb21uuwNd7TIKirOJ4b4DAUpk010oiDBhzzXshg
DwzESlTriXV93OpKEY69cDOgimO8sxyVHPwrB1pvCJC/7iX7CvFhN5grQJz8Vjn3FLJ0ipKaQe6Q
CK5ETy9lB3UiUYGJ+u4EEZqBlq7i7Ssv/q3lVux2eZnCg6eV9KT9T0OC2qQYCB0VGNL/b2UVaNgc
QnBWTl+5uJdhUgBDXXQm9whOG2JUhsuzWcAyIpP/YQq6jK6Jb19uTOyS5o4LD+2lwdhLzA9wIox6
JP93uDaowDK6jysPxPo8bJ533F43XrNI9rvsKICdpfmRxULSiCnIq+AwQBhnonmbNEeE+1KZ1mep
VB/JQh8lrfbVTGw7v2JkkFEwpGVxA6+VU32qpQzfTZOkwBL/YPPTwKHHzXcvCKJgRaZoI99ioPgC
WST9SnA7UeY+aFh9NmWZ7SA2g2Ch1i9Ty4mvnBH+iGHZjGzMTAXGOEZrIK/z+6flXcYCvay0xP2D
/FfiHHQ9L/bCU4JpS6Q4DfZD/FpnOCmLpATel50Urpl3/LrguOLKHPbw5z7N5gFaxJzORF8Sy4u2
QyCqhk5OBsufFFU/uve+7q65+sr0sNvzK4Lgcu5Iak/kCBaIiCoSXI5kd5rRQRdSeOsrxmfuxsRe
qAhYljWnmeVFDKKDeEj+cHy8lY7uOl5Ofn+2usfBPEWmC7MqYlWrJjci9GoCKdqpuXRoEWp6a7fS
vZEhttapMjHeAbObLRMiDUtVRbFQX8BF94KZ/VaDMZbbPHS9uHZemFNVOw1KuxPxEoxucaArbXov
golZAgTx3b0cdzwxEQdgkot5Hp03TpmtZo37TDrNwtqV8QNfLtkQ+Zvtru1jaLP8/DChEoZVl8bu
1DMjp29PRuJSjajWhJtLf8sXgjNLCtYfjGkjJPUmefSbiKnls+IJWEpCjPuSCAT56rwVKqML6GNu
p+OegGcrSaFvPLPu+oSvd9DMR5w6IJcnKSb/mBu8RgXt2f+86/7EhYKGcq3+xTNfGTF8/awVYezg
aKmKNFE8JIkMrthtvSZ2kn9vpzTuI4ZZwVQGXJ8CRYnAP65qRPXP+KuvRl//hPgSDSIdGaapE1ly
iVq0Ib8u5WYpE36zkQnpIrrrf3p/0kAyLewj1943oVvIwsphJW9075iihNvSBVzbs0y8wJ9foTV7
Ml8JBUnB29tgAJ6VRucgWBku/c9h2CH00vQ6PihG2EtunOXvfhy8zNKcHWRgidG/UfijJ6bW83hW
m7Trn+HmaU2matueTCuaA5YAHMx5mdhqLm2BPVNFl1Hp37Bhf9+uy2yCwCyrWwA5bHUIUFY8t8Mv
S1r7iCdxf87ENU764mIUIQ3Qj5wfXd7m6HIQ+kvllNnnXbSn0iGR5ORUrn0SnipxvdOOjZR0KvCD
2CbMLADTiB1lmzapfZLNnnaoZd81XDrq5d1EtdWKh4tyyQMyNTm+5ZA/V9E32rytMWJpZ2cJ3t5W
tZgg7DsjayEs/7DrYRLbicNjf8N6GMjXAaSRHbD6YRjlg+R0eIB29sOyuaQ1qsC9syyh8PgH3B3+
+qUqvLzMtJfWhw1cjacoqAnofUhyboUkf+XqjcQfnH5vvCL8e5KMgBDVw3J27uuwZRVKQ+51B/6m
zxO1zSMVfzT1P0TjXFzpvzjiP8LZpO18ETJtSnV9VfzEr42mGLFMS/YiEucJ4Ho09ZBj4wIVq6sq
sG9umXtOr/4WGb8Rrj7o9Kqr4ecPxQHQeef77fAh9ODi6zVOL6OQnVoIO4EsKJTHC7cE0w/tVQME
SkZbIOmar3QkQuFPTrqP29S9h9EcvVU3YeRNVhDKQJOkgzezgm+rj+zCXYleMXDdd3hjn5A8Ls7W
73Bn3wbUlsuJl03Peg8mc7nLIelJZUvyu1GWjazL/7guNPVV0oCXIBFjodPiG9qty1uaYeKEPuf8
MdGePLnG4KW6g+8VvoPSd+aFZNWhtYJet32mHbwnFmtsbkfy8v+jZG8JL9+CQ23lgyw9DEHbo4ZC
+/c1JlpQjTFATKJx8E7f00Y54zpTRRNYtieWOw1rFzeoRVDY4v+xChxsGSGkvtKXqT1IQa4sqib4
86WdYQsXotGu4g7EvrvdHQKo9hUqsZ1PTY1XbLkaJ9S0V/IkmqC/9eK8iZEENyuMidtEz34nj+VH
YGDrrmA2Rr9Scg1rRxE7S3FDfDMyozXcDOZ+/uqLcqO0KOJtP8Jqaha1rjxD6DbWLhy0KTB/CwNW
PJZcqncPIObtiBw8tcvJFYtdWSbn34vn7/LlXgKi1GYYG4DXsScnQYcvjM4JY3n5fh0rqXueqAwN
rKJgcb1OKLau53rUrMMWJ3zkVvaumV1wRneHDk96natqB6IsOuYAuROATBdQbHyo9QOekRWf6CQ8
na2+MKCq5uSzo+YL+jgaI+aOUm2tvFtehpiZof0bqM9SX5n/+EwgWYV+H8z/kyDEOuSuEuEYOLaT
NsCser1W3cp5w9TJO/juPhdlX8klui4RROd7pRscXqGZIH9MQ7mO/OZilpywKz5ZqT3/qv4ZX+qM
WFX/FLtkflshPKmbLJEomwKJZT22UbSfqntreoHyLD9ofePIqcMo7i/rWsSCmRJNJmGrq4ktzykj
eycRGh2sKr0vRQ1lXE2CE2MscVw2kLzd8fsVIGSwL/pJh/thRBUo8n6gxrbii37XqMFimoV/jkaz
p/lYGtw0Y5BoW7kgu8OupmKcI+FINgHTl6qHn3pe/W0LxIXcjekmVMeS1HRwVWqmMY/2zn9qa4+K
7KXZE5doDZNrabIAg0/JcTkFp3yKHoPCQKkYnTL2a7B/ue7VaRlU70dg+DAnIkAwfTjWv9GftCeg
S79WnIYUlZtc4rMUdY4EqD3vi8ljacdL7gCbLUuBI40ul/wJKLr1t9ehogiXHcBs4aR8kAxFvjpe
PsA+lEuGompSUTSm/7nrFA+Yl2cmpKOyArFXF4pstta14W5LIn0ef1+gkH5bEcTuxp4902n3F5Zu
DLxPX6ySREBlGewEAm2MVDpO4q4j6DRvemIZu7SQeK9KLgcq87+m7xcPNgVMpddPqif2YH4PhohW
drSOfgC1iwfllUxyWvwWVJGw1AlYli1l/xPYJHzwB8B0Xz94hOV2Uwl/OdgX7vDudyToCOdb6LSZ
y6AS9zz7go4I92CmrGUaAPIZW89LsCDqiJ+72bEOAp6+JhOrXDe7fs0LJ0UYo3Pb5+dDwyyJG30o
ACZXveJLv4nor1qS7XIowJNjLV8yT39E+96GFJHKXazTfTA2ZjtO+0fy95zULlSpuCZjQ4bdX7d0
aXFbg1aTXsy277a3wKPr2FIagJRzUclvH7tOA891oqW2uuPcoGDHlwiodtb62ZPU+WJtpfIkBuBh
lmGoLUqIR15IYo2OzGRQTuZbUH9OFzpMWc2d1FUl5o4kwDJfUgKcR3IBKt1rZdYNbhXMxS8xASF5
veSawnqLCEDipDrR9H6/pJ303PlRxPfP6YOA4ZUR2Lk3sQu90LXNc568wqSivc+2D1wT0YoxnDZM
zvToVdX5iWWEOny5N5ja3oipNOfYkBlJI9iEopCVL7m2ILeBJ91PUrA77kMiP/JluDawRMel24cF
++eijRFDnnXtLgYxb4neS4sSy7dVI6wfSDlz1FzAB2RytNmtHU6yG/SN2y9SXo87WiPnul3BkXKS
uxuizUJbM7LuLspVB/9e5ssrttDEQ4Wf23imkq0u4GMD5A4dT1BiQfJZ/hjh5P3mrKkPmFtI7ElK
fYZQkEX6lQ+R5PlgQKxsOXaDK0kNI+fFSnt3W5DV0huFVinJOPpDs4XJLRY/22gGC56snK4qS67l
+hd3MlV1MLIOm2Gj0pGCyJ31l7IYlnwpGPQX8/GVzUgd1wi3ar/r7UwzHVsot10mJsoo0v1n2rB1
Z7Uf/izV5QBvnX1Le1kWM2FqS5XuJsfo+5XIsD5idccLAivnZ9XkVc6w/KnUXseqqSlfeMHFzSt/
7u348wGzAGRAKU6QpF6xmxsYHeg/weC0smhqEVWE9x1DkInCgclRTONzCBrLJDj90NptxHs7KQ0b
ZRYS/5Ie8kPUhoH+r+bM0bA0xPX2dc3pYLPj4ikOZpZVSR4PrUoksF+oZxKVBb55lfK6CdqTJjMP
MSNfl14GaV/Fb4Q6rmVzPQek2uxUSTNVt8s6T5LY6WwvgrU9AToxjGe1KR+ozsDh2pcB/aVma9t1
ziMDpdVKBOKNDRjtSRrBqqPxtc+FdLK8pAfnqp1xyISU5JzYF206HPXqJJvBfGP+EmKEYeT8R4ob
Of3fP8IxpS+r6Mx6BbfSBzLBxH1KJLf/VxdrJ/YH2beVlKdX8qFmsohqai2+Y47w2HjKKaXWlI/I
SJ5AhF9OIMw+KnMn/rdFZvNMUJZyhVlr6BKx5vMkiCwEC+KPZEmHC5DvHyrlFMLUBxDQW9b9PYG7
9q+e0P/DKhD9VO6MT3CZO40fteJgzPuQG4dlOJXzhXaKw8wrQeoZarv6oxDOn++lW+2+rhZoBZxF
medHTH0KtxVPk8p9QFEF/yT8ld2vdVr5JVo3lOMcZo6gAF5ZGu37MxvCOhw4l4u1lvMjPlohkSyO
thQ7gXYHwKFWENPDJj+LSDfR+ruXFVSYPjse2ehdcca3r1QhgAb0YMfe3U4wXw6oRIQV4jKxq+bd
CHkEyk/Hy9C71oVlEZJv4dv2vCzWrQ2V0vCkcxws+YAvaCPMuqwJguQqNakdUrv2AcYrm4pazsnk
mTGfTrywuAJJeuRW3oOuOOxN+zuhoq7+q+ELVWoxsG80Kmw0fI+iHhj56sO/ppnAuEexmkWtxjX0
4ZBAfM6v2i7Qwgy95aIjjByDnA3ezhTrxdsFcwcoAu2lELza042IN0w5c6uWNCbRG1Zn+S/JCa+t
RJSdkXzV67E4rYdukry+OAKOx2gspW5WqEU1f+qu6zBGpk9tXapF+fXIzytnfFKqTXANgVrtgfyD
SWvRg9FdzYtUJUvGU81nWyPVszvg1bZoPNzbYz76dIS3xKn5HK5mcOtcx3Guiy8xE/mbEJjtIItA
fUJaeD8MwaEkvOkPwA3Dl9IM9fjE/Cx0TiGxFE4kS3eX4bRZd67xIsvxo8W3PhaCKYH+gB7ims/E
tV5W5AxbrmENu2MUfnUyHV3kMqLvLk9tq3Fr9/O4gcmxToexDdDcfHh5iECnKaeu4bFCJ8OY+CFR
uRdWDW6Hs8R/KnOD+qOU1UFoK8rYoOWlrRURjKG484EkyZuHdD3E6Em2e32BebCN3WAt8l99HhPY
stWrZmCqdfKGff0XGkME1uKyyymyStdqjMwgF43esUPLl23j0pMfogVDsiFQELAVn9QkhXNPc3E2
YCYqOPBulqu/t4CtvM3i0IdnjAzh+u0exNJBVxrQbteBCjux0GWZTy4JKffNbanhbMSVJE1GRhMn
yNcBJrXApeC0I2PlQRx5+m/Qnz2f34XKTYcHds3kox/VMTLEQhbYOVgVZ/qtyjI564hImBdGRrqS
lvUk6KP3zYfSVNZLBLKuayt4HiY2pzcPPu8HeYD6HnfvWivY5SKoQa0U5y/z4+7/xDUvkAUzmjyN
ici7KUpSjhqrbRUMMLUWifoUrQq2nrij7k6Af7BDklrVGlN7ds1dt7AypzoUMaKOoCFf4qX+DT+I
rAgeYeFjdbIyb0JalTZ1aLEkayWolUw4pDHvp6lmhoXxo4+7Bl0S4c38In7X/foe24Ad5AXbzYF/
B6SApqv/Pp6kK/ipqdHu/TzXabCmO6fabtTIu6Fq8IeMfOCT8zMlY3V9jlRx2HHBZrXt16C2Y9si
t4UdNEbTLiPWhloiGXvJJC0QEzxbjSSiUaK09l4A1ekIl9pIUM8jmrsv5CjCjbIEiieyDzS6fU7j
SAdb3LkgU1LmraxFA3P9LrtNCH3Y9NzQkz6nNxcJLo3xenCAFEeuRe5RTR37h90jFrwHsEk/04n1
W2TZkgCtvA8pAXcjmX7HjZlVG3hn56bj3PB8YmnihzqYrKG6HszMT93OUGzyMN5VrcjPViWaBTIS
1h7SWtoHK/a5iPdqFfjInjeieYtokgQwYLIU5264Xi5CDYu1lEhLuXptZsyG1oerIYmfZnMQD+yj
E5VZKdUlwgcZSvqQNxYoUr/1UfOHwE79EQPpiIXVyd1gZ62WANcAgF+BbDbRycj+k7GqKCJgUb32
HDYKBuq9Zbwwk0B0qvCYgNpGog03taHjYX/CNOF3G9rZDImsCjjVZXdZVIZDi2A26r+eKnx4xY/J
T0gaPPjD09bcKdrR/Wa8Yb+B2Ly1ExhzxRaDEV2od8R+JWUTuC+2eamS1MtQGrE1q0P02RBcX40O
oph3k0nNRUPkRcyOicJ/BPdzlstch1JsVDrKEPTI48ZaFVC9xIuaDly0W09CRA++QsgYWZHoOXKd
DtPOGsBZbETsBm/FY2vyucZ5RSl3+6G+95qmcOlL9EMPMHeQ51QUiooNrQsGpn+InpO2wAesjdG9
r7nJWBtkL3udYtnXpzNiiUtYyUXRcRCcxHQjGF2KxkSUc6gd/eX4bBLE8aXRdE7ae7BHmiBASfTY
m3FN5FlKlghjRcIluGra3XZuXB8w1nVJEvNF1mTnF0SPqh//DJWpEFEQpegCU88yGUtb3elzJmVp
u8ZFlDK/PiGu4mlZ/yFl0qW1/4qMc8bLSwemF7r0bJtyynzYEnqYOyQEMnZmeVjVGv1Mrfvjrki4
MUcXl/QjVOWEYBpK9C4lWDpC9GwAjQMIf8KRy93N2ddfcS1sDsNgjz48gr4Om5G/9R6XJFx2V854
GPf9pd9fL5g/S+oSsIx4BmyGd73KwIjrwbU4l8duKaYM5SjBio7290LaUUn1Vjk7P1YPeaDJTX9E
IS25gTm6h2jDrpcNhvCkpGDV1KrxbKMwM23eVtR3CTkEE+Di7QnbyyvpULdUThK+A6+vGTD6Ym8k
Z/qJkti5FGjLriXgKVojaS4+2fOmnFfDtCgSiz5STX0E4Z381ZP6RtPkOKB3qUJQjktJkJ276nUh
vV5fkHy54TZx9tW67qdfIEx3j670cD7B2EZggQfPvvuDZoy1UFVQEGrA3E7ebqz1Fl0AFcV19ngJ
7C8OGsG3ZOtgf6OZclvUkaem6etRH1Rt2q+Ekn09OuWcE/2fzl3+CDHLGkbFdYZdnCAM5tQcaXF6
iTsr9SLywc5I4TIR2a3DfTmMh6+QOY8s0B0dRcmbkVO+pJwwbDJYZU3yKsnRBx0Co+6xX/6lyAZs
KjrAx6vZ2IJcIcK7tR9byVdfoAGo1bkc0oBwP3DJQAtj73shiUDcA2FVMhMzgXd/tDpCLYnfBiEN
ZSEXDjsiSLfWNb5X0RjgjVXcSfpp3s8yFrzzRowpPfUG0R7SBPzb4MY7BXof3nUvvU3QNqdd66Lu
cmHmV9nc1MP8Ip/R3q4HJcb/3xsqtMvhP33wLNFzgytyYvCIWRZeS1Kansgo9VB2tCEV7QlUTX+N
umV5uRL54yrrTmw5X8hm4UgTPsk4CoJ+hJD1NIpSZB0O9kKOr9cJzrMzVQGeHpwfsroNRUWibGoe
kZfQMEaCRqwEmDUnKCAUgPwLsh/Wio/9+4ujJwax8v1gjRGzN0+6vjuHAmCj6VDrpSEQvZzBtu4I
uKP7rIAda3EiwIOxnX1WmtMFI26DXj/2twLzodB9LD0dYHO+/k8jzXs8tYhSFkdrQfB0eF0ALWAk
9N6tjQ7H53yaerD0HbvRk5ObKHbMgmxsXHB+qX8W26yryNdXlOsyLOq8CnCear+9N86tPdw26o9Y
LR/QSt6OYvb6EwTF0DeLEZrpVkrFvj8j4CL2y4c+aqNAy7fG5hid44kqO3+GV1vFpX7zoi19z1QB
o96jFfj/90TqotBT5Tlp/4aVTDVxgNGMCd9ifLSnK9t1K+WOJ2d/5mmyUngNp4Iic37cplnZWZJW
1EcCO+wRTLibdZf2pF5pjuUgIeV8Khuujqa4kAnTw7pgqbh3rqEbvzeYXt4FRHSihCSjSU0aPThs
KNQVuVQ9HRGCD6Ec8nfGQ0iV7Ourkt3dtfE4y8WrLZB6GhAuNvLDv5CQJe0yXdT64aLxBUcmlmcA
uQqnOyIxW1N7ThWDWNBSJIQT5bhvM6knt63aAcc63WjXzZttVnLTu8+qHkFFIGPDfe6ePuU2RT09
2kMuWenVYcv+5z34jD5WAxVBRXqyMyJ7dXszzlteCcHXlkssV+LERXja8lKNUIzQH8PD5ERvz3aI
AaOOVr0y4GKmi1xaBthfpddv9KyimO2uPrRftZbfcPYUSdmyv1O3jR7lu3a1dJWICtC4uujPWAGD
4IXmTdCBi6C/J1tKDpzj8KcwFVqfNIZGxTo3Bk/9wRcQFlIJ92Adkxvo+nFuU9B+tI5ojDu98v9k
RezNecSOYTpw1O5eZ44e9oWuwCumVNRT6Fp97QSDy4Kjn1G3MByYajPn8fUH3ZTzw8PQqGpmaC0v
cQ63vtnlo0Nr9SwvBbuKkEQZUOK8soy2ZbaPe8WIipjbOu+TCrlEOlNtGaNJz2o8tLp/mnuGQd4b
INLROvaO0+k/2Ml8kgAO4lnfVIWeAGegeDLZCKQuVBAvyrbWxwnDiToJxLa9WBu5XiWJQWNe8Uge
uge6D5PuUygellykNQepqVaTUI+SUPlJoRzeDzqj+pN08cm0qxwG0PbyUgJxvGvzmPn0uetv0kPg
vzP9m5lDoTpKOcW08tZSvqxbIAFyu3RCbTGYOwt78rOY1w3P8wMghROOaaaz3S4GOoAvvhjZvV7P
lXhHDhpfDrUVzPIEh3+4zAxfSoaGpbBff8XTmITy1p/tGH3h662FNLMZuX8H8t9+umDqnvu2HdT5
FCh83jZbmdQO97+TMWOBvZo1QLbcowuWX5vuIfhEzhTYQ6iXoLnOAZbpfvfuEwIFC9S9XrT9l2X5
RzTmgz74ycBjfB10H3NYtsl4ibqp3jvMThi7UuXKak7nDBOny2rxQFyh96GNyG4VlJMcT3kumT+h
sfEJQ8yd3HRMx/P+/oJGmyUhOHADtjxITjC2qpMHu7pb/nIVmw6n64U2mtH161H9iwpOnBgmJnbH
Z88sHibKHUEwYWlj2S2LVApxBLDxBYSFm2ifiMNNQSe6iJaT+txCYZYbB3KTBhVbn22hglVHdhrs
Nl9/aD6TcuZ2hu4YD/AWOJC2DYoE0AwMlumufsFxrPRWgDI35Txw8R7X0FbSu8r0Mk2RSIc1483Q
iL6HivO4vRsn+4Sg8PhiGXzdW34MaSGmD3wLy9WW2pAVEGRHSfrsLeVDJhKsvRKDU8RHuCH7rALw
qEViTkWJsjuTxFOWoQyHHbMNDzZrK8LYDyneWRvGE7xP6iGaymijaS3p0ZZeq1qIrbctkxjjTdZh
oa0kOGV03qPdKChVIsut3xY9PNIam9czMJ7EaUrdm2iFgm7wE/qg3JJzrHzCmb0yXE4BKsXRRcC8
2XNy7BUnXQEkFFPQMvlGp/WZWUvRXoWYhmRguLtlNC0dqJaJITqVfxcPhulKUby5n1Oe6XBOXUlO
Z473+32SAmjfvlSWYoQge5CiZZuFOjd6JUvFdj4f2Dq4G2oCJM5CICLrfXuc0WbFDOMmI5HnaBNJ
jau/bPeoqJBdYuV5KmRk7DV3kYQy5TNmGQqSux9SZ748ZZ764ftv7dDnJ7IXqGtsV0ELaFBkil4Y
MuJvT24+YWgxWeiYD9rWcC3bk0wcS/7dsOwd+7qKsEa55y8qhS/HIrTgFblmN1LhzHFTw2u4Qjbx
ttQiV+MRuPeUK46cxytiLmOWVGu2E8Wek++BdHVDzCaSJSWppWqcCwuSOdZ74KB8OUIjj61/VpRq
pygQOu624KWErxYIlljfyTM+lCHOQSOze1mnkt4PT5pbHLMUpZ9REQi7poFzsB36zDkG4tOGWI50
TjuYjHP+8iPOMZjXh8F16u3HPH7lpeWrofb9DrH7AWcQClLH88K3Lwcqcc0+0ls9kqBAoaUV5tHC
krKLZommANaAWonktW/pbAjBWsvx4xs12pYRAa7KH4vOGuhQKmT5hb++OuPEUsWxHCIyxKiavTtF
FBMPBP/kvAhz9J0MA/T38gWPt058geADJkHw1Rqc2yRG9vq/mM0NMS9zXjfO4RLw43O0DWS+nAsl
2vjd01lDY7pmlBd6fKFsUaFA7CumD8+GpDXzvwln2lDHPbExjOY222cR0Mno0qudpySEC5sRIaj7
dfh8uAAfUaS1cbqAFoJjWuL8EbVZJPqkEp9DwrtDFsA1HSHoO9tkPmyiCF0PMTjMi7ACMFVMdE6M
0MEwPuKOyEjnytgVXAWaEg8l2iBE6j0D2TZAOMomxdI6vZtYr1BOfOhrJPYpCMlElioy6da2fxf2
CLL3cbPXCmqaY6ymuLHEn91yjbcouD0e7cxyIrv+9L/esHIUyTy3zhhzWn41j7uxfvMD1Z8DbKzJ
vjk87wwurB6OrBYCDcWMjoXVK59z5LHLjNBG9UaumbvZFdlvRwpVgrZgDpW7TTQcdlTwxg+6SWfH
gjz6/7NW3GsKClkRYp4nLF3pb00K9HKN/CTvANSowViS5Zx3UjDf4B7/T5ADWa+tMnB5e3q2X1ea
kE27Snjo1NiRbIKiPxynzIOJ2LBx/MQad2xuHY1C+3hJ1xlhTYCwTcx0l0nSXWhSpip1qQ9dQRV9
TdHXQ31bS2cKw1xxDFfyzcIyfMLz5mrVQ+4IfDWXJLAk3yLJDiwZUg44k8jVU3kkcYB/vouzh899
MUltEJPlsDJlq+54dbjiEpP1poO4XnDarBDWJ/DvtyeN5xFPwjZWhGJE+DxDt9tgR+OkB/w66x6P
nqya4cQcxbmXjcOC7B//pW+1O0Y8U/iSJ47DDcVSzqIIm+Dl4izg/7RscIQBPGej7ap47O9WgM3w
Zfe3DLHHQ5hKDr3UFy5hLOurzPkF4fYU/VvgANaTqZ/HmTF+5ZhPA8+mKWHlAV/WOHR2L6Looy8t
n+yW3/8+7IaNYzbOhj6h5TljberdUaaYlAPNEAwXZYbEQNmIO2F3EPdqdEbmy7bof92R5LrUFjvc
myEcTsImqPK+PY+ghK6fi90HSEbtiVgIhMuHZRMbRJEb0OeWiQCT48fgmmzEFbDz+tDr2DK4C5jz
wMci6qd6M4JAT1o/660J48iKMDifNMYQGk44KGJR4hzHLQbs/LRMzOpOtdwpleUw3nT0K4ojiq2V
vAn1WvHCGzrtlToA80yhqsS4pTxoZC+WDdCCwB9/eyoazvDSHIId6PxmfQCVbe9nnK7NTEc6mB9N
lLOCZ4riG33pv1GhcHWQdk8fgnxtWbRfEwg6SYHee3PA3poQzIgqVIkXmSPaklkhVVTEUtfLEkDO
Eu81g2ggL9XNY6oI6N3hsMmaovSPVB7x07XNBQdgnJ+HUgRiaWfNI7JVEtE0e9iV3sGzWTkk11nZ
LB903RA8tU+MBoGuPQ9t1sdMHqaC27YlpFwc6hmW57eDJehmjjNDA45OcsyImGU96RaIq5noUuoB
BYy+RjG/zddv9IvhCh+io3gK2Ub9FstromDDKdkH46DitxPa9ncj/PvwAKUqjO2/hz95RgsAsYzj
xi2wXYRVMinxpmK5BzaJHsDJ2kmEs5WvnqX7rsd7TL8re544pIW6SU66QC0dTCGo548k26RtRDNT
ssVV2JfFjMFFganHA8UyKfdKcBri3+ZQNT+GuRgJ0NhP8yu771nC2a9yrRvRKWqcK61cH3YaVBgr
1KnJk7d6bAWgdvKzHQc4yApuhZy0G7STCfZE9wZAyAFqN+uO67qZ6OMEQUYUhv9BYpPT8W9c6Tr2
gu1i/2u4XzsXZf76ZWfE65HKYm2co27K++pxYuQkWHm9rGvbNHuJNawuBUMNCm4+Yq+iGhL1GcfP
0KCSrBNpjYjfmdAdI2VO+PpqE8ZXEg4RELXOSpLClnJesA2I92fHT1H0xEJ3N7YSzSEZhHvGWyat
PDDqqqeY/ElPXWADXnmT8b2dSU8ST43QP5goIlXMD8zVRM/3iXsotaNCtxzV/7+2Cq/y0p4qyG21
G/BpXZdMYfxtCq/ACkTbjm2adKaWCXFynorEtz6Aiez5cRJe5PcFZt7mNClXU1qeU1hHBC5bzfBn
pPRolXaYFrqnW5jNkW952EZyCT1PyeKEEvn6gAH50pE4Lojb018j5Jg+G1msFNgpZ8jiQNQij1h4
B6Ng0kLnkt0fOz+Cd1RzYFEfxUrrl5Wp5Gc4pwZdqJG4sroKUizT7mMnWCg8qrvf//PXe/mvVYy3
PXJizKo3Gwuowem7qE2Z+2/BayyhXihXgYsJLLn+pnMp/HghGIcGlk+H611tX7b20ViP8stIxZ3W
HDrEnaSQzeytFXuO0zw0fr/u/0RW3Wp2/N+6HQHbkQ9qJJCiXwHVO6YqOEQcDpPaUHqOf4R2dUsW
b/fHkKU8Yrl/OD97S+1MKta26OKJdHN/MdJQHMKYF+5U7IqH21rfKRrJOZwFPbtvbdHz7CZIi5Uw
cW2yHqj4zaQ2WLF3RLOuAFhpUzx3O0VIozSHcqouUQKxLUEle+UdUalveCJzno1w03z4G+ApmU9f
BjxPOXHREF4wWHd40tO6mpDJjXHc1DI4goZpPTbfLETyAJTSS6BsmX7SiYq9UJf/MFuU8lNZcww7
zdh49hJXEx5fyt23TzvEVDz6ACzzZN6XBJvS3itcQK0q1Qt5XXBIae2WlaxcWZMPtNdR64DWKraE
MSi3VDDQtHuVms+o9hOZ21d15NzQWsizKLP61j/fIZEElTGpOVEKKJhCmlXSIdfrnt+0H77rfp1b
+BNiOg4tXZ7VnABApcv/n2ZoUNZmmrW1bFdYgvmAXgcA6pzalBZzahLl8YV08AHqUhZ+chVI+/EB
NNYoWwTwYqTRw9aet9zwOaq4PSWusGpjVeIOQNfsm5t+xzFytSJA7WJeCUOpxcGgHw4lQHS4h9BK
xP1DK9GwJIKmsTS+xefD2butdOWEJ+UOhw30nCX36e0MsAhpoRLKs48oRgXvotjZzAloYDhzHQ11
okTOj54ote+JG8jNBHF716ZLMIxCrAhg/jpyBRSomWRxkb16S6CR1gaS9w+grGnwGE13CGhsnuK+
ka9oWHG/L+RKdMx13H/DGtllYrR0lL6VVQl7ogHsA/mc/O+RmcPyMSG0DZpKt6v4u3ciKNb1gmIA
MeO8+q7BPC+QmUSp4qRne55SXKKbvIXfAzT4kWnE+CrhX5P7IFbISMuO71ETCg3L4v9T9RzBJ+j8
6expIUwzuP85hQXv5iYEHDl1nIaUzE57DKp9cnP8AKcfEso8p+o/9gAgve7u9GMfjo4y1YUfzKaX
D6/3unpRzsJqIOFD8dLueOqBwBC8Tjv44AmXAAFvJk064f6cXe2rffO9+pI1kx3CIVsY9bKjV9CA
djCw0QpdkSDlrIJsDsnmqkLBUGjUC9dnLFwNKvqHL1nejuooIyvNCilLyywS63B7/jypCpzRMkzQ
AFp4xlQ8nPktsoJOMXDLWoFUStqMlLOjSS9wktuugiVmfNGdsmNW4WjKI2LwONy829KXtusdXvHl
HE7xhumarhk9fTggcwCyzH6b/JvkDxb1ljj564LkU5IxXCJiNja56jzc0Q3uL7625K+xoYNRljUV
vFxoP5fmHE8IpBpRwnpIYX0wTsTXl938iQgMQbz+kLOo1ODn9WHUYwsuDNb7FZysNoR9qALJicXe
SAIYBzq6kWNxN0sLaFTDJyx+cN+im3v/GU3TYuZf5jtvLRbxZnDww7iJZShl6wAF3kdSIumKTlgK
ZyWchieYWLMs2wCHpP1+AlKiU4esAqTFwBXpOQ3vzpf8fNtAYnTHzF/uAZbsVeh4jU8uVCvuu1cR
yqcec3fdC8QQzzCDHsrKxXsWMClsbHsVm8ZcBFJLptRG7u6IszZuk0fFuAP9vuzjdBCri3S9nOUK
Gq7gz7aF1ohljLQ64dUrHwmH7lMrAYb8TM/1aOK7QT7oVEsOLUxtPoRFCIHgbjKJwrAFu3ul0DEe
3MeteoPPtKUTuYt0rvqqM3Wh4JinhhcPMoEES9xIYEXl6vke0/8xfaV/U1GID2vBqAlbciNOyG/p
r0qEs3lXaLT/+QUpbVcOf/5tL5s3vtd6IQK9uPtaU6/eh3NlQykqGims9oTzIiRwEatV1ZJ50afF
dq/Iy+RzebJf7ahqQtlyarCfWeZX7Xu/fFIk1L6SDlpvztfRvtlxwmqRIcZSx4xOzC8o9pqctf+N
h872fh0gKvbfBxVDWRDjN01UbYqvmcJKAKOvmHHdyj0+2WDGy7DXEKYsDHZ8CWVxse8DYdF0uhNS
vZNu2IEbhG5cmJBW9VvhaqMwgEBQVfj3CNzHcGD2Nxw8kcbHh/KobGTS86rFmW/U+ftwL248XBFu
D7C+lY0IabuBPnZdV9hRPrzzOatJh9G6xdPjjxpdXHaisl5stCXymZ2FHxBHDeHHgHvfCjA0vtCB
JW6msw2duFdjpdjDFiO+H/t4USLQyWtnzLO6NX0JcJaL6gqkvyKwmPm1W3TJ/MYNGtN/bealrQcy
rCwjMjwKA+ZNc2jzzxRcf7W6D/0UEoFN7oxFjv8wnKeZBgKdqm0tcMpClPqLfQx3EzOuyWvneTwf
vjOoM1dJ0OOi3wBWKo5KiyvfyB/q0uHOxAY7kmQMW1wdGVsEHzJNzZzOQ3ljYoBWEWIVbfE1TnEg
DNNWclnazX1oaDMMtnEMqn/pqt1bT3n5YHN4JDv7r37srfcoF7X2f2RKccy3RyFymwu8UV6sILi7
xJPOPmjtmiGuAdpm0Y0q66ETONZ+JCdfbRMzjXQX8ni6WIDmFxY5/v+aY5P60/9n0LbZCx8TGkX5
uPgEsxZ6++3uGRrVe/HVtmtaS+qvlhFMRyTPF3GkkfbP0k32ZFvyiakx99qx4ZdyINnd54Qd3vzG
jY0U5n77g0seGqu7uQ+MbTpXHnv7Lg6M4RlOoB+C4LrljPeu2oWtC2r/y5j1kf5697uoQgoPgJRg
vBWRqVK3fpB+pSi393x5TVzH6vz3/JnQfUDtDNA/8b96jS84koyhLc8wfdO/zkPfXudGrIuPdkmd
M9vaalP9XSi8/VizSqz1Kd9HFjhAf3W09pHEmJjiXAnaXYX9rVtpfaAM2yvHbGcczcJpkRignPd5
Id8AKAspvTosZ8pjG2BXwOPWW4tLWcIwwHBk/aNOH6SprGf3nd2D0ae2o5SWzLiJZ8ZGSVyhFwww
QflOloCX6+bPlpLfkmy+xyAPuq+aedKcSD/0GapmjLrxyBFhI7PFWEDnIdB0bK9Bgnaa1+0wZ+P8
DNhLr2s3giv077tmUl1qYWVxjVlfH59Eq5A9T+MvjgW8PSx5JBfNDI6muhoL22aCb9XvFQAfO4ed
zv+EMKJs034wpwYcBqPX4MS4VeaWJWzQ2PjHZGLAVYd9mwK2ny2ln5FnluWMJwjfu+0NV0TJpbFa
E1vxTYgfsvh566SEipcDZVJJSkvwj8C2PGjLs4yuC/HalG7DYG7XLMgu/usyYd+ndjbwL0Y1a062
euhiSKmcWPC13OC34ua4Hy9BhQ5MLL3u48XNZrUH/airRx4mg3akLz+20IJ9cVYKSqfjIWUAk8jo
08Q2igyIwKnAV2rNa4dS/yijjNgchbvnf/oqFlMjDOk8WQnCnupT5NfwVK2MJB+UmYvN6chnGSRI
hS+tNmCTkLWS9GjqyI8ZqFbDZ9O1FuRsEuLSyVpf2vlVBePlLDz5od0574aoCyIyBXxKiNP+k+EQ
u1YGEm10EO53JFz9YVdBztfgbb9CACwYFNhjsFeBq9AWmo9fpjzbjbcikdG8bq1l2y+DihCUHbui
nz3NRGW/vmGFMUk1eOrSC5I1PDApAP9157HnyT8jfGCo1bQkBJAiOC4ctIETxIjFzyG5xGjH1BxQ
bKTIBUMVGNFw1CmWplLaHLQCdm12j8rykUiGyV++ZZftYnet2/zTCsALrwqavAXUEVNjHM6Qr+0k
razeP1a/dDmpddse7iLcqAXoDdm1VV5uf9R+Cbq0jT4PVTNiYzuDaJkhRyptTI+L/OB/XxLVIFIM
wpqxWxQMceW6TjlT7ZZHHkyX1tqtkgnwtW7ClYU7cNkcLeVfBopeSSHVU5lLBwfTtdcGnMoVnBzv
5aNrVaCBPntsBwnevatGQTwHQhkXvjk3YCPxIQrz+u1o+NFxWNaL8OaDy6UDRNtiABLYcSsNYT4B
+DKj2msw4VxmsGGqZ4ucwv1CPSnaQfWRvEvrNVqGL/va9P6kRPVzV4ODLBryChWKc+t1zQO31FkH
n1b/b3dvo/swdnkdibSz4y+QWq9vt3khn5+s9Ly0NUEBKG8wyjQbZC0oJp7jYdTKXo3KV8GQtUC3
Q9Q1hvPEGJ/EDebNz3D1V3J09qz/FBjq6JSOFqGfE4kJUSuqDIYzvCxPx90Pd54NzgOlro1j5gzW
DC+oHvazfnS6vihO+mfc8wZWa1Mp5iZ0zLxjvk5B9JKhmRsIiwymPC9ILo63KD/OZy1f+bL03IB6
x3Gka9VF9mSZ04S9QmRLXNzZ2LwvyfnYNq6rWH16mF96nTYMHrfSJ5OmwweEs1afRqpvoyMcmxI7
j7lMdOfOvjb891MpfzBFve78E+a1XygPKi8akozN/rm2iGcJcbZXeM4tMrlr0rBCtaqDJ2Du96U1
rmytko6XhdMHbjNdyEsrUeZav1wvYeacvpC2KFhocFGO1pVD8gXg1BLp5n5gczdAlHkfZRFeqAl0
/GxzziCNaR4X+5x/+/pleL9JtJTuGnMJn0GiubcH1YGNK5yqJN7WAshh22S0UjEefoMgIhht0dFA
IamBeK4zo80gkT+oId1X725l/SJ11kBRZBgrExGo8UFqavht6nFHTC3Irpx9nIqPjh4E1NzFVxN8
uADnh3PSBzb9srr8ACLDDx54qkqw7J//0gVBnStllAD/9RfUxj12bpC4ak4joItEXB10BXzfaRoK
rkMV3dLOc08vGYWczYHfwlFLW8klyXjOZjsIberPBVDFhqg8qgyf3IqvWtRiGYG0dxDAS39ZZ/mF
KZ2+CplAHHR+50vf1iqHEKq3LDlqCOSbfT5NcdoDUQ4ssXUm6AlgJZzB7zXtnWq/aDQrQWx9s424
2ljP9oo8usgyym06XmA1fD1I0lfv7EJqJRLieAm0UtiXTWDjqE6GYNNsNxfCFjRMPvRYDRSdNY6D
zQkdcbwDmF53UQrZQnkyqyyp/O/7hUCxh96GDrxWZoCXUcBRZYKKPfvyIJ44/qIGQJLMO3yqmCsy
aOhzmuAGIbw0/ADDlL/55ep0I44jgJzIANRyRTm6W+mfKTSDJJx7YY9uIhhp2tHmPAJ7/0abt4cJ
u1/A8CJLmbw05LC2EZnSgOWFRAqftiUMfT+4AMsIjj1qf7m4VvH30yMW+G3MRiOndKnAJNhQ+60j
rc8IbGJldrCiwUf2F8VGryuH2w9572yFB5HV8iaLeY66YT0/M9yVxJEZ5rpMIro1j9DQGy08/Q/o
rN7kHBDSk9dkr17EAT3NnXqoqy6SDC79vdA7O8IAc80r8fZ4IL1YZnF0yT++NjRrsxe25HlgQLv/
oImn0ASwKZt4sn3qvqtWAp/HVsCc8DinxHdjJKoCB++mrPt6lyJZzyHaOvxPC56RTJT5CY5pwwVt
tIw1Z1/ZAlq3fWuNYZZwoJreZSV/x58X88DNhIcsKPATE/FPZzWlKc/g82RdfcraguppmMrKAaPZ
2EDjadb8X2glDsUOer1VD6sRj93sqTeITU/Q/1MqhJJwBx8JC7uRNDgqSNkoBTF7DAV1ePJIdsww
A49ISceNwp7aYurYxNWez4aRbyd2n5dyedqrwQbwcpcLXaQudIy+3TFtwdG00E3iv4wxDYhmc1rg
/gC1y49wzheDL4sjPq7ONmQq2LqebzZjkyi/GQMOl2IeJIbXV2Yy91ys82kcrAnRGJDGDH3y+iMf
1qOb35UX4yENIhVNL3VuY4A/GT61if+q8HfOUv8tk2lE+R855eYQwyrWe/1ziHH+kjYHHzgOZw62
2X6n63rxVKO9Ep8JIFgN4wZQoSJeKAj/mHjo5osVRQigfcEp6am04IyV/loN6iXG44hcptrBrELd
wJYtzEwdHaDjdiAzqguKxgH/qIW6DEWdm444n23Gdduj6Zvyhb0b0JWdicFgp68YJg0IQ/L44WWt
gyklUTsBOZpaiXxlqFDyk/qXZC9+hnMASxIeXspQlBQcqaSi5nxDyn4w4UqtnWxrwjXeOK8kUiSm
JLUgYJNjeDpjibE5Je2IYPUbDuHH48DfZRRf/yy15Aux23aX/tsNIF/YiGqRFRd+tkVbVYYAiqHw
VsRk+4qoGrTYLHc8oPg9ncltPEmIwJPNwmpoBm+CKYf5CLQCEjakMX+o2JgQlWlkqEQakHHRT/JM
cMrOp62upXHb09cip8qbPF9cXx/760Af1WPr1lBqXAGEueJW+DNPxfiQ1wtPD7y+havylg+xizCG
eU2TVw1I2toESH5TVc3bzJUgBdqtIi4pZO1Rc4gFfWMVlBtVTSyLlgBVZoh2pn6rDsZ4XeFPF4bO
6t0yqy+egOE6eAit2Ze4IDIDRF41rhgDpxu8NVIavli9YKGqGm7OHLqZou5qgLvW+iLcA39U7X8N
DjF1q4SyrpfLm09vPKivCezeEsaS7vX+QUR61X9Rx4Rj1JDaXsYwBmWngpFm5mtrPCO1eu8nCsP8
tvuFaYI+JQXb405MbmdHWiWPEwhE4VHH10yNeC7GKgmlFObcxTZdzrEAlfdYr60Ck5Q9mv9FWOr7
vDqkDWwU82RGkvADQdO09ivS+HvbOgkxS7LRNkh/PWNDwC7fyUUKu1BkPHFp1QD5fatG8qbK72Nm
plIH/9YAUVBxRepOO2NhAVBuadnpVj5Dp9AlNVl/xKELVEHdIVr9dyTkHkif3nQKo3UYw7DeeUiq
cyttxBQCTK8dP+/HOLcOuED/08hvALhySknDovBW3T82P06khOgWho7nnBYaymWwbUnBOdQnLOi0
Rc6rCXf1JkUj1FXUH8U4g2bRfoe0M79G0O86iuXQRBBhfKa3DxidH7P5KdRBtqO6GFhXn5NOifLd
ZQ0zDUHGHPZbuAhz9ZyjiVDGAyxg6KH077ExNvoEcDKR29uXQ3TNPMi0UW4/r/d01WDj7GkZzMA4
fuXZ3JRutPVI/ogTjNEy5/GTOKwi2kyk0bBeptYkGEEJiL6pmphlQkEGCK7qBK2ksc2g4LSNUqAH
f4tiPHr2m6LpDqxRQfaU7zBA8Yw22hn0BBGkKvggNkoxZCFAMSEXv1b939mPDa0NE997gwQCF7ft
3xvcTXQLeh2yKXq0vc4EZQ9x6iE2rWDy/gxpA6viM0lfYwSBJ3Eo+Inuhlu0WZPjzdTfaqmygX+L
c2dJ3eqYeG+/OROIgm4+rUJbfEtD1HLaEVL/KgxBhMd+SeIJkyAcjSqRp6oirk3EWL84ctmnoCde
kV070XxbP2trqqB0dN54dl106XkDbQnQzNnSNQqlnlkTlVgXhANtwHzj9Z93uC8Tih++sOb1ylF8
7Jk02iMxsfX8zbyRmexYWt46Me3tKcDacZb/DOt1s538TmVxz4xkaxC9mPa9Q4U2HSpACdlecano
tHb+DkDXxe2jjhuU8KflJSz3GsKiCD1Wpem9+QJxAyJDVNVUARYiuSA3yX/fd33AmZWbNrM+PIwm
pe/JIYnDF1GU7pMV/ogr6CeGJdULycgnELQVsQ+YapEHl+2F8nQqbJM7PRpVmeyu/srgHD2KeyCM
4dYyWr1P5AJZTjwwUy/KUi0bWiVbnuftvrrQb0fe+8ne/vBBM9rGy3Ej9Hg6UVWKYprqOfpqds9+
yZINxHEfgvWL9GLOBH+4DOERHUGt5hMC71rfkuhCEsXxuXkzS9pY6hdiXl77UTTCK4g9FQP2RuVO
9nd6b7ZPwBnIYZxUo3lsa/+o5UiYDBD2yJ+JmKU+ZVDm3qx/OyxaPbVuB758Yufmsk9Ugs7ZZCuP
6Hny4y+UgyB+LYXgzjfuGSeqBPa3quJFpVLMLXOuAQOrnutLvNbyU8hPgLaNmbSkxNNiE8swP/LP
Jml7qeJta6MCocLXU1hKNwfAAJVGTm84wCn6TYm5ybKW5HApKHh2bp4mptRXSQGrCBr2GjvwTtl5
Y4KNck0Rz/GRd3WLbDN7TsCM3dJ1ETXPQGcydMF6ZVsJn3qabr1Qrb9zy8XibnRTCReyxFxGncNV
WK+SxRzHZIPOnflqzmTzPsqqj9hhBqjb6Mln765kb35cZNgAPqCmsXiHNSIZuiApWHW04yZL328Q
PESBkwlcweRgPLLwciIYklO57ti5PFq2NkwAl39LO7x7qqaAUPqNaGaUq9mRJ/ez0Qs/QxjFpxB5
BKkPhwkxP7bJfqFV1jlNH7dtdRj4gdpsw7WTXA0CiyKKqHk7na0/WmQvOz9zulM6I1f89SjXCznn
N5PWWIFJMI9n72aDBhJodxpK3KxT7Kw+5RI4mhR7lN1hyTzSrp9UeV6eNgudA+fH8c0D0kiPeW1h
MUTW/UvPzeYY0GpQM9uwVhav2L1A5TJhogU88lx35Zpvy9e9O1eNXtr3UHeywjJBVXHUOPkomKSU
3JHp/+X/3vTe4MN0MqCIIwnIjITRiRtNchYhMKzFuaAObQ5aCFeAaiRl7RCJAJWKIUERaN6mJa9r
roBSHPxU2Vc7cFo6biP+WrAdrmtsNofv7qONHuXR6Gu1R6Bb/ZNtXztHeTxkPwTtHRJRaGHawR1u
hbr0LC5xletLC636v3dW4jMLlaNqBssqOzlioqYrpR0d3n1k18GHT/HTlSVGYOe9muBsiNKNBsOT
R88Ml95wc3RZ5JTKEa3WTtTfmYMoJwO8QtF5feZ1S/lyIKnv75uT2KQ4VMxu2qi022A0hBmla6JA
YvaIJmS/W6N1aGlGOmE0fRZInr9UoCjNeKZGGA0G6rfnZYKI0HFrCG/v6e4XGfmFTVz1AkNL+Iwl
MOXRGr52Ze0C9yCyfz6kqmVWk4TCol6PahRIO6hYLQz419TWC9iHi8ecn2xv9N5VjUrPkQbcyYjj
jpPRzvghwCofJHFI9kRDbDFYArjMDDJ6IQQQ3c+J0yA1ejpvbzqq2oQMSwqADTVcjwjqCgWtjrEl
elHMLIybpGh/GnxUe6kg+k+VrCSJCBW8irNBvDqrLQMfcjfti4lXR6wCGevGWvIC7OZJYblnwbW4
EVu3TafHTlw6S02LjSGVGLcsLyWn6IE0S6kaz5CBSdgOWZJB3OmcZZCRV1zISEmJ/L7SqfcZJ2Z4
k+SGe1TPYxR7WRE9Z5nzl9iH66gL3m7m5wnb0kPD/uJXP/sQ6f9tQ+EAubccX3CDbhOYx+YNSA6w
sQ0he1QgHQNX6ypDLT2x3k6+JQDgbE0Tm7KERcZuDQHXQ8/l2v25pl2NX7R6wQI9FRGrszv2iwN/
ylxre4B1acY2ia6crEWwSsvHWwQHjvwKjzkiYtHJSUwwipkxuE8Z67KHJDwI6OPJ7yQR74H2IyZo
zTQd59sBLrIFYR4OUBCC++3giDc4sFPuGnDpLvcEOYBMqEgb9Gh7EUXjTD1AUehqPOOEV2PHc3M3
adBdCjxKe0xy8YMo2U2QUZKB5pUqoQAOBkoiHAWG5Ns2PWZV0rQlfraKiZmwOWHJQs9HoF54t8Zn
bHV3mFAbbss926f949JBdQDKRWTKFjf9OOBtVOF5w+RfWZ6Ojf4InMDZsCOcoc9lPfdvjkYQQDcD
s8kZxa/YhltfUuM8zZcMqWQIYNFKmMhEY85gaUiMjW42bWRhpuK8+ybq8yJbYBwLPEF32rOWfS52
KjtLO3ObG3lhrd9kV5Ajw5V1acYbWweuxm9OrpBHEeGRx2SBPl3R6PU1afJ06PaUkFiyhp4TJell
fVI0BL1fuH4EqMpo9P6segGkMQGs39ZoI4+2H1DFihnhqepfaeCSm2cdw/2tN5ShEbMagDdyU9nh
0zvA5sO+DPPWgkoimu46+HKvkALkxrwTHupASEkaybd8GP9JRPiUvSy3yojZXC6GCCtZBGiAdXOJ
aSupCFypjeKMOdEQMEKOv4NYIplr9TunNST0YJLnf/ap7Yvvsys7uT6aK06h1hd6/ypA+KsTVjRs
VQAq6MFGt6eG3xQoTadcUXAIRTIDXH2XOEKiD2UHqTH+LchlumC4Al9IeK2N2W4+ASA5KR58Amhe
FLRMbtUbuw3a/yWHOAMSnR7QWoLzSmcDBMqhmxI5O95bNDb7EfTByGp1PlIulgPgOwagwcC8V1qI
JUi4iG/Dl2tIK6CJXH3plzgNtF8h64KnjiEIcLqbrVBjAQ5jtb37YzZGf9tRPMuakLrE/Fn1xxZU
kCRslYLqFZ1TgmPyZKLocDcHI0exkZglK59fjb0Uyftq3PLQz6BV4sW89+iyOz9i/3zJHpsGqPDr
4WfY3gEZ5y/cneMb6ZOfSC8YwSIqzjLHp2q3c0Yfxl6YqytRLJOoduXAJJAauo07+42Mkyp6gBtf
DKy90GajRkPTxSyfpjEHyUdt8hlNPdwwZT5dDLlVWTLbgPJDuxFlhWm2RJBbLK0f/RyrPwVm+/6Y
WcHiS1JYiK9g9a6jbxDSjANEDHfay9ThHtZv2vBCQnUc41BJFty4BlNyrqXYirMXCf7cdwf60yn5
rGXa9Bx+UanStwviD6R2uB8QNRMQQTR1pu1ivqiaTuZ8VMixdYLW4FdxNJqHKdINCUEHzK5HmWO6
0VoDBpz9iy49tm80r7fpbyF9o2CrNH+9RwBjrDCbNntRMgfCgwgjFyBxuhhLvaML8YOWdtm2rrd7
5Hq8k9UbWzaOVczdf/cbClcQUn8trqJm9IewybPae0Y61ZkX96wbgMRoUzF6V12GaxDT8/m/8aSz
jEk5As3Z/Dd8/KWW8iF9Aj7qRb5ARPMi+fqE257ixD5z3EE6CYGfPNOG6d4PqkO76FYqCQ/Pp8HP
vY5m48Oh7PuYGpOZvBpHuyVUmRjKysysoiqnmRHZIzFCYv0j79r54LfaC8gJptw1xp89d/lPwdQW
3uU4WvcCc1IcGKpjxPUW9kgYXVWKurLYqogwFB0rzp0ORyhMCjYD2Gdc7eZpjmWrI2V8tD+Us6UN
edTNCBcAi4LBhrb8IoHCHVtHICeJT6OQywDPnOcGREOh+Q1CUchtYgwKX7h299QKNFlX2nzqP12v
60HL1D0YZd4Rrz0soUQNUGdOfiZz2BtbqqnXwngw5w6s1XozceXkuVwdsbLqgwjkxPSGdOQQVO8x
s2POi4CYyw/5iUNVVXx6hf7yVKA+brZoSxPdyyl4c8MR7q89gKBl4EjHR9RCTNH0mUP5i9A+1DgR
bHDSeEs/b17nvd8Z8DfaQHXxDJSzrDWka4LlaASKoYxt4NzsRF79Jb5dMBzmGAf8YNmPBKFo1tol
0mV5PCCbCR76EmW4csYBwEfyN+fyheK3047ABw9kcCULjyXYXrr68shAW7DUSZaDeKkHbI5n52rp
b7BmchMkM5aFetGUaRL0i+A4hqM/2k2D+ynmzaRKtGO7ISnl4ErXFFuvvEOVGC0NWkC7xiOjVs0T
bUgGMpKJRm12puSeLzG+vgxrxGQ7ZfhWA9zoZ52JdHNTFurTSLCRCfSrc0y1YuyQlSu4ki4dWY3M
ulrny6wBPdltf9O1TzTQMKsL1E/ilRWOu+cl9VogG0wdpJkITmci8MCKfUUlnQB6hPsvEfcTMNI5
6xmDX9sWO3UrJirv8ZCmhb2F0q/rLsXF1foT9MbDt7nsWkxPPnqdDwDkfWGjRF48sLyDLW4sonMm
VNYbNgworyQt33FnfFp5boQfh3N79JZMkfqgPgFXuO7HsmB6PcDeLlr+1Z6uLfXQhykhJkx8U5GL
aZgJ/p09NchAVwoo8DKRBfOGgJubs60jBxT1GZZ7n0PwLqdH9FW0QKRVxb0lJZU0DlVHKx6hylvh
Lp+MC5SVdbDInUP7Sk71JADKZRTLVzDGbSOM/B2kIYQ3GUe30kYfwv2VVsGU37jSco4TZWT2lidb
HAU0yFfPQYE45xmJnA4T+aL7IPfgn0MtS94BEelDpgIO5TotsCI+n7xmrfmIenRRTd//svY71MjS
DHXH2mhEAbagq/vkhaPcVO3LmltC6rCYrkagXbq8ZhEoteGzgXQQK0CwF+aEj7OSpNEIqpYJgxVN
pevJxKgT0Mu2WLhkdjsVfZr/szlJVZv+5mSM6nIDrpUZNXq0yrnD8eigvAP+9GGPEdUxbwi5eZxx
BVASo7MtXiqHfCkCq+Abno2Tm8NkRzXwW/ShqCErEakdgxPq/+PvPWnL7OCqJId/LedlsaSppKxS
hjB7WgH4xGF3gfZv6edm3/aQHbCelxqHp1pa/LgSObMdkv6l0wGO4WLK9JLArEFSrT8FeJzuNe2W
8SNvAFdbdTAkW7EXSNqzitGOSs6FnJ7ho09E0bt/n570tdYh8NXwsLwWzUG2zmKASHaIAliPFp5N
xq7wuBIPEmbu8rCuvoifOSpOH0hzbLykB+4pdaMemResUsDM2g7TbQMGEbXRxjGBqbn/Y7gEIQ4W
L+oyYCgWrWTD/i6rDn6q8QFUMypV/5JZzF53H7W8xXrkGbYVptNE7Algp+vQQ/s6JrPBApdrVt9K
VzHn+xUcLrlzD9eIPOVuthaWUronK9lPUFqMtByVlicXUVyuYQhDxlSzi7p3Z05Fp7rVdOD3TuHb
S+pnqe73eisTeMVuEdRBX9JpmZtXSHsIpEb/I5x7iEGS/RiB0qWzjS3dKZ6ht7BEsIM7WO4giIGg
m5TkYGV0F8tk6jN0NPB2c6qKOQX1HLgvG6oOlqaVjOhycMzVT+XQFhFgrmpef3SFS5yBBNanbFAg
ipBx0XERL6Zy/ndxpiwRWoXZ5FSR88wu6zeoSdXt/M2jju/C5Ihf0LWXZuIWjReflrxtBuTtTUDN
RMpDUoEH9QIjOyyIpCQeh1fR/zLOG+wtmvF3+HxXr9FC+OeQCPEdaOxjQt+K+Ef5ozC15llZwvcg
7TymYf+LtzazQcnhuZgcKQugO+6OtsuHLa0z3tfDzzmjrTHyCWsdKRPamTWgdNZqV1BhaIfiqzeQ
l75hQVdnUftu78jpfg/TqgBsnrAx+98LNI3StsWUUnNfpGcPLobPpWgBcE9I1L3thdPRkggpEu4z
hojb0VpJrdINSWmnunQgIb4nHRSctmpbB2tFlTGhWhokpNUxhoS4G6URw2dyBeOVRSbxL7mZhItJ
xLWRpC3oEvgQJnZujYjCk1OBe7R7O9Bq3i4si8lmwvQ8CrtHk8bZ7tFjC7EwIQhldNYvj05cqpzv
+sN4/lxQhQmAdrBRFMNz103heWjSImgG2CWtG+BNY63A6jbszhyCBhsS8rj4GNXPJny83TLNEpX0
FMSwRzMCyCI6gDg1rNtdK9Ww025Lrux9sWaFVbEpyFFtKJXqinAPas4dXWSPUKMU3UZXYj0eF+qS
Pig8DtNmlkiefw/NX9d3wTl8euO3UE8fu7wqfHhr9qXZi7jGwkGFg5flDjC4dytSwVrj8YI+kygz
7jng1l1G6MGjwVpCTRhXRSY+GcRaO2SqT/ZqPCZyDL6NJHOKHHxG5xua2dCVBfpE4/o03Qo9tjx9
x7+UldqnrbjHqCnuAk7mgT9djqlpgEQQFHAkB3ZZoJsHRAJBcy7wSVHHq771vusyCf/osJ209bMI
wnrIjGURIvf2WA9iYnSoepN4wsKpIM/LFe7gcu12+lDdO6VmcWvDFdpSJz3MMrfXM8nMhCOGSneo
ijRin56E21Wxd9ym52t3usgIfVWK1sju0bAGl/EOVOaXyaRd4I7tev2/YVDGX2bwhYRgHxRzlCde
8TYqjo7NCfB8lisDTHSkNQittJKj0xQKPDFFGEbbMPl5jCqjfN24ypYiHsV7BRfszVSir0YkKlPY
uEld2InkmKGvd9IRre8dt7ea/McHPttO1bbQk9RijLrlP5gjAtKU7Lg0USSf5TvV9jm+zA5dSr1F
cmSdDVteuVsfIRUKaDdg2KIvbY1KKWnIU3tuCub++XABvVN/6DgZzpVzHVAEG7aysIPex4erpRWc
RpxY3ldXiqXtKv4W3/T+cFeVk+7FbN1kcfU0bi30Uns1Y/S8LdJTFXNlahmX8phycb1d7099FYoA
BO/eSe5R/QA+MKfrmMMFlaE8yTMmpCLis2DomXM9PalK3Jia0faifZgnSPWkKjLB5kaIVgM6L5oA
1ohPhgQvuOD/peIHXq7Hzmx7VCtWLp+lz9MC2zml7NSuzS9NaBRgrFf8xnpN7DhHWYjC4S2H5rwp
22vFqSYFHhBr6SZYzhGkvrE420yWIH6jtGSq+gTMMhKCKdGxU0Gw+wZ4mOEniqx8+Cf7qF0tFuIG
GkKhV3k8y/pZPffd65Ek9PWzDYPEY0gwkEZI/wU6Dpsdes1Sh4PJf8S6fSdoDI8nOZn/pRjGpx5V
mpmKYOf56dLQw0p+vIEiYC5h0eRFjEv8ycsQmqfiEGEry94Hd+eIlFhNSLNQWs/coJBYaAjhbzoe
NWx7AKxoXYDrno+a4DGyvCPHG4zvmy9IppdUrWRh3EfzNr9tKgQo3rHUO/sod3G3XQeObWotbUar
59fNR6csmh70oE6cFy9lXllmDr6NVMzIlPVKtyvZeP0TAuhk7F6wIQDOliE5VfT9UcbdO4bHFgyc
8BtYPBqI6lmFK06ZSYHOLCTxHTO6rX7h8pqA8e17jlG/fGNGohpNr3cY1ED6Ar33Jo0euagCCMn+
BdS+MCyiogGRvSHl+Ml18ah25N3A84prWbt4fGz7zTbOPQP8RjTlNZk0vFYTcGPaWgL1FleBDL4M
+OvMYwm4dY79EVxRb+/Bu7zLjEYI2ke0R0/Yt1Sk0RiPqs4s8e8MoAgrPxMpNbanSsYAgO79sPAK
xlpDTYRYTk1DME/8D4VqFhyl1F42XGUfK9pd9unvW801L8d5HeDNIHyCSuU0DUjQOqJDwflzT3Gd
oXPsJQkL8jZbc7iDJDdSjhQUb6rZKXzCCWM2N8WuNPPk0vG4t+4DnQlFmPKsN6BMbmE3um65zeYL
Xu6OCIK2bUERftMrz89h/AwfUDMW6WmCcYBdUGz/jvlbqXOX9ACn/jRxvBmYPsboLmopPxCpKVVE
uFMlt6F7TGWilur8seXga2/0XsxSXNy4ox2+drPuVx0bWrjKVNPGEpME699Q7mjVj64CeJNA0ca9
xPmfBCp/FmmQOhGLxwjFjVbh9xg/wg/4PWEzNj6RphpIA78GKbn9ijKrGR5FvH7HHgJ6fAV2G5q3
TyApBdmley+tOxuHc2FhXd8XqwUIVmaMCTQUCfHONteLubzWITKD8l0pRzTBd0TKAwFHeQ19xKYb
DlwofpWF9Zqd3TGW9YKg1Ml8XqLZnMtObMB/xIlqIPs8p4t3dx5znZgpiEuh1dKv/v4ypd2fvWNH
aHJ+sg3MmB9Xu0Qr4ccjbjiFEDWnukPHqMzvCHt17ypa0t5k8L/LMyfcCMPEse5HipZzugePfdyM
nYn9RZh+6Ac8mDFjAKEa4PxP34rxf744UmN0gIImLOPK3VTvQBa1C3QqX3YWlZ7xQYnNT+OTJ2z2
RlliARkGWqhfJzLp6BPB/7J0HViM4zxLNX5q6Sb9m4vdaUCA5ap7UOgzAH3C2TODwuYtp/2FEnT7
OHRj7tz22O/VbI/ZSWS0NqL/L8V0qm/eab64c5HLf3b3ix4Jn5h/EOTtq4cfvlljb+PXN4fqrUY8
7XPhMmKvA4onW8R1lZf5mB2cleFZrYjezaPmx6OWe9ZbP6j3o+KliUaD9CP2jcdQSStmZBl+xUmU
1ls4DIUpmwctkdpa0ZAgzd/Uncc7pgPEBv2scSy8JmfctNYZQ278/OoS4hmg72Fi5WvTLUNGL3ch
xk3WuK4wsL2L7mOWipR6Jr4i+lJgnR8HFnjiGkekZ5S+yY4LLiNafTSinB7N0owANb3HrhdtqtR+
/5iuut9cqAchG029i10XCv0AOI2djV5CoM8Ems9R16ncBxvuoN9gRgWHU+vxUPRZp9mrY9tGCpJS
0Ld4cZ2h8FXud2BsutRiv4db5yO2xsGgAVWj8RlmRjiqnxEeseV3RjCZWPhKJXE6PuaZfGf0kAwR
394HOT6QuEwj4iHKaglatgkp2R4vqTbDv0ewQb3AK7F9fsbp/YkMW84w9lTVqlMOkaKX2/n9XTCz
NHilVSDJuDhgF1+zAuw7aIYaEl3RPPrrCNX5t+nwynqDxxt0RuuQEsQ657XpLxqKiqtCsB4Q8Vod
Agg0JpzCmfIriAk2bLYiFcO4gGkx+QOGNBRFsrXPBxGwmSwHeKDK6Bx5McnvyfCIMR30ES8+251P
iii8q98Wvh9LLmI/Uw3ZNsnTx2sg1kONwpVOiAAp5NUOo3uUVQ/kzCH9TbWf85xLifga8FGlg2r/
7yp48eHdtyaQGnb9UyNtf+ccrkwkMi9PAwhjjlTNv42CiEZzAMahrkp2PSW9pOcwisqfmWyqmp2Y
xKkfnsDswQFhXiI+D7lKmD1RxUUyEswnQaYAqpjVdM0p9OfExkl8o5MC09IJ/eys1Ffx9T0BJOTE
ynwyISqpcDsvMvfwRv19KdB7/tt+LZj4feVh1WSmo+2FQj+thlhWJvuPG2/BXHEwFYBNW2J6Qpi/
giRmVCwBUFWqTcbagsX+ZL1rAjM8MScklIqaZ+wiTIeW7uXWOWF9w2xGAmrLVR8ZnwpoZrTRzup7
kt73Q4HmYXqeJh28gVNrJ9+7eMWBrHaxRuT0ndKHDasIlpP1FS/ZrM0es+FT91TWBMKbpyi6KDeH
lI90bmp3GWmVPMXH38eeVo1U4YXcSrmILx+IUvApCKjQ1Iy9IpA5bZTdC8FqOcAt54chTN4Qoylw
a3//i5qmy5DL+1CTB9cIjK0S1MvVNHHXpq7h3OqdBUNORMYnYMUAJuiRjeP6Oszc8F+YUQXje7yF
whj0fEa5rpynGdK1IhtDNfwDk4fB6UOy9bMdmZzEmbm/NMMUeni8CmpYUEX9uwW/R9DYj+iqLmQa
IBTnYEPDFNpiiQvP8Ss0amQpLGUWKg2yhaQHilb6kr/Z/KRbfVvIcBLMFodvI9TyhCTMiZ4M0BwN
uOkSg9it1SOWUqZZj7k3XBckI+nPVZwRb/A99RIgRwE+crvu2jx4Qe62nvN8pjRJbtaJkRRFjp4e
t2LIa+g632vjlmsVCctuRRR7OnZvdfgp/vRg8qGOiekBMT8JLFc5uNNDrIVMuUnjMzlcISRhmiPy
yHekU/wrG6PR717Th+muvnwcEoHwij07l7XPTjeW+5WwYB/nfc2Yw+xVuHqARcnPhpevvPJ9ATd9
BsRbcd9gbqwkRw5X98KL+zLm5Ghbq+1Hje5oZMWmFZRBDScSAxsFO5kme+krLvVI4oiRyGIvFCTu
iLgsZfgOd7YQ/KnVawo+Mg+laUiM1T+WcUDh86QgXBWMnUH6/zKON3FZCM9eYceKUjYNa/ztUvIO
b/7Gf+ysjZK38mnjnL9zqngUqhC7X4FfB/SZYYtkZknj3V3VXnotTK+tDVA1+RqRdWPa/yIhIC6Z
XQFxd99ZJaIqs+jv0/RjLCQdn+tqWA5Pni4a84kPemIX4LseWPC4Fd3tijBRjskFDecbkJWW2BBr
wfcz1aPU3p36Jk0nRubK4NpNcy1nUpuHmKZGm7VDNTFq8j9fvPdeZ2DJsSlKFvQx559mYUy5g9DC
cJ18/7Ak+zKh19S37TWrHvS1Ni0FqctI71ZllZZmQNkTMD8dHowZ1frQJ+usxKmz/qLMQcmCZe15
ZqNzYz0CrIAInW4gPqoJdwFbBQ8CfQ6TafpFAovos0UQZfwcDZlFX7PGiXdbFIimrAsU5iDpqSFZ
H99so9kSWjzpArnz4pJHh0bc+v6yK0uxX3zGz9YLzzeZvHo8IZSuTrS20skSakncYD6M7OJFrZNN
iKD2N/aWi8ikJZxzjdTp2E3wZcWep6TwGEfFlxo9I1Xf+vd87pGfbPrsbVXFyWMusmn91+DKYFjF
xTqLCsFZjKxjg39haR/fJF2/AMCYG2OY+A5bc6i9OZRqFV4S6st93SOGbfXHjtDV4cnvZzLP4d+C
g983pH77m51JHMp3sHYkZPZDy8DJ8MIOfp5T8n15NgHjvuWr32Jy7FrEn2pFq6vxqV4lGRJX1LnV
6Rc1035JnUBV6HGviMGcG6Fj94beoKpdWjDfpa6rtylc25RyPLIFOijW/ATKeVcEM2rbnBqhmADI
cY6rFyWDa78Tf/S4ddV/oE7v6UyFOqkdfHqPdGnbB2kzObPj30xz2Te96PR5fH/vK8HpZ54iLi0V
OzxBA7knp2xQJc9AucSAZ8hNNoC1iEByXmhYymfF68Mdr77XtMLm7mqM/uRmo08ghm72ZLb2F30s
68NKKiVySxA9FiUA+KydVa4haW/0/Xj9Im6fypNcyX3zDNvm+mRLdJe+pxKyK4T4XfP/hX1ntDbL
jUyg7SMg7P+aNnsOTx6cPeDFV+vdJoFrQvI/Sh028exDkR8N931vmRs4Fvv/JEOakGTuuubj0iQR
8UGl1VgXxLe0o5Z0lWKbIUl9zWNJm1mNgv9LNUtcNlcTPZfLmj2MlJKiCofOcQjgBzEb70PYBjVR
G6tSr1IpN6Sg/fk78c30NnFfjMbTlU6YTBgkpTVYTEMQ3IVGaUupU3JEJRC9OWHbO1H1eM8dhaN/
Ks7LzFXNZn9S3emDrb0ikCB6Ieopw9oyuLOGXLVn7Foq9tWeZzB2MRJIuzbjKJFIgSIgyotaIxyB
MGWHzaMUvft/YElEmU5hxg9cvspwpaf48FNZ0OWxCy9XH72SX9zugYyqgTYJ+chlVlPhbkeAyCmc
e8cTNmg1GE1if6UbGXh577ej3LaCuQmh0ksYqUtX363MNTkpSOlruP475vQuOH88UXSc5Kj5J6IS
gJOabO1xSa/ITq8kPEAT9M8V7X0qH4OamPi55dOyPNGMB/vjNQuq/rHjjaEFyiZS+jaMZVuS6kWZ
j7vbJ2FlMm5qzWM0StkgHFRzt2TvZoZHz0nqvtE+CLgLfLu7JQeCZLszEt6jfuJE3D82MsaxhafY
B5dNG4i64/kUStMsn+eNLP+dKwHBnEokbnwv8yQQ9JTcNh9CE6+EchfCmOcFzuMTW/hM5MKLLPSm
WKWwOjT2w1yWSmqOM33dTz7V6w/CEMa0tVIGI3EQgVXyo4350uNguJ/UWno1olWOJXvFmT7nzwVV
Iak+rCRAiyCLgDVRE4b+ZxzgIRX+F/CXBch0ND5PgqVChU5VX3KdPuZHiu1HP6AZ0v0PeHHTt00g
Ays1HuPMwx5FBGA/xwxaQDPk9UdLAfClPUbSgjiZGkRWU1mYAxIwevs6vRSd+9sHu0ppOXnz8wmb
7RAG8iJrC6rapNYDrva9gGV3h65ycSbPQ7Z+jts+Q50tzv4N8p3wNJkI6r47BwTQb+nIPE9NZJ/b
1BBJycxCiKYVhphMPJXVgH9RRtMm7Pp3HWF6RCUQ0n3A5zTFNIqe6+rtMNHJIzrvitTKE1tbpT5T
udUCCys/Nt9OxxxOHK28h4IS69RkWSivnpOxQg3t1EpsRJamU3DLXqExlaDhbgGqkfAtbKbZa8Nu
cxLHop18HxAN3mQulaiDcj9DhaugjMbJ/JyK7B9cxvTVG74O4GW3Oi1atlc0hJm5gsm2MzEzpSHA
A9diBGUg3H3bm4dl521HWLlyFDSkErFquwE0+8QQAwGAsYASFdrCITmLfClEcHYnwAjSvRinvxGH
yLLP0WGobGQnDg7iC/3UV4RShvNrkvWEyOlR60/7VCDX9lmQq2FwjRfPUmtYqS/8wvLfZ2SLu6im
tvwihZFeEydloZWmGEge02S9ewKBijjroYltNUbQvJzV7/kHjd6G6Kv1nrIRzh9+SXOOPTYbpDD8
fXzD3PdUBPBiCQTU661Se6O8/zB+Q3c21ZBsHP5DwsPTPd9yKgs/o5pOnJkSiftrKZ6s8NJbBupc
eq7N8OIfhJ4J403GAKcLcbTE4dPtTOWH3w4Hrp27Dr7Xb9injOB90rSERz4q36c6ZHi23iuyW3dZ
DPD6YVVo1mC8v6rUDzm7YZQGwuMYFhqLtn80D5yTxuhSPeDHeIeOr6xapuJIVAd3mfC0M3uPFdj+
uMdbJ4/UbZl+R/lG4O+TSw7x4hw90Qe9T8mpIfetLClFVZXNZnHg24zXIA55QI9sLknCh2Snn7/6
nXO0mjt6zzdyhYwy1DDE2ulR+m4A9AzJaa2zWWhz96wT2pK9f/2r5A933C9gGwkjNgsweFJhEC/r
imwXVIyMhHaTrrGiZiOYMb2S+jvDqrSdFh/y8mF54bsvOm781XzIY1asQRcX43IXlWKn/wmMEi3l
8eu63PoL6S83nKWKokp/MboHQRu7/xjk5RrUaTg9SKdfhYU7MllTgiQhopyvj4aEHVHvN01oxp1p
UVI/z7N7qkRHo+NaYctCZQPLbVWjeJ1CdNBqtKGZqrNC67LookNH4sDEzqEg9FL+zmUP82lYdyXn
IBzxwfOt4dSN4xhpOXG1lQaS5Oibgwf5OT7zxYD9cvYpGcCPQhVqD8iZe9A/dl1amL+XFxf5kdN6
VhJeroFUmvTIO6+oD40270+2rPn9JVxlkZcL6BYJGGziETKP2RVWvWu+pcPqw7FXk+u5XF9ezgAN
4eZogGskBEww8wJ1Vwig+IW3vKP6lBMp5jQCuVx0021Sv2O+1OODo80SOWK3EFGCIf9x7WbriQiI
++/1/jHE92mCUz4mY9nBWdj6JP9S+il489sVvC6egu5St7ArUt+8hfmbPWLrfzgOfY0zGKX7LZs2
SPcJnB8zG4AlJc3jvHT57Pn+3y9RNbI1MGh6G5BXWWYEeIi8aXLieVGD/8I3pDiWFVcOB705qKc1
i09lhE99Ni9uzfo+w1AxMltEc9DMI4ghj/I9nvo0APRM8VC0RaSkPiQU8Vxhq+NAPLV4L6NAr/Vf
VoaWJHsh+fKTPNbZ7BzkL92qsYZxyiyCaJ/ajVvd2RAkyL/5VJUQsG0wmqfLsV5QMsOelBvKT0st
sf0w49f2USoux9QhW1FWpWi4F9RsKuNZheL7ilvfzdSdHu9kGc30Js5SfjGtd/xRE36ylRmM6jwz
OwJklNxQLG1eTAvsiJyNXir1TrpeU/RTdZC77oq9zGDYcpUqxtHmgbqojX1vNthTRMcnuCib13Hb
zUPTZ5cShBYvVBmd8WVUYFSiufrjAtpLGidFuqiF00h6zWQ/oClQ1eFzPDms1zkZIquSPNADNk63
NigJkkMwpieRyzSeym5NwWJNI+w3MTzApGAY8GZJLa26qrGlUpe2KcREJJWSwnT5Ekp0XHdNTZ7z
ToyQG/HES/RDuxssvcy0XtDCJEc8+7BCMtaS7ftkVzevMrexTGBsJzUW3EwRGNhmMryCHvlWuYcz
rgEG78zHW5vyV+jZoeRameeoknVbWcnqqqV4QFLqhk5NjSfNKLbhdkYl5CxQSLvUt0B03N90Qhin
HAye8xYsHxm/1G/2bWfdr+xKBZajuqUCY2vp4sMMSPfy4F2r3d4CbRmuWwSN5M910erZiIR+KWkg
cqvce0f4R7UqLYcLRu8YH0dbtVK4PltdH7JWR1fSLhuqNM9zpje4Sruy+migb1k/xanAdtWrMwRe
nhWH8VQigCeFqUAWKHX/NPp855M4JizYSWegnDwRgQIwa7ums4p7JBBwKh6YGu1NLikDjPPEm9Gv
oKH/aDg/wbd9uX7TIzplZzqQEh/oSJQlILlvIGqzvOexOsEILJS40x4UMThgbs68hfI3gC7kDGyQ
h+2asWdpspoFjQLlBRBr2XUNUBBXxKNzIoJsD4AyIjifV//YiZAScilm8GKQUO/sSHWPBwSCkol0
TkuvQeUijxZVQzlfKMdboDsUTmuB/PHGSbGWZ9uE44NDvnRBm5LcUgCVoyg8bfKjpuG/upQcwIBX
ArntxYnYroIaQrOc7kE46xZCgmbXxoySgUjYRJOI9Fb6K6HNeUy0ylX/k/z2wbh/svCrTSUa4xoB
xpTGqTjc3sfN7wCr1256dT82kBj16K2k78sWI8hZN9Au8mBEK7M5a25gNOi2xhSA8MiMRCRKBoeV
AYykJN4yRSUVrHvv6RYTsiVTyEb7vDyamrRMdPjb+HHuC6s5a2qaTUy4ERmkqfhNEyaP0e0hxfjv
Arxsf7pG9h4ma3BPduP83m53/79raUGd1zS9DanIFeuq6NaUK8XRAcysCH3QE218MJ+ZzSYVZtoT
nEWcOhG3xrSxPUBkmuzT/2GIjrBImykDhDTXTSodRRGimsZmUXZ08BklKe6wIEVuwmdd89C1VIrt
AZtmGUOQM9q/nCid/5an8mpEt9WTy95HcizrfJa0YjgsfYfYzfkMFGyizzAlwUq4Q1+4ccNeeay6
Sn6V3HQP9CQSwxhk6m9A8KSS2drtVlY3psTVc2vklF0gtiag81WnQBqnsaXBL/yqif8foUP/kfAe
oAkFDoSRb8qJF71yJoAjlFPjD0o2Cck9UyJCnBIsB/fmZHaC0XcvNwI7tvgeMqU6TsgNyQ4PUD4O
2du9PmYkCpv9OycseJIhSfDCnAldjR1716y77DwJya943x9uGUL7+Dm+ocgZtfsi32amz25te65V
FcAAtKCr3tSJTTG4BHU9HmydipGdtA+2ml9dqgYpq4+4jrbGbzLOiQpaz6c7ioaOJInPlefMCH7Z
ww2Ur6hn3BaOKUT3IABpjRsyE9yh2Glpu7dTZP3spwnXrPRiZHYI5cxhNrGQeGaVbGFAEriBhLyq
zKrBFEJNcTQWeYwcIsj898LSVSSU1UhWGRfRbf+3N5xOBc7pMmY9JUC5HZo+rRsrnXu3OiAnzq32
RMzpFAJjw+Z9tv6bI0sJ+mqA1ZVgKdlb5yqwnDizFQuRE6gBG3UMb2cqVw/yoWK0fimllTm1Of9j
rrCdi/5TFuHCuC7GcS8Q2D7NA59nyW0ao3/Jw7RAVbYr0PEY79B86hTPBLA94u0OVRpQdbVvbAc3
cyTsIOmBK6ogFEG5Vq2H4vEeRRsE35RSRl5F0vqA51Tn7i701BE0eWoIQf34n8qKBjfcx6pcHMck
58KM/3Pzq57xUfqrvb8dz5ioRdot80besR604BfSq95Z6evSbiU4i6LhWZDAByPsebf+ioRvYOfc
mIu3ExbJSA2BevATOYn91r9YFO4WTnByxHLUuPK2VFaJwMMl5mzeBNyOhI4t9GGaSxSROxaESJA8
I8UBdUsbv/fqA/UYcbE3LOJ6N8rJW7U9MHH56OtVkH+2EgONs5m2yNSbryHodmKBq0ZLajTDiHDe
D1l3hN+go9y3XP4jOGRjMxV/Ig7Y1Z3mIrjelmiHz+sdipUqhJ2s8hfyx2Af8J38+QIciyE+q3EL
BO+e3tas6REGRgmRU8q4c68OysZh+ces3GPosKJljCyVbDKdRS6dt57PjCKWhjmLYUT6hK/3xckG
e11zRQbTjlHZzfJo3WAhJJGmNiCsQonhd8Ixg8IOr/AYJk7Muv+ic8aZdoAj/C26RySMADF+Zg9k
OodFGNiHGDqGnZhYTgKpIGPUcOqwvXhmh9OgWTQ1tFHN8+UNhuoC/OfF/VHk5oJdwAX8Zvdh2nex
h6y224xYbrg31T3gf1obFZrcllX7nS3PBGYoxAmoLTk8VTHcS7/QdPDsqP9fuvh4NjLFgLdNUtwi
JSxVgimnk8eNr2Tgdg5T4VLvsHOvXiEOUk6YzyVWzieiOF5goSqvvCM+hhVCxqh09Np9DDcso1Qa
DP3SFig4wvScIB6dfgNMPfJEutdnFnNM/StgSop62RH1XWWZoCfybaIFEogTr6UNRqRpzBsRR+cg
6JSTTkjS2jr14EwQTerRnrBPwF1TM2F3tNybFg5ENrVpmmHrYIatPqBW0ytmRUb1BaxXy0+cNgRH
yV4UjVtY2I0WThzfBsHbOHDFs6zt48F+TYpqxGmHVQNxl0JxahwnaExcv8KvppOFVpXC236tecfU
VTCjZKz08V9+8tvs0pRTKWsk8OSKEsdv0y+UTPc808zmuYz+C0s5QsnA53mtO90AQPw8c+BGiDJ5
P4wE8Z2257RPZHR9kuMmk0OhaSFG3u29ikpoNBIHRWjxJUIF7GWXgXp6Kim6ykbpbCo0kTgCR8h7
b3xEILnTHgAQ5sLPeMAPtk77MlcVi9Avas7znJBuGTKAHRgZHi3f1U6E4qZ1Oyq9scvp2dZBjAXJ
lyMamY4rxkqq9ykevfhmQCfu+oUd+pS35TnOQY0qhjKdyLUKZsIZ09ajLgVyXHSnx/6j5fKvWkRj
WJcsTFC+PTxsl41YJIb3XNvPfNrKjnHuTAvAHce74H6GdRXWfgt0u/oXgKFfW3yUDH6ZGOsZ39+4
EXteeWjOVzIxgUw4kF4I+HwL5B+tB6o7ui9Lm7mFiYQEr8P1Jw78WH6zVqhseXJ5orOtbzOLl9jD
Go3N4h5iRk56EhOCCoyMDfizW+LBVD8OWLUoEzoxd1dfpUNKUlwrVyNLiqTMmK8X1aMxxhQIpAG3
1YXixiVPxCVMiAs93zHBqWUUsQHIyZHQmw1CNU87Obt1U0Jib6h342R7VUO66Om2R/b7Wj3DLvfa
Ez3AAR7le9HfE1b7sr7XINtp9yZr2wC63ylEaKPdsypE4lBArl/9N7MmiqVOhHtoKiyfR0LNtjOD
hZBAfVfryX6MZIzVcnoAfz2u4jFQQ90FN1mou1zfNBmzmocihx9FvFHHbQIXRs58KOSF5h8CEpab
Syx0/PvR181STOk00dGWAYc2XEqXGGTFua5Vome9mAo1dRuPLcRUO0CUEoebg3uPkg8I+287s+ks
9aiej1c5VuGs5au77cuY+LSY+k2UX5rrTTlU4G+eO3yK4p67xYNPM56x69Ue8kFYLDy7Os+FhXkN
HHD+tvqxeGQF4fOJUA+ozp/ylCPlCF9VPHfS0jF1E7m+6bsushYa/wxM3a5N8aQeRlb+P2cj42K8
w+78s0KhrKn7V1WebuHSCSEMWkQ9BM/xX5j/IKZpkURebbRh6Qq1XV8VecXqNUJghDr/2+sJqG4y
3IEL8TglPXuGmRJ7LVj4nMbdVZyJrg+vdLkJrmRrCtGdmN5or4cdTrG7S/tFQyQgDaNnb4/fFjta
qSAWiQDwEOpJ0Re/K1CD315ZImiR9t2YnOhzEZX2AMCsLBn607gW7t15fA0NVr8bgGey6dXY7ZOB
4MB17wvSrKX5UcQj1+Glk9bznqG7Q5DWlCGEJPvQhezQmX0dP0V/6gFg4zWqkQ2idBxEzDqERoR8
SWFM6Awj6IbmQ+sOePxD+9o2+PA3d3SjFmORZdrgLOitKolPM7Cy1DDyyTh6FkkfhK8yBgJTvQy2
+j2YO79HyuS6o0m0TBQmWSbmCZMDtcvX1j7foABCNVG47oNpUnaGcAnbcKMVqSYLvQ+LiZ2o11fs
yePnIlHnikIRUEkZfQmCd3c5petesU6YZQ99xUggyjkwhFT0g/YDdCjjv87BmKvbpte556YXo83k
q7ft1B3LWM5QXAANFCx4RH3QrcGIu2Hh/Zy2mHbxipInD/XGw5yKoPvTpWtCnhVkiTVizBoiz9gp
SQ6EMQggNToyRuhfDGzY7NN9q9dnu4lpQ/7CiJsk/gkCRfmhauORvLKSGaHV5nDjgPsvXzcpw3gQ
4z948NeKdw5Z3G5qANFXuIfFj/rs3ntF+Jicto4+kFLV0ukdqX3/5Y98JzJdPca6EzfGKvPjtb9L
6zRJbexURT3nZBtvQLt4DsENasVRHYpGP9AvFOkYlPyKe1RdxZZOKpiZ5oPgbHDHvhNAwqDwFqzJ
B8k/r+4VAL5yE7Ix/RX0xoo7iOVI7YAevY72rCEkZS7g1b4ImafzxGd1mKGE+BURMjOJUa+xzoxT
Hj+UaCLgpA8LuArB8Lin+znW5sicz/eNWuD6YLVLS1zVq+tdBJOMSYrM3rYXoulQFbrOFEdEEUw+
8aHDkL5Ox7t+1friOHCdZMToHsL4yza0Q8htAgQookuN+aLhfoYgLL3dfcU7Br0BsBmP0/zotK0e
Mr0iM3kW2LwMM+8GDDMg3/t2YlOhLlvpjAD36Zbo63YEBMtfouFL8qlFvErpE78kDu9+8BaRj9Te
Q3meLX+JsEJz3LiNS/L7vjLIwt2RIT2+HmSWiEMegk+X4lWt9kxVgP38Gi/qAH8KFkXCkRigX9ju
zkSG9qblpC249U8WRHjyWzGB02hFHuCDvtvb1epieAbgrM1x10WLgsLnWfxCnCm7eAWc9YsFPYAU
dkeVHgrUexHUr2u3v2Md45G0iTPGnA0PRHR8sE19EK9Gt6gVM6a5X27nTCZMSApbIWbgPZ7KEkHz
kAuZB1dKg3qy6EVSnFH2TYFz34+6FzKHJG2O+3fyL8X03eUfCBeG9iu3T1fxVxRaF/Gn/YsRV3+/
CGFbEhyeqtKTI+hCB6JN2eZG9mjCI2Y/XErCf8XBKsINWgF5QqPY/CurE96rAx4fncpLRswD8Ish
CZZzhV6ihjVBig+tU4SejS11buqoT9gOahknlo6+dBx4vDFL1c8I/FzBAcMa10hNuwXVeHV+9a+8
q4KbM5Bs5kUM2FtqOSkgPVyIQOhMply/7yhtVfLKm7nq20J91mGQdMd1OichPYJHiPiCJi1NcG0T
UMNQpUmUp2CPxJoqbC9t9AHSZMQFR4k9oJuwg9MgmqWAFXfmHrrZ/9cBst6htDNelVkLnMIwNCVM
2pM0N3EA+xBzdR2lg0c7Smyd90+/DWbYj471HHA9Sqm0xmunXJW8oAELDfAtispDNu9ZNxxGcAUg
4javt5oEfbom73k+lCD1nsXlVJHecPFLx+jLneUMj0ftocIR8GSuP5YqJo6KZXIR/RLPGftSwhK1
+dnIbXUZdZwCu/wKW5uZBPxJcEc2zePJLB1DdjzBPPMMAmhz9eb5sOaN/mgWAXJOAvZIII+yC21m
/97KYYepxLjyyLaEcGWNej1pe8eQXCtXbMh2cREMW4EBfHB8tgTid0pAmIJCc4HrwACnVDjEvSGK
X6v+TUwcYWB5hK1GBhp6Nqr5BbuB2M/S7EcFaC5FzYOhYKUsoLL/b6mK+t5UTW7rFrtufUxWj7Re
Nw42/9zmX4SpaM+DSXq0A8A8QnsPIi0cEcu3ZzFmQDCXbRP+BoDvoB3v4IS0rD5i2Bm8/QWioa7h
EHyGUZpkY3fF7NcxzL/sjOtiQxIHNYGbp52xxnzubgAcwAPhMEWRjbEOVpQBcRdnF8XyeliwxE3x
7xUni4OUn2aa1wYuHnXnVBbSrat2aTx6JYsclGTlcT10jR72j55Um7S8Ox9dslGr79rfV6NnRH6W
NK5TN/6xuQuls7irfiqmIwwaZTufGdbmW/TWTMLT/LqB+/lxRTImtF7fH6v1K856h2jGZkO3lH/n
i+b/bOlKiwThL0V5TdZuuY/0UKf2JJ2tCgd1+bo3/mnFqJZXMw2Xe2sxE7ktwxocfaZS8PlEAXTG
nsy4tNb2fSSt8hGu0COOY4l4traipQPuHVA3nIQcS6la5kI8Tj5Kul5TFus6OsxSN8J+3agTcaGv
Su7fiaxc6OJ7SQrQ53j3GF2w7vj2SfCuxPmQzaFlgX22wZIr9JB4MCUqMd/NDtF1nccSwoTp/w+m
h+GH7dCT0iG416d5K+aK2A980RF0LDTafaG0unDxEF90e58Vv4lqaHgfSoAaXOWXBTanFj+eJq5t
dxg/X7Gxi0DZOAxyzFd/Q7fguGIqyy2Zw93YN1xS9g9u6UPPcopNLof2N96ImU0ugWUL/83r+cLU
NHYD/1uIU7Ai2W9JU6MUgN3OKaRLGz8YDvKKkWIeXXRQSZeib+/oeMvMZEqOvM9cOkfH2Z1fvpcd
KszDl6HBQknMgmVIzyDwU7q7bu5qvI45RLx4KGik7xepJTdZwwdtIDymykuC2EfERoz8n3pQa6WH
/4MeIjwcHfYtSpgh8x9ANatwrzT/s5A7mVZcyUVoR2qGUwedRSQLpakabxwYjh1KQ5LCc+TfL5oi
Hy+hvvTCk2nBp0rtfQ+RNLrgw1LolMYbLF7zqgvGg98hbsGSjFJ7qJPX4RaDmGG/Ru1XlTil/f1y
YgvZDH29OSawoMit+XEBQkT1vIW32zoHmbKVsKK2BJZkULv3P9NOeXK7yvVWYv/AYHsysC1O/QqP
XJihhpp6bXEyOQcAzr5n18jCrGHgeuX3z2HKbpn/dFSIfYt6XBrCYauBhmPEETFfXZc2NujooVhm
8ocYPBWWY9nzX9j30+7WONMdWXEyrZCTyWtRzQRjxlbYVP4sD7RteSj9gknE/Mq8RSWR2nQnoqZf
yjwYUtgJdlWj8Y6Sz9e6vCtHU7YpTE0whUyrYNlc7OD7jvXBqPC+T6blfXdbBBkR0K49anNfNMSn
ZigEsuYYEs4m3X430iLCK2x6/Tw6Z7CVk++7Iyq/W2s9nQPSP/j1lANE70QUaM2GFxRHOu6Qfu62
n+AW/ERfxfP6Vji8eJaWcu5WZ8YmN4vU08tVSqLQ+WRUeCuA5UuauvvIi+FqiCPe/0YQ2zX9fsgV
0W9YgK3hap2R2VLq2xZrOXMLD7J7Dfv0f2RBKchAgraxu1aoQsv7uboOMnsNU7wio2QkjVzSAUXI
uW5KTwAYsryxGVG+zca7DP/QqHJ33PTxyhyeNkfSplCmO8YF3OPbxLgQwLIIefIW2GNelEGPwUtp
izVNds0dkynIZdLHlOui2NK6I1jBWXLPkwbNN8hkUqLNMtMlPXdWGH2KGEe4bZuNBugZ9IxEFRdo
2Nb5NcHlW51s1xLGhdfq/qfdXQWgobFJEkDCeXfhaZ4hQV53wltY2LXBhwk0mA/aIKlhqIU1ftZ+
bbsnHDLtTx1iyKYejAhwO7fzV+3Zq1pf55RnMLiCOw/nzaLyYBbzol9icLXJSWHpZ6EO1+NniqQC
+Jo6Ftg76Qt+PoYNI8GrhuIeP4d0Wb0dAQEwnL39NvuxssuNx3ugc3oWQ/4Vk81qy+Y+8wCfWoXg
Mg5BRbhCLD6oLd13lG8u9+DzaFGDC1SytMMy1RF8OtNX+X9U21b2jkzLp5c/15SZexK7l97+DfRF
NrqGtjlR/gxFZrOjZKd6DlcipaOWLOF+IQ1V52zFMCpKbDWUb9fPol35UyHwrKLZ9lWi6Y6mtT/e
wk3WbdLr6cuk1ncfeZSInFXxqhdmNKDZZ0xYvgIPzxBy7ItSHj5aXg2mTdqfIASzsoYinLsGuSda
XQC+36KOsPS4njCcd0OWFSA2K9ZpdkZDSCJUYefYtMstkZTxFbwWRANFmGzLY0eGc8gSJ7xvVgbD
MEAa7B57kHUNpWU5RwxDuQCZdZ0E9muMl4FhjIlJutfrUqxTxi7OryFxuss1Jzy2qhEhNbKvJSB0
xfxs/5eYugUIlxjFEzL7tzw8okEWLDZZq4MZYEkCYVy+W81IXJkm/VCuIAfa6oDgXq2UNbj8VqcY
RdvjwcDzhNcTIUe3aaGon5AY4/N0ONGKoOSCcDYdeHWTxL/ZbCNvNqJpHjUSBuHxz+/HYRDkVX2x
z2NF33/iyXBHqkWLUESysNpcp7I0T4omjpOl9Fr1/oJ84Dw6WnoXi79xpqSRUQc5pHodhIiZpkWF
a3uNVJOPVF0tkCHSlkpYVTt67ADsCHLu7uYDYElvZ/cMA4WVD76gbVpVEjeb2KTeLiflBFnCKrK0
DTxrKifI2M1eh3LUzw0YTZBv5w5pBmOyR21f86+5FSK/X8iWsyN88wvg6fp1LJTyIa7TpxVoyYgp
XEoOgcE5VARis9W2p1Zd/VWkYSzwYiKADQShPPBw2j7+8720BZVWdV01DKBJliiw5XdWvRYX7B+u
oyB9JhCnfxieUMpF6axLo2MoGjTWUDwAdksN4Kdrrbd5NJXZrueaBQdFOYt1uirnY3BeBnMgNFs1
3+k/R63nq7BSIQ/ul8iTgfILnZTmOxRrXMDtX8WDssuOrh+LJSxEaSIy4v9C+D4Fy/9mCc8Q3zPi
Qyw5gENaLjXh45ZBmgRbCoFv9I12G8jcIsUjFFcdMpbZRNaMwfqfq4wBCUFgqR+cdo8wzA1lcDbA
vAVGkLItxDptfKrvcTgoSWk7cwzek3tkB/VBYtGa0hxayqq9Y93kjoakbZKH7BBp2YCLNZgWBejp
43OfrvJGA+gkBIfPGmD1Z3Z9Fz49hF9xXIdWclSy26x8NnN+P1fLNnxRtI2ICdwXxS8W9/q+CSYn
AHSd70Y60stKg8nK3zSoBh3o9dNlG0mSUiktm+V6RuF3VYQxxzd14fjJ8IUJmNMQ3I796Ptnsm6s
1s0kx3ZvVwO8FBOe4VKvdLnlSWR4YYe28bI/Hdn/mxQyRBRGL0NgPg3Va6vtRJ+SQHdoXTfvyZ3+
R5st5Gg2HIKNx9uCiNZDl+DuuwhR8QVPH9tr/XFvR0BI4GlwFt2/BQoH9ga9R8tRFAHkGgTb4b7c
jlnwmWjenR89KrAU1jf6jL0zNfOE2T9voo3KzddKWoZqIrjHa7TqbtzMPTSm5HdZ8+YejtYkQlGp
u9F9gakhBGjm0QJ3Fu11EchVygppd5HCkWFDsl8ogo8ZqOC23iwhS2pG+bXuVKcQG5dqmupEA4Rp
vXhUVPDIDrM6Mgt8EVGSpw/0UVDgCOD1rDs89ubbmd7ahB86rLdPcCLMCTP9anZ/cOxHJnnb2fIg
w4v1ORQCp+Dh6km6x8XYr1PkROM40a8J8olYJM4NW6GRvkSMlriAQSuFJB2hJs/E3G69jCqo/c2+
SZgQGKiY1CB6CH/nRtXYiHaeIZ/UXCh9nWjOFnerUsutdS0Kd1Wo7drgELo5vXU120e3c4WIk9Tz
RtTjjnpWmefS6Hd0dUZWludHppzwpwETwSet6aw5XwujUCPVyr4pgMAXte8OigKGHYFtxbnCczGS
gVME+pQHpf4F9jS0PfxUpm3P2drhXWNa88h9ZzI2lqL2QQwSD9SMm/LEcm+Rbh116SSXePHo8qd6
ohRDYWErSKrQVbcFJAx1e8t7qChuWK7rM5GEjS/faw1Y683ICVx4KoGKMWZP2jdVVXNhwX+O1NVI
5NK5LAEMSm4q3UUEUfnC9lP5aZuE23exxDwYJig4Le0oyr2khSbNc4WVpZaqzsedE/GVP/HjXrRu
NaBwmzmqn1kCA5iQk/fSq4l8JxBXY2n8llgBvLACIvPBidAxouWRuAcoHhzbmix7DAl/v9v5tsXo
z8bp4iDSvUqI9Xoo/7LZYm6QxYrLpI8UqMzAZclV75f2d0H8cnDi6wVC3smBGisOEbapFRcvFYju
w/oOWHtUiTpO/Ck6byuoZIsfh7DRNYz3Eo+qi2ouJD6+uvy2dWposOhf0Rq08SieJJMDOChs9iJJ
JDY7lXI+5wiiEz/PI1sZke+apZ6ntfL9f5yf12T207DdJl/3OVz953xWUmX4yvWBJnf7iDLLsvMw
Oq+Ft5qe/2e7CDeNNp9/hE9F1ddI+RAB3DOWM/OD3OsHk8ZcX1z2KQA/PuE6iyfHmn09yrJnAfCh
iT7psFo5tue0aiEjvpV/gNS2a594QoNFhYYiJOdb+gbvuJdzvUnY/zMTyYIG4rbk9ctiFs3j9xNA
UNV76XmxZjEMwrfX/qiPTsgEaxCFNGFF4nm75LDf2JKrwHD6hZaxBDGM+XAukmP9iAwY8pBn6hKr
7H3eNBFMMuZR9a5JL9snbepQORYDDotcJZFTAH81DcFe49w7WMUv0oMkBzDV2jZRx2XNJLB/zVFd
+M2jiz9n6v4Qkjc33xMPx3zQ0/32Ew1VSWf1AfER+hYXCK+6ISUGQFO5bV/hgIDl2y3XmZwquaPU
7wPRIDtPRJqDKckNNRl5go1HUAIPKY9p+4VBsZflLr9Lm8q/eLlwir7tnOETzdHeH29NFkJuJ08A
UaughivumrzYbHt8Y2bAzALMr5Mp+xTkw6HCOLmGS8rCT2GLZmWvbNU9WvFp30v6qM9/hAHfIf9E
0bQNWCG7ocwPrip8V5Bik7hKnc/USVnnVOwTHj23iWIqU+adHujr2w6V6bf7j4Ag3tXbqaxOmMp2
RZ2MZztnK9NE2iPK+8egnj+6JVdNSdNRpUoQ53gw8AZk6GpIdzJpWt3Rj+9qPC/Z/SgskxWRuXUU
mKjYB7lm0kFSxu+2hshqtf77o8p2dFGctoihl/UeWkcRfxMRbmv3K0JoLcli/Qt5lJak9Momv0x4
Hb1cAwnnbzt8JSHT4qQGsc0zX5X3K6BXliJaBCH43TDprUAhAdSznrw8u0xKOGyAadyXUpwTn9kS
+Hx6RGthp1YFzd+okmob7P3GCawSslQlhmHpwX0POv3n5QskhaMp6sXdbQMhdSzXn0kKw/RwHq19
ZkWlmNNunH1apmrUAyd8MsA1k5B8GIwSinOuhh2Em44p3b1K7kFpIZvFjyL48RmyHh0VMFdSJYIK
kHA+W+AcjD/TSg3/a7yVa4498kLZliKIdfp7Hlkq77jZ0fSI5JY9dJ1rJ6H2XYfVM3rPTpRBXBDQ
PhYfKI9UUOaSWZzITy+o+SVl3TAEmtfWJkaxz7R6YCuHml6kt+S/f8OPCDM+mqp6ZUYapKHS+i+w
Zq+wP2CE4Mbs2g0GqwhdDWxKu316nHm5RizmC4kRDO96nZ+jTPumJT/Qo71AcBaT1Uo6asShWKLm
/wfYRGPuU+Dx4PNoK5ijsU7jkJCWxtWbQfnHf/mlwx6mAFt7fHdzfFL/Zeui7QyTYoFZta6y3fqJ
GBwRENjbrG/iB4x6oDPHRhx0JjTnxyYvLsmm1Kbse3IQnOu1gRoE6188g68DdFSCexSE/aV8+FHI
kWnpaQArygCNTA7pQE6G52RsyP6+hxPvOsrqzS+jNcRRyZdKXG/JJI83sNOuMF7R1EHzq1kjroEJ
v/Xp9UCFomlkjxgFLXocuVhJZnF+6Azm8Fvp/KkguJzZ5mCN1iUOiyDDuy85iyfN7bZtmdoSax2L
l57FHguECXC1IJutkiEOFQdLR5KC0Jhfpbf+2qFXbr8418Dk/uwyo7MLp9ezAmwUKmP7E6et5dGf
BwM0/upbU4Mxt59MTkjppLyQkdF34HIw85fC6sCQLaodMLWbTbGDCeTIesAqoXtZY+oCz8iJyype
UadM6Aoz9iqDTXuQkFPub38JreXadBHvBO06gOoMHkbRsXd6xfUH+lNmiPbV0xChIbqu1JtLEfyl
UoQdYwIjaW82c2OC6LgD3oPEx0vgE15Lg8XygNykCttdtlYG0mScDkPJkaFElUbw/rDTjFD2fLdd
FbzUtI7CJLHVay7huHaiLzCiIyEqeY/yea5lM4o7AbLE15zf+HCEONsiOV5hoChf0+aI4vbPqfz/
ysW7Qco+i16jnMD1awtCSo5rO0pTIZi0unjjkwcFfoxJDcSVdMZBlDK8OGCA+8vmRL696nAJO758
dUqee3mOCiXxB2c8rsYkejhoEkko5o7MUFY23pXNcj5Litmu9mGl55+7KIXLplDp4RkoIACh3Y/6
+p6WB93ynUDg14vvfimo1UwxcaT8LSMS8HLnvWUg6ZLM7vzp+R0fTeMQgAJBY5GFDJwUTEIoFqmi
lwDI6uHiZN4eBYho7X+KLxCoSgRfFupeEOuTjUZU5sMJvKHzd6LqQ44r2C1B2lM4PVXLrT90X0zo
v3E+rnIc6fOCmD0KM4Z9xLyqSWEVeIiKFrLmiZ/TkkXtKDw7SLSuouO4stGUGXHzSSwuhcab+Tcf
FYtwYS6I2wN0MQGqKLQkBpKfwzw3qWaKFB9vkc6mNe8b+ub6A7JTaaWg2Jx+rh1FPudI22kaZd2J
wv5Zh3LlrwoRbB6pvMPClRkLPsYu1dSkVnDzd6kQ4cb6az3t5xyc5jtr8EjbclMu5ow1OyeYthr4
b7GQ+G5ioj7P3K0t6pF41Th+zmTFEgvqpuJo5AbtmCj4sPUQdLeW4bUGk+LZwzLPV32Dk2r782q/
BnVibHieSgnO3j0qePULFYGY6I76YfpmPF0KmVXY0UDfEUwjMVXUBv50FHStvCPZWaBDjtoZrwFk
1Yc4I3+hvrk2Xsj3bwjox2PDCzV0EjKkwkZAMo6MrUa6QxE4W033dluP+OttNr1rAa3HVoNLnpcw
3EyXRUpM4B/YZ6i0Kw2a/mWhYPHCRJUGE2htb9e2srAGqjpYm+2q1RaeEaOpbDQoBsjuuiVIOmwy
VP9zsYVl4D023eTURoWDgmmGmEgS4kxjKoK0TZMm7dUvnkefajyKKYzEa2Lyfs3+CRO/CvSGz438
XQj23P3wB8VLfDGxr6aq4gUiM6UPtJKuI/3kBVWZXM4mpRaU7hYXsV2fXMMFAXlBbiIykhXaCkWd
2HBnrC7MGuWstaGSbj95QN4QrruywTFn1fjYU1RciTi5dxzk0yaJuAi8MUJyF+IvyxYiIMG805Ff
tfPggkBA866fXw3nwxPAyUs2HpVANuTTg3qBSI/Z6s3u5CDa6DAzioBQ7vZ5kReJ7Ra0UCxLSozm
EDAoOmYc/2ruMBZs29eyvbqICYldU3hcW4HUWjAb6FDHNzmBmcXweU/zFp1AIbeV48xk7X8+XRWw
zogBnybGzawiGYtZMWxj9LwlxoTcXZM1bcFeJ2I2r6Gvufg+dfzUObsWXnqhvupJKxjRyG3MAp9Z
IzwXIeO7XD5oZ0ldaWJ6ydzRXfeNBfLb3mXerFKzI60eBGQr5FiAi3LA0B7DjDzyfiVRU6MtjoHG
7KBFMcB5LwsIg0cHlGmfeBIcKGIBSTm2oWo7MRASaa5tFLdA/ia/2PZ1xCU1t3+2RiiDJF/m+6mG
XehFrTpJKqb31rnN2YlhTYOdNKFlcM/fQ2KcWMPancWvQdAYmbVgYlDNOJthhL29MLv1GFWhl60a
ZEP0GrjCkJX6oRfxPgtl5ynH/2es2zswknhSdeTTWarbb1459PDPyfcZ4tmzGHvGbWHSKwMNyiXy
sVwOYzKfepH6SkzTubPG7o8gMgSC2hkMx+ZaTq2LsvCl7t3eMXu70jHoNAiNhNgEAEIjOPy1WZpo
zGCOmuAMkMQN+Gf+ZhXx8EZoPZZ8fmk109n3k+GioC+0cnMoqdrdXSPILt49s/HfL4gRAfe7awvu
Gk3c55RS+Lv7h5xfIPcK8zmo13lv09d3j+/pUizh0yV6DRObfYFSaqvNCJcLksydCESRKh5nyqAs
C7NiubSHxfq+auEulTAuCAvKBHbtmKTeboJzmWg1FRp6T+BG4T12qvGxTtjExp5GRfIeXOHSiBMj
cEsNo92nBkBdsmnRK0qOkmlGgoeg8rVNeLUEAHeBVm39KDfwEY0xo5PSi3AhsHVB45hNRTZ+myM5
fjYV4Np9gDWVGWyedgm1wAbYePSFg08pQb8pv9Jsgbf174i0D1ykDiTwOw4efrrWuIw8BlyHXRDQ
gxBpXhBYGtK6phjbrKptzVcQhYI+biO3ZaMdwXrgIBxsjB8qItWvQflb69NeBCOMM9PaRc8neXzR
6Ud8/6d7PWT+owQ3WTvULXeBp9NF9tabBylmXdYphk16oCkHrKEYMZuNghYfzunP3k1aLYkrWiFx
vPcUxPuQdxvRhHK2VowIU5uTtCHaifzH+dzDnhBi0bkHvFyUeFnruFUk79ke56Ms6qjF99WHXohr
dA+XUanpcThMaTkm3WbAjj8jNWPKB6tR4AhHo3HXcOBZha34b3wxHa3O1yZoB+eO37QEgS3RhNHC
G5d65mT1as35cXTzctYkpY0AHbjwyMA317X3o/rw5DZI40IxTIu7n+CBFUwYNlLiSN0NaSb9pGEw
6QSHHXutSQWmrSt8gDtvYxr5BWcyNEeu9nPqhIUrFXgbawRfQiJ7GPW5j1S2dy5bAyoKpInKT+43
v7w9rj3a5zjg9I3h7pBDRv+XS+qMmb18BCErdFI3mpaRMhGXm2pKmGLQ2im+UrWGeU3ThoxXvZhN
iN9yqz9yEoRdF/3DSFcdpYVqzTTI4kuBfHCPSFFQhn84vquPccEbqYmowMUObK/q7czNXYC6gY2J
4SsQ9RlWxVla+HJiI1sNeiQPL4UK4syNINhw1uPNo+0UrFUUPoMKBJl0vHXSFiJgwnTpd0v5fceJ
oRDqpK2WnpXIoFRQyn1UcbEqQyEF7jUMk1u7DXKqpkODOLqL3K2ETiq2kznQGxkT2bm00+Yr/3Wd
nS3nOG55vkb/3d3qqZZYZ1G56SA3KbFmf5Tx2n9A7JaJzbtlfl7CqJ3txC/4JK33/h2OjLZR/Cbc
jLeBEtO0vGWwYqUaml41qUtTbHYSRKsxM8QwZywdoCZvW7VetAB5OOARL9SuIlU+1bcADNvD2sl8
y6lWMh98mSIHGpMCL42vwFdTs6bb41nKcu3t22NY3lw1fEMLjqJNG3x0sVSyVp/OwqP3zyDyHw6T
84TTFz39OwgqedvFn1c6IFhn8pgyI+bucELWeTIVgesuVsStAAVFH3oJhDrLtqRwns7WsnaQk/Pi
oY4ePtHGrf5rmswdC+jCmqIAsbRSvtdTJBLTJ8nKtFoL9+dZpty57nxDQgt4W2k9yuVr6UQklaLI
mrjAAkibwb4ZpN2l0M9nZY62KBYrOI0Jx11zNGUxxbVrKLQWEV/gSh8oUox8c7dABEi9NhwD2Qer
MddUG2b1xAhmjM2cBxxPdm13JySSyAE/Xd1jHHzV+wAZnXBE1dYOFB6nqfa+R01YQ0uOusQGcUxc
0PkkFCVm2r0HbN7z5rC6OhsPNG/BI62MrD7NbSN2x3wcoK2cmk5Dy7UBsDFPHlP0R3/07SsYyxMh
/bAGopEVqSIv+Y3zQp19Z4jHV71E6A66+aSMl0QH0dQPa7iZg6rSgTt4fLcJRdhbHFTksHroz6Cb
Fd8WsRvdcO7oKGNjtWdAhw6dCvgsIy4udHxYCqLZXtKP24sc8UklE47wDs7dPxSgB7JCslrqy28r
bM6bXT/uDv9a01BWnrtPRck9nai4CmpnDL0DnjDc2IkdUzgfGP/uxOpIsaADBiKvhaFjK5hNjSYu
wRBXwJCenW5vzCpFE95StiPNgXYdYckN9Z1UipOPElRQXWZz/20kLnLDVzsA4tEJw4XnY2MAJSf+
3o+IWS8E0E+v/OdYBmeZikCtKFUzfovwMTTIH6ej9lEc8J40KjizyVzp9AAsxy2tH0uv1HpVkXo/
KQ+HHdNjLZVVaNRMVVC30qxU2gBcSrl0zmdtmm0Slg2dPoP1rqvgRUq9Dj5Q68PD9uFLqXyHDdPL
GfvF1tNzv/OBLuiJFGk/jp++8h+t3RI/moSMlWDCkgnngcLiT+PQpeyvK8OxgGi8dfeY/g1ho7P6
ou5YRm+FYL9vDGKh21tiPOm/ubzc+EGJXbFfhDnAA6yJ+VPCxN1hlJH9WFuv1vRsRM45RTIJ3eH/
iDXy3xcpCwRGxfEOsWD0eDf2gj6C1a8VpguwsOiY/GmLen3F6gSwFqvfnoXWvAB7xmqk2jjCvTSC
aLKuYQLuSTZKJA6haUVFeMEcD97Drj5zUj411mwkRHkO3OwYtzzR8t8eDMW/PIMn4zwr8aO+7PZ5
EIaott6Ork1oRx4m0Bu8yl4RkcqAhmO1fqVdnkmaRRRuI4NDcDkdWFOWKTZrEz4Gwp06ytoiXB3E
TWqlLM3EqT1n3jN1/sDPMU4BFUoaN8/A/h32lJb25Uk0CC3HCqBcfjtr+EoylInWSoqibFMiy0ye
0dXQT1BNTXD7jimXzaN0PDasoqrpfoucLKXA2dzxrSzWaMijvN13+SPOmBVFR/zCWj/jkzx/Y/Uw
WUcT7sIKQn/VzlLtJyFoMGoWa8NsOSEYdFzkvVgeyR9W+hAYrLGb89lYASSBlaU0owgTXU6iWZ0Z
kJn3bgUtdlFn2QHThJvp47tODxZtEK1YXpI0YHPSRxJEj9cOOOw5aR4/rzBdd4D81WhkqYhnzcQ+
kGksziRAlQWcqUvJdDL1qHpg9TVMU4GSkTnBbdN0fjZGsDqLWNmr1wwDKcj8UH4pEUEsBXrqNOAc
Fc9bgyngS7N8fibmfb7BnIPQKLMvBQvQbnPatLNECNbpZzmmxp1bqUApITIvENIXL06bzYDjiiEI
oFsNwZn4iF0KSk81yPXVtD59lmKG5O+aTNKiNjPP4uq1C5/KGHy5R6ZBuqg439VlQBx+ri81AeU5
GY3q5YXX2dBLf0Er74y2lZBpOdH70TgDLOCSFzXMlGZ7PdOIjm2HQI0nONL/nf8RpeUxBKH1Wn1V
zbsJnMWRjddVBjJwQPSYlZ0J/I4oSzGKdK7tPcA1FOld45bLPda5QzjQEtTKNTVfDUFTDjauuQ5V
EZrmeUxbsYyYV13N5N/PNProIwpToysGaILHvfn0KPYkNQwpXSjZL3wZ3yvD0K+2qM70OH1LGzVc
aOhgw6PZNzY2o3GNRFdkL+9QRoRRtVaPCrpBNW9SYr2A5PDkshkdhhsVdCx/ujhCxQQwvriRmchj
3yazPAALCK72TB6R2tyqsbEUbMfo9yKkqnHLOEXI+XUA4iUxUI9LzFB/51onMfVJ9erqV91hDNSa
M3haQBstExI5ymxOjNKK51tZDNBIUuLBBTX+V18H5zs/lTcxLokvdFfv2rE/8+2av3Y1YSqfTmhb
8+dn0tNdlHiTsukFxrISg0XPjDirs710zPHKQZz/EgSwEVbwltUm9i7lDpGu4cEoLqmaNYbQWKMh
1uSl5bd0enu+/iLpdy2/qdvcUnV4blYWJi9qjNjpTm+etjvICEvFjsd0SpKCkjePN0pqqDXJBSyn
68NTtnHHdDxZH0RhsO7wETM+Jvl3f8iGNvlrz0RszCkaQ9983qnpeYiCqj8OdBox2YIjS34bClZC
UUfvKXDIcWELLd2sDv2IoTmC9LyuAPZd6u+olGLcoRlSY4vuqY3IrSbLgNHyHhSGmK0qwhT6Wr2D
tlRefPjRxL4C3JwPoqVxJxEFnIcFVc3jXeHSbumekpmxpYuq462PbNJgcqeTkHs47Gwd+CP/Ziqd
aiEdzneqpUQDTI2rgzTi0GRaiwG8Ga97aW2UuHE9wWjCi3caAzMZm9RG99CE+okHaXZa53BJlJlz
+VWNjLmQuGxavQf0z8xmujDePj4Ciuaf1KplRay1jG1eWcDSbcgwyn/gkounfZigXUIHMEbODl0+
rqGAHpr9eNhfZA+Pan+Wu79ys4wiSJmko47wyUEVvbTzYL46p98JG6CrfMnpUyR9PNUTEcaRy8r8
0m1Llj4kJrv1w5HwWkeUwq6Vb9i/mlfhGa7JQ8dpe8W4MVHpy8ZsjwJr89UEbFEVO99hU6LK9lGy
HkolYzyTLPkI67vQM5zCphTaiSIz3FxSysLv5PS8GfbUjeuCe9HKQEDmoaWwKpJYbXZfIg/ixNpM
RVYDMxn8sqyuvSu2B+6wdQ8lTOw35AErdruhG3k0iy62vg++8y2dKHZ3kI/6VRG5mSEUBx1yPAFz
WApk85XeuvR5uJyfXrRC0bSC/JljSWDj9LNcVUQDgWR9waEXgGgzzlOAHstTu6+sdANcJgv+ifHq
kkV7/sP4g1FZDdlP78VkcyHITLA3yXzgWyJwzOVgekQPOEcqm/ddZjBRqBxY/B7hhcPMnwGPiCfS
fHbHAO9V/37HVf3wSqD3hN/JVNgKeTokHXA7xpCCsiTE+DrxSPOy8Qyn83knC2JENEF1J8OcfS+6
izqiOCgQ7rwA94yPUn19PzSXdauff7zlVW2R0kOgYKOSe4fSiotGqCpPOZriWOr0Yj42WlU2Mg5T
Dz0efkp6mT8o9/nk6gQcQm2K4BfA5i+fUeA7NnM5bOevMUWllWK5PzfmE5XAwX+0emtatJH37iik
ZRFL+Oi3MqbI1miFkAcapxsgqvbIa1bWJmik70n2lloxyUWQPJojxLAEWnkiUGSM3eC6bppCsCUj
nvgih4q+eqZTb5nRXQdt+DscXVhH9SSNVRK79oVwA1ejvSeI7Soeby7jDPmIPX6lhqDVf8Rrn62J
FakuZgVSNFNOVPtxh1NLtOJS6YCVvpWmaOsAY0/ADk1RPq8HqaqaWg8O9TpeWwiaE3eepyrKeIfc
TYhSy5WZ5qvghRhtI4eOCoAQNwN1ARXTEt9U9jZTVS9l0uBj1S88BAeT3tLg3sZEZXD+HCFrAW06
buvjSdFcNkPZGjDPeuDDs82u/10ZdxCpxmzx9I5OX9nxMmCM4HKKRe/34SeWZDfvl8bakOI7+hY8
1E4t/fq0yZH+Ah3BcGk3fmalzmMDf2+wfuI2ocvN+kH1/6mFsjNbdFlFV+uhrlPKFByeDPXeMYKy
MpIyzFmjmRf0rpKEW/tb4RpOs6mHnIHvdQ41ABRh+l3VBsFWCt1PFRJE1KPWumwqen/1Dh4p2QkG
A1EkQYtN681cNXRT5WHvso8Tu0+B3qfoaaRHDVL176K4cM2c7sM4u9GNABvEcQaUa1I5M/5ZUnty
+ueAhz5jdPYSHJIfynCXYrULQ4rzvNs2aSvR3e3VOY+MAkdWG0nJygQQVgQ4wLq5j8mqa4zBBVdP
1kelZGDT21fFhLwUIFOR2JM7vORGWGsPSA25CZbRJvufgH+99+T+Il8giUhWllVj0M1Bn13QR0tt
tpU1l63+0be6BL7fJ7FntW9IyKwP4TdMLQsYkFg663aXmwYmFVqmkz/4dB4m/anfHtNHhFyoxRPw
F3o+LcdL1P5bQg6Up9xjOS/WaiGieqlh9Pt4JXiV+LlCpmQOqWOC7TYGcTUe2RJiIHc6bP0i+SbJ
HefBUNneZ2Z8LFAq73mqkD3jEFvYs/AHUncq4gK7Dz0wbIDQT/feUSHNgSFjY2p0lEQ8xWBKRyTa
tylzPcNaVeUgEl+4Dc5JcB2tCLhNcKMo651b3oXoBZQ1mb/lwxJc+oNTkmOh1Xx2hi/wlVDS3I+j
0N0tzAmiojQf6HsxBUg15cMRkRY30c6Ff+jUnTDxiKA92oKgPlLOkxj1TwDJ40MpOuytd9hiQc5t
vCkfLbEP/HaXAs5gPTcqtIEgCP+yqF9LET4vZpzL8d0erZup+6UiK3S4XzGQAx/SsMPz53HUSJK3
eVeOeDc3TJ/mvRJ899X6M59hqviM9XCaGk7fuJ5W7q9pGCqCqVivC/vHF2EJrOA/tvIBFWIoRNvE
/2HSYU4TvqspiLXFvfCifh9ZyQXVts1aBW97d7SDmbPY8uL0mxvCA2Hsop9cqhzWTo15xF7HHO/w
ejc1aqO8ySlRiaLw5E2On3R+mW/bc5O6eMBiGzvbBrlREjfAJxXAjJwb9OgCQol7am5aw5ybj70/
3Ru1k8Ta36ZdLtZBUNp+gzQGEnbkA6iHgqpMc7OUNlb0qxJbFQ1eKrQhhedAFol9KZT/vtITgVMM
QNNs262Qh9XmN9oYXOEmJWhu4Holr+6+GBqnaVjGu3Vdfvkf0M4t41jb/CS+E194T2bU/jTdAI3l
xECbTeNOXDeE2I3AmMP4PLTi/H5yZhDGWl/EUZkV+xj/Cg9Sgjy2ks5jmYq9VaZH/QJFBQ4l+2x/
fQ1vWB1GsJvPESMDrJPbe1wzDj47X6AYDhD/cwFioMEcp0SysLOMMOJTsC39gv8KAW6nQA333g5Q
XwymK4hBFG0fxm/0P7h3GtzI0ylBYQn2qlZLpS/LOQhpFFIzLbqPIl+oJKGrlxRhsx+v/PmKB0Ix
5MlCBjq2lt7h+C2N9dtkc6yBUwTwXErTC719nnopcfJDAiz1oZ2BsmUN26Adl4VIWlEdK5YbMw4X
m2VH2JHYlwDWglEY63OGL1IlXwwOjc0HoJUg3gMoR7Bgyn3/qjXSnNyv1HTjmyD6Gew6YLwv/464
JfRszmWM9wPGcRYrL/tC9sKMyTc088QZ4pXDq59IzZodrJRRRTWAXla/QKd4dAPVrvNjmU2g7Ud7
CpaemabZGWdvmSnocQWgMO2nS5xeq+qVUAnWGfdjKcBQU7iHb0XcKi+6+4uT5v6DGEDh9UjXiKQq
4Ff1+9yaEViRi/ePmn0mVSktl+EBQMTiD32JjwSzxlLuODaIzWDAJblMlTcVEaC53d9F/fOfmuWn
dgs5dNNIaY8sukO3LkSMZkI7J70t+iuiKh/WY+SmA1nfsO1C5DTzKMwGn09fEd3MSAQk19/vEL/r
PX8bjKMQy1bbHLfxBRdTowza83LutcfuSLmxOgy/1KsRI8TsYFHzW8kCzg6WL03kCtJNPWQ5Fnui
nTzqhlg+ue90R3qthbsfTfgRRye76wjfkLuINP5IRVNzF+ZRnVv4XZEnTf8Ys+LnsNVRzMg0arP7
+7etCE9K7ABbRBSPzqQn8hUEYa7/4bP0uiW+sp4PVG962AMP1O1vOUzwaFYHkZQTE02hqOtg/vfe
3NfR7ihLmt7t4KKm9hUvg+KODPzB32CVnERwyun5mdsNxbNBUBXlzV9qyPEnbN4Sg0D4gL3085z/
RjkZuuM5hXV4VBGd+XwkYYBZs7OFAVR7r1o5KZgAE+3/tNGaiwtE/YLySh7nQkLCBD3uGvRyCAnA
2eGcP9H0DH/HwLvRt6SJxLh3yTG6UtaMCRQ0IspYHE1D17L8zMxB6ywnPX8ayF5bTn1gweCeJaz6
3zGCXwCP+vWtVL0WP19AYG/I6qBtwkcJVL4zNCSQFqzFyjXOq2JPQSsftwsCE9iVriOdSHrb0Lrt
uC1ZZmYaC/Uy7ew6Mbp7l9oaqQeYI/iY6/LflW5LwZoxsmQuBV+c+l6OM4ky5vaXX5clEMKmbkST
v9OxHzbtVXYQePI9+lpFBJOU/5Ae/LbhQak3d7l4pbJGsdlOYjJM+01ppDcY6hCik9H4IPvd7/Fm
19kOgWp/gaOfmtSiYQwm+D/eNJ1h27vucg3Dft7fcOAL7oeWlPH0jZFrWm8SkqgXzlCEcMtR3BsD
2FYdfhs5BulC2xzTDuqAptI9js4vHaRGR3sBxxkhtd95NCd1aTHCb7s0lLtTvx7n3f/alQTHn1YH
XO1n/6LTuTlZ9F2iRtL/58P3AtcIUnVv7lLMq0pQMaqBqubtejnPKtqTYLZ++pImV3Ll90xsJDLu
NPa2pqLZvLL0VWSIGKTKDOY8SRk7qCD5w51dRHbC4vG+1raFOpwhCfzQFXbbF1+5WraTvIU99L4N
USx/pE9nJ1EMFoQHeVY7NGswHGMjqzd1jeSHCPIzuZgfGmHhZmaKJd+Un8YkbEPSTSjxGOgSk3MO
YBnQ5WDGgWFjKFtUEX7FgNLemMK4UG5lur/pjLVYOUp8KX6dCKlfZTm8ANVS0uMcoKx+jUC/A35o
83VqXe6cO+Tbui80VwZCEYzRvgvQzfNbTuTGsqCILE64NiLFR7VXGe1axZFqMoPi1TKHJpKJ3kXJ
2+79B8RQ9L5zhfbS/b0mIa0F2thTFJbRLW68SQSRqCss7idcNRVzXQVvL7jAFtx/ADIYAPkuIwBq
viXcLd+c5VX9XVLbVeN/AMLmC9Ibf28wz/u6nDXjDvH268tlqaNMeKfE2fRkZmDS5WW2TvEbgpN/
541V6RCenIgLfz+5pKHpPZg8n1QjGOWyXExjokWs6UyP4PCTeF0Yd2y3A+hq8ACjF0y4Okm73YFt
q55lLi6GByUwxm9NbwzgaL31nBs0kGaXBMT/2Lk7XZ978xKxlnX9ubLop22K9BqLkKIxHqe3QGYK
8qeaeeh60jCV/q67Kb7TsfOw3nf7Z0RP5teSnWsBbtPhmEIgh4ySFg5PwETDjFpzOpURnicrIV5W
zJYiv7zGtpuJIWBszVrgNh4442pGKXZOlQ/wHf39BwKVx5N+yGo5TtuVfWlqm86+ZHnBDj4o0/EM
iUpOKWVJNgNLojS5ux2CDbTRCHzBXgkrSC7JfwF4J1wlxF+crj0C51zmC4bnTvgwXhpV7UeQzwUA
ieGp42iDjru70gR29aatarJOZA0hI/0MMfiVN2/5lkRaIV/MfpHBp4W//C+/X5rC671wzSfxp8GC
aTgiieyrKo6DMQzb4wNZUJyUAA7zjpRfAYeu4+TjimMbwD1BC/ky8TkGy6ZeYYprZUSDwW0umJi6
rTPWiOtPi91hpo+7hmBogmh33vXA+LzfUDnrhGmMZJvUx87TsLY83tXbzDt1YgxkrbNr6RK2fmIr
X4yGN9AwkEsXdlDq3TYivSL1nTMWGpvsjIRrW0AnzCqejcU6fySZa9N/D5061zjgDbi4nrUHE+dR
ECM7xfpm8TlaZfXtRh/d1p2pvROWIuc51XFfY3ldmAcBjTptYbC6XHjlHUrFwU1ElJpYgvd4vw9a
V3frXX2p4jYjhNoejZoVEMu5GNxDgdrEKBs2PA2sQ2BQ91VGDUSSTwJnoYoScnKJ20GZJNWKepTU
MMKUsBnA9kXKyoqpxuufcwgE5z4E8iI9S/HAMQ+lxxjFYe2nJYk4PYGp4nxpbV1t3fPaTwAcp2cK
L7oF40A9BoAvOP/Eda9DYxMyWdGGfmDilVCKLsFItXMMnDTwgMX6oPN9t0YpK5/qw8+bklQoNrC8
ugWiu3IoFWIugv1IB1YmnG0HbTVpeXRDtphPnTV6dWAHVH3KvoYFXfdhdcspBMgrrwCi+QKEYzal
MiiPWJ6Ks/83tlT5E8QDNYxr5uwkXlbVF7DZHGVXa5zQqCn1OkH3UkKxRqkHDOwpLOUfrsM6VuvV
oduBup4WuxqnENgE+n0cBL7c/JY3HLnlTQul7WZEwkh1m517V+mtg/719vZfoz0xOgXeeBbICi6r
nNsJWUhkG851D3aFeLy3UMRNqEMG2xGXMil5LY2j+flGiFumOvty6GIGCG/1GmQkC56uapJjzdfO
MLar1M9jwVL2nPT5ACCkk6F5URaX8FetU81OPE3e1KIzYGSq5iOyR4Sgfh4/4+/tgSV41wXmHwl7
WFQvKxR6+RmXVjoKmyjG5ALO0hmRM2dY0A5nsO43A1lNwl7mAOCAMaPk0W4Yj9SP9ZVfc+CUq+MH
OyzbuaCyb78wve83em+xZGzY34b7I2F4KB5mvwlGuePt85u/TsNBkPJB5TptytUxWo6J7D85Z/AR
sjlTXIk0z3tXSXhYc/IBj8WzQIJakbhRpnCtOq4rEI95oRGc6T8pVjvgu7Kcy7wZ1qfA9W/OjWVr
ZnV4468XDe8WQBONc8zCJS7y2VZPsj4j2U5OK0ow1wK4SlE8rkS4AgAOeeVQxmRM3y57Vi2iyCid
66tnkXYW+I/D+u4epMFrAwCB/JAiR1mt0G3Fto0a04mwKYbOm7n8QeX/cOlRJ+6leakjhK60eAYr
e4g2lk9cKQRIlrKqXTGwjRYYw6Z1+pv3sbEjdG4tMydNomj8ZJK1qdpIffjWuC1RtzG1ZW/TBj0t
Sb4XNxwlF79Fz69C/3e8ouzoVoo5MFqhxfKEFEpAJkZ2cwqG+qv4FwEu7tBz+1612KkcKSj4Ddyr
Cs0EGV7M0+8vJtNIody/clwBFHLN4gPmeKTNty4Favl/m4FonVJN8qqOq5pkm10NpB4R738BXbrg
A7RJ/S0HcKirGFw8zZXMr+Yd4z+szMJkJgmoQfzFVXmEWy/GFvak4GlVNosHVvcQI55zSJTDZYwi
DMtjoskHVHL6kcfXC3dMKWPul7nhff/mPr3OSWvnNLSx4/zF6T9wp6R6zLgjojoursaeYpCTcCQv
OV43HbikVuphwoiR00dNjTQT4sxinIZ1XPwjNr2COxFVOGjIwfo6JkFIv/24dhQhw4RT1k/iwKRk
XC+awcLmdO2zqP/TJgrSnj71lionAN9uM04sVe/Uqjc4KCMB4xBzDTCkzejVZ7TXlxsUm2ILcgvJ
yLrFnVUWcloC6JGFD+xtLR1E7MaPz72BaSbPuwzMCaUmiGP/uzGEFHTojbjfODW1S0qd85uRnN79
NGm7g6M8G6Q8S6ggMQYC4BekUnbw7DWpK0nSGH5zxNS5FtSY0OP7Oe8Do3nJg+OWRjHTZ1iwfIeP
5vLBklzsvd+VaFftsgd2aQvCJ+F/VvoSWnoqgJM8nGmBerPOl/q2LEZJHzHX3Puj1xcH66CGSr4+
Y8TaeGf0E62OJ3GApsV3aWZlH92k74UrsAEDVI0PEWftniAvDME0NS/PU3TCdFdH7giNTAXXmKjm
ztmdV4dJVQzz36GOzKzNtsClQhGmI/slG/zLiAWdXmuLPMMIFE6xRLWNMIPMWTi4hTSWITuhHdlu
Q35laB5/9BJPznCKtFrWDgCIHcRydkHL1P0D3Qyoq6CeuabdW73XetMxTt4woaDzonxD6XXxfHn8
v6Pcmq9GXsibEb9FGDPg3qBsmeCE9AITJge9LalvqSwpteMVhTeimA/+lpNyL3NF+y73N6KwF/dN
L1GbNpD67tVh57StAgtjY/FCIJ6xJBclWmEKsCxxNk2nmTrRYv5BWuQ2mmcxUbyyA/OIEeyDQpMj
2Six9xvpcSiTnz9Tb8gg+/aQ+PKosthBh3N/3hBJGvXr+gKa5lHmE3b8AXJ9KYKnL8EsaROnlm6G
Ho9T/NLrDnIpBp0SkjfQDqSNQmPbqsxDwyCkAyvxs3TNMpMdr1i5HouKiUfBaIE+mGt1z1zvGy9V
HhHcBDg59MJKLhz6aIJ08rRrQaZNGDUaixrGuDdz262FPtRUg10brgs/DLSfz2CUWOvkV6OaVvSN
wpioq+tpKMFc0D/rxoLEa4jOEi089HwKnqTkxEkcib8/fM2KhzeD1B1H//77tSMwhvHsEQ++xQqa
ViwIteSrxyHU6+72yTatQDbN2BKhlzGn1tkawiHtZeviJhvgqN6WDtkeKtI/TZ/hPWJeZng9/PV1
hlVlhv3XjIyKq5N4cpvjLnPuKieki6On8dr3+j7WDr7W93X7lJf3gB9JHqKK9nB7jZwwmzq6OTUU
JJWb1LZqw3DKztm4dQRe48z8DcsUWHiQ1xxXxgxsE/kT8tVmEYdWIuOnS0pb5q09hSLiDpeuGniG
NzXhRBliF5pJ/Beiv6WFCQyYsrHH9qYxgSuJmmJmMes4Lh6wSuzyaPUqsvrUY4UY/9dCqwB4oKlf
IZbNp7iWE5U3gDFSQ3W+UKwqFQhuunGRYKS+Zq+Iy3PzNMVWSVtntfvx2RvLCnEhOMYn04W/mW4r
K2HtZ6ippKVa2DHtpm2SsEobIxK4bvtB8QMeYSZHCJ9FAlbWE9w4aKamSKLm5HvmXGOfnKcbeZH5
4OXGQ82T7VQqeSNBQIrVGCCpeAURNt1r1bvRJImcsSQgFN6n2NTrzH1ovR40W2LEhQZZJzEV/osw
EIaAMXhq/U/TW5ujF+VG+htmGLGvUa7jQ8KOOmi1r2/UlvcwRaIQb7QPSMBsXCbmXRmsx9gmunAY
dVhz0M56aqoUyrKcqlhCif/GDxoOMSohoHQoLI21gy+i1fNrM9cXXaVRvi31MJ6pxUZzqhoC09iY
WV6f6crncOwV/eJbaLABRg63pJBSLlMRVEYqw0n6iMttWVy7YXX/YWukjNne7alIR+F8YYiC7WPz
XPJE+UdgG7okbo8+TGg6VUpWdSCexqUUFSDScdpv6bndKCmp1nXgZ4CHehx6KJnvhidWDSP6vwzK
V8sFu6GetwS2A2ayZESmo1NuC5tiEqpuwPFkhvr5Do04O4n0nUdmyRt3xuxb1OwSbPSjXPaLfAZO
8Vz5DbXB2Alc/LD5D4Xu3wQYhLPwB/o0ckNTi4wfbsDqfBwprLNLN2Q6Di5x5bQQDkJuVJwAQv9V
djZcH9H+3IdwrgaqsuOhpW0c00b4NVs8T1iogBCHy9nt0QxusZ2Ir5YAjDpo14XAba4sAM0/tTMm
wC23cWVZI3XPftxEPZWVytfI8yL61WQ+V9qvjcbWYm76r4uiFgLC2VRE/MAaHnzgwTXd/N/fWH32
Xd+WrtKMDHd8bk+C2oIwJfPjgIIB5qsItWLN7qvXYgpz98bnADZB5RMp3gdfFRlEwKoD/Sz0exFV
hxC9/JZEqkarsusn8Qx1l7x34MaswiyZ/eLwm4ZpisGlJU2DxfkGI0xnoXbsDifO1RedYSFbofUx
InBSuwHu+R1l+MHLy594zP9L9NTpOX6DnR0UESUZkygi41/iXpY6nOqt5WqYR8DNEY1UXJ2wC6rD
UooINK9hzs8QPF119DHm/qVdEf2qq1H5NEVqjbP5qxXNwv6sjlmwqivVWQhFKVKbw2cSd/IB2vBb
sFwh+9FAjdVe4KmojAhH/htTUUL42e0IlFqetafhuoCFTAAx5n7htc2KZYZVNt890IyKCSoCxsfJ
wC6hq58LnwkpMDqOQgprysImlqJaQZ55NOf0ykWzyOMKpBKjT/o50xaex8SaTpV4G48W3qvvIHl/
63ZWk7i5NN2d+xd5tfj3BNGXOZK7t6eph4mdnA+zrBcehfZdLET8gzI0nNA66ZXJCZ/hf6vU/kLm
ao6L5+/Irs1zCInFJfEFykFvekSUxiVhMMo9vq0GSCPqa81nOhkP8OsfiYIw3/e9Z3dWEvikZKtl
McQcdfgsO8k/qynUYtEy1Qii/VRbrI4qFwDKvnJIMnLX8ve9j2fCZ67oqotEmI/B4zNwf1hVpHrQ
2aHXhnfSnPpHmdh7IpbE3AXzU50c2wnPXsUL7n46KTw/Y7WdTNoS5irZ7vl4ZH/7ArPrr/D9Sd7Z
5zk8ZiJ8/up5zZXQQO/XpajjErBUOqGIyHfBVFhm/2LWMghwOR/vyGg2sDzl3NV07uDx0jqa2sgu
OSGJDY3IpfIxCa3x6bcMR5yPM+xnrYzEJZktnEDsCPi3GnoDi0MCZP67WbOeXXuHGmZqqJlhZ2Sx
yhRpuFOsm12KOoWKeJa8clihQyJ6zsY8ugjheEiQNSobbx3GuR3teYiPDWWL6Eqkt/e7UWVkL5Ux
WRiIOToQ4aWEMYQLHDMX2CEECV7Nwo9ZY9oGwnDsJPE/PEkXexvsLYxIlxSR2/oZY8p6dDEWCszT
7OHitkKeNZQBYn/lipx9iL2Cwle35SS/qVBRLDM5anAdgvRvvt5cVb+AC1Nb6bEyTTtmqit1QR9c
d989AzDDmOfU2sFXus1KrAbp484pgB9T5VrKd5PgzySVdElW37JGI6kgJycAGtDVGa3fXQffTF7I
htsNvQf7UvJJDF4iwvyoWIwkmgZOZIGpUlx7/VmOpyKEdg8WuWGgaspofPvO/4xlaDH/wcblda4g
CeOfjB3z7E5vqSXH0XEPG0i9AopNT05vHI/jcCSanfJgs9XrAbysYVMcaTtTaQBD2kDSMc1LVh2S
itAUkSy+zgUHQx9+go+XFQGjVle2ATbneFMi32Ymh09NWl4uN4H+EVd7yyVg7WdhUJQNovWK+zTl
RW5kgQgkJ7pJGrk7LJeiwNdU4B5p2cBQsK2rjH33rfmReQR6o7FmPKg0+fT/2Xh9LqMcrhJoVEQ7
bL7lrzMx8X3tbowW3qMkAq0mSvlBrByiTi9qGa+/jBAZjRPLO/SurLvasbgub5975H3XpS8xjDM8
+lFalU7eV98GKgS4/qAA1FZpoR90IF07uYvCjkAE7J8o5n1N1PBvZYxVGJyjuwkcevbwPA+XKQsp
zDiXF8LPnAHpmyONBAEFnAQHa2eD2DtKxBW8JnJp0ecBnWv8xiZhjhbFK7QHuS10AufeXOh+7McY
NjPAhtzgxgiQBsPe8FUt346Moz51vTKi1fSi/AuXdjArahjoVgMyA5uHyLK2Yxvp/GEREQrqbXaj
EMIhHAYHfqyE9DSVQFkBR8GM7rOzOn5d4vF+Okza0D8gzoWKFSQid0xBE9IcFNGGlxK1AQS7Pmzy
7pZatRmKOAl1E+ISfpQNzLAOykAX25bmxFFi6M0hZ8lnFovAuM5zuo/mpK+s8M7OFzlQ1y+WoGwf
rEZtcPt/evKjCCfL4CyuPE3chmOzTbn4FrulUj+9j5RYQPCxkW0C2ycnt0CHRBTmanvxP8B8YKUL
dmPkV2gjxg8jPRRmig3MrVri7PLLExdeelo1+/f1vICK09+xMZLImd2+Cdq7lBRuyszZGMzct5V3
flkJCndhmsj5PvSdNhgtggM4lOv0ohRTm/lKXAI48SMhyiJ+Iw2ZFH3sdn2uD8lqjyXdAdIiTBrC
umaWiss7DeMNEEiS/mWUAWLx5sE1YsE5i2WsoJZKAJzF6Vt4V6FSBPxjd/qM6pcEhVidSCmZ92Su
D3DwmZZM9iCFdEirb8eKQ2IQzHOn9KlPWjO/l2lET2KLfnag4xC5wlGXoD9kaOThaSvNoIfrGVmk
MX4xbEQXt9BJ/U/9j8g/bTHO2qOl/2XELp/wrSS/JRE0sx2VO9KZcBSY12vHCgUWTmq0NqVVsIog
7CYWY0V4ITbSeIlOAQZFie+6pe02P7ikEu/hCFubzjD/N9kIvTzbqVAsOEZ/IbP3qrWYWapO5E6P
8uKTV3HHwjKb+nYuQqEvGv+nJuTg1A3TUXPAmFXdFV/0E1ApKcq5YtJHjxoGBcdBac3EKv+k0i0n
cx7CSicEsZTXYayim3R+ue/XU5hKQahVgxhRK4O3RnusIhVG4j9VEHBskOgWLoosYvZ9zivoJ6RO
shVd4gWy0I1TDcKeEtYQggjiD4vqBlY9emS1ZFy8+T5UiUOvsF5NmnYRVPOPQAj8P8POnPWUBETJ
cgBEMaFkojNViZjNN3UZ+LB2fgjCXexvsi8+Tu6qxv0N1zlvSwt244Zb5mtxMv10fTIHYxj0Z71G
LlDGWBRmeMlFVa6ra+btXS/vD4h66Hkx9CzAAJbjGMkL8m0zXGHDONh5h7XhRk6yNqAe0wArik4P
rRyaxM3mVrDI59tIn8/TM5L3wGuMaFTHonv4fmLvRB+RoWaRjoqNj8JbDo7Qq9RKtT5HaPngkbVP
sG2Ynpk6CLv64rW1pVO9gS8y65p0xtiU/7G9IcbVhruihRdFMwL+nklMtfh0OGm1QOrgnIFbl+A+
LDosj843z9v0CuuGI+gLJgfL+Frz2mDdduPNTThLhztk19xSoScyi+ePyKXWCPMaoo6hwQuhnMBs
OAdyMZoSkGUz/TZEZ1ARYppflNOsfeTjI0B6HgEHE7KWToZzXtGgMRW1hjYY8d7AGRPBMUjUmnSK
eLb8hbVzjulZQnCoWMh9Goif2pYdaDoT75Nvg4YP1cahACA33xUKvEe3nitaiusxpMSd2OUj0dLU
4XiO9Zt70GUg7PlTI1KPQSVHtPvaIKlLg9saQmvZkZfOaWJkBLcHrVsZKnniKzxC5vKYxromH8HX
lLqtiDxsGJnD1vtgKyJEUuS1Hh6kzasG6EBjVGYU3HuletTCLP82T8iQjOfcJQygW0w6w5oc8czc
2p//C2/b7zyxIx4sY4qZZeMDkhLPqIWpH6PXaHhlUlv5s8feTqXjNTKAyXGSBja8BtOcA1n8v6rx
gECe8+lqQHEvuppysRlZwk2sFnfeFsLagAzQweb9IdeEVa7JpXQmh/8TFIq0q93CdkQVx/TQ5Ezk
iHu0l3RlqlSA1WQC8Iz37TmYwWfpCrb16Wa7QIvraHUaGdotVn/G5hC6ycPTAR3U0unOUyS9/TPD
EsefsEWa1IitwpeB07jO7igbpoIyaBPBj53WUrEZQnvMcoCabWgy/Uqv2q5G4p2g5dJoIwuVLhDH
FESXYr9sYge0y8N0kVytrtJ0ILGj1l81OLntuldqTYRwrTMfUwA6FUyZ1QNbtfrfnRrNKcYNY26x
PgMLLmwMA0QqN7tEGo3BhM9vPrMDFzZiDEfFsNXNK2kdp8rgYZks8c/JuwErjyTymUWydYdYMAM/
Aam8axWoDQ7A+4RW6xvQxMfHKffhSubCsFeuqdeMLn2h1WKsEgI7b9XtZJccIAZy3tNCXNXwu60g
P93w2pu/RhRJ/7P+pZ9N23VZ8b0Yncy8FTA/GxIQXqSS1qEAWWEFzKYFisHsgHNErhXZLNX7G63J
iHZLlx29G75mUKSbol0+Lu67QQOEZfP94r2ClT187e6RvLFkxroVin+m6ejM/UOuYBo145pVqGnJ
pndcJQHipNl5gITpx3tw0opKI7i9eokfg1v3VCTV+Nd+zNzTPYxuW/u4opD9dBN/ZnD6km/VXMXm
grAELqVY1ZGvNXEuf0d2MJwJ8QBE0vTlCMnJvHVcNXtPfZvr2zpv+7GcQI6EyKXgIOs43rv/Ojx3
sItN4lDTSVgJJ/dPkm1saPde4vVzNmio8FNHjLJ0wEZ1ZqPLBiJHpZB+0+2bEy+GlSc86MkVrK0a
n7JuSwIYQgoaiX/b3yBWkC4S8hhATC0SnP3WBmh1NIWaJvVHGzlQ7et6cEYje0W4LtXIzklF6ct4
dcDfXocW9ghN71FNF7Kc4coKMxM8AX2ZWCgL9E7HFIOZ/s8tlc+tSaqIkAKURXgW217JuE3XI5x6
K0W7y3MZSyhAjGdslrXocxo7BsJa7yuE3BM5OiPgaVZzTY70XhHvZCsmoUjPwZ7Gzwuc8LYSmHqc
O3yef2htZtiqU4SifKGJb4GrLaNU4A9T170Po+/as4huYsXtQmpSkBuv1YazACVC32yc1fWdseBl
QnnWoaYDWWawflWx5MADbFV54jLAULQv+ngplXAuK123vutzWGtTMk8P/MPMHX/8OZIPFcz0auTd
OYxkjMB9105ibyBdEti/O3rJuH4aMuz1YzOAvtoXYyt/P2ahNQwsZlZDk8quvXly5GN38ZaXnjcT
avBp1r/kx9esOLmPdbh0U3GK8ZhZiSlkt3IlRPYY+99BEXrJaN33zoRvwGoFa5aXNhr4VExYhk+E
TVMBuk91eZ9lMPxVYfEaOjY2ACLSO5FgxEZn649KFh3wqMGmvvbbWshtHzW2ihjQGPYYumDAs7AR
nvtH5V7wt8p9BJUxzWtRZ51R6aIexuhENCs463vBuiOlxNtscwYSbEV5dQguBfCeXurvxAmo406O
CAUvOVO6oBAkSjLTogfD28+OrC+VrcVOjdfKEP4hQ2mfILdP8SIoK9JOTdhp/PaQbeuiQLU9I4q+
h7fRy60vlPoJjUnyvrNFRhjn4NmE9QWozuHCatc+sUAMv8QqbTGHDHUBtDkqm0ooVawAOH4bhB1u
djTi2o1IKdisU7G6iGGSnQcwuH/E3SnvYLPZsBqRk0ZDsFog7tWTvh/VoA0jCsS4ykleDm7PPowz
9yNtoUOMHutuoLTCS4dJ/JipEW43RqAoGzqK7KVcTILPP8MbR9G7NR4TO+ow6bAxk/ofYHsYHAgE
oUwSntfN0FzkKWxs5QwPKie8FG4Qtspzxpe5Hcv7jPxt8nZ6SzJ66LC7qrh7meYbDC8G5MhkwBEJ
pyd16x+1XVWcAPIoPjgVvDS43fxe8wA0k+0LZrAziLCeWDnyfWgzKCOolX/mYjQiyukUyp3cbNYJ
V5VPvNreYTvC8LF8ztLJapAc4R2RWB8iNque64rRcRou91Kt4qkPEfUOJSBcbAz1++2zFNr8yoYO
VU8/tiU9q/rPEek/dc8ijDmZISk/KBtbL2yehkySJH2ZPEwWzB+qsdIQ2zmEJwBhZLa4umtC55wr
jrXj4Y6B0avXsSWo6tOYNZt42e/OvjAbsQXnWinF22Igd/DSdaq9a5TEbAQ4O34c7Bnhc+gOV0zx
Vop/ukwQBjQehSG7do2W5W2fWquwJK/B0MMUHpEufRoncw8c7bGXpF17+UJokwUI6MdAlIfyXF2m
19XzJ1fvJuQ5fyiEGYoTYGE5iyaiaPgDYqtMBUGZjO0zGz3oHNTPhL8kQKXgJZ+xAINAkns2elXe
LnVZfHe+Xgd6vin7L+ba17b26TKSYqmEot2c83PA7nFcaoMymINDI69X9McwEEEKdtiR6v07iwT/
Y/SUxgQfD5hqsg03KNYmADMebPoB2nMZ98qdpO0UnSuVYVRg/HiOUVOaTZGH9sPBNTWvTbKjGUqr
Bq+V4V4Bq9KBFZajfV5ThVDxS0hQzwGSQtHLfCph7G7bUtbwvMazNw8R2q2Scz3ytuyvJFSWoIpv
9pN8WzwkXVIlC50ZoFsEmxUUJ8y2x4qpZmPmwzppV752HJRsLWxsw6KFVA5UXCUAMgBhTD4ECaR7
P6HBqV5adNAPIcQqztUFnjsJx2QSaX7/OYLI/8L9155uqLnW8gB4bbkgFgbHBRUL14L4mcxnboKw
DMjLQAmip8W/iPjVym+zR7F7gapFCnpAmIHD7io8dBYuGMpFvWEtzFkNZwmIhTIiKZRQ66tq0fpP
qkomL0SQ6W98QP3QRAi//IE+OvrAbekSZbwQBucFDoP7vc39cEpRoTdXG5J6Q2jt3380MD20a1zQ
9QNj6qVghT9493lZQeCceyx5Ri0NEwbs2cYj4vVcLNQxe6jSHuL/0RvV0Gs/cqINcoadm4SaWfjg
DZv4lKcdh+HZnm7MtiRt74mLswsLZD6nZQmOoo3Tj8DUdOSmNLfh9BPiYQAHZGVHjd7HCgnPSDp0
4iEOHMhCq52zto1cENzTI8daM4ispz4rBP3emOUET2n/JWcS6Imz9c7F84s27lU2LGg6ywFHdZNa
TZrhjygsldiOnLT6slVynvUPg0UlklfpUAcQfLCqP6fpFuPkQ4ZIHd8iby7x1XdRa6gjKIxG+avj
90hDWa+5N41bT3RxuIwmcyZGxFL80u7c43z8/wUnvjnK5JZ4iCi0HDyDrchEjiwUPN9eYJG4K5MU
fDPBqhenqdO5BLyAk+J7AopwO7WGeuXBst0X0fOFTs0dRAbjwjgouVmDqM9Upe8ePhnkc9CbK2Iu
opK7ISX0ri5j57fv+IeWJubEBxF8jFDtGfdHk6BLpFZY2/nnzsyQOg8YYctjaXn5Zo44Imu/EpRS
XwmXQ+o6+3Q8m2UAKURETXpomB5IWOHVXr0r12DE/hWuJzX0YdsMhgVZyf4fL3VHyFWLQKJtLxVB
YkzwM8Y2L43k2yflroYsdq4jKeelpNX5TIvmnT4rHuBDJTWLbbhMGFfFpXzvtuTL5kRqgyhTfaCf
Six4SGcPL26+kSoh2ZbVRD3n+M1wOLUkmfU1l8jMqdq/Qnpdol6TOIdDrloObY03OlKrEkL+mEjs
ENGJXMHRiBPRlBRffX83YsRd3JbdklY5vWKFtr3dS3O6GT7ojcQ8EcDJ3P0/PccX7qHWsQEhWdnR
Kwy69I/1ZXnWUjeCgcpihAn3//uO8gphnlw6njr/zJeEkx5JDXdbU9geJ3K4WJc6M9cy2u70vQx5
EcYFM5qQncjwNw5Gu2whhp01jDnIRENEBJs2b7KsDjVEYmDOlH9tZIcm3ujyLuHjArqZrACmlLq4
fp+lkxg20M4d8xpIou2EwnJjElXCBwED4GTQYSBSPLvlGkIfS6hC6VDCV685RiPqYtCpsgLEdmpj
/YFY1PzaLHX9RFKS4gcGEuoz4biOoitCyPCbEmV5v61JUiDql26fIxrkb/BUVjeIPb7yy1GnDnGI
rWrJ6bI7h5jxsptMHTZcmRlnUbnr2sNZEMscwx/g2IQHQ7dMxOHmYAwNz+mnJUNg3dKLLob3r7Wv
opm1a6ZlM0VCvWP75giJWsaBiOKgXZBMiCFHwZljf9TcpqZIQsqAr7tO1W9IAvO52IILv3+TBsM5
TWWrFX5YbvtI0lDeSqfRK80ITsgyTwVqP3AJ9Az4phVi9dUdwR1OGH3GhCXXvETT5ikDhjddOpS8
tVgZJqPc6oCJRS6e3p8RSj6jtwm7+igu2JCSEKwyHZn6+na1NZHRm1Up+4NuNFfh+7/irg7Vc3y8
+laAfHHyq2heGdnhykoWq/12jJtcUzXDhOXuU7gTazYNCnlYvtKbWMiEZjFqX9PRSc4WC7fTwJfD
fl+8kPQzE84zXY3Hq/ubRDVcDUXxl6PQYN63dMBzdAcAxVt2u5VPY9gO/P/87emSVZm+K3ZGlia3
BV5wnGGhKyubnMI0LJNGqNCCCOjUXAl30pe2lfiKTtxxbFEftXqSfl6InB/G5XlqbHyiOcipE7n0
xmEpX6xK+VW09pNpsypmvHgxclD8vw+Jk5OsP/Olj1JREwF2vaIB0Q4BHbpc996VV5g6UAY4Bx7J
bEv3V9AgvgXhtlSJcHk5vkZAugPBZWDVQ9bh/bpHkI+qYDkvet2kki11Z5CD6rbjO+h/myfZMsf4
UYEhZMoobdg4wiqRdvrfnvKTLCm/VxTruAmIqtTz213DtpDPrQkC+3nmV4YuGUKxY1AbEa1ng1uC
DBh6c3QM4nip6ckvbAy4I9ul8O1khB0Xp/BRr1V9ojthvfcr0unnXbtOVutYofJyYMQbyZV4atMV
sPVg2WQ5gtg90aSR3d2YbWmp4lptZwXVp3f83eOC7jtWhqoRfeR2HTFDtySj18SfHEd4bTJRbVD0
njwERkqd9OYoPsjsp32QgDXwnmswn/oMsLayVwKZkw91G5N0FqBhj0m7jAw7nFMRBbwbSnXK/Avz
Ckz0lpPw644vn9VnftWODpX1ou2QfbvQ2NxKDtRqQFkPl9dIGmV9/Z0on546poZLiXGWR49M0van
HlIb0zOwuKNOrG38GIFJqXhj+BGNsY9Sh2/K6V0Qd3jjrxMAi4eNhWUJ1aCRWSHV0CeFmpfLVrDR
4Yk5IV5oItkya6mzXVxF0pH+y9glAWoiGfJeyUHQy4DpPGjaz5M1oeW0xhmp4wJE53FvanDsGhal
NTiiWW4KEIx0RcrNf6jx5ZVCi7vzo1PDV8wpvyRj96mmQshoJ1phexKGMMatHLHUrJsrtdvD93JF
WKaf7KSgOhs8lPNVTsoR2v+gvyf7OyxtnPKIDCoG7NFUGJeGfR345s4N5KwWwigaYc1UAR9nIQzo
tduLM8ExRNklmwHqhUT4fN3WnFdsIy/SVJGvxgcjQM8PN225axSiu3K1EMeJ0LUuGJhjwbdBDw6H
Ig8ZJzUoGGuJUcQHEUbV9l/CWEKuz1Qf/UxYxFs8eLq1n40I3EtTsfglefdB5YvLqAgGQiRknmHF
hzyyroLP1B4NOLPaKMK2Qu6aWRG/bgHYIHAfaqCd0WZ/TKYOuoajVJsnuChXfpK/yS6G3212O3YE
/kxd0sEZ7p0vHnL3nFeDknHIkL/EZdvPRXTeDvGXVBuk6cVMYs1XQ0jyLwAnYDz92vZtm9vcnEoD
KMej2URbyQmoCgpTW+4OMI44t285IP1NfcEimmVFRybNkbuhopFC0RWq4/Qo50WXt6sE+qBhGU7R
YBKqnJSkq4f7+Y0Krw9/xLpW8U4227P0R0HOZnMOqSrG2RaMEqlzdYlObTCozo3pXkca4oixl+W0
jVrR0fZUAmyuaSESoKLWPuKge1m6AmKZTbgSNrK4cOqRYE+kG1Yd8xslQRDuifl2AZeyVKnn86PX
YvnLb87HsDsugdpwY+Y4POHdjEvtpr5AW1K+/pxC1zLYzzJwEPvY/DpwyB5iQYp7Uwo6/dp81T8T
ZZOo49CqbYD7zcG50EAVzidlhPwaWSToIlfAdDHtFtO2m9Cg2ZcdQQPcdgDTLF9fo2P58PR64bY3
Ri7ZR4p/Y+N9SX/WckND8LT7kxCrzIsgXDIhpRWhZwW+q95wi26NlNNhU6XHpOa2e9WdtK3R0Qt2
D7Pc24BsF53OCJOI7EpF0qkFL+9lZLRkCNZPnLdUO9j1KLH8HFACWlO/vMTs3RlOhARsh0Vy/oot
/zyTRlay+ZRT07mXAshzv464MsI5tqfVLuIvl0wZcuKZN7ogM8Jad6Lez9ytzSaGqBrACMTug1P1
yJgjP/Kb70siAezo74Yzpkm7/dyaxNWKkYcoLNv6IfchkW6frzgixtg3Dt/cFmhfxcBgLudcRez2
s71BWTUaMmnAN6bdhfbqmHrufnYmtzXDwbBKoqI7v7q592oGjv9K2Hiag8MpPOoWd14mZ5W9FeKm
aTb8IJKqUgdZKW8TUA4J7vEGtofkhs28oGSlkXujaEQErnD7GjIKVOn2lBH4Fdty+tWf1L93w0Vt
MFN6SDPBwzWsh2Kvq21bsYLM53LH/XfO4VfkGS98ebRvOTyK/KwkNPVv3iO0kmh3ZyC191Ypyy/x
5rYglsekeOHJ8gcOgyQHZ4IMgTbz7Rc1bankXo8AE67MYXdNrRvv3lBs4fO9rYl6eCBGmMf8tE90
NbXuujGz5Pp50NpUnSFaVQpBlY4t6PIhCLdmz6m1/qLFp59vSbrOGlJN/tTHhjH+LvbgS1l1joGh
vpU1uVlswo/mkxytndiN05l2DJHv+U2juoptihrdFjqkumQt9QdJQgF1BJhu9dVmet9G/ziLYtUs
kRdlyyPTeX+/I6x/c8qLgWpgDyjq/8UXbjd5BlcTrO9yPF90y+kXB7iz6GyI4lrqTbjhHMEbkOGf
EL0Bt0H4q0IQW0TmodLFX6+aMTwM55ylnSoHvJYpSM4Jid/aZXRoz53+PcprarHH/VM6/S9luK70
yS6uXiL2K+Anmor8QLvJfASZE21al//UrDKPCldzH4x/vAPLqK5eVpiQoldFJDOnqMMpG6u9dmk8
FRSMaCWI30WsTrSsRjr3dRn6l0csA6zspQQF3F14ntE+0bwj3oaZ9bs8E93jFAovBmKRF1gbfSmn
gxWFfAfenDYFa8afQS0TjNaslPAtdQyg1bIyYGOUnucx3jsijskwFY1RHItR3obd1pCIpXTpq8Ug
dVLION6ftNqlCqv8QR7NJjQjpbIkNZQV3eI4WRy/Cu9Wk8mVCspPwzORfLc7LJUfqGhQJEo2w5Un
H3sB3qDXw92n/YLqBCL0yxHrnZJTsTe7n0PFDZQHTfcWB2oUsoOWU9/BgZ1ZY7nANJYeeT/JkguO
oOzJWytPFvrt8dLDhI9/nqIKZIUy2rfWZpLvIOBOWor2NoK4Sj2cNuKwr1ghFSCNF40xSCohBRri
NwkIiSYunJmFxuzDJNHvg6O0Fc5h/8yxJuYX8fiP3FN6jUatu3FO1pY5ZLYPeY0r5p7C+Zm5rI9Y
QkuUkEMpH3QNwApsOO5nEzSCMVwXSR1WA1eiXQsV0SwdnPrEK3raVHKT/BckChY62yBcm/OHF0HH
9E2JN4xLQSZIUwoBpci2oYgZolqPvRl0FnJXI/NscRQ/Not1uRkaYUHIvvSyj7D1kLgHm/xCf1G2
l2S3t1ScE4RgpDwR3+miTE1p0NuDPcsk2Mj4hV54WqXIh4x5xwbVRcLf/GBpPvgo7Vi7EKKLtRmn
BG2HfV3gzkpBlnfQCrbden7+1e12BESM2hH6KBHyw14eA8OPR50mpcJRycDqqYy+pai+RcoUFkgS
0Z5Ecbi0YbNdLB5nmB5j6cYxTjdQQQtVmW0SI/c1z6Jo8ypMhHZrJmumoAEhkcSNL4euuMgmuuWr
CrBqd/u02Py9DrWvQnFnHA/RezXEUt8jSF6eTDCrbprvToy7mSjiWQ9GbaPUJzGA/+qvo2fu/YUz
LirC/wPx1J1Ek3a+YV40Pp3OFaa7DmpvQWTlvHwXs0pItAaM1E83hH6JM8GYshDGV9vzhA9WyPp3
902W9S5kb9AI0JWyoIe6Er0/fQ+nwsicOaHV49SFKhambjKq3JuMkMctANDdOyac97rmOl4gRMPd
c5c+ZhrMJvupC/kVgU5XFWeiunX59DDeBkcgBpU9crg14G55tA+CLvaWPeX66RAKzy+AjBcozuWA
/jJ1lH2VuQfQ6QpxU5HV39oZ9Xx6p2LokL+Idj2jx24w5loOzoDrz+yxKFUXn5XiXXhDbnpToYFW
Ew1Pw+hBYjekQNsxuv1lMOj9MbZp0Ch/++d26mpPqjm73CJefEp0ldzPB+MBtQhVvn6wwr/CGUOC
Pa66SIWnMzGDJ05G4cKJTUFqcZyUOIu3mBTYE0Yhtb1V3nLto7TA2QjJ7dSL2Kk1dcM+YLuKF6M9
WHOe2qxi3cw1hEkk1bLoUA5fRxVZaA+hBishwwb8aM/LgN7a1sXspUFHCfnqjZpLjifm2TRWvxBE
CZZJF2KarJ/tltaRc1oVNWkhKA/x4Y4Xs3ePYRSaoHTXmLXx1Y7lLX58J2DV5GUhlVz4Dqgrqi2S
S6J5kEfyM9wqRl1s1yIVdnrVP3l5HbHw4em/S5boNH7E0WE3FFZcEYaztlSGuOPKWT1gxrfIROzC
nKmZ9PZ1t0uJ3Cc8xapaB05TZ2J4dFTXwfr0X/huqlSnnS2RzeHVoku7aZFO8q4996Uq2hDcVbwe
wm2INyQcc26eE7LNVTFIkCfgi7ZurBETxsarTG50iVziW9AFvxWkxT1nDbrJj8bdXQOedNuEuK3h
dDFkrjr4yNoPhr+2srQHWv8f0ZqSOz55UBeNf30C/pdziYk7sxCEbKj/nYVucLruOzz0G6jMkMqb
DYeGlpvP4BY38vqCBD1MIO4UaVMHmDwtvNDlYEEqbXo3PxHtzQnMDzEnKmNt0fYseQuWYOn3x9ek
Iten3FLBgar0oUlGLofrdeJ5yLtiWDSCpNw+owaGLaGYIR5wUqYUSq3No21XD+oYwI6rJJ/qhN6U
0MS5p+Ld3CnJCtwBbliniuKcshAtBzlvpe+N7wzMrNU8FDN3EddYw0ozuXY/a+5vtISI9NS6uw8B
xsJut3plyfyQU28FDezXhPOTHHdlyjNPYJ8wrDIRv4FoG2Z9UzbU+dHmLD3afLHQ7HuL4MD7mGDO
sPyKapZiQ9oLrWUZQZRTtn6UlxvtUvVnLmnrqEYmpY2a60JB8nAyPvpKTIL+rTahxCulj2Tp2TDV
F5XWQ7WPrXWMaag0tHrK4OlmmdzwUgDTT2uv8wNE+mzLnJHBiJdrgmL03Z6rKe14lEQc4//52zV4
hltXZ/G1TiPt5STjE1FZjBKVLI/rgOExaejTE8bWTV9vvKSswjw+lwdSHy/KqoielnHoDPF5unGP
tzh+dAW379xQ6fxRpueMmbYvzyj16SDmspXYbQXEJWLlAZKeN0rSWtOfrwxUdWCggYtk41v6LIGm
5UvZyxMOoP8TFjNlQF7BJx3msH5F3WliSv8IWdAL4VfwoEJv6mDC/jxXz3K2UN0ubw6y2EzHhdDa
Z/knLgWmLxfgOiCNbNTF75eqwqYH0qkTSRS36PtOG9XXo51DTyEKl2HPWN0NXruNqVU64tCUcRY7
GFVxfKUiM7uWn05Xt7eg/p0preJqubh2KgM6RUVVCZs2OcRiOX+hHwT4vsCelFeU3PopkrbGJgX8
8/82Vu/81LI8NrF44QKCtrocH3IdFqTNmnq8I0ZoN9d27sl/vP08J0KcbN7snyHswhM6fuV8FA+5
Xba3aOETpTo/pfWWwYZ0cW5gvr4f7HaGrU6DGdkeT+ogL3INow8Vlf7WleUDoh9s5XT8LTY57WPQ
IGho4WuuoIgYmkmvz3bcbcCFP8+hjlzfFcxfR/5lb9eIUX6+XZ8kz5ZbMe0jJEzSU734tbZZ9GFm
j5RP9W33/hsZhAMFzdRYB7wLQLD8QgkETFEPT0zWGxb06RfsjpTkdNuZsFilusSL6xcmgqN+pJ0T
3epMcjU60Ke1u/rS1/D4Kgzxq9Dtg5/HJ3MhchuX45x3LFkQe7nYwnGB9sEboS62NV7bDcJq624O
HBESHLkLWCAwubWSIiiHjTItefiM/ZfeqLNtkMzuxxCRUVhvD3CawosPmrvvNxJulArFaSP2u46o
fg7xylmyj59BAGcMdMZnYIkFRMaVUHmxVjjVt3q85pU3WS5YXguyqWdOVQOUJIQ1gvLFvXxGM9la
QlEDbONyDfSs++cLPgSoeRkBhCniGdmlQ5qP4Cc5XSWTn9OvWyoTlU+3Phqrb56e1VSxHF9DMbW0
GMfnPz0GGCjGekh5l5vYG9jSLktHB7tjlLdVIcIsg0i3s7yiyuyTgb/NeFHk0aNvhEeZfyuMX0Ow
rfCszJWinkqwR7qmT2mUSS494n5JbSw8duTSBWEFXjVhK558ZMAGVFPvv0N3vdhbpB03bWsN435a
rxyNe5Zx5nximmjyHIByNYUEAHbHZ5aASCocfCVvp8r4nOfAU77pO7434a/WgiRo+DCrAJmdw854
YvCe/0ngiaLpQfAGqHth4do++7Lxl6+MZ+VotKKa9uVqSoJJ1Dc33ArAp5InQx7tpkysZ4QsP8mu
qK6XgSD8hA3rCfTAzPJjMHXSnKWpt1ksznxlPaAK12gGrGAdaj0Y1dRXJ6+EQVoHB9Zwo8nRFSEq
v3LTsUdBW1AdJmd2pRMQpJBpzSpoXjQM611+OiBgcWJztqfYEFhr34mXl/Gvd9lcV4QIBH2OZ5nZ
WcqQ87hsZ2PXCD78TTWcIWvFXZTXZDa/eFFZAO8NlJf20ugvH1GMpKHJv973ofa+l2PO0jVK7Izn
3A6rQmj1wdeBcwouM/GWZULF/QCC47h6Y31beJi147ew2FB48+pNpZ0A7ZMY2FfiQ9swvvi+Ezc9
d1pePYVqvzJ4b86YZIxfX3Lxt8rj6jsaO1hU6haHdWvIj8X/opc7UDrlsNqrGK0EmicBgajM6mXO
xWF1VJoy6TePQZTbU7ZbSwZ60XzcXxiiM2yTu8taEN1XWHDSHzrBOivaM9pRwIAbfppDIgQTe36g
oY0yCNhGfeFPXw6spH8iYP27gMEjOh5XP2FNykkzp7fsfhZJpiqi4/ADcFjqkT8qs8lJi8Vz1EBv
oqI+JX8U8Y3x92d2jmq3ywcXuHqz0JbILHpYwSatCETKmJGVrddh7uvZOQMmjIRPmePvMtVfhUZW
+xlobPOfjx6doBkF2UdiBanqEEW1Kc0+kLf2Ulpna2ftl9kIHCTXLZ35dqxVBTE5ewy4zmX8AhKl
4y32TdR0qGGasNdzdRJtNR3nDkofofb+R0hMOLZnNUfPCvE1RUUaqpS8aBQfPoW7UapAtRIQDwOv
m2cjGValepBfTLZf1Gw7H/JcXvipdSt3ev8LbpSrwePOcddQooVOt1EbHjG8BkLQGon57bAFN0Xq
dG+wJDvfTKQxov8XKz7FWIpdJeFc/pomOmAQT4jQEIbijwM+Mb6wtaG0qTnjjryCdKJrzpnnugiC
+ba5wq793T9nw5SzQzAtFYh4mebP6FPx9dDts3l01jKmisEGwRTpsA3i8DW4fcQo8ak8osiIHezz
aVffNwsOQAc1b9SsnFZ8NTSHy364oFSX3RUzqaPYJKyyXlwTJY2428ktIxe4/R0tl9fE6N/zKjaB
d+Jee1EcaUrFnQ9iZ/2HUbNIw3SzoC4MYZDQuCdCodT81N6luDG33FV3SObNllGIMdG6IEo++yYJ
MXw99wMZc82ukYZqZM3WSidU6Ab31LpIzn0yuvqsvzzAH6KNtfAD8GLekJTgNB7AVAXGpQoJA81a
7j75g784nUn+q+j7nBwgxaHjMeobdn6saFaLnRBlwzZSqvm6zfdK7M4uFUuUWeKCG4LOZ4pK1eGd
rU12cNnyUTYkJ/1/TxeDW9LPwEyghca8Dbm7FW+XYf5v7M4ksoVhFZwy5xPDvESwdv6AiuEPESkT
ZIVgHUXjM/hPDL2aVrYO+poVI3A4Y76T6Mt9eWWOmQoTfTCUQQbP9uSG2GihOOESnaG86I0jyZRP
O26DLfneMVQY7OITfQx+HXS0LtZMjWbcExj5PtrgtyBaT/VQUHKc5xLHki2wN2lWmASgC27O1XDx
hcXt11/HO7B/ejEkD5JtCGaL8jgbgGA7ayLw3QxZw1q6/ZE65vUmpCOv9B/Uybv5ZZYmS0QUonh5
eyPU/DzQljcRWkyt1o+R9R/FCxGGLZ5qqR8jjkwEe+M2ajh32SMDX5P8OkIvOSWPVg7zRALBqEgy
VMl3wUlrHcop1wFC7QfCS4KwJ6brWh+1QifQunBgiCR8O/QToClSHN3WIbDu1JkYgQ/ZbnpL9sKt
CHCvynFvGlea8d3B6h3I4TcSuARMo5hZgGWHzQKA3n3SZ6ev8+u7gyhgV7fi2BkUwXEiqW9Dyf0W
PtEPAZT+3xGTnaNx9+ncnetWt8H5YHVKHWBYFn7+WZjxxZDA33GiKEoqmNYoiUuUJK2ftR872v6n
YJtfF3HdJIw2Z8P+QDqNZ5memv69hVPp/VviQ2XbPxg+d7yFHhdLhGZXy8dSyGFXxX5hgCAVTF0E
KltQ81bGjFCvo7mDDgJC3qqkMwfMLCtL446SA5lCD50ZvMqyWbByw4+Ib4ySzxlLr0Jc17Rgo5ft
gDMz7mQXbr+QBdrv5LMxTyXUznDSjLjxfm8BkeX6S3eHjwuW0IvK1uEiiB6PeBhSR700U3Y8YBiz
N5vlld4JdQGN3h2xwNLJLdevthcIidB2Ip2h+tz+GYTz9ITPNaDvW11XhQKt7pT5wZsRTHikAaR0
e0g3jsLL6jCAWWAtqp+OTZxyycyBOpSwivsRiXSHPXpE/83nVssAVvP9ICp8+/4E30dVJv3D0d+9
6LkPMbb/N54ko7x9JErJ3SXdp6MEe5zW6FLrYnyFIiJy7Rdxy7LKlxHvz8/lHgsEaF/6RVeF/8if
GcFICaCdoEf8c6zghM3sieKQWyA0MjoGKjD+c7Gj5TcOzl0Gu/zgmh50ruwDp4r91YRo9we0yMd5
J3PSHVIAJ7wO4Zw1YnW5SmRs5cyk1e8AHq/iX/TTcHdoUSQEV36FR15TB0FyZSwEtAVacHo1+aY1
O2ytgrVZX8bJXQlPrmeDLYZJJsHYBHUz5B+Jr3xj4xPxk/q+ZC0B8s6mHKA8ifQToNm3dKjMYjRP
17mERvaXEqEuW00PFCWdij+96NJkjnoTzl52fyXsvIzTrfpVKU5gRtHs/I8q3/D1Z1uh69Gf1nWz
oXtl3ein0DePVnouWv+Lchq64ymTAnjyOOKVQPEsKa25Hy9J5kX6AiprQsbIdKiqSTU3dJwORqb7
ZFzkW6b4urBFPG0dHAPAVODRHLZX0T/eARfvlpu0jf3n5tCyeUtL47nGZukJwHAQha1ciNoLfLjW
jjxhLoAK4SA43o5S5vPyXijW2RcZgI98m79ADcgHDY06nP+XhchpTulH4WWqJX70saqYJe+c/7x5
tQB2OhjpBJkJoTSaKN8M2txnoUQrmIe3zPp6GZRE9Ab4Hvk0nR2NW+K4UQIERUn+YSnp2vZ2Amkj
7NwyAniS9zxGDSwR05e1YiPy7vMqBAHQYbigp0ARaIrem+rtLvoI/j8hcF9EabRzQj50I74apq+y
GH6cy8qk/bT6R/pkd0sw5awx8C7lOtQZ2/jwBxtOp9obzN7Fn9l4BDj0dXs69W0J2sVmrHpIJ5Z+
DfG4KxAVQJOuw6spfiF3hUUnZs/X7hBxZKvt94YuMpgdxN9U91rhqxTqnlJJOlMVaWUgK9ELn4LY
jV4r8/HXadCdzyHR/whpdWV0Z9weVXY9NY2xel8hLMJ1jIXAk4/lLybLTe2iL6nuOxouTPyM4qg0
5M6raKYjU6h1NfecUU1hga7fixFjopKjvfg+cw9886HM9P0OjQBSS+JHQRpVef7ERqLLTAe8xJDE
+1YIHDvpbpwuy2RbV9QBIUYep+aEm4YCijn+aEt7d5HtszlpM10eBQfoPSxA4AnRzPEa6IatP7iI
4dwUf0NLSFtO/1UyCGpUfoudXblNmtxq3+oIBdtU7ombF55SK+XG5ppkouij+RsEptfsoUncdN3p
lvmxnA5/VmU832RDNyqPRUzqmSSc7lKQzGeitb5r0wmIU5eo3SUR5mHmDlu1UViAFke7XGzlUZOg
mhKXa0XXxpixn2XqQEfI6Mxi27BG8mz8w1xtzYwjja0qjPckvpVbtLn6dioCVsh8V4kaEGwRm2p8
j5ciiv87YFaDOt954U5K6Kj/HMXiK4/SXdDAufJIRDzheT+HgJVOH9XDEFy7Pnylq29PCqaxLSUi
25rS5V0AKehzENnZk/xBhNWywsvtgqDOyHRUMyJTrELMC5tZ8Hz4XFf2Ts9bPc9MN/yrqRd37adN
nu4hqsey3nLdf6W+qUEYMBSQNr6NSsDcVBQ4/uSe3RCEh0N9oc4UL3ALN0CFTOQFkGaGx1Fx/HWF
wC4Cd3Tu+oKds+oUqLZ0QlDMl1XqpLu67IBm20knFWHCBUqByJHLKoRA34AWgPdwIHd7YaI79cXx
X/K6LzhDNhZuQ90hZ0RkyhsvY0TMQ0BGwa/qTvESTtyMoC3EMhVGMZhqffRJb3SJzGincdlR4DUP
M033bjbYnRnxorckbCaz1Dz0XsgG3ZScVqstbZWi6fax4oIhNkhQbKfBLS3BHLzPRHkDbyQAoo/2
UunPbH5k/pNbFQ77+tKyN85hjjihHLLSdV6QsjBdkTE+PKHtkItZ6Chmy0lY/pL3yAIV3XP7paVp
7mXqG+jNb7zztlx9CGX63UEyWlB4r48Z1O91mXl4xzV4aGplVawfQpFZtY33g8n4BA+RUhL4bONY
Pin+ZSNb9aaFt72J4qWzqPLuGoeVnLWRsuHCSPgIhGcF1A0xSFbMs87rskL8B/8GyYpFN0dbcVoy
whE2mOfiaG579s2Zbvd4IQwRsO49OgBFAIURhUJAZZe7UZBvE5fFuHY2EbGA/QWhKiB5vJYmD5Gf
h4aAHfltHdspUqOChtXMjhLPzYMoZewj9CeDXBHlErn7x57SBQk8CjU4GMMTVD3EnnjoKF304SbZ
PvP7poZU6YEkeOfk4OTQzzp8MdghFIkcyME2t31xcJMNnFlTBw9VF8zTU11rtlf9ivLS+bpRJPEF
Me8FcsZQ3nwRsU/EchYwiQR+4rhKoPZ2Ij7fNodRzdKBTAtLwPjOUVXx9GUKchGwCKiQ2s1s5CWo
B4ybJRrmh+GvqrnnKHp2iE3dF4W4CTqwARy+N5wiIBouMYzzV2tlEZuYZGCvQELnMa0ZR/2mOYCz
aV2A1+eGuRB1sMhn38mdU9P61xJqZnH4VTYxEr97sf879gA371qdPgeMg5/O1UNPAIpYfZGAoarB
aJfo1KIfNQV1CoJs4bIexAwia6bN96FMbYXCQG0mUrdv4IOSn2jqxgH0OixYharvTtIGM0E6HWyV
QFJ0nf77AE2B1P2K6GnJhBC+x3S1+rIh2aVLyrPYH2w7d7rMTCRFKEset/I4/G3MCT+tTVpAUlu2
2UST7AwYxs9OqxnQrlWdCetWyD1qSVpmb7ks12Zsx+GCHQE30obBO2Rz9jxuZycaTp2HTpEoHlhA
gm2zWKqpYVQcBad6Vy/W1rCnP0jfHdFWizWmqrxpDPvv6CJiT3hbMUf6tlQu/ey34NGU6aTAEJQj
oOO/z/lit1gfEtRi+FixGAOktCD1oJqFcdtfOVXhZ2pui1S0CDE4n8xfKSo3Ks4+MTSh70WlpHqv
XVCXUisgKIi5dqW33xpOxnaF9zik9ePCk843uZB5RPbjyoW/3AFvNRm0/08pcNMJpbsJ7smUm0/k
Y1phqjGC1SAZgLdowYNvDfss6Fnxfa0s88tpgXLA4KXIrz5HNY12eCRim0w5IjwfC0FSjTk8gFRd
8BC7Zb4gD3h52bA+9s+1IXvxScDEnrODhEYQLLp7AibgKP6Lv8AcWJ1jkKOpQZX8sRwZmHBmht3r
uUxOOn1MmZINue/oNUhfuvj8ot62hSXhHXiwy752k5E+GHNMxWKY+iiFUJS1B9khHWvhLVxib6AQ
rmySwqEhLdX58Ph/wiSDiMTDajE8U0tBLpsKtN3lMhiqBefipJ3DzyDyKX0MgO6iBq7vTNK/EXV3
NzWRue0YwHfuIyFas5li9oHQHDnxFv2vNuGXNbTLIdrJOd9WsOQK5XQrxyoVMdwFxALZHZqqG1P0
J6LNZvxrhZ2EJIjRZYhJYH0QHNf06A4GnqW1XSkY3LDvX2ZDvqXWeTg1vN8M0Vp5FBmnDYJhbFQL
PpJamg2a48CujRGVYWGLD0hHnV0VVrXCPq8bcwPZvibTzELUM1T0NylsYOAJGL6qUe8fPYXv75aP
N0+IQNAVPvwnd/Ay92Dj7Cxv1SGX+S0wB+mRvgKZRdDQLpjagHgNkwmG2R9Dd/7mu70iqQj4ijJa
G29E8/1TRCJ6XadjyW3CWiZ2DAgYW73EHnpZN5HPQ7rwAPR4ZGcnMCrEsSPghtbOtuct4aiZGEl0
zJ2Tq0YCtZkYXdNAirq/3N4B0SM6udoSZwugfm+BJ8/hGc5FcWihBLsGgWW+Zqz558pL7sbzWFHH
/5WWTwfL+e1zHfwE6AhWsicpR/GNsphVqQJqSYa/+EiQbI8iV7W4glHf7AAEqzZwI8qj/w7+jpX2
DHTUB9YO0SY3uYHqOOtmgZtyRw4EVJVF91bQy/Y2uepxAslTPIszBrNhhkV/vkaxNButpRVOeSO7
OtfyTjApwFKD7HlVlbTW3XYC9eUS/mICdWK3Lzl+RtAxOIPD5Sgva7zMvT9yEDAI4MB+UDO3dlrf
JfwmvvCIYOFYey5y81qcPODdtupAjz628rseAFUrNpZLBvNyHm9dVEzqMzhstPpjk+wYz9NYbMWm
S0/J8U2fAo+09miKOzdXBYt4lDTfGONTPCri/qremBLISC1yCnWw6l5C/TpO1S9UvcELJ6+N0PIh
mxY3MZa4c8ROKpfaonrnbpBGhFDiVZxR0lxLKaD1/ROeAHqbcLPon8kkr6BaxnL8gTeGJO9iUJeG
Zf3j+P+56l91bKIy/6qoYj/J4oJZRspmqZ2V75eg2rP3AK4HsTBlf6GG37lCGA9y456NfXdlNqpZ
MP/tq8u/Fd+fa1tkkGJ4CWIncxwejtZG1C4HNOM8Tf4bTLVoLQeWnyyBK+sj4acNCXqBDpE18fUN
lHT5TfrZwywFMqh1YSPfIKLZ/7RyeCHm9fx/kfeN6hW7Dou3J/fnySSJFvWSczgM7DBrFYl7n4DZ
rW0UVb5Xm829pOTPBLUme3cnkivzn1ZSVsfbpdtjMr345YrEAv0EXtxY3z6Xlv3ARCLADFnTNsbl
mlJFmc4vj0jlkURemMHX34fgZ529QHIelDAOtVeuO+nwav4IP9Af+VpF2BJCcpNrwTTMBXbA8p+L
z5gcR/BZYq/4M9cpW7VXUUr4OqVGQ0XL5P4iUsPviHTDak603suhupcsDDu2gdFXRyf2yR9NJD6U
DkDRfUgO57COz2Vr96QeHPGjzRIlt+G3SfvBdYLNh1aIoYz+CoBbHXhSwna6OOfHQmcFLUoTp7AB
2mTiuqyRMp35+bw0cdgl5k6WsqT1Zzqglb0g13Nn2Tjugfs6tKWN+MCXOLdcVbI9kqCkxVIaoZUg
7pC1fjgjFp7t/sVmBIEK9P5F0DJDuPt5id/PSKiTzDzplwmkxwMX11GMLwzvBbMp+gnCc7AWWskk
gmYoY6d07i166ruSi7EE/bYPhi064hfgiu2qzLhmmkmhSk5qiIxtoG7KQbJ+SkKdXMQFSBHTOoTM
x6TL4UoAGSLRRZ1lJpe8AVXmnsN57DXhBfgbYHIylQ7rVgt6KU5uO0ZP2fWxZEcjRM0rVP88eE0U
RoMc9LLYveOJzhQAz2idxruLwFaXytkTywLpLZY6h8iloWoGSZ2s2ylcCfTVlqXd2GBOZoHlISUD
LmLrKxZtDUrWN2KSm3Fyl9sxiABD9Ex56a46d3mjwuPU3m5LkKaoZW3/AWVbPmIsMhRy9cTEFLNb
7IyAfJkS5olIgcD75pWyGbXKq+UFijPtF1qsxVeFzC226DaYlegYZqWj0oH1AKAlCt+PHwHtQOCI
I/cCryvTjl7x7VrbL0JBTS+G4V9tm5S9cQ9ikBoOYieCQzsSY9CBI18wRNnq2GkQjNZKBmzZXfRi
lGLRHCETtBxgaTJ1jnjNwqvgyu3iUHr7ImvorvnKF2YlegaSp7VHn2V2MAS0CaN1e2mDSlRePxKB
SPQUjHhORiZzH2d/PqLn8oHjUeEV10dIbgk8EsDq2pdxzVzIHbunYrnLRHVYOxtMqiGJTo012YT9
xHMMwknc20X2RtaCh+sfx4rqhYwNj/j/18prOeawTj5ofGu+5ykt01yy3fQ4jB4ROu4Ikc4EHua5
zgQRkRb6QT/IFfeEzoCidIdUY98ZIze6CzFAy/7gl+AoSdWYC7TvSL9OLu4B/RcT7VOysX06cDa+
Uq3m9Ptp1KKWrZuKKUOma8Pi0Rwrq0LTz9MII/F+i3XsspLI3P1GWHRSaephp2GeoKgrGyD71TeS
6dFnb1fKoDquPjJWkV5TZVyxSjkmLM2k45LwRBvNte3fGVxV8WIByTXTKn1+0kCWrLZBrFkfU77W
ZnpX/I94r/N+NaWF319jQOI3xdvHhd42xWwgtwvauLyLE4EeFitzXDTZjWKPdRQn+x2h+VhGQ5qu
dreOejORC6Ni2iDcI1P9Nph2dGHYckimHN3Rk4vtCOVMgDJ708nhoO+8CL6+vEJMpB5b3Fi+lmoO
AwqnNZMQNCqMDSILQOP1PW6/ewrMD61WcBJHMYi79pdmS1cc2KoNoYabXVbIhLFqRWBigTq9MBCt
J4iiZxAdLfgtSfXmuVY7cmtgJZ01nWuPDONaXkD+V1xGqZrLR1gt/TEEfZeXL+kMpphiUhRnfIxM
JWvjKceNjvLvppaGd7QyQ80eyl7WzMeqE1O1mej5PB5y0Ml+08K6Hjq90fi48KJKbcYukX3lm+at
Nk5YzVdHIN633nEOI6U00OW0Lbjz3ObEotYNqdwrYe75CYTFSkVLsHqZippMgkwDavmPLZ9X9ljw
SxiB6/TwH/DsJOIif0ZRPaWihRA3ebLR/zH4XGgbMY0thGgd5OvyAuqvm76ISEhv1n4sWc1xruZt
jiA42XDIw4pF5YFide70AgymizG3VqWdtC4ePZDzArTbyTRDTZRIUXhv7+EbMBbMHIW+8rjQ8UvC
j/wl+pp7u4am3b8btQVjD8udIM3JY7AVZyuyxfBni2Rf6M7Oh74WcV+57B/EOCBDto1M1Iqego6o
u7qMwWv84UHbURFDHkByHL7/8d6qviTuNcHU4q289hiNFkDjxcuGBcB0N6shIyF0F1fAcDowGvSz
gbFwvEw17Oq34XzppIlg4Ufq+CmTPuY4vLx0IgBKvUHFJXZHVI0dp3PVlphAta8zw9IyhY3C5qxk
aOzhG5oaoUSypr25l1Zubc7DvaqKLaGJ+yzQ+akXBYBx03o9CgpByU6QKO5ayIylngqOdlAHXqMq
bj3JTLMx+bPq1bOiyyc+3lkkcAiaDYEUdPqXboCAb9thDu7FYK3xODDytRdRejE2YUsc2pM2v1pj
EOGiVe4JDXcHI2UN62AUSgqe7EEku9pug4NH2D+cZFCRgEgV+31hFBp0ZQ+6BRGvbn/B+ZD/gfBl
T4K30/jbBsdiyCtu/S6AmM/33aDM+nK3em7jW25Q4OTsvkpOL+d9H2Zeqs+kjba8vYE9v0VTW93d
2B4WqekVkfL5/ejL7bwHk3fooxX2INRAm5nOvUt9req318EL9MRJgM/rdM6eO8QdrTrz+fCWkq/k
7CWELuW5MXzJBQimH+6Nd5lr11RNgyDXxi5z7GnFerEJ2KjH+qzcySvAMJA1L3I69O6e61G3o/4e
bu2wP1lU7blF8qwz+VONi7iGT1+PGp1U5uPuBubQQSDNH0IpQtnj5tf0FX00Hv302DlkfvHLT1uC
VOPr9dE6erA35sFibMNnODeUj+h7jCKgzpQGJD/duAxwrguJRVR5fbsVYyL6Adh6W/6NwC1O/MSs
bkcD70nVoKnPolO/UBPOp2BR/GUXv+kinDXkV74t5lkSoYpEV6PbsL18QaA5CCFZXQ4Hq6IYrtsc
YKbnfExdneGsLN/iVavITcWik8jL92rAkLDjZ61Plb34EyjE8JNvoc4Xi4V77ghA5ftFyYnfVhX7
u65MGXul6jj1aHB1NC4k8KiA6BgWlLbD/Cx7QlWOgRdXl055K9jycY1phEo+m87Lyd8GlYA0fHM4
EghkEeemncccLAtxJoZJRrWlxc60pWPSu0G7BqP7AqkNk48hfvApGS6gS5kZ4CVZLYCiw1Wixm2m
8ASSiMt87cGODYvFMqdYYJJbEWM+Fq5rTzvM/ZSOWbxDTadv0ETZiOO4o716syd2rfJKrPnqZXoG
hU4umVrBcAUPP83Z0NXS8jtlFeWNCXckFV5o1EDQ8Pd5JRZ1pnrR3YcG/UjmZlJ8WzCLTYYqQ2WP
epN8AXtGS273ofHr2Ai4RUwdF2os1mjVDi5OW1tRi7uaOEPuK1214qMBk2lG9gp7OAZG2kPfx4oK
Qsrg6m7smFAzZiI2QWVJNpl5CQnE/zQtMtDTzlYVuQmZka2oH9ttvTePP/ONoVpuaGEQVGe9Hhb7
uh1v2t8zgn/XRy7LdTtXsm2clOY0sHk5Sj3A7DDsq5Vi1hwRS3jiXb4AXs3K11PaSK//RNqvCf0s
D+0CcePS/08tk6s5idgUSqGsCZk4IWUD+Ywuc9iGiaPbmRW/ZNPGM72u7tYT++ryYb9vVzDA7jxb
KptrSD8itnkGIJjIy9pvyia0NCs5cIjcrKkjyDlff26F4V9MbbIv6bsHeqQv/VF/da8EGGM+d0eY
wbWKEwNWLKJXzBiYfL4+MjDx/fPcEaL8v4nFQVi4J/UQv79J0A+9I1ZCuEqq1tqVEpf56oJtM5yt
CxQ+0pEhuEPvFYlBZAbaBKCZWc8SUlTuALxwaoTZ+XCC6man/H/ztUW3MTFhipfAmQpfkY00/3cV
NDww3ADrgI53jG71iO5vbrVIV/6I3eQ+IEydbhwZixzn9STbqEMH9ZbuUNAnMSm9xQxKPEPCgt07
HJJg3XbF7yEQBSTbI6jceUDP5eQvhejKUGymh7Tln+UltzYkDVreVvyfYIvwOMz2+ZNg0cod8L6n
AsFGcgWm4f1xMnpPwiLxnORHutZxC1rW0bZwMfK0VAKCFgOqEDix292JshQeBOIB8s20kwmt8IP8
a7QBOBdzQwgnYdkjt5SVSnQCFHu6rH2vYH8GXGNqVJiqFjGvnOk9ga4eWXger/GNWkcJd+fuwgAN
Adc9zFZcZs7k+ourZWXrsWw8+g24OfXYNcBv877U7b48xPTcr5IXuT6mXWxNLDmF5nHnHBYG+ep5
+Mf596EGPhHSHmGdXxQ1wtCu9iD86bocmcmgeE6qhnjHqL/w9uSC5zw+rCG5hWzr/KL3iLFI1v+u
ETmpWxipfU2LJfjxxPDq0l/UBDOvXSUmUVZh3b/6UTgyUcir01oequa9zo2LNltHvg1GWox6Ez6v
V81Sai4QnsSGJ7TzgIl+Qq8Ewejc/286kdoVel+TsQfh+EDrii3G9q/CNu3WpCfitmuyeq+e7YLL
Y6B8nnIvivFqjnvZDw9/Plwqk3EpHjlqX6RLRPrWyFxE9i0upO3nACTD7n1BZg6sBxjxH0RvO2jn
5oV9OxF47Bs8HfRrcWf2c+eawsfYs6b4uePXUq1Em+bFCBd55+1gJSjbE9XVlzig3Q4CG69Y8YdT
YmlWwZrVDnNB2oilsfKGY1gz9fMEhJGmSkBhCKJo++Y+k9/3yC3eKvqTnM8C9QbqkXC5pxA3xRQo
6ZeYolliltpPAl2vtU0xkz4JDNLkiWJ1p4ZVqKr2XafuUVLGfXP0amufpMtSNF8BT6JoIltFs6uN
KDtIdnha7eZvTtWaiHOEnHuZnWmpX7tRdPz1tWGt109RGzBJGf/4ZOphuYyChO4BMaqY7Te1xafY
GJ6bo0fjJQetUdg+YG2icdEcdnXO1UftEf2MXTpM/S9hQcGkT8kMqalvdEZTW6bBKcB35yKbc3ih
sQwY6TGoEGfFxbTGDSHyqNcHslZIWC8yEaCb8q3wUTm0TQkXxZhjS38j6xym/yiwOC+wd/ue5BS0
04Pcn1Oorp/vS9HqDoJnWAbURs2nJaELnF5UhIYOsadFKpFtqi2tSZUs/NxBJ7EEUhaoyx1gmEYv
YgW0GShy6HtAioxaCAbaYyg1VP/k5CQbllvD9UVAaxle9PL7yQpLuGaa/FW40UrVfC7Gs0iX+7d2
ao6lUaXrmC7PBSSXr4QBRoFx5pm/s8xFOjLo6X7197oxlpkQqWeYUXg6g0NwnuxIRv8zFNBJzxar
oo4XRu1jOuQ4qRzmOtgBFeZA6eECOYTNy8oqMBmjcVeI4xlXQ5LN3ReKmqHk4vDhQVQeVRLJVIoV
Tjb2yKf2fXEbhkxagvjXWXWba5uT5uFqsAGdZJ3jsXdWycRTt9x7Z5RGfuD4njrX3pfP5v4kcQjO
VDmgB3XBoWtSu1BCFvbkWGXq67SP2lCY5pmX3bEk5uObicOQ487ZVPZIhGPR5Zx5dkre6Rkg2+es
ze1o+uAQLanY3QqTzmG3/uIRS/zMjgb13VSAdtFycZSBRB7xU78bwZUKYh1+PH7PPOwUYK21Cd1k
ZJ2eXAxyLWe8zEHr6J1QEQmZgc4EvLXqsn1uj8uyFC0Tv3cuBfxMpqyeoBAfIk9qRjCz0PC2hQ9q
wKy591iRMCAL3zdLbCN2eMN4uWM03/2p6iNZAQWdJlNwtiJ9kmDkNwRnxg0ag5SQ64xJEdOZ1yU6
qb9IAq+btZJUNluVp711MaA8DO8Xwp67F7B7SjlQg+LaC9p+vV24qfxczQ+LnoVUYBESK+fpL0RV
ymKNvP2WhasN8fPlrTtfmHYJeEVhLub/LrTp0xlctJYnBBX1v5D9NbSveGCV+rbYqOmZ53pVdlVG
98xebEhYXgWT5DHh0aNVpwl5KBBiFQmwwYUHnwaZDdyjdgnQ0FdIvCG36JQxISFpdwikB4VOXx+y
Rkh+1AhbYamMAvFNPj5aD5UXRujWGCkJzOcPSCOPzoBus7wFVHSohFkZbuoFjmBtatv4uCNodS4P
NYraeXIvdF9HHwMyn3nEVNqMMYQBDCSExIeVn7/p0LQUev9oNuHHwpVxupvu5mCii+M4eJIZ7FNd
YBz2waK0gklVkO+l0dtlkghBdXzQetMRCZcaO1ZRIhVBzN9AL8LYyhDOyz95AbWvefF1xjLfkMII
TxFYDCudaNnl9Qx6IeUr/f7cRlxN20FDjWz6bwXrcRHqn7eI9vvgVpE1WtzViEHLO3BW3XYCOx1b
xb72NA1jzIA4aWS82eW24Lp0odP3406Mg9v2EZg7DnMGFSDEQN6vD/yDmN5mhqa7Q3d86PwD4lLa
Eno5eGSuspCkX9bKaPT/6idg3Eh0pJWxq06QGo/c/RSjvZDgnVrUDcq3zECfdw/1VH63jTXXetSZ
k1DJlNFmRShdgvDbhdxBlNJd6xsuh3OTMZV2d1W0WJNOpqAty7/qKwGN0mMdKqBB3v9SES4epQVB
5dUiFL3s3b7goy9Nm6MGRQYOxn71xFvw9CeO1gCZtxKNWpHeaHwMQhg5GPVSazrW0zsv778uHhh5
dXEyiLGExBMGckfstjmUt1Kjrz8RToknZ1oc/mIMSWysGBWyX0ZLhqNcUpeLXECn/sKqf4HNENl0
O/oYzKn54qwjLqGGklPs1I1/BGKzms5xCEQt4uDzmGw14SqPSoVDFmlI0J7AJFx+tM++yqckGCsH
kWn2jkyGBwnwtWiJnqLJ8S68tmP13iFUUz6WC9LS+BvpCl5refucv3YPEYiKpfAEajrtn6MsJMl6
cLy81PpAKLBdfqCEQMcLQ5W0E9sSP+T8Ge1tawUxlcwaKtfvXfTu0JgFeqqGG5TJ0xdhG+CoFJJw
/VkHXeTmI5HaC5Nh0WAl0LLYbXAG7Jhwq8GgjQj1bt2qc+iDR4RAmveGrFHuOP2Gy3iRVuLwl9kK
sDMK0KEvMPGurpc/S4oE1miFubtjcyAmOADNSx+WUsFQXQ1eL11hFRGTfUKzzjs0AD+HMEnW/4eA
4PpA58JrZ6nJZHZrcJ93SBSZh2/8pj3s5KOIebOHkzsdP7MUIPMNnmcPtzpV3MQ9EZtYzvo7t5Bf
VL6ml68TePCwvNvpSrxxBfLpr+yRHEL+8vej8hRGw5a83ifW6kuBfAzxbcB+WOd+0Tba9zluWxoZ
wha4QyGahLnwxLJiafxg6u7TXQrK3A6u62a0KBSyKvaB7Eq8ASo2Pxt5QWHio4aVqMSQwqce4t3s
LUzcm0qUAAGYrj06J4/8c5L5T5pUUAm7n/zT/SOeQDBPD90FAhTGf7GHN5xx3AkyFtKfrwjceos7
D3zPbnduxdsrCIzRwbn7qQquz5/qDQTDgUCZ27y9Av/o+dSXUtcDVKhLXOP6oeHIM/IH+ssUzw9k
ZdYL/AG6uuD8RHIsWBChxui8dyMPxQHIgZqU94kZYwCnGlUiFRZIHZENJrePpDeG80aaI8o2elRZ
j/zv32zHGM1MY2JXL9RCBjVshbPLgqUJsYl3+043am4b1JLCozezka4qxze6i9jdcnE+MU0++qQp
tSM/GzNYiyTvG01Ko6S8XcwEo5Y8Hvf0NZXAHV4+2V3ASwIPIgrt9nZeCKDvzdpf+9WHsGAVLcQT
0XdrmnOA23MGSXxgusurVJO+51r/9ZtKGLwN0nZ+hHKUH6PNjYj3j075/NWseRA5rqbZ6MJDMIny
VPf1ZABv6wTIwmaGVQcX3A9lRQ7jtEGRQqQoaQAupLQL0uC+MceBVYBmkhw1AZmxvsb50SFjGeju
fB2KXmqRyVpYLoopT35JBR0T20xccxr4r/al3aBC4H1MRqmA5org8nMS5DfssDhcT3Kdm4D16PWy
5tteRu0l8hZ13GU2OyvIEH4MPZYQ4AEilsKeObOG7zDk0wfcDTm3B/7Zes1FCSxzQ1b2fh8P+DsU
BB+TmkCpcFNEn257xl/yPCeN5xJ/NnxIU2BmctfYErGsh+i50+BtDBVofC8G3WDBUp2nUQ8CGV5U
DcDzKat2XqDiPZCAn7kmwRHqAubrv2kzlGQjGHKtmSl+5yC2IHtil7m7fonc4jrlNg9jLWZxufvU
zsyYgdkxLjr+SsYMEOoLySI2+sGSuUQlsBWovaL5x6F8aKaVGJPrGsBO78mRHqfBcUA7O3rGcmMh
XfK04rKQr4Dpi/JwtiC2MRjpZBFCykiYheVrRvG/R7ts0BjgkUa9J0KUmloUz6UZLDjZnyCI9fnp
YMFAf0DJ42zh+xKoHzUgBFWh1Re2wPY3zAq5ISJJN6SL408owNJXNkptb15AE7vqyNCudMg7qKBV
RcKRnLqhJSCcICKnQp5atFY2JblT+84GbKTlfUXdOukK/QxyNi7FcRVUkAhO0mmFscSGmgRRgTnj
Rh+GwbGr+VyJWm3M+1HUacj7vOM5BZ6kCxjZPvEFpLkKPPS8GU01zGCi2bgbz2HRkEaWqbYYs7VL
7hUY8KHQubLRuhcrKxA+7IdAcqbJk9kbuqyVPlcA1hnnQrL+Skh+oeO8bWk+4Y93SUpe5vB+nsGD
9r6D7WaEUPaoP4BMrOyEvmQ9xw0WLG1pPwnzRLBxWBcLtB+FU4+etdTSW2k3Iv6aKgKU2vhu+N3W
b1UWOculJ1KTJvZe8/TIzRFQSSfumZHqtGHOO2ewKFtsMUJCHOO+mnxJ5REZV765qwwsff/ybrMw
uspYn+Vtu3IW2XVhIolAfiofjq4KOIHMbcnnp+JEGpDGW4KSkIMNB6T76z/yr5o8pXm74Ye3C8Rb
d+ffMh3ok5pnrMLpN4FGh7TJHIhDItAvhl8dnOVMbpoE/3h1+BkY+zl0B55AMH6Bm9NZY8kaMHK3
g7/HvHVfXuvQC5akhLWuuxo4TKFDMN0tJX9N+y7Q1wUQ6QKKq3S+otcpeE9uGiA2bh8hnjmwpfVt
YchzP3bQ9xLz7sZjF4XiagXPdUGqd3iKhIsjeK1cuWbXOq8FBmZptpaooDq6scJksukx8VAz2zhn
Gx/CKM5dpZhVo+HMrXzOAhX1LTPYQztXknHotes+s/9pTtGu3IBzkszC/vfH7fWoiLUa2mAM67ZX
g6bfMpv69Yj32eAsJugGdDjL1JN2RqFPtttf0IN1mdQVJBoMrqQKE7D1JPBuexn1w/zi/YIRYDXP
lfg+PmsmN5nA4N54e8mSG+m3hCa6s6odTw0EhiUnzWFlvezNmKp5Z8tc0YqDZT9CWXdhH76b5eds
cid3Tvm7L5VJbV0xu92hlQWfBg+KJsiXEJMJEVO/JFnVPslq7MlEOJojhlwEIT3Smn3jYPpYek9S
9W3j+0KXeLJzrXzUvw3wM9M3RrXVrhd3IbzSsBijokcOINuR8sVGxitvBjsb7Yi8ZKefwCleq1fn
YVB8ENTUDC1K4qjkS3LKKNJrd4maR7ERRAY3rEnbkDZcXFhEJ0wdHNxoTpZ/iDFR1GhFywk8P6qD
d61wLZiMQeQ3iggBeg7E/Ndsxwlb4ZdmOHSKGfcXdi4Qzai781JKiqgzdfemMKjCKp7AxTDJOcCC
DKlYYPcLtZN2lcw81G193LSwpllylGMCLB3//9SapcBfTIDcF5ApeuwLxhSPqMr/cyvqmBp9WzF3
lm3hhO+laJodJFw8ox7G0/1qs53q2Oz/x76DgBySSzaJQbJcWl7s350Ajcum+W/gpMucd4F0CB09
yXO0LD42X9L3PSK5kZcGzyvV6CFEGE53ivyffqWRL9rZ0tXjlfXEV+UPQzERtAySU68UOzJg4iX7
SFamQyqcsBUgIfd8/rWMckkH2mb0qIZemzmZStvFbaWGHaj5Pa2soTTWrwlDvKHhqWpw3AU8dbDT
QSIjXbpHzJNZBZYpm9O4dqpi8eIKii8T28Dah5Al+oIJhLLRRRZTga5noFoa2mS/5qRS/lgL7t/f
U8q4Yfyi1jPQxxD4CQbJowymKVhPOxRBgmXkIZKtsGu7FmhH4ZveAb/wgxWWF1lD+QnfY0eCDimo
b1PBRiaIOITX07y6JHiop0as7MTXsIUDxa0nThhn3auBuWMD9oQTlAvSj6S7uhnGRef7xer3dFh7
99/1yBbwfC5m2zNy4hX+MUW4d9HM30YcPf6COZaBtdlY5fuf97+X4bCDbsMVWbb/SerUsWnuMnlg
gn/Z3OyFnmBp3FZHT120/OfB+WDNGTWobQz2ZG1mzKU9T6klFlMxZPgUEpucU7cK8iWmAT1Z5IiB
kWJuV7eTHMDxNvH3aekNRcmnBnXMwTFaIgComUM9bwYXOuo+zqJjWpcDAMWu/JqJnKwvNYlXgmKq
eoyVXLiRqRj0khd3y/cR6YOE47XKCx5hhWB4vSfEyefcm0pfequLZLyP4PAIDodESDgCPCi2ytjP
nLVowc9YoM1VS05lKTLlCBRNn+s40y2ZARaoyK3nzsftsa4Uqt0hgi4kClrqDEbzmXBNDmkEHuob
zTcCeE74HTY83ol+lPVFU7mzmx5iH1CPl7+sVolV0JmEGOPuGZ5bZD2JbMREuolRRXYDPBIWowrF
XdJah4Hw191e0RUjIhup5GoSNe68DtkYUYuFy5YvHTEhtNr0aVRo8n+0YytcV6B6iRF7VnNs27bP
UZXg5B0gMIqn2Zybg/pM+M5B+Ru47fghM7MDcmtbCueuGdJWOjDmwBqNGIgTbEwixK4G/iyw0y+1
DMYPxBbftDryV9dvwDfbNZaDgO+2PiT9yQA0ZCUQAdwYGdamg3TOD3u0+in6rgJLuKlRtdtTxcqM
VRjwll+oVqIf9Gys+F1o7GkIvc3j5CeyqKhS4E6WBs757jcqqH6LOO5lTVFIOaYt03W9KfJoIMVl
k/ntrckdWZgU7fk7rUKCFEyUolk/UDiQXXEOUToqZSfVrk7z/uTWT+cSD5XzYNfNNaLwGLexeNZM
sSyaglmqBul9ZtY39pyr38nV7SbTs6Bt2Z+bI3udMfgRKcWWvse3qMHPW1KAAXtEXUoP8KszbSoY
eysuEEosrYY9OiM1wIVzyCTgnJB2yWyVd0RD3p2mgv86ZjHg2icPHYWfc4qrCqfDf5JJemuL9XM+
IUtsTAtl2QpNpAs7LeqdcEc6UERy7m8Y2trL5j4bq+y0jrH7Zb9Pbkysa6r0tP3yGkdxvhjDU9xk
IfEPzqrSxapV6bdfCOONcWvEUORnCc+BM9TqYuJ+A6IxFNdv3Jmm4VyDMITN+73EiqpCnba0fOfi
17fNsqlDFHmcKh4v8HWyV1uXe0NmfceGAb/AelKFQRUPLHOQZ6FtndbgiPCZBOv+ktu3Z6CiQKDS
hSO61kWHg8I8dnjzYs8GSbwTeUocTU63YI/mKpTAlYtD2N1nucKAvvJ6/3ABaF3sVtOESDipMx7n
/Jz5KNol2B0sYkd8FqyURXh56nigMoqzodt3He706Io5YsJpzGGGSBT6xlNONp+kfR/luewMnf29
EVmXq5jYjqA6NSHbUYFpd+g1a1e9L2sklOnqt09DzXKk1DBfIQGrsyxDXNbwy9JbDpLXDA43Unwb
DS8xjXAmMLiWujJ0WohPuDnAekaVpHU3hbWD1PiqS6yRIFf4m86TJaGGQrurrxw87PAUKq286gCE
K3k6GpdmSD443DSBOTNHL9CGcu+8mcl/Xe20PsIQxN6xrjl9LnnwJV2AFGl/GS0+FSL1A0aaysCp
sjPiG5o9wgT+5yw4lY8qPsLop9zpfaaDOrOG5QgiBTNdjHW4CMITlOIwgvAT2X4Zb8n9PJhuvTnw
zmR1+zeMeETd4heTUiW1ZNqr59MQcses2FxHql+uXvBfWJv6t8z2cpwv8cI2u54szWqkOqDNl50l
cgv3l94C6tp9J+pCvcjhjjNNgWw7+38rJKCRmoIFKNcrgwXTp4OGL12n6R+WXfNT9QEEDVaRFQ2c
MyfmqgA29oEWWPF79M/LZQvcojP7AIbePIzAg2Wekp51dtzWoOeuDNAjg3gYpVkcTDJD8O2mk0R8
B0nYpQMI8ozsYFpCZGsaQuPEou24z0MM4qMEOt01mnKOeHwcB3d6DZXKJJCCxymiB0dDXCrbOfeR
85W1BvJ3jW1kVu/TnVAe2YzuEEfy5khTOXmlw7ycuaJPSGTZpgR/tAP8QNSUcJTX6X4+NFYeM6qB
cBfpH5M8l0ovUtPu0SHlvb2SwGjpwfrT7Jowo5D2LfA8FFqq3AKnEcL7nPuFvtQTfjxx+r17PWLg
Mx4rrNf/8U8kUeXU0UAMv3Yc/ax+Yh5cM4Jc+HYvZ4PTSwMlY48/A7qW0xJ1VTYBETovFBLSJWNJ
WH+UzwVvkZ+5kVtdKmPfBjev5791WLztEnwSXEdz78eVE/ujp+nS1BQfej6D4Jv34wzYaUppP1LR
mLZnHtj+lbLvo2c9weglkfFNZLT5/RPMSajX/oM7Rd+4MhtMWbjLZOqSkoHvHgVeyUD6GRuDHinv
JVd9oU1RRsDpg3Mh/PGj+Dt7aYm4pLkaAPej2P+6qZSg+x7ZE0lQrtww2ed111NHzqYlllFSmgt7
KGLWK4jBSG2q/jUD0WVW02+/yjeYKfd83Ib1pTkWwqg2MYRc9tqbXXYH2oarowPSCJtqk6oJo8Yk
EwHIFROsgJdT9TR0eFSX/ntzg5N17R8y7luziy5a/unrEZCPFbpD/dYGpLDbfWyafY2puloeV+kf
Gj85Tkph5PWbeA1aRKVoQMDQkHgz2wumQwtIR3PEEx6zEP3mSBS58OnAcFhq0tXglqpwI6lmDOjy
hz/N2Dd0YRUvtF1fN3d4rg5Af3kh0RTOBty2YI5B4L+Q/B5P25C/gfAYPsF0OAAfZoyWUV3ELp8z
1Y134PHDswI3mIQa5QpKJSSORYVBVp6gjulAyUc0dN5MbI77P1/TXJpKyGO4EEAyqc1lHOOswH2x
befyKFkWgKx9j5aMr9s6OOtvsIet5dZqbtHYJkRt7SSXMtnT8mkygYQF/kmFbor4xF1pkwqVQ3jY
iKXOoBwUKziW+0M7YPgwC3n9GWrz+dZ2gUdFbHxyW5bZS0ZWzzfEZR37B+DI+Ua8GqrlK05E/atk
SvfV0idFKgQcvlYZJ/tzHUpS1mp2yHayOLL62QJTaVyCtCFdzGrjBKcL26QFX8dMHbWSqoO8cOuA
tB4XEaaokQuZ9/CjwvOgb+/UWh8l8jZ+pfFq6+dlFWgkHBUtiy55UZIZPg4dRx9Ts6Si2/0sdEn/
NaRbOZzXJebLw/bKXvQaD7+K+5IirnwJBVJLxO9OReTB29+tRXW/wRv+hut4oTDETA7c1xHtcjhH
70Q6m8FeDlejsXy0IIw/QocOp8F45uWCRySQzDfW8WH8YitkeaZKlmPGB9EsC3eaCvEhdOAsEpyZ
Y9AWd+vprD/nwH8FAJgzVkxHPs7SkjFV3nE8bWDCb+fIvix5SFycfBsweisND9fVFDU9E2qnUcdd
64EJ5fcUuQc2u8HH5crwY8C1HV6cHT3dAEYHCPI3VGFwNqsW1va8R5lAD6DJ557m8RwTC1uQmheE
jz8dZHb8xpy78DMlcqcD2M7Vw2m6RAKx43pH73fiGtGBfq3lT8mhFOqA5TzVi6zf8bsOPNfeWpVv
onExA6gJp0Q5tFweSnBQxmZ2Yv8dshQ2CxE6VErlqQzOy1saEzdZZ4W6vEEUMqULPmiU16HWEQ9I
2SZaUnM8kNyjSvcfyubNSRvqyF9mcZyRkCUcHPWh+Y/FDX6z9WgRCjNweIitC3qvoHySG/o6kEqM
qKbrjkH3InJXhbZ2EPPnQGwW8NTGHo0yq9s6yGiMF3tgui/hs4w8yEbv+C8xqp0Xgv2Zw0uC6G5+
Nddvm/K0DE3hN0Sya3/42TXotIWd0xfW01OiFDMcqE0dRbKfyfPOO3y06H7wkR9CI5wUTrP0M3IM
R8kH80avt/iXQbfKJE21EvTNDdfOChVyuZbywKxLvJbF85vRCbflxYUbpYeW2l7R9BWnqR5eEglA
uWDrGWYLnhjlGDn7PDww2/Agz8PUSa2GPf12djA/EJ56xHvvsZL8URzjAOGF6tsRywZEri4cgBT9
xarFXt5iP/8gONSVouxf6yolqTgCs9nHjv5uMIBscOvgber4OeB/NYuaWMFBItaZJVc0MNbTtSTz
yAuXuMQ1LbEk23WFzkhcQ4EtCjyAzg7Djc7TQLJJdoDstSgfMxeBB9/UrJolKEZ0bMkdq0t2PVFc
sqafBVkS2EMBpckDXnKgt0BZQlejlcw4L+22vj9xHgiqBP5IG/O9OX6deNhpRJTACP9xBV5Rh9D4
SQfmHRXhN1/WXoA52NPUyW7Mj5pQgwciP3rX13FhYMVcTbINb/+JWwP6arBIjwk+BqmM/EhAvs5K
Oho7HTMNaJBVx6PN2m/hZTo5U0v+bUj7y/pHYftzW9ENw0VMD+6gPzjD0NIkdK3CaxmXOKEQJ0Es
JwiamLkGnxCu/CtJ2j6uU/ZKuoK18mzoClP9ehtvmeOS6pXhBdyMLfWk0Vgg+oWkoR1yHnQViTEd
YBYjFRWQmzihlZSpvtoISxBC1pMQXIkG9T4bD5CAsIslYPWVj55Brx/lWvVh5I5dPA7IbQbRJBaJ
pc/Bk9qbr+i54+Ec5G+vId+2y92kE9WZV0gQG9qMi7r8e2g3TwyfHmZc4MGpRrjn7pSwpI1nZKwI
7RAb0eiNmJp6ydHYGqk+GLd4RyTzVP6vnvQ7ATZAycHNDpj5hvH125r4iQhvO+JO63QZCSC2wJ+S
APTSXuHI8gTQCKdRaWTP7aQ5ulDlb/w+7AgSM+d/+mmt5Ug9hJzAj2vEh6ljP6ey0CG2WUKvBBCm
TWy0SDyR56DrwnaTNafk7qbsw19RDDfixEZ549bF+4DqgL9Cvz6YXuOY1h8uQTYfflyEWJqrfZ8l
Xdja3Av42Ik+2GYWORxnYhpRhH91tRpxanSL66MmXhxssHSC9adA3Uhw/eZ0meJy5WVKS7LvmdMH
rALEjevAaDmlz6W0vgMx2W/4n3SPjAodXiWoWSEfbJdPMxH9wUDrUwfshekTEjlsrx6t42qKAkcs
bwrKHAEdPZQuvBZRaHfxpugpoGShlE/yKtKKRp6wOLuyie2+RqowfAJES9HhsKh7mc8X8+hmWlc4
ECqGFrvtM3aC089P+K8L2EJmo10KhCe/gqAdaLMRPSKhb/usepP3DgccSbMugB1u3knD6/ZudwdF
kPKWkdkNT/gWMX2IvbqRzSvw7QTvy/QU/0b0ym0knr/gyQ8Brizjrm7gjxRwy2nkqf/vOPk5+lOU
pMJp8N6YAbV1HFbut/MCwj/fomxYiNF7sxweok7PAZTYctM1z47anYAhQVpSii+MwaO3iOYKT/9E
+64xIsgfErnmgxCS4foQGsPDm80Jp8n0S3sLRzdA1YRMaDNLAMwYFvChX7j9EbBCXsoXD91B7sF4
lxqL9QC0M+NQF6qidjKmubjPDtaCLmgg6dkziQW/FWq1YsjDg1AqVxue8DPsCreeU0ohTAzB9lUA
I1xso/vd8qv5iRyqK4qLmyg77APHcxnvmkdzk/MT07VdJca/BZ4GDz0pn7t75/p/hb19a3SgC9gY
ax/pbmeGJiPHlGOm/Ob92lZEfOg3/j5JUjXACtzj69U642KzZrTFHh+MCU07GduzSTkMsEb4+FKQ
z67ClrMNk16YD0gkDO9b8nlDbjSuYf1PLCOroF+el2gSuOBB+3WfOqPaXnM6+5lF673ee8bbN309
KJaP2VQ0AO4qrwwwEgoPS5sTZTHOMF/wwaNYcR36FssbkVG3UuOEAnsA6vVVJ26mF+/C0hOq41m7
QiOb4CKyue/nP45NUxVfPfXGpdwH+4Nl9mv1pmYD4F/PeC4TQva+iPHmXYNAzWO9t6lyqSrfPd+v
w78lXLghThRXtZrhJd0O2LXTWlwj8HelEWmN30AOHKijOsxcGgu699nQxDHXmhhmXcxUwC1pin3y
2Hm4w6ySei93xmfLTSOsrpXmvIIDsiUBiUkag1FT+ZXVz0at7xbkINgkCX3RijgkUBP3PegRwBwB
6XADwJ3v2tX/grvW0CaT/qF78ufG7+ftcHHubpGzw38gnxHlIeByoX4vdztxVKy3YyZY1UydLmw5
0OXrLtR5djJNIWpteh7OdyNVNYs/SMdqGAYetcQBkYttoI9+B03Lo+WUKWL31l0azfYsjZ0HPtDj
8Om2tumWbCiVHMWJ0wmBZpZSJHMH+fSWpMmvC+LJdzDm1adqOij1BiHwV3AlBv8G0/Lkn/KCi2Aa
dNIYkPaqe/Qj0spZxOiA8EYxHHQbU2TVGBxlewHTeUhZcf9qRiu8aqRhE4G0KlddPSXRdLHlhi/m
CvGY31RwLSvTzHi6MDdIrTum0krA4Q/R+HMw022nECY9xJuJah35u9nEBmrZjDZqIzCk6b/FbvYY
4dDEw7diKkvhozyDjv0o4yqcGlly12VC/hmJl4lzqvny9bFwveAxc7nMdhJKMOTA44t6Um2eEvoR
SZ6uVpadnmubzXmXcRcnfoCivPWBOUEBSq6NTBGJZOIrEiQHyjAaZVQZ3D9RWN25n8gMjsTFmRyo
RMJ2glJNiy95pZVHG202RNUvZeMT4pY5An0soEeSmqzLK/AaMBV3EqoC4j9WOFco3HvKkTdmtzW5
Gep6xa1xYvNYHHp62btcDvF7Is3n2hM02K0456Tqr/GP8es5zHr02+XuRuCm9QGkFmxKjURX+MH/
iaB6Au27zlO4ROh9/fL0rmYnFDQa3wvZTQYn7JwpchmJPvT3htx1bOVIymAZ5aa63LklDG3CG4GL
cpzYMkeFl2hSckoJtaVTplZPQJatVBqgJ3+sWl9j9PDTyvYXiYCpkm0flgdRTvDohZ55c9KCSNEx
p7t/AfBp9l7oAcgF61dWnjdQXIHEOopkJ5BjHo+fB419Zm1s9diGWOq+LpCNtZhAWxmmVIm3kdvo
DoUYYRqpUJ9tRDLdMA1X3hKTiZCAGTAhEtfepq40Z5nv2Q5eGCd2YuA1WvaC2e/5QUNGItEGE4Bp
QSJyNxxzWe/oO58v1pqrucqWutlZBRUDvh6IW/ff8X/S8tWS/sLef1bkKS3Kjuq8SGcKX3wQv0Ro
QjTEqoW/erl5KqYndgwQgvjZipW7tvlqJpxgYTV6lx7tSuJjh6KH7gGsVcSuwiN67lOB9E9mNR/L
/n8RUttQ8Y3UOprgZyrLCiBbJ00T0bfbRF0LPNl2Pl5lNjKDiR7YKy/M7zMNJ+8N+Y41z6PglfRM
Dy/FU/EeifkNetwODGX/cgqrXsJR33KUuesvDhcrwy86wDtFES2NpLvdxghyWErNttrIBByBUceE
ZT8yAAbmK/WOJCzbamsq/QW06waOx9fcLyYiSqnrucgTXvNN5RH4FC3kAyky4vq26M84r+X/tg4V
RWcrwjqj9fbG5eDvvCHU86CNIuN5OnGDIHhbr6nCegLaXwPqQa8PvIFh9GGROe8ZxdQzHMapS9fs
1y3la/64SNCLyztof32dyWUMb8t4clpabVHVn3JlcD+RCZ3Eat7B5UrZKv4ML16hZqqLg3DLdyBU
cBbVZqnlB7WnX9YkmP1IFqNNyxpeFdUFGOXSGcVqmewDdsxY93v1EbKLi/Bt9nBiBs/FLXHRBlyd
RKEWn6uWWCCJA4vcbKKu8QWw5/mWx4/FDnRkFgiy8xJnwXK+qSyH9MbmN4UzxxFCVptG4I076ZNm
tG/6/fpOXXnAOw2AYrPtTcG39v8thOLnVKGgdmdIL6kH0SDr+GEp1TCRuG9tZWmXbIxKVTL2c3Nm
oD4V3mdLsCakJFUEI3JX+SCdYGMjV34qkec26XPqmP1mQW2jtZchW7uXFBZWs0+CEX1rfUfKhBZL
gk+vY9Bx+AT0/hqFDXwdgaSedAh0901mvs8EmTIpYlRKzKC+h8Bx+coAzB9HcJfhR7Yp6lsMTcmH
GsfNiz1Iz/BE7fgcCtG1CFmzXnUXAuyUBEbw8U3sOi+FGbLJ3fp9yYYWihwB1IqSdNFhWg3zLyiE
EjvOav3l/Y/hiQbcQCuky7CgqpVpii31XUkFpS606GYX4JVQToO6zFDnn5s5l8AInG6hBeClvtq+
WjQDqiFYqQXJk5KZBW2pqyNKJZ6skDhOUAcIm16HGj6mUwzdV7DhbDyBLYwA++OhuP+bwmfVf3VZ
zX8o4Z8NsK218WlEBf3W1uP9/DWM//M3Nn7h9yqRCxox8THE4Dtnj2ZNCJ/oveJpZgo2ReHSpZNC
px7zVYRVxA1Fj9NO492DXZpP2hnXHyJ0t770eEF2g98j35IiG7NQwhpYjnYExcmaJo06lSwqzKw5
1oTrx6fpD49yXf7X6+8QhtMjb/2TZx+ESHnH3l0uZpViC51jNfRYtGqq0ShXgVNheWNTaf3WmZpu
0X9jDERQm24qnEc8EEHn6VvNqTlwLWMAAudfNMnqWBLSRUdcZ5DGcuMuCEdPBi8WNfdkBp0M7BUz
OXXxz3QfGiYrDKyqqC+Gt62VFV6odPajT3Ginxdu3e6GKllPFulavjtyQi6TH14js+fReakP7YkR
vd3AR+WxpW8B009gayZQ0EcyxESpI+DPZ+zQvlUHhD7+BNLzC8/YdFOkzYYqZQFiu6BHcWBCa/US
WpyDEtdCrb41kZaVaIvRRFLc/y2wNcoIYiK2U9nDXE2bf3aduDH+bKlgYUxefXdrTQnhc7I76ZGm
sTFUNM8UeRe/fwqpG3DwGGJyjIYwSBxd+emT11AYqNUmVmm8FZTYF5ljUx+eeKDP3+58yO8OHx0D
XtETHDVXWOTidvsT8UY+ZMJMuqMMtfsy2uDs+MlCq+V6Bwroi2XCIMr2iZXR1mim2Ku2j/0FfGbz
vcV8W3SHHeH9tYA+Wg/vTuA7eaKa+UsnOhlt078BzKBFkZy/pl2fOuxVR92wKcj4i2ZPHkaGvSvZ
RTLXLM21XXIxHOWwH5y2kfqBBovvB1hy6M5Km92ndmPFSZv/+RW6OFDvQYeLFyroCI9JttHlbfo1
GN/i4fn2PwdJDGcaW+JS4W7EGoJoNM7qXCUPIQsPT+OhK7DQaCDsoIq/qSzuZB/wGDPGiAFcXHsn
qXYa3yGUBPvVU/5isyme73ZttDDtJnCqFI+6ygPOQm9ec0IvwJgdG3NoAd0H4NcNAUlRwnMdXVL8
nVXdRDHapCcOsX1/4bYs71bxXOEei1b3u0fG8a+D/rs+e0z/sHde8NK76f7Ko7JXav1GDSxl+ftW
fyTIonhRieaw6/irs6lZQjzCgjyEkRRYF3aqavUYebRMtHuN7d0+ZCbGXdEsqagesnYzASpIQil1
zvFoaqp9l0+HGUMcHaImKwP3uD03dzsZHP6i2L8LQSxDhLoZ8hjtLI2HYQPmTD8m/VN1R6JtkmVE
EFu90dwScSzZ5ksRDAet5pjyvex4ryW4AHoKMiUIP+WEAm//df5+MMwwUbKKXZ/Pjm0WUh+wIPjU
Cb3j7k1AVY7/6+ZmYOiRV8LnBgu5OGJEU5GE+kSRVuBq2d+va+CocYYDCvN/yHemYcar/v1eu1ad
I2+ro6sRWqi1nLLoeOuBwoHhnygRxFNHhNlvV5XNL9FZmFGAHDp0ExRoASeIE6SWNegpwaCn4Y8/
ewRTm2HUlfXWU7BtgVkfrLNS6Lt65etSb6an1Wl3S5i+Ua1yVreQSt1ELFh7I6XDRsm0FMo2vvvU
eFCyVdIMaDkXXxz27FZNUotsKcuFAzA9/x5cXtOIcdUZaJa5iVlsKzEdw8dTq9npBkpVZURJEPic
xRPD/kA6MD2TUOxwxG2750ZX0l7tVw60LaYNBEucDT3XFFm7gIyj1d6ZM2ybDLZykDjpaDoZWRx4
I785rFiw/rK1xPr5nXVL4de5EenM13zEmXayVn8Fp7JKrdycytfc9DbDKp1rugo5Coh1GPEBi0GD
PaGvGtR+eI4yWhPWfB1MsVOY5QJPSAngdkIYA4dYuqjI1e3bvt/iHLQmEXFrjItZq3oD1R1CA7ad
fnMZl26ziOTxGR9PGSfRRApFBYERT9SmIGH4CCR0t8BN8R0NrQzi4Wuj50yHOe9bBqersqIDzJOa
RKXThViVZUrSUugcLWVnSIrGsGCP3skNHl691rh4wBulpffHEvOAGzmEYfAfhD33zbFewTUUZp9U
J8IYg8Fo5zJpliu7rYm/5qqgLR2GyJ2DLY/OUYgM7qwYbgaUAX1oj4PtikpxnBQDjEjGEZ2H8+aF
P0ZtWbfBujjp/QfLZG0VEncBqc5VIKTre5/sLEtQ3WEsPa2o4sJq02Q1BjFs8uALPyXGn5tqXc8i
ecFxtzIc9EYl2LJJwec/M59DcixoCsK0AAKjL7HTB7/tBWXgZVOyiDz7xsM2MR4jQIsgMnMx4rYJ
uXhiM9lNm53U81zETIZAdFXnUZW/2rVIQfCmCRAty/4ZzNo+DalJedId2gIiM4sEsTZD5Xm+0gD8
YNT1FdcQJPiBNK4J8NWBg88Yhnvz8y6fjzeaQWJ6ul22eJ4VQJSWTzl+d06c96wu5qTfQsOuXmiH
/PGZybts+ODHAi6APyYWB3LLDnbbEgkIAL5tU2Q5eEm5g8uEiWB5lxthbfg4i9XzpaG18rPFdTvX
B+7TLnEAZcSInCUBLDt4hv+rhhJv/7XpUkNfe5Ow/GsnPB/8x17WBrYJxeWh70M/IPanHBvC1Aps
WeoL2l2sUJyA6kR+XWAvbGyOz8co17kQLPOHSkT2YEgZsSbR+TkVAF+iS/uZc+Qp+gLYWP+TUI6c
5caDg77+THAb2nTMsMIpctmigdDH9lH9dWsPurUuwPfoxDmsjc6govvtu8B79K+DwXRNo+bvq/Ar
fKtfEDzSC5dFU44JneOR0+mx/ZgNj9Mt1pZb3iz7pfN6BH/UaXtA+P4Gu9Zv32Ybow0/fXFPxHhr
mbx18OCoFwAa1eFco1kek3CrDM+FYgWzIb9YFDdaljE0CTlZrTmN0yOlIxnNm4lq7z16T++fLTDV
yqr7pP3oQOLWIbeja3hx3b+pi6XWV78gz6gWMYH1L/V9eoGZL0VPYuT3U9DFuj1xfFEt2PNk39CU
UlXHTZNpjxhdJQ4h81F9nFyxujZsan+giS3elTiHCp8D31Q5RrDR3Ss4v3A7LXVBaf84kF/q++VE
AMtFWVJToQkICK9m4idbOpsN48Ue0zcUvQfvK7cC3MYnQHpf5u3I7GpOJVqr6U8GKP0uuMSb+sS9
pVTl/atLn9Del3PanuQIEJeBinZOA6uMZtgRWKD5+of4ZwrLLeTdTqXhM67ltxoX5YQPG3VkebXB
0hbQFbsSWC8CxSLpEWgZmsocIk/9cd9Yn0Mh+BnhH1Ji+GpEww2zpjBRc2L5dvrLkMsokLoBDpEN
qmeYQMbCe9ZNvjiBnlDS3hzY/XucsxLcb+zasTHdVxM4dxunkZF31U0JIpnadtGfMVQ6xIgt5iai
w2IRx+PKiTJF+tPCmhYI1sbke37sNVxyzMn5Fm/LiIKzrdYc2gq6jbGrcyUzMPFWii4ZEkdzzUpN
v0PUijVzG90Yap9CypuE5/uMsm9a7mt3f5sSZC8ivuHzQ0jFqRuEExyCt30SiQdqc3uia1+sziY2
cbT1OnwEJhDZTBuu/cVrskWiKX2OsvHcSxMM62Y1DYeasDHOx1EgEwk24x2LHFEi8+FosI72q+fg
gASlnB3g06dHL6Ry92WnSf7jsZWXgVYHN0yZH4WxHfb6Oro8QOo0rZVgzsXCL8drJma8xzwS46b9
ZXFqSOaGwbY5foAr4pcouKUf5hQ0fGTV2FBL0ToP4/9T5KqGdSpXA1CuX7rD1RL7tZBXt9kEOens
PizLph06hz5+K5R6lOaIZyZgg1rjqIcZrxbPHgxQzwAwV1ndV1v5pPpF3oQZEAxTOblB78SqB6qL
DZmUqCsvyeNLb2k8ym9zd0UKJ98kWRcLTqy38DEEnKYagW3/F+gkUT9eXTWWkW2ABH9K7rurOTuN
jxlv8riH7fofFTz9dq08yQDd4eGNRFWYPIVF4q3gkb/Sv8tnF2G9dj2ghvqzp8QGn+0TH1EPY96T
Zkenkro92ltncyM1kWpmxLWtrF2CLTPjO/yIIL+t+gEhoxCY29dp8kodf6wG7JGtn4RP8SCPZT/l
l2h7sTr1dk3evLnyp6w2ALRz5g4JdgNOTnh8wS7GsQ78RxdwmRKRM2vBliIVE/xGcYYDWvJlq7T6
sqN1hpRkC6WdYH3+ekUycn8AwuocdDZAJLbb/RS6NiatHUXzy0v/3sPNnRNJDU6OWJDdkOXW2PJi
YAmnbGRUHOhsWrlnfM7bXgWcZYQsXwSN/Gj4XDmh0c+Xy33SK595j4ktYemPUz/8lgRvL0vi4NB4
fHlIANJWJ6oNsHx+iXyoOX4oGFsypaUeC5fHZ7DRxxS9YC5gAjYQbf5Bs0tC4FXIU9L1hKpYN5em
1s/cXOA1SBtoj2xlHo+VBP6LXb0RGl0kBz63cOsfKe6Xd1Mgk75Dw0GGA6KHIX1c8oKaWNYvcSgQ
+tgIPO3NQx+lA0OxVnBKJUbzrSUH/UDUGo78O8XHRpEYn7ZuyY7cOGJQ9+FABp5Zie2LU++hMLKx
v0rNuIZHQIoUPb+vp+LzfZbD4QSbsijHdra2TDT0/WSd52W48Hs5Yysd8LxiJtQTp8/QfnBYilkq
c2wkW5nbI864sPQM1PZZn0ba4FFzpdt4cgR5jcweY/rNzI8kamGsViZazuTsYNFoq3RjseE9bAeU
fTbnMo88bWsSSP/1FWsS5aAc//caW8hvghq/V+9ARNodcqi/hd781C7mT04CvwkdnBLbCGWhBLSj
tYXc/j+yvmrCWgI1yadZsBO1xTLo5ZT7Et+rUA2cw5G5jzRUtcxeDGTlgqRfcZQ0SJ18k5m2LpoH
hIcW+3zQBYT1sio80h6+YA/8Z6kt2gNyp1otFMiRR9wGJ4FjLtdlAJAQ6UX2C7R7pltIKLNFJ0nO
dJdUbNjKt6AndcBeDNqFLgfRHsAGmdWOXosakSkNPFpuW3cshuTfWLISxSXhYYYxi4HrUk+l68SZ
uBgGrxkC9ceqBekuTX2SxOdQM9ffe94z1+nJBSFzPxZnzn+DUMAA2K3kCTeicARk9y92nFu8K7sO
BQBtbhtqBbHgwcVNiGiRkz62vD7hsmVmbXH2tcyp2V9P7SzMUf8b4t7NGEwreLuljRRcZWhcN94I
Z0x+RJ+b5weVRicWFsKqw2tvbUp3v1MMF6XgOMjizIGXlsVegwkMMetK7zfQ9KjE9bSl63Wo/Ew3
bBs9FMe4UeYbWf7hKBPIN3pnOaZ5iRckLE0w1EAuG+seunRxbkyF7d5stpf7J8q7pt5rvSJuBL4a
t1xsYDid5zRms62NYV3cUr2u5qnloSf49SuUrCFfd03cHzS+D0Cq2SQepPgdPChlFB/JSq0kbs4C
sVfx2HRrxuWrOX7JWM+/d/LEwKuIE0nwIn5lqS9QeO9TOL97qcWW99UMdrnTuiLN/idx/khi98TA
sieG9cJdTXZo0DTm5rt1ihLl61dmkpv3TnlXbcFRA8ID350JkwUdGBxeiFxzBSMI5ZLMjTUdFK9y
LhNIGoyP+4topSZqjbzIi+I56n+A/yk7MrMp6BsVQX9i0cfD841l8cfEWEmsGrqjWzcfuWEQDKZ5
lyhgQ3fi8yrLt9XsoKwOLMb0MzI9ZolsdIrhTkNDFRdG5My7ooMBLpduK8wb/cM3J4pNt/GYi6nN
Ze+KThBTiryFZ0Nb7UFbGcmYkUuukMvSxOX+QKmAoE8AuxeWYpviL2QvaT65Beg/5F8oYHptG6as
IXXiuSwpLUY8pYOtjh7MwpqnX5XApLELA2YsDn1+ZsyeUZ+Ox8akguQvTRLvzWVL1+2/fP1A0Xi2
Tz0fS+whF6GMpz/XOgv3gLD9t/grFuf9Kp/ym1mkLxGbZGNWxEslG1V1L5kKD3RztJodr2eNFKEF
3H7sU3c31UjemTyt4lZ9+i0HfWXNCyt/EH4zILHGzOa7xaynzGgtMDKvL7s/oqzt5qX35qP2GteG
hBZ3njFLSDO+GL2mTntbI4S8YZ5cx/UeAZySwbJkW9hBRO9tTm2ECohJ7GZ8KBnpG1wn+qJsunIX
nQMZuBnCTuX/jCsW17+lpQ4nXcuKhfy39YdxUQa2oKv51lajlD3B8Tz4+e9nMXGJDj9n20yMwpVe
nOfbhaIPpfdjuSung5wgbfJNWUqXB0fUDavkxMR2aE7sKWnQgdyxfFUmzfDH+OlmYMyMqEGaponS
ZvW2cuOqxNOQ4U0rQaXezJK7irvoRBzSHP9dr4oo6YyjTzNnLxYllDvEKYbMAWNfDfg6p+K7E5+K
RdASGBb5ganvpe/3pVEyc5ijRY/0HSSKIuKvp6zFbYQvWAjCRHupIgL6If/tDCeyAB9xcj/rjG25
5Q0llhGlLz5FIY3O5YeJ+YJwjiJmpr1p/xRNj04CU2CvwUo7i86KM06wU59jfEM1EzBDiyjATSCK
mMWSM1rpDNaodgNzniwdp7IiZk6B73OMFcjRiRuD0UwBhlHpNOnwpoTzJ1EHm4e0rXi+nDUTxuZe
z2TaANxjqCc0dvfBSxInxUHjrqHsXAeZTj43+xI0B2ngydWx18BlF3893OUfrYfc9cbjU0GA+f2J
Y37RzUbv4XXT728SdhAKgV6WL8mHdOaCNDv0bdzZIWtgvdIw0w+WBdBi/qkxp6FTUK1r3ac/YLdQ
OIhrtf4FN6eCmgd9MfDCHiejr5JhPt1Cp/kI0HBCBi5PgQZfUmM8JkZvOiF3k6CRS/3XFVfR/tuh
GUqSREGhHXTrUsimDs0GJGtBltfD8qzw1X7JmoLvgU3OsoQbA55XaHuO1wGLwVH3btpo3bSB8BH3
uP5sUCx+qFKv2bEvMIoV/73DUZsDM7/JOyPlDGCdu9TbGwUUOdhRe+HyP38J6GlIjxLfHzyqkfA+
LsC3bUwVEUNe/fROuYLpfzl+gGAqpXhGGLghhfvjs8x8YMBmtelztwt35CvZzD5hM5GnicXvBQkO
aACdpAhWuak1OpeP0WqC82R85Ms2d6c2XjBd74l6ktg50JkYe+2tifnO6HbWweE1ZZb0TM//lEmx
IqtfAtJUA/BPF1dw7FwiWPhAP3ZZswI89jmsqyGusQy5/3ARM3zm2ICeNHLlXa/kVhbmSxagzLMh
XGnsQM7IWXLTxf2QYIKkwSD/BBhEQiSVyb1T6Q2zMt6sDSpdN6Ju9nd8ItxiorOv54RVonQcror5
unSHP8T6xAVjvAGqvexKtUFahpuj0UWPbmuo1LBDRWEzsla/nSHdJhMxeDgT+8C7ojPTYsi46tF6
d+sx/LpDNm/XWJb7htfRtE3rBnn/WCs2ewbS+vME0MsTeGcoZug+zE8GESgexICtWH0JPVldIv3b
ng7al8ujxy9Qoc9BTtXBeziFma3hXlRmRhr7SN0KBMyonumT6aBIExDr9CBkoQoUvRE8+O2x/FFW
zPpfSb6ZOo2VpI3kIFE4iKhGqkNZiLRkjW28/m/CRk348zMWtHFQmjH1Z9uyzkxw5iEoQl+QTisP
wDKHGaJXV3jlF+MZS06x8R4shEmnejvsrlv6OCMpzXqa/lAyq4WvvSu6wNk35sgyj7RLsMac9sUr
hO4iHKfUxmycY3gJN7KrtvGeE8BTq5fPTthVzV1mYTgMLciWgRsuwm5UxpjAuZcg4nLtvTSSyvcd
wfrpnwRcWbLY127DhnbiEW9+ep9Ez1pwHSgqMwTLIOKlXQ0NYRzkz6rX5Njw+w0xh5RnSiyO74Mi
HX3NCCL8iF9LJI/ZrDBlyaVCv3xW7AAYsej0fMbpWG96C7lYNDGgr2aHvzhhBGC3ov8xC9Gizcah
I0hweQlUmQtJZJMKBuntB4d2A6gLCFLCDQtk+PdNTqCTs03SjHtGxCpHhCgeF7Cnm6PlbIf5E5X+
zV+Npb2RuC8SdorAWCSAw1oY1FyUwBrIUUsQ/r7WNuHQX1tTawrZXGMrJaT1ALEMOf0CF18k8ehl
YBb6Y69Gz5SBEeM5dNRtwnFay+Mte1/KoNe+VRe9x3dXV8EDAmGNiApb9rGddkz8iKH5IjR8ehv5
DkrF74n5hTFEYiFq0tw32tLueUn1T7qQRiyINxVKAT57ONKhzYO4V1NaaGnhFwaPQpS6ap9Fx3Yv
hca/lQ0t5r9xsOP1BCJJGnGHwAIuV4Dweos+NyVNvNJ6Z4mAovFbiICiODV7Le7Ks/JEHtGPJpaq
yCfPxt+XeD4T9J5vTPfVYyELG2b9UBzTQwwkyCt/l1zUa3jlH+lGuplv0X5ElI0I1HsU3MP69mll
J6t6YmWEDe8JHLo08W/mvC9leLe3fXILqh1z+1eBiaF5eSARdtf6p6eyDE8QhED01FonULBlhLaN
U+/zEoBTHy8yR7OneeUqrN6t2oyMGiLl3ePC51ejaq/TTFqJc2lHbA+gqnrFL6uMhxfXY6fHZ9XF
4So9k+kFSmwyyn97RxnagGV+3L75zijEFUEI0Ojafx3HEZ03QHgx5IfbAxZFDYAu1+WKEkoOuOUl
2oRgSgVRnozWVestN9hknBBfqxD6w3nIcqgGacbkIbWzInfl0655rv3vAugkq6MK8b19vWO7lTzP
Rz5z/iIqoW8+yzyMZPYLQmTo1n2UfASiqq+w6RqTeumVVsYfog4XSUsI6UXuzKb8VwBGVzE5iaDh
veGUU1vHQRxUr+2eyNW1J4Y0I9BOM3VXLVVGPw5QBHV3itJCB0iEhvbbj9kMIwcc7rXR5DbetVp1
qBqrZadAcajo5H6UBerRBX1jOCa93IfrW8coQXvtcNlpY4iS5MIwxoWxpZNoAQ3t/R41SKCg40pz
qVlp2j2xiq7YOt5NTEJqlA85F4Acvub+YZTV+cuY0rCuhKcTUpQ+kLbuVagVKQWgjqDPtyBYJWDU
mcYrGa6R1vMXLpCwsVMe68wZVTC+XrWlWiKY33zalUMLB2fUCb94RfWcXaOt8ldT7oz1rVePZMWh
zINK6UpXugnSLmvtX7lin+mJoma21OiLGm8fNDf93l4GMk915joC+J8t7C9EqtBiGQLEA2GgXSjB
8jAcwyubJCHNo1cy3kK8v3Qzhoh2Jtz4QyylBprqA04y84EFBwewyMzONjtOXpv1OV9KCoV1p4Kz
wMsI38HSA9+C3IhDOQBo1t/RD0LBy/QmysWrv2l6tjE2s9sbVAmwTum64DLj0++RZD1MsU0PEu7V
wCRYfV9/h/uUdNNdk2I9DOPPtdgcZ3Dwi3qYBfFBQC+MyrdQBWnKZgUNNwgda1NReTLa9yEbn5Zi
hdahkz8rDGb1hct7TqnKYAKF9IN+YTmFRUm+veUQjAuz45NqPeBjFxo/YRVfbCgmaDtWD0SX+Rqa
O/ESQZSJH8v3IGXmslqpbeX2VJfnDURdzv3qiLNFfbnedOjqLQ5LQm4fGppUl7QYePF4n36j2a46
1yS/OTXqUjyk2eMVGBfla/sbjv/Lx2ywb/P2WMBYCI7Cn3qsWZsry4aqSmeAlRrcBYkAmz1Gem46
XyZaQuPMtotn+7IAKZF2cdv8ppGkuWpWq7pDYowo5lYA76euqs0UTzmfBb95GNRjStQvgiU90lnS
SCSOW2w9j+RoAZxbr2MfQEi9D5qlHrZEA2XoGSrhl2PvulURLQcCaNRcPaQ3msJNOHM0lW8zOUFA
nofeQ538t5z70EUo6+In+5Re7kG3SFzx4JRfDFBAbh09lqNVWxGceW61z4wq0be2hV6aOgxHoVBd
V+zthINOheV66PqGcYXG2tVjwglBsfzLhHMuxXPlXZf6ajnOKt3d9OK85H/f0d8+JE259AB4NMYY
Wumc8t+fZU4mNOFNM0gMvsYK3wmAM+WTx20Z/0CtGx+8mGeA7hx8I5wqCeDELGaN80y4W67KvGy+
7oNPgc8BtGxIlYiV2WWwk6TT9r6f5CMMPvEvRYmqkm2pNlZU1VXO0yHcmphYfuXj3rRGtR+pWcM2
Ld0tW8q/I9GFafU3RKF+Py/o8v+eUTEEIRndRHgkkhsflOibQSEV0x6hILPsSS7KoWyHI9jTe2Lf
AmOimCY+jpzwoFK6JZs/glY60uWko05rVZG+eshjhYMJDGL8bYZOP7NBOH6zdnxwx8NCSjK8ILxP
W7Xa7NM7+cBN2e8NnUXlIZq/6cXgJA7d6CmVDeZbdU2J5GzrdMfyAu1QkfsylRM9ECZyfoqDXvvD
k0Yn4n8Cu4P6UDh6K7FcwFFfJG27/mKihCqiz6ouf280sOn3cIn4BQTMqy9uMNz1+tlMySEoJGHD
LzWNVNimwnKxl7OVhwdM0PrwLiVbLAlhrMSf5i1VRnr6UhxYyNR7om0lMxRxMBZkT5Jr+ayg21Kj
obCJe/RYKG6F9qWFNBpH9drgFOfm0Luc3N/Hb9ERGUdAg9YUHXMSMfQevxKnTQb7J42KiT/jCMea
qlZtPuD7XIMHhlanLxFL1PAvhlMTrmPOom+WpS1UFbK/a0I5fHkwlMaUslI3Y+m7rb4sSBmA94UA
36XkSdYvCsGz9INZ1owzBF6izXxsF8X6xrnoAFNGB/lCTA14ZfJ6iD6SD8/bWFAMd2n3KVUwy0s7
PGC/PYmKtnuT+K1wWzLmt2VL7mpNiJChhCft3SD73qsF91cbwBGBCuduUuVP0NrXerA3Dmt1JzW5
U9FrCqyYNZXj6PoA6D62Xof34zjv54NGXJ6929tW4skndZBy3Rop65fyXUusVNZoDvxB92K/cbkO
mMwUKTazLyPJAkt25to0leP/5rb8q9cD+Sm4VZoHzntruHUAorURMlfFGJ8kh+PCDOZALV8ZiP+Z
OOsZ8tkyYT+CDdrbMwcqWq8LjLc7H/PRVY887eySSuFZkwoCHLyci2GqHtq91ysAnQPWQpcI3o3T
R2gQwJu4yy+otz3fe/xGdne6jJJ9znK8s0YlZIMjcfT7U8EhM0VTZ99y5ovDv70L/pzCvUOpUdHy
wJXqUR8zZ00NkPtPGKhkyUXND7EHinSg0LsaJfLIRSj5Ip2j5MgNy2ifgTmp7Lo44PYEolTR/pnr
UsfJrwVmm0ENlTI1hkCM7gy5uhhro8TdUb1IOmqTCQblLTsOjsuRqgvZ4yseIZXZSQa+cT2WvhRA
u5qsKrc/3pkTfyT73HK8UBstPikCQfX3R9wd1HigBDII/BmqFkeiuNlCaAbDapi7Q6A1oV0CD3BF
lcZdY5cFLOQ9b5JaF78NtzHvy3wP3XarybxnBWIwigYldusKr3TR5KYvj1EmglSuXytnSoKwc+c6
EvfKmgqNgoMzw5i041F8j6n9KqfVOH3XBHfrORW6AqyavTKXBg8qAD8zlA8H+fohjgV1dKDwIHye
RXKo2gIc9vtywrsl60agz5XLYPr7JTIMwZxpTdk35vWOJpGBDr71cS94ltGk6SMmwx7LPPdIhdx5
TcizZP6vqqnvZwGwnj8sjJ7RDn3lVFoOfR+tirmo6+MX/ApnXxiPksG0YbQMJvlNF/ZJzc+gnmaS
oE4wHmTooC5fxT/hpfjd1Cl0Id+9oVQIic5XFednBL/flLX8mgU4PpfzmJ5/2dNyWkVPtcVtB0jL
BpqFZWQWFnHeCivUhKaTvnCZ+8qqV+pw5FVj09PUBQczfjVdTZe11biHYkprOqC8PU1P1EcFe0ef
KI88NllA/d/t26Fei6vrLIU4mUQRHIaK9rZvXQnv+rvHbnJ9VdXk4k9suRkPZ+DUrossGl22dFR1
m5EgZL2ZJFFGUHWQNku4f9XjlHhBoAB1QZpAjuRNuSf4nDCRDs2tboVsrU8eaaK9k4zGcHfES6cA
reIwHMyW59NDDBiB0cOlO7C/izSp3FaRIG4kQxnhxeJcvS2RLBQH7VAkdf0t0SbktlQiWvHMWuRd
U5nwvnaQzgguXFhS2wvm2MtKR7hWf5HUb4nzMcz7+4qHSOR2RszSkrlnbQoI5CJ3UJ26SM6F1Nrs
yIzERVtUlw0I7HflO8EBeGnucyFXP9g4akizLht718azuu++v3Pcu3hpjnRbnLqUbZNR89987ygW
IdHfq42XQfUuTMP/dJV9p/0qq0upcYMW7MkVOQ0u0GsHvwgaPHvUlbmHBHfkpjpbucVR9b7YK54n
bqpXv0uL40mVytBKRTD8TOo7vbFXfbzXDmZIqyBHKqAxiCGgj+kbx9uEws4NZWD7+wAKvdSG5GNa
oP1xBzf834m26+tmYvZkmrzmHsp3qs1nc7UgzhK8P30cng7T6K4bpDYVmFyp+9ok81m0hJlh07Ps
LMm0fHhAjxvlwazZmztFbLAbK/1AJfRgSplMXSYPBRLuJxw/5falwsjNkgx6hYKPzbGvW089w+I0
b0JBNZDzfTRGJaQ5KEar/Vy01Nvd36dQvnfMzHZBK1B1+67EnXIPGGjYYnL3px9hiyHp3Ocg4cAB
wSJIbO3oR7iKGBkOv5I6thliV6xw5JnDsvSP+GlV5IETfXuOhnpo6pNUA43yy+sRZLL/M22oOSZp
zhBWpgXVyZ4Bf5b/XTDfEQh/rYyHbnBUwvc9ByXYN/OgWOx8dWTqu8cwsVuXhbh5oqo/5Qer+1bl
Lf03MxgAFpOZcLxU1vfJYU69TOG6phTASj8xQevJzsrnvSS+zmKpnEZnYFGzajdxFGrz9fwLyqhW
jKdA2cROSiOFcdhgsbpw2XHAi3pg4RXIMg9ab/XnoCbW87ztJO8YC8NcycoSfdkYFzEy5bznMfFJ
mvq3+OioDQqTx1Xp3avY1Arw8Axg4XlC1/8jVkxn5zj994NxpCyNVo4tlR2Epl4e5sSEYvyMlz2g
lvT156QUKqTosg8sJwYO9dr4kaEA2oaYB5JRAM6YyAZ4rojVZef4+ybi2Wja5sUZd84dlOeXkLRH
5619xnCRw56oEs1fSCEyarDq5XgPu8b0RN4GLNW0lxxKeoBJWVnGleOK3CgyeTTRWUO94htnxTZE
DK7U9bEtjgZ38GBi594UQA49J3rEXdwxteVNZLgaf/I0Z+jWg6ry8lRfuRmnHlN65Eg7KV+2NnGs
eiNpJUz+Fk90kCD2MKKyGNcX9hZSm2PC4zdIcDjGlqlJum5lnNG+C634Ku2HPuEnP8JajIDZ5Tdv
a7mJQfOY34derXZ2XvePwmZNqdqUMy23KrfJyueJs76iExJx6PGUQirPwVPzdQAL9u55UqkUiZLN
E+4LkGGaRuP6jw5yHyp09u5xGJ3SEXLg4pqvGVO0o+lzLiwSZ2tbsyE3/5ntwV34w5BxWkXkTGLK
4tNK/jpaLeRL4dN/YGg5hgCciyyRapij+A87i9ZvKv7w7Om2Zxhn5DMNLFcjD92/KQCKRViv4dl3
GOpYz2no1DopDOD+XRaMpePdJSqTx02xLavrm15DaT5q/I0paJIY5QjNcHJxdNEuj+tuxt6/Dqjo
1iqhhS4gsinGomUwNzO+HBe+WcbkPlqHgzh8dPl17lWC/2jba9a8EasEFBFTNh0ad4y/RbUp2k00
usBCEd8bEkLq1bruqanpe/wZ7+IAaIEqziosCeyzy/i3g7SsnRj+srhrB9eKc72lk0RoNoUNGzdw
WCmStIBwwCDkU5YnTnP1xNdnlCNvpp45WdWq8JXyeY2KraekeGoN68Lb8lGMl3fzarQGkRrcHW0d
dJfJ+yIkbkliLiufUXcFmZtyFthYnP2BTC/nJfSSw2ZcJlTO0R4JXHCwC2CtGSVf+iYWnwShGBlZ
Ga06y5A1c8mXrY+XR5h9Tyqw25F/keOi38hpSlY9dSOShEWLNSBdDrFrRPuRwoWV7o6O6DY8kgyV
xzYBdMlz9Qnp0aLos3i3/ETU+r7s2FT+lufx44nyKNjgGvuVrxW/WR3RA+upizq1Um7oj8Kpj5gv
cSrKvZ0z2oMgtoYa7ZgZxFY9zTV3RwgvPX311vKioL1I1jEgwmrARQU9tl46cDXTihrcdcK5wrrd
Gim0svclB8Jw9JrIj52XI9uUQOtbRSRsFL7dVROFLWpBX4x7gJPTaF40JrKWoVYPeaD6sLPOJ5y8
SE1Fn57p2pBx9eVvgv3EitGs0QTnPfaJURhpn2E/Vh+sIXorfmjimvDaP6+3OGpwM5gKkvg43K9P
nRQmWKsIL0hBnUOhF3WJbFCAaUDwxidj7n74G26JO0T1Y8Qw6s1wvs10hhR/LBRaIVmnoZ5Ae8DY
ZcjO0tL7urYxRtfovuUpxX1mKtufdayBzrhfoe9Haxuu925II9Cfz4SCrcE814t+tx6QIIRIpGWy
MzufNQLwAEXVKvJfFH8fho6oZfy6aTYG2WEAxmj8HnLGUVVKjWmzOaJ0nXqBvnSB6rMwTTWmWY5F
9Bloy2w5BPsvexI1BQFtIHNz32UIUYhJ7bK0fC7AKVfb5ighB1TKbjGRWuhjmqOL1wK+BuP1mDzG
anOYC6g/59M1TbSuUUXzXuFExMYwe6Mz5yoGXMJb2QbSQxc2ir7EO09c2baA/43YoVzkeGBZ9s4G
668e+h66Id0ISR6W6I+6grkL1imTYT/+qMNyXHp+Uzq3Oe81FnrD/Hna/AvVxXgSFsDkrt0TJ3qI
lxaxYvPnBOrBhXEWOBXG957/3OjpagRLNEMP6KiXbvhAz0A06UiNqpoVI2IKtsicvfatOoR92739
D9kS0LkTVPg8aar1BqvLf6bMrYRCiD46Ug3sha287GS/ay647yhOOcgIdTxFLeBmOIHziVTZCV0I
M5zojVE1jsDOvrSrIBnw9jyM98ufatVpSugXo350SEvP8lY3ZUAMtIeWWMSUM7ohqvW5XUaEfBXk
GunXbjkkHLX0nBWGvZbtzvoacBXTBnb5IX1YjSXUaER+daWFrmu/l/2TyWXZ1ED2NwQSzd0L+ibW
yc8PIb0uDiEFNWlEVtinAb2tP/3b2THjDHU2wJoFiBg5Zsban07vFw6yBavf+fumRKqSghUqLWV/
wU1VonfIA1ho7WlahEv+8loEPG8qbWucxmcRrBYI1FaZ6yiM/e22Cn4xWshzoAWJrX/rYaYd82TP
EPddQlD6eOJl9A2475ZX3Ya+YkNrOAtqYw2g/54oq7SW59/KFnbbNodtHiykQnQw35Jr5XCVpkbb
URKzlCV7FZ09Au/yVmrC2PpFSAAU5gaR9Ruvq/h+t183fC77mxO/HQT4H/8QHgUJDIAiTKf21QvB
uKOT7leCjzEGW/V43VLgGhbGQiXrT2snc/cGgbkoXrmzyg/bBDMX3vAHNDf3jC9elydrfB5d+ti6
LMgMmu8Oz0R5ojs4uIhq1nAXSjiwrZCWFEGW6KsFPb8WPyAbXlP5JYF4jg8LgrExAJBqT8p2sjtG
DnOsCfEQldpY6ATqPwR6xg58AC4bsENHCDrH2O75SlhmAZaUyKNA3biFdnnobfzTl12W+/q183/h
K6+SOeTd6d9Mio0V3w9rPUCeX2TNTRAMmcf2kDBSlCdrz+Oe6PGxhxfT0JcilYBvnpjAffEXfNXC
8rT9ZJLX1FbfBEtS2m2+nWxZV60W/XhcaInr06bYfeWd4tFZRXI+HPb8oWn2ixuUCt2Z66PDlCXI
L8v7V7zxYULoWEY5eIF7JG/6sV/bh4hdDL5UWHXn0IjPUI/hylW2FNQExPDXYhbdXdJPP0h09XmS
KT7fg2QsjeWxSUEdYMgiO7TM4VyzGtGSF0glo+i76lK1OvCrkC1SySuw8A+fOE1hEWlRBIg1dujE
TzbsFVFwXcZt/KsDSH1NbLcID+AcR/QEydLBSHMUj55WqBNKpOQwH7CZy4Wf64bslTcFEyFnTJUH
BTU8iCei5wBun4tvqE9W7bIE7Ih7G+roO0F8zJF+AiXB3l76gIt5QCg1n49ht27HD9YVDAXX78Pj
HABD5J07ALujNPtdkAk5qVoo3fC3IgGo3bcxLCRrjjWW0a9D63VH8MwebhOelM/wJcz24Qau4VvU
H9ciPHpqhoTExevTM1CJ8FAfWmexYfoOoTmEarTDmzsv5iFXccUQb3myUcbT2+5GVw32X3QaZEfi
2ONQ3XYkR+2y84zWvCDSHbUh3vEiXxNQGFJx1lxs6gQSZzp3x2GiwCbVWd23NhDdqsyV/D7bvU56
+8wfnlkRzp0lkpRxq4lirex0Q2f0k0JvyQRW6STpoA4CYvp9BLdYf1/jRDBsuu6M3rlutbTu065L
qftxRwMtnAVaC4ImbufAhLNkGaThe92WFlK6DQ9CvVLbjlrhzr0aj8dnES/7WZg0Al/l2SazgWpx
k1NA2YxJVNrr0TmxkX80D78I/afhegfJ0mr2Plm7MMGZXwrvTHtVStup74FqXMPfbWaZA6R57sA8
0HWXETWRWZkFv3bAJPKDzBL/FonfdT3LXcKDdDuNLnEZwqAulVQmT2sS04omkVLmu96GYu8thivc
9Lkbgq5dYsjLt1j9p36kk0FZTAZrzchjT5b+YX3jRQ3S71k/WbiGBqtF1ZP1CuvDdOV85PKh7a1w
8iCimsuo+H5xy5AEtez6EY5cPGJJxzQuqu76ViwS2DA55YaZRTMbIRYBCuE53GDLyKwVK++f3P+6
M6js0VBFJXIOt/swYA4hLMA7rRi50luGz5yeZ7UqmdVx1C6uXCCBBsHDqsbceYMV2QJEW+kFzvpF
oDGzXpLeip0PqHp6st330jlEsaEBm5ilHBzzerJG55DUzao1UdTl5zjvQeBECOOWUF73fPgPWm5B
3IVm7xhJNjv0sINre7yYsCB7Xcsj969HajTbIW4nz/lq5FjaQOBFY7+RN8dktia5oEqJKLkTBZGK
AIgzF0zzxMVz3ToRNQYGQ+hAU5CmadtrBOtwNGMbzJlTsP2wsVotDOEaGSD6k04TZHHzYjUkewKg
7U8F1FoSIIdGR1wVJHelcYDRoG3ACb+F+svkM0eMGGf923QDzpEraDaWUKlVD1t9nYDppa+mOUBt
t+sUTTuzzViOL9wwQSBkKgHXJ8o6Q/R6UFJMEm3qWwBw0JCne0k07BdJqklKMuAHCl+M+JZdnE0k
ic5kgYYEnB24YcG1NvLf1rmhYLUTTgcOY4wvhEdYj8JMb91bGsM9tgCsDVPNVf5JfkAsB5uu3fkP
EHCmRKKTri9wc4otyp+7QvBU7W3V202JVeljtYP67B8aQPBOBMXEhCAgaRSYrh3y8seQ6O0Kt592
d3bdeQT2JPYVO2noAqID0guux46IGwZPAUqA2/29O46bIV9FMBYCzBbUvvFuIfdWeGB4EZnhgsGu
iJU+6Zv/qfhR5taD2URUknYui1BCFqGoHASA7ICGw4rt8gwHeqKDKRk0c1Xg6fdDAPy+F8/VvuHx
fp+8PFXRkXMG3E4fDLBOWuWrejPTu33HnbfZ2Jp+NLgLIrNdBdZUxsMTWJa/Uv6muMuGMK+QAK7j
/aOrLrVfNPiewwPqnmicOsTkDAjsDELGpXXcuLq5Yoypl9/sIB4qrZM7RrZhxbCmgldx7Y14Ga4J
SkcntBwS5W2h84hUwDPTJRr6of4jXXtvw07tnZ4EMmircLLlYAjdk0XYwVg7jCRBs+nEvBe0v/7E
DPXocgisBpfpHkksz0k7cQuWGw2/7lPc2qGtJsnqNhafMH0EPrbX2tJbLtmK8r7usIsK0wRzuYmR
VSRudXBWfGFdqZscw4nUE2jqtED9fEOlEAUn59+X2nf5V1gAOEOgahUOMCWeBXmpms2VPnkHnXIM
Zba7X15dAq/fnJOazkwl8f4hPAc5S4wDZmtehPJ5S5NHR//ruaU+Y5qwpW1whsIGcPm1H48/nZ8e
dIDi/MuTf8KbsmXpMey0+y37nBWL73zTVx5FM7Lk1QBohdSqicf979MZYMoYcmkJzmtXCaLqB0Oi
lD3IDROHDIf3N8Hsrc+YwIAmZF9jGSxi0aULEo1O0ljEfOiN+TyaSkVgjJ98m+EHDTOtD2QnTX8Q
GMOafWTl66fNsSKQ0gIpOrBivpmrTTt60Yf1natYd4X93qUU2UB0999st6qeMsu4Jl1o7MmOL7bz
RI6th2uES7qhC6ZmKvYFTbp0f1l3YmiKyJz9RN8sY7sv9lqUruQlAkjUtCFyTVmiGQh3xbty0y+w
WNiVHbXWhXYryxSZw8xpWC/iCQL9QyrpR8RgEqSOoKylUMNWEGnDgPXJ/PXyqF4+u5iQcYaunM+4
WEs3JTjvi/wsdJtF5lc5BvL9R9GLSHsayOn5tii3xk3a7TUwTx1moGFqxu/tA4mmK3FKU4G9L+ok
tJ8Sx0DfWKSNYiY4b1+2Yjy6pHUM+7V4xwidvrz0WQOqGimOfd3NB5nk2rvF4p7ej/g9nl2YgO5k
m2X/wDLuEs3CJ2F9iOoIwGT3IHOQtdFI/KnrE87o7WL3lqFNrTU2IX1NzfwrJ93fX4Bc9kdwtdSO
0xtPRIPV8GhFZI/8iXykf/3vpGGlEysKT68B+JCP1CBXOqrNX7aP0RXcbS0dvMCX2J7LKajfsDTt
RirfcAy9IHwiCfu5nqWCYSJle2FHzJ646DNDFbbesuOTfH8+6Xs8TEQZNXxI7/ch4ySsqUanLh4v
s2ppnHOAQOAMyERObZf8Le5oVBYohwiwaPSnAAyxNr1ujr99vhgdbWNA0LgYEhpJJzzX3pfeFffZ
ixpWGlHtbh1wJQRc+dlxKVyR2XqOG1/qMZJJBXiP2dIkftv92q7tHwzANKywrL2o9T/SUnDoX4jW
wSYQ49DMXcGpxqer5ZJXTwkwL0Fom+NrAjRgbWPddqp5yRJbWqxAK+s3weWTs80CyH4ijDZ9K6uY
VhZ2baqbbFuC+W86CVHbREH6KIoQu0rl0lbQDeE3hblHCgAvwdgLgqxQAegGWR/9e1WknVAeQzQ6
xhrML6xNBXA+V8yRRxsELCiOi5EYiEQB3vuXbEv0Jl4ABMgkNJcD8nzL5c0+astAJJLAsncs6naw
tlbd7mO72Y5cpxcMrXh6FSh3NZEdmlNnvjSByb9YqtM/YYm027cwBBjBE9u5/je2ecAtbDKvkdF0
m5csF5D1gRUYnzX/+HXc/vcwkBhgr0VAA9RBeuGbfIGpuA+odbyAKSa9LL0Aw7LsN2utTb3la0ey
qqnrupp+vXo+a9xQRpdkooaMDrpsmY0FO0kRzUug8JRyHPVPKOsmWQs1LXsyKIw+uu9BRfzXXG9t
WpU1Slsq1IkBO3pS/8YcwbjnEaqBhDQmUnPSfGQslAbpZ26XB39ZuRsGn7MdD4Q+YlCwo2HmRZ3I
xxnwOEg2FFYoUoYxvmBLbeYmQ4fXMKiD2ECQLilyjoIdjkWDhB4K+ofqkAhcNqXvVSWdeiHKecDP
ALgEQoU7stQU2ebvC3l7Vk1Va57y0GdFeuMJRiqBFBpf6OBP33q9+8ChUXNwkWegxILAV8meCwgP
RpxDHc0dAOMEZuUK6aFLYtoTE6Kyux0ME49Vu249TUntKyogXgSfDcq43XeyYclSAVUj1URUE41X
kXcDtt3cq7cyOkB6IYO66j3oAVF4wc4kPfhoXnF6ug8ncy+V0GMDx9BwCw19wAReSkM4kDmOLS3/
Y68Kw5q5Chx9c+lGkCxuVmdivQt+GWpYDNLjcUCkwgSrh7CU2X9h+y/w0ItzXif3WVgzd8a7cLKy
/ioO0Sbh4YbQdnV4YRTDL9TPzrrj8I1jsWl45kW+UZ3TPU2Hx8aPAPmWCzTF6Ln4J/F5WLJzJBOT
9XOsW7IG7lH6ZVO2lr/TlhaGIR4kY38uZAcq76X3ed4xSzkF09jXXppmZ7CMiryUjnfwI3z/DGbl
OheEj52lSfEY5k7OWPF22IRyuQ+P7Ctfk27l3ZGomml6UbEQSEMOyn+UpnfWrjy/1i/Y443LNsjp
Trd/MOGXYic6O9KsgeGJhBW9bjBgZyPacbBZ+yeMJzVPImSv5ifVYXCMOfZhdLAGILsBs5wRXvsu
E8EmUwl0IAG/qTKWghr2YdytdwEbLZHhkDBlSCzOdq6UR9jtR9/i8dTT0bP5Mxotos1kiWvSlSFb
jcZjSGiJXPNcxdP81Ru7aiayPmaq24O+g5a289irRvM0jJS1+zXH0wC1fZqCmwpGTxJYK7OnplrB
FuY8nzgqATMRmF0JBz/X/C/OAMCt2CNTgyif93S7CN9lWD2hU4BGpJnV4WKaw9edELqkogzEfCeH
++Luguz4Lof712TJPOhDHq/ukWc6g7C6+MRP6LScu8jSoPT7jTyGjQmE4A9iZoFCWMRtmChQVpNR
C/vaxzEBsikT0grsQ6RjVrdweRCrJbfzxswTNzBMQJ5HISlXKQm7IwmxKCvhELJVdGRHJJErp3O9
AtfPzZ2Irfa51AyntSdoQ7tO//45Th2gD+ttP6VrzRb6TRKCLU6G+KtVLvpSu3Tuyk1DUMdlTpFg
BL0spFikF4ocWwo8stsbVAsgCrdxaA3ODmM8+wN4leFn9BqYdxJvJqz03NvxsrduCdBTz+JqjKNE
3svT6WheUhccX9WM701WaInMOpG/3KnP0CR/BnKP9LHBXZc/ag3hn9mMJTt5ck1S4R+a1fdqa+FY
Ekiuf/c5HgWH46ONEVId3TDmbHhLnTKTRlj49z4ZveKFt50+s2wWndG7w5yfbiJmaMoi27sjK8xP
wWposAEMG3A0uBGXLtCYcPt9VawgxmBzaDBIyv/Cm2CxZyA6QbTsZkT5AjYKL7KCEfJD7LaQNVRg
Bf1Jcc8cR0RFf7kXEIEPQghzrgbmIC+u+8CFEmqAyY90s3grA7yGEBiwYZTmA/sbU7eIb3I9A29X
dLdecCHFJfwygZkZn03Xc/ZsKWdKAkQR3jBGubmzH1L56Ry4xHNZrGfYZ3Y9pUqb4dZrkLDC7ML1
JSy42aZ84ToHKBm+SPoKK9n4jiOqow4TwosKTirh2QniWQL2Suvd1uYDkyKgNUrkorXFnpz7T/uI
/BySQuq9y+DsFdob2C8NZJRhLpiOj/Z9+TtHb4gaMhZAbdA57lXHEACIIuIy54VF6H5N0DQEmsW8
XrPJRT9DZ+eDGEOI0RG7Khm2qt+UqEHfaJx1cZMFIIDJws16SBbbRm5f8hcFKlwrvOH/aebacr2Y
ed4nxfrwLDBqj+4wUDwJFw+yl7xreCcFjCBguBuVHKpaW1quXL+ToJHYBRBaCpu/ayBb9Ugz6DKM
Ot67kXyuf68kequlOp/CVF5mxx/gXN5I3aVpVsyI6+IbNu9gJKpXsfdVuuz1Rnibqkd1VRXNcTRb
VYGTqPRAzBnH14kAJ3oVc4+8R+GyNHtLdN441oPBQjRzT4i7VDaA9cY07awhWatPXBMk0pZezKVL
DvyeEnRr10OUP0FaC15nHrGqHnVUvPeOmAJt2k7e042TiyZPNfm43wAI5FIY8u5UgvwRAL80wJat
y53KZbGk/a0UWVKzhe4/iEz7XTbWZw/jG/xSYb1RN2bpmaW/BO1+ss6y+KZFyMTBS+jq+4RGZXDI
eqRNYi/7KLWMKKTCOSwbnLrDe7yzWCmyorpjdvlezEh02PdzDuEby1aNu0yUgJ3sgVzITRgNUmve
DBRfdAQQil7JorWW503txvcyJ/ACs6CTW3BCbPJ8X96IW+l5ZHuu6WxWp/Y0vlnutqWwwGmgYSfc
ohdeXnqLS/U4g27t8di//ngOtdE24L8DXuhoCX7y7K9HvTOgYzZmVTgWjK2fCQDJ0xkfuqAr0by4
OHxqAZOTvDafHyUzNgJO2OwoyqlwxZLY/3GrAPLGsZo2EQ1fqd17Co3qVtkvlMjW1ymVc9xWODN1
6jFQScEOwBwGneplw3xykIxg1JCOLGc+DNr1rf3p2tbskccKh+6XQWFYZ9ewzymiiTdboDFXwAZL
3Z9qZB5Of0o/BDZpjj4deBM83YQEAWaEeB01Mczp4b5dfvPZ8fUh8w6Ad3sGAa5/8yTZR7wkRPkU
EuVhZE9iqUZ+SB+gG/cq7qc4FbDcq//Pbhf4OcjLos5w69qj/onJGX6Nc2opAEDA93/IHJ7sEz3e
pg6MFGz41AjH38lPJMKHXc++exGOvSjFZl0ORM42FlMQj8z9ghwg0vZPTby93E5Xh161Q7g6e/zM
lga8KVBdHEAxg05jf36m7LHNeMjPQlOcDZ/cN2d/OxcPARoTmK1WY84wk5AEIUFcUPggWYVI6zp9
+Wt+DxbfV2Blwolta1OBxlH5EngvoMVppro8d9DuENsDPwJuA1hc5NRsJKmdN563n+ir6E1gocGr
d//H572mg44UUp6HfpGqxMpc47mxe6eZcLhL4D28OGHah5l1/p13EkN3tChCW4NqOjqfBkuKi5PB
CESsE0nRvrIL8ATKmR4UIm96Fq1H0AMNRQicOsCVAgXHUjjc7T1eCtgUcFc2Qvim5u/OTMrICdOY
BNs9uLhKyzOVYp+Yx1oHljl3WjJSGuQI7947E90hr29xD34lj0pOxB5gOSFbHV4Lt3PU0mwzKpAX
mYnQ0E5RBx1FSQt+98q/XFx2FXxTcfeM1OMBJ5ofp+MzoF4mkC8QnZgV9R/mUzf9RArjlFQihhSo
PXREoocuCJpTgeUjR67uS/O6oiHsFZ+qcr2GFHM3yIMUVhuQdyddKhJ1P+MEZfFzLWNa8NZ4ysqj
fA7s+91+rPcXhjvGUYZFgsKmh94nus92N0ivJ3Py9tyt/hgRiBJHMPbG/HK8vi6j9is2toisUPgi
Q0I1CQswqYlCPq/2z7blv40EvcTNgNMV6S0BH1O8nAfX+fvqJ+mMzAHqjhU+C1hobFCd0Hd4KVFD
Fp33qupQnrNJvIYQ6FnZonIjQcXqKSzGUDpBh4va5UNRoAFYR3wfNSkmM9/sdIYPOekFD7R8sP0B
9PEZzpaoxDqlX/WmMOi3Ftw0yLIBXG+yELWofYD9g3dczpZ2qWm33awuji0VWilmLFym7obyzkmC
j0w1tNgagdQLbYqPLvQVBAPSxH1M1G9uXMc9s6YxJdcFEuqNaIitMw8k/P5yZe8wAfDpnXFydox0
g/k2aWsVD2z6vR43LorkDyJLjRlZ9oR0F4KLWmpdgFiDk1me89S+lethWqc+RWkk5SpF37oeJP6P
fDT3Yyhwd/4dQBhnK+Dgigrv2biU1V9fDRcGBCw5AgVf7+O92w6ctZyjX9LEj+f1Hwr6pCV2aDb8
/LFFa3KF5LKuWzJyr8IBMKzQEZdUdO0ELbX26C2nktu02TgQZFKxuA7gjNHS4KSsdLZu87sdyBnR
eSQ47736roqP6FPyklQNLPVXX5YLcbhM6xPo2SEw0Gu3uIk42aWBPtcrzMB0tm06cx3I8FD2dnaQ
Q6hZ43sZT5fdHH4A6DRxEOkDY/3p9IfSBaYCYdhcTZMCfhk4MTw5wa8RaV4/QiGIXH/rZsVU9HkB
VexqmSZ7Xxs0nmPLY4ctnKxAhmFcLmlAOJka4FWBkI0BzwoFkummbaoZM7PmnfhaQ+iY+yoJxxyn
w7SezZsRhm7tP6CDVqh94S24r6bhaApXU3jwOGIx3Fl4bF2DZ9W3j2dApOEL450WO948lJf/GI8c
KzwwLtcw8130cwG7S3jqivbN0CA++skxCvXKhpJzarkF1/xXQ5i+mMm1UJ4idF/XKYNcE0ixBfs+
7u1IQ5iiCrTVaxS3n2wHPqwtJS63WQh4uzDfsvUXU27PFeR8rm7LXI3cW6mCPmMlxs5VLs6iTk0q
fnw2D6va3mZf32Zj06RJaU99tgc8gfWfxR/ZuAf7lE1TQ0v5b+7lwxef8eDH3Agyu1UKNLTOvvFA
Ir+44mEF5teT6RvkJ/J2ZT247RIg803ci2Y4+DAkjQ9hknA+ljc+gVKgtNydDyoxlwyo2OQd6Sw7
RPkF/61oyJgZVoWMq7TvSHzS3un56oxVgOZ3rRtUAPn8Q5TQqLz5Amt8fvum4G03+vawgbCGE7Y9
VbY8KrYa3KwdqZp9KwmpHOu0+VWjGc0Ne+kCG40nrN8MVBzP/smd6sgNSktuHLIQcFDaPb/UCcXo
rkt/obQZA0UgzwRIudyDwkP4HRpKr8CkmDJpRujiP78hzEBkoOiehZvnqb7CgQow1a4Z25L1a3Em
1e65QSy1l6XCJtKJzlZ2jTi28u7nOit5jFIiSRYNXlhsB4nZELSIIzz0T/t06xVZDKhlTNv9fqoQ
LYN99BYUc4Seycewpl58g/PST34moZUy2XrioT2wbwDGjXqZsSPLXGpCdt1oXJEyg80eJMTWRUjR
7tBEW/6QUZq2OJMZaUjOzbLO0g3QRT6l1SPwcoBPALXeiztJn64bLzL2Tg8j+AyHhqe/RwJJvjFA
rvITE5EMGaN0NTfSgVYoJtntVsRaMr62Dir7u8jqoByLcs6lCp+bMzexKjDp5judqLg3+4qaxCMt
tjIYUvDNawcnnJ/rbikrwiod2EqhtHcmL5l/6+kcB2+tX1bogKE8xgalRBx1vC7aTY1AvzSnu9Ri
LFosYzU/PjPbfBWu9eqzbGA8vmbi8vKI5FQk8iNSIbux4puy9Afzb5Ny5B75A6HtWiZOrwAz7ugZ
WWxy1o0JKH3iNULIfi1BAYAiSF0qsuuCNxUzqED2vUsWcYIQIUOV+xC/ap9Rf+WOolizRIt4s9+q
NdVaRIo0AAfQ+ezQA8IqLN2LsTwyXkzgVPRRqNrWukgAoiUDbzHWfGgHLmBupjOszvLAT4liWIZM
O1qRhkmwNR/wQqaxLWhiX1JFOMWVgmJJS2NoWleld6AH519Pt2PUYL/VtC7MKVtG8o4Jv0C7wWnk
gyTNXX9vopsDnrhY2glfLRhEeit+Jl0oRY6HbBaIZmkNqlYBw17AoH0iGR6RxrCOS6tcxF2sI5t6
o0gD6hOT+V4Ytft0jYrDSviGOGYThm+e2nde26pcNeqatDC8yOLNKv+cCXsoomY+uKgCLV5A8JAK
M55xmJ7tz41ENtacSUUhXclh7i0eV5DHyEh04bDbwV3DoJ4P0qEid9zQ6dnVtsslHvU7/lFut8eh
xWZ1dElGmk76t/oA12E17MWLeSzoeYuvGL851NUs/G2JB9X6n5by63nn0W4NYnAekh52IDWw/Oms
5thymwSLr4NPhFbY5nuyrmjJiR3l39NtxR3nsUS3qA744WjX3l/NF5+VUXz0YvN7vOBTBxgDK1j8
sqbthkmSKL/csob8rDKc2HxIsY9z8WteEoR6pvSD+wWDGQ7T6oMfXV5Ch7JdW1z6yvClLc5dOhU/
O2r/IHgQc8XmKHqjVxtI4wnk0F3wgKV5r1lnjLP42my4BuccnUuazr8SM1O27ymO7n8OPs/+cnRM
vELiGqSH/gOtiSbcbFvaoxnL5BTp+j+WebVIUphEziJz/p3NVq2uw3IZS4N4is8MDv3e+isrcWLh
grMJga5T/TdauRzUhfhbQXXTbbWIh6p6V0vVHcsggK+a4diQ8f38G0FBncpHShsdRlmwkI+4iF6n
ChgUoXPgP1BZ9chhPsTDYabC6UX9jS46ukjeO1AlL4EWDb6iaZBFooR5ssQVmYbqVRhjzX3FY7+Z
4wA2T5HjDYu5BramDp29KZA77CUJxFc9jvFME3YyyZ/QKl/3ZrtX9tbKVjnwqy1BOx+Zz8+9JrLw
di4/ORE6e9JEhC3Vs9SluNihcw8RCHcDSUZMYjwHD4vmGilgucY4lhHAPLRxk0EH0ZrqZaXKdGe3
Rsi2li51KAgaiFUPPWODJ6z4T3t1sC+n67DQlh3rF5Rl2L7gHQkjSQ73879JvJA2PDafetlQL1NO
1qJsP7U6bqWjpovrWxoeOqC9PKKEtRQBtjakebbch6r8Hx2avtbN4Wb4+oBJmQU3GoQx3JF6ywCi
LRHnC5dRW9tP05REePRmfrlu8DVp4n3PBLme55QNRwLt9DwqpdBoGZn67Wyg+oa/E1jgE3HjB2YS
4H13TOguy/zdGT/0de0fl1epNMPYs0iPjE9klXieaOpLlVmCVIxp7aMAbdezIhCSD7bgHRZBm8au
pmksCmsPrpEthyQsFZCS+6i1WKyewnnW+v2e+13n+Vb6HXQa/+wPeQ/2Afy7XU3x74JvpH5lKIUl
uxPeKhHUJRwvcQKtjFGHcLHem5hqymHXzrT928Pm9OdQ+7GL2ZnDZ5RERNok5n3pSlBIrfVKIbF5
/djyVi3idEcSN14aLuPWm3Rxq+dWcy0wqqyMGXTYYsJD4RX43QbhiDubhYskMXz5g3qx35DjK53D
qYaWKmDP8TTBO3CgFZt4mJFUHnqKMHCsUpzSZU8kOJ7Djl87rc4MoJmGwn3uGjc3f8E1Wl6Ti2aF
82Ni8NtlisfG6Pv3qJOdIovrs8PKfyj8F4REi/Y7H+AVTEs8SWjVA0IW4cqihxap3yZNEu6wtXi6
Tt5rXF4QRWNK5GUNl7KLu7wFpu0CVzko1rTGwh+IZ1UFCQcNoQxWxOU/mCZ+VV3HiPECKppGyTy6
bKLYzZGAEcEO9l51JbsndTDLgKPu0rcQGr5v7LO5EJ6iS8JaZ3lANuBhwRjuHFhxg1+MZsFgEDpd
gAwKM3CiOuYvWNce3IFrknOtuFvfdWjA/18BKB6g027OYVMaJ0/xtBgwsSJ9+9AFnBr2omGBzZNy
/P3tgsPQ6uZrC+Khx4MDaGG/mHjCpvNlG7BApVEqcu92yzQeUJPgyzqC2D9Qatw9K9vu7wySpLkm
04L6gOT/VxMPrDOGdn5MfXwd0ev6dh77i+PGzwMzFa6yJySOsdv3SLMmbHwkUlpO82YBbYgGnZlN
Ysl1q43AYOUOjcSv9tJ7Isuuk5H0QvklEvrYxecjFzlq9/XicYDlvWXl4bAcK7e2EQb3sSTxnGXo
yZ0EDikbm9e2tCJ9fg1vbqlnOL0ORTzYbU3M/wrwXPCjxvSiAVY08m2Ng/eO/lOvfbiKpoti989w
qRPxKu9M+RQOWNY+i3SbYbq3XcS3zzOVnZnB+YnxT/nk/e69fhpgBoR8iX4LstvjLyw1BdOTCoQU
zPn54Kgalaulp4IhZn3kDvZwZWAxWcGZeyYxFDfxgHubftBQy/sxzoMOpvhfA5E50CxGPDB/06mM
3/7vtSeRv7ud0xjoGbiQ/XM6hjmpn2QsUWwf49ohvYjn4vAkj46ZT/f+bshVfWAQSFmMXfZ2T7QV
eDXWCucnJLSmNwYJN4QE0hK0cqLZlcyRgRVh/lNPXACHKbHKF/mahllmHfgzZ+L541TREQcaUSIz
DDICTdMxali/S0+l414bUxGfSi5C15ykcJUnx9+KxVAMU+vepiNjumVQN9Ep/CFQXjZxYy5Snu5O
PFrYBHugBU3Y4cnjWMNH4oe4H9M+2VHSxpC2GwpGxGMeICDVOv7bhBQI7c5rLF6Jo72mbVhtZFXa
FHHzM1XCM4ZYy/JxsUYr74gSahoedSHuMTwOUvF3IrCRVGgijpaMvleP73yH/Y0VhYei5/mIu1pt
VBXhAYxBbN/4ak2eZ31wsae47ldIi+qvvLsYQTrjvv2JsxiM0jc8d3TjBe3HDwGq9RhGbhPjChcj
mU2xkmtoxK/tXzTm0CkLfrUbZdSSeg+NvLDVGewfZM9Inf9wZIv45aKcVLnW+a5CsHjJ60BA3uRA
9ei51gdmP0lpsC+u+TYvqSgsOOacbp5RiQug4GZwEyAFNVvIdSdzBa41gZWAlMWwXSJf1/BwA7Rs
5jn0nIj+HsF3DPFqRjXhRvAZDY5g9OE9DnfupgzJVR2yJ4/K6PDqXhNv2xHl+IQXiURb23UeaGAR
/YkKfvCYhfuzFclAkcZXN46gSgE9iETf5Q5pOVwIIQb8gqMixzPfEEjd3e6feHCZZLttDBR4Vxf3
Uz0MDuUHqaozVJooW6LZLCD5h4Hfu7lhB10aurD+e9sJ50xyqLqugxpBdURj1aUCVV24k9/7wqSk
YUsW/sCrxyn6ERj+hFvcVVV1qzYvj59IPYLiK65K55NoAY7IDrKmMdkUEBU26tVQCVi4rXuY1faK
d0F/4yBBWzbgciOgdOmXk146lWTGnJ/R9tu24H6/gGAwIj/HQYjxnRiB0PZ5FY7Ck0TWC4AcloaE
DZd4+W9LQeBiIwNxQsHzlRCOvEf5wHQRVTP8F+g/7Qw5711VN/3/RqCEcrr7Y6PNSFIeubXRQrlG
D1BiiFB2XD4b3+yBiR4xiUxjIFyllO95g6rVROIEzySqKJWAx1KHFKdr1nafKvpUcEz/vO5YyRWF
et54yOA6Fa7fI/1HKo8PpywiWDYENVGCfAWm6vQAK5VEOqesuvBbR2/Td4sTzwO04UfdLi68PKI/
e2Z34aD/fZV1HeVfXqoSxzbbAnqzZ9k9VcXfsH7c1XgQwJ8nH7OZL8wbNhUV7qvy1/zDl07EETe8
Gwpz8uom1ryYEziHK26TjrZvBYUe44ciIGR9mQFwm+3FyEMBY6CXJLXm5YiAisDtUEWtXlgkZkrI
Cd2dpSxCpzga24C+kF3pPjzLOIITLfguK2amVCfN0V/GrIdfgH3EFE1cAZ958iBLcmUmhvDfSY9c
E2HZMEsawqBMAoImpg/Y8GZxkzWK1MbdShyO7pH2oJ5FCw866AahPAsmfWm/I3sGd5XuTQWiqPVE
17/4LkJlhGX8j6WzD24GbQiT0710TYRWKuaTPhEl6f/t7IxBxBSJqeBwzoYh08PhZZ7sLQacR6kS
F/xR/bWuEDH7Hra5Y/OfFxGB2SlMGwOIzlOiu6MnehKdfL7xQAFs2agtQG/73nsfQeEZzch2mLqs
iZsJcv2Gh3hRQTtRm3AfWLswDmwIHCQWp6EZHIKwb6I+KP+2hUfvrkIE6RjAmeaQoLgpGhH7LMaj
5p+p2Kao+W5C2ZLxQNb4CToQsegrm3SDX1bTEQYKEMQwWbC/B+zF02mn1kXMvse4MSTkcfYh0a2P
hj9rhfbDmEN2YFhBQ1raAuGQAYLk//rxdMKjf+ibHCkTQUAUOnThwnBMB5HqQogFRkUo3xECYoDy
nnVKrbvcdoXfkUFNICGUI2Qo0E4maZbKxWkZh/Et5SpASfAL4epfZqOsaoivBktLpnE8yKH2i037
xm1gYg8WjN2ewaghlKMCdB+v6nGi2ozbaDh4ZDNGVvnUf5MxZlqL4LfexL1ew2hYuRY9xSjXfHU8
uzLKuuE7F5p4jD8vPQZHelrUi5xkH5F0qUrlhBtuMfUB6y8Kn5LnPB6sMY46ekXCm2W3aMwod6n9
J7wwhvl3bkd8UVoAMELjD/BWY8PQKieZyjB7yhpBv3stg2X7yBWViE6d/LWaFHeeeu4gWcOavx3W
lQkuzmf8R9HnMkXudyPEw3rtf4nRQgshbQ2rxpf4zxCdwVMC2xmDUZ8sOyYjlZDwRWfveNPTsj9c
suiG9jqlGJwbdxA9BvaIHi6luF6Le+HDo4nG/IIhfSyOD5s9s+EdXSV+mLXaH3M1drSEafAEooPk
D2fdGWF9DqdntEVHk5sUD7y1qEGc1zGAaccLYyf04HTquor2xRPsE80gmypoNylhclAsNV7M/TjH
mRFQBHbuvdArU6B1vnqeU86kgT9Rfh0ZacHxeAPE2fuF2jaFdhmrepds6NLtfYLR8JK7wH0CPUI+
ITguWxzvDX0hWB5ndy3f1C9QG4/445DaqVtIYzI1745MFk5A6CZ95euMmSQyjXIR5O1Dt2SEdzPy
HyLmIKd6TZTelyIlQGWEMxmMS8bOvKl1tKdAf9w1JcURmYYWUKnxDIWyRyBmdkottMvrme70KSYA
SOY3fzwIF5413DI83tR+lyWPlSje0OyVfVTGahHD1qav9/hjCkLWoJyPvfUEbExSIGiLpNr03S9S
mBWeBx8Wzhe+fzJrkAiksqFvsOBn9+tX/jKAWXDw58kNRYthMyIE82sP7soH1IEq5dbg8cvEB0C/
hIX8Jcgwo8n8lvFtpIhU7Tez0fY8AbnEiv1eIJlo1/s9qa0kI0izr7/EAXU/d6Z09fmD1Y/wLZLB
RHetrNDknQxBRwfuu+rdVavyNvbL4PRagGhIBDWvbt6KF+J4Gltj4T06m/aGNzJW7iIRBe+NqZh2
szse3VeW1yl50lgZ4BB53bHOpNVa7EvR+bTuuLEnMRDpNutuMpDZ4wdTXUzcJBWRBJkGTybtW54q
DSaQ0JDouSIzsm33TpN7hZ9+ntvobtuKTvc3m8GMdcgYOdTJ8HDcnXiSJPaL5o1w2eDwd49mr6TP
J63g4SFJ8Slh5P4dGvlH1v8NMRg8YFLoTr5T8BCCGYjDvmBUDg+MroX4I9gik/isWsiTfmaG/oNO
w+JYyjQYtDiWzkdCcxvKfhmB+uowyTttVnMlnA+B2DT8keG7D4z5Ga3BxxhoeAVFH1TE0addwmef
O8NklMsVvUuAeIiHIs5b4bTWytK6wH4wcMZveLOY9Po/fHnwzN9RUhri1TanL26hzovU1jtZrYWF
/WLT2iWPleyRHtuEQ53w+VCX+9jMZoV2uV5DnjX6tpoCG6ap32dzcq6KM7+7cpBVdH+MSN2qVth0
//K8T8QiS851Zb6icRAWu9OEhQX3+nFaLpDfEqyII4/2ycUMcKAEHtbLtT8iq+ctqJOrhIRV4OBe
V2utOvGOOUr1oIBqxQVWmYSp9GScLTi7EHSRQjpmoXGPu5mFycjoFkJbxh3VkpO4nPdCJ2FPHMBO
xy/hfRwE+h+YaGj445IPl/XZOhy8cKEY0RCPv2RU6wt27xn+35crWBMFDj2f3HsUvLvxQhc8dJo5
MIbT3KlSDedcC0Dh92ZB+pqL7ZYVEvZNx8Gbh6etsrFU1UO32TkUe2zZ2je2QYrY+CxSdNoG/O/F
j0epl0KDl5pIOGNa349MFE75J7YXQOzaWmRuhffCyUjxS9LZpjCmfqBjN0KAPBAxHFxpdjDo/kyg
t90pDK32Y7BqJ5uGREFLFAQFcLuioZahkjx/Ze/IHvGXBgAS8eqEFbuaPEArizVN2O7NIxQMSD86
XZ+rUyikinGTgc2PV2QXbP+qq7vDk5nsZlQUaxYcZKqhdVe2RJQdFj6GEbmT1gGtJ0A9qIt4co2r
ixHvfHauqiD8FQtacPqcIvr+G4pl0jaWJli8XlU0/XZrxhZ03tw5jqzKrAksr1/Rbs05eGcxUfh9
lxkhqxo8uqgi+f7p+qPSERGvnju7ofCIi7gOAt0y8ZXwJXOsdlJTfEjZvXguVu9xGPtIvNWX3TO0
d8YjF2PcR7j0SNVfat+yNfuSECtGrh5/y1YWA8DGMH2g0vnor56Vqww2vq7Mn+EQc5/wI2+D8GNH
9xu14n6heMYIWQ7u1MIt5yxXy/mO84P6ux57gU+nYy6ziCiUgZt/qciCz1mnBdE+ZUgUm7x6QXuJ
0o838DaXwWgwOZAU8d5XydVFXKWsxCwjIQRakgtsX7AdRose+R9RZYEU6RGP/avjvATnYbBj4lit
aTiDq8wsdEhJy7N2pPPdfS6BN+b6Jv3v3iJkAZuuHSXF6naK+eBjRPEhfd4Ja0laAf+O1udtwoPM
ehZjMgiaZuWzoqSQDDMUzLlTTKQB0TZPVTawG18zqngvXtjRa6OkE2+Hagr+uzJDFruyFZQipUEs
IhWhkUtEt1JEqDGFy//iwmqtHnaOi3GSYfOH/p4r9sTD2K07n+jQZXZc77Q+z6HLqMaswahVM83y
qKiOEiQrT2Tr+rj9SAylyjR/BEyNAeeqBpOGnhwxgVUnm7C6F4Wj6KEKqhQ4he0QLhoAf0sN8gm0
CRihjPB1Get99zli3EsZ6XGa1fCl3o/KnzhZZ6EPBRB/6qRJgmv5NcJMqlvOKinn1r9pvNgEsh9x
pRFTkKZ7ZkXe33PSKF+kVEBaMH3ZWsh9zvOyjvxh+CMiv7hTaXH2XJ/PE5KNe2kDbgxaiCx8Sl0K
LgCvtE+G98oJYz454QMva1uvZXaLeMrb2TUplYtIKVb28CDXbqmr3EJPrnKLJHmjwfludMF5VSNF
vqu16o58SXy8bN7Omg+FbLvxsHxVB2Zxsa+WPJCZuICuT+Bd5zGuhQL8xCRxAdubHeb4kBsLRfFA
+3c9ASCwVoeN71LaU8bltAk+jrNutgp7q6BnIK116T0o/64mqD4UYL0dWt1h/IN8Ol2ccL68zgad
oxwslgg4SSOORFpqZ6uIczHiNorHuI0OlnW0sVMFF3Iokwlz6d6oEj2+c//80s0IOAeLEedRtcD0
UF2kxS8Zw8dGA/NXTg0j/tfJId0G4CEOPAAoq+AjV/AW/YphnX7awXwV87u/H0nEFb8zHMD1JSqB
9qpmKjlMd7WDznVeE4GWQhYHACxOtNvB8ymzgRGvK8UlHkFrLozqDtmRq7qE7EFIaB3jNcRaTQsC
JOW881fEGQELchCL7s2MSxYp8Z4LdRoWE0Fki95lZ8ZlXte23KE6C/ljJz5StLmWbxRG+CbAAFem
gGY5JOJU8KwTm2PHQ6bRfCWJsfTFWQ6haZEAWNgc3L6uROn6WenPDieX2RkYcyJWrnLGdAaYRGGf
+4GfG8Im8yd0txS1xZvW4Scw4ARvni3GAA4RIQhcsaRGUXWwzwu9vec73ONkWgeYInxqbglxQKF1
1PR3CQSbR4SiqR9FBCQy7BEF7q64fcQmdyaeearQef/Uc6zyVbxG3kogcXqdbkS6JPxh1x0a6amQ
GrMjC/sFtDijNcvk+zoOvBJhAytqkr5hAI3O5WjY8lcgsyIlfEoefkaFlo5ibcf/ypBcP2ZGW/IT
K9KJxFP/TVCubmo4mx4SdGm9VBD43heUPgrrsv3xdx8C8xFbxwr6FnaAXsJKF114fjBgfiCZ2Tv5
07/K6HPO9jbH1zntAPwHHjwoYlCGv+INfQA6iGVlPAjdAzaJJ8jeopYBW1CfjZp3EZhXHJPSCE5z
CesxTCswhQf1ooTAC2rAAVt5XGAJR7lqddzfqCrQ+HfPsY1lBPFmcLVHxEthuEzuTXPquMbQq/l8
SV2NaylBg0txHcfFYd61HiWbZ0n7Qa5AZNdX2myrAVvDU9E8RZcGmnvVGJ1SlnOaRiS3Cw5d405m
EmBOcX9nqKjTzCRCl7YO99R40J1uuXVzNY7xjmGCTGY8mIDgf0JV7SvdcDZkbTFA+jRISG38OWOg
bHyHzbsplS/mS4saGTMCyynfdwEsFnnN+4ZT3JyX9w9qgUXKfuKYQZI0uM+3m7OoujHz1jkzKS1m
c3WXun1+GGpyFrAZMwPOwFWbZQGxecNxY6hu/xA3QzJFjEbSQurkukVtv49djzM0pMIln/wOLSNV
/iRfP4CvYpXd/QCSrY9hME8YIBL3DHCdpsrj2pT0GMjBbDyEQgJdVg+4vuufyiemu6jnD9pT27K7
kUS7pxB5WzqIMOpBOHhMnrSDp1izXl0OhGVW9LYJN51zBO+zXOx3qwZuJmuCjt9H1ms9xdYZRDdb
5KT3mDeSyb5oKcQFVMPQI9Ik/15zHmD/WNKn4hXJgGWemHHbyY8Qh7/D4sxbNhAxdyZYeklPxH6S
5ut7Hm2nLUy4eGO5dVBXv29oy+QSQlKqID3eke0f9oJxECJWzPa46N3sgIcfbDuxs201usJHC3jI
OYknOWguID+CM72GiN908kVeSB/CXM/KFWoYkas7sJqY6DOXgn3Bfk4jH38Ii2QL59DcCheYZnqk
9stD/wxLLLJdEWnwfsOepTtuiMJSg/HlnmWPLOljboMEu0Cr43HgvinjpavmCI2h/vfnKmDTjuCj
+YXeXsD8zaUHfuuDkW2IFK1C2iR5thBs0LJeks2BAF0NTlRmhqZZum97lHUrXe+mQBVy4TLWkV+Q
/ZO8bsS/V6kKIWBCggE7kWx7KuBRjnnz9vUEtwb8UG3xi3Hs+ohMyoz5VhJ7uvYdTzOM8RkukMzX
iymheAtEogJV0uMQJwglQwNeW7TtAz3Adi2xQPASLlO3phZsCYlGKlioqZN1LU7hNHM5m2dQtD1Q
IRMbXYXIIu/69ct6mYlzl2MJEzf+qJGYPFF/sukP+TnxUSj9KdHKfQBtSe607CEHTFGqq+XNn5yV
jlSeJPCIAheMSYvSrpbIewGiJ/tO07nXYAWFNrjCgETDMYK0+0/uh/vQnENTFl43z7D1XnKpl0yv
2Z4JY+N2ZCVg70WMtlDgGz8MPFLbPD4D+BL2dfkkRR4Yl2tciG/IkAsk5ODpfdHEEJ1E5YtBcdyt
A9vBDWiD8dGuQPAOJsPIHIrIHGRUa0rYJNy1RiUtLxfsTIkI/RebzxBPwovc25iOq+glygrzxJcO
huW+bXerLpTO8SpOsdOUN+MlhQRoWN9ok3jGHMNopzOIJH9z0c//0ZPtfZGSkFdNCJX5nHXe1I14
K54mnfoSdkLOA3Zlxv6KL8szIf66M80/rsBRFzPXA5DnaFPhCuzL4LkWUJAoECLq+Vb+9G/tG+Qn
chS05R31Qw4upA8e6LD0Aj1eZBtURhbjFvGJoV+93upGdSJcO2aNFJRmuch0WhdAf9yQyHwV9wgC
4PFkSjgT3somGZEYEwkMYIDcYoUvKWS8cGxYf4/b4DlelUVJ0tz43FwzmZy3Zf2xSmyI6jc2DY+K
DvnqJO7UyHYqURjV6ukgO/XkdGez+55cKj/pr/wyW+X9FlHmxmykKNroM6sq8fLsaMq6x+3rLkbl
HtsrFdDxU+olLDLr61dtwJIE1++8Nu8jGOlAZ7sdeDHvCkJYvY4oRW3qmuTgdxuDNv/2ivNzyj8m
Z5PjLpGIQe+5PubJ/4QQYarXmWXCR13bWQx+9zjolgM0e9tJr6ks6wWwodu05G9jTFdGZVthU/s2
kfiCXODb3+U2uc1wdGlS7osZqZxVJOSy6v+kC9Iaszc/dOigvUk2PSVBxzR42Np6bReJZxODlu2e
6HKwOLXsCOIznjLJAFQz8+xliUEuKJDPpdsFUBNA3dO80D3nE1BWQpQ462WEEWzXBTycb+a52SV5
4S3J3WD+BDbBF1fEwSiaIiYhOgh7bAlxBVzjiK7qjMdZ0ZzfJsLwrN1dWnrjC/T3PoD7lS/KP8sT
kToAkOwHyZS2SeXlaYLQxaMS80ll6FohotIXWt38ixlZ/79l0uwvfXoe/kpu9jJ1T6daxwN9VJoi
Sh7pje4WEAEA1QaAbxI+jSKHdIjjnWVhO5bkgH2ntvCHupmD1wGRhTj6Ex9QVZotz35mFFWYG+ol
6mXijBNXHCdbiQdOmNeSBCzJSIwL7HtT95c3VZeul8RQgLADFJ0P9goxqnmDSeiV/JoOzQqEwdBJ
40BYCl4sMcZjPb17A8Fi+kOoipOmhkOpgY6zWuwcYzq1Gd3keUYnn7dK6q/bFfiyOo0RtK7anCc/
DKSte2WPo9XD0QOrw6rM0Jm8UC57Q6L1rT3MSV3rEkW8c88RDc+bfHvZcu/LkpwqzeWqDB2/f8aU
mzCZWBMYDabj1faxPfHUlzyQ0QGbz02cGGE/++PgGF3bCqyc6h8qZjd2PCBT6ojGHrPbgyWylvY+
ZNDEHUeXmpc1J0h13ePdEm9kczqDhKEcU8Wiy+f4y64HtJ1maz97LKXVAF2z8iWCY2AMCAOxqmjY
TxO7LIh17KG4JZSgLlHCzaDcIr2X1AyyRNtgh/VfG2WNvOqeqG1IOZ7s2a3yEuv/lfAQpZVabR0g
Y8bD5P0Jstej3UnU1pfDP8fPdQcFuG3dxANwkHkDvU5Y9b3nDp8v2BIhYKIKn4kGQfKh4MO/JAf5
4brw3DJ/DTitpBeX1yCDPVznOjw2RkVaVc2KB1v/XhHxwruiiUiOlgLW0YURnJgio5YDN1TIbDOC
G+oRWAE+Mqe2nLmWJ36DmG0kcRPIqlfBydoUR/VK1JHpFY8l+vuU9MsLDbE/yTRFwMckj4fLWEhY
2anXKKgw8hOIfq6+nFGiAz5UadmiAm+ya5UZq4dGbnJR12BIE79i0auWM2WeO14QpekchOYxZRSr
kclTYCAkjIOOEPqanzWb5IAMfH7xXjtlOa4W4kWJjAKYsVbRSVscqRRpOkqpABzhQCBDXhqakr6T
SX7RZ4T6XY99dSBGIEYS22QtU/C/HI1EyyGL9ORdT91Y53L8W6C2hs6yCb13MKRT/iXxNIdT2D8f
fVUQK97wNUzJd2hzCcqVq5a22qMNoe9w33dmwP1vv78C3rA2Rg1EORDfEmisWosyWgYH6RVe43oF
FvYHUTOEMuAyf2/PUk3gIwx1R5fmVGvd5k+91JIyE8tlQPQeV9uQzzRBHoJwyy5szDr4/xYym/xk
psw6BnVkEn+eqbraZHAwgywm/ZIhgK+UL6vFwbzy+w6APfaA5oJqV0hZkIgf+LImhe3XfJfjxDvu
WYwBfJtH7QY/M9I+JdFjtrcKkHXr0KTMij+TdYq5AQ/DYeesaYXUZD1JO25j7A4HoJ6eE1bz0cgv
wLJirkzs50f0Yq496qJQSSJmTtqlPlIK6LVI8JAn+o+Egbo3No+R0CN1Z4sHLEgvqfPUxlO85eyh
GjPSWCpPzCpjyTw8oz0bmIeGfs+Ci6vTn8HnqfFUJT3zETdsmeVAknF6VKlecqWwnySv00vLeBjc
1e3V/TnXPpGazM60mWm7dyG3lZm+gTBpoDWYz2HY2cNbnIMGd5tMAql2GDNBnx9g9/YI/EwBKn4b
LUGa9V/BsE7ZxJF/HXUL7BaRbnRJa/nkBVRLrsoIkqeccunnkR5e1MJf2TH+r/HWI6ojt2D7BtJl
146Lht29sdj1pvG5aAZUFuYB4dkMdnLM0vhaFVdseM6KGFoztMVmSmYx4XAjHWey1CX0bIh+QRDi
rozl75vSjW5RaisnAkrNv9cnw3CRVrIZkExTEWrh82Ir3Qh2J5ZpSguepWvpig6cwJiWlbIrjLur
BbLZo6sN0QtnliMkz9e0AuySRttzEEq6hN7L4heasT63c42GNZ92oJdR9pB5M/QnJvMbh/+LU5an
L4sm+qvwmVdkesGt/46eKLIqV4NJdaP7dGqG2mvJU56KAdmysiQCS40UPhThMXukLa3heWrh9Gsq
UeQ7JRFcGP/wkrMDedkjOO3nFxqCILlhaIqb+vpGDuACh928sR82d63ccAiTbmVZWA6ZOI2cVtUh
UDI2g/tAzkpj6jRJtWbUjKbHn0FpRyaGR2wQ9SNU48fRCzdPg3iLX2CkEMwpMg601aHNmonB+wqL
QJFnpDUHJkPX8zuEk2g0ZKr80Jqzo5CPcHULLosOFRE6B1XMV6XK0Yjpr3u/N7P2BmgrSAA1tVft
lL8uLqwl9601JMe8DhhztRrQeewSXSVwin2NFwMeGYV7ibYsoWq6+LUwXOVBguMfEln38VNPVYD8
cz1Dscu/aZVkyCHxSWQ5iG+coqCEGKYC/1bBnY3p8oIhRQwakQTiFV6HUB0gLIFQmYb+1wHGKv3e
zfjmLAKSVrTy+WaM8gTjFYQb9JXEVKhJjf5KCa+ZsyB01MFqWn+fX7VHLDKYJ4OV699gpdHtaCov
sLPV4kNqW38vt0z38r+HBy6+RKa/s1aiZfn4ue87e8TE7wSiVRzeAI62ql2zUl3AZ8scFVcAlc+r
S2HrkF35srLGhflk3AJxLY9W/u2cX4o1gAISXEitCXcFpJlf+v2mca4Ts302Pa18oKMEnY2EIGNw
/4pdJdvMHeP/No1rhyWB/vt57H8xfLuOLbkkFvxZk2M68IvVxBlXBnNOVoNwe2lYFJTxthXInQhJ
Wd4hD7NHPJ4PtCS9qWqgFewjKZXn9Nq/9ard5QInvfTd3Ukp8w8zUtJV5OenlbogT76YIZMn/0Tm
AfPjDV0hz62E5HvYKHT+YNvsamnrAKwaoEbJJk+tHy92UbBhZZe9Q7mARfECt7b6Pj+N5jsa58wV
a4a78gbHJZFV6kmv0O62lMiER9UwhiG/Kb4evBsoDn4HHbwTiGex2uQ+DmYmPhYDXQaq2bHs/uqn
EXbW12NOAzJMV0QeyMOttrXrfxgGGIdEvO8uDX6QhhZJe3OvbiemOrRx8vxc7U+uXgA0bWEp8yzs
Hg8qg8I3vB2ySnOvm4UHhQeEUgOre1MeIns4s83oI/E2Se1QKFKRRmDpw54uRzhrjp6AQXtu7AGn
z0C+j1lry4clMToM9bLhdVM8QnsTV5HRXCbBOaZgH4vjWBcMTAG/qLO2g8qsUbQ60FAt3NUwBdGs
giNsSMH/cy51TTWo1SxWElOwBbt+nydnHy9B8g4J/sDd8qGivDaUU5oUWxjy6tC6kV1nQZ9Z6+PG
nhvJhZQBXtW0QbPb+XqsibQgC5I0B/RaOgbQQ7EGWU3ciz9TmkPEcOXWDQKo+7xBZvZIqqNQEt6i
FfbG8ElKJxFOe6UFuBGjB7fLb7CTappZrBKt0LyGN0r8nktqD1YFEaFnzW2fO3uCYo8yN/9fyi4g
j3C9AmX2gsdKYT+rU8z1j+9jGz2ORq7BlQXtkhUU7ZpbKnlGuIIi7pUH+qj/4gJ95BVckRuH3Xa3
bFcQuv6Phj0BCJHpvouZZLwz4CoQquB3/5WWwXBwtEdG0iOJ7cQn8KiUksogLYK6gHuV1QokRvRH
YgfuO/AHd8QfFWjiGpCdD13fb2xy9jeO0MbKhp26dw3Xq74VdspQEgUB7YaFV+HLmRW2mhQcgJU2
hE/OPt4GxN1BFLiSPaqPqgoBEq7EaAdpuWt3Nl7X2VZN6RMJkQm/SGNB1Y8YDLc8BuIVCv/gBbT7
/XaljGJIPwqDf7hlld0EQbqsXN4GFxuuXQ7aQ6xrE7qByjMHDBva/bjyTFXMS9wE2pho59kdffh5
AK3XFdUWVNaEyW2gE3y3B6+kTG8vuOk7AFDDKz4k72uAylG4+S3LXwyfArdSajM+1ps+N5lYiFSw
lEX5lyPK088rj+Y7OzmQY0t28PIsrTA5SLNfMq9Zb6ffgMaSTfouSLnaCfExEfNOid2A26xAIUfN
k/7pLLxqX36Ajav6vtJ+aynxJSzG0E5oT2Xxof8IAVwpy70s5ztTlLf6dekCbihWXR2CUXytJjiF
j6sM09imqImdHCDgHCXnkrvRGLcu6VFIfoZHcpXiSZJI/vT6au+HCnpQHwYDCYS8rtA3mORwqsnu
fHxIWZ4A0Cu90OtBvDbNrqlVvswQaxMVzhnRx0HB8p98/upZhhASt/wbU5EbBP+D8LsfFl/Avqu6
Y7aOHqGrP9bDniouhL4iVaqr+Pt1TyBnY5LGsiVsM6qZyJg1FqWvyCiokbcWrM4KVMphLwWbmbsr
6AbjmMNymEBKRU929Tt8l+XChaRM60HekM3OOAuV4CAbQSoVIgGPs3zzQxG3ErX4tY4QfPxaQVl+
LVRijYW9fdyQ9LO+guGqCYUYZnduIse41t6DTsAgIFvZpWNpOmfq+PlZrdpr2+a0HMtckRwM7ufu
YtEF0jOs60ICEa8JQ1aj1JhtICyi72uhWLeiPqzNWVDeTMuzSoDT+lSm0u0N+ciQVTVaHfUTekzp
+9+JEpXh8KfKehXqWpHWdfVEwcb25J0ywcuFEVil+ZDjkqs/l8jfOo1HaWuAq6nDQNKmBZHI/TeW
WbCghtNZ6vZcs4tB+tIZKLQDGkVfbcX50d2n13GgUjOlNv4u3dxi7NnLx8G68upat5ac26Zzqd14
f7Qj+PG5yw5bRrgRkVe3tvmPi3zuZPzhGMUAkJmRoFDj6lj+O5ZpdJP7IEl+99J8tAnCwUKvenvn
C2GluUpmpvajfEkRATQN22GFuuFF35RC2RDq9f+KaCdylQDs/gvhRCN6+X/Jo0sIDwra3cWa6MoU
DSxp7FMCsXA5qIq8VyjP3fAX6yog+m1oApAiWMwB01y1ZxwiCRXR1DFy5wPlt64WHn1r+/7FLFIV
0Q6vD/xe9wkuLWWYrjFP9CmvXyhHAI9tN46BAQgRYC/sgDokEifo8iib32vlRtiGMHnM+o4t5n+p
lybwMXp+87g0qSwlcnzyor/MrNusdnenI8yX4I0oplZeqDqaK5nTXO/vs3woRsUjEXzgkwqsDIxw
fP1pF+xJjL6ooBYRQe8EtyV4boJHu/BtbiW3Uz+pPn5RKdFlud7q/oxgTgQF6X5EdaAstQLNHEM/
ckCiHwDHQyZrPgLJqMCM5jQfShZqiAgVCPWIQdy2mA/zvYF4q73HBQgElK5NRpT5CcqV0masZIt1
Quuki8RL3IyyMCtPbbSV7nVH6T1+V0gAZx4dAYw2OvvgsqkXUCPOo3bFRoQrU200oTK9C6A8gipz
0e+UikxfrzykjqATG+lhO2w3Mtwwf5hDfp0kFGoI7hZjNB9G+GgoH5AQv/Bg+UHJO/BEtDkFCADh
1PKyvSWhuPfmmN9yQxJMwk7RjFSskaCYxwJPHJRBjE5ziHIsHfwAjFsGdjmaz/YARP76FokDlkiS
QjezPdGqmZLP6sxzdRAffyttstPnwfhTgs+3kDa8IOHWk2JGgJ8Lt6U/K+prf3t4a8eJF3GGiyT+
Mp5j9iLaw0d4GzG742PGZQA/5rLBsgJz6TrHHHiL0Idc6TNarQOL5JwulqIbGXPOaTqcCTVfTn6G
HpICrubRvVvW9Gxt38K37GyxvpPVJWHkjb7EKoqWu9IjuBC1rjkD5RKE8qcm+0s6JQkNQh21S460
ikPd5GE8cRL8VodqwkH8DZo8fsBbI+igeX/sCsl0SvobD9v12x6ZVnH8mp/Ge7oTptce7Ka3mASi
CHPtFr/MOeyDY8gUX+F0a7p3yga91MuU1i+m+xJYmeLEDyYoUZhdQKkPWn+/7sp6csVl//BVv2ZQ
f73L1a7yTQ6TSSBrPXERARyNMIgidU4LvecWgKrMg3DGmfAP4r12rkYadx03deILx72TlwcHicPk
mDNvA5DR2G1jI1VJxAV8THkp0OqISgwzl/nto556f/y17BRIazyWexat+/qJRyNpX0PKMcFjgRx9
Sn2NsRCTRQgs4bYm37fUKhXHGTdQcyv5BFqgxZNxndiVTA5bRR302OqyV/+S+1g43XYZL2OxwBvV
iRy6HryxkdRJnjhrX74pAqesuaCJUubcWkO4tK4yauMthnsBh9CzBcrvMRskZ4PcXy7IbZLlOBYq
U4SY24RW+tpL9b74R6pilaj3K1J3oGiF33Vuu5gblGd2HYSh6HdGoQqxxmjX3isKMMEjbinI36IL
SP6EaEcIFCUqfTORJtzGUnb4E2Fpuk5VRcxRf84EU3a3mnV1EbD6EndA3DXHQB8khFW/5D3ch3+C
nfbtxp7HX5mE3PIEoGP51Hzx3YTOzw9DxGVuVdwCOFFL/1EKBuRS/0jQ5kJVSi6WnvxpmPZoaCns
KrFBWHLh0WrG+3LCW/vKiiWH6T+qTR8UxpekH2Gj5ZIJ0ahHCA0OnMfRhwvsj0Q3fMQTThl7OqwZ
xmUjjeSn7R2bIxz61U5QtyjUxKrFWVikE84olF/QasGYZIbCiVvZRL1sW5d4IiVGnSfEtShVAVdD
VHL4/iCD7lIAEU2GqAGpoLdrlIAym5pyfCtJ252tmNcp1k0rl3h6N1mYAkh28w03iv1nCL7S+kS1
J+VW4mvw5KfoMcJYmtQIrzyjLMkJE2RRT82gPbDMRJ3Ztu59Er58YxzYXMZY8adul72CnD3xyT3F
sh/NSvffPdlvaSPYEC9nLWt0NDJ0C+axeRu1xgZr1SOoCvwEdq/uAw+GaO+2v8s92xh9nw8OIG2t
bYzMnjfGdhKttQ7UugJSl+J8+qYVZBWHzyCLNfcqVmmE7VufAxze8oYNxFIluWkHsyPg0AnS7G++
kb3Y7L9ibNH80uog6E/UIgih1t4Aeb5a5YvbtF1MSPFgJE2VWfxk+zeqPGeXKL1y/S4+Q/UHUbjc
whRU80WNRBSMUQv3YnBq0daR5Gew/RwlalI1g7Y5PPHnwm6J8gkkLn9M4ELC+IGjTl+p0g3keLJO
aN+a2rdHh5K3HR9C+pY+oAuqP3eZ1rZpNX6+RpWX+y0l0Y4QnF0106/zp/03VBqnqsEmtleWS889
nKVQjjLQh4H6RC05TCf8X2aq3pP0AKD1l5pKi31Zl0Dh9d3xj+0SKxvx5GIlJ3ezHIg1YtXBrrFH
DzczQ7wr3Fy7kHUgXWRaFVVfDDGDqEaRe6sTLuz04XE+x4i0Vx4nAQgBESWJTVCuMTMr3ep7vKeR
4Ao0DEMPMrIArtnGYwoGsB0u1yW6vICz4x31jrTelFWPUm7/KLj1RrsoHTzSDrGomVvA66+WFC4W
6zH3sV1prVDGgcPlOGl6BUgBJwElvnaousBbhw62tqpgwXLhsLydnNL+aJhUSKDDwJa3BABoYK5o
Ik0AhW1c/eo3IdwEoDJ5IWJZp07qYPnTe6fwV8uY1BjISRtRndoa8wBCIvvJfylWGfKcdVL/22m5
IbfI267Y/rJLEfyZPwuHtGTbYaqAVs5CuPA2QxBiSPHvQvMYM0H95yXjkLf5EFtdSWfVZbX126jr
O6MLovkr1FwHxPetuy7lJif6gA3RHveWaZ4Qw1IG9BHTE1N9jbNYHSHZbBNcLT0nb0gsLyo/ENnq
Ijo+hxYUKP6Hp/mgZMX6w3i3b13Suyb+vYEHcNA9cAVqF4I9+qCy8iKRWKdnmZUude9Zlbq3I8h4
lRUIV1X5pbkB3hfTZle9efOdbHDckXySBuE/MCMyOZKNN3FntXxMGLbs2p5rIBdpbPTssvwdFJ6P
bAMGO87tDkWX+OLHSS5SKRrffmQ0kjVPQ6ctrh/ysdPjLPQQW2LEY5G6vd1P6Y8mHoEWfP+8YNf4
jeFGA4LBL1vvq8sePJpiyKaK/isvxX3QngF4veqkKNLvjmpNJ4HDeHkHP+IhGNLo0ZfvPYwPurld
L5QasUkpdG2YGbae8FXHnwOcT/ANUoxSJATp+R7vKwEj0yAMg56r3Qtrk6opttohp77lkrtLKICs
2AcgQTGn4iPlDVpBBBBKI8y2NcAiZVm1mpzDOIHSEcZ58EEgO4VUbeokHeUIK+iVnJm6hVc6riLn
qFWX9lrdUHVRQHCwy9lQXOm8Tq0qWwopaJEIbZqQnYNE0peQR50Bu503tDOmejSFUgDa8D0VySiA
H/X+6we2eVJVl8IvdCZ45K2B6j6cH/AfxWe64FHMRz13cYGRtulkJ06Y0wT+esoPpu4rqTqanZoX
OVIONtVvivsIcp/AUPody75Cjb2gaeSXJgaOkSFk5Cqxojz9W13yKvj1TcJCeR05/sP3yK145i+6
zjRJX9CkYQJPJoUUcPCbfM5lrSXw+KlcqHz/HqflKdXnaarBApSUAT6MBsxS1ZLPxrLCCQsLQAbp
3906av8XkkT9873Vptj6iK2fEbzO8sxKGatx2XOT5k2Sj9qlwGjaAiMDeaNWR2P9S6H9nLDOalcp
trzs9folyOhjc5LicmT5QcbkqhYahIHmfRiSuQXLBjVJBq2Z0kQs51PnQ3gczzUP3anXcumJNGQq
0DsMcnI2hpo5IDhWJxdJeBe6IjrWjwHCBRmTtOR2n7WSqCFiyNhxFSX5FwM/ogDSpuDvdPdtekfj
Ca0m0zELHsMQC+wn43nZbUFKndDbNsm1TPzM/RDx7oRqqW4DX36BWs7EvN+rA+v4tyRSQHi3Fg/q
Me6o/U/ckIxBH/30JUkGGQXFRrP7iSJmeW988EPX3ambfqrgx1Ky5LlE9QtxsCYhHW292U7vSDcz
SYHp/uK3LLF6J7ZGacheCO69V6aUZ6N0bpRqQdmNNWC8/maWisBLZPEtodqAHqNejEHkez0pUYUh
J4fIgeN7ObYLsnFtDDsC/ZI+fqCHoWnu5fjblGhMoIzBR5eb7r4DTN81MjY70Ga7Zwy85dT0amCq
fdAh9Ce7wueHmcORGY9CbXl8cf5dmAtcq//D5Xi6laEb67fOKahw7MKq2/KoRJr4G3rX3UjYfRDR
SLEQvbgSQ9dn8qLjIcLNg/tRRnL5y24dN5ukkBqLFvPFazqn62+ZiGSVyXTZhQX+Ir+Ce75zNxxA
cu3reaz7l3IxYA7VBi6u8M7JaErN9uVkB7fkSGzkXSTSnHImaGjdHn9w97qWDOsuLGfMtbBoj8nP
th4Sv9ifBqHxKCK/5RXIo8C2bnUz5wP07loAtQIPKDiXY+NTcw1nsqR14SC+Ud4jxfJaQHG/A7FU
pr6dpvr/3GwXksQVsiJBnNh9JPiHOaD29EXJnvClBMhSiXTazu7roqptWHwmTooz+1c01s4UCfk0
Gn2UK4VXGhC3a5noAWD6WnTQkRvDoHCil/gGItKCWC0Cj55nNYUk5SFXahTTkI/iUgyEK4pwTzR/
xGSvYQAiy7hcrS+3SOlNvknfamSHBOwkN8ILZ3jzfcgzxC4Gh8FoURT++nEhkxbdhe/jp1VbVPhf
zdFUFs5yA7ljSUa+Q2p8XAY+Bs0e215YOya5ryZx43220ZWm1Wl8t4aRpiTB8gmcdGItrab/JOD9
bFgSpZhnCFQbhZdLjISDqurxjiInyrl12lS+tiZ4hO2MG+Su7tdISw25ujriV9QPS/sdxb+RtqLU
dTWF3HxqniCYqolNyAyEHLDs9uGPEHWvJ1/WEvmjy9jJoQlYc8ldH/UBqUfoAPjkB5jpDF9kU7eQ
HI3eqeFDHaf34aQE2Ng6CbulDTTpr7bOfm0bMznyOCl1RtzfJpGPOAHeu71w8r6c3bG/snCH4F8y
p6lw12652WEA5ma9VXLrOl5pXb9u+a08AmVfVz2UsbnUFAWIpJ5uyAgtuPAINrGu4YHEjjnxq2rR
zvE4uTc1WDj2CVyTC4uaFC/tmcmXAEeEg4ctOjeawYFfVMrxcQm3n6osbEdCPqNaUWr9D5PlZkr7
HhWCcOq0rVsyvGNaZEFbKXgZ9wkkP+Ths2CjgtPT+Rs4vGg+TUZ5Qhcxn/psgj4LaW+lJUWdr4qY
kFmOuz8744aSKsAzesde7ncRIlqoqIxAT0EfuzlM/3RHiVBlsqOYEkERKkt1+z/a8M3IbbT/gMim
0g3sGP7jLgcNw37iGC5ArRv/WxvA8xOYiNRdpKRhM++uHAbDpI5Q4c/9dQ/OvSwMjONBWXk2NqHj
cw6pIiW61j3SGAO70FcinhCLJkZZEY2oHQd6KCg4XNeTFEo3XDiQ2NI7UKeYN8nCMt1JR0RmZUsM
nrneuRtoyLtsvsRkyl38UOX7q1zbb65WtzZVdLTl+Ar/bqHXy3/lLO5lFK136KfCKmO25vULABVv
daFoCAp/KwZjPk+Q/7sAtNURqLTwHAbDkEuYJuzfAaHpT1Wbnsk9mDJUjJx3umLxi/2rBCYTtJTr
7VzcUHkz+fLUtCKcLkPNXQMnygIZBXmdy366nBdgp4DYwo2PFYT229v3cJ96WARGmBzYpVKuVXSO
R4PRAvh9JePJ6Cbox1nmzIEvlVrrM0ZxLbZMMb5o7GQp3HBSTKmeG6TCicnp95trCSNhHtpRK+pw
6EV1DO37OzFCZdG4xHkXbK0VYLMi9CgjZrAkklSsp/coEwsZ2lj/C8E1FYqYk0qKPB47f53CGDJ6
E53bHSDvJ8r6QO3Hr2CWKgTWVGG+ISiQxu6djnM4ki2rtINy5d0TSbURZvHjoj9MEgsDBNnaJK1t
UU/qrJm2IYfmg68UjHT2BYCd7uur5AKvd04LdEWtZuRYIvlA5JWpPcGpovOkM5svdqWOGpoAnn8B
K39mHBUY+Ybl6AmTq4pg7p+29HNdh9kh1TbwBNc6cooSld3WW5PCsLMtmRnvMY35Anv2FbFPHn1q
wj1RA+twHTD6NOn7MT1iLC7IfL5Hu4MkscwSmDoMWqN8gSimd/dwYPn8aQMXVkorICWYtGsa5KB8
S0Pm9WucH2IoONvYSl0et9OScakWNeUXtRSCG+Nb4TUm9/R1gaydhw+Vu0+xPyw5Fyxk8fsPjyD/
VQ8PiMviYNxDd1EOGWX8TfF8Lf5aNCfwsKSGElKLcfwE9Yt/StZ/0vEQQAlgbFXFfMr/1N7KepJi
kFlLQLJweXpqyLzvu+dVdh+CwST2zxiYI+AXtQVH9jPb7QB5e44N3siyIk0l2pZNjptXSjEgMIGa
UMEGkkBuz2RU6HdSjk5Pb0OsVRAQ/k03T7ud3+umUl0hU0VRYlMI0HpNhlIt+mNOiIoMqJr6IU6v
jMlhMxoXwClRqHlYytK8Hy8PDdbzMaavj2VHutB1uXMVXCB5HgUgkyCoDyhvsLMJslYiOYXAkw2I
AsC4UeZQA7EgETaz0A/o5wssnyAFLxcPwqzCodEUX5CK1O8RNuU1ibxplOIipGHQbr61SyTdhVIF
/5j0Pn6pCL++v/RGgxez1Xsk9iNL9g/i+jASLsSAe+RKKE1rsPINF5rKEecO2iiF5g3OzCUFuuB3
1+lRyoKK1l+f+H66h19zCHJ4gNeW4mqQQ25QEcbh3J26kxRseQOXjkdo8/DELbDLNd+txyVEQHNG
nh5sadr3rgNR3ojzK6plnQwycVpUIo7+Ra2Kfo0R9nj+dZrC7sTiMCBCJxOKnHEd38Ho3wE/B8ec
qNI8FDmxMQCg4rPv/hy9NiQHT81qwDwnSY4Yt0iuIAdds6ZM/93O4gBU6+vYq1K2JfuR0Z9LhP4m
kLT52npdghy8jnlPbdisx0JGBrID1NJdbKrhX2AVPrGhUcNM9Y7gbYm3xNGYYK9if+RdYnNt5wIr
BOSjrV66Z4VSBgJRNecmuYev0Y5EahmrLoxpHDSxb9JHXPTcObqrlIGQFBAcwVpKF09dG5LrQQj2
GF55uYs1v84K4saplatipT2rWQ21sw3fSADZ6cXq/rHK1tmuqo5mjaYG4GFCPB0KG8HAHahReI1Y
SZu0DwmWIzE1z1bs8dIFyC0Oyyu7cMFHP5EpTDb7L6s4MOH4JeZlGDIUS3y2klmzIFbsnd0ZDrM/
wJvnk+XQRY+X/sq/L/vPsTae1cMJezPWbtvq4sZzjzyJbgGN04Bq7fkIkfnEKDm9pqcAPrI3Lxtv
PuGUuAJScTn9GnXl8pRfJSlX3hcZeE2ldcDdi6O2WvUAYtXmKSefmHaFD2oeCGfauEluPUqJ6PVM
HCrnWT9HhxWnl648I392rwEMUflC5mtO1pNF58qfO2v1brpWLByQ7vhSEPZka+j+CIt27dfst08W
hRRB2cmhCM3BqfuyzWuG3IMC85ChG0JjmQ55QxEl5+clo554npYhumXTBv6z4gioY4Rt7C58lk+o
w60lBOKuyrDQwq069DZm4TNiSUdMukHZBOk+qQ1VCsoeA92gb2a+8utTZ85SoHN+Q/KMWECsoQEo
UQ6oKj+zt+gOS3Ak8/AyZAqcjA4Pta7rs8MBXEL9aLeFX4208cNrIwObdZfeUetMVOIp4JSLa9W/
wmggYlIEvoPF0RExWphGSkdr9w6+S799gVPoA0J+bF/LDPiqlHqt+9VVtiVAltDGgsDXtcHRTuFn
Zsw+WTPhtXoqpW/2nKVQo44wmqJWcvqrmbrZc74Pym9UQvw5Vr/NQXfTD4RVqz+RW9ZcDJNiVepv
tcT6FaMw7V7xNE3XnxqSYajoExqbSg7mKjRSYs54UZAYGdkThXCbrGyZW2qxSOKvpuTmvNkuMZge
mlxi006NOPT+JL6lzHD7/0BaSckB//Ac1/eskCPDyadMXLCYzInY04/brzjtSVo6Ts+Q/MZbM+gU
H9j6ESWao9bfk8qQqiRsCxKAC676gRROyP4yxt1OwrWupMEH7sSd7n0O30eOzC2DICIT3IrqFLb8
zG7aNT9XsaS9gz0yV4v0m1FGFswbSomeAYqPjAf20DUMjHfsbGTEY8RlJhKxOaQs96TbzgJP9sgA
zQ+TlRG8+4pQ2ZCWDJA+98ZXZwuu2HPhpmTFXRhgdUuziT2lKmIoyBGliOvlsnxaHW8/UHr7Whf0
bD1h53O0z1Lcju+iwtwLlIa1cFNpbs08dhsdj7RWKMX/BV3KKumvjq98qwqOf9+zomazWAeqs+zs
Gy9TFjXD2BYjeWdNHBGr1CwtDYzguhM/NTSc5JvvOSzc4JoxCAVQzgT46lwkMjiKXpj1nxz3nk05
jd3nvnHmZAjRhvC+4rgX+cwdreiwS7jQIEHZMihio19w9VF13neVy90kYBdAhT0SoDTPexChA0Xo
AifF0IiJFg1ngvo5vJdvIb2blv912f9wLnHDN5hjJPiWWCYZfrtHmkoj0H1uE2bQxi1prbs2VH/k
Rgp4MoQkhcqYLX6rzVE5Doy8oTfBCaUQ/iWKyQzHMbxB7lW/N3od3TxJ+TzB3Ol/YJqU6psqJDK4
gRRzAGrbzuCqfx68HUYimUfrbrk6pGCBpvygpIDysie3czXGrkAY+pLjuUo6ojqnYcF4svUd6qkZ
zwwJokNG6haEKnwp47u+jZE8DBA3Ye7T9yLTbLjLSzmeJi+1egqvPJk4Zly0AnOwJoESnLUxzOuj
k8BttoAL3idmcmCvx0qk+70cKRDO/1mu6/Hqzm6YL7f5OvQrK5r7d6fsIcFNWixIxZP7NPIYfRV8
SBkXnAZ9FPWkPis7PKulBsyXbuvZDopw4UiiNoH6K3WbnwRl2O0WMMKmJ9mJnFgVt0jXFk/LEEhP
M7j+sqWQXqCHAkMh/9fXLXebQI+ndQjGmuj/yUgFMHhTTpX0k35ephGZ8x1Y1aGJhc78dNFGsEUb
6bkuJPA6EuINVQmYuWSM85mb7EiCVPfNSztN6GfkZgk9hznwf44cjDq6Nd72qULUmFAjrqXuiMub
4aApe+8wQkA/al6EW3gskGJUh2NGmk8BpjkMkafQUyoKzRVKLOg26ZFiyoFR/7HaTfTNANC8ngZI
ZHYO2GXFWeLVUwcEywKe2oc9ZM9MOpdvRE7S0kGL/+mLg3Qeg0+3cYe74nJCnp8BJW+UHj6xJE2p
h2nLq+xo8S+5JMKrxNaO4ic8tsJtldY0ZOVw7qY1s38iLeycNm7wULguokgtwV1VUZRxu0Ah5vl9
F+ufy54ayZJu4PvVub3bBW2KXvB4/G9z8QlP0gUps2P80lZGv32luVB2Pji9+9+/aamcSTAwFnB2
JClFnZJRy7xaKnE3ENOxO1BKnyZ+xnniiBQBfV52atF+/JQgLvg0HZg9vA2w9IL81ZxfLQpO8e8s
9XjsrmRcNB11OL37waGtR0rfJKngzu6wW/02qfnGsxiXUpsPWHEkB5arG0hvx0ygpKJ8WHWKcDec
gN8xsr4i1mB89HQZPsObz8kxVaSr7MNbE+4QTz//nrVIlt5J46gkrWvcaMA1HQHzj/UWGOhkItxZ
mWzIL6+bBWzIjTHhhK05lzsDpy157cLDStFQyU1IgO2Dtx0+lzey2bhLH32f4wTIRTjOJnlgq23O
OIyBqGCoKLFWQr03vr53Uw9w0g17ESHwKURpejcgSQen0rCb+DAuJ9hGf5XzeUQDzOFFueSGe7bK
W8CRCB4JH4yJdjrIReQ7r4tWRzRrcwez/io4JFMV99/QYEjUZhVJYS5KLGtnXqLGYIyiPihpLt7/
+4tx8Hg0siuEQxhBdd1/i2YO1ti/Dcb1wSbRsvjCH0YJUw490Ui31ztVvTRRww/LOZatct9Sx8cJ
SwkOegPSAtGOICiKIMvc0zlGsmiWYfxBcfz4CB9U6D1CKj4c+73b6C0gw2v1Xq1r65HXpIzV6/VZ
ujUtPhxGfkmhHA3Gc/i8U/GbZ9DW97Ml8OFb2G0eKRYM2dompPnwqs+iQeQTOvhz7IYFIONBKaO6
TLYiog8Tyoclcq22vEdigCADP5rK2Lc/3w2sr4f+QvcV+aJK6esUuQixjea5OaRrJeE4egdvT2/S
re/5oopWWeDyzRxZBUfmQ8A+ypM0NCHuD83BKeuugPIb2c0q02h/heR+Ppcys1Trkf6TkKs/lBhy
87TNBNCdEE1ZHKACFM9fpmENClJ4FyhmSYPSgXl15u+2iYkgBuk/u1s4MPr0RfWXdedIuEgSeKxz
uZxWFBFWVc678HoRQDTBApK4mET4/qDZHrYIyh7NiKjgZEHxKlK8+y4fCTxCLYFj95Kp4jWHT3Nk
vb+6cDw7nxqTlWLYeNP4fxBPssvwOnL/jyWTS8SScZ9bFdXgKCi5R8H8+S9/D6oob8/DFm4a4otg
kJ9iM2KELU75j+Z84XWso9HBycrmGKr4HykpIhrC0VW/tMQxObeWiamIf4jmYt87GcpAXmn/niS1
ODzbdjY1Le+0LF5HCiJikTeHipg5yaC3C8wF0nJSnxZ1k1G/BvCgzAHYQN4imHdTo34NjOS3m4Sb
NqCW0dKJ5b3XJHS5F4jhQ5vEGxE09NQkxD4tkVdMAkRDIUITS7Zk7Hqe9rJ8xlpL2uCSptNG84SZ
Rt35yD/iadRbYncf4JkE6jobXAAHUnbY5kxNB42+huwS190KPlqi8pVGGknofZ/iRk23KXkPUL9j
wMx4Zk7EnKpQtPsW55vZNy4xym5B+JEbT5K7kvxQDtvhe6K8s9YBLLis5NDngf6yP5mUwnU43htj
QNV3Iq0fFI751RceIBm/hszarHpVXjpa/JOBm6FgK67Qbmq83ReW3XVpceXQNm4aWlDRJAGDu1KH
gu9Aihs8easHWTcdW3+HrKQzq1eQzWwS35Rq/xVlVjCFUHeCpRaGvxloCsT/Ph7lOEmK7SXjpv1z
gxofl2hO20hpKQLnCm6kh0/ICsa7GyCpSDW4t97rfRj792rLjGMXqCBHqjg6yy8a3uvpTOQH2f/R
50ryYy1WQIZ9Qyx+hXbdrAKBL8t7AtQaSAIN4ZdjGdbBWT+8+kk1E1Na1AW0FytVhX3cNGVLsqnz
Eou0zdiwjk3jq8SLXiu0zJ+JQ0dbEX6dXsZf+iCIuYcfiexwcQTibQp3IoGbdXef4CdviFPFQ9EK
4C9E0UVUj4e9dG4ZwlJdTP+JIYE2NC++d7q59GUJeGYvAOD4fVKCFLEueCr6XdyxyrRdXAbykdbr
PXcZ0H2KQjM03DcyqQnkyQ1GJlDUiSbiaflK9ao0PSyamvdyRVG2QZukmYuk+LEpb58fQsJwcIw5
pk3zA0GF64B+gMvg6uvc9Ud+/zylO8gHt4AdDDVg4UWpkus/WDwE4+QnKZrjV6m64jVtWskAUvgO
rgysT2ONSydyr5+YGX4aiHsWSL8mOGLeGjebqX9Z1ZcrbCYkvkdPe0hiiJwEunyyygbhzVQf6OLL
WurFKg2iiwE7AzqXnhioj3+pMt8KkA92GeKXY3WWei1KZ5THwc0Crjc9gUHltVE1KywBZEQSHooJ
wsCDdxin0ROKqZsuDwZW8a3Gu8Iu7eIfMugfFa9SCHvUIRgoEYzsYFSU9yhkN0TpgPaMhxSlsQXY
8YO8QaU775jTpeUWboI1atYaeyOcWnaZKP0Il0qKmxJamLNhZvno460saxxye4CSt/1JWalp+nxn
46p/kVn0Jas+sVz6TMUxB0JQJ3KqQj5tbj80iZm3ElKMOedyH16ekPSytfxtvdov3W+rD8+Ed09v
HM9EIf/mE+GvqdxBp6rpqG4FrwIL7SuHryrgIgQs3hHkHhf+W8oAoNvHKEDLYU1xQnb1l4q1BXng
uwrEKL5FwKSHhaU/nVQFkt3kk9CZVdKI7u5oOyUP2KCt0r8G9w4vmwMpHXe/W55XwGg9vgS/+KiB
u4XfnNvkoLDCduW1HT8oUnnXmSR1RmLKMugku946tj+tXVlz2+rrhxrZd7Iv96iLutytDpAoQpsW
YF1vZFQY2sV5O/fu78Y6bky+pj0vxVp+nj238+eKovbJc9sRrU2NxP88v3OLA+VSGjr9GoAfWKHq
rV5ZZ/g+X1Knlb0scGqCOIrClhLo/Pnx64mDmCavqGV63tDIdgNxNVMdjhaYGbhquK07ILnR7css
noorFoMGWWojgTEuXjURDApzb3SWj+BQbScGsGvYiVC2s5EoxNzPBI8vlr7E+bpFWsT+ZYVxjBDZ
tDf6xeNB9reIBZwN02+rmvSJuvV3v7mKv7mBE09sc/8KwC6xg5E9BOdZRDgZ+z7UE+TjZCE8klUK
7fbJDw+G9iVKsW0Ju+ykFHEgd31yEVn8B6jY6gBSaEk0oSEmy9vBukIBilg4amnvdKIXYjdChKT1
eJvT/3EzGSI3cnnuQp0oS0VCq5KjeORoKrjx2WpQDmHa7sb9OB2l2RsbOPeS9D+yYsRVfWPTJNAL
f2b/ghs0pEjUE53l4qthSEbvnfqGBZ8XxqzjgfOKhmzh5Mq/I4Za/Pzjjr9xYrCpMj5Eimh/WqOZ
Z7ovMoNfYENvoncEmnLwGmV+FfLSUc7c3UADZ29t0Ztn8cn+DQjCwh5gOdVqXU+RfqDgccOLRFy4
a+74llbhKhXrNxA2ObUAcqch02eIkweBl6M8P5TfbmzqEPavukCdALxRfoYY1kqdUJ4kaQjntKYM
TLV3LopgEW044yQxBxak1r018XU5R+PQOUD/Tsj6HEDs/2BtuXMa0XvSjfJEFT0M02FPClEC6k4o
VZ6Y3UOueNO30OSwzvPnDOJaVyvj2tPVENcKLigOs4tddQ8KXlWqqoNBinG21Y9ro0tCO95jAedY
UCq5PZxT+yc5y87zPJ3aBV67v3gIda2DPtW45WbiiUtl531UybSyjvoZl+VCOaAUoKUvqI1PgMnq
EF6o2jYl/kp0Zaa2yaa1t71gNUS15AxMRP9y9KIlfW6haJ6kx2/5NPOdzuE6v4k7ApWmfwBbiS77
7lm20fTUO9pLF/UY1YF1nhan0WTPFtCYkz0Q1o/3hF9bfZHquk6Xyo3YWQ12vLPz/h2aFwVKSIX8
Y8csNsoeUsp4JW4kfXz3alcx+4sNmdciYHz/pIjRVyXMU7g0QBxTurLa+4HmHQM5rOfpkuBChsls
HsV8CWheIwHickCd3KTunsyRdGOXvOunR7e7qKqGwZMLIp/gdQkBlbNpt36n/Bdc/MMZWMfbf8Bo
lK3a0Li2kI2wGh1n0SxRHJufVojSaHXDsJg4AUeV/pUQrb2xTDmqbHsEsGSy62FZlCLZoUoQHX//
6bOH1KJErweZ8ATN+xKdZfxK3xvuLmYbVIpoHeTKMKN4KxLZPFwM8azElsqrH56djTZndFHelUQh
T7iCs+4UuDv9kgthxL/eCoRIBAAn6izCZOf5eTuYS/7bkO85lDraFBmLP5EjlW3k2WKgtbIrWfHi
GNbdQifCP6h7c5/nIcmqbXuYwjps87B/pHgmb689kSmexsuaaxmT0eO7lwV3+XkhUqlUumwnkxbl
ya215bTlfmc0a956lj4lj+Sm2Yz8P9t8eqbIRFndd9miUype8PjAmGovWAeN1v9y0WfMCSIj+3t9
G2Z26QQHqdLS+R5p1D5ywAtdrZ1fVEBmYWwZFYuKbY0rjFb74lGkrVHPorMF5MCfHWpnPZbue5dF
KtIpB5tK2RBkqwakpM6h3Y/5rIlkE4kVkZ4SchMaJO/iQqfw1etflfH7hkmnPbxssZPPrU9X4wlE
UP1wFjaK14pv+2GUt4z7lVKetsmRZdQ/UIVU0CPfgsQuZ+YPHzLfGvuVpavDDF33ntOJH+jVZ24C
ef/qQpGI/Uoethx27h2W3Wdaq2xMczHJS41VPshkRcKe7R/ivibRackiDIVdsQ+sm9GxG4HVTtLI
lO+zL6Hmif+WElJW1ONMQemnFQUabQKdMHP2Xn4nX1nhEzUe3O/3Qw3m85AqPDhzPEXVwqm0zk8M
en2laxQqL6dMhwY8DHXsGgQEoh5mFLZ38d0x414kGKWC7yGAsVemQc4/GZWQZ8qYJSUkTINx9rV+
gxKO+a3ZXfcZMEB8qJVawrjucxGSkHOSM0rRVW1ChqizspQHOe4DAXs3NmCcyKHUdjEK8qXQPrt8
9iytQzkwEE3A2pRZIOwkb8Yfke0x6QNtmWUyPFBTkgyhuGNcOgm/6f21ZTwkTK7OSu3XqaELk8Ix
uzbKqL0EI448XlpYbElBFo0IXJzj2tI0aUi0c8AxYVScEF90kW9xOk92AHK9DfU+deJKpJ1Rptw6
6qw3N0ZTzGL1TGhVeCJxt1rhTPnp4wFevKEXTHVC7QgRLTOI+ynVShiTDcHClMKz3nWv5VS0Fwtc
2BCbO39ZObpc1XjjDRXwBjYd1Rm0Ytm7t+dv3MGqQcZJe8D6Ksr7wtfYJmd0MbyjLJvUrj1HQChn
8s6ak01GSwq25kQbc/2Bv5Qg0mW9Q2TMpfUx90zpAgCizmFf7KP9MD466UPh495cTwaKwDiQdStJ
0wqoI4EAsAx+j7a9Dkwpu41cT0eDEqEXyvppy7OSEJBvz8rbzARHAZ9+ZX0D60rRlo230GCRCU4t
kGl5B5uGURk9sKkLMSCzqsXQazfZGoV1XkfdeRMLMx1P/J9ySDGLZtW5fNjYJzFrth7LtwrQdeAD
xVczAOxxZtWh05qEVJDPaf2TsF5/5pecTNp1xb0N9dBL3XUY5LHikhlqN/T6ambR+YKYxG3ZXqJh
Q4AJjWIgTKIpZUbhQrKv8eBz7J98dfIDsVNxeG7OD0r5ivCF7MZbiDoe+UB9tUATNasD5WM1HqWP
Zg0v2pNsdkMitOrEUTvgoBt/jhBM4udvi2159kXG1wBJraeQlk0Y3HdwCK238cb7fb+lC1QQyHe4
2NGrVZHVeGB6oZk2skSjlF4SAANzGnb2WM8l8DjXbTivUW7U6KxpjXTjjV114ESMoYTDLV2DhhUe
ZrFDDRo5jd098k6xNqCeywhlBJYvbatOQ/RexOpAXG0JDP6goIQfa4fAvKle+8q9JECs/trkRSgL
YdspzVzxHdIJLtmGpWpwV9khcagO3KNco8st2xFGn+uvmC4ED+OKyQT0aZFksEu9Kuh/ZUj3FcDZ
TV+RU0EcuYXH2ZEAtPRwilcn6A0NMIYK8VRutA9FCupwD1J55RmTf474hsNSGzRdmpX58BSI/j5G
XYlHcsJHFYQgneJAqGQTL7MF9HaILBa7mRRuv5exORljCwdDGL6e/djcFsvoZpdUPZfVeercg3FT
GFbRSBI61va4zfmV+fWmTSqQINuuTAHu7tyAs73FkpWo7jDpVu6B25T5potfMOkNW7T3l91Mut7y
q3sFlOaUXW+IEugQB1Masv4s3bR24AtKTdpHDtWrFDNv87m1MDvzlA5e8JCJAAD3D5wP2VAChGcV
qJDoG3DjLVOJ/hygAA3AEYMchecCG4p5i8669CaLHena61PurLn1PAG91pxCrFLBmHt6oVemb4XY
XMVNKcj4+6NvB9Yj8TZLSCGzFJU/sRN5gpA3EQstmOy7uhMY0Dh37xNfUAT/9cp3sYudeACKzp3d
N2SqWMxi4ooD4BSqduyiOW9jvjz3KnVn4f66HirNDI989sjJYSbjn4BC/Zn3FYRVvM12Pn9fcFa8
dLLk2D3scj73t2lIfb1EAInGC90WU2VdyJ2xH3rv9DSqQTT3vet0+sKjxaJbIrkb8VajSTk3R+XF
x80oEdkHrY8jCypyIgFhhbzXyucvrbs5BSKaoW5RAIt2fQep0rKjtyWUj46p+JR3Ks1ahU1EHxqA
sr35xXDkTalw6wCEBRUWlHkLxiQGuuRCHRkKcsk7VvmivnSk5QWHwQM4NXX24n6Q4ld+Y4LighEF
mnMx1jawWJNVN2siugoNOTTMdsmSZvu2sNNLPmUHDVcSYMq7ZhTnk0lr78+r1MO1RmsrEZ7b5a7U
fwn6DEebgWShGd9oPRacKAM1Ni2JymQU/8Wgha+CrCgk2fFmUoheE8wvPRvee4Tp7WR1VMCqQ2I9
OgQKznEwXbv/9tSblRW1ac1JnYluYbQnsY3J7O91yBFyaWEirnVhu+hyZvaLHnWqANYNT7Sswgvn
ogwpfC4RshI1pXjLCO7FbKvbVpJx0SLip7ncFpQPSY7bM2cMN78X32EybJJZNMMFYFBGZTT8guw9
r/QE49+eZrB/x7a4D9JC2/EOg9/y8u1AryzCewr6llo8kXPzUJrgGdaDSJHjo72k3XP7UYGifnu8
aZn23zrfVBN5663jJmx1rNLO8/3LYEpT5vvCpJhE1ENFx4Z3wtotB59Sp6sRQDJJfkd9J15tiKIl
ScQ90Zi4+ExhqSEuQaVsEQ1lVyhEb/Gfu4q1t45TPexBTp9hVrzAJ5cX82z8rGlOY8PSGXxWIdMN
uDRelyU1g+FP5FlMlT5uMT0F/v8wN/hVHP56DoaDtXZmULOhfuvyGpJzeLVbC5/192A0F7TSwz1q
CaXlVIblgTv41VDM6nRZsgBoZyOBJwGxxcGa/CakeG0exshmgvR/rOe3DankQPhzwZu8G3scaJV+
+JwFk962Ll0qln3Yq6SjadjrpKwyZ0RnPpmv62njMRFp3JKJN2G0n3ar9QD3OWcr8/OPt8YQAkYx
XpAVB0wgtamsUI3oL/vNWBpDCuERuquu0/KZCIal7b42SPFvSJjE/0qdW3tMzHvhvpCPtySjz4Eu
6xOeVp4t4UHkB+FJi+FQ+tWN9QgrCVVTaiQ5fn7/4xdkyLlTLyMOdYpB2YjCC2hLD5SKR0992U5y
3g3+DO8EyjWX051CoFIn0JGoqB/m1Ta/HFK7Qgxu7foeaO4qxxvQ47EtCmZniAIiOg1+G1OCDHLq
wzEcTCjlZ0yrxroaYYWqbGruSFcSZTM6MA7iNuJlUkJHZPHJILOyJVNKUoE/F1RSQcE88a3IUX1p
1O3a4owevjQIXXCPYKU/7jCJkFhwokP29vEwHakjHL9nFxYsB8xOEjHqHIBmQErw3Bb+TOHgtTuP
dlNmcRxWvYTX5rYocEi+p4qenIfTFNP5joTwwqMX5Yu59qbqMSV2HG4yqfTOW8WGcyhWDOY4lmaR
CO2gaITj2KuOm9tEGxIaGBByuszrTgCgDikTtTfDpizfhrqujQrrZ3zzdUB2QZLu9nHdH52sKI/f
haAnxp1aIUdf39upmbNJxoqk3i6FERi5lwHN71NZwsTBLsoqVDnMK9W2iK0PAuqKWsrewxcaEKGe
DoQu9GShbKCd6YVPK91nMADF2OWCrl0OAWO25qOW/it/UwJMVHPZZRFIYSPXGJP3TgWdnmVhEkCp
2TzZ40WQmS+jeUx4yiPKulhFxtstY/He4F3f3lKZUfuLKE1K2NdF7F4FP5B5HiJMhNOLwxTCu+29
2lgqP1zyrkK6jHQbDQsemDoDhJcr+rN/QQNHfd2wicKxgoEYFyHTAKCTNskNnP7N2/I2WVZ1NHjq
MIgCbXJeC8nSA5b0xVvG8eN0Z/4IssLQmx4aauwI1mg6C2DiF1HUuMDAX3NKBtLcKIFSDOOwqEKy
g114Z9kH+eAxkUKhV2UxGeVh/ts1iiLSKQKdqW751wZX03vqDEUnwHj5ALUtgBS+lh39A/qP+qZS
PunyUJJBxHQ3TwfOcpEKSwgZXi+eCb4IDRE81ABAgjFKbxnKgcyMI0lyrzvZ8+NvM1zKQO+mPl6w
3b61dKrypPz9cF3TzTS1j+wmgwAxlzKfbMiv3MxzUGNQdONhMwqM+c/nZf0kwTCAL000JzJN5E5g
qGnX+tdLazspmhArzZmiSSnZGcVvK7ZHLdRpVPDETfZ3CdGKT7wSU2qCD25TkgJYhtrZYp0GO2Kg
c5KMPnVzVtu6KzR8C8x0wJhg6PgKkwJD9r7ptf2Ccr9ybpC8C90t/KC9a9Dd1Gvukn2uc5AI2QK5
8yjsMh6iCW/6srJmFHNqLfDHOQoS2EpjiaHzFSqSBNIn/fchUcJWqeuP68gHSYp2nmglwB+UAhaZ
Td2Z2if5XtZ0/CUM245IfKwoobrlFHj8geliKVv/3/lE2plSec2v+zQBJ8rjorrSBQaDQ8T7VWiP
jugjlH0XhMopAx4t3HeKBd2fiGRwj1x/LRwT3KW9+clHdobt+RvDrUIreo0ktO3uXUJjc0b/Z5eq
HvqAQAk8NDdavDVCsY29RQseOL5Iv1guna6hirUvy56WFqblopatJMUjxk5nwmN4jktERDHkjcGU
vRyz2pUOR191GPSiHrE7a3mmWto42KlmRbAa00gBZR2lY7XUTyqEv04fUMfenXE92GosFl5PngyB
cE+fraHeAq7ssixxNhm/NFlRZ6sGy2d8OR4aEHKbr+MuvtGqP46CvCg2tcB9P/ixoMQwLG8F8uU2
W2+wov6OZgPnLqELImzv+hj9kng/tk6aogbW4eduZb7VzvIzo6OUskYOTcaRHHxMNeO7IfKuLd/d
YV++VCkk28KT637yPYD4MSon2jfJCIXUCGEnibG7utcpLavFswiTKVLN+zz9ob6F0UYoBskEKrzr
VbCSnCLcdNvwyJJPlDzDY6NeDi2gf9UQSXL2A5vMsJa7nW7WFB1tMsW2GBbamC+5XItwJOhfuek0
D7liJiTnZ6syo22MX2V2wADG1orIw2Wa9nwVRDoieM+wJxU+TuUAh0s1BhcNaTFNTMWHJKnHOae6
3DTsaTyCd1SIJpdkF61QnKA5/vuH5s7TrCx7YfYkjJx+XhnTLywFhhauxa6V8Xun9rJh0GuWxsbX
7UBYJ6832UswEL25ymqpB9GiLfKCrWwawU0pZvfGmLPVpKxQorRxAu7HhrsAaniSdgfwSF0X1rB6
eK2ZtorF/FR+avfw5Ddd9QIlfZ0et6gA7D7K1NgMHNxvFD3h0XAW6gb/xcMFICB4yUooutDn4CJl
JO9u7Sxzt3tI0/Anz9ag7z4ibPVoJFOyALZ8T9CWdll1DX+PjrpcV7Z4i9gX36gosm7ViBXAJGAH
YO0RSVxPYYpW+6SG73T3g0pZW0YinyOtG5lgq7xs8NaQPMgDFQ1e23l2+kjeVPfOLxCITkcvdIzr
/ygzMgvddf9kqIkJiBWwwj7nvg367rE7N8MjNnIc3oLKYeDqCRCT9ELgFM5uny+EVL5ToMM0bQJ9
Lb6vPkH34m3lrR97QExKzCnbcJZ6vP1TJ0o6ZOZbyWX0ANLegwH516PUlCL9FcRxP5yGphoddkJt
P/ybc4aLVhtCn+jD8I3b2tzX47HVfDCJE3hVtKbbEeDV5UTcS9qQLznJHTH+CHBU+d0mL7UKbUYc
ku1+fUdkmztW5luIly454C2Fzfy7PX5pn0CDcsTroDnEAM8SqxmQg4OzqAbnw2ApD50wrtpVu964
RwEYg/zLOlP/TniK4u2A0XONf1WH/UWqOVoJZqopkifpb7Rat6PoUy3digibde9gdKbeuBq00ega
3Rze2XBQ21XXCTGrIM3ankWem9w45arrM8wzSYMDcciUA3m5zqDVVw0AtndcyBzBupTyQ0fFLt0+
YUo4WlNbGCA2k9kRmwSxMEnlBlV7HdrWvwJUTl2RDPc6aaZvzHv0lrd82zjCo8JBVkqHzkyKD7sd
/bu2EaEMGkLNeqkpWQrifIbMnatV43KSRf0aIJ20ll1694cKUzusVP4YjvBZ7NyJAlAA4MDI2oaa
rvbtL9IvYfaR49DeX23eJZSxChXMKwktBC6HPVgoJnRNU2RK1pSiZLlf7N4j6vMk5co5vBBBla1W
9UKYb8rzaoNJnPCNsT1Mxi2OFMl+sI1zTuAuMchWImBSxij2GwiClQoDqtGYyjlbUk+sCwfCYDnO
p5BQVnIHWg/SCQP1GATf4ImofegabwACS7apG3uWVNPR8AbYhELITsfor9m6R0iqA8Dnoo/eEwNf
Z6EAL161ds6D1kQt5Paf5xCczV+3J7pGVkiPzufZ2DJAKFVwlzj3S3HAg8tdWeoCbRdqxQjdGnr4
vDd1C5MnY8BG0sh3XNbUHB8usXZG9/0B/dP3e4NrWp0QuNlLdC6n0696smKAb2X68PkAYGzUNAbp
25Hg6i3LaeQdSV+axmrWOAlRiTCrjQJevW5ZS5bQ1/X6vPeUk3XQQj5ROI3x85YGCLU1uu5xQ4q7
+LX2Gx+2ddrgv9SM1hRFwM/2JYYgplRNcjkeSt7Yd6qkBRWYAWIbyE3MMm5p6Ppz2I4KIFKDNImn
+myVV0okBn4fOL0M14tlWYg6r0GqUlp9Mv3Djtwi+YF6/C/uolc7mwzBGC+DTmfQsLQ4b8JMELvB
bXdqL42CIYmpFQg4/XdA4m3P5I8VtTPbfCVj+7uVJtc2RYG1VnZoGJzLtxEYh8bGSFQ2sXR2+QtZ
LIJSl0Pt4aZ2h6H8HYGHes1opJ8/VbUCIQSN9SwAcBVnHZIiYGN5VnqPGX9JeReK/NU8szHtl3vv
DJtR3bc3MWWTgnImVCMW0kr3VQ338r/AZEROxuCIDG8Hobr0+CQ4R9c9h6KeLTqkMyShvtRHJn8y
bgBV4eWGdNMuG9RBxKhzuOq6+yZ/KMClV7aa5zIZBDxcryzFN3FwfQ8yOHkZI9AiQytopHeI1Egp
lRowFAk/WVs2hb4uDO2LK51K5ufcNhDE/M24vZQcayIvISOSXQcBs8J1oyMmsYPgo0hdJzeM/MEg
PSYqFKsTj4uIs89WJliKLEWABVbPhQQnO3Uda2C+Pq09d1+gLw+LJdly3v31VyKLC+iK8MtbkHhR
feDUWQ52DokCYK7tqf+9r2+LUoGjQ33TSpp3T9gbU3rGithaPbMdHv82NjyOK5mYYpO6xTMqCD/3
NngXMVM3Bhvj3bWZFILGdRWDo8MWPT+VSDW1jhzCT0nhOJoed1GYZm7oARLi80iHu7ZpX3I9gM1X
E5iGtIG0gRz315Dlo2dCad7J5SCKkl9R198R2zzjHJgX/7odWHBUd8HLRBxaBPYBgdS7TnszDTKN
mRyfJ3RcTQvD7Tb3NQaacs0o/R6rW86Pc0QIHQ++pAYmRRfYzE35/Fb2HEGlTG4P8ZUO+HWeMPdL
5qVVtISITLj3xwIE1StAxxHxoldaDWtu2EZpLsEb12sbfwHteu5ReI5lzrJnRJU+A2utVaFZ724j
PkrcTQ5llrl0LNN9ZMRYRY8rob/pPwr1J/pipZxkgweg1TtUAgDUJwiXowp+kYjDcZM/FAkzWYzp
I8CPMwjO1I3SwBo06KGMhlpkZjhM+yODlj3AV/xLt9cPQtaBsBHalQXtwQt+sumZojPqkNZnOeje
TOrd/pT3tqg8QeO0b653Mucm3RE33mqUyW/UXI4BAvMIWrZtvhXV8VIcrvpUcvQRLd5EjpJoUnld
ITTxoEMCSX41Z4UCtyKEdA05YWGdo/QM1EkDHjkKnFp+z5Btr4TtWVOqIBi3aJkIbFZOKwEtsofC
FE37c78rCYxNgaZzhPh0bGygVyJjanv4OxCZL1lg9C5I09cJQQ40UWrD4vjVmKBoUX8oOCfg1fe7
EKrTAixYKHh6NmcsypQ5xiflVU+JXW2wCpytJ0YvxRKF1Rl0hqY8bYvcMJSa3WSzzU6U9nZWj5C2
BybAcBa9cSQF7pHM4VWmv3XTLYoHefr9OveCQDiRYl18O8ew0fRrgaSMPNqB+O8jv2gTDfkbUIJq
oi4UeTvk+Xq3pCs7Vl/n3AYGVE5ABYb2vm/4X+5BEmO57WfrpAwpwde6WNFGoQBHnVHBTL1VuNqj
ieZmdhepdat5IBP9NM4RptT2Wc/8E4HOM8XyB+JNKxt556ele0uKV+kqe0x14YOYk643S6krMVJG
awe1Ec+/yP+ynVeDjggBBzzqDFdPIhmxnEwcCntFFRsQW8ERS3TkmyJm96NWeOxbQ7FpomwDegGl
sjxIWTUVqOa2uOFF45lbTp+fEf1vzCLFuFHk2GXB0u7AFDxZXS+MLUNJV4fJcpu1rXIDefgKBY4F
ZAt5wvZxtUXaMSo3D+s7Azi/3uz74vBIdVysojYfEET0f347MzLo6rwP9BCuaqKL2arCO5c4JyWs
jVN8HiYteN+2t7SfnztgU3SGRIxBYPrP5apO+cCnoEb7Os/GmZ6NfKVuuTogOgVuAflIDXtCGWva
rluPIdHXjG+lPl+dDoGqeOh++ccknlPeSIrKvHA+i4HouMhsBTxpjTd3cr2xJd3GLta77cGlhaMz
Cs1TLeZASdgb5vkrG5SINfny9HTtJLfkrR780SXHbzVjQKmx+Z2P1aDRfF7E18H0z/xTMdqRfnON
HmR+9Ihls7I5j2TbMY2ZwU3gXigNcM7AtVsCVDyp/qs1Ch8OxqtyAm2/v+7ZmZ6BqLyZalp0TjED
WorG2e65qpMdVb/kYQNr1ebtSQ+G5jQaMLYFPsQDplmFIcWYEFGRCcYR270j6yTfyvS/hOnloCjT
GWJOblfZ+IfqmfC0zbU8EtqdftYx28NVzvpSctrbq62BYnaQhvTNP16dQpOeAXobWpGPd8W+OS7m
QdkuxVTuQalJKev+XxkEFTtmhHKR6VmKZPOOLCYMa+trDnlWrObIPa0oT1PAazRjxVeyv/4PPb6S
sB6+SSz9OImbb73bkf5UEK37iiGKB1VOtzKuB+D11YwSSoqDsFbirHCGB2uW3Dv1t/WpCQ5WDmX7
ZX5fURNE+im9gF5rAWSu4wJzljJrPdU6JzoxY8vJumJF9psf/nX1HVALP4M2DRYwNmrvfDP+wOKX
4OF7bBZAvpQNku27H13e1pBbT8boXPc7K2C689yu89Gem+yvdWrSX/cN1nt1EgVPB4nsG9oQKHIw
ft1SkdgYB44YibmRaDwzZKPv1qC+BrluuuTN80BDSZW4Q6cF4Hk6LHhB3Vj/XwKNOaKIZiINfQs2
zoC6PenBCgAS9EVVziXWGpOBa1Ut0ZuyyVlplbmmTu/FKFAZVMKlSaUnj55RScG2DEmHSVGuQ1Di
+EYkwWNcozJqjR7AZHUANPcqMVeR1TZ1dTTtsnIfXiHv+ImPpkjeVvlAUF1+kgVyLrrgtddzpwa4
QoO2t0Iyl5uweX5yrRu+Kut+MYpRXazYyaDYO3BQ79SUdTtjpqnh1qoUNounaRrxyNOCqRELjlHQ
hZaRWTFQh9vQlqibpyisaUHVGrz5npVW+YnL9iurJjz+wbTO5AqqWl4TpJpBmtks/3V2E4atkzdr
ts/yBRKoeu6vYCxrg1EzP26h8+LI2LYKOrtBhGsR94Q5IIiBaQ+4I1yHQi7a8yGPzLDzpJ5TKINc
1f6MBidR6QYxQNaN0TuS3vV+MVpk+Xohc23t+RNYOge5dss/4ZsKVyDhlnC/JKuGlh8UzS/JmqOU
NF5T6tRIyQ5XKzkRxAbMIzvG9Xm8hioFDBLL9I0cF20LEJiiudMIk+nndnvgqKpqvSA52EHsHrKx
7PF8gb7p08KKodlpNmykRTXl/g8AJRPgiZQ4CxuyZgGeK43jhYdKXz0Ah7YcIrwbb668gZD30Fbi
hgJZGisT1TsIdT7fJj4NLcRc8Iuf0E50koO7JZbcLP6f4c8Go/eBIBZId4RMJL69BiJAj4mUw+fo
525ElgscqKw2fUpQaLxmA6NTs2naNviYpFxm+7qrlDD6YfLVgxXY8vq68W33aKMGlcEdvP1PD2e4
dD+AJvfNBuh/8yxgioUKd5lPUetVP2VjY+hJQCKQodIo3DLCl5EWmMEC7BLrmITwcUm+IvB0HxPy
V8IvIKVOipraULy4Xw7OmOnOGeiKGGArGOO8rFdBB4BiqeWlO8XfRl5cc61XxUdp5nbBr1S7lRmR
iJgPSJOfYdg9sIapr/LRHAtmUUWFEx7VdBr8JLl6XssIDK+NJbYFHESC1YrpYGM/KH4oY7TKOZwk
EmUp1rRxRGiLyevAM/9RJ5AeIOIvw5Tb6p8zfVkywI2VqCzh6+0dQvWXcl2xTJj0+iP45eFhWVo3
mnUsIQX70O9O6EhXwDvebKUXCzo2fAhZn734AYwgt9ShOtzPEMVMtynR6C+I59nwJN9zx/QLfHpg
13g5yn9BmkiP8kEdHyj1jg8BPhceCxY0xUuVgPr7X8aYPdfNLhKHAbCZG/MTw2pRhVaqnpmj/iPj
5gfaqCN8Zug5U2f4u0OSp2muKpNDvUDUiik8p7qNQvdkKykzBAtRSbSVSsWjOqqPv8DbTLUKYzf6
tLyJtiAy6ETCOdc5jz7cfBtJ/zujB2tlpbaPsrB/E6/bGuyWts1lvEF+yq4v6JKb5CDJDEGUAXNV
xUV8crLRmJdqSN01D/Iaxa+HVh9e/FqepKvIKbhKfOg2UPzlIrGzU/cxG4vvRDqtx57VmECo7SSV
QArYeyJDHIj3d2bH0rZcgsxgXdw9ohxGVVLTCBbXMAN8iz6aDvrB3FU76+Dtltoavam9hVSBD0zd
VNuwRTyfQd0Ln5GdAuoyYMtzjwvJtRJDvGMguh65IUuOOKmsUYPvhYz/gKXIfnwOd4d33fJivmRC
DILjLColl/htLdzSCaaI3od4WJL2LkHK3yyKGDqKNKg3U9Z1/oxJRX/7YKfOFK7L3P9Qn/Rq2ve8
xvF+GGZBRW00V8A9FkqLLTD8JMdwLLA3cvqjmdBVyIOHWoMorX7AQa2Da8khZQGJR1vinYQj75i0
Vr2TAn0OQo2G6lnQi9jbXiDL3cjiIapRqn/VOdvjUQkf56tk+fDdvAqm8NmQLmJKimaUfvcNgVdf
JVTQpwN8awBHQ8Ye4I6HDuvFX+Y/WUj+c2phu17HAGRQaXyAdFxjOM/Y7ADmvX5UlU8kJm49GzRu
+ri4y+eY88oyMPwinNrhakNSZeeTyBPadSPJgDqCxmgchgQW3dcBcsDmXlfuTxDkVn166umnDcrq
uT8zqXLjSurXMyXHWE7BetP/6jbb5NJWPNuon0H1VXn5USCMn9Nz1730U4f8DB4dbL/3L55G+ue5
FSWgd6GyOI/I2t1EoNC2cmR9fmgbxMs2Nl+YBirTHf2daBLQ9bA82kRr9DiJGdxk6gJFkxRpliP1
DXD5IRQfejvrxH5WlG1kRt95qa24v7HwetG6Ovm2bl2bv1j9T+mbWIl2GbLQrTTImKurs0KIx22X
keXGpX0P7/IShgs1nUZJ5htGHHW65XhzZ63lEOCCMhT5qKigZl4YwoezTWgxJwpNGh+ZbFDqYw2Z
B1J4wIynCsO+J0nXhpcij+vNu5y+kuVM3KntxElRnBjZCSV0uTsd5cc37TZBOJUE/f2PfivnLIrQ
XnOQ157omn2WcD8XscD2I954cjcWMbRGb4YmPP4S/vKCPu5BeZpVIYAvvWnZJ5jCyUHAJUdQ+dAj
qGVZ+wMwhPnmCHXyM66zX7wxpV9vV+UPykRERMT8KS5R5BYdULdN7bQki7s0T1+To35lsXBeasQN
E5/+OcpWJ4pjZhqx7H3OBRlfsfycN/pRHgXVXMgPnj7NGLhmKDHhVpI00ACICYk9M68RPctnFOYl
YAENaXr2JFIITz/IsynW7CWkZZZGSY+gCJSGRy4Mf6qfAuYTYJR2Aa6iBjsV/x05qgeky1niZkuE
FunQslLGYybFIqygYDum1SIFmB3Fjwj0Tvsvwve/NK6hV99ZdsdED73CMIwwyjUyZkrcuv7eCvAQ
+lplVYxQipWkeSH3gkW/4V5FZOB5uc3cPdf32yUdhaUmIydIJUMEyqoNtrxRxFkgDHAnsFJfqsvk
Rl9n3tI+AL19F/WmeEsoTwV8qVIxF8osH8AAOSapYS356QKHzHVBsdaiW3wU4oMh4EXDM6k+IrUz
CSyHJTiJtnGEJJX2sGpaQKxDSQX31Wn8+WEQvTM/WvAhq5Dd++qFUZB0JQao413uCkoRklg76ZtK
I5Y6I30wGekpdgILRTb31yGVp0+l3WEruWj814JxoIP3qZeuuwXLVer4UebpB+TzP6YGuMPm+EK2
5ZzUW1D2da5DpQ/7AWp+dNDwrHdQECqXxeHHjJt6rUFz3fBZON9lwAbXERADhu+bcJllV+q4DzcN
jfZ5snI/sEom/rYh7Bbq6Tkiv1moFnn/N4Tg77CLIxhrYEIT/5flO0msaMF7EZ7BiTFxS25TTF3b
cjoJW8WSv6JDHxtEVTybA7+gUlNZDJrgIvDJV2te2DamRYE5R0gJWUyHof9Jc0X9oZ9TzCKJTwqi
xYJ0zRsu39Z0hK5E1XRti21z0kRkp3HhY3f2hq3PO1xaLhjfgM/JGZF7/WIGodVKgxI625324xMY
7f2m7w1/afSrhtEy2OWN2+HSfxPYvOtO+LqQAROpCLAlpB8RkNpZyncEaz4D5qb9rj4YPIZ+6W4U
jKz0kHLh7j+UbG9+BDVGawPARIgdoHSANBbavZc7s5gtmyDuM3xqXq9+8199ytpdPYHWEDs5xUWV
m33UXcO/pbe+p3ZjY2ZbzzIp+mkasEYeViK7uyX5Cu57EOXE789661Xf0NkOSSGB2YSuA6GpNg8V
N9Cff6c+1B0jlPeUwUOdYc3XkF7gtoiRKCLrwYg+2f082F+i1QvMC8kokaOuyOphwjBbwtVn4c5d
b6tVVw2sMJKpV0nNs4JHHr/F4mUu28j3AnT1rEmxCs4nviAL3tX5TNzzSyPFNTR/p7Qx8T9ckhb9
c1D4FKzn5BOR08K0hmPgDmgjpgoG5PVKoZe2GXNKVsOAKqsyG34TK4yrLcPxzoq7WPC4lLOP+DAL
wvlOQp+UKcTViQDBP2Izcd4AKStSRog65rP5TYeTE+vQcmPzkMpa80grH8s8YU6NxQIQwq7vwXCu
nkVFtSGOKBQViVpnVnHnrZVVbLbLBb5F72HFum2h69X0sDqJ5YFG2mezUcH/w5QWiQX0K0v4nF1D
8mYcpCnpBNKuGTqHK74TW8+Jz/8WeL/cmZ30GwV06i6p0S2kCjIGZYa6FqWSWx+4ECgUE8dDwy1a
jmpDaGLFjeDtbYHH/sV4pwGB31ngw5gIK2UQJf4aNx85EZtCk1plpRX7U3v6ih6t5+oaX5Y7zuBg
jBorYtVybzPqfPBwfotZHqWScBihMSPzTSJCP3FLN/uZrNyxwjGsItdstAHys8mziHbvZDcNm6sN
FcY3Csi9OEYUM6GvPS2zCDWrrJbqI77hQ0XT6H1dc5SxeRIg+bZDc/1JA9XaIUT/JLgCT9f69Cgk
MTm0NTIHTg6sHtSx8m+VaVk5s/xUvznarPkAb4KjnWT0V3HI2usYYIX77+SAn4PKm3Z2p/oRnKC4
BDYbBtvzfkGwzgmRKvV+ozBf+abHI//qsxYIEVV70ov6Dld0SVYlobEBpANq+DSKnl/057dQiWd8
mrC/AWWpQtG/Its8MdlQKdscITANeNLlgCjKzsQXyJtrQaiJQUJHD+swUeIxpygLCfveDr93Nzr0
Yo3eRsEF+gTKZz7pG4oRcXxMApgUQf0vONSSBdMHSz0Nhgbx2/RJDOUk0qUweCCNLDTQorGvqsg8
XUbc7fge9X+zYgS0nxIoNkfjnLjDAhLgYhgjKqxQB+4x8ZRTIApWdiHw1hY63R7IRE19jNb2AapA
ebTeSPQ492mM7EX3+/jdykzpeK812sTOhLpuzgA+4hQ+wx6JC4FSZ/+6dn7GExUgnctnUyEAL+KM
jW1CV2bI3yZBl4hR4wv3rK4jbbJiiBlRsXM0gTt9ZfLdqj5+YseFKlWREl5Fri+G+I7z9L15fy/m
ZvB1BBZIhng4U8jQRKYFLADJX5t9N2q/ksF7wrBeJJ1K0f6X4sWxGK3F6dhtn6yLeitMsjOvbfNY
Z7EfD5HOlP/kaJt0mCIyQNRIzTILLZvu60RmwgeHkMX+srs5+CUlLd3gRM6dWdU/TMM9toV9yikC
7uai15Ppo9YS1t/j1TZKUajb+t7W+lSnT1BzUnFH6mqrsEubbRC5wXP/hIclwQxalT4suhYBcUfo
IIHbZnvjr6aJafAHzmnnnrmLQnL7cfcdrUDXD003MMYCLHfPtSG5sGWEkEXGxI9MxwV1iR+3faWe
rRju9slg6yZ2o7tWX6a2b6csaJg/njRGfK9Y8up7JUuIxePLj7ycsaQvPWTq7gWS2w7fJB6EZdvN
0lVKtpksgetPW5jK3L261J4g0DS5OixHKDju4+aqUFZ8H8dFYuaNKojQtzZxpKbyI1c0aSq8dlP6
qzJJ0qBSdO1Nx9DYI2AehtTmTKSzRfuiNAEattwv+ERdSRivJ0cdfzhk8CjmXPOy7N4yTQLuMK/I
lzUMyNsJpLE/Ult0Ytvke/BL4TZ+P8cHvoCY0xj6MBMnvF3K7aST22DCNQGL480wg20m5j6pMqF4
sHLUb/IKZ+NmTY2BqS6oHt3vQPdLbhWomKcO6WLZpPxil4dT51UkrzkY194kw0n12U5q3TeivMr0
NZILqVLMpvSKyk2jUYLcrAHBXTW2u2Fnror9NEG3fn6J10sHjuVGdZJOA+e/8yad0lFItEw57f0e
PeqNEBRzM3WBpiaJWqf6Wjf9U1+H4BhGbhUEp3PWulFUEwPzz6pp8WW9fRtI24wotfpr4oaJx5zb
IZk6Puh9D3rW/DHHLFCUrVIdRgWZr+R2Dc207D1RFKYtEEo4FUyL0x70Fv3DQyq6UFsYtN31TcWA
8lTne2drhFt1HlOMAfdF/JLXFHsr28gPPIf9L/ErWnYGKy9BDAW10eniyF3GybneohtZVC7riBrZ
iZ+tyvydVImGaOECtI4uqLeDvlfRSQSQytLBFmd/AQWGLTxqLBvt7xUzVBlxjU2StrHILCDYbaNR
e9HN8//jGui5wmlRVjgiQaovGvfyOKeBy6qBeRAZF1TEazWoKSn9vkPbM+TIFtR+zO6gy9vjbvHc
RYnSEN9yh+STEiHCwSNEFqpKoStmaNmGSOX/WyQJLXml+ArAvZiRHJReXDM8ZlJV2WKEJg3FgOA0
EWLlq63+19lrJY6zS9L3BK2mZ3DFhGVpOC75Uu8eilTEi3xjX3mYh+29B2M1JAx2Nf12XtqOxKJZ
YTZhcqLHp86k+QFx6sXnKr2F0YwBL43y44Gp9DCzHoXZ/3cVFE4/xwM78CZ6Q/6WTwKGiFfI+jpC
Vd84fHStKWECMwxPvTsX3k471LmB/dQzpD+hRrlZgBKKdEeUE4krEVmdNOq8gy8dbQw6RqYBq3fC
97kRfHgJvzWyGl1eLKOCBMGOshrUqFZFse0qmbkQcjp4NlR2NItiRrJFiMG5YoocVwURCi2RR3Mn
XClN9swCcOpysdtMsg7cW1pg2+9snfN31GZhf9GsMjIfbyt+2Z3PdKdoaAoEqV9wTQdSHE0u2R1s
Mt37sI3bmpHhPD2am8g8PGwQf1NPGFf5mx43aGSbG+yIRTYib3cCRSQ3ckvOaiPSxV3GJ3f06X8R
l6wXR1Etkusof4QhzGGyJX5UBOtJzdUU/FToPWMXm4/FJP8+U7xcfHzpvYGlyF0RE/sIeWCcaXZ6
pp4psDLWWXQgx+QhgN8l7AcBhYm2UiPxoGhN3X2mbvXSa+mYR1Wd90idePnUvmA/6krjsLnFBMdZ
XlgNoKQS61Nsg99qm/qzbJquMPrzq6pZy3Z9DNNY4nuPuePiNtBG7oPR8ra6knW68leTvumcHGAi
HqnVOQ8Q/IpWNXebar0WwHBfWpDA3+sfRN/XE+oLZC5PTEjrXUByd3K/jYEw/bWuOV3/VUT314p1
HTcf5Q6o5Q5SNTZLEJapvcrS0qdp8+4iRRSzegIuzcpKRe401WRmPaqm9+Tpab6nR7CeIn4AuQcv
cJ09ccFCj7AjpgWa82hCmfLHfNR5qWxiuwjs7si++J8eZJXcoSPoRg+GP6syGO60+k6JRKtsflJj
Y9rDJ1HeCbfot+G+8ygbOzIpzTj48yfuYoTiR0nJ5PNg7ykRYqL0w1166grBP9zG75fcgUNfXZeY
o7XPdYskg8Tlgd7BS5FVnZtBHqbT2UMqD1WZxTOx20Q3YxrCBhUZRtHcOkvvAueSST2+ZUa5g7MJ
ZHITuOcJmtQCZWIySk0z4amIHZ3Lz6+wkVelQdYW78yqj5dDt38EY3ifGdrTN5HNNWz2hDphBH1c
VtdWjW97Xqbt6FwMOVdUuEjOR6/EObBhE/NBHGGALkSfFrmYBmCaWBcWYKdOVs4mQzGmv0KmX1Hl
FWlBkZDTXOKtlo4JW765edVer4T34G3yIWrML7uCK1HHjrsJg5dgT4nFwpIPfGF+oSszDeWNUGeD
tFEU9gFOYK9YcXYexIqj2v4PbVQFYFwr8TJWbyTrlJPzWd0q7EW1jYqXZJcPZdP82a37poGK8SDr
PCoGnd4CfU4xx96RSpwC6vSI9wviprcrlm/U7IQa4itY/qPqe1n202bB9uJltk5PpWaEeqxJ+c4H
u7+ASlwc9beITIHafO08XvXyDqXRBUBuFWvQ/2CZWa04jXUFDNLYmbLTjzPlK6/RPImiQBbvLMFi
vkpfIVWXMEduFvIUZAshnTZz28rEg5y6nZ9XDAyGVuXf1Q2OIi3JTv7QiAlavxHLGbYSPoUEkMLp
6UEgkj0CzqVBo8uuHY4zbpmYu3fzTMbbRqdZGlJupccvmKe99znAk15kiwJhEabkjoqLBpYi7uUG
YcKseEWYc6lqCKbGs/e0zLNtX577nrUcJTaEOUjFG7fqsGl13R14Zi2Tl7K4pV0HgR0tMO43VssM
UF6W2gQs2oLeUmPxQcvlTPlACXL9yqqTEXPMVy90kER8YSvjNNlBaE2vmTWEYmy3I46bIhRfIbRO
+vaPgSXjLv+4VcvXEa0vNIBhm0QtrSJZJapDv2ZAbqrSdDbesv/kr5ehzTLqZWhfk2CuMtERcFxI
9KN2YZO7VwYcrfoHl6DgFlgfBQZd8s763+reEmaRM9dTvTTiGbJZd5gEXIKwgALiaKuQ7E7daKEP
StKo+l/T2Y8BgtdDmTQlVchscGWeNOevwxh8IFl9+6I8NOzEd1k5ATwBa0vD9eUvXgcyeCI0WVdZ
LeC+Z3UEXI+k2X7+PTu7wpJ1Ci+tEcjW8EW4ns/rjh7fJf8EXEtsnM7zTFaDQpyDN+diSXVQJpav
I5GIcTO/S51b1VcFAvo6iQJVjzWWZ4pje90GF4aTIFewgM+blf0QhkDcaM0caSfSfwOitjyUbIPu
uzXATkjIRzwTxjESaSnBwrfqWb6hZc9JbmDA7/Y7aLVlqGfsCcIzvOa66App8PokxJbaQjxlmd6E
yPg7S6DsLW04CFCze5+a4g2HzWosmPL1nFbeqCdN8mCbiTR8qpA6yM3FHyQeLjLew01zAVS68cpb
dtCzEsmL2zK83zvGU4iAxeDHuj7hdXRHIc8tfn0h7v0YgL6qPdfltkHy6ahWIDKMc1KTS1jcIKDn
oVv+ffU0gIQt6Z/yAhf2H3zQz116q707GiZ+jqwfTeTUaQSG0tVYsLOX6yUyCQatiJRzKkxBR8t6
0hOEsMdTVg3nB4GGnuHjXZb3c8QaSEqaw4Zn1iive7CCYu8hzJsLaAwgyl14W8qyyua+X28tbe8G
Zr63U49pZbLulcqvhm3Wn3FXDUk3D0WbYgWWwKtPamkfonsJiYlgrbe2TAJsjgb+YxwEsDpTXRj1
UUxmBTCDNGIe0xc1arfdc06S6SaWF/SGBK3sC1Z09xIBW/J0bGGISc44co3z1oVxZGsJaUQLoH5w
PMrdzjLYtIxrsiLaV9z3AIlxth/uCWggMzslpfGJDdBJLHcXDaxLBjAA8AdJMRCDBiKKZ//H0/Rc
IZct8eQepMa/GgCQdIGHRi9+XyHoRs27hA7p/BXHBMg67GGXBMSOfx/9bVvH7OCSGPpBFAdJkg1m
0pSH1pHZ3b7IIKG+t+apvpkDnVcZBI3r/uWLqxegC3c9d7K14T9FlE21WkQqaJ6HEvfScr8cFTCY
t/va0TsovMcbSSmiX1rsY0jhL/YAEgd4CDV23kkujwXw6ckArG59Gef58LJnIrXpMCtYtyCTL4Nv
/v19OMx76sUZjSy8vcoZb9W9/HCIVc4kQuz3Jsz8IhYsJNxZ5jatEIIns3CeXSryXLmDPfQmaJlo
n3y6X71ddje9cGIgKuB9sOpRdmD1/mmFJq0PwGDOcQFQED0x+MDF4g+qwopqEMSoBnVotnvQm0UY
QdcrcGPumrQVx5Krb8/L9h00H1bEhwc3JI6hy9Av6TNrB4qEB/pbs6aSe2/9hBLHpMr3KlPN3qcE
0yaUOHQi/YleIU2snao6zDvQHLLvjC2704E1KwQ8+gfDV4JaBpq/KKNq8ZHOPI7qhXxygTuKakYu
t/8v5dBxWxmwWDTbS9X5I23fC8+Vd7acso8iiviaRAdpkz3yc32gQ+xfEgIoQ4BRmHwO3DeLteAA
9XPKEF4XifSYbaluVaOVzXJ2CvU8g7ZUYuOZEiexLycMU3H3osZEHSpcAFtQ6EKwkBHFprxD9SfO
PsTqFUH/ETf+PXDLH05P/LJEuecJco3J4h1nx9hiQXDuJbdH9hoPKfYFzaGoX191hKZ0ZF6OEH3D
60DNFzjjbaKTS6gB9pEcD4Xh9PATQaieBYI3bnzJczJrmcH3n5RF3nr6pLp3WX3kpKCK9zh8Snfv
fSoRtBF3EeZi+VFRjEnJPb8/riKt3fJ6WL0C/5Bf3c5hw6Iq+3kzFFlWvrQqaXyirNi2JAJuNsgj
h5xG3q/G65Sao4nmdcileK/2mLfXs/SvMrEmNs20PAHHQRgPdf2XsVwmNG5P7gRjeEuf+dtUiEeS
O5QXyjZ517RuzDs/fitgGKFRP9DOU7TtCNBE01FHdMC4sN+OKttsQfTKRdxSlb61iU6C1Y0rdsAv
i4zYMdUUmzNRR/0zP9zBQfbDPmh7CRxeBWDib6pdP2j/H/SkY6EeqYGXoWuskmGg3Yz+f86CkNNl
21RaD3nQcppNGt2eg60IZunDSl0iiMU1w1XNu3Qyee4Ir1HW7reBexpTYzuJZAMbnVWNkHa3LWP2
TblsUmL28h1N8x95w6T+dPYr7UKJvGk/TNk6RylpyqZZF12LiqbyvKAM//8P7NjX6iJ7nWfjUmrM
OVx1/E1u+XeCwjjTe9TF12ykQJgzSHYqOTbwlU6kzjn1VXSseF16lRJTpy/JAr3M4iOgYID1Hlzd
DfQlVAuEAYdcVVA/RpBvKpaUR5xTnlp8xpWSs5ZLcfWOMcHIKxQpyCMz8NmKo4ePTT3cpqJ8Fo/O
U1FPdGO4hkiLuvSMVWHrHA/G4gISSshUcj0BQrs9Eas6YtEe6WYwJxz4A0r9cWT4q0WpWo6jqLuP
ZCEOjkz4MoQHOJYp5bEkqpbPf1Z3yji3AK4QRoCL/fxXAjriGinn+/edVE1RKVsH+ORa0A/usRFb
0csBuNmdxXVtKp+2RBvX2J9Eldaa7P6WRDnFdWQIwVskKUPr94WWLnrn8zn6Xq+5bY6WJ1fZ3SZz
osstZLnziBMFGEVRBM8/INCa6hq+6k+0laefap616kI1tH99ZfdDo58gbNqHqGv6BAf+1N0DbIiW
vrYWMiyk4kw90CYfjoGLAJlWBHLwWeoMFjKRTZrbCYGgfNcsVqUnRU8XLjFo+akOnCb2sDah1Dxr
WYhqk6MEtmmVif8NRgfkiUPZM6hZHjJct+4YdMTSvEOCAHQhFnK/woGq7zW4eDrfq1tFcUme6VCm
iDzo3xLskJkUp1Hwk040+VZhGNtKuAUz0LWhTOkuhy7WnsE66pZt3b0uytHwK5+MlkYOVjSmYN12
+iLacE4VK2CNyo6inni1Bu8kbJEkkzIKzhSwiow+URJFJ2A7KB0Yrz3nnR0d20d/gPIOuAFBU/Kd
fdBvfspfXATUaCf87uUxYuB9fRK7kKjf0NIhVMUGuEr0BBh4jwETz1UtEIWz+3SPklti+MG00h83
XlBtJPCiAUX2FuOWTzPAoAFRzmO4ubkiXqQDsUdO9O01AJjkHHSwD1pn/u1pmxsfYZc9GoxH1F3L
AtiC9UcXYXCxLgpbORkww1ATSDzmNLoiAl60lomOJa59ZGWph+y+Bu3eh2NHr2fx19OECrtUO9L6
bT2TvgH3DpUQviPNskyPOG1f59+cBeJBECnPuiZgSv8WqxwvwJEDgPWUzKzlpZJUoPQkSeFPTHdA
pY2lwNIzz6HYgkWCMacYRAFm2+TAvWCdQtO6Imi76X60C4pfbR2r/s3izy52mz7ug9HMOFKqDTiV
nbY14PjEUyGpUGJx3EUq1DRK145TlIM/wpqwTRzIOfLajof1L6QrT8ieQy6IspDeEOB4Nj+E/Ra6
lfQ1JjJ2BZs0wFSsI/xIQa1qEmvgwzer8RMztiLX2j3c357vrAaXYhr5EmrpWiVfcAKLk3iWE3JV
3FC6CD4k5P8fUH0cesUB/eR5XCocyHYVTEJjjqISPuAJkkrFE/sBqwy4NGmjsfCw1Btoscuj1i4F
bX3sbMLka0l0fZUDmcE4OXfzHC5FfQPhfEZvrYcq/WiijtPdPIqH2hldl9wtgLOHTn9JlHvOqt5w
rm5RD+oCeAWjj1CYtc7iPrAEycrT4XiLff0qjq6+bB01eBzXGM9gC/ogNdLsbowZed9jdFO4gbhq
/wzRKV6+luMCXhvp22y0SpcF4y7HmZ6omcv3eABjiX4DrxcVMm86tEOeJD6ojhLosPkW1nPq+U0l
XJrRYCRGEvizCrAQ5zVgPWM2InNm2rOjGXDPGuH60bIBS8Yw+4AfpVVbcPn53Psp6zI8VrYrZS6X
SOEVnJHSZ5p+zHN5QGDOkiV9dzwl7DnzbhVMuSpbyb9vCqM1G4YYUmtgzJTWOkgqGguJumGfeuga
/Za2WAgY/BkpCggDMBD4YooL7Lb7oojIoDKr7YGv/q7sjgNzHdn9twbbumuZMSYd6mgoP/A6XlMH
a5aggLmNiURvWLHdsPaYDtV+quBE/tKz305rBLAuJqH/+IUcqpcVKmJab73W6MKcP1SW9aCJR60u
TS5MGN0r7UuFWwJYbe0xc9IpV774tirxrww/+7/WevkyZiyz9Fq9RNjnZxmvAXEngN6tE41lW2tx
bleKjfUqGJh4hxa4UlFPSP1ADbVpeZl+LWlBg29GxFfRGNLXERVcvLt5PYxQ1vMg3agSlSrdi0F/
aEPJG898EaimMpMDTFviH/wgJysLuyi9FzmhXOQ3KyirUZ5WpemJhAUoPhQVcNfyN4DZKR4aV0mD
XIlu2cWFF/hfhziQR5ezhd0C/iN0CxXsrYcuQOLza2FhJ3EYvubueareyv2bZKDJIGd+ePHdXVfq
8GCuF4nGv5kZ0tmhVqzI07BWW2FzAKRB/FWQOTU1O4oUkS+HrkjHEA0EVA/JzhK5Q3qN7hJxz4WK
IEaviypYpkCUJ+3ly9lp32kMYeUzwpSDjOib9Osbv6XDWUtEpt+ecodHpx8gqvozz+2NJ7EK7BOQ
lUuGlMhKPLd96ZN4V4qsblF0cQUE223yXMmAGeLBWsTY+D1gjNjzCUTIEE/SG8Abs0UdGv0NAYUb
F2B6+3BUOJ6sMDHIHDfvgTfT1MhpAxlAW8KO+8ODy8EDYU1/2JRjGk1TCouKCwQZ+nPxscGJDmec
fX9Mk1S4AuRrEsgUSdcJBIjb0YpYKOHURDCwfaUo8wSx7w66SskAUevD2ekTkmf0xtaz/swOjygq
7MzKgp+lwejUKuYNC+b6ilO7btzHTMkF0vVrTE+mWzBynHtWbjXz1A0PATCtr26FkSO6BxTyZdct
6KqVYQ900FI5OWavkkSdSc3hM9AW0134/8Ff5jZc2wgOwGIAbahlJivT4zIfcAIZyy2giC2TxU8X
/oPbS+LMwz1CTlQTYEI/tSIB5yRJBATF7YbK0g7FfXq2O+/c982KNR9hRwdHk7KzG83+SzEb/f10
xUwsoN12oTvsT2iC2UtPaixM02qzl6REbNWko80sbDOyJOi1+Ipd2Kg1tqKYV0N2tukEBh/LXTgn
l7d16mdD4JQ75pW0BamMf3kI73DZg75u2X/dQFarMa+TQsfAQIFZhB/3gSNpevuQI8phQIxAuWFU
tFdKhg5p5ukTlSG8yywACkUKG4WVYjSS3sCyfyaU7fLevFd00j6xHsTeHiA9Ww/H98cwkt/pUjhf
hueq/X9Q09oLgdxvotHucwD9bTqLDcF1IEhJc9FLsC+v/nc9RW/RyzZncTR6tCAHEC3lHgkgxbAL
3iIxA+B1H+N9sgPiyC6BvXWd2Krb1+ZDzHc92ssE+pdu9HyjmvZ1zWw2s1q0ASY8cvw0Dq89p8ZV
xLD/cNIFOKY8d4bH3+804DEyNcb09uBF9pkSCosjPCvpESJJVrPGNE1H1nTCYPiHHzo5qQUjDvPf
j1cT5J5qHcSoV8t1qnQh7GRhABE2uToqa+0cFHf/Cctspr3yDubIirid6DzICib/jE6iIFclyeOc
Zhto9NNP+ah39AYvhnOnJBFotnw+dN+qjlVeQdb4U0zYpXgDerbJJflowQ1qrz/z7Y2hBSAwZX5t
afuolBpakILslDi4pZpol0dNAWR5NOVfDEWDRiSvUNUtNDbr6kNSi9+4y/dnFD902y45yKljWdTi
agRTXT75hI5PBlX+bs1hy9SeBkYtdJcZ9Ft2VcOqZeTtpQgrWqo1kCbykczcAOqZtO7VX9DJMniv
bdXJwDqKY0yTPvrNvOWfps2cKUFf96SQtLfnO5fcxdThVAkSsWlOynOhRI58M5Q6b5FFwR6a8V31
ADksqPvfZeMZjwFtgOy+8YHfyydkj+3nx7UnAU42z+xFy7ATLLWwYSq25beEsQ1Zb7CeZOiDWhq7
7DS7hXBp2PVFsgDINpZ+MPgEjQkn1Z2L0cEFjhlF8WnndRq6/nPy/AHlhdMe4jL0xIaTS9C3v0Rb
vLuNOIPKAFA8RDQe8JO52a9IzxcegQ7ZXwsn29pyPGpdnop8Ku9zSdqfOyrjF6JWdiL8EqqKBwNA
WgrZ10wcL4AKUANtuV/kEaa0q0HUSwDh1c9QzOgh404frsk0zXblrmhZ97msei7PHWYvDwcWRr8O
+nj6FiA6+Df/39ivwxv0v5XqLIHP88ycZoRFINSURYv842nwwLohY8KPKQ04f6EQFZMjk4PUAUQP
neOpCWolYo69h4wWwHIO9KCZD8VyxsIxE01ZnfXSkzmQMEBC5J7Y0pTL6q2FrTVl2UOFvM/UTVIo
HGrXKwRtjwyZxqRyRO+kTzhc71rEHnUS7PZvlDQGiquqwwxGDDS3Gp3jJEDW6SrVfahzxOQzCSFS
AlzwWNG3o1rOk2TaiaYMsJooKTkHFSFGvnuNV9Z/EbPi91K8TEjd+Tigp3HbGd41JDZUovFe4qZ/
/IOZpvFoUGrOvL3PoPDWoEmxqp/X2ToezfrVZc6cOEe+B7HjTGil8PC3Em7B4iAH0XhmXQSnae7V
5nURB6ClxalEzoc1lJ/W3u8yUtFZQ9wSdN+DMl3W3uHV6ztAyPEFWYGUQiEH4w5lJZuPlftngOQe
od+6of10fmyJLVVu2riT192h08fayiFmQjy1JVJ8JV+oD5dMMuu1uj/ZaTT6+cvg2Ano9cbqy9Gm
/0lqAtBL9peEmAdoY7vwRRWUusXJhLMI1yUajR8WbykRunYrMp2XginhNUMETb4RF+PJ0ilHp0Hw
oNgT42hOxH4xs5U+nlixNzlth3Au7E5eHCBOIJPIICCQzOvwZzg3FLV+fA1cOB0AUJOle9wiR0BB
qQZ6pWGAP9lW2EJANBDkKRZ9dagez7M17l3Tw6YI9y1/YRajPJs+3+KH5bBUntkkuwhfaZOrmEmv
0+thXfwRVOYdF1n4WGeHs8rP/r5bVWKDKvQSpjPStpe5UOgmZw3e/XP9iSWCCUfpPNtUEMxVbB9Y
+qXyfKl/caKIbRV7aiSW58dryGu0ev0XKnqKb4JREp2i0pk2HoqS47Ykg6ryR02FDABWSaXsiCVK
hn4tXxTvSmxqpf893iOsYL4xxt3ph8mh+enzUtFQWMjPv3TatAeVSxuNW/x73LAtLCytYhDLKYwi
L6i8ZsuLB6+NCdxucMQmU1kcgOwZ+cDnMD4NfryhyOiJIyG9L+Ai9+lL4zfWdVNrIOhjwe5L1X+Z
hnJ2yagw0CX1QfNj+wvBezsrJLzNga0kqPYkGD+P1IZrGRvj47zZBHZ3toqhBfiSj782kqs2dFcl
es3CT4t6KrwfDtta0ItpeSW7PWIXgKZJ7Zrde6jeUh7R17RWmgObohURIhEpnLjYWN3bCaofHF+Y
Joz01t6XGLyB5G+SU2tgQZybKuxatD4lMpMbFSpbLlsInnx791nUfe5q9IJsBLuwbUHMDMFM2U0T
YSFg4WzuB4vKUgjI+DDN58Ycno7oO9XHGAF1JLVIwzKgF/wg8QZHcFYq7K1fbKuwrkcy9jh3CinV
ajj05wccTpklS/XkWcpRRQE3WomeaOP17R23lMg1jm02h6DX2bLhu8qwWwhPHBwVFqY3zQXGRYSR
lLv+TeCt5LoYIDBl8ekCeO0PErIn4kcVEADe2nt/P+TfCsMwCDAZIcklK/aoIPL0LODSneJpRu5x
ZowdUQ0GI+5ikqe+JXPIYPuark2N5NzSdyE+kB2mE8h6wEA3+0PVx/6X8eV+8amjPZCo5fUugnpl
80PKAa0MhQMsPxcyqXr4k516cAiL4mzAHF8DYN8HZEmv0JK6+or7lhyPfCAyKLvj0hry14qaZWkL
GJdp0FHZA5isD+MHAW8e4cFXgxOTGc4El5sMIQunQAp84I9dIOSm4WLbp0/8tWBznXDWVl8wqyI5
cxJbVhR8qwC0yBjMPuZY7C8cRTgoR8qghEFz3Zw3FTku1aT3UIZH+0Vfu/8ZIh01XyVo9bquhhZ0
APS6R1+csRJOJG1awf9NlRAbjvjaTXJHnw9mvv7rT3SMDdWB3TmRxS8urljPBRF50mzHSPxb9vS6
UhYf2gZeuE5nhM+Cnc1qCVubNEuEZ56TwQi9G3xen9TLFqTxniYzIbws0McSrzC4bxwzgZcI5bgF
dzradxcHPD+NdJ7NiCnaiGvmscXp55Nqd//qw8YSvkRyfea0JF+YXuKTFL9cDsNwHgXtodEhT/PN
3xlCTZ61es06hRh8/jr7/mRW37PK5Da39ZO62+vQOTff66Ah99D3r2IVrnVcC2Tm280TDJm2U03N
oW1ITmxhdzY3ROSJAXpdbwavOvyieTa/LNeEeomQ82iTGWcq9rQk6d1p08PvvKJOcTOIie8Rl2cL
vmSbQZspwNG6bYL5PTxbA+DI+TYqkRavidPEZ/4Pcd8+EF2VZKxzQQbpdATI7PuNybDjZN5MinA3
W3y8uV8DmGdiRzzaLHCWQlsD2wLdIRQOt0QmKdFiNHis4rtRpJWP8HyBbi7gmBy1GfFDGWwFOkBH
yQiV8T5CPiGcPeQCFiIhWiSUFuzufaLnu4f7rLe30Tc/EVIqvndW0bHFtHOKazTKFJsj4JAX+hIO
PjpZjC4+GJ/Gz8rW/J9yTyFrUnYN8mi9cqHeoQ7WOmK2KFL13p/K/LJuGhzXK5qIJwI9koeHrU7u
XM2HfBpk05wUQxBy+rS2d1zFR9GYkCFSXHu13ohMuFxI/SYiM5rQg4EXOkUUmDaHhkp+UOU7rW5d
gLx0lwsWaqcKTO1kOXDuLzLmwDUMYceWtq7sUIz9+lF18sWVY2WcrxCen8PxKI3IzqqqBrRJ7Sjw
WewUOisqfc+rJ0nOu25i4Mxgr2A9M38GTgrn5yXM44aAxLEba7XEfTE+Dlnl1tQ2JqAIO4/kvug7
xsBNU9AJ3Di8IHhD3k4rL3ctkYZo+ZBTOtKeKJVPvQdnsEpg5j2ALjcEbt7DX+nKo+TTpxKHdKti
dn97JIUdkQgtKVOMFke3DBUOIWaikpezledTM7DDyxWlvq4NMVgrdCF88kchbuYEreSoQTyjSe8g
NnaKvPrdJb+4xFrTlSne349jrSP+YYwcp0UhgYi5hOn24PNQgm+yygevz24h70tfWkP1stDoL6cp
/mpMe8vEVuszznvsqjVI9SvfFxecYeRyX/TojAQdbo4nBZYq69Hrnwvx32+idWecuWdgGdC013lb
n7mfxPieqmyyPbSgH0FJ2SW2I6yDWv6Uosd0EYTT8oyaE7VHLy1ZvQ1/RvPFQ7M0Fe7cxOTT/rPz
FoN+BeyMmSdCiPHVT9Hl1nav2oBpGYA1vhX0VO0S3wwYr7yrJY7m4VtIdWHHH8vJsvkYIbRmTzG0
3WXTgqGC47xjS9rvS3QXQZdnaDLsRb7n6sRWdByHW1su+26nP3NcKMfBscoFRCpNVUL5s6yzKoTV
EW+LixglXkx5gWdvGGwNkybVa45FlfWusAist4o+JJy7lIwr/hQ2PVrw8XLJEtRYIieDYTN+R3Zz
PCqr8XOiub16K5MwTT+baVDP26hhroFprVOwEJRKD97j847wxW2ETLxheDwLlw1ygLlPWVu0Boxe
k4FX4JV7HPSPsWVK2v7Sz66zKtflCzsbhE5Xy1zkPfr0ir4nq6B3HeSTeO+bO+XZGn+7gG8z1acI
0HU4YOFwn+EG5n5wjMNURBRNb3sw59UP4Mkfrrx9qvAXuA+IwwnB5+TT2RTZUNtL6Pi2amgjtMUl
Dx2VLwWJXTIljIdqgk/xDKAFJS+aB0+rjInsuvQ8nUlCQGPhJaXg75PN6M3xZBrfvixzzvYzF8sU
ZpthEmqmwi8JiKjxIMf9OPxtBYQn8lWTnuDKKqIsMjbBOIac4F7lJVJLSXeqemJ1GyF8HQ7Z3sUr
RXVX/ktI3YOG+4YVB2yqViK/J8OwwwdlZvhbt/pFJkzQpVq90ZGzfLGxO9gxcp3caBPw5biKfRBh
v3ibDS2ypz3uAuBRyiUlqONuFoZkAGRYXRr13zWd3XYVHSbROVCk+kbvu86T9z9CxilY+RZoIMx6
GyzfOMB8YXWJqr2WyevXwICMilGhcioqqV42+8oxzprBMuuoNAtX2cJPJ94epwcVA+NhOkq9MXif
a4VJ1qojQMlemTmsTfWjxb9OGFNE/+3Z9XySai8tI97YMeqLmn6eMmY3hwmKROZfHaHlTQNYywT4
lGKrFSRrhdBX9tOOetmFr0o5imlpmp6VFynE00lEIKmnQ+HzTDbgBE98Ddm7msCWtYgPSnV26HU1
rteMHpDHLEWZkYy+a9+NKkkemmyi5c9yrWP8vcyVbJRxmdIGdes/i53NsvDkeKtZxF5DhECTcACT
trwCMUGi/aZ1gOb7SXQnqhsJ1IBc9iLEb8DPk7At2C6XkzaKPjKtHXMPcL7e9JZElbytCnl9jvLS
nWup6Xs5eP1XjmNq1AZAsvmwzgApUOEArsL4nCLdBmXhA+ZOIUL2odvR9SrDNUiMbDyCQIxVvZz8
r202ub5UdFPRAMOYVSDhVQWZqbPynDEM2+9p4kguyIVwE8Fu3aECmi0+ZlShJYngsxXOlVFpb/Xt
RYStic3SSp/9UhoZq95ZWU+3/CqObk2jugS3duNmlTtt3TvcBw2yu9Dxkj3Ym13M/1obKeg5Y1rh
h+/PK8fEnpnH0Y3xjf7iFSwI3eTWxu85x9QCat/vCZ9CEol00ItX0R66qwDMbTvVGkEZ1hWStCx4
wEdfeyjG1fMxsSAFnizvPVMRXZey/Cb89lGuluDnAbmf35dakxtsLZfYoC4DkrJnoFiVtAfWWwjv
K1iv/b9NZUd3GJ7thLcLsvay1wDWeYWOKUH3Rk3AxWPTJuZuwwF1YwNM+RkaF0cIS2mVFMwSTxha
w/acQymaqXqvZLQXMQ3mVU7mwsXNYqmpULiIbqv9i/ST3gWbDlL6JZjftiz03vQ2Az23aVNmeZzz
MWp3o9ZfNb3x1Zh/Xsj3FyGbAP9IJwgGFV6+evzPtMj3/6za+4rmlqxHl0DM/Sb2goDF6l5vs3he
qUwlHdKRHLG/c1/3wrb580Ow4J4OmhgqlNgHFlnZnvVwi2sh3z2ePlHWq47mGQCVDC+1b0We2hjj
ogdRFEtmEpV73ULAIHszIvZ0HWriLES4ry/rnKFiujU+xg6Dv0eXrYqmGHYcXeyLH+XDFL6Chh8l
3NOEUconJ6XfMPHhdYa+eOGBE6UfTobgPetnAJGX+y8id0+9sv9pK6AIMRMU81ybtWUPFW0uKFXA
ED/1MKk1IT0hSTztlF4tJpF08zgLP1bG0+s0rUkqO/zdzdCojVKCgZ8upNVzRwGh8sGMXUHlfLLx
HAmOM4HxzL4LMfLr3Elr1AW89tAho1ncnZ03aEUBS0K+fXlFA/TG+xHJ1qPwAPlf/YCfYZgsSaTc
Oh88kGtLUzUcUccSqhtZC8QeTEvsIVvuqa1au5G+JHh45v9i38+O4Ho58J69XHwChI8vtJyp0kFJ
Cf9q9YY+J1HzfXTY7ZeF/WK3ya6Blg9u5bfc1apobShM/q3ZPKEWvJTkN0A3l+ErpV6lBjQGFla9
hnBEwZMKGewv5v1SLbZmuNfcnoju3OLJnOef5z/3Uv6/stRkPCYxpQ5zG0MxEi+aj70YFtVc+Nu1
R8XkAO4aciXBElsboqMWx/Ge85GMlL955vTSck3l2Sn5SAG1tp9cn1XYdl2bhC9NfZM18fAGkkmN
S7rT5nTn5noyAafrONHAg/A4zrkLq8KZpugdCwpDyRW4MfbHsw/RySRYPcnyZjqBNrK3cnqMdh/T
KDOrq6H2cRysYGmaD6XGSW1kQ8e+2jrapLOMER5Apbm0yKIA1/pW9rYry/wkbvO8D86cIW4OIrIz
ZZwbevsVd5GzI+ZwX8xZ/9fFQ04Q+HcJuKp6xe+k+u0BjBsJba4uHXanXKMkp9JaVnzJvd/ZbzZH
zPn3tDirnuYiu/LXwT/YpTxvama9kubIWDzB0euyQj2MDiOXsnrAap5ttwzX24+fKCZme77+D3pn
SAEZpnUKY7vhmRWQkeIQ1cv+e4SReRpgSBSMvY77QZwEcVgXeWyK6wW7LbzTiYEDgB8S8Vf6/Qji
PdhF8VwikNmHY0ft+P9zaZ0iTG9KTyEd9aMbFoQa/8KBi3mdz4ao/jQ5EtlvjBpxL/rp2oRwJFyL
T3t+k97hIDps/3vWbeLrLFJ8V5SMt8cMwuCQeoyJG8O2FYD5ROdlTuh0FHajcgQszSv2CJ+TVDKc
PsnAhtljaWx2e7Lfl0bDWMS1mYOYl0s4HPEyhxH4A9uwaqrr6zUhOskge6hRvWw0SiNQVLgrRmrY
CNr7NHGjlTQ5karzNGRGM9+P52JrxOMTKNMG/bEzhPCJZF9Hv4N+9VgIBaVrJx/VfGdLfuSWFEfg
Z3GqaGkwkkb9fMFHVk2ne3upHZOswNOfyr2JsG4iEXucR4G4e5WmHLzvklDvPojbQGby/oyGuv1F
plQLDDnJmDQ/BKtDiauNc+Cw9ZGOm+OWPMzRsDwDCylANgQTJk9QlkZ9IkCLAaek3+oMOxyBPFws
pFLFeQMfZXes66BaUMCCPxlQpOCq/EgqTchk/P9Avz0H7d0WTxKdHczxD4r4l0WxowkX/8N2PqIP
WMkksdn4EBCN5QLAtd+/3C8rSPrrm6gvyF1oad8/U/wOk0Lydo8B5xEwHtx3BwwXkVjMkgvtGlUc
8g4shTLDlQQWBU7+JdDsrZiXRBBDOtRs67YUOagyFqVsQuDbE+PzpEaNfABRFFne4Y31hTsaFoRg
GpmjyQ2d21NaQgniuZzpBBvjlgky/Gu11206AgIZEufi2LGN/sAJuz1R3l6VpVNpr7PgkSBVOstk
b0SOuoeXuM2721DDGC087EG2kKYVvPcvi90VShh8KzDJtDMpDm/ODg9fPa9IF4yu3ihOZf1LQ3Ky
ioe28zQruHBRK+JPKtEnzRatIoEnbPcCh9scc4SnY9uyW5XjK2eVXstYCmufst3cSBQfsBk8rxai
4GffJkzRrsW0gN89F25mOurtVhbpAqc1GSDrwkTlIT0ezVgjVHVg0dmzybLaVGsb9rk0xzwN/Sg7
TB3z0+7FKHxOSL4Xj7lSlACVnvpUYv+iNlx7Q1nYJxWUJgZudQuIWgc8463FesWtDYHm+Ecl/UBm
fm6t6PkonqDWg/Yw3NdjuoLicK/S3LXtDps94W80cpap88l7rAlX90TbVrxYgs7wn5NDVEdijq5J
UJXZAQ2zZMooxFefW1D0b1mrq/D49W6ovgjWKSJv4g5JwH4aVBcZvBT0ZlLH4BQe8RWNGwj/4VRr
JSwoQTxAyuvFr39qW21rJfJhMhKBE0ctwJXu2drigObFHfBgHsw4ZM2JrxtBZ9qWhHw21OyfGfX5
N11ZLiVUOioCzXxVzb9n06jYEeUGUwDHM1Jtghgpy9dud5R8KsBJ8YTGlnS6QDR4ZZ38zDz7bgSn
IGNICWCaC/svXHNF2OhjmqgzR1oZ/IVWnptLc/bZn3VfJkVzy+C0zR3ZyIxFwvSUlDq6InLa4RiE
4zfWFnyau63Zc8+Pod2MI4c2wJlnYHtaQhRENxZkdvS7C+QeOC1CEA68Ah5AClj67EDof6wEM0x2
8qsYlg06Lq/h0XcwkQEnZ6s1A/990GUE9N0/k+V2CgctGsiQMs5Qpo77Ap1ZnspbLNSQFvBqxrEF
N5c9qZSguPcgYnmwu3NXf+89jkdmCKBVL5HN8pqW97jpGkExXVs9JfM4lvh56S2FFMn+s6qv2zH/
MzGtQ84ORHTGN06r2qyNVNYXJnyLcQZAMnc7TdkLvECoqWDS1ZdCIlg8hhEmA1Zv0Pk/dAvFMxS5
lr3THFmcW1vhnXm1dFUko6/XoqpmcTDJMPIQpc4W6dzm4JQZH+NT062P7CeHzaUrbYTDjOkh+ovW
Gv75GZ829FPFhBUJabK8u7IMU6wM1mwf6r69anyu+Xq58t0LZSHPMoHbxhNzPwm1X1kWo8ERCow4
drPshjL9k9TWwVfXLXi/oaVvZkZeSMMadzRJall2J/Y0tbhG37dSzBXDQOxxy3LyeeCSSioI6VbX
TstuPKcKPxgxTWp0d3yYGR8wAKEetY2QZLw2LDnntogmOtEw5Na66Y14ZXI7t3F8mKVI/y5U6ecM
lfwc7iUQD9o011zdB4VkCmfr8QNVV0B9aRMI3s+S4DgN6ze/rTq1VNEdb8Je0dFeF79zWUa6Tigp
rgNjFu3k0sijwsvLd3NEk4mYKlGWH1YNmSMFW0IdQ6OL0JzHNybK4Sanq+sanZ3J5GgcIz3EARHv
QwaTVsCKN6TpU+rlSmKogRa1u92yh21FZxQ72FGTAsLm2YvbJDJ/M8E8Yd2ciY3Cmiw57Grruu8L
pk2+IHgAGuTqLtOmsq2wf0g6GPbnuvWMCW/JfcewhjBsQzHLVlodjkOZWGqVNNMUv6sF3cKe9ksL
rURqwtFDf3JAWBjx0JC1OmpPnsHN17G7bq4JqWd5GxNkkVkNszWDdDYfBY62hYqe+1gRPXtXm/b9
gT5pKX2SDnUZfOZVVIGLo34BUSaOOy747h2vOgVER02RXBkgzWSw/aLAS/YYqp/vrizkemjV3VJ+
0ghxEBU22VCuKcn4xpLlC8EaA3SeeZhp08vQmrnSzW/OMx7DPPwmWjrkozr5ITj9fchQL01413YN
HyaincdTlK2DU8aDNYUrWrUNOA0M/UxZI0bR04SgALnAhng4oM9EnzYtHqlV8BZxqoG9zP/jKESh
VqxD8PtatsTHqEdlQcTchDTNeyR2eB7fhX6kFsFDqGYQw9LndT5lXQHAEwsnECqBGDwEynX7N51K
m0sfKEwji+9an3xjCmAaWaP/z0y0PTWDbiUCHxVcjQgj6sIbnNFJEnqKcV45QG6hNiFw3YdIuxqZ
Z7CSX+1KQHVhCSNrNe0YxvHkKE7cjzH7RtTOd0UbxemxbnbuijShBapqe10r0bPBHf25vA/Nh9e3
f+Knisgl0vMMg56ltTyUvBhbfreAbMr24bVsR6jKaPTGw/d91a6hEekyA/i/jcMHNnK954Pj1wQZ
oTcKKqsCjNbIdRW1++gOqEQCfg3rj3lkM1pY/vU3Bzrapk/Tn86fVAMdfqDbFMfN1UG9nigp7xzV
LWRuFZ082/V+gbwNTiSmPCCoPWHNPi1AGOMgqyFt477rPA6+OJtauKqzdE1doX94wpLPtyX69On/
iyWpaEENDaJpKb5rI/zSh02LijkXvcpwEupBoPyuZ9SFTG2VedHAAq5vzEgkIhv4E/yyKhe+noI1
+h2yAsC1NnObXRPMnIjRt3CHavMnybiQGUzrjpEKiQuIQOHNYk9uY62q6irFBZRIbegFT//D23g2
Ki7kVwHhwrdryDQnqKq7xWQ4lsP7762Ez3Pq6jObQrynhv2KMwA2MPAmaIz2UcVjRi5iJiLMSDkz
U4t0HS4+OsROV0ncu2aWPqPThCWnP0XVFatAMuGlgv0eOCRPSV+vm2TZiAqfrXvSdoFZZHc8Jjqt
jyBAB+2VbKdH8u6lT+fxLkm0Q5uL1gc1rZZYuUBN8Zb1fLGernmvZYDTEWNyAO55hf8kaY90oWmI
yKuHI5V8ZvXdTF6PtrTw8kIVCac391VlF7S4psWAZnJ0BqHBheQBWwDI2yOe9fgc1SynVFBSA6Im
Q5ZEjo36+JL6hMWJuVLA8VRKmUaCctgyDJ8djcEQPnWKbu2g3+9r5ENcAhjaE7Ap28Ty+MZSqg9h
av6MVIEwSCfLZr/opwc5Ouxkk+deBKETJSvYFpOBXEwY6EZdyYZBclU26NVu8K3OaHfbNqNtkoFE
Sr5Xx/HaCwZwwp1+/m+c83f0dkRh+TsxG16/FXPrLEaYU+QWxJuveL0F/lDyxda83muXV7E63xXR
gwTkv+VQuLPk1UvC6GagQquTOr1U22H83qi67NiDgspGrayfTCVCcOo4uvL197dRxipP6tGlQ3bX
+tQ64xkr+3/2Fjb0CjBR48hyLcDj+gRKDY+rh8Qz9iewiPQ9LlNum/0cRGwsVLy81mOO7TzkjWnD
dWb3sXMKs+ENk2i13mVjUSHXOXN+M1E/HyVRSvT/WogothwuJguEbuELQEFI8qzMZfGzkZWQ3hYZ
Y/Su+5tUFUoQTZhKwK2ZirzqLOyzINBUMFdkZYm8XrezdhfFeUcfIibD5WJ1zW0CrzX1rw41rw9U
9UM4gU5Loybze8ka3fN6Hc0K48cUxBfzd9YsIHvNChK/rQwwP1kXStOTi79Rr0tzhvRDxY1OPC7S
M43ZAxO/z5dWrCkg1ceq7R7/k8kS5pU1vlu8jbOH3guVtT5Hx5+jDRbJNV50s16KGlYPIzHn/TWO
1/kiXKBRHt9ZkbtXlNi24g78gdQl364BDuPrVsRpKNYleRfc4YdgpgNSAm2u8mZekmcqxJ4gwjbF
KLRjmB76yB6mN7wuwPLdHzToZII15IxI/tZxXscrk4EOiHwDveIuI4MCeErfQ59IO510zp87E55x
ucN39mhPdgPewapBmdrWPInuhJKu/C//ArLmFRDMwGq/gRUADMevVZRYjsPJDLJgPkS/esEL1/o+
Sote4zpUh+dlsOylbg5/U95jgMc2C7phDLcOu5xtDM5IshU2UsvlRKOkE9Wcr30s52l8mW6a7fzS
3TciBKWh95WgUzGVLQzUrjNmHsMb90S6QzgMdUVTE8KcE37zHDbPHjMVYSePVppxJju70TEqVb8t
hyWMPn0rGJzQdRr7LgBmfqtorxynjiCmjXS95pdbNfSR2fm8zTD5pYcgBcxBqxOSfkt/SWmsQAF3
+QJmyYD3fw2+qWsepwHa1cjro7GKg2mVvHt3uG2dVtH1WYtsXkWlw9WH9QNSuoIEMZJXTHDdlae4
A/Ksgt30yUPUNwQN2n7viEHiZ02EVIv6gVrwgw7bnHUzd07AgSDj2Zo2ZAzjA5XLRtlO5Ta4oiO4
QCHZxaz6YVy8B/2zgEiPpMJ0TesXG4no4gLDsg4a38/vDR3bxjHCNwt1juh6zdexOlkB5ZpQE7KU
4ZMHolnqMWAuppLuYn19r8cP+YNmrNvUoJyqBzA7B14k3bJ0/qQ7wI0dWS8x97iX6Qc5QA/4o4V6
DSimzrGrvg6Kucc9CCmyVleuNluhLZVRD973XtEzwK2HYXmFJdznDNDjy1ueMsk9Uu99AOAvLqfK
JbhrYSySXIgcUzeVv0Fi5ui+NNRyCR1SaFdOrJJMm5axd2VwG1DtkwRh6AJRvopQwWx/PEH4uYW3
em7xndySKnzpzDBbRtPcB/Zv0p3K6z3DK3+jENGT7D5L6GJhC5GGaJCZd3NoQq8PodmgMCJBeves
6hpnwZmVUAprZrXuYY5txgxgBqfBnquMfuApydZnSzXxii3PWiVh3vWG4aSNGnRyxZA1DO3+Wv+9
OkR7PBXeotgxpH/JDtjqGeyd9i8dHLzGHZzT6+PwdAliRGFvffelBjZvmFfiH7EOUhx0iGHElHAj
r8B/NkfwQ2GD67n0UoArrLbUSPB3L+wGGJu/N4I0BF1XuNofoaBxd6Gj4QuO+1mIueQkUpBnllh/
TgI7QIlW2IveOgH2u12MhGZSw4IK/NQabiFwbwvDETm4LhC4PUSVsu19T1WF6Aq3LlVbJdod0hfB
JXeeNQFJ7Mpstt/XKV/GojfMAJLA9o6R8RXTOdXl7sDEuYGe4T350unQCmY3lOOJOXMMyHT0OS6s
fRC1UDX1zsCJh90t2/SumO+mUVUeuPsWBsdweDDZLRpRPZLSjNtpltxBaGqAozbsoGQitgVKmbjR
m7uHIQSCdSRfn5VLuWl6lEECNiHq9gmu7zCXWLR+UzQiys5a8N4aNMl1r50ghovkjc0bz+MBXQs2
GACa0Ke/vEr1AGQRDqliuD7nD8GYQ0hnbLPK6usPaiBeGcmzemOYjVqQEIxIotIx/CXANCgDyGrL
NkvjlFWfiW2IXtzkw1YNWLTurZVHEHpLjxXSxJ8QYgCPvb+LzPhYC1cOp+iBE+Kx/eUGiBifzVf8
S/thqYeGrQNviHZlIc8QnbYXYImrVaWYVzLTudoan0hSnWmqT8ny4Q4/Tfn3DU2hlOISPuf44oRi
nr6JTSnHUwzJyum1Y3ts3fefhcaAWKCxcRUFIfdcLd0IE6eZnJ+V3XJtvwU6CqnCWJchsu18iInn
RC1ovS/8vb9I7q5snNQxd59YlXPtAVleyWlRpKpL47UwoI/ZUDWxgUooKKJq0x7xKKalRKk/9QNn
tNksWiH70Z1y69IFZcl7zlO4ZtzpHWeO2K8fOxExjTm2zVVeNwzvOYbfkfuStV75LfMzGF4x3rhV
docfHayGh3CeiItXBdlr4DSiElhYnqizVefdIY9NlJBDq4ArGwLDKcj5nxla6Zi3TOZwE6S6arz8
XSUxOFudi8ZfoYatPvypw4DOF3TPl7krjSyyYbpp3y628FKqyQUAuD1ygpINBFh1WDBp3x9Sy30h
UjfotI9LE8FagsXtYR+PRBeO8DCom0ACTmgin/5kGXe0bltKvLoKI2mld0+Xhjgkai/ozal7cTuR
Twal6/2Hope/MfbhiWDRJG7GJzs+BDIRGYkmccfyxlIWSRUgKhkLEaY2BoaY88zZLRfzEC/eyeyx
eooVTxJ++bTFDePYAbFvisN4wpWkmy4kkfxJtn5JwGo4Tmw7XB7qqVlY73VkbviuUZMlGNNT3mp3
L7sMCFP+L3ZBB1bLjhjjWQb9xaVLCkUnVG2b12B0CbiXl841Jc4b0iV8oN8T9kwqVG2Muz3MCqK2
tbbbBCe82ADd/t4Xy6e2d4IV4rQR1UgJlQmnHZiXERX6R1ZqYc/DPoz/RzTngvYtSRU5ENjOnQaD
I9fUUtHe8cNWPajO0dGr0IcTCbRYNnUilkE/esozdjWzXs00HAIBy7WfE0WCNB07C6GU3jppRha4
FvJKsu7nL6R4+6qT0hzjUDK8HWfzTO2kqV18XNFyW5euL3N2I3Zz15Lz2NepL0prGcFIu42ESJrh
PmGb7JQoxPv6OaQoHeiRIDM2RbkM9Dvnv+JC8S9Xm9Y0j8U4BN4YU88JnuJ+SVX8XlOdMWdak/pI
4CcKu/AfT1McEN2nSFFeM6CXlcdKQYmkmnhw/OfG1wOGWLwnbjuuhhYZ3nAGquNxat1RKO7MvOR8
YxIWAG49fiV3KXgGRBGb38Ax321l502v3Ncl6ouykrRnVwwrkbYHNufXn5E0BREI+Qd2qDoVRfQm
YRwsDM7L4q1RAmwxn67fZAxgln4ztE2DssxnvCpjcApiX5g9B89+u+Mffgjho8IS34yLfUKZkk0N
objqoIG3zIVx/3nIdSfqdVsczTHQv6bEY4D2QIJtxwfdi/wNc6+dlCFO9uulV54og5qiStpYheEw
cXn0mimqq6jj6lJAKUjWRZeRvN9LJFhH3gFKj1JVptUm7c39IuWpBo5XhnZl/UGtGfB3e9DQ9pup
iWX7VVGDmQn+FH5p74oHoCjcQe3qlo6Mdgy2ebzj+iuXjFFIUKkAMK7gx9Gl18pvLO3pxuuOY6Uu
+JDuzez57m6FQ0RRg0YXwqmh/qmTeAMJJwAyg10C2+jLdyIjGSuaebt0xF8UV2nhC1MOasXc+20c
71S2cs3j0n/AhKm0AqU3NMG0KGkym/GJgDJx3vuG3pkB113rNz1376FbJm/3C4y83O2SkdCWf3UX
ccQ9pTDg9C4BVG3ZndKp/1cLxnHC2P0lXdGl/5/3erQkPAL0RwV+ieTV3kyecfVepuaL83GJxpSm
hilBDKNg2teJTXGG/SG9azB5nCBOcrqFZLaVx7MAY2MlEJsTDVdlUWQ77jYpJdg98nkqPpqgMeBz
LTH+gwDn86WSlNwK06xUFTSLELRxhG5Am4f/qGNN/8we4H9IR2IGOAVf/6r9a7cn4yMpatT07GwJ
M9o5Apr8cbyKKFiDeUOTauvR/Dr5T7cXdK2Zx529o4GZo73n5Q63pUqGq3q8ChY+w/lCsCbHXASs
vxc33WWtxACcL5+rXsf6wmg+q1ceG/eho00daNU4b2iOkKqgJ0ZqVWqmuY0FoDu1LFNM9To9kWYD
Z0JCB0bDUuInEgN0Kl+OKc1UDxtSJhnDjcYhennhtEED3ndJHwC2lGjuzdDRTNKQ1Pgw3Sbu6ZiL
6HevW7mkVbVI8170sW917JXegsPlTR8OaJRvkBHTQs16v8Fc8fLS6Lh+WDs8awPTy8Df/h0o35LX
I/D4+89j0RJSvAKl3DAL0VcTTY5DvXcLcx0Mn22qf6CvjlJmXBL8EFqc2yQbrbUOqmAHDMBuEm1G
IBsCTGrAtl4EjcHpoQLgF2/eI4SlXmeAG0+pmWCeDTpoIUvx4lF44YVHho5yOOi9UfCI2mO/GsR9
29x0DSA7sUZvntr/txe8zSZwP+D6wHE2uTKHtOm8Dvucy63lpev3fEpppxo8VE8yLPwjBOYikTBn
eVwdRt8FYWxZRQMI7KWl9FT0Lq7s1cylagWn1vOlkTJ8sJmsrV04Bw8bSRD6b/68fW6oOX62QnnA
3CBRvVbskJLKcfpukYFnSFPiQXd/0Hw9QkSqrjSbeYWX1OMIbXsiHUDor/ImGWytbjASjdVGmFd7
vo+QayFbBMqbijBZyYTv8mLSvy3wbmDWOSEzBIrCqXqONkD5BeTd49QOMvTjmkuCBNjd/bnqJ44j
SpeGNHNhepmQxDMmx9X2cROctVm+dICNKawoPapzXpxuN3xpQaLer1kmYEPFI5dxliJb3LaSEeiv
qfY1qflanH7gSebFVpRGMpU1Rjy0sJCeX46cP0kmcj4ZVU6o7AbzPt0t6y3JI9AdQUphFpA04B6x
TYFd3Djh2vv1Kj7QO+uEBVkizQIgqAJmwMsODUUqOKYV9wJBzKATLjR+nMg8IhMRpd5MvcYlQUiN
xIMVyx+g4s8E3SFj0KlA9PwHQcZY/4G75wxorxfQkwMVPXcZvIOMxQWmHhP0tzZzXZ3wGKpGACI1
VCtWgLCxaRlhHcU/a6AadOlgX6bwG7n4B5O+TfNxPxO7cD4mZlhXWq7SZR7M/kf+Zt7d8dscT8lx
QcuAgsoep8diVVLzvM/HOMHc4EQjFR92dOy8CRfIkuRTJyXw9Jx8vvMUx5Qa6IZfTp3p6H6R8cce
QLQ+E1NbDikigRlgaJO0FzG7qFzsEKdHfgg1AxyksCKpI5Q527884W2qkOKO5IdD6QbJ+m6aJ7z6
+cX4eEdlzrbe/DozAI9i3bg/5EnIJSsBzhTseJJR8qEs8cnjgX/ICqBxj7qHV00X22jpecl0QczG
tTa7ocSjbGgA7pt8DnBiIwFY/RuLPdVygXD4gXBzS6JRHLTASY7Gh4mdaFxUDn+P3zRD704HA3L8
Gum3fmjUI5RnHiRTYal4qizhXexVasEs5ZUg4aQs8Aa15g9LOTfWwq8giSyyKKT7M9GxViC42Jrh
dAPSnTDHFbxZRXdtFOftLn5QNkMHt3PnvxCtCA3NkdPi1v/sisXdxEh8J0Z6R5T58IXzvyZdmNls
p2cp63pWc8fClDexUNNOPWER7zjG/ReOird3sHxRrwsrfl6nVoG2Pc5YKd1xgem0x7c0VTKCpnIF
CWiEpPQ6XmFSGL+Z9cAN/D+p1THpbth1poRwtp/47mI/BXltVQy+tP3tbU+RBXD9d7Oqy5Wq7vQK
6h5WFK8b70oH+r4/VMknmtdVWRWrlMvet6oI7AjqkAnQPqYP2MR28E2EuUUl80WSXO1K7d/a+YqC
LK9DPoWFcmd3llV7fhxbSq/vIQUqM4ipD4qYA9pPk8u0prCafVgMcv/VkHC1I19vZFPf9MW9nf94
05q9/2iB28I/Q1kC1LaKXaOGYuu7XBF0wCGMlomcwLIEE9DxBfn+lcPzTi6mPIo+t3Tui9Y+YMkH
yYwVFs75DK2z9MK7XHASiQyK8foiaUq2y4lpuPY4du1B6p63n7JTCC5O3yaPgjN2uUlhE4B7bz+9
BFey9Ls35ueZvagxxJuUypXSZKh2hEos81fY4v3U0ZJe+4pc+tqASPkcijhHJzxl4FlO000Q04V1
+s6eWYCLgq95VTunjS2dE1kL8avExYKgFMpo94u9oPSFG4CqFXPqKajZ5vuBqTKF9Oa3Tv3oA1ND
D3bRswdajC2dCJRckO0W5xAE0vagQrV44+yadnRa1tok7tuc4zp1gFjGiYHbhJJ9oO/f41btS98K
bhXS06wchTu2MhXbhOxvYNxhIWveqOOiD/YLn9I3svNii1IJFHZNn3ufVj2HcRQAf8DE47nWpapj
zpJqpMYMbco4JTbQO2XHVmhZ0ieOtoTqUMecTKbS0pqMBRLhYhlPo7+LsAxiBr3vwT2v40zdmc6l
++hzJpahJnY9tNcY60q9rfcjwSSHq7KLrF6DIiiCBdmTjpMO0putV4AGGJwozbOuD2A8gJARrgj9
KhT97DnyI+9KHuSS0EfX/hkLf98adDu4RP1MCRqL1C5iLilqcCkBzUlbxQX6O9xm+rr5o9IOAIdy
owKEpL0jUdPhUcQSfK+DkF32AP9g0WEk0S9c1DTw78f/GrQ0CpEB6KI0OfU4RhXUg9fnuOaaxR98
qQJqkbHd7R+nZ+OAndGq2COs5lxDOHVd9dSxzWJI/5DRqYAuM1qlfiNgk+pET3lv0smlO0V6cauX
0X+sE5qoaCXwcc923x/aOqEkDDVVQ9XrxjXUFzuSXJkRHZW74AD+4iYYhVX6zOT5LDxPNbjthh+E
mv++VOshcOhVjeddmzP4OfqeoUBtYcKOsZAdZDZFVgL4GfdiCky64SP4nmtvePvwUzU2yWjk9E39
qs1lNDJWEXc/EpVKlTVUqTVWabI8Ev20iVXjDxCAm8fseFcotx0GEGYhSf9L/mEuyhjki2LtDHdH
lVPnOBUQKsSWaLJ9XBxyloFCq93crd9eT5qoLl3aVY+bwPVZAOtGVduUwmpCQfl4NcRPtASw5eK8
lg0slmTj5S9EDcCWyqa5PWz5jahtDmK4P1N1pmqKbZM8c8taytjKX0m1uDf8EbOESTYR2Woo+QkA
hqI1DVbm1it8UkxtZqvrq2ChZ6XExrAlm5U99ToMWy67PEO6bvI/53lviZL9KnN/igtwjs+XUYSM
ilAdZcubewdNGW+/oX1sbq8vE1ta8jRpUF14UvxNZla+cSxwQ5EYcyvUEjPZi6H+BQQVIAppFYug
ihwriTABE9OJc9QOVroy/4YQ1PAEAEE/kmNRg7yW2a6ydOBFqdvcDO5fhKjn3PUv6mZtzqfAGHfq
0fWEofSybDPPEvlcScV/wcAQFLquRTsL3T6huEkc2IZtAPcFGBKuUyBNe/x59x6xi5Skk8ukK9sh
i8M3lnvfVYzlLX+pqctpu1dvWhD96mPdjEtBCUtystOMJOyxAc4RRzYwwNjv2FrqKGs1LHX65Ouc
DEHXxR5fblBvQgkEraVcZiHMCuFeqUo/haIAZX71ct/Yr4zdX3gHsqgM2M+G6nYdlWd0k2nCvx9n
9AX+E5ktmktxYJe2JW10gN17uLTs1EnL4mDrHonUXI4esW7SmLGye/2EmtA70Xoy0uSDDN8fmHh0
9kHnxSFS65rE2bKZzRtfMi5VJ/AElD65Ypz2BQm5arTw5SwKp/ADoBMpSrcQlht+3Kmh5JnwNr1R
L4Lqko0UN0e2N4UOyB8j8JyO6HaaoeQnzdGKvDeo4DETolE8KvDc27p9fdvr5GZCW2Pb6aAw+zRh
2385ri6nIM/s+UidBU5Ay90EA3dVYwqGPfgzhx6gXp0PAMvtw9NCxt+c2mliMtzMzIJuwMErC2X+
IOG8aHFkP2MM3hYm0r/DbArui2WjMqqxcwOrc2MkUF1pQjrZUPG3n7G65DhXBh72JzXhJsWkSm6P
ZbrMaQgmu17yErxZMmazmEF91Gcv3JleApDBbrk15vAfiEhyrOxoNdD2VKz/DZ97e7vwFJxXJMk1
wc7cgPzykvGdZ3T7DVEvss+V5RGVaB90S/a1m3OPsi20iLUgA1nh6e1lgYmq10EESiSEWnHy7iEe
qGC1f+oFC/W7cUmoc2j/h2S9r7VeoOcH8r/HAq7OoknElQcrwp9jpR1Y4j998TpSt3nLcoN1I7P5
BcBg6SfjzKbP0gJ+pMB1j1kULVW1jz74MXzlxKJV2PqZSKH/b9nomOiPeAk6jmDnTa73Zkypjm6e
iG610ST8mnAexcDuCztUDoDwpnZhocvAQVJj4mrWAs9GZaJ4bjjwxIebwlBfGbE4iYAHRc43WMxW
+r3iLvgE6ZJou2Gqx1/3SCOySYUw8Q241Xfvysbqk6lrhjVIRbx8bdNj2p4MuGohKFh9xgBvUxjI
8UyGTsfJJ5GnIQWxpTa8n0earE7tXSNKoH+NhDov+QWxO24WAjG7SB7EF+jGg6UyLNP89hU53JY8
00lkx8BS13U0OcKyIBY/Z/I4Wv79vP91RCr9guL3X8GXk3F6blU9f87j+hgVBqL8M8uLs06iyyBt
+9hqrOfnjRYxnGGFlaL8ejGQ99Qkrmz9S+vVzV5RdN1AmPrYjDT/jV1nRMvX2QAvEqaYMLb55Q9H
nejcr42uQ//VqGVaiPo3fXYgZKx6IwUfK2H/tyvtdiOAX4AHMcKkQ5RBYQU61ojwvwzkby8WtdS1
KPMxATOEagh63fctLp8AAZ5Tug23m5N95UtuDY6vzCC4sLvfBiwv7mDS7PMiV0+HDoBhFqSN3c1/
plMBy1aolI7CUsqpMNO6hpuiRCgLJzPjvV2dEVa7jrYgRUK/Y5gi5X/TyhRFrCDRG5cGM7fjdaDy
D4b+VVNrRZYH6B20ZN/ujBEMRJAqBbdrjZdBnMco7Ujmu6wAC9tpqor2hCR0N16wyjhwMVvEvTg6
s47E0QfhcvtxqyoTdxARp7POwiJ6q3mP3uVfoNGtL9KUBrN9kA53ViMZrtKMb5OgmFFxpDDD6HvN
dKDNlr2hHY6Sz9KSsvIo/tlK0arRWDTc6YlkOtGLGejFALXYuiEfDzgcf5TgOzn8o2jXhcsr0uuX
U8csZryXFWd1J39Ngr3Au4a6OV1wp6AbrfewTnn0su9+LE5JAzpGmyM9p2c+Els5YmIFmB87JwQU
v+5RMVDrqkyMN4MuZm9X643TxSbdbEOP49LfAKBrbbKvEsY347XuxaZf2/Ie+y+QYDmohM3XjxHA
u5NYxvfdcQf9QaPUQyj3RSrs6yBW5VTyvf0tf8lCLHgRhUYwlfsTQX5VOEipquDEu6Y4StRlKwWF
ybeKP7NilZ78KAH4wa//3fESWKSGmPv++7ONRJGOBzjE0SjvSCGK4VmJvxXIGhOyfDIuH2dtM43O
vucbSKavy8kyXRKHMTE5uCaGv04foMUoUfcDNQhywWHYanhRlCDsgwBcSWQYhgg1zBeM7DGsMadR
5JK1ptW6hudLevGhXRrIAx/M+/OlzJ6nD7tckgX4fQ31fOwoHvnSMa+egyhLunlpJxd49Hd+XLyi
50AJ4YanVOyGWnTFo4uwFRkybbM7+qAmlzxluKN9wCK21UmZ2LMzAyxjpfa4fcOSpfRruEm7JH+q
Jr4nQ64hlocuEbTKMSoCm/8EX1lf5QU5HUe9BIay2zI8sx0XQ2LLOFVjf47kpD54xHAFZ3eaA3Vd
5/SsyHgD5bGXe6j4PjoymVZn3wggKsx7926rn7s11HIsiYnXl3/gkd2yprQBL9sfg9EBwh9Dufab
uls2pnt4b0Q7Z81IRiudc9b5N/9uaYx8QTeEZ5Odlp0CmGT5MjePKNRATGmgA/IIgOTwvs4lVbph
GHJZho2xPYrGhrTRf2U0StocFu3EJRxKy1FKbqyRMhU5oO8owpDviA2ctHtfY/AmHdD6rfz3uPlR
+ncbTBQdlgZbe8r6qVIB7rJ5EQ99JKO4BuhYh8EIk6Vr7EB8DPaZwnruaqQC7J0rB8+ZSU3lhAIo
va82wth6248gkJQHAFBVkBDiW9r3N/aMtTSot3ZWxax+LlGQ/3WYGROMgN/8MBlupW4bxi/3SXCg
N4Ae/vPsaPSZtKarGBPMMe7NUXvRqpy6u5UG0wukYIh4Rwwfmgtw24FaO7Mtr645FiGtSF5dsbO6
PzO5CsZxpDAjV3epYf3S+EXgUvSj8Mk0KtX70ILjud709JLbLQIaGXuM890DzQ7FOR4QHH504SbB
QEUPcNyuJkpoMwglQKer89LgdEDLaVwEbllXrmHJIur3yODI3IWvXuU4rQeB68N87kgGuOZaXnt9
dwsowPTdB96Q4QYLi1c+gRdALtzhFnnSfj/8WRAt0Bsr9tIAYeLm7itV1772j9bukC7Eh8XPgVzR
LNonHtilyT1M9XHtDqdAqZQ7hOr/Rwn5kHhumd4hqQPR6/0ey5LpRmF9k/Spgzg02g2RiIjnBGGC
6i/KnVfVyWq1PvjhI60QVamKLbblt2wwsmdtIkpxMCHd0iHoaMWYbDCGEKXiKkhNaD961fDKdCRY
Emb0z1tqmPnK2P4sanKfvQ2RWDHN5PNMsE2VEUPxaibuSRfoNRBzW9HIGqGlurifx1oGJn47WdGv
rLRLDWf5dFXqNw6G3l4wAY8Tz0BeGA4bF8JrtyEomEyVhCMqgw178lZUw5pbCMd4AutewEFE7D9V
ayU8JJ3RgGxcFjidjE/xXyTZTF3WLkFnOixlXSbuTH6q7K8S1zpNbVcOrVAE8zsTcyM4El8xi/od
QI3vYHJaON/lmDoUij/GBZuTRCtKaISl/eaE+PIEcBFJVeyCaZ052zs2haTYbrO4f6gxxMBCH1z4
zEwE4p0aXFsz60XKjsSC9NY8GQUcGsK1FFL9+GByZsgNNQ564wgsphtqtA1/YGK3n91BQoZm7BCC
VAvLmHiouexokwOx39WApyYmrmd0le+evV3cUkWO01kExBM4ByX3P/EwMpkDD/Xmp/XeuD82egZR
prou9W8OWi+Npjk+1pybTadOACS6zaHU/dYehZtoI0oyMakyr6SUdGVxv4AkwfEZIV5xevpjmrE3
UXuzRRfLXqi3de+9GMK39NTjzYef8vni+qQ/DLrhZU+ggcjxlh8xiyeWap1rCZ2W7ka4anTj1SwU
TiBv1/eNe2EBh5oaaFgi883jzNWYvrwLOwQ1vgHkqIOqCyMK1u2xdM5oymyjPVQrPSQTi7ykQHQt
5VJ3KC1Ltd31WZ79zBSs2K9RN15rUcOBVHVLUGLZSsa0MSGv6AK5b2x8R2gBpriIYQekPf02HNR5
fhq+9hAxBubHn9GsNvbB9Fjj5GhD7LBU3riaz0zUhNKWn1vLeMrszqsbET9AxNnzkCehHAx3cU2n
8tsZlcqNiWgGdKeK8tIu1xG+WmnxUax1/IIfQXUn5nu9U9sYHjr9cAWbBBucDWNepz8sV3zosisE
xMJkMi3eUehl8v0FK1LL926tcoLv2XhmGXyf93cZe7oGe+1do7YTZDOiaUeSIRStAuzgMBkvFyA2
5L+Js8ePRQ945y/olHkeodh8AzNc5u/p9enkuBOBkoLbTwkCfGM2tl/hvPKPxsiPcKqu34RyV9MS
+a1ZrOAkDkjLDFnAmqvVekMq4HaAICMIQLWyWry1Vsy5UCoseshjjqiJj0HhSRRQPTqtRuHX3tCA
TzUnV8SDOVFu3o1Aef21KfHxGHkv3/WrD4V7f4qbFo1eGQyf3XGO3TtiQ9oJhS6iWVMLaafHqTX2
057j50kFtlt6Nazi/ifmqw2fLFOpvKB9H+GYIDyJUEmHlMkZwWjkZEtSWeG3MLBz1VMSR+ICWjcB
VDVPcxSrAhMgLMEyhl21IrAY959XSHXa60US0YW7HvPDYbrSjY+VulQb3zJiwe7yJQZtMTQI0v8M
QV8QHBwPYklDLIN2nMvpLc/RLsmA8mbxFUPDWSrnw0HtCPt4C/JZh+S+h4dsPLkZzIogEXnpMMVd
P3X3XhPT7aoT4q9uersK1hKEHcoS9YgN3PIydFiYELXlsq28t/dPOC+dnlF+riLUu7RRqOWyX8BR
VHmNnHCoiQnpZnwHqfOdLS9HErjem9VLwAGiKFrdprJLeKf3pAmqfI7W2qJOjfGk0mL7q5jkFx0J
GqKL8AsDUq9ijQVA8Eo5badHqww0mJnmez5Y4Y6PzaqI8/YgEopK+udlbVHrj4mh8hAk7srUfjrV
5r7FAJGSBDYfWuQ12oW+GGdMb/t7trtP4oFr/2MtIRyB92saDQdg8201InNz9KbBgwUsMXofeaqJ
+YLU+BiuBQOWb0XnSnJE1s92USuQUiLBciDj560F1cHEz6Iih+4OyJHyuI4/5Iz5oJTXGYaRibCN
I2WSKUztTL8PPqdzpCJGaP86+70Wzoor5updJ62bI39SWFVbxGen5VdDmpjYkBLl/xLpl9Rx3/MJ
z2sgFaeAwsNdkvFqC9oUheYpAC0S/cn/jXRzWsgIZYxPqygafWX6J1FJZOUmUPKAUOvM9nqOzuB8
ugsgRaofMcCisF05JBTMPU4UD38tXEnOnESBEiO/MXk9A/u3EbWYN4IqXEtirQaz9+Bk4eAPh2AS
QYNZq9PcUCXiyHsJUkEE641W3NIRVy1acH3PIWWgLsfXPxTtF1UEM02L1p0pLgth4qQB9fiXAV1Z
i8xt8OqqpY8ODt5+vwz5LV6I2u/4xGzJy8JNq08lVBj9qQz4euOB6tA/aX3gqur/6Jshmmk5rAlv
Z7GHGyT17fZlnkNbCZ2mfBcWM0orUDKYgvOREOBZryNFY+Z6K87uGlMOvpky/7c3RQXm/Aaqn575
4uqkOaSGZsiu5Kef+mTQsnxDnWvTIB40WJeyZKG9c3WXYcJDhv0PWp0YfawOOtvpe8mcyHtQSP2M
hrxxsCSqOjGs8n1dSm+9OMgxgmR+zY1iHQwfK8C9PZyrAn6aW0sDtLFNY2XGS0p3U3d6FL+ovJDn
2hvAu0Yjo8Ft8DlA3EXMVwpv0H1G8f84uM2qrDRyPa7sL+HTIMw5ORQHtuMBkKMBgrC+tTIbweg/
6SZ2L+QFyUwOFQCNCdEP6Zo0RQPFSoyAI+AIMtc6UFBavgEWYSLYrBZofaNSYd/f6Pu7suF/j7pf
AgRjbcNSXXOk/x5Y2k5dqs+3zlaBwMom/8v+kMsmpNUzpcLZQn24v2znyApe+gZHPh0E6FCjFCA3
+rR7i93Arsd8UhlveuIISSCxmxWUDXJ0IE6MeEV9wL9YcpaA2DrY3Yo4WfCgX9uEbQ+91RMzg7J5
yXz2+ZDGUQ7ggHOJUBsUNTTFnZ0fskbSwNeFMxqdCuHo5cxMmpjsGU7ThArRWm2+thGhGBYe5OZD
fZRGHFUjJ4Evkxgzu3iEH0MHGysxsZz+4q/4PRqR9Psnyzc+njlsJ3AURXOiDn+mXzr7zfDI+6m9
FLRloA+BWJzoKkjU2Tvt/RfFJamJmuJfiWwieAqyVkwqMaaX8QrlmvK3DaBw291/y8FAoVMjhirT
LEssW9HB8YdN6hFRWLqdPtsrKOo5sYyC1wnGHtXNENQxehh4/8cY30OglrSdX5Z2O91E77nrQgkC
D9glij0uBjc5fKXvgQvKnQii9ZZuUzWYC1w/oALb0Tzdcf0zU08BGt2FPxIFRNMLt91wnAHNncbZ
pP6udzFlJkccBN+Qchv7GT1obAJ701ycTAy7nyta6oMvD+VJXAaX6kCs4DuCt9vdkm+enTD/w2TG
Dkn6iBdE4WNZzeX27S4T/DRWsWahF7NbN8siDxLj9F2dLNdnySjnWM22BYoy4Do22N3aD/JX4DOe
sVTXvBaC1JwXMEoLqKl+MOh+1ugeeBW9ii5PhpwYzcbBNUGha2j86GNbmW1S2ftcwP3mFi5OYclC
FwHmUIK6q0nVzvPdWPMFkKeGK/6NY6t4W63cKsFSr3FlVPPSjHjVnZy+EEalegGCJTzxn4wO0nc7
0388uOszjsBR0WThkfb6xd1FJpWZN9VhDHmOaN+aIZ4bOrpvQlk+d3zaMRgJxIBpfxGc8pve44pa
9f55s3s9Tn1QjFRCGQ8LwX6qCPktmPRjDoNSvKuPKdtTCC3ZrPl/twLLe8T+FZXLdf3N23Jjsk61
DsAZuA+BdtDbI3R1+OOXG6Kfr46wgEsVAjo2ayX8WhVcOPF7DIQxoyJ4rSRFSMS/gpnjrvhGosw+
celSq+rRyfKYRIjuj/vvIWIX3HvuVhlMn5ZRoHMSY1/uHCdSPWEs4Q3QARyGbIxN8ksxXS1oj3Jw
x+oJLJr07vA3+XYAsOAOPaLvUAWNFgznXATxVy8ZP0r3llncrWTgFqqy0yE55VqJDQsCfx/AA69l
+TIO4/EY954NgBKEB/01Tx2xKN9ZkXH/MpvAqf/VMdWmis30PUD+2+8wZtc2fxJn8dqHt3avGHpW
KQlsvSf2xd4NdvYTjOi8HrqssS8/gnhEJNDUSerXCZYbtLRtFJ0TDSc9dVdyUGYdPtCJ2CreCDH/
GLipdpejDpWZ4oZqLxLGrhQ/tCSaV0rtl0670k0Inf6Zq4jyxDRGRvBTLzCe2W+hipj/NJq+ccmh
Q1gKPQHx1MtZPOCAhLTPDAhnaFVr0NBf+ytRmC/uj6Yvf0hiREJuSJfZzUSMnlnTB5iVrmitwuvZ
K8v/QjRP3sz4/hq5aeZxhX0Z7hqk5TzEr6yd3JQKcOXc+wAAt0zYA/5RtrPeJ+LW9H78EHRGQ2py
gHfg0EHDCfC+Jhn/lWLO5H0ajFUbRUvx7dHuGLc//fl60h5iWMObmEHXtfks+B901WNzpH88ry15
pAU4oEyXXe7wh3mmzPFsLr1TCDsErLZElNEFQ4GGNuaD14EDV6UO1YpN50qzrLBiqlHc12noYQGb
36NJle3DUngtP+Z5bR3qLj9yTJMBZ/qANV4HjpEkfRszgNXD3vJ8RIb+ugx1oiS9dIukDhySvTL5
bVCZlMC4uxRt4dWlS5brjqQsB3CpqdnYLGBWomzyZ3Scp1uIWoHluEYC2nlaJ1UBPH26T5O5L8aB
gClNbjeEzuFvfKjTXzJRZQiEH2KB4a+JrufQRVDF1t+HuodpCxj/XoC7b6iNie5m7NwXMVmPaUey
X1gDqJK6o+AV0zk/8c7Tb8414Gy4/kIWtAokt4+LX3raoPfjjsBiqOm7KqjpYeGnKWIlcSCJtSUG
/iQXjkG+p5O0xRQCv2DIFzHEZ/vRu/dXT0OKaxC/WSi1NN/3N9F6d8JTbTBJLmReMc9KoVS6587H
2TCrhHT6NK9DP1bCm2UNPIhcpgiQoXvqMlVRNWFQTBliSGW8NTtHnqrK4b3scUwRj1kUmcmhBE2j
sPFzCzW4djBwc15Kxh1fgRPF6JWuKSgqskfy+Y9QOZXn0sPjYuwoDtVVhyHzteGq7HVlKSjWhZri
Ev4lyjr+tDaL5iXzZ8+JiIf6PiRh9pLDg1heR6DfwSxQ+B5IQ7jCvxG3Ol98giICNn1W6uTLkJSg
lbKp2zmpDIGwKPWVfIq8yGYRwZTXTkNbme+ZiVzHlqBE9v7vfzQ9tx8qqwDFcmOpZlxTP8qH94gV
aebwmJ5/CWLVtvHbE5zSYEe4ocr07s11z2wgudxNDQ7Z/BP9j0/4mCeFbWJjTG6gPUd4ZXtRVLH8
iVQJUkM6k4/8SObtf+tytSQe86zpPpm9wqY+iO43kAOIP1FEDuef2ZTJvLQB6lYqAAj9quMth2dO
cHwpVjLPPJLjAsnzGgEP7mn4d6cjYCXPC/e5Q92sahviTpW8IPQSiIwZgxApqCigF4pYEYD5x//X
EX9v33cRtudflEw/c6H9RYskewRIOzp8ilXI1dQQg2E2U2p1xKJgwVU5WnVMzp4tL7eG+FsMjIY5
vMSLfhjqji/YpTiYKYzz6K8HVzxDYPsTsdNf3DWe8bmFKR4gCqmxvt1AJKRj8n2MhudAekhUyzLz
l+o9r1nzcAY+n8wSVG3XfBLjpH+PmlcvxJCd1hGnpS+HlXZ127SVTHYusZjjJw3BPztU7C+TNKXl
MmLYE7Z14LqNTJ3BlDZe8YzK24hDH314Tt0LxQn1BYjB/pcESOTvX0P8sLJwKb9zAvQYllHA67+4
J7F2aktpqOzPlngpB1fa1VKFQX/Im2AoFO04bFpx/iSQEBg7j14wNky2vAnRdA+1JLjZrmNA9Q0c
8j1cvUnvItx4JxZ9/KSsza+WLw8TR+wk66E3QWnyhvlUm5bgdpwEtae1IcoF5UGnDLk0ckskCPaV
I3lvyW8Wq4zrvOXohWC1tX4kYUbsDM7zgbhnTpwpLGRd389Q3BFvSQNkyPWVkYWt9a/GjWnpnoTd
L3rPm8wfdn3Ei8QOicg/yVIrGtPM/R1xRSkvYjIZKEbj0wiKkvMBF9i3GMYuMqRcPOgP3Tjow9zO
S6KdI7n6dLeECxqToKBjBx3aSFiK3nOnqhd44zOpcngDWB2mdkv0n5Igx17vE82u0HXV0vdYAe2z
KLoSoIw2pOcQSv96Qi/7FtZR/+t/MJd6XWk9uhwRbCEOML3LydH5N73fM+kFU++ZHrT/vDOD1Siy
EkzCWsz85H9fIilK3GIacWRmdlwZfZ9uv0cihgBsKiaGNkcdlcBWVi/DErXFcvOvxfYVkm+1UOs4
DPTF2Ylwv4QZfcFfSe16tT5OQKZijatmufkZaCwhjY/UhPTKlkXI8A4amaAbNEzDHYOu5zOdGLlB
A9iWAJRo/kqNqWoh4huJdOkvSI+4KRQ/YpRCX5UqD2sUmCVTjXzCPe5IAvQ/soX+f+6a9BnI32gW
sC2kqJZpKiXgUyLrRKHL9qfIg6h8esOoC0GnJSWE4P9tWqWivhIi4m80r5lKbHihi6SgUrnkVIaf
4Viv2GKPBi6+JFcBz/iHuYUx9klGJRSO3kXCjwu7ZxddHW/gKDwUaDdpkNK38/IzFncRBS2BQIal
k/UFJaaK9lL52KB/Tc/qVNHKCH4jaI6JFiK5tQwuptGhHAxBLDmq/g/zVSCM0m2fdOqy8NKParD5
ahL9u/48cqLbbqVVXvwx3xqtRCIJ8X2J1UhgJ89GPZt5faRx/GgppwZYG/iGmldlG/EjndCi9nDU
1kKk2ZMQv5xE0IhZiEvLILpS18ffWRK71iy6OP1CBefFlLB+9kwKq5TVCFH3Y+pLK+wKUrmw8ECJ
8sH8ESxBvjkeraMgO65Cd1qt1Ab7vZjvtwscwQio/8edJHZJO8g0ItyIN66gPLIX5xFGxyw4kQA0
sZLOr/JX+mWL5DL3FpUYfBoxtjC/JyBh7q6KYE+hmAUPbdE50Er3YZDMcie5EqxG8MOOKXadPK0A
x1mWpaIiFR1gDWgJmVQjoTLKbLTfH5TN0APQ+srArgm1AH/DR8lv/Pjts87+0gUjAX/u2ZfK8mq2
/gWPVuRncTPngZCgT8QGcRXiMWOR+B5OiMndz55lEIqHZEtEQDoZebZR9DR7OcY1k87FOGY3JVkx
a1X9v0+omQIQj2o5jEHquWBZqdk2Ig40R3V991MvpF3s/TPk6FZaq6y0Aq3EFbVw9Dmvq4CBtnd+
afmDrVDEXzWKg6nZ8r9rsli9KWVZROPkcEleUAV61pYvYa+9NrrNgc5cwnWSNbtE906qqhSweFQI
5rvrp7gxxXYKKanLySyftg4fDqAjapk2JSFfX918AKVmqp9zS+JbFkVAzKt/h+RzPEwGm+u2QH9z
au6WRXa4Hgv1M9tkf9ZL1xgHmByI1ZJalmAXdSSenc8JTKNpqA+zXfjNd7HN8lq2bkvPLLSjKdUx
3AG/B/8eIorOZz3t18EiWqoqghwXyj6Ew2S9OPQGbuXbA4M00cWUJbChfSxSUH+ckZdGMFcwyshP
Xjk6EIzWwQVAyw1ZS6kZkX7wBBelFlSfBTk4ki6/Kpn8gZK4+92fMkHv0cjPcwpLvI77XL+MMR0p
epK81YZCxeGlVxEWZgtKA8KanEsOuI/Mf2IatsRaGKt5GB0R2n8LoAxxL2iPJgNMBHtt4uJW3dFg
FyDm6HevxU71JV/dfkc8qVD4eR7iCwzOBs2hXM85tf5lCqvYU0RgH3NxHkUXqzSYmAyN0wDzU25j
7pX2250nSr70op8/jrk01FVXRc2l4qXnghh8h9UCmqOhwa3lQuHxEy5SLpfc0pctD32NmnhhFVX+
1sudw0TuKTIUhevoN2xZvvilO4+bSas2yITjbEVAWyyWGkmQ49rQpz6V9WFHAegpt17IWLARKNkD
vxHdDpKwmjzGRWjnREXr8nFmVWhfxDtA7RhY+HATRlNBDVVbnjvcO/sEctmrvVB/6uPV+2uhVDJI
mWOgFo4m8v24Iq6SxPek595unvRulynFzQI1upy1fDab/J7gEH2sxi1R1rZ1KF9SQ3EUi+6VFUs3
QbD4qypXF+a1kH/JwKkRiJKaQShFhUHD2F1Qdhsz4cq0j/tgilfkayNUcivc24NtbNGYWCV8zyJz
kknk/wGuZereiTYxUuASIog6GE5oGENdKZJd9PtUzMzysYA5e9bAW6S3dPJ02lPeHYevg16DEc4s
udiNw2ZgtFR3u9u72QA2gvvJnZAWg3tVn3lrRok7RE5JPfdlCpx4IpOO3gJIeNiBJla1JKIOmnu7
jssZtoCMs4qoPb5eNegdXIeWTiNubeHp0YE9E/AT5UThyHhUpBEmwHkxURIEucMlVsbPOI714sqs
6WZZxx5KUQI15oKdJ5YTpLTv69FOLK//CGpuown8U+fsVCe4aLfFF1ZL0liGeRheD8upY4KNHoFn
dHL1rI2lQy09EwpA48MjY6ABLREbB+xkuuPKIq6nTVYr6msyC0ylxGVrYl77vxImL7OT2X+gOB9b
TmKPdgAAQjTTRhEuwah693VdowhtKBkX7nRVoRR6EsvJCjEdATOcNbGi8AkBsvPf5mx0yYiwQ/Kj
J8HI/Q4vtFA5RIjBk6s6dO0AujXh1ruUSIMNVd55ahxpvS/Wo6w4e/rV9aH2+Cxo+LBGqxfb3NOU
vQQ5RBIPrKuNQ7ESiYt/5PPAuvYFuBv2K8eH5POIBHaTd+b2ubYFazx5RC6Qsd1TZ1vhyuUMSyxc
tyiCe9KV04iyaCq/ddjht/PkWkxjqYSQmfchlQe32EvKLxNlXCzqABq44Dop4Eiv3sV02KUqi8mV
lljZ0CJz/hu4ZhYx/kYek0KwkCC5fgaiGO0dJMWtTOVfMaf0PCTZ31Z6bB3xQBkaMSZzyXir6Pnf
nCwmM3wLL+IV/+QdSfGLGFqnRAZmTe83Vq/CM4nhlwHmhEFUD28GJjiI8arrbs5U8AEefaIwGk1r
tsjD8t7WB+xqebTMXjEfS0TJWKnEFzJ+zxxfGQwFGkqMk2CHhKnuREHsUJPruNHjLTnxqbnxv63l
+c6adROL1eYAUwIQJ1hHyFmBn5Zm06ekFWk4LeAQGfwpFLy254njqouwyeo9T/4vkbpkHmLEcYJ6
zF2R1IdH3DL08XZ16iwFltTcRn8yrKWo/5AUQsRTquGR/PugwcpkVu5ydayhGytySD+b3L1EqKBG
rNyITe4vSHUqweodnc6g2zbbzDxr8B0zJBnCUQM01y5Awhp73HTXjMDCc9rQOVwfFpIRYrN2XSBC
r/yBX64ILfCfhbWKFH0g/yBBldHGWD7xql6+QTthjx5ojRwhgMT4AQLRafWNM0qGoinD4I+mh8/X
X0j7gup30XaIoo5vCoUYUshZ+FIUISO8VEpnViQG+DtPpFrfNJklFpa0iYcQGuD4xMAu0D9B8qCR
uGmz70QBf7ag5WowQTcyVKl6n2Uz/JSKXvprNv2Ie9lLkoY7mUuDdoMz2LKWmCz7+qoFk4IBMIhk
F5oPq8EeFf+fc8UyRPrroS+aM74P3/137eYFohCNTMJ1dnSe5IZ0gIagr53MvbStU4d411UUnxDR
rkAn7XB908l5KbMltcfTl98ZS2ooPTxkE4V1cKbXS6yOC1rbt1yzYzrTH+wYKICMmaqy0Pqst1wN
GWzxp8uAFpQHKOfsnAHIzVmJgyBUzo6GcU5qgcI7YYItoiFvjMfpbFq14ktvcHYZEu28lZXfCt3t
mFfjQCpSH+IH1MyR8Ym7gumJHug6GZnw51GPWi6NcW419+PaPTTvI3+/Ty0i0NOS/ggtd8Hpv+s9
YYqf2qZyG6fCAcguo9gOgMsILICmmPeuGtXxWNhRJQSmNW9XZOOJNF4Lk/0CSqaBeUcEnnJAJZOr
kNKyhxAnDgpVulnE8cJDF5uE6uEzZGs7Tf9NpynxCdnRMefFbK6Vaa3RShLIlN9xxBNiKGL1llbZ
Uc/YfXnC8ytCAOnF1CrfTYDJREpa5aodb5YB/E99ZOEx74/IHIzQPvR1OUlX2zfNzAkTDm3k71rk
o4XoZXuSFbsG2FZliHKHFdsgI0+dP0flWEe7zHUwjmcpZ2idkNTFXltZNttaQz3nV130cxjzSBRX
e7b75/jKBToDjmfRfNr0JQM5wbuGQfbGiJCpTlpHAiwNVc+xZ0W2DJRFgY4CmLGoNEseiR1yAJZi
dmBKNwbZwQ8SpqzcnDEGV/2tCpIEw024mWGqnL2JSBLNf9gTQsQ7fseImO8oO005X1+G02sNT+m2
82uzHLD9OADTm9h5lD1ewRwRlfZkOihzePznInfB80Qy6PW6v3m94TfItV82vVSpagHa/I6yr/bb
V67aRL+TSBiF6zvSJ7pEGOI2JqBLwdRsbduSMEat3/cOs5fWm2zD1fToHs3PtBZRrg+Q53FZmjqK
DR5tJzR24sgAeZdPbLKSb1Om87CIEWCZSa7qqV1ENHzbLhmdHl4ahzY3OwpEGbH88iY+5Id8yZYO
YtCRrQmAYgxqozKoQcNYeQKD+ZoE7Ahnran08qMTRhiDjwBxD7BkEzrBJw58UYO6hWv5OEVIgpfm
fWN6XAtMpTL2N3HuCo2jMK04gYvx3+yXlzEpsIYYy4D3Z2qkEhAlrPA7OaX+RqWHYR+azQR+T9uI
TLWC/wpnC3/fqVBPSDgGh6GICw2i+zrqybYTnosTZ8Ha+5Nzm67n8sL3B5qyMV2tGahqg24PzDbz
IgfznXT/6HRu4kEN1kSNuWIM2rgW4rXfX0dXPEwpe2AgyL9Ej2yYKj5ByMty15dUbsUwIHfZzq2c
U/s1axt7Hk2IJZZSEoQDccRJwPg08SZhzlaMfx5NyAOZlSUjdDYAoe6/YSxhTySFDmn/UPI72mGu
uXGcIUu3E3byQvin9fc02TPEAGfiTQC3tmnzvtc6V3JpZ2kiBtjGpkWQne7Pi1oCLcinJ8gRt3qq
x9dY4Cjs+FNEelPpJeKfFVN1eRhoAqNDlekTNfv0Gkq61Y2ZqwYE62Z0X2qOKHvp+1mf8qki4/4Q
TB2NkWm0PBy9/paEyi8PwfoFg5js7Pwwqn9UZcOmEqBeP04aYCVoEbUxyJvhXnv1Cf3stL1SUW2L
9dcr9JN3CYGM9rJ6bMLYTLsz1K3kCK0WlNmK7kXsW/A025iyyx0i5Frh/CzMSkbNb4XZG4lW94mI
frSwzDfpgogskweFI8rJtqrNBxOFBzAUHxrgJnEgXhjCOV8PAjuZhCDQiNQ27Exm5gIfVoXK1FcE
G+L47wRRnAAcTCWUcXr660li8OuK35TMiyFHjrfMqH/FGPTu+9kVXTlyqvK9SGxQ8FiS0j01jM11
blU9xzpYbM3kfvXkvbKzQB3LIUtKWN7J8Pdzgc77A5WsqTyjSTizpVKc6FHcQ9M6mLZ380Hb726e
UJv1qCGZwU5JO23Fr7cmUX0WMwCU4kUctCal7taOt9xjAvHQLCGhSqJhKsVwe8C9eWI/vHm/oFa9
nLlP4Ov9vTNp6FsLfRPF/93tHNcXrHyH1IMfApLIFRgT+AJGGOpUjoIUDq0Gw6VpNkEX+xNJi9+R
bvHUkgk2aNtSeh4pQL0nuDzrikbcwKJkRTbdMxI42kjlN5xJSJbjp2VU/oSQaqaUpfr5wCLHWinJ
IinCRQSuLpY5sTAzfsvvVIl65O8Weqj5ioS6YQ6uqFkQ/ycvltTIBWBxCsFmxm+yXqRZ4bOrbBcQ
3AmUQbmYm61zb4HDx7GDBPuzoUzwuRh7fPqgIo4U4W+IoH+263P+N/+Ks8PWOPD6Tk5py/KlJI7O
zl7jQzRM4v0O4WpD1F/L3+NxO5YVyGEUI+3lC4ASHC5jvZWtiLTmkMHyh7D8oi/bFblEN/Uf/6xB
UiLyggsOwX0PJPOtYmIArzw9q6cm904Yk8BnuTH+BTIMrpixm9ux64fiWprSe2/4eDDBC3xX2j2a
w6TWOxd0XI0SI/edL7BC3xFPaYh8kTXKWI16jwm181XI697GLB/HNFk+DL1jh4kRI5mTdZa1FqZW
fZN9SL3a36aqaZPpcv9zSVZn1VlTLEPC+loNXwNSV7085jBSor3RHLTwy5AYXfoYvXPczc1fELCW
UME+BDgaVp9u43HNrXyY3OFU4zb53MK7UPAXvtYMO+Kw2MQU7bsieS4Z+R+NIEXInPwmpo9bZRfj
kXowSBR/QOdCLr0HTBx4UjkMlsuyD2CsWoTQBXIB+jPBccAo9naSWvJfmig2Xid9Ot2hyeoBjYqP
sVELl5QehGcmH3XtMoTBqUZAgPFYnbVxl1rZmwgc4SHBs4Wf2S0fCH0aHsA8SCl2OCBtjwIi3kis
YCo7Gy9Pq99pCa3sE2fqyOuopH+pKRcRWdIyHgCrgN49E4TKe15mf0lBXMO0pQO1rOVajqGuOtEL
CowpOAX7BQX/sqEDjSPxHHh0Le70LyY/y6cnk355p09BH11rWeAQK/vzZCtRElCLDWCzxc1qEQSL
i9VqX/6sPV20DI7ULMPpTAIm6DvIrE/DuHJgdhqNSyTogf94iZkDkEsspdY53i9qmwzrCoL9EQ9x
Sat5IRCNWdF6J9jO6LQJuL72iGAxCXrbI/PR3SvWZteD5Iu9vvmE5gxlsQhG9WB7R4IEaZdVUU6t
PJnUj8wkWBpgJRMOTvWn8wGlu2Z89rhBgl4hoPL4t2WChFsk0NmPvAC6+YeGd4gg8D7i0kTHwOho
IBRFg7LaDI+8VTc8dO4luYaJNJSKd7w6dPFRrSBujlN9eAX2EV0xx/60HYPkoGvC3bsOf6kC6yXD
Dv1fffWxBZRlKO3IrHWgw0P+7XTT9oOBTCaZa7YIKj851pybs+aBXzk6JOOo65lT0LHVxafwyx/j
npOPIRGPVi9lISSiFnmjyC32Ys2nmWHyMfEgLbbqbbKsDjOXZ+XgMFYlj/+hZp+sIb9iRx5NOCyN
6lfr/v8WLV3p3saDjQrv8hHqcYGbRm6smr5Krc5Uyl0BtlrWMIQuwg86A7IRe357b/P3/li8HkSP
JMIXjpSffLwcDaWJU3Ot9ADFQXl5raUheieczTrLJHlfz98XX4M2+xn9VnoH/y0kcSNzNYFjs1DR
/RERKHvOhXhBK0Qf1Q7JWuKtJ58IabSC17WAsLPDRG6+7TYXoSCkqH9VH26/biGtfp8o0+aTPe7F
DffUhVnmv5qoP529PcutTQNw99cQf0XOv42fzQZLgVKRAEkVCxNaU9z+BuLdypIAYGPbi58GiuHL
duH5F2xg9LmivgwsS0khC+18KFwTSBinWocIc35t1kFI66G1Op1gCrrX0B/umYGYtSs0ox84L23S
pt+qJc2+NMo7JCEgGC6IYEhMXhchNN6v3FTzywJDt3CL+q2vcs1qT9DMCZfrGvt34UlqAwzdwBEX
XwUVzQ0c2XXNcufW0J9B1WbKQ+gcU3LbQjgpwbltaaT4GAOFyBrWLk6Kk8k2YY2ayDDS5XxRlNXe
Fwe3VsFWezKNM2HtnjaCZcPSaLTCExwfpLZSdtolcNu52JmhG6vyndfNHhogPkMz2B5BbskZBEvb
GzQecNRQXeWox6CSHegWk4xC43ezLxQ1ctf6qWn5/R87Xtfi3tL/m18T4s+oW9xeLNSrYIIGaeKE
VINcMKMTvvSLy34UrRFPnJdMTHXOgDBzIFyCOC3bDDH5kiRnXnRZLWopAe2srzsHlHzOKgA8cJe5
LdwvKjibm/4ykm0FDxR7ijht5KanSgpM/EVKyL8Al1+OA9RPhXbOBrlxWlNxszYGDP3+V8GoAYDM
nRQI/AtNEBAl0KLI7F9nLdAN1TF3SXOuJ50+KZml5IysCmJGbEBOGTVwmBG9ONftOThXzxQsvflv
60g64gtPneSZLe/b/+6zFHyCyxZBqt2l4oFdG6JRcUrcpjaTC+ysCvQQgwpWXTyAwkMqcX52z//H
4r2K34RhRBnNHbM7kkLPCcT8E3mPJhHnFozMdP6kNKFqc0vQOp898e8wBM/vMqRuobjZX0dMv974
ViMHb6AJRhPrZ5rooP0srvdwZl+pUuFmPoG06pRSbpJRGwdMhmweSTFBfE+Dd8KrxR5K7mySuMqW
raaFQml7Q2LKdsRqcCQY+iniLhensusb1kiOMjK7T/5621nJ8k+olcOI+XQJkcDUsKmuZcxVgXtu
KDMzr5K0D2xP6fRQ70Rz9xOKCb1F3KIeSREj8HiglbccBswPcLvgj7A8u04GvBv21VSWSuKb1HmL
MWiIioIHn248sTi0DFBrBpfglgsYEl3t8NCOYENzXpk9nVxPFlRJquiA8CXS9oKQo2Ji1LNLqogQ
NjEcFTu2yRWmhx6bqarFJi0NWXd5wGCKc83nsmDEg5zMED6iSf4l4pzX3/9anQgZ663iegfWU7h5
GkZ7p+UVFRfikZXUf5Sr3R1QLjxpAErOQo4usA5v2apmjwF6mfrVbdr3MOZGvZeI32Hl6lorydKx
+dd5Q8vdN1JFQnOiVj99m95KS6AggJRx/1xgET6zKJMiyd5zpZneWRGSHwFaZ1/JI5teVYFU8qTY
L/xWkOMGASl23VZK6+0yZGEUsxBahZg81Qbpv1IAVGMEXNCZOdFlp1QVzPzQB6VXCKSZviz9OKXy
eaSqjMws5Wto5azRWVh3qj8dlkG5woxG+Mc8VKW0yg4NxnjfwzucDqunGrMUXFjkWx00zu1N3inz
1FkIXAl+WPplRUFWleNGDcAp3oDayTpoWfKO4OKmUpZGQZg4Tqcuzbycnicd+MUgvcXqf84fS9wf
Ssk3qh+W8uCDYPn1hGDrIh1GTHKqnSN1z/E+3jtJA1oNxaCbww0YeoCa/J5Ls/gc4jEUcvTykLGp
uTPpcWLFxbutMlkUqTgEnHNpBwEufG/UJhRtm8h36+wbU+jUBMxYkGCbemhTjCma9gYMQsagp1sA
pcvJcMemjCvEYLoe0v/DgYM3fDsgqxX939vX16EZI+UIyBn3Pjo0iGnzXx5fcErY7cArlYNNR486
o1CVGa7jTsnvSsjs1ZABpQ7pLK7OxQeY+PQq7QTwQLgS1vmAHVDRV6unKGPHCPSwTXuZjegSqaQF
7s/lAGGcV/8pUNQjDGuwFd0GfidA4toulFF42Tv/FfauZWGfrvx3s5wG290fLmBcUbyE4vDhEk7O
Di18iCbQx/9iu5DR/EfWp+YYaSqfxhxI7Tv/DxnLjAOYLFoPIHvZVBnp+JixzWhyNMes1hTlpFgB
VgWAzwX4R2a7hf3Dd0gdrnGVWAVA0QvBiJu/cG35KhpV5uLNf3Xnwejx0Z6fLDVMv9SwxYs0kYPA
HJnhhJXL2hburbPdBB+vpEHa/mypwQXgNQbRL2hSaTLvdCjJrUUHxLgX8oLfzZUl9kte1WcwuCFy
r6xH8zGthApqpxrAh0xQMwMGr5WTu03DGj0pb7a2qv/A9yz/OMdwNEPdaJZGf4mqJZzUUDqz1O+P
KkPP2sND9XHT1cqRSi2EQewNPV78sFP4AXQ1BYho3CrGR/t2abSCQ0wk+r8QWBLb4qxuCGMo49wI
LyhHeXB1VzHSP8ehi17A5RFM1o3Ut82jjAPHIyFXOySlriKWiQ8Mly1e7JgWgYPNwegvrboMfmhx
XFoKqWTujvBBNElZ8gVVF0bTlHEZjXtxo5ES73F8tYYKZV/NTSVV4rmxllxKjLFu69Ro6VFnKly0
1B8/OTvfczn0ty4rUvgOGxp4lWL+IcGwkUcfKnf38kscz4W9eCY1UnON82CLtLu6MbEwixi+Bc6o
MXl/F+Wa6l1pMS3weMfQtG3zgcFj1IzoCf1meTGWFQhymWgFgZxcq/m3zDIAyX2cBIr0Fh39KnsA
Hu2lknd9md35SlIdk6AXHBubCuzRtkI3pCq3v9ftuyr1gzje+e6xfSve082Sgu7b1aSNZIInDThF
brzVDrD6ZFb8yhJkLs1T8cWT/J+fnbj6tOesfFu68pXDoCXNj2Xqo9H3iEdiX8zOwJ3GshYdHOuq
j/U0UumptlATF8R2rwWnlD+m3xih4WUcnpH8UNwmSyy6W/GIivjvN28tc4LQqn6DAocJnYkN6nzR
7efpjHFEGxx7jLG4HBz/nHYi1jhDnEd46fAi+86Zpsiyu6i8pjHE476IwRQ6KS4bG6gJUb2PdZIo
cYNrX94hHQiuqWEqoIpGNGhNHZ6jfz7dPngc9aZXJuweeG/EPXGsHUePdetcGGJGck/Rx3zsJMwA
CFSK3bnQ+u16socxcIXjuEQapOD0+5AsNV4wMiXUDpzecaYsAFpTfiplpuerbHFbZIBSNnqBBsC+
2WVsrQrsOStvdPyeWe/ZeXNctSjQqCjr38BqJbAusZ5gHc/tqe/qvUlcyNFDGywQ9hEEfrzQ12Xx
tzXknNtLx9iw0vZD7+onyIy+boUpXBeY/whAIoL0HvmT0SnpPE5LyMsHMI4GH5KRr/rlC70aBiJ5
6iRwCNh9fwMbmSuQkA12Blou4DtwK/mdffVS81EgxIQkSzgR2fcYSHA/0Xcnfju4CFd1f7fSufXA
dr0pvNM9tYwPvQS/SKlvD3JbEVG3canNicwUAw5b7dS9lhxjSqutYJbMT6cydg74aYuTSHABGE98
//lrV+Ep0FVle3HOXjxNR9DPXwKzSVOObRyaEM1EKrN/9PpENloZO1i7bERjlMxSUmteIRfcyC+X
HD1VbUKSFj0pDTi1MbEkyovuRl+6LF4NZNP4H2vUq908xbFYwoz2RxSqpZrtbkbV2r9XG90tnUYQ
lT4FYdgX2RTBiPX6ugseW0RlosR1rNwMeS96d+/HiIWSxUAkyvUai4uYsRk+6JJPDCXtlHypjKMI
RSg4EtRl8Gd2AiB0oqeubDv2Aeqf5BLQ+sVlzQFwDGNw1NsyTK18nzdbVzXfWnOnFLO5YzCdOzTN
lDsr3cuhCzBEf0zHaSlppRKNTXv8+iF2bBBCJ2KG12yCLyMCzI3/pCWBy6Ax9yEwauSyWjgdr0W+
g6GbSo4hdiDWj2DexcXsVKqvgmeHelf9GpXTDxBKzaE+BH7W3xQKIRfl6xUw3Ue76kHWAtr18yHY
X0oOyZ0849QYbUzXWaydF2Wa3qPgFUlxFsKuc7w5+Z76SJPtBf7frAIy6dSyIlJaCqAdg0X4Utum
+1285BvL4C+5kHj4NIV1iMFzpFuKl53lyZDE0RTJua2emlRFmhnYu9X0kgIuOwP6t74Attd3Vogn
w8mJOOXJWVZfz8eUBnkVI4g4a11gHCCNnJ4AIn+wyjd8GYIwoZMpIcW/YBIhmafRw448ecVwSBjj
DF1gIzXXQ7s7rwpKlGidgSC6ZOI+I+uV1KzRKqc5p+PAsihqALicZPjWMfMIVYdBVX2K7jyyZNXx
sB9VU8paPVU6Uk8EDxOa+lC0cJTA7ccKE9NNM5dyBspsnM/J4IFcISo5LKnx1qm/3uL4kozaVY4J
apqg+tNDfBl7mZUIy6S9FQkrMWlPYcufc5FBoOSrZcxn2KH9z/QJETqgDaDQKd54HHaCN6AK4IS3
tSO46vfnKqpms4p32xem6NS2L9TZ4Aiha0CQG5dJQ70SD7q9rWZW+ml/2wOpNMa5nYqOMS3GIRmS
WDipvvv3pGx7bE8quOqGrfgWN1I3iwHMt+0jXO38EfQlCvauIWGLfgGCz7QYrbz9KMHMW431f6tz
BQt2cCJkhf1njIwKaeAv1/CHsiOAbGj+WO3GRkJyDvSuWkBHCMP58Hc6Ql5+SWDjLcnE9mAgxbmH
qI11KDv5N6LcCEtMZaQuqM9dHsqbHwwctoIgycEQHhp0VHhpEkNuKdC1jnrlfiUaqHMGzX3ivsx7
XVQQ7QrYBp5AHtNOKMNYkGOy61uzCDMdJq1mpMbuCbyVREEMpXgssF/7PbgQAhQtJSB9G3rV08S6
bggaoEailvVrF/hYdSCULMvsMtK/0hzuxayPg6zl230RbQWPp1IsWvogXJcSSItjexsU6EpxPNaq
7Ie735wXW6dsuz6BUviWu7gJWo9A6MMf9pTOVh36SOkK0go4Pk92+nOZiJWWUyYpmvjGcetis6rf
wzz/ayvjrvOG2l14CHlRq1spsfx8TFjT+zi4rsqMMa/zpwEtjyMbwEc1IH8oFMow930zvJZUweaZ
faGcgtxR5hdPIXxAbUoA8cc3/i/47TN/7mbVVjACtIeqEVXhME2z0TkWgBoV8zkO4WS/KKDzPql9
XBq/VhC6Qul0XGxvBTwapTtvMbKWBsaEZfCPrnRHKoEJbVjMV3My+vPf5uv4d3oQQoyENhYVMry8
P9RI/8/+KZJIhk5QPv1Wj9K+FCY9T4ZKGHCop2yXmCbdUJEClxzLwpSzlZoADmOiVlXD7cMv2dCl
WpGRGTfLQRjyQgigwqeOr65X4+67RwXFwn9ZuiaXBNlHoPqqj5GPtTHCiBPvRCWr/Bje2mgSkhHG
9vse3TXGvAl/HdZVMmY+1p/hfaLEojhxNSt/LCs5XhIuCfCnxsD4ChDvoC+7YleuMyqXhjQRUhPG
CBM4b4PWEl+Ukq3XKWPeb/VTD8O/qOwa8aktACmMoq9FA2KqwSHdQPc7+YtOMGPwNgiC5RuKLojP
e53Q/IzzdV3lBOzNGo96wvnturPtdybIPV2d73KIDPoHMRFpzvMcy2/GDjEgI37PudYSPJGDe8DU
wkCC7I+m9DIcnBMp5wZXzfyysGcdXNsnx0q7Hr0uN7LCAFK3YseDsOhS2QOyCmBpFqSTdxVv3myK
kbcZwrCmIOr87+GgSdfLExvpt74Gyzr1WAtXXygf71GclzR2yfpXl0kAhDheAZ5rYkzp3biM4ceW
UzYjRY+tKYDlQy5rq+OLg/jImy1LspqWXVDZFJx70SPjIKSI+n5J1QD0g2smMc9m2qrmxAdVFrcl
dhmQFUOZgANnejcL3NO0+HWdvEZMs7Qg9iwdidaGP8OorM3h3crrQJ5AoT8J7N8aenfl77jNEOEu
BqZJnCy5W4GVej82u1yqqG53Lojq76t9/J9idwj2fuXbvadWStAR99zhZbJoglNUGxgOYDkaB77A
PUs5NAa+5Z4h8FuRDq0g+iwI6F0t7JjO73i1ycnCKDg0lxQiSbRQNUzPIju73sg7NaHEjzhpfo+m
7rnR7p2yWN2zUCvS3Rj4ZGiQSI91ERWILdRjK35pSIiMQO5xpYfGwyfl+kkBOP55s57156S1w9j5
1RfqGCSCFaB1Uz9DcbLBPP8wsevo9eSl3mUL8S0dn9Gmn4MmXzAslQY1gAxRib7PnEr2HSca1pzv
/OUBlVB7z0L1IYB8QfscUYZNIqVI2uFsvG+zIxqFUZ2w8pGNkCQlgqDNFqW602QP8ILJ2P/brmBv
t4Df3uPg1OTyl14l37oM0PW33zbuDeAZm1a1bMPUoiW3MNcOhKIJv/APz/wzgyK8FM8duesCixDd
DXc9fe/Pc2FH0GL0imWmcvzuE7pxY2c8wYucRSr3l4lo0bIR6CH14Oa3H+3oBiVF1waADD9K5q58
YSFhet/H36xpoiw3Ug47I3BUaqxXEfPB43lbUMGcg94qVvdaybhqoZfq64U+znOrxuOBa7DgEqhf
9sqFFDyFoslAfGJYT1LNbfHXUZJtnvcK6N4GNs8UEH9UCBTVCuVxViTNDlTXeVMUDhitLxZCAYGy
Ko5UA3/jIs0YqzZ70pGqgWwgL8qUKHNp/M25kyYZ9rNZNdM6qwOPkKNtM8Z9P1qIptwvhlb7jlMh
vQM1DSJmM4XmU5iC5AFj9K6WT49piF9NAeHhKbZ2Wm5yDqBvL17nXKBkkSDvz3N6UdwT8WNf/W3x
uBqDvsy6ono1+kLdieH7TlLwupq+wqqCvdCqjQgsoYfCJxD2dfq0m9tZk62HOtQLPer+dh3K4ot0
WEzUhiz0X0tpqRqwkeAwb0WYYTko7nJYLiacvLo3F9hKRRqSqxxMYuMHiPIMrVHPZMLnzkMsISAl
YB6rohVlX4nawwKQvAN4XRfLsIFNzKNtKTthmAKCWxO2LEupnUN++N3n2+b7hxk90fCVPDpgDPWh
5QXGwogp71gxNx/yHbwIQ+gRedn/+pC6YvjOnflwoiUJE7WMe4fV/fg5tRMH+Akbvc2aleDN/7my
plqTg8fKVSiCjzbVFehWACU+jzF/KTx99FtIg/a0ie2kXLhVcr+HihqCqNWF4zLBk3+x7hkTabmm
iLlC0Wx7Ux6BBER2GUcLv1edNES1POY21VeOkFDM9cZW1787yVquz5cA1YOpKNhQ08flw1kkcBDc
RleJ7C+LwUvy30XLoYbrcgJZ2sX+2atX0FXd9rz6U3Kf7xHUDc2AB9VMWaZiAhS3xXTh9UJ53Vlr
m5oXmnjeHzBjCyWF0UkBgVm380G5U3qi9UiBU+ZQr134zB1iCNZyqvHNd7RQZYR3k4YDETtmhKK1
0m8BAnozI6Joav6PjkVSrcUxUykPz4A8bsrnQNozWibbwl6eHNdvFCLKBEFaHac/WD/WijJoDioo
PFM5yJK7etazocqH/p9TXsIyRPeHK4FOsBcXV/yUob9GsgpKTJ9xLrisSBJqYfCSjQ4WUWAY2ma2
I6LaWNqDRQbi+8bumNFVVR3AFabJ/JdZVxfq9cJ383zF7hjVCLKvp67a1wobRQRCnwBg7Scg5n9N
69VDjcOahtCT035BvSdj3aO9+N6Q3JSa2hIiQYsVVhS2pp+Uo2oaxlsFCcxsUqzAWsHqu7fmhVHJ
5WamIZuhuc1XRDdSa3LjVu+tzXs4dk0arWAchkL5ljD1pIp3idjCpY78i6FuSamM2pBUlgj3535C
+3//GJr/5I4AS5h+12OeYagQNiOUIgu84jLv94hD1psMJJyaffClgfJ1AFIpNLF7ZG+F32Bfe0YT
7fStKktIsByB7nMDDz2VSi897XADUaRpQ7/mol73p1/08c8UKvOE6tlkio/Ywcg0YP7FnmO+elri
cXr+KpgWYGzJcwajhZ3rNRMl/R5waHF7MVBvBGeTOyW+GWNPsT9lnafJIkecqQSYxoWk3He/bgQ8
aKzht5pUyEOHLNhqmEd803PDF2Gz/E8GbrTzVkgkfmpZKBuV075Yo0APRdIrN75QFHo38cVAiF27
wLLWgfFNljttKiZqAcs+WR9UMEJo5TbueBYM1t0NppHT9FNm7EVu4Z5RZ+9TPTnL4121F+DmcJ8g
JTL4pvac0zbMzJZvm2iPi79cwL31kUT1pxy4DI6ZP0b+FwyasRQTXL/f3gX3H/8b7XBm1iF5Tjj+
AaosVlOAv5ooAfVAsDj0Dmq1/opapRZhL2hot40yGuPg0z3CksWBM2HTFIpTHeptgZy2liW1oqtQ
ev38qiW3h/NaRMMwP5O/rZ6kN7gH4Yw6IKq1IwLr00zKAVkfXpYMGlPzQn/w8KK6ocNSoesSpt4Q
+kd4zgJrjMGx8iZrQZmcRM72a93ygndsI3DFlrE5wIYc3MCRT3D6dr6wa9Nc2ed3xj1Ea9f1Fnfx
El3mm7ZVIVIZUZk9501jJxADuxPGDVdHF5tHPJokgt28/zjm87GBt29G/zg956ZiF/dLCQHOvyLi
DJgL5yU/Ab5l9j4N4BNE/wsA2DHG74Ji4LaSHzNJoXdN5xO8ZJ68Tyv9OgkNiDcFmWpY1jUnN8vJ
+g/nTt8vAf+PeAnc1L0KTmrHwxHIRc4vvo9sPwwlBlxnRC/utR16mD9s7jNdeVsXgMoqjnI87epP
juiklP3RyC8iutNfSxPGn9LQMylklXhuH95Sn6KE6ghF9zYzq71D7D1J3k5IKiOz67/nSAV+V/V4
I539OJVEeUgxaLQNnf0O3NolQaZkNrqZ8Twebkb2mNpu0PvKtZ/IAh1KkbEsK1qtek/doXNJNSKT
JumcEOfLOEFbSOZsWyS2Z5uPBdRvkFiWe3/nPiwTF7V1JzGt54K9Qc+1ZPKqaBGWZceNAkWWwZjA
S3KinvmeNLz8Rp9h4WV4lNlOM8lzGd9GECvzhnqvgnXOb8ex/Pn465GVZ55oDz8vybjcrZWpQtKS
p4lLarcwPxmhaIJYgwfhZwoivu+Qkj9FPiwxQvvYJhtsGpDkinu+j/e01Ay3fw5hfJVWEJlF6UGU
HB7bu5ELugVbSVJqL+0hBWp2oZ/qoXGlUffVk8WHZmSJdkoUu7SGOHandpnTAmjWs7zV7iw4kS8R
TYS4AIw5I0rppUvhFAZ8iuAOYaXUoW/M5bPbxU4FoE3ODJdBiHabexmI/I3R1h8jS0wAxXxf1iqu
vAp1URPO7h7BUV8PdMP3hrRmprbEwgm4/YRlpoemZzyxJSQ502K67G9hcY9802+GMu2vDD/PbHyP
2NaWDBkQKO7OvwFz7E8rziHaEsnyI0+VCR+lag8KAzbwBNgcAOAPsX/Bzzsipb46GJl8u0ZRSb+G
bbTJg0yPDpZy/fBBOkiVANfF5w2DSjNaElhy33GgirOGYAReX1K2+lppKh00IYxNpEO4BX5VdO/Q
Zo5Hb3DM5A7qV/4R+qXaZ01KFMrt20qybk9AN0qAtcndQNT7YoMuI+R+M9ctnFPhAOUAaLdbkMX3
xAQuTCzFM7ZwJN685zkcSBH5gJrtQrwJ1bvW5rnp1EoAqeukkE1WgCN5NelYsD0U8oHxJNFRbz8+
IS/PYO/mILjzTtC6+j8I4Qr1oNXxr9zH/yAImegWFr0hF1NUcwEzLR7DyHfq38PgM9L4JBS83iUv
y5CGa3UBbj6HU0Eb3uqBdCsyCzbwKIsnjQ8H/kjAYTmVyW8339VhVCqJ7IQAvuWBz+NvlabcZQxv
gUuz44oxuR3MOa38+soS5nxeEfX6GmfEE48fsj4QG1Zj4A3CfgiAX/ukHT2/DFfSycIMzXjOWNb5
14AMDGB8/dPI4Dm2dx6t5IcbHxmiSsbKktqKEvNchqs5HJZzg6D1WsBOWrCaXCCaVBXsWpWkRiW2
Z8gvWd3MzdzlC0ujW8aJNY7yqAhotyqxgx3lh1mQgj4RXC2xQ4b7RkNfECEO8Gp//5iymPUHxvkU
Dn5DUoClXMgs78EayGByQUpB9iuWETO3P2WK+4Ww8LwEEtiXy/3oWiAugoPP1qMVOeLWCI4y3xnZ
AJnCmto1o1q1l7j29fBBi7Ckd1UdQq/oTaMppv/BBw+tx6ChMDPuGvOsZx/om/0Wp/Mi7x6GdDic
7+//a15DNOmMAEI02BXVh2IrO5u//Blc+WHbd7gBHKHg8GiXIY47iOVnVCCL+IbgZDHEYaL1lCit
WjNJLAwo2UT68AElNdO7wYxFFrIyx+MYSuwrIbuF+31nF17Ac8CJy1rJ2DZBKiox+IybAabIxMl1
FSxf3qkYA0ARr/aOD4DaI9Skbf9aswKlUYkecm2ebp1rYrYmTr8YxGZkXxqPifLcfvyiw6pDT1Mu
SVbuctUo8qVGpX78tYv8UayuK3w7TaNu437Rz3R4X38skOWMy3z2UQexN5gMj5Lplf/ZTribZ+qW
wx5m5uGu6Rb/4C+OSBxl2xPZUIbjOp8l+FsZ8+52/7mvRUf28lq0BC/UnO1z8h23UFjt1TqQfZkg
abLFHA/H4bUnahCzoaCgs3cQMBVPs1pSWSWBFLj58SiVRWq0pODoMKkwJbIi0jl1icae3rhJSi9z
6iGUN8Cp84j1pN27VqzakwXK2Ee1V2NYjMSm3nrq+rCLlDM21FKZGSMdJo5/8zHmlgzL644DTvkk
7vC2FY0vo1HGMPmW4Ov+cVWkufcpLFgw9r0KK7AZUO1A7ko+GY21//c2q5y15uruG8gFwRPX5gqk
ttG33YR4DwQOw6DspyKn+ubuEeqUgriAUE/pQrl+8vEbOa3pbtQVDR4KEvz7HHoAhZQr7Ml/Texu
4G+j36pvc5X5PLfzIY35rqu+mcAMzpj5UQdSYMGL5mH/XNBfnaP0l36T+YtwN86MlCqfyEkOctgf
t48Dp/1z+D1LOeMllM9zurDUEt4laxbywZvgTQRj/fYd+wAdvyMu5TpwJV1C1C198zzwBfG8vLZq
lE2I0wA00Ag8b26PIU0LY4kP37lnMuphh5z3JorqHMN2ASGXIm6/0I57Zqz1mPQp8UEOiB0EmebB
VU/OhHF8skvB9uO/+FTAQ0pQoQtCgXnh1zmbOj3xbIfCA9frPzNymqMjxD28Xmmqvf0Qb7XWXWr2
wMbs/FyOPalcwMyK74Qs5VLHLbrjVYT3xmIV8igfTjjsRzOcQQMt+PnsrQrUe3NWT0WNSxUokNJD
JQ5ZJUyOmZRMwhEkkQ8+f/GjLtrbLQmlM9YrTJ/kaGJcyl39n9guoINokFr/uWlzlkVgBakhEDuC
NxGm+colGPfKNTuDVsNTeJ3B8k1Jl/wuyww2BDu0peduxXSl93Zs9vJkNiGfLKuTxx7i+rUDbmgJ
nl3uBmlWEOhh62HjHBdO+u+Ab9Sdb0/SMgBYqPodzk1dl6/DZjuroAsCbIUUBQT/56xpbi+gLpyd
miXwe29UAYBgaR8nmjJrbkxq6YzrEtEcsQG+NtcrdodLdzRt7fegF7enSDaLXjcqX6dQc3xaBoLK
BzrtgWtiG7/mDrTO9vzyUwK4EALjaombW1/imUMTz92iEnRiUqLg/8FjcK0ssrvEB+O+eZPZc3VL
ksBzJr+27C3ZJzirIHbG7ua0UZ9c9rYLxbm5tKFl+zpGxbAKiyZUQydK3utDd7M0Z/aLmAhOFAsb
zWrabKOqG9koIwOdOmhr82jqLDrGihuyAIlhySmGKo7hs5iqVsD7q6mMMHlUphyTPuTSMKc+kK8C
q31vBeOJ+7Hs/UPtpupgb5J1GpYRCOygoXW7KhIFkQ3/6fJKfes7OfkaNMv/6WYwiBhamOvrtoj6
Gz2FhUpXF87Y37aOQ5YbGqOLZgue0iQ5Fpm1Lj+OLWfFBbt2s4nlFt2cYneqZe0j3s3OhiWtMdyk
qrCsYmOmKnlMCZ6JbKX7L7NYjapd1851hkYJRlo/7OjSA6EXrhUSwg9KKlfxoLSRRchsh4E9LOmY
cqrO0RUIskwUbXKXhjVMT9fmh+UXdZTer2esnWonUm5RX6XqkvVNruOYXOs+p+1A9ii2DyVQp9PG
PAp+PCXUNrsrtValVy6qB6/3HBMnk3Lj6P9QLnz9dMw3ZnYRgHwHY0YRDYPpkEUdbhJ5FEJASLqc
UkV0VspdXdEBOKhBOE43H/I5UOO9/Jykb1GvO82Z4zP/vde/YN1FFsYPYKSJ8roF/dB+j2uGq+ds
N9pbBSZPwf144raVNrXPCRnAKjNhLhQYIsuOGdkpF1kXdkauYMMPTVuEBbHwVC9BiVRy1+HJce4T
FxYW7w9cfEzGFEqCUHmzVO0iOWHyfoO+OdwViIiv9K2bwjtrksayuwGKQlDuTK6LoN3dRs3/xFdE
6b6anL8H1Tx0bQd535lOAI8/QqubbDYl6IcEyv8rF+C9tLXvAADf5zuLfBb9bJp0v30D/rSxWN4M
eGIVeo2VNf6mUI7tQBg3qGqf8Hhj3RLorNWsG1JC61ROD+cWEr0yMif0mE4cppswspSdmd+KEdC3
HOnOC/taRQXNO5iZoW1+MG02U3LTsro0lSrouMt83JJzZ58EfCC+g2b4f0jClqN/V66X7YQ2px+g
cF/r9K1STxUn19U8pi4+6fp8smBWXi6akKEs6KYKj0i6zvUyinewKYnr481cDZ0fBufJJeIltryc
DL6e0Z+Nslo3va0eWWbI7xmHXgj29Fe33HbXh48xD94k+C1IYBAaKWcsCmnIwatd2w1Ou5PEhloh
Y4scIeQZeJ0NFuD3aWi7cCG69Tl1tBbiiS5YFQnXVTOpcm2Zgak1kb/7PvOagUXX4qS3tnFxUt66
b8aK+I09jIC8v+ku88G0zanLvhAC1/yfmMfu25IqRW2u4Noux+OIV/a3eHLGbfA6dmcnY9mzOUmr
iScqj0dxs7bvFxwW9zVEoc4kOvvkKga15q6eVm8K5L0blKf3KbYGc+OiEuGrBWpGBddBFsgy2v4R
yvgmzRVVCfOdnDK977svBPFPKOCqrG3b2ciMfVF85kCwRpYGUoR91i5aDTrvo9nE3rHQcVA3X5jP
Rs/xQj16KPahb3AFT6ejVVvd+wVYdSl1XpTBucEsPrSNOEQ3N4fLw9PvmOkghMBvy5dnmFAD/CdE
yYPlaAY6Ix1P1lBUTuh65v5DCg6x3hOcwzWJjrbKZYC+nMimsGDnpXbIq+rmrT8HGLGA1V95zdis
dtbUP+g14/Tq91fpzfKMa8SKICOd8u91VgivJkL72IVoWac7SDe9ODV2AeTZ64I6sL1uXbcwswgL
iqx3xfJPBmcAqswFrA6JFgcLTKIPfGdT4AhOaW7JDoniUsRlw7bh32tfRjkGpBB/POjKX/BjHule
ZGDTIwaVgpji22rXY4VP9Gk+AFZsZJ2QuqXAIPr/Q+xoagf3OFRS0oTLqckd83MQlBl+JO6v/Wr6
/Jrego7BeBYF/3E4bwKXEpGeqb8T0Df5zHqkIklzfLTKEhM/iNVGO+GNUUmtDTuLPHi1EzwHyJq9
Psn/LafRqEvtiu9H7t+5vNrafY1y34BCOO6oQu9w8/JzzEym9BUCIp/c1B/fQwCmd5xlgvL3py5K
D1cZrb1OXm8ikxoSMQL39xXXJL0xUwBu121D6ljvfdbOj4xmUz2tCHWxnwwJ7N2OHC/JankOLhEc
F5fygrTBmML+x/NURp7cH2IHu8W9x52YKBmBITb9n3cSYJaVnTscwV+DvD+71jY9y55IcXisV6Cm
0sy0WFHWWac2DP9GNiphTF4TQXWG2q1tdqjX1fw4eyVHIlfnkK7dZXU1hm3Ss6Qx3RjFvZmJtal9
JxqcUnAepyy0QG1ADWYniemhcBcpnZEiaaddZwtXu3g/KnZhIJeNrfrbtE0jYc1DWyYaq2VoFWTb
eRzO3J03Bz8uhfA04ZFXMhNSQXY8JtZ1lx9ZDEukwK8PD53d7g38WvCoFpFsJ03kAxK03B12DwnW
XcrSjrIVdU+ZkYDZ5lYfOT19pbmkTXvrzSZAm/Wfg2pk/Csrh/bvuCmXMquGbtJLtyvMjH6HQCim
uPr0emtKMgyB0/L9v7NXc30+YBVTwlrvrIukGrQNMeY8PRULK43B+NPCxt2FjSf8UWQPks5ZUJK1
rEBRDe0FRQiND5XX2lbU7rF3p+hvAxV38PW105PTg5zrUmAIjz2Rj21y88aV6v+c1WvyBu3LchPr
dL+txWCqyfq5setqOKHOb3SJYpjC+AlwMm9oDs2uepUieI5sfGJYTdRDe8b9xKtd8MfAyLuyUTOk
layBITUjrtNpwBwHDjJXzXqi+GLHsvuuUJut1LK/zqzIa8b2u3/GmxUqYD2T0T/1+JY8J6tdKXd9
27tdoQ50QgEekXwT6AZimBZNUzqCKy0c87haFYeFpRmaIXL4qHvFzSE4DUHoRjlxtCVQZfzCPzdk
KmbQtbLqkbs+oVAzPtPzMgUZ/6lVKA21gqD3YdpOg4VmDZIYZ1zaybCDJCsAmlaC+sh74mcMFt5Y
PiOFsjYuwdyu5oUoxJFU/5L4efDrIuVcxHJ3uA8Rb7dCvErO/XemGU3aO3GlmUGB7k4PTkTVIqGc
1Uu0GNhacloF8AasUYAVGdbeZ3Ujj3wFepPQk3kktNVBTwutzi8cP6oQdIKn6iRI4yGrXnAmqCvE
BNhto3GwV90xXXzwtn3OH4FDrxARM5aGvqmScetmTWy5/PEnqHtZSRER/5zSZQABkcGrTY12izti
ayrPG3RV/0DYXX4XIaKSnceFTzC4jgRtilHEtrZC571o8CQOtbmN5xbElDHRnnem1zHiBGFwokia
YAROkLY/P795hgr2oHfH7gZ2pF6saB8AJtgkBzyqCPiWpvIPmydk2TAbqtIcxanXjT8iFjFnXJO+
5cPsJm3lFuSTp6H+3xdLoKH57TAKcxqvCG07UUwYb7vhfBsl7/L35zO5ew+dSRnYQTScoeiD/tC8
rKNkn3fugn+WuWVaPw6v5X7ixzmiuk22iKLiXdsxL92SWGNPfPzVpRr0UsgBuob6vcC55ZvZTHap
YKtDP7TOZuGHe/8TMd0AVM5IaA+sfXCgfl9n6xTWVqKYNylLAJDQ2z4ISgkAz7oc/mJ3TR2AJOFJ
dvmBtvTos65Fq7h6FJlfRjgNHcTs+qiz73FINQTJLr5CQXDcMXkBGcvpWC4VIouITlNIzvbEnhLG
j1E//yg2UvBc/4CvkkNzDC+mCI3SawellX7Z66JNUQAlcX7lv9R5UOE282VBkoufUEz2Mq4043iK
cj+CmqPeWVFfmEdwUekiUxNRgrOqB79bvgQ9V5l+lGDJ1uqID2T02zhninKWZrdLQJ/Bd0xsD5ys
XJHPL59WkTvbW9nJQz0sCTxxd91zhGG5/miBMKiR4wLrnHJ9C2JT5TxBOxIeWigfcOOK78MI0yjE
hGuXAqKHV8EPLfSFvPKzC1ZoyRS8WLfsed09bDgpfnhxXM3HCQc9nL6gbxRX1XDa1XfaoVDfpWeS
EeX+c0kB8DeD2Kda2xvsklYaGeLoRQ4+PCJ53ay5TpxFe+5HIE4YiuswfZAwhEuxxglQY3aoc/T9
jQaVyJUF332bnq3PTO3HQ3jdWgH5DRQduEbduG+xEI18zupSH9wHvSsI223wFY78yeHQg3+pWZ70
1iDdgq9c8YHfwAMpUUClj6aOhIr0rL82XxhVtVT7qsvuNiDaJqdp4Z8l3UIx/jbMv37hUNMG5IYZ
WVvOe1h0dTVCyj74C+17svKDMWGLYUyTnS8C4BF0Je3HHtfFNSMHQxG5UVGdzQHfWLiViE8CePkE
Wo9b6+ONMGhlMnzjRthmtT7pNgb+v1rGXk0c+92YWJTMQeTJE5Ds0V75ncJzwhbdXuml7txENTBZ
OXdaJuhgI5HcZaYKTpR6MIgkXflZX2ryvAuX10T0cKO8xYFtipVbf/+ZGOuoHUEo5zPI/41Yw39H
zl+spYlkHfU2s85uOS5NXHbOz4jbRC1gQpPjIKbOWJc7QHEcBaL8olxeP2RGg3cnvd2TSDs5B+lm
2K42D+wCT/BDOqHuvOEx4s/+5SYl5FLmm63wk4Kv1D8NF7EW9OA4za/ETcdev9V9tZT/xfWX9vUm
pkxpH0omQHIyFGHOxllgJGLJOotHln9AJV68SjOxLUTHxcxACewPopT8NfbVe0XjnUgbKPKG8AK1
ChavOkQkzOGkC1Hd+crbTLyiQmTmKpWmx2+Fdmf77SBlis7tyk7V07voEN25WbNjKl57dzGk5Md1
9uee7txI+L0wMBrVOklxJJq26Gf5fb67TzUA6dHk5LqaVFa32v3ee0KjbmRtAjzxBlpDskGDrlfY
5g5fm5Br1gu/SnaohKjJW+YbaJBq8mAyIjAH6VZrNVGJpNlqK/iWiq+5KsLaWOH6c2bHSt3tC8z/
WfpzToxTM1jMnMgPMTcu29UlGC1QTsZexhsREmWQW1kh4S+KovZowXlPrEUFJ/iBDcHqyfmec+91
5B4UAyaUJTGz6v4embGlJHSL0EFWH2M8iGlDMUnOO60bB2gYEbNx+6cnJZjapM24Qf/K1/+XG/8B
klxoK3HsdUnN8kEUIGPjP826+Gc7VmZUf5ZkxM6jEwswpxdKE9GSvF3z8xghUcRf+ZDFibJZkn/N
k3FirhvFfqm+gxHZUEGq/uVXvaoqm6bZm619KPDESUQt6GbJV9BS+amjw24rpK1E/WkhaZ8bv7WC
sTPsgaNs+PrGbK647iXPN+t/1t+OoZLN9CVsfiOBknmKY0uUrSzxeTiO0g9yMxMekX21w+71MgMn
qSFV9aNDXPJLC+0wdfkN5YKQEWbQtyB2yQuuvkWGNsGbpv0n/3le2IklJQwSJ67/BgGO+cKmUZz3
1FKECYcetw4wmYMXfWUbnlHZWP/Sqs5N7v4Kx4rM00qV24bvYrVzltaXYHEZ4qW7YfN92m/EW8oU
kj7z0t+riRCQm69r7YUInGCktgmaiqrBAvZh3qqAM55weDTI4e1oz1ngR6bXrOQbHP1rMszIJt8i
mGglFxcqTfG9puUPH4y23wC50nIFaDkT8o1qn20kdacDIt5uP+MfsJE+bZM9EG58rGeQPxyib2TL
OC14Y1oNW5Y/ypU31KNw191M7shU+uo5ktjaO/mQp/OcIkNGsbkZtAZvzlE1EyU0+6DHIVXxm+Ke
DqfDoP9H8yS5a2/wPSkN+YPgfftWcIkH9EGATepFGM+G/lySzai9zNxMeYkM/ICUkO0tkxp8z+Oh
IJlABh/4VVqODaUvTjmJ6MMuGol9+2REM74dgZsVndAT+XJkH4MB+rV3wk7t1vffAeLQqMj/gZ5U
Y/SWbCa3rovfBFeR1xJ24AGLIFgkl1Rapp0clVu10EiEyFLCt4rySnW38tSsqgku4Rki/PJRYK9l
0sGcqHBWyOzZC4+Ki551ohyihamtbQWViQhg3UXOLcPDYEWFOfiwJVB2qBMJu0cKM6XbqjqJ+qaH
HlaxfvtXYehuFFqxh1nReR9AGYPmB69K1oc9aKwStths6hY/UXoa1N6iyDCDx4LuZYcCEeqGo7m9
L5CBeZMt9yO82hnBMayenAvCbLKJ0nvsJzbAmjAmvSJBUsYKc5FnObHwHg14aOnIOd4CcBCPxj/2
8FuWF0e1qQ7eD6cKOoMylHkP69x91z6zV/hJ/QbK/ikFH4wEdn651egGbdYCLYu7tQu3nlRmVqKR
QRKWzNa/beWXgvSwFo/E/OmvkHIqjoZVUF/lny29rQOtedYniX0VfomIOo9/w8ROO541dnZwfp7w
zgbZmPNBEsZ2n/CHIqtPPtq5F3XNQ5D4aUeVJTVp7BK1bCbaWBl7Q7Oi5rboTwUDFGNuiaH+AVQe
AI+qnQ7EBZk0BaKMpWgB2zsd/4I4UFvsXBfYM9fyRWbfWU1m4Ynrqy0JyPAl5+E8bflU2JrLpD4l
iNM8vVIlqCheQbNXhaVBe59gER/kL9vTh3vQLG5nDdMoJmnZnm/HT6upyPZ87JhpmYG/ZTIYlPAx
mVQ1918xuyMt0dgviuFWsgrA7yoyOxNbqfJ+uQIy9ortzAjS72kMbx0RbLK1LApSzDyfGaL/KJis
MCtbiPlt1Tkpzv3lPY3uYc8UqVDXOGpdhRTXxovJKyhZDirjiMkmHG8bYoTWM0l38r1RqP1pIqU0
1/qddZBg9i0ETZfWeEucJVPvuBFiQMxz+IuW8bi/RlKt44sxopC656alPJ0dNHeYmxFGMOxHwUIx
NASS7fUvMYW1TYEwh5qAKWHvuT1vN1GQZohWmq1w0fN6ixr+lkEay0ndwJ/OFI7QkPKHkFbmfypj
NImsdD2yhHT25QJqQ7jcCTx/1Yout7fUsCGKaRyYvjsUrgnPCXCqLMm2844Dx13VZt/KbpcCZ8Yc
gmvXHnfQmc7RqBwLL3bNnp0tN8T000Dwso2Vr6afvYW4h8I+bnYnnuSlpR28P+WFVvnESXTHs1yK
puPN5CJUKN7jzNKOyPDKBlAI21y676QSG2nLDMIvOgxhHfElF9Fif+kAbHNhn6NmbGPMDGDe82Bh
Hp4Bb9AToGq0KdniHFfFaqSRPq4RoOHo+bd+IGaFCC4nhYZ7g1Tg+rQqrxMhebDZMgX9OL6uFs+w
1noYdiTxZAr4rGV6c33vLjiWubpg6grPBKH0SPPP2CaUxkH7JmUZ3IVAqel7gdgPDejwiVjuLuwW
uRofOMxb9tC58mIIhmKZS8kaLqvKD+uI+z49/bb6STXDlAjwArg/sOD7/GT3vEVaKIBHuzQh7IAo
AAnT5JLxKOK8CrToLhNBpA8EfSac0lYY6nct4SpmrccuFIWI3u7YKgSmECx5OwcLjkTF7ThS8i8x
hK93TlhRKVnnUMPxn8nZCeblMx2764MtB/2pWPjoZ6hxA9nv52Nv3uIyDxZgdKBZ+db3CVijSsbF
A8fIhcU728D2K2+wRKTnZqN04DZVyQc7usXHSNy5vrqiLyq+wRwpsofC8t/SxU3LgA3ClXO43o4U
MQucVrSJHS69Rjs3v9o3j2Yg7CIrawZ3d0i8ZWEWKOT6X3gEEbdfcrUW/qJxoIwvL519kyyW6L95
hN21ZH27FGROLhBR5dvc5dpRAR9omrjSienMZ1HILRotbVoe3Sk16vKu4CdJIT/8s/Z2lUFpqgRH
gBZH0sXevLGl4ULCVqa4Fq9JtUng+UNib6+84frgT26itVTPSkQG1VsQGNqZ/0y8yy4FTV11XwLw
TOLkY+jn3KXBNbBD8qdEtxJEWZoj9r2fh+sd+Ym9NpfaGAfb+Bxyw2W0ZZHv+u59XRBQcb2D+GTa
E+mbAVItM10hLN5RklEx11XKTeaNPLDWw5iC+9ZvzSgsWmD1A8rjHCq1C3R/AlcqQZjrZst5AnIE
abLHQ3u4TqGvVwgIilQtelmK4utan4jBIzdNN3rla9mdQVaACnbA+4WnJf7CXP7JtDAJZMdjokF7
8xJ4waAbJ/OS9d+PkRKwtV3dDvP/hFM6DQ3lAtH51ewnzFog21T5UFbqr0GaSOnAYooTDaKyLfBw
TY6esYSHrJ770hwvvebyrtRYGjTGP/glprMZXYDizpUTRjuzhf6KjdfZVkqihB+DEutBpJS6Tk7d
3BIxlzoWj0NqX4nk1tZaYjlDaqdFDY8HHqywUg/7e/7Lc+Y0Hp2JFJ3TsbzuTLZPr475XlmRM63W
wN7Laby0HrwPlJ1kdP40Ckc9NSy5wo66n0XLHiO0+AHZ2HRDk4cfBf9YVvP35K7vAjeuLTW/sjh1
Zenksbcpkvv5eNBjZJCrfGDi4TaIDU00O9vfmtIm2NClTJvmxQ/h/I5NPxCSxuqntOgBuHTuOZpE
L56SeUjwzviTqgInFmJ+rS8m7jHBo52AKFGS/CvUHowPB5EE+IT3crX5NXinrkLuFwqq9uvecsBX
vkKrrXytjRDWD7N2KBDjq6EHhaSAG4kadFihb5m9uIttI43sLNJ612okHMVBo1iQZKMfwZaljHJJ
1aaUCiT2y/5t2j/icc4wYAb2PKMbYuOthyiW31i6W3kaEePKlYjYpqM/H3r827z8HhLHbjVsd0so
UX6fN2mfNTom1wgZa4Mf4wTZj5yhp2TOdrldcPDG+cZrk6b26OQ3dz9fJwaIAdHp2h0G6Yhq3f2i
B96Fc15+BFhyM1BQjkCGzMOy3aqr5WjPI0+vWXBUmIZvUdMbzAOuQejGAGKGL6X6hvXpE/SeWGIL
zKtCbGQXuV6/HuJm7XX//cuW7Y4Gpw9V3otsxgjZZ3afFA51omCp3fFmjbGQ79IhArUfED8X4/XY
gCxUlqTxzWhSPCS0PsSJlOm+hqwkDLnZSOUIY9HnZ+e8pGMN0kF2+3y9oGVadftWJyfnmA269X+r
BMebWubkEnnt6XUfAqs4giL74Kzy3qL2iKRr28kc/Lw5SFTKoVigDkO1gTisoR4vS+bjQWYQizgq
CnSNxQgY5sQmqlj8TW5NsCRcDXSahKRZx/2Kdc4YEfNC/uOyIwRFK9isPRtPldoRrTDgJ/o9Yq0v
Dsw8kbMVw/qjv5xdhC/JafIt2+CuoU2zLsPpmoetV4Mkb/lEN1FrEA28SNP1Pqy6MF9b2zHK+27T
0+q1+r5K7vV97OUjoycVeQLxwz71uVJjihPB3oB/B7OYAIEQ4EY5k5Ec/+UZGEZkiABQZG59AUuW
FarwpH/OFEjwof19n0hjVZnfHXWqow2QOoe7h8Mkoi6SCkPQf/iKhJTwKoSGX5F6kI9Q6QdJP75f
zpd9CD+H4ioZj9iS+9bW3Uy/CzlHUpRWBlU+rMH/TUrRYKwisBHJV4E5M29D+E0K2tSS+aawIvju
X/cr9cE97ILdjXoVaPSrTLjpwjDJeEcDV4JX41RFYjOUQJ0ByqZbwMR0WvtA8RiwWz5mJPgIcl9C
kfwZyYUPJq86ZogFpT1OKGRQNLw1zjbaTPEmdwHphhe4pSNXlyUhVmrL0kb+1kSkUBncX9dzN0VI
7E/TT3LL/vYQxvkw360sKMifkHvjtrP9d/76w9hzMJ3M+AUN99Li1cmjhVtlo8t3Z91nd7Nop7o/
LnSHGwJsiu+D36hrIAwm0fVagNaMv48FTmtdyCTyWF9mkYOfmWQ6NmHf2AfvkfovIxAVdfSCIbDH
16OZmnHd04W3nhOrHCz7dTUzNtGF2wfvUGq/QSY+gi1z9SCzO+5M/jX8cf3Bqez1coF39sGBdZ/7
UdEnczF8mgWtTkzgVk7n1LWbnFFmhMHWUKplVNK6Xr3O2f5dbmP5MaN4T/zFCIGtIvggLvrfSVLl
MyFz6Mj2X3p5k4dGxSflKbm8BUSNd3mGvz4wGRymVjFDU5dyiknsVavstMKVW7Ln4D2mQ+lnu64L
oPRBMVhQAMcwAT7mhMehfski6deq6aqsBGAjkkXSsGWyTN8TvQu/s1j/g8GxlJ40UeKasDkbhr0V
nAhy2eD6EAMlcmB2HTZ87tpE8161Txt6EwvWw9hhE6CRGFcCYVwFrgg7+s5XmXMHRNlv0h+RaDj4
hzu6u1/RLNAHNfk1nmJ3WmHgPpcSSOpimG9dbjeQfRhK6H7PFswsnnc2NxYoGRVGwJGs8lS8WjM/
y0agkU4y7SspE0L2Bk7U01c6cw2hP95bKXCvBR0Z2+JHerqIZEfBZ5Lc8Q3JuMkh8izC8pghV6rh
r7R2oeZOOVY2JRgsQH5JsxFAX3EUXQZ6mnImgfGPDKYlSlsVyzh8t7QB084hf2V3exZ48LbapfcW
jH6Y0NvKB7OYZJuKxgMnYcZT8E+Jyypi1s8movJzoskt1/YXeRXaQ6Qp9uTVPvc8IfgKlJIFxxpt
yA4u/rG30TDwZpIM/JQjzJxfhOr+Q3irW68xcQj1F08XI5xCLfV0nHgqeYyKK2uv4n5QjvjVPSg0
KXLlktYFS7dYaJW3rrQOnDFq8ybLWGukMfE962T/YJOfKouBPfgVcRH+aF/eMAMMALSOfSDKecNE
KBPK0WmMiEYJm/gSIeE3nQOP6XXGw5JmlWnGBBfpAoE/p/KP96KIFBFpcPMpb3JAHWJvZUEPo7GY
EZ6rxa5PnT9e1+38wn29BywJJ8fHa2YaJskVRVaKQyk5YAcHluoDSUC9MU+cM3h41O1yUvKKcSR6
BANvpgw3CkFIL5TjGon2Frs3ij2jf40M+/K4vcdwZmWS59gXC959F9Qv1Cc4g8b1zWwX9XYYVsGm
jMrXnrF+TwENSkAd2EVjrw6qQZld4MO7OigqBd/U8YbKf1skxh3H2Jx71B0qr5uF1Ta3VZzJvv0+
u13ABVgkmOxd8ju8OfVrsFiWovYaunpjCK1HQwXqpiDuJbpFxhg5lqe697DPSxgn9hve3rqM7biP
KwcoA9j4BwiU7ga/B9YlYP2u2m5JQcyyC6wucVRnvisztuFEewHK8UR3vEH1ywOAiXncBBSKkh2B
m8XeC58gFHDfujtZbjBH4+OsrGz+weq/jYRvCtF+jPr8hIka1HU+uG34EwUwCxSizWLjBEyFOv4t
qKVKbSQAJ4GlNshjiMeNnTlEjumTz8ttrgnq0QM/o67n/AORhm0LqGxlWPE0TP6/0pcKDnoyVHQU
cbB/XEtEwiOuQqu+t00vLBgK4c4OrttSftWw9RL7YWB+gHijDLA1FU3eMz25lOJ2oZagzzg8Zn+o
ZIseDes1PG9dpPfeDcbJa8bTEadWAEQ0wze7mgTMob8tkqvrx9gBLAtb7seikqhOYN3nh+67VP7w
PQSyNe10SfaHENcsL5XFNriJujv0KqObUpUkl2GFCynKj2QGTql0LgVdkdVTF2Cuue6yTfQr8G65
+exHnZOCyKoR/fXIqIIKD5QJTpQaDPKkPHccqbJguAADDF9T0fKzS+MtHu+rcntC90nTJuu4j6+/
5EpW5HBQSX6QVh/lVbApSkNsRNfMfrUzkbIg2ebcPUEwlyPg/n3I61v1bhkCqfJ7BQgHt1JuUtul
wJtyxZsLqdkg/6ltG3QlxhDjGCzCTmvfJCgUSS/p28AuVCLuOs9NqC0s+a6qIbFxGYVqJXIXbVUq
Lw7+CuiCK2GYH5xztbkJAbU2rNP66ZGhsjQgWw3N66IXzLz9mYL3yVNPEPCglZcQaaD+BXdJEN2K
tLiDmSAFWcwyGxp10d6yceAN4tf/9l1hTu8yXQNSbZfbc03ios0meWxkaEdt3OSuPxWnuaE/fywG
J6sRN5E5TSCug+a5R7FZutPSTVY+9tBQlkaNoPOE51g+lxNvjm0nllRJY0nSjSwEAtjxD4wWkPPr
mE7Hq9WbhbkyoNGv4O7TbLwYiIUGdG8FOegL7nxXrF7GRjlNeY3TPb3RzUbtbbxKmRxpQegga9F4
bUdrVv37zPdtJcPrnOPtf9hFquAZPolIJ8hxBzngxkweAwfKHjSY259y3uS84Ko4shvE/Xc5cwVO
ziZvWnm5VXjTmWKiuoQeJPncvrnu9Jhl4nq0Z+L749eEDSXLGdNrmnOICH+Z4hOQSbm2BK1uFqUH
Y73lp9MZgLdghHvU9I7IHrQA2sDdn8qjFJxAOkq1dnoe6s9lypLspd782QbbV/1lyqUj1ov+5P39
Ns2CcX1CxhrX0EZy9O3l43xCTsxYyL7Vj43kAMZK/pXYPha/h+vCzSvSX/JS8VHnYYngQb0D9W2b
f8naRODFJJEVw4pCBiFmFDuFQ0VVry9u0Aqw+PAdJ/OQ84yiIuxfOKDdK4EuQGyf0Dve7TlH1K5e
XyOHZIs1ZAyfEASP0q+FQDCs3iG8dDnP7qV2N/Y3ZxifWvr7zCD2mG3xFq4wlT/2gmckN9tbvlr3
zLfWYSwFSkeyys4m/z+ex7YSS7NL/8m0pCUSRHHlpuvzrOZmhQXQDTAbZHTKjXYw8i9Hu77QVILj
A+qDbpAPCh50kxQtVHS36rBJD7mUCz3GSWqirYqCabl47Ot68mUTYKxSYW803KDHMpTiWO1KnN9j
l3UoN/L0UXF0A26QWw5Y6sfU7Aj1jutQO8tmQL2ReyhdVwSorXaleY+8l9pJfpvo0E/sfkl0pPqY
BWbJ2gYlUoZQwpBg6YObXO47lf3l/+2FgAlQaza1X3LdYOH4kUxvsHeK1KdGXukyUcwkWukoojyv
2jVdaNq4ckhXDRZ5aL8fxRFfWjbJp082Q3nHoUAqHh4BLld/W2ztnQZ2yqyg5jcgQ7LpYQVbVUWs
Yc8vei3t56tPbK6qaeFwc9/bYJVhCGl44pLdDHCRZ5itR34cDhtqRMojPlkhT5MyqynR2KrPjp4W
gsC01h5watUzB/Y++s2WlgzRVpDcUQWq8C1nXDYv3CfJk+2f9mKb6VVmRQDGOzA8y2LEO+xsfitV
e3rOQEhqGKfXfUmwOJjEPceBhKEul9zZ1/1+ADYM9Txo2vrJ6vptpUIqbi5vJ1dAjt/Fr6W/Svoi
0UnNoaUb3tG7vBlHfw3Yf6oXxJXQqUIlQCSr3pOD7DPObECHBclMSk9GdlcF0rxlcirxDSRzWj4C
wsJs+mYErf+6l4b4AfIWit5VQg3ofUotOc4JX9m8V/H8ZYt8pAoqs3vvaLXOTNIy6rxyz6SmvWlE
R7XRTXnStuTRPiJ8nJ3JR+0B8wcdXg1LUaTbJqBtwItPi/8cHvpJN84I0CHm+WygNd+lUqjpznCe
54ypB9HlrR3OJGuCrm81jxqzK7Y0O5Yx4pS6qiSCiqpLEeAqmQAOyfzohqrto/wTV7KYgMROQG9z
b0SNoSGzZDJ02oky+Ln8akSqShARjd2LacQU23BXbM8rXv+gWYz3Ah9E4DTElfbQi/XMoV02+ZYB
+fraWX/Z6d+Wo6lxYvCuCR3YqBcepgNKC1TwF+BiO2h8vgl76U/oGQHh6XTrgIrwjb7fJsLkQ+EG
O2jAWJihbnl2a4cJ0p7+WwIIWDdDUPwksYBuXiojcIEm94tEMBoOXmiU0MaKL1VyUUxi0pBgB1Yz
YVfiwQ5sX7lron3TpSdGA4Ij0e3JltFeSIlpYO2qGFwJ17++eC8by0tbWpJxMvvOR0vKDbhjWTns
B56YYMtp4usRL0G5Visn2/+UQI4SiZNSXcqczyyujywdVAIMCwqXQNankGScIGpuefHLTOK6Gov4
2Kme9MMxUacKUPO6qdJhYujgP9PFkanWb2lslKkb6hsnrXfZcw/VEnde7kIA8qHk1ZrrAFt2YsvW
wwnaXLvY4IiprHMG/hVr5CGdCo0RS9BjkuJw3PUga1W/JLDykN/5X/uZ1IQxud6iENeCkoKpPntt
srrOq6iumq828BRA6Wfuq+NVpaejJ1/45DiGP0lsvRtZISp8JaWBMsW+bLPufUdW46a4gpe4C2te
2/dZY50ehHU5Cz33Wly6ZGITnYT1Mh78rhQzGjd8MxMtYqd24NNQ2FGgNC5F/sNsTR2AB+5UUipL
lQuYi1LNjLJB+GiuD9dBVGt43Uzh9OSF95E+3G61r362yiSG6lJaWOr4gXf0VUcZgagiw9t5HRir
BMIBk/Bg1f1m4Jcxw2k2TKXowkN45I3DIwsy+NA079n7am/ws2P8TKjU8LkBD0w6nUZa0IyPBjgb
J3xJKP5SpszEst2npZxMHIyhn0zJErNEBx2cqMFQklO8xspm6nxUXmVmZRnEOWxWnYtyM68/uhgd
76ZztzA2QqeDKxGz/ZhU/7zTK7H3E1WK3EWPZCueBIk7vxGrE/DCyyc90CscCKCaIwKtBIwwjq2z
CSezlLvWzrpiB2kEZzFvmzzW1/EIkPy1hjVjpq2CHbmaM/VS5iikDKlmENVmIhuzFG6l6ZWsXp+h
alzHKuEIodAS9mxZ3DP4U9Gw/om3wAi8Qh9GBKl/ze5k7s0rYiWT+oqRX/9VA3ODCKuBjYDpbZHV
MBV9R+sDm2KvvK+j452T9kNgyijkAIdwFYv3h9wARhdoCAY0sHTOwYqh6Qf/q3xSVn7rcggogXke
kib5gUyFk9lrAa+NyWc+StOxq3rJaccN0nGQdCTmadVCIDGKmxwDTxWTtjcSRbnvsULg/2bIbMjb
lMTsQ/YB/Ks7I4rLYHf91Pv/ZSAdNUadJ69150Rcr4Xyf7e7IVkrKsrFw1/Ak6I0tzVK38EkUWyy
QYX2+OfSU6owhwWoEFAWCOmhaxXyiuKJkRYXY9b4YAoa3ZuS3hVlQ/6dgNONNmb77YeKGFmEePxf
jW/ZrV4bJCDe6LCjxhMPOUuILH0w+3MiIZgaRLSXazxP8GxUQ5+Xejqqh8GVGKzglOOFCOdT2MmB
pT395U5LK+I5THGQUl/lLsV0V9wuVRXfboTapevKikMhFJcnpLHfEuRq7ILB7jfOESInW15ki+Uq
gwRXHilDQxEA5HNX2H9MIfxp0v58xJaXpwbUv7ymjI5tZE7KGDuVkSNN+pWTYzPFfbHMyvJsx3ph
AaYeRuNZSCz5Xx/iZnqZoKIdSywpZF9QSbjPvjUjCL0LKQg3pJ/puF0//eVY1kbMDJmf41XBFdg2
MJGq/RElE9DKnmG2K6EyVcyHXFaozfwlKP5qhJ692Hd4AU6SVnhlhV21qgq+0fw0XEz4tR5lxRYZ
XTugZoReVdED1Kq3mbQtvJe7ttu9HRksf+ntJSlLxLQZPoNobAj7qT/s8jlIyl25TiojLM1y194B
ye9w6Dh5P4jvwPDZl7ZQt2WkIn1sSs6CrRYylai9rXqB21riwQ8vG//2NysXDaW1g8ZcUx4FzmAL
pndTfL7gxevsl4ZsRZchU+Gu94Jyq01x4K+uKyGlYhiDs2nu3n9gXQykIyn1FUxrdhuRe9OgindN
nxD4IUXjORyGCAAUVyMdi49ivMGO44+FJAfyAVP4ZWgr76uoO4udf6bCqd1fMGzjAktj/SPqpFkb
EJo7zA5075R6TGI/UK4p918I+SaAFTC934a0bmLYQiLBn2txd/6ForeCL2I4uMfJW6GFpPbMk+jD
m5nIW//szAoivLsQWl7zkmmGEeNmgO3vr/90kgtGMlPPOaBsvtLBr60M6f+7GQxixqTqP2xDgbLm
M2ZcNA+3dTLsXK8W+QoMvGwMndFIWf+VypbInvuBv1od4Rh8QB30aqL3SanziPh3anQO+MY0Su1j
t+tn2lL4rUQfV4ih5xZJEWm0iMIv/lrQc69bIv4opHkgTfiSpz1ymg/X5fnfu1dxzILkqVBCObcG
G79wNyBwVQ9J0dwB+0fu0VLj5gO/5hkJ69X+dy3++CDPm+6ihdrXmsNPWruwv/UjVmr/QoM26//d
ljHclKlQuznRFB22epzL9FYijWv6HA6uVXPnWXQdnO2uj0Dm4beG8zqeDq0TEHvKp0kOEDXxIeu8
YIc7mCjX3HvUkkwYCkCsn2YZGKpxKRZQWBhTIn6ZBk1ghnDw5pjrJb97GD79bHZcv4kfZvoPG4rX
rj56tULEuQ2ljtGiB7AGcpeV/TDSFkEToICCz8JlMoqkVQ3FXhaUsKMZb7Tb1nN9yBxaM9x3cSig
xmGec1bdUgT4iWUPDo2zdNYDWltiPJ6Ui7pOZP6QOfcfE/fT2GOBO75f9VnpN7AySg9lnXoGxGzC
i9ZvzmvYZEGBCyau/HArXiWWLKdXNvX+wHsD4Wlm7z0czSvT8h8zm+YTTS2OV8GJKM+6VM/fNOVM
TCp+jnyBIH5WP+t+rvJdXoXwDrgT169uwpX0IB+IdrzpLCVnn9fXLSWJVyVFUVwlkk1dq/id8/1p
CWrIehnWo4vvQqFfQHJyVQ+Pr2rkWig/UksHMXVJG3COLw1RahUqzX29cAn+weU7mn7dYdxuRDsh
HHwnCn9sSYYcdNqS3YophEINyI6B0oxtvpmE/2exyYl6gCx0WZ1OrAaW6EzwEWmvrwIl7giqsXSj
e2K5k0nCVzKoqbDKRXj95xZNtBFMvoOjJkx0dkmic9uWexvo/javKJUdXtCk5PCPIQVNtu5czav4
+uymA869/CbA21l7ZaY0ljx0uAUlmSUNVHPHgtNHDlsKDeSEaop9vePHGCUBZsDmh0mlRbVv1v6f
7NYEZmdS1QFEAXyWcyN0xR9Fp/zJUs1pKnvl2cZdxQqei+nhwJfSTClfYyj+U68pkNA+uq6sg9gW
4+mIaOjv4D1ruJOtRD32D/oNnY2V8P5bjdv1h9yahqWW2/0413KIOIE5/PMfdsub7kr6R2TpVpSG
GyC/HX2fUsW2j2zUKkvks2pLikrwBIXCtF9o6mPtMbhFb1VPRXk55aEO3BDFhQeoS7gr5t0yJYEP
AbcUjiWQ+9UMxRV1sE6ooc6928oI96pWB21m1hDm87EZlj2H403bOYiATWaWn3Rxp1uyYl0JzK8u
0DB28NLWZWUc2tatYQkoUgC+VNT+BkVVLlY0d2AiY9AnnYE8x0ldhHHP5+o3X9phBDlrm6x+VWy9
iF7Qaz3HjqnSyLePQqKbu+6gUD/5q4XVsVXX5ioSWQUmj2g/xrmnLOrxEKYwP79BlQXZscWWCDNB
Lk8c4mTucRNEPK68zQ+PZzjpraoSEcQrJm/mvQYuieMHW5t6YqbBnw1sepMYeAjd0L4EBIHga6pz
eBblHgzWdxfePdzWiR1frhRCXwJbeXwVIkQXSKCD3fhEyZErkA4QXa1A4TrgkwH15vFjq/LMc0IK
4QMOoq+fhdE0sH3CP1PniA0pL/3fcJQ76Tfn12rNmzc91li+cCdv3DGnUtiObpZoXaqFIEnTLOPy
hRxNxAhBqnr7RJmCELk0XKm241ovcym2jTBafSkssddvTk4X/uiDIwAzMR8YzHj08iIVJ8RZDg1e
6918x/B4VqrMC8L7c+KXlfhTXpCVCtCHZRS9GvHmiSYrSJYjY93n0fXoUHXbRHvNOCMRcNeIjfoO
2yQAeP5CrhfQCXv4FiwPFwWvORF55n4eCK+dgbB5cwKPhobAaVkzumPOaUf5zPuEH0AW5ZPZj9kv
hLM4FTCyLgVaex1zf0v2MKAg4ZNh3IQzF43B2vydi/eB/ueVtZoEFVf2VKPK6hR/w17fhSP47k7v
x4OsXrBmVRga2qc1UVhNVNfC0aUgWc4P6YzevtnqiHe/Dl2W8serKxtVWcy8X5riG9xFyrY4sgHW
yz6dm61QS29Wx4Ep/PKuXlPQ60fJpN7JxXRyJm9yRcAZTXSPYtjZ275dxYAjDc5AI0pc+849asGh
KbuCG6p1RzzCIKdR+XtBFLnR6eRSMDKfE3lLzUZ0IBr2tJw1RnzvLOmCXWtoxDBCglag/w6R+x7R
hq38p6lxetNE3VgtYYoor8unBdwkIq4w0WKZq5wk/O86XqJ7Yf1tH4bUKwgB7vSdn5fRkpT8tvts
nXig5cwosuy0g71kwNN4oRSxZvRtjWmr7KD58UVYEoRV61JYA22FMay3C81lKzZv55Z6O2HjMUQF
kIrX+sfrotiTymcm4nXf7Au3vGqV6DMggn9EK5V/mYQHpDyp7ile2S3E7ye4vTs7NFImN8f+XeUn
HPBArmoh2Qwzzf8RHevD1fRlKmP4SS3U44xQ5qO77wZjODu5j1qte+PdZrT8y3M268VZphMf+ENm
baoGjlVcW8eunQEvZp7gSOkTG4BeDywnd6qt8f4zRE4RvayZtr3sDwHsPNOgZozP3cPB4zPzJUwJ
k22ZKyPk7g7OsOwW4WE5gxa4yQhHc1JbsfOsHfvj5+gtBzqYLL8KF0ERQbctudrsQVPY/WLYUSfE
iRL5PlNSEEMTHkKi+abCYOCS7CcnAZ9X7vr+esMDIpXNjNvloqBhu8RT2HJ27khXVx5G1JZOlyR4
0m0kkbup/05F6UZaMmKjLOwBGIeP7Pxce6YIavvt0vJCT5WI8nEM/2tYtkdADExlS673JpudiF6F
tmibFxGsTdRakbS5p8ZUWZp9COOdemzPt68B0ukv9iz3CsqxxCfvJFoHBDkFoqnImkMkfEFfsW8j
iIMRemGJ5O6/t7LsLAH5Hp4uZjKAQgGv9MYn9N/9kcEdNsrLIDEQzgfFqBgB9962KpjLTnATfXbx
h956KtBlPW0jYMXZZnSdgi3O6RytkSzUAgEhKsk8Fs5kxnB2cB4JSvb+cA8K1WG+LzDqWza5VVCy
z0xy6hPQzsLPBcPYYAZgCQ1J/V8Z4mUa2aPLpLRDlRnv0kohZCYYNL4CSiTp+Iyk343vjHqLF0xj
iKw0bAyZ3HzK3x6cyrpGkNaEuWEg+ihaDFolTxQJPKEiu+G97UpQgMF18etvNdiiDAdUW99u3PTg
QeMBighwUTkAPQ0SagDfnYmuRpSjqva3K+PkcMZOq8YxT+CjSddRcm4L1rhHwhPwrOQmxxSlud8Z
kBFxuvz4nJ1q7gnr1m9Om0RCdmHhw2URbwPtYP1Qz02FmZZQuhHGoL+xwZ9/xHiAO4xTpHPsVJMX
gzjGTPC9iaZhmLRVFl8Yd4+Zg4iiiIFBOE3Xp5l2E2C14rW++GVWOrwv06FnYUE0kzwe9T+HUYiF
vhxP6mGCR/p6AB/w915gnz0i0/baWQxP69/bEZBzoy276Z61/oaHvuZbiNTfhaXpapeUSPDdHuvR
Oem+2fGmwYmeKdYEo8uSgPKAyjBRKdQY5n9TrdvlyF+G3C0UyvL4Jm71ZL+xRuWl3J19YMPivUGa
rtQaKf5MzP6rID8K29ai8HbV5CFVPrF0pX5EKPvGspDZXkCTtoQy1u1LcFMRVEiCe2VEUE8hYKIt
SLXuy/zJWuiuNFA/+8UTpgQH+DduiPcSaS5sc8Z9HDJhkuTQnBbOdpaopoioL5pnjqiP+b1aDmwP
xjcHjSQONIriatpmM+EamKZOPJ71snhI7lLTV0aktqIeXevDEMk/8SzDwenjiztFHmnHGguxYKmm
BIogQzLmitd1UUFy/WxWxfyND7oJglKuMdFuSP+DIGa37AqsbjAZEm/jFvCKcFUVw/y9N6AqYjdK
hD5SqwWJXHSp4qABWXRtNiNlcpjhp68att6TlTtCrNSFjh8urpAuw/889pV8zibajznGFGQUPAMp
eLHoJk2aiZ6LzaTDtr3Y3wL8SHdklGNGvOlF3SPyWOjaBs5M7SrvjTvHCmXyzCRzTc3oVTKXds6j
ZWYsTb21npLms2Ur05YPH9Yw14qC1iemi8ObHpQSuRpnU/8yn1EN46YLtbBqmSEiuAK2/MeXM6s8
yZx5k3IxD/1fL7GnSCgtnysRGkDB4mODHQcWSubs1hGQiolqnAX9SL3Zs+CQ5pwFydpfaWkXVI4C
xAAInZQ84w1hh0FDo3mcqm9kL91IoO8YR4P0rSrwzuBUEwakOl1tZDyY3ddtQlUD1WuR+rzyzRjD
sw9loXkpM7ffAU8jZVktOOf+5DmelbUn0QGV/WvWdDudccDZ1sDD1xwrRop6X3G/aEs9cnLpApZX
Dxa75EmjLiao3vGTe+R5TyEfcYgKj8bi2y0uNBJ1e1jcomhRfaj5btHCfFPYVu82UstDpoLs1EAZ
iALI/w8rKLBPtmFc6V5M5ecK//Ab5fJ1N7/BWrudd8UKRarKaSDG1oYRSAa2ENfHuOj+2hA+91cD
qmvXBcrslKQWZ1b05SZsP6DNd0vZeBwnWHZr8gEnRtu+lKYgsLiCYE7cNVB0ZRsxTuvVikGpucu6
ZHp/OS3vAngNN6xbycvj0ZCKsfxahHRGnxgtaLQkhAIb8PvOn/vWBdBVBIM59qgvl7Wami8uHxIL
SBcZfMwr86aUVccgKXeNHQxQI1eoSh4GU7PEWglaQMGcTjmapR+cwrAr3QnkO0+ZUBTiCz792zvq
TI0DYszAFhJQQ1pZw62X2eSWNHyqt49lVmaDndnnAGliyMl4USLRcsY1iaLY929A1W0Vm+3aEhk/
XCqTMSSzmkhPLCiFDNV8jsd4E0uQA9AET+6hF4ILMNRxqArJE2dsi0K8enMh3xm2NZYQ909CqbEd
chceVEvMvoL0/inysy+y3Wnz7ztiZ+8ByVLixD4Xi4elv7yZV3hiSFhWqmI1EsR7ygwzTybfKHgh
8cK/4JJoZn1LMKxWaT0zFOuDsJbSL22pQzQHrzHTewfT0F+Bp/MyRfSXqBmcn8KAp6s14E1fCRhU
3uWPkggo4JIdnlaNeoeTZQZddROrnczw7n8oEpT6LpuvIB8lV7JRRMQ3TE8RePjPiG8afv2CsPDM
JKaqkMP2TBikj/o/zGYQmb5nF68z+ZXIRrC3wSygkYhRzqupimwrtnJVJy4QXa3mG2AaIhThAjfe
cGSAhD1AhgQOq+QDP+enBSAwQaJm1MH8CdRWqAsVppWKJSN0UeUk7wmcm6A5AcxMV7ezohEBMwFO
LH3Ly51TdR0/iBQVIK+Stpg8klGOeRNkCHmqGRCHkInc+g1jjmKYpC7Ju7H8aqomxao6558AcSjA
n4H/S7oTOkBjZ98fG6kgVMe92pPJqW0IKEGr8qra+VBVCtCJjWQGuAF42IG8Iu0kttIbllkQOqmh
2trdC9rytoNUQ/ySObtXlSAVXN34c32+N8EBTPAPccdy+IdEZQXreU8Zp16RLFJofVfhSB7OSyqM
UM8bo5TTfohWQxI1eaFp03ix2NlYrd8iB8N8nPu/OS9CMa2hvDw/giM7Wlwz21yzaWY+BM64ZNvG
8XVBNDp97853/lCtIB00e1hngi2tMLK5a95/ePdS1pSYLI2k5bvNF9sK29LyEabQmgWMU66Qx5kS
nWSDvurmPJ77tiI/w//1Wr4LMzP+5BpJQvAbjYoCQu4ml0MmiAKMt3oCu6oVQrSHUhfQI/otzV96
P0tpEYQjgAxUy/dUS3lGk5f3unht13BIflS+O+JXxi4ZtNp8jr4xOtZkqS7HpLSwQ00KuR4qv6yD
WQDt4/Z/tLNHGkFHldug4bLyUGPMfNkGbYE4RYLqMnnbT/ZIMDkx69U4dVBa5zlbpNlS6+5IVt1A
TGWSgAkPvM/tE+RrDhjPVZY4VzC/pjbF0YFRUpuPLWaDIokc/ApS4Mlc1CvyLSbMTKWT2qubMUA9
Nvxbcq41gCMiW4Tx+kwR121EXR7izfS9GnCTtqZPAyVA3UryvtHZVtyl1GVudqv5Jm2N8xGRaJOR
nLJW8Tud9TXz+azRdFJS2w/r4ziipYJm+3IAQpzFlaw2AZ+WfK885ZNxNn5AhiB8B9Ej1E+o1BSm
i7tUusPGy/Y5N+xjloe6iRDNejD7CQ3e0EENPI9wQcDSvIfrqi0zX+VyicLShzGt6fyMWZ06Bwkh
4EUDeexHGDbnQee5HH9KFpFLeNG6bH0+OHujaHIH5yUxm3CaNxnrzEY4u90/bfLTBvjIOstc+d3x
C6Rp3jTUzHC0d6Sjx3Z8ungR3Jk5avVsJJY6BpOv1gwCDikk2b4WE6aEIC8mOPY3xag3IND3HpbI
vVWMDD8m5UJp40i0jD/tITYdh7iFHZpDWQAJhxWeoW7K6qrA0FS+j1ma8sWaLJje11CaTLeebv7D
t9K+fPcRZ9Jj3zDCMh1FwmadT0NqBtASneylDtFJjfIHTSU9lMpuQaGAfZ3smGMxO2rnUMuten6V
u3di7hY8qG5rZ44893pTwjKGwoZBrrV8w2HHZUcfdsdC7D4KjOfmaLxPOwTuRYMwQZ8nd/CffrkZ
jgu4I4splPh0/99PI/1zNI08xeA5CR22dPLDsPijCBQy8qGJ83g2xchcdIEjxNoUUfDxGoNYybgW
ANGncooGdNDD2vqfYFuWmk0Y7e9n+ytJxdhPzJ5Y9NrcHFI1EZWp9qeq+9Qw5LOFDFTo60jx0a8q
OkXHPue9cIkBprWpSOg6Z7UGAt3sXkUrZPemlucWvGWcMmEgvrFa57vQmpyIcToMhMEQgEnN7dno
CcQD5b/HRro53WqjklMhXlcC9xwVlDMW3nGOj6sP7vyKL5iCtIifZUUZXMhvnJ83DUaBlC1q+N9W
I+SPzbTLwqEcfY74d5hlGDZ5VnH27zJUjU9zFAuUL5EgqHYOJDB9Amd44KkyF4cJrUT0iSDfqhc5
4JhqAUT4JbOopw2KwXE64bp2Byvc7930gie7GOiW5PFWotsW3TQGeG2EmNTkDH4YZSiP/ZPma3qK
Jmuzo66I0ULxl/I6tuHt5q80/h6a+j1Ia1zh0vwNLdBB7HTh7JfTXHyNcukGb5Ia5PTK9M2T+uLA
wQL8Jz/zsVNcseqBDqbiQN7HkWRh8wCLpJjtkcQwMLUg4KSRBapsAJJSFy0FzYzq7pctjovE1vKZ
4dabUuSSTDj/x75UroPXJt3WUQjZHvesH3Z4n/yQD/KkCjmIpI6ZFxHyrXmpwep/WKZmKgcyatn9
6JE2V72eb5BEpQE9cf8Ohj9Uw87FZ36McQx2ZirCzGtO/ifUPyGWmAzdsxxmn1cOYsRPUrb2Grd8
ZXq7FDKudO0dAxbTpSJ50IcDqMfJahBRRibHVzGBeXgkBA9SijQ6tio8V8EfqQMTo/vCvk+upxIA
cJGUMxYS4j2t52w5j6rDmDjhxQOg6py+X6j/+LA8SwosKHpLm+NM4WDChjAOpp6k9i/mW/nJmrvi
Of9jvdryvzvRX5HjOeZKZeRnUN4S+snTZTQ/CxhHvXfSaypMr0jvNQjCjtHQbFrSo3kK+24CcQCf
Te556amJV8RwspCzEpIQrG0ZLjBbd2/HhSBHjayXjNVx29OP4ehDofrj0gcv0WAOamVVk4FjUs9v
u9Y/Q7KexwCtosXC5pduEnQjumZNuW8cG1vrEZRBkHKFPcELzusK1pMwKBy29TsWkoKR92QimHEY
K/Q0SFQwC/awgbvbCqXCV4ULtNjCi4yXEaMR+hOP/4OjNxsoGSfoATR0LH7IXufe3KcgzaJZEk/K
Gz3Ox0zSrOIb2T7Cy+wudnjDb8CXvI7G5gQsyJt+4cenR+fAaLJ6m/PNL+KHFIG1uqMNUnrfhAf5
eFWy28r5DIJIso1ZtKYwP+N7UJ/xd2oEocQ/mY7iOj3mAHYL3J/8Fy13SjsBcfDnzdIgYyzlGNrv
cVb3nHptWANZBFVohfNT8uU6+XtrT6JXt2ZZ+kzmgVUKrCWv2F3WT3DJdqaUBoFNrS8lNKS3xfB/
dVBKmwP4HpnF02lCWCGvG+ARl0LQTTzbSwB8grfj9cio+1QRzClayFoTpj5mwbZ43ABuyTXJ6uD2
lCheebil/5vIo2Aavi8SIC3hmUctuK2HgPnsOW9abAi1Up2cRUTzz9gDIi8z67fUlVNLfzsDBToM
Lt+DvzNQx9wFG/VOIup1pjQeXI09emxgiD+Tx8IaXJvoVHNfk0EOeNbsG+rK5BYk5kLfD4MetDGl
RpmU4OhCsY0rqetpNfZjqFBCSnLHA5JNssmYy6NGLMhKReRpx6AfaNRwKg7MjmNpYoayB5+HogQn
sVZWsNUL0Ddfpbs0jHNRiGWFZS+Td0tx/oaOpW9DtgSX6Pjhbqh6VaGlaVjX+7WZffTCOQLHUP17
dBJCeGLHJPLhUoNMkGlZJAPqEFEGrSeHiK6ebggDjWW++7bycAexRX3qGH+BWf/L+DN6XthYj7qD
9EskVSVkqUKSVZ1fF4awoQgTXGlt4MQOm7KcRAmVYu11R2XcjNLCb1mlBh2U4fTw5KdRatYsxfhv
8KxJID7FsGdZE2et6ZLhViYwZ5abNc0GFOZJsumt8fdBHJ50sXZkVjtP9N5RCBvw0gCeEJ43NSci
OMcdlk5k45TaWSwd6CJwZr/K4jQJdHTgN6Oe45fRInOaSe10d9lNSa/r66mgfkWBW5aueDi7FAy7
0+UmML4siMNya8OzN4NUrKLDyV4IU/bQurH+mIk2iJHwuOs3kehUmjhksrfe6eXIBlAJzTG74tJx
ooFyteiFQVtoK2Bl/cTPO1aKIkl5NhFJTSGI0aolauWiJl2RuxLz1ejjK89t+l/UwQcPtTLQ5GMR
Tfhm/Fkq3TcBMn2xoR4ePq2zO82e8Honi7uHaV0EPVx9tdawI1cM0TKayGcnm5l7HX/8Wo/o2yR6
xDwBu+j+rXBdTref3z/dEaeEDsDbitlsBLnT6Le+p1YJYn6MdlU3OiTPiz72t9kIb4NdvFaPBbb9
0hiDI4Mrlyzkn9XF6E2Q8xppSAjt02ZDQwDK7Mjlp2vSfehxeU0Gj7GXqRgRHw17tHj16CqO14kw
XnGPIs+QCm+1vR0e0TYYsfmMjTO+WFgUiwqFGENlBFP29Frd4Go2BeLPXR4YSg9kGbpTWj8nchxo
EMMaUlKZA7o4VI34SbhuPaHpQaXpBsG5qv4flK3QQ6CwcgrW3n1Ii3u7Q4CAItp1bu38tdpIovcf
obSFUsH1jKWpcqeOAcsVllVaKBrjooDA/hSJMgvFbyGSmmWT3Gu2OAIBkGv2DZ9DiLZmcXldb7VV
pTg4eCqYbnVuaUiQs4KoPwpGac6/aZnnPG7DS0tj2Q4Qd/xtufi4QKMyzvJPOVfhmMiqllDdX0E3
aZhKJtodbcwP3DgAjZGUpevl4DQbuy5QKGHmIDHoOGhaRraqQhGd+/d+m4CZx9j+cnsM9Gb5PtWO
YDY6Cpe4m1YYCV3ljfZO3kyO7ISNvO8uffw9U7bMeyuzEqphUO9au7xNE0EX2NDhQfi9UgHwznTW
S+tB79Kvqtz69v/GuwAiQQc1AV5Kz6y1cv0DSnOzQVueIPLLFGJK8rIbLZ12V2jzranBNzvzE1sE
ZJJKPJEoWcCjf9xBa51cvlZZTsi3v5ulSejO/K+uxnSHf4Im2a8OAxmTmm6XTqmTxaNJdtK8vD78
PxfcNnkV4nCkwYKc3MMXAwvg0sPJXKy57NYw9l9/fxnQf5O3eVF8p2vwd7vfaP3LS+JBMZePUE65
tuagBqt1FrXIJqlP/awo8k9JwzxnYkU0v8Rx7D/6Z167xD82Ifo8UspROH8t8aZriAt9yE67KpMT
IA0s/MAHLm7QzHlMO2JQrJRCVy0MMjp9ciTYur0tN/3sM/xzIxQ613Bh/XxlXjZD2UdXiZgpxMTY
U8QTclGpEtkxI3hz/3sATU+oEntF4dNR7lxMFalUDXMizfV4sj338g4T9wi6YWkstTvAbaj/zud+
46QNoezxXtnkVGgpGcr5BWKHaZVE4FGrmihsG4l0pMTsiLZODCJe4cLwAS5ARzoiEx2smXej6snZ
8WwNWXSyrvQb9AqWizYbMSHKG+GAP/qw0MO8qQi51fTJBwQBIlWFbsPMmmofpRhZIcQ+nT5V9+dI
OTCfijqE3RpfEZeZZLdrRIltwYEfSqlNUBDNQLEwaLB9OSZbLJt/U2WpKniIVQqll6jXKjws3a78
Cjhue/6ZKPQ73Sc+7tP5lVTBWhozlAmddf7g2YWYVP1d4Is/OEJ7PsvWNEsb/RApBPqBZt5a4i1M
AAjrNBY1nHEmKILkImajvjV3EAVPicirk/+IkA3gxSh4Xrk8GcwvsSjz8f94jKGwGqEa/S9EPFqJ
T8lPgzQI+3bc0XUnk1Sgy/ml7W49D9CScUZwdSrFZLI9U5xGPTuU5o7cWYEHXB/eDV81G3NhFC13
p1H3K2aZda7G7G+VBzdb2w1awnwmi9tAAEGlwYzl97RoMTjlaBqhKGt9lJRZMIZoMJqlb+/QHAyP
ygH1Shs/WWY4FFmmthpnzkBNT7ZBUd8uP/YnaNTnneUcWfhHkoGd4RAWmCFXCWkzwF96L37HovzC
Haon8Gal9wKNUgzvDqMtH6pB6aY1AfHRzCiMGfnkGm8XAsjZtLF5P6a6Q4r+pT/QVhE66WIEni0U
lP371A3HWOrVVGojmkq6+ZuuCRm82mHx/wv6EsmD2Jf4o/zUtYvmp7ihGW1tBBRp/ShJMQn2yOBr
7Hy8rtwUnjTH6aiqPBj660gXzZZd8vVC1dR6sYSP9dXDu30tpmrooYc9UJqx6++TsCPNKJhdYGjD
3p8o2jrPjaYhnYXY3wxrGthPdWQTELgW+Kclpk6r39F9ZqlloFF4ZDhX4Bgvv7ehpx7ljqdgGGHB
dNWgSYu6+78dnGrG8u+oypkdBsWwdVYZVNh4VpwEfTZsWvkXc5vOvDnNYP2yO/2WUGiE5c+QR5UO
hwqCdYkB+zBlMdi0WvfdBDLz9pzk8n9sN9jAucqWWB61gmQrYUWRyitXPUEJwsmUDUot6/r1T9uc
3Cwoo7URu9PuRneYJheGJkRu9KphRZ0P/FAHFs7eaIRXJW9Y0OjuqjyOiH86OJNH7ry1Pm7gx3uK
d0FyFBce2fMZ/yfF23F4xJJWtT3zEGqtr0ag6zNPG/RhVH4+AbyU0b4j2JzamxiTK6DdFq67eEvK
gJJSe97qhZ6ixD1K2irvNPix8pVDJ3n6drHTXtLfQXEwKY4d/l/WGAKAEV9GphQtA7H53j8R5TGS
EXTJOYcHhQnwTgX1Eqx3qtjOR/jUUN76OfdsjbQhbLo00n5JM5RcD8bOaN21ExS4brrR9wZ7DJ2/
5ZI6V09UKSD+Zl6lEdiQaxa5tRgtaOYm46NyToEzwl2dRHtkDnJFIugJONix/ujQ0AbTsrOsFm+w
xzyJov51z78xeTduVAU3Jx9CkskiG8qv1kUFG9oLDaXcC9V13Q7VhGyIA3CyDPafAi/tm3VYVMQX
XT9J/D+2x8aZr97PXXapWsRhbpR6aUQfW/YvHb+M4693C1/Wical1MMsN3cVFu0KGKZoqv5i3bKu
QZyxp1wwdtBMH/belDslNrM1K4PrLjmFJ+bQBG3HCIdGVgMBdEM3xPEJuOjxMOOKquS1PyFzVnvA
4wBeGpxbEeGzhLx21pGs8CQUsXLnVS2rM5EHVQCWcsQYbfzywy62WTMaRNSfK7cBQLNW9xR3wQDl
q6E8Oxm4ITQqULlKir83E4HsT7gKs22YvZfKyeo3MLnqst3R9GJ8F9utnRmU6uA0t3ivWblWOLNm
UNXg5pUHDyrcMHUnqPxXjmQIGkvba0neoDcbSoEKpymRbbcyt6mga7aT5taHHdi2g8zBnrZVdWV+
QCGc6aSVaz2CeACi1i/ehxGFBPJtbVkZ8JDpXPpGlYhzutMyJeVD/u2Ai2cGVVq9jeeskdnTy2AB
LjumR3/JndtvGGdkQm6apg/clrfPqMdC8UWgEHNtbO9jRzXwSQpA5USBb/U8f3xhCqCBoe/AFWR6
cb8AyOuKRqK1Q6lC8n3mnHBA3zIIwKkVa/9/k7Yk496EV2aF5r/JQawLX0YHjQX/+av7088NbN+6
fuigGh7WffLFNMHszOQhpYvee7MVksITRKk5RUxgyfCtp+wK2kEe7DH4Mwp0QAYHSJ6Zhrq8JGeJ
aK6B8pY4ItV+djB/7p5UL9d7T3RVN3XHc3rr/4P6FeQ8qTZivpOKnyGAhBe/4YZWMaWPuuEXp+xH
pLhxM0gft5nzcWYpiliCj7/+CB0XRzy2qun2DOLq0BgluDPmpFfIqUefWS+gfwgi6CeDmiJJ4M37
XakcKtz+tkXb4RhHyZohqFaYJzpIyeyn7Mrjaj+9VXhv3BbCB2xA+5Aq+jH2No+9QaNDC6apO5p6
+KyK1a2OwLpqj6OLOYy9qMOkD/gx6VF4gJhY2Zj5ckQnemtIBKqGDJxZX5WB8l1CFYSdF2omXyC5
nVbA/0O551ykDrhbkd2xJoQC+RaVIuBtq4xuFS+eDck5kQ1JuQSUgKITNY537xzAjbcujPz9JnHE
4PF+pzM0eOvzJZYgXSZ5Mq5N4bMLUG2JgFiPfOFvwXAGUddVFKoWJ4ryWYcnZyg4IAIpFZuVMuWb
ntD+9+Q1t1vOBdDUuaF2npaBX6DsX2kiKteohoD+d+jBPI8pdMwYo+hlK+P+qVhjAMOzK68p1/59
MhGgKlw6N7ebHIIR4xMbYX7tmdNKHxRXT9wTJ4BMNOf5KPoknzu7dxi47oCDIRZ9CSQQYFdQHh8g
PSKjFyXNumYSN+r17IPOAg+45bTP3FOdgd/UFxkEy+erYap8ecajDzA0RGGf/w3SeeVnJL2qGXka
DOk8I7Giqa+ZX0G7BoBlZeg4lWhBpDlwxakE9OoQmY2NJ7lmSuNmgz9zTcdwrQnQtTac+VVuJ2L6
aXh3r9Ocd8/WzCPozSziTpNqE2+XXr1GagHgvfXu8618bjtZqJRviayYIYFr/Uq3RDsLOdmTy+mR
6VKJkIurPaf2AKmxwz6xYUcqLO52hR19LCf/sTgFk5ZUN+msD9aqO0xjvbHI3DEJFlRwEO9xTenH
oHJbj8PiEnh7lnayhJ8vvbfqrEnkiMIwKgbBNmMGxohsFNjKc1bVpR9E6yIuAT16VjIxGY7xjauX
n+z/zAN9wes3G0WD7elnaw4/XuBA4tIN5MYIWXOZXRQb/AFy014HEwQRoyJX5PLsMIijvS5frkYR
dER7KFNC7tyN3OUt3qZX/K5q2nmgM5QqyEZE4YExHwAiPrY3wTE0eAvZTp61JgOweTJCcDlmz7QV
0JP65kzvlzy+BFa9YJRFSDyJBgU35j0yRhwbdiQaUMyc2PMXcNSuIMM6zsaalVH3kUYSXv6oEPpP
O7PCRUOg8gj+Pa9rKsAcEsWicwoD7JTxiOfjkNZshGHubPBG2DvPBj4zwbv7X9RfTD0LXsF9hQ/F
jYx8hfo/mhdBjeClViJtEvNyU0I4BbWLSl/26ix1SQUyiWGSbkyCrhE+NVU5qIR0ji95Bgmxg8wb
Vg5XHWjfcsaWV6MXliC21l1CucrrGNShrLuXBJBbwfXNlQbHq7w9M+DEafRgCO8qeKnul/z52lqn
lue16iVO/fY3+450JjMZdM0LXk0pO0FPEZW4la+gWyKsFQBqpe+vuKDZyd/RwkzuPPQtapr9rNIq
mrswspgsmIa2CWPA8ug7UxvmmEP7dns4hyOhD1GN6w1fSqd4/3rFAR/1V4ZwX0/j+xgVlB+sTIh1
5xBrcct3Yue5lbxADxQgajmwU8O0u/hOzgdi4w+IZmwIBPhJQ4hhjLL/E9V9Hm2Zh4tbh570dpPg
xZAIf1YzmbF3sGHTXyAzQKvsBTdWymJ2WwDjJmKWo8SearX9Nh8LZ/s9GiotwSJeeuz6YgZvZTWC
9Jqj2KakJtIxJLuEIX7GbxchRUJZOt/MZYbznKqSfKyw/ElLaX9rqZclfZvo8QxBLrRUGv9+1r7+
wJXswIGjSgvKlo31ArwdUXR4cWd6VeOeruY27m/eP1ufs6i5YHh+soiCELIM5nSs3UFa3EON27f3
KpCvDKgGZhFEv+esT1gbkN2Sg9w1+GEHGbOYUNreYl5Nip66ZZC94yD4Hu1fx+AE77g1XTBqdchF
0kppHubJu/vmyRoi2k0S2KG1YP8UfnegcJJ0By4TVLKj8QaMgOYGIefTxoE+Qf9relnP950UqnJk
+3X/eSLRPVIXrHsVdD1cAQKEIk4EnAD3yKEIFyFYRlzNqDjE2h+X4AJ7SceC8sHzn9f2kyw8hojm
tfvrj7pQREpWHP9TWZB8IVbsi1UXc9Vrih3rnoWZvEoj2r4+LpAQNZSL6rZBGN++gWMgsPVUAQan
nTErVuR9R8OF3h91TpNw7dXCmFvMHuhF/OkIgs4Xe3MpU1VbRaq9ifdBn5J2sZ9D+ysXs7rbHsVh
drD0sG7DIKfK2Il37OWVTjU7WmPKQUUSHOlOXUjbyt+RStfA4Tsm+1RGx23jBlUPJ2CCPYUKeWve
UXpDkhnx63RQvBiFmnGhERMIrJIW3G4U+kuLVMps4oru5exj1O9UUF8XxMuUAHQfHb98orMs3iNL
zlz+wnGyPRr8H+x4L2B55HfRlcnNN2Z5vI9Xpek4eSrRINIlqRODgJeaguEC/fyzrc5i7IKTg7MA
4UO3MBkHV18CtXu6ngmspkgKlR+qE3/x+zkbIK1ye7hEP5TMFz70/+1ewqIdXv5HvWIC2qJjH7Io
qrWug4+Pw9HfrC3buTMFHZMUSeLW2h9547+b0bUklhGErekMREOfc7qf+3cfYNwevYJECzq82qzC
3HAQ6uJ8Sspslk2jY6coQZLYCJ8MCXg5xVoK4R1j8zhDyesa6K4UGiWfJoBlyxLIJEGwzBWZs5ge
vLbEBnTZtgINRQY285ZSgR/fsZd7cOl7ks/S82/pf+NmRmcgIP9ZNX3HCl6Cf11t33cqUhFBBj74
02aWhOJuatSfBrmTJOKbX3VGhiJhBKmu/tfgWvGHrfZ/5IKCKcO+/eVOwdOrF4lzXXqid5BzLPYZ
ILNa1hteW8JDJSnOSQgsnmVeGTCckY4gBnvMs1ROmYluQkFW6Ncq5JuKTU57nemryyivJ+WzYN0A
mwhy8nu67gPME68EgscHLfUzYPvgr99o0nh90FUI7hxEq4uqd4UP3AZ+wJig/vku3J6wVVFQCtqU
P4sOOlfukn+u8b6gi1s1eenvPNNqIcmw82q+P6vny1aWKzXwHsxfDJO6jGhoN0qrgM0FuoiO9ErV
wGWSxmXgpj+dQ/7tBk4jz4InSHBHEx7Nnvth1iMB1qqksYL0z6Wjb9IzaUKe+bFDTmZrSRm37kRk
RQNdvqE2mvdcn1GkmQt36J6oPL4i463GXHa20e54msnMdqMZn3JhjuwfuxSaJFLHxX6XpTTMm4Aq
otRLA0KS+wqlEOkrdXP1cypQ0VBocDkxAzDKb09yGQxa/RwOjlzDUWWAHL9FrVW0IZQIBxkgpLxG
A6zyjMXVFUyNuhXg8ofYGqQVaIUB3uoIgVzZZ68V+0p96PL41VIdCThVBGEWeeftOzatkxgz6Y4K
5SYGLIGAW9bFD50T7kuNh3iK5nbhpCCi3dVVprvkB6un5fMAckV/2v3UdlH+5DLWwyE6oZj9mfTQ
X0DHbokgEU9cv3q1SrSi1jjIZSSSoYk4Z5K+vxbc20fC3FobQTTqfPdaFwIlvWeT0UOswEfn/Kbc
OyN5T0KFg7Tj4/zhd3SwK1YuatPlwg5pLGRURvqLx1TkXEIo2LeI8trQvPirm0rIhs7eykD4tdcA
o7SLosZwAMS4ZOJDwTtqfbXbtEPpRTASXxxpRaNo13DEntP5y8DFy/RPK2121FtdCIQ7L7uPaa4S
/aS0nVABi0tFJ2apS69J4TlyvXUuL1PhDA64IoHQ91bbBaH9EvX5oefne1jTT9LZfg95N36L6ZnD
3K3RNX5ARwPyKSkSfTvs4ePQDv6gFZzsqQX6kEPJQMuREHl3IKi2HIj+KAr51d9xHWKGwcFlXAGB
Rz6JgSXOcyN3iy9wwVaqs97YUZS2bGLOVQKgaLuIHFrCsppDlT5TTsTfFXl8h2+4o4l6cJ3K2S+p
Hol+lojmVyunXmKl2LL30IzBgHMfD8lUQPVBoJAcKdM4Fwt4PZYZOmryBGr0CoLPerxo9jQzyTaS
A0GVbcivDa5UYRnlr9dD+p+w6rr4rPX1EG8BwiaWTvgL8Xht7rjvUC6MDEF35BclQpU9iTtk+/cY
igogNxJ72YKKW+YfZFzqHF18KYTZ7YONZ2rDOGx6LjOG8Na693oMqUUnO3fpEsXgQmdXW00Uq0wt
e1HC7H/1rMow2c3V81Edw6SCEgZyadrfgRfX28OF4YVX1a6AOzW1PoNTq5fUcFWgQgQOqRXnUsxb
Xh0YJvLCsSA0tZgieWp6cAoJTuGRyreNcYGBHeGvknUGZtlskreTCmBCzXgQL+5CAaXnwQdpkZE7
suw700TEV0TZOjcz4AAsaejKDGZ1XIMWLg1bsN41688K/itdiBBfMWAPk0Mg/t3okaGuNpPTyJaS
P/YNdBIfyvZT8Tu3YQRBh9tKtoB6JzyVaJt1L+QN0X3VyFBwnvy+W49GlAjzDqbpuBbcsXlm8U4X
8U5P9zputYepATKOfmpeRrcdbT5BYgqgxwIdNOE5ydB8eCFtph+Z8F2JHjB8jGjAZQ78ZSNeS3t9
R/Oen/NFbQL0fqx4ps68WSgp7QCSW5q/011O57FX2H5vnxRI1spEAUFmgm3zWxAhvp5u1dZeWQw2
bzssVO6ApCveKnHnU/tkBb6/YinQ7yKEWTgjwNtvehMlvd2Fqfi1JpmN+1iPIe7AmwpSRR3cQNQB
wsSdntQCDgX+/F2lYHFWyKvuJ+b/BPpvFUiAdsGui34NRIVIMqY2cmvkAsdiw4ObakMlVdikwDIB
flbgcuGeMU+JWG7uIKabg3S7perORRlAHCp8gOXGQnd4eUfAequUkx91jz7efSCAZiZMsR38Sqcl
3MxVQhpMjs0JjJ/tla5C8OfT/HSNGdaN78Y7RltQg8X8UNLgs5RqAqFqzYW9/nFwuW+I9dG9PN1M
0vvA3uM4t8HuXOvutpZlp4EhTzEkunW1XXZh4C24Z7/fjtY9WQpi0chzMvLt6w18BeKGPhD1TVTs
cR/PPHRypcnbwt4pT+C6YgSeafhaG1Cf9dh3Xy16Puvkat6S3IgJOBrA2kuo/1o9gN+JGUHQ+myC
in6+tJQfF2wCH4T0E7ypk1Nxx0jyOydrroeZiLnEwfpypI7zoazlYbU7qmu1ACCkZKvQCJ0fx5n9
2UPDVccr0wii0iWkVHRuMjc/Ew1bvEUNCgMbzYWmxVoh9+DQcF3n3t9YkEuUv9wnZYHonFTLyunF
9BvDnrt2juctkcNFh48vm0HyFfTYyDvhm0UtumPQs5EL6DpfFfANIGqVcHmisqKVS/FTU6WwATdb
aJOrXj80KHRBuyGxkTTtKJp4xVioJ//1UNVc03SLrnz4qKwilxtkZwa2SBsBCw3q6GNxxHNYzrjg
ylB3m0ZROccernb8qSF7995o4pV9+/qVfxhGiqrUMJWH8MPDNHdhY2bSwer/cvXUw7zAFWYxDozW
yPMDnkpS7nwZtYzo0XxG9qdDGucQRaDD23dscAZaiyv1XB7jaaRp6vTyJyAJUqvISFYfgAsKqpM7
WbmDhOzkkdg3nQAZecipcGOgm+JTPkByZ4QFzIRkcsreQEVFm1pE0nxe+Zg0mcfZQ+JpkkquQXcG
I3y2lKLjRU6i5jendT3eaR+NtX9AxJJ0UsAJ8VFscf6yIxCP4JZgeX2V54kXdqwl1ZOUlPdz4Xmt
BcPvHc4ml94OHYcDF+wbqCjWAF4QNqNvkJoLanFAemwWsi6/54HXYtxCYa8knT6SM4jf6Esmugv2
DbYQZReX8vAg8+V/QoJIWMraPnnnOIeAoA4TWNp1HrvnIgSevVlH6s+j4QIBoCZbrW3HWOHNd6f3
t0wu/4uDankxsRyxELhWUrUb6IjEtPA+BOCvzSDMZNEwR9ClCk+0A8CaWqZXObkvMgMc6lAMxfYM
Sa7DfxP+rYC9RIikUdWH+8n8mTGQXEUeCVB2qgktL/5trGboYgNG49Tqdqw3vVNgxNWMbmKVW8i7
oTaA27h0v2jX4i/sWzteVDb1czjrZftjoe0lsS0kz21Up60ceUJIimYyI8BXnuxf61yoYscFRAw6
789yeui1V4mHQX19xVXP5U85l74c3EZsgXFLYsICL6oJJhj1sPZEVMNHW/6ksCov5UWCxkqzmW0k
FCxrWuy3WBgBiVdlPttaJFt3ihuIsftMdzIQOkhl+K5leTrdSeSBpXfADRu/LHKYlBwkgtDKgr8q
kZSjt8xMi+cApCcFX6e8p6d/mm/+dLxifrRBjC19cyX8brgbWUvor4OamaA+UwQW2DnNjJmxDV4B
RcTejPZMu8qfhNIgUUgNZdLd8+MBqSTC0dtdnISwdlxxULkCs4tBE8VLufg+OmwCylMZkkSNK2F/
heXC5CcyroNvY0T3Zupf/Ap+GieTMLQrfwqLO4IzBS5L1vXvBFFoI2e3V+PbAJNTMldVCZ8vO52Y
18k2qeZL+P0n8sCBxJm+vsgL842zq0mN4sSLDrVeFKRinY3iswRwmAQDDt61UhuN+IUJEmL2kg/p
gj3qoBZYq3nUtTceNJBDf2tPxNuHYZSkePBR+eCKMyMGx/ojUgdwFoqzsIO6Q6866UhNLRMH9LCt
qZyvVZpSGCvyIs19XH31Hr68SoarnEN2mRufV7JCcBxDLU9v+Fb4NBHH/nw0PmMIhekKuknIEFz1
CXx8RGlWkfNo/FOLnqv3TOaUuxukz37HG1wxZibfRNxZeHLq8AIeQwIDycpPg9QSf8kkagvot05r
hDTzzduvyEiZGmhc0id0bwlBfnemsNcN1lylMdXucw+IQ4pwNG1rXLag/XzRh3JckaLEaUxIdFNa
/uy4Fx4kfgJhjQY9fvh0qWB5pUeEp3l+B9fLaZT1RHPPu2VZ6Rzqgtmwg8/ZVeeJ9lofq4QtsXSI
KB9Iz98JbIwi1nIghMeWVxzZEFkhVkNfN82C1KpfY1lqQ3nIuKuSKlv88oubhzjlALpEjY/tZHz4
Arny4esVNC5gMwGMZJNZBylrHCwcyvtUb0P323H18UDQ3vRDPL1jEcNjHPpWTIZMq864tZiA12kB
6fPf6lHc+s5nk0xhOY9s8HWN5m4TrtkobMVI88nylQ35qR8LsTtVX7poXhOFdvXztlixzCRdtCgM
k1EkHzZLh8Hh+8tqOMvUKjc0LXo3NogULuHTFkwhKKsVQYOswNO6sNAG6xN/zvIlxT1kLqywWK//
cMlh2Aw0T1XOV9E25UT/xKsLGtjz+ZpPswi8E6iXePKDNM/anY/dxJPEsK3U/MgievX+9687S/gf
R88KWsYdoFdGNludpiV8bDZniaMZgqa5dhhotNCANUHszqRqbGgodB9SMAdDxdO/7SEx5x4EZw4z
RyYLl0wd/1xITjtct5ZGlMlzP7hu2GaBiHWcaUCzNusyz04WbN76RrQX28GD9bq4xt2F/ETUmY2Q
/Kq49MWq0dF4vMWNy6s3RkWCFFNQuGtgMbm3sNqjpW0slBC9Qx10Ets8Tsnwzwe09bWdXkSX4Imx
yiJGMTsF6r5DtFDZaH39Hg+N1bNrITjWSm2FTj+8OSCRTtK7dRurh1jEgX/athEUvXKgmoilSje7
66BUxs1OThzCCSyAuN+6hQYHGBK89iIQwlVKx3sFeq2GHEjZiU0pAjmboIWPbm1rEaFNsS6LvmHl
uzeQxxxzwF/1s9uNJvsRvH5GJuP0y5d81Purff3odJX5CUnGYbmsXNJYmYbtQkH5AkOQa07vEXA8
LCdLd9mJ7MdlOZimHKtbMlKzWfYdKfJ5Elnb0am1lfeLahONvoFhxnmVmwqAT1IT0KUZk+0sBMeM
02eEe3Rh7HfsPvlIdB/un7OPv5t1L/0GSvfj40DIcrikrR67wv6BID1dKQ3GNCyWEYO8iRmxPJ6x
JmqUh1ZvjKZ1+bvuqKszEYRnhK42Ei2m0iOt0oD5zpJHbDsAKbS1qwKdepk2i6UmEmea6LXhfeJ7
z8hRjQF/DTgb0hqG1XJLEZPsDzzjIj4bFfUFoQ2wg5hhCfT4wvTQSEQY4JpxlpMGg1u7lKDpNSKV
pisNOO4e1nfP29uk48+xOWLhgqKVWtrpQe/kAzbOrSq/u913WwVe3Dogqf7vMJ9zwjTnYWClpmIU
H55qLS5RP1dwl1tEd18feZ4aomRm66EXkgx3I7eJFTqU283vn6Ka6xJjMJXK6rLehgkFYjEFGinX
JocM0iqGowF0Exyi4z9Kcj6R3U6HiMYDMryrDdZoB9s6v26R77ZlRBVnZhfLRxxRtWdhY0vAgg6E
MTwG0p20DXw24h8BMZKigVDqu1OygFsSGGijYQsnCM0PeW6M0GwNF3a9NCc6nsfoaR5YoQ0hHjT1
ARc0cb2cEjpb93GhlBM2iP0ZAoOoNimSgmsyhwwI0QOF9/urGkJ2GOJ8Y0r3mU0jDA+8n6Q/9K6E
idkOZAOK7E0mFHwWTUhPp3k5orDT8s25CM3n5RBi4daZlEdx7wGzMmo9j+mupf42yAWMpq8QYolv
JyvFymbOWTrtpSQ+npsOkmvkHZT8OGkYyj1ZNIEZzlD79U3O9/1gdMMLNGfcb5BMmHaAlQjnfY7K
tmYQD8e9bC/v7jqs9gd3rLg9IuqMtKm8M/KYw+a0XZNeur+VcjJZUbFN3TS0s2kqJDmhziPTdEYm
4T0NK2yLleCL+PjwwPn75j1CEUW3NxlIykz80RH2ghbppEOnfcbs55Rd1tPMhnMYBJp8EnZeg3lm
4GdyQVK1d9kt6Fyr/l0BPLDNvVdb0aSLegpeWVAX5TQ/DpyUbavBir0PJs2Lj8WTqajZ6OUAJ9lU
Q4ZDCyHLYpNcD7YQLYVWRYSwUX3iYSmYGzeKCzymxDI19+MNAiAsoM6exJhhA04mZP0P71hFYfvh
O0EFAXgt52O7jvr12909zeY6i6dwZUO70oAiqzcsuJYuzCfFhs8bwh6v6OElxGrp3llU+sKrDlMP
HmzBbgZjByIWqUbzMa5ouoOvmbrfiLJNa9w0yZ45m5WeWoqwJhdYhb3Y/5kL8iN7MTBNcgTZAta/
NJhWqXkozXo09a9stSETesCZgWE4eVMYwYDZ6WDJI8t5YoOz9B4zNntAfqKxVzos38TzKNux5Pm3
0D1mt3ORSDbZveIm2Pk36bDzGFKBjQFazSEfX0GIRY/wI8fyL8clxMD6gSan0N4L24P+2tAB9YcT
6i/or2znSaLCp3sPWqlUJo2iV8Ntz0aXqGjZyti/0iAkzWDSVRjQ0kINX+YSVx7/rW5mXmP1FYfs
ptPk3i1R6AkKDr4mhAyRnNR7A4A6ShEfNLjyb6e/4BWTJOxF45rFjUWVHEZbr2ZLR9zyy8NufuKd
z3wDe0MYgYHc9ucFNTSGhZ0sI157PLL8cL2ci9TB+nGZODFWq5NBdU4gzt3GfnQC4D19ohuyBg0c
Fo7Is/l2qQox2Yw2hVvC2tQrAJjfXwiOBUevpWp6tr4nKlj0CTXX59KK8f4CjFggzo0GKzt+f5ob
wGjJfOdkxfIUEMlw3Js2tkyiNZhnAibh0JzsiABfXlGqbYOwUzgJ6tM/tQvfaxih6IEWPJSBhdN6
/IsAKOswblNEeTzwJD28+SqtAwqc68Gf6rqoMYoJz8wCwXYWTHdKA3g2f4V8P0gg5v8/tpJ6CLHl
7ni5JzuXIhgam7JyKH5Y+Lf8sO+3ib2i9FCGVSCh6ZbJNRAmMkmg/of0Z9ITNLmDEzJ33mHlG727
lkc4St58lN7zjVLQEUuKf7aK83fxm2F7/MHTMzLQz/APo62Eb9f9bOGB3SuOOTDt+SZPKg9Lfi11
vN0m/DwhmBSFUsFFBOK6KZ3vuq5qWl0ddpVxdoK44NUvKX1/pqMZpv4wh+0nsLynPPGdRRPL3L3d
rGtDby2wfM8YleFCuQx31i41ZWN0OYIafDPrYnyNj/s/ypnaRjSi4QfdfSfxo3N6mwJyF193MvDx
X/GkicFQpBC0U3WSB6YOQ5MG8SKL6FGqF1pMskgp4XV6e7VoFFPJgOwEPdrfz0NtcihQ5JXGX+uy
pSeUYlntIB+xC5x604oQykVKUOqkBpH24/I2CWiSed6owZrnhQQH74al1DYnf/ikqzQkLjSsbiPF
M03Ur2lxXHz7NsSGjTy6oZ1Ehvi1zHdN38fHSyiehH92RvqH588AcejT20Hax98GAHa95vqnZJNX
2hZaBgM/dUfEE5enyVNwv+zCUZJCwA43m8XPZLT5no6IzpngAait7sBzIPSHnVQkeTpWZcnNBRqv
voxWZg8XI7PtLM4fNCVFwhvPxeHT3aoVPgQUp7xWWvFrS5PZHaxX5BJDtdb1GlisWiFcvzWzk7cY
1t7xTfICnlM7bDO5vlXSgxkAh+1DPcPs9CKFfgUKESAky/JZqAczw/VTS92k6QWhDx2w4AJVoDlo
y0/WpzGfJ/z7AD6NxUXZH/UEpu1gVeNShwKDfSEnyFEwdmmX+16FuCFjkv07AsoCZdPsUak7ridc
LYDF8liBFAikLbvOEUr/yY1qpT2mHfXL3EqiE4EF1NkxLxRPnmgzj0NDGy4m4plasxhQ9TPjE2ku
ZDn+BjVY1De3zXpW0mNhjiotTWT0Tfm17CS/45KkeeeBfjskWKxGqcjBH7Lzyg+A1B+kgg+FRiwv
+LS1UvF5WtPJPjWO/DjkeZjH5QHGqoeFMAzZP8ArsBrdUnELj+ejjJOv4ffYQdxKpHK49RtUKqAl
ZArlnuSLY88SHd6iefoGXtHDj1KwzsWXJesSJr7rsVcaSv8qseyM/33EWnYzAh44bLITPZR5iSwI
/wnps8+U1qHefPbxxHFvfmjvH1D7YIIvFj3z45cFICLcSfB/Meh4iFu9tWXzMrnORn7wqlo/WquO
D60Ercd7eFEZSSuRkPMkZU/mVi3l8TCxftLv3SyuKK2ovgie6VVv8Xt1TuFNC5pDeINf+TkaqTwe
pJSnjao5QXn+QuGW+Y3QZ4q2DDpQAPCFim2uPss9Y1Phuj/ZI4vEPSbQ/V/7wP7pNQV1TmTqqyEu
baaW/wQsKdmD5U9W+XIXEAGYAwMLTH/ia+EbZ8dgd2C1ibJWkcaz6mPk5ITEPYBAX1ZI8GK6IeGE
JvE2IZUaQ7jrUxMJAKfdmm+4+08GJD9c2x1ma12mXlz1OSzSiCptvno1LD+pqnJisdgdpfOrL4W8
mfgSfSQQtBP7aWvWfh//BEtb2SQixnMRgY3hA9J4PI+DB9J0ldX+8cg7B586EoCiU0+NH04CqSDS
Hhib633Q4kZJPNrdxzsAVXAp28xQkclRn2FPEw/iyVjmErj5AgXoAeCUIfn0t+yiLDg2ZX2KxOfJ
1RbWO9jWWfN+Tt6S+R8X7tSDLPvL/nagFESoSOJszhhRKn4dktfKQD20/S37a9u8N+K6ZV5uCloi
UnQU7bsdoD5dg55POmATk2lcEXg2LRCqngmhQJ7eaSDAzc06q4h3lgdy2lNNLfzX/DcOY2nVvcwy
Q0oIS6pjIvS4mebvdgRJTscRI0HFszIy6xzgIbDbH0kZhundX9PRWmgjn/WhAGtqEuiTO+etHRRX
bKUrllOQit5osnUxVdN6oBAKjuPkVOJNvO33GPwQ6t0ABym4qIRTMHcttECJxoUwHicisy6znplc
UWz+EJNQmvmj4vti+2quYqRxoR3BlYDFDS9hfP6Z155073iG40WMB/mdVO2QN0JAZZGApA8AA5k1
wXmrL2Da9nyZhQfK/1EJRNNxgijzCHwfa32v64Aks6OX3IE1jgzwBkfY1vCcDayLc14ZObUd5awT
wZqs/PxagfXKh0Nre1TUUY7yyCA1DEA8MsG/pENLM/DNB/ADrVbjDOz2WSXfuwgG0pbK70HqnfcQ
af2flrJHgkhpHJL+5DurI6ShzEC/6Hf/l2Yo/SAdhbhvSBIoGUUseVveq2YcLvB+BflfRThmQCQv
CMtxqIHhUl/BqUv2q+qFy9QSmazX7OGyGxBlwM7WiJ1tWt/wZSg4xC2cfuJXNP2U/5keZR1UVKiw
hFDIJeEmMMecFKSu2dWzS3B5dKxne2GeDC+rmZgQ3OkzzUbxEUNF+T1aK5SBdNONe4cL0xTKuHfz
jcFj6K5uc3YNMQFa6jzc8Z1UBrfB2eCJBEl2CzP1CDi2y6M7HmXCWPDfHObsY8iwCl1jA2LoH62/
DvkesIjMmuvuFFsYJ//+4mO+0QpGaenHNLDHLcQguhPRsW0PPbTI/VA9igYzhtl4k1kYwepwHygb
5wPskvzaS/Jwwve8aVjUZ6WqyqWOoCKIXb8bEJHl/C1IXEbXIun972I0r8tBjDeIfevb3YQ2qMiS
rbBOs5KLl4Wj6pnbP4PEX07Ep/RKdZD7ohqlbaGi9c64Aqvr2iekOYr/PjAhKlCbXS/+uGMv8/F0
9yDCEvpaj9A4Ru0qCmI0BCskPWD3GhH5vkz5YVL80DSUyhYDE9PDQDExiVNCrSymkTnzZOeCWi1P
k7qd3CL9bRu6k5d8QLfEDNqUNCw2gHR5t7nUl7aTHKveN+55NHMDgfgsXaj30d3wJwTm/enuGMcy
FO895kNvRn3Wx7103U2wzfbR2Hq/H6o3LDbwj27sDG7kSukimMPC9xsYhZGZ2nH7SHPEY1YzEs8K
OnZ6U7Km3qkhggSVauZQRwzxRAk1JWNijpz1JnIYUEPAPrRTV5iR83jPnt7ChfSYAcExuti0DVt2
4YvLNKy08ffI0ovjd9REGOo4W7aQ1tYs7bH2oqYEZbNK3j0OfoIOABNvGrQUv9LZ3NK6hjYQ5EHm
9JKoX89mOuvk51Y6ShlGFi0IeOdfEebh/hNufR6y+t/Gfz1BsI6D21jzli93XG20ONaxZvkrWQFi
gIwyQ2iN1P1Ql939NhdwzvHz3EUyfwnIA/ESFBfuZG/LUWLA7D5HDa2upXeAAsqqtT35o9kVObE7
GalMkaodeC5H28UtV3+pyh0HS5s3H2UnN/hkXiFT/tx5wAnu/wIPOEWGf58NuEGSeppR2xZZE1cX
kb1lBHgRohH3YbE4ouluL+zgxi5gHlobeb8HPUa24loFgK9U9aOv/EI8gNFoy9gTE+3zMf20zpBG
8pPXt1ZoG+2lQYLUfiSj+FQs6wi3/e382RTM2ShQ47r8y2bvEonPSw1g/7IZIsgqHkOqxbDm1843
Vxyd/sERz+15HMKTucs8ptQH5nmo7t5ieMCt7r/Z/Wor15cCcpDS1+/Gj8ZDL6Q+2SHvil575eWi
91cdRsx2RKpTDdwK6nFD4ozWFdX/DnwiKviC+WnCQJGIdDFtCtmqUl85GseBRzc+6KDD5oofsDn7
XGJ/hn79oLOzIf8p5Y1Vbnire72eTLUvYfpc1gi1WyZ5LEyvIdkT4oYH1O+p+3T0KblVAbaxS5Am
jV+/ikL89l1g+Jik0y7jBVpbTF1KF6zNKJGr4My710Lm6C3MVOPIOBx5UYlGnNLX/43mL339KUI5
MAcG30xq6Kc/CpifXgCOtRy7GfGZf7anzNrJ5HMqZfM+14GeULXpbriPryDs+6zbbbxRZb43cXpC
+SVWYJZoVo52auJlf+Llt/yLWRTGjmgOM5j9vEyyXw/aivRqXRZTeCRtK//13nmX+Uw0AhfH1kDG
fhcJScy3uHEaTYnIzZTF5Yg9zCdZy+MdWzD+R+o/IcHz7kFe66HmnrimoxusiXTkVVJ6IRzO3MZy
RlNqBRPwV9H9Or7q2QBimI8kX2KwwnyaaIdTeACd0dK9bLr3kuaMs/+pCcdCOUoiUcuxD5pAcsJ4
HRTQxsRgz/Y/0xqebFKML2zo2zThmCC2YV8zWZ3X2FIx2MFf/GpbmVc7dk03871t7rbltW403U3m
5EIwg0oimnYzkl9udVFd2mFljGRLjli6KpvN1LE0ClnBjWbbbwWgDmvaMIeQnyZK/dt/gB4tvmc4
TkTH2pk6Ro5yEDS42oVflL4jGszrn3jT0P7QdvcTrE3C3ZyALEYTil+1jjazWxYp6lG6VuMLZVaP
A6NiGBUGD7AVjNJozmM2utWAzcX5RFJYurDz3ImqWWPCj0tMfACdHGU/ewUZjssYAfKn0tZR9eOx
Y/AITeNOR3BdM9YUlEXeXpcI7P6cdN0UL+bY6SVrrxWMKe9YoxrTrqXtMe7QhQQlA/drmlmvlqVP
xVtG2my+U7k3EwuuXFipLg9Q0BQ6AfhxR/iCWn0VyE3poSQgmbkAJ1t1liNlbwDc7ZTdmL6vsxBP
6TArIfQ8SPcaxadFzDXscx9omwTOxVoluM9JX87aIfqO48vgQhSRbYMmwQt/D7uOm0RTtN53+QOF
a0o51oLX0sCBmwLtL1Sq43M8879MjfS1LM0OrYP9g/AVemmwkSZz5h7o1RUtryqYPYwgIkVN+J1g
RP9OqMErGv6EHtt09DLqwfYWeGXsEQfUUzdk6lSeMc9YSwDF1zO/0yOt+A+SmVlMb8JS/6fVShir
3UBmvLWHyENOj5ObbkH3vKKIXxXXH+ry9y17piE1ONhqY4eP8qY0Vipk4w6j5ihYHXn2Aveq4eYZ
L4bHLf+396vIVNZXhbAVWmNOjQrHfKilK3zRIwfEzE67A52WG3LrjagkS5LFPvU2L7kzgsD1WZPC
BVE61+2SKtGm2Ozgpo78WK2KwMLfqZET/fDoci6dbnmY4sCXNQiBZG1kJackFbVSE+I1IrO7tExs
kwcJ9Kpla+kfF1szpwf844GkRWWMkzLtV6MHG5op9Ne//tZcXlxc8OeFrkV19mv4y+Y7xDJl/A8E
1PjEJDKCqtuiHJoV3cdlyTtPoPQkWoVukVKeyQ4JsMybrTV+8I5tKFAxYbcpAR7bqeGQDgk2x800
50hdrbx7Zcr6v6RhkHDjiKiALfOZn7KL/HbFGTIMG67hoYOK2RfuyufvEA1YazsFnzkllyivjJ8U
aihcKiVmy6qnrgz+8pK2oEmn9mTwH2tkTvdn/X75NHmu6uZFEWGA6BGpX2teIqjPRGt0tV7w/W0O
OOt2CaCllryT3ElcLqhr2Ojvqylxa6f6MYm2j4uDqoL7adXgoNUt6BZclOwOiABsXLnFf2bMOcqG
b4loRMcD5+Ubv7kHtEWzULI0Ps1hBEdW22eglixoJcDM9vIfsChuhv0FEYDGOhd1CO4LXZPj8AbE
T+f2MfajbL5TDOp/FY/ytUtdregZkPpotMl8QyuplPVTCDb1+A182tXjmSdCTJa9M3mojFxylihv
jEBjCuMZWK9MIrIYJ4ITQd6coFqYoB3qS8BXYIwd7S0lHC0n6niihYA2salUT7L4SFSIfm82++6B
ZSM5xqyseIQko7IieVHZgAVRpRhFESE5kL9ZnHtrWMPsOcBdiAwjFZU04+63E3/3uJ69WJh2GEys
JtI5BOr92jJHWEp4LIkH1k6tWTkc/mizaJxdmMApYVLLKKPyN6GqZqSxRu9S7ZsLjy56EFLRYvC4
wEvwtArIE49XtnWWXl733GkRR1i1ETj2DBmqHo3NONqUIPoq/X+kdL95mlsDKoUvnM5Qq/vwdi3Y
ZkXPEbpuFW6PzsSK2sVnGHUljZQPaOleYfC/WW2uSi06Vt8ix2zaMwt5rmjB315Ogc4RQKP6GaUv
7DLYLvImWRKTVRWU8XSI7Cdt//spEIqxYCSNYbFxnxI7Bep3mAZ2x4csxkuqWtFmTrpeQ7iEsla2
+GjsRsMLPF+rjl8k080AEsdMX/aCZmfH/9Ha0utMR8jI3oQACK/6yZlDwFrCRrBUB4xjC0dimNMU
iuDuL+M4shcNVZ4BxOBVrA3HpN2SK7RIyWPLQzJC2IZmaK77eN6m6c1SZwZrAevvxP0DsBa8+Yzp
rz6aSSO7PtY8d2xmqPT35ZsDwoKcdkwnpJWlJN4P+HL7YRPVA5kVO0nyB8yyEfKMCsCmWtc1nlxa
RrkWWjaeMdrZ7NTaFt4CcMqesSsdIZaZT+1R5hCRxMw+GLRuGtbq1bs6bRqMVV3kNdiaPyX1iyzd
BYlJBUMgp4HrrrHLzx2KNIb36I6omPeKZGEpLEW/kOv6mhXVhd9AJhdJ2EKVq0awdwD/3FPcganG
bP+27XvPTqbjUaZA2Zqoc+oN2wh4oHkQp53bYbJZRCBR+Pj7Z7IxFxFLQ5LYtTIIdT9xCVVvfsGu
Vc+qzTazKj9XAnKAdvVam8knHFy7HlJfdKPHevI/PPOtd8q3a1smzYlliTbCOAFYs5QmXTgSEJcR
I/0WSv67hIM+XtfO7NYS3EaoUeAmTBD+fvXUUNVZ16V6V1l7uPYpCxFoRULI67LaFzseDZoRqrpQ
S1elJESR7MDxVlzMEzyHs1U4uzpRs5tdSXB4F94OKi21iX4Zp7vJ1Hs/HhHBjSlB7EvLYjK2hzri
1qsijH4myREDYLGQi7fq/KqAS2nakskp8rhIM52Qfa2uEbweGCJ3MKL7jGrjraqH2NA3RRRQfn51
IOi5DLyyRpWvznpaqfG+MCEPyy9GTgMJ60TBSYEUJAbkCOMqOBOukzmKpaXGUQ72S92OUVrmjN5y
S5D9/VOGLyAAZXxEM0YMevRHTjM/jdb106sjAJbOAXZuwXrZKUF4t8ZEkM0odfzuZBxkuokXl1bW
PBMHCXdaUKEvnznsMdHKQTBsB9htbkKMGqC+C+DspHmzR0eXdnyBDeiaVHe3uLIfOmuixzJeT4fX
He8NREdO2I0EIKtB6Gws/5dh+CTBA9hLjYTnOEKI9MxwdZhS0tWlabg7zIQgvCqU1Vvstr1ICIXu
uBbl/984Yg4z4ElTYWP+0omghWTZ86FaY6F74sSTEF+O8+24PGmF67lLwr0m6tb7AOjDGA6IKfpF
ldG4oOTfUg+KeIVA87bndffKB5sDT/fVrcrWijdpVV8VCyLCtpvBikYw+WIxpnkW0t93Ibl9OEYu
GFNcqJoC3eLEsuELuFZNm1ZWXkgFA4keMVDKH/vsE3bG3IBXrdfs2XOwOSm5BO3zlvxBNGtPlt3B
8W9R5d3NdriKwE00zcePVWE2klS5hXQ0iQhGqsY6n9skhrb7foZDv7pR0AJ96yMCGORDNzCRt/Tb
+OoY1ffdmH/0CL4e6ELTHTWlz/mDyK/N0uz95Sp6VDUkGa/kR/bVDdUsZ0HpwOoBjTnjln/sKa05
Ohl3D2PkSO8OTf1NIeWIQNNtQmreqbMAOTQ8uxNdJUl9XGhKnlFPWvqWI1Ao7SvK1LKjSaMj6oRD
3S8uE/al6oSypHHfRATRO7oGoJv/cNEu5qdJd97usGwoJnR7J8gGcEUie/zQlLQlNNt3JgFIWTib
v4syhxzZ3g3upbIABlCh72NQh0inGdMb3bNMwfjO/uXyqVC0abh5Qx1OVW2cBokWBwK2gHfSBwpj
aBT0s/D3H0va+2SqhX2kCBWlGUxQKylqhuRovO/uWr2MqM7Ss0oQvFs8wqn6w40ga6h9oJMlhVtI
rO/uVT4SYB2AbTDbDyVdKIakskcKIhvojLBgP0lsYhroAdVvdSmX2iBPu36tGuH+QHlAA4C/PcFu
6pNWNgg+Wcm3dB/PyOU3x5DiFJ4TMYUp4Me5T2KRhSrW6u9Jehudiu9QtBvsKfG+SICjS7pxB2sq
W2OsSeZaIWQeeLmBAVNGPFcR8lIz0jCsNjMXvjV4FhoBxo8+4oL9WxIONZ9H63MNCfUsaTE8wmZX
+fMMleVubrd+7/Rg++p3p63FAYxvn2JTxta9jtQ9scQvq4Ku9X3iaMEPaHDIHvLZtqkLUESi901+
aWo+ALH1HOKvJdQnZFHUh7PjmCqThCJ7kAMs+kyDGNVHMogdj9R5ViOQKYSLsHECnURc7+Vm5iT5
0TmmNTJ0t2HQ6XpfAl/waGS5Fh9RLcGrVB4CMNDR7hII+6dNOM4jM/wmuLhMjt/wjuDWjt/6oezL
9zlMP93eSR+Iou74bqhGTXoLyp4IxETXdawK89fU5tGTtYL4JmadLtVSIfUYAOFBJLeNemgzmjzW
ks6YHfdl/2zFeTNZzTX+FK7XYyP3c9Nuf1nBRRBWSS7jrOtnZsQevh8FBad/DJTep9j++mBhaIJq
e7Bgpreo5klNORQxEwg0Hdxf/KoNL9fs851sXzy66JZumpIwoXD1VH/sKskuRImdUqHNT47LWROP
wuE6K5TAr47m5eCrpmAjw/m6IQ94ZroUKodIXBmfUj/nVhOkGUOI6N1VFQzS5wQC96ZNlEpeEev2
8YgKWpqJjmiB7gooZ3waHzIs2PsAsnm55X0jaL2Qzv+Mw0/KE64t72DYiauYSRNPNmD6lbua2sNS
8tMYMhGT3aqhdhnsWYD6tMULMp52K64R3zfxugfF9Uq/C3H+NILOBhv58ZSDF/Wmvll3Idyvpudg
/MRcwJB0eqUqN6Pp3bWdoIkTk4UCpkkrtNNlRa+UN+OP+vxJi0g2XA5LsSsI1PFG/y6YyYbXCtCO
iTLvVN/52h6GcD2+Bbb8jnSHah1odu5DSlzXbo6GvaPauvQAbEBeOamdzLtLR/5dA5yVGOmFwuVj
qIA85XVwTlMH+Oz5uU38PWBMPVNaJPwQIbow+LkYp/P/Z68gpcfZpNn4VSnQYrrGKa997ZkB0m4r
Gb1bFtQ2SNBu6b5q8Q0Wo4q3XjuL9/Hr2jOvvRECNMf9QJ/PyvgCMcUU8HbFXp3uiKF3O/bN4wFw
NJSPIRJyKqjyhsym3F/kT0BwC2Hj3cNicUQnR0a5KnEurKLpkzxoxlo5WA3lGKKDQ9/jyqPFcnCx
+7Zn4u0LFDUwrXhhVqvrRYF6jypN7iQg2/qVcKW6MLT2M9JdSiW7kQEume9g5W/rXKB4SYs7zB0w
noJbviarNFhQYkI9vWpD2NO84S+i6RR9VLOiDG9uSxkuhCIb/vU0PNVPxZNmp29UkdCrTI4TAdjO
6ZGk18/3TVM4aVoP+e8c0Nbvc/7c87RsG4QDBgXZ/z7+lB/N3FHzKF19hNQhYj0d1QTmeaZAsapm
Ow2R0ViF3MNdj0c4GFesLLREz2bK0ImcOzDrRlICzieMtMi9DswQL26EZAy4YWEiDuPmPUnEkxz4
Jk5A1WGYBYCdieWkBZKjtHE4ud5ak1zPjFwOWGJ3oaWchb6nAlsUgoAtimb6XwIrcdpDDxhQzywh
HwntkWGgf2AhZljvERZ6pOGUgu5G9l964soJlgRxIo4xmu4ZGU1iexFopOqhwCC9mn9nMwvtMaS4
RVbWjGcgp8Ql1jQ7hXfl7qEh3r1Y4/cVi07Wwm7+7Vdssw+8m0wovC8A8FGQHKhagpK3Psf/v02a
s/tExJ356VthFaF6aOEb781bjIRWxQzfgIguQnqlTfXkviDkiP9yvR6zaz6FvOZXZCJWbCi8NM1C
6PYJWi2B2PcCXJ2vl2+ogjotI1IY7kxnD/K8KV7GAYP1J7PPWdQYyQFtDeKXEBkUZg3pMWxhOv4Z
/0xt9yLvu2i8FQSdsqszF5Y1nMRoCE+xfpZYH3n2LQOZktgya4AJfHMHYmDjcui2BcahMDyVcIfB
S24/k4jk5R3k+kF7xaBLZoV/ENIuvYx7l3EvU942cTisRK5WuIih4k6amPVE4PrKz063Yy3MDjbt
x+dXZOhK+w+MDcr5OQ7TZaABJdL1r++x3ivpCKGCGetsarImNRnRXKU07n/g9iyFL00svc14EwYY
ttXRZCtSzUsD296Emz1K6Z0oJ9C8ZmWVrbjmy7FLyYM6VdGPCaBJFge5sIpg8CfoZOHGyfBv1Kgq
sKuHK/jaxj36onM7hffEOkpcqf7wFlpIHbhesBBqErKNlFd+5NrChcWDWOo/2FsYxKrQdr6iGNVj
8lpiahkrYOssKV9rVg7JmF0mjM01x9UbjQz3EpT0GKlSbI3nOc2AXa5ESXEifl4jeNb1IJh1FRdf
IbAU3PTKgzqemCdKUQ3SBgr006ohnDVYiVSNKYAtz9cGiIlUpPY7tslV057KNuC5Jl0noWIIlB9Q
UqnhrP34N7YE4tDlDc4WgXfmGT+4T9f7kZBlA2NQQr9ddfbNBAbSFiwzGtU+J8CGrAybFYWAANMp
uGzp+gGOhKU8f2s1hS0Wd5Gbl3Lx+JjQeb8tzfPoAg23VFvKi3FHJYlhpuJ6Iv4lfg9pXDjfcYfZ
04/Kv7X5VJ104F9n7r057buWCLMkgHvaePShzClGsFZSd9omNtCxuvV9023nHEUnFmg5ooQDlBwa
KZvxUNjZ4dqTnAzCWYLDMGg5UD6vVB6pSQKnY+nKWcSE0NYIRvH+bJJ7dD2j8UsmFhuZUmw3UyEF
D3MkiuPBHKnYty4jdpIkEyV8z7hQOWQJ+PI8adBrBjlZ2AyPeE8BEjIfG6Hhuk4Dm7kgMPoPhlvM
YvtBuBd7CQSNfRrR9jhMK5Khl4N4gBenwKemejXVHJTZH6EvUYm4Nvlc/I66fRqO0c1sIo2Zm6gE
uIgNfAWI87wUk5eCIJe28jYZJ9U5pLgjmgLur0AmmP5yFDb3jSYB13wKeS/kzbQZObq7IWvAcJxi
rXjRY/1U3D57t6B96Lc5IAxCHD3keFcpValPbAF3yekieIq5CfVHEp9h/pYutHzYcIP7MUpbeE0w
+dr0T/2UtV4lMf1h8x0t/D9CPP4+HrwF8XfVCavHngSe89kJqDgJSGQn/MLCyCwOYjLBLifsPErE
UNd0uYcRKIHDHtcupDWP7WyQOjUGkwItEnzZ82mUSO2d01AEcTwq01rZORed7a2psMcEGy/iQR2P
jzAEBjlSF7R9ZdGNptrYvqYQ6w7X1v/V1uwhh9EAZ96oeZQGmmbHVn5AVpQMhDOYZzmjEXIdCRho
49uMfdggYUP3W85hKjmKrKGOHueIhGD2Fgc6Fcy9i3ZHcoaCMp8Oc9YoHSxr90zOTBrzXXZppK3r
ykvIiRRIXLggxTapeaZWpW7XG2U+F7Q92JBaX3BynTdUIiXs+vp40oLQ+8MaM92yZOMMyABmnv8J
6bSXjwYmwLAFA+gett8zDCkqMImTImb+GVYYUhd8Q9/iT1nxvmm+iBkXcOpYYU4PhpmiCnRjX64l
31mLJAyOWpnAO1snc+BvsGEIvtfB0Q8UJdD4GyB+boSXkGc5586PXJqU1/aVbs4p+NUsWkORD/Pc
YmfNtHwIR5yca8CaOnSoKDHW1I1xk+OePl4v1IRIXIxgBaSIsYfb9yzYPnFcTB7xwN+Y82tPaxbE
BIK1BDEXj1cBUea2SE8fazoG0AanSGpEz+vWN502/keo44PF5sMPdZBFovw1wdYQ8g/SL0Xryg4C
M2HQ3OqzrPYdUqcGa3UUWGaZSBqBmK9PIUosAXHEDePc56GO0vp/0tL3pyXJkaWw3/xUnCAqed/S
LGNCbB0v4eSJWLA/A0bRLpJ7YIj0YOgYLxNWBoewgSgpLwIbOfhviqgbmlPn0ZbPU09lsRNZNxTD
zNTPhlc2l3bByuUlhE8ATYpvPVGscMbZYybbfrC1ZyLABTxQvh8zqKPRP+t2wNkQxxTFHXvzOMpJ
Jb0QpfCgPTh/6WvWYSEuVgHF6ordXJuSKaYSTxeHuSC1pj8Ld1AgVFnGV52YRLQBYzS7KUNinB2x
UxLIxgn8AgfAqC1YiWAtOKHbO4+VLsP9Tvda/OQ/dSQI3i0c7QCBt7e5FiGNo6cqtaA5u3bMxjWM
B8CYN63OpimEf2ZUmuRnV3v9ddwEirjFqU280GtFuniZzT/NDLWOZQp7MVcO05YxRLRb1eHJCkFp
O2iEaF80Q9rn53vDUgMy/KWQXYccuHhFjxhuWEkud5DJnscuJmoqyNcxWbl26PclMVHVKF2neQOj
Nl8l1vSOQYYeIZkJPTiPx5pEHbUfi03IBDHZin7n5BaILnG8Y6QzsNo6DvBg6rP580HAI0fTkSlR
9VtBPwM+6TCcer6EAE2HQ8I9EWvNEKKYlHtAX+2hwAZ15m+F7ZZiAV6FhqDQovZd2hZSM1ZXT6gK
9bOr4DNoQULVJ5ntyruk2CEwwHLizRydClYZFQUu7ZW6QgRGUOii9cSHFgngEdj03CClzP5dCAuN
R3QbJc9y1IKsuzaKtSnu9xcRDb3e/NRWQDg+r2rhZ+tegS5EJkET344ZL5TEhxYTrcuov0VKB29r
k+EhgaREF8nQxYf1cA/AbPvTpDGAJJCLRN6NwQ5s0Cb7XLOcZ6r7c2M4WX/lYd/tuNt/1m2Jvc+i
L8oywxDwdSO/mta2ROZMZQknctdBf3JTuObEMqCHM8zfWckCuTGFP2UON9/r03U9+bETexnf34jk
+pcjOScEKz5Lpt/m+l9PeV0wbAWTR3997eV2Xvec562/jyMThlGvd/IBCan5W/rcgrEEng8dDBR6
W3d/75gMx+kMdCcDhXDNPlpBvV227UMVCU97FCcVMM1SmfRrhJnePk8TU2PITMcEmFDpuATfFUfW
aTvvFbKtwLuRkFxWjDjwptC9xVWX1pf3zPiPSAxC5pWJnDHY6/702P5jAGk+h0zCTgmtxfmETqpT
SHH/XrjlF6yqM4nphrHST/4ELbxYuvctz6mxlYiOJb+pj4CX3IfPT9N+xjzQQzGPybTU4X0PceFA
M9bmjYeZsevoIOUj/CnLVWxLMEcx1l9sht1tYGKkG/UsxlsNbYBSOAuwdY7JomaWrfGXWijUh6Vg
85ECPoh+5bxJspQMYuxGCSh8Twwr9uwDlzWo1yQQufOvxpj1N4hrtZrg2ZeNK5TvNHgEXruu3qHV
nuzLz2fQObRMr0U2i677uEJx675OLu3ewW/onrThjsjtsU9IlnPt1EnzXDL9lw0m1K9IhtjfS+GM
v+w8wLokkqOYQRMrHdTZAN+rMRYgWG8FkWX2eUuhfP9YcgdILTGvIsnkgSv6ePmAZqpih/GyETgd
q2JciRzwbnVytfWewXiIsR7H4dDuRZPhVItrJ/vPnaaATRm9YPkP+Yf9osKSpMggfyL2PvaMiaxp
fahz1xS2QfZ+fmMnWwOyMLiktc2NeWEItC/fi2sWIaaxfsrLOaTke9T+CgSup/Ecp1EGLZQxIDhc
JaIr6tn6ntypGYTnvtlh2YmL8Z3OZHkiRJQDwSlMzyhKtKIgu3JDKZ+tmvD1Y9SHC9OziKzTJbQf
R+sGpfCt1HA1W40DMC7E6EBu49nc0eH3ofxfAfHVd3RZ7MVXeSXTb4ted9rGNZ89BzjtWLN8yVsl
THp8o5kbCn4KfTPeyswmVoxwTwfYb0RzfcVWEITk4YhIb1whfo4yfdkc6kwtFVv5tyfVRFN+Gw7x
U6T1q9hbfQ9D1l/LmTI1UkG60O05LF1ImFiA+TAOPMRyhcCSg6jQgGmSxnegstnTixZaPAJFpwsm
ai/szlqSIu91z0+Y1gHm1so7dSqeRaSnORWH5V197hBKjM6U7WoW5ZKLadIzaNv039PlxiopHxZq
x1X9fcfjzbfwbjmaT1V3Thz0myTs7CAqNOZEkZNK4Vx7FpdVKDkJnePMBXbABfSKVfUlDoVwYIdl
HHtMb4ALI/Wk4JGekQ3dxwWAJjWCu1FWQVckFdEHGmC2sJF1voGwj1I6tTCwBdMHUIUq1dBe3srf
jh8uhe2PFR9h0y5nLkeRLG56AEgl68uHGd0pGTw27RChOzKBXjzbsN4e5V4KJuSeXPWpfnvoZzK/
9TQT2yRdjHfBLA/76IgFgLKMcaAUIocivhhG8oKNZytSHnGPedtAIRrRTWt7WB67JZ4yPxp6ROIT
0cId0/8kPG2xCV+cE3yGVALOThkP9yNDh0NjrmHB7Oa/qHjCEZXmWcBlvjkuVDkBAJRBCtBe/QgD
cNXxFamVymGDzbmPpagDd9X62pppckvoTh2XRZYojurptweRqwj0tO+ymK68HH/zqOIoUejMWXXp
kv+zkMwjTESlyoxMlFWxKoOzkNTKn4LLjU81fHpd2ar3enAnhrKOtlltzV7oksoH1Pq2+AUoSDBL
BQA3UOAKJP/MWF5cB0Byo3iKxKwV+pC7m0548IyHbkucRxVf490YDHmXwrUTSpAcwmAC7oxzV/TG
qlQhQ7u3KK5oUdBna/sis9moUC1jwMpJ95XUCYb9l782NKl9GDG8QAjv0MM9F+Er+pAqDjugJ913
UiOO/SY24h9LZaRVJOwRsR3ZpQLFkwIVOUHWI5YB772wrCTfYPRqatoD2x/qH1y5qN18Aa2BkVng
xQpNgW3zwS4ExgFOcZpJn1qV7PqgDSLOUEIAJ9CJ3kKnliZ/u4uAuaXGuYF+NE0z7RKL+QxlSEoW
jjD/mwpT1+yo6zAaIDZx8MjgKCz2vEQuYRGhgl4ypRqW5TiL1mQKcdDdLu2O/YnA2QddfE/4O6cS
PhnW+3+XqRO6EpJktT/QF2KhY27eI0FobPBCrZVBaWapRAXK23PxUBJ5Yk6aFChSej4o2YwEvLoI
8ls/OdjeG/QkmvrBojxx/cJYjplYKbA9qpvpRin8RKpJ6SthMQGEl0dhDu36BxSvnTXn3bRtQu9C
9m6KHcnfi5wLPvBRJcuh/5srwPpAi1qGp5YPJLz6aOBhJkZbPu0Kt7Ld964cQYPHxFRcjd0DvU5f
cfVBJbLRvHT7Nuf9Q+pG7aXlDZtArLuKL3o+fJN+bEdPiflE9WZCfUobWFd6ce8uLJVc/9XwPvf+
tdo0O/vM2JtcXQQZmfxlCIteWZvOxIWjFUtypD396Xe0QhKV9gQoIKjyGuwXGRo3azJI2fn1ZkA8
bV45QqyXuwp21eH9McB+ZUUGEuIgeB6wx4gP35JPKHfhS4rG+7jxR2NgqUPfDjz7Mb2y57r1Makl
yv+XsVBnHDbI5ZJOoPrjeY+Zd75guKRiJCyDmJoxKkKeTdj0vTSJLc4j4i6RftRhqGE14Y/iCV2k
G13mrjaLi5Ugc/6mCpMSvwPPQ8wMp1XUtSeTtLyN22vUFQumM3BL2aSZ8Vo/HS2S3vbn2SZoaFiy
hO9nI8C67ZKyGGGIEfXaj9+CU/TyN7vnHXjMa73Sbz+ejxTj1Mxf3VSuOi6x8n03nCD5L0bAVYW2
IS8rpeCgGWXTry5q8IxAzwd0B/IALy2V/5vcpm9/u68B875Ecgnm1kd78hFyi/Va4b6DN8bnCqnL
wrhhhwtKhNE1bvBs6C0e/1ZAvx7uC06R6wPgnwRYBiXSnUzvQeYdnE/BuyMkC/GnIjDDvyZnLxH5
1NMcqXt05eUN7JVR7ZZsfzS54TJx9whUMVR37dGuNHs+AGcKmdCtpXQjmjV7lgK5Yp6ySmw5jvpz
qigVbrBx5V7gzBnBgA3WYhb1W3o86H7a3hxOpBuSDOxfm1q3i/oi3m7DloiWRy9djiceqKzdRmvt
okdnJZl7wLe6Rcct9jYUKRZVVtlhzAtqHwcqSyL5neNv1Zi/X8nwFu5DPgqZkZk+c2exn+i0cOmb
M6THLL6zWHiKvQfW0t9OJ8ZtA+uHYPbzz0ad+6B67A6DxPAuJNxzOhw8dFYWODup2DAlAFXTIbSu
WI0j1HWXry46iIsIE8VZhaQvJk68k22gh0XtcWOMs4Xcn6rhmVqu2BsgG5sQM5hwyeeN6pQuEfCc
vLqiezusgyIreLBrg1OD/sT5GJB0dR6KN5sdjAKnrViNsatar5HQnomgvFvG6NwwH9LP74Y+aJf8
S0ei19M5DGiVeOpTqeKBKxR7oDLrrtg2y2dR8nkh4B8CFqiUpG8ViOWxOAk9yhu2i7OGP61fpvgl
EX88pjZNh9htlZtgV0FLoNQbyhLa9wCE/3CmTt7F/Qi2B6FaaxvgZbokscPaEdbAA3lWVKlzYMrP
wgyCSMlOJwxiJTQKULJsEbQmEBr+783TfbFeHQ0ZGvVAw8kJViXgPE2wyIjnysk3JWWsCiqHxqLr
F5Vn9iTD4wt2wNgcNN0YW+3DpeXLjJKemiJlCNaH9ebxu97pB9NzkbMYV0wWUBCDuhL40dDVTicm
f9XZ2A7Zfc/MSyiOMp7YMvd38AeLdbijACQgx9whXX/O/9r+JSob/l9poYOVAHGRt5X2v+E2epGp
GKnep6zWG3MbcHnwLlq32paA9Yw4qx3Gx/Gy+6S7vzX0j1aANv1rx55U+6e0Zqfo5xPuyQOeLOep
0/Gqt1+b81w/Kho891EIb/Yq5riD32QoNku2USXx7IDsO4oN9NbO5G4E9xK/UKpzvD7xPS3nAzsP
/M89kjyVliFcrpJ+xbtdPxw2HKlHzlidTFSiCd9qIJpzSGK1vRabDZBQbAq2No3TiC09o7q8J0cY
47DmokDruHetSpeK9RrETQ6fDddjYHzq/vL+ELPP+OJo6tSGA6k/elKD0g06ONGOHWZnnjdEDxiW
sAyzq3j72NFgVmlcDHTNybXF/13OZqH4ncCORfnv5u6Hqdz0T15aoXXye0KYS1au5PC/vGQUpZ02
gYTCezHECOHh2cOtWSOZlp74h9FJx4BbXGjsGP4KZB2rzJ6k1VzZzbr4f1rA9tk6VAeYVLDB4ODI
4rsqwMbbneaLQ6dIAUQdvBB1m926V6wHdK16VZN9YGS1ujAIqEtblwLMQGJV94eNLQ9GZPbZTlU2
2HJnxxKuoJX3vxwHc0HVOXFNt+zcuSFT2jZtKk+eAhEyHk7Hhwifgg+uA1cXZmyEDV6Uglxj/tJb
PlmqykAjqUH5aOFeMG0JVzI2rCvsR7bC2qNsFGI/stonRyFOWSxJ9NJDObrs1l1jb2JLJJCBkbKf
cGTPrnNKrx466i79o6PS/d++q86Oauvjyq83Ac+dp7gTcDB10OEU3VZg1BLwzVv7pmR0MJ6O0Xhz
/smxAmrgjeY9GqoDglxA/DUjNkGRDI2sSjjFXZSo3a3mzLDx8WlsDwHM+Q/fBRS7BCZ7HiBckaUO
tDRYONJ8Lw9J67JKU1Kb5FNtySWCssl+oOO3FAXa2ELQJKnFnOALa0BdmI2H5WT6wyRRfOC9Ir8s
AR8mGPR+oRwmTAb1NPD7mSmStkTdi7s83aY0m85fV43cQcP08xPRuc9sH3HReD9/nE4uDLP9VhOR
E37okajMaAMNCkR6j7Ynuzz0Dx66iC2A4QXCqGJCwJN1KcnSjQQsmrPygFjInOEzi2aFvxS/QOCo
VsBnmP24AX+jJRVL/9x6YCBSCXaHdMPDjmSZyV8d0UvpDz/mzGIG/l/ZKENjl95U/cvb3P67J6Wj
BYwXyHJvqGFHFlzOQOZxWpvTuo2J65RDkwlTG9VjWoNWdyiYLYeRq8Gou2tmzzOrd3u+N0ueTcdh
sJq3j8Xg0te3RlOukOuk1VExsOR2XZrPqlJq5bp1L0maJgZBmm9FY8KWJzKCF1O7XbLchBeyr9Xr
e0Trc6lyi6k2TowNj9LpYJmzaYfd0F9W8P7W8lrvk1QqZSwBw27k0S5Z0jHQE7pGbDwcJQS+xkD+
Z9VPQLx89xyZKFSVFve/UU/0zzDWFRyIepsdqLfiDIykVMkf70RxoX/o6IkVzLjCr/n9S4Kci/P8
NDiZQTwjUIqGndUuCZI7vloQqTbzxrTiw5j/90goB2UrhAdAI12xBQBFZdDmxlK/LWPVLyFbXFn3
sP+6SL3DSZMX7Oqv7+H+r+MBSk9bte7m2dwqwJCzEsTldEfoxPg4AHsT4efEfmGY117Dn3VtL2lR
VYgOxiydctMH8T7bZDhx4SwAEHdjQSZLTgH3nCB2Hm+kp9aNx7kY8p52Ggp+hZuftDG+JqJWhrWH
Env/hTiT8diGlq+wohUFMFmTLKKR9ZusdBrkwMdOY4oWkB9pPibevlGrVos5Vdash+/QWPeDTfEo
LqY+2JMON2xj7qqcq5uOaI6E++2OtdEA243dfFJjOeWoSJeZebUE/gV6l526kcLNjEhCUa0A+oO7
ejNXi04jR/iQbM9DfJ8JgfXYWh84GyXs+7YAb4GZFC95QBHmOacR7y5W7fcTOpWYmUeACEbpdded
I+ryqmFU4FaNaTbs0ynbyPs02NhoMA4Wz8R2bQcWKyYwTiUxX6bOyorZdx7hzi4VlgyBIwfIzDwk
8I5p7FgPod9cpM0/7HOBLOcA4sYs8q34qvps2KaKyGA00DttCQAMQCTONPVjn5E5UhHM0jUmv+zp
wzSOt0fj+yqCz3wrAvG/aiRJHanlxX0Y113cuDLmzNO70Yvv81sxhE3O8k070Htmxg6tg97o5q5o
ee9XcQu7IVmzOIJ7dbWE5YL62WYQLryOECLRhwmR2+AYQ7pC5HiQErcIf3KhWwchOxO7mElEvMGO
wfhSc/qnK1+SzJL+K8tG4SGdLzChPEaZaa4RpSLSRbWERF5c49tsuFMa+SmhVEwn8FWsrqHN5R1X
7nvVTeqMLQiWSLYvAo3xOAnBHxqgZ6iey5962rXw6LgCO/P80ovZdptv1aW81MWEMe+2zIgVO79y
h6bE2PpJKXpBwmPo+HMvgNucwnBuCvFAluhdbUy5AOQbpFQPLoAFOIKKyQdhMVS51OejmOvR5PEV
3IeOkrdC2dit3AMxm5+ETsQ65f7ZRp+klyFb63VSpZiIJvRbhnLx1/nXUvL3InicGRN7qKRX44Xq
W83OHPnjAq1cuXBmAhF66AKZAmnA95ru8Fkj0ic5/bTGZSMMDjMyFEmMJLdpsRStBmP7XTT+QIIQ
fNuAjVMzOAajMGaY23Isq+M8acoURPKBhbPbndfxPTtDG8rzQP4i1PrE2cfk/gA7yENx8JLh7Wi6
SRqyWkjJPqetf2gH/t+O6s2lXGT0/eUL/bHng2TlbCKxOqdfpNd/8XdgEWpmb/sKsZwHfZvCcBsU
lAF1f922pTHdWV8AKBcTGg67wcRlilZhk0S3wbbLFF9GlOmLxe1k0chJZo+e/YZ8ulEYrPPAHJyf
Psrnsa8fjl/TQWZIQ+YMeFwjAqQN6fcTTUBoTZ562StujAWNTfyM02QJzN+O/XCZiWUS3k3u+NdL
r8z8SxZaUK5AQTqiY6bygYGv2wHA8mQxSumSuQ67NT9FmJ1CTGd/TuVgqPupQ/J8gOEmnsXE+FBc
AOfDG2tHbyWzWF3Zs51z481NCodDikzCQlfb+E6usY4EgTTOGfSDiqtJ0jbFpFZnYwQ8Q9kygpwq
MhmE4nooKjzaRjitrlREoCl45ki1o8uVmuyp5eE8co3pIoPBNyKAGPKMudNIeyD4cYWI7jmTOh43
Rzesgnu1pU7bfsI5HpTIuIWRPhZ8UMsi7JBd/kd5mirBP/zC+GMPaN9YTbP3/krxqvIJBnrrpCgr
olnyduzVr0Tq1/+GkpGieXsZvvovQ3J1122aQNIZN9x628gaAu+ZlA1JVx4TMXI9IbVedpmTRaNz
v/jDTjwvR2A8vS819K/HtALhEp3reB55ZKX3GLNmZWh82Gx620tcqt9QsOGNhZiGyNS6P298hRJr
naeI/DpggKRTH4ql9iq0RFZP6iNMHnlQ2WWSvz/zcUHqn9bWtDpZpUeOkwlT1z46qxovW+G3NoDh
ADRQlwrO2cVok3JVkGSF1LsdbHIWavyyfIVlsajzp4RF7OEAhYOnvsfTSwOTLm/fm8oB04ZS3zcn
w4eisBJeLWf8pJRMlLL9e8JertqfI9jJpEc6qd1iEyNSOIrthr9B+qhjA3z3MMZsbzCzCZc4OzQY
sgCWmTAlNZxQpqa0AWZJmwQ4bjm3+OJQB4NSFXSCvu7IZcfTcejEjgoIYQxm6jb3mbB+5QVuhqFN
O+rW8CLiggmVxOQp1Qp1JZFtovwrxooUIJrlq0z9czy5TL2E52n60e7uuKFwFeB1y4UGKdfdyTuG
unkvo2nipBlM3f0/Vf/sqF4uVqgdO12saOF02AVbmF6ae1vhm9oDi+DJmCW++NhovI9H7qXu3mVB
LNK2Ip32RNNYPQtqFz+6FCvpRP0GKGgT1ZCjTFxU80qrvx0DuZFUe+cnC6YyCrcIwv1n9o1zZo/J
gyovm2MU6DtqDuzrBxUSsQJauI5gEyfNmFFARWuYU+U20huSr3TxjYYg+kHoudqUJ35+x4AmI55u
p1LSnPcvlVy8W/6qKLQ4wPqVijcluRKVfTOF7aPnp7DVIXg5FTQqn8Ix7q6ZcYgKORBDhCRi0ktI
0S4P96UonG04p0dyc6Vbf2ehPpkGHOPUfECqjyHgvkZCZn93kTN4mmALwTdZHk25v8I8F3gWs5eL
nzP3hdAKoIiX0a/NdC5hRTKoKnlSfh+pGlwiOPV4xwA94vK+hJwmOvkudp2PgQsGXX2+XUlZESU5
jR2O3M/W1HyI8rGwzmcjb2lpv+uGJgb7E/Hz9+Ahn+VTZLq9hGcdZoJgTkD9lbU8U96P5sgxdZt2
tmsV7ymPDOZfoMD5xBaH5O1cnOdOhTva2bBfG8MbZqwAGRqwa5hKia01d2DeAhNHDA0UVfvOfJHJ
NyRxU++WY4kNUkL/qMX5WLpoFTFCAvwLVHufhKVoopFxTWFH/S6he17S0BeUVslFosaYvQa+BVgR
Vm0x4vvlstoO1SkWh8hchT/JDpYYyyRgDlhK5n7iQVhbJylOh2kzbL6YL2of3dhLYNqt4WYPtg6r
jRn6BDMhWxEe78IS6qog4f6yyz7b5pF0pWpd+UjdrCF6kMScv+c+/Q0MAl2i6WjfJgZ9BygCXKVe
O6SjjVpEIFxSGhFBkdo+A35KzNvk1N8tKJKa2+s5gGS797/fiNDiunksD6wKlgXD0d0VA5I61thB
qOlRbgWkTxoZvcExeF3sahWWu0l5tn5Jy/YxA6HbvpdN0nF42dOG7t5GM8G+ruTd/oTRkwazUWXQ
ihXmEiPPneJUF+AERos/1jn/6pq/UlnGKPAdjWs8iT85pbXlNdk/1Iyzn9oaqcffes+9k4CXDhbo
lFE/e0gG9VTw7J+hKm6tEPrqOrVSjlaV80pdrwvZiQrwOGS2wCnJ1SeIZTZk7AVZyuTAV6r7JpdH
YaUg5n+662a7ff3L9GX0oAwhsCR3beVbWzg0VIppU8+z2oAgXvfSW/6DgRTjN5GH47B7Z49gzRRX
qREVT6W48qFPH97K0wfNCEWCxwhdTh3KzzbjKuhe0dClEj7CYFKShXTAs12JDLRj/WoEFr7+RnZ6
slDuVpJUeS7xm7l0glvewQMcDpefsObBTif6Anh7r6Og0bxlEVLwBuLF9Vyru2+nrp7VzxQmUpx6
3t++53DrSqVieJmxURv0VcOsVL2b9C18IfQvFH7dHwTVm99WgE6JUOS4GW3Nw1WkPCZh9XMZffYf
HHZ9x7rJSfgXisq5VdNqi1vjipbZc8FHZWrtgEgT0M0BLrcwazg909MKphEEjATuz+ZdS04Uo4Fd
ns7k8fyR/xelodpg1TPrhh42CXjrEbJI2IunVqNznispMvyIWaTW92CFEZHwxxanosAfISuaI+OU
hPR3gpbEAiO7x6dcl3NBzdFkUpCLKKoqizI8tn//1ryn+rTw8yLYWYhviB3UhQeGenP/E5nCvguy
OtafiwZ4qveCs7xoUi9Sg/1japP3XKTBfMli0d4VQjLp2eK4MNbOfHQTCnTRW3jjgfkSqiMcWPiq
hhbcRA7dttNFHw7x4Ud+KPnYZe4yTGpwFQof/fxZ3dPjAABtmECZR2dJE/6/pfgnNH3wsl2LYfv+
rYLzmJpAp8sa1d2k2gTLJLFJ5xAWOJVXvfdA7N6V111J5kAywb5ZZPFe0jnbwfCeYS59k+iuiN/1
QeeA31sdj+hntQQ+Dt7gRLB/VJHRJwOQu8on1cQXEOQRCWfYc+7kcOytmyK2C8i2EMdsublXJUGI
+dZtziw0ulio/dnDN39hf8zHd8vYwJsMQBSNMVFKUq/RepHqWCXZpdCgWaD9i0ujtmIDCHppTEJ+
MUTUdhEjwz9G4ZmjMmfcgX1bbjP8Ag9W/K2586aZ1WwAthpN9+WGCcxo/+E6R2JCzFP7R01O/LVY
TEzSZEgjuDYOqVO+RyYZeFoKXbVTjWg5/RUCpIOap6esHqF+e9DBpY1fI0aCcMYO4zmW0A3YNW9l
DLwG6ebb8m0ScctXJzUuPPtUJZ0fe1i22x/4y7LJdULdFw2kWFtzeWHi8A03RBcQBeiYk5+vkuOd
UmICCzhF04fLyYyzkTJ8fKK/Xd33F3v8HEgN40uPtreUFlUmorj8ACrFOQo2b92yvnZq06R6KWjH
GBAGjwsfh1apkMoaOEhyJhsk8IDaP2gMrDlVu1vYe2513TbejwE7zaqQQ6rvvwJRi5DYDqmkdqB5
eOsZvf0j6f1M1ZsoS6sbVjOzLOQNZjLkgFTw0M0QRempu9qI0pZWaR0DsApTiDWrPN0Djn9ahqxX
fDUDIpfc1gqR/JQa7sghoyou4uY6sKBQLdgpmvyjZpwGDOwyaW4rNZF5FBdgm6x6TmKu9ZEXOTYH
OhQ0a8D9ytWBxd9hPgzqs2TVhLyt8NAModYdjGylY0I99cg93K9jiiPag8Xq61Fvp3vTLS8cpURP
x2clz71DIL+Do9EHLOIhHvKDHSUIQoFgXi3ANnYNkPnUsfaNAmV3pBoX0af0+azbbUz8E+WheF5F
iRFriqgw4c/BK6EbnOF7zb7s6trLWr+mQUtVPQcTiXIXw6D+UjksWN7zC3fK88k1f41vHKUhZBr1
xuoX4GV7jZpJJrgbunsttX2gPlLrEpnOikCa8o/LilC0GrBVP4uNy4Rp15BOcTeL8yFDV9DoGzB1
VJDY4UQnrGI1kGUk0uiTCEfi8taIwi5i4cBd8lVsqvpOF5u9Ho1Y/WOGmzAnajYwhaIjOZHiExGr
N58HbOA3sHCFv4vrGz/cqk71RiJhZQZKle9CM1SPt3wM8HYG+6HgX/JwuNCin3JFlpAoPfwXmTL9
FUB8h5G64daQdsZc8JbXC/c7Os0ntfppD2GFZDSbdT2XB/eRVtu5ka8h00Pc4T5ZjOYMVa6H5sSO
A9jACQ+ydTEaJRZTWj3VcsQS4ag+dp3A93B/w0LVFYgoKGMhKF0+iHX1Kv4lfxJuJ0AOPSbjp4vJ
Afrwldq5x1d1X2XKoux0hUmy+BGIQIC+Yw1I+3hrYqTjs36RL9MnHZOl4F99l1MvNLxhU5+u5RWs
fJpI3IV3n7murmuypHUjKiEi2t4C5VBBMtoEEqgcHMnWis5wUQtTKcyvkb8BSxhgq2FnxCw6UymH
qJ+qcwXZSHeRXgIsoyVJxPUDAWKGe0Va2Ncg0lCDWxLTaFZGKZEcgwTnTbctSe6VCOt2r1uzxaNp
Sw3rUFBV4SXaZ2vXyRzDGvcCdUKKfy362wT7ol6wzIAH1JChsww1puyhMoIHKEYbhXVFliUGcu6g
bSiF9G2GloqIRMSzpO49Ekd7mF1RUhYLTLBZr6rI9FTBzorjftRMOcnIjZWVIRObYF1xP4BlT9IY
/ycsTkYgPbZ6CH1q2Af42DhnZKeW0WmYOK80otwCzKeiXU392dzjlkxSwoMj/+3+4aJuSaxhkNjz
OcLz9wPlh4UYGzXph5I4+z573G2JbFJVJ0eCN4O+JUT+r1eLTgN+3XVzCC+lUIWRUmKJye6UnK5i
cxBB2lqExDd6zCUi612YXjQyBGJ+VVS0PFPa4XS95DwaECgzqsmHlOxQTimhUtg1DqrzU3CbIJik
8IkqS4jEBBRhl0MOuCh65SvZ/Fwu7KOKB38QUvhm1Wxr4PFQl1aPGEtbhp3wkwuRZG+KX/BP72BU
dxVypCeI0J8WtgLcR+jSq5cQffK0dM/BAd1FfaegYYgRy7+LKBhYDLnSgwRWPaFTh3w6Poy3JjCU
U0nL+V6/Ja9Vxf/CqM4HgPhSNS2Bn2J0ZP1UOCoIpg97k2Y8jzVywICTlgFiihq1xUlzP9jPcwFX
YkNRshfK3XaPbJtbj6gbJO/75o0uV+/iOGED//uVIaW/sa1I3KYtM6Gkpi7I3oc2TmDV/ZuFOzdL
GyoseItpmJ8XMd7h9ONXYnHz3NPMgAaOhpC5s/8xNMihR4jmNSL4nytJvv7IBHrnsJ+xRMc9MmMD
ADktDJnZ55dwTj9Gf0ItjIQfZMmupt0ytZ9e+LOarAEVYNVw2hJTraxQD+rd5l/Qxsc/zEBFr3/j
fsy9udDXBz1BfOSPNSGzMmInT2NKhxfsLa6kdKJvZFOtlloBt8S3OUFZ3l0TDg+xfXBlDordVEtT
ZPzvzUQfs4t9R56UjWWIDpvXnUiP0sCmaztrQLYffTqreC9TX0w9UHUruFDSBnc6JD6wmpzvrJ0z
SZYtyngAwx+qoF6OxW5xez9Ug/B54PlWx3ZHWrwj0JNkQAadx4VDAJlxm5WDyz2bgy90eu6Of6mj
5eCPVKLkMVgDu2XoDTbitbJDorMw6h9ZjlEiKyaOlbwFyCTZhBMLf7xxkZIvKVkA90Cd2od9DNfc
Kwzgro7PXCylwrec3firBUXYWm6LMLPodFXzy6iX3vGYSHkcGDGSDdL/8TurP29FKTxTqw6I2qnU
x7YjR335lQ/mcpLbXQg2F9aaUjtvzBOyOxygNQlQ/Y0HMZzLTHfJKTK9u9KDAKNwQ8/PXvAXkOgV
v26pFK0Ghq4QR4wuxsKjvDThU+k/E8fMJhSBgAA5MPrxqgtNzvYX8XqWE1y9K82zK7MqIz8Q4cUn
7d3cZp8PfGu5C3TTZu5F713BQiJyJ/mv/Wtp43dYhHGrpONgVp9aRFu//o0GD4zHh2gN8F5VLSvX
NU5FXoEdhH5qqjzDmFbbscmdlng0qsldMM0yFwGxIbVGx5Y0NQH9n+gDmDx6fpoU2NCzvypuIkcA
2do1Ior5CK14nKsf9kitQ0eHBN6mqYvT3plMfp/W3ju84jM8lFKPSyggaAu87VCxqZQ865KWUqTu
IS+uw2y7ylDVywM2bIwOKCJ5dr7UBu8pe0xjD4vH4hiau6Xx68nJrIgC7R8GlREww3fsp8g6GSLC
Zx7zmyxCmFfK+LmkdcnkW54jpilF9D8iH2h+ul9TEkF3v80qOTiBGm802X6fkA28HYGApclQ1vN7
NN/Abr4iIy0uGPSDnhkel8kRhCijDX3g8bNFoufPcF8k9hmL14jYTZoe/lyv26GwvgdLT3LafcC0
69AQvb6CTk7y5oZnlss1NrarP62PtEohwchp8X37Kd/6ipn8qXscuk7bLsWS1S9TnSnjIXzh5VyP
40lsU+L5CV624AekNpJeUB+rFvudHVJRBmV/K4wYW2XQWrBLe+VgTBbxhRm24E14j5vo7nbmDHYy
IP8KLbqHtCLSC5nJPryHCzv0qYtqXiKr2mXnGInZATZpiWJD0zysFpyNRFozOde6exLMMrMov7Wk
Z3mXMeQ/fRdoRuCxQEOXgft+fBpzzkpMpCnPNWimu79mZ2xrDT0uNtNtTpJcYmtIxwWUiTlpV4JT
gRr+VFGnsx9lxgdZw8RZ7GXynj1ThAtd1EIRPzkpEaPJnQ7qFSsMGJz0lowRRvzkAE2pcI4I7rwO
X0sp2QmTKYX5TcO0VBJ4nsOg/7Qrj1PCiYUsiIl+juRKWqU/HNXJ03ywEN2qB4qGZgBaozISX6l7
QDjVVtGayJxitfRUCOSwDfK1CElja3q9kd9rvLMUlCJcL9QBACVQuZLqAPpjyUIqrrxS4NVUElLp
DOWpKkd3pKL4dRpnSx5p90FtLTQlhQR3tnxvKR3LQ+u/XE7N+KOuOWkcry/rweOudxwp7IdynFAl
nhqCFP4742ui2JAI9So3kAoG/afawzfmWzLeRMoVS4S06ulNYTImM/qT7iDOZ/8WpaDqnY6TBnzd
VaFBQlEFpJekmCT0KFsKaKDAXEYlE37DYh5wJj+5njw7lPxRHXwze5hgdLQD0dqTJy0kz2IjWFvD
/LyozWUBxBpCsuyktXQakXRDwiD1Mffk7OOvv66g3Qfq56RkEoIGIPqHLb13ipYv1Kz4r9M0w1lF
htCtcbn214WF6CeMnm+/VORXdTtYKBkOPtqyGOgUk2f+K5SN8ZtRM3MEf9C/7ccTCymU5jFXzLC8
uYue2Y5O2y/iN+AxTl0YhFr2Z1ZUeCJeCUG4Nbv7L+RoZDkx42F7Wztec6Vm7daL8gEbl7J9vaXS
2obOQjdH+69MNIMusATkMobNJCDNt835cW9ipgxnbkWi28lZaXa1G0JK424diauY2FrTUgy3TX5i
vuV+WctoHKkf204/nhyJ+SuwlC9b3AG7PJjn9jnU/+bZW3K4LXVwka0O4fafr5J/A5zwscLRZl2M
rdfByCuwuGFrotmsWrZWWKL9+IPuKhaCjC1URbjIyeyhPDNxbXrDUhrdzWNJ+BhggQ5sHv5fFYvx
RNpNPfdjWUz6U3Dmie7nKMiap3on0OKhtqs2HCukTziJth0c5uKVSOUy8/peKFw5GkW5M20r18hR
S5LVndmNDVJ0Gd+vFlaVSSn+vxyc40xx1gptFFFD2IwUO+s6lLNCk3aKTGgmNttE3BKTvWH12+Im
PvbdyWsLoizzScc7yI/DvAI2hq25HVrvGuZL++0zZGPyLMnhUdlnJ0P6w9xEG+x6EWsIcltIiddF
xSNL4CHb30yXEr2qu96JH/ysOxHMbsOsQwYVZl/yjBr554e8vccIvcBZlUQe0KORe29rOLm18+Pe
rHrDT7nR4XM0fFIs1ICZlf5y/5b5bKxte1nQng/voNJTuhbr0ZlGHfkqCKBjFo+18n4aq1ej5SSO
ruz0VPp9ymd2F2m5Db8Splmz3BGUQs6ND+Dm5l5HbsOYxxcoz42A2lJ5JKe2ncss8JqMaJIl/Kpx
0A9QAgoL9OpjG/e8RNydPHrjNSOLTL+Y9tZVKUUQnyhERG52H1azZQDO6hJta+sBB2MBl/FU1L59
UbeBfe96RDTFqTiFjp7amgpaDGtpTHvOo2Sru7ipxovbXYeLnjRbw1KLHdgfCuBuTDmKPQX98cZ7
NRX5gOS2Zqle7MlABpi42Mblb9d9jqokFyIEXzlO6JlBR/nETiQ3nLgFgWQqHQprEHE1o+I6/cPf
YI22/l5kzzE7SnGCv1Rb++vbWq9qg0VarnI+R6ymA1wnbltRRmqicGI/sB0R3YQ1aHFBTxzcUxWI
z7IfA6bHpYLVSbWs1ZGdBDaMM4J/lS2p/v6EUeRPzyN44ubaHBCwPNZQkG9TxRMiStScKR8/u1Qd
YQQuL06s7/HCiMwoYtFw2B1fQSsJJEpnHNkS8wWTDyEpOcOtdJyJZVcsZJrrr7xQ+mkZp+z+tcZ/
kf/syESTLkffkndjDSUf20NvdpesPnOkqF2QoVsljwZcJ39xAR/Mmczdy+j8x6nRaG1fr/yQt11v
UwUfhwb3Am+mJ3L/JuVqX/Pryom80vKWfoDrnwCxLR5yIAmiV6HLjQCqx+xWQAeXkiZC6qosnrZZ
dXsAo3Ch07Jr+6Z5acdSmAv6kZNr6IrfD7GezNu0TSgq14SkxryYyEFbK4u//GmJgKuAsAvla3xq
ZYrCzee8y10grByU9jGZ89rqTWi5arBrb3oltHodTLjJtaPx0rIiSRgQOrrl5QkrtsLuMYW7pDiY
4TFzLTKSiIXZFk+pfLrUXGZz1ms1UE8rGum1MzVDiEeIHVrcmtZCPEckZoFo38HpQ+PTCX8oLoDA
g9WkWYRvwiG8uLZK47vjJfj1x9PkUILgqdEyVsYjsy3S8buD7Okz7P+/n3qtl751aFs8B1iV60nJ
xpIPOINlQ+gOBMLgIZvi0GrJ4RQInjmt6qepTbOhvftn/fg3oajt+7WulV2G0Vz0CF307D5r7DUe
IwINu+wMakI8GH1eT2fTbGdT+0EY6kJKIjHtEwHBqWTJUjPN0VEUDvnic3TGNe4i7Uhc7NKqr+be
bjU02cqQyMlHt3F6UT6l0DjvQJJ35hB5qUiMeYHq95Zk73+3lDJvj6kBG+1j7de9ix3L3rYglbpq
BzLLASneZ9/3xKVEkL3rwuNk61Yf9MUBGgM8touqlgUm4fLSvVze7a/trVbZinL1kPG1u5AfL2fF
5BSOUdC0DtpBui+wJYW6mmcVWG23YrnTGcyUJS9xNEQ3XGe6n72h0joocTr3G+BdVvCxK3AOmV9q
u0zjCm6upakEEuRUCy+6ktTHqwoveH9Vj9pD4Sel2KC30McAOD+f2ZzL6bgZx4TV7U2yRnWqFVIl
Sxe4dB9hXqOOv3Y0vfWDgi/BaER0KJk2oS0Oj38PloWRQHHScNP+3l03XWVdZLlkmaO+BtonFj6k
dsVxBUNMB/iq5H4zN3rSQOSCnPaCdN7hlMhpuW2HgCBAue9DU4IeZApZmza+klForcY4Vm5Mmukk
vBiKeUyruz1zgYISKDj8hqtEhuKcbcLDoWvbv/OipFoSyvsBm2vyhiyGnJEvK8Gl6y6VC5w4IkTF
dV7PfiPFsCNfSgjH6ptzqek/4TjJ60zp89SWaEQIxGj+6+OvApM7EIrr7qks5fvKpRDE5JPvS7jk
+/TyicQWMgKzU1GoUtOpWegN36lDLi/+aRZ+wRSIPlgvdExVnQaFGx0L+a5N//kShu72Uchmuuub
TVWLOGvQd2B1TqbKPSq7E5vXHO31ZG2Ou4maMVSEvbw+yVyR1Q67FpOVb8YkpSOCZEsvmtNs/XLu
TFXiTBcxFPkFYZi0LPZUJSFRrGbZ7+HVPYLl8nst/SVEo83TPkZVj8UnDjhM5MQpikrZHZAmJtNN
Gr53NtAi006sg+GTwRYIEBExBIZt6IfZQRQWFrcZocxMzjfxem8SxfTPmyLkctrHP6PP1kdRSTLr
qXMDklVpEB46XQYRGRzREPdE+3vq5/tDbd/K5IehYHoMTWP+x2shzoDFNK6epT0xfpFfiChrvLbf
IQrLY2O7mWW1HpvSHFVconRP7p/K53Z2lSPJRCD1o4wCGBnShtuquTXD2aQ2y1A7ouLSGO7OS8xU
6jFGC1f7fcxMppLI2Pi7+V8umlJOuTcoMV2AmJzlOR7l/qURr76aZHlwPnep6mBI/swSMUG3cM7U
PJoJ/KcDK9N0jdoKqOy49ntFGy0kUWjwBawjbWSl/6qGvqX3WVXv0hoYuAhfIQrto9sZ58otAf5D
fLmYyRzgSqLvohAMpUUtgnHKuXmeQS3lSDtxZruj6m/6JXEaW4qVe4hqtYhB/qdFtRRDfkdrnqOq
4Vk/nTe5mkYf5NPhPV6m9Yk1P9fWQW8i6ZzaCXzPeQ2nNNEiJijj1t/XaVCXicGMh8c7EGy8G29J
ZhNBDCGUiELxpCfEzofEkkc9cFg7HG8RQ48grv2qNhdGEPqCAqqxlHxM9OzxQO/XAL5rwiRbx+Hm
lfgImdS+fc0lySq3m3ksSmpD2pOYkATSgfJTkGJXXduZGtT4HmVdyIe3PXdcdGvBGVUhnrXB4Z05
YjWiqqpOIYUhOR6YA0Yf950OWes4Pd0yY4Qymc60CCc0wwX0rfBGupzPI2MR9YDUm9P/V3PxpXr6
2McJKE5gcLKmZ6EgYbf4baTu/a0gqXwGUblhsNv1hmxm7PvzSocCvud4xsBF6LU2vfydnRpYYjaq
0+RiszhxQEd2o2me0vPy604jIkkt2PMYrhraR0RN5500O61Mqrr1v83HVyxmpLfvyXfE4Hes6OrO
ASSuI9CjSgba/FRX6r60nnUMZkybtNxLHstesyCUjfNgzhNogLO7rXhjFpFbhbZ0EWdXAFhdmGpo
OYnTVHkRONOmj93Rbepo6WFIff2QAXimawsxGLy2YljuT1/SCK4jhaAiCJedcDZfO0yi3voOhg7Y
cdeHc5jVOMzkgHQRfpg9lYNaQUKYk45uZtAjw7TfACpxbbLUBaO14LqxsIs2ynhk6RVBj4BIkwgL
2qoamc/r9YoCkEPHds1qIDXOWApyI2m+0n+ofB2GfmTazUQTA8aVh6K8HzR93yd/lmvT/MQdir+f
z/57P705VDXztmiZ+QtaOqIzVWwVFP2muk5vBg7cjXcKPimcrlSWf46kc4Ro/f/C19X1XiYqB9dk
AprxHiLotFw/UZpZEheEgGmybAoIe7N1M0WLq1t7Af7i/oTtLTXF8pd6ijf24RVDNQi42ujRL/bK
4QSWnM7STr870/WfFDy4NdKKzpYu9ovlyFuR9xFpbZ1Jr0SgyJDy8Bgu0W+XCKkpBHf7hc4nNjL5
pNUsYkIaHI7dkfP4imGpAP/msEzJsMbpdts+wL/Zm7xmKjfHoTLZzM2zosMi7hxzYtYYyx4RVKPw
slxx6ReAKkdAHRrv1E5POGUQm36knXrTQuV/yKQP1nvxdPC+MIYb5QoDQzn5E7kGvlYiCdmG4F3C
llBRT2onisjC8v1nka9rHLvM2GjF5S8cWFQfKi8JDJtf5unzYfHpu3l+9A8YlkB+RQg8UAuJXqYy
Tvf3eN4+cPkpfgCP/rLF7eCmfpssgQbnZjRhII0RIIWnkn/fzRjR0KQAxEPuzYc1FwpvsJh0DCPE
NMCHpkhGes8HazGGYpM9w4kPeIWrtVS8LyGA0H8nLX9YYVvlv43rYwaE0GUidHw1bNfHqw89AZ/K
K3yCyfaYe4UqnEDEq/sCo5VqMHHjK4F80jvsgqGZtKcpRHAKCKrkdfh9AIyY/ZeuYGXnusyJKQW+
F3RKzwGKvxDumlbnTDnlzYe4pvuGXE8257ZzmLZaJoozrBdofuqWA8wyXV5UNuR38sMzfnKJp4JV
hI0QimmmxaAoSLWu28YMwLXCwoQnVAsUb0xrfulC2Jzwh5rZkMZ78AVr1L16Vldtcp97GPtGMqCB
RJsrZIfQo1WP0D0lJfQQZkp8w5EbUbgg7yIVQlMvXUXdx+LOCIu/NPZ2ZYdDZgLZUwp1iZFl0R5N
y23Fme/Sy3IdONSWx2mVIL7L+bAgWvXFOzHd65nOu1+k/JIXWzrXPw+Ob4EhPoiYAKzVoUDC673A
b92B6M1O36X9VADiMmo0qq4Z1d4tq2Bmg4jJWqiKcl6hKyctlB+xH9kJTQITgDYv5pD4LrIuLprH
mdy7aJFYEDKJxHIw8n/cCo0V1uRfsMfekqofykycW/lQikJaxq6/066U3NuKDxr2n/QpOMSAIT/V
PSdPzHioB91qBlz/rZ+DmnqlzTQAKKcjxAOK52N9Zs7p1z0oYUz++awGr7Ftp3876WnLbWs1/YbV
ridjslrJkWwh4WrMuf+0dl//yKnjaHjUK/CmlDP/gQK/NmPqZ3q+h0FmFqWeeViSIksxcsAbGX9t
1yQoFtI5wp5ANp70n+W3rfQtwxRrNwcP/IMk3ZcWjfyu7BhH1KNm74+JYO9wm7iEF2g/TVsnoUKk
ACKgw4jofLJvIhUm2voLeUw8FaAjWNwMotFhE48tsgmcf9Iup2kDEQ9iOMmtf06rU0mtDK6jxFbE
FXyLoQtUvx6TS5lcUX/8ooHEvCFe+ZRw+9qeVg8e1JpBbTFyZ2kZGvv4NtZhw+YlLd9nxp2u9Z7w
4hxdKLC2BqpyXLwVFfEEbsbhnaueDe8jIKCtE2+aBXPNsZMWgWRiw4F6N3uXUoG5anovfDkp25De
BpL8qNq5XPRy8NdrTQ8vOv8bfHP63PBYniuTD3wpP+NtJOVocTGJnUwiWLfZSijdCLzyoIZGfk13
crO+a6oyJ7QxfIGX9cRgjJ/7m7XkiLCu9wrraL7/CoP0r2lqMd2Fy0grrQNO2xveEmoaeph+7R4R
/s+1B1wOeFBXMi8JPXmbG/LDHsj35UuAyXkBvSDnNKKQDxAdSzbfwgbMYYOF20LlpugR9wMo2jxt
j6DEY3rxMUB1C/1S726GoxQfp7XBBlMJPtySIxrQyl1bRBSwjBOepZhakjWLj3a6WSzNjVeYfytb
7tsjzXko7Sqho9gnjY1AOfY2Vo8hXOdV2GbUFIugq1SJg4KXbbWbmyJ7krkPlVsX3Xv7lg097NaV
vvdiJE6J3AxifGNS8BwiCw92ICKxpeJj6LFg6QYVuR4Eq2mTs89fYsIQsY4Rl9dzWEK+S256dt4b
lzgBWckkiZ6uic0irh32vlBrASg6xz4WE3uq8xLjb8Cdg4gkyBCMPPwmMs7soSyPRgQS9clddGzU
MH1AYXZCWhJX6H3UazMrKFuUBR52G8YBz6bMLDpZTEctNK5NopI5y6f/9SnKv/ikKyZze7EWvK0n
K+ueEntALM29fM/s9VmxnVGY5BYJptfOBsbJ0FwaGuJqMWbLO5pw4GH0DJHVIV+Y7lwtNXcs7gYu
wkQMz5clQEsovxM1y33XhPSb6ITuN5/Yf3jiZoIaWXW3nGqJNcyLnJa/wm8oTT0T7AWRVHAzzveC
NQHzzZ/me8ytT+2nVdjeHnu6MQF+3XH+yKqN833GYYrK40F1hRimsC0c96EkF1nJMGLvRN0bBYBF
QmesZoKH4Z6NXxpw1MG4jMT8pO5KltqbAPpzvCVIYC5w76u2dxwSitp0bCGRbzUIIIL5auE0BNX8
i8Wnw1xzLNR17sPJ1zJVAmSpA7Tr0OR7jwUfkASroKxPMitrqDzDEoDHZfJ9mL7j9Xv2BHXblIn6
adOfavn2TV7JNasTu8bJ/nx/0X/omRLPbWTMqG0po2FfB7onxjWs7FN8NBegdU1h0EQAg8By7NeJ
exjee/a5kpGxa6pTmjq/KmWVu7leZROVsX8FUZHDDmG0cg1gSLcwa/qBrzDnQUAZ34RJ/okFBq/S
Tf/NTdDzFGWbERmdW3+pI6LGGIl8B4A3obG30rNrL0z1COXrbp6BrK+CvF32f4BjwJRV0xrXse+h
VxzgJ6xgVRV4npagbq2abU7rtMLh1Cl4LrT70Q3136iifsF3dUCnu3Qy+FLSysa3ZKZSNVLeTb8J
F/8LXBXD/7oYBxtjCXhh2XSAC4TWlGZeHT7vimiVtRfopMMkWITG/KggEAU2l5+6XUfkbYUosIKx
/jiRUgMUDvSGso9bvFBjylMm6kaBQ1Be6jp8QgMAAdktHk4yOlq4p89AywvnV5d/aUdonSZrfcOV
B0s7T7Vsf+RgCtH9MLLQ54rX+DKUj/zc567FL2oKstafw5dpof03+NsxYiQdETEpIvP7ARDVg4Vk
vCuB5iXT+6CxHDjH05K9gX3AXsvfa2nckfs2KYaqWKuDbiCjEqbdhA542NeaBoXfHe/m7sj9apJD
tjC/1O4fG9eHEvVWZVUyBpdKy6zPon2/pNOOaM5TH86CGhCFeNrujrUTMVWGygzYBx0NDVEIL2GJ
GGJc9vl6/5scyB6/52cCmUREgwCw69M9AyQJu7gFqAAmGJiFatzqY9WIy+jhZOFulEiP02wDXne9
sX2D1oE431W++OntAaz4VJe3aUaHmb/4nEtmPdw5Asz+1vmUhNkffNS+t08gCYlQ20pVeteDQUKi
c999pNKaKnZjobZ59o4R6B+Sff79bYQVMrEri4TCI6ik70hzSM3rVRkHUr5jPYiGrCdgY+6nPgnp
NBybZVjAAB1K0hy7oHgibaYFPSoX9rONCwvji2unTLIub/v2okLlnK2xG28EFFBReAwVRXwlywl8
4AVUyxhV8dMS8E1F7TlV1E7tCOTInHDUtfoquQdr3uA8y10IOO0J/XtKOKx13blYAOxqsrKIeq1M
8cJgF+ZX2mGxOlCp63FDIo+A3zTfeZVBWMDdH/4s0SK/p/S9jIF/73J8YQbKTZacnktZl97qdkpy
2O1gGMVn+yDEwzZh/i9KhjcxpEQ6Y1y+wIOhgo/rzI3utQw6kaJYkzQI7oL7zXSwVfXhY0YERzMf
XYfZ5l1MY/+CJv4uwk9YD1xP2xtYjOaFKxd8eLipH/Pk0gUKAvixiBxHqDz7k3hbC4TgP+75bD79
l+1YvQp0otVMm+BX+3483MExj3v0ghuS52BeD9v1bbSwgd4uWkcANBZiLPVOT9SQIFjxah7GLHd/
CFyggROJ7lIahiz/e/jobWRAVYhUvYM9a3exAxnfqwTnjPBKeCr2aI9xmg+2diXn4AWEHyyF1xyq
mFA1D0nZdBbCgKI+PJHaXapC4oZpLklnyYBExPfzPou22WgyXE2erswCCnMYu7DER4M73pC+UXA8
ZW+I7lLvbN980wRsDUQw9LfHwA0XodimU893aUy8xxEOgBbMoYgXuFCjZplp2dGaMtI9wtmNBhcI
aXEgbfFl5AMouyc0T6GAAouwaeJI3Nho6VUjTiH3hlweSwf+Gd9heEPJ+l2hUtLkJJdQtPXTF42w
M3D2YMF+wPoQR2BjBsVkBJq/u60pUuMwn4NrtlsWvUx1ctKyUR5AUqpjlvrKg7aiDSkHatUVYx/z
jaL7qZFMyT4Uj3K+v/SQDCLhtHfTiR/q/eJxQNd1nJhnKWpWtJDAhCfKT2R30IrQ5gY/JPSg2YOP
6Vjw9mk3d9ERhScgP8q+8/yVmnJPMLyCAww9KbqY+FMwSVea7n/MAcqWAAKsewKxBH3VfqfALRHY
goRMIKPyDYnp5jlxF9M7DNMDYC7w6JqAGHCQXtRph5ijNxaFcCRcH8/vDJlv+YOqiCEITJWv91tS
RiWZMnw1nos5gqCFu8gT0G2oW8s23Qv8xO/JMmmScuFVF3Dh9yugFiJgTbD5OlzAIwLYqLb0R+Jn
3Qibb3g9LHPuJWgfQOJ2q5KtMucZDNs+mYLB8EGk0ZrDBMRuVdN1q7CY4gicb1IO9Xf+4ZnOTQUh
8Rucom0P3NNak/Q7DXNqCIP2Qi3q//iCdLDgKKG1Lliq7WhXwdEpYzmePPXItlClUwe9lWFncTYe
iKwk0hXdYKIiIw8ix601yWmcRkLaOeS9rn36uemI1/ep2FOHS5XhQFRapHRxjHXPu34dUZmnvNsY
eTc4DjilYROzn2GlBD8WFRQ71YtLBL7VKMK9SYgfDS1ocv5TIqrrbqKZ8RFPMMfXEyuYPkgunee6
5+whKUoyTtwhB/w88AH7b/BzgZ1WlLBHWvVTF52/0CWtve5g7+mXox32xy5Im2kng2EHaSnHyiU7
F1ZLmttSS7U7Q97SoC/+zS/WpODTY0IXWCUJvWvubqVdX6dDQddXO6GB6OT66dQ/bTIg/xGSiXvm
gkVK7WcfXA2v/fTf8Zf/+CAIWDufUgMS+d37K5D5R2V4ypayefaKWmN76wT1kfQOio8tZWAgJ9pb
8rM1WwUnzk0N9hMnjywFbh6XUIgCWTOkDYlS2QwXPVRX4ofgb2R64Q2s9uojAX/WXjNA7Gtx3MCi
NsxzkYII0KoLM9ifY2gREtOUpKw9c/15t/VniVbds7cM0ztErmvnE14rIRtC4nDxR/rZ2zinkUa+
oxQaacGl21iBxFgE4sTJeGCciMcFrVRooKiP5adfk4Av2Om6S6vGdoq0cjVo69KJK8lcaXkhPaBE
m3KXJNCFFawgbud/Tp5qjSdj+KspEBCJBlPlqz2tat8MNTTS2tMHwptsqPN7dPXQ+8dLm3efGzT7
AB2FGMBvxpPctAgKQL1zo1Fee9pMMPOIOEILLUiQpQ+XtRvUkUjmsL1DZ0TE6264tMDifa71svXp
W/mlb3rInERs1aTbiv+97gUstCM+cMeWf4mndnICq+nDU/0ndcGRjJOHdK82rdKrPIjetoHoi5IS
BmS1TPmr/2RUvYCvrrH5F+RIlOTju/oca8wftr2x6QWs0wVrxoZTBOC9A+fP6Nkb0PjdrqqIrKBT
mpUxR2Bex6Yy7fERK8x+1tJCONcpOiqPxM7sw7kfXRluEwLHMGhXxXJ1na2HlGs/f80xXIzFBx6M
jihV4atK8ieWyyN87sfQ4TjZTLoSbiRE5vbnbfJEO0+GhJmAWCtMRnYggVZIFRfC+CuKtvycaYs5
wggEzznEfLvcy4ZJ9pkuJCjmWb8gFG5VWf5Eif641svTJSFbP/8BdKL6ODESnOktN4qsoGCQFHNk
ENa6RUT25W/gKlNWCVooUAdkfRN90m10b3q67PcEyc0kSeRZdkPnjj3i9CeESt9PmbQoGni85q4q
lpf89l/MHw8OA/M/EE0BRhthNc5Om6Rs7ZjbWEvEIjsCZwE7cY18Xax5LYG6qmM60NzQPaKXZ7J9
37hUwQh9rrP7dNiLUGtBP3wzP822MLVJiC79ujHfZp+1UjbvtPEk/i99avpB6N/NwjdK+R0yBrvb
9Jn4PKqWPtFUyL4lX/CiN2WuXyk3/wVC2RQoxofq/7qGUEzZVRdKCSkggGdEMRFC+8Z6IudBXgfq
c2UdF0bEJQvaEkCShVOwGN63EHwd118ZOnftVyE2rb+0126SdYn3tAzC4OKnBXcqPjvXQb3RGHTs
o3rl13WbZqMy+YefKFCSjMzIoCKyg5A11+z+8JEfJOaDUf2rH7dH76S6U3Hn8gzhq3ovSn09kzlE
7Crthanq4NLLWjrJokZH/ThkddduNjGBkWY0Cc+ha6zbNC+mkMYECUjoqwxDcP44JoDF3eGYnBE9
V/YskYbQ4BxrJV5OF3UOJTTp8ieHDkmNofrhzB6jwRQRinn/YQqC0A6iAKHDj8x3b4l1okTFxM0X
sHBn5MDSh0IKz6+dxLfPCaC7Fc1Z6/+oTL7Wmp5FnE0isOrwsc1HZ6pqPM+JGbzSj1swedC7+5Jj
zrKuYWKgCffQ/dBQz6cKgJILjb7B9e8r8bJkVxqpIAl7SNSgLuD9u/5RnXVCdLBzMUHavjdknkDd
WYomWUm8sQM+mRzGG6R6R1uafqFXqt5E/hAOFPVHdXaojUac5zYOWFELvRv4qgJNcuKgxCJTEe3c
2NbcCioZznZMngs+DgE663JdI0SFxrXAcj8bWEuLkH6UIyliYZfrfVgRyyYevpazqv7lUECTLPkY
yeZWRbPtRhbcQUWltjhGp0pXTBFfPYglYukxGpMTOJVG+JllloSFwLLejec3cI99lbKO2f0HBhmo
/nyzLoQeX4QzBavTO+Y2qomZhH+eW2VHq1S/sB/pw3Ah3+MX+1hzS18ZvhyUoFLU0PFJ+OnCjSI5
l2g2e65EQOBrd2L3jiN+WucbavoRF27Mss2frSiaV+ZEHfbTkSg20ei28NZZjXkPh72vF54Lo3Tx
PNhXUTH6r89qvyKtAVHRF8VhjtPjM6whKa9EgWqbtgiLZRQSIcgxOj24slZ2mmQcUrFf1moCyBPq
5HLjIiuzAwmN7h9VgEtrklfBTD1lSjMbMZu2vFaH0nNfLKyyDwHat3uzye07O3H2foa8bhHjyVIG
+YAYYZ8CMbYQmZyplbjmDs76WTPVhuCROK7TNRIGaEtaubjYTq7IMFJ6YcyInh0v3O8xJiaFz+8R
JjlzPoTJacIWzjexOYTRq87zicJiAfLF1kpT5jYLFAw7ijsDSkDXjCvHHNBPYz7yi4m2TX0ms33+
4yJem9gr9P2ItQzEyKrb9Zfaj6MuMyQSKhW+ax3g45lYyUN4VBIW1JKQ7+sUHdZT2GwHOK0tmGEz
KK8Vju+MapL9R9FOID3BmcH8f4aju/c09IUyj1tbR1FBAjR4uyzrK56GZj1UHBjCAask6hQpxN9k
Stdh4SZ6j1yIvSK/YE/XQuyXZGAVFjRLVsgqaF+UGSgzdVDT279imxdKxKZIs9tF3OE11572uSqK
B9wfBLPdt7ZX7wgcnRu27BoknvIz45ZDyfWVu473VoeApysEtkpwhIGI2unOPRtybl5H2Rx4yVmm
ORuXgE1EIq9IhWx50E/UvBsYY4qjYdu/mcbDUv30ZDAhHwxv/cfAUZ/QGo5Ld3bUpkML81H1aSY+
A8A5LoBMl4Y6P3Tqf8I26EWTDORSKXadKRDDYRPkEpaXo7RInj2VeCz8pJ2Bi2QkuV15rj0APZrk
eA/73SxuGdIZqBDPovFJmuwIyXjBt+ii8v+ZpdR7+wV9hdprUDhf2fh66jHLL+pCOFtG+wn3cH4j
YYnzaNcA/b5GTFMErIRadfovAeIpjIrsBeiSt+gw63bxbikZgDg2XYqecnUtFVVGWElWD3kgDBwQ
pxyYxesMw7K3Ajo2Cqb4h3k90u8x0VFOd7l0LjgvQjoAYck1l5IOcLth3+ZwEGd2fc9XuEY8K+Gr
ZCzfjAf+KQZ+ETsxwE65+Ll7m4T2VcsuudPOvxPaBCS9mQbBM0lZZrNywkC0sZtdiBJbhrdtiZCr
tloEU9xcHc6IP0lJQ3taE8ZCs5RueXzRVu52OYJpJTljUHoOETZsRNcr+QQW95xQZiy2tLac9WZ7
G9P/MUZkwvb9LgTj6vDaqdey9HWNSquPwQY6PAj0uRoj1UwEdjhiROkEAQ6bmaphs6qb1i9rK8YU
qlbSLxi19BE2spLlT4xQ9BiZP1Ccexn4j5iagtQZtmjia2xhaN82IWDJxrqr9KR6bO4DwUM20oIs
8mH98OZwbDzniSA9JPSIzTtrG4er3BOhtPSfoChFOdbzaUX7x6G1gaDzFqCmZL3fjV60DSUKCE9J
gFLHeDovENmgFPQMcJtoaMUQWAvDScazzY+oep5YkYatXG04AtxMzI1UMf/RHkceipoPLKXkdU7D
ISyDqaFqYOi4koMxJqLmhzBOezbAEd4x2YcbbBXX+zHpSCNBJemTfROm7MnWPIvwcIqHD87SGV1g
PKRZNZInS5TZTm+UFUP03A1LuHKvy22VyEiygj7Hlf0PbxuTuUJgN5zmUvi4QtYYrS99M14LrER4
0lyHFRla1D2sGFEAZkvO+BJoHJUH4qgEQwm+3bQsyL+XDifkyHNU3hy3NQGxbcXQkqfq2IN3aA0f
RHeWEOV40S8D0n/XeExNovEDE8eR22WYguW6+VvOxuKrv+tGgXo/3fGEduCPgM8aqi5RzwcY+B3Y
1kIqoDbWCDEwsqb9HhEMsfjH+3F//tauS+uD9IXeQPhPd6ltrQjcm4pysoFbIWguvQuVOWUXMqkV
LGYDyNqKzdk5K4Pz+Nj9x7Vi+wN0yBkAG3garTmlAg65HeFuRUrSt5ZFkWDNraysve4NTFsE5FnN
WW+YG+PFNllXvM7oLjD3tQsY1x4iLo9mH0oStIgf1XSrypuT0RELQto65vdme4FgwomhmnBYuHgR
BVCj+BxY0xHsqayCt+DAW/homNKsZiWhiCvkdblHlBs01epy9I0lOsBZ3DaRcfVfrUxiENj4bmN6
Xy0ogAlBIFBmohKeBldy9oYJBwEkKShp3P339BbP700wgFqQbliAXYbnKprCif7IM+yf+2guooKi
40CZtfKlsidQDGOIH7OGmswVKS81qhHevTngjZNGCTTi40/+EzIA4J3EZuF3sPJVgeaIVCpmg7vG
S32MbPs2f3PS4cezlh+UbW4+UzL7E2XejUrBn5ytteY7cWkmYuFA3fZv1CokKR53hrLjMkc0sM7V
XV/fmXTeuxAeey9ZeBFrilgCofUIYpGnMCOT50J+uI13sc0Ba15bPIJfb61Kdg0nBYHyPp/Ct3MZ
ciKPGLZPQv5EUmVyWpVQK0dBmpAQCj6hXHieG8JScLu8AXh1TFbow3BWO0zK4N+bppjEs+M0i1yD
W9hMRhepf0eIxRiyzqh3QcI3Ljf/FzWxuRrXiVp8kaxdS3Apa6BciL9QfAlrWkmbgFIL+S+l+cQ4
QT8xBUAmbCbFm1CxuRTcQnjopBK6sx6T2wlS+WrPysXtxhV/FP7sfTpdQir6BInryuvH5ILhgbpy
/xSQ4m8zDxePgwtUGv7B3PGTFdovE0hhG3aPjuvZZRSwRPVWXvE+L/0fSCIdgJCIVAqqKA11h3Nv
eKCB+j/c0W1dIFm6fjqbuHenmoea4EegstmiQL9n114vVrWaapFq5KYcbarJb1VDML3WT+rXGMMd
zgzS77Qmd9XZKLdIbd9e+71hWqtygpG4TzsNPLhqFQjd4w8dTbyj+mcB8eRZEmSfIvOAriMQgfLi
HQFHWvANzpR9dtoLhRMPbrEb0xhnPAFxfxaeB74EQ4hih8UbDNh3IvhWPdFao+xjwULDU/yKy/+q
O6XArddi46QFKQ6HKNOcCPH5dqtpuvgDwGzMWGbZgCwEyewYWKtRIqTeKPWPRhTRekXz/pcqZX6b
Bw9NOQxyBEiCFyDrJyx/wTneLO1ojD5Nth4TvWWB4VvYFlgtdXN6aL+IAIWHQZgd+6AZppxgmAcL
v6jyTGd8GcWTq4RTz+5/Lvk7CnQTuV9IIEzEbuNnQYRb/1PZK1KmJ54T6XaHesa1Qp49k2IieBtt
M+3mNp+JgmfRENf6ZYb7lt6DW5iQXJUdPZQvDCarAh1vQvC11Jk3MdwYmWSzni4lWkzgr3koJzQI
fJ4VhDY79QLvAXkCjMooHqukXthYxtgTZXf5OWdh9pQ2lYb5w/1zPYN5Llj+Fwk78N+uj5X7SCGe
efI9g12wXUCU16sDzKIBJKeB/GG7UOHLjLsFlYb1RnO1FTJb3mccWPG2uRaMivPq6pmoLQCLnve4
MMiHf3j5sOK9//aLbGMybZnFZLas0VMA4b7CDQa7SBXh9kZrH7Tt2Kqoo3Ds3pDcG78I2Fnsi2os
daH+ulgh2bTZ/quNSDbB1Y2uMbjix6stKVbZvaSw/gvf/66PxOwRU61y9uU7EJORyHZzeVk2TEjg
a/d3IaCbdkTnKj7UUqTjj1q5eut4sDbW7jtaV8puOfnPXEiQ3XhZ9gm3q8DNkcW51uY4iTRTMtFZ
jXPBm/I8408Mw9CsqeHPA6zO9B95XhMlRM+bEzn069Zlp2EPjdSmdk8Z///ydqhasF6YIlYHnzzm
tTiQkjTFmAo8azwdhKKpwwtdJGhFKaref+McMUWmt8hR0nM/NtxGdbwMXTwmKRb4PURgpKc/GDp/
WQW9+ZOYAPhCOvyX3AKJKLYR7YJ2jAKZM5rbh9LLOpbL++csdOMOSYhg521Qu2CZYORt+szYCmHo
a3HIzTS+L5tmF9VyFazhSrpg6D93VuRx5tPEc5xmkzFUFOJMbomiuAw+2IPfJ79r2WV7jB4T05CX
foB/zB0Rt4lYyMR50C20kg2KtlxM7jx7RvnZUDIKsDTHzN8CYAJ6yWwUt4o8SnrG0zBgzllEY0wW
+g5NlaraRl75SmhCcdezfoVm9MYqU8Dag5UujxBWNGIrA7elOHHHwzbWR7bI384zWj0KAtwOqxsf
hAKhfNWXcpQkzESSoAEKHcBcD1mvbjZxeLkVOziBx9ElNd5PBBXLdTqZ66C3MEpfpfP7U01c4KTX
Uf/ENEmfRn0wKLLOjRLJu0QSqq8D5riKH8YC5j7M9R2g3y09OKDTYXujXEay9rRpBfbh7mmWkHX4
W3beUYApJbCYcRp4KM/NMCEGoWyb67cpmc2/i3svzmtsEGchyYt/po0QOnbJwUdYqpFtox7YGjVq
CwmLPxnyMB5HjU2U3lb/8Y/bAE0mQDpuKm/CzeflR0asRl5zlappBM2iTDSsny4E9ZitmI+EGFcO
UcjYJku7NCTxnhtm99LR/hPIuqEBFY7MomcLLYTiR2VJyl1qHlOTYR9/BUV+bNNfp7Feq+STU2kA
EvEj9CDARCL2B0vDfwG7DltX/yBhFA7r9dM9aNKVJ1EeDsiFfLnQ9dD1TpqJxZ3jeh1wz/3RyhGh
AFUS4EiwehqgAauwJYP/QLWiSS9CGttnwl7iNh8ZWLYuUUA2GoXDtgS30YiLphZpKXnEEJdAE4DW
cxn0rldIWLwQaOIENSu6jNqgHpVbxv7G6UggoQdqLIhub5c8A+pxZL7FHJd8aUImKke+BWtVNhD+
ffnnhJ+woUAX5fMvnwesVg37NkCObO6Ix25RUUWMM/syqcziGkpvLKcR1DA7dJyMTlo34IR7Y6s5
XKflZFxmhveigF66Wv56DZBNRiQlKAsEfoGwAtCWORoZ/f5UCoh8OsI1FnPhtMWfPQiK4xo4gWjQ
apfCJe+M/Yv1mkWrd/rEzOr3jGXPngJUPhAbPglpvS3pwbf55Z9411dGnTZ6FPhxqgM/vgE396ZK
P2vWt8ldEtL4e5hugY3+boqI3/+7W+vbbzg9CBwRSFXug3yNpAvoRDouJFLCmod9EHpytICoscUU
rpF5s1F4MPTB3G/2539L6JvGrLnKg9JXPnQZB1U6j7YsvB8oZpbzJktjHMOxgntt3YQlAGnH/1tB
wLAGZ9vgyxY/m8IGzGqAay8t/W8ZrSdaNv7hzLGORSlZGO7eERUSSDXfPU9lxMwA8e0d9G6E129a
fS5R9UIF+RPPQGxurN37luo3kVDjk49M4qBPl2C0Dxg2CWxaqKi/UAKbMEFQbok/adTRxcBD/nmW
SZxt+Q0/24IkBKkAzU4MvfhM+smOXUmsq7vDJYZsqdanAZdn6HkqMMq4qRNvvqISCau2Y++l0D53
ThWECKdvjg55OlHi284bUq5xLIWHSN/VK+Jm0iMk3tvtxyeFBOsqat5M3TA1hvxApLN9Hy7VzjEb
ReoePTT61Ol5dsZ/5lJ8cUhX0zMBjd+sPeSGkmICjGlyb/mpwdnfAybgqg+1/6/0ha29bfxHYz8J
6/hynbYvKPDqpJHbPfB4FCVdRge0rm8MZq8VEYy99yGRvr5Ko2Vhzlqr9wKnFWTv0fi6KU0lHyp6
2MTC5Q30r8slWnkr12Bkcblpv6zlaQPzaOeyH8lybpIgwuGTc0X+sQI6qBz7f/eqFzctWGSJIuxO
hZqtcP4H9x7joxYOkHPVVcCACkoAYLnE0yVTyTnLR4oIJpY0RKOndDBUAbCPT7iSOtK59zAytT8R
D8lbhIBxjvR2Xw6jDIcZoGPIH4Lkll1NrC8jbs46NWMmjow+0YYCatz6T9ILx1bOcREPxDtGKOda
ooeAyUiZ51XbFZ1IIYc/7LNHlqsB5sXA72foY4l9+S+WKf1xVgn3WGDO/pJ2NM/tKf3j0rIm+FfF
sxy7UoQULblhIpLkoNbQ86YtXA4G/8aaE1fmjh2H4jEuKlBA+rDgS4NC5+6l1ym2YJqbSzOvxaV1
F24yYt8aFKyCBnldn+qTLJB/sugqyK/QmP9ZOWdNIXM7UUvFfEvxoJSzyrghDBUcqboW8wE82qpu
WJnN/MTkowStngvW5VSI+8dMTWnQkL/vGDqgB4PFyS0G1K5vcNF4hQ66Xw1yPMJ9xIvYrsVv5Qe1
Mn3aCWhDOG4TvY52yGTRL5LbeFSZyOczjassD8oIMCEtLYTlmmRhOAVdL/ozBzMVPAfLkGQ2aJxC
xPp4PCJ5q4j1vgIz9HHO9gt3OwgDqm/wej/c5soQd/R85Krr0FjRmTJ3C+a9YWah2EsOpT7iOOg3
H/Dy/9HP7j3zcxeqPlkGiogbtVmpXYyoUv9aM6/RmkTQWuvVCduXca9r9OJ+7NIc/xv1PtgYvmiv
CLSMKsRhRVb26ZrM+lgavr3q+9/ewJc6hW5GDw+B3lJpWToRSgfLO8NtOCqbBJdsJ2f9Ls6rOtSN
yXMGRxUOW0Ne0eXNQipaF9lGrqYAIpOPeXuvOQnRDWkmuDcjXLRRFSAcyS6s7nPwmlPt+npAV3EK
OFIHTWUZQnJNvVtBZ6w6TPT50eMk5CjOsl0egfC5RFyWqvurr8pT8mrdT5Ouh9n+/xUQqKVu3Uel
PDYdAJdUPeRF12GCQBkGogvO3sCFLYlmN5evma+MybsfGF+cGwASQapZPRmcvY0MSDnf1BGdcuFV
sOI30E7De3qH9lG1oLXApXFB/B9irM0zw0RztNWJzyL5rRyyoaZp3hlr6rL4w2QbRBv4VhBdZffI
+RJ1uclidoz4pCxSqTmVwKRFv/z7jZx8CzMOIqd5gDrI1v+p8MfUMv1RjDULTo+npKGQXgxRAmPl
P0QhwrCIxrBKzkNpvR7IKY9587Xtl3Upo5VM2+SSBmhvXR/YaOLxdUZeHXpCVtUcLzc7rR95jWBi
lEG3R4n+6LSFXvhd4/LnIKLG/Y7RpmMLZCF1O358cOadynkj0GCHncoErTpy/R33U373VYcoTEtk
aJeR7IEy7zXXH13/0naBAIk+AZAMaZPZugTcDvY9Ioj+8/kvR7EiOuENBMFE2GsdcKRTKCbeom8P
dq7eP0tlacf4rHtKEsPVdJGDRHFCesiFknJGK8YwVbhSkI6iRQHE8rlO7Sy9WO7TlU1KRH8J01hZ
CrUj52NI5bksdyMSywaCtzz+qEYVU1iJp8aXJwJIYBo6/fVVMJIG/RrbeO2EXn3002chyAz+WOYK
2bRAs+D0oNGTpiucLBIhKPF70knOMaRA+OXbB3J+/WUYqR3Sv+hyhjVFZh0QFF4bANzTpYSSUYiz
n50m/p/u6JvOVp58bVjBxTmMO9vFrluEqhgzooangPsv+A9BF9dJeCOEwPMKOkTrJL0nH465VCpi
OiK5vgiS1LVudEaUbKhE+RaKBEVMuUx7YvSvAJG9YyE100pUUJcQJbORObIXS0UIt/1ezX4eOfLf
eEzrrnDsnhW4e6O4US3kc/gsJ2nuyt93J+nlUH6hpXMUBtYGbitJrsA+5gkLr/u/vWjLEU4Ehw8J
FjB60EGkGirIiW4En6Zbn73eXEAgz8yaHUcr7qfRLG0WQJfH4WYu9hg9Ddik/hJrJa9xyXHUHyQK
sx1cM0khJsdFRjp4g0OCuUXAbNa6f86ZkrDhpt3MrzVNpkCJ00w7xsfjpsRKJ2Kh+NBMtwCZyNVN
Vh0dIILhdY8M0d6/Eje2/q+GWSyDPYINKeHR6s/wJPwuwpFp+dS8WRVOq+/YewJUWM4jPxLUx8bR
8aDI4DOweRBJVKp699HFxdwbzxbO3+QzYvqGtT/3Pd8hehp836FOawZKmE9buMlyckSj4Phz2UCd
NtY4Hqq0OiV6Rn5/PllzZLEvWWYwaahzW7SvHGkEdjmOkAslvk4/dK53582oxvHOrm+wwawd0lyl
75n7Iqd/hLo5EbPOnMoLZrj7Womr9vVh5OIz/5sAn5ou7MaqhRObrnK83mMvgknmgW78V2wbMxPR
3jxQhVN3AkbZ0rx8Cs52I3KO7DTPCA1I4sCmDiyt+IJ36+dflAUXm689hgqRJ8qA/Uq701N/mcJd
S9mFw6N4AqpcmSUFzJg0hZcFhzV0n7LQ6bA95PvMoYLR6HYEpdTLfE2mnf0BQyBg+sQXrVzSbJE0
FiuJDaqBOQoL6LzSh/KXb/LnGm2mWVmVellufsuOFPKWCquTBq5UUY1Fk1DQ5mzOHoFN7O1LiscF
9ksGWM6ktHxZ2mpAju2opZhLYTYmQF/6oY/04jk2SZV4pWfu6qumrBtsD17w9eRaJRYyjiP56FKd
6X6z3KQ8abvxRpYaY/HvpHBOBy+iSxQMEJSzJDe/+VuZ92e2Wyl8DLKON0ehCQ85igD7ZQX9CTGZ
j/xC3Sm3K6og5vdHYyHTqwuwXqKugvmkdCgwA3W3fsDbNvHQFj9dYdpUBPWcg1rEsXpkS2aQ0eV3
WoOTzmvb0V/oot3o9OqnWYNwuJcTTcQN6IwQ1YEuXWaHzhMOF3DyZNwIn5LOR61im3Qf4qPaxVVS
uKSgKF9PN0G2pG1o1/cpqamRNO2Sedipi3yp3vyPgQ1vbQ5qUlCpkzqw0Yq2JMsRGDuxXOze+08F
bFMghtOkZH/PXSTfXIa44f6+tpfpHjNVixVnR6vPz2OS6Sf0fhMQQzaxNsCJ20f7CW5cHWoCRj05
Y4pGOhSGGdD0wjpHk2LKMtcw9tjP80cXf4XiUigN/TRO9zYuWyZAImOFos4Pp4Qzs9BXh7Aqnh+a
ha32B1WulGSOw99PcesLx2G9Uu61BPQdkfCjbjmz2Da6Qk/DCoD/Eiwr73jHfqH3l30hxiavKd7I
Qetc14E4Aw8jQMBEC+3mghgoauR8XrR8OLGUg1GEGK3YgLDuiWwoGRVinmtff+XAfRRGR9/HUgf9
5hKIoXGiwxevH/iXNT9bPpQCRi7hYAbk8X2FHGmW9ke/ajYDRs5zEjhuBWyY/8O2Jo45w5nrAuHu
Gq8tZ6h464o6tkH5RcOSUmr+7S4qLWwSbH5aZ+dNJSacCEg9/HljTHdksTYPUCy2b0wT9mqnimV8
jpSeWsyqx4ICW4+KZQCz0++4bwkwJQs5HMCsbgnpmIIGLemt+VC9kysUA5pXtuekNSUevRX+M/NZ
SuZ919uFPPqLwhb8o0evd2LMYEVwa0iBqbGWmPoHF8AN82jBPJ9c5D9VJHGUjya70TXYZ1SX1mSK
xQmYm5/9D/aYQfmUpctWwgogO4OON/ylvq70bB1RhCZLEHPL4AGBUJSYJCwuyE0FziRWORg/Nvd2
poYx8dkROuBXEBbeDgwXjGCbL3UdPT5+IPWnJIlLZwNN2zNWlDc1P8GtgiJrlXrkRhcy1hoOdS8z
//umUnUWRPXIVzf62+37ZK6RIrUe6MUfpyR+zKHmCQ2nszpCWyWqXs09rrdgkdLmlecgfnl5QQf0
C8Fg1iOBlBKrtlECni2SZfIET60wqXz37SANF1vMVBNOz8Nje0oWa3715Re//H77+GyIYSsDhgBu
RAtVB6C3XBcMu4i9I0gMbzS/h8Bc6w9Rs33H3tzuWKiRkbdOSBugNtADcaWnroETCFeH7wQ01QYX
38iNxr2WNTeZdJZfsO9McHsY2tSf+Wrs4YVp9SL/GtcabF593AQurtJ56HOl4cwfoNabNmDsLgm9
sBqwH/jAGi6jSCVnr/f0kzytzekdg0aeF4AmlkwxaVD6B+j3Em/Cx/6yuaVeb7DCI7JqALFGWzza
wj3eI52L+VWkWhjxOqB2ktj4xi6f52lFuU8ACSAStnEadBU3FWPxQvBMHQRs+8Vc/BuLeceoAn+A
ZTxdqSIouSMdWPhycDzE2L3bru7kjcH2Js2mHSyDFcX8woSm0QqMxOlKGM+QMEGu7Uwdt3XH7zLQ
3+FhqZUQJUoOQ4to0gc0WQfxNRXuSCA7XGmRKj8MYf5cA2rVsgcN/rVQUkzKYr55ZC8Y/iXPoDYs
RJn2IIzDbgvbh0JLr/heQ5nbXgA7DFjqfpBi7sQQ8KCfrA6UdjmdeqLDNntubtBGyr2RGiA1qAq8
QROcu71y31OH2MrpHRpGSfmxAVm3Sj4oDqmjCeGAuT1/GkeBBUnHYXlQlYKYeEvGWNnlRS2v7D5o
5LtKhi3HH5df23P/wv0O6yNiH4NxnQM2NKwK2FesB5U0AsASpvjWfg4oYZPzYYMzgf9hzI9bLVlG
HpK6MofEu2m3DKZnhUHlvANK9zvqC2TUHob8IvmIVPJikViHt6XyQE6xbboP9nN7W4vheUJc9FdZ
CLZFu6eTkxsQb+e5TvY6H1lickbUX/gci2scr8CrYEtjWiO8VPl659GrM++8BBFmhmbt4ZeesA7s
FZTRZCHVwgNcxn/kQ+xGv/5fKu3pG0PZqQZYdIFG+TnUdv1Ds5J3MOj4P7FtHEy0wQNfIJtwRgUE
Y9HM0iRlhwPk3vpr/5VJPI2cRnB8E4mKkCU03u95a0rw/Me82MTa3itO5bi1PX27m4yXcvMhf3l3
JFOxZzONPZO6PphFxyKcz9RbH/YxwYlRjwIeDcDxSX+n+TUSO7eiG15cjoULakbymhti+OZ0ZNhO
7PJ7H23TtXp7HPjVYrtDS71hSohhvtVqREG3g3j8FDLDhFyN6gXyThg4+16D9QiFmkVZ7B1fnEUG
lyPijUnd55m3XTiHSOCdonnVlPnseKfEjVwslBux1Ff5TtXf7o1ejv0/1W38SKWba3jhTmFcKEvl
p3GXL4bsUxMUm7ovOu8n7oIYMR2y9rQ+zpX8xEtAwb9y8zPKHFfGZiD3D+RieFfUw8FeuH8EpHp6
jH41Tb46rEmA218K8sqJB8X2UiqiJV8jvy/oP+YATu+IsyHYz/4x0E+Htk7KTvweO6VhTHnPg43G
k4jQDrYT8Tv20P9ZgfOf4wgT/TKhfJxwOQIlgn7SkoEVMuf0wD/MUj1qi0aoJ/Hmr2MhBZSQqDFm
D0e/ohKfPxeDeC/N7Ear8+QrwM1FVdIxwayhbnwini1TLEme7WppIBdrX2WzRygaF0h5IkzhNwde
AzDJrH25pIseFNpbC/gQ5z7RdeGKAEK0+56kGPYY8TCyt2mOfzDCFmdR10DYJEO16wEckM/JESx1
8OlJhwmCoIF+7xg2Fkl8o+89lCEZIaLSQVBrD9OG/1x9P6RlfCMOxaLwDVD2/Q6Q7OqhvNtv7+Fx
twmp+bqMqLF1xj/2Sjk22yDqa0tZ5IqaEFX4Br+2M87Rk+o6eLtlDwYqk4e8+7mQdx02sKIuu8iR
RwNboKZNbTYsWnSWh9Vt5VABfvBhEQSlC6BP4N0bsU3NdemHI8AmtOLOqPFjL8ru48m3SoXazSyW
SJ/r7RSwlIr87J2HxiMAXbZtJ6z58W/1vsPI0imAAkwjmSIsHyxpJGVfY5VTSnarefK1u4zM5HCC
jxPyDxZDK5O+2CNyr78CMOxMu14v8Glg4/2cl/AsvUcFLoJjNdpRyUCpqi6ckiJ8lisOGCezJ+gt
8dj9GrJclOZKmPGQZwSt0G1eJqq+A+0Au06+dTN5oBr4dFj78djzAzxaOcDoW0mfInDMcl8M28eL
l8t6fmU+UKjgvsGZ2Hf+2hjdOlhDT7HkHj00S4N1mFflk9t0standwRdnI0U6kSiczGfeAcK9qMS
PqRIfajHFCrX7tJn+6Hn43LsD91xwducLDnZa/qJDFBv5iUvAwgyoiFSNab8tTOesAmxy0MMZjO5
yaXM66GGSuneMeMlXV2or4pZKlRj5ivXBtsvVGO/cpRZgdSlhzUNJQz14/LVFcqOrncXnLjT31gm
KMrVfr9Dy8XvXIyVQ4GSzYEtJx1OLXSWezofiM8xl8l811ToTXZSjDCbZ01R6lS0NdegPwq5eilY
rsYkkvDW/t9H4jTvNWK/QYPzjxvVbGXr5TlZL6PngG6NZkVokgzU/N/+8qM0PslHhElyVbE7JCWi
pCfTLnpjmEcXz1AWcJf9zL4HVn2CQTGffrUunDPR/mPI89VlBkP7lGo5qYdn0z60z018xBEtjd3F
84MoY8LwzzH8HzouTY6l87qdHxMJWpBN3K2gsNxTQ/+j7EomknUze3FlHiULRHE/Q+uweScm1uo0
HtxH7MhnsVpyOgFkTNRK3I6MAQ5b+ffEUltxjlV11RwRDX/jbD5Cj/Msj68GXOBodMjaYHyIThPq
Ta1y+mL+WOUon1c8B/us3whULMwOuDZKkw39hM2I6bvEqJHxAafNjYau78Dn3nO0/LKaIRpZGOCs
2oC9SFCnTA8N80qKJLdh1xtz2sZ5W+902JqPSMqSGVhiihPuVC3kggfyIEvTArQf8gWGqTti0T2S
qxa2zO1GrFBuOAviW+yLzw0I3uxspy9PCxTVCfw21qqqZnVBsQmAfqIB1HQXURnkSsZQlRPePxWa
G1ks7QZbSUucpWqtjpwMHyFEHDt2ShiFrK/wkZ8FiC6sEf4YNKs8SGb9tDCIfImRt1UWrE9Zklnu
UWFqDT0FE89UE+/KPOq3bqlMb3Zkwoh1/shMK6dmnUcSWpgP8N8Df+Y35pcZlmohLSK4ROiK5s6P
Lj3oenmdcQwjFTyvXKDlsKn71/csciQWIbj2ITW+DgO7PSY1PAG3sBjzk77Vf3p7egtMHYh7B89X
rDLCViq/G9DN5sVw1B1WhvPMqbKgKPjfTMPHRh4vyfqz4FCW47JwGfBVOnJjmUv9IJ3MHgybnJ8W
YU0CE+iQXFDhaFq7eSxll1S2PMx6MFSOX8Nd7fo3sOXZRHGb1YoaTPnroRUSMFwme0BNhFcNF6Rx
QPMUB73GJspoDT/CaeQWj1DQctNqvOFv9udt2WzGQ85nqLs1STm3OETMTVYfURaSfa17mkFDiqlg
ZsdZChso5+iT9SGr24QghUNJcJrJ/EhyGrDmEe+aKqO/98f/Ahqc64BqpW+8uGjv+EEQGc9YBIKR
EUGrkYANTuk5+yR+qRWw3mTctvA6fHskiZnmgJYjwWcoPkL4k2YFbqWEEuFziGwDvKfe/k3Mb5C5
xL5kc3XepjuusEd5v/lAV0icjFbgpDWJapw357vwdOxrECbbEFxSQeLUEGdc4Y9gI+gEl/cWpawe
ZShnAAVgdMyARAoJlzsGOoheh5mfwBFUaJpbU1lzy/T9+ZNY3lRD+b/o/C8/HoMKZulIiTCjT/oJ
nSDqQumSeshUt7Cn/9n93goR+zHOwY4XvM9KnMSEE3XEFwIiGWbh8/R3LdPDAxgQd/meB7L87rtf
67yS5m/7TnON/Qa6+kpDomqScF8Q6UPX+5vgTa+W2HRIxHwuq8RucX88jLlqyyLKaVbJ+VlGV428
HDhtHdSd2IsRTQiBKaP0+6tMNN7VhYpU5LR9vlPKLdcqAl45jXDWMVCAfPcgJa+h8RHs/v242v+z
QdP9Hyzw7BxwCOfG6LiBZw2qgf0DOISikmIv34ZglgFYyUXfQaQySHiJ/ioqIahy15eKfzrHO0i9
yVrkNryvkVGKL+YgZJw1fNczmnUihVSg69LQ4fRkYEzNx2ThN+YEMVotG2Q2YM7/qjy0Hky+4hZX
eRpYgwgeV2F/n5Au6PgfkNzEdZXnLtPFVkiE0w5JVB4XPyiuPzp8ijbUmoPvlj2bqVTOLAImcfXK
Cyhx8RdB9i3ZvmSG0egFhdNEmj+Nhj4yD3ySAARv1Dycas2sQmSy9PRJ/PcAaalf7Wbh/9Ai/na3
FLA/lrWPNAa8gQVOM5cKgFfD2Mc40gPlZ0F0+bJIrjprxuuan8EwP3BB+t88ooTKEaI78c3/Vaex
T4rXDsf7ez+4g363IdV+yf1PnfBN6kGyy9MyJZ3Dv8BtriVzZM4kfMVL266cAp56MFfu0ozL8KIk
zTEHFcv2AiYSP7Q1E+qFdleAQzZU/xKbyHPTYNXLlRW0gpHXxW0EnDzgagdA8oiLkJ7RHR66Qwfr
4ub9KUhLhKEGs+sAdvLVmMCmbldTA1B3k2V5T0/hZPSuNUKeRZPmFc8mMwo2KaRirRL/UtHim8Hx
5S5lIrk6Z9GVmQqsB7GJefHpDse3rnG8juSEy9mO/+mBHn84xfu0v8lwXANaOHzs+yWh4O7cY+ND
FP3HsOICRGkrfQM6qe7D/3Q8w0Soiwykca1INo9fGx/YNuaOqM2/gF/AKvrBZjFXwaLl4AIi89q0
pOvVFvUmi/OrBIuGmg2ATQfBU/CUvCDS+oa9iq+b/tYNckG2BzMWRwYF2jHSpQxOtUK6ce2wmbgI
R8K9HpuMgFWR5uJ0xpvhbvgOJ80eWo1n75QNUb6kbi8oOijMREz9tPLOGuM6jLvI5vVITZ7EjHf2
qV1fz/Ae+IApdhZ5xiXlctDD/LafoEbYrrRYxXqV/WTScVtNG/N6Rog/qfoCunKoLNV9gv9AR1ms
ua/PE/SCl5pHOgdn7jaIcAcoJj0YbSfmTfFDRgSx15GCGOpMHbVMW7ngZ6RYqS8UuzeVL/hEd4AF
mxL5E8g1KJvSG+7GIrEvjmoOIKMScxCrXJ2FnRYeJct59RQ/1zaaiLh9u1P37V6W71dXY6Mdcr5D
JNn/pNf19fvx3kTyPcmuFbU4fhagDPObL5lk+9qpMA/vaKuJfOZoCkjSJgvmKlPPBvlf9YrUsTEK
eeVkvOPi5pvXolGr1HH2pHtqvijjP7Hmthu4S5UFLdlzTKrlOV6GAp/6mcRgi0ZnE0qfgPLioO9J
1wpNFYuH0DZyNrJR8MI4udsJ5D7rHULucE4tDTaKfMA8jEWsXDWnhctjcaPEW6wd3Wpnh/h0DYmX
bKzCpbRe5X9FRdDChF6KlKb4Ib0Qj0hMA0jlYRzWW6avv9tWU5rAw8LoyuSlazbgSG6pdG0kZ23N
zTN4TPvKhsBoF+LY0pPSX6PmNT94SqLkR1ZfX7uQjNWPVzOE5Qx4oXzr34QzuQyt4eGqtXgwSyiS
MeIEqyjC6WfSltNie/MoQxlbo6MD3Pfpy6eWZBbrARPhERX4gQWlGfkakWtL+Ux+feSr9eOJINkg
gLvRPfhO+MDT3vlik0c2ovF5h1I5Mpz22uacKP/0uuePZBYtLaJEQdh0D/9FOo2otmrPyF0Vxylk
29YDVuuFT2O1+FA6KljwFp/PxJXQKwtNdsKk3HtABPh48QsJwxiWANLO6aYSQcmfMTpNceX92zNm
uyO/uZFBkV+moqW/2OgotWC3SOR0H5vxvGTZIij7DW1aOvlrzD7xX3Ustvjj1rL7Jak6ZbzzpfOr
vVbpZ4tHV05zC42BM+sWYwXarMZpFhM8hJYwHJZHJB9daIQ5YJOSgXx63DkTlHOgKRMJyxT4H5QF
qZ9B/3ARkavwgz5//Uw6toQBdmr5owiBN6EVz0Zcjs2mfvC3Gjgcl1Z3/XRSbrXv1v5Ye/2eSsu7
d+RqQHsxHSly9fH7EubB7x9x3oRGo9SvMo893FO76GiC/TrUfd6Y5ZAOIZ+oOcHmNzzf/RjBGv1f
eJOqD/c11qD0J6n82N5BKq2WnrI2VBTAMU6q2NrqaF+hRs+AG7rRbqm3/UfozXPujR5kKwrV+h0w
pQ9LC14y/eO6ZsoHwN8hV9B8hq2h09EH/Rre6MKTtlNsAvP8AmWy8CstGHGxDrbX+la9d12REyL6
CvCfrC8GXkeWSFKnuNhb2EQTcUuAT1uQaIKHm61NPJlqhX9icvAjHcgNRrldwcBR2gytWx2QebG5
rzGqMqbNk8NRtJWXfIu07ETdIhGVWNBHmwO5xr6xrW/s/obhcFjpSiUFn3NTBRPKRTSwxkGhzG54
KNCJFNZODrqSMoeQlflsyJ/j5j9t1Fbr9FF3HabPVo2XM4UKUvKsLqt5pfa6OpETtvyOA+xRlmMK
MOKz8Zuxvq5PVmFhUNuxUtyGs7rDCjVdtVKK4X/hAXRHJOgXLDhONRg47b77msVIY3XAbia1VRh4
K6DxCuKk5Zr6KPNHHCIFM6lLVfOy47pWZ3qDW7/49qNewWINRJXjSPJYtrFyVbZbyfYFiQD3GUJl
KkrZYmlA/8N2nrrz6WJ+m5sBcbeYh5dMjznuSpn9tDNSyf56wEKbPZB2WByhz38fzKJPhVVxyLtV
es7wodeBaQbEZQrMofA1r4E+7MD4UJqn22pArvX+dpnkwEA4s1m/TW87XKD7Vd3EnXYW3Hkv7Pgg
ouqE4jwyahuQt9kzd38WufYYrbuUh0T/esOy4hcwKbhx+NvXv1BQoBVjwvzzxe6crVXhAOZrn+8W
26JnCSghBSD5eZBQf61cjjV25hHgbgJXwmtACI/yfQdOqyF8jrFtdGhiLnImtdYz1dNYtJcDrPVQ
Ue445+AQHZjrQc6Hx/52CXT9gL3VWSV7yjK/AGgUlkZn8tI9lUf35IWvLbLrsv4f9dNp6mH97h2U
DfBYKFBDebwG+ixhqEupGpaXu6dUOi2fPZ646w2b77z9pmqSr+FZio8Rnr5WH23S8oJALgFpkRWV
BExIwOzjbZOf6PB2RRm+UqdyTkCivpahF9E4mPeWNLgWkZMyRkdXJTVfSBgSFp847MlcK0JqcbJ8
6CUR9JFlB8GORBUPzFzk3x34YkJWWOIKSEtnYc2Si424SEnypA6cSZ5x2pKFhHCYUXPU8yfz1Qjd
mLC8U7do3+GGdXPBnmPrz94Eb9qJhw7zy+TcekUbwK6fyJkAf701vD8HNbjJVwQW89ebozdwfFah
3Gcu26iZVJc39sR9UsncoYsvYCYEMBJeh48wGs5QaWSZz3ywaO/7wB9i2vShW27hBOyb3xQG9sBR
X0nMocDkk5i4/3Mys/ZTOdWCpdUk7PmkK/DVmg9Q+UYZq7QixcWLApaRACJQGd+GE2aEgSbnzPxK
7yGnQUXoJ9iAQiFezB+dVWonWBF9i2slpYc49tgDYxJ1XnU5md4ZoaEA+RsHt3RXydeHo4Z3oso5
bFf83ye9WYu6GrC2tU0u1Apxjh+DoErOEeW3oj00ysozgQacXuAKdYInwlRDnwwSmDpbmRHy+1V9
IUpPkSsc/2oP6rN5Pe/TePkLMXKk3+x8pnTYyGmjXkUi90TdQA0S38ic4/w16IIthd+8u6SYtGaV
Momx5IFGkprKl411RTOVGvKxcOR4b+eZLCyHB0+A0w5Cw4rbRLecEKCOwVAZEe9jtU9f/RPtH5V6
ioruPWGMNyARbBoqYEmt12g569O7QSK6aM1NhC3y5scAchWRMbUncaxbSmLMITDOvayizSKt5eIA
qApVdnI5pLI0ASwTp1KhGNGKhOiQA3lERX+JbF37h8VxeS5gno9pMcUNwbiLEuavZQXq+4Nw0NT4
z2hOKeb8PDbK8yboHrRZiHZwMeols1k1siGgPeyUJhBgHaW16OXZCPbOgxTB+nAMFWNn4/Jm4tAo
oms2fq3N0Zcshcz+KUGCxDM0jbhbVQBWwIt8UXRYxRtLTRE/Cpu0d44UOQjyoI1aLEiY05xWVEI5
GL/iYG/o95LFxqvziJPXR/GXOIV0pkbXmes43Y0TmAL2xqHf5vdieN7ejlu5ro0CpgLfx2R6H2sb
VtwPh3PpoQWSogw3x8vWujbZwGNVF6ixNaOblVO+aCX5Z0MwQsuxn/N1xZyMwyhsY8LQD/eRQs2H
ZrX03lRQ9xy6LvQkZYjBeTKr9H7uhUfRxzr8TMjc1tss2/CRyyTc7HLYBvZk/B4crmSpNLCrCe3E
/T8i4d23gas9ewuLhXUR7ZQA34Nvs3F9arl5a8RFC4afy0OoVfdsif+FujFzC/ras++Z6V0Q2OjI
/h/mtbJFQs2eAdvpQolMakJajCiq3VzYTf7wDhKt38iE7xLg2yQ6fLvecpfrS/jsPuK6ByTnywiu
UU/kVf2OhKCjlQUwV8t6HlzBoEDTvD9+PohKotC1lUuJfaYiNOEqAOIybAQT8Y/8W3Arl+Ib77b2
Mnv1RvoUAgkkOLgOcTjDPn63N+Z+A9/1AKxgl7E9gwqRyfu+9l0svFlzHtP+ODUhD5lo/4Dk5bq1
x/zA/dhErEw7tW9YqHL2rtxW+tUEPoQcg9PgPDTj13BKeHYDoN+W3vWldHxGGja9/wSEnaXXY2rX
hl8toEkmxK3eSYikgeL4CylYsVuR9QEB8lgNfnG8svZAxeDpVGl+0+T8U+xpq+fO+Y5Hqo55+xbc
80t4sPEO25YfkcUIs+Q/SDEmSDyJSlWvavTSfEqp5b3mdCL+KcCEeGiLxlH1EgdwsjInnZYvFDL3
8R0VBX7hUIaT2i+2z6f4GZJvDnI1owltgNhqxfJQwFRjKWljUjOLtrEANgLHJuLqle43rk/vGNZt
50a21VnZjJHbpn0m9EUhqPlsKlwswB7JG/73bhOtv/7wkuJw5+ORucvgHlyvN/tKjAWIu+3lLGUO
xW5lwP2yMCuGzVOG7RWTwDxLPp1fOz6mZjvu2ps+9XzAjg496TMb2UNVXB+iQKlZYqFS+adAbgFO
AX+taScXU5BGP1YAN2J4fUXK7ap+eTHaZSql1xM8BVROVn7V8kLLflHq3zIhKZcYc516HNTBWshP
xK2gPmbCviufgzmJQ6cW7K+oTN+wIz3x8KLH1iwzxlYXj7jiP4LpbhQi9XuR1A9vTXkpSgQySBBU
6X4Hb8CWA/SmfJskhdFJfC9NkhFA6Bp/Q22E4Ga2XPzwrhsyerCWkrpuOt0KZlxOxkrDPhTjBfE6
aX9t+6Nb5MQIuEFE/iiyyLr2snYGSo5YhViWM7YC+rOwEn/Ak4PaQOSnff+xQeprXrG8gaOgPo0n
v/HlPpA2zkO7ErboDL5Kwbt8ld02y0ZijOtIX3DZqXK6+husRJ6OSL8Jup5qgxieOZEXKm6OBSXl
rOsfz42pAyqjCARFufz7KqPWNeYwQKuiQBJr6sqwSlLe02aE3OTIRx5mDcG4p7sw1W/GLjYt6NSK
iyuK7r6dwJDdgUQ4PSL4EIpTzm5rye+7pkoFxdJwelbRlFvVl/BhFj3DUpg1PgYhLAAvzeSALpoN
PBwFKdznGH6Diz/Xpc/f0fmnR0BRk2XCNtWqn0XDgN6HZzGx8ew51VwFuLrIhhS+Pg8keLm7ialk
ZzAhKTkiGa7uTZ0fRaz4F7j9UHtE6m98bRYtGnkNRwAiRqE/sybzrDxY5ZxRtbYgRu+2LKzfgt8s
/ebaAZIBZAk+VtyLDN0vthW+XGuYOogvAqYgM67FH4K21mF8xe7OjtLwpR+89qbtav+PDQvCQtaw
yn3vF4x7XX0AzGReY2RYMVIK1Bzicj4dF96oKAGdXJzmDEgSfDaRF5RqSJhKDeQtggKrc/72H/s6
cBX1boohCRpDfqhiDTJtSmAQKcrcW/0AWzs8SLy9mzpz255GlXUdNKjiXDY6f+gjmZXMMcJ1jiyD
j8sgE6Xc6PI1jv2VmBZxgaDDdTF5r6alQnvdXF7XG3LqQqrSGxMVz6KAQUhgLjOhEENBnRBUtyjT
xVsOwUlKrOzNXKf3wRWQyy4Esy0sHno3TftZTsQlUdRl9e/1fEFaW2ESeoXeACWf8ozzgtItOS7s
oKfAyNvPQS9P3TreRKwBmoalY2Dzs6iLSGs3lNoZ+CMlQXQ6acdUcZQUNuGz5EY25KAXmr8yQKBz
sgZoiLvuxyAKQrgEAGgtpa5wbhcmhQLIyVo3kT78bzK0Ug4BzIJoYdholse3ud3B9itvJoVMZMMT
TgyFPDIuAugl0K7Y5NaJ5EAynC2jh+Q4Z9yBKtNq3LJstyucey+RWVxXskbBYUmbFpQ2H0C/9FIk
vx399gBTSnG37y3QhPjxYPGzrzI23I9bMoX+ua9xhBa4WtAI9aVEf/hkT7yWxXu+F3rkZIpp44x5
k5UCRBMJnno2+nxhotg6r6aRtUrzspfVlMenA9/64BspwLJB9qMd30tKgL3rGAy64JwJeRCyE1vU
NaLPnrjuToq+jxjiohzluLRlWHjOrDr/9t+4ObgMRHPc+uIsY9LnSJ5/8a/+SAO5M52sXhFEMK3h
bwwsEWn8TigaN9miFvKT/z+GBVB0yBSt/0D/Cff2WFzN6vY693N6mkbyoqF2M9S75MwTsPMu8pWy
0mSLoJhpkEEKk/wgSYti7Agt0iAcyQ6k2UTh2t+MYeNQJ6Fv6wzf/qN5oy0GZQUGgPqJG9/omDtG
3vukFJMTcJ/ps1BBmpcWeqO0oIJbll9tXkwMGTLFWOKCX9Fg4/f1Nu3yySQmAqgHEQ6GJZnl1jaw
ok75euRPPO+JZ8lv3XzKmJ+i204KxuwaE3FYdAIL+LNNXmQleSrNt1EUVdkeDzE1xI4bsbTsKbr+
Xx6a4PVq+FkLVtCO61tMql6jANqW7HhJ84FYCd3uXnNBZMAeqJJMuPv5i5+BvPRw53vdVaHvBasf
IKZOL1AgovPKPuahky0D+WbjXrvBjqPvrAkBRW3Vy0FIWzTM3MshErp2I00Js5dXcbkrf7Hy+PWy
obEkKBXf4kD3rLZsT7VG//nUm99yjVMGj0yHLiG71g0dnvZ+r6vvn1kE1gzoQxQXsvSVeiuy8Msi
t2TzuXJjGudI8YzIN3lk9fc0Z8cS6LlyZZBh3gPQHd9Xrc55YlJx24J3UkSBQxru+BpgLImwS0Rn
2nuUAf46MLJ6F87x5lIlV+D+z+277/ye8cqgKAMDcnih4nZ1uiRSKdXhfXLWapIL9pFZc/VR5Wz3
c+cpAkcU19q4AhK04YTpbiOKMmJT0kJy4wxVZ0+RqBnxs2cEF10M/e+Db/zRkjE4AbIlHkE6yKPA
FbSKy9C1XtdPn2OplWoIbj7RprAJmGRTp2nGdzhKZkTwPh3bNjvyP1GndR13FvzSBCkKJAxByGcT
SYVzVRYGhsBcuHiqU/BCL+homCoBCWNzDPc5of7zAPYkwfgOfEld4bcAKrM2D5MIHtQBK2fdg3kd
YMHcX4IxOMclnBqEHtlfbfkuVY0DTo69WM+98HBAgGfn1xBRZNeJ8JsQcVAKsi+oZXHrdtlQ0Xet
5lNqB2rbLOAt17VMbCPbRlgaQGR2W7SZTuexJOPyfsK574CreAsGNifx5ubmMDB5v7wxTYjlRpti
EwAZTTf43QWubcxPl88h48rvRsI6IlStDghyERf50my/yuNwfT+SuNLa+QgbCYbz3XdTNNwDoUKs
4KzCoXtX4rYLzsuvlsy4AL8VFfABtSf0Pj4B5Sve0Ze/BupDlx5V20s9l3+XyKlH7LISg9haCXjv
b9UXzNdSiJds4kILIoSt7WGGobZADMhskcDvPNjgvVXO7Im43HfwmmpGCyHNl0k+8W57omfWy2pR
/5n0Oyv4yjUO15enhwtR6iRkpCB4OCQ1t+Af3l9RTyUfcyVVr3AiSGWlk01Agq97dQjJhBAY4AY3
YjFw/zPnC4+C5kXwYOV2pgMNbnTLvQmSesD1ShgFyUwh1eJ4BdvlulXMxR6sXovuEq04Z3hP0CRs
f0IKvbf8CZVcC0VTrjom7kPaP9YRL1qhbuRfeBFhOrzE+SM50q2S5EamOLKAgcpq8yi8unfja1sR
x4k0VnQ48VtYZAFbHmuJ/Z5Zc1viwVCIFg9+hKC3bTuJcGsAQ8MxlwmM/WhQJM2gZw6hgXI44tLa
AeL6TOrUDJqyJSU80fMjV0SJ0GufQcQRzXjWmqxocVxwQS4QjXc19+UQiD4S78JZKxYN+pmnxQRz
oH2/MKNdlke0NX6LWkESBNe+/uqtnMUB2ElnnGFUWD6EpEWs7250IeqUAzDRgr4VgyFsqgYUWG5w
7qvLd7NE2SBT9F6G6mh0wMtYyLw2sszTtyd6CBwTya3VoibiXiZhcNMAcbZpDd8uIpNSqLIcMAaq
LhsCx38P00srMdhx3vqjCxc4sePDhqn/0bbUWZgLNMrp477UiCrog9NeaeZ/Q64jl6+dMZzQEy3D
LJkzroYgEe+3gPuVhzLw0oloBN2nUEJnJB3/MUdX1XGMu8Hk/F/PgA2iGEfMShY+vUpKNvVOG7sv
NFCSrNzAkT+lGdvuKwD6MpsISj7lodwqj6Ia+z4oKjtGcN5G3H3HjlRpI22ia0LoB27I3qwwIM4H
S2v8STmhQsGUXz+Z6fZxTQoa79JvbQemvAZcYAD95RxmldEFSaF8/Z/6N887OIgCSOgGcJ+K84TP
Xerx8w4BCq5pFffOrqy4pM68JlKm9XlnxmfDeHa0ZLcbCab+GGg4oDilOTaLtwKKYkHfwjX3C5cN
plfQ8xZ4vE+WWzu/E+skkrKhchDZuwdj5f+0SAdEPE4hJdrQYlIl9JudEtUOpX+FgLpcMstGfJ7F
WbmXdyEZ/AuwKjv/MRHTHjjsztO2TmL+SD8lFdXxqtx1RK51f6ICfIG5DWcZqsVJHgUyRw8ZnkzT
Ev6NGdTYqosm3Rf6xy34w07+f93XjxGNNJgmo7Yllz18sw0Mm16hRLMQZgCTr8JqE4QYa/FjgN35
UJk3hbTk//GPcQCNTp7Kqarh/jxfr2zWuqwY9FQbQ9zAO38ipg/95IEBxB0uMfpBeWcQmZYnxODh
Swn8oOTosMK7UgSw4HisQ7xB5PKo1pLrI+Tu7V2+3S3W7ZyhNYslC5BH9qEgNXX8l126YSqdCtYU
Q8x4zP6ASX+qamYomLO0slW4Tqa9MQ82rGbzrlQOGfZiDDqOBiLwjT7uL2eUTHults4rbLKIOVEH
Y0ixlFKlLnJWDmCQwjU+mXOr1A0Hx1PRYqk8heyYQH97tTAUGnkTmsdieTSLvSdnLhp81AR6HkAR
Ll07iWw89p58PEiFXjvAoUIaTeFuiOflaNn7kCvhNKtXOHS0E3QBgp3/gMjJX2kiAiA3eClDItVy
flGFrc7Kqlvl+0tR61GTqArzBHCFSfUNOpmg+m6lkE6cbtblGFY65H/0LesIFJgIaTTgQw211zEt
AJM5Rvny4YAUtgaJSbu0OfBEVSJTh4l0njXNVE2kx9W2VyLkTw4TPoCquAzF1h+5MdbsGK05amij
IvqwVcv7k6R6XIB2Mrz/2Rs6BtvPLeqU9B9a62d9BFk7FLM2I7PDXhjxk6QG+Bx3NNb2kfCzcwy3
v4volmDKhDYHlkho8RLpYG4D5qecIVlNQ2zHTEQxjxk9oFDgiwo0uPCo3LCeOUhjyQdUZErClbN0
DQNlGZd9zKvE0hYy26XIKLHr6vjSi6yvYauVZmld8xD1Fs+Xz5GAqG6YMnGcIgQnkPV05su86+iW
mZ5GDHMYP1JWxPX7LxOIJll1/1cQS7yiBmLzg8DhbFmr1sKLkS8GHrk/8m8ujopu0frqyvFqz6no
RoRfaEUNkDHD+0zPWY/jaC7QggzvsNAwmuMsZux43meVetKcimTcNh1x3+svzq1Vxzz5J2akU7ng
TLSOIWEvRxGT99PEMHMOgjMKWezC3f559RhPjw4F8+sIKPvvgz2hL5aBQdXalyVYKVjP9hoELO/x
j09QHhYrMDj9TaDUg8KWLhIkZzdxZ58MGeBMHcLtDLXpKtlJFKq3sueZ27sVep2maMa9UTu+3tbO
lfbp19CrQvGUXfZ472Tr7yVomjj4p7zhiG5tA4k+2+YkOAg9lMaOF3TtWAzQDtqnlHI8jVc5rv2j
99fWPFWHfOt8sAo+oAEtN9GFjud0z/pFieHbrHC+OsJtwWsFOeIysOx+c+SbEpjQ4EV7ROCggr2v
NYCMoqpJM9C7RNp28hzSCBsGajmu0gYyqz/KGeNC774GM5QRgZfamZlWyBWcfA6w+fC7xDhx5LFU
+iRvwIU1DQPmFUYlG2/M3sk1AMYvO3aBE6sWDTcKcCKE5efBB7QJnGKHSjieAhPwnHL3tliVuYUn
d60HNDNh3IfKt54M8dwykc8rAZFjO/Bcu22sF+pzTj2BA14uWZmf9DzRfK6qr2L7Ag3RncVtCmsD
pOhNFWYuCBsucj0jigGOQciDn2sndCgxTdN5Bs44nv1vHj7eL6WGSTt1pio9RlHhZFGTS/dMeFE7
Bfe5Bsbvw1K/nB+g6oEKz0LdpgJog1BPVkKAMMr5WBmiiGXdVwz7BQZnp06nfcu34grfb4JjN5l3
Z8RAAIenC8XUejp22gBE+mYuQOqq2GO2oFvhxpc5Ke9Vdl2qmTRtT6kaa9a/E0BVuFW/wt1Gs7k7
Fff/J0wuKlSRUn3X8tqmZccY/6nIqGAv7b+7r2e6HpIz+XTS9DKhisWAiVDnp5RejJ273eoP4dZs
61el/g51xVAcn3+dNnGwLF4qPa4IVKpGp7CWkzidk812u+SM4eTp2XnGKZJ6Evls+XrI8FSqQbI1
sxOfe9new/+xPQb9h2d5iBpTtz2yMull6VKnwj4oMC9Chod/fm2bbwD7hsYhGT3CyZM0tt/k/Ups
XSJ9Iy0sslOZborJMIqms/aZdy93TSf1l9hbq9eDX5b42csMbxhsCUqvNaeFHVW7KFum6D64BhNS
qqeJO0ounPhyCE5wHqCjT1SQflJ7Dip2V0GDv8lxn4aHhLnBHrXG7CSXc9MxMqc/kUado5wqZM9w
v9k2ggz5DEqFF9hKAUbfFupzJD0mu/FEX2KjSZgQfJs+gVO/SKOrbF/f2xzYy4ELT3P6iQnFK9ap
r0/hdBUbcM3leMkizXPBmjiohgV05PrmEwZuGLsnd05P0tHNMOhhzAVoxMr64oyKucDcZgjoHgkC
RuuRsPkBPAJZWUbPEyEh/NG3y1cujYo7UKSqGBFRbtWdAj1mty2VyImyDgz7CuP2cHuatkE7dDrN
LAu+Bc5CzOdcsATTUjLdVw+uV5BdBvoENNCJroT0UKjoyUnqQgBvXzunXGDVGxUPcnGiCqDBCViz
F7U5C7xSUjgB9BaJ8rlNVhXexbidb1DEZD7LFQu+GXYBS2Rkcn7rNQNDPO6dePGtAPsPyl60cWcH
r9txWc10slz0KHwN5sBGkr13lDHZDrl50toWbw42QPIjbs93UuL1TUjbyvG1nIHHlGgTefsbdq2l
kVabwD40kAcU5C/rd6bDkzwGk0yLrVrwyw/f563XU7OUVrognslph/zwvt8O38ZummJp6rge0jY1
eZrnhrEySBtlv/+wX+Kq4PbuEV27OTVoGmgT5VUI0KuX80O6FQ58bG22FICDIHNqzjZjpwHyX3bE
z2ZW5bSBKTmKNWG1gVthbvIK/UDaCNFQQERONz1rJri7GBFNoklUHSpXJTj8Bm8LsGMmfREh8io4
kEcmHIDGNrLU82gJUDIEDTCSx43d1/n+X8UiICVaVPrK8hFtKP7vJqb6LZqfqtQUh89I7nEzLfu6
w1EqJWcMpCi6d5VJbbokh6ZVg3y5siOSfN8duPcvm4L5SQz0l7QNmdwZo9hZKlz7ll+bnFzpR5KN
J4TlAtwE4Xtn85JNYAdWnYZMCauQeJSlTui75ftNCezeJg9akwFodim8L2pI5RYk21EvHmCigA5n
UtoQKw1PlCXp806MIMYo6qLXvpIbrSauK5L4ecQ+p0L1p8KYzVK4l4NEBQjVjKE/aepuNxQuQx4a
w8ZdG6aD+FsrkM25dzgdNlqDddWW7AwXHTyi0Spq1w7IKaPPSSwHKIFqRUeEHwKzv0ZODd/3dvbz
ceniGHEICmJUOY6Kz6ACGVXMoNR0GOlJpbrdTJV64GBhgfOFn4xI7lJaAkfOuX47PQT38Oia2A0W
b3uroChOO7pcoO6xC5sIZrN0o1rLzkITjLUv5ygRgym8pGw5Ngbg2I1KzQ+LCeYR8utMWpWc6fiw
QiYFwsjHGQaz/w9ZWmSB7kqwmTo3jzbWXnZRcTxYyV42LGSOSW3zErwlWaZxQu/wL97Jnu0L+zEe
tkXgz6BWfLHP+4Eg6uOQn4d6nj0/kBRbvoqkhxexHMuW/cN+sr6DAmaK5Muq1wD4FmlbuwNJu3vK
D/179r/UY00GghY2w/nUQalZ79KcS2603mjLSSprmuLe5xKWqSb66W7HIkA1Vwxn0vzS+AL+kxNk
yeNEKTPoVwdHUEdKYE5r3NcswN131kH1cVA9FuXWJujc3ggQNHv/7Kfvicy1VKAnVNwbgDNqXUyG
UJqA924ufWXdXhd3rYBQq+eLcPhcH+cQsDptHbyV4q2lr6ThpEjld5KTOlqEQPOQQ0F4bFTZ5Whg
BhMT4nOGqp7SuzLLA3FDuQsBQDNnXpdF9IqOuAZVhiHBzcwS/OnkfydVIgQQ53/V92Mxh0t6kdWh
oUomoG+rv8YOyshDJXxQobMXAjfIqoa3PrAyuAE5LXM5uLtTe+MgwBBLa+WfDbhIXHqK9PLVOH6X
Deh5NvpQLY8Ou/n3FmilQ3odbMUHod2MUjiAlPHPW8z1jLRyFBWc9rt6yq9b4BZCouwERBUrgvj1
aFpZeYHSfkCmTMjpidc4aLuTTVL+setcsIGNaY1Z5WGLzxZw3EXqc6cvvVFzs2mteTS1udHrKIlc
UurMNeLeNMkR3GLnBzX2uPxINy9dxgR5H4LEcoDxP3UZotD0t3AmKU0uY19/KDtryPoHG8b0psj2
u5eTwQCZqEQ4yBJ1W962fgB1XbbQvmsEbI9+H8u3AAHVilvKYCzBn7VFmHo4slVfAWJpY0eoa0bB
JPlL4vtl5QQ03NClpv+k3SC+RFRTguI0k8WKQvTXVrYqAd/CDRldgTdH+jsEHIjA1qEbucZK2BgF
X4HBs2GksIhGCNNGRdRALeAFBgXEyi0+7Y1q1ym5VApbXCMvHiXtO2oq1P2QaTI7/2sHpJY1dtxT
FSN50MGNuY6S5LfnFmf4h8O+ynp106uqeSvtJUfakB1MFNA1RdfCgib5N0Uz3XUahd+os2K+Jv1M
wPvRMjTrFYl2H6LV4H6IgZpn9azCHAF5Y27VlEmToF+LYJqczOMf6HZGK47z/vn8x9IaNF9a5+Ty
nOVubX8pdk1R5c/SgVUsYD9maHqJAAU/DREYu4KqHS0ym3UvDQ8c6ujbHu3qRsQYV9ifgDyzJsHr
dN6mE0eB8RHVWZnP/cgPBtQ/rCtQ8qvhKgDTYSf9S1zh9YNKI+bVfeqIE40kxbZUvHxeD0jm9rmf
YqfJUMfmsFKJt1X97yUhYvSjkvIwoFotz/2qUGWqdLhIgqOHaRuyagKTsVzgbQJ1j/U4VE0M0/V9
q7Ag3x9T9JS8kKM0FDM0WN0lHxfrw3Cg8eRJPAc19Az2WCkyIsceoapAIKbuCVB31Rh+3yJuvXwm
X2433VtK+TgqQHtKuCQS1J9n+oktq9SoWGRveDJ6RZP5a9LhBh3f1UgSi+KVtTOIP+PFkAorqRoF
QnKkeDUx34TMmCDDWMC1iz6FlA+R3Adiq7NWwges+1jYLOr91SJiXLgcSaKBhfn0dNCOsmFS+Lzs
6k4y501WZntnlb+aUa9BUdA9vG/4Ak20xO8zlyFtrfAcwITF3xdIR00hRgkyZAyli0o1xr+PjmRm
u32Lt5w+ZTWLKMLL3lAcC2kK8nc3TpiYAyDmDalPtPdayV7f1almJQhzF1o1D3xcBs1dyHbpJQQj
rbZd5cgX8tRWAIZjXayhvD+/cn7JL/l0pth1BBEGBUMMWvlGgdR9LgVAHgtQcaFEJr69ryWB8iRe
qfmFKj26yHy3+97LZdCzu8R+tw/eetMlPBmlRP8HAqU/N+YEnmRNKNv1sxg769wZb+UxzmYpWMx1
0w2nTj20m6OReudojJwZngfmZOfjiKC0FreuUh63spRGNXOTF8Nr9SiIQ/tQF/Y7WGd1lUjtngV3
6RNEAAjnPZOTWBa7tp1UUGgnjapb8f7yPvmWaXczWYN4AZTlC7g8lqjcLZpzcJ6RGD875h04hWY6
M0Cy/x5G01B+phbn+kcXnD+F6bg5jtodAxygUCByldnRKXVJtDyGcrPR6Jg9yMiHWf5GPbkfgAzp
it15RceyrX2vvpTye8pPAuo2TP72c/IUd9HuebgfL4ZiQVEAqP+LSW2WgOvXLjadTTUP0vk36uOb
7E2AP92MAn1rSgQm+bUBhHoDoE85gih5WVXqonMHjyXKJb3rLmyZf5V5dwUxMLGdX4YPomD05XsK
1NT67Ws8iDpJMbAMiXjIH0cXSL7XO/myQBGJMCOAWrrpb8MoKJFc+tmII6ZqhlJMvjVDSTL1eSH7
wXSJmjeoedquCTE76bDLnTKRIKtQUNFjJvx1JAR3mKQyAXHorOYAzuYHxPCOEjnCyeP10M2NKp3R
r+LgeL3wI561ryA1kIixejSltylJ8piNnJLr2/DV6rAxorjFxMXhBWlXwYfKz1NL2EUQhq9Nq4Rz
vxUePx2rEPFDVW6ar/r2/VrbvNmPKPW1HgW7solc/fq9PQyhVKY3q8apUCYLzrk9zUgqIPRnjDH9
3iIViC6+5NG+lAwG6qPESVPAdU47fzT6JI+OJTCQokbRejWnKxZ+WEi35jahkxYpgsIRrZ3XYu+P
cl2tIV7lzC+WTYDGihgtl1BPA6PEN6ZytesPCOgjq9kIOYl/1kU0JFPTXmQVPclWPI60ZwRH2dcN
1qldwNblqGQ19zfHbsrlBomp7MWfC6cIr/kExYAL/nYSKLDCzh5LPDC3+yW75Er3du7m7wuVktcT
HJdncph8qGHmXmBeH0ObH3iRRw2A6/CPyAO6uvffKTwKBRuZOCWR3BLB/502jPZG3CFoLmZoZtk1
6sFxTk+2DJVBAq3vaNwbnIo+EACH+OV/kRfv8AGXbHX8Ai4t2kcWlH/08/QGBRkPyUaazH4IFqeh
wB0znuhoeSIn0lmdA5Y3MikscFPUi9qJhZ3cBiYHjIHUG6E8JgAIkpUebNjYtmQ15ME6ThpiwLnG
AI20UsCS06f4QQeU5qqpTIvlWJbhx6EhAAwqCroZBQw2VgF6OSzmupg1MLgRXgtve8MuDDZMr0SL
kl6CJX0g9gVcLQJhCKYZ2iqAgLmOB0pnXLWOq3qNyP+LMlAmYOj6Ffmj06W6QmRenzcA63PE3cSS
U12MBx2Jmd59oWgK3k5ZA8dU2UqxLNCb2vdJDeng4Iu+iPr5SRkkp2zm4DlI8jYPN95G6mhF5eRY
c453X2Oc060g1L97SzpQw+DmZ+54/zpcz9olcRRypwqGO2ZeYdli4tFQ+rqd3E9m+lJQVcvJ1tKb
Bp1rbVIL7fitSou3nwOpNab3sfDsCz+1CY0Kbf4332u5Cm0+OuBXh9C+6f6MelFQRC3sXTZ3y1pP
unL9VWnAMjPZFUkYrbgtTCuClBl6kU0Uf9Am6176yCJFnDBro49RoEpWPYwmHbJHNoIyjEftkOPp
L0L3eU23DAltKGRtYxHFJoogdN1ljSDrUI0/DrVQKliyAqTB0MOZO1O8Hr1E5J0sgWxW1rZ8KCFr
TPsyoX9mlxs1ne+IXRncW+rBl635Ug2mu3SMaKBj3cLqQZHZDtcOGtFuxSJ+hS0fVx9oopfMB9DB
3xuZI4x5iuSjEq1bX72HCuPRA2OgVKszzZOUdCMbkHNm1V7xp2m/YF28jQa9ic+BwXipTL7n+ajK
IG2vbM75UlYlZi7iTfBOrhJr/P9JCQmMLdRCxq32ftyo2cTjS3/2/HyoYuXQWTVg4tpHkrJu/hlk
8mqXNeqowIAmbQ+2PxixSYtKP13uEAYLm6cnCs6vOv9TXVOO7sBUX6QygEG1u6kF/K01S5mIA+as
3EvX2urQHcwESTAljJK01eY3rNbtMigngwptHl4qeIEUI2ZLUKz+rspTsQ3aniAt7HrGKCzAXoTd
D5tu9VGS7IODisd6WMoR9YEWRV8bPj+e/5P2spIfJ7Ke0wrqIECR2a/LNpyamCx25mz2LUiooRQ2
8FrQrBhPRAVaDSgJQft+Eyecq5WwVVTfaHpK0+K+Lq9sesl7oWh6A6RJmyWrfoKggzS3FvLXcauX
GGyDRSRSRtCRwxt9Pk0UpRdBQoBHJvNavkCkzGBc7nPo46cDRYkMxUZjDfu21TtLxUoQgcKLZ46h
UJxOZjErdVHJ9xiSNUgTD30ZRi4IwYt3lzL+Q6CzowOSN1jL7vesUxYygPHH9an/jfBk+aZuyxV1
C7E/o7QqbpkVUeyHlMvzwkGEkWbxtxuPwPopZaYSTCUI/FSqPmg89i0Ui7oFZPbm9h2f9WhuyY5o
9frQf+UPoJ6+FuDBu9qf9Hvimmdrv+mstvmpKhneWBrf6uQ1CmPJBjinEWZZpLsargmZP+DfAgzu
TScl9Po5kV5oISaQCT8EEqpBFdXjyqFg8Q6WCwyiXa5pLPThbnSc5RX2R+m42/MApAGSy53EeBDu
oImbTVfO8J0thctl3dY75RnHjB9qDPcSa8Y6g43aVMo7tK0WPr+4EA0bRD1nfOqeDPSZ9LmZ1tyn
ZW8dm+vnmDxwfcEQCv3F0orFmTzQWoLeIPytWLC5HEcEqujA+jLKC6OpnwxG3Xz5EINsRrqydyWZ
JibZ6EhDWj3WdojmR0SK9XNYP5YmgFv8s7Wh+L8+7xsFGLAf6ZujL9u1rpTitRdSVxOtfq8lNNaw
GCQEBTNTWmZerL2FF/rA8hwCoohL6Of8alQPAtCJkugEPDA4CED6KdVYRWM/6iTcKlvhpg18sQSV
ifbgmbOu9RYp0Fsv+pY1Hf6NbhDQ7luHvUZw44BzJp2S+ltlttA5FyFnC1qNtJFSbxRjvXFBl4r6
RNCLziDXEUhQECKANrrGTmZuDvz5g3EDeplju6sVQJ3yjENVZgNh2l38BmqYHBI57/cBwinODaLE
IQODwQlXQGLsDVJWRRstToJTj51ImTz5OkXh5GT6J2qK4eorc25OncD77kZ97hG34V4DiGZHFapH
HVTppaqQi+nV1qUE1NxZPs+QnefucLtqKdXS1i8i6431oxHFM2Xxd/HzVNbOXpqW0HY0qkQFUlP2
veebgTx2gl82CkFJjJlD3VZWqyHDp4jRj78TCf/aPyF91LUJh6jvjEzcc/KmthIlf8PZrh3QmT8i
YQA3IWNq2p6w09BrzQm4v1BStJp5SwfYG2v9EEcd34Z6pqfqZ4+xBbbjwddVFFpft4+MXlMOFrrL
ees4ZBlAhCMjw1wZIeFi8eajJODEc1cSdzF0lT+4uG0MYgPrFx/ghdIT+/XUl1//ODnT3K6KBJVi
JidsDxpsHSCNsouX1ym7uk1TP7wMfuPH4dID4Cfu3pcOOXqtL3fKJHg8vzip/Y2lGqcsdAiXliX4
GutWz9N2IW24QJmvBBFiQcKC/o/ncCqOfHoJI1BgTn/NVd6Ype0ja7m3eLpynXgYHEDqDnIu+0YK
GfwXeaauGgZ4eJZvGkXLVuT6o1j0flYmrL/CYaZynQxTODHwX1BecBathHa7bgp1sJ/DVK0BfMhd
CDNq5yFhlr863BzfOKl0DswnBFM9rFZQSG/04lhlpCvqkKgdddwx16g39bAH8l/0AJJWtKeAjg6B
pOpodLpMA6Z6ouM+o8lHmOhSMpPUqpfEfZGW+B9VVPsus4sNfCP8WrHJMGuyjaT9+ed32WWnGlkI
M5TtXRbRi36n875SzQ0Mba/Di+5YA18unEAMFBHAr0FkqidgJy4w7wF+dzalXhZsQSeHHyMgH8HY
Y0q+kN3rD7qq01gMrLADqK18wUsv8V4esKu/Q1VH3iIR7qxy6ysqo2WU1b+0F/mXdfyqOnhzdgse
VY8TN8jCH1Sr5+EZiip1E89aLw70IHollBB9es20uNxXuiYyxZAgz2BsoXXTAXjiOAYm6/VdPGju
8JPp3ctQMd4bYB1RG9L4c2JbSdzgfOW4C662DK/Nd0sEc4yt6ICrt4DEpBPezY7OL4PD+gBfbybb
D2xwho5spQhgGGE9rcB88A8TuPBqz4KOGtjcGygdEL3CRFGd/idY5XQIiRxgAqf/qiUrKSxdrAY0
IvXilG3G3x5nzvxaqRTr66Vj8nTO1l5jOlXc7ccZvK5TCtfF1AoWnZuJ2HC1hQdUAsJadvvCc+AP
RfFUL0lvqfVh1lTyZRyUu56oXfyRLcAOJ6HLODxN3+3+v+JwpOdu4TiF5EWNjd3IEoSbM0TYoJZP
9WPTVbFtb8aLyiT0hq6680akqEHXI2nSAS78ew/ZJuOH0TyIFO/UezhQw6kz/fVPBkcN6a06uQ7I
/74tTq2TyDUEaHeSgwuG6ENy58Br8QdxLomaeDqJPaf8k4zvLSqMWbjS3UABegyXYINpkfD2ikyn
omdXnpPnklqhyZP0LX+ChwOMw+NcQAgAj40n3YWSYfWBIgUBkPIY2i5WgMXSbmL9uW5LAjqaJ4DZ
TuFt5FlFooRnc1z9OiA/ppyd7NPIYT3VjKo5/hmc0bIon9Q5SdEn+ktbEd25lmhC0bdCmcBQBTKx
Yz7MSK7K6xaUJKrbTeUVrH7vsnqIerxZ3ncjfUm5kZ7ng/skB1G35A12rV/w0Tu2hRpI4Ochlap7
gch3ynMVv8kEGxRHEM+y+Cq3xvkJfkMfOR7vp4aqvsLskLY6jWLg1+4GCDCjHFnxjVnW+O+/K5iA
8+HFSAmCqHChivCSCMmNQrjR+9x/78BQSTJNheUOjxU/RoY7c3YJJm6QR7GGCKxUfg0HKessgb1P
lrOVHNXvrOSm5zPUDdhY2dVbukj7EgDOsQhu2MOfzoRSljEOkbwkp1CWV5RV3ctEKcdx66hJ9P9p
enD3dSYTFVQgwvF9jdJRREtGwEV20Hozv0gIaJEFchMmDB7liktkFVibUB8+rhxUxDstte0oMxOF
I/M3SiIUPhQJOAf6gme6mGT6qgZMOH+RdjOvj3Xrj9N9BH11WKAfw5NAquHl06XGbiM8ZWcOf1/q
0u0qgqYanwhJkjmAjDvwJkV2jmie/edYXEwuexPEXbIh0LwMyQZ2wCL/teePfas+FwjUXbmYghrX
85Dd0wC42tXOmpAtXsj4n1dA7vjO8g==
`protect end_protected

