

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
CWO2bSovBvQ2ByFi3vbGk64Kz9+OlU+ol4ZycfRhtc5mzW4spj2ZUNH57Z6TD/HWbssYOjRT+UqT
ip6xHZc7sA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
nB5KuhofnITTIpXOtfG8vxQ8BtQATMQkEP+DmIE09Znrcw3yJd8Ym9iSaEwPi49QFbQ4UCNnUF1p
Ci6v7CITkdmn7C29rKsxyl5fQwQ4Yg2Y9J8sH3IMncLyMWd/eC2FXu2c+nIyMZ2PxTUPVrUjVKNp
s7scT7Me3sAj5vk8vEk=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
MNNArzGZfZxohM+fQiY689sNLR2SVnrB6IH+/5sMb7hSfawQFJxphTI8Kro2JGGDqNxumEJLUYrG
7mZGSE03rCaVpdhD6Rm70zB4CVRXmxwbIpEK83cCm08nMbZ8k4fK0avkhJQjAW3CnUztsuq7IA0K
kdwznIXZSyXH6lPiqjIN2Skr4/LMpA0PrKFOFlQVuPkT5ZvNvxenTGhCq9p/EpzKYQA/Q64z1Pcv
8PTscPeWEIpmqBcuycpxO0kwVqiQNRqP/TotOuVFkjYLePFpvLupJo2vDdC4y5SiD3RT9wZvaSz2
Bb8UYdK03OxRsiXtjWytUX0MRrf53QlD+4mRvw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
JO39BJFIHsw8fi/kSg8TBE7CDuzx+VxY3tt2e34SSpwe1+CidGWrS2YpQSFw2o2o0JVA8lhp2pEl
VW+YDwewZ52gevHf/k4qIWqrG228k15Q2kpUAiHbcd1YG0RCacsRIqlWdSiw7wc/2b5Il9la2dZd
yyMNm5GMzs0PBGaInn8=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
DxfcLsCbVgOrlbX9FvTGJxwVAV0OB3tR+6ByNYT/Wivn1M9TCrq2dM/5FWlDqpdxHIYJfhQjjzlJ
F9cbuhfluBOxtIUuGdHg2uX5LqlRjgmnPZ6fbuzAGkBvSUoSqWJpXOKWx36bmV4iGY/0e23H2hgI
ZyfwOhBcKKufNk+Nq7xnSV7GWSBSiZWYhL47CEdCY+E8EYmyeXyXT8RcA9zqsfKsEZqdz1rU0vql
DdxwHxaE1OVS6MuW2h6qgK3l9I9LyDohZgyoP4VpBk/e9sTSLxcSmGiXwe6zlvuSw8MrBIn34Ezs
uAteiO0K8WEa+5P+7J56z0wy1dst9IfRzCpYUA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 45648)
`protect data_block
FQjvNcyL+KY8EzFxEhFvQgJCTJgk4U34C67RxOsrpJcdum4ewshYiukRRXYuYVWafSoLLp4vd2xi
Al6GjcW7l1qG1kiLv8yt4nGKx31XTU4VG6u04tXJFKhFvM/9+1YrJPyDzCCb1mTWfXky6ra+cWuo
4w2fv4HSuWMp92r3CrFzx3GIwMPx+f7Cq9EdHso/9lbqKTsAsqwXI/66EMiIPDCF9jNkKRqaiCbh
KQIlPoSj9umDtBiBORr8FJRkaVx5Tmf+JLAhW9G5ysIkAaPfM0LkVpBPujOMu+tODV3V7g4264ih
q7Gge3+KFRQvTGLh3A4WfaGTCagL4rS3qlveN/ZviHvHKE6QiFRDhR0jG3iu1xUFQBEzJj86wecn
m+7bSQ35FvgNjNG3e5M40+sDzUvAOa7Ex25Dt1T3IDtre6U1j3NRbGFFTYu/deXtR7aJE1Ei81jQ
fCM860DEJK6mIePNvr/IKSQC1V5dRxTqq9EgIa4cCDl9p4QIACKjmAKi6Fz6I6fHu6egUQyMM3rZ
6jUN9vi6rhwZlKFyYfFsZa/z8NVNpvT6zBlXCpjcNNUFaLRMaSHhmzPsoIKwu9OkAk0ZS5aNr9XM
X4HDpfLy/l0CfS2rf2Fwhaz8LXV3VUlPpQU4gCsa75zeQ0dJjKuwqfVLR0IvSA96yTcXl4VYg7vT
cYuE32N/TmmH9/4Dr6nJkT9pWhdBpXKW5B2rfoAiD7QtZo8iFohmoR3DdNkMQD3ylhKTJl9qhX9T
QMO2A/FLnX+YuraYcadgPwlhtirbdp6PCFO45uFcu1LAn0ztRMsEb7dr+yc0F8qPbGza2ob1boxO
6uAUqzgXrHyedYEFmT9jrXKO0KJfYk/jp1eAmy7CRnQYdh+XhpVONEfaCBc04IcD1ASIWL2u4QWK
pYZzzz4RA1xiQul6ZRWBPp9vfls9vPBmsEX2jxPz2QkcxJqmunZiitcHCapFcN/mlcCacD4u76Xw
YOBVMANvPIe/56Bw1Gj4QkKDh4B+zBXlWwRAHpZXjqCSndkE2qMsrFKR1jvq96l9ZcZoRqmJPpfs
sA+a9P02H+IEQ8pppvPCAAwyAmKLbrv5WwwCcrR3kpsEVKXgshrFGVns3gk3unB6EQLA1CdDg4xC
IIDfGI09Do+u7hknOpOCxJSM3w4XvzgIPmqRgooxpIiZlWsboU2pJ5kWGijiLjZ+e87KuVXvJWoU
8XO736Q3XzdHUbc2LEOdJ7/l2datOHMuLE+OrjYUXOKrXKPCbnx1+bB/2o3N6VTZXAa+rgVC3Nys
d3yBrwLOUW/UMhAA0XHJbPSWQQRSjseoDBGuFm84C9TS5qyAGQDJwLVT0HA56X4pBF/TzqGnivZL
zNn1hX5J5f2MThmMjaqKeX/CJndsWY9U3M8ajufONhsnUEVwe8fhUR5x99ptxQYxEirxvqgsYx3q
kA0OBIAKaGV+bh5lvxRem1PQkgUQqeSrWWbGuTjIuPiourmIBVjYa5b7Ur4Q2vUQgud37U9SRY3H
W8/xqg6UeDJ8VNWBUshw2zXaAIf2HlKbRS9h6mc+ThW/nmKWW2GNNuZDg142mKue4u8YTAn3NzBl
lrwccX2DFfFk+rI+8K3DpRAims8LqbmPtIzXgUhUHP0BXrgoLmP+F1Bv2UKjbX7ynANMmLdVYdeO
fzy0S4VvvCy+fy7C+LCtbnB12Y/hkXu3WFZl94pUdc/WEccK6Bi5k0+CjnGNdSIpdwu8nATRBbBz
ZSN2CG0HHGaUDiFihfZkZnRUh9luq0hF9x3FnwwryYn3oo6NxqE1ilC9nj9qDzF+uLO30iXK/c6X
dByi6jTE9NvMisbMSh5ff+AWeMrQt3TBNVAFcpsy3PIUW+N30JmXUx/a0yROJ1ZlwcxkzmeGmO3d
yp38BYSRJNZdYrNTZI6XPdbvzLAIOgnmUPB6zriEFHakC4+sAs4Cu+Wx621k5GuYy9PA0il+i6Yk
LSLa1gq3Szi4ZuT5VV1dfHqnyyyWlSM5A/8oWIeR75Se53mD3kvqpZWKYJCvojFP25j/wC5FaJ67
iBOkyGA9qiWcQrmoUtAcnBce5vFFmtD6igJ06l5f1igMVcEU84wU1kKeRhuBRPq06LdVRCbB615f
pbcYylN1MQEksziGoF9JABS16MnAc1fbVvfF7m5khP30FKtA/07X8SlDenYWdEywmKJU9Q5E2xuR
EX1m+nI1PyUDl5mqOJvq2outd012kiKSShqzAIZoD+EqsC2ptGrC5CPo8Ygvu3C5ypKE45kKERys
/Gw0lbGVi+FYqXNw2qGtMGD6kJidlnfq3OAXF+soDSI3F9UfXdaPXQM/6QQzbW4+wGbU0yGmM7ms
QzJj1LVYN8AiHetXNk1+mUn2Hul+BHXku7ijJeyvQfoEqNrSatlKTfc4qUhnq6O2oixEEwlTw6BN
IxWwoJZ7yR/Lz+QaoSWyFk9GMXGtC0hi0GQJqpWwN64dUoi+PJA85OOplVTX77V07Bs8iHW5xAeL
k6w8zaqiMXlpfLNKakvXpWh+w1GRD8CEkPLlV07G8sZa7K5725uvaa46MG0IJXKg5oow/Fw2hDWF
jir2w1fXtuMOV0LRqMiypreaddXH5gXDGegWy3uAKFbHG8VE3yzvAE+ThhQBJwtjgUwnS1RzPiIP
DZl7P94N6fLcHKKxBOXXIRUesEBcXDoOGLVbSaTC8GhYEddyO/Ij9zdsy1Ddq/BPnC7S11AUQcpV
Fw3e159oq9Dpm95VzOkbuQPs4+aUf0XxUobS+K7D60qZMRv1uyLrZZXuPrO/jQQcP/Aly+WPKCtH
94lVraGSkf3peHmzwX2axAPniCL8xuCs1UhkSrAiqsWeL3jOWrzmD4ZmqoDpfIFoZwmNG2CUhMYA
K1Cwx3rKB4JbXRhQzePgzaya5U/XsGkrZG2Dp9jQfn7N4HkhwgGt3eWuTDEdBL4BDYWM2akZ+A8b
0uj8jM6EV/v5dMXiIOCKk/p/RLZ/rUR/HwmBiPz/GEMaMbdogCMAS8wKV/2trckI+H+Wo/h7Q0wO
1n6a6iesJn8D5Wk08TKhB1cs0oKTDXu458j/vcZ13YZq5JOdXJ+C/XVgXyoCcnNO4SAjdQiSjx8t
ANeyJIxocpJN0lsepHz8B19aoMQTqB37JVNrbZN9SzyxZhbID8fbHgciC4wSMHJ7kAL2xYxGKGRb
eoM4AsMuqmCwpgk4sGfZAKBhKJwrgDCIAYzDr2TxSGhaNSmxXtSGhxqMnuT4iCUDKZg+EbdfjvUw
jZgXENEy2+2mImbcJlBxi6TCL5+7vVWLFKXqW209oFZA3Mkx6vk61+zzlr2TZCamHgMg+s4NBFVE
zLx35ODPK8v9i2Nd+kMzQBVQBnrQHdPQHLWlW9dcmoVgb2z1UD7ATBhXqYL5E1g5dp+V0J7es6pA
LEGbcrjQhvKwqp+QpYXDUX0MnefxnV17BwNPQN706jnmcEHLKefx4yDGzKEArlIGHeIIu2mdmElF
BbLLaiyWisvj+nH2nddG7PNE1khsinrWjimcbpW+xfXcNMfhoOI3HPrkMWP8n5Sy25n4KWXBJ9rZ
saK8JgPONIbiPAIZ/XQRoijvDi9QhrHSE0G6PO+fZ8BUJgLnbJt7yU/Z1z+JUVqDqY8mgxvQyMjV
jbwpvcPmSlY3s/l9O4S+zlJg8O3EsXrmsvuUNpbE1ciqaA3/OFvDsVXXA5E5aV5F7s2g+qkUpFJB
3ViileW45Ztmn4oyq23W35D9vtmnJ0SAiYmgFyIXTxZZnoQ1dYhpd0Z6Noi/xH6urYMzWUGHMJq9
9NTE8iyqT59rjiKHpT0AjP/yDxYDFodjw4GVr7AEflHlVx7ge3iVQKLfi9/k8wLRbiYTbDixlDv/
eVr6VtUbuHcHyhUDKjxaU+FbrwoiaoAeiYoXFs4tH+YFX1iN0GE1zbcs+OrpPjp4di4+Oc64Mjmm
1eanJpP3fY9J/PXm8suFGn2fFbJJMTI0l4T7SKF6vLS173X6Gsew9xbOHd4tUdFpjS+RxCXb3ddH
efBjk8IEh+fpZ8V20KJpzZOUv4ta+Ke4EImyGenoaKY/yJHgzv8z9U33jxFYQdoUlL0S229LQZJD
aa5PcyYuVAfGg1bq9vI9gQbvyK+HHWN5WJxUG9Pzp0+hxxCo/FOYCfEQGvEnbMecuIbgwxOs2vOQ
OczCH1GMCc0YJuK5bQlRx3cLpAjyM9djvH7TdptmZjHnyFZoR0nXturCSKwjzSg6mEeZ/Wj1Z507
hg9/c8pCRmonWjwdMObZu2YZ7B+Ri+Dnfl9ZhZGJDD5JEyX7h5vXMarIz46d06wg3GLKwf/lPba2
h0+xvdHRKdfn2tRWnMMBpAvlOBrY/vstdeyl6bTYO/5j32zsjtP7tvV0ILWLgRqqstFoXVv3VVrE
arwt5Kr+Vzg9SAjpUuTjAl7ohXp1pCIyDdro3JZ2Xb3OmG1UcnKoIyTizM2tjagnOY860hVXwZj6
5zddNnMFKe6I6S6WCZs3EO/9VO51z0dSXzygA5dLJN4527ZWs9Gc2HpWaRDxv5pJZ3QpfMyITMi2
O5dENZVEk2IJPRHMDYw+eMVSCb5+HcsEgyVHJ9uWsbOv+Rs/sUpPtrEpKRCQHPSLfxmAG5TyqM2A
lZ9U1J+unfe/0mgYL3L0FLxWY2bTI7cUMMR44VF8oxYTRUoOMYIqnVgoAQ9mINsidl56Kr4kh2+T
vc9GS1ZWKjO2dBvxOx1r5mNQVK20nWaHOjzfgQLAK5qjfl+MViA/Cb9XaZgPnRKaN2A4ggkjdrN1
oe5Z1YYcpr8seO6obSfPZjOnooTHqOfcrsOuqimcpoHU/vedGzj1hEIh++N9QJCbGEfuOfQ8Lebh
8XnyZE9zFMUeMklBGqeeLgeTfQ3zOWU043KjEV+dihVAqrnQKLd1ddo3rXUWTbtdiUVL57Wn+P8L
KObmONAJywrM+/XeM10FeeYZoMsIrZO6jhpd+Py53tzVmG8pUeuBMGb1ch3bywPbSVzACGzxycap
9Gw/2Ri8yGmJvoOpirppDFCOtDDj5CuXgwO2zYUT6hCb3r/T90MzXw7xCZoQKezO2OF4JiDephdt
16TK/w4G3QldJl+w8dJPWtv4X1JDmkDhfPGyFBxWGpPIjDFbFxge0XQyyAVbowtT6uLxeGnhROBU
yCnUEXcbagdiG7LsbZrtjhmuN/IpfoNkfxBC9GJBIeja6m5UpyrGCaUkbefp5F+jZCEJHaeo0deu
dg1/MjZoNog/+418/MqzYwOtay3xGm45lcRyitZr16rbxV+WQpemvJFqFh5A9lp+q16aw3/blJdg
aszWsevDzS8eyGsd5LqUO47wnFdlpoQuz//ZOF/oRhyglH+wSGbn1KMGC+FYVwMW4i2nHi68xz2S
V5MCG7Ocja294kZ+aIW/ueV98P0SLTudo0UeUjW3gCaW5hlNCqaTCbjVQD9OypHg8Ebu2Id+Np0k
MzMm3N7FRxAbzmc879EwebaNkBp+WGBvzQ8PRNiFg2+zAbm0hD6lZdIoG0TEo5EjhmvN3Vm06mbS
RIXxftMzaf2IFbb8DC5FWfAf9r+zcajPsX/htjvPD/+0jwuSg6zVD6k2dgCER4ttHkSqnI/HPZVj
O6PtRxuvIa4tkAd3tpI7/3P4JIgdtaG5BbuUV4GzfXFfA+qvTYR2b/+nTUFY2JyqVMwOMNaHxBbZ
5wShmIHTxHmpv8uEKTh9c4BD8+XP18BMnV9bd8XZFYmRueokDM+6E3q2fzYwIGRYIKP3JR27XZjg
HQaMnpCgE9LR7wtM0TZNfdX3dkzvhpjyvw7SUZY2Fcru3uCldSR9k6B1j3RlClYzC8AeEOZyy2fn
8qGLvN1McUdiMsHEIa7Ve5OGGDX3hrpnQUoh7pXjDvYBmQafZN31mZH7LLXNAG01A8IbcxirxJe7
Gw9saLt3tdwV3SinIQDg5mHIwuc/ayRr8iS8/CYJi5nyC00pQpnulAVCW2I/V+WkC9TXon1VwcN4
hE8hfW45Q30NICEpT208ej/WkvVqwBKBVYMyKZzozGSvkrsvIGFOLXRAImRNPx1YxgqZ54gNmZNL
HGY0TUzv8MEQjk5X4Y6v395Jjgzj/XLXnNYyQDShoqy5NBUWryT+ZmV4E7IXTCDL7JIPKdvpUh1b
JOPM3S4ghhnq+XW4q6hPT/jkQn0ePE5Q0LwLvFKA4y5TtDSrARcyGYkcgd5b0Ak5e1YkomaRakqK
AL5Kq3Kv02g4HIyVBDXmLJ6uynUeZhG3Sz4U1o+d4lJZnwz64AEBqcckkhGnC0FAQos2J/yio8B5
POE9qfINcgQShHEgtVggkZF8T35JYzru51anEKtNp7zLWyiGjL8A1IA/lhAsUqjilAf9z2/x8NwL
e7OQG9uCbjmPd6S9fH7ODK1GqURSIN1jegwvZzKZ2mSyI3tAxyoJIvRERfvFwzt+X3xV9M4IekOL
9rMaurIWKmWSmFlkzgJgiDNkTgnCkfIH8hru9G6OU97tAGFwfnBuLZtqXmcD8xT+5pxRWbFJ6T1n
XDe6AjyfiF7yWjatSAwmlBcvRb7ecxa5J2vS1ltFaH4AY2S68OkfBw1pxPd1Of/MJwWt/Du8viVV
cdIqNCRHj7pes2hIXMSHXrEyQ0YPKU+6LZIAACeESk782GuH7tAG0UBEou44R3y43/o5avFTICaM
rGp/57HFqHPaIX+QVxNWuFFSD5ysOU9+7Dl0UFgT4P6LTCHnm7+FVBF7ficAemHVIkl8Rl9dkhRC
SYc5uj3EYcOTEiM0IUODiiktRkHeS+xXZq8jGbaFHsoz60oouGBSVQSmmzxCoSC0pvEMQVJbSRKf
TFydeQ9XxcySTQSes9EuWtiVrJWVNqt63+lZNrFb9tDZEiGqt5wpQf/fyhOI77KvZoqWLpv6CA5c
yveTPosRpJiyT2B5tFkNxMMzKZTjztCBBfv8r1d1YYlfy4iGUWgfxUamaqjlbV6iqMnDxdZbUEqG
FKX6NyqzKadrBN/Sr1SLED/9PzYOVrxwfKpiXF0Noh+Z2cuzuxHRn7PZOI4Jmpc/DaFVcC2SKOW+
8RTOKkrWFhOrRldky7Zm2/TcDSMHGJ3tx0Sxlk4HAISHGa4KL62BC9wTeSZe+z4yVF0nq2HurIVc
KS8dEyDy6u8J7TjayNYuPAuonfj+IOGJKgk9m0H9TU8UGDxumfvbUwuY1rjGaQnz+4o9jDdS8iVY
txaSqRe/JK0yz/XW2Z5o2pyNfBrRGTy00TxRxbQOv1QtLyZM2y/pSadr8OEFI3FEDr9E1Rd+EepC
5xJkhGWsLZXb1BAAIrJM0hy2oAhZmSnMWMXjYvommn5Spt/dBX83gBld/yc2Jzpmqo8QXmsxqts8
b5UciBgYvjMuA1uoUOBnpFXjxDaiJ/EZ+PB8hfiTxUJHj+W4wHwqjBHi9NIaM++5wajpUT9X59X/
5pD1aKbXoYVqi4RJBFCgOO4LgSYD2ZjHSc72p7oRiHqsV0+xIjuWCkU696G1C1d9WetuibvfOjkQ
5e/hbUBlCuSgeDDsje0Zs+ZQhE7+MfaLah3n8oiqW1+Er59uoLPY0TU/b6c5Rlu5eP6GtW/0dY9f
dtAroolywhUXqNMBMusk8n5sXJvzOepaCJ+oXWRGUOi+QYT8blbiBaBbNBKhlKCYjqveeMGRkP25
Yl6hRY1ILFKusUZfsD35LeUmeW0K+0IlcyYLKfdZqwggHgGnJTkuHplcwRWMshZxjpmrtLWAGvIh
8kJq5AwhpJZzqZoCwsUvRR6ePp0uA1eWf7AvJaOsxU07x3seWwsJQ/zC6+l2hbV5d6a8TCkt2QF1
YwBNgygZZh2UNVcqHIRNeL0Jab0YXm4rFSZDm5XUUkSGWvFXIA/yx1h+RYhgf27mJpVm9cdQzkuP
rUOqQcKI298ZGwvnX2Q6BEIvz6Ux6ccnl3tlYBVBIYvPfnWUsfLpj0cDG04an+4EfsEor8OvF7fk
k1RuCsU7XCcd5nBsOiCFftkGUehYnFIchOF11XYQI/NAA8p9S3qu+WwYsea4cu6xyiYPhOrxTgzv
bla83i07Y2KLIaj8WBfVUNPi9HVGKdv8T6RfOBeDqros8+GngMeHbNnHEf9Zt0VjXb6Q3wG1Rxem
QbbfbCEeXZKhBNKDteUc21tTYF9FDMq4Ow0FyEOkT35gWR/4H6J3kDhzYyhG5uBOyVsV7V/uVAzG
Bv5tH5THJwsoG/K8KZ1FuvekJ5+S8j0pRt+0BQW/KaNvQ1lmNS1utW4mxkct5Asl/ohGVqB0q3df
EOyNzJ4N0nfUx1odWreFpAvvK2DRMCbwuW9zQElTsomNBUu/WhsDzP7ywZfNuZAo0oirvlOyQ3OB
MRAl5XXdszXmO29hhV88GorvZuGZqIg00a5f+7lCUyoDvzJ3qu6xI7iwO86XtZeE3+qBbmAT/yLd
XnIb6EJzDqvr1Q47GkUPXO7mCwSxujVNLLFTop6LX0Bf9/w+/2v3LmStq0fSmnolOe1pGBaIXRZU
cLkM994b28RGbM6W8GNsA+7Vb8pC81jL09YDyYKUYfmDuDotU6/KbMrHDsk0eiFknO875CLyY11e
eGz3FuMT2/Ean/lrythvYXCy00LVcdMN55l2O5YH40sWJD+qkn0bbi/uBEPnl+sfKIXE29WaV2mw
DE3HhLFxcKbz9d/4ijHr6DttMjy4I8MZyLWUenvUxU7YV5aSkuPVJtZpRIrSg1WYlp3V+pyFiPeD
scVPsMNoPfUnaZ+0KAp2xBv50DnxH4jQsurOj7s5GPNaoqglF1+4rE4xwWREM7O8pE8NcbWKmo1o
KfkIN3EqY0LAHwDJNjCgVgWpZsE6v1/Amqo2kOWuWurqlr3EoGgwXSWBasT0Jr7ugFxZYHHP24SY
THblRRX7nwvx8b2IKUb2mLt98s/0DnrGU7oh2Gd4yd8UV3HxuFoXuWJoalo/SGUkdZCZ3LU6u4Ih
QrLcPU9CVbBjIHDgnLI+TZCT4GmqyhPjxmD8aw6DZ6CsQ86ju0VNnDSgKI094SDGXCfCMdQFl1aH
bSE3YemciUhigD5YYqSLH9TlZFlzVQbiJcvMRKvaEtPOHV+cm97DOHPNQJ6sJjWyOL9IMv+dJ9dG
v38KKD+HjFuqAR4UgnHLjMZGVUuZlTHuNlUmiwn7OqoA/0A3AS+i97CPU7sITN+7ahmGGhglYVDx
CXhifNuC/48lXRhh0MyKauhKJahe5nmwqFZZmzycDaZ28JV4FC7NBQQYnQThA6iY1t+g508jnWPt
8Yu8CRLvHW7hLhE2edLJ8RVhWZgwOrPQwjICqXMhhTxK6b9cDl+v1fkL9iRE+DFgWDqZaU5wekFT
9nXIF9xuhjM5pEYqUdK1RqJExRxwjQlOcNMWejf4pPPS5po3WyCEcwjfFCD4dqvju5oPBGvnvx1D
76vaVQlfOKdHpwY3Be9oWCZitcL6ypGP7j9U355gf8l0cgrC1fg1r5qWYgQQKRfl0K8ITkvNdj1B
/8vsmXfGohDnVkqGub3l84RFGg4GYEaTkgxeeqlKGtaVXNh/zpQE0jQFerUVrMMNluFUBS3gmR63
gLsIy7J+8Uw6gfLMiw/emKT7Rl+LakvSX6s8UYZkk2mDvHZ1yIT+tQozkvP7/W0vCfK80apSJAXZ
ErCvMzsQtFA8JxExPCyTsJSgw5Au4QU+CC1puJQhH1knUQ6wl85ktSEsjvcSX59IpNa/PoYt0OoR
4do5CZGlruglzkTMI83jAj1af+KIEwKXJGr9gX9JKbazUt2k05A2FfEfKkFPv37vu2sOVHAFRXiD
/wJ0j3c627yCJQdNbtZmxZZiSrcpeC33ofgd8rkkqnAS8XUpq235xRQoz6DCzaM+SHB6bfgM7QuY
ON2ElI5eQUI5IM2ZCnzCcTDzBSEsJk6bpw4cDF536zVI0G9NtNesVznBst+vXyhmn2kn+v2nwf0l
Lv1G5nMOk10KUgJzvOK6zP8FzB2Ud+/G8T4xSiUYwxjTlpCzUkfToIbmVl5Vm0MUIQD+x8gcTdJ6
b3k7vSb5EHTo16yAp3vFhUN+iYgS1e7qYapCX/pScLZmDVkHLItAo9tL1JXJMYoonJ3HShNC0w9M
MW22ZA4J93e98kkkeEbLAVdFUMHYUBJQmzQM+HAX9uHpSPpfq8xftVkrnS47LlCDZMnfAN6O6pTb
I2CuMaTQLauy5GO4+QdANgW3A5CgyLg4Cg/Z5v3GdhshZBW+62roATOY/Di/F4TOq0RUbT//CefY
pYjAjYcUcHTtF2RwQbhUQruMtz/eFgwgIwYvdP3ENRZwtZDPcDxsI0fptET6F5hLu+dZXcefuCIa
WrVPRUxR+4d6xzz9MaG7BfO8720BGwQQCsNML69y8P1y2NC3By562giPs+ALgs0CdW6x/UR+USDp
fEyyjpyOMSKv0+Ddu8HnB7bCHx/P9Lfhwk9BvgxDwYbINjQHt6/3y7jeYewpDWGCzDnkLB7or277
SyluR4Psn83YDO1/dIa8QS4C9Y0AtHiCscyjGzbDbzj/4DwqwuieqJTS43HvkVlPcCZ2syKRd0P1
gMtCIcpCsFzFdtDx24wF2hIAMSfRMDEh97g14Htl79k0PhfSjz0xTAOyS9KLNwyBlSNwm5EV1fmq
QJNA3KHYDAMbOBqrZuvUZC+jpiat34/UMk4baaYcTIrdde5hXLuRlEAEUq+Cx1L4rfZQHHOJJFot
stGFT3Iv898ERkXQXEPaKHHWMy7FyLtahDXOEGnnBcwMLcRjlIcJTxgaiGpS6YSi1WeYLL9f1PPF
HJxNhh+5anP8GUxp0FNZwbM+85/vPHFfR0DmY7l5DLJUymEONtvtsPQYe/EkXiMLIN1KStaV6ee1
dCWuDQRng+MySw0wtJ1PFk5sYCvU974yn0OGCoBv1vT4TroYSLleToCPaQfJTjAJoHN9V1ydBzqd
hA3vv7SjPGnRCcvRxnXq4pnjBOTC5husu941cFTBDbpwfSc3lh4PPqPKn68zgWcpLoCWFx/P62F2
YkdDGHlUDHhsg91eW9BIrxPAyiSX5GPeTC7guFnitaBQkSl5sctcsq2GRtPqZUSfTJhAcFDIwR7r
C/sN+cGJ9tE3tiZcQUpVOZKaZ7WXfiTDmOa3mxu0IYH3IAoZOtgRbeipSFErc0uWikfCNn6TpmPQ
H6xJ04zNR/QUNhxEnHP7zU/sdRJ+RLK4Fr0HYwohS2QZtvLkuywxkbA/dVE68HX0jdvqwHz1SpaS
SsardlHgMryz0V+s67PSpprtzEoEXdR0qnDWhUWfa5PGOEYsECmGrwanFIROQEg0Xh1vG/e8o8Um
hWtW0rQsb+c9FjxleLfCao3TBqSAkoYvlm/Msd/lTDaGRnJpU0H1Gp8OC/xukYovEU2NLrBuZkaU
blabTMAVdH33y3TmW+f2ivWql7MTCJMkb0s6v/Z+R6qqr3Fm4yoPEj+yTdknXRzappHb4/glu0jL
gmmMUXd1ndBAu8FkKAT1S+ofNMHCV4YTAk8kPGs3MDlEVIRhMW2SEGnGsIW9Spzd636+L3AZIf40
/MhVLqiNmTaaXpIVccEJn+AaVzxbwwhHy50ve3g6CB2ydc/xZGvTRoQKhCXg34cZKq/HY8Ni0Mm3
ErsG0rzMM18aXPCfTykeIPLYpNkgvdDNZ6u+6bGLY2ReNfOXv1kxrvBY5uBNzvLlFRodxciq3fdD
rqxfz9aedSak1TCRqEP+wO1QGlNXbSx3wcQplPfr06CD0QZnS/MHLcna0ScgI2T4c6lSH+Ri53HY
IlCdvME56KsIz/TNSVyciTbsfmj+QuBAxFi7iOB3TOvmPHRNg+gkZAQ4X4x5sdEwd+dzqXRpAygX
uoMTZKcf8kvTDMyC+f3tEtwQurEvWAssnYZFF7EdWumUj2aSDHyq6tyMF2dgVe+eHR7j/jQiLvKp
Up7jqEvkfqy5PG4XiGVMgpiI/xS5ESAek/P2PqmFT45hM/98twBtv0hksDEA9VJbh9OEtas/VO/G
U3+FBEQ4GkVpatjFBhY26/wuIIjhVexoXXFyl5OejCxa1TbASvQ/V937o+3D4U5ZOWzbNbUYBXEo
fJ04H5wVuWBt7XhOYO2ZsdLqaCCNFCgLOlcM95rLeG78Ieek10mrmiDqCSFiok5E5mOoKXK3aXrE
mUzBisj+fYzCGebHw6JyTJjnYnwUJFZX2OfuA1FyV0jT1i+CQvypYdbmUinx/M1db3V0KGfa7Xy1
z44EOB4MFEqqoyU0kA/KRKchSNQirUNYLlMrgVqI2X+4LPRrgelDAVEi3n/Vii2qCyHFUumLnpql
rUWGZLCU13isrzk2hygC4bLKeI+f9l7z+jvYRRm1IDivotnYA1MiaEt+x1qspGsPRmk5NjPsDOxg
LdywCbpT3V1LYT1hyqxLfLBa7Lsz9AdmK0fOh036mzMDkKZOm6l+6sN+i4tT3sGT3rHI0Dl1dN4/
q2sSG6h+PJClnE4u/zmoVM+VnF/7GAdnCxxfFEpQZyIa3FxgTP4UHWy+Q32STghbLz5TIRlUphUX
7EOmzImac1lQEKYdm8hJ9ss4lFaIwyjfLtVZ7r5m2dR/LRtYu0Dvzo3D0dJoSZRTZMzrNsDoA8XO
TAy+zVTEJ+335kg6GejnHxAZWnw3/WfgTiSACRtccvoF6aspkHd6IaGWES29LkwCJ8mQ9a4NGwgz
KCsmAzDKsE4MuXjkSe8hdMq6cXJapM5pttcTl8DCaI3glVd0GnTaKnxQ4nNtMfr59x8KtZVI6mpb
4AqnO/8g/mpYMwfjheotWtJEPmTluqqf8FICXQFkFPUIH+xdohP3MLQ2DFwYhgMC+B2aT+0epz2X
vzcTmkAx3Bb14lMpt6VbXQa0m+T5ZVLGxbGv1f3wftyYA1qB0OED1oeQZqAOEBCJXOJeUnSYKkGH
msUFgIX+nkIKfWiuGgoOMg+4mC7EdYeKNHzFJ+9EDCI88PNLSRN/x5TJIPu1ucncqe+kFcKizYP7
SjIkZZw0TdFXWfnOCJ4FJ/9neX1QHzRfBuRPVj7gw06OPABv9ZF0A2nxchnOtfjF002UWfrL4DSk
cdRv/WYtfQBa0WAfDrIbL4qP82NE6KCR7kS/dXBc6Zej4tCYGHBEFZrICOW+ctiqKqrq+0ILrYfT
PDzIVXFIN7xANcToE2+5JWiLEV/qknSkurL5tlvrBReyu3IMsvoKj/h6fs/tZDI0JtpU64MYXJ7R
4smErLrYSo6sFJgGvs4j57YeLxvQGB/SEiC4+TdqKVp/mN3v244bYbyjytCUbnE1sjObdd98+3M1
zmfHoTCMTruY0J19NE0YyCxlvgrw6qSuu0Q8KyG6UxWYB/o3deJAr5QISTb708uHoL973mnewijF
E1ugovHAvb5YaHZ7hJigr/aounUxiktBi7cu71fYenwbfZhClioeAhDH0NSx6ekqfXlBXVCG5G2O
Y5+uysr9/UBGZCJQP5pCGaFavwawrXqQKCo/ROKh4gxPy+UspfNxNtZGstXWXHzWXrd7lGAFmUdV
E39jVdyCv+b9zyqfdYa10lWJ3W+dmDoIMSvbrwE1NNZGWRlXwlDA69UKx8chufkRjZoJ/RhEwJDv
vDzJW9W3FyvAQx5i59ngHVANO8MZ1GxjrnHrQ4XJ1eMz8pgkpkNnUcDUPT8TSgQOtQGS94EGM8P2
OA5ZZEiiDjiXKxKcQt/V08y1tL8j+SaoAKUEaEJBPQ4g3bGVhpDjr67Btu9fKXioWrTMyle1X2cO
AUWiiGrSGEzTEeQpuklk5k5BXw+/4TVZM/hx2vgJnhdWkbx34f/C5lzhbP1deECX9NJJWLPbCab5
2Ow3PgjRhHTaU932duULR2+RD/tozDNhdi2mokIA1/llhm/8obZbNJx9aOpKo8S0UVbYMbO9Selp
I+gRlSEhZTPTROszi2zKrGbzuyvdruAgSPyBDvO1t7hM7MUHUoa8Ahniw+AXCcR7oeK+LCt1H2NK
s4/B0rlx6uCIVw5vzxutA4yP0Zw+YixAQzMqf+G4nU+7JF2saIdSorikSMTbl6lGXrDwwuHRUysg
5xNzJVadjLw5g8dXVHjumMuGMs/VOCuPQ7zzmGxBZqlKdFInXfdcKTFD6ntn0FdyPRoLD4M+PvRT
89rk9uqHn2QPnK5Flxf1O/iZXqj9ME+6levUCsZn5AQIyb0mIwWd63FQoCapwm3k5U23oTUuHzFV
Jb8P5mk23t9hswIdIQlrsFItBfi/H+enSnS0Q9rLrr085Nc87mAQ1ifJ7cLARLJDbk0GRchiJHKb
yJm6E+iBMtk5182YAx7+e7QiuvryECu2rSS2Js4bKn7jRgZNIb17IF5ULrI+UuAzV+mo/OjBsP3+
nBPvIvz8NhulefvUVEQvD4G1XUU0Lu4s9RsLcp6iW/2DlTl00nzBlSgOdHrdi9mQ6n7rMcGiuCu7
7vr4Zhrs3piy8YNhEw7PaCSfkSxCYgIpew/068ljoCuN/kccRSmDVMDmQRAiPiI9m54KmYQ0Skiz
ltflaS9GbskHrhEmHkj7eNs4kOEnZGsvfyljU8kHKUJ4LUGGgaHJuPN3zUTtEYKbNNvXRhJ497C5
LWJBn1xOxCTCitX/ZxWKxDJBJwflHwlaTSxi/ghbobpDgeY3DHQVRwlM8eF1QFVQrn/CYPImHi7U
4ZToxqZl/OrOdScSyHxdO/yRSVdtGIDabuaFyF9Kkw0Z2fng4KGcd2b5E7LIP8bTqbeJegeLzqGG
4U0Wg4mvywjcg/UIWHZrw5ijJBnxzM+qxM+zBJm/a/u5Uw04TnmTHWgnk5/MAAZRbx08GRa0B6dU
Vn1fNReg9styol9LqkhRBDqwEGS5gi5DBamClHl3+q2OFywFtNsF9djxmOcABb82NWOleNfCJvgG
Hiw5wYS06SwOMFDGuOlw9uUF3O9OrbUAmOHuK/AgRX8NTVwGqd4wJXkAUag/m7MLpaOJkcaN4RTM
93aQfqIMmwvMZrphqLqXBaldJEOLefbmh29w7uHrnwsNk8nc5nbCaDHwAN5mxeIUwuzUHxq7IjBZ
8iTHDf1XSQCAHMF6LZWDe7kaddJ6tBzbfVyXGrecGLe6ireOC8T59mr5toLsR/fpdzdmVl0LkOgr
KsoORnXlJkrLcqLE8nMjKbpAx8gA1sgaqCz2BPW5p5skVq62JF25kgv1vcNT/NwcCW/S86EIm9zx
611laF7SbmElNjaRFljws+pLfR9j94BU8Ea2XsXnHcnp3Ohg7X5oT1PI2EeNUk3WNJDC7HzZEotR
NIgpZCxK2LF+xhhbwAANo0k0CwFA3I1+U0rKj/PpOag56MCVmjf9Wq51xEBRIyLIEWLmyXONOrsX
cdSGlmxyZ57mZgPrqApFuAZglQywX84FlXOmABf4+/1R/p2kATlcAKBoZDMXOThTQ06KIRD3784/
r9Jrd0QcDRZH7B8wSB91Icpv0ebNLyfBAGtkowQz4funL29BsX/WO4M9ShngkKtj8wNZj/L18Lr6
qLjnTOwkJ/WaQBnP+nyjuyp/aLQAtxuRv3pA65BaSb4jDF7qg+Dwa1pljQJP5lmYm860d9rn4v3H
sGoSMUqGxBDmmvJrUdLEvtGEe4V8Bt5dfw4WZ01JVvvaMM9EpWo2Bdy7d8BvpdWQyakwXRMsSKOB
A96ljd9l3x/ZdLVY59kpDGbipYdVkjW4KJVaMfjyW6Vyao4TjeWQIL9r9JLo3iZm8ZyFmOth1Gb7
KwnpshEjbN27n6IUmFyoz4CWBQzqx0CMEwJsqHksmaMxRqjDQng+d51wE3y8gckjL+ySGK2639/g
tjcYQQfYUKBqVd2S66Iui3ir1v9ENegurhbMJs09MKwBKyHpV1lQJQodKoxYRXfV7EW5VWjxhi9P
1HrneF6Dk7YvNLVK9I38SgG8MMbgnSY5SEyfus4R1loQX+LOEn1RauY+s5a7R7Z9vof8qO/y+NWC
6Ppmk1lds3mSbwAFPAqPU+qzwAGDdeiPVRbgJDS9HbC1Bp32NXXVGspX1ipKERHn1hbUIB32abL9
jBMaQmEBW8Kw/SO4PpHROLewTZbT4K8i0/tNdyFRDVrkNx3i8C3pvuH5/QPrEEefAtgMRFTxNXFY
a71NuwKld7LPZWmmkBMKE3QoZHrXeotSqvA4aq4jHG6ObunO9/fimCgySYS0Y9eeePMfu4xcfhgL
wKNe0vzS3zQK+PEOCOlY2bPbPDsPNhTvIoKrmNl4H5i3oyAo3sJSDX0jF/DX9guMUuqh3f6iCbkH
zjsENqwoujm35yFyjVgbSkOQ6cgs0XAM2TZDgz5IPk9BiyYhCFihbncWQEvxjoqMdQJkCCbsIqMV
0rzDGjur9BJ8XzC8nifc0YeuivPeDHGalDmfMy8OGJHrdXTiMxyRKe2eoxg3TlLtOwZ+kY5dBCzS
QgYRMHoCg9Bs6vufYSwRJI8+UXa2+XDxGbr1W9Guch8S64B6w97hu3EfsLIMDh/EIv296jtx5F25
GUExnHRASZkZyIffHwFfOjjny6oyfaY1KN4cgGbAyiSxyTmrIFKOVZP5FmRo0wqDopHF4LKcAeUz
UMGBm5MY4Yfq57NXQkZnfV2mup5mgXzn0II+pJox60PzFj5zFGNtVPNUTxfD7IsNMajz7YS2oo9k
n1HOikoA7zdZrDhcw21XGf4D2bwWzK6J+TNhD5zgIXJHIVDfvXsXStY7r0nz7WmgFa8cKx1Q65r+
qImtZm2S1vsjH8aLtt/KIvQvyDRQBbtcsj2rxM45IwXubLVNxJGZtPT0aGaYTaohBMWfyet/IDMX
iJ/8upoknnjEqrmg7qFkNUEUhR2zidBllPyfjJLPZze6SdWeHoQbBV+5+mZ6/I7CEsPbFYwf8iys
7jXEYYHSZ+WpyRi6gmXYs9eM/YVd2Ixp4JwejNofcdbWDP6KfcnUlqKneanSL0jDLIWbwDlfL4SW
bTjTzqEzphzy4z1H2QLCk/rGe3GhYbHWkcGNbbXwLHwFbCfcYB/q+SPfIOx3wQjp2CWcXoxjtZWx
aRs9J4xctSVg+1+PBGswxW4ZTKkdnuHSP3mkuYCwLgdrRvxD+qlg4V2DvBrgMRLNAYNs2wv8kqSE
Y8NPHb5Om9qLNB1ChIdIfkn7xZO0wB+hxfQTQWegexv7fK9qFbCCzBEtEfxlsqhElXfXEqOxl4Ov
djPowo0OxT5K8aZR3yV3GChU/XLjTcDdzStlWZSuD3hQdF/RiQUsKZ8+8PeXagIoR0ABiZcz0gRr
b5FT0ZrqcO0XZ2onKjw5w86oKhVt04NMQWN+a9MwnZLSRGJnPHctl547Rf7ElXXA8XwyHIC9CQRV
vEVlbmaVyIFxP35BEnCJBecqWM6Z0eZF3z8GPh7dDuz7Zm6JugTQA8GziAOPnIYqKsxZg8k/WgxD
OJ+asGoJFSVXcP1vT6F/2Wc4TUrHPG7OuAwNJLflEmFmLP088sBLNvLOTVmFg9ETd8opKOqHZa2C
t6sDI2ET2KS2nZPp8rCGdbjbrzueg+DbFn+FfcvDeo1TntskxIkSmSsGHPIpsqbSG5YaIqHvrGmU
u1pyZCwGkbYegqi2a34rUizd4aKaRfbhavjFZAAHiBl/Citcnia9m/cg15oLT4Ls8GTvergcuGLt
vMm/9hboVuwB43h6m9Lv7w36SDo8D/RaBY/lHSuc3yJqu+VSeXSSjVSsxq9+1Mq2qXp3TJP6ZaVx
LCtQ3pmyflB2JhUj8HnrYc1zb+hmaOgDLkGIEg77x+GQ9SjW8XfnNeurfwUvH6feOynnMdALPRcb
O5bPi45ltdW74EQXJQeFi5NkMhXiRFvTAcKvZTSgoqMlTEYEb4Qz7vFu3GmmBd4Mcg2icplCySDc
VqO92i/Koh5PBKNP+RgeuO4S5MMIEcQIneENL4Tzznc6WKTD4JrcaMdS9HOKkCPWKsmlo6MBEjOs
RAIYCRW4ziIcuSiHY6r+RXw1ud6yDUuMktvHPsngkUMYTgNc61rxHWJ8bn32YiZI+PNgmB0ZAtHR
uLf9SVnhEuiaURKJXx38jckrMyhNVYSO14VzZ02j5oqAOUoccQ1dEEE8SJM1bvlnyANOTOcHLena
0SzossoA8xgyX2UD+w0UMGuiPvhhG25VHPBWvAtSXhvPl8tnWca7Re+0m8HoKeHvnhPzkw/j1905
AAxQlg4lvBvZ58Iz+RLaERgsU5gXe//gS+gppEw4twfsaGl8wuMqxlBoCwRe0y1ZRC7QqlmsAY0u
taPeDJofSO+NSbuEtA8Whe7aTQoP8IERYFgfsQ7HQGAP9/kFuQDEzMwpKpCgw+OI/baHqo69nHUX
jVuWn3ocpXjn7//mOXCGWzm+0EVxskcxg/fgIow+Ro5ZwF/CAfLm82yGo3RikUrSuO3I0GPjn+Cc
ng+I57NhgB/6PDzg5PAj//vikmiJK146/yv5NfVmzUUhpuZNY6Q/tr16PB4O5K1wTDjw1TiIb9oB
KIeORmsb6DtL0MoheaH6qX0DXcgkntmtytY64uI0StJUa9LMTtRthRjQ+xT15IEPUQUJTevlx6o9
9130f61Thbrnar9SyoTtsvEW/NXS2ywnWd+opn2o+jLJ1r0arKui+CqjnuO91I1kpt/uUr11MOP8
rruYPE+bdSpUwwmEmmsEaZyf5ctWQ/29ddILuxwe1r3nMSCjYYBpY8CT64C23AITKCGeHpWY1jB/
XvTWM2dpbHArJ62IfE3VrC1TFa6w7Oem/Ixgwfy9vKTaHdVG1fHxglDJjpOliChCcptq2liAFyTi
WQ23Q7pvkld2pLmeXYOMngF6ZCjOugBlJneccBhKIgAGhF9KE5W/Sh9LPlHlUeR5psfxyxEjs5L/
nQs4d//VcbQmSCQNjvnP8/A+9BiOtOL1s+iJ8L+smz4uJkqF+shAEkFMwtmqThYnFYscMQweoxxN
aNMEbrH8L6Mop087Iu99OtxPJy+vsAW5MU8t7q7t8BtLXZ4vMPNhVB8x75KrcntdTUh3i2SkVN+4
R+4PiNoFIIEGe/yfrTqeD7lsztJGia2elcllIwmq/jXkYwQHFfzwPmY4EdEs37BzGnH3K5dedtw0
CSoOExE5nI5ljAzWeqIAJUqmQonUyC3f/shEmRPUYNoFZgudFcgMhDLE5i71Ok0r+v/LcSt4Done
wb0CktEvGC5r8HY4j0FYMthS/0JOU0eldLTOYbK9Ycc/6qMgFgW6JyuwUCaxVzc+r6mx7e4jp4gR
3rPSsgHrjNy+hERGzOzYcX/rVSZO9ggDfQG3r5l64PbOkHFS68pkOd7wZEVFPCPq2NcPEYMS4GtU
6zlEdzlib8UpJaiiWZX3kYXhNugHTOfowh9ckqFYkl5ogL4jh9maObMWm8IESkCiAy78wJJV3k9q
be1hlBObwt9XJX/YEmDmNikuBbIr8ra1hW7V5GhiTjTlKqrsUNWX/qwOr4owJKo/rcPqNNWQ/Raf
C9Yx8pgjtpF8jllgq8Y62ET4+TofR0C+ZX5S52DBVxtPu/inJg0AsSoN+qrMI6GAAVl4LsSBb9/F
Zofane6H0SgzZRcsf3GJarz+dRhptcdA2E5Laq2bBwstJi4VckZqqnV8KoUfmtTLZ9gZG1BsBy5f
XxIwLFf7fbzB20wm96U5rmGGNnvabBieUU9tmA2tgZFBkkKkiTxeP8LVdQddFw5yJOfJQcIU+9uP
EY9iHgVrBaeLSZk5u85LnKGflHXBOPuefpksONGlPs/EdahCBZwDZklJXQU3HMGmsj9H1VSyGpFM
hdklFp7z3bTb+30ah28twfKwswoocLAn7zhTMrX03JCGs5ffiJ5Ic1Dzqg3ASoxjOBDQANjYnm22
6/e8GuIhrB/wYlXW0pdzCRSYu1YJsgvbyUEg2wF+qF2yjQqBF+25Y7lnYkeg5tM55EcKtxcToqCy
O46qeuhFP6Df1Tda/rKoxQQ22VvKLzKuGsyC9dT5yZYxrDZu295taKgDFY+SxMx8VrYyPduNL5OU
MubaR4pEegt7DAG2e0YIeX+kOGD9eyPdkwNntU7jNK7HnsRBYuDpw6OqNThZ+zw2TdnIU9jId7Kb
RPts7178w/nnMi3VYT9wD3x2rnu2FKJWb3M58ND9+iJxbQBmCc4VGpPn+c5zqi4MUenV/SFl7YCJ
qoiZC9tDU2jkikn/eX/Wpz5Qh7PB5VEEQL3JtmZ2UzP4VBkKejHhNpgglECpnw6sZKUQS79QWfub
13cma72sIapSsvNcAG8WJE8JJUInQvEAszaJ8cqmP4cl5AST6CiwHcssSBirBPJggWnMrK3bQKsS
zkce5Jk2uaWjQiMQAE1Jy27rKmdZNvAQo7eH7qutQtr4MdrNQ4x3uVRn4I4+RJ78mH+fMFdr3smh
dBi8HQXhFQquawqo7VzQgUkkzRXXs2ELjtlyn48rLsw4YeJOTTxazfG3lJXmGmtl85SK5uzlYm2P
LG9gGvTwn8/oUBjJ/lHqq+UujprPvp2nLdqQaRdX2jl7I0khINWHDls133DYxDMEAOaNrqAh2g+k
WqsYu/YiGVKSmsQINxXesdgbizuX2IFJaiCenKWnvALXBEFfh4YxbsOklP6N+UqZOqgeBp2NK5l4
rIw+n1MUU7N3epibAAQGbyEDvcH9jUKUlPwwywoVC3dWg/a0qrZSV5wuV4Qb0/CGOYvZcR3uA2Er
U0D35cUoKZuw0jCanUscWCSN608Vrx6xoHyXpw72y4NXEr6OXM/ERroVrYh9PjzCy3SMQYofY8ny
1Oawqvu87gvjUm15SH0MkN0yBhiJKAlVApE7KZCSAiliuM0eBWoOaNdFwZeQId9EzAGlCfQWG8tK
yeEmGDgOOqNiU2xIMfIaLQ0U9uKbAgFToGbkK/cUhmRr4iFoBNu0FtF/9OhQkn3/uQR4IF0+DnQo
myD+mGyVZVHRMSa6xKm2Hd0KfznmwVE5Nb/GcSiLx9MhmvyVeJSMoY+XTypSDFPtKUqn2GBPCe9Q
kZC1XVUvbEBKg9rBJxwQcWJZFrXCVUXMufiwa8TGanndjVm0OiPFFx9ytn0HOj8BElFHZhW1zMXL
VdbwJCU1ZzTpgzguztOF/7Mcbbst9o60/+vWWaAoKak+Bw9wV5IJ5HyUGMzOz/ov0qv1AeNpX1j2
irmp2xy1+U1pqmNvLtr2313l5vCjqzDZCAKxDJB2DjM6QSDO0hGNdF8PnvMj2P74E7DVe00a2Uyr
VAh8gHyBGU0DjfFehnHnN5f1ECpW4+N2DrVlw97LDLsQQ9cVJ7SrPIAE1mCI9f3rDPNVFO2rPZj8
OYojdy7enq/MKZ3J6vAjsJ0OtJgAvAH1Ybe/VbujFytZBf9P6SRED0r8zm/ddQp0MnZyzy6br2Fz
bYYLzTHK7bBILIO9W8l+5H2OwZ9My0J8vwr7beqwAPy2lRWxyAVRg177/crQggWOmBDE5u6Pyw70
KRfiZ2L5VvoB8hPxqyE1UOKSJCCmMFD+QC3//bu/saJytVjpo9mR6TMPFn+F9KBsf5cxYwMZf9EP
AtkkPA6W+y9K1gx+zx6z6uJJuwfZQsbjh9fGKhMtSSqJb3zwxZ5Q5o2nGKvV6lRzR6rPt31sjV8A
q8/oLNOQ8mRKtE9WtLNLVDUOQ3Xie3LuWSGBHmjEz3i5nZxId2nD7J6jEkT9sUUFcTyPL9qhR7wy
Fh97T6RsH5S7GIeUKi0PzUYBpXwgLt0K2KNUbvSvqsNW52Hpxi9jslgwblo3OuWeGFkafyzNn2fg
aAm/aod5jzy6WAGrUvrAsehZpnfdioz4GX/7aDF+yzArNjOH2VKM/LyisxqlXpASSd+bLtHClHqO
7E+eayan4cyizeokqOzz9XGUce9BPTWq/NSrdQIIKSQ/T1ceLmpyl/T/676rXiITpbPzgXomwJce
nUhXaALiW/axHeQAioCdWvovUqrwUGwQzde3XX8oY+od+i7MI8QEMoup2Y5nUgp8gJCQgVG67q90
E/e0fRtLfaFZJxwjnY8Uwj04rd0Zr8vFxNavmsqBhim/IxHT/bZkpfkLbPDL6cdDGu2HhByG7jwF
DUydm0VvqMJyKb+zzq0Iwch/0j4V9fgZFXBoi/JmTwtOeZFh3uTVZMtQInNAIaRVh/rBcRjzvpnA
i2xryLoLawgnayHw1mvDuN/Rg6fnOAi+LLnHaFLSLuthjt4DZhH1h0a7w87k7PDjMyJxNInYYE6h
hCrPK1/K8BYEMj4zSqCmRrhlUyyb5FxNIGZ/3tcQ9SQAqYPbMBlj+lVFCvkmDG9LWedUj5+aOfWI
50BeZOD0ENNlPKADR2c8eJPJE05i1u61K755jxGC/MoTy8MXrDmM0FbEDWI2IVy/olfhfZ9teFsm
AD8vPwJlZnSVXmHvX/3s412NZ9vcjZ3DeJsSuTf9gY/IUhr6lNx6t28A2rLNTgPHWNEbHQHmmY4n
CZchF6eYTodmSGK1OQZ1u82viJca6z5iKV8Frj/Xan/c0N2zIQhkYBhRkCJ29T6Nu5NzNAjaxptG
NhJyT+i84QCb1Hqrr22gFWzsiaDG1Flj9P64d4RoZ7RYIYkg1C7zsLx330r0C6YB8sbqNzewRIFv
59y41HWvCzNhs8mPpS0rTWezHV4h2iVWcO16EH/P7Zxwyahb3+cSzqyYhFys5wVA2HnF0QOdkwOz
c33SIipmQwprhRrY9YrOoOFpH1rrG1ZAIDuhR+4psZx0/Cck36i9cQIiV9setzv5PIjQsVorCGgB
AUoq1BuUvY/lMe4uyyfSGu7MY6zxsC9uc4KGWL/LlZIqejAOw5hWp3QwGygsOu4ZOvJvKLA6WLOK
YjvQJoJ83QakT2EjC9FzXDoPfl9jKJiM7gNrl29qiaL8mQyvsCySmlW1dEooVRGxNuCyL/Swb2Nc
GJVEZ2rCVymFYlZSQokJChg3V9JCUfT/6CQ1D05flU1zPvGgEYQpxt/xs9GuUB2m+QvJTR5phSeH
qerzit92bxoRkhgW2duSJtywjcoEh8TzNhePQqy+R39MeJcSVmRr/KLhHcNImfhlzIbjMTaKpHrx
emaXDd5OvWtUWLwoaIFUe3e57HROcW1aWpJjJQMLGKjnln7NV0VCQDvTDutoeWonszkqUO4RarCJ
ZpykQiGfYff5KIUTIpfgwMCzsiSDOBILp0po/vVF+2pyBX7Ctp3lVAhLLvyBkctc0YUedfNjizNZ
xPzxkDBRX+yJ8F48crX+1PLv1WRUgeVLSLoNTxheWWmhnwymXVxFUJwPBlrR15Ohu1E+7vBNUu7Q
Wkvl1tO9UL39AWaUSxevxSsLGpKUb7U62PS1I8YGIwpBC3N4HFAxiFQAHE/31GIRKo0TQB8uCM6s
8PSj1+AmuVYUJxyflj73jrCYKddy3RvfNhzi+My6roMkmNoojJUnqvGIYQeX14+f/Tcn21MRazzq
slPfb1SiSLB1KgqJAx5sCyULk1UTofq5KFT3V5cTR0AgHo+n7bs6nAXq6tiVOmm71jMq0dzZTZov
caWfs3Ohsd9iGTdzDCBbILtyFpS25WHCEKv9WZOc4ZtWp8EQs8biBK1b6bD4Gb38Z+yb0cdAOKv0
zOPve/XMm2RI0dMgX26iRuWRTrGKLdzRdDV6FDiDf+Uk+KBkMO8oNGpex7EiNc/6RGZzKZ+CvN8I
AJhfY+vRFaQs4qi5yJBZqIH3bkOenEPNPy6l3oQs0L4wuwBmV6pWAfN9wvGTFDx01QHZo9WRXVBD
+GOwNxQVxvQ57rHQcwMLmNO2SufXJAg8eq738QNqxmoH6m1QpksDh4D2IQ5ZXJf/rsXgE/GVlPqB
ZRQ+f8Ar4PNKqWfsxlyHbu28RJnhbo3ySGnWy2vwQvJ0ryEiDycyUBQkeD175FM2t9srlkIea52a
tP4T5aZXNgr552Ugm5L2T/8jb+ZXeChPbpsAfhzqO95AFuuUAJHE5l9GFkZ2IJcXBfLRYxVgoCaF
iX59eaJSyHCW0vzUHz4Qysxb3TjvVTQ0VQ/eAVfhWARrLj62uLHgfPUsvlukOVk+lBbj7LRFITNw
dilIWAaR3XOueg9ShmtcYMHTJdZgxwzN28GQrHDHxcIWhvvqzI03cH54/sj8ezgNMrTDMD0OeFhR
6mgSTNgNXJpuQmB0aBQfWDc8wp0Tb6yA9N1X9ZY0/U/g1G0iMbkpnPMqe9kxItDFbsIVho3OzZyC
1ZtebYCHXeG/TTXxA8Y+s6517cuAATNT5ZsY5WTOlVyUM83PxUr0zKj2axx4AMyK3z4k3Qy3/Jun
BK4lvQvrDiXjkk8Gl/FYJFw9RVKFpc86719OiCyBn6Y65DUKsIwjcTVlE2f0mMI3gj8QhSneKJxr
VZgq1dSeT9HUFOnDsB6aHxl6Nne6+HL7ZncoryB5cE1gXqy5PRZ2MV1TUveFZcevE3Wy3rRabA/6
ZSGQdYChlbAxlPdXOL4pkl1lMcg1xXFDHravESQLK4J9/oUuZXz7lb+f7yC9BoLoNv9002medFo1
/0PshvSQZUSwYbbh9nv5sdYXiQ893Sk3pK93WIxKMg+b+PUvSK/rFCUTlon9KjWuBs2I7UwrqL4z
K0p8VOCoXphJxg4uBTkDLiVbQ34c1Mn3ExSkgap6owVvRroF+uOM+F1RnDfGzdbtvrrgf+VKEHsJ
W0N+hN0hs4oPls/NjyFNM/tEeU/rc0M1NlJXOV/YWXmtbfbABMBnLwfdDaGsjiqFtsquOGlwXFbW
7ofb9qlpABiK2NYT3aj5syO6oY1jIDZAaH70d0VAdCGU+cPGNqWs7AjCRi37AoxLcW8fi28qOIVD
7RKwJ/yFGgZNQudSA2Jlr8lEbvZ8oJLOZIxeXQXChrGfT+ZrTdo0o+sb+jnKXLlzKkFANmWJwMlQ
S9KmZ+uBnbzCHNYIIpiExf6Yq1KyxzNkyEKyFeHw8zTcIcVJIjvjy46oI7DMyiphl/PPS2/w4LHr
2Lie1xICHwJDARJm67IkXXlMjxyFsfQqNynzDYkcgzCKmv5uHCltkRjpKRmJEoElOPvV6d0sehRb
BM2DMo5f81HVT1FC0+7crNyfQKWd0TGwkQvd1LlhMS94HH0pntQNLG9MzbXbcyvdbuSPzRyIPzoh
D5mD6qYUwgyTSLgEYGPUp9bvAmMxgixFqRalqDjI1LoN10NfMYLcdKi8VToNcVYqsahxXtQudQXn
bJPksjw9av5/731tvpsudzlAcqI0HOwpAZ6m3e9H/XlfRbo3CGsng/QWIa/PYVceugvTUA+H/Fi3
qhvg/O7bvqJCdigSIfNe/EU+d9WpT3g0x+DYyPUyU8BIjIJvvlfyKppfD8d3wdbPyTGYeW68+opg
YN7B+7ED68EjYKokK5gfMH6DeFmMdLl78+iCOkZtqYyDEiGqN+8LDLIxpyF0DCBXPYEDQp9+dTTZ
PTgMt3tEpaUxwydefOR+WCpQ/7QBIKKv+qBjA/nzoldDFVN4ycdwZdiNUSnxSDePuEEEaLm5nGmL
OR5ZAq1DgNfgCRDcas+0ExMTuYgIEpeXgwjC4CKYPP2BadWJd/WLUys/rA2T25Se5Jbn4kfJqQ02
yNohqaZZQWLiIlWRdN0anmiRmoGmArjl02hu+r8U2FkRBOBp6gLtHcdQ1liCDBilIoNH661D2jGL
I/P5gcAmuYJ8Bef91zRODvQnz+p1Abg8MI8T6Dg6fCytsFnXNcugwYXcKyRjFXUoajORPpuK0wVZ
rrKpq435XjCKJ2Fei83lh+8x7ky90DGNYzpNxM98w5PJpUT/WxoSCyeZX+Sna4jglk9NR6/2ra64
X/j2X2SE8peQkaSnU5eTYWzUCXWOGMpl3n0MCMARNtLG6qhqoQyworA3L7fCs9tDoRZADytMJaUu
eAS3Fr1pL/cZBIdhDHZHx+7kJwv45UaUIQuIGkXEdOFDEM1OYMNxF9P0FURP1PEhj1aTQVE1xXGJ
uVzg27ePGJbeY5flwx+zlEvNllBEOv4lHc4g3G5ZWmdUgRgN9zgdrQxxZsYN9lOGNA7A57/0ptaA
PJFEC5j9CtsFM5Ls8k78uLAVVl6jPlj16MwT1Jay7rIT+TXZElDCR5837A7Hfage5vIFIRWdu6oQ
6060VnX6cIG8v4H/BExWqQUS3q2nEM+peI4D/MCLNitV6NdaDNSE47QXh4h78BNjIejF/76LDLPw
Yi9LV7vZwaRzyt5sqfgc0eAPbsFNITWen0mZG70sU2gKyc8GijyNdSgOjyfso55OqybsEiOq72U6
y5N7236JMerIdko6mDBSbuepxIM68DtktgMbnOz6UB7SNKsXKcQutF8+DPHYxu5QcdOsUrRtwOwJ
qrtPuxOiLCDEBewy1Ga5xB6KBv+stYjVShdQ6UqiCiQmlMhVlyRxVa+6U9XzGiwLv//2uvhoV1dd
2W4mqX8LR1ihZMEWv41ZS07Exkh6OzKbUToXHXfIG1NOW7TdaeDhg31AiJe4Uh4KjR0VJUNJqg6E
CA2RnK5isc1ExUZNYWNOHT4wJ39mkdVoEDswBigkVrCkZRwKCaYJVHNki95j/NZpZePhUlGzVDRm
QVmJuINhlSjm0wXgHURtYp4fbxCqlKeG4Z1bxlkX2/05NkqHHoHaido4Vr0/OHlq4Jxef3F2vDhk
L40oDS9Fr1laT64TIGdleJlk7xdehktk6Tvw47bEE5s9qOJ/D2r6VgnAzDtLExXFWwj+YtdBfoMQ
ZrbUdpGWJayY3C2VM/sDx6u9C1++GA9J/v00qj5J3mMRVZ/v0/I+GZ3+/gBsoFjQA3zImcn5wVFu
SRo0Uc1c9B0zToO5DBudv/7XRx4L5JnIWMjlq8XwBZhqB2zD/yg+0tkESLN3yLLZ94daLItWINQ6
TPZylDebxGCzqx5k2nb9zsOXdo6LUjIYUsBCmhQb4tI6T0Dzr8C6myX6s14fRTYJ9jV569W4sZLH
kB/E71D4DgdeYJ8qcxpTQ9M9WR6rrP9rN0TpVDByl3/Zb4HB9pLIg3AL0wna69FPypNJDzvNsj+O
WNeIT6MiQ6nJxZf5gHj5Nfsx0GSTt1V0RFeYQQ2SNBkzG+GzxuCOSiOLAgphA4Qho5BphZwpgYgM
2VWuU9zvouAPDJKygV+QinjcT4SrkLtPdJvo6NPVNPZ2WM3+zrsaIS9bq1SYw3AcRW5iZlK2UmZ3
R5hLwqmudKzXbhfBmgA+/KziCh1CTbCLPH+dX4a3BtbRTQuUO3aiFOnxNsm8NSSNy8D8dLUn0Bmg
L454DFNGk+2UgYOyXdAi0Qae2/B7DULbZ3LqyERcLyPFi2qS+UzIJ1ZvECg/YNpQSVqoWac6aE16
QKbJCf1SxeiV9eJhjOD7lLS6jux7j/JBhQ9wlm4+H04NjnXcLKSSM8xz3xsXnleeDCHMMeHjChCp
OCiTXnAwS/hVyBKkoU3njYA8AImYfla5y4AWRevHu7qceT8UiDYBY8hXpuygWJC6g9mxXPhoe4A2
QpujOY5yl/i17Oa1SkyFMfPcpClny9a4BqKhQMpT1k491LBcTv2FlSOqk/tHoSzKBElAQAZh6nk4
fASXJrzpHgvPBK25F99o2zwlmhs+GK8djS0WuFE9aOFyX6kvjIGwQ7Vcey0CI81uD0s1zZJ9T6r+
6TJumt2j/nzWEPeUFUmmrC0faqr5nPuIulEAROAr+bIuTaOHMkQCfnHBlTBWcvtTmnVM66YTFhld
e87lOUIyl+dnXIvX+jq7jTopTl2TjNPs1aLisxt4alGiveOvipvxH8QBakDRgMk7+Bz9DEmo50ee
GiGMGx0WFYydVa0ujx1/j/vazZXHXkh5SLw2M93ZJGetFMjrqyOmX4Y8obJX5eTePD76AFZ7GVZU
Zt7yLJm1g4IZNYXRcNrDDhK4KPyIIC0FVSHrxYcCyKyXlHZz8vWY/r4/LLcSLFZ4mv5XV2eZjQKK
bWlPWcRwU2cLNwtt298m2X9NN2bVXLwmKNn9zwyOSt7Wy88VbPTk0xKOZMWZgltLhjgUJQIz8a3e
NuDocD11A5M7pDMA6HQ0c92041H3nm1rbBSSh0jhPjTegPbz9Q/XTcpVkbdmL/7ChvcRJYYdW15Y
0krtjpyn2k5kLN25uei3fC4ipDZBXwmQbylaCL53rJHDeFYsR0tAmm8ILAmhxWrxgSfkEJI5xZOy
5+3BD3Qud6WoxVuqsM5KJPxqifISmPKdZXzJa/wvw+tuW5TBsNlBHRh0qkPK1n5qt0kzHGe0q7Sx
9pKJBmKg106y56uZsliTzxflKkhq+MM/fpSNU4zlW++9J9z/Z4zvZQl4Tr2SG/FNhUjaCRrfo8Vn
MvBaitBYDvvVidgPFnCM5oDC/N7lxMI8M6uiHICJQ/rWSYFTU8hUVP85V8fmGclsHhySEQgmIPDn
ECX+l7X5hicNms7kLfjoTt0yE2b2WYJuCuGjAKDUbvfRMg0SpjohcqPSYi8pmpW8yYoivUMtdchJ
WeWkDbHZb9VFsuLTdL4FjMISTpwTL/mWcJK58ySKI2TiVcnZcRVLxQyddZ865d/xQrqYeC5eqBFc
jvANR+7ewUvLQtmONw5q8p45MOwoRY8Y5uQglSFM5LbHZnEWf8EGXoyN2fRwXxTyaiGUFMzCZjQI
UwK93M2Ib8WgMa2P4/JC5WzVZhtK2P1BsrKn7/xeR1H3QnYbs3rAfrPXJt6+6Sdb+Dd5Ji54U1si
IkAwyFRMqZ6LLFvDIQwkarsTsE+xGgNngqFjS+RxFLKe+5QJj1wN0kJOVDX4/P9UcBoC+drHwXT3
LwvUiXrS0gRfc0FJZxyRQAe0f0JR7EbSv0xfPUKm3gRCqvxjYEZxR4WsCs7OawASo81ji+2rHz8x
BiuGAlrRmPWPNR3OiCQKUnkBSinOVYt5NsLb6H7kbRsZj0XSPjcgl1zHHydl4pleaPw3nGReX9DS
DUoNtbZ9yKEnEPtGVhQ4BrqzqwpVZ8wxI3yYog0FQKMz1H11HIm/DXkoLPiWc6SZKRkrTJHuArd1
wkJuTGkvosOWgs2wQulRLxCMxVK/ZB2Tv6qRaEo4zPV93KfWarTC0Tf5JRbQrbXbTAMNdB1/zbCO
YK525A50uhRWTnoQU4oA7UOFs6HH36jGJexOIpeWgMvakmVBSDfd8SPByk0M9wd6L+lZaOBlnJ64
bAG2ra2mj0l5Obzd6MQX8uyDyJr4O089a75Mid6aOvKcfDPQm9aRjCoEacPef6fR6rZM3jjqvRB0
NRkuQXaNqHC5YYxg3XYf/0HgXknv3npwiKCb5kze+DQ7gUJf7KpS/JqZtHpIpx7slfjPP3Pa42Hx
zBR3mWS5aMEewx2IlOnLSDtocJTeWkB397uENvjVeEy/DIOQ0iXBfdh7/vbdWp8gFreKO8RATxGW
x+DK8howrLqrn1CGxvT3S2EDm91d2TGT524mhJhkEbqqoWLAqsKyOa1R6U2oYP/wEY5RpioKJlUW
175HJu9Y2Vti2aDfc9pDfGVI2OTBTB49Cz6CBE+A/vxNchXfYKEmSqXAyHiHl8/X055BeS+mRzh7
JI0jq7XWjxKvczq3VnP6yasBCIa8sRrI/iARXzVBduUBEsExvYfYRlNVP0usJ5m+6x1TuSxcJonE
CM42HETeQjz7aoprIquhE0p0vc6mbPpI6pbUfwFlxXm29c4ITqcJpvH+ykYK48YpG8Q0bjLywkKD
gx1c5T+N82LjlTiRPgdEx2mP6luA1kuq3GxZJSNXLi0p/jgMgryVc2BnwwYHc34PqN2teGL91gCi
T60MOFX8HBZrk3jfTMnWdH0IMPavnIuKa6M1d9+J28htqhjQErpHTYWmDqm853mpont4W7lNeEZ4
+slVWMXtXajDGCcK20D7dY1mSkH88BzU6v9+SjpWQFcAo9/Ze3DKLYa0wgeZr5G94mEW5xG4U508
Vnsdx1zEhF4h4bFvHmi1AlDIOKQrKqpQNKyIho73n/OtAQEPcCg0XlBx1ABqJjzPVlXctUUh3kMo
DFenwruA/8bvGQDNkJFAXRLlaRPR7grlVJmOeNNKrvISXylcnls+a779L8pJIitdrtjHJtdL+0M0
yzDtoLbRrG9Ih9Pobezine/ghl/P8kmw04JScKpPIDQsskE580HsHhaGoA1GMxd95EX6o++RB4yV
hJf49sLAB9HjaOhV9CTxaisF28W3LkMyr/rOiC4Jq14DZ+3Fv9WQLwNHkwYOs1FNQ/ul6ZFX4/jk
cV2H7AwlCNwP1ypX4iyE0g2Cr9xjdygD5oSMP6WhHLRHyKy5pR4jWhWxF4R9HClsFxAqTU0Ikoxj
pqHxg+g5oQp1xVEDveIU4Da//mIEhlWEUgJk2qA4eHyCsvMV9AxqWmvg1Iqo8bGfpa2bFqJLq8pB
a2JZmUH87TAe1Sd7cQ7AclBR2729MxAwd9t5MPwHcoacGDXwlCjWlCb1lQR3/2uAaYfnAtduYHI5
E7QcJewh/DSfFCUddXyaAGL4414PjVXR4VMarcQwQkrZCutPo0XYP1RoN0THnBPx+dNhOiH8tXcC
D0LJYOaTnLtQ1mtW6R6EM69+ECP8PWSp0F8sMPZ4an55wSPYBUGI2HfhOMWyH5ttb+QiMPbWMo80
dQTa46yrTIG1zmCk7lCSWMsKzACszj6YNo9peplENkrvmSvKoM5XbOOgk7xz0uYDfPUEmAhYKGAE
6JN+Rf45IGruu4eCqey3bIIZDaQzaa5thNWCk10wp3W+cV9gFJ1ll/G5FPI2ObrrJg/tf8e8va2I
SVulPC6lnzfGjAymFauPwGdNoCPZo1yEBmxwvogwhnWGdau5eSQtU9xjaFopWF+B1jdaXvWVohGW
Mcq2qZCun1XClzmBKznO5Gg2ILGChFcUKiSEd6aN3ewRdBvcKGOOtbWXN2F9vMLBZiZkDCJnwiYs
DlTeKkBrPM/mU+fSNahf8FRtwH/eJS4HStmrJsbHM1FeswR3fAtMMHXT1QLosLeKx5yS5yEr7mtH
dzm4P+OBYM83vLE6anmKzsJ1+9OGFu0IOGSGZBZ0DpfxtmRwY8Wz1hgsOdLLK8A1ygdwol++m0of
xJIaLZmuinXfurqOQ8B4uFQqCnWzFqBop/kc95llDF9koSB3BEu9rgu/bZ/GpWUhMO6Due3iS63W
nnrB77Ak8cBHga3LlFQAp62y/WNOj9f/qtilMhh3ytwJncJiPiUWkoWDgjH0hAUVR9v8+c6lXHHU
+v11+72wjqIACTfncZTfI1UJcM5TqUl2IO3ZPVxxrs0Dj0u/To9W2+FBznPFr16U3kbmimvpuKOV
V2d4GG/z6gO4tcnGvRM7TVQuSUyZzgKmBRuNeopntMoalx79bizwnRQvD/o8c0RhoGWGTLbqb7Cj
c2YaN0lvBywO4K2GmoneTqb6jcmxmrHlYUg2gH7mbwKh4jeIniT15Nb09cFgFTG+DjpL0ke/WdB9
fbz7OoNhpxCfSxOOV2Yev8O3uxI4SDKjuA7X8uH+khG2QjsuLyQk5RmfL382hSxyZmZg9e5yRo8y
WKEUYb9Ij9jTsmzQpwiQeGJtwstTB/rQycm9SfIrIH2VKBN4/RI47TNmb2fXtyc1eBcnUYQkB3F1
dbz/mEneRcYo74nOiqADqCpv/yFrFICQJT7LNTEi9Jfuu/CXD1pxBCI4FvjnAKK5WB3clK1V/iZ5
8E4tiU+w4fVetBqfpu6HOdC/udO3SyO9FmYFAQODfi60Z9lNODTLoN3K39yNp5IRSMmciSN1XR2q
BDshUj0PcBshQDqdN7uCizkVV8CSU66l69OcynC7soUBGmbPBXKowGu8zlVjjjeHIhtJRgZm7h4z
Y3SUOavlGsEdtJgklXVblSVVMFpGrJ7Nlnjw//8rrT4+HDMOaQdeTu7xQNJnk9COH/AOGwsogMLa
+raf9IccjESWnCmSZn9HeUgK+OhNhuQrTYVUhF/RJ7zHeh5N67/ubpjWpJSUEK50/Q/MmzsMgU4/
Q4mBuN7NW1BVw2nSVjdJ3G+FPTpfHA0gLOjC1tJWGxhDy2Efh3HTUeF/kmD7MqHMCPXKMGvxdV7C
D7RqOKAE1X8k+8aWpYllIyZmexT17x+Dj/lYuWPTPqqxjEApHEQupdAGPU8Mxd9dDsJ1M8JfmYh9
vgZaS5KUk62dlMs6tp7WJGlftQgaAQEdv76rJ9clK0gR/wfXi6x2GwiR6hMxSRe4V+lJ0sRglEdU
fSgCa9li+nom67LaRbniPCbyoXO/xUPwfxoNStf5u7jklNsaTTdlBBSUTMzYdRMp8SgjgcfedHXb
o7hiqG4ddKPMW/1FyfoWzYxqf8tSw0eRBRl8zuNo3F7a2TKppjbiI6KeBLAptK8LVRa6NwWFXGbV
fAjnIle3B91aaGrDgE8at2GhAXoqefXxIB7/tYCot5UICQjp9c4KpJ092Wua/8TBrFTtdPdmls5N
ZxcSn6tuqI4OrlErCvVxaHe12h+VNxfXLwYsonLa6WSmO5f1I9LxBqAsHRou+XqmpWfk9nknBHWn
Gvvp7+98sqO6d/6woCWTeGSlzRM+xoM1mrF/98wW/zXzp+PTM2xs/sMb4gvxrAQiNLZRGwGdud7G
vjYAyK0U1xv87Npym9i55z4Cl9kWHiP+dqFNiQVxIREqBSsXaWrgzW2Sb5QXAJz8N14K9sV5WgWk
yPGHnBnzvh0DNe/kHbnDhRBQt54/GwCBv6PV9F4t0Z3jiAFG4UXq57749/pFJhuXMdEEG0UJQYDK
4u0ang1RCptTbzmweZUqpaM8c+mb0E1JtcTTiE17Qa/Vtw2zOqJqDmkivhdR+Dxai7LihzG2atOf
wiiWB24ZIUO0X409YrIaSaMZpkblsIt4Pr1MS1QOSOpFTNcNqAyo3CYxhkNcaTUBvqorF5NK2V9/
mkH0Z89Jw9z+HW9MMm9jF+TrVE0kWJIfhPkCI2B2+mewc6x/JkHh7kuGTMM6jcxtkNY2M0p1GaMY
SWGvdG7qaPr9vnByNGDMD79kxHKwdrcc1T2n2r/Rqj9Sb06g0eT6imIrSv4/9Y8guk3a0kt5NMIg
sHkIFFe0l3njCWgIhtaXlSH62dhgh73B+I4bTkqYq7Qd2+DeeT3k8roy3jdDZO8DvzHlf/TZ4nsS
CFv4W+4S53y9dISNNqU2sRO6Ci5Kj2Bw+QUmvEhKalydttRq3IDm7vTOy8Z8m+v9ysoAvsKygh6G
PrBYm22bmzfH/596yc9esLPcigAWv//z7LT/td889r8bUAw40Ch8TgH27pzWv/MPTt3cmjI39BZR
KvSx3mJQDPn5tBl+vvBQJbrNHHBia5IXZxeAXR1iR9Sk0d/k+Z0PKMxz9qC0hA0BO1qah6gGzSAQ
WgJOKG7huDLPxw+eb7Q2otcePxTj+piBAwc9yBkbiTQWLq2JgeL2k9SGEhUi3nf/B6HC1dH2wS8T
qWq+KV8Xgwv6M4d18PRmUW3a4LxAU3ocaFBKyrRyqlI2vwCW/5Cejg1tT6rzw2kcaxjBu+zmYUFM
zkx+3+6/SR5tRx948lUTAHAUHLI+Cjhy+Aegk0f9iKsxCw4XHsovX4e3g7uM6te+H0VnbTVRoxnJ
MUCPdtbozxMiH3dShBUJft3YSRhanrJtfY1ru6U+4vbkjadXqJu0099LY7J08ddBUFwle/91MCG5
zP9/as1hC5na48lQ2B263pRWiif+qX6We9sd+f7+wcvliYOdCGWOfVE2rN9jTGOKxsM9XCV4ctU6
bSnKrOkE1BHzdZuYHoKoc39byS4FOO//p94TDbZDsRC9DUkoqndVZTEYnDHBx1tB5xCZalE6jgWx
H6vktt2z4OI3p4NCo4Jqx9EkHuAAejDy/BWdqeZ+qYdjklpGHX+S/cUziTirySKkxGZwNbuKsKsz
3BeTVu3wJVL60dSJejPQjkFbkSAdeONA/xgMnupndo0Jo1vAHHtNMefIkh0N1xeGpaVU4JaihwaI
1d+7qK1vl+V0uw5x0F4UstPRUxh5YtqLR9HDjpcBWUqqqnx17nvnnG94FCrfMqZkEboMYiyds/aa
KjHcQ+AUktdWWuhL/fq+t3l1Jjcxej7XdoXdYIksdzQRpjHrq4/QF3q7cB0YeJwf5qy25L8hkn+5
YjIFo7Oi0sXutyo5UavRGoW2zuC3Y+3lvGfBf5eRmxq/NS5hMjQROd8Fhw+j1BM9awQeglQNxmJ5
n1dwqGhSziojSJ+QOfSRBmmkI+B5za76iLLi3BUXgkD7JUMEb3KSsAAK3nZ7sKVYil48ksQnMxa6
2JKQw7r2GoTNGnEmPBy5BZjHAeTX0031QZXKE8wJWF1yPi3q9Altgj9oOtzVdAG8p4OStQk3JBcT
VTITuLmqjVMcUyuPfWo9qBNX5QTqXXHvcYc6+dby7hp258yZyqT4Mj5goOvf+CWgskTJlIz3YTfZ
RlCB5379EhVqoUQHyDvDGv8Y32MXxhi1YzGo8Vew1kb9ybfMMk0lQmyDYVBA3rqWboF90zDtUORV
7KhsAxuZwlBemRmhJ03PBHxegbMDdvsUcMj20Hdlpyxps9Fikba8b0C6lhsnHM6okj0+cYBcrKAz
d0U9Jp6UcmSyor0KpS/rp6W1L1WRErt4+meVxerwjNnonR6otw7zTg+sVkXM3LeEwTvNz6B44v5+
UwsqNxdYKc28XWglN+SIpYftaCI4BIIb2kwumwcYA0ZrjXEgdiUYh5sejQOnf/VU7J94feh3nbdE
I5nesIIhjHtg9X8/CUpD8asoTCPxLfTeimr86UGmrKiII4jrHzEUTBpZvJsiM63OAphznCwNuC8S
kKiNLUJ+83oLoXXCMiWhoX3U4VbR4u7nkAW01etXQBYVbUekKrr8VUIXRbUeN//Z1HKKrrGdmKkg
Rwd8mj4iGF0m/J/wF+9vIUJDWgv5vJJfPZ4gMDxZhdeMMqQogeX5LXJIvwxk+kEiK1xZDVpNoO4c
blCjJvQsPiPdp8offdOuwcbQkLnTkMBq86yXkTYtpmKCbDhynqpopuI21hkYox7Yqm/sWY+A65MF
8Ne7J7sdCI1tlS2hdkRcFZLE434USOCe4zerAaV218HDVOm0z+u4VzwLh/BDXe96wmaQOmSiSIrB
CBdMA5PmyFdn0l5fSKizfIFGEo2nngntj8Pdbla+LMJ74ZhuB1awF8WMGl3TqbkuRlZQjFspd0mk
/5NqP32XrzWQ/9UPXOj4clF0lBPRO7mNu+og3+zUchQ+ul6GF8E2Uqnkms7zGrpSCKD/gcNsNn+G
uHp2hoLX0kPKbDEFWGfzF0dQPQ2LdiEKAjQTw8AVUgoVMkL6AptnQef7MgNbJMcDZCxt2tT/MfHH
LG7nzIKye36vgzwERvpkiLX8RUNJmH4gSPO8OxEt+MtXomL5bFeT8P9oRmnuZH+ARmVWPWnfhoiw
KBQsuAK1n+cT3AyJ3emJZevw0EbALypmDUftbauyIXr2CrgxaqKwq9RCZyRqpi6r1hvpcAtc13ud
R6i2q1LI4DZXoCH3g0+jJbVzzwfih/XZwpTiDYpOLw434nSqnHAx+2pqv0e824p3P0F/lZFqCr9i
K9LmyjNa/B8u93TGCzO7wifNDK0YTqxABbwvIyVu/1WKnfalq4Qf5CETPuO3Gu+6N2NTqKqy9G7H
nVgzfwUzfDiv9d5BYe2iESpqTjk81fO1zYPbKfCXRTw7DdwwqsGlKaMkBIKhDraSP1TWCzVcjszq
Dt/99HUWWq20opH2N+asRNdYHY1qWI36xRBct0kTYT5hY9acDPz85t/j7jbLx+4JCZRoNDkL8e2O
NdsW5ILAPPX2pJTB7ys66hK1I6TpBLojNriaDL7L+nNUfdweaKDEcbY3gjo5t+HF0gFuepp9weyc
oCQPMTv3TnhYREhmoOjtlvWL9qa/BlsgzlkyuVAoakRbA5XOnqzXfMF8xQpiCpwf6FvPPH144PgB
qyppT3CLNEWv8vlDI9gHLF24Ccr8/CI1wITO37JngwwMO84Ea3vI3kGTQCctIq0g2ILmDM8OnYMs
Gvr42Yn2GisU6LA8dYJqqzqzZr66o2Darhc2ChiLO0UQWNQXnrEA6ao0TB97GLY9ursMNkHiUInl
tKfF801dybxVMJRSuukjt9Z94Pk5o/R+L//j6+ZuNTaYPC49mUuRnlZnmZqpnaIaGctOcgF6qaiI
LgbHl5DQw5K7+Xl798iop3VG4ftNMbAI4Ue85iOQUUG0E74j+Nk5R0Vj7mzXCq8+M7iAVZrGOiOL
hvUHIOMFXrzThbCWs8hya1/xGnNzbv+020l+O9anOEy7O/77+QogAUFMDQP/muxby7fCTkAPp2Ng
SL1F+l9m1rGd2enu2rSc5OzTHWDTfcEyRTWBzq6ZRbP4PYM+a5AARHw97KQDIH/S1O1r+fD9tKYV
tNS/QUfXn3rQNjjTp5eS6Nl5MHYAFQNOfV88PacEOLhu7zoguq9iJNjpk5z846BFWK3J5Zd3wFmp
/8mlH4/OWCPCvYsZQpzaIENSR97UILk1y+61oMkwOr+81HMHIjD8JBteKm3dME4lpRPn5KMWpzi8
sr9kRGmtEPwFCWFs6gSY2Rq/dd/RULqB6Octv2iuO2bmqjYxGH1N3DYb/gvwkvReklWacH/kYPy5
P49tacJbjPsxkoMea+M7UTrdnjsAVxev3J6nsIPMw0ocQbnCEtBclFEnGpKOnCjQWVSwfSU7YdVl
kj5FzC0yrI3aBqCvRxGcHSgUJSy0pwCmA2LUs1b3CQmryibg/yKbcJT5TAiR0pE6JGwoLxjVCXoF
FnCxp332q50ohhXeuCr5Wmvqpj4ajow6aXSaqRMkZxekH74tumuPr/k2Ia/BDJ1FxevM7rvKMsdW
nhn6I/GpCLRB/dcXbuDeLD5t7zgxpVcGDA7Myh7WDlLeuAExyZjij89AktCu5vrtnSMtsnVwGI9F
lNDkoqlONm04jJu3P1O+HW8st9XqB6Q6aLhgxc128zcPzL5BSaeIi2SlYG79SNLBE6zLRMdpoXRJ
Wqd8J2vBHeBu6wDxLEnDTLPMB0dKvXVeTzfQTVTSyttxISZ9ZCphkWOLPPw/tFMPf5lAbT/idtFD
2lOD9H8Rl3s50c+UfUG/mEfdzUadXe0XLgGr7eu0QBtavGKLO2L4buidDjPay4PKxQRm8/Ns0vlG
Hjhv8W5ANP3dFQle8D1jhXY/Q44natTjNZRJ0qK54H5ng4GCmGHBlXFo1a83DcjH6MjyGQJ7kysH
quGb8cJIcwU6eEQWU8W2v5/dwYqZXhrvmNZQFqlvb5xSko5jQGHSxWs3zgogWpXe1jbxYqODZPqN
95Qbq80L9Nf35PrhlnIdJEdyLM7EMwNFKrJ8SupiIIA0GOsjaZmhjS6k/0XbzefRQIpehJla6fz6
JZBLkrDU06H9d7IBgY1p161wT3dSQ82ofSqPORORHCf1Yh5/psGqLLC/khgxxZCUG2z5MIxQWVNS
44XCOOOTaavAIsXWY/qIYwwiNFBtb426hDDFSmRO7qiycQ+lWoJKcFp8Cz2fkawo8iEEFSRntJId
pgy9aAdK3PV+M88fso2hYZoExchjiOwwx7WfvVfvkqRV11GdKUrAEVHCE0zXJF3hcZNr5xm6tFvb
g1sBXb+cm13FO7TUKi33j+av0/SldalVHwgeZgq5OQfWKW56xAsCsqHLMCM/RHBbdbWxRwFV0U49
2Othba2fTF8qzae6sTd/5dnjN9h/aiNMSM5Jv7QRofjvkPabrds0M4bEuWrVOynkKZsfca9nDj0Y
1R3b/eIJB+jF0x2Yz09Sld6nD8R0JMrtHrWjEOzPnGBppDmCas6+9VjiNcW65FZNO/SoCulxSIBb
lsHqRgm3y4rgdFSBCpr5xy0xTvY9wT5AD7yWx04m86o4xB6E0AGv6mPg/yX0T4DFprhXiKW5gJXf
4MRIyiu2OWqoyZGQYglzIqZrJgsoYenG836PZc/WRvnmz3DXdO6EbYygdAGTMYoOVrfwuUcGPhrl
11lKuC7juoGDcmTvIXI9Pg/MtI7s62KoZPXn4DCtn7hR92zTvvgGWOlrdZ6R0L3fhlBEORgvVdl0
M/DXYxOQOzJEuFOt2ZauKhZxyENaEYMCJxf5ZNiMqvzBzg6Ywi3sZbE8XWZUvhxL+yL2etjhXKm+
xqDkS/sSPwp0/7xWR3cn4KbJbnMwdCw1ZFno5L2VNaOojPt58Hjb6jzbfevMaqH0ilLWx0T6wUQ4
e9Gr2au9J/gBu/45TYwwF0M+NN354C2Pn7KJt8x1fxDvGVQfPHrGVdFuLn0pF/+dNlYmW3n1PweA
VmVjtSG5etM2/2qRGZAbChcvaXF36KbgjbQsvKKNjBU+iDScudUG72Q1oArMukZ/fLt1jdqhJGj0
jFoKfPM/AiZ3Ar20HeZmGr8LH1/6ZmDBDY1fS0hZjECvomiqIqsuvEovDc17ZNPg/5zhmxJP5bl+
0cbA/91h/jZJiw5JGlIemiHlJPK7sJ38xl0GfOaJU8FxWWPP3pRxRWPMjoRMjLsP1JioD2zS19NN
0u7BvSHP9fg3+XWWNCmjMYY5KJU3ebMbfbhvI5OT03WgfGOW223OhTB0l4onbRcLHryDVZmrtKg6
vHagwK8TyIAGkH5ny+amBjZ3Sk+39S768Hc34UBRMLelnU59GlOFfQF97vWHJC0FIBS0J5473c3h
OtV89vr3VvMfORK5NtD8ZXomOZVdS7HXphip2e74tHXee3H6sgokfvu4Grdz9vGjVPqqPKMSJHOl
xlalBW5uy9kxky93aBeNZZvQBIn53euTEHt8ifVUcUmwKUD7id5GNM8du7WzxFX1I2wGDAM9x3o8
ro57gaBt7VisNWo5nVlV5XO0PdFJg5LX66qWA05jSCxeCK+jNXrmDsF3APa2sh68bJCrzmf7u783
MsyDrt9abnts/MMclT0PbiNUTveQQoVbOzmVouORiW1+Tf6FrmLnLR3ZScJG5EBHD5Epy63MwC/0
GsiDJ9TnHzHNDhTziGGLV551e75wdXTVXR9dgGlDENQ+7ww1Ajx+yMOtS5Z7ReMfbkeKJOop4oAj
KQmz6CfRVz6kUnRjRqYCD0cHMe4FQOPSDDdI5DU/0mAGHgQhB4rfjhXp4iKh5gdKVwYaIEMKPQwC
U9J73JD+ayNg4k7Z6d2YidDR3vzAXLGFUIYB4qdMPPoeEiLlfVhDr8zOqlbNdsvQZxVa3oc7w4MT
Z1GXF7+PA/dcW/JCKNIun7OBAD+oOALuhaePAFp06xgD6tUK6px9y2XbvwFRx3orRasoKWpbixjb
SaogDCJUdFIsO8I8QdNzVQJoikzScPgjMMtFU5Dh/W/iTeeO7Ehu3PrglO3/tn0CfiN94lGCElgm
3rkkSAsdLjP3YVc5f7PpHyt5Xcw9oJ+F3cj20z/2z52yGPBMg2uGvYGONBOXX6TTp5caO3ulfR3M
e64M47P1ZoABQJVK7Rr/+NVS4PKJi2/tcKfrnqvjhvFzdI59QlI+18g64WGV+xbYwhPl7mq2ytEb
ylHD1RyypR6JKb//XrRE+iIiVgyKfhDJU9T/Q/+eaiRsk8O8xSnKaw1ZWivzj0PzWfxFC+tAvRbE
FYs0JmmotvWIZUvRnxfjmO2zpAtDmh1FVJbqxBIGGGvUWSlEci6KIddFptw7cPFoqXJJpGkgqSEX
fPgI3L6KBnVoln/BbwMkX4FFj+NVuq1Pzu31xO9FQDm3wqjHWmuFfn/2iDDBe5Rhe2cgZCmuQJ/b
SW22cKpBQNQwsCRHTsh/uPV6e+0piuxpmFbAnlfOJfVSrNoy+mMkaUCYn4pM4ax8ZsdU1RCSPajW
OBzhS7qLOi8eMHB5ICt2qJm7IW/4UoPKOz+0F8xwB3of3BuWN7KLpDU2o48bWyly4a6L7ytpP2Yu
vPGmLOHWL3MihovgMxpiVYa0gyuCooQ8Y+W2+D4sZpS1cRWrQRNZ3vqZMIcB0DpFQPDi4X7egZeO
2zUAp1vYDLvLtSUdhNErKrNjXp82K1ULlEemeMiQVg5payI/sKqo/4ZQjG6Mz+t2EjBlhbNa62Kx
vhRRX/8jt4k7NkkkNsBj6s88E7sr7vmeJF2HotPevslChPTNbvfbezUz/SQ5tvemn40mgvEVqTbe
QYZU5Jm7TX3U6EHSQQt65bmNy2mI7wgv4m7QbRJzQvzc17rxH2FyohKPXchEP1U6gEji4osIRPtT
MghQiaMFvyjdBHNVeMwmwsi/KFe/1r6eTLWtG8lhxbxPphFPnVymflPL2xzE4dnLecSJfV0AjNIc
sRsr0uU87Q7qnjFp8MANg1EEWns7kuM9oqb2Q4/3Cp7TJmI1WkK/cbGq+RN5wpXZ9KsUldnBMbx0
ZkewCSdcQ6nDd287ctN9qRMZKpX0Ub3HjuuBBF3pJP//kRbHUecRoLOP0g4kxXmjwkEW8mxm2DMC
3QLaDglJFySFevTrrozggkGJg1QuQshvOAtsSMxoC+ZbzC6C+K6QUFyR+ATwzzugjWtnsupE4coI
kOOxnFWI6hcso5Y0QI+Z/EFyjJaVzKPe+TE0C8dtRg6h7zHXo3yaeOOlo8GRiQucXnBb4brROw/c
oSLDZyIFNKx8h1AfVA3py9sCgO9lm8sN9r+aaFT4JeWfxtH6TTVqHD6SKY2ht1SOoY4zsm9OcldN
r79FqGwxzBD8FX+QhR4grn9IBhBj9v4wBOkoUjHqsKOsuCz9pQx/+1rYY2YGbrJkFOyJSut2SxPV
26VNz1O+jIt9Uz+AhOWYcMPoiVYlaq21mIjn3NZusKrnWmvDAofSmiWgw4R05xcARzlPWJ+cC6OG
/QxxzTJA+RhJYW3c/+tRDGLHxmIG+86jN3q7euzjBw/yt35EQUbqVROCw7Zqgwx/BBWuE2DuiYe7
Ycwm4DrilpA1/qoZKhkGHJxGfmkovygPG+UvojgdWIEVfENv2MLj3xNz/I1YnXVY3hdnk/6o4vYC
LZfyABl2F1gY86dLgSwhKKek045pL7zOusg1UQkviEsD47O/y84+f3/tqsDwJqGov03rvtmCVd/7
H3eTJ19k153OYJ7D7keIeHS0x1IJe3OqOz9/0vLt1qTOIuszGwpHMMMtFmD8uLIFh0IbU10DraFH
pn1XemEO3jCJGLoYBo1zjmAn8tEAe64xetYS0232QyuywY//ZHB9oMyECjQCOCX4HU16bB61B1CI
Ss+wbh9Zliko0C4KBQXpCt+XDohPXEEXoFCuS7S3RghhcG/QaNuy+nBAbE5Y8YcCRAcrsrNQf7bd
Ib222b/2KGxVCXMS/DOf8dQkaxQE7RBuE9FxEhihdlbniydPZkqWA3Gw8zxlpbdVO+LozHL36yP5
/b4VOs/8z701/YNOMvMbM0sWdEta5y/YWp7nxnkGLmZ0C8qe5OZaH59k6dgo6aY+flAoTXtQSvWr
iQtMgpdGPJW3pIQCYOu3fE2sQdZe+ICWKxHG9CZU8WVMqG4BOhBytp8c0bNHdo9ZyWzM8pNI2NUY
YPRfOLMwt5hPoL+qcCoePKQbbyJP170T5+citFGZzl/cgAGndlY6KcbAFTDqe5mUd0P7sKaOuPLU
GokklPTyOywxipB3aNnvTnsYu20b6EVXq1zfyB2OHIHwzQDuvpH8HEE6eKempQmqrGvlSpRAqv+X
vK6zdOte+Jh6bUrxpsk5MJCzAebEC1P/K1rBZpTBhE7OAUIZSp3Cd7346LfMpzeRBzcBVD8IuNZh
PS0lD0zVNlkUfCxiTqTieGCBQxBZK5b/Sej3oc4gvYCg6fZkGA6nXt1I0OZ1X7iWfZKuxqI3iIvn
HXY4KL6+0TvP/K0MzVumtnATaB48oLNW7dgKFJXNkVc4PREugOCjmg8rTQYQppAu8roIp+J9hffn
NF1HwyD6wpoGVDUgdbzg0kl8BuMQSOAwWmqo4Jn7zKhM44UxMnW8IuntkEq5c30FZZVhEfYD24jF
o5aCZum7m5Eb8IMq8Zo01v95WvwPy+VdEiWb230A4ARdl9iXYoy7SSdx/xfzHr1UBBi8KWqBNv7p
RjqWponYCb1iG/7oNd/lqhG3/wGg4QiZk6b5Th11rQxcVTHJ3KeO7+y1ptaIacTSOntWJKBjvBjh
0cE5xpbTTtC1kTtBT1tE/htkMvytd9QMhA4nNMaj3urcvYF0np//qygejtRNJc0054gEmQkvokDW
0rArURf4jhVgFm8dcmCCDIkBJbnKjXegW7l3IdxlItKOMJIws+Hv4Djt+1dzqCL8Gb2trPPKl/jl
DMaOi/k6qPhmBUJA0bO6cyCWPCz7e23XXtelC4991VlJxM9KQtczvsVEtex4+hl8wJmXwsgWdGmz
3sXkh8wO71kMBH9gOivY9vS2atstm6GMUeMbCQUTiQVZGwhPuWmGkVSeyNpNJM+EhWjZwSJ3k/w3
M6zrCdig+NPgbIWpbHXyaTQxxRF6293eIun910QTVMpMO9pHIUBiXi3MCRshwUDE3+eV5kEoGqsg
sA5mlIGFTKDlqdxpW0RqeCF8NUUdEGyOpuHO3fXLTUnZErMHtaimJNgZx5Rfu54MMsuR0tSzc+uV
4Z0L7garGZeoi+QqxybjXPTmy61RGVTbe5/QvupknN91EYyR++WWgYLw7Qi5HuqMPcqglZqUMLKq
uWR2K/yG3BZCggsMVbUteaUCABzQJkWcGC4U4VWrvTyCvAB6ShRlKZ7u0RY2E6sy/wpup6jGnkvV
4OKAEYGUK66w0e6dNaMrL9lrTwhGHDxB/82cGocBZFBEnXD91png90CSPhz8KHqYLGMlO4XnnjMA
/hltcdaKxlKT8EpRpimuZ6q6yAb7Obu7vGVlH9JQdRWOX/098IrQiUnbR18RBYF4MBuNfzknipG1
BOWT/dER9jL6V0BFG/BeB8DYKXcZRETbENfI6qkYtwOEM6Z7ip4ieUU8+Nk8vMej5uaHDsgsPPck
+YnkiWFxhPtIPzXGkBzUjuNW0N/S07yutKiZpHvcFo3HxV9umSocqyWT4LzjxdTsG8iNVXYZD6nT
iY7IRY4hIIEIsednflHhrxP++m04TBY4TRVz6y7W7T5/mq5YIDmz+1MNCoz3vxodGOFw4uKM1A/0
q3t5nRomEe+a7eVISmj4uPN95H7KiII13xZ0dpWhUcTF64OSzcOZnHWHGbEx8nBI1OgJa62tYbNH
2n3u8X/so0yo3QHdRTOKYXXaJiApvdRMQeDLcWGw9oD4O6/N+4WrDl0Ykc3lXyDkg430a65Uj4ke
55UoHcFgxTpWkMA/RbPfTnZ4zn76yHhasZP+ll5/j/j0iTe+WyBoWgeiM8XiuGBvC9ehVJqCtaKl
wX184ZDaozgK91eUltYX2Go9Sg9HLYM63TaS9qJYtUu9U3bzsvT+QRVOvsITBjjbBli6RwPfWwOG
8TDmCpBSAXDI1bMs36lMlVy3hMIJF8QBdt0mE3mEUTjsrLgZ+dbkaRJBQ4N1FEXee3ulvqK4iFIC
BwYkQfEfqJcEKQOj0f1dB+zcc5q9kdSwKEnJscx7Moe2ELmlsvvnUAyU6uag+RZTCEEOwY1JhNEo
Wv0qr9EKj3bkHv8Z+rBkyIYQ3q0Fzz74RM+ZzXIWDl6rjaI5wN1z/FzfTbi+3YJdNpmxGDfvKbnW
gsEsCMtajmqRHHv7t8/x3Y136YQVxwX5/lDGyOk5XQxvCGec8p0QWBjCiNayuQp34HAX0fD9LG2F
6uKC8qk7i2HSWCpQ5PovqmEufTF8VXBTRTKhcsGJzJ6t1xANaH7vH3VcKejHdQDQeeEW8up476ST
3dIPtyAS1Plgr+N+7OlAWXGPxr468TOAX5sNi43NnTzKNkNrPrid/di1pf4FKhnpXToVXXr4uEX1
+BaWX9x3DdLsy6pjnwkN8YMIHx1GkjAhQerWHk37kx13CgsVMmMJGAsGgLTyRY1gdjF0Nozx0MiE
b2w7K9KQ3dEXg9eAV/fOQJF9YjLvveb/FD79r20snUpsbRC/TW38uVFiU+izPj7wMVLhXxVDwG5O
X+3OvHneV2gZ7RWIyXhjkQT3mpYjqEMHYpVXhAjXJPl48F0s1NhF0Na9hFKPtznvLDR6qU19rpHE
Qm3PIWXsRtT5+/wStr0wxP/wG4yXkkfOm/+zLGv1yNi4+R1gq+4WqvROG6pjfvhAkM7VxK4diqSM
T8Wx2m+dtm2Ne2RqfBhQFHB6gvmWQE+VrVGgvjxfES2P7c6gARR5yHARirbQoc2wwRqiwl2gdBhK
2JxID8RqyLzQL0p1jsnPE/66K6tqkH2JRs9cFISCB9C58GuVvNfY5UVbwmZGaxhW+adzmHRA/48i
XxvvlK3X0mUyTQahsqYX9JHCNTVYiy63EfTHKOZkW82pddgq9TrdpqQIggJy9uzH5w48OYsJqtBw
o88xo1kY9aWSrDmB/6iLIPFc56mlQEOMogWMy7SuBPuS6tZe5sF6vEuMauVussJg3soX0ZSa6uuD
fpxp5NgzDCtnOvG1wImS5ViuiIrxQDW6HN/h101DdW6IdZzCyr+hRP3p68YXVra+e2Dxsv02x+rY
C6jXgYZY4YaoU4eJgv5PdQWZZ2rW8JYH8iblr72seZPufUk05ceomvnljCtVzbWklKGYCdit6xfE
S3plmdnM4NRVyXkOYV06+m9xhJ4K59kfOpG/uvcapQDOgLM7Ic395i4nKeTZJmQ9sNKUdyoRSAx8
erQmwZOiPgjoSw6IP7BYHGoo4+7lZiyAN/l1Xdnkg1yWjKrVqAn/gw+JkxkLvTcBYDD+tpt63pIg
aDrT63QyWpuYkFhRY8Xn6Nfma2FgRQ3ciJP8E+eBVIRkCIIzXKXvv76k50cnE4MMg4xDFtLwzcEp
Z3CEIekYHePTFAVf2kHkfm/uZ97UDPcktayRIVxnvX/krOPh8WwxERnOLghTmFzDuZawDruNqWxI
s+VSt4ysRFTh5h2lUVaqFu/x/f+aakH6IO7Ok0A9qJZgdn7hOswLvqLw2h+aQY69HbTErTl1BtOI
nXIviTkqQ0t4ZrsXEjhA0OJTGHYHvs2oV7s5bQ5XkGhgMCNE9VWqz0kk1t9HzuR15L7e60Pn5XFM
tZmwtDN3oJOhZuSDjG/txMfo9GNoqvTwY417B5fDgn4Rt65GM1km6DfCRrXiq/P2kmkSs2xlTlzq
mon0yeWZHHTY/H9f8qXxXq4CrhuHqQUvQ64h7Nx7rArUSQyNaRps6bgOSZiz1PI7BNYuJKR8k3ym
Gu6u5Gg0zMvrdzFPH5fHGlDJtk5dWpxzwiRo/SOZY+2uhUGN4IVyceJPWwD6P3ukaWH25KcCDIZl
oyLsdxUKpoIK1QbgUAqcWzASd/Ay3/Ko7wjrdD3Qv1M4blZLgccJ14cA31cPJA+JYxxEMu1CaBfE
fvePy0QQOmDgvcjuDVaI4DanqnDm1g2mnhUCWkVwlRNvS59nrmb45yAx9WwTl6ttZvv8k70rCj53
+a12OhgvGMqsCgxht0um0Q9ftaREDfnax8WulE2sSHE5jDeT1LOspUq+NzGWv2dZihHq4PJxulHr
lJZrIexqMusd9YepfQLjbLDC1eTA8WpFL2ofadAybyxZ8F8+zsnZfg/d1HS2iAsIIcp80La0qOHW
VB5fpFwGDXEG63V9JUwxh4XxQIdYlMSWjFTv6hyrYDa6k4sBM6DgNU5rdN+iywyYfMysx0LFQmkV
uOpwA+ETTzWaNOAnp3njC8GEdmHwtGqwiW35ST1PFoVz0XjXJWJJ/HxSyT2eMYWk9AfSCELPWIfd
EgBYUrj1OwUfPudLCwiYC0MB/H+ijOIZnY7XcDGEzwjuWcToJ2Tpn05pfGIy4EXMBvMlC26K5v4J
uee+xYiC+tgvG/1NnPRivW5gmT9TBqCqKCUISvMCVRK+81uM5EAi8dmIxhxhSq/Te5kWeipIUnc/
NKiVwYI6TrFVyIvs77MZBPXI8JW4sqS5YQeNwjAvYq5iMeGWkhZ1zZ3hmtf96wr5iwaYRLVd/NqC
zP0kpXl1G67GADzOy6OX9f6xxOE2X4ykdQVxRqgo4zKbzAjeRVM19fwGl8FfUirg6JlsL4+b1TI8
mRnMnWdU33QfZDxTd2+oksYwSUGDwk0xtqV/PNLX3ui4E7GgLKa0Kls/GQDHO0iOw5GsDa1SHCo8
C6QZ32p0MC0ttsu1vviux7wdDNQiwgI841TaMP13RPaVLOyFySqtzrcjkf0Ti2OHnShIPmnXvtK9
tbDw/ICoVYLh4hUG/G3bmoOLnyLppnv+XrKEYtvMTRYcf5V/l9CSEm7HemrCx+MLT20C+d0nEfna
KKqVS7BxwG8PEI2gx5XAL5hxwAhDHc11CXrbcWhQjUMXsFRqX3GG7O9yzEw/oXD/QLrsg1JdvI7g
bsyAwIxMLc1GIjIS0ZVKLN+/IJzAr7GhTrwXYJDciklQyKw+1y0Tn7wyH8Fphk9x4iZ0unRn/3qv
2A+T9ASqUN9TZUYFBJKtvKgY8hRM5NXd+59x4ByKhFx00jlpmfOm6iqpFkpGyLr9JoZbG3YAUL38
PW7Uk/teqtJVhu6LNaOT/N+yjHMfajgx+UesAQWyoQEO19DBrGLp+8SlB5DJO3iRJFijJvQRXL+Z
7/7F61e87w1MutDEqTVqLgQG4yIsBRfBIGe5XqQh2/pYXKfPWl9hMihwpad3P8dCF7788roVktuN
R+BC+iVAdfkJyO3L3USpW5Xt8tyf46WQmrsmoPRsKfnjIv27vYCdVPWEv0BIVlAReNV0AQNv7a4q
TFCi6mGGlT6XNIm00Wr4EO1nT/mYpXTlU8+rlq4OaBRf2QM4DB9j80VOWM0XHYYlFdVwYmCJidB2
CSGZsWnXTbgZ4qF9DMRY2ckuTOdXxpKr/zVIgI64wl21S0ONY3Qk7I/EV3qGIcI3VcsrChXOzpjT
So2iUYKpQgD24ubuZHbAVVGnrIND1JFmGKyrMmLNrAHyeWP9YRqR1Jhl2n9nLPRqWTTn7XUrU9x4
mpfSUs/RvaFa8t2VLo+smtiIjKqu1G18zUlcnb5DT0X7UZaIBHFBYbAmIJ2tAOf8kaXtuTP3BVFB
+XSmSX6ObYzdjBzaNgipVlENEbCiiQzaNdB9a8P2HONu+TV7KbA2ObGKQ7kEwfu5nWjYOH8ZESU8
BQ7RFP6p2Opw9FHEb/VRKHBR1nStw2L1NJBVVx6LynRG8etOzCfxArFS1LRAl645kNCoMxUwgvks
NIaps0ZONqBli8Voo8TGsw+OFTLi34CxDYkOK3rorzfK7oiz3j7rh0/gHEJxZk62WOaMxgygB8EE
5ATz0N7/cpe1zCcMLlZV3puRra1IZmgzPtNfAlOHlszJ06uJSwsVssUjUD4HfuBilp21C/8dkNJg
K3RksjpprZ66QI5Xr3Mz0j6FX9Iia52gpocnikbXx1UNoFwrK4PljQbIUDh2g8iIOXN6XfZyvHMc
B4g5h9RF1nt+9Xxk9Dq7M6lXq3Zsv4PL6eiedeZS42PP8uFRnpuf2huT8vGK5SVFKTSgP2XzriOY
0uEp3Z1f1a5CNdCELwwRfPXNpREIq/nAnKhDmQCCKAo7pmxvshRjvJifMNdxWhrveugcFWE5dvui
WQHcZP9cZWpntyiudYm820Bumwzsx+YopNAbzYp/D65qW7cyDh9b6MDWj9hb+Ir9rI7QCdcvHC3J
EU6YNgbKeF851EE/VrftqVdxyD68TyLRykRqofg5VP83BZJd6pUTkM7LKBBDptCWxR9Ywrzdiy4U
YF9/EAY4LkClplJoRwM7IKTDYkht7dX7kQhTLECoVlbZWltu3L2ZqCgyQUOthCO52v3XNuOAD0uf
mF8xG0nExlzujDW/tRg00yLIi49YnYXCQra4Uh0GuQJeq1Hv9wjr3inMIH3lW3PkLN9l7MCc+0/b
vWcju+TShhzWhIs7gH62yAuUXQLoE6O9TYuxkp5SF6MvOe0gIOcDoS/3VzXuj4kzGCsDfB8FGw2j
rEjUMbU3qiAec07Vw1imgzGTJk+3xBIcsSXuVltTjcrmuum2PSeXUxX5P+JX3nRecC8XCwb/s9fU
h4s/AXk6lF7OIyNZ7wAjUM4AgI6rzVpPxKssqLnSHkjAenuUaXP6JT/pm7jiXxolQUICyiKMSPOg
d7yXCMH8EAD1rDAo0Iie3XCAV4wP3vcMGM1fIhluRA/EDfmhXg0wftoWeyDdrjiARoqqGM4CZJ7H
isjl4VLO/QuNgHwoigAdKi15I9XlGRQZ3l8nPMEA2fX7LzhdzBlB8D8lczUTjgXZ6HLhEIKtz9Mb
Rj/w/QYpDLUH5G5YSpg7iMZTkPjwE8Q8wmKAN6zJNpDZxqBMOjllWp1JEn9VoJug6/kZ8zJgen5Z
DiBJSL+/JnMG8eGQsrKM7XALGEVfmGTcr3UJLdPBDmgCDaaRlD9aPX7VzF91+wSX+UDtnunV/99w
kcj6/QpemBsB3GL27BUZwh+LvxMFN0BW3jwJYtJ3l+oly+MU5wieKqRSAg6RYYR6AKB9OLo1x2Qc
grbmbvTQzh3zKgtS1/+hUrfLMvn9FazNmpFc5x0JTojXa+x+i8b6M5okB/1I+0JU2Xtczxumjm0Q
ObkDqMI0dajv+MzZcQKBYneIBX1B05umsvtLJvw2nuP+gWPgysb+RSzyz9PIDEysFUUF8/wMhPbv
saKD1C39tWyD3bpwUn0EcjyUfmQEqGh5i0RrbnQLHpj1f3tnFLJ5Kdfc/wnRJcdewjqFLbgry+s7
4VZY65DmCNTEP33lOnD5M+Buq5hR03+3uTyfrsldkFjSRSkOSnb6r7gbjMZu5QQeSiXSP0EZcJIc
J+IVfsX2BhZf+jbNO729khOHr28rpqygdDFzIKE5LAtzGLCPiu7wM9QvtnOTwu5dXaohK0MYVoy3
HhOh677rWRzGqQv03C2CItxNLK9RPjJw6XexuutEYNGDySITzIzyXjlyxvbhM+2Suxzuc45eS2RQ
d5XvGqFX9Ek3adyNUYjByVsqhcVuRSjMXb2rsgeWiwbFv+M1Zqg3OzRs+B90Crhfi1aGEOlUp0wr
bap1GTCU/nYm6tInkCjHXm6WnMBf9d7u+F+DkALTzMuB2xKy4K4+etpWU0RfUDBwHh6WaNAj6UO8
/zFmOPGYvYvEZw35weGb7kJNHqvdJTF6VE81REgqo4SOcMgXcC6pti+XXK8tGQioWhfWPi12vc4h
ZQLM49oRhDlrx2cszmydxFjCSJh5K3/3ANcy7hMSxzdJ5OdcBkl8VlA5iSHWfJ57H0aexv4bsEqm
Bi8MbR4Lz5Olb+/zqGQ+X0eNVS4dqohiskPbaaVI4z9YsAHNqi7Qd3xaunDrCJM47KYbTfRZ/HmO
Dn5Wbem+lQniARAtPYDcphGh7YeX4aagJ951vNkx3Ex1NhZyyLMostC5vI55BaRCY2np++xLdC9b
u8wT/9R3bmtFzHnduHo7d/h98md5jQXVSg0jywx7TokoICRJcDfVFBxPQcYe+iOhb360MHNmbNZB
LLZDSDjiuRsDkN/7zaaKdr/a5BT/xL2gtTEUh3UGG6+GM1FoR1NoVWwDGHEiKyUiO+tL7vD5he3A
uWc5+UU+ZpqzJnFNQTJAX+EyDlDQn0qa/6QeIJqAC2pr0EuUP9b+NpL+8gL54ra5OQbelk4jxKVA
qoEQmA5tofFa+guZNu2zd21qK49+ah5u3XC3gvtBGQVVCAG9DS9js4GyBmHoXqxVPgorFGX6wCjY
kMUMuCyfQ7LDuqbZCXzOrY8Lc7iAXNdYVcPjs+CJBxswmax1s1+FRKoE0LxHpX7/MEq+Jh6N3u4v
UywDFJt89mmZwtkYkQQo/utcUiwLau/du9u989Aw7XrH0yfj7VuWzlhTD8tqctd//eFkqaz8zppm
SqHexODtH8WGowFxRpdauy552nsfxEXoKJIT1V6hDV/HlBCQD9ms3Ri9yspeqMMr4BM5dSoxIKgE
dL5h2OXN1PFUxz86zWX/LHtu+2WlgFxM99aC+uhwoKtcgaMClZkEY5RNWgGQW8BOMwds0Jzf7jlR
g5jt0tiA636G0q2DSs7cTHUCjSXYr3bCFrPkGPoN40PMKavEcxbqxLfQn+gg2aIzdPXsI2cuSo7s
AZRVEwXlGEzs/DsmLwBOsStyMsNCleHe8LpFhtoA1MLD8PrdEv7LLXPAflZTN6SS35tUqr4zxcKs
ciESQPbrsDi2aqlY7nZL8RVRw02lDXD726TAFJUN5Dp5aHCqWjn2fyz6jM2LS+xZSHkWId0YO7bm
aLW9SNA9hHHf5oVAogovjLNLRtxWfw6Luv/NTJ0DP/sWuny9eMXxK2HCfaU8TZgNBbKGL6ctB7NQ
4WYXD62OJ91KsLmDtgKbrdefFfSv71B4FSrEiaNQQHZ4o0L4mnK40xJq1FNPL0Qt2Ow40KJ098bf
EUONK4nHmKEcOFRuog5a5aRXg6FO96Foiwq/6nV7OROTMpzmDBGUMWCSEOh4dT+bwM4v0qAsZj4T
Bu1q0d7VQOLD+/55nPKwx/MDpPYj1ZY7gQ5csLAIpArAOg1roiSMoiQiT1Qsuhm3W+8rW/c1wkP2
Qs+0LY9jjHarco4NfxCW7hc64SaUQZ0zOQNWd2YR3LYXm+B0jfec7l6PgGTk5uWUnqaQnmJY2Ww7
3+hun6TNW6yRS9nHziztjeyciAeiovxAFDoQpOfGJjiu0rYLWbb2HdHy2+pkgy7Qi9EMKh+acB6O
Q89kSP0WHs8OjXOiMsrMRQoxYUI4PAFbDRvkresKYytuXlcvxw2d02c0qBijMlM02kd4Mp7Ol2GL
dp+1jEWZYXqTQuXSgn+kpn6YawEvW7eOCeJeIH8MXYB4jJWLaktRXmZ7YqC0rIKLyNfHgP04K+Kt
cnwf+9vjGf3eA49lJO72EqXy8R66TAB/n/OjQgY0jrexpEufbbVWV8utZXux/FstQ0WsV8A9cVj4
IR2Cp7wYzr4/vsqmxkGFQ+MdPa1Gb15ZfU+BHIfoDSAlDiruFpxXFT/XXV3MuHbBkuY55Hx8FfZs
j6wIoRzk/x4iot5Gvw9JRC8IJksZ9nezhdS2l9g5J+MEI0d7VipxvDSdwoqUfSXXajyeTD1XPaIL
1ohVBlBuDny3AnJmOaF7pttGxQyQwsFkr9MC5p1g735bkHR1BxR56qf7Qm5GDcukg2whOn6TNh4Z
muLfhkr7pGRZc9KaxZu0gz9zaud1p1IOSxXCcnt2FUkbXmD4COYDBqJP6X9NilyhVBxZYeKAGG87
4C6lmrjdF/q8CYrCFwMiRdeGyAILAP/9BbyOv9sgLsYKCqYgR29LGISg/7T5TFF9WjTc6uPcJw+j
adMkUkEm7iZXMCo3zdcwwsNG5FyZApGKi/BAJH7Rrtn1zfnvywS+lMo65DmMBgNOZ95pk0gupYyp
8gnc6fhi/kSR+7ybrw50ySNXuuA2QwYXn2VIP4o3g8R+g9xN6ksX72hrubehzrhgFhunALgjABMV
oDFEqBGn3CDpPsJyR1SRLDVYSmgBt4X/DV3b4putdxFJfT2RH20NpO5aULSncW1Dazb+cLw+fDxQ
rH9rOg09XxqHvQS6HVoiSQPZs37mS8FMYMrR/09zBG4LMjDzckiv2pkquKum70OlXn56DlzqrwQh
CdjGQ/g7yS1oCZlAMEsK6YRR7E1KpUqwvAMq+nuBzVbILpUeUsuSSjQqu0/R1vMzyyzkzWaTNZsn
Ys/18t08CEulpe/NFiRV6Kt0ZwzwV0RZMeUq/bqBnSdIblCwvb32Rba21dVgV9A9Q1HSqSrXvKO1
9gpmhmPWHS8V0/W6oRLWjYifhL7TAPRjIo9FgUabEgnVOr9RAJ3KOu8X9rSfKugwY09pwjLd4iuh
Qpg5BlecNXbxUQFsnJRCPd9gNecKMD4oxluk8zViXJbiTGVqswX95bi1td3WBg+iXauzCxmHMyeu
wuGtVYe4qieXN4KrKjmCD+j+tcLYJOOY4KjH0GJ9GJEHvqoCCbboOq+K9YTuSfsDJovcSHMc9FNS
emXLIuTjQdJSCPO9EglxwyYDA+4wYNNCUq+Jv/VUhE8Sr+nfstLG8kbfkKTuQcjui/LPBT3Dw70/
nSPzLUSdu+nNaZuSsdi9i8W/MyyxQMmXrvFPRuMwRMREfuhuDs46VG+IqxlPpCmvT1g6GcKZvHBa
+dY0O5VzOas8ObkVOY3hl8YTbigy+OyZqUHRXR6EhCK/1qM9Zw1p9OH0XUhChrjRicxFM2qxDHVo
B6l80ui9j+P2Qze+QZck5TcbuwW1xWAuoX120jRLr8wsnyM4gORcIBPosZiXe6LN/PSIRv1E0Ws4
cy8SCpdP3Wv6tSe0uD2PYMdK0lTKebsok+Z3lCsSrW43L1GsAL1m6+Xjv2eI+eqdUSrCiPl4rSwa
5mxJLfoiQv32Slp3/rbDwgcB+ruGCrK6Co8cQezl6XyiZOw5DX4epy/dAndluW3yfxhXTuhYYg4b
fZRxRm65R1gbY8nUKwD7idICMpfovlVAs42qm8ac747cdz/gktpeRNGBQhWc8Yz2e4xC30YptNt6
6OvygcvOovEyUnHBcwa2KwTZaCMLvUUHecUiVBiPmYXlbUjlrAQc+k72bHBeYr2LP1JY5AxYfPbI
cbXBVkdDBxdEY9QHtdctYcX2SWivXd63IN9uhsDzEhZyoAnclXIhPH5XlNt+au9NYMhmus7AUL5p
rgZAwj2e+im0Y1PuW9ZM5fk1/o1vLqv7yUJcNeIqmN5l16blQGoPH8KW4EkWzYBOvnPyPtpg6LFk
4vgbKIWZx0W/M94tZS8T3Gm3qPdPSv+2yS16jNTfYA62LpfhWV1VvInXr5r+fgrVApKFBT5xCiPa
4zvV+Xd07D3LVTKgUwjTgRDjz9hlCnhO9vy0H1mEpJaOlTf1TCkwCAxx5+ngKXMpyvALqdS5sZRO
FAbHt0FkNf2q1mXpGvJtcJpLjQ8RfFCD1AitniRs1I/vlLqoPgTYATnkft6Mf8y85fpEVIclqNvr
slURAVBAZfTLF68MJyTBz70WWcaLSwo/NtP8NggeVT9vXCgN1sssj3myXSCtCG7nrt+4AuVzXSLd
3ShrPcob1mM+KnKXDhzMXdlNidvoTRJJ8RDnN1RBhmMKxuvAHYgKfrV2RDkmOjZ6ZkxmKt11vfxy
Kq0PfEP9ZxrB4h9KB1M1f62SQUtPNQUDTv5YPboW+OwesESHQOg3K2NdiLNe0jZxObXhHmssa66f
wkMb3stChWlDjc0bhx25qaISo2UeMfCJU1fcEtbBr/0qWstGEK0kejzZdxAF343dXiIkD0DK9FjO
qTh5jPhlBfZFyfvfZUao0cuf61xiLt1BvLYpu+rEpAYzuXZImzGomtO+Wl9T96a9aK5qNCOjudrj
NBptB0ZijBDGWf1eruyak6UKDZXFu9FY553Jc2BG49z3Y+JNYj1N7yanMiBG2fP0OfdEHHDXMzzf
ikFXjwzAl1gFsEWcUyvN8LgVe0/OMfIuSE4XXYs+3/QOn1+UbhnaXdeEmzMQazICmvbd1kp2LaUI
4TYdPUVER/97btNSM5TNqn1YnAyzoS8NL09RqINZ1yXuG6Zn10PURY+eG5F4XAhuknkyQ0DQ5Bnm
ZifmGsalYlilkKjshZGBzf/IlFa8OwqvXlIexbjhEZyCAppBLbSYuddNURp7T2GUItH9TTkEyvuB
PJPqyTm+yeND6Alb/DRA1oX1Y+5+MhLQcub+C/dLZIc79fhlxy8BNNN7HoaDuC5yICZChHLIu5OU
69pQ/JU+oc04VrwNaRqN5W4ND6rCKD5LUPQmsBCdCm3Bo1s8pBgo7kQLYxbjgm3XPUdujX0BTKlh
m7FQNZmdOMQWpwI2QdINXYU+dEz6pCOrGg9D1EWu7O2EU9HeBLQvCDoHj6IdTq2yzEUEPAU2tUFV
UH+rA6MFK+RE7j4qsncKShjuey5dkH/PC9ROenTqMbqiLX/TWOEtZRpnI1+sctNwDH6O+/+rubrr
VNx6HRYOCBRYil25diWURIj6Cbbm2gvHrYn2vo+EAUVCfvSaSWv2pgpKPP3gUzzQRvfEXpgSCSim
oShMZ070LDp3n3KCcZqS2EDD4xFOvyWdqEXeLtZeCmd8fQIDCNROqCjUR51rM22+MjaFQ4+0F4Bv
9WWQccl3sR8XSsKCyv90SSLBxXuSiW1L4D1+WwxaQK2J2/fyaQTbhBdMfLFWC6/HoBICZDBCK0u7
hJt7Vaeahb2wDvTa2ZZxBo27NtGxIZpLOhVnOyDoT5bzxdUdb/Y0OuXlUnf47h3c4fLnkofkxtn1
wuTAXSeAzmC0wmv+2Ld+Y8++PYDnvG4B99bY3fK4p+b3cln0OgACMvaRN6BJ34brO3DVEG7eb1Zx
JfqfRUmj5nVgiNWoJ2miOFWodl3m62yVJGM+LpKUT7bZADHqlBxISDxz79zDeRXzp0DAuO8Fqrys
KS4e8hAEHl5/bS7MG8z1vf4U2DHVXcL154yNQ3LlGY7UQ+ZrrujL78fm+JKc/yPqx0ng77Bxy0Fi
zNZfi492DdWhABDo5x/SfcaCbBVRk1jC3RC8GyoRdX1FlkmoEV6Dtp0NAManNdVZW2tJ4A2ABnB5
Vg1zQVF4B8/AuuNzKop8YMTX3I/t8pB8fPu7xTIckU09+Rp4DSJxw/C5Kfi7/2WqNIPbBnbxpkyf
REm3pQnUM8rvmeAVRU1BatwSlF3fnxtdn0tOS1rXKvqvAKTu6yHP+0im/Hm7qXx4VD9nDeBkIxBQ
YxcD9Iz6J2ojNjVADmpxgi8VDKa6xLHxqN9V7q/NZ6CJMxrYxaNk0xThXZgXgsjgKQyBIOISvr4K
YMPdr7R2tf3PRqxqHOKnDwwNrhv8QNdwjtV6AhOpY/PB0VL/zZ26yL4JzWGwpVtrOidiDUNs0E+D
KjYzOYXNVLPQ2z0SRQp46MYF4r/Mplp9HyNfYlI1lwNV3e6D4SyL5h1W63zetkYSRd9g3U+gid7i
b50d0ZZe7et6nemBRZTYb7LDv71cSudNbPpNkZ+Vr49WEwk53huES4mwRE+8yaY6WIJU+WLRu8Z9
DYKg1U0YzzFDeADIXhByPSV0tPEToOszZ0wDSsggFjKne7MPJGrHgQdT0VXdlZdGLAkgddHI7Wm1
5nOb8jsw2osq0Gkmjvl7rbdfzd5wZ82fiQa8iK5ieOJrr0+USU7X8qu0WJ1Qv1OSePkzlv4fBHvY
YvScjjZueOu7Z25jji2IlQSNLhtPo9FA42mmY+NElqNDmQ3LNV/HHMBOHMUS5GJFbOe3UqDgtU46
T0M08VkoN2SOBaTUBRmwdNEBAto19T5C+zcxyHMFlAjFnEAeddWyh74CCBbKvhARJZma6pY8WsLe
dQd8Re53/9HTJeAQfWnlvuMv+1AY0sqcvCULgSlEswDBgUHK6AhKJJeGk/oJw5Emw5kn7cZGnyxh
XV3d1ZujyqHWZO9954h3KclipAA3AMt8S4LZwOcb1g7xU5Xvn0f3o7OzxsTbs85skeAGVO0do4vP
ouRMFiLnZFqMb2MW+9b10RPUuh+5pd8m6h4eQZS37QQnrE2Z7eizOGFs1htUF6ikfiJesUTiZ2dU
BTh2VyyjpGVYu2Jhfeav5x1pa3bHuN+/mafiGJPYbflv2N/wP2Spg0pnwjCBQdEEcxGCMwjPZTh5
57A3UNKQwlNncBMIrmOHsGepx53tn6fyLY3JfbV6awaXkH9MTedBXXvyIRc462rWcZyj1cIc0W5o
8bGeI0YKWQIaFL3NtvcQBrOXWpNZSQ7shh6c490XOxh3te+CB2fXyaryX8ueXg/M5sdAAy/i/DW0
4Om3qdDXpOlB+Ae4UU/dYEJE3nEOgIN1o6gn6ghlqoBFrYWsf2KDy8E91uQqdi/sQ9N5RgK3fbqu
hiOOQbKdTeDdWNG0qZ0CXtnx2PFFwXhZgzPaSiT08SjRdF7km5hDx5wT4WlKgvvZlQzd/nPHM2c6
t9TMi7UVlgfd41k5y5gNr9FUVN5SD8SfKzMXDnE4G0aI0pkBbr0qAURCp2rCKrRhNtnfdKt6s1MI
SaC8ZYuTK4V0kCko22R9joYlKsRAKK/Y9or+3jAOoFATxr174xwIAp+NhzhL2Zfk0spQj7oolunf
inZ0WPYhl/Frz4ygfWjkGhHOmXkBHkmcs/Ek8Nr6oiwDyMDepsdxkX/ewsWFgfgPRqmQw6xk/PVx
s+LtRrR+hmfWVPMJ+jVm/kRLWJIbEm5/BsAjUqxfKblnE6GcUS3TCT97s36fZMp1hjM8vWSCinES
ToP7LQQgQMmujpGgVFfXSZD8uwREZv+00ZvjpXme78gbFVBn79zHxZ6SLcTIKsTvaxFDjg7vLFAe
o3pwlwSxiQXR5KiwuO0NYGrO8n6V9sji8oNFPptzHa7H1benunLMJ6kLRqh+eS99chPzXrcbQiI3
lVhOLtX3j9/CiA/cuo+GpfXQioQB7e2HRV6HQWPiW/fAtRpJYrr7GzOMnHSLOLoYMqZbMdos5rIk
N2ukg73qY1z+Y1a9aJ/x2kEsppblbryySARoy3aGsc13ffPQR2wZdMt5VsY/5hx4nOWOtiWVBzVv
Gxw8nrQD7ZgDmAeHvDHp3QT8o3CZ6wS7llPxjCUG+jdTrzuFxUqexReVqcpm1mX51PVH68+eVt0u
B6gWz360kjZUGMW8WxTLsaq4h2swp4eOPv9L0MOL+iUYvrdzzzy3u6ZDc4aDak0TUNgkhNG5qIN/
MpJUU2sRIwRtMAz03Hpe4DNQM6CO2FK/vgYu1S/7oRdgnKX4cwvJnjapf9/M/7sRA29tfcQObJKJ
MAO48whnAbLJeFOYwHnAEsXTnQkU5AzEHv9a8t8iarxnukEXoIGig8g3AClQKQ6H8RvzEwzQlP0P
66SDKjzC0jToAzCmkV4uvELyDYCnJa6hIQ7P7fg0H7ipfMVgIYThON+qkT2QsJGMq7QQzE0OhoxX
wQeDpJHXuZAYgy03RtPrZwBG+S0Fbr3TU+Rs9fHUlqw7CGrA0T975AMKKL8KP6QxXJOLpPiPqRcY
DIW5rDHF6sZavTl26B7X70duX3ZwQ2Qst+Inj53B8PHZmLq9g9YyJdzKAFHZwn5+lGEuQySkASSc
t1NNnH6s/e9+/OdtpK+4r4RgXTBsPgVt9HpYwyoKQj94VaguB2tvkDAZYwlU6/hqavEZgXUFnXbz
jMQeAF/RUgTvAPhWJMwfMmVHGbf9rumOaY7DfQOH9D7z9uboDvVURimT/ZRHSpf5A2LCx5/+Hz78
Qe00GyBdmcJIT4jxAznJbCmknS4158YYwnzmHkkPhQ3QeX5q93fMT4tnp33kJYN/DGehP8fqr2OF
O6KYiWVxSPhvIzmlrTpLPLhH39HpU6G8u4EBFsYZ637hBwtEpOK25m59JQiJIUDkddYNviv/iw4f
9gm6wgfl2ge+RxZk2LQe+pAZaTFAkwb4u9WZPqdbiSKuaXw66Ke82qIfkQIVk+VeKaXbOvWfyz1c
G0JB5htxY7qLKP/Iu4i3zu77WznQFnPSy4/0M3um9l505T2b0A3/o4Y7wxCW/Xb1EMmyXuUjFJ34
bj1xMmwPs99m+8Jx80UDvkLADa5g9VmYZBgSaGnR0Qa3wWZy2DT2913p1mphxeR8yQh/oxnQB/V6
AF6DxuHMNmPtJykptFG4LFGiJ8Tz1sAHUBdYQRjlcUggouu+RbZwgQxgYS+/k68R59GPbFNTEfAu
18aiKoDh1EuEqCbths9dDdhZOEKB7yof/94WobGbOuPFS4Tyk5/YT97wsmkWehjkxaCxoBPZpC+b
r0hI1pyXC23e2TubbywvutKBg6g4PXAry5/CYb5dSS0huNXefXf1+4txv82V5tphWqWozrziiCik
JnMhCeKIJxPp27NDV1ZURMBG6WGDDVIeamFi/lmEv+uscXUU2whWY6f1/ET3mkKqYoUfsf/If6k2
xwR/Saa2C4dLgsIl8Wbfi8iyYS99FGhJliLIxMGx1jjVAe/lgCce+4RUaZvbHTlAOXVkJvDiDXiL
9ffsxSp2pN5Db4CARsWr64QQobp5V+6kQzF8jL+VMFysy0IeCGNwS74fnP+cRpuctSdHUn9d95yv
F716sihG0hojzaiDkjeFvsm02J1589EXc9HvOGddr6Nxvb07pchuu00Mzb9C1K4tyAaZ27AQAoX0
SBp4Wtks0IzWMp0RVaN7HiiRjc3nRh4NfSp7XvpOGxRguLlFx6n4cZxhIwPPxN+AZ6MTiX/5pXcG
qrgIPSRhWOqSl3/P0/b+dBkc+CrgbWTsNoUM6fIsm5oN6Du34WGKgSTHNN30fhyQqulGW2fUT3v6
QnX/enZl3HzpG4BH/qrXK/yG73FNSM/beoDwD/SmYRI8hv03nTMPE0OyHwF936HUeuvbpbQ+EsPt
ThS3XPd+nEH8PuPiVAraT/3MAyKX1lNxxtUYgvECp4EJbC6XRsNn95TKnFtC1WbwQ8bJsCeqMiIf
ORVlkMlxKf+9Q2HP8gVbpA1Q8vo91VGLkvfVKIhOxVkveZKrRRlyef6TXg9j9KLVF6SeCIld3NjX
CjHBOk6AWCeHEAYmp3OqfnYTkO12CFSKs60A+jOZMfw7KFzw3p3cCjQG4wYuK04RgTYcs/4A4zfR
f7/kzmSYAKAtIsre9DDQA3Zx9JJPJjhX8W0oCuIM02eyzVchFD81rViabVmxkMTsoJ6VXgPoulCt
/JZB+U4+A8+Xi0X2J7Ez5h9j8GxZGCJ2UcMcHuCh2lo98zPXvT6qEa8Wx+5eVfmCWuds5M6Wi4i9
sSR38zVLHuAJ/tpRoT4N3X821/RrYhHknS4zjyY3XHpQ4odtgGbFRCtl30eU7j6XCdyupitmxt1i
TS6K2LAO4dF/ZvG1D09K8qq+k7JqQQF2LUJK8n4LUKANEuTb0VeyMS4hBqlJiFHviypTsm4d86N7
MGfCanSezeP7uGFxKqFIz3EQveJu+fDnlA5ny9+/PV/VjOjNGEfWD4x5zrO85++ddGpMGCapie6z
qE3EX9py2XVVUIXI2z3OCaq+5S2mh2qknKTxmVnMKPgtNHdUugEj5QGSg1fPb99WSqYXlCW6TdzF
raKtQbKvU5agNk2DDGlnvDnrClad/ZT8yBPk+AiScZUBA9QTrQv/Hza2I16E4wEoDfbCetCfaLZN
DfKEvWXNBtzPWoQbYIj9Gl1V9CgJi/GJfQ2e8i/fLMPzlJLwTkkjXJHDWqp3w8llev4/ZB3AgcZC
kdcZ35V4ppJ9SzBUDS+mPDbsJvXyaNKDSzmnxjwGO/B2y5fEQtVO4oS1m85/Mmqn9n7H4SzoYLlA
TPpuE9FdXgJb3eV2xtyyVQppZEtqSVqPcSi4G5yuAlEHtjqFV1/X4V5gHz6mwtHRHztHGsTHUyE2
FSQJyvtetYe9Qmarp2Xx4Yz4VeQKgqyv/TSaWtO6X8vGgb3BC+vOv7zuBZ2bXlE7sPkUywkNxvZm
CQNouzP4LGGDtbT7jhTXltuhf1OhWtzPXbimGk2OgzTz2pujJ1gWbJvJs2h0Xa4rfatnDVwa+hO0
1veg6V6uwGHU0YulKPGN5v8s6XsjHEBgRD+Dbj9YbKBhq1vP85SIBgLLgYUWIvqVfrHyLFItiGAs
6V/MD6JTnaNjmQYsRCozMe8Ci8ZCIHOr7ire2CIiO4uMvz/xulhKQ4KKb7GvhbFENXXcAzttaTsC
/4TtvoftW+Hdk6trzsEqDnP5+l0tJ4Axw0gRkm6qGwd7DmFF7xIHXbCokHsFN3G1a1yk4LUlPtCC
h5sqUFqnhEZunPuG+w5F2u7xhaKbjLOHjKM8mPLgPjnmDMT8sRkOj65KgZuZFHKE/KCT2tywCmmp
mKuYHz7tUtDDX9/MNqHRF3lSGNDpGO1qm2Y3XP/9J7s0nnd9uAYnPryeYYGWiHf/1LA+kqn2zbgs
WkBXZgXzBh3k9NVJVKABtpkXPt5jglYrwYRYHbSioa31OoFp+vvxyJAz+7K3XNovIcLnfV+ZZJk3
ReqDKVlHWxGdoA3pWQ88LTiYM6c5T8LbzURja5/aeJ+mudto6Ps2GQDuuJmun2IMEOKlPaN/M6rx
KaIm+/m3NLimeDROe8siW2fyt8mUkh6WMKlvvgWb/+IqBDS6sqMckNH0laQ42GK2Kt+2RfTlMwYp
a0DaeJ5gRNUUktv2p/EWFm3IkEgm76tk36mYKM+JL+lgNyrqTjdlg1cMrqlAmfHP4X6g0wyo7WNK
I5xHKXaCkQ43EBSaFyDBdFtyln101VCjG/ZMZLH6l9YICv9Dze1Oyyg6MnjskOwALNSr3iHIhom4
x/2ETgwBv4izhkiNcp35KSGPJjpUc3PaiIOuTcewBZXxS1/cXWFO2XoMkTpqg6QPMFMRTaxSjVIb
vhp6ViJb9SNDTSa/tERUrhCZQMv8EzbMigFu9uc8h0Q/aZNGpir6FySTEbkC21xkL6WIa8tdJ2uS
7TdXbVLiJo9GE8KQ2SW+ZCHkGYmoxiEMt5lbgu207h4F522D0eQz1RbhSYqygh0EaKcrz68JtZ/9
/p4d0zyvTAUN9ma/8wKU9kZeAI46OYftk9cj9KWVy8yWFZI7w9EbyyCe1fsgALrIEX3nORVidT3b
swyRjJhn/iXuTg2J0C98o6LgwEDsfNDfReVvU7fwnS+unv1AUJCdMzx5QZgn+KJYW/o2seYVaKMX
DYedWkEXFUAbi9x+6e9w4De898HhNGiQHCoTo/MLYAhBNCH3vGRetDGi6vtkFT98kSCFqPknhzSd
onqicCiWgbqb0MygipiW/nsqJUcQdZWrDa4ExtHjKg1483sqynQ2Defy5ZWIDo7rxBpvv0272OBD
KpTMF629W77o9paaxc4vLm9fYqfhvRBw819nid14iWpmFSIgg257aLvFFC1uttFNpvc2E1F9JKV1
kr05yJNeUnfK18HAXd6kuabbZdpYIXwjDJW++lSXW2KZFRPzHLhi/37k4BWCkbXl
`protect end_protected

