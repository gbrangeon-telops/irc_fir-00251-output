

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
p7Rd+JJS6BPhm3C8uEMSjtB2IOpOZImN8ABL10O7dB2/wknTrPPVnggIUugEe0Un6rsHScVa0yw8
WbsjeU4skQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
bancDuzOXzE/C1Vj5QpW3wyih2C6ymZ1vv70urQ985WeT2kXc7KQyN00fbod+1ycgrcEzdZs+OxF
/cQLUqqV1PAWyHyEqXlxABFUHjs/nxBl/f/B9V0jlBhAzKCCHBVtW+DFv8KpHE75Z2lg+r4JTjg7
zQiXYHxUisemJqUJdhA=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
rZMEEzwWFXOuo5snJgtfZx9Urf7eZRBCxLhuSc3DgaT16zNB/FC6Qo2PLk9pQbhTwkt+6VFrAqaq
rIuJ+6NqrQaj6tzRnuILLQxRIcZaZnlaNGPM0QELT1/pgSpbDRVs/w+jfcFf6hDgLWdb7+lF2lZt
EzdkUS2z3RzGxMw0dEl0kPzX4BrObwXWpUb1u4DD6JMZb6O50zBS5jLIs04xzSPqxA3PuLRWpuc8
zAMmWK1PCPqsF6JmUA+ToDlUTA4DP+Qb/r/OItKXADHbpGUiJXq85NgUc8TOMYazRmcSDk09joNa
rvnt13K7ONnKnXu7DU1cLEZpB6zC/Q33/JmxrA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
fSUvPGwGSOzh5U1OjbBgxWaXchd+ErSm3+d+gvsNPzEzvrhBDlsbz7cjXesFumQgP32hemPRlsUr
lFspe8TkimNAMoMtRIt9Rpr9MJxdvSAJ2AckK92TaQKYGICYWnAAwRZdM4hFhKQynq8onwVPOItS
8G6qhIBnq17qx8rO48o=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
MVMseSXR8Gidb6hUpBeQo+a3Ho0qfbo2cQ4XmaaPwOf5p+bpngyRNVgFStTGlS9V1Gq9sxZR8m59
KVYbqvyTG1F7VywlVWjcCzm53JiHqc7770pyh1TFlHFmlBkxaKOZI17/BbAJVPtrgC1AFUgqJIKl
KWFzGNfBnaqYhwSBpkZVKTp2N/RCKh6/dORV7jPLmH1kXSt5iI647oKA/xzmV2IPvCjRau9wfIMP
3BcMw9SliL4YOeA2gPuyEVJdJ+sinBGqyYpGCshGE4syCgACrJDHcCC8bST8+Ee2RwROkSw85PvD
RmNqdRJR8yBkuN8MggDeHwsPe2oFAGN33DaQEA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 56304)
`protect data_block
k1hnGr7++S/Z4MdL+7MS9p6AvhJSQgFyWF1k7uP+xT0Xl7wwYr/WVrcllDOu7oka6BnHckh+5trk
muZ30ihOa/3yGVx9sTmiyvYRHVPEvQJsUQdPaFhXDKfjvU3VNkwM929P6jKtXVkLHu0hhb7E+n5l
msIvfgLFWwwJAT6md72ZTJ5wtO5/6o7zf7BuXhJ4lfXkDqeJ3bz53yUl1fkH/P0S6V2XPU/V+IKY
ADhISNuwuEThOUitF1e5V/GQZiZKVMyXPfIKbDCjgcqAw2ORZCU/vOoktNKYzbqJx3xVycz3ufd+
4pQKLaOvIT8uGb1zUdhQu8hxRVB/DobD8NC7Qu5GzvMAvxDVlgXAq51Y9SJtRgxbzEC4eWILl0mb
QFy/4MWvxTuuWMfPR9R+NRuPP1tPv6fvsVmBypBxWzXyMRqDLCdUqqAe07ZcPwWm8gO8TJzxW5dL
s5iYFozitxIqc+O1sJI1UWxCOkJr4NlKlDZ0bE/is04WyryoUe/TDYTZUuzhMURPpsuECXmqQuck
Ryb44B6Y3ZAeyqOPTt0WP0MgGH6OC3GDP65LyCwz2WKnCSA9f3zUGvlY0Lct4hVwfylA+ApTFYqv
3IGB4gVZNzTN1D5sSN4WHP1ltqWwCbsuPJaURMkPxGYu6wEF6ovB+zEFL8bEpfYZKB0v3+gSX66z
zqO08zXpAqDsXwmyHRSzPzyADXdZIkImfo8wJWDIB7gzkJRcn+pndVmmPY+ezlzz6Sp9Rn2ROhOv
d/jA+70kgQ1V6avfGbI0ARXjwrrwAgZp0qfoBpb1U9TEqTKAWGvcKLt7YZ3UyT/RgIAwvXhT7W98
tacgmhUFj1t/xxdE5P7RWV5RsDA2DrJP28aZwa69qr2OpTxJTaVoPuOiNCbibAnWF9mOr9MWhcWG
uLfGOaRp/8fvRh48IqQc49b0y2MxdVXyyssrPm6bmYFmKADf82e6MFCeLr3DiM+bObb38NYcHz9N
OMXwkpZ/D+1oFAB/1+TITIsW//jIVNodgFAkl7Xb50zOrhC1VUOjua8gcWDho70v/Vue2sdHzKuO
1cwV9vs7X27HNESIIiGjJYh7xsMRVlmUe+NtLKFdXzbByXyyTy3nn++5zvIfedZmK5tFWMk3U9XR
KudLgEqkCjVvHr8JDjOEwKRXNN67FYTIqyXD83HW/KuHBCi5CBWbfu+xqghGiupAKAxgn4bnYUxo
XQTfITM0V7wm8yvmTIGe2VeqtPRHF3IVJet9Fw8gGX1oY7I2ehhQkm1TNnTd3mog/vx0GKxAgQJe
NIbDQl5yc37EyuxCHAiR8/PWH0oVm26WdeuiTSadWFSj64jHBlh7408H70hJEOFLTxUBI1QDiUcj
YPTL6rE7xT0OI4ygX7+TSrjSJ3piUn1wVgyPvI7uAvrFB/XxYy72FjD+6FP/bKGHacarA7AxNJl0
UZcGjBudrZxF6SKOaNGXqbaAY+9TaYWuaP1gnssjxYcRrmm9DnKqaYWdDAGzkJFhToCKkLyFYE2I
3z1bKMAPTCBR7fPAEd8VNYNrQfQeW0LoiMiqhQ20/0WCFA/gckz38AitoR8bFfMsLbqCWAlgqW6A
3sknCmlxkON8d0yoMffmKkWdZTsoSz4PcYFiztY6otXhPKQQQKJXT6Qrqnu/pbhVZ3HynwdaUUv/
+HcWsIKETza/1arTDoVUFJARFb3sAQt+VvC4RkXpzQMAkEyhJRz4KTVwAoUvqcy+DRAMpr/8074m
Dox0txraPcM5aGxMXWkUOTB80Pga2UXJVLl+ar7Ll2ZNOO9+2UrAmW7dsr7REXV38g6WPjThqkt2
Y/fJFNlrRKUj6Zyq4kaJTmuTiPwXEqLKjXdGYeAXlqzpv+IFSnegcA9tyyzYlhNiEiDZE6Gt4rJB
tbllpRISirW4rerqXFyhfpz2zDQREgKjbdozQk6BUCsdc9xr5ycbAWPblXx2pdPKxm+p0dMIjI72
DEMk7aAsZu1HNN8FjUtPt3fqLO2YJHG/W8JZeapQOJkFAiHv27fAWMl+nkzjIB/rOQh69a1BynVT
dFTmfUpjRN6lqmJIzCmPmFP/KM9jEIEpqJepiyH6u0Wbr5OOZUDg2QV5L9OwlK4ZC/Y/z+o8WQwp
t9bFlK8DMhorTB8czqMMWu0+SY+Jctfn7+4b7yl0i8zrGOp02kEdTr4KPTJiqbUWmFwK/vRMLwd1
Vx4LnN/is0XxXzbjmKvk/oaAV/wPozj8kD9FvE5O625dPrB3TruBEAPb96XRZfuP4dszfaJGkkPz
0rtCkLxeuJRMtCflw47aER+MhBF6PFt5ari3o0/YbVsDy7a034EVs6njvvxhBN5lBQHyLH0ND1RO
cPyr15AbXZHAAmoovISJxARhu9rJ1fgrYSoxubPprECMv3Eze++Sqy7Ooc3on/1JX9OMBxKi/4B7
ewVQ7UjYlROHLOpNxJQufpv5a2AAOkIp3X0SJedGragVBV9r2oC2OdjD1ThpQ6HZ6taDvRdYV1/n
mMMJyxk2YQghMq1yOV3lA6pcyhqeW75QGellOVcjemmHZcRnLy1JmmXS6mFn1Mll+fdAsFP97/G3
t2wdUJ2uitdaW8XHMTmt2e6H44WfUPgjZrLqZHfqqF2UJCVlzsRSZXZ5qXOPRC3sk5zHb2tD1qn2
cvmpSpEPvkZ0/U9BIehiXYxQh8wL4pDYTHEfYxEpV95g8aYTgTLWSj0iTxOGhxUbCXf08hBVSJAg
YJ/pU9ZY2DdAmLPaptb9h47tb24fpZ2K/ebmoLOwEq3uzsCKEnk6CJq82/odKLEmBYX/FYbKgqik
JxYFNxZkw3Y6BRhocdQg043WhvK0kQo+I7Vh+fPvp6jjcXxCLxVKx3CKTgfCwhfpjjFTSCXAKLmZ
uFJDmxPso84DDz1i9KknanQKCIrLsEPFl5TJOyPQ6OfznZcy616o9ynjbQA1nNZekQRwn2cJqve3
Em0G/J01xCk7steroECDXXHWfF1zV1uzZrsFV3EE4ZUQIkS/pTlVXBEfglpKyiCzpd7mdWdz06tG
Y7S5/jv/EZ+6TdgakADr5shkCESndgggyn7JgoPOSyVWMhbBR3RW3RSWFDmzodb02aGvtU7bM+p2
CNolNmHoJETEVQwcKTUi16giEDGWPhu6bf8F1lhUDXccO0jEOef4sJAweBkuspUNUNnFSVo3bOyT
ocFn9/UAWiCF0tZ+vGJkSWxxbOaPgJ84RJh62Dr+EJPo/gC+bOPRqidFFXY6m3VXXLOcK+dCUZYY
Jd6HMS5XCmljCCFsA7eilr26D7Aq0oDM3LXzkJypudxhvrcjXIZ/MZ8t4XR5DwaNYjrBo7/4lsrW
OmTB/0LJ12bcMGeHR779sjIA5QBu4w0bJTr3Hq+kd2gTIF1Bc3wjy7BDDeE+cXW71MD2UaPNMMzH
UTe2X2/zzzJpIMkDsHPUmvmJyIGcpnArlrf5E8ipatfvY2Tf3jY0GSV3IFcva0M8+5Kt4Xy6x4Z+
mgsaxvBQA2+GGVVMzVKivOOH7KWe0It0TfOohTWojZD4Yttr/x12K1tDeB3iNSpjNmOLJrRK+77+
CEkSw6zEP0Way9ih0DI+LRGD3vMKiAIeAX5VxLr5OI0IcjDX4k85kca/1XDj/yqWl3bUzLVTy95M
zEGLf89wolweKiK9zInbFNgwdrn5ZAh3kJJT88ALaEDXU4Q7+ASShDgu59aFTeJqGeib0MZbPYZt
MiWxZ4VTYMxWcIfIaL6w0DO5Fus/YqtTtlYKX0ZRk8r8zZRWWGyCA3qE56wK7nM2cUpNcHvZg3bS
no6fIMU8fCIMrDq97HbfoTegLGM4urZi/GbmEpx/13DzMlcVaY/YcFeiqonvibIbfUdpdXRryEsR
u3g8HE+NiXdFyg9er77VnnmPJQ61k+yLNv9Odt+hliTrVuAImPd5ToP8nt3hfarzQyHejOm9MT/e
EPbDdKEXMG1vlwvYachAC9J3L39GuNGr/b6D8kzVTdupq3dufU5fswJTJn6CUSQGAT2z61VrbjyX
/1tZp5OaS2GM9du9KRRBOZHdblPExBddFwQnGBRO/mihlveyVGbhgdR8allxQ8DQA91hZnkpCt95
bOoyReDPy2jZT7VblgtlT4T1+E2c6TUct6xeF6oHXlQBMeAbK4E7ZKrOEWF4xcdvXGviZTCGJ8Ae
sqhTqaimIGkePJ3aKlLHZtYimUXAkJAXOY+Nd4Ox4DA9oyqwDkuxzuoFtM/MivPT6IA9ZcZh2hAQ
p2O0+hIapJ5gyLQrzQwbTN2DptkFLQDScfOlrQk9XjaXeCs4jAyqGQL8BXbb4HWqSNttGovFCIBv
Grdz9Mn5tiHjNv7LivM/HGdsopu0Z1BaNze9YQVz97yTh+PFdhxMys6HGUU1KBd7CEbc7mH0ZtBT
m/nQl5dXT/B9AvjLGHEZhHHSEYUyD4PK/ZwDnZzmbBsK6U0b+7GGEBfK8Qcm3NcERYByVMyabdMF
7kgDinM9cEXlZBbKpIaDWwr7N2pYglMS7LXqGBQpKIh5cH7lj+EZotEEFoDykmummSr84nK+5jCb
JFyN3namBzCz/y7B8MiujIp18HIVJ7M/xk9HKxbXljlXBHI6TxL6uaZBD9WTjVdmolhmcsqdFvG+
UNwnv3Z5H5PUiS7W9eHYsCTrQeQgQLGPElVmbzTGShZMvRjbIQfAI2VGpr8hRWq9yCTqV0vWebd/
epgEUhY3CAYdxBn1IF8RBG+8DTbDPydWxqsdINlBFDuMoGM56ccr5zHTNy5A8nqNtcpO7e3Y2gxa
WEcZsVdCpp47kh7hstVyVRsgp33rC1Qfc1wTORwzph6WWvKjAcC/gsCpu3VL0FUZVQRDwqFQlhPS
DxBQwLKiN52CGTgtTvEjesZBfMVw9cR6cHCURf5m9nENroNElHwgdR9AKGs3D0M05BEIYWwi6P/m
MxOpPDKWLlK01RAuxYYfTABEP/t1VLvK7x704tI5WZZNbcAO51LyvupKKUdOder5N37kQ+Fw+TqT
eEkNJeLF0KE46uIMfYjldFuESF719fXyZI25gu7mzip6Qg/WwhZSOmNySHHRKuZhfvTc/UBXBjvu
X6cfUiW/GRKLy4VW1TQiAQF+/ypJNB76cGq//434pYPobwFTGQ3YspV1hF+Oy0aOU8vm2TTbmftg
gG9Wh9AZMBSdnD8oWO3RbHaityBiQaMhS890gpLXmfHJ4xpQI1TYhqMQbKjFp7AF/DfJIHfIwv1G
ptvk3B447EQf1i+E304BD28N91mJxCVJk1JKdDDuBREVQ3GUyo5+TDgduu5egiPz4a/3lu94Z3+l
pXEqCcJWHyfVXFMBn4XK01Bbrap26lpuXcMHVjhhBNhmt2Cta0Cq5yB004A28ic+3Uia8wHb+FqT
UnPhhxWTnIhoXYpuNNIpbuVmCPkkmgaJkZKGV3nJ+oA2Hij/NQTGY4h2aY9zZWr+nMqi8n2ab2Vi
cA9CzLb1WOcy/0W7vRwMUo41gj3r72GNr+dGzXN1MUd5fV74h46K+JD9UYg98v6itBManhcmU49X
IcF7UoWAiC36aWj6XgCS+uFZ7eiH4lWq/WkEznIoTq5zEG2W+HIdHAMcZNXdAIhZ+Sf+yeR3Wk5p
Gs2iADBFCGwtJZNmRc52ktBDi5epz0WIPtLDT3qjCSG4ESBxZHUS0ZvZ+RrMa48hGxWjV8ktQhM6
hkjWTtQfSTDwZvZmtAQs0XSsvs7fCOzeCo1jsyOL0dohtJEsaDcjcnx9u/8/E4v6QZF3JTrDZXM8
XrPvcMf7dcXz9+Lyls4tl91SDjtPy/0Jc6cR6nQqMEEDjxZBbku4Q4nNKTxTzvA7Z+ZXQnleWnbh
JoV0Iz8tQ4JnnEbCMVkUJLSNBxficZ0fyQEwBs0zwuxcQuo9HpNj/sH0gitn/8FiA2KniAF++63e
Y52/r3u+DsUrDUiMxFw4zkMbpaeq8L2pTNPG1hXTjq9t7g2PDG7qvJD19wOzVswRtoHglW0ihXR5
Rj2crr/mQRTRRbpZ88Xw9yFfqUfPymycmITjLD9uBPVivyHlvJIB6EjMWQItzjzVP9Ta1n6IkrFp
f9mceiEdD10Eiu+T33p1fCmliwQBYYcD0dWAjv0tRK+AjLoStl2YN0phjb8hGArtsUB9l9hf9gea
CmFRkx2/OzC3NS/3Xm/v9h+q0U49NCG6/9e82uCqDfFsAkwcdXOARy4srIs/C9PHxuXB5idk3Djw
yn2r24Wy5XdC3+5Vs8KGb8uVW/WvsLtjQmGHIH0qaEsLY52dN1qwW0DE1C61YnCy6g1U3oaUrLx4
w2WHdNPPKKm0aTK++kLntSLAZZjnqCw3QIHRArlXXJ7bo4YzMcLkEPF54VEyMsZrXeYNeYU2Y7ej
TbDqFn2MBpH8f00oOuo80rz8jpgxRXX1BZO+j+D29tvseh7J5LFgmfd2ar0drNGq+YJ8gNTlKQss
zwnb67mjuxpZyikVeQk+doCVI8Rv5Q1scXVj/OSx5ABWcTnP/7ndcinzx0bc1dS7iA4dQJkGRbfG
42K89XggHagCYnt40VnlqO2fqwg6LUXGym5MVaLfeK9b9bqHehtVzmwj0pHGBpfkT2UNT2H0c+P9
5JcZxHRyIHGRn2p70uBjHse325dvfgm6x85SgCyBXzZANKwifjkyRi1hesCft14OeG2f7OJX2dVb
cYs5VLtLU3rg4MnHQfSK42Ziefde85jNHP9c1XseCajBvAULKq6k+C45qs0hdZIlEKXheND004on
ETvgFaHyqVvSeQnbTCgDJHfcddTgKYnsLJNy0XCSAcDtBteA2dN3BijTg9yFvQvih2fiuumBgGBs
AorSQ3da+RCHOXSr1IsGn0/W84+3dvba+3qGYYNawFGkeLOf3bOqM1BUilZfdKYNgup2TVq93Dl+
8b3ozzStplpEhGiz4+TGVteEX60XMKuyu9osIRbHuahH02VZ3PCWbj7/dbTfgd73EwKaflyOYj6s
nVe0IrV0Z7SExZdxz2ma9Ow3hhg8d74YTJ9/xK1rZtwSVGcrNXs3p45FxYSWOE+jwcD65BHSm+Nu
+OVRUh3hsHzhD7ynwaQp0JEY2vjujk5wnoJx2gWqcQ58n5N2cfo0Louys0RsNMVCYYGC2FnNm8tL
scS7aAHzBFNLdPZ4u6cUiIwVhDq9MYPJQHIY9nawHCEaFW+5awtWbeLmdRLHW9Uq0IxHqK0VmSMr
k1AxHD1vhk/DQxz+xb4+1vuEplSTpGDkmyl7u9iKXZzfn3WJ9l5BsQ8AUWia59CK7itlHdnd04gS
HAynFgF1GRpl92oZoB5M9cyq9+ygaWWOpc5oI5om7DcpgDjl6MVYyWEZUSyXY3XZSWlhyvCvcCXw
8zUPrpt40NSkIjNh0FMNnj5Hb9qorGvn9j2I1QAwhMS9I3wgDTL+K/ALFVGiqf60GVUKTwuMWRdu
3y/ekGGZYlsWz92nsEHyLhcn/SNdaV0FqCpsFoKtWO5p0HVHD/2B8GmYtRTYp1+hQNRzXO1feR9d
ZvTfMlO3tvDPbl69Z45hja3lLy34eOyX4/i0IVDuSoYOQrHOjJW4Vdlz/xuqalv+xKhCy8qDZTUP
XMiBen0bxePT+7D/PsZhPLiHwjKEgA0ZrkPyeZfaYlMqN+SjTZxpHa5+g3pInXqPRpWqJOj4VlwC
4KZr2nV0l6ymCFZz73KfbzNf7I5w3dERHT67/Nl+VZifbLGJQtB0S3jIh8GT3SyVJppbWrTUr+FP
SiggAjDaAEEAqR6f6k3K3Zc1TdIiNTIiFZP7FIK9s8HDw8IWf13e6EMqidDxXqA8MzCaFQs+OnkC
dPPLpjGzGf5ZHNOSdCPLLIyICc6oBDajbPmKh7v3jDqwqasdjFQn3Dj3XLP1v6HumkcCyDgdv/wF
MWUX3oybQfnLe0dHJZohUkGo8DjMwY0pKQAztlcO/FuIDscUX24pOh+Mss5wEsfyWCZX6NmHAJbx
1twAxgVYu3ZGGAacFQHdX6+xLhn3RzA/uWoE3LaQmay5AifbiAMg6jIJZfI9KaSX5bgBfpMNhHST
GS+tLH947ERq/UIjnBWbNJeWDMhOQtDCmQcR2PHdWD5A4n/bmNCepKNDQza5orAVZG8tR04xX3Nk
YuAMTUESZSoqXLfmtkqb03ogPAZOEn6XqIrCFwbwzyLSDH4aIP4HTOWhaHIM9pOwENmCrx1kltsp
jGH9B+TpMQvCkfl7N4nNFp8hWJU6MjnOmnEP7NxjvWdc5B/OGOry03eQB/ZV73gnUkajOyA1GDMS
wlmHvUp3s2RktMrHitn255k7ruyMqVsOzGiGRNNL94wUzmFaz9tAUjwHkecPpui3CACxdF/P5QF4
1t3FwUvlhmMNNOz85nbEteC3/kQnWQD4DAeihYDQL5jfBmdsYMNxYkmPsEpe0szWG0EmSSvxDV9J
NIsd3RiuqxmHbrce2CpgMpyqGn8YM/C8l9CCYAwHlVUGvChrfY0V7TitgrrE/gED3Wndh/aHHFbi
w/JDMyupUNHQ6CIPdyqnxXq2Wtwiy9TWxzU4tbJeHII1rGGxr1SVngjuuVLvlBjWfNjIPxTBWGkB
FS+9evnH3uvoMqCQU+N3XJYmGVcHrgNeay201y7kqjNfuYegY/Kfp+qq7HCsZc96N5/2syjMxltX
omtFI0/uvSbYZE4LpElz3kR/0x/IBHCHFckyljJKlLwaeKYIav2G/ZnldqDCPOufL0c02Nd2AaT7
2qTZ1Pp4GbEozdL6tOuSGRIMCsA4ducc4cSOXqzm4iSrEq9uGkDaLa4A/MgD4ejnjKCAjNrK08t+
cbKnX4l+ICvXEEF6N2DC1eMOX02uh5ageXTgqSF1+1a5Bnn9TKHBXMcu/fMv+mpT+Z3uyhrY4H9m
aar7wqQ+kGcwRLWFArrCsYEzYGL/Eo8OhiEKjIEKJBaw6A8IDLRheBP+vKtIJ81ICAWVXVkoGpxF
3cjNg9EejuMcEEmUV3lsP6WZbpinJgD67tkjzb7lR9+NwW1JBsdfNOgUdTJ4UNMuXrfT/0wV/aDn
6pHOC1xfAKldCVf/gYbuRnjZ9CYW6VI/E3lN+DVMgvKVJbq8cUIHKbgoPqGdKAI6ZZtEdXYdJBRq
GeeyQfNPvsDjovEZ/+b+c/7sNKBiUZG/q1jqJ2dcX78QHl4waVbdx1O/R7NiCQ7fg9nX5lUfqDsw
scsOmY8lrPuyZ0kOW5qiZfUhno3P5zrl0aQ6D8bqd97L/U5lcfcqfv7u40UfAxTnDwTOtVdOP0R3
R6XMbCbpPOqRv6nPP9FELvbsqbynYeu04d20WYU6Mojm7yBx9diJudkrzDzu8qpLPG6lEyqypqOk
RpBTb7eG94HGQCFru7/ITnq+rET5v8p3Ulj2SRWKrt6+7u8+9HPGTevJMZKilz1tXinoubnm08bn
CLS6UVtWOyGEXF9t12l5WoHhyu7Bxu2X+epanJ+4NBz+sDgZQWc1AvkjiF+BlXXlkPCpEPJ3NJu/
c9+9+Hr7t5BnyCCdskRdinxNpMtrUOsiKrJsEtoT2n23DLKq6Sp6Z8glapWY8JRCqSoYtoXk1N63
0QgqFPMT4WL9bMgeKK6N76ouFmPLr+Vx1m7povL/5wxMH4qtkYtTNiheosE/WTcdV+zDCCN8T+n8
GXy3tNoQe024/BbtmAzr7zKrJ346pJhcD5YMZsNMxz+vi8u+opgHQbBP2+42MApUTh/TerHxULCa
ocIR/xK/kEDhAiQOR2+GmWvbNZqpWJHvpM/bJuhkBSjjtUzQbjfBqi+E6VFdpS/8C6Yrv7hUljjL
SN2sOGwUVcN8WhY8gTMfeWRKuu0y5SltP1Kg5KFUoGgJbmkAO7lAPEQttJNdmt7JC4TCHHwiMMG+
VM3VysORlWPon8bOCtV1mE+Gj0Q/cDEiQVdfjc/N0rCm7y6uD/JSEA5e2RGtlVRT5Q+D6JP2vwQs
qTAV1BWPs5u/tpFy9ObGIA0NObdJt/Q6DdYCeWCJNILgIfgaeRO/eYC4X7+Zy1psLMOjDYqDYght
L1lUByeQ5zpdPXtjyA9qaOGIm4zQue/2vBQFHh6Zc3dBanMM5qpJaXQBDIzZDFLkDOu4SDRqwWLa
naBOWEIenGm3Gu8xJ9VQPFqn4C8acr606SMd4BiG/Ulvkla+Cl94sargl+HgzeeWiHpGeHUeqRD7
ARG0JNRbJEPfuUFAURmZiV6GtwJo/cI+jr8SWlvC5viGaN/KqyMBdtyOawriHmDhmO7I7dBk8Xm/
nG1HaBJWgBUp9ZnLnyWBemJYiMiJPUzRO4NEoMW1o0dErzDhmjtdV2IWRVNWdKNzmH1kW5YZM+QQ
b0Jp46ww7CfHJQsMvWqeOpRiKxJ0HGgEmLDNNh7lFX6qE6ghCIeOvbMWD/ePxYKgxIcwCQ9IOLsx
74Lsot46uqqsTBfMj94ff/+nKSjTCcROBa/oZfQU5xnWm5DihV16vaPIRtFPnnuBa/DCWq9nLay/
/IvW4muA7adbd/sw4YAoiZ2zLRp6/5Ctso9H+apVlm0d/kuz15elNsJqPZj6Z7UMw+WQMiW/Rmul
ws6eJe0kNJVCQ9GgGiZ0uJj6Sqcdr5+URn5H2qFmvZ70T4C+ERsHqZbfbP/hCnpzeAAzd+GRfoTj
/3Xm2pSAq70TyO4XybJJYtNu/H29hTGLzMpjZPKVTRYHf9drBnWEeh0IR0Sh7AnrKeijfUP82qoT
zmQi65F9l7ulYX0O0Q1U/bzHpk6DtjJ/kIjPovywAlFwjC+kk45sWU4Hcs7ihWT7fy0NJLIgiLT7
P33/Tq66NZMRI26izkftx8T7aukdernEZWRbEBMe4l27HRX0QS/uEjqwF4t6V2tMU1EsP8ViGzH+
I0SpmDZMCq1+pE6f1pSZwL5Fm8plu9lAY8XiTHgcE2DhEaQgmi08WkQQ6hmPaNwjtyGKSjj3Pnhx
MtcBPCennjpxL37VVchDdwU8+Upd7z3Xco/uLSatd9F+fJ9PmcXOEhT3Ejxn52dUdwTw+i//vpCk
W8PaUDC/2OBPJ3VCbvzGL909nA5TTFAk4dBlwhbXkD0P6kiFFpJFaWjsmKWpa99llCt2KU1w6svK
hUh0DBV3P9htc3NIAZ1StrjmRZznA/1VQDtfQ6zGNVJiTH/yCQyKmTBvuirqXXHwHvdGAG27P49g
Rp4Ku9OAhyP46lNiCquHRr31zSDLZJLyTmzK0ZmwHCR3u0AvSDjlzoJXcRDi82GK7oldAmyZ3dwr
4akJS3Gk/2FFQE0pP7VEHpZniIw00FxNbyOWhzL/5ooF/b0Z6cpyzvOezm8dRFROOw9ZnxAK/6m1
2O5TMJht/mHAq92NI1lo44LnCZtwk5ZLApoSzcfmam2rD9PcK77d33MdN41jaE3qWsvcYcGjdGTI
TkIiB/I6xH7SmqqvNguLBhr5SvaMj05anIP5XK6o/4cqgU6tzaZtnoQVxR019pshJOgo72CEqMuE
pL7VTa240F2hIBMOtgsO6ueCfNP42Y8wr3P4Fr3xv817WulpGN0pV9s/ZWNt9wrKzjrTXDV19PCK
LCV9pPfqJtGI4+mN52MMx23HStXaavxiam+xaZUjB/U1exqF4FwcVBXZ0M8dgHvaOeGm9KF/t4z5
B5v7TDJgFgsJZlI8sGS0Poj+fYQBX5unmb6OO+/fZKN6g/Ehn3rT9EKGL9pcF+gD7mUCfuPm4roQ
OzkdEvqRYHjRwS3/0YOEHyg1+VsqWgYh+FscsVcops379fwibU4YxRiBDIukE1JW5LlCfvQrPsoY
bOIsgN6yQYkknL3pCmUERchckIWEwcms7v6H3cppWZQI43wysErPHGaEaZlkjV+4Q/ahnQCiE5x1
g0uaVO7N0r2y8aN5zry7EHk0/yNkPvXfe99lq1vlN2oyASWhEQxrtuJigCHjb1UDdORyD0+OdOgw
5CTCxfBAzUDw3/T/A6BFk21OtEzs+t3cs+5Ho/u6cbgjyuChALby9c4/1WEotRqZf84vSdJctDCa
ByjA6zqdEjIsr3zvI2oRDQ6bUfkcGlMK6F7G6KOjCw6gtIfOZa+IodI0BiWJYT8KMhCYQIoFrwM7
ZdgTrDm2jD8mPHfF6uhYv15l8bsmSpDjrGjWLn8kZjvrKL9pNIPXurkkTiVxGfOHzwBunnMkE7Vz
YlwolR0PdCgoxSDI2Fcg38ucy3n8X0odtHBFG7AovK3kiX+rau6vyFnMnPRCE86wXIQ7quWAaYPp
AFZ5myg0EapmpjEH9nDQvDsabgxQOMGXtA7BDd37HCvGLl0VyQAMT9gKqj1CtJ+NghIW8Y7QXJ07
hi/eCTa3lE5sFyUBYqBEALlP2nqbOOll4y6ukjNjD0C0VcPKgeK/rd7RjXUCGyHEOZdsPI8fmOSd
8rzADsXnGsV55iuShUwjON6qQ8dreLTXzn3+VtUQ+NhC2b0kNCKxpYBh0FAGI+Ej6uTesUZlVgXW
h56mvg9qKeQwcuItoh2iFtH33Fo3gGZ82DZyvymZJitxzNxHJnlvEO7d2AAOTVDZ0UWH4Hk/9qox
W8MwFrvhazoL+EQ4U2Hp9X96LoOx3rLNB+IWucmuFfT0uqv2/nN3QMcEe3S7Y7U9KUpb+SrJIOAq
35G+lkT3YOuWIAvS3tzgzwnGiH/45oMf59iyjeEJIJwSQLN0Kn/USoXzCQPTHfCcltUjcugvWkg3
KukjpaI7wAQ8OUIzAMekiIMUKsUL6c1FymHXvv8G+8FWxZhq5UEaes+EZ0Iu73Iya1T1ICZgPeq2
BPXIe3/3zE5RBY9MA+vqycriUx157busQ2fQSjyxIps+yqpzyOVqc96YLRd70+a7yZ5/toYMyJBT
7zBMI8+YAhXmGM0Vb5VrEcZXbGPsE8H9FtS1knF5rMhL+DbJoWAluP/DY6vu/CTRPkb+VxhTWWZH
/SGrC2I2oC3lsBfi3Pdn4FW919YN6RW2YSw2ee0MrPPm2JHiOzRa/lg6yn5JoYxR1LoFhBlQUxev
KEoaufKUXR7p8nOQMAryg/YogRv7fZOCe4s6YxRxKgZUTkviP0BPAxKIm3L960SeXpquGzL6vqPI
C7s78Y/m/v8ZemckpxR2rtAyHTHUDRiKPxzVzDHxcqg6RvT60/yfCYtklHXzgcDldk0+tVHXQlOw
mSQAaQg+TkXtuylQlnDTj5HuFvUh35UPPk37yHa2chnIEuReNNnInGklsmXaSHIOVC3mxBK5UG7x
e4U2JTsnN74USCLGHSIZIy9WravJ8VCXDbX1qQS+L67YP9qE6J1a4sRlZrXWs5dlt2uFXtjhUdyw
eO0StVPjG5Z+IgYmxqGVC+GF/DaHNRhHJWiVOA2ngla+gx0wzHSgGQS+FFakAMLI3mqSIO0EgZnL
Lj85u/WEKCfJEe+qSxWn82LrZ2xw8UFVJTny6Hi2j5SfZNxftYfNb0jcdDcweahBCYfY4HoZtcJi
74C3rCHbTiNpcmZ1lutZxvgSzU8616QvlvGIdcGzVU3wc8LhplJGiPu314aLHC/IZF/qtFj+4daG
SBxY3WKkF4xciU7urZxt+sRUl9pg3Dd3r8zlVVqBwpnAdT5ttEp0260cUQHn9BYSr5ja7Ezjo7mM
XjnfqDCiuTAWhONYMN30vX+7VXitAmJVEjoQV1F/s0s0/VAaLA9zx+OvmSqgPFl/2crYXQiCFWUC
YJNd52wikDPHOijpjA3ZB8Sg3XZRTdoI/3pLRk5OzDsKji2JhfAN8bpST5qR9rh1gRzkr0XX/pG2
IBgYeXJFgiEJAE1B65moAiw64b5QvjFZGMN2TOvt+GAtwC3nuHznVORFSVoifqAlVq2SPD3N8XxW
dz5ASWqkH8EwPhGinVMQ+N2XRzELaP/DiZHjtjuGy/Hb/ssMDoOwLxUf1ZL4Wu1EF3iZ44R5dyT/
Ha1m/mPR42McknO6BqbTMi86k+rmVvcU9mMhHX+JzFJHIISSN61bxOrxxBMXb1HswLILL70NJxMq
G8hxoWq9eqI4rBGryFlxNNehth8i1vZv9gHvYRqxnrdYXgnHqHHIGDWSIzhIBl1lZiianJnXQv5y
M0kszC6eqQTO3jKR3LZj2NvqC/acyJ7ehi/8QmnHY6GljgQrtG4yWtCCcJI6XNFzCJYEnNIDWKS7
s3JE2Mi6L8B8ttPwQiqpo8sBqa4jppFVEHlyUeUxkqGmWQmfZ0jE9sDhoNCtN8bakUhwDitp8K4X
wadfSoAHZQDOqqs3DzJDY5mKKx/LPDbtgF1LaQBk2Iuyiu9nKOYkpzerqymJMRhlUv0/fpxda3ny
B9/jNNGSRq6nrAh1csTNl5Zp5gAejB/jMyW1a2gO/WnGAEJ/mbcAQGfNB5P7FtaQ69DyYdzB6lw3
zoUeVFUszQrgzwfM5a7lu/Reja5BDhVzzIg/yPPKI5RL+qnBovxl+GMMcgBgy4TqIqbDTE8El3v9
rJ+uXshTN0m5dtZ7XuJICXB6KoPY37FkfNx6HwmeEeHHlrB+001WkaLJEMqWRvA3RA1meqY1duN3
qeIymp8iUAUJmBVDvScxDsthWBOO6+E/GhLrPaM7pZFQNFzXYndvY1kYu91TkBhGuDIIw3ArLWMw
SmtHhi+25DQlZRc+pyXPcQJCkKc27c9zPg9NWrzeiTE1CgrJBcPFF8SVxnzm7K+WCfozz9DyqOIV
YP2ghkkntATkAEMDid79oO0Cn0jVmktyDpiHm/0ycrrxzoVwOgaPn9AMEKv2i0xc4DjBI6Clvl4u
oOM+cNlb+9ni+djwDBmTua8U4i2sxf+QHK6uKXZ8n/O/+quxyBMLwFL1C8xVG7t/7C4GMyF7Aqzv
2ykBJPKokPcV10ta91lAF6q55MRv44XZTmJNhQNLVmPXQBVvx1hm2JtGD0HxUQYx0l2yIcgsLrls
grkvSaUbxiXZulF3XFCvd+ifrEjozyIAMxHvXZ099zx9bu2RTStGwL4zPcAsDy9nZvauuga5NPV9
XXfs8s9a4KZSdbMrh8wdEF5oqKmlMYsfAcbpP6zUzrk/+hB44AriPyiyxAMsb/Jx3+Ftz08KEy8N
ebDhzE2G8mi8ce/k8QuaSplvW7EIdY2L3B2zff57WOZu1l2t4Ut+YzmmpVaiLkjXySe/f7OfsSTN
iC5IhT7seasIOnUQELegiyvC1JCH4+WhETyClT9Nvb317TGNvD5POf4xLjKhRyB7SG1T/uMo9ViT
Tm0GomZ+6DJb4D4FxVffQ3hM7uFaL26V2OGeth/n2dJZRxlukU6Z2uDqscvhbQgblahxUdTCCigb
2/TMKaYmReutaQmzy8u6s8Asz/OnzUAcsoahmGBgsWpPX9uqFu/AMuu+dz+ETwG8Vf53bPk1WGfz
drwickgRB504FOEIvG/3vG68yxFleYt6e2ELpvti5aKwXMD3XtLuU0lnaMw2CBchwxepHYjHFZsB
wGUNi02GuNaDTFJ8O/c/54wmQgroqg1I9sagJ+uUZQwf2AQVvaJ0kVPJC1WfqD+Pf/CsTpeCEz2o
lgdrPfsVcQSOLij3kufgjG/Yvc+NmFqXQIkiLTh+BgWHj0YfWCqWmmYGI/jj3Q7TyGRxAKZtxpJH
7oHXZnScMBpWgSN+91DDdFIvJJPj0uKljExtUyofXjHwIDDPIC+CQGDPPZxAfCQtO/4mhJQ2deKj
vAlogaSLBtCqtEhfzRcUpAMx1H3P3Z2Tk3ec1SOulApP3WNuub6Pi0bW7l5BvvQ/Zvp/yQAoaqrt
ArVVMzUWp1yeEWoB2k/NBrbG4StOFoLzam4taKRuIlrx4Ktnfwjbt+fM+vRg8+Zv8DTmQI/F0Ttq
FYN69bYg0hLPsd6F0KvCLmKt9PtQKiHLJ7PRPYdc/9htpycLBrAxcsjsYDJ/a8gDsBusCQ6NeFjk
dgw0uIWP87BKXfsUfQFLFYI3hijqr1k4ZZT7XwAaYicHd9R8SbyZCclAyANXCeczHEfXCP7uOs1d
YoaTl48IAutS1+6x4QTpZWixL4lRJCMvp6KjcSkNBPS+QyvoXroigkLfpk+ezW8Bg0eYURYMXm6f
2vVUFGjVJZ2ElcZjN8+kXAMqvrxGm95g3HSJEk/AOUiOLjHSbS3PSy7bkCbfAkw50zCNVXySYWpM
T2fBrBIpV4B9s6QzImgiGV3vYj7+nL/JkgBujt8nG3kFuSsqNplprHTU2qMosRtqSWp7LtN5LoWa
/5NMUF36MaaNaRzgOBRccrs9pq/Z6+QWiRPhWNcApjSns9LHBmRq+hKiD9Wm+i34FLfP1l105v5B
9Cl9ZX5J4ZCCvRUEAMn9F5Q0KNS3KfukxbaS2fp0iXrTwBiS9i9G6ZWfkUDA2cgPsTZsMVKxXx44
jjswTe0tiLvUqKQQHUEW9OWJQudhAvI24iMyQXQ3xQQjKtVyQ8dh9ctIyEBInKCSxWtAfLMwDvVf
NQwr6LparnQWBD81m3K7MMg3Aw8nZMakCWQjfKCOv//jKlzWBbUPEPkRLPO5/e9MmP8rwce+cHL5
POUPL9jLen8b9Gc92pXoVlw1l3Nhyb5skFMic3/EqgLYE0UBLvYLkqOFPbErABkXsYShY/yUSxUB
hOUUkzKsFignbcpX7Z9ZwRWbrmNzWU2YRBK+4m/yDWASmvwzYpiM9aU1QGnXHDpxxnJTAZOD3Mqc
/YJvd3aTTNaq+Edcoyi8XUK3CAiebb+9/wRLO9h5UHIMys0Jkt0CgGpUuxVNK6oP2HaAaxAgoo4O
l6Qkrcu7BomKXopbf99dg2WdtxboQf0qDTq9w9T0ISHPTaF/VU0AaDu83VlaKjp/183x6LlHLzIZ
YvTf+GLXvlYtINYlKqhBa9q6vOaHc8A0Wevspw+Ee36sbZtYK+H9cWH+4nVW0efTV09ntEg8g/vF
8uf6G67ejPq8won8VXsAojDNX6W8B+RT30LSldBmMXILXDqPLFzbcFDGD0yOiKPNpHo+EW7lOFQk
aoA4ggrIfASJvgP/zTacus9EH7Vk94LbrzAWMsqwu0N4vh3NXnAZfFpycIdh2ge6Wnl5arvsH2VW
DwEIcoXrVAVTEeUZoIIdsC5J1VHF9PrRp1jXPIllSaBcf/UBHxDkgY7z0lLHOtNR36bjCUyhzyKn
/SuIh+TWPrhlvlhpwD96iU4DBnlRmWmutgBvsoetyl7LoK8ay1tpe/iKP/KNSWX9Uy9z7jMuHHJB
RvL5nR6KMKXtYlQleiQyBV37xDWq3V1mEauamo40aNdFsCWK3Ko21oTy49DrHQgdZaFN4ePbCZ6+
0e+xt/uButtSztT+aAKx+bbyDgdKu788hIkqPaSytMcLResVt1OP7bZHB0czDP0aaSGHZUs39Mbi
uZm1niLFGLiDawmDAlWIIUh4/N0EL0OVTPXuNlHbXAs59gxpOR29+Qc5k5JRcb+oDlibMFkGCsNj
MdnjmZT3jeugVqyN2h4yCdMyDiix8Qi2IO/OEJ8a/xFfF+PoORLqNTdfBF402YAwEn1CvtEQS1Rc
H5JcXS20dPrSKz3RkGmkSQ1F9LcpZI+cVD5R+eRsDoc9rbaX/XIm4/SQujsWaEUMv7hfX9xNGf5z
zOsMm8HaxvhnlRKPeCKIPsXutRXUvgQ8z05AzQXQp8VafB6hGkoXJYTOrDi/msamgP7lpgMmdB56
MTaWdwAV0DWudajqk6i2QSige33rv5B8RvkaVaTkMzMazFIwvyr7DmJjH6F3/tfnQdcjSwbF1vy4
wbfzuQOB8uhnNPpfMnp0LqDlJWzOr5Z/BtKGiRlwS1Hs/rGlfusjatqSW+RmVkWTL2TNrHkIeQ00
Ys2VUfmMMkTEv45jdm9JuJJyh62GANTWd4M4JVUXlorE9sFkOPeis5+R0YjhK+1EVne0dVoR2vlX
vKIsWG+/QxM3WtZgreznqUBohEooMoL/u9kxdnywf/XPnI+7ahXsfbU9gAtm3se1aRYsp/wSbPDe
h9YGwaI3s8q+u1N8QOH3XWQudpB/IuagWEJOk/eGbgaz2LM2sd8t886G8o9dY1Ix56Ce8b1PoKfT
MOIvNT/WQ4dsYyZcUPeuXUr584TP2La5OoyMVCb8cc9f9zJKRWmg+9/Kyf6iLX8SKU4kn8JQLiM7
fDP8gaBgOypFWiPYmHJCSWRdvMMOUYMKAH/qEAmkWNpKz21aoDHYoeAntekHQR8+N0ymoHzOf91k
g93JzKlbMq0NYDKm80EZXp+kjkFstKKxqXrPB8TeXikkacDxm4hBAge118RDelUhnfxi7lywcftI
8CoLYgbHVPHBhUAviPOWLLwuVTWf4uimhgvkM1Ix56Q/wKVoxs3Uc/EouTK7flkPxKKdmS9AhS4k
ll4jWV4OWIIL7tg5mG6ay3Jqz14ZgNRXauEORmWsa2KusFsRsK8DyyJGu/rNmpAt0M0eeM5LAPk8
qXe5IIUdYhx+TqZNt2Py8FMtehlrDHZSfH7MHwQYApo7Xyv2I07SHG+Qs4VwLtiW2bS0BsTNhKJ3
KPKxcQclAVR+j3LDYIvx+U63LXDLRX+W/AjHQdwjWKYgiqsOJF4L4a7pdR76gm0DcH5IsbyczXaQ
oC36le4AinfzUR8peJgnMAJ4wU0kZKMMr/+bafKdJbuiWvXNPCUfLCdNu2ryfgS99K+a0P74XgXw
6O39ioqPJxKILo3BIdNS3mJg9B7nSAI2a/7LTVfDmSpIaTneisTduJLWI6SKoljWmtNOnAjALVKS
bfVHk6ujmEoJ+4oIVmNAh5uMPKSq8M/GtZA6Riq1l2GGP/vxkfCUD1Ce2voroCK2vaH6jtS9wYwt
/u4Ya5LwaphNbrCImaUzfTKiwMx5IZeLGnoaWBnAZIKZUKHyFeoCgTP0VgTegmEgrV5+urgd3Kos
OKfeB9BUkdWbE18im3JKJO98oOLNbXFrHET4edxmhYZEzRUWzkDnlndTOgJ6PbN5oglWfYYTaNJB
FSZkCUTRXZWPIY+m6jGLdwmx9jeWCbjW+hLEPi0eRql7DnIde3g2aKojHXlF1DL2ToJXKMorzbWm
m7emEqqHUlUX/RBpxWczEJ4hrTWHMeu2lzSLexlKvugUJKLxzmMCO3hwS6YNBAbSKcInH8RfhyXW
uSomv7icWtfglUj9Qarf/KDtE29qflEElsIEJY/Yzu8jauHPsOuJ6gvnM85iWvZfkOA3JLWSM7Ub
wBxI384GuVDHQcAt/kb36Se7TAwA16MemMtOKwGB72II/FMx2B7uTbnNrqru8fe8ag/Eg2pXFBne
i3q8aJT3BiZLiAHuVfF2yp7lcVfTm79hoDTstXqqLKazSQqKyAKizPhWW2mbtGC3REMRLYAimGjJ
Sj7OClCCC6FXCY4ABa0fyFlJ048u0+px/nmUTseuu3oIVhsQhzn+Mrb/CW+kiQ11FgzFUa3q3wtZ
OTUhjMh7OED0NuBngC5ATmrjy9E+EZRAK4O+3RN9HtsUFu0eoQNBStzMM971+0DSeXJS3SwKuv8z
J5SfmXcOtO3jO5NuNyBpwFPjq8pnk6hE/MBZgKsr+E3yhMv6GA7PebQ1QQvzUkV8cgtIopuyHUrh
JvdHapNtcTRiAzbNf6HPaTdum1QILsTISO28Krm5DMuAI/VyvG1r6/lXAusvHcFBiQ1rbJ/Vr6O/
fxdAhVNRvnOsA1FBMzoqT/vLehOBBunObimyT+zPyWWzE7goLV6dfh3/ImYRJkemSiwjSrDyNZ9B
+vB7G/vibi04xyiCejDW9kCmE5kDr4OuGAdY1cSXsYNGxwJcv97kS3t3WM1ZFGaOu/H4+ZEcUvK5
lRL4J0iB2Rj5MOCajHi4ezN+fr2/TDu3uvBfOMtRGoH1TKWNU4mUGdkqVJ//cF3T8GApaCsrvKji
PfVJZnH9aUz7wb7ReHbeR+xF2TsggUIBlRV8OvtKjeQJydcgKVSWKx0Rs6C0PppnFrnG/rZDPK5v
aYR2dFgsHibEHrcEFKMaRYNEnKerVvqqvtbH02qfrw1E8bAsD0FY3eSHHJIDIAe8tpHC7+s9qknP
NAZqG5ekOAhXW1vYvB8h8uOFmIJfj+D8RrYqlRUDJJXIVCfFbfoDFEYSeB1NUAzFxdQbfykzBkpL
hKzcd7pCIPhDHBlNjg946J2Y/bflrAzcI1LA1fLp0bUh9cqu9KGQkBuMkSINRAK590+epAutohZJ
nEb0tnoxknzNsiX3nkRb23xHhvvS8GDOMwC2ye1S6VRLl/qAtT2fiAfkcR4YlIrh7MD4dSHu8pBs
Ypc1DSM9OuMCdSMOpFbk2ruiXUUkPZCEiNEunjtgpiYlLV+1Z3pgbrVZhjleVp0iGIOa/4r/7VYB
NI7YdabSCl+qCj/44FcN4xSr8loLJlh+w6H/qf7frcr//bdn44ILx57OvLOkhxMaUfY2IyhbDnKS
cBmeaJ8Dh3Vx8K4DH1opO1ZphCAj0oIN6OXQWD4xYFV4Gq11h48AFlwoys/FZ/dQiepBnCzIYv4q
vFpoLNWoWVB1XxcR/ESNGtfASXZMoq1RnQ/5uefD/x6gO6a1whpXsoMCvA8zpiUTPSvIacBq0BqH
5dvByNy9L4TCKex5Cs6Ako5aiUvQKODs4H+LWIW6mKuBNLoNEgOWQuKWU/rMnZ5zQiKGDt8ER0Q4
8VsfnCrGbU4YvS21cOv3fJmT4T2GTqbLS+IzBkpDkxY2JZwl9yIg1O1i9/xYYjlB6Y985TKHkVlD
m2l8JdOa4hBdYQlPL5/ESAdKYddUuFXD9agUlgtJkcUYIwGYKFahOgFNvDZofDR0Xag6cuOonAmG
MqLFtaG1KDEA74MeqTfoIBZrQbUmk4HFPay89CTzXvVhux/o99BDROqJNiBU46qY1AWhYDhvYJuH
K9/QCgxQQGZdj1ei2TjT7Ad/DWjna2xuiKCaBe51nSUO/7xj9EDQvENdo9dsO1QDTBkW3J7vmakp
fEZnLuv75RuIdIDQxyQ4wAhXK4QHUY2IaN0Y2DSmYoWiEU827zYAqRLjQr3htFKR0asazr9pDdVt
omoNLbE4lK+tUsd22jftkeWAy1+YM1q16blL1MYkO9c9F9QN/6ih/tn+fGn5zceLU4UseptoeIpr
KzhJw9NhKBzk2WlO/c3H1hCWuEBKIY7VmBlD5YooHrRGdpuGRCd4Do8DNIyNB8s+Ew4OoEc6NX1l
SDG9BMNjTRmWVTKoEpOd2hIxvz1R45fEu5HZLXtWC6IZVuUxs/jvuzlJBBiJLiK/06efh0V7+1+1
0vDlQSLM2WoER7QkqMuDnmKKzVN9CVyjh6o8X/ut9aSZfyq0Ick89ltHGnDzosm4bSlC4DfacZtO
nQuxcwb/GOx5x0K85MsBzfiLOm+SOi3yhL7fLEDMWuqTaJB0VgqVOeCsmUJlU5LanGHKT8aRqOzP
33ynwqAiXjI+EfpHWBPnsYnZO+DoPtB/jowBEGBlkR8VclmI+2jGVrJFtWbNSewFTOneCs2A3/0u
vufpY3Q0bWOpxLrhKTCFrB8JRNDbqjhbWnt9IypcJ3RjSLtjYwdDPWx79jr9xeWmn+AqQ3H7jmLZ
++xieF2Ba/4tDzn4AMDL11VY9wbjqcUNzfuGStv8uK4h14vK9f0kvC913Ke+Z4uR1j8BO1cF9cTN
p5QdGWmUeLajTWz2vfvh66liP0ZbMGTSC8vosWl6R6Gi6PSo7HIJN5WgUnYdbdIN7fSnoXD52vmb
LW4+dafzygcSOiarY8CU4CXSxJqSJGkCevckEpsQ6sHL+9ItadHpAwKEv+8S1V5XZ9lVQKUoFdgw
Ct2ELtk6OVAvtkdS0L5LQQendjXq4pddi2k1bk2S/+gJvhbegdAXz5uKbaHbGEqG/PD7gAIzzySt
WXld/G5AUSDXnCC7xA32FnVHnTRv1zv7JcdAul5ePrjjdT3z8GxEUnASrtg5wONSAcYEIi4Omnat
6c6DmUkjSGDXd+fpQ4BD2CENOsX6gtvLQApBGNc0aMGnaUHBcaRqLXxp5yLXaBjVqSisoYieObye
9o20Qm9o8kzIiNtKu5XrQwAGGf0M1iazLFzamStukEJaGRjkXMcBwPobaHVMfxgfhzKw2sJ+tbt/
UWEwFLiUSiVk198ceTgukq7qiEClIJQLEzQ/ZOKsLEF5kJsnH2WmBeDkSxJYS0OV3QW1F2adHhRj
Ca60dGcY1CQNggdG05PckiLtF3JKB51Ej77DL2CYGEwonfzzNuSiFFgaojbxo9wcQkIaiekwZy1/
P7jj/Q2+htmSnxWVedFdI+//ntW4USWzcBOzzKmbq3TVhBRnnmpkTMKzdAMY3fBxiuQAfYDIJeJ5
rcag3nhg80V8CKny8ViKQ0W3F8UT5a1LdFRqF6CfpGNaUrRiPUKtuYbVrkX+j8XMoug2KjadH3cH
NV9XMB63u+z67Pt7Lif+kPiF8zC7xQwfrSdd1/Fq23dPEzLASLSqJ/pEAv8A+Y+1/2hEPZaDEZyb
WDTOTvUdEzM7xF+y/CaBroIXO4DT+6l1SGqaqTBoBrzHk83/TzAnKVBfJJP5idvMSPIBBo8K9hKw
A6epN5fuM+5P8ID6Yps7ZhORj3P9RcENDbYEJrWVffRqp3m5PMbsum8vDhp63H0yD+DET1WP3vaU
zJdrhN7z8ZcIOhdViRPt/BjChBTHK7rYyC3396hVd+z11/H30asg6hgnhoDkcQn6vUway5O39V2H
hQm0LYtiTYUsfPUq3vxRHyIY81utSMYNL4mWazrOUwWnNpiixYv9jTp2c4vC80dip73ujJJtciIW
UkKrbyDpQT2jWyZY0x7GPLu2ZCCURy+GHB+AST7CDoZGrS+iuv+FnPpWKrUIk7E5/y5PZG/MaGM6
Jc/kNe54exaCLGBl4YBJF83lzTBJJnofHHIfFEAUfMJOraQ+AZw+bRNf60qKfKywmhjE0SZbUt2W
XQQaR2bRFVxAxA9pUGXekhgEf6ZLpHpcY44A48ExcR2CmYHyB4LGuFUMkbLBgzMhqvJHiusCtKJq
mTRfHBf6+PeP9hsOiahGqsG6dnHsTRIxpCI/jjMTuqIwf0HK3ylSnmofmeDKYwjKYD004MBAjrcT
K6MeC26s85hs8d/eoKvk30hhGD57FvQXLTi/Vgksr6fw6XtF3nxc10Rc7QQiGzZmoxRV0o6LsIpV
Y+aFbtdfhR9gGqZkeYzuow1QiTSVpZ75WyX4M9Kyl6TmQXIkioAsBDSs/kxOI4Vo29H0GpoetOmR
jLEhW/4HsL+/4X9OKI2AsCa1alyi4u1Eaa1pD5pPkjtKcA7nEi+/Zi+V9LxVTXleMUW0tY+uOavJ
voFdPOvSttBPXqN2n1btvn2PKSNEo89uQyyW/9+/H6jPsaF14+EtIxYozLqOQn7jpKEUAkQxwQ33
Azn6RLVSO04FAhHYaeids2exfl30exCqkpi55ykFqH9SUMoS6VdEiTjKjYNHGZlwEZ481Tu8m+PQ
GzxgLlO7TvWhevvnHHThtqlLCddGiRAZAipEYzUZgebV9stJLTBa5SThgjH7TP5YhucneUgu1ZHK
dFNeJQHQnbwhXi2ZAQZHwPuxfXVnTudy9/vq1ZKgOZ+U5q7+W05X9quHo69XzR+qUb9NXLU5ib4F
47pwLt/vYuEberI4bBCsjp1iYQKzBnkb05LVHXIKcfAe0AYJblr9XKAMDssQJPI3zM1mL88trc7X
ni1DpjNyRiJ+YMdEyMvWdqX4HhEdWgpzJu3mfTJP1Um1QLpaHev6NIZLeLpOivJOPeZLNweCwHPw
Pi8Ow9kEUNE43OSbUETkyQ3e8bDuDZSdAk44LHXdbxUmDiDB3rw5d9YWq+RXy4QNLrGuHlfD//EN
zgEEHLwzA4M2hC1/0ls1XQcRznNDDmNlg5/CRXX4ukp/551STDIfIHkNkVDVOS57Vir0GqJ8vOFD
F6DgOQEuS/LgsAOXi2rw63vhjmN1iOB1vCr2+vpnrepnM9uVOGzm8GOKCtOmv77F/QpQmt3CofK/
3pLE+T2ZsGh5W2qljokxrdLhYiq5LVzGUHo8gnA80sD2OR/fah8le/BlqJpYlPSJFkJYlwjvi1AW
kxoK5JarmIRfTztMW/6DRpDce/GzpKjQiTwbY4IFpJbw0i82TajNv70Ma+TpNXU0GhANQFp1BBov
ER2rrSftv9jM5jP2OP+DBo3MO3vOkSg0SYVDWuWt55u1ObqfMPs/UOKiHnkt44HyfHLSATOyxtsS
H3hs10zcLKp6JhlCZWrg+M2DN6PqWmc38eBaXQxUA9DXinLesCkHwG6oWHxTgcmNGdlpMTJzvGd5
z7WGJ1EmXIHb/eNylE8JLv0+8v9KDYAfWWDMJ3UiNjyjZDWvlEySTUkKvKmOSF/9cUhhWPdB4GhB
Zkb6CgDfN4iEs/INwlZG74IPjFvnQAaoOgI2Akn8D63BfLGAYj8PLAOqUaqWBkCK3qjR5RGW3MFf
qH34Z0vsPc8/T/U5meb5kbLo7+KPPFB3SnAKiKX397gxc0FrmWmuX9Oni8peW3LPmJKCRJmU1oIq
gsO/Kj+3f+wxxGxsITosNeZWyTCAweA3EWr1/qFSYeN/4EBqj+dIkCbBMsquDiN55tE+STTDQZLs
IQNwjNCYooAQGMD8Bg7FH+165cm5rFh2vapbOQ0KD8ovnJ4ko1Q8iokJX/cWzhm2g+odrO17NgsV
TVsymPOZDddX/oC8G9YJwz1J13HE1/wQeK7VGNeW2CEWf/ipUQGvQwH+7YsW4uXUGSOxyjH5TtI3
5MjWfC6kJFSSgcFS8h1mfuX8rlip+wVBhrRQ7cRS2LtZZ92Al6WpRuYGQG8n87XzXiXbaEPmBibN
lFy0Jnx0MlC0ThkZ/g9wSvaNWRN78wnnfwxAy0MsoJxF8G/mF7QPNotWb5OVDk1pIVoYMKzPhiyk
FctZX65+dlM+1j1t6emzJwHNJwlRURl7RuWXPSD7JqdvmpVFyQeqJn9JF2PsCC/9h2YgwsVaHhc1
lrDO+XR0X5pZq11YEoEiOKvn0gFNcIJ26EEvN6Q0sq8qEgR5g8eSoaZagJ2oXpAh/JWTMc7hUFB6
Yn3z1hUHn12jve0um6flpa0FhdWhwYL6NClNph1YyVyoNsrQoKdxQ8JOFYP14qph3LoTpmoUSnbK
z+THbynLmIIdEJTkAfsSdNR/WS16f8KCt8/G/xZug8LEpld+OhP5XJNVjCDJW2qQrZljJW3YfUYm
wjMWHg/ZFpOV3wXCq+u6sWMlMz5pZ/7woRXH/2oAZL5fI/F4/JJZFdzACfaV3pS2rTWxTDbKT2of
JP3CkIrmBtRDmxo29yGd+4GRu4ncbDLdnzZ2vNbY11QQoe9TAoHIuswxrGSyDi8SY5HFTeyp9flT
MTd1XG6br7zUNwmwjiVOE5jRetBf3CM41evSLF2p44Q2RiK6kP58NJTVqtbX4rjTsTMa2RqC/0y2
P44QlVrD+ZVIuwqdpCUL+GH5NkXK3cbp78+TrYVJifthgCHfRaR15rLglleZ4ZkUrfLz4XKoydMH
2hWplgT/kQVJKaEP0HjzaLNIA7kRmd91k6/UdjX7Cm9awDs1Iv/qu4RdRW69Hjoo28O+jfp4bIFV
A4IPLqElrEm0vKfcVnCTtscGIeKkkxiBaa3Tsv2S24LWKvcRe2dg2PI/6inz/uFhDA7fUsUNE0V9
TT45aulM+AxH9xJ/ryjyqgefACA+vAJnBDo27lcO1GzmeMbAbkfXXR25rddzr/67ktOkxuhioksV
k6aH/9N28USKrJcTq/lr5PTKc4AygVg3opWTHcUjxBQs7UUmLiduSIIYWNynqR78mS2EIo++w69O
a3oCj17wk92ljXNlzWljtduRjkkRkTl6+O5tn7zLOgFkVlW1a6vil8oPjA4x/Snpa61jZVD+Q9fq
AxdT3EmlI/d9YW0Y2JKPjqKjsaYG+0j75y9Coi4xfKLHlVNhxU7ZWl0Sht+RiMiltNIU32BOyCek
5oo+b5hO/IvfK/oWqQLhWRN5aADzEW8wYLo5Tr/egvbdDln+PpOhdxRcfwhPZdzR0Wm5k1J9akxp
PWDTtG32w3F/WTyBPlSUQCW3TnszStTsTjNtLPiY533vJjs2XnBv2vzN0DTnka7wu+Ov/emYA8MG
qkG9x1lgBPrl2xiRJMmZs9IVxkhFObzk+ARFfKZZ9e4q6D3epRVofT03e3AnIWcGEOB/Lci1U1YN
FISDe5ao0kx+5T8VbI3x2krgw0hxbH8Rq/PB3fSF+S6sCdtao98TA/bgkAczPWEuAUjxKIqNNCxn
/Adqxe00EbO+jSUCLUOzlH4u4prjTXZ414Fmo+6PEu/tqIC/cIQbaOWWcRVo7L0I03TbT4eOV6x4
4JjXSqRyL5vZMpt3RjtLeYNZ/69JjGzm7wl+qUfFvbO80uOxlt+Ukak3dRdH06fvNy1mLOrDPufV
nVUWWqS9tYuA2fub93DMrWO6x+BiweVLT7pl/qhvZf85qibTu1ENVLk/0O34qkUdzPFyQqJUJB7A
34bj4KpoGPm2pMF72hAOdAfrYFFpAA49s9diDKqtUQ9pjg4X97E0CPW+lzFdJUFIo5eDNjI6hSsj
+ef7VJNBGhJADGnDIe8dfBn3lQcGiP3HWUEMizr1XJJHAou6kkor8ZrlGwFpIfUbGVCPi7Z5/sD6
n4kvb2okGR0u+dE7+Ewx5XmLIptUR9QHl4+F4MPSRDtukzqk0KhMqwOB0cDivy4ALcMxIwsyTw0m
b5Tfj2NOq2z54WvtyXUixx+bCGTp7+e4jjJurfW02u1sm48tNgeIhGPBZNJRPNtPexQghy+NJX+t
tpPhRRsiWomQg3wDyvzBQ0KbCy+QClqQqWPD4ShrXAOn66/WZ6aLGJEKCmjR+4U/76okSDjitV5X
E/KAy6moren9XxZp9XINRSqGqTIi7klJ125I+WCwVBUZg2qVH0p9cRDpuC1S+12q7qGQuNy8QZ4S
9To1LnbaFhh54DpSh75rb4T5MEw53xEKZFpLeFML2RYNaY4/SNhjtelG+FNhtEhIq9Nf+Q/1NW3Y
RfW/re1yUZb767Toh5vB9EPJ+WrgJn1dTMB1Ip6Z0HEXdVEqOB1ZOqrRISZBxkcI0DgtD4xcuY1G
bGPauTFDGKuCDrsCzUKWm7pn/jI91ZoUwfElCCPLmBNwDGaVfdmYutxs2G93bP6G9NJP3LGT4SPy
SN2q8ch2TF6tZhVgR3lOF7mILWdkdzAu3ERSiVeW+88eJbPO9WfengxTtRZdzOaVdWX2jlaeETM2
mC26CtoeEDotjDJADeEfGST9zFyJiDIGBrnBkxh85x1bnLKY1dGASU8bx3BmV3tl5zAJwom7LG9J
6bo5EX2XYKH08/mbYHX/Y+0C97yOJTKTjZyRTmsR+2RzCeO/BvdIkTNzIGeu3JqH6wzTdFEdrnHZ
V5rsTLa3md3u7aPzRxGn332K+4MxH9rgyvjooFf+tptGg1fTOec3TlPgVnrYNDK+pz/cRYuqffoY
MyeTAyR9XkeaCAfuioPfVjxm50VFYmWU0DtF3sJNC2KXb6Cj1S0mdDUfqBG/zrmyEBhOZ0hvZK/4
CfzH7U62xar13UFH75wH0KVlrKWIN6/WZNX9eqkqpvr9KFJ2grAE0pOWJUhvyhiijDlOCluGCro4
vhl/9JxynLL/mWcMNvYtPB9lTdFhY8ag8bgTykHDXoF9yNRtSuxIqy/8dqk+hzvWdy5JYkgQNNtm
sXYBvXe9YvZ7ljPYtUmmGOgHitaL+QaJoWFz3fS3o594UZm16rOdBFKeyTA/IIkoyUo3qTqthfgn
rUsWiBRRfYWdfnVh2EanGKqAEIp4Mnq4Vvc5hFettqakODl+ByidinSAM7+/5y4/oVIFheuIU/N3
2A5tl58ZLQRSd1DTKKUX88KT6t6e6wS0BTLqQyiAa59SgM322mSDZO9853B+nHSD561xAQ/rKCac
e7i6PBqoXaU143Yv7Qsfm2njXbNE10adh8F5rsoyhES3vOfH9cpHMoIPS/sy9FELbF1nwaKKE8Z6
6SAE3jD/vdE9TFgCjo+ob5IV7jkGZIQzHEhZlQlJL3c8um3IKcG9IxDNlPYapsxgPjVco1gOfkm2
3PBhopK2CGVEcmViAs4njKe1dBxOo05Z0m/FptzBd0KHC3wdBXh0XbMutff2Ry2iL2BTY91gbmIM
QELXwPrhzDfeGLLpJXvJGCAh+C69Mkeld55Ujo5hFUcEAyHBRo9Sv28tKQRIu23vr7tiXwm9jVVp
IpZOQ3jfYxkiWcL77ERvGTkC9BV5yAYHEIA0YMJ6ESHglSHD71lKBssgESGCo6TTokl3P4gjZnrr
/JLcVv3O8YWAw1Sx6/rH13GNCXe8HprzoOB5p4efifjUBOmfvhz4j160LtWN30zPAQ5XtUqBmk7R
LqfHRuaHip75WX9MzWwlbNUlPA2vgs9R/OcDEqyAKNrCOwCh3MEGuk5Q3KZQjRoAiRCR5z+zRNta
6RowPpTUZxcIN6SPPp0DlNf6G9oCSFsQMw7KnKtANvn3plrW+5jY/fyS12jbQRf6OloMm55qmlvt
v3cbuUg3JUgrBZOKIUtzWLP6oxhzgh8GWZXiMrNubX+hm8DME7yjvGoHoI2VdHzekzo4ZRmnOQ45
Zg36wCJ77CJ/RbK1E3DVJkrnX/CtRChWdyAuQ0Isg5thbtVFFKH3UnAZwqvHevKIVrFgYoj2l3Na
BYZGNpQoZR12VA8tl5hF21vtP5BxvM/NKH/GvtN7fLakC1GbpG6iJZoQpjzinzH8NvYnaz5GPLaj
GwBWzDmvTbv/QhiZhf5o5IpaOlP38ZiR0YXpMxtqJaKmxZUtOQFYGUrulhileYJbSEOIzmru1ipx
1Qvv/1INDZJ41+ZLmZ/2JnQ72Su6GIrwmr4tRBi5Jyj+yuTgmtUcVIGAq15WUkIQj6Fo32zjw4eF
Bbx0mY4E7Ye1ExB3jbKmVjJGbbVwc2lv3Wj2SkWuGrYLOFYr8QWIcvhEntf9toEd0eJ5u1SIwNAp
2J64MrszRg7/qyxsGK3f2nfeUIPTvj9n5vdRiAyfmSnk5qXHV78BToK4Pu5z9GW8pH5DJzbg2ye4
+JQkdG3iO5GI4BoL0GFaBoCYtMvcexjYS07uWKIjdYgzikoI8rX6lKr0QxQmQiBFOXW6H9IK9erY
svamRXi2UQ18/RS4QvteZ5JGRFNF0ewyK83AqqaPPCEUk4ywXNQTdS4R4AX2hhHGd0mhzj+9n90G
A1iSfT6oxURuenqJvQLl6JdVD1x1Pq+vJw2MsjBwq4Go6DOMZqU09PEgRUZI14kifxLyUUlkZF3r
XN752AJRbvx08SAPzPb8IfL5Tbjd8wvqZGmDUVYemjQhAL3pGixtQA0CyjYERzkBaJF3net670Sb
6Hb4hM3bWU3yWL5whgFBcPrTb/z/bZ98KTPk6GnZ9OHJr4POqoKUAIzMWAWe9GcgA/lbqVOARpFi
1ZNS9+0sDlE/Wn/cwG3PG9aKVkZbVIRR6uDbFRzsRyMe18Wo6zS0khjxX4OTskJiIdk3kGpqXHLs
ZZsv/cR2lx+SiLlg/XcWh4Rg4E3CPL3DNkzAviJpxO6piBv+1kO5YferRPVPimH/XAEP6915RSWs
86nIY6SV/ScEcvS59O0ykAhtXOkabCdVhoIB0JNk2CF+EMmQ97DxoMtwDK1pll33lUF120rzPji0
uqnXz4QyV6OCO4B0KjIlJ30of/IMg4aLJDR9Y12TgxPzywBW4M0V/bRxOK1ehpPMZVgx5BEFCEAG
Gcay9X1C/EniHsMlwNuZkGk+cMD1S41bNNCfMdL6W0CYJyKIYunwVvaiqIr5wBZdnuBCO059mGW7
FwIRbXaULkgbV1wpHbQq4A5ODQdT12ZbxyALqN/omM98AZ5hrZdAvXSaGm7ePv41bif5ehPJnGXR
48cMZfOAd26ibJ3Wpshcatl+/oQPOCUembn5hi1em+FHpkbcvLo2aPQD4a+YxWaDenUbyHigXPVs
Auj+3nR44ECW/k9evl9BGjMKj8ZTUrXc4cdhdYq6Cq/+ylrWBb9Sgo20EnN91kebkLYOxy6LZri7
hsZ3yGsaTUQBlFmaSR7HuUQ67a7EH7fqtnjK7qbysN1BmIcvqY20duoeyjdYy0OYARnDu8iYB5Lh
sN4y+RRkOztprbeUTm/GeksSycdSK9Ogc7g2wAmignCYOKgUv/zCe239NAToNfnOeApNtl3IUM/h
lCzukJ52LE6LXc0bcGZGfX3F3KlWwe+JskcPeU+VuprhphNeoPkqAC02ClId0NK0Y+yFlLaXENYg
DKhL9m5EA8BwJX1qD+Z8aOpaWnIanBSkXTEohIe2udm56cAddr5OCdXd9NPqbNZx9ngNgqtMILjO
UCkNt23GwEczOLkGYKlszhd3tSRe0t05KfIlv+sR04qks/lmncczxzeDvUWcrPcrTCNB2oazPEkb
/jSKn7BhjnasvNNcKKaSNqHtDtO8bCiMMUgIRPammYt1q/eaCqTsDXWU4lZpDTOhQFRO+ruoAKdK
kbwRPfIglZHOU5aD05F3LBPMrf0fSToi0w/2iznx7hdrKiLaaxFool45y+bxW+1mYL/XYkjdqFBI
eSigGRJgVNgNmzEGYfCW43pTHdMmAZUKBZfrsJXjdT1/j0/nKjt8OfFukZG8ilSjW6+p8sweIUsp
jNi8scBk0mBqYCSFpj9Cm8WSicchdnmxZSWonGMDNxJ0/v7U4FtjXcYRNstANUUHVdCB1p4fBPlJ
ezITTZzXnA5DNx2RvM0vOuuidzUPnVd3+GLDqsiEfmpIdvm2snV+9C87r9fRQ0gAL8XsweDEni3u
XJWyGIs3FKtNYbuoPz97aNDvUDofrs7+Uyx+AswdIki10IJhOD/WTk1ZnZl2JhwCI4O0SC2AH3sx
PAd2oCv13VQAU5HaGNRo/QCXo1Wn0XLQYdOx1rEo9+kzLD80q8O9YhlKKBngPv7dXlLpj9noYzsu
mjDf9xXMQCvBSXfizkssTtQkymjBRvV1YYAdOalutZ80gIf8egJ/Fo3mJiPCBxoyQHGV361y+Flh
DlpB0kelpuzwizloZ36ljfpXJn1a1dOp76z0Y/fnPacZqlJjpPnxl+gHSVrX1l4kVsd2XUpukCkC
b5jD4lJC+6fmhSP5i+j68nRWfL4U8qJongYheWxF07hzdZFYfQwwj7ykyQvJEzCqRoO3Po0ZBiAi
knzeqCUdY+ta2PMTE3bQpPU/QiJCIoNFeanT4pNovXQAkXLSU0O0La/7FV5giGSG0Ees9l1y7OWC
0Sj+Xxl5EFvyy9qZb8NX3u4/dVufvT/b6aldnmlyzwXpFJj85Q6VGYNwM+J2ZLSXCiD0WU8dW/WQ
zjytKmfFMhgkbV13n7sxoyny8m7e2FHeCp2JB8DilP5Dm2yVFt2ojsbGLkChDVUFZzUE/M/4xOSs
n9oZBGsizPLGugiqt3rQC0mXmpN1CjbyZ+T+fbggLB09H6LkG/YdGe4Po3Fh9suc89yC3DETgSP9
faIaUeQl3swcv+sA2CEaQyR1tLZY/YGCM/3E5jwoq0zoo406VA6U7hyhhYjbduHEznvhvnT3lAjG
iXkMpv2cR+N1Ub3hlFdq/5dM+SkTTob5AX/F6xGV2SG2uYwLD5nbzxQASBmvbIrMmkx8H1QqfuYU
OYEfrECo8ueNgMMXavfn0xfvzHswuSuvNF40SDjuQoExUY2OpcTR/+3GI3l4xwE6009s2ptqMmK8
wQCZrKXdvyhkr49gvhU57oNWiQhbTYlGggunWSCaB/s90KlgWhKdlEwzmrRjhe/h1F44a+iMnpgf
QHJd9UMFDMVqVy0WxphMqqMVN5gOS58r9IUwLSZSej3UrvKCZ+nAJhvUg77h3B9KkigIBvO04Jsc
tCWAXUdfX+hEWbvDauh6fYG6AcyHFFmEBPSGjQbbatFpv5jfaDGIDyg9dx92jw+n8A1KoPZxnacY
eCFmSvHeHl4dla+00oQTzHLFc9mdWSQm3S3tfFw04uHQe0//PFlKtyvDn4dZudpTArR8W/fDaD+h
3gT9adGQNBiZlVJX5KxH+HWykOsDjdN7e8xCrUUMMXva620qIyVuPLuh3UkvuRAn0pab4kDFv/xW
CoiHJ5gmKmNW+IR9ha3/dF2HrnicEZ5nf/UsOVh2e8SucRb8Qmf80cltuM5MyKkZGsxJTvKm5vrs
Ld/j7ymQxR5YaJqEsvuPR4/IojFleQ4CQQbkpratFz0qEWML/MNCl1c6QUI10MXeHUclAocomp3f
94lGfJQsbYF8yyXxzGZo0AMwVhBx6UUrrVISlqGRVKmrWzVfHRhcQwEi2wi1csRb2KMrOXxZr3hU
ckDqEo02ZnucBfRXJqriboUb53pV2j2+s/SkGUTbG1/jDplvXO+5Dauo+qd06gLclb4BKcDH7URI
q4JBsGERdBrIXMpvgN264jCaZZ4pKXi1CU3RtMQBBbxQOEWsJ4I9jQB+ZIlpl/MM5E9PllQaAfd6
3Uw4VViZUCG7ik/rHgZDRR8OEdffqMSTVptVxQAdMtSsSIAfrbbmsT9vtkGFk6hNZs0kcyr9er/U
MbL1G7zcARhstsQQvSO+Ngw6LW86OIoOERjP0X9VUzJNEoE3Yui+W/mvqNj9xyTTgtgovjvTng5m
KCij8CauHexfMIwUl7rOf1XvGwIji4dKdgp6F2cnRkIjpa4siL+PDfdxb5T+SsZ9Lculh1s58Wu3
EcCkkrAKw/fcBDXAC3TJnYTw7ou/BUHfU6FAeeO61KATXLTk8ZjzkIU87pmB48iG9wC5RDOLjJD2
BzL82EssM8mDmMnpKQsojGDsLVYh0q28dcHlSmGs5Dj9l4iIaiWRGZIyMSM01tMecPqUC6Lqlxfz
djnFdZNTwVQGni+8kVVxAlhZHRmzhasnVCvgFnrjHy2+cAwlUc+ScMUST6HQQnZpwkCgzom0FMkk
JwCtQjg1mfvNZ7TgKHvNNFyzQsrGuJQHU0lXelGj+oZ+93Cpcawt/ziTtL6N0g9QzY24qJg2Vk4/
LOjUZjpUJIrpvHKEYUqqGJkcUeLenbBFDkiIY0kmQJ+9SkD6UYJVO7l72Dx0amm0eRyweJHRQWnr
1Hvd5a/9Wb41Yjb37k6ghD9NlVO5/DmaUr7C92P6ovJYHKgcOKNK+6PZ4IpBPjHtzxZcIf1BugoL
IS3h6n7bgUkx8G2BE4pXvn1fOFFy4Tlwibsjayy1xruezlWfQ7ytO3ynrqykqxJ6YAE58iTrRwpG
fuEsWR8j/wCKjUK+Bnq6SkCpm97/Dca/PFaIuoMQp/XXip3mVSVJYolhTbmAb4yy3MZ8Vs4AKoUz
4yX3WHonA/I4ksCmYlGIovdHVQF/u/EiT7kf30ZHv1lLkkibv5O7/PxHMX3jYbAA1+1boPCpJb3a
YcbLu8F9qOQof9gsqQ7IY0RYWTnA7N/95P0aDgyRj8iNdX/+Bnux04U8Gd9necWJRgk/YuSxL4CX
99GWsM6CGzyPlUKfrq9KIzuAAHpJQKfeX0e8Yk3UAsm5NyawmIR9GZJsqT3thsgd9ec/JqjdnfMb
2XB1dgWUoNBYE14cQgBJ8ldCHppcSdY4cuvc9botUVG+EfloRDozLt3eJyCWMSdngWp9eie3+bZy
zjnfaIy5IyK5rvkKuHcmR3/fXqMjwncsx7Ss9tp7wzuopne1/A1+nLBg12avNQ/VUxDB+mQhP2QV
h9gT+vMJI60/zSHHINBFg0ES26AKPanPhI5xYlEAfrDUN5pFP1m2F+Mj0k87yLvOWYwW1PZbyRXU
Fw5mLvkrFrMcFFcuDK8jChy4gd8jM+BTTWzXDqyO1gCMTmwrSpyH2/1mlJze6xlaJDIaA4mvdZLu
j+kLuKmMFKsJPeKFzwNRHXFLuc4Pk8CyAGMegArHLOgVvutee8EspMRbt71PoRvjPGL+lXiI09Jw
jCMbjoSNbTjkcFDCvPR1osY3T63/oxcqe609B04oPJKvAX6z9b1bCeGSuONjD7/ANmVnEXX8QOqY
isyaiYj2kot18sodpp7v1j1qnr6hNf3hM9pfz1sdIo5S6VCnNzwGCCiU7a48PAEpCu0jWOZou2Mr
n7ANNxI/AoHcwSbN4EDJJcMOA54NT4phMs7hkuJIDgxzVQOVuFxQAACdLxvhpCSNTT8qn63VCBDS
r/zyciAD0asQWBrDEhw7yTMS0y+9ll6Sib+VE93MsmGJyLLmWME5c69ViOe3hMF/8p4upYjOQHRV
7YRbBFTNL8rQJIItJvHd+kC4sCaTUuOYlFw8y5UOC+ophCl+Jb3GdpQPk+OSscbx1Qc6CRAsNbN/
Uq2tbTWCRsOsUnZwAuBBRuGB3Uuqu1UlmlSOyCcQTFp3VOJ/OCpX2FTg1lAtRQ3MqifC9DA2ApXX
jDyLxF72JKourrVhqsMykmxs/dis/fP+C2EOJvsIPmMsmgB0Gzp1yJO318rpKR3e7PIBvKSk+0PH
yncJ11KNoC9TBlxkzmB4U6Q804YGC/3I4EDa7E6awuI4pQQXKGVzEPZYSQK2QOj7EUcWPd/w5dwy
NxloD74QLUvsna35Bmlmzk0/wfI0HM/7ekdPeahdTnEr5/oZ6Mm5MyVUlpkPmPFSwOevfBft1NN1
6vFycekNxHMvo2oXAn1PXvnIDOHtOXMRgxdhbrwwWjLuisWsByvpwa6d3THW6CzyVMBDqNimnY+S
k/zy6f8HDqgLMuni26u9aBAO/PooXsaD50gKxcUQqw11MujOfY+FitW6HKuAgrVvIYLQdm4m9MZj
uw6RLOg1/EprrGUV5lCUzwumtZV93g30gFTuy+jcorSOHl+1x9fCDUEl+gzBDCNlQZMK/kyF2vOr
YXPvoCq1PaF9/6gmnu3SjD7vH5/4H5092z6d+cKEivb/43BUQHNLAdU5yjd9ghv/NSQ4PSEi6d85
T/mU1O4gEMuoTbs+cfSUdHd15C9Bf+UpknMaWBzCMkmIiZ6coEDnXI4matn6Tm9E3xQ6CjpTi+dt
RrevvjErIsN9sT0bQCayH1c8dsUNAbSaY8u5oI/WulAo1K2j8ujZYphHcyN+jl8uDX65RbTxRZaA
yLgu+DPMOyxa3rYe5p5zPYrmhbFyjWydv3rrn5S5+WqDjmHeJwpP+E+ojIrGjiEztZ74xz7jt/Id
DSWWHAG6rAu5r0R8T2s/S4fnk5alX8EQMwRaAB/Kay83Sbvwq/+CuD/KgDNtzX7YgchH0/83vBJo
PCP5nwkdid8xrakmleJPH38dYDdxEjV+6WO2Uundf6Q28TNCfwKqu7J48DQ7A62gToD+qP7fS5Ej
vAPLLYBLtmqO8gKHf54kCrhmq3fpx7wBLB8JHKfmpplJc9eOO+ydZns1B/vBR/vx8JQWPsGNYYOh
CMpiTo3KgVM76zZSmYCnYH0EzHly793sbMSXduYRx5q/jbnD5+A5jLsSxLW6xk292LnykUj7F5Fl
MvvyCu44MHfL3MaAwn7Fn9PPYHVPDurgk14+cBxlehvJZRZXCih53AKgBipA2eN3RUxz5MCSDiWi
phacT+m/u2PGE8WG7QNa+YXfDgFgVXvmb7Ba9CsudjB/txoj0Ft2UnuS1g8lcAcmq6U+xcpcYtD+
4jkBPE9quiXM6oASeUGlhGUOt4JXGk2KVES96PBPpOMRuW03wvLn9zbyf5Qpll8ouyB7IecCEaRO
fhqOrTa3cfhEKSi6+mwrbg8wKABthoitnDyzq7bqMdz1UqvTb9RsjtFtSr/Gyn9VIBeCBO04Zh7e
hUXoA2l29OA0OlMg9yDufOTEnaFu8AEPrGW06GKm0CSrmp7nILpXCsae3/0DlWinXL2FkmbJaetp
2UgcAUiaY0lnoulUVp+X5q+w6lyKMPFkoHPg99sdIAjXegk1CAz2mQ+upV3YEh3mPIhBhvtv+0SV
PjRw4adjd71OEhul0te95os1OjA5CZ9t0QayFrx0hMBZl+Xki6KMh/05OqV/mP+w49mfNk2HOMsp
42OMF8gL6AYUmhOSe58aMAHv9XWITT6m1thUo0H4Y7298THmIn8D9+UUZwf8+rhPRTGRVuwtCHJ3
TCN/hIYnE7rbC6+ecEaHFlaAqtyMw9XpccIOwtzTIBe8SnlRPc4i+dYTVJzSVyKhe6UgBZhOvSXJ
1OU+yTJeciZYvTd78IKvz/ljUz+bJNXMdcH3ayv5uK8270beTp1TQkjydC7gf22Qb8cIWAS9n54p
v6wWSaItAPWowRYdhaWSKcIcgSxs4NAUOL6xNsNrIpuOfbmyXeMSOQo1EuhbusuNqVjITFyksGkJ
2aiB/ARSI0R/PmAfUrXPbz2PS1i7jaJuY6z96TAt+ztX2veo4CfIqx26nCbieNAbbK56MrrgcPaf
/nkFYXVUEYe3ydMy+gvz2uQj5Sgzj5wBfUgOV2NMrxN6atB6DaMzJ8kp/i0Vw4dF8n//9Zk6RiVS
lo3Su/fzhGo00I1W1BWV6DOQ/W0fEKzIfnOas3QYsCOhREGDUn2w4SI3aDx3W+jbLK/k3z9kzrI9
RPWa1KXwQOz2J742jPmiyYrqYiJwgq+gYjJq4dwsrLNN2QDLUxu/8NaXkbFUpxRb3FAtNmtTbDlc
zi/eYb3sJ5J6bUmXFwTNWb/k9neSJwxP//pp5S35V06lJ1HGewqsTVnRuKigUxcn3VPswnZaembb
oVjExosJlq4whqyL7FhOU2Pt0F4UURCY/kEqFPdgcm06mRZGx/QXPY3vgRCbWthVJb/dwfV35U9d
/UXBQD9YGOdfyg8r87QYA2L94IVjxe0SyaML6HUKXDgx3ftzFOtiG3Ztpc6rkJGgVUNDp+wpg961
plVDNfdMyCZHuiMZTSDjHp8r75TVWTOhFvZsxIt+ZcPRgHA+06VZUhFnD7mmQg6JuqtRioyblCvr
D/STMi72w86xGnn7jp9HPJBJdtEU475ZaxCHpfkp9dCxpvgtI7D2kOWZ4I9kYmqAiwtN5PeML18Y
GMAkaI9+2fqMJXKtNkZo3HNBnpQQIQa6qqcOPB3+j1NzsqkPtfb2h6mupycyVRNgkZ4gqSnZ0Fit
3Fclzr/OLy6zQB5WjwEPsIXngTtXMYslWJ9T+5wAwhp9i4Jfjc477hVHA8XVUP10goOOytAEgDjR
XrSDKpXzlcNasKMJYsmZLdjwaAYvZa+UJa7IUGQXvmdScUshKw/revg2T833Tzj0Uo1TMy8WUHhg
4uo6zCy438O2uvafB5DViOdBnV0aH2jhFiub2DKAYv/mX50dAzkhde2Ixmk0dY0WbOCxSc3Aect4
msvn4+A9SFsAxarEr/acj4UL4+C+hci//06xMZCSN095acEfySJ8H9jbjjh3b3oIICLKt7OsZZHy
h0VthToIr1/SEX+07XbXA62RlCvWCN3puwqHhzF+c0Ka1AysaYW7cgCAA2/GvW0QpBZzySZHjq0T
IftS0P2heA90VrNzOg4n0InOCTyCrBu6+AbduKY1XVrUMfzJL3Gwbo2UASBwiBSeCS4Fu7Po7UQ/
h8+IEH/dck+2AJMdbd5Ja4UwwMVGqiJ/TQ8E/YkiivlAQ4Tui869VdCJhvQPoREWGWsD7E1baIVM
RG78RTyV+JNXqp5S7GaRGMsTDSkzQhrCcLnwvggk3EQLJk9GHpAV0x01xS/iAMNsRh03kmUBSh3h
B1SS9CvjQshKRq5xa+BVEZ8FHmk2Nha0vtxuljsvZnK+Jf6D7nRtFSsRQFfXYrEpbN8HcprkCAT6
bPH8Kv8zjVSVkpVTFT8j7u5PClUIh4b90h4b3uiNW3qTSTHYnkC4C244WR/xIZCzpCwmDK76AOBt
VEMy/KC4litJtSmHq6frO2t/8t92dypRik3ccot9SKtz4DIa9DP9HzhcfcPd3OmLLsV9wfWSDVMw
839J+15U4S0O89hAhy+84xgtvhfptSx03cIiW0SO7/i1ROdnUMhRBq9bKtNKpiIv2EzxOmZCzGk6
bX+Y5HZrC5IOwcUAVqbhKo6gCsFhZW6/XC+eLstE+6TtItk5ArLYT/XaD+TOCHt08jTruUOEB/VW
W9KxaZB99so2eFIPbbIM1fdtsMeqXxEmc6J7WEOpyi+3qSzFghESGmXrGDfBlNIoJf26YF6eWRq9
V2r64vzdNK9rtFgjfbyb9BQQcaHse5eVOmqkSon07FdWxCFXlgcQmCX8hIZur2nE9eJgR4xupx9A
hFs1D1LSINZN/mXFazfRlWSuJkevCvwagyXDgERYxCs/BLEx3z+komAGs9GO4Z8yhZmP868wIgy5
UvpdLCUaghI2kN0QOcCtwGuQMo1+7k8/ppR6+/KE43buIOTHLnTuef3bLOp/iuVKWPvMWdv5pxeA
0ca5jsf8TKEBHBeWO7ksOzG8r3uG8A82aeXd9SoWl69sqaXhZbJxwoKd99g6L4WokCHKrg/CxZSd
qeYyQiwD7ayw+oWNCvD0huOkzxVfpmS0Hc2j2Xn7DVs1uaEhrnZ4MeFsmLmBbyITMoO/eIkZkj8a
7y/GyKGBcN/hA3ynQZhF0sAdq+ppAmcuptHIiAlr3i2MSBPCp0QCINYXOVZQw3yDhi+LujiF1jEQ
flH/htMmAQT720aowtd1FNvSMnPz9K2PPc/iROXAwN2ta4ONta/cLR89jw+X1ryMe8pjl5hen3cF
Cn2+pbS+aERO8lFS8noTUQNCP4CSw0tAMJyrs/voqDRmlXt36lRKGQt3eTdVdllXopCh8m0Qh5ue
UFf7vXAJrL0EIKSz5gVT/FFrUasKMqS9FARM7szN9eH1W+yUPXEdWWDZ2y+XJXAEEGqfrqG1Mcwt
gz2cU7FyvLCj/NMvK6rJUMhrQglhZRXJjkZFkaxeS8H1SjntyzJfcQf/sdgM1gKfn+ZP3nvc5QoG
kWp9KH9uDs6bF4cMerU56MmFbvZ2skNFtsolKDdhMhKnScGVnMr5/xZdsUNlj+OrAipfMoNkN1Po
8V+Bqcw4W1FlJIlHUBtsNzcVNOYm+0m054HWp+5fCsmgeQWfUla20eYCjO989WBXpXlRMjm23S10
YbuSu40HseH9BFZGg8snO9oXfW7ztnJB5apITagesBCCXmXbHT8hBu1F+wuzQ2wnYMnPD5jSTLl/
55BdcjevhQq9b6DXvxNJLBNcuwrzYrlsk6vG674XfECR0x6anq/GmLxBw8R+PfpEHv4+njjYz64l
5GLkq1gCERV91FCZEeV6SdtlDGOgWY7XZ0qrRQcODvnT0nE//g/ZkxIWzlDsh2XLcnjVgMSTodxa
7x+5wIqii6VWRpJsdWKafzPN6ofALnXoCzl77isNM7ORu/4FnX0nzsNoJzUmmbht1BSm8HRJcUFS
yaJS83iJR/SeqJj5oUSbqHgbP7q5mJo/FDXCJdU1MoofqCZ4TuakYKHLH3qH3iv4eAZ3bgNcKWAQ
37s18aUJUXen5jLFEmszvAcTMT/ADLwXH9GsqPJnyHTT+sGzGqsG92S76fievf090idgFx3RUUU0
9fLb4LQu6mSumMDgTeUOO8drWHsTPbm2raCzolZ9nlnw355uAQtcxZgfqbXfZoZ0eq6YlVZpjwH9
LsazsBNxrcpMY8uqpNqFo/cQuHOvoWlwXob2aSPWa3ktsUttHnmPOtjbdWamO/ahUVZ65u7oiGeL
YFhckngsxAvW1XN/7ahxNhRakecqwamuroeqbqn2dNBKkE23/W16oSrcAlROqWZo3jsmJHLvhODZ
dEhiOzGQNrsYzreWHC76VW6hqZsAVHjx0LSHUjUtv0f5q6syi7fPzsRxm+dKNPCDOEzLC/Mv9T5l
Gq8V6g/PG3Q4LsqdNlcm7cq+q+XRA9jT7Bg0bf9IQeCRkwNDUZI/+gFfQ3Eq2NcjsjvxvhWbnDUS
2H3bXQFRxU8s8l5AzRHxVhQagFWfEp98Af38hpVY2nXQVAR3yO55kHUmqaz8Ob2zH/3h8Pw65qGk
onPmFAU4lIcEYgYK7YgqBhcLa7D5OJ3wjLdXusQY25duKFPqQk6y2L5uvHq3SuXhU1N2WvF0IMgg
z9umS03QfAsY+tfwSwAZZjY+M7DKhcxHI8cWBU5vnMkUkIzYtyd1CL2MCOwa7DWlznXvGzwNz2EP
8rCJs4kr8yOyMSCdkHh7Tn7ltxRayez25aTicQdpk1z4Hju0cpuB5RfSX6dHibQn/fohAowJDuIm
R79bsKiYs/SKjGk7SgN5hTyE30XCNepnfIFI3+gzWQ05c9eRKUXqzP9kG0aUsKvFb+r/P3rTIEpz
+iKBfUkPMAI/T6VArYnMXhMuu0rk11i34KAlCxrtbQp3FfE5gcewZDdA7ZxVj8EH45uZX5gP+TQ3
96ytJXUUzPuTsR1+vCSWJBMeZpl6BUznp/E8urNexmYz3Zh/6aMrz2A5lY8yQK2QuqFjSOIMts5d
mSH3IyGlK2jAimHxJPzbRkwGh2Jbv91oz3hGXsrDUzbR3Yrn4/pLTrtCxem8iNT0pKldbg6ESGiq
7F0D1jbW4aUImTTNaZ7NWRrBj9vZcdYYvp8zgM5b+siMmKhTQWowqTYqWfw8545yKm6WPwGpXwbt
eWb7VX7L+ESYT7DNyldaMxuYYiYFTmNTaKDC7XpgbosgDBU58tvhlme950k4s6My5X96kvBN07Ik
yFfKQBaGaZ/4qf/y88NDJ6krKbVSW1BpmsGG7D7xZXxkEBqwRwI6SKZilTH0WpIxLDpUAlPHBBTO
+Jv7EjVh2b1fUh4OqMGiQdoYwcE6m51qbSdJNUE2j9XPUzUolpgMWx2haahFYjE0XL64/BShWQ7I
wnxQ31JLL/aa9uvH21oDpD2rYoTBeh8DBTOHwau8P73afvV3KZyedonP3AgF0GWkRzwjF7UrJnnJ
tf/6Gaf46w96wJiUGt1uAc1ONrFy6YunIgqhFe5JicJLHbDkVAzSWlLSDxDdvx5JDGDomgeg/9xd
p7sFSnwluqNAyW5UPny+b7WI3OY4/eQXRGw01k3MzBAA9DvybLWOjsWlaX2T2G0mbtI7AxCS6iyB
MeHFHf/x4y846MP9wf1d8EzPkLIjZ8GXIYay2lNgIwRftasUlf662RPvYqVxqnM37YqbbB47Ugcc
8Uyqi+IqQ6mZWjMFYEdy4lBsqnyDrd78LTWJQwBZ46E5OEHarj6yTMP5UCGuuWfGK+x2yqlJZX0C
QWcZknunWxmv5+U1VkxiqMCfmiBtG2WkU1JyuPo2itHOSAz1Pb0ow8VRU583IdtahVZYjkfqsK6D
kROFtppQVtqosw8c4ALXbroQ/ms99xsIiWpbL7kvvkBO2yxN9LQVlsoSNP4y0qIAEIMc+p3y80mN
pS03aTyd4Sk68ddaRHtMairvtNWJYbje4pv7H49wZFQ/Ub8UqeRS+z7PJmxLSGc+J/m/8AYudRwq
khdggAiFVo0ZnIkphrbhRX55V4IWRIi/NvNDUUNVu0rCO/NHBVmDq5JHOFuvdNZDs8QNoVevR0bQ
Q0+O7H1+jHnXhbTyY4k3fK0FsrBBDqTRFXArW5l4g7Fk6nIWjPOS9uRIYQ35tEqDYlvxyt3qUBlz
UF0ov6IyMBpUduiFdZoZOVEL8pMQIlK52yJ6N2W1zT3k3ikeRb8CVGB+Ko4vomjZUyvYT8b9s9jT
PyWGhf+Ft/mkMVa9kzPcR7jqCQt07aIsC0WayrGzyqG0AjNMXhiMjtXJv7y1Gj+Z6gZDx6a84DLT
U1p/6IMKqG26z2lpxETYjnlYGo51HwoAeBpUPYIUPHZO4tc4/fTNFsyN+8bt4fKcFdTJYvmN0UpS
4OdQY98sl4husjPAmm1wJvKfsyRKPLB8cahFJN+c+nJ6NPKbOOfIy49F49IKQBQIymvJGtZ1g3hJ
anu8XnDxHolV7eKFhu7rYLvpc8n80iQFTb+R7Bt05OSRoRcmT3KOFqsDrGoOdQI9AASRw3DOh+5m
8MSAJ1g8k452mMvrLdBxpgrT4Z7wfuasIfQ9znexOXjXnaSothwir1YeEUTHGFuXZaudp0taQMpf
FOl5LQvYX/iFkJkXgar0dTgj3/XNkBlcnk7MErK97GKsqet9QCFp326h3UnKpahN29CX8RI+HmtF
8kYyAMgN04IXSrjbGJ8B+tU/C52IbSSDuEq8hJV13sg+VR/hfF2MPoc9frVkvYor99CoTI5XwYEs
m9HuwIsvcB8GURFI0TRerF+8CDbu5r//o4c8b2NIEqtsxmTHjnAUIIQ8PD8HyaTPNs/c+4zaiCJl
tAMvJ+jh1mtxc8/kn3aEOxN6SdMptuYE4gviVY6F5ovB4MU9DtP02T4cQl6aiiDRSDf5vTV4K8YX
DQHCxYvlE/tTMzv06WOZ4zwkSmeJgl89hslV0V+gvlzTtdVjgTLwv1bIfeEF8sSoykxuqmmJdFb4
Ftc3lo5QmTfdIpr2QUE1JHMrN3ay5ZsZa18YIomp2gC4beJkaOE9xQRf9mOKLtpwHwyKCc0dSLRp
e5zhRqnp/97+pibYAxQJcG7DgK6YfY+8X0/tUyRPoFmES6y1NFaDCCnHpfNoqAKrzYGlnk6mP4hl
RrFVu04P53N+RZRTXddkABPYLY1VwkfKZ690Y8hYRhukdz4rzoISKejsAiS/KVE6vXQnaweftMnb
yCUxuDyt67N0WCqUG417N3H9RvLVdvEg2QidBZjfcmNRRjUVBgqrDk6ru6him7yv9tycmS0tOVad
cjiWxedzWAd3gkIABavV+F2QKlKi2I8Mo89eG590cyEZ8AFyoHuhO7i2YYQGQsq4QiVuLk/TC+52
0iEP5LUZ3zHThjulpWM4++m9GY1JYKzlVqrqjhybewdFuXjZQi9bDwidwFKopqG8y4bXaEHGYck+
epcqkVvurTuc6jS10gOICWkvQLPPFMO3FKab2F3U1xPb1FXO4kIBQiuwaDlSTrzTU0Kd5YWgTMZM
cKCWe5Nd1eg7Ezb6SX15IM8r7f60Y2DcUi2/SsnV2zfvjmGCd8t49tfEW1cTQBDdPNefshoL/O7X
TwFPiZtHAs+NcHOELxtfg45xc0UewhyVcND5Qu0vfOFvNU4mtS3ewbQJ9AgqoSp8MVS+EiCSrtQ2
kegWpf6403jcUnHm9JvC2Rs8IE/m7w0Pcu8H631SR9Dr1mQE8oWmDG8sxILt+3hPelznMBITrV5r
xEoOgaRs4/WwbFWIf3L80ZkY5npzuqorarj+q3MV44M8sZAqi7GgCyj292zAwt9oRzksOU3IHVwO
dTFtd/QQx74wawU4I+Kv4hYM8QDooym8xhcTj1mpE7UFJJImDCoIUkcZEq8RwHYnjmyLDMKPz1pI
rKZQSqwrcrXv9WStPSvylOgnt/B0WkWV9cHffGanp49mFimDiA8eR9AklEN/7ox5iTfUgu15f8uP
UuiMbX223gZM5GBwbiREe+hyC/Qf3CH36SzR/BBIHkbM6e4KkLH0gvfDbZHNvRPjDxHe7LxgXY8Q
sD/FklwHWgYxz4PedGP3H32EIvsyFfF+c4ok5eqcFPLjRSVtZmLUt6amCr+RwFNP5gl7OCRWqCl7
1F3KpcCsQuQhQGthFC0NguO0vHJKIoED2wVUUKT7TJtMKaC1WqdhaLlMB0yH2Lo+aB5eHVIn7/ym
DG6QOHJTwypq8N3d4JGQxye2gfGm+1TLfqdzIYfRmofoleJ376QzM2N847a8OHePCG+ioVx1IMiZ
c/u/4nop540w3VITn4lrqHwtj407GBGAE1Tsb6t5KNMqiT7eiP4ncbu0S0bFHgHjZIAdt3pALEw+
SN23BE/wDY/GWh1Spdc8B2oy1yWoNfdEwatNG2PB0NxvAI4WE1yFwCz8mVpWpqcCjKfgG3zYICPR
qVneV9+VQJcQ4ui4aHE8Vga5PB0IScGZVQosZpr7jO6o17GkAdOgL/dE2p4wGo30YgoaBFS+RKgW
n/NJ0ZUYZf6RLuA04c6kwAIqBBMGEnRY11xfqZHUBJvhaK5KRsnuw/veeM44Yg25Lu/nNLo+kYZ9
joXqBUNOYraSMQk+Y8mfKvUOFsjN5EdOLIVthbPj/SsnEthWYZfpKpi4RxCkXmKE3GqZsaFTv22G
gXMe9GPY5hN1LekQE2YV9tbNj0mro9HauJzJayDdBzeJvOsZRh/Og+J3CH+SNz8Ud8UhQmfvdXbI
rvZC6w+mvn8C9NKfGevjz3IgUuCgHiUC1wEabP4CMcfIDYKCHb0ic+9I3+be2hvOJyaJIXUsJhB8
MS4Jij/gXYO+O6cC3nYaYCHfsjXrfjVQ3z1xaTancSAIVEoLuDR45B4M2ZMULkNoY3M8soxfV/NY
j9qyQdqiCt+3JwmCDOFxiJzSP/hCo9dZ8E1igggsWC6lHJvlQ5Ewy7DGJZyhnASaa6fgNERCcbi1
8/WDOCNzdTBfeg4G6/afzv2VqU0QxF2QWj8yfGRmkIjZcp5ZDsP1pSeUfj8AZdJrfgiqwh8M1n5f
CmilGt0cZ41qhwF4c8ymV26MW3lFeMMsb05HuZ44KUjsGbAeQ2adh7hRYr12fUlABXng4M9Xcr16
X/RvrKneSYXby+QSG+wopBa08mewddhF7UGGt9/5Zd/kYr5FJ65TbBJ/kTDh+9vKiShV3+eEpeM1
f0tD/pxvKttPxX2dH5jzRoaFXm8VL4/KPb/7F1Lp/IRGN0wMef7iFDPZ5Vme0U5Ov+QEFFZdw8S1
DDWa6g1RKMJaxtLmjIxV0OTfjyiFL1gqYZPostXQWcRMTCuSkw+rShREhCerNRF5wrV9cwJQwI6V
wkFFPR8++JW9O2QNfeWECNbCiJIqzM9iNOQtFvCUfjL/feGyjhAWe9H8E2YEwDGz5CbBykihD/SN
HFTYQxdjOOAJdqUTFHDDrbpb6sbiaaaqnNQc3q8uf7EP8yvDv+/Nq65KTLTNJEyH5EJt7JBne19a
umOTlvcZqXStWIUxm1LV1nUM7SiKDjTRQ32zkvPArci56wtUByRv3CG+R2oIxyY1NtuCKZG0UuMy
+9g5VLz+uteB2CSzE1PBtFGk/HsKG+jZABEWkFxFm3iaDs+FKDZg4peTniglmQbpI97+Yqh+hCp8
+V9MAwLBAB//gVpRRAKUPsbQ6xrqKop3zadCqfzJZcNd8qhv7r3iiKlasGdpXFsgjQtVYSvHTnai
MvsGKpMeXxmTeErd36h4tX23fFdfMNRJTGIy/gm6AILoq5nBaQ0aSmWhK3wCPR2wkZNiLwN2Zi6C
Xzwns8Ch3iTZaNI8Flzo8t+enWgIWIJUtFU67Wz+HXpMcaADwTJ/d03B93RvH5Us/W5EHapsf3Nj
GGhGNsA1Q2IIcwATpuoT71odJVpGkRVKpCsL7cHjFSdcqSkmD/p2KfsTzch6G1j8LmhQ8E5rZXDg
1KsnqHAFfhZtWtbAQfbOwAHtEj683+CskzDv49MT6DlrCukDpY+wLMp52IJeplC3zRpp+F7ETEsI
w9v8nxd/XmS3PcpdXZg/cLqe6rzBUlwtLET6pfXik/iBLLes9M5OwNe2ggoAJqhKryvlGFFpQNZu
cIR5IKkyeAclF5SZT6i7MjERSlQqHDxIiFyX1rZEUerFkBlM4LX+Jcc+4yaqndeaq04uY0UbZsEO
5MOnsgKfRPM3Gb1JarsKct4WR12mf7XOSLiiKgDfvaEDuYHGk5IhSEpfN2aTmmgTVicZhemIpi2N
S86a5L0WzGxkyBiRnlAQ/r41x2QkEil4pIInKxxY/0NMd2oaK0Lln9fZpwaB6gxkPcsuYPIVBUGb
j029Rj4ez8UvLvmqyby0DZjT27yz5oXRcXd8ty/9SZsPVdRQLAe9D25cJ5/8BR2DVq1kV+XGqPaf
L7ykpipRo/oR5mj28g4dAdmXFuSVdwzqOT00cxfO66pEf0cfwchGvAnh6JYaztdBhQjDO2vlvFrM
emp1Q0sqj5FfLv5q4LKyxq4lEKi/T3rhBgX2PSqpFbzmiMKO9LpfK2AHIO/pG+dBTtmmSHhBuMlJ
wmDvNf7pGvmkyRuPJEaRxQ/2sG3za/c4d2v2244IQqEgjP8WChYTtvMKjieejVx9daPt0mhosveM
UmTXq0dIX+HJo5GMw3RhpeWRKGpt1OTYBY0KaZ5YIBNwNT9HSq220q7Np+avqtHQExEnFsRzuXQT
cf9XfnkcOzY8ldqBx89exs39H7ImIirUopCq4+1NnhBi1yQucZa24oawBThNp4XJn7LHTTDtnygi
pbh+zs3yAdvIgbnb3vpkPcM6AZEA8oQ1t1VBmciv6xuPpyfpc1dWGC9ygACBzxSYRJrDOxMpUVLP
ogo/RiHycSwz8hcpirQa6Tf0EXv+zj0J06fHwlmg2kOUj6mIF78WHwM5593swi7FyEvpojo1FFOR
nmEekgbr00me1rVo3wMJ6R3LPP4huM0GXtA3lUMH7HwIHXgAXTWwzANllWKDxQbc3I6OkpMskVqk
m9U8pYWlRv4WMAMPxH/m9bz/wzH1878iFbpJeNtisTcwrnMXBZ48R8cMwKNDCkjlbMA0OAwhRm3b
RpiHm9XI65XLntkvfk5KSRd4d55MDByLdNfPOnoQ8wERMbBFfKBJqakJJshhkKsLczef7rTBegDC
zNKlYT/pUHUYh0GKeUHiX7MZvxdrnJtu91wV9vWvMbWlzvnxeRb98p6Fc7oS+in+mNtQB0eOSI0F
4u8K8kN8XsD2lt2UeU/5V2Wq7O4/Zu0V9KUmSuOHsN7xNg/pkU3ZprUX+p4R1L9GUlXBIl2FE7m4
kFJdkBn7HuF/APJy5RcT7BhFMwTkPlsCQj0feJFdIK9RBUh6kFikpBpqBk+ED4CAOFx+blwkT6Cx
/KVt+1iLTZfmZ6oCoMT5MJUpQfAHDQYySATvcZ17jSThnf2yEQnDLSnzX8rDcs/mnuvyY41r+rcO
bhr+seFCpJBqEPUiQQKJIKLKYif0h4mIZ35X+nqk392YDswcdHmVm0ugAt3SBZbvc44lSFZBuuAl
XJrzaOauLIOmV1d7mlcM1kkoLh4H735g5gSv5yBfakC6H/uDLlgZzaHr2+cC9ixk/BYzbCz1CQs7
4VIRLxf1P0rB79eUK+Y7gg1vCfPRUmbqJT9F1zbCEUqzZiyfh0lzrAEgin869O/RaSf0bTKQeZwP
BpJoDkKtb5YcIiRPygKqhonNbG+iVaHP/3iDyrJrVinfrJPZCogMfs1AxaZUjomZV6+/ySry2D1o
MUMkjWCUFztKLKEAr3o1MQktrWR7BGuTouei1oDr0lA2eZwCV8Xq3krC+Bq80qsSVjRxw0GmMGgL
FqsbHawKSw4sodtJvs4PR+tWU1xqd5wLZsJN86QemX1d7CNeZhoy2JVQhJ8eJHH7vswpFHk6XIOQ
H5L1egUe0ke/HD1mrihSK2JRjhkXIoFJS6tBh+F3jXfiyjmvSUSZ8xmROHm7Imsy8GW/CahBugj+
0/Ed3TB5soBOEte+SQ/dJMvXYCMoIlEBB/h1UtSgwm1afhNsJhMX/3U1knt3hADu3JdkH2W1FvYG
xWrn/tggIbjyKhZ4CHc9lQH7kUvbpAG2xNt2RJrSI/WlZkt3bJKRFH63bKIw5Qsj7ehgAdhknQp1
lSes7vd7R2kn1QrTJAkFH+DBSQZH8JLWSSflfJzr9hMyx7CocwbvOknOiCq9BQnlK34qFSTZ1VZ+
4h50iveWtECSJ+9f8kVVs5FgtfdZrITTcBLnwkl0vkgtHfBKBt5ohslRIt31dl5Y2wGTvcSXk3xq
6cNYdDu7X0DmBIVLZ36uk+zgSLkbOFTVa7vPgUgnmerfqykfSD7rL/2KiGrh9l7xTJcRO1dJH8O9
0tSEhK3AGm+RZq0hwJMe0wIdJsdk8mImCdsflBtEklv+r41Mk3RAr7Bt9ZY+ORGazllAixKCNMDE
N1IwQTXwXMc2f8R3lrI0p6AgtIc6acorUX9mLyQNA71r0S33C8nwt/CFTNQrNnvB3Ssxm4vpyxhI
Wf2NNYcVrhKty7j+EEmQBtHME0/pbjjzfwJ17hFBFIl7V9dPL7yVsT6WxwWQQzKPNFEo3FELcDF6
LskGFArCXMSIlRvLd2iYXj816INMgCvURklqxm9PHM3xSqh8h/CtXovT8DDuAYzMKj25xgUUKdT4
y0VmYem/DRQErV4VmbSu3fCbpq5ZeIXxuvE6W6CEhIda2U2aUXy34a6YVRPN7NW96hZggSGfmAzT
DvV3Z8YiRCkjp3lr7NyINbXWbrZPw39klQQwlwfT/WTLtv4rviO+7wrZWXuIys3OsxT44skPreUa
kaayKY/McX+DjI3X5H+HrTB3pag+G4poEzgc/pkgOpNqyUuo1BHspIZgvOaF8OrrrTmFa0oq4jiP
TDWJq6wEnzv2w2Kw7t41dw4pnZ8e+XuF9AdQGKF92eHEZpTZxRREmdSgKOp9ieE3fIYfwKqw3+xu
MIvJUEuK99f0aiZJnjMQiR7kMwmi8AWmWsrPIWDUA12KNwDotn+ZZljYUHiE4Ip94s3PTa69421E
xQAXvyDneHoWMHYOLqi9svScI2oYvcXTuSHAW+cvMtuDkm04gST31J6ICXq5XC6GSUj3bCl9Q+CX
v/rymEsRRj3+h5mIh+bVdDpxNs0YPNZK0RhfmdRDkNgOG9RX9j4mwrvQcIBrdbwQ8Xo23zrL3AoJ
1vaqzrwxIsk1a30FuWHGFAAOuRlKpEb0aHbeeFHNNIRAPNmm3G0fAmMRoPOmAfpQsR86OPeAUM1V
cVW2Lr/CJvmIK3b0LRmEr/5HHGceV+dtMeST8hQlHuYr0WINAMC1iIoIaTbl7QWVgQwpfIl6L1rW
wtGHRXdshfVbKJ0XTfk5W1HZtjXVAM9tmsI4PNv5/57ZR+RRTaHgyVVq9Xdqdhy1Cl9jaUmkckSb
wm9dIKiBwuWYw50nkqHghNmP3cNhu7Xict9JFUOarMZpEUG3SaCzJIcMbQKD+A+zd1olcxclSUlB
WvvGnNjDRVF2cJ+nCBCM4ZOe4oEDMBrZtdwFfrH2t9rt/X0wF0NQam/z+4nn1EethQ8mfrV5e524
etEnEg/BrcUpsm2FigciKkdQmoGXTdkJLpeHe4hn6c7t4neUPlQEAd9bW4TVu5n0oiuQQMTFSQdB
GUTCmst+/T82xz1G2SPt8U/akEu8Ne6fNj5o8VcnNZDSnr5VMt2Nqyg+UJmBOF+hYbRH1Qt1PAyt
SaoSYU6iOqLNcwqH8wdboDWiLu+q5ur8cnt20tDscqsYuCSDDjxbiBdvV3oXXX89WhtkTWUW6+8C
ZW1bn3MGl7l9dHrM8Ug6FNvQaCnau+rEZBcGN3ESv9wio3WNze7X3FvJ9IVJKTaYNPkEUpwxtnYM
k0n3G+xst65/cOPc5B6xr4SQZPxddVuHdi1UeGpkML3wr0U0awXl0ZjP4E+rza0H/oFWTEp3e5s+
Oa10zzCtUHZFHr9ywgadykaUOonwiPiKyOHqWWyEXapOBwV/i3a5y0w1WHZcyUNBfcT2QBkJ1pAK
keSGtzhEVn8wF8I7CA4f0bkZ8CZZvz2SFF8FNBWL5MR08E8hNUyXE2AC8SNJmFm6FQJilS7TeU7f
Iuo7J5h81c8ro3Ha+0woJW0sB+nz/n3o+EbMEFs6j5x9mykPvIbBf23BImE+Aove2/yx4KdOsXEc
fKPZw5HPmSMbYv5AOJZP/X+ZDLp5tYa6Q9MOrcsWc4qF1O7XG6hDChRccb2wflXAhj3tpBZ4u04U
OGjUPwNQgU7HNOgfsqvMnuinm8In7ohOFDtbxG9t/JhZLDAzdd0burWi372Et9gocgqDwKg0hw4E
CGgYNY+xxIxvktE5ALNWwwcQA0k74dDLh02i+WEMa6ehKd2o57qWc4TrqTlQ1+1PXcP3UyqKZxh4
zmwX7psqqP3SqlnhZYET28ieZZGzFdzPT/EYQUekmqt3hcFy5awn9qgbKXGNHXe6N3POYOn1sKOr
CtI+10xxl3zem08OarKbDkUT2xruz68wGnQcrsGbFzPGVuEWARxOeX3kJyMtBFyxfdMASdMhda+z
NcH/3CJyUHQTDW5ojvE0UpyK6XX28O+IKrmNV8V7tbRK9oRt2MF2I1NQjnCs0kb7wf4g+dApLKmc
LkrkQG+VxNzJyU9KyU1u3OcWsLgaNfaDxVuJFnS+LR0n9dNmnCegWhU6W/pewweAlPSZ6M95OuoF
FCb/f6tNw2ct48H6ed00p4DuVjRaZ0KGJKCBKQujShojr8erjrhtfz6cUaxzjfCDpoclU1OZaCcd
ecY+YUPRI5u2N5eBjb9rO5z5snkCXUbuQf1V491ab7BbOazaqhtHgTOVlMPe1+pAX9t74gvh5ncu
F/BbBqalmBtbKCkpZiDlIKd1w6F9f1sMQkeX2Rxg8dDCIlI+dUNjGiNZJmJR9OaQ7AKqYHHJZVjN
RM+hHg2jaxu2NAg0PuJ0ftS5+jAVJfNlQkcgdTxJjhbXYWfxZz2lYXmwh1fqe7RjU+Hj4zhHWHdO
uCNuTtsSswgQkudjMmVzCkklBwakKXSHtbMTUwzlkiScvsLdLZPEo7lAUhjWqcA7KtLFaMaC2VDd
yQTVghkPJ/GB4h2IxrZtzGeIKnUaDHJ4IqActry1GRhGzaheeF3Hi9vDJ/FaRbikWnVj4YWKcQ5T
97tz2ddW47E787+2KcibPLHvdf6n9B5o5dF1JZS+abDVSVIp17MZTidldrwsNm/83BrHIUeZS4mj
V+Xvklc4w6ie/TMW6d7AWvN6J+yMdVkDE5VgLnPxrWBQgo8JKExGFlN2gDQ4snI/dYSG6QQiI69w
a7O6OfR5qTgvX9NnxnZL8wykwP94PZQgjzWN1cEqy5yhj5rQydFXrf6+wvWMJKOLAmoHd+Ky+RLO
D4TwjGTS346/E4ZsoWqltokEpNbwuXUA3cHTGpm3aDWvHc/9Ydv1UhjZMk5/NDl0zp0Nko1uHNmA
C8p+vWreVveA0T64Okh07MQl2JHnoY40Z1f3cFLc8n5vqMPQuAeADph/qz9g3S2xLl8qOxMZvzo3
z1gXP1n/kftmK6o1U40PG8ZqMvg/0r61qEx4oCLd0ooAfFqwmMT4qM0Zgb0wPxrY+G6ez9hl5/Fn
7UIryUh6pKkB05Jdcc2Dj4GY3MJTElEmkOuq7VB2DLa0lbssgzE2wonpFXTbmwRRc3KW1iMYFr3g
6csvEi0GAnjsFtYKuWpBiEY+fiTe5nRyJ14Lo3nWR2k0rH4e9zRq4HHWjrGz086vihs9NRXql/gn
caSdqQWUKD8PRSHvVn/y+X+JEn02CUac6vRnhCDccBeWfonhCI1/4rNobZ0yOm9PYdt3WGXnMwZu
xIGG9W8EBjH8zFKddD+5Pcxrj9TTdguFTjXxkYI5JNAVq/aP1MbsGuomvRJ7RZVKbtREvQGeljl/
hS1iFO5YtSFDDf4i8AubW5LQh1MeTauOgsjL5zYY3BFuU8yq8WqARotX6tRr5xbwcDm6oa7zzvvR
fWrj+sNi2TPpy27v+jzr/EXkQbe/lSbM7N4jbrwR9uiKv/3PUPlI8CatXyddam/yOmwkBK0uSxXs
U5AlWFsBc7f5ULzV6gNF0nfqWLfDi0WDxHB+vviJNw4WlTgJ8zKaPQj5IrNBHShmXypdVibxyYY0
9q/vA19jQglub6Vla1mnMIBV9EdGbPR40oT1dZ3/9szRrAXor2tesc8GhgnOlEngyO5/ebGmlpjY
MK1uVMs/1KaNLAPy4jgQ6S0h+vNJaTrYh/VEC0Ht7RZmYsqe+78ehqOGmm2GnMX4C64jUb6dg5b6
zmAvETb7Sd1VLXU8ri7qorkdDKxH6atlDClas9SiViKV21cbCyGb1hTYpmabJ70usLI8C70p/rdh
NO9sRDiYTreIJZzjof2ZbWXIXo3ExYBQyQjWakJA5Beg7q5Njj//pRxOKCjkqKOYtwLv7g4pwHVB
wzBPf8EyVW08pTDNCFDM8XnGLMKPcLO5FrsJTvB5EVL7PmGqI4mRLDzndPG/mloWTeksP3DuwwnN
NIyh4wLIPH1YlAkxKepfDTDBa3huk4yBj3A/AIbMOUU4Zm4x8Tth5QFVt0OW1EPmsf8cYfC3Fdv+
RbFuM8FWyuLiITwZOOntpekANtHiGoo3QS7MIQFKCNSXOr8vwk0ToC8eTBH1AMdirW8PpqZyUA80
Bkgv3nXJbV9dFJ88Gwu38rdCw4k7YBq6k80Vrb6YRlM8skzvujok/ZD4qqLurR3Uv0GtC+mtP/Nw
S6e69LYi4GxDEkjfA4WUOQXgbOlug3un5KIWNhmT5tpKcowWn362MWSesoH9gTk4Kc+CUJ2RlFPd
5D4Sn2fWBFXdjYbu6fw5qtQgZpfk1LYkPS+Q6mQiTRDRzAbAp8foDsDvGQfWe/HY5HB9t/eIjiOv
BIClWNqEt+DKgMLCxeMnR7ovHBzbD1WHv+0U9Z745BqDNM4WqFzwMO5BEY+v6Q+ro5bpR3b2tHUs
UbdWg3RCgjh3qhUM6D/5pliQMQ3iGOD6WwIr49dszhOzVsFsADH9qz6YfgFWO32tSApUu2BSCYoq
3ORkV2lONKGZb7OyD5CBqqBx8CXrViocrhRT9EELRUT1fGkVY187cEiblFLyE4Yw4KOoolzpyRUb
x+sTZnW/YntJclPbVyv4PHXxMvTzfgb5wKgS91ECvCtpuQLtB3iRn8HlrFztJ/xHQVd2k7yPn+2u
KV7SVWut60lJLbzd92c8JOsXwL4Rum2smrwR35wwfQMMV8wq0MEqIRs1YveSETmY435c8pRJFyqK
B1Skr0pUfnS6HXZ2ZF1d25/Znr3Kn4+wmJg+uqkW9cFtCKBkKdVVhXppvC8/ZaiB88Xg2+/I5At+
nsFcv5M5xvzF5b2k+9a9R9SqeqKalK0yCL7Ux/6v1VcDU1aMAPyfYAkGvVGHtmH0jCvk8V9L2o6t
7Mucv0I0Ms5+ZKQQFalJY7TVl1NTOAJtogRfB4AmMQJQJtc72fcA1wgFtoAOfL5sCbmUVDNBDpNw
Aw8txBN+UAU6ci//lHpgQ2J4YlfzJp6Ui0FSMh6jKMBaLYFyCoV6T0/289ApNHEWyMdHN668xk9P
Yb/p4zvhAk4I4A8ybjInMLAOBdauw0sFLPD2T+YICp8R0Xm+wYsa0IipwUckCyHsEQKEVRLBOVAX
hdLYZGWCQfZXlYjoXNcNmShVHCjnv0BqL3u6BShvmRyTWQ2UKg/DE17wUDg2cxGp7fNGWnWAl9pz
EUeecpJdj8Fe+tD3Q7RkdXYmECx3mC9RLLgL/cyZ6sgL7cpfkaBtp2K1bEvaTnOAp2abQyIp7A5E
Gm2a3xwnRVkkRmeRUjrn9ZgSnfgRzkcx+PnSBqRh4ZhWbr68OmFWMcsQ9E8lxdlmYLjjfqHwL1xs
FnR92VyvZ20iTipGILiWRug0kabhNIwOX0TOYahta+5PM/WNKf3Il9XaEzTMH/XVxTfXAB0QyvWk
ZBnK5zpgVhmMWwlJ8TOK/jIPoEkWe+vofNl3w9p5tIe4JvQUcGhwYDsrTUMqHiQYXwW8hkn0uIP5
L/3GYUBYASE37za3wPrtb5DfcTwK5+NAkLUxs3VU5NwDjk6SmcCEiuOgrco4xT/uaGxUBSxB6K2h
Cs6ECLniH2JefK0r3Kitm3lrQt/inzDnRtiT7rba6tsOKd297fWY4Jysa0MIs1ZkowjMoXodY1OG
oYUSVA9BBX1uuMA1X9XorRdTW+dywr7JEvdm9o8lCFZmmYWyzjoLB2EApDAG+94cl6e6rg/9FHYc
7WyaTZmI3zarOCwFStKGjdSEQskO87gzV9Q71RQxzERuSnIqBtK0TpBwIfzHB814CpgRgzEy31NL
rkWvHnlXAHLDp/r4VHtSmDoHYc/3A9aW6UI8tNeWs3+NcPhhE1wXWXaO64pbinMHRSo9r9h2aU/4
ZHOvqrXoZgswe7ckSQXUS4KF0z4jdSbKmKu7Q+K6IOVqzKvRtt96mQIzWmFWMJlEgTFzsfejfxbY
GyALDix7M3gUfw/bLboQhLkmeQns4iggbC4v9c49T/kmd6K3wmQYzst1LpnBvfp7RAF+qXqkiWuM
7Fd/eznHUe7GZU0gauTTaz4o88HRrmOhitPubp72j5LulMlIYbx8MYVrtuSAvd0YQVl36cQAJnSW
Ih9BRP+1sITaWkOu64g42a1AMLwVfQmrq94Ug9vGRGkgemCsxuIrON00zLhO9qS4h1HSCBGmWqT3
9HsImERBcizku9iXIpP3fFdTQnAilZYaL2umfJkE5enSkZPjQES6saWDY2hJYmia9uX4fAC1/Vd/
ZRds8YT2lA6fSvbxA1dR5EIi8gJyVpfOJ/VGc83f4DpW5YM3opzQX92xXLsVvOh2IgO7RI2KY1o7
dnLbLpPZyDl5lx7rZgPPbc3Zk8HJWJVrcCXOUvSVnBVb5k8MW9Obt9VE+JeBawygYKTAzKB1WxXt
sF9ZecpsLp8DOR7LLauux3gMswpKqSM+cl6GMI7bBNPft+TJdp6IERcXJG5JPadvbOUEycVLUN5p
7gbEmSNQ4Qz0wxplgq6QguieSmAMKhS5uA1fOzy+6ZQTfwV6Pv+uA+DrqFGI1tYFyhiOQzL+SrO6
gigaAjgXXh21XynhzBabEJGrQE24w/vntQTpw1l/33oroXUU2bc4k/npslG1hydFSmuiVpqGtn5O
VyqbstH9pUFWKvNJbpGEVP7NCh0jybNgHfWwb9G8u1ET355hlWWNb43VZMmed5vnD64ogdPDSWf6
hpAiiS3iUXWXRSgQT3dOS4QcQafUdabEXcDSGHvNNKWKkSZig90BPU6ZTF6lg+8PeqrQFKKEbY8g
KvCtE4PjrcEg6p2fRx1+kSKfjPpfiucq1n4RNP6l8j4veBPjK0qR4KjFb37AJDX+W/gr82I4cgWv
7o/JUj12ZTrd4vr/A39vSx6XO+hYWs8tmSizmXDnfFvD7Wb3PU8GwHBnX5Onv5KhHAlser1X28Je
S/ndOXqTpGNMIfH99H1Cqj4GLbnZUtRLbd60f5XwvLnaYjPFRKFLyT3T+Gh0pnrF94MYKpxuuWrH
orT6R7CcxZGeSDi7fpZtWvStuzPWhU5QaDQC6gJrFb+PGrnlXPtkJRC5GP968sq+3acHAkBlZqoF
rIBmivixrT96pilpovvOlIr7SsWqYt8huvluaUwYv8zvda2ld9Oaok6pXrszwPzHJb9cI9EuZQQC
1mOUagTSipYgBoi+Jd/GC/h2KPMjMRGwNSSSfUhtZydXcMBBF04Azypd6xg0zZ3h678WnwjEHsMX
bcMhl8RJPmAWr4q9Cie1SEu7PCkf3/wpMpkL9O5Yea1rWtmv/dCUE4dQq/ij+W2G7SWlXz3OO9Wv
8Oz/BcLC9f7q78fMgx+G5NSEx4SSHlUoekCBCaoqENMIamCvySm/TXwzkAhc/cgK7rgxiU+R6bDY
cXK4DQKka/LKNGYFAJCn1Hss+Npu1cmjtw8iV33EZgRoMcj0AnPOXXh3+Wvd7iKMtwAU3knrviaQ
XyVWfb5sqAoBiVetoUid2WdqmJM2qRhxxom1vGr2iKokpGGfZjklZQvmfyON5BIDiQxJzCbRRvlI
tqVWiVag+eYQajgrvjx9OrZDvruQefAJAl89ApcUfICacT+8RCPpfMXJbHq2HRSQnI+/eCDf2DqI
BEXNJ9MO02S5CAIlpV/M9LHyYg3gy4yKD3qMyqV+2LOIMstR8Z8BEWB3PBvnaFqSeFIEFqpt6C1p
IzlsTojUfv9txvW1LszxTS+8F8IBg9Eru7FAmnP2P9odlnVXAVZWJcHZsHFR6+a5B2jmyag7ajTh
JhqCa3We4M1rr/bz9pVr7FR+ReTe1Hy+7ZQsH2TUFeo5fVZFy1SUnzKVxXZPV/Uc7Y+AokmGusHJ
F8IjsjQ3EWGfwwbBSn4fNfPqwYZRHFTCEZa3NexRKr+1cWhkcGjxu1ApvvmuSw8vPUUid1wkfooN
UVe7G4/UUTGY2EKIfmV7KJJa6btc8K8iTwUs2rhalICIggvxIX+GF+kpvIzukKKCNm6tl1EHj92G
qH4SEfebM9sOvF450AJ6BhlYh2WSf043CNukt/biHTZjOKgaBx0VVlE0thkV+aaI1L1R744a9OMl
zUcZxjcunbzAXiCjX836FsP66Ja6T4ZtO7zxCOLf8BIUNyJbeOFY9Rwnf2xvGS7LlFtDTwl5raJy
T42H94nd6C9ODE5igQmH98BxmU6vvGcLFh+NNZYqtNbSl0cSd1WKZA/TLp2Bg98AaoZdmv0TNE2m
T0hml68Dy1bJS6OtxS5aDPrndm95htG/1JCN1RRE6h0Wtjr6rvLMBYjqPRzKOvQRXir30iq8Eh6u
YZ59aN3B3imL5eb6ZYrAc8LswU0AuSBQZOSnx08S694QGn0VBOAcmExIZJ3cC71s/wj/JydcWxpk
T9b83Ri5c/MA1rmg7yhu0clE7JDg60ANv/0oFYgT9rKwsjifgCUK6Ek2cMCzKUAuCVX/rVDgVzFb
uDndxzG5pzlCIc2Gg1hHMUJj8RaEK1ZwEXiFHAoe8Wjr1HGTFMX+av+w7Q0q6D68iVMCZI87JruJ
orVxQ39aL+uX6xW5tYLu5GpOVmgqfhyXyS/r2lmKH0E3SaFCRQgE29RT3PkrAzJ0RXwT/Eh1eRCX
A8n81ufxnFvy9nsoixT+sA48yUYKZpQAF+mM9g/Ab5pMgjq//W8z0OY0naokD2G91Ge/ml+A6xUo
0JoMN7IsvSs5hrtRkoIfeV6ED0ouSKPO77ZiV6O5mZgHEBhVkklUnCHcu4pTvXuwBLSO8iFmMb7+
/iZiDGsu5qjYLhZ1S8XEzBeEbap1hlqcpm2uLkQETtYMOqOotQWdMfshmoczxYwCbrdzAbsS5cjJ
y0w3M4CnO891Iggytp7dz3x9HP8dRa+jnNfoA5Z9CL6Zdzz82ULQesrFqHZ2RHT1lIOBcXFcbosZ
13HtEANlG0cddhRJqh9qVu7q2av9ptW0mHUR49d3z/ypDwT7wvrXaIGlViyH8EE7Ko6bdS+kJg8V
z4S3Q1jPirKDxU7pHKwjWc5faQZkJCma4WnQp3tCvZi1qreRO/6FewuQiErbwcSCt0KFdhcVAcaA
ZFUn7h5U5g7ypzR8j6ytve12uQvEvGuqadX/90C+/Gbv4+Rm1KzuQQ17suGI7HKNOYk/HHs3vFsS
7BHK7kAdKpIfmNLfA5XmWnhm0+ItTrzKpHAl8W8NmKhVuTZK0j8LRelxwV23kBmwmn8RKUD7ByAM
vPYAic33filORWY9E4YleBnZetCx8OmM06RampUHEbvYCgdstyXFvxg+fpIwjDGZZHt9DR5LoutK
qoUn/fQGLlP0d8/jQ26TsQs35mrJHT+9fPiXUnLie8LRxsJPmYZ0Ta8cE3eSKO9kMaSqDKxuDIK2
WCXEYN5qS+TMTzXBua8WD6bguOZVDCRpSpzvhu7lIkLMJDIJpgm7XctpVJB/vicxK+vLNnpsUkSE
kgsI/ujd0sZjMmC7wveiQnJ7WmDp21/CpR+s+wcqKLyILmJniymZRmLsEaeuG45JCieFgs5bnDy1
1fxuEmk0Y48aCm3h0o8yZgP87phd9ME5fui5/gsMLdIPIGcAo+3PJw2nJaF5OHukLFraiRhPoxsE
D0qlbJGwedWCqxVKgGXLcTY0O9xCkS+/39pWBffSEX+yjQTEYlAvsfsyFoHi59cEHitwX+KT0YIJ
5F+cHYTGV366rKwNy4piQk7lezj7HvW6wm6McU5hGPntRAFbnmOqS4FHZQiSdGSZdx3skfJI3H+p
SRRpUz3VnQ/dyp1mq/68L8L1nb0RHXEl5LlZ/PfVtEeGT5acSAx/bKPcVgMzCOMB4S3kZ/Bb501x
rZODdcjKMX20s6jy9QX6Rdw3nwMrP6u8p9TiRCOZfU+IZpF6KM8qPDZqimDcyKYNIJf56vtqllrk
vQya1D/IDXPozta1tS5Wt1Xtm1FFxzlc4+UOqb+T9XI/wMSiMUP+c8wpZq8EumL8w0Ssw87fCHkz
lHVB6jiYT6b69MZptClkGbmxUxzkgMqwpZ8wcnLqTNkJxhw1kSkSKVGokO6vDacvp51NRiAth5Cn
/FE+/mjicGWchsnoetGh2+uCaMGsO6ckf/3y1YgpJegKE/Na3Np9AYTNJTVPlqXWjqD9i6a+ul/2
PjXX86Mro+ErXtZhqpx7bIvGCSonMvvWAZTvL5fMTlHevMVoeXfWROGlI8jYRqTa61LMX7gHv3eo
Yg5EDK2HO7w6Z7FVJZRHszh+BgjGB4qAzPnuXSBZzEGd3GWTwvVsLaazUY3PyLKldFB7fWTEO17E
8UHdm+NvEUz5Qx5K+smknF00BVEvBs6SUMHbVnu7390qBuiG212M/hamZ8zcEuhd0IYcGTDXjcJO
9xwOt/7TKSiKrUwa/f44MsQU7HcPtOB0oOfFG6ew0H1e6aj0rRcD+pc/KbBf3Dk1ZZ+ouZBxNOe/
vlQoHyVty51ySRq/Hm+e+iwEu7wHIA4O744nd6JeSWFmPrRCebpnM7OfUvyedBdvrOnTr6GGvCIl
WBnV97p9MOk+oqo1NcuDEnFFI0w++InOw4perTXpIcl8fMwmu9fUbOo3tO4EDNZ+1lwTYTkZ0XCI
fjPvfpeHbpNtPBF3YfEYdO+ZAwrqx69OOPk3ez2+qN3SEHDPRzcfDz1cXFR8Mh2zlCfiDCzat5bm
RTlgmP6ocZ3FaU3pqi98EeNuBDyZa4K23QvnvunmIu+egE1dODAoLHJpqwnlTakIe05/kflpGES+
uuo/tBpJ+bgjV5v0Z0ujNh45IDcSgmh2WCkvVEH+lTADPMwOrwmAujoMD1W8s1zyo/OhGoJx++AO
9oWBfCsbs6PEbw5fMufR0N3HKbmHiGuqc1PjbriL8T/VrV/0bywdkr5dvnzLy8ZJEJ2p8Mo37g55
Il5H9oXVp0r6udxjrVgSqsqtAl1WTW9ETviNmhKuA5pCoHn/MH9jrQkGoQjTQ3a5pyaSoe5nnIAZ
ciWmkYxfFaYrvE8YmCk93uQr4HHuwLncmhF1hGzswTzKCuc188Z3MqOdGLCzm+1YhFv9KN/+eH9v
ea9GubgA8ThmtQND2k1AdeYBAF3Wc3xGCIjBl0oJD1aYcx5SH5NEUJKijfpQizkojfIm3xnvnrKV
nc/DlUiD4xddVJX1evsztRXcG5G2pXs6n6CiX0rJoX6frNvzMr0JndcHa2ZciSPGOkRg1M1cYe2A
3TiblTAoJvn/MRHOYzTEnjMlopOGJUBUJxNRzZ3VmXNeRrxn8HrCQ0tVbNPjUZ7SFFWV/wnXshqi
9ShMcaf+apapHeIi4UV6Van9IJW2ha8UIPemy1OAWO33KH3I9uSgX2cxFMkU3CCwRfhMPC/8Cdi5
rJOB+RhwhPfZ5TiIzzib5WvTn4TF1H06cdSg9IqJ9hsqbH0x2hECfUasqvKEFulUAlFkzesviuO7
TkOPFjnIw2hZg8eKx4nUWvuc3b1MtTeGlk/ctl4LphbbVahoLFzNo2sr950qfMv2VkHwZRK3CJc8
QOmHWVmuhd4EAsPbtQDl96bRV7qCBv+uEW+vFSuAbI5n8CnWUgjd7N66X9j3hhxVhsEVb35cB/sB
FwEtetjgeZMPXOi9oL7x4IJ+VMdvjSP3yZIwgvayudmMeCG2QPSKho2L5kuT2wKtU7KrVfrWin29
3PQXuha/sWuGXRSxzizXXYHk2IIB4++0/Bdc+0njdb81O4Nn3NBQ2agVu73oTFoKcbEafAlH1tLI
n6PbfiE7rRPLHBprU9t7r7/eqrmFaHdS43pia8ls1pFxSznXUvjbJBNxSNtkCsbsvkRg5uJPeFg4
2xHxt1FcZPGAzDk8Ul5ZOUVsiV19J10yc2fLo6FiqyPOTX9g4msu7R13qxcX5zE2KDLP5FXG8wM9
DqOsAoiqhAOjIdl/j61HxwLd9mLKwrUbdOiDaB/UzqUcyDkVzBKxqf1p4yBHemiy83+Ls3q3g6md
E+AkPSRtfs/Hn9B/I9wmS+Zcqi3UxWYwWCmGknNKXxb2SQrgjQZ1VIwAQQv0ArX7Q+KLgCtBaCWc
T4XvEiyg/dOw+/xoA4bZcQeD9yNPRhXxZe3+WJRxrWs7gumhK2E7FFd47R7dKduBKXUOigMb+cIL
73b0DbfOVdsCHycKBhStWdhz42ejX5Devcml4mANESvipqDf9PPn4VLP3c5wDZcbnwEOxeu99a9F
0rPGErE9sKKkZ2kTggok5COSCrmA/OTJyatEsjJpfh6N3NF1SBC6jWBncgpPPwtIc9Kx2KvOJBWt
8/pJT/HqLK60rhp3Qn4TYkvw1MBRK2dX2gKtcYHZqM6fKJEkfCTqVNFyCjCAihJm+z80OAfw7TGh
P+GwCbKSgDtMl4Op8p2RNR3cOsv3AogQVds7xYaLvn4Lxe+SUpk5dEbJTbElARtiR7jt+ZrKxZT0
SeIHzhj238lKgmcn7sINLIz3wFAaGEiciFNDHY+TExsMlYwVj4CdSA6wvjHaAD1ZdU6B0o9nIPkw
66vcjSBVRMsGUPOyw+EK41shtB649BvsEd5xBoeLC2oAIfSuoiOPgZy0GlJB9H3EsPgSnRWEbhPx
tbhbcoVnaE7XRUUTLjW7p1cmftFqspm8hGludbZz8kYtedpYE7ebsIM9Vd0wEb4er/X1ZUCiYdS2
64X51VwDxDftFLdD02W4jfgaU+hLVfpscB5I2cWli7Misrhnavj++VJeaSGuivtYaX7dk7FaR//5
Q6rJ9hFohlsgxLR/kMKHPrr/9cnnxG4ZhYyDMpcJ9FFHvsvmff75gh5B2fujc0v6xiTKZZmYwFCs
xjns5ARKUwH1wQtuELL66elQ8JFoEXAvFFZXYvP2KH/HvbVT8cF/400j8oVytY592kf1m0121D4n
GySgOuS3v1aTJosuZFwN9zmHLFJjm2IYf3/cAUXpaF1V0TRwkpi3kGfBMYFsODEAVF/+kTrftWQc
LTxxfciKF4HxdUk9S8WHS5jNpEE6GvuLRzUVloc0GuBaJVc0WP4lCDbtb/vx9itAkbHnLXC3oXe3
2HFglgxDOz5dDyHCRlk53e0KlqidwzQw1sFHV6kwkYEzWUgg6G9Ns8B31tD9pz3YED7zQPOanph4
EuAzzqVyHxhIMj4PpZxyBhOxaIZH2rvuokPyW+31Tp2DxT6J6tqdpBxS8a4c4poWI4EfmdpaKqEl
PwyPm3HB1U1QDSmeTqWrQMcE0RtUpIa9M8B2ZtbGW/l0ytgfqto/rQePFUvnj1VOdz3akzsrb2bC
lBC1G3oFdCRB0CYd6HDx0jfn+XxDpJ8XzFJKh6h22x4b6Mzv8FEl5jjcTuBbKAFQQWyGPi3MWJoe
X2yIr+eghKgoq8GvHPJN1y7iSzy5mSk7BshLqzLHzN1iMBCiKg2FOZyDiWnMkHaXvCTXNPZUtol1
YKEdfqPgUXvPiQF9mMiOqP5SBAZ33C4r9UXr82tz3Wx2OQoKqA6A4+kRSY82N5WkkkJT1nZAexgk
35G67XW2zQXWOs7sPRa62iWjyhqlgCoo0Vit4GAPkuTldZM9pCngopMrQQBunCD9DdAYmVFzRpDi
znqjjYLTVe3zSDmATYfHd3IGoXFHWBWO+YwRidQlBWyvjt9y9Ik0dJ0ryE7r99cegSmpVg+WEIOz
8AlteLfoToX8lhvaaTLAuZKN0WEaYLaocSKjzLv2/YzD1URFQEbzO49lPtJ0q1SAO0QgxZ463Ma1
xv7rwFJqR1r7bcbcokTUa/RaqaYNEt8Blb9UAE56FwDGDPwLq65bwVuAetfrYs0XvMe7L+23um/U
qSFm7Q5/Ll2AEDEJ1n7uRDIckOhmyXLQPkwk2O9UE8ii7SWWuvtsdhxfUIQJb4K/AH7WfXLyRckk
7eJFjqmpMnFJEMTOdSy945RocxguqxFT+T+8MBhv80NK62qnBT+rhoH+l0jcB3PjU49HcDbDok6g
/LloU9Gy9mO98RedAEEG2btziuFWOX0sT5vJT/rS4o4KuvrYXkwxoEpI9vZy8acpqGqhUORGcrR+
7IecwFDunpEJ4Frsw9Z4N5W7Sx7WFfz+T10l+IOmN07KUAwPKNmjPaFp/6fLsbb82p9fj+JAb5nO
LBMwtrWUMyraYtjsiuL3wf+JBBqePc0oDm0n+rA7pw8ivaU2B6Lm27uHO81SX6qNjHpxScTCnVI/
av6pWuo50Wy/9Srh/LEq4SnoHH4mdM0y5WSTz2/fz99cdVULCEoEEpbKs+nCg6KJj54mTbY0eMld
aloMCYNoCPnTXFxiPzBxo5/9bsCLKMojKbYkVRO9qrr2lPLW6QQvihhq2nlQrcjgZ4mfjVBXf6CJ
HWd/2uNVywJAwcC4TO+MQ6sw+0xOPCbdjQ3IyKZnngXziiH1GRUqFXsVd9+KrPs5zKLrnynfanbB
wXz2zdonUdv1jNiC5mtlQSu2D/unXAlBBqDHLKqOxXHyJxqKZujzZyTwpepEy6TkRN+jHeSwakHY
BS9rDrOut6w8DF2czHZ4nSn7Cn74Rw4I/kf1ER2hwfwFEz0ZnRL87cVZExH298vJ9aL5zs3Lgq20
g1WtaFFxjc30clfvW4mXDfiKfyrj8hzX51XUi0ltraoZJQShBw68Jpzk2FqW0j1q4zbYLXBAXUkw
mTzB9bpRhHSBd1zro65Rxgo34JBih+g9AuFEuf/bLKhcsoa2xQquScdxmI0SWWA8o8FWVNYBeDTH
lCeOVcIG2nx6hop0TuwQGKEnr+GUiPOLLdMbh5WbQ2JmK0oqBejt2fOqg8WDtx/ys+Qz3D6ggd/P
/w7icirQhp1CVIWnmp8OZlG/RWOKl9kvsh8i3ho1uJYeFI3LYRrKCGlR48ykG+EHvwp+w/o6NDKC
lR+gZVkuNXtT0qEt4RrKN3SBWt4l0dKow2sRyWQBClj+7Gtu+07sMnnybtgLdSFT0KWaY33R9QWR
cJNq298pPBlfHZ0qkiddzwrAR/R8c8XI5BCySCjilguEo4X8ocsdqeO+VmYUa+LHVHj4VkBZBOHc
qX0llcHd+R9IarT2aTsFlwc7PZIKSsSwnPap1oBl49zgUmVpLk/I0X42JUkFZBzOMlyv9VlvM+YZ
XUkH4oeX5TEkkExeRLStIopMoPYPrQrl1nv4zFWun9nJeEQICGvCkc/YRlTemwZy0ZobppDHikB0
BXEi5qKjj0r0iA0+808DFhK859XNUTysmJTuHVD+jeEjBgcf4jKGmufYxHugguVWijGYH36pdhsO
ECpIhjX5ZgWMnvE3BxjgdpfZY7gzzYJP/us3tJnD5asxRAH0svOCMlzxI2fjX8IBclUCp4TbuE12
s2ZU3SdYLWaAvMkdmomiqqriRvyoHQvrfSbhiL4N2cNZAf8/aSlbMjAYssVT8B2xEwe/ay25Oz5o
0g06Bj+knlBiyJu81RH6UTGLgJi7CR+yEiJ4bfWdN0UNpUKOiOgXT6jyquX3d0hx5OwW0usBKt1W
PGSPvCVErvdh1xVmvW9U6kTiLw/1g84QCK58/c4TMzUpuGTKhEstA0JQbQ0nlHb6UMS62772ZLyH
rRJ9lZ1q0AANNjr5e+bQMGwhzTOoAHJnEPHTc9AQtMU597IX0fLq4Lle6/Kdff4vvoUX+vovu+Ls
36MEz1yt2Xz2ukBVaiusxVTePVtycLA++Nuw8i3ZBeuZcYckknjvSCWNS3oMFe8giFP1mCXKNDh4
iPNSaQIJl9owHzlNmtff7UmRgFBAGNchyE1OyX7LsLtWWwpq6VD/vKmkCZuDJQOEYalR1MFbe/EP
eIWmT1GTixu0siFrwHZusF+xvxul3/zZwgCKNCuutuS1GvDVSXK7JHxRA4pi2WyOgRSW+P2pyo+2
I9rOiT0RxTuJlMYIyKRTcyaSaMA5BMqlFUkWhTltJbmJsWwQMAGkAL4BapnfGU0kNTCB/ymOhYux
nU9UdlD3xIQkPuZNZq3ppnftNLuybKmoQNeGif0QVUxQ4B/eyLZG8HNkJ4Me6dciJOXIWEXw1fEa
ZTTlf1srVZnT/KDB2ZsjeHb0tCHfxtRob0vvyWG5htor/Fcj7gwOckN6MDFqTYu17wb4bGlHdHk+
Wm0vcSfLVHBwqT/pieHlK1Krt9VpnJ7Rg7JToMgj9t+xrUP2qOsKFzB1Op1YLdnXD5Q/VJf3IP1f
OvwnMUlliwqC22tgdGBSQw09W5bhRlTVI6JkXn0lSPmwGuggFBYLbpXhfSP1oygaCUK6Hd5Fh0Dd
BJCzBujwonQjRuldJKb+kcOOt9iTZMUB6xSrtlWlxIOa1aLqZJPFTgiDyca4Soo2T1oqa919xWJl
XlwySzOtwuQZ6Bsflon+Tadc2DRa6t6JbtXJrS5igthgPl+bqtIZsUNmmUD31ThAK38f+Spt2P0F
xItdKAWJbC+bvjpEdThmWzCgFLrsgzKGAd2j7jhoTvJMbFdpVxH1a72Ch/qiGvRMfu1MMz5Oz308
ZilzuY2xKrm71ZqnSY0ImnMB9aslFnPRYDiw8OzMKzi7pqGqSXfKq5dGyyD0kpBDxq2ouqynlHO+
2DC1B25OpWJwYksizej9oxacvYoi54kyERvT+yR51SnwLjEdu022L+ZLP1ShqR6BmO41uAbVA+1m
5gNlSxhHCWWqKNKPrO1EI16jQMZH91oh0YZIPYTopp0JSAgu6XYDbpvRl3YQ9Yd7SfF42VAbfQ5K
Wk2OVsqu2yp1shm7E9DcSJvGUouOIS06U5i4FQYLdkPgKRilSWUhipHQYk2NkOVht6MOTSVJBWLM
2UbEFKbrrS/H79btfnuqoVxYUPMjtwDUaDduOYvBRfBHiw3cPiFn+sNyxp0xYmPMkFW6g+EoJnXy
WEPlYu+6JrauN/vCTe2Z9DIP+8nhSvnXxXIm+JQhD8ot5XOicpAauFCqUla9LsIZPJZ/e4ZwroGe
OjbGv4X0tZ+FElhy3AtFgB4tT26IBk6dTPSLsB5iaL6nbYonDEvMRWvVg1lHwEZdXwd5O/epaA1y
yn7C5UCtAe8nZEY0zruiowrzPa2HgmJ6HzUxmQBTQxIntnnFxVM0wJeMu4i9iDpAYuO/qeaQqk0I
5omFORIfgdJ425K26OcqzJqjU67to6IPEmPNpfzvxR3dciVqT3c6rx36vnEkNLkKp+d4gFPxaG3p
EdnLbnjKogn1ATkfTgOrGSIyQKM77LxU1dHeIg9lGlwZzbPHI+AFyKL4BOAuZDvDaViP2swVrVg5
BKaEb6JRsRjgtvyxzm1YVWpewhniFGDfaNn+7QEO+fDboAsbYtgNk0tb6MecnreF67J9pLQDq6u5
5cefpCbvzCqLX6MGApBWG10zj2pghPd/Q/zVAcXO9ux30AtHNDwNXzMM0LVxJUa1+nUNxTxyfnf5
E441o9N+9/L9aDDirvthH4se/usKp8nwaL2AsUrqrvYoFvzZZXRy+pB4TZ3Odzvr/NtCYBzVSj2L
F/y9wzaDRRkNXoIbOj2Xz8w19iyxFgpKYeD8OtdpbOU2nE1USsdQnKL673cYYe3CENQbUmXVZF5D
KpswdttKhIu+ciute3HQsLfLO57inrK34KlnzsOBKdTGD+wR7hXua8+2k9xV133/0AlcwD6uM5sm
HCYhIrXtYpM3zwAvQIu7vJqZ0INh0Aq4/50k///OxB0tAxGGwW32ZHH97iAvqh6yiozcxj6t+k3l
camu0G0BIYTCwb8J/7PQ6bJgO7cdg2+5esNgSidQuRQ5ota1tSfBACsKIvOoMy5XcJsSyP71XxS+
DaGADWUjZTG24bHhacfob3fer+mJNlVqypGI+Z9Mu0VvrN9ZFQvDMede6WkDXWsayNglJuFJXJwq
tBBprxVhJ/wmRNkM/k1quxcNYlY/f6qx/oqpk2zucO6mWXfUQ1o4PmQ3Ud+YNa94qVapxK81kwHq
ztIs34cbx+LaqRCcSifjCMykVAB6qo6afYLHlBeah3rQQwsqZsERWd+uJ9Uh0kiwyra+OX9phnNe
N+ou/vxCkp2J8eS2PXnSlXdrCMyk6zbf0ZULq7CadbFd1wrRVBjcNg/VMcygNcIkq40z1NuzLEQY
UT6UGKUC2SfGjyuOrbANE7E1QWiQGmQGk/ZkrN1t9XAjyDpxj0ejEHH9LnF13LBO9XbxkLq5nmhO
5ZOpGH55z/QWoeGX8FOok1dmtJ42xd7pdW63A2bDLavly29DOWN44pv05oIf9Y2VoKk4sTvbnqtz
YBVxJB5mFcqEiiueElwkYBxU1C6bsZEEXX4XB6w00BpLzD+jn+F9SzALDKxtursYP9vZo/qQmBhu
1zIYR+jQrmcmVVbPA6/Adlqilo3szk+Bh/OoF/K96CqQ9xwaV95U18YjGB8VEZtjOTQg/OyoP84P
CCwKeVlG3g8a0Le/pP27ZcHEqUk+ovQpIMMyy2ouQIDB8SiAsqsxOBX/e89nC1kIFf7PJNUS5SQE
0q7RQ21OmfoqAeOOgnd7KnqiFeMpQWxNF5n6C3RKnnIae4IIPcxcwlG/31DBJz1vfSx2gGbV/ndt
cf8nTnhOVkWlmYy0SWRxdh1mOj5IOyIiffw7jbf6cyupv6YIeRiiG6ODsZOZTC+vbMluFVSlVhRw
02Oaa1etmJEmIqVeKIKvUqFm2Il2wFyuWS+S0VvS0SOf7B/1250zOmQDIMo13w826ymAv6+NVbV5
Q3tDfsn+4E9yaiKQW5qYWd08Z/QBNJqleElrHe4YJ7w9lbC6HIsxdFJRwg4HHy9305V+Tm6W3BRv
RpPW+AafcQSlCrbDBK+0sOwcT5PvwY4q4XF457ixKLVUQF6X1xYfyH3+1VkIZY9WbXEihT6TwKpT
V0Z7JDxvYEOUEXl6krrPngGPtwUd9g+gLBReSLPzI+oih9fWBDIUKK8Ubha74sAe1G8h78/mP9ph
eNcFtLxh7a+uRPEm5ce4ax4uKzdBMF4+6aNrO5K174ndqfFKlnWWaewRiyXaReXqyrUGbTXLNcBd
vJfAncKQwkUrXEHQZuJUl27KRfe0KyfrYwImdEKLxDu2zk6smFTMdjXDiF2LdJPhWkJK66IrfZvY
whCqZaKkEl1sCsvf3aItF0S8Nke6gxRRIFC8dJzdbOMWk3Sxv1Cdzwi7ijtDV7k/msq7t49Dcmqg
svTLB1cyZspEfUcS0EwNBJDiEyI2choyJqVss51Zd7BZQmPtiM2Cr4jujV3VjgPtESksmvUBz0fC
OUgdDAPSnEkArKHZhVfV6356Jh20KYXLTVJ/Ig4xtLXOeoesLUPmq6I5OsNsHvP9N81wnl5GHaPt
jo8Ftz3O2swPmUsBPqd/bmWSnJGP98ht9a5sAjtvhWwVk4Ojo3M3c4IZvQHvQZ7kJ0GeKWUFx19x
cMhBmmgj2JpWxfgzjy339xhl1+0SXDJdg3PWIbLTBTjAsfbytcE6xll9o5pnlPXCyvXC8BWbg7kM
Ae8PmUW7vYdldcXDuycGCTXz78kb+9BtlxtJhK8UlboOw2Cq+w3B4jKOIhdZKqhdVTHYZS73sH/p
5QczgMtDBBf1x2iMZ4OGhGMmWmWkkFeN9QbspDPPCZ6qoOy7uvpUuh97eeY9zJx9co5A+0YfrxMa
3bvsy5OC2YW/Xvf0hE2h+xV2dDukz3CnBKr+aoN6dvriGHKQaeEWYXoBpaMTRty0dWBzFItXi6TR
R8u9rAM06nEQJXtXJLMLPj73+E4VOkw9yY8o4GKIjGJtSfB2pjQEq/3Gde6qACxRfagdBJpyMDsW
EG33HyAQElZ7m2V35uaQFAJyUOCGOigl42N6Owp17V7Z6RwKzbBXQmWUND7+cV/1sgwJjWS8y0mJ
DzxYl+6r+A2IkStv7LiWLPx4Yy87kWfAwJnZjRJ3NzofFofaFao1RXR2K+HBSrjdZFMy+U387ZHd
fozNPL3Is41WnMSM5t8tavt2iFeB9P3s449NSXnP84gD4SJ/B1hjtxPHX4MjOJ2NP99/OfC6YOys
QVp4z/8gHhOBtDzuS/hPewcpz/6z8Ka4nTcYGXVQr5uTKpn93WhMOy5nXf+2VrHqQH4id5047Owj
uxq9BSECook2YFcP4qWFYjgW+faCPevKOwhNqQMBaEnLpsNCXkySsVDTa91NRagCDUQNsHSRkMPH
qs9065oDdsvixTjV9FzoHW1OhVAi8VRmQt1kX8XufZCwxL4p1vs4LWYkuRZRlyj6TM4trPGr3E61
+yEi3zMISZmeYF+bnck8qMfF9evHvsXCn2CiYbjdGF3y9gANjCqEFiTw2Pc6RbbO3AOxUvHZaYSi
eGnRAmtDMUmEcmG/M4j/QR2N5kLYAYySwzt7Q66CzbUL7NDZRxtsws98A3uPpCSE8ItV3NabCWf4
GQ1p+jOGd7QwRZpB0G7xZuJiCKarZ4QFImdinjdjsDNft8x2SBl+o6J/KooArMEvat6GoeW8PTLL
RDJh9k8vIOvHSCjjit7JHSbanGKqFYrAWHn/87VcbMiiGNgohVy16cpS4x3X091RwMs0f+NQ+Rft
ZcnasYG0QNrfOiRs6/weM7B+9NQaEjTZ0cgjZBY6JllwuU5HX08Ol0KIcSdFdFzTDgwXtvVnsqzt
YneVWSGikl/9STRA0JD5+GJ2RhruKzb3xdLc9+E++x9YEdtqOrdzro2Jfd4H6OAMcFnmxu5VjDVY
q6r5JfO1FIcRbpAhGypMv/kwlND/0hNEuxRV5s3guktX34j2BNWrWHs3CES3DbqBedHuQH6qYsf1
HVTicIA1wwUo8gxnqOFtB3XZ9IuZgPjp0VAJZjqKCJCq7fo8iT5MekA3We2tBjgDfQhERYZMcJtJ
MEnmxd6OiTjzwf6ZT1t54oaO2oHknhqF1T32nSYqNcMPW3LQSW9+5q9BdjADMPtgpYAOhIqrxKuA
e7Oqx1tOXmVog8B/1gpT7Q/mf2tZ2miectR2CqeV/lvzusVecZW6gZs8lh1H3QowCGio3mLy9uAo
hwf7gBbTdPaMbR7bbFVC2ybnQlFxs0P/oLKbH/dFVymS/B0zccaS9Bnq9NDA3xSeTjr09+/A/7kh
5WQDEx/hTBC8qnxfRiEX2S1LC5xSh+UziyrwqmQPezJ0ZoDT4GOe5uT5Z8lu+SzUADEe6cptZYRf
/iBdUUInjkb8/yTx50XE2HOhsBhYJHabQTu31M0/yt/eOctqfg59+T21/bYq6RLJfADcdxFryBHq
cXpUEGmMSG+wrFTcohzqSBVb3hG+x4LQpB3Szqe64K4loOHlUM+Kzt/twHzk6ROdzj9nQb+NcRMi
zyt2RfAg7a5oEJp1ClfB3QyH80jVVad7XRv7ZaRdedbJv5UHQpYvf8IcANLKRTYFQIeL4/w91HpE
NChNRXsDsCYzE7LprQnzMzf4VayKcATaSiRi2FwjZkvHK+V2ZqxAux25iP7TGRPQJ6emj8L1lJ+x
B0Fnfmt9UFf4IEQHAKNJqU0QXBXNWaGZc8E8ikXww6bMHtO04/6Ze78+GVmE5BTjdBQP30qpR+7M
mEyrRdwMlOfKAfse2I7a/UsFfQeLfua7g2BQB1LgxAmFyKeIunme/c21/Q6/Z+LbdSK/Kv7BrzMw
liLb6j/6T0xP5lUmbJ30Ykd7besYmQjIeBj1aVXi8CjvyasVPG8kb7nnFMJwij+mRsEHar3FozRv
i14fKrjhtLonljpAkJh8kdPbnMcUOWknXAiH+rwHGVq6g0gKi9fEyENdF/ZWLDnbJpqA8K4L6tZ2
zdy+ldNALdTfgR4CfhrQYzK1R7tBOXUECrOaGfMgMF0DfiWRtCE1ENWJiiarwXdSUxt81y77vfmP
Xg7xmGQq5mrtGutk22w3jFIPS6rka+X4hmSQOh1dLs4SEjGELgE79pSQf4FCOGp7IiewhcXznUy0
mikaEUYyTZgDQgvISbqXrwhmO+n+ecYJmF0g8I+F7lWEkGSffsYnc7Zlvo301DtaE/L4HY0EhxP8
qStt3sT4uI+95hOtppNIHmL9Fy7MHY2NAf0tddAX3wSVjaDwl2dgardkAC9fUwVIgcAJGnA6507v
ojLqEFaaTZjm+jI1xGaWMZK4IFEhFPaVioqalAh6AJwfIMBY6s2Bvhc8tKYiIwlsmAmQNCePQN5U
hwhTniAZbwqIVJBQsKj5LgyAUTr0BeQGOfwmU/f1AL1cUjojyi9IFsMSwUUAjQPV9pEwYwYgbo7O
IIhtVCRZPIUa9al9XSIAvvjDYzdLTkHjf2a/uNiy4CoWcv2p8P6c0csaMkoDTNc8bTfV5oVeabFj
5zx/o+UtlyHPYEQ/wI+Ip+W/58qCXgbJPvuymxrQpm66tm0muISCu7GrkInrmAKRWrfdhowymhta
swubfQI1p+d9nCNeVrOrR0OvstJQjSqqAWYQyF9XDDfynzMuBg3ExMsgFH3O7HH8Mk8XzSToXGT0
h/6muu0RoslVmCgOkSsfmmLPTCFoH46HNflVwTro8wiGvi5VuySH5G3q3ULiZ9y+K0/wIDyn7qxi
668FLL0zlRIEY2Y1ekfoG38Y7iTZxf0wpBI6sJaZKswJKWA7XcqI0UPXPeuZIoVespMZv7JmQcsV
Bg/gNyts5liiWW7HjiqiycUje/zNcT7e8ktBXHBTGJ0BCvjxe+nYzFauovF4nwhAww5XcvUo4Y8M
35eUw650s6fjiQ2C2Z0fBV4WY+eipFsPFlEW8ewPN0eYOgzoXTMukr3o4yUc0SN5cdGElivtJMZB
QUZ8nBqoJ1Wvizksi0eByBmY6kyJzstOamB6Ncbmd/4bkjo63WcsAIs6wHQXHH5mmnjt6Hi9dzIB
xXiKkw0gObv3jZaLUZUy74dOVv/U2P5NYdj82NNRgleer0JLyY8P7AxIHtaYmyIU1Rw2ut/sFG2H
/wja+VlZq8DHtpis6uWxIQAmcVvIWDpVPhkhOb1cojwIj7cb6TkwAoLkFtQJolRQsMWZwX8C0Q9H
naySIp2yPj1x8kQSnwexO5T0ffo778sGWmApvg6Sh/DMLe25V2iGNyc+FHrVWXUL1a5Lc9LYQcn7
tCAW2ZzQchDQqesqFhe2/KyOGGW1yRIU/S1mGtgZGHQ27VESIKiJpK9rWMiIGR+N2F4+DLAc0+8t
1fBpA9wDaPPmZyMNyslkC2ltx842nrKrmURSE6qb5Uz+La6QshGeUvjjIDjopy3h+U2sx6yj+idE
XmmuD2rBOaDJYa1PVmgkixPbalEnPoF9H78DMU6m1UrHhLc/PMGgdCYnmUJWeFj+hGbh9IGt0xsE
ixR2ISbTnTfUDEdydiI3DUSe5TE7toNChaWhqXf12cvxdK1+jYplAMzLYP7UNBn8PdW9ugE+nh3X
44X7fvgKOnC/mQFrI7786k8vtZ+kcZ7KZH1OogujV6fqDuUBrUafRmVpsBXTIgHOkjaB7FgypUhm
knI+FfokEXBD68We7fwWCq80NWFMHv9XBzrfEDzxOXZ3KogIKLeFOx40auHs2ELoE+S6KB+h/kT5
+9UEjS1NgZ64tTbKEx+6QiIXoSOJ/5b1LpfqwHSyfGZv4wS1Uef4ScfS7xpcYAbot3hxF3+GTpUn
xWqfivxQzwHFgyvxLdp6FhtSW2mehtGCWsUnkxKKyuhoCPco1figDhiOVS7LZhOGwdB9L8RwRcpi
16HjKITbiPA3Q2zqtDSj4kDGbfS4SMTUYMwVPi1azqfH6CvuyZHiFvrfgOu6WcbIo4axgoND01c1
adE6HoRCS65Z/eDtIXxJRgfzal08Q5FqBcIsfA9xQ3d8JoXjfEA06SII9hcXPOGVp1ne2bMrQAaG
Yi8LP5vWpLqjYAzy/Mxf3AGNYpeWwresrtTbzx4GqMv8KR7Hn4Y3Dxx7A407wRp9en4GbqwcC/i7
ButXsLgmwgYjjb50OZVIEeZcKb7GGISCZF4EobGbbOqdU+7NU7DiGcRG39W+o8BVzz4MXD1tdzna
wlk6TepXIflujkm87FEkPoeqvUm15Y4wKu1Ro0pGiFqwESzmraa8TUwkIDJWrzutwmlv8f1MtBnj
EpJJNI4DDyS4TPQ9o8AbQIfHD+kFChJu0UmOJukFgr5n8X1daiOCZOU8zw4NfGDNEzmpr2EDDPRH
u68bzJ2jWL5kYdAS4S2hUSXS1ANlebGNtiRt6HOhVsq8CeaYXZ1E6gwdOKypTEz0Ok2a6clu6+eL
Kq3C6Aw0lH0ctGeQjBZIp063IssDfHO7X9erUOMN1iB2AoCwO/GEAzFHP1bDNJgyKJk+cxArcQlL
eB7CeeGJ92DdLf88552ivUn7FCjiAxmKY5C/7f4iu4bK1F3Pi8dGPn19CrfBFeJipz3ymMbDC/IF
8whsF7hPFw5JuKlO6YOxJkJD+OkYyI+V3oh2uxUOfuG83WV91aRGADX+f4tKE9T6Jupj6M1iuF/5
/ZgDwX8JGJ/M+SgW4A3xxT7kvDQpWvCHq8+tUv56OFiQVTTkY8cU+CdFzOmYZZ0szOAx7MCuWrP3
ojtG1uD71zCo3onHQE5xndZBmsmXz0zIRF9bz70ekxSIknoezom3BVKYexJHiCSEgBrOblAAl1m6
4PVaaPtiEJv4f9aaFEAExDCCHyNfVA2BF380lZqPS1+zkE4ChxLnM5SpuQsj8hisnHPisXjJ4HTv
0Vr2ZtUf5ywTrt/tALCNH8RdVYUpndA4mFaP6qEBFFFJly0Fcd3CsImCS2c9PkstEl5PbstNGv5I
V7hcNHpaWZaxRzizNL+AC+IGZLAUA+gQ2c9I1rFFOB1dFuyo8rPvYY6b5HZKrIA0sYMZDAG6Zl+6
qhrnErVLxu+q8QNGqtKqCTmF258mQxRegwGWsyOppON/drJ8GIFa47VRajVj94U5eNT5+HQPzdvV
sRQi0sudcHW72ObI8Gp98CniglenH0a8JLhiC5+gyoeLYArjcxMNAnsyci1KLFoQ7zlhGqrfZGoi
Zsm9BmuFqoYNn4kah93qZlNunwPKzuRhPp6juHHgeiW43PeXsB15AVR0wh1TRP8tniCkXFttybzJ
7/IxVpfleXvE9JRlqQYMN3TG7dKtuQl32nDGUCQ7fex2+PMYqPw0vY3NsFhC5bnjcpS+FUng+awu
a1Qo8xT/rahtoh9juLPjoCr1h6N/I16MCQN/bwHOXk6JLiA9mwjZ3OciZi6wKtLk+Fbb5r5XERtd
Xw5qzKLzbRgktLFn/iBYmUCynV+Z3TUdCtTh3Iw24yRmWA4KRoZ69d/xAR/Jd6LzUKbVIBFaEMMx
hb1teF4kf9Cmcu8VmJbsKZZ4P7FXSP59fykJ/LwSMzCgWwuf9Xey++XM7Hwn8BCseMTD5uJs2Qtn
RATiO4YbyOy+i4HLhthv612U4p9ievJFF2qsvWTI/H36F3WD3n22g9yAkNo1JFaboaKgB1utwJ/u
OW/+o3COEgtVPWto9Ly9zTnSIdCs4xcHLtFrMZ3FzE8E43ggicZRbf3OLz7x6OvFvBxpNrGTmkmm
G+oTLPNm6yGXZcHco7YY+FxmgTaaK3ru+rl6DlfI+l6UHIvTGU0fnJ38JcvaIfnjsU/vcwOTZUkR
jy+ZGuej30Yt1C8CRQtgfb3RLLw2E+7tYu5bwM9t4AYtnjdgYaWp4z2sIfLjtCcGUiCcMeUrktoe
s/qylfCf03++sh2AxGK9NtAA1nxh4duiT2NygYKocKZ7Qbv7AL1HHt7FlvAnFyFZQXrhu01xG/yW
vaa3N1mLkV+Cy4Ga0eKYBNVzO6XpqrCvD4w285cK6snOQ/VhemULIiDWocyqrvV+vD0Yf383t6OH
UJ+eI6DmknpGzLBek9Bf8NdRmkh7yiRaP+ZwCd2mPvv6sNRtF6+cRFE3HfFEA5hIQrSKxolTgaj2
LZjqpRNWmlZIe/GUjTuyUaNsSvoQuyaoGYVK4DCJWdZQbD7+pNP9phAsa7x1kUJh+miVSL1WlSh3
u9IactMuiJZxH81D0jRwlD510rmNnMYKD/obBmFOrHQDSef99jVbdtLyvEJnogTQqTL5IKWXfA4M
XPo5wNbPaiWHu4MV0Z5C59kZYA5k6694ZXrFi5qsCWEiLDVcJjSajUD4qYxktyTGz6n5Oe1tfBFC
fJx6BDvMGsfwnRqhn83xRwJHnQd5n02tekLNFPnVygKYVb2C366y/JOPqatrnuteeZpzSBAUrJZj
+rpx5Wcor+kkuFAnUYvjCpRpgCu6EBVjufOij7A3BP8d1BlgMlx6W6aTAbg31+S0O+WLfiiWTGQ8
hlewxSgelZQm3MAtAsndF0jL5rGE6xCxKLbc0hTt5Jl+Q2aD9VlqMEyHAbJfx457QB47t7PqFWwx
qFUgz9ucYOYAn1qcdylej2wCVmgFRVwxNexjnUqnjkqz/822ME/5rFCgVqVEyZIY2gTH2eJNvCUg
eQpgh65aJYem+pfl9UGigoI+hjDHa5hAJxGExHtgpejwR9eXEyQPDtAnFknMnYQhTbQNXS1Di6Ci
iHK/EeSaeJFPRbijUrdOO8i2L/YDdUxLScRlFZrVjyRNbmm257RlyV29sf8GTayHJSBVYCGyR/ba
p7mVPC3MLbMazCn7nKAvIBen6jUH4e2GdkUk5pWAI/mQqro8KMsdatRcAkhJvr+n8HylLVYMaU/j
yMVAXgo4YwAR1OiQy9xVZb6CNForTOcaBnIh4oetkWMBTgV6Yu5PNhNWiXe+ZWkCWkas/3Umj/GL
pHTEKeWJusKgznfhm8E9e8Zf6/5npP0A2H6HJLgb8buKSO2BZqCR8p8KWtuu2NWZHjIMrI+YJS1F
dTcp7TJ5iRtCBI5l+8YigNBMVc4M4d/CHF7Ep101PnAN34cVsbD045MmWWY/uEC9JJGb0khUGpMz
VHtIB3GvUJplXuNR5QCb6rgqd6XjP4VbpPaznNGhSXWthSVRucjDgZ+0ayMZM0vnixRm7qGzS2su
vvKJ8A/owJHYEYBLAPjaOHQCGBhWdw0EV1MdwxOef6b6uslBpxHWhsaGnapvD4G4FDOq7BgskwGi
CRaBkSQuDeo7pGPq2I6q1smCn0RM7Vezshvk8ifeE3UWC4bxRPoa1RmtHh+orl7GjuAx/Phmvhlo
N+pY+fybWTdlKqlWy70VWWO8StOFgLgICd9bO1o4UQOchqsxFTKkcCDlL+QVpU2bc57FORFd7gi8
1zxI5dmQhkZCInuQ6WJtZwmIp0PFvq/3adKHZp+e1ApdYuOcMRB0EJ4wQoFQ
`protect end_protected

