

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
FZWxslbw+U6Wgup1K8ZmbZ8ZvAwEdSXoQX5Zxu+YDpvGpSAvyJJdij56SPMVKmhf+X7kxMgvbsEm
5B5AiAyVHQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ntA4Op0vLLt6gLQbdMxO+e0Bhjub4O0zQAgtU7SVthNE2o/5St+SvTkDoJ1ve5MFs/Rgt4JL1gtd
IBaLjbwdyEGV2JKFzmLfNOLgk4U4bgeRTGAx1e+I5wKQlcq6qarG8xv4yuzAX6jRFWecgDUKdkZr
uIZCcXBmuErGbIdhFKI=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
I/9QBkeb84dQg6xWUGWLN64S2R+IIBcNXAJuDMwqYLTsejjUFtntzi/OgGH9xu74CzmvMnJuiSkZ
p7NF+AufXfE0LUxVeYNmvB8UnCKeswDMIWMuVEpX3XPk8OVFRqBWCRJ5c38XRjldLuPPEii8dq/d
MjasuPQowI9n5pgL7s7SczhrYfNu0A0XEQTAwaUPGij8aO4+LpdeoyqZwdg7p9EXJlysFsw3bvdq
qHiouBqf7MqPbKppmCVMlrH1R0q5YlTlllFEZblTUq4IO2ZWi+5zgGnEERNaNBZQ/na3tnrwOTGu
mqAR/EaIPbn2R/AR26ZYNuBuu0Ym5XtWJuqzJg==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
jRGmdT13qAzfiT1K2NPIFkj82nI6QO0hHDoQ7U+cF5NSt11k+3KuVBnDKOWta7RjBJSeiJs3q5WV
MSQx2R9/yJGRUjq6DQS8PVF7sqUyuFjNc8w4wdPwxcG0hsCFj/tEGyFHTU90BhMVIeVjf2WlERXd
+UzGn82C1ATZxC/M3Bo=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
c66DzsXEGPMNOrzYyBeymw4AV+RpL9x7eTO9Hf3l3y/JxC1wwEbipw1XtleybcrcOfKY/ACDBUVi
s9qFxHBAPyb46Eh9l7EGLGzxXJTWMed4eJI910mZ+WMPkBgIF1jvUqr1JGStUHDdUjBjqP5Bbe3m
2g3HBNLeS+8Ciq924vg/jBwWCA+G1zUvjlqI48sc1XMFszL+AzQf3r5t6tBvdkd9goSPiuISrM7C
eaSWriX/kCtr9jogh2EYVx1Ud4JT59uRVRlS338jlkF39xoR0AXtgdhjpZa3Qu6PtAnEwyq9aWWk
FBo+MHknw9HNH3v+t/wWSpyyW9f8/AhQrF1o5g==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 12512)
`protect data_block
3ZGowwgE2kmSnPJW7wBFzV4uGqfQz6qFKsuDdjq5cp47tQ3EZgyJKA5wMASL2NmFBqf91Urz5ZsC
enBaXVhXyCNH8V90EoUOlHKjqpe4JJ7/4N9PO8Pv6oNousI7uPkIv7ic0LhLpkLU1M7UO6AdHXp9
GIyzDaJhE0b8qtBaBG9pxk39QFuw11p2100sG9aNOlczkwJ+4neAXhabNIv9t9HrkVw4Gk1DDrCp
uWdyKHXxFiCX5wLKMr8MiPp/GVTofcETX+GxFP4WAfT9VerYl/k3u0xXar4O3AuadSn3hNFqZUib
N1ZdveeJzeHfHbSc8aDE4sAbQ/dH1vSqBy8m0pC3kPuf+63SdY2sRaJ78yCOc2us6o4z5VwmnvEc
YloPC3IXx2SoUfltzlqxhnLmleGUqrLAg4IGjzojoeHJ4W+CqGCdnuu6ACQp1PNRnxtCYYW8KH2/
c6xEtNxV0eGYofA4UYXFSkVpcFsETaEW4F7FWaMNGH2mIzqDxX2rMQDA44ssR4IpFsP9hU7V5U31
mRhs/80JUWaQW49Z2Z3/oKa/jtcj6nLlUwgI7s5/+jI7zuTXtzTTaq1zgozKe0AsxEzP3Y2k/HHk
rfl79NeSfWm2zTQG+EN79qMP2U8aFUbQkdZkujIH2Ey2tqbrttjZM3vDBxwmsfvTYpyJfGnOdXMe
3/FvYmJ47PybzOZtMC38pm+4UWS1dZhmVLy5zHEJBu3HdOv/kWZu0AOmMnsWHP5jUhabR8rq9ijO
yrFDbnOde5TggDbJwXR4b6Vgq78vWI1KlPycikw/CuG8lxRCLhboVcdr2SVWxk9Ub/bxTvjt3lqg
sMShDUdYPL/25bd0ixQaVpZ20CH0leG+H48xMjhiIcY30nozJdFNDFksBQAO1HQT0D+OmVXpzm4v
JBHIwBw1YSTYBe+G5cXM6RGW3rfWipI1c5TjK5gG+Aek4W8zYKih2iSO6PmkWQkranY2SZBjn48N
O2RGY/F6JAb0TpyRi2khiBt1+zzg8O4rzc1pYJUyHS1zhZRSUfApc6IUN68pi8Ustz8Pgv9VQv2S
btorL70nqPkco2+GmIjn5c6y35DxhasnA1pmoEzzsqgwPr+s+iGuJ6BK+hlkQ+vb3dYk3nkSnlzB
hskIgiyOsSgoErR2iSjXDEH0cpCTFJBQPSKoPAI3GBz9oXOx16AvuwjZPWCc9hxOUhQrdORsxQg7
62Q6h2eBWrBqUg4GQhdR3OwakI+daHDCf4l07OG5Tw3rgtwS9imAKRSgLM2cuVuJfYjvACCQDBMM
bGI4xeVu1cFkjT+3X6kxJXwDT9ZsaqKta+4w2KBsTUl0LfibBZcVkoMVGZZ8vSZX4xBeBBbFEueC
oAAOsUW1OKhF/8KT07Ovl1sA6Xbf8lXu2ZQQWC5hIGhVQan0YTClplDCvgklXQEKnKLR+1n9dOBG
62EqQjF7PkGE983SykVfzgDfuPUKnuqL/5gjjeLUiAuDr0x3FQD5RmDoVY1zFqTCwkBu3Gyd80wz
Jd7RuomZlYdxTX53efVksuv4+T9pIwqYC3Nml9FiNUehvMx/QGsTcS3ojyTy04W5Xh05bHO90AZt
bZAxFUK+7x0lZuNaB7a0wzaEV7KVnBdMw4xr1hnWpTsGpsthnvW/jRgKXpgfruVqLaWjJZMYiPe5
mvESX79+LZFsVUnDwTc3H5a1Eqz89UEGg82xUX7LunJpfSJ59DPSiD0CbQZGIQnjSIT9RdsY4znZ
h7bs/AqqgzLpdqjEH10lFw5prdatN4v4c3uMtjb0Ksrrd9B+A7oQaPIKwXiEOKM8gEwFFkK+1+V6
NV+6rP17hC9deQa34oFrMmnUuVy3Aido+1DFVNAGaup/PbqDr7NLjV2W0DOay8ban5vuFUOc6bfW
0bcNaKyKIYHdG01+eTqTFMTtgQkKU0CdvDOCqooeTpJATZ9G/so2oY8aLhMBDLlEcZjsL7Hq3kml
EaJ/rQoJktBAT1XVIIHEcUpnLwU96bZbv2lBbACZ55y72XvEDPHwvvCr6dPuRRl1cXCLIQAEx+ZF
fsaYnb/x0OEmohfjj3nutVUu1chv6nt+0F/yYnswrAWCjdEFMCLfZR90goUdtDWiZtxEwb3xFwVU
ekIoxSRNxUCBwpv9peK1ujilexHUQixL7OLVh8fnP6E4q5HE81vZVCaYtogRF82zX1x/xbh0R6k0
YN2yC3AZ9X+CBbkmd7qq1TdXFeiN9sc65gdB18A1HpTIQc/+eG/huy2/2LLmBc+wlGyPjwWuW0rd
FP1qmnCUesCqeQkzHrofOlsF07FAkQJO8xVeQBqP31MaNiw7JpQgUp+NNJ8n8491SyNJgLDlPdkv
dGrp6yyHGj3Ie/YnlMcszHRCu3ngkbiqdbdGm/6F3gd41uUqIQTDYc34QsiAAPvApcHWSkc3CIa8
mRFOHQABvDqZw1pnARDBnu1CPR2F+7umKkF8SKRLdvkg5RKTDILbKugjbfR2MLUc/Bo8mgcDv373
OdaJx7Qb6PcsaGnUi9qNKicRmch0zeCz8Ox49HSK5b4uL/qHe8CPlsKLpLKG/AnOBTJdR3Kj9gbi
AlYE/QbLoNoh0ijIm7l0VCmBraFivJXJ1+Exrqvj98P/gjpI8r9rO2Qz0spMXr9Sj34TYKDrXCfr
uw+Is4CkDg/vogpyKobzj77uXIQYqGdmRYSIe4gtFFCqqz3XjGaFNpU8Aa9tpDKo9VFeYGp2qESd
HpzxjXJM1JN5J9rMBwM8XDVJagIhtaK0IIzN+khfbD3zHRtyZynJOIv5sZZFlP2X/8Z/aV44vi8m
SPMY/coMHmNYJG10Z3pxkwqbw2qQH+BuEOrL0bUebW2D5S4UpFcC3NBKJwSxuFDxxRv33baX6a63
v55NTAj7hx+gpoReaX+vePAHsAT8inJu8LthQ5ek4zXmd+6m4NQCKhSVQjV8LlJCH/HgEvFX+s8a
dbJSbYitgI163jzbiunioW6pPbH4xdnFaRsfU/HxIUv9vVteh4hwiQzug70r4GPvFbG+jmxU/RhB
S1n6WbpZC6yHfVSfXhRecY/4Igwu1Fj5rclfLEB9KebFqXRR5UtQP6mczxLpG1Eb3OJHwDHIR7vV
BtRLJspP66QDiPNsTdEB2+VpZBmGmas9w9zzUXzVDn4ImRjETwAcYx8bvddPz/jCeogqjQ9oTRLm
FuomL0gK4y848yhXstNnTtZkk0oCgCN+HdMH+cAxesm+iXRd7Z7gB3aR+oO4E6XE7nteqO2/9zNq
yL1fPMFiPSfCO6m/CRjM2b6v4Hk1dBNDfO7mFmABnjbCPw15PG41ncTyshBNW1UJ2bZ5ALyiHfWp
sSRIIZ6n5i9FXLTiAFgmT1DuH5+oqO6MT6rYh63myTRbCqWKJja4rtgGjPSAPY8PDusdihGk7+Xa
zWyjAql6XzUkXuUM7SroAOAvRLsJnf6thlkHJvegflXr2wTicKmoSG+t3UhYk5gh8RVCsqUifv41
hZSK8DJOPpCK/2WRtfXXCqWxqPGvAJ0vn/7+zRO9qE92apNUXKkNRyDrbdx28shGprXvDa4XNqRJ
VWwxXfauEyR6a7UY9Np50dlOHOMmEVJyR+BUQbyMKkDW9PG5jCHtvA+NM+NuxvU7PdOIYDsUhvEr
l0IKyLaQzC1J5MG5EKNal0cHXS7PJXByFmjMi4Z1fcNxIsY4YGJGdI1I+0lkUBaFjGQIHdrBgTxn
iBdyI420pRN34ahvo7aGUDetOfkdsJL0L+dhszE248P9nKM3f/AYltf67o0JMpsKONoFPiH+EPXL
u14V2ukTp+0Qs5gPnZ7kh9GFz9QZsTmQg/l4nSrUCvIAZSX54nEEsVOal0jnd1ZZzfN/hi14wc7h
5V0xBTfrPIfydNndUd3AGuEY+ZLdP1FxMSMJ3Zw7oKTIe4JsNxytY86d/3WaICVcRFPGkaVXoyco
WqsKtfpalIakZMeLxX3CZuLHQ5uX9XYRTy/CdIq/3MN/ctKySczDzXFpT4Xb47h5wY3JXoX4JZfC
nrPOBinKCGtcdC76cCTITMSgcVI0DaHAkHsBlxz8p/CdwqvkJ8BYyOyLXBUhTYA9ZYVz08I46DEp
BAKDVd7yCI1Q20zp5rpXZg9ykvG70GAboWEYNoaFOSVjY0Z55ETKdBvYYXRKB6yPg9h09tAU/+ql
s4yYZTuom2k4EeJIj6qcN2GCNMAJ5uKIwIpXJZPJyqY/VDTW0NMe8cJPCL4gZATRUHdgX/k02VcW
/gtzfB4+E2E2ilTPfODklORUfpWs5DO4+W3f4TjQW0fIEHXfnrHhmQNJcOrtlJJxfNz6VbilaD7O
dL0bwt/ndF1SBpyAr4QPGXRCs7pFKf7+fNK8ANCG4WHU2srgXFtFRv4ppDoBQS5XP4Kkd2JGo+8/
nLqN+hhHxCAoqQgSge2kEco23gCzZ5MJzmdEcQBzDOI0V3ML3+vpt1FAS+pipONTesMSEkkwLNDN
EKATHFUhJTDEzGVIbZQDTwB1rK4vm6faf7HJyajjRVEsWACiaVaZDjsGfxGeqbguv8zN/OzfcXtI
Sb383pgwliIyb/zst33GVIq0FLIqrWxie1R2nSyHcpba28Y8qDiQZT31KEao8DZqkTG/YHbXjM+k
pqbP3/0A3xdiVhnmWQuzH9k8a9CTF4iXbhc8hJuziabETc0lXKHHYk1Xa6EAGqztrbRcoBxSHApk
1p4kL1MpYQinZHJPqmgk97f37ayLWRMBSQzOcIKog8dZU4KShAMA8/qVluwyQhCNGQxMtX4o3Qah
6Hf8FfahsowQOYZX/OS3UxCvPZQVPTLTONma1+7gCU6ueJB2XGG6RAn72oaJ+hZGr/sPegwcQ6b1
Q4m+coWrQr3oESheBVBMvvc1YWZTvQOjVaCaPyxGqSD1omhtNle0l4HjcDeWb6ly+a9MR7cixR7+
kOf29cCjNpZwXfGUKvLbeSTDvbdKa7C7fFq3II7BJKY3qIi9/KCFW9vFoPWRUV9CwnnSX6UTNs8p
7JoM+lwXQZZNBCVhKcrZ/I4pDmi9aIr2/daOxW/o+lqOoVVYRbs2PfU7VTIfY4m1DJqhBElCZYsQ
rF3n+TezwL5ahX84hefPjlytFL9Mrz9Qs6wecVi5QSfYkeZUVfXGhwWVdS3vf9gB+qk7qUDcHE7x
OBtvdaQRa/zi8PbDVORYYkciDablmJ+fwODNBuimeAH17iPq8sq0B1/L2tvGLBfIq7xG9yW7uuYT
ZBwgGmELXzR0csZzcFsCwmE0dRjKJrRQAewiiZClYwNk2IUsfHbNda7O5BDzG2eRl/ePpFCKu+fr
hOEvYISMwuT1F3LhQlTFlNnIO6FH/HflXNUFSFwQAg6vjZ8nKcpme0rvnd7JbwiF+lBrSDzHK5nI
i5cWVmmWYtVNDEIMQ49zkaXpn8mpWGASYdTpAALOdXD7JWSG8K7sAVHjFYWxJSwEQuw1JJPzCgFB
QEkx7hlaXHa+JTJWHi+G9jGXoC//sYrD7T8pPudhUVs/Zk+5taUBhHvVi0PY//y7hwdazVuDQXn5
XIHd4J9n945vC2Og6BOXqvl0rms60Y8o1nDAZCItE+eu6sIDPQYZeCC2SOzJhTtHxHLGrTSHrjnU
PyDiKxo5EtfVfwT/gAkbXUYfAhy0MbJPTCmiLKBAHQrMwtMgpczbIKfCCG/IYZ78qx91j0WBKNDm
KUCRfORFcKmIRDY6ufqH60dgQf1zA33z9kiYOhdhlxI+TVlNsXlbQcMFOT9f5pWEAanHYWL3f+XQ
BqA3XZm/sIyFz1aOAOAilMM6SPXjR5ErM5R4WDs8ddtyMzWDQdTthA8mR2TF3T4Q4D59oYy/qMdX
G/KbgEv8NQpTVNMKjEl1SI0aPXRhVIsQdLYGq7a4yCmJeYavsCOKQcwI4YwhzQyNVNbfgrwUzxNv
zAiCav3bpZ2DkB62xW8weln03GU8U3rUUCDTV2srhyi9dfRCQt6xpNnQDThKjc60SGJLYB3cvsAg
X1xpcHBJrncLYPKFcIUArXF2DE/2aUXyO6zOhmk8irbKL4d3idVF2ViZfelzay4AGj6PZ7pkbLCm
2fnrFebq57lnYoMZotVnSSqNNYsvZtGxvudEBbUAO6s5SLmKGnG//G0z53+Rju4PJ6Trgfl43OMW
RkNu36VK1d0jcT2rNkKXvLKRUpW4xwBmFQI//XoWLhj8l1Xupoqk2HcwdH4F0MTqe1gWcTg4CATU
UqNNw06YqRSWU18grxJvwiB6YLdgEsOLCM3M6WV5nCDh+ayqfgwZ4m4WEqw5ZYNeVHa+oxSA5rOB
/nGljwUseJgvfGQp5e2WdIXWRdfV6CO/VAehwqoHuKFQL+z8cNXK8W+IC9ThpUCQv5diz6kL+sAU
lCaX2EA9gjQwKzzESfVMoWkbgif7q3SQzqxXDx/Xi+oJ1l1IfsuTfVde+i8SS63zFNjp+DSm1DcK
GVQyq4LKpwU8VG9Xo6UsLAjd35h9qrSAcAFxf9AWo4aVhysSaOaeYT7iX995Lu4qnAUQpJegcBqg
bfNbKxSpFtbzCoKfXWwJbx1A9ZiPkXCzZ62TjNcnCaSobqbh46/vxDh3WNf3q3ubK8lSSdkPkugP
GmDN0ZjhQu8zIGH1V8nuxSDHKF7FUKDnXW2esgNaH0mjMyARnWEhWM9yPng1KktyOnDpUlTPAOnJ
aSh8FpzAtSWnzkDZag0O0WdVXU+iMeLeZIhzGpI18+Aq5ULRZGbCECy+T4BFOrrL8nCnn5bByN5U
Gs+zDy3bNQBZqoCIsHnQPfnmtnG04Fnl6A6PclljYitLhXoFMjjoo8E9FUR7hgXXIIk54lvZI1gH
nTjCgdoArbeHnasrI/qVzAg+bcb8GdFldWfmRvcrD75Htm3gX8OKEaymcaFfQAPYsCjA6qu99Dc1
PGNKWVY8fyppukM+7meRa/Pfv6L9yQHw4XSo2ss/6DFixW/PIJmB8hGGLUz3PdrVBcI7SM5D0kIQ
/1H+OquNk3iRPxjZNVivUdOMCif97PSaflT4GYfxjLNUNYf6/lIwESIPuIbvNGZSR1P6kR6UQ9hL
n4qh02fBpdoZspN6fAw76HbLd2osKbGiH0RNDuQtDth6kRm2ImWbRDgCCEp99KPZbwuDb8SernHR
+XMDCoUnnnxdYG+49Cf+u4/fuvEcN+27y2T6u+bKTQtdO3E7WXV25IYsUw7bFCU65vs/4UtcOm+X
gfoAP/gOtAbmBH9BhEGYnBYdBdDG9ebH7NUWWHAsmlwLIdgul40e6sZDfuh79uNBWA5aY4/LU1wr
PUgVhFRqFo8MidmvO5TjGdT8vfevxN52MxIsUnxG6OynmUzRMqA9B+kqJBrUqLfwbdK8luAylkEb
P3ezHb2EUP6QpQoz4aTwmZlcEUpaFTOzNWh6efG6cIfR2G+qJ4UyJ6TZA42zYWGG1E+Sv5qkvRWd
L3xCIeHzUPgWfSzKT7ktcf8J2gnG4kRNFRF2gSsVaukPeWsaR68DpuMuHX8QTgcUBijqaMqvMBpY
8tkpjaMg+5BthlG0Ep6BoV1bsJ3G7pcTeycfK/U6+b8LviUBaPvomwcZ/m3Dsg0pvTqufKoucIMW
0PHjvsAMm6JntRlbNGMOaxTu85O5Ma8Ko3wbEtxzMOrqjDzadaDLa7MfWNXX8USCs6fbNqBy5ThI
6h4JZtK1tJkAqElqw1vpsTMgVwa59uZDh+P3LOL87cW6HTfMQ14RSjxr4MCBS7JVVLK4TUUXAl+h
HFzDC/HwiXfkiTjrz+3V/q2IotTCPoOVojGwuXuud7rCEWWSaJLwEUDyASJC1t2nnw6SGRs4S3ue
Ok5g3EBnZYz3UhkM1e8VPbbezjXbE+VyPhLSiRdjZFrufbMcELbUvCbfdb2eD7BCVCENIg0UPYe0
oFyR0tiF2NMxkFxPdjIrSpnkNWZdgynhBKa9rJi+JjYaWHWr7OooEKgNLMhvvRKY2YMsr8ZTerdE
hChwSvKRikLje7jT6mHPIAPSreMqDHjPl7pUHbOnmaXvnIZ9c3Cp1tePgUJdVmM5emdr/vjFGvmy
K+JmVXz17JnDWkOSF7XLCdxQhIYcjuf3NDE7WScia1DMgMSPcBtXbSgaezFG9+k/8gH2hlCzsyiF
zdjtFWj6alxBYhZOiEXkFZzbyzRySlifmbU18cVepfzmaX6W2rjWbdyxy98mFXs5uH17scqp0mRT
NDJdRPvjlb2vbnjH+vPyX7BYo0IbqACNnVq6bxi9uizvBIQvqdmHv3nFAV3anV+So3EU5vV/L9Xo
pz6YLABKyWmQy3WibOuY4bxX5b7EcP5JonwXfn09EGFAV+fo0nwqGl04TLU/Oa56omZG7A4c1klL
u5kgvsyyBJ7F+FGN+bXaME55OqIUlMlk5y7Q3xqMpEccIXLKsGDHZm3tI6nT/WTIHHq10OBbAImD
MEhzHmw0tw3/LEN4m1sXCs4+dY1uvtS9qE8TOIzhJaYeCLxU8wFcGJiOCFA23egBrQrR9SWs9Vmp
wTB9oP9aIV5bE5uTRPAgrt+av5k9mpn4Dc+RJpS6hlkRS3s2+53nh6t/6mFRnhZLHeqF2QalKuue
Ucr7tKefdPEoRSwr3k9IDWHlcpJ0KeAKbjhZW7XF6R89YJWdD+a2mWRcbU5tXDvBUbGzMvMGzHUg
B1ROvVmbhck0Za0zjUCQyk+0suN6aVvRlUtH00JHtBB/JRg2uHEFvz+QN2KlwERDTld7/YA2gyxP
e9DP/RYfS9+D2feJ0lcS7GOf+Qg5Z29BnigngUmaiplqbVarDlGaJthvvLl2/K+pcbZYqTbIGlpx
2+h71dNdppYX/YHOWkc/7aOU9W+1xLTskR9FDvJD2SdMODeKb5L2/JqsF+CyZoPn3p4RganRnTgT
//dtuq8OSBuFCqK5ThooJ5GJz56n0vKfjU7KEQzugl9gqiQuGb8wDdfQFUTAmOuVULIMKuI6VbDK
Sw07bG05TXSgex2C3sYgrRwZwjkzfBxFgV1sPV3NCRThnncybt9BgD/unyiAMthbZibV4ZV6R/wF
hWMHxscR0pJTch0agK/6p8JDOcVdabz3Z+Zt5knXDkRhF/ELz3gWLQJzXKTAjtE3DFf5gAHnBoK3
FlmNsVzWIJjzmYcILs4I44kZ3O5xJo73x0rvfedG7dKpZGPGKJcFSpMYj8Y7WgmShofYB3i96Mr7
WfRxTu20X+CdazDZp6PsESIKAWpl0hUPqQs0gTOeJ3MwfzIGLar7AuuC2Uk80Z3RWqj+yIq43YrJ
P7iZlX4DdPrY+ju4rKfj0uyjgUJkTmA77G67HcAFaGdiyE07ZJS9Uvzm8nJj4Sf4cwBkvDPoKgRU
HXq9jQorf8SY4PrtuqYchT3L4M4nbFLjUutGtpeMqN+zd5/lNq2wGHa44jVEeCH5BlG2gHkPuoRg
U34623SO1qTVa/WDvBIC8qD9ZejqlHldY18knSglEBlyph0D0HUXF2NV7GpkAAKqO0g2fg/AEqU5
ZPmLXQJAk/wzYQ1FjYJdCL0B9S1yLSBYN2UH2h0XS2dHqEsIFj4Z0RaEHVHjFVQFsRXDqLMqYTeF
VmjoPjkquHqgzfuAONatEJhUGMKSazgxEWqtyCMn4N6Vcej64Ax5KIukL4tpoQ61kWvmOq15vjE6
OeksQ0RLtxEVGpM95ZWzpJm4JQbZULl9nJZEu+rYlJgPpYIbO9IOkaDwITRS67l/W8s/tl8v5ON0
DHEQgxfg0OzRIeoFcjrqmm4G0QzaBloorrQMgC22lXyWFrBrJAZrJEWXOk7sRlGuJiENsFxlWBdz
5qoxgZsfSQCHbcf9s9058Y0vj3pU2qxXTLLOIjwtd3BJv+uXMG+hnVTrlFpSC2heV9BbmaC/Iska
WfkVwVCzirp9RWl1LUM7YRlyVXg+rzqrjhFN95ZZghjkZVhFP7zBha8hMQiTS937SmvU/Z43e6cK
K+DUInNUlqTcF5/xfUp53yrsjZx6Dg3ZtPAeM4hfz8CwlL3jSJzQ+kNcRPyQyB9s7Ip94smse+EC
az1HVbiRA2z57A5qizhyHD0U+MewCaRv2zn1ewSNE0ZOgReoFxGgEgdDYS+MPfA2AGO6Srn5I53j
uNbBEKEPWvxwy2eq6jA9DXe59uyFwEwT9wmlcFPZDLBC4HIEPSjO7WYtrz0IjnTQEo+HK1e8r7xU
UPOqvt/HR0IWVHCioFaqelXoGt7NcuLbDrTIUdTPAQ1R8+h3XYfQ4nOljg7PMCeWUJjK7u2LnYPI
GzS1pKwZTGpO5hO9BwOWTHYntOluQrOM2WKrS99KcvJp3yX+xREwAFNbxzSkfrOKZI5daNsDCZMQ
h05TwZHbWL5Mj5I3XDNpEC5d++kSoj3zA+GX5sA6ain8Yix0lYv6PaFLocu+oSE0w4QZdaGTyl98
HSq9jCkEUWYefyhjjnpFetkEBn48/mDNkMR+A6ythA4M1ZPnfnPwzYeycMQu+myCZO6CHDeiu+K3
GhYgMWZaPpVzVTadFA41ukDFKnQ4kOqR87INOUBWqCswq6gr3Z8WdvkdIP9wEw/MpAWdSbjWnRli
Hu7rrunFsoni3Gnb3puzUAR8jWlKbWupVxQECN2TJkDZ1LVvXx0e3LBQ0342H/39xWNatA1HKgYC
Jb6nUVd8CU6zEMEmvig/zAOudf5FblnTyn3Lc1wGKvli3gkq68IOCES3sH10tBv+V+e/16TB7X7L
qxr75GJ1uSToZTK7gi0sCA78Z1I5PaPsjkX7uJKf5/dASD0wBfZsbgfoiaBG03RMphfd0WPh7B+0
8ygJjPlIeQCn0G2tkmV+boScmq6HfNngMtYPzreUbR0BIe9h8q1MyC7f14JXpDBtCftCYyl2letS
9Zt5gbsZEaLCD4y0If8qjjfp+jJZLO9XU8V3pdcMLM8dU/TMmDYvDIM7cuzKRTIeUACMMqw+dbtf
pBFR/56lf+55D2GoCzV7hjEHorQBtORKj1B2k+glkXwbXq9+qhXG19lqIrnBvhsNL6HVWCH+OxoH
7AscGhaEfP1jokQ4R831F4yE4q0AOqGwuJlLuiBzFmcf2Og0unv55+a3EtGiC0bYjRM2GqCM5JnA
VXACM+epvr96urQ0gS4EOvmv6bQ5L3QmmnthVP5wSAikEmKhX4gjYpOgkRVM1/LMXPBfrZjNKQ2K
68xyrzN8BUIEveuNUjzYOJHrfsPL3ONREVsjDtjjldUk3umYokIjqKFQueqWHi6a1Wjrve32Dltc
IQjFYz3cca9PqiVEwJTTIGb+9NgTHDG9vsbglEA+Q7wYr9li4JazJR6Szvt/Aea9uOTvhJMiQ5gj
4zBwslhGfzrUIm3oSeSCBb4gv3x9ux/o6EHnUVUtYww2E2nXdoR/ehP+p7F4NT47bXAUNRRSpoc2
0k6eQw7tHUMWSvvP6if6H1yEpidlbyCi9/45n0y5VBicXcFYAiGluKEdcq+5iLJ2n/TqbEzrwiV7
9JPdQAJtAWX7lbBfqZ+QbWqVRVoz0COs4dGKZNqbDzb3rh2phOMDPywdlTVmvWWg+bEnz4n98Axy
cnffsgN+G4UizSlWRvSQsIPR8f5dFSgDZmXoN8xDI12zl109b12Ev6gzHkIs6A41ku+dsRLAPUk0
sxQUf1aD4a1NqERDI4KEKxLI3sfV0IpptVbizvDxsi1AjMvNQ5s6tggHtmr4776mXpSNJjASHt65
S/gCeUNhwexhPE+g1TKKeWB3AiYJCup5+y8qkcAGflHrxaIZaBNe0/GlZWjEA2dWJFMi8i/x/zdU
zf5Bd2s6VC7h4c1Mt6W/YuXo1h00OMOFBe0ch6Ca8BIxYc+ZPN3YLEwADUxeKfaJnaFCouNHPv+U
esSL0nsrQ3jXRgMAOydg2nw/qdYOCNdnTD4jUADt/K4DhXX1UPcLDRb3Gvc0Ccn5KF1J72iNILSu
S4MzcJpL3dFaV5iGQP/lCoUwcl0jzmYdL9C+dsEsY1JNzq6ArsXrcWYgiaiHxn+3TRPGAa4rowc5
0GCXt/oTveQLuKTQfi23Xp4sTnsvYtyjGcsLqdbmLGY9bdF7kmdPjCynUbH0LjEUL5XGOd9DN5Wk
sE9qEQELa6HVM75MiNPzT1U1AGrKaL8HzcUHsfAkFkomsP61DSGPjSOwSsg0ZC/8tw77WbwVX+NR
39ewAcu4qqhkdITj58uoMTCq4X4tH5QF+TSws1qkefEpYZ54gJSRvcQ27uauLUamy/Fqgaco++MK
a5soeiNtrDNmXQsUVtg2KQJLXFx8Wuwq/XxyXLQ88Te45MBB2FwnFOzbGdWpL7tysBwycfv3Ad9k
GvmLAFVvNNBYj9oXpIT2MGdkeoOzhNl+eXF+Ys85JXEZqVdRwvrwOQHFrmvMsw670E92D5WrOB8h
q7cbysa/p4jOPRJ+qqiwO2HJQsvrmxDkgM4hOPpl1sZMw6LXTq0B3gNEzB/LutSSbGOVuY3UlD5V
XGdfUm72U7E7wZ7Mjpslz/RneulINTeDbX65MIEt0aQ9PUBj5b+zxVGxkGK0QXAIva9kGR34Ajnh
aPF442vXLDGCCQw5iLUhfkzQd4MNAjs8Tzae6FPU6Y6NAtBXBAWTYd7fD31bZDtT24ynk7hwehOW
x7/K/eTq/BwLL/Wvp62qY8U7asvmOz9wI9g8CcWgm2EesfS1BEWgiNVwAI+77R8T6MCfylGQDyBz
CByhW619jGFcr4g4wwVedluTUGl3Sbo9IF6CM6u60nZ/OSqb+R3koyaZhvyaXzKfZGcgnZ73XrXk
NdhG38Fy4L8KQbu1lZ6cZdwj5YUibwTZy857En6i3fIyiixj7vUkYHz6cDsygLRjafs0Rq+6NPfo
IwU9tvja3I64Q7CMeGebqBCloNL/XiadznjJ552XoH6r7EXa4cMxWIsZyoGqZh4xibA326ND+R+E
Fkjtu2wMnB9TDCsmKsoAIeyyi8j9dlTrI0kjtlUpwmOgMtHQzML2h/kw4889IyngtokGXMsLcH7C
UlIZRT2zVbakHbDPuou+bXPXtMa1q3l0ZviayKwe1rpZmwL7TCnNImSQmh7ogsQ9fwSHd61awVmw
HsID0PFK4m9nNNvaX9sbeeKBsHjlukmXUWn7CFF2NGmEQZwyuXDbguDwjwx5/W/ArSozsOt0Lqog
50ztx7ro+u/yO+BXyKVjTLMfntTjqeu+bFo4++qdcnEqXBkJ3KvUgjFT0Zw10hTfVQlNaWmxwqA8
aXPYgBkvg9Oj0UQ1SLag1jjmkZyfiibFq4cK4PWytlDkTt7bDmazQl56fSSzrlzsyHcPHtca8xAJ
TpBE/NoTihWWc1x7pMqZ7wadVRF1UdWVXFBolHnFquyJfEewNRsoCaee0hWvuI2t+JkeP5iyPFn8
C1a2qjFo5/d4b6XgmLbauAu/dr8O/e1wTHAvVS1eJJeVOUQKiSHU8zKIYHHvcBcqPdVnsvt6lEt8
oFgb4k9Um3jp5djBX2/XmgJL2ll98kUAuv37wjl/eCvIC1D87o2IQkEpTCbC/FyPhCkC4Xm59ZqY
uEKDALCEDBWYcIIob2CNtK6Ue9BqWFM7OVQxeDjGPS8dyXj4AgfBTwC34RtT5s1hhCWLPKXG9f/R
ECnAhuwMGI1RRl9zjn2NhQs7NqDdJEOICfkoyKzU8SFoMOUrEwy74RDMdVvJhlTClEGIF1/0Bgla
bvXXaLL/7Rli5KBH3ojqnwrpv8NG0t4QosaVU5swH28S71RLxXgXUflbGKstP/eK0rXh0qeg6BI9
EZmvMKJj5yFcjZqYPdhFba6cnr5wvpo+rBd9VKbgSnSNPLXL7yj1mpYBuUtjcoWecsgrzIsebZen
f6pHCEa3UptsqgA1D+/Hftvff1fAPG5KI9DJ0lVdNR5jUFICEt0djmsgMycdFb2skXwA+jNG1Jvx
0uQ6j+zp/DwcPUIo3W1Z+80SM95nnK3lGAV0eTFvzotghUjRfZwycMXghqdkh5EZwbYdqZQsx5HX
9/mXlZX3S5Tl3jxsGIZ6YTb3qdbkk9JnHC5EbkoeZxjLW6NBJrJYPbFbvUAVGw/RiavLkfWieWwW
D7HMOHTQakDb4ckcj/3cUqalKO/jmZKFuA+1XopzMAbe11lS3YutCyuwyDvkcIa5a7+6Vxci+4W8
28PXBHK1K4L8hEU2SB0tvUPBIrRJgPppcHOTb8HhBWGYSv4jVpFv8hoPJaQ1GoxQGlrEJrxNyW0P
sEkCH5dBWb03CO/M+ESPtUcQ8FuibhRmjtLCcispcIaVm/h5ju4ynJpHIHLhCcLD9/0xKCyYFhS+
tiw+gDr/Vd6H791Y/CGNrIlzRyKbOrKro5393Zir833GcEAq4oRXUJm5f3aVRkUS2+8rYAfXIIe5
J28jF1irkiarV1mpGHklK+XxqKJmYBD91WN8BnpmTnG8bJIBeq4rg6Ra6Q8Za+HUJ6xMGGvhq+6+
wqwl83db8n2VeMVicn+En8obIJ/4z5NwK8fYl5VaWZdA++RNEsNuu+WF4EhtUNggHrNSpi5Attoy
D2osUNyvxFB7G34Uz9P7NvUD1ZImSYvaEOttgmTS2/7ew9LDqR6EAEcoE89BmzUo/Yf+gVM8hsQK
xfSLQ62H9c9N/3iQQp0qpx3wx/INtcOyHNwz6gS7RS2Trp7oguIlSS/eVKvi7xQ6aZj4cl8kF5Sb
Pkr2+T7EJr9yocXXr+SvfpGMyU29wGy5zo3jBRg+Imy+k7OOsBENSrEFotwR+5dQqgLJ2F12nLLT
BAcL89/Qo/JgCGUglXt7woj4MKl2dTj9rTI6IUWt97EhYdHAwptjF2HGVPRKSb8MxX0oNl6ZupQC
orzC+ovnYmeM1VIDfXOfWfVIYEQ6s8wFTXHuHxtD0aXWO/uwyjY1sRygwSfCzzILgWh34jDHvXbR
Scdxeo8EAHsMJuzS12XYVoeIukY3URyiwX+Ah+DDlQMnLAs1UKrR+57NfwIJrAUJa0SBs08Tf3T8
9vcAcGWIVF6ei9D/ziynvFIuMpsyx2/Kx4n8JAUWYSvxPF0xD8SZfP6e+Hxis8jdLvRYSLMZziz0
L06zny8MsULL998n2mge09VVqgtUqVY0nw+z3D1maacwbl4WVDXPAOTzM6CedGR//81t7oGWEVP2
ILD6Jc8k+6+U1Vkl0bc+P4gA8cI9Ak0/WqTMCb/v3yN42TfZ2gbXPuXPMsIwMe90aTerVKSUKZQ0
FpKFlJBt9NYZtEWPGPMuvXwnWMrWnO70V+rAM8HLBqE419UujpQ+O/jB6MsRf+j+XSm1fwG9/j5H
xQ/lBzbQ5HdKzYA6s7DhkVL4G8ZFJn073RlpsVLmAx54w0kMMbzOoTyesW/ql9wlNEyNeOKhvmiz
snfv7ymwEBfLGDrF29bnqXOqnK1skd83uyeNZoKeTalzQWliheYwHwT+++sfdiNKMeNs1P2qG+Ov
7aupIva9Ae+w5fc2sBHWgE8en/uTJz20aOJSJ+gpHfJKU9YGJg0eZxN3IqtBr7Fet6fAQrvpGXZX
+Makr3vV7vA36hrmFcIQkC0a7aqHRFOYV6PZrTaGw7ZBVVo7ZPc10GQqY2L9tN0wvegq64GduFgy
dzEChQShlbq+BvBc//uiEFL76OkWZeWBMINiKB+zTLTx2e6ZO79ciyIlN8zq4GwSalNyMcbpE4hA
fN6Fkm0LZfqMtY0JzV11kALFXXAgqFhyffSciMkdf6x7c0GAhbYCGsjAR3rKmXk5mAzfrvSa+BHL
PT8Kde3utvggfGlP7wlyKiIK9G4Bx/+t6dlgICWnf4BmASDRepBGR+gBGeZi1D3IRypAudex7mp2
fy3nE9lnMLXh/rE0Ua+mgZQJHsXTyWslqv4ksqvJFk6DIyRl2Ib75543FyTpV7ECb8WmNW+xM7sy
gI2ix2cGI3xHXtbSME3nuqBheIhrgEAdLYvfI3JfpZpJty75U5T1030KcbceNyNpF8TVJkADUW+e
qaKZQV0eRz0rM08gKJ4I0JPNmeDm01Awclp+YEKqzLmD0DiVUAfI99kWkHfodd1ltSdtK+BfY04V
grA4FCFKFas2RMK7yvOKutJOWXgQui5BVjmEkAhAVbFoMFbbGahYIoWCVO2cme6kXmAT0jwdaBbF
VhpBcN/IbmMouGNChfo6/X73NicYKALMqPg2e2T1Bm/IF4kOA3XPKnqr9Zo39wQ3cAsh3l7nq4lH
AZRMMyRgooG2XUrI4tXJlzqHcvDEmiXRa8EllVKpZVwLHnqW07+IHrH/XqRRywLQE+M9/wPExO9A
QFq5YM3dn6GXtbNct7EK4DhSIsqUjyn3X0tGDmPKJR1HzxSUK5uzxFek1xlxvD2aOq2/7uviulSa
2FIp/GCqqR5vxpMJPNZ9Z1/VP3bc9a+xPzWxTNN1Q2MwpovELwDHDtenMoqYPyT1s33KltOHhwxa
fE+a5eKLuBUIRFlwW56w3phmtNUSOthPFSe5hsGr1IY0z2nGX4b0rfaf7/0XBkrcj/GGMeiJTu9L
EtS9xfei4/oDSQf2V6sbaoQ2/VTYdkGYTsXe2F66f1fgjDAiI3bTVsjs6ZROtO3TaEHCyfq7fvlp
hQnCJGEiyPC0aae8AVoJqLC7qrBxaknXAcRDnARhUwFyUe0s/H8BDmiKfx8JyT66W5KpOYJhU9UX
eoiq9hRfSblOaOX+TAEqladw2WNpw32DWwRj0Sk=
`protect end_protected

