

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
iEtOB5S3Q/0nxxj3yhZWc1e9CYVNx9kxE38Uvw9Q5GTpbeWA/PaP7MHi1hZ25jWcWTCQq2m6lqXe
j4/ejpW9UA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Xuau91ineWkILAnXNctj7ghjv8v9lVNvmGeO8/qKPRA098IIoEEWbPkQsDw9y8PN0Kc6j93b9RA3
24AkaGw7vS3twv084InDNHpEnlN63djkx5ZcyOiUohe4xecSmu6QA9TFBRDs0Woq2jQD5/qd0oJL
/BaRHEN9wihMkCnRmi4=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
DukDx60lt5tRoBa9fYOjxQXcMx39PTzSzi3mfBKPNtGRH42SBSoh47iSUDQLozXc9RVtQC3PW07a
TdEl+U9LI0QpSHNQLVojqhahZCfYOg99dtV1mWPojzxtpV99k2zYX2J3PXN/YbIzV8ZxTpLcq1Jp
CAIcrPJ/34KYVzvzXFRsvxEfk+CxS8lIGg/nVz9ZI/SFfi31TG5Gc9nsiydQV6NxDLfMTIZ9geQt
WjMt/ZdcVbixfIDM01Blr6PmvrTG06LX8uxL31TQuw5SZfsZBAh/PoXSzsMleljAYXIhMhdSUOnh
qfkHi0I/YHOxbZGvwoECi6yzPk1O8e4p+mbfJg==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
JfFouWl9C67kV59ngW+xbX0i0eu6h0roaptqFtm5oV4WYkqMJEDqBwmHay9e7sJ9CO+K40RDFIJe
/eeImbz2XS0Q6PwgmMgPAHRoOg4fHkGIAEugmb7hj+mXvk7iQo09CaB7HocKsvGcx4nu5U5a1pLQ
6UjYczksNjCCieDaJQc=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
RNy6OyrkxjF2nMK7NTVKf+mkYRQZVhnkvdhxFI69h+pJImlNAm3GMG9cNkr/rYPBFr0KpngtSqYa
zub6qdQpsLCoZ7qDFdEc1+wws1xQHHeB7VAyyByyPc8Chu9XZcfd6cEAYC55a9lNvtmKoAjppEfF
hj3OtTTwZQDicoWmteMIzi2n5YcjhwpDSzFHpmKq+NQje013CABovpP0/TVMHv74ZpkyX30HW4tb
0iH2SzLvUD7U/AR0ul2kht6wcMaLE9E6bQipSYn1DEnfUpMfQgGpPJCWjykHayljMFWfI9ucuNXK
1XTo7EI77uCstdWwv1uP3ZSQ8pFNDP7NXG8mpg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 9552)
`protect data_block
xoBOfNo7GjSs0Z5LmLib2e6JmgAiLdpuKEulkNHBRFWzT+1rqLFWP2/obnes3oFebaCXTWH/e4bE
0UQ6sAOFKY4EQm3Thavx7/E00GgNmnLtu6x0affs+ME8zSTvjDTj0jfzp0dDGKnAAXfowlaZ20WW
YNPsavXt/R5TcxB5S0n79Ovy+DLY4/Uaa/GlCxJOXp5LxsfQDaIqhNmHB6CIR6t9fv1zCnMGnoXX
DeYLuVHje3Do+EG83BJInngfRk2xlZ5Gn2yuR7R7bQrFaYZ0GMRd+VDU9LekpEwfeNXrNhQUkf8H
2dtISU3HnkY+D8aqkCsLOY7TAjYt9moIvqE+z5FkqsFR7t1rXkaU0g36YDSKxXJM5uTs3UUFk9Ss
aZa47qTHTGAQvg71k60HSdEaY7EMbXDztIcD2OtmEusSWlNwl7Sp0iUCaILIm+QlGUntFoCqYdGe
rkaaDFg4QwIzxdLWhhMi9bJEgGK0x2u1SrMgHBSZiLlJG5bEJDAoCMtXNBmyXC5Sn2OunPtscnHC
KRMCob806Y57yZmkTND4ZbtQu0KDtKzSKqw5DgIsunNjJsZNX/qVC8t7KBx/ALpwYL7zsJUsrTi9
TjmDdWYd0Ph+hykquwp7fpZzU12nf81sPAVFhtfatoXEMFYS01pc3kef/JfA2yHq7VkeIYRPYwwD
FczRQjGfbbzhaMpu8zaiMgpLA8kUm7cjxvVymYXvNfqr5Jyp5TDwOWceiX6ie3o1Fce/Z8x4IZmn
Wayxdo0CHLkyUEyOkH7o9NP+vv+Qt3jdYhEeJ+bvNRBrkkpJb+5mHRSufC3oEXkd0IXhuDfLm3g1
JmFw8GIGpRWu4stG6TFsn+vwlvbr/19x6ax6P8DZU5GZWqTrdLlWNpCnJWjFzD1IkaXrLVxrz8cb
l4B3MyXHPnoLAB3VSOkQBgN23cA15m1HFJuU9zNvR89d/sTUyaSaFrGZWcmBLagdO9O/r8mcTpQg
2y95cBXxA+eAItwNUsg3IDc5jQ5OkE5vSFHXPnSzEayQ15LdDmgwF91fP+gtS+6WkjVI3oZjcliM
S/xYOiafeJWb7Ax8tG20VUMotfitncRrKLbvIVca6uEYyMmSEt27ma5usfGu08sd6kOw4aAy+cFU
xJbkwhIezAcjhbth/5UrhElbZ86l9QGk8r0qgpo/NsuOzpAPyhm1SihHT9m7tuex2tlTLY/quj4v
9fQtNyuO79kpBtfISjB7CaY7t+C3ajIQJqGWr6Wn36MPbvHz9kMTyBnGffAJ+foqoEI/MA0bL8kX
/oO+OX4gppyk7JTBwBQ3NDr7IO+sDsVRZZSkewq74d20HGULpPxe3ipQ3W3zsu0u+rbVp2wof9LP
cFcOJwukw2lOrugkS0Uqo6zzVpMuiGfZZvrJ+BZn9G1tpKYVOgveXCgLgd/JlInXc3ls7ibhVEh7
EE26ab1ZfjpaRQ0mpPiQcmnH/lnXvw3/URopMMickixv7DoldEka9vMI5UguL/O6IMFs+zSK2kCr
yqRvBdHb80gJqXo216uulFseVcGnAEsFuCS4xY+/V1Ij6RT/ruVdfA+FcCU3wNaunjGn7NQY6GXG
slxc/fo6z/UkmukzbYHAwDsKiEby9A+guINaq64PUIUgppzYF6sHkdUWoJIQESR+qg2j34keHWyW
tTobInPGWH9rXtL3E4kVN9KIfS/0vbiz2BYOM284glWgHKqo4gESjHdHRpU/0faYlruNAq3tf3PL
vMKaHGBaZnqdfiXt37NShlg5VZmI1osUVbtdwmt9C9YwiAzcxpK8oi0A+823dPONBNDUaWGl7T04
HkA4ohfw0KEhOhmzqSHgWy0hXgwZFSBWNIjwgPsvo7k5q9UqNLH64d37+5XYdz8mK1N3ko1a1z2k
o0d2q60vMYuK/5KVDZgYpskXS3BE7ogGKlkQmwwMjIb6JYRfwQds5Y2nkJ913JTNrZtWkHTAuP4C
Q2Dzjr/gFSzXYhpB5iYWrIgOI7vdfCZNGwseS+KQsW6PBoj2xuRGkctKe5ZE8nouE4FXIIlSPKH1
kfS1IqDw3mve2LWQvHf4YL2ZGRx4+B0RNLbddmWn9hae7DiwSlDiZ0JitVtp0kjWuV6fRO6nBJqF
HuNenVFvXIIfqcv+88fTYulntqtOLbpzEwOGEoCucGxBTiRNmtPU12iLOKfrE0kznXvgyAqc/yI2
nCsLbnK6ZPeNCUe4o57fW1SUw/bUgaNMRIWez6k4ENsssJ1/y30n/OPX1Hq4jiB+46E9XujBXmpK
3LTk5YD4RrD5KhlVBtCPW31wHXnLjtz6+1IYpngPNq2M/1j/BRbsJXCQnVxCaqADnTyeqVxogs2o
tiyCF/98bw0haeVERYK8bsUKDRZgUgrpddnfeAoWa2WdUEEgIwl/2pXf1hLO47VGkGE16QGrHLUO
R1p+tq/F2AQaBDNkLvwY8gCLIVgrQvdJJl399cAnT7te/LYMH/6fp7WCGPe2UD2k1nmVS2NPqvId
O4f6gr0JRlx6wqyTuEzSXSSe97cWdaJfYp5ZmX3ciVAuS3UT7XLUAhgwnEVU2mVpBatZyKZuz9ud
/YcNHTucuZLVbsKMjA8maR+VizRSap+qtBnBwnWBCtX5IrYq1lGpPkePGPHKcqdMcuHPu9b01KsT
sQ4vdnGbwAH0pNUudM74314ZcfH2dQ3xL2AIhqA6t7TA2jZ2BW/5ZiahA5eeos7AtkVCtBM5uAN5
yE/anUf1LBmXuGy9k+4TAS6yLDrRUiSFavS23BnZxgq6y9JMrf+lH2IxDzTgyK10c2IXjE3hLCx1
mNN+5yKQgY23WA+x86BU5NiXiQjTTIy5v9GoGKVjvyhkDF49/LHp8NqMPGNbg2sStR8Os+RhMN/h
nAk08UYfeI7ghol+aiec4eJ1MVoHyaZ0icPpJSxTl9FpGVCLjlyFVXid/mPILD3X+jet/9FeRyEc
iHx3XHIK8YXx2L4rN/5t9zOR9ZLl/qN9eyQSXhCIyoI7IRG9n7AtIzdQZTREE6qmMdYDHgGQWFHO
Jz7G4e6RnLYASTTW6bme6P6IH3egRrOStWpTDkuljDF9nsz6dLcMlc9bHwdUizIQi5I5xZCSKjyk
A1I6/hKGvydECnH7CKDe7VJW9ekM3ATU6kTKXFfXevZ8SY+Upk51+vDOdXVFNGB6Ag+Hw+mhxJL4
pkQrRDD25LOcqmzHmG+972GnoOUEhUU4zeaahpzf4ULXxTlpP95+RGdAhfYiVkOkmMiP5A2QXNY5
uWblhD/ng9+/ysS7k57gYeQMkS4kkfNWKifmvgiN32ty+N4tusmhdNk/vaXp0w+CCIrYzN1jgrIg
WlDjEYtalge38TuxqETCAeJSqa89REWywo3GDt49oCgBctq2iVa97Ujtepc1MDbDnANCWeMdOLYA
QG+Zh1lYY3q52BjeEHzs8FL0qhIHfBjGN4+EcuvAyf7DG5mHKtLs85geudMw4ytwrf5YhuKdyMF/
1fS0aaVEe2JCbUQS2Olt0aSCVbtJhNEyj9cIez5Lg1M54tQTNqWc6HjSTjOfhOAbtbxXCBw44ZT3
Bze6xYiW4A2ed+422O3G74WGl87HPcr4zX/qtKJa/SrDIgz/KlUZqu1SAtsBPdeCP3mGxesUmupt
Y6n1hTw0YgXMQndqVMMgp7KAntQR/FFxylmPoLfIhlPLoflJHqnk0B01+24oWXv3a9UcRCW9IoBJ
snOWniuCCZ21PDFUjWIpZuXZ156KRz4ipYfutVJKU/3Hjj/Zdp2YaA/wkOVpwqBm0FBer+vSB0aH
lpWFNsTlylMc9rP5Kt/JR6pjHSAsKBcYX2g89GDIwCH0U5kukR0vRB0Gx2dkHAjo0fuyELo/6QOo
s+ah1OX5MWX7WRpKsTIY+pZDjkGWf6Ecaijb4V/kFVRJwBu7GOeEzz0CV1Jt3dkBCPgE6nMh24G/
mO3FcXFIVpM/WMxySpRdVACzzmOwZyg54WAfqZHAUxjkkRICCIN6oP4VuwMwpWE+RVYtb8Ruzu20
Gqvyg24ZS28XNGEt4goAMOCpuejl/jsyqZdwTLEe+RAJ6spQAm2AwjBu1cvUGvLzdQOxXTKOd18W
qT4b9vdgk5mV0zirMFCEds4O9xiUKp6gZOB5auoW+LaINCVSlSe08TbGbT3qGbW4y4QkfZXuKeEr
si9NJENRAhGiRdJMp6Cr3nEl30/PHshQRYMkdFX0nbWkEMXGlLfuCBtUUN11YU3oVxpPEI3r6dL0
Zdx4BJkF6MOGouHlcItmWWaAQTTYmHS3jy4J7ojZUsthmorTgSnnxtvwwjWl8+bqpDHZLhsdiW7S
23pFdHrD9ts4WuAVtvJHAMpdvem/3nlhZYV6oxJX/lKcEO/Ed/YE443Jfa+5YFyXDGyD0xSL7l9K
t9R6Yo5WYGMebhFKqvVZtd7ggCMwFwV+6vBcIK6CDeWgVTwQ37t/8imgoI1qnNJdsoDyQ560ZOZo
k/HWoH8rLgjkF9A7lEdruqDJxrLpHmzDoWcerfhUp8nuy/UckgIWw2Z84O1O8AKBp5l7Y72B/bjj
kOeefBamnD5FuOiKXHo2TUSzSQ2q/+fByqQi+WXPeIQab2k0wn3udPy05OvasfNC/SZJMHpj1rMO
wzqMdLEs4U0Y7Nw1yE2PeMe5HTYnE4GRrBqWqVHSOjVkIixHJkw6qPN/Sj9OXQRIBoldnyx17oiA
f8UMmGxSu+K8gYkLtd/NLqcVksA8f+K+VQXWN2raOmMpyYum1UY27GfqR7NR2UdflhZ10ileXj25
dsm6mIdwf/mGj0FFDumCixq51JtcWjkGCGo3ve8bcecMnJ6HbAZ+vg5q/uUqktpN+c5XNgC4eJ6X
S5r3VCYWRqYXpPqUmweH3VHQbypYNPitYOUP7BNE3pmVcPwGTvI/DmZiehFt3UkOGk1uEDn5gpb+
rIISiVdwFWh7I06uK98A4H7EW2YKsBoU7IS+q4vZVjiVLDWzijjjopCeI9cz2f7w4y3THbnMFgoU
yZquuFWKCDQwnavz6nKCMWlnRoYmbILdfxOnlxDHf45xU1Qzb2ecEvBu99FEdkOkJUhKEPrCyM3L
Rh21hENipWsVZTa0vHADVPCoxLj5fTGHRYNFvhfzQ/LMl9e7XwLF5S4O4NHo9riqvDgQVjmMKJDP
10N9K6iVBc5rtc3LYO8bJxsbxxnoSseWmokIlzTSjN/koyVchK+tm/M2PJx4L+Cu7JGGbFjdnRgY
l2hazPBCicA4HE8DqcOkXD8Hvzvclv8+GV0M3duSI+vPW0siVeQAkijbu8rbWVAcIzBaXpSxZGlE
IBmYqjaNiUM3d05ag4RTOYQZrQiAw3mwzoOL4FFGv1FRCHhrH8I7eJlJwMMre6LXI6Xg+xhWUAK9
FVx+qNQySP/NRdgmsxAWTxtU4CSQcl+JZFTO9zvEWg/XcsbEkOlcKjeHupJV4wTFZsf/UiDqn6m9
/cgKt2yS+68ZyTaBrqlD1qVCZ+tm15mCuVh7N1QdzU7xOxFFrkBKjg0JkBdUUGJtinStdqFL1RIB
82PzP9U4irzRA06378FJTRnptdAZMLFgpgbqTVghJLcNwZY6VS2oaG56L4U3K7igyBCfbfhCIMfy
n7EeyJyLnDzPK26/gpP+d7MwZ2cldQ0aBwcIY1ZCrAqzG240wvxozCvk1qYmlT5UYo9H5prOLvJP
1nLK4dnrHPKRsFU2gCXvijVITN459+WU2/w0FZStOdzoVMEVz+T07d/71cHF3rBtLzFLCi7HxiRf
eKnV6uY4hNwHS8dYAS4uvs7yo3YgEP72+zeAQ54BhYLI8B+gnjDy+m+uMpPsWU8e8NlDoxdAqTD/
mIeODJN0T8ipzwP98Trq7PJm+pX3/b+SWH+NLYOJgd/l5lXPw483c/h6j6/QszM+qbtnYXPn0IxS
Gx7QKzuJg+2Ml21DerrnqiV9wNKZOrHJpXqVoAlXABHCsngY9aVOJ4DR/P/9dCnyxMSa3hTWPdnH
pFMW2Wtf8yKOv6+xCrcTCu1otJm67aTQUgfcVg+SwAE3swZ02KiXB1+BiJ0MVLrg8/LiwCstLs+c
NXdQP4+qEU3maMBqLNA4rrgcYwoTkA1+0h92OdQy/UJdV8qgxw8/HH0kzKoHQ+xGF1MHNPOZtT1F
EJDKhBLG+ks1RPHaOYomrQl0ss5nrvTkBlu3WapxWvHq3J/2y1cFkqxi+gYhyoFexEF8gpa62xzU
axNzSaoFodYEZCn0DrCqLEdM9zjzFPG5QUMXSm4vsmiI18vVF4CGO1KZ1+LclfMA1ZfEosDmcI7z
x/5QMU+YQPyutuzNHw4eVKZe6sHKJm4ikC6s/gwjrKDiTkGFynkzPVV3Re8bjCNKtGJrM0WjUBEd
cxRWeWByc8TrbBBwP4LUHgIH1Zq+T0i9FRIKYQK/kJNSrUHZSSjYK/BOHiG864HU1J1tXrZLsifT
RJDQFEuimlcWSI+ToMy68lwdFA4M6lb2ADeyJ1/5e8ceC1BHlMLczgmUhjAhmOKKvUVFweLzgiAg
RMDHETuA+ItB6e4ZdNbmGRLvu0bD+Ch2lptqa5edgrykHR0FjvLiiPEg7fYfUY0Y9hSQRehbPiPG
Yk3gNAPlkMUVhoWKxjRky2u9+XY4pArNwbwbA6X501oaKYYOqR4UQMcd8yikbcb2QJqSlFMYntvu
dT17XiCvpR12s7k5TObvwn0ifiU0wsoj06BciEHKu9FnoQ1Gp8DrDJm7lqNjgaVjy6P/cJWAgQE9
jNtv3Dma0ZBvjrV4sdSg7YgNS1FvHit/0JIrv9/QWFFkwu0Ytkz625ivbkwO/FiDH7HMWtacRo06
tvFQ9wBqoAgfOe++zeH8v07URYH7vlIa6WrBFcJOFC8oBxidp4qY1c1RGi+T9oG2bMK8YQpBNzcg
81wujLoQso8xpBHmhAMcsyA3o4MhdII7hr61nDQeHHRQo2U2b2zApaW1IgvIOP7n2gupX0jrVr3Q
qejxKAc2ps6G5Uth7gjq3ixy9W3N8r8hEgDs4vOPr3oz8gNG6Qp7jHV75zN6E9eE5G45QwOv/Qgy
2tMQaGs5K5qxOf3sV+MzpjQiMQYWy1qxXatr5KHo8KmqL4PMEb/TednT6bj0qfpljidchTAMGpTh
vGvrZn8mNhF9F3J0BspeRlShbFx3euPl7i8GkqCt8oxex+qfQ0xWJynIR31R4w1E6ts2PYjG82q2
/XS3NkOaV7iQSh08SZkIR7V4X9mi5NlBz64n47RZd1FaOv93uS57M4MS3lr6nGHF5irdATRV/y47
yk/XEb3xwkckG4flePBNOKDQ41qw7zGx97xuCoyi1Swz2SbdGw3hGSNUpCwDLIqWJ5Bl6MszfREq
Cbmh1tpv9ddPj3YEc7MlvrlyBlFTSrbL5wcYs3MSXplWbHL2YX+polEj1tUKwNSAqK4PWQgoldCx
JqKYC9a38XWMTgs15Ae67cEtsEBq1jjV70d3a+AZwOlMdvH8T59LbIOEu22Jop0VrMc5JF0tKswf
L0okNS8kRTxxAX530bPIBC6LL4kCAwZ4MbMqUqxdABkh2awnx8c+vsvGExmzDMiPcOdDSexZu+4M
V9xBURPU+w6bjxnBzJ0V3jL0yulJ95uAK2w/JhPKNbE9F5Hu5opgPZ1RQjca/Ygu5n0d36bawncA
nDaxriKHwKo4bBG/f1OiBVOwt2wUspUzMP3//CMjpH6K/rVAiJ4WhtMz1H3SaklbdsHaQuF8kGrt
KMLhGfYLoFMxY+cOlbwkph4HqapXKngo85s10ZaG1YX4+77HUlIPHWtWcZ9zOYs+Pv2QbTfzdiXW
aN648VTOoEQk2xVFzCp9RWd/Pr2GDjIFo+TQhstuFWJhJbWAEVm6zMl1xeSLh3sIyxU4AH1VWKoi
UV4s+H5Er1qerJlo3QDNKdk4cfLUEgGZvAsNXc+eKpWZTcfFQ4eLKDQeREbia7d8YaIeoCSkw6D1
5wua7h0F8DsBX9BO7KrbDtN9zTdtg0Hm4Dv9sSxHWk2eOYhsSb+a6pV3KAjgh5PGhVbkqx7XBi2V
cDktAyXLkYdP4OaUPah+ssozAXmVTnWLp4AogllRoVz+9T3QK5JS20bcX83QV5h7dgFwZhH9OHAZ
hchJ0gPp3YCQPXJxINzPTWvOsbnm5Pf/UHTxNCJ1woLH4Yzny1h2TtuMB/lLFuXR8PjzmlMWDcMq
xbNRHBMJW+8NZXWPaOCJQ/lO5etkWTlPEQ4okYbQBlCD4EcGdkFNb3tuOEMcLVFFX0Ri0nxPTtt2
bOIJ/T0DwOA3hjpxx+p4AMFbcK1ItO292OMlGBN7pBtmDG0M9h2gfvQCUwOcXjfQxIOgn+4OYlXn
x0XAuEQoNx9epiLMslI6coQ9mWY63Kak2sRfb+3VpiqgLDBbeQq5Esf3RQjDqCSGBuNzkYK4qM7x
/X16E26jtTpcQUDA3+/IsTgOSzw6aStfBvtezOQiYZ0JGBb8onDzCRmpXrIt5H4UcpeVHKWQLnF4
st+0USAiiQQMQsKMHeRlvkqfe1qL522PJeTmLGldskUUO+NvvcQyDiosRMsgdiOPKHrZZZRH+w5p
+bC0Yq21SGxVjgtoQcmo92H4pQIY5sCMHHXzmj0/+Z7xoJiwz4kCJSgYt2Z3AeG8wXX2yG0MRpnn
w0N2wMbPmBZsoq9SbNyK5BTvHUSqe9M4ZOSGx/1fVn30RuG8prFbSXuwAriQ00V/1VIkXQ22D9nI
kOmvdmG57sqSgt9BS7i3jRCBO3vj0hKniDblBnOkxhKxqj73D+sVwLWCEAzvIwyVpAn2TpNqRnzn
vdJSFY+AEYEX9lZKSiRBRWywcI8KQNVUpVPDNSz1bwaBIFPZTwQXVCIc2CNI6vfd4OhQxYO6/oqt
zJmaRgXSnySIiYaBe2dMFXZ7bOooHJxUnyAFqm2e1JWFOGnkgW7kDhrRL9+Ft2AjohZ4+ClaSRl7
Bo90eTfpiCIYkY2Dl6OE9DqQo0I7kNeOf8iMlV7afF2q+jH/GU+4PU8gNlw7uJOAfBrnDN7pWr2u
1zBmY5I7ncasVvdtUNiEmCSNZCnNLVvoVeVnil/fdKDSCRkbunjpX0L5Xdm2jHH3DLo+QiYqSdn7
MakkIeyApoz0+tZ8w9i9Gf0oiTpOdfxwTACosXhmldOGKqDPr7XOQnXRyHmUigZM5xmDoVcrWcAH
E5OeCx/WeXekoUaW3IJvSnI8PISmfS8S0c6RQqP9iRl57Uu/P2dsti09rRcF5pi7ajByJNuiRyku
m7XgQuNCjlNpbbLINqltRhsw5TVhb6wUrccnuGYKq8AKU95AyBGcOQf+B5rhAtXE6hdWKghDmacs
VPrUDoWtXSirvI6TF/wWTIyfgmKI66Et8+UuzFFuciubPHnqc/7IN6AN12bT1sn3QVn5OY46VYfM
bvM9Wr8SoWRQbel1Rg+nmk25Z8VCCaECg8ebDMhryvX+56A383ACNAK6DxqLv5ohAeVWpodYimBl
guF80Ls9L7lg8CQYZlgJ7CP2+KNU/gN6ZMqrkww+beesrtd8jzF7whQ4o6HYhAOzZ14PEfhGEhy/
c5cSjJGMbhIou4+NtDYZWHrohylDNyVi5ppP1oJAsV+QkBuJq/7jD34tkzUi6gkCMphU9Ztzp+ur
WQNHihY052reU13bpEMnRJAjTC9BVZu+AaBAYhu2oS+6+/nlesQyPh8ew0AE4f1YXghCrGMNuh02
PWuZIT5cXx+X73wUtAjQvTvoxO8QZJyg8YhIT18y9XFxuUbNmGNUAG2zwamR3SVOJ/W9n6Ympmpu
CMvjS82eK95TBRhJgd1jDweFG0tJRdwPlVC5esfBwskXcwDJrPhuXFnWIqIZYWnZNbSNbYlMPZUO
skU61DDLtlMU5Im75QNtoZZ6mYjqK0ExpWAgA2A75vd1A5s8XxSLU3htmTV3isUXAragZbOPnJmL
yjHljM7WJqSSWpc3PFSzJ9HrCW7cVJpROopYU95Yl/e+vhzd00vwjO828nVsf5jY9tchV1IpuZrE
LJTbqmmkCgMntqe37LyX/U4o1vrXDutadjVQF+gI/2R9+LHulE7xtJvqJ8qGOg/GclkPQYzl90wp
8ER9L6Z38Yrtc1EeBV9B1piyFxJBuYC5CwQjlpgrVyuqh8vxMxZWPDqDoABFK+mDRHiqxvTH8hZ9
Jv6Z5CI0L2Gouj+WanEcb2n4eW90+0U9SJiJY+wwKnrBra6ccEtR9LEqwiiSmIi1n1BgxSvOWTX0
EzGemDMsKFjqvPoa/ffkVEpxqcgh6vq71ySCVfY31TSt8bZdQMlianZBjVXyUYadz8dGU0jJWhhy
Xq7Ol7jHdV5wyLQI2m8XLjcQXynOZcTALIeeSy4q4LHd2MHAcTluoHZKb2AlCz5yRSHMdE/yBLkt
vawmDnFaFsTSGi/M5o2nP21XYWoywrMg0+SDOtibhhHpUK0DLGYG6vtJMvqKVjyI7tdJFGQfRDpn
UNqKCwNUIy8bBqpPSGkr1oa9pITAIDdIzGaY/0/PyymeLRMC4HjwnMfuk7Yg1uuuxHWSKiud43iG
6Tw7/gbzqUuLJD1awJ0QtcIIiqOWmNVP5N160p5ZLVH8YfSfHqgA795hx29puDVVkDNbliKvxq/u
IIsasCJhp/oLaVB1SwhOJsdD0fdLoTH+ABh7wbltwhjEUjLL1e+EiWjuJiUg6irBajIQQXBvUuAN
twUfrL7LfPhj2/6CIjwbb3M7x1V39jp8GZrHz8kBlgnETqO7b6ZRcQZEVQS/QmibuDIXm8LRNHP9
64rCn+rq9PeOUudTQ64XT5BuecPJNNp6OJ8nMGG9R6/matN5bkGwDI3RzM6PkqHNrkqpDG4ne93B
oT2a2i3j8CDxRmVWytlZluiwuLhvtAUY4IHOinTz9Ee08McQnfaoZukeRfUY5O+7gAV0lzcM/FPT
SATizntVTduJlz6WYaH+WdTR6XEg4y2LBoFepFHgc3CcgHOGKwi/ec78oNQhRBmPSgUE0ye99Wz2
03r3gc/ze6tk7AzMmkKCoKVQ01h8oQaColjhItG8fVDkcuaNbG9lVKoP8foqe9l2r0iIdQyECSoq
Gk8UgB48b5vdB7dbzCMsVIXBPsKb32mC0MhbogtRlyvdz4GExX5fQwdGvmYtOI2Wl8yVMROWyHhv
HYRp2TZC3aNiGhw/aU0txK8Cb7d7V4aHzFybXAe5zSdLcD+fYAGQhDezws1rTV2lRjhgeazelch1
GGOVidlaCf9wAjIqdoaOxU7NwEhOswoPTKXWSOuoOxcOsRosBi/1jKGuXLzuuADrR+Eob5RbWbIl
hmjE+fD+hyeL4k/QZN0IJBBUVYPV6wvrY5PVELH5WgIEICR6zOW2fRY85NEMYK7YTLHnYqQOACMv
NM2WwKyurSW6x2nMXxu0AptzWYX9QyCY/GaAVq7VpJmxksno2aF8eSW14kXFI9B5tZdyKFYgSYMw
9ZC9238rSC/RdkXvNyK3xqWxiSMZHjlK9+b5PU5n9jUrCRNTvgXZ0HZVvchP2WX9C5yKGs3z+dif
UaSuYHYBvj4+94yBYIQ1lehtBP7ttUda+uKh0x8hysPFkPocPE1kKWER7HE1eZs9jJdukjscoddN
rndS8fMpS9WZgVQjWIsFD/q4Hossr6Qdy0RUCN82b4vo+EPwH6Rj14B83wJx+XI1sh1KpMegbAxL
N9+cSPaWxNy4KniP5f/B9PfMF2nvxdxex6GKOWqQscq+SbEStgdJ8nF1Tv6xU3dCYWVU0u3+2NjM
EcfbkrW2yjtLSGrUfO5uuZCqzHGamS4ksSnoWBlEyTdex7Rr61crUcC6UeUSAWHXvMZc8ytjuoj7
NRK6Asx7U0IpCGaibzCR2OjOgfMoePmpFnXY6MX4b420TjAgZLnTvHyxtDYSEMZ1vBN8fDudjfsK
/axrWhvOk6iHdX6SkQRMtqeEqQuA3nVjmBMe+Vaq2j04lq37Ucwvuc4ZWvvvDZ1BWvQO0OkcoHi6
C8cZNU8WRAKADcgsMLt1BujEtHdzk2frwUdjnIrOmhjwCELFudkCT0hocnlpi7sXGH5WodlDCZOh
s34byNSKFJLtk6jFM8sCqLuasf9TDMsxcIWUDfOsZo0doBm7WD4az3sAH6rwPH3DrVrVkymml4ND
zBBqEN9BzoZy57D5wcPe31x3hhaEv//ARrXhgEYaP6Gf4aNz8Y1qJQ+L3JqbNkKY0Rc+IQCD9sEI
anLlPSzcXdGj7aux/y5oxs4VTYCtzOJfq2ok/cvHw7cQLMRTkqpJ7Ll7NbphmjFVC8EJ8WmDiNtY
/r9okRxsHSTO6TbYoKED4ASqLnkNtRRAwHx6lIU5SYifbDzghtsJSq4tlfdX4ga2JMmOf1IwlufP
yl+KVCSmJaHz4ag+KGGNeTHvmDtyrZPv28cxfB75p6I5PXCiapqg3ivUmVDiBIj1LyhHAtrIWiAf
Ld7qGixGVhgUumb/punrEVTdMx3uFN7MmzE1tsjOcx/VCS2/iICBg1X1q+cZbG+1fDEu1YJpCAGs
EwViX/CegUqrc5WsLCA605UVZZJgAVYITep/E8yMNx3Ia6mschf15QQJxx3AGw+ePTj5ig+kg67V
Ha7lszXsp/OLo4FF5J5aM6oEfSwy78Re1XFt0NmR/0uDWGsUWMHfQSP+cEOIwHvjavsIaLgXgW57
VYLQZ5Bz+dn5Za6qOW4pQAMMIpnwGy4UmuGFdJLiXE1m
`protect end_protected

