

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
mCyyeqqjg5/0TkdJEsEEwiyDfrhah9gG0fpTMwUWGOKZ3he/dpUva8HsS4xtl5XP9zdNgeOXA7QE
z8wIFX99RA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
X35C+3C9De7vC0qODnacg9gsvk+3IzrNpqQYzh787Czr0LrIg4SN4n42C6CPfkCBLDXSXwC/eOXr
yWqN/Hj/SYBmrS5kjeF37AKShalo68kYRaZgUNEiNvBgjtaJt6WRpWYojbh+ogFdK3xIXCNq+Qxl
K0+QDwwSCDU/YMofxGE=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
n73jcH3HYbuczKsWgG6ox7VZK1YnHzJQ1B4KxEg4B/kZylbLOe/lb0i8/kn+CjmMlUuMK0WQWfed
hITAZaScEDQ3B6jcHH/bNliHMpa5PCxNetq1i73KuqIUSMzdaxGWTSuFoXR94e0GNel9SANUqOYF
vTOS9qeLaefJfWuMi23yYpmliTIg3f3fAbSdeAfef4vuNm+0XcFw60RpJQs3nrsFq9KW/GfqXw4u
TZNQUQbt6cL25X91FZ9ygQq3zmgha+CzhVMH2888hx1Tg3YKoHcpCHNpnuDfIIlbv8c/WTDMb67v
IK74ph/GlcH+s638TtetKCgz1jniP6o8owuM0w==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
lgEz+Sb20/Syw0As3tLsdRmvucviIYGeDJylwgde+NWKzNiVP+by1Maor4kKAxxHjnI5lkH0wLYs
PhqSC4UmzjejXWlU17tjRxtRz6BbrpAi6gmDH8SRbE1L1vIa3LM6opScw2kIKRT06DZ3npJLvb1L
GQYpSvbMBpeOoeXBKyg=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
cuBsFlva1Z5u1UA+GZT5hw/3RJ+t4o7i70J4gtLUlv3Ik7QI7QGdbqQ4mg46AQCjs/XyJI5tDPDQ
SIWqonbFU6W95Sa+82Fm2FOLny1XsFw2bfUdFeJCVtBal0R28pkG/kXPwJRvcecEIrS2a1k5PBE5
sZrJ66qcp7DI4wbfzpv3ic5F22QlsAxZqXZEB6lBkhSRHmx8sxDYGL3gz3qyqFuTzoFlxGj0D2l1
7IJKcs+gQikUKNCj4QKZQHmP0x55BD7tR2tDFNHuJwLQeErQDiAmIcwGhliqTf1RxwWpWFh5JUyZ
nisNHaWXl8SFhFbWbHjUNb33VdqRqkyTz+gZkw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 49408)
`protect data_block
GrkGi+IZVBO5YwKqm/kAXlMmjzPTQuFLExbLRYfPiywG8gM/lzCT0dZsNU1sYdMFz2/z+UzNq6HQ
dMh+FLjjBwwDAvrnWnvJEF8DhUuLREyaecVC7586sRcr0/0lweRzytaDIZ17YtHv1bzxQFmpvoWJ
/y8sMwUA2z5a6eoppEXhusxQfqIeW9fb+lSh0ewvidv2SOKDQgjrWXnF/K8yPadCSKf0cEVv6v8f
cmvdEzOYfjTXWSYqnXPU08EQMui78pSWFTV9gG4hd2I6+QzNm8h8ALme4ToV5fyoJyswX9unYJRX
lvxwdteF+cDZi4rhsTdrpBTOlYszYT4vDAnQg+YbVY1j4z2iYCTqZu5+MKYmJ8HGa/Uvl9hfzXk2
NjSDqnDc0vnx2yiS0Lhqsbj6NHNu9hxoQzSVqs0DGL4eQs0KizsXd8H+w27xgBdFYTTD4wB6p80R
cqsoPtCCR2rTf5GwAL8+caRjVNCLo91sTw5MOTboYOP5EiT1RLFf3HyW6SNYRzuejx8JZjY/I1sM
l2H02xf4eQ1Pz2JegzIu6ZC6TUlZvYPprbuNqUF/5pd/9fnQFZfiR4RyemX+0CJuEZjEB4X8sVZ6
2JwEJPcJ/WQGSLYmpTqrARcqu1bXqgT7hiIZKyunoysoy4JlMRDHjmkwf84S+n5szEUG/qMTj6Pi
VKDZHYpqI0W6v188Em6NVYDcaJVSxQEE6h3m3DFX49wBqGiGLpUYYPkqMl52vJLSpdjFjh46imQX
OgTFzLPyso7UIa5GqRM9pbFFI2pEwM+cpdWa2+NYUyef5MsG9Ykab0ZhiihrR3G3vufSPT91vyzZ
EvfWN77QUuW5zeXS/fULKdx3rLhRgRy2SXpK2YYlllrNyLGWXM3wOYOZpn3w6Xh4wA7ZlZIWsfAD
OjXSqZVgcgVSJG6JDrTgCYPEU6Qkp7dDBbYPD1QLr+kMNPydcidLnShAsgzp/Sv66P7ruAqAcIcS
4OvbJi7T6902+8T/23y0sevTn81YmCRy5hatsrH1mK4XsIvwNILFpyb065mPPKts/hHaWPBM8fcS
JR6rtWi5oUkC6gEh5uIz11cK3PoTDmDqyOhHA1CyM5go0Oi3mtltlxKvbE8CwWaGAEGh/+N4vepJ
MCduTLMdHSQRVq3oHJgw/Hgu5+KzTvE2Jn7l8jLEjeLXY640ADGjuaVPkDv0T5nezhpCN//iMtsU
prvNpMb81f8ey09XRrolm2H/qZTndneZ9+8M14pw+G2YOMb8Ey9KIurrieiYP83fIynnt9ce++94
vdZ3qn4wSjktZh+yvv6NxsNEjmukNX1LShqpupePOQsxV/p3wC/XeRhvpiEb6+Gqlom9+6WXEF4R
LU2sjEYuc9G2uPFWV2kx3LZgb0WiFWoo29uPyAk2/SuyB49Co51sbDmE/VpBDhf39lG+wkRRS7M5
FAay7uh0q1iGP8WtBKInmKqhRGteagA4KhF6BqmGMrhRLcE9uwBb/T6NHJCicVinLkzlmZdftRW1
iq/+lGVLPsmzX0AbnGlQZadngCgVhLC3pMVvxnHtFLYassruNam9DC3XxlO2XHa6TcXQtJ4OouYE
uxv910MKw3fK9F4DosbYDyMwAgQuE+rAQza3ED935TVtxDVcpGIfyB6ueXXSCjLu06Xe5BTgCd+x
sF56aef8yNsSI/k9uYPdf1U6wYCH0fVc5zJwI0P94NYdIFjXDG9qu4LQOhIWd8eFPqGNFcEKme2F
A9olMiV3CTs0I34mJXJ5ILw1CDPozrtORtM1XeFEx0hqtkMJkdSQI0K6ImyrTPyeH3knq5Wb3LJl
/wSXRyvDk2YkCHGC4t1wpnAOt6TVZzlr4sjiUxEFRu4aGqVa+FLktT2dIkf7LGVK8VUU1Gf61w9/
fWYDqhhzlvxcr2idz5gtA6lX2sN/kegndObdoW+DN6ol3X6yJ+nwH4VkEn+d1Ne0uO8sNBwX5fhv
Z+uRPlWESc71WTEycVi4qn5WKRDFSl+ecBaNyGYpF+6kse8KRbJMbWAjiFh+tH46Qix0LFQ1Vfg3
9KUJwB/wAXUL+KHvAvfwepsTudTxZgBK5GiAhFP6oBg3sYhRbFfcwYCrlpJtfPnOyl/kkAfqZk7T
93TOPFLR/u2/BlpF2onedHlf7NO8pQRAZUdlbhSN8iPgacb5uJqTqJNuX+vMNUYG2CXWtElQU8z2
vf/QXlGhioZVthcSFP3V9G9ljVhg69r259J4foMB/aGGypkERJTJU7Y+n6jeWdqO4u6hArj2lC3U
zFgCv3Y1hj8CggaVdXbnSB3WX75xuwglkkVX/ktZO0sm7PDPNEtPHWGFWRjlKlxXTxK3EiOvxhYe
6v7Oi8P0w+cOrJ344jJBjhNN1sJ6Hk1SenXR4PP7RkfQWbIw2xNJftMkWjFZwBEPwjFDH0DYyy06
SlrWZ6CGdgyKhMtyEn7kFl4Eij1xGcs29R9gxBG+F6hIeEi1G/Js1iQz7d1R+oLJOEKtT550ThfF
3npUkUbJeoytSJ4B5sTUMcdrxorQFedFUwhjDz0lrabz4+h/eBEeBWvafoHQqiEH4xZZSli/ua25
IKNO4cV2lMICaO2D+KITw5KHkRCEu+r7V+YSerILQYv1rjTr9KE+Xxx6YrqxCd0Ce8Jof0uLeD5o
ee0Izt8NqiTgvNimhb1fI0EPj61xTTz3zfY2zkfUyQBCNgt/1KEco9bisc8zIaFscA9exIxKiBm7
yYl+vU2AqMdY80SH0WteziSzNRUqQae0cIrjTjn1j2Wc71THgaFQW/4n5V3XkzDLpvhj8nZIXQhJ
TsZ2H8TTaIFgRBRBjFefkHFxVdRSC5mJO9eeFvUsgs5OQraOKNtO/4Vf140aEWBBEuXoFo1nZi+w
uvXUWK71pZPWbjIXt9efBUdxpaMgYcGNWbj+cvP4kMJFxnJhY7DvHqCJD+74Rj5ydx15H2c6Nv6C
TcTDobAjKqK8vsQOTkE/x2pUdVyQKgzuKf9Q4HwHi+yiAF8ya2EAslNUCMEggyLZDPYj7auERQDU
DBX/Dk2N1qRFVZpyioZvFlMK+vUWowrO3hvIs5d2kFBUGdoTi0H390R3KGRlF4TQQETTdfF20UyP
AHmtdtq0zMkoC/5QgJi7B0RjCnS5X/wEeFZOsy/U3MpHH1ifmUdhlFyJogqi8Jb1sTYfMPWMlNW7
NBJcJCUKbdZzOwEzmBHDJdpRNdGi/Wm+v8saY+hGm9WW3bcN2vD81H7b7nKYcH4yn2QMgU2RB7rr
WSP9IeotmKSa5bznj2gb5H2z36shcsD6xTwiA648QD+SlNpTXcfuMyZNfA1yx9O6vl83NDU/FcKC
Oq7cExV5gHvwFYw++EmqQujN6m2w9RR+EY4QNylFRRfjPHdYUIuYnKWUj4Tm0tNULO1oUGIPCR4E
2nKnsYeIq9uII7rSV8oZb3Lah5VyMm/xmfnL+NYQd+vEY9JdCOHfenyHA6GvGWwEkIYtTpBMx2Jw
KWh2hMv+lHCfRBqsjhri8AYu0GM9sLGxpv2GtW5pI6SVI52jwfTTLbwJpDyQxQMGzimyzekVA3jd
hT+cl2LhQUF1sz055Cpp7ZikR6Cthyyc2rBXx2VbC/q3SMybreF9PLsKhF6XkWiqJsWI2bd1P+1+
e5gTSFTqWjxxaFc4uyRWeJ6PvY6rRnQ/hjB/fkWnnDMMcSP0DbQTqBM8xdn89VHLQ5mtt3FdtZzV
ES8ut9u0vkCkGN6PQtWB7iaearogM4anCVSk/L/EhauDcGVqhSRBE9RdeJYhdV7eGhYJPcNn+fss
RVARkS2XV/vlrg5yCLiIZZ43RvSY3/k6EAxRfV1GFDrW8Hb0w0zkYl/UKsyV9SWjySowZqENSQZf
Mu91BLTSY12ChFYZ4hyzopQrdpkk/YyxFUTfVXi3xS06sjEQr1cdKPb0tP2J429Acpj5ZCBwcZW4
DBSCkhMA3wwwem/j1MBpQzj12GLB7C/Vq2OhGtegkvzyRHZdmaY9e7dF50h83e01DAjELnyADT0k
de65Uhg6gD/YPHbMwj9T4o5EQGpDtUp/8IoTLGvGdEe5Z/+HljrE2UN4aK548RpcYSj9nYHJ7Dph
V0XaMS4i4bgtoz7FRdiWTviJd7zKICwUOEgR27kLILbOmE2xJlZS7UspilOwlnhEfB/BF6UUAskf
V/VI9unVJYUVNPjkFR+bnIICm93goi7xfVXOKwH6nPcnqdmr4TPRH7omK+sC/tz9Jzam+r7N66Qs
bXkTkNTIFMHxKttV9m1g3I0Cktu9PyubdnH7wD4YjcfPOvoJ0MkrLUtu73YU3kR83YZBMb+Q8K1v
tQY+Kpb/YudS5RryMzmfH4xABcr+L1fp5deXBDDmLu5SgTZdNzm/9MuVcmxOjB7YQK/KunM/SEfI
r1oUDi1aIrJ8/xqYrppbybZRjb5vYhLINdNbikQugWqxVM++HSZRePL/RuDcao08WVTEsWQ/+KlX
UZmyfOuoCdlG3T+2S4ec0OeZMGxKba7WDzG+/LoZrdlVQbK/jGYCU/HugZNnQJJEfpQ+2cgh9m3b
pql7UzKWyLSHxQg21qJT06eFSEG+hVgsRURfuAehrcVFrReZ1sSSg2ZYcyeGPxdueqgbUITrBoK2
nJwyd0e1eqduIMU94gAcQEDXnnyvg8h/gh2Jq3DSTP9lNg/nAAHfIKJJEjj0JCgQ8HQd4zpG9Jj/
zXZoE8Lod0LAkB257Hg66uZuUEiRveD7mM2hHF7pZ7cj4MfMydx6bp7PFzS5ehvDDfQU1971qau3
ioCWNX/kJMj02RYyCavCu/5Ndh23nAfNISd40Yzr2kbrUbvDrBxM8LcqlpSr65WpHrRXDCmQGHe+
PsUBcP/ODrU0QXSxwguT04LHXwiZIl2waeivEHAghvxkvi+zhWSDO+kqF0wb7qQpLKBH8IMG56Wq
iRf2fi2wY2zu6TKzeCCjZcHo+PaPg7lWy7b9yUBWqxbbN60irYvn5uNQ4lLnwqyn/zjh57jSf/5k
k670YWZpgk2rTKck1dy7CAix3/5GpSIjta0R5b1ojNK8uCcieubWunLtmBnSQwmY0hHlipyM906r
RxxuA5EvBUMHH1eGt3PM3m0tfLovv+Ugj0ScjvVLVvsI2IRG3i6I9jnQ25byE+hnPLKxE30f3fpT
lqihi4tOrBpomwb11CU5iVc3oi9vlW6q2vA8SXfHOWDLCoMcAlHMlDGHWKBcZzsak37rwWYIsFcm
RJE5JZnNa2eXAxPkr2b0/3pRRfYQefbIZSSsehaQ+sexBExsI+x9oqUQ6u225dW3wsGKfF+BFiWI
jN53VhU3MwCLLegqzywSRBqrKm7YCPQBRCehWOfkJ1Ze2kfsshBFSyYvbvy41vvZ2MCQltdLgTvc
R1IN2vxpSWB4IpKhfEXaYE0KmlONVjRKAxy2Nuy5Tvjh/bw0D9SNiyzJvcTGq9AW03cF9teHRi6c
e8Id9jCe23u3EdnpvzEuNYr0v6D3jBPBAYw+nLLL+EpeN6Yb2/MiKO4HaD9wiBDH3Tr26auw4Jhz
uIrm32kg90uZPnuzA0fQcSQpaU7s48Wq844+4pjrhtI/YAxOUUk71DVzYlA2UMp4DlJWQD7hRGnf
Y264e3xlUeBnh2EKtzrbmI2pGgKtu0y+yU0NXBzK4ukKU8jQf7QLGyPEoTF0QkV70L4eka6jR2rt
rf9JYOlTseiBtRfR3i1PmBut62Z4W8KPVchXZweLl70fGvdachnkUUl0wUJjRnwsls3JuuxiFL1/
qkMTXZ6GsKLowTY4C3h7f8soCVbIj1+vfxKEdeu00FjkJN1cdlCSWQmy/SjY+yXKh+r0dhLgOlxO
+4UpGpi4OmqpG1brHL9dZ3MRGuKzSMysZ6x2jS3BlxPVVjf6jCCH7AVSBlnI4/H8aNQrl9awsgkW
Ec6y3dBbnkgmsq/KYcs2IaOoVhs0Mn5YcSqnVNn0SLDSdAshVtGsnVh+OMZelOlYc4HKLAYHtgt9
wZ7IlUyJ4sF/3CMTENALul8hnvCefoT74F9inE90+CQxNePeHmkKSXceqjCtgaDP4oB3FBQFopZW
//ztUEG7TOXUjfO2yyXZNfVOaSuZCrTBzg3fP8GDqxkJQd/g/t1QjbmVuBXlRQAjksmMQW5DUxlY
yaqzz3Zh/kjMlDWm192AEQ85RoGpgbIsB4Qe6q1icn6srrMoPAOFho3o/d/WZbnZuWLZm7hJm7ZP
kOWYlYYTA2LVKvl/TrkJmWTRFbI0YOnwAeJW8H7GiLhF4JdRRAhwc2/dnThIh03hO0nZuXU5c5Kt
3zz29QRHaZMd8xTEsw6PmkKgqACTNns2NcmCjWNVJQ6E7bTFCEBvRPbJKM2i+FV7TwefPO/OBMpO
APtx98CmLidud1Hd9NXV84t+mW0qPJWo1Z6Xk6AYJg5+xqp9qAfItWsnsj9RtEhLfXcSjgqjVtOm
H6ESPMRcJc0s07CzhsATnKkULXCY+zsUTx+H3lX4nNqCkiLR2RZoJnusaqXPDfKNkUXT8Ra/xawA
xLZP6ip70VwubpsrfdoxNHZCmhQbHk0RtM5RA70xmrFAThXJw9PiGPgaSJtegAL3Xy+DUu75qHuA
V9aKwnkiHXq5DrHewzfapZs27CCR58kmP7HsJgLP5mRmpw74fy8cZ0+nksm6NhLWNJowq+BMpAxq
yYYGfeM7dBrixC9teY0jTNwDrPVINNyZocFzqyfmakjXO7jOnlnsiIgieyGDieW3YQX7LtO9FxoN
LozdVAtDC3Dc2GaSydETdR+5ZmTJnqrm69SPCvQnooj4mxvA2LcCKx58PewRY9/6obm4O/GNLFwF
sqBt+ScqAZGfki0TMPTuf7y5PsJpQ3snQtCETJdNokEfyOpES89kZVnmB8cE/tU+qTheJ1i8K3XX
hekaBjYuuzhzPKwMbzDWTpctiAi6JlkSigIDMsjyN6lVrVatT/J8TI0e6L7lq5f7a/6HbqDCt2ii
Ey+B/O/cwDhMqPbWFjwb1h9REU64gt0FOpIa1SVbeowg0axhaau0CMJ27UjEoLfRmXcJPRUDNMIX
wwgO8/3mRH+cgkfAg2LDKMIfLj3/MHouH45grxX882BHesAKm98xxcC9msUl7Vvut8g56nn8l56N
AEcUxHNg8IpGZP62jAXC+QXQlgLuFozkmA1GFA66FUkgatNFswEKpdrfAU1pcPhtqiYqv9YyTfps
MK18d/fLC+yeIV7/DL/H8w/5+sGoFMlsm4si1McyCyejH/8cSDRBQhcnTQw+HR2opyeJFi4z6lSD
5oDRhuUCbywMBra1W8XxQI0A3Wgmar/3Nx70AgRNIpMTvWht9Fdv2g3XYO8X/8laEvSqRcp/9CtC
b8aK2yjVPsGkd3mQ3WMg22yXbx1wmDtcK4uJtxEq5Gz5cfnu2FjqZxKJeCRRDiNU9B3zE7gsU7Mz
Y0GDja8vVG4Fzu4zEiewTlyD6zAI71IuUGxjjZL9Fecj6g2yLmdebz4b85CsZ8FpMrLDoZOrKG6y
jL6QQR8G46C1hzRGbBL+Jx3/C35mnPhX7lG46lEgoGa0OPszojkSP8Ts+gtPS7csnsosH0BsHAAs
Sx3t6nnXVEjUbQRCt98KxeOALS1IU/7cSNoMkZ4jWQ3zvo4bZZmh/ccoabhHhwLQ1BZFuLSDwTYl
3c/x2onJCm2x/V9v5TGPZqz8XnglfCqxknp8i0CH9u9tPynX8XSb9kvWAcKoTwUl1g9mPnvV88vm
RQWD3noN+mk+2yfG3n4lbOEEbd/UquSBY3cAd8QeD/3lGrZU8PiigS25IXWr9kRVGdrdg6E5RoJI
UeGANLCEiOGieqcBfLk22dCwwzrp228yEaogrKYixyAPAPPbuHqBnrciMdvuj9G4m1rGJnLQV6FU
BXarEig3k0JFLZBX08HRFB8co8/QwrwdFUqxrB1mGN0GxVC36X/nOOFetk6LTm5ShlXz5v0vRASC
hecRLRI0ti41+YQWjhqflDUmhF+vr+X0yYdL/SL15yR2yMSxoK6SibBzKcIlKVgBDF7IVjRzdejx
m5XG0bHqnMWi0r8GVFRhdMG0ZswsLg3PnHxiDntljwjjhMbCjm95O9fKDvDfPPwOJOWVb+JXwbEC
B8Qw2ytCsVn7TujRfeIXZmsDgIyrl/+XJcSJVWtENb5ckFFomPTumbosF0zcKYwNn3m9wupdjWON
v3bRkmCrT1QPqXvwE1/THWkUR53HUoESMYyj7LxHCAQo9P/U0euTJkwOcw8yRTAyv/2+nFlwzn20
YoAadIf1JgKsWMkWH2eGleS81Z5bAA5qKTEwu0eunHodJ+dr4KK/yJgpJbht17kfAK7iBKQhl7Iz
WIBBGAd1J/9XT0tCDUM4yvNwtrb2yaKfrRyS/jXdI7ef3eJerWPye8yyV8ehtjH8l3GNi/ICucQY
6qdxqGOVn9KiBRe5Ki+wu7/uX6z966VIXigsmndbIh8wuof+qSbJy+EE3jn+s07JmfihlPKfWLB7
SCvaubWPFh7HZyxoJbRUKFFdBMOd5ZQNR8ELFiaSaC6v8u7A1CEf8a+6hoEX9uYTL+i9sUpTqK7F
sSFh4XBnadGeeme+spIwdsLgvBATCxpMMnFTROrH8l7msnPK65NIr6g1YZQyDRJJvQgIIL5IeIvF
qaJpmgIt0BzsoRDjk3iK0uYkMeZmrKtvgE2PIs2e+82CzDboFshkpwtfGXRao7ZAGJAFa30PU7cH
1SQWRIuPeoDN72hTAR6bwavttMZS7tWleDyQqrVomGJ805X4Xx4E8nXFctveskDSYyEHoiNvgtQE
NcnTIoIYR9rEn31nQPrQYNla8Dl2n6WHicTtu22oRqyS/u3rORjn7pGXVsitg8pHYQZnZDYmBk5w
axL0PlVlZi1ntKjtsdunIg+BeepBIeIK574wHxKrzpvffB1gkbbscRLAt4KI13R/edQqzT8hSfYO
3GbMW1NahuLlGzILrrv2mBsRG2U1FjY3k4MQLeg/5wbNoiEAD18/RPElteI0JxrJc+RBfXduVCXj
+zq3hiaYrzaQAy2I9y3x/vJcNsxiSzjJidjyMkG4wNuK0B7R7KSYq+2LVhUu8LD0pCI1Xv/9u4kp
3+8Vm+DlDVmpJFcyKfdBLJN6GP8spirDFrXH/U2Y7LnkIoWgHpsDMitrAtwp9r2sxNvjqtZZLal4
12wrqHCptIcC3efsrmEbkkX5rQ1VlZ761KPzGZUZqVNmAno9yM7Y90PNRzCMcoKrgfgiuLHCs7pS
Et+z+ljbQ7vcF/QIMhAR0Sn+LHzZmDafN5mrs0610GrDm76LuoJ/sol4h87sNv2uUA26Pt4Ay2ki
kZBhmYQUiyD76xUKioA93WyjF3Nw2hbCbZiUrHMe56pve15lrp/MhZk/tMR5hQE5v1XlzmiUb52X
VpuQRC1YyiLqpPhrtIXJAuveCmPOw2d1A+WU87IsFNH6gHpcBhKz3nGZyadnqhbLYOOr5KdIjNBN
T7ghCklkU441eH3LhMcIlEwIrZc+s8hU8uHJAnMnRBodQJ2tV9qiskq1D2EuKMpm1DQRFRmkTDJP
nse74XIZc+m7XLObConFa4ECzrxHP+uQuAs1gJEHupZnsqBP1MEY/hk9wAU4/5YqaNOIAKBP8JFR
OFcvNf1R/xe/L5iyFm+2bdvzGkTh4uKAXt833e2Jd0i2AXdOqwPSstBCl+A01C4SG7QlOqzw2jp7
R/3O/z+CyMeQP+z35zXGZ6j25yHYQiMFs1xBds02oUyZ+Wj3sZ0Iu1+GiKWl0z8LmJ8pczHvxiEs
xU5jivfk2tBhq7b/+Cl493I5fF7D2X9y1c69PeL5kP7q0jnO8jYj49EkOqCNxe+4fUAmyO36IVVy
1BOwRO3utDFurWnp6hFUzhRI30rDa1HvZA+lb8DVWc07aP0aQerZhGvLSkYFg5TlNkW2kAuDs8rX
cZbYzoDqqJHTCmI2O4i3b9H/8z8nE1dWrVPLa/UiS4PVYCCoAJFX1qxpcPXjfJHV0s5iutqjNVSj
Mf5v5h+K8k/v/fB1Lo5S+fBTSgX+kU5n7pvbwKcS7WYGupVLTjLL9oKJymk/8PON4Hj+u8ww8I9E
HXdy8CzM018iIXmSHk7Fw65eee4aOf3J8dvJFegcuwq2nkd5BZRC8TzyEPBDMeA+nxr7y0sLpT2I
AUy4zdUIPyiOQm9TLmOSMYS16Au3hg+VSU4Lbw2njx9ozdf0wFrHLCjb7rV/kC/HE3cBOoBfW3DV
884+4qDJLoZIpaWyp0ZXDmpnUt/xQJkjqIaerB/C0Jdv7YWLdmRiLQKIaDWYJuf541uJZ27R9hfH
tnXOo+hLdgctYFTfXqc3EIzi/EEdyIZJmmOo35KD2iXtvMJ4JG6VSQAR+zifvL9HFe5vXPeWfqe4
1uI59PUOb37XTLjOIce7e1fGMymmlkqmHr8/8PKktPaar1MHxHOnhSOzZ0UtaelmkfBidgDxT9QU
vLO9EAHVlMkN1BFB1f8CB6AWIavV2kgxGgugV92cq+y885bPec6ryaJv3IfZOLtqKHHDCduVjp2K
euhi4qpPp7oCcFc9luyqc8+SJx/cY4s3phkykL7++2MRh/1uckoeQc+5mIIcHhHfwMQjPYgJhZ0U
FSOw79sm398MPZ8qbmUTIxLg4vbzRLjEN3GSFqv76Ah1HRKpmULJaz2yXtxlUMexgo3a6NTwICfG
Ga4rVThOSqlcq8eAxSYxsttZpvv2/mboBz5lu5spsO4t0SJovICV3g94FKUlY2u1t1adWH5nOgba
+RMhQsy9gCZ+AXjn/x3d0VJqwfUtQyLAu7Bnl4Gstb5spX+NmZIo5Op4vEygoNfZhAs0+FyVe53P
uxgTcBQ60BaZrw5pVFl1wm8PniJzxSeUomu8HZgnpKU0/dLTMvGt7yJDcBJe6fyKmbBX9BXTMN2E
YJfRpbr1lfKDatlITtc7AFqyPcebe5WYAYY6zH8misAQdwvTmL2Lm8l1116xkJC7dQ20j+k8UQh8
7bGVBhZNLUOJu0dzXcYgVt2kYWHayHp5QpXseBKbDtGM5R9aACInYHB1vznk1KTUnT2irv7T/JVV
mwxzSELcUVhk1x+sYH7rB4aLpIWea+erOWPfrSP9bjzcbZb1FeAg4+0VFuG1/UwDAdFmFbOANRe1
lwkKlrX7tdBWFxX66H5PLWuS/G4Vx0kIAayMPEWdkSHpDdMsxvvfZTI/nwh76HOhKI0P5wsJV2nW
azmiGVk1qzRNqZeTgfNe2ol3Yig4P0ewJziNS5u/Uslvah70WcX09rRHdPJq3o89HLqMel/HCfhh
hDO3sbN8e17flIf/Bsb4U0WYVZtBWaFk4iPkDmSlh+CaTPS20axDe9lQWgKUl6n0zkPBokIGftWb
gonCpPv6wDjHgPTTENZWWKjK+vOKwx94pKYQfMkPeocytygkROWOJfxMD8Vxbt4mokuHAgfcBoGn
+kDex7q/4EV+kVoxHUFmYXjFGtcUMglj07SsnLuSdDDopqykr5sU0Ks4uSo6qlDQLPRoRfaz9hUU
8U0nLsmK02YQv2CvepNV4sj9i2avH2t7s1tebid38H2yyOh1V5dKJ9iTqfEYicYyzNZxEDTnwSqV
EYCgtTkVXhVsTsFKMXU6bQfE5ZjixtD2MCm5Prc50SULksLIh3wBh0r98R+Ye+DLEQcDLVOLfCOu
sUcLbkPgnIDSvs0sFUoUTiauLQPHv2vR/k222kJRtVqhsHLWfZHv8Nu3sprWPJbdxarPNgN5D46Y
ybFRVhZ4E/JnO8CBJ6JltMbIikqDt5b5sTvAJAhYZ3YFZKqnVFiKI5ryr0ksKfJt1oLWtUzwlQ4+
yjZxGUoxgfy5FDhjYeMyJy9zOubHEhZn7uh21Y+sfsOBjeFz0txp0TZqqLiYyaL3Mtd2EvKhT7+D
hyffktcxKD0BV4tZ4gi+2N8V9Ii/C6b1wjFJQz3qkcISIJEzZaS4SgQ/rh25fKkHBVFxlykVA/2u
EySrtCAi05/kGOpZK5bSBicafBYtOOgLO8ELF4iNC8JGwZeqJ/su3P1IOTPakGbiuIOuNcZJIquk
B+YuaxsB+iYejwkPi8mv7QwYfOG/B+wfeLLZM7BgQwWw7tUOdWNWp/ESE7x348NOy0GPY4sL0xhO
K0HqaC5iQpksZndsHNET8ZoJQW1QZhxeKtKCJIEoQIoJMgdw9yyMbF4fNN2C3/n5bIZUFKkcDegM
/MooTj6Idd6vzCCKOx9bDia2egS5vXUPX+dICYvdhSeEBNV1ssJmav03hJBFmvmWOrc0Wzuazgrb
oxsqsahDHJh5aa5rMfHF3uRZvfLli0SLxh7PGxaxFucHeim6dqUWRDs2hLLVPY92OzTYtSK8yhIZ
gGInRF6gysREaAZMSCMAog4YpZSTxaR4eaqpQMidY4LL5QxOQaoZKPaPD8cg3cg37FDID8StUllA
HPFbJQAL/uHWyNvlqcoav3ZPceyhGLfxpKMlmMrKUjE29k8BPZ/ju7UWTB/YcWLuM2k/XV0lY2Rk
3VmJNVy7WayOQ05ue1ORG2NAyLxRZx0YFDaXYR54smdiGxVe4kynQQb6lDKg9iX90zlQr/UxjZaj
uk1bUOF00uZwwfLYZn0S30tDXrYaIEBPKTZzSq8kIs2lvf6MC/VJG/mCQ/kRJRRtd+mCbGBoZrbQ
jF/UcLWt+V8OSncMTAV2fOIAZcaiCMht9Ts/ThqRmiN+laFwwyROPuV3ZGUzv1BV4FEXi3cpPg9A
mlHjU/XsKl2yIF6k6NPlrYnMMjyOi1RfhDI+usnBJGY2Yqmnd+WiJMaQqx6gAJEOtq2bCV1tAwkb
yAMHcGLtdSHPbefUT+PBIMDu+6DEtsWaY+i1N96Cd63bCMJUgaqFianWZT/xgb5FjJrI5T//zhJ2
v0UTOUhAzI/7QbHmTZqPgeOhNimNXlQfTgyUFZAeeS/oDZ7kPQThyM5QdqzPboQxOhJ8j+BXwDtz
IDJeKP4nbqNJi3IGNae3nhyf0uaWZYgokLZ89KewIIkMSP4Xclm8dg8WVKkah21k5zBs0JMKBdZG
Ttd1NOVJ5ZEv7DVycqGihYjgEl3e0KhqC64Sfl8YxZfWfqXk0lDUpIJ5gy8FryhA45O/ojWy1ff0
dzWwXrf3Jo5aRGtTXv5WOfxqFtV6mw4NxtfL6t/Nx3HZYYOLaDThXEYiN3HHDX5yh2weams81PY8
m+ZzMDYa7wEZ35EtvoQri/02//plUE52p7tqGDMDcwLHudnER0Uh4MwnAN3EtLgPn9IRs0lkbGyb
n7yOcaG8yR9cFVFosdBoXQ6vtwuUCI6E0I4OD+L8ObcvT5szByK1XGurJy33FROkyM1rUF6oamc/
c/cuqh+ly4ZfS1F/O6LYYbKXTgtMgo9laJto7fwjgc0bGrDVI2IEghqo8P+q4P9bObbeEhWOe/Ge
ry09NVlyc0rkltCREEr2s6aXE6FCw+fIc6d06vnjsXX7sSdnogxsUXT7AtExpuFMg3WYx0FVb27r
M6q5l4aq/m0ZpJI2JLG5I0bm5NNopup44qlfWdMJSSpNP5a+IHip4UPzks/qoK3hFKzH6kBcpjG9
bbd8BXUU5qmFJ8Dl+Sz8LPfsQrcV4KZCIpNsbDZTi2RMsbY0R2HOT66PsfkuHG0CMq6Nqr4jau5D
uDw/EySoIfgSQksVszREpngxYzCLjN/oQ4ywtTjLZ3hR3sK8LpfEZFRMY+04NnSicZPES3U/sl22
YcQ3//mWeMzr8TonkJK6uCsiMlBtanU9YzWmAQaS/bUOOAqQUPZxXD0B/1XXOpBqDm1qUwBMa+VX
SRr6rSggQeB1jWfe9e1YBeYO9wm/NObY3qHbWCI9oGQzShutJkpCJETwKAFlwHy9gxcLN4dKIbF+
9CWPohfdNhr+3hsLQzE0pKazq3c4xK17peoHGaXHWfgaMIy+okVwAqG+Atf08H+m2naFfro+2o71
0aP1ea32zWslxaF7oCLr5zLtSmNKMzdedxjso9zPBLQkVV1fjidtVSl6b3YiaBaX7YQdjKSrMi0d
rVkxlRX48qWsbUshm8R0ZtEyyBN21oB5p4G38MpeYEiGVYobflWcs9Sc4FGQjWG4EaffLi4hBtD1
ITEGFEjdhdc3AzgWk6zNKaF0UIZ86gwjvR1Nmg1Oodm94X64JTcEnJFWZiuMsbrCh0Y50emrViEC
oEXwnfQHk1WNRe8VFp86f6iurfDK+SFPSJ0eX+S4VVGXaThvBTtYnSQG1tms4D1Gwb/cMFXxi+ys
gboS87fp8dgy630tzHghZc7/YzKJ8LkXLAo8dzAH+m1d10H/tJFMeJ4K9ZQU909KEIbQYSl+TCgv
0nTWqcIZWgGKAApbBjoW+xy5N4Wt+dR34kd+CZ7ysZ3E0/8ewKxywJpD7KaVuU+LMQ+99KPyZ/gW
XNQU+f8sHCHzb2FVXiAfSoV4gQtkqYf5RGDmvji21mfYQ9l2dyIjYwuYN75tsiBpA24RsxRC3L5D
ly5qQ55WtgoFqJ+oCVWGjp88j8XxF6IGU4cMplhjK2isUzEPtkBR+BhjlvpNhc5Tv4W5qVVkoZJj
rIQL8dbhE1zAHxvOiooElzWtgX2ucL8jQH6alA8O6tEYqgQY7sLtcjL/HkkIzXm4m6qe4bZL01pU
tqWQy+46VzFzUObPqB4etmemSYHt+CgRwdSHU2S3YKwjOUkqNpDkMsWjG9CaBOWOC6VsmrE7iGhL
1kvv2V6YbhD1BdUMv/dWbsdlyM8X2IHIHt7kBClM/Chdo4iplI9WyZAmZgIkcXs87QcmBvxEiGNS
BWoJS0k8yT3Ewk/AMrIRouDppLaVhRbd++6J8A6D9o6mPcwQYvF9zFPyC5H2k4oq0tFdbz2BKd7O
h54syJrn6NCbZPngc93Ll5hsfzywP/bFQ2BsZe1166px3RAk/AXXLPKlF61YkTNf+aKyY0AAKNEg
IowHS9IdmG/mYWWJg7Cvjh/SxxX3fkXfOdqFBXXKpoCyVzKh9IKkesYUmKOnsZTCejawhx4CPBO7
+XOMnhWechNkHdkJSonrAIInksz6x9eCQ8jXUSZs0s0l4Hgc0k1xARFJpfL+rNNxloEd5Egs2j8d
PDPARDhTJkq3iGEOKlUl/w4NOchoQrc3mxNN5CQvYXkM//lhHtjmfrBI3iGcZJpyP6XPvTkWCkl2
8WZ5WqZhhomE6wg70f2pX82rs6d1R0LZj7U2cjudU7GZ5Kn91lwp06sOswCWRY5THQAx7Iwny1tl
a5hfd+rlTpdAPZaki7dh31DbilYKd0QcsHxDRmsI309D57OVnwRO+OSYHimI3mzaTWRFM4HDLak1
P+3vuvMeUl0oUZ26l8syJCElZDPZbg0yzfer19ZuQ5DqD5NrLPPZW054bmGiSD5dvSzxnm8Hj1KU
YXLSjUnBkLP5Qg0tB4PfvGkDx+LYFfI9lYZbWlQPmLCxi69w/EIUHyRFUXaan/Cdj1oscDDUy9eg
iRVvyLhqPdhZYBSi0IIV3/zE3sGgF05UvE6uqdahzAACzaK83J15Az0sUt8Idd1XtlxyEfP0LzKn
O6Jc2OVniYNWsmQZaU8pTm0xVY2csHcArCDztPD8BKEmmM0+gpvutnLx8iQO8badQCyl4dDlZCY1
E8vLWdJ+h1x1sRYF8vTFYcfWkeFN6Ud9eFN70yAGlonTOGLwtK7OWmg18OS85CLgNlT2nGFcZkvb
9UyqTb2guRG0/noMbjRrTYerGgMR1xIjRxzIol6cf1BY+AM1IRhKTnYJxgDaxrdEcCWpskwLvEU/
Bf9yveaSV+oHITKI31j5OaLagjXKic57YXcrKqkxr5bgnbmz2ZZfFOw90Yw8chTQtoooEJNsyVCW
TfNiTjrhlWTopGtABsAES+jthubtQtO/CNjYYg4zwTTyzgqO+aiwgRe5/3B1VB5gmNi6PWt3iYPe
5NzE9eobiveNNi6lVg8YQUO6S2+K9rYIGzy0+/okCEm7u/iV+xpQ2ynBNC76jlBoHJrXWY9zuTMn
0wxiAJLlssch3aAAy/Qw1aimCV06z9C7kdYFh/mF67GWaeTuruA5oowIOo78D6YvQomDUsAmAxWg
caZjpbdH02oqLJc1ujP7u6Ewk8DLJqnHYepEQLUIULZ3QXUxTzcU3R5EYI6LNKrryHSmGJ3hr35o
FAannG/Co6E+F3R58w+RcRTyikmV+UH8MxqS6IMaRjslm11NGEy0IgORTfmepWiZhNc9DTHnP5+f
CF7dj6SSF+PhydfE9x1Fuj9EpzPq4EnJy0WurKteNRvQFUrhe72oFOQotNC5eKr9SUEAdLdPxPhp
cgUg38CFoo3Wp940aBGcVoz8D9sokgf/RPDLheOZqW50+fnBEV/8/Dt1PGbx/xeWCgPtHjMyIT4s
F6lUMwCjqfb8YUEdceamHAPR5Go55SbInaUFYUElaSwjsvyPCX9ud41WSbmFf8HTHM60eOH3Gwd4
rapcYDRYnQUv9qN2y+vxfuWgBCDmlGq701AhjXzuIROm8YGvdA2lixcc5hDsjEHHQr3cQ+a4k58O
ZFTpdYW4zWYH7GCPB4ahWwTHr7PGYS785TSOBCoUxnDZhW06kbjgRWAWTerRoWTBDGf//QmrAywJ
5Al8LwrCaPNUt4btmhMPms6bFRhUkMbc+jCzd5o/ghP+dls92speKVPiwkG7u5KXCUu0gKdQifys
Zoc4BA4tclDnzXbNoaOtAP1n9RfuWrHgbcO3G3UpI7boB82XdMdob8PUbSwsnzpBtXO5TQAGUWd4
1FA/4/XEzsSkLlEEfnotCAtwKMHz7C6V/vMd3xnyCqwOpyoSE/e5YjlRcsQhq02ifYPRniSbk0Si
H5FUFiEP5y4n0yYtNKBKjGt4Fbk9cDUvrFYzz4Hln++BIy8Wst/HJFxv0oS1g00k0ZVxtsrFZXZa
5guzEYtEx7MngN2EocxJg8h9HFPUwfraObnT5/KGbf+1BVnFJfxpDrmmgkBvMxWbsshrm6NuT1qT
KIUfKeZZuIz8gsA7b2SqLjzbAFhL56l2nLCuoQZ7UxC+V6D/nAm/iiKLybK/NwNMKBsjlKqQS+SC
VXVx4/EOeS0SuUmVv3ZsGUXX7olKeNIAU74vqgwieExAyvrNNQoLM01PfVMc7w3QRwrHToLXh+FQ
IRiS1nLCXY8pBZ6rNNG5iYrOlGzdgDFokV+t+Ai3BtiwnWtx/iymj1hjoqyN2i5PHLIzNtw3Y+Oh
LgJMTy+GqlBYYE7L+dj+h9h2j87UnrtX6zzD9lAqffrNh83qxPBPTBZDmhaw2Jw28HuXz50PYafG
5xU4hYlCWfhl1LLUEWw7zVB/2n6KKbZ14cyQ5JqAN7eUxlBTN9o3op3rEMux29F4B241hMmg2iaW
6ya4s+T/hcrudueZNGBCKN+DnO+hyA+3SwnhDBx24kImwIOyX1BOfOwH+RHYN65UooUWoCIIrOnG
BA5TJ2q79ItPMSIccV6TAvX82VIgCCuB2vNxtfj4JWRyZnF+EtTGlzhXQwc5kIFLB9j08XEWQbwJ
nzB/fa7HNmhvk+I9sZabiIhMcgE3vdPpE/76UPKw04d00Q3ZqHln0St5BXipfQOE8Cd6uabqTrTf
+IdrkLeodlL4SOC1v/stBRGdbJw/ByqAm9iks7JUIDBj87zDFOfMoN6P+MbQ4kf7QVZmSbVtGR6w
ks8jqglLETlXtj3/w2Grfb6c6qGeejdqu4Y1S8JIQjmNjMSneK5qGLzwvK3q5b5O0ZYbhsvmEJhM
gn7kicyToAdfj/k9q6aiLucUIwUF42KssC/bahHdIoliJ9M0ovpmBDK9uFBGp2GipcvVI92pHQPH
oXJDBPJbA/tA/o1qIWbkhUWXO9bhW59KAP87grvX8anrpGP8gWk05BbflHwBxPf0ddmDOPn699V/
aHWr6cGM9HSO6TcayTFSsMbrEjo/STB3HzsSjr7wGa+d5ycLmFK9OsyJpG4acz+U1M+/YCU7fn1e
oNysiiCMaFrFuARnabqCvFcgo593c9sT8Vl44nZtVZImWzxldTjhEhYJpnNBI/uXGgSXwtgW6VLI
QZ/GaM+2SAKS5uB1W22mOogcVwAOWyXoSLmJcS96QjjdXFqA0zLeozyu8tpK3qxjOXneflDsy8tY
QQdYKP9LIUCenCw+IY+2L00a5YXfq0R8Tuv8ov3WZcRKq7OEXvOly54yxacA+/ncpSOKQn5In/Be
Nv3F1mB78CMbDmP88Zgzvi6bl8bpGDSruIfdhKo4rHD+JhbdWbYN4IgZ7PkcnDpdQQ83RItTfr6+
zpp7uRsTXdVY8rKXEvTQ+iLY1pJgEmeFC5hzOkY0h8jsCCCd01+Lcuy62GeANuoyJrc6NYlQ9vs9
S6Tu7TbdcRIjRaUSbhesEAxrYa8oSf7sPgxbjDf5w92xgRxAwORuTkAXkidZfFkzYpfE+SVXnWnk
Ti3/HsCcK/jfLEwRd2NwtJn8PsdDOWNEs0hajEGf/3EMf5JrteIhO49G42qRuCubc6+CpuE5nhDJ
4y+JSinEI4VUGstnui+WsGIEKanGoxJuA1+Uh6rKEKNznT5U7lGzSlemDeZpid7OYm7+3QjbzAS8
dZFBE0lHrJpAvRIW3799ZdilY5npD7azx6MyYYeINPmFazBHdmQDY7/qpo/KoGCqC8X1Hbwm6z/C
aZLWlFavePVXTwyqqqsgSq4R8thdyOh9CcXna0Vet47+BjoOnLCSRPxKzRwdEHnAP64Ni1jtFe86
vKOksKn8amwFsXX24+mgywZYOAtqr6Lr4bSMFaM+ENmsW085NpN1efN9pUt9efAUFZFdoGHsZXc9
zfxNAGOnVHJfqENs5FeHFL4jrnmDe+0K1j9x1/E6yBotM3E0naYMB3StE9lpvaTQHTk4Mk4YdiIp
70wuWGEEn3hq1ny72oJNdxYJ3+HEGO2LEf96mr/6VuRvnU6e/aBChJ27/7pNAFCxfq92CHaMEs7t
813oLW70zJolTuF4FMVLqGURO+2ROkItVKKEEbPlJ3c88hoiyaOOCtN2p9hejt5cV8kGBA2DGDb6
8nDbJdjvw9YeEgXSAzAcA+sEBUvZ+w4AgO/egTgsypdSBcrd64H0f9U37a/NgVQew8XAJ57aV6sb
29ClhfZwDkGSYj0I2PlT36rsC1LnrfzR748LgWR1tWRXCoTXXQqDMbYP2weiy5tSDom9pZE5Smjm
h8vnXM05ekoPrIxf4SwZS1ON8IWk5bQacnQOYYstG3bCZfrPqn7QG3eDIKnxnnFu29C5dChYYRG5
pZnmCDxuSEdqMuTZxntwOL5cAYJ1dpR5JLQJui3EkjhZ1h302m5kjFr/ZlZfnM5Accezxg6A/XvP
hMD5FVtO5UrMYHI3sr9wZhIlM47FFk+RIdD2a35BhVm/MkFrrV1AIfs0yZSZ2D4NW/KbiG5Mt29k
huryP5iU7/2pfoG5Kr2wk+ItE9P/W9/iup3bKydEc2iSqMqJroXh4Co82eShZ5ioGrabnj0P/bVf
67uWNvVMLmDzVOs6M6ivwjPWVB2tvdb/l/YbCtURwQJXDoeJBLnG6o96r+JpnQGndoPjav6zfoPo
Tb+4jdoO3qYi+ZDl2N5p4dLDQEgZGmRs4W3yO7CB2mOFEZfaytGGUKm7iQynWodTnzPFHIbFYJyj
qdRKn6HNrTb1b8nhM5Y+D1Llqa1yQvo9inAZPpL22UexFffsYF4WxjfDz2D0njjmMw1K4Bx3OtZY
urPqZSsngRPUPhTcKZOEKTSsGHsKGmAWM3/mFPG2HElTuTsvQP6vALXO9Mw84HFf7wHogJcSg0d7
yoidAeOYTlCDM4m9ZXIrMF5pJHAqY/LGojlh3FyLy8EbCIteyrJOO3BGZNcn7FdT4E6CsSfqx2jC
/6wiTchyEuF5GT476P6RHwPv5jgQEeQeKQFIVeLpnV7C/reBYiKc+drbB0PfJaK7w6GOlY9I1fBo
p9AmtIIQRaix3oVfA+l4aBJ+nfVZQlDrK+1Ny6e+kUpX4Wl9gtkI3MqRTmNd2h6Y8yD0cqYb6oFE
t9ExsES3m/izhfWbz0nPBl7rS45NHarr62vr9crVx64rI6PLjhG9ApDHq/b/7Yq9NCCuGWV13H8K
UxFaiHggr3+7aj3T5wIFNUhS8oM7zzK0gc0MLhoS1l96wRJe8bLgDTEn2xu6vbZ8eQJD6Q5xeqtn
TMJZseFlBnQfyuaPLivSZvowIQGCXmTIoar0k4HEumEhGN/vvv92HgW2vooBxp2A7ScZbwUDLtQX
KLe48j/mXtiwBPDKTQ8WUvjUlbiaG4ajpKcPr211U3gpp7GYP+cqCU+kjfE+tnnAdpu8IVkEyYsp
ZrrNVnMAG1v9d4fvMeCtiiaWzswC3q47XkyvxgsTIKDUd1Wk5iFO1/ycfftO7XNzTVKxl4raXdik
yb5G9Dm3dQxpzaeSf/X4fIX1U6CUKQHRJib+/K3Sr2R/whbLad5B2Kqvn8gmxw/XZgWDFAsX9ZmB
b8eIpUIjwP4jb5deT4YyoOdeCtjNsqGZbsw1tMoSzwLRQaedg/C4bYfg3CiOr82NEyXO/1aaJNMO
SFxTkxcgWZ7pEHjoInSCndSzli8HOdNXJKffQSIqYTas7/FEE+IH/sQgHM9i4ZnJZwmXHV+UYPFV
9r3Sdbmg3eNE7Vn6fOZr/IS2gyuIQVUAfaTLljeUEKfm/CSy8QoWdrfM37Jy6d3fMwNau3QWaxjA
kCESW4Q1ejdVOClzUhHFGWNM5AJhEXj3vKe43c9GVjxhofPOHyojS2uj0ld5ZKfVkoX4W4hJwluG
4U85luYMS9+p8cdS5FLmLJB4QB6Z3Xj99mOCrPnu3b12VAy9r8ruAjEoKQOEv+NmGivcJ4TpEOQf
MzFUkJdxBfHQ99gK1eeZ0TJ4vtttCyBI1KgIxrlsLzUdx13THoi/gv7QtALvSYxcrGDiVt0NjP+P
jWpdyhghWPjkw41QYv94AmyQk+PrZg98lR19LDkl4hC05XUY4+ooJsnCpswL9Po371vm6lvD7mp/
JWMy+AhvFw3j7zm9aHkW9o8DmKHTVR+eZ1Vn+DrIMNMF7iK4qR4p8oozg7K8goI2C5jch5siMOQf
DzyBIiZCgGZWuPaO3oHlsdG5uzdxAB31AXwgpHVCCfnKPkM04Ny7AbiGd+YtKZ6bg8k7KThBLuyJ
xO1DCeAASJe2yFz9EWQ6GGUvKOn4ApOUP1LNj9N9ssfujeaQJm9mPBgsLb0ohMRiOsBhfL13MfTc
IsakeGmCm7W6sx7lVMFDAZ+ry5TNVU0wF/4d3FB5rWrOap5pPcgJJrh/C+3xyOcjR1XzTqAiZNcC
3ED8hNtqLa6oZEuzXssZYDjhS4PH72l8TOM6wuynrIM43Oz6DzpwbkKXRUru77n1yuVYe2ZdCUdb
5WY6sqW8bCb1IUkuHljabCehtotnog54m/CSjBwHq54JlMLPFEEq5D+wgl9jEyE+PSyC4x3zcaQA
2dpsGaW47rBHV3aMxl7/jBogOdtyfXkquiu6GtR4y1Riyn/vXe4BOJiwEIBSb+3Yt+HbaJ3Z9STs
/Zizb6sGfyEdawKVGUB6PJ9MnAiIgy/g/GrEUW0RhBermn2uB8ryEK6YRKH6kqCmvFpxNx+dhizH
d3zyk0coc/Tm2k4JgYYicTB7F/AbfsyTQ7RdDp8iJHIkSTx3fsgdIsP8oys/zMM2RPAQMlxa96uR
8/HvCQLChe78ARBFfPkK3Y74tTaU3M7spojYr52rVIOHCf3rHDdQUPOP8p0xvX850RwFF3QoebQ7
yIWsp6/qsjqrnzN8rNLAGAGlGHoMS1GDNkktPnFHBqifYN3UcN7cwrHV13u/yVNuB06wKwlY/fbE
0i2RCTyHsZuCHo5eCWnZ/3P6Ufi+EcJLYZ3FDbgjQW3ZLh/oQmVrkshQTLRTMKP9rOROXhrQ8N80
0acKQaOiNWsFQt5BnWnDx01DQghQ3RV8+VHJOYO7RprQLk912BrcPblTTFCj0qHwt1hZPerxMNOK
4lKFXybsDZZblsh00PVSx+G8c7iQqGNdR+rTN5HyVNtsha+ps8RvEqzLezj64rkcZr9Kee0SXRvj
8o5cCdNRUbhBpZyM/i9TV66SttteR2IHbLuOHsxq4I3JxIYldjE3ltMLttakvuHKczwBTGs+/eGK
5/WPGFT0BQUODqSEw4tsKpXZtdr1Z2tFYv2uW4x+HwCXKoX6L9OHbr/gWyYTY6sN1obZOXcB6V85
k29ZispD8FeZDkdpXJh9QAESxCIdB9rwsmW6T//+XBChj6liv9WAc0X4X0XmpTYhpEAeobvfVe1d
aXyKckDYzC/C12i19ZjC6fCElcP85r4vwnODHbFO6U+ursffVQPwdiTWWDDt9KBfStD3lHAEq5Zj
lY6SaSmpwRAJNZH6H+QrSHn8axf07ovMTR00AwZBMs7jGdBAPlXAUKgPGB4SawwwDzS7pmC2Ok9f
NP2duHxBeH87k3BQo2rjIL0Ilu9WeW7MaQ7/wwhnkXkgIzk7LWauuIqhNnzrFFQmjQdpbfQDVH0N
wTXmBopaXbMiXAN9mEVNL77CROX8aCQUZ1Iei+YGKvsUJ7lVjz8YjR/m9y6BU2drvbSEoAkN0T6E
oPj6jWaF7WY/WX89hJeYYd5NjyoQt+iEZYwLjGz0WUpbz9bAFlMEWjHxEqDz74Fz19Hc80hXHwHi
ziluZoCYsCn4gSmn9TyQs2SAVJo5uDlVCoDgAVIy5+swMJRUzUJNd7T4VyzM3fDCIqWxrnH4Kt78
LTdfcr/chj0GwXCwdJyx4xFtWm9+201s+UmYI1m2ZBhs9U4U3l9Xv9J3oREr1cpH5lV14/BJIYV0
EhOflc71nDoQ2sBz+ni05r0aSKygN1QTkAgWMPIWvjQKl30Lwq9A0O5gt6Cr5NwQ+yCHuYGgK0wV
VUZETUitGyrwA8Nkhv2Y/EXcKn+t+CkC1Ny6GAv7xhYrerg5TieX8NyAmz0CWmvsvCoXWk3al1ak
xd0wsTaKSIIT6KmeBECq3nldDKy88O/Mr/2nHcgEqB9PU0DOH0IqiCsaU9hgflEgrY5GyxXhlIfJ
EpczzMABjS67PnKbPBWF8PVUMUXbwVqmOhyWeQd4fjZ1uSCb0Ng2VHJj01C/wB5lfT807o3BYWSy
Dz/2udUBvMK4bvgHXOgYKryYAj4LYVk47aNiRrzYXsKykJLcN+XGw2kXBYHnrWfR3lnPy2fOa1Tr
bkr2PrxMk1dsTyQBHOEgpK60aVVllB8iIUufddle7DEj7Hxm/fJAZxorcEm8qtGgUhPJZvGFJNsW
PpySNR94sSds5WVkJ28/yKrhvu1bxsC1OlaHJlt3xSYCPl/fpiO6zBK/DlSlLICHrA/uTt4V0Grw
waVjKdxqWwwKW8wNNWFd12w/vwmClCyE+huvWxisBEgtb8kV1UbPIICu9KKoQqGVkgL7oT7H8Fr4
ulMCv5qj0EwxiQ1jzNfyD75mAwpKyNGeGN2Weyyz7nhWfNsH8BC1eSqsCa98TsxIq8IosKGuJNWd
NdYb06WtABQ6BKU9rdN5MRv90G6Ln2UnMNENgRdsTg/dRWIhhUslNF1kATSBehuBH4iPkiXVqGna
/g0/ViInmFd1AFXbECRI3QhXLWBVqsY79WxfbiNK7IdRi0F5OM90sKiB73IbDN5hCr9O4o/CkkkU
fOszMPz4BY9X9/anx6d7+tk820Ijhi0iZkGCvlZ7z1vGRfOvFWKZ/YPjZqgUof1rQsJRQnwDc/bj
zvKxMh4Chhi2gLAR9XCruaSzRv1stlL/msH3M9thdsUoNdx5srK9w9JQVAR6T3mCg25eGKio/ZDb
LJCVT0oIpd74lX+y4chQVaRsd+MsMAWHOAdwnUz5rSetLssfHXSrV0V80FjBLRnfv+3C6f0M/NmB
5QWa1esRapHI5d9O8NNuvPSl7pltaWcYVUlYV727xLaBk/p6/K7Es9WsfyGqqY56RNh60AB2JDZr
2vfHRo8i6KtEv1G+BvO3Mdh5G1fVEMdK+3p71/eMQriFRRlzxhLKG5vz+bFRRrC3t7UyjCjwrEJz
nHoPi7aLk3UfJIj6LwTxmyaKNUV8mhj1+mZ04kfbxmflcXnmxC2LTY7uQSoAHz/CSEinHeMUUScf
coYTXS9Ifzb9joljeZvEvD2AYhoCe8ByVUVJYe12Qwu8FQB47qpZUimUI+HepCLspzwO0uDYrZK2
0fnZtmQU2yvq+eRlQZQKMSKH0m6xERuPvxdibxRnZoziFV+8d+ZaUO/oWpAME7v3CI2NDvnIFB0e
hJREVOa7HCAjuhsi2hfM2Sm2x3OU1F1/Hm0YBCWSCdEUjPpRjBLYoItyZc76EcbdEuauSS7dVlPM
DYgGqo5fPt/fiEcdzHZSHuWS+mPROTHxTb68xHAraIV5iGdnceST/PELqbG7qy7rA/J4quX/upSr
YTQTp+qNl2VjoGpF0NMroZW7dUeip4ngL8R6GhY26peDIqB8avDRC7X/fQpkMR1uH1TodlkpgF8m
Z8KHEdEj1C0cHH39vx49UGJNR4jvUUZo9EuEWyhwq+caUs9YfFsJubB3Cz3UIW1i33s5dfG+N695
/JcRJPDwilfmo4fJkE9zxd6aP2T5l3vzRaSvtG236nyPDBzmgNotNAsWyqxBFXXlnGYzq2VlEIbB
pLdWXd+rKXM5esrRSHzHCjR/Lh6VycvZVkEhVNdCr8J56U5hTyywSsdYqWHH52Otx6OQp0R6uTC7
7uyNd+D0Kugkd0J6bIrn/7YGm3NWuc8LyFgGdQbq49zJPoAzpJdL55EXi0rmKSHl23RSPbaTXuUm
6bKAw/EEs5BS8q3KuQpb+/c3E/DlS+DIg0RrY5I9XiRJdDAtO4ykJ2r4twbIqLWPVTWBIV4238pf
4JNUu679gJDHVFmFqfYrxqI+GgPBGsRBcQ0SfFWjXt2Qy2Ku8rW6UYEwPUWS+iCllpLT6i3He9Ry
q9R2GduFnSGknp/Q3kOa//u47wyXUiJHIm2N3mYQukRsOtk6JgoKyeEyxcn2PzUdzF/Iiu6PS9Vq
Zk92pQZDQr0WdC6vMJ8VJZHQqvBtEAXnayGmhUBtMuj/UOunPSeMHNd7Gf0eewPdljumqfoprXPF
BHmcLrf5kVgAkMf+DbO0tSCn+M1v+xWVB44jUlMb3EWUbIp6bdo8IzWcHHW3RCWmpDbNxSNmSNG4
BUWVHV2rvoOAhilXkguRH/0m7j2jfqzXrwd3b8cCBFNsFXifs3LdgS02xzrerz+kVZQEgioXkRrh
DMNH3ERMSCnOqp1BeiX6rPoLt8nmPbeMpocy5SEGZ3zDRkaViw8r8hYPWryzz+zfs6LQXo/aXA3j
cyk6wilTlgkODXYyLEpZ7VSMFZshkeUWmdoh6A4mju6JqxAjURB/7uDRYOOEa/iygTg4yfSEBmn1
mxbdRxkMH0Y7rmGI+2BCrPMfw5mwlVYORJ2W1XVKuNT45kADzmrbfBb8/zdrRqgP5RgnSQHFm3yF
uRRLkKTcTCitm7uFP8lSJEFYuVgMyoJgOtQDCvO9iGlmNT8YqK6UUj/sTaisIz3DiymLUmm4rvwE
SIc3WQaRMFXTbs4ZW86MWKkAnYLD3z1TwoDC8ySpfs1S5StPQtCG7DxLnvTfaMb4Zjmvx8P0H0S+
KtFbFlp1EiGf29M6hgRjRKG+jCh4+8iOLREiGNfgloKaVJuCyZvc+0QONO/MK9KNJ+jHbBQ52nSW
nqwSvkFFRTWvba9jvi4t50V92uyd84uxSkLhfiRpTdfoj8t8q1CyaeiGvMjdUFJVxF1VF0tLrlMd
u8szCK3xiNhJ3xRSn4GelqPlsHMxVnY99Zd1cfc/0WfbfbETmBt/K6vmx77FNroR6E0GT0GQkz4y
Ym1L3EijeLDndUxrF9Cnc8r62tEFNrTCalTPt9szPu0XTmc4PxVW05Ewz9DtL1PP3d6GwnleESH2
SYScRAT7v52UquaCVfcgPKMbxnfMFqYxouEw8oAvUb1ZZNRQzrqTBNW9vqMdu555lb71JiS2nWcV
cFBoezy1fzBoHOlK2BtfqV9jmTfOrIY/NGk3y79ALZSExG0Fm1QLacinc2Ow+VT+kIdFbG4fiVjq
4VBdJa2Iq85uwOLJcg5Em4tdjXqil7w1UU2TDueokQgb7AQ2Srgvlo0FV1aJVoe+k29X8ykrD9Gt
I0KHP7i9PQ9ihQMF5wkcUcy0ElcDZ2Umyx7sVT4koz2lkCoHdzRJ1WOEI6N4Gsj9PlGjMKUNHcvd
KcCm+ZVCtV6iRoYR+eYVuXnzq56qCqYYvoxDajUK0hf/v16LSePzh7V5deO8kGq0e0lY2lGDNJHF
en2WSKz/C/EW8h6XdchDb3/jtEn2oNsuN7QEZu4oyxs5LQvHsCGg/35eGvvbW/TKeJopu+h60N0U
kkx9t86XVrvp3aB4R0iVXNgqC9E6aQw7zPax4/y8f9Z3f9QFURUTEbAQLeRIlYy0iyLnMPKsoYvZ
4pDVtWrzltibiTbvNEoGsvAFhuvfHXnyzHbGjAXwlXKK93SUgsopjhsJdAr8YFunKkIxBYoogUO1
EMuVE6MoTmd4JGeIeiWdtucoMMG8kKi3o8KyCT4HeoKw2niojD91MZagReapigu//KV15QGCAeL5
mqte16VelNSe8im+8S6pBeIqMDfdzJV3mmtIuAKH4d4um21oY4tdzA3MwvQ0K7DO2hhc1ZrqvqoY
6q/cJmHIpOHSFaCfcTNfZNaYTOXJOujHQW8342AAEUbLzIlc5C478Zuk75eVKzT5XJNBqol/Abmm
if/ZT1N7ufWExlZ2sD1/lSZ1128ugWC8d6zCOx74p6gVGT3YLPeakkbfAY+mvVmWHziDMeKof3sW
fUZWgs5uu9OQTRTG6w4W0dmPIaxWOSNdx3UxiSUO2SRcPP1j8aeNk7ei/qcHGCM0jmof6BLngoE2
gTmz3Mie8r5ZSoarwXBbVw5Sj7JhWUmeXtR9mFxTMFVnQPdHSccrycMK6lk1nXQM2oybkidBbYPp
IIZYT0coaGSDesUMBjxzaJm2CigBFAY2POiuzk3pAWeBsQASdB/Es3zuH9Qj3kzvehLtMvgCsE1F
ewVqzT1eMlIz6E8YUzGdYzBi60+9zkWDPtTDQYaRZnkOTB0rGYVoSYPgOAMZN/1YmTYyErO0q3hI
5r+EREtupzXL60S6OQPImnUsDugXrZXd6W2KLQNlBOVpmJ5Cwv+HRPqVMq4Ua3FE92jmRB+IjOtD
byWoCEpIo/AwtuYCysJUQUtCTdGzbYMq2U3PlwiLVTkS30uErYBnbBMyvxgUXNUh2+ezKtThFn9E
PD/7RnylEoJ7+YWSH8nyGKJDpditOZPviWcPrIQFRNJ4o+Ok7bNlG46ZAB0AwFqnnd31OvsdeMz3
3s0N+usiBE637paCIZKrmQlUe8SVMsyfgoi9SM66Gx5BTuoYy5ZJXxtGZidhM1dtSMVYugslb2ZV
8R1I/HHn0KHi70s0RZcDYgvd3738SdPRZSadNjxbj/N1nrY94utbgDuzqPeJOyGWhpz9SV/xphGE
jF4gukswddQQ2AGiovsygxfZtwHZ2u8YZh1mPbWxnuLNw/mJ+AcUxL005vr/xtUFhXneY3648T6X
nI5eqpLa7LMhOOhluRBSPdZJtOYUCDQSU3guqYAqTjeuwBIyN/S5nKbn+//OCCJP0B+nTCUjZ1rC
DpzvC/KkMhT/LsFgXN16Q0Fgqu6Unl8QtxHExr6D+QzdaFPWsBYlC3oDA1CqT8L+fquNW/Iix/cM
Xo/+cBrX5v4zt1AkbRPogkjL5kbWDaUZlDultYQE1WzaVbW+QFun0XvOITtMQYBX8VC2epf9kjm4
DGbdMb0igOw5lezT3pUUVXjSWkEnHuBQzULyC+21nZ0NVtgerzri9wPPpvNO/Qk/mRRUp8fhWe+b
hnGzhfE3zuNRP0LGpHcpJ817UY4XnHnkVRNMkqaF5vExG2nq5FPMeIvGYcu55ZBH1u0xcHnTdUYt
/s4Xy6Qj4/4p47tbZhVrcGgoTlK3dkJi9JYhZw1qq30CXqRrZHgJM+Cq4fHEVxBrqBBD0OIAuWhg
j3heAbufy6uQV23YFNIRvEVaEnJaMSa72fQF+1w3RyeacTwocKBdUkf/rUFZIp3Krwy0nWl36CLa
pSv/Il4w/CFMgOBsZnSKvk9gn+uZfRCsJZ0qO9e7ZkyFYXKckXy3bF5t8CH2xzxo0GZ+0dXxW3c3
rsLOzpX9FCEImtlff7uqpZzsb/0JDmYd40TLBJVJF26NXiPIkpJuSAlsZX2QyarLpzfIJS1tdkWT
nN1JWmCPhu8Gr/YydE1q74md6HbAkZ4Yf/ttZy6G64Er7PYyFCtNhydtlQocWuq96POg8i4eI43a
/m26XNSgF5ipNdT++N6bq44GLtAxrXVw57Zl0u3YhLt3MCS3IKGkf6Wp1IGeI0ono2qPKPwe5pfR
YLlrxSQXGiqJrntPsVn72UBzKepgB29QjaVrjaB6siEeiyLhvi8igxFnBwe+QrsOKrhBI80kSh+2
F5N1fiQMvoJDO7VkIRV4iB9AF8VQBCkziTegxQy6nvMWS23IWAlg/5YTyNhAsuL3TEa/wDOHUGoU
lxizmvgAZmCFzS6WLmobsShZshNB0GNiSrgBl5hSBMhc8S6H9Dga1Q0/lSBZe8/Rc2Digi0+YGLC
p5BP9c5IkVX5KP94N7A60GntF/99iC4HX9an/xoBWYkdhhJVU8eKKNqnNNpY4UCxSwBEStPaQ0gh
T7kZscbSHGXRMJrtAgOrbM7Kh+5pFFxzK9oB1qBoVUDs5adylCMOWYhDFUXBxDEwZL7L9FlroxYt
Bo+Nsg66V8riWIKWGer0QQD6nKinn+wk+s4ji1dSPFNdJDlq9U0c399YahoS4kWccCK5IUfIYDaq
YcbCxhd+bQ61cF9EZrcKv+FrpDQBfDmWmtfURkiO6uMtsTWYzgeGCGJ5fRA+aaoWB2ut4jyVo03z
CsT6VuPo4GDBBISjT9XWf2UgKv0KvCQ9tTjGVhCLymtz1HhrZQKtj8268mq/4S959yNVBAZDN/zV
qPSCHC4qLKfHWIPGWx6HTcB2td41tb+pUVTilfdFDOdpHxXTuj3TFevTL8wH1QLCaFnGNOzsq0uV
bbCDaJn84eZq2UQ0mG6k/sYQYEkQVuhZ8V143FES2/PG2hI4qYkfmFg4xgOY4YfgLec/+/wnsdH4
7jERyGvymwO17gny1frWE9sos+dzKx+T7Lp4adXaoP8sQshm7ceQMF9IugAN6iTDYVE62yJ3aQtm
I6zkz/NFBDEcn9yrxbpdj2eq+lHvL5I0jftMiniPpULPg/wpCFozeuSfXrh82N43MAbOh86GAOJk
Iuh1srlB2hqMK26fBNc0ceyVXqliWVMH+zTzYRvbBMrEfMfZi89PRV+CMdOitJ6LX912mhwaU9RJ
QQ67+va9TExX6phbKVavyPzZio52y0mXJpP+Zx5LRBRWLsaOv2j41CiMbcCOYQWCtQL6K37xB0Qb
TPQY8wx3o39VL9w/7cJcq0e0m4j12NHxSAiQsk3DeBv3aRJ9/mm7sntw+qrX7IET/im+kC1D3nxA
7tUh1V+knzdAI+UoenueDySkZ13RYPnIaZ8+w9K215JGZ53iPVsmLgMIrPuSMsECk7KlxN6YPFnO
d2MOzRFPAH0ONJWNPUX0u43HQshXCelcRZWX26eijHcLyLXACPIjPiwqKONi4UyIIaFfXTfo/xtU
TTdx5/YkXSM4n4JQbuHHyXaMxP5BOdgT7THQ63EQADmTal3YCpl4hMp/x3n5RIR784uujKL/Wp9z
bDRtpEOpok7IBcMxnoJpvplw5wKYPXdEqZuVjI0CExVAvAihuyZ4Qdg94cPNaPru2XNdoKBUCesQ
Cypmbu54PyR4doTHjbh6w9KYTRiFS+zKQ7qCjecxKs+JyuyxVfD3MILeoY6+YAvbwrdGHcA8KNyQ
CLcULKRc700M9hI1y5yc47O7+iq+R3kmPx1k6PYSxG5N/Cwr5hLNYVh3GPEmK41iWThuyKOCNLk7
vBv+VmNqkbH8THTIJ8zAaRtRcoW5MxqN+ROcdiANghOHR/X3uCTWVJ8ZWCQhRTxvw18w5yzjtx6l
RtvWo0bzGlC8Up5HTLsmbTr5gyhMIMai6u20D7MZoh4XhuO+cm8XpWF8LtekEkY9TppRULI+XxwE
TTG1NdBxPeyHdRzJThH9tG11hxRJ5gIQwks2a4IkbzmdtSEOQIX2mSH/my4PGUIgWYhNwIQ7HeAa
jMyVJ2e6ZCzL7P6J9lwsPr6MGlhl2V56qJdQGIeH3+xwajM3MJdi6dQw4MvCrDIiErlqI4jY0iB2
8m3ckWEboxdtHlZkk5zFFAkbA+oSZpewzVGM3j9ccRHwdOWyxEtSa6aVr6zW+afOMatES6o+tZgW
lDPhlrNitOjfLwrrzCZEibPIKAkvoaFheAlUadiy/rQGm6DN24PXf/b5AEiZhYEoWoB5PYXM1or4
A5Hk62coVz8qtHGs27WGzxoxMqOp5KxHHrvosJUglf08nrQi7BJjOumlmnqYDkQ/mY+KJv0cydNQ
GI43fNkAE3QrLjR4J5lep7RJ72XWB1cKgm6MYMzSsSIGuBmJq9STdq5sUD6/NEdKqu+bJ1I+U7TK
5gvVn/B7sv5orznsUtH+NGwdjLCPeN/DMpyPaKQwfakRy44Q7fyMZw3LsyMGJmWpWHRxrxu3irMB
Cc5YFHR781G9wd2eVxlgF5F53WNbnnXzQHJor5rW2p5Y8LfcrTQlMsaMgI+60htHRy/CzC9DBn+l
aJSxFStY3Y2etvIDYpRILjlJPpXA8ow90ot0QVr5jHu9K5ojYkO9D5VhrMw+C488mgLIji/5KRly
jec3+4CMdiWgpQD9AyIR7K4OvygQX+nwBfJVpGuxJUjPTAae9Kp2vCDd0+O6auYcj/ClvwZRYE/V
GTmHiTD794japOH/fZRUCqCYUotmJLnk37srNnUGkSJNFRBkyTChr89NAWYxzdMYUKW5fLGhjtw+
Y0XhsXbZCFKOs0+f4g6Q3MTdtXrQLPSLt5mKTdOT8onZ5Q4xaUyRh6iRoDuMxaZ7ZZl69XFFx8sc
Vrl8tV8OX22mEycMZjmXnmVzbRsXvvtCQLT0A9Zv890alUVe4RVZs3cmRy7opW0Tm7FQR573Glo/
bzejvP1DiDF7+XFZ5Y3zcGX/tyNEX78RRHiSLE6UvbaVR1tAeHnMqMVHgyVAxwDOEO4GTuspOpFr
7ZYYmA4JWCBXoclzEMAQtHxj6hBUjID4IY5MC6PJM6w+zTg+avIF5QHHoHdEYJJoWodzmlbmwhYx
TppIPSukVRgVZfAV0dssBGlgDkpDhFEx5pwskJB9uwIl6/MTE/u0Hw+mKnrRGJG9YWOcFXTg5QSc
8KvUIOwrbs/U5fEP4OOjVq8O2o5UMKJc8BxgKoFjBcrKy2Iv7KbW+tZ9pu6aaBiEEqsnQEeCXnVO
q04W1Kv3B4j+t5zTKh/vwoQ+F5QR5VZ3a7QaQoOg7uZl1PD0Zuyh5fujfOEr8orWbF7Qtm9TUZaC
UkriFLHyHJLeKjaTE+4njVH9BuWt3wZkVYJldQDPcNvlhMHVqOnv4ByZuqn4CNpTYOl6ZNOfdb4H
bq8lr6HotaCaNmzc4/5KPh1sZT7A5xLEmQe6r/+17hvqXEGt2LOLgWB5AOfcR3NZ3aTIfSo/wp5K
vOTceKbiCwa2xre1jI1BZcBRBGbGYdMK7D+pnC+PWWSyicKTJlv5qMLeIve83giKMVEAGlQGXhvN
xu8NnEgiWLVIOkxLrQIZS8Bnm0WrhZoscp/BUyViRhp6lbYbhSeXQ4DQD019RuQ8TQeRUT465MXK
pf/USqQAFTiJgy4UohVKemHGYAJU9lZtBBpAidMkovOg5xCje5bouJj4rn5sm4/xU0xbtSQgzkh2
4hIZk77tDqScdWy+PfLnR6OCSZQM5MehghVGhqPksHhvEA1D8vOLoMJEMqb41lABF0OuYFvdqv8D
jhpKqSQ/vmH1WVWyvoFljOC1jajMhReRoWq37tXDZQJ6TzCXQch8n1fHLApbjHgAg1cGrE7zXZ5W
51gE18ikZXwoXKvcbAeZoB5TGY4P+k+qGP7ZoTvEyDLXuL/KR6ftwCVwwXmfpEO9MX/5FES6Nei+
ct3paVYyE23fn7CvJPql7qoHG0g8aGAWQKv6oBfiJ/OTH5db0+1dnEczWGlIfy7dJB7KPUS3DV0U
8JrZIEkRRhw6SN9SvsDE49H6PO6j3FFkhUkk18x1YFERWCxpjCBZMcZqbYk1fOamPceq+Eu/5I6T
jTtg6SuqTylgR0CSBxBh/XLarbl7F5p5dFmfzUaoN6Qj9rMl44wJik/+R/jmOa3aMeBcwRbANjfD
RvjuFPvl4q/zbjQNstrnX0yH4UTDq6N7XJIqdQHOHtq1xYxuMaR4f1i1ZObhC3Jk24b5zvPtV7De
TU/XhrH3fdHH7ZYYMokatiwxBZsakT9jGeDIpVezEXpHlaIjmkRWNK9B6j9+gflDomciPBX+eaYR
qyYbOesNmhFend0ygXQ+Fb58WXIwa5IipmvqZK0LEx9fnTES2dq1+yEBlXVIQ5zw8rCBUa4vuwaw
tQkFmzQyhY2MagWX0zP2vVrV4velVou/aJxhVPmF7eUiofq37pDeVwxF3HYQYFnFVP7PE1oK/M+f
k6IX95Q1PxQDSjPgmg0kRvIpyojUTATvDXcItnaGI86MaYLO/+3MV7e0dUGdspsJXFZthOElaDt/
FGUY7NEsQXv+VjZB60mSQANdOCvwc5JbPnqFw3qb66VOzLvLAdROfwzIks6aOvMP0E4Vrn/zyBA3
6U/BK3Id8ioe30eoQEbUUbungmkPgXSbDOHdCWDubRE47H6mgViu+nCS7chDFfZFnas1HzzDxrbx
/Jre7HVNaVT5MLnCmnOUEJfN/i2ZZWOz/gIVlM28A17NXgNsjPNr3I43YUb3Yd/gTcPxy23dLY+1
WkfN8qL19GH+oMabFzq3VyduHHcAvan7gfjyRB5fAbPr/68D9R/uczEhJXdoho65rVmRwVdB2ejV
c7CJOlVRVu4HrKrNCe/87L3QtnSm3y9InwruIHAtTxoS1KK6myZhXnhdUcCoBSyWpf4dkO7DbUOQ
vwrz3zwcIh/iAqgiBVNhrw7ZUMPjqHuRQflcine5HoMkvRPc5eVddH04g3H74TJHTPz0tE0ZD8Q0
ujmtwXVrQMK9xeNbYcRZMJ+0QZ+1+7rtMGONuEIZSp7E1BDJyJUgLxFGOK7knqQ6Ysc7rRI5ZrG8
1p1rjskun7ANmPMzUf+/MRJ6wZypdABwXhrpKU1A8T/gSdjbOrb9ZG5MDEdHL94o3TD/6ceEFpXj
sXc81Rzr0YO0NYIoctaypFN1xVLXqV3u4hRKZruV72UbnKEfFdZDp6hJMjqeJ6PTdgUXM7J214K/
4AMTENwxQM4dMfMP0TKk9rNxy4jAUSHifOjHtgcIosmmN2+39EJ0I54nymjIf8JgfYf/bXJVdN72
XmpkBDMB/M2esd5i42zbZhq7fiqcrSOni/QiHPmhmb+FyrbtA7EIOc+bdx3sjftw9JCbYHJqkFDM
giY6G1PwfRiVXVn5/RrOCi+Fqw7m+Bh+kUhEm4D3M6zUk7OV/0WWdgS8cj9IzGYPt8r6oYjJg9i5
NLQ8v75vs/rkC2bEPAZTrYccZWfa9MABYa4kv0RbmHe810OlM/Wk7M39q7z0fKnWFFezrgOlNBfa
NKyflBC6GD+64Y0vHAjiGnSq6jnuikUu4UQpcgPqRRMtkJyV4EKgTdq4exlz9ItCXmXMFRlSX2K2
pktt8odxGXnNaus8qAGxS0R5iBPy6mPyVHETgNzipZ9qAJS2/Khl2ljGBFLKF/wHSkv5uYLKk7kZ
ynpTobs3Ogc+rWjGR1SQhr3GWsRRXFYxJSknvbOitau6/iGTPugStqDNuXS+R8ECjBSOqjJ6GBpV
m2kYud2PQ7sYoGEFMNBR4wECVz0MozY/sbqRaDke+7MfBO35VIU2u6X4fM5qyiPH0w2GdSa+c0zm
Rspx94C9v53f6EBP4O47m5Fo2imnKl9T7oMvdTyfsHmzxXoZ0pV8KalOPlWWz+8rTvIs1hm0fsnh
7N6iRcdxaWvdQTB01/JFetBVt0tz5doaWxCzDXetQIVikaarE/ra8zXjuFRlhNDFrBy0GJpGz5/I
cvfc0u4+fmzAHrZpON8/dkV/9n5emnbjlnAFMpHSybG/6jaWHvbcYazi3nw1zn9wxyOYdnWuAZds
1AETKZR531IN2vo6oxhNprMBT5Z7yKdJWenOA3LmhGbcmaCTWj7cktnVWO++ENcjX8FDYkORNNqz
wnc8cpYpUpxjZ1JZrKdgrOKeRboeAqoGuvcULJO6G4+YiXSdGEwoQsyUhBVGxYBZQKnhIxojA/3v
A9gkP6jwAeDYpddDN1+ocjc2n/E2tcmXB5QaPPvDKgnCGEmGG1hZA3ID/4M6X7TQb5QcmvWlgV/3
pAm7qAkjjlAn6/yvOt+i4qj4Oc9O/HDykSbhixOEpnj68/pWHAqz3yGPoMKdugT76y9JeB+/EJun
vwBuwjkJY0Rw467aPZRZAndvGWqCFmqVNO+w+1NYbsgb27Q8j2H3WxCCWXTj/5pY9IvxJ0/9ULqA
JHcZo7mWygSxLVq/Cjh56bfhvjtabwnQ/oPbdoZuMlxWmZpcBZy9b750Rdd9vzbtHlyXcbVfrHvF
dmzyQIbXdHDSke1dlu2SMaZCt3mxPcCNlSZenoFSiXY8BjubqEd1WuFQXYYhmZT3dvVfoBU+aH3r
wY6tZnYfPfwOaq12N4n+6MBchVN7xTJok8cGqsm8YqPuNxegfgaty/juPZSU3g7A0zpa5KhvEuye
mzxAoLB2NuOFKrTsuM0hkGiPcwXgwRo8rpo1CGDNSr/aMISfpFJM0T2Ph9ErZtYjJTX3w9mhqvaK
D54ivB8q+cOT2WZKal5LWhKLjBgRmLVG9WjDJ4A4JtEKB8FgA8xNownoFm9bAruUL9V6bKcj3KaR
Pe0H1Qret/wfvF8vNWrB5HlT+glMHs8x6bZo7jFgjpwQ7szAhhJZ/6/2ETpx1bRX9zo+9+J6RlDL
LO9CRcmGzFyiH/Br9fcD94Cuk1knHUlaDZ+CKhV6dDTdAyTLCYSvkZuoJpp6TdgpIPbQRJbCnDzo
/Qbu5rXGiYUlPHo2th8hjesnWeL+uWQ4kQ0ccXlhBPQmxqqoHq4IqxBXsKG4Kd4fH6CNw679WNug
/nk92aFnXXTiw2MDu0hW8Mv/GO7Sft7ouAB9mYrKBcrrFGIDw0OCq0fa34l4eLYh8KZURMLyOU8H
pwWgDVtmcGbhTnp+n9d8YhNG2FR1SEy44Mdwf5L5Po9rfXXFWFXu5gR3XJOzRFAHT9LzY+ZulNoR
DnlvU/R5DE0abrquXke/e9chZjo2MlWEMs1wSoitvXiTSMuDWdfNQsWNaCVGZMsNhzlngrVauSa1
NNzUf3qJXv+7eeqFnMQOyLvgbLrMzMKz2fe7FsYNMgzm9n/7wlPJDeDPUyTeMOHoopxyHDdHOevY
0xnIA8enH2cIRw2sTBGawdLsySQO0qDT2TaXtK0/BCx9QdjnaFGxVcfM21ZlQCJ22cfG1bb/2NOX
KnSL99uiBejFChm95e4aRcDZ/p18RIEbvFJrcnMbKbcC7v5TiTOiOvbVQnLm6o9NmAgCSCF2biQP
+ErunDpbRTjLzzTQBRmNJv7XoR+xRqUHp5srJSUu29/zj6InJcEJKwLjz8Chyi+2wKDI8d45JL8x
vBNKISGjk22FGOUy5eQYdJY1Zci8XJ76vXFdCDoHZrr1qAFnByKqzRnjnsbEdrFL0zSOkiczr4Yt
UVUWO+eLt441Z9pwo0VY4CXziAcB3Tav250KktlgCBpuzY2dg77x9sV8pdJLIbqhyRqh0IdtHPVO
04jLEWdVVbrjMBhHH4kvi4yrkLG/C5HoJ7JscKWupDkAvunC9MS8su9WSOz4hLYJU8FamwjZn1iO
0IOBx0ewjue/76jdDSA6DFXZnwwDfhIobm53RM4jrKc4B3Oc89IvezVTaldbHEZjAdEU13+kgt2H
Xpe0+/VENLtkw8k1y0EyvnmaxdAzzlWKOyMIyCWidPaWHHOpngkbcOq7eddNflEBDe2ZJ0t/cLOD
U+ordfMdaCFC1bCrNq5cYhYkVw9+KS6UgCfVBeVrJ/D0JyS/eb3DbKEyoTk6RDkV3wN7ckHxtTxw
6fBzs1WaCfsb9l9VjQNsNMvYgR5sgZjX3m7olhQXdYWRgykSqYvIuSwgo6+NSh6CB/pECs3OiGb6
u46la03vN2f+7fVMP/7K7NYbGsBz/EyA3F2mR30bdv3pb0iRFn/LNvYP4pvQQyiFJiscTfo74OP7
pClVn+Rb+jaFkBBoCHzM/0Eo2b2yLbuTaLv1hbczSo3DTsCCJ/tS3cKsdEJaYNNK99NTE9xkGRIm
FCLJzT2BdGi1VCdDnmj7iAbQV570Uxb81YADcUKapz+fp+zNDbVWm5tBIAltolyUt0D2cBzCsf+J
emyTG8DMerYkXOnjkxCg5qcQWcxRQ/56qDSwYqTQVTD6gcWmrI15cp7ouTCQnOhPErau1MQsJd8M
s/oLKeScBO5VDHzvvgk/wSUlAwdaI4ewP4LA32v2rsBstwI36CSXrO/rMds0lAEO/nljKBW8reIU
BpEHhJeGKFBPeClnmdsZ67f+k00COANSBJXddD0zk8pqosoWKdc0YTl+Ch8jpB9orRb1CBSGeQEu
NzUmoBR4hNVNoZwKavVUs5d22may5leD1XH4aNqsVliWel7fMP9ycNWbhl35/FNCRz1YZ7I8jBR+
peS31ppGZT4RgL4MLH96uUMxJb5l1unFhB/uBfqaBmIkG4mpHLZ72beWwjUcWFL3TI2kbIPvjo5p
Helr3gf6bzulwwOx+MFJBVmNhTBlhOH7u4cKOjweZzK0VbQIaCQyQID6kDQul+g740mEZ+CL9MLY
/ckubNg5hR222Th+8dRDRh0aErPaCHfMTE3+8c0Vvd9j2ksHfjhYIl9ukNblO+iBqlShAqtuNWUc
8qU6Xj1BRI/PU7BtuWzXEUxbtOKIhkRcRWFzEVi95W2MMiBmFTCiPlNKq0jrr044arojKQXR6USg
9pmS6Bo0td+C6S3bNybn2qiVAiE2UMHgBYwjssREd219aWs7c1sSaMkr5Hr91wIgKjGPolLyDHFt
yD4K9tkbFzsGARbscSxvBrrSFti3TXu6VOwpgREbD4WxAFSkt+PbxXqovFnfEfxFEKmiHT9H7zV7
7a+hWj+Ht1pqDzoMHbFOouECsh56wOmBy3aO0qR2kp9520ql6nGyWkse/HaD19VwjmcOkMgR5xxv
rbTrRnA9kxnic0lDQ5IMLjs5N19uRlKh4wnkEEvS1VXQLr0egaHMyN7eLH4W2ddPApmVHQDq7nsB
WMH9ES5ih/2RGznkBg5ZKz2fQvB6cpS1CvKsgnBmGzdu41eQfR81+IfGtBB1ia3C4QmH8cnMPbzM
hu36jg8T3mKxB5r3EWU4/HZLEVTxIibDFp33mUEmdcWoEJdSuBmnXfZgbzXNA37oMO1XQuS2sxUU
/LXpKFGvBLxiIJXQIRiP9s0cicS2W+jJLp/ffL6khvCD6lnn+J1BaIgi1wBP5CiBoT2DROwaS6u5
IbXqLNtxL++gtD0c8uypfUSl1UGTstcPepL4lESx/Bm35Ype7aR0KDdQt2XX7xIvLbLFAAhFdWm/
c+zno57c3fgrGzc/6HEhOBVNgOJLcFp0Oucj6lFNQawD3g/LwWlF3/OBrfL2SBwv7AGrfg1PjEgN
MufxViiDIOE42Mg7cPKwGiwRJfrH8UHbO0dHjWcuCXIhVZDFskmXHoRqmsMNev//7Z1zWkK7llDz
y+4pJUsuwewFyeCtjMx3Oug3es6mSj4SM7XPNmYmjpzWU6xK4oq9L0N7nj16yi9fBGIQ+7vgMTdr
qJkmNtRbFXOCcJ4oJmYM2DI58wUBn9de17bzUNOXEv4zZiP1r/jCMLkEQlS5PQABaKBg9LBclBh0
2NvqALdd5uiIa6kKEQGY7MmfrVNYbMNg8fTzsFOpYEGThlhu08YGRaRdgsmvtU3JzUCq57p1xkus
0XeL1SOsPKjUixNLqC3VjCaClagZ8a0JRa2CT9sHsNAYRPZsk313isxXP2yKeed/xltzvjSqRm8t
ZVm5zjVLkpxOGOY5VvtSZsoQJI1FBmlLxgodoLX17/LYQOdUjwb7Rn0S9qa3hN7nKzSjciT9hId1
xNswcP2tHB3AGfmo5CW6Wx9t78HJ1WMjhSXIbAlLb93wQAdVxAG/2r8W3pw20n/CLCzUUj0ZGoqp
EcnCXvHeS4xNsnlTQPoDJjaSIbF3S2IXEGnzTRxxOxImyA54PMdm8H9SZSMsC3D8ixjRyrMe6XyY
QabIW//c/eM4mJbxDnd2LTc2PyU+lUAxtTftwuev5q7wBqYs6u3aVqIrg0p/D9vAYj7Z0D4EYXxB
TkE1jZbILR/J0+ZVRMeWLa8JWquiOiFuuUc0Kz8PL06NbSTZzemmeiqDQGtA57RjXszaadkmuxD/
8daGKJ8n8sN5ymfpTz/oFBvh3U19cS6euNNtqp6VXxFPJnY6LgR+xIjBItexFQvCc+7F/c55WAgA
TgHNVpulzXYKnBh7AN78nAWWBCyKG2DnuaL4QQ3hw0bSeBSbvldO5lhSiId/loSblcNHJHZS6vNG
RRRceknJLAfsw6h/og5amyzRbx2tYgj837LCFmXca6pLf3pn6CRleAVoz7HXb1CJCSxh966ZIkE1
bOPoDdncduNSp8iz/UVynTu/810L1n4WZcxG9eg7dmG3d3uvZZtfGjVaMJla4tk/dGSuReCu7RGT
yT2kfxqJrH6bZzcGnOlQDbycqqygbPx/NA9CZyzgEidyq2lTniZ+RB+fHytyurz5gm9Bjw5Xsr06
W8k/xWdrFlCNOD48/bIeJIEpO/QSiT2glGBFd89LeD22NKR81GHmjhrxZncKjTkf5VX49qhDaHVS
LGV9XSLjFH/PBsXJtn9+L5gAXVJS4gJ+OLjCV3uRHMveTBFgaQ+wjv+Sk9kHxmRIiEo8BheFXKnV
uUOdmQ/huJEBqDf56MJJ4EBFa5zz13QWBy3uxBPr3inqGTqvUsfdWRDz3stU1w8DRwQ2yUv3lniW
L8gu77TaU2bZfz/aKHcbPhivXzWvJgwbpsByUvWDKESFd2Ph82Lo1JlCF5uct6iuYGDZ9ct3zy/q
bRGXVUNhlU55YyW0EudiJOh5YPGag4ZK2IIIxTkAbtxK6GBgY5no3tjVr0Wvr4BVm8TGzPJEA1nw
DXXk5Vm9gKxl9QH0kGrfhUgSUz4hHS3bcZ9xFTp1RQTCiqgGFPW9Xy5tyIkYy/MSbb4s2YF8kjMX
j1+R5PYc2qGFr5yjzOewLrlclmGLU07L43vz2Xy248AUyegMGAKIUyANO4igUhaqM6uIhnk4U17Q
l7sHtpAXKVMr+QRl25BSAEAHHdXUht7WoBYot3Ah0iqVn5RjkCtpwu/9oSp4pD0cTNFcgkN4Bn52
kzVLrPMGx/DgyAXv/iHO4+rnzREh0kHcVtOe2F9b2drh3JjQv2dusMSoE/u7sWo10WxSq87VkR5S
E4rpnQ93UJb0o9+9gRElKEs300PMbrMth8r5XDFcMJtWCh04QWkg3rffmrmIG2YOVUf+omOcG1YS
XPFAU517O/G7Jvwu3rZh77pS7XuaRLyiT5rj5rzjZlBXiuZE2Xxi3SsAfpMDoHNutpw4EaLtO8Mz
e6dlIwP40PbVQnQa/LAsz/VN5k2W/zbzXOy2rJgdxB6kn8ik62HZtpS0QxGFwfpSLEDwkByyLOC9
IqtKsdwd/uqLnrBn6s9Wy6BK0/HqAM53BgSKHyERBRYz3ZDPA6bLVycJltmS4zwAV3uguSmYKyw2
xnQCTChDVnbhFkg1MIUrnivh40VJJDWuro1pOYAuXGHNWEFnQu++OeW7QH0pIYScvutotju5rA0E
h6WXcNX66iJrLaG2Zp7fiX03E5y6mqvhjJklN1a2Jwl2AnfVcjaKRLGN7p+HzSV5APKTxWuzNeGS
AQTCLkGODD/9ndeFPnD418n0AW+qxTb+F7t+ouPIBJEQtTyRVGLsOWQdqZBB0BG2fHDz87Y0bd58
Anyy2oJBwwHi8/S87ZlzCg8MWKYN7t9XA7TAh4InQORax35Q2XpcJfnjOVXZXSF612r522Hegfvl
DgN3G+xLvTGMieBBPVvBna60Q2BssUOcGdv02VTLii2ph3iTviDbHg/nD9knDX5clSIwDifOk2vq
h/9ndJ3I78+MeABIiUBnI2meE5qwYAlk59khREoPS6NVQKhspwyUrbUK0vtIAwMS1m+iWyxKLQw7
L+MMB0iTV2m4L5EY+ZFUwRLdUFRq7ENHOImnHz8zmUvaKETwPCjVjVwbG6xoE/MhgdRFaWVPxQBX
aR9Z19uwCXO60Y1W/K0tHtLWleQSwhya7P4OXfnaZB/xt2SFSIY1pc5wZ/HNmp5Fy33KHl3f0uQS
KceR1dVyOrWoyG5UPsq3DbjCqBneSPP6mGneHSUzR6+Vv0k96l2+fQc4zET+5gDskCF4wViTJY40
yM+AV9WuGQW6G+ecKN2ntAVmoN2kvwNeYJbbpWg1HR2uZeNNk01HwyyUoNUuvnMPrEb0Oqlk8FGf
K07Jz4FLR3rZmzt3vbm6chz4yV1AX+UyM1NiCmUi2ifIqUdKlSVEKLHeaTy4zxSSOKcsCLXaa5/u
Wq6ZhnOGf7O2xEah/2HCam31I6A4i2H8i8e7jtL+R5UsKw8LvIoAZxD97ZCGJHFlE8Tk7hUCi54s
LWVKZr0Zb+51c3qNqajqZgMb6pimApo+UtVJ5rmln6WdDKAq8lDVxsuYLS6Ytwo74NvWlkenIK0Z
dW36UwbatOw81yllXjSzGjcJk8kqtvWETV6qV3RUn6+zqaJ96bXLU8TPDibaTVAyVPSvqYWWZ4dk
kwnYU4Zzv94kFgqBcf8H8cp92Nv0Aq5QznPzIqhIeMBI/leyBhCmaSX/w/aSmXQ3ItEV0MCkF2ut
YMmFN70cMhTtzoxZoAWbW4fRmHpMREKNCImA1w8Qzj0sfWwkLlPgrS+ipYhhph0Jz+GJ5decILhj
AlITli8bns3mYtoSmG/utRlzV/wZ5mcd01A05r95tHOob1KMzEia/sMdgjr5PRrca/peCluBcnRd
ONQD+NLc+SUTsiasZFcRGKbPhg4rL7pQN0U+yiMccqJDhwCTTXtQBx1GJ+J6BDHgfQs37Y056TXz
2k8t1lodVz4P2J5C1+xafNGElaTo1ZSk058c9lIPkj7YwoZdeSiaV2qoJScJ0vpr+GNzQMDNDCMA
+GYSYpRbCo3s8qmE86xqa113+rVlvDZ1N/ZIcz+/xbkOlUJ3z17t9WgiImgzEglXLudN/f6NsRc6
c8QwW3Nz6d7TLrwbMNq/sgwo+OcyTHwRE7bhD1YUNyzKHtWHh5aYgTSdq2amW0p/hJgSp37hOdyo
ZC5nI8QHaTOayjJQfLjJrxeXlGFFw2fk4/0eXzsLJLpErdgBhmmk8FB2SPgcJR0I7V2f5MJyjmWR
x6MfYpfwo9so6hzvqf1lhEFiuk8aoHiB/E8HfkR7hn6gTW420h2rA1bXzlVqQ1CF+4j8Nm39d/BX
32X77ponR8/B1CnB+vnGEAyKUJe/WFH+UaY8Nzedal/LSK2/Z/S0JuAORhgCi/gM3Ltb+xW7yRgP
4j3bbSAjAFhB869xEKsr+onvPuphYnC5i4TalbcXnSLkJYaNx8GM6JowjgBkrAPL7fqEgDTZzDpo
SzCwoLLdiyHOJ3l1oS12BKY+S/2kfSbax6x3OKDpJzVt7qiU/qavS8z1QJ0s5K2v0cFntfB2N0yk
NwBY28vzrw8oup+PaDd0XcC7UuNAyeaNXD+6kWyc6PyeiqF/lN6vXs2vPp/ZESJyFtD0IM/NsaRh
inmPWksTP7LzsZnfhfqS/4X5vKL+YS/kgW4YFupkWuH3zwREJZKFzCg2TRIe0P5nJ1lX3qnWgF2C
acbeTKdLib6JNf1aOB+zeQRnugsS+O9E5gzcRga4ZcM/XQHZcmkrGf5v3tsKmCF6NkHhNjH+PjoO
VoVvqxAHo15KHNXZhicDd0liohphnLmyAI7UZue9S3ustNGhydMcNdQnDQV9ahEY1wPtpik5BbPN
g/UM/nKZN+x/06lp5Kih6XVwchqF4MGKKtaux1LUu9oIV1ii1DldsdQ3x3g/10+YELkFuA8tw5vh
R4GTMIaJgO/5u105KYOkHatvYpRrNi6sq9Co+OiyJx3Ty9LA2TrseMIdTxK08fmoHxSPydwpgVbb
ZRNGK/CtmIO2q1JpdBOr72XErikAH5rtzWbghyAw7sPdYkOfOJYH34m3wlGvuSwMS0E1WmknOk/Q
IVHb/4oU3rYnUI5nFYgblUqA1bDHtnHRRhpMQ402JgMgoZWKS8sAoA2MyI29L6GueHiPQCzCBpOZ
xTlGgq6O6/CdPHkAsEBMUgW1dW+/tzZcLRR5C4lT48Z56l88ZwrXDPUCYZbhw73hz5HyU7GrfI70
UqGwD/XXk9h4O3OTTKhy+O+dwM1zHTjfCQC/yQGSJ4o8/bBBFdxGrkqwD5qs158zUmkQMJNxi13y
GXzZB9oR6plqB4wRIXGk3LF6gDe/ffawkF15GDy7RZTzGa6meriGxI0gON+sQ6adZhi/HoC9iAT5
az3PrgQyFF4dCl+qpbdftBp4KrdqF5pkmAjQDu9l60o5eHfXR50gRIKt5SoHnZlAJurB7/eUl1aJ
bCtPzASfma0pAsj0JS3QbMKl5BTQej2GZn/CQ6Ge5niflfiP1O8XeQh3f6PzD5+0rjgJTShiRQE5
bOYlV/rJN7DhlioISVMVoCt2iBqvjIdpsnSWe+MvGfITYcljmjQzKdQyoEN/Js/fxHZ9+CQmot6s
ElFzyOAnSVslq5N5vnynlGZ20VfKDfAOuxolKmovQvcJtudhRVbh7wFAcpycNELB10sHjQ7+267R
f4Jz3WOLP5zwrKbJrFoAyMPq716NWuCY7H1IDQQc8tpojEwhVsvBgOWrCyfJpIQvewg2uCz/vlwZ
VGMsif8ElL4mEzfNr5fmNMSqmnu66sQITFleP2cZtzIn+WMOnLAICOha5XEtU/dlgzGOwiyBl3f+
AIKRyVlkDlmP74vLsLlKYAKrz5C50nOriebin+6Pc2vIoYu59vjcF2BHrwjtQCgD/c12eB0rK5IK
z1L5rqdxsF7t2+OgJaRLnwW6FzuWFrMyIQWjqm9XzEiEoBWys6fwoqoqPWfH3ue+yOHVfvMscGdB
+MijEvwhDwkxKB4p1ZkVEuGYhvIg9D2EhV+c5wCIuEvHEi6PvnnAcMfu1aPEfg3ZP4MXAgm3iZAa
9mMifOmr0rUD8h1dHxanXhVvQrW3m+LmzB30rXejnb1ZZkRAc7BiB8Pfl3h51dJkJbWwNehkmFRR
h59uSyewwN1Bq5horG30LPqhA3JNi9paRkNm+aVIHKiZfLO5zJv/Rkbt4J425BuxKLKdlFmvU777
qtkoc5A8VWB3ZAUjHNP3P3ObhzW3o7tcE24Girc4j2mO6dKn55pnyeYODnN2bBHFUCXG9/eE04M/
exUGTcDy3hcYWy12hpAi2z5ZsrkCtpJXx21UrT052TN+/AH9SRRvpKwARYmH7BbKrx1pRzDF1KiF
Kf8nlfTOfzpMrCK7Cd7cUbC/ysr4No8VHRuE6rcNHc0LzpKdZNutD+VrcRwGJQn4QpY+vIZ/8JBX
wKNRNAmgfl7/bYaXWv4zg2FoI2xXa1XX6RvMctP3No3ZNrWyNeCj2Ta5qWz1T8OUBERjmSQWURGT
SjBHNWFo8Yv6esfGY4E4Bt3Z726aJhSYO4V7zlFuItuV51Kc0hDojKClUzQ4xtxnul58WCn8P8TD
3oR83rrKroealQ0AxZbDy1FI3Je2hmnRgVIx6gHYQipfmEdBXgte9+F6JclYPkhEgObMnLdS0pZ9
J2v2dMO51Iq0AptdN2A4Nf78up8cJHmVYEIqc5Pd/QiFrYyPv59cLDH8UrfExWc1mBijDpLDAE9q
I76bWT6qXWOuzOAVUZiPJ9BNk+LYTnllWXLTjX9nWuPqhwk9uu0HsolC9QwFrs+Qc+uRWqPql0Vt
FWAG4GJzhl3nrR1B7ZuFdm9ozFgNkhy/oRWDtfIKwK4Nv5xGp5Z8HkGyDHc/iXCFT9o0N0MQFvEE
yhErBCwUBCYD6G2rhchLu1uKSqfZZCsu6N6lX5XTyoahwgAqRLJxmNowTq07T/WLeDAnpZ6+4Xjg
gs51OJkL5DNHafZxG/TKdGC3wF7/W37s83myVPpnEK2FKeQG7x1q+TahnJS5ifi7M2F+LHM9MP27
+ObBJU12xhvy35AoNc8cOH7+1jo8zR/jwnIQDAfMCb88+vPtrRA1A1mSsQDbTuZs3WzFOpkvhqIV
5aILqG1MiAkl2UrDtk+ICP5J2Xwam95od/WgSj3TxsftYaDZG+J5EKy9N/NeI3xn7LiXx6Q/C66K
Vq2QLsHosO+N/Ws9US0sOIYJFz5+Or6ZFKljm/8rXgmxam1H05cCSLX6uKOZu+g6FVC37KsTTAJD
nJpmgAp39e/U6c+aTatQ7I4+dSmBRSYnkLJs9H4QrM0JjjuCzB10DbbqoctdcPx1X64mlYWtJkDv
v8yUZ8hg5/8v7QaiQSaLi1gZ238400q2v0+bGk9nHyYn+ScihYCaJ4ZNRPHKHjbRLDoyEEbIQtFb
pgkiqB+42IRGYxiitC/SdzTePWTP1IONsi/ZHoPUiPZN7STQYZha1+cCRYmRyIhzElLP5S3hFVZ4
ov5DdYFjUGNeTi7rVwFNNEEFy5GjcvUgcuC7RajfC3ZY80anuNcY/H4w9aaaZRSYfZkHamKnzQvv
harGeGPe1ijZsv0uE9yDEVjCak7VsidK4jEpYGR+Hj2/WtEQWOo5i2YqaC+GgYUolcW2tIlnytsE
Ia/sbH19s4IMp667R6nj+RV8mGp6Q0GxEbSOS1lbmz3O0Pcguem2eiQ2LBpRaW3st7FBm0K2RxrT
JKxOAQrh4ymokKcu4hkmW0acFbIHjTr7L2jsXq3RucQbgwIPh3Mo0mGsHc5XQvcYrFd2gCdvVUrw
KKFos4tKmXOR3Aril0GxmDfv04UjyAn4bJuBVH4DPG2gEHOvhIq5Ray658nyOuoIg3o8aoZPxOGl
NZQ0AQYf6GWcbgiz19gCtBGu3Q+ZljZQQGN1D/yj09mHRFJyfNwymCtZ8VFGPuxC6qHPn3ItH0O7
4mqcgVrawu5qc4toHhjau83vvuV4hzHLYiBR09kxRCgV/6cNvZG8b7pjjJizCxgT1s1gTC1q21FD
8+hYKhWVpdHVvXg8KailZXa/8M2v0s//mGXWD0Vp67uxjypaQXIwspuJtvX67tB2sSth4a6XbUfz
9GWfAgUH00fKYlmJd9XFImp6Ys123JYiCsDSmP35hHjSCSzqQHIXaiSQiFGYgNBZgJcx85gxRLhA
fs4csckW++EghgK3YbdvEy4WUEygnAysmErMOQMD6lWcZcNuxFFAuzQAHmLQJFAW/AY5wsR/qWUx
xkMrABvNX3KcBTBNLi3eqegaq6Dp80brvdiZZTBs/BPXN9gw85eqcEO1XfqWiZIUpL3r2eXPxkLx
bhrVzxDCXSk1WTCHi99fyUQjZ3X0AyIIOjDYKJ6ocnBsr3xY9nvf8QOJv0vT7Cnj9ZwHypa07Ljg
NknFUNVthYO3+NQd/9SqHH8r6FitwBBMaU8Fne2h7uSStRiz+2jxX5rSV+Bb97rp8I3cH7rGkSWU
MTdJlHvs5R8CpwyDCdy0gldpt2cEMAiS9kGniIM3/U6V0Cw07j01TlX9W/3zwFnAwdWNIvGExekh
8S5JDLXdFj1gMJWDytNGfJW7Dcmgn9bIOZ+0dHs6GMavhXYwNYt3mqpZU7w3tuLASwQ1SNBzmYlf
8wuHUIvDX1OqHCC9kn2DHdxPuYiBu/qMNlFQzDzufJ4zDKLEDE6ERa2wjufSEc073vHqfc2n5Ib4
yYkniUIJ+nfOaX4tmjMPZIsd4BQNWEz0n86EYq6+2fjhYtClx8xVbqq0C8JGiKXg7rujV8Q5lHBz
Fey8CnqirQ1yhirVg3qU0OrNz2sdPI1gLNBwedovnibQA25s9ZYU3/4m57tJ++94vwUUohIzLago
DIQ3h+j1nFJCCScXq75/vkf4YFk/EMU5EWeuAKaT5nnGTmBHeDTekZsfWaIhVmca+zzWYlVbqkwv
fYnus9DyuRBqlMHVUHs1s94gc4M58J3baGex6DdbeNyUy+zqqdZ41mwKv1NXiZoGMWoUNYDeRvt7
nheSUgL/vye/q9a5HDENITDV5nuJtmJ8hUoSyjKkDGL7PyhEG1B7QLxrO/du0ZOMhs56sZ80wa8T
IiHAifF1ZdR1CVNq1aflJ8zYJ4wigoLf1yKW4mtQCVJAf4CuEDNiNiJbVdtWJZyhXVj6KVK4zjvq
t7Yn50VDo8HsB6x0z+3orMDgHZlrZQfs2T7LlZDlZ0SJTWs5KiU86lDonaIp7AZ/t1vKRogUIqme
mJyU1vzXRe1yAkhVuyIB04tXuYS5wS1o3cxp4Rd1XKtT54g+5TH/QNHg+gSfeOsFDAZDO18D6hRw
aO9O+OUsQU0+a9VJvi1MeP+E7w4t+anxDrHKWKbS2T/KKVJpUec9sY+AFWI5OSOunD05FMJwlAkH
f1eaCTI3ZUv6sucvUGX7CbIFBlBcpUJQsv1vmjWWaTkzA1x0itQSLAH5bNITLM64wpDrraNeCyWC
n+Lc5hCfnv6iIM4qdsQdlkKjsaY7l8yK2IAQiUN6yMkEFFxsUPkh8HQin2BvJvn8ool6WJy1qYx5
bjUSDBPCzBs3SeGwTtDlxtaCaaC56T+Ecrn7kBtGMZtmOH4doIXe/OmOgbLWY1OKGSmy/xLMbcrP
0ajbG3Xe5p3W74qzJuyoFd+PsgAbWjj+PPXCGFByHSvso1z0U6fyl7Z8N407Du1ZVTUgtXD21RXO
Wna8WxsNYNl/EQZ85zJ/bp/LRSJH4X5S2xSB2qvxNxg8fsrjHL0N6Xt2URgeEaNc1VZf1zGYFaBu
ujcd0NPhGu/1n5+5XMrrciSvdm3QO+dB/uVXP0dN4etRMy4I9PJN9WExQNwgi2cIUOKaWpM1w2i/
kPHM9e1kzfWjlrp/VQxTPJCZ+L/apswKnRXO4DpKbxGp64b1E/sNmWoAzY5Bc15pD80oT70cZwKn
Una3s4vO+aG4uQE2pRv2eI88hOAqRz2XLMYaA50zOg832TX5thtmjN8docUBwMLLI6Yk7UQI412y
35wPCuIzTveiWewPqiOSMJA5SkdZmljK4Kqx0H+7Hv2rPmdkhw84Vc43RlLO1jbIGAutimCofylK
MrehOcfPWfSAp7QuZrv0lhP5BIEgzXTzD5/F/WxSx04mxrJWEYKnBHolyFWTXYx7ro8YqMjxpYlH
bgdieI49ccQUMeRq5SlEL7kkbEqX3cfcXC8hwq2Pz4tSh181GHQcwZNpG2u8QhCDH2LN7uNSYhCI
dp7Vc8xfHZKQgf4S1KqQjrKOgo5gdw1zRdppAr9DYNTzzSCdhqz/OCun57jj5oqg7x2sM5EDHlNY
KJDtmlHmHlyOID0Q111pFGiDmWOza+kLJHl6VIu4Zr1p2uDQJ0mqhMF31ZcEZ5xQNh1igVb6xhLH
Dl8azfMQSXkiiPzNxkOXhG7S3WwFBOMPTn0cANcZtmMb8WvYRUJs8EQ2IbNq5AB904wqOj7n+my9
DzaGtpVJ777SWGQTfKCyi0AE+F/Q8VoXTKW3x0HXSpvKT2dzVlsfGXrTvqBb8rwwmqDq8n/ORgg5
DMOJYXCExmhdjXOF173HTyyR2flFYEdTFnQlk9lLdFIpaYb+b4D5b0L4da5MdMoCfLZ/677slIBt
rwcJm0rj0EQVnsfVec2VzJg41U5sBBasoCbq1/HQLRCiXkmbZCqCk7fg0Rk/bY9mJdA88RLGT4uK
zrV+W6qfrWvnPp12LNT6yvbsKAWO5mpnMMt9ZjjR+zM36tcRvXpFZ6GEPGXK9pfbWfQEOaukiKqJ
v0uVZu47rfftKFspnNqjJxzXIYxw4marSyFjhMtOHA927Q9pMpSxi5rT+/p0mBkS4t4+i3nZoI8e
u9YaJLv+oUq6h0peF72RhV4f/7TfEWIR75ko2LLenXsqaBUm5P2ni4uUuSNtslJrCtnHvAuwekC/
/ITpRGx8Eiq+J8npAo0ffW9uO+dy0Ft4GxN4rbA95cAzQHq6EuEYJMgpupBe0gc0KXinmgDPJm88
U+qMPEerx5YqRHLWsWctQBmliSf/rWhVvWS24HCQ8gVVP8woEqd3/Xev58S1KDuEzJWndnL+x/U3
ZgS3OxUNxI2F9l/aWI9iaR/Pmn4d8qYto6Q/7Vin+MxsxdtuEU8xLsNx82K/QocZVme7OH+R42Zp
i6Wl2skFDHxN3tHlhnU0HhqWUfvnYd2zIYJifxfqbmYVuqkgMiA+24luKnlkZnAu18nCl6F9Lo7x
7FbD2D7jMoQLUhokBq0kmg68otPT6CJROPBAToe6QijGKXXno4B0qb8gR+YWxPn1n5HezjmzG3cG
/hTnbV+gQ5Tbve0So2zc6Jca5AygxIvN7pzseePfYAPS3dbgBe+2sYIez7XhmNvbPiotCaReWcgA
7SVGvWWE9xUYs+1XrcZ66sP/YxYUkeEGED/9oX/h6Cxzjr164SwpwMCWUooELmyJyHObXp2kMzt9
jBTBULxTBFqqeJZYnlEx1XUfkSBZeh9p8E/7Mvsrs0bWI0qFkkk6NNuoz6/O3kVx+dcWkGnsVfGu
Nh1lPVs839KKOi181k/KEArqyOCbBkZMxzpK2L2WN4QQ71s6UHK0LARzCKjC27DUqSMa3Wx+dnFy
VqBJtT/c39ctAGAFTCDCv+XFkqorMUgxqg6PA4rSY6qO615Cv5jE8mwqSFzyWNzz3wB/ua6cmVr4
qhQYcJzikQKuASm49m/e/nAHIcr1NCQQIuzu0B7JgAgqo/K6u9e4CUL2LXd9ImEKBR7lY3lwH2p5
0bPpWg/v+5W3pgS6CCwHrt5Yk9xDhuGfuoOhy1iCF1FtPdATPa3Qc4zdoqeqwFaS3NdkQKggFu+7
RYYnVaRb7u7lSclYWEatBoasMrIzynGWJUSKEfPSb45Xs/6ZcVbV8+xvIu8OKB4bwzaDx6BzVFL0
K9lAfaWvq+ceGDdF9kp1tlxVmeHY6Qhjxw9WO16ov1XgHGR+9BJRqA5rGotepC4cO+bbe7Eglg5b
iovrjeXWw6TC6MN343fc8q8lDnhuBTWKmaXK15vly0VNwpU2EwaMcViSvxohShvIVwrSVilt6j05
M/g6+l8bX1JCRzlChrYH6HgV9yoHeJqSGnzOU7CbPpiACnheg9+Z0wVTG8YvFxcU7aBpFkytfUM1
QteOqc2yucf4b97XWGLuu5DOFB2kr76rgntEQgeAzxdphArQagy440cTUzTRbAqRYUtFcJ7g60ap
8wDYhdtnkB4b06P6imRvru2kXCIUU2UAViVInBgLvrApKfCKRz+1v4hA9vVU7nWFdYo3N3G+2j25
Q+fiGZqRbzVlZaMUtZdiEAiJvka1ek5hboLnIAfRpri72q/a/wzUp1SUypi1+RwB8UI9rlA30eoH
Dqx0sDWP53vqay4FomubNQ1gDZ4Xkl+sM2VwKwA85x6UEZlJ498AFrvSezxwiONJgIGQt06CdHY9
qWo7QXJNad/GmEmAIDg/Qzl4cqsz102k3g4nTm8B625PQXjDlf2hQGot1ybmgDufnYde1FukyxBR
VJWFtKb0lZMuUowex0DhUedhsC1IA0yyDHjn5CDuDCzG53iKMTTF1b+80Qs0UGNIGcnYEXXPSFTK
ViZVFtKVMjGfNgHAiXjWHRHJim3ZbFwkZfnVZ7h126E2Wni9ckVm20j6Cby3EmUBs/cWKy2CVBMO
hDkx/pcTP2SezKxlK2OObqIcl75mncEjYGtbFi9QWH2n6nXIm8iKSx/1U8JnYvBA4E9NyVl+VU6C
dd4g+0iGIDHzr7Edpa1xgGYAcPZQMAI3xlgJsCV0YYcZgNGxSgZn8DwCce6V0ZkR6Kpjy8rzx99Z
poIfag5Ia/TskXDhkwx7Iom3d0Rz94nHYBJfVerdggZKRsNgqCOMmesFlQX0zal34qgZnd4ABo1m
nxo76ZbFUz2ux48/4Pp1q2hhPooiuwbd1r9QG3NjJDb9FGHQAt6NA8nuBpyyqEl7L1m2OnuEb45F
VE/8kzHBOlTI1YGO4KSi1R6GUseFaVj1rdySiaC2rLhx1krmX79RlLdSmwj9U5NhCz3oKOEKQ1XQ
TZCb33zVT9gdkL66icuUzj9zOHRIa8tBHHQ8CC1qCaE4PgJvb8/vzc76dKCHmsT/xlhgSuoEQvyt
DUU1eciWUiGajVBchi03dX257637mFGH3mgxczX2svksmz3KdB7muVqlqmkY5q2wU0gYEEgEYYRT
4hQ6MMduZsfQ2ueqJVyfpa59QokcJlaFzIc9G821+qA/DtKA0hGJKq3H7z1UeEJqE6mmLFlmfwrb
NilTnOm3KL7WDPm8co/53EhohaJm4MlrxXg58Nm3MOccGtQ5ew+2AbnKttehTYQzmf4C7hFzzROn
Qs1F3x+BJD983Jie2jbUWhNZ5pzIlz6HbQNk49MT5B/97fmdCV4tnBR+03GN/H45lISW0ZsTTkyo
vEa+5RD0/b8LyYgdkjX00/dJ4WaaGXCWKLrmZme+3MCPpqlf9tJB3962F/d1oJlTWqtbAptSk9eM
L1FLS9u/PiXboieCk9gRLNABMuu7KpbIFCky9qEm/WkkxZlFLsKi5pvp3y9+s27pO1EPrdnm7JnV
eG7N4vUlO8GiKAspnZXSISzov8qtoIdL/MXdZGMo/qWu6NdO7d0fJ3fnqX1nY8BW7xohbHR0FCaP
y6LpCd87Nf124GjP0NtuSkiB8ruswc7rlt+Tj3DaqZO5GcBvG9LIDeUhiaHQXq401OBR14GbOcxC
rTklqoTtqKYOE9aWm5TI0qwRU9tAIuVrAtViMPRQY7wlE1N4PCO8OkF64lakKyNUZAw2KO33xs7k
HWTIaPTc7wNcAMj5nB9xRLJcpdWAx+mn+IilKsVpA/t96NGjr/3ANW2YXS1sWUZLxFXBZ6Q6RWBL
4R9wkTjrqERjAUPJdkQ1Taj8HjAIfKDGn0BjiOjoWvTTUlxZ9G35/gcL+1pwl81inR7fpnhSfH+3
Wdami5KEYClgLgBdCrg0Hh1YtDxfKl3mJlHHxJ88VUnIRQBjoT+vp82i12R//cIPZBcsGCwTAQFJ
OUXQcIUvhQLe/Icn9SUrfXiVbAYdffKROy3bu89xC7tLKbNnmwCzoPjYe7AENDRIHU628csuQktP
jkZqj6rMPXNbBe0apW1KKtvHu7FeJx2RF4eDuPHFau65wwtcVOChCxkAj9gcz0To3ePK58x0nAwz
Xn9b4FO99SVxM8EaqFt/wDghN1hN84b02pFUpSWsIG3mkODVN+PmBJduYprpVkQinyAPVh4MAO+p
Oeprd5pfsrnjJxd6M0wBsUsyIK510OKkMK4aYiYI0pXLSNnGmH6pGY70mD6CM2+c5gB9g/+XWOUy
hMj2NPjItItQZ0CXzMcZm8IhFxpLmKPeOflx58NlFAEwbKZpblvEgFK9ASa4Ea1B7AbFQv29UaC7
S1+eGl/EvUYriVMeGkg6ETpNaRsY0o+7gEe/OPyKeU9woVN28b0dAiM7zdI9ePxgxTegekR2oudx
DaqVdpCqNHWW+RTX0dvXpAD3+LH5/s24n7tgoQYm9tedO/PMFjWm68EX+57HtnoMsHQjkqV5ZxBT
sP1KlN6ICaPaEJb5OAUz/dy0TEQN7yDX9b0OL1S0JaL3oYWW/fxzMNoWdHXGhX7jGty2HSZBkIQA
le5CL3IFpniXs9+yfW6SuTduMHswaMatfolBnHsH1kIz/RS6HjcKU8YaCGtLpJ+4/Hya/xlksBqO
U0gGfzS9eIjPfyoc6Y15L/za8+oiLwKh41Z/dUU160h4NaTIYxhloOlwrWPfQ1dmddpfuKc72BNJ
KJJ908vniYJvIi0ibrZy6FXwUfTiLEzHYvFbPTA6miINh3kRSawPk9XR6OUb3sGyR59vlhrEoYxb
MvfUbq7I8/Wuegs22LaC8vMtruSdsMgGc+8sBhXd3n0EEPpIvRObPeRd4UGlRFKmQgd8RBdK6+Ss
cftiR6InHnrEzYg0JjrkxNCDGv83srYcs6VNviUi2i+4TZC1fgGxmSR2cZHQA8zOw5DKUThlUlI0
O26fZuDJbqOFOi+HHpCJXMxkB+kTu4Ja34Bo/QraA0LZHGsfmdSaWUttnYD28Rr1cTLQ9bCEaWo7
x2x8mTRnZIXCWExoEyY2morWfL80eusDlWQwFnxemCFWVcRzN30vDH1dz/SHIo26Ei/DEe4toKhq
u0swV1/H94KujiStdg8VyA0/VneQPaQ02VJoEuzTkcJSSlvBgcOBly1NfZCLN3nHfyf8kUJyu0uD
gdjQwLDnR2uP5rNmeF2GtbupxM1W0ioB6GZnJ7Rmnl2WBadT+yM9yliI4vHOVqimnGj9znU+ec78
1pAzZDCAd3lqeBQYZoHRwdBe8eubreE6x63CqOnEVm62Iu2GQhuVlmN7nt1Gewj9X7l+O/DaEvrV
hfKx9fhCXvWisedBNZuKYnfU/TGsywdP6ZwAgAfdqtcgVYNBWpVxLLU7mnENIR2VYZ+H0++3P2UE
9mUv7MMAjKqCx6HAdkRmVpGv6hGZqPirbKDXdqrXTNF2hleubT0GVdKZzUr7Rbn6jKIMJ6AkGB7O
HQzB9jvBb0v62gOh857e/oSQK152HVW4euuZs2/TUneuXLOHOKvxxOiy4nQZrfxVZQAg/xg+vho9
7gnW1lHdK/7olCveCRTwxhFSjTcB2oJCWJNGl68qxno2XrCJPmXHdMGT1WXtTcv8rxF7r7AiKHgF
7qTS6gukXiFy97oo37fL7+ydY42+r7+BZA8VPCnRUtyQNyIx7v6y+pkfpW6o5sNk519StDd4du7F
hzTbJguopQ5QN46o+I5bMKJxp5DsJSID1hERchIinFoaAOnrtfBBBWzp2fx1EEmqc+bbU0b8wrKX
LTS0SN498+BJK3VwU1kwWAyVTaSjKYyL3D1WDJHC4KQZqdJZDf5G+oURbYBKSO7p7v4Czz6LXneV
8O9BaDu6EKwdt7TikVA/i1LIs3TI67j2Gl4h7fgGMLXiydeBNMNeS7s/tIJ62nuhWsD0113qiMQK
rGU2ckP7ZHYGoKac+tS9kv63XLQFJHWmH1k/kwp33MN+u0zXQWxltmLf6wA4uUIbip7WsAikVlMe
8Z6p1coIx48hRJWZ5IvX6ykPbJB4PT99eLc4KuPxrkOkS1LLK5QN1Qn2zsHM2op0G1mhxUy4uDP1
+vba96U0FybkOB1yqrcb84SJi/wDRuVQPeP6N2LqsFv2gg/NjwEdOVz0PFuId6GV/7z4Xji+r10d
mvTP5ywmOE8RNHrM70WKQHlC6K2O+cv5StV6IPFHMQOeSrMWVIqvs/rkodZyvzaZnOGE3lCJeSBd
P6Zn0Vz7VEF34UqlmbwavJD3zWB9+Tis+sPPEPiX4lwWKjiAEX7dh19iMAdii5wstm03ohJn2UYk
k3Baf9++IqRTNrQ/+rtJZLG6mfAs4YJnC0LkBt4EOH3ME3XwIFzkUiFww/l86gifk1c5oGnFNJ0+
/WysaddgLp1tLf1/RdOmUBe1qnkCPH96K7VEg+LLmPFe5S1kxypfzQfFgCnTynqG7VVb3ZWqh3sp
IAhkGG5zrEjype0GBBD5+VbZTKwXnsQ8Tgl7M8DJh/sd2f6tvipC5EbYKoxMilWhbX2FIKsX6OKa
l/uHSq1w3ydKuY5a5xLOYTdN6kuyQdhNORN3qwo6a1MYrSxtlAWDnLt6vC8BCu8ib6FmeHLCsLwf
Hyl/kVEpvM7ukRgmJMVx4MiM6dZCXtPum7pHxVYNRwCzqcQVxnsofkqLDtWtilTG0VVIHG0T/oTF
TsiHKlRkyEbPQG22gckyIkyROc22VJSSBBeDr6ZAoW4ddkG7TKcZDdPWOckbF1PTR6aUtzqgO5pN
TYqwYIv+osjxMa7TecAfHjenxwTFViC7Uf3FMDKwcuuUvTZ7HcWsrYJTvjy6BTDGNggAc6aFCTr7
7XuDGuSd8kONne4PynZ7a7fiz9ZOnhW8vdfyHIZ5y8u7GZlG+t/P3Enu2Hl+IwVXQ9MJMawH7ugh
1dAGxwCOvsz7V48wTXRxdcPJ5pFvpCaSCeA3qon2nxYjC6N/q/R8hYVkNs4ytOEeGbJTaUjMj3hN
psrEAeJynz+PSHjfU8Ku48tCBWsVWbjax/3A3Y5lrBqF63B0BJB4S0q4o1cY2Hg20huESt4T4hD1
EC1cngcm5lsAHcrfO0w7SV/UJhNibPov+Ff49ymbC7PD2Dc+aor9z0CnBPByUbxQ6jvHA2+5jyS6
zhrSwZ34+bbedDBr3mLhyaliLkwMm9O6Pm6DqbPmWVlv6uqJyVXREwuwlr5oCwPwiSejgAEIvPR/
emEtpbCbe7W9MtRNw127MDTu4pLoA/7BXJLl/+YkxUIqgaGMJ3ZGagXrANrxaXSrDUWPCC7M2KBW
7znZArpLPgrgAkwvpeZZ8B5ALFRZ4nN1sjKS8eyTS/9cTCX8hq17xLJD7uXptCnNajm+iXsTHK1s
hCb3wSOwrJbNUqj/haDwBe508KtfJ8ZMX8KSJRxkgNG0quOpUfJqtOjBgB5Qk3NkBhuGmjJED2px
v27wwg48vr/yxgLH6FThLHgZuYjzgflxB4TBlEncs8xcYNPgb13WZcPTmGI7PQKVbbBeQdKSEftb
Cy9P+vpK0a5V82YnGO9TDtHMu62r0WZ4TWftu9FoGj862t63Ike1oyujh9DJwwWpC+0xtuHcNOIf
8/4P/Hxc9OWMYVvGWRdw2tgY29RJ1XymqtDDwHQUF9khPKzr+dkIPC+M9DASQa4vOjFb1Dcoda/8
ImkfcObBRhXoQ1JOvsPlIZc38rXNylBzyZoB+Ynk/fqjm0p79QrOfMinX6f8v7qgwgbrlrHcsD1W
n7IEw2lv6OJC9UDNpYsvme/qtlnIFOVE9Ha3Idkjv6AeP+SG9KgLAA+TPVy/0jDEwMARSOQ7MvOm
fuGoYtnGdf8LFxrLFF4nvxqYo9jY7sM0U7EEeE+6NEmNFos3iQtM9dsE/+9sTXUKFrwT4yVIAoiG
7rP2+b7VVs1zlF5bfeyjUZH3RzvgdDChrVOkPqiJiSzA8hqKym55pJt5aGt9p9WEQBCT3Qt9r+a6
wK+1BCDywxOhjDjKZsrlA6DGMEWYoObiGnEt4TY4YZrzLYGlTUbMZS/pOV6F//KAd6OWKizfZL/U
lU/MLQWQrsY34X3S6Mj/6nYWKMv2R6fvuAymMZet1ZwSX1zXoSITftbM26voI2XzZNiTpHE10uin
8XFtNe6qN3i6dgxPpfA+65XcWddg3nM8fywqaUReI60acl7wuX1U04SGx5vJIeRo1BVUZPzMznN6
4IHLaP9mheKZptNvZco5ERAHWp9VxcigCIl6zj4LJc45EF5wXehwQAjT8XsKaeHaFO/37djdaJXf
Zh9Y1VVQnDNSmah3/LGpuPLyWg7MO0GZbcQF1tq5sflgvgnQiMKjlO+583ih15yo+f6fPwCL7B76
cmTSnjZJUxyn6ttKYuJknmNdLF+bC1Rc3ppvbgXaENq7gR48snlgYgtBF+PB9o/LwJkAc74KWUPv
hyhKdX6/vuDHvqMxpmpfW2adpP7ZjZ0CgX6GPaKjOSRh7Za6ZyRWFqYFwGj1kyfO0/pMVvS4ZgPl
p6qzljcHhJFsh35E/hHiWocd9RfU9DX8mfkRlwgbIJWVu7V5J3eY5qMs028r3oxtDLLXx8wrn08F
cvUsbUDW6WWafmku/sP/9JYQVfoNmfE7nlXY4gygmM9XPl4ka8ftbCaPIzp5LYQe/bA8Z5kR2z+E
mq9q7YKsu9IsjixfXtG/SpTdvjYUudqRpXkDYIhMK9VLqwiG+UhKW+/ezhjKQcBrVI6WvatRn1yI
bLBgYQZ9OC/awqY4ElKAAi1Dxv7M5OStwLO0fVDUKlzOEO9hbZaWdxY0/A7bjmh3pJjOYQk1apX4
SWIHIJSC44o4d6/G9qOBIsCs7/n58do6lyPAIVTCmLnpO0xqrwnEPd5SsllC2KKdvFi2qTApBjrX
K6BdshpOEFuOO5fMOInNAJlRk9OauIivb7xSZP6UZyARTiUMpFSZksnTPhGxhvInovPuNao0stBP
OrtDaWoWQdcCh/END8xjV4MunuVs1lPKrkiB4zDhTmN30fIZR6PGc34ciUUqjulqR2cocEFK3y9U
af9NIYd6gvPVHpHKcIS8AwqXPTsNzlL2YqsBRNM9uk0zr7peZwcECcxBc/fYdzdCYjO+aAOGc53u
faVt8gCjlMV4AC32avwhMhgtCF7mWXdXJfZDBi8UN5cmz1p14w1qd4nx/atpOTGNq0eLgQ3BMEc0
t7ugyIJuym9TKULNlNLttRKPgW8BoWzRLdkoIyJWJ7o7TaFJZrXcT9Ctcjgc5XV2yghlRmErXUV7
G8nZpm+bvgP9zeypdkG8XPWvizbioHB1++7TwSJSNP7wzX+QAV0+WvvSU+448reB4fFFNj83umbK
8mRWSL3e2lSAL95Hvtesi2Ul+pjZ9hOgNz2xXQ7E7D1H1x+R8oeBbZ6VEv4gJ6LFx00bkkjHGBud
A6dAGqG6ehWvgy4lS7DcKeZXx4qzYxR3TK8h3Ql+7ftHyk7UfjlwTiptuyTN7qH3Ppp4kqhqym8q
1IDBq0kjmTT6k2YzTT/y+OfkReloi57u9W5Bs+aVTrGMvHgDgk1EDDRBChFB7xg083VsLyitLKLn
SHxVTpnmcIkatXCnYNhF9uWmpQTEEpFdZ7WLAMzcsU0+RLnoU9rJIptZMqOK1aMTlZ7S8TYAKyvx
PbhOqUtW7UYUEzdrNSp+bFdLGvqEBSFJMaRq2Ylxb45sCvdw9jeTV6RRNCkSVNbPPuCvnhnDUZyl
e1VYB2a6G3eisCZYt8HMli1ZxC3z4Ow8ft1+K0BPwUO34qz6fwD2T29GnW8lYyQaqpSSggFZFhGj
BIu4Svh7oVd1HGl34XC8/iQH7DiyCYelGFj5gfDBo8ojkYCT0TZ3GYAwe5F3ukmzSfTMFLgcI9kF
p+ojHwaSckLGU2QjeMevyWt9djkyUBty3Wz9rfowlPp5waRGWZeDYNyXCXj5GQlVXrAZNNndySHz
bUgXi9FIF7R+4N+95BLIcC8xqC3wNfyO2lvz5T1FcAshVKZHCLnvn95ess9MKPamvpuv1IDaBRr6
nQ0CoEx6DTWqah2jbXzKvtewJm8WNNHqzE/f2VQeaA8LbahuNQFhCGKr+7rIbnsFhRGzk/qUyc5s
bCUOOe3xwyRZx5Tdno+XfJepdMcj4GdWk8YROMA7dUNqUfoIlV/GjomVhEJNcHG/enPn9pqqBJcw
OVYs1q7oD1oFr4F7ZJMiccHMO9t3iXZKWi1jyKYtPPI823RXICIubD5zxfVE0c/cNfpbWYmQ5tIc
DtzqO547L4S9+cuvYXmbvQ2V6WgqP2gVSlX2QlcWMTFGwalo+HRntasiCZvmLKHf8Gc56UyrcFPs
hUVauJZ06x8s7BMN5sU/T07dKu4HUu3+A4TklBXZUeXRWnb0qjbBGCo8vxMNQhsID1LFj749/F3r
A5sEYqJpjEjOYfn7IszWw2l17kmqJp6SkXWhaeV8fJfMzTbqJ7ZKUz9odjbkNji6KlOk8a71m0mQ
TwSHoPj8e5cJA9kcUpyetJPdO7kS8uhJ/Ix4jQsU5hBV0/mJ9oJkZ9IswdYxPOjEnQaVtVtHqBpS
QfeDMgylM0OIboh6wUV4kXSPVbBOL6nBpMc5LifWHuD8xl3hfkCUCqgYWawy36NywvHlFnp2mpbY
xYMZVNyoM5zq2KIBcrBjYH4NCHaBy3pvHiUqw7kgFSQf0hQadRhXhS/uxU6IcpsMgQAc31XZfxox
mVmcw+8cknS3Rxo05VH692UWKt5TF8j4lv4RH+9TJ+vTzGsN2vF61fiFNVQrI0Ial9Ia6I4IvWpT
cppq1fMoDJ+wTWTavCeMRQHYbc2l4NYCgpgDPQ4esUUCXW3ieMf873ToF4eiyopyFpOJr3EwsQoT
zZjHe5QX91K7g0o0LWqaRahBna8jeCmDNY8NHdCg3JHlVfxkbkZa1NH8X/p7do3qK88TObYiQEty
QZh34js3Vsj7tMuemG4uzXZpycaKKDA7EKkCH5/sUDnhbHABWSjx7qDjAyh+rAzbg7LfmHwi9bIm
2zV4zjmp7ND7xlkch9TQYLhakSnI+5sGQm1HTSFj745bU6gPTuEtY8TtlNS6pBmf5yZ3m3FK19VN
XjUpmq5swTs1tz+d/SDiui345UCsZtg5g/ClTWYAfX7/OKJWJ5Y9TNczlCdQDCRJdlQzEc1VYIBZ
59FjU3zgU8nSHeE+tjRNrErb/htqSmZfbb6sEYqWffAMFL0Kxz08M6svtzdnwP7b8bnyerbqnZUe
WtJrNjvDY0No97xGxxDNywclqex19cLflwOiB7ALJLx80PfO1AMCM/yCRbzpDfKwjQfkBswlJE78
nEe5l7SmQ8sOkvSuigXjQpPCwyfynIJG3DaJpLDyxlfu9ZPPXdXeyWo5OonsmycgwtDmnNl7rbfb
VgUzR9t6Y8HOvVxu2G7EhXNnoVGBL9dQw4YhBqjGzcdRBQjvux8D3yJgyk3+/xRHzBAIdD5OWw1T
vcBIPKYKCNWJxaeUG4rC5fczleRM+tBXldA0DbjH+2uL7Xa0RKW3Z0xsxsIlLNAgm7sFH78+uaN4
8TSWPRZD1+Z4+NmqyeIZaLQ5/ITG9ciPRHDOb/7J5/aaB0urKK8AKn6C3kCicU6DN62ub4s+LnNh
WyLZ0WhH4/7X1XVOINRK29jaRNG3D0dOcP6JHvPPrsuPuRagJK/40HbmRulOvHlxk8vqhGkZVXN0
LNAlr3g3elGTR6jy9rC918MhjrLAjMBGjguduS7PpMHyUEePK/4KCa8o4UDEpQjwkmbKS6i6ZcfN
1gUUy3iQymApH4gAziLQnQUtDyrAyOanVQcXYyKXOz1YyBu/0DjEXNuiUwCGAim7064pyeb5TqC3
kygRlf+WTYUKu0Dx+nWHpLPbq9AZE3CWGfgW7RPHeN84pm1Jg5CULGRR6oblIhKmJuqMvDhny5gl
FkpOlUIc+eIeQ6G5FaQ3kSn4Y3xh8GF/0FWcqoG/SOHi5jK41AOcWjimKkajsIXByu7Ko4R5/L6o
G8mla9n1j6U/H0DvoFusm7OjGnKS0JlF/GgUlDrTO/72OlyyG/R7AIU26kGT93DapEvJkT48Tvqe
mrUIwnLPQr6vzGSdzVdzeSWfByIbaaiYs9tI3duSDq+0RkqLgadCeakOGLYEqggKBlXv5FCDTaLB
PmFmq9LCFszswehfswHZBS7lnc4KUAU6CjHSoH5VoNsKdgcX/KZZdyjT6qLf5VpFf4vwwjKZ6eMJ
k83kzzvv5/PcxcxvTL02jHvLTCNv1tMvG47/gOgEmaw1cWKClKSZHV6dE4Vkw4C2iOadSSWf+lWi
W4c0T58IKK4JlMrjlfP15+FHUg0sIpH3SZ6AaNJuquFUZjsx1wW1OVQH4NddihV3mHrHAMX20CEE
8xA74c6UqCoRlKGBhfIsR4gDJ0jZNyL/rUn0RDCwJd1+NxdmzK3iYE4qYLwY0FtXVojyc8My0Orp
qVmpJZJK8UA9vF2f+1iQLoxPLY1c381O2vkqzn1u3vwK2Cw10W/Obg2GC8BvpeERJaXwWCIP7P5a
S0L+RdZBZyq+dglBo5pE6KwQuCvCGh4YnHsjSylWlH4sEU36pxINJtjpei3hgnCQ6KkDacMv9JiX
niFQOs4xrEU1ePGBZAuHE3CEUnEkQAzri4WbXmz+IUfuo/8eFQbcZPNzN4LviKFKlI/vRp2Jt+y1
wZoW08yZ9+RN81EPV74QKZgVCa/d8GQNE4H3zyg2JCODKeWjQGleZn5mxoeDOZ8GsPS5Iimu/xOJ
nytrq8cSzW4wBp1AYZsYxK2eSUp7ijR9Lo9+3TxFEUjMJ6nU+XeE6B4JHer54Bh6nz7ady8BcIAe
HuDUSBrHNK1tY7aL702eVA0XhUq4BTfy2g6MAX8TljfoqQOwINtCpj4A8ULYNjweQs2PiSIeb28z
7qcZg2+WWwSWOlnleLDrslWFbECJAxISjg1pQoqkWtkfpNmol7yf37xGWmIL+ZFSFv/KUcLqjZLN
Z56WMB/FOBtHxVdcUeMc85Hl469qqrahZcUSnQzAMmr4mzj2kY1Khq+Lt5RxTrEZ7yB/4xRO1m0H
aCT/CueweiY2YzBjh2tzgUOSExvobDqBK5gIc8FZOUCZUQF9QZDd0dWimGR7r/l/q03aAk5hivfn
HHzMGQHMrOVJjJUskZzNE7LFnthOiE+vbM/e3957vbk7ECYEEJUT/JQWPvakDHkMVvjU0BOQKhCk
ZySQME8ujIn0QpwKDk8Gar76mhS4cHU0wt3gbGn7ngNB5bVTkfjJ2Iv92/gmQCEz24M7v6+b7CPg
JoYSVINnTa5ShC4491QsWtMpYZOz+B2GSe3J1WiBzcSj+L6eYPlMRCZJq3kjLhdSeAwM69xHs6KU
WCi3tnYwfJKhur9XAU5961s+FAHsRxGbd7LZg4vVyYNrx2OHA6dBR0dr/eUYEv8ce3LuaqkITk6D
lB6FcUxVfNqmrnrXnlBKAG7XTDoh5vBnzBBFqwmu9OOwEjWJ+n3f2eC/vtBiZL1eWk+dGbilM8Z9
E6CXqSjGLnLKDx526g9ch5B+RfCS8fjPe4j1Jo/xDo/KptRfJnM3b1R7Avy6b529WSmH2ny3NvOg
wT0b9fhLpkc1iyyVk+F9O6UaaWgXYNh4NLkONsb0t5S6w3RJwUSNbq4p8lctbup8x39QsSKRwW31
tP57SkUoylIiSmVeJMdXJDWyG/cqcSNJWQTnsm1vF1+oT51U8mloaGaVs/WrfB3NUssT8IMqpfH1
Ly3AmE7/b/OCTTsUPXiBpj+1vkl+Ye1GAwVMKN+gdHi7N7/Uv1tZu5bROwWuQ6wrwioBdgfkBcSn
CZeH/3GfNlYdURcrte4zJexqL4QPu8wq+7AsS8y2nSlyhtpLkPJm6EB4LIqwE2Myxw+0JXf3X2zX
nnLHOWvCnp+hIy9MnEGsVxstRyprZvzvuCyViiLm4BtgxdcAACwBt3GuHPkUujvGGcNwDNbC9m+v
QDkRAMF+VbNdtslM1PuYiyjtLEGI0Nxea8/ehHvHW6hc6Dz/kiCi19Rv6qiIZiagHDzz7M6kYDly
krXOkG+/eGenZHAdP0Yec0bxUckLe7fs0rwnpXR/bRVp02lkBnphnWJ7gxMAGe1gYV/oINGgM4sU
LNCQymxGW9lc3mdw74qC3HQrKVELZW0uQ830AP33Jqsad1gj+CEj8VtPX4cGT89c8bEe0bEi8qm6
5nlsRM2YxOfk6EnJasb5t08r/eTgbUS8jLu5VrgT+DdEL1jNTMzTeHnygdf8zBiSUDaEVYfV/Arl
elR6/421zObJiP2fvH2C36CiMI6CH1r8nvqNFEr6EZnBhvN0so+IhiVLnrrUrkxHyvNa35a5pQW1
duM2dEPwbci7lhuSC4McsbkNXRtK0Fs+nc+jI45Yg0xYStc61WxlF7q9c7m5TbWXnA3n0BQuN7uB
k1RS34iq50eRuOGVNgQu2/7TPjcRCXGq1G8+fJhMdPiO7MwSWKI1QXpyXZM3ol7zo/N733tlA8jj
h5tGNY6aWilC/7T9kh1KkSTzi/1WFBL/EE59uZ5G9pvJCcxP88IUjv/16WkLrr6BSJaCy/NTfpXR
fDJqoeb80HBsUPPqoLvOiSno4tMU+k0EYh9tlDPITBPxkgfkaqn/eZYVa8oUyIwQnNlW/1LS3keq
wCY86WcuJAPJ7QAmTuPsdEpBFYKLMY5VtcaLgYGTLxaCeU0EKhthK9uwYPCwA143casB5BIIicZg
kXUNA+M5H7rEfV5r7VAWo1pdCsYYDX5CEIk6CBQ7Fe6AyojVNB5aAJm8c5yZeb2NHMSDpLpY7/HJ
VHwt/oqVcayjwhLfBGQpN/+CMYnJ5dcsfdyorUxixr/wzMVBNTPw1lIgtT0jfFh+3fbt+9P6DNoI
ou5tzGuwmTy58wWLxH5W5wICxIOojFk7+PNRrBvagLUh3vIEsTDC0ceo3MkXQfwYNLSL6PpTZGfD
dTlcajFLxUs/FoBEltZzJ0IJQN5G+gRd2S+bQ//MHpsOwZczc+0t0RzQ9VozRNGuSDKitE9gkD9G
60hOBN2/2k55fGQqawIOAUn4rMgdQIPLbCCe++tig7Pjqp70/X/ldidd4blpr6MNPILVmxrs3sgp
osvTX7rszaY75PySq32AZ+16L2auKKetcD2yuRD6ZXQOdGU41MbgGQLYo52bjx7MgnA69Q2RBNdh
+NnukSQpTnRQjJLqTx9fo1811qhQGVCPd3iK7Bnl840fmOlYBJgn8EvxdYalyXBbyh8OgxZBVtRA
W/6KGzBxmDNfRoL0q86IMekCiNeREVFJZXfC5pSmToJZFuaXaYkbM6S8x8nV1GiqkKJdsLyjkOFk
D4euN97f9MKZueIiClpXmjebDk2/PN504hY0znLbcUdtvr9OevqXbPsgH2CUroYHkpIubjuCWIS9
Q6aLAdSx8UTxO/eTG/oIYIVgEkK+YuDbBqhVaG7lmyzClc60bYNT4eROviIos4Rzf8wCCusG+zuU
IYabx52Jif/qlUTX0Xkb5O9gRXW5GaYuvvCWl9KE/uH2jdlsi2Y3trwZqqhjT09DEv9UYvY/8LWr
+511M/EgQ0cg68oBF+igZiftkglniB2eVj8X4Q1bRmMN9N5YdzhuuI+zUJiOlVDmZOINXH4xKFkL
BtLV3FAdiVoRsGLWyxmRzcicdVHvs15bBl0hurh8xEw5N3eTLI3JSOWdouQrtpGvDCBCkUq5El1J
nbA0jKs3qd0MOvHZ5Whbsml2O7ql07icJyqC7kMqCF6GrbaCRz5Kw33s3ITGyRgN8bpCHZ4Etpa1
UfXlxDQmonQkB6G5QzvPtir+m2hCpZk5su34N9fitPe2WfXcOuyr2zny1F1r1CdJQgiam1p2Bgfy
MNOfO0jA9j0+oVmEnzNmf+BFjmvBA6+dW5e6QdcjMxxk5u9ym0Jy7jRWLkMhudN+aa5MLm1JLyBA
zYGz0aGi3H5guFPUrITZJo3es3El5dHTgP1flyqdpX2a6AJLSdDTPov7rJYZ3vrkpjjVH8Qn3N5I
4SHy8voiHCtHLeZa4vJd1pGTpfqszBTXN4TORjFb2hQVsQHOmWnQdqkJK2jfhbMWqOJh85x6rATy
5RZkoUykIMsHTA3NIx5URzSpMgkb2Uv4NUeOLd2e+1karAIeK/9G0nQ+3byvECGO5IfsVgiM2aeu
iLmlOILHHnQPkRB91fN0EfMVFTA4Ct5VFe6uHIHK9s9MWkZM8XEZ5kaY47hA0UJS1QBhnJjEF81R
dYn2jQ3YfuVx9x6bhu2ryE9sdQVKx7UUt/sSAHXZoEuBzqW7uuedlki9tlppdtYJqzfvqJ0SMNax
jb9/t3KuHpCo3TkTbhGOy3A2ZVhGp1nClo+yBQeIZXXKGRs0v0/FTZ3iY4qxhFqEtH7v9Ecd9sf8
1OSSMlGAA7vv5c210sMoae3Fs7awFa29x3u2VZe8rl+oeZTMjg4TXwt9OIsj/4IBxWWMoJyaXntC
lOT3pwXHDsa4nkilfavqprJv+/Kqkw1ps75Krw5ZshfSC4lUJzRarR5kaywQsRJ2CW+CZXX1A+UN
J9RqMAmTJKLnHSLQymj532Jz+QpOG3oqENFgcJXcnxAOENT0QViAGy8Jrwcwku4+H6PwwM091YYl
wM2knX7txLWeeFIYKuFCKDFdeVRorYwDf7aEowGa8o3tuIBbRe3ouMHUZjx8cKNXqjLuFeHgYyuG
qN1+Cc0RqQQsRsger3SJa6i6Au9Z2STd8CD8SdF2k/AGCRrQlzY3wErNX2YETRnQEthFwZd/2Iby
jZDlFVpDFjzbsa1brG5Dz2X286iq4xAvjsq9yyJs7dC0jE9b/ZPr+Mrn2Q5L7gUbcZ3xfn7z86dV
FCJeEM317Ab1aMD5e//12yRPkP2jEzoF5/JFLCCgxFwOYvDC4tZvT8UHzYAnjIwhszDsZ4+NipRG
SaNveFvWWz5sCyU3q4PNP69LXZn3m8sw584dDtMPvOtrgbyiAq77KEIqKZDbFQAe+3bJ7THs6Nnv
8nP5AVjVg14tWhpccIRK5iBdbPnCRJaCzyfAeIy3Sfpjz2tkHtFXkIDmakcQ4z154eEda8jfVjun
7PJQvRYLZkAlTVZenSH8hbDO7UG0wyaf0RYoDT5EJI5YfnFANUw7pWlLXtpdeeyJPOaZL7XTTh+I
39ShnhexvJatA+l/LiqnJvaB1LgOxTej3wez/iu6MRpnh6ylx0JsgPkp5/UbT3IR5AWhrJeGUZF9
oDd+6jqpXbEvcZZb9GtUMbyBMnsK9ZN5jiJMBzYyEcf9Y73uRIDePYrqB4iOTE2T/hZTF6MFniEY
SgX0OZeaVJosbP5uVjgI/VnkdN+7XFcz0VGcfRh/3AVByCz195NFFwCxRBkBmWQ7ueRq0MkEw8AX
Jjrfvs9rlq2bYpqr7qmaIL91wabOtoqrw3Rxhs0XkgDtjZgZrged1F9U1UC2/i9owClm23LGvJ2e
tuviZU7PuoYKufIM24j2XwvRNADmmINH/u1c/iogQaNM+mvNaukFJS+fSvWRxiIzgPbFiFo+g7VC
W3VApaHF7UX9/P9UV+erwNG9e6pegdSnxKPSdejQijlnqRn71rBB2gcnmqffoMRJFKrmRcl7D7sl
E6zJaih2GIB0Zds6vmn5M2hBKD5wJBMR5kkCtqpreO43rO4B989VgAI2Wl6L8+EYc6LSp9e68G4f
ArS/czObMc3bcQZDo7hYjYslk1tehF2rCGNJoT+MxUOazGJKFa/nGTPB74H/nQTdhyOfqAe2XZaB
+MLXZaxxSZXgqB3pnpyisHoaOWAFkkLIjcMqChHy/jt6nHv4gpH3zrvwtUi733iNL0y8wCG4ZWK0
hZu91K/HcwFuc40Nj7ktOm1jHt19uOr4n+0s6C7MMAINJU9QHHPrLZIiRJteDuhWC4j79Ogd8uL8
chzL+n8QQ1vNJo2bvATT5vyfiaKJQgiE9KOgfGiiqGkK5u1qf5n6giGxyyhuwXK6ZNB4AwEEuJbY
S6gcuQLiDU8us4L1B7mJvtjrA+zE8GoBwRqUFy5h9Vdz0eaB/LzQbJWgEmybpQ+jpBI8pUMixTm/
4kIQw6k0tgM67Q3CS4iaOpMd5loRWncOapEmuCBnZ9D7SqggpZDVvmB1DQpfTWr6GEoNRRCLQOYo
cD8dXM2d10BfrpxQUlRU+dBoI6DxLpPYaPVNTs0evgiILJVCEJfyETDUBhEM3tQoEhcjVV2bfTOl
wpkaPheKDG1Y8ya9gp4YQ6tSIgwbByDYyJGxwvW0pqEWau8S4OXg6Z61lBadRA==
`protect end_protected

