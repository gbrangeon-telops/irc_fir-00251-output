

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
OHeaBmhw2WWXga/8pOVTMIzcYutI6Mhna2kzvZmeKvttg8GRcsMBDXpogvkdmdxp1KLLzWXMAKSV
fUAOBPVAvg==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ao3tKAmGrk9jDIJ5tmEl5p3MIRphIc7Vg/SqO4TER/rFDRMS3J83CwQ2b9YFrnde65FSvizCvsTV
0Knxkw8zoIma+TSgIxOnivhI3WBhgKeA2uGkUI4h7aI3JKyXt+ar8rATgfMIjtkwwZmXnAQdFAm/
DhnKD9KmESp1ihQZWxM=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
tIRCJBwrqw861TllYkYZisN+3Hf+P2JXRGH4rS3/mIyKaeRa8ciKvXh+DuDwE0CQ8FK1JKt0o7Wy
5niCab0pNdgMIWoeJTN4M3Yv3mIYHhxe/uhUY+qL9dbTdi1peu0ypGwB+pCVAaCMnYsMP87ovoxG
mFxz/aWHoq6z5hUiOqs/8QctFGTu5uGrqo/fDpwnQByfUDzc5kOGUXom+7Ix+u0CBnUzxUPMVE8H
FW15FWlEhZ2/WOv5odw8POvTaQir1St/I4TCBaM8Ne779Z1F4E4v1nyrImWHcYGt30Ex/kdASWup
x0rIb4g/F4zfpMwk2F9PI0IRzfsxsXBx1PSZmQ==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
vDR9iZfmcKoc03DxzsUkjAUcoXZpLGp+jz9oB+bhIzk9fA1B+YkBJ4B6wGhxOSVsIGzj0A/2+sve
cYv4/y/PnMWoVJu5GAXMXsNWS0+yhRlFm65eqZTnif9T4BQLUfDB3Poe8t8+8qJraoiNha1dShh9
FtnafnjfaWlgFCK4DSo=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
P5OVsGiC3k02pbA8zjICborh5BXFBySD3cMhIIsNr8DZdx+UrjbiVbqZMU9Ry3hJ/1iX0Q8zDyFo
F6W3nmvV82n8xeQJN36fxUpz69izOLDYVC7B/XqC5I6fwrewIKThxTuK9lZtFdQHHrzj3T2ZDLDy
Z1+PK2wQ4cNjjft1DSS07aO+6gcWXb8X25cWmNGk/P6Hl0pzIcfFFHwO6Oq+bJ671kKmsX3jUKAg
DTTCgxx1Ex2XG0j8cWCnhZjmetyd9o4fKBdb10goxmIXB8/8Sn+4BcUJVLUQkMnRwy0YJGGtpiHs
ZxxUU5IU2sy5csUBb6rGbP4ap8jLGVFhtMQgiA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 16944)
`protect data_block
1IMweyZ6CW/CcaZofhrWbN6Y5f/fkt6O2tbzM9UzpqMKvZv0ALBJy2/yBoqAn8xwE5dey09R3GYv
w89mV9S57L61pepCOW4cnkow5QCBdsoc25zgMLCfdoR+Foc2O+92jpgQMQo690RPnlsModz6ouY3
yKQEZz24HVkeyogShB7aJcSHNlpCxD3Geq4txm1LNWO8Ov3mj+zf5DU98F4VC5qJhAzMaVj9cpkY
hSNKAZBY8+vo13HLEhvM3st8dWH/xQ0Tw92ws7150el4xrPUu3QZYhT3cEB/OIq2aloM2gbAv5+B
4+6b0c7SWfVVif1EPN7Hby6ey1zIq6jc3S7MPHp2APZB3iU5lIRgzqrAhOwnMvazatkUz8QB5E+t
M9u+eBowtzU1k5WSfQYE9NapdjrFV6Oeo2clZS8pIFSjq+9S/LzPIdbLWSVNrzTdLJ8BktC+OOsH
q5/IygVtYYmtS7bXTbHZOnJ9qlS8enB0CocCrQmzqMhWrTsIO3jXJAoCBv+ve7j52ec58SGfL1eg
32muypAiWS7/jTJmkFDC3J9SKmHiBHhMp7kD6QjLm6MOdfjp4V0EGpyV+V4RSlr7io0lxtHncIaJ
0qv5GT1oT5msmq0RgnuzP8Hspy7f311nlayDRkrvdDi7q+UkkJJ+UipLVpGCaGT5CLeE/kxyOZ+Y
84rM39FHJMp4UKh6J+fksKurKhNhEDyMRVW7vVEPWnVX/RNtC3LgAuBWV8mNJ+mjqEb2GTv/y3ki
D+pt66kLGWD6epkdJKmGqK5VoZC8KaeVr3sD6rns4nKZHXJ8I0LhJQ0OHV8DH0tbjmGN4oofgmcG
z0J/cb/+XfQ+AB/H/l3G8K+9sOr5/UKQ02bM9KVxFKIkLQ3LuDIjOCkBKn4I+l5ZeDpkq4vGn7o9
eEsUSnqPZh9lnooo9Y5VT0oin4jGxH40XXctXttaNhw38buJK0AWb0BOKQXHVMR2G5K8fKZ7qVnM
fElaNrCKhX/mGUlvw5mY/sHUKfMArVFazN6icUUmUtrjZWk/YiIJfjerMKZTCDXjRq6dcxisJmOj
jZ4auttnAZI19OGgedOpDeO05RJGD/WkG5VFEeNoTmTq4RbPn0q9Wr6zfmKaGaPrdr0fOaxzGgpg
A0qMDfMIcJoppmkeBnO9J+UO0kay5wAgkXhvfYmN0fUz05xJXT4yiBs5V7zIm0vWvvNhyVc96WiN
LClXwqkYp6mtlE4r60vnl1VzZDEk0mfFFrdxFFBqmJ+3AHfAGihgZfC6NFxJkXuE2NEZj2DWK5W+
0SRwKktOBoLt8OmQAPufWPvAz2S1w2dxVt944bn4yQSikqq69ONX9Si/dbm5DsGuIB8hd1y41w98
ttv3Pe6qaJOLxf1VCamUeXbCJ1F8yu0mp9cIkgjtR+hXrvkMYsroumwe2CTDJGuvUdWiPFDCYmmv
EdYho5OpWFwn+q4zJYNWtPEcuUm+pTEFHZRrF7T3dl97zCdEVZ18aTfEBKooTNGUySNh9cvBOiIo
hB3/QnjtdpB2XtQOMDQvytac9bKb4UVie8XxKkk36aBVmr9Ab9M6ANlR1JjFAQqIf+Yw25YnlShT
iUc8hdfEzWmksP76MTPuVQMoIOcOKZyZHGM2/JlVr0cnNWhyQqAh5N53YAz3CZ69Iha5vNG1nDfk
y+zQie5YQISc+NYtl/mMbuCv7apy1HKv+dqmKCISXaaLTiPjE9DOCn4070wC2njSredUpBSzkftT
0mF4dVVogQKfEHXjd1/6oEX8c2fwpTdeBkNeEjmUp+GFUEXF4ZrMQUBbDmw8McKYO7UJ7W5GfHSl
OCzB7508/lZx+5kJNiZu/Zqbuo0dlwX6yXk3aKv0kOEbqJL/zQ447K9M2CRfYdo9AgJ6SgxQs23m
Ry4Qhka2128XUdR1BQ8iOZJYqFHdDs3ykcnJBK7ijBD7pHABZuk6ItrLONN7re3XD7BL5da5Uqp+
aRyGWgkwnjl5xsyi0uWezJtv+MuySQi9BqfEKazBDgCgielz4/yavjVTdCScryjR+2/sAbIgp5J1
AfrLCiwR0081A8CxGFhgaALZ2+ADB8dlaF7B2mZ2S5Mv1hHdya4aoeG8z5cTAyJvp9r1V8UzItJh
ZbaYWhU+6X/LVA+keKzmbd6IMKePYJvKp+Mcs9wRUCn/o4dvgSnlkJRb+zK4QlakSKNgyoOxMhdq
+UYuIIfQBZQNIlkk0kiQI3N01NhuukgXtKMC8wS4/6QQezde8fIJOX3p9QgSJRwQGCvCaUUyV93G
VfIyiNVRvtZoFf1jKhnixSKbEZ1uifc4RQoeyqjW5pZ/fdUDZj/K5otkpFII6jHXgWlYf8vLrjX+
xNzbUvXwlotA3j9alA153n+r5L/slUwUVB/L+zS9sU5aeqEzk2fZDpVA4B2jU7fuuHmFD/F1UiUJ
5mQNQFFnXD4DcXzcpqe31tB4eT7UZXPa6lca8H/kn1hLylUH4SyuJT2jyDHChzwaokec4s8KM/WK
bDcBZYNuYER1wQVZJ7Uavhgpei7rhMH27O7pkLo6ROiOLJoLNUB8u5h54C6/D8PDg2lftsn+9Dcn
8Mk6dDID1qTOvyKbOETbKuB499wF8tyvWXSYYUSwfj+4fHme2mJHPodB8M1S21trwPgqKr3bQ+bW
J1ZmTUQw2g1Rlv4n2LHQifBc5jVR4uTiI66jvWk8ox6GpsRyRzl6cr2YyW2XfWwMBF+o7ubt7NuJ
+Fax5iFiD2RsA8OQUDddD8WVofsxDAg38V1XGmdotR/0stBP8t8zAkks+RecIXxmlxnxc05sv5WF
/HpgfAuZS8et+aYMAdROIAX/jblBao0yZ/mF205ndSXeA/r8pI7/R3ga6ZUJBtC8wJflUa8xY1ON
FetML1DUi4w+FWasTbhDPikE820UYSt/LNow1YMQKd4qoDoy5+dFmtMSEvQEF0ZEWT0sm9wjpc4z
w7sJoYg4etv1hs6hzbV6gFKrrnM+fpd1Vlj0gYpKYH2fCdyuqJZ0AkVtZQgglWUfIhDjiSkvig0l
xXdFxhqo8Si67RTN3HhnvTkx+cBq0Dtg1YM00oyffnMVwQjE+kVP41s+idamcqBxRZ6STp7zrLaA
0i0CJlEEYfHtNqnjAl7NAwCTDFff0+0BjpqahJiNvpiJwMrmnlM/PSJbue1/9NPAZu/dWikElhvs
E4xuP2SvxsAyHA7mVFBmcTvlrvNd2pEHAg8eZf1lu4gHi6Fp0AQO22rEysRxYjnH88k70m1qDzZc
sOTvIlde0DGe8ICQa0VZmQQviC84vqIFwW8Sm+zAm3VGPVGzI/5Vb8weexmIxpYl1qr+mIdl1CAV
ChRl8JKtsQOeyU5bxlwpe2BFD/t79dS+HQMDHOPiXHEPuRdlNqsg/aLoCEpq923FJyrPVM65OM6Q
nite1KmIZrLDVPYTund3H+oWGN21KN0lYYDopiRcfEP8cMpw7cSFYA6KBAvYBqRsXU3pIvbxkuQA
h1mcG7Goxnfh1cM/+cxDlvFaxKiTqBb8+1ajHc0S+4wdw3OwhHOANHeJ9HypG7u23l2iuETYwGzD
DuUoPE3bPXD/kzzdavjkMqjDO56p1M1gy7mh9MOVCZVYJRHagjPjd5yTximOYb0+MReR0VPvN8HC
yrUzg9U2lvzyW3DUT1wTNTTIvORZn7+4a9FjkfWMnYdQXvY/NleNJ4SNSeQtlAqb+kC0La8L7WhM
aXfmUCX+4rQYM/7mjpPRmlM3zcfHwX8LJZPfhFql6gVHaQCEBOjeVoaZYCRUlnMxC/Gh6SsTF1NO
tBmAbpakpPo4vDUMSUzveeMzAUxL+8N10npxpKRlKvnmgfW90bkKGEz88CxAzwYdLkVq1LOuxID+
AI3CbNVTMrhwK0ThzRh7vCayt4TYIDp+cVRKfmmPlVrK5Grb173VpwJjgIQQtAPFWOn8x/bRLwLo
OKobn7hW4SMMUOZyRZNgINMDHXDq4/pe1he2emoeRW7fGqwOn3vH9UmHhWySTzJfTz55o9n1a7UP
D/wDrfABPk93sLzz+8xDsmPBpySXWcc53fjt03k7UxovAJyFd/g/CwnVYcdMvQAXBgMsK6GvyedU
dl656LGNMBCq4Ja+oTV6hPCrlUvS4SAp6qRtvg0eVb/KbZy+hnRWrfx9RIP2ICZokAI3ZvlomuXA
2Mkt8UjpVJEtd8dxcotkx2ixfTUif5ifdKq5luJ8orraiKcx8hz7uxBL+7wwGbdLA8dWQCWXAdoM
usU4ivsX4F87/oyRlkcBQjtczVxh2mnkX86umP5dox/62FmicXmU+9cIFTWJiBfzKV7tihzQcAPq
9q82NyYvP+R2cXeelVTrNwahsxmb1tcSrLHD96HvLzM22QGsiaO8ayfAXcipCag3nfyLMv49hUzX
+0YYnM7j8b9QA6AoJ4lByB7SJE/nhVVpXiwU/lxR1imUujSu9pAWiVw6dSYhgw4LWWPP7Fe4JuI1
K+0auosY2980ULsFJ0LTEfHzywlSZ5lyhTcfGn79f7qSa6cOKtfn+L1R68FA5Ap5XbKT0YdD3P17
nyuK9Jho5/jnFJeLEoKGZxWnH34kNbipZPubSzRVF/ulOWizWBgLhMZcBxCQDj9KMvJdkcZQmO2M
mLSsUgnQ6/zODCszFugoiuVacjCh9kMWRAMfmQ/4EqixZUOW7CKF4DOtv65oSkqW8J7285yInuIF
GavWvjEFYMEqUCkRbfaWt7mn43XosofuQPYmFl3RrYlZ3VXdM4ulH1E49qvday+tZli6qA7Q0Oz3
ikkxQSGb3HHolby7jRhpZkUgPY5jO8o2oLCDfV5/46v4FtYcG6kVi59rHD/Z3UX3WVfj4Xz66Z1v
yVTyLEtDmPGyrogLK10b9PQTS6xcm6wYd4LHYVFX4LsMSxiJi5aA9njz/Bl5FRi7MWNHwUuHMnJE
Ex5bT7sKEzzp1MerBQqBr2uQoCcC95nL43qb71gsEYzU8qgWvf78MsVLgeXNz8xQzb1RN6ekuHMm
RRUbd2byzEJ3F+1XO+ezbCZt8qpE1xZq5rzh+K0n32jVq4euffmVnTVyHWIhAQ2UI7yL9Q1Je8iO
h2FCZKoG5bebiYODqLB95yuHpfebvhV6hpQyAd5r3W4qUk8G4VS1ek4yemhxo97EUecvSKpSYUG3
XcFEpVveWRDfHDEA+RTF1MaXQbq7iVbAATfc4NKUtm12p/csmHTExU/mAPFDDKHgPijeMreNzAiF
kMo8yCLwI5EhT6qdURF4OUQlRb678UPdIKMqxjc7Sau1U1in/uOddnn8pdtkSCCcsu55MhZwEegy
J7sMhwN2t+CN/xPKMELU1uVoCjqPjmR+hZLiG38I8urJxk6oLWhlYAbgjZHtIB8ITZjd2uipL9zR
Jc7JiHXxPrTKZ/yO1N7tjtVwGtML581nC99d7wQt9WwGohkxFwDJiU302Y1Dtw6wuZB1wGoo3g+B
f5lvQt0mgS4pwXNDJSsPve4okscIUN8GaYkE8+dgkOmDgfcANkz6t9mjouqfw1X0CsgaLwYsD3LX
97hE696puAAS9B0MXlx9QryWtW9jiJycFP1KbGMwsuJL5vPd+ULBo3IYiG/bw4xYUQLkl5LbXLme
qgYa1uVEKffqttgb+m5N+uY0RlvUt2ag2PfQUgXFqngyF+kpufrJXDPkRCpCEKQYNEdvFw+Bwpgo
+SIRaPBe2TDV0rO9b4HqMvpoqJtr7GqblBl7s96YEkbxS5W1dG07b2HLaz51G4apQhZ/ovSSryRI
1CYim3D+5UocqdbAU4ZfeTrErpKjNTz3rqqF0VkQR5oeLX4TbNenjg+LFopv2ZXgl6XIIJM5QmP3
VcNr3fPk1ZphCNN77znzTuKeM6oxNbQw3XH9qJklvk7BXW1fba9IgV1ynWWJBbKCUuuX1KEVvMMJ
eHwKPUsxkzoAk5rgaLVSSosOKsqZWtNgT+cK5dxgTg3jpnJCPgB2YUx4BzXFZ/vquW8FyPDBJXlO
1KbedjHqLOeqPcLWXcvdNWZPJ/31OQuY+lQGBJI/g0XHyY1UIQgAdSqYcDTM+PhtNYctZlaKkK4u
pDmMI4zAgioFw+5o2O91d2Y0WHzKwp2UK2FBdzBvuT9GbCwcxWujLgBzx3YEq+sqDOmk5hle0MUd
1Ri5S00mUp41CO5HP4FlTTtcspP5aA/bSQPMLWTo3oAP08mDFS074iZ5BDoPH1fRa73vsGUviBpb
ntWqhbMJn6r05ZdUPonRwfHEuQQaaa1yE3MopyMihhXfThzeWeWNnNkE5M/4XLMu8X/O9JKyQH1x
lOsXv1uGedzs8PYq/s8KiwJ7N6/a2J+Txnn0nZjMv6lsZkS2BTYx9z6zgPk0zMTPY7ken/2kyFnd
CSy+gW1kgAo7ItaJ8AQRjaT+Ta/Zz/Y7vhETGDdwcsxSydCwabw2zaMnak8/rsaI5pDOJCuJKiCM
L8OYlFvZJeXYLHHGLRt3EZn+IvlfyUqeJK2y7BEFF5srWSbx/YdWWZ7taiRqZCnPHATtcxhHDGGC
S7AEggOPdOXuTTPLMt/Jlpi2W7V8O+9TleFALbeVWMm7v6V2cTOhVbOcnNv0xzqsM3gZ3ZrmvSA1
PEYyerjqb7BPzb4QXdRCE7Chn9K0bXng6hBghZdYGnP7yD7R3YYfHHphCShVsdFb/SjKSLDqQWrx
aNFD830eJBWyMk7cMGP6YqGiJhFaqpPRJ//TEiB6x7w/GQFDkxeaF4UgKiWA7kIvjKsL1M1BxaAQ
SmA/lQBLoFaHT0GOMDcdPvnwnid+a/wRSVsleVdzIyURrnbHnowTX9RATuF8SYCjkrVlQOTWUmsz
O0QPC1c9BtaB+cjRO6jqZ5cYPJvKhK7qqQYrJnhROTBZHPuE1VW0KbKjmn2G6YIbFzZ2DBRfi1nE
Ka6zCxk0R1XyWiCg4ftJiSHxOrIcML6GhsyPATcHN0p/EssKDkn0Vj8cnhBXfb9txZaNOAIU/b2Y
KLfsvWUV6JyXGy5dsLZAQnGipA18R6ETe7WSPOLt96esDj2Fk4WrbTJ2+r8X8cnk2tmNCmFLkXFy
cYtz2//QLBSWNdgBmcSHiOobCSBG1qSk+ge9la5GQ3MZYqS2VkJPLpZlTI7mJAyRY3Hk0GfTYWOX
ZiZAngm5fX52/H2oyOYnYgYdGp38d43eyTpJM4CLZthYbDu7p3R+Hv2BDXKkvkg+bs4VX2xhl7Hy
qbyBLXEgS0Rsf03KecwugIq2pgbqlKVxOObfL2/IawQbwCu66LF29g9A+ETnIPsqyoPpeTXqWqto
6UnIYfjpoleTY2xMFZZtF8jIGSEmSjqpbXzLpxZcY7kuQqA/F21TN19DNQ8R9Zjjulz+kYjSIvVu
bj+3y03a+66ztCEO2hJ81w/VmFcvUslZaIZzsq7OzAJ+bTnmojo4Q6K1m7UoFHM8OwKQhpYmlA0R
jZgEGFQUE9aOcoOusuLM3+yLb5V0ajrtqcuGGYOGW/L6ULvCqko5y5MjC0f9qiUzdNF7t3MIagqi
NJse4R5kDcnzorIG2AhWbJsFmVKyKYrOpFd7+uA1pumG1RUTtmRN2zRJwOMJVYVWuWu2MimFCvpU
stmY1ZTxslt2b9HnwPI04BHXRGqbWAxVws1pOaXBpIDHIow51oUbq90ScBpORkgbRRT6gIqH8jCi
rHHP4YxuHS6bM52zcDH/mdwdVaDMyFfM2/Unc/WnNE7y0sF5+sPXM9WJNiC+maM+wtyM5nhbywxQ
iUNC5f0PEEVMaXav4wtS3940kr36SomAtm3y66sRfe67qlZE/f8U+8q+KFc27xGRHJqbsdGsMgHj
swIdLHuWStXJQi6PEJL5j51lCtNTg1So6ejj+9q0WHSGpeRfobV+SP8tr5WP8u+ixkm1uOIiaSGx
EUBhRoR13/KgDApSVQf7KwlQn+d5DxW09RxDnUhPE3cqgC79LiR/ZGoadSRExHso41PmLF5WDqiw
CsH2+bU4ykASej3Cvbrs5huhmqrELpTTkt9lEBxUWd9qREK3BnOFxYL6v4+jynoQzm2AnlhauBMA
1VhWgoweWNs9EucyDuxObJ9x8eWNhoH9aAQ0B4q7LEHgrD/blGDXFwKGAPIcuj188oqUq5Daj5yZ
q1FiT0c60AXtA7hvgEperA/Y4of1P3eriqClr+w6MmQPUrcfrc2WQN/D6VCn+mt4hNUA0Ye1iVJT
M+7p0CMxCMi89n0aKl9uU5HqiB94CCb/KrK5ck1axnYFWrdgyQZCzyAeMQXUpS0n1whaVDLaSUXS
yrGo+5S96TAaWhdrlA4p2zkDX105q61/GlWBiGzIllLJWwMf7KbwQqZWjtMFkXdS8Aq+Y1IGSFVK
4a6THv6LHHclkoFuke0pT+wVAstAUjpUmVLV6pz2NF4aYzBkQovVrfPdyf98PTAvGKPECAld6AEd
ZIZC0DBwdZ6wANk6Mq+AH67LK8SUQ5AgAPdZWg4dlJoeyo316/EbYE7663Xm2yo0OsXm9WTrTIL5
jJPiiVIngK/kmK9fhoulUjrxz4WtfoV1lTnrWnodV0wV/krTCOVmbBgbXIETzPDkP9N1BJhh/Qtr
I/JUb1WX+z6YA2AahhsaatqkE5vbMqxXbk8jJ4I2A9UuzAscf0faD43+bRu0rpQR6MIDEL4U/yFM
PStPLJZldb/B8tPRANH1P0RgWcRPVjFru/8WH441ope1kS5Wib/RQmKyGbWxGP0yx2HAETcg4VPg
JjyqF0kZ1pBaIzS5noLmGpV9ju2ZXGIG/JoPliP3rLwUQXHjinsRvG1wJWr+9wHiKYy15l2FwYM5
ctqgjraoKRSg91caxDZEPok+u/4FhmQ6vVbUyW6gUhRKTuPnWxBnru13KlXASHwuI/HpwCV+wXeg
ocLoag1bQORiLz5BkeX76s4XG1eF3bUwJQVOpbhvrLMyutt5ftd6NhZgQz+hi5nja6sURM/aTWfQ
iNM2PUZGBZ0I62wK2aQ/zIc8yKXGUSge82GaYX+A4OSP8NNqX/+FQjf3pSagb8mtJwQj+Pyds4Y4
PkMoFBZO64nRyT5NC8mLDOnrmNxFXqWa0Sw+56D6gUpXGQl6147tSE9ff4OHfeZq8BnycmcBFnYe
SE2gOUw+uRD3gw9c/V2+ekK5VgKbNc6yrucaIlw0NPmBMXqH5xtzbLDnfA+dirS7ov6MdBiFhLeI
LkvgNKTGRrhKIHEoh7ZX2PZIeuryJGo9FZ5yIiynDrl0tYM7sg4Augnn6KcwIpSFIBdPYRJyTf4L
bWOcJ1PqebROsYt9HTR59Jn0jTToYflg+70VgNUT6Qu3HQqmlTrXYD/ZPQjZ0jyfycUCQ2tNvAIF
868Ay709jkcBWwECHoL49LJhcrO7L9YNooENN9eYEZA6rMkDiATsAKq/epoRCb5V/AaaCSO/LmRO
jErMllfIa9/Rlx9VCihLkE8BdDGZ/aQremC86Ss6HASrMMHiBGNvKdoTJnnQkXacitbRUUkUG8oO
AV6QCkk7MOTZcuVLrmtsMPItsydzPDiDqm5AoZslbp9V/hBLkk2n33SDvuna2H4rNHLNeM5Id27r
5W8vvFCRDr41fjqLZIkDcMdElxvnelezS8n4L2Bg/I49JYV+R29ky7LgjMBPTa2VDlL6mi65P3A7
OhnAPvHjMSENrb9BsXlBNrB0FR18dL4re1mXFK1NXohj+Q4LL8Zx/4Gv9BXnzab661eIyiV4o+Bg
YGhnxIcOQmvrfzoolMbYY23mIUSeRdzOB82gbb2Yww7fy7uRX4plK/7aUvyLAsHmnKUL104DE6CX
9TEGhnU9cCU3hbNh9Gft/FvMG9vhTucAcddTSHmm5coPpkyIlJB7AIORIZnQSh2REiwbyL++xxiO
0Bkf2YFKVrdUyTYOpv0fnT8Y7YF/YJeuOb+mBQfZg8ZzEWRp9EVz5U9polQ0w1njzgqs/4J3vGMJ
NBnYw2WXHm55oedElJq9BpcRTnqyGjzuKpGXecBZVLigqN33UbfNs8kxx9Y/rWn1dUm2K+F9dQnF
GsZDcJ/aYbvt4w5mVd70qGx0TreBmCZFN8jHFiewzZiJZ4w9evjBAFjdIlWSC2reLBr27PbQ4ChF
32aDI/QwkOKNKDhOb5my3tncTTgnM4tSCq+xp8y/z/ZTgBxoHQA08vsqTp97tZrmkQST/lF5nxeG
bTUziwVdrRyiLnFPteAPScKratS5PhcdcMquTp5/D+ejEU65tPSHGTZBoj501R4LBL5MRXTg+i4E
htCX7Chg25iRym4L7JQjX7hCpJBMQDjTsrunODmdbommu14CSruXYQigNDVnzUAtrV8KG1sjqtW3
eP0jsrOD1qw5r80yl9J8TCSdpL7gJJ7VkrQLYU1TBKwB4Hrm2r1JOwzIdFRTKIEAZF4hYDi3S2L/
ryFcNnHttIYCAbPmlejjDZsiNPi1vgGoH8oUEB3+v9W6yWtgXd1CW7f2gXKFR/uWaxVr0tUFYQ4v
aD5XZTTZOvUhGmtCoFCey/UQIfSTYHZgtZ3f4pf4DWbf6Ar3nkhDoFrjzQm+qnhs+Se4B53xmBRn
nwmAh9t5ftKTHnh9F9TEU8VaQnvU6K/1PPGxF3VfDIyoD8fq8x3PD+99GpE9HtCNRzrxHZPoQT+c
/dPbKVZO6ptKTpEoC5BLMuI57AZw3P0MObPPjFX2mJ1e8/zbr6Kbo7JwhZie1V6DZVOU5YsmLuu1
qceENoU3i/BPwh+xCcgaO6In2tPrnPMSqsAo2NEVqOLY6mtcXT+pJNO6q2oJCYeOJ4SUhgx4sy/3
UIQxlxK05Hu7LLdBXGAoUcmMLHto8sG/97qcJgnpqBkIqJ/TssMZPfmrHkoOJW0+uc00rkXoMe+E
mUye0VmsDgwdG0PXKX44WLn02Gw+oTZgI4lYDBLWJgbH//p4jWA4wXjADq7GpGRVss9iGRhKmCY+
/JrIFqyADpxZmI7Lxs4gnvhu3hFq1qJCHBGGaYqYiDWtbZj6YD2hPxwnukNJT1B5H8GnZIxcPRFb
lMcGKJYnWCARExxyK37CksC8iy88KxC6XyVTcOAK67tgfK5mu+CXzpHRCY47fDQjqbQUxSZPG+78
qKK366TkFMEpjWCn2dR2E4FvDAVujfw0uwfgOXVpmqu+7rmBcT1mF3fOg+3j0AWNStLEX1udieE2
2ClEYAq5FnqGDx7qvhKrfj9thGSe9kl0yDggX2TX7Yz1B+RV4nEY6DA8sQPfPIutWbIPCsC6iSr0
+ki+vqBT63Ht9wu0A6RkiK+JjlhetMgHohFp0dsfbxqgwBgByX/vEH0BoHgid0d1zJyzosEFPerV
pZYGSRCtsw3aqSzkmfcZplxWGWtmOkXW6DghOU/FCH0QtF2zRvUWLeBrsVWCwKnwgxWWplz6bxez
SYblnci1TQgbkTStiXStC81unPLgJ/NquqKixpSOaDAP/ZElQG1TBe3HlLVKl7t6L6y5wbpYOe4x
Y+MiG+47oT/748dGM9C4LYeo+/61w74Qr+cLw0MQJIevxDXXzWd3Q1zhIAHblvb7COgPnA1Oe9tF
BldzjLB/WQq5JfSXnAx5yu/4jEbAoI7zmnGRxZTu+EiWLN95KsXnFTtzJuBLihvVxetieT1duWWQ
9SQQL/tQGd+3t09q5tfV71BSEagvO+Gk5K0nMueGsXAzWkZi0rUrAEvKJ+1XhcP4sptVAwBi87fe
RIRq/gH0Wnzd3glNGdbjpN7Px5AhcIQTVJFKUR5ku9tTc40dEOEmnvAykFR/SpWjc9UH3Apd2rst
QiFmqOAeNg15OdWJ5qu88Pm6imPucaVMjIKCAkF72+zpP8njCj/lhjFQgCdahlzUycLGjAN8rqid
gaFAbC1TvudRyRHmBDuUDiBptxYcnkKPbCNJ9Lw/q0TyKWhUY9lnkvki2vZUMtEIPj5Ky840xcXL
4bZbxwomq437Y3Y4MAJUXwJz7z5aqc2YvefdWKpKqhW+fqKQxNjOYyhUoSRV/G97TEebQ4YVWV0z
Fll3VZZJIqnx3+2iCnGtNdnQqiUzcuvNeil31pwe5b8ndOn7t60fGKPKN7/Rs8SrmF3wvDA5bdkz
hXG86iwWe2mUfEagK6/rqpoI4pmrMyeOO/KhcUB41iI4Ujq3NGw3gFRjjSmMKsw3XuKbi4SN5DOE
0fwx6QLG6Ig2nZoKGPxWFWOioeboG2xtdg7dyaDkdYOnmkYnc/69huhcHIj+qMcDGVNe+U9RblPj
wh6mNoHOjuK2lLJpka0uHeJXTQT5GNr4yW9sW1HzxM4+CgOOXGTkRLlerVNWH1cdlc0DmFIHUj0c
Y7Im1cy6NutCGu+WAeRGImTjlt8+dsbuV1rl9vi1QgoMjnIJI5ecyRT2H5/tzNVzzsqX8raZtT0L
ivkBE0E3M9byVMQrVhc70PZS2ohQ7Mt+xnqCnHTi1eGrtl9t7pSOEDQn4U7Oe6LWofiZ81BtatGO
ms+LAivon91SAGWJcAWWGV5acCOY2MniOpS58jgJYaDedKJhuNx+++M4uz53iDK7zWfX2EeHKg+C
nvTr9bEwh7L8BSjHCP0Gwc4AyimMST3HxVmAiEjt7bfO0t/JrbcLBcxMlg00251wK/3gHoqG2z6x
pDYUsWckyfWIS/vLcnYWL0l85TF2IAcmwI3KXQO3sgEOQRP8TnMUINlhXcInyb0e9fXJj0710ySw
mPGEKEBhqQjlL3IGRYXiyaSMU/ZpNCmVJ3RSnsWD+yuEu/dkT7kPIDyjx57ZT9hykNS/HldAciYd
tmtyBblEkwgD9R3HRbFCxS4t+KyYUsPIRa0tyzIt9QnXL7kEQ1eDmrp46u9B6RjVE5wvB5ecoL/f
zINam/LQFn+qtAzeIN8DWqXS5IFfalgZeB59auuXo0JrbfqpOMBxnqa88PuKGLt7VPLX9h/yOdjX
WbG4dP1gNhKoOIg7YLGugl9/vquBd917pgD61xWxMpMs6MEEvlEoHfp5uBN4Gwpj8G8gG7OHcIot
KMRVAPrOuPdg8ijiLKpi6S5meShvXNHfiPrzrKFD/gFs2j95oRg1HjZSblDa8fPvM+9bUs1rixwY
HGvjlqfMo+/ele78YcIZPyM+Ou8blQCXCvogKl8nacywTzjOoShTnp+4xEWA9A7fOVBA1pxnnoXz
6JcDLM2nUXjHzdvLfu/yGpszDgvXdH+7ax2LvVX7h8oU7wAhvlNCAMbXWYHijbmdmV5KoGGJYFTp
RLjiurqY0+x76s6U+ljSwjpgqxOIZAmPcN9Fjza+BzJnNGFIrAXvf5X3dQdQkq2KVpvdilE6rkp5
1MP5KO5d8V7yzwn9ucZ3hyArVKG4CoqyZs72SwvVeS700CKvZJ7j4Df2n9CUWi6sjsQEb1EviNBc
RVpX62B6SsqbT8N2AUFnLfvZrsIV9ppGgbyU/jhCu5kOoOPAhJvnEedFLxwmpqqMN84/E64kBslQ
9juXcFwo2f5QIeGj7mumDmlLpcckMbY6ayGD8hHXkjEna5yvCRsMRRf7cz+NL/gylf+ukMV14tDu
9IGbKg2YFcWRmUWE++0rsNiH5vhZzM/q/marD9o6aAKWIGUt2vp8VOsw20sFLS7twHTOBF7h0Btr
JtQQqtwRZ0dY5PilN5Dhy5Xc11QgQZpSc6gXdd2DV8lrSoFWZjYQ05QXyGhhymlYHxac3+RYlG4f
zPErnvQ6+yzXGI2UZIMqYWVbiGPakHkLKO8ebzhp5lx/32CTPQ0xwRWDe5QPZKRZtd3oeQP1SDOn
fjLQwtDxoMHpcw+k91MnydNiWxqEu8yueuxV75GFWhwWV1uNPzhJlHXkBfOdPnxKUSKfgJwUdJS1
dkhw+8gKBGF8TVArl/DFHqrQNtzNaBgt+HfmLkguDEr5QBxh7PdYg6Yj7Vs4dBfcGB3YDgdPpE2c
GwkU0fFrOz1K9TdqsnvhZiIKDrCpOe9fWD1+8jdy7QKylVjXiFHUwdJTw/qmc4b6kGKYeCMcjkSI
iLF6enEYShEN1UGS9+TFo55/x+LLd0fgvkXUVNZVHfeRaCWYXHGOpvcVn1kJi1RP1WY8tjTobKzF
0nG5hek3LYYuhxe/axSl+G+AgxALhZQEyTRAOJZUJuWgZPPUkzzUto3fvR5bY+dtXmvN8llT8nlP
auStNHXBx6cXkgPo24qnsbaaltomM43GWtwpWhRycBd/+xgI+LykaHDXiVWWvl6uT2kWnPf2BZ8E
5C2HADOvMIbkRdOE2aybW7UZUxaISOi9c9iiPYGrkTdbG3GI98ICM2C+a+GNGQoIrfYw+UGNHA7R
lbuUIt5IPn3hjiuuZFJoft3keLp9WeSr4RvThQI7d81epQCMQ8htFYQIvQ8QdS0Yulhqr69XzhJ+
MzUdiG+AjEhhjBnGgCvYaBBfQ7/dPX67H2eYIXifwx3rQ1t4ZID1Mwr89er2SglHpHhpM7tcn8Jd
3O039DXI+3Lz50wnJQLGrElGn9r8gt8hpNiWRhVbp9Gb/yIQsjtTq5GWxqByRiiOUy4JvwfT/6nM
wJY8v8qG2omHuOjKqpnvm7XSsJq66RL8NRH7QsmAtIXmzSTJioUzXXaQsmBMJe4aBXTOa+ZtN3bS
kSnTEk82jjvQWAw9TIcOZ9p2dsqNJw/zwQMBzGDZpqYYcIQed2q5F2wYykgmLYRtxM34TzuDaUYA
qKfL+dw1y50ZzHSHmjf7TBEuBtnzOn1Zwxt2JbtwzvF6s3GhSCjjqMcE5RaZPknIOIKjU35LyPqg
jpkQLkBP4KxaI/8YqEdn+75R0mWXh3WqD6Z3BTbItlEWbUAAzeUFoZJSD1VQ3hI8sdZ8bgmyG9uq
jJoFSmnKzRgis4B5MBjI+FJvxHmStE8Xha7IvjqEuvFC9JZjSjWXNdh59o7q3g383x/+1oEAYqNT
kjun/K8+7Qjhiq1ENAS2V6zG6S1dMBxVXd6LNluaiPFj3yRgS/QEG7Yv19niaL6o33Vd3Nn3JSID
AmvnJ9J7xex6tSxi5zc28zfCi/Z9BCbyXQICx0eY/ZeiMCzxaVq0OtdSrUk3/8CGAvcgsYcxii8P
xgLX4rpLDx7dXhuqIYzDQ/gbHSasWXenZOMNAnkqqgx2JTHzwBmomkt9NdMRif27u5Uwjyu5V8Z0
XFes5NpzhtDV1DEmbqbyVQenZgnQPp8vqkBRVySv1se1CczH4qN+dLENJkz1Zu+4+oU0Td0y24qf
j6zO/cbnJnmAVF8hIXFu0LHeM+h1gc9Q3De+KsCi+wr7wxFZrtXX5woAKkPN+xUZQ8DsM0ZFaWPM
XpETt79obMBVlMKjHDAqdilZOlDIws6IW2AERfWgexw93K1enAt57HDxWLKosqXpLdzjyoLtLj1O
oGhwnZXzufTsuVkj2FFGBrXGRbS3k0MfwSIKnHDTFw5xX60Mo9bhSf34a62zoqKr+Hw4+JG73eDC
7lyphOCYEM5IKq3SPNZLBC4VIP2o6eD3HGniid/Ej2A3EOQW31+h+ZjfHkHoy8A7DYtb8b5QKbGO
AHe64d9O8xWJXEK8bC5Y5BYFnXUodRPS4tqsDg1JTTYEksOTUpM1+vneqnCh7ASEcwkBJmb528tX
i7r3e4B3EMicNxwPQLYsjMbCM8s519rHZuiLNZHFhSm2EguM16P6aKPNDI9UsoNcuEax5ov3BTn7
zDAkmWeT6A2E2op46xqn4ShIrTtPNtPSlOJUgWBV9cggCKKscRoFA9HJoe5lHEOgs/8zd2/DjpRR
SrclwDwGir3BXqoOkszkyPuDVONN2rwKG3E7JuxvG4hEnRjzUrTHdZUL+fKpfXeyHF7ceJL/sXSq
drIf9Cu6IAP+QO+4fxOexLik2L57cAul+n0YWkrWwv4fnqe+1NQrSClxFBVpB8Rcy4NzWRh7SFEZ
EuY8n50kxM5ntm++roRTopli0dcD8zlpMHwRe0i8uXToO9RJL8oV97NQeIHV/6xKqZH3kSF3HRyX
gOfesaIVp2tBPLMY1Z98O3gApYa0bShpeqP1TAJSlneN9C58GRihneUCEG055B58hbhmkWH9f+Qc
J2WQLCveDuyOvdXAAdZrGDTeQHklQ6we8YD5jMMIjsV6BgTbzCckHF/rf6u68mZeXpNxdb10pKDW
+nQzSn5jwkVDTwR1AHUdsQq18ZRFlBamcorF/LFA+cNyD9flnqb4HJHUKwKhDz9XZDIedof7ZwLV
kl9kCGG3y52j8sJx7N4IDRK5pTvfToKvlfpJ1IgiK3YmmMkKJ5/uD4H31Yi+gCwkHUCxUiSEN7lt
dUGKOP4lAm0e1P5+0Ybbp8eFVtv4Nr3nOLu6jpeC2DtjflDdwsSBVJTrPYlo6x+ab3o4T5e7/zwx
oQv45fjGFGNZ5WkvN38MoxGWocUwfVtQCWo7xA1UWq3YBL8tKM+G0IHkY9o+ZWvqpy0HHjkRG8/h
o6QP/iqCwzR+xs+MSHpDDb0RUHAnUGcQp11XMvimJnM91ZzvUStgSHQJZnT2kPvAEeCl8FRbQlmV
dRJSwMQxmm9c/1qPT2ciiV1V0dTbzs6Ga926oq2VBOM5mBlRx1vU1XHzqWUY1SYXznFSXo8pOU+L
yu00mnvPFnQrykoHVMbDRk8ioCgbStlFm0WJ41frJ9T/5gdbk717qqtcehxawy43MqYD+ga/HrYG
NB/o8QSxhdtOcGJZMXBmD12KkOJSwSibPGthdIKe+U0/6k0Jgc+pQFeG/mc2H7o4pf5DYRulp3m2
kgZt62aDVqPRnVEhEHkBnmms7bR/va/+kymXu4uz7YJRLzMPmMuKsXTykBtbIKHatBa4lnp6r5AF
2e3d+rsaEWQlYJK42Zh9vgJ4fzAWi15up4uP8x8GNaHmqRkS+G6ADJgGacdzJ2sQ7DxIlx9lfUVc
v9iHHYsJAJShcYRMsjPZ9/3n+sSGuAeqIoOx88rbl3wRxgE8awGYmFByfCaOnhKJXNZXW1eosmTQ
1Y59HPOEeN0UuDRx0TKsb3A+gSwksHuAFuHZkGWNI3JCdXREJTkh5hIRx6FjxQXtylOBv0jQMcX8
zrGDTotjey4pgaAvj7/Wo8X4Y635JKz3w4+0dQJde+Q/gkUj7W50WRcfqjSy7T7mf/R1pmYC0iJH
wjm4sMxObl59P+EfS3OqPrnNrewNcEz40zDU1Gn9yqhKdU1KeEJqXc+kikf6MUZd0/SHAsz1WSvY
hVPZNwAD333QUBEArwmHaVOg/wbKSNbEvjiuojbVvxCYUlicDYiiYwlF07C8XQii3tYW6q1I6pyv
xJzsWqiHENanVIJXQQuFwyCjzZqMn0PtrhLNa+UAJmeNBKIYMVpIzmQXNE5EsscmG2987kxS03FK
jSxze4m6h+fmKVY/XTcpcYWz8MFsdr+pK25ECk8+LjChqQuHY32H5PSpM71v8ziPeUzYJw4coG8J
72eDGJMY2GBevn62/rGxrCgJq8yyIH5PGsXUUQ7kjq3yayuyiabPRaEkeiPeomgHB9gtnTsLPJQp
KK490D1mSQveRujZZBPeGdkefBKCR+A7itreXHsNlFhM5Dol0dkAV4LZH6nllNX661jQ70z9teJ3
7RJR1WkF6OSQLM2p2QSBAKqhwKHS5bmMQSrLHdE8Fhskm/rcBR/OqGUBQPD3PO+wCmRxn31XL5Kt
LOkDMkpdRi+jRVS3Ki4UBwGmwTil/1XJakO3Kx/lHgWMmXWAn5yzQgQt9kNILWSM8pIiSsnwAUA1
qm+LzrScc1ie3obhAYCubpobvePAYGhprsWJM1j0Q3j0Vw/ubj8sJcaPV8GiJhHx+I4H/RVv5pE5
NoJWFlIRvU7f3knERiMYhgrp/XD1a/D0PchjguKxself518LjZoZe0NYses7r5xaiAz2VLd6xCPk
K8C8SZFbxARrz8xRpar8nJEs9jkCB1pmFmKALg1LJyJiuTytyfD1a5nuhpFYO5BJsDUlTGaz0yo9
Lqd4UHZXa5xryrypVBU4pyIYhE1Ucxb1boSmPdCiOqgiP+1hW5oyxzKFdAMZcEEN6Jxup+5qD2ho
HaDbRNliXhjpvPvyfyamky4JcypKAAem4VYV0Bbx41s6RCNMxEXyEL0vbN1hsF20Z1gnOn/0tffM
JG7bBj2lFaA9tRajR5f6Q6VCbg7YPG/9/8N0qfdkrKM19oOntw190LHNibJO7HLooWndT+Wg7iwT
fhP5DNUWg4kBItKlIiYOTvLiUwn/rZNjoz61aAGYl8CKL/KCGQ6pJQslel2Yqd62qehYRFqBVJjo
tJipvkZGoRyrAiz0nsI/7VjX9sqOLRsXWn0Dh2QNhvrmx4hgAhcgoqpVIWQl71juONtELFusGLEX
thBlJDahxFHHKjh0lV+uIQiEJt3CEPBcAXz1CR95wimlsTV3awykmx6oXzOsFF8OvRkGO2wH2zjo
FFcIyNyPrSxzY+YRb0GS/R+qlSlpbt7BhwBZjARPu3h/fA/fuUsCFNCN1VrTiYtttMK0+V49rxx6
o8Cqno5/so7A99GBAGhetSvz184XyLbbmlWLAm9fKOiHz/ITcObOaNSzBe4n8IqLS5Tep+62Sffc
+tomCv8vHdsQRqHdx3GYaSyoWjtsh44r3Ro0jYSXBIYcUC64oLjyz2ABb3r80ux5iV6V1Cc8LPW+
XgYND/rn56c1FQjCbdi06GzgNzNyDLcVGUqQjCftLWknxrg8NBVPuGZtxMrloocyMACDxb+Dytd9
LsS0Ke61jJPGxL2SZMda5uQFlawj0Xk5KDr1SrR0q/UjE74f5YNCviVt5EYvG9aP3cUYNsLp0JgQ
rzSyAEkWqNeQNSERSaoXmLirz5zvUDob9k55agznc1e+Za3kG0P0mJbub0sdVdHrq3mHoSx+8JsE
NBgUyfQHT2i/cogPgPIsnUhoMwbYD2fy7939O85vZCiCtxhczLVejFYaVKT+u8nRtQzTQXk7YLpB
I5RP5NuE2iyX7WEdrHPRWrT6mOTeAK7witf7xivfRUaT9mubO2ZjqwV8nU772xK3kENe3ZkvAKS7
cAuEOjSS3zyW9grT0+irsDnpXDcMcfXajIcb2LLIlRC7y2LetOKZzK1ZxnLVcHsnGDrrXIwQMSgn
ofkNmx0Sm8CQ5W0wMQWWp3KzoZQabT1YVHzKaOPCeLB3rSzqVURf+y/GWBMnEzlP135pXdJX2qDy
r3rDHA+UUD7euNZeUJILm+zoBM8l/NTS8FGxu8VISoeofQ/rxK3zRO8AG6QS5l4vnC89T64fv2ad
CMRJOOi+ngoP2bXSUVKJ0pTVbRAjvwMJRQ0zG3rEO4TNonQBd0j1OZQNghpyHfmUTtZ2owM/DUTa
smSvyqof2P1xzw/pmKdfDM9SFR/1cW8GPP14+4GMYoZBkAiKYNKL3Y9I8D9SbV/qwqWtfFHtXT6K
+Xej+Jt0lqKaL+ew5bt0npzi82gyNXAd+OhUWg/rIHhUvw01eee1rZXujGhWFB66KPu2ueosKHfF
KQhuXaoVQBBJ6rVVuWz8kXgdKtlA2MDxSOnCKckvM0SWfMxHv2NF2hKzBqbQmEYMZ9/GUtzcCkgy
MeyEzWW5ghc363oUloj80RxrGEb0WG2Lxb04fwsDUvoljffcJPczkte6Vp1C2IpeY/O49uwYreAP
BE0AdjNdfRBK/Lo0lOXFHnOWYUqNyVecbLgFITHJ1botzqmzSsa6X1Yofcv2SVSDF5xNAbBa9K8M
0wGe5OBWADgVSItEr/X6wYBZ+hCGaglzo2j7aya/UGhSW+/oKVAA2EBJfFzV6WQK8kGbfpLRgytE
HUPu3kR4FoijCSDW8RIuU60muIL42OcM13c8ztZHSkAgdVzRAanoqId6IzbfUWLtHU3kK/OYEgd3
+L0Oy64bP3x638Mmyeb0o/jiyt1gIz5ovgLvTVtAO4z6qsDbt+y6Egd8ujrphJfsSdlXRD0L0/fu
KAGKY3TBXm/p9BCCIUtEGDHv79E783DvQI6D7t/6l5tmg2k/ZAsvD0RzdRT50uLd437h6e3LUp76
bUVMJ0Chk/eaPWYJUrabO816ixftuWYqj6a0hArZnd032OTZQpE7PFu79+wq6CKizebKM0X/ipci
KLlYI56zp9keS+76ALroJbKxDhgxDcB1qhBVDxHKyXdqDqnvR4hd2rzV2SDqgzPCRqtv4rNd7CLq
lDPFVuXoSwwzvA+D6YpRrW4TiLQ/mv1t8P6g4i0NhgDYu7ImSG8Hf+RtaQJisV7El5XS+3LokWqv
SLSFTF8OSjamfzoxlmE8Py0C+TcfV1Q7/HM233gRGkA9COn0Z9pG3IGU/qyzHC/iwnF4lziErKrJ
uC27CY47oZagwdAi25Rcg57n4eyM/rjC1HZHR1x8ovJywi9lFW97gQyU4nHdpNVMwMhfiuZGqPy5
vyRh7Bf+uBtzN6PAn2+3YgiUNLlvlGURappruXcR9FoMFC2hhsZNEwIe/BcobDxlRywX+ftnOmeB
pwuKCVM+kzejO1EFozi78ltr1PqmVZa8eY1o0EFy0E+ZIJFjYDdSiepUrnmllfASx2dVP82tCVlR
cCBh2w1wNsMMZ9B4Cti/XTRrPNBFYn44zE4UXzx9haY2OvUgY35jnYrBOMygZP6waRhYzbZbgC7E
JoI8u4OxdVxu2v/VVjnEwS+BiP2Wz6M0mQg6FP591nF8oi3L/BrC7CqTuxsl3fdYtl2SZaHQdDBd
Q8BirzDrD0XZfNNXFSzCkPAeE8ZU7r7i7ZhWmaxyrhjoZOIVivwPR5owF4Nh7fYLqI98t3GNli1a
O6GJUfWknUsIhsXGx1Ky9oqXRukOMxrgExqcku7NYK0KYeFl0iJ5SUUPDu1Aq32AU2/gPDhxiT4H
4UkrvNkwCPe/2HFsQquuLdHUvWUL3XxgKK9C6dzHao1fRGlIWgVh6r7wIIkQkLKHqK/sIINDs0ug
b3ofeApJjplz9x7VOsqaoro3+d47YI5zwwLmFDPWa71cRIDm07wFBk974jqaQkw6MhGKDDaBBJOg
+sCZz4KtEUSgL75fPnORocWn+1tlAsWdZcsiBobVbz6fFPzynCuIxgdQaA0etKh0pK6VwZxEmnKw
pvtUQiBHtjkruv6yfpEM8byPzGfFb3Z3ShU566TLOVXIXbX1LEs2u4itIu8lSpvzRyM7uc5KVM05
vq1/oNOpZuuG4vrYP6C+U6GF7E/N/JZUVPaLJleyaHTVMq2MPYCsGBufxn5ptGjMDO/HAFL7JRme
SmHh6DJ2zP1Ui9QL533sgvP/fKMnNsOnTGyOeS41OukGFBI9VnzO9GAhRLn/w6fN0xB67xlZFcRf
AUSilNEiOPbPvZOJdlxD8uQBLYeocE2CfGMwPBiesOiggQJn4gYqfWcqUHRLdrhJ2haz+zEawaif
7vqABxzHSrCDdNtiszuJ9ZruLLgz8bx5i2v+jSypRXZx72EE60ysWGwpI0a9usruJW1bC3YTbfLE
T0TEaBbrOWtuHnOV93lk4tqiT7U9O7ZbtGcnpoS7q79Pa8KiFXsp4nq5C7Q/aLNbJVqnEAGnH6/Z
Y5kiyhc4lsrtYUHwa5a9jo83zjyWRwSVDmHjT+aCttJD0u1/nJBLs+rmBk3GLYbyhvQD60QwoYm+
rO9dRdX2gGWRFNgBiZwbTDAqAL0FgBTxlCGbHgUqUjmSsK0VnD1EdduJQJeU1eWv5N0hW6V1Uhib
iS5JQQQL/I0xpiJCAv+LDf0q6+YI2seg81d88S6p9l0eZ0wtxhiXeL0LW20ygDdyJPiGr1Lk2kdX
xRolJAaDptimuDo1Zoi/mGRG1icqhKYTfbzJRrfHgxA2TcpbVsIz6h6cQC6mOhz+77zYa4qBRiep
EUHZfE9zOeo5U2HBPmwLj1akvEn+WEq30RBvYJmshtS9J86T3ys+ocda3Rv9soRzY/j2EeKw02ku
UA7Pes0qYLPjhss+yyfWoGBLqfOioR4rEjEwPe/MYc3Kn7Gw13kGsdKaZjfqAnutnO5znhTGTo+9
+uYmugL69xecMWW/E2Sm3PIcujengZCN0wEwu9r1XhervZDvl+FNeVMu4l7In2QZ5ce7N9+KdHv4
wrtkhbXgfV4vt6VIP1nWnZYjo0DJkPnyb07glS2Ye3hEbzeQKxnbTbzooC+mOgM8Kgb/fy5kcS/7
pd+RbSLKxk/7TCqtfoRl2hRWQ4QyrU/z2P4JoMsADzd5S3TMNm3wXaK9CK5jfhWAjmffPk+0BbWA
ODWFwWWC1ywqBPMk00CNt/ygH+ehFhcqbOrs5xFMHh8x93wYLV0G/QPdBBcUXWTOZGWTCQ1FVIPg
gFDX7d/n/BK9lUYoNchvm23pEvEpiqufIG6UKukEiLlKnSgaKjCHbxZqzoMz/2sCUvVHpNRFtRIG
+Rov0ViApzwlrqVTZn/sbGN4Jn8gtX3i5kG4GpxZwXhZd9Wlx1vMsZZ12RVnaHHD2JcwDRuyHK1V
djVw8Fm5gdMq67O9azP8XLDJAlVFb+KFq9TY60XuRSyrIfQnpbFcuMJKHaUnEng457KYlQtD36vM
FwcMUcAIs2vrF5Se8a9ZBTpAivHmvqMIReanA6K4NNMXqnoHjZL1suvdJ43FBHGcFk9w1x+h6Da8
xzUgCUVzFK6zXh6C646P
`protect end_protected

