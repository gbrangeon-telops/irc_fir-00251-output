

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
ZF7Gp+JQYN4x6Hvjz/p/glt8+Yhfw+y+NSJwSgFAT75FGfBEoCi9gxGC1aPKEYH1nKSH9HDVBmjN
jVYDQh69UA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
bCrwACZO6VlyUjDp7F6NflPANkTfGVm4hgH/4AFvgK6LtR4U73r1HOWXfaKa3y3uaefm3opyWNhK
nV2TI2PpMLr9LswzFSOsgRzHCqR+XBS+8LwZ+lBVN3PhbED4ykAJBbHjWQapS4mEVXs8Bors5GDK
A5lW6VBcepABjdMHcOc=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
sWMXC7ertaTFiCso7MQnbVyuVSvzDQRw1zbA8jCBUoJcGFv+Da5uM/ZInIx2vKnorpctjF+RfQ/I
vLvHJ4hFA7ai3KLDBa+osiqXeR3vvyAO0dNGGmO7GQ1dYRUzzSKKrGTJhKWqDfnAsYaLroy6U3UI
uNSRIQtxv1ciGPzcMfrykPy27NH2CEGiCobfxP5HXDyrOVBqWAZuLaPzQRv0D8Ie2O70SiCDKawR
vbedGBup6qqgOpbOuoCX/zcbW+qJ2FxQY5Zrju+0WyLSf0XnZd4src68n6rXZlziL4eo4Q6lUGQv
gUEyqpp9Wiyw0QLmYTxtAKnwwMsfY/jCo5ZFSQ==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
d4cZTzaonF13oHTIDZgb2oXxuKQXQmTrHOYXqYqbAU6BYAx+7y9fxq+NNlLqPYeukSU316ZJ2R63
uH6wrMfXFW1V94ov6Pl2EeLSPre3P4xtwdLCKbJrudZD4i07Cl6ICwNSN//h6MJD/kwUIU4k7zeP
ni9WJs+GmLVsVx0bOck=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
W5Ic6b6KWpsR2htHXte3+6CjlmHZcuEa6WOajuu7k286E/JIlKxSU0tNrXH7rL8k7QTBc55tiAC2
sT6Jtn2FOqn9b4N96SwTUIbdNrh5Ew/7EjwCsd26VOwpEgD86kAwm7rEEtRCtStJR4p0yrbCQjf+
9+YuvQ3Ab1Y5fgtY5ijqZPgs+knlZZFAxm+NI7o8f97lEMTpHDonVgfj/KtK8xhV46JSrDB2FPhp
PMezRFDPcrnrGio0JnUe1oPbSneaSJZPAFIoGiaaxfjjDJIOa0DMtbVjecaL42P3+sAmOk0R5Mfk
8MlmwedAmXWwr0D9NdqrNJ68Zt9aVa7CXXiS/Q==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 7632)
`protect data_block
7JrnaSUqLTEpIWz2ebtJQV1+A3BdqVx/+VOrMjpRmBby/1YHUZKKZ//Zxq+yq2NC2oF92fu1rjt8
enOXX9FVEB0EUBaCsvR4k/pJjJkCp7XWdW5oMb1c7T5mHiNd579ZO21yS1tEmT5lve9QQNbOfyo0
Yce7LqhZLc/F85YWg5EJEhpJmX855F/6ygsbTID4oNtE/7t3D00pI1vo3QUpemiilgFahacqGDfZ
Ua8Yxow3MSGMGXkpOhmuuWoY5vl69oKlp8slZKGDeOtHUaOhd1FCyy5HsLzg6DDhqLHFvww36olo
NJdWcgf4eaekCRMmG/aFkm8+CrnE0YhQt9MWg2NZwBqSDly5x+kl6BGhwgiG5E7ALApGkMnPDXd6
/1QhplPxtX0/1scorOQG5GmdkQoNShWPvvAtr9+6tQHFEL51hMzTilLXg6Hx0eiR6kSKWQcmgihX
6yscmzXv1MbpVE2d5KoirI34ICMNU32Tivn7+v1b9Cl/uvUDuLAAVWuzi2ggTX/5VUIX1YSrdz7R
3KULYUY7K5ScJXEXwGXr7rtzs4doeOJQqQj3ca+SpgYGTHFpBGNQ2WNGotynlPK73F2CdAwfBIJ/
EaTI3y/JgfpWrgP5u5OBrwzY0LjiWyBDXvk36PgXXqQqT1aHegLPp7c6TlO6AhhqPn8hk29Su7x1
yK3/S0nHnnKGBx0KeJyXBcKPzFuoZRAko3bFJpumF2RyKu+//KN3UxmXenzY1HAZmjTvndOqYzYS
u1QReZJogYsjl/jy/CPuA41C4tHwdLY45aFQtO9Rsv5Fg9PC/zIWI87rRMcmM9fWgOg6hdZG4IxB
vi1h4cO0HvV4sd9F1laef3HzIjuTxg/vbiegNejJNLGj4QnR333zFYnWqt95TKPzUuepaoQ9T9Th
h7iUUJhqhvCCXKX0CX/dtsirT8ncvREUfpWKDeA8mZXt+ZIBjjx5NgMUYsAyBQREIfy+phk7Q+zr
db9kARKrWzILniPlqGi1Vc6bqvB8C8Zlivi44vqvnnry8fQma/p+6FbzTFLN54gV2IP7GICMFD6+
TI15lDq90ntCYSdLpByHP9x9HclMAW3J5hYktIvkSzsuJXVB0HZzLMtgRiwqBJj6tZF842Ffkmh4
PV080vO/vRikipxZl+/1Ur7/QcdL8QlTNoJiuGo6NZclZqiuY+v7Ypqcr7BCXxDfg/8NFWO+alV5
w6cu6GZzUoJTzIaTXetkGDQRrLl53/uh8zWcrjhFx0dLo6fuDz/j6e9qCN7IoqyMJi7W+3Gxgzic
mvRcVCgQOnfeWcw+w22CHW8I4O/AyMQdNRQ1OyRooMJSc5RxFzo3+IGMHMInUGMXHGeJTCspo7Xk
jLr5Sg7G6PRatfHSH78P7KNbAz0CXeSPGsbP8CrUfI5dx0BEcEj1AvfiEgd+VOG72kO//pWUCeof
dijfLQwEQjqBC5Q8GXqatG7rB1w5OGrRAbKp7LHPh0nyt1IRkfnEVZ04+yqjmFUEQU5B2HoYJgjQ
g531cS5baFXXtz6Ajn1J/9jsdG/rDC2ArAS8p9pLp0kgS2uk/geltPwHwR+YTmxI1ShKWKvaOVJo
5DwE2+eCz2V594pmAo2VEKZ9H2ix6ynEHTML5EYpRHTMC5dFOBHKt8iuvvh955S1N/IYHZlukZqF
oG2zcnxWA7uZU57h/kN4JZaYaTGjQXyMZ3mIb69LLS8nhVeMeA85atRNHkQZVw6CYL/4Wg7lOFQv
I/mvCfyf1Yc8zwxE/AyM1IQ0NN4QZfpUcD6D26423bKT6lOaz5HwKYAJMe2pFA61P66Dz1nSR7DG
1tMoT2u1EXH75uXkput3I/iPgObnZR2ajaPeCy7WJvGjgVCbkTP2udV+q+dFY+yX4dVmkHxkJXjW
fy5NyFjiux4EviVyXSXh0oJwXfM+LPIcAwk5Or7E3y4gbjcYNuuR9bGraG6wpg0MVt7GVr3cfBeq
RCiOQODwKK9x9FwUDrW3rK/QdRJClPyEJdj8qPHxhJyhxQ+BrIfPt1163SrC8Nb1WlBeX5bDq0z0
CD5PNy3esstIG24P5QUOsFRNH1SzWK8CSWLtAaypcrPUHJUEydOin4zjSKRVvLmsP8Jvhz4sui+T
OOHXbucl+we6lWX8+gw6MsWuMqPkrpkgd7/djbpRxC4In/1epuDrqUr7pqN+YE8MbFOGdS/1B5ZY
iTZn/cyxca3aSu3wueByYfB8eOVbybwdgUX4npHPvhDdSkorCvdOWvREwqWuymgpZwJ0iYRm90gB
/sK7hBglUxwUhavQOKWwUbr5iLq3W8i2oWfhZ2/uvSEkzRdIFeaT9W7Tj2aUGCjIRC/EGbJWA4+l
eet6geqH0KifY3kkSW1rdZWz/RkNXNQoS6rV0oZ60mKLnaQArku929agrLmDDHsOJWjbD3oJqUl4
fMmsZ9tHzbHVul5IKO/55wykZIOG9hTzogo0XcSjIv5CBRhPEawEJy7o8lcDkSJW3U+3tSVProjf
5sMXYT5JtrMtNaVRaGL4S++hzn+IDsaIjQJZBHOjpG3GrNUSublGJpJjzRfXUk2KkuQh7TxQR5Co
NE22J+KPEEMzCBaPyBGM5xtuRuHHB7FMcTJKVFBEt8CGVcwCXLS+CFMf834flvllvIhHmAivf2ed
P74ciHTWaEC5mghj3eIrCi3cuA9t3zp1QYzah3Hf4n4fvzXpEWhVDkGIwD6RM6nT9oJsmzeeAOf6
Qje/3tDs5/JKcJaQu5Rr8zdV6F4Yex1rYBVtI/UIrvJN2IlhyotsAiHe2v5Cg3YME83fjf3OlbtZ
9gmvxt5AQkNHdeGLUbFvvfgyqzoUw+H+iJ8lQ5aZCpgZxj2bwxnds8WVTxMShGFb8UrErXQwpQfR
MbNFwpDA83PFcj3lUcu6Ud+NDMPE7LSMkNhUV1a93kol/13BEUYqBPwvZY5Dsf4cdk1Bijmj29BO
JssoHkDQizpYHz0lTaWkRW0tDPvFQ9Bh0gQvBvu8mNWXDmdpnzsXQxWRe29EjvzoIecznBBSv07C
/80pY6SeT8KxqY6ikgx22NJoE+cF7PVtkrGazrQYCkWK18T6+Qn4r4ZZrAlrdEsjxGhNURYqOE8A
8zFwVE/5Cuq4kA5VV0NVxOVqNId1yiLUKlw+cQXYxdS9sdyzrXFZwUGiJiR6pDryxEpzxIuuARqm
bQNetC3nLlmhHGaL50bpnHHfDGdLKObZH5TAnG0R9IsI7A3NYEJLTfW3k8wN+zH0cbIgtiI12igT
cvn2qvZ7zY2jJOKgYKXODh18CUx52fl0wbPlGifClI/hJddC5DvO5RE1hx7RlpCRpRuDq/koikV1
0RWEvK2St5Q/AHDlOj1NHkHZ/LcnYC5LexEsonsvQsx/D0VdawnJCzKssbcl/bNZhgMQrOAJwcPD
hZGKGSLkY27e1rcmvn7A7BbtrhhiZb+ZlWou1XqdL5dogI+F039wgwnP7tMXOx1YJOvXZAChgWaX
4fX/1ByGGJ8WCgySY4j5QafwDi7SzlQp310UZiX6yMMBtObrE2+sKNQBCUTN0ymYb3jZfB4Z/CHI
cLy++hRjEOINH1TxQrCAmmQSBbROrdJVQyVb3cfyJWAoVHGDCB5USNh0XJfNxieQdvTLaJ/09R5q
wkIxxt0sWa6ukMz079hWGy50gUGIDJzdQWna8RhqbZ+L9dSRNnWSNVlY36RlU+fuFYH7RBGfrwEo
3KiFxDidQJ3sWgN91mMC5AFjbP9d8cSRFXdMOy168te57ydeE0k+gDefIZyhfehR9SsbvjXhpDfx
Dvx9cE+PdJs7k1NoZz5ZBfOJswRuKH+/W8DvfShcZo5oUyTtHuH8DuQG5i/UwgAJhNpQ1lqUjFos
VXTC3nn+0cjGvSorh7BiWaxsk3yR9w9A5NqJrkwU2+xss4eVn0cyrBtV3Vi26SCQbJbyuXYN6nEB
KgZ3qikrNKeQ9lERkvbA/VgyJ1ErcZ14KR8etJmK/Amf2csM3B3EWqFnIVOThzklWN09qv3D3JuC
aqcegcaHAHdvGTg0XUzCoG10UzvAkqV9RfuqcCMGYHHUCmIIUNu4qqZdIeEsNQ8u8x2VgEcXp5Ei
au2xZ01iYi4wrtpkNqVG2P32y8HMYspBZMRAa3iy7g8eHxAYxqgqoo1yIzQyxx8Zdhp0mFXEbJCR
YJqP0VdS5Ez16njkhEQp5CXVhRS29l1RdcV32okzCPxcssIwPzdKq9JkPkxqRUi+FwDKEyfLo0Ir
r0g7EB/GAZyKf5a/jHXWK1M+t29tOIc2WtM6w/Z5TktH2w6e14yS7qvC9jsDuL356OcNSPYjLU9m
k4nRLIOsnQStu+CiXs0Cf1GwiE6hsE79aXURob1GLw/lpzR/t/ce/NK9X2kkS/TlpN0M5CcjoI8U
04wUSfoKkoUUkQbRF3bcMgZGWI0MKxRCu3kB2We7mk30rwXT+heEvmnG0axeEYnKfqerxXJ3+0Aj
G4RYM4YI0Xb5w2SRc9UUfU96hgxuhFltNrQk3cNftI6BfC03KPYm7TjOmjXVP0RvS7onp2LB5y/p
gF0+yDr0OsV8MARlwZ1YPvaytr1Rf1+nBaBbsWX5owuze7ayS8N6OS0wku8WDkTi5AUCNucM1e8+
Lz9QaWO0Ug5x0nmS7VhALXjqOlK2tv63UKykyUWt7xPTbfbTfO13qhcsrqALXnRor7I6atkwHc3Y
Lz/P0Uxdo8rRK27pEc2PhNUmJJsVFAFCIGTd0rNu+4p9wdOUfgVnZWzqyXJHvqAAqj009fjaHixs
M8mSWrGvvCAOrDecrGIb3kWtsCGBQUjiVQO/lBWddO/wq7coCLDBmFukG5dyPhPpygn/qBBtRymc
Fyndhuc/BW1HF+WUeTRJYwDltX19g5qtdhoY5KpTN6N42db99VT1lv+/+3wfFsE3WRy04JSo3hDK
tV6LvaFrPu9tiipsdbAhQrAvMC2r8SmaPR/tg84jOgBDoCeJubgRcU1mbKZ4qmeTej/99Gh1o/bb
ZMdZbxQMQS9zEJvJSofda36mBQM5lcZi36ku3SCyGWG4SPGe9djWHp3jz+cGwFG8fGZz5hMeYf8I
/71U4ryQvTlIKGgui7J19YMqEO14j/zEacUpE+wzSmT6ComAh/k8Q2zLkp/P/56vAoMg0RLW77Gx
WoKWffLqtT6LxtxHKHLn6lvTd83A13Jxcm8G3LfNlEisfBTFduqaPBK6GtOCfu5FsCNKSjpwhQBA
0P/AtYCUtQEL++PClYULde6ubREM4FDgfw6LK5/oDkBlqNajiAZaTI85g+XxYNaV5joGk/EHHAO1
bUuv9GlucQ7oA/aiWzkr5JdRuHw4M5zj7FK8tsZMrFBlJ8z19lS8UwMcMqQKGdBNmTPaP96JGsqx
lctAhPU6MYJTo4ilMMNxcSkV1IPW4gXg8kHPSMfjfL9Wh05a+ERZ2VPTUdp2w1UQV19orWZOczUB
fy2xGZyHka4e3vrGWiZnbbxPt36Nz9uQtmzoI8868o5hgqkLeIjYlj9i/zGhaR263JVkYvgey+Ie
UdpbLxd55gknG8XI+44qeJrnxBc/FStEZKSuUQMfcfdj2NQlVAesmSSDDe0ZMqmAgEbaF4jVbDQJ
cdh7g0G7gmdYRM/5tYVLhcPmg2S/n5cXs8ZJLFM9ZdKcqfpFvG+0KcDaXaHoiuEYYRCnbM+dMxlO
yAEpQWs67cSGUxouamDdyVfv0BVXdeDzURoJY+WSlV5WXD9qimSkxMFpNM6gLZfHlRHU2FqPTKWU
kLp2ppg5Foc+YgZ0do/bDe4hUB6CG3UIm/Otj0hW7r5thlJPutYHnlnExStsMlLNxRh8tNg5rZEh
vaEO9J2hL6Fptj7RAzjfpV+Vp3D0kGfWFeEE0sNmE4ADfHefUnD4tt0Aeo2HsyrzP87cAWwpQBde
iDSv8Ym65LS1+6qNBTaAOwz0ZeHP8MAa5XP/AEn4lxUsdexQDEjTxDpgc7CDpTiI8pGdr3yMHf9+
9sAP5mmZVtqcM1c8K9WCyItmpYlE7MOHA5qxyG25B4PnEKzhiIJoZ5z8rtnDEAQ+gMRW5tDTI9hc
OceXiWIMR4BzbUujrRVupEwFcdEQEp+CHbU8gO2yyFm4KaR3JqFhNPg0mQEKFu4Foi0JxRSZFsQf
TDMgJ6EycqIHqFQNwMnHsumSTg8Sz/bOiqytgZBTpnicX48FBVbylIhgfEzYDbOiSgMi7Jeffz/C
V9dHODXEx+KvPeKbnzNaBBBs0BZWuLXBwbG/z/CqVvPa+IJlgpK02KqkOiGMse9w1V5EG2KcR6RF
n15DLcBmX6yhNGLEmL+jWMHRy/bzxiMXly1gqXg8y8WWlzIJ/NAIBjIYD7tCkYLOBmTcqx3Itowv
0G3d/GhJlWUYOhL3TNbgq4D1Dpopk16X8jgnHtG0u3R7HDotagH5aybGK4PY7Jl0Z0+rr6AJ3Vnx
FJXu34cGmQpdstG5bPd0XYnocLsMKhzS6OlMSnYMFjvXeLZwl+ye1tTRYtZYPLnuc5/may2EiUPp
s9UpizAgxqlYaR/kDc1hymAZ6kB+tBlO4yc2yAuymPP5QSIXpX4iX08QWYMrUroUARYOHUQQicTg
CzuBLaooKYQi3b8y8+75ApQS0NUb+jtND26atu3z3X5pKbgdEHwVnimmBNC0tg7UgOZy5KSNTRkM
sUJsq9QoKrdJLt4U/+x5sJ82rgK1A8fbJQxFOo9kL/joVumasW8YKE7FpXBlkVlpnHXuJF1KOZE8
7YW6WBL9m5QPgBqb14Viu/sTYgpEZXBEeIJPhxtE6TTmEW7gsC3wzDRn3qu/Gl4z0YnqsYy3b+V2
IWUrObtrVkXLGMAwb01DEWcPbnU6miGYTXJjJ/F1mt3rtH82UBIDhqwW6Zl/XOszE25DxWh4p3k/
H4A7sSwsRsqDYcAfQ2xQseDEMV3+JVQiamI4gsWrP3fCh/hfxgOVG3JnZ0QyYlZ4f6brWGouyYs4
YDW8N/wl79EVKmBBjUDdJmuyrs2Ls+We0l1D/IouDS6fx6r+89YM6CDv+kgDmpPN58taYVCZ0MP8
mtYtyvRv/4rfEYz81KreZzV5mcLxFH9rdLIMLF7v5TQXcASdAfua4COH1hfuYRQNKxE4uD215Nix
IratoBfnpZwIucMR3Tbcsq18sRn1kx7954Da/GU/dbj0CM/7nadapWC68xhjgQYBuVXRSJ6+MV+l
zVS4hdHHyPos+C3iwPObedhOYV+jvTc2ZbqGRDZkzjUgO+JShcoNXLo28Mx9t5dHUm+Bx75VDeZC
RO1F1STdLy7kQTB35/FlYaIi0kI5mXiIaX9wqd+draTUDMdJIo9EeGwTqXTVwUoslgdpBOIYHmcb
0iEAmBHHEXSow5c+1ipWFe6uv/yDdxUVWpPdKj3kkJbQ4wAm+1AwLeWqBQWAFSNNp5DBr4MOuzIC
z4nkt3Gj7CB7JRWOBTSKD+te7BWNKCFGkumkzPG0imjdW234DUW0ucc7SvKRDPAoSxNQYUffYsfp
PhrgL+BJHgUNMYVE1F/inrc5MAo9L8iu5nftq9lYh4zF75cJC+Nv2tW1GVpyOZVy+0YCR/vlk1Ln
8f8rN86j9dS0oliPuB3wgZKt33I/73dQXviOWP+qfTQrEyIGEeZAABCG8JD0TvE8vrt15TSaZrdF
prxPZY82wWJlK1ghsLR7Rh8Suqa7V8GB9MgOTi9gPImIIfZV2qrV2rprLh1wcf1fCPWOuEXIVqdf
IiKBbaghoNGX9dEb2dnoQ28u/zb6YU5gw0tpnv0wVfFvBK5qCnr26+zCKgY9vc0kjxGRi+hS0EqP
KE70I6O+96zM9jIjTQs76U09sXAccVqJaP4i4gW4TWGHQlw5cHuqDtLGl0Ule5jzusqJNHZHEyLR
iJQRRAbvSLIAtgaOvhp76ArXQuXmsztxwCEXSWZGSi457y2RhPCW6fEoYr7vpXyO0B29WIa3+yi7
B+402tkThswUxocjANlEEV8P0zwfOpAdhTfWWgC6296DEnkpX7gm/aNOmqqZJVWzn0Gepfp4hQ/b
5KI5rLAUEx1bSvqm+AEEbUr0azLm8YW93IcqaKLlkzE7pDxLHzNH4gtOx8oTph2Z5z7zw7Ani8/K
MAganbwoPH2eIWpe5inKACHUjpGVh9t+zVAPVc7ym7A9xGZI2qnTOSplColhiIKJNkvJm32ywVsj
+ZmppOL3WL7CHKs+B1nlz7XRgXtcTmVeyEbb1WqeftZp3ZZ3ZHqzUBMT4toTyqAXbOp+7ilps2GZ
+BKssnZkYN4jq1AdAEwfwe0LDAExStaaoTDzQp8kJm6AL5U4FGpXYcr9lsXaKFcG6MQE0PgP/aWg
sqktPgaPk7IpEPA4k1Mi4WKPbeF8ff3Ds06/hKYYnbPkVUu7UXuEhP0nZrXU9qgJHKI/eQJW2m79
M6pm3XpoTeN41jHOGY8enCbRR8oFMpq+A85kqU5hym3nfHYTl0uIm7j5w2bTFL+UjyjDH5Y34IiQ
KTSiP28MT5UZ6SmpIWI4Wcek7j4C7UpZtLmxNVHZ8QSKUMDXk0IFE8lQNfF97ySalJN202YAFmSb
ZU07t7gg/H28AOiu5Ls6J7R/gtDJvXapSicdW3SkUlT9TUBYi370XvlHfjFnWFFig8x18a5QakHc
jBGiCE4XoaqtulOkaVsXC9y5UiFfFGKDtZT9PjAnpK9rzojTQRb5abaK85KyOEWGwoj5YS/QaVFu
rR/cNKRPtCVFZYyw2eJj8hEbzC83Ref9rOd1/5tOOUA3nMUYlLT3SspZ0a6yAzyjFWUTFGmG/o9Z
yMX6xHDfFQVa/5QNR4831mnMU+eLmTbx2gUb3CUppoWkykASRq3YLCTQCC4epzhlQAQX0n9ApX1j
B/gobDfFGAPv9hSG13THMm0YDUo+0r+zTWs2z2zgM4SIskmrI4yJsha/4ug9sEh3unA4KryMXuGF
n11Fa4bMpv4leoxvIU3mTdqXZBYxfWLiDO4sy2X4SCkxncrLTeTpOPSHZ3Qt9c6HdB7m/h2A8NpG
6xCPWXT5YAzjPa0MXPWCR3hAaLyBcOP69NfFe3ng6eL+VOkDA26BBdTxlQAcv9/T9lqtvjStHI9G
03RGk2Ln4eoaS6rEOBkcu+wYhpS2OSDjLafdPddynb4IIGQONZs5QFWj6vPisNBY9bCQBgWwUWs6
cTRw/RYIdwtZh7Rnls9L+TTBDeSKGin0N23DhMNb8htITlTmzlmy+kd2EQBoTCXaY66qJS3SRaq6
dUe4fDaPRHE75h2/90PkK3zorpnY20GekCc0SZMVEckv1d8dKUIydPiOy5vuW8z2h31HZB7KZFcq
37DqGOMUFtTzfoID83D8x7WsdDXXYYNSR33CYWLdD/th4PQAOeL6xxs/dPEXAf+fkItX9V826EDq
rodfo5KsJLXIqXA9pFgY88JP4rA2h6n5ALIQyN+eXH2XRmyzR3OJSoxQLGxZn4eUqwQR7gv/2jbb
3vcH9Dmd7qVYaX18LzCIfUI10h1gOC+Cb1nq2N4C59/L7K+PbBzg5SApc4dAD4sX2H8ZVIX7z2l9
k/js7hZFgdkndpaB8lwd5yrZC2gU3Eyzee12Tig3xkTI5AKfhCx+9UKuGTvXJA5jTKIythO771YG
/WfOfM16U7R5Zczf270pjhzVhhYfIXUABd1JB1GJ4Kvzyh0g+cgueNme30OU2aLpuPZydJhHA3Bh
xWrdTzr90FilUckw69w+FH0WrBhaXXwiMZurAcmi+QH8vdZakeFhttKJPgwWeDxEvGNOH+50n0+r
+PUsv8DRwOTS0iro/FOrijh7gxBh8v754xwWiL80hD7SMm2feS4P2ilhu0gkbmDO06IfXcwQw0hR
jVq99LIFGSHSF2SMWXcW3M9xVCzgIAKmC5gtOVL/Qr0Mr5/HTcR59zdeQ91951fgsNsLzdImzvb5
RCyIxUUKc8C8XpKCORaXG80F6JzLXx613Jdt8m3fspnHTR92VEXXKJyTN/drmpINdhyB3umDXgj3
HgmPtX4VtY4NghLueemV7JNhc5crlMKrkgAZ1DkIQIRCCjHcYXgRafUxPOqzNFo34jCh6Ikfqkxf
yVS0vAs4UYxuPZmlxl4fve6U/RM5kWWYDRuqNgFnJGGzn4S0l4R/vVCdxLk+q4QNMMtm
`protect end_protected

