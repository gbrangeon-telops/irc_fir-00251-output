

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
FAkw7gRmEwDx0cT0lLfFXgH94E+u7pXWs5ahSt/pzljIAtlVd5PhOu9ztNGUELVfoO4Gol+zPLUh
TN9yRctY4Q==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
OsI56UKE4Z4O4++RpLw+Gr7y1Sd3eUkdDGmGZYBu0aWjoj+iDwzKGBcBG0rF5D+4LwCAgnpAGiys
xLyYTz/ObATK7L0zNe+Mx/H+/j5j5SXpNvpcXkGCWx3Mtg6EpqxneRyrD34svh6fn9QBg9AkFvdb
eTcam3dZU+Gacfm2Ivg=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
qc1VB803xD7sVBXVT5KuCy+daGAjeSNtMgViDKH2bpJoW4aexvjdVOFa9Cn3ZQUudsfzbRtbOfND
3qwRkfwGKGa/rWJp/b4u168LG7R497q3mKgxz4wZrw5VVWth06zATVCPkvVwwcP1aVCYV0wxe3+F
BcZo/LoE5dzRftELWM1hbxUlZMlSl/apI9c5DLD1ZPtssPXqyfH8yGBCJ6IwpqThHkCcKlxPWOFY
XBErOYYrcO+fou4DBovYWIgQB0ZKOhCR4cvN3q6rg5XOYT99xP70Y8jdZqXKRq3PuDDZEya4uwav
9zgp9xA7sRjUN5/fcIvFMcfDutvNPIc7IvkzWQ==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
xeydwtnivo2IBZhciZFfy3r1qoKk43zuwlyfDAWr7E6QmSwqVQF5VHmc7oNu8/L6oqsi8CW2guof
n3LQZ6J8fPLN7CBNStOEImWoOU09vnECk8Bwe5gJEo2CSwnqojJJlM/jtH5jKtWnMb5YecjpsAkT
3bnS2U0oIgAvNLFItdk=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
QglgmN/aSMz0M17AlWb9oRKStkdBh5nVOwe4/WnjlbCHuTNXWcMIzqLlv5JcAmIdzL/13EAMS4W+
LbXaFXFMcWHAzC/5AZxX+CZbwE46qfB6uGUmUBTFEckk+Ba1aO38uKX6EDual9TqDkiz6OPrjmC5
MifvdDzh7mlaB+rYqb5sjxUWUfJCpXIOgO6lavL3535AS2e2hAYpmi1PB/ejGTuva2r1NRmDkiUk
Uq0oiyBI4sQwmU7gFF9pADJRyzpgRQuSICfI5NAGRTR3by64/5TeOArBdjuY9arezL4gMGXoOIu4
E5vrAQOLZikLF7X3/wpaihrUarYdJnuPPVXNaA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 48992)
`protect data_block
NgaDwLYX6F9Qw+D+gyBMQFEDLnwdvGSaFeFOc0LiRHbPoWS1zIRueYgypyYgFTBM678JSf5MRCIq
8pHomI9UpT4TueK6pfZjxBsuesMf0dFInov5UdJUWOQlPPFEXZGaVwE8LAkcd2t83SgNiGAQ+WIm
hLzO5Mjg5QgFsRZAN1EWiOvGcqQRT8BQY3yeArUEkmwRvIcnqaS9/CoMVklgWS7YlNzZqILayqoS
z7TrVem0+li9/RoVIS0ehPzLqwZI8agMSj0sFPLlejyH6dZgMls012CjZaB+Z2bop/C/ikPzJkPa
HpAQOTTLJO1/dQjeQytSUm6/qdcPU4LWAyWSuS1UAIxugqvnR1cHsq6azqvBZkQ3KdCInrgopVVy
ut3noYsB3dXcDXGRV2Z2+x3dyo6LgjMvaIRvwcOXRW9mjqTbUdaHNz4m9E3PkNyCPRn17Q2gerAC
DLuuI+VwoKcp1gdH1y7j//E0MF+mwPplIbHDF0F5m84HywyJDaWinpYf8vnZu3BvZfoeNW12FFOv
JQvjoMqI1i5q/1XYajlcJgYXacmdP/3KV0q9MKDGICqm13kJhy9Q9QqppaF044ygt2LNiKl/1YLr
kVYDMx7VvFh/dqgt18ICBglLfnX6XQDlgn+pRnMDHUNiPj7oxRWlBgwaSwRyE4sZGD2kbuLbB5EE
0tbGnHRv+fFFDW4wSuCzC4Na8G+AyCJFUH35It7BdIaCsxxxt7Ts+30TzTCX/Vhn/bdY3U1abH2d
ArIGk7/bX/Zid+WEeCZCTqrisagcS+knq3GSS4V+JMj5hjuJpE8wznLDUtcxMYBlrRffxnprGD6f
OXNSzVRGVQE9lEUwR81G2zfTUfHCVwZox/gd5lkyGi0YSAp88gm8Cac6YFe2KEkQMpnu1G/ImgOD
JEQQGcigSKpXPt4csGvKLxAvrNfHVYm1dAqpGdirc34LYQTVL4VXVjf2YLC/MNb00Lumw32czL1w
+a4bAgbh4MrXOVi1rRR8XCZ++ofWeC/AXHrpAzjFvvbzgNSZ7pmOm6SovVvBg2Q0+xCDp1AIAnQb
blKff4n0/zmc6nAA3KJQDDiJFLViu+HxiF7vii3j3HzYa01vSCB9Ga9p+5hexDfAvX24Ke7NYOhf
0x+663NNnrJtVEOEDPnN4wZDt/Roz7xHs027eu/mhya/O6qyqZTLD6AwjzaEfd2zhjTfjcZ8TV2n
PSsNtwnPDigPcLAxW22anKzYWFWg2KWE8SXi2uDLkpwocnqYb600Ck7zRgiY56aZRQY1djUgILfr
Ykvi5OzNI3BUeSGOoDhjnnI+4UocEekzBvYz+YwLz9gGB29sDiaFYtMwP2rZWlLJ6js5ouBwhpxW
PpcwmB86HYxLaJUYMQvvPcdp16LKKpF2yIsJ2wJVAgG+4EeQK0vum/9A2Yv7/f6m/vbSTSsjaH9B
nm91fhBUX4OvxP5S3friEAklRm7kF3CjnoKKrk62f5DUaCzlysMhilzC5vVlhNxPJ9gyT8W0jMrK
LSs00G+a4PnArY0pQDR4JChvg8SunTsdVXxZdm62kvZGKb7XRYuO87XcFzW9CCPQ1oOUNjMhRKoV
nKqnL3IspFAyEiljYJow3LbhROCKTm91Vbm4k7lTvQ3cByymvvC1AJIJ8Qds/5D41uq1zBqNX29I
z7LIJ1JPCQ+HexgdYzM2Bxcm8tEo00MgcONa9eqtn6pKuhGxqZcHfJRuqyLA5XRSrXUwHsVGdyiS
tJ1gs+F8sjBGVGr9ndp4yCzBxYSkWbTeqt4JfMC1zS6fSfIFvNcheAyElcGbd+WQZ6+OEeveQKC/
QJG3otM7NwHKR4McGIVHGi31i7vtvCJgqMqCBDL/RLJXMZ8dX5XEky34C/zGvv1M1ZQRavK0p67M
ecoYcXWOZPKl6DI8w6As1Jw5idPJuGxPcyM+HA1uSQEEuHjSrMZ98dJu0EaysFsxKFuRwSvetFcW
Scmtg9VTZhYOirOGNgKKLAiwiXA9xyNEoMjNxvSNr+iWnBWpSrz5CYDua+u+zIiLUfoEkCKmZvIN
iyhkQjACnfBED8dbKy/TBFWDXltvwBQvOYveZa1n7i1hTVyaiG1kQSrSSMESlvy8vmXAu/HVdrfu
OyugvZZTNVVMpEtKAM0CcSZSNMIu142B0FLfAI4TZYW7pYvzysBdYEQSdi20LgfrTGJQQXlx+inb
Ykncm3Baa8YtaX6vmUM2tLfRfBcwyFfytRJqwxl8P08chl9eb21J7u6OYJ1SQ/Bz8eKqlAW9hygz
mhEFaywrczfUSDpubj1s5+FwUkoSNh47AgtzYXtN+MCyN/QtmkCSSF0wAQpBUVL3xYmuPmwpT34B
vlhGwkJ7LYJ5glM0UOxP0n0fQy9vyMX6iURcOv2mhCi4u3eGwnhPE1j+KAva4ZBBYR93v2w67nPP
KDMM05mAKFYBAHnJjdbKodNSKOvQI3VpTgQcwhCCrQFKFZ0r3XY8jXsi7C+2Sj16LWjSVz/UY2VJ
F4QSVik9xiLvmvcZ5mUrcHc10P1R61329ANJd+UzukcBEQ022qQOIt7PdU3laHzGcidgSQqVs9Qx
2TyME9UnmyaqdgftlY+A20iDa7Rrzuo9z+9pOQtshBwx9McTtGVAmtUi3lnYmJuqRmZ5Rtpb3ZZu
WLJlKm9VoZv2fdxHoZSNN0eZBoySAgH1V+dyD3EtamD6qkknTkp0B5HZw9NBYKfV/Cg6CKfQ5lgS
azI+o+3LVmFKyhZiQeBqdzfLtLlPRlRYNDq5fz5rjJKXDJ+j8b8FUvf4Cuz+WmTV+h2HYieqdEmo
gF4PiIw5pPzyVFn9yelZnWFhJTThmK4CcFdjUuI1Bd56IpGvVnorKRADe7T4RLF2oy8dtmmZC1A0
BpV7hjjKWIG551XqiHtx1vzFRdzJ1+6PSClt9tSDyw1+Z6po6Z3/X0hPGbZQiVAxFJeX8yygx/lM
dut45QPvQywoCTVhMb7pzmc9ogVeVcsLch28AC6r/KD9cVMzporg0vOFWAkdFJNXbnbIWduTmDdD
JottLLu8ysxQ9rtmUIdi5kHkCWfg4f2qcIjtDi7bs2ofMOCjdye7GlkZhaujbYSm/3OEhYo+nXvV
o4Ic1RAeThm62zmgVr4AHqJxUBZtg5JMQM7xHop6MboJkcfpbv4Ogx5qtM3HiUTzzBzg+vWMfMJv
fzNHaYwhFmyYcP4Y7+xT6HJ0MZNrpPhy07UJ7qAS596dHS8+8NV/AHUglpMWMQz9ke7vTQylp9Va
eG87q1jJu41Or4d0PdmWevzdfSaRiQ3lMYphfNanzP4rqcqELwW7P6mYLsMwHYRfMWZckrCIas0L
9zyqdDR4HbAdWPfQ62dsJ9QhErTrTqBOtcTy65VMkauDx1+uQY1CsqFBNXRVL6u0i7t3iPoURqly
kLXFSZ+JlygjhmFrBWD6Y+/VnvLsMOkp57S4BiDg75lS+HEYzJo0ZIHNNqijWfw6Q1d+VEBJ2iXr
97oyh16kf1LwyAHmgUhJPPoa4OkHd/51lhzXW+8Sr0VenXkDQwu1flhGVh4ZpdHxG3vnUk8EPCai
FONkHxKqYR4UMX+zi24VryKoyrJdE70TNlj4KTH1vun10ncNR+/PRXbK4JL/g5oFQf1339Sea2Nu
2YYSfpm2LH+1jTYhv+fsZdkX+p4atzttRJzrK6zKVLDrsX1fzEJe6WjC2Wpwd9Nez9RqfAraF06E
AMkZcwJVHnWyxnJsW+7b99yNV7Vm1DCB5KMKMIFUbiPIXDD966RqtK6QsRWE39G9xvEq8/gUDzqM
RYSZ4o8VM4+qJwimvZXVb0TszOR3N/IHC76ynfftWm9iAhRDqZLUM7AR/ymnqQPG5bzJvbYhMaGE
MsOFi+r/QnMMZ9QZP9t5gW6Vty7lVY21Ynbto7dDBy453F04v3v+zVzig/2UhtHXBtuh29JLeThH
ixsrK+6ptCnCRjQU9WKX1b0tB6rSBFahOgnWnGsqRx90CV72eDc9Bphr+pEK2ObcVTcN3eZH4pBA
zlrA02IoZAaYgVbBmv0Vbt5v4DozFaGYmFXrpxAyllvjXh7592ePdZrjoDn8kmUTe8O9Dd1yKjAe
gzXN4B46nqrFa4cENqV2q0J8kV1QXlwahrPLZiq72nUHF5v6M2zJlNWHc3jVnBMM0FgKG4oChnwZ
dJ5LLThDUQjKh+j/evvUyfXqBu4l5A+vXBCY2rU5W6YdYRPlmvSCB6MoJ6Bwkq5coBGUF9MwlxX6
4ssZo4GNB5McNx9lb9dusaE5Sozdl5iUUqOvGLRQL6Xv68V4aS0n3XQN/DVJDlD6SdO4UISjpVS5
JHpqUyn7kvhtxC64Y5scafgautdGDqwFbfVgg9GpS1fgPwXgE5Trl7d7S4OFTEm1gaRvy+zRNKW+
eGxfpyI1LeGCXImruNspjfisfKkO5BwDwREzA4RJY56SmtDSlbERg0CwzbSpdLEgHAS2/LOS5Xfa
MhIxXV0XoeWpZ97smEN0CLGyHa0HzfXB/bXuNgzo4/rr0kut31IHiyTs04rBHkcYM2FDvwcSKH37
Z1TIdD4GOlR6aJTzxeytLyXYavDmb8VadgTdaAcLaBC4Hnp9FIXCQrHJez32/5CHXnB8wDB2qfDQ
MH9xCuLG3mxNBhJWVX6QuCRnDp4BPEsQAKwu7K3kut4cX1s7XN+7DZhD+D9woMROQogrB4udPSZL
kPasF62I48JnfXFFaEfPvPR/qeZZPJ6c05UQIpBKv+ZLgnslgjFGXoB+Rej4oLEMUks1ov0GeGTL
CEeh3fJIx3RZR0AxnI7s33frR8ndhFjCnjAVfqqzT2sFea6V7Z9/Wi15gg5MPzdK1ARbwtY2sMYo
vozwMGkn9w0HfbeQUHNX/JiWTPFS4b6LdSUX76G5J8+cHWbyZLxqIUuJdpggcFV2pyuCshdo14W8
DmhGIpZO+gjxAtpQKTtQKICynJcqTWCvq7VZFv+S+ZStUSjvDjxgwTVl0CLlImzao7q9JO5KpBVX
PehJJldpKbGCX6ePkldlVJa4ooLzjFh3OyQwKdBcWJpV1I3jzYy6Pu3li/+f8NRJpmhPaHTEPx7V
sAeNMpULVwVuDWw1MluO9n7iNSilW8cVxCWMIBnPZ2bT7jURZoQo1uSv17hH3cNXTxYnodRTjt6h
6wmhfRoUu/K72CoPRB0S4CmO/27EQquBGbSKIPat0UgCwgu7DB9Ua17pQJTk8FAR7y7NDK84WagQ
1Puj4r+xri22m+hL6NeaV2LFW3iFnR1JDzdVn/51Xbm40K9xNKK23TrPoiiSDDNgWIsZgta1grzI
3H19cLyu7sZ+qUVFHn533vmg/JWxix7VF0cNeAwuO7relD++Jfbf1hiDHRDRknVmCZ0Ox1v3/DC1
0wqCikyFJ0MEUeUNUueM4nu1slpSnNxHkNZgMIzEMCdb9FyG7t/ladDWTpcdPf3vpsD3eFWwO4bl
pVkQTdK1XlTszAHrufUA9SfwuWKI9aYo6o4w/gQ/IvByDSyLTT1w3jprHR9lyc0HFeyGQKRDzepm
Cq6/GJdlQm1Lv3t4B6DoqihbrNxX1TBI4QgS+1PBe1pz18NY0qDxKSPvxZt4nDBU8H3xh7zIw56k
dEWCUtu1p+z1OMqTxFQnX2mFgcw0d//tHc9WW1798eJMKmSSuatVGCvIkwmilzP2rStuVknEsBvq
jDJnYL5hzcvvJJ3sfhy/kFoQOxEQdIwwArL4dYre3RSFRKXCfbCcahbR4+wjO3250qf9G4BXCBfq
m36fNwpSzPUlrCd4cduz480ezxEZ5MBd1ZdkU5NEb06yIhjQkNGdbg5i4zHelEPKRjqyDqf2ZIaD
bJ1z96fRNS52RjTWZfW5SbxsNdPfjR6cHBHFZAM7Dxw6UBZA8jCAVagAhKbY06+6w6S3W1VhQ34+
33mLaK2i3Pu36E7KMfoxLnNU/OL8E4+tf/A3tT58PZGpiLxwsu8H5lQCXFodVJ/3B/B2HT1OYpng
BvNxDWYoANzjDnvaTb1GiNnq/uTsTbKicYXCmox1RxXU/5SLce3gkp8laJdadTKekR48ZIdTWl/w
69Ycd7kmZ42CFf/Wm94s1Fi/aQGXYHb+kby9hOEiJyeREK+j7TBoGOi5fvFckFb3b84yh8JA3gaG
afP5W+mDX/o31yPUJyIKH4prQ5XZRPX5GEdm2mOHtcTJwcTvBVpfTEGdZkc8AaHVB6OTWcCZ2JcK
AG0nzG6hIbc98RoHOe3DcGCPk77PMFgWJ0NLtcel+iWrkV6Jb89eIuGRH2HyUjQbHAjaXKZ8BJww
Yks6WwALBdfO7NkKFLWIhgzWESwSPY+r0Cg+veU6pWiFzqymyFAQr05QpP6Nf3o7A0xPcjsY+9sd
uTgG450QDtc50BzqwHSmAgJ8AQ9hhSCPMT8DxiFZ+KFhF5nKuayvf/KhH6pt/58xu0kaOo7tCZQS
E4NRgBbyWYQaZpeaHOrUI/fO5GT8mc5p6WOMNQmieNl75K0eJxsq1US/ggQnbUAinyVD/8hZRxkT
yOI8WJ3vvEz+o57ZK1r7U77ufCQqvlW/ZnJNazkQBkgy3APDdEFK+993Jrn4ZYWl+YeBFDoJCwuN
uEWoL7CqH/gOmpFPyb0JDwqWkHM5Xd1S7lAcp9GOC18GuVozsUkhh68jQpA30t10mZrngzMG6O0W
LiKZgM7RZ3BaYUc6OPaHr7OHxGdtxDOFyrZX+CPvwT3gYCdEnSc2rmOaeUqFOhpFQDKUOjMfQ7cl
hQXAa1wQr1jguiDMLXd2zX6flkSb5fia84t/OaTmAMZKqWvfMVUieIUolWVWHS21skwGm5jXvicJ
g7qrIeQXHgh1QpyrU2o7v9QvuG+1eZh6Al7v3rANjI+jyhujy0tvFdfsgvhivcIDQOoSCURDBx8+
oOZSx3+V9Ydu5N9M7EJHqnErt6STgIZUYjOkdTTj+IAMoBV6D6uL816tZX5nDr4zgQBkhomUxPfn
TWuMoEfUG6KymudLCV6Yos/hGZ1Ckl0moYsQuWX3+0IOVUo2/z6E362Eg1UP31YeMHqYhpxXuAgY
SyHl3NH2HfBkP2dHhQ7CgmZ2MBpjGHsK/onr8VqsVzq6CRU984K6Z52GE0qLyKpNcT6CdKOj6GGM
x1eAb+MIiH93Wn8rB8ie4uxaXFyEUkg8NBetvRCgO2KglJ8c9civ60iFnqJkj+19RY/jzUJLKYmE
QcLcKFvdcKcroIH6YAUhKxWZc5+8vjxcbbGgqKj/m+S98Hd5BNAW6asaXFn7KujPSX7QxTWFcjJt
Wy5HskPEiCytxhAAJ9tK/am917sJXT+2s80DArBZKoFJ2xFXyPMhzt8IAMmrLvm29vMtxZ1Xfxnu
SZ1mABQps99Y3nF5LjRYAuyppLEwgQHTOhkg+bsVFiJBRBi+dE/GXZftkThUMSv0VTriy/6zrE2Y
Dt5hzS4+a6lygIPYwmtoxR4DZA0Sdxx4Q3sdsCFoThUfCf7jq9ORLEAlwsbYipyAW40zTcyRtkpw
U96tR8UrS0IQGmAnTnJ7qnbGoR3Y4RpqCDmn2pP8wE65gNpCeU9ZfBlACEWhEkS0bePJuR8GurIk
J15FmnycNC/pq0tOs07ukvlZrb8KDEYPcECUcoKCQyUerHZstpuTKdZudhlkQ9FLJmeTkC7MvWoF
spLk4vUhOjT0Cn0l7es+q8DL8YabkCnO+28U57HwA1jgIhx9fStpMlD2e5a+aAtGHpUWvLYSsRzn
W9lWJHhjzSgplQanfty7Oco0F9SsArTOC9G4glKpEV7wkWJcQfoG4fw3AiJjPz8/r3tAoZbj8w9w
ipDJfg0aL97q4reFRlaNFNjcVM0qiFsLKZ1x6GpdFUg92SPYono/A9iWgU6TnI2K67lZR7nkZF7U
q6edkuHhlYRzGv3S7Ori6rMDxjF96bReiB+WJWROzhlJHolfTOSpDsRou6TRrMUhk6qorp8OnDxm
HbypuBNa1QONfdTPjJeTM/cYuYw7heACTUvatxB3poewNuVg9jNNkc5KGzKoYaPORQzsytfddMk1
eHE4Wzm6RxdG5S/qNxq3VRYS1a3VYoYb4JvufKFM1p3ugHXyzAeItRoMWEGLG8j+/wZLk6AM53bo
Py9nrIl8G/VRHRCJCOIEfLaPe3kWSxl/Kw3zAv0IUWooBFOX1zGmRy1NUb7NN5HvIMBmRUAf/YhL
+TU/gOLX7O3dig5BZRLhxhoRSxZKejjUCW/MG6apLFwL6QFt4epQwSOhkxpJFPucbem88vis/BAE
qz1AuuYQ+2v3AC9hPJK3dapVrny9GFxIwuj/fb3Moa2Pmd1k3OSBD9crQM38c4KX5J9yUJs9NsIe
3w3cLF4/lCX0k5L/tZaSmoUZzwQFoWsDXR1H3ZLEUgxwZ+XuKAlHbrgK6sqgNJIH1HHiSW8Fzmip
9TFeFj1XrxVq5HatTRupZk8N3g93Bqbl+bxUz317k2Y/qeRIJRKPJHUzmLblsWd0EcQefRToAE4g
1KznYM7c/eE6TyzYyyUQ+Iz0/zyEOirbc6x7qr6T1P0FPoBnbt3eAzGS4cgIRoXEtLjDxNbz6giO
4MouLfr5dnhs0qMI7/pRx/eP+g64/b6fhmHRaZz9ZN9b0RjQNov9o3Sq1VpjQe74XKoJg4IjM5/j
xSOaiECJcJXK4X0IPiTBzzJqDpCLz19otWWYTAp+jKuIYT/fO0fbXiHvg6zNn/uNh9Ew4SZvbJ7o
2DYUhg6/4w5SLJt2quDlU2gRSmkoYG+N/+FDheZTbL5SKSrEbzb9NPQjtoWlYUnk2/wtb9BX8RrB
xf2dDzsDQQP3YzUwPVXLuoif2Aec/LHkcZ/FDDAzUh+0dNUbKs32puUahSOjY6n6UU3fL+vM0zx+
s/tWREDEG8BkVlEi1LOCqBaJgQnx18OF0lkE64u8WiNO8HS5hhdVeUul7YssHFoKXGtTsFq4/Xlq
Y5tur4zGhQrFZXOUi9pealeMSY0KlTSp2FAxROFs4olp0ifNOaYi4UhfwYsHbjhWZMSxCjAlcwPq
guSkuxac+jpp/nZJcUcs9MkBiPN7MBhePFTQXxSAJOX2ZgUTe/fO8ID3eB/2o7/qdbsdMMzKpyEV
qWh4FtDJmpxieDto7Ty022jY5YRV0hJURGLuPiZdfBM9wO7kEvd6Kat5vux07RPqFBHbyv6M+JoA
Ebhf+gmFa/T5Fc/0Co+iKLM1ddCS2dGmZ4n+HLKXqG2VrXM2O1Gc6j5ld96Af7706a89YXS3bnwN
POTGsqXfk7bk8kCTL8gXH2HN0JzWESv0RpbYRx8lJ8UAIXKk/FTINLF2S3VkRQ494bJZ18QGeYAH
EBrYfP7Z/6LPPQXzFDA4AxRETbxpCuQgpi3zhwZ6NVu0U4GVavvaKoNVFA3fzaE7dzoMT50HRtA+
7IadF9LsQJhO1BgKXOIyctgmEx/suDov9zM88piM/RJ0JMH1Hi0/tnbtacFHSDWcRSuJ1LPG9LOA
fsIUOyYuRR7p04bBzLhCz/v1aHd8V1VClyoXHUHlNBVw7MGFGO1ZBiTqZhHuiKG0Ja3GsuLLjw3S
NjjzTiyt4+LMCsVjahr6XxeFl/xxKnr+CiVEx6x7thdZqsar8Y+dx/uHE+emYPuJX+PM5sRsDNyB
cZmtF5R2ZH6hGNDTPhuJ8ghhXyIXO9/huj0iGkrj0j0hRJ9vl3E4jMpqvnQu2apMTq1DpyXmMHI7
XBdqSzK7dFML+VMIg3TL9BiNv3dZfHlOl3B/lgeThJHQ2pel+H0SL0xxwzbDI7l5IiXr+fzxqA1j
jV4XWMBrMOQgMpdWVvre4hG0DS2JLWfxlWUkC7SZhH/hK66gxCZqFKZTItsqjEaxAUL/TGs1kd+R
ZMmw84oyU4Wo32bDAuJx1KzI61wrV6N7wl2iRajxUwXvbs3ABz22oFELl4ZHaIJLWcEBpS9/PA8l
CohomF0dDAIXyGUn1vZ4x/aT7noEzawL+pjgOFDBRiUocJqfPgPubXoy0DoJUUuLCU0rFQWJvE4y
b0m/l0mpALlwwm95+rp8woEz57w/P33BmR/sC75mCMbSiMzaVlm3vy/wAX1ZEos+gFe0A1OqnWA7
va0mkNJgLnbwISVrthH0Uv9RWbTpwimx+Xuske8Sn1dEFEvEXTXgBi2pA8B4jBa0NvgnGy83sTX2
vKiLEF4hlsHehJ3EokN4ZcQk5EL1wb3z4vCyGf8NVczN8Ur94M3y3WPufyKD5WcWrib1dTlG1ijC
xhVDmjGd3M423O2064A9y1NncWGW7kWR+tSsrKcIxNixzodoAJQDSv69w0zSIzcxcG/lNfeksSi6
C6wmeJzU76dOi8Cnr+Sw2KKNyDzTDHG8ODCt81rozZl1UltL/QRzyTHLyEaTak/giedqAjfTv8vP
1e369+hImkXK73nwcP0jL3NPmDGT2Du4lNo3hBDj2K21YP+Yj0QevW9MVMKepfmrzgllRjUsU8ca
VvwwI+YgEJnAJZQy1OxOUxgN5RYtQNIvE45K/pIVrB+UgCRxcGQaNJ4gnTWQZGvOerr2KssR6O2Y
JfGancJAI24GylRGq3/RyszfZaSXI5/h5Apn9UsPr7Ao5VBHTXNFmVqwnZSfo/yq+tBv+EceX4hN
PKv3cPU19QOjyBPfd1MQJF3P47l0ZLCXyiMqAIvJxT1/z2oJpyQtmRjh0f3xD9x+n1iYdVQ7vu9K
bxCMkvlQGUaLXNt+BIdKe/LS8jN/Gwiz0QBnATPK7VX0ThClLFZ/P8wMl4V0UdY4hCmur/saz8LY
08k+zTegQPnNp3J5KYkJTKBOSRmmncG6TxOXAMZGfmBRlcoWfiFdQbwfRDnp6jGiXPiTeHvVoq57
zEuYOwrCbllIleIYiW//FK27OsaycY02ljdt5ao+bjeYSMHsKePWTpXPPek39GpSthwgwOd3FyiZ
RN73qqnq+sjlNaaGOAfR4nDY40jEHM4Un3cPg5M/TKZ8pssX00FUVA7JD24OmbAII5PqfC3+bx5I
dIum4O5Mxm6iCpVLKQFuBdL9T3VJ+QvSyQ2zo9iKTZOcJjdg1PRtWZazrsLKnyQZuZKtQkIB34cg
FMm0ud/zO5v3EQb1QPuw06ayalxCqjBMZVxc1L9enomohxTUeR7CLzOBoG/hqQ3Bv/UniRpcWKw6
R9rQLv9jj/uXm5AETkOCvFizF9u5r28NIhWl986QOsbB6RWMHEAqIVoOvD1RaI/S8DKp1fYsQZtG
6PQwKHRx7exj4+qfrjuze6VG3gixJBm0ElEmP9A5uc+8aMbjd3LgV/lyincbZIfsrSAQYQHMZVHl
4QG0oulgvPYR957zzCp/X1PO45RJV5iZVQ7LAXiWKN4HAwejcfKtYPu5gkw8B27mp78pSnx3Z79k
ld+gK+Jfn1LUscGLHTUuuYNm0gv5uY1Jg5nM4mN7clPpWRyqx88V/RDsCyNW9KW6JBVH4DxCOTVM
eOmKXYpV9PBoLTFFq+4QtQXnSEt63tGafg/WGQtPyuE8aauCaSeIeMChJhqmvYTWMaYgT/1nXcAG
OmdqG76mJPHsClcqgwzo0V9snMDKdyunUYhhd8Ovny99fk2MHPqgQgCTHeqmTKwgV8mcWx6cSzdq
IVndwjibBAnqRP1wTxgkj7vLy70BkLMlubgQQ71EnzM+/Pn+2uvUO8a1rzhRlPFqW1PYSlebejX/
eCOugQmPbdsj15UmOfZI1wOxqVgx/JxFfG05u1d2fK548Eh2tOBwKKcUIE/DLRp+e0yFoyj3zi0o
VyKGTsb5qc0pZQNz1K7nJ5mXnulSmXr7fLpsbTkQHSn5Tq3rWVYzXhI1c1fG/bxZI6tCQHvj8uaf
9a7Ax2eELT8L3pCPM8/trCF+eMpB4sx7i4aQXS/2mF63oRRi19IRNzBGrEj/rnCmn8jneDYBB5A6
KzQVQVgR063ULwTvCE3BrD1Fcv6qKv0OZFlBtjgD5EQsvKTgJxI5Q79OZAmqIrpg1aj7qhZS/xOZ
pkPVntHBzk82SLl7pJYF8Kg+B3TwIf1eqsrvnJg4fgvxgYRDRX3SHFP1zGupbNXdmdY74zWWz4Od
wonux76C3E/SVjJ20ETAGgOPQK6yLr5S3V3sYGn5ncIlOSm5mzmesb7byw2po/CBs5lPpZed3rYj
ptq2LtC6WBz4AyGjym7lprUoovZ89cHqdWI2Sl9KRo9UNRMP6QFl5QrTKD3xDXLg/Ym6Tab3xNC+
JCxhxLl454V31fRCO720d79vBLirtp2oSVO99TXKKxsfaTnGADnkAeV4zFcJwC2q6JNTY/tBWSLF
u2iA4G/00MN+ILRxURVDgUGSe0PmGUDTQ6exLfpUPOJY0NARBdYuxNWywYjZD8yZQQ2QfSBEl0sJ
AtLYKVD6DABYKIfAn901mYSrmDnBeagJieUCAwIOQ4WO1wc1Yil1lZg1n2iojRQZH0HmeXXvfs+I
TyMUIt/fUiVefwYWyn5abZnBE960L9ZGJbqjMsM4I9u3yntgKpw59J2v8EDEJ3sqIC0ewFCbPbY3
VyNMghnNj2nMpCiG9gJpbZ6om0t7PIJ+7i0eDo2P1fP54uXY+hKe/al5s+wIOKo3EI4UKgmrO8gk
VBsdcGK3TVHYODPktYynwzoLmH+Sk9ZE2CGH/bW3nBjUMkPwN7JEGKKRAkaz4Cl5r9i30eI9HqcA
SIMy0KwIouY6yJyKklcxa4cDLOl73KUtEVg9PQq2UTqXpEcs484XAZWQCknrAAA87tDGOTPnZQbG
TYnEIhYU/m6sY/8jhfdHYKYi9QyJXCqw/dBqEZ8d9l4h4/39b6Uw0/duG+lQXNSnHpHCX7eh5SbO
H+4gNHSzBPiFwj9st6fN0YjxyqqvMneV0f+s2cBbBDg2NVw2W1bzEu2UBWHpl7UXK0VFiDnMRVb3
DNKIXiwsdt12sltc3oV+3GXMT/LpGVfCkhVpC0mhEh2RnxMq+iVYBQJKT/yVjPkWuc91JEoMT5/i
KIDWEGNq8NUJsgKIY1YfkDJ1f+dcZu3G9j6qRhqnJhhXpq7NUrax92gpYjcTMaRinQRcSMGA0AuJ
9/SVgJ53j5X0B57aprMxqI4TGWu8yu6XtzbhESIjlmVCpwzE7d2RvQ8xhHJ7HJX6QV/1EysGOiG7
skibecX4xFILBJL2MV17CncB1b2WZ+xPhg7x/ys25G7HFw57VAveeN7v4qeoZZQFpp490RV8mXta
BxFvKhef3b59K1R84ZeLPwFrQJH9lPjWb8athBG/gpKsbgso21KSFMNPurNrZZ2DG0KHVqGuq6V8
bZUsaTRehzHlmwTG6NNiC4OOGzlbrHUrWLgwfBekDzWuYVE5qhf+HfxqR5IFiC0xUq4Fhj2MNsF2
m5YnxYRaYI1B3GF9ro+U8htqqiIHcZSEa/Sq1iep1f0wGj2U2xPVSdghRN4rLm2Mb9WTsOX/uLHW
iHazMbHh242HakpnvojlHGMsBzPJIhFXxEZX8ZiQC+o3t6pb5ecSI7xoQgRN/IRVXYHNs/H7vYoT
GmciRh44IbTE58t8bZjqpWU0ff0RvmcBT40Ogzz0Ir8PVLzoeGWKOydlYDDVgm+OLcDuMxhBx2VR
9AV2WMQdX+RKDlgJHootRjIRc2JapM43lhq/XtD9dZPTd/9q35zflwuJFOfW33uj69vsgvibTraJ
yGNqzfxHEovFdPyKWHk+1iqou/WGhz9L9Ob2jgo/oAwAlTOgc74q/6G1FbEaDp42XcK44i1CNfxA
yAgP0QKSyG/+/52eQrNoiNMp18GzOiEgjgFXjjZItMyJnFLwdIdg6V7axMUfPoz0PEmTYlqfUtz7
It9advY2SSF+mc9iHWE00ekbrcgg/UM12+3l7RS/xgcL6LL54u4Ib8cJy5/XsxQgwlVvB2V66aph
K4IB+zJIDINzIqaq75EcdxojTpLPqyV8PX+YulsX2o8qMSRvVmI24UBUUcHe1ydZ6OFgk7L0rOjv
E5mDTOA37a0GQd5M5seLB++x/yUoyIlJ3ZHHqoESWt6/5Zioj52inwFhrFBhkY0dtNQxUQyWS7+j
ISkkZqdxP417Bak2UBUOttvBSrf06EgyUytfbwSV8FZAzk+l3mJIawEY0xYGKIekHCt9/uDqykWJ
lWXZsaK6wSdhBjO6EmjKo/8pt01WiiLxNv8dPSlCIs+ZgKzeFAJIwqdQJbFY8bB0LGdC3+Ilc8cp
Gu0typtMGm4BfNk3zb9hmm5yK/kCjvjGPjJG6bRYKYeP2o4Epc4xjgFpxPjHDNVeSzLlHzEowzhO
aaD/kAJMrUWjQpmHd3UO0Y97Fh7ipQKwH6F3PwaJfIz/XIM5Z2JFmfME27jYdbsM+mARhH3CAPqo
e9BoqQLrFUCHXbZg/j8Kumq2W2oXXreJcrXsVU0EQvZtLylL+eshR0ZzCvBTFEnkjfYNbIjWVT7l
4JpRmxyu+DgunDviO6MZ6IIMF+PJEvEEKpuFTbTrki41c5gbPdui/WyvZVTPstc2FcEMjXhWOTn5
UvHT0F2WNojzi1XjRMF1xD+XAfNhuR5YoqqaXD430tGzXeBV/5o0dDI2qxEay37rnqgVS7uUD3j8
zBkcJubwKycDN/oRFwShBqzeTjjb40Y7SCEaOSaaPCmod61hd64r/ChfcqRQoFpIJEetifigIOWT
UrhQNjQDgTiQHWC1BvIZnUT9wjYH3p5xuE7hAYQCBpi2Y1uqihFo6QjubU4kb4HAjkUnuJ0KM6Vv
b39hS/dYqk+Ez0qvnCqsG8rHXvefkewuxq4kJYewEWKPQkDjVWg1kE9698xALENhBXCfZi2+N/8X
YGsfH+AcbhYueldmrhnDhv69taKFvFRDWES9KPwnS15CrUf1tDmzPmXrsch7eyJRlvDLzv7izPlv
7tDMkDmW8+uQMPGoGZxVwOrjoEOzNk3lbXLifzxqjh0QfZax0Hsq3wkmny8BnB08/Y4kgtV6nBq5
W32nX/m/U8bs6imiotbH5njyLV1MXMoggxF1z7WoFQKXgHqYabZkKbc0fkcoUvegr4kYFu9t55VW
RROX4oLB9hJjx7Ad9WSzAhdsztOGu0iPKu00vuAwQlvGZRdLTDxeC2AX/QEFXduIAdtc8KUKPUCU
M8Yr40yweMKzgxgtgRs2pd36xc3w1VeQqPbxEw6APw8GewsjEKwkNthvMPUeVhFi516I5+IyP4XN
Uv8N4bFT9W4YD/mPWjJnVZ5ZPI49hTgdRwzaEL45bc4/5tRFicELP6t+RElz3qkD+b/7g0+NLNY5
QdvcpzH8DjwEMVyB/YoeSyRhPnS2gjOwcyuwafDyF7sZjV+weZB1TKcwlQ2GtCc/20Y48IsIS0Nk
TshmCqht8Thuj5QIP0U2Sj9EgWZZ+7j1W39NmDwdcjkJgaJrnNgM84AiuwpkRklvD9HcGGWjUzYq
XIW8YfAa6goLgeGR1IVS5IO/EW8yS374bl55C2kf8Jl1iF2X21NWXCucAOpOxfKgJDOmguoillKq
WYe9ldnRjG/TeKYgUEhrYxchdj5rQHAdmfxqSLEjPvtw3B5EMT/+0A536btyreUmKeeoOWtNI43Y
7LrkKYVahJpX91J7tInxPtIVeOBi9SHK9GYPkQrLyzvqjAmrqDXZJKrgyfOVFEn76I2zGExmweUO
MjqwasMrBqEA9+Sq8oPx+wz6f6dpOo/N/e7Xr11DkFsjP/RBWnoNH4DDVZYjtMsRZ4DJMtkvKXmL
8dbfGa0gQ6Cx400yef8yeUJGiMpiYDMQaHLHohLM3Ujhu3tC/waaqcypAOkn6cInf61arbBkUWby
gdZ5mclcbPUZapjWlbnN2/uIk/FCCo4XcdDYYVDdkfsuD1kPW9MInDjXt2Kydu1sjbluWsbrB9T3
bPeQdEuWdXzJ/V/mhic5NmAWwWJaRgEclhbBHLgdJGG+nFlWHg/9EfKf12y0uo0J0p5GH6jMlEIZ
bfsm/EeXsyme36GvJF/aTSP2wN+QeFTjz6Adqf/4vISl9LaqVy2/eW/BM4qas0w7zvoaRvch9xFd
gwChV9RFMtU80Z48XpNLqyjp5YJBVofNZFO+h8AyowgyX2TNAkzboXTcnG3Gh7qffOuNRVkHtmDZ
75yzHOjdsNRk/zJDDGLgxE1Jrm8PFplYpgYwPZTR0zkUx1+89x40NpNtg0nDcFnVFKHfsqlWZzw2
NQpKfrifPswafeg0h7z5OKz25+VrSLEUk6wjf8vSwhdnpSRbEXEsF9edcvwmdeUWcUFBgiAZ6/V8
A7FeJ9ECAWoLnWe8RfGwuyy9wl3NcC2OqU6KFFll16HqIhPOb8dVhtFe+bSiYIDrLYKtMFbiK14J
xLo0+afm5F7HR57IaiFaC4up1rpEsOG2nrAdvxUzIn3BkodNoK6L/GTWM8rUXQXiYXCTv+QOWAPu
X32vrSLQfdNX9h9UvHSYJghzPi4dnitPGKwSXJK/n8RSkRMQenSRXS51KdBjnwbtzYs3oSt8tw1s
a4874wt6D75wSaWaLPgcHqdU7YpXKhYRvFDUajkZUqlcEu5fgRAE1DKDwNquhhMC3X/PDsvCf/Pn
0kghx+eDjsJSgcUNKw5FqOkLJICVcpQV1E100Ry3UH7sel5mhhwIqM4YZlS9Sds4qe7k2Zkkm+3i
Mr3ZDLQnxokeqS/7ujPkJETdeSCLZITMnFf+9Y2nc406W+ZUK4054TKRf5kcSi5cBSmo8a8kd50+
OyGjGZkQ06R9vBT6h2y4urEAD90mQa0sln6E3p19Mys7aw/bXDISBNM101ab3+3ki6rNTJ6lWPDV
75ckL/cKmSsOSK/aSsUncavRvFpRqjx/cuicTdyw5n8b39mUtHUBF1JvPHc2/wz1cot3AXoxgqhE
DvzTzGgBdH+kKCiLFxOX858jKWdpOc9kUU+8NF5k7EVaoBEsc7iFaGroEVv4XjQVVjZdi/CheyZ7
VNMqSYG6NMKfjoEvIFFUM2yZ4Xfthoi4zSveLoctK/rRavP5tQWAf6OB56eSJECsc/y0HJfYChFL
Txvwj6ZfWGB2a8s/2eHSHicV2gRHz9R+VBEaRugAdlKR0HFzrALk0UMj5vCK8ymqoNI5oMgodKi/
fzDB7gbobFLqD3F6V1u94GnccufXchvof5CSYIRNawPNatQVgeez9agBhXs81ADianhLuxUTq3nh
MzYW/xqVLgxumM0DunWeJt9MhAaNsXC/0xLgvKlipdJrAkhbVK9qPxzty7ZcMx3hS2PnjxyiIchb
BpDL53fJ+J3IygykHSzY1J6g0kEiahE8JY6ugETgttqSRCvnmOg1y+UhI+7T2TMEyXWFojI+7mK1
/u8ByWKbTLIwv4NmyB7B8pbdHVLIIDGTVPh+Wan8UJty3HV6EFW3iAxmDlNIO3AI9haco0jOFyHQ
DPPfePX66Qbp2y1z3InwiWXnu/5lfCKTYMXoE60I0YFtkuLM8T9xn4Bed4VvXc7rGidwva9/EmoG
HWpW5u3bEaTABBmCU40mDh7xGOBUe5z7MowPTldblEFMuTJb2pfhcki6gxCqWICQhx2e6QTQZqQR
q+hxOrHNzCwxwji/P4DdrXNu2jBb71tzoxmcIlLyZBLZUWZHIe2ig6UJIug6z8W8NsYBpxgtZcYX
GqqnvF3vyD1JD/8Tuvqkwda7CE9c0qwbtwFxUgNmSd5JnIVIfGM4wfhQ6YSq8XjRZQqxtvZGCIk0
Xnwz5Rvbz9qffNh/f/jrZDrktL6kHC1OqKeDLcrN80jWsP4HLCGbKSzlecmWYwWLQt0TfTipdDbN
VTqbLEFK0PbpXKAYGPDVfQEoY7VR8Wrboexr+QVu6xtqRhYSf1z4blHEj0foJ5bCayj16pYjjZ3M
hSg015UpqEfDe6v/1wJLIkTthQo6bSa64L9WTx6tUxj+oQRtTRNJVjW1V7cQVQZt4AthyJVNUNXe
juVAE5Se0V4w+ggS0D8Lt5lsRDo4p6GbOPwxubtqkmyqF/n/M2aLyYaqTtTq2MbTeAUjm1IxK3f4
aizwGeglD5kdk4O8BaDoQeopEuwW6dDH4ihNbQ7o0qowC0+swCMC0vB1R1olCgtW7Q4HsDa/Ps/t
+qM6Pd7uFe+j5N7SzARCgVzrJkXyY1SlzcnBJkGG7yX8BFyx2xpO332y/iKdW+rTYJsS7BDYQ2Yt
eSqvSdlhwueT4sR6bASISQWZHEU4aVhfuyp7v8isGROXLdRMtpS4RA34TKdr90/KY8lQdFKyiUMu
WrEOaIj1hiCnrVRoD+RfC09qhxVQfp6dlInIfFmRBM4B1SWjnCpuwyxGL3lW+LV+vYP2nzHJu8vI
MXoeccRVcp3J8ri3FbxplmsNhZX/eDybmtCBW8wvzFmWk3RMtYV9A0QNmh0i6pzSDwgPUtDYVXzo
13kh6IoTff7IrR7P95p9nW3vbl8wVNrFGKky4WvWpD1LUiqohz/QtPdDxHd60t0N6zQVWZUjWXYT
Wxyb8o1NqeEHfn2uk2lNEVnKEHzAoTahKJb7FxAH6qlh6GiXhf9mWTdJe7Vh8DPMJcn+jIjayxQd
DvBOJqV2sL/LlDDSAlKNWkMm2+1dp06euXLDhv1BEbwYP7CpPweb5s8sW0AsBKk+jwBIvh7pppJk
2CcJLjKcSgYXv8mKdqztCnZzuZNMDcqxShq/QDksPfTz6aFuaNtVQRhXrmgm84W1weAXlBvBnmQL
NpE79SDH1MP7ASG+uGc+tgwpXxbNxUvQsxRccBKDUrUbNG4sy/NcIvG1aXSt6IpsNUrkuo6FJFgs
0kiKZTH929OkqzyZPdKh6pguGih7Xj+Tp+RrxynrQKgB2MX0XOk0Emlv10vwLpDWS2lcTMXDkicz
TR+CD9FaEOQfustGz2IdFiRg3HUAdZxC83ivxkMWa90gPsaNhL18ScAU6rT6PZl5KPxB3KKxB/Ap
Un10aQJ4iO5DznqRmjzwR+rZ17TOtjL4N/qwTAYurzZ5eIaqZ89bhpxrv0qkdlwQUxLQHIp4huzD
+eDv/7RlTtQF1Ws4D8vCWVrjW5bhGVeTqfKo6/JJTbPZxeczrWWIdhZhGlPu5J9AQ3q+VnK+BnHs
ceihVzvvE6znXwViH1o5lb4uflKm/+sLtGMTxOAKYEn0+E26LT50XUSLpGKKeEm9fv6QQf5A67Aw
SjLKvNN0B4/cervLFphIr2PPbpS1Je1TYTtbffr1UJ8NjUMHin7WOrAlO9B5vVRUTNYrgEKGo4u6
ZTLvTuGAAai/mMDFw3tO6aGfeBiu5lIJkt+APICRhhExak2nWQdn5z53vpgprfM+EyUUuRIcFY8o
bP++zhlv6BQG06fdEcxptzQ6+ruHVQMTgg+reRHeKOp7tfftR9hhpSuwSGKAoaq4+0zaNHS2jQmR
FU307WNVmiVyUCxqsN+NZJzWm6hx6MN+GjejLZFFrwbml/Kzcphup32aUpe7/CA4kwuyST1QYmy0
bZv8ke5qVNO2SZfsH86PxXGSmOdQW5Pw/a9QnJpOClyRujoFiaiIeZCybEmL1EsmgTpZew8bARvF
9VOeg/4ZPKVroLMC8ucP+qy32JzXylixtpUnQqim+7i5uGLujcXk8MYkXauBMlfsuT82nZyxcl/T
vHT6S2VG3euiNKAJGXnxI5+U81CbkjsaU5JWWihAO7Mlg5HyTUQemYCGMuQ6LsC9TKjVPNw4ax6V
PiLz7icmylbkfDdp9OQ3lsNF02jfUQhYg4YHd1NjlCiUflESC56XG0p7bHzEB/ZPsiAmwlQuY4jf
AF3jPuxA/ketyzO+0altQwwCTCvBvdjlj5PMtCQg41v8v2D6/GUYFA9NS22+nYH4ZKvpSo9KFr9c
gkUw+yQ/s/riJ4Xa7SlTG/9nWMQVbrZgWyba0O3qwYYVuDObOZu9T/ZSRqnOpK+1r+Kz9SOOXgPY
jgmCVgJxIw58ZVahrWQ9WzmyQ+UBOAvBTEtpUVb4Vnyfy1s0ZJcOpHejt6ifHkyawLujR+7xpChF
83E3yfGW0CpILetyIlAvpdVtDMrCSeuVqfjuLY7DBXvAQff4yre1eBCL54+TM3au71cQ5GOH+P9/
lIExH26e+iEAWCHwooDWzi2QJNMoXDXqHprwEAIuBbgALDUHJQfQd2whqEDrd76pGhdX8n5J6LkX
nZ1dViSoNcgxPjBUQzL9YjWerBc16N6RNKYS816mg/y1oA6KLfw0kpT9cLrtYnDTF/IPkZBZRGgn
fIKUx/curu2WjOcM3aEVaY16Qh5so/1BgvUJIP9JeieqDT9bXJkj5EutXbqLchLEAukcCIVAEx5a
h4s8E4jP5YrdBi2WrUbVnP93clTYX731eLNtVrDP9GmxMQTya14Drkg5bqYex9gH1V2pOEGbjLdQ
/yDs9gMIQ6E7dTQE4tmVV/N6xAQpX319PxFlTtkI7JIrVs8SitQnsmomk/qYHmeO8jCkMGvab8IC
ltSUQCyQ7kedWjqLbILt5vrxMMy0RX5a/Ajj/wIZtMAogk4M0sxNuKWFF0XeRg+ANLj7NJ8CRSiI
jYyzz79VI4XEvUdOacLF4xLBqjs7nV3clfenApyU5LHgnFqxY6N67ALtzX821xeIlDX2SKqNR84J
dwbUdQLe7X4qopckyM7hTlfqt31TUSIHQ1vYFug5rTqxLIktjQjsqETEQ/u3X6A6rPBwDUPhjspq
mGySxntdXdkEDs0Tr1u85jiXcci0/YY7nVXQmeGks8lUDQqe0x7SyvNkayjCisFR0WympEBFOWNb
3QyMni7m2HiqfnhOq3l/HFyP6gYkDBW6yxFDo3p1S5gdHbliCusajVuh0nfdBtkipwVsBzRADdA9
VaQT9IbT+EhDqq+F37690/8PgWlOEWdXhORkow1qHCUAOTVMi0H+8NFOJXouGA4TTYexFyGX1RLB
Vs1lviYpWOcdH3folyYsCoPak5f3GT6AgB8j10iSOLmdrj7KLzso0Z5uHKDpQ2gUg6TMiRxPOypR
ldgs9+9IBI/WVCYTyawomm8lQhi1p0Ujaa2dOO0jgX+d2NzyuU8k+BPm/4vbnAObF2u9tKCMMUev
+NQIjORXJLJ11OR13TGlZShWzBJXd9brL4uhllmuYjcpCNC+ij32Yqt5KKVfu7lzTZ+QafWdBeU3
KjZ89ZNpcLc91WWsa4d+LqN963MT4sCKoeOqhUz7H4R2rjZJ+19VBnlim9OztZgB1s+xcoLpHbJX
W2FCfzOZ9cKFRjHcbiA3mO6hcY0PQoEhuoukudHWKIbPY2k0sN5tvHACk5i4j34u0J9mu/xJmXq6
dDr8ht8phUHoecfOSV4anMNaHav5W/sVF30tFpXB47hEk2b918Wss6NH9Sy/vTMQ4QCap4UwGWKc
w3uZHwoWwhen8Eniozkxpg/mBOH8JXDALR+XOjQ2kC7llmL8ERiRhJpnCNM9D7HRNd422up5jcjQ
1rWNDApwi3Kb2qqnIy40JHzmFdBFY207ieJvSwv5TuVwbmlnXWYyt/zq1sS1sZjZhYH4IItUwV3x
4H29AoazBaqE4151jLJDfMHOi1QVBdP8heT1YfEYpGuJnCWcuyVEc+B9cLJ8hgV47NR9MUn9qOdU
gm+Ey3U8RvDftmcgDk4LqjVdMaw97XvldtBun2iJF9s6tmtq+VMp275xLZAoXrhe7Of4K+sYUCcp
stXD2RiMk8+hKrfk3oHuliCbSCqCN+6M48i1SwQYe6Wzt8RvILOe3N0pVzxca//msGidvHPx9YyK
2BfHOX+tvLnYA8bt9ocLZ9vRGA3a3hmMdB2o10F+hhIgw7aGN2ZOoC4Fzdwlxov9H5lW6ltVH60I
rpcAw32LCkOFKJwAoRniPvMONU25qpwxhd07DD9c6jArstnapcwQJH2sJyjHYBXCn82L6MB5SyTH
jHsjYoN9QHQm3WwHNhHYhU5v+9x3H9wMfIccc2iAQM2MTfwtmMq4RwnVRSwD4QhwcpP+pwh6w8LA
/7zmYnAlsJh84G9YvpcSMEBwD8Y2vYaD+SquwT1IaR4DS8itSvSR4IIxuKdrbD0SU20Ekb5IgBuD
PVIPF0No0Uqxa1xsSCAm4xmfjqgBguVgC8HYKB9CLydwWfQ5UM7Z/4Sc1HcveR9m9g1bXsGO0QiU
ViiKbMzvaoxjXoqm35si51amPeETBIa8ZgoxTd+qvEHIuZOPbHKYluLbDluGXur2a51mpGha36PT
pbqEkVzqsTZvS7x55mQFnNagtynpYbsK2mDT8BdPpWgLvz0pq8A1rGi669SGyNb22HN0YMW/oYvr
Ai5r90bVzyMH2WEqV9d5xNoyTKyZsShLBSLj5dnCEeEjjssjg2Na+nAl/bFMIw14riXQSRRFAb+f
vsLYtHIh6aGrfvcQKk2iQT4xS82Ay5suQbqMBxB5OW4hH4wu1hB2gm6sbGIoNLorbypSNCE+8BE1
SfTZb+Lgvr2PNudZbNEef52IkvVcsXAHbBgt7qvv5DOcXitwDK2s+f+bm7Lq7urZmjjfBlqVo6d3
w0K/HJX/pPY/uhYZXb1psH+RiaTFjMupkTbA4w2mEXQvX7yrIqCbVE2jeX1cG7ON/XDDnYSqqCxE
cBhlSEYAjaKkfCiZ2hWe5iEsHpFRRMj/9+AK8kcd3HV5nxyzeLFMs3JCw21lVX3uOYiU0NQ7T08r
3IQBVyhOIpRhw8Ws9TfQ+I88Engd8NtLP3WHP3lKlFK35dyGPJPGz/kFSDj4KBwZhKOlUTARr3hl
AWNuAU6yAE+rz4sMs0pETsatKHB1fmqQvsy3kjk8HOHyQQ5HJKOgVa9/cOBJ7MPlPfJpsTDP+3Td
DK88TYTj9TVcB58aCGgGde5laLoywiaiQY6uMZ2BGJESF82yZ5faBcBMlZt7sbAuKaeAG3/Nl7Y5
iEDT4NmM59azMKAoluRldgz4JVoo9ZVhxoCYjvtIG6WCcoml73gBIiht51U1OQ4XRNmlkaXYA3nX
/bk3CbrtfApjud7mIurhyGNc3Xhmf1JkG8j5q1KXm3ogP70AgocYon0/BIqHNlMV6dt4suoE8WlI
N5JgLDMN6lmcgJhAOyOvstTWBz2ceD8z1MwHiiA5naHZyMMdU9kfVuW2P8YvDznEMRKtSYrbedjJ
sMYLgcThBWZlSLVGk1PXMw5y+KDIoGH0gfzIcV2pUkTl4GWTv414MVY5GZKTA4OjPBldV5BoaT77
TXh0vncjVCGvw7uZNlrZJLLAsMVF+FAFcOUjIxb6Dk7PKDKk0DG19kBFoinMspG1Ye7w3JoMj1aE
GN7Id52BVO3rH8JslO9NjoZRaQpiL9sUZlKEkNcaxFgQ0fHoB+8AsMKtf2f4S7u7QGNfnhcwvInF
xdG4jqtC/K/f0CWmv7eR4lWyALgaYD8TH825w3Rs0B8ia88XSFE83hkOPQzTpJQ1p61mwTO1Gr5A
Ox9qNkMNDW58feTeTX3WOrO+0xwu1Qw9ExknEnYm7F59fZ40RqbOrBuaz/OzycYoha9gyuWcqyQI
c+XH163rIJfaYyuvMAQCtniR1FvVkFwRT0ohcqVLykpJ0GJRqAhO+0Xu9YIEOz43W8oxc8ajBm7d
pxQgFdCcVyTr9JqoLW3CG89sHilzrEFo6GIz/PhFGFm7r7kOuZmtRrBZIaLnVBnkxnfMLiWfbQt3
eunZ7wWONtfErp5Z/sCEET5RIOhIqVW6Rnjvju/kuCd95rMIzNob2uyaGSHKmVs7fSHOnJNHcnlw
N/qSKlaW2YJUMS1MpefxfUuyYIxSk7bIjXpXM+yGZGmHu3lI5DZhNveNYUf5sW4J/AnMNdSVxvqP
6DSAGz8w+cOyg09P0uZ1f9T0DSXOjRzzq3lmbYyOKdLEKdw3+ukd+4rzVd79tucqtPggtGV4BJpN
d/3X8LKEn9KpidN+PngbrmNa+05R00SUX2d9XHRc/pt3975ZHTFnxlB2RaQzRnF0XXMBE/Opxpth
eJkYPc5JFBLwOoKiUGER24ZkY37GI49er2sQS0I0u5G0cnFtlr/36a6GeG7UMXOaJyfA+J7CyBFr
Hltw2OC6//bvdkaNDrwGlVczaHZIw2pdbJ59R5/6RIsqmRoeJQEkrRUAWuJIKMPPLE8OQn+8woru
kRfGCXuvnXef3O1sE4+H2URSp3TNnNP9rcpvRygRtN9TVxjNEQ+QYUH4g7G3NAk/ov5WRfmtvGLT
dzKLgAp9pOBZhM+zaJRqSd4DGBoz5XItqrwMIYwSYG9meS46hvefpph01kJ3pNlmP6jPwVT+rIGy
Izj89b611vnFKibjl5i4Pu4D9e/l00in1PgrM5PhjQvpB9ygCy4GsC+5UWai001qiKHV9S72wQ+G
1r6a2JrhMkEZLduGiUy/6iMVjtV0Sv7EzAkymMSVram6iKpACMRbSMHIFuvm2Q6aUCfq8/kgmnUE
IPsc0uafrW4Kr/hOHolwMccBuyET5OpapGmQY+SXJvX3DaGmkXeV73L0FIJR7L/jdGyWZ1guWngz
4zw2oEfonkw+czKa79TXroHm3u7cLAe58nqgZHNURn9T3txCOpnSRkSbl6+txkFekEBuf2N+Lvlc
n+5m3ALmYYNZDDX/8i4v6CEG9SNYSqEGbxEaQV/IBUnKD0cpprz/QgOfsg69uYNOTdqdsCz0yQ1w
JKQ9wjZcoQUknlFYqa5xabfFZBdW8XK+g85THIvK68Ka3BOIE7NTjp5sfrJdnNlDLZI6zqJa+qPw
CscXSdp6BAXzCeWeG1CJSE3dublPo7GxD9lGtLFKmCvMNdDyxcF52jSqf8wfmmFx7zU6/7pOXWPn
4IQpn2WMMbPPT0BWhcpl6Z+Iviqg5fk1pIY+dO+9PUFOeapeBaylTAkVPa6Mx2yd7S8irjufUIwL
UPgObyduAQ83xsysbzmDXu7kcLGWqME6IOKMlLC4+1ebiuH6iScN0/7BPV6T+Tad/6TB3jW69etH
V4TmnoJCnt1HTgSFTUm0MzZuFwfsW422vCXoCTbi1TUuflH3dFuQrThLiFGXCfnUqW/Q4ovuzz8j
5I5yHKWS6sSsvgg12+TJu94E7C1ss2usNmENAzKleDwfPDDxoxusZudV28KM1uufMOhPQMTVhEjf
8x4KasjaYfUk+YbZ5mtAktjKt9x+RZzekr1SzIb8nEmH4EBQYke5jjRbCx3S2ip5xMtx5V3XRaJj
1KbELcg7BpyixrSmXpVLlMjUdUX3Az3TUt4Os4fCgCvzgVwcBOF1+7xZ/GFUxPjnsWmw88/YzTC+
4z6COELLS9OKGsUyB6pm9kPsIwNdNcW4hRdiNE7aai2zP6A/MGR+oBJ/CSFbmcfQaC/k+z8S0X8z
TR7S+9GTEixQTFJ3fSihkuA7/cx7DLap3S8BmiUV8CwudFJ35l11RjUhKT0ZACj5dvHgsNniZvkg
PBXzqIrtGxQxAewZDE5knpZFla5+BlpwGkADqH5hiiA/6In86RSAwM2MmacWrvOWcgWkroostFs0
ylvtcT64xEMwTidKSRte99cwYe1+Nj61jfdH1yHDaBCS9zwH5k3RMTHXTBCf+xDWcIzxkKyBwz6e
8rPkD3TIuyjUl2BoTg6Eger5WY+97YnqSe/zMv7e+S1mzo5HXet+LO7GdsfOV5ivlFJroegcNf0G
cUqWnnBeV/nB2lRhRHteQ3bxB1Lx2Rx7j8LplNEPY09A9+naHJQmOQjq6Elujsb6HqcpOTOJwUOR
b5fa/nEdaR20YP+zeaZjsmfjaYQrfZiyTcQbMDWWyLRKxnmhBDTCIwIW7N2gLGVs6KKeksKRGmc/
hWzDAQkdIIuPuBtAEKmmTliP7M4lmgpSEqCMrZJLtUsFYAkKl46oz0bu6Na9+KNBqm5mdcRA+05d
1nAGH/AyeIAJRkIw/ZLeF2Ddwcog2ZF5r3Cal0r9XR/wE+G/+J7yMY7Zn/peqEjpreaRvYAWwKeR
GizyRSJJNRbdx+EAf3PR3YfZexvHfRJKIg2M3ZKvkW0augXXz+1OmVjiEkGnnb2Rvrj1NfWR5Y4H
9O4U96ot00TrFVBZG/vvmoGbxk/e4fGiBICUW/74u93FA8RUY8dPmg/nHRuaXqoVFRxa7XLD30Cm
NtCnjsTkOBSwuza1mL1EEfv6IMqjA4w1Pv6w7uZ5eRVgkYJBLh3XWG5tjbLu3/oDlqybqpYq4B6q
n7UxBALYCdCpA1HnmD48c87gEh3jnq0rkLaw4iYZQj292f8C9UncDpp53hcHOw5m/ploG9WHUPH7
w6eP9FSU4LXeXmnzh9gXAR2gYRlV62SpbQHNK9WJHnk9p+wH9Gq2LOePFW3qrfDVK2+ScX9JTRUk
Pe9NoUVnGPA7fatE+6qgQptFFfEUSNj7ez9MWaPXBepmRJ7Bpw8M+9tv+mNelKqigvbF3heoQcCu
1a3+qfGyhP42cH26kfvzPusAQCU9DdDY7h2kHRmwz8prbBKo1NoQ+aPoBe8y5lZraspXJxclrYzn
yxW/p5nmFGz3xmWEa+lI15CKzNYsE93Tegyi6TiK7fqBxUYsL3kHKAsDyXoYQd/elLCBBgbyjWGT
RT5YjP7NiosnwM0hd2LjOcDb/jyv3E/MK8bNk3Z6Hg2vvZhulUi7cqcu6NQ5yXZl1vBBcFTlstgB
z5KE+5d8C4lP4CdOJFFtdio7FQmiizKwM3mscWRkyRqeY1M3Lj4nxSMbQRxCrFkym+DRGeQRUj35
qPFw55ivLTejX/DA84DZ8qEhSkTiSKWIaClGS4ytIwDJvdVNlol+qcxSRPrb1XH4latbRAt0BJJQ
u0fcG3QrISDpnM2MDezc5doW21xxcIqF+1woq0yMsByOKthV24DMTmTjj833T3VTBN54oal1v/0X
O5TaY0B1TwZ+XJUxc6BAZ4K1oIw/pWy72j8dmiIBHmZmpW4oQe0+I6s3sYeyDmqTrfO0M8c2A06W
x312+UvAuvqws9iish8LEm+Nzr+bE1hjhmnBoQnInsqDpHnBHyBngPSfhAgf/L2MGvbz0jrBz+Au
tq//aqauHjibv00vkP1eJfEcJ0NqgOVP7I6gnmj1UiNArm6HzAv14xMkn23iUPWy+hRZ0Rs+MZZ4
7CZV1x2eWx7qHxOgLd1mac64VVb7jH9NHiLYkw3kAY4iDX6Q1KWJCxHvRdPTsvz1Ovzad7NtrCol
O4Dcz8OY4pI2JkmCvXur0lIr1VvTU6T80xCvhw1iaMM7qwRx4wcJ3ue68Vvn40/3TAyUVUtKbOKU
84u9sHpefJBHcgq+lT2YsaTA0gN44nwhCbkKqMWaZnz7wVzdpJirjASMtfZ1Ox4PpZ/1BA4ebg83
6MuXGTyPRD2vyjcb/8K3sNvIrh2HDVpGcWGcpcR0pgSdfNNEm1xSShehGgyfIcz357Ld01pY3v6B
AT6qn3eN7MBKuzb326bLBgzTOTEAbGYGUeHoH9P+F3yg16dYuo7juPZlYXzPP7m6bA93RUbzcUfd
Ssfj9hejIE+Gnf04JlmtANIH0++jKmKyt7KdtVI7AcTbcn1/wNbvxm3Jr0bpzUxUxDbZWo89kaOJ
qDOX1Zy/3MFdjXUgty+cIXOyArTMbW0IjZ+UV0cHZfZZJ2GHwqjFv4i5g3bdwSh0RfHNJaZq0sZ7
BSidx0vqcYty7zeHLUFvVoaLt7hOhqCd62FSrsKZXigXzeks8W7hYHkaEHqgEwEp4UcbYZl24q5/
4mXcVNNXXxlQEJZ/gRYKUVURgxXamq18aHpY8YQfMymUCrimSHHZnZAU8rT8gAezp6w8Lrj4NnJJ
ISPRZVxjotq5J4GTrlOjv7d/eh7zpKn9Po/J0FOANTRIB8NZ9iFKSvhppMoxCvHiW+JBv84+PP5a
x6qgneS3y/zQ8g7JMfwMJQPG+R1fr3SzGJbBOwA2HSz4gq/s9uBE5cKqnGsjLTwnXqF6HFMgwJIz
Me4v4rDmJWXWzkHaxlXJWleY9/KTmpdysSxwUNcizKp8hhFFweTtPNKWULqKIiHWRlhYeqEX6HO1
xMt1FQb+fFAm+kKUfbpLtGcO3qMb1TbagXTgeBix16gAu5IQzjxfHspiEy9zNEQoXricwNRI7K2x
7Q/45FpimZC6d4dnmlJ9iXTCSOHlSE8FMilFYtps9oI0J0uDvmqJxCA10zq8uijz7FmgntD1ogTo
WflPwoC0Ts1NTrBOakFMLe0bP+4gTYT1r3IAkVWbhvlDS8SxYjvtgT/mUygDHYA0e3FCg5PItqKM
omtTXPdvr0RvR2Om/cv7DzZJJcXwVWU+X+tVrgtrv712LpFyOSPDUWF6fOMlYTZq7YoyPz8Eho4b
75h/W6lv1Kq7CQk3YeOD0ScpCgXtvRqX3lIqT9RkLiH3ESMr+y6LUXFda/Q3S1iJWDbVh2+HMFJy
m37zVl5EwY43EZBFpovVosTfKP6oenichDN0P0SSL6SRlBpk2NPsVbJNdUenhEnSic4ah9oxEEzh
wyzhn+4heokACY1yWK2VlLFlew2OirisXezcJyecGViObCQUXk3e9iInMLeiIc/A4kK7WD+7rV2/
NLlvJwouQ8CoLPG9KIDs9yBQa+ZTpmsE4mgsfiM53CjtlxCw6up+d9S0p7MU7Pd9S2GmWFJSo1s5
hXC0H7ZpRo5xBNbeLF/zoteZvvzA/5X52iXTp4ieSEiLrOcmW/tXJZ3iMsRnyavzceLwIg6m51Ln
61pdkMhpVxgdHIrd2/30sgkOXdywxig69p6Q2x4tq8LWmjggCwJin3GI1/NTHANz/fCF5CCqWc67
cUqLlwwvkmti5LVBgojgZ7KrGvsoZc6cama8UIbV7uHoMV/BZzen4vt5xJKKyf2jDToTBiFJrnsD
w/BdObp3yyhkd1pw1DWC1AV0kueUxjC6dxHXDzGsgHngnudVkzsj58j5W/h6ZsFEcfhmI9PTKot6
tvpYfUa3HVebcB4cmdUJAIG1yRgHLnh3RHzKo6amNh6v9ETHEaxxpOgmfgQ5++lLw8lBLiWRS9gk
MUKw871PiI3v+6Yr+C/eQyvZYbxmk2lQHmbEVES9bIK+tKQUZNR40O32CEXZ+2+y7BVQ9YRQaj7E
uIKF02DA5OOnr/kg1uSwdOyQfw/vIWZ2NDUiOR2R8zIKyy9Sy4g/T5krX1dX/VNY7/3JLxs0PEz6
fisd19yg6uOdf5CHoEpwXeaOIXIyyndj6DcV3mfsJbfDJW3vi+H/6KRC+W8qkrp+nTWucn2s8VMQ
R5lZ6wqlN8ARzh01Cs6Qv7KQSK1bxX6/RgTbRiBAdtk9Kima8uTY12+2C8clIeT8xV55wz0PPuOg
RZOwNXJONIf1SXC9iLgC2ottluK646TdPCvxnMokD56RB2KLd2/1pat7xzWDj5hrGj0pTdGHwgYh
9FFVulPwgUVmqutc70pTqWzDvoZqn/6Gpj6tDy/a3LDr7LN/ueSJR/3eDWm4l4J9BSj4yR+47IUo
WJcx1kAWEDGjJAvmnyN1S1X/2WfrqAVIrtQQS3UjHU2gbqRVYWhtvyZVR9tiyNR2fPX883vpa8Oe
jgDDsT9cg0G9StSSqp1/yd+XMBOau2vQQCf1gAhsIXjkBn6KjyQE6SFMu+rWgoeG032CBFbstZpO
3HaqIhIyRPyMC701KJOPBql7/IP+HzKckBuBo4oqlHdeEzRRvtcGlY2u8jfuJ87WNn1NsudEYMP9
UsMYNXfGDUuHDvbKACv0AJYjOeF3K4KRxYDhPgfGpaoN2E6nbF5Kx3+SYO2t8agUCw4jfLYsXbGX
a4QmcR1Jcy6z9BxZQ/hwXDSrfzTKD03QF+2fLvvHULmkqomOJ8fQE5r5yWq7zvXXaHIRVgs26vq9
XwZ3qhJHqDymfo4Z7B5a/6CngiDHyhkNcUWbkgVwJ64PhcYyuUT4gHVcZTnbjXrDTXl3NDlaIimf
70FJ+1Nx7eb9euLU78inTRb6E0m0BGGi8avMhOAgP0ltbJUry2sh40V3h0+q2eE6XTjMdOlHcQh/
mE/3RCWW7kYu3nL7OD2XzmsxpMycSXW1UZJuCD/o+7MKU3UTeYfvb8vx0ltznp066t0QlEL6VvAJ
zY0GqQ2cu2k3TDBwHvI2XcXBPlsc6/jwAfKAIp93++fOOTaby+QZQj9sffhxZcsG0NCo4H9yERl6
+Bo31HbERdpPB7yh4WtFGBeEnrxd02FGZ/WlTr3Re05vLhH0uUcf3DTtr9ZXtGo+QhNVEinOQS8A
VGy6WMvtPfoRenMyrIrY8PXvU8tUeaYiJZanWQVEFZKcS4PY0FQ7KcfkYT82UZBoHPHrO9ubmnAj
23Xmsslf97CCdVRWwLvsVOJtJCXRIAJMAFWOAQnVzdVvots5VWnNyTDgCGJmfpFyKo2sopk3DB3J
3240xNMtQqgVqpNiKEOuUMfbR6Oa+8VMVRiu+RQez92095JUPXyccm+pYQF9sYryYnAbTu4etELn
yT+luUQXM0PK3IKUdT69TOIqxzbVeEUo8wJ42xvifYPF1Y/MiWO5UCzB21rJ2aW8j7oz/2UkfjZ1
/flLHn8SGSUcPMqP07zUBJV7L3UR5MRA1r8kdLxd4h2V80rMewctLXb3zUaawkeeiTY4eRykIovK
3CPGS/gm1vB9EqbZBI3C31YmBBySUafKKx2cjLJ+SSkUcB7oDCzHFF9j110ELlvM8tL7e+9uSJTa
87FSpHdlniZaBftF8GsIZJiAd5YZgzyYXeDBO5vWKeLIfDMhWkq9UA+gJyrXmAR4561iJKJaX4JE
C7R6aLbZN0n55g5HlDHumyfC7k0yqwGt77LKruPZ71Sgr+eQqLEwXhBowfnbKKpH3ebzBoM1elz8
i4Fzyhp3tI2Jy6g21uP9KPdAbGcMNl50rO0gSIohLaMrJEkHS4xi2koN7ITdIVS/dJo7xYnatxS/
8GBWxu+A6Ckc1NIojzwFy2Ve+5D46ZIf4Bm6zgxKaNZON73kTUMXJddVz0mq81/21ie+Sw3N3rlY
/Svw19Mu0a7fQiRU2OBz3TqfK3NtqmRPzq/2As5vScMX9zx5g9B67k/0mYM8gQW9SYxDqdCYfaFJ
7KJF6GTwwlH9kwAv3rbqbAUZb4lCoRdVgzLNfS8voOLLGRTqeftE/uXJfdTZe8S+DAUEuUlWlwbn
uT1GZ1kA4JsDD3MALeUnfSECyadPkw1FP8meFiiL20eZgIFEiBf0az5KhGecjWoU6aA1FSxy1qGw
96wm0y65lMOYRBUhYLoYxURgSDa6UkAkaZhvmHWd55qVAUB9ztyvYnPEXt3iKKk5hhM9voshqTbY
gIAep4hEj+qwYtrrM+hx2JulyH11+RYr8tyxMB+z6UDlJT9sbCue3xDifRd1rXIrBN1BXRr194FP
vGX59vMMXlN6VMnmxzL3lTURkFqsLSU8vXE9p7hADzFiV6lX0ixN1jPDPYJhxJeldDDHDcsJ2JIE
DTJ374lzyAD4JqFZ1P6hgpsWSiylzn5sAnX5GWJkqoSno4RvllkzDQhvDcNl1hsAt7l9GB9d/2rS
GvnXmv7zUww7hsJQh9CbySQ9fesuIGzuQXm3IWgcWmcTPCfILUbYNUNXr85KZRvD2J5cT1v01xON
ke0lhWexyXjDXbW9BKCxd9yT9qKJfvMiarJXthXfJQajiy+LTuoBuzcgEnl5r/7X+vgaMBqG5epB
WJiCTn2mL9/VouNDgOg7IoaiKhSMDDtQPR/T/pVyX2amqbg/TJ8KlZ1o/Z1JN8oI9iUMvAgY+zgS
dtU00vhNxAjZQ/qlYiwbb2DLVpxE4hH0whB63M3a3f4EoJEpW2UOeQJZ/hJCnjTFDJbTInR5Ixel
1MiUdgiyFsme+F+JJAV/UVzAihJbRmwwxO7iUPQssdIcxbMHfW3uPTluRATVwyEZs/MhrRVaQPgc
I3whlpF1zURsnHiPVuPJI06uUTiseLwD4bFCHRPWb5ekZFwWK7561oey8h7fOtb1WwFTjNIyzXm4
2P2edrF3A9Pv2jAMQy0Ej1FvyYAbsTjQ1+7O4LuIwAhu5iHaENMZUehhmTKIaHjTq4ce78O3dTFa
G0GWAYbFsBkqPBfhKrbT3yLbUbc6+ScBm0fXsdSTAlDziOuiJ+8iytw5WHaoTBacmSvEPVlDRcWU
2zhVJx6gdfjl35WWQtNu240ds9oO2TDaIbVSHmlis7kDQSd7QKIGK3w46N3X/QU5B9B8A7X0P15v
mnN5XsWR8R94f1mRJZuv8A+z3ecbFE5XwpymtB/Vba1XNe36EMhifK3Ed7bc3k68tNTQ5X7IJhNI
FTBT7Az6Gg80pHeqtFwWMgj5YmNLKaCsncuRwmLJvbWJw0xoY2Kr5jn9gU2wYvHNqOYq9mJ2jmEu
7KgdzyvsR81KjvDS7HN0HrN7ZampZS9WdHZC3hojeS/nF2t+ExnzpquPv5Hztjc9S7XMVn10H0Tr
o3yKCHE0M4bdwlt3iGKiKpz4ykYiIj+1ECeW12Go0HDZODpAH+ULrlIp+n9kradOEYIlPYDfsfSt
++cfKF4ZDYO2dB7QCGOHBjfjRdMj94UNWN+f6YCAfWS+t0vLX6t3wug3uZ4hwggFxVvwI8NtKML+
G8SNHZYIT0HWbzk5FU5pa8L+FjS78YOXf1bRpHUiCv6BDokWYZ+IvG8Kldt+YLIgXDrvqi4UDRvZ
WxhY3fd3Wv1NV3XljJeBzQAUjkYskrEClBb7imQn1Rt8Nm3oh3tI05gWS2BJlljyW6ou8U4HR5Cz
NA7qLOx5sM3tuXERCZF27Y/69eh1b/1QhsROYZIxIwyWY+5jCEaH6ccUb4v/bQrz6z37ULt5bVEm
CzkfFpanLDAI/i/ySHEgirFRqN730eYnCY44XdB67vH4m3fpaBZ3aobyH23BxPPfz6dpDMEQVEAk
jyTdQzE5ENDzyukQ1Lrd1C2/AmaoRr2qsH99XQOg+jtKSpLgfgvG8kXHpdASjkAYvxWHwQhu/KP3
cz+D2ZNPYKRwDpcJhGih+sg39dFMACIt8oosMRHp1IBh0xUQ25SPvk6BfD9MHN7vagoONEMmY6KA
Jty3JL731ShG5NQqpxDvdtWHq71pFpe2dotpmtcj3F3GHiffwM7PV/XMdF+HrfeXxp4rRh/bDTfx
+eShzvqMrpfbcwQqKSVvRq49nJFi+5AxVI1gNMcTc+UOwWvBGk0uyVoDACGr2jfJ8MElaB/8r/iQ
3f0ZwEHQqhP0/Xy5wt5eBLUwuem4urXJ0mBjfxrZNI2Bcx2fJxR7Mc/bRBgOwGrcfUo7qnofMNUU
YIpsRiKGGxXocqf3H7bvadGCLIRMOUol73e9rzgdwbNBo8pvnqqAa8Tb/3Oy9Nlr27MPqMbfrkow
mFqe6qSZLaRWFmVFtXn2hDNLvz9JEcux6UP5COfrWbI9naYFJvkPK4m8sw65BsGEarSyK3SCjwmd
/oBiA/PcI7PwyhGAtBk5Dc9vSHqcSEwb3PukaNt/Ko6Db4RBo3QxS711CtLQ/dDP+KNnJCGEZh/T
sKRU0X/Y1KO1w2OTMVVA0rwZIPNfEvQ6CWM5M8oGPtM4kAo3ACI8QHBLHYrFwFcwg11HZVxn0kAg
CqqWCtAdE8qPSyPZxXNJHF5Uk094FdVs9OD7+O/H51g5os+LmLR17CwbmAF/LXnV+191U+XeMoVy
n8HiliF3QnQN5/cw1L7zyJMkIyv6dWCHWJyd+jQ5itSFMTR+tvF7MgtsclGcBg2cccQmNmmoYm9H
RjImtHh9KcwESJhHZyvufHp0z4wYvlfCc8k/inA+1ztJtAY0lX5WKTSDG7rB/YdY9yfCm9HRPpDm
tl0ID1vNqOXAYuR6CNnMZ4l62Xqk+Ajh+Yle8ZcZcNQC7pBV8lLHaTQ89RaMCHGW1nWlwmXiFsWb
NDk317ymyB8LRUTInTWnWMTf9SFBKGg0dMf/3PCAgnfHJ7c5Lu91uF+wig1JF5iGnPgT52ldRv9k
3XzP0asuspuLFe/Tx+u7PSOD/fkztcuFNSRSd17SkrMZRu0fH9Kl3Srsoiq70uE2oRtqDms4px8U
PES69nrhwB8t79w25u66HznQMLd3ihrnyQ+od+7JBmzmT4OF/cRRxRBY3QpvMR7XJeY9PXkRBBC/
BS+nfzqpIpiKdUM4/j1hjR5zeAFqZKZYveqBRyvTj26o2vIS9GjX0XlLNnmUPju3B9Y/IZ6aF9Tw
a9h/syUp/XfSK7u5pQ5KH/SeZipVCuFJtl0nls/8fT1YfPpyN1T/jIoP9pC7ikZoFioTviLeq3CK
tSuOegWdJ25nGr0Y5yn4hVGvX2a1QboY6iL7ATt1LfVeiaUXQ8FcY86lfHD7JPLHCE8PMRuXD1Y0
9J89KpP5nILUk8BkQeYYT03r0TJ+/u8Di5zDxc5WxeB2WxByMHy38nEwJy2N4FosTB83Yv6zI4Yu
w6Sl6qIy6qK1MzQCgThaCsHkfGN1Ek8O4ffcipEgUV1mEl7/EoqZ6dN77VIt2F3I3g2C5/4Y6T/s
OZMnxBVINqEJFSjMKZ8IQS5423EX2BilyozitVJcTvWG+IjzagzUVFIuCCDARZJBpl5U/geC+RrF
WvX9ogQhXSktYZsIJEWqmhpKwz+QmJz8xszPJNhNtFRvo8i1wE4LRtKTwVDNn+Ul9FPV4Djufnuu
7Kair/tyccLPZqeQMYd1bH0NuvzFlHJCpx1J9Auw07ctQe+AOBQK3qWaaEvMqQu9U4fhRSc4Wh1B
zRaMMZ4RN71it6DY+eytx95Yspgn8dS4mWyRpJ2YM1FzgGGc4iNsEex1i2kJZeISBLKoy/+wAoCV
8DobSoutqclBvIhA1kG0VGE37BvGYs2WthM+pZSlnyoBrkBsraWeeBCTBNSF2NnEnkQX75ey4sLt
ZGZgoHIPYsi/C//qKTGX3evHGq+yoXj5Wo8ME0CO/ubTtMR7fBLj8Z+Ryiy6wJwZYWFLptm5pefs
9oMuh3lSqP8h1l9UehfgbakEJNn/Ay88VWXPvf1QHzOChHHTKVymFB3JaUhAfyYdOwJu+1UDqlN+
yPSObMIjT9/HkiPecAsqzjpcOK2ukJbknx5Zj7dcBC7yv8xoia/tvoPEiWE+N95sIQZmxlLeaXkX
claeiS0J+EOMH+FkbmRTDmlYeuvEpESdnfEm5V+iwKxueNRZW1jp1Grpcu5Oe85rcTxIqgXt499J
MfZyyDkTxKLkRlZs/NPbetcLbStJ1ZRSoS0IBQQQw2lRDq4pz3iwFqj+v1d7z2P22JWaIiPfF1bE
IIpkEbNZiRqRhaq6rkW4t405B7ReMD3dDCTNAt/0kntcviv022FSnWLt6g+/T0XQSlIjfWZvWVx/
1rStFFBI10z0uepU8HBln3khIG+19w0bsxnEmcUmI5WKI0Tethe0Vr1XtzN5LXEDi5z7l/uAWwQJ
L7Ra/dQ/qyUX1nE6FkgpT7ey9R+VTAOCtg4nMDgXN0HGqhC20lU9IgzcnT8QtgUlAQq3/30HWqSx
pRBS7w7IWvIYiZfLoveckyLu8Egq1Wpw64ckedCKYbcKjT0uu54w5NO+tf/tZv2gqAhZ3/r0CpMH
XvgLfNGfmwwTTeRiABJuSFKg1OE4gKD30vNqd/ypnvzyenu9DwVEjka3s5RBZ5Ja4mKEAnMgmVeW
E/mBOSKNVjeyR3LUp7CbSbPf9/iABjrEKMlRHiq30zfg6dGiLrhRNAwsGYfe18cmG8FjWXK1i42E
s3F8DJlykJGO55njL+DPc7S4YYCwhjlj+JCA67NsNSs+PT9kWsCjKiCT3DZZ5yN2VJrthJlcbbP6
PhW1dvTL/8A6OBr+FXF/LMe2cP9NVa/5cVmcb+iq/q1jfe9XXxgnVBQXtGiAjrvS9lwT9A1SuRSR
n2tQGSjR7PtPy42QwRGAW5BgDvWHYsG8/pGtOCqfpG54jLkmr24X+UWtb+4EfbzL8buQr+zZwsaj
Cpf80FYcbSmBZlS+irDYlzQVVGyJ7Op0nz4LzrIuS3WOOIVwgBD8fxvzCfacTSmhs9wRkKKbOskR
h5dWNww019lRrlyiNfOlWhfCbi7yxXbzMb5RlSSNg/wi2cPZhBNRBO7neRdu3lznyKKvk7ZsoBSV
URhCPY1pfxNFgCXekt+KEeczX2TAEVA2VYlQ5RsfgXvgz974/Jvw4vztE0+uDNDOe3OaaQ46RmxX
AMhS+ILQaOd1dsAOjnouZ08nHo93hq8FnEPCnzkYDElJlazy/2n5vVwvsfTnrH1DOnsBUmMHQU/j
GTqXejxjwOx/1LxOM59yS1n3pUlDjP68wPoky0FdVuFdFB4zaQE+QGuiqClCNxYIi6ciV+aBHDj6
wUaQebFFsvRn36+k4tbaZAqs9mkc+uVky7OHg/NZX5B6+bjcguXQUqK4myIHh3bdSUBUOSjwmWN6
3y/acP1P4gh+IY2O/PgBy8ITTCmnE8Sokvy46e6S46GFQ3lPm9r5uz0GGIObvheOd4Fv5My9FJOd
ssE9gkFoufAjhOLsXGojIKMZp68A7eZG2Dl0xkeCwZMRFPHlAVZEs5c5nTYPX+q3gCS7KluPpU38
RZprFQLxWGqa3DVeGGgTKP1u1bGjuMMQ+DqH2hVjhq/9vsj7guFLlQ46lCVZP/TJSLJMZ918M9c8
X4kAGbgrLGkQsIwiyyxg6CaUCfwcQKKP9UDl0u0Nr0hlZrA1LONv+1qyDdLvyC7qXlwM1SInc9h3
s/8SaJer27NBXBmPHDNmTjQ7R3GR12PdhrWhtB+EF5eJ6qtndByYXgh498LMBp9VzDhRhnfJGfu+
uLYwI4OQPNyb52AXIoc9vg4MKvrN8pgRcINsrZ/ZCslvwGDiVnGnKhHJCA0UWghfZxuW4i9mFQ39
uuv/k3ZsZ8pC+i0EVL5PzTd7Ol2LYB7ddwkatlGDMxV6xTbqXrPZWA3nBvEber2vSjH58izZSgqO
4WTMfIMnsFWY+E6h9B9lMIjpv+gWE6mLCCF9rjhd5z3N0sG1oH+2gSN3KGgUDR7QzWYwhkAwfNNg
mCaTrr5CW8QlE1q44pqkgpbEzoVEgJ0xSWL3jfJEl5xpXFkJehKK04GtXjao9JqDa+A+xbwJ3AZL
GeUzqURweAPxoHB0O+R+eVU6KR9qAv9o6+RWP/U6yJrkQxkFneoyrE8TMGcSIk4O+dufbQ/VOP8N
i+LDRpDS1pk80rjj65otYgLRHcl4ppNKwRSSn2eAceFVjb9b03Qi6CmFvjUIcILIIL/ifTDn19qC
b99nSMFbw/ceEViwBPVE5KJdOIE7pZ+AZlAqRCKmGQYnWbQTV7oTslDGv5rnqMV1RiMfY4bdBLbv
k4rDDjY9/Fypm2mfRPYttHqUYldLNks9qQeH5ZQfkxrjjCXGPfmB/RA1Y4fLaH13RMEifdI3kHOZ
XaXIyW0o7PUJIfjBFYguzEORFiHgqILaxHeYygAEpHk1e31gBfxKrk7D/EI/obt8ne0nQi/ctHbx
dbz/XxHLPCtPsRoLin9j/CpWEKhH+a3ghgLGLw6jS+p8w86ulCXSgrGS5IrVjiSuuAbIA9X7RFz+
Iowgaq7ffuNJdvi/fMx9pwhU8nXE3V0JprTmu5B8oqrVHQPrOBw7asMRyPL6DvGoOUlohNQXR7jQ
lHPzfuv2+p3nC8PqpN2aaTPATGQCOWnRwhztlJItAaW9hUtBapS6sCdvR13QiqMxsakqPe47rsNJ
1jgMjlQO2VNhOofVRb9J3ZyojRziT0CTAOZiNdyd5CQaeRWTToevVXOlsnL4b94bQHdBatLGoYsc
1in1FoL4uYNJtUibc7pnSFBCRguIHFyjLM034r6/1W8ZJPGFVK8H7ea7t3smdTuvZSk7Ei//cuYE
PABobDUGfO5Tv5B88hXcp55dcUv6ZmvcKACf5JbWBzhndHlMTZiVLRi1JThAuIHDahWYsyRdaRz+
puTT7mYpuKK9ivJPRovsOABnMa0sMgsLZwyMGo/izxT1XZ9tlvBOXw4Msfk7d8QzokI8Fsj7Kf7w
djAmswxiwKIp1mFFFDFN5sF27h9nd/Q85cx76sczzWr84YH3VTkFb8vfPkn4cvpBma4yK2Ci6Xf7
u87ER497RTbzvr2gw4PaNKIzoNnYPF2uA2oz38u9PnRidUmoV524QSyC2kj5/MWpQCXnB+xsYHIh
1PjxMPK8Sxzj4yzAcPyg/Fn+acaxSIAvjtzhX5TPJexYuUJe8Fwgam5Yeip8+ctfXsCIPpyYzFVZ
t5V21jBwcI6B2UeghDVkA+6kr3M602fIktVLx4qaP6g8ox70/AIWic67Ad87VBtScd8uGkGOPS29
85qy2axRPL3kbcLlOzkRBntmsUc96DZQ01cO6iYfHVVV3IMB37X7LRJzbM6vxZQ9CNyVUqxmB+YL
MtYU3WI2OJNA4UF1si9qAQvSI73c/5zlCWk5Vw/N6RUKLCyV+xcEdsgGrqUiNh9R09FugYiSq4vS
wPj1ZD0uai8vBssADAXEWEJReges1tNeiISwSzStwgb39OYZfaahBA5XtiKLi4Srewr3tr+uphgj
PO0M+m1xUL7x0EnCx/O52p5L5H3jGFVs7pLNRdF8HgFHTLcvlggvz0obYykpPuPpOeyIcdjBg3EU
8wZb7nwci6mHbMVXjYpLP2oM/ZDo5nbstP+ixKbCzK4lzDrh91vzT4sXu36TUQN8vVTbZCvqWfNC
WVkUS9LoEai/mZ8coLoeeYmtUcph2lWd2TcW9GTlhakcI5XQ7d/W21jh07+ShrrxbdEAIVPrQYd1
vbU6QfbN48FDukFz4codO/BM11SBF8HMDwmNwgxvcjAF3OmQVmM7gfrncEAGushXEe2igGCDVi9z
s2OAJ44E6gUCLIM0pJiLHWZ3/6ygPuwo8zgkzYfKmF1Jpqk+z0Zf39t9hd+gu2I8RW6EmR/LurK1
BR0SJmd9Grkt4JufFe2UoMjJQXhQQ216CUPoDZnl54udUmyDkLk2a3rOlNjiXyITSNhVbmFT6WYJ
a+OQ/CPeqcZ8K/c3bIVFGI7YK1xhKqDeB8YKdNA9mz2JVCWCqt/m9xn7QZEUmcf7gJrwdzTRHMBg
NFFbb97v21tysQW27vuMOA29tZiwXGtvF0PGWL7VEs3cjDjsuHlg/I71dDZjVx4JEvKSMrzg/5+d
Y5y2hsQOfxdbsmSdBwSmyE/K5eo1caf/7akYqpq7bvDmghhQ7qOCCUM1Sxxr/dbbNY0CWLq0vEHl
Sc5tpfHfO+6KMRb3j1kDsWs9InLFWLZE60cgoMv9b0N6kSI2IMUm9ukSsX0CB43+MPWDW6zcX0+s
ZguehvY8gjgC6Ug5Ni8HESXIoBNaiHjphAMtR8Z5KoAKr+PV85Fd/iCGKzmpcw7euZOGZLYD/qrH
nLj7LPyDfRduUtL1skniBNXunDdVhW96z7jQHF4EYmHz3oX4JD6yFXiZfI7spLOvSSat+jbUseMj
9lKumb16snGOpLHotBAy/xyBg1voEzjQJqFDeayIxc2kI1hUKCfZyBurhUOY9B9IJjmkghjLA2oa
9VHwmwliI1NbZO9GG0mQ5lWnAPxiJ4mIc6A+yIl89xQjTfMKWHv78Z6g16Sgbsjy3piW2Ae14Rwn
mkU9ojQqzPOpF090xtLiibyyErXnTJtE5Qo7b6Z2s2KaXAjfE59N9/YAyQaAQUNr3gzGMMaubCre
GoX7PtTnkGPuTEvcLK0Ip6TnsWo4xKyTD6utVD1foZeg648Y1Cuh97S4jTpEqdDFrAMIMpptliSs
A03B2srq9FOMf1+U2q17Un4jiqVSPO59VctFdQi2YUboRu9Wn6AmSZ84GytzkroW2ok6GQiq/7Y+
qjbZsGG0V3TPh7mYGBBadYYHFUjrl4rTpIjYCHgFphkhHg9ZFMMNThhzIcTq/MZoVX2CvqolFITT
9Zgo2eT8Ptzz+1CVzRUw/aE/x+7UpoeK61SckOARoWBvsHHb+dFNRhYUCfvAi9f8/jTJUBhHPwi5
nH2D1pWnmxGYyYCTimK+G9fHf9Fss0nZaRzVwzJzkVdFPc0z8WXXvsB3cbdqaRqfwhri0GA7Z7x9
oKWcnuFnkWiUC2vC5k5fJ15IlqgqF6GCpU+3hsPDcTNArxDCSgq/f6efu3yaNN9VL9qqDzQ4GL35
u2G+yz8yCIJz0RDRtVk1PJgNfrB1ZRN3DRiPWYoJpp/uQG3kweUjBBpBe97XwV5oJhP0uK46JfSe
V7iUxUIgu8qBByi93m21X6L1/uRBmGnd1bUBNccshnjuv8bdXwSYKosEHuaovzjzKHGSuWsvbvF/
7wZA8u+LgeZfQsgm72ZyFmbhA+W7iLAWpAl5prigMZBIUFtYdorNF7HyiM2YjKhOSjIieXPslPyF
id9/52wkVKJgDeAvHXlh4A9TX64Cv/AW2DlQMLRdi5HmlSiqD4QTFGUA5tRsLYA2cKo6fDIPnVXh
iT98x02NuQuyQghIV+JgLrlVMn7SqhynkVBetGKqxJ69mSpvJMMNqWkTOet/sAjhCB49UAuBu65B
HyGyVKm1+IbHX0XaBjtFCxSi+71xz+jIsXpHr5wzsJmbQZrV2RWnLGC6dk8I0vCUUeL8tUh7nsA4
YHE1pMV6UpLmmMz/waR3cdP77ldkjVfGGz9HM3X3YASKf7TywFmk+kL3MYWeRJZjOGMa/ZZ4JFis
TnW6MTBNZs/ngooMa6bVhDdpTuXZRZF6m7ioltyt0x+SRp6iC3/eClF0fpif/y5gvzjt+AX1w5o7
PzMQIehXHpcd+hpaZplkRLluEVTTxRYNJV1Q15p7eKRvO+Vb4SXAVDa0XItOhvH/3zLWxksXFhnS
1b0n1bAcK0/qR/vxDJTD6qtFuhCr46TMQouGp9asVIeXSCXcoIaw5rV52jRNiccmwVyIlX3S70gU
eXCRupl8aFOi32N6G8wbBGW+beIrvuFiBX9tCdbDSf79PxZD9F+b9pEkAqgy2x8jZVdBxRhzyS5+
sdjCjyT/mJOX4+rhn1tZM8vTBZCJBkCXtpCI+gZ9wdYH2Qdnef7vBIJyYRYq0+4uhKs+X+RS5WcH
Ja3chihAGK5aWUHgd95v0W7kMQiXLyqwmIvG7hwYfaqaQ42YYLk1aW9IzLblaF/wA17WcmNgYpTM
wK4xu6b/6P04kp+buiZkU2Y0Jw4QuIxeVEl/+WZbpvG7sL+vqT9tiEDMLbWYikVVR5hmOuJOYUM7
LPZSvymwWjwcXXdFyAZetK35yBacQiSioMvOMTWYznq67IIM8oZVeIYYYUrwyBL7qySdxoZh7Tea
b6FGkdBlbb0ZGXT/g5HnacYFNWx2xjfCSLqLFh0yvhPGwpexIbtCmqYGCuSKsOJ94KxgNnsG18nu
+Vmmvcjg+e+5Za6lM+Ixbp8HrZdZcTTweRLIXSIaEay4Tqbp39CioZHnh14EK3wjSRRRRwQT+NmV
ngepKGPZOSNUI27r7TTODho/T5BO530/doY/dK/DyXmzq204eze9wwoNHTd7/ae60icKBKFpnZZb
YcLoc3nigtMb0pdsxY9LtdA30AtUnE8s3o8/WuyEQBL0kMCNtV8cYmjQ1ma6t7zjWQCOysD/IgH/
MoIZe2VB/1tHZuAylth6Yyr7Oawi9pJTGyTdhoCswLkJpGIVLxEBXhsmwXT0ckeFB0WeeztKLei1
Xv3gZ+yJPccWprsqxBrNA47x35/yQutMaTShTNwMHNm6pDnql6LZDpdo8Yf2IOP5v+AFCWrZ37FX
t5PrciwrfLXEX/ZZUajJxuEp1xrhI9hc+uOQBZw8IUuHNy/oMYrQ9qhR1izyvgIW0dPX+BWKJISQ
yXpQYSFh3CkZW0TSLjQws/dnklj7OyGj5VI02mr61Zv92G4R0PiQqe7aHQ8LDMc8omt2BAYFgsnr
w4cGlLGq98oo+3BkJUcQqY2xDSU4IYK4D799QW5+n8mCnBTGSvYlXm5dVn8mf+lAuEOhPKXEoA1a
PR5CpW2kxG22B0vJ8WiNDIppDeRHwKe1xBqkN3/4BSwfpqJrtpoYrAFsAomFNNyNYKQVOw9nY+bP
iC6tdsxeAYbIwV0yekDFxm0iVTpPLX28oGztxzv0bRGZdBnztBSLfahSN+lfWzJSxjSR7scGmsKE
PZKCoo2LHVeCQQcR2nEShPR+uSzwVAMH8k5mtN09DxXtqr9go89tohS9p39ou48WDb2h7VEaNRiM
2H01HrEfUVfyP/ZqTpmjeb8OM3Q56yEFY/bhrpdKMcURe2gczpxGGnUFR/f6x0qg6y6uE2T49Rt4
5HBS+SAJ0uiAeeBJFk11+QuutyTR1q1ObBH2K4uRTw8tDquDfwR/8/4vOVMtDQ/oL4lV1uUgmYeR
OgzX1E4VLEdkIdQoTYUPWQR4IuvWuNTgTXgAvlTRQylaxV75yDUBJ+ThcrzF0hwiIoIkqats0U/l
LNcJS3U6CsjJjq0qxYOM73KdeLCwaya0cLTb6LPajlUh9ncnusWJ8JYUlnXCPhyVT8FMKCAaxWyq
dJ2pz85IbCHcQFwXwrAXRYvTpOtjYG2k/GLXxkY5kSWe0Mjl8Wg/Wr82+gPHzs0CPePdw3F4ku6i
xRjcxgAwJ2hJiGe2tuDM6LIOYESNkA9kTp4PXDYWUGuvS7tqAWJWOtqU1nERhLk4LH05Ry7+/hAF
dS9V7qwJygS9I1gnTDRpBDWBjWms1FYdcZDneOUrAK23L9k68z83dIMTPwW4uH+4t9jApnboI3kF
RAeU2ppjDc6hTB6/8EHM1YWF9x7WPA/TGRna1fLedDhwzsc5VPvZ+VD4BgenNs7Yf0BnyFtpyUsx
SDbfIv/d2z0MV69A+hdqAVxWYFN92IrhJJ1GR7gahg33Th8uEJgfw20HyKDlU2wYCXQtcMVGvJXq
/SLQJZydH5zMXJ12ahlJH0k1pzHhOTLhtWn9tMoOVxmY6TNfrB/xJIWMCbXM/c3xBcFNxElRs9Np
FxJ0AVMMEhfzTlo25rHQrINSzgmRnoQZfTXH/FWgSD5QBqoOzdQAOF/quxDLb04rbQcHLiijokM3
0XGDPqrvLTuJBCU+Mmj3zeNvWkKEwRsEK68ZGMWc0NxMQfzq5awFDrQH5pRKljiv0RhnSxUU4MUc
tgLfaYmaWg0TrIZvqv1c5QLh2zSnCM/XqhTxxW2zWiBv9YZAqHHEvPQJ1Al3ih6vhHShq6Jrx/sV
icTvFbgb7Sg3WgXKphILzrq+Vmm+tznXMdDW0PuEtxCpmEwGAjH83BVZbxtqgO9qkhJBIv9dfrjH
mM+vNNbi6FkVvMPwsL5Q79L6LNi3bwKMxuddt1vstmgDTTp0lsAlNkDjPa2DzWpSgtQUMdfrfsWO
erXBZbwfIkb4p1YSxD1PcjUziLWfTNnhz1YrBzX/lc0CAToRyyLY3HEgf3XL7mMHlUAeElbNr8cF
ZyP38qhyPWnBj1IOlORLdCAOUFRZLifUIKTbpyN26kPhViKEs1k95SfLd7oZZb3u1hNnUOMD5LNE
GZswk0nymzoxOCg1E7wWDyGvP93nFtk6Y1vxRWlJWXZ6YgEg675xlsCDCMvD0JYGiOor/PDTTyxe
VIjSilISDU/1vUoXQzSw0rO0iMa5BCAVSKDPnbirYYHm0lZPtH1g3Uc45axe6MsddGvp2yEY4GA9
YvHbREyCJ6u1q0m5pRVU09HQvMdBKenZWrdvGx5BYXAhsE4pJN7Y0oMKQWgpUOSckyJLivqhCxkF
SP1JFIeBqEH3XstsPBNt3M2lrY34WIJyIi8dk76BDUdNuKpnGP/eHjosNxBY0Y6UwjQDaSApTrKO
EN7l5AWtFKYWCAawSk+1F6QTjlMkprOw6OxrkuAoArEuPpZAziFJF2lb9w4vpKWTz1n0r2UBsNno
Jhei6aPRtOV7t4UA+aCJIPQ6vL91FBdeBI+GL0fRD4KdmvYeCnRHFctuKQP6hnTGU6B1njB9wCgT
Cv4IJTNiL9lIJQ2oJgVMgfCvNQSWemwl+pke+igBYwvSKtM2VjDIIcXPtslsKyeWDCHmLDbZrX8i
owKvkyYs4z35JRZM8P9OAG2uj8mVmnSWLk6JdMM4ss9fexRb3KwezfxOh4jF5ngpvNbUFWeACynF
JnncFD6CKq3Ug1DhtkUI300VLOUtyoatAUCyykUohzVBdJVubFgX4/h9hY30DlF18AlFobvOW08j
kdWGgoFWwk9/1+NoC5Hv+GKlQMRj9AG/cDTzTQcgCNi8JdXXEMQqnU3LVSaVmuUgB/woS5PNEeq9
09UIktporcf2AwOFl/TrSR/1ggKJ0QesNqr3isNWYORjXm23v6G0NI8m1kM9JcFPvZs5zqvNv3Wl
ij6WLApKOAVdbRWU+9x7wthPx2KBOsdISNSDT62oC/b4PISJyVay4fWzX6dxkmjfhH+2ADrlicZ0
njOwcG1CbA8VYhK3CbDP3MQ9LkH2Ykh5vEf0jidm3q14uXz7RhCw4J3tepMokbNtosFtxFo6P1cV
F1cTNBPFRWs02y2nDeDrYdjRcVaExaqc0CUP5g8RL6wgK3HkFZrMW1/2/JjwvbJxaVEu1QzwLwaD
P0pySYrjoSrNPqA7gGP6g1DZPOh2Hkg9zY7/JOOzG+j9Iwxf871DXhIqESxifYWD3EAb4X6Pwjo3
2euXohikitKI0ZTel6wFbFcvs2MKiqJOx2VixsXjzw0iVktfIUBxZnHjRA12tFTHgUagT2ZHJzzI
15shcFrNv/FjcMU3M/X1sHqxlIUjoa1Kxn3PWXzr5JtNXZqYnCzplbOZ7wkZBTvWr+iYRiVgTs4H
B0+H4XlPPrajTgDYvtyFW6I1Daex+UFQefl1cBPL03TjFTsn2mJRkiAGuI78CzlSPBCdX6RvpJqc
SE1vx7TGGb/xbmuXbL2/TugKeiVmjwgUeyAzKCMGgqg2A+qutRSf+SGETZHMOtguCNECRxWDHlwk
L9ERR79omK9gXTtZfOkCFUmmO4mo6AN4avUSll6VryysFwu2FQRnfL7VUbgbzUQJmLNn3jlvAesf
31eVvPqDQ91IsyvkYuTZkyHH1I88DanQ4oT9PnW6I1ojLPcNrTe/zEf1JmZ6khGg1t4+skiUBA+9
GnjzhunVbnsIe8opLQCMEcS6SxUp/h8nxa18h4a6Mls84XdmXnG8svI2JprJ5FmCMFYFcFKTBsRE
qjt8IogBggsHH26Hm0bD021IVc8VgOpjbGU2k1GuvwSZLKz5ipXjOxEKcCN33kltesyTN7VxW6x6
P+rf9AxxfP8YSDd1MrkjIqnn0ifCkfaDr525BcSJbk772qtPH5caVAjCUfrx8mFK8ZU1yshKg3R/
vQWc7mujklwjyrmn2z9FEc0AnJ+kONj0tUqafuUbtNpgDQxdxCLze1EpzAFq8V3PzZsoKrN9fE21
yZexWciTslaN4DH2yzlBReE6dfsiHnvkqmszfSrJ98G3eUh7fys5rlZGQMW/ReocrwfgptWqrEHG
EMsX5XzsYXjCGe6UOEaQTHnG/bFwE3ChxMlplFlwPwgMKtistfjMvJ/ULFT65NaJXCCMtLKntSNm
fKA8u+0iVbLR3V+8gjmwWoj22HbiyeIVJ1GKUoeXfDi4dZgRYgo2V626+7eK41NCMEel2qEQqNvP
iSIrYJz2TYYqMcVbpFtjXEduMiePliF8/HJq19UcDb2wFk+Xszpt3A+t5YhPl6gEMbKpBHuO4Kii
cTeLU1Wffa18iDX1Rwb8iJTvd892MInugD0p/fDPE/+tb/edtLOqB9Zv1E9acRsLYFh/aXfGyvX+
mJVHeQZIA/roQ/Gv9Yay2itqrUtTy6crj01y8SokPpdNLz+2J3+zC0ncc5dKNDoEl0YzscWEfivH
jVpow/5DSeIwQyjBSyiPOJ1K/Ir3+3zhqOrpgExlHN47H8MGhqInTqXxtvsLnVcUWrIXRCfLojnR
P0v0hyKadHIiI7K8qm5Dmgs2Ur5ZrgjqO1lz7MykFjdJWtgOIuGsCKyCLkpp6ofhay/wVlZKcmVT
fb/4kMqtt3SD1ZzpwIAAfJuJiJRMfdvrMhc2u3ldm6w4TEhe/K+z/l6OdyDU7CBwTG66JbyPOmun
7h4nVa/O1Yv9T4kyZlsrgm4HIEIOLTgww4wzrN2lm2wrj2z7zRkIOl8wJcbyjj0oCu16vxAO8Fa3
sdZ1AWbOYDGDC3n1+SAc2Z/GMLhcx9LmKzuTvtOQH7+XCtiL9Y/diVTljIKiVUFn4gRzfscpprpn
KE25VFLUd4/4AKAXaqO/YPjCMzPZY5oBcFH3pLe/BRx+dsr8ZbihaEeGfo/TID4RNZMIFaVmCq2H
a1SIIzyN/pkjTnw1M5h3bFWvSkR97qW0sRLaEN+cZQsQWNWnKz3aGcOv65JJkBMCmwSeiXjtfmlN
OpSVNUbsImQd+0g0xd2fdzZ+1wEBWr9etagiPlyKJTRw9HzDCg7LJFIXAHok7gZMyQiThtKp+tJa
hP8FXcE+DJE05A5H8QHbORbx2Y5p9gECr3A0s7OuFTkTI6EOhNOdZRb/Ekv87pTFeI9llf7fWobM
dNqwHjeK/7aWUhWnh6xJInwuqgL44o/42F82AvHPtouA6LHmLmoQOs1P4HS+AirGCioG+5u5E+MU
z4I0fGES5WNUhoZI1yTWmVKCKUvx4GIOAfOwxu6tYfTv3jNMKYI9pjmpCGPUO+iuvXh6qj1+Bqpy
x6JQPle8wsLkq0gel1P9tHcJ+wTzscx0ur8wWInQvwtp6/zcB6520r+9tiusYGe9tUqNHnWUQjjj
DW4NopJUBtagLAmLt2TX+zfn5DItjknA1GysOVnCJFA1hNXoMkDDXoIFmpfPqE8HkqM0sbkMXX9v
TamlqJnlawu08stezfV+dClhq55qNaidW2eP8m0SAC2rL5rw8S9KrLei8odB/oKwekpZo/qX/DaN
hVy4gj2W6SETHHdD4lWnXRkrJJXco0MJdTqm9F8pFsspzEYYrtPCl2O1IICzqdsxYcBO+oWSrYyc
vXfv8DQZuAts+orm95E/gUa8vkh2TPHyb5jwNDqSV0yrW8IlA+jueWhBSxZ8iGCoCW5gpPwI969r
O07FlWUQhcemN7E3ZCAOk5okYOQX37M/kmdcCV5GgN6Q1xVYlA5Xcc+PzOOjTtsirGg65c06odGo
x7UaHQKyw831nFiDYgNO3fod8ITiaMG8ddd4w3L65lUJSXkLZ5t6/GRp2amGhviWNLQRFB+fyFjE
jYBFDWC3uSFyjp6cCii47dA93EcjE0z78m3txJhZA/5Xq6AQhwWkJ5FNEMUF0s3eMG10dT20GpJV
Vgxm3jjCLrWHBdQ7LGYuR1V/pxWsxf6d4lB0VAahfI6ON5wjyBhOfrRrZBUpiipMcF8jwBWKt5A2
bTXYf3JEQ5raEsAaNkVd1G7bD1gj+sPCWJPN4XylfjIqNiFjFOwL0ed2LY8U5INlBGGuEdyOa/CY
qRZCDW+BumJRRGCiqiKMIP2LfEYloEs61z6eD1CrnimPG3JRduulI15mPU764TYF+HcZySu37lHO
JYkjkd4m4vfw/zMj8TqpTsmANDsyHTxmqPTQUzs3H9UXW58D0alrJkVA8kfbZBJH1MQx3WIIRYzq
+vYPmnxaNzQAcHyI7h5H+bUMSRJuFauj6PzsT5YO8bTw0PHF6VJfxn9c3YEyzf5k3YwA1FrOO1Zz
ctrCIWCNgDOqpie8b3gwDWpbphPkm1BvqPTQr3BU+wHi/hVjQ78g2BWfA1N8Qy7jdov0VN/BhXuP
ZqVWVTZ+qm6/hUq8fxxtPBfT/4Qx6KiOhvE/zy17HsJUcb3B8dIud31VYf1P6uuQsRdV92kBx48c
glCr6IjNp2jyb/1FKDJcnLIkjYcewnijncmQAZlaAne8eQGeGGKXHj1+XedmGUnvuAjykVKOOk2g
5P+Fy13eUs/P1nU/8CxJxVwPr45cHtCZQrgpKJPptsrJMn8qVWNXUbxLzO0u/DVp06MEQayVTo7F
c22H2SavVXP7ia8ybe6TrXaD9XkpP1niYcZrflbRfGd9dhkZuf4yoxo6b/z3iBovfw8FOjeMKwJp
SSUlHMUQRFPakrPiCigAgsdjtXBnPvcpAvsLN+8och/qAbTbXfWyfxjvLuyUcxecze5nx2Yg2Abq
5E8iBDHOOaw+eNgGpHMPR7UJ4upkIJmaiVUM/g7gErijWp6faS6nf5DOU/YHfzpMSC/YNEZBJgM9
BDt0802zOYltKVUrR1cLn02HyrY8lLNYhReJMK9HiUOl+bF1ASMdCl4sbK7N6cpZfjoZPkdGHzTd
yBGdLrCfV02P0RsFKQrsJImn1l4tWbVxco3SUpuING57Ubd7+3HpaHnt+uNUe4t0qRjEHq6B6o/X
F5iBUJftj51HKr10Cru0rcTN+oDYaYl5MHEJKHpUpSxHUBS75BOn1aaIYsxdRu4antQT9DF5LL7V
89zwCOVwasnKZXOZBihsHvg3cahZdBQLs0N59MfaCj5+VNY98J/Uj2wDFMkx2ufGXRe6R44LYJbj
LaXshC0zZ32OhAHBFYwjHbKdg/Ikai/fXfrhiFw0yB34b26SureRreft6mo+p4AlKDyQjdM9SFR7
RK5S7eU30tMDozyZymjT5Sa9stWkuJkRdpMLchITr+0aKxr1SkYVdY2pcpj6AvBauH8F0siEV1F7
qPyJ/xxURtOpYOmh3L/oAMqvX+YTBUCGwltKcNohWv1AKM/8c6IYWYsielGX0dtlmkM/QFgavoLb
0Pnr6npECV5cIPnZnWU4EUV6CHs0cJhwQmezXAdH208kC2EWw4iHth9PUWD2gHM5z24Kinz8G0gf
k3HV8DyJBFpwzbcG465hju7Qa4Dp/+or+vrF2pn6MnOOwdR1cPNuDsIS4wMD/xJw5fHhBamfQDUK
zfdBG/YjG2vAkBczoVy348xmoN2ZWky8QQyut3ETNt0k/5vj0YmTNlb8mFXfL5wZ8amgUMIrafec
8c4rTLahF+iYPfJOwAtbcoW4fkIpotIi0Erq4+1JUQjQHmaVxGKyGn+RS9hV6NiXOPvK0p+/mzCt
Av1q4p9BQpzA3NvDSYBuo1z9PR20RdWAGNXDnvUfXBZIbWI4hY8sZzG5aRO+uBRuy0WJ0O9Qwbbz
yhikvDhklmVQXk9GIv+rSLU3i4MjpAgQ4inYw0fm1ydtIBAOjOrfGrryYYUethw7jy31ZTClf8Ll
jnWls9RDPhvlfLrJtRjhYFdMWivHixnk+VE5esn4kH/cJkI+HlyU7+ggIVbe9Ke6yR6Qt/ysoa1d
gBKhb5LhnHvOZF3LoM75CtGRTdEt6b/t6JF678KxQvdnBkn13Xs7nkf++XBC8tD74XamoViTZ9mm
Y8DupKKeVJ7Uodg+8Al7fTXg9tf1K+AWepFDZdQep3LvS6W2pNOVpiqaA+IhzL6n7msSBDIuVGVb
FG6rOsfN8rOlZqc3pNvk6QXCHAzBOJXSRUbDOmZTJYXV+fpnXIS+yN1HOS8arr4D7ETvnpL/Obns
6uAEPonIDt3XXl+dZ+8jRCHcQaDf3aGnCA1egq7+O7p0PtPhKON4ewCBbt/NUz3mTvg3ItAEo9nn
683yQjWgAzbjky+FkT3OVSlo13Y+hO/Tk1wS+SunBwgAQkw7W8CQtuuOkq+mulAGwy1Jx+c7sntJ
EcOwcW9bXAqyXLtrvxb44yr9FX6AmJ3BrTGB6r+O7OAbQUvWY9cIZ6133nN2OgJ8GnW5wE41pAdG
YK+KYJzs5GDWYtKMc6mN6zklPjdzqIxFBHbAS6bG+C72HsCZj6tecTrgYV36rkkbdDhqTJg/d/iX
QP7joCsjD4GfFGV4mElbcCk87wA6k0cERhV6010Sr+zKH5bAkEnLODGCvgu9mBhRmGZZZ23I3Qp1
Gawz9RpO54fujolphTo/o2CoX7AllnVWb43a/5e6ocB7T5Iyau4KFQQ0QJwcF8qK7ErS7GtanSq8
efTwpsHHBTkmMP50Hq3V1fIMrBE4Npf9JKDbERy9nhkPqIz/IQoClIGOBMt7QLJO+HwQCfeORjxr
o7dSPV1iyayDejY7fTF5UFeqrcNQ+Brj/DnS7ApoYlD3Ge2YfHAgDCtpcd2rLKCe49FI4jfQL42S
FYQ/Snw+c+559DdMPku4+AARgc/uDyuzbamKg3fkstPncc8HcyDCR7vqow7PVF3Kj0/G71qByLzi
pEhRq20sMMXQM5RKucJaXiMcjxnYFRyiYQXnMnbFf8DzAZYYHVnXmRrtZhM/O3eashmyXGp8N8Hu
zG98QOpmQ3a2iKXvAadSc/M93GqVUDdEC6FbuIbVmw135Vh9mnK7u52AjsO6UoxCKcoORr9f1x5H
OoRDR7LOuaSYfpfNfSbbuDkytzJNRFhc6buZgaIUjL1eOnYKB9JRifHu7htx1e7RARQIvp8C0QyO
bTeoGffcOCdhnuvM8naT9nB4MJ9AAuEcj+p/CvkeEp7RW9Ko7XWIdY+aStUE6FJ56TODsKT8p3bq
EQ85RcCZNs8zxP1bXLDyYPo1kkH3sDezkoMAj/0lZF8hCn02/efCHAETDpFRO1xtOQJnGRwgYVwl
XZ2YK6qcskDfMy1b+9vOvXg8aOyaj/J948K96rjvVHGJdroZ24gmNf+J/REOiwp3jXyAq7RoA8LN
TH2mJj9nCNEw72MaP7fxSiklehUZPS/llvRJvQDD9ozn69Sj5lA983X2pyWHKUflp8fM3dXgp9QH
zsDm7iiuWtJw0IdIP91/V+/QuJGKTNvluh8RSXKkf9UzjqbP5l69Mfg7q1eX/Aj0oD55az+kG1Jd
CO9GYjTEBywcVxf4xWL/thcrmN6OsMBadNbuB3hPXBJP4Oz+m9/3BH9SEqg2fQWlj3mu2FayEhwS
JVlnO9Rgpx+YOfGXE3LR06/mYMsVINK4EUB4PhvLALYVs1lb//jTuPTNmPbkZ91cWMLCxvAaVsDw
fDkdYdc1jUU0xBz8DrBdZ5kHD8JsQGLKUlfuyHPZejUc75lZKDTNpBGDq27tbaoSmYgUauZg6c3E
/R7gsSjl8p4oRRnGem4qtR1eB92Xk1ObDY8yrPy6FGxdYrM9QMRlyoJBZ/djwgexkoz6kx+v0H6H
shucfKV24lk5Erb/2koHdNDfVh8m5D3MKhNufJ/4VRfLIo2SsCW15SFFgAHxOHmB2cDqz0w/9vmR
UUm+uDR1h2YgzZ0f2vx1i4GX8a+FVuNjU+7zAwKr3AJatAnnZoDWpHJHz8tF0+FU6dATu4qZxfpz
F0+CZj0fahLIHGwqioevti8O9G1gyxiCHP3a7To6FOpCE+MuwzPHzfSpqPA/JKIrI6grYPZ2fk1C
Cdl7rlASB9ZfpT6TqdeKU8On8eETzpl3twHG73ea0QMCkSw70z44wZsYIZj6ITa2OdnVhTZODWQH
IczCsUu96sb+ZoykUWolB5BqFSkfiF9OKtMX3CzUacihq98WlzxestNnOunkq5bw0WJWMACdWwKF
pgKsv2iI+BAbfVE06zQAKC13JCf7teCkBuuGHsJ3+gANQ7Z7s3MUJiuew7xg+sqsNdKfEj2UNiKj
i5jdWv/EZu/uk4KsI7p+BzP7NLcHoC3Zs4omjH5ymJNrLWddpGXK8660JwFCCleXcHhp8bVtplr9
4DbZv8vs7YJHDsJYCHe6NWgo/Sle/QYuvB+PSWIJZ639lJddruuRYNCF6TOscUvYKeLj9bvCQ5eL
KNf8XQcGZUcELyuKZUjev/TIdoYUiHco9ZsUYM865mVDj3Ou+Dt0eP3JPBFvvV672wOUIM384s2E
LubuNhxcN+Wx3zAtXDMC6pxZvgrXByzw3m2wDRQ8t+/9VCbgVxlA7YNL44pV4wtyCupHJHk68eaH
bpcGKZhGlr9bqKuRCHTH19m+23fkQW9UJR8bbFN0pcrNOQLT/Dt2ymVOY0yNHdMXpf640zvC/gQJ
VNyS05jXar1P5rciyk4YL+Yn+cyey1+/plfmSGFed02uF23skOwganoVl9V/Hq1KeFttHX4TZ+dv
EI3fQm5cbtsGjNFN+nkSaVOX8L9mO4J/rs1aro8Du0WF1Kx+ORhY92enUmFmGegRCbyMT3srGsaV
RQA4qWRYGsMIqkzsrm8QW6AZ9Lg51mhXUOOp6GpVx/RbqSi2qxMP60LIHxhxutE2SalLkW04J3Za
j/0sMNFpoRGzrthOx7arUfgl841SutFV98LxNLUqEFFGSKaxl5ZrCKbvvlwVQVUhZietV7dX/204
UZq+h+ERoYXNmS/cBUT5mw7jNG7OxmOy0Mn/0bT3tS8IbymHEb2DCQhGUuHqPDrkBPZTG1g4b129
SjSy2PWYtaN++SCMqPa3pZFux0nnuv2Yxlz9AlPwKRvFovpc8Uuf3DhfXB1yHWtz5O1gz8fLBvNt
LTDOZaKxtX5SPwgHPbyf6spvhfTMyqlKUiX2ebGS6Ommx8/UeXrgjB7Vgasoj5uWFpjT4zdqeSEW
mSUEgjHE2glYlIRTXbYuh5xAaXzNWU/EO9HK/Rr6Ke4sPVRD3umw7MQAHMgwu9LoEdTLcEkDpk18
0Gv98fHuND64Vmcg25M/bUGC/t5gKN0fo9tKZtie60rJzTIufdNhtqsBzg82icErYGuTglLMJvsR
AU5pynrRqqij7ZzxNVnUNH5AMMcyR3rMZ6KO3Bhr9GRmuzpHC/h+kSNR0Ov/V5erzIgv/IsnkoSe
835RxHpbvETJtXC5Vlb/Hp3DSmiJ2Klln25CDtcmkjMDGQL46ArTd8pxDztJYUdLsxbiZql2UGtI
i88/QtD07tcIrFFK4lkS3bLmJ8G2QLzjHDLfG7znl4LuS0P0ojI1ujdAiuVhlnswK4igwAiIoDc7
NmwhKpSjSqBUUU+Hus0XOWJ6mJjAyEdddzWw72iKHbDvPXsOFmxn2z6GRLy9HHi/6xThsEr4jKZH
+zB3xZBJNYMHbI0UN4IXVpk8B9X5rld2AMcVl0USZu0vH9ehYPWvyn7MQpv1qe9TwsxZ2W+Bz2hD
sEY4FhGxfJ6EbYM+/MJNUXDSN9r7XwqJgxX/0WUWhfKv4UOsKq9I6ZaQHSH48H2sze7eGNagtyrx
GuY/JyDKyhQJlZc1DVaZ3ToIWlQ/iRpDpiWomlG5i7XGDM/sccUdEqfze6ut975O76D9YfNRSsRW
hO88ZbZAHnHsUvaYxD2HN0N1b5otsyjqrlOLyApZJYWQ5tvB5tZVdicqe0oKpMpdyJJqvPXFAWBs
M/czyyH1KEHExoaoYT4G54TwLYeV6J2YmLiXDNFfjzxbhhekTGB/1awjt9oxj0CZH20I/dXIhaah
AKqQVgPqkhuvC0+gFev7rtd9Zrp1amhNdXzQn+LTX8cPG0dz9y6Q/CEwJOPYKfKqS/xtzAmTRE9C
r996KOIZgwzuhMRqFfX0poVaFwCEZxxl5gTSijHBk8Jv78PRczHEDs0ChvUMgfj8tNbwEcjhy8Vi
du2cp6LxgtEB/xSlr4BdnOCNdKhsLKq2ikK7w6d++g/5I2KTj6kvLdAWRiQgZaEiZMKkid8/+/Fr
30dXROlUifgfqqrd2/7VC4haV9znMtm5V+sNqUWt5gQ4+OSlhoyVTL0902JKv86NisaYtDAC1Vmf
F1lK3Qhc7N5wmmpzLjSdmY+NxDow+AxcpwLxs49N+2Tg/oMxEw75FkbSgiB4pMcoDGKKiQuLwb5/
w3AJIree7bo8aYax7zdBtdY5jxjCZcFi0LA2hZOixRN9pp9cQgvKesiu558nQrybOtmeezQK/nEa
W7Ck0r3WbfaFbnCwDQz2fYzrF368Drt4Qc5jXDuJ/z4YpFM0ETyetjt7im+kDqJVv+TGbZ+YRT+w
etYnQ/lGwe7oQHwpo0+gDwu9TpJ7v5IcZMA8s8To3RqTHfv4aLi+0iW6LWpSeWy0AIzzPBv4In1h
fB4A7Awif7H/y7tY3VuEr8TYlsVnrBPY1pFGRF1srtepZs8NpTJh6NgBhKxVCISqhjXaQprSo2a2
cpSCnSkP3hw/5MLJTdtDnexIv4amcHgMcszFtdGH7DGCc2JEvdv0X2nKun+NyHSMGUQgoNWBTpLa
P8TEa4bsRh6CMUQqjMIa8J89AOpeMlvT+5EIhRFk2yOh3F4+11Qt52fKVj//8XrRQbz64LoQieuE
nuUFY4kI1NbtHjgAsDp1JTXHT+4ydXC1oJbqTHDFx3TkdvK54jugUFExFcc+4On3GirBA8dQDx4F
1gh+y8/45KMnXehNYJj5D3UrpfcNy3SQjeEqmMTn9lE42iXDwiLqq66jG50HumTcNohlLOBPvAcG
RYLcwOA0bpEznB3/Z6+bGqAaDtqCX3Q4CMcR2DkUPBGf3hr0wcq17KDItspH5LBRyE7aTd3FbCP8
wpv2epdXiX8zadK08qmjSYM+Ij9jJwmAVITkAuA/43A36DHrZ98bspeydt8d+6unpZCeazU6aWDq
vBvQoB2qtLMuFyux2bbAWtZq4htrBQ7Iq8/px9hG9a/kTr7s6M1kyoXC5ZXWtwihD2uguiPoFqoL
yuacEK2hWkpZ1njRYdswd9GzucFxB6eCBtqRNyZ2WX/i5NOJ8PIynK9WaxghHWx0Zg4/5xYR/s3z
ooZwzoGC4BpZ3P3ZuIaD1KWqdyq676pXXKy92mS4p764FO/2QjoO8MHsc/s2EiZO5iwfEQITqy++
sGN7dBHpPOlmXoWqrMgBvmH0d1VCir3PoFz3w8Wm4awl//AHtTwiaXtRbanOUoFl7Y7bQjrsr4ko
lDQw/UGDLlBcBtB57Q0IU7Mm7xyizfYb97FA27VdS47ffbWVARr0p1HwVizd0O/L6s0lb0NnxAOp
fDDQQuGgfmd8FDbQFOzPi7TGRzKsyctvounBmizKsK4sMa2powyvAXcPXrJn+W+bufPwiCpSUjIU
lYe9HhsgQvNhiwM4lorsXHI3AnvcTrRS02myFshMbQiJbS+fqe6OdXkakayFFrfuZ9i4uDLMKdxW
SRmxUSLg1letH0iNvJ+rgHR8xbk9nmZAp5tiLzr5DEi02ptQdr3tHbID1a2LL+fVahsY85CovPwQ
3pb9vAMuEyHsRZywT9BYDR99HjM4HbLh+mltd/bKhAss5ecpANAZ741EmnRLRoRiKJ5hXx8x2KtJ
7sw+898bzwcO59vBioAvGmD1p2tucGZG91MJD3C2b52gZ3UCx/Y6iG+5aDlxlOb/gcluZ4X+tJPW
5hMQBRoYjzkUr2rjnbj6gfuxjwKnteNRnWZdvr7ozjANxHDJgbes8o3pucuiLm+uACfnNOBPHXKg
3rO2Hhef5fvOJecXKfCyb2DGyd6SVxqqkBBPJOf9/CSHMuo5xD96iPCWA1zByqhuSQo+zCkNkG2p
cmujV0vAVvgt9IjP25ZF1K/mF+OI9A5CPl/HE9AbH4ozVbwAUZmgaqdANZ0r/LwZlpshJS/j5oRF
Ew+DSN3ETM9BL9g0vU8j5aAm8FEY31RUYiRioC/M6YbtR1frm7y78/0xnQLUu3KEZqa8X+Y0uG1z
PBVVrzZ6kqJm9tm58HO9nrIWZlJkIWhdv+EKSIHkjmLmBM0U87+Y/ULsuFadWiMgJ8Oe0PMhDwc+
W6hj1WU1oGbC/GrsbdRhCUSGpDJowBrqAIYpVOfyqcvr3OgzUWHxVuBHuZoLpyeWQe2BindzUCiG
D4BBxGR7Txa+ZSenEbcuXPSfow7pcI+rvcLtQPvn7n1qwwaFuRcoIWn9a3m4IU1zm6yIukag1mCW
aQTKcNErLfbu5jzaOD8VvheTEojsZwEUoZSCaaLBn2HD6/W0MW6jqXILG+ZOpqlyuIdNM+gAsxZY
6cNL+/uqrHTGQ/RonzP5fVArbKG1D5PY2bJprsPGTD9kXedVGX2WPGjIIU3K0tU8zT5f9IYa1G3A
MQXYPtfpy12SHz2vbqiK8vm09NTbZ8+IXVA0+vs1mJpJc4D8lGuFP8MJwIoGmMN4PKio4AK8JgHp
pDMA+wIU8Gj7YT2v9gh1Y07h4wL7YLty4XRaFthGOJ42CephqhGN1HJhhQ9VCff0CY9e4zWqAjrB
AyybfYm9D6ks+/x6+ZVe3/oYA5Ln8MjQCFbXT3zpgune3cdbQVCdr1R0XJX/dZyIO57B6jgWyJ13
rdsrM9gxd+i1xcOUQVP5A5TopPr++0vFGjxQNZpDEior0KP45Ack7uyZmghQEqT/CtUI+gpfZhgP
6hV0xDioIMG42IwhvPRMf1DJoT538wulgnRwdHDA+KsU/iSEhWJAph35mYi7/3Bm0aE9kbAYTIKr
3Wf7EGOIiOghy4MpnZjKng+JexyTRz74ocoaIespPyCnSIGdPYogjXGvQYdqAeTB1oRj5vrJhAYl
dO6zWWNQPrhxpbricY5qzth0iqb6dKL/yGLaVq6D4fJakqfwIV3DpYDdtqci5C2I7qjAMUeevmCu
T/rplyDWr31W2zmm+cbxM/49tT3LuPifqNrzaJktmcqgoL3RdZp+1ybEH5V7jzCCCguLpI51fjlP
WiwSxZmlu0anEt8Mi8ebNLhI1uxXpH66di929AjPw7T8H1lEC+BGjLKQYUkzdkMTXXUSXz/xIBt1
oeKcaZBFZJtp0uwk5bTOrUxgKXYke1hPMrXCOy52SOwIIGxWvw9ks/41XMO+Di+zO8QZ3rJSbDa6
kCm1BRCMKQfVRu9w9UM/4Q1u4itLOFIVlOOjlfZv0SCc6viqH8Vx8Dmcw/kmKQFRuSOoge4ktOYE
JeFCpXXKc/l8m2J36ZaBQJG7OXQeXIk/mgSJ8U1TGKbhPDGPMd6iBNWBTnWvA1/Q9IvldbpEsBMA
B08w62B52MqXdaFMbGNMa6kKccrMZwsBE51sXErkOXNGvzlgAZmoDunYNMqvPRjS9w3sO8B+0mhk
IGgo5oRnuY7kRZ9GqCCpu4dpTaREmR9gmScABwwGmcBelHCXyFK4V/5k02UhhfBSUJ1MhxpmCkb2
2N1zCh/NLP4oBC+xR+LJdGtssZqdc/JcmSSwbrfANhOTphpyRSz3jPvPWiujitH6nz6FWck6oVWb
/sPJWtHLaLZfbOIWqa2+m3FzqM4xHp8H/vWaaXQXsNGnpDyj5X2zvgOdQsNjVetNVtL20ypIklnK
fhaX8D6YCDgi65CCBXsUnAhRgKZR4gP6dorzMPN8rbj70T7R+lxi7KhF1wW5ujJ3mW9LS+A6Y005
YIbkYwIVQZJ0Qo76qLihzjeKyXkvD3TQ3DPAu/xztEqLhGWp/9S0fivkfVvR/nlEtwNr7+gSqarY
T813BascBYAxYgINSeRCCIcMM4e9+wdbYHzHT6DTRiLjkpVGXCTfH1FbVO1SNdd2DEzsKsIJerXa
5MZhzPI3Ot3/eucWIyes8mTk+6kL/nhGaqa9SEwmy2G3Kkf30YWUyUzh5CdWYQWn3cJX4KNtUIoq
raqnTPncp3/HKqIKYGAsgNoeflk3/GVOe/VkfGrLbmv4sS0HeFMMW8wu2NzhsADg5E37/+3GqTUJ
/hfF8yzmAt1UbxlEC+i27CYZox+j65rLCHHxrOFyWjKxakkl4L0dqylDeVl1MbxFyzbaxUEATvrL
daWyMvwE/swxU9151XzxcLENZ5l6a/wfCzg9S74XfEagUxKGWeJyoEDn8vJco656k0yDu08wEd0s
0fyOUafO+ZWaDi//NW4XU+hJjpMxD/sdnfE5JvD9fVBwgBP/wHM+vUPIlwXiZESsx8HMXvJt7vsc
9EM+vwlrY61cG9We/tJNNCrDKZKzpPWg2WV70FFDuYuk4Zy+2Rh1eyFFnK6vxtaeKYMMHHRfSb3u
SBObXtwXgN9EjWnmvD6T1BdByb+3WBc/KQ5ILTQSZv/UzLhFqjuAy/S18iWvFvFJ4XdBrYbWOWYU
IiKEJUZJHzKn/rdrGmEF6jsaOGy5qOuU+Ca8gBRl1+qw/+3LjjfeNUnMsc9hfa1xrOMQWI3BjG3r
rwK+zTkAVgbkfpmg9WYMWlnDcBdt8IpSxXYFXh6DTMNSbZxseDwjuWeeYbOq/AePlDHm1iCEBBTe
kAOOqJXjTbzkC0QZH8tTJDTFuhHkV49djEfYed70JsqCna467zBpnP8lCt+M+fOFF60QfxGZy2X+
IDSyVRGgCmOs+aYDqdlnUL8qCrmUmzZ78XrwvfQDXJFTPayktaGPqXcFNbXJnQVPEL0qFR0RFgCT
ju4kEEunI8kvev0Jb/A9VFAwiix9LvwEgOH17gsslXssPmjrkCHOvs9ocL/WlVW89vZvDlcsSg8u
AvU9Hlija+pfv96SW+73ZGEAxtq7PJ3xTeNoO2gwbzmfX1oym6F9LUFJYc3ISfXzmgRfaseXjFEs
xpyrZvneYqYdLOM42nTlIcgkZIbvsS4EMifxjXI3ZlReZdx6TWq9tVr5tIKcu6I4xi4F8UkEwnQ+
TBnCXp2yw3uxPzcAHu4doEbgbrG0M0LHh4JTDGZlPmRtD/dJoBJynBJjNzr0iV6jh33GM6oSPJe6
yLj42mc3uIPzcmSEiN2wHtSwonNynuVWYMAkUwg90Tb4vTKhU/CgzN4YAQdxffdrtC7KhBhUPo2+
9R7bVEcpIWu7z01riYjJN9VjFJ+TP/pkgj3jYNmxOECN3UWHyAk21U3ubkZqcy2MvX7kzOv7XnJt
upBtQaUvjiDSiEht437gxng+BF+32QRiuShcwEyiPnTcsRtVZaKGq+ftW54UeyDMtnHkv6SbZ8XI
5vB+SiZRYO7Zch5fsEjiYnfgffSkiYgJ1xfmiIYbNyyPYDOKrIRA4tBFLS9gJ3mNXFj2hOnproQm
elJsYhJGpbeAR6PY2nI9/x8EWYV4ldanEXuAynCvf9pTQKPq4Wtyu1zV7fFebb0n4JuQDIWJPJDW
14pnySTjc5AULIpR4xIE2E4pwcsvfB3C6RtFajcTZZMu9yUSgAofQFCDQ25YPA1MkNnQ0Ocede1Y
iYj/HUpusEDF7KSp3X1YbmRcPkhOt7p5UMq4AVaWzc6k9o3YRKaShBBFLxpuEnNlrlC38xi5MAtD
/jUId7q7+gBahGCjQ1sP7JieLUpcEo8gQ/J/1ePNGRW/3v4QQLd20hBIz3Kwy6KWwje+XXl+fa9d
tC0i1ZD0ySLPT1/xhnzzRBCeaWqiPfAHzVr6fmL/FsfeiQ4EPJXYKhNuj+1xOHeyf10eI3WWYW7C
N0Ko0njvdrW+8Xej6c/ZYKBf1ckyZVa42JCStmoHRdZOR6ElR8pLC1xPosKMJBtxN/szMyOXHC2L
6JlG+049ZzexfrLtgLSH7NebYKyPQl07CLR2Ig317Kl+0Tma/5n3deom8C++IFanm6JLanlXWmMY
hVQ2kAk3qEKPimhCsMEdUN0bb2kXP+RxuJF9DEZfGWaKWYCvy1+4qV55ZHyz77pKGHQCk5tgJost
qwSQiQ3d25JBL0WXIqbh36rwN/jxyq4nbDJcl1TwIp6Hjycjxpn1Ui8gyr/48BwjTNLaaVySJ+Pa
AvLSNP+ta7c9efXdbxbuSSY+if6UcRh0OVKkYy+FxP4VHsskjHweZIqmX6SGDh9ek20lhUJI73QL
xFIMLWPkeHBp5OuioeiSxM6uYfIt00dxYYKdr+bDqSWO3Q1mpxA/6YKLtne1RL/gHWAOYdFgiXax
q0uW7xeeLBK97g1s97zTE8Wjoe4vucfkyf2O+HRLiIS4jjkhA4agSZsVtjxSLlySre4FWHeXOy48
mtz91tsz0dEC8r/zmM326rRZgJZNKEs4ICILA86ILi9PCokpnrlePTlfNH8dkYVOV20R6hQDPqyj
/7LHw+NLGC7qxEZQimZp6dHnVFQqjF18WkTcZBVYQ2OYpdeqbDXczLJ5q6LjDdhwP749vbaVtvji
SQOiEFPX0u+K2PBJUZdZUGmTUP0wOYWdK8Zc13RANCD/QqcJhaKMk6KuNA/IRjKa1sDrvX3HReom
bzSM4TeFJBiyGGcPUA+ycT+GLu26SJN6tJaUsq+e9xbhLp1CM0Zol5ZTeftxhMV1t326sLngMiq7
fHKeA0Y5H8VMtP69IQdb4SS2Pz6dvhdBpIxeq9CcIAmaIIN+oXCyf20lZ39sWQhyuyD5vPVcDOUs
1Zv+cFg/ODYaLiU6v2Fqti9IMAPCZiE8MFTnNSwOjCfIYk7HZxZiWORceJ977TLUDfV31UPDLLcE
E0GxEe0QOIDkToqF98ehSz/5ihG7b8pScxXqzniByCizflw5XegIIUeR69D1C2KgTpUXQIOilrKc
BrDYQadAIiQSYkMQn9JEw4byJur80rG6j82h4ONfHOhCMW6tnwz/yYBMyPpB4dX3YJgkbJ8XN8+l
VzsBUOFYwrZQ/shS6hZDL4FVc+e9ZJVzks3IR4Gw49LfvlscWLNZ2yX7mnWgWrXqbvLTJzSc2Oc/
a0S8cg+RINjqtqhXcIREDxSQrxSuk1txlMhhUHfvOgi6uEkcmsltJTPTd7YOXjlXcgKgiRtSH2Sb
83unbMqkTZT23v7qGLY5l8g8QIMh5Yuw8m5ettd07aFABuhAjSGlbsadNkddBz9J75/4JNCceE2a
TkEpyF0gkPlkTimA3LaT2AX+u9MLWbPYpPhWi0j1wfA8wELt1c3Ug2dc1ONAnsO+LE+vrJttbxU1
K8uAFMclPXAjJAyGFnniT2In70df2a7xjwSU57wRLtFriGpDs+xWB5bDQul+veuh3XBgz5WX3+F+
1wSxwdLjsVGBLokmJbTPEreai9KGvSfnEDpbgW43brnuw+nn8ghF+O3WdVS0FbXVRkIoZ+DpPTeV
/FSOgsGbiVS3Hh6vlgryU5GpHTtTtHctMbMcA6+fnqNIgIjcQC1iItg3xXodADzcLuz6B2vbmtyD
qshSlIoXGtzQusK3KHVIp9iMN9Yr6Ope2k/Dn0seQeFKmp4Bm3NbIP0mUcPfIbIlfUR7oeckfPYX
xiPFReAfR/7/5bN37MzaUhFnr2vhlAMvnDNNPoQdHXMBekKjES9w7KAfwuC5MrTbsw5SdaPZU4Ru
+X+jiXI+c4EL51vclREhDVg73sYMP27gHiqu6yNk1xK7D5XP/GG4LPI2T/r4Z69reZO3QkE9CIjR
+CPG2yMuRCj77NyHa8t5Z9UVLTOEzY2eMHJIvvOCj/5KuDCW9ggS+tDv+HI/kMv7NR61iKQ1R/lc
JeVxgT1/3fXJsjlxiuOJ/Vrg2DGf5Wny5an7PmVguokjlkLQkVv+Rge1fxyH4GywzcHx5B1Lq8Lr
KEadhN7ZObWobVpekCd3Bab9ScjZ9ikUbbuMgpZQoSSX0Eh6h2H5IZQoreOWCjW3SQnNrCwA9x1/
EIzA6C1vpi7vuTxUHyzMbtiCML4xPJiT/gzLy466uKZu7vKCFNpDzr2YFOET34HLb1mrzlTFmS8D
2ARIfLDN98nMJ7lOHNHoUe9KkmD0TjoBCM2Hn39WLYdxVTPJ/lUnu9zGmwS5EHunsA7wJOptlDug
lOHvZk2FCmxCxSbMCNTLXzd6TgQomTm7e7OMHDq/9kbWmuKLLTW7SGQjp/ymwif6PZgDMBF9L32l
xnVMJiORd5iIKLcXeTuPco+GfuTdMnY6bSWY116XEcMQZLIdK+wr3CKBW1u5j3lO+GkGlXBBxQYL
hF3kUPJPYWgw6MtwdfJrQDeqBYYYDrQjHkLN5xEfiNMQGimU65CDJRZHcX3Uux1p/gC5bnf09srn
YMoV22HHHKx0re7qkt3K9j5LN4PN2jq3LhPlSzEWtyx/CaTJpZ8kGn0+DoWXL4fjeuDm4NhHREjA
WTeX9nHyIhE0un2hTen4ujKYMmxE587PI7PEWP/oFVqZSeutUE+w0wEDwdjxPVJk39EzQlid8hTs
dDiM4vrNcPRNF3PRJsmjL/9rW+PJioPN8E1tTUALatbIhjD3wjcPoapJEpxrwx/x/yflDSff7tCX
b+b/v8rx6VsNudPqUDZzfuaQmLu48xYVnbE2iE7SBy129i7V0R/i//UNavesPHYW3zReRd4mXZPT
h8k0Cmk0FoTpMgTuiZGQtYj8ga5/BKebr/HVHf6iIlJIP2nsBm8HKaKmA3cOkBA9dZFQT94VJN8n
0ceCLqpMmcUK6BbsyBrMaIwZT8KFJXy1OHz6dZUJY+G6Nbog6w6sKMFPFztdJtUc5707MgvZaRFn
Iil1O1Acopty9qYXtdwVA6VoRg6CJ9DZIQKoRZjEOi6oWeRMOY+hWx+SsYhioi6ETyPcTF/RwhLV
bMePu070P5T7eUQhj4rIRdGnd5wBIcS2nWE75Fp9b4MsE0J2kzA16PSmz6q/ZO6sej8W19IPGETk
4CLCtI90FuKZ3EwZBJC/3St+uU467NvZFJNeL1Mv7MugutPKEkk9txkQJkxF0yoWItOCMMVywGYE
dYLFt6EZb4rHQw8Ghcig3y9xNiuKG7LsmuWKTiU9wgkhIPuLss9pdBY1UOIK5Fo5DHcCWFzT/Mha
+i0144aZhvYj9XiIXbGoIOHIGGVyshKKqYpN3ssR4KpQCV+OIk59pypvg7AINk7pwtvQ9zq1pu9O
madh55eyTmx3h0f11Fp30iQvLQMO96BFJKGMKRyUp8S9/2Nuwt8VqAmLcjojuwEILhFLIdap3a73
x3PSkMcA4AWotcRUfbkzUSuy0+c4W5F+Q5jJN5jLpUa5HHK5mQdLrC0paHQSgrS/sEthE9msCunS
41ywBh8fZUQtcVj0uSBx/ab5kwpGIk3wh7VT/IRBMO3UOo++QaDwWaDE6k2o0EjmV3A9Jcb6E0gz
jU3Ui65w6ZvfZbJG2M+QaDNzBitQRrlx3ddn97xdgxoIKjhdCDqreJtyQ6/0Cjtcm6jZZ+axmSxD
MwWhPWa4ovADvV0aHkWmhb/svv/7+M/BtWDgnGgiquRDEW3h5PSaEj3wNH2jF2jKNNB5E1tXgVE5
XfZJQAb2P5IKOCVPvoSvDa4HR4dHk0jd8EdCKem2omg+cyv2bcmil2+wa0yFVbCG5/imao30pwOT
HnvqL9iZ+LvisiaOFj/2KnXuKLrBpFKPuYRPsm54dE3IDLnfzrqTSqHXpjuGA6ZL5lbXMU7MgHqR
Hdz8ILxTP8e1jOKDBr5mpGBoSvvwZRTdZwZDcsFYOrNkOYoB8OtWoTce59yXuuhX7tNSMBkeYgA+
Pk9XJjSc9XJ607i9/4ryyriD5PmtY3XQKdFZJHeiTtlasa0fpn7UQC46b9vjReWwqTS2I4l6ot2o
L6TVcEJ5099Dhu01aO5HudjJBcJbtUrDyTprndjKYK7Z/VdJAIHkC00VylxUyjgWTLzgCA7vy5mM
hmRgK6tXTtjJOaLbyhoR83AzMUgeVNhKQ6NxR4OuzcW+L+g4dKcom6IymIY2gvSwHNty641Rs1J0
SMl6UHknHemU6X9bxG6T7sKlV+A9X31fGmSFrKPes+CyRleqOEZicaf8VAENSmDhkZUFgZHsvJx4
tf7c0Q0FfLEAtcgVfw3eA9n+1iFlbHiIJJt2YgFV2OWWKUzcUGV21ghF9UzynsotsLw7vMj7/08c
PFwvhthAhcVvdXAcUtWT4QYGe0NYPN02sVVkR3ckut36yfkp1NsOFNqiOj1enRmzx4X3HcwEqb/u
XFTbxXNpUwmCEdItn/Lkw8bdtxk6AcA3/5isQCgm+GvIZG7L7/kaVQrF7N7GGDYv/YUtMeppzCLW
8Ch8YIIGLs2f4yfF0Yft3mUDL8DpnoL9YxXJnBh7w5PE3ItSLwMuafdCZPavci67yG/AvlRj5lND
RiP+ZPDHRdIvqa/km1eDENQr/RnZIEWb8Rj8q2HU8KMUOoI3lypN+IGaBIR/SaKI7SzAUeF+/5C5
9GgBbZVH9ghuJfcITi9SGXalTnYlb6WxXG9ibjxkyVhzxz5gx9GKBQMK+kIRdKEOm44ROQXQG8tC
wpaviC+h0zan1nzawAfzQs7c0mQWVr/ZXB/S5jeQwWCQZw2AJaGYHQjEfv7Lv2y5w/1tm+8dYjtg
LXxKCBlxpW/pM+hg3xswT/rmpirnTzivvA0iAwlSo5Tyo6F8nh9qon2kslstR8W/NpppYZjCV55C
QC9FBWLSM8vOrQg4aPKvI77DLiWqA+lLy1jPyhz9JCMqLTJEMBJXFbWfQ0C/cv1jqRgBl46ryz7F
fxtuY2caOYp0ijFMpszr0H1tlpxr87ZwjVVRbmWb8ux9id94dtYC3putT99BEc4SsfvWg/SF8LhW
K+39N1zjZ0O+uJcku8ROM/9qeuCoqWhwVxvu8neY7TmLoXSJ/Kk1CWZEu/Jk7j3WUnqHuN2iy6du
br74ldZWifYmgyEyRhANC8cSbl8IZPuJ4p3d3JNoTBQpaNqmBpY9iAm4CLsJpa2RmqVxFTI60UZD
w+vs19iWhqRl5ADKNwY6mrC16EmNvy/cS/KxlHCG28rOwsoqyL9D8lJ/3oh6H9aS1Rl/TlFEswRW
AOUEhiWlOgsSSx9a+dh8PdtG1lBG0PR/YbJqQpQyZBi27sViv+yG4/OqxreUgSPao72McQDNIhEI
VjeH/z13jE8ib9d60F2g3QiZ6c0GmAz16lMWJckg8+IKqrIzDdTXmsaql9QymEelOeUWPDHH5EdS
98gMOtlYayXjSsXF5lmY7q35N2JDOJJggWxih5c3dOh/TouSFkuQ1Q1HFZdzwNIWAgA9JK/y9bv5
aLW3ctiZJQfJjhGoLqqEhaFG8Lep02mg/4f/e//5rlvtwwP+iSde4N2eBtvmT8R6XUktnbxAg1GH
GES+U4YqF2XPk3X0Lee7TDk8yF+553cv2Q+Ftkn6ppk1deWk7ErlLhxZSBsJk4WamD5bEyuXoH/U
bePkF9LnNzLAR9SJ20qWobBHlRh0lZZVa30V6K46vrrs1hgDefjZFLAyC9aADpAyRBcOEKZ86rQh
giMBCcelnN/TTbg3SDnXxBsAa4uh9zI/XhzWkrXu5usjSN9nnQOCmI1+0eNX/0iQq73N8UI+bm1N
yuOt8IrRwOblPlMlf3icO96a7uTC2km4wFK7/Gsw4WDkeTs1NDAmxo3pxX7VTkP7WhZHvvF/J91i
frz+C9W2TFkVizANEczsLfDkjxP55OsYL4Ij63JKA3VP4EI2/aXxDH9o6ahlcM1lEIzK7VHEnwJn
EEXkkh2E5QXmIBMVd/TaulZRzpAPtBuh19ENXH1AfDy39sKVaZjsNjvPGhm10dCR9pI5an6T/NPq
uWFpmBqzjZ5A4z8H4LX6f/yw/L8b/A761n1Bk2Z4naljb7VE5eYQeVeZpi7tcpifKvDpgFWZVB3S
L44ZHj5V6HTVEidW1WZi/8SezW1NalX76aK8RWNe9o1ggLZyflKXAfim0HRZ/5/IIvFQhmxlvG6K
22LJoZvrtrhmwpzvrhKK96ORvtsgINr86vPqqN3BkxDSE0XvpmZe/KP805LjA0NUA9apOU3MV/Qn
eo3eiVS8TRZtfbvYN/BUq26TvbX4NazcIXsMRNM=
`protect end_protected

