

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
BwHHaRYHij9TGTVh7NqyF6fPKvSJbz6zXpDQ9T0CSRjM0Tr3I2/EoB+qBgzPRFij4R1VpNLIhF/W
jnZk7ILw5g==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
EoffIvgX5Yh3KSkMHr6Fb+Y16CSwhqKyrZiel9vaFNUa3EtfX9ml680qKyH6k7Lt+GT7JeOZ8tsv
GeWg3Is5mnBMAsR5XkmKmU1Mf0hiU70CtdaVxbMu+l0K5NkyBzps5GWZFbpBi81xyWc3mZBrsdOP
SKFV3jiPDhzIXFusLNI=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
pC+fmAQpqkr0vqse1A8SFfJnAErWB2cTBoy5W2fu+Qfel2Cgg+f01SLqdiCqUwM3sdVOYKq280lw
0KlccFWeISj6EGy+UhrlckR4KPE0XJ2GFpTDwr6dIxS9OpYPDM1MXlxttLYJRqT3qA2yEzsidST6
0i31grVO6qNsjmpW2d7uByo9M65VEOheITjyvjEpcaFShH/Xo714T1rUj9u+HOahJ+Y/IZt5BXf5
ifgOOsFSC4Urhn+vw7WBdTykWaXAuPqSgZ+BAzkf1tn2a5qwxdC/nJyffVluJZjwqKsS2qOqxdcW
lV8I6VmHkVrsFF7Im+SIdtLtq6ajfsK+Fu41Qg==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
sjA1wOpImDpYBBRjnwY37zkJTSoQvS3OSqKSHwre5fBAKnkrgUJxozoTE8i2Z5d9g73A+Dh1Khan
8gYd3xbR7Bt78jJM+PFuUbVx7c2wSRcHOAp2KIXVLTpuc4ycdBn19YJhb2UIFhm80kkNGNgavUsF
mOqFyOQQiDU6WY7JVI8=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Yt106ecWVBUI4xOZZkRHweGkZD2nlI1jRN4H6Fzc3EkfIh+DLe1c/sY05LO26DhXbTC0r7f3V5kn
SKvkly14VHuR+p2mt2PXxY2kZUcL6SEF75Sdud7O3qeyYyxwzbLXhAk8rv8ESHYXdpJzGlAIPVhc
CV3MBlzutogOhAPHHcbRbukDx/ONHomfzueq+JuKHmbmSP3Sji52yPtcq4iLW/WcLghIBdR8EZ6j
UoWFDA94p9C7hEbP1WkZCFdBxukr8LSVfTsZyILoNCYLGaM4SAN+KSvY/r6FcDftOrSTK0VkVrNX
POMgLw4WpJ2xpIx+qCPH347wGbfYnUgOpgfHdQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 39232)
`protect data_block
E3AapY6Q87eJ6R6LMk65EgVVQ6vKvpy1Rn1eECzEi+ImXdVTW5BzbYmQcF+WGFAwfSK6oWnNVXdY
JPHtgUsfbWDEdkS/DctbQ5JDymE6FeSPBaYyFlbwTkc2fOil1qQoGA21NymmUvxMnMwFXVi2XIym
2ZHk5qxuGPUgWX6+W+Td/Pu49WJKmfDbCNhT+yaomxr6rgo5KvekguJQfqVugzNgW86My7oeHtX3
6V38fc7ymH66pG7oTJG4WRXGQQAnOFhpr2+gScnZjnkflNP3aESKq5YaMzdXQhk7ZCJqc44Fjv6y
aFz/4OJlxJMphIqheIO9H3eXyewc+byl46V446+qcmJ66mei1L76E30gRGcCCoqA2aGSddnWn5sM
3e4HG7aRGoaZuRwKYZEO0YaMmc+ld7/fJ5vmaI2VtC1LmstTiVHl8IXJO9tjq66iZL2+9hV610JD
RMVB7OSU5WinCXyZM23xfE/buDzznM3Mma5+aL7HqIMpUvzpHjhTHZXqh6JqvmPzoQ/Dnp39fHRU
Q0q4yQzyJe8Rikn2MyeGxRxxkBbBE3mIwCb61HON8YCNlLsaLtuQkfFy5/XP3+6z+kg0Q/bXjqNX
wraD/352Xew231MCQByx8mL8yLBdRxERoGbZWu0ZfdkNbo0/hcvDEz5btrRPEceHTzeUh26bc3xO
3Jze+3SNYjVr9C0t6H1KkqSmKDKjnDowEf+FS/xDIA9SJmhuC+pW2qRuY/Kt+M6+e/3ML/+h1s/y
b2IejbXrAUfDPRLFdzP6rSK7gewv8MSMKxQ6bu+NrCH7/rtMIJS940sO4NTZAm/+j3zmMsMPh4hG
fImH6Y5CBmjPyDb3xIAApG58y720r/sI5kPQqd+FwmDh/PeYEgmVFkqf7s/Yosp4zWOH94SckCSw
dVYpwUjGBwZ7s3cMW8Fw12XE6wdIiW1oXzp7hCNjJW7u5xy2K8QTiOTWj2yqrvpYtlT6qeWCd4je
nDuzp1Wk47kYtN3sAmIKeU0E7K/wurJ7BiIYblD9Ie9T7MZM1yWde2DIgxtnPCT+7EylhZbxEYPS
n75dRLmRPngW1E50J8gg+AJr6zOWNZnQv51EnfrVf7tDA7L4qSADDN7ymwy+y3lR8NyXqVK7cG3t
s/iYIJNEvpQ2y7L6LvobxDv+p04X5QW0rIZwDvSXtG0YFeu3/CXw1HdQxwSQ+zBCgyJqJ/Nhf3E2
JKRD4AZcVjFf+PYrIMmX3LAZTGWdGjBhTQjdKbZ4tNFMJ5fiJA+q7vd/9k+h15AXAk8cd/4BFGBp
YxDZw3DGiX4pwmJZEihziH4mEMIH9NJohSo5zS+MOL+OF9TWqQOr7t5pnFBamEASjI24ipqgQHis
sHInCWxIrCBznuEUrqj6fSE9NB+e6Fognm3fZtBon0rfqJBvLXwhFrxsEy+LIS9X/jP/xj3o+Cqu
g3dNiNcPYYTD5FgIpPAqymgAtQpkPlQRgRielYpqPanU5GKBDx1UbyPqcED3p1y3sLU8gsGNNT11
UegKrLeEpbO9VftKh4Kwi5t9lyaoG3Qw/JicdUZjdm5wJxLDtn9RS13zsUQTffGClZfua23eeV6/
+Cl9ldXLn3fWOVoosWL+dLfI6fNrNylQc9uzmyfL06X9F1TRAq++FhNDhUI1QqJFPFb/yYpwUzVU
nRYcNzA81e9pib57XWXGjTfCpGGKb8EuBM+QmdNkkKBePiEfwmYf+k4aCDT1M8L5c6B3peEJ0Bly
6e5dkxM789e/Sxc8tIzc95O/gAVCNdPq83nN50SjmcMl0lSQl8R9wnwH2MOAP8uEfdo6mIcKxznh
05sm4hE3wSzD8osc29CaXo3g0Se6pOYY6x/vfOfzqzBUnqUuSwcF5svoyMSGxblDsFoIIayMTI2l
I1fwLUoHtIy+9q/W3u7+boeZa5i3b9VQYAxDhm1E4zfOhNglf+RgeZGDdtfMnXHOLi24+VET+eNX
8tz1PJ75XOrdhhWx1RUqYPu6kyAO6BHOgnUtsraGFAqwofEFbMNt6YmVs206v8aKP9tqB7sFIok+
RBpykutQtLBW8Wto39jLAzC6GK8C/zbuhPsscQ3/XgVng5GEvXXcplQU1nu+rGa2qQb+W5xOg0sB
oH7jq/+NA22H0NJWbY6gm9EzreycM4d243x1X8Ra90SbltOvx0a9uMWqKhJh/97hLoHW91To/Q/j
w7b1ueLEGVZnlyZL95l35/974ppN+ItVSSARxIssTn3mC0aheEzq9rdD8EoZmFxYt2Tap3j7X2dl
zh6lups1KVAFaPdZ0g1+VabF5asDowrbTFaRrLNPR5HIJntzWBwXyW4SLAsR3TgrvenpzR5GHGVM
KuAQBExmYEK86PvKOW9YqBeWPSEOlinFZoZ9HD/2h9pbgjMiJROT8JXRiOGrbyq/tkoeijl1pTy9
wdPyY4/39dFaC1IiXdqXe/g23bPp6JlAl52lgtJdM6XOFi/PvOFcfIysQQEVKXj3vR8TP/dkLdsV
vBDE95p3mjHcrQURyTRU39MZkwd7ULrDlgF7XCs3rVWoBVu7gUVLpRCrbeAqJLR7bDRy1V3JJhEc
XF7oyjNTzfn7qWTslz5lNCa9U486owhE093wvRqPnbQNogr6h/6sl3oCpuksOCyILvTmC2a/+xwg
cAN3EqCp2oc7p833rESIwwbSeBfBi6/CVgir4X6d0q5Zz8YdUPDpXcAGiZzNaj8hYXir+MLs48bQ
owvIiCrH+h9zQMESw32Mxr+doi6fUNYvOFPMi0tZO0vpenReMndkSrZji+1vu8bxKcc773orfrL/
jkXkVRb3wL0hGp9kfZ6cR6sjbZ67QFCxb/hpBe9Pjqi6Xpm4VgRYgNR2PS0DE+v6FUNJZy1fz6Aw
kgZKGI6uEj3nuCpIvgVbtWvzXzEw9pZprmLb0IVbzKTi546r+xYhj4sllBwpfYpYRssofGKdHNz2
C9OBJeKYfN+KqlXAfbKNjACgU/Fi/7T3cWzaccpX28iOBz8e90n9fBOYGwFya6r2aJUO7hMBoLye
SyyHpDwqh9Q6h21gyxNHymYg/rwmlILaBrTyFZo/p21d9VFUZSTQqjOW0xWJttsvSZ9RftnobpPb
AgPw8ZTJu7bo0rE83tydKw7lAnrvh7FZi8Ml3Nw7DzoEgnnyN3YIYbdZ/CZ1D4XrFKB4ipZFjpLG
IITGjlb8j9eG+7QUZasv4gLFHsZND+I4nbAwgaa6gFOVP+sByP3VuncveeSHPB5F8c4O6XquFvWm
buKOwREdcXLx/cw26VDmoljdQ5NIrstlpA6FrNgDwxws8yR63BnN7IPOB14hwDmHIS/eUICVuTXZ
mlk4F/mSFnbQCCypT3PBAIeNw+aWF+r+XCdR/DCvv+ocJXHvO7nwQXzu8fbjtontcO91P/kC/248
m0AIS1XD52d8D+loXbaASiua1iH3NGsERVp4hF6j68ehe+FYBvZBLZIPCCBa1v69O1D02Z2hdAPb
0QlQ6sIk6W8tisFDLDJCn8tSL9qTJSWSr5SZHFJJjqBJolyPj9TwUHDGAf+7MS0Leijr/ypRpxH2
Y2ADTJSZt8KrviQg3tno/15i0+LYVnRcJxm/WnfCbQKwAzt2FURRipP+hoYnQreFL6Ho1b6xDwuY
1Bz6dY6GX7Xyn0Jw2yGwBq9h5VS0nr0zYVEymxuIPCX9ZFsOP6b4rU7mtxvFUkHF9QLwG5SMqUEk
EtOlk31mJq+jzdgZrK/QVcOscJ6ShbC5z8jpb7A14x0X/W0LmWgolJ8KI2YSkH2OPfzfC/eL6Bo+
L4AkHHq5bL1dMIfVwVKEE0sP3RF9GXrTKYz4BS5V1v7TYxDVu9HqA4GQFi6KLnSdCSSXWrQWcsTb
rgoCeGdw++DtnjYSeLEdeIYob9JUQeP9z0VJJVuSs7QMMJMcTNZaL2g22jI/Y/FPitpNEm4jcQ4g
YHppTkdVUp40W96OJmmRK0zuymqdtTAImTEE8/8vB8OI+kEzY9mvCAFJIq2UPmklJjfTYQCG0hE/
g3isNQoWhLpsF7eIPVfMlwAxqRF8JudkDjc5EQtQHv0p0RYY/ZrJHm33Mgyd5yYV660CFWiw2gCE
9dUxKYQKcee41R2IKxsxdVhPT6U2lw2YMVHbCkG8vk2axK6Oa8bydy86JwKQ2rENmGjOIGt4uqUo
fNQppHH2KTVgGAYhjWHi6HO3B7E8vTYfv+r2j1v1xx8u0tH6mX8kUkFSUoOwFfO2Cf8DodOnPHmY
3SIzOqDS4cypbZksYU7XVZMHZdLrYqv8N1s8LKM7LSuNZZGDC4sAygVZUA3J83rItbJjOkFHnyRU
GzPzXTt5X1zeM4Ten/kgEmNSZcxeOE5zq9DuGrDduzgEwjLtJHYNCn7gvD/RV7nIyUFn9LSGIvRb
+s6PYewGQ/LWHi2nwjkLfuXnMYZGIWTH/juftnIjX7fSBTI7YQtp0H9i1BkYvdqWbZMZp3Xi7lR+
SOIy9vly7hb/F5uKhMJkqAEcVBpmrIOowWszJY0prXGxen9cbVqWYFp1yaD8v1CrixyKPPJTrdNV
6s/gz2Fm7Mx8rZVVTR417HV1ITE9l+0TWhf0XN8IQSmoSX0D7MLzTbKUk44H3sneqKtLFiLZtIPA
y8VvGxQE2gGx21c378Gd6QuOcfus4P5sUQ9HlCOOAQobRXjFp3thSLgROGuUds8yfeqVEkJ9Dg+w
oqKMDpwqwFMIqTfwaciMR/cPUU7rcID3Ic4BVkqzNs3hy8MkNF3+haefBAVGD8DqVTa9pwhSvVau
pD+41O/r1tZuFzSahlenvpuaf71Eu0rU7CDYvXXpfszCI6XJrXt4NIibIsweaEJvqmZKjgDnSVXY
YvF6A0EHCahm32h9lkvBBzllahWiLyoWIJlfC/FVSYB+uvvyKFTkw+3C8hV1wBI3cCHCPXX3JwJf
/yFv34iEDqXAONkitrzvVijSDsM+oaegLZLKe2H8lCs/kbnp31FWhYO6TwlN2COzpeDrxRhIKRps
03elzkg8tEOKaeancgLHET5lOYrNdC13vbh4J5Sb9Myjery91RJCqmA8QGWkhj77erzWMDW7YEEE
xW2af3DX7GduoonhOAZS7nBEA+WsMPJsOZjZ7WeQ4AY57+RaLODMQL9YsJ6giUNqAy+Fq3B/F1Lp
YYClCv16Jgqzm012Cm6mBW+N1ZT1rMWP3HLz25YU9xEy7UvXiLNY4G7FObFQSPPlbnanxdHUPf7L
elFr4J22BoNvPS+qw9KRfFTFt3V8KQO0vujxKJXWqQSALHX+OPfG5P31TKPYnJe+CfxMfxeyb9Xj
GYZKsL58aAUrMPZNoSK10aBI67QuUGduWzqBSOuoZTudGs+KEFeiJXBXTvu5Cyjww4NtxqFydZ6W
FSV2swmtp4X8m8StXqtAELLCXI9ulEpnL6nLNFzCp/cNuj4NH7grsvUKJ9zwgmb6VhkyY4zT/6oS
9B0REkXtIUhMTJRso2alDO8kyO3SLvt4LgxM6RSLI9LZoYmTKhcrRySnJ3ExbkUXZ3VjLJXuAUjC
FStMpjqflSP0QUAPhnrf8FXLYekqFYeZXVr2lVa6P+33/ATBdOHZXHqP9Kw8mScsVkbvhaB6parw
eyaag/uOUC8fzEfxW+T5xDOA2k8ARhUWJuWGWE2xeiqXJms2GdFN4lFVYs/hosEZe/JOTOwYeDlh
6c+mI8KT3yK4vXRL8b3eumTyMWK/XBQLcrq/5lel9Jnsk943bXsImJ7TKumRUUVVR2NGTqavs4hr
sVhEAB0f3OaTP/sw53Ej3S97R0IOx9fGnWV4uhNQq7n/2qhWH4/s3tKKVreuWxInicrb+uaZJVWX
PfAo4VgWXhHENK5uLRNPepmr9L0I2DsOU4+sIjMySovvZXw/LLjrJVqLt4psWZvJHXIqwX+ZShyv
QtpftjTp2dCjJsOWwMtbebiA5GcWDwojb8xrm200WgIw3CAnXf8Y//5KR3KW8Jv7NPVexq6gPuhz
aX9I5ny2IWhETcoi0hPSFyx185qB9UXj2Um7KOgHV7ZqUT93EU1ELrfeE4k07mWW5P7JTQGCNZpQ
PI1o+lWxvTshLenfQ2Y/w9qCTZwcJ3J0vH5km1ZF/Nw6SQeeTAMfehMPVCWOWIh6lWI/VnlxTwlN
LIK4qm4ePINqfJVXQ9qGUvoaFKE5mWHDQJQiYpmN5b+C88Y4e5lVDxOhJZbh05nWUTira9iHkA1M
QPbVAzS8vvbl+1B9/lcq8cfsuR9oHdhsYhSfZkUKg2fnARqWPrbTn/Fm7TD1jYV1FxwNZSCXfJ/f
0rczr3gDc69QmvYnTZWQjshA+qHmTWkilSdUM1CpwKi/0q87SI62VxTljHuAE/iQM1tALhwzQVoH
WBz+fZWODlDz0bfzLZKZoen0Kdh3A5jARtt6c4uZPDdkAtUKRRdfcHR9Ro1Xc1TesJAm2B4b7XZ6
3d1jH1z5iQkugC61T4W5aO+ZVV63zB9D8lCaYMROuCLX5b/UjzcFIQ/3Kak5lduXmzV3GTD9j56R
qfnP1Pau/MUoMKmZFWODlX+hc8PUy0cY8TOCsQnlTGKiNtmPNc0vXnwEF4bc9cpk3ERoCjy4qtlF
JQoA0/uDof2N5R0MoDX+SNnzb+3rtljp3haYovXGO+cBf3EKpc2oxWChZwF1UtoDemtTeNkMhtpv
Hy5SylF90ZR1so2oge2mOzVT0EEFjXWiskxsXx26zDUay1rieL036gbvTvYM71zZuLjyetSBJBj4
bxSykR1xh/un5qYs5ayiCySH1T89SM1PcXaE228qhySg0d9S/Tbxr/tu1TnGeL5a51VWYf7YbqBz
t0XrlhF+KjB9LXUEQNSq6LefsydHCQdzxV7lwFSFeXVEfKR726pbqw/05lt35/T9LUBnwSPPJXUp
l6UdOED9i5y7cZoDhM7uCZQqiCQU96d04EmzYxnGn7bUDiiXazU0Y3V5rRK3pMJnrzKBb6Dlthf7
Fqp+heiLOS9DNgkgkDwHG1SShPJE11WvzpcWKFCuQH6FffJUEYauMsA5R7X+999v4XAlZv2y9A6t
3gmwb4WO57wBqyGk6JQQc4FfuIHCNPouFe5I5iZPb2NbsZbHFwl3Lpcpn1ilOTw7mbZgUtMEQngy
5s/2x+/sYDq+9eihG0+hr+vntaUC8a+l9KKZ6J5v6OPqC92xGtrFWbQspTfkvsBFofoJNSfE8jMB
Y/Jn1hEUy5nwXDgpt48ThH5lDmfSBjP4TUESIEoG1DocOxOp/qEBUL7HPk8UXGuB+UIe9HJTy8G5
nKLRBwbXyxRkCUI/wtAhlANgBLGeUg9twyZKRwcYHMyuILoE59GubA6QgVOTlbWQou2I6QquZ47b
cAeqF3qC7L4vaBIHdlWKqJfYfqVO4opRG5MQ10g4/HQZjOGCJ1woH9PTpv7MHlqJ6hS8ztMOnwA9
R6WorqweS9WsC+Sssy5j6MLbZXlqZzuNm3k1QpexeYfmmyCWITA4ko5iOoCuog/jox8GSBMWA8h1
DgZs214DxapG2HIZcg3CwL+Kwkni+e15h2vPVc2I/iNffY6LEAPkErkwhLgbBhz7YhnZIMZdRrAR
3KLox6O+opWmrxZbXSODgRQFq8sbtcaiNAZwxMHoGJPb6QWsVMvxtmUhO+pPYzcEfLE1Kk07ul/O
+2tNClEX2RkXyd/gK+PQNlTETnomYJPq9Swh4pXLERZa1Osu9O0VH6XII4vmgTyZvC4QhXXRPS3Q
crXkjR6rowVVRG/xZ6IA54EuaQjBYDP/a6GN1fCPbVYo4irOkiMxZGgEvK/HCxohPHRmsnxSSFtV
WjXhatldEF5oE/jRN9wez3chldwNa+AfXotM2fcIJ+IiF2tII6N0LzQIVDrU65G81ZbJ8+/FhdY+
u4YlPFxPUO8Be0aEGBXHDGqWRZAvYpaumQZPdu4bL5cjnoI3ek2sIt+eiQXhFRzLDH58kvx9l7y8
0TJuabfmZa29Y37FuE2UDm9I80XvaoNix+tth7Ks4eoRNU18JbY3V+X2X4LepdZ/83T6vHp+Ljxy
XrkmwR0Y78T2RYYDiTNLsuA9FmvPL3iuwLmO5R73sEPnyIIOw1pnppV0WIorTpytm6Z99uOI1Wmz
Ewqajd+GXkg9+SpQ1laavohhfbRRuRwx0NByw/973XXtVR5tC2dQNwm9D3YehKvicrE0CiXdHcOs
1mAHCNZhPtRjjJsY9HOneh+OGZxltWsbARHhOgPX4MpVgjBc8GLcScxRw2eRH1ntkOhuwbdO/XxH
4lm08G0TwCqZqKkGb9Jzd8vtOCclRVRxRLoW9jqrLK1FGowffjVNmiMe4bhGEheU0sT4NRUjshCx
h+J5N7ETQHEYKCcGhE91MGl4M5uLpQZWGYCj/ghpaicerXACiv0OzVuETqlOyvlNNNKD9t6i1npO
6l31NiiRX0nmv8FW4RwtAgFvsqGvG7VIKqeG5RTLuffL40fYqPlNP7xe33cs/P2peTrj1Pbj0OQv
vwr6KiA0DZCA/od+6BCJsnEmEFDF16+BVIa/FPxk+hXTSQkjFD+O8Nho+L5Xw8vRGS8jMsDuxfK8
S/l0uWosHbGouM8UHc5Dqh2zujuH8CKbs2WBiR+JRHUXaxGxlaWFctEL40MVdmYgDGsdPh8qe39s
6wy0O7JR38nP+j0hUScC0fV79+vkEwlPItDG77YC6vh8F/IiP7rchIfZcnBX65GxqY7f3aqUzam3
4cqlxjZ8Le3cuPu9cChY0GJJrcNpMbT+0HbydN9BPkqgckigHcxktLYxajJnf/TDb+AXpDy5MuPa
pxpLfaGV7z0V5CXgQruZq41dt7FAo9yRuv2Foxm9XK6sICiy6T9thSTvLXznuSygOGQdTQ4XujR3
LRabkVqZB3sxCLvQR/lz3nxGOSk0yKL5s21Y1fIdEr2gUfz2eorA73iAZyLhIZQwWgDJtAq7l7hV
5l98yMZ20KN369Rblhe7oadBqcj0FSpSkyIOokvmYkw2RKGjkHRhFtuK4VX0KzLjat51cpSltSP1
BXX1pms1/R07sbsa8skjKhbrXS2eWkkaaEcL/sbZ9F04tFiZHDQoIqyJwEu4QBbYxy5rMs048+kR
9/0xbPGobR96VKJeA7tT3GLQ8c23qUkeAAchHV3btAR+7RxvNZV0iZK+dEgquqDQkqLmVTtgoBVB
ebedfMEYs6+r9K6cWD1PLmev4lJwDSh+XM54qZBN5rT7PZ0VGSMyBd6SWB0CZHif1CUFyWNpmghe
rk/Pruk27yYpcSOsqEDViJm/KkRHPc4PPqUV+eaZ29ZLcmrSdbcIDATQnrMA4RJXFE6GYTjgOIVk
KXDI3ZPi5jaoLUkkZ15LK8ChChOPUfm4RlpqU6TyzQTDoH3VLRY1+sezW/C1GtmZfPvkw4OhooTu
EjV9vAngzIwJLuLZ+IyCOUYOxXS+n8y35nul50qLXequz3paPxE1jOb6CQ+ycCYBvu8xJQLKCbI0
pOLaiFGuvs7gd+eZF8doC38BdVvCJrm4vO5N15A8QjInERVczbLkKVnK6r0DwZBrduSklcrjQpoF
6Aflm/HpOPRMZvt92M7NkF90BGSbGZabR8uTXN26s72QRGwCVEuzaBM/dSWI5uY/ZMB9YH98E0yK
uJp996uyjRJj262f6lcPFCikWGk6pGVVRQeFlLx+NCFBJraOmYUIX9vJ+Yrvi08g407YwGdMj1Ys
5Ttilqiqxv9U+kwRNYTArRZKTrb9Lev5EtomyUe6/YZsKKcnXZnQtNnx1TQlKSA7TIQ3BEy3VOFO
2sIh4iWv6xX69chBn1PnjyTJF1bMSAcUUc7M6HJ6Yl9opzpW+rvKanaue0Avulf0dB6jjPgbo7Ql
0tuxd5UPBsdg5IwtIH0vxeV3y+riUN2+IVEmPY0S+t62T212BB+7LQTRcV8dCWHo+uch1zNNcwbd
iMHXQCqQzANrcrT/S2R3SOYG+7Vn8ac9jPvjB9uzduGhqb3K9864uc/UMkyvDRPTFVGzMvcdTT+h
6f1cTlXCNUKjagsJCtKOp3uR8VLwVbHw12Am4Fboa4qJwq1r4hEHs/HGnrClfmSbWCuuHnRlsOfc
lCECdS8uedpWgUgdCBVCuYWYFXs2xOIbk3aLShP0neJPxxtfCeOOOU0xhkvbMdNDVasuZsWamz1a
yH5venBa8EvexRvOrwu5bFORFrlkXgM685Qg9AXRUFlHXGzCWInTnHN3PleOlH5X5K71LTcQFRqR
11FLbkalCw25tMnlqNFchfdMTAqG5ilL/fS0aOqZTkRs0AIt3pPWBCbmCOJWqotd8xQnD9Lc+0Ol
R3iz6pgtu/pDZwXw3tt9FHuQEUo2AjhKUGjBXcsbi7BHlONyRarN3ycVfSnfrPE8aeUq1rt721Un
CLVWC36lmty4m+wrtkdG6kbylOSgYfl106r25w5QXyYYLm7S38bW1AFSpKzQafRvB0iD2PB4gtSD
pYWs0pPbCrcNFfQ4f85AEE0PwBaP8syLM1Y+A8Twi0ZrhELTqSxz5kuQpYnJgYey5ywpm0AprC03
S5zRsGI9Iid55UesrRQjGK21aAmFlRmCZvFzDAjfSA7gmf7XTZE5oNPs5ta4FE8wrVvmyj9KI4Bt
Dg6CUX/cqMRX/g6mrU6vnSpApjHOyYG2oTN5Dh4MhzqfVqyBlu/5ffqrGMvFwtpXy8jpbWIMm8jQ
DF4GZxVaHBRsVK2PBbJ9R5AW8CXowG8W3lfuxX0Wfu0YwizuUQhBczvbF45gKLgWS1eFIFVNWJOx
RthMJj8pjznUXFJsg9we0EE5BzBaPFOYo32zTeTSyeKGe6nm3InhpRizoZ0hC7Tzw0X4BT/PUNsQ
37QlybK8TU6Y74ugJrULgTRWv0IQWBuoZB16oaVz+izNFuYqdZBb3sd5+4UhPUYUejxLO/IUd52t
Bc0tnRvCW+isHZc9OgVNTzFhXvwIgtmUeCl3rUvwF3BKunzM/xpx7dWIkRQPDGDPAacHuXbdxefd
9SgI8dnrTMQAgyPvm7qfD/VEa6EebEXf8umC0UYv9F0zHmcvZ6I5pDdT7N6Y/DgxcOrQVyJaVNXA
TpSCx1IFjBdlXVxrp7zhl3sCzhGqYjftTm86aqFytj9PQSJrJYJQGp6schLcHkgz8wAYVFjL0YW2
6OH+XrThTbpqm3HESGnsR+4yMcmewl6/ZkPXKoXT/AvYdxOnLIrovMX0I7DuBimmRwuAXBkIijXL
lzC5+GENp6G4IM7B2hltWzk+e7X2I5A2wgB6SjqmaB4cCMwwkerw2bRoXapgbuI7H8bS4MCdLxR0
FWxylkSETiUDhcNSXCXwQaBCJVnq4shdnqEFoA3869qrWSUJAvSpR5naZ7IwtXjtP5EIHAMq3q+T
fblZIbSnpCyAcXdD+/IPArReUXrLwsjJpagTe5yRJxB3kZxRoeQiq5v9t4B9DybMZ+zRW75RC5lO
CPyw9S5YxrreDHI/DDOF1qPYC3H6Plkg5ASeoNLmlm15VFOVLP5T1WL2Nf217yS7+ufBhk6+VcWE
oxMfR/5H6V13s1VsAwWcAaAWCgubs++qZsmJtIZx9sXvpI5kXOGHini/9mgyVUPM8GseWqR4KglG
+ks+r/DgBt1iuWmON9LD6rxW7cfGXIuqKbwRW97IX5ROttk2+L6QarBehkBPDKQjoIQ1vD1XhkL5
Ka/MvS20iW23Ykp/Xoetu7tvOOteXHr9mn2QwXIzFP7QqCfc2P2gcHfcjGci9Y0HicamCbFla5IC
1GTm1eb+4ftKFuzd0pzwhZpilhQSlN3It66u+siNRIMUzxZEmToriPeyMxk0rDC/b+zcS1/GTYOw
3yZ4Ng+K/ug9Hig8UYf0POv1edGA/UkW7S3sccw84O64VRZDRpDh6ZAG78+3yT40eMCsYbXFRiNX
WtVJ9POqyd2bezB3J1w6kh1cPHyUBonvyNvz1wFKGty8GO3l5Y15YRa6fKoK+c2Om+3Rr3hx+xZr
/fkUqh4iqc8HefjAefl8k2ZLYilBjTSuX244NzMGkYUNzixQOg2N5EFVwC9vjYkomNJhIr6KiHR2
rOu3tiARc+c66WUSx2C+HuZ7lr2o6LF2W7E5Mp5jrXLxvKYTGcuPc13RgKudjaKJBePeDyQ5rgVO
VJoFl/VqVLkY3rkE2wvqTFzc7kJ2fnRJ+hDA7gmOWB4GFukJ+Ckk74ptFGEQzf/1VhmQllwtsumf
/3uqoQPHJThDKlGCqdQtbHQ0YEnenj+Pegne30c6geCzjOrqqvoSTC8w1r2hdDmPJCax4rkNtIuf
PXnBM3n0pG9qM/gZplAx6sU2nIG6UlCkrYnu8b1gaNJLfb4vIXENS30gYlCPNjcANRN2DlWjarVT
vJo5zny61Co9YMKVOZ3apRCmT7LWUqlNKZ7sLBytvMJ/nlnl5Hxz3d2UOJXX+18hJFyeK+wZxX0c
0dOnvTmarrVEd0Gke9yUbxp1FG/ooNKR3kXVPZszD8eeRkrlrvTDxohqrsrzc6uSL2tB5ix3I1xO
hd/2yQjmbse/xdrw7x6uTXLU7axtxtUVIGPoTRpLqc0s4ReYutZopGQ4h9F4TayMtqHpLboavtRp
KcOb1Fo8bf5H0Ow6TQpfivfoGRQ7S5UoYynElsL5plLyWaQSeyNDEszIdfDd7ZSCcKVqRs/xL51p
J1tuAoezbtM+MbDn+cakxuk5GfHls8sVSY3Lt4uR7iRb+o4u9x6f3j7HuBW19zp9x/5MVOb0cHh5
EoGv/SDSWYQ3SNBPgUSpRGf8/BvsoY9u85QgRtEvpDnnTjJf43oO4JUW5VxGNQAjzjsS+HoYDe+Y
pRUfKGp46wGkeirYWA2jpfcMGYB7As9mBXeP37JVGzI1QY7EUIeRmJEbvvcZM53LNeZWrjAmpDpg
4hEN+V0VhtLybFgTuozxuCsa/rB1FFEVQRrhrYalxRWRtwvWFo5H2D0tRwtA7S97TGXI5ZatEh3p
B869GKuc1p3vl1NCPv3aNvvGRahBboeUISTmTdQG5MNlG7hljyvbj/QG+RXxHWYOAHyGWPobIo+T
/SGNY30X/ws1pC7VnGyrth3KoJIxYR7NoKOSVWz9ZOibo1ZyJzrNFdQz0Y2Sn9n2vkKsAfIXCacs
BQS8gj+UT+f+WVH2IzmDzIYuoSjr6nMv72lUTdkgQhoxdkBVtOJ9+BUsdC3TwfFPzBAWt1faPvAT
F08BOBXpZqttolMSP3DzoUu2K8I9DX0W1oeACzn6Xzr7qrP5Fs+jvIy7nFe5CtB1YHw9TVXYQhwN
SvSTAeFSq3vjxZCNzKQTU5Ef789+ZvXtFego2I5cH8O2gUavq6wlPdayWnRAc+APsICbVq86n47m
7QpHcJ8encI/HW0Zrio98U64mvSEa6/W3Do+0lvj3x0nLAoidhoQHwFXVpKOKBAGd8V1bOK0WonP
KLQ5EVAw1oRNYQjXtF7BGwHykVUyh1/cTsey9LEKeo3DBWQsrhuZ1QJVJ1z/12ooD/g0Hk+anVx6
5T5VWowFcnp55xtXp3EoA2Qu9B40hvCyzNS2fgfMkrE2XeUS/0z3iU+hxfZJ1YH64jXZoPkege4A
lplHKlz7QyPBjErAyJJ3d42ls/fdtJRS2o4cnsPqJaih1BuPzbVO7iFOkruEhy3eaFVCE1XL019K
oDYAabvwp6WY67ClI30Z6p0yhiHm0OIyswK0+KFM0C1rPLRaNGgdB+llL995KicS6XYI2EN7ku1a
X+aNbldlUgpAnL67Y2Bvnj6bYClDoM038OiSd63szc2k4lglMN24TaG45UbL6tkiJubOYKFLYgJ3
Auf7qgsAPDJhW8O9PE3SDVCsviGZTe++vPkaRSPgrYC9dI1vR9Y+e5WWoMndL/eJmtQFN9GtWYoh
gCUuJYkoISB3tDLsmmSrqXnguNwSrm7NcutGhPZ6fDvx6feU0LBiMUbcFoEX2Eo7PxKXamFbppRl
NfkkHTIpPSmglwq7ec5lrhOLmJj2jaTdpo+OdiEHD1wQ7eKhEMx0XmPEFoiYyU3Cao6vwXNCA3P3
ejB7RCKZkrCpmYNrWHP5FDcfx9i8OOnpIub1rgfFYxohrFGU/L5QEU/c9gTu90ZkxnFJpoBvGUeP
mYOhXxqZF1mGCDxr+hp430Fda5/KILswqt4RR1yERjktYSxZTBPLMnYJWjuKUOvJ99Ls5Hz8NEFm
OOh8rAy/d75ZFfO/0YJqpD0IHtZUW2DT8TE8ODoHS1NIqbQdTfxyAjjPcptnZa0KCWt7PMB7/IYV
xxlktout41XXckDFCt2G2PpsEQxpFZE20w+YjeLTr9dQzzHpPRG6oVrzOuN5Uq8kzohWBAftcBXY
anhGRmFY26LvnuU2zkR0rHJYOeX53kKdIjDP2Kp6xxlzxSvNMFeGpv93W0OkRMtr65RyauDgAqEu
IyfvM+u5lFa0E3XNwykufuFhbkkHo3bWP7oQ01embfLaOF2gLEFtK2Ps/mFYABkPjfBsnoLg6Cj9
ntM+VdPPGbuHv4kbY30v4T2lfnzBecHvSNUJIIighVHPFy+yg6QTlRdXVJH3fZX/zdA0utdTrt1m
iqOZdTU2B8O2PZgiNe4vu4nyNaP2UpUeo1IdO5yzD8L98+qXMSw4n4B+G0iSq/pkeM53FZ95hsh4
1HEMu/UUb0bYH/QE6wAQ0tVBRVLTqtuE4/AqfkY5xhX7wgQZufF1nOtnvDDuPACrU8qr2Jtj/H69
Tc5kKY9x/3hADRCobv1fwDDHw8y1tTa2SjfZhx9TqoQKRit2SwGAaUO2Jf9GYh5C7f0dJtZCvKeJ
t81e0CgM6+DQ0zm86fs19iTDvJ0BTbDy0J7E1rBeDhgApRVn1Az8QMtlYkJN0zT6Qtyj/ci5T0Eq
enxZAQZInzqz5fn5GFEpP6R1gyRYWReKSZwAtQ+1EBYSAyLVyHPgouzza3hifOb3B0c3mja3e94F
w2BAahwOV9HumPAssrcVuZuaEoJIvvhh/Efg16m8RdM+SVrXs/dg8uDVebH/f+1Z9T/QilqN6L04
SvEOwUOL/rs1ZU+OTq19MCWg9LfjXLiFUhfejnV73grK8vh3Dyn+KtbDeaXZzPiRCTu7l/5ZZXOz
iECSQ+bV+9runEDdynLH80RQs4/ox4JjY/7Lo/Dnr97UIosBO2M0alvfRBr2yr8xjnF1A2lk3bJP
nG+OU5Bj9/ebgRbNxNBdh5Ssp2RfeY7Us4GcgAPzUytJLJcAEBJRDJB6WD4lwmOVG5Vf/MXXvg/V
x3vpiEi8cmkGFj/6PJ/IFrROY8CwhL3Lfd6b0zmXyOMjEsPg0w7Yb2EXkEl9CPJ37ouq4SMeCrDX
0rybwMeMujARJhaDCoEc6jb/zi+vVm2hO96X/s7iUF5jJCePTkj+uI6JUpxozeWkdZ0RZDTlkIVR
kii/sDOleHRkREWizeVTzc4IuxPXmBAoZ4it3K1MOg/X0uGzzMHJlfAuO1rjhX6rQDFPysR/ylQd
BXxKS+6sBnsJehbDAtgUg7TCkV6BgheE9c8/Ek8m/SHEPM4QQjermMP0/dieB3pV/1YC7jT7OXhq
d8/e79irbW8z/aCXbskD9QIAz5lN3u0Olq+BNQNusstghnoNsV27BIZTz0kpOdoscxId4XzZvGZJ
EWvXPKgF9UqURCQXLEFj+JKhbmhI61/ItHpjMJZhXoME6Gu0oJG9kdthza9EaYEV9+psXMrSrIn0
Mk6C497lHj0AnZEwkZk9b2vdmPGKPs4bpYJTiF0NykSf6gG3KWKxMLJCj8mAyUBCGDodpdrKw4qR
4HNshNuE3cV8qNzkD+DzUtlHOFrOR8Pu9xyUB+Fqk3974KXVmuNOcDKQyjOlSJvbAg1mQh33W7Nl
jM7nFdtHag1O6t1GsKz3FKb7lwSOA9PfNBQfqtLRx+vjdXr4y4jYKyy3N/vyHqs5fzi1z9f5K7vB
96yQFPEGPain3ETkTX3lvJ5QjLgS4rNOc/gwTHr3oMHJuT9lExPmg1755wUxhryE/4k4AmMW4iVx
hHuMExqlSpIT1sARdj2x+PKGhi+LUnEMrOzuvz4kWE/Eo5Q6bPX+roscIcDF/S1immVrtV5jKsm3
jWJtr5fXKfQ96EW98QkOapAnCeiIu3w3b6SWfXjww1nXGhJTxuNzdfanuRqz9nAz8bq5HMx1tY30
zbZw6FVI6825cmQ1wQ1RPoQQp9rKQOuhISNDLhbOe7yDSVdPwgWaK5o4NqhdV0CLPFUyQyhOkvu1
ERo8Pe3AjYyCV9lxHX6hKDPc+Cc4yiA6EJuEx5WebTJL0BfwrBOLcA0ClalFEWefBqMZJa+F6n2V
ZqtGvmAfjsGtvf5H1SfNW770xhC3gCbfsXFqqbqj82J4dCUnt9RqNt3nuCPgRzRKgNuw736xmEXe
DUL9Y4fNurYu2LsSSmbluHdkG49Z0k7Wap8wA7NhRoVKweRDDIObHLUIU8LGAR85rcjQLPLu4Fty
Yx4/URU5hf8/+iqCQqpGJdPCJa2XZobzCuQixYREHLKmfKvu4C5JnAGr7ZnXI1DwneQgQZGj70AJ
MiXdJ5DiG82nxwKxaigK+upEh9GEmySJdHKzmAE2GSgqXlmuJ7uOWt82TwW68il+Agp2YNo2yL4I
TRZhNBklruDSXwMt72lQvRKz6Lkw4+kb/ND3VdsgXYxV83sHu8mRJxbw59wKnTK5mJ5nbVvbAyHh
ReKacYE+/0B1OCU5GbteXe0QLD5zVJO/5uW0rbBkA4sKFkWKKuFc/3E0ha9S2Csp74HEuqGHO5gy
WWj55gYmNjF2YKEJl6YSNVTVfiZ5/4HdyC5RqzuzZr3VcavFXqTZPlyF/Oqig76UTNnsFoBeFVtS
QgRjCuFF+YHtjQdofbUUOag4OISQ8pZBiCMlgkY/Pjc2fhRAjtnkDZTSj2nNva6cETkVHmv0NT6+
PuV8rob944qC1DbXkMSRJtlolrESQBP/o/ZdT/RGJFOvzdIZ7KellsHhz8Qxn5AJ9quyBuU8FVUZ
ayZi3IfHoU/alxQan/vJ7UvNz3CV/tFeLYnClogI+FVp9XkXYJriINPYJjaPbTzJlQ5ngSdaBbIg
mQ/OnSIIqYAYkhlYlXOUaHWWmOskAq+IqK0eIanpJaETfj6sPrdt5FWvwn5NW3MkdESlrwu6iD5B
y9kTO5gk60fZskTniG1gRXfFl2y0JnmAKjTQ52WJm7QWoiaFXCgRM7mXdKo2aD1FzevcOU7L/8Gh
5mo9un2CwM1xpgyNRDJP+QJ0M+PtQoCiE7by7sQKylfkmFpNb7L4qG+C9/piARPdQtmHkHD/74t5
87dkHHg2zuXzVZgSW8wASo4nNsdIO1yIQaf21Eeh0T6qGd4MkvgmmslYjYt7OhOVMIhIlc6vKU+6
94mTSG4bJ2/xNshDMANV/w1UZK2Eo6Q+uZdfMePZP6XvF1lq/VMRBBUQHV1P4x5nRh62Z0zRzZlU
HWsCRaNXUK7jgTB2L6cRTbVVjQg67y2idHH5C2w87ENKEaWlXgWLckvNSgPOrxzONuiU4UIy+cyC
GHocaxF8PYxrCBkhc30D0TjLe9FIC/VGGOB1bW9Z8rQkdvWx/3YQobLJYp2TQJlTLNWkAb16yZJb
e8z+Elc/7NkOOuH6hu2ktjT5ZBdSXiRFVhMD7lR8watZml7X7RLDXbQaWlMcqVVs5N6mU7ckeSTU
dDNqbQSsJLIyCCDcRgR50TSLz307tOHtoWlE7oXGSxuGyAZqnbvA0lhxw35+Ibb/p+vkn2Fobu6m
5KNxt+cfc2/r22q0OqxmAwq62pHmHKlCHYnlcjnw7dasRiJA315gibkTY+g9VJJT1D7ZpgtY1l8z
afm2iol2BiJGEomaKqurcQ7zStZTyC41EwANgj8n2HQF9TZ8w3jUrXTsfLPv9oHSm91yzMkVjlEH
+rAThV0FuPXiEI2ou2v5vSigjbxrgxChcgS8JUF5jFuC9zpavd/X6yIOHbBvyBXOCwOoHg5wmB2r
k17hhynQ9wxFzZ7ozp2xcRgTN/yWJprjkLQajPsbb87TNm38Hwi2zJOxW1rqFaWYiup9wP3gZhdM
T0aSto/ybh10IrPvMutfu2YGosYcs+jYGylVgsuMD7ZJ1gK3uAMrpj3YEkXeQCgp39nhjQRyhLJd
WcdZgigWlIpLEpAb2LKa1HmQeu6zeZVTmw0M0+dVpqW4a/tuJ/HZiad82zG5A5hAFdfBCAHr//0Q
XOXh9kWeRDZIr5Vi/cWXd+TKxFv7X/7wCkU+Ywh031KjoQ+WFMZCjnU/rgYipDkIK+mr0qCp3hEZ
EGxmJWAyCsT7gsrsmR92n4wKLXLKtnAzRk1OLnUAVakVj2PF4bUSQnJhTnfPDxrXeUzWhE3oSZvJ
ZleDmS58LSB5+UQ9RGOjSTrBAuWd+GgZ5LnNp28QCTZ5Xuun9PwdRqd8GjG2GUEoHGxWIi3K4+Ei
0lBaQf4dBXT9wwjNzJErpz7FCI9lmlF+g2iRL9L0GjO0Baf+JPXyN+/Vodjco+Q7bA/1MSgpLCGo
L0fhHhwyecHECZd8EZDG6KsLzd5E24zzc7cdBSYw4rWFhlqcO2SN/V/hMm0BTzAAnsSeslcUAuqW
fFAtpSac+IXFWv5yZ+5lKIGCDlLsgFyBPgcKxez5qzmSFcPxmKVoVgw3NCWQrmxl6ZOf14CGGbc3
PhjURCnQ4142491HSB5vhR4OMtE9bE7RMt9uD6cgNG25r1fwYhcZyoozt/0wYNeX4SbH385AyclN
aIsTT9zsMJWkbWsPm5mc0YJUA7SLUKhPN8bSeGWahAIPltLPWybedhRnPscbtD278iFk0Z9Xv/+A
X3NhIyXjBEkmbfwHGk2AZomWKXeLKA7/WOEplDUKZe1a/ZVof0V6DlOJJtCe64HWP06WxZrbgPO2
rTfWHsOiFypSWrmOfSqr/JyRhF8TQex3WlGC4eLwYxeR1fg7VS1C5M+AdMk71bn+r+SskQ+k9DHO
2Okd2D9l1sp8aCLcaYWI+sckjDR0Y9763Lek9vhaw3Y4ezemS/eNYZ5B7l/88eHsEEPjYoOy6DWT
G09B+Pb/jTkItO1C0JM1G+VpMMD4yY9iKBphoseA8zcAtuVBnJvJ8USPGYbybg0U+hGes35ATHrU
ABfJi36MomcFvp66Ilw6H84FyHusi6GKdfK+ANd5MQvm0vWWoGxoR+zNvgmowQ7tvhM22RDscaIg
bGdRmiLSbk661xDgK12SmFmacIonf45lnBZwoMh3jyE4a5Wy3kfE7OrR/1lh0ePFC1SoblohQaoQ
hQEybdaYTjXY4L+8Vy8XCo5deVVliU0C3TdIrpQC9EcKpQ/NPTyezgePW/5H4/1v8Mg/B7Q/MPX8
7A03aeLaMMMCmEScdd8tNEA/WFcAJ2eIZCRz8D5ouHEEzckcJNbNl7aRPPyr3cCu+CGy3HQMj1UB
qYVDoLbY6jRX0w3E/Ip4BBlKdKyPRfQ5LXo3Dzc6Uq7dGeWWr9mpy5OUKU/vkTweJ0a87LBfUyUG
owP0LAjhdsJnV/S0yWiAo2g4HAPXVDB+DbtGWB1IJCbkVDWZGwIC/n2TD7OzIj0K/J+NcwlbfZzn
LLEUNhnsRLmNMRfgpxRGnRdoeg5mBmzX1r4NniM0C2HYGhH6AxAf0OZF34ANkhYqTEwGqnWgoyq8
Qh5SJvKtViy4BMDYkh3w/SPEyuuwlRI+E3Q9RfmDaur/abeO3q8oSxBPYznOlQ88jWpWVwlB/0a6
jhT9ssy1d2lpWz5Za0zoT+8sE//QTj32/YDKATrwSL3ADjyWzD71UmBxQ0IMEmB1+o5QBMu3focZ
QIcUOVll9mKdjUQx6Vkc+3F9VbhJRbCen4uO7G8YitBAlBcVk99O8GllbKVaXdFVzrUOQUTUKOFJ
DzO0Jscwg2wBHFGmTIA1wSkusrZnWuMyT6NTNbjkx9HFfn9WhslTj6ZpBDBtXWPgpXp1RflMviZE
A96ItjRyTEZr1cDckVB/qhFjAiC8e1SS7uGFhYJkiFvyoTCz+QgGCyRKdlOOLimqnPcCAp7PnGyi
7Q7yNBZ2uy7NwG9uXvN7hhkolr/g+24I9HIENv6QgQxi5Mv44oUs5kxps0MPdVI9Eghb79ejPHt9
1txGrnOTINTtvCyxyyoKDPGSL7iObB8QmWHDkOn1oLFnJjubMkkU4FXAVtt2gbH6uUe2j2vMM/d7
ken5rEzcKKzdvX7NrZOTecvF+u+jJao8bhw/LiM3SsRgzngl4zlsIWqyUUDNiiA4P9alW7R+cs9t
S7uykSlDiC7LNrkH4eiwhxrfnfNVO9SDj+E8TRh34btGVHgUYo2pUoS8+uQnoYUBNLxjW6uqY83Q
0gZF3u5GeVScdxRtncF0bhXdmXb9e3pL+FM5CRUDXwBalMV39tjqAoZLDKF8+b8BOA+BKPddpIfC
HQsYmvyLLAdyQF9jBmJqLKocJVSw4tf/DZZDUmsjiVZudhZQ8726NdfcP9dIN1ggeDpGFXgTzvEk
PjPTw5HI/lOg6N+y1zqhofBOXvX+xHD7iA2ymEFEFxuxOisQuDSFltR2PEDlpESGAEYXY5lBy7EJ
qi+ooOtsmtJooYVflwk7WfZPJ+zOoYCnW0pB6e+5B5z6N4dBiuYlGh0FzOQUaDvLppMoyYLF+s6Y
ni6MnaPmRYL/7CyiTYW3Wiw9K5u7wy28r1o2IjLss4lHvKR3/KxO0iGs8FRMnFq3oiE5nBljOGDp
+MYcFd9dbRDjfE3XmqiiJ01+8yuOSRqT5wc6b3JWUVa9yTD6eegcNd6RXY/K1Y6I26ciy09uangW
CTUfDTLGXHkFo1O+7fHxZ1Nm5ys6+COtXbM9vpscpwqJA0k8nZgy+FCcG4C6bYIO+hqyjfL+AmE3
KkH0H8kmIwGos+rS6Wy1dVsDsdt7f6rPyNhihYjnqdy5yciJbrvI080TYYnQ4duCYxRN9LepCO08
hFq5DeFV/0ZKv+RhNjBAcc3V8FGzOZJmmk6yqEV6A1LRXyMQt4vJCFtRzoNxESBQOpsZYWJ6ZdlA
VhywXXIilEvC3jenPLcUHWgh8bQ/BdO3Y3bz4ObFLAxqUs9d5xJk8MW+j8Fiqk0CTu8hYJoymhO+
Oyw3A5eSMMZh65Q5SPTz1JC39eIWG3whujptKcb7+RzqPdtcGS0tTvq+Dw3hc6nECTZ4DRvU+1aD
MFT/Zupoi4RETiFM4gQpsbqERWsWD+CYJu5iYyAq6LTejUYVfAW82+ImQE0bb50wc2yi4Cg8WeDq
yodsHgIF/fzM7+MF/OPNoTo5XcOTB7qEJnwzzp6srvScRqKrMAPs3TGrJJTygzV28MC0UNlNb3eG
egGJ1CPCmOYycxsM1j6vCaQy1x4psLG3ab7adoeBkWEbAE3V+ehHUd3/n5lYQ22ZbX5o2YSgWW+d
BWoi0WqAo7opXrkdOT6LF2IK8wpaqu1S644V6HDapPvJPKB9j6OxME0P6+tINCUOLIzLCKihJrHN
JaCGlB842dKEOOPTceZbUfv3KMeYkYXRphH2U+lU2RjjNzRsBaVDftZD8E2sqs3Z8gWOQq0GZEqe
c3rj1xR1z4MiUza4YU1kChDqFNK4mTsLMp4+0eVTBnVF7Ea0mo/Z70zog7apDMSXqAc4d/8U3VRi
EsYWhF6vMHhhRNLP9MAKg22xn5USxRtgZCkxoJx5iwEV3hVvVSF/Al+nItFaCeXeFNz0pmjRxV03
lKF9z/QSd/3qc/iMH4cMRn29hPpgkj3RX0N4+Nk/UsZ4/+QuS6Qi08uIoMq73X4/gRe9GMGm3aWr
sjYrBC8NtmOpjUovjdViJvY+YIn9Qw51wkcGGM9yhfCE4H2jnfnH4KpK4LH9/x2VvrGl6eB5fayN
fvNmm1USFNQW8qXMFZEjggon4Z5gqpd0aFDiu4KGdfAT2xjKl8iit24PZIAm29J/tW1SgPlcRTQg
hEqIkIHgYgSK9NbIECoT3kmW5WLp+snRlVtutrBi4X9cjft6tQ3sAQi7zc7jDdF1fFQcmOy6nTb1
EJIdW39FvGdUaEUMMWbclbC+L0+PNhTCrwY2/82v7bpHjA8PZmwFkPlik2Fe6NZ0zO4zQ1saD4Lq
z3KnrgzBowRKvWGZAkSLIpjRQM2L44B9LKIhqGc/oND7Bb6wTk1RfpC6yTjjyzOBAO+icN7CuMGx
istjid2Ggl6PVTdVVut5OsC/bvIWx11qg55zXvmWeCs04ss43lHtIcF78h4z/qSYVRPRZngs23Ms
4fxNBL33ZNd2H9laE5P1BtLd5Mh6Zso49g8fwSkxzXaTqbOfrH0SizCAu+IU4GkZhFJmTA1YT1wF
vtLZj2Q0yaqpeJ/42FC1u+UytvW8suDNwxb52+5l8He99x+ushNTvzQS1yK2Jmf4bum4Gbq7zG9w
4x66blVlNBJa4uyVnMVNqVUsPvE7e0szstuqWvvl7edBQd9AOwcnfqYV5AnIux92bef0eMYxTXDW
Dl1CptO6uYd+PyLXUIIPrOcR/9eaKiKTYASbUkd5i0fgcpXlp4fQ6DvVuJ1YWLqeUJgvavRnSoSj
lMRObBLNFgtc5pIT23yf7/ukzWOrijTc33sbYzvcX0bHdOqjb3dSCVELwa2ilc0QGnqijtuQ5q9R
GvWn4FUqXx3mo2uCA2RmmSa+DhnlDHf9pndnuUqHVj768VAM5IcpUrzwDNS91p1y1rsWt07Y4yX3
03RGKvPzBxqH+ghWm0vgLUX5hVLbiA8126FPYLi+rnf5qSkGcNZ0FrqYGjiOvsucfETw+fVR1vl2
VtXr6pzJDOPAnd38+aVJY8Q7ILXPqYuiaX/yVJhEI1DqVb5pMdIArZTBAFOplynAvXSBK81pFNwE
8zxyopOhzo6ZuQr8b6Gjh+cTu5hgkg/1aapKDOK+13sZt8z3OkDV4DJpNqY8EOXgFp31ocFgLa8r
Jn7Jk8VXEFs36+3DSiGEsEqtihxaNAYy1nM+ap/XMpBGtl1GKDLo31d9hWbcCdncR9Yt7DCVzj3Q
mlCtAkCg34CbQLTzldBNOnYH97+OjCtUr4TlW/DUaVpyxtiFNIyYJ7SNsC/SaUk0jGbQI3kArqeD
uoyiOfRomjJPuyx7S6UvXIdKrJAwcEO5ALAZkotvI9661oSE7c+KXVO4LV34FuEsomf1AFDM7+y4
QeswHL8lCVceJbbGWBIT1moDDyTX8cBLsNtG6DgZSz15u/cembh9yXiZDAYsZXTaPiNkLU/U+myZ
pq1uVBncGRBAYQSdqg8oKn/ZhLYrEa7TdN4zCSiu9NSBgvVSYmd3U5xGM/Oprrw4R3EkbjydIEBb
+NvO/88OQKtIWH3KpSWU0A4aLaGVQvedYtotiT7v/NDkO1vHgzaGSCsAafM6ybPREOuTjNVUBMLn
+pikip6nqXA6YZMk4jQnT4PZRO13MRjbAPuuGg/tSwa4Ok6kpeUNMjC4h12mq4xKxqfiJcDeiYst
c7I19ibJRcx7XoVRxDeUPgTGbGR04Yr7+O8PFfKv1y/EygDkw8VoZbLlzC81zrq9FWpqxfOIZj5s
cndaMsd1q+HHr9tc5jzmK2x1kF+kUOHnUNp9MmIQrx+9BZytRU6Lb19bWemfr7A3gTXrWDe0fB+p
src/sKctmIzJyaysMe/RuXXUKxL3iiITIpIELoSgwHsDdoGWwNvzPsynX6+3/+aFQOELMK93UCCB
ZxF4Mq7pQv7IfP2aeK+C04jf47iGW19VjMAMwaUXOEMO38y1RlslRrY0/XR4Lqt+TkslCt1EE75S
RTPOe4PNVec6I3NxPpZuvL4Q30srUcNla4igJZlp/QBGG4fQZEPpRwDZAP3Fp6EW38I4Y1BFc0Lq
Hb0Ep4ecWHwcQA5AgIYcIftSKHE/ZBS7/v5iAAPbvX9rcRy5Z8tr2yhX/wfXUCI4g2mPeEFD7/KY
/iHXOLl08E65qaQA4kS5OvKvE5qdcw9KeY264radOzF3m1L1OrAVp3kmbEAQNa81OrlWngR0yCXT
uEWd6guid0QJ9c7xhN2c+OEtFbqBWi0Fq3+KuosULakan/jSGltw709gHGOITUZEBz0iA0CgFISm
Af9vo00KpOS8f26xSd03/IKmFgV3Ac9XwIZ4bYUP9ttVljiyPio1ZSC/npEFjx3FJHdMHAYCqUAi
ppnCg/nuIfKYf5K5RavKx8QDyNkm5qcumzSMNa3gl7nollgLGm/Lz4riFwTUf8m4wwpSz/V8ydxL
sCfZOXNBJtkPxLmecXbDCurFem012HUbfcDKIN9alzZt6yVnxzp0fLi9MBqFvjonKDfjNaauv8jH
/WJ31Q8hPmuBqq/2r5jymJggk/AS/z/uCrxMGHxf5SiQl2sAIWqny257/t3DoT9PgSM3cwxJ5NxQ
4GGxF+DljF+2jNxBJU1Sfyvlw4h6G6uLpofdmXTZn7TKJ7PB94kN2cfZaoe2lg4mReLzcblnw1+Z
v00Tnoy54MoQIT1mHAnlPiJh5iAPeJCzdl31wcp2BgtuST0j8RdWZVJ0wwIk51uM9CeOEiQ4MNID
HwSjFB3Iblr4sVSCimRP+wmSHm4RDWTnRZvsnmeIa9nw2Y22aOJ7cMtLNfbx6lB3JWALqK3TRgoy
E7x7BJrUiiCzuHv/Q01Zunw+bW1JBrdcygh6t9ph5+KWVM3zs8GzaMNJRUCA17hmXfFEJHIx4uCT
PKY6wWErcLDdeKJTrx1HJFYuLmcBWw0xTYQMnaLTbTBDXlU7QexlUV80BUDZJKBCs3PJwhHiQ/Uy
vIQ+UCjU0MlCyTe8eKuraH6aOTrJCkbSNGrsAhHMUZv583dmAxM3i+MiZ3KbujF0aJpTx0NZt+m6
N2v+xVu/+zQhRjcDyRjqGtvAz8M0qaqVfQltz32AhUXRE4UVdfQHUFUxlkjdxzwb8Q8op3pVAsgm
0/VTZdzdbCKFs6PS5cdACwqao7h2fnAtGKcbqCSp8DeBJ/QWD9mPAwplAaB75lb9/nfctx27nYhH
kTVkGPdv0NcUjAgsElr87nEXwVWMDZZL7dYHNhMUOpdYvyNgqFo6V4R/IG/Yjmh+5Vg3eOhQIz3h
5sOXlwIk0xVdwnkAP2Y8t7kXBKoIueSZZZqSop3PLWpi2hMID/N3UAoKz1YNdI7kLEFaJoHgMTj4
MTCOAY5gmLzydVzZlY03lkNbwytJjAQ13iTC64JHD5uASvv1xa7bYJTeNfKGDnPf6vpLFb7jurPI
uJ5cqsdUxxW4mAdQBRkAGLxMRrMTXLLc2Ry474vechg6sr+ldxFrTPw7sfW+fKHsW4jw1gqRmgVT
YrdxWEVa+u0B+xbRq1nR0hWNlyyun0s4lcof21yrpr67CdHH1eY37sq6boA4boXPuHckqjV4rgrL
1ZjDYq2H87XDEVz/TN7j6xiDxWCf/c+WBDJ0hDOFA6XfGgHTSEN43r3SrBEATiXOYTdybeMB88Wl
poQofx1unI40AEmF/MIxUDU5xkq5puWdxcb5NRfAA38jdHV/rsKDslmy9me1jpN4wx3VjsAECwcX
2GDq2AsfhiEdtbX5iN5fUwV97xCb+bED6pukG2T00MSkDjwX1zyqt+VRgjFlxpoi40+sZKNs4Qfh
Cc4MZjLf4DSqVXJ+I1c54IjrRABxCyO4wMvzDXALvmvKy09fBYuTfg981onFO35Y4SiYOMG6FLOV
i4guishMCg2sO8TbdNmBFe2aLiIxojCLOtcZk3DY96/E8CjIfkbvCH74e7esNT6RS1OltCECdk6A
lHBMWmoqcfWVzpY0JmDqbTanY2iVXgIkFXJZ8SdGeh3RQlWJB7vtRJHDZ3FHeLu7U7DSR71Gd8Xh
mTKzeWuZdn/ce0aMzo1bZXWYrP5ORbqpEPD+UcZdOlRHJA5nympCtuQbxLAFf6Ox7h+2F/PboBQ4
S0djM9oGqPD9EdAj+XmOkqmohNb6dfCrOKzQFC59RJE98NIjJU5DxbOhEC6qEywDViURt2QX4SQw
yjTFXvBVYWGW8EVjEiwZK7Z7LRZVCg+9odpejMxiLXENDEDH7SX4pAmhYSvsHnwh0UtrmglUvhJQ
JNf0H8mdtkJF1k4U3xE3ISc0YzKiXvkLbNwXADaqIooY+amvDI4SfVbtSxkLSgO8xc7oBu/s+TYT
dvVHGyUR11hRQRmkiC3xyBuIxin21uzyj3P2jROL0dbzo4LXuT3orNsiO5zUQtmYBZhJiUHLovGO
a7F/SwSyJ1qontoypMQaZJQb6+IBEWdPdGiNGxcOROCpCcUeiwjKLOF8tcQePiJs2NGwS25krnNf
aTLCLPEzg//DQwIASVe1GtcXMg0STfO4vMpEPPactstk+lJ9SZMm6uXN+e0sLPTAzsFfHKBV3O20
LYRiEgyv8fRdp54GrQqFLBV213NQAp+Ot0uWiAlLZ+9HSIseFCzpRGt6MCmBXQSJhwitj3QnvxBE
+ZiY3ryOnLi+JplIBedH79hXuS+E8uBVsE7/1ZRuf4dHSRhRw0X66uyhpBlyrwLG10UsTjpw6+m9
BIgFLHXMABDmfZjBg94oAfFdS+yz42XzfkQlhtnYnTGnEgixMCvYMtlzywHB/ROA7AGDWeiB46vO
v4cvXHT4G7JsZLjZiG5cbOW6cGfUCAZNBGnuSyHiFVdSKyMe6VzaFndpfiAaHIMucDkr+2NjulbY
zJgOW6aYiTS8AJ/dEMgOTSdQKgirxct5rWFIaJ51J12XG2iJlwpGFR64ZMPLWydxTeawHxnwTbDZ
hbszgosJanXVDImCqsaf6FlbvNrIySlYS25WhYAWxEYQ1nJPK/RshBlVH1Ed566wdhI1SrXBnYLM
cyZy/F4zSekfW1BhO66RIpVRO1qc6Nf4sScRrX2ggdi50gnOp6R6MxfYGQYM4ISsGHLQ6D0Ub7MH
WcnXHEqjkyLm/iJEUa/1XzSjvinLtY+fYOWQDDKYLLi3n+nzoyGUEMn7ma228UvRHsMiIC3Z4j1j
D0aSf9xqz4U/Urugs4Hc2psaJYdEqetzkVqaWlYVcQ4DempXohPmEvhNIp528vVHMEukalen0zJZ
KaJBjGg3IPOutU0Uh+A4vh7uLlvGBfrhNUIfkopKSc8bOl/GJvMsonVb6aNJbcPMiVmbmYfvStDe
aKzwOiJ3Nwgn0w/wjGPXmMBa0gMvtlTRAWyQ/Hpw52Jzqanh8ehkg65e8EX/7Ew/XNgoagg10NWt
0w4dp7HYqR6v+t9fnhCZdzHJVaQkTWkAkP1boCzdSTU9GfqHtOTWZUkyBflxFaEYUPBDMgnT9Zd7
yIPOJm4JqBGzwKZxNMOGLD8tZPCgbr6/oq4kL5pzPOANBfquuJZqcsELVGV97PH2nTPWVJ8drsTr
gyugDMqbkkPcQ0f28L5DjV//P+CJfwNStjiOVAIVQEXE7EZI1Dzwz4W59NtXfE8QeMZti5E5TbFD
HML3LwB8y8WwgJCWQG3YSJ2Q4RKxWh1hL4WLEI0hdfUrfBya25y7/V4V6KgoMgd8BTRoeAvDbir2
L0n29RZDFdiKhd/c0He0q51Sw45rdjvSy0g/ojRuqkA43bC4f5zuX4oRvljiu8g9rKTlaVnfUrYj
fXkTmSIOr/X/PlQplQmhH+7US74B3bGVy2fCqqTAHX1pp6eUhd71CxBPJyMjcXHHbD9+IVUfBxyt
9RBTovcPmx7m7LinCexEJ8aTVu9/RR+LwasvJlVGQ9YN6z0Y16ZBqKtXmUj8/1dSC3uRqVYhOHB/
YfSjJznT2XxMMBXwhN6/DiuMZaTQG7/ejxu5iGRiCkuXn1SPbWo+HtkH1pDDek/Zcpg5R0xPTV9s
qasmEM6fsERvIXMqjcKlsyl7TmAovns1nBMPuuxU88dh8aHkgIZQhXNleW+T7NbGt/XbShGKQZyS
V7clfxKCcyTuJt7kS798EJWQQ4krCXHR1+zzVA7EaoNag5Otj3J0ZuSwW2gs7CHF6Z2odNbQk9WN
7MihZGb6d6wGifgXvW4vRWUalcl5CyqTbUkrBkb+udvnmeZNM6t8FNa8wqYqLWhqzYyGjQB5bW6z
2iBTggegLVO0oknwEGUPfx4V6BEBgM2LEclRMGLvnTwSvHYrhVarM22gwi10bIb0EGk3pNo412+y
OB1dWkgNZYgZ0an1R8BBOhV0nJVUS/TZwPQb6qXFtGuoyubYlhaAuCBFAh3hF/8oU16FZ3l7r/b/
OoiOeLyZTafllpbyZD+hdKQt4ACAiv9ehSZSPm3kpid0FSYFz6SOK1tmOsGOvQlseBEO2ehZCNMj
mhIb/s3eXmVId69ZvLao+2qOKboxCiC+rHuh6owr0sol2JmxpHBq3lh9+Z8wHidfVKXGeFrE0Rog
IaC8CU/0cpzHeEGl0JjyclB9P+B5yvmj3N92TWY+QojKzDKn4AGFVzsBNr6e874JT3RN5RfTOHav
eEv1BWPe7rlG4Lmod+1mxQfOqPSaOXUALTJtouZkPbhVf0HjNf7FrClDCm0K7qrqFEBtqjt7Cb9g
LLX8kZR3/XbD+kXpQSDTMKooK262ixc8Sj2e4ybqGxHV8eWLB2FckbJ8847itzLWu/kBoi8Pmj+P
WRIfI89PYNRhtmVtP1ON+wNLguw0rbvOQ/ejx624CVXVTlwahJMHhh8o83b22kKJ+A24R7+77mcL
UKLFJgKZMCxTcTVgyl4NwMIW0B8Q/X9qDIZkIxA/CaoFSjeQSoZPS+j9ExhnzXf8I61QwzznKlUc
BTRBHhlVqePFK4Jlp/7MaOWwAbCyilLZIOsM2Xvae6xWP18jhXnr2BtCSYkRFkeTnQUZfPxYLe7X
ogJYEH7CaYu/H7hOpIsNSFkWr6eZwSuaHBq0IfEU8sLCAsZNJWhoWINDQN7TjqsQrbRjh26n76vN
KUgNPIqMIDQBMqtGjRcmh7YCFuAeDlsAnKU4SwpRhZruRY1EsKbkK9wsNycrbS8Zqjv9mfynxIcN
JFqPskGvRwAcC8z0w0RnjEMnHj1CxdfukEqS4Ym6MqDEpzGTlw2c0Wp9eeNxpWMMFQKGuftM4ku+
NP3O2z5YHgtZNN3Rr/PuIwsWnYyoqntsxWMtzIcyqMCntd3myxOIwYI91tVfuisSno5Vf2ex4QsO
IKQKh5DQKLHf+amAx9jKYZfOpJye2PsQKW8QAbxM6WQEVn7tCZCQysL5OZRrLyDjAykFE/MvDUE3
mc1mLye1TG8IGm2tEiVtCJUYGpCXSU9AHQt1ytcxibE8Lq+nKKUhZe/GfYjVFoC0fiHJYpzNDyox
+pCbUD+TlOnc99MyPQiFidNZKLZeFHvBAwQ5TElh+sHElctnJvAMG9oZBioTKa4u5Ex9fvbfU0+/
XGVnKakK2oeFO6ZmU6TpM5/oPXCItsDL6cyAir9vPD8jnT+8/2NS9Rq6RuOrA3jBerP52+Oe71Po
/oXUIlRCnYeAn/6jXSDZAVu7xv8NXSiYZ+9v7oxOI2+CW4F4tkqUOlG+Ao/s3b768VB3GUnLNhaS
vI83iizYWi3hgnzw+kNoB3g6RzbsQDVPhtmowPAStU0yaZvNiiSD12G6tlBlM5hVS4r6MlNu5/Ok
1w+i5fRI/HU+rRcZe/yFlurTFe9Sw+XMQ2eb34SjIYUMGMpuPi+xPzdMBKMwyf7RNm1Umh9ucMp1
x3Lq8YoLULrmMSr4FJENCpe/LZI63ij+1JpkPFvoNSNOLjLGYuYl7Dg9cXZDh2sVAPSkcfh5yDZZ
TjoaBUwkV/SkwO0To36ucItVEt3Rri8R1zSgUGYUx2xka1T4ZT0JNgKlNrZ9y/5GrD8OovdRyH09
IL4CcHSests4Ee4toeGc9ko7cgswRfcSal2rEaTlIrikXet3FyXT9yRoPSlFeOg40T/ZTgbSp49S
TuEh8HYskY9Sf5HvvPV3pOmgylmHGRaiz2JVmFuszMfnrCGq6DOlm2Jpb6+3MUG//nA5vVJtzZSD
aAE3nu0h9xfL6fJEMK8spKn8ufy2tGTPrGMdiGMiu8W8cNjjTk6VlM7ALC4nzmKiKrtgNcRYtmzd
ekm9ND2yyw1CX0LxAHT1yO2Cjh3gJVzowf9M8Q75Hb7hmtacEvQSUlGRMn6k43RFZ7SAXUSe6Iv0
MNXc7CTLfbvnDgUvqLG6/Hl95O3NR25Xl+c2ue+UzuX/QATDYa/e44XBs5DPAMZOFbg5gp90lGB/
uYN0G+kKU4nVpYfjLtPFUJOPcyXIMhFXBSNFKKst8XAhMASNvIdHt2+7WDRcUenKnDmC//KQKLZJ
j4t+7pmd6katzZGAj8I6qzSE9P0F0q7LEO6WHMsL7IzHtNtDIZZJ/4EHSJUKphNpaX3aeGX9ksJs
40IXWQUspu++bWnrp+JZOeKmCzs7oGbBx4ODg5nWJfRyo9QQMQmMeTD0XeHweqIZyJtOcTYiVR8p
ruTiv4Mh1G87WVY70HePYT94sxEpd8kWRR1SoFsrC/OXZ5L6SNgu0qUx2MjRlcgZqV84lGBmTUa1
dntfDp+5mvABiFqBgarcldaLmC2DujWs7ipnbj8I5U/NJx3feY5xecZDhPQ8Lu9neOfDrWwcGDTr
4tHT6LkWvuH70wPldK9DMFBX4DGSeZvy4pmFWeCzyCNqwPxqjL9jSYKdIlgq/uTWVzptxK+ELkJy
UDGLw/bHsg8rt6Z2z+hl/Ko0u7BKafXQVOTf4jRR9Gagav/o+D18LIuAGnalTvJzDmI+WdPV/IWJ
+AYf+t57plO9WYalkZEDqhvbhRUbSmyNpH4kiYX2yK4FDEfC4LEPTNFWVjDPTO+OUBC0+dM55Sil
yB5xHLVxrHkgz4wiw7K80zfgrtJLQuc728U4xUUH4UN1MjZV/lOvOHmXZs156S1Jt/iY3f9kRLZr
Qpokr55VNZ0SDFNI5+t5EK5dbs0t4+WyzSVJubm67d3KNoHAu1HbqdVhRmLP5GAzibziFSW+gRpd
nXGNYgI4IelhXrIgogTrWgg9oxQjXLE1yfOilVkMx+YGvXR3Mm2ddRKpCeoAZNvfRb/m8Y9V8qg3
hs08p5QvRUeHpznPkRlmyeQ0vqUeUhV6zBhURvK6trGQDQO3kuWGLBg2B0+u6LpplPZ8Ga3tZlfn
OcCersYrxLR1qM6muC/KYN1NwaM60Wqwbbzop9pGNruQIwGSPgVrMO5Qv+tea9cDw10vp82wp7k0
3z34FODUyJgZPM5dWcxBwvJ+f0JzU0gX3hoq9TuRaO7FJGIl0snK9L4UGkYvQAeNMVUERol6iCyH
atUBEdTsTjU9XHs3ugqiFN6oKk5oCUv5kMPc1KVkwU8s5BQFnKXbujTuP7UDc3LbO4b7/ikNBEMO
3tNTNxfyttdY3vM/mVB+w2KTfA8S2yuMbSvA00YylwMuOgiw3LSG4MQnD8rjWeU6GYsckfwkW5cG
1WHla3arpI6cL55wPtWuG3wcSSLV6FmtUmJL5g36H+/0dQr+9EwlfB0kXFSbn8pcXS6EzQ5ztP5+
Kke9EtnEX012Y+1T4dRgwC5oN8JXpI7c9zImyIqQfqb30pHRoOjBuXvlO0NlbVGaDsijIRX0cLQo
gOcR9iOuMWZJaTNO6RhBRqLo69Az9G3RwP6e8SrUSvaPziCULVOp7SJSAbgybgHFFZxKc3RTGRRB
KdA7f6ljdpRL4okBtwfs4ADpfuqSMGVp8QFP/yzFe6UuufTP8WievPTMrEAdbl3HLLUi/Qn7tMFa
3dYVK8Xpa1U5u3KUmbpCy5qaEV64pSzG8YrkjasgWclSqz1BniwP4zWYr5Qu3ha6+vtmIpkHheCH
kPOZ8c4MsjlY+LzqYLkCZTKE/3KLtRUWVtLFyxcybFQhrjhCZPVHGdqXHotifXGDjQzY6RwuavE9
tsKOUHeLnYT8XPyEfD7Dk/KkwQ6yJRPZnue/KB14FzO1Yn1G9cPlDr6OORtm6u+X71otntiswtww
k/HKMAae7Uzf8L1fE/2H2aobDPgkXFnNQAuZ/bURMSHWmkerKnvFKeOTg6gf5WIVq3+JL+XJ8E4b
HeKuyzjv/Iyk6wqUTDAeq4CKjdJ2FHZosTh7y2SkMabMmPZ6AsfmuE7xzyEH5X586oM9727Uimpv
tm1vqpnnVWoE1JH55gmzClEKebPNosS8572qYdqWzGnVr1jqp+qHWZC1nxnFMxKKkJiY8jMIb90O
67twvRLIS3N+JnSNYl3wlxKcRcbhUn/jW9tC9qavNf9p6OVf1tWH0CzggSCuEk/YQXFw5N7j0i4K
t61gT7IA8srm2aDgZA/nJzzxAhOaCFvWjR0aEAqx8r4F8HZT581YdgbaGkGPnIOCTqeUumFbVKPw
Y15ephCYjdMsIlPMRS7jyYmltqil899v3euveGXgvvlichTPFufcTxJPEh7QK4wpagdvH1KKSm/o
szcRNhkhnbXnC2AQEo0u6Y1pbZ95yegv3HJqqMWP7+ShEly9z3LxfKC8ii78xELKzF5YrEFPZMPr
ATB0zKMMEtfSjeORAKv2rQTx/YvqW1SGFYKZwy0n8rB2YXkTlbYGKys0d264LH7CRBwP4Evk24A0
HdikOg+ft0u6F+joQdgLiAmY+e9S4nRi1lJYzo+Zmqc2ZFLHvBrhK8EnU0OMnCebGT14Qv0SIJY4
dP1OBhJS3MB7ewhBc2JALKMAHMUdVkkByDltW9sMu7lr9T5YZQt/uNu7bq+y0tSKTFg4zM5IjxCG
+HGxZQIAg+TGthFKINQ7hUguxTMYdulVxYsh8QZcXl/MoPMHTYxnbVxQm3qTb3UuaK0r16SRktdk
IMQhAW2TNj8Dve/j8VPkJVmcK3HgvN6GHtatqiK7+r6iTaX3wJqrsYZNV1MNOYxOhYkGw75W+sqj
cRTTMwUFFbqfG6OuedHS6oNumX6fVM4T0eSGEHOGuS2sj+uEn9BmPqJC/NK464R7AjzLfD/JWJk5
1RvNckyz9ZCIJOLFikx3JED1UyP0PBOoCzNe/f+Fk/Vw9g8dmNwi5BzMyQ5KazciShI3Nne+Zk9b
utDsKMV4JV/qM69wptLQ0X+LUi7x7pgzIg/vhiJ/171ltymEtp5W0sFtLkn9/KrK4uNKQsjT7h47
h+zx0ewYXW+ROlKmf3mOerLWeVgnQcaw1SSKQv+pOQXD3981SibHQwYy9FrmLUR+3P0x3kncB7go
SWUJ3B2piyPwZCk9zcdkz/PjJJrRBVZvsG+21HA87xx5hon8tjwuTUINx6rm7CxH7zADbmm3d00S
vGcugSOVoXldrffs75SMGXGDz5n4waOYUjkrwjqPlT80UXqPt413xd0Kh8A5eyqQ6AXOniDXwEmG
n1o/C5ovT/DIs4cwEN0DKFRbcIs92DaPa+TVPbFgoip8cDQO//ojoZ0mGf62CfFdvAJ/y3W1kkoH
7EDgcR7w6S/dH9PJ8eXXGcJ6VqRAbZ/gI2fEUHCD1WZfpsC8X6kTad2+IL2Uie9cQsjenoNXfTF2
py1kx4+FLws0Kin6r8TcIS5v4BeIYA+oUuQtxsx172vzUawLBtDgp7Mbbg5mWds/cRY/dF9EAlmC
178BXarwHEX6s/xY2x0S8cG/GDkYUqOycougzr60JDQPT2m0e1YRaZ8rveqSh+RK/yTmT5CCn5EX
eI/jGFpVnVUagNn18rqJvZlvZNaBjBv2rauMwXJ9ELGOfNeLwtqSqbkL/UGLy03UXMm7STjnMqiu
/CZ8pmnsCYS6aJw92w+/LL7uVAc5fi8IWBjn3dxZ9kC9oIbuItxzNR1qZdad3MvXIDQnAwTvdWd6
3Y53QwFETO8YoDqXLEak2/H15X0iQiFAv3/ZV97vOoLj91FnZKlleyFuOrw5NxyMqg1sb3AxCDud
UdzRYD3ydROG9zNeY7w6sUEd4cRAK3D0mTu68MAwTc2gGRxAIUxPF7y3HIcHD37kr1hejaZzbxb1
szTi+YFdSKzPtzp2IYzaRKpBOR9zX4IIvqvKGdGj1y9XQi91Xbjqgw0ZrWIsUALaGkvf/vAO437U
nBsvvZgQXzt+0V19Cs6K6RvCS2+Rv7RR1eghNzr3w60hRXDaPsifjaZwzM0zX93Ww6aiIuhEkzT7
GE5qhzQoy+0DHNaepGxLckpuc9+7T2Bt4vBwjHrRHDPWtlWz2XZazavblq60nlIazH7x8+J3lH8D
UCl2nsCiA4ZBwXSHGKfK+p19X5XvXwq17bWuL73uyEq2lu62Fg1k3tbAJm7imiTxNp4uIe4jarH0
uMzBERu/VYSjeOq4TJltJNFyadC5BD0oG/CbXrt78hP05pVZWV4/XIcZPYTjjRojU5pQWk+EpmW+
Jm/w6/lPw1OkuGosHSaKwsnl8v9Yz/GazmNXIh6x1oWJR8hsP47e61EeQW3M2f7DjSA5HlVAyZt1
O0vAE5BiRes6NZSSPyuSqEwMCI2ld1KqqusHkK6HzY31CouXQ0A8bNVwtftu0KC1cWDXoR4YrXCm
N+TWNqOFqdVBXzVXBq3Y+xrZnH5Zaze7ehzb1VXWoRcnw83429UfrZodPVMKheysckrTxkyVhR2k
GKgylUsGZn0L7pmQjFGHUon71DpSHoBvGSv8mHCZUROkWd5x1OWqZZNyer4Amg3Ny+FkqxGixdqC
QoOMab4xhu55+V12fhMqoIoG/hRbpv3bsR0FGbWaO4qETis0vXdvAOnni7vfNpClTgKmme4ehPgp
YiSSGyQ3/200GMQLTMwOR+tp1yQhR+yk63EcUuen5EnRKMWWCVN2GRQkw4F7mrfXlSjItrNPuGrt
yb2eobnMrKkZhs3Fgbap1qJZAfpqMadVMxsIYULJXO/KbXQOumBwNJwH89mAoOQq1gC9HOnt8gD2
3vGQvJF+mr2DLYj42kg6xjB+yf6iC0RjW4N71cEGMqiA6YWuGPDT1i8bL4zn72ogRmXouk7eGZoN
6XAdcks2N6V8dh+qvrW9l1odnj7qaAjPoHidnqjemYeS2oJl+ElTS8RGmFGBHC9wrHbGGCaKPIqW
O5GKc2SsWUdS6ngNiYFbw94upbLdIo3TDCLN0JE0dTL9ER+c8NjA2aMlE287GqAUb/jYp43lWWq+
SAqFpCYk9iURngBQT8lChpA9A+UVWrlfKYIl7dkEghpvQdygX2oipMu3s1LuiNWn3a6NeEdoVnuL
A0M+DhKD8pvkTTqBX0/eJ4NzcdjhUfskSX1Dl1D8L0ErsLFigRkjwJ1I1o90eyoOqtUwiqQoAoki
u/HW3dKVX9iHKU14WMSPSpdnMzPCkqOnOnu4kz6E256t13QEjM822fsgGJucW3tvwgUcLyFWaGRW
LAcKEJsl5bimXqb0MyuGza3a05MKbX/W+n0Xk7iHlJuP0fxg+q7B53+Osd+umNItsG6YL0mKn4k5
PoESUZv+sPKgSC536mb6rGWuv6UFng0bdh4b3Jmuwx3xsoGtfPeqCWZZMeZS6ysatM/k+LuEDrdG
Puf1C9R3qdqw4I7Ehc8m9Ot5xq/luYpC2VwKhcQVYUkPT60B3xwNKm4sPR9rDURbIidvIVT+7E8j
FP0MKTPeIlu6E7S8gaiI0pQEqx/8PmTVOrzXd3nwVJY2co7v1kKPQ/qL+TzEN694kYLWpYIuTr/k
cYXObSNBtg9LBZnZgJsHog1ENr8yYGDUjJXu6YKF7+4Ll+DRj0XTItr+son/cy2xqderZZwvt83J
yNLWTJFbSIrxCVR2cfvF5FqJ2p7wPRFmSD+t/DtyNReneulRe1Pzm6+5kDdN728WYWXoOLDGy1PB
YI/Nmn6dnSCSPWJ0QXtv810tdyX84igBfBthnKhr2P9yMNxiUHSS9XubaBIqsPrspEZbXG4mRpQj
vMkGCOZKJbiOM93YmkNdiBG6QWX7xSdeZY62Q6ItaWQqKiX3rbch/NRShbeuB1I97Q+uuffnWNq4
EvcBDTaj7gv28220/qoFsUEvB6pbpx55y855H3Q+3btVEfxW9+YLBImFTIo1B8JMx9qIsfHRJmTq
54L7z+kHqaPYRAal3jvVIG5SWU5oERvs7pBXYThhcj0Ajeb7q+VsVYRlFGAc1V8/t0hAFNLE6KGW
t4UX33zprHgs9W0G7+R9rFBlZbwrwnKeMb43eRkte7poBkp/toJ/glzulbjkO7Fc6XWsR/9cL3le
8QRku23IwMKmqgh/2k76lJd7gELsSWwN/Pw28SICE9ucZvskdtPYvd0LlhnA6P8mQblolwxk03B4
zgSjWDxb7q7tBqb8gpY3jimCM7XY/tvCTtQJcvAzsS3lB/3RRYksFzSe53b8Qy4QdqeQY93P1ZOq
IMxvEZfi/k7LEFMbPoOyK5o0A+aXYbuvhbKPbRfMurEDfNxlt0SfrJMRX4sjQZZKasoA9ej1T27E
Pxf37Yam57uuDqxQxg5yPCYsoIHV3TYqKK7oWCiaIuslzBX4be/3Q04l7j6NpaZXmxLjdJCNd6oT
x8GJnBFl4jrE8pXHg89DJSsEq4u+mwkwTLDt19n/bMC0NqKjYhsGTCQvXhe3iajxcWJ63Wzt5rTK
6aOZPguVYT5xKkK9FilIkr4ro4/0pj1oRcEfPqdQCPFKElFkLYLi50G8jUB2LWVd7mEmo71X2xZP
skylg3IF0RrH9DveybTxuPdows7y9PppszNUAEhaCpi7Fyal8cwRqJtQQdZrozv6uTUH/s0tHxE4
JEy54VJLYAPjhJkSkYyGj4bNZ6SQeKMtw8liLn9N80ObI4ArEmSxODx9AEHZ4VueDEn4gX9JWwxD
2gX8jKeeIZz+PNx7fcjdZpn07cvgTwEv2HUKMcU+zML5C261OGZZ52SWboIVDKFk2ajWqP8J9Yii
yN2/vSWZQsKZLgbMmFUDKPTQiLnGDzgL4Dfy/UMlTfFqmfwK860Gkp+I8aczd1n5hkLCEPtpBPvA
KVdNv7mhkzyQZePrIaQaABjoHL+ZsjgnFeVSMaUotDUbnArdp3+auk79SBX8D3N3v/6qf0XLyjOa
VXv7zXQn1boH18W8b38tJu15xmMoY0gY8b2Z/9cVFzlWmGnBNLUdqQe+8ZsG4hI6+SXT49au32Js
+pSJEVDoIDxhbfgiSFGGbPWc3KyywPesyXusu7Cx+t3O2hwvpJ9oQevoeEqb8CF99Dwj+fdcbi+S
4ourzYN79sUo72V51o/7kURhZ+lCBBT39+Vd9stO+VHQcamZpGsZZiplvO/wV5G7DSoDVgSAfgvy
MdDF79lOR0PIYs/AcCKwm1p+ZFx08lDOa+ETni27LHeX5dRax0tM4/5sc7CVqyAO1qQHEjO7txlr
aX+Bc3DObxW49D12BG705quBHtEKCXSGxXwUD/St+LuEPtRzzjCGySab96uTv2Gg8w4c7htHwAQP
nx/1neh1Wx0aFltKEHNlsWew/UDJinJj0wBRm9jqomGgRBGwUvI4vG0PBFR9Un0rlJMvngS4H/Aq
YreByYCuefZtdcHNWJ5kktukueuqMa0p6oDzx7jtcx1lNp4dbAHQH6jQ+h4JLtugZVDb5iIE3/XX
u2bTI6jSp4C8YLEFD3zT5TIIjChi/ldWU5QQqdRzNsO0+q7DpjR+FAajNMw2Lr9wMBRnVsPK0AgU
MYRpt3AEFCPF93OfPGmVF2aKQc3HW+3JuIOUEua6Tmulj9xAxNaUUTRIHddqwJr4WdbtjuskhYAt
89/DDpyVpC+Zi23I/3Ho6vRn6VH+8wCeawBauo7fSANmF+CnJ+4YKDJamhMATjAHeE1A4FyZDGtQ
T80K60EAtnhsB5gA5s8/qrKWRSzAuFIZo3iByMoEOWqygKm8q5JqazcSa5p1+ncWfZo43NVj+fVc
IHTjmLntSmoeB51GEonoqBHLammkwydUNFLFLEmoOs+wckNBvp9DY+JPxs7Wh5LZUcrluWoYyWq4
pQ8iVL0s0NPPUobzygB8d/ql3rA/J3IoOC1gij0fkqYrhPScn8guuSnaEY6TeYRXZg7unIcKyUwU
nL2XwMgzeG/cm81MMNC51VircOKI11rw44pPKy6cg8J2/C3sjBoBlCNjlmuQkIBCkfsSw0fMGoCk
BZgFqXa385lcH9NNyj3EbtstKCMZy6T8GrtCkHtMl6jvJyCvix0av19XPApTx+k7rKynx2KnpH8x
IjoVYMTbLN4unJpNio87yupWHUoZJy6cCUbqSRcEAi52llmQhiM+ijfYe05CdjwIlA66mKqJR0+b
25EJbcGDb2pk6MhsO8sYAeA3BAAT/SEHz/n88TJkAckX3hAlU4wk5fXzE9nvOX3k0pXJDW4iFIuF
W7Gq7HdyzrYCVFJpvdFu3CTdDfTDhWnHIp+2Ib1+C+KtOeIZ8FPBvX+xNh8HpxJzAefLxS3rntOt
YKruiTik9pFnMkSskcYpf1HoOa34l+qBlvqJJHFRgu4rlJOpKpgEoXNT8XuDXs/toTk6PFy4yK1K
BXqciL2KtSy1W4c7z+20MWUXn3C8WwQ3gYby8a/cE29GbthfPWTCbBLgtvSL2FrzJQyUbiqBwtw7
mRa/vrwjRKLu/rdr2P/hEopvouwRu+sSp7ptie7z52mmMz//Yx+56NBRYPTkYQPLiuHaiiAlAPT6
4MARYu83kc62Pz7hHto12fzSvEsHhUoYzwLGMBjo+DlPvtqBlEDEclWqX3wC2JW/9emg4CPk2qD0
rIeNOYezJtN2wdsAG2XT0HcwAvWa08EWBREjO+610mXzmnqIAedEDy4j2UoccOHYNpn7RVoWu2wm
MiJXznSWgNxlxOV8j6qJUUeHJISrZoMMKiy0CCuo8qVAV745F4zUgY/NoU/Gw46a3Ye6zn97Oiie
2rlj457dK9ccRJ6pGjHEuc/f0S7sBmnmIiD2CDtNBhl6nHe/2A2QgSbVd2oG2o+FNwUQWZkRzGIm
Cke9HPVGY/g4F+ymgYS64Z3XZ2nf2JUOeduNqyaoakpWm69ZuwsWiGXKFz8O+Ds2R072THhFi2ih
CSl8AvVQwWXlN8jlr7WsSheUK7OYwds+66SMvXadDeS6Ce0UjWBCOIMK2Tw5R4bCAnJCMBv9UxVm
RF5uPn+f4un2KVCOycUZuoD1OLFdXyksYi3pb5qvHysvqcL4d4qV6VuJvLQC92lB2fJjr7J1W5py
KneueCTsLD4eetYIrThq0BgtRjV4cEToiMeLEMN29TPbNun5Vc9Tnp0846dHy67Bmq+2gbgHLa92
UjM+gMZ3ccX4E0xm153hIHdBAISml5SfV0gzPSTHftDNds0bdxHEGCvZFm7PZN72vhY2PLWvHoE7
1Qa/a+Q3qlOVX2zrI0MSWQbowEnJ/vx5vs03qqWJeKlXt+f5WXsp1yfCUqUZE1tnbJulkq6O0ZJE
LXPOEkuw5A7bMzd2WPwzXxkxm1uPvtbiETt91Vh4DKiX1rdmbfkwqip8BB+vzFvFgDIAg8U+6vjG
fSOGQY/XgeOnlGXbRClmwjiMWdw36PFsoern8RmnOOdtC9T9smFjALhZimRj1lGrJBvqErW/kKA0
EmAypj3wUNl9JNS5G4nTfUXldfF60m1xrwOkbHWeSOZTgLBq2ztZ0OlW7ipx1XzNuR/W4iMaG8Xy
G+Rfp/e+RIsI6CwmMAHTgf1f4A0bRDfrTaJ5f6890BfO7+3EyFX2EzBGY29BU3JdpXlKkOQCbPnn
S388UpObd/T9mWXfB84tAcmgrknqzb6f+E+ReizhlScLYWvEqANU4lBbB+7H5GMlH+tUhYODuGK1
p+J69DhpHucu3dGLcFSuk8OS+h1Fr0eXcfg2aFroQgv+dhRyMMZ3YTu7lW4DE6CsOfZwsjZ7n+Me
60cU2NIII9n1iMJgGV/EpKZcqSvCpm6bb01s5romTHQAga+78sDPcVf1q17A+y9WXnZESUkRGUVN
0wpFS06Tjyy2fKOBMwDZJWwzgAduhHNNHj4qJ8lfywcUrko9NBpOzp/af+rwlWXxoF5SRgn4Rsv1
/stEFEigONZEXHUhjCUs5MqHK42uP9Tvx3oD9lhjDeyZhh0vdEtqDgw02cd7h4MugpBh12pizt0T
E4DZmEPTvjGeqolvQb2S1UUulqBWPb8sFZxuah+pkfXCKXTE34M5DkcVwphG84jejz/meGJeN/+A
djhGB/JBtXVQ5GEzgO7/YaDXnT5IWQEWTDPonKe7QoHgWK4v2cyyWrk7LjQ9rsffI1CxDfeEZ8WO
dFYAD8rsNbd9IfcWPRJBH/hwFUE4i0EEEYXDkljffe5CxB/QaOcgAHyZ3ukyO/sEaztr4jpB2CO3
ioxfoVlnYTXg7f9eddkjyAhtPLQAmmGxj3jc6dMCJ7H7Ky1zre6jcE27+dKnoloVxJQzbx+xuqQz
eIYwGy8/NiejAq+WmG1+fULuaOp/31/zUxBim/8ZgmcdJGBRnc5KUHr7DvDt/GQ6OB51oTNd6LxH
N6a2b45CRnivVZI5GJ5OCETn5R3CcgCw1xi1MR5YS2eQDnso5He+oaLh9E4ui8rLy6W4HsUfneh5
9IHCgVEFxk8VMbTxgFryWYmjuDm2MkWW43U0dwxdFbhY4/mAAUk7rOeiRrXPTomItA1yuMHd6H9V
QLJdOlzF4hLR1K8TI9sRX5m3Maah38542po+0sfoSYnFstlzke9LtvBS++DsG9Ylq3owZ8NDWo+X
xO1Av+onqoK62XojciRiGTuWrTrtWo7GHoIR+W+Dn+r5QMy8wIYyZjqWK7VpEsQAnEMC/gxgy4qu
HNEGsuhs8ZUY25jzq3aESoyZu2YHlzQlInWX9vj98pGtxQotzB6H5lc2BXZQiKIY59mNaZy5NTdQ
VFJMXbIeSKV4Ya3vWyC3Ly9gP/+leyPK1SMWfEO1cai3Da3WaNlCj0XtFHfcz1RhiWFJSmgNrJ7f
37SeO7zjPCHPH/XEGeiVKy/wAILFuQk0IkeWC25/XYYw4inUnITfT5a0H3Whex2NH01HNZcmuRtN
IG8MMTSdFWrPnmqW90ecv2EQhG2sKpklXJIYCiQdr8HDKJ6/5T6OI9S+XdIcnAQ5RKu9Gq5e243I
dHKrE6gnWWVJENZG6jQyhJ2694vDrwLzpmRVgToa8zR1AJetgccDYS1Au3vBtScuTVn3O1m8Uq0R
jJ6Up+4Az9eGR4mvnD8itENvgdOPoj5xcd4bRn9c25sGGcEgvNpW9FlOXibj8HhIuGTa9+0SaLcD
ZaJ6KbmH2LNP0MkwlWMz88CUvDwLPXGxgsUrH841Tp6p/VXvalikjINM6ut2m6VYd20nOMHPI6ST
/PpYmZ9k1kGUofFec/N08XhVVqvrPTAttVrjbcGAUonEz36fbnPkGtHL9hWh9qf7K5T4DBHNY+3w
DD+RlAvlHzTViTLMMZ5iLxni6HWrn8h+eCanIh0jN2Lt2bKTBw6LJb688CYRLD0+ZqoC+tPjWNZr
iO71vwkPXxH0zfwMLZDvYFAoLXBodIvJVeq8TpCcfmdq8M4eBOU6IS1g8zRF8oT4Bco6ke7u59JX
Ttng2vJI+pGUtpBYUYlkESvkFXHNf1FlGEW1XCME9xnoPqME2PSaSLAKY1yKwBpUjd6smLkYZV1q
ITjqpcW0V4qcsC124CODNAQ3qmjA2Q6IX511vru/GY8fvSHmZChD9JPFK9Dacc1/37jbjyCnIXQp
ob2duHPQcPs2x7cJpuJtGCTywSpm4J+QfsDcH2A5FMYnxJ+mJZWfXj0UzJmU7oilTDKm6T/Y4nz7
8ozfp+z5uVXYnMWlAjqGnlw3ZpVp4NF+4pFY5Xx49IXdqCe85ejvuHVZCc3t4jz5osU9WLs+XK7O
lE2ul1FXi/8VTCjCJ9lCqNUS4OsW10EbJ4KCo3socfXBRcM+LKlvF01EIqlyl0J35/z0ymMpOxOh
jxDgzEugFD+RjxuYeIav2MpmnLBPdTdpIqHt46KBhr04ORy4J4D6aatBAlUPJ9xdJhy6sid3KmDK
Wdivoh8knBaIYgGQmR5NtuBxeX6XD7rg3JsvfrPHMh3ewsJIovBpfA39JRs6UZ372gEAWHnncCNR
eyi3CmjvYtnqhP1C0mIxsAtR41kWMD7kn8UQD1CGwBN0IxI5WkL/iGHmXPna3kZagalM5oyyCcxN
SFQWod/TKUMoW4bWvmV1dwT9/oeO7faXKlwxfRAXZ1cSSS+lCMnMuidYdKrEoXhJKBdQ47CeZzAg
3nj63Emp5OFWUxVKpM0YFSZWcamWNUnHMFprmws/GwqTVJssyB/3XolaFiYN5lD6JuHzjKQSHj9X
gir71MHrTlHwJmjmNGqv7k05RGcFnTIsIp6EJcFAVbM1E2QJYAlXBhy9DjLEQcSKmyHKNA2hDlfj
7jagWCY37ZiRdeM9i9Gwgu/r7iyVG40CA1mmBb3Kt2rK3sbJKO/ywO0mV5KmF8Y9X5KsukIYIJaE
rzSGCGlbtmzQ6uhySHxJ9TTtduR3SHWW03a68B5jszP/aa+DuggmExxPaQ883EbSHcNlkLoK/eaJ
t0TuFf8UqjHaB8Dfsfpt2sOP/R7dPCy/lP8tiq740qACdCCq7AkfMbAPBTTIjmJnNzGtJJ2i8LVQ
ESstTMuypIyvb7qRBSx/VPHX52OwmFq1UXWdrRTnp/Aa6QtdNVD6M8W1dmOLPl2K1nF1EMWSczxA
N9fcciSFEwcAkwXNIUnBrqDO7aNWmJ0GNj1GqPSlMY/vl78NCDh3EC5uCU8Ea3HgQsDg/D3mCpdK
VQaTZm976sV20LL47pisCi0VVzRbvgRpQExPWB938lIAxa8sw541BGBcXYxKk5iLV4JkBzKqu0IG
L1YkKJzrVoBRUVK4WtvXsiSFEBfk5714bOW+8x2VdB8EW0OO7QmOYJ52Qd2I19qfcdE2rxUZuNQF
M2DhjrkeJyymnIOHSA9WwcEVCYYTNHH1HzMj5VnvIjRYs+nOrmKSXhECbO8ac9x/p8a0dlKw/uWH
Yqwhw7leZupaRIYg6te4t9u7+j4tDkV6If9DPM+feXlFi9fU9oauu3At6ZkEI+rgA37WbOXMZNgJ
ZHNhGY7qxSpdzb0uxKv1RrTksq4Tyv5NpUXlOLtzEpgP9ivK9AYnHsyXtled6Wzro508iN5plEZt
0W96LrYKC4Mzdw2procpGygUMuVm87dS9GHcZKKRQistTO0j9DkkP/Ubb7SZtH2cMRrT298TR48t
CA92lx4lz7Y4QItKN2cB8cCViMAmE5riuwDiKDiTN4WND5IqJtkt1JfbH6J8oUCt9DiQytjiWCqR
PGpZnlyxpFnBMu7rm/WCH0tX9lNKOBB8potTM0yQcZHnnuMVmGdPpp5WIXn21WBVuFtdeDhAIsar
lVYovj/lV6YglyVGssBystDr5kzFLzKuH8QL2V03bQyGzWxwgVfxfZ+qg4S6m5bNz3xkn1vccbKa
ItdrBpNJWnXv8XVLdwAxOCRYjMnNxzlTJvawmlS48GHp8svjk8pm3cLasBvkG3ddbKtKRUhSwioe
LXw/aiCD39iCzfRz+NOE+IN1DOaR3gIj3QvcEyOSR9ksrTtk04DA/oI0CAxGrkfhol08qC4jc7ha
mfqDDcKL/SF9lOZX73GRrZl+Tark20ltdjk8Y755Im3nf6lMFzKtyorAngheriwAPP92cFi6bQKl
driEVOIIyhUojLc+QdBzreXTROxrUscEm4QeGE1BNjS3O0ghLuMbGvTlcLei3vVLHlztLaT42HAa
ffg1J28MUskTJOwILnW8FhySGPW4Fq8F7s/uRg9WfFSvxLuXY1wzFcfepFF94e7ojrx/iH1TN1Fb
qvgiEZzYS0eBLcBxc5FPt1i8DH3CZ3NALt6PohMTDrcsrQDoC6n7C+50680si4z+XXocOU1nZh0A
38yN16IJGdCdLAi/hkmky35+xtEOKRid5n9d109lb02C/K9yKuuatfDhcevGmAhYwdBf/Y0JZokG
ipEum6yGkb7z66MltwE3XDzXnOfupA9vvxSwU4zB/t/gWtu2BFLI+6NIynF1qGV+k20K7FBKmDGf
gFo8lMwHd55qTb6CBh6lIiM/ZtRoSVUiEMmwVBsUHqEAsaUtp2p2gA8noz8AuOmqA9fQDXQkoTEa
d5cd7okhZ31PTTrDjuQUHkqyiW24EHs8Tw1H8TsRIHeEiwKqSLEm1aI1RHFFvbVV5H1YGJb1fgwV
n82vC3NTaY8wqNSeNXtH2g9KvNzzQivNxLE/8BeVqJ2ONHjI90gxBEV5e1uJcFCmehee84m3H853
ab5TNcklc7/i61BlK7OfwAZxvMociwboAiNrntlgqGLYVlwnE+IIlRfgfWgPWNo9f4nA5GMyk8eT
LnrYF6i8FedGEs+kvhlRrk2ujgdMQZTBkOjNNgkw1F4+jRPv/AqdJcXHO9BmWMPx1R38hxEdQeLN
S5SbneRz/7dclPhPDoaZWORzgbgZral68IQCrUITTkbpscOeaUNkmx4NKNx7LWR1OAwVz+fdZjbo
L4Z5Poscm+Yq48gQR4GmxeWbzevPwosLGUTPUGs8Nq5lW+VJpXb2AzvQJsnXz5VjDeqpbxhHKZ5b
QyD6Jf7CR8bSzWLZjUqMY4QXxNnBjCqo0LbNejhhsYPCEvuQ6sJ7YdhHRLSIxT0bQngS4kQjP3Vb
fU/1mppOxFMZwfoYcusDKc93DdwUtTc8D1MeKxg+D/6yAfgCbTizN/8PwG7JLTGMy93Vu8NgEa91
VrfGdEy6BRhX19tc2v9LGzptLED2TSyidwTfL9MZMviIb9/V4DY0yKEq9fgXtgdYa3EokRoK6iK0
3qo4wytUrPNR8e3GCe3CT/p1rj+JT8RiBi+RMsC0UAP8bqjCtBs3QVc5u8X1VGkKiOULgbPM+PL3
R4xZfsRmq0HidWUfMBI1Cipv4U+MJeXMS/dovmcxbs9K24TDuFetPvKSkQkFFybCUD5Lm41u4mQ8
hrAikABLE+d5V/xFFgB7pvy//dtjECTFMwa9RExmPtDfnTZRvQTnoThCitrdEX96wgZN8kDiL2rS
1hEXyOEZFpSO7DeZGMK50ybL+77n3U1Iro6Y086fo3LyZ1/0ZQh1h/1Xz5gW4ucAGuSDxofr0OH3
O+n2vL5Kjzk7p+ePuIXBb5eSGA1q2HGVg3iDhx90iTbQ7NOYOaoszkd/vic/7rKndz2VvQafVhur
WrLpK0iipaQ73fvQjxYAM5Rg/vuPBiWKAg9ZOQ8L6+QwZOBcgyhOVFDTqGeud1Qr+20vk8Ydy5mz
Br+MPedTFFtaNWXnYnRa5187FHnRGo4iOBIWqCN2VgZOlifL8aS8y3QmaLxEuK1EuHebRLDJln+e
ksRIRZ4h9x0dR4GFAgNmM99dyZdQJ50U7OlspyU74PiS6Q+/3Fea0k+Lkou67Een9euK5JsRiJh+
gTODDzLUTAO0dxXbw/dlEwjP3tZJxfQOaYQa6654GUVIpXwNWnkjVh70Zy4dWiJHBAYJdROb/lgh
frPuUDsFgZWfdQyjeU7JOuMDc6huTjZrlzBLgO9vUl86mSl6MmI7+jM4uQ5zgxR1x2atYXFphzSk
fOPIYRppIS7GwAAD9HwRrQGEm2t/Xp6P+AGbhAl+d4R4iYp6r3dSZlTWz13T0LHNJYV+HNV0kcQV
aijxARK39VLRbOP2lVBZi3WG2fEKdwXNpL1239BiFTcMloOH2x9Xq1AAL4KYLB3BR+WwHve0Yu6f
eiWW36Y4X1LfYgNRe06iQlTMwso1BeT6Kv1ahyQ1usQbn/tE+U5vj0/W7wCZt8gBvnfyeQCLnbyA
p63i9cdC/7kiwrWHzTJhecCkyOtMhfhpBZDdV0l78Iq8XL+JwCDMHZY5pvaE0UGoAGYr1Y7sE/o/
tKqIhVYRfoNxl2FrDbXCHhsIt1fA1xtBfg6J0NX1NwIFg23QUJjipBABe1dQ2dHbSBFBxNHeZH47
vkajYtXbmtRkaTN8j7t9rUYCgfatz1flXDEB3L7wB/njuYDP8wmsmUj0B9RtG3QapAmRm/jDu/Ay
Jk3nLMf2Tq9K/yhAdKMHxY7/qyU35avCPVGRcBEbIZqyvArk/zKbh8wTpPENvhUtCTRm0DOIDDsW
WJs0fR6V7o0IOiJGRnafLSLMFp9Xl4RigENqku/XafWXTuBzozoI9areI3S2kLhyoRhvIYXRDbHx
9NVPdokcsDWrpg6ZV7yres/JDqx5HwbfjwWrdPg1o6uiaTIsnmiYM1kijk9sSxEZaJDk8TjOTCEr
WNOB9ZEXNJXWKx9sZOInO9eXRw4ba2Nw0z6PtWUOlx0RqhpDuI94QgPY2NMQ9cW3FyQsdcMlWARi
72bUa8vVzDL9WWS+fgi600PQv5XBha1fzbm9c6PlbAV1ZreBrySGtqHKUSLJytvRy8niO3qjhyGn
iEUAejBG4QeJA13jSK415hgLCa6ZxGAYYpp/1ayQDXCCP6IdkXfnCI/0ZCT7djqWMRKA+EwqcGYW
PuaAreQP4J/FTbjW/GWVDQqVZE/LHKwZR/4Ste1ooFG+YI6HMLR4R2QBVpx2cn+vM8m+0bciq52n
88/QtEi+g90aKlmFE+VyHU+1WCIUpt6PGAxc7MXNw6YqIQL9OXwi22hORphcB6krhJm2itfb2IYs
766Kwu0VaygSxr5yH/PJOYNG+TG+PusalvhHpkHYnPIQwsq1H1WkRyXrsutXQc3IuTefvJ7IahNO
sNgvUtcVCNgpxl5u9Xoadoavr5evGKtCmnbcIRDyExUITT2pCgmyaUsI57MnyFZFJBB7eE1xZCtr
GHy1fIXbdn9a7AP0b+jSShTpGc0jP4jpqzKgb0tfIsxLidosmwMb/GKkuXyLakO0lNIqDsPx9Uyz
C2pDxH1b1ppZd0NfGmJloe5D2uUhif074VUN9XxcYwVKiSNC8SiUH7+A2ItoknVVaWc1D/0qD9QR
dhsfZ/bQClRVUsV7OxqApiDMHTSkt4Viau3nRRNe4FKP0QmWlwjjgQ7MgfDSeDrATqypfLXrEnYh
QI3XGRpFswTXo4zGHSiHN77FmH6qI0eGQnlYu5Vkwdme2fA44e/k7pEYlr5OebN4H5sOXtgIRc8j
dSjdGhT3epWvURzaE9RMRmoKGjLQA7WKBiduwtzQGuNHoBJN6X1XX7J9e8Kbeh0rU4goaoAp8gam
X078ptelxSTss4AcSbHWJf2cth4UOdu8ndf1wM9JNZAIqM9Io8T/QQXaIZUKlJ2uFZMS12VkzAeg
Ehw9Al2uYZMi4eCs+6gsg2JR/n+bG/D1cjaxnQO8WLGg1zLf33XJilBP3HThofLQJMf5oYETjOn9
lBNtBMrXw4x8KGQzOhdtHt9/FeWLbILCPFz59k+wlioPT3b+UM+VMhTt8SmFkXau+Xc2Mz9L/h5R
tiIGM4/Ps6QksiP3BmQ8Fei4U4jSttcfySE0BHYr8pFwf6GwhS+xgpvP+MwOJSuBr5YzCX7B4Pzj
aK9K+zHpDAg2t5rL/+PMM89sXgmtCRYiiX4JuxSVhamt52kop3m/cm9RZFPxgqy97kgVFVOv8hzL
Tja93cc/3i5hm1EwAGTiAxiMyzkeB5RSxfdOzD+gNausQn+idPalTYehVAxz2jrHlA6oJDjiPRt+
MV87uV/uUpPImH0szgEPSIKbMhgwfd5suT6X4d3V8jizNoYz9Zrdi3ATrRTTmBN+isnaMZ5iVSfs
sszqmV06LQYdh7iQjVwMuuQ2+iwO1tZfK/t5pP1RAnFk/3HXH3bCf9r1+sWGbepEplveQMC1+CR2
wD2sRPK6fJricB42YpjVRn7G30xsu2vn9IIGsrvcwVmdBxnTAsslIZH5cei69xaaZW9HrXl9p34n
hiPdgdvYPOUi+Hbc4LN//sSxhDvpvedYx+VqqrqxqfAiqWV5uotJlOtCbYeZmeCQ+XewbfphzMuD
BrM/hBzVQqN0sXe6IGCQ9oVOLKUiSt0O80VCqcJ0v7Hnt3Bmd+uRaZdBYCxSzmwwpGtRT0eC20fd
tB4EN0hOcwM6OJgJTC6WqXgrd4M0LFHezdFMYCStKUNcJG5tbh+httNVv5irSxt3y8fB8WEhil3s
pNss+imgiBnkPweS1ECvM4Kf0az+E8dSYKnZRH0pRGcc/iZVKJkijnJMuWIoIRkKIMcQpzExQ8Ep
ZUH6KnTtphwPARm/ji5NRRW+GLC9PgGBj/Kxa8m1a7CFvZAW+YunQH/wPT9p9gSD1H1BpHiU9iHk
WBfUXUrMtOmvP2bMB6Wq0oBZakPZZOr71I4A6K9iTMxpcf8fEu4LV2fdQhKIJUjHdDj8HOAl+ZaK
1HrJkncIfXXaDupY6NbYC/7F4jkyrGP5MY7CnROwK4WTt3ggKLQt/H+me7u9tpXknrc8X80LFpiy
kONZecrkNSYNGGIcKlIvfR3WQiyGEUcovc1Ep55zXOGTvWkhqc9+rgMSrEq+kIu0CYvBBwY5t3ES
xcCRrbf/yL9dPGz11LNFLo/bQQMk/nsOr64cJyRdIufcovdPJrmkA7DeQGOTl3w0mqAuAcmXOAZ1
uxoifXtEMuXGgjGnqnYuya6Pa6vC8qEpSP8FUOShI6yktOdWblIYoX3rsflm/+oej5qMfd6H4qVu
CxrQkT4q2s4BLKbtA/DkavtXOWZAnJ12GlfA4/p4zntIrMpQqJt+5brWPjZVXtMOsP2p5HIrDCIJ
Pa2YX/DZ406YwQMW9p32gMlkzbmCxBIHBUlgLd/1Vv7EYpFzKoZ+POyrupqlF0v4o8wc18Z9HApn
8dnhJwKDLuVcP326T/FC3fLTnqj+RWr5VchmymPQ97KR8qsnfHkvBXsGeE/vi1Hx36nBjAXEXhCL
uuVFbWMG9G5QZsUqSb53/jebGRYApIDpOnvSWh8OSShqmQWopEJoOjEtSXhP51ofhQEWvQ8SS5J7
TAT1bK5/iFq4kAjQuiASOBd144hOM9vtbkRhlxJo7vXxpv+uI5C73w4E8MbMyjL0hUreRvic2598
qNkI4yBGHLZh8HpPEhPImuU4u1k90bNMUTo9Eoug4h39uSyNZKpmNqoQl2ZOZ01cSdOkjOiTz8bC
yt5wR8Zy7LjYfYqCi+1tKtpVu6fkpTFP0IxoftqgmdFE6TVc/ytHTFi+4TymRdZKFjlUKawhdMK9
QDG+6B9X8J8Flc8w+g9lhzOFlnxDiObz+9b64VE5x1p782I1Jiy+KAL+tAwandNA1bC7nV8NwKHZ
uz1NMdfUj3wPzSfwcyIjVxOZWL0++/jWBOTXzTKsi9Cs0qsOYoQpsFSjcKyX9vX/GQvvVVoPLNNW
zw1fnfDdtrJoH8JFnORY9Kkc0FTRHvMPCU5ZNG6NGL28EQhiJIVQdMEVGMZSrubwwGvcmdArzOw9
+CF/tDanbzD48BIuYPq7XUOXeyTzdHE0N4lB53ssYdPC5UUY3Srw1PZaLRkQZBpOheeop9E+Fc4+
sRwRyz/cbdGEPy+WuTehLz7+OoEWeTVwq5vCVEpXtXoO27/KWi3Sbir/W48DvTIRmvrwwyxnEL0S
xC3fclQanvn1QZ61q9lbOYabeypWVikZy3ZX+O6FudOC/IvgMsi7Cr/mEz/oK8Htl35UOt2ukRJe
nYDrH2F5d8O0XfyGPPfO84InDP4/eRNmyJEl4EgnhBL4H5MxfOT5TssZ8OJTZB4zBuC8akzKHocf
ywAoM2ZxzsNLv3xHNZoySkRRzKDWm3wWtYBi3fdB2qMZpPVqPoQsND4V8e08b1XjmlNRmvw9KrvG
X/WOi9f5TRvsl6YLn89QphpYF5z67bskCdmfQ2gg/ub8fpmOydRpCHiMpo/P/8nwX4jpIx81jaFV
wpGUtYA1HVHlp0FqeHl7bI6FTpPNR25N/TCObWqiHaX4xnrtLp5IzFn+8wVEeTXVTfn6IrVttfpv
pGW1G1thS6WSqqo51DZW8fYDrijKdqSaNcdgFzzKO8qT6IEPQ3Pms91a0MLzhLgNXTFzLtWZ6OBb
aRrR0NuoXYErgHbonqQJLvQzovbJgrJdhujzgk1fZ3c/mE7V/1tFfxSbjOTwUK3TmkTE7qaDaysA
9+6jASgKAgSQamtwUEDgbvAE7Xna1qZaJk8nNM77KzzkbAto8mq8cRBzNFogQU8KJrkwWsCo4Tj6
CkweUJp569Ovn4Ff1v+otArk4VXbsSr7iRmGjsu63QpdjbF433jUEtM54wiGvdli0N1ZUyCSDIF0
eDnMqn7cXbrBx+CvVS4314VipoH0n/pnnc5oJt9VlkF7A+/YstuYgf/QkWKshTQ3GFjRlRQ/jSBH
rnTVNDzUqx9nng1cYo1wVoQB+whrGB3aTCL5Wckjun+lgBgl1sjeE7t7SYj3dBSg0HWGOlj8HM0X
nj9GlCX2/uKTyjA2GECmJG36hcwxQxjFuF/NdMoE5hm4lV+Edf/j+5zuOE7MSuSosFwH/xI7biy9
jyh6Nnc5RHgdeU/WuZjJc+uuSvoI3bjQAp6jZNFaLSUAZ/fhMQ5Z+9psIqaaWpl3TaE5rW274cRM
RUxN00VZaTgFHI5soo1KeI81/QG/PXTMwP5VRc/fMXenPLhwIJur33G1St1WN081LhcjXU3SWBvj
FzC1PtKFx4jkpfsnbbJ5pWLUHITGclTYrZtg0TQ1EQjK1ljF6rMpx4Iv9s3S+xtgcvNwSnNnwPNV
tCIv6voZVu49DMmL/d/JMk/by2D999vd2FyZuoS8OGdmbJccB9IwAvK2FycmAFlWHyNDEqmE3qSg
mBuEC9Y86UuZJRyl6iTE8QuM937M5clKNYZYyojbWcDkUSmJGY/Tj1j28IIQxShKTP13jqDQ4j2G
4XcmRlXdfmmaERjj1QHxaFYHUu1ZoTkc8MWmZ0Q146y/vTTn/aU3meJWezkAhw3bC40UwR0Aollz
Cw8Pe4YaBApyvNZCSLisr+f0Ex7I9yiYNIdkXtXb9t9Gbd1OWdKm94TEOMKBi/KpN4OOvk/9ys8c
ij85B+PmrleteLf1VTrCeaHZR+/pU/FtXfn6pC4bwOrbUmVaZ0drMg4q5AOyzaWTdp/x0bfTc/aF
seLPvfL1ZL98neryevGBOG+15UPEq2x0zrmDBl0MCbR/tUCnipgeExdUPa2Hu9UYKQR+Ux7l9zMf
iCotAq1FF44COmmROwBHUeOkhz9TQMoTbBUohn50qzGS0Mgj8MUywkLdEdFisOHJfF0HJb0u6MeQ
1soIXSX5pXxjhYOgA0b43IWmTx96zLvjPMdg6oOFDRa2BVzoLmN+YAA2RCQ1aaAkVZE/e65lIYps
Fy95AScC1VqWsZKHICEL41V63s1utCE0/46J6bsX7gLCI6R3qgV0I2d0fGFPLenUwZYEW3fX0ivl
hrg+YEr04GjAFyLBQg+/rdowKJQW7sXL4LavrPV0kkM0OvDycrl0xUZpN2lmTEY/6x0iIgJnw25D
/AqOu3aVXdEYt3z/LXnpbvqzGHKD+iKXEG5sjMc1RGrtZEkN/VvpNlUfeBy4/KrpFtRqWN16H3uz
usaEdLAGPNLK7JL2KsVkm689e14kQ8ulawUPVkTToaJdGQc96CY+mPKbZkQ7ruuZf1+3+ryCYoxy
GkTrLx+Kc8+8K5xQPmr5GtvaYh/TBQoVx8uCtsJohuYwOX1orIAiVEQ0F5vVkkXRTOCV+yZNjH8b
RiGQztuPp29CfYRAocmR1il7IrI34Xv6OarwCaGSEh0rerGgT/ZN71k5kPDJFJADKN/G0Lsllpbm
n7O6YheyowFZ5kgBXzMJNxFc6SPIgSNNuwXBhjUBH3ST6wIKSnwVmOxX9Q8Z3Bmw7zpMyJn8y4o6
UZTNB5zNgtWM5G/kJT4RTejUJ198jEfyL0Gtt+r82SdcEExgdwf3YUzE0VH6qxUcg21VInOJYz/Z
8yx4ROkZW9zZMJSWFZZES55i7B5HoXEOLouwRxR3Kt/J65Wk4EG4N0AyERjoztN+fZUY8kobE4Tm
oBG7VBb7EXEBM5WocPYzLRNS2JcxiLy+17KGjrIHizm3jNJO13NmiurO67d76aLBgMLKPSFMrqG2
neM71P77qPQ77EmLmUj+v5fShjD0Y1E4eHMPk189jtIcf+r2xwz31hTMY9IemQjPpNafkfxjNRUn
f2wW4YdkQ/9ODM7qKcvk7OUvEY1D/x7QKzzdtBQ3+YrKsQX2Kp1vG4M0Oat0nsMLpTOIzhSJhS7D
41yaQ8d/T4F995wlvMtXDnJXd0g7ZCcCUdA8QtMcQHWPk1bSHnUYKgVpCxGDE9cOfU36QTQfUG6J
oNTip+mFh6LS6Qz7cYa69ZHxoLWa9xrDUA8j+JofIaygIFziOo8FBmuAIvOoSgiRttSZIWHVJqRn
6aiYTlnFvoBhCP8kg+zpBnCMqKpkyYBp0BS5wLibl02mgWEUBZiVIOtWXYoOGJe/tV0/DJfS/Wzy
Ta3lKGNPs24e9SETY5HD3w==
`protect end_protected

