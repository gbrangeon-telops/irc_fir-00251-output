

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Hz4PNZqDQYlRQ+ken68CUlKtwl5bD3KVcGYwK7pLDyYBwi6Th9L/PQr7ts5tJoXAIQRYcIzRxOvE
bOvIjO60PA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
GP7r+Hw/Nq0CwA10fCvNkrkcgK45iHUPRmPqoCkPDKd3ozfduaGFS4NbQcQDFEPry0eRmQ2gSn3i
AGkmBiS/ZMkSitJxD/EIgYbO/fqPeNo/xyESKAW2O+T1ZwGwXyv6qMAp2gFqycRAbj6T5U/FUq52
EYpn3NB0sMc8yOEFyQo=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
le8HFUmlytAxiraEF0H5rT3qqsng3b8xZZHcvlli3mx0SdV7s39NBBuklCsi2z+U5UKSzgnk8WIo
w7XOgbkBH4I5bMmtC280eEWQOIcj1GSezKn8Kq725OUTUl7WIOM9hdaAEgsyYV4aegR9ufM3pfv5
jM49vFUeG7XEd7xqdKUxYcrZmsZ8CqQuOZKMv7+xnku0k9eaKv42hAQ7cL1uIXuIFvzDlZHyC8MD
e2+jTkJtzyJMk7U2Hncf7jaM/O2gSIFGoRR2sNNwVB0ATLYzGBnoP+wY1MWKJdSoIbDQ5r0792eb
YO5yRbe6PhUe2+UdG6sNzgiR0viGJQ6R/9i02A==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
tSJEOPsqlnARL2Dz0wpm4XWyg0nGSs+Wnp+fpstkJG7juRdPH6snLi4H3YFLGcOIteaUd6+0+nV0
HNDEDrgudSIwom4ffSyyotXElk+U/5goIr091+0B19LyBlVHPMfovruJJsH5yPOjkIUbE3z//OG/
9D90RTj2hDW4+5DRikw=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Y2U+pnaPqDjEYN9Ag4nM7UfxJ44UWPvMFi6W/IpytPtcFc+Gta7bvyNellM8zINHBtaT4/XvwpGs
zz9LduYm/i37u/eaLh4notjKL1KlEzSl/RQQCOAWEkJvBF59EPqbeUalx4NMTEi6gApYczcwU5ry
jjndsvqks3Obkc3R6uXlQHIzKbPFQM2kj8SV74srGUscAjTY98txOVHFhIk/okWPW2x7ScPBZlnH
/p6enNTFgNVy7YICPLQQ9SjExe9hKly0/QrbtcXPdI2+m7HVD28iWrn6JNqPDPmkYTv4lqGhGruw
jT2AigpLW8vV0cP+HITHbLQV7l7eN+9WNmGRNA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 126368)
`protect data_block
9G2D/MDaibnDMNJnqQkLN8+G8C8hX/XZs4XwV5b8DCKtxNZ584TvzPOa+Ks17qmWTvmjB1cdHPJ9
1M3UJM1R7kiU0vP3tiv2bTyBFmsxoizOcmtIj/0i6/h9LlFuUzfQqp0Jjxw67YKz8ZIH/Ho0XT8D
7LnEzPqDMP5CAspiBPya9DvxNQL4BfyaHUQvMfpFkPCN1BYJOmw612dm2MTS0QHsO09U73lBP+km
bk502l2iv7fMc7nPiKg1/xXFSeSqUWKySXh6Gc2/HBGLWObQMnW2onire4F/UvoH8qc+y8wAu8Ea
J8dWaQnHC6L0RdTS3HcmnTIWptyJ0dmczMjTjX+LhAqLLM4HDiENhrCsSa3FsPYCaZQHV4jJQTMr
WyZxPLyg7laeU0Q7hqomE7W6LEtC+u8eZnO2Sg1eMOu49aTjbmpTVqikXthiorAy25h1m3hCgE3w
ryxaJCeZydoFP0Q5bJhMjbs1EQ1JkS6y13u47tSTjCnZF2RtlNDhGkoKlcRhTtaYdvMUr+ml5C/c
zFgszE2MGJYXYeVVoiskXHNTW3YojhSmFKHG58A8CmmKm0LLjOo7rZUckiV0odglFXqeIwR8mjJ+
in6SmQ39v2ldQpq+i16uZJPFaDgH7W/5J5ic1YYysTDJ1nb29p3yjiPbhYL0DReRo/EZ2M9qdXPI
mX9c3cr8netwxC8SocNcZkc0WwWMnBh+Icx+TSH7a4KUqjfGKzRLxmj3WLRmMPPySXiHQQA0oK1b
s73zXuCNN4uMOmxIp/mZbODAdmsowaPqPNZxacQ4x56pg2MgAzwwEFiNWNNxniO5VDsrLq4m28tv
47Y1jsxdjZ8MRSg278Kd9h+DpQodBZyKZiEsJ65niUPoVRKnWSCLVKDP+VlIxCzWbDVJJtlDH3+O
hVsbtn7DLo/E1F3BeVFUbEKyEK6vKF8f+Ygeb8Q3MmVVBBhJVwWMMLflg2fUekU7FY8CxJRSMxZs
Eqrri8TUYCnT/lQfAGt+BFwCsX11LpmWzc1mXPkGyxUgOgcgHD0f26WWk/urUlQDQpPGYKfp+Vl4
HMKqUStGRi8NGpTueIvv0pZxFg5Ny/BX6Adzi6+zR+GQM3DXtUl+Gi8YKHRNS2z0RoLU7/Nb95bq
ZPzoaeJ93ZKkLyyZxqMOjGeQ1B0Css1pCyyWjEQg4Dq8STXjOvaZ7iZS++y/gmQRN3mNuyf2whGN
ITAbZCG886bCRth4c709MX8bQzx6NjISoFr2XLwYJqRJgVeyd+H+sIIonJJ6z/jYSMg3cQwRWher
XZNlmYg2EUUU3cy4fNTDA2uq0jFkyXgev8PSc+REt2DZDO/gPOxSs9v+9HWuuP5zhr4DWFwnCMB6
jNZEetP3aZqsoCzuE5dQ3C+ZdY2XutLpQbt0j3bliP35cRx/SG43XJwgpZ7TOw0kz1YUI1SMEHJ+
FjfHIlpLte5NRv2PriM8jNBxStPv3SKCxamXkV6SiM+0GdkNEwn0lIEPLyiyWyjRSxy9h8dqOjSc
gYeCz//EKSOlumrXdMvI4onGF7Zef3A7KPfypGTB5rsu5pWerwvDZHm87HwHVLIGZOiJrPLXLTun
pMPe0vp+wTE2/OrQJZd2ORTHJ/zjOu2+Uf/UAMSdJo66Fhw8NGzxPo9DiEILFzpnXRz2Q5/79qRJ
tE6GOuhZLNaYAaBpzpRWkaI6ceFK7MS6i18eCIIYtCAVjBEntVwODpXnqu7lvWjX7PWeiAs+pPzg
DVdsYquKidaOzKshQNwVDxT+t+bdnJkD002Zqvo5FJxKe+9esCWDVDlbiYN0fJpwuDMYdwkMVqYC
NPwBDc2ghTMCExpPEyXG0Hmw2AOVEqC4uSjvmqtd8v9h3rtaxljeNvKHeUsFPkDFokyfy/IqYhW7
dHQNqfTEX5scrDGoWaSdUxvAZTjWWGd9Vg0ISRSJu/CGDm30bgnifyXtf6+gTwcCKbzFkNa9ftTi
R0bQ3LBHzWIX/9jObWTW+7eDOp0gUtogB+Fw7/xDgF9ox5VXq4UnBTsgomwYxyutwp17l0Pjc0KN
Rm4qxz4TegkHZX3Y9wyqJcKCNDhlEUBsPgFdonWAEF3iSmUqX9mxHXEYmbEz1Y7ybfVDnv/8aWr6
/Fp88NqhV5ZiFOJPcDvbPQlFlO1yjdYQ5ziLkt/6w2mXv/hf844ujzvgAIaxzIiefcyup1CqQ2hR
U4DvaLeU0yOVys3sX4rkwfNz3WQNWRbEG1WMhlovhspGUcVFZVw0BTAmY8j5X+QsOsiJVzis3SLj
Ltugush0kWL3ws6W7IJI905azatdBZaVlRJhHaFZpHNbhAx7N59Qf8fAU8ZbIjLiVXMwJ7IKQNAo
yysq+AZZJMvqAf00barA3olKtnpBHNSEesIQbg7MBZtTJhnSNyONZRfu7hm4ktWseJeQwj2v6ZaO
OjuSqRXdRJVz13Gu7TIl/x7es6LJEE0p4bcT91maMesnQBINHS3T5+O640xUJ0iizFkgZm9FEpf4
AyLhY2gfODAWq4PJQGBtDp/qmrPrX+hG1vGbl+kWDe7wF6v6hzYY3uxgvCRRs5+VmfhoPiMBGPSJ
TBqW1Ea4ZtlrZ6IZHR7OLZxjKh+R2J9XOAOfZXVupG2fIaXXO/H64zHwZ5ys56QRh+J34xlCbe6Y
GikzXrQYOX4XXCYH2z4Q0GU6HBotEdvf7IKtUgWaLCW8gbx7sV8UMlqnzbqp/72AP5u99aN9oaub
44WIg5KSI7AnCFxY94nBPv+IUxnN8hE/c7KYLb1c/pup0tyFG/A0/p0dw9C/7ZIRhY+lE4pyXNKo
vOiImFmmkbGeB7ojlM7s5hIwOdwI97iS4IdzDzoVRN5pdsEabC75QbWwneXcIszoxG/7AAk70uIM
979Yht6DsuaJesWemDUSNcEomPJ/yJ0Xb0TZU8IRkYdFLfWUN16lxhZKDyZmzl3x0ap7VXFkFyWq
0qGGkojyMg4CwGxo6NEopW2nBE5QJ1KRfjG1UAyJsuMVeP7vy2TMRFrldrDxaZU/IcSLi3ePd9n5
eAWh5oQ0DJjC9tHuBi2LFfWg5GMDWa991o+LqNy/JANA/5sxd+mzbj/AE3N3P90eN3XcBHcZgRF6
M2zEdPiZnMaVlHakbbdDoMIDj4Z70KeLipC8RylZU49qeR5ysZ1RQLYcxegiX7mL9XkV2+rVJyzW
SaqTKAu2cft1EUF+x2WY+aBIyhdzkXlo/nfneUxo1aaFr1SGx0Alw8gM7T5A7l5ZZwJreJUoflbd
qZwd9t2e7n6cddqqBDrVAl+8jEsZCm2I5XVlGzIpI2uYyRo3P5DWXc7oK1fC0Mudd9narr8xdA2o
HupQQffoqnV76j+MeL30cBV5EymI7HhC+7XS815xjKFDz1Uulj9l8vF1Xf72x0orPGNxNNzvE+yC
Fg5pFoHOdqv/YGw6Gtfrho9RiBxFf0hrnSHP1rLmLDmkmg3nG2TUXT4bM0hRRMr2Fe/XXJQmAMPF
suIkDJ4nhikr/3G5aZfTeFtlIfHJpoql4zNAKawFxs4g2WYVKfgV6l3UCcl0dIkN881X9jAzSkIH
NFks3935peDXSuEq8bFTrRj0RpP4xItdUrqCIxFwLS7lI+YWdFMl8MiTIJCnj8ZbGICPWH1Uy+P9
ol9fTnR87Z1AcouLW2i4PQh1QYMVf28g4KSxgSPSbU1FXBp5N8mtx1XtXxmRqGN5Fy2xKR31jzXp
wlkqxkucuS3rfeLSWxIfLj7PfD+xnjKd18WwdbNTi/IBKh4oLQL4L6+bZ0v1AVi7u3HvKMcvI8yb
zRVM0vuRx0VnBiv0M0mXimxQbkgcbYI/PM1/zx+ZJs30bvWKFG/KfNqc5vJ4QPUw11liuo1pei6u
cCV2vK57Y264sUaFwZPk76d1orajdoKxik3PnRX4blhsBH38xnl13VID6NgYvjiLZ1p++JYmgjSN
MKiQvkJT3o0xSTPLKlwdp3hpM9iCew5ZIcDdjekfpsF4oQQrrSjqtest9I2YS9sax212JFuZ2WnZ
O3415JNPIMfZgZdOaqmZJg7toQe5LdKA1f//AzO6TplNyWjZiPMUronWgdoaMFkQer3DM2Dp0cZc
i87XV6Thc0zOHOw3SC9CmjCneUzTLiKEkdw8YbGbZdqYJutHgInQEUXbIWKkOzwYQ1LrJh1FBVqj
Em/Z6njjw+p3gPvaDpjafFK/sDtjtCjZyjHyfFxf2DYqZT29e5lmBI+vxZlurvICkjIrzDHqtGwp
zAQKtzXqwFGpzlFMNnZMzmEASnQwsy6Z7ldz464Seeug3OzKl5/5JIzNFIg3oyg3D2FpGzo2XdTB
iGKTIUuVbRO+zNs5Kgh2jx7U6IuS4csa1bjRcehyrwNV06KqM9FjzozKdCTtnTTCfa5AXLzpb8nW
9HMr+qOjkk2p0u6vxZctye7JQwVD7BvL3YaZI0NE5nPFuYAe/z8yAX6sqBH+P4JMQdd61olRihL6
nZT+1qePN4Q+//9PCzMMlGSAOslSrpzvfqGztOypbO0/gcsBud0QsDbbvV0Qo3KhAv7CanPThP+P
3Lv+jtqaVNaFnR0Al6p0QoQPRbQ2TsS9HmowiDUBi80hkoCdccFlpeqFBj2DFAxPRtFohR5Broqy
NiKEZ18iwz7ru8V+iMQK4FsYMuqC0vsz7z3E2EM4bCH4lsnFzMBB+F/pcA52VsW7AmQZDSXABIVN
ZDGtvp5LxIiOfqo18MQbrmvAZDtuT1CIogJnNd8hDZDlVwgExshfM/a57xZ5gngGX+JoP+NQ+xrm
tlmCKiym0FyWfp58dpNxVXc6OVqz0BAh0lpNfEZuMfw1pGV717WpG2YUv4LW6PtexBrsBWMXgBu8
sbd+L6lvI/Ijy0SAIXx601IF/KHzHTRLH5piM3JT9hjD0dVZQRPQCIcKcqC6I86WmLIysHG4ykww
PHw84F96KZONnkrNTvWqPxspSCXZi79p9+EG+glyea5vt0pMWAiL929pn/UKjLmDe7ptAJI4443P
YQgh3LG6tsO7YuEwGhvui7vM8BNJSUjbAyBxHADSxevD36rAeph96UluYotqAGaTe0+sa4k14YqN
DJSovyqmUUy7jpjVcS1toY71aReXSWv0LffiN05y4dqcieXl8eFEmOYKSz49foKHOlIwbn/khanE
8zri5Q8ujE/elaDo6FmjtaKDDoFI9UA1q98ukeNncHlEXOmdDs4NfeS99FYMBDE9MrfXNpfCfu7G
S/03Ck7l4e2vM9ucW2ht2XGnDNvL37Vrvi9Z2+j/bEFOTwI2IcGdpd4oxP0DDeLiYTlQ5ZfALneK
LnqXCEVYSn8+RhGNtrwO5xCJ4ANyX2gCy8F5k+FNcjXJaF+m+jnx2MpD2zjgF918x1d1GQYoZiD/
xGt2uKNV5sgCa7aCxDiykXMnnqVeZ1eWCJ3aPq8o7gaS2VcXec2szdgVWbnLRAZDx9QXcqDui7Cu
u4Lc6Vo3bYd/E1iTQ3mPbRlmpTpKBS05RWJ6u7E95c187RA7RLlpXXbCD63WAyPAW1rXu0VWFjw/
pDHK+jBfbazqLZPRcKMcyDO0vfERwZ8DxpLCG/9hPRbP7L8tdsfyg1+2zgu9Kwqe32psMh5cwSnu
e4ZplXnM2XzPdvhZfVvZi+MuKvgSkqkRNt/tssZFpwD/jtFbNakXWS0HavzYCqiDqYGeAN+VaR4q
s7uLAbIHc376/ulY47FqueKdHB6GjaBF9iCUw+KNJN3EaqhXE5mWlOJ/3x42SBfyxzrnhifHwuWk
lwcyTl9iYPEK0Dg+xxr/Q6odpVXTjpkAzyQLTMQ7h81UifutGR3NekomSHWC+iyT/Ljdvc6tYVAn
dEishLWxQlftrGi7CCM0HGOXozJ4TnhE1YB3l4SA2DggFkvOu6BguSAvBkozvjNy59l7l6eo5uVM
d5RTBJnISXsITTsVTz6FD6jJ1P8JtWveO0cou8zYxoWwEFWqpdYkU4ezajCyMyHC/IT5uZVZCnF8
uWMpjR8HOj2jSy/0T+geF+aUbguy6BIY4Rb7ewIAcNnF4YgXkS4V9szX1Rmkd1owZfKTty/1gULU
bR870XAD9avIMQHWzy6Sx03BZVR/bjRtUnfuvyx7iyfgFfJZmUWciDHTqZiVroQghV01oxy84/a5
DoqYkVz1QHHQGqciV7BoH2i2WfdshTYBe9xa3/BEldSVUKcbPRO1sOhWh78zBONTri7B2gfd98pA
AshTLlfn8aO40skAhEEwLiKVwDtBphLC2HKfpyRhPUKVFWgh1YkvwIgy/VCGfquk377Kmf82PXJJ
nwi1Gx/8lq1WB0MfNRfgB99A4d6wIpMGrcOM3LJbB5CrSfyZxQBqsqZzeB15vey7pqH5RrKR0ulV
Wln6LZB7GWN+p9y2IoFGL7TQH9jwN2j39cnv3dHZFYSdcDp0Xv1i6N2rSs4DvO3qfdN7R2OXAsci
HC2ugQIOREwrGQvhkRucWBBNB9JODu6n9AHqNHMTUsvkjpqVbr8tto6YRi8qwtRe14vrgFqELUWo
Rvt8KNMzk/hDeSSkIDKmFN1PFLGv6hHq7s/V3EFvluv4US6auoyuLNl0S0e5Hgcb3sKjPAvJ7Y65
532hg+S8k8oBGWpBRkS4gX47VlBTRToGVyJTw7b1z808lJHGP7+uQ1JYX20LBO0L3z24xw/r55ri
8WMGMiSWyDAqYSnMgrAWVSY0SKKAZWEBMYaMb1uyhCXi01+8Uyz5NSNA7vsoyHDIQciE3RtFwigO
M0K59cvv6lXm7r/veyrrqVBEwdn6Y+pUY+uH/8WadRxl/fyOhgk8IpLnZlQGzSVkUMqaFc0xBeVF
LfBMD8/MBfvKlajAmartB5beGHE6RFJnba/KfxcgFKiuCvu17Vgbm9FQwDwLlaumwBJqLKz9uz7e
ohiwzQSdltwY8Scu16GmJtdCIRNMX15gTygK60KtYA9XHOVPki0pWQLran3xgxMVMBGb3VNtUUWQ
MJA35rkqnJn8YkvaiSJHMYarPRlz97As31u75F6lJeyc3LikFiX9cxYw5dDO3qReiFIGncn0umI7
DtF9aRm6rNkN8vZizP0Slv/jmEi5eioceORE1prqqBe4YvQsAEHJo9ZT7uX7viwQTphFMejVVrs+
YjI4xzoRYRkJK3F8KcbTtOCEsIUL7Hd0IAH2+JP0A0LQFU6WYtn4bz1Fvjnws0x4zD9EGtW2S4Uw
L8/Cbh5d5iDbxP/tKbj2GF2V8XiZ2QEoMO1wjVIa5YlhOd8Cte7D9wqM3wNrurhVFJaMlmvrB9a2
MikLolxxkowRx6GkcMIPTjeUIX7oeBikM/HMQw+1H1pbCaL47ywQD5QWsvCii3RCxzjrOoHpL/OG
9rXozdf8YfUGUgigGCdnbwT+FzO0ym7QwaAbTcb+Z6LOHtoFT85ldi6SF/37TQ+/x+nBeB6K2Xav
A4Ew0f0OtzGsjTtlvHUPRvKqLjFLLqWMXhgY8gMzaHUsxjssJm4GrjQWgzWUSjRnMuOEaczPOA8l
HjZTsAOKmhcom5Gfkg2qUKBP/eR295VGDIJnJIUnzroHJCDX9y3huv2OmO4dtJvBQR4gnUto35Cw
GF4QsFcsSXl5oUbWN7ypcgoeiY8OnS4z1NedjBC1kojZtfq21cfV1AMy4SwDfrIyeq0zC2Re5hX6
kTvCHoXmh6UXCZnDKTzskZZbz1DHBxZbuXe1JDF4HoER1yppiZ2OjOOjeK7Tigc/F9UcJmFExcV7
yZfxzutSxM308w5m98RSiCwoc0XdpkW+zqxxfMmRMB3ViOzx0Jd4zKHVThTCsGb6MalImj4Tieyy
3yEl07MBBmGVU1vvWpjbGAOtaC/C3eVfPeKzWrGUw8vD+vFUZ5lVtacLo9B+AWFTSMhMQY3h6d0N
k9U4jRrv1wm2tp4koE6TTdYMs1ug/GOMUATOnMlo4pa+KAHdjmevkJyZZTuVJQLXcWLu6Zpk9fuR
Iu4vylWxl6Uo4PhEQ89gKVEBdPmxvoxWJEbG9J8i7CCQMSuwi3Cwcw9bR7c27JkBWlr8UM6Sp3Lf
pBUrRsO3IsST0PuMdNBP/bhZOEtgkTIWuvKTzEakRihOUPVk2VIC9kEVMbwkFNErRx3wgD6sMU0Y
cJUaDvI9y/QXbG4u/Dj+eNHj1DXNiarNV9TbFzluy1LOaXoQxgYJSfgG9Ebpah1p++3S7B/snVFU
W0LDEp1NJgTaJKjED1FBSIqf7yvMQciC+ZU9gAEdHYZD62/q1bzvQuPuLQq2CEg7GuVBOAQk+Vfv
6KLx6+MdVDwG3lHrXJsScmajXKM6H/rec/H4jJBG4EMb4VWDpa2XLeQGt6D+sdxhskzt3Oro1xJ+
MuehyVNbuCxP4SIrLDWP+rOzK1PtfnV0ypaQRmAYLlzj1pi9x2p5fv7ufrExGfQIoNtrAimWWDZ2
4R9je7d3lyXvssR5z9sjDXt98TozPlXtS+p4quOc1c1/JGa9BQXisn8XyMjoHLboXuTX48i5VtIl
7WTEnESXKIJ595q6/Cp0/GvUzTNJW2xlKhlMS2bXJKAcIRtw1NONKvsQcA9C+GJo5cf57n+afyzf
GYJEBuF69QpJI62/5anatMoHQoAAUo3T4Dr4ajNZ26FehVmfQI17DW6/HxfhL5aUxrh7+2EnwKIF
OUlvzmrQDlo0gk5iDenrhbVx0N+TUOZYyr94IL8s4BpEqPalxU3DTvwLqf/2pXoaSkbIxpgFiP86
+bj02kbhshBlA8EfN6LGhPuIAnPLxecOE7VY9oo1qyKMGzKan8Nh3hBkhFRwT0J1SNFCkVwdUOHt
pMVU4VwRvq8SxAtMOsOQuXhXP8l6kkHhCLjFrXzU4rzNKP37ZqykbCD0SkbLGZImrvaqyfxiBFM9
pa0d0kNc5r3/sfOgazycFDXaAQM+MrUzuCkhPZAFNBofi3xddLbTYItT9kTsrz706lDqgEVOjDWP
o8DjX9ycFoV07kRzW3KE2k1mByo94nxldvStzCZcYom3ChjrVvGXWfqzlw7NyZHlU7T5npmrN6YL
oFpWb9f9ydMRJXP4LXwn/4SPQdtABGn7uekjfwFqAvrVXcvghUn+MZXW0zjiz2jLNObxyXhAGZIj
B72oWWgFd3ThVl7IdUAnczeatNuPnNFXCtyyPw+JsfQn0q5t8GUEf7MVhbZPhHMrxNNVUxJJFrw+
8llS6dgUCaokxJndy+sd0KHNjZ5qKH9r9fq3C9erSZ9iWZDsSgACuJjZ/2TCkyiJ5ZmxI8sf7gyn
c5ksW4MMq0hX1mDwrARyVCkqdLs3absQ8hDzNvZLKSi/o2L/beIpSOJ7BJMQGTpGQKkF181TX3tg
B3RyP3PnXUIhOK6CrAx4zFOn2Cn1V55REYRMnMsDuEM0ZXsDQXTFeoaKFlMv5l2YgffeR25NxTmq
zQuwdZ7EqBsw2D14cI1DuENmbkjakVDq9VScSX6gu8S0r5rOvrnunRq7yXcHwSTRq7S1fGHGpIGq
o60lVEWP1xHTQSHq1X4SKVm8s/W/6grVPidjuIoZM/ynPYfJ+ZkkXgl3RX+LBFCjFfrIGwLHYzWE
8w1/uct118YYi8v2TJ1RvXK8eUkDiVQ1vpVpmpygijTxWILnoqztI0NeHAbdFn3WTZ0hhiiI3YUM
jkXiSrDH9OYrdUgRmcEWpn024O51Pw0T1vK/GVvA15uKRLFYaVS7jGW3Ae8dQff0/N4p2pFCiHqr
PC8RwQoRekeRZnl5Eyi0hul1KFddy2TXxa9jOH5js7BRysfzWdYP/ZSQHJ0yMIXV6NTdHyneeUl5
q/LXSPwPttdp/FYf7kNyJffWJCmAC9saLH3qL/fV9V7bErNnQxDBv8zuDe27gUMrj1F1U7VCLliF
3oaq+AGXpi9sGKqMBka48qu7pEQ4cc+ZC2lPELVQkYlCifk4UqRPHvfnHzUiUstxtR22QKbhsVqN
PsDYa2PbuzGt4xGSO/bwplVIqQ5o1HncgKYO/NKTb6c+Qo1/trEDaH4LK/pIDx7kXLFeQzUGAJNt
+Cerz5GsyMp1v0doJofv7GWS2Kr331ReqUdQWZpc6miGTpxXz6fOQr57oVW4Z44bknwr/gora80U
I2seTb91hC91pgUAJfL1+QjzqnAF7hadaODqwUmOg7EGn7q4/r2LKRTtjo/p3wHYoBf1KDvRqlUj
ZsONBFpuO+ODLAmKdfkZ3HItP+U4OU8IgLEiFCquFpV4auyFfeg2yhf6yYT6A/UA8wxyK+7LiVpQ
DKlShXG0RVjsRexgsm+YQAqOQFu+pessuUzrrz8VoKCsuKkRvyVqRXmZAo4700qosV3QH5l0m9KE
q6GUwFsK7r+txwsAEUBt823OJNrcHMyHp2xRsMZQflqDgkGuUyIA7vifqBdw6mHHnocrAjvSaOYT
4nvNR/gIQA9iXppbXYpz6WuYcxK8jmeuqBx8AwiZUUxYcw9DGjE9c7kj9V5VDjW7UVp5Q5EVSjLF
iYkrbimKSCIY2lLvBhaxK3fvnXs53QpCZuGEFmu8FYQ1OHwKsR2yPqtxJEq2udrteWMugW9jHDzs
mZyny+YW6CPtCNTDDV//wiVBfGz2Tc96UYpJU3eYe2N9WS3A5LXqUEefmzc+1kJqgCYBeO4lIuYf
W/cQ/1tu8FJTDNt1sbUCF2BwD4DY/V7434PcgaPz8fE6amfZJaRZioGmVDcRCt+efUM9RCt0c2mW
E/yR+NLd1R90bYJTsc2hLGRIng6NwdmaLek1LfH9E680DFlFvOKjadFn/EhBLCuPiMNKEO6b8U/N
sEuXOW2KwJvO2dACkzLJoKEfKovJuFWxWT6R493e+Ysw0NW32hYljVRoESdlqht3tbXXZJ1V25zb
i0GOofBUWNwIzc4Viz4aC+ly14H+b5aktEtxLMWLwEMvDqVUtZGA2JjwNTBTHGBO08dtXKmWtiMc
kFUHyh171O9JnIEITIrDWXi38Euk+M1xZBvLCLoNavQVbtEVGamwjtH8In8l2MKpjR2ZfcAVsIid
xzub4jiUxJzV5hFoz2MxsBIslUycI0SfKpBU6Mb44OBJmpHD87GlNV/fE5vheum7ambLs7eEyjz3
oZxzxdWcXLYCOUlhZWUlqGxfiZjvJPOkomE18/nStiWuXpVI9vByiNwrpd5gD5psEunE0IVQ6jHv
egyfYpsrwGaSkJwi9cIIRmG+6I32AvVLUxRCtgbzCLlt/2ZXch/Zgvd2bZgpBEwW6JfTWjOaeOJ6
qNLdE24hwoi4ELycv6wVcXMr/HYcbm/XdOhYE9TkjAwm5RW0m7+L5dvUdH430kPsNGNrCbKEovC4
qUrcmjciTp3ng6P0d9dLshqRqkRyuKogo7Pi+0utiTYo9pnxg1O8wBPS80pgj1vRwb3Up7plau0L
xu8uMsq1IFzmkoCsyHlXbhqQwARykvB8oljPUuPJypmF4AwdHJXnehee/xEaNMt9Elv5ddOq6WPP
E+qymnNXjBhIxLNtmzkGvuR5+2cK+dhjQyyS4u14g9MQxnn1jAlgCRY0s34tFxfqnM9Kpd7BWWx3
Bnp39m7xO4FUYhyYj0TGywAlL8PIJGCn2gw5AtML7kwL5oNM4EpI+mUuNBmAtPMYSOdzoLK4J9Zw
2AFJvs+jBX2orxYR/6NBtO8g7OGoa+uzxq/jFFsr4/HDFCgLM/fdGJQGflT4Enuhh8In3ObOIgpz
FCRimXOFDK4LO2I15UEV3MA7mVTI2O3WnnazkhN8Q4PC/Umxp0tGgHH6t2Sjuw5XfYBQhZ0INAee
aI69im9Ocdvwc08GZZ8B4PpNgRX/x0l+plMHuMdvHH3aCOutxcbBno95zG3C34UJmk8IsPDkEIqI
OcD02ivdpWlwOzfiKow66poer2wmPZOtzXgd3DxO72P+AXHz2UxOWCz81pQSLvnng6fnhUlAstOR
5UTlcfgWSsU0u75ynHdWqsgV4e/MSRRWuQhgQ2LMgPenEAMmAHp1Jr1M3ICcdE1wx6ZZtVmAb6Qe
kV8YqYEx8/T5QuF56VDZhvwuzVTgJt1H4XTqN3NJwail0nB9WACrRUsDjH/L9X9KKDD2UjV2t3Je
R0SX+Xe7pLsDFAlA5tJKrJb8h7qbuj+uHZIA7fMB8rBovtXl3cDT0SnqQBbPYxVPnWrDN4L2QFgO
4k2Ho8nozg2iH9hHhjW/yIy+gxuAk3+qgSNN7XaLM7DUzMsgLPWN1OIj91O9VEgA4mnX4YbZDkd6
JUHuu0d+rg/BnKXiIr3dKkzBVq+b5Hx0gbYvBJBfOam5UCurNO09Fai3UsgZrpYCTZN+Y8o07YAO
HlYZq1Nw9STZ0g8GOW7F5akQ/c40zxEY/XBF0MavJMiaoMYEkkuKuztW9ubLM4FXZXDqMcwsDq4I
t2O18qSNWDISZNFZObBpld8n3BosjHQQ/G5W8gjNClho6OeLYbQeuv/BiMR0+pC0HUFsmeOBL0TO
orNPbooSDgEoOh4PdD+LKIBNu0G0hCk5th8ytk8kwV5bu3ioJzdcW3IuPL2ZOeggQTrdK8Q00xGk
G94wv9t+Ehepcg5MeVs7FJDgLu4o5QgYh0Gvxtc1b3oXCZz+R6PZaQBYTv0a4VHhSzmubg/gw1Wj
jLxLKXxfrvbLtvPXHF2dfSzdgQ+b1pQ8XXvFJ68xNg+PIyi913J1kwm4Z8CiyUKtPM3ac3nErAHl
3jn/Ja+Tpbnu69t6+s4crL4ZvV2Hx65yPnmUHPdot8unGCXUbTP7QDPSQC0MWL7rgn6WQpmd2PRm
Edi2vgyt17WgDahX0JzY0sNIxQuvkIpsSFir8cxT9sgdLeWguoglOAc+TaMUqMKKrig0YoVebcyQ
jaq8K7VR87I+v5Rbzv75e0nJzi8keniDC2VtEPa/reDxaaj6gOC2M60y70svD7SNtfHL2KkSs7Bk
kdAZiPbmyJ+NmXWHmad/HUtQnDFVTGB+TOOCDYgHEkEorFPz6C9rudQcqi/HumJ00F+r2zCH8+8x
lVVMSDo2I1O0Y3qFAZtSo9F5s7VbvzQcMrccq47/7PIUFDAgYUE+KgZ8NEH0KIfwNk3jGd5uAx7M
E0t119y+2Yh5ZwoF+ZjsLMXUduJoai2f7Gts+u4XuOr2p/6cxMWhWR8+goMDcSIoD/oqHlmpeVnz
DaOeb/mTCR8AnWeE8NmbBe+x1F9fIYdWlj8hid/wc6lxQeows8bgGkgHHpUlDdjcTy/1XXoo44/s
+4n0nwg3dbcI6DsokKDc2KsSVodB6MobOHI1eZBfgaJLCeIBETi2V12ySrFwnNIXNXfC16mycB7i
F+RiquL6Sy3XvL80y05MjV6Og6Zf8iOrT3SDy2Wq+s9WDVywD+Q2eMzwL1ngvyXrmVQyQWhqUVQz
UJJhWQJHWat9xN/oOsSfY4y9eqAyNDNgYAcsiGyn1M1Yi2LfQpeDxSnaglYnBdLgzfubFN4FnJBe
wHdGCRnP+MZ5s8zuS3SAwpzVov3SILJ+xVcQapj4og+59/+DiJK9suNPA46shZ4C8eheZuScB4pI
rQc6MDQGo0PNsiD7I9MzLntXADRUPDxoRzOC3c/OvlKomohLQRd/KxENdrBGnlBNv38knFkJIZ/V
5B6RU85vs3131pnjElVMcS33Ozp6McAVCRleC6r7IoveH64bF0M4wsCAUvgE9BOuPN98mZkD3VaS
4obD8U5URGShp66JeffCAoAgPIS2AOpG9b02gVwbH5EfbgwpcXgE0V2jXvkNFuKbbFTonGkP6We/
qQy5/mhrC1ls3izw9XbqKYAShiub9CntsTI6MKDQIkbEV9BOCdOjJIIUdDo52yCAXyReT7BTrkkC
34bc22c99eQOo94YOVN53EqPYYPfyAmFl+14+9ov3v4/f3Xr7XywRIpTyNGOvUlrfc2Kxcy0m5xp
EIS3fYU5XNVYRf4Nl1C4c/w7Qk9AwSeMnOdkH88LjgDw5VLnOyszLpy3cKol0XCWrPmGjaHUwNdN
1YzaRsMcpiY8Bg0K4j5KdM0XL6C/1BK1Utpif41XwZjMVj2QW2e7I16omej4LeyPy58SLpOqcSq+
ZM1vFWJrpnshCFruLigxFottMjSmr6jG+a7YdWg0vzxF3XnNCnauk0JdxE0DIB7aUHeIWeeyejRs
PA457dnQ49J0MY/eeX2Nsv4wQaYRi6+oiongGH44F5cf6lJJqbhXPMWKdaM37zLODcPa7p1/fNpu
Xq0R5VxcGsjsUut3Troqf4LI05LVdmFxjWHrhuYnOfVvbS97u+5TIUhuY3qCaxxIdPemQbM7FDSU
UAiPY7649EJiI+Z0/Nc1pLaQVJ5u9BY2BNp611vr79SIAoPPouG8NkFb7TFY/ipd0d0vv8j56VVu
AwhwSMe8aIxf3mbCCOeDNi2ogAim2LA0A+dEOj5ibC3jJ5boOCJGkmtLnT+6aZeL00/8SWS+odn+
i2rosoQxFNndunOQb+2a/HhswZ71ZCi5Xvu6lH0BbmST2EW0hVjUlw1QmO+eBErqhWH8bqtu2Y1J
VioRwqC1Mm4aQxIc7zB8K1yTlYjjdaueAW2kYt2HHKeMSdo3KKrioHVN6MLaHBbJlFEOVGV9Zlm+
Y24VRf/efaQZdkiMuwnOqk21c8JXleF2gJrB2ezUOt6xMXC1gr35Nx4TMfl/3+eRVqppajhnuq9R
16lFhVwlFGMMWX7XkEN7zKbhamCmX0oZM59dHvFq8lXfYHiAp6213RaqoNFlJ8zBLyBa6ERSDhnK
NN/ZNVxXHW7YK4UljSWD9ruVxRlHZOlxtlHaCN9VUB7B1MoAaDhMr7y7ecJ8i/7dbhC98qu4KfAM
VgMcm8LOh3abtcFQcSDX9YIxLhRwoKw0jbrtAR2HPoOsWOXvjHY9vVEEkT2DppXAkU1EGqt2WCMn
LyIuxfWrdFvQz58H2vlkoLGYUpq4VdlPIliEiWwfl464Nib89E6IGwB6XM2++pW3Vk5CZ5phVDUH
Su6D+nCzRXn4nvEb6ughZyTWipfISC6MYRPgAxMzGjkaOqslFEqDdVoh6NegP7umRLp+B/dNRCN/
xquDvFMzNU+/uRbmdYd15ZKtPfAmh5vn9x2jX2srip1qXjgptwjY+L1WZQHwX2FX/3DWHo9l92/q
CkLxKfmoY2CkapmhA7oFxI1VZHZwtuNZ38PR4G8nWeJtsb2Bct7u+FB1/XBlQ/4jzRKyGgu5pg4b
jxi9o4QfVS1iIrzv+3L6ooi8p9U/tHbqtoMcElhakRWWhpuyXVa+Y/10XliKKnD6l5RXjrF7K69v
aL15PvjJ2Vf3Zkw2Kw5ZFb8KYNoEbQyRNVyq+CfmInJC6BLd78drVFbHL9Zm7t53WeB+w+vydimb
KuWTSVOuyXWyU6GsxRfSzAYY3maZBWskjuoss3cLlgqpGs5K88zTj0K0d+TUPnA0RyPQv+48aF/e
9qdQCyU/ZIlstPAwdWPAfDxYYVDT+lcQxFrO/OZPk0sn7NjARrbrSiNLWVPxCmT3D6Kt4y2/mvdN
KPTPywukoB+Fdof0daduLJfQtzsDgBWk9eCkuglZu+XalcRbAaR98j6AJCN/W6PGB0Rut3L3mBMJ
xOKSzyhHLd/LrDF0IPZkV9o0QDkCpCrnPMN8sg009VBzkwleiJ69mjty8eYM46ueREF8IbfI8BJ4
WHIC1NGw3p/5KliIP8CIjLqNDAb1jFwnKaVEuzh0310BHjPqL7PqOoMmvwZ64lvanZ4T1RMKf6KI
2KqYpXar1sUXcI2qnZ8T2Ybjrf83iEpj20+KVd+sxq1VoAQA1HFFtUVTTSQBOhFg/+Pn/nKmFD0j
KFoRpQ6UC7xUBv6k10lSsV5OG2w2u7g2ItoSffgmBNSX2kLladF6+D918U7MtL9bN7LpXywK1gL7
qGTRcE754juwXAoOxSNAE8UAGg47YOHIDr9vMKW7TH/blIb4DqMpMNzNLtuhq/+0i0s7gMkinew5
ba9+ytCig6G2Jkhaj6ruFCbaVFKdf51Qpif1uYn6nhmzdioLThMNm1GgyGdteQ9ZtrTxAAimaPrv
BQiQspwC3bvbLIYGIWy0ToJeYCKgptRhnFqh5pMeW8SSBxTu+d8BxnZ6UyVcLSLfDl6MVFMaKZAM
yR1tZuqYTdkLc5S74PRXj6RuQrrFz2LVuFwByjE7GP7lyELatAVr4VBw8MWjWbq/8Rw1/1GA61OM
bj/QUlbOUJ30bUWVQ/9nuO6pp/lbTkM0dd5J2EUag7mfcIXdOY+G6Lyk+77V26ObLxFGgmEIV7cz
cdAK/dUPZNzMOvCEcI9dP1qE9EWXrpT0tpvzM4wcPwpxyhYuiaTJUt+gTv2JuHEYqV5TN93N5R8O
InOfcEj3+DA97VN4O1OkxDF1H47+RWYKPNxWgHxoneOnY0hPS2lyJNUWfkK3J1sl7xiALwJB4UMr
IQgcr9XPQnm5MzxL6ln+NIm/W8jxVJLgVENZ5FmawCQZC2pCB3+laCgzg2wy+br7O/R5uvg1RlKw
ePertPCROACKUmhALuh2gY/5GCQw4duB+jcz0/O+0QcBcCjcqmlCnIp6zh3l5OTKDtAB+Q6ijCET
HtC5gUHxeYlPIMG86fQrj41kE8OEX61DoJjOk+kYep5L9Pc/bJD0+QDuuZNU2NlhDRs2DIixKGhv
RnX6g4hlRXOVr4FWjh4KobcgGC51/VX4kFQakErADZoKHJD0BJXmx2LHzylgeS8PzxFB07zIej1i
qycv59joF1UDsAjsfkxa/xKYWETwDA1zFqnyTMhR/1X3Ziy4x6eZMBkyjrDz6QvGeNuzjYgL4IP8
JQg5fxkcm0MAAZtfFY2U8tvnxBcadVJq04ODc9yzbvgTxShspTgazg+gma9w+1OE+1+ipfO4FJly
ScRj6pvWfzy8TgzkZbg3JAM2izErqsZZUVrW2gFDhH/akCPRteUm/lAgQC3VhqWqfOC3y4Tou5BC
4rQwinoe/agpfw/2jywgPNR/GMlwsIM0+ywOE1OO8nasBOrnlt9LkCE5+ivDuNVvLsAFsW5sHpL/
dJBoov09FKYJ2I+H9XgePTJW75wgKfO5O6Syxp1JSptF5d2ns0tMHxrqd7hXzWUxYrIcV2bHhx/7
PG4zfOnufRE2HoVF7wW1c0XSgM/7pZrPCLWs3NwT2neJ5/MzJTJvhurOZz62fvpq96rr6fbXoCoY
XCs83iD38FvSmAl6V4O8FblI1TpD05BtsK9Rv7iXrgNJKMAsAwS5Az1aYwBcSFc4WNCLjlpou5GF
ufPzwngEKtbCb1zMV5+J2i/jcpnTayn7B3kmOZxgHNyIdbR+/zLJ61kIH7SNUsukDjX7WypGTOqE
zwRraAYWq0+YafY0nOUewvGAN32qZXtQRtmG0GcCP6L7SbHRG1qkRJUxwb1upA5qxeGo45thoz74
G+esq3cyX9mjNzKVfX9XsLLnva/fVpuOMp2u3+23iy9svm8Qecr51fLSc4XXkIyORhXEczvufHIG
VF4sH3TAY9jnt+n2DpFXb1drdwFsn6j8VNR/gWZPwvAf8SxS1EZsYFQHJ+wke0JQ2l9GZvuD6PqV
opbeJxYdMM1Y+OsUt3Nl5jv/+Zu+6V4kPRdePuLbm127Z5xmaJA3gts6zUMIau35I3ypfwQzHMpk
K1gNZXihrZlj6UYWIUfRd/r+MSGSNNhjMG7TOpSjKQw5D7QKm2q7L9SmaWvw4tK0Mb6sbA1Z/uee
DTkyvOnMnP9NpCMUMcb1nFIA0onJM239yfzBxPXjCQ7gbg7wa2BmlEcJ4nke7BcpKHzVKNB6hkxJ
OmT4ZaSluk4Q3G5L13uvblA+vQd2TDw4ZYY/4ZLGV5MjKMNV0EVLQOcIIX+TuLwGin//EyM/gkig
mx5fRq6NV2rE9zZxBY+Xti/GgvYBJSUS6RCfMBrdtmA7dHmFbw3VzXiMkqTiqqBaN+QQNezskBHw
LQtPIg2eD8Z4whfMPOP3wU1G2r9bLhno4DnMSAKx6obk7juot5Qsz5V3KT/lKYzNCz66d3CyIHOt
QqqEZ2uOXkfZ2hCKhLexsElwLVI29hyT5eWnJL5pTpNvCGqh43CCMIn9iyCTToqapLJbhN5eEVtD
taMXXvwLoNHdszxi8FMavvmE06BpwTaOdgR2ug5tk9PF4fXlRWdzQo3FCAhKWQET2KejmAD8OJOD
a2NMJuSklLNlF0YQEdBMmZ/jHnKTrABKPr+pXnuFcoTz9CgkpGEXb7i/CdLiJ65uV0wvw3orH9Rz
k7IAxnTCEgw76hH8MWF03/Un7mhWyj21TYYdpEEpb8ec1xBmgY73mIfXMygUMNwZS0JxP5tG9ulZ
kw6d7DJgKRgpVwjQIZiPWjQuZFKvW4TTNoSssyr0fGl0tuaxlDhrElNEfVEjI+7zIjHCzwanDpPr
M0haOwBZwl4po7styLx99ymwH626e4k9D+izao6cVf+cN+kcCf9xObJAQVYM8Hpg6hvwbdWufzKs
grYG+s03QE83sDclIu0QYif7MJ+BmXItVYeYA44Us8OWNyg+9wIH9O/5z1yQO4yvmJ18Vx7nurO7
FUPWS4WpgnxOpWtnrW8QfznlfvlNffF9rsczUL1kcIWAhTCB8x7RskmNhon1O3/zHDjwn1nHt3h7
6GZV0EIinK/hvmlsoOMG3uky/k82Brj3mI/yGO/TPoF2gzleYKamn2VuoneRLP9LoRFLNzeMxmCr
Ws3jNFfMqQRCMS8fMgq6gBY/VKzcBj2JJOueXDLFlIcmuKBofmn+4DDt7XvN9kZYhAIy+AixqQD6
4RjKpP5RxTFMZABXmN52WnSvgRRfEl7Xn4XWl4cPm0DuQD4fwhhKc46ezgbcirZxuOSh3DgeWegF
dIZKE+YdvpzMq79r2NAoGTfK1gLrLsUeGth0pqtq2NKSjok0XC6mJy2wSn4kHFMzyJo0YWHWjAd9
5n7QZN2DrMTxgHEMpUUi+GDfuN3DjhNKbSBbgPgomrUw66AkMy6z/VfJdmbUtbokoa8PU64XJSpW
06umXnKZwKIj2cwxr950tpLPJZYdKzsE52mgXO2yKijW/FHPwctKyG60QrK15RQiFnS0R5NOj5B+
yiL5e2ZXCCfdvJnGv7wIZpBzbPdVNn6XOkErXxSNdimVnh4wbebwwYoWfW72HbbI3bKGbU53jnKn
h0DC3hUSYQMTl2EuowI0c8uywZzzPXeJS4wOV4CrA2TozE/rrSSALC9Ymu9nqcU7eDQ2WeAYtW2e
Y1kQjYGKv0e6mEqaIe6Lc0IDkbSm6ePNnj1tL8X5ZWmmHwaIFSPxNM6tYCIiRvT9WYjxOT3W2ZEU
ToxkNFIQpZx7UkSFJdNZwtCirjO2Nwkd9IlhAJgNjWFsaUf6reZ61qEUZ+EVVbTSle9J3XaFlHWK
XEOFCvs8/3CnMerdm7Qv8Lgd2WD8VFHULeUyc2IPUzRgE9UJcMVz/UVjWjlw63UkJx1hkqOKhomp
0aqshoSRSbe/J77eqeDp/ulQn+a/FHF8Z6ACevcfaXtRmEAeOxDQRdj7oGXjrDs5CkB8P5ux37Bm
DsRb4HqeFqWwm68fytbplw/a7/4jwj4kbAKnbPYz7m2cvO3TWKOF8ZXE92sao7otKqOVszFxKx7N
bw88EijHIWPdPbeLQ2UM6SDmCdfQ7L9+mLF99cJ4Bmn3qMmF82x4A3hvD+KXrNl5SOjXVygYsFfL
4AWLTd4uJ+WL7nkaJ1lg9g94CiqsLCWu3fdvBYSmsS4T4VLhTOGf7J45v7y+2EjrmxmbOdXkiFHp
8npCQK1lbRuUR3Ee1kpCwr04vosFbUBMRX9by9JpgEVv1FkyxSGtiEf+RqkuMDTmKuRUsEkU4SUN
0zk3eBB2QDlKUm/0+rtRJns7+u3fncgQnHodrY6Se87AJpWNH8NLH/p3VahGpE3TgRZl7bXOGvj3
qeTWlWktP0rYpVkCTnh7qc/Ink9G8VMlPECD2rNxAg5QJXO/D+CzQMQkHRPuzxhebIPGr4g/amiY
qrKrAB5N1kJbDp/TxJQU0HwGA/XwPASZc5z2DQ9AhHud99NzlzFx7joQc+cxCGFvAHmyHtK981l1
CdTFSokJFFxSNLTbWufMMo5qqjX0wvNM1dl8JL5U76dExuxBwJnks9JqCqPrn+Ngrgvm93RRWgQt
ZVbnqYzXXDX0AGREH1zdTzjYDKdywhJC1EgQTxTKaGvoNHIyIPw8pC1+X9ef7GOlhvIzcEYeZZwr
SfKat3nuDcL7RL4YPUZdvi73xEw7ZRmHlkztyZuhPNMfkXm3Sjlz8vv27uS53xS65WpbXmdwC7kg
xMhjymYMl5XfBKkv9LV5dDwIQ/KAojEd7/abA32HJbxgKWTxhhvplfRVVvGB4+lw7dFFQnJPAASQ
DgNJmePsfMThAkXCD2GG9uNOyV+jjBMJ+6E4bF/cz5oIbOxgy9f+L9PgDBs9UI04DEpcnuPkQl2q
NFTnnU0KOoKDoEnLN3jsFhv+vO8VmD0plzJSJh0OjKS6gLslbV0q7EcsHLtSyBdB5p6+3jOtvUa4
5l2xQiIIOc5Z236jp7TLoBTBRlCIO/r99J7CDJQjuop0k20YYz4PS8ULmxiCtWOechkZ8pgVglm0
RhUYj6Zg0EKacT2kdn/jWWlQUQXckhBoaIeSMSSFfTM5u93bR5/hZu/8gLr1LtMqs0J6LyX+D/xH
sQfi9nSjJom97kHD+PUmotXb63g/mpe7xFhovQAZRRQLpLUncT7m5L5cqZuMXd5kAKj+Bt2TexIZ
LMi2kcyL8+NOP956Q9HSAQqcLpJundkyl7Phdv0m3/n1JhXj/nXYb7I1teXpx7tPyKXdf5SCmR5M
0cTS5fAEnF7vOmNyXLu1ZJW61maRJfzCqmvFRRwf+Au0Nhp9G8gFbeUL6iskM20c9PV5lOuQb1VQ
TwqaXETfZrDFdAZzXm9wweW7Upmue7Ty52h/Plwo7qsk+lJQfjFiU66oO73KLXRAAjtvDjBCPA4q
UnSLwHXSLIvD5OxpOi1dcy5az+I7+RFmZEHviix1/DLEVMOKBh/XK6QfH7AU8m2R6K8gLs4z+t3d
Utsh02t6shsBFTTcfyDhbRm+DfMU48F22M90JM1+172zisKtKjAMVOeSn94woD/gLFAU8ACKnMXC
F8OaJz62dQL/WCGvZkDoR4V1ymPgt7nEedaJeblCLlmbWBXBan77gmVid1OuUNW3V/uX6XlPGl2k
2xXZ67HQ/+4PeUxloc+iAdik899J1A0ayd9pd0+FeP2UaO4WcQP5FtqYbwCgCp80/5W3MCO+aTPU
e7dNGQw6sLRHNwd+S1foddqL5y3NiUsRc1JKKL7uKp824RTuyUUkflNiRsX2181vKB9s8c0ZBpxI
Agbzr2Sfnmt1U5q4sjdNtY/lKuWqQ9piLxV3+gICF1TiUOImpuINcIr4Y/d+aOprvBcV1Y/vZmfD
oRI4wqJYOKLNz6ag1qdGzQym3UP2vcxNgJQg3ijKmQ9vABU00I4CapGyx2385yNhLA+7hAVP+VAW
BN36qcUkxSeeY5ClA/af/vcXbwY2TP2ERsghvh7qPbNImSLGUz0JEnQFv15gWHWVux32raLFy6dK
e4eu3CcLOx3shx+udwdZVaebntotZUlCcRnMD5Ms8U/TqIajR69x+8Rp6WkRis2xiwvDowVy5WJN
zgIpe0dUrUIaOSGLhdlWxUH6kjE2LQgQ48e4hEfRCEhXoI9hEUOwG2ry6K89CabvALbt521yjsVx
Fek0UBNTseSPgHaG67c/EMFzR8VOc7IgYEHTqicSUokeXpIuktE4fwivnunPoC9jE/++8jkQNLxl
h+MAaWtWeidNmNk7QhRGDqmCGkBsxXV84XLyfHzv2YXsT3d1861Qjnjsg2grW/cT7xYJ/LF7uMc4
/QZoRQzMQRW1nHwOgSOVosv5HaGeTY0SQ4SlxeRzoOYpWPObEp/+5LnahBRCA8AF28GaIkpzvrJ8
xzxhvikRzLmT7ymDstRYxRRzsaK+SnJb9TT8Hqy4ffckgzRZ22hHfiUAXjaPHC3dZBafXaON3QCw
Y+dkGXhmW8g93KV+2kxW3PJBnn/BPQ5VgClcSbAarS+g3RHyX/Bd9ZtPkczqVgYsfxAcs+i9Hm6+
xr5xgv3jvJvlaN41Le1fMYfV0EvKEG/ZUhGYEQonBeeMtCB9auXqydRXAkCfaBWLOSNcjv9BmLat
rpQzRGwRtF9VGmY1MVIfFDIWGk++7229XockCzf1cKmITnQdhCGaj1TQTEKY6FuqC4GrSaAkdfx1
rcsuD+BS4Vzf87jHRnbRiOOxLFDBR22TChDU9Bo37hsNdUdFQRdckQqCLykT6AhLZOZgCXw4a5eP
n9Y98RO20PAwOveeTM34Zc5cUIjmeHR96L/TmkCl2l4zJG9gfq/Pi5IEyKettpZAK5R5xosJb1We
YtdGachDVucBlb8tsL+L3JXbspKK+V+mae/9ljq7JNQT5TjfwweGcAO/EnLsrMYiqfOq7A2XbnvB
9wRqvUpAbzvqyR0gVeFmQPiJPP4BiY8CAAF4WJ93oHgAk+zY3Brmgp7oO25D5keXpQ0rw0at6XQ0
PYnoIAfEocV0uE0V99lz42wdhaQvKBcxkCowys3e5c50DRuC3j0mhVcSzXAzJv9/N9BmVNGarz2k
rmkS2mWtfQpUBOrdRiBT2/lHR3qA9VcFwzSFGBMYKZbNhBIaF0rnUi63n6mtPczuT8/3U1mfcuF/
Z1hUtW4I11JcgowItXC087CDV478ffxnZDfwVZzDAW1Rd8MV6zdiER2eS8OlEVkmSsQpiTFGr9Tz
4UdPsLe7KMo/s6kXT1j9zbRO7DbPYPYSnRGQckggu1Qmdfbvi6/7GUBEWSZ+vfiayPlWn3/eFe+Y
QJxZPD6KrX/9vE+V5rP7CA/6COHLjLOGab1VF3hjDkE5DM38L3tAPX5yoJJwYkysFcmun9UcKSic
/WY0IVvoLq8Hd+o/GUbuE64Ebx3Q5d90DarO9hStgAHFUWfA1bFM1Xi6rCAqFBNrlnuBIsmEBhNX
dUrC0scmqrHP5w+vJGgY2jzP2yemEZjqI+uKpomfoBIkeSq0kiSre+r9GawI2c+uvkrLrEQTQ1U1
wWdYR8si8VsdwDpHLYvmjNf4Pet6QyAkXUafB/2QwbSlglcqvztK1pdSHpPayUtWrMuao9i551f0
Ypdoqi7XfH5BlxGfb3d6Aq4DF3WlJPqwgYsPqZrQfgZ/DLSQFlkw4SZMqk9+caQDrlbKUH2FLNFn
SIYHX93ijMYPo7g1PgZWdc4suk/4Xmvuhs3kHvG5T4WGxbgIfROasRb2Z5zRGVsNB+ZwfVZzPHkP
IxESbG9tuqlMelvVui5X0J2PAlXU8oKyhjFvaIOr0pq+xau0r++H/gXiE6+v4Cbgp/k93vYSx6BK
gKOQKNHFZcLMUFiu2hRRr4pQsBOIXVqKa00nSStYknnI5jbdaTCpBozLNUy+80l+Fsa1RP8+3+/o
im9zOnz414NiNjA1IzOXBSzWjxsYhEC7Op7sdXZc3GnFrx1Zkna87ReOwJXlMiio3mZHkcCRJDv7
6VD2YhbzcLkNvU1k5b5PLwwlRvO6G6D7AkaG8DRYH5Rgq4R68oDFuk1D5gfs/6UrK8+Dmh0q8sdP
Em23vzBaaxnJjHX3syO0HSaoptQRViwtOypNFzrX7NyvDcZkAOTfOgOULnH5RX/qeMIledFO+9mr
2x2yfbYNZ1y2j5ZIZeJBhig2SUU44d07L/D2TToE3h9HH0MYoVXXTjhg0WwTvrx1QuN/jPnxShj7
zM6ia7Sp0Nq6TMgK7QjTPVoN/W1UPZZcr3XEgLTiew+0BWUqiVmeg86HpqcgPIr4FnKw7hIWTnG1
E0/l7TNsjFpQbk79SYuPNVVsXv2KIgvjedMZ9MulgDUb407fpvjVRZ6/EEeIzfe9FS/+6QhwXPcZ
AgvwnBQzz5vnZUMVvQU9E8RP3Jxw8+eFRD017gQBVqw0gajh/W8My4wabWC7P8LDJelBJFrMwS50
4OtNCuzpkiOFmSzaZd4UGdakNs0qIyVzDJi6+kyiPr/5l3hJpxDmBP0A37Qtvn98899vOb4OlwhX
fpWH6tvTIC9g5mgy/Hz3hvpRbmInkyaV9xYEiMIFrGsoCEwYNygip6dqhiiNdwlOv4jW0I1Lcb8Y
3O8+CPGpbhgDCMrwv+V7FAX1eLWo96GoZZdgJy6LVrEqcfUlSMW6GmfRRGOdUF8ZJR6/UBca8ZxJ
XHq//jTeeDDMkKqhJe8wckRSebDfz41d4kYHIBrEl0tl9BKV8r5go1B6NuO0HOITdH3RvWE2+mDl
NblKAVxXRfyPIsRu64lgLmVbOomObGW/HajUcCzqGzGhVqsS39L45lLbcD549j8un6BrwmyiO+Bc
CAPVyv7+Ooef+xyaZ8m5wF0t3KE1XQlGsn3Buu0VMeqY/39ub8P6mWee1/qS7JtITfjUC2/jtzez
R9p6s+NLUze2iuGdzJHrGuX+UCi0Vfc7HhT+NFcvDbtbsVLA1Z26SyYmf4p5u8dylLiZZTP89J9e
YsCfjKlw1FnNR9CUSO5LEIXBbQWocGnCY4s6JB8b6RJK7oTHqTZqfenNtgTBwfWCySZ24dSMtWkE
7m4U/kJgl8hJTCGyii9snpETLWkUIHtwGKtRxQKGumHXzQGPMlbQMo4VtVj7koteuUieOnztzoB8
qgTLWhJsJl4aRLJVOGLud8QV0tsaB/S6NBGCboDfQ73Xw07027c6bneyOK6S+Gsk88RMpGr6bkS6
AOkbKpdPQRrr0hfDPJJ2G/t25PHn1ly8LhgVPY6HiJL34Ff6gm5inTagxwP+hakEoc0bCeiCqTFe
4x+DGXxIDlL7XA575JVyhL/HfYcIubgetmotBcTPQlImDpP3qzvlqkGw1A6tEr3lpGa1XKbKdqeX
JubVzeewwgu5YFAbYXkIp1CfLkwIHZwEZTCwgTkKfQzzcDaa4i0+PhmQIPPDiJkZFTEi4GnAuh6c
REru2s8ko2ZH4TOqQkz8RJxUwKVwoyRj/iUDul48lSTv0Rcbtrcn7t51o2bF77fQS3zONTsRdiZ0
Io+EDuij/JIxW4MfSJo+RJ+sSyPSUtMVRZmFCtBBRbEyOeA+8+y4hlEIpun+pHtx2O9MSPsJsGHQ
4JRfljWbFiJKJR87oxdYO1ra1FdChVlqjnBoYU95LjhOoF2c2M0M+bXHXrHAiLpHlmCfh5rasGSQ
Wm8q1hjEUUyJ+PSsMo01OG09c5/2pu2HCK0UcCo5HiVU2UR6zvuXnQXIuO9P68JRI1dIMOBWEaXs
+G/3TcUZogwFstmJwa1FHPAAGUUUkbjAGLVccJp8iQ7CJjMsgTZgXHezWA+zWrZVzl+2L7xTIMYz
llNCRUfTvjQfUKgAcaz30rkwrVXYphT7VQPaNr3Pk2wcM3/wClsoBigC+qUsCzCq0SwFtwB5YQvs
njVMlX2FpppF951mQzq1gzjcLNYgVGL4Qs0Cj3UAynAc2g3OGUrE8j7E81/Vhncc3uGEG1leBVMa
SYJ1i9USkdFuDPyOkXo9mlTxUFAXqdbhysP0ifhK6u/DCroyCMrdfgoL1cYO7uqeFQ2GKYqk8gD8
d2pat7JITIflOjLii6xrJgJ5tveNIx8TyGtitQ3T1nfvQVhinmJNMK8IY3CxguEMAed7PPlTP1si
lq/ACPs6+G4TYTbZ1zboMGa0rZqwQ040pIGBPGIJvA99j9f9T7S9Y8Iov2dc7bW2vN3jxv4S8s1U
pJ7QzmniyO4opcrNrfEJrTwQ77xDw4wGcSy90naxlBDKEcSXMEKuhOLC4QI/r+ypDSvxQz8dnJHc
JG2VogvIzDJFVnZQIUrLB+sqJaaFzuqeJOUlR7/JQeaDYurkayA9unoRrfqsaWdsVHM8pgKYxZzP
R3FkSIJXHLJJE1G2g3IxcPQBvFPlS+o5y5sV8M4ueusnsb/K940wyRFnDYDL0Beu8vOe7/++UDR1
jXgCHBjyFzpYOyUYKz/pZVQgSXYHCWiCPwgzhOHR4/L3zY2xJkOcOdbAagbvwKmaD0ncE9KBXetz
qkcowsqb21O1qPPmi+ps/y8f7ksID4ddOoVIsPdoBCTb+1ENmo7BvxsXlwxZWiVYzTzhAu+mvuA9
ABHOYOYp8oFcMBtc9JsqbJiakQ132+0Opd6pMRd3FFJ+vjQ4HXmVBzg4Rymt7arhdC6l9nZUd39G
28z7I+Lylg3eFXNPFs7k2N0xWp21VnhKi8c/SsGzSRldmZZJfk0reef1lZ5Bu3ilO+mlLeE6/0c6
nQebk7pB51WdSWUsz9orwwdH0Xu6gw8qvy91BkaGKalIzND2WnZwl6ywvxkAA5drZDdSk9qjpmwZ
r4g9fR8QbNYlET8nR8FwKvoWSf6lCLiC62jSQk+CcEwjnOS8LRiXz3r/ZiBdxBBbt27Fz09l4pYh
gM9iXIUymVFwph7PG2qh1x0bZAlPdBJWHZvMEd6Q5I7tbEtzZgOH9gx5NV7zqyixJ5Q+ahYBrt85
GlnamuY32m5+Co9yrSUqbnIo4FQmMJi0CAZccAyDW5sDiEQaNOo/hmCStOBJRcHfflZBUQe84O+T
CoXSbrlpHXArnVfUz4OOeFioBmq9Qmyqsa1cyADD5Bks0mOoFMdv+NZSkVv9iiSe4myE6ofP2T02
7AAs7t2YeVtD8HWDaYi7gfxIwCEM6chvKbI84QJLzgAzdprj4CBigZjmzjzGxVAFFEPQtjPPz1B0
Je4unZzA/ZjzH2RIYOGrCtm67RLoJCxKOqNs+6OgtVno05A2cRecj1Z+5vELMeajueh2EbchkOoi
Phm6OjKdy6cVBmnB6o6c7iE92SA8qcJYpBBtYGlw3zJeuuD4nbUkq7hJgnT411kwUaEXb0XT845u
VKI2McV0yupWq8jlryj7T45yN6z6N4saQd7Ewb2kNHBn7RHZSJQVcTn7T9KM7BdFBkPVc732h3kW
maLuBIh4lR0SgrLO4NEDZpbFJS2lIdaYqSgJZejTTsry8FXP6XJDgTur+rvaPXw8ZCBBwPusbVIK
lwsQ+XTMCO7vu8A8WvX4utzOsK0TugiNWd75CANLejkNyfWV21viRYhQ4W4sO3XsmqSPQgbzMW6F
biXq1m2Jn0VWg4pRWArFa54D4jHQgBgyCUWmnvmeE6nzWwZQEAXyRFuDUh2Awem+JfEywXiTgAWv
fUnVaZ5ZB9gxks2/GumuYygyPNZ9RAi1p+ppiNkQ4+ciO1g382F9mijs/GlpTJij2WrxkehfJRDj
75NMe/DJVh4cwVbbvOAS6LmyFT/4Cn7Vm+0jbbQ1F7pFvMbJrogpiztiHd1+DYpZY0frnryv6d8k
yU89K+oJogZ9mIeRRJuPgFfTbjyCod2hM589Sk3DGnXTeJxuCBsP5v5MPFe6ihYhh4K4Gw3W7yTw
XKtG42lDzjQsf7jBOIrTuKy5i9mkhvZ/sBMHbSRes/fc2f0Pmu8PmOvhy0tAe9f1Gjw+qRr3RZsO
fhsD6dwQpk6t4Sx+dqoM+D+zxmwaexD3matOnzXP2V7xljpsn8DI7PSqAOLZm9J7kp2oewm0WK0T
OS6JBnuKKZPz/GkDHDXNM7JrWDeY4oulckRVUulZY1QazlzfuLiUiyU6pQAFKewKMecrzOB3IXz/
NHrCod7WJZnsCrRZlI+4vjkjE/N6wEAohrHbG1J2Zx89Xb1rlP+ePaveKthuR6M9hYG3uakBUSgE
FdchfHRovHuUEuvBLb5Mew8th3lKumKWMglJWgmDp7DnVlnOpC1w/8+5aE3UI4ggXg7OKxE/p3av
OVIlgijNEl49UbUgsFgf7MlYCW2XnRxjiouxcE3YhJCcM5dowqBGzrENNw2deQcHgBOmnT4SfS+F
Wbrdi2OrsNDuvEsTFZt7PWpya32SaGGimGy2xY0LBQBui9Z+6j1AmB4D21YrmdwPvIRxCOIH3afJ
AAF4Dj938cr9L5rIGBiy9+Uji3qCtiztKm9urX5S4sbJF3R0zajCqmgkrXRrLiN4ajkhtgXGAhcX
r+2ddvOx7yaAB5b/1Bjj9GXppsfs7oHPfivs8Mve8X64ANbgw39zptWl7IRDmSKfAwd5ZdecT1Nd
hLyCFZUolgNko1moc2JMn+PZJrJ6RdAmozwgtbPum16GHPCma07kDo5oX4YGaimrQ67AuCeBfaeC
0+MYFqRRbdgzhQUUBATwXuUnvqmV10w+CS4XO4wPIoxX7IgYWT4UFADJYF0dtd9plYpvTG9E4GOC
L3vL8YCz8OmRIMidOaaZx329OZl/vRInqZccQH+JY7YJYG8Z+sgXi2gjeP4dPC3P72mQnX72P7mO
evs+xMzkYsDsKWlx2KR127aDId/4jbRZw/WWMPy2C5v6fpoNQn3OLUf5tKp/YlqYmFEqC+bQlgHp
lQnC8XZQpaCwIwj+apPrQlijA4Vxt3bMXi5XwQ/Y6/43XVaVcd8f4SS9IqnjWdkJ8zwPSPyww8TW
Fkeh8IDg2EAMBYr1CL5q7Q7jGeWZYyqouKglBH6Xzh29XWUI9lsrLodSQpOWOGp0wVnXp1vo3IWK
KN+XR4W28OyXkNC2jpmrXwMyZ+T2u7CUqHb4G+7UzW9KqjXurgnD0IAnVPw3Tt231hNtWuz5W1em
EaGpvZbnQTt361VQw2BSHt935imAYt2QX8J93nJJfA2dCkKAhOLtCkpbeRyK/M0McSsOFZVgQYqb
LxeWh516gbQOw9HNaeGqoqc+EU0BB3+y36zY9YbRJUd6HTXOix4XC0lT+plgYoCFcKw/gKXlFyF8
1HB4IWzFmCtfMh8FN4dnyM7VWDFYTQFZDVDOOsDzr3k/Hb8NQ39YNlXI3ee7Dz0Hzd34vVsueJVU
3y75nNc/Cq1Z2rjjYuiWEOk/nH/a7mpiogD32qyi6DAlXE5RMZSelFE3bcLZwsPtI4+VXhMVkss0
x+JnmpipR++lETsrs5MyZZpxYa75Cm0uW7dSQlUz7z0k2NG3e/O6WAIW2c/W0aV+vJds01w1UohP
xuXWRVYx65O6gGdiZv+3cUxaDwHrSRZQYD5g72EIBJwtCDCqlUwxNJ8qjVrEeg5o3p5BcFT5Q2Lv
lLDA1VXtwBlB8NkNvmVIak3gZGvBOxWFLkZI2gsODfGUR4nYWCx7lOWdRy5pLTwlpDI4Ep/CwLIv
OJW3iklsXUcZi9dp3ai3aCAbbLwWhjnlo4l2KKfCIOlmrn+pNImr/737R+P3zphLjw7rr1LYpLU1
4FV0A4c7p4yBFpIlmmYU6DRFvqkApbWT3O5XVSO6yCZCKnWk242MHx8L7aJwQ4aOTXvWKBgMcTBo
b0i4gzOiIFkBhosKbT+WjAMQHvrjmnMwBUVf3UQpyIBdTt0FFHncYplKGpoLLc7of4hoS9lEU5+s
cwcFDg6PggQrxSyRWfMWcpoT5Kn8vDDnEpOKU0yPQIUDavEL0lvk42PqdlgnkL6gqaTReHCidV+1
LTbJHxbSpEK8EXP/zcBX0DZJvFr5OEgvvBFr2Ah2peXO8JujXMmLC3VqnjJEiaiHTFh7GjAZHpQ0
Bm99oa72xKnHr5a4rbZ7CIpuw8nECqcVIb5ExIdBEdra+G2CvBdEZmHfZXFlZbb8w7jwmP7V+QsO
zWxeKLpFjP+qaIy5MvWt5yVZLEQ8tjhwjPscZIExSl6cd1Kke+kN/b+X4NLkKXxixDZHQaHzl6wP
g7Iauq0Qnm2pg0OKsL9ddqlB9RamrG7f/cGVSomAFDZ/vnlgrpgAxf+xi5YL3a2HD5Hrh8LWWXfd
d+/atI5LEVR6tH9CkV+7R96UKo4+gwh1hsu6UST9gDSKRCykB8ETZwrEOBoj2IXCoA+5D+gb/MjO
plTYuqoZm9eT+84Hql7WaGBjorvXdAdqh0JdTopSqHwnkdDHcL6+rI2QoENZLEZ9kdoWakMK7ebk
T6Nca3Z6D3u+X1Ov4JSxrPKc0u0wrW5mtwaqpF7bmBAlOtlUhbDeplHXJWZM23TtusbxaJTKJiKL
ju9Oam543cHbhWBCF0fbuzUwdZi2Hu1JTCYNwOvS5/uUSYYctpIVRorX5m6Iug1E+cMsNMX5nvRJ
xiK/KnNvm2ZIhCI4PT0kz9a3+Gh/3BxScanDBtB61WqZTxKO9d6IukOwJ3k12N0SuvmB3CS/RQLg
HcfaWzAkjLMaFEW2iqD8MWSCH+MGi07Is4HEk1jN9s1KkTEPpJy15p8Y54jd0yvkSXa8SQIiSb8u
G0vfJrpn10ZzF16Q5YqOu+srIcO75StJUOgPZgPiNHqDeTlXiiMu6a/7sFIr4SGolWjGVpvEI9Zb
cDx2UGKoRDtv/r+jX3pfpJEOrE5gXKwLd/GGKCZ7HjVxhsBZJwE5/zI16ScyJ6EwJnFg0D+o1LOP
/y4TUQ/PchXqYNvdkBCY1Z1QGxt7z1ik+I6v7qDoOXrYRrzQy2gY1SkucO8AIdwmi30MSp1gtAo+
ruf4O2TgzH3xHN/afGXg3fgVucXnY/6TT7bHak8bBjJpsUuZP2NomrqknxD6WtGVJynk4tr8Imzw
HUgy3KIK8TlZmG4Od59A++O6uHq2C6IpPTi4p5mwgnxQSpkjheLHcVlZwYJsCjzA6a51e8vqEcyQ
4KwcVYF+UNMXBGIGFJb8qS7OUiE/8tv21X+3gSgtuBgynmIWEax9bwFoNKxIp5Somo3dsyQ4IHy4
A+wUbojxg7a2rAUXj1mRTObQShO1EuAbBkbK/DMLIDAuo0EvpYzVyroqbGep3DFcQhThv+1soIPC
HnNt3oyyDciF+wpWo8Dk4NTlsX6RJIw4Orl3+YApaihgnGRagVZiKVszIeKFHcs9vRnJLAgc4g6D
ui5W4rJ3Mp+hUql43iNnhm7N47THuFS9q+VLtsUwzuxQRbmpNAgpe/mcgJd/hQeml60vpfN0GwX9
bF9iUe/Zyw2NxsaX6QZGgMhq/Gd0Eor5P5xos/UBhbe/j7UnA2ON1eqHdeuNczF1j6+t9gnhMaUL
MBW6DDSOIMlFYq9I7CtZXnK2Hl+SfPSx590M0VUrB+fX1eSLSNJ/SszwQ1o+GQJsUvngiel9Sqd6
QBSEYUcsPzpAVajk0731vz95ItDwale2yUv4EJ22oN7V8nJANEj/0Z+xZryZqD4PS2Vxn55/Atjf
g4WfnI6P6JqAB4u3qZHqMny8H1hwE8E2H1OBz5v688jT1KTKdvjmaSZ6AquGzF3a/dGQIMl36p7o
Y7YDp/tycnb7xHr+aZOoEZlhoWbR5IWJtS44A3GhH+4ayummMEVaC0kTtsxt2gyD2OtM99cLHKrg
pWbQCv/HQOueRwhVkX0app/iHXHgjm8U92Tuz6ZYYSSvfLLls5w9Qw9V2XoRkdRmDzRfcB0qmdmr
UTQmh54v49KNAjuLnZRh2trXyLl4KbCAOfuHMnD6BlP4VbOQ6uRkK6BzFbE6SpccSO3q3QlImz7F
TTMUaJ0rmitzJm0LJHUs1v9rQz0PHhlqbKXaBbT1w1b1BblGZxrns5NOqVBMxxgs6W5RtDYKVV3/
eJdzRVJYgXT+2fZ+mkVVw52lnb5ANYRwwmRszZaEu2QEoRF8904sJaJAwRLc74KcL3krpQ0Q6TqB
Xp1mjQSmz4Kgnc4iTPb9vnPXIHHAtwOp0JTod2to3aNtyuWep+lQ4uLmvyYsSBnc0j/e18xNJBfK
lVDdo79sibZcRxg+nc7d9mQGRmp2u5RfsZ+H9Xt5If8hHesxOW5Q1W8dLnvtzctou98uIWr2krwn
VILtfx8aJ7cr8knFsNEHczch3UTCrnQGVJrnZkXQ10XHvIvsMJEbbN+Dc0sDTrZa1mT8lJutXZjz
w0f2rRUspPbUTKS9aIDbNwdRgwf9IT11+c/m0upkLGohfQwbCy5/Ay28I9rtTz1U7H5PBxO1/Dso
wEVTH27HvcFGeSGVUeGLABDCvq9X9rjijJa4QEnV471exmoPBsDIRD1+2/TQlrp0a/r08S+XXCtE
MDgXPvRmYz2fRViKaM+XnMxn2DJwuE/7zu8avPoNhhW+MxUra8+GUCLBjDhNGvSzvcgInCkdhI86
oTy0UFXYo1dq6GJz4OJdoee2N/JdiQxd2EO0sF55kc2ZnaNRXww9hS2UV1wbaw+M7zMdEWZE2G0y
w+6vi5O7C+e8RbFW4x03v9ylyl2zgpbxUFzkhRvfs5NFPffGOPI2qcESlqRTyf1mX6Y06X2m5sQS
zrj+t6X1yLuz0H12fYe79Ig+kFxQE0ccupqDiVackdnuMlqCNmh0PtP/9DSn4V7uHvTH+zqq8weV
AGMiG5WF6Yc+xQ7Mc9FIH5uvYdAkc4bmKb7gnSSuyqQneKU1MstjLnRyL5tTxwsvIRlL1MplSnm5
ntPJ6AQdnUlbBAaoUZTEkuDb8KwqmcHbHkVD6xGFEb1rCZXp3t7li67ut5AwQY6mC5ec2BIvzwnU
jwlHWRSDdnMpq7vcrZtygP0X8D4qpxyDz4eu1SRvw8NbDuEwsLp3ifzQsc/cJZPW7kfHys5SLLGp
mJ+fqrDhFVOaZ8J3OWHKUPAkStYgmGSIgVoN1p2pya9S0yXY0glQ9e4D2ySuv5DvtYw3Ymqb9OUq
EsR7UaW1JfL5yfgmuB0pUfL1K9QD7a2SzS0plaXztIOjknr5xOM7jQ4M/9wuj3poWYqX833+YE5V
sN6QZ2vOs+2wkEDoLZuVRZXO58CumBHz/bXuBWSw2LX8S+quzOsZgv29AZg4GlmPAGHZVAKLCiXm
oM9zztbNcslqQP6nanDc7bTfwj3nBQV9MYYMV9yPN05gKseUZwYt+j4h153fuN8QsfUMk+MtEcrK
ZuQTvchdMG2ghkH8H0X11osChj2EXKUHoYFZmAdHWxkHBfHrfULqYoaCwjvNfC1389lNRvlt6TSl
q3FPb2utmnVwbEzLUEvlyBc+XO4hfmwlTa2jrpk9/drZP4x5ss0h2EAKcmz/ucQt8h0tI/jHxwMv
cC37GQ6kxO1Tp36haqGWYWHkwGP3iAMqPK8UMOST+dlNYHXOI570pS+efXonWFCEp3zazFGPBIPi
GzK6y28B/wcF3cEPfJoMaN+FFlsQFB8T3lPKsC2M6jQRhD/GBHTVclyatFM6RMxYSw+tQzlqaV1U
QdZWyr+jEpIDN1chAHkbzO5ADkaeCh+92NQTvwMtpMgXq66ues6pcnWgzgJq5cjMEUFub3gBThgI
UUR5nntkn+ifH3RJ6tD/63Xfwh6qUJ+NzEPsQAMERIGql/TbPgA8p7CzUKu8tn/vHUNfbD9s2Mbi
jRUyy7S81PceZRCnS/e+m8KPP1aTtRmeGu4GtoR79GnLUMvdxHHffN52wuRC8QlcUQ4L1ezRGXdO
3YvtCBbR4BeD+WMeKYNfprNCHi2M9t5CjvXSQsXGc8gNozFH5bU/OqsPhPWiwqTHaF52e2z3kRGE
bL8IKsoVvXsmrOqA1jiSBtooMCGwbT789qlcXt+zBglTIBjj2s/GR3xTjg0MlIWPj0APptg5XE3K
x5TL/v1otVGZf+rsHS0yh8oGBGoZYepyR293PXB2SJRGYKJ1Mn7vkNoW+oIhOn2/iz2ZBLirM7xA
6tcCBnH3rKMYDU6gH6ZM1n7756dgEaf1h97pEFip3cHVpIyQqM1j4BXaz0w8YWuKKLbXaMWbOVhq
F8bv5I01TOWT960sxE8YtUFaNd7vLo7AHGs1kTu0l2Da3n2SfCzxJvv5FdBG3hBZHQ/uyO4qLEwI
LKWr5sgFU7C43wd5jnGT26nUX5WnytQatrKXMi7GySI8kAbzgmNZxvmGK7f4/EhY9xVs8JjOXRGb
g0bZNOtXuTTx8ECK03RbdnTrx97I0RZnUAAR5pf4AWmU0aS2GVwUORUnDO3wuaDCDhzx/t8jFGlQ
ggQUa+UiGKkwXkG6Hbi7i9px0DJejVF8+4VshcPxuuNCRe5xqIPOJkTffo7+293fxv2KD3aPFz/9
3jui9icAktvXtelA+qPuzY9tpJXtLjJ4H90Q/NGvIRyshPc18z/nOsRYYeksKwVDYt9xYf/ClH/o
CevPB2HEEBwKpU3nitzddjeDyWO/3qU2rLQNp4HgcRu5Rht1LhkzfOhjvXoL+kg5YoG2ChXHkZk4
CJH8M4ML8/RA6IchziuH916mJKqFnq+VlL9zlw2LaNyb8+vvrIHIKuhIhuJMpNPzkRmrZRFaerr1
dJr7lsNyIV6h+1exYPj1MzQIFLNJ1Jgyeys/qkpn/z8tQhzecUi5szcPPxbOoG2xHHIJvjwp/W82
ZrLAsRVBDJzhCcjWEGjO0dOU68XYA4J3NMQjniaXvDo0pyk6PiY8N5ngeyis5dvR7/e3KEHDxa46
4U+6dbNuqobnNNaBUE8aW3+yo2TcrxymCHXJkK2oV3FQDWHwmuG87xU6yluYHPTCOqRJRJcZ+G4O
lJyGyPz9bwq5IAGGQ6y7/sJ+kihdlN0BT9wr5jCDKmJX/57n3T0VLgthNqBiQpwoNZa0JJqJFL9x
48/TuzliUdQeOJpUmmc2OZ7T9tmgGavvpFcIDm6WISVZoojv8n3pXEPXCftcIjJZ+E5yZSSXZGbz
wabb3dirXDoQpGosfQX+KPlvML90vgqxbKPiaV0CJIBF/MGy0/3T9pMQVVld2BwY3557hW5K+KxM
50LuUyKGXB4vLkMBSBx0PvK8zFbb4b4IHTb6OZa2nj6ir14lE91nmvzKrzWf82Sah+ZJNO2xWfC2
pixWDkZtYCcVmgocBx4utEyobZ9DQl01l9TWeApsq5JWJBjsp/LonpwIPe+HrFSo9ztO0eTrbFg6
fK6/KffzCPirYOQc4x+7SC5f+rv5JdxS5U+iUxQdAYNMRiApuZ9vS7mGxnU+39elj2BjNXfG48QL
ktgpeXiIjSdBp+gwmrVBgg6zoj/3veXNrx363/mvKJrgesvjhEJptWc1CynEfokpEQG4H0Jp+3qQ
5S8Ff5/zwPRETVQxrJJgntVkwspM9tzSfhg6IH+6hYEPXyP04ie9aSa6ZfmoEOSqDV8vPUkvVW0T
3uGh/FmIgYfL3i1uvTWhOHw+64RAMDnnGwIWFTleCmpclm/dA5IldRoGJrO0qqoh8+jtA99a3dEO
eHbjPPpWwudpajE1k07jDA3KV5kTuoRMEDF0Nz8PigoTU4mDDM56Rpw3K7iLOw13h4VXh10W3uA/
6Gx9QL7jBK7rA6HSVF8dFnyxZGng1seg/8QjO2GWgO0i6ygvvC4K7KBQOzfuJsqHrMYzCOxkhALQ
ufyu/UJc400lXRJCkMRm26lyHcXRFkTWXN2qsKma/6f02daWsiVkkDpbHcrXTXObjTx0BzLqw3dP
byOFy3H/vRSjxUMBL2Q9Cun/KqDe4hGXrWaqLLJ/koxeminauXCQzj5i616YkuCbaQrZctKt6smY
OMT1cC65sca6APztvIUzQ+4XkQ0P/hX87cmn3onoUKFCBQ/EboUv/1iDTqAB32UaGXrlKyQ9cLWX
karlaUtqkf37nPYSyxFSQy4qr8sNn4bOP7xh3fneO2HYFHs1SlyxK0P/94OrIl+63rZn6ZS7/mZh
ZBR+2CURK/tSUtcr/cCpWSS9zPwNUeInDKP6ct66X4ctxQrtpqMyQXUJL6ZmdXVeIYCcm17ivnfV
iukHzzRB/gFLWiWaEgN4Dq6XbDJZVB7HXVyc9QmxD2kmMpnZ0ZkyAb4FECFzOt3PkbAB7sEZclgb
2K75EFrrxMCsCtlNnz4B0ifgTXdEnIwb4A+4VEFL1kbxpEJ4WMFOjXjt2w0zU6rMTdPv20nHIyYa
CVbvKQb5qM0XJJl6QsnjiYasMAtw0UkZyCxboIlhYpLl80SPvdPor6DTmXEEJw/yugWd7qTvb55i
fMTTv84vZ0Z5nyFf/BA3WiWHE2nmVMFSeSjDd0uTHXyWZPXx0jClCwIBD1hHaUxF+T3DkkKnWNaF
T4KxIh1he9TZQto71KdgU68LOfnxpiRSCSCL16dYWM2ULC1dJuMo1tk4FsnTwmd1gzxImCvenRcK
SMKbCCodq/qzPvvHzRePfsQ+g5zqLkaBrmky5C61DvJE5LZVgngqiEXFBfmjI1bqg8P8UywFRQ5n
M0p7FLiuWbPVzx2+Z0cZppz3bhDseTexAEjmkqB8/i9ZM0Vj0unsKP6MrRKc5ftKQwHihEASZb3s
0gHuuPbpP/fqb0l4y8Pqz818nXRpTRPX1ueeLth2ZpgWF0X9sUpavLJ9iA6keQwv9tVDrqshUVGi
Aaze+CAlPp1OQ8PbBYbjT1v6BL9KbGmDlC/75HTtuw1t1MVmkaIUauMPF5UPBf1XWC0YvJCpqiyC
bcwJIO5VHImjAUHVPJHh8HrIW9/9FKE4niA3Tpav6igoQ0aRyIdkYfYc7LZjuLiLGY8WVzgbBP9s
LHyCB9OWaN4TkVsaqwhe+9uEqNVCfwUQSHk3J8Qyw99h5ZdFnpf6MNrTxxV9ZDvkaDtA8w1VyjSC
Ll5iPhfdtOQt9jy+uOJtjvK90BshAnw5E9x6UDcayhGyjDL277Hp6+R5VwAXWRu2JoXZZQZn30YN
VK7IpFtRqOiRqDsO7M+wdsFam4HN53qT8L0NYNMzIDRfEBBMdcm+Ybm6W+cEpJUiQARu2LRb53TB
GXQy5l6iq5SBrKx9mxLWUepJ3SBdCmUyglDU/hvqo5CKnhpGPgWekLYe/FrgYCA3eNocffvxVd0y
xXn9kzcNe6DSB9jtp++eLhS+Yhqp/6EvQG/+oymxDWIFWgyFxeMwABp4ypqx99doCQ1PGYP79oTy
eN+TMu09NwmfXuW8nADcBdLFYWuVGaq1UHVJi5CmVYea74gsxGU/VS2BaxmFH93V9y2bLUajE4Jb
+DAJEvq/fxtdqFg2GbM04Ksjk6xIASckVgk/7ec1Am2wXGHzVgWn5DidRtVhPCqmhwgNlyU6jwj0
SEavfjuwDmJvkkjRIJGM04h+o/IWxRZhRGhRg6ezKOYgQBHHyVYRGP7oysNBY5D5UiV40Hhmi9EV
utlwlelyc0JN9OUYnLhSjrh46e6kM4VhWlvO4txMHauZDLASYNzTuUU1TWeAlZTWiRy4xTl+3cXe
s+vTofZWuYH9DbP+IgTUcg3gfG83IekeP/EdBEHVyJC74WUxYfOY5Q+/7hY37VlRH/DzmqL+HLKU
QBG3SJDwtyYMgNPrq68MaqVTgiifzVvCq/E96hIxEIVgOfqvX18W2wxe7KZakmSB4LGFjMp3EFQs
kWprbZG+VmoPzgNYwrmfA3LV6G7jxv/yL1oiPxa4xaKwVaKPMiHviy6N6ewKL2WoKdNIUen709ZF
1HlzrTBxnjaSY5dgp12budxiuVv9ID2wegTAQkJeESxS7SqjSArvmHWdgSqa2iIsJQMStP2ygJki
RTbTK8xD5XCZA3iqJ2aUG82xFmL0LUvK7oE1EZxtbUrTH2ZV6qNf/JhZrSPnTXQvuEo7YLpE7HI4
tHwMiCJ5KiIhGIvt6TDMxjUSXI2JdE2HY1YDlA6D65o76cmJz3RQ7ydfb41VzwSPXEIkk2+4IFUI
Y8HUSdu7w7W3qfR/3ihjaG0ZtLYSXPxyJ7lpqykYNQUP2SkfZ+zUsu/lu2BcfnhUyUstMXcaUFuV
IcG8BG80szOa3tPoqxvCYA/1ReoYJyE28JR19G64VD64fT+u15W9O2Kl/258s+u9nR79c1jvRerD
p4QkENFmcmvA+o0yiNtcDqN82zjwUc9EIoZsXYHAOZgTY0JH7Vl5XcDctNBQYyisca5OF1oT22ao
66/ixBGFTXHZxx6eqakDqqEE2swBeU6g3HCFvD7aSkHHbOFSKL5wN3gsKhlJuqqBf6+CxYZ9sC26
UgfJTTiiSE50TyCHt9Jty74wWF26UXeSxMYn/LwCRRoI8RtzcUyTRhoDVw0in//Nq21V7JFWQ3zB
4+M3CHhOA3rwipObcg2pHsoy7Rlg0BNbE3tGM/+nTiTdsY8jqcYRgsYHuNqUSq4ugxB+BBI/9Cds
9fUlJCwybOPF2geuYzqQOPv1KBb0xS6N93xRzuEmdwkumc6nPONR449YhfLg4WM5pCKWgYwY2ELa
9D0g5j3lcbVMPclnwiBJbNl+nfBLXuGvYi8Ja8ZJuUjM+iDFIH++m9PdCeloPl73Wh8KrRk6VrkV
8OzXFJEDafTtfSIoEk51OBmCRGBkc7QaWNPPlFPNHddEKbFWmSV0ZZgxcBBCsnJZukNDbroaD7Dr
HRFbad2FCh8heAbf1Qk5SDog4oEMGsCiGSHwIO7zezCY22P+fK8TOekd57Sd+g4M+MIEGAaj9Qxg
X2RU5fFFONe22cPNyZHAoFnkQE+xqj5wqg+fMelC+sjWwFF2HCcxA64+T2hcKVudmIIpF2AjiTmH
mofUlGhWYPiuP/xEfdLH5DAwAThg3iHh4eQh4KcQt5sMHukRV7VBYktD1zdw4mr9zojWsweNeHsz
EVvwrJyglMTxo2yE3nqOj8SrC9AncV0ItxfbC3lKxXdcTkHfJQHqjYLKRrREKbmklx9gEsp8V8sS
a7DjuBjUtzfN8W2xsfBKtZPrhJja3XiaHJI0ufgV0d5fnNq0VysaBmVhr69XcrTeiJF0sz3RPOjl
hffOTwwphok6qMxsl0mgMQMFiXLz8ze7TfIXGdwcsWyIONAZM0M3cxb0dN4Cioa97q3mMs29Jkx6
LtaJ1xd+VuAjPGP2x3HmcFWgVVpcOUaVqYzCno+KGdt1yBOlgONYjOKQgdDR7HIIXzsOOA6GnN0K
yKGyu0v3qeqVkrQtxRig8RoIOK+FFehkjJ2B6NwbtssvxkxNkG3Pr3fAELGRR58fM/57c/fYlPnM
vALVXjTX5HRzhB4yswEzR7OK1KYLDaoj8qCiUlZrUxUGvA741QYjxUx+MdSj37kOKwFtFxlM/zbf
TzEnXtAc+wGtQAD93K+bbmAZT2UdadmepAIkNq7G/S2QBj2YT7j+HqFI0mXYmfBvOsOwqUROoObW
z4LXcGiEv1Tu8tRbN8TFrgSViwE+eyZrs8pchxk3/57Aw85M1BJAWghk2BeKovOVNPbAliSdLVer
3yG8T9437HuAirPQk0JoL7l68ViIwYYD4Z76DNi5+qaC+sJZblUie18w1cNbRB59eJQWiy/egQ33
/0tL+FCLlQY+TwSg5Q65Ub7WL07zT9VLPhtWK9DYVFkTohx0NhI6HWgA3vaVDRJscJqVzDA4D26I
8XsuCH4Nygk/47diMFNyTrC1dD9ayxUZMfVPS5NcRLfbjK8B+RSG7fCmSZFwsJwmQZQJMzHlHuyh
Y5IguG2eDFw8nsEc11n5hslfqZhMhQM8e+JlMcvqeJTrdxHEunaGV9CY6tcLD+K4dzyMbaElANsl
5Q75o/wlErPD7ImjYzTsDxZxnixktA/CGPVgHf25zClRVBqyUXQHmNHJkAy0HRhJOEUCmFZJpAvq
JTF9xmXQSzGD5GprDos29XXXRgCRRQSbuwfqnPBco8gW3xZYGmya7hFpcfKWunyxZe6d19xsPR7p
bALfX21VcTYzULhTyPa59n6JnoIIUrppWIaMf6OSbC0I42hFJSl01sP8XE7lY1ua/NpkHAWuQ1lW
Qq/Uct/bU8og/mHZbdpamnJyzCdPZFi4/8i0Nt35z2kd55apQiHE1AkVNOAu5eNpYsGZd5PwrhmX
k4WkIdYn98f6P36+1psHVXotJvaE6oXZhD5d86UbiwSGAidsybGNxnukhxAHxUa6NCSnH3Tl06GG
PSRLZvoTXOuBV4oVdN05kOJh76L1gpS+19yGuKrnDzhnfcG8cby6esnNQdZkKY2ASTh9uR8/ROYS
xLszNHEmhY0TGHdyX2EiJumQB0vdGkzQ5RdvWcfBIRmDmPWdYCLyxTljPiD7diWu42Lijla8f2iM
pYJsJSgPqQoL+t5qTjqOqslbVrtDBxpYlaVtA2Firj+CwD3B6DlxFqVjv00G38878UFHREJ5khX/
2DRiBQpbiiIeV4XOUXUnxm5rGQoggWULrmjbn6lz+Gl1CDX9ypyqwRoxu0EA2piYJ2bYe4J8bKKk
NCAYCxH3uR8Qd+VrB8Z5/w+E8v/5FhzGnQx9M2SOsam90dQDspGnWiyBfTmYcQXGfK3XsUiFtzX1
pmFImx2DogefE73oVfDtN57oOjDxMV90s1qXvwdGBZGQYgnbvcFo3IQHH3w6SDHGzcNVMmj+doW8
oAu4sMVF7pcmgg8IpDvElVTGgteEuw88IIsfEfihyOAgSQNZ7ro9Z8L8tMLh1uk1PxCda9CL1K6V
rxzVZQN3cHwtUe7bKcdme9Z+3FMlT/6/5t00gqEBWAWG9WM70J4rn80Pj77QmqjIgkr11zMHDFc3
PuYyA5ZE7Ucjz2HF2vApNJcqu6VmMA8v7c6Dzp0ezFETcsQkfhmkO+aSngUV3mjn6Ok5vLUpZWAz
DUbvgTm3jmHuTpp/iWqAxWGdnDMCJH9XStYjL3ymm084DfLQluWXrnkBg9SFrciClML6BBfXriP3
TEC4rrLru7hDLgGnF+M2J54JGkYovKV3rR0EYXXpgW4MPoF2v+ybFAc8i8QO0migKpOxcICq6Qhf
ad1+AGniTHfGrZ3uGSnj2MK8C5n/2uiY1A3h/+I3jIv2cIOzgd4i+P50qfl2HrFTj3tXHwiIVwMs
gUGTzNMlHy3VufvWPoZXA2/eu/GflNBpmkVKiE+8rWupK2C2AYfMc42KSgPFBbmUtMZF64QaIGAD
/dFr/HgvU8J3qx9J61GYyTJK+KsbNCMsQjZ163tUPByji/2pCTySd/k5MM8uk569/HtM1mNfPHrb
vt6VADWOPPXnbfYN/9rWxYXZBbk3mwB3OuAjhukP/WB6abdHsgacAeWnAuTuNbFTtXtYgVNEkJRa
rqtqL0NLt0xEw24vtGH8cEfVZCs5Ob1LDUqNip5/5Iccdua79fe2P0HdSc1d/2vdHZRsaGMAmkjD
YdnhLpCdaA2C9YHR9IB+5Z2drqxNa3/GB/b5EZEauwAxKmEjw+I1iStWAYizrL8x75CEsADS0i4q
x0KiAN9+ULqjsCaNVGs9vDiBpoRMYIl4/W7Ij8G+KezJABOwaIOv7U50gnv7YGA8EpOV0B5Fqc2R
oJM42KlPGCxYttim6JSfy6E+xZJUwkZ0Gb15YfxZR4QEwvOe+qclakbkNa7a07qLZMs285eVaJSO
N2d01As82/Iz5EBEEyM+QuAEcolG8fcFcULXk6+EkrnAI0vWr+fCJTFr0TBQDMfp3bnl1ptMs9Y7
xb5lL77Vb4KDkoe2r6Lon9S1veEX7BNOxZkD6SbTnX9W86O5+vE3S8r0cWW6AFchcs/2bJdpMwct
b7v16HiI+RHcq8i6rUDMUL3Zzqv6NfUa++TnBM/9EED1VR2r6qzdNLfW2/p9IXRk4jhNltXAHrxW
P1t9aA77vXwtL6sgTXcHjTnZxIbHSMpNPPskQUsvAi5893aTW90Lr06QW8WSQ1nVxGIiH8zWU8qa
g1B4Sexxztb1RqOLxAhD7dxruRivjJaB8qR80hl+ZbDGeWB5/Yb4rIqGtUJ8U+UtB4NdQohn1bnI
vdcsIXk0nVhPQ3gIevIjq08FIcopF75TwqMXQPsLvymJQrR1nPBHNeJf7KhOgseevczIH9J8Lmc/
l+fo+VHic2tED4AkjSJ02ac/x5h71CqbFSIrGiNAp5YsjRVyFm/+pjnkZWce2zvzZeZ/lF97zXSO
0si6aD5PdDxCMLEpAqn6Rw9WtWzPf97S9Tnn6YYf3+UhAGUKYSrLxVPyBJ+u28gAt4MVbup0Ha8L
qq6IQaiozBV0mqbaJFZsdfraG99eDJjyRGw4Kh7TfgCje/SAR1PMLYZzQlcP2ZTgNj3Em3Rchrhy
6WT0P6Q+Nk2+IHkaXwKlvAMz5RVXu2ORKgN8qeR1Mj6DHRWhDlFxihPXCdIKuUpDwnuYR7+YA5tg
JRb3J5vHHigL1xfkAh9XPvFg/HogixmISYPkXE3ta/0WsYyghEo7KlcZI+VWN/CnOuNzH0yTlXuB
hf9da/iPOwRunUmkcxNrn+Q438VFWqRte9cFt+eNj9PT1LuaBcCYeq3Wih1K1sVsO6Y8MqujFKSv
3/wHd8QMDOGIru/FFTCDQfixcY+flIXNNCe6fj3UF9W/seIOTUHfKHDNuJa/o/ZYqg4OwlNUgabm
jz6tFqodIVItHfCpMHm5V6mVRDW4ldSmv2ngLBBuHhpWAQcSOznf272uu2z/5H0f6qs50gjMU43r
95goHqHCPPhPVndflnoQyGgz8BTD1FEGjAJzEwGKa2yasA1HaK8rVaLWuCkeTDlE4R7QJbpnyZmA
hOsFu1BUf3GN32+TJg8CANJOIlzHplNN9T9eiYEB+jAsJGnsBU65ZGRVYs7QZ7DSds6VYex7YQqG
FndqQipT5/LjURz9FisFv2J6wyS3yuOsnZlzZztGg1tX3Z7x+JVqqxlrZfUt0vL6jys5ISHWgOhU
94DdE8GuU/rnZCZ0kQYXi29oOnYV2oKx1O2jzkzsFjSXr0Fcp/1Yd/R/BaMGQicNRpL7czQ3H7FU
OUz9mUQnkEc2TPk8YTi3GnKRnKLEzgcKK+pjXeP+PGcjLz2e++1aWt3SpErB/b1U67gCmXaeM29N
afst0RoI/j1yHo9IyTKkYNGOjukKRYq0vCf5W1fTqdwnBTVst4Dy0vKWg82IzUENnrFIk0QM7GbD
K1t+BVHh3OdHWdUxzwVF3WwLgOafbEYarqN/oqq0aD1qg6DJtI71gJ/F93Qm2pgFohvQlKYumehd
FbUSwjRzddGjh2mElDRan0eghMgD6gksAE4Oyc5TR2EwvjhwsJimwq5GvVj36Gn51HU2M9QTGapu
ccuvjHHhUHPf/U8XicQZhBi5+4w3PH9dNOSRIRKRYe+KUMJ0/zI8tbTh0PBwEjqnkMLoihrASV/K
kfLXEttNOuEAnZzMAgfA1egtAcPd0ambeImUqjo9CGvpOBDdmVRGiaGBC7pjX6qvXmFz+09EKZba
TiMmIYQcpZT1PQfBIgljq19JmmKzokbd36HQVmOv7gJlDttACccIqnU7jKE2svNxTIiN13gD43DS
BuCTYEQqDXzZYHx6mQb3S6csjQ7WZj7uD55TSjYYBLvLJH5KsMEddadOAunewBvuEW/sy5G0UYwd
AOCtnY+MJP3BAtmhEf5lEaEjoEgp9WSA19nTz+9SR4LfH2JQHzQ+tt0CogWmKM/tqzsS/cthAv9A
3h9fT4Y32p1AqU4EnSlrWMm74mT9xxT9r0LAOdvM7HGyw5UTdtoOmpjeK8uaMYiPsdCw5tuEF48G
Q2ybl0gKGrx0rWG6qiXh3qEDZqDsG7s/lYJ8OslZqCZ6ZQtu5HJjeEudiXcx33Bcfvx55RrS5iRd
D08oreihw2vJY2x0UsUzv709L3SNoPXnRnHIm5e4XmLQ4SrrI0o0PXNeO7J/RtPW86/mNF3m3fSu
XHws/QsL2/T9w5zuInTodE+b3QMv2W3MTyxRRAxJiQcmVgMgF67u1Cw5FCz8DkvzDOpIRvOx8qCH
J70+g4yN2RuUrV1eVpBMb0SE34nAs46qiXTNtQZTqJwNpH2u7YjZ+3QgTCryXcT7s3ZVlIbflq7j
aZN7+sBBSj60WqS66ruozXJDRhTcMRdxayZLyt9bl6TubvoZI/Gocxvr/754uzcVGHezuDp58CGc
WdCRFq84WNGSruF5k1zLlVeNCq8nyBk/C8EXWKlQZox0vNz16Ag9kYMD40TwHsk1LpQ8owQaB1yR
lNlg5Vkka5kGgiviOQHMWJRVrr58ag1lrxniZRvz1tBWlK1uEgu0Um2kGDnsoufXXyffAXu3Q7/4
+Qf9UgyEK81TskiqxewS5ypJdOEdEfcMscWsIQyp2RcHnWwAu+lA3S1VDyY8Nnwr02Hl20oUrjjz
0jJBmnjp1r55W9grHHAiaf6XIkufWgvBEHkkYQLO1nrw9sTpYG2/1WysznzL7o3U1rDJNtRFgkym
K71f2+zVbbKsyIveZr5JWem1ph3aJkm4v2HWDboyxm/8YJmhXuqEnIGXVOwoqbpRdMQttYe8Gei2
wHyQ2EWPzyEQPSaR+W6eOvEcZoasWtvOkWvlV6yXL94x57lmbwNwjp9OvKNS6M9YFBp1iE2wQ+FY
18jQ0hP3uPS50ZYGwCSY7kVTwY7v8xALGSVVDEygUFBIBP4ouAf+XoNSVeMbKaJ/ZEliRO91zEY/
qJLSlmChqJStdS5YGda31U/P35vBTn0JIjs8n7sy1PpWSaV4hzqeqWbDmVYMMK9PRZNvVQy4YsjB
j36vo+Zq2gWFLgZ2OaBMmwbcQtiflCsy1dDr0Insidi4yR+mHjba1gtt63JGcddRj9ffWa1fOYFj
6KbqmeoQ4UW45sBC9KkCVwBvIFJaGQ6utjU3OL+XNOsduOerhfxZbkr2NbnW+71n5lGpwqvrmSGL
Qy3Ea9+Pfa6ZeFKv/I7TRjWdRdnAuscMDYnz6OfN2lDExxdmTx9Unlij3QoPiufkfNjQM5JwIN05
/7mn/kqsarKZsz/J5HdtbI2ErDnH1shyEGLTVuCDJOxmaLgK21f2RkZQ/O3IQmMVTJ2CdyMOxhbA
TqJAErR0aT8yq61WJ2U9FIGSKP5jpKMOqUykQK4ZoRn5sf2YKi7BnTAW52ydIU7Sxcb9YLxhzSoJ
tBDxf3D6SBujmzRAXR99hzk+3h7Rnd87Fjuvje+ykJXG1nzx2rMPP124upvWf1i87K4kiRrop3Sn
Y9BoAhCK/kxE8PdMZhFQzL3Y98szfRvidcw6j8FcXMWwXqM8zoa5f5/+5Ykr0jdPVxtame1rgycu
1ttqURUsrbz7ENRA4365/Iz59GaTJuWhamhlKKsiap51GZth7chodpS/BjJ2SXDYTbgmQ7/7+cRK
qOG5f1FXpqaLd1RwJTj5JATRTvJDWr1uq/a3gJXHxaCkUp5ifk7ssyRQX4T97rwhaKpBEQetdg0f
EgHTewddY+W208PiCup/UDCW258s0LQCYlgtKNo41JURC9ZqHcAYomppnbciWF8WO/SDO8hpDxI5
8IPPKqgzpRus5P7NfA/0O9DTdQr6YmQzG5WZki/oEinmBm1E+uVK11CoPVmk0tXtYcUksdL9RXIL
eYu1H9PJPDfQ+9Qn1SrvvegY1fHlLFTVM/qZf1biBr0uQHI31VwrYfi3P1gfOBWIR7JpH85lsIGf
3LAzV+/yFnU1jI5Qnp0GGMlcfcBr0cqCc1NF8C2/jmOUXMBnkuD1n94tCwzI04JPLkpOPatjlceo
//xk4+ZB/ERDzR3eyMcjyfTUca5JOFwFWp2wG6HIf+E1SS18YLLKklXh1QYOQ5F4KMO4QMBnu69A
TyTY+78AUPkd6IN2q8s1j8tgsQiGISJEiOihyHsoxB9/KJymibcYv4+72VD5eBu/Ou68lebury3E
znK1zeRrztJChUdvKqEOSyv2qAKp5SKJKZEB5YhKUosDOvHNf5QUjRbZofeTi6jBOa3/PDPhgzQE
zUwy30InlFbMJ0hO8pxAG83Q2JKBbdPZZsO/8EztzMZiGNRN4BVDn/+nghECyf3cS9dhWlqqaMWo
0V2KzPKzBEZk3Xl8rrwf1fxeTiSNZFKuH2j+vGqDIV67/n2YkoOSbPqEMF/vig0ZB1Jx1DMR82xW
dBZK8IBuCKQH5ij6DTEgwrujYE5o2ZxYlymCArtoXuLlE4HiTH/QkMXwJXrH9pEVhQTfPdzgiSdC
N9Zen3xo8aVwsqcD75kNBoE0Nl61y4GdWbiO/ZLbl4+KECJcFA4hWihxKg8V/NWrz4MQfYWc6yUJ
kBtjduiisqk74Y3wAg3tKwInRN1yvXd7fJrvOrRlAmaGRjSLJ8DVEoRZE1fVlAX4ha1g6fLAOroG
0EXTt5AZftdqTC9vLR3F6uWKy+MDHtis7PMxrUZRRVnH1zfmJMqPSEHTmJIfOYVTol1yohThdulJ
PHYh1ZOLXwqd/1dPT0i7JkeFDR+O1XUwfqr9xxD4jjGuXElkvyRRXegKKUBMJ03AsnbFKmSq6nmd
6GjUFAq5sVLE02BUxkkKQuNI1o5yj5fqA79mUxRF8lhzW3GkD9fWjQ8BY21O0P1PROj9yT44r+4X
d+3/hS+9lCZOWNyQB/rlaPWKLhC5UjBka7NrqkVZmXikdGJE35SOVqZ/TU0/FldKfFMbrHMYxP54
i2Md01oUpH1oevPaaICYS5AVzD9hTk7qDhI3vCqpSp6dIAP4kZvr1lkXH6CNgOzo24SGxs9MT1jN
VyioE4kczwY2QneC7V4x62+H1scb4gxDFS09DDxaiITekzH7jKWD3w5gMjDS6Dg4lu/uhdQqzCph
//GS+ObjjZZ0p1K8epwiL7H/ZQv7p+V1gMv2CAs8TjgJJMwm92I/P93nT1gf4/iMfW3agx5jURie
YDSeIkPbSxvthiq+Nv7ZLRzsFJVBAFNV74T/Ai9yCu0ls39XY3O6wI8yMCu7/t2mhfydKFUkKTMj
qIiCCaUbs1Zude8HDqTEARtXuJ1qkP8oYjPp8an0PGamgVvkRQoFBIqAk2qv3a7QyPjy3JGQ3wXB
6Va1Q+F7nffXDGEkvvxGMCBDAXtWUtVOvGkJAh3y4pVdjI06AaFDhzsMg3b2cQTAtZAQwXvrPMbM
OyxnzetsYXf+zHc5rVFODEQtaVwJOZ6A3vKG0znSBEn22iWRmG0mcLFknm7GB7SwwI8ip8ABQ0PZ
5hZyfzXj3TZuO3Zu0e5jCHokXVzo87DGq9XEaWcjL7KaxdTQUzKmomtmyzgjT0Bu7GWypO13kBDX
Xr13mkXYP4ze6m/LQkecKopKaSMWNiiBF/rqkfbdVgHHo0qIBrZLYDgRBXIybucBfQ97afnm7DSm
zTw3pnoLs6ClOqGlpg9zvu+5z5pQI6WRO3xaOwOe4Np80z73ZONZpv7z5CKGeKkEPvFCdXltvsT+
fEGz2LJUTY9mcaX1mgpQodnGdIwLq57Ky8n/KoUtSzWqALcgUnvSGO0/tgsc0ptDG5lqqe5y4wqb
2lRAnJpaySXiaOZvFsWgkTHRxMoWWQXaRxvk7muWEy/nKCMa/25S1MjfhRChnAo2+KEHcoo/CcAK
ko6A653ks52dTJa6Vv4G+tjt7VsNcyX9z0yeLyeYHUxkbiEW4DxOrFuSSX3wtS4hH2EOtcwU3iCA
doeJnJV/qCgkKisH/a8L+TiFqGFhvcB1IbJ4IxqR5H+MxLXUv0ropYtoaTnCCzyTjtlncqToXKb9
SK6yesDzTE6m8XB7LJzljlF9fNatn26TJjy+A9NkcAOqoujAIV8sdqglqlVyYyE09dAMiHgFEQDf
cSUGR39UBBIL/ZuLXb32bHwrSXSrQZUv6hRYL++mRlws1eirTqbz3BZIgf9y2vJDlcm0B/BlnU0f
sq202tEJih+szAXykHEK65akzCL99wCOi+EqOas9a8RDp5k8zKtjgjY6tBWQb/zU/hzFWr7DkxQ2
ZJHn5brsyap2vKZtM7OdL1FO5GQdTgBgUssUkwr4JPJXMSOM3kTRrAHhUjPrhXJPFb0KYnZOMdA+
KqX1TY8srdTVFmMIVsbWEfb061RC8PTgPo9m8edKoDLJHPqbrpdTJfGVS2pDuzQebj4AeNxtQ55T
RFNrKRh3MIj5c2rYfgTi+kTdhhjQM+TD/FdIby+XiM+BbR2EV6OuF8KbY1JR6yPKakhL/WF09QiS
EK+bBxYNcpgoysqOlPd+LhngusY1gJNOAJOsFGUMKyV0Ds/yEM4mJLJBStMpkhQ0p5/yY8/0as1S
tZp0ufvbdgrdWZr1+ArjYU5InEjkyYCwEkUCe+jX95mhAk/Qx4UFyXcJ7ji71SUiMNQDl7xM6OwJ
zE2HqUsKP3vmEciINboac014YBYOpcUr0zUHCbWTfB33iYD0QIu5eGQg/of5UkHiUOlIMqaQXUkS
mUUShP9dMkz4s3BZboQaLqPy9AzC/1bLBxPX4q+gPTYK7yTnsMlQFywC/WaAXn86DrAHmQur/qEZ
13LCkFuHdP7NNX2JsmZq33/YoNwpEnl1RqQU5l5PuPjD3kyJIB7Lh1BitENLB4/YiCHD+Sg7i+s6
KtIafv7zaa0r2VAzjeYCb9niU1NswsgMDPv9M5MPRyjJKwc13N+pWgoQhrT7GSEKxvE5r/goNHw9
oOQeUBRsU3kCnw3QGLWIeMOerStDw1Ded5A5Jcmf9TVshSYhw2N4SerNE/M4toSok+DZm2osIFvi
iW+457Wd+Ej7dfrmpE50ICUH2G88ayQqThGyUpjvXChiX01ks+9zLi/qfb0JZOTPS9p2V3Uu9K/d
reDWS+IMSSnX8UXWocSWOnWlZgaJsdgtFyyrq43j54H/8KQUhXT8EYCLwamww6Za8jX2sCXPuD7r
iygdx1T8YU2vbNjxxdDwARvkrqYCvGasuvhZ5ls7S6vdqHPHRi2g0nhOEIMZrUvPenagP8jtNQHi
/uywXeyvVc+ETFxx+HTTfpTlT+qYnc1JQacKjslw7GoAM5sm0nnmvfNajjFEwbPo+Ox6jd+iJK73
PRrz7rDptOo/k1m07GHkikf9tje78S0VeWsD4S3zjkPlMfD+3kMlP72jxIYy3pwDKCPkkptxCg/G
WMRyCV/Tkr+y69CVJ9vwLru0RthHDQeP7w3/BLFtCvkdXhfFsxaa/wbmn/uqnnae1zYTdEPG/Jjk
lH2HEzc/3n/P9aPKT/Jr0R4UPLn/SAy+AJGVsPyUjmpIMIh37RU/Ey0NJUTu2TVPPVMJjRk/ApfU
F+JQqjpOBmPXQdbg24vdhLiFAny/GcpZUVTMgyPIADXwvGS7XWS1BR9BYhZ1YkbNQst33PDTeq1h
KpJtHHLWPnHWAOOwG6bOPb8NBV1aPH715V/9wZp/TP+A/wL8fLm+RmyB2kePGNf3zjZ9txBHFeUC
MlRhraNz4yYmWj5f25vj3dicuSXPFPkg5HfCihOXqMAIq9pg6HHjJZv3kI5xoi1k1BR/ZJj9+gmV
ngdaEtkD0B59boKZwiuxB7989QQn2WVghg67lrTVnmyJDkWssX4kgFsUbKUKoqO1bxKxE3EctJ//
2L34LyI6KlbLiLhtmc7kSxxXhlkP8I81JMdC2Iox+CPacOzFqDNP47SggKitCzrmLG1uTFdCdLRv
dmpkhtpLZ+X+YAIpz78hMRwU8zIYSU6bauhNUoykvlrACpMYsrjcGYhn7hbItQAuq1oCtVvC5aU0
1KAmMLm/Ha20zic3vDtFjs+vdXiJQFg8MEsHiH3O+LB1zv7OnFfc4p/sTrMABPQrR35Kkdp/Q8Fn
UrzINVsOQ4pqXU+LlthwvB7tAvNBny3jvpTkfehXKgTOrP95GdIXL0oj4r/9zpnw9keJo1a5waA6
9r3We3qlevT+DN1sjfzsDozFbKCTqywYqMGubmbdptwrludj1lsd03MNvGToRjboRKyQxoja1HH3
3sb9nFto9nKkIEYL4pOQP17TvE3K69twKpRF1gEEmLr9k4RF2by0v+vpn4YbDBMGpMJWLuSMlWcP
j21vXSmuoi+gCnLI5qhuzuTqE01MhBnmZtVwukGXYKxTttZbTjxgu/72i388XIirhnvDbyWPG3So
zqaqKXWvO26xxR/HIFYEs3yTgWZzz3XiN3MXHknAQ08TAnc8eavo+GPgU1pD2vRVFSJkzUTxSNEV
3aeLxiwgtuQ+V+RF9A58fl+LzG5n2Lvu351E2rRbUbJ2JAPUcjpgNttoyh6Dqux2ixSprgqtQ6p5
0d3FFRKDoUUcaEFK+t3JwU6hbeieY2Aphiz72zHLuZK6ZXcj73z7Jne+vrqUQXcUWUBqlplehj/I
dgigg0kMlT67pS9urI7wYCUO1/NBEfWt7iRc+t2wJAtHcjAQJLX7gy/A2FMcv3RoxpOUGGmyf90a
kxkk8vXaSot8i5vNweqEDVO9OpuQdU3g1wsye4jik34RQ70TqH8RQyDBwC+aRNZDUTpHN8kv49eu
7GZns4VIwcfD2C7htoZ2Vf1ANB85J5a0/6PIO5HRAXKqf7XEMwlPYpRsYqo9k23FYgIGdmmXCJAJ
WftMpnASU/kE5+iZYxmjK/ilWiPaRnqLMT96CSogZ/Ij+0tI1pxRIlcaswIz216YAQEbBRAjcY9J
ey3PRdn646Y4gt4xQ5ibHrCuWoeRn6qdS6fGFgu0EW5KwpiNVj0RTemFj7u3zam65XQkcfgAKPjB
BGSpaP39XkgPdm4yB9mGh0zYxzPvlYMNPH7tkk0232JoOVeuq7fnU/xNSS8rStYd7cElb97TNMKz
1p220Xxy2xVh11yp4ksFMENdvmxZ+GJ6jFuNfrPZEt87hdgTuA1/1wBSxHHSAiF6wvEn1XgpMejD
Vpxgk2wGopOr4EFBXSS0NH1godPjbk5WMi3cinpPEoynkWgXw5kP5A6+YVRr9oqIpXMc0bWCMQw3
Jg3IB6WeQ0kN5SV7zT5ursux3XkPUb++KTvschOYetvPQfr3JtCoibM7RzJ9MAVijWQB81X0xj3+
+8AMC25T6ZCJNXQ3zUPyKSA1MmMgKFClgbxl4T39Hb568P7piwP+0idRKrcYXmBx4ewLZWu9kJDg
KutHqFFolETtxRPNBxEubCYfpI5dyQd9oOJnESWQdmxUbu+j3y+tSKWc8kS46IgKdFr6L2lEaL0j
z42210sIkfoTveGDAC/kNOJwXX3HsKgyAhLEaRMMori7K1m6V3esoucE7cRIsrwhzG6HW5HLDKRn
dEd2C3wVb+p5i5IVBjFLgbsuQqT1l6YyTYcGkBRbI/EQLm+q/LRKmGNOa86s76wDj+uug9ZaQB+2
5xchlUKuHUc4Tg1WVJOvUdYy86rdwONMpqPISpu87v97Lj59964igBbHDIz1ipAnlkZsX+TsXseN
VHugARptmQJkrIknBNh4XzvZBaOKKIm9eqGofYRCqZ1kTGaFcSpvBcfAmRu7vHJLWKqn4bubkGXO
RpWwJBluR4n6CSeZKaGfPnI2YnZha0PUGvopgyLFxsx99nG1yqxa/MRZomIR+m0M8PA7Th4wySIL
CgOBS1sTRzmLqLjCzY4QyXRrRJievGBStHldz0ZSVPOTjmnG49nUz1acOhJfQJwigpz4uZcP70i3
oqCAo9XoMQlT4peTO0Tw4vIs5VB9sDg0Tyba2oCVVyGIGFsmXk/bapVv7Goil82IVAhpk6sdvZH3
38MaSVf0PEkevoRX7owSrcv/rkXSMFYhU2of62BbVkBRzQI3OIzQ84/CPiaaiESQFDxSLp3A5Nht
tKRAZsFaC8goC0N/5lqB+bwJziiF1UlTcAjMEHJqwiU4afVFo0imnVZG3cFxrwDMW/B6+etJiWqI
m+erTekaL16TCrYt1WpZp8J9XKqw6QqR4OrnoDNoN3x0RcjtKymYd32IFslWf+96FvjxmXW/okWM
HCfOx+yP6f4VHylPrOjxAlHZ3ND6OTlveOSDjJDVf6qI4DwJFGdEMIap8m3ZOEG53W+qLVDW2Vzo
8Car5HPLTMGYmmDS/45C1ytt9QbaUTHBlHxGdLS4y0iiuSPMjRBb2Nlm0l5bGfVHrUQq7WBKxLsE
kucoCAkbVw5d/pRCALdPyJ1SPEpKh/Gi7R5cAYaGxyOrrUMmv8HDCgxw2Ww3jMTUe1Vahwr2gmnM
wXLzdERnrognnaystjzR6wsPcjGfxA0U2BRhtf/4D+zsG5Uo4A3Xb2GvGxXHiTaMXJ+BhSDKHYJN
i5aSgtoJO2VWL5khCYxhaLxGr1fosx+3+Ev0X/bT4FeXAMwtAjM5guo9hVRnM3h/riLzz2bbW13K
IrAlAV5DNlbEBCri2vJZ683ZwqRozWuI0OUZUrWvOiKOd6HpZjGr18BxwJeg97Yd0SuNfvKS1/Sy
9z+uSABgcgWdnTuq3HzlancQw77ztjOxSrY/L3qPtrvS69mcAs1ZMrlE/m2XJM1wJP4irIUkGyRP
NKqVQm3NHSSWhHBhJNrlPOS9n0I2o3QGgDnOWNcNBQJJDb8ZlV+2vLrrJ7HTLXEjIQx5xBHLTtIw
0VP8lJus6u0xrfkYofKfzYevKYdaIb2iO4iWmEAeV6KJ8zkvhvuGdWxCn0uPY4h9rnmHtB8Fu6rA
aWBJIQWCORgsKX/38vwoPlwPC8FSL7gRAWsrMlFj5hBbEYF4J4llK7x3Sl6u//f85rCCng+zcIW7
LfNMqx+yyY/WnmBmBolm7trOXDUWqnxjW6QfbxRGq4BoIXJMLeq1gn3/GpX//6nMRTI/uoovEO9k
Fw7bTXjaNtUxNoa0XCxxIGOcFjB33vdvCVNUKl2//CCWxOE387CLck9oOVKycVeWIlGzw0jk28wl
/c4scgl7/PBgURN9ndp7HhvIUAzUy51acg+44gUj6FpsGI+3W5qNTqNBkyDwQzMgFpZBIGDgcskt
i+HlY3jGUjpEpunGNiwbyXjNNVBkBP19bmZJhcA2PcR92eD7GG7jG8Sq9LHPSwH0cAVJ6PpD4h9C
2jcsA8Xy46l1J/q9S4HnEEnrH86t86ZJ36UzyZvdkBHbnPx3ifi8Tq+y/p1Mx2reonLdRJcrT5W+
pZJoXv54vNZ5NvpYRzS2CkNnGfTYFnQNJJbGmOQm//ED1zXZRHyTp9dN6Neg6dWYTWldDB49dBk3
EWJKZDs81mpHVuMMVhyMcLTeEcuJe7ti9NLeyuLraQVHAvpNTdx8S9LQdeXVHYFZZX17Q6WlGnK8
6CuvsO15+U9tDdDzf13tM1wBinKp0Ygoi0jtaNb8AgpiioKODOclO2/DhitK3wCcpeVQ0M7NoqVo
9C3H1qc0NhWZknBuR5+SY3C4kJ8Hv2ZfUaqOlfoGplldOFs0r7cGG7JoR9eBxCOUgmvzew5wJvJV
5zANb6lE0mO2FV5gZJ8t5uUZQHF8zUWYY3LkaQxfKjVi2tTMKMIM9AC858NTZjGd5lTuAu/KXBhW
dgYLz23vJvQMMa09jpuvtiiNGDKPVkKkUVRBsu5vKK9GCJvP1WbnNii0XddoTkvI6XSTfd71LIfO
+HNObSrd5oQBDIfgtevM9DXiwqF2kBwAWZNsK/D29ptKJvMR3fqumQr/IhKzhgwEp+6hn7ESdl/g
BfHBWG8KEklqeNcPeiId0cwDow/jJZcOcjii+WOiOgJuAMvsItwKe+BNDP8Uby+9yp4UYvQkBAd6
g8b+WIvIizq5iLSoXz570lvFO1u7b4GMG5mojYanpQa9PWX7sWqkEakASp58LlChZHFSbEOqY84e
vbkkCovIhl6jl0RvYFaXQkdmvqHQuKU+QP+4mWwSJjN5nft9BDTslvgt5IY3fEKQ+afPmsUU4QQF
WryTBzv/YPXf8j2h1iCz8hF6NVBalmcgUGEWpJJNPr5x2WYd7r1P6q1N9+t25Oz6TmdTFf9t6AJO
WBmiSObaajX4xuPpntiJ/AQQaIrolXWao3COVVJd4L0Zfvtwxn5I0oYFA7vMucY5yChC3QI49P+O
yc/7S4G8gbR0g7BynTechRo+XRC4tEY0TDLZzN+f1INRx0dvmLjINezIW9tTMaB08BlqYUBsJgm6
KXzPuO2/shHOKyJNEpOYYvSX/lCRYyeYQpchpE6rJnxQHk8FqeKCQdX04EDgfhFu9XEYJ7SNnn8O
jpNB1vh93gFA5dmbRL2rMUCns0d2afIqeJrHIghSbajvAddNZ3RVSyqCGOGMQczQD6BMq0+DZ1s4
BivJnMv+RH1fcBkeXaujYreQ3oDSfyzZcvMttDlc/FQ+K/myST55bmqX8vKl96Fx3t/1llRs/c32
zo+5KJMGbB1OZCWbOJWzxnKFJXNLwsfzRHrT8xv1V6JNHOjdzg0fFh36RtmKkpskMMcyvHZBpFGU
1/x5Tgro3uiqcU8wkSJRNUtZpu8VBhJcCWmX3waPWfd5S7XufssWG4xzn68AZ94bz3Qh6CNKIUNc
b2TcJqfvosegoGWjR4pdGLXrRFvZXFIPIkFKaUSeCJPHJ0NogV/iXz5GYiv/Nx1uW/2eR4Gb5b+2
h30F6gIl1DYTDob2lsm5JCcSX+ghMOin4rwOY8dGuJrwxeLeXUwYmWBKjEzQ4I/vKOybc4VZEJDX
O7uTRFKsO7HA7l6vt/GrNBVKaWz/UZ3x3eTaGYd70yjnchMu12/QPJz/rAmbJmUfBdssOIuY6VkK
R+VOef+Ux+rxrvVfPwuBkRmng4J3GdK+Vzepp7OtxfYpJ5KHZVU5MeMkSyfg+5GBVgA3or5+PeeR
r5/fAnpolBXY2U72qVk9xwtdF1s0u3SYG0u4LleHVjBkaqXbQjF5oR9ShclOv7aqpmFuqdUmBXOh
U22veoliGjK6rPJIU0Uz/B9a1Eka/KOTYtjSYfIHlsnvy8kDZViX94MaFEgqI5egYXbpgkm5U0yS
97i4dKjqMzLaJ0vEEmdRcupsTYy9UaKTyDNaBXj75Xuocm6JMoSFx5g/nHmcNyEejcM/hdjSkQUJ
k4rT2Wrq95aELXQhVQx3MOTMSCbAyUPL2KJAg5P221T+wPJ46lyy3YUUn6irflts7LqnphC2t9q2
WR5GHN3bUSFVTnbzXl/SXMbqOlIaDExFJSUStR46I3xozyobSGl+GLzd68h2OHoaOxdMO2cVFFVT
rdAsOnSmGSvxB8pey+bZDvvSvzjmea3FkIDdHKfQ/3pjza10HLUrLh++wkRQbdv0Z9YGZZzV5qmz
B/7pIRkpZUKdxKZUkwlWUHJAvZc8fkd9gOAQLCjnBtznHxN9pycSS4WMdi8NThkFHcE2EQUHKtY/
PKVEABxnkH2KupCvCX/CA9tBu/OMr+s0HeyYUPyC2XSUbNZC3Ag7wDPuysy2aSqMyvAfNF/QXn+U
VRdYjaCRena1ca5wYUwBrX7XGnPkTdAvrG2BkacZMPDqPuFTHWiLzAGlc+BQ3TALrdw8bY7jeWb/
JgXqAwwLsXOPLyY1TRWVuOAIzwgocT8LryjsuVe8aMXZIIBdYgLWXeZ9E2kntSwhs0Vz12Kh428Y
+Dgquxckg1OIOPvI7AiC7ZgN6kMtUoumKPIxPXEJnucCbA1X3pSyx44yURP8JBPtksyTLZgSGA7U
9UQGCvKtynkgHpYkJWT7t5qAM/7rMsfP2gmP7TXkKX6w3dIS9KFbUwpw1DweVNEDFBus3xwMUcaY
eSUIxYdWhdU6FnpPwkZrA2mpbDvWX7Dfk2BBCPE72DfUJ/E1glI+rMLW3UrWOwlxZvqaj7bWqCzq
eHBf1yajUhgPwLKWDGaCn2R/4fTvHOF4GPOdnWBlzcQU45BDEXGUZ8lIEzKp/UPUY0QaMpoljoSq
2SC3+yRv9a3Ibma/EnXccdQuYkyVtesySxsmr6uWkcuWlb/hWn63/PHWhZKfrD07AqSEEgBaCcsi
pyEDow/u9xMsLEPyQaU+mDDzrGhCgCoiHXDlK1u49gpvli4Ez5XDKKNjy3oMfRMpCPanCXaWR8OQ
wmg+iAsxnGU4tm9qFhdhoNOqPyLcwOFDt6N4Km7k/lMxFL/tpKLgevM3ebE8ZzCdMV6hq4A5BEn5
X28Ck6VDsKMWMbPTopWPSd6esvFqMnHLtaWfmo29L0cKftYsiy6U8BLEa07meSz7lfMWlmn7H2Dq
snas2c+cukRRC2fEasK8NGODRYxMGAIlyM+s2Es+FTjUxfcDYv6aP0Y3ySRac307TsjZB+mYThBS
LXXL+3k6XsoJqIzVRLF7r3+VXYfhbHTIajBCXVDz8anDEiNRQZ+RS/DD9WkvJkIFiIjMSWdIl/SA
DOm56nrXe2uBXCKOaGZRMW0N0cOVrYU1UdNkt5T/MqLwW4aOwIhWhNi5fkXdsNIVnuREac7ASlfL
E8OvZPwBhuz2Yv9DlEAJGYWhA0AYJoYvMlE0a+30/mSu0QQNKAGJXNiUp0xY9/j4vEwUapXh4du9
xMLHco1tUXTq1OTdj8SQ1L0Y3WaRvEsXpILMGg1iTUAUiUlphF4w4mMnY8mpPq8r1Yj2NlnGVpLB
apNyLJTHLiCYEH0QH+3QCzcVY25OGMFsLC40xUOcbuAHmU9ZfdD/gNjiHv5784149XrekHo2vmpg
3fy4+B3LjOitujGvW07kIBPMmbnoUOgqFq+85gXpKkVvQ89E5VABRCSPq0plN2uvfS+SXt6I3W/T
iXlZuFsSMnakCXbyjg37qYdBj1UxunqcL5fRUdqyaSHOR2jIBs66P/QU3g8OpxQqZCOMJpTjpMLO
FbOLSea9iwwHKQzHGpTPJUYJEJRCInpgkAOhiujp/kbV81jJcWihKBKb6cJ8fu87mJ0/l6bEqrUY
QvWfWMw4c1PdKIJ4KBHDKBGHVPvvTS0vpi/WE5DnteKEdSbYI8A/ActR5TkuS3lt85fl1hpCzLNt
Kp1ajvLos+uRx3in7O+I22sRxdroF4EYvNg9ueSLct3KoSbslSGRbeFKPLY3ZQgvaflR1mAi614S
BODDIsl+2adC/3Y36uQ0nB5HhzrM1o155lmrS5jpCPDD9ZXb6iukBUp62cnGnLqMm8TM/ik7b8i5
cSDVfbRBnmHbL1PBuoiCd80oU/5bjXTVTUhaq8LvzCwINgG0Rq6PvtEu7LfcnnKaXvwK9Q+1E1qw
m7n9+zIepREMjADZhKiwiW1dPhgwyK7So8LwgboPjvs3JFCGIm3kpC0wts45CLbncFDreQhNySgV
h8Gu9FhfKsdb1YdM6Gij4ZXx+zOHxTVoCP5kKxZSwsl1frtLQkAZ58ea2Fu6mrB5Fc7R7cTRHu/+
nBXU9fFccfU9tnICkYY2bVWCmE8oW8vH09QWkE3s4b7H0UKwNifsxsvVdOJBp8wM7ye8U/zKgS/0
yPoMa8USsN3VxbZuCnIJYJHjd2G9+67Qy+mpAZMTcAL5ksqOFRP6+T5Idy1EA2U17MWAdCTfWJ8I
bBFTqITAVuRmjWASjmauqy2RsGCxkpOITFn/FEMorF03eA2OIPhgBr43owjgWa790H4eInxpYlX2
QiFPu36rgqWHk1duOgCBgrJFUoSo5jx1I1cqOVTNsD0fLeKi2VgoAyLuVFCVymvIRSAroPzqwgqO
1NHokZ91BdnrkfT77aPdVZg6MwkpmOTFjQiWyUvofu6kZyhjsGEUOpgjLboqxPsS7cwwnQUZ14z5
j2oQ6fiBbcI7j3Eihz5KRFF1SDAUEYeptfmkRpfEkHB7MJsZtdL83V62VU8oQkBRwLk2xo+WRd4Q
tuJyi/HJ2pJtxrRdtjBXR8S7iEcL8+TyLOU9VBm5PpGvmXZp1RF2f1d2JqPFB7pVT4I6EjYsnZsB
gqb/YxandbNpMhAs9AOsbm3/W6uNk1wTw9z3tcjOSoVIKedmAPxoEOKr7w4Aflo1h4hh7Ra8xaB6
Y7FxxMjzieW6fXrr9qVYeHPbbgyKYSsaQgBwLQL4LwxCZyVzCfRk1HhJyRx9HQmCxBT6OZX/iFLz
ncaIQOqH9divUWz2Dt5d+cgBGlJ8eVoRhysWGaBcwYCRXUAR2OfXPvYN8Rk8zPw95jvakqhX87aU
66J0ZjU3A0V1IcNqCHT9lknoeuKLDaLWP0/wr1uFFoOTBn19t4I+rHDrzYbRo2F1ZIcSNvq5LW+1
wVwT84AfriBMC51M3fXby/hwvs8a/D8DpBLXjw+bIkcXPIbfclCMhCiKxLtNEwKPwr+qi3N1Uey7
DYR5340FS4GfNbiWz/nB5U6VGQnWzkeFN0JhUUiOl9vhOY7TK+rsuiFUXVUKbLUmXqZ87X3822xq
jKnRJGjvZteloch1qppSsFANAcNqPt+TeQ47p90sg/8J/vAybBOz1/MdFlw2rc05kgRjIpHU37l5
jI5cKDcIY+g76+W6DCgCNxeTtgBU2W+8ckbYWaj6rHgohAGVt3qOwWyl+q4c4fRNyoXULiw43KNm
AYXITdsCf9RnFQsdy+NQT5cS53nHYwYXG7MPfwDWEo4zVK+eZOuOOXiWFmShn0qYqLYXESn+mNnV
PFlwxzSdc5LCgGtisR6wnmiJxtvZMJ49c/XItUXBrVQDRdt4hfEii5MccCj0rEf6dZ+lY/O8Hg6j
O20MdGuC8FpKC7nybdihbI6hIzCX2Kq+ierrTYNfS3QaXs5bGzGSpcHTCj+cM1S0nJBhNh1G36QK
ot23YcBKintt0JpnaAfKbSVSJYtCNLi1uMpIZlg4WSDfQNRzfzVjrge80LRH0KeM2wPY0oJHWmNL
oCWkmZt9k3QqkSUyp8evaDovZlfzwbLGw0ITwylMwsmdngG2vzPfqfsiBvfPsHlOaF/IPxDmUr6C
W8IrPsfE/P1HxxIHKJnO36C0y6cYlR3jhJitC8DMtJzOIOVf7zX+dM0UPr5j2v7rokdUiwAtYuGg
18okrHlfe5309HuV0Q8xIlDnduY/R5zOOeFHb/A7ToCWS0pmwFfa1nuqtmITNx+wUq02L2d0DPDm
Bvsk1aX+VYJVNFZA49lMzn2C8OxOAeHU8+JCE5gfQSIugbOMe/IATWTXq57eZmeR3CkmMKYq77fm
ekE+vn+fbuRan3pscMa/zMAxo61xug067N7ERYPvcaPJk8MrgoyXNT09fSgXmqmC10tkeis34zyW
xsbqoCuBhY8scpfgnMtHx7/0lkVpxBkJ3Wqv93XVt8S10eKjSi74fIigkZ07Qwq23rKXG7E0D4Uc
x2koE4uIMIT8tVTjOjtudQOArg6NnR/5H7+11Y/al2b/UrxCI9XmEOwEulHRPOqkCTdUctJS1Ijn
E528cm290X9jnbkdVKusywSSh1zMYrUmR7SGrQRRzDxrKyZ3cPq0+QbzVPfJUk8hDJyN+1BT6bKg
2bMH1xjKxzoj5BN7g6NSTjykZzFtLEQ1QzgeQ2JRBVwKsgSekqxH5nP5mvxOXhD0eF1H2G/Qkpzx
4lyPV0Gy3qRSmeyjLMYC8TYzg+sl46G6vtFd2hzK3sxDD6wvc+BDVynvHdy+HsAnSFLnrLqq1p7J
cpEqwc5QkaaKKLxW7yLwAgxb4iHQFEA0cSsJMnP3xPCnBcdJRhUfQbDgghdFI/BKoIT3rDBcunEA
d4KM+h1Nmwlg5NwitReu+0tkPeF51t/ZUXxD3pRbwXAt01zXkZqPQagd3ZuJdx04YJApEMiqbYR8
by7eehoF02UdTuESC8nlKU7wu30DZE13+XuCQdG6VZKMbwZNxpURrx/uJQ9tj/lW+CFuMTyuevzo
7rPNgehRoXhgIoyhehAVKjxEo8O5cBo1bIiiMoE6W/0EiPL7LttWSyQ9gldsinFZVDuhmU+P1Zr9
gQP/FeCNoII6zVZzBc4kHjN6E8LNg4ISzViFAIinRcr7eNsRHXm3x35Vfxj4FWAJer3oZQ5k+G4p
LbzxS1aYts4X8Vmo85adeywh83JrQ48M5D5CyGanwAtwkHAwhLOKeCl/x2CVZRrByqJaqEyxZXjM
VqsbdbvV0hdrq5TwhP5u28NjnLYmQJ7TCiLbpTIaJOy41PWiEwOsChlk2Dh6RnWLTooTwQGzGLr+
vUMktqhfkobrqTTbRz+3PfEtMPIyzMgRR9Os1pfbS5CGZcs/xhXfBp1IeV8NeeJCpqxytVTbdyjm
mgSBklfZmthDCck4Q4gBmdPK+pKb7BneEOYziB9KpIbyw3uTrD4s76R8CSrrATQZMnwNOryVFTvc
Y+QGpElg5K4EwotEH3L+g+QdizurlmSgEKuEf1Dg7PWD1HoOLzHfgKcJvWiSNmcGOd9sXxOIrSs/
aT/BBX7udR5Bdt90r8uLZ5TFQm1zJRskcNDFFfJCdsvtwMtTnGrQ86EyKm+2kAAZz7VFhISAi3EU
xCCsBci78Lj3X8WRUTghP+8Ev5s0YgJomzXJkr3qIvmAPhew1xo8LI8oz7qmMxzCPF4LprDY62Vz
2J7IRjCBEZH290CapMV1M/ZZKXxnD9qV7oQABYYkhM5gJGNa6ZQew5lX5u0FhoijmPO8zccAMNMz
jsa7kD4AzF/ZuWApeqs8bzkHgWe5WcW9k8XgaIu61BrycIT47Nq37QMwapKQLKDN6ORC40MsI1K9
BsH7VZgMh8dNm3hKy/X0xDArLTsjyqa78bcWV+6HS2CEmndylJczAGJutSoDa1sdEz30rXt6KD3D
xK+bzHdALW/Z9kYXpIDrKQmav924KRMQzVLvYZ+T90ZopI0rk67mGMxyFY1EtqTz+AQHVe0ND/yT
WRoQqj9/6vKkwZ+KVFW0gXmm0C+dCCNitOz3I21qPlNsjM8w6tmsZxAsXi/M7phC5qbixUjPI/ao
qjT1/hQuYA5iKUlsMN+jOS0I+t0Fv1SSV5+WYTPvQsmc5qvfjXInXiRyBzJr2GNaAfVHXW4fQwQw
cO1ugiC/m9CgCqT6+CqV7a7o1zoLQ0PzlIt0+u4t9HUH4lx237h3dWmJe/6mpwfk3Qltd1i4Cas6
lehnAGKXHGg2veNDrRSpYWzdpsCJ2JOoBfeJzTTyIfX5bihc/rM1yIEaERNNjDQYZMhpwilVSIEY
oEJ1ERpOnAQh/XWGvUzB0j6MvDbErHQHhbNfePJ9ioxJ6OCQQzn3XH3/CCwmbAMwHNmQCiMu3LVt
eTTFqAMb0Yw7PdV2154uxjWLdbU8geF1adZY00o8Uy3HAmXssNfobVNaWCBRK2oq1sdeTls+eMkb
hIATDF2mpHXJ+4kMLh1N0tR+YrnCTV9tXyq2OLdkjur75fDMQgpgTRhkzHw1UKQ/CE90CvVi27RT
9+rx5ZTKdago9XbnubrXz0A8Mc8RRKsMcKcYFeP+zvCufPjiUZNQR6FvgcPXXUrpkGT41DyaZ6FH
1+DF/tKdh1f2OQCW27+gmDBrfZVhGEz8yfFn+IeL6ZOq6w2ADmSn5bpJK6iWrRZ/ZOqGKoi7fXO1
itDlMFa1QIYl8zn5YUcdrejrkmebFl7f/xrsX5MBkYopnKBAEJynD8nVzgKNsT86wN3OdiLJmiz/
2e94+g8ipZr5XGbby4hMzgJBUbXzYUScG/2NBVhSO7eV4i2cvQJonVRtSGlq34dGouWZ++IChc0e
FkOAxU7W2QqV0J1s7F4Vh0x0lASVkBv8CBx8dKz/3BDEtKZv/vJL/qffFm7hq/RQL3kJACXICjpF
dDNiv20ez0W5HqeKO0hxsoZwxdfx5+yvzy3fmy8TB2Qj4TkERapt6Nd4/hzA0197CZSkqoNfQU54
lFn2qWHCFcr+1o00OFPLYJnKSpqQVz82hIQzXe6+iTldxSRUAlHcLOAYKQBQVM/c+pbkWCuZQYJv
knkNmvnUFzAZ3U8WcD2lzotWvmnQp1kGZzjtVvtMYWsGFPoXfCceA8RvXY6ESiBQh5sg77yiIu/f
yvfpIAsbIzWL8tHdqCvVdDNGKB5JHIHqFD6c9hL89f+jAJ6X8xgqWlQurkRKcBLYraO6g8itHgME
lbH+ItA04UsT5cXZEnvwtYZb2DkJlT87upRiMFEGiZ/VdyOX+BY7qckI7iz4H9OFUfRE2vcOlQuF
iryjyBoNsJGmqSlIORleUYedRvdI+SorszybE2C7TMEYAzsrJaRpwRgwk/dcXQKx1mKfnx2Qfvtd
7YXZ2CGUtBlnK2AeQCSQsn1Zobbsa5Mfiba/ecvgp7ryT9bv8c1wLbYQOt7P2ZzNu00N1thnwtXQ
3qThVIixJq0hNoWgVhBWN+Py6TX5w3PQXPNZRDE3i34RPqNpd4sM3v7dVNRfkFbxqomJjVo7r2sS
tCFebQmw76F5pbPZBEpHr2npfiXXLEIYaro0wIV3JOw7aMGCGJpA0rF8Vy8Xm+Og3Z3VNxVFGkLV
ozgZzFsQxUW2/Z0HgNwQkPnG1w4Km7a4uybiWbXh5C53BWf4emZzYHGSK0synfNWRSvWWhqKeclD
OhAHdMTNcxRhpM8vmnppB79suhBTc3UxDLsCP435LjEABK0D9Zcl1uy7YRzyLJg56gKWBCcURBZ+
258jyeogvQ7KZo1ixsKVZrwRHUgMmeNL4xfWQu2vy1ZMM0CDLll297ZHecQMfwdb7hM3Dl+Du2xu
UBmxBhnQgJWS28C6xvnUzcImD4bec8syMSaDZM0LyYkWOVesNnya40I9bDqoc+kItN/V6Z5oxg7q
hjMjtdASCk1p+Yv8GlY+iVrZeFkuiVfIcm7KeOvW3TLIf3ylzwQWTJIQj/al0F8toM4J5bNAXhMi
Tc8tYzqaHUiZOQSo2/OYY+kgCWsmzalPmj/emKtnM6JZmjHe4hmwlDHiKDD5xwlyhHmSFooi5D/2
JyRVzzf9Hfas4ad+SZz+47CLni1mfIlSiomEk+7m/23tNfW++bbCJ+DTg1mEQIDLHgLPjbvb4g6a
T3WeaThq8eIseePUiLl/FXz4QsjrSxUZJnXmtlW+60GEXp0lCtsr5UV8Abazkq/5pgr4KrhjwTwj
J/bde5DlUJlE8DXzI+b9gGYd0e7fjBATlsi3ZPrngkL9nB2bjLYGUbrOcpd36lXlvMyy/M8vwfll
RWUVpYOpyEyliksRKSDuMQma79CrWtK+xw2YNhvn8bWI8ORNgTqaQ+LJWUmIIRuFE37y4w8WBKX6
TKyYLvtpNReJC//6EtxCiJXHuwbwFBHpg7alvluKX1Z9lIDYfF2N/KQJjQrvEN8OXP3c2t0qsYjb
mGyrSZUDyC4cn3WYKY4OFDR99fa+rMwieWSeU70kpSzQ4PHnfBnkHUSLmA0fNSEa0Urk4becoUTU
isBXzATfJUUH5SthhXmlfm4mlYUBmeA7goBVubZlm2ztbphVyVroKVnBWZfsmyJqCcXUPKxWTxEr
CFKHSOJbBt84b+fG+j3T7WkcI4Wsk1ppo/oGuN7CaqtvgG7CH5i+9I9PWgDETlqcihqSycYUrIEX
Cytdyz7l1g6mF0CgwHtZe5PjupR/RvN2Ddk/6xlTFNmJ0I0PxzMu1IjovT2Dlp7uFyOjCZ4PxDob
g7+SJBuBNw0/kK8NacjqXrN3ZUOZAW0xQEfW7YjpKKZudl/obRzEioOPRIXesD8QBQDf/w4Y/J0S
Ka4DRmIfLMQfccmcGWRnU3EMI6bH7ftQ7gFs50aHhY9b5dEfV+Y260i4jM+10Os//rd4Ul8ScBZo
ZVLSKHlSnygPV30xoZHb7PrA8r7kQgatmarJbpBm3hmdfY+IU8fn2qCwQx/zx+5zv51vtdTUCYCq
g2Z8dsOdbh36RZ/OqVvWdKuKjwKWY+ybnwCHYEcNNMaqIQzBILmViLpmX7Kfj/N7OjT3umWnEGyy
8lLaP2iBy0Vdn3V7+hb3lVbDGCEeOXqsZcHRohFtpGYHKm2Vapc6LlXIpB6aHUHvY97R2eh+w0aZ
Muq5XSP5GGvooFli0a1nxQyJnLUtLMxUVEKIbwb70SqagPNkFus3HXpVZwyziUIqFwgqkA0C6vo8
nrdB8B8UlCbrGGwhewIPEifOIp7QyfcvNTp2fB1Dmms9gEpdxFWDnMa99D1A9rcgz6DptaJx00ne
xVehrYCHIU4TXUHEuBuf5xow9inbLvjVh87hUteRm9KDlerTs5/0/NT114fZN234Hn23FrZlcz3y
6qPpdOm2pddrzFWgzi+onFEdMlf9eB+AOrvDdphUFAwiZxh0FvWsEfMk1MTE9ryZi8mdCixwoU2j
Hh+QQA5EbB/hWZmEisCxSIZxN22kKqC2ziydZDAtLXz/mlAiVDCornCVzBVxG+Fx0qEWCXmEJtXq
kKO1yepZCb4cNw666j8EvqibBRMr169EGUQS2tffLP3UUs+mQgzXWw6W7omnEaMAkPCDys1gTtq+
jZp1R7Q5Gz5TY0xUBDGJRAABZsMkJ0/+UQqNiSIvkYrRtXTikxY9v8f0lwAgpaHe5BMITTOWFp0M
G3gn0BzhrLQ2GanQxHeI64iXZmClnvlvdmqmNY9hedtgHNlUVPRapCrqQRAC2BsRPtb/U2flbBwm
Q/Bl+YRZdhmpA8uY746YHCoCMNcLYbO9GwWyQSWZRcXPkALQr0H1M8AE0xjDBlLuEC5TaZiirUOa
eLIi+5AH7392SB8q2aVv5yxSFsrAv8VauMj10IiZDS+AZXVTMvOaDTlxDZb15mapeYdfQcGsr1Z3
I2sk3AXxJ//uf4cChiqW9Xavb5q173VIM7jBYVJ54H6BKB+xCle6x3x0BLZ1m9Sk+bJ22BpWRtKU
+jzmA2na3Q+HaSYTFPaDzrF1oBq97t/+/vWVl9rtVVXMey+JYCg2YHE+5VrPLlyh04i1UPGKyO7i
G1DI5J3OmNITEUAL33Y3eSbphyHg0O+QHcOsR+QmYh9n9Y/IecrfzMhcnBcU/cwD/stcD201v3dN
k6fN2ApGdgdlB7CZN4/UhzJApjpA6C1ZC4CkagrcdVx8V1CuL5V1U3drLPSkoPM5iwbFChXYW/MI
PLE58qDiFIW5bqmGAGBKtJTZJIWzOadbSdOgG5iBEO8sfB58AiBTi80Bm7Fvorc1obbavCIzRMtU
xHSbjSGnD7wqUese+HACs7oLsYpB53sFllIUI1CbG1Kxj6jP0zic4LbEdoR1LiNtEJTpmN80hgYk
saVlLsjPaIARTc4EHjpSi3eJMrwEhaiCHzRSlyI0wtYA/pm5wkqjobwo1F9Iktub2rgxkqcziJ5g
j/Z9biMIyXD6DHJc82l/JZGofDqxXk8NkDksDTjKHlIdgZPX1W2CDA14MQNQFWBkWs1p9lrUaKVA
fssIS13XgIZlx/QkfjaFgOqiCVbTH/st0l/vzvb/jkNC89FKlu5DP0TBNfsB9Ta3ivwFT7ojTwRX
XWCMAtSZ07sQgvLtOB+nOcaSuTm4IJd6utkbNXV3DhkT8k4QL3FFWx+D9bOTmh+eqvoID+paXS0/
20TQAS/9YoKgPe3A6TN3cVXMwvoUYOlUlv8PaVuKMomHw9GHHtdif16PJ2VHMPqbz1BohpNBqe4+
Kbicz3X69aRlQ0FjU448W5xqy7ibNEka6xKHLMF36Q6rDKqq6ZRv9wTTCv0f7RVpXWHVoXJWCsQ8
oRxgn0c6SGYb4o+wJsQR6/AzZeHg1DPdq6/piFXesDo2y9K+FCY1ixud5OH2nFgyIWyChmwY+uD3
eP35AyYEG+pObDaD/0MsdHjAhzq5koHsy56kBHu1h7J4jZRQciF5fbDZc3MYx+FGnAHLKdv/VZ8V
IcGl6CmNfmPRcA9Fmh5SK6Tb/ZI0Qw3QhaCVC4hAbfCwmCTAhUvIgKWf3MIFCo1AdlUbUNA+JE2r
IoiD37u67qfr9/2hOY9dX4rgaeKWpwVdEAdiPQAe/ceQ7ybuQtaW3p9EaLE2DFbPJrhi8JCLWfh2
oIpLdrTTYqG8mfRmrQW8vfEM2xQ+XGCsnRLPqrjPsFWXF2QYmDIAqFKRTwR/HT4HcmT/lj1td8O2
n6OsJ4bbWPJk5clgtkDsay6zgkfU7QsqbAvppxYyWrzpRIMgjdTmaoxppEaXfjSY2TP3zJ7AO2bG
G3G2/NVMl6iPAityFsaHxK89lJfZgZEE9Ij0DcGl4WOUkiEgpAEKccebb54qHZVemPm6OILWMclK
X9otOCtYfXePs4tK1SGtX610wEYTT10epgYOtzM2mxR1sMWtu1GCzhAk425D6d05iS0plR7v9qA0
ngOcflibJbzrQAjtrM8j5MuX2OGheVpgavPFRxcQiohsP+Xen6gyd2/NiwgL8n9SjEkSbcqJW+Rp
YuH0LtY7Wq/lncP6NPopJ+4ja/75IJVEH4+ccWW/FV2e1IbKr8MqBQsGNQ8UkPbiGA84vumyQm7Q
E41wVWeuIUv3ruudafzm2YlZVliEagZK06gDU5L5OQRae/ZfHuPpJgAf7t4+IPFoVvxiJs6uoWjT
p6Ur957YzPZ4lZvXj+0QFK+DJ64mPqwvdc8QeM96ItG+ql0Nos23Y4xpO2GE3/DObGvTPJI6Ezgj
ud4GPB+DwYP/RRjCRuDloMDfKCQqFwxUfiyMiXAdioGyPW+6r8rp87bvXD8gcUI/74YzJtWNTbZa
qfjwsP8b9LcCBpNfByZf28uMt1nPSFawSHAlm8NAngZVFrwJDeCxvc8RR8GjvTaf8IcGDBizBvU1
PwJjiUqwZluQZfHefEfKUWU5HaV5ZISn1RbP2oom5p0A7r6ajsFKRcOJUES3KGVi5xwtQJas0qhc
0tQCbDEoXxlGASzRwPUZ8gV48WBGWXUxs9MvdSk3hoPEJiFMrgZQ1xM3LhohFjL81yC0/T0ojwgs
LSY+d3setEayuYGboil3+IJPQ7NIBm/wVyOnFw+sxLJDsg6VilZSAGUPOxuq94hQOeY+Xqh/UtxU
KGZrqkbP7fIWXhgWaYP+Y3Norud/+nr87VdD+8wubWnG6TApw/5kjdj6+OmPu7yJcuywzy3mo38a
6iMbKiLqnFbh7H3SXu8y0pOeZIMwvVBEQzV4aY9OU6qbfkjQtj3QcTMXOF3navfhbReBmc5wZuXc
iXfn3JInoXsa7hY12CYIL6AF9j8GA3IpLmjrde+3OVKT/T72hA1OeCFU8N+SffCyFbTkp49UwKfW
i5eb1QO7Sk+N82uUOMR1MzgDyC1FpUcB5tOsOgKJIs5pw+FIjHDncTHE83AW5zwmsKMmkFGSqrRA
gZEDx/QICyyjCFe7V6ePLU0syMsw5hFFgED7xZJVTLwWsYmTyv+Hn1OnGTVd0Sb3ZOZbzbKrRb/y
4HjIvW71rhC6lTTWCSxbsoTXtiGgge5UpCSYCMwe0J1iwYqJyqcBwcG3Hfir9PYj3w9v17XGsXmy
JgLZoSeUYaR7BK1qSdgoHwtWMI/V/7d2D9jrzP483zbyPL9kNd9dKHTcL+ksy3xvbWyxWysw+4hT
JDUrKelfUlbrVnxNm28ng32vDle2svgI8qIp8VNqQDlhsm1F8YPtD/P9tHVG7QxkavbtyF8p4Gd3
DMuvHljne2VLpF4nq1/yqyC3uOClqQFCe4iwzsFdD3Pvx1jgbRP8MMMefw+6nsg98AaM7Tb2vE2n
HvNnAinR9p5eJsnxWGbv16xcKmkwixzReClhTfeL26bGNDSQKxjFrp3J7nFw/ZHHcMkAsBwvIKPi
ws3vUiNhbyh+7ZHqPr4YFaJyKPJUBQ34Q10D1B3qVP7rC6Tp05gGfFasNgy5ma3wLVCFsQ7IWLaq
ZnUgL0Y6p6ELll6HhYkr/HYh4yR0PLW6PnXrRr7iuCc1l9xnQG5j14C7ftLFjwzNDVZ+8Ak4wu1t
QsRhqi5P5mRHbQCz9HGaF6i3Qn1ErSBLngNJRLLS+MACmq3U1YoV80PpIJ+mfxBbSvMDR0fhoC/u
GSbG2oZcsdGDSQmrZqr7JlxbKVFo9tTmo7ipAgtUuiquiz3xkV4DDJVoG1Q6t79UoYer3VZeYDjQ
8G0EZuudzutpNxwytppSy0TAuB81ie9MkC1qROlSiXImXrGWiIzy3gYfs2qmatG2FegBSrScXnqO
WbSFg6FlYP5JjaA/xq9+Jw9Ij7rO3GHXiaQLtG7j4qsMyeOtIO2j13pOQoewPVe8vvYpdtl1Jm3K
6hRG6heMJYU8TwOxJWTRoLH1wKlOQXMLZUITrncdzv3OpdyTTt3UNUzb0X52OjvX/vdrvo42Gy1C
l1HiSZWnV6yJHAgxtjGAL7YaYU6wPE7Qn0atL0FTLWlZCOmFfH++0ihU4k3Nrtv/DSn9oOdd+QCr
LJyI8WRTg1SzKzV5UWpfJ4I4GqubuT+vVbk9pT0BJ8iA6/2m+bmATW4dcBmGVbgtBYIvjA6ZjbAC
kdJ1esrxi9UqNrA90FabV9GoC5u0/Bxn7Mk6Aa0L/CQJhRy+rApprF2k1tVaR1PiVi1VzGdJ682z
n99PaGgGN/aPV7R56T2e/17tDCrl18At+c+Y4BVH4Jw2pDVlk9ATpUqRYgch2lqMq0bBx+kiPIuL
S4uKi6fPTAMgAPlDvEeAa7vLO6rr/nO1BP4G62PKqpyvKnyRmCeKuY6wRAesTyhCKMVvVTpvaOJ4
UVjWNBD0ue2vcWrjgsDCQRnkmOS5QOE+FM/X/fj2RAi2t2aVwNMYUAlhh7pFQvdMqQYV/5WU9eel
9XLpzpyQiZ7ASeoGDqi7Hhg1PJRfCq3g+YQ94OyVVpM+PY/++Zm2lYxDjJZ63oPX9jfREPNuyLU5
N8LjvGjLFY/NxelVppBW7J8BxqZmUth5g38P27spD/+u903rI0eFsDrWF3BqMOs7koeppkTJwG8Q
mZ3wDynpqXxuzOJjnj9Zh9wcHrboe8T6IeDwNzdlJw8GSbcc41t71Zvq/eOjCDu4jy0oLFYmCD8p
/e9MbbYguuEsK5cuBmLSzCgEUvVScoJ8JvanKMpYPgZyx62B+WRGXKpnWMeYp0XNlNwD4ymd4r4n
fi2RnZhIfuEmhHYXRVW1krp6Ceagg9eHXDRtDbRFFDU3GxY9KwLlTdnBH2HYivUYJJMvhDY8tlNH
k6xsLzFvRVBNL8b9t/5S4lZS2Ha555QKsK1rxroC5Lsas7nkJvLGNYp8wLD5ug6mDe52dznV+KKU
cyLwACmz1XibsbRs9TEcD3cRR6GumdJXtv8/m7uZaUo7D2iVOYQ7TeNSo9T4png+/CYBlFKVwe5x
dP5nFNJFFug+WJeV5r2qKLKfUbU0e2MzlUj7nfv+QwmsYg7kl5cJxLyczXDDH0TIRCOdgtUsEc5U
rybP1YBNluoDdN0Man1ErkvMH04ghgCGlkHYLvV/8uYFei/t10QzA4g+BTW2vWEH9HpYhWt0tZNI
7JVTAq3bfWo16iFeMYkbEVNAcJjrGOsoGSqXHyVCMqalGbwsDicDvZ1rK8nez901Xqywx8pJW1Le
1Jh9Kj+LqF86nctr1U04ZodTqAO3HmJDyHDinnAyq16utGufrJ00Cs9AUXZHDIEjJ0R7Pt1lW2GM
nXTqgGm6f+deJVzuMrEdAJ0itewRHQasHxRJzV1mX9dNNfNcUzXcZutM/7zOloPlNstjQr5Al6/I
uq6EC6WaLhAqdT7fhvoC1Ad+rRpsVbObncvJ6ExYvP3StAbaRSY7K5eITfIlMAUJVQi3+NugQ0uS
43YWOUGOpmMdrJ8DNEwgXhbkP6UPja7Y3boKDCo2jlcgnw/4v9AFv6WAMuRlEViaJx8a7blv8Fff
GA5kkmMBTEcPh+Cr1nA/xF5H+SwoHGZklGhgzA1fA72x740Z3DbDaKQRJ8TvFoB8LdnJC6EVhjsa
vu039KLxZQkjzbDmXkyNzlu+OcU2kt6PLMg86SgiEv8WZpOR1Vkd00EqBRpJ23cuwf7WjiujtKd2
iqTrJ5pf7nxtKQfgYLwIZnVKCrUATW69xdxK869+6hGmPkjevEJm2D04v5SndkkFCm9t0mdWpOme
xL8QjZWn1GmpNvNSnT6Q7e7kxQZ4Ww6jFmftoHxuAeYQ+uI3N4615W+kCczs1vZr3QDEo7GHE+pQ
BIWmzEPl7EyI0mSXxBJnjF4rxxyr4mwUPNKWCQA19lgj6F0c3uL2nSANwzyg4IEakfDZflhgMWkY
BBT/N6zxGN65fS9amxJQrqKGdnkyx0PWNYG54B2eX/+9RmZEnyYlCty8T+ibl5mioTcrSd1KmtRK
sMjmMbdYDogcnPAeSfaY10pIhHTlSeDOAQZHVB3GzjBoTqbhjY/3xiRrACy6DdSLUVwGIVMp9T7P
RX6zElcS+rXSql5yLFyqkQRaPpm0kLg2Y/lX5Xv7mRHdo5G7nwvYXpBKfb2fexFSJVDHyRRBbJ6C
8ttW0Dt6/1TyoQ/+X6YdXpUrQ3ENdSzMwlg18Q6N0A+kk8hd51T2g/PTpkK0I7ydEPeddp8Arbx9
qo52yPF4G8Ac6umY1quD9BlpQXI1HBpzlFK8E3KilcZjW0DR1yxDxeiZn4xqomzraZHVNKRGyq5z
ea1JMXA5fIyvjRaEsV/SV93RMlnxHzTAU2ARSxT6MoY5FXEYG+uMdwISffO3DhVseMwUR6B13BDI
Yl0QRvUdtuGMzHhN2Hr720JQp3JhGJy4xajOKQqaz7uQ0lEPfTM/d1hiS2r9wTmEI8fNXgYT2/sX
hKHcEKdR3U2YBUbWWJL+Jfc6OD6LEecNlj45jW8DhTZ6dhbcsrnSP7cJmSday418BK/VZfPtdexd
Vvj2Zc0q6DZPFK4KjonFEck8HwAbjlEopcWBnRT4SVU50T2OSJLdTuN81KlXqpBh41Z7btdZrX4U
vyCKLWQKE8E6tyEHpPE3oBM/wjlvDdz9ipE4qlQXmH5Hb3vo2W97ZHkQTg5zIlhM+mZ4j2yVw4QR
RftV3CbFlcueos2eqI9XXGtYnaco2XOAsqWjhQIKV9ttktyGh5qALJHG+qDp4Yp0WC6HcfcXocaQ
yMimov+ycL+99CbTs+0VgjwbzGHohnUlDlKILvHVRmUsU7FINcy23n37KCoxy87eofzgHu2hXdOU
FtRlbjoNx4ljZ8qGE8BtKH/+vJRbpSbX78YRcqMOoUMPS1KivyqUVkgrOypgeOo8if4pwsowdrM1
cDuXYaiBlq0JXX2Iy3paf4AMeQ3Qlj1QDvji8gsluoJ0rQPnAbmsmeRCPv1f2r9P26ejtoG4P/gq
5D7rpCotcWLZXRvmUEgq9gxSt7UBPKUHnfAxrLwa6CQvp3pH1KBy6+OX+H6sjfqXw8UKBVNWtBpv
FDqT12hiw95F1RaydlppL1+8d4vs0XUR41TF5OIcA/cBZVLyu5lGhNoIe4/zwENe2Lt55oQWY7aE
Bfl6TZZgOLRUFt0pQgFQDcPWLvIrH6GcOv7rwwZLgXzvngIvKxXMvdL22mWUYHPu4c/LdsB4voCm
ThkF4B3m4BzGFH6265kehIGIGk9CWzOsXpYViEnPDSn9JzXvO3DKhqfnWnP7hd/NA5VGlMw/TRiq
aM0n3eGbDotqQ9dsfyg4/U7KiIhVckzplK3Gqwe6BMuKugEuTlyh1vonEmtI7kGD9X8Qn3d7J6+l
GQrA+Dkexcyec7AZDtD0Y6IkygIS8Tqki4FMlAbsBjK2hAyN6FGFm2D1+/JTZxkIIvsL2nhLamMF
ffSLEAFTvZ7fGBE/IwEeYLZkhxAQa9cI+C14v8kH1PcnUXksHvXXGAhf5l3PBSonlUj1y7nSXqTy
zA69Rqg9T+cvvnLsCQBvYvP1sdbObe/RdDx0mSFmZYt+9zTgM5XHU5LCSooADVrfrP2+RRo7qylk
q7FcJEq/I2XCH8ZCr1CjMzsgDakEFuKAtMi2F4VIQ/b5B1iSyr2Sjb/dWLtYn//6o00OVrSsPsTN
bUNO5mLBos0FATQSohRpYvmIgLS9C7krWgU4JCujmsVRNxNjuRcqKJQv6ym+auaKqwo4SanFZnhY
Njm1U8FKvIMBbkZIx8idxlblLVvEG0+EV9+62MiRocq6xmw74rYeB4zxbwydpf1O1mRbmc4gqbYu
lHwLVIfMoA2OzWMzY7fGWSTOLWttvSTTrVzgAjeTHiwwjogxLDVY2pXUNoo+CaybIuRAs+OkRh4O
imWtpq+nOWEGcef0L8QN1nusoAlBRpdvwVU9A0WQSkAhyZvnzstIsWlDzVo81wCrQt/lI0u0F4Yy
7z2c6bQBtcsTwHnQ4EN4BGYCQtfYNt3Pv83OEcMi1ulexGfyyGpn9hPK4aCBnVW+EZ+uS5hBhzsb
cpcNsdGatZ6FwL/Q1f5sCpk3Xwuc5HhhutBOkDijGzDKpUFUGTRitmCYcvkdCXuQxscUbIeYd4/f
ouUHeHRhWct5iQCMyXFzakwhgQ86S/dcMVdx1Oy6uFGWR5mq658nse6LT6Ea/H5W1sTXnCQADYxR
G3P0K7M6r+3y/LXftbErQoyEWQe5ktgtvgrXYPARNx7obvscNkr/l6S2spOzLOoyFtbWmlMtl8nh
ktB6nju21Ma/go6vp24zhR8pZBncJhE9/ret3qXJuY/CK+mr7uTaWnxvLhBfGUGT3g+LOJKCQw4a
c+kEaVFMOLRf+XleCCm6U8GjowbcoC6Q1vwvz7XiumuuE2Pm7ihZZ67eVAjhtgd6ELhdRuSfwqdc
02FLZT0gaZbo2u9lPH5iySzA+oI9j4PzVo8PCZs6Gopnf7WA7M0XZJnzvVmpW2wiHHRSuVJ51xpT
elkjF6uG6GeuoV7tynx4m3BkbF4+SO9l0n/rzK3erK6YiP50J88s5hiL+8/KIkImWbJLBRhG+XVY
Ne7xLvFC+cm9lbDQWlDkEAtbRa6hpkxAUkhIzq7h654fkbljGI04OsKwgtjYXJQiWI3xaEAQiOhZ
DQje/CUCRMFxq+4eAa50lNMJhpuwp7jvxac7j/vXM0hZXJwQW6RPLH7K9gHTy2wj9yejPeicFjjc
XzO3AT8+i+Gb9m5MEVG4tRtdU7UUl7WcAMOp2vEzOPyKZAW35PuftlFFsrJYC84O8Hi+aZHC5utG
yi2W7GXTEL3uDo3+LQif73Q5cHPu1tTVo0JzKfX7DMYnQLmtlqrC53cuHjOIpT1x3Y2+9QfNf21I
AitkshIQgWkHDeH/MWE9Sm3r0uCm68KryrmLr3CnWn60I3ynx8YRLdAA1K+ryBZqX67TGOOqDd3X
SaSO6aaeOJ5K8Z6PgbKc44ZBtSvvyY6BUwma5KdeJaKbttyuypeFfTkkt8GkGbIRfOuyOvm70Qot
Sftg9i0vRZN2LzLM8wIGw1grsPNdmhtj2HeXJncPoYMON2mGqvbrn3Rl8wMhvW698mBQrkzNJKTd
23dpf3WM3YfMuKxtqi5cN9c8nj4/8++zESxwBuEZIygVApllncrM2faT5YyrWna+hxpUUPn4Gsd7
96HdlV16+8oocMPT3mztxvI39R+0JFxLKG/fKa+CZJnl6g72WtQ8rYavLIVY3gdpBirtWlB9mP9O
D/ctx5HWsaeiay76q6StQOWeygXI3z9Gb68BSVx8B65M5NiM74yh/gAUPel1kFuQD5gtLz/lBRvM
e6H385d186iydpa06aGIPYPDapBLiRjXI9mhipu2PjVQZ+DRskyEBA+05xNHRaNYi2irFW5ku+R3
yGTE6Di1pmX6DEH7X1802cpXEKX6leyo/VYF6pYTTxOK2GDrKzOWVBS1bTANXmySHAtkvUXSk0E4
RTqOAzVTsb2Icjf8HHyqqVQpMwGIJpu+FRS4SbxzTd0Jzy4Xy6meTn2lgOLgWfR8K5tlQkAnHjTj
aENlt3iupc4rqmnAXsS9pFC7U2YQbHtOY80j0liQSOxRGm2VmGqohKhwsTC0SgKu/8HgcK0lXb61
AgSO3VEn94gx60Zf+AXvqGwlDhIKtLzyW0SMWL07FzMqcfbVG7bKc5oIrPtxTGPVBNPfrUK55zp2
Vt+V96CFHyhUK6sEyMHgt01iOmlWwyR7sm6f+Q8GsepvbIiM5vRnBRPdC6Rf/58HicTdelljaMd7
m26bhIDQl+GFDUKrIYkZkdHYogHwQlJhhGBZT/FZgl5LtNVrBasCavZ4BB1JxSTOh8rYO3Iyk+qE
HF25G/N4gdpHG1yAn8CCsY9EBgrvlT0++mbGpoBDYb5HK/BZDTn/mjv6gTyZuK2kIm/C9qQ3ySwD
pwRptD88MYWo3fhzVymlg/cBiQ271g4dltZ7qBTzEKqvweq39PYQTyjn1Gln/mTpytCKLFVbOaAt
oDrVVdwM1vjRMnNKQmWV7J2jynyAjHgOOFMj2pOyBmFHrvpeDSnSx35mLfXsqIQ77BrCe/O5iyQo
uarvLHfd1yXJ4K8R1cyY7vcYstz+pyj1KABIGz0uRkHoDwPXe5K4G9yYDrKBItmwZytmaBo6ho9T
EubKCzrHFt+hwmgWnS9amPke0UgAiUIFbgsueFN5UT7SB3VVJIUgSTFkO8GjpOuDlH5DvnGCTxcX
CkGo2FfZceEiXCG7xbDS1OtAW0ACozHF98xRvqbzIwne+zERF52X+WJT6id400Ga1pe/ftjJ2FRJ
AqOEF5qhgyk9LmDTOtidq0EgVZ8g1FG4wpiyrYfMT8p9VZZZbTxmzhz2aWU+mjvEJbkbtIX+grF1
XNVuGI4n1k+xl7HqMu9GeFXbeENdVSP0kOtlnLgW2NFV8AsfYWpDQiA8ob8aW+Fi7hIsu79rib5i
WxeEcuemzUywcYRzFysQG0hPDY0t3VJ3Svb4nOailKTrqN3HB50SPGy1UkhR8/Hb9roqkGT5hsQz
Gz1dktlDIQAJ2sirO/Au9DAbJJdEfBVARVvEfrexWFi94gxKTkyieUc0ZHrTkkHJJh14awGfPmkO
1I4eUXNkT9J5SDJ4opdJ8/CVm7TUC2f2lddLC2XuM2R4MsMTNe5xNdbo1f8rLfEiQj7BoQtPYIIm
hhZWgCpixjS1ek02YAfKXD5OjmRVvtKgiuuY29lbj2182D9QX31aC6pFTiPQ5mhBQVoUL4DulPAf
6v/c3humaDRB9HhlSJmOD9OeShUvdOkZ3CqJroSqj2RinSn+8rKFdzzbQSCEHxfgMKcGzNwsErNZ
V8PlylMEPUi0vEUpDXyUianpEfNBOY1PBU3+jgzdmOt4kTi0RAxopef/e/3GtbKxN9RNcgOULn7T
at88rL2l6iJlvzHH2kgh0eLLvCPXSO/hXlwCE+oy1vFhTHKp6c7zvuN4dD+htTSEP0x0jH0lRabn
SrwfXKNjNJBX6eGouMgaKEjWVJswXEZQnisv9BcGZ/sA5JuL7lgy7dEW7UXYR6medxOx7m7flk6V
iHLu6la/cldzyqJyQCF7AI+gI5KUn0GBtVdWu0Nci7Hke04ItBUG5WDUbWgntGjBlfU+ukNaeEdS
CQrurSkT4oY3LR8G0AbSVdNm35ps/XB/LeFDsZD6vfknT7neOX2ZO0QVte0Cmok4zdDu/8JbEAlc
X9XG//1dTpOm9PamVoHaJQsqbhQQuSvFKnf0/4n1c86x/4ucao3Ub9W5qAeGk2NGR4HAX9cBVFRZ
CrvfwCZEFqkugzTbR5KPtlkhlxoq6oQLLkuEkxmiWLJxu7sIYbOqfauQicWs2fShiTZ5d735RTmk
4eQ1XBV5qt3kfHIqoRNdUtAJGBMl+8KBoM+UMADO4O3HqPT+yKN7zQmjzl0tDAvzU3QTSAY0N5dO
KDKvLcqfnr2/hpNoUHUCBD0qaWTVge0Fx4w1ZC67apUW0g7hz+92aKGtQ/vmxEUi575KBAnGy1v0
z6xJMIeaikEjqyWfjRrDwYUnTfNmZVw9dvPT7f23KPH4bavwBrSsFxFOFnYcwOpkkj6rarQKPLyR
nSLAstktde+g8Q8Lm3PP1L4+2vJw31cSkRgyr7hIScQumY58EQwKy1hTdaTTPGQLgQusHLefGgqu
zUT0RmD6ZzH/bPBJhhj5Q0RowfzNrpjFLiVHaw5sUVNRXsfxkSVojjTcFqLBq+LybCUKQE5ywFJ4
HAfCvRcEo9y/lqS7kjU3LUxxNYFDdbZX5uEm9ZB5bhX3z3x6jrg29yp3zijxQg7H7mcMXnu+oOEa
3+Tk+jngsloG2q0qtwiDSbAZgG+ivBj9LM7qoHxGXTTmjujKTTYEzYulwnEGDR7+rxZbmJXbr0e9
7uJz3eROXvyM1ycheF/ksFVEBTPbl8Uc2vaHG7BN3Y4H92iajwHxtv5oFJfn4SgSfGlaYSGSRF+0
th9jEeyx3zqWopZ5wvjgG4Ze9cyggGGDPWgO1ldwSX1UTqVN8ef160GiamOG7zL7CZghkHKJ4Spe
akPHEvhGPuVP5uA5MKK7oQrUkf7m3Ufn2N3E3DWSenq08pT02aWUErxj7Xzx1sy+XuIdV4YgwxQb
iQx8MWX2+DiLD6eIeRHMOR6/lX1fUhNz3sXxYaYz+jKgHlffW9nz5CJgWcAGICrAcg2MGqMpkNp/
zpXMNOTSMc20mLSF49xO6HW4Jdgyh1gS1CJx6T69WDlRkCOX0HARk7CCxQqr0t1ZsLwgvcDB9NhZ
JiOq6N03Ofz3C6O9+VCNWA+5ZYtJj92aK4SPc4dvdPFGVqs+VCOoYlWvixSPNdtB0vZvWz98CJ3d
oaFRM0d75ejL+HCwgnFkzLlG28ApiIqF6S58nqM51K93pKKNweDwjeOE818JpgPrG758u/IYlyTU
dhtrHQqBZx6JU2mtZtScagcEgOwOjT4FXv9CE+0oBzVD32/JphZaERMjUKDxkxRS2nivOuJ5qQNI
E7VKqIxZb+t8tAAbE/zoc2Yu+jv7lpREBPTJpLxG4HR6/AMY2Acbg5HF5utO9JcAp8er4GXDdrIr
SNytCGpf7XPk2EV/IPtykYDBnRzCXYlnbOBBsQhWAiMZuqDkJHDLoRFDBFZK0joF06oOEeDmYYCW
l0HC3kbJwQF1G94WOKlzO8vJ5ciyOpMwU6aW1v/6k4MSbaV7Fgr4YlFe0otohD6AcvrSTItVaZmk
isPfDOaFG3qN3YQEgiXIvHTtdQWDmaF90cUDbcOTNvKzd255meeEBwBkyqX7vdVrFv9lScqbt7Ka
p5XXrvIWqvGwaq+rG+eXS1gQBZe7AF60xPL1alwUWWCZNYLV3mlJFnGNULwVBLUBliP/jx+YP+G9
7RjeJ8kbFnuCVKMK9D7dqn+bHvBlV8GJyTPRn3XwJ58UXjZWc4QpMEuOfNSXPIVcejHIoBWpftsO
fRlV5UYqWbgZYVKyqSXg7T7i4GRO+KJe9wzkJHpQKvWxO3W8/yyPjM+hXXdxcRSvrLwNHxxc1Xt3
3xwILA8ddSSlBQKXJpa6T5dy4SRvam1DcpOTbaDwLwXp7LNYgfApxf+YVjVPaeztTFJROXgH2UXD
OoQfuTfgqYJEQVm6q8XttWEQeXJQWU9WZaMLjSaK+MBNjw/Zao9xoykn7XkQiGCom0nCRYhU/TLi
tbaN0jBqGaNj5r+iuyTNVZ5mw4K1cFA9YgLcvQT/1gZ0MYcHXKuXw+sG0br9x/9QPQdtlfY7Tll7
FOwNFYmCLcqppIzTydPVf+kFPAp8zDR659SoezTil1a34L6sXleneawZTkdw3J6s54htpaiXOc+P
IBG4AzyvTPISxUPpUzQ5dgYCqMF+Nuw9fILjilmLnqfPtJtaOp2B6uLeEFoM4K6ZUa1iAme/qLc0
wpcJUYnxP0i3HZgggw6cGe53znM3wSJVSKB3wZOyRQjA+jajeEqQU2iC1FhMPFZcADaj3SPEnko6
IKViRx1wCLaP7zzeMPjoCzYMhEQvkZrUyUd61qkFBcgSzGfqTAytcuxSEXKd3B68TklLstjbLmng
61KJchGxuG3AIS+frFxpCmaM0OocxmMpE/DbaK47/JOFRSjM6bN23In2WMfBx1o6IAa2mdHjUe90
6QyNIbz4aQWllWoqUiQoeIhRlFen7DD2v+LAhzEV3rf3v+NxEA27fRAKOf+W7LxYJVHAn3WPio+o
ZcRFrr+daFmUd+i/BbbdMagCfgxanZNkJnDImrqPMiavMN13jUjIxZK+qr2bEthvc5EyxFw353PV
P1B6ktjcc1NuR87lESeUaUla+Bm6+98HjPG2pgs2kwY5IR1A7PcekhEP3CkJ7Th7GO8aJuxtgToA
7yAtOpNyhaxGS7RAoNoPT9uQERw+pLZj2eXqxH44B9RE1KsLgK+D366USbNq+8u2KNJ161MTNQhs
bB1X+daBC5N7DW5VEiheNDgddSvvnCg7y7/5UD+XEY4aWmy7zzlUNYeuSY0WUsFanuk98Quh+zlA
NzQD/aeSddeB6ZTztBCWd0ae1h4z3KGF6SF5nkKnMGzvhTUo/sOOXp5eTrMQpRdJvZzCRe5SQ2hz
linKEi5wSLtl1I1OpWnP+9bJJZgfYN9iLzwDuSPMuW11UPuFpcKNRMvLJHl1ZBMdTBjlKwbpVD8Q
Luv8GH4vyarLdUcv0kooafmsYfrfbZIi9KMnFoMxg/PpHcJPshmwQ4PWwP6sWEBkzAQmew3ZXXRy
h3oYoAxS8GYQeBMThKSOjH6LLpxHRgo7TFC7dHfoNFjTBZAaM7CtqubImiBPdYnp11rdEyDMYCWg
uzmAiaPBg/GU2vHffUeLOmfZ0uK1SydqP1Kt2T+0r8hmsl5D4v+qkhla4Yxt51T9iR7ow4DhMhd7
Kyg7c9cGy3L3USzlXNuJnOCOeWIAweapipSBeFNsHaS82b8Kg62tDdvECUMSoPZUI9a0MA4fiXZn
Ykywfzaw1tzbC5ApQNp9s5uLnREsqN1Nc6tzUdZfr5amqFme50BFPODtjGSxzaNopI5M+iiHxGsx
lc25sxNoC88MTccWcSTWSYXWxKVRmlJ0PXhZ2Se+k5pDlUi2CjaFZqW/5IcjGWaqPdRf7cIRxTwL
pxmK6v9VAYAeBVg6UTUaLo4sl6ieuh5hXPawNvSJj6GMoVr7D9vZEf9XcxcUPyTinmeEwFI0ad67
1Q/I4xNj+n1CG6YiZaY7QCr8dVxDrFNps91vW0J/DrGsdfAGrO3jrOh3jkBwfzF+OFN0UjVX+vYc
PkliAjDcYa1jlaT8JGT5PS9WKvCINBYe7Z6ZSUt+KDuwq9ZYJORivq2u9HkFSJ4BbSFo85wMAN5J
iKBg4wl9qhjUF/rSP8AGn6YwEB8GFgnJaxid0iox4bq/K6RK4OspIbdE32zXmGOACOFdSzGy2Hnw
b9vfokaybVCk3bImifYgrieHlSEFems6lPo8OSfI+Q3LbqeGTwo6+ZoadXSLQ6OHoGFc7IKmKcTC
b/tftrZi/TC+RUtmdvfCQtF5EtljXL7Qs7ymay8gKocrjV36KX2JnL5gMibbXlkPBiA2n9DCCvfi
+F4QPj5t5w/tJlTFnmuuMt/u1Z/QLNFgRaAF7OEE1zzRCeawtt7idWTPy+MG2e2a/pKUTGFjaA7k
9rGlxb4pnvis7WzlUwWvjyjkYhNdIuQ1PjdpHFIwGd9uij0L9uLAp/BlThwvH5aV9xkdV1l+wrru
gYK70ROrmKxzLypen0r03WOBe/d+VypzGipdG4MjHGpI1ZZuBrDL+Zk60XKFpqclvd2lDmQDAqfG
uS+qRK0uh+XRT991OQCCeND7iDBDbFA3DYA9ux3MQA9RTFBLHBPTrZ5vfnL/R4yCY+G9q1XnkE8M
38FZonqaF0v/xIZ6+hr7vkiXoNtC9lCZzjOh7phBgeuKWeJWN+GgIE36XFu7G0/r3pN29N3Elfrs
eBWmk+LPd6G4CrJKNyvbpzUUFs51fKeU9N0cocTSMVfTkM8pPb0iIIAj0jlTCidhGEc3jkfEu8qy
HD60wQxPX3VJ2G5CbPixzRyJK8sc6sdmltiBm/a+RUSLcaxNTzk+azlyiLi8gbFbR6ONOnFinlbj
NWVjjEON5bwKlct5YV3O61n9u16QkHJ+PbyLxQeD0Xy14x5rfEgQRYDdddT9ipH7nelsT6T4WC9D
SLzF2bdUk/o9ia86EM0QG51oSw4DSXFeIUcDkswuDCw9eLzShWBtXUGavd9FyTTrfpZjdJqhImEl
Vm6LwzgXSweBb8F5g+oFdcHDTr2ab7ah1KfygAm81ui7k6C8TZjmzmh91heOLSCHqG4ialDnAPXf
eGAPEoFVQwCjXOE5GV79hXmL/tPmNh1UkKWiy1EEE13OEL2SuJI1NW1cEsxEpZ+FMZUT2Xk+hnPA
LY7qo2rbiIX6c8IvSjk8EDQdElaSiWzhlcZwAv8vN2Qmjjj+EMjLrwXZFNH65I/9S1vK4KWavv9t
zyjxI5Xr71b65uvgd1KgmntKeVEzyafLyWUF9nYpPxuuAd6TycqoFNbswEPuHX/DSUgYn7w6dTnX
EDV0f92/aY3zvJXNssNbsoAYCXnYb45f7QdOp0mZxC/EY3aaSf+zXHru5p1RG1DWrQpMR9Kup2n/
VBSWU2bw8M1Q1ZWpPLy/n5yY3F+lqE6KVF790NZKJjzvd+RL9ry90GwsgCkhE/2lIFdTyTwcEKgB
fNHOv95VC5iaoL/H2UEPtpmdQYchplBJxcIxJoOCo+V7jLcsolRfty7tmtkTaVjWAyZ3k38U3pCR
WGNXWTce4sjSOuMzX1XbHZu7iTiU5PGgU+vc/10ZEoEmG7QHyn2Jri79OgMqoY0ZPzER5QMru7Yd
Hhm7q/YGfBYrRQ1ApIVA1YBCza07R8HswAAX/2JNwua8si0jjdYAHVlCMu5Dj9yc5bbHMPNjdFj9
Uvcm1zTbSUOH+wTtNBmgQyGW43WiW1uodnbLlA1mJvytghd/NMq7BL45S2YpYJ39ul26i3UMFFmY
k1EiQYzhgSFSMgJE+RA9AdYvuXPOfXrY+D7VO4+9bjlzgKpvwiM1EL4Wz4NrSlLHou73djyvsnsX
A9/OrELA6VwQm+dR5K8USHIv4ebgzUS0+tpXj5PQCCQZknSou/eopRAIo8pU6cVC3H+y8aWSapVd
FoSd7Yx4etoVJajpHPD1e6uKpiRtXdV+fY7uLIqMxdmyplHfOz8YuUviNv2gxa15+njLgwC9Yelc
S+s+XHKcJG5ri7uPUVgUxiBcXltONiPiQl+QuTlKDabtJayLHnZK2SPlkf4IJfYkfbUi2g4rnc59
8AS0hz3ymAAddRAGjUYHNRIzvcknm8s8uaQlFKhejcHuuwUrLU9Lp+LxT78fmd/85I4kwwgQHY3e
/H0X0o++UGiy91DZN/Y0L+a6Epsi/jb355uSw9XPVryWZ3L/HHNoe7I86Rmz0dnRDWtjp9kqTAOW
QW3Nssb3hmlkFf147uRg1huBwcA82zNvCyz3zAG/qyjTZSmkC869Idgm5dkZRo/Ol4ariw6FtpE2
8x6vz77bBPXyedRIrNpaVOGgTxl2XMfgmyJHi5QKkrAzjwI8xAd4D4kG4P1g0Bl4XL17f3puq5V1
RIzJ5IaGOPDQrjHoC7S55GuVAebtiiS79Mpg1H8PBOuEcIm5YfQ7GIr0qVnaUWz56TkkB71hEFIo
gQU8Wx4aEX+8JS5F4n+qgCdZN1KOanyb8qKhLyuFHNMc+4u7F/ul+Wdbf6RTWS28tZJN0rbxLCkb
/SIrhT+SBI/csuAyJfKr0ebeK+E65twpZyNgeyoTQjWf5wn4CqSKgJoFwx4mJk+IrfltsOQVZ7Tp
R2UQMElZ/jcshzMl0MiHVbTRTuwXUiBzZQBvkDC8UoMBgkuYmjAETiI0IWrU4arikfnD3Am8ZUQX
ELtE5xnblvC4n9MeEbrU63WE7GGPxcGQCwljVPdeiGmu/trN+PDdmIhBM+rfxnvvk4lYixfLuB9u
i3acngSAGPV8xPgVEC/0pELv0Oe1mTSP2lrK7kcYXImELkljSICMBFsoEPdPtYKYCCZal6PoEyvE
FgIX5wGwe59m5uYWYhfgFNXxw10zLJEbKULHDfdF+Dvfc74ioRlXgy9pmkif+b4L4ZY8HcUPGV3Q
dd6Kvbj9qX3WgtebT/Vnj9slYu/ag44aufY/PF0b/T8+h90WQ3Fr7QOX+dOU2+7GY40W+DVYp6BP
AGTCZsRzn5SgxT8fjYGL2RABapg/2mJ3EbcgUJMBERHQkXOwG6Y2WCglNyw/aScpcNwA7nVCX7C8
1FPqnvjZrGqjVvhlEKtAzUX5hOmNjW1QneEl4TZdCzm0g9wL9adPW8w7iyqWH4plIADi5JY1buo2
CIrDA4GelziciBQbXDJUaHwSH6efAFlCmcWJHjErZnSc/1R+eMF4VpJhvovPam3bPjfNsXiQcZuJ
IPBvg3s2CEBehgIsxFip3NGtH9MAfTn0fIafGBe5LcD4E9d9AXbQErItpI9AMwvXiFBn1ycx3GV1
ur8WwKvU+CJEVP6NnsAMXP6rbWX/UVj1ubNkXNZlwOBp7pmSP8Jgf8tQBBe+U6VGyqHSI/sx+++P
5cKKCIjc4D+hYilosB9swhZGYCkBuNpbBzFx0T5AxyqxwpxHroAPlqbIipgLz4juQ5Bky0CzN/QV
W0ghiG4eHysOyuKRMvjfHwyajJyqsPCCcSMR/ZEZDEDaQlQDQ3JNljsR01u+vNW9YZ0sXcnfIumF
ovt1sp8NtuxVxDh++fGoJCl2z2GIe/ylOyJXsB/Z6eKK0cLqhjsAMuMbnhsQ+pK2UvyRAQ+s07cH
EjuFVGsasJozbleFpfpynXsz2LajK/mXybwAcf7lMbgjW3y4uz3Hw7aV6cfx5rzhE6qUTuOs6ACZ
XreX5id8ugGh5qkn1qo+1mUZ/P5xHA1aC/xRDRHn5Bbw27vX3FcP8/PwWoubFMGiSjqqX7c+CsgP
lNxa7QeKNe2jIAoHglwkGh0OxIiqJNCacSZ3bPafJMTaiJbZkqoZOYG5+IVqaOnWRaswcXcvvnnw
hcV5WqUn9Ok7goKfAwlHsQqtz3/6fiJEboFiAmfvErVfgwBa3q8aT0KZOpydoiGGULgjnrxH3n8J
aULBY23pzPuwpCX5PO7kSh6zhrjQcaZt4voKagkXYI7S2FN1PbEydPTnL1scn/HS76n2Gzf8emt9
QqL4woKd6Ii1kO+UjcT3Ib0Xjz6ttwl1AvAWUJl/+bMmYdzP4wgIIId4hm7bV1AxuQ5wXeUi4BTQ
06OhNvidIHMsDPLDJk7ECjCFKpLBT5g0R45sVEzrqlBUwqLwiYvwTDvKPkcWsfVkQpAh/Z9oW8nn
ZXOcnTSSutN0Kt/gUEOxLc5ZeJ7XhJedk+WyD/zW2QYfq02dd5ursKXTQdGoOjudxUuXVeopdy+G
kai7E4uXkSkZc+WJg5qtiA7hKQfIYR43b74hU1NUtbk1Ra7UtgivO1IymEq6bhNDFrP7Sn7OT1aG
8tx4agkICib3VAlLCfze7F7BPboEC/hZtCxUQT6r2WQv4XefFDbFUW9mpLlP/lz8UEe8DrrGFh+/
UB/naMsLyO3eGZGnJkw5eUEogDpz6kb3nEKCwZOoXwr3/jy9CRnKRPZUaK90Lh1xZVqxPosagSxI
SrZb2AnJS9qLJWH2XUg9FmSOYRugVwSAhgFGLjqIjmCNxmNHJzTLFAF/rXSNAefB3t87rf5dgvBr
8uFVrAQf+J04hanlSlKep7cH1y50FfoPKd6x+zfNf4nCPFjMVADE68uCYmTtT5GS+MWk82LdKByO
Qdi6oj6xSmwIYE594tqW6zAQqRf4IvvyUvjbCJ2dBVpYull9kqcgMabAiRNE9c1y3MwLVU7IppA4
mbp8s4Yfwl0WMwwUZKO8Y/b7JMWBAaIzEWUk+NT0HmmR2y/uNH8593RRYskLgRWVdS9KGhxwMgB8
0KXHFk0Z0nSQrngXiGppVog0JKfws17VC2KEGDqPpeeHdL6ITVMhoU7unJLYNHGudqObNCY3mEOu
vRAsAY7hFZtfXctj7o5FKkR2R5NxX69aq55jUNADlWoa35q/vRoJj8+FeYVCtEu3bHHlkppdw6DF
FL4r1dYJdLvwlEjp4y7hqhtv0ZsGK6GSiskKLwMTvO+F0erbWhY0EUiZg8XehTay0QSPg9vY0B9e
xCBdnLyL7taDWj1Yg/S5pejObrFj6Xv+Fyz5PS8dmCYZrsSJZelF9SNEXAE4OwKyflk9wfKbwp4f
Y3yxH0KtJBRKkOa1zJAc65EKHRvJX82fR7q959KK6z3Eb1em0echJks0Y44k5XOZWAowVK1j5eCp
gedVTLW+UQKXzxBxlk9uovG1LZCvoD78+GrtKqStj88eVAIlYiRlcNvE45Uf6PUb7MsYSpLHxrZC
8P+0L8mschIE4liiEp6Z9JnP6Xfwn/zl0iqFuc09i1/LZo1R1XQE9kjqxge8n1tvglnX2Tad3K7+
O88TyKmobxR+MAhcp8lfz3f3AdvdXyu7g2oqeJv4qikVFm9ogyh0KMJIBTlsy9PlAzyYk331Cwrw
xqN4hQ5IpshcXDyPu05QvgzydplUIQsgppsihUsbB7zAH899peEnz4C4uCYN8XCgdk0VAupM+QU4
9xz3YH4KhygQngTh0kdwDn3ql+v3dzZeGQq0twrxr6bzY63uKekZ2Q00nNKxPsTikD4g68h2w5x1
mCwYQVdRDFxcGwlwhCCDtwih94q8YRtIoxK6+9TWJJ9E5fYZtb4j+kGnedV/riZPIng9Vv+OPa/a
MFuvK31CEJp6HDxbZlLN9tpP6BOSn20hrLRxwmPSKmnH+3h5WFyNJMqTYEMD/3GOHpJvf2TekKHg
f7+ht0QBfyzDkDuojgZxrs+vw/OIqO2m6N8axQHL2l0S4hogStetWL/1AaGkPoKvHbm/DgpA69Ry
p3Httjfq9JK0Z/gxRClrEPxDFfALkvmB6AkIPhCZuKNqWGa5EN4XV9Um39un1Eh4gUzvS0lN2nk+
nBEbA6vhI1KhTIknuqufttAAtmSeSG++ZzcPHLU5dkcIn7tAxRazJRKWBeh5BRpxBe9JtAQm2u0K
0GP4EZxvLqrAeCrB6ASvu1TvIkUkx8gOmCcPTzwLzHTx88+6zKR/zI0j0mnmu1XA14MkxQ2I3bZa
CYDBJrJVa5j77dXvwgLPF0uhZTLo1XMT0glqBUL65cHkRyp+rV3mVDiKtKsPPAt4KH16qrndXU2S
sMYK/nfciIFzQBJhJtqfZoKn5B3GS6l4t54DzITEQBjFhvW0NaJ6BYPl8eSa/1qLOhmwRwilvy0L
Pj8wGBZigf0cIrKYM2CTKNbvqbmKsUe5VVhbms1NWFswMWYD4YV+8Wv7HDmF/UXJZpRzPu25Y6v2
o6jxWpYsKRRXncqVHQl++JvqoDTHzxJF/E1tOzIEIzYXTOvntc6oBj+saUbQfy4DXpgDgKH8iNKW
YvfmzjOKnXm2f22oH2sPpkCYYQqGyGhSTQepijXEdrMU/SsiySZRQF4QkNAG2I6eCff9UEc6wnSD
iD/MCmEKM4k6VjjGv9xfAXB/1eYhJ5z7nxyI9lkLiD3/rBQAc3AYLEQV24I6Q0hzzRQ10VBhx/qB
sS+JzoTaMVqt37ryyiSHag82SP0e7drvwMxgngEULBBR1H+yAG4P89gB2M3Z4i5H2aIK2zg53PVd
SOnJQGxsQ/8AtniEE0TkUWzjGjWjiMTlRgkEzeLWB3hNRT0Og8vlJwkjFgIbdjKYH1LV1shE40bq
fY/F+knzzWBz5qbOLd2GcZ+1yEpVRQkyKeRXI5H7SU4o41NjUexTdp3XhEj8RRX8RkJlkWoX3/qv
IN/W/WZrb6/8FtEiODJqhyDnlcLgOtR3pQmqyBP8Ie+nmY0OoG6Hp407WyluhfrPKn3lZpM0cwZ0
jcvNE/xKszd2mk558vxoWX7h9LG00VefWz3UO8F04wu53s+Yws0plm8M8GWDKMI9mBY2eaX+iQXs
gNCrUBYf6EABjAaP25voAnwjpEZ02rmBrMEV+N4/2iv69BRYLp+C60HUOMP6hF8AP0bqRjU+FOea
RvNJBPJsMQ3OTsLYge8KaA7C8tpHJsB7KCdLvhTaNwyvcQRGLuN+j2xV8cZw60N/cCsXrxFB9Zr9
8FB9pztsu2aHazr1kuTqmMdyJjyO796ND1FWjTaGg/ACo8vueSwR8yCOilnmBKnTV8XPINbYr1dx
pPfNHyuGBQe+X1NLO5Q6/8oOGLj8rFMDYaMlXEFa0IvhTd75J4989DqQFd6tKLRQn/iS5Q68EPz1
bfXxwG3ir7mmke8X+cSvoptoJsqZgy6mOJm7+IiCJEKgFiMKCv5yXl/WQrVB5EysBM2EwmOBOQg/
87qhmjcwcZplcxg0u8+pFgJBHu/HZ9KIvHmkUUTWbeFtZWlA8cWJT7xQH7nK1EKCi2xJsgQj4VOP
BswA73lXhANIyyNGJO8KEqFGaUyJf5hchpSpQMnLlmzuq2DMDCM4LMSveu5vV70bERrvHhJU6yx5
AN6z6Ba/51pvLZywR/zjPkwlqG+4te/8ddwpwoy1fNwjdvEqAlT1pOvxeTjP4wSS5ZdNoWt186h4
qSfMMvmHEQn5kzknZZIboyaz/n1OBDH4QQenZAsxPbf+lK9YRRXJvS+9eCsVPDtPKwmCoBcDMv2Z
tdyD5kyFrAbpWmzzXR8Ftoc5EpSU28rX0rDPQyA+K+csKuWOdvRIvrItuZAayS3bs6j9nCF+PRt9
kNrjluWXrb/A/I4uzgD+RbY07jVmWNVXrj/B/mZCjCWuX8BPdGLy6yZFrGYLQtBpqKb5BtUmIW9/
u0rcrq75lOXtUh+zgACyWKmSfIeGmcWuWMMP+YwhWiBw30TlMVS3OsmEMika7JU4Rn6EJ+vsRG5d
m/nJQNg8BkoVTuvkfGHDH7RRm9C/3bMPGLQ3dZBQfT1yVIAwxeFX4Wa9jVYrGed0S/HyBCvmdEq1
Dypr9HLCsjtotUVHmT1M6VzM8IgAfkyMq6Q8ec3eWT4Gb2941YPYAeMYDaqXE7Aht87o+aD+fwrX
std8BtOxnwLuhXoRjNG4Nmny1KSOOdEUzLj2ptnt7YlwqEfl1EVEzCjyNIi3cNia+74wrpKsMIJg
tuYfzLc5t95QnKadWgpgz2WCdYn7v8/XVE1U25wXx/1jGDfeQfZL8u8qjzb23FoKaBC+cmx71ozn
2Zq9Qhl9MX4lIKgiHvMPpj35YvRMKTuSXghK6z/8va80jegUM6HYU8BJHUJOZbgt38+IWM2P28e5
buHKtLmjjwvgzv/Flh+HyHyaZwaYFHYPsGHBrtFCxwaeYpvUUeAKfUbMEOAWwLZHhJHeAPRzGivT
AaA7cnB25H3WS5aTBfmfab33aiu5Mibkna9SaAzhYsoj1ql2IgoBABUc5EICFImEH6UI2yh/hhST
sZkTMUqVxmE5OBuuCpgKHGpqpnFL+GCUnqNT/PCqzBOSAHtxv1rDAz9RnB6BRgGjnyC9tluZniH0
pJyodWwMv5hi8FBk2s9bteMgE3ePPVY3iTOae2u+/y9ZXRsPVpXShdWuxRFXC9cS8B9uuCJk1aRh
GsBuMYRaGALgSuRdwvsWlxvNh0R9Jc8eeVnuRPw4B6Xj2CFkkT1eNgLIgfMsf3GmJz+Lb4oh78GZ
dafC4nckgIp1uRN+Zs+5JIhuBiYh0RGzUjuUz3jjZiccu16MLad5Q5eSc7WyYiOajTszBH/SA03U
TN68lNJ2htj1nwXi1fGXH5IaEu3162cxW2nwXiv2fIxP+afrvnRQEkldS94JKAld7MmkJuQ1xaS/
2plnjEbu+wTO0F3/TZqsfeKbcCd3KhObCW8nJBfPMuDCUxcKW0oeo+tyjFgUmEg4n0oss//BkS+m
sOaYcID6t16zOJw2BsnCwP8bBDsY6vP5bqkKSqSMM1ohzHwlj7DH/5fyMEEBDepZtuL4WDl+e7wH
QgKkVby2p7Qp7asU+4Z2fmkxoy+kIGm8352yP2kFVjphvjqqyHID0fvbBfo0UHxbERSPAwgYyF17
AE1CLLoydkY8A7DlYl2Aer0D2ymMBcuY7LXIpmEUgEwjzu23+Yvmx0V2hROnbALvwpIPiyXolcdP
rds/xfo7NqSvdQ4BLZU5gbwZOcJ5fiRHkWo4IsP6uoQ0K45otq2vu+4mu5w7n51EMO6cUAAGaDz8
k99d6ilTrWdAGWb7RlRoKm6Pw95MEfLB88SwcJgLqFAhfv/tOHQH7bPpCWP504EL3xkFFpskD2wX
lZfV6VvJ1uYqdUD6j+irgvGSvb4OfBqaJRv6f+ffo9Ym9KAf3EZhwj9214sZWxUFqpaF4vNr+yiL
VzpNzQM7DT4qLUry24OTJaGuOh+mbfmAl1Qq1G9kaz8Bsm9zRqjtcj9AiiY4LErErDoCv0fZh3Bx
EqrLAgBapcb3yUbcKv4RYHKEfuZ7B6F+qEJbGrZKyuWFP/D1nvR8kGcVgI2gNqU+gvdZnNC4ZoE+
tOiPSozl7haL1BWjDA0rJzppKNkmAC78mE7h3NMX3hIRdjCIdZVDOGh+uUOF8EyxRu+UI6zAG52r
Je1hBybhuv1JgThak7knxqbEZsylLhjD6KCmZPaIUok1oVFT1jawkh5BLiVn0wLg8Sra18MEnSmu
Nih85maRWRRR4pHQwIMvPaWmIWOIxVfMIaAaG6Vhb/Nz7CI0nFqnhZvthV63jYO6vzimyFeJXFQo
gcFOGXvQtxH0q+vD+bkTv7uxvt5GePT27JYR1OVkHdZR6YUu9b8MohPu5Q3CqyB8KqiBMN8cSE4m
XDqa4r/6bNzuLrXVGxRdPyHQRZA2A5yOlx042gpQKtLnwaQE+R9LN1a5QoZKcsPX4CKizYyVCBAS
OGGN3X6Z+eyVwG/VLF482IVAxcbCSmFE+0rVV/gennD6Tgnhqm8faX+Vto/P2QIHggUBqL6l30jn
uHnVKDOBC2/3goOo/CB8fMC4DgHXvgexVJHZ8VLhNGN+isF+TCfgwnXkQ8CMhBDyk2FWLhC69Tdi
3GGX5RTumrNgdxBCUBO0ZPFeEgApE+onPQAwLfj0i2ltVWerjSrV2H+qnofSW+JF7dcW4AjOMXbZ
0KGJvIlY/g/91ogh24WHZJgpPpNN+n55EIYhz46PyzcVgizq+b8HP4if88bLZ24oUZWREBJP9bQ2
86MzDmh791RHCLvZhlC0xVX5hZIa2ub9OBdNkPqehdQo9LJJuPTJVIqK5zsm5g3p6Ct2M2Niu8iC
0pWloccHpW/kQ+hdjxK6DS/kH70zHyVP4H12a7JIGontGhXjgzgT8v5Y//7JnNRaWH9iJwVnnU4A
aXLTkMK9CFxwvfBZEc9/FU5y7lkwx3m06T1D6d1DRuyG2ehR0GtRsZ+YTRqxkkaJ+XwsGi1hl8iE
cLOoGraCacVR8OG1ftI6AMMrd2vTNP9WFzlnBelKYizCdeg6o9Yw2AXIK+riuoaZ3Vd5YuMGfZmX
P4Xj4rgDo83oeiDnMCaB6vSeHFGgKV+aYStcUGgAPyC3ZBdqke0QmQPVxyngMlxoDK7Gd/OhAkoC
TUNekGnX3v78q4nTzEpsMn5AScoMuFH+VFm3W+Lr6tDXgkEAJQ1rN/UT8FNYVuhVG7NS8hjEi/rp
l1dCpRL9o0DDB6SgbrrcqiHL239/A87jewckhsovGsVfHWy6c84vUNDakJDO6kIkQXsiM9b+2kXs
nnGZbq2M+KqhqSKmecQH6UTJCrwHy9GiN2Ne1d0XnajauE4glRXvIlC6cWeeca51COYGA9zpmZKq
VOefWDiSwTaCtay9kxYXG3IbOfHF0/6bVRHLeVz9H9RHUT4BXUqkPz4mOuLf8YZ0y6d5OPn/rGwC
TT1bOQZAPW6W4qRHv9WqLEP53eNtffpynFAVAU6hlQ0P/loV+u8+e3Ejac+I1UCnDOvRrkDRi19M
AYvtrzCvXmgMOdO3MTSIz0M4LhblwCU4CSsag0Gj7Y5QyZ62Ek7znEkp5XtPIkI2LSwNsHFVvTXz
rs7c5VY4MWgaTNZkiMM9ncXGctabQD1iS1g7NPKibNimyNrJc+1plnEvrL/MiJ43TT6YH8ifrm9k
oy4cvQPfQ+/J8oHRft/dsC0Ghi4jjirUacHzwOlhFSAMttEEhcvLWI5xqqtgArYM4MpnUQuForhW
Vs/sQefShU519ycJHEQ4NDztwS35M+IrChFqWcyUBL/sfb0Ne5FLMKETuJ9gwTwWZv9hGBB5kBq8
afVE2st5lKnDzXm1YZ960xNfjFET0txlyJRdX1PVrkmgUozp0siLuHxsaxDqbyqCZXsmbU9SJ5y8
KO2JvbCdGIrYMVkEf2Qn58XO0/HfDMe6oMJo+7NtDkciCeJm45JwnMsQ73DiKP2Bs1KBt0Mk3ES8
QYkN3b2tjF37SO2oVS4MQNuxGqTAYPvJk64ANVrgbsiyMN+DpAbAPQP5hcIt58fb+EjRmA6R/TJt
16hgatKtyXZ7xsFsizoYdYIrBdkTzYSFbiXEpAcCORWpkQKIJuDuwAV72TFiBWfOVmNy/QG7xbUt
vlwCIOmiiMAHmFsXYQC5dyz6rnZfpRcU3eR+9JbFoRNxYaJUyOaBNVSoRWYEqe+EnmWa7K06u7me
HoesN/LmBz7Fod3CVHJ0EGv9xR+CdtiP5AmBrx6FEfYCYqNo8zYjJl7ChbjmgtgpBIF+MrlJfs4h
F4Qri1ATqGuBLh3KF1WZlgcm1ESs0ydNGbJ+tBddanHfX/jXCdq+Jb5D6gbKAwQBuW6Xfc9ww1p5
Rnnniqdjjyhk8igfZjHuXMF3eFfkIxh8dHcy/O8yWeaIEhniiqc9Ql5gYRIBx2t3hElm8WAkasvq
hYAnRZS15EIH8mZH3VVq63CK30LqNSpY2ZcIePSNLLzpOAy6tqgOemZvTtUy7cSgqPrP4i21TwkF
HAWuru/06W7hFgp3BnhSXLIQXZqhxecfcaxysgDn6zRC//FFV7fPoL1ht69DjL0bf8+QRvL5mNlW
pFrVcTEQMeFL6/Fhp/s/s0o3IYz8exBTPghq2c/DNgqKcmbHdthF1PsmzC8nOOMoE08XBs2osRZg
XezaS0LFpVRTB2XfxvqAsFL6Cuab5v1BcBYVSIIGfFanVVULDMRwL85/bc+C9OObIbVOtOejvTxA
IsuNQPmlBzobZtZgd9q0Gxo2ywbrAagVkDkZ2LgxqRM6AO5THYgiXzHm31hl3iy3Gh6zecoNkLn2
+a8t9v1rEj7NKopeshckNkwpV4UwxQ6ue9lPnBZzoUnLjI75sHTEsHweZU/+hfLYbJKzc/zznNUq
BiGplU7068TVXWq/4b1s3weQOg4ckVqmG87Biscfy7fstaoErGts1L9zXOUQm7+7xf4dkKUqoySz
Ljw4AYj8QunzCWDjtE2VZWXHuN7cqv+iiUU56lwL0f2YUiLG29tioUc/BNWY7QjJ32QRYtrQongO
WT18JNq/BkBs8y6L9AbKF3yytL5trQbwB4VcSP4qbHjDWzlS+s14mk0zr1AvT6lAwKlmDaVeaPjX
65lSeOQLjJ6ejfx11oPds+tIlE+BCZYK9YNY5JgMsWQ2FCywP+X4G6etDiMUA/MNajx2zaxbqe72
F5yH6aH3bsekSIeeM/g37xT+leDkY1HBOd64Gzcglbhq9Qv3ThdmC2rAmCPvVHSXEDaWqaFqdKCb
HVQpwXtJWn7jZs/5wXLjduWC4kcNKF6yFVAjsCSvddb/sPzQRXlI8QXnIMMq07qCGWVgJsuWg8VD
/SV5/3jpf4DidWUF6UbBoFe0OiIZhgE1dXi79IamMbMhCuPE/gAASVsZzQ09QieJ+RTP1gGiH6KO
cC5z3rMUHnydbjJQ8zHd/iiyAfd5BspFsDb9RNahQPNfugIcIZ5/sNTooUiAdPsS91iHwYOV5cEb
igL/z0Db25JppPXklJSIYeHceegvv/2AY/vCjPm35fuLO1OeC1/o5woq9wuC/dj15p8YAmld+gEj
+KqTsTdMClCl5OlZ6KR210TUIOB5qK7VIahcHNsNPbbCbLBX4zA9cRocVXfB/ZmL4l7Goi88RmIA
njHGmL6TcOFiAW1kxljV3bBnlHg1fYQFJxG4aeBxo9o+b+ODg9JDlInOEmIDgul+GghYUbDfZO5K
gJny0Q1HDUvnvmyLtDdSNyxZF+E6+O1hOJX8qvkfZeAol9zwdpLqUhj/xITQhdFmWi1WWeFeBn+h
5g8usFWS2YIJyj7k1WAL+yYuA7ZZpp0vF3dWHK//ZfZX7IsjL/Me66Mt3pSPXMdp4yTcrHpLu+nz
VlpGCiFZZ3NbRffuAYN1OcQIj0TEwMbUFm9os1OxvjbKuZ2uCK4s9c4qKg3rjbXDiZ0fboRuQJ6M
Hj54sAgXV9lCjSGb8jlzJzUJnbNap69j2cfs+bftWwJnA/vv0CDEJuB8a49FDjqG7n0E9wBX8nr+
BphUbPG3vUJYJ3c1qhGC2uTLWmZeLnEVcYNGnzZV4UEnkGG0UMwWRyzjw3wgzeAagkzrMQ/cXrtM
OYQToi4+OKQgQLrCc4ny+RfTk2bGwXT2YwVa5g6cDiXNVqXQ8Aj8262S6cc9d6GDmE35ctQc3kgw
HpIFAjxdcQ3zSmEmwA4i5XaC8YeftJffWt+ScJ1M+T/fnqCtQS8+aqCuSzrr5Lh+u9Khl/wBiuur
mjD+gMLrZo+sr6DT948OG6loD8nAtLLr15KS18TmUS2PgBhizPGWeOk1GOOQj+EFfXeYgt3q5nsd
8oFtRxMh9mkOTY/8n4ctruPmhfgeUKwJ+AXeRGEOr99zysUKXAE++Nkha+Op8vzHWjuB8uKlfjd2
rkyYVzX3PLa17CsaHkNHdvTiJqbQD/Zqf7vBhPb2pG4c/S3xm/+ZIBM4vw2NjVLeJ7DYgLb1JDkP
YL1pBl5hq6hloQhyvKrmmTggaNSp3D3wJm+4mFa2HFzv/naGOvDJrC1hXcN0CwohFNFcrmhcaKK7
sxx21ZzIu9ie6uV1WFqCRN00Zfe9+U3a+Aww8CxMoLtwOZaI6cvsSydaW2tsAvkYFxHC9M8XIf7b
e+fpIDbVsqYpqpwZjJcBsRl45jx7wkDpkv9xYZ4rxJgkDQskfsmFmTBy2e8yDsxZhrrafsB7mquj
eaku98PRMK7pRuDhWBsQvoVIis3zIdgor7wOmk3qXAxeaejBWxXhDRJ33Y3SgKNxRtXuMvjfUWXz
lNg2lXfdavcAWFaPpz8zSJu7FTTPKQmCbpghxw8x7BTxTIK9auUN5uNw8uYR4pcOI3TSuZEPqcfA
m1+vFaE48rlQBWKi5PhsS34kOxIv+rIqWNFJcPkF5OLEsUdlDQLBCYmXay3e5ZYApygzkEAh9p/U
6KALrJPGAB/u+EHhuug0aVCDRK9gxDoIhLrTfBzu8oNX5gV8CkYSec0TwbISpRorwT0gbL313xhg
vwVkEv5wVKLC4L+a+OZD0f92x5qdSHbpX/4aVMFgidjfUOXiND2zXoAcTNUZog8YiHoHhvLKXyqG
WHDjLXZs7oc94NXrkEEjz4OqDJ7dA63yuwnygsXUjHzvGPHJ5zAjYSU+8WwrEonhwlL7NL6yT4qL
iJGPA0SWAVQMNGgMACwUnGdJYo5ygdsnbqcY1DVoU581Jy+LchuGoWdOfTIZflFL/8RhGvVcStnV
LUeJz6Y0dVDjgomHFiEC7XHj/n6tofZgld5lGGkzbn7cPWfd8bDmYhUad2HedtGIsYDN1R9nuie7
gpTvbWXGQm77MdD13znxJZKiRVy5JU/8Np7d/p0uKi8A584DjhB0buVM+aiuMwcdBZNRq3oJhScI
9xNolyPCXJDHxdPejKhWEa8t9a6VRM6NBteZy/RRPXYOJ1RtspU53WvdIQzfBC3yk7NEos6V479X
WtAhqoejPNT0oJeCMmpm6qUgkHq229DGB1BXL17WqXo8DKgmOfmsixMi7p2Wd0PtXzJWIJASfvI8
OyT5no/jBJ26FzfShPlB1wJpMUjdZzIegq1W1hMJRsaK6CPJpoOLsn9TeN+57ydWApWegbNZs5H0
DFJ1IyDnLaW4p1UjZ3eH37SJCIUE7K0OuNEV7N0TTai/twnJf9ZGyE5A5qtPs/WNtXY9d6UwQ6ZF
dFsG7ltDiqA5NmwZ/DZxqE0vDJGylfYXIrqW+xIlTgAJgE4pFVqRdQ/81VGChx2VjgnHqvUjbLr8
Kq7dGJgmErxDsWYGO1N+RMV7jqCk0KLV0P8WkyffVN3xIBzBfwcOJQKNIv34ABwJX7xOoazQpEgn
QgLsIhFvqdoCMDzHFpBhiWs+dbnFhyLPlLpuqoao5JP5qqyQJtlWhj/OK1XgHzMlrfj/tRHkyC4F
murxcnyM9RzXiUaC8ZBC2j22QDhor5S8zj+KHSgqB1UYMzC1BQMXv3WToI3FiFRuEe8W9DybxvPU
jbYLujEknTLK6DtuwZeeSuCwsXVrw7hY7v72x5Py+y4UJRsvFVgop9vNQRGj3ybRt/h518Rw3Lsm
MMzhak+XnpY1RCOzEqX+IYlvJbLHws//lcw+TmIgsZtXFtsDZMvNttLqmZ0gjPSJt/5BjCStA/NP
e1/zj6xMWdujfCwt3MwdrHGV894MwU/cDR110RKGwuyQkLmgMt7SG5tfx/wmO1yjOvUbbOsq2d23
QVram/chaL9XlDpZK4D/1plTu7GXnC387Pwa+LZkOwdIPQYguO6uFrryBov00Zwkzgc5/VVaI1ey
U3wKXVbXvWDSLP2kTJAGVkOCwwJeirUivZxm0rdSsaGxT/foOqpAkZ+6Wo1kerJ6C2gVLRtNTiGP
ADIRleHudzayYkp6qYXUJYYD8EKWBK1v4g9yQz6HPMt9qO4Txzxg3elPyiW3f2AAUXRZ17HlHRrW
+ZaQ5/RiuvEiEnKAEgfV4D77T3eyXFpsAdmuIJNQr3nea+51P5C6FLwDstjadpVE9B39lcuFD7OM
ZPWgPX6vXwtn0wV90+xYqZMg/I8GR6zk3JStn1MOUrgOaMOMlgAUHTyuTrg8A4C6tprrIXoDPPnC
hCM+QPVhHVkKxmKFFTw3k3EP05Mot3nMebMrQiZBpYjhhn7Phl6nBYxFfg7fNJbcODGSe+9TYFTB
6GondkmO82H5oE5tU/uZ4TO+0NB6prROaAUiC77mJ33/TABftr68f7PKS5Y1EnzxFXqmC+6AZYYW
LL9hU9OBQe26xM4Qwa9/qMVAeeqoGhPaEsGG1x/ioIVINe4iH9rJC230RyySvtWSN6iQMGfRg5i/
R8e8FafqXTEUSQAI3hjBT+JVAdT6mWa1PV9udOXgpn3PBuEinepjMeEbQPjRDBpnd5GGkGDIJ6oi
JxdgisiaKMhSgO56EoQ8/C4oTOQ7rcSAdRnuYkIZBHyXogykHlNfvyWHan3wDhQxAeqCUzb4sjXS
ezrMf90A6Xb+mcWXyAkrxTyp6IhEaoqrJAEtmYZ79XLXXeKvcUpBsXbAdWnEkoD9GTuIux1t7Ksb
W3VJXC7eAxEEVwQKvqBmdwdML2XmqAzgeuxeGpTggug/1AR11K5xu19o9ubNGx7EfX3WSSAs+5Lg
7D3yGtMhVaMbmTySkcCpP7q7fe3TO0tjMYaZE+KZl9FzhXpSPUdzCmlDKi/nRrAC7VKs0TJ7UXvY
sJeXsF4RFLslsiF8wnHnE38mFZivL/+LZgVCK8lH1NZjJdm4Vfvwc6VMG3i8AWVAuVn5/IjB29R7
WWRPtFIS7f583wG2mc2CKX/lzUtZw8raDNPh+FCJ3+zsFVP0PpAOmXqHxlwNxxrNeJqFwnP+N7tg
jKMsbYQp7WljGhmiPniPs9N8p+Gal4WLPBf0Q011sUSR0yBn4hU2jfu9DJ1JrBgU1q9A8JaAOtYg
xbDLzE5wcbnbQ9GCnNNmWMTVEGMjGe7QoJKBU4fTrXwhw31Jmb9JfWNaMYJvfspVoJk3Ev/zzJFm
02juIsVnQp66oRYvQoUVqRc7iN3Kumgmzl25uJjFEIU/t7o1jEE1PGvnQqZx9K9MZRScspaMyF6/
Z6d6ajA/ukv0ubNPwQpQYjpiFypalZ9lp6R6KgFeDEr93agG26UV/ZUAUdr5SvJ9KagDrJqmbGtf
+QxrRTQ6Rf2lPAARQ0+lrmcZvbbPn0ijdEy6zdai9eWnUjBX+QyvApAEjnjOYFjm7HEUfW0HpE99
ckX7BEmFio2hhaF6+B4koaHH0Ewgl5apd867R3ml7VIAUQBJCEKGVunkcDyNkuCp3PqbUPsm9lWu
64fxjMREPYFv0tLboqpffEwvZ3kvid/rH18NQubkHxCitMD2mQd7zsetT2DwuzkdXWpcy9GH9Y8W
7fAN/hE7awFhnZNQ218Y1gHuTL8akbm5e0F89A1L4Zk6Z0Vz1HiTYDslBtSEoBwp4g82oVXzgkEr
7gcJ3vipmKrAtx4myNsOQDrKldLXbOuHAvKjyxm7gthVBNMquLMJWplM9JvaXPtvua//CiNtWEW1
oNAuuZWTzHLVyGDBxC4Ixgo+A+tvaenSJYb4HMUUbyeBj+hLm6xClXmhQxq4rpbOsNzZPsUxZHYg
c4LeWiwXRb5upArwpAvYXdDz0CKQNPUb8q9FbtqrfmqhAHP68bwvMlW2+US2C3LXXL2R1mHPbS4Z
gg8rF4ZcIxOgsPxBK/TPfgxPN3b7vGXF+Fp+bgBzQVa/Cc0J6mlc0Y3uH5tXLLD+wV510MCwf+WS
yPHiYJjW77uVQRixzA1ZK5/Ezaie8WbczJZk3LprCoQHJ6txV9ziAXoh3acfIiTksshlDOYG6voF
rXd4dYSoB0aRp53fTjZeouJEbHweV3Qn/CdGuX6h6lUvHgONGT9dVfvMAhJ5iff0v4LTOVckxfOn
tIUuUKQIjAEzOsGQN3zDr0T1PWJEwIWiBYzD5gkYd7QiJyTE18ELFyqCu672b969oOhkGJVw6Mtj
/0jNy6ApXwFnUjOpiiFrSbH9h2BRdwDW43q1vVXF/j2xnAZ37FSk4HhwXGEvwisW4pzniMqotNxt
xx+hMtPoPHwbNLWi3UkHRNKXRaKrPJ5wjfZcq1bfUM+0EoZ8h7F94BhJJm2tNGTDMtSaSUba2s8V
U1ilNi5VtG8V5XO6HCUE5Ri7/cGRC+9giqKzr4JQn4C/2l6h9RNDCe7pu1Xq1DvUCXGSv5awUARt
OmtPQT3xfzB7LRp6TyEPG+0zyK488uLK6pdaCpGQjX7pfT81QJhAfO+JX6bma1nKBbg1jLrRUyKA
AJ8+r83HgRQ296ormXsIr+JgMGfVx9yJpGaQU5XtUh/7U9yrCn9DHTeeY+JPLxZbovD9Tf7oBlm1
Gl4qaZ3duxD8qWTFNtYJIWoV5XpZTpaK+UXLjHTs+PgK23smWIW9mQyjq9eA8uQhBeAAcbQ0L27x
QES7BO6nGA4nNh1Cc5qdbsFwne+lqzLb92XmrVHgpr6G2dbpCcWCd5HV8SBaX1No1kc02RjazVhr
5IWBVRSYV5R3LQT9gOZK7J+kl7oKrylK82pWUtF6iNkh0WXnWiBrytRvvHeMX7KjYCEFHl4Gs71Z
4rN/baotWcpvAiKFn0wQZ27A9lyqjAUst8bGIDas7usMGGRkOWJX1iHhBVDucHfJ2DjhVWb+l1oC
7GBk8CkXFbdUW1q/2owZhJF9lvfyudeW1p327+VyDr4YK9PDC3wo00TeFOLt2QlVRhpvTR0iRrHq
2CELqBuzkx0QmeK3qaN59auWTjlC0kgxKdx824RFv8USa2w56sHm5B/JfgNP158VBU6aWHeZVVxY
5p2TdJFrLA3fZg37Ww4rredgZGkP3Z+ivSKnLL6w1IKW5mum34h07bCRX/ejSiLt0LcoBFTATLS7
JUzgYsimuVYhLszTRpnbeNP8fGRSEdutR18BmPbSJYPlVFud1R6p6YPotrNanZs1iHd7ZDjPZ1WV
zvs0m9QFqYzVWOTIQ+kj+RE0jW+jZIzfRskvYj0p/W6cg6VMIgq164lYtjaXBGw6gaeH2i+ubyCE
PzPNABjPP5SnEHMXzDF8MfajRsK3Rf7ZLKLQa11Mc0rFrJTMYMcjHvDljW/YxBcNGU+uoXpZmwtD
r94HMLcYyzFwEJrTs4nVWUeGPSanbBJh0TwTaUjQtL/1PjpUeBix0mxI6L85uxASZZ5FN/8QTfgV
h0U+Dj0aKTA569+ObgrPpebWhdigGVOnBOPAMX2pFWtICProokprT2P1OvddRxgUSRntiCY8w2N2
jH1Rd5IrinsnsIgaKLuI6cGV/lmdnMk74biLGiXYkRqdgFPksx2xkl248nw2QQQl20R/I4HFUtbE
qf/kIHwSLMzD+jrnUFIenllCNxHiSunAu3lznR+nPiwxpJQTAgayQ6X8/lLONh/i09jp/oypeeYv
n13ksqIiUVzzJj54H+CPDchtkiB70zaLbAGez0Nfe5B+b1YS8eTpe0uq2we+QOm+3bHb/5phAuWI
ILP/3fwuVf1wdbLrPp2sBAOYZGd7WvMk8SK9kk9bhk2pPpMUfRGSKXs//dWKBTBXf610ZzqEXs+u
5GYFxkxTobfDrRfThjIAxmneDdX2urcEZubV3Hb4vqkfG5fyFOnLs85HUPb4gf5j77CVxVHrJbej
atRjXBcGzoLJk6+vg/tCiP4r4/OtQQ+HzS1lSMGKT+KQnpc6lpQ/F7wCBEigKjC79AtTnaWxURgR
PWZBbss+//Mli1jLl2fBwh4IAUiqAD7isUYyWDxUP+hPWUuVkUplonLPIO1zwLHtKNusdhAmyxSP
6kWYDSqieUNpFd8tTYKo8Hi1Q5SoE1Wn2uvOWPxDJSDiEvhu8BbFhkMarfzjmtJPlj70ZZUgYUo2
arH5DhfEdkAlRcuO6DJw8dMqlu+/95fOBVgMRS3dn43D371ZJEJGSQbltQaM+M0rJK6JCqVvwLgg
9fCcFCWCZtN7YbGRpXUS7Z3VV56n8qtdjLBC5IY0PKLRq2pco8RCdtzmGZsZNvUo/LdxMACsrmXf
dHkyvkB59A15Hve6L473GNlhK5Gzk/0JujVf3mWXGmwrKS4HfpYuNax8//uwBR/7raHASoL3C4IL
8J7y6bC7vaetmQDiqEHS05SWtk9uPBqqsky+KKv2l/Cv6axMUXtuNDkGkqi2qcZs3AStoxJD016K
pWTMNbCUq2v2LzDTDQDA0yvhRGMF9s2rPhD/LVesEWVSgQpMBE4Lvil6w8R1kx2tnIhCjdhs9r5a
xeXFUE67jDW9xTvv4MR1sXiIXoksXfNG21NcQScy+fJky+YnoKEaxQZX7tK35whxDtSOB4E1Do4U
oU+teh1tdIaZIuq773E8x/Iu0RBnC0YXb7/N14Zue6TL+HelZnlSdOQ53D+LTqndEsAnJvaFmkB3
Z+cQrPlVhdm15/mhXNTec/vnowRf7nfQn/HuDlhNfbhq1rMX0o/R8x1OINfYRE3HUYItYm7xZtTC
SKVI6J6ZJiKijNB3sbcx2sPldHYA0s58WBcojXEeElYC9RIWn1FoO4/bT1NIDgpriuClGlp9iCJ8
9sjnt+Ml6XX+VrKn7/+H+Z2nltDT6yeU16EnAIhFfIzv3cexKxsWGxo63dRzoBprg8YTw5TWKkBx
ZA+pB7yCMEe96a8DiPvx6ChTzI+S0RT4JeqpmX5NKaVrkwWQAP3S30zVNsPYFE8xSRaODCl5eaB0
nE8li+zZzCwyukeSmNRQeKvXP/Fj5a0R5TGsLuQibEEXOcW6w8ikWpZYaxozGgHzgliktbASEtjZ
2bnoDaa3bhX/OLRvTcEthHpMV8QBXgCW6c5Y8Y5MGwzS51tHrIS5oK9kx4FO/HgePLD99CsgW4C/
9Vo/XPGEpf6uv7qbhEPBKsk+nHnZcKpi1qb/sCPUZ5gAEYd/oIoWblc5G/zy3DZ1yjgHf3rD+du5
WE48T8yDB/AL4gUAuGqAfpoAsIKjuzZUl5V2G8WudfDEh85q7WGiueQzzVr46KCLstodDvzB2aUK
CkdjVU29BkRJuwjlUSMuouQfixCngdPVG0PTvnYOfGWMy1ZEiG0SxSJber40ESjge48D6afVW19l
27pvZRmvkHouJi7Mffg/br2AILtC6avu+1iYFyDpFG19Ve90Hn0hKN/uYxChIPv5Jys3u3o2J8Vt
CUVJXcWUIu4azuyO3hzrDcTBxxGRQAs9tNzcmC8JvYPnO4kUsXkbWtxf40IYxQGZ+WidSUdWIkBg
lNCbEah5APFV2tl6IzQEXLVZydC4DOZTDrkaibcBz/xrKvz0+Ya7X+GFEbBf+RTzMcCTKBHz6cnp
bKspvhsXNjQejLHUWwAWzAalftyf89KS6NgWZoRcsv/aNgT0E2zFPaCpZjSWzIcZsOZ6mdnnuzon
Wlisw7I5iBZuLujVc+nc1voTpVLGFxWURJ44LX6p6LBiw8mv3phUty/190yohqk+RXO5aX1sqzS6
rqIwxylnSWygtgAbMs3Pcvv5aF/j/FauyvQPMYqn89IPYzhQAz5bsPJeZVogRRbOjRgGobV5gVrf
LkCc4uoA6gpXp6PTrq81hCy12qMW8Q0IGKvdfJrRiYv3R0A92Zb4/gohm7KUKweZL4FDG4OXWNav
nqUJ9bXDmekwOv/Q1SjuUZzjUppxdHyjud51AKZYcvzlaU8M+odZt9frmKldqvJAXFEzkNtELE8q
c/RjRCKiUvu2msizzfT+hn/wWFtBCihcFBsVqCtcco16lDEz40KSAhLUShaOks3gcXkqijobRIP3
PF59LIpWgXzrkfd1xBcZ2c+nt7r78vJhbG57KX8PCG1jux932+4l5Zg5bOshsPZTCe/sFBbgC06U
+XCVsU8r3KLsW7YiGYytyKjGCLYmrCaFlnP65zoDOhprJnkvf9KKO1qdUm+4QeIjm/2wNCMYh/VJ
NLD9kuiOSXuEce3zl7M9YuBx3PglctgGGCXgz/PWi3XLaxj9N+Gu7VJyuA6Cv97VM7r8RZXNg+G2
nR5x/Wo64dnoY+MZ9SNUQSKcEIVTdnoHLxfOpi48l1+tWjxs98ctsFBuZ1kpsqXyzw+5+dURxijd
EUA3z/M+dG5Aj2pyof8xKUTAWAO8Npfvo6oEqzYRah4ZucSwlVRljg7cZ7+l1wYfpL39ROjGxL3b
ftdzH/+OKQ/lEq/EyT6F9dJ1NQPr58NSrKuKnHVPDi9Fn0gyD5EwU0pKRDnwtTSe0156huEFgL9F
kBaqoFhsdb4JN1VMPZxXHy04nWfeYCXh73WNcp1WUbRcE660DXK5jt2H1PkDKnYsoE/kanAD+ni7
OCkMlrmTOOhUHtuCyoN0UZ3B8YAX1ixzwqLNa4mCTTz/PoIfDhusW54WmCap4t207osH7XU4M+9x
C/pvH6BtANjO8bF1Ra4KnpUCw2Gh38Az2xvIXGIH+F9DYTCgjtC1QlWWOgKn9fO1XdT6FPtIzlL1
NNfQ+fcm+verwf5TpDtN/R7DpvLjo3XkhDCUbItTfYeFegkJF6eOlbzO/kOsF0Vpk9nYTDXxn9ML
/fffiOw/h0FnvzVi6jKN3+KUHsec9wSGaOWVNzqJIA7B+nfuUFPYM5AcdfVlPBm7INXEKGlzT9OU
61Zb6oQK14xVCAY2ygp1mg7qdlWWpw3iKybLzy3EVY29z9L+REiC0+k2B0Cj+jznDMnyYudg+r7S
eUrkKqcCM0k2+gnbqbDT8Xh+m94pRH6eZzIqjw3czqQZdjxy3keVwZcz5IVLceowQviXC8+Du5nS
6zprEDT/h0UNTg2D5C3xl/QJ/gSAUUehuFiM/3oHLSDMHfhh5TiqHt9+7k7tf1hLOc7CfKELFZwF
ZxXBaQky2uGVj7A5e6b5R8MCoGxiKDXlv8enYiaDcQd9v6s3exqzkECcXEH37c7hq+3IVsaWYb8m
R8tFjcFVWEqPV9xp9lE5Uxd8yEUEJic/gStRL2wQL6/Nl3UUTUkm1hkJ42ElQJC2oeYy3EqMKWyw
YQa9pi8MYGNlf1WC2QqXY+H9tsLBpTO6XMshPQRgPRTI9ukYh3MUuHn3G9UY1jKWjQRcGHUJNVld
99Q2ic6Kr6N1/iRwBPiSivPUwpQ8aX3cLAf3bTq6Ohz2+qaYBoquBqJatU1c2P361uBooaYNVsir
bKXq+eDltxdZ5AduZhveqMVa7xGahgEcQkHvina1JDV4ZNeeWCpoJii1jWLBKnIEVWigKSWF4qly
nrwuK2xpBS6SwDfouRVcoTOEGk6wBITaLwp7KMnB/HTMvRZYZZAIs3ZYxj6kXPJ+rPNP6nXdmo8x
k0rIi84nZ2wgxv/HH3ZJy2J656CdrgzyAbeLFVFrA5GkEI9uWu9JIRG14u9kuDOxSag+Brg4Fulr
SANGxF5Bf7R5snoB3aYjpO6UJR18PprBQ1iqMEpkUH1mf3cf6PE/mFJAYLqEALAJfpUCXg0r9fa8
tlkga7y8k26qmOsZI8+j7qN7SMwGixKGFll4Xr7OWJwUhCvuKvLSGnS0te6eQdb9UsQs1kdZplcs
/8ct1QmeJR7GJQEaOlXLW5B1OLx1gkxYMchWr18IDbMVLA10B81C2KAb+ByqJlwEdNg4Rso+slUj
iRW8xLzpxW8kQ2h24cranQPByEpdy2URAOvWjJ9MB1nScv0kqv5wI07Z2N5qaOfuRH6b7unFxyLO
9Tgedn7LCeu3v7VVnobKRZiyuO1h7oJW0n2QuPy+rhIuXCraxFZZM33WfHszLycdcCW+FvMPuCrX
b1YmGqFSvUy0ppRKEJbhKuHx+SpUDqCixtvcKz5GMU2tpxPmUn3bfuzqITtbcyiNwn98oXjD4I5+
Y/NSkkxMvkJKBoV5QIv1tqGt0lezKRZy8EvXt/wWGqsJAPjXkXKvvvnZDIh7DeBYgWKGkhiC/fsR
r0YhRmbddUfTU69DcYDP+HOEMisgftaMErBJ5Phwr1tXDQlgTK5LDt+LbGXn7V4PcoGHK6iWBSJk
iQzoa13QK54zONzXYPAKKaM4Wm4Ie/8cXFUK0YyDTaFCEHBCXZ9mFCEWpyhmHAm1doAfBmL5vCuu
4XBQ0K/7Mi9sXfujpdyst/4RC66nTbWlqMy7h7wcsf0s4/VWE0WOIZ1FeqjCZwRHXcnboqBPHrSV
lGkX+4Bk/lR2n869QNG3H5v0TcSol9X7dXvPc/ZEDOWe8ZX/sJrlBjJYXBTvHHbjbV9Oieb3k4Jg
UQJ1AiHL7PiTH52KflZh0bobIvjAMWgchV0t72EjOp57juCj0L8k1Cf5gu+ZHa4axoSzh8FvCNuL
Bic9bXGJ9qdgsAPqRlDwxbhoPI96S7lVK/TjiyaO6vLRj73k2MJjhhyITjopsnWBRdh+j2kl1kPV
yzKfIrRPucotu/8Agirh7dzonPrlSPpETxlXMlkLhmI0/tbwm3+7nNDJdtz2ioxqM8n4wOInsUiW
dthhRpFPGUi++hNsJFsRlCL6laD82VINdRORjtqwR+oFkMW3yGDn4akcA1uj10lh3caz6DFbmmp0
hAR7UKJWYS1D4TgUS1WfWKOXOHa+AH+LHSX5Z7pQ9aGra5WN5owSU/CVKGzVk5Xr0jSNgWb3OXT3
U40U8OqoewHrEF31mhyN1lC88LOiUgAtiyjCNmQLNPpTx4uhDgk+IXSUqM0OY15I5u0iX+H2SP9V
vrvnGvr8GvO6a5BTnXsjfZWUG7AYCdI2KqsOI9PxS91Pdy5P337X1uW1OiIcCABefGY1zDOB1Xtj
/R+1O8vFj18nev4z5LLHqgpl6sc5lKRusq9ClvMaPBvOmu4iEk3gyT3kzBAAnt//S0GtVpKkpWug
ranLwkQEc/IKjO45eQ75iFTzrS1h2Z5QAMtmbFGOfrSkQn4cZKuWQ6Yogr6kf+Bw8slXwprBfdj4
XUGXBiHovHlUZusf//8CGcUMO9zaJ1zWu8wx4nvK6/cKPw13JdUYWikLOruDGT0W88k4z781nscp
rd+xQTwpTdANW6ORYOt7PiSSjt01SHQAgPNra9gH2MEkbKKqiMqcbCJuesXCU8pCaqwUGNhAgRQy
ScQUderx0SNg4i5wt0jTp4ZGqlw3NQkBi8qQZSPsNukgOcezDH+3JKlYdesw2qvPjvkTJcsMZ/Dq
MXiyf0eFiUATGHCf0mCEvXJmTPH+JwJf2Qr3z55E1BOY39fVomcchUUr0nPdYcUHlEcQjwg1lC5z
dz1D/u7KS0C9cdzOgzCB8oznuiYsBpFLWYwh6SDeCF5E6rDNiUo3SJ/HrQ1TgsYZDEoV/ffCJG9f
mo3O7VRlDqb7Zqu1jD/bCgbWOO5Bc+eclD9RBmNURgLVmshMQZfD2YDeol3IbQ8xye5t3pZNm6/D
65TOzeZDBzgouyf+6zpKVz+ZZaAZrzQOUymKsmYgdtTcVMkUzBlRWILcvaYb+n3Y4Wiuq0pwrg2O
JZPYI+CjOf6SZx/+pIUTzAnZuabnqSQ3tDk+6ZsMA08LEeC6ffFuhWzwZ1mzvI/VgEzkWJlCAUPh
tyukotiyKx5QKzLeLx9K+sLT/81X5Z7/nVoy/dtIJSe3AY5WlyOlhcyOybblQo19XGBYQfl7e3UF
i8pmaIN1d+toSQ3MhnxYclzPa4aBkcSsLVg+pK/SJP0QJ4dWhDBRKY6ES1M2WK62VpSFT7dbtVIB
KSkccGISdWsgfE9gP3elOycyP0mxpujynRZA5UtWTlNNP8MK7ZW4SBPbxY7C2OIPV55vb0L27T0Q
PqsaAzzeMEryW1kUOJpjdSPNIxraxnb5tMnIVUE8QAf6s4HSkTE2kjQj5M5xcQ0xwwZelCvnZ583
A5FPAwr5WG/q0XBkM2GcxL8FNWLSbk6cYmJ6Jbe7UiYsQg63iA1ehAkOFy8mKF6G3in4J2Hx/Mil
hhEFeCAr4oezfDuix2MDpAd01QkiB0XQ/V0582XkYFh4XAn5KnyIhtAUGkp9rEpZBtveQiT7jiDn
uCrygsCTX8zZQ1byZwbtVyDqP8SZBMGbhyYxKFNxdZJC0m0C2f8I2VRcNy70ZGFbVGgnXq3QK+nv
BG5mWsE5Hpordrfxk+oQS9LzI2esbsBDdJXiRSdY9kU60gRJK15+ujwAdbtOGDId4nJnOuW5vgk6
ej2QPoNSuvSMUR3lYKMS04E0o8nB4bp175K3JlPYy0Msy2ek2/3WZwmRXK5oUSckST/CdEH5wck2
AFKjyxs0ZYpoUuuik2mQMcZ7os/wkzeMHRAzH3VlymK98qRSPC+Xi+JV+5mIneS23sFbrEe5z4rC
/Lj6jr3R/no+spxD9vurL9UIZ2VZ0QH1XFg4bDenBV6hrVVpoSMmVKry0/dkwlic5cUal/KkmBp1
3L+1KZ3PYsjK2Cp5Wak834zFvfk1wtVLwzQiIuORi1AVKCooxgjAefOkytD2VsWQeQWhIF0C+R4V
V7u2TP2R/ukpzId6d/tEVRbvwud8iazEW8hDGT1sT/GamHkJjwzeQ60xMQ6+OX5K1u/b3JQdqa3v
d6I/zjxnAPIscPsu+QVigq6dSBybTfOdi1K9cybycH1OeeWQBJu7kNn5Pe8GXn1nyCXwZznhXtTC
f697R3urRug74+6ZYFcisPCc86DKXCEKQEaPjwR9kJYsCFebdtiOB/o9xqTnH018VvqSww+TXDw3
GwPexBGFYCuxY0nXmgByf3LP2GvDP3EZ7+ryTWT+dexfeks2KiY2uB9mncOv766aDeg5pCJuVGd3
Zz9Coie+fDpNTjxA/gB6vwWpvYbqPxhq/QNg8PVWwGxRVkHZOQx3RqAks7Q8YI5Zt77PpaHONq97
mliEpg0/rAahu37XTWhUOVghu0L4qQLRUm2HICNB6puyPelfwJx54yTrTj+n9fx946c5d2fsHAOn
IEGg7hgDxTWxWamPxT9XH9W3TpcQs8GjI8dHczpH/MAxitI3hffjaWieADxAWy7ZQxypoEX1PsU9
r9huX+fPOviidAc0vVL+CJXYl+mQTlZMz7eP4dRL8wWpbVSz2KLmkiUCkDxD9oC6ZA2wwMQ2PYun
L6UOFX43Y9rmfslou6KLC99m+ZDl3buBWrDXeuMmg+LH+9WkwXZ6jI55/vgdxUtRcQH4COtgIWMK
/xkilI2D1ydB7jDzO1VxZokE8vbAe7+zRsVrOXdkW4Bao1rr4VoJ1kXeb69OojqrNtCvV7gRXX59
Qly+8B+pRcdfIKv7pGOvddirih4kVjTjwAEQtvzaqCOMMxD7bfFua0rOzPWECOy7lcH9kLu3aP+b
1E1cLG7FmCOPp3eIeWtyStKEDiEXhNRYEdh4Aa4w5C6s6fsecGr3fFMkngBggz33zAXkJgaKxeAZ
GWMJQQBEoXExurtH/lHiwZCCfAQo00myrB2p2VE2H4rmb1YM+1r/5FsLi2lIf+RE4C1R7RM8uZo8
LXlugy7wkXTHJQ61RDQkYlWcP8DMH5qgJXy//y7KMLxIgtnCFdSLyVOY9sRpoNumQkGjMzDTyoGe
i4fexpbIHc1nE9DbNlWhhQWzMKzFHgaTq6b/nyA3lZniMdLTwl74+j6w3r2UQTagvakDNgOX2bh1
7M13+2SSVShtYxtqtU2S6sDRHZTVHA97C5f4ZjYCkg2/N213LAwp0/A+3SFfiXdhHuguYH8zlDze
QVZD07V2MEAa2W2vaGEPx6B4kjL4dAS6vXcPfRRS23mX6l7fOY2OyGgY1LEgLnhI2Jgvh3oX8woE
e0W60VLd+LsoJKOGpm56IjMVKv/2Sjm9nJQTaiUsD3/wGNnMy0zPlyZ0+sAbsPw6hjTzWiUYVjPF
MvGnhOxrmwGSRF3rJpT/EXerb7i1HYBbnWfZ4f63+dqzG2okuVHEDUV6/9fIW7NrvqqsFM0G+vsa
ccWkdVy6vKltCiRt6n6lIPcFdVaSBvoSfv7hHFRo8LqeXJwVJ+eWuuXtI238b4Y8SaDt/iSDTIh8
yut++gsZQQV/6VoeG7O/l1grScVHJMJSxDQs2xyJw7TLAsjHyLREKDF5cktjikiyxtx4yOqanBz/
mHbv6uPChcWUJ6fD5yK0/AjU3Gfk9/XR0Ji+5uRVtg9s0vomKZs0TRaR3JkmFFdgH/KYQjVFYvH+
2bfr+cu02k0iRY5ecM/SHOsFrL8VQjrAKFH19W8A4apaNNGxjn5YS+xO8XKTLOBbyJoWWZFPAW6o
UUjEP4wAFggVwQ5lMMoH3BT7eZhJVwsITQN1a3tRUMN52JZU4zR12tEs0LY+g2H02CIe0QwNOjen
pfgT41KVeyyceuvhW+EmG9y8kc3WL/kqYYBCg9k8LV9qBiadA1MYCjm7wuy0qeHrhicZuarI4mz0
VD1cz2ML1/RvAoNFYQaBcKOt7JENTsKmVZMNLMIrO8tIeHap3b2SbEe36JDzjL2g2R9Fsy7iYBJ9
G1LSSISYOGyJ9f/G0zJ1Su3bBVIicEBcKs442aupxYlfEiGjctQqvxntd/iTiUFY72VcOE/BYV63
qvOA1fwm9e6H1og/sggn7dnIWHmrGU2bK+ppSUjD8I3yByI85ob3jbGhLO+BFS3rU39KkNjz7k2b
G3Ww+KTL2ccEZfYKNbhsV3O3klZZ8T1J6HxC35Jy5Gu447x3FUkHiI3aBeNYKZPcjLn3IbCzmxLg
TjZEdjdPB71+b0X+Oukgtq0mAYbpw0Era3GFwH77Cu1UXZoZpeI81L+h2gIYe2ZqYw883ZZr+Yvi
EJjygYotxx+sT5Iqo1uKTzzGUO63NpTs4d79X4GRro3wK3xRlIS16lqQFEM6Fcv9vQbVUWsitnZr
bYvFiJR60BD05rM+CfTXvBqPUy1QjOmYPYGVX3miOMgkpAyUCKeFDG+yaGOD07F98CzE7FJ9SSMz
aqYPyWHlAzGRAtqzwImTHqiBk5bTLaGyns+4uS0oHFMHeGtb5nfRd/88g7Gei/Vyy8W/ZNYp/Ffx
8GtOhZmwXZJ9Ba56h4aAyANQxOFQj8KjCIdnbWbANy96E88OfrXnZPVHpjYljZ1PynYxvdBgwS/X
SKkF01goAu/HKiTlJjVjc4Saw6EkkP4MXlK5/h0cAOeLg2IufIZeMhkPlLc7yMFVGQc8Pprm/KnU
18XkOR8gu4PP9WbmeS4Cff3ZpR1ciwzRsEsMDkvLWbwK7FpjC0MM2mJRTIoKwVLaEMFsLmm17uA7
T6XxzczIs2a+D0aJb6WfGFRUMaNKxtaJ573OZxKUGAnRklU4QvWo5eskk0FUeX3ZtSL39w7VYFCF
BkGSNQf2+yY78Ez9YEhVYmgXhw2xNAj1Emfvyr/KrzAEitvmP0RLZUYir7RJ4hn3BJx/xUR9RlaJ
7gBCzJlk3MajlLGiTlPL+DwLvNlag8vT4JUQcgrZ8Je3C0l3vanxGYM8DvpGbJiKODKfJFSoMRHh
1dvbZuZJ8Mx6o6z8zXQSDhLDG1pD0D6pUHiMU/c5ixa0Bu3/bGqn0PEkfYxIkzJgAbSYK4gGLznw
8m2nmVw/zDXPM9JtRbxV70hzQesrukSa+onRBV7WGB30hXtkHu+QULbTZ3D08bpjmdB4MOT4J3vl
Njg27lE2fMJRkcrkbrEAP0e9962wiHgK6vnDo//HG71KJkhsOY8VhuLZCMdHPB+fAb7hblJXmm0E
3mJSRY8A4+Saq0bCvSsWOB7+e+tUPh0bFMDC2lqfXqWTQewUtb86W63BGoKlR/6+14SZWWx+/5dQ
glc437VWfnEY1YsjJy7BcJNoVIozyeYT0CJWzK+/vzejbT7kxQJyHjtStrSi9DSgsoZUgBlpFZ4o
8r7uGHGVPYtqQ6x3E7NJsTerghySDx3jjsg6BTz5iaXX6FEYeWM2NIIgs6wjbDYvGYQOPsphSi5l
nMzBXXNevCiJZ5rZ94yp3YRzZmFXOcNUaLwhNGOkzVTzz9oqZdUt015clLl0H8yT3RP9rZs5ejAV
krZLoOxvkGI6isTzEjhxh11oRyRMUQ05DJo/z5uKzj5HQ4i3uh4ZDU7eAniNA89mg8hJpFowD7L3
VUwrm0M6/yACGBP3nW/dUacmXjv6bS6hQLQ35s4TJDWmoRa6NowaZdPUtpRmILHH4wdFExG1sNxQ
lR/QgNgg6+W+M3NndlGM+EcZiXl895zQtG1wQrBq3BbCc6aj4kpaMuF1gYvj7NfswBSoUOUp4zSp
AE72zs+cEiFenKTCApPYAl5Diukrw9qY+3zTyJXqoIMv2Vt5Xt17xBPuRF/xHZtYK3JwSOJw8Lto
aUe0V1dkzo1Nr5gUszh5KZk7OX7IBOpK0kdwBomXOHXTHL5sRgN6WAnjh/9+L8IPIb7eaDoD496O
v8xTl/NBxi0Ss876DwuLwdUv7tneQgDkGneJWVavOOtG4nvSMzg9ytXHNeZ02UH3jE73jXYfxCt4
S4tTug0zu9DrDE07JZeN3h5FdP533EWvIQLErnTasuPZ4ShtS4Dlwcz3TIO1cWgSxS25STjSG2aU
2XpwD/6/l2RRJ1h0ZD+hYyeStrouQ61lSlx3X7NhYv3p7uQ8505E5jcPeMRJtObMT3ndu5G9x7rz
cQzLGfdZZiBFkLM92J83ky+Yrnu8xQVDZrqfhuivfUOOJnqfV1SudKZfJiBhhF/+XyAHpL2pThbp
uHQEwdgnoiC/756a/EfqyP1FCTFvQLXInRvUU+Fy/YgKfKztleu2gkXJvWRQUazqjRz3YDNITSXg
NBFcPleuCI9Gry5XXVnv4UidHeodqaBgwYbLKuQWdP6mGm62VwFkiA4HsXIK13dglRLdcLvIZo0R
djUjtxF0Pss7dA6APJFMdDBtBxizbkLMUbjG1rRK612K5t+shS5p+gouGv3Gv5z/mW+G0SLVCcc6
QPW302LqDuTLz7dWCsxuiMWa8CQi+JeIzxliYAzx8CeCwEAzaRT3Jqai2CWNPqVM+FujA542b900
IN1smcFQP9IrLAAhuVjJEfxTf9/vBWbKBKD2dOTN+49sfGuuSpyiGojh+pn/5GIDsnFD+s0e3Y2X
TTqNIwgH/w5MTzi3ujZ1MKClLM1Ij9CJ63/6I4xh8VSKw84GiKVprtDDuLwbrkyOnp+z5XEXGvZH
JCZFQHwrOa3CIwO/q5R35Y7v4wqgAOqJO0ZNWG7nidMRfbDdBkr+Kg+Z2PANYMPPATbwMt581+5e
F7NN8pNWzi5WGfOc5keGpjALoqs6zDMRAUCNSKoBJSki8bKG7yGOddv2CWLRLXDl7N38BFGp+wJq
IWkeN9x/hCVPCcuPKquooO7udJse6EvL51MtTbexi5njcWlw/rSjt8HGVDHw0kJb0Q3MST5JicoD
PwcQp96Ucncwu5gvpBiHB5lUdmhmcCSmlEwkNB8vqBrtlg7B+wpcvKLD2liHpUlPbXGgc0DOf0n9
PsDAWmXFrM7BM+IkA9NxwswFW8Ss+BvRSJEYmQicQdmV9MkeIDKfkedYldyLLS4vBZBhJjAjUwOb
SZMWpYIsEr0E05C26X0TUA4qcN3YQfQxFGXiWzAX/p6GNhQJrJLGZBQZ1sooeSYi7ndFGHFcTMKJ
qpz+8aJYHdGxuUHaa7551770PkV3nz0lLAFrqKkDrpeqI9EbXzKp2E8sTd4DenrswLWgeeDl3TCi
0cfjFacp7gfOBTvt0XOMI3qVEjXfK8IWfMhY9GZsL7ZX6VJ4+XV1kotIf6QP7rPLVomi0eLI+Zlu
lPoa9Nye9bKYFlPIL8R1QDsYaz2/PW1wXzZBi6s5uvSkQb/ttiSuxq9JZqZ0H2DaF0C+4g7fkLxY
iBz0fjFJAO72mtXcfURIu+HnpDNNb9glWC/0Ztjj4L6BieeQbOTjifv8JU+79ChDr4cSboD1v1wJ
vRnaXSnBZTLKW2R5GQMPSCquIMJxMP2QIWKWKLducPK/A/gKPOWVQbWYR5FZyWMgtExx1F7Jwkwc
KJ46EgsiI5LZCQVLOETEbQLRxQSIsA0hDFwCRGrSklruo+MCez7vUze+ceWg/O0ylq8ztsDCUokU
FOwyyQrJWOT2HWOr3xnktJ/9ulSfHjw0uaIMIa0Ck8SrVs4SwjHyQCpoDWT4Adq/nXMHvhE1CaV9
n57ZedhSOCY/ThK9bvHB1zvdLOedEPeNCm0OGOQ5ymXXyWHiI14M0YxXgtSsCniPumVi5X+XMhAe
OFY5G4482Eyy1/HmCVEuqOJOGM7S+edf2aicwZOO05fuUN6WOPBLYElcl2ZGUcDCjUpOaTcsx+OU
fq4x/nPAmhiy86/je3WaiPcUtuhQ+3Mda53xctNlcKv/mRJmNuTfAgDp+9vFkyS/LjKZvkw/P6df
Z4QDkSq+nZrGAETixEbn1OMTRyw6chsKZ9BQnTg/AmPuUF0ZQmbxsC5/4JIM2KNv2ymRAhvCK0+/
42j4xosGpTKV5IMMzfarlCP6GjHjv71KcLb9SqoD3OKteA5x0HHTS5Yhl4OzK+6xa3ZmrJMO0hG8
tcZ3jhNNPKQZiYtOeZhhnvM/m8Bc11+2k/VCx7Q0ev3lGRtp3Y9WcyNd4P2ioJ2uuYcwXVndmW+u
KEdZOuNZlJZi0F/NR4/SgQN3kRD4Rw8fucVR5Yz8QnBIfAG8iBv+tAs/hAN7NK2nqH/tzXhYoBSD
sJG0yfyek8jUwN9IT8FpPxI18/jbZnZw2sa6OBaxlYXxefcKSBAk8q3R8EjKVH6gZAW+87JJqNSK
+vaR3YDCDdlXezj8PAjx7WPh+sn3+CeOxaDW3q8FpzjlEO7FvhDqF/79mUNfgPiRwXkrlaAhKMDa
KV3Pco08gEcDF8FVICdsEDqnWE3zAT8kP2OMMuUZsYgEGElDajmRApQew6lS4vU+mLiJQIO2GGTn
aO4Ugk8VcXJOe1Djg2tPV95tABSTMvApVCQg7IsirxTE6sgAdcICpsKvqwr9vaKv9YxBBpk8YsIe
nc/mqRgGRmy1MCXP7O5g5lvvjYK2UoSK7Yqqg/y5bmyQcgF30z/oLtRy+6K6gHKQlisMTJMxQuKb
Duon29qLQyV0I2cpmNRpibvE4qqRzlsKMukdx7Y7IOaYiKy2Qq3gYi3B2zuqbdVcN7udbJCrTUbS
uctmzgtQJkQk5c5Gr/oEMSQeJjYW9rUdPFWjh2de7DM33+6/PRnjbHFOFbGenrD2E6amsO88D/BB
Ib8azfSA9aRtnZYzac1cGKN0+FUvjA1Okf8aKSUOK3cqJWbrUHvplX0JdiWXm/jBQadtUSiPsi+p
GElllzJR6+6PWa9YiCSnA/LdO7Ph8aWWXXB1kSAP3fjIRx66GhElE+KjKRbK2WodvmFKuE3M3dxo
006ghUwFAwHG6dKYEO4xrJqJEdTcIoYEP5aKKtcB9SZb3V8ZkVuhMyYnC2/tnL8TB604WnRIxNdp
Ju2OQOvP4eBzqQcsXiFU+eZpkPQKnwaTZfvmnc0EAO01Vtch1sVeTNgB3Syh3LA+6FxDvioGGIHl
Z2sF1ykqgH/K7RUrN6y0NkxTIqqrWoSX73T8xYbJL0sCN7NQ/N53WGYX6hujCCWT2ZAJzstlchxV
lFMBUugFqkXK3oni2K4nJAA8xuQfsHEOirW3mKvUxwWQb68WXItg58ZvmIqTVsCL3x3/9lG4jXIf
pVoXy0LpEY3ekum+tFndmjrTZkQSXipyNLyMSDdAY5Yqu5AbwmPT9e73DH+PRyrRAwggKCR+DO7V
TA6IergtUykl0aj97pd81oXtaKLdwkGBOZCntgB1JAl7OSCF5yq1vUN3/OsJdVl9j5xCXcb6qI/O
D+l8xz1+AqtJrhP8OAuYkShviavAwsMqeYcp6fLa2RwJGMOjBwBvru08UmFZas1XgbClxSnfs9n1
/fyP1t3BIxMscwzAN4TMOTwG6LHS+IcWguvl9lCT/PjqE6y01dXmST7ysAIDe6B0yNOo1bKp7/9A
q1I0KPu57U5eAXHmExMK7H0vf/Pw6vIeMmw56jGTGP21O7G4royflHJVDxoM+i862FSy6+jsATSH
Fh6xtu2UJOFFyBq/VAZiT/1uHIczk4uNO8TZokec8kV0vxEBi+3rXOA26J2TiB90idmkw4tM52GJ
tWbkHe3HxyKYEwy+sfd65hzWXeURTTvQEuM27AgzCYqoqHijRwKOuPpV4xXvaBaFMmbNGtkuSYxG
gXKy3raO8uRMHKNQsy3raGWDEICmUdut12FYB6fGpLeMBreEzgEYX9E+9UiAv+x42KxCoQW1qS7k
CDeyybllcfLsDVWxRxtSGcAXQmrB1WnXaaBUGLjsXdyZKYFruM/nNQ8TkWkkwwnD+2k5HfFLcNY9
+tbwyY+TnJaaCUR1hr4qq/U3odb8tATMcfiQu9ma029mQOuO7dWQWPH/4ceUJqfw85E526GDRUky
C9ZFbQFQqEPIHqLp+aJ7US7EWe8SSx3Qj/h86LcHwZooRuHWpf6Td/fhAJQXdGLyOFYIUYyjPSnL
XGEA4VeiFMdLUCcTCanWO+3ywhfhlfQAdfwFvVryWs2dDXKEqDltjKZ8py9akUS0ESolxawwdJ4q
JYeadXRsuEsdKD1zqnlmOydk36ZYpbd5fRCJayjxrZPwowt3HGbFJDCzdIIcGXnwcM34Ia5ebnXU
24xFDrgQa3cAM93eGz99pgxAH1NBwz9iM+Lo79F2+eMmFV7O4rYuL+OnFXyctDXGPbS7RYlkV+k9
kKOU6BjMSxXVaTq5a6F1yz0lRfPRLebm8RSv2ilaKQUmsljG5aVrxl3EbobAebm2lfpJwyEJsnuI
jOGPmkLry6I/rU8goCZUzZg/aRErdIE7eBBKy3+o6IosgTaK9rscEjvqDABB8fFWSBD8D/Id9zQo
5Pyp9dt62GiYdQA0RfpwjaW7E6ZYnvz8wvQ5HoiX1QOYQNtjNy8HZRvPt7oeuY3RICziHuHPbeqm
7nhptZfXVPEEoDgB41vfaLVHXgfEW4D+nFA+U8ZyV+Xngeae4wsg8GCI3SdNrvlXOvXkvUJ6sL9d
CNbUYWwJuM9hev9m3thKy5LTQIbfz+MS+Z29cKByS4urLJn7Ijzk96t8DGQxbAhcAsFMr5JiIg9E
TkhPv7h0C3pGJsmzb3pTL5I93suZjmP1Pvmc97CGvVkxj+n8IHgNWHVeSul2RPf/kM5MlQESEjKb
YaHlypI1E3HruL8P8ExMB2JyRqIuGuyow0QPTEX7aC6XQma1j2ObwGnJ7HfmfyHywR+ORtaGNgSJ
xhZE/qMtDeWOsCvxaZ8aoP4yz5CSGlXlKozlcUfcl3BnVBARnmmwMcSHFqKbFSEjtxtMJRrIEQC2
UAI0flq7r3F5C0RRT8yb7HjT+ySRhYoUzOtJKo5eGJdx1X3lusUlvpSm6ay52d8FFAh9MHgROHBL
1Hx3rl8eq4R/poHOJ2WYK6ytFn3RAY+PTV2qquUL/5pASP18OkRtyzG0Reaq03Q24sV+jK7CIW/l
pX7QW1IMOXZdeKobQzRgtg/WfwDIPOyyseuHStmpwhi0qa07lFaBVx0D+hN1v5aHYut0C4uGGIMd
LTFYanbVpT4z9dYC2zml3qtBHlLI6CTZCRdY+N/NReDudSzRWraQzFuycn95VsqnZTalbNkkj/P1
AdKb0y5FLaBIhAkSsVxjPcNO0QX3KOs7nVF/0Xe87n7rsO9RMKiAQd5+r8JDIJDGAPRnYP947neo
LPqw70gnwhcJ82/V42XprN/sg+7hQX74HMH9lq1YXPQjF5JTmhCwmLvdYwJWE7DFUgu7f8YpBAOJ
65Sy6pH+9Ok8C02jmYQCsjGs1s2CBex/MPeN/8WKEs+TNXENH+9Ukcf/LbUxuTI30MCerAZp2Tt1
UkAMmkYbKYwLRV1xlVPVyDP0UZYUO6DhklcDIjT6i7XUF/R6KVN3N4k4QJFeec89MqJnR1pwvMFT
b8EaAyQpI0ZeG5TX0lFaUA4+4zTFRpnFuimCu67xbW32iCyiNgyIWSyB+cFPS4/QV6wX0cYSK0ln
q06T94LVENG83MVSQwRAmIGMo0EjgCbekkNJ7cgbQX/EZwiSNLSY2GiG1CMmw5Xm6DF/vKtPEzFJ
Kg6n+9DXJFfZ6HFd3vh26qSfDCC+n5pQYs49VmQhG6rYaMPfLHWbed3o2/bQ2lOsp7MpzvZI7iqP
FLNnhArjTYT3XE10fxbOlxlY1ucm5hn6moxye/alG67cEaJirgUfyFSjrXeTvC8fXUs5jOK+hFex
tg20OCwNeHr8Mhxo6b2uZVJrYP3geZuBwHB8EWDzEaeeE36IPGARiovK9zZJH5+O8CR6aZi5h4x9
c1Hdv0HZcW6iH9HY3idxd4jrqnJdz+k+uUu0os8SY1nLIvD536o5KzK5WczvWG5iI5bFukgSQuwE
4gYruEVVganEWQWffNZlhqRP+YmG/CkBnqkCXCNdA6O9Uxxe0E2mOgXskvawbKL+r9lGDouLxKTe
4L+9OG2yjR3JQn3iiAZk/bXCQZuce1ZVWwWAPxTCwt0Iw6zfF3MEOyY9yPzQL7muYg8yyhxY0JC5
+cwkoKHgTe6vMzaIX6egTOFTXO2JARgkqreCFo+6nlT1rz7kAk/Y5xnuN0k4csiKYxulQcz7OTW6
GS2by0ZgTeHb2oL6WjgPsB/GwZol3dM7g7RWo06Pkd5h8bE03WFhvDSNiXdrTS3xbE0g2LbBImzu
wlniNg1uxSa9Ht0DWgOndhYbFhOXYVMykrF44hlDFTv/V2mzfphumK9bDEqTEUg0bhaYCdhZLTpM
EhjCN1HBTeUw+9MjRkomMnhrcctpgt5IDZGjgaZIDcr2xd5mpUGCGcoPyHL3WZyaMeMZn2lh7Rbf
uO2O8aaNGroi39+tqNvavtYw4q3Un3qmgv5d7Zp2BEGqoUOjgW9mLzIqv1YlPj5w7sBTvsKhHitu
B8IvdXxwiQpOyO+06mFEYArNLif5RsuCeZnjqUQ8W99T76dX0Hjsof4cfAEMK2mbDm7bfI1jsteP
jZJGwYctouZOa2p7OEEOMd9vsu20LovpNOptwQRUPTL8k7/hxMFB47C91ycop12LVUJgTOBz/cMQ
pvKOs14yEOx7mhnlfTZx6uYkfopOixhjL4sR3KVseMbRiHg2k2nf8BQbRxF4dkZmdgUOI4BjfaEz
pQJN+a8UHzh3lpTLLFjaKT0Gwdt6PYMJfI/Bv1aL+wP5KbcmW/j46d82sZxCz4fVscXv7PtN0yuN
CiZvkHBQFBgkCsd6gfeRqCttVNVQZ2BeF/pc3ZRi5I1BOMQzUcmYrYEEbVrTilWxghaThqQ1W2cf
wj7Zb/kFOAocRWwvrRqqUJ3pp3SDd4BJtXwD8F8jVv9NW85oTmfA30uICYxEKPasE3aadXGIBacx
oFLhI32QHND1OUbnMIYuNw6D3E7ZUmKvxDGOjV+d9gBaVQAyJrsd1cqDD2SwHQpM0JYGvzxZRs2F
oDxStRngOTsB6xLaTkS06caQaakFkd35aosyLvf4tNhvvoEe38nDWrFZoyXOqm12XxIp8yYA0Cft
xcHeLAn/wGU4RHe6Y9Ev+iDdR+5Xfztv2EpUHxPzZEl+vmnlPM4JPG8Jd5EgkWs62gzURLnusZco
HOHnRTyagQ7iDEp+6qoN2FcoKAS4ihWekijJp5ZbEbjB0Y2S/zYXu1nr8mLoWahQMAeu+WHWoe+e
2gmSi0J/SWg/XV8KZsdK1E3fby98ZZcuUyB6kHV6lnSOHNpwYzSxljJ5KcjiNW93PfTJIDFqbJvs
fsRB/Gw2V3YarP+Ba9YrGWiPHAJf4kR+PV8KclPMUBPyH0u8Y30RuGE8QxieghWs0ie9PTBTAPwV
pNtfhHoVxYcFQd5FDUs8syRhDSoI/F3qNBQSz0voJ3OpHJeXeo4jcUFcdl5wGsbNvt6gNa8xdt3S
3t9/JNGhVTq39+Oz1G1oDu/Xg1PUCXhCNJlOwRMVBJBKWoNvKIRkKKKvxuvZVT42Ms0cv32tkKu/
YhPWjhsikezK12pVjEVxD6SQQG7q/X6Y5Q77QRPOkDe2D8jhd0rgJaUQZ0oKvQYIdoZXsW1hi+Z+
WIDWZaO/Ds/UQY0t0ndvQ5f8o9DyIfqd1sZEMDXpk4EMpk8NTUqo+FjJGArSUfK20Llzco0I77Y9
GEc1cRhIycl9RKwFxGhraQ8rVz+6ODOxs7eUkzJB1kt1v7EP+QZpJt1NfY9k74cHlSp+wOsGaS94
6FzRO1fHdJgJ13IaXt3vg88FMcwjzMFJR7pA6HeUwJ1U5mkXgfkqM2nXe9rnlkR1uOA5Iy8SZkBx
wjDbbRqj/L5l7TAdgNoEjuJvFbe9WVhnESJWEiIQVJR5Gr87IcL/pb4Nulf2WmfMAUCc1dUFgIRa
N4DFKxtSJHTPdsO8OFktSDMUHP9Pf4igSs5jHfmR93RwtPOpDPQK5waYY9U5Y0EJONhZ1xk4p79/
+DWGLOd3J9by1o5/yF2/aoGT9cUZGYkegptxnD7xgroFTRjIQmT+Y5YqzM7DofU56OJmNpMRKNcK
kM8bvtLV6NTmtUog+3J0rMMZX8H8b2XWMdd9SMoXH01CuTxZW7gVr/h6tPx08CFBT36iWdT0ZI+A
7qMIcHCpPb1s4hPexBIliHLiQDFiyQEh0cnh+w3mJd78X+8j55tz8HrE7rRwm9SHRNQqjd7AcRit
D6rkKpAziQRqIPuZCO4/oQ5szCcYef+hOSgFJV+lNhoQjww/IxPBOAU9ixZ2Z9Rvb8gl4my/wylt
qNIoXn9fsACPX+2Yq51eEf4/7QJIRWdAjXu4EpXl3qQCSezFw+ttJevXWmz+pASg3lBhVPXU1bvz
LvvC5qWoIBFuGRrwUu1fUn5g+Lg3mRi+GAKDAyxp4ORJjvv7O9WZFbHL2plN9ZRra6qVpnVYyGAy
cQRWqOSobJ2u2K5w5VyIgfeN5/1ih5pXB/VHztSI9Y1DGZIhifAy7tAJ+Xzn6Wq1LdDCXFCmdjnz
iNfYIgi069PlEhfzEMdL+HnqNHrwKjRb6q63rU03L775197Bgjm0gnP4J7h3Omz+nP5eo4JbvEkl
RmUv8uHa9xt+9J7opg/mwhTgHEmK8AzGhidzAmPX9W1/St7l1GPyBvjoMCceTFFumYKfH/g5fslh
4aYQ+OW/eEUQfHEMr+P284doxnJkw5QbpXyIo3s+US4wuWSlX8bAfEN6xson4xmur0Y3ejckX9rf
h1VuNpVwMGlWN2F1YGgYwRRAyzJMkZAuDsQ3/El1AqXlNstXT608SJfNj2+PdyDqgXbRGHTSn4QP
eW95zZknprlxbT/zxNCePbA44Cc5gSci/7UvucTd8NAOOLa42alsGoqbkp+GH5god2ch1dJ6/b/T
yOU5GvG/ElZi/yY1cgIELXDowv/1WG6bnfObYRdIacLmZhJ8zf2CA7z/iF2zgw4g8P/VDwN0K2Dk
Ye8H5GpzwK8d0JI8bYnnHBfVJLweArCwotMfNp+8iCbHwaqOJzsGJbHGq3+6UeS/+LDWDwprElGm
UG3RLyHHZH3SS8kp+AuloRtvyT77KvQYIchQK4sQfGCo7pZXkxb5viMiBvhCvLKNrk11r0IrH/Z9
SpvnQroCeBoIT56dETJIik5ZTGlhG7kKUtsA34FhHteasCdB9NqJBoAwK1PlKunrWUhr38hYYLr3
BISBUY8Oos8tjc1RIiuWjtF8qbTVnnmQ/Yq1ynCpKbjPOPhofhHsdMZs/zeLq4CKC8xSbacBA2ao
0UqRzdUrm+9Yvn/cnbocSMf8HiCXZbqIQV6W3xIfsU5AENA2ezAlix9qwQBBV5cONqeNSZpPIitO
uoeKDRObIcpOhwvrtl6fr/poL+3SbMJKOec7JEV6JS2bpvPQjK1drmcDEsdQfxV0s1bLMN2g07cY
1O16wM0N+74TMFTQzOAtYoCTbl/ji4Z+MlV6+2J3YEV720eOylaABQ/Zy7uB1Q4AM0ad3ZAKuKGU
07eKSBkMWTwLmsPvtAJDFHyhYsO7it/I1MnTznO3NwjRSuoyP+sX1QjGVh82RXsJEpjTDnBgiK7h
PacSHM9oXp83xL5xHSgpXRLOR8hYOl9cRfxxE4J3GoRHp+QpnuzktokXV8n9pUWbXelIKorBOcMs
nD3DPp+4VX5jDt/uX2yzhq/EjkXGqv255qeIzGt0uzi2pQqcrrdQOD3xtnotMCE9/81d5l4bAqA3
/lWXtPA4mjc3WkKCDfS3NPk6X64pvOIAYOiKpNTDAOKY+1HMViaG2bobjMc36eFkWQhJvVIUv6jO
WcuYfzhdPb0k7NMlF6BZHQ5SwxRjiA+7rntkrnV6h5labiTzT4FyRD73n5u7DV+tYVjENCg6JlvR
vAK+S8JDAxMUqI7vXCPSnDJWk3jzjpwd4ElgM1JPYjNZajfYRuXftBkHb7Sbm8nG0gwGZD9s8O5x
uHrjoRRVwKTWMmm8DwTW+fEJ/PEpssF1+bbKIxL1uUmyHTGOa/guVVcIdr+OSgOvxX/DQgMdyDAE
NXDX9ToFH/AIT6xQdLM8V/4LSvWzaiecfov12BoMX45K3VzSMqdFW5ynYFkqJ/5GWCfehwf3TWFV
o4afBOGSVJPYMwgsYIFg2zUmWUM+VrH3Y7lkFLPqF/LGGfhdfOHN7rOA8akozPwA2AxxOzEt2xT1
s9Pj6J11bRbz5wkqEnoMv+lFB6BBkLyD2tXFDkPjvsieAFlcXcNAo92zMUxJPFDKGxN9nfhOiLLV
l5IyqRhrmmNPMw6R6KUddeGPF5cdxuGzOctxrCLRglpYSPlRRoHrhxHZRiTuOerdO+GhV7RDqjeu
0m3OyxeflRrbHy+Huzvgxv0wmXjREf6C1x2LSgKeVkVmXfNF949y9/lnrUFThu6MR3QHOg+c3CZA
SxowgkeIvYgL/pyp2Lr0VfxICfQMGw4g8SGCAqYGQ+2Ds+UWa4v50regi20k7jbnRXbIIPfB/3ng
GTVrMEiRa0q+VxOkTyKkkiEPRJiwY5IQU9gXIW3h66sPOgaYFhRMWiaxt/zXbeSTbo4esspTqrZI
FHZrUP6X88F9wyG9dAGTDaIAZ43Feg4YMhXPfp13PRIrzbd1RaD4mzu/EPywcO6c57wna4UCIOLD
8OeT1ZKQLBQcmF+KIhWZ5cxDU7RxXlxhBdSqBCeI0PSH8IAziBSYWgw79hJ0Y2y5ZoEJJDB3yVlK
4vnU9oTPklCMd2ATXjaCx5tdOlpT5NLD4SyORCpdtSVXPLa5Wnrj9LtxEK9rlTtAmHK6BJCbHSK+
YvezfFfuSSHKebKgeNdwneIONoMX8e3gUflbjW0P4jOQZLf4uxHMimMT+ZfUIZE2sYEO48n02Osd
VuVfqtRvQRVwlc/Wyz/99VlQI9+aad4kd4nMy2RwS0I/v68w2S+qzl/Yf3ptdReO80EXdQSfizXr
x5oRmH6OvhqF/Rdu6W/xSC3837z0X0T9oUF1MjGFB2T9Wn8Gj4rhck6UYbNnoFkQ4gt6jxnKGVA1
OphFRdDUhe64xdVsxNZhKJTt3xMgEVLouyYqDMZdJSm4T3Gfm3xIOh7WlAz+HzhslqTXlRsuCxiC
WjwLX6jiaVDzOKj43wSNHm2+CNBFjhtZkgihK+BY0o53L+qSMou2iZI1/zX1c6Gbvi6VXkzrtdUI
ierV8MAa2tNySLYRYmgpxK37v5dUx78Oe1zS8Ninzn3Qp+Ol1x2Z6uo0PBkvBbfjEIwPbP+Uo4gi
t5yXUgUkZeLOtjF618zE2KztCc8GXaMsgSpIiGm1gbk+yuzeifc9Pa67tGP/KCiQE/DAoG1tV8lj
tmr7Z7OStKzKyqjYHCcdt/2hNHYnNY/h5QL/WtMqMhf3gKl62gJQ4GBeZFpOdAJpdX1dxk/A36d6
Bt3BN32zCAZ/FE+ZW1ARSWJH603y/hS/UqWIMAGL8qL92pFHR3HSrCG00pCjjodOCSXVOb+P+dod
Lhw/7F2BlkXhzZ4kRqDOJhFKhDUXz2DVTR+I3mWqxfExA7+z+NjaTEpnOGSFZ6QuAQE4DNMoY9uX
peISd5XySsqQnxJ4TbYlVgtthGgMA8gkn+Knoh1mtsF7jIT8maqIT1XtwPfHNVdyL7sSEQihFuft
JzYRt0AhVPCx87HMeRuTE64fbmblwTCHjd435zvbq/ewDci01mMy7wDn/yaQmc/sUzuCoVYwMppc
RNKAcD4j8f+arf6AxO094zEVKzRiTfoW5CStNc4pWUH/9XrMcDhcZDvwdMYVOo06vlw2/u8J2pkQ
mXRwAV8uEmPtDy1s20Yjfb1lxPmzwdAHGiUXzrluj/QG4jZxVARZjLj5n8ud7vV5JcWj/1NZzDdx
UpaylZgGHriqC2XGbmqOB2HuWsDW+gpSgkBfq6d529/3soR6I3siMXTMUQPc4jrEfPrXC6UZwkql
gD9WGO+LjG2xfjQ0cGC1DW4Hgz4EbFN42sWJFr74bkROuGg94GAh855QYWaON/LJQMwwoFp2faXX
FAXc1KPpYr5jzYnHLMkM5zffY+e3Z7hcz0JGLoYMNfudeDFN2NdGcxClRgJ0BA9THSVz9ExBS2zH
MdsgvK3a2Oomf+1QGvJylnQ/qbIIFZPjgSDlWo6uZW9SmWcBBfQBF6WW1luSFN1OjHBNTdceDkzU
RhvBwrXPHEODiByYgx9dzGDfZm8qUkK1yjUP61RQ4eR2GEH+tQuZYEH7SzwP5MqOzlTMspzfuqBa
m3gANBjeXlRomWRlgF8OlChErh6ik3JqZLudJfgriW03vma2TINnOotQO+RgMIQ/+s6t0ZQKYmzn
/iK6Oi0qK7HTC+N9egZ1KHpQkpsCA8mPxz1ghe2iJfbQiI03kao6vCXGNgxANZmdxMl9hhbaEZU4
N7j6tgiBJORQRXbAmctPfJpKw+h+QGS9yzPnq43rqwcB75jRZjl7445oS1+BD7Rge9k/qJnkSZvY
rhfFoOLULoMtxh8+PmenvdeYAnOUY5lhmsYAposXOOZ2o67ARCcZl/hksXWIVPEHy9uSZ+OCAVaZ
MzTbUfEySnRjDEF1hL3Ci6RfCmNtyQh65IuAoLxTnkkaoPWu4MA0jQkqg9NNENRLe1DaEzwEL9ku
gS1KdBiL7299k1yvDYf9T34Srnj/TAgRzpDSNvqnpIPSdfKxXwpqksujiJilqUvzlCHgg0JNYqXp
kcu3KKXCIdUZmNJUso/ItuUQTZQrtt/WvPNxImSZBawDtN5ILqKt2BTg/6plfOU2FGIek1EsbCAh
bsKoUMYVNclfFs7+9BPdKM4/XeEuARflQA7Z/iOq/wIcfY9OGYjyl2+XD4I2OvFpzJ35NqPV/udY
+tngUcJE1zh4+cK8AbMarjG/wsVZhB4bLKc6eIOw/3nBgb4iRiEiuKcvZCy1NCB9ZEbI9wvGLk6m
0vN4LMjxgAEhxha7ig8J/2LL5f1wVulse6Tqs0xS5XmsHqD+5PLe90NdqaHp/3G05zplYqEbkZL2
a3Q/DviffoSO4vErga5Zt/czBIBZXNzSHeYAo4aT/O5rgIetFqJb1T+dHRez+qz5bLoDU+C0aXUl
Kg6yYXBQpGMvvVMEAPI0L8/uJq/z7qkMNWTKAxgHlxAxA+zMl4j2vFOtuxAMhPlKTbd20eAfuzff
3/qbewdETuUJTw1F9khu9Wl435NrO6vNNm2+IuSJ7GNy5Vy+Wkdt1kBYOy1ju0enI+IYYOr/ZmC5
XHkDnB0VJg/h9rUzYc9zbd0h3DCjqdfrlX8nj4mywyrzmFuSq9fpWmjinNLEpocUH1A/7fIFIv2o
3Zg5bVaC0lntLnbYGEtdEaPOLsvYbOuzqofSCEicU80JBdT0MAcURcRonzhnhCdio9CefTJ4DQqg
ZUwEwox5k/VuvrgPQOZRr4p6C2GnryO5fVyRMjldKvg4I9sUFnVT0g0PcGESuUkD49mAY6p7fk+s
qjRhxPVmX61bZeAxNSgZmIPRt03ge2Neq08/mB1X2qkoR6fxiyUjKmgKUHvMyXc93HUMxBaDqHNg
8B9VM1Sso0o2pXdMvMm4Dl+88Ba3mAoWRNbWgCvcVRPJ9EPYTOsp46yUV/4BFPSY8at+zek8AZrB
OUQOYu0KzuqrJ8mAi9qBgPIhcXZ4QRGInMUlHbXKvy5rCjHXi9Rlq+0r/goYGY64r72HzKhJ67sJ
6i0Co3WZa/inFefewzrADitBcdN1zVZhjcQuHTuS/DCwlGAsaDD6p1hfoBR/VXAbJ42l1ObJ7sbK
WQYMQyb5J+GL8DfNrXjkBiS4s2ruZxDuuX0/8iQDjycpJO+2q6Okl3h2whqMkzYzmDvbvaEXxaTy
VnVjvgFawdT7074c/LFvhA6WpdRUoyDhYDfVewJtWiX1+/MXmuUYUOQyqP/teAexOR/Fu6tfip2J
4cXGoKSTX3/IX6yfFn8vMopa1kAQ9YlArNlLm0nY6HJsXxWvuMVLnMGcCiluo7tZvfz4Ubi2D5Kb
WikNticGESF3G64pzuV6E9Fj13SEgzGfKBpvqo5JaXUpKPGzs+mtMVaIFeTu7kV+fvSuyOfMe4sO
5Mkbu0xf9TA61OwKXDFgFQle5F6qsm0v8WlOIFRPSL9FVj027qqDmhZkR6++yAt6yK3OD63dfVby
X7AfdLZLvMyyR6dIfRLoUlnOsVrr+RbA7zomd/dcXZnTTgxYSB/CWa/jI8VGsM9XnFz1BI9MfBJP
XB7dhY69cGqCUHpLwvgyflYhmZ9Hkm5XAlBoIfeUxmpA82XVSIY4WX9i2xq6UdTv9JyZ1qY4kgPC
yLnCLsVqCpxhTS0jX1y4aXthiMPBhP7TMD56kuMa471BQoroJir9DEYSvaeju69OvEVuFy7xZPFG
9cV4T5MzYB++K7ifNyMN8FOxh9gP57AcBVpJXGzjLn+oaeVuzmJIciOo+afHrAxEKjqLEGUArJwS
gUak9Eo/w5Mzp1F8Bu+skqk+YwgwO6osqRWyDjlkFsXS2++92Sg6CqDpsJdQJmgngy3ySkrRoS/a
gunGIz5QiiGJUsvLYAnW0DvXzcmUsJx4xYgTLvEV/z4Ln4goi5Hh9w/f7UgyRPOAV8riPp6iIePM
9jm/2IT7RjxhoCkw5ivBSitYQvTR1gBvRi7K/IrHhgGGiWggf+uyqkYSUHF3+Xk/JbqDCl4pS8E5
6gQdS5+E3BIarrh87r3NgvTblIUJ+bWj193Wx4rD7fE4ZMCzdX7Jc5YR7VWcTrFqtjy2Ge8fceoZ
FvgYLMpjMMgRb4yjZLkizRWvy1HNjg8nvH+xdl6mu/dlL/UPY41I2CoTCXVy1ALq9C5cLh976Lf4
vU2rp4iQKXZnWKUgYCOAX9uMwf+dDhsawAcqHB5MIF/aIdAwM+UfcZHtkoIlfbRoQe3l32lmFi1g
QIYAyROVsFboKu973kcpijRX7Er4HQ7Zk4H+ysdDVKet06BkWwh0jO7ZMcI17vUx4XRU1Ev2UhZi
IhaxoYuJpjckABivcmUpsdZMUpvMleRBgMSbE3YK8FF+Pos4YCkgPFxNZoWGMU4mqTL5l5lH8BxT
l34I4uC9qwoxwoUv9Ts4NqJlqg+2kadbpSFohZReV+ECbAnlb0j53fpFO9VwbPR7B4Uzr/9xeacA
LwPG+7mj/+FPpUOHNGybnFtJA7M8LQccDbGDs8/Csdocikqrkuy3UKpASsWP1JXAo+g6erbkoXM0
Xnd/ob+XVREaLxk07dyJWCqu41Gu2X0uDuT7jNjBK8uT9Gv85mSNcFcp/XpZzW5/XeKwuXpaAW1Z
yO75NTUebflxF9hP3iUj3FzjN5BbEja+bQ3xfplXs1fXFYSigToPyzqiuooCts7WlqyHdatmWueG
5CyelQR53AZhqw3UUC/M6TrtxsX2WynBqCF1AMIyZhu6FbvW00sJ2xzpygyh4bvRdGeQDS1108lj
3ZUd0SD2z+25XK71KxNyXjrilN3XJ34RyE5oISZWAEFttuSF2umpRAbncTe5SBIaR+Sp/ZtxZVtR
559I5SYTVoqfGPw40AHbhER0tLUkzCdFsO81IH6XmIwPoI1HisGeDqCON0GOcq3TwQqNutcRQEiC
MazNup+gEilrSe81xGlgqjBpyttOc1p6FTW9qWPay2VG/6J+o20KzauZwTqO1oatEw1Nj9+EMSgL
yIEsZGn+hfajghVJPVytQDU/BEAvstJ62DboaMaImCQGdVmeCvsqow5xncIdUjp7wlvQHxKx5B/8
LkwY4ls/NTxmXq+sOG6cNU7Cggb3MQh92+1PNrD1rWjqnqxC/+Zr7J0vqEEVPwqMMqqNvUokG87P
5yOn4o+k8vCJcCVMRJIzxYOhI4CrgbZcfIgvIxDCctI8p6zUiTewQfLsVTk8zuQIBxWmzWXi0Zuv
9/SnM4Cid4Q14GCILwALXpTKQ3K1MftBxub9Uz08BHKKM1DYKMVgpzyI9Y8rw+Ox7p+DoSPbzrYe
x6VvQmzoeW8IyHeP96yhs+KXjiX6Rktk/amvv0iwWFQ/Y/0k0KKQ0J5Auc01Nw1f7FSNVIFINjGa
4gE/93RvMcQgVqxKUoS5EkS2lK9S2ns13mL65lQkErPBHnb1C61FVui0XSrfHCBeWYFsFRHFvFXM
3hufV+TQ45LFI7VsW6PIAJuVgRA3GVCKza46Od0pIAaUPwKGb/gLOwCIbmf00lOEKxLdwNxox7JK
IV0VPoLheNGtKNF0lYp/hbNKjJdlLB6RPQoS6AtMWxJfwz+2tLVuAlwOrrGpH8n+K2Tkk5vSKEeY
oqK7hFPsD4flkjU6wJ2N5whD4mbNfwllrs2wi71gLglP+drAvnlti14LYbIjKDeko47zxEWv7eyn
34m4V64sVyxxhceRBkG5lFKItCRCdS0KNc+p8AmK4lfeZteh0SodT72UgITVJKBrIOgxF52h53t6
7xGMNQ4AjMEKa48Ql7sR0KK/tn1KwKoSH5617IsPc0c1lZrz5PZ5R5p/+3egiJ0zBhSTeJrsKHQ4
qvqU+DLXQ3WYBawFF1JjKM5P++nr79W1Ttf8363caai1+XkMz8UCyDa1t+k3PckqjxE+ZVjNzzcq
hgwZq4cYjILAxguc8OKVwI8qa3vVJ6F3+aIS6BKfzXOafSzIq+hG8aTohwuUKv/p1F36pu9nqeLM
j92IqRkY4cKDu2MI31iPz3EyyggJRJDut1tnYI58OjZgbEVoueC+Cvb7hLe0ZCWpEXOX6mM8Wb2T
hxDp4RjtQtv+fITk2+Xat0vOr/K2gEVL2aow+rwT36sFNgwXXYMbKSGREonDu1jy0GG35PHYIpUk
7rqTotMOaqqyyMFCB0lKkxMYoYpoCfJUXoEDR1hzASK0SBwkv66V4lTW1vEKQGNCarvp2+ejuFP6
ftcThhDuIHhgx8s67oXEvu0nQtv4Jncsbyn+Ht+bDXoZiMxe32aVH0TP71+7QbBvDz+rHb31pAoG
G25cMTWq9zVwqhG7qpzJosTDkodBNTmXM5YnlbOE4Ojphyl+Mw/FwPJmSSv1KFE5Mq5qTZAjCpoC
jLyK5ritdskBLb5bogY9u2vAtFSv8SP1KiVoPMFKuAAiqFtXaw+AN+JDrw+eCqYlFd7HRr1wBn9s
HWV1maLu6UyppsjuN5YXbk0eqIIcsSQNaTDk8BOibf2E0invBWPO2+4wDc+nrqL2HErmbAyTWchJ
v2aIJPcC096JTo+0YyQpK1UEejgZiVxWEVB+faGHUTS6bsi4FRZCeTLf1OYAfIT4CpfgHTWLJ6NZ
ztLQnFjEgDumXCMGMa0eI5e1ns8iGc7DgsyaAAI6pWvsdZhx/xic+2MlROv7jlZ7BxIAVJI3X9a5
Ns8egTbmEBnkcSM0SHvuTntAwPmuPumOYwYps4ngI/dssqjGpaFm8YGXmRFMfSjTd/fcpmBzWJmV
MTHxQeCWAGV6Zd6xvCSDLf84S2169fyUADlE4SxSAMSyugcnRRhwrjtW6l8uKBBO18EM62s0dnBI
+p71zLBS1aflf4XPFyMfBRh8dn2T7tdwSo3fq8hMt9norwVFDWTH7k+a4QVeFrY4brfK6t7Nyett
v+X8TXal6e9yADzGFtxg3eZeuNp/9px04lTKRjU1UlgOSbKFvoA9LqeBAPjMa4krZzACG/wYH7Jx
1uUwD6wC6k1mUjvhmHDGZdq/wUflmQed7qr5Lfwu7/Bm5hmPafE5Gm9b2Cgo0Wfk+16EMXZFvJkV
qJFm6l3EwLOhoB0z9x21QVSZ8DdXA209XiinJi3izfcAUsOGaialm5oBzBSbSpfJ0BMhawFo11p5
j0L/LRmxn7T2aojRIb10KHbMFWyfkrjbRKZpeW3yYxqY+qD6MDS0c3o9TFqJy/9H2S3/b9uPEQ0K
VtFtbIdAd5C9iPvBc2LeuskBt/aO3Pd5753L6NYZBNffaNqUJ2zuQX3xytZplBZmzRfGjmYzGZ23
Xn/6qecAWe9cIP0YeZeSDQ6UErB67Flo4KmJxiBui7wMfxAQhvLkdO0VourgHPrC5UQ9Fc6zGOwa
UlXmX6U9mQIHelp91zEMme20Yxpx5ORs/n+U/Y2j+DUoPlBfKqd9OZb4WepRl9iJHj90yAxNXjTh
IBlxjRt8AyFc4e6LD5C0bp8NZVri9PQTkbzXflgU3Repfx9DUO9SfCzoeNH59+WC5fXqIkIxCsv4
YDIFQKz0o0kRiOANraceh1pUhSOinM/ykA5jf8KRdwj2LRMD/8PeHmJsHOYXQuygPEjfIzlbNx3Y
o3QFLQbYRrBmrDBUG6VegbGRa9FebSZIaJJU1cxu46MvdsdzeqGnMklsOWficqWKa6GgI1uXZ3P7
SeW3TCEvtjXzlJaUgQyqaqSBd6KMd4qXxLZSKxc417pAdWJOr1SVM8f1l1QFFntnVwvEVQIoton5
2AzU49iFMhLXNv50yO50sM2JIwwtVsUNACh00LAmsvQIiq5V+fZ5dLzpXTrnAw1mwGLcz+LCHX7l
Sms+c6l82niLaL+wNRj9fSj6JmhaWef5uEn5We2UPH6rDxJhs3LABAv6+r8w3hs5IDKP8uN21lEN
TIrPYPj7GbtMQagt+xwRzal/DLPGgVIXKTrNm+KsSiRDwW/t6Wph8f0FKtD9bpjGy1ABJBLYpmgS
Sd/b5kZlmBty4dXxD2SFAe5ZlxZ17CgaBUeE6a9Z+JerWfxq+eZrieeL29uttvhCP9lh66I7z0yJ
hy1Qz4sOVY0OS9vlwzp45Ujy6I5L6wToQXzgKNesYjo+rx+3/GFDI9S9buWtX9WDGRcsZAyaDKd7
hZ+OP20zC6Amj3Le5dAuvS1+voTqB8KxJjGu4JhVpcWzBW1Bt5+Tq6tV2S03Sh3J2VN5+A3epnJZ
r21XX67kgVi5rbUNDo0gH2Th3aK94qzxr78JGrApiNhi3aoKKWAfDoqIpAtMl/fCofmbcQuzZIl0
qysSpWVggNEpYlWQGwYWuS0lCQOv3PyhrhVepAqeW4W4G0p01sT/+ya+ZethHxYN7EhCwaP/6dmP
+JoCYBhfsRTDzc1a6UOygq7bc+raHt+UlZi8kFh0Ols/U2QP0fKFJVL9DPzOrUKUpjukg8jEA5FW
BikeP96bdHxrUovwSVehhR1xOMc5fpchXd6lcysTe1dpi2lC8TywbLeB2M3gxANdd5YNKK1Qa3Ze
BiAPnbvzQse89dumRuwhbsAOFG3frOahSFN8poqpfbUpn54Oumwh6Ixh0024aB0kjZsiz7XHY/fU
ThFRF6qHLe0iLzZ6iHPETyBYyBaIYbLwX5Ud/5GxACp2rGG2+fFblSCXYo+sX6t2Wrm9t4rWh3iA
VjfH5gGqloHBHBYkUlXfcEWrxtgkJeo84jUzcQO1yYSVHdvzRaBezF5jVJonnGwxLi+Dz5nRNg9U
/eH6lwvaaA0Nyerey0n3tZ+7/2N9afSp36Yy/k4Z/oMM4hvGbYnEyELmegg3o+GL/ZNamjSubgPJ
kTiTqWdnD3P8AYDIIsbKOUBTPUVjqx3lKHX8NdUpJF0aM8yFp7omkD5Q4ptJ6AZgO690gfxCdNp1
/j9kkMSXE/JZpQNPgBgKbd60gAQKnaXiOlrjP3Vh/gvZCOoENKvq3nxMzkIKY17stJFCPwA0Emq/
GKrIPy5SoLmwanZbmi8YY2clrGewYcWDaePjBWKsgLHndW9IqQIC7TVDdeqrX1hS7G6z+V4TDze5
Ln0BFi7H5DndUoByMmzIrKx4MpGb0TNhOEHnWdu3/s2FYTzPpDzc9d5m/65TQ4X6YWH74t81vc0Y
tKxeGLm9/EPcnzEfA9WExwkEhJy8ixsa1NiA7uDwO0KuAAzbaYWJVfq/kvsh0/++ZQGnlOrzxGfI
1jrD9VM1N5hhtEOx2tLjwyA/1slPN10+GUvU52Dp15gHvSE4Mf0riok8IuIqEWgM8srQ4syMkSGf
hmtrflAjMbng7ZUPMTMrviKwp20yNE+Qf87gmujBDjXA9B25HcVrzAy5y5DtODJKYXOa/UtexxUb
uYCi5FhZG8lofAbv3QaT6YXMa4ovDsg7HXzOZOwsPGhrJO3jW0GUs8CdTSExLcST/4RIpakPhec6
gfF/vKbXSbpoeswu4lIgcKTsV4xRqGBiLbKPZuybSFNBOKdMnBbxWG0uCaz8JhQpT36NTNhcf6DO
7FFBpmpxG6bv32BVzy4LLaXUzyXg9onjzt6ns1Biwvh7xdvmWp1ZhsTVO4AFIFqLFZR4/4id2AGH
p39hWssvWyVaGDw6StBpAnePCHu/nWaBnhXZs1o8RHYFhZh1bQXQZXxp1U8Nebdo+L2Kk5DbWhal
bxVNINYlBMi4KKdx1lIhbTdFm+tXIH37PXCa5+ye/ln7LfGRMtG4w/XbsgQoFZcPYKXbzb1k908I
74eEifuhS+3vWbpYQWs3own01KkpHKnTyhY5V/LwwuVy0eplWoKTBMfHFkzlw+LyN6xI2VrASHsj
aUWxVHOTu315kEXv3FzpfFnHCom/iC6rZ8JZAKBD/Tj8tyghGRk4TGAnzuytjnJqMjySWJN03ld3
3i78ozJOzpAIAZsY2J5QPOX1kSoQK7kuEyLtzwlMfxu5UkV8F1X3Jjw0fDbsfRP0HqC0vKcKhGPC
4Cb3WDHKNxTmC8XWZv/AENIZxLEMhFZz2tM2xP253OHsmsCN7cBuLy3qzVkztTFgiW7ofiTLbro2
a2zg7PuWEJhgedjOUaHuwbkiF7sF5abTLL7j0ybGpVMLEnESW6YtBBtPIQ0CcdBVZz38IuKHB11L
lnJ4sQ7/s6jZcb8AMjnWLoDitgbNR9a/qPOgV4LiIGbmtQYB6mgAlR0fib1PziV6xQgM87vtzk+V
oDmemiglVU9sxvXZptR0SzxmZm1zVZpVstRLRicMm+Bbp30zhLSJo2F/Yl1yv82pdTzIHwwTcPP+
eS7IW5lcw+HypL06ym60WxMRfdhHZ1BgTiBgNprNwNClEXNTQjwgWzXhWrNGGXk1v8GmRxD/w+9Z
NCEYEL0XlYzS4gYoKOmtgiV5kBu0tX9WwuyPy61E0jTVDHfSSE+xfAZEFArRwyqUUb8N8W47hgNr
wkeqCAfUcoVNDMyBDdRgNtX4+Xe/btkMsOw6ck1h5w63JjN/7qEwRSblk31G7iWnjHq5Sdk8kHic
kQB9qx/eOogtPRqNjGrbt6k6G4Ti6/H5lkxKruka9TMeywZPhFibHyOoo6IUxdxCGNIUuGUXvUXz
UixdMuDH7r91yobF789mT611Wh+gkc+Yhh1/v/2WixTRHDW/XhrcgbXNcz6HizVTkPfAJgXCfAN3
9bTtqNvdB4qpVlnDNIvUnRkq+e/XRh5M2dB8JcHrmhHidiDmKtnmU7lVtqXwFCFAVniyu5xThr4i
jWsicvYA3gYLLvN9o+ArcK6WRGo1H7vEd6YiJy0Io7Y+vAv0zadE0p3x8hKQYyu41xjhfFTAhx89
Q62EdnXrr3a1C36OS7h5XSahPQi4JVCKeILv0cck0dubSyLeCmWosysmwaJRPOn/zmFHzKCDCrFv
T33YgAvSVc9xVFHbuBT3FBdOyTIFAOs1q/hQXG9HnVmvAZz+vmLHnO5xO5G3ATOSqdOa1uaFZio1
dIn/byrOHRBhJ8/glUX6n+78xD/Up8RuhU+OlJ1mrdCF2ZcgteS7X5qPmWsBLcSbhe8L69+T0lyi
AKseZMVsoYdbYp7qAHopgNadc6pN+mlPkf3laS077VWGi1ejpVLQVN8zCdciDVxbja3s8phYu7jI
GEtm603raubyazpY4XiZLGh9kjXfnLxhiaKOQG1oFlzvaWc31LnlpfPCBp1lBfZRdLpzlfN5zZLH
8VXZFlLKDAFX1CrHtKt6QDAhGBOfk2eLnUn/VfQG6MDdz5L6Eq5uaf/nFYNhpgRBA2rriR1ycKbi
UPEwbAuPV/LUY9r2NnEl1baF4JsEs0vQ/6sW/c/eb7/ACJ0HTn8QkxcfI2YHVxu0FbPdjVhiHPkr
DJV79Pm1+vwjc5tn9rpTaG50X4kZV3w7nl1cCubfUJgUs1+4jhn3a/63R9G+VHh6mnxyEyG3UBz9
VvYjReR5covw/xXHWjiWc9+DQH+bu+sOkVPvuhNWUDTLfn4FM75ZCA9MTbwETVlB4wlvRrYcotlO
9GVCbBk6uz0IlEpGOj0LTU6tx1V4OGFpwbIJ645ccpbwpD8SaIAy2HTBNDNRwvtD5oSftdzQDTtB
yTV7Ss1QUimqVPNqusZkPmNv3YuFwelKU9nJ4WAt5aHfx53QFBV3Tc6sHTCrbDFKvOlRzvsYEUCK
oyUKzKtKOPTp25SMF8TziJOYMmphdSQjm4W5TPhuLYw0KwPD2YvKTdzNCc2Wx2T1h7Kz9rXaiX7a
uaE7U4SQFiD4bcoOWqOXoNgFwxQCQj5SkAHEZ0moE0bDeORA4QRaQ/Mt7u/OX9foOuGkqmkU+iPF
UqYGk6EVWpR6dme3V6WEwi/JAsQzqbZcGs9PUzbJhs4ccVh9/o1SrnPvSQer5E4F8B8T5HfrnBT9
bEl45tFCYqluRodMvKM+bdLVc2FRxLzkrV1jqKCQ+FIgayXS70813VuOWGXY7ynOjIX9UbxbfyGF
6Tld3vDUK5bNJyAJNu2Y9VTQnm4nFMcQhC3JgZFAkr35llYpYY+oIjNYxxkndiApB070bWo7sdRJ
g5qRy1EGIG2ByS0WK84OFgTKumeqZ3M0wbNtP/zhElnaicgKLUUhsZp8BJfjkuelEFLmk65vlD9F
YnxgLzPwRkFNGLDsdJLCuDOr3HtV9LbTlz/64RGOf5QaNXOXjlOOMl3JG73xCcY2X8YGjxs46cp2
vq8WDf5TiflMgXhkit/c/r1tWGNjHTijEFZ6JOL1/2gBrxf3PENBxv1FrPNknQ3I11/9xFaNGn5g
P8nQtbaIxWkSZYFZCXdjeUp/FT0qNDrLVLJfVAw7Nk58t+FZg0PoH+o2zENPWj9u1quAsmU1BpQU
cza4FfO2ECD62rVEGKrOSIy1+C43z20AxOFxdDV3KjnSrMrGgQpGmpadLP3xK9+Do6QHPt+qbwhu
3g9Vz5P1LVlRRbHhq0oVQmyXpvcC97ySAV/+GBiLXyE44QzxiYrnaoxQpX7+LpzcVy85gzgg9All
wYvb6yr2qsKZLd9OFTmhsygawHKxf3/XYFFIg5q2oeWpT3IqVt8M/8gjclf9AtpiD1pZkhGVqWzL
+9SvGrdWv/1854mOOoTb7qrPz1kXOOEbvwDTo8arQDZTMmccNr6jEXlZLpnPlXjao0wqF742FMSs
lV7Fu8Gh6BFguAB6dBz2GzHVrGitvVrVQ9O2QSV0APp0U2aLVj4QUiN+wkN+88bWE++Wn84LPxSi
IMwTCENcpQxoUj0/PADL7In9GbNSecNYE3mPM4Ya6YVTlpiZ911B7/JCULUy7PuhOe8uWE5xMNOe
xF0DKLEwGaEYZXmi9L948HVE1MjB+yYhaqlcszhm5mUalHLy/Y8mjUFEUrnWc6K+tSCis5E4V1+l
/si18IcwiSMT78CUc0zN7JG32dQD/IrHD4BfoWK291JLSo89GsFn4hTs7EjXXLCyvIxKH5Ji2za8
9YJhcx8KIEmCLGcXaGGGqPWThV1brtHo9EFK/SE9YX/eAZXvyr4gGlnL03Zm8JKpY/meABWIuNKx
SDgVqeohZi3MzKSOnr7LHbJ4OzqXycKqVuqRkwqD8qK3lYmmGHSq4ujJpMWlxrUyxbmCyMSbPY32
En4iYTLRt1tNDTV99EL65Vov8HXj1pWIyx4skcLyfFNInmUCg2mFJLKsYj9XAExYtMwXGGWHQSw9
19f7Nu3cvHosC5jHlDcbNwrt6r4NkNJ1XWCF9doJLidNbCWdrxLU3WHqLyuxqt+8aUp8HZNSh3OP
ZEzqXmRTRAXHr3nKc6q2QJPzzKV5byXDVXYYIFlWx1en/cRZcxi6NGxfWDyJRD3WcHpNAWjPJCHm
X9//k6d0rAbNf8FX5ux13P0WlgcjqdtOii7OV6sBGAh0PnyCiJqREzuijUMbd+P7KFGqt+uFuEO1
iXiVSJ82681DCBgDr4SbvFk450jrKb1JO+sjxyBY+rq9soc02f+5yIeZIsbwzVETOnUYamHUEBcC
ifwXaUUhnI6xStpn53fYdJlxS5KqKkBZzipji9wGgIgvotXrPv0nFGPxOsLfcM2TuR4YXm0LDoXL
ugX3DRhJlZAEVVKvMY4iUKGkZqkf1ozY0YWqTFnJmqerOpB93AF1wmw0PgvrTS1OCKSpq7N433V6
k/DxENHbfT/+UDGLAbBQ0+2hZ5vvCpZleVs9Okdm3IBVZ3ycf3KFOMfghOKS0nJEiKlLz4ryskrc
HDceH1el4KFi3TBVyL9EBnw8kHExq4618hlKGx395ltku0D8Nmd8lKN4WrI7dv2E921siVZi0XdV
oAe0wuH6jQjzKQTAfMVHNg1uGPpXjV55ZgTlF15B32Fd7eb5Gn0w6UWVS4j7NB5wSm4luj5bXNpV
KnFPubo69fO0TbwXXR4uyBYbWGsoqbOERi+r3vf4kKJ25moqEH/kv4aKX0tYJGyL9Sggr6xM2H6D
jqfSfJ6jP6hDL4WvJImf5ZEJifS8/NXbpHUCbj9NdtNisozYOLB/wlXIqiEaxw0L1mt7TGTkQaL8
UCQeHlmgC+DczJQNEhDjVn3Ilmr4CR7k0OExvE17mpNmDqXiA2VmhIrOmBtEJ/HQzlfrAxgjBJ6r
AhowclHge8xgEegZCV7NDomXc76zc2VN7MrIbdKHgeVNGaDcGzbvFU1CAP5b76TTOXEd8of1cTj7
Fn7Et/MYabI7yk5B8DhXCL5kZB9aZlRY9eGAtWAGugeYULNvKOvO1ev7bawt8fLUYPhF37K8NXSW
Hg/wICKzs2utBCTMRaWUz4fJv0sBPVWI3S35FbLzo/IwarEaBInnxBGIeKc9k3tRtLaANRoQUFGR
7Gadm6w9EmmFe9twcphDa7oJrf7j8zusy+oxt7QdUnCwJ8AkNfeNIeDHtmk9FWycPIBc2ER/alUA
KoFeyvqlWmSvJuw8pJq70OGoHfm4XsD+zYEjfvnLPkYdRhNi5irjnCjkTugTVryxCocOMMLCYEAO
EhlR94l6gOw39IwgHCIEDaQidagqxul1BtJTAcQV+ivQo6euFImkwQ/TvYo+0orvF6u3eKsS1pom
hXMlUZjVkmnfsBx3FiVuW3jRTFpvVUsa7nJ/+jkZzOpSTmzuFo1cJh42wrffHLm/ZlzoVRBrMsH/
eCfYJzUlsRm5PzXAW5bKITYVef7kPDlD5h+7Ov5u0TAVj2l8pTGnVpJsi9xGGfDbJQmsTZePex4f
m03LoGUPoN8ZCKLrjihKq7ria4JuKrZMQOlQq+dTf/HFy6Sz2+uGCXDNxQ5FPxxIntIep2PgITtf
Re1REiS3XZWmHpIQZQ4lI2a1IKshqZiro/usTTVDPVkoZ3CcL6eTXGkDUrJxh1YQGR+cK48jna8p
ALkItiZ4be6MhpX5F/u4F7dkNDRGQHvt4shgmP2HLX2PqsqX/HDaFPf8gi+s36YOS+3FJa0sjUpY
kIILhrX+sMN/omaPJxHwLypI4b25fDmEelv2+Dl8tixBgNnXJ0Kqr6wqfS4IdeOwtNSdDB96D4me
AaDwhZfer79gSFDNsXVT8k5IkVSvvc09x3bPpwsNwJ8i8SttnYiciAx2bA92FucDFX7BX/b8osXt
j0CZv+5hVll5bft+5rbBQlkbto9tnA46LrH7A9Hm/fjwb9IGnlwFTPXKb43uVJOGNdYJHG3eLbue
/eIQJ3S61OH3M6YL0TQq4QfaQO2moZaeNNryXdNUDJpuTd1HPMxWGEoZg2DSRt1iJS8TSZmaYw3h
PmtdxYLj9nyZQGt7cYJzWvqbQDyChWmSgAWWoWYo4guYBlpn0luO+hLwG6D1ke9rRrF5wOctPoTU
M4dr2o9xRfEr16RsMuSJ9vr7dCOJUsa8IQcI1TZyE7xsJrJcrbB2o/2nHAYVbEZotM8+9IRtYQuR
ZGUNzpDbdMLDbA/92MtiHVyJpBz9htTipdxuarm6DC1ajE+/7NLadeeT3ECbJkioaTvbCc4VdqjX
pA8X4F4tbGr6HBRF8CYjlXtusOQuXyEKSQtKKZe3UQH6vNgeUEaZk+c/QLQbVBnEDfoFLAas6IWJ
1r6h3G/oL8XOcTVb8jSLXtYId2xmtwqEpDcLsp3z3BYBHAC/8vhallX35S2k+XknqOmKahhM8YmE
Fh7ij257jr8NLJ6tj4+uhK1mbygV1mFkFfQdd+1lAkQVM6UfLrwyIkjj7biTlqR0IrzvtUDtIbuW
OtdnHeBfUXTvz5U3BKZHHLDkA8qMurCQD8Nj9Z0ilo1vdCnHKtyUaX7cF3IfAYd/SVbaTof+ljWv
DQ8PekFSQMG+EtX4IWQhUnlQHK7iINGmlN0v9UmzAWsJZqG8iRB0filmumib/0E6qPjvbA6JNYlG
dPR+ECxAw7kFK/xD7o0lXE+rt1aumcciqqufKubJHZ72NEyY2g/xoCcvEi/FYuwDJz2CKuKxYH8v
4OPxLjzJ0CZpjxWz5Eovykwijx4GuA3CDHOfjK2H7pgP5TAz3NrHV6uA5+nmaRiWiWrVeM+9axFO
3yefJqOgPC4Sq02UvfiQOrRe/vFcbhhguvrrGoqRZLnhauG+Du9GacX5W3S7sopNTJUoZ1Ak2dwd
63eOYR8vMN4uXPAoh2wIF5sB87UfLXwzc9KLV32KO0cdIEg32/vrW95JVGdhG0r/zNYr1ktoigix
AvOy2fJ2JrEmq0EoUNkGcCH2a2MAGHfB6N1vqVNBwRIhM4T2qJ11LZ12MKGTzhL4JCKllbvj6Vlo
MnX769jcLQAYGGniCKy2W++b7dtAEVUPLN1TGMNT2Uazgprjj4nCpbnFFLNBr2xyb3mDYbt5/hHz
Wwf/Td54i8JYXUEe6MCcDem3141knVG9gB0TiXYoUJfcKnEqmMgPbfzh9ADZs8Iky0XWqONgePGJ
YARy9yzVQDo372yU45ylrtRSXeyU6IBQjIzJ2pdiab49FL/bL00uPjRhEI2Mwqu49EnTJX9fuMFS
UvUX77fVTodYsExJcf2a6odgGUSM+QYRX61vfjcmcEWvR61C6kB+TaBjKw3NhsCVrK47+cILBbRL
3ghKGNbURAABhtNtqp4AsiO74zMSMdvvn+ViYAXwURlLmVVDP3LsyDst3ekPXwvxzIOE3coc5WNw
r0bVGPnZSdccLVWL/HDtCe6DUSvslgkPXVho2F5RFU6yRoZB7ixFYKAozLT0HgJEXi6ptPjs5657
1bh8GE1ii2we+ImIpvAJl9l+agASLnAdMZAK8uXjBIX5IyLVSC/nqoDo1xRaxdOEedyVLVz+tbhs
2R6qu8D6I+cvoZK7VRuO1urqsqbF3raMlu5uMUpMIuiomDfa5LL5/35f3cFWgnaztUdo26zotUYR
IzwlvXnps4hUmGo83spwLwYaBBEJ074Yu+a/9vYFMYEwFlyiyjhDbdTsINKZ/I4uDPt8/eHsxjaw
3d1aYQEmPEHgjDfsL0a4MqSfv2vNn8P9Bg+siCeMXP0rz8yvjBpeShIYhVECb6DzZHZaouxNw4vS
eYh8s9/00Swjt/BGflJQM+yD0rtioQR2I7kj014gJMsExuzuc8rctuDbV/U9g+DT4/DEQXueTPWK
SR+do/nVSyUSgnV8XATlBOPWWMqK/kKlJ7AE1L+qxqvGelaDHGxEfgTFkNXa0ovTdu9y+pr6PFL4
XtRqZkOHAg8Paixv2m8m/RN9s2A5BugzaCCXkr9FiymNxDbvsjKt3DT7E3nrKd5iubxBVoI4uuV/
mu6Zm8eg46sQFtJc4Xk5HzrViLzCQF/ZkkbVg6Qi9qLXfg8Cfy8f68dt94eOz+aGHr58hU+y/rQt
q8L5V1LHnxC3XXw1ATmwwJCuf6MRO22FJ50vhzLTfbtLeSK1Si42NDQnA762cLu2VOQYkF5Yha3d
Gm7j0Obhj9ls5f6AJejFXVSuhUfS9ThLkPr4Fq58HNarRUWZOMF1ZVeES/rMqf4KEv75BzNvz9hI
BibVNfJI1B7ArvsIyu1nhax9FQ8nJNK/q6uJ0qNySIh2qpJeFTbRuCE8RAJGaB6EEPd2FeZbKZ4f
vYnfaXGu9e7JVf3wc5DghmtojsyKBPKDgIY+2/LDvSOs/Y5Tbc1KKrYlf5TJBARj9GIWTnXLUeXR
VVqDqyagvvSux/E2alL4dbYhJBhSkj3rxrMOqG7RRjsFH8/iqy1Id4TEPRK2j2bwnyN344AzOOS3
RxH5P527xRwArey99VsWtIkQlS5ED66pXsZ9oUCt6dAN1rdmO0983IkRM86j60CnQOVfZT2adsVg
ZD9BRc0t7WU4Z6rbwkpc8Nt5U67fS5IsBq1GtkYeKULgRTz016EPDdCgsHUXgqLYH4oFon9YwsNq
vYAycrZXJ+A235zwwOexLJ2lbLuSWQlcydXQgnm5D9onitnJ0Y7bHvHNFjHk9tjb+3t5EPwhwmA0
dRQwDZPT1IytcCHtc2D+t7bWEfxd73tiWjiccBTU0sBlcD0irx1tXBUHkyjSJJWhWvOtITEI9CbF
dEAilg16EQE6171ieTjH4qCzGRaFoe5g/NNgUOmYR6Uxbw92cqrtwmKjictUiAqH2o5izxCp8GZl
OgFW9x5kqOn/+fQm/A3xKZcwf21WmjIFIbzvVmjNxpJxALqiBDUcNRonUsdda+V5fTURlQ8c/fyZ
RFbXmeMJ5OxO4x/TYj9jafGIvvIao3/RTcqIoYfjvo5r0/G9CPW0ntRH/WuxaRNlOSJezIgIHwc7
kOmsqHRlgqe/tCKmtaze4Dtf0HGTeMnHuH7S0yXQUrnmi5rnKvgoXszDOaSvTZ4yV2a3+ndvhQrp
7cj6KgxJFIltP82YFI1NFp5NFt+igGMeZSROwQpexHqwevM0Ps8OS5y1Iwa6TTl6ApywPlLuHwSE
IIpWDWualq889iE/7b1xYCVk97IQQGkBacowJ4yTTL+Tp8fui52PU5Z5s1E6rr/i6FFsvqA5VHfc
xG0h/eq81y3eiFOl1fj3ffZCk/x8sspT0WRMNAT2de4zZNChUySjnn5ScvcVkANs3Xba3KpbQfX1
FxhVy0O+r9NA44pNnFXYNlENw6LwlqJcqeI51HGZPzoAq1omvsVvAPKFiZMZMNCRlN5e72j8soDT
KaLkN3MTx43Uwr9xBHraQLfIsTXs/s5VWtoKz6938w/j6KxwzZ69MUrIgS49ppDtBwZ2G8jiSWs/
2+rWKPNJfsUnQ2Fq8U/P4EUIJ1UI/fq9ORxY6D1kVT0wuSjLzSJTAXRKuRdoWEoYsK0BKlkfbzGc
SwYQRjU4fb+UNFg5bXzbO2uIlkaRW5SqJnjUOZkmv06QuJPNBTFfCc5/3ocau73loQtQvF6clbzI
K0WHlJlBo8x/KDC98C4AQoxq05ZZeyNiCxpzIaI+fkLdelmYupLVYSyef7CfqOjpv0sDAkQ5AAkY
gX52Y+oS2IB1R7aLcJRw4FsD+ZAMKhRphPEBFl04gBWeNdU7Zrq3xDaxMEonk6TxBHNfQBP8CJ2w
Vg7YacjTH9ur8z/NnnQojUOTQoc/ateHbP7dWgE6/Aeiej5X8hb2i+ntXPz+i1ns6Bxv58Hpqrxs
IPIo1ZgIMrOOdKyNTm0iguZO+1JFnPPafiZN1tLSOqR3dqAyBrxDlbzzcE4Dk+jmeBnsRXIvdDN1
Zlgd6En3QA2RSqdR3Po+ORvBRqw0XrUHpPrIeke4rVvE+ALzAtGSoxpFDBFg024Qz3w5PZr6Ucz/
o3xT+DEv1aICxvtgMRARR77fvxNock7roFvLZcnh0Ca9znKQDD+kmxuQK/t07YZASzkClYoCmuyy
w8MZpbM9moCe2R+shEBnKnCpDV0BUsan8hEqekao8sTfvVxnjRBSChu0DPkvwp6s87j96ysXcoI4
CV5H/QEhKxGHk9sn0/biqNlxM2ObbGjRcdR16CgfftIcQyNgquM0RhAvqvA41b0EukOa6jNR2Z56
So0WQwOhIM7zP0Q0AGqoN9UyHVst+vzuEw9kXNcIh6ArNTueKTD8ERvPWz8hXvJVDZ+YTxmuutk8
n/O5xkQggusAc51NvBZsUp6eiCu1fr/hhc+RrPDLCveImBiBIeJn3Jc4bY9Z+9pKePwMdnS5HaGe
RvoE8Oy01hjn9KSgfHyx9TOhpxHQEdYDfyZA0V1gu6RL3W71MV9qVNebvLnGJBovKLlGlOSqsX/8
l9243bWSdUJD7fFW9rXneVIm0VeIEm+AsHRcuUgmImrki1Dbq5q3QUORsjmWm1tRlS9eU6BDAO7v
CwQSIaTrNWyOfcTbTDJQqiNuBr+CU+mpLA8mIwM8oX92OQNPIEF/qTKkrhcUX/WgJrZXqc7HSvAX
wlRDHUtX7g2eCKm3RXGECcBW7ndrj/23NBgOZTBGp9LIwNasqnR0Xx5TWi4snWs1mnH7Bjw3Y29y
rcsF/7UxS+KqrWO7e814DEN2pnHrdQMuC1pjmRIKcK3tIsUm3GFjSaHncpX2G+K5Ee6W8HlqliiG
+FXWIo4mhikzgZb04ZmfC33kI5hNiLMvZ9KTxoz7C2yOi1MZbPXWJTyb2xz1cBn/I7nR+iozEMEd
H2bin+qd60QgkIEjXj5pUjn1gLZILtli4YYkWT2JuznfSODH4qJijGHbClvh5jGZ3zlteA3OyNWv
7tzATd1xPexSHWZhiHg4O35mMM9LjmWuEMrBY737LghdaIUe574JsyYYSbfiHPx9aygVchLpRqcO
cgy2AIEH2FEVt89z1OZEJEOWE3cteF5OWk7LrgdNBTuM05jS3e7kGowCIeEtQcE3fVpQzqiF5Q/e
UfjJfLaGDMJixZPhQgWW6WUBxoywnQAWbql8LPIjNJm+BzRYCgu9CS5EjWz8ElU+sekrRsFLa2HB
9KEU5WAB1YI5kHB8CTQ8HQSxXPJcE1ptFAk1odN4ub6LdXW0vk0zmjWo/tF8OamaNTk5FolxG6S2
Ae0yZy8se4c5aK7NfupLsq5RfdP1gakyXFfpDcgFKfa437v5HnsLc+BD/bNpbHZXd9XwPZQRsg4P
ibNY/ts2DRxiTV4G+cwfL/JXIhsDVGskqAtxFG0GYAx8OOuIL+IC2A1P4TmPxZnphAYsUmIBDX/Z
DPRrJWKWE0a9hOzxJSwPFCFvUFkmBq4lkdFlzCQwbHhem/gRiu2upILcXzkQbOkij94L6X5jRqy6
MpPbAac51IXF3Qb2F3xhZhahk6pVva1zheUmqzycrf687+kXvzHULAqWnkAbLRZb1gKSP/NVGhGL
feWMffKTVlG9RStwNjOVBcNewQoD6V+MOGQNuLveug7Qx66ncArjs9oSggN1hgOua2HRnriqGGzZ
V7K3s1LetgqUgKav6Fq4ikrlgD9mngwmtZI0f8EzJr2vB2IbwTAd9OgpFv9WDPWWgTvU4cM7lkgM
IwJhyUEwAl9QHvGXdKIhh9cy9DhBg+/1Im8Q0E3MsOdbL+MwqpKbeyxgulku1U2Gz/rkSN0IMb9Z
UDwxPCD9e3HkBnBH5ACVVCE5oBf2EdVjGWQHukjeb4YEa+0+KEbpbkf5prYP3bIdppL17MbLXfdn
HQwo+R0QrEU2i1iMo6i/W0PTyVjkvWAZFKJc2BLenbkVe7tlunwasEBi2IJU2Fa+ja+TsqM1T2eI
VNLEBXR39zNOqqevgXvBnIzGUMemz3fKe8GRz9Q3n/L6WGc2SAINVnTZsKdijqXhoiz2QwPq1HlN
2GR3U/y52s9K/TUcVIqe7h0jSeYW68HU0dnH7zPZHMNceXv5saoL/UKFosqynRWobvbHpzWQ9R8z
bOO08rm9fZiouaUJ15ZZPO+AAKsJgnSj12DDExoHE/7ZHlnWqBHFnluWGBpoL+zeTeoR4UihgDAz
sf91ERyJuJ297pg4Vje1kxVwpkgKav5BU8lU9cMRXj44LQ5Qn1TL2JEifusoRcgjFr+wj5LfKkzZ
jX+p+C2njwdmgoCV5vf9WN3G/MoMxcrdqQJ9sr7/rJ0PkgZaFVBRvk/TmJzFOZFf0qBa1a4ewsNo
8fvj4ezUHjF2Fcip0/8oEuEFjbd5mrxIBL1vR1T73ZX0YWZjVqgSRtd0IKqoKEHrY4l7I4dISDbA
eiMV5+0UYGJlkIfyYt/XW4ALiOyxA9hTuHis/1c/H+DzzusnAxuGnmfqwzy2YIrSkCgj2iHHKCv0
mE+JzvwxdOV55Ptzz67Vn6DgVGfObPhCiUs8P+eCGzEImm8OsVUXQwKebE7+JyC8HCxPNLJxP6pX
Sz+/STLhDcfFsq64zky2gVQN9Ugi4Tb2SR7TxUEizK0xIqpDt6C8VbPQtmiL7Nv+kBuWKWUeyFqE
tHzrxhtZsaZ/6aw3LCXSdtrWPcgx/qumKs6IsHbqFo7MKWlTxO/Lc777HXdKV8VnsNUwWYjR+IgG
j0DToys56PyP2MtAmKk7X7HlRz7lrlntSQsCOYbfPmZb9eoM1V1NehHsAF7jV7duOni25fFEYJDG
3ml+sOThMJd7HXGdS/x03GyS14VB6W5GzXfywhe9WWyLZMU/9+1yvtJe97T7vRfHBCkLeNWsWrrY
cLwJWsK/MghTp9dRXMFbMlInO7gHloZ6Ty40YRCxeKAJCxlQ9tQgu/zurNj2xhYiqqlDFk7XJo/j
PWi079bJM0s3c7OI+CWkwYLPzen6JIM6ag56RForlWK21UMfQET1XGaIFS0EEV7Ft6N25v8wf2y4
L7svapntuLA5zaL76CbEJ9Vs08QkVMUV9uucyy8KJ2t80uGbP+HaJ2DGSpc5k0JIErSmARR2V2K5
FqlXZ+3r9epBQApbrQf1Bq08215FvL+D6TIcizRIWGUX9RYntxtjDgZ06LxtUg7VNES+u/tVsGFJ
Vhxg4WOfodkvUlhmdSLqNYrUAHPDULKTvIi87OGPemgNkoTsyJ2tv/Mcz6W+OVQrrBmSvPI2GqPm
MF1SiTihlyDq6vicdy1nk4QtEEqQQUwj7G4+OchB22YQRllb3eS210ZJM2lpWi95u1hLGX+nB+bQ
z9vBtzZEpWNlZFah0OvwLVB/CwsVW07P1Mt3ama81/x3W1sl6urzjqwJoQyWXNYI0f6ArBbb7Q0o
52N5k6eUTJfToHJh2tWBqvl1RHqUIlWHI+onV6nyejjwz9A2+0zPBaacmvitjNpZaZzIB4dwZBT0
rwIak31fxrO8oSJN39wegP1wvqSzWVQWAcC0vc4TkSY7Vxtc0hAHU/U6ekUHGxx1fMqHUK6Rj3us
3IIGW3WgZzVwq8CvasiXEldmrHxHHQ6eKnQ+cVBIATiPwg0NXMlNKIYbWT+J7i7QWe2B0le4B8sS
pSEkXV2gS14oDf2cCEOQkkZbY8XVPsnkWUuGFovmlu4S1MHeMBCOoBOnZQ3b6YU3dgDrnspMMN2l
b5PRne/BXg/+bxphr+oNRWabWvvkG7xkVOR8XvHdcgZhygfZRvAlHQLk4EZQeKPQuzQCXRjElWM4
xMr/tEPAcGBVzgSvwhRFyXLUq38rMK81o5MR+Igkp17TzH9TviJ/kGi21qsP5/ofHoKt3EedyBvw
DgLCUwnUJPUV21dI6GYeCBYTJb/3B6iAXtZYU06JiMochZRA74R71pRdANU3OsNUUTcUP224xMIL
HzOvnNV8aVUcaBXUcHcrAREm+upnDQR5wKhgRAKBpI/Qm+ZhGFLFBm/nnWYKXwg5NVIerJyYTugB
sgebu1CuuKxsjmxelOUlPm3dOUYW3kKHCQVGaQBv/AgsVWPFuNLyqxgjjHqpcHZ1/bL77PoQxQ/Q
TSdJEPRI7Il0/xDAhVTFK0eeR0KjMWZkDIzfaAm/PaWgQ9o4gaSYfmEDB6PNNT5y0aYrPXPrQFgm
PypRBGKfDRF/eBJ1q2oUZDVWNBnq2qQuIPHYHBhhoE4JILijf4H8roskPPy+uKFjOiN72lwbN/yU
Pls6ZCG6PksvLXuykEP+79+ZQss8UoEBUolb+f1ikDBYajskS6lA82G5o3KJ6lPB67RwTtWhhlIq
Sb+rTyUG/6+l0aTqtHFM7ZKw1PGkL5jbciByc9Uz6C1zhvOECe832rvzXfMkMRcpEdalyzsq2aeu
XTB48LAL5RfB0smx4b4MGGEOhKOqat8gkSHfalDJar0JtA0RInloQ7wrZ/vR8NT6j+Tmw9Smij9D
1sx17ZKqLbnKjOux1y04It7eSGFdEuW7pIeKevD+Xq2uWOsS+ts5SoMd3InJbqerKbfwv3RjUO+v
SV83lKfoERMFen9OeDxZ09/elPzPP4VBpjIx59lnGpBBOmezfBQbTCzbBPRtfWJehTtvUKmgUNBA
b+daySmpOmzmLj14gYfu6w0a3H1aQpK51OQp0MD3J5B9y2WqNxKJSCceLbxVzAoQqwLuyS8YZ3uN
P8H2ie7UCK7dydqXVeSSh6vOVj2NOc7jbuLk20ApXNy2QJ2CeuXclvTHZYLp03pZGKfm69KO+FEV
5jKci8tNMIyVYEurfWxy55asWgI0UeOkef6b23MCRjnYkXdlHrn9RGOkc6/ADIKZca1uVn+fwNe0
by+DIeOoM4xUiQDO7cD6XqKkV/ojSWqXFCryR76k+EWY86iQ3KSfFi5wXRINqMNJEzVAldUyXmv6
ZLC+ud6DiUIMK1Jk8BY0BG1/b7KrcJXj3+JS+o8/MN7wyURk4K2jstvPJLDhagkKULctHaMuonS8
k71rN6DQLW/CPHpLFA7S2ewHiQNHBkdPPCNTvP5H5u0g/uJM2yTN83JxggiuA4IpPowzvq54wsfE
dBiIvfU8tb4gLx/4QfhJb2MoEICe6zDkvcgWWfo+DNj9Nrz5jngrMKBo2sxTGYzP+hYjMKrDoD0r
st2+nbX9g6s7npUWW+007s8+ykUeAGx07zb3cK/dWWNrGtA9J7hlLyV6XCcYI5xUJutn2Ifb91Wx
eR1UkwlWjg2VJqk/Fr6/cDvS9/guody3gm2PgsOnV2/YSBSv8UuApSnacL/xCp38a5A0E5kiIlCt
9/61ON/1lmAUFgh1hMHKNRf9pxMtkVrLQjk8nvultUKiZOrXJ/TDTiyELUhpCtIlyjFARI8cb6pT
VQLIl8Iz1jmEqJu1LEfJOlkzvEXbf5N+Sde0s2QzC+1UunCdEvH4/YxbbScLPUU3hLZAStCDJG2d
tw/7vTpjtFElx+5xWuxRORH7YuKibBD9Fw5EXSxqm4a/J0r7zBYMUoaQa3h0znwsceea+FZfjImT
i65IXvVTTQeLDXFbNZP4Up+d4tvg099S5GQJjdkzf89AqGGNKbrGikzEjonuGkLCeNAkBcXDCvqg
iYJ+U5C6/nluc0i7mIJrh9LPP0JTWU0wi9b99vgEbl2bey45H0Gj/PJLvRsgJPQR1Xivr4dtBkZo
mGsOgDyhBf1I1KJVtlepd+p2At6JgJViE1bU4m/uSxBjvXydm9NneZ3WAMUjwWoCsjXpdYobzPgO
qaPlr70aF1ZLMZ372QfQcfk4piZgI+px5Ztm3G/OeDtJFZ2Qg91+kWaAYS/ZVTsTZjfp2mYRdMM6
1TQK6j0ZYcFDKX5Dien7nnAM62/ekQ9LsYrYOFChS3MBTr7oIrFNi89rogRIx7p1g4Mr4eJ7VXk6
pq3kvdZkHzMMshVtcWPzZFPgH/jfZrJrI8+p4IKZDvSilB8Ca0EOpkCFMetlcMsoIXxm/fVHyGF7
bU8dUMqp6VkZgJAwG/eILQRaiMQydoWrf7zk3nYRulHOTf2SsdomEWNUduzJbVcQL3LJ/kMKuS8S
4l73kzDjqrV4FEOSzpwiZocHWzji7/te2rOlR8/5TwDkieFmOJnjv/GqCdA/k8yqZpJ5yfL0pPGy
qk4DQN60mhuqWeQ72wczGu1V7baFvQiu0ZVaIwVhqQ5KT9SkYuf+6h9howPoACW34VO6uaIxETZI
H/h7QGCkWFW++lNtmqrx/qUOOliVABbT0PeqlKo9qE6WMzyezkGXhvr0gg7VWDOCDOJRTIvOQOlZ
2w6ga1Fr+mhNYHixjp2EBkfgdOvtdbqpHJEsTs/DEBD+ilFfFi9FlfEBcIhG5gsqptdCanxW3oPV
hnCTU7L8+ASv08OQJzJVOf80cJbueUXJ0pK/9FFp8fF60+GSbd9L1nI892VcRrsdZXj12tqQh1Pl
VzZ3a3euu2A9R0SMKmoGsC/4XXor87/XKIv2WhA7trEyd7jRQuCyztwaAQsEzO4AI8TQrkTgSxB1
skZoqTL3reVO1HO4iciFsaERJD+ik2um8pzXfFD0cgklzOYNzOUTtACLP+nmVg1XJEF4g9/bzqSh
iYnpWDGfDQkK4PhM1dR1bpeWW+ehNh1zWFS5Y3tDNlZ3Pyo154Znha811ydCIPhWS1YDoGBx2j+b
Y5276HOeTLLBnRq7BTu0kTILjNmNCJaiAzeHtamaYNs45u8YiJC/ChZ/C5a/M4NRhNdv9szjC5K7
vkebuelvMboPrxySMre0eetiOooRIKbRyFLdBqfgUwMK7SBJnpIoF2/CSe7Uizoo+7nyZcniy+hj
NHCbExNPaUsp2VzZVw2j95C0b/CFPRxKwaBSen+ZcEl6lhsynWJaDvcM2oXPuX9uJVcwvnwvwkx7
z2IXAlGB1oh3RkQ74itUNMo+s8V7CW471TE3szd67zJsNn3uXuo4HUXZAL06kVejlcPcxmc2WYQt
i0q6a/rZJMvQam4Xn087Tud1nREedu5f6B+jP2cmZaquOX80LoZThoTkWkl6Dt7wOtC71TwX0ps5
mtclXabk1B4/HmXGr261EHOu6A41CtO8UB3+eazMd7HobeU4PxBho0vwTCTnmcs25BLCsypWVVRK
q3Xi6vCwsqK1osgzi6Iik3l22CnGvP68VKXHE5y4RDbj6I8NfO5W2B48hc80GSMLLTD6XKcJn1SQ
XRmLTVN2uh6H3D4cCnSS2aKtZxxevW9I5pL9Xf6VmQPs1quCnYvplbQFaL4moNZDeVoqLNI+L+wG
YclOy4feWentS4MzdNAGHsT541m9+u3IkPZOuIk4KEaZrZkiNM2FptM946zWCmiIWOeIVahOTjfd
Fj1ieMsYCgm8TmKXz8Rl1JuWdRjdI4ErQkITxBDIKhksstYdinU5Qrdn5bIMWozBcLm5jD22zYBF
lxPltExzfxyuntuRx3Hip9jTd6AltrmIdiiEayUSxbMBYD1AsW+mMLBX2hPP6iK3wOlDB/W9jW8a
L8IBSyE7RvUYi68RThLIIVUv++cubUXDv9d35Lo++qZ2n08Y7bGeiqSS4AANSYod13dTmsBsx1EV
LVIBGC7DUb6b4v+VF+GSr9r9Wuf+mluaQmp6RBGt4KteC8GkgK3fqEu8+in4qk9YOyLTBNfLFa2E
lpDLiRK1o2XW/rWi3Ky8Wcn/OjvLLnOeDEq2/jauDpehy6fvim2fke6McPkKIUYsCeKByzixeNaH
t79ZOVQGt8oYPjBQ7UUl9ehHH5OWH8TH3Vhh2cFeW8ijYOLhh+Nto1AvdJkatKMYWlI/p4B3oZar
5P/Wqv0SoJpT249+InUUNEoF2gTyE93+a2icYVKG3zTqu2AepuRxQW1ErENPcDXFJ0HRlkk/QaDj
Yp8UDp4ZF+UiDvXOg6Qi7n1S97elrJyRutENADHy2xwst3SPOoEHu4BaPtRUfU23YVh8XZOBbdgz
iBm6JZNVjYcgLVPzF5sY0uHWwGYYLudOHLrQ+o6FbvYVvONCnJLtGtAkeJiS1LXzJ6J/thFWTxOU
adpdDpGtgD4xQBaFc1NPUJu6hdYzGZ8xav+u+A4k06N/OgeORYPDb2vsIx6FqUfHuKbo6qw3NS9A
dew3z81zS5xW8skz9RMH8BMxUbcEBL6cQU72XQWjPPb6wITwMMoU/lWnAeQ8YYXSCYunZilnYd2q
UsDaj9eyj6RiZZW8sLaF8JmP6TKh/+Ayyffxgua8dsTca+wQsY7nQYfvE2tgJgNSX+vHDeWaH2n6
lSvnGxgfGS697CErYUQovvMv7gwVgYrWj8smMB1/6ZMs7VJ6NrjlbadOaQhzI8XJ4xdt8TkXLKOC
42mFyAjU8bOWSJfkaYH7Q42z7pQm+pQxupE2cPDjMpgKqQKD+FXU6MZZdwWtL3yXuzoUOJ06CcIv
R6O1JdePadi+MNsLGgohIFa3E4Ll8bx4jfXSdbCf1IbWQhwR5FRWk75Vxecv6wG9mMsENqoxlmp5
rfKhXOAUvkF0asUyeceHPvxu+W28hYHN9Y80zbToUYaBtVePC4aZ5ysrilqtHHet4MTylOoqu+Gn
OIyf83yzpCb/h79NOil66jEjimEPH7FzcU0zGCcD0f+j2dvzTJR2Yyuf/9Pq4qzdxoS73DL+n8Kd
Os8qTzs+FYGVH2KQFKc/NVm+NFb9b13ZoQobDbPO95tjkphw5VyYLcxWs8F6kHx2JiKyju8KuIA7
hxjrBNPk1xOvpr9GWNe9Q7x09diWBMTHIkiwArvz6LBxtp/347JUTSbbVnb2mkMGzrE2DV1Di7oz
9Ul9aYp6uTAdRARD6/3bb6zun4HGM6VnPDfVvTRnUAZNfEVPRFKRAosNH0E8y7/ITW+0pCgmSHY1
zgiRWgJUFPNEEfQbqUk9+cXUoiiEb99U1wOEmunyr1WFeyDwaxwqnT+/xGE/c/he4UgM1FszN9wX
O41mziEFGPuBIIIZtmWkftQ3HuI57xdnL0jnBaUuV3NdFwlY1qGhUKOVfudPhNQSH6yQbgDKZ1z2
YvdX1+qMPyS4g7uJVqOybHOGGEa3aTylKeIKuaO64vEFTXnoJMfqFNbyIEkB/1xnV8vPCkP8l2oS
Wl0Kr0LR+YFz3bop4K+2JIx8/sytebtj6n/+MMXgHuc3KnnTp9cMsZbj5qzd9pA/8apy5EAFxjmG
L1kMIDshp/FA9XjdAEqbTq1EMOVTt1hPLwGt7PLbHQZyxxiAsQC7V7IWf58vy6z8tcTjteBDR/dA
Qr65ZNWWISxhmHG4ze7kH6VLQKI1mqiyOxLDiCfP4oXQcQW3ArLu0lAAs/cd70Funacml9lbf5Ba
6J9kzj05Gz2aoqPIxpd+4y7ohVpVKYfynZaGsac+yaHgAfrWQadrZgW7LXq5TM11Vpp9uX8yeRgV
z7zA+BKZhKjibHrAT9EX7LV29IJRfGYcbcv4drWhYo1UnkWMv1e3vMQEqHLYdX7QSG56xXW9x8NJ
4icZ3lhPcHBV5ETAa2hUo8K8bKnTkckmdWLpPy5LnFbMfmNbish62KeswCfHVVRudKuSfqm/6IVt
fyU5MulwaG6auIf+XWmT6mw0pZWy0CtwQbkkJeKwvInnhYX7zSSULXgzcCW+g9llrjDdHPhKwHuh
QONkqJnmfcAVdYgvCscBmHoCn7eUTefTiLonEXw69M27UUkmHhWFomaOhr35ZgmLFfvyTAsOpvem
wwO7H40Fich0zPrhuXCV8zc8SiQmf/TrJVg6r9EwWjt6LvglsHwvAuHRbS1u+6+XdOVOtkBk+Bre
PJ0UNUGx1FVcPFg40+3BFb3LwK/aJ5SJOYh5KddA1B7Zg3wRkBg8q39lzVr/oUlfl2qnkUu3hVHn
e/bMJAdg6W2i1/euWo/we3WqUg4WgYi7/AH92uxrwKVk7APwaB/sAFkPTh1vVwGVQVwvlSjmqqYB
XMJs5tMLXfDCz5qQ3D/04/3AGkrtNj5W91FywTyTtlF4BxwhKVca1MS52u4w1xrUbJJiYqj+l74C
gR20rE74er0Ko1NZt+qnQe38cNt1KR8recPQk+h9aoVYHs9erJ0bc+9q7FvW6QaHz4RSHlY9jRc7
paxH0P1EKIjqWu5vo2B5Xor8jQ0OPI8mEcomJ2sE74hQgaT7IQiK5EjdGtnFQSwcFweS75a1VgxY
OamvR9pA26XJ09oA2Qd0jh73d/Zlr9pIrBM3y697sze5HTXro9Htl09tIIG7CkbBSv6tGgQfDTRh
k49RW+rEFrHtC6T0PYPPZA53RLzzWvYXMxNT3VzB4Oz8yHnzXA9TzQm/ulOuti/EXXKIn7mfEdNc
ItL6ars+CPDNMWHPajUdExocminmcBs6rBgRhhKFsLQfZzc1E4XoS0pSyYMXS2DEo99Btts4bDp1
CaKsoj87KgPJgF6tvL5CfiCLcwixkqlXHZi0TnW+xw8Py60Pthpf7KAR6apifuO/+X+JQy8fk55C
9/YI11QA3rMODqbc0vqz96M0pN2hpd8k+IR7aVYQSVtJM+o5XtNZbS2G6G+8ZD3pUtvjBlDdtO5I
GrcM9AGAZgYjHu7A5OPEQfESamLcWFHuR3om+IhDAkl4Vkk3ZJlNhSbrebkFq7oAsXtCq4GnqZ+Z
uHeUH2IzoGzVej+ARKVdOT9ybGkHCBMGEdmrwseoXo3D3KSsLQGKt4B4mnEcIaPKZu5GVNQd70Fk
zG/oTUPmoArYGFqkelJxcyqlt12xPY03DrWdVnVkUU0Kc4lRPJUz9ueZ2bwLyCSO+dKUmbv4xzs0
d849kydaFOQXQ3z+A98UJyHdiBJawxXX87MJJQi3K5ZVst32pFA8ZlVP7NFLDnzna6QXgIWJfgz9
/NZItgEIQhqipXTlVu4EAuOdZuU7nncqi9QK6tAfkznX8u0uwbqA7mXJ7+ot8pdvKlgmoDYVwUYe
LjXxI8/R7ZAsHj2oCzqFbGJLJ6y+7uIvppf6F34uCNFbWzJRpFEkbCBefzXCsXkVEThdUTt5M3qr
z4qiSG5tbY+bCmYUem+4UWvtdA4N2w0EBi+vIhQi3K5gBCcVD/zOS+YUEBjNHvRaU70KcJeMLRgo
n9RzmsF436iKycl/Cnw445dUtDosoWVYl6qSTYATcz1wWdl1TEf313BXti1c/N8GXnhFqhqjbZAz
EKcGgG4xUdR3SSpWmQBkfH/I4zWvBHWBy7R7dyMzgC+ZtDvfYxh/V5IY19m0JBzoaDqt171l7T4Z
fn3VKVo1s1tvXaQNsVvyl1ZYVO8/ZDzunjXRtYM5g0LfplZOE5KtwcA/Hw8Y6cFNwG0pb0G1jigh
dVxoL0ZSpu4JfmukNI/aMAluMdY/FFiBZiZlzk3qIecnMewo7Xb2/CfCkGTryn4YPJ33SDtYPvOB
ZQVg6ykDuTTLqvSnGYa8cEHbH875cVFEWZLeNuGzHRQC7Z3SKtN94WKpt7CJbi5Fm6RLh1eEH6Ph
GrooiQsShmgMn+Fr+bmm3Mpnc7U0/ScMM21gJsk8HxzG7I/eCbP1KoAUTCnUzaOyK5Qr9JRtGzBi
IXyeG9/d3zxMvcN6VdiPmP1mBSsOZCH/6nDsOmW0oX8waQOQXgcDkRDyfjPvuZr5YFMm5/pcRWsx
YiErsms998mG/ouzUVvCYaKhirA+NuJVBMLSCyXrh8ZDovD6IM8HIrsrodIalsXY7AUgf8V8ctkP
/tM1KQib/ErR9D4GcDIGRUN4uQzwGSvd2WXokd4/O74BWvIPhQpl4hvHMpsLHERb0XP5B/EvYNIa
QPD/svRn+k8NMedybS3CAdmI+tNEPm41PHxsAu0jjPNp0kQNiAX7lVhED2uz1UsjLV0GfK07YwhT
swwSBCWTbZyOAJu6pTGnlB/Eh6yQWEWT6YHZ0oHAspqvye67T53eWiQDEVcrdGXtYsAuvadqdx2D
UlrCnWvaa3ZeyLQlxRRI3zIbYPwGqcEBd48t+sndke0mPCrQlt4xQYqh7hNDqxWFroPvGC28pOL4
w0yET4EVfhAzeF9SwnXjARrEpDyxdSOHzU4O2EVua2DFe12SWD4Dw1OEIeAX8Cc63Insv2t6zfVl
FoBY0yQGWxmu2uemF3IcT+B+6DLi/UvWtnvAFpB1xPAo8zhVvoz+orDDX3hZIyzr5lq0WpU3REtP
wXEpmWrM8urTpyaVd6vmo2zxcnahup8W2+sh6v17rtHWC0nmggORV8YiWwL0MXwj6hQloxR1mTsq
hCRvrJEhIVJlA05qU3vS/jptlYDmxaY/PULeqOuvjAzh4gr1tbJwNiTAMg0WSHBwYrVFw1+mZiPw
PZ0JbLfYbQLLrKzlDUjFLw1eVfTpgUH4ffENZrzE6B0mSkqQ+RhIOA+AlKinUf9Uu3uANBZ4kAYH
fd+z5cUw3aO2WDBrffgZhXnN+/dIDnHTFYk4jGq0ujs7Eo2cEH1x+7z2cW3jkVdbYxL0RYwxD2KW
XiPrXqL3XoVVkOCd5gB4DD83tTtJ/j8lV7zFL0bocDq+t67WwdrOUauCqBoEsjJ3U0N9BdvhPc31
Z2jNGZdUoOLa2XRGTeLjeBLbuWLW0kSTaWe10Hk4aY2tY91Idn/aTi3XcTDrQH1mLFbJUZ4o1Ezp
PRYcTXy+zoiSK34GJyAnNImSpA9Md3erGdMDh6UFFCB/AnjPlHfJJX6sDA8dke7ntL9wvqf7pVt/
SeC1OdKRp0qzy+r62qFRObclI00tr+Ra+e1g3dzBxS7jCU7jDgC79Q331oyXMZlmWKE82Yw5rIw1
GgPHYUzU0F3HfLFDR9R48ou5cj+ejN79g//6ww1AYi2Yl4DUuWcaIauEjkqJiqYQP5n6xrXuuQrX
Bv3PeEiN1sL5R5TBuBzoILdpkbdlnPXy9tnpPBz8YPV6cqx8VR2Bcs5MGALbLaSr/aLr1eIXNlxS
hEtEaYaUAdBXpRDjMfCBKxY2v+00ICyFp7TrCTnj6Ql3UZw4S6rdU8HbS3bu6IceEGQiB0OSH1Bl
c0oBsxIkNcPkZarfxIUMNS8ioPs8HbcsnsHvWJ5uU6/2YnjcaVEAtcwDqjrVr6U7fORFvrZo6jtm
k41cQlgh5J2ROY0cYBk5zwq9UNO1sGVeKKUlyOnihP+hdw7IIGQLhVYcTQZOU+WEHrmFKyMkp3lz
9knuZI3lAFkxPUDgQaA2AlHs+5iiHH1q+lSSFiSZllVuCS7G35TOaf9Pe3S8f1SsE/KDS+MaLUy3
5ntvce4Ep1x3R1snoqq7nSHK3RxOtOWb+/f+0ztfiuN0feY2gSLBJ7MD0ZxeFL+bRtyRjwLCROp9
OcSco4iqK41jlhbYnqrtAcJ/XbF8t4Nq7fbyr42P4ij9XrsMXskenaY1/drJOZBKvP67+/luOv5a
5YyxJl0VgRM18bEEbsRjkingIMu6pbosRAYjl1P0hrEeF48Azl3p+piOey+ttogtWQvvuLKGnzJl
gqQtiNFM1RqlSDEPE4oV2Ydp08soJ9dGKlRtaMd4GculGL8zlUFsUqTN2qyx7tYFD8BMvlvkHftD
THHpwFygXUyc2RaBATh+FBDUl4174CRQUdD/5MyluGNhVTGhuov7L2knz2GXs1+rPXqqGs/Kd2UM
EJUwsf31d1xzGv2oRusfm0rQbrEJKQjBbzrcCJ9oqr+q693SGwQGuArraJMu648OzWbekF3rP9jc
AL4q6zyy1sUo8oH3S0ShFGSzX9waAdafCeQzv8NFky9T9vQfqkEnbCpWIBW9++jjvin2DxIWfnad
q+K2ps+dsZNLuScqeYlkZzYEwE3rPfiUYtPlyzYKlHOMzx2TDNfa//0es39rCNKQV5K7NhC3eszB
GlXY38hSr9JXrthRBMPW//m4afX4k+thfdFreV3+YVAlxV5HSMdx3JY0omUJWp5YcICfD3TYX8zT
9lX/oMZDmID+aFjihwWxEx1O3L3paj+OMYF9vG18cc43DYDE0qbGFp5vWMdUjXiemPiJaxM0onM7
lufZzP0+LR4OvPkY6nLF7XaQaVorzkVLm+Ab8fhJ59Ipc91e8Bi7UgFcQOQahqisB+poXh75ChdM
MQhb6sXICqTvro/9A+3CwCedH07erjX1z1H0Ex+qKvRpm3V/2bD5PHvUPeomzsn5CvEbKOhIsT5/
BwkKnUxtR71IFjcqvsITQVZYhS4VduX9LgzBAY37g51NyrB+ffyi9VOWrzoC3prMZ7YJemQ0ehqA
kvawCre3FcC12+1FobYgDFlgKQ3+e+TQGX2i5fgpDJcOFJDhJtou/QvQvAimaN8RHkAx5Gm1uMTw
TKeU955jjnRJEclw5n3h8/HJERPTOLZglBgis7aviwNvLFVO1wYJBm3ELAoXmCM8Q9vs793c79iI
eWa4+oAVu+5PkojhX53SGD+/lQyzBl6iSrrv2MYPsYS/11L2BSrOOkw7nbOOHdBsUs1j6ouef3pJ
O6m8eB3T5aH0mPebI0URzn87fm8D2IIvyME+sQ01ik6bOgbOo8kn+8uTkUzukD28Q22B78GItr1t
L7EpB7AI2I4KXrIpam/+jm9tuThKNh5M5YPwW4cvg6ZVym2ZD0gKxAKKPr0e3IQWdR7p0QGapgoL
rXGPljyLTZbAtdxvrzz04/La84aOAQYBvBkQsbmvcim9Z6n7LI6MmY4Bqz8sWMyYurnasV5k1Px/
ilVhlOU93yQpsyUjahSG9RvVL5JQbDadb4WyAelHgS5MxO7cklb1E9+s8/eXGJ+kmUZYC3olnT/z
n88lLv9SFJ6zqQXgCOztIFsMc3THYPMPBbSIofD/ZcJQN/abrWgEAiieVbuqyH4uuZmGntk4WPlz
GrxMtXppC8ktn5Joam4dJVwe0Ot/DqCT1V/ppvxSD5s6GFMDdti9OxpqCdUmC3jfSpYO6Q6r8jMX
SN3H1Q//GcEzQaPzDTkAO2xkfmz1HnRlP5oTaJsxVGr8dSB3e/wE47TfnjAd4ssF1KY4SttjxHzw
mAgcojXOHa8AlRXMEz38KJgfHZTZ20nru8C4R47LekVF5vCLjSWm98p+N7Eqi5GAfEL4P3BDNecy
v2f/bIOuyLkpAAG3aKk+24TMUQe3cEtZ8D6Rj0uH8TV+Af7EOvjcg1FdmD94PJOOoEU8JI0eCVen
3DmGkOZm+BRAduTsDOdXtlLxkyOozXmhL7iInOPYTaBofPqh3tcWSWbU0c+srtuCa/k+31RQa06V
ySzk+U2zS9M9ij5DOXUfxUg6VDpvjWZsHMycfF2871Xz0Cn2b0aexPKSiCFLvnB+RmUt6myZFNX2
9pfkyz3vZAC7keCa8KyuZO2uFwtRnUfyahLyXEAW84WEmaU4ZpjBfDvp36r/VIjkYdVw0pHyHGQv
18HS/tFZ1bF7X5so9vw6ZOe2/tuv4qubGJqC0jqskflz2pYLXzBMzgP9h9iNbu+D3EIpApwoAdor
3xbd7hdniNShFw7HSDf82gtX1xc2jZO23fXjG+Q0shY/PgQq8a0Roi2Ny7IUGtWVoZm5B4jzWTZM
rPN22Yd+aYCzxZ9yCwZHiNdCruE2z4hckQKEA/jsY0m4pbf3XC3g8znBtMxV3OioImAXmXR0luhh
BmynlaXLQ8cEruYWv0tWogvqoSPnLydW7jIVhez7rgAkjnmxfv9zllyuLmY/b8RxcHySDvBddHiK
XKKx9uew3VaWcRM4ss4pvDh4wvjM6OtUucf24n2kgm75qNLkxyf1LB+1HHapvG+j9vcKNvnvPtCm
HAsUb13ZXNux2B2tk1R2Ya18CqYLo0NObdbpAJzWcn1Maw2pglCVVZ19P/fRQlXEVi6jglpraCpX
qqLMc8lEam0liLqRPnvZF152oHUCAIjID0D+zCwwZCFeoXToOoaEEMJHI4qy3egVj+OWguNF2xmY
yOnfRx7AfHe5nMguoX84v+wsgZa7s2MJ7hXKLsrmpRgfqd27g7FiW4bZj6Yx4LupAdXok+ZGDNyO
/5Di7GZvyGegrnzPJ+ivD6K6lLghLaUcdhTaJmsufeH70FZvZ+EztDS4Zqky2nm6rcpBVgg4aiL9
7oS3RivnRpVduyYEptsjfxuljAA7cZye2Ly9XEpB8PaeZX+VSaY6ceavCYXAGTZBPY3NbCPBgDjm
5Ek9qxTn+vdQQGbF8pg26Bs4rhutn1BB4m4Nc6C81DuFz+InNlspzBCY3umXA/q68I75Fd8eLOST
j/PCTCI4iXAYgDeBV/dQkuXxRT8aFFBGfD0WfFrJrej4E5iFdtBb3uTG833a3zD39oj2Ofcnb87C
h4w9Q9XRCubqsWuyOQotMSliNyIuuQMM/qA+2WznlUIVPSMMyljq6YfgP699+rXsygHZxd0bevjG
T7cTrmV3uPSYuluw0cY3zJ5o5tcaAn7Bz8FWttRjsLRC3dkZuQEYGdp7AYQyEgbl7mbchPlvfJLr
b3X6Ke+srCQKXBHpxtvLV30FvyelqOtzu9wUbSdw+kHByNlXW2yShlFuFUF1U9DAt+zF9uMFdiJQ
YYAJ47AYziwpSfJEaWDGFMmQNLjY6VhQ47R3CWPph/DG+q4ihFG+NWr/lyllg3ffiUr0Tw83EAIr
1/kx+Wr8+j3Cv38cksfwVW080BoJ5RKKwY/ls43MytsWy42aawmIyDBePr2AnITgfGQ/4M+ADyKD
h4srr3QmicNftax40Lry4KgxbFzMFeYPGC0PjHqufrX2FfKKIIFjYdk7ox48b5Cr6OOsAIac77u5
QDRHI/dBkD24By6o2gN2xuNDei7aFcHw/JRbJh6WOnLlLPDDgLgvqYfpyt27S0Dvmvjv3oAAke4M
l34TU7LG9pL5ZG78VhtEbwcwrmM0KtknNUTLHV5ZhKSRjdM8X1UPrYPBQmmhISRAtAgR1whIo0JH
iJX4fyaq6vB5mKxYlo6m7tKwHQoq2+8DbbIjty3se2QVBUr/SQAxPtmQ20ZZq72DGqzy2j2Cmduz
MqR4mIyNeLHJD3eM7gz99QGUoCBuo+TqohY+vZsny/7i9t/9vxnn5mq+oMQInMc+dBeRzNORC2n7
2zR74R20Ow5U6n61iYGWAgCmYCdURjvhKYxrSPU3ydu59CHLLg1+zF3Q2CS/yslqP2VIzuujPMLp
ak7Dyi+qoc5MX38TDJNktv7RP2EqgHVLnXcOf+DeLfg4K3JUpz/bXgt2I9NimdjQUve/DN23xAjo
bpYQuNERtUp1C8RL/Q8R4gsr6Hmz9ByAEwMXMmRNIBgi7tUWx7983IdGyBUUO/d6OuL847D0CJJT
aRAbEx6pt+gHxQ+UaVQI0BAuCi39QWptVPM08WCPZxeWrfcHbBObp8WP7ie9ylFkfrnI9eOiO/KR
vGvGSVbxGpJc/o1W75dEOtv0lddgGik6htQJZQfjsup2cqv6mW/RmtYzfZrKknNjzfOgJw/jT7au
mA9YVC9ZS5gwHUnRxaSQt8G7DCNU/CyjmWIqJtYPt/4firD+VcAG8VYqq5BqcfEzIS1rcXvASHO4
aw5AU1hO8VtK1OECWkTrIH6c3LCBebQubKR8MxalrxVTR/1fhUG3DZgEKv7eFj8o6I5/j6j7zUNZ
12Dsz+byeWms3jU+IsyCJcTcD3Xw+TYKYmv98BzCzabii103KkYetfteexPUq7ZFFOorXSCHNyXV
/3Mv24Mw1XitowUJr8rNzFZUtwCHtbUvrMgTOhOU32u+TZBjrye9YwRZde/aVX1fIvLeqvqe1bDU
QTN95uClpvBdgJKdfSNkM6B2uRlATqurPSHTE5nHcVfvc4WsYC3ssErA5APr0aC+ZSkX6fR3Qc8r
UUQXLS7EUzalo72JQUasMC92bh5+XIftyKQAcwwFjBaATzbZBO3X59Z9reQ76miqpeNBtUHl2ZYH
o/ie9BIkgc794b+nGA3+C+nD01n2RuGyHZVYjjc71iXQhFO7r7QisVzyhrBnqVxUKpbe1HtQRqrX
szCgTpH2Rkt+2B/fxu9ip6AaxO3CQuzJ77PHSjnDyvsgCTzGa123jKzoxLdCoAzHU84FT9htwEGK
pDoPAvmO/ceR0EShhW6/Dnid4j6SoVSxqXIykcvgAtxtSNixJ9VNNTpXm79PpS/pF0hYfzKGn8xE
nD9aKnJmW+jaJfzMwzWzepivxqgY52lf2QA7cdGUdVHZfVW2BvOSHO6+duB7L0TYOT3NsLlRWlcv
+B6VROx517JGCHydTlG35S2kgPs3LIiBk4X1Ri/QGJBbat3NB4vIfIxTDAGszBtMhkLjojaBeTRJ
qT74NSXKpkPsAxAw3HaBwvBPwFxfjNRY83EzzeSVq9a5KWQqwczZWhy5eeZLcbTadv4d5TQP591c
cL5wb+ktIzLbQ9R85mjG9voGjBFH7NUzVJy3Q1yVGOG+DUrRW81Ody3lGhY4UuGAFGMs6u/6O8fm
jema7ZeuqZBzRBGodvlG7/JBEzJRo3Kwr+9Lnp22jCotqeroDF/4XFS8AnM8kvBRQOy+yJ8JHjhv
n8AeP19W13b6G8nMAL6Fm1et/CuYDaKKk+gUWrWrOUrXcXonFQgBZ7+d3cfQVNvGr5Lud2E3fuJP
XWD3LDHvDBveUOc670fa8RnScS/VZDF1hNlm7QskFCWygyffxCiI7RpcCBdMUxur8Exrwv2SLF1B
qWQbLgK1dW9V66CqWmYtMbHQutEPhA5mHzlFYjT5MqlYxvsC4Gm/xUZwGOKjHtZ/o+a5Ot8UBqrR
wurRTLWKfkTFvfbmt56nzBJSpBSXBVHDWJQEsF0wpvYCy+ZMs3cAQQBOUYEHqsa3I6FTpUcPW+5K
bFmRYoSXmPU4VBtiAsic7wJk6TxUhTOttYxNyyqmbKksnIKamg0plSGcXg6WuUZgyCPqpxmP5sIj
7vZffKVhMmnpALHjH5wB9eh6QLsDmn6YtGfVqNZ6+UKSLSkpL/tLZZ6BGRI1JMpILgwg4zEkwyy6
IIuaoOS3O/fJmDFU/voq/A04hwjamg3Vqu+c2Q7RTQCR8kvBBebHla8Mr4mzFVWvVTtCXp3Mz3Js
lV9zk6W2LuuhdBxJMlB4bREo485P4Vb6eFHQA3EqmjNWE7TNGQlo8KJE28Y/Z+gHIg8kBb3vQkMT
eLzw8+Wv+vY0OXDm47mKeZfRj6CBFhTk7pkWPDppdZ2KiFXuC+qhdt6upDFMhMOX255PTtTzt0uB
P1CNmqYGOJKNSBoNbJE/QvkPJmM27U+uAFrai4ip0JBp/l78H5pdzm9cTUQv4G4emOQGHZbadoFR
RRE9KMecukBxmtwq5xGw4K/jblttENvtOQXaBMsml55mob8d/yZ2rmDvcuWD38RrCWA54JZjGGLV
6yyK274cXHiOJqNgKS6bbRyD31lLD9ZPMRtYr+feRje+lirECpAzSgNec63Ozr7cgjl+2f1vu+t8
AUgI+XLtAaG8aq1Xake4IX5WuoWjLBUUnsWUmxMwbdEhuI6tqKpx+nPSDWZoq33prFlK2KtlRySp
AIifvZ8mtTwMxWxhu4oML7rxHlZPFHFEPOz3EFj/Ubmida92wqxzLsiZuIvIVhELxeeQkInSxUXS
eOMfRzxIRGJBVu0nzO626kngG1XQCzgiZ2ekWSAOhST/SVVv9HmTVP1RjDupU6Yrd6wyl8iEasbl
J+Rez61H4tz0aPJvR2wNyJxJ6Np6S7bNslBKNXiZgJHxe9Wu9L9G32E/djeIINzXywB2Ed05VdF4
T3/82CcIly1Bbtob5sgBGmyrJuONiouZWFZ6xH/iLyU+FUbYuM6FIJFjtJyhL9H+CSet0jNEAZZT
VL/9usSu4wRigvhbXqCWAbWdugutm7plEthbmf1blcweQPwAvwr+DKexi3NhZsEpDl5X4Di6Cuk8
i3qLckcMUbJrxiZaYUsonlXM4q2ltYWtmHJVZxuNaApB2w32vAMiXDTymZqrwLv48DvHBXcUADcR
aYUYwPUgTbdSIkCO8IajH/a/McOlTSFdLYdsZFoml7Y3tEv37pPoFQQ+537IvDIWs/S683wUdpS3
gnDnQKpQFrzFBmCaTTMPRu0jhoK++VFe9DtMZiiX0nsTho9VjEsQVbgWvcWjM3XGlUDoKvpYaFQQ
zt+qbh2nxW8tza7gEmXAtfzuZgYWxSk1QpKE88rcflHSGCpzgjtQ7fQq0IJ42XqVTCN8uJ2CVhi6
rSI6Gux9qCRycyV28WEvtbeJYu70083bk2Rpr9Fm0xcndSQNSi/sennStOkjr8EFvHw27Vc+zakK
1tBY0W1amMJwkL+1ABzAjLe9vDPu0QGzEtpPPB7Tu1k9tSSyEbsaFHihwEravEsYdbetIyzJG43e
YITQsiHKVo0dW+1FuN5Kfe7i55LMyv1KU95Khb/Io6nuI12zzjKd/dH/uMl5b/kFq5tyyNV2+9hV
IINjSdMmsIT2ofiyE9SJCAGRbF0MqSN37eJrKcCZT9tUSlK8PH61kX05IqCMamx2TQ4n+vUyQcVn
Uk4C5ZPRH+hPZEZDMXQiPndCYM1xfhjKyDqfxV9aXUMYM+ozyNr/oYkhU5wl1BNtzJIVu0X5FkNQ
Vyr3QkfTBOV5IZhzhLHSD0sgzKpTup5YE8jWFgxKGwWNkPe4cRm0K9WkzpHJ4ipvr+CA+knIZrAw
gBZAlFFw45OpsGfVaNHNJyn5HgnWXf1jcurbrtUaRxVrfXVHomrdYt2zZOlxLhVfsKGoce0l4kiL
XJ3YDNDffIYaL/d934wjcjSctEdXMHH4/OSWKMWyVlELmDXXViOY9/rjGnHfUTa3v2kS6LiiN3o2
PaNOIGjTwrjbUt5Q7w/XLlitdurRgQO2xqpREg4wGzZTGEGCHL/k4lPyZIMb0Kdox0bVmwTAnnb4
syHFlTWobNN4fz26WAwmFDI902mGMvGE0brB8hl+XXybPgKLVQpg+FfuLxXNmX/iQOqoUSChAY4z
o7w0ku563S9q9K/4iilN6SFNPzjTNDJmqvl+YqAFvHI5iPr8G289N1EUVX922nFFSzJkJ9/QWjYa
gUybhiySWe1MxrA4G9xziagRy2+f89/3MMpbl3J/d5HD9iaT40pnSQ1NZB7nFZQAHya8iv50c7Fj
RK9yZNLBCJRwbdlG6MY0bA+XfxCLZpZ38LeVt50lMQ9EVNWF3kEsG//NVlkHLQEbMzlqUVly2CvI
MrZNtOaMJCqQ37x1U5ruJYrz3BbxmIDWpGYuCMOHDIjGTZoX244FQINtc3/he3zUo65ah9iAMAab
QXHinIBSH0Q2IlX0WSFyS2h3YeqBwkSgPXblINvLEeNow/+vlUaimtpCqajyGGo1hAQm1HzbpGNP
plQE5+Agy9NTO/veGOnwK6lIqBesSxFQcBj4P3xumUILpFn33QfK1JwwLX2FnzqU0cKil4lXOoph
cVKMsd0F+Byf4/zG53WGn9Y9/eWmLUUAJXtlifFd8aOUg07+Ojny/EzYg/CDoQdjD430i9Zesx+N
Ve1mUCqGia5N+v8Ktxfwn+i6sVm+6BUlvHcUrhzGzYL4K6LCpJY5htUas8UcRT6Vf+H2jvGmunAF
Ri3DdwsXCEogRz54I55q7hjBivzaNc5pn9ASX0nJUUKelGWunJSl4HQwqlbY6xAYuGW3PU/8raxK
WZMIvj5FmIVPTRANu21osG76GTwdDTEtUqbm5zPCHjPKmEb37tJBL0VWO7ejDyCSMBkvjCYMSi7k
uAmc4OJvyXdq4YvfLcljiyzMtGvNr5GA8q7vaDA2GnN+NBGgwWV2nAO/F3mykN2G888xEHPVOMKP
Yo5CAEBhDLDk8RU8bX30cR7EVYEeoFSK5feZBd+A7NO26KVKESRVWjZeeFGl7ojmwdziUrYAXR8j
t2Uc6Pk+EjgZTfDBD9Nt4StMThFUMqJKep9qA//HiI2LfDMSTPM92E29ELiktc2X2oEnYnDYdKD3
tuwCkydk7tsLgqrf+wQoln640oquFeE8myOUN5rmUxP4apzeTGUd/3xPaR4WLw0tWXGpycIMbxRV
24HnKcQE9/Y9JWe1TARBtkYV28v2taJaZCsGs2juy9Zw9B3wdKoGcMlYiT/9uITSDWLrmwDPPT95
pat8B7h1tzB3Z3w0gTjf87XqEjJBuUAt67L9fhbSyP9oAXVxGJM7dKuD0UdcE6rB9wF4HW/P6/Py
nCqAq7iX4cX6Mf2Ji59T4iiYrrqbEaMCu3k5di8TJ3e72I+YV1hXdlojDSAtg/C9Tb86DZzY+WLu
3ZuF9HzqSkm31iu7ySFWCZ8zVAnlxbZOF4JuuZZmylwgk/CuH1IUb5EibU+i71v+HXLdvye8x50n
zbecFcUZ8BBkhqFmpTWwB5mnTAzpmKTSYZ6C/Qhf7DuK9K6DYb4QhXnzaSgEuTZ3DPHzBL28v93M
E89gg/qafq0OrPWWuuSw70vmhVsfDT7AoubvTGNpivRlu3Pf+7t95+3vJbQalmeBMCFJOOeqB7bQ
lgQ/pQtvSYjp3tliApiL5EGBO6Ak3AVphn56JqAHBkup3sfQkC0fsGGijkLfTXLQR3NwHvZeXRkr
SOEgCnCh4gF6lNy0Ltjkmf7w0aWAwiLW2eoEuwo9AM5DQ9Oo1dgLDquGQq2V/DtJNi9zwTTy2Lhb
qA7KBt6u2Sn43C/qgyGBgZjipUUfWlv9ZsARxHzNqaKb8wsvJGMxlnQ7+jQZh9TYBo4R0Bek+369
gOZKdlYbt+2xR1+AQ7VaOqwLfuxIfiF1TYNR9Lv4sATcJoDXK14/9Nd7iUvt08jSIvfdE87y/Ggw
EgTPhkHpA+SVvv0Qcci9c7Yvfa7/G3nb/kbwTaEztd4x3rGKD/8wLbKUWxk2rFpDKJB4Rd5cF4mq
nb6pbMeLCVsuPf/4BwBwIJoXbq82G6Ax+WxgL19aKlyn8DkjcWs8WEU8Qacs0GaImspPjtpp1IJR
yufvRDbpWzljAqK4M364Qrr6Bt25uPf6piSnE3UP0kjgAksxBm9dOgFqgRbyPXt42XczKQgoO2ml
1Q8Ruh01Y5kvv5yQjnpMP2HvW65f33s2EYPVhoxwZPJfxTIWu/hGvNxY4xx5dT0Ou6eN4VZ2zbkf
aCCiAvMyRsmT9slprwn0LcJq8rVxHKPzOrdYj8BeaHMpHDZgAvqhINnR21UxX0MXpcfMMcONKfjE
Jq8DDnhN4EiD3aqeY6Rt1jkToIVTGqkxfoMnvDOOc9slxl+gyTs5B2xXUf50hJ5Brwb5CrwCLHaG
RfjZNB2q2HHkQJyx3N42XyLZ6kbNhChzibeUqPsZ01iM+PKZSybHQgnJVVNf4zI9X5+e1kkPksru
2E9Ru0XbiNdRbvLzJRbxapWKJ2ZGpGuNhhRuwko4DE/EZmIpzaqV/a9iXkLG2u6ZrBEi+ec03t7Q
c5IoZ8fSFsqBvHzNat7CrXHfcsou5YEYNpulCrI/QfyurJ/N89YtV1KbpE3ip4F/QGL8ijimnl1w
Wdn0VDrlVX3dlcXv4DdzOYU9ovFPP14oBHd4YUATfdtS0HFf5b8pEYu1TMYV23r2OxaVV7EYWXGN
T7dl55n/ACIKgJdFp3Xtx6cADQwXQv3AmA/vnlktElhaZJjjHjIuVnqs2RgZj1ZPknJxx6HGav8B
dF2Je23rN7RoM43ZkomhY5Bl3hLLpAwrBpdhnA4fYqU4Q5Nl7kn7nevUTTkFK5a0Nyfq/WUD0K4d
SywerePzxxNLJ3vh8EYq1NAuaKBPC0btSr1Gl6hpKdVmlE5ewawHV4XhUlmXOnF27oH9oaWQcmSH
CFRxKwBpXjk6+uppYF0DJZpIsVt2GDlrykx/eAL6LsSczAIBLPgLJp0pFr/58AR82vTrOCwgQEZL
czmEPLkN5iQYOkymexyg1/FtAl3y3Iw67yBo5BOiMtg0dq6p0qK7B4t8Zc9t9/rtFrneHbdv8Axh
c67NYlEy++3loxka+riNhAEfV9AfPt+Cz1Vxipc35X/Pn5jKGfrSHAnSxnpheT81KClMRezifapM
JxKdIdW3PIyzD6YfdKPAQGHa/FtLwxT9h7aXyEQcaqM2UgZ7Nje+C/qQ+3SOI4Nq1OCj8j0jB+fn
dbcFzxG1NKUh1LfspooSRLU4saE8Qg4mMN0MmfBJIxRYWSUcbit/SdvWu7uxS3yy0UITc1CHmpp6
+hHCjCr0OSdzq0lqNHjXCuoMPBqFWF3PLC3a99HR74wdAYuWB5VllJYf6y4FSM0Jj9cR7SN6Vecm
lUVbxGIX6e5Bv+JxAxYfZ25O0+fVvy27ti6F9y2Go7u3UGxKo+QdW7Z5ilPOWtF8Z2V9DcKL9/yG
891AOoBqYYpjudNl4ArFI1NPrisbjP1Vki4ewO8/si0WLB5bycTdN8AhPplmk+OP8MKTMoGQhrVs
e/9XBV/UJ84KrGPToAk3eNrn6cxn22fZhVsTlaLg6igYWbn/DDLaXNae8BBs7+IV3L1xvQDtT9nF
sjQQHCbdsDIzRRQlBxQ0LL/2GathbgltCAh9g2AwOb8UBsbHSD9hOBR4awvaa7J8mwDBMfpwZHtT
SaFG0oQtFGQs20qZm5lkY/HUzGtn+kRjcU733iRE/mlZX8MwQHqYehKmQ1T7mNwmbY3BcWY+ICGz
fJekxY8JqP1I1k735fTEl0qVQtfJHc3vnvJK79/qyHuqwgWA3DEY24kmWqM29VrxMYv49g5V94pE
UjDDg2b+zFmAAD8QXBpISV8md7GTgNxot7hga+TfgzU1LuR7MJKENgBnSPVputJMvFNuyB/Ofseh
QUuqwT6zIE6KyioZxDyo79UA1MiEXGEnRYcQEZJovZVyt9IQHp39VqefljhhQ32pxpoj172Y6ptP
yqnQKPkOTcr2F3Y9kKPEsVEYMX2LHLEDDttmhY4HYkxKVs+dE1qbb/57S5L8Ind9LccpjHg0rhS7
608s7k0ZzC36t639CDo5MsWXYfVOOZqeLln47CRArSBI3SajFFqi5kNYu9wFn/At9QQt7WOZjL+W
nQZim4LazDzNTm0sokch+4i6WipNIyNStTyRYGDoiXpIFR8bMdeVPP8HIvTKb/YcQvbKwqj2IBwM
GPgOc71l+4mFBGRZtj+m2kutKHXlwcdnJ/ow33DNPf5I+mX4bMpXtDQGocHlSO7y5BqV99zr00y1
QGvIBvkCKsERRL+AJBpwddcZwEoLOBAkEhDjEO9dy3/cxVUDT69PbpB6dKfkUZpWvvAJzYYthJaM
B0g0DiwffYlT8XRsdqf2TrbkeSXdnLcQkA8Qqqv10J2wrWNQaq0WU+TWpmqbgub2osiDnArfeKVh
VyuWV2wasUwcFLeFnSwmnrdMEGOn05+A9fUqAGOYTrtD8DGFivqxmMQc8c9xRpytiX/BomefbT4x
R45mrofb8r67DP6iODFYSu11GKNk1ozhj3R/4egFK2wzemHrmlWMjDQ7GwanjdmofZDtlcIuiMFd
24c/lC48Sbyi/PXmKueJESKSNwlIZbqhhZp7o62KAX0HZMYL9UY5ZWwadZKACutUaXYqGGHMTXTL
etBeKOL8W33Gt6c73u4z4wbUcpN/oZ2p5gfuumSYCVs2ap7vPW++3C4lDNTD9X/a/xf9xig+hxI6
FNA3J8lQZYDX95GRuAzLVoBy8SSocuJgs+XlDvPjprlxRfzjRSD88UFpkoaZPAQ96WsSAVf++g0Y
Sr63qI/JyoMtBu6d7ELfpuJjFh/HUiYJ/gOvDQDOeEErnjeLWjJG0lH7feutu7/hSM42p5wDd3Wz
sQQP2oSrDWlYM7pWkbGHySsOoM17TPRSszzeBaLTHsvaxbk4qykReAwmT7uUygDCg+PN0sv/kwfa
4xQcg9Z/pz2FjYa/Pxg/n1yzArl2wQLT/SfseCGs5pbDTS5xXcgY9oi73fB+Yyoz4aRoqkuwVnCj
+E/c+pTYlaJjyWZblA/2yP6OznsNR6omkKwgGiXTgVEbkJJXI5O+3MGIFLDgykYlWYsO9JTb/ivU
cr2mqZgOj/Ck5rz/xkkQ+d3drNK7dmO5jT0cf3KNQWNJVIo7BPkGsfR34JwriuNTyWh5QE9rUkSA
GQXpF4t+2qelyvb16SvhJGuyBIA9C6ShvI0aVdM32QO+5qYDaRGTbf6Mtil70b31pOzIJ708JXiN
/x1G9yO+gk/vPjIn0A6K3r2Sorwqi0OawuVzRrO4tZG5RSeBnhwHdLuSeAV8Ycvtidqyou/oc8Xe
zH1NaTHMZbYwiGQBTMeO+I4yMJiLlqcZ043gpbNDTooSDXGTqy9MKE/t79OiLBCq72uh5ZVJslP/
SAFs02jLLiBSuA8aQwejuuf5SfatT9axIEOvV6RO91HQxdwMfOLQPPDqMyGfm1PbbOeAUfbNkU92
psOF9b/FtqdByYOHILTla1N2QxUBivNqcjjtosXFjGR3ZY1iIaFEOpUtUWAeP36Lmz2YuoqxswCv
Y7Q7U6KjhzW5YyUGutlLlEqDu9D/jvZYYofVtSIltm88HtxD6H9MeoqmH852U+CkupUcX+KXwScv
k9lJPd+crnszobJ5sLBqiVbUyR+keDmD69BynkdX8oG5ExE9uDOXSVJZCtirecSXmyzrYgseOy17
Azfxmn/d3Zpzhmq9uolR4z1Bxkt+IqCmFHKq/6JLf2zAYkhKd3W+AsGeDzlQ4Kp5NU5ddPtzgPVJ
CNmM73u/oyRn5nO7+KVI3/ChD9RaL6MwtEeU9tjNdF+QGzQN7uSmKFL+ymeQQZAqFCtsCbbCTg5Z
Eb6IEPJokKhm62Cc4AZ8TsLM+t5WqwvG/SdjS3y1j0wu8oZPYdFLKkC9w8li/Ro81kk0rFpIHKir
2r9t1HrY3Eam3cU8p0BCOngJsMz3gHnNONabNlBeNatIReimOAIOMJby5w6fB5rSXOTfOfBFEl42
Xto4OHF6sPnALU3C256l6VvTMOs1IsjnKX1BL1XbH/xomf6QTXYXhn7sqhbLyPidMjcTARcV/mbk
5tQoiFWwWN5q6NeIF0p3ACYjyuSJBfCaFmwbyUESQF03cNEfVRNwX24kZdMLa+5fP9NIRZBpqXdp
qa+3WCWUxBHJgUXvEe62IJb3oUhIRfvRkOd7DeF29eSL71BZaaeqyBX72dnu9cxbAGElHmTwZrdT
Nt2dk3MHZgnMItTH58JnLkxHuMm3856BFH/+MbEvehrIP/VOsD8icyHs4ITbJv0GO4h5rMNBn7JG
lqpE5Zblg9q5jNYRgEu86qgzcefyExkpb+JQtI7p83KKfj24mKkky5iY2wuQi+S2tIpKZbixEH4U
VjKgXdUkG6x8gUpVLplgJOm68VPCr8NID1sKgYTh2PbjyzgEERUGT4C04NQdzOGvT3GEYLfFcAGa
tiPzsEN6NQPiJEuJr7K0+G0uZ6uazWfcpdk74TJmwynzHx93bln2XsECcswxZfA5sAzEpN5Zi5TM
AXIEG0gPzWxounLOSEnJRk/HlVuJHjbqsaqEoFIA0lO/BltL3Z/phewTDsAb/Kh6vF/PV3DNY8fK
cSuieX38vgdmxN4Xkfu/lGI8tBq3e9XhWasK4MkxtrkE7EzkVSgjS9nrXqmNmlGkuYJRuK8h64uN
pp47DGZCkmS6iflBruO2LUhWSHbTvpoaBV8yJKDdXr92nI5pKbWJMp49caZGiWXXCROPzC/QFbgd
Q8ku79aXc173ZG7EmgQ8ZTguEYEtYb8XzLshJ/NCBhOaxzNpnkc+h4CttLmCKpUrVULaxaUbOjtP
H7ny7tPuqtawqyJ1c+IvUtw26msJCONTFtqnOPluRdz3Ac1ojCIK3qt8d02y+Q6UmoX/r6D6updL
fcdJMHj/hwlNczKlThjjKS5KzqaL2k+zCUPJ/ZGrJAenmqldcXtXbJ2+FVJ+14ugtI+1jPCaVrKd
KFx7FatpZ3dq0I5INq9kVAQfksMJBnb/jF+rDAuHa/T7HhCMrIfq4jZofq6uSbXClOfLc4xdOtbC
GCFfjj1DgvVyErH1421h3MK03ytDiXOEhQ0/qMi6vWHzxLY32V/ud4QFlBscmLM5JtTxzU1BThVQ
lWVY1Z7l8+JpR8D5QLWRt0L4ktCA6/y07MeVjI4x5eHWG5A6YnmUu+bOM2X4j4h9BVCgxKjWvNIX
gQx3LXYTueOv4UjNK5Qd6XTyPMf8VVqh2qt0ApqBVl4VWCs6nzKqvMtC7E+FG/2w9Gj4zBZ8YHwf
uNXcojKxg1oPvvcWasnDqxdelRkYV+XFUAZ4HvYcHcMZuPLcCqQ4TLQBj3GvQLVlNemcE/b7IYWR
ZZhOjrom3bLsaKMqu4lMdRcGifOFPY7EMM384Y6kO/fYl+R7YCtfJYDhHWiHh27y/Nv5srKOmVTD
k2EGyB0AdyEEKOXlYeuqVpdhjfUyOF7w3hFFTCqoV0buyoEg6zVu5GiCkDgbd3q4NA71E77b0Nlo
BCLIN1K5KnUwUrlyCIucu+gPL3zJk4RgoYPPULRzUZG6C0SEkX9Z4HnV530fjTN7Q/izXynDnHcZ
q4uPM0ZU/+T6sWUVyJLx28gPwQBDtPcSSldhi7S4hSnAGckS07IVQ7mjpLDIvfK0aDZT3iKwh+VS
cxEV1n2I28/hAW/x6kVAH+JwPjj6c6DGDwzOiOHNAfy8RDKH+R56TSH/NJMYp/ImCqZ12nsgPwAw
fy2zBFUyjHY5ejmza9yQv2yTzesNS45U3EpSMZELZpCc47UZVZEN4xGRb5TOsuNSai3gVlw3vNDT
lLel94k8Nsb1tlNasNRkHYEZ5h0ryExWInJkaw0YQtphW+3v8mkwVOyyKIyR+eS8nVyjH9eIifxp
Iq5ILZma0zZsZCNx60FwkHcSbj3yDmIn+piqb+24hSd4YQ5ebiXA/b7FAK5pgSOHm/ke3aN/Hi4P
Xm+W3TlfISFV3jaWaDZYm2TC77Ni4+TjBzfgSuq405JFpCGkCSF0oZlH4Egjqlq2km0alJvIiHdi
IsK+U5bgze2mrVS1ZeqU5xubn0x5wQmLs6rJJafrc6wOJfmbQuD4xh2vmhstMgr06c8pW5x47JRA
jW7BM+LPiaAtrB3LMTWq2137tAK/W3x/mzVXgBYLIclqFa5yZ0RxUGBK1E2+d44mVY7uJcXkAJNl
IE3vlqf173Fk/U4EMB3CLpgr+JcLNASE53m11KyfVaECla1FyhJ6wNRqlTuGpPCP/YwdYeV9Oi29
3/9pV0YcnXs6GcuBCRew+M4aMLWWj1ct4hwu/qa1AXFzbNkytoZVFoVidPRwnGe5o635drvWetzC
cD7CqGd8YmDM9UP+oOJSqngoyWGTtq5SFZrQqZ79kcUWIlcJigHp/YewZtZMmGRrDMjzorST4Ga1
wReosueY3JIyeeebFJowpRdcB+u7v+rHucFrooS31aigfBGl2ZdFTWiTykAbOLZ6y8HhyfeAF6J3
Hk6yvLLMhhwNMfVUIKUBg5yAsIfzk1cgc2d7CoHt7ITNvVXMCaefWNo9oCURU7avXSwzcm8kkYFI
QxI+4MmvxP6B9fGzYNeV/58IbCdbmzdCM+Pj5wrylwuzqHSLgdyDlE9VNCzXRri8r3MSCqk/3AmB
Ul8qpOWjIjbKo9VVZFsjSweKAYZHaPLlJU+5Mkx4a2g2eqLzkLUekUlTvo0OX8S4dnVk52sFb3MF
qParo2ryFXUIT/qT5D+j2tB1uyMR7WEluv61wPXLK1XPeNH0ygTrLlXlPFz4XO7R4y1SbEtIC4qV
fGtyfdPJxB+OynWDy9Io2A0HgzsM8JHxUuiHmSHxjGlEx1V4yLT6raJOOrdX5vWOo3q9h/Fnu1r0
/JFq/5Skgd7kJq5gcd3c4TCmfG6gRPzo/HYBWPtpL97xONlXNaRlcjOea2mJ5GC9qUS2vdcgLHLu
PQoqb03ENjRbExfJovZpP9CryQCTa6umZH3ffQ/ZxbbcUGSFWpcFUjvDy3CWaUgTCSe7jGTQQx+4
rSvURBGLqLTCByE1fxoXt0i13u8jwl7dkjshWWlT8X3+L77eG3lu0TwaF1xHESTX65U3QI7mvhtl
bEmS7wrsNC+1lDs5rtaFiiduO/Zweuebe0Y1ySG7I2wW3rW/3tad3F/Kq/0qGrAyEKcQ5h/p0Gpo
TgmEJlTFFermnXNbcUK3Q0Xh6sk+i+yZc8zV5EzPOHs5JXfSLAIVrvgrLaykyH4fWLDXYpxD0I/6
2hOySvay4lOIVQOWuBGKSyQdpiguX568u1r1DFGYFvl0o61GSKJodMiM39arCVrzXt6iuV3w8EfH
FcDEPaLoiloZO7gre3+BiwEKXWuI+1YD8is6zShZyGmF3h8ZW5qUNAlNXryeZa92uYPoDbQIHnbr
Ky/wx7gncXkP5XGH6BvKNfxTyvskcMNr6x3wxmt7MKQ0H+BBh4NTCCe88YEii0rDTCjTzrixt3s=
`protect end_protected

