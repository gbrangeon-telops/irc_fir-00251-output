

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Jjl8vAn2UJruW+pwbvMAIo6yT6bQgTl9+ZqbT+VaAP/dcMa9HxI5w52bG1uOMJkKjbI3shaTb5QH
+WA4TEmwBA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
jY7USlQiP9PR+LALAEYZsrKak9VnF4tfhT9SQb5jLUPXs+eC5ZbIVQkPjdV+4wzhB7b7ai6shnHa
gEu6kUZZsMTRIotEQn7SVZESTAIMCGAU4lDLU7RT30ySc+gN3y2heOoScYVxVF3kYNcbErB9g4iU
iZLVkq3ZU0fP1VLA30w=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
W97r968B0QPwlTs1emSg8mtee0qHNpQ+/n5wfXS0R66Akqy90VsNXhnqLJjbnGJNqaGSMTKCRNVS
ox1Z0rkuemlJn0dMgZtmRgHM/NeyMTSbsBwVvTSeFdA56k6PzciIIQ1S8150Bxbexnd+b7l/UMK+
JO8+KzzHPEIPqou3srZGn9dog9HSSfTUIqvBgloCeGmDxxwlsFwQ2VsrffuE8mB5Kk9lHG/A3rMw
tbJURgYaS/b69KLL9Kc/urEgbRWHU1HQCQDL4hSKE79WXE68MZJ00kcWMfNfAOR1zytQecSerjXJ
iVVvnEzEtzUejpnuhHCRhS+b62dMTzf5a1Q4Dw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
l6IXa1kcvqxcIuqXI9bELoLDvGs5XxFfhbXxOKBitloxuDBS5IYgW7AXksTedGB5rM+6jbAr+PVa
4ykVDtx+9n1RZQ3HKQZNsRywuW0+Fcm/MhmC5isxnEClP56JmzAEyD9l7nmy9JJJI11qQTy86iSs
hkUJMmO3Ph4Kz8ptLn0=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
gEbAM0PoYz0kTXyuDtZRhRtQJeO0ezbVNuHzWd2Q6Djxe3WZnx453sNsfBBqykQPTu/zHrWi/wfe
VIPTt4c20XjDHHTidMXhf5YGMYpytIjNmzV4g6PhJehJgJTQj+T/bAmaDaXLcqMDTjUNont0w58X
XTjVYtxQgjqcVftNf5PS5GCVpRxSTsKbT4CfmHhBwwsNC5rLtE2tRCpmB6tKw/7xf8VLLD8a23zt
cVvVNX0bw3bWCGFmWZjC/1fhYI19WFrjQO9Y/0zq8T/b6JCoxXV2HE4Z2dJ8uXvV5GV8EStC7VCB
DhBS/R4IfNLPojIIJPxvrbzkKlmuEkhgwflRRQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 57936)
`protect data_block
DqjfwJ4Jf2IG01gq5GJ7K3wRF0TCOw9rPS4myZ9mre7SHP3FqAcmzLFN8BhTodduyvy5Vjjb8xl1
zPQtB3Q7OqaAV0wvgQe0KKEuH/BJi0qiguGEwDfCUaY235bGfgqkXX/y2UM0Fs1+liv/3koDxNGh
0lROMHQ7bsnJ+z2HJAz5XTSBjr1anODCHyN2TPLsEfAAQ3HFkOQqbaeFECN7U+o4Hc5UFXjrC185
RiLYkZVyrP7uP0JJTXmllpoLtItDusQ3pRKo5LIKF75qR8GtFt5uETbStWQQ32luZWYj2spdZNLj
ZKkWvBSfe5ZjseNyR7QAWSbyAYePdyETfreTCyDq40cU38HRM/4O8aVIIRIUJeaAojQl8PWfZWnx
wUHyZW2LzitdTlXn6liNz1bjA56u+DCQKmTSLZzS14Oj8lojcR7cczIfJI/Hy0ZYqxZKpKOUxPHe
ek9kkWIU06f18om/NjJds8R8XxYQas7HW8b0LHm2P7apQo81lLERAcpbNL6nsSBptMCbEvW1zrPw
OWLVxTAtON6YpdrfsV9hoDSuLXs0DkYs54DPRFhQdAx3CIy6xqBi4lAby3cHibgEHSgnoGPWCgSQ
4yaoe//Q7oeMEZdzb+dBLiQVAQdZcisjYHpU3qCiJWBcw/qJWJEmBizqnxZQYZkC3nQZHzhUsAQW
nsmhswt+UwU69hRM27yzVqY2ocLp0kJ5lS6uyZoGFtLaItnqCj8tbpzxE/51hhnhwl5YMd2D1/rR
DwlEgtaxNXGJDSoibkWYp13q/Awb9T5jHp0xu2gdix7jfOl5qX/BLEk1KqpegehWjMSRN/lluS03
Ql78MUJJ+4+FLEupePvRMUQGlsvG32akRDVKVL9Y/i9gDd8VsQFbLIt91s7PKxZc9niJA+cvpH8H
+4B+ZxyFb1HGLA5OCn9tJTku/W7/eYW13AxQtutSNBw3+f37Jgrk1GJMDIP3H4atYqDp4ciwn8ox
X0kWv+GMVZJnhTxELH1xihhJ38Xj+8hqNmBIPfLyrCUFU3uPFdNS0kWz75k7dAHTU0Epsu0AsXqi
jwIs6PPlI8VvO1omFpSoY5Oa7sBPAyIhcxebQKnoJHBQiquS8sJOFSxgTU9/HXAaS+2fSG2X2RH6
BYzHEqXQANIyeu0ZbpkwQmvi+Fa5V9zW3BdyB0zMRs3wEhzRGWdiIED3pMK0Ia794L1uUK1fhu9F
G9jEqpMKLAGE1IzVJVUVHK20NXV/NDBM2JUvOJMh1idrxaFaMDhjmlBfah7m5aKgm+UnJTY1AC/N
jYNbRBdwq3A10jXKLTA6oYkVQNQQpW0Gu6BChBih3D2k1bG4F2K3XzhppzT3Jf6hWcruXYRhvSC0
WrlxI9wSM0l8rRnYhxGlAypn1ejW92BHal/oSMoLN738XDWBzlqdXe33IlEZAHrcFdnYKGyG64xd
PGwCCxRs2D8uzaPgvovYOp9usT1wt0JBHKwbGadj6hjGyOk9bYxMppF1ZOl5zcjjldj391mgexOU
i1N1WcaswYDDSJzTpwesuxuOsGojsaCVrlG7m/N3OMtlRW7kK09wMbcrqD/i1usndC0vaayerRV+
ZEFGdridmc8ABirxKZ78JNDCLE9u121HhMKdugUOwnsImnqU/69IGfgGM2uB0srFfnFm1ylmV6s6
ETQWO0ePm6EBUoEkrfwee7lfMsHzZZQpo4kLCd0OStB2S4rmJlW5cHfxQ3rgBgfdY3Lh4KQ3v9yg
efUJuaEiPk54r0HueaYZariMyrEix2sofDGAjtql7MFINs9IABiocemzFby3n/GSMH7pun8ESzGX
lnfolSrfXxDuRpYNFHTGJeY5mlTPeq/2b8I+ZTTVx86NeSdDlEAfKjSM0nSuJErFt1JYHLL6xsRs
gDAoVFHtq0DYgptMRIC2q2NxmssQuDvDyRArF2DbMHzJCnGAwxNwcpkd8AhJyTGh/DLYJ/9CuLlw
UpqFC3W6MhoKsfv9AjDBZFZGN5t19A3W9wyhhm6NhhpnLZYMMtH0/DkuYR4vb9++jaWA9JU4on9d
tlKm4UdN1VmUaVWyn0eqpcu2BNaGQwSUEgysAfu7+96BTwcQ2SbvzEy51ns+XIH26eD3mqr+2v9d
xP4IvAMmQKTbcUke2407e4buqdbl1VR0Ibchbx6u/7atLWPoHXKf3alHPTc438VTiA3d1iROf6aP
ocfKLYV9+DFIu/5TRW51jExJ1FBqS7TVj2xMdvkdL4SXT+OwNe5JyGeeMsfYQ3yxFCiQlxuIpax0
94/NMLjtJ9TDaSVmZ4paPGKEfNkokXq3l1sL8GclEzDGTF5h0OKu2pwBiSca+5j1j/bZdUwipVyn
6foG3MVRx9Bypi37N54oA5zel679mqYuqetk7rp0CagNzpOTcdbQOV0Oswbd2c5LutnHZmxfhv6q
KtdjwVvX/p5E65Om8RX4uJh66ose3h/z0x8SWsux8RQQg1QeiI4j9MdYEyLK1d8RzOPuxtStrFGP
9mUm0XrXKo2WVozyYbtZge11HxTDfucFrYv+KomXiCdtWoB68zb1TohCfraJmEPMMoan9u4HyOKD
ZibwgyQNJXyKVdCm3k1hnwvk+yBZZ+kkU0AjgNYXvN259QXQIedDs1yar/knb3flsIT+7D531Fyh
8m3HQNIGxufqhTKHzeUlY0RVYmtGXT5HB3n/vYakW6GZt1/J3W45gfNRyBLn9R3oajqqnUAaENQt
emUO5mIphcL+cberjILJs0xfIryBpyk33YofnDniyPSmsuNkVErwfN2LvKf+CLS6b7qQFiiTrDG1
SOurvejRh7XuOVRy2D84mNlM7qVzbxzG/ExpOVqtjdglrq7PgZJ47xf5iUtX5WyxJLjn/uNRtYu7
mg7cKa0FTW8TfXzeapHejo4XGGp5AuD5xpcJrvkV8mYrTFYnm3n+GNH3EJmwgUG7Am1DdxnSmVzr
c2k8t2cdQ91FX/fJXt4ltww7+2J8yHBIXGaKNT9muOG1McbZB9uicj7LSFBc/FmmPpPS8yh+YaOH
27jcxu+Tx281qPYQRW9WXzmm/Gv0JPBu2h0hgK5UZz5/GAax1qEDtuZreMDKtVhGat6unbkMyaDi
b3FRoorMCiL7GqJNdJeGG0EvICn5uKWzKKM8P++pGaodOPdmIkQ/iwnBKsY9rCoKVk+mjpDwQ6nx
9vx6tPPa5C86m/4Ui36mc3dEPzk8C9pTkhYW+X1bSHFGh85hwwL3ufGvmEJ0bO5enEkH1QuRPguV
XDQMvdt1f+vBR7f4tn0tcDt/RXSApF86/DTH0Fz8F96gJDrMGqgQ5G7jX6yQMDe2oqw/cX8FFy+9
gKA4QdP+mJsSC+GusaRmW3ldyYR8co8OpfVGJLUkhLaGdXVBk8FVBEQovnz057A4U3reVUsuBFEq
RA4m5ViXffeYdWe9+ka0RgVKRk6a4dpTDUCdZ6EjX7OqSyLIgudhiBK4Kyp99HiVR+4OFwgcnxh5
jWzjh2vvEvU2FTpfWebx8Z7IbhBEKV/XI84N1lotsgS0U2v4eQtFT043d+ItnC6LDmqzvlzXDZbk
nJZf+OTpyzVyRM6k2yWQG2qMxRahiZPoxyHlJvcQhouviiU/SsYdiq4UMam+KIpe5kye+F0J3jPQ
uO2z4a/fF2ylqVYRSruMiSYvZA+oZJwXXUUGM4KTKCo/viu9fySl7zFyFnHJkcZLPxqTMidqyIxj
aGKvDCvbr4AvXyCCUmJIvoQ8sbZYYqEfDy177VOpFlTSK+D4uebnHVKe9lD5QLJsXeQXe53GYxSx
5wrQFQTObWouUKBG1uaKcRr0P0Z7clB3LnaXgzJRvQT7UCMWZMQJSWGMiBVuWIrA9L0clAbHF+Ek
tsgjbaCnAaWQNuzdFyRxPt8/QZUsMMEBVUkpZvgS3w8KHGWbIGWq1LnxiVq/t4VoK6CE2/yVELlx
t1oAQ2dDhJah7a3aa39oWgzCIQ7zCvJK8941BB+NSldgWQHVbqtvbyKObVikcdaCtmYWoHiCOGm5
VN4g1b0ABvVx2m0YPkFkOx+1/c3IKE3V494NXNFmtBkwDWo/SLTYWSIARSYJdpSpygryuFEPwx8G
WP/usK51gPe61+npUZVFgPvslBGrRdMQWYvBGriI0+OdYl2IxBL/TsHCndJ21vTw3Y0n2yuV6vg/
3ghkMjmRBcz6XHr4fq1/bAa0x5fkYBNEJBxBCpybrLNF5xW+0+VEHjka2rmLa1IvM/d2Vw7RPPhN
E2S6lV18uI4p1iSFda+GLxnUSUsnPE2t5jWBBIWBdnCZVuYGqazAbt4ZaP0D6jxlVNIHrIXyZm1H
GY6jv2lHeajpGLUvyGpt4NNx85AY+7UPWnZUn2IbgLNUSST1BmOTrC/3qiFgRBD76zB49GhtjmlH
cEGWON+UdUMiluYDMV0ISZ8Ss86tk2n2C9nFow2vJPy0zCW+DxA/YdgctZVNxgwdLhnnajLfDkXB
kCv9UPEaggC/kMUJyOeOczt6DGJbcaEzB1qVl53yu4lKl8U9rQ0ZfzJcU6NJ1VNtkt9Tmh+1RRZ5
A/iJBBnQL8XVcLArKM0mu/VC6cIshT+OVN1K4seddFCwXNvdwzPkcjyr9xnwCM7BXpH8CyMJkfUM
yXCprjK9h1cg79iNXihpe2a68Vx9FuVg2U9s0R9fJ0AfFkVG2/BUTWe+pDaCcbSxx9g1u1tHTGB1
51Vtqgu84OcRMcnOgROknSfGWCZ6Ar+kagO/vvL/6SApqaXz4JXwRIsp/pf6TvmkIGocoRFBt2Y/
ZsxDIsfm4rs0Nrj7ADY0Enc9X71TM4aIhnq5N5r/DxyJoRyIroxp9GkzyiKViwpyLZdvejeSaqet
zMVP2/n1OKdvtQyZ314mdZJ2iLhjTpe/GojwG3ZQ5HJk319T7UHiBct14foJG8T29S0adJv3nIio
Q3oHegxaFLUv+wYWe1tPwwoAMNmHz7V4qk/a7Y0M4aSpP/GfiAbK2N7d18t2QwXk4AsmRx2FCmMo
/L1az/2gJJyClYULdx/0l8lmZpKcei03/RjgHi/UOpnfjN4dZknwsl4Gr22JJ+RxR0szHimNGznk
GDlUBDGsyloNFK9PkpnCpIc7izC5kVWSdn2/8ireYlGpdq4KRLrud5l1CyRqHymZfaGwJdWXyiKo
uasu4fk2Uj786WtvRiCs2IOUzeFUQ/qNGtP6OxDPjbFsc5b9Ct6cBp4Cg300F8Iwy45msabvEojW
suW6plyaysj2HsuBGND5H1ZZLz408qt79YsbRQM9IYdUvAEToIEhW+Dg1PisKclDMf3DH6oMv81S
kxM/odr3lWFBpxGsMliSo5c+4G6cxLaPzoR/MoxXuBk1WlrbpHQvmrmE3FbGsjBXS9FQWfbx+Tbz
IhQPt0/fRSVnlPr9wspngpAwKDjgaeZOIwnB9bxdo15NWBjvgp91R8/Wm1OXbGyrwwIkGh3rZ3l5
urqAmJXj9qGXCdU1eob1tuo47yPfQ1UnRRxoKQ65DHDoFg6Ngb/BymDGs5astDnzViNEnlZqv8aa
qBUs5YtE0TSM0YI0v6zi89ip4YxGXLWL+xRgUK8fHamdEG761MramXV8XOSjfLID3VXMIWBUC9Kk
EgkOQjXVlJB8EqVYQTaVL0hccRwKsDIab4J2fMhlRFzN+KvPIchHaRjsk2pPvOt2GYO9nLGXMdSC
alc4NBCZaP4uE84srnm9JqJ40UUmQGhvFv4Ohxp8KHGBEL/xPp8L9EmNGdTj2y6OJmq9mhq74y5R
ulvlsGwreX/VaUXS0cRmbmHQP7vTqVdmBNruA9fzT68aNEE0XKW5/lYJdePddpHZvvNbodhXdnkJ
2PgPPeYSMRaPbon9J3yJI5VKalo23GEc6IUs6XxOeV5ZqwOI3RntGcHs88VY755isFAkdUNPYC12
CTRpEBfB+CkKPmsn1G4cvYAXDCO0Teg/adN8f1lsq9GMATEZ7YM/iJr5B0yW0mq1mc8o4A6Ny/8+
5erWkOgJxsVFcKvbA6KcjdWx4WIbdKJ7sZlAeCyPKsB5zTNSp/ToGEJZpoq+Abnz5FP+6Zrc5nAs
b3VWyzCB6kpk8l5RrQU+axu44Hg29N+LmoSvNu/Gt6sd5+cdtgkbHBlPXDqV/nLXYIUPQz4/xngq
GrIAmGxvcb0EoKXyurUr5x2mNvp4SkKlMVBHjHBQj1oYUnfORC1y/8/YHL2wB3Q/luVdk/GTBIh3
IgRT2tQhWO6I38X+cnKI8FFMQYCmaClWJLA25D10OqfxesogbwOWXDwbcWXAkEs06nA9mNSohzGI
/QYvrIfHCkuiCWvPpupseLesidRJuTwBPMX/MNmgjPdvwaVUmhk0yhg1wk2hnwb0sEdo3AyRP8Bb
LvfQicxpzJ9ghlIIRLQTvsyieIMhbwDUpE7mLhaZxDWpw5pWVRkrX43QfwI+18C0b0VSjsK1NaQt
a0C2I8xLRgqJU1kzXaGiEHrB9283sntFuvRKL0gJDU8IxTU8cyM+oSoKfycjZ0DfHooXLpgGFK/w
5bb9fygIRC12kkFIpX45nHHN1v44HBk+hmVTjRAkRVcoBRMGcegY56JVvddQth7GrpMKZPU2j0y5
zY6HjLnn9WxyZR5onzhfuZAXTM3FO5I/XGcrk79nZBhwv+dxSlMXWlZ/HfW8BnKoNSJysxYvU31D
3417y5UGMKtDw2UFoBUULn5kdUEh8c2Wq4+MxYTcVOKuIyMMeTQy7WfvuUt69qcV3Nwzfig0m6IV
ieC80AOslS7AdHBIDEHRM/o8gvx11CujDsAsA2o+S5/G/RR0Inq/ba9f/WOXfoQUkL0yifsPxSYo
NgPBIuzgNeSubmGkb6l9/Pz0a6j8T9i4Il3EGPOmW7elAYU6lwUG3oP/X9ufZzQoKs7E8p+jAGc4
biLPpLiz3rLyHPKsCs6y++MEYfA/M7TXTS73kzUrOioFQs0Tw2bOkWDkYJk7noYPw62PqBaTD50v
2xICv83xM2F4qIzsGeXxaQ9qsTcyXnqztAh7QLuvgkS79dTPurJY/eQ/+HlCTAs4HPbYWXCXyo3f
tRv7Aub0nnWKcYHMAL1vg/58jUhz2f2U3aMSq9r1iLhluBMMU8/PRZdr0odJa0ErniV3VoGp6tCE
+q3EsN0Db/jp8ASKKHe9mF+9S800xvX3644hm1ZkQtTGbVXnjMvbK+PqunrDQiZpLb4YnJeqvGz+
bdwNcJRKwdZMzWVWDZyPBa4SKKtX6SYZdWyr1WJljorJAGDxvb48KZPjwcuBxBUWoz5k9tQkrQjm
pdEytCk830eRJHsLYDIGFh/REUx/gT0lFkA4jfg93wSwhJChzA7irHl7KSlDpfxNzTlXSgtn0O8X
qkoIy9ZOtSPwi0gZUodlVzGgogfISVV5TZqE4GlE/7peZ3oK3C/ndLveOE4PC02lL3+3/p0aXgDk
vMKKXPAEX2UAb1D0w9FStS2g6pqO3MNIQvMfbY5/R9UKj5FPRccywLqVeVqv/1Heveby9enbyakv
/oB/MihfmwNVl/KcyC0pIeTsgeQCW+POIYorXutpncu41YjlAqubzWGCAkHyoPIBdr4GCSalLud9
RMMHbRHVYnLMA1B97MVf0t/zwQ67ZlSzFRa1I6KK/Ug2DXrdLRlzfsomUoGdYCn8iu3jBwVtn3x2
AOsq/vR1WM9vXhbCYtyeiN59QzKvXjtTD5xIhsTevCMwxfyxU7Aa+yqxgYSCG1klgaxDw9xmPHzY
o2RRNRGWeC9px1f7v/Ud/WpBlSFNqOz4c3bZMIsLo7kjtnA0tJn4A8ok7V12+JmkNjFh7ov6vBuK
40UmKYk/XM5mT/TiUqggsTJA5qEUDxkUSroaF3AOAWJ9r8HB+H77nvYXmV0T6JEoDXbKz48nd06B
lhR20+JRSNcL3OnEFpzv4e26C43dnxqERvrlYhaJobQ8KFA6N15My5SXKrbVCXTAVr07ZBOVGBhz
M6xgPu/qvsJkgf097xq7aC2J1sZPu5xMPIW82J82OfrYc6Mgy9B6Mf2djhKEwRAFhMyoWMrCpA9k
e126SQdlB0rxWeeTwfUo08wZUXcRKBKlgIfFoqI2ErHCQjc+H4oic7kCGHVNIyyIywwyuwcGUM6v
X2mWjppbBHDRABAYBv5jXS4zl4s5uEtfd/d9gQ/93iM0FMl0f2vrqO1sc+w/nJP7flRYYJPBTWI2
KEGPm4kIgcmwGCVdkC57KiNw5sBcCaJOR7Z9SEC/y9H1S4zdnlMc7ddQAjh/zq7y8ZEP4C7kE1so
d7dcGFe1IS1vpipUHW5c/VeVw/QS/Xqq3Io01ll87j3kmhRprbC+a1n4c7KmY7DMUtdKb4Yt9cM/
bLlu77d38mluCzI7lflfpRyFwo17gmhlhymPqnFE7OYs6fbDpd+mY9xskX+0ugpWCbPw7zNUPwOZ
7VP7QQthdovKyLxvcNZAPMTanSmCTNVSK8JS60vRuElWWvtwyLfcxwmsYVV1ScBlom6MrB2+ZFTE
F8gcNnVlgCgOSQp8LB/oDhFS7wVqHFZiTiZpw6BLt8ncni9c72jTicvUBxgw2N4azyhE5zu6DN8j
pDdaIh8EdhKx36V54hKx5a52Vd1xKOP/OoBiiydS3OdOo95YLWWpu/fl7wd6r3itlwKvDMTpWtI+
hCb/jtOdVrdf1FOBsVTfTcvn+sgkZFA1BnWuhGbI8gvCY40v9LzLS874et+52MwzQHBXdfsj8CRh
azrKZhNMHCPZE6i1xhMy936NMnCHIRCICucWEMRztiYd33w6dJyVysIrZbNe829SPWDC/EJftLIE
CiU51d8eQ0CLbxtzxHdwT5g/7d16uRTKvnlmnnxpv2yiBfnLUn3cGTovWsy/uAWwIilH1QJKkc74
wdPWx5L3FSPr85L72L0A4Atym5ZT9lCkA7CGcb6S+xArYefX1wVFkhcPWHW8mvPsiX+eih+ma0xQ
14qtolmx03NDFs6UYMPv+f4+ULuAWkHJUaFWaX+G533J8z8Er9gV7HsC+wKlEhCkgUU8TkosyIKf
brRrij+eBtHr2RFMZ7quZi4PQUFrDG5xKLmUojEdtasyw3aTaRT49ZeD7qjlqGAl6blQwAovM+Fd
PGWDpBTAoclrCKQjphf+ZYc544CsNl0LFTd2jBhIhVrmufjQoqyNC0s1EeXUoyO+a7HfmiB5q7JN
jw7Y96PpTmCQhKhI9TfKyWSE5XKVYBej5wsLv3LhnXa7j70i+2/+lP4XcddFkIK855Jdp9ZTyzm5
xeHn1oha4jcXF0FFzwnCmYlK8KFy/qZo3pIBHTToY+FRXLU1J0+tjxhbCaySDiv5ckB2Y/a85dJX
NWoZ3gfVxbK/neijESl76ULPriQpcGj/h/VPGqX/ZiPJn1egfw03LvT0PF0+K8v3zJQ7NzOPcaEM
UI/Xs6SWq0FpgCMluH/720XwbIMQBfviKu8xGzNmQiiNHKdbz9URJiJLqfG4lLp7JSN8RqbM5pUk
hIe8HWSzf504lSOoo/9vwb4zTo+XGEllgKesMlF3S2OoVc+s2ya8db8M1iqK0PHObD2K0GLXABIg
Ym/u3G/8cKg0kUoPdCMMgu+2MRBNbUqNS0GKbDAM7wt9jmalOH6nwG8OhJqB0fKxyX2gHU4WNvb9
q81IjUA9RB5MEOOhR6/Z79Lx3Ku5B0iS5rnOURqatBpAkJ60VeK+9m+sSrjK/zGW4qP/oLGMWkO4
LPiw+ouTdtbWid2z6/OzdyV/AymF9EOHEyeGF5DD2fYwvx/qEmCZlYMulIG8Dz2oxWTuRLIO+ag6
ePa6lrQxSN0e3LGdX9tW0Ps8zqW/OCmxu9ZMsEh2m0F77XyZgZMruPcsHececcWJ3OwnRS3Gxw0o
M33OozORdbjhmud1T+DNVdrNIcZzEO5qzyYoSKfGe4P2a9iuQ7KML4hmphtKRV24SoPCkq/KYi/H
dLfU76rWl6ddDMAuEQ472QjtBy1c5oxpjm36Dm9g9rAqjdv9m2+Or7a8MP0UJEYqmzCAL41DFbIC
vq4FZyRz98MBZiuoOuzO35THtFBLBJgCXRCTImXJDHOKfl6/bOZdpMq9mZqxY9LqVBH0iopjAYNT
NGYrkYfWudi8oYUeP5CbfIe3SVmOuiwWz+xrJhyY5Pj/qF8stvw0RisWMs+/qtf5uy3khyByMlVc
ItuIooPrHvNlYcyt/urqPnEema5IEQ24y5OPFhxqL/vQosxhwsNZqD8rxk8J+qK3PRuh3Exdjegu
bCsRQlDwaSKrIhFMDD5c5YklpE6V+j8kNqRyVFILuAr5qnMdU4CN15108AYWm+swFrIikm6J0i3J
QEzYXTegnPBby7vfvm6MZd4ZzUNngJyGwMWp8Q/9ufWpHh+n2qJ2kvXTQGu003GmlZXb9dG8xt9F
XGyWku+G5ZO/Ey0bS/FA8F9gwLEBll+2QdgPkNA7hYJEZzBBYugzcxKP2Hp5+C8C3qB6UWPVkquY
d+w2fmauF1FU7seFGPd5oEEkPYgnSqJexxVn040i/bwh0fCX4vdzIRhC9C76FzcOLt6wi75Z2dpC
Rx9ZxMCC5BwvAYCstIbOAMyocHLOeqKuAvkNlHzB5vL7/j6PobBtHnhSiiH8OtigFTeE46rUEA5f
/DRYr97qdj+6hbCKkimezazrsySfeUwte8qMmhnQq7dsOtl5S87qI6Lvo3nU2I3Tk8qYNpL3P092
0WmUB8zB5jwrjaAEtdhp6Zlfar6eaDST3Ph2s1frqzKj6N6sK/K2PSrxvPUFOFsKsc20Z4P9R/mZ
zEouo92BbA1FOS5eLnIzB+N2uFYxzfM1bmE40ltZ2yayOSCKwlPjJcv8pXrl8fptapLa1earPS8u
nd6udndDb1ypi9gQZ8E/HyoSm57Mi9vPUYYf6ygrdkzKJFBh5C6eP6LsikNjJ72b4ULU/jZaNyoq
3DSJqwwMweTd+68dRaO++azSyMGrQhmvjUI+H8ZKUzIocWfSRhdylkNlHngwJuov9wnMOn5dvESY
rfCaUWEb4KyZtxZahmM7lkZbs81hOcjVdk/pgbG5HqyOJQkDgqJnLizeeNm48Mx+zlhviKuSf0uR
xwdBpZWKaJ6zG/4zVim4zJsIDiPA5MEPX6OBlxFWlhDOnyRhmqdb2O8QTYUUsTCiD4aHuYqYbuOo
cVZFFXywnxL7uRs/ra0kp2dzZRaTninPi1rmETpIr+U9bJg4RNLh9XVXZuGcrBS0vTOazLZO3J4d
+UCll1MfxZxSWc7Jo0Y742gmUoCkjLFon4yhQjlTxQBqGnMw1fXVu9Yii4hUak3K/Uw0KY/uwaYT
Y9JnIHhv8Ii6Yhjo2F6gJl2m9svxY+vSEE/ovuCVIGQIQiKH5ihEvyNyIF9ow0309jSPZN9RhaqR
StQjbbKFuQnhlNZzJtQmxtWa8+p27l5ZzVo3jyMMuN7VsNt0heU/ENzO8JPRqVUqZQEmtCxRWFeJ
C+gbptMGKwNmhry1s2nEShsHHUx6h0S3zShk7Fy/sTfcaXkxl2PjtLrzC2diQN3iTcMuNAsOgAJT
qC1vZmbvYlzsWIrYTluEEfGCC4yDXyV8eWoOkHljWSibnzisCMuw53h/OgwskZ3YOGkhmMZVKXKA
oRU4FSoxTVUAra0wVsL1gB4EreAFN5JrAtXgASk+eUaSOSN3dZc88q/KhwnhLE/DeuyhUMfH6RWe
D2551G8NkTKrkC5gHM3Rk6aPENbp7jO29Y80CTTJycq8MrGtofq4K/KRNDXurSLBsb4wC4Qw1nnq
Sm7ueCOUkpUMmWzQKv3xvMYzA3LUJr+EfatntoYN7uDB2lliOxPiSAmHUYY1RrtE0rF+tSFovyHF
y+iCqT0e15fdclg7ylUVlMVeNq2GFXw0+Gn2C98+5c22xs72tHI49SvKlMDu0AQio4QxAV/89m9U
gdCwGFLgbgzRkv/KphT1xLSCGEkTAepqr6ASpPGHUvTIzT6YEYoCHKO9PsayStNoF1CPnzrkWlRZ
ax92AaPgkhzNA3EeAeGCii1vH/EQm7VPrGRapOoj51yXL4PlxaQsdN03mbzxv7tSftESanfcms86
z0sZxsiPEuaTGDwB5fFd4DbSy54kFhH7r1DaJ6ZqY5rtVFj6I6J1g9RUnsMPYl/aPSr+KCzrs/ow
31NH2JhY4OOf2kz/rkJCI/RWYxvwvmHlao4uO21DJnWcE2L2XwuodbgQcOnc7XR6U1m0pi2ZagX7
C5bKKgr5ZAUL3lYkK9UcA7XqeUu3ls63Kmw/yuvKz41pPQAOj909NSFJuPighO6znfLPw1sDz25n
nH2QL/52hz2P8Jn1mdQeLRwGpfFv/B1hdC2S6hNhAREfTtSMgKG5mmVom9IpFd8B1yNiMziLl+UD
/TBj13yXw7zVhx2aGBlNZ6zaaiiol0eg/n5R+RXFrLvDkLhzuhdeQ6FMIkAlnbJ0mCAzn8GL9A4W
qKo87k9Hk1SeIYx7iLFvjczlCifYaufQPZ8e3PzprxsDiS0lY9Vh4/gB4Mx5oyV683yce0vGXhD+
Z19aakp0jPHo5gOL0nW4qE58iwEXq2bIx8GT4EkTTMA7OAnA4ASReurojTszBtWIB7SEpCm4nw9A
vDpsnvMFdR93lMhFnBY5LGq/TEQX4W6GjJKNKHU+/BB9XP4VcuT8qTHWyJ6vvtlTFqK6hWQG88U/
cBeldC8vuVLPSmmK72QT5CLiVGciLlEr7DtFgJ1KXr/Zt/Rw9QNM659ElRLj9yL6lPzZlxxmllRC
nZNHVJgyMGzLf4Ako8nFc8wvumMKZviSOA7V3HkF9aJo4/2to7LPqwIolfe7o2dsh1aC+8I8rRrp
E1GDC+rY0QeXYj7Yegdx5XpNj1ql/2a2Wu9ZkvuXBolx3qKFmiYH8+7ur4x9n3xSkIDK1Du4YrFw
C2yk+0Boq6W2GFfNLeAb5MiricD2VA9S4E821adUIItzUqqshatMVunk1yA54RNOboSTuutnO1Fo
DNClWfTZnZT/uKT4Su6t/obVyEn5fBMAsHyc+J7m7AtnlkrMWSC17n5YUYiAmzGQQAIF8GZzLS+F
MwC4xoYkQxslFZjBZPmpSwm5WQv/DpfygRO0VSiBYYO3FVmTSgS3D6K0GK4qZC0IRU1SuacDaJxO
S0464+nldTuPtvqeQ1DYbbHXBLQwawB1lGFanvblLbY8xkiM6Nev1JDDq62uYg6XrjyAkLl6x/ef
jvT+zNRcW0wEMJ3G0CJLvqPjfDOfPOyG+/8KOYrCaZxVvuyiV8E5oEsPhchuaZxf/1bkM5cBmo/2
+efkuXO8vyYJQBU83mEMumjw7xGGXFCQjsOUknaESaNvTqrV9PbCEvCfqswQAznXxLHHRiqM0fK+
m+59mXDTxSQ4W40n5AKQ5KW1ko9zCnTx41bD+L7OhwXSnnDZ6sW3x+l92aUjtKBkhAC5q3StqBcI
UqOXCMcSTkKIgDLS5FLXkQ1j2adqMVGlDboKjYb4+KFlvg7wWuWRwMyUCDGRJUV26DTXpwXFOwRw
H1tTJXLV9aEvpi6M41fSKvjg8pkXay6IZml6+E8Yx7EPDe7Fv9NSlomA+kkZrcarrhn0bZfQ73Pk
Yw0gxSG0VzLf2AgQtkCdBoIiIlXvvsKPs9wnNfKNNUjwGeeyFbAH99sv5NLeCyZJa+Wwd1SNmU9f
gPRwuJtFeJFM5qEVRFuLEF83+MjFB5SODItCXMphvi2tPZX0H6hV5ZbpyOrU4MC4lzQ7GCiALvZ5
HMheERkkcd3ZnO0VmX9EfWBoRTkeQqx83cuki0rOsl24+nV6HPGKw+Wf+FIzJDWj3ktI0Q5NNfRe
cSJ9LE5yeQflS3mk6yIx0D/kdSKM7ZHzWowavSlyc47t8YWhg2pMAfHf+gth2GCL2PRwc19CsuPc
961XEgHi2dpQeTZiAlQp7dA+4fD7HVQUeoDJakYGrp5A11Lod6mn8kamBb0Y9rkYpt8lnIeSZX5i
8LSzsLVbdUMPXJFEUzUsQ8iqObsT3tepgem6jEv5RGjspmZL3Esgwb4jczXQOr+8SDkEqQvWW3O2
z00FIzhAyAWr0kOwZ22I42DJuW6ZOYG5kzFwRB+Nou+7epEv5IfqhUMsTDtQ0rgsCM9jmlTlVUYC
DWmE/jD3rFo/zyXcTV/rRUMS4sascXDuBQ+eMdRYBRFgfPwcywaGGmaYOTfH1AWtA87TP4PT26EU
ys1Ip5saQCOpAcIDa13C5uY7RCxRxRku/kHiBOpCFun6/KShCUUiLCWs6KDqGcH+qbN9MM9THUCf
ppfcnUa2Xr5nU2ESJmLdHHiZSvYIj0yVLa9QlPSwak7j2QtlLHmSj7cN/nHMpuDnT1J7MdOk89cY
JnizNF2iIL0J5QdCR4qiweB7Kdabd4H0KGYhxsZbqVdD+mtJmyDDVfH7gqyMKsHRezKSEUB3SAyz
UxlfCUELn9OCA0W+EWCqndqvhppx1UHzvzexzp/gLLwhmXb1lX1G7fkpbMh5TvDQB6fv1Q0wc7DY
bOgu9m3WM3Y8ycHZN0XYxPQFNOcmOb4H23OnAyJ+lH4uoxZnZ5EN9962OemMQrNed1vFtq1y5Q8h
O7LxhpeI/zRUhhm7NwBhx2VSOQ9gVnWfQzd1JC+nEnrjQBw9XNXClicaIqPI+SuHt8hhbrlgPeRv
Ij6HDIcw2VYmm7Po5qm/iEmzuf1I3Sjl6ctzNhT4oUj+fjIry+Xq8DL9vZsOXvGvtsZlf8a35MYr
rkINfNT3/6vs8+XobMwzjlrwOyJN1jJtbQDdRN/DG0b5BVikpdj9u225VwePWsA0q2IsAhjXARgL
oTm7EkVtnDQz92jWshTZ2T745nbYKP+28aMCTgdRDkxWgzFmIfXrfW8ZmbFEMferiQSNRZxb7sTt
POX6JsXiarOMeppHyHHZrQarwAR7Pzjomq/fgH3TCNxLLbNpv/KGN9Gz0BxmCtvta7JhycUzP0rJ
VOxBlasvs/ORBmTF+G5uYvXLRoYmFIQ0WyFj2OFCr+3euJqoPszlUTPS/eGqNe3IhZhDsE6Gt3Zb
IOmsV/ekzITlHIKQC5VI8dkVh3n6RQfQ5o68ibj7qPcdzHshnH+w+YS2DF5ms1JIgZCAOAHs4Pf7
eD0vYaEqEsqswa9hBgeOIBnjmJvlZw5hazbhr/s2ab5PZ3Yv0WYJPB3W0P5qsVOhXhVzROWBd4du
LYJgYkacXcdl3i6SzezpBrdhqgfZvm0Ld9+LUOWZKXBHsAlvip0PSkrrwRzBJuNWmrXgg2bienZ2
2KyDKoRdmIvS2Vpsvt0Nhkx4XwoRen+vlodCCsfeSUhh+ODKlsRq+1SQTbAhGIzFH9M2JOipaxrC
sSLKpvSLoWnEz7JnVi3KIrYZWfwHTYKy7ExnM4YZRtcb/sDQ35vzAtPEnCud0N+rRl3KqLhJrkHS
ko0pONwBlQqvU0budNLUQGq0oPDYcrUBRbbTLTHg3iOtlmjgjNzZCpl6yIEP6Ps/lDZqb/BNEuho
vfddf/2U5Av9Aom3GeGghw49kqs8uRKZNnJ0AsbHkNMxmiZCCpO8TRav+nPwcKlM1GWUrXYuNxWW
EujDfogXK0NPUH0bF3Td31ZlqNugf71UPgzaXx7bHBjfDqUeqrirgYPPDjkJr4IE9cnthXk81t4G
U+vPUw1JkEkFUVYNTKDkA+mC4uqW4kC+PPrjJRrljoav5m3+tXBbDUQOMIWPjovHyrmjMfyVz4Xm
qp47uui/Au6DRa0Ck/0wkGAYAtqBf8s3JlfpYZkx6XUdeTMLa0gJTD1l04n918FPALphOrDN8WH+
rJR7/G4GD4qy9EjiAUFRlN6HqWWGxw0N+RlKVs8+k/BzClNXH98UIJK88WJ5T2l/0hlep6pF94aY
z8cf/7WlLhwjoWJ8R7eUrw5tzv5Mf0QeOQ2UvP57ft9J1JaUFRvS/fz7PyvLXu0icv9UUDLhx4Ka
rliDLPrJHiDzlBbnYUh9SIggtmkaC2eJb/wCktRQ9co5kBK/jjb73/XqpwGxAVlvPkNtyyf1q8+E
JLYT+w7NnDjTajGZF4ULxYLLx2wjvFHH2GkVBUOuptPIl3z4p4AzhZ8WtrkJ75X635jv4ah5XpK+
3wAlxxXQ1HVf8A3+M13S8iI0jKL4IqsVIApNR7xHpbfs/iwAXTonu5Ofm/FkdTN45U3gHoWWphMo
2NiQKaiAqqMsNqqwscrIBupeFe5u1ua6v+/AQ78bXfoU6Ca+kLR1uLqdHs0CoPhy0AMTZWDXwW9c
mFOAw2g+69hn4psrYN3+hDlhLU5QAM2JnUCIMSoSQ+TiDNi+i8AOFiCaA1+wLfTg3/UEClmAn+gx
HB/4Bq1YTXqPhDEdUxLRN6mR5luGr3K8QnYURsYJuJ4uTS1oGI4rzPxBs5c31DS9K9CBb4w6rPh5
cnY2iMSq1gNZdPw37dhSV6S6OMLTnLKXYBwYKP8bpN727VFNDLS7me5OsRPctmoiSxZ1uAgMx9FO
LI/umEdkMXEqkQ0bPHX0nbHASvxxmVGh16A8d5SH0mp6f7vODlBLD0oc8x63nxhaFc8Qgbic+Ewo
tFCx0SVcA4euIShMRqkPl4bLfLDZueOsLxglbE0lzcFOhRe6oAufZn2SSTMM5AqWYXu4k1AGrYrK
snMcaV+fKQRsj2VumTHumi5JXqf+LGleqqL7U+SOLERBSugvKUktC4tOr8pcqDJpz1nUDvFH9P9X
fUqSsSFLMgl9C3fZOc5jr2A9O8PJGa8pdFQyXbT/bDGM0suojdJSOxn0+xA0jzSjOuURbaoIRefn
FXacToNfSy+Vbuwp86HQWOPsb5A9coGdWG/LDZf5tUsm4iDQ3PLXMm/gBBhI/eyULnmgEm9TCC0x
LwFp189O9jOKXEIyiiv1AMpkpvFIuTikBGT8/GPP9rkrV+Qj+QNEEh3jm8cmCyc/w92Suxz+twBJ
VNbcpatA/KaQ8FwMXGYux+Qcic43JPOzrvRzfk9RMzGu3oWjVqFRwx2/jSkKeuUOu8yUSVsdbBYI
pHOBSnHqtBJNn/LzY3LQMKCxQ8x4M+UrucK8MmqR24QNSuK61vC4aojJ3tUSpay21/6YX5lgVCep
DHpT3ltrsm+4xPPXJMPZfAUUv3qWJ6RZKR6u3YNaM1awiSECb3WVn9KW9QRK6v1crw9nPIUvwMpl
jXncEZ6XwgzUH1cJO8+6jmo2HrGzpNC3bOU58RYkYwWZ/9mjpIOWzY35QoDaYGgDWFl67LROtiR8
SF/ojbBhm8ltfKPKH3kqiCSkfEk8WST9AvcCbUQzaaTD+FoBYWA5Mq6/qPGUG90BLiB2OQ++8N0X
LtRtmzQ06l0GqFQFYQswPezRNFpiLMvAkFqqfi1F0LrbOOnGfaFGLSg9LKdS+0WBZIr5SzYnZlXM
91en8rJp8Ewe8a4NN9aHZPIoFcyAAakWvwIpvnyYK+uNR3LG1eQGJwpk4oknY14p0WSHhKPVVE7Z
DyFh11jaIMs3HGZ4M4k0sbN3CyG0sS2chdeAVZ9jwAAnn0kK3p1QvaS4G69CJgT29T/J0+skuGft
sdlGCsFkNQt9VckVquVZUIAsG26kVn9JrEppaAdVwokzZvRT9517D/tBsFlW5UIV9q2RU8Rg3psl
zRqlOk5nq3yaeYyTPj2v21OnB6mcRqGZlpB3dHLgINV+qnUDO4nqSGte/5RhYWP/LoXtQtPSaarO
NX8wRzLEXAqWXsC4ZJj0br0WeWzx7gyrPWokcM30kZtopJGpylvv4oeg0SsMfagFQ0cUPB09u6mT
aREEGzl/mo3ljskVRMn2LF+vQeYIG99MkkILW/oSHrYNI42bRi+umYhCP47/OfP0TcfKyWsRt7nS
HpI0u3wQ9B7xFbnUJ8iGr/vAVGKyOyH6DHn1cmxQYa1CU1k418gqkuE7aidPxlwoOSIfnce1Wyv2
SJhiF7Pnhodia1bFq37MsDtEWLLz52vt5hdPOabdMwJiBXzXJNe18z/TKq+mvC68tsf1mOk2hHQV
lC4XGTlZVvdf7HeNPtYROkWLFYUWbiMxCag7ffE5IQXNe/JIB4GWKmYiWxTXIUVMozDOo5hGHx0Z
HSSkjWWpBuskwq7ZEXerhAioHc6vZnT5QgCtAfz0ZqH3PXPBSQvTb2XyRi2aic3PeQH3AhxGCYgs
5p5T2xKCoP16kJuSx6KdZourmmKrXS4m+rDIsAi/6kCldb+5SqdT2gwycEN2nLhJVkqEFmzynYZt
2fOJ7bUaOTEscKrSAdFfr1N92lFUX6KAJDuZ0bF1GRKKwtp8SUFuqBzKL17SBCEfS+gtCsrtmw2Y
tzpWpaIp59xF8RNydAxu5c2ybD5DUwEDh9IhvTRa49TvXwLHVQePkEHngtlU7prAo04D4D2RKvdV
P0CfrKgNfNcw0f+BI/syn7gesqXhJxtT0X5k8w3NFgDseDMBZ2h552iULSLIsukYW0dtOH+nVYBM
NlaeoLI+F8IWpKeIwMIewTcFxYVNHPbHzxiFa9yIvY+rLd595t5jJZtMGnsd53a/AoiFv0SEIbKk
wsw7p5TLaJCdHswhLi0E1u9HlQzdzDa3COrvBzV8yvn9qFJtF7AaFyYpNxr910tV9sprkgwLxfop
hm4Wjt3WVEqf571frwKwKuOuyrfngspJgz6oqWA+Uytn/LlLjlalEHL/Dm7hsqSGkvs6jeih2tBm
Djv2bU6VqnfRNgsEf9HdGoTmovoovcTeju2AhVlEqTytNiTyZE9PUfj06yjkj9oFo7lO7R8DVMuc
2Zgb9qXkeAbs1a+eBRpByhxJNf9rfxa+4EnWj6mpqEslH5bz4x1WJLTPFHPTjlYK4uujeAuHT+8X
rRJD+ylhrjjF7C0bWbcYk171KfnJnFCnC4CUli4kN0MH+OhyvX+hk1R65W4i8v97BtenASoyOFWn
9vslxElLGs+wPeyzdLKUaxoxt4hcGTP0jbt4o6ep6vOZZP6MILT87mtybkrQsil0GIm6yHEnvhaE
hMMxFj9nd0i+T10pQ/pLNo/X87TUkd9Io72Hwk/ClQsuyWtsyssmaRbvyFoZr73Q3o++RPqEYCwi
m7IUyITrs56SFTsVaxJbMgCw3V7xuo9smCV6ipq/mjqM+k+iFWnwPou0SWrRaw8uMGMvnPs8aeb7
e9gx6/zL9P1XeQgls+DbN/qi4k863BYUWC9shPvdohWaw2v+75NHXlV+QlHJjWiJKqCoQriqe8Kd
G/SRE+IgB5u+PAvIP2tZhbk9SyCydwYAW3HpgRRuUsHhK+irr/3EOmrANKP2bFjm4764W7ej6MMG
DY4TnJVi1s6Qtz+ir6Bi+UVXI8Iz+MTJ//TDATmaeSEjFRsk5Kkh2KYboAh/7BWpxxY6hVdelOOl
mU7AyfMQ3mDLLNLSoN9awxagx4U8qNnOwcscP3PrEMxpevMTSn2myiOEs6bKMafbkNUhh6wQl1rj
3OEezCAdpKp/ePDqI8HmBnKuqj6AymYtOzAgwcYrA+pGMOY6jVmur7bRT9xAfgA5ydLA+SiITfTT
J2YlOQzpI01//QBZm0Fio8KOzhVg5IUfVvo0hjg7rkHIiqcdamHdmoW3rMFDuXvO7vTjK5dH6bSa
LPD6YtTjNGNuJ4pSwvNoIwx+Wbe+zRrjrD6FCp5eOb8ju1uWuty5BRQv8gA1mi3eVrd6lBLK1xPW
pq+REx+/WXV8zkvmA2edln+26jRD92xCXnbz6FtazvPBqVaj8WNFrMKLn9WGWXXdXg78s+NbIZBm
E0jBSglDx+JlLWA/ZrjKqr/4LYGmVUAAPrg8sBoXE5EyjAYt1H/rlIecTfQCOOXZMJ6d6NpPVkGl
aGfuBAmPINEaZtM14XlNL/9xn0xZaiHCfWZPz3KWL8RTmV7UfA3VpUwm3LT9bDd6pSJP3Z2PUiSK
BgEWS5o92+0YdXHaJ/BEHJbLLOUjcVOG1KDG9N6To1fHa4a2VCk6gWWtulMaklNYoKZ32i61HmBD
Rqwocskz6OgI9zMxh/BMGm+V9FkGvF12WFw6Z+yfk+U22inSUDGzXuDD+yP/Qc/5n1MfGObxMm6d
DIyslRSvsDUEij6OKKwviwrRUkxEPAzY3cBYU/kFpDtlt+dYSCjaYmadiuE3KBC+cU/cDevEMYfE
n/waC1qdtpKcmocizFIwtdFVTrF8JpS1qJ+lqbGrBRLjsXe9+cvACJgRjk+lOMDhQ4cV7f8fzXHk
3eXn7kcF655z0ViUOTIwkvAXebRHaDtA7oogUDDsWhcDGXYjY/HpaPmlqb8I6dWPpEiJq6nLUOSF
6TPK55GBriXxJpa6bHp+DTPP+EIjyAH3wc5UyLKVZXKHz4hQaXeQc2e2ze5SCN3Usqo07pqCmUgs
CELtAnsfdE5puS/ytc27wWZt5negHwo4X0u08Na5Rgzf3g9Bbj8VNetRjlxWkagHJFV0RZpmPfHh
ocde9JVgyfrrsh9TkcrGzTvQgBHG6OBIVL4BtTSyg19Ci83piTmaZRO/2JhqKwxKwYOiClJk6lUX
wX9sScijGep4A1+LHjQ1y7qXlCrLTNK8pB21M6YHyTTH7ljBunA5D41pNTnbwYpJ/8CG1RpizCuH
/iKjgniPVbTaIM2Y7DKpBRQ5P/+kdyXUpn7x981XVfaKbvAcOFixHkZir2rn9nciXTI0aVTQE8hq
AQH54AfExWxhX5KhGv1/Xypmc1Oixpj/syvaPUhcYOhB3bCdw2G3OBNFlBGrIalP7oATogZVtIiI
nEQjReI+4iUeXBPgQ33dDuA3tTZF2wHO/IoFfNvctoouyspK6UCrZvbrXVxoLLdAZdm7KobAoJNF
aucAU5BC92mnbWTCKza4NLYF1UYihEcGRhPuxGhG4KpzrnFoowSUa0Eg4sa/qVNoXSy9KuXIy+Dz
Yidb2vl2jd+vY+CRWX1I4SIj2G4eR9Jt0tXZaQjVVgkS477ei+Sm5F9Arn+A6bVlRP2vrFi2gl1r
jzwa3pB2aq+fgNn35tBuNB3DRpGwBQ73qEjh1aDTFqtQyWJs+Smf+tTIGAoy0HMHcOaVZukvKDu8
epLTdS2oG5wr50yKGqMfe4N07LXBwk184yHXZqf2MlJeX7HxHuAZNdLOOfaW3KYJDV/63s7/WuXo
MTSLctBaeg42jh9Xz0LoilG3mwz3fkgB19j7bWw/XQZ8OYefAbcW3fo4EUzVuQ2aGcm8LtnYdUXa
kyO/MdX0Q8+nFdrQriKgdb2tUBfddkNggG7EicZ69UDwJdRFFICp2DBfY7xlSgiV7sc135/86Sdq
6+HzT9uRKmT2xWs0qk/6s8OTIWwDYYjQgIT/fH00MzcQmtcCvsliEpCw3qIIwuhT3Nio6cX0kElS
7dNT5UTeP852bxTmI1d7qJoGXnMGwdu3mDh7ys73nwFx686Tzk5Eb5DJwHV7IBpfR/wo1APhOMGz
75kAlrMVdmxM9F88Vujvqg7YDhVvto2wsI13M3erp+rRXcZQUwtyIxcVqP6Pjsu21mCgcGorpH1Q
qfQ4ubmCRp3L8h8a/oEC0iwNHz3pAfrOVdf3lVPaB3oaMHqFjx3//lJtgyBZlpdy6n264JA/LUR9
5Xqi0WVFiQ3U2MvdmSwDZ4h6cemaGB6XBxPJqrH4xSUWZu5oTxLuMA55MSfwZIW5j4wvtyds5Xqh
91b0CVm32cOushPH5WtjRMh8tVoVuha6lTlCSM/72vxLtbyVDXxC0xaChvBla0hK8TRGYA5UG+cd
OKC8I7EsnSIkYCuJnkRVpNo4/Hcav50TBtoL6S+NjQalXNCuKOFapcdSWmcZi2Ww9O1PzrZKoTbe
pwoymD+H3qrdt72+fT5AEKv8L9n/+w4Rqv4GhwnCkKd7q62iuDSghQP1IT05ly42d0KLWMZYTxsG
si0lARyMW03SIGx3qN9hclpG10okyycVXhCz52TQ8iMsWiS7C+ZNCSPGtXaGHUAWMWjyQ9S5268a
XG/DbWsYiKSX6OX68KZ9yD8UoL5nQMtma9Ee988BspjrYSi1mo1og44CPVDnXsZdbaC+i+dHmtSJ
P4tAG71VGNSxYe+q/lFun+2HqPj1+SbtYzFqBMGDC/Uvta7gJ6EblJ127yRkaZIuGJeZfnuyut/E
IN4/B5/TJNHVSoF9XuAMq19SNWZ4aprhOwLjdWMIFzY8Ruv8AGSvq/MPY+5FFkC9ByUhGeOg7efp
oaOsfPffmK+WlLckBjGF5RdempqzUlcryqf5nhfmG7P2QmrmfdfhZfIgjGC2jYipNobZ9hOzD7Xk
b9cIEJyaNPWN2bD7INXtoX6j9eLaQx+10kd10dyma39uoIM+9uq5tEZ9z3/R+E7b1nFAuzKEFJvn
I6xO3zw4DiY/ufgraDOL/s0y++1BvJz16vDpYMAsBbB3VSaXffUMJItsGeECqOn0z1F7DCU5C0nH
/x5t9WvP2eMSkgL/l8FvC69w8Ij6xGY6cxZbeTIkieMlYMeqT0eYpgNt4mCWHXa7oMClCAQ8o91V
6xHV6/c3tkK5vqF/8lHaoxCKlvwdL20uhk852sqzVQr4aSJp183q/GRIyHE4s6FSsHyMIpGJkbBd
KgJAavNjr3930S0cbXpym7MYKPL0/ahYBOTDn2Bf6OtI6f2Nu5HkC1iySxvqeC/OkjfAn6leYfOH
R6P1MJFUHBdqkaidS+XM2QmtSgBCn/i7kjKdqGJKjhqoNmOB0Fvs3K0nO1+t2vDD4M7DbBNAZjbo
c0v9ttyVzqtl+9NMAX68HX1eMFPNDFS6IbAS7Yx0PjUbRa/1Z1lvRrsCewkMxYuzntHiGGfJn+6n
BQIv7d9LhwcUVvPX6yym5NTDVf77STrEJv1SqlVKIIc8AXqRNeI1pdrVv+ugo6qIkLw6SJ8FVAXl
lLVzjsE3OUsB1WuIhcYC3HStndLnehhCDsn1zAV9bYNeyxA0SsYyJgh+X25csWrb08isqI54C28N
OEzg0UBqHwfCf0XS5pQBEL6Zcmeqwqt1obrcpjvE4dz5HWQni3OjkKGm6qa8cJv1ulsImjGhmnq+
FN2zTcLx3xTcU8DiGgRxwOdfdeYem3zXppn7iFamUXFU66UFIza0Zupn1n6vQJOz7iLVp8qYbTXN
BVOcNkTCctcVkk1z53EhMx7JkYZoH2ydZAi1zEcoThsImsn4+75LL0Flr/FK33UOeKVk/8koZMzP
wI8lDGlByW9Bq41rrvv+Q6wdvvcYdypBXiuTONEtHeCEG1Gpo6Tby+NM8WJYdGcO+w3fPkgzJZi4
Qbqlu6/0/SzfjprlCG/plmUJ5qmJM7d74PCaL2lrc+a+xK2IUaKYm4BYDvvpKnyPJYL/hvlRGUt6
6vkchsi6RnTVEsD3pOtN2jPNAS9o50YzGuaBwR227zSqaf1xTj4Gpk4yzWBaMujYIc5iIuPc700U
8akHqay7GaRyLZoKr6QKjeK/k9D59nvTbnGIiK0CyEz7IZREPwEqx7raqjGjrIwCqHjQqwFAnf9X
uRoJ6n5ghEKDYwLUiBpSpLn6ukSwyRfJrzk22qHOn2JyTc36r4PAMvmdaiY0+i026dnYJIXcsJe7
tC6rdOIrdaEERrQvtjaoL/EXg+AgbUAE3At2yhRDh3NmWjqvnnwtEcFDw1Bns8zJHN/4gLZkYbS/
2yr6PVL/Y6UW220vOW9Nd8PpiNFZqgWnoWTxRLfGzqFmfbH4rrWi8j7uu+s1JLzYOH5veWBSHa74
0/E4fy0RX/quzmociYBbdbl1+7MeI07cKz7Hv15EeOY0IQin/BXRsDYr0HZEEJBRM8C5Av8RKVAh
AC3C2vrcR6kxbEkdTiqqbQRoQGq5aRmMdtGypm3HcEaIj26v7J9+em2/7haNVSMwRqUUknXaEKjx
YPSTJMUlp0HcDL0M2b+iHH7hPHrsxXl9cCOTif70b0S+OX1WoILxAH0xRskrHejaVqwH6m8UMIXx
rKhxLo1kkrSMhC5IUznMJnH0Al9L2g5Rv12esnQI577WIXYPKYWcrDFMIKpZNnUDw+lqIl6Ow1a0
CNqIu+hVksJoF0JpLRTqdixASrcn2ozrviO/tt48SyJNi810kcELYwDg+FN+fy2qBCz3ZySs2JNv
T74xWzeFdx3i6MTU+3QnieZ51jYmIv5q/D+wqQdruLvE1Hb5PNZpbbmYl8sfCX1WirKcVNXmM1jL
BawFkZN7Fn6DflWi/06xJvJfpnR8RsMqWNHspuzk81/YGTX9QO6avHGMIDNQYEczovV3+w51pLxC
z1CKPVZsUUPkuOk0/oPeBgG83TllzjvLfnUKz57NVw5Rw7my1w5Yw6hAppJvgoO0h+hubtkKfrET
V0hkXKQljAAzbSVfTEX/v3pVPn6024Aw0+ETygLkOELdaoamVZi8diqgbIZ+aIBgeyIUptp16hbX
rvOdIgpMnAmwwC6DzyEYTpfMCm5+U+avWRbdxmIlqktv7fkcygj5owYt4ZAh8SVVYYdMLllPBFTN
/ixir4DXTxcUitOilvRJYDu868fERlZwnME+cUr1xHvcOBAmPFvAThWgjzvMjO8Kwjqwo/a8GBoG
UqbMw1mtuvR6SYtbPRsUXW3ET01PLzskTMFb+4CU/6acHu8p1NeX5Bzgu+CpWJtiskRtWWtFFskd
uDgYp1pvM2XE6gUJmQTIOWekIs2UsaI62iibxmDK9A3EDh9/rztzliJqDncl1VrtKkNLUuD/JKdN
piFOTR7nKOImD7hydC7KlWoJl45grcIEu8JPdDMqyIE2tZiJeCr9Ro2CNpNygxcM1nooYh3T16/c
QJ5TFA+DmeOOTqbQnpeIrujgZJuU8/WgA+r+r7d6tBhkJLg/ntu5WGwdKjedhslXt5toivz5163o
cfudmQG4Ds7a8Aj4w/KnxGHa2mEzEGG0qMhArnhMmeyZ/nPzxanAAQdi/bvTSl/pLvhrjt3EVtue
W4RS/G24eXFG3iE5mW2rU3//FaXTwWVFuFN6nRnGvsR/etI4PkC2kjj+5w3mceXu8URlWZ96CPlw
4PZX/Y6NUtHuHItXQyfxB4kAFgmUY8qDgsEFdCDex0zSJh2WYm5/9T2PHRC3THDJ+Z0/1JahM/ke
bjWyF4Tu2MTg+BQYx7Zv7WWjCi04XZTSqusBW2Z4KaMlBqeHsznj+2axxSsOzrdfn/YTn9qCuJu+
GO0gXNCMx2WLYCqRr3KzExMcTK8dIQozz7WzHBqHoikEq08jbKGcJGcbqaf0DSog7UWvlniTPAcW
QWqr/bGaTyOBD0YEzV6+uj7b2dO+o9VEMmT5IKJA7sLDJ17aQx5HK5ZfWxDuuM0amNY4IPW1AVP8
b0SmMDkbRs1D9bN97oSIvj5Nc4fTvysmva3QDZWUnMenYHgWb5KpU9xxgRQrImShnrQ2JgsFl1z4
69h7I3ou1M1phbjbyjAjFssQe8EEo1tlveZNZzVmIEKTxQ0K3usHhFm39QyIuzdcsvjbIKmpTWIm
3FZwZMGipSzgFMI2ArVEaJVgCjqOWcep3a90bbGUoebOFZcbc6HLYiab9erBIBsZbHsh6/GQyT1s
0EpCK2UBtVYo3u0uycELTCYr6X9ZYJi8PQV4Qi6B7QWEiup1p93z2uBc3TGmV4Tft8AQseNI8g8Z
5mSPmctmqWhM3KeD7EAV+fTkoeZD42gezu93vp/4y3DbNoyzwyCDygKoKsNSaE32K9FXgnakYaHg
494HReBFAX8iwdyg4xo41x/bd7upihtsxaMPxNi0Lz8RVjeFczghjEI1DbkUOn6hJ2nxRQtKuVnT
WIyAobTqQt3qNbmKjvAmG9zi5CCzVm3ij0UgGnOo70Ukdsml6WV6FFic154HOkPE8cugHJ3N82Yj
vZZT4YxbQeyUEbFWBwWVj0KKyjhKUw5yh3m/epaDtTDHAWsnvpD4MGRG4HMz4LVD3abFPqGR+p2t
UDiV3s5n6y1u1nWJlFZ8ISlWNY4juhwspxhC+Z0yNb5tOxn5UaHbBt683Sjl0IH3j1alT9e25A3U
YF86LLJreeGkHWgpTD1X00qtqKqJnX+XnGB9LhVQ97vnm8lp3pVKf6p4PvJ+6LUMKfe+P6bCalEE
JgZ21tTwbSaXMk5U4Ml+uMbIir50amQ2YeGJ3a8zKLK06StTccx4IjpIx0NgLtYuyEc329GEe8/x
Dcrq9sQo3TuGgYR4juI0pu2nZkyw3lhhcpHcZM9jLIjyOCq292nwXl05UlZZgXwxuUWhCa8nJHLQ
ms+VqX6H3KTpC82eXCUyb6Z68oqti+te9pmHUuQzmLM/NI35NipiKYUDN0fuQSWnL0rr3lXlTG6Z
cUwzj1uHQZXDGxjfjTaCFr178kqmyg+UUj1r8kvVvEwwbEVtlzC5YciomsOZ89/ZNDPf78G9Rc/h
FHMK1qqO4cB+OWM7o1L2jWGhbYpjqAGNnBOqCFXzp2/jjx2j/HQXeYp1dHw7aEVIiJSx8EotlLS6
2ZeRtr4qUP560IMGMjNAv553Nk0Tvzfi3UJh87zUC5dLaV6WEI6d7bBiLitJ7FzAoBqwvWKqc9sQ
haE/UPVHn/fl4ODSxY2lQ4ll8HWCuHrH6sPi4eaY2zm9xFcu6prUOdn1zVLsk3m1HPSckd7jz+7g
oggnN9lbsuIrvg1nouNhJx/i4Fxt1eVYlRE0BZmX4I8EMffYqTHc2NwfJeUWpMftxeSEVier+LNF
GqWGQ4x5z+LLzveA/SAw1/7+5nH1eHQ2hlOLKZ4QOIUrICuYV1eidZhJ/0mnKqpTckHjkd/yGNdn
45l46LuhOZZ2lt9d5kRlL87RxnlQ5Z10dwqtoVWYolgOnwAqT5zfnR4IUvlokg2bUBJsD2ldmMYw
tH64paqZGgySBXm3x3M5XFVOKsaPuOI6M1l4yN1qYwXZw2VTkjLfJr69F6zMvk24TcQDd8G8fTtv
vCF4WF3xuRv+ACmEX6j2TPDoTg/RBx3epCaxisOXTADkgqiKggFWLS9SqMSoXnI2Et8YobeGIXM8
Efdw04wrNQvPW2H7GJbXyJgZJ6OOzJZruzy+DjrIXQXrJ4muNYU41mgT9S/ZCU6Qz8nU68+WY/Fg
MzGzA5gwRKsgrfjFg8JynD7BwtqouzRW5i/eKTynWYbTTSQvS+0vr96lEkNT79u8nlV6M3lAbz/W
UC/vCl4iVshATdlrDMtp9Ds2XZO5zqH7UW4xOa4l/d5AI++GbOXLYB69d/7r+eS6d1TcS+oPQ4lD
S629YiIJKW/Mj/3FYkxzZ8eSEshe0d6as5C7lE8QDvuTiRddxugav3HFZRg7mWP1rX2K7faWp8z6
ZgbL+amkh+7bSn57+R48aeO4aoWs+2+F+5LVKRvKX+DRh1x/oToAvg+ZSxA4SrXUmkdj44fOtu8B
K5YwnnzvbE9uJXPrKxXOVaHwC/RIBKLH20f0R5SlkZxZdO7/ngfU/eOEUh82m+CoQFW5FeuJWOSZ
J+bl2rLg2M1FtEt2lW8c8Zs7V+R2dfX3Jb3z3pg1jemxvhKFjOG8BD1ikCVlu/Y0T/y2M3Vgej0e
VnPe1HnUcZSk/80NFjFo7VkWpGxyCW+thuVSQf/ptD3dbdp3fWq0GGTzx8eKup1GDIFjN7gH4ksS
dVPwpBSrvtFIVWSghtgLT4w1EhdD3mSfymccrOc2OU4K+DT0RFSSO2fSx1AjbddcsmoclGwiLVgG
EtK0ODpZp3w4KTpZDeBiUNJ5gN0FrefEbUDZThNt4WTqz7CthjqK+VMEGu1nLCNple9K4jAOWqQL
n/6ibmpDt7q5qIyn2pzNr1p0EscBioQBvGGIgWWJdM9HHXI/gh9GUyaCPaNY/+cREZxPnkbYWRte
QraK/ttJg716JCL2SW0yg9Xfiqqh3JB2VM0QbBjiz2QniYTYTecH27/Ge9qdWXaqaVuTW1cVJIKn
xfuBooOPryO8+30pDEcri0Ped8JRds1NF2mmIZT2K0/H+t04SoAtOk9tfhQlQeCmF+rkjtMljuGI
0hXIyCzF8KwaShR8Oxbmdrp3WVbNIgVEx+ktLHE5Ca3ypSaXZmpQKxLx+IF5Deiy6ou9+jnFIbl+
o5ja/p6eGLPtHSh1+zPPFh76GmW0NTeMcuQeUf5OrI2CC0a/ij40pQ8U161rwvIgbUiAFz38MTGC
kToE8h4oRjlk1LzyRJ7aGOxINHXqub5IrmCCrEYir7f5yjyJ+bIM6YSAGi2ilR1ph2GssefsnpFH
jwvNo7qE+c+X24aPPi+7iv0paA6XDh4WzICBquknlKG556tjK86TA+5d4QljlO0lOpEnb7xRBKlJ
TjftfeM/dtbEnXhvIX9WERrZPv4OEqHXGVRHtL+GF5AOkivfX+SE/i2JVg6zv1hXEWZBAqvN6jcM
Z3To0tL9zmPpaDsTD5y/UDW0hJebDwmU5DxmkGj/pfmF+T0AHe8xwgWp4b7vW1buy4CAlQj8nORJ
BotGPNvUc0etv1kiZvMVwgVPHGhzHCfbZR0Y2AIuPIVX8+yf4Rzldj5Ksu6eczms+b5du+IQCNdg
mSUUOipyRUE6k0pN6P2ZLMAbDUKbyAVN/rf0Duv0Txyg3ioitoYUgm8494nN+maMCXDCO98EU2YP
Fmp7asqNVoc1xCds1lyPuBxJnEuMcDBgsU9WfqSuci6OhlmNtGC8HunZb3ok9o8njW1VOi2w5nly
3bkp7/s64gVy/nq8Mx07WBjgbD0xdZbyoA37Lpx9tP4i5jlUGb4+fyQPjqQ1eGuT4DwhlNk3IRE3
4EKroY2Mqgu2x0ZOP8iLRsCnQHfwi2q1uOHRQOnG9ryNUQZmO2gw8FXi5V7wZQT2/2I+zkXQpXp2
TXUl8+znMLuS8DAcuYEmJ/QXI04vSudMNaf9Bzw5pianupP3pWZoDQ3a3PY8fBmuI55p7Z1hWnR1
jo3SPsifkFMzZYa7R3R1N5xXqoFeTZPeVv1d6jZacleI1qVCbAsEftYNpdAP5diKZA2u7UDCzflu
gd4qEDM/sIIrf0UDr/XCINf7lWrXFXxhqoOgL1Tmi7V6cywdzmL+ppMa3uaRVqrmNQH43mIpGcmj
6JJFPQvd3DE57Gdhpv3dpbyjk/gBVh5ah5jO3ueprN9HlN4DG9l1Xpwk8BU/OAyiDEaKc04lRaVH
/CM9q62kGpo3vQ3E0sqUXxBeCZ5qGy56J/2XGOnZe5mCjAfPOeBSzJlcVVXJOGtUD0Itsie/LvCN
p/zRZi0YPK8HYXXXVGxwbcIoMthpFHHe3IXDbkhzFRyYsz9Cewp8Alzz4/BKfju9osnpefi+QVie
uqbcWPgbjdUTf7pXrD8/uIS9n82CjMYoKGei2NW53WG3iZDZok14TmYCC40W8CcWE2HIc+bBYYxL
cQU/A0VKAqBJb+1rTc/QcxX1/oI5Fjz+X/V9NU8kyullDyOYShjbNT5QdNsKaveUMvJgkNXJQP9k
b0Xt/dtvgX8GGxxjaQ0fgEFn4U1tcBKGo/DnRBnbNpdu9bqVrzQ0AyAI6rvTkKkZV+UZyWmHyUZq
cQ+uZfBnte9H8xJeUqcZL98CEqQbmGtrXpEzyncKTtq4BFU4/yZ8gAbb08KD+2k5IIvIGEsVXB6n
cH48RkxTfdMqG6uuougMST1vZVx0vGaE/aWO84OpuSc7WkxGTSTOrsSjKjerYyAqFh7cFfTReAqz
J399JYEzZ9xQ2ZrgzNQJZX4rgMzhfKpvl9FfNz1xad1PN6dZhl+J8svCUbSfZ4cMcs/dqtH4rK93
OKsR/EAYcHyImRCk1Y+ff8/e5lbbB9qSFqx6Ir+nDZu6iwL3mU9jjpNt3D7mxOMRMaYSIcW2E0uc
MtC04XXuH5ZSklkG9pQUrxNRxRV44e2SRIi9lQ/dQJe8JHoEgqOPbA2SwYU2gFutBU6LGTF85AqV
c+KIl5QL8BNBfFN8ZfmlF2Bivrt1Jb0hPoyfD1qhBLP8E7Wwhq/xmolVkK3Jwe1fT1Z4kJioKNzH
afyX8oB0HdprbppDPGIznEm2jU7nGezKa0w095AXqaeexl1SCn5OyKs6poomA92ul3UWGECCrWFo
FPMnju9RIk6caqwznnTGeuH58EBetcNCPR92kcXCchdAK51ALg1SOlUxjK3ES9zukv6EO6y8BkOQ
0v3G18T7qlTrXtL/KCKZgu3x3ZkXoDO5oDpPHzYENmCSiCsHk6uWiRJ1oYu1qv7MOPNxSkjNPAQ1
3vJ+UbfmCnt2pDUTIgsbjHI+y7jMfIUC9MeKRPXFeoHCs80l7V8B2hZSDnC3VOoPKHwMqTSqZBC8
7UeTtqlbKPQs6EBzl8nLECwwxHyRQoGvKkcnfW9cT5aSJgDIs6g6JM8lw+ENEPj4Y54Tqa2sg1mQ
AriKN0BQlaQ4ClKKEsnvq7ZbaHXimBlDKt/5WbaWHYLyjBGOKpQsnBrlL0UoMLnlkdGWTOnj5K1A
ysihnG+Y6fniMrc8bCf6HwniuR4lOM2CIDIaqyd1hTi3DJH70TCIB2sESjWs1JcCTP0RuqsL65dc
Q5KXadpHy/+2pKXT2s1vpQmfhqAypS4fHMq/bESodnut6l8c886Dt68v5RMGtFad5EBBvyrHjzKB
Zh+CEV5+KG1nJTpa7mxeJCdq4QxaVCIFmA4oq263nU0YgcWshA/0JUWl8nJQBdfmVdlgnw8chjWq
9ooMblC7+h/pBWoGeQeAwt8BfHpbm0zIyeJcksUATso7YKcis+2ESFW41wd5xpKpeTATVfmddAW/
N8PIrQIoZL9819WabQZkvLnsl8R0Tt+0M/cAQylb4GU82Q65i8vbYRRX/EoiQE0WjwW00R0boodL
Y1SLzEj8fD3aYT9dT/yaGLj2WTWS5MnHe3VIulfq8my81IIqkHhSfrcTVT6qXrVS3cOzBdvWvNuf
Kx0Th4CQj5EaK0nD5bxcufoeEqC6kdEYfmzHbr8lmlXG8k5yaIPG4gxOh3eXm8N3n3LlBJSZjvtU
o51YvXQPptpwQHs9/iUNNdrdqVgvwfZwEx3ZqUF614o7hbUVWyEpCdpD7Ib2sKItpajHqIZLxwGT
L5ZsZYrFqAibwU1NHXHrTYd3j1O5gbVsd+/M5u8jfcWdD6s3osHhDHD8pTHjfVv3I2kg143caRWl
9AxGAyEGeJcaP6oOLMeWQEQ0FAkdKuJLjElU6rYBSHuAGYFoBzv38A4eDaAgC7uyZNmzaEJeoVHa
mZ2RTt1G1NpK0NRNFGLef5GCZl53QG2GBEnO9K4DrTw9+NSVbmX9nhschDebyiWrLZw/pXjEZ6Wi
LVSb+r/Nk4+oAqeTg4e/LyC6TFRI26yEOX0pDGkl6g828Ap7H5i9uQCUmDX4daEm941C5r/+y77X
8BrBU8OqscLciIF37E1aQkrUcpZ2xdtJrkCKadtQKk08bfdvYDK2mQjQWWRpU9rz8uN3RZ8PoW7f
OXVIVXcoZK/nZ1M/Te7FIDYmqRjOjROl7fCD3tYjE47V681ejwe9Z/TH9NdYERtmZAfQ2gzpZl76
p/TbyDx6YGmjfeJOPVOjJ455JgRl+3KiqqpA7/HCfhVMM11QgcoaesE0vCnLaC/vlvT7WRPXYvw0
q71GrE1G79yt6y8ow+Q5lTiOnN8DtP8jZDHv5hI9qT6GpIc2jUhuUV2IA4XgpUkI/SjkT4nRe/Sp
cvs/zrvCrqhP3GgzBBPxfN0xlsfYJsf0XOWOEvO2J1KtNmOm7/+BPNLCukD8wwKtiAS6Lae8Vspu
TmwyqU+0XSifEiTL8lh+8Vitzt9qmS7DMfWn8LOcQ4UQe/mNQa60D0GB0zliw0v0XEKEKW9CWXVp
4LtUlf/lt5GiyO52Pu8P3+jEyrRz4qX7ofOizvsyCeZlf0h9Dbm9qpL2uYBax81UuKO60b4C3MvD
NNfuNr38AGT9oAusPLIQrtJUcfLEU03Oksja3zSdO3ImKbni1YBuZcNSNwSe8/Be3ATOwtyJCO6P
7tDdFuvzZcF+caIESiw+QGk15/CHtg6WjrgJA7jChAnDQAiB8MAJlkboprlFdMLyZQakmgAW7z/G
LO4tjQ1faY3DEUYpbREOB0+A4R6HkTOxx/TUwCmLxlGTGgzUDnzlq2P+LFzXTGREEUWZ72P8na+Z
wZD8oCw+QiV/K6K8BB3MkI2LgNfJmHwyK3uww6vj23kS5btDEkxcOBszrplIhSgNYTtwEn3tdvdB
P3zP5dj7ZdKF5k0HFrqZyzgoIJ6UOfcOI4EJqoiqvJTXVPLAq3idFJsoUGR4oopp2pmvsSIfPQes
ur3sLuL6NUYOd8cC7tkMg767yUgnkRTRZRzTHkurfSwpsSCSqjnIqwRwTADmCtGzZy/xaw208xTo
gkhmvQ6I+3TkKJgQry6XZvoLNHd5gdBuwDfzBr/K2G9PKCQnXKef2C9Sp0D+oKZuKvmPtPDL5l7r
oten5LfvAP0+v5nRXvvbHOLqRDVrhrtV3j43cxrfAJEcvQRPuXpUZT2NXEt761+L7y+atA7jeUxB
UaFLL+wfPY9r0eh+H/hqs/EPLVse6bK2RoHEMCzJX/8Q0kUKhBPYIqhNsOJ4njRgzkyIe3bw3PoO
ZgpsxTtmYSVdR2OmouWsjXSywD7Rtkt7csmSmWo3DfzJRsNW8wApP3BqVRfxaqTnNz2mDSfxaDWn
I+v9vOdruTNjxwFen5bZaF3MJIKXcaAnBn+I0KF487iEOTRHaz8ptvIR9MSH7LHQK3OKWfcYWmqx
3X5jLIfpoHMYAnEH9JPC9kQLLsAt9QmUTKKhfjOMwlvEJQT5/iBNlmSvfh+dsrSE6CvOGuhi2SWq
hfYd3mT+AImcTIJnmxc99vpET9jCjPGDpneADngiSwWw+qIr0MpRysL3bu+2U0vBoevdfA6gMXHn
b9XGyLaEcnfonqX21m8rIwi5ddgZH9hpZR8E8g8FJu7tt0wORdEzzvSyhFfSA3UfGSiXdcuKiwWi
CEkmYvPqRk0D8DvdvHYe+E/kQRNLHwTXHq4znMkUsjhgKedOJYGcfqgMTcqrzfht45H6urwCqi86
oamCJws95xbU/xHWwA42dblOkcgXflVCoTouskNA0WUWL6UwIxZzkW7TZvJIPJYJlCbCYYmFfVe7
IzLDwr/nZlsxFV5TFbeBfF/2Ol48PsJWXdOX5FbQqXUsdVuATSj8R7rKXOmVR8WalazlFtNUu866
Mwo7pjNQGAvzNheEeBeqg0PLOEyM6EffyWrfXYkVVysrqw7X6WuXAywTc6Z7UU4IQc7Ai3ExxOxf
y3M0gJWR9PZRAPfeDSLuv4sWrSAmqnZYVUO31YKKJNiFPVLnmBjGXgsZqfWKAWUwbClRUSOmUt72
8aWwKsxmCXDYVaksraH2BjrazfbRRB/3iSpw+ZfFsP9s+aCG8x1x5S24QsnYR2XtzF42DT+ry5bK
b1xI3wnC2CkDlk/k7kO2cYXUa8gfJtilYgvClkl4q7wWdsMW4sjsyXlnqnibgTkqGgR+TSiXssr1
+BdAVWq3EXfL7ittn4tiMvlsUwsrsPf/gW78PK8fOA9Rv9NnmWgS03Mgetekhkf+S7Vy2SBmWGAT
J2s9EwNzaG2A4DnzAieNbHr2aers7GTS83wFyIwZCSKqLwN8rElTBXH7+MnM9JlgvEs19StczYms
ymvTrYcXMMSL4iy2/JghYlTv3B0nxQS7pQaALm6aB6/YbwJhFhcY5Ew01SDq5oUy+KA5nFWRCPMd
4pskLo/g/GHUT+zt10jsh4NUpC4p7NgPB4oue63tHUccDFS0TSjvqm5JB20APRgLfEBPas8jKzBi
QMaY6meV6LD92hnq0o/6rzXBIv9Yj2Y/+D53OW3v/qoDi8e7tFup/HAizNv7+1jNqSgRHoIgNnSV
BuD0HJxtg97lgZPgIMWyoHCYSWYRRAk71I4ydw/rTRQCA6GqoY7txC5d6CWyVyeFYpsxxrVpBVPO
D7ZlWOQ8/zjUy81/KWd4AlwrBLcloKLprWRQTYr9qwuI04LlPW4wwlFJgZOxEjJ3PL1mB+AsHAJZ
6Of2kqJjD/tUVw8St6pg2OWDsVrkIapwUMS29bWGxz25U0PGlWQOKFu3LgkFBj7UQJ/p4z2qblxY
5EWfEk4g9H+k2wDpvO1XqGfwd6HSIYdsZ92HomAmVpIUGTdnNhdT2AOa5CPkyBrqX0na0QKELYf6
u1TNxYDX8IMlqgYdGv0MkcinUhRnxBla9SxkSRMrG8QCL0/9Q0IUbwLddzioMlk/XWBaoApWqCTp
0y3Nyzk7cQ1RCTIELYiuCssv80G9n0VwmBeqPqgYhYgSFIZPD1cmGQG6ImBO1kpAetXEF6CDa99U
Bvnr9absm4z7C5eb/HiiZQsdVYW2X2/Hlwr3zieaHooGBx8nL6aa1eFXjd133ahaHDUrpSe68krf
T8YJta68lwilhYQEhP1MfFedVpb9lpRd+jKfNpR8bk5X/wbesRYm+V7pLHHT02aHG7U/qJi+I4MZ
RYiQm5S86PzUo9A6iKW7PWIklyL+Y7bv8RDLcdXVSNguYgiGmRLZhh6t2T6ZmPgJHttLLGSJ6Mbv
THZNR7hxuKvJS0Y/qnsSPPVjzcfpLnMcbPT6GLPywvAfZB2n1a/yrwjs25prEQoJqnGpo/0rtUpW
DILlKW7V4oITouUuuSVBI8SUhwwYv78UcqZuiJgfALxIOY0ti8kOvXWmfuIYNzl0ged8YC1Zk/wa
PoxkQULkFnjJ72h/bdncnZuoK+SDSmlwwrHMlSJ0/NrNY4bKMAHbemiezDHvyTzC5y2lh/n8KGYH
sVQfW3uo6k3tAMeAhc2TBEeFNyAXRfBiisoqPg9mKQGhjG6RPsNGHWmsfcdmNtPjXOXkJDZK+vrx
1p+OZazpDF6JYPrxs3cB4F6g1WjKwkhLhqHApnj4zEl4FfgSVzOslB26UnFjwSJqq6OIDXPoqOZ0
kmplYWndEgVmT3jbwIW4uQYwbS75LNh3WJfiMJH80XccN82kp4gRv1AVrxzmLCMnqNcs1VyA9oaU
YL/6SiLnCgsczH2gOFrKSACtSJaADDU3Z9+y7brFVaZKPnzo5eFTlWgNEYPvZSgE92fnF6eZW3C1
LfJdvEmt2uNuj9LUQFa8b1XYcp7NBCzJDHwDbLN/Fl12RpOPclS6MTdJVzw3cBiwkn/ilnv9qZGE
6IXuWHvR6qqxaEmaOy+YeyDC+UmLvgneTpUubt3WQQL6j8DGYITK3/jIy/5MDe9dER9VprVwOGVs
qz4hg4xKrfxoVn2zQbLQNkYdGkKfN5N/BGpoUJf0Bfm/KnDCq06NG52iyJX0BXOkvwGTVWknN+af
i4PbweuD82nxJP9ETspgZ+PVG0i+qzdmHnsoiLINhXHqQ2QSNCjB9oKWAt6YjcIlXkkK70G77Lbf
je3lGYpGwcZo84qgoIgq7omNc7y3L71y0+O6n7RINFa2OxCXKIYxECmSRilLurHK9jtcwGdMfKE7
qvfy1ngob3bhv3ui7daVsPTIn/pY294kOnP3oHLe2Z+wVgpAsJgBUDRIDJyt9RO/YrzNzyWHnN6T
moEs4j6S2qf0uQ2OcIKxi68+quK9i/I0AtCL7QaVwDAqY4zAqbdY+ON977DNon+rpfCg7YLfwd70
Z1Yn6K7r8DglxOlhL3/sBX1HFmC7QrO/vwcnLycisORSJIlM1/lCak34TEDto+y7nWr/4p2qm0lt
dRRDtHGnZlLAa8++ZYkukX7ymRvmK1vRHx7UnrZz1c/xWZZMzF0j+unNo03z98f9qmd4nmJODDs2
xTQGcYCV+a3tlVw6IbipvtzhAOTlcJ+y7C/hqW1jbcM1/0l65hvfOg1IQj+lqfjbJS2RwRS3eVS2
/BUoo1YVB7k3U9OO1VN+Pp8gDQRl11CgK56Rzkfwi2bIGsA5E2NeXJek8ebSPGGCl6KtHG7lWaeQ
dQ1Ow5lsf+IBXGy0l7boEUB3JewYzSpg0xmSxYVgG50tUJzejGhLWVt6B6jGvKE3KgAYnTTbi19l
RP03bPHS+2ykFkrnEa2C3f/mODobuZhEfsZ33iEUdHeoX1puwxbIdX338JE26eCk8T67NtVuUnTL
4f8cC/OYwVqw5E5Rznx4l/rNaF1OwyASubeX8mjNXx2UmuAfmY22gwZfP6B3Xvzag0zxLaeW5RPQ
PyY0/IltI2AGGJotNJe0uTxg5Aw5FFJ5puvGh5Dv9jssbRUZWnV6IWI3U3VSjs1t7IlU2HEM7/v3
4gH8C+xUkEMjhegAAZAJ7U1SxF5DsrnM+hzrUIXiHirTi7KTn9+vAOq3a0A4hDxb2Y0gt7EPWa4n
14fQVby7fGwPawWAelxhXFMfEt9M9C05dVSfnQoXw1YHDU+YYThPInFWXgbFJD2aS9q2qGtzIEFE
gXdNd/7l3NUeDPZjtnv5uS5z210dZtq4XroFxysbY8VBbKtl3bp2TG4IfIcgQrqtkwXbYHobqmCo
F2+cueTLCpFqbRQABsNShdOfVy/hekaesxLJ5qYVPuYUbVxL+bosXbkBfzgXmv/xAq1spWzmeniH
Uo/2Ar1cYcAQRrpPsLrsUxfs+wGbl0Dk8MZgxIf0s8lHtRwwCNTA1JXgv8AQKbv0oOW+nfNLsok9
N7n6bb+1UB2ntw5/yuzVojDYwVAwXP7qLrmDLrDWjznZTfq6unhscO7x/oZetAq/SlApx6C3Fzeu
AZfw5N3cvEM0x6fP4Qo0yn9dB5myb19HxlAOMLDnxRxl29MDhTSL3MZzFl486Xoom4Mr1vH/4Bif
DXu7UQTjr9UTSmBH5Y2xa56OzKJbaL5TKkghNYPb8BhggmAFES+LNxChhtsgOcW82VUEX0cmHM0h
EjBr+d5rWPr8n4541pGjMTPwAIz1wB+QGVe4RGjexZBH4tSNdpgsKlStKJE6s1chQBMTG2kkRzy0
9AygiK7kNQ2SMbggMltl7au1SDBQYHA/S7H8014yAWk6VffsAIUxJQIjMIdmrVB63egP3HGymS5M
vmdq+xiH8VPBE8DnSx5yVv1OWn3EJ2Goy4+89mpeQeiZtdQaV+toul4EG9wl7PUnn3xiEo6HW6iG
VRqgPbeYcBWzmUSr4L1pF3uMTEq5Bz49nzpKKxJxLyzJrPIp9Vugh3yEd9+NJF6Fqc4pvmyFeeKU
7ordPj00yU67vNi659xInXx2EQoe1OL5WoIY5DnL+iUTf7yfHWWQQy3ILB9sGvigxwGOA6SZw1y+
aea2GOzqrPx5SGNDpV5H3zcedkk8ytesVywStvgyS3V95c7GRpYWXpm+tHF7qiV/xF0EanlbhEGI
Sq9QoXsuy4uoNZ3PcgeMR6zXudfvdvzzQVKMJSnG7Mp2fAzW8+PsAogtViYfZwlYJKEpZmnVk4s7
yDj13uPWFfb9xnuEv7mKQ5ySC3PyzeiqiNTFPb5pOBLWPE1lJBQ3Hb1egxvvP3C+VVgjOymjUkhN
HxrABZ1EZHUuWtiYszrlQzYe/8uL+jonV+Nn7F2vN898gxNN52lgKV9yf8OkiG3XwNEIHy5kwWZg
2MaaE7eFf1+3ZZc7+IjPEfuyrJXAUmM0xjcN7+78ATVNTCmst8jGCD1n5WHQaQHYVwJO0/aHZ/rs
v0pQRG9AJ2fwNisprtjhBgLT1J3mLpJ4rjwQerOuLwGO9JlDnZLKp1F1fIpsx7TARg7/2LIQHIeg
kGdrK6epzSriWgwPeN4UQvs8Ru8pj4+Is77aFqaNLZObr8QtnNq/ldOcVMaBErWOknyqCUT6LKnj
bdFn2WUQjrhaNvcG6a/hoNkX/1JM4RYuSyFkqRxf4aqC7r1XZ78hJYTJ57EAG8o/Ukp5dxin6tN0
3WWO68O/dBfTz8p9Z280/1WT3HSaUli8DDdfTZPBS8r4K2zLbfTvUeOTtWBr4DBDk10yjNN+ul71
5WmZSAdo32obasHVNIYJF+agZsLsYlExJ9X6BO80g/ULSxbRLKLNdBpLIDXkUIpH4PlzOlkSfEqb
shtcOCvJWYq8BvB2VppSLWUxWm6fBYcp3OB9kPBlJFuTqRlATSeo+kLbPDxuY+av2ge0SDv1pV6v
oay1se7H7q7BYZSpPiKP4ygZFAAcwBAFdKBSw44BiiJ4PyrZnOMRzpCEPCse3gnn6oMFbq/tmshJ
mFUhx4uK1wueyfrvwvPGA4NcNd7dHGTNrp1yZ7fZ+4GooO1bh6/ZLq8RRIKMYnuBn55H8aGx8B/N
o6ui0a8RN3laurEkaRnS8v1OJtsGxh6i2Osv2fHQomIBYf4OsMQDFfFVXBZtFJPS/wXtn0JFTVV4
8jBUa5GCxKKiWemfPdRayVr814wmcrHFDEV9NEv2eOmSIFI2UalFB/4rtgmXIRCB4YABoEgPoenl
04bFvkWXj6ecpPbSLeQizG63IQtV2SPO0kPjSCy4TlrTSJ2grLdIH+hgHALoBxAiXgPnoVkjw4Gm
VJwyekdPy49LU/wZP/4NC1wEfaUbjFT0PkPMpVbxTVRF6GfovNp+BM+rLICWCF1MuaRUCWbl2eEH
i/cPJnuUCK07Cu/7XMffoQtaE3nAY7Yplj1nY8rEO9kJNTzQdjY13OtpRezoTdy8Epmo8l1Cy0ZS
Mp/e+GqeXM0TiwYBi2gtqbU4dM6ed+WTHbDAX1tOQdYtPQRIqMA/FwXzS47WAlIZtyRb24dBiiHz
2XBsoO7rwb+qaZCI0CzZNCTIQ7vzBRgtQqI0kb8k46UPJYr4eog1kNJ6wlqCO/8lX4YWz1Dby1NF
tEmQGpn2V1wla5hoqczRYwJ241u6wrEQ/BTnhaCbHV7gGoj3fJeoOwCUnDh17deoGP9Mr1Zu1i8X
wbZCpBmEt9/xX3y3DQHYa630YcmG++M+w2D7QFAWmEF+FecmoJ5tgqGnEmu3qcr16tHvVTiycm26
bDv2HUiI/+pcyHNiuwR+jWcK0dA3ZmwqA1JSC51pII0AYgOMfTHRIIM0tl9nDsON9p5sFlJNqmRn
4Q/99rm300p3eAINuRChuwWpZ/5e37Qmp9afP87NNfgwZBmm+4rNRFm8SIbYFKf3p1RRu77/Khi/
Tu7Ob4K5sPM1wYqmzkq+z7OZvIAaKg2FQoexjFYqabU7Zjb+Is4plGFjgahujOnpcV+jRfjg3MdD
rkeq5TEnribnXZYqg3R13hRYNDx7RDhMUDdCGu2LsztuhNzNOw2g+/vGoNtyeDePRpRhJ7FH6ab/
F4WwQpx2w98xNReRI5e0mQhCdQ/Yk6LNPdxer2TJY0cNaCw//FswdnL6mDmT9aRRZxdHBe4bKcON
fWgBbLnvk7FjC6kT7xgtAPG2d+NFvrfUf4zO3WymMxGhd48EHSzLMI7KGSmFu0b6JzIJLOP5wcjX
t4tKq4/Q5hVPtLf+RVmxZ9E6KdSKjdA1t/+TiauubQegoBghc9A1rv6yoo63tkoZvlR2wFmw7voA
yKo7NLJjAzJoXcy7chl0EC86b/dj1+iOwTHJPgw2nElbPaxPOHMbe4egphNQGZoDfR1HGnqvAtoz
3ZWluHmRyr9A3J91N8wbCuq/KRJ7/i5MALXHc6HyHLEIr/iT8EyKI16zcD7acsTvaT0WhcFOnmwC
xbhHd2wgNjrra9UkKWHhIPqmtZwhd6+fk+PkTNy8F/g5rpHhngiB3R+1g14jMgHcBwLW1EetLs5f
nqiHRDxilnTEG6JZuH0ebj44h4Qx788Z+zGMHF2ERTkSClv5/TXzkzShxyadT2lt5TAmRLqglQ/I
scgCf0Dq27rujTXyXTtEo7cEPLRTvolZ+7CwvtsdHpA65GHz6JBgeWC0AwfrvQ8kHfKTH37URDo9
O6hKqTVu3i7mTRDn1lQEE+EU/jGf5fZz/b0+HVPANaIrTfijh+HY6iqv8EEQ/sHujB8JjkDxmlF5
H9qNBZF86G/apB/py0j2KNEeZvg7y8ZY5DKAJim97+3wIrRBnpM18VjaF4E+76+HYvd56yOYioyh
tfT9I4MdhAV5idV37FRUWnNas+e/tfL8uORm22KYI31QjxTAdKJ95IZ7E0i45NAxQJctOifw1n04
E5KHveHge6TjOGYAjWnFeXsIKe28LB3WnOBy84kitVbn9j5wy01uxAVTwOzExcFHAkVtzv2fU2E1
YV+52Ojf1cTiOdasZDyrJ628ngzkGCaDZLhiPGjvEKB89zKHs2qnkomHvIqzy0E5618DFp3Nonus
dbVDdHUHDfGXz0h2rH5NV9/HSW1q6wEfE6uWKUitZMB2071zzvfRoELe8aDc2T/3Nz49bQu8+ltF
3xmRfZQOdcAV9CYuPtfCfadRim53X8lX8TEWqZh/xdkLmxGqw+KGWoyFI+hoGJNPI/E/MgtEk8IY
zM86j7f3y+qu2Li2hzeTn1bR+rBBCkko7vvRX5Oai8OVX/nAEQKVQikRkVeSejsFAaO5u4AQuPB7
E+H8lulwglNQuZPYz2mHw6qQJ83wiiUrNo+MoL3PV967ACu3AlWHLQt7nljbHJdxSAg1AMTHfmH9
dSoKD70yX5ZbE0Lv34uTkBvn6jj7q+oXqS0qybVocVR+S4+Jnn20yUWraybMhzViNBVU/ZRCNBAK
efeIuOVW29t+YTqtLVE8mkufAOBVpm0UwCnD8PZCgh66G9ZAb1sp/+en4YMHe03JrSoXXIGWQCNh
1xW1VEONgUMS9KiyZLwsLCORuAQhJmocoI5FvgoGcG6QuZH8uQEkL/EuT82y/hffbcJQ8TzpcHn1
KieaiwyV7JckjQWUGMP1DHvyxSvP1nRq3AV53YIBsHZCLRQctSRPra/zQX3kg1z374KCrkiOkMcr
ZyiuatfdRrYj5DjwNReWMWcaRIdxDdelT0PyC02/jovDfurUxbm0wnmfNIMF3zP05rodJGB3cHkR
f+RCJpC+TQbFJpeYYIYYN1rUfwsPzdE+tZ/+u/fzB/na+UlL5iON164tHUfCSh8SHgTEr3QoxHEL
iMQ/LXjMZ/ltDA7mmhr0BOFoWmz2j6lThQmM9NvvwxJ+Rfl/gTHtDaea5KobS3cHdsdj4lrvOniA
nKftX3iFgVeRTvrsTWt6sheuM36SA5az/golhiCDTHwf1OtED6eQRKyLKW/YHRv5/1cHbUoQSOb9
cqSAmDQQ8Kiz/b0AH/qROVTpAb/aX/cIEUvyxdvXVedHF1CkhHq0/v4FR36mpr2okl5U9XlFqh3v
3gNDuQHDyq/yu4ZhA6DDvn/GeC0qjg+I1DI/qMUL22ydsc5D4SzGQNswUnr9YBGIDDvjC2Ve0RPD
G0qJbH/bpcHVdwd5ERQKR5cv+KUinEaCNtBUGk3p9xI5gBmh2hscUVowEwAJOdLYhQigssRM7vcB
zGWFUm1NWsGnToo7bkUAJuxU9sswiNhYhgSq3Lz3V1pTKv00ei91cj5wLesornyI9KRwPcltXGtl
/LVtFcGnS3o3eDhvHNohE7RS5OIt68P7EwxPJDfk+yqlClmrvP4GjkHYDNnnu5U+aM5nZeL1Q72z
s9JosRzaP4iH8L5pN07qmdxUmmcHi1zk4g74WgB9c4xr7yEON1wTe3xwWGkAyM1pp9xg+Ruxt2/p
Fzm04CD0nDYT6TTtpgcHTBFzGjt0JkYq+vuwHLuYgq/7hrdVfhN0f6MymedYA0VMES2Sdy24yfzR
ipjOQGPjZ6UxLoZnZl4cgUWOnZ1UGYpkNdIRTdkB1gYS9/s5/LVAqZUNO4z5kL/hD99jDNabNJn/
ifYHg21zUOjsmq5CJveUIcSEyqJzBf831J2l3+iREfKoJ7iwTWuJj9gI7Ah1I5xHiIylg2ryzTqp
fTAgzpsWd30AL6X8aEFII8MjCG+mvwQ8yM+yYzmKO78awYLe87ZZNj6FfhuzZtemGUcGGClK5Hbq
Qy/hivpgFzF4wWlFSU6/358p6WxxZRNZxG95yn6uyROdTada9jGctf1ZcRoXNN++gaWviArPdZm6
PO7l/vclW/Am0wZ+hJ8X9ML1YM23uLAbCnfYyfpX+ZLvAKkrMBWiABEpUtJmIv/1iNLU2w7QAceR
RnCToxaPE1kweeglmIu3dZbHS9xAaFu0zF1tflln7pSi7QVk0AKlOWmn/pl0WIogculQ/k3zFwqz
DzrVG/+UloAG2Q2RHSb0lTsddBn/GYbzRBGmzw/kVDpCi713ABAiu2fcZUN1Reg5C8bbaWYelE8z
ZCOMoywU0fzK+j3ympo51qQkPG3SJhlcMrJPg9tK6lq9r9tMElrdUpv/elUflYmR74bATkM7IiTE
uPs5L+pSKCHAUsrdaycUof/ss4QI6+o3Pnshqm23I36vv2hp08DilLnmdzDjM4PENEacoldX05W6
Ow0cqT9R/AcimAsjl2SRdqBSKJavlmShUkD0AUdCf0EGvw6C80Vf0/q12qIqSXN1DsJp9Q4YcfLw
F2fDhp8Ci8+iYdH6kCvpP4g96xhCw9IVZMBY7Px5v0tBkQH7+ozCcsyOG0AxX6vFxg7ILd004rpl
DagLL+VlqqQkK0WIxtQAjPtpPMRzNkxC5nSlKc0TcC6rYuCLg6KKO2KBtFo5MacfdZxyXbHdRr5m
MaN3FEfGMsqtXw3Q0SlY/pxU7aeZOPDAioVqtJH0FSgytWL/+2QL0Ovv6waS/K6yxvOil9w34aUW
dnXYsQQk7gF/1y2hiohDRh6SXvommsCBRsP4VoO/q9p7H8OngHI0EqviGGxEEKYD+yOqPHfromTP
1kH5j5JWpUurRit3RbhDncGy9uUbi95247R+bvnCwhvmMCGVsFDBYoCdvj5efdkN7ZzZw6VVE3Jo
w3dC5EbvIgMeSi7FTDwrSarlcMeRVrSfKmGXoT7mYu1pCl35u8Cl21FrCq22zs9EdPG7XsBp9Nfy
YuAJNvjA0jx8ZMhloWRywM3eE+Pgk0Q8Exuu67jx/YZwaRnacNFEHXR8EylbdnyDa3hb8UX1PRGf
U8ahCjFLBGqSMcEzWiGkks5sc4ZFLUOh/3KOUYXJ4FVMuY1vzHYeG4FtzL3BO7hjO0S6cqKA1q/Q
8d96ddi7sCCoka1YwLmrcAn81nvlyUh5j2qVV079eVgiLCjAbAhO4CKPW3JTh4A78BK7MGCgGwrz
P2N9cNf28xfURlVoBYHCP9Cgcub3cC81WXv1dNOciULXkKeRo/2n22FifjCxLPpZKsIsUfvOoVGu
eg6GMGF+pLECrBB5bkMS5MZZPqHLyYU1NP4dfE+EH5yJ7O89nCKSfwidIVFCfftWX4q9pWAb/yRC
eupEy0ROmljWY7IT8z7eIvOBqdh8qJwJXgDP1HTJyIfUWvnYkB30N9on2ppdxiaeXIs3jUS2TJQ/
bA5VJE+VOgWJOOJxdColAqLVFZHeF7izGqKNWMpSUFJ6I6YFqiokeVY+x75jUCzST9nvNenMcOKp
/YeKKGfnVZSGdmDf+zby9w39DaS03Z8P48WSyYXyeAFLKaSCc1aPV/WMFS3YYvJYYJrBIwQuGMUW
ZMhia7oyo3rUTMvJbvJWCBmM/rqj7OS5gOBM9Leg+xeUtvhqQ6tzWudcs8ageTNS1czfz7njEPdo
osVMWtJjhRp4KsRq8SRTaB3PxhKU3lASfu/ZfjJT28+MR2mK3RIa2RO2cJOm9rZ48XPvkmenYtwF
KByBMl80q+ApFlPUP7BufObbBSK6QiveoHLMgRCZri/z/Tj/7Esiwawuyg+IzynrlHcMX6K/Mucv
4/oJP9AA17p6qcwQPdiAFNS68G/+Fq/PCl0JjoIqrOgq2Il0gi3doKlHbASkCWdiQRKLrPOclYKJ
iLHyS04GWb4I++xQPFx3WopN4I0L5Ew1F+o56B53yRnqyDbqVMPk8xzrZqVqhha4NZBELLmUKkFt
uObzUOllXgRgLvRl9Fw+wVsRCuDFEOqVPvZoBR2KR6JoCFFh6XezHWWhYva/H2KesZI14lEhoVvY
t/CO9qP9RTW3bkyZGwyiqSgFAb62IAdd92RXOa3/j9IhKThSNmA8sD4esWpHXckjbvyV0TI2QAJ2
D8AL6wW+2/HQFKSjPCZUGttqDXEWfsXaOVo2+LFCkWgYRpoN4Zgb1VbFF80yiBlLStZJPkITUiRp
Yb86SdbMLN9n8jZvGo/fYYBVX4j1B83hSjC1ceB0QEfHh0j2l9SUZDZ3sYMHYOP6+fhppVlRiQFD
cfl6TY/A1dn+KWDE9C6GJqg3Qsxl1Bniy6sY6HZxNVIM+3hLqgdSa9d9JXAMvwtU+//wa7huIuFE
imuT2Yj6EcQHpd9ekrXJYHsA4lQydjV9sPWn4C3W42U3TlaJye4efQxR1wiOm8+zGei75XUM09tB
YI8ew5V+7PnujU/f/UmJURtRtQOfXXoIKGpwCxE2iOq327Px8nVD4yZiVkjmpLfDsqrMqkEgWZ+E
Uj3NLgSbSnsIzJs86LtADsxGVZakniwsl3Z1tFlh9/vlS7CtZwCDINhBxICZ1gkq7RFtkA9BAd8K
zumJSIdVi7TwYzF5a7e1BtnKjnNIbBYpRvYa/i5VG0q3wdzhjwFrWjiVdTHrplSGns2e4F70Axzn
kf6w6/rSepMsqEWdoxvHG+MImYFDpbKYRx/xeeWz2WWjam5+RfkFdoFw9kFuK9uZ+AGXrHNHjP8c
eZLShxGJrRBfan+NaMb1NTtjdLLCHrzomDCsEBgsevGOcUOr14RijJnwO/zCRjGEra8FS0R10vVv
1r9aV1fw/eHIi2XclqiZvVbFO9Q0IY1kQmIpINpHGejF5YQYws72ARykHpLBrG8LrZ63FSMROlRy
BSVZfNl/cM1o+s/4RrAdEPwuA0Ppv/AgkVHvwYPn3fjc4p4PreSjN0Qa8uVvRkAOdQQTKzuuRBQ8
RONZ8wcaAGkPYNuRDX7H0uoH2HTbj954ZC66cm8+JLopnpIB15Dj/+czeeGMh8TusjoiLFmmTVNY
1LMVB/SldVf5GsenI1F6OidUmqZJ15mJu92hc6k5lUEFGlhldKFLY0uUegF9I8M53v74/8RCBnxD
RLi1nuv0Ac9rAYUoMjgB7/KhpCAjU3cukVUv6RnBYG6O29NFb5qwalVPxvKTD+gnk9160EQq5foa
W4l4PyndUhy4O8FqCch/4MmijsXGpz711nvHF1hFCaMJoMDGfcg2kAo7dJ1IJ02HyAtAj16eAV9m
LK5I7/Ppxwpgmmy0SmtJzSOCGHtZaiYENdU9JWhuOEOSEDijrP1jRwcR904BARrO7SZrRdSXMWk1
5WOxsEmvp1XcwPTLJ/UHYLX29J8eN7wZVuLYEiYvkE44kd0X2i2t3wxB/suhgaueAdcshXv9msrf
5MExQHNuEbsmnyn9D38pDsEhybjuoZ4yy8S4w6oL8rR5CtGG/hTn9ajRR1/X9wvoxzVWSxCk/Pe+
vaz2v8G4D8BVl/+mKIWcyIKZmKsd9XPJ78iZQxtx6j2/0ti2FRNFDvkeAN0qcOgbMydIPETJ+qdk
lyqtI5Mz0wSgvezMxwlyrMUWlu0FUNxbkpcYkqRxsmBn/thjAOEEJQ9QZyYniliQptgbDtU4fHit
6nfCqpzTVV3E9P2rUyKL1XDWnrxsYNhLGZ0u2x5XxWZvyPBKEp3heY95NiaQfE2i1TwfXearWc0U
WJ8DdCm69ZIjHnuyFAWTWfJw81HVAjRZwq0DhtmeEHwzH6YDonZvgTwkgabhFVQH/xCjKmnHAwoq
PUg3HoqoZdz4aMxku2PtixFbSfgTETRKdIlCho0RUUe4L1TfjzYkMmuSw9yRkw7O7a7vKU6bWbig
XZor5N8yH/TjGl5H8zlYxbRLR3X2tGFRVyT2uJtz3x0VB3ASjoAyh7WW8yQnU6TiudhZ+DsgSGPQ
nPYCkUKenjkRaMTeHKuQAQdt7zkRW5jPEnJ8bCD97IOV+yjSJIjKvFqAFTwcCpMODvcs7HRwiQtv
W3VCVQyI8jpUBKQpgNpiozmlhAuW/w4zvt7IBoMxeSb7OZYyRGxmKoEA1ck7L/T55OQRQDzslKO9
E+l1vlU0yJgjGCUDJmCrpuz6ii6ibBHaMElVDLOxV3IFiraEkIj3Ut8GDk5TFvFTIDZ0zKKnYoj4
vUCRV2svK43qdfEi/kLHJaKBOvlGtRPQK65qy/pwU4vA28En1tds6RhpD1kxIZe6dmEEtDjJ2w8b
5YrPyr8OXfb8IQf+2xbeRpS/b2CdVqYdEclbOl5vC3WEdf1HCXxyoc2uaen+4FzJv+rBLqdTV+jy
UpRVbH0XGtT0tv0ZbZg/CpCh/iRrFdQjhEWV95XqOcY5Mk3utMFMN4TIVQnQ1EoklO9MHRFJzrVQ
fZaBnQzAGQxbpxlxJM2HdgE2JG7MFOjmUH8fAD7IN4XCkaKEqDfgatSbrMIML8yextf9mIGtKVjv
o4goY8OubKRjnHksGklT60xP5l0pcC0FOKwUNDulviGDGInRaB8gy3haNHhf3+vqj95u6ecxxq8C
vQRNGxQtgGoki5YUIAl2RkqsQZ/t6DqHkvum3YY377f+J50JEClqLfJGdZGH+WsigM21YFlExJw0
iFSS40758KZlLc+q+QfndnUyNRuqlkZoLnDo5wKOCK3IjBTGNv/CwRNzKICCsB9aRTWi+esrQPpl
gd3OtD/XZNDMMDNOteF6udALfgSFz2PnYcdwrIZIhy20pi0oAtPhyOw5hcgxlfA/QbxJhItN748Z
El8qWsqvb2fjthlY61bYbq0YPwRv6CmCTITKzlb4DZhcyiC967v45dYhlcklElSaqH+gGsBbV23O
ANhuSH2/HKJdSM0x0TGcvD8n42ERqrjCS3w+pVkZAlVP2d8lRnd1gDXVCUv1EOJJsVCAT8reLFgt
z6YOLj0/JzJaiCy0KZL6K+Mjz7rzs99/l54hwg8aPJE+F+rL4IwabqxspWlb+6u5aqNJUYSD10I9
iUvJb5qf6dCLLRFk9Ovg34/C5ANNNkc74KtdiMUl9DcnLKYB9gY0jf4Lo9w4A6W5Uh5V6NUhi35a
gpS7tl6v+N50bH9MhhgiHLNU5TFQspPg6s/VAaVL+/3MYQKqnFA9KduMd7veQgX2aGVX6UwZ0SA8
hod9QYSzDxmsKCQV9UiQtyOK/EbNpZ38lQHZrxwxaQ9LSza6WkKcPJenlZlSlPDhHy9ZreAavPX/
IkWn4b4mf8f3awyFBWwdBGQKXStwU7zi7ajMGiIz4cRPe/K6UsgnxspI2eR/A+DAHMYjvD8aqrLm
MxfiEy/Wdk2A8zpBpiRQkF3JpG8meavLCrhttr3aTwsori3lMoP8SaYW0VFFk92fDRn3he8HZ11o
3WLT0jR8QoobtivbLt8HbJWga8ZUIjKmSujDJjpIqztLLyq2Jn6tG96l/ESrQaTIVEoJBmJ8sBdo
+6fMIDxFB+EfD8vw/h0kEWzqpElPmMVYLz3imX5eICzdCfS0h0FCWAenlYK3C8Vcicl5aoIPUuv5
1r+RJHOcUPk4KvgPXNpa8O5QiYVJ0CKA7u/JafvodIHfgKJF3K3l7dRtGZiq1Fjwhh17fQGy8IHX
YSdNMstoGG6p0z6whMuAFKCKijZA4YKBADgO8z3+gSDE+lNrllu/KZq59/z8v7q65AVB8Q0sroAj
K+gDGgSOjBSzax+2oSCsC2UloqbI7wILd8DykQElKj93ZOGXLmgI+vzxD/BPPI+6jlZL30aZ29vb
1TS0RTWZjB9qD09lSY2t3HtzOX/a/GTTWa8leUn3iiO3tAEOpyJrAeWTNMstC1pDnIHJjnGVgtHb
VC8Hh3KIAn94W0E5ouUO3JVE4A8VmfXXml027tuxkDdGPygJwrClrNh6E3lb3OKlCAW87ObO/GnF
QwmmDQlUkYRKQhTevih2DO/FRDcWeTiX8xXN/CoAGeyOP3YM7Q2xoB2xlhZueCHRp/EYU9ZMkalN
RjzPsfmhpnHO175JaxK3PRD67SQhecxRadcNK28L7z67Hwe3vBIMByfa/wIljtiCgt2XbwExNboA
SqIjK6oGaXalBQogTs3C2qhdy2pQtlk2Dw8j65MgaZcVrMaaG7sK15rURxM3VLwqbskZGb+ovWuT
ecsfIwqw3XkGmysrbqnFCpWfMJvdvIo/0JMR2r5590nxMMVuzBgmGzbK6VTB3cvk95MQzqf8Ybnc
F9MaHU66icm2T2pkTd5Ut8gJT3M8zmKQWGgO7ENgHgq5i0+O6w2bjJrjgzrQzI3FGNMyJdDoUBFx
nApADCTSjE66fZ61cUrOwdFPJPRnjegbQGWyBeuhchsBp8Vrn2cLjf+3mB5izXwHI3SSyVamk7EV
7Jd9z51cz6AG7NvV907+rUPH35oldKG+CfrTps1dKET4N8ABnQV4EKoboHFD7wIM/9bY/enIMqSx
0Lk3pZ8+vjCkflcTqWws3GbirwewftnKy7CuHRhURb0qsd1LutpJDerRwbIOGF6DuMBHMMUXzfuN
PqBPzHZ5FstFkniYHC4W/QkL2zbWTu55kIBZAwAD1UwI2tGPmhsNGDYqJC+/kIUrhyoC+FVhpku9
pf3f8s8WiTnF8Z3NH3gXJlHc1wlv+bfdawbM/0ZWwiaeK5MNLviIhIut89YenI/2UdayKJvmZG2Z
egaONptrV7ENlzqWGeihKRDnpk5X0OBK+iAaarcdLEq743U7z4vjQAyXC9LyXtvOhJkF5oDQw1Rq
2+YxPR+aDOK1XtaJ1QFfjYD9/45/bZH06notPjUX7BPUsc2AnyB0ZVtLWbub5KQYOmfNyTKA9vky
zuav9Tgqkeiyms6uoQW0VRuPRNL4oCr3AKqPdtL9dZyEybw6wStvAmpBt15Fxlu3G7TJwsya0A5X
M5QFy/QSgq+kVLQ0mkACxSg1xZIcYLizsDGNCc/nY6UKuPFqOH2eCPsr/spUjeCKYW8v+TKgj5hZ
APvPSyYkSnkWAiunIK+ulKLVA+2duIwNv819oohpSIPJWDPZXYos+ZCPX81W+7cqnQP7WU8u/Yrc
sHODtdaRBPTMqAsQK6E+fKcblW0ojhXXaIiPvJ/5mr0P+SA8bFrbywtarVkd2WLBTWGBVcvbtZka
Q+rePHaCAEgUua7IrauMcstJ2JcbiNUe7XAwYBfEeAAd4hXxxoKLT4vaXtVitWoY1PhilI6eKBYB
dcHo8KG7di7odibx3Te4Bk3NMogFzAc1/AHg76eYc8Qo/ixRKEVqOWIqiNu/b9VL3MSvfstiTfWb
GJCaOIT4rBuZoaT9CmMhtnmJYGQXMoDYunmxetVfNkQvmO6hgc5abDFlRYVBvBfTxU3jVrzYAzoZ
9tWg5vxdU5d8T+MEn9iaB93zmq6Lk75DluMgf9eQBXLEDN/8dh6ua+6G2TFQo+NXZlWZjbI1vzHM
YAfgixLpqSSxcFK9fod4E4/50bFfcIsR+/Z0Lft1ANzpkBLcvaMvwdgx0fhRj6yfpkOGc+pa3DbF
EmT10Sjx39eyzqPpXo04vy7q5cf0HGsR2ha0Gz9ooFb8KkPwuRU/Xp4cZJ7RWe5Lkam8SbaZJFeW
xNdMRFZPVuxJLy+iFGLkGph27jkqXNv4meEr4I9gClg9v5Fg41VGmsoNpHrYGsr42ZfZuYdwWMr9
mQDwKS6PwyljXJuSMkw6sxMVXq40pJHT2J1UMqb4rQQbQ6o81xHAgPlZfL7zsvyMXVCLtWNwaBtn
uL0LSBz2FRAZdz6PBpsH18nqFesJYQGta+azkt40UKIGd4UZ1E6sEzawah9iXapL/t+UoeWDRT9p
Gd2ILY1te5yVM4xmyEPeH8AVdGTegVuOlGvVx2WxYG6+DyOi3JmiZ5LujTk2diM5tGdl19vAZjFe
I9k7EqEHLpM6CcbZ4PBSMTEuTE8L6QAORoYrPiIE6smSde63pq2Sc1cPCKhgEkQkm/KTinWokztd
PCzUYgqlT+SgV5DqCbIFYJLIzwgKKuBzbaEIsFw06GXLUdLJP1jjfeW/t67SWVYqeHs95QVqQgnB
9YByHZ9LR0bM9fKKq8yPEc8d8zIsbbjEjgZJToC7sa/4Obhp5Xo2Tu4KcG9E+8RMXa6/GyjaSK+q
GBIkAK33daENMQ5l8ZwWZTZNZkpDFoH1+LvfGiDiUIHpZSTvIXS5XU0zjsGR1GwIPyU1i/swRw3o
94LKU/Udq5ZmZHbBDCThBk6yIZ0vJgL8JdXjb/MAW31zc5jJespC0GpcnNTd0EovWp9Bq0HMA42B
wdEKPOdmowPmVIB48yvSho9LE16uv5ZdToehal7OFqA4YoiUDJwwW+RLrs33ssbtdmDS/NOSnPdV
o+RB5BErZ/ClZasOAh7tfll6VcHtUJqUwpD89lV5LKSDqGNe1YefIMEJnsFRAtbVU6B8bZf/Z8zD
dOQJhtRkQDx14zacZ489MUe80Tnnd1ql0O2btNhFoSYRpLrZXatLCBqUJR3x+W8S9lcGNBSCtgsM
PZviqEpPBryT/BkL+8D62P7zawAcjJUC+fV+sNjupCKnGqox69Ck0WjAWjTimcBGrDREU4q1a5Ff
Nb2mlBzY1qXsh2vwOOe1xTeLLb6mrv1ST9aXpbbuSA8+ktaSGCEz6oW6MuwBDbRaAR1+fHT8wX0x
RAtNMvzHC9eYoE2E8WbPaj8v1opGxC5zlrmGLpNSBVTq9VCBKWH2GiaELJTj7Z/eK0tF0MYW3aKc
Z2uVRwK8ZnXeJhQz52Q6ihqm5jWeV6B7YZsi4ieKy9O8vks2o1oMzLlXYwoC3YXkDNGOKNOe9PvV
7cTIPAAq47ibNaZ0NL6LNWfh8asxGocM08K6UZyh7k5u2I8RyTDC4tB3OGaPBAjgwjWwHRMiz/Ud
TQVq36J/+63DW8NYYaCRug/KCI8b5yCVGvc0Lr8tx1cmuv4bnAbiu7r7++4TsvMN6lJzKFW/5Oeq
hIq1HzToontN2wIU8WeIk7QcX017rvcfsIwgP9ltF4NmuUS8NOUMcKDkD1YOQNj0hNj5Rwdk103m
Ch/TfxPP4ONQr+yofkfgPdV8vPJMLGvLxti1Qjn34eFZh2Qr2+Ikt4My1bMrpd2Tgg1ouz4PpuHH
8ykpOP47dT4mpCqwKuPvvjlLkjVVqN9OQKnRdg+wGwIZWwYO2vFmoYsGsP24GOnfKYsrkUzyn2Fg
gXBaxXVuLBa1j77+gIuOT/fgYClUNZ91tpMFmQ/u/Xmj42/XtBHi2glr0HL/6rX0Bx84nVCkV6L3
e3YFw/in+AjVi+dO0gETyGhl0dxKIyv3FDtVNzPYE0skr+l8Kc//9PhNanw/SAG9zoItVy7ZWGQv
+PyCunQzCxYjtnm/aIHCCa27q4L3T2QWcrE580W4nmjXYwAu48cHgYeNmPWloktpAGuMaw0XxHme
NuUYeUPNv5OPrPItcnUMysGNxjY7SWW/ZVwzJ/BMXvKhLkxhQI7jXj6gHWPDNnn34i5N3fVEnoFC
FwCr06A/pw4bXlrkcPs19SIVXKWkE4zb50a2XscweTi7BPzO8g5ZB57WR3o674aDwNQ3dTxCbUdt
clMmgYRDCikK+WCeh/HWD2l7zT4UKhzIyTxHSNy74ysCL1bJhvDUUUYGOC8nSbqLlR8DkQJev+ur
Xp8EXFDwK+n4/iUlG6AwuK62VuNti0LVn/8nIxwYfU1zK6NtIy5AH4jxjSFOMkO27ed1j0GFRwZ4
Stf8P+ygCwYuVhM4wo34yYfTrGQxfuIAgeMtCO8oYMzKUJP2FxxBzb1l2phgeZHAe8pVmHnCFKP9
JvnqPsMNGxsayAk+X5QewMVnyeiAFukVHZFQiqsk5g+eeP2C0mj/E7wDKc8T/8aFYxg+jXD/aF9W
y/QvRxGBn5MfAuclB1QZFp2xp4aMOppchHLB4TE8ih+AUtgxYshdW5uGNE6X7jzBdpTe9xF5l28z
JDkKFE6lFgSPFE9MxA+MZfCUxRUSEGzVuwOvygzqeCr50l0LH5/ZfmljytTKjvTMkVKBGKn44sU6
5LehnGhHRSsZD5JwhIKDPA7a0fXQjAsH9bXPRA/EnyEenlmYwy8bT96d+No0JjuZhVMcTz+pcNN+
pezdoCVdaxxRYQ/rA1LKAWEaKraFcY2kkq9uzI3okFtHi4TshL4Npg4Ne+FUZqgqW3lnfeAoxvIz
72in7fIk+IGNLU69B0jsyzfbMf9OZAW7YnYgvav+sapBYWQVl6PVU9qwAAJK07VmTAopjgu1HdJh
hqKt7Oeg8npTlRCOxCBwUGd2bUW+PIUB30ppPU6fBoGhHcbCQvprx41/66VGAGq+1x1aNy3Jxkbl
y61wlWBj8d7Tpvrc1BEOX72+HVkGSr4C/Cumi8qBGfKE9uja2rglvthkGtEh5AjO/ntzjJcQfnCH
2JeKrs71q9qQ5rqScxGEgjrjNNvspHx25yd5sP9n1vRUXoeb5XJJPHKOiBslXYGS00pft9RJGC3U
DTr2/mOFHF90ESjxIaSwZkdEjhIK4Jk0IYIro7KC0BQvw+RtsIbSYG0eDQwDpKJc2mFz+LrnU0Xw
zWfkCkiqCoZgeqjhgi8TGvWfJdfyiP2KNLUs0DElrh52+RmhQ0dydJ5CmQCQoKjmA0JlrCSXpfTy
vv8nUbyPP7ySfVBsIYqDlUuN8QBvzlIpm2TREZ3m8yFUpMZGIvBSfmIavQ0I6FCYiN3ZT8TfUGiN
CR9urYe21IlzxHPxmTOT5W2nN+fq1wZiaaPiYFMbIhJvPGVlKuRGmohtssPjkzMTUCbwLIVfQzLR
fHXEvRxOG+08RyBZ8rmK3EfvnhEwYQxuZRlg68SfskohiajynxKuWENkzkm0nG2NE8VrsZN/VwbG
oxCQqf0WxT+dB5fUdEe+a3ISReyvriKY9gJ+GxboYvShpBvNcl7kyj50Hxx7Aw2eVmwzCs8V0suk
8hoGhqLErlmMJB0q6qBGoSO7yDZr2EA0LDMng04w0VTjrdhORFMIdh9bygLy2XLJDm4/AkNm4Bqn
gEY0MHTOjxlV5TzySHbT/KwNRh9EctsuuqgCBbMLe66ZpRLLuYqaw9dVsr2TsRUzAlCMkNtyr4+J
6KCWZhEm9kewaj6FOqHRkfSO8uP6bpnkTSQNnoJ92FZA/GH7MVTcRGfVlUgmu+Q36O1mYAClrgyf
ZPrU4B5/Jiz3R0kYzuVHHxaN15YFFbHzxN7ZfAFhR8fXBdzn7mO2d2f6RIr50htakWE/4DOURVMy
46+WUlf0HYoO3jOtOON5WNm6aAaG82Ur2gRse+asownwaJGaF5KhwA0OuBsIIblp3Oo9zYXbAPVJ
cbWyDj1BgAeDuPc5jG0qmTppmZX3U7uKZrWpm0xSpjgNFYMzXYxiOil/SCydd9kPVXvhLFRti4/i
LCqnBUKlBgPd5Ixv1L9wTBKLCju4S3lDGdEkeBxGLvohMuqN5fonktGZ2/9G7CjTmLXcsEhTMIm2
Vjcmby8FOks4cFTmJLUUqhbu5lvS+0eMQUDx4rA0wkYvbrGWDHplGWsKETuOwKn52uaPywAvSodO
EtL4O+I1Uyp7nFQ29PUCX1GLRnRTPxvbT+3plw3B1OvZBswsk7Zi5+uVkV0jkICmjHKlOsXK6Awv
qsxSDxeaFe/Ly8wSg+eXfHEhvg3UTyNsmznDUr7Bx08ox/8uzpGYAvWGYSploKty5/5ofGX2SxDp
Mj5OBys3/rAL/oxvEleI9TM3uifzVSUA0nnfeXO5Er0w4VZVxSeIC8OMdsU+e1nmtdQX0j7i1SCf
e55tA2GqEdrGWB9W47ICvsQrfuJZkStiGXgJcDoD38KYwS43XbUHpD/nO/vXm2sT9ZU85Y5msfij
s6Nxh63c49pSrgBVjQ1wVuOukrtgSIoQQR7d7WjWKSmG5x7iXpyOHBDsLuc6anZCXOe/AAY510Mz
4qvG4NbOKqMS68lRrjRd9fXds3omtBaRbxnotBcgHt38Rtl/jsZ2H2b/HMj1Ilmq2f14J4cI1N1Q
0ADjAVfxFV5zek2FQWNo0Z2dzEQFihcoZ4Johj5AVGA9RSFGp+Uqg2xo2LUi6K5WiVXS3wdQt8kv
1AqoTshspIkjjwwa4HPHL8bnWG+2gbWZTVJ7zBr3Q7tBBd694vZBW0/jzDjwo0HpSZWkGsUcDDGa
VYA/yg8y8ogdp/JlcNPoTRw2FqUAnBeli5Bmq101ztlxxb0+PxwNXHZqN9nJUDZHpdsKGnEgUCac
Z4hT3ZJwMMCmSozlCCbwtL/WqqMixpHomx94yX1gFeYvBQzPSVGrX70fC3cbMHjS24k6qh/vJJ9a
y2+R4iEGZ7Q+aLz48X8kVX3epxx8Rsjg9GqqIvFkm9xPbuzPXq1X/IXmp9ERzj69bzzn+lmpJtbP
seBOfihqB7YHqd9yFqttqhUKEy+Tde0/VMJr/qAicz+B31jDnVPYcsbGDax3YQyB163LQ67F+mJl
kHYmz211B1utWnhrkhdlHR9Z6hcnjnHyhHbVFYm41R/2tq+1ulic4Yxetr1CRwiYo/l0J8MvF69b
LpJDNbPpFAOeVAha5WVv2A+h2k2ItMkEOA7pkHOL7pPH/EUji8iz1SvUpvwq53HqdsYFryWW3l70
POTcFYsr0CbUlj5E4CR6nk5mKsKeSV8vArOQRExH2ADF6qGuPbvNwUk0fueNKK8uo4WNhOZQ928a
z8LFq6hi5PWpjW2agTgfnzDdd4HQmnD4Y4T+9LU++wn6tf9US7fvkI9Sjp2o5Rjp9Irk81jGIY8o
i26nQmeb61EeoXR+4dG1iW/bDaQ5SlLezg7Kn6WkEYpZMyXtoDl9v/jjP5lRYjsjIdHUXknj4lwj
gY+03UzpgvIyctbXAs71fLNG9sPFgqOjf51V4BnNQ8CYt+DlBmIZ1cG+j23+SFdnbAjjHdxAsmts
+U8gpnG7KEb8qwQ0pEnWgmOYn0S54XXwdF3NjtEGi9o499x107CS6bccZd8Q+Mt7nSGJsXQrUVKs
u2K6UJwXktGOq4kJxnK/g4jxj06xfcYyEeseUPCTMlORzK90EHx0/bvNtZbqvbADGjzyoy3YuanJ
McQsuzfWC0ycLd9QJScth5tr7yd6+OdqyTGuiUleW6Mw8zbrDe9eg4olcXFyfqaaWPdsNwF2JKXP
Yqd49B8za0s/i1LBAILdOgRG72YemYQOUEAThtBNHI/wyNqBs+eL4xTLNLxJ7saVNzKYO6I9iUN1
z1h95x0jkG/pzCl6DbOaSAp7HVwaWpHR7NBvc+dVU3lhlL9vrDhP8wkOJOIXGSRR8GFcQZuGWaKf
mpGz/L4FOpDkt0S8vVLMd6JMzJwpRUdODY62NqcrC7NZSmYblN0T7wdqiQdznpyuRkOmg7pmkOVx
zSEJFxr+Hmxdq+mZcQapXyXUVV2bff3HfTAD3HnFynQvcXR0yYFdxbfCMJK6w6ffH9A6ZJXkvVFY
PiRfw+xWcboF7yA6gOwiwGhM+Aynb9UBjWwBdQXwR1OA8Fudps1uIU7pys8YWT4DzMG13dRExN8R
FiFAamA0RQowvd+aFxGus34YIXnQfP6aW4zRSY6w6K2S6dz+LIquuvKiPpq1ke8L5WCFQ7/2tjqj
ik7vQzc6zPOkfv2iNhnT5wLbYj1AJBhnsda5LqMmtBwYEOmiUrLhHNmWZf1k+7L/46mK9Z8PqMoq
q3w5h/9uOsBSIkWJqeCzXoiaO4THJ9mlFOQNq2q0S/45RutjiRf6Hj92VGhsHfxFDltN2MeA1uUf
mnwLGf6/8bsMUy/x7rsjIbuy/6Vb++Rcb7+YI5hW4GXJ+jPa1MPXNL7Dk1MoF0bLnGB7aI6kCPva
tJG/L3215Y2ogLbJiQ+uG693miPIWIbsjWabPSjxJJr51rY8iaJx1tu6KBTSpbFqn7OlKAJXtzis
Ft2cShHGPdTLWwQ8QNC4hfzow8w49AxDnUCeJd8ov5eW2ZVCa+OOlxaympOwiCxSWb947sdnETQh
hnA0/MVzuNA1MyS+bgccaJ/RWMP+VnAE8+1h/kpljtyJMrRj6El2wAe7iEjfYJNkohaupXHTz/NM
M8Bk+Td78DZyLYuUq6sThoTHG6xLoQYaJPx/DsJwULSK3F2qLsJYWa2VsbgcztIceEU1OWxH7aOR
SSf1RorKrKmqJOd68Zm0m7MZuFXQq28+/B6zMKURNYg2Xb8BEDxLkUqHFDCbGSmKRPj4GfatIje1
tZEa7Q3t3pZTY1uYs2vx68DwmC0lTKokg6PvflCFdn997DJGIJ2c2GMnVwxCyT20Z2PxX1aLCIWR
kwpkSIceHL8kAdJAcryoh6Zr2r84YkuIKJSAA0qeK9HaCGv4JCpYQ7HVweNhaIDzdDSO+ae/mXxP
pMERKyCxIaAcqLCyCEd84ya1pwWBjT8o4HjI1trVPrTGBVaug2mKj78QPVM80FlsCNMkBN30+1yS
zTOxdSpWloU3oXM50rTCKmNpfng6jk6GpI9RLW42kI+2HP+0/y9VIOz1/eVsdxe1UOKdNYZNDGvu
4Oer8zvK/9WSwJslzbgOs4sjyfMB+5kk62LeV5++VsjT/mWHnBgjizuci3jF3hRupvJhQ1c+Vf6J
+9YeT0jgnOaJcL/r20LaFopi8MLubCuEPU9EKoSsFxBN5qK6qMH6+xjPVElCzcp/DBRRH8z9jN+d
PP3IUY7sQvVKGVyfJVMlFGW6WZTmOlipxSGS0fEOtqr6b0MRjlUevvUunABS8me4I2RyAeMoj47k
MOT7VXukEzTpQxWb9NNDZIYnceIjeGd2M+GJW1eRA8XqJh/DU3FpLTiyniqzLXoAMg6l7vlgojrO
dBn5VeWE42Bu4LTUbbHzNj7Uvq3jZbFAPywnt+Q0kfpzMz0pV6B3o8/HNReCNbwdbu3gL4HWSvXh
p2iWX/N/1ocXz+ZC6NM8K9PMeLfi/vnF62GUNTQIdFYbpiQnnIHYZH3JXiTCnCncdWFKySWZiN4V
k99pwqfYfJnupmw5HXzHK6GT7KieCgSY1Trg7gjkscofyHPfjkfrOCOEW0uSrtEOE23ZQimfxr+8
2ZAc9QHZwCYZUMGJ9mL11rQP1ZWolJ9uXrABhDQ/iKfAuRe3G83wlwRFx1fIcDmWRzxmG7THC0ZY
vnfg3Ax+9yMXZZ8+/TJCuDf3iUEtM+H4GMTNRGv13T4YBsSq0U82VqzlITxrU1SDYmauOUYEHEJs
+ZaNC7voWvIBU729KBo8/2005OTadUYpUt8WUPAirnIGk8tU7oSJbNB0TxgXizEPX9ZAYTVQ8v1h
SUiFQl3VQ4gfE2Xeo2s8hBG4NS/XGqtf3+LoVGLlIMcJWqZU0BJlCl1JNUiXhbSflu5zBB/JJpJv
oRxh1YpeQQVby6NPRgjc0WzS4dL180HcLSrYanbuY44GwYgskRnhsyD98b/EDMTUTq9eXNe+qevG
+sHl7+jAOEuW0w+442FRlBlLw5pTlK92rqRK6+bAp0mttAtIfEUApPOLcso0gXDO9U0pEw/GwmWz
UObdpk2N/uEiVduwlMLzw+9ghAcQz3UZLyKCUK9JPFMp7iPVBhQR4ycLX2XdmwRf/pXeVDAZPi2q
2BzVl/uUECuV2ndDRe8mpf7VlFU5pN6lNEnPigWyx/D6CMbA72yL7gzWpS4CvRn3lRRXTJK1Vj+R
jh36BDKfznzAJj5e5vZAemC4BcmDGOCyrRfeY+tw7XIYFn3uWr+dZb4xH3Z1osM3dQF6bp3yojyw
Hy6BDq/sg/qUw7PDULF5IpOBgpx5xTFPbPA/5wVa3WC4fxf4Yw30WS53rZ772ssSsDrtHVfzlMRg
RmcUFsKQtsHmLlw5n0oWeezEc/iH9Qo1xMIOHJp4DVEYjP7T66BVpqlRKjCAeQUB8oasaMqI36T5
7b6O54Sd2kOKeD4kdtogqMFXTYNoGO0VVVKQMZjpwdMyk1TEQdNq47Rkh2XKRa/Y+oqmy0u5tw4l
2u1o+i01tlafVixLFpovM1hefOvQKAcceEarrC6vDPgBrXSLlEXrze8O0V5IleQDlsWEzFvap56+
49SveDfAik0854hYHrAh4UBTbC4zQXOyxTv1+hp3vjz90QGM1TwbzHicSD9T7UTxd4JoVgnc5+au
JvMkTqrm8hjimSm6+9ynukdCiAOut6GA8IFCxrsKLMCf32UFWr49jI1jxwF23zqntMIGsnYvMDCH
CFtdDEJ5zrckcdSj+cma7e+4eds/MOc9t2YrqOG7abS3wfHbchxhkWOxhjeub8ZQKnaKzrejC++X
wOsVCwxMCn3enmZaUJI3zbKeI3zsDxA/udkvrPol0K/axI9G7GS9syDnHTxyOi9LGmnOPXM6A7Ea
NPHIiaIy85sQFSpdmFZb0WOfMaQDJ2z2+ufZTShP+9jBamCEvhNJ4KrRwzYJm3+SteQbQxDU9Lmm
uMAUBmoDu2Saimt4CVPq1xNu53aHo+BdvB5KbyFkFHmY9cyFAhLRqy6zY9k8I6dX/gxYNSbZDZMg
ZMJzhTjgFGWefWH6NoTViGDax44LIGmVRXzk07cbwBBBw3Y73UvyJSe+0B5l+8SNlHEvWNWRAxPu
mzhOS0DW4a+gvH5tvAoydxeNaJ2ryWNhz7ETUDdBIsNHPoSRssI1V6S17BSB05Y3DgJhG5CC+dmo
4cMkb2Em/HrCypS0bjZzOHHbLy25l1SaQKwWdoAzwUURbXkTRMfDtSfCzlZOAPQHnl2r18TtcHU+
sWRD4iI3OZ6bdXhJbk9xlpBwzG45j4lmphKH/qkRZvgOV1Xs27hycJseu9DJquTEj+/puNdBiFhb
ipQAz19K4ZXL4h0OzsVC5xMASZaBcW4Vx6mnLwP9aXL14GX1+hxn4Oqs11sa9egQMLXEydBS4gQp
CUkJykfosX8lsvJJvJVLdmANmWnRVr8g1sXnIWRmQ7jQJuUrCNpuNPK9irzvorgNopgH2uIGt69g
xnBturMt6zlcnfhw1N0AhzHCSNR1hzbk8AnsVVrlRwURbHlNeU66Nv1BhDJuzCi9BXzTK8EJ5KrE
wXghsxCZegXhXtljszYuL/nJduIh5m04Q8/WMQ77DQVUkZ9l7qdD5JtdDQPSQZ+5f9woZVZfJOvi
ePGwSsVy7fRD2y87eKkkrWhwCZwAiaBRnv0xCMNWAmO7cIju5kKKtdUZKYEdKgCISddWKU4+NOrP
oC8Jvxfge+Ivyn3dX6FinMghdxdvdm1b2Gf9lez1RMU/DwHudxGRhE34w367VXNYpE68kyGcYye+
IMtqdHxWQrONcInky0NMs0l/4RxfoExBP5P+azos/Ow+V1uBDfX7l9mBEX020GWpPzg++XzcReSn
8dM6sbf0MxhLh46iFb7H9lHS+DWeOz6I3noVsCjob4JFoUJayu75FP5KofrL0+9w/+1GcDpeHCtA
sMgA86VHlw51+D9+iTUDHLB8KpuoI2fb6jlzZ+U5VwGb5y3A3qZt4LkI/8i+faohXau0fz4qS9Mp
Vgs7kKDik3Txo2lI97jO+cRr27r1MxwDBTMuoZbXNaiTDISgiy5fbMTt34N/dy9EGOi7nfOjmt9H
kU1YPIgxxMxoywusGm4DCB8/i8gkhsxzDf0nSIMWJNABk2UaMC6woOK6BNlnRBlypmX//Kko6SRY
jG3lNiK1W+PvVeo10kNs5M6UqXV/fQmb2ENIMswo500xsRs9pX5yHEGmGps6HeDHjEWyNKHwfFgA
4M1pHLM0VHtoEzdo4IgW8ygOL+wBZiCgTth9dlJcOMSV1Pl4av+T5Oc652hF+7G2A9u7xeB+pSSz
6iwA8KeiVxjD62LYOB8Fq5j4UdWtDMcsobH+Ps72yZz8LHjpTz6r89VAD2WwC9DN5gXOwjGiLBBk
+2fqXuUyl16MTIQAMyYvZwioaEBZJBNZ7Ef9b8T942j83rQ3CYvKqhPt9myY1WGNN6XSKqrvnU7x
F1TmK+2pkEU53Cux5lwxrdceAbkHZfI+FVzWG75zpGam4PnyUHXca4gEwcZr9XsE1iB25ahkk9l9
7WpvkT9oEI713KvGP/yHE5bTEK39q4XAGFEubj7hKmPj2nBjGrJ65S9ncgMR9sl0QrBGLb+h0HcN
66IZb3C1lYc5Vy2abe/BydjKP1nObRprsCv4+k1V5P/LjkAPSEtaDANaMKqOPFrK5IgxBseWhLo3
MDqLJ8iK84hAxfelbbonhcWVmmwFWfqbH+8pDqKqOL6qiKcf4eJeUicTnPa4W3DgkV6/yB133qW3
pOBb0Lj4wraCZR0GrKizyjcg3OKofpx0gXMWlkn1hsSCzp/eSLXKqVINgBGD/PA46ygsHEvDRjq+
ZdrdivFpbIQYHhy2vQyQ+g6j+WPQ6rdGXXb38wkhINCwv933X4XrtdqSudbCdt82KnvMRvpL8Bka
MmQZlm+VhdYY6fPWL96mraTTYl18T9L6oWfHY1SWvYjkt/OqDFBOeDd92aikfgWNmFecpzNH7xJ7
VCYTz/Sim5wkq8zhpoJCiNfsOOAbFymjLgGK4+pZ9lJdumhyiZ0W02b/IUtLnNwrrwEHKjH3t+zm
W4bY5Zw4V5Ee19pDmzl9yc+YUJUIcrkyMAAOH/xwavgjOt8gLcAkoyGrkS9Gs64MvvnhhDJvQxvT
N/sUuir3tGsaGWkCbE6RPRr9OEu7zuf1OBAcJ1TKhCcHIuTedzZicHg0AZEfviXZ2yoHkMWj7QKt
HJkbO0DE+Em9vaenBOfp0PWpe/FMVueXpjms6We3jbxLjLp2S2fxhNBLu1CLB/6avEmCzENqsOEE
IPcvtW/MelYuHF6zKyGDvuiLv2p5INhQQj89DJugDZzrSgeNCBIEy+EXWtIV5OB09u5Gh9rCdxl3
mwsU4m+XxzF+6rtonPbcmc9+vHc5HN5Rcr3hYesyeogTJz+B845hz0ewUlFx75zb/EQIlfpGgnZm
IvqLgq6KTIJsv1bKz7PckW9qRiIAAI3ee39O4JDaDItV0iSiIUWWXSeQrn2GVhVL0UlIAwfCmNzo
hfT0BK1dcS43dfUuZgO1ATf7E5lK22ptdLRL8v6cedBTr1Xbcl9oJ6U+s5TmdePCsxlWQfa53MWI
M3C3uJoCunpbFAhDTafiR00LqaFGgqF9eUwUxgV+ZVPUA7OhWOh04C05h6TZc9PCtY8tXv6xGtBx
RdT0l3VgQ6G0HDF+ij4VSTr6As34i3xUPKUTQSbxxgZLUXEe+Sr2ocbxFSjSR4rXrXSgMkyuD4/q
wwkKWff36zSqMHj+TYxExEHmZKZjbxNDRd7Q6TK9XG52+gcMEoauxrFodMaF+EFj/qGJS68JVHzA
4ZpkhO97NvyMhy8H8I93Y1Z5l2ItiME4oa/2D1mj753dW5XHOsNaMxH1g5lnJ2fEfHphTmqkWTNA
WXq94aUi0X7rcDJKgQv8so2UaI7iu7Zwk0zsP54T/pWECr8+1iIpYy4ILo8JdhTKaAoj6NYGhqmB
WDCLOHZu8FpJMXbyM+hWgokvg7M5z5tW1l3Sp3eVEpAsS2e6cutntVyUGn7ogKqhfWvLGJ2ePwY6
CH8OqPBYciyKnokAGbQI7YgzUHwa2ioU8zjtuzt2n7Alonwiv57bsZ988FnG9b/KMWgUngiPZsWt
f9O5Hl4bNMsYt5NTRMURHJIVU1vMDdyWATzHT0WgIJRgxBx4+AHb5EFux3tXUNL9KmEvctInIMUw
vcnlfsmvaxtRs1o6UpPUEPFE6RUA4J8Kdq+u+ZdC8Tt/HgOirnrQIxD1GxwXLdGJF6+Sfn2V+gJs
A24l0xIz+NEKXG4Xz4Opm+S7I6/EVws1Ud2jey1OXophcR9bWILF2Po/PNFySXRH2krBc7LSuyrm
JGLTXTtHyJYiFp3EwI2xb05JQCXm4hYljpn38w0g2LlyE4/bhIZ1E1ngi7SsOMpSDvRFriBO3IGg
BmhZKh5kmzNkYMGg9S0C0ppXLUgYzXIP3oymP6HPvG044AaW8TwjRztCu54NwVvWv3rOAKCjhjuP
BqEA+mASew2aAvguunhXSYZQn8vEy+TORkCnSMBX9fSZoOutXPDU+S6Tqvnm8vEnlPUNB24MWfKj
UmvZxKE+VBLpRjTCgTZrU2pXEPJPR9WU8tdMfQwEjjEAR+YKhV8hfrnnxyOLACXvkuz51MF9kij+
kcHukM23xz7fob+wO42NJiX/91AW/ZsULqgMuMSATEyqD7u0E8uUyPcpGm1Ura9hBmheKMz+uFd0
kk/B3/Dxh9aiFcLUwqPNmNKuah2npRyw/Ki1pPW+GTNuCwp9P9VgiZHZnsbqALwtOhfDoD/BKST3
YS0Vr0NW2IRhI/ZLOoefNPTNZiPgDwvLm6oGCGaJhO+jDrF3aRkyTltJaO+wJAVPrn9Oal3CNKDs
CJuHCkN/exfDRuj82t+diO8OIu2WRY4Qogv+IbYulecWbH6F0MKW11HL4rwPdsP9sJZ/yhocZsu/
q1GQ3LmxZ6QCrs70xdLjM4AU2KSGqA4AvnLgj4FlL4ZUaZpQv97a+UtOPceO6MTsImdnM/Ge50d2
t7+HPXuCKaM51Ko7xdg6Ldn/JPp93vVLZyvQawybYd4MI0Ty0DwHKavzQaUPvMlfvkHvAc8/sh37
SpeEAJbOcm3OoHcY82uYEdSNwQvRK8UPosggOXQNvOJJnrU9kesG3TKnnSaSkoEQIVPjYqXdDkve
beYbl6CFWfMQOBppVZSYCGLHmrGezfud3J3yi/FpmkUzmbKjcLWP5Kc9P7LoXX9fcxxHeVHa5ouE
uab/ctJh9Sb/Xds8/e10/NtbMTGnqXG3q2Nr8mWkQyJY+i7vWtftAJF0DElJR5fPIzGs/QpdhM1H
cey5MntnACXY16mt9wrpOkepUPBMeL/v9BJDWI/UqQF7y7TMmPQ3kjUKq8ErmIEdGCd9OSIiRM32
52j1VOiqAoOlJ6VReQt4AAlJsXcW9QKUo8+MFigObmWStLySYt04nLXBwaF/H2X5fQEK5PNb+w6w
yY2/dtIJmQK1Vg6ef/ovOjnHdV0DofG0nr1lA+Bw5RCPMPu2zoxQ6IVqweGA0gurRV0UhgGSaDQQ
n8Nfd5vcWXPLMO7F92aUCjed5+DlzKHc5+PM/S3XQzJmfeFydPmM3w4h94dLi3jxt7B1JuZ4LlJb
tJ1/0+SBAsEceE0UFu+UReaDQOJMaI+iAS1vQA3GI9rJpPHUGg8jvkdubv/Kl/j71AB/YzbboNM7
3DFuIVEm7Ld9aH3lKPnFyur84W2TEfjrkjzL2EOii/wGO21AiLiw/0qofNygkrwUD9/3SrHmtOGO
P7BoK2uP3iEpHdobZJTaPcap6QJP1sQZX5t1cOqHQ68Q0HO3nDNH/GNqq0n75XzBRRL235PbnauP
F4MDhA7ThWvP4qympg+haNjnz4H20dwEvXIBM7QqgYE3u5ZvNdwqIhKjk3bFyCaVmKQrc7M9x6ca
vrgPl2CkGDFEOXfyTgceUf8+mrLLPFPGHUe3AQVx2QigWNiZ/uqJnrs6y6K3Okfxe+FlmRs0r8a4
JGasGwdsd7qpYLdhECkXFphO8gcAGW3E8NPZoEoF53pNTfB9p0mGh1dRV6km4kKosw1nSmFBBveu
XukrZOi2UVY0iwZBB57PsIFYRvbXpYuLZTv5wDmBFxCm0pRrLskjuH4QmaN/bfIfafEzargYD3+m
6X907gPbXLENBS3pPrjr+EV5x86hEjQm/ypHXrDhE4c+UR4j/hXfnDcKxOYveU8h2enL2w9GGlD9
/BSKtuQOl6sQBAyDnGpQOu1SXAkkCLzFAcWtx8IbZ4lDKeHLSyqQn9ptM17rawmAmnWbCgCPah1u
Y7aCmkhIKL1YV6t3HChWHYDYPYsZODrNdjsKuC7tEQ0LlrTeLy2LGqOBrnuG6GqywaCHEYhmS9vG
CAfX1vsPtsqiD9/4RF90vYTVPYv9wOUn7g9sOUbqyeEBW+vAoKjikuzIbGjKVmwt3sRl/hgpf6gh
GxWK2inWNMZAjLISslbjLe8L2aLDR0u33lnE8+uw40s2MeXdK3+1oipC8lkFoFCRLuQQK3l455/+
U+sgmXYgYCEaAHSAhcbcho+PL3Mxf6bjC2sJqoPuY0+KFLYIum3BgGWtR6oBkDbGCNQj9LGc4hAE
rw3jzk+uyx37c7I3DSM2gEnNQT41uKpgZnvBuQP7JpY5+pKunn3JGjQaxY/YjpZwxxfFeQmzGwDZ
G6ur7OmE1fylKWuY7SY3StoUPF4Wr88oRIxRN3FudtOPeyXlTnJDqDR9AETjqkGBJZXeTPOmt9f9
8yyby6eCRL6bWS7wE/D2vruDrR9VTkU0GfOHuhvGjc07uFOtxIMxNCKF1lkC+l7gWiZHVONXxJKv
DsNm69QORxUbgPujD+fayKbX6rePmMe2ChLOZjms87lJd09A0TbhQYUf2B7POj34odBp7JDA4/p9
23cRMaBcAhM0B1gx95Amv7MVEnkvsqINqXIl3FaSUgY0JkJXD6n94KHbVcui/V6LteTVtYdclP6o
ZOtSirKB9GMPc4QBhZpJckRpnoBMDYUeal39So0BRBRUVQZTMSUJM6tt+Oez7H4V8imtTr80/8Dh
GnP9WkH343dplWHjtBW3vg+hGslhuuNKNs2c0Z392yKwzdaklRhyYtnCXJjkIseJFbguuRSaiqI+
Bn/MWBtSFHM6gzWJz7nX/LsEfTtgkFHUGvQWg4jL7RqjTqpnFUIR+/6EF3r2ctvPq8eZ9xLFJMhA
sFHyoWD83Bxn6cSHXhKZ57O/7YXLvi5em/2ojvFfPvfYY0jQIZGLte/Pa6f5DxJ0na3WZhSgjM3w
vOi/mqoWtU6Rz0Njfr6LRYEG7qTdp01Kn6Q9ugybK4KyHZ9DAG+ea25AzyVsv9q6oQrvUMsw4yGW
trHLEekCPRRjvmm4e+MOCsyXbIA8HL4W1juMkFttjnJ8FkIIBRrE24NZSZ5Bih0WfauiN6TN8Rkk
szxfPb7wc0O3p9eeGbpDMqcH7rUF5UMlaM/KYVco2dqqUYjVw6euG4eRHZdzLX6fpPJOzaOZLAfQ
a/7MojCWN2rf3uE4JQVrqkA2ojq/P9pGkbMWQusWX9XI9guRodxyK0SghK6vhM6OxkK/BPQ+6pmF
YH228doukLsMDmWADKqOdFBfrhyFS4qVu/XJ41qBY7gzqzlaDLN23vX/yJa4qCWTib6hGpj6mkrf
ikWPnJAiwcMID1r5G+QqT2N5SEIDruGxMOjX6zHgIDeye7sP/AMMUbK2nSXngwspMkMgi/mv2mc8
1b8izocNWzRvqtj7jAL7l0yquPg6Ti3aXxW4TunOUhkxdjfuCa257bM/hkrXL2dM6D45q0mFcGJ1
Ez4yiqozRAAfk91WbinWCL9Z3X6Wqp8bU8Rld9Kfxcp9uLv3dNdGjJLUzH+83P+XMOvjrUDHJKFn
ka2zFtz4ylGeX2E9TyHvgZM6MhWXZRlkf3belcmDOwTaGrpbApiQOYrKJ4Wj+kVwB33NFSSeIxpO
q/hcGIJNeVOxocUvQFN+zoiuhMFnOUJWv3y1OzzoMoDicP8pScy40jqiqWlngcEYnAvEMU95AuYf
Ys6X7AmqFyAQmQ92BOTUI1bI/uG+o97Tn0shwVHDwvPLK8tiyH2+f9nXVoZnOHiv/hs475dCkm0r
D7SfpWPK/GbLgTRnLDc7e/dJddvesRMHacd89/U5zerBTW3Ch0ZHHKOsg4cV7Jt525S+GyejSs5k
zNZ80wDYiC0S8250YqKlS3fnNqcgyAiZx2S/A/RMIp8tinRPG857fQaQIrVP39FaieKqmmJsNvLY
l1LiMuzlyeyj4CXudftNUTvespL1aDC5hKFL5RgON5k9xMxGIJrJ2C0rL40Pj0PJQuJzguWgzVUA
UJxuG6pIcWYVf5uKtYYTnw7POpW/yfT4QXNejOH98xDAQAQz7L6CArG4AX7LS1abLXu9BpCpbPLk
6i6PPdZJYRMISDq/THcdxn+6hUkKJcRiOeoifJRYtMUmwjfWwWWkqpSsgZommQdHvv8ogskBYomx
HLw58r5bUXSz+BJlm2Gq65AbuMd6bYWFfFuNvCJbau58ccY3m7J30RZsHu8ZgwtrmK4qd9I98er9
DeLUBylDNuW2n3IPOwYHQVkCozHI1SIQSE4cteBikdBIV5Xkqs7Ra6JXQSwSGhQuMGdMwDEmfJgV
2YCTUzABjko6VhQdZgrv0qsOzaDsKstSonBED8ZrM0bXF5IJ3wxQTF6QOlYCPCw0ULwcyFufl74g
uNoUiBxYfkUZXwcD3KJM+dzo0+aVxRMIn+BEpxqJmd2cdlNONl7c3xI9Og0hJbZyJkBVqxpd6BZY
OZ0T96NwIPOk58F4jIFd+asqjn8+mkKxql44UuW+Z2UtY610vpYd0EaVg8neU97xKumw1I1Z4uIY
4MpBk732Q8DyI0ZNfdV67VcVix1wWOiPm//qz/gcAEy/BlFsNBdxyF9IeWK8xRUZS7ExxJ7DnVak
7OX/ObkrcQ+47QB2YFEIzwbZICw9TKnT75DbjEN59zFPVN92IRXNe5Nu0kE4yUUc3UBCflEpqAZw
Neo0ADCtBisKhjFfzSeU1Q2pkaX/sQfwdOZy1eb2NDb+rE2TD4lwCSAlF32scoVgBAxggYpScLYC
1Mhj6YLr8i8PGKkYlOglhkoC4pDTWWlq6lQprdCc04RYA1V6HILIitQVmpckli6RfnYqJeebjY6i
J/22mFOAmF/gzPn5JJBdfPyozR9+Nl20bJrHHTUKt868dJ2frNmjB3ofO7sepd8HlGq41lrkBbAL
1hUo4k+ShlEK4T0W9HpiLQCsJVLFzm6Ttie0UzvHqRB4KLY9ygwmWwYiZ2zzrUyUu5I0jUSlTK3V
V1FlJ29tfN/87R0QHIkqKqDU1UMxwTxh4E7ZfjWUvpiTC3Ex3xozvV76Knjh33Sy5bEYD/X8m+J/
4fg2TTqgSsoNZPESnOXTa6XKPX/jnzAImw9gO6u8gXO5cm/fbEH0piU++hM9LI/nRonbw3OtdMvY
IXH2WraPce3qvC7CfuJaA4lWHl7H/DuDNU5iG8iv3/AGn8PHHZadhW21ZiHKWqrVyk96SvtbNa50
Cayy2hkb6wJhCy5edZabEIuiMAW6cOvO7oOtrdwRpoZQ8NKuIcVnEQT70f1WkMFCpSB2szvR3AHz
3THOUCjUb3cm5fZDFXCz5tLLDs1cCNTlHVM2BdWdD88YRVkWeryIdXD/pO+zZxatd0F4IRjr7xVw
xEtlIBwUtbDb3FrY5kUmCEb5gwg+mefWyTDb2R2ePWO6yWm515C/YEe2cM90IZqLwgGsTLjOTRrL
jOecULaCKRg1lxm59Ugnww3NZl0mfjNcsL6uqNuXlzItukHPrWXBFHkbZ8Y5snvcPhxNKxedCOoO
OMYW5A2qk+p6yj133gYdL2Gj32xQ5Hvdy996NW4nWsGB/qA8DEwb+04oWoJBZx2EYaUB0Ay1YgGD
7fSqOt+QtAaWiAHL/ST3rt+usOrQq2S6hnWc0XD1KotwkVfUXwAcsp2IuPEjvEJdGFsdNUq4QzFN
QlPtzga9pHC3tCmNHpgX4MLQQE3R12kt8+qcuB/2OCwUgyva69V2HszMWl9pGItr1cHb7Oyl8C8A
GHLmNTk4ygVPMkdyB8e11uFKSpYJPLUNlyBWpQfSbNTvJP44V16fAagFl23dWHXXdTUOsLwpWFhE
mIVvPWCm86K8d49z9Pch5v+EViDtsnsDZkzNxjz4NxUncDpH2mq5j7sO4hjxyyC15uO3pgt62a/T
uvmH6695iOFezdRx2mG6NNNo9ccwlcfV4YQO8KG75EAlksbxfYGCaaebWs31yXZksLw6veBV5Nxv
5wJCUk1y62aWBl7AajlqUKk9WBnPfUJdELxvwwbtcbZICjkmrNKDa3p+XrBAMAM4DROgO0P4Wv+K
RmIMVGqn5x330q+u+nEpZf57FOUl4FNRIRhrASAo++ptESqq86Y18ayjlq3S4qlx6T75lhvAOLUo
UmSSnBHOB2I1PplMaEnKBlOZcCc6COdhlNmi+IM4rraU4QAbHZyBsgmeiOt4YppMZR7HT9ZSzfPi
0KF5eMpEJ9etZLH4LpnxST0GBXeKADM07yR06tbbxIZ2HcYhIbUYSfBLkCWA7T7H7tGx2Rl1l6BY
ZRcwmoiPwQkm0olvEx69l/NGlI/vo9JzAKWLrIn63i0oFJVkAOFLreO/cpqOf6tzzPicVNN+v4Qy
UOV5Y6jr1ZzY8bd5FyjKcYSII0epF0upYZNy+D2Ps8y8yBrjURclqUmLLiuL8P6N6UTml7QGawTx
gh69kIfHuzXO86dc8LNmaIdm9a6LVmmraye/BHHoxLpeGY/MxfGCcVSgqCkNU5/RMlNGn4t2pWlX
ovio8uqk6pJaO/5CB+vKbNUeCgiKzZ1xSzGUDmeu8ouzwbTWGeMXUo1kRWg6GQTysq+evPB40Y7S
yFt5luaAoHV247FNEYgHonSLu8B1/EJTXJtTRmNYPDOP2C9nL6rFsKFbrzsi9I6xvWvOxofIJt8e
MCjGyaZZ3p0BN7s6xQwjLnoeIfROLl8E8Xr+COFjnYmF+jbxfdHYL4rVt2eqAOBsjeiF/qdAjBR7
dcoxNGGKTV55ed1z9vGzmocYUWG8E/mlYvlyRPaxtRL4E+V7rSTe8d6wx4npMbMaU+gygXQzR1Wq
fayS6v8dNYnVMg2ixS78SIeWhcYZ+dRuR01tLCPkIKGTVvVrYznInO2SuCGBUIZLRK84rFB2U1Xx
keW20B97/MBW+d36Ch3OvhrwOgKiR7ZjQ7HpX9gw151/oNyP/j9w/mSkGhrPeSBLVxVJO97Z7wue
StP5r5GBr3dLFW4GYaoaAG1J8+1ewHc4N9GR1KeYoyDn95TUqNee5bDpEb/W1gqQhWmaxw359z56
s+QxVTcUOf5uIJNwbHai3fPgSU2iWz6+OBRyX+1RUnoaFj7rzXgfa9LBQYDniNwnpvQkiCH4uU1A
A4YA6ePL5Nd8GSGcm8u+7LoJE9+2SvVqpEhlQODKj+p21YQgKSrXz8DfUNCoQeJpF5/FvQxKKO5U
ylmbNI9Khodsr2QkvYusRxfV2WkhADpEfmF936NmPcUXCZ+M8KDi7nSopPCYBJdn7aZYOuU6HzkG
VG0oC+NOlZWPzVARWtwKRbr/6UuYS5ntv+oMlgPIb63InhrOwPWtucLj3K0mElk1rONuj6yUFtEy
ZHJ4D1WhoHBHE5Joq+W4NReIu1+dkjm1/UcNT14G5R2aXKVzD7YvKj8RU8r28YIUQwnh1PHNhFTv
y+MhZ/C89SaYhp3qXjiDnCClzXFqcSbOaFURYsMrmgcLFs4HhZpZsk9eIANWERf2XZ/hEOfc+LAF
+LaXIzKTKU4Fj7m4+r9X1HaPfwH/85bg5ker26Xg070ALWPB2j9gzvKLdSbglLlZuKw02IWwy8VW
Ep2B3sklXuBevjMwna6lLCOUW1gVjQhyca11kUX4JoF4pDIsrAsibVx7iMrv2EAwd97PiPIvMdU7
oGhUClyRW7VSO9hwwKewY2YPhfi68Pk1DC0SmF+/zl1Es3QOw0bFJEdqCDhOrZv0kljFTuRf5Ips
L7df3IR22Hmww/fzIuEkZl+mL2uGMgzcd1x+RCXg0E8WJbTJO/PrGOkND6P8b2XmCQmqSYcSxLUR
yG5a/L6w1Fle2BjSv9exIjXk0CUQZU7SJV5xh0TjbzFI3MIBs4M8NXsQCmcitkgVXnR5Oh5b6Jht
8AxPb4Lz8Io1Oj+ykmAes3Rn1OtwLf9kKbjrx/dTed1j3xev1WB9amQyZnmRGU1bWVcM80ul3uQ7
Cgo87dzslBCN38XjppczLTNj0B6jLZ1U4d8TqX/nfxRCQ+3miad7DaHxB/vp7/6FGYW/1Sg2QdyX
OwYoMkN5H8STdsXUOq18+LKTmqiNTvyVBYNdGoBsYC/Y2JTyeVcHtNHNXQMQUDS+mbOJbq+0rFDe
q/oyzc/MK8tkWPdFlqGANyMXjpBbMLNQu/IhdBUzJvmK2MZ5PiNkLu/KWKmgYhU5Z9760PxGiUVK
8acrsUo50vDRdFMjjtXPy/YCVr9JAI1GL53Em6E2UKsMbEVog2UEf9gB3ZTSMSrJxpCREpTfPrBq
cZCmxGV3sIUUH+fYpsmdUBs6aKdzXdoPx3WvKoXUdLG/62yl7GRXiOBQYa8UnTFp0ym/MXLE9ogG
gHBfKuyd2cT+0ftthdV+v1zX1Edq4OgWutoaxxLBgdLAnHkxgSGsVW6XkqZ9XiqYhP2945ffAcB1
u80k8khEwNnay76Vx3Nr4ObFcnbblP3djGBRGyHGR5aRXWx3EqDDmtyJ8tUHaWJhdlpafsto5CEp
SKeisYBOBBlVxrNoshCkP/2TlSgEtnqq92+GzZU2SSVo01tYjFZNzheLq+ZrFD3godmJYXDyvxwt
0E1y+cWEfvnC6/uGbxbZCaDOFJet6G9MoCTkbFRci+uiLA/opRtWIlbtnGekCvJYfSKYhUKzvTaf
VxBSqs0vX8zY7sPTZZJ3xzuTXCdcLXYZP4Gp6Xjid0Nzmp3Rs3WvNld5L7Cic7DeHMcGPnciqob2
xQ7gBzh1PvcU9ZThSLhIPUYMm/jpHi/95nxW0N4/DK7jkMhGr2/nWbp3wslpUojh0hThPz+at+eZ
0eWn/eyQjP41u0Z78gcpit/kc5ExkQzyBZEZASiQPMD3Cy+G3IWEapivclXefbeumLciPwA4NSy9
tUZ7EV3asAz5gkGJzhbiFOxIn5SppCB06N7oHce/PmMpf4HgtvLyigZqrDHI13uV4geJizVVyFLb
Tyt5MbI7qXYqCGGa7tBCdkGyv+ElVaNUpDFUBJxMO2K6A4J7fw0cxWrrUsK/cw7Mvt+0Aapa+ARO
euztpHymWYV55EZ4oL/h90ixZXb3lyqQZ9C2wTXNUBMe8oJWyRzWUlV4uWv1B2Pqo5uJGKbCyb27
DiNtUHgW22xEk3+bhEhon1zSL98jia+KgiKz2Sb5w4HRoyFV2f3zVXqXhMzgMJ89SEEHCH6lN5pn
vq98BRTOD/+fBnMVXqa7OPaVsxIizXAyVBXgxslqAlqDB5PSxeNuROmRrWj91tursgxDoA9oMHRk
aUHnuTizjYuCa4XhcJgk2vc/ApgcuuI0tV2vwTgsESrDEBo9R25GQk62bcamLL1FsRxpUtmnYxM/
kIAPEyQoGlXWNpRX46oxwOrO62KPo8p9hPc/Ts+Sz1/tkga4ZYgO3vN4OnWTyPGG+TS1fiiLnF2d
1W6Yu1B9U0QFBd3YRYq2T6nzr7MtVf2vkkAuZfiLT5jLH4TeiycsUxkhaJJSPVAAIujYyiYELL1e
5FYJr8ScPbtViKqo59ltChs/E+LRe9kb/s225Ecby317M3jKanOPIWT2sVa8ENrj7Xwc8veTi/Yu
hmbtbo+/5WNhtjoN6Gk3e2t/+0yfMj7HYtV0EV4bJdqBnTyqsP1o3DtRuj5t+NzaDEERod9CHgiI
vKAyOldDxnqbEgLxO2Ec03Oi80CdDOImAoo6qg+AdLsJyVLs8LaYAyIfGnrvwH8Mfi6itFd02uPu
Nymh+3ywi/nK0C1ZD0rrOEKLHkzyfuVyz/iKSODVcGDbSM/zXeKEvi1vjlLqcMy57PDI9UobFI/y
wvf0KGFJCrGmsH+bECwgPGaVw8WXkKX3Xt4sAPzqDJ7/w28Ch0XJcRZayXMWk8oF0n9QzjK23RWr
p8z01MrUyMrzdbRyXuoaCpJwUs8SJTn7HWs4WYZqfXmaF2BnugKyzXvxPZF3l88ZV6xg+ZiBieqI
x+G4tH7iOmZdhQs7PzINl+VzVslldMWuX4IFqVDzPsqjTqJQ+ZJsLFGJzyo9dMqxkKX09p0ktate
s5zinrlccqRymOys/zvCD/otDMS2WuWosznjVug7Uuj1otKSf9/KSabydNTfqev1zC+4dB8Z10Eb
uzidv8ce7b4s0amWq+mh/Ev/6tNX7Cg8uPWbsF192ENSnFpRyEBvDqjlLuZa93od7qzyhapujuYR
ICy2OWhrGT3Gh+n8jWaUiA64lBeiB9g8ZT7Nf/hG34d8xZHTvI+Ti4Wj02TUpOWWqKoDRHdO+qdd
BOd1KkrTcVzH72+HVmsVRUiQvp9deUXVVgf2+3wXjicrScjSYjWutF4jEOyBw/MUuKuyu20cKQPl
JvoiEqJQGm10Xh6hKizgs4pSmE4f2+VySSWC2cVPZkrcCgxqG9EvuRrHMTGh3uDyHrS+XOYPW5ZF
b+CapeLYhrTssu4yQ5Wso/U1Mu85Qm11I4zwGGIqm20yl+DTW3FBJTDvl7gPWDtBn24RQX8ggRF0
XllQXE17pEGW1psyvzr6T6BxCrf2krVZ21otWh5MAc/3kWU+cijRtmhvW+T8H3FhtdmYcp3PAudX
os1QE8Oi6CZVrMwjp9no2Td9iN+opkPEC29H9wFcICzh8+8U/ph0943nlxYaQ72nPGt2JHZ04C43
uDgPc2cXPWF6EqNoNGzlumhBdTSvpWR02fsWV7Jv+biLZ+hTBisCPJ6284fuMpycztlmtF3c/JN0
+sP6pkhkX3PC6X6eyvoZ7rEn+tD0jLpRH3j5wL1Tcpb1hlU5qEdiumXopnPpSrmiOMSbrhLwwPur
bmxaCPJDDzFWU+h3e49rZ2T6FUWKC3Gvas4KZwKom2rrnWv/zTJVKhFBWvIlBI4bAW5hXJV6zs1P
GD3B3IA2P1sYaN5n5xgdFhY0V2SNM4OTMxcWdtDnTPpg0f338AYT104rTP3hf7jy9nKX5F9aETIm
Al3lWWiHBoTL+tVgxnQOfcKVm35jXnB1/5fB7NVRc/DZzYrtjEc03MREkHP9Ch76GAo85R+6ndyp
N3dUQScIJmtHpRnk8hsFEOoQ5g+Y7qVz6bmj1ApQwbFIE1Tk6DaRfBAyptqzxPR6AIuElcBkdoAp
q86wYtoK63k2NTAXcPjvFmUKvVOsAMuW5R7bi/j9P0YX+8csaUXG2KOey3rbv1m4mlClnC4LggOA
YVFUooBF0MsWDcniK3JBiLzGurGcH8YynHEBenP4K1h6r4mK/GgcyhRFV5J6jgNLc2yiJWU/9VeR
ky8ogesCjwHad4GVwuFciB95CLOm050frTej/gYC9XrPULY7g2HSJt/R4Eo47GQOcEaMbeHyCINv
aidRZHkSszos3chKCg51XpuVkwwdVq/PhQ+z+CXmNd5At8jt6WyFRWrgUbcGtCDt9JbSFPsROXRK
l3IFddxLcQy3NItUY99D0cuh6/gbwcKy2RXbRAOu55YWco+Ilwuqx9H9RhWPIbC1nqKMzNhC13iA
2VdRxysrG73i2bSBajCTJ0UFq9oiOuFlllygC2Fx9UtNPfhI13hZ/c6d13IHNalEH7knV8JpiM8D
p0zVLrAHDj2im1uW/IyvrZz1AWN86vVSCVY0tw975CoqJLBCHYUCYE0g/QnnYn5jQrlrQT2ybZbr
THcj25fb8bKZWDxdrgUb1N5shis8V+uSamxRkYFncIe5Nqc6EKJqUTXtgRtHtGbx7O1ja1LrIHpu
UCe3jd3TTkYhkniwZBxGZtysA8nDUdX4RcGqdPTUpmZl/Sxvbx+RecdjYVXbnfFw0cPNx+FUIQf+
q+td3rLCVnkcJk7yDpioRSJFE1QtCp3r3xyEuWbG5RDy01OtpJiaR4AmUZtvDGz9Un3i1BuDprko
AGBVDNPGHkRHB0uFEGCBhLWFxbsW5U5PvMHKKyciajzjHs5XvXISEkXHKcDxATyaDSB94mtgGjhU
Gea0bAXpvLIBcIjFhHwwwDo7xVJfbhF0Hvtg3YI9e8iHOusDiIHdQuaE0TS5Ffqqe0Qt2T+4Mmk1
VZSjBXau/L4rya3bVYIoFXSxJbfsOsVGuFJI/g+Ih3c6vZDW02X65Nwewd8f5eMd24vhJdwFvT5J
1j0f6lsJB5xFZZABFpGCtY/I0mrzuFbslc1kPDYxTDMPF73rz2WLtQCyBb3fNkUqYEqmB2qGhXoB
mkZawL78LpcktPnLO+4l4yYSdfI8DK5CYiuX9nnL9xjV7AA9onDcosffN6131BAO/xiE+154Xp/d
UfBshXQXM/rrQocCLkcpz0YuGZ+IoCdN+aJ9InWM7jlXHie66bX0K8reOnuIvxmRadk2jeEM2CAw
VfacUnC67UCbKOgt05lMwrKc0Pyp0t+RdVbf/g20YDJBMKDEzJuVw0t32Ece4ZR7bMqStLuY2Vuk
4qAi5FaR1sGzWxQxKEPgospWlaxlh0BGyfaL+nXaoY8HYvhpycvpEWK2nyAeZRu91xahbU7skfD4
P9klK0MfRVDnpNJ7LftsrasG+k+Kqd9qf7DxpKaVZ4hEWe4acdbKl8JvwHis3WL9KD1xtx8kol2h
HsGZ8KmqR0jysDC6cXNuE/iDDs+I4QFLJGr5eCQ8HE7JHiW/1eppX64TGSoMLDS2CeS+vU7qUPce
qILaRA/2GtRpXWXAyKEdVxkHTPqi+Bc463u21azLZMegqFURz6UMMOTv55FAVNYzKXmKPFCfPlv8
TBPTCQ0Umh75XRvDhtK4QKNKNxzKEPc2EyhWkA2ofEn1TCzoXfe0samRczChpecmCp+6bV62D7ZZ
Ai7aoNotLRM5a/5S+bqIYApPw7WLvDe8OtVmlwx5YpQCIyJDwNfbfoR3owoi0he09PdoyzrNA1Pw
MfE3lxvzGNkdqQ9EHBv66IJ2TAMqHWgZUYYMR78nrdyFYK8Bh2FUAhyOK3LAlwpqJnO0cNt6MHZW
vBo7z9vU837FtExQn1stiLpp7yAgiPGD/1aQ6XN41eP0a74lIor8uBryaXHww8qiSWhXw1S09Tko
Tej6zu78pv3LqUNIRV31P6hYCyFo5GDL3IPosKDLhjqrr+49rSR5ep2QqKM2MzRXmH9NvSit1M8o
7XCNn/NSmQdFn1TyGp0bKsNlJ5lue7UC7xSVA9W8VMkNOCAHn1dHFW2GSuvSnuvlHlsQGKlp1lrC
hfR8hvVwPdI48UGskjbTho1f+fZdoQpjUPdszy2vC9PvA8PYoR8ISk1d3QMe5ZaBQG6y17Z6yEaB
3lkT8K5+/yBidyZLuGol6lwrzmoA3YWfg+Zc7q2IfnPb1pW+5Ppp9E2nExXOH+PcoSe4dC5M52O+
mKCMprUz24BgjBcmqGKU0RqbNgJ/f8Ei1els1fMXdFQ25CuZ7lLXpzJ+oOFYOU0p9dASJUTYmC6I
6ViRZuBqD22F1Srrafh3uSAcDYD7w7pASZAzYzzdxG2u2x/UiOh0BuGlPzVD2656lfEBfMz6N0nw
gMT/PWjGNNu7DtdwvP1Ec2ZqASu2yBIQzVtAx5VSV0w+Fj9e4Fvu34kSkiHzZtsnZFcrQe2rpg3m
pvRXqku5tJOnhIF+dwETAuBXPsBCgF3ZPFvG9deZWUrr7MVRYfIac0pj0UFZ++WYwnV95xJnvBpd
Jq9xLWJGq/KJ+20vTt4jMhBeQfvKUz4zw70VsDCbNjhGz1KNQQ0ijdvO7L+h5f/gtTOTWl+TXykS
hW9nRHuFKrA4ZARq+kxsJe4ZB/eyc/f5giYJ+h2FEbWMS8uqwH2SdEnPn+EWJW1vSGn13tm9P6lg
A3BDTFmQqXjxyFWOTzKpF3lCuYnFPVbwgtH/e7n3spCCTstvJx6VQ1uFH3QiYApg7//ck9sSj2lM
jf8Ttg+FDkTJHluGvDod8oMkKqersi2blxYpUheofWeYhS3Iv2W4E1QyT7fthTt4hQ6YmO53+56Q
hq97YC0JKZ4LM3zDkChct4DCVLYQTv0sJ7CqkPeLva/D9V25+Z+bWC+2BfN0LDv/Eh03C7te8p7Q
8fwPZ6xW/j3vWEywGh/Ug/uLcKOYVJf7DaeBz20liHzLTuL76PMUxJX49ACobk9KX/7ep9TqJrIy
pUJ8/S+AVA6EaWHNRiilGse9gU+w8jAhVw+HqHyrLWlouit133Srv1Ql0E0KdVE7SLSPysw08cnM
QFxPVqLBBEe3THXSil5oyHTvKGnpPsxiFdg9jYSYC4EEC/pXsuLmeFrE5u/19YwXJVq1lnHe4sRv
DUYa8MEcd0J8DNuq4F5ZOhxj9A+u2mY9Grjsr88xVLG+eJvlfHNoEk55ZA6wozw4L/MjwOd7+5a/
tH6g/GYtqdpvEUDeJgYsqB4svYgiLnoevehcb/sp0iADny181y0S7UdsqHwOXPJv4WLVVIAKYujC
dSVUJzxy700yakz70Baz77xajMF82bVnEHp2X4KZTryRpaaZ1XukEOVByrcXtwTJC0327XsUsr+f
Uveuocx3SASFhhj3bcIaUa3nJEe4TEu/M/9lgvBGOl44WBp1fl2dyC6LrH2N7dFXK0MXfb90nJ6U
uqu7D70g1oASIlWMheRYX+ou3/LWEIcs73pbNiXBNTk0oxWx1UhENkjdNRgfQRTsnvhkJhdFwwi2
rWCaxEkP3yIs2nX4TyaJHlnmpQ49A33E3mHagGlGg1H8dCw04fmC1uXgE3u53JKvMzeHpFVb2VYX
avqX+KbCWZLP1D2MAkVL+MNVfTX9cEqFz+nzUm/nxAlcUgOgcPDqpd+6Esk2Ooq7DecBYGox6Vvi
BJvUQm+0DOAuEBkkvdvCbgiI5XqpryFzp/uUVA/2wRpb1+97l3ZO34WbhSxp1rNDsWqTnRT9Ost7
MRMGEL+W+BReGlksweIa5k4HK9J2oOZsIzFdfO4okbUndwQSf5rmBD9OCLkNhSaH0I434DoQkBuw
Ngr2ruJUsU53gbAHhF4lHx2ErgALpo14hZfdd9vlrSv6RH4Lq4KQ8AxhyUlULahG/WXWHvtnFekS
z3iOW8TfcWABaqxlrFq+kpfKBBdux41sER/GFJ74VQvt+AprJrkVIp8losMxgCZFaaPV4yAZnI1M
b+YKEzGatFfs1RSreV61LECikOa02APGrmSoG13JphjvGRi+ihwnsNJRPakQUr3hJ2a+DU2Zt+wm
ypHJnhf85/X50MNTbOVEOM7HPUMCBbYdIK4c4Att+KSrZ+tRMlMTu5PoEf4JViOH1iDh3ko+mhj5
dVzbi5ca1swyrdN6MkswFqor2F36xyscrRLpxqPwE8Serg2g8QUzB2/4kjF61SE0BWcoBbXJ1GdN
RrNGdw72/GVc+BG6WextajEXljOQ4SI4DWXT39OIblOzlF3YdSFH2Zwhh8rTJ2oFcthwF0Tk8mzU
hrYKteef9Q5DxlpAadM2xZAFY0jOaRHPRTDBW8wd8xGxzPsVVI3b+MeB4QGGomEMM+0WeZWBw6ca
M5GfoDqgIFUxBWOvjZMAOcFte09V+izoSU4CZVVpcl2apw044coM7Gq+QHJ0qTZAamuGywSgt/9Z
dw2tQUZ5krT3mtWRUPehX16wvVlORgE7bkRWlUufLv9GzJ5mDOLErg8lhdb3xDrbbOtCDqQCBulE
XM/kkhAFZLii5ycCoTYAT05RnItcL6wy
`protect end_protected

