

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
J8nZtW1Q/IGk5bZ13EIEEDntauAKqOlRji4Tz7aOFZMrRrl3qAAP4lw8839dxHbOPehATkI5mWRu
O3oQzXKv+Q==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
PO3vY49rlamMYJ9pWAsIelQmo4roKT2hFecsbIIwc9Ce9j1Gil9MEDKbHqn/9XWL2CZb1+nggmfu
MhGokjjD0xhuA7bkrZ61EFG47AtPbrzrGJmyawEAJ1PNLVKIspuVYNxaD9rI6pyGoENRti8P0hyl
/TLRO8J/SzWO1wVCE+o=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Lek8GlHbeyFgFk70bzers4fkqEzZWIlCFJLfSucq9OzFI+lvPoCv9lLJF6jbu+G/Gu5TV4ZuNXdu
mi0r5LAo17AD7VicMD+MhRKb3DE2N3pAEqyDrMS1jasKAHiVpH3eXVPN2AI+lDAVZoDhvjSuQjfy
us+5QMijcCxvAveyXwnL06kT9i9dtQ6hie8/MMqHXkiG7OYqxKm0Iia9+F6bzSI9YxeA8Doz1sM1
HWlzlbYLDBCHp8//PX7kMS2bPsw5C6UPaQ+TKox3agXXgpP4ea6EVU3GCBe7nIo37nZIVwI8YFKU
1lK2hwoX/DoWAQ9zzkBtnp8rOkj66EFG574xNw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
H24CFb/lxJKnebrcZ74EB0cwdvz2M6JUcau88JBt2iuFL0aDDA6OprhhTeP6OvCciaaGRsBEok+U
cbANkg9G0zLP53/WvEkpdYtezlQI3mkakzT3UxyQr7e+pL5MFVi19R/4mD0m4WBOiVFQ4vPfnILO
XObce3WQbGcK+NGRsMw=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
RFnK9ETQkPWYtdMW+yKQ1MaijPhYXOMfuPVBKnsFVaRScaR6M3W3RRHlGeNOaiw0ukl3q+66K1rC
RHUWrifpwoSOSO54nuXmCv6joF0+cR+UF1LUkBtOigSpmJUx9SscdsvDcBNzrLmtogpoKRScYdGy
LrKeBNVoMEblduWARlt0XQCFRD4X03OLybCK5/hlbwAJA/OXY8QP1rB1MFXLkjS4zFm16T1j7dVB
psuynNAT4Rwsqrw26xpeXem+8Ft+gBzXVIL10rNKj0y4I07ITYInhk/p/CsNH9FgAhYM9jsWml7/
R3A8DckKe32XlGviTUqdr3zXyrsrjZFSJ1kTGQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 107936)
`protect data_block
5wArtbHo9zLQOlZ8YpbnmdjCG/XaYKuJKRIBzDgDLGTjypYQLRaiai4UTmkr5DYyrexI/Kh2tzbZ
s/R/AJxJwdbAAwnq65+xeKXD4KPc4UI0nalRsr8RnXJ6hSnP+ihTns166l1Pj6S5msH/uMwFFYmF
XtpNv8tUrDpgWno/IXcSckeX8YWe6UbsxHVlluiYT4LqoUvhEB2ahdiiWNFAxC1L7iz7X6FN66eT
Utoxqj0rA9Lq+gJMDTDxmzmYaaVNc6URngHJOADklxmcD+1A8RhsjrQvK92gi1nnDq85imdhfyrh
76h7O7lN7N3eejm/SrZQQWj8Par/uLktzISxjR3fQhBsbjMALSIt97BsEhKT42HlG11WbrUnYCOJ
WrXPNs4LI0B6bmd/oi0wAyCBplik3rW7hAGmkcJ7OildYaYqkMUb5Nyl7fNHNHetCJrHQlgy7F4i
KMV+613h15wM+e9SLJYnrRb76yJ+gvYqgz+uVdEjk4ahV5pteeK2Lzx2uTa5IzxAcQOy8cvXSb1D
jCEe1QkO3xxh/XBKkJyvBbrQm69yCQfBl1zNxLHXMNHNfkA+vA9oqdvkIJrR57wHkYH3rVLlu8sD
kpjtYCHtqjR7jrvKwr4xzQP0/K7E4hX6D0YxjrcqVEDVnHnLUyc/2aDn+KwGiq8i+9/PjfVfJPav
cMwjIIFvZ2t28gNVKZegULpdkevNMEo2JetQK4dUD0+DiVn8IuIylZ6RUKWWNhaCw3PktCl0tULn
bxMB6pa9tO2JMkK38Ph1ERjP5Nwhx4HUtXcEb7gCxjF2RKMPtWWK0Yaqh8uymKa/RqP0q7IVVDd4
RsmFKSF5GJonrB2rG/uwJlxRyKHYjRVxqwtgFbsbT3ysVQP1PkxovZ/t/VwayzRmS/pdZNm86MEI
TFlfRDywjZF0uNnZBy8Waw7pXKEM2ovchgYnNbBNAdVbpPnr7ZEoaeeJrMB3pGNEvItB0aNvK2qL
s5fPvNebbs22RA5GCVgzfe4b2o6v645U7zE0UeqHPSiFD45Ov0vCmEoaSovSZK65xpl1TWoPn1kn
KYjHJ5xIx5ZdXGPLXb9p2BehG1uHEjc/xJNbCDmE+jLul+Vp56mto7v21CqJXFUHBe+PStsaVqKS
x3OcaeHWZmbsKumMcEwR0zIPWnOCM8+dy4NYpSJXmi+fmF3wCGr4CPV9rzg4udWN/23PIMH3DrSL
zeM3i5z6L4PdqX/Q/i4g+mTYGqz8LXj7B/CvA4Xo/wP30FJOUV6uf6vD7ePNa55Tvakx+/lvH5A0
tOHRVnPaGnPGpfFd2unXCZ7YIj7FJaexCIpCBZ2mYSHn+dORvgvdEBhuYebs2joyXH1fxqwcUbbr
h800oI+FThMvi32YHD/RY7M43vnju8tvbAyxv63NjP7DfNVVw9FPLyXh8HO60Eh/woNEAMa6kLoT
wcqcOVB6M01hUupnROGbcwB+zEScEmqliY/pamb7M1z7gLz2qJNR/T9gzaxlSpAzMND8GcUd8hkm
s7ry4bXqqtMmXI2oLPognJ1pmUMR8VX2RlPjSicWZJm397J5z5fSjG7oDinYSz5/NMQ0PIuVvS+9
OrHzX9ET0rGSWsTn4z9B03Xzbs8gi5bW5soHuI8zBmTaklaE2aDib42tEoMScnXR9GNXeSDjohBw
heVltn3QyxS93TfolXdmT8GUS1m8CAcQqeyx59j2+F4eUDqpa6mOzn7SsolkGNWhD521uANhokRJ
xvsJFCdkafMEU4S92oFOTW6fvOpSVjwpUjb5/hy2e6mRtAYL40tsgUw8Ou7KQkPqNG5MsQKKcDZj
+nNCCmSmLDAeZ+K1XDGglFFoO+Ok1cZ//rjzZ17gf/qYKgnAUgFwwp1qfxgd6ftCRdAGZ0UG37xL
h71R7PfzhmhDih/fF6j7Whx1GGCI8qUcubUmhvYui61QvtuHt2Iqp1XetWJbzR83WXpzPl3pj4zd
wf5zHDao6hMKf6xyTd7qYJ1tjbXa9eJw7F2w/KqXEH1H//FLV9fnxDvyXLOK99bqe04iuiFAl1GP
DwovX1JxW9DirLIMKFE/SFZK92ZsiFLU3E+A5fu/NS7wftWwJPMRPqPVF7SGFi01sRcW8hDncL7g
CsYYUygqB9IacxQ3mB8Cbqpir/h7g4FzaTJwHQu2RzpTuWJ9QhZHdTVuRX+d1ad+w7lnEtXlvdlp
WrqR68IDr32JlP5CxNFQehxkphG3tnRFn4EkJkq/aaYwUXjtLFSN+aIUBg1OPPksn+Q2EAeDPpry
C8j+tbRzKOgruyhdUGIHMX2yRVfN0/L3GYfpAwBo02r3grVmWhaou8uAFFai80cVMf7RZLgrpCAq
eZk/u97jLLKNULDujwWLCGib67vUCxqPlHJA1dhGJ3HLHWqQskOzDZukrFUwhxRG9Yy4HVr/Tkbv
W2ARzRZjOmX+QNb9kwtbI0Zn2ZaLEQFXDAYJ9TmgJQJVvz8MyZ26UTwD8reFHWDjG8iB6Af5hKly
VoGdBCYMdO+7PlUt9mHbqvhZdTpHRd9VTuR0WyXmgkgghRq4i7/RGvkLGOoEL5UmWOuPPiJKlr5G
OsYSNddW8eUTyNduCAEB5HZNSb7aiHIqqeqjEhIneuVL58j6vLSQivUkAYxg/vCUzsHpr14LWABo
NibUWxirijv6RPUbO5Cvq5OqVd4DAiGhE68Tz4mDt+OPCUXNXxUK3AfYbzG7/S/E+v5WzUJXpKwA
0FsYqu2y3cOB1AiLXmtlf9dyQuMmwHK5rVkocoEQGkLTHhdVSgaDuj3VmU6p/QTWcex/PqrSrxKC
OYYZn/qN9PQrZxaFTO66nMWEuRnp53V2NIxExhIq3ZRAuqD2ZVdYCSF33o9xR5pGnjOpLs3/soJm
vPNJeuejiCbNMWSb3aAvkR9Kj+kkr0ACWSO6ia/pv3/HH5nTYH67jG9c5eKUBn7/DIY1AOx/6GhC
MV9zc4z+j5wU6n89uSkZ2iDVMLD3hAoM89MqJ9a12H42PN7dS53nJO3oHR7hY9+Sicij4Mb8SvGz
CtZbs4MEEMjr3PSk8ClVgnGyR6tq+GlyrcfKJirXNrhCFk4TDkOWy4BEYsQtYFQcYyY3iLKPqvS8
P+yRNmYATlB8nwweNaxvu8meDGnjtkhbRZqgAkKAwspNaC9wkFxiv178meDPA5TumZ3loGQBVJZR
pQK80Bb7w6rnvnygUdsbd1+epvV7woLITrq+Lrkup5QNYMc7oWzoBYU8TFmrhhcy/V5dR3EOUJFU
FGuGXRDTKAkhSc+zrFUXNuf5UGue3PmEoQbnrFDlGLR+S2CgbTrcKxUK8C6e2uizRx1aJzvwMiqN
EH/LgaUozOuZS50ejqrHKbWaUBZMWRkfO+c85BzQwdq0FW7aPeGcPZU+4tpaBKegP627cKrRE4lv
f5gvtygScOmsXm5zVNS+kHG9AgAf3xpnWidqN20+wRCT9UtMcCZ8SzMOrfQaon7NYZnyiYtrsYk2
xN5+LnUqUHalwcSgU903JQb0ZtYXeoy16Qo4U7ubNf08CpZ8Jo4Vzm1Pn4sZAsnWb/sn2RiTXIBg
GCh0hYb3I7s1iAHCOPPPuRzRMs87WqHMUvag2coI0553EaEUsum+zZRKieOgVX70BtpC+gWxdSQd
3VrTdLlcHsP2qbiwuR3ybqtxjXuqjDAvVHhm6RLf0ImBabrHvQmhAdfZSHC37eskAJaU6nFPkNLT
c/Hi8GvqUbs6w79vifWa9uGYQcG/3sNfSXf5UDOBDGL0mOWt4C69+lQFjAb/gH8NC4s6JNbxwOpT
SVrzgHOfvbLCTO3mM/KYj6AY+m2q7guyvx7pEA5vY9oGS6XIK30SDHxYdw6vWIOCHiPhf1qAUYkv
DZOVO9s3xOIC4kScxL2DBdEf+GYwPK1T+qqDj12Csivc8rDgKi31DLKYoHoYm68s4l6FvbUDAMZh
qrgzFXRUjVv232HHebUtHpoVwjeDLZUphpHIM/JLc8vMO6I+E5UM0Mz3PxHhtLaTAbH6bYOh6mdu
HmzuSnY5S41dfMObpXOeX7y5m20Npfv2YScMJLDQoq4ggJLYHWpes1cGJe0nMiHRxs7O4Opb3NnT
RiqlYKvwnkWF+usWzGMM1F6UcLZt9BXK3U5EHgyNoXu4q96Nw0SzvhoPDLpIsdGMKD3+s4/OaGYl
oNyIlkVCmlmLUN14KjF6KXDAOaIkuTlWDLFz8HkGXF9NYsZqi5x5s10d9sQ964dv2X51lrYo/U8E
cToNhBOMdO4cOlSpLtYqFC22csfc57U67ofq4NgGMSQ9CdwYas994pmeVrDqFpMKPonAkrz08lFK
9OZFFWeFJs4cbl86jJlnjmsQP9HxfnI3KNKaSHWYJFjK6KurPdIJ9VAiIJNc99QRYZf2agfS7nKp
/mZM3iONqlZhVHCWonLE8/UlxQifWUh5djwoGZkCSIruClTK4PazwNXLdLZWmFBKTckjx+n1Iw5v
bmgJH6NORESYZIgwgiwhlNoA+VfCN5GThUf7bs2qsMUslC7RXErhL7COlIH5T01fTGaNGbiYG/g1
/FnqR3y3nDiYTFOmzMedmxkkBAGN7RDFlbc9N5tzB//euyOBunKVDI9mg9r5uCyqe8EgdGC6C83h
obLcYXw0P52L9E2FksBRIOwo4JwLqSzVw71f8demisiPZp/j5zRqjj3DpwhloFT95eDHExqxGTWV
isaUcJo3Wi0122CRL/MQilYjewNtPMkKxwAn1VJHjrXMfBj2urz9Jyqz1YXclV1rEoXpbfjlpzLl
ip4ZDhvIw9QcuPEuT66a/o5vB2H9+IWkZTEEzPB7ODOOpLvT6UJgSEvsH8PVaXG9abzCE8uzzaLN
5WQx//FUKYY8hv9DNjthip7Zmyla76KWi0uOlg4qXixhpiyEnTJc+JHMrcbLtvxnToN4QI79KOA2
HXxU0PnUzDY/E97peB88NtL0l6w+11YQHMYBD/uLvd61GEyU3u8Sds48Hcg1SIl+EZF9DlS1lQOk
nBBYOYpyX9xo+eXIqi2zqwnxHv9Sc5OWcjjtdjMwIOy+uOhH2+yXkqqpiohgyHvpjD4zi6ePunZe
XpHv0Bm2rNfguwZUKvH/a1NkK7D30c0sbm8+oO7RT/UnnrouNIkuqEA8ectPQ3kB+dlK7Xz5wp44
uFkDkhcADAwdBdgP3th+A8MPc+yM46XzdScKwh/wqrjnf2vQmaCW8r1e494Vb4te7AEgDFwyPdSI
f3fPpE8VfiSdfwWRYxETw7E9W5m191nGwDm/2ez7A9EZl0D9Aq82F3Z3ww1WNyMaPSr2V+tahF2y
50xnHnwH5A7fvyjk2S7nUvRPZGTquGf1v9XSqCdUSaQc5gk2ciGR3xKQn3fhzYQmDdTpm8Gtv0XT
7v0COmmhtILtvIxo48FzkoOKfFg3m+SOELkfo4EvbKdHnQznDL+rP5Zko4HVQqpADQtUQx6w1GwZ
N4ICpLyQstiZff2RuxkjBU+YR1+Kgr4VVlUu6LXma31Y3ibaCQ+a0FteGjecdRGI8822D+81ryLe
u6f6KxulPBnqTlMJQaXSzpAdXc+WN7gWr8VQ+h4kyKIYdC6cQHkX8IzdhEkrU8imO1ai4EVdGXJs
OoK065Vgca3LQXGkvF0SwuTE3DEC/TlRrOsR9DX/vld75CH6nn9VVbwB8l5aV8z9Pd7+TjYVKHc8
45HuWwU/2slKBiSvbiP4W0jxKE3NRYKbsU6meCM+XTy7/bEF4Noc0J3AfB2Do499e888tXAUyc+S
re83SUx+f1gU7QLX+sKmmfgd3zJf5PQymQX051AKiQ7TlZIvzDY9vEfNOKTN9GnHRt4ykOlzaxmw
ESjzRSReV0PalwagqaHKZyWFCkkGLSK2Ms2hsinAvLdOItLminNgnZv4YrIMHYu2XV4Hhp1e7Ze3
aXL2DJP6KvxI1TWY50lHB4GRale+ji4zj0C0paohTgMNe4So1Y+1Gm5u4kbNcAmLnq7bZw3RvV5i
QED/Q36/7qt1WqDcVGlZAvdIJ02cpzZUv+fJn6oESzuVAItm79dktgTkj2Yb0f2m8WBjrXXngnzn
lEJjKZkEclWPNjvKjnhQLwuktzBoHGAXBsCJpgHg+xmh3Ls2sOaXv6e8QK5LfgX9Jv0aS7eqiihP
3O9jiLDLhXL4ox1g69VBlJso0/BUGX99bfZ2lGEY/D7qojBu3dP4MhGa/nZcD9T9WWVsTvQL3RWO
svLNPtki0sS+LW/jJFj/F+EPe2wewQq4GfgZIDGJ+Z1RignV0E+NtTzdPuzNcfqnlU3SXr21lR8H
eCAcP1QGvyM80K0aVJ+Ec4cOt7MPWoK5LEpQTFfB5e/seamkXvHw+QnGw4T1Yqg1k95JkZLX4H/p
ZK4PVmrHsMjO8CebNWZToa2RXqEkuTyr7o351QGZxNYgbjClMNfz96yYD/tyv6fKcJ6omLTco7zA
Mstzc+zuyi2u6SqYqxlgpoU8Fouo28nJEQIH1JPxdrjHEimkUIesrrh4E+m36ZU01YSfgF2NYybv
MQWSddcgPjAE58cgNcbu/VU9JLp4F5Qqfv9NMt9m2Y3FfeJJLTh/cQs3SIL5Lpeh0VLR3jIz9v/8
Z9rcE/NC6OhxW5txnmdYTrx+PE2kEzWktAuF69LgE65zaNYBBhzug+nYdMM3cuY0QfvuKZwryz2P
e2kQv/2M4Du5yklZj2zu9u2MVZtXntdzCnUHD1YViOSJvdeWNtGCMIxEwJLzG3XoAvUNufeSWM87
r9zqShazje+mGpKTBoU4hxjZedZLkHnfFG2VXk4TzFVCuS0kmqWzpkoETwKfnPE+M7TQxRvMNIPt
fMCtT1oeZmZU1nUWe0Htuz0zbuEa7q05pvm3WI0rVYu7icE0fOxD+kWe3UI9hlgUaDnC6p0pvNej
HB+4w+8z/LDlv6nooO7Ran59dK62kgrokl7IXHz/Jg2ICs1obmWOTDwxpn+Qz7gw1a8GmlicFCMb
XvKdcfndTJj/yIj52PEcJUhr5iaNLODyQVDxZnFppgyA+hkf9aRkiOsIND3SHw+9bmUF8GUNPb6s
xpsiVPcoQmx2Who9bar+leaJSQWMSFH8/31/O9p6XGaRjgBmHI5mYGW0h5foS+Z4QvkcCqixhkaA
Gr9XCl1aO2aDC6SXfQlB25vD80DmTh/IKhdRyjG30UBRo6DTzweJBaIkg4rtpk1bFPKoB90c6i7B
mChJgb2oRv6ENubh/Y7TwBazL1HZ7Hkg8QhgUcFPnzAa29Pu486zfpzpEBMOU/kBzsr2e9jloPxr
QlZ1FnsnKm19SI2YPCqAhCZ0Aoi/ay1v6hPi7ue33/b+2Az3x2/iHzUYEiUn9drpO8BfmDEFawVB
LWGaoZC8ZtjhT+/Xg5S5+s/iutjNiKne6cfKNLiv17v5+Pn98+Zg64GwBc5DYKWyZSeCSKRQgccr
0T+I2gOD9lmlzmcfs3bgp5ge1BSWQZb8tJhJf2xVpIYph4bsA0Rpn08ydBRYGsnjSmkltc9mgJRl
LEeFr7POny8dNsu2bBR9WenqEZIrn9GAAjib1SQAc1o6oS2Z7C5qHLeXi+V0QR+uVWkVQVA/U2oP
6WjlrmEnazxjs8OsLQlDJ38MPFADYwwI2iQpQZPlCIN6NbBKDpLGQY2CvkTCsOYPgIgnaQpv4xC+
2zJ51ZtAwq+xzmDq1USeWTuB+7g+zfmKDCfk8b3NcUAGmf5xmUNO09eXjSd6OL+MAj1NLKBWvKR7
O/wHrlyNFACV85PHrFAJz3J4+0fxezlnj5V1Ebah0gI40kPtT4T/xptcJCfIc0lt/6f6ZVNl6kf7
leHA5g2YDiBtlPZi7HHn6u/gwGB/wrAmWjHH2Qq48lKBGGoGHo9XHW+yk3Hz5N+6sfqKeBceSjSd
Av4OQqZznd97blRlK0+YWkI2MSQfIw2zxZ89IbV2WhYGGC/9Kpv9OOZ46MeWtprkGOvBk6ZGCPXm
9CC1anJPdT6THhYiXl6zWNn2FeUPnXjcmAmGfA65+EME8F+UoIUGE08GLlap7z73Su7sQqb27/Bi
EjFYt7e4EmL6v5z+0ZYyqSjSMqWNXW7fE5mBCIrMMUwd2ZxdVLLDGPaF/VfaDpDmj16v2m2c4blo
zKhUZKL76uUrprjrVPtf0/OXU+vY/nHDRzc9PvbcCOBvegFTvh/9BNGoHaXofPg0auYpfqMNxRM3
LNV7W43rglWZxhJizcf9Jhu5cE5VXy3V40nE++SizWR5vI5KIxoOhVp9ydZ+jlu9XxvoGanDk3u2
rAmZWg6GM6bz2UoqI/PxB6O62JTnbifpKFSYPDsEsbWTMzWXmNi+tEKRtpH1EDaEER+hNGtELr/u
4SSeCnGWLaBtPtwGOOT2PxEi2g5LhJ1QO1EZd7h2HvWd/rzuM02iQxHJuUoQl+VqPLcqVzEZxNeW
2Ej+ll63qJLnV0Lxnl1XuboLOWoX89pHAOl1FouyPer1d7ihBdxgaq1Zn3Gsf7/fGyKgLns0f6Ac
b/+WBhIhEzyvd4sf8DZ6+uk7jlTHC5lJeGsveyk76eqjpquIDwrNDaXe3/kEnq8RmEMVxGnshVO2
zDbPo1FUogvNcHs8PFKlk4MSUuVWIIwsBpi5Ut8KNMXn6NVKlvhqRaOLeAa3lakkj2SvTRCe1vkA
NGs8vhMSr7A0z6QwQIjmjVRRO0QvKHFkyNNV9Bkm4nj3//iay3EVdmcgWwte4uAAr3KAvMem2eh+
TDH2BPKhMoQO79B6rjaxMUrCNEV7QDvjDqC7dG8QbeATI1Xg3/ONQU7PWU/8NGhDcYpBsFco2/RU
TgCOSSEubOuMtGqNFJMJbbFeyAV80Dwut8876ShlxbMRrlZuX7RmpHOhYsuzXpvsw/zuNEDI/n4q
BNm3GkqjvwLzcydoLDTM6LGCyRyU///2q8GDrAuVylcxXXsXDXz2oeQlxP/8Yi9OXLLAkansCd1x
jF2v2/+TW0uNP4BpI9OBzg+Q1F8YRwQVvkGI4mZwRhJV5OaMJeJwBUjxLfn4Oqdk09rlXjlQ+WIV
Y43OhNi6u5Lh1WhSF5MgNUsPh3qVDcK/QUgva6Zmzdk5T/F3M4CHG6YrLKDUnmBSfh3UkPVvruTL
qY55DRbcR7vDT3N9O5QLr7NfwlynsVmIXBVKpz/d1y2lqbhKk5/uxOg9zM8vnxPd4X5R+rX/AyY7
pnyfnN25YgZW4uGEfwbbB5SlqlfIUjroN+XGjddUGjDJjIuYqKwNa4LOcG8aOJKB+eNmkjNkWagM
SetSMx+/2BqQ6M2l/ZnP1Z3WdlScj5AKCzi/MRD5d2x2rQT8LKTxza3XJg6KuqoW8ocRPmVRx9Sm
435U128M0cMxX432tApg6h9jvBLuuBA7WEF0Ze/XL0ZqzASk7Zm8EtU+cZvJIgv17ZIEQ/7pl3pi
F7m5UiUOjIzOLxcEXkKwSsv6RJSMMI0gzMq2IpDOZZlOj678eLHYvQ93YUm9o/tVeQPds7aWJVWR
L2wJuyOBrt1QXYxZJCy4U6Yv8hQBsgr7qjwt623nydecvBc+Rylf0GKVnWTJb6aA1c8z2jBZjaDc
/oP8bFbkiLkDJ3yzvO5WliVn6XTfZ/PD6Iu0jL2/vMxrTDLlYzNMlkeFHJ6IFIlpRx6dRCpqOjm4
pui5+1/3MIpujz7e899HTeTDxD2WI7WidgC7rxW3Df0mMEEjBju6EMehVIGMMQgrfGf06EHEU7p+
QBjVGf8e4r4ELcq8yCABqxAnCw1p09ayTg7bezMj73q2Zzkl2S5DHBwFb5YGJclSeYZCUC8pYiVS
0Ae0B7xz+W2weJMUdUY/cVlLjBTEx/7gUk1gM3pygQ4U6cmFkfMBhAE2o6EsgSRaqkU92f2FK0Ma
nuI+SXsOp9CzVdlFrbx2N5iZWGZjBH7rMs6lZopAaLa++ywSwVOVBmQ3wpn0OOi4SdceaUxW/wQU
hi5BK/UFj8JHAaoLAUFwLm3sPnrWRwWpQPt+SwZgZ7rvD6IaYtjt+xJHd/AEeLluHIVrZrAT4Fl0
96LJG/zBP+0P1qMb8ieDBYjMvhBDCTX/u9xenAbw574L3std667d77Jp3DBLxKHGyh3+bfqA23zw
c6Vd+vcQdhguI0iAuWsAa0THFtyNdp5kPlV9jCrK1aXBLD1fINfm505PQoagF1PJ+pcuvssxQaIw
MHxDZMylxyhKpHcRBigDVqvik/7cFVcY3OG6MXBlq7wkOw7w2YFmU/Xzlrws42B21jRZcfUNxqEQ
RDeIDky0g5cp0M5wATDB3QLJ+SGKEdOiYkhNgzTtZ1qx05gWhlJjg/rWvd+qPpH5NsJrILhEFbVA
4kjwZGp1shNTx+BNs+B2a+2hrCVosDUhd9QGipFrVNyK/gKSpS0tlJJAySM7n86bV1ReyRe4jzHv
eFDZPZvWkKU6ObrJHLxiLs1c+QZvcqWKsk0u31Ojdgz879OP98wPaK/B4GSRBRHsEEk7XUc6Ftuw
D4TAJIDahLS4F1J4Xva5bSi8xrkpeu5xQoVL9QO+wumXbK5o3HwmFJW2lx3MDUGgrdL6EikBFbOW
aWUcLB5w0zK1bzT5gePS04bUOlw8HmJvWFwGpf/5FdusYEMr8EwTJp3mWTpZsFFcUKC92SLW3+VL
B9HkkugpzA27PnbazCi5GAAsKLl9D+fi+/WcbHaXv2es74xRHTJxS8CHa3DO/ZDtndDEhnNLdQ0Y
YcV2bgKMKY/wb5ez/FbCYKjT7A0tLV7ZKNQorBV+RjoQ+O8u2z55mmWL9AQ7c4PfNWJQom/rKz/5
ey6qKOumOvWhlAk1hg5zaWpyDJdDemRuZcw2Vi+jKtb9lV0CeWtudXb4QJfUn12Fyn16B8TFMQ5N
LjOFUSrHQIHde3eArAdG5/NOduQZBwSgA0XTJ7Dh+GcFLiS6u3YAxWW+sFRUM1mOPeZZ95pwho2z
2CKADJZKEszz5HwgBQrGa+75WcoRDic8uy/8/TECk8DhsQbzZDOXoONuKKT4rwumd7+N7pvi5Byq
pCvDXMQFJeOHMhWvwOwKFXTsXG6MlxqAmf4bt+WDiYap582KwXx0IgkUIcuuX2NIMJgWknkPt5bk
DKgoDJ4mVgMjNPgJI7CNVeR2f99ZgUIPGY32zeida6Cq35w57+r70J3vUHkdhjbibckTj3JWetva
DjJhx2sT0SbVUvJNITW6MTGYfLHeyhuzF1TK7ZyaM2gBpbdEYzFMsHPpMwVX+tMeaYeCkFt0f4nu
eAnCyGdhJO29MUeTAtaWxgSaLSXm/sSpfvbcjFKNzCQ2XmbVT2sYPH1xDYI/FKERs4WJowLK7sV5
ybdwE+oaVatym4ajjQuDRgoHnJxR1HvLNpYnya4DbfUu33WG2g6OjtYmIh+C6ExPbE2XG03e+IPE
XgWIPGUPBi+Ev8D+izWBVTvTTUHh+tFpk+Jud3yy5bYfOVT4Peu4qURF9JRhDGGjN9uxy6Mao7yW
ehQ/uiJjW3wmUYVg5UaAMSwmV0EpkscPCm5/7xiI64kYPoQlXiZl56xB53Se2r+GI4/8/kN53CdY
jFmzwCe7l5ZlTEuOLhXyVu9avsr2swTtyDStNVNN44JpxlykpaxrMI6eCx/DjTmKgqnZBx26yrBt
C8ky/tn//5D95SCc5AHgHf+0izIvautKFdjqTW5AI3n3U6cbKn1dWWWBAQLSxZ35V/J6VSVaLakB
BeW42QCWY9DN4QHlzS+5FWgRmzYrsBC8KzaEo5A6u8A44cVhaSKjeD265jhiRaYeF46ODZGW0Yhv
hsqv1CR8cW6ilm/V2jPisrQoc/99SGkwe4Ps7PqWie5fU/FkBmOckwjMZEX1c/AYnoIF5amJbsOh
efbSPQhAm9/MAqz9crMETGzcLlHjZhuHfCB873y95yrZat+Gx3O+5V4qjhNoJ99FMOZoeukVEyL2
nsHnWxDTvvC0e4x4UQpEYzzaf0VA3RVhb1KJ5bSAigdDUOb3MRCtgulGhQsQkglJUggkBOG40nnW
iFaBGkVaJgHu7my64JCgoySUttWkEBJbQ2wdnSI+dKwm+qv8xZEv9OO2pE72iQi+E6M3qYCrSbld
tJfyb3KSMLFo56TMlT9gUO7kEmZ6pgmoMhboPWf7nVZ1RhRGTw2JFejZYY6PI8MBZWDj0pIHvbY/
ptBilP+f5J3izLpkAC2wPiSDIxYMlRpuydU2voiqp/hKZZLqqje2VR2C+HOKLHq8Hn4YvgmQOy/x
LToGCUN+M5AaKFlZMMKUCWOWHzU49jL1G5yJ4jYAWr1VySj8I953edC8wwVnJZLjaysn+wfQy/Eb
hro62QT62ykAbYazLVfenqGtd37sIqmPbpoZUqaJIRV7XNckJI0pqWHH1UJFUcDXVD8b9IJtqgZ3
XOvY7qfWY9awE78QezsB8uDhHCNvYm3rJKTfYWrChnVZdSDvvQcR1nafFw4xqOl9zqA8zW0Ildil
mmQlZl6qKv/qKRkZVFeIVOUrSnqG0+3nRy/jwr3MvxET28BL2/BifOJ3i1evv0h1ROsVUKmFJr5L
dZ1RXnE0jtHMdmoOEdES+4XD71mpedkhSU9V/73ctrvIAUNQol9w+Y6Y3n9ePPL9GEiLLs9wExbb
zz2uc42DlL6hcLpRVmW1rvlEO1sUn+cylShM316hbzJq8/YRNWN2hgiz48XgSIVR16qAFOVdR4Xq
uehyrWe9lD0mnviVgLpuugwu7EXCYlTORyFUCBfJSq53auVwinYtpRgOgGOFkKpdTvgI3rSVAC5T
ZAGFri1C0GokqOMxs+t3LW4h+dvzJpjZCMTtdOiTQ9sPzaspakVHbQZvkSfKtrVe+W66ZixO7pSb
qSSiWLZu4kQtdWjrpRaURYQ2VWHdri6bt5QvbiPLbVyIiLDEjsXEhDJmZTgrC4TD3GRgp3Te/Eyv
1cibYVnHsPpgnmYeTjoEagH3AiTu9v25Z+fxp88cB9jhndL+MeUpVPa1lGKnJ/2Mf3inb7eZq4dB
XuNSiLZ5SipA+Niqi/yja4oewkvV9iDwz3SuGCha8DXO7zUL8V7P7pO3PSfgJ80gsMf4D9oKoSuX
kZoKuBpPafnG+cFZ9gsAdn2OO5M5cZ+GPcweS9FNmN2lk3P4+/YgDIQIB2heiY0fCFhu3x4y3n6m
XOKiUGgW7/o9dZox0O4DQgfC5PXzy3lfxGhVsNPSRqlTwAofHbH8NeewOAdUWaN9p6jVo2OJHKHd
qw4B6D9FMIOH+veIMXo9KAaXXZ0nB7EpGgfmesn0s1aqJNTHtdx6XJkWkmo2PlmHmK4BX2naqqsg
AxO49Tk4tMYq94dAOdbVdGo07LIWiNaCMFKTtejLNaK77omwoirPCR/K67LlA/Ldgu1xMis8Y4KN
xGIKHvMhBxbi1kMQIJzbZUzoQVRcIdYADMQ9Yat3rXl616KRrx0PaRjFiXpoXOkbb4uSBcL0P1jv
LiRFIQNUqab2PZvlLaAixZtXnPV6cNV+JSSTeUarDPmjOy/gd/o4P/jKLaWntQ/g0g7i7uKZfnvh
rvhsO2XRLPWcHnzQrJEGhrIiN11HHg+MdtPgKxU5QKpCVgjMff0aRlNCTtU2MFzW0jmUi7N8bw/X
hYV7tisjIIIJUJH4W2pzMvNywVLkdKMR2cy/OlMJfhO7uhXXoRMOHHP/5L92XNT9Ns44c6csoCxx
YJncQ9c9Fec6ch5r1JZ6JWK6jP+5ZF2FAkrE1t2GtBImdRZMbDUTlIoqq+Y/MkObdHZPndQYKQEC
hlVYEKKMEXbqZdAIsulHt4hrt4IO01GALAfTs2NUQEadqACvkh91Yge0RGgjgZn7uH55XDI/mO6Z
t9+KhmEkcPeTN9SLOQRIZQZ8p+m0PWYixAVnEtIoX2K+o+EpABKSqZzr81/F0/JRQPOeUwL52+kl
y++PtvGC+XfAYZr/mUFRFJ0OVQ7t6c4SI4TjZNt8SPf8RgEFNeDDLV7nikY5bLuY2KYaBVkS+Hof
LUNgwp5lreC3olAB+kVp31gGXk4cZJrYudkNn46+O1n1NUc3wHJyT5XpSIpwguNBWInGYojcwDQz
Q4oTtvizEeJbENCM+UYqP4iIxfvLOQwffM/mPBA0VvCNJp2FZ3F+Sqx5GSrRDZHv/PYKTxGNxLOQ
f5epU0L89zcO4Ni/4+lD/pxAKmOaTU2VK+Fn9/OUasQNTTB8mdpI3Cofr9ezl+HjwTQvPIUjkd05
2V62rYREpCid2yN2aNXgc2Y8DlojYzJQzyYOWmEybdYDCiDde8FmVml5HovWG9Eys9/Z1H47hKmQ
D01LhCBbX+cbKH10PwKxvJfZb2ZgJ543eWZDbbZ1vJzRSUD+eiAz6a+tUjoPR1tUXqMb1zJ3TQJp
s+Oxhu+dHS37yW9MjA0yRQdSYSvc2jK/5kB+hvz6xfH6DVjx9cm0i8Df5Vmo9s+QmUGaMF3Vup+q
fjFd8YVYtXN815RvrE9GNlMOsGkcU3sE1ugBCCs3jjQDKlAt0Pc57uU4XYDuXAbvgIUxmrGH56Fp
9DoiRgJlf8qmssTOMyalFdnHcCiG087FiH5oo+F5csbYD5QeUR4KCyqbEy+ZvG6YDojqLEG1wgTG
oEtClqJiQ/7uygAvrckIldbgQlPq9UgPA7o5M34W+XZsbO/HxutlqIuyNxQ5NKmc/2HHhDzmHH2J
CpBbe7rt6RFPjqeVHzARA75hyllfOAHk67QzmaQ66xwu0iPsRWatUdZ+4Iy+YdJNEIMjdPSeG2Di
gnnP2fmsBfFHm1tCdfM2rPJ3NKI+b83wESrxOSJAeB0jB0HDnL0PLZGjI8w2jFV7/EWABgjw+8UT
afkTTX5jwy35s0fQwx9bCgGztvQkyHPfIG02ZXeJmInk9Gh6f/oCDFO58rT+lECSFxZgd5e7zEme
KhcMxsosld0hgJXBLYjcohm5BNJTnFtpGdH5tOXdmFZDkwW9PqzyWxitHDFR79rwFx6Xa1AyZIk7
JbjZDimumb/QIq40Fr16tA3hr2Nq/pUvWyTzLwF1FywhcxGUYa+JwOUFHhcUtxYQPMFN/9UT5VLK
ycc/j9fzbD9PtK78aFiX2uuO5jaRQnsp0o/Xba+1IYgX7yYHoOfj9I4EfN+od/yJdKBLraJGczU8
oenfI/NtaPDAmY4wbMAidRNn4WcDSrZY/6PD6e/FeGBXqPCMShahLWINlsnQrbJdbeqZQ61krHog
6kgg+22zTSXzcC0Pd68chNaPy7bv+K+rGBdNXodiIv4NV2G/X6+HqFlzB4n7o6Eu8Zq7coj7HvMa
5VhcxWZaU81Mw6Ji3cs33TeDWkLzfmh/1YzDbJ4qwgkEfWzxZ1cAKWVTbaq/Bm3tdZRXEMt9GYHz
I+EK7wuzhl8k6IWZe650gkSNHc7v23Lyw2kocKMuDv7xn4EQdv4v8E55zSNbXdua/JxKWPAnK9yD
25eyB6R1F82qU5vhpUOiS7dhIUktHu25ChUUJLszPVYbEXf8IDx6FPfzUD4xXx7m1utSSFAZAwz+
2PcbnzRaahmKOxIz2zcP1Bu/YNRlERPJjjoz20Chi6lEWVaVsGqY//2p75DgQmjyCvrAlVNoeMvk
umL+t2rQoxumSrv+aReKEfueXvwoQk3qBKEoAfEV9r/wrNdlL6zyfZhWBbyUGxA56SXtuPNS+gtE
Xxc0WGCAZsu7Pm7QLiKM8B9t4H8LviRJ+arBlVrxPejmKPMmKJsxIepwSXSlrjkQBUvBwEL7/8Ym
nY3iBq/dv8eloV/z9hKOxgL+zf/wtgjrWwlt0vcOaKLwVYMCVs6gMk8Im7TXZokc+5Bc7eq6kGZ1
Lbh2rKNfVyxcIvy5hWQaI7Y++2QCGFBhx8eH+rogoM1LWO2rHupROPxaBDX5+nGg+c5f7BY6xWnT
5qzHn25+R4p0eJMUP98ghbmXvMhTpPK2iZpZaxzjh8fwBWD9Uc3F1ztQWy+yUfy2/sgg1AJGynTE
52phcZTr1Bw3zBIy8M/jUj64ypvVL4AbQLQyG6fy25MFhr1jRptrxXI3BiEmlsPn2IL+zdKMZaw8
bCL2kl8YA85eAhPpYyWbN48XFFHjNf/+yRwcoxT2jqBV+QHYNwfPZoK58pGyFFq4wLEsr64rWV7z
hcajeSb69VFhxRpRPikK4YO9UNr8ltPrgA/7Gx3SeK9Nir8ekkoMl6VMFuc/YaWhxWoKyQihjv3y
XZTMlRqzUgnoIeHcvuWT1S5BaCYYZNiQPEdm7HEPXVBH5Ge+cU4lzX20bRxMcAtIPjctohy51N+1
nYyaSxXuEQqMDksY4fmPSC/jNTXZG/iyyORj/p8op5mCJv0xTNtK4p1mPkb4UDIc/G6i3WWVs2rQ
QynMbg2egLv8aZnp8H8+ZymoCjJjIL/qEjpvcyfpBaBl8sT4wUXDgHDqdnNEyyLlRll28ACC4BYA
KpsNlSQv40W9m4tVZZAbyafJwRlcfhlkpWx+7w69O4qCMWK9qZnvjXHckO6ztJuHmM2PSerDGF0i
nsv2TMC6ZbcegOgagNacSJp7FqBGUKPuPScKUKg7i7Lt9XYxKb3l7wxxv23SBs56RCDGNeYnHpQ+
whBNI4sQek2clng4EsgXF9BjQ4qpdSmPaHuP5/OIM0H6hPVhG7H7c7lWCCW6e5h1LC4fKL+6SBI6
jFKrkIsd/bcSInmQ5K2HH7ECz0VagBVsLnN8LbHGt2jWINVBiQd2q+BdSZDDgYgPy1t4fPtSMdks
N6JkUO1uC8ey4N2l4Bh99sWS0R0UYgH0Da+tLf8GDDaTOEoKQcXPOc7WI8VdLRI2iZ3ui5w4NU5Q
fGvwzu8Jbc/G0jZWmTT9PkKkXNQZPVe/nqhtuytrlxqQ1HG26SEkXEFD7niGnOrof0IWVnqAclKd
nVRwzELUNKh2nI6zMfIbLkJzdf8lPGKMstMR8+eIzAjhEL3lcfhImai0Af1tc6XuVGWINdGfRTH2
PJ/o9p4hfZKYVZGtd1RRAvJvvrvUs6PEVBds3cZbcj+eCIBXkqP0CHuxJtcvOFhj7qa4rSHliv/s
+fHBIfMoHTk4uVU7HYD+o87RZTtNRaBG45DJGiKs0J6TudoMhyNWnfHu7qSEXS7xQFR38xuMo5NE
vHsyRXl4n/yIYUh9Eadrtp7MDLz0112czTvoaXz1nXS44MK3qMWiwLDKHNfiP1i82QBXtuikS42H
liViFhkxuVWQnZ9y6nr3lx4sCWNJtYO+G0fzpn4FJJmbYkbrqs/S34k5Kqic+/f1wUi3+lO8wT6s
RgmPpFRCCVfZt+eRWK0U1O/yEt9Dnh9ZuwyLhAqFidCCpqvTobUkB4alvMaHk2FNl8MRsVx7Vzd9
otYlxRSiQC/b1meeYSV7j3TgY5LS6tmkRqzrMR8YRH3/tdY8tTedGoWpDr1VQadcG7xDRvtRr/f4
v4JgUafSCgeho7ceEKeiwPDnf6JT5TK8jXg6qZA4agUSzjIk/TqI0gcrVnTB6oiwPC+4A0vbMnyr
XPDgQmIFgUDa/sfJFNCk5mtee8YzY2O2+W4TqVrQ3rhV5WIF3Hl9oPJFHieqyMO4S2I3VehLFPlb
xHPHQMBBrXFmmgk+kx3z8hBoWE+t8ScnS/FjVDwH0jIj5xE8vFwF0d6yJ9ow3SEpiX6EGFIcUERk
m8T37o9vlUvFP/sByxII6/PAKizH8HZSZh0mkCBKHEnQPExyNqiWBE9I5HX2CZ+JWCNieAgS989A
OcrbvKQdD4mdGPX9j5IZ7mEorVKl69GLXKNRdHwttej/xcE87mSRVxqEDTLLM4+xNuPPTG/ttxEf
E3tBziDJ1B7t6QaS/MDFr6S81pdeG/qw8IwJJon6NQoAwD3zgMGIWQkIpnTSmy6eOHx//h90TO7H
NJ8mtwq2aPJhVLl9xgQwnbEvZlKPadneb5qRYha1wE1GcqVoEJA3zoDkHm/Nu0Z4D1QYFc4vFmJA
LCJyx/mn+6ydI1fxVtwpGc5Nf28R0BM3CmkDeqtO1Pd1XKT+RqpyCeUV80q+RewmRzbg//EydjBq
7jWQjnjEjmFGA2krhZK8OAehTqaDhreJhY73LWO0zpH9koXFEsBu8xUvOB25jtfIHWw5RVTJ9OHj
RPjakHHsGtGQEzlsjqa1nI8EGoVLr/JKtqMnQwdhh+a/HpQ49rnL+MFJjnYpF2VvEycz4IQB69ti
PWfHn3RWeFZ/Qbev4xMReiOnahnc8UY8c+T1UC4DjTrgkzmxAeEhxr1POV+ocnTY5hrsKV49Rgte
bYj4xX9ZQrWzlRrZX4RKtgWmimtftqpx8VAGnDxe2vZ8nVms79ftWbWuer4CF9qJsu9atMmuwBNz
/QWS6tpVjZkkmR/Q/JprJz5IHbTG5Pu6FLHTX5sGktK74O+6NgTnvYr8bsTVLIm8z7mAYP9HLFYC
nyLlzCkEy3RsjTBnzeMC5Mq3wLatI1vvZa5CKN3Q9U1yh1UzHMEVWLfWM4r7YdxqkPVwDLlMTITN
l6N3byYa4Mythni9MgsL6TbKCDjUMBiEGvpAsqpAdgnSkUlHqnuN931moc806Kjot1GjHFfT4GNC
s08heWGjBeKfRjZcs3hsd4vM45GxrAb5yuh8YTVf3NZVKA0LYrDFRYMXmVrRvRaFHi1+BUMvNxGl
WV9IHtOf1PQ4Q79iQ9EISyNHeHiLfvjRdkfOMC7mINVnUp8nQZNn3Xg/st7Rv4yIwNzugPzG9p70
ISyj47q1y94Mp8vqdc3EucUqpLB5SPgNMEpxsfAoxNirhTMM/oxL6xuBit3yoTYlXHrBn9rk7jT6
Q1xrIt+6Qdr7vD0uy4TFjDb+Ju6ytB4k1RCzlxZptx0oPupirG60pxr6Po8pCF0Ua1qIQNOq6M55
b1IbI5azkyK9ja6CTbXRXNLdl9PCS/xHxdRx62K1z41pOeod4SidgZ5nZy2cwohEfoMMxmsUrxuu
8LP0+gdpseXuz8lWRMKVsVbqYJDjmMUdJJT1CYAFYcVrG57XRu1DbK4BlV7YbjEoVq8M4LFWWNjY
TySevp0pKCqphNiCBwoAT+LRUzF7ddOPJGDg68Ijcbq14lowGU/GksR7q8sINfmROVIgvU0wfLaF
ezwRUaCIw9QOszUhZjbV6qhvnt13L3oxyQIeFG4hUOf7mStlX8ORNHYfVcJwtXINZ2mZe/qcYiRY
J3Kn7cArv1uNdCFvdYgoaGetkUcXP4Zo4t2vHdpqImKCwjrPHLncWeo38XmU5FBUToEeloyUN6Ru
eFjoetbTr9/M8r7dFsJkIlmsrpWxK0OA6xvZlh/AQ+4rzG94+XZfOggp2neoAysFgK5Getn6ApMk
olYRK5QKyixxv0m2F3/NkVyWeHhMeflJ5A16/4FzWf9jRYUdJbqpky9mfP6BHLJzfqLoSl/2tum6
Dsl0dSRFAfceUOJ4E+4Ae266oG7bK1U38OlwzNDBL/4pTD9nJeeacLTfqAQ8EfmVmzxXrQ82F/RE
ys3Dn6VKnZ/zJqsOGr40UQ9GG64r7iw75TpNop2/td0CDLPbItUJV/CCDV81Fs6wSs4VYfm/CxnS
kXeempcsnYXuSkjp3QTLYgeaZPjCnfj/3sicxROgtBwM9bPYz7H3dXbHIpCwNXecq1zuVkG5Fb22
wa2+FjfCmlsadaB2UZwqp0iYqMCteeoqQB9kZRinemf1SnI0Y92FpPBYvKvzZfl3aSliO4b6G6aB
xf8rpuU/VZevPztfoNJq463OJgvinloWxlEvhf8KTkxKIIP2+LBbUjB9PwNM64O5MeZ75oR0FzhU
qDTtYJQA3/FR4zdXtvYwjOg4w9pHq6DLhsxctxr6+8ayRS2UQNcxLouPDVPepu3Z2iW/2FfIMBdn
NJn8gfJ4X5rEAAvE7wA/6lkV12rruguYZtuS1ddIep+XBbRXGZVjb5qHSA9HO4P2uumIB8B+TYY6
urLhZE+Gdq96whMKpwQFJvWFzIXQfwc4CeBaG08m9/p1QGCEgvTzA+cmRR8Y6HyZdl20NGjhK/ax
qV6bcqypT8kR6KicMM/4ca6HR5layFp67tf/gY2xIMBceWHb+q2lRzWrcfZE4Kt91PfHu9Ij29j6
h8c5aGCmGf+bUbaOQC4JXIhSlXJE1iCpeMHB0jHPpJkO8cAm8OXc/u3ddXVK81PdnFOb5XffbLBS
BGwIon4qmAimP3pwxlO/29bSjWP8G5tesLtwunp0qAlejNZo0KzgUoPui8yJdQ+uKUVtcLDFVDZS
vyhICqH178DATSvyCCGxJ3jWgx+3PLz//HBktN5SeHHMHGAKvWCbBGBiZyVFBOq/8ypAOC18ece3
lUQVyBEAF2vcTKnMgyPt5EqxS4VdK4oeSDiEDWhfVIsQqK+ksJCOZIyJEbd5m2EIC6MmOB/cuo8y
wsNFfg/n5HaL05xXoNnR5q7jscjc+MJ7h3lbt8WFwPLOEbTrl5VZppYJaCpy1YTvdd1lcFJT3Aim
0yzkqVkHcGyFSJezNohj0MytXtx+xp9FAihQ+vr+xOiG3obEG2tUkRwwNTLBh9yCnq9eUwQ5l3dY
ki1MqPs6fs0Snn9RPtOh/N632qeAOhI3+fyIYldxAIkWGHLQuwkDtjVvW4qvr71CzXPKpXS4I48H
k0GXf6RSSjPOzWOUE3JwQvyIR5RwiSURrjTdH1sGQAT7haARyFx9pOM84xM8NCkEqu0eJTAG2b9b
Y7SbPyGUb8A57B9cgJCz5HaLQ1m4HJGkGugZUcm8cG7vodzmUUliKOAT6ffW3lZUF0MHMAe369RU
q6mbMuZ0qLJ3yAv+WRP16NpnKEFyN/S1MWLmFIDukEbVoFu7ajaaXi5gxHR99FtjPw0D7GLzwhn1
FBJmzxLGPpE0G2jdQzZfpsZFC3qQAFfhKV/0K5rHj6vDaIgE05LlpAr8DsjILVVsQc0aNvmltNAL
6M9X/WRK2iLR7d9C4hSRRD0CXUU8lKsdWuzcaUNe8secq/k7xaS4nRfxSmC4voXm/kITYentcIlH
v5RSeDcwJB6h8ucbKLpeBqVQ1eopZhbuP/UiP/7WIdFl02B/Z6Sn8Sl7K6DOpaeCJk7XskRrIVeY
3VrJQrZKqldhyUxgPOzs4XMOpgBeM2Ni68u76/IBdmRrWc20TGMtBZ5Kmo9aKk8m702vHNMuE9Z1
9i3FFs/TF6YuQVa+BoPZVlxMc0RT2MG+zJw+eB/xYDIPfYz9UGltnUmV6sScAMilFlV4lTFHZjbP
gGYIJF89X5p0kBM46IY6L3sz6GRsLF/lAG+qg3588TL+ZCJisSw72AkR014PSqJ3aBhtGRj+m2tH
VpulijTEvI/DO/As2OWFqZMsgJ/niEd8TPbz/siD0xuSM8sPUSusz2x9zhSKjxfEohJAiMspHBHm
fWMKBtjAGn1Oda0QRM5h/eHAnJAQ/TQIvVfhDOvpuvQ8nxF0y/qjLwU6EeYK6+bOgc+Y6wW+jxA8
//8Njbay96eKwodHPl0PqLhp/ouCHNV3VrXVuhT18LdInLnxABEamfDg22xm2Mh2W8PNj1KwzeF6
ORUApDbDEU97wFSmseBgAJMgxsb7BNiWgRtZHEcnPTTokSpC968PEtBJ2x3HXTlAzfN0Y34idN8K
GiNBZ5Ub7mgRE6H38e8N121dWr7pJ9Bcpa9/OPo19DBLzPfE5keTB7N7EI6b+AntFqVkW1sg6ReY
e1FopxVQTsM2IQK0zwAD1enSoCTdj+en5qBL8qIRBtRryfv/hxJEOfwUVuCQKssD7BRFSiwgxHnC
EqQQslCSudfv1COM+p+Lxda61ekoeTKO79aLwXntsuaobTVpPrFP16yKAS4ZfT8LXAVKaoEHzbwf
VgdLcqJYYZh72jyPgEnYqBgKVaIs+EhwMRg67QLpsBJUR/4UA1JJabkLwX79RyFsfOufvQjy7Nt/
U2VjBHnl/HcNv4VR8Pz6iERQP1hgLzlWAcWwBoH+su9EZ4v7CQrTZiPTqRM09tDcsDH2W8VBpXYw
6yDssvY+AcOVIPj5DZmZza5k+ldz0eR6D5yqodPS5kTdpyJCago+7bNb7/+iwYzDB5k4yOn6IOdo
204gjeHQmykdEBcf0rgquV60g9bRhnyRD/IMgswb+4T8RY3g7AE35HG2VscdiaeiiL1FkinffA2a
Qlf790yMkTkGtkzUdSuY2mF7o/YQS50rNfkHps78F0RO8aL8O244B3ESbX9p1aZyRrW6cJtqox8e
KDUQth8rwaD8+1RUeM+Kj/A1LKFvx0jMfvPWH1OgPFY/CRPxFjs0QFop6NGEjqy6Wz6pSppFl7IJ
1qOB+/WsYPt9hI6gnHF6dDJqoWRIB17MiGc2gUMThMNWWNbrSIYqu18aaoTyYTyjRwEPOUSvVzeo
C0kxurlIlnfXcQgydQBpKVYbUXa6UZRQdeZlW4/8g0utgukXnSFY7OPax2xjnjS56gSi8HUyaRCm
HwEVAYQeNBXuffnrxZ1ygUTL6iC9qerdLY+cQgLBufeGfrnPUaKdrPMvvhMZYHberlsO27mEDGMu
FLjdoYV2MzSJRyPXxxG5GltIVyvs31XEvOis7gH+KpE/I94qXevohrQMJOeWSBIpPPe27YlKGZy3
7JGgxiJDejODGHnIMTlxArNKGF2N0cQQBtUDZLcWG66aL3tmj3uxwK7L8XhrRHMl6BHvmstPPnqd
O098mstWcWs8jsHIOh8/zyqrc/tmhprpW796iAYmfvXATC1UCRtc8Iuhy14HoO7ZrgHwThhKOAt/
rWdsOM9jyVawPPavNsdLzFNf+QGTFFNShMPhYvYs9UnKlYtAYxR0oYgRGcCd580KY9uny4hoGWqd
mUBxAgphcWoDHcnX/2/5LhWrTWqJh3fR8lT+TpQ1H7O2Gi8XdEXP8GY602/GRgjxaFjaoZ0Ssh+V
hvq74/bn1ugnStVjCDJku+E7uxLVZGf6A/0+vHkl8Ku1/KyPlZF0K30hhvUOnM0qMpH5ryK88JC4
4pH6IKWc2w1Q7+pPZwjXwatH6kMP1MeGnqL+e5xRl5JvDYEXzvsrPZLVN9/Y8lpizrj8iz3KrmbE
Ykx3+Iod82VLYDzjZbHvVNULfXhdb5z+CV6qK3ATQWd3RljgiJofYaPRp6K3ofHvQRMKzgjZBcvu
xAchVg6mkq9k50EFT88bpi5GOZDWmt6UyUVVWead9qSx85s//5m95U09IPrv0lLI2SfpLMLcGqcw
xiISwN1/0K8CLdAYIwsKiuil48aTA2642tw/K6+v3oYE5qHp1tUwRw7n9zDsEpXn4/CHa7HZ0V4j
IjchuGvlEflQlQkfHpzWUnWuV/OAwC+T0VP5GoPin8+jj6OLDoXT9r45Kkg7LuUfGB0cIphOgtT1
SXdR8iVkOs4sbvJq7K+nqk7NGBWZYN9yv2W+Whzo2fsnKza22ley7pzQ5GO0swufuITknSv+/JJs
1dUGhZfq7bZVaA56UekbS1R75o04v0qFT/wvfzmLcBl7prUHZG1QDkHATRNBVpFm45qAChCP+0Jh
DrfodcbtxTJtyEkWXcIeuuF3CZIC278i4zkAL12wkSry+XqoG1pa2piHgLmuHtQbKV1u+mlWiIbl
BYp7JA3X9tgDCBE07/DrxC1hmPTDy/oKRP+W0jYIGQwzDaRLUHsUoZoTQiNaSNDE3ZClQIB3PLcR
OixVtTnhKg/qZ/J/45FVYBvvXzkVO+wRuGCrbnKxTFh+kShTBauUH7t+84mKsrpWLKj+QxfT5Eqg
ZQcvqU4GFOJR6jF0C7ChsnSSF3t6vSXXGDltE1cRMxY/AkbLWeY4Grg4Zj8IpRYk5enBDu8628l0
rakSTjTDxJfFuLzBAJfyjaAE9RJud2wSaWBcXfjZkZCbUZLk09VxlEUEJQdJ1HQHUin+E1Cb5O1E
k6xAkn7YPAkho/yZ1NHInVZDQ1Vghvb9c4vbAWbQOvDmfRW6szEhM7sPgnBa0cmtQ12j6wxk98eB
zbD7fikDToHCtSJHWHRmBATySbJPx4PNGiD1c+hpxeOuT1OQc3KfAVsdWKUczjBOOfgAEIAk02wF
YShSlKuUMq2cJewQJAB6FMdRBwZ7WoOQDZ4DUaW5hNWuSDXiJRSlX7HfTgIuwmvVP9ckuRxTK96S
874wxlz9WGflXn6BgNjKUfK7UUykUBnYuC5LlV0NiO9uaeM8w4u7pIF/mg3mecViW97ptzn6XFIj
g69lM+hmQrahg9seb4FKnn7EqRW43HwSuRpTZcBP90SHeRVFdYLsjZh3Sec7SDoXx2iCtr7NH8ly
5F8Sj8YyXyvjW7IHmR35NGbLMPd0zvk7EQ2Tivci9iv5SxNdLmdd6PNY2KuWzsQe39WjSFNJJYiR
m1X7ARRMRSSz2sykxnDw0aUDU0J5sV/YixddPqS5z/eqJ1oVW96psfpMgl/AUsNPiZxIRQbmVmGb
uuwEzrhZRzIkcFxfS15eh2WSGD9Nn7aezOEmG+txOztUidRIayBdaNHtVaFAVigQbOjqGTqPRrtJ
MQayKzYUqNW573enxlow/g6xGVyMJBgj19plewY+8wys4JkUpG7rSXqpl283DVTM9NwUwotB5Jnj
g/DUk1GH4hj0zgCHJc1RWwyEufgm7rVZ3pqWfczMSe+5DHm/w4oLHakw3cq1PDJBgoh6G3okC6Hk
LSRcZ85q0QG6zO9b4Oz8mHn5Ast+BuaE0K/EuydMfDyyxSrNlUGMPtaOeMflOzeR8MuQv1qZruC+
Sn97+q07OrXsVkNDudHYttEDrQPdr7pyHDEYvc2rVcPfBx30PRn+znYWs9BxkDWLkfWC5o5sNwe/
Cap6BkSBEQeLFIRWRikB21EWRgN01v8PBr6PYrnGlJThqC6cNVlA/e4WqmoW+8rM02Vo2G8kWcKo
i5+Tb7SV2NsJg1F6cdEPB+ape+wUiVDTb37gPGSSqe9Y7q2c2D3+lVeqBZPs+u4KDvHrpsJlxRah
ubrl6liwnnWK5FAjFLfnQHSs5gYlJHOcZqbXzjb1iquBlu64Ni6I34b7b+01fPX/qWWsE9nLhLBp
EnBWLKhI+BESCLG8UWnd81C5eyRjr5ghiLT5AxD1eJ1dCHrEtgRuA368WZAP9ISaQpmhdJ9A362w
De6XnKKxytsxpkmKmF1jjau6+1yD2L49aWfI2751224wKMfdVxa5U6KbAFw3i6uPD4E5rU1qMyDr
7K0jVdyj3ArCwbX1+rxLjl8wAOqbAZcEcKnodmtaYYHJk9Q8qC5cv7Cc9goZN6gYfnUJ4Pid3mRQ
9KrFuXwdXjrNpi3oohtAVbSD9xry3Pt/BOQ+8PJcniTX8NncbzxGmG7O+xcenobvhJN1oLOLFxjS
KF6voWoPgUzMlr61IdTzzjxXPvVCGmrY/gyI1efY/SDrmfyWR75ltR5MCZ/G0sp3jNpPWvrwVv3c
NiYmWfo+M+JF5Zdu2G8sjclD/2Gowlxiza68y831A9xn12xhNIp/dZXDevQ2270HoSTV36STEwnK
sBU2C0kqXYD5u4mdkq4FgvOyqseirslzFzieMVo+/ga781G4pqShaE+8OoVej3C8wGf4dgTfb9IF
z8oDQcNHZ2q+DPJgnG9V4Q3vKCR13+OL2nd2XcptxZLZUFTNYwm5dvZwe7Khp4BLjTsji5uyJ4Jo
EdBhvkeIOafLJ/We0rZztJ+q0Ls/5J2S8PdMsdFpYKRCHdPTV///Ov51tzQeJPtQrzhjKGAxov+9
nlv2i25TZ9368t3PInbrmKCuFocOQMVdAk7xEkIN/IjqY4GF/XEBR9TPGCsB7sOeqC41dHTMs4+l
Buk9yw6ZfRDi862eZPMqeK/sKAUuhACyr1tWp0H+2QCtsn7/h4OB/tTP/Do7ufYwRWnfPcij/4LT
VDLUF+MPOyR6Qt/LWIbpE6WUGYkFNqOVj5J0OiBMcBD6bOINIEsZHS37qtAjDCv8Bokr2xoSjZvC
GMnBRY39I7nFMlDyhj/FgbT/UpG1F7i4dNeVHAj2IqGPAf3Z2vkmuBKHH7NhT3H5V+uJAzsJUeG2
QRSbviVatVjw55o8dWW0n2AP1boyOl5f3hY3Rm16nps+ggsM1PdNIBqMlE9J1X9LGOVQJ3YuJ5eZ
LSwUw9483Knl8PJl5BV/W+qnGglWk5pxFLrg2Z2KiprOSFVp/lKHPdSJyBgL6UQKymSdnTE0jtTC
PfdIcBB5lwt8WrZYGFGkYmPVoRAEUnK4Hn4bP1YJEFuDKXLwfbdNAHff5pFKMnvX7SE9Q4igrJiR
AgkQOiM78izaar7nJZNGXBbig9swAIYmiJ3TnLAUcp87tYa8pQf0s+ivciY9O3ixGVjDr6O+UP9q
8+FHxbD2CKg+G7ZWe+E2SGiC/r4MTusvcgVIzxr9INK5+1wuSjVs03oKchioX7KAWzHuYkpNY1d4
dW/xL91+fsI86aMf9lcJV8YtE0nuPDYrVMgCgArJvdjocqNhq5ye4HwJjSuYCPdDh8KFi85IOwgC
mrLVG/Lb2Gqpa5capfcAf73mYO1fJVvbfS60KbXZ3Ik8YLY6jqhJMq4dQlZCd/tbUu18z8Cab1+x
y8JUrjTfs2me9IlpoLxfCdZdup26vE+1e22h++Ho5IqqbMDk69S//OCEdTKz7iMtvPeBzxs0f9Yp
SIrGXyU5/TeYzhgdQBBty5CZeGYC8tHBty0oAtpVtY+XFlx39710fMDszwwYxzLKgj/FcRZmnKYr
pr2E8Uom0DHM+tSnsXmRlwwWxel6rYUzLlAK8yW5Y0CdKEmST5W1hPMfTuYGkdqrEDzAGuvHMv89
bl2agoTgGtVvuLeyP6auZelJ8pV+mpJFcAkrrKes3p+W7EQLm9NtYlgTwFdwOZJfIyn20JKFexQO
dt0Yw/eqLNX+m7DOK1V4X2k6AJzmwHxxcG7GpdYLp/jEJORJj3ty2N6nxSK2cRFD2lAaAAKoXcBt
J/zGUcE8VwCOSatc6JDN7z4R4e8ZF5itxAChPFoW1EGm/uprW9UjbBVpaiBDJzi1RC2+TeIV0xix
g+UpoZfHcNf9VmF4hsQ7xeFLd0A0wB5mnkOr558S7oZ5gMrxnKQ9P1/eMkZcp0Gb41h9ey5DcLIn
hacHsGMrJdnHO19RpriFH0DEeGe6OhIsSFs1XoBciO9DAaI+qA73R0t0RSdWZ52LYOLiObfXtsxb
CdY8RDNw/dpZcvWgbeMG05shSMgILrqt2/PqcJoYpfwEHX5t/lhckY7lfh4UBg4/x6zEzH/NrGDy
aTBER6hA14BWUUPEwzVkVG5J85C/N1pFqldCB2Y/2+1Gj4IDS+Zk8bKmtkFBknTxA+yAjJJ+Z60m
jFiFgqQYS+a9lFYypJp9ncSveQXQzAV3Pl2ZFAlmpzKofJN+3dMLS+SMhd8xQGvYFk/OAqf/mHeN
dmd8WT5lYmDOQAhxtrSpDhi+GstHMQNigRhsud49Voh/KCHa4Cq/Oe8DmfnU9f7XU40cVkZ6hFoU
Now7gxAqiF5PfEwlt03XQKkrUhoH+xr5SFcss09r791f4DKBK6Svq/jC970HVrLZIKbjLkqr98TN
WFLPv+vdOSJOUlh4FpcfQrrCZOK3nnhIeUnkzPpfSjviLnHlS1CoNxHfr7qEE4P12a1BtrAhWFCV
pYiJdhoUa05WimRDTiaHbQDMuLVsWQ1cehdc7ZzZwXjagm3nTRQPlKLa7tsk854jJbOqFCTk1BXO
0DY6lAVNM9nzEj9NL8RYEZWWjGpmhkYmisVrBURB2awzZu47RdNXjt4pwvZyxecD2AQb/Jq4ddMG
qzXO3sXQovdVTQm+hOAvmrDltYUYOrj1GsvaRmOS5GbH+5SujhCc/WDt0HibcjUVHL004MXolljR
h1mUER6YUMsxSI5DpnzhxdAKvi9cLJ0hvcBhttyRFlacEoflPuJOuldEjXn28zx2yBfXpPhy/x9w
RBghIY5UP+Tu19egn1OAoOyMtO0OFH2BvDV2qtwpfjV7+lyvenXIXCmKxw8HzyF/wX6Fr1dMNEmK
CWIe35jE73nVqFcsDBJi3h3j/hbFc3cxUFNy66QE8tt6cZjV4fDw5dhsiiQidelO/OfmtUUKG+7w
69tUhAIK+pjXjoXf0hBYhrx3Lb+ft2yUHMw0TKyEbiBnaobS5+dnMq/BJIixi89SAjUfgx7nqw5e
w8setkGzoK0Fs+Lx4afWxeP5cOTzBkhCqRypQRPXo7XBTSntgMTa0YCVIAzqn0wlaIBCjrRO12e5
BPFgfdgLZjMqMAxmpVrEFWtLmcbfxcLfBP5uNtDAaX5EHr3pkuf1YWcKc0BR1zLtu/0g9GGhXwy9
73sYAL29Z9WZohpxam0vdH4oQF5IwJDgK7QlJ1J3RCORnfQrpXPRbiReTiR8/rFLMqPaubrNMGgE
6JvJjd3Vnxyqw4N7JQEMFCJ/Igru0hOsNyIFWAxwfGWoOllFnz0C+DC1nuop72POMn7NBw9KVl0B
WNtYIVcDpMabEfnqW50IWYfEjOEZHeUZ2v+GrqFovw0Rba3KGzQrnFPlLac/SAvt4gTTyjZ3R+da
pUQPO4EWkmQ3kRX8LaEOzRCCul68GUYykAW5uEf0DeaODmc8iTB8pl5pgn5qCR8aF1HZzMJv4K3Z
Vo4OSh3RMndtcJfuSSQAAxjXWCBX4317SnKoGhj9dUdD1hHoeeUFbJ4N2em6VjwHX33EsD/xSLO5
BcRXIR7NTLaEWkkYdRF1T15mNBEEK7LpW3UGiI40VXqlU8yDhdlfWf5vgwdkpYuG/57G4Em/XU6H
s11FpalVp0SbUB7xRCEUsX/6m6fmf/CM2SFHWShYZkJF5e9LUa7KJeHAPdDKTKC4KcZ9wPAg3IvR
IYWk23JgB0In1kqUu6O1prCkAaoQGn9oGGR2tXCEjmQfarUrcA2ppHTt3N5ZYCJ/RSs8ORxX299j
3njw45SE7XJDBXnLB2PjM8xf0I4soTeeuMNgKLHa0XO0Ib672yl+Cc9+PTPH3d0WonH2vWeqCAi3
EnXLm6RtoaF3B6aw04zIQCdOPYYLURru5/vXbDU7Vv6XujRdy3NI/SLGLroY+EgnJ5NX7VQjEW8s
5K25sQyYY4/9ha6T+weJN0242J+lB3yrhrH2MdikL4sRf9LqM4PoAo6YZvQXdLc75Om67FOFiFk2
q7azYFxymK8LfDZRIxN6O0y+mbVSmE2xfmRo5TgGdzA6RztJNBnLD96rRJopl/f33HHdYv+N5E9U
8C+1B4RHM/ElCWWC3Tw65nGpe5nIF5uQPjMfVtHqXA5TJqIKS/Orss8IsnYKDxKE8QA7LdrTscjr
M8WzXYqvZdtSWUhSMP7YGMuNTgHWEP3DuAR6ihvLwSUKE8BVstY1QOoEjHBDdi4KaQPM8qvRdXZj
6qtyuzbkGQGsI5m7/kc5VTIycHGw71FYWL6kgf2kcesCWO0t5aJAbsrs7kAA9ybN3H4cjJbMYpvY
d93tgVqvV+Nt0+iO2UJQtajdiDwaIfbBRVakYZQtzHtpA7kKxXEKmix4JZzhGBz6o/7eIRamh7fP
gXdjXw8oWRwir2DHlbuNqtp/R2DRJmqUxZ+JsDBX4IJhKPOfBkoaDw1m3OIl93lCgNTFRIX6wvaO
dFpJjemFT3ovloZOPczTUJOFifZmDgi6tKHzWqO9NfBTdXr5LnND1fFQ6Ez6VfLevgOXtuftZoVd
R+lxOqT8r0EukzKWbl0VHfbvGhZq1/AvQVd95DLqGPXQO8u9FFy3ki+7N1JVjZhsxvASndbOV9gq
SnQDlIdMk92lF2c4P5W+ebsoYHPMxZARfP79tXquafoCdfOQRHTTO/znr3P7KvBVuInlBQHU9Rm1
FscEtLK3ENhJhlpjks7K1Gwy1xtn04EPI8J3JDwQhXX4qTWqQlyqVh1qhGKFdAWmNnvXXVRXJ8wA
SzQ4r/huYWimkTR8vNatWEpZo0dZeSBMGC2WpgjZO8FX4NTrLllMfDmh0E9WQFAIlGco+lzefMGE
SymT1L6Ks+hqgGMG2fJtIMSc4ockSHdFffkjLZr4MI/RkQB2hjGu1k4o1lDAczN+tv3AyuGwQhZr
ImkmTWTBC0DL4CxzoKS57qTslVBwngYZrDWrdrfKYQyOS0s2opbIaweZCCIxeg0LA8SrfRHLdCIA
JN7XulXiqrhaV12Jjesqnduf+fpqmWRsMpoVav4ARomzPpHNQamKydCrT4HXG95O19xiUyZppnC4
kzu2zk1WW+Ccxo/MHviMe9WXLdOQKyI/3HY2fDUHhFRpJwkHVTivHcGRtYiQxbBF3SpufhyBhedN
f5Ubz6iktwmvqH+wTzjQguFKfnFdcy9vexaF1p1fLs9iGX/ho9PuWthMY2OPyEr3p6BqfKXiwzMJ
AFMZ32pquFrstzs7hoFL42k2EZYNKqvTRzsTF2waLCQBfnh8cdEFL7Ml8/C/4fVIlxWXWWG5b+S9
SrMuyJID3GgaxlAvVifacCtX205Sa5DFbT8nNWI2SV4G31ugEo5oGntwDgS4mB7oK0/DSdUrs+pd
rGGZDS/Mjbh1QYQiLgvm7sUwc7BsoRxNxo4ulvRI6rSEcwoR2q7rJGoeVpvX4wcX4emlbeXaY1Ps
ULlrC9VjiuUm8A2z4Y3jyA++X3SJ3WHw+15jNjBod5MXd+nQ8s04dukOUeAL+PCPwVe6hcRvNgDH
btlfvIuiJ2lidvGK5g3JgtVrvuJqzSR7FCVUoPJ/ftn4rF9WiKOfw03Te7gOlz8HfA6bgjOPlRAZ
+oNxEESUYUHm+9YObUC9cbJ9lqm8fEY3dZHyaFQ30d9BDRLJ1xN4YEhIT+g+a7gqLlRjm0xidvys
H+zjjxIdJGp2VHTPkwB5yDrLuaqBc3E1P+Mi85dMd9jP7scNHLRwHD9VtcI/3YozC0LlyGvjxElj
IKWKSJJh1GK8nj4Q6vTu4upnn2kRPOojIQRy5jpCXCjAwSVkumFPLWLoqO9SRu/iH2QL7Ye1r3ot
zqLXkv+kFcAIpNHg7GnF7dJ76veyz0nqlNOv25MndQJWpHaTQ+msSE9AIO9Jh+CrkJhzMiTZ3RBi
ekjYV68Rei65+pyGF4LF2zcU2vSmwGasSn3ahfcBCn/HQJm8zoO73C1uNlH8Y9juqASeNBR3hEnc
ueOIwjKeCfMm3tSXud3kVGne6UTN9e8fp9vy/gb46PJnJwZdQD6aMLXMgAJIUjpyPcq9EQbX3JkG
IT2aTkULdwg923WUCc1lIJ/ZnJ5rhRz++Uk3tZ3q3Mo/OqLMs9zyTN6e1TyEeubPQnYYidWNxz2R
SZ8UW/8ryk6p/o1GzeTiobd4skZ8UGod44wseuoVo6R80cwlCxQpBs+mLlYaoW0/emz79tyoIHYa
PcFrjRgsc42iyXzuwjOVfpKWvPLJ1yU2g1LwmJtaiSQU2T62bBEwhAfAW45qr50SxmheYZEs60Ox
GgivbaFL0z5K13UGmKlQXkL2mX/Pw/YAc4/XIK13FU8VY11YMlT1pWREAf+nk7TuOZ0o9GqkMY4h
I19HhmcFPCR36nMHxTNbp+rnLFtlvQC5tuIdF8K9kknN9QZ2QzN9BsIvqNToY6X5a4Q4ZK8fJFLZ
rwlKOKGpWGVutqHLTVkRq+IIjQqdA3n6i86XjFFKTvooYsb8g6OwM+Z4b+vbG89DEevoFFTCCBzG
z8Z8eMYiMqS7FRGFRDpXcmUV+CyP5lQBh76QAXqTI23An/XIW/C0O/YuLExBrwqwmInC+dMrn/OD
Kmqms/eAvH7tCuDpzVoL7CaM5EUmUwIRMGVHAca2ZzNpIQAaAte09jGKMRdkASM8xgoHUaGC6xnz
1sAcxOauBr4GWXsaij1mozvarvT4FjkUzAaEX+ULaCUx3JbvTtXXyR8ZmhKande9YChElIppwjcW
eovc5MsYD1CUl8WvPySy0/9ltHq3wDiH4MUeC6tneJ4yJ38YIEj+nLMI3CdlMcQ4UgjD5aj+Hr/w
yikSvbE9kInhKSpua0nL8qu5mLZTvKwOrWGnXJRF5D5pnOF0igXz6SHdThwHButjVnKXWWRbVk4Z
tFo1jmS7c4I76vNllLQYi8LMl1lzTvq6W3a8c4aHHTBiF4/5OYG986UxDntAlulZBiu3unBidimE
p1o9ua+7p5H0jtSkPlhcnj+mQQeuAhn7PtyKK7JRUs2sI/xfnF3s5NeaZ6HnCBGM9Ta6nuGShDZn
qlY0V+QEKZNSRk0hVWUz1h9gf7o5tjFNpMUhT2j4DTo+0ZQmyoVImYDNRG9m1P/QSKmg4vz+x2tm
I+Pn9rngsGFUkCXjTscSsbbJb7a9/LwZvaMnsb8mc87qpUB9sDB0Jv1oCWEU1kB7GiKFkq7pNklw
YyDxwVqJSrAdoqZYxMn0wgvC1UN0vm1StQx48Ve9ZU8k6SkQ4XOrBBf0j+Ihv5OHKmOjprlGmio6
oBPsH3wLTzJwJb14EVKlR0zC7jxLZuptvZbUBn33xRLIElpEVBJC+7K0rqQcoh8BwosAdpZ0mBPv
7gdees/NEIpucBqogiyYIW9IRUlccz1fqO9QaMQuUv64hImh0nANyE+wgB/c4sEcL1SxIitorbdQ
fkutsr/WKiJvcYrCbD7/5+LkkbYmi107x5KbetIfFRMGIx8ikZVeNqC2M6CYtZ0wxFPGF6OrGAbA
s0MBFrBlYf87vl6NfvIr2xUODRIkd/Jt3sB4IkNcVuwE+2550onAB4YP0mfAgxoeawmTEOMAD48D
ci8GxlE6qO3SsR4P3F6uuJVLblKNSedtZInlCm290hvclq7zHaHgjWSTSNkCBvCTi3N32asY5g24
Cq3lBtZmXHQewGP+LGqxAcwLH3VJRZIlHOjqLIVgqDLs6txbSME7GUmrjgZmp9fp0U9H/5ljzvNE
NCUkX6y4Cw8kNf5dkVITNAlLJWOH+mJFXAUqNoEVdVMR4EviAlwhs+Ge2hmCqFsM9CV9dSLIs7mH
EYqZDoQ5MB431siP1nE+9m0jV8N0qp1JBxMneUC4XQ1Xrodpdzl9tr0HHdYTxL37pTDOYtUWB6yy
Tqscr/STnnpsOPx6m0p5i6xnw6isTx1c8HvEGgFeHQBKSf/p4bk7B5Uhuk2DDHK1xuQHNRYmPRnY
li2gnEerCepgC5W0WW7LrZI+/oPIq3LklNozog0XXTnE2l595pBGhz5ZBOO6D0c2IAgEKTvpbJH0
4awEN0a4pEj5047ClAVkTKWgljGX1rYeMHjY9G4u2gSs7jtokSM2nJT8IAs9H4F1f1xn9B16nQyI
fdg7sSOgoREWy3Gv3rsG1vIEtFQlkksVbHqO2am65i8U3SPpVb/pvIZS/7EtCcawFc6LdTztQV52
xTAlYmXrYdbpWWNJep8l0Ba+F7sdMzy0bqqIc4V+A5uT0kkfz4PwNqlpNFf5jewj5P6KPSc6Rq3g
ziX9gnUpOmuqcIs6AeD1vazAa1/1wohR5RwFCdWbe4GnZvvTDYspIMocsnSSuj013/GefYfZR/ZH
yP2ywpybM3ZVLXDK5xgPj2UNmo54KxYoiiQH1hRUiOoY1ccWlONbL6TN6Em5jUbsKOjxC4ovKeYc
nCgRzVjtKj/xB0yDOR/xL/7V96zqv9TWzUx9N9xKOvRuoROz786V3xrT/lO9aQ2UjD6VHzkH4RZa
zdXjgCZkjP7EQz7u8yPpdlknBCfyn9AvhmCfa8q6senJRf7dYgvmEy4LN9zv4WeJGrFaV5UwgU7S
ZeOlRoVHCDxKW2xxVSg4r7EEtW9ZPZe1Vgac6OiSD0Bmo/opLMseYfCTi7JMPIdPfc1XBiJk9Zj9
SfZ533OKLfMuX6zW9ETGMzaPeLlcS91TmvVqaVR9O2wDt76+f5vWeTay9CalTi98qeqVs9p9gRri
cV0X76/WfM9g/PgkSJ1VACsZLII7isWeVFH5Lj78mRGIZi6rZJmABVMYX8G8FaBVjHnBF9geELYn
AEqxiWkAibKexme2pEEEUptV5PfBNsT6XCV4L28i6sKAwAnGrLU0qIJgMCSqV6dsOnT//YhwqD+K
Bukm6CqvZp2NyAVYUOYr0GbFK5l78Qs6AE6Cbr8N8foNdbaD5mpSPm7XAyYfscYcN2WEB+C+UJZf
2pHbmwWsnLKDDmK4cidvBjWae6j/XKAfQvk0pM3kAbqjCGPmiMquOAmOMVy83YP7YgTgSLUJJGHE
yWbvoXDhX9+cf72vJ6uKecUsTr8HYF41CMhzkY2ACe7zQ3x12v48tSXTGDUSUZuDmVCEJxeSSnV6
8cbQ15Nn8Ymjb+gneRGiKaEBIxmJtgVL5aLgNn/71yB73DfpCkuhsK452P7THWeIcAboIJnbAK43
e5Ma0Ez+liiGT+JWuzAzBQNlAvQj/vZjqEj2w/M83d21Bn5Gq9UKfY4p5/skbe2LR/w03Sm+yO52
KxqJeRzNWCHB3fMfK2JWKsXCBqBT1c+T5pCj9BExdAQEAsipuODv8I1sHDqyJ25bViPMBO8Clhql
VZnq/CKkNa3VmiYM3W6APPpzj0BopbS92KpwPIM0Cw+icrh9dF+YGwr36hvXEE34FmnKFeM1Kck8
Cjj6rzzftHhrGbgtRh5IUa3JDGRR+RnldXRikEGJq059HvoFbRh0VRyyUVGORgSJ+F9qicAsSWB2
9g0j4ejY4sJ6se2gGbBGg7bjb5U367vrlKVNq1W+CdmcOJDzainIgj3AjEugXvx5pUw3V6QZsLEf
U+2BDSQRJM3Hi/RUqcUk6CJ7TyKF3KY6zvCPy6axKV+44PJ099jvNuCNbe+qXz1t4VsUmmjLL11U
jECYzSonrESZ/l1iiRt8BpV/pTCYOaNy5CQCZ3gw0It7ZyR3WsO6vMcMjedJWcvP1aqf8rJktwRu
FQLPb9D6ADeMlMwYeL3jlJKPd39o4pZI5KbAZN8MtE7u+p8vZ3TyRxApzjp8AJaGdEj+2E0mlEvu
zNBz1b4VZUeuNhVT7OkMh2+bNVNBnLPfTrruBqmDcA9h78KRTcbpTDOrXM343tDxHM7YtbMHF+0P
oOE2iZOlaq0bTvRvuPwUTbzXPjxPaVUbpYFGjExKxr8vl0b/Y8E94Q/53fe6qGap+6HBKkL59mvy
NkTJa5eynvSS1T1V8XdLW/65hkgGxAljc9PCYuvv0K/wm5h3B2iO15kf9R+gp7nYbSNpIqY0ZOEJ
h1eBnGzdfgH0Mad/blo0iKnnrdT4wUvU9zq2DZNX7KGNDIWFjXI53inKxfl3bqaX+IDyE/eBhcHE
G9TPzcfNql/lIa5akA3kpw6Yt80OPcGk77al+cmtDpgz0rRu7unBxZ0GMs0H5k43USLxNRkcur8B
ZyPuA7/6pPuM5nmEsTf98jWgcbxUGs+TsZb8lgxnMK/QphcigulGXLtk19wRgVvFF/wpBnXa8HaU
4nO2Oyh7clCSnSEcoEexWbu28PeAZOZLnGtfgyd0avtHI6kYymbsdK22nlcAY1obiH6AoQ8sgIjt
AjLkntMtypAR8+ABAGoIr3Ydh3H+infUHGg2rs5+5efbyRvxrTcqBeXMVLd0lPx1zx+/zPYYkBt5
HAKCQ5hMCtmX7C8BOpdj5Vwqio2IMCVHQf5QssSE8NKgnr/GysOve7P42tFbzUHw7+6Dr27zD1qi
fZ7B8XTJmz5Jyh0oAsFyK1Es5QMzRG/0pGNkNYxy5IIkZSezohnRAD7GM2aiy+mpLk5ryA5/C7Dp
xfKw4awwTBYMqF4ABSjPChtJSBvuHQM25TNBovgxU4uNP3iU7jyukmFqs8AV5Q+aAm5PshkRSVGY
EBw9v4GsEVZ5gROqQiqOOjqgKVOcTWrgPO8hg0WxCecFhiVhosYY7+sV1kFJSjKuhdH/Ss7AkG8z
4yJB5I6mc8Doumg3OIrahoxNgwo+zM1uU0E/a8Wqn6er45U/9IUQAqlitH8C6L+rppEmk5P4tEen
bQG9MLfmtf+bApwQk2In5zEqlzGpl2eONiRjuKmNtfqMbz/Eayg3z6bDqCMji0SKa2zS+3N3Sj1A
btNjN3E5ndZOm1nvfBRNRMl3wkuC9AwDoFhBq4E08e7tdUi3jqRNRYZy/9lPiQGPWaW80r9sXb1U
NL/nati8+iGC4BYyfxZPfOdy4CihswYYWn3qU0GupdtFUmVYzSQiJRLz3lWFutqfDXJBxgqkQ8ed
ua1yaA5dMe5wMfCq4EGWVe0BepSdolOyHlI4J4H1IU6Tsx6ljVtcBB7mUSu3qk+PHdFpuH9Nnq5W
kOffpM7RB5Z+HO00G3I3F/u5DCH/ZH+NLoz5N2+fAef1sCBOJjQTl9KvVUN7K4pELvIn/3KsLvlw
Bf1F1oBKsJ7iVdrFdLcdWyKG3Fui57V5cI25q7wsGbxDPQt2suUywM76tggi0iS+2lslV9XXhcdp
RK9AcswqDtjAMC/7aJ1gAmp1BFBDf2mzVsKgtQ5NJnnn+5FctlBhobjAGke7au/VmkncORvNn/Gs
/ZwojGkJSEn5r1A85mcDSq3vDn7Yy4tL1b3o2lhohiNr43dFnuiZvhnvZy8STlCs0Z0M5x7d/pmx
UOmHmhvt4DTTMXFnhktJ7yrJ5EuDMbX3CUTA4FNgYnjb9CSRAphLejSKTtlV8g9h6vPRKeZBTqWH
iPcY9M47zlOn8WOkEWiFirJfUUyNiHU2tbMTxApBXMoiYjBPdr0w0Z6T36yKufCo89CNgaLdFhk0
WJhcq4rhnj6u5FT+OX+aPuybPP+bvw8wBrBs16DPys0U1MB/L8gc++6XQLDDuHz9kt8QWg8LTNVh
7SlD6VxBQ0e/fqSSxT7xzxVH887oOSag9Ig3KBmbqwnEip6zGcA5PgKgAvXhkxCXLFziTkxrfcty
0Mnhz36Vp9vRlVlIDpG72+AsGYSsKTncYDU6AssD+wBfioE070LOozADsHoksKo9rb2JHaeoInSs
gYEpMZXb0cH+VXDoQVyOgpPIn2iiGHrqQqRd6y1u4FcRwHDB8RTjIPjqqLhOcmzrv2HeNMKBO7Vx
I7suGLioQgq89rr/a2YAlaif8aQNz/vqDHDKbXtPm9aOSyXC3z0N/wxTq5UVKIIe651QgOW4Fnf/
n5GudMHAbYEu+BU5UHe4mZ6cMYh4XB78+HCFusIGv96sGg/YEN1QO7B7s0VD3TeUO+DLrd6VzJUi
dvcza3CkqFt8bo1TYb6eRDZHkKv+C84j1HgaOt0LZmgj1cUEvIsxrAf3Z5UO/NvSpxOQ0yrIqKVd
n3WOgNB94n1o4D/we3+qYRubWuyvyY/pUE8dpwz6+iAaairs9sr6XaFpy1ZpUOrqvS+oqYv4oDys
hSt/fzdgx5sGUbGZ5wVF/NnMAtdUWcsfkJ9F8YOyfBuK0KpyjFfP0YhTXN2JZ5BN4Axj0ZVEGqeN
OK+DFWN5vbXNI3QcrJoMNO4StmIWjJMjNexPuEbDDGg9Fy4MOHS2DcHwBygPkaXeIe92PBeYYJL6
ALVp16gvYBndAR+r8ut+xE8NrL4DgkmBxJUeDDYUYa09EKOlgfVACc7fOwyeV1cbcqs8FeWm1S+h
zvLZL8hZEzGBCFqPc+pdkPbA2iw476KFKuR6o1q+IAgnqG8w0HEGb+QkgG+QzAB+qWQTvNuGNxIO
goumH2MZjWVvf+lp9TSRapFKDOJY1+yXwcFjUInV3FeuaN4ZDNBqWSZOJVJV3Y+9usAPp7bAaMGo
rxcPYjTdplIJgIP7Y+RD7MjT88eq8LS9R52Fg8QC7AYnEOdTNP/gwOPBtjNZchLRZXM9h6CtAS1Y
4s289wqsIfFIIfODxNGGs9PtMt2pu1AZEjH+amxLEHbbs1Dpcu0mQ4VVVq6UpTBWdrOjCYw2Cius
ngeQhVKR1MDUOBdUS739TKT9x3XgU3g1j4BSDg9Yv8i3ZPvRU3VPnpEbWDiMbQAzaE2yQgvmM6gy
sLFekmXfIqt55wbHqlH5G650A5qTgtherrVS1xxFN4vqS3DF8XBqMcdHfY5+vo2Qn1zps4lLMzDy
3FqHJZW1bQbAAHB0b0nKG1qsu4+Kj63aEQd4VsiKQ1q0Emfg1j2YaI4/BqvuYx+iJh7ybUOerVPw
dxz07psa7s28JcPBqTjAHNvXZJ8GinY+k6TufUDLeF/BU6QjmL1EfN+xJVxqDwojRO9VJYDPirJ5
6wKEZjP3zkhWoLXycmOQwQ9oz1NMrrVgsMHwlI2tz9bnSQiEeLVJ6Nqkp/N9aDkSaR422knw2f3b
96EXn7XwoC5Kw/Yp2ZvOI3pubU2tHPskmnXQxsPZmtZQGVQE8SNOhT+9NYh++M1OAii+0VyBY8K+
2Qh9P8GAhQZ+WbxXdbBEJoZT3mrGJg1QhqohNBXRcR1IbIm26PymmdBu5bPInOo7QoWQIT8G9jU3
QCdVBwnHOLAkwn4EYelI9xrLbNOA5i/u5UGMhHTFUNSC9sOb+b1yDZM1ChO1QzXqAjphh2rYNjs/
EFITWA2+gw1OUJXd2GkkaKfyHoaNiDyx13ftRYBod+aEa8gU6NQIccSdbxE0gaJ5CNfH4doZ1o29
pQOaPS+R/FhFyKqHOVGX7GhuCboBEU4nwEwY5zse3OiEwLLvKhkisZhBKHfOoPU1R+JAma8Sn54m
3c78QA3GHbkIbya57Tbu/cUMOTi70NzVyo8g/M8xvavSxXqMMoiQgdAjEtABvuL1F9EsUCxUqzaI
LZzuAmFClYx4QYWNmbsXUyBGK8NJaGJ8P35XHFEat4uAlWVL1vU53DhKasTMAeRomt+wcck/AGcs
Emav1biVAbR043fCAtHaIdrYuAuw3JgpY4R4SH4kN6gGVMSvfPVD+Su+iTpQ6yQzn9nDe44bYjRR
ObDRFS6DrJJKat5T32mOPXhaWCw02ZEHyUQfE+okwVI96DyNXjxFfM0umpIS2Z4+J3JfQruV3Om4
PytmFCnV3FvTLbthXxq5SFEvaUAxnc6cb/sorueePlxCPmtGcSv33JbHCf/8ptBPymbASNPfwsVU
x7Ax5EKgYx8OIhCPmT89NayEr680HgsSdvdrIKTVgdbawdk3QxM+UkLVNUxJS58VLi4iqm5BQVkY
zeF604ngqj3/D+gmfCOvazfu0KhOtll1Gpozu56jsUr6Qs5vYYLAsq364H2UtHLuOKQWUocrF80h
mxy5kUw6ecN/wvRgUVXUl/5YoW6fKIoXFsxz0mL60HSofRJW/O/1B7YYHuhPd+4ZXm62UOqAXunb
VfzvO4ONeLi9LxmgBOPpNv94S6Ghhfvp3pgwkIKaVu8KrPfTxUZD+1mze587PoV5Qm5D1QdHU8pH
kpOV/UfVW/O1cfNZ7GUr5m4trsbDp6rxAhtS1nyVMaQCe+5HlgDJQgosbfEkWloUVV21QJu8+iEk
dXz6PCFnr3bTPigZYJQYS8sXZUEyP1C7NK+8jKtkKp4vbA/cRntT/WU4Ll1e+pWGkNufuBLmiHsN
XcjI3ZXYfsVAe1Wvk17l2OipYhP43EoJe9j16eKQTKlW9kvJTAHvnDth9kwZsR4VRmoWtfsMA2Ec
dJcKVumQ0fCDicTrZjHjDAaLqfZGCwaqJeoVEcKbqrvPBLSZO4aIxjHIVkCe2oiqKmelYwX2wUQw
ggjhxI3lUde9NWQEZbBT9efjNWgbKWPGEEft9fobL6Mm6XZx5GfLskFBIaT5vdfRVNzyWLKFX9xc
Fa1RZLc8V31lwokJNbumLqovdMDplo+TMVjmGOMnS7UmiZuQFULxCo762qMQfxeBU3h94Cjnd++J
yZvTlhS019DkMsufZ5RInREGI5eEzyujhEzjZ1hG+lXdwmEf0ICi/HJxN4BF0Zriuv6PfYrHwZg4
IXQ1plF+nj3rKB8ENWWP+UbeD/kC4Lih+V/g1hniP+H7usigXCjWQ+OgwZ7otS/s8KFWS6I7WyhE
xZevBdqwr5w30B765Vv1lZjjb61P+y3uuv1fiH4D/Ba7HLFP/qAExcy9vYXsD/hIQLacDGI0+5+z
vEz5VePWtuNBEuC7I7sVtylod41z/gVUUHxBiKHEhRtJic8917hOJjjhPLlm6tchXfsCYIoXYurP
KD6lSTt3PHaDRvgxPSsVmvWZ+ITRnGNFsGPgJg2PXUqSgAxEomMi+f+Ui9bnXOS1Fsb0kf+TuLo/
tRqk/LtDs1WQFPl3EVBkxJN/h3vM+Fccn9/9JjIzavmXZ19yZ+B1Ocp1RbQptUKw/t8H6PhkORXB
C8ntCF8guL++4m/t8Gbb5yhvXEgVgZBcfyHHU+r3s3F+zcKW83twibFa8FoJmrCITZsvHuYc4Cc4
qhRVHAyjjgHDHKW6852mBVCH1dYg+KzJKliKfegTKgvi5GyuxJuUJ7Ed/ygKuxD9lXSw104vRKh/
In2ih4A/YQDmthQ9CsXRbij9LBiytI6AwQCjBqxsc5aUFJM5daKtEfbO4ea6N8pPsKRWbzT2btwK
4aUXXLKQjEvfWFIaFAMYxQXTR8Qr6Z6F2EE5ZSIDV6h+7DROtgxbis8jJ9vE+o2GJrIWe23c70BP
XzsZh4M8OrdoLaQ55eYspTgYDQRgdHfwm0M/ZyjBC3NJJZDAbifDm0HvfoWpF+BsZYrkbrKQvwj4
PA4MKTRTvAHajrzlbvzJcHmkJRScSlYdev6Bp+RkoVSJdM9kLs1XBlQHL1IvU/RISoKmtqz4fNzE
HEC0PbD8rHqTdZ7S0noKfjFNznd/dF1hJF/SQ43hQw2/apDa3IaUETgB2QZ/3O80TAm26mgfyO4I
IsDnLF2c0Ck0VUrLBWOJw3TJRdY7Bs/+8QdEdSPTDcw/qefgk0l5Ayx9zAv06T1Dcbdx00DroggW
UG9bXXPqoW8KxTOCRLMeDkUKdhuaf0khZ+DZG3nPBy7Be42P413GwVMFIV/1bg/9W5oEQCRZ6m4y
IoL18tj3jBkZNqsMNSpA1UN+jJGx0VK1JopBcSWaVNCEptR8rHqv3COk+f+5gBmyQHPitVtsx5+2
h8V7S3QiSSDHYuil333VW4RD2EQxXh3Fo+MqXzu6k42ZetCjphEuv8jldER3T9TlHiPgCEBSVWqV
G6YZc4S1DAylpmnxlTDP/YoEPjyQdNMb6spVCT4nYzUehIrG68qVbetbQmn8BUInycsTrLtPcahY
d+4xjtbdX3M1eofNs0wEtohoGs0SFZxX4Q/G7udClq/LBmT7ADR2/6moCKDDL/fy9YGQvpnzUK8v
MQDPSeo9fGWc4Wc2KMp6XqChMe5Q5SUgpC18+cBpvs5GFFZEx7i93ayzBtwIveXtlu0APKn0r+4G
Nxvk8LJItnO1xjh62fykeIqC8sMDn6Ig6a5G1dyyxJ1GGlLf6qgEGWfFj+ThmUAcVR0kjasyNHjg
OYBhCZnQBJ3i6qVmY0GRKvPlIT5/rG9/VR+GOfS/kYy3Xl5TLl5Y6Ufl62iTdU4aefV+9wobdCQM
nLVHNG5x2Bts0TYuAW6cPuYiTCXk18Jtx8ibtzxOEKT6BC5aFtPh5lStdYItsm48xf3vFW5RANso
kodDHMF4QhQ4307qvU3QJ/rPddfThHmxoIxmYWCeTGa1H6Zg1uUiR5Y4EkyGz9rS9U53n9ippEQM
44GaM3hGT1iNqZnEDJdzFbNgTZuqRHV9T0NK6F0grISSwkYTMw72x8qeFx7yh9G7rF2bwhPPvX1J
1BZGRQ/6A96Yb4oihBrgdinvlzxSJAbU6Qpqvyfc5WvkKf/4Ysgw4bNTDfNKZ+ibftwTOVRP6qrK
eewBK44/EldG4ffaRG6+qfMzu1f7Xcb36/J53AkLJBPRQCA1l47K3Zb4A+TBvhzubcqqhX/UhHKY
iJ+j5QXAyV6cETooZ+JsXYGMpqfmgjzot2lMXduNN/JqUI4y5fZQIRPkDFGfpGVbvXRTBwOTxDgR
d1auChgMz+d2pC5SKVfA/rlOl+6t8hHqPo+JXfQzos9Ahp3inAgM0Bid+JWgKpAaVfBEnLRm8d2z
cB0+iwwZ1mCx6NwSG1y6JIzRGhfJSj2ipW6r5clKFqZrKXEMa7jCpXZ/2DYZyisuDBnrTtH5RR+/
qztKgvCXeZDUrArdcef/XXbSd5kF0SqxBR9twXkCKqnK6rDbXbblsqwmHgoGFy1VkcVy/01zfsjo
qrfOTBBq8nXJwhsYyxIHSCKeV17FAQMmAdUtLlCK6glnXUAYwokGmko3lXCYZ9DVlIH7N0xcPrBM
NIZtZXwydC8/o/uCvdR+VfMvMOdHQgdf7qPxajbuPAevFePr+N7G/nKgtCGCvQFbGlmBfSpOdKOZ
Mdu5bj2k6ALeC9CMshLLR0FU+WTwqIfRqIZFEfn/xRyr9U92z23LMT/5j3fskGFqnvep63maIRaV
1tDN/cY26kluBPR4main3LVganjywexpW9mvgYmiWXjT5wojPq09t+BpAkmAVaPVnG6e6GQvBbUC
xDWo2Pg8QGmSnWy9EgxigCgDdgDqw3Yp+w4LP14TEi1BzGcTj7H6avqqZO+v8BxfMrsY9bbNHZV4
X4Mm3AMbWw78wScpJeN9R73x4YemGm1KCrs0EVrSd0nTrJUsAmXcpUpNU0y4UF8uhRpiSgyDFBw4
3pT5Wt7Ljrd0HSnBP15xY6bxEbBE2hvstrQbpRG1aAe8qVuoD4uaDVxq9OBJRQsPKeMXX6JOvuBw
S/wG06GGZ7iOE8HJHtUVagJKw8zr5EBODzKScn0S+sAJ0xoya8EczrQYyk9/KzlNJLXO5Ff+jjue
Ze2lOVuIXAR7O24ksUHDde73BeGgEC7a9qX+GWy6XecUuhck9RNeASfnFH7yojbKyHeGSV8afPpM
0N4CIxVK6mkp4LrREFYNRUoviIvPA05yEZ58WSEd712W9NXqIDAFiUtJ7Vj8pPD4D7rFb5vQBl5y
1phFKXh2NoJlZRlrNTPx7hygYpvEblAG0tYuxhmZKz7MPBeuzcbJg6lEWJ7G43DZIl3W+VphwhJx
JCUS8S5wO+Kyu+vbhHWwIs1ZFmmbaJZhCg3woi93pFLTLdtTqe+2JlAGrJ8/+U1Ale5V/j4Udvat
adlHXOpxcPsSu77GFyKCTUZessTG4aZX1RrXTlihcWXZ8bk0h2CLlJGwJfcBXfQtkTB7ardRlKlR
/6qR36G2UatFQK0KDB/LiLc+V0I09SFLvn4V+UkuF+FixYttesQ+1gv48wtuUdSzgGvBbvVVxlcO
jP7LmGmSsO2WTS5jrPmCweGPJh44QcPC6LgsqJz4JHy9TN1zHy+AIHx5Zsf8joKT01+ZOAWnRs5S
22+xjlthGz59IoU9+9oV+YboS+Yjvd94M31RyGT3gfA42jNNIu3X2QY5K4dPC74JCduXzyYp6kBN
qY1T/M1UV92xjC4hZF0YIpRQgmT/6CJR81fkpoPYbxODC+0RV+7SamFbLi3WXwFuLAaaR3GsrKJl
ykLMD5MTXfNzCIsse/OObcMn3c1pUwdH6d0lm4FbBkKSenNilA6sFhZ6hyP3Hwv0TYoxMwvXpJbN
gomjJhvM03zloGojEHRfEFitEGFOwUZajQDJoUKBJ4LvFRwm1i30yoz8fc3094ukxU3UUquTj1Po
OTfbj5WYjjihfFMagm/G0KqiWOwqH9dtXV6oVHHdCx09QjFy+2VDeUws4wDcg6oqOMvcBc+w5bYE
vJPjcDr5/j3+Cc3bYUZpKb6s6rG0YjnPEMmM3D+PMOsBlAP5TirjVMHDcVqEZszEkcYcyI1khqgS
uuKB9S+GyGVAG167yed9lsPWS+UdWhF8eOPXWd/KdsZavcYM4EmWbKHCKm7W7pR7LAWllv4XpFOf
zXiK671QOQZqDCHeFvFqdkCLRhDJnXFD1MAlloB04bTLMhH/Augw4f1AMVg3s1a6MY3dCy1hPLoV
S2iF/e6hsQHVaOws+GD6+WUUiwDIxvhuLXqjdt67rm4qYRcMOXXBzBpx9GTdkTMuicj+b6EM4Ivh
ZBtkJBsEtFTj5AqJYskjFosmzmiGuAgvANkUnNB711zuI7Fzihq3fZvLc3d9Ok34lhpkPG+Endoe
3Iw37maz+J/MzQZqoIWRV8pwA5IMpsb5w/AKCnCIf+S+lz6+K8VK7lWJQEwjhFjkQt8nM2OMtoU1
oQ/9jj5eNLMCeDzzYVUUYmJEu02thzdp6TA36Tq07uf5O26ptvMJXjDGCF8IcUap9HRnbd6gej4S
fnHNT/7DN+swtok78+r0g88+1zTM2n+g6YGXKfjDBFg7lWLbW0Hl4rYDBWVe02mpAtWxqF/BCsu4
CUfTyfZMV48+G1Kydq53DX1vy25ln0BBV9gxvB0l6jR4kJFZxWv4aVxS9DihSWDMpm+Nb5o4Myk+
CQuttxHfU+Va2+0n2ytmwSt+HFfi/qiGK2SeRZwgv8E5w3VY8fUJOAWpPYHaKB6wRoeyzTtoRTmK
dD0TNs6s4dFIMaO9HN+Rp1/2gQIgA8LAl6/NpghAuMxqbYK3ctrv5m+6SnrIYLnwOQas327ZB+Dl
wANuiCLg+fEJjD63zMqzRNz/YLzm7uYncDFfs+lrTmEYsRc2spHdvz+gngdjcLR41TYDmR4LitxJ
dcZZXG6WJc+HPB/hj+yi31jD7xmUJUMZSpPhSDmOstvvtdPxRnCzGDqH/HbEkHySosbmlODq36T8
45SFfjW+GJaspYjnO9T3az0KdmCjsGe09nb7dn9MwYTdGk2Do2fmFLIdpo+ugLI7qiHg0Xd24Q8z
FrQWdiqXafR6+Av2GUZIsbgSspmAIdmRKpiRsYEmRqJySK05yHqfuh6xFvzGItXFZ4JbGAA5GwMt
EGDaW6HKLudnEaUYJlT8PvBunk94WyejJcQZBMCl4SjjOVjOvdh0yoG101rB13KTArRCrEGFSb3V
iNV5AbV6Wj19fuAZ+a2rWS46aCJogk8dte1vSkazMEimWNAlW+SDN4o82ck8C5WkTF8h1AsbOr+j
aaffXSLVOtT1u6I/KyGtXz7m9plDCmn/Rz6dKLNxNNAVzcaJsoCO2Myfax/hgUYSb2V7Y+g1Ekad
hCUuWCcPd6EHMnKPkDo/Y/+P5I1na9ya90O2UboiHWGbT/tWF9lmJv4cQHcchpQaGUilrNBOwxRn
S4sH9VobBynW/z3kQcreI2oq4NqTz9w2F2pJUpM6QcquFQXr1zY7+xhiLMIosZLcKgCfr5zFyx82
52vOhcMkTLUoFr/XDYUSUkWK4nXZkaYnegb2iIityumiVKcJJAaoYwVStzpTFTtv7JrXqgmpornM
pEHnSESQhgbXsMBnh/rQN8K9yP3q07pcmf4RXQ8ICy2DmYs4F2P/Pqs4l7qihNaK8aMq9CXl4Mj/
hOoqsU5ImpEJYCWZNVmedmL99ajRFhK4/vGe85JKCLuc4LaBJKpzaNMo15DAepgnV35yQ2/8fXAt
6ub8P/F6r0fGOEX0MuhAXXq9stZJvdF0YxVj/tzDwoInceVgdOlrzpwkRPpkqUGwJDCBq24CCBxY
3b6jJeBLJoWfcJQYiIxmM6Krm6pXn9R7mvo608/Y/j0az6GHr+hRffTNAEF5TpkrSn7E8jDqApxi
MgFVfmIkIATC8ga6Bm3ErP+feapMVXMU89WA02nxLsuEf7IBJ/0B0UPt+pfI/cLc9JKlhP10L6pB
E5tASi3KjBp9aMOc+jn7LWUVXZhbvhWfn98bMlExbuyh8c0djNhOwGPniCpNAjHLiKgqwVvJCefw
OVGHX8nBNoywAO+8CFM9GDFGWzuSOOZ7ZO8C70ijy9x7sEGZCC/35xZWORyKWEfRNOVf6r2a5jsk
gCdhZGtZu1swG11KG0ZJI8bQ+2ecjocNpELzXhBBWSR65ECodqLKZEpZFJNZQ4ixo5j+B9eH4XOE
EnnH5jiaMnLihEBBuXAC+biMT4PlcRY8ObSloGtdbeI82eCCFP1q3gqOm8W7qBrl+KVupo2QSuHf
fmI1/MHdAd0PEzB/KqTiRGSdbWS7TsQc2dDYU9u4gjpJpHLywwgqo5kV+o/lsqUFSsQgmREP/n9D
TwjVIZEsDyBYqyCZprzHCH73tSUBCLwrj7Ta9FES3jLZ/PmhwJxqR9f+8s03AsqFzajzb4o+h/rQ
uh68M4q9C3sjbYeed3lyMSr1S5GrxqiCRkXXmxQhUhwzSCKgATycxqDRT5X3YjeR+gaUQhblLX/g
YsLxBim7xajF1OlA24ijvVqQycLNksVXktHMqVHZzqP5K9m2Xb9MGSlv7t+xw7Agj5mHUFS456be
SHieD0hywdZN6AsgCpcdKYvZ6GH+cX05kJkj0MzbqpJ71LIOY4O4Y/rjEzPcPOFUmzNU7ZjBMYWe
R1iCz8dkbW/a9MKrcrRHLq/+sEg0KOnSXz6KCRwgN2pCs3m6FiJOfQ2KVseOuwpcNy4g4ZokwblN
aEwtPEHoWFpCCYDwpNCIHzp/1fkH8g1p5+MY3qp1X3Ibu0+w9lJc8NcVYZPIsyh6m+UU8i6GtsYY
Rulj380Sj4jAuvOrMuo+22MeuA6l+1otZ9GfQE/gFOyXype0SbRNd2YiCR5/8Tpu/CEVaSMiAZtm
P/7GUayoy/p5Jfzbu97LDa1VV7fIwak5sZFNgw7vbTteBNUT5QpYtkv5xS6JQugtWiRJLLFBDxd+
eLHlO7KU7FrA/NdKDq4pvT3IcFKfEP5Q0zgOlhTKYQHaWzrz615DHRmBrDoAm+cS9e99YhHsqEXg
HXXiQmzXjY7j3xk+Wuxg6eJum9isw5bWXE2da7sGCWSyoP9RzdW+xgtPaoj0mXl8J8uzG3/fxJfi
nWKnPYA18scTeakMR+OmvWHiMqC+s4DvLBVBDYed/h68SaS3JTCcg6JrPPVFL6qOcoZg3f/7KEbd
aZv+e1kZoDnZe/6jC8IWPl+/Pfr0vhRxxAXiM84K/eiyvl1Kj99akmFn8XTk9iv+Mu/ye1F1snXF
s3eSPNEhkWS2NDh9BbqqrxHXWktuqg+lh/61MdB+CgXgYd09bMtZr+g4aFPIRCY5rILkJttjGG7Z
wheHSulXm7PPIVfgFxRqiNKWneh+bQW497hVRj0P2kBMyEu1/gid1ySbI4wJGK4RBQaEHGTWQONj
OTOGHMIPu2mviMP7n1BExSoFXegmIE+QFuFnwJj1t+6D2GU8JhCcLdQSS1TZ51v7tMp3hYzRTk2A
JMoIrGheZZ8XEscOWmJVZiqpgWw0bqEENhhG7X631JMFxEPip6V0Hi/DG+vM0tIhMhRorrlOlJdA
+Mku2HcyCFOeXFT5e1HYnOtUHjQrncyJJds4l/DLNiwiD0ZsBod2OPr4u5bX3EhCwZm6gUcJITFl
mCmjebCPdp/f89WtK5xjHwNoTKf8AJu0trfLv35XWLjq5wwy6JXX+TTfTgMrpwqza3Sp+ShGhTBT
C5WyqO8M1AMiRzUVEYIyMYflavS7LAC1+FKBFEAXYzYvLsFvIs8K0eOgzYh8gN9b6Ije+0sv6jSQ
XjiKIUhEF5i3VNcGby13Ilq/1tpVV1TCJgNSktmYlhRCHMLLTL8tBN99cIXgjpEtREnJCIkMWQPf
3LUSTKYnU/P2be8Z46EDyoVna9YK7yeg+GnQ1JZx9YtoRB6pWXCPZ4FEU4HqM57YQmM01AxdBsfP
RMVEVutyD5iGhG9/Lcbw8AgBUM6bIWv+8lUuj6S046YXpIugjo2TYzGrhTXEgUKhWxLoxQbuR5xy
GBE2kQdoQqgD7pgpgFR70M2d7xmosb+/MEpdqEVzq/OF3If9FnxfnCSBlkVWgmgQ9csbfYsBJwjD
GCep69idcciQDHPTh4W/9jEK/5EXtyarZrJpcwt2R9r3J97wywMNHxLRcM2fxNboRyTah5Zm4PIk
kAHkyEt5nWAy4B9gsM7Q8F2nrqasJWbUHDJo7repX6e/HioYvDWlZV1ckmoO1R01AZjjLjqP7X5q
gGpd95CoRPcRq86KBjelHyy/TG6CmmFNTWIe8L9gGYZykJylOn7SfpiRLS8JxJQPVkrHGM1NIec5
Zn/O6mKPJzG6qcIBPq+ll2fJKyqU/PJu2Wbv8XdXtJLTtYlet8/Ie3j4GMXjXBKThZeA+OFEERxF
hTR0vNP2e2pyCmhsFcDbysKI0T9CQIKZZ+VZVPGAlUwTrBwxpvBwpCNC/tzRYHQxmxKOUUXpA+uV
JaXuQcnZsYJmEi4bMj53HXJlw64BNbCp+9+MSvtBrhgqCU511LjcNdhb15hr/fdtralwRQ3ZQFTq
EK+Tlyg96okscrqPDaukTG+Wv52vV816lHhFmXDSdXvZothxDDhn9OvKF5s3yzVYEun5Yq7evpm2
tYekN/ER4QM2IlHqGVEJ4d9GQPmwPKWRkU53TDGRKx2b0J88iTOfJqRSWHhJfJAGXg0hu+WAZMFu
lhaMzmmVUGuASUhyKqXg7DXXD5mNROJqRpyzCzJukQ1BcD/mxpd7lRkOQdwQSsaejaOQSM/Ejf8m
inzuhAymbgUkWqRbQgehMmBQKbVtysNHCAZGid2ajIg6oXxvFWcAIzELfyc31ugUsO8Ew8uTvS32
5KXf2jvHarogs9z80XXlrkURSSoJyc7uuezOI4sYYd5ZYsb58ShSvHJV/V36lS1oovXk0BxHs4Y5
LT6JU2Zgl7VHJTGzWkzIygiW0p09PMl2CXiRyu5K8eZfR1rG7fXkvXrsMlEXS/7A1nbTSSw2/EkE
gaahLRgTg4ILGaHYM7Jfgotut/rlZ+/f/Z2ladOeHY47WPx1rBnpp+dwCdgcd8R9aqvq9ao6izAL
bqOF8NTKICEsiBRnawEUzTbeJj+/eUnFs42jQ5qUzv0kiYLab+9JT/Ak7T9s4wMFBoNlD1ms0DiI
Mi2EmHOcp3XvpWa2q/y6NaYcXHXmppq2kdmbytD902IgbF7rOHXgO1zU7Pr+Smo1qFQSFomQl828
ZnCUYY0R4roptSrmmfXyyAPHbgiTeUSWVCvp1II6x1osencvJe0FV/AeimMUqY+3lUOYFsS3GRl6
/jqeUVUE0gEwJ7rcLIiD1jbA6j9b/qScm7o0UUYS2DSvl9+LgfeMA8h5AJeb8YLWSI6//2PV6AP1
7dTqoVHcmJgIj8kkK5ywmEJGz1XjwaG9R2WK65BdXHJJ2CzPEIg7zDFiBwNv5a9askdAwnwIw1Nd
245ikG4jaXLn/EimjA1b94dG+YwQzqrZJuwwOK+HSfHbTktppXuOHs0zZUZcriikKbRVHvrdyGo0
kuCXH4gkR0uUu5tEVPN1mmP9Gl4/QUsI3KILHtQwmqIMuBH8TbSkC+5jzmb68rNfMcEfcEydW2J/
KiUKaIYdXXkuJpjAP77iwHkUwZnKS1ONR+VUFOQb4THbTSvxi9gLVCPfqoJdM1+Zf2SSuOlgCf4u
kHu3wr5wn43BP0hvY/yJr2ScJeBYTV3dDarMPNnC9CzTkSDDa/gv6pznMFFjNj+vJqy3IjfMX71M
B6QmPHLb95+qYfqBd5b+umIiTxpxi1+IQnxKEV9q1npHrE8IUj8BJwuPpRZKb/6O20kNMpiN0742
VlT1JqmG4nVpimKEt+dNFbHYhBYStiOwc5QWThTfVnCkjWvycu+IOKTja5yLZ87lX9Du7hSBuo94
bKywhYwKRCEPFt14RVEMA9s018cmIcaPvsvXsKB4wcWodB01QpcHUqYT1/ErjcvcK/w2K5W4UjU+
NrSDUZUiSvM/ySi9DsYpxjQT56cqhZOSDulXwD6J43ZQcIQ4pj6kVdIMrwAhM0QlHz4x77HUjfxJ
a0Av6aYktkukbN095tRZyx3nLXW3s6DxBY5IHcN9l3MAxPqY0RBDu2lhtzv7EA7MFjF/5tDYqSMv
oylKNUt1qTT7AsjiAxyCAgeTre0M8X2bbOyIRi07BbEsD5JgXTVbYixJmEX785SZRSWwnUZu+J3K
P2qgax5C2O7N8mNIV5Snp/Ba7ZP8YtrcoG+jEcIq9KY5INXc1iOa9Fej2S2yqF0kZ8ysc719V5d+
o1UmnYjO/e31cw6jjOgE7nxRGJ6vm6Y2gj38RKf01iKFMVzG97M5mqfemOb8HyhgKqJvgWX+9zrR
FwPY7iaCor0xsshLOUZXrcGoMfYYaJx8B6EO6xE5geOou2OO41jKs+yeVfMX3mSJxrkmxycmCGNF
yEynapxcBdTrNVao7WDSA1P+4IRRby28Z1JmFY5kP/N/a60L/zl+fdrYgVdxCvw8wICdYf7DwCH5
rhd4xU/eZ0575ABRXSsL25UDQBi9jlENNjp0UTeIZWZqpVRrgExSW4EdX9LrmYIdl9oOE2xFpsBt
wHsU9uUobgKUC8IGU+adV3pnPoEXH28qL+dO1r1M5qBY3Cyv3YqFspdWgxY5AqiTH75aVd4trjoi
yOi4udRuirWGm+R2xPol5yl6+7WCpihnGyndKVSdXmFc3dKE1J0EUPcW4JYmSb9mecv7MRXYDAS2
GElIpsY2X6z7uo+cFnPyvqYD2EgPgOwAFhflUcsaEumttwom/6FjAjr5AZCIpmyvgmzZuzGxI4hD
1Z+B78H9XfcON8FAknR6FMiZAS6j0Qqj8vqs3P+vMIcnrGqEs+SoASfdbPXTDWqMegTFSnKaKH0N
6ZnUDRq/XcYWUyUk6WcES1neQkINPVA7pHoRmeWUYl95gmt3A/lb8XZnslrOvyi154ZyqugSM2KB
U6W35AhvVec5GOesCKGRDitJov4+nnepJED6klI5o9qF3aDHg/Sjl1qkr9b7HAYLEk0CBt8xXgn2
3hywFuyUImxuJQt5Jrd1Ccx+nAS7+l4KcOxK0FVJ3G4eZZrKSSTbVBM05SCidbvpAYUVJUWiuN7f
HH5CtHjbANLLjWdUx56RTkMQlmMBiie6kK6ymiH0XgHGvuEt0udJswQAd0nbFR0ZzreEdpsK2h1h
WVrR8HO/qPU8RhcGjQpXJucvh7zEuugvDtfQGx32WXvKSLc5DUqpV91ICNEgoFx46O5x/PnzX0a0
20riJ03CwMVdq0x3SNpiFZSphOAcXC2YCIpoaBXrSHsro8dfXIKyYYwOrdzEafXlOCdLd58eftYd
JLBuB2UoJFsCm78zFw8YWBa+6QxWV/l2SN7Y29gOcWSaFLGSI5+SFuYmv3oaHogEjwRENOsdTv54
lh2Y3LfDNY4LuYBj90dWl8rVLvyEKie3TnzbyKQHWckquJLsRYlJQh+dp7RKcWzZa+IY3+FbxMHM
OV0AU70mDnk3LImSCwlVFWa4A9FNl3gPgA97UShvZ2dy8ZwOM8itTczzHbi6OWx4Y6N1C6/rZc+r
e9Hh/q/okq7gUb4ZQHQpsv7IgpO3ngf+FCIfWwAWaF1hstJV7ldyFU09q7XAeQNJdX1ixUCEXta4
dyoHAkAxCfgaFGEB/k/2HB4LJhE4Df8TpTJ21ul8xOlY3yhN9wIW7U3yhV61fNEPVsrIghEqGJ7u
NmPWYkQn2H4e010NyBqP7pIXw1LbgFoJQ1p4ULaxO3egdtbrRxKXlVHttjAYpgliyBCmOGBTRvXa
rOr+MFOSXQR0zgdhY1SZwJMg5kKACiW9Ltil1/7ywuG1OMDQKcRgPPMy9EPT2kkmCI0tf/S9gwEQ
FiYVNJCH0xhXzI+NOqIjteh8ajxyUX5wMqgtNFrknCNgZYbUL4CnJNo6t1g/o2/V7Ps6laBEvaQo
HIq24Xa/D0vwJUNlN4dL7DTKwqwbeyNPeEJTcLDRQRnrGjL3q2fInKy7v3EFu6Dk/pfOs719Pc0e
oXTv4GdTKpBGpOKGmpCli8d0D06w0R7Z7KuD18CTPSjH5gFFtC8S4cG5b9RX9cHnhwOMqrXhOWqI
KYAzTQMTNHfOKWd9yXJ0NV3lI7OE3x0KV14318gzZB2Rue6icbZI4TYR666pfgm9RLYdXzvpssVF
2SWu1vMOBqTNdUbW7F9poDw6F3AtvjveE2ldehCEydGAUFHfQs6GI3fNlc992ZAnh9Y2/DTknaMi
3z2AnV4oz7ThCWOHgfwY3bTAqyLjaMOAJhE17C48Ck21KerQBkDYOm7pe+1nYHI5Q0wKTXh+CAHV
iM8Acr5j61Z8QHI0c+o9KCbmELDOXQIWacadTvvxRVBpkc0PEcEXLRo8T+axIoLRlGNovKipFDZI
Rs7cKQcHf4VJ+mdFlnrLjnOmFWZJyhtjHUuab6joHNqQBB8h0dWNk/wIKB0b6i6fWsGSBrfnlAvj
3zo089+aCqGkpV+HSELOJqs0S5Bde9uMe5stwWbho4EFWT09MJQN84FMmBmvpUihYNBsDnr61v2S
oapzv2FZ61Okr+k3wrND23W9AGRxI1HL1O4KU3DMurQMjYwXdzB71eVVtXZWTqpz001/M0gkHfdA
lSNbjay/vI+aTUdVWzfam17mxAGv0R7C4olAdW5AuOVhc+9AKnW8gJaXwoOPAecipjV+MpQ1+QUi
tofC+lN1dP8DrkHmrWypqix+vNsD9FPXJxC8LmwFzbXuN9YgUf2aaWRgFfU/3PrVLlW6WldcKmMd
iSS3Oz9qa8z4d/kmZGLnJplewE06zAssCcK497Ko9UqmcZcpTnWla8zwkcexmHWm8jZm9GqbWNX/
43LnnVrjGXcXGBKNfId8iVcQq7GJNSJAwnWBdXhpEdqDYeglWZ9sZT+MLUk2Xw6kS7ZX9IH5E6Zc
S/0LNvkzmabWsBzXNMC43FMo4tCMAfBHa3ZvkUNDen/IM3GCCfuzxFnyOyveAmI9rxLPDuSFbQoa
uLkDkwUrrisSVZ87bzBD+T5eoOu4x0XwDXUS6dk7+RP/ss5bvBZfwMp4Z4CP/iDDtrMeFMnjH7YS
YW2SP6RrkFmf8zqEYvgCgJYhtBBAz58njDKcZIXfmqacgcsVOXrf25KgrZ2TyBLoWk+797xeXOFi
vELaxHtdoeja+jk94zCVmKtC+LpSPwoyMYyJ9Ib4NyxhVcKec4T4eYN5s6GZ/5vvFvRIIo3GNGvp
pnxleQwR8Wf3nfVhxvnw5+nuIOU5vJtTrXa5ymkOla4jJQ8FgXa7G/c5wdI2vHWcEoiK9GQF3mBi
FOGhjygESdNuzAFBQP/0YHdPhYKZ6GMcKfgXy4e5koqHFNl6b40f7C7GDtamHNM8c9Bbb/Yi4pbk
XX8fsqGLI4G/7W6EIT1shCNTevAnVg2/MWu0RUSjAkpHAXR35uXdjb/UJxdpMumMUs2fJ7eW2XXq
U3c+Dou2fd6DESdF/XHvnxuI1efthqDYXvH6loS1O4WbSAN8E/CxTCBYSSPUcPXgRCXLUqYvjJgk
LD4uOu64FQ0FT1zUofy0PM5jLgRDqt26zp59NyLB8NOHAGoamf3Rawwc5QLxnW0KTold5Ds989OC
pf1kCzXtOJP9bLjBKAck/jUykYm5UIUNl46L7hkz+nkhwWAGHjgJXAreSIhS0phhelaQtRjcAU+0
cInJaGa2WV4l/mFXuzsnB/kP98W5YHuadLj2yoDdF9G1WYsXb8R3rk63/v94tDjM9+k6+boYa+gE
qT0vdtG+w+Jq2XEpZSfXakd9vunVxutPMZKD0BedleO5qr+CaZA1GuTb0LL/1XwEsFQQLnFLziO+
wruSHb2Y6ErGyuVoO6KOM5bpl0xjHdSIw2Zl3rLUOKeiKBR0jIWTA20ZJvFGBQ72Ti1G5IxCG/u1
hx/6J135vSGfm2Zi9VNClBUlhPGoaJ6n7gZUMIqVX6kkIsH/ZwnEnr3qKYNaR1Ddct53Xl7d1Ywb
vRXLLUHB2acHQhALzuus1SdTVc8Yh8C+7i73XRiaMgBR/YPom2cBBRwTc2SG/fX1Rcmzc6pmJR/r
G4mmftQB+aBhtdzlXrL+OH+riyVcZvXUX19ypoGOZwo/Dplfn9W7oWr9IGn+Z8g4cH9jRGrSLaaZ
JO/dt3yrGbCFiowK+wzixXXAbIV8gmlXlUlyHwH29oBuOmuNhMfmcJQuQy6H8Z0yjnkIdzeTMgbk
ky98N8xU+ugBQ0IYNosfTt8iqoIljNOM26MUG1Amn+uGf9BhA9HPm+8zTrCWfBeLK4AcnBKAmR1N
jSrmsjYZ/EJ8sRA03LBpGeVPZnbiXSUnY+K1fDKhlPy1qjZzjaryly9M53Uv1PZjW7pHiJp5F+2Y
VC/A3EITQidyoH5Sg1c6KZ2ZwxuZw9uuCn/lBKyYG9HWCgCAB9Mz1MhqXoFFhPcDnXHEY/j5skq3
HvbB6NWD9hm3Z/aBLslO0z5mqbINrwODdksxAgdubqyfYGpwK4nXHwj2RsCrHF2P41+QU8zNcT0e
j9m7s3g6FfZyLtdn6mAhEr6Kq1ATJnFQYmlgsaxvfEbpgHp3d4SQLellMaSsI2vL1zpbw2Oucxyr
of29wYHLzh41g9a+FkSVMfPqP5kmg3Z5WBXr3KUCtHa1H9M68R7aiAAX6qxg6HR0p0iNYYaXFp1I
IxvLOKofn6rrwMVFxzRL5E31qtK4YtrCx5v5UWbY7deMXanHTAyDA3yj3JH+cMK22qLlMOX+CA1p
72ZowPw54yBy27XrPYAjtBwk0xqFenZGB+JekEQQHhWoVz+9HHP1tJZoh/03hVOr8tmom9iqpzam
8FrSUUNhmL55kBvl3Ps0u/qgaktC2KzuixnlmhIhDb0GM5q0jW2McZ62E0OSPJbLmOVwVgUWshxP
NJTMWk6v/r3zTkM8Og4Q57ogyvylo3+Vg7FrzfoqxgSzarAnw9M9sURVUV8j2as3/olVzymfpJGy
2JNVDhQ8kHr1/go5J/2y1O5ZnDkC2SEOstUjfbd1uoM84S+PpST3FmxIAm8qJkwAWssU4M7W5cto
A95egaGxhd8iXPuuoiAtcyWxTlWZj3QrxMs172/6WDZCnOK1dLFiDll2j8tUlY2a6QUq48zV1k0U
3mEJPHVWliL8BTba/cvmySJjuoJtTkK56lEDdSi1Qh3hZWdBJU6oI4vq3jC5dmWsgx40rASAkNHa
RpbMo6e/DOlT55Y84k2wai3bAeJDaLG97tov19mMmTFXCL59VfvF7oAU8iWWUu5z1FfGWGX10rM8
HOyk+d+S/0hzKG4MOkgIy4KP5D02WDbk6WtHxqFknY70F1jBCHMOYCuPapTPfdhCCiOQV2mXoPOI
QmKiFYTMMUXuIfeCDB068hbU5q0OSXDjBF1pCT6JYSB+SxbPk6cWe4X4PIDOsqD89+avpUY3TLo1
OhP1aogtxycBPY21dv9DHs3ntWCJXyXvFNsoTr9whFrRbDth2IjGYB0X9+6YRr6usBE+zx/4d9w6
Bk4nfaSBLv0QA+Tp2JrW5Vo66XDeUFQ17byQ+rBHJTQ98T44HH9PaXzl835+7UR8SxeF9deElrw7
/JssL9vFyXR0XrJCXWn+GNxdyy/cvIdImy1p9m/YimlqjGdHgAjSGabKY0Rjc1GqqtbXz2KihiNP
dKhXBSFrlgco6AUeaBO6O4yeFGgnSi9JQvzwpzdbt4u9GI2t9q/nLeO6VDMb7jdigHwwuDCY5MbD
BSm8jwcy5T6K1VIZny93PnFka+y6k/B2Z00lcku59Rlx2GjM6ZxeX1M06XquWJoGR1cKfUDj4YWp
0UoeYBYhFycqgo05afYtamMiA+rTxpf2epvfP4Rd8YE2NgwRmqTS6wdRVJ6Z52hhF3+T9C7h4crD
1SZUlBTRB09PvtM3k5GSI6ZrGOw5avAlmoi7atc78z57Bo3HugyAZkqGkGN0Z/sytB0WNg8NE3n8
LzeSJW+DIObgWk37ez6LtkzRmAIXlGWEYGPEG46UTxN/XsfuhILypj9sdCNtMpw1qXK2OQypZTIg
ofdYcjQXnsLXozQzTvZzKSeECdMaCt4S8QpQS87DsVArHZO5jeiW3IzGibTCrgUt6CWhLJDvPM5o
L/K1+KfQokEZsSWUU97a+vlx8C6IjLmY3f0QVbdxqBS6KYUMzR8TMNXPgs/ugtxFFEbt3i1B5AAl
C/K5crj1bWa+OpfJ4gkprYSX83weI3hZB7s7UPqCsVmyAWTKG3PfSl6k2+4Ulvr4CKDNXklixZzE
kituKKCyiuzzrsE/TXeHX3gZKfthZLpeWbDduE2ZLXAydWaCo887U5+D7iBN67uwMmZdDN5ZgilB
SFe6GJpfUbuaHcoTa1IdsVBQfFfpBP8J4fdpLmhmkGvxsI9kmwP/XJDxpdQmrY0r7TtMNhg/wxHm
DOSRQAKBi0tGODLBMVEZLuVr4PGHLogK2bdnYhxMcWKTp/7e8A0WH+yscvh0b2GFwhArN/dV8QC1
zGV2SQB+TsyZ8aaEye1wf6WBJQDcJhFdhYoBSlopO/SdGa5ddUKh2CiWkEyai9njcqYbrjxPqazR
CupLH8VsdKy5oo3xkYyYYyEeWh9nDlcSi0SE7k1FZ/kz7mlP6d6W5/1mFdZzb3UoET2hq9UtnfHR
+OlReJsoow0S+UXOmL053MvMXJT9wwBqp/rvTTWnXb8bbqSO+4fpwBCxfEzYpW5L6IxxLGtQyfkB
dVgw1fTZarlgsRx8EqdnHxJ5aGOekVeMxSfZNrLN/OzpTtpxdduE49Wm2+ApblnB/Lj663jMNjBe
9ie8FbF+gJV0V+qtN0uNXoKnIXEUK6PYQsrsfBW8RhFytx37GovQa/0im7dtxxBo02jCGMK8mxhQ
9jeQv5EIez5Srllgai/xMSQamhLpctAjkDiJki0dotTT4oERO0E91DKYKY219RNz2JR+AtF0suEr
RSU/1oraA5UvjuV1FeCxP88DGLR9uh4nCTZ905Yw3OkHOgonii443GGhM73xkgZA6wfIgLnBnC2b
U1DKemcq4cJDTr2S1Th2vCUSbe0LQHKTY3o1CsiLq06u8NxRFry55EL2rIvSfeWBlVHJJvsjDPiv
ttV5qhtongWin/ZTitSPQjhIo6lj93T3v2kmGr7/NQptpXd1XaVGogu9cGcP0/QocJ45U8wncRTG
0xNgsSCwKR69XNzS/piP93ozqDyGaePSdixrBViyQIZ5c9xyNhzJEE3fYmcKzsLwXeacnyIHCobz
ah0hY2T1aVj6nO6OhLdX/hdTdQVO/Q9Ehgaa0tkMraUK6fKMG5cdNU8HoA9VtHPVNyYrjTipSSBR
16JdjASL/qnVHTt3Wt0/g02gpJWsP8HfpNdmoNiDftN8eVVdM9Z8JauCNje3hDI4PcV8agMBmfs4
SFPj8oPngahkm6V51lvtebKKSsyr411w6d/E/TF1U1OuU88N7kwxui3702UhEWKXDYAbtwBuVXr8
SkX9iFyz2ubiGmsv1BV84Jtd2goAaFj4mIgj9uCdd0gxs1ECjinFQvHuFb4e+PYlcLAmNtnZwaSX
PppZJx32g4JQKABRaRsdDiIMpX85xwh3PcPQCow4k3CkjJuqLQioauQ0WuDTZnkr1KuAkxMtVGDy
2SiY2iWITvBvbz5Eb9XEv8RWKViFT06xo9Je5A4v4V/5pJsTcZ2GqizagbbILFnskKnMoENWsq7j
pTNHthsDX9m+DdRAW3ACzvjO3cajEVCZYqAz70LCHI35UBtg/CWg9NA6O7rkP6QHSlE6lJROkwcQ
icxeJk/PoIxumiECxetV9/DV8HW1hVELEHywTTKnjpTgTI5BJTUArPKZGpXP3vyPoaP85+rTSU/Z
wHa9i30r/FSrpf6bJYSiHL7dm4HMUsvlIqiKZOxfxqMUjb/WHiH3tA7ZUcSMLthe6EOhZ972fLgY
WHWCVtezPu72atNzzJvrsjh8LrQFhqGNllxhCd8HM6roEn+c74Q12TYMVM/kPZ/hMFCokZWZkFpf
EVjzUuF5UW5TWLW7wu2n0vatFIcxCIdIXqTHLoR9gE+R12avbiA9m0Ocjw/HbiBE8fQBbKP2HNuZ
avcHvBFaMegh1wFlzDX3uJF2zS9GJKtk9DUfAMfzw9ht3WFMqDSTS3iIlw+bZPG/8JX2mVjEonnM
1HwZ24/b0KsA/dGVJZljmc2ekk7JF2oPjAY/+JNVBSgJIltmDq1bAF2a1KHrzIYGim5y1CyNa8y3
8lNSfy2G0obfKs8rntjgHaCM1HMB2saOjgRpa+xVd+BPTulnR6uPj6yFJMXtk9jW2w7XHvHyZmtC
T3drbNIBdskeBCPRPPCghS+n6OxjmhyxrWjBCW/sg0qvI5D9jg9+5Ay9S7k3ZOynMBqmq1JXVTX4
o+BMURBR8Rus7idIFfjiGc4D+4UR7G2mQ9M8gt3zIUY9b0KXCx5ZgIMPynZi+QolpDQTgoWFuneR
nNvZH7pORIsxBbqlOPZQmKNZgxEuKgLmaKaRkjbihm84y695xNCJCprLnft+OHkSPr4IonCnJkcR
bdhdSB1kRHBhGdGdWSUARRAVg12n41nPmKzQso0FM1U7Waw0pH4i0wgbdQbwvwOG1CmwgRk0GzVe
M2WLEUIcnrd6+0NRmreEM8gjcPlnM4De4E0LlU3f35LvkWZeYuB9xxWYWKugHZ7cnJXaAMzgePBp
7hT2AYtBpRzCiuIs0piUKDqksGLEELgtEc39krL0VLnya3Qxs1AUKDV3btZcoMyLir4uS0o6IZIR
HpY6U+W0C/Wt+ecZlN4zPCAXkcsNnNm/z/8wPBztJD3RE+HM0RG2m98mNL777kX7pzYH65YFQqBT
MLAzppQvoTxCBZw8BexUXdCZfsceG9gsJp4NZRfMRKyxLWtQSw91u+L/wFa6eDqXfTb2aI3i1Ew6
Evx72aM2h9smotAm4mzKgZZT+trki8RO+S73jZZdxAzJNOrEcyagcGUrbmcXFGA9I8ILI6zRKfCT
d7OAV61eHzzJO5wMCi7HcmesCS0Wvx169BL4uGgYdRP/u8j3dPmx1qQ5nMP1SkUZyHN4pmyHOcvs
/+zI0TYfXnjeCPsY0JrPCH0RX1JXcA5RAZ+4uXYtjaAv5v2Aq05+4SvtbuA5x+vEW4DNEMDD+Y/n
LC1+EpXHTWUCAnZvcXx0D7xHwPOZoBeMiNe6RzibpkManwL1ozgogzDNg0mUwKvj6lnqmRIPXOmg
MDFbdti3W9jh/ViLSx4KvJ+Ut4+t9hoehQpZooEgdW80XEeU4CW4AS0fkOOPz98CqWo8fcSonj4Y
rkhkNCH/wCCiAjSJ+bX6ywAYYeFAfB8cVqKbg222YoKG/JK5iQ2dc0X38Vb1r2twGCH0yEO3kCiF
JRNa2indF8C8ILhtLBmTK3ROC++W6Kq9O4lg/921xYAby2zra1fzZZW3YW0t4lCOMvorurKxPHCA
o64DtbwyLL8JNFQejMh/xKuZ1+33XSrGL8tk/F0yldoqGmp/OhC7nRppaV7r/9zOpEGFSSHehA6z
mJ3KXreJvcB9DTRjpdZBB2c0kWKKaPwD2USANZGzdnbeiLGYwplYVWogjg8+2m4aJbNqYDFhqI8z
m9JIWsm8KYlfRB3EZtjglqrq47dh9/XPXKDhRqv/GylpoHwGCCHfaOyQwylSNPwXFYwePKF5uwAe
OBhQRAeCNtaS1Tr/zRfNMUfoXg8YLaH8HVfYlFaxdmkOBe56Ozxi/rcj375HG8eey4LbTyqdzkfu
rCj8g3OsXX8tu13EFNtW4nryPMgRuo/Z8Ii3JGkIsP+Zce15tkCkaFX6PFfxsvd32NyOR7fE216M
j59ayHdAd8vDFpHjDaZhCStRmyv9mvNLM0mHbqElVwlqHuo3kbn24cqoM38U1GJLhm8O5KsP/XXi
e/Zs/tLixQzA+Xt9w6XOoTlyCCudkr7efKHxmdLhSc2ta1mBoXpFbZUElVi0JQdBC0LiiYsj7+rd
RpSct8gkPB78SvryN3gcWcNcc02empK/2RrJFsBoFJZ9hkX/fyJwnS0R9htrT6SPH/oHe8wwvEKx
QW4b2uo2zHti0dJwTEJXpy7OGuU3sQNJotC4htGdNG0OORn9iqsVbD5VNHE74sBfVVMwSYdTKFpX
lDma4MkfoYSh9ZeqR2LgaS74nrbqWxgnZhqSPfafrzdKg/v0dDFSle4HkwC+PEEt4X1Vn/lyTcAn
b4f2vGMhnUQW6YldsNlSiGhr++fXs2v+140TORH5HaNFPCez8VM/Fyg5Lj6gcOz1G1j7nB46/1EP
tutMGxqxF/mT+GA1Te3PM1aKD37614EQTlv6beWpI4h/uJeEMpvKhREjJ/scZoJOdF25kFebR/bu
K1AkXzp+1S7AJUxg0GSvTGdyCIksOmAAtu0kbyUwCLWTUwRDWmQiGL8X/3WlJyAipGxPdoFb0sdC
j9Y2GM8YHnV3GrhVjMH1ICgeq7pfAkURnyDuF5ukf/8FHkuiPSK+M0XID4tnccq2zcQityQJb5+b
6zILfMDYVI5KZVSwr3HJrqZVK3frGjIMyeVoFLHb72mmuQRbqPmnNRff4/4Us/2nRRQvvRrkOxvo
MV18+3WdBrwtu7BZkWe9o6wtKiJ6oe1LHstsxcnnjm9RmlkZh51nEkHrWTDtHgpQYyU+wSr8JrY6
2OahmBndMBMBfccQaTBh5gbjMyalFvLylupgpWDa4QfnO4KpzpFUkqvWCav9fCRMtKyNnbCV3Wgv
KE6wpm92bmpA1Gxa/s6gaNFhqtL8p7nViZBFqJVOKO1D7rTbQWOLtuQUWrEU8pfOlAdhRe4AfVmx
7578GJy2EoXrG1/FcdjmHLGIehPA3d5ildy5gYMVp2WXaxBEdfO7aXm+OAeyHcOnzPUabWMwIKKp
w6KbTV+jkNVZ5+ZsPqtiGuIe2rkIQvrjciXiStkgyoDRHG2XukSK/AxyecFXsAHGeu1GPn5BGbln
VgjE33isDO4zSm4xAXk4Og71gSFdoFazUyk5W/ZV4xoGHbQKRgkNel9pwZGKj3QDGMM/tvK76yFT
zjGlQ7yb190eFM/lN84vgot/VLbTRkX2P/tFEX+rdEbTyeQVgLCVXETmyrwynqkFgrzbdHGg4wD1
HT7nFM1XkMG4GvyMuoBnyrYttPb7f5MvX0ZHJrwpmr/WUt5gUsR6HuC2wR2fMmqG4GfvKBy6cSlY
PNPdselYH+7pHvF7KbTRP9RAc739tq02KWxtt1Ze4O9S8JZRU4FHjoC+qNOU4UQ4sUod4+NCDOTY
Bv9PNn/Vw0ghtlOZyRekpZpFvWfRBegm/sTnjfOzxeH4E28/AT+KlMHagbz4zIjS9XvoSmkLvOgc
ZqeswtjW4YT20ulWB0ORUTz+q1/FpvgEPeQaApt3g0Hx9FR/eWGQPFbNurMOodcSK2oe9rC7Q78H
OVlzPH2K6JYDBweJB+pZMGnKMhwQT5PaaPlTpWmp5TyiaN+sl8T74bVw+myd6rDm/YEUdXDGqzoA
cth30GNqWkhCX00jappnBJV7902sBVbc+KBGKgFkTdKkbYCzfTNMMGsYzXzU1TD/gGa3LNR4JtN1
NYEY1LXOLpBAcAL6B1e/cWiHe3Y8WUjLgb/qC23Py4ukG2g2jlqgGU6XoQIlh6teoS4erKGZ61Nv
gAEqWx/IhweBRd8ORergRbr1e87y4OMR7KxmlxBYV7u1u6YRKryEDf9MZez7oleKutnpu24Idyfl
h8sZyIuPS8pG56RxodKeKPu+27344KypJXI4BdW9UiYJMaRoJXdG0j8Vh5tPMxkr2N35Fdxu0elQ
fClNHSYzO6xb5a3Dl6D9zeihEhHKMaEtcPucqtkyN2OuF/CWJPBs9PsQvRtSFDF3ahWHsBJuEpDV
zC5up1Evp7FMx22EIOU6je/qcEw9tmP8afDB0CD7C0nYPIUHv8pOaYgu5A0Re1g/ExpujvZKSTsP
MSvSSIaHeyCsJZIzyiuGiXkxy23/jy3Pq8AHHLGt51z7TKq/nN+kZwhJefvCaya4ikENfhsWaoui
k8nKAdM8G0Z8cHbrlEfxskQaE47Df+RtH0PIsLW+1C+vraY+62aG1ttUmUm4v21BRh51elacSOol
6FKGjdlw+TVrcUbDzeuRDbdWGarGVhzXJAsVaVM0nMOSIGm6OUY5skmm7hTj4Iq15DvLk2tw6nzr
VZ+WQ9MNnCkddsnT5q2IGzNHHpuFAJzgfiqj3RjqJ/yeKCgx+9Qre1iGkn3HxrZNVYW/3LzjCWGV
tBfoU+j5uKcXfsMB77qdnLri5r4LB4b/TN75UAyosMKfmgwasQ8Ilb4XdeLsEMOuRCO+ExlfmAXD
YeDouPPniXn/G7tUiBdr7m7aXN0ZHAsECXgN1312TieLQNYngEHq3XlDMs1WnQGN4nyVK6P/Thzm
Hl4AkbE78WYBG77MU5THsm/H6H8fMpEticGYIgc7GugJT3dRiRh1NciNMitumatjzA6SNeD1TRtG
LWu+sBFdR8TNmWPaVRMn22XwzhucOr6iu5nSnYG/52p5YRxSsjKIM67R1Afd1yyTrYr6bOfYhAhQ
e9NRDfQT5hOFTJ3zxTZVAvDaP5b/ZolCzEJomoiFUSSr7806Qzu1sNzdP+i+7b/Fok5mIWRILmFR
ABmALNEWy5GzAa+sn4p0waUETEbT/iK2KWF98zQE67xebV4id9rTgdXXe8upBISs5DE+T7yHYBaZ
dBtFrwybN2atAYB+cZLFgXpR9W5AvnbBec/EYZGaAMLnWL1s6tQKGQllSJgky94eye1wNNeqchLx
d26oDOP4SGIWjuNpJRLbomU/TjHcu3pDwIptf0H7vQAFGFJbx45IhVMJZEmG+3NzmkXM5GCuF1ti
uanz/3uq4c+erBw1WRTrgcfKU5eTa+6OEIHi0OfFgj7boW1DxrksGAzrNL29RBe3IW8xCju6mJzb
cIe7V01BxR0i8sdoMd2AnbNycsAg24ajgfxzPkZ1/Jy/D8WL4hQxHOtNfJFPybKnJ+PRVkhC40LD
L7oP0xXknd8vY1zV2bsD0PEDbw8BYiNCuTC8HPGVJj+c9A5SynfwXjP6xn2SoIJuNPW60sBK6JJm
xmmF3D4ZI6e0m/TWKPrqjEYUpysuEg4zHoiWSQlkr7p5adhltxpC1cvpjq8Z0fIIRGFbBaqlOp4I
zxiGI/shJ0Y5boQAZaoD/pptIzcE7iCvxy/qrh5NQaSYQHjEW12xVL+44CiuSq2SoyRZ6XMEcQfT
a4qmT5jmzcW6txC7+93sH3ewN3inGCtwrQx3t8pF89xhDl3E3eKlQHfnPQt07a889GramOe1/7V1
b7utxQ8454yuYPECJC9T50FL15P29P/AGFTbtDVD2LqEdvMVLCo3tQNIGGDvKuvMNZ6fSNwkVbrK
DByN+6wZYbvGtNtzLPaCEYxfAeXNKGjqVwnPj3DryzfKvwFjVCdKZd0WiQt/Aj+HdJsgACKM0jME
zdeWDSKaus/bQEe7dEZYWQtKRbboV1DPnSMfbtsyMSBnpth8oTf0D+0mHxdaqjjR8MvL46SEGwVt
w1kuXfsW7EeF/986cwMkth5NDMzl1N1v4AYFLGpkVi8OdlVlRWF3BIGyPzFcQGiUnA7yA3iMJfVs
lTod3iVmiaYuptwXTDeOcRNB/3MVDTF7JICF7e2Wn9Fo4Xari2nQDAfHgvmxV+7MLbvR0UJMhQqQ
94GwW4PDdmEY1S4GsQbdNf/dVP8yDailG1ec+fG0xS4dRtIF7PYNlqzA3yysl5MASbkHk269c142
1NiQRZtdPejwpMnYY4SA+eC2OIcXBMVceJEqDRK/W2z0rkRi1VIsjdtLYJF/GUJxd7Q6LuVRMpYd
VRUot8vQpBwMjJIxSBBM6qlC417ytk8mLEPnhrsD/3j8AvO7LX+unukEKo55c/kTN7sfivD+erok
Zn4QkDikov4zc++A0lr548NTiGjmP6s6iAb2Yig17Sy23/IRNTIDbsyqcr/WFesRa84d/sMvFSMN
INX+u+mIWKPOP3mF2mfAYfkxddPt3QmRbZiHNfGzi1zRIj8dqZ1xWtb7yaG4clueP7LRT3l5icE3
gDzNBqdva9HPTXENuB61C0eStQgChti3LK+0+jDMlcjXUNuNcaeME/UTz91hs7fSIdWBsJ30nuMd
9HnPpnp5O7rzLGa+JT12A/7OkXbNOMKlUYp3AkLkb2P4l+Bb3U6J3gRIt06E8r0e+swcJV3utNqo
Narua1kjram3Kq4UILvhPuFt13LM/FYJEihbNXYH58tMWRiE0t74n6zbNAJIo9JbyT2EyawtS120
Zg9IDDiiTAW2AJeiYFAfwO7WvwUioCbDElt9kRWlK5/87U1e4xfEk8fxESx3Y8RtsRITPI8RiIQl
l8p13Gt+ayijDocc+lOIV1kfh2iK5u60NhTSb30HCSjJ/EPywKfBbz4YXc7KxnwCQmZUg5gghNph
OVOS7SitPeCyBfmQX9n/FsvaJSTa9FHubxJjTmharQaHFC1m96D+aakb6D/g7+l8zINNxrM26zUD
1zUa0xsLBetj/F8z9EbRzZr1HFCPekr/gqVN4cw5K+Bvg/vI6lv+73iYsAOabSq9Hj5PpqKzbPUZ
4PsDryaB41S15MKn0B3VBAjdZbnjLbRLGaXPIt3ys4qMqbhU9o8eEZ7Ae1zNPuMK0zWQyY8pldKW
BjIrmXiXkb6GH9hVDuaFRMAKh+u36qv8zuADqPEosCE3QLmMgYywlZE3tfTHeLOyqTN7zp1s8A5P
7vA6k9Y13LxC0SHHRjcpfC4Dmt3dK70KqKo0/gm9VP6E0nLj3BBvx2JpIeuDRbK9A/goJx3LPToc
N3yfk+73b+LuvMhmgF+AzBHIre0CfBx4kPKxmuY88zYW3/Pi9HwqAvgeardBbx7QbudQ31hdEnAl
t34eeTzYXPq0JBxSVqopQcYtxfxJeHH3p5uPGTR1HKt1hZlniFbp4RCvccVXaSetaivoahnIuFXo
M3150L9/d2erj6LcTczuXsz+4KL+RAJlQ0yS8i73aQSJ3vPIryGxRtpfpiiCHZflsRAUnspTQwUu
kxYV2jN7z0Nr5+Jh4tqWHWF2khrG9Ywn7sZbAc+CJqOvqM4+1G0ZIE9H+WXbBepSP4CXbgU+29Ji
vwUJUMuBEBNMIEJXYJ/Cmd8/aSB1E0D4YwNozY7Ho0SndEgzMJJcfnWA6OOOi4ajWv2N2RvPy3U7
vOSMEahJUo6+f5ESB2YNTN6vRgo2JwoG98FOm0m8og0EhUnwjjdFqo+tV9E94JW2yHDVQdxoPFpX
yzScwPUui82lI6zc9EyubHXVTaXLzv4sRWMcIjt+Ar7ksEMXZZeQLK7zbUKdiftXhq/FFt0O2QXM
Y8HDfRcYhyqCqymVjM70sawFlSQzKOv7YYVEA7dg+t1yIK7jL2XxlWF6iaklCf6mAeVwBc09S+/2
OiVBVWmBdVRopYz/ij9UBLmJtwc76djQURcdoX7nKF6JNQcc5h+GwLVR7drT5s6znvWC7ZYDGOfD
aC1UwS8cjW+pyrpAExURAK0imc9N9qnKXiCDE/GbJV+n6u5jz6wDr2R6+e1ePthV7qTSXSnBvjci
1+LuzsmrADoU3zaW5HjsQD4w8dcy9RdtcOuaku3Q3FE4NGBP0/2uumWEyGSSbF1SZHK3dmBTAyLl
L3DFgGEBW5Zpm70lopp4bxbjP71Z2bBPtibYpudCsRGV7FlZpcqvmZH3KqPK7J8jCBJMHDLofYtw
U3iNUiYlOTGndBVI4710wROXZqjS63jYfF5Ebc1AI5G2ZOLDsvtQu91Yeon9CIMFEVUzrCna/hOP
1saUwEc6ez3LGikvkQnLPoj224A46sbfiXfN44gD+Y4Ejlpmrlb3u5KrvhHNCo6Exx+b+UDa5xpg
/GT4u3l8TXd9XUG4Qls6KHHatUhIvvryvGBiVOgGlb9F4w+rZ4V5+xWunWOa22p0oUlMNZ+jJUow
kvnMPTonxPbWUYwzl4Ex6kMgFGVT7Z/2w2lfCSO/vEDOgFVWK7YEr+nnOXWHzHBUp/N7YmdIA1yn
sx7FMef1fcsETsof+H6JtFu/ctVuH1VKD1XXsk8jirLYKJXXfr9Ww/1rTkyYuTk1G8MJmOrrygaP
xtq6cRCOXQxkmPk3XLPj0+f0XFD71s5hJtlvpa4SOkRVKe93h1fvfStoY+WNc0L9qNg4y2F04/pB
5OKDHK5Qdczh/MKyg1IA6XDq5v0xMXdCIs1UklHvhq+dNDOEa4uGl2wEMVdRbkVHO90GsmCRpnBU
AQz2YysFYk35XsXCx7UCA1FoIN7X06H0D9IMKEHf1hi8nybbe9JEe5SgW3+Og7xjNHiSqix3Bp1o
Vq8SOu5p4OUJySKY45phYzjzjb0oCDUC0Fsn0J5ZwZVKXhYUfV91NAYNSCoi6GaTGfkvQ6030Cep
QE56SpQBvf9GtlYwcyoijMcapxMeD+ieybrzeIgmbSKJ3I00fYztF7IpKaPl+Gs5cjuxt7IUcDH7
hzQrorr31qfTA5LCd7uLNQLQxYX0fH/Y8AfafjUHAnM3XE2jNrA+FX9d/hoXuGb+C7GFrvLPn7R6
XFqZIiUTfXWSt/rK32BrY2DFPJKtC3j+Ikz2uoQdQRWrooAUcEtiwbzIQgfA5yiQukBnjMQdONhP
T+SiLTmEutNiVkXC6BloWbDn//rktZxX6tnt4tKfCBPEolDqTUaISB7O6l/jCAbiogAEq3Oex61f
uIcjvLEGGu/u2ET/a2udxbfhne6sWF5ayKbNNGgIHPCAhOwjlGBLIqVfR1VmCwwL1MfaUjLRuYfw
FCbGvG/lNACP/M0VYE0+v1C1u+NJNd1xhtpOREN0v7vo3iKDKcAAPHXJd/bPcXDWAx6Tr0jsJL/R
UUzW0WDakTwBVgCvPvb5wFzcqNtwB6Y1KINrphCAdkmulbtSs4E3s6jYFiLPZhakGrRwehGvm0fe
uCXOQEGvu1h4qa178VmSntVKTu95OE2NueEdpuB6omUjr8IXtSmaYty2WADL/zLtqu8UG/S0HbBn
8uiWICmIajJve6av7GWRkrTKaVvWaz+jGu1/dwjalLni/htWnzFrkdoUkCqkCIkrUF+xyOi70374
iDUd6sF8Pg4Qxs1cpLOyZ8W39k0UDhuocRPMLj4vdcY81nuH5pWSv+83nTakaMk5WVzq/bng0kfk
cai2vbmzc+GdiN4+b9q7v14z/nE001W/FddNeuQzq6SpcnIFlDgJ6c2IkgVYVEbGlei0jZp86z8o
edGYAQ1/T/wLfKJLwDboMOc50syfWd8tpce5W1XzjiPntRO5XwA8d4xjM7AMiZyAv4NpL1XZKj3I
agKDxWAmNJUAv3baHVrUXvNFfVgAlS79dTZW/CCzPNa6Xei4xtcJeJhDPtl5fTxqeFqUMf0vOTtm
S89X+MY42/6U4Nph3CIdb+F5WCzRi7SZj6qkRLcGbCWVqOhC4Gj0CqZ4T9bsNWPsy5cQhKoDI3Tz
B/FZUOaxVZoDP1BiX32VQ2SC2kGhioetvsziQsFx0lcqDVacBdD8mIgrgXPu7qQmKcWBm3CXLpsU
jVBP/VsJb0k0adTbDS13CJP7Nskpb3BnzbQU0vWbxXCAqdSpVA8QQMORnLJe0phYNZUjS+axoozM
z/5U8dJIm9Ec3T7aB2gmYEEpTbJRqfIYeBvHPjy4xyzGc8gv2ziXUBeFI/g45losgDHtnx/s+vt3
/qMXFaqoTh0snA2VNXAzxWH7m9tpqbBo5xl4f52n4ycaX7Tf5fC69UYPv/FwdHdxxlPmKazD7klM
4uuHDe6SXEEjhUIBi0meWFKJ60gIGdy4B7pFCmPujNAS35qAGj7M0ibAJZbwBWbwIxwGICEM4Bga
ZGY3OhYJReBNacipMbU/GVO5t8XovujYZuFNtm52gL3MBxHhfFMrIPv6TKBpmKCSzP6+0Jw34VT+
x0FbFo9L0tev+fBm22/BiXQxLae7mbXMfFs9l7b/Ly35Nd/BdxqMi0g11YYHtZrOroXhnJSvvFZ8
7EWR1tbhkjonvf+6sDS0TWqgLAcJcP0rrS+B3dyjfE73pjspX18E9c/qQhU03sPqf1sX4fhDFg2e
Rgo+3s3//55wxmH3yosDC7tHBp7Goi53ac63zWhX5sPtWjHkhJKShJ0pubhKzWXZ48t8WWQVYQO/
xrM3TRGqbeNCJ5s7jyIXRI9ebY9o0IVyWvphR9hNlBUCXPrySNPLdRZygYiWpIT70Ak0GH8QYJv6
C+/rf94t/ciXVEM7HtnjpZhX2oW6qzp8vMUUW5qiRcP2gMxN5MMAi3sQLxeKDmUgngfmecztISLD
ldB1q1DUXTLuDjjnogZTh0x/0F7kN5aWWg4v6HnuG60VMbYSydd56AWnDgq+HFG+wKN+sOssG8PH
i8lc2hLve5j4ckzQv9l0H1jlZWgybRr+owUMYjLaTK8gJX2DParPXQRoFifR+QHKry9J31JgVL7E
qUbXmYJM6dIme7NPsjeKwaYjVUgp89/umo8Oa3f5CUIMHQDgXV+112Phrpl1HL2SnJhO3VWMnKI4
K2j5vS10D0iWpBI/Eakmjp02LGMpZRJ1AfHJe9tgaozyGcBwBBCsB9O9M6zC/7CdHjfpPyLue+i5
DXhY6BcVO0cE5Am1rCmzOn2kmCxvX3wES3obVG121ZHf7xpdgDAFwgxVJXZsjxuAV3HdebSmGLzG
Ek07EexsW6QamM/il/uOPVT8siMBlIR2eQaVcn8HObwchC+KkkhjlSvbF7pRWPOLR34HweB9js1Z
C+QZbTC9VyB3HABHl/QKGYeuYdiVr7yrQKM8mIoaCdj1tSDQkK5DKnhSWxuiqSAEQBCKXaOGFzrj
qK1gGE0tKur+88FEM8fqcTxlrP22TYPaPCPiT5TlE7kwt9JXz0MQFli4uhNNOKBLQDof38lW0la7
4qn+ynnJM4GgYYXsigGUh1YZdlqPykrnjS6dPF4wtzNrEGNmyj/4m88teb1293sz5ry6CjnHySUz
yVTG3bgMlExNFYEc+pZEA1f3lTnOfBFOuHpUzyw4LTnpIi3BwS41BKOVfCYuJfZCTka9of5FtEL+
jzWrZVDWTfliPX9b7Pxf+h5jzvcUpxKAmUgFq1/uN+2+DAzXm0MirfVgT7deW/d+E3ZaQFeV6HzQ
SOf79yFCeQeUgBVHSSxjjzmmT4mUckzZnqLAfzcVV5Osh5ZCDO/QcEccGZfZhNkbbE+K+5rUWdpM
+nNCIo4/e+TR+mxXxq7opU1KQx5nYUIhaFY+3ugRGKvNL6BHyQI+L7Y2dYjgj7RSTh/i4aUEI2Dk
BTF20CorHvgNZuE4888pT9VSxKDgIi2mbKA+xDJr8xfI+LHA2ik6ViGaqv5diVnwvAPO1TuAarTZ
0a9dYhAsPXrmb5eyGUk6Leoy6d6svfsZZdJeFOK9wCsAk7ku0rqUDJ1eRqYWKg+nza2PHdlu89Yw
4L32RaK4m3W+ozIzlvZsV/9BkoMwD6EC5tLD5qmwAZieLnYMyac9m+Rq2XxEDeYdlHF/j7870Xjh
Qnn2CLkngTy3yaHliIOxIYyuJ1WQ24q1d9FUzQ4GcljGQSfLKShxAV3siQe/uhjD/UGG93WFNJP0
TUiDeO2/qYdmABoTUXIIFDgQvdkvdXqbZ3H2qIg/s//urI13qkd6VFBQcfodzSNkFaRmdzVZnI6E
oc7fGDYY5geWvHBL8sfEvOe5j+QccDyXDBrZAjZnvQt+6pjr9wk7KQPAVVqCx5E3RVIxmnZkwWS3
mf7T72bE3N/H82f/niA4UFHME7cdhsSb0JAn4gy17tZvUxdnIXSgpMyJZTl4CfnvrJAla98Ob+/e
YmQ64CgnTLcbakKqH6KlujU69Yzb4NPbPxmHOC9HDKbLyS/iCbmjmcF3FWRebfYVlr21HFfGB54G
8M9kixMWFvQmTJegBpk0VzWPHzAC2CKl2SEYGx2YIUCdQfvOJzcEHAvL7j6BEByH6H2tt4Kz1/1b
wT2RAAderol/LKkfUi1n6sze0bRGgf15TsR1qNuUH+dOtuSmVB5StwGICPBhPNcUzjKgJix2B3f5
kO9D0xyUrpvrWmloWh8qOS8FKCKA20oVziUDgTGOev1+2vrM/5kQhEtZ3WJYTF3TyfY2YxDnH1Rs
fglJmyxbYvyzHkKVJUKzfDr46Gi8AmktIB9NqoZG/PcpBp2G+jEhomwEQz7dxg2Agorzup0fIQIa
ASq+HeUOdh+LXlBvoCNEKR/t4NAPuo1dI5HelGJRj2mP3eVgWUX9qDIeffa+OtMVztyMyDcd44XE
rSWhIzRcmGaQqTHUVN0u+c98GjtbpDAYUQqa7fisHJibE56rdnGzg310KU12CNhNyyJIAPKE/DOn
FLqap9RZKWLfyHpOXFwqVFrQ9b0J6B9ggJo8is59A8pU2RcvM0Bco69hI4T4uLxnrOGo9DbzwgNr
aXIHsvHl7UnFgxyDOH5HoPYTAjG+B2InBUH/3kRn3F9KbWpaRTvNu8P3rW2DcWn/mh4N1csXW2vY
PopLHYv0Q3LGa272ZxahXZJLpkOA92mE3Y9op/u8+qzC6MRa4KN+rgYO8RXdacsYt3jXBmxlGoz8
qCtVZ814sTBIZakfUnj927kqlcbqQGm1l4ghEglBEiG0z2fFMyRbaboal43TCsJP/KTXcZv56SUT
dyYIZtP+7iFaJEX5i4TJObxpRlHVc84Gi7tfNyvSGBQVR42U9WJYPZIKex6ozQgmyDJuatXhZbTy
KwN/deOLP6qs+B29RhdBOu9K7En4YaykzrLjA+g6eZIVbBqbIvf3Ksu8EO0IF+A9w7yLQPYqVA5i
yrnr9XXlp993Cy8eITBicDpZZxGFeBM4wB/GdYqsroZH617HMdhuzhmmsVlsYbwj+V/OOgFk/ePm
qIxba9pSmCmJiEudUGksHl3Yk7OT/xrkciy1SHCZh//7AM7lFfruNJ1HjNc9eMifXCHhgsun4AyC
xVA6QY1aJUKwQeZZBOjlGesrTu3spNhwE3Zjb/w6bbAkrCvLWJmiqOVNagEqV3Tpw/4KArcQKBuX
8sAtNwCjsg/1stCJ0MRe3B+3VYQ7bwJNEsCl4YogrZEgWCZojGBZLE5iVwBXFsn2LWDeofWkncQh
kyp49edeD7tjhwc8IFBbg6FenTwP0ONSDe8UgSG3+cRFDCgobz47q/uKyevJjndtE8puMA4dzBlZ
Gh8DWyI7wUOfFrBT/CywZ+K+1A4g5riPjYDcoIphaSkX1TUfDzI7J1NHBTzcwn7vD7hVjNlv9Lwb
Fhl4byrHFq4BMk6DPPatXKhqujjpHGSbXmEKH7PO/zRcCWQA3ZtGJ6541kcnbk6FZlUoSK3rns7D
Cz1qaAC/zvZB1ade1HW1W+llx18oF6FP1H7mUAkFaolMlqmwFI5+arxNkeJ3IYVCb4604VPJmTRA
tfNei+Y2OrpMYMSmHnJczG0Tcvn/4qKEBGsO1kM6bVsh5A2a2Ms0uvl+inbkSooc5aDT+L2kUphy
P8Msy2dbdzO+ZWvm8VXIa0n8IjKOx13F3ELRj6hWbwx98O9YwntXwdbDDKgY3JTX8xmw7mGlgf3z
LVhk56eoO+DJ7wpL8YMEO71gL/9r0LhnxOyi5st3IL5OoPnG08y60LFyuwzSAQvukrERbf/QydqY
GRTFA4a/PCHgMMngMzFRoTUWI+XaCjulKX8uRVl6HJFESgXYQbInIOH2gU1e3Iw1YnM4C7nU2Hj2
f1vBeyJwoxAa2K0ehWFZgBnVUCRxvbjwrHwdzkgGyKjy1/ZoFS4UKKBVFlfe78cPmdqQtvat7Jf1
j9+q3Q0mN4+azC5OXJGYPZsWxU4cr8YJdZEUEdDRHk6MuWnN1dXfZJ+CNSVlUmTUWEjtuAbDY6VB
MTGXmf8fSJKPQvqtDdHhEJp6ui7qZI5hxX/kBOhz9WhCKkojQMMQWoQowapH1AhAbrm4CKxeJDx7
4hs0ifGOdQIF5yS6AtPoB2VGb+GDrJneY9CPnusC5DxEwtUgRGayAS6w7RQSdvskI+9RK+ocFl4f
ISKmalWhi4yreiiLENyhHVADI4pWU28E5uKOdb5U/e/FqUmmirDHEapLcqT9i7BVhBKjfdNUWWJk
/Ky7VnQDS+7AE86P3A+LUZkYTQQyCsVCHU+ieR8rqkUkIitZH8y5eCZsuRU4gFKry/rwONkUGLll
n5s6Q2TdV0eJwhgN7NZsoZjEwOiIfXRkRD0080Qbh5jHwnJPlVW0GFLpcuNhiMxusXt24mrI4fbZ
cBatHgo4CYtxLxCdymwZP2OqfTyJp0efrzjVQ2aq5RU2zVHezcJepBc3WzhAjCj77KDRVaKb/WCX
sC+QNw2K8zR3j/9DcX7LvErGxIYwKDxP5EXQkGcuRv36vkvx9Ylxj6WaNDdHbKkXwsIgrCn9Svyi
e3wAJsFg61I6bsczurDRpnPsxBUlyL1qBIk8+Z+uLNA9kDdnDi5J4A5Mdm61H6xf3VDqvDKrttWs
8PfUwglDf/rxWKxaaigYbSyhdRRE0fbbKAmMt2C5AeE94Bjh4imWfWvK4TLl15puBntLa/2U9+9C
GMuemI6tE8/swcl3wQzkgCj/NoYZVbUU2QqvPnEI82CpzI1AwRhTSUIm7iUPkT7IafjXMmC592vK
wfAsnoyrrkdws43awwRaP2N/9OH52C4hY3/q+1Dg6uZlIEhtjeTBZSU7zkkgdXs5mbT/IcnrvcxD
JRhY1A3GvQGhStKiaX/hVjvnng2sFUdfla/WjdnYKSgMrsy0DwCV88RVY2UrdXmSP6iIyHOt3nIe
rqd/2Z8dewK/kfxmd7M0F94Aj/YH+hPKakiKbek5T9gKzBx5PpfL6C2i/uNS84TlPWySfoe0eW01
XNcu8sjlWfOifdjAJpVMekVWoKk6VWbT7gfBUhfJNUlEBBksmsN/63oePD+K+ch72XTahT6DZwHD
4HvW1wc4HVsTzzG7M8iEBE0RhoIUwcZwrkcGHt12oHqqu8PZOt5cRh6xOMxFV8RMPHwDCNEKktCf
ot+81eAdsryM7c8VpBu21e5K7kwnk2VH55f4vGAXzjr2fKMoIdtcgcywmYLO7WI1/5GufwbMqapm
s1ptjfC5U29Cum34CuOAqLw6i+Ed7Mx7VOxvY58uOJLlw/22xlr9rPvMFfh8PBNQDLQ/PM8muk29
JFG1NjZMd8sjZ1RwsOiq4T8pTjISd8Gs0cgZ3Det1N/95JVRG9Afm/VOg+nYZaBoVkkk5HE8eMi7
WDlqnAV49MviKXi5syWLe3FaY5D4cPuhQ52RPDubxnx7uSNRYNI5xNpxIC20Qkva79bW+cZGA4LY
IaP2DUfsvksBtYmxyfHrKzSXZ5SlvB7j3Po2N5W1U7lipUSqtMEH5KFoyPSr5FWFSc9L19Gf1xpP
Dbd5eFN4w8j0q3tcFT7MjSScDb75xwbqaI3KmgTw2wdf6Mmt70i48tGdzYLSbD3/hEd1LK9svOJ3
OYMsRv9ikowl7uCzGGt6aEyTNtfWvodPpZxRXF32X/PZtCHUm/+LSNOpiLRK6A5OSLmztJ6Gd99W
UmWuZBFBtkkgZu7l2K9Iqsg1JEg/ERy6uDasvZuj1dREqg0teCkeZQqvO4RXj93LWqwmD9LayGBj
HkPYJqq2/tAApWPOVXA1CcddVTTAZxRqh/fUWZP99SAYjOT1qjlCuUOKj0vH2dF842iMQXSNvTDQ
+1pt3u4JwBchfoIPa/A4T0mBhw+dGPnaBixaDR8EpNrKowRIv0GU5Kz+/bv/gthHZWduSV1Smtbw
kxXR2hTrpqq1TEy9LNkAsdy0WPL2OY3x4MehbGGiunCHVZnwA8xOMxAVu8bFzWOXarZK58aDgyIU
K8jaKqNbeFo/H3wYgvm/HyY5Ij4b+Bs7AimO9WvWWOUp8tAqUic82rUpQA0nQE9A2TaGPAOpSIza
gxBHbmKuaXemTpQo5HBgtUe8X8PNl9gu4xRhIYMqb0dE7MesUNFnvQqSloZJkS2eyaMuCU9de4N1
eL2lVvKsppG5+vfjOgN4K5Gexc8LLMeMPyhIAnpUPgf66SoWc3O9HsX0bU0Khb+ce0ZcIRSfhZUZ
VcOYp5OdzDHGHTgqhvdS72VMfusS54gSe2NM0AspdNvgW1e7BOaLlH3I+cT0gRIp2LaykUJaQBzW
dWUTTOpNtzGspbM4TRE8u6wQdpzr3MGj9k9n7zxf+VLgsy+oCYPd7ClvqDJeGLv09aUwkiJgZIgn
L8WUIA+IIA6hFaPT7TI1O86BtZfpMJcEp0fCDmLxtIooYKmikaSPh7WTVLwPlIH7fHfdwa5wVjj/
deQizUo+vouzlqvybDta92aZHtTCnK/Q6g0SxPMU/W7BLMxjG91WkKlvgmVgWijvCtkynnqBxDWo
EIMYuvxc3/YLeISbmpdP1fNVhTgnPCFgieXPkc9k5cN7sJvmuDnNfS65LBqsjTQQcyKSyl6jvRv6
d6ZCz3aDcdWpdifUZeEYXg4wCU8mW/rjDwthkosycRiP3RHY6m+SI4gvDlc/0Le8zQZNc1t+rvE/
RtHwQzTC+SgRlcPW+nfITlHSDH2c0xmbPcBzpI/H51ihfBaRs0sUK4rNQ3lRxNvPDs0Oq6fzMV/6
KxW4+kOYzc79VF1gnFDN7aL3ZnpRiAmEt3/QOUqJ2h/eS6/O2Mp8tLgY5B2mnvnOCdh7KL79rU2c
k71Hg62prOBaySh4aUQwwEA+SVJqd1zrTkZNxPm3dys9zZz+fZ9qqJZxGvVChbguZk0qjh6uV8F7
q00ISNYX5bNlv+RCImaMs6yJ+g41Cktet7yjY/ZaFVs23SdG3jM2GaCJo7U29sUd1uRD88uc+NTI
5lvy8R84A5hTs5wwVL4MJ6IbzsTUOgvUvdZ6imVOhSmt2Suo1DNV/7QgWPiADg2tVHgzxJvpPz05
yQhVzV8HDFbl/XvcJ9I15uh8BOPxwADWo4p+F7z0pcW0AXaZzmT7IPui8En+jorQiVZEpZbzRQmv
PlQ+6x6vOGZhQW8VSAkl6W/S/JqvNr4KO+XIBrCYBiW2nncLOudiQCK7z/4/8ENu/iVpzSYwQDJB
ljA9LNUpHttVQC+kJ2cLYY32NcaA3/TsGBTT9Q5440F1wtdrl3sc9R8Gp2a3RXaz+AykpEEhbMRH
O90KnkbzDtIDD6XWGvXKejwt2S5i4S/OyJbj/bZlJwJ1ScluVc+YS/klzN7AVX/rXojPDwIE0lJf
M300bwKHgW0g8fPQQsmW4Ki8pyf2lxu3ED75yyBv9quWAGsRYOct7UHg15KotSjUBCsvzAzBysha
ao82RBKDRvpqBXkIKYpHn0dFf1YjxvNJDEFNWsj2DY0aDMu9huM8Eb+WHxxZoe58en17OSJyCRwE
TEb/ZKKWc/kiBEbf0ynP7jRfPNyzApo3oEnxKylblWY9PFjCOhTPSwj/r/ybFkk8EfQ2QwcCBI9u
rIeN9v2giHt3GSGOcYw7wha+pH9j240yaELNkAtbq4e0pSW8yAINB6WkDTph+OG/0VlZlT/K+A0s
2Z6coWJoqAVZ9CepbGABYpacPuyvYzoP7nNRc44etu1RSM01KfyjBP2ngYFDxI7a2nlzo1VrsfYY
mT3pYiAZmb81BXYxFYfwj6JLBw5hjKOmRt+6xkQW+189md0s1SNDpy/+JWeZR+36W9WC0EbF3ml8
k6Mex71P69ZwH0K0eLUlCBFNv0XdZo5uUl/BfXsE+1lHHOlXRRMGxfMPKy1lmEFPriVtoAx9A5Sq
wVU6a8DKzYJ8VaPgDpiAlpwFsg/luxCH8gWRDzPAPSoUrZJtQJTGagNsiLC38+krMmQd3uKeTwK+
c/8hP1OrO5oexI3hjQ0i9xpnShisevl4bZQH9uvMsGiFMM7U+/MtYVDEREPoAlJ1XO4AUxI8LaAe
jo2iibodVb9MdfeWtbPosA/67QGB5yBck8ln1HMt3SXpoi77dWbtWMq1U5J85UpTj+H6VuYcV9Sn
11Sf7zBItkNx+BtjcCp86fUJGO/OgwL4je9zenmVOC0e4Dfq8nrdjc+sXjLr/+ykKJVJnht7pkcS
XQ4WIXCsr2SHrcQLmh6bmTQASrdmnkeqHGLd4dt+CcCrmKNQI9Les0zyOoHFXu7AgqU1TMW/kmbp
FXidPcIoybxcRZaP2IM09Tx9Dy8G0VHyzSz+/RBapx81HSyCfXWTGGJ5q/9uaehEBHqSvqTiz1+v
YxzAzg7rnqcm2SuMOBjA7NMTclnma09i5Nh+VNpJ8VSYmwpV585oem334xi/OlgT9pYFJWgx9bKz
3FAlYmaQ+WOsbgAEMuipOqizsID7bpIP2egSmdfvVEpVDddZeHBSW+CjSnVoLVLJDxS8y1pxP9iE
eX2de0tHowz3V/qOLbOVWbZeyv2XGdncfR0MDiyqtF4ynS+PoXzKyhXaZ9jFvDkdZ68gidvV81Zx
dP8foD8gFq5q15+qO05oThIF0uF+YuttopZn8hO948n7MPOHorRNN/7nnw/khOtdFLwfliu7yy79
clSiB7b/RR5Szp6lg2c1fpadFrsFfxxjAqqG2sGL+z5mqOkdXLGiOHpYMiIQQ4zOQ3InX5JvlMBp
yK70SV3yuIKZ1lP68UdeHeH+DuoUu9obHNWkJQ1uHf3lruImFB8YT3qco04oxRbHcpBsYL9zbABN
ce/VMiKBfIJqQyxSVyHUgjkkH215z88N7/jIziF3anXgP49/UrG8M0o4X6ckT9kWR4Ac6LD4Olaq
njw0mbOVowzwd9U6Hh2MAcGgtC+UhCMJPY/liWErnK/idg1JxKENA/7Jkwp71VPZLVJ+vkeADomP
bLuq0VuELibJgJStDVk+LIDOzg4qVJfnEpVS54Hkq74/c2flju6Iee+66KBjToKSmxRGP/P4piLn
1AokejCXhilPChsJpKyp4wf5VjA5W4ga12sAAmjUaGpyjBrI0Z9pootAIt5Qf5QWhfE87wL3hTzP
MZJylZr7Lrm6SjVslSm7661uDqO7BKbI+5y3VE5gGN6724Xgv2AH4i/LbowOLZjXjrM3aUsx1dGY
KF0mMH+aAuCxOPVWrGWIDnhntevlv1B6zb+fvBOC5QEEJa3jRIpmSeC8VzsvenDKwLQgg76XVYww
qGzNejHxN2TbMGjD4vKrQDDH8hxi8x5JwGPLGaSFT+dOYNI5Mrdo6tpx6SvZO21l/sfR6Ky0d/4G
FJHUOUgIgFkB+8jzABFVCA0aqSTsOCAcr9rFOwDMO8KZh0SYEgvDXfAeKUyIjoV8unr0U7DIPp74
wxh2IG0RIGn+33XlxfJ7vTDfAon8TKGobXwnroEtkB4AWXlIvpW5QuJ50H1HFQHOsrsoWJhtmAQX
i4WoNaRwYkkjv6Vxm2jp3nEwsQ2tOnKt+9RAg3TCJz9RiAPKz4yWGX9ZdP7UOWKJiozNnSitiiag
nNGMQAaVzDbbPJm/TJHHtDO0zUKuIEPPwae89oI1ydWewbyezOhwuP3FqfTBfetqfnLFlvIRKCRq
AuwTk60eMX6AChcAuCUE5Jr0ShtXAHMqpJn9QqG9J466rrbqctWDeAtDSQlN5JhNAqFMn35cHALb
9BPvAlhoOf/zERys7wgMQ1Mra0vrKLUNSC9GfW/KJbN0juCsIqFCwUOdAKCc0AxChTNmu8UC8CIG
9Z+0475LNrX0za+TuHuO3LeogTOgngnOa/6wUWacZIUAPG3bGwC1BLO/yZ4ex9uut/D5L+DtqjHx
fZy3rb5aX2EfXg+tk4NdX1zvXsrFEy+ljz1at0vpEoaaZZJVW5ymkmgOSz8ntM21vrUF6NuxtA6D
yIeK6+ONbROlSPAmGr9wjCuHIhUj4mbMbfGykRBk9kwswi/TeaSFZKCxBbAs9Mb87M5RQAz9MD1v
d9v/3IAfHXyJiMix6x842tUO/TtWTZ/ovWcNqFivgy0semeusFNMm8ise24twOx+8GFWmIysBMtC
WyAi5AjdVFMdr1yrcnUtTT5X+eO5qf89K/v8h8Tpo1eDbDw9cYwS+FcdqURLXPG5oiOcv2BUJ5T8
X343s03nrKIn2q2G5E05kkMH6Oascm68gnMGnILI7UeZ2JPGC6/79ghomYLKJUDX56cXSS7HKrFh
uaSsDC25jnip6M+I/N8bxdGgEk1CUNIEJmwrz5oEUeRFK9XzOfUNoJOh7voYS9m96YL03asjhIBF
DGyzZa7hzKeWlde6CojQHzxOd2YHL1F2BZ0iPOUZ8EJCc2LaSKWrul33YCZEgG5TPJDIKvpp4yWf
mlWj7rKbWTGEMU2l0vQHXoGb87CsM5yFJC//v8LFwGXCLADnOe0DRoVMmoVREPLo2EgdpocTD1fU
yxtL3H3xtfAakI/aDTXomYige797NjC9UYlOTTO439GqYl0Jeqg2tK5VWUXL/MolaJil/zFfsZxk
eLD3twenufaDVSO+0K2aheXpo2WL9hGIbAejvWBOlji8Qq6QL4moNIiW5x9ou1DVws2aK21RZoXO
DUw/IiWFke3ahQuy0Unsz/zJKjNYy6X29paaFKdHxtWBsu2DdXJoX08vVh9AWmbK5jwSQscxxHvh
hr89RqH8O79Ym0lHq0hzOis4lFV9pHeMEu7Tq8jiE+NBAIGQZawEplONXfd7Y0OuAPI3NnCK6QCM
IMOI3+OkmGwHq+jVrX6MzfOoPLyMomsj1gU4Qw4hh4XsqQoX2VYtQvLJEAvP34WliUaCRcypvjPc
tr+h0cktYLzRpD7sM81CGNytjV741Vqk6ZwIHLlBa6q3hL/yGw6vIRgJyvwbv0YhDrUHCQqlSmE+
bBb+GcWH3dAHcc3ZrDn9rg7KXK/0PvvxVHwvxDkBxpzFFbI4iI/abd0Q9qulIf2RIoKsz2rpbhGQ
558k0xln+zxgox0yxDHJfMeT3TZ9GOe4rfE/+2oK3k1+QIs9qDHtNCsoQ+exqMJW9MJdwNEPhFyq
u8UNNsd7vzmGSfkjZol+Yd8uqh2soOrsvFwNehgiTq0aQo+Yxtc3LucOSe70JV1CBwr/qBQMlcTb
zoEXo+2S0+vwHuuMo50iCzuArx6wxsSJWfYpMo8+yuP+WxfFUwG/JKETHuikjmL+xorcub5LbN5N
XTkFvlGcPpvjneYXwerwjuzyuGfn6jvu9Fi1vszZgThzgP/C9r5N8UwIR0fHjqWstbv8yNmNyobe
5PO7rQUxF7H+pcG4LYOKGdYoixiVdoeHnX2dDWr1vuLgVLV18lv56FTzrvgP/RX6by59H1ZEeP7o
3qg5kOoUsnx+k6CQabY/MtY7ZMJuSou17Ym1Cf+Xzq50vW8OvJ/4cMw+57gvWVGat3YLlR3pLxQT
0ApP9jTmae17M8//dtrdACgIOel6oeA6EqQBwNFRRaYJkqMwkpRVi1hMx/lTFBJv6cDV1xZL81XC
fmrlqqN2cq8QDabs4H7Y/p+rIiVmdcr6UlfpuNeE3ga/9Bd0i6ous/bawYKtR0CSZ487H6m36C6p
8xPVEZ5n/nGI7HG0cXGhZITSdswSG22AuTr01IHZb05pWL4guvoKguKz9iPAool+iTJ4QpJHOy9F
DkH6cR+RZz7N6asTC9IjIe2c/qVPR3KqcNT0W5ADP3b1VlM7Xvn/JAfl7p1QIX4xUHlYdXFSOHMI
7ojNiaeCd0xw2yl4LmgyjlZZwjGrHCmJ+ehiGUAgMx0PLsO3R33iO/Srjrjm28jQLQzTTuso4B6D
9lrmnZR7KVIh1XUJ/Fe/X01RP2BKf2NuvJjDypH/lAaRXUZFQp3sGrdHX2XqNX01+11urm5voc3C
3Llo302lIKKzOoPZKrupGi0Egmfb+fpU+ZplfyMK3vUbnvvtibX8NNvDcaed5qsrG7soc4ZGzuPS
M+bLi3mIMpanwuQqtUEQMJtX8T+6UVE1amjbV/otLZLiF59fzXw6zCTheqG8fRyhcdgQOxN8DwLU
+Town6DNahGT3Ej8vAA5JebMJj6/4J/MLFpeMiI+qofz/+vWSvAi23XPHY47YV3O2b0wNxC3zFNB
NWf/iZ+uZFj+05Tv4zAx80f2T9cDZpc5o7hwTEIGv/GDe80AKaM7NVQBbRPwkH8jGwzBdQWtdLOM
XGwgWdh1FobIr3F4OCX/6wT6DxNQAixz84M3BZLz+KE5DOP+FeUKEorLVW4mZGcxPUw9hr8hoD5b
AK+B+ZHNBBBYqolaxfSQNi3rZo4yRJNXLPnmvi80JKnY5lq7RNQXYHkicSawKwLpYWVAytkXeE5H
pFdgdv2gSQsYVyC1C9wiT4E/Y/yIg/u5ah7E41gdydjb/BDRpdtevOmOmrgM1J6pCkGVc49lr3zP
371/F9HvfHyWpa0cJ29ZNYM6PswIy+NL3sf4DKo1gyMTFiWfLfT7rrbl2JW9NU0uEonxPKmbgZ1e
hBYXJSt5JRi0t6jEdtjD0R3wIfLcn3K7lvD/g+rMaYgk3hZ1+aZlk7cY1SmdZTCXlCIIHbreW6bp
9KMlU9VXIyAVK2O10E4gYRl+7MkX8+XnXfx33OqZOLyE0zCpr1qqkUPr2/HxpYTnidNUbkioHQit
czXIO8rK57FQQEVxeiV+ilS0CDHNhhm9t0w0S1lTt707TXjh+RIaNIWompPIqZLFWzNB4evrbz/X
Pl07w58BEts2PiLLiFMgzjjSPrXkXFdYZowO6RLVs3RCDkmyzNPPDtcoywIqbR/oMrsYjHAP7l39
EedMXdqVP7ZPyFcdmVvOBxTJ2hKndK0aDeRcSpQJ1Ey3sDbNWE2ZtRqnH8/xsBWOrQ7CnXRkX8Fa
qLiQvaPZixMKINH/geMdSUXgOVJlo+GvCk1GpHVeO59v5UTZUP8huLptmrF2beUkW9HFmP01Awiu
+224h9S9IY1HCQthpIsnDNiUtkyZKitC3qadn+xbtMXeHTQ1+utuucJ0CEbC+imwzzzpJVBmcXeh
ONpahdGW1EqMI/uVp47agM+wAXcDUIrX04f7WXjnYFqfra6DU5OsC8C+tkKw//lI096sWuvWej0Z
t4VlW4+tfnwO7n0kLMpR/yqRQAsJJvSnLF4Hx/gyD4pEAbYmdxhVKfaMO8UOjeoZVkrU6d5UB54F
7RwA1IczAa5RcN4EcZ1FsIVuXIjvyKRfUGTAfnIDH/qX4DEcjI9C/Jn67r/GFPu10j77207NWHVE
LhRn8KSp0sCFvrgvc61XJuKCAqpLEtcO373sAWB6VlEzEAJY+gu/aVKJ5tBAyUG5Vy+g9Aci/Ba2
SScSCDEZ+2LkH57rm6aoD8jzUSt8yTcuXcYYQnSUIbIJu44KCLpYbpn3rNuyreJm+1AzzJrYV60B
Yb9hYC623wd0nGx/owlr1WFvQiq9J9+5z9G/4JdLt/Np2C0HblXBr/eAxFXmuHvGh+2tpnOw5cZz
2+fg6L8/e110fJPWp9WU5HqHNaH81N1xOB/DVWhKgH4CU42NQJ4hcYi5DB7+2VTMFNRwILRLbEt+
bPuLpyPacM0sVa8vS2v45PoDrCOxOdSybNo3eXzyKaZ23MSuqNjXtql2Yth4k918qm5RUfaRYWB6
AxDDfHVGCiLwRthKY8PeWg8Rf9Q1RumJXDPvrGKr47VL6sx9JT3bUQMTdNj7h4AvYAokMq87wPlM
RQC4t9A1BgqLB7P+d1uTcQJ+UpM5t403tnrnScfnr6lvlGnjhkRRLbFWWfYktzjqv95EMdaH59Fx
KDYcZP05n0MJU6uYExFU5V9DCqFP/YZDcLRP8WeeqHvt9C/iVMwGvy/ynPKa/u6Dd62KW8FVsWbz
OT8WCkTT48s/mHcw+LsrnInLAUi7Hdl01fyNmivByBXuTmCdi1+nE4cGVkYVVU1uY6pSfzLtl062
tYfCtazFoisk8M44Dr6fZ/DpN/3JvZhkDMoQHzbOFyDIeryVE/9/YZDcezSXFnl9CYVaFBjNCMWS
oOL5ixxYJtJC8BZxaR8Poa9BqJDNAnRf3D5uNbXlhOWAJEVU6ZnOChqAH1iQ0upKzKS0oceClp2N
k3dYsn7T9/FonkZvdll1Y7HOQnmOQcpxcXSBaDKk4o+ksCg22q/6k50OCq0VpBumqoQ38DZxwte3
oGysdsbu84MLPbtsp18f3tpeUUiFW7qxoWc4G1GcpeQdEWmP2H8dYwJ0iRayL7G/5Y7m0GBXJ7x1
cuZEbualRQPNyReIZkPXcg8terR3GZOQGkqs2rWMfxiPW/b2JDc433UIANB++MiBJ8tRwkmi6cIL
URozTSDOg0YVKvnDNYZ/wKdU9PK8kqTJ17JqvcL/0a2eGQJldkc8QSOLMCBpv7r7JZmXMFKvi5tB
F5u7ciDPLHCOPdlQxpwn+fsa76/jtpK6vSmupnJwJWXfF2x4YwoDSitIkREbL6Is/u00cx4tooYr
Gs1THwePeksGzC0M058UAq1WxigmIB1D0oApG/ZNgQYiumWaZ/eyYG5OxWhS0jSzOcsEOCtMDxmd
GAepPWUQJbXk8oG2kx9RRne8BBRRr3vcHK+lwIfbS6qOilS5r/f1bQeQwUZsao+j/Yp90KoNxGwI
brSZ4ojr61oenIpEZqg3w3iaTSKUAxoupnKDzbGFIcn4EtnlK8BfAP9xEXo3kvpSoWTM8J3pvvXV
6yaZ69veAwK7y2Tv/t+LyRKzoIizL8qj6jtqdg1ARhLgaP9RLyUjxryVfiGjwjmGbm4RBC32LCIL
jlQ8Ody8xrGKZ3tHGZudsvWBgN28/H8dUyy2FUHA/edpdPOaBdiZ77IJXqjdSybO8ITVN42dzR1G
C99Xr/2xK+QHI4UZ4cTPNffopiPCasruQYz4CFi9cKX8vKTOiHBFHJQ2x6iFS0wl0oP+tBUXLGb3
IeSWJ9NPtBVdMtj58aPtecIuEPRjcCfDSrDIs9XdmIYsBNrhxed3ZQzMa2aChIBmn0EZVWgEY/cH
l2sZZyi5/S+6fCN05nbBJGp+TpUqVx8f9GParm7Chvu2glsBqAOhj2jaSrYHcC8aIe9SBucCnQ4P
FSlipjwm/cCFPCX+xjvZCgAYM6d67lBgRQB/a7F5Hwx93SCcwvdXaoaR6HVEpWBxNeLlvVHHfO0l
SFF5QYbw5l7PVTWIjfs72sUFjgJlsPB6lxND9SDKzgbH1UKGnITYTitoI+NmxDfr5YFGKBI6XbjQ
D/WHloqL9qM7rrpU0pV4A+4QLcaVbiSu1uQ3IwK6k+MdCOVFcU2r8qXkTOtrqEekUobqvDh/NAK0
/ZvVfLLarmcj043wz9YsjRbbdgAQ/o+dwLboHV1veUFDDKXJGE9ToVVtoJaiLP+xB1bTNJrc5ldV
C5uI3XewBGMC6qk2FfEcoiERV1GxSaXoahNfAn+hLMVgg9lCrVAAvdadfvvOwS/QpNTjmBd8t0DD
0m4SZbbOcPn720ceTCBBMG7plRSCsWRMI3+rlzkVAOEX+H5OZ21kAI56zq9f1UD7g+FSTAA7aJEw
2jJ4KKYSZ80WQ9LntFoGF0FsHOd/LWL4qPQFOIgXNkq0vtG5+9GRtUh9RVJhmAzn5S6RCZk4+Ahs
EbHme99m1PogiHyj1kfUPDOEuBiO5kV/YXFOhwx6+pKqFoTkew4/R1j9wBv+A77ZT7lgoVfvLa/y
NdUHbWkWBUOoNqt9iFkxCgTv7EPTVizrYNbZ98kWI8ox6SlKC0hp58Kqwi4e312DqZg+1bXoD7Rh
CLB/gX/cil37h95IuvvhCweEqUByN/trvKhe+oCh0sPo9IbGhZ15pn2IAFmLS0B07Fmt+lKpXA6K
AfWR+DSOBtmuvV+cW/hzfQmegnRRlGEBifXFnwyMTRXsggycWh8ATp1bttxwmjBqYKGGnALB5DYS
/j1I7z3OibW0TwH8wcapjwo35JkdtNaxccRqvkUI4Ko8wtvyH30pmpZNnZjR4mz3VVKvt7KczNVv
nI3SnO1n9lQLfdPGd5dCbeing5Uj4VPVMXFiyBCH/eazXvntZc5G/E0GhXF/yKvrK4Ve2jdZataU
LCYE2zA7nvFiM0Sz3rLz9GgpCocMZP/GenG0Pc3GL1o/6qCl8KdgRRreUN/Ql4GIGDfKDaHFX63j
N7xjDYP7oM91FgID7vHWO++QZZzL3NfrADBZaPjrBH6C+zwctI8K6qZGlVd4rFhQjNgR87OsKik9
ZaUMm95ZnAIo1UM4JAA05SmPYcCQzQI1Gy94QitDAgVIyyDJ7+tO15AHtCWglHbe40k6daf9izxp
2gFOj1ut7+W3EyFhFy42qYgbWwS2Hn1LBDNUEL0StmP07fkGjxXDjLeKYp79dPMKswvBiSLhRKam
22VUoos8cQCJwR0mbzeeGI1QFLVKeII/AwkxxIFW+COf0QYxmBtklJCp3YV9YpvqPeg9+0xgG90k
OTiDzQfnISzXS9w5f9VhifiPeZHi8q+w7ocT/GXXLXtCCN/dbf61OeVCLcb0l8l9dgY1595X8+66
raSFsGeTDdCdw3rOk0XpkIPwB/mq4EiI9KifEQaL2q//OQd8J2PerzNPUyLeZAzvK9THtZjbxKX0
FmjDovkV9Um0yox5xDMHvDxkjacl5qP3AujVXAN0fbyEyOZfZDeV0lkjebrpM+MjXCJSUTxSDINH
0wqF7Ij7DdkFYsGUWSLCijNb99zcJxZWlFA0pexGSk27poc+EpV9XW0CD9N2S1LDEMfr3/VBmvZT
/SE9J1PWcGCB1CqLSFUaxD6kuqOJNxDZRhCYGCANTlJBPRnY1IJLYNRgLoMlu9cAv5EgFfog2iYE
Y0q+cCv3LzQ5uRhSaurBFhNWYS/bAJyUA4sLO+c8D86qsxFkCAq8nsKNKnfCKb0e2iIMOB5/BK7/
Li4uuiRZnfagyhS1hEcKaSHyUp+imOFK+3sZlC/QhIGMgnjsDGkSbIpCWM3Ek/R4k4bsQtW28XAD
UknkoAjS1MKvRFVN6zg//eIh2QIVczO3844DLu8O3LYf9Jxpp7tRbOTedNesMPJykJriD7OPNf8k
R/zlQSdVkr+9biHl6tgSA0vTc05EmgFM8N/rOSrB8lnfYj+OH1QWS6W0oi1PcB8gOIZlSdI0aIhP
hOJX3jszbfR/KxrnL44IcgUnSDWf3L3aVQKf422/PKqZliXCeLA51n/bJ4yCfygSh10YFRiyZZiX
Yjdaa6lJZsk4+sppXYkiVR/6FLodWl7bNazldtGxT3AK9KfhhQs7vEZCXPsFWsi6TEVAkExEgrmh
qCC6vx94gBz5C02ByAAkYZsIa70Z/84GjA2Z4FYitWMMHV1hyEZguaEcM/i1gKGivg/bGZHGKYTZ
xUIyBUGJxkfaHjyfBjDojeh3lv6XBvUUEJWCY4adfwXJCFb1MZlYni5ANmimxHUFiKtD6NNGHFsv
hxSBkjnGr18FXgFwcJPyZMgHdvFqciEVB2ek/lbFmOcrOC2uZ6CnF1ujVjFiDfPVgSdS5B4S9z6g
VHRimdYnOvLxS83+O8+yRX5993bkC53C6tn98a73cF/EO4e4t9x6n8GZ08gYy5vfmXFRJuCAWNUS
15qRElD9sijCvqrQ8SXibxKyp5sTtjf7t1aXVklyjpImLLWmDDuJPRlmyrpX9EiJB+Dt7AqaLr+V
8OZps5bzH6dTgfg1rbkq8TZi669/mXkvaDr05dwfz0Cx/rlqHSIOKlhvi8qAfKr1QzX44kD/2VbO
X/q1oRODJXK22FHzBhJ8yBEC18UVA+2od60skp/g5F6WN7JLxjnU1vF7ND78AE8H/Vx+gtdiun2D
5/SpHhWSKIQhp93B6wdcEQ28GukqPXGEku9GYX0GfQ19fklNrES4rpenKliId89ieQ/phDrrHYgR
l7AiWgtd3tDjWXzdGG2HV6Ywu8RojDTeYtvAemHarVO9EkwEXzZQnAxStFJDVtqpMR4jHHrYtg1b
yOu5MPh0qyKscsQD2BSSpdb5eCUH0EfBCXEG3gO1whk/HP+oltTcVWflos/6HDPPlhx5dj1dq/S8
64c8z4cbQGtcYrb+onhqHdTVfs3CVk7mnQyBI7yv4WadHHjW8jFAW6vuCK1ohJA6x4WFu6RaZPys
Y+/3AGwpklQJgi1JkLOXORgiGbAIdXZCY+MHCA0U18llV8xtPkCHf940f8XdqP438Nkwa4PX5Hif
d3KyXBtH1NggwOVDmcRZaBmL+jDCUtMnENt87cbhRVw5RL6g122MKKVBamdNPtHMWJqFk9Y7Etys
fM7rEivIAAnbBqEtO5+8eNPIAL8u5Cg4OVjvqIZBZbYfXoy+pKtcsRpBJdqyR5c6uq0sdiecfa2U
Akm0PPblCuSLAO28DQspE8AGs1/jL3cjXr87RJ8HjFDlZlYJ5w1tlHHNjut+/jEKwoXWQ7Uc4BOL
zLSLa4OpKVyzkuxhNfzx3SGveDO2rxnG9xdnF+pwU+HllP0W2SDJ24OheL9AHOFMxe2PDQ2oa4E+
5uWsARZ3PFNbXbHxg9eK+VVR+223AF81q9UxILwZI1Dx7z4MohNXRdgk3ZHdAv43QdU9aMV48AkY
qkHJF2Cm4E5FkIYOSTCw4Soqq+zA9NhJ/iWMdufU7NaoMnt9koa9QF4NerDA0xe9dtslNRKdtzG0
yMKFov82foQcVtKCZOR6qF6rzG7VT2LcnR+4A9B+nVD2zjzrzhg7DhJPSYe8DSdlRKDjm8Kc6dqT
nGQHJGMukD9FxBAqX03MW86S71q+8/CyhrHpzRdeFDonmoUSX0V6ILpDRNZOLcVGH30zD4eZ2oto
T51IPJMVJ5CDe1ZJGnw1+GXd+yapkp/mUQnR2ya06h+I4HxsMJOVFopCNw8Ca9CuLIF7gO69tG7l
MdaqLfs15Nk9uSH5Ofovaxr0tRFan9LLRoOOnH4da4DSi2sAQUMp/BTtrfs+fVELIKROXXvlg5cE
rJzwBnBY0VSjI0qoKayLoDIOTMNXKghTl9eJNEv480gyPooI6ooo/sKa0JjfJrePBvDw+h7vlmYR
Zo/ErHnvRtuZ8S9u2rGtXityjeDaKMi0GtiS1llLmO9xBpCYrcfCuXsCDvQK/kYKoBfRsLG5ZXeB
8zC8ws5A+wqZHfFzGyrDmp2w/gUsPze/JN67HiqZhLDMqrHmMIe+ATvGns6IeurntBvNgKB30Uzw
0ATFEBUBsleZaT8DeMIbaNS9niTyfOnJvcOlM9Aw4V3ZPqsPameXuTBtVVCDbVpeZeO/1oYzEy6X
dZ2BpK+Y2V99xmGH4ip+3njx4QP3BCoBFdJtUXYiD/xGN3iQCIQxLShQJcA7kyDkrZVHEiBbaHkm
piJowwH9PbaH25iwOafaNaNwZGhrFwkn9FdnvJp3Fn+QHmt37kazxAassw0A4OD8HlxezcmwHyIN
ho2FtvaMHm+l8WVBJiu4L9wLQ3iUJdFLLJbXaBEGzllEeF6FHKy8wJfVhwuNcucxAyQncB4kpMDg
oiszOb4vGb/XFnSrrzHwhhlpolgVgiNgwgaATEsOsEWbrhCUiOf3Y0Mz82vavFgJMskExmbqDARU
ChwCdMIC8WdaZp6M6nLxMA6arH9jaHUkW+blHaXX+NY+bwli/GlDBPWn3Lnvqfwrysc4N2nLuvg5
/5eEl2vVu++kSvHRPSLG4M1fQsLB0IE2mMspcckECJXH0sAp6WRJXuOFXTw2ijqeLluDG7qyhxVp
bOaG7jZhBm2wEIvGvMm/L4ABRM8Gs+GMsOXk1I+VVgYhXcyOiidco9BvXTF8XWnfTCjqn9/Gp0Uu
peGLSGx25ZCwkvN1tpoXsx98QLAbG5MzA9LwmQ1FnPuwn+pgyXGddWKXNh3CBEV4ogFwrDikb4Fd
O6QJoViaz2aTI+CdIcO5hPHTnS+5jp++CoJ2h3Y/grc/hLeNjAEN+lKerR/S+FOoEvjDjpceybDu
dTp2ttHp9t3X3CQ08tybHyUSRpIUWbmefkVOryT1lgP8MBO3NfoQPsuYWIZ8JPWIqiLa07f8JQq4
qr8o6VskFVx8EXCVosM0DdpxgJrQpo7RIZjFpgVrBqlhbk+tiYc/NjiXPdNRzNl2fbajbYu0M5oC
DG2wGkIdcYqcFu26bGYAN8Uf0MLyAVAQ7Nhdj4QT9PiUj0sSjbdTCcH73NcGxxMXXPVQjzz/KbGE
RE1zb3gmYbNpDAaFtauKFNC05IofK7KR7Xz24m9ENroNiTozXOHO4dNjzQhfcsVlVFGRM5ab2CGw
e7g6THMCM7YbezA49BG86jD1RE+zmWtt1dzNLhfEEgtDHmskPC0X+pGWEX037v2VjVMJX/kWxCUq
CKTMDsSNgQJlghq+Lv7vgodWgrLcTR2UmG69GG6thw8txUIpbAg/RHPmP0lDBp8Ko6zgwMLco8Ss
1bjKBCp6NrQXxbQ5PFKlvVvIqdQTU4xzxsP04rNPTvkFnLqhNBmvEsxnUUV4mclNKn6s6qWBwnFM
SNoevDug/fNR1ovbSaCNTmk8OBdTkju4Y/kxInqWEIoPMwQElkKWwTEzXwFQKJSTzX0jS5gQyFtI
VRgbvQKiH/HwYB8plw5HQ4Oes6jkhd0vEJ59QVE65XJownb4brMKuTDacHImkHPNDeSUSAdua10M
P3/o9ejgGjBJpMmrsKxJf4LfErdG2OfWgjEKk+7bwF+5kR9oDGdbzNUuZLvShEUOPLtogCoY3b3n
FdqxjxPOJkTKY+0YxGpJskEFPW0Jbx6k+vHUS17SHZwIvQxOTG3zfsEkeGuCGWHjfID0nye3BG7z
6kZFtD6KlwAqKtkeH5uMX6kD21GGI0+5VD2cEeihzuXuuLN4wuj9WHvJy97Bpe5Mtup5hTSoPZPO
7zGWhW+Cq1OaSR7DbXVPDnCe9GEiiELi/C28jSRJpv607jGBiOLVg+IqR+Mc9qAg3iRPl74uXs2k
BFHtD0WcaR+QXFNjz6INpDAJr+S1MkhTifT/+Y5XZjJvIP77ZttCV+WG4Ku72k3n8ixj3yRZCaw2
CU7WaMJBZ8B9Bqud+jxGqfMmdBhdN6aKR+E6U/Lzc2q1+DwAIENRQtCAEB4L4aKW48apjjG0jez5
GDDEO+JsIQcGcflwYrC3atf2HnFpYKTE9jxx/p9KQWU1MCIWWuK1ueT9IAHzQlw96sAaNNVGcjfl
WAh7i/2fAE9QRDjWZJ36xbTI/2KTep5pZ9/j3Hsglv15PxqVLe5xKFOPm7nZ/CctXm1hjT9fwDJk
TfUxOqVDb9F+AEkMBHN00HRy50jGHa6rFXS36ySoA8owaJ5S1RONKDxBFVCA2AQpFm6cVzcTBju1
byDFYH0FdZkq3YxChKy84I4VBQHBlMjJ6+xIzrlDJvVTO3pSmodpKYGy7zIaxj2GEJ8i94ekjOMN
xfA06aJ69gy/PbWji11yWgx+pCs1d1ckD8dP8ktwfvc7jypa1y7TUQe3lGXGdGyoBJ9lvduZoG6V
HwYxUisy1dC2ceABXgSLk0gG0hZIfCRFTT3Nbe52Ts3V1JUDLmQYUHjKdBLbD5s+0Fx7NykFQS8d
uOmEdKd8Oi8Mh9/opy75DstBzRKKjlxvF+GZQ4t/KYmdUbr4BSMWs7ZgmxC1L3zq5kFT/YF4Vaen
r1pERJZUntw3kUMPeKGL2uINYrqj692Z4f+H+o+/PwY7wFZuDPKZGx1DENmxE7LjNNKwJF3uBIrS
bzSmcrHAnTI1vGMW6RkXwTncufW982yr4gO0p20aWoK3+TL9Yq1DdS7LAijRLs1uQm2vBLqJhfa6
YYh5VmMzXUQe5MRV2GSZH3WmLZYvGuNPbKJhA99IPNsv7e528EtsOxXuwqA5mUXCfk8djHwZaPp0
v0Ss1pnLIiVQSnYYBph8XYHCIZqE+O5wr4tpYn2c39sz8DRkj6uDq0F7ej9rkqO+7+IU0B6kz3RR
crNoJZLowXlm5pEKoewt02NnC7IIut7dWyHICYSg+6u4yrwzwz5w7cNwaDqSVcCKrlFfZXg+scg6
4Dq+OVFRexvBzEhfkjvYSWjUFb5PkLMnI0wOkJrTL6Zh9ETnWJLxy2m55ZTx0ZsluITet+AjwHbp
uNdUsyzlWNxzGJMKG89P6WWWRh6XdjZi/8tRSnrAaXByVhnJSk/+vLuugmKYtakUmmAeKpg7FSVY
Rh7pjVSHTpZVx7BIFlxM9lJ2n62mhrTI6rrEOLLKBCTSSbqUhqCvBKVRNws02WfNjVfZNl2oIu0e
WisblF07D0TgkgBcSyNvXQTc/c/z/a1Lgvar5cQeZUZZh0W8KnqyhFJoo61ewo4FDieComxdidk4
R80GAfm54JF5BzE5zS/B7IoKUDhGBYM9m68HziDgtZH5T9SgJ0xth1BjGDXB8nDJhyM9Ik12dtyd
5BMz9/06LDeV0RRRmADm+x76V2Q9n5NRHB3DfudOU7dmCWdBLG56rVdG+H/jv+MmDmQDNxJ3xZo9
k3C3TiIh6PpIBP1Mh4YwGpUl85J9bQCC7/yOGA9ixIYlBKVZsXmVD399CvCPbOjeO/m0zRcEjoeN
AAwlziTu7588vuTwnSxC8flG2CHaTJClYwdpgMk/5S8dKJWMfA6pd+eB2lnnUG9tLE9pUooVn88d
ea9EXyYqKnc1QPC3FNvF7h3eV6DR7P8+R3rb5MrdzA9Cef/u/FFSw34lzCddYxH5rVgy/661vJ97
tfAnDKaoOZANOyKjj5KRG8TMnztirB/hLBGPHZXtTnXH1ePmBELWLkgK31tWzbjWXi/eH5qf6gEj
ntHXlX1npg59Om6/zmifexMRhwGDL2vL+y4Im+1o6k/5k3Wx/urfuRwWBo9yNjWv6wENapgX1Uk5
KWoBqoe8C3T8UxmFSXi6+ME/Gf+vMgqdZgJYW4RrdWNP9qqAvdESwMZrMeoBxCt16stBiol23huv
xbVwMrcD9RLewuuNIta3UQgV/ilmivvS+5cC5Nlyzi9ZWl+ehWqDpFaIX4MnRsRo5k3MOEplzvvl
cjBj+WpmfcjHhh+4RrUrddKcaukV+ebNa9ttP1M9jv7b2+EcBD3k68XqHujnAoyMrKKwUOgSLfoM
BIcFpro8O85QTVAxxLHV4uCylyVI7C2QPqcOnIantGFuUzJcMzykdwTVy4auIHfBlRYi79Ah6I1G
lvE/vrYJqOI99VEDcrB2hn4s9qvXFXw0HMbgjVnDRZISJwYmQ7msIRdNbHtgckcVXcTXjM/NKM/Z
8QVJgcsCVpXVneT7tr2dU4X0mE2d4ngL3SuWnRJnj8DVGCnxQcgpFbWfGLiA7Ddp9iwrIFANS2Q5
rMYmtWf5vsYqtcOPiu1uhNJT0xdCYHnXuzC7PB4VCPGvxtJPyCxlsW8xApjHthgz4sr+W86supap
4GZNZiS5U1aqRyjqZi0v+mvevaphPyZD/WmAfdlPStPFOjTSuoxFWY7K87bdPbt9w/Sn0VohbyQV
dwfU3/TCofPHjbQcctaaHsTk5yeYwHX6sqs9k/zuRnEHd7RyBFpACCGiB9kUXpAtKhmVln/fmwEP
mOXn7kSrhVpnGRifLQah9Pk2+4tonLhDj9eQz15yeJKJaOxI0zzKHITR53LjBkj25bBFfZVa3Ul/
mUrqyvRyyZvKOFyEdGhxFUqK/V6Kf8JERgPRNX/DAzaY/t3dp51R+VXTIL9m3mtTXFacgXv8Bs6F
tqHkADOz9xYOhnCeBPVWuN5G7gQwLm2WBWKTNYMSjAB/cx+ytvNgyABd9VtSEsm1mfQ1sPJhroxr
zIM2y4prrDV8PSlM+9sBjtFLCD/J9Kfp5KJXec+6aJgcZEuKwFL+5nt/CBPDtrg6ODVXqqGBeGxk
mv+zkm7qFbhB5+MNZZ3Hl1euQT8Cu0cUm8ViHnPO9Dfn3adfWLJL1ZrWjX5QMByq2yjC+BVwbZTr
bYlbo3TobI5UiNMZiZmOaWgyqqmkGXNltJmyqYWDBqjLtPexmFFXQOOpz+euVHXh2tRCs/xdrj/w
hJVAN6fDV+yM8YzO74qowEzO0R5kLVx4QiYs3Dq16cuGTBmqiOWElnrNQWtiCFvHwcM/y3joZzwa
x990mxiddLi9nwphbXzE9pD+9MvJkpHVPpdkdQ1jN8uOJPrSUtee+9fyKtWSBzQj/rQOk0J27HHU
kwvJohMtLGSiZadCPICWGrqLRkXWMwwOGQuRBsh+gfpSCeFfeVW3Mqm7zGy1Eg9NfuuNQjJ6DsTv
upsqq76icQ/P9f4hdHGHm8uEN5vE9eagOCnKEMa0sqDlymgglLrh2jDRtFBPogi83z16lwFpjHGb
eFmmfxvKCBZXxwhzMxW3QvW+6+KXf4ic95nJ1rSNR7R88YlZWmyg6AzpdCu/p9f9GUO+FhhcNb+J
zxbbWFsTudBa0BxKibd+vYvBYJUbnmQCHOhXyvjSQ/5s5RfLHl3Vbu+E5fpUywkNc2oGhwEjAMZG
Ts8U7e34R36uJRN0JKJgCw62KbHWT1pHNCB3dk0T/DD4dSv8XIgu2WvuC+SWAgo86mFob/Kf8JQm
9txJPf9uuqsQdwOT0aTYYJNEe+VJa5V/sHubm2Wycbcf9a3IYQHGZV/DWFgr/aLt/X+/tr6sbt82
0mWuNGOR/CSMNdqNDv2xoEh3NlunGezQ6uY4MafSaTO76lPwj8Ge8blrm7xHB6JYhriOp2Zya7br
LvAuzDiCeEh3WlE+KCAAoQj8x5Ue/k5SECi9VeycdS79swP/PwKDfABUsYR2FFuDM5j1AdXapxS9
31SBaWUqQDtdi00vbz6g+OvJ94oMCWPHxVZEp3NhaB8hKiACUiMSzjF87XDOKbc4AZzi5JSycScq
kx9g1YFVKR85DHXWHIYF234Zl4mLlH/Z9dHghBW51gfmazLzHo0w9caDILOFsXboWaBYunV2xmD1
AI9WcGfg9uMBbn9mXYfEEgf5SuDdvYfaeITyD1aoRYvqjSF6keuw0M7SS/2+P8yi3wx5NsvxOdEz
b73lSD2sDFtWC4JjcvDbakj3h+EpYo/oHjuVMqP5Nl00UcTZjbRdF+bRRtVL2VLK3g4xyUKIXShy
TrWDRZkdg3Bn2ObzGodYKDhG4fW2fZ0O2FcQj2PnkXtA9W+1c/mUr7L3oBCU42WvZGeMFGC8/+xy
jIKnb0wghe781NYRJXj9CAX2eWo2m24GSdZ1qo3A9RvWYfd16oRux5XrrDtBhsxyC4+F9SMv+65A
CjN70ryi8xBvW5uQSWcSXOaSChDuG9X7ia5lV/9gfPnYC43x/OZbkrNRQ49A+2JTsjMU/uRdWUnp
ojai0cn3yj6BJSUNK6geKz1erqX/CIBerel5pqa5CIWZd33DjcrOaj+sH2QUt7vAieShfqWHkzE2
kMPnCXIPpesR5TmnficcyHYIxRgH4N0DoWhdZav8IU7FfaEjcabW2kxsykbmvI+HM54H2lvsYtzM
lyXG6277FdknkZHSRFyvSNdBIyz/j5SW4Mozcw5lFFGRT+f8oTvEALjGxUE4088byMrQypmMEwXo
NeKntd+AaR8f4caagWxKRBqrWESYaBXbNM4Gb+JHLldVYkcOvyxsg2UNn7nAovqI07kP0o8l9anK
tlBUXkue1X2xrW7uEpXnWS6159xiXquNuoLi2tcmqudyweGFFiXOE3g1SHphEBX+nX4YirCYKhBs
lO/l1oZwypTphV1yLoPx7o9bh1Y4S+3LHxHx+mXW1u70SJ0yx6XbKsTD74nAqUUCQoeK3R5FLUiX
QMxbhOK2RXyOONtasPH7MCq8uEqSKLyOf3gskEm3+eE35bAnDyaTrIjenVOskGeB6diEIyZmvVsq
pLmg8mEMU3WGcneOjIDJuTIgtpoVIm3X4lS6S6TnSDeYyG1yypaPy7Txtz/ALG3UCUJIKjRou+x6
SabhQvX5IAIuhAM3vT1dz5nSRAlQfnbYL1dlzRFfsjU4ALuwBVjgrHRy8FEipIjdSYuXv9aDL5W5
A+rlhmukK1+wPdJx+j9ZyVxN00eUKTe0nYrMfgdX+2zr+jrVSPMuJnP0GIGyY2vOn22SLHFwcXqs
zc+EJ0N1YyVRZRrnMXuy3XfjkHrC/QBI91StPOdxHIKq0K8O4piQNXZXb5hsoHairEA+qx2ATtHm
t458Q8kkBdaQBzrhIBXwo5jDEwif3cUqdLF0YSJ6Uic5GZHHvcOHdelDZc4mkj7soniWijP9nYhf
lsvsC+MaUB/gKCcfE3y20OhgKfKMLtaxNV00BrdywSCXtJAqTlU6ajVGOPTfdq86nV0j2rAtNVRk
mPqEbaT4Y/gpuIWxIwxyFMQDjd3fO6Ny8Ozr0V694bdyLIz624ZTxYgJMg5Uuk2jXczvrVX9MD7D
gqGNA1y9MxW9yYITvtMJVoNqQFb+gcMaDs6XlQMND8uq2cZu08t1ce3sq8VMs9tgLUbLR6yfyhiU
5sL37onT/fdiCyEHxa/0UKtG3nIOfhBmUear24U95Z2qK7/LZr85Mp3jdsl3CD+O2XAUWgGC0bpk
/yhXuC9clDbeJgLg7AgSp0Yq/ITnNEM/Lde96Bv4ZspBeNt+Xe0ifKtc/fP4FSoWzfg3+AwQgu3J
CdTxEEp7DY63hXImaAH/D+I82Li2PBJqnHszmAA6wHZSaqaskGGrIiRvK3zVSIB/IXvrddIiLLCV
OHFOqADaRUrxp/KGacas6BskcUXgcvWxOJB1AsYAAIukNkR6LZY8/swLMyEubgaDvENF5pm4Db82
63dUu0tgEFfYQp6nVFoUMKWHSD7Hecrsx+HRvVz3XqhSvm9mSdqReA0foWBqpAS0/S4GRC3VhIO6
hAEEig1XphNR5s44ASIadKpwaZAIqJ/kKx0OoA7wlHrtBu/dwtbJWO8HZ70a7WQdH2h74lzY38y1
wsXmVjdvT0tBebqSGvKG0kyIjiwGWAph6364Zh51b3eHDmfqy/lW4fGGfojLAGWnhfgwXRbegUJR
MMTdzCMhrSE7cKpPUPpk1I9XDl45S2JAp+M0Hm/NPMNj5tZ5Pk21oWgGsn3hQ0nYbLbGgDsJO/Er
3vt0H6D4yu2JESZAgrTZ3INtwAITutRXjuX92CQKA5Pm2GqO4pQjQP9JpX3XuvvwWEx44poUDR1U
lNTyHjp5JD2t61Ny4d7jKXbiC6NfibT47HamC9ce3W/a1Sxpc0WOZ3QWnrChsK4cZ29WVCKhwZvl
IkRjMhu9BOrV+wvSEcBNYH5cqRbQ4TTxxKMHBVYcTQ5QG+Qdm7izgRTJKrdXFTd9bW4bWVsbGVSD
Ds7flY6YeeOKWuoLlz4iGXQd3rM4tnWWDrciZ7R814igdL/8/csfJP5g2TcfApCjuH5Ogr61XSVJ
eM3lDhGeSTgp3w5aW2xFWqVwgOBbnOhjhQtTbNlsAsQSm58aP4PpOrc3I6f8USi/oxJ+91jqpLT5
K2zA3XpkQ/CfHjPDw/gxdcUnTWiHjmMwmXry/RTDfG9UQzOHRy198E7l4M0jmS/Obywt0alNefq0
wztWEXLdFQHVRBBFP17FniPLs1yhHc+/m6fxHlpQGbXeVlMrGvAoV0CPq25BJDFT1HSxPr3XdNmR
pQLM/+rd2cXJIjXTJDtKuj67a3a3ndDH4/Vtngbb+FKYnCgQ+GUrDkm4L/b+tZFR4PiVqZX1qoQw
ivm1Drir3cFWxtEhkllNJae8dvpxd29qaZUs8ctVnwAHC0k3ld6Va4xsMuG+HxAI0NLB14Xq2j2M
zXiEUed0HRXihFCD3aIXgGQOl12LGhHd/HHBr2Lmaicc2TzqBEto69+m9myN00H5WiMvubh9Sbp0
Yg3kqqeGFrIemsLLR1ajim8SZbU/gY5dOmBundv4/p9J6TWvejwK8DZ4w44D3TGUI2TqIe66eAh8
T1Q61iHPQxRtciiUwlX8OM5wNFMhF+K68M6KxvyIhl2vdBqIcm2in7h6i1w/OAHZLNpX7KpDr9BV
5/WugHlUaQWDkLFrJLSlk7BVVxoXYWTgEmsCv20q+QHBmXJDX+8+slJIEowK8q+vP+aZmv5rVc8r
ydry8O3CYxBOyF9w+U2YgplJXII/OCL2pS4lT9KhJX2e5Bj/Pgf3BHTuYy74V4xOmSrWD+bFFE/V
78mQqtsFXKzQwkiqPuE2WFAHGxZvmEP8aWgdK3IBQW3QUrlyDppnOsM7XgXL3GYbl3vIbUYAEHgQ
1uAWIkT8+UgDWyoM1DKkSN8xW/963RjCsikI0vFwbYjuNqmLXQ4rCTSJA0/918KxUKdPVIqJ7htf
oCTB9f+T82IJZ6Et94+3g0ylVbrDdSvYZ0fu89pVYTl2NRSN1TXssPAEV6ZGRsonIddywoEZkAg2
YPCEfyApU2qBnIHZu++94VF6KX2KJNFYzX7Hr6M0INLHhGeWsOY8SWHc8+jLvJHpSxSKMfe1nSLV
TGCwYs4jekrq1iyJ+r08F+jGm+x3JkX/8nd8QMP7TWQOI7GxSoRmO+H2hx9+PJRDjzWGTEZg8fQR
o5Kg0jdR5gKwGMEpCZEcwL2PK+06flZlys3KMkkpEnG4wIjyhuwUtBWGDuVzTEjceYQ6LSZboTgU
Lw7QOoicFn7B5iHSf4O8cn1jqzL8Az6tby9fdKlu7GIYwNSM5Ye71C/fC6nS6cewbgdMynVVkgM8
wC/yW/d/jMq19xyXmmks/4YVlsGvsKsxCcxm9yBYkD3Z51zdjXZoqqpsX5QRJ5kU/3O6b982Ohag
eMwCxZ9VWycDQJahwuFx6M1q1Iyah1Lo5hBbN/DL6obyYC0KlRxvb8dbZ+kQGoIT+kK6U303ajX/
NRnT9jSageIP6IavKRpH7dsXz5h06s6ECE1Bc2OJmbtasr7eXgth1E9DKEBKLwIuHqUGhW7yqUW7
FqOuwyANS3+KF1vmc26QJMuxmFOZYxI30iBuFZ0UN15kiB4CslUfIyzubrcN7qm92Dw7NfR1snbk
reSMvk307ycusLqTgBoLsc/vrUSdf5R1ZrLnwJGBq9metYqa1yDjxJzbVabhLDU4ZJI4KsPsoiEh
GlB0gkFUtuFQgn+0wnKo9c1EGnvzcoHyfq5gET3F/mWfLrCkIGNva7MqEmyiTremZWEcOcySDA3A
TMSB6q17n8nV0w1S8YAWWKoW5YX+uJOIVH43kFK+PYMb4e4VDL0uNVpmftD8l8Bih+Cc5iua8nw1
rLPDqQCXuBj7dceRIrbGSACjaKH6fCzbVff4+LgyPB5dfN6HQndou7v5KqMPfXGA+wzHHsDDagmO
v/pTADDP6H/Qwu2JV8u3qE7ZnX900uuzpIn/88BRoXGOrGyVNO5v3aPcjAK6LE3q9ycIhIUa3R3P
1ExDTaEXw8sUEexK++2ByYNRWCelZC67PRmrcyki4b130oTuTbaZG4uLgTdx+DL5mLTkBC8xT6Tt
VuSU5KDP1cI8Zl72YdHsulXy3s7FjbpTzTFut/0a+xwssgzC5efRzWUlcMrL4U9ZeFPTMmFMsgep
0eFe9lJa5dGP1GOb4q/W0ZBsdfbJF/VYUvnOx/dZXzJCc08CAcXiWbug7ADSHh8J1YcYAlqfOCb8
33W+M80uXY/rMZxb++JFzVlagd5+9MdTvkx5pZpSPowgy3OxpZFDCG0+ULMFSc056VnBFwuYjmeb
pq5YboKFrTJMe66bhputuEieEQ//MfGxp47YtjMayAW1uGnXsuNuhZiadZZrrJ2I67tPpFaOMK16
VwTOHAPAeO5oo5Vt0at2nLkn0ijqEqmDauTKJTH1tT8P5309fpCJZWg5BLZP+0786qZJXBf99FG6
Rj8BpQ/EiOErPWdHXhdo2kbhDe4xLyltXYpDpjFSqmAlhEg/6Ta49wR4VVxtslaQ3tHu8PvW/D8I
+DxeOyBxK0lRa1Xh33lG81vO5FRuUIm80Ke1QSl1r3PCSNCM9nyrly/1mzq8hnqhMgUTqpM07IC3
hRLIc3DlUmYbgNGQGhFuClOST1LW0zdpJhNU/ngFb80aLk26KC3Lu6bUpyhw9pxX/yb++gt5VljF
nhoglUm3EaIVPU68IVx1w2EA7Wxu2PMMsym12QAPqLzjegsH4TsEO+Z6uc+3Bpy5/aoHGdNA6HeN
U9rWIkpHQTeBsCsI1CrAfzc1OivwtNOyYkZxrO/W43uC5VE7iuD5do6njLfFWIoV1F9/93Hut03t
LUdcT8rabnxsUj/dh+goufQTjK7Rgo0MAKWEUnTYmgtqoeSWY+IQleeaAsyU2ThKv9a/Wr6NU4xk
DWeh5PTPfUHnwiyInWWg8QXySDU2wtHbY7jhoCyX/GUG0a2YWIUjQbxBbQsGMP5rqkaBBo0UwdIE
YghagwBfJOPyngrW1qvswuS2ViX5m2wStlibxKxz1M5BVHhuTZouyBd4KFETPusNUZLevNx4pT8Q
flSsxjDg9sFzGbgn9/S5tC8AHKwSxzyesAk63W1xf9eg5FlRdur+Fo5CuKKGg/Isqvzg0HtdbgMa
I6yqM3NBL7MmrQpPfFpGWh/ch0btsb3EOxCWAJTFol4g76tuaI0WPzVWAS6G2d6DHp/9DTlqv2qX
1adnEfkC4xpoAMWH0gyk2ZtCzs3SVCGGkdNFesWe1oKMszeVOr1e6nyyqo55cT/kHvm573gYNFmq
kkMyPGDTK3p2VS1eSep/zs1mHpwEb3+w7F+Y9ckQKsB4VTW3FUq46EYrFu3+gll6Qqiyrya7jcod
Lafs3ZnPZHRfoWuCHcRiRLkqxHrWw1ZGaZbRziAJ1fKX+39jIA8FuDYXuANuRuu2k8gBiRHAbpih
ElK8xrn3/AjhHKETRPpE6Ym9XCcgkBgFXvUqUi8kXAuElVQfYOUBlr7RjydOPSpDNpnGPjcNzlfd
1MYNzzSTr8N98QCcdhGhTKvwCpMHDNFcU1ngPc3q3aI3ax4fj16XNQ5QI6HKF4fKKHaOt7Dhii4D
WoAAeMgp2vOwL1AHj+wjXeu/pKzLYdrowyQBOgVJvZUEPYKyYVxm3HZTw6IgDFx8cA5tjbGfUChJ
QONWfrur+ywQf+fhhWwbup5eOppVWUf8r3hlfhB6TUZz4ZfkGj8hGNJAMLSTabLl9Ogtub9UxlFz
kXyw/PG3ycFofqaHhimqce0cTN7pA3untpMg5Ab3Xxt5+H4GmOKBjdq5kMkixFa82wfDdU5hGfn2
XSZkIUzAul8ADLkotmhgP+1r9UWqF/sY9clNMez5nzdWjJqV05Jx4lKcBfOZfdZpBI4VazMd3gyR
EGa7u6D3NDQ5kQPVQfiqFtNXbzYyePwKAv+37FzncZj+SdPGksqb5RUmsLKFulGzml9E9QZeoIHJ
j7GR0R6hTOCXD9lenJ+bGxNnVFRvYWxahvjyLXAIDdGILSaMyCT3cfdbAmLP7lg29t+MczSzNLZg
QtTcWm0ts6aEV1I/MOrZbmgPl9U9P9GmuvNmjggpTNSeLl2aqo1n0JkQ49eK1oYodY6z2xjuKjY8
TbLofPwCbQAMg/cg35EKY32TgyfA/9zcI1PXE0sRiau4vodSGfeZiNgIS/YiBw1tIb1OofFlNCYT
OglptsA7Mj41wC9OUjznBcUluYB4g4kT7B72CLgEFaqRylXG8pc04r2a91ET7VJnlO9ZvNREyv61
Ph7oMeOGT3xCmkMfSJsgLDNMTfB8yJVqh4deNvmIVwPVZJ6xzapgXqJS+fwC0zgaRW2+dPec7WZr
TvX9HCDY4iMXD8Ywo+r9sTiuZY01iaZlsmYDmOhPYnTGEeDsWeYbkyrNKwOVrulIwgRxnMszsjuE
N1kO2mcVlzP0jbpFCY6SHqOMzUR3N7ZfO60F/tZr77VuWTBLX/ujJudk+SXG4WJue/mJOBO86DHo
PtP0fHj7Pkh2GRWBfTgNxTIC+fTS7voSxXZjin7shzAqqqrUiIppcKlm84FCkx6cMqxp4oy/38PB
L2zXluEE/IRpmIgw6AEvDeSfEwmeMR2TOx4+KB8ap4JB+srUSkOq9ppNpzGGWPx8LUbhZjoctOIy
MwbvS4A+2Zkj9wzn7yJfVl7HtRVjD9vCAX9y2xk3i/cRU158I71uJ2shcmgRvg65MSxzIlEOogiW
V+c4tih7tUNpWUfgzEigRzxGfeAXKPXO8MUA8TwLIuciwgOgXS9Dn1CGLtE7dvc5ZjlYaeS8rc6s
ADv8/YMzKHhzOdN4Q9ML4FHbmLLhFJABD555OsXOqB87BLmueprwKg3UfzsODDH3hUd6hT/ZpGZS
mlUPLzgjVfGtFuKLX5j2qyUz0ETeOOUws09Zn6swuF/QlV/NupIOZDX2wYc8zJhc4ANXA6SH4qiR
rpXlMoCNbQWOd9fUVzGgdFCZSLUza7GGmMJsVDGr9XDmqZIf8yBEzvYLwlMPtZ4FipoD0KEye/Dp
y6eUfDSwXlv9euhdiVvgvLImzoJkR/oYi9RLVT2Vt8KEnhYkwjILsAFzon6RSyVXvL8xy0LTLUQs
PW2aMi38fw8NDJSLamAkV5EQ3jJr2bNyptXHh4RZc3D76g/0n+EZ5xYYlseHZjJ9WhHpNyghXWOm
LsnX3ftrrwCfJj+Hb9feJDWxs2zs5avbpcwpY2Z8UusDwz+XgGAQvJ9q6bnAn5qkEkK6L3A0cQVx
GaKlakBHLBeLgjIC9O0XSdaRJlkd4L/GUQWZPaJe8npAyKYSlqmSlVOPo6g6cETnhIQ/lpKyURWZ
U0mZLfowTstT52CNr4PlFJ7Zle90BqIpz5FgpWK4OcKxhR2Mb1Lds30A97awKdUi1qIJO0Tdz6Vz
T2AtvXMYuYq51da7loiHzNXY1uLFe8kf9Pe0u0t3+fXMsfgsBJSpgXHVlO1NO9y/rK4drOf1lGLG
fNzmWxGGd4Ojk/4ywgp23ggoqPGGeGhxCWJeHlH/YFdmV6JU0+6povfbuzBqP4J2Bt4nYOIMxgIp
I6k4zoMNv4DmeCaIQFtHL8qQSWW8xCetUP2Q7BWkHBjugHJ2/LSRexdjkulTnKHAbcR9UAD6OJjt
VynaCuGu5pClc/hthub/dHnN3d6aTz//KpferMlSwgZLodRZChJjweIseMCDMZBW+Xx/jLmtDw8f
cCibkTDT0rkLDJCpk4S9ZXSVq5A/qM4jOyqpeYzJITF8K0F8JUbecNkTGt/NwGwsr9NmETGp3P2/
ozxvo3U42Sr4mP9GFvw5IQggculRH2OmRYIXKseTY5dW5rWyJwupxz1gqwBsb+rfmaOuZ30PPS8r
6BCrQemmzdZPl7T4azLUllh6heDoZPpUSG6sZ4u9wAZlk/SDPeeqsd2TE1OIzyWqCvOhG6CEYA9p
gwkW4XOn2NvScEQsu3afOOSsXi3TUA+S+UFpl81aanEm6v3csKm3FEVLIIXzB8ZB6251IHqRVTAi
Ecq7Bfm3HD8xJFCE3P0mbvbsQ/Ne2wZD+UcYIxo87kIMb0JppX72gIyDr2gTHDzmLvlG5+EYsBtb
NeFCYDbZyzSAaV00kybkOVxRHivzHgskFfRLxK3yUfdYDIrMCbVIm6XzKC91CpG8e+DFTzyj2dSK
spWbXY3G3+wKODXofsgGAForUWBwrk9nLiGvMHYa3+7rvVYuh5qFchWNxd3Fdqh2MuvJco1l9wIr
E5xxBtKgnQP3UfCkTVrNJEa6ibWF4JU6ZSHBe6s5NpL47Fx7hFFIlSWLuv61qMGmtyUbxYSEbWaY
SMs4pRiyzyhZ0y7vV3kQLI84a1Ib2EJC70KjHNDbr5mmaYyx1bTw3QsTs3749JsTP9/ybIPcNU2S
bnCXYgKnAD2U0bBSb4zRrEEE4cHr9AuZxHJmU6/pZor+AVaDhPANPDeTPyExsySC3vgXl4/1LY45
xnRGebyDEA10453ogzKRDP10acSbzYDFTGoR3eJYVLicqIHX/lhi8HWwPbSwactHw80QO6NMmPxs
kbb76kT55atnoAYqlj5fxHMZvtYriB9QRGWQzpktsQzS9TbJAiQlqUmBwheaw4VHCp/TC/Mznv9z
HwwAdIqGrgzvcJzalw4NhI8LUYeDMO9+6TN+O0dJmEhWTKa8c8fqglNXoIzH6bZjlyK/Gqml8L5B
dmtnABfZB45nSY6YEU8ygOIT8Iscmx7pQ+9uS6hcoC6HK8VJLCB+/k3r2S+E8jCmJdzTTKjzInFw
kVp5H9EPn9pXmQ1VMjJAmsKFn+srcYLhXjE9YRKHik4WiAXVC1O+37CF+39SLAW9I0778MgWO3E5
WLPHAXp+I20FDcH3+hQobvYHDLQgwfy05G39cEz0reZC7iTeKZ4vy1GVqlU0TbwU6heQuRpGDOyN
JY2i6G2FZjucVh1RVifOFDAi13p1/iMAJmqTyozplJkjYsWkIOIFG8ejeUI4gBELO4IZtoow00NT
lkARFzhLE2t07lymFWWdS6+GLVDxUaeMEjVBRJLSMRhkZx+knwEiDgnPQf9qHBzKqx32X4Kkf+6V
eLBKYKsOSA8LvWdYNgmtdur/wXabScJg67T1uF0YCCk+4snIlR4+PHQ01hMJhJnmaiRdYWbppHZ5
2ecFcR4gPp67uB57ofhOZ9tKywcO3UhQ8njyMzt1ZFY/JXC7ISBBybWse6L1+llvMA1mZZ3QOmys
UCKf5a9YYY6b+Vs66Qr37WlV8fIoGDYijBJf92JSEXkNnWLhvFE7QUbXSPqde7zfw1T9xp8sb3Iy
oLIoJ+0qoJ5R1+3Wi/IPIOe1TtjJyXThDiVlI62oUvarRURwTMZ9axmECZeyT4hPAYBoTwqvgNnS
f0ZF69Jt0lS+KWDVWN5E3WaGY8329PAezv8/SeyEJ2j68FzGGPFtiED0biusH3auvYgpkisyFi4V
PyfcDhtdrkK3+rxD9Wk+QJJVXqIrO1AFN0ZNqJF6Ca4DMYPjAE3txMD4VepFXRPV25IFcOfyCxYH
E+/1v00iSvC+sarCUKHfRUSM7igqW+8chGt65rWORmgaiHjx31rAwBaLiDE5Wq51YP5Q7wRqGH4D
BJ/BZ3PWL2ejCuEocyb4cynQv4kG8e3GDwxtoXCTLT7wQyPAhXrTvyuqLUfuZPT+++0hkZUOaSy7
Uqqm+xZFI1d0to8ANL97RpOorzOGiJ7gfhsNFUU7h2VS00KrIw2GqM3t1/ZMIPnhM+yZn1fgMwyF
GXotR/uafr2rMVYwmVDcEYKP2zwtIEcDQpSWIy/q/vjc+GQJ6g3TCh64fziQCRTqNgsc73Cm4xGI
QFgJ63IQCJ1msp3qUFshIZMnqr35gOLi8EpQUbF1KrAPxa5W+46eZxxMV3grbAGoeN7eNieSCYWa
Mdtar078QSkRRDEL4clbbsS67RLFxhQ4Jd+kwIOU5pzYfKqquqVCtFb9BS/XKkh7bGzEZ5pvMSaT
VosHpporJvdcmfgzUvyZuNOVXxWEv1HbNLba+kQQ17HFwtUQXclAXlyzywKJBvg3T9Aj5RVtl2vG
euXqAYlOQhehL4zVaLa4mgKo0WNB26ePw3L4E9BkGVn4tBuRdrvBF0uxFil5e+5J4CVOk1fofhKW
odCI+Gap1dChhcjkavij7+RxPz6RThxx6CeXbGCkpe0z/8eslzC0xcCYmkLr9M2hwCKRsprBWxXN
pjn+Hv0aVvy0WKRi14yoRYTCDoWI5g8WED8MY7JSP5u+/cX1qY/+dE1D0O7+THNAleR9Y5uoShxT
cY9xCWw2pyvxOnz/igYpUZuVdFLFhL79MENW31HbKxm4yblMtWGZT71sGkgZUtPUuvJrU8eqvIkW
P2dYrobe4IYQ0xU56j5p4/a35AQ6HFtFVnWq8GTOQCwzN3YKlvM0laNNf1gfZk0YzF9/FZs6HwAV
+3YVM26aQDOoMzGovTSuxGO8zdeTP70cghKlfI4cd5JnqkwVWC+pjB0iNujXojwUJG5hP1U97dl8
0wHO3eMJ3Csx3TVPMwRtsQ6QriDN0J1bkeenN5vVDlRg5Hbhjw2ZU1eQSkqLbK2/WdzMVtqZGur7
WDxDrikD47mKBU9Z8Lo6YaiMtCQes1yWdWtEJBwteas4cXEQoDR55EiGW3nnJwBsXO2bmTo1Rd0v
ebDzrJrG24kqttP74Fy0iIppx0UipYseS6tRKAaiGC4iu6H2LNUD4Lm8BtZgB36sLM4YLd+NqUKS
0ouw09gNQZvI549Wsn5EUMDaitRtDMgGjC9T592X23EJ/AeswKzBQV1S+b6hZUA7UoyTaD+8trgz
e9kSUGjuFeQxCX79tFV4AK0fM9D3TFVrOLeJ23tB1U8zHwMWwjXN9PAh8Yjexuodnmlq24zQu2Nt
lAOlKCDYSNxatCPnzQ5UA4gYqAdpJBd2zqD3/v2OMmIgTfbETrYzfXnbiPVnQxyG733w7ShK5Zd5
1wLSisHxlJSKSrdpWJnjQ0VqwX0rhRysYCT6jjsTwoc24P+fkfMvGRF/MkSiTFNFCazq7/LXCRf+
meLW01TQhAfPBB1dG5cB2SR1CYx5Now3lBrFYgMyV77yaWHtPb5UiWXx9KAcUHHLDJNgfQkAVSHG
5kWkzesOxW/iojC4IG/wtLJjht2AneGM0hKQKDhEf8FXyEdMJRFdtOD2IwpSamr/euEKUofdGehl
zm80ogZO5prnjTSC4eHrw/2MhNLc1TKvse5l0lSWhgIXqHyTUQqyFRu9WP06WKkfy1pqghctdBQA
LhQjxYkZFpFOutJBHYxeWvlyQXbTPBafamEyq1FbBXaYHUKJH8dBC6e5xy4lZ86Wj/ZUCFZE04oz
axVwKM4EDoNAsVGIEBUdQmAdDsMJ7BC/y+APw6mAyMn/osn8NHFDJpT55u1WGUG/Qa0zDRtsbOuA
fJOWBtH9MfCXLlrPPjLw5ctz/D8OqGeTPKDJzOQkM07rH/udEPusZv16SKQoN15WI4VYL1NRGn+Z
ahsIRsn03kvckhPYqdRvDh6GJ/hqJb2TTjTemG3qvueuZiGNjw4YtiCInzJSWkDcXMZwzsNFLZFi
ODIpG6JdrRroPo2SvQpqIhfyhO9q+Gwq5uNDxkqeYXyGVEKWPgoGkoq542x4D0f+HIF9DpiaVSM/
+7mA4/Dec3FCVS1afwtW29SARGDkPTh7o8lP+br3RYSvX5RkM7Dk5nViOIxS4oN8rt3LXoec5gCY
qAmQA1pVmWLaF5zAEoapJWbT+ae5EfFKdxFAZVoSxg1uo7VLHGvKaje7ZUcTe3LBPMj2SraMPdB/
dMiOSj9xYWW3DMHuJjN4jiu7+YcYtZ6x1Tfpo4s3Tsq165i/4H0GEOQPwpVXE9FXICV0K6K3t1xd
O/CbvAC86mn+Iegdw+uo7ldE6qa9L7NGwjo5R4DmDpsBNgKIOiwjDXegUOpRf9HDoXqkYySU43D3
IuXRdlDeX11X4KpO7RBk+VTd2sVYAnrTjmlnHNIpH3YKc0Pl0WVK4aw7ne2ofhEplSFuaLFW3JLK
xIw313WB8fCRtAHR7o6iDEmMGp86TVvQYkj5dnexFMFh+XCCaYKZAIgYYi26zShMceGEiSq0krxh
OK7RO9XC9RtvSkNTaQVzusSiKorXh7Cr+TLYPrX88b/uYiRm0wo2nQk6Glu8QM0VDpBea3S23QW/
mp4ePLDjyEchKjZmV7/4nnAZArEO1v7/NEIgXw5FonugFjZ0hkvMCFgdhWzs6kQdMbbUlasIGNku
MdXBgIcwWJa8jnnHkgPFftJkYmhoFY7EVJX4cmfF374sr0utGu9lmpKmVJP44PSjjgs6vsgFv3I8
ZmZgFPkGsSzvVQQUfkKQcN6YZaJ0XpFolXc6wo7di6fFn7h+HzE+8EeWWJvaxqqDNoqsic0M/8bK
0ak+n+0HnWBnC4yhLnLF4dK/my0qJlT39lEoagcjO61x9HiqZF9WhAOmcFYGmWfyNjdpqiSrmjct
XHtoXF3MxVmuuNVPdcrEW4DXK+ePjSzZOD8NScxHgP+X+x58EQxDULW02e04Z80p5LPsJ+fPE/vX
ATixk2PD8xg/IyM0E3gTDsKns0S9OGAakYI8bQJu9ibhiB+crb6/nEoPcEtaNnm31YB01YUhFsiX
8oCq02TA9P4pA8mvF1ESxottczBwYnDvUUNU0PA7iRefOqfmyNCDP9wHPfGJV5U0MCTaOlRfSxF4
YLoH87jIi8DrZ954WXmjqUdIDKhle6+NkI9aghtylmc8EJckXNqTmPj+r8lS/yRSu46ZNEmJfj/w
19AXtRTGI2kS7TApnaXGtvdX5PQwaznEiKhdryUQdvoAe+SXy1zKZ8fxSbV+iHi83nmtMKGHHydu
lD66znqmmUKAe1q4wPUPY0Y2Djls+WgN0DnyQOJ7nI9WWXK/3zLTZ8ss47hm9MN/GPW/bm5az7gr
FWsIETOHhahFEHmKxDpw+sgpLn2g/N2Pw7IJ8oBld3V6j+aOc5E9rD8Ki0HrjMQtSxggHn6teM+/
GSNxqBS+uzfrTrgteP0ltTKpiJgMmbQ7VvXrFyh3r3TyRgl7fwr00eJkcXTyNjwc14EVFFe7OS4J
G3DAA4qb9AgYALGp5S3f/LBGHQUPaCKEKX5Ux6I6fRNa4RIfzA1NgwDRMonSq518mN6x+ixbE545
5q5wk91Y5T1oe7ids/AkQPaKP9D0Dgwxgwwvis9gaL+LiGNstSTyHqpQ5Fv7J1LLukH6MoYEULzM
ETdrZGd88Ea7M2utYIXqcyb4X4Aw+E/iFbR/UQNlsZOEUFaEPDP7hwCYA/CCB6BPEsVl78lB5tMq
OKl7veDZYujx12l6eZA8HNC+6XdCoWGHsMvQBJBXTdz9sV//r8/ZWg6naeIQopHZhNnX1vkvXHY4
hdPb9FFNk6h27LxtfMbxHRvUKxeVyBN/X+VjdYYH7tMBuHDs6irYJ/mPgEsG2cfIT8iGzqJSaURB
d9+sE51Zdn7STJEdt2JPx5t1jeniK/7VV6m0qnbRcSSX5DL0rRp82TCkwOY+kdTF4lGNvx+QlU0/
nL4Uiqbw/F0nhON0A4Mmzkm2eo2Vrbt6Xvq6G0vJ25psmNfxZ/OoSHU46IdJWLuOsq0QVuYT37D9
1CiiK0eATiG4m412GJUo3KL6jN7nYZ0XjGiSC0AeuByrvB5gm9HL5BHYiUOJKSw6a49i2Qq38hxC
w6CgFll/I9yYK7dPJ1Nj+HMX4MgNgXrjqGAvynJRo7Fwt9uDKNlQAnclSBTJiWLQ5hmJDsvyJoBn
DtKju7nJTch2HReXGeIlk0ojmutRKQRM+tx5mMjsUsGLLF8ubIP6/Ddw5DWvW9pJlOkKbNMNKq+A
hUcNH0fwdXzK6eHOpXAO1WOIzrkrbUWiYMx9u8pExUQ6Fmesw/UV63/RBT0gCeakAzQapEXvNa2O
yCsyeFpQgTiCpK8nkvglnhiID3t33J3NrizXBmhZsKbs4NjoO4kkrTtT/WW4C8XcQH3Yh74DJVST
VC5fO/6/eq/aMkcYNLwiZO9gWdgS8Csg/QfDeak4vwhTuc+HM84hfC57TeXUQVexSHRnTGtSfrxd
FClas8ovOyw+zg9llLZyujnEqu3OKMBWv2Az5Eomoql24F6jfaYJ+LZKN2lY9aKC78EsGRRwmXYd
VKsgeLnEqSx+ZszMUFyHIIsj/GWBV8xR9VuiLwvB5ldCtNzDEx4i+Eq5QsxsrOuhZgArgpDMPv40
O55r5sQ9uWWbU19I4s41wXNxRLZ0BDun6Pyi/GleB+2NcxxopI4Aboqenxh3HwXV6SGXaD3vHuW7
4Ig4IcCXWmJ3GcVifgubnYrGtdQYPcwXSbYie4GvkfJJKh6aSDfE2GFd5ZZ5FuSkC1qNKQGRtgMX
gjFrRJLzEpChx0YyVKornf5rhy4R8pB0rmO7TQ2P6NQUOtQj1+aBc4jx2yj7Ds2sDkBnAcnNLBV2
DIhMJS+Soro5Y6/kauoy/PexvmANE7cizYLUcm5ya4oEpyfFjf3smLCLcv3Zvgzo/5sqHdE9+M2U
2SFTRfU0WzhDRiFBRRtJ05QEKbIGccBna4Nz2zGm7BkGrkZF8Hd2OxJFpmd7MfYHoaWo1GErYAIl
5OotqF+uvIUn8CjT8erpsJBc5fmeawq1n8UlQilHemGIpS0tI9M+OIcv5S+kn7/FLgz8A7SGbNDz
VITBccDNFD2znGYppsUGP7ZGDzDU1XSGwFgb+iXp3jzmIGhBlsxsLEs5LwXuQnJ4Fxc3nWFoBWJf
R7S9LRdUPh3XO0327lOCIeOfJPGMwiQYpW/MgSLpFO0qMPxUEA29V5ilF6D7xercugAPAcORV6An
tnQ6BzeTjmy4DKfsoFcUU5PQamh987rluEbmjen451rEamOiL/yFEZUowWPKwIqi+4moTQPJhsSz
/+wL4Xd7XIGXN3jDCvXu99XqHZBBoNqisiYPsktbUA1yTxjKQb/VprJXRHD7aRpI/Tl40uRJqsVI
HKP0ZLbbiwsBlTsth6+Ti8viPK9VlMSZpig/wJpSFCUEwJDl+Cam5jzFrfJ4Kx663CRZXxrygK8G
+ob9b1NErY7N30182lf31Bvd9o8gPdtPGJzYPq56acvUJBNqj0r2JxdyrG97UPtsS6kZrB+YXPjN
PX16s8KGGluozH5ymRtl5/abT9VSUtAfZ8MTM3/LNOKjxbfsfdXlzBzhqJ0Ju8nRNuhB8ATBmUFi
GbxV5Iyat/CycKbDe/+sEs1SFHfnhChiaqDXSJOzsYXKUH+7Jv7a5TN9bJJKLv6KptY9kwXRHg4d
d0Isg4qqZo9t1QUeMTSTBu6ZOtMB/MXBC86q5ltUNBKFq+GdB3hOG17fZMeH2RR0mDWZ0orMrSVE
zVgLdp0RMKB3mT+E5VUEYDCLN8NeYyL3Za2h+AP/2KTSj4OS07J06y/qyWd6iMN7I9JseBpKCxin
ElcmE5RA4yiH2ETxkS/TQJQdzplv8uAIJICTn6OjKd7zMyTP6EldGwdRw8/b1VuncSPAIJv+P4H+
ZeTQq3Qro7AS8NSiiTMp2LmLQIZEr/tcoTCcF6vQkWrB5cRzNvW2wUzfma9otpImVX3T3unvVjn1
7Lm3kZfoomsLBsh+/ObUhIJ4BtM25+9vgzUCyAMbLkEHv9aNrdwTkBwF0J+pC3Ie1IvZMWaDzQXV
2VXxljzrTAAXPQWXYV0SlgtrAlT+GCHhQKPXx7uLutxGcvzbu1c1rpxytjvYJDdz4gXWp6xUKWuU
8GG0oyJ8H+0+Ork+HYnskecRELCWTA6sdd+QerCqld4+1+YGrH3ndcxqcR/z46z3FywRZkWKuMqM
VNQCNdwKINbvARoHIjDONV+JXVV62WOPtZiHM3LAObJalV/IimuRVGZbdiUjcOtqedsE1aKwIfRj
Fs0hivLeyXWYlkjNYkFSCHcX/kyxVBjXcztSzU7CPuBhvKxUwYNtJaEUbzc6sFy/NKM/s9LYHkrw
Xk0l3ur3Y/W7w2um7FHvP+1BcGAduztxI/6fqhsrH9fORFR2xbO6BL1CfZpesOgr5dZAxNraqHYS
L3mpNmQc6nncdyJ5QlPqjgYgPnaUOG4G/Kt5ZRR6gZaVmNNjznqTIJvk+ywxZ5NT/YpDkJewvDkb
rh9k+PxMNbx+3hc5l8wpI/2ZOsm53+pO3TwMsvfuDFXuJfm/VvGjwVP3lOPdtYh2nfwmQzpvSgDY
wFp77riNVAMyOTfSuySWqJt15v8M3FF144SR5MW/0okNCRsTIFImDEP0Jt58mKZgnMxlFsgkYx4k
7Geub2ZwDipbYYAn+hsNb9OcEYjM/459awJk4NyO53y8w5RPzBTyzEHrqVTb4FAd8gi1sb1glyxc
FlLV26AFXGueIVmlVQ+G7T6hv8MRXS8mRvCFGNbDQf6N+jOFEzXMBmQJqy5+Vl2j4+WH4S5uGcrr
pEXkOU9OEBsQEiGqYriTZ5CIvcWE/D+BNp6A7GbHsLzJje2qQj2mevwYaw85/PMIXlquuAVF/uqF
iuL0l3AjBobkIFGUpEGd2a6V1FbgGCRg5xaoYvr7SH3gNiLGYZtodzo1fKh8KpsBLVzdw+IeQR9o
gkoxKmY2goH6/drf7F2Y6UJ/VtIfAGE3DdIL5bT7o4wBwmdjzo4gqVq3fFy16tAec9CQh3qlvG5G
Czy1ErVE5/jXwy52MX/gv0f5Lde4cnCD2ps/zkORf2sFubAyinjmsQj6hd8D7rCuQKCYYPpBX4rI
6cTbWQxkrYkDFxVKL1s6pHP2wW/eeCiaJ/W+in2H5OQKHKLgjLksaMvhuMk8YO4w1TqiQN8FTg6H
41JmwlqoBu8yl4KF2jLQ8V9KBC/Vhe1cYkSDiUGkzKlqrd6fNgmSGwxtFYoqOppd3oesylQKNAxo
BBcQyOGmubjnw+L6gOWX4TBzLL3QcfJlmMEUvXM6fvMB9+zjQMnQ/aeo9OvEvGfaazqIMZbMZvKw
IXhjB4BxqJW7BYmjOW21Eg56N47+fMCtxU+235vHH+hs7XQGBb2GUTK9EWO8PWWuCwqddb8ToyA4
uGmFR0G0kxMqddart55nfJd7NCipGS624wn0qMroP9/Un9yaMwV+mPxG9J3x3VxJ6rq5ZyhcEuHw
VQxUJab4P0+tQbP7i0pL2Y7U39H9x2daqp4/BH1IEwS+6w4TnO8IGdpN3TK/9PEWsKpfnVGUnRIo
W4xEyieswIVrdnig04W76ZRm96H4kg3VwEFmShT87bcV6N6FzI8jdgLk5HqQy6xPI8n495sbczgi
6zE5QLVYn7q11VHBp90s3ngKrvoqUQlwwyEbJtKSZPck7RhQhWNysQGoxPzwpNgeq5TMgA8Qe1ow
86dGQ82Bn24z4dDRRpUuAynEUfsCWUNkwxxwhf2BLF8Dm2FkH6AWwj7FoBL95wmyGslqOjKDhFet
Z0Ym2A9+c+ULTqPCypQUA0emCsSQjh/Vd/H04fvAD26sBomiyTcXSn1/mnQ2QEYsLfspUOHKHQj+
1F1ju3W+DC6HeZ5VwqOvJIOXSvciVlo069GDKUDphIj2cYbbQS0iWngmqw/zEUYyK765eQaHPnlp
EZNDxy+sfxvRkJXgR+9Kx3Xf7cTAXBy8+pYdjz+PKhtZcHmXxPcXEQgmSC+rdvNxuatWK06/YiFi
Wy1D6vSaChtO2WTb6dEXFzk4HgtPxe+2um1K2zzPBdFgbxAT4/fT8BFcMJ3sA12VRwT/Hg6EfkCc
IjsQ6LpnMEHCvey0jONRir7U1DdV+w/O/U/HSZZRRy7hsW9+t0rE/JtuVFNaYBzy2ZU9kgcTkgiI
m0XsiF6nB4Rqog2LR6bAQX1QXs2IUFjanoUy0FRMXz71BD1ZYWpp9kVYWzHGqqqwMkuALF/65WRw
3MIsOPHrD1K1+NCKG4L5rGCCXxsziqqM8WEWr+m23HWxym9T7HZI/3D8Qhx4CAg31XRjlm4H+03S
y6XMWsJ6vgPTs1VDM4qyV5gbV9fqjIwkE0oiFHXEmPvyBxZR5Gc18IPb9y5stKnSjQzsU4nXDTS/
Dl01g4Lru3b1zzKi8aCtXj701s73gApBXy8sxkz8BRyM/LJqo75E9fhWNlAG61dUOGNO3kquDJ5I
D2E5s7sXpaFTlp3RafqaeEusSPt0UCemb4TWnUa7+hZkL/ZsK90HCiyIomw/UJunzB35wBZ4zIk7
Nfr/xaSrt5eteEhHoKJ4kp7jRDJuS+nQtXto5adj2EZefpO8YynSizpHFXn4Bj7E/U+94Rpc4CgQ
oIbbi+8sshP2Ga/icgM90UbsR1bh5OfDhk7qWRtPXZzv/EfsCxI4n0gk1hGjZim1am+BMWuorsKk
3RsRW6srsE9CPMcYEEo7fn2Jc7J3wgvs9smKvYXatcMgsFrij3rIGTuWtPYz+Drm2fYoxx/5rbht
r0m3vL0iWnTMvRWtQ9aSdyD/C4LEivdiz1X5MwEoRfTzooWUnj2s/G3c0G3DlH9VXQ+e70R5eehy
2mAk8sJIbs9EOEghJdFKU1ER0BpL0eHsX6uDFL8rF4ah0Lz77kcpurWeIUky5+6VQyaLlIz3ZM6v
zLM+jfnIMHizpZfVmN2DKj/LyCxb6Hz7bneRYlSrVDneeesX/T7lNct37HR2F1vsy3M+laAjjurc
/aTORI1Ri4kdUKDb9a7+Yn0Kv2xBBD0cInGlf159tgcrdvMtx+eU5ob/PN5PeFH4bNIdOyCsYfiG
mjmLnm54xGyM5FarmvqcozHkwL7vOYCoLXuhKpfGVI+60VayeoRgs/04G+7EzdiC7DkBUc2WaXUF
JQlty6m2ezWd262z6aFZEOeLpxI7Rh5sU2F/bDpVi3cdYU/I3al7YMv4qVxfues2Wxmm5jFtVrHe
+hE6MLTb/nS2zL23Fi0Ssv07QEntNaU2sOX4gaI03eaUGr2a0E6rNxoHJfF/EE8rSmr1Wqg0qGZ7
adCjWrLGlxli0KaMMueqSc3IOVCGco6b069B3SR2Ja0CG9H/X4eDDZwxAmV7xNRsyS5TrOy3yxwR
yZCPLnxJLScOSgybN5gy+UbYBWb+pINUnFjGdVscvRldirKQ0MFomz1LJNoGmRJyv63tcRgjxYPL
6a3CKhdlDhK4sDXZ4Rvta4PiHsr2zsEk/zKh76ONiImZnZoOgVkbbaUx3C0Ymhi9Aft2mjX6acj9
Rn5xSgTO1A+eH09DrSfVK6Gfjwx5vw+cB5FnEMEPiF12AbvHQS0s9kStn13765aTJl0iLrjTxiKj
Tz94JQKvFVOycCNJb3KcngKHJSFwYUCkY/F8QFHO2VOscxIaagMpE2F58n+Iku7PtWRdIRopUQxo
0v7E1oPzUYFLKUsDXtUH/GnprKdUNIestNaKRQvrGRE58qkCfQ2LauvRnvnWJQDk58MaB6/9sTIe
lgaSIx3uThHvxHGBtB6hNjmj72ih2yDz1YkWkbrf1uNID89FbnRcgKViBqIaUWcgzLT3l0Y3WcCk
vHG6bbJP7cVeKijz3TXBrzWhmUp/UsKq2UTKy4ydrmRfogsEsYLCGKu67yuHzwy96k9nRIiI5GBl
0EYJuv/QatzyP7IPBIZ+cN3qpCr0Z5P/r+ix8hgmDM7ipuHHERvUE40tJZtsnQ7lLiM6MWm+WZO6
ewtQNpfol5xpqH6qLc9E8q/I3ubGzDTqU2A0FxeaA1KrbckXF71anROcVUlg8XT1YdMtjw3ssWnW
OFpArusH+nNqfHCmX2B9dML5t99JnyXSqe1OGaA3z11ICGBTj3DEmQUnL8h0HbLkT0gzp2OYm/Ui
FZFleS0pZnBLXoSjoz2r5rzJ2k1DuZi4mP+Jt0ybPhCaDtHa07qVkdQnsoR+bF3HdoQcvVVO375o
+VdIE1p/nCHmHFx1AcCACMHYI/TDchdz3cxETRalYfZ8O1/ZaPBoOFDK+7eUhxqVfB6/qfumMsvO
usDOJ00SLkYDU/Iggt7qW8R4RUuKC9mCITEuG3gFkOWpm4/jNrdLgxPcDHGDOhFZJKKbpU8YpMQa
SAUmnbUmPvV+B1fYT81b9htsbgMhdpFM1bXcEo/QInAUnA/EjHwg01XCvxAKRiv02maYkx83BAqD
W1JbMlROymQ+1jlVYBicjV01AHsytZLgR49nx2bUCcTZ/ZJfrvUO5NAPZy9NywIpgATRNXm21iPD
rxpavOQJ6cy56PqCfY3Z6JHC4POc2C0/LYGLKORsu4xuj5BGQfDWJUQWQgDZokLA7bPcLiOOfBc1
yMWKaemIQMmh5COEkw+wkj3kRvstp7YUWXMgWMGREjsmaAr7syavNddMwVnC8oJHFZqrw+7BHgio
odU0/mn5fn5UaFLihHOvSGgZZXYVSDeQXEi1zDJvSLFF3fsFxPgs87LBHO+L9bhLT3zayFc7pog9
xgBdzJdLOMsfJVjefVeRfiHov4Aezp/DkSQKcgVMB5BvFzA8T2rTudb4plUhiOUmWjMXST7sa1G5
lGLPYWWQdYUHDKArTMeIxherFxlQfNkYdva831mR2D6CSTdgRWG4MGumuWMkcpmskeiwlDiL1cL8
AfgR2NnBe4JhSk3s8cEzFJ019osRhMAfWfddH2JvTxq4heeTa6wY/M4OmOQ+cvpi00WZWAuJYbRX
NfV7dkuPfJ+HACpVKbo+mMspNfsVP1NWQbYMKEJa09Y87sX8mqX0dfBF30Rr/9iiIIie++qvBuQ2
K2V7c8vdPdZcsyABE5LOe5g65+oyFMtQNWl7BtZV4I6mJ9mPBai+gFYUT/ly+i6nzxPFY1R7iGdx
y7GctjcDra1u3Nr48BaJkna2oLNpvRfAUfgBhzeKUK7dLDTkHxWe+1HpmZA0EBaBY6anUjyoHCwd
idPM2BLsgIXkdjzzrW0Ef01+vZgUTVJV5Zlw+n/Kryc+dKKVEk7i1Lo2Zw7+kZ276c5LmRFNMtbD
qeYCwhhpcr7yfkTzNDxganIZQDLIUDLJWl7Wl5lYEA2CB2EI09sS8qufYMJJWQwtVYYvRJMTx0/u
QQGVmDMMDNh46sHJgCxaflleIdIMHFvX4kQZVtxSpZinIR3eye2MqDNT1u4nVoxzJkCeulFS55E5
hVsy8PgNbcPmgaxs7jEoYBXdGcHrACwAt8Z+bYJUHyP1ZHlToEXgbxDaRCFz2JgJ8VUGZkryeL5b
/oamc9W9QFxEDDmmp5nb5zexQkf5uIFOppNAHKCy3hYF30XChI9eLcCp0IaBnIg/4GhYZHSH0oeW
ddZUXCID0k+LR/1bDXNVuFcngxNA6j2njFsnkcDhsHPT4hh5IyCPrKdtrooZ7lCMqC1comrFQusE
C4SoXnMcl/B+zpn1ieAEw5eChfIPINYcJGmVXePZDoB9xBJHRVTOkoLwYzX9pIwLMJGj1ew6369E
/X0ukvsK5zI+RmjqGB7lJJBk+Exuru6FHEObtOWKlkKFNXVR7t85mYSEXiTL1WmINJUDJTv/cOzo
XWzQZz0JE9bcejpOCHcDIlqgSieTgWGO2R8NDiKUmS211XI4wpFxLJ0rJa3kRO2P8cWBm2K8GDRU
VHkbccvuZb0X2O4CRweACsvGrO93L9ReNzvI/sIsRRCcBUtnor0LRjAbE6u+SXdFfspWpPdfL9F+
bKvgUWR8mAv8MYT8RJDY98l+j6mgyWHkueHmaa0VkpJzZ9MtP9+yq/C6n+vkeqUVcmWxRB7flNGa
OI80czXCWwrqo24E7g8IPHVVnIGGuBb0F15VSAwCix+HmEm9q9/8aZJ5+bullc0uvEabomuBMUuV
/SjN2wxXvO0AnFvhckQNtZwyC7YRGGaF1Ou1LJYMTk+JI5DutBvE6uVu2dqQ02imb11MXN5BeUFu
Rhph0f+q1xYS9A8eWCj/MN3B0vpeIw8gT0mpAc9OhLt74clxCXwt+OOk/2Hk0OnwdsO6UV4S5KVE
WQsPHIrTAo1uWM4HT2ccIWFkjnUXAd56tXSKImrtRvzNyc0qH8Bo3BUGsHSp9H1fxkPhlTvhOe5S
stEpZBpE+K3aV7qh87CM8Zsnf0S+h2vNuKsDzjeFri7EnsmkTV2FzmSKQZmHaB8hAC8H0wLV4z6A
3s5dUnYeDhNjjUVOpm4xcYfE9STFeegvEzJefS5Dl8HVHscdDmFLiOLv0kaAtliJoLOEVRrNYLT0
ExqSaQzJaDGpDxaR3avosG8Ah+EIiV+pZo5GmcNyKku774wp/9FyvXigfk9NePKWNudl+ufzvmdu
RBJPfwXuOkcr9yKbrnsa5vix8DKZMiqL+u+73zG7dfxYQ/MxTgGbHauiuSp4DofSdpFM/Kk56n+U
4jm8qbKORSkLd8bLdyx3ioWYGI40Soz/66Ya5YXJ+CrjN7wXBanH7iVfjyGtBB7gjoE8b937kKuh
4XlZodMxjJhx8+2FxHsShpv5itlay/xQ5BZsdN3ppS39CSWwFK21dybjPcv4s7xOQU7ZytBKA/cJ
UWBENofrMud9tnY/wr+I4nxme9PVtXzxflmLd6sJDM0voXdikffiUWMxC504MBvPjkPe4NaN1TI5
+LLXqv5YeBm9XGlXm28F6MHqu5JEJCEhtIHLwjieucD3JN+LP2eXy89G6Cp8O38zvJWDVNHm2+Sj
zXJaQs9zz9RstV7Y7cwtd1kDTj+eBKdOc+r6ok4r7D8XyTOAeIt6f+BYhF5GCoNSChmCvsnmMII2
NI3rr3TnQi8xqdyKq0hQZnDRU++1po7PATaL99KRUkg79YXRQXRbkZrxehN6y770HeSgCPqrdbSF
ek7xfks2aVi++4FQB4g3xoQmKI14DByFGL/jF0Orzk3SWrJncTw5SiwxSpdo2PeKHUV3YZw+1j3D
j7xlbtJJADWE0+0T7fMaBmAtrIlrGn8ajvEG492D4nZfqhLOqCYgwLeZFVusbnRdE8C6xRGZLXCv
GGHVmjatWHDd2o/ZOFku/6S32hkMh39/lLZ+U1QSDosNN+y3XPZ9VtBeRUvUE+R94S5oyhVXOiWX
9MZ4oamwJ5tfJIxYZonDaXbdXuR9TCANUzBWptml8uw0Rjapp096JOsm+oV1hdU4o5KWc4WGn5HR
2AKgEsLN5JkD4h7pQVApbydQSHlZ017lf3opKeQmVr6cXK882LsvEyvs/NsnIFHT6f05Y2X1LUH3
pgyxQ39DlR1xwjoseC3uFEf3C7iRbtXkLoOIXEXbvO2P7KYLxCDlHJ1DgejbCht9rUOkHup/wqCx
a2o3n9wt5RIhp5GRn+9iygVAo7KpZaJFQhIqd73bSiSLo74xV8BnAkFG0R8/wzoHAyEcoqA6M/FE
SJ4vXwoO0iIgccyaE4vp/T/M3a/Ys4BqrrAM2Wsbel4InzAFMAqIKaT1JGGXSwS7qH6Jvarz+nCe
XJDB+p7Juit/5m3MBDVoFCz7BZOLUFYuD1BdhY0pKTYah5XPWx2RfcpwHgNPJVCz4cpXIFTMdWvB
zPsHv22Pt9A212nJbPgkczmgtVBZ7UMIp3PndZXaz5x/RvEgsrtLKoSIC/dAss+D1EtD9IEIFTH+
GXelIC6Nkp6JAgmCGHseFIs4oA3AKSwJNPq312PqNZbpevzaeKC0Cebop7ViXL9XyEAu8siZgKUI
xoNKZsh5d0/QIySoiPISnKm9terQbVKaaAk5OEf1rQwEOg4JDPFJVbMvgpHu4whYnDzyq539OyY7
ZvNp645DVDEIrFRVf5T0+LLHeOLxvh5VN9HqdLBknVjWSWOjwDhlDHYIF+y4XB5kyjnyMYqclOXM
+4km/ORbg3XDYtTgsfxNJe0Gm56+1ni5egM4boCjAZGEchQ2V5i+D5fnIm6SUPoNWbw8fb+6l/go
a1z1BAhJKsIurgUlKsPWdNahT7WlM2jz+h8dbqVQUjcrniuz/+sYeSv5GmGXoJ2m2d5Pa6Is4Xtl
yqUfmc18mosyOOcyFMPvrhn4v92T2RzOUV6pfP4NU3erEcVJQaSrworZOHsqTvTq6XHJPFf5WJaL
LYfisZF0t3EgQbD9p3eaxKGJVK5tJN8ZShQtTSdARHzrA2UKJKZhi2qESq5f59076yAPSuAVAw2E
9nqMv68CRqpyibAIYA/zDZ36zdNAnNgSE7tXcJjhV8taf6QwTYrEwDRJHND9LPtR7L1Nu9bfkv2a
gCum+LH5Rul1q8mIrFKPhKLCW4fVg8rsaLze05D/AJ4SikciDeED08vSkUQ+nZiYFqce5vXWmSZ4
z83Uw8RSPAO65FjtoVIws7ZN71Cgzz7sYxZc1TfRkXLO6KfTeHqWRu8qLXu85WNb+n/34tNEa1MK
xtJ5hBZoHpnlp5oQvtnCXW3D87SNaAgdAN3JI7otl/bOlvakfFCEofag/izKBfdstmNtTzljR5rZ
h4lnsDjD3q4SnfFTOtet4/nkz1bM/RjPFoHY4zl8fK/RSZdOWPJUumHwtmAd11sG8kL9NFmEmLja
G9Q8IcUkLBaRrzjBMlBr5rgqZmCIEnOnntTWR32G5ZePdGoCwthnQ50DZkr+zuH+OT21JPrSpMX8
UNdJYmdANaM9+UrQYkJxmRYA7bjhzV0Kc2ZkmkN2iZgq7e6MEsndE0jcwFb9qUDJ3nQyBMHe6mYZ
0vwmxgX9FJ33UIMN4UYsQwdBnJsGJmw/5AbEVHs2xtGCaCAh2x6XPb4pG3GsACd+Iod/EolSNx+x
k5+MaXzbgY02aNO9+lZAEat6mKTY3FYkdYr0Fs7xPHnRVB3awYxFiPpJUdKtlg2E0Af89tQLHobf
RWorhAW63vtvEGkTqlI55Cqp7lL1KFeLW1EbBQJnLU3ZR4p7VahdqY7Y6ScYfmN9HIhhUPGBwfsj
/Kuo6NzYmSjqfL0TOmfHfuyPvIS0mLxtS2Z4dqjFt9oASICABj+r+vZmSMrDXBIAt6t5lGx6+GHA
+SXSkfpsApFe8f5RbyW8m4cICygkkbC6Cqf5jd08Sk4hXK4pBG+KBgTSGcsmlLyMf7SrRcQnbt2W
p/H/XOPeHPwIbgOxfDlaSa4OTupy9nrHz7z87z5Zh2MO4GeZ9zn+xLMEPsrSqPt7FahLZe1H0PvJ
SxWwwypZMuZHr2VtzjbyPQAQr46OkjtLSG8yJA5+7wTbMtL16noUKgWtK87tUgBjrIHGurbPLt0e
4aYLA8po1z0fEDUQei2zFrt5P4xRjYEmxiyxMWaj5x30LGdR7aTcYDJ1xxLzHwHC9TTm8CcPqK7R
dKWNDYO3Bla2VHWeBZj+ZJ5OaXTQcVuc2KpRnb00RhbiibNWWY7oWmNuGIneBmACEGroonkRJXtu
XqD5yrVnvJCdsw+MCli3Ec+dXIYHvBluxuou1l//hrhMGjwylh3qRxGYE7Gb8XxKojxbndeC5QZn
aTs5JDdYyqbgwaji3LeksKhIZHdY3A+dn4V6+AcgFv5kxoKnzYEcFZ2jAXW/0wbKQrvUaCKz+pzz
dyqRL+KzbvLaI13XaA5MPvX6U0AJPzeNbKrsyRBn678y7R0uY6HDNIjt25x/9+x08YVfrHTZk2aY
HqW7bMWDCpQPn/MYlAIdRLsB0HH7vz+rDVTHBkzpikK0Wl6GKmCxECUpOE385Mx9V0OijxIReinE
iQcNc4bCMPy+d2YpYLBBRJ1G8lUZ1dtppob1Fkv8UtPQGFmM+Uq0DtqLDLDFjG/FOUK6antkx5pU
H2tO39D1dJMdOEnUj2gSVpX/zc5tUSnEbaNEyKik8GZItOgBdsIXCK/xUYDXou4S7oyK953hZN1H
4kyuwvE5R/6DULGTrRufnwTFU93BwnOY34J3QEH6dWU9O2g7QLmkUb7Vg0jWpFiiJb+hsdFn57se
mEfKxE5EgIvEMb/erAvyZdllPHDzkT+5dJiHGh3TymhHAOEmn7jjnbHppD21UZpQEMAxwyvgs5nU
8p40ImAvEFBBqQgBCio6vCB5kSpCPauGG7gI7rOhuvd5DE4Y28VpzVQSN8XOW5Ex656JjnCm7UgI
vDMTROiCFDfNCBC8GiWkFjdiQJvEySmZ/AttpelTQxeZpfIeDRtcITiHAogxuE/WdqZKgNUrpUOM
i+Bil2ntUEjoVIn0W+ZtsVAHcgd/iYeu4DeJW4Y9mAfloBF9fYlCAx9+LkjpmeTITc4RyIZYAV1W
bI6A59dVrxPtVDiDiPh4hHEjuwVDNm/81ejDjNV2or/Y7dFZ9alO/LZZEuKF27T1kAxhPfvxY+8F
b00XRYOVRsy0FQ638ni+jb7P1KpQ2v0guZ3/mSHnk9y5fkaR1p2Hh8Jc4TDTVOA6UErxFfVJBT9c
U+O3PBuMgPYiryt3KtsDzRfS711UQfrfHdJjKQ7769VLae9IglIqt1I2rbfkmGJ5vRVoHhbgBXUn
onJ9XwX9AaNBh+D6VHFUa29ORFlRWidrUawNdXIl5YExvBtA9RD948s4JDXWi1bsi5i/WMN49q6c
Vc7CvIPLwUo4/1DIQuZaUd/Y1LRm4nwGCqWgmidXnFdodwq7rjveZn5FANadKPJER5QmWlEggemv
xiEPUg1OSKsVckfP9r57HD+hoJ4v46l0hRo0QfY9i32JPdHvBD6TBHKxj0m/GrmuOXTANVng98pD
KCDC2CriLb7s5jSYVng2gl3ymbjma7xgy8gXKu9jeTwT2ybDhLRd7QXoVTteJ7dkkY7iJXYtSpKs
9OM4WoFQ6ldxiRShv+AmX8vmMaQrQPb9/lGFnAQ+vWKb1Rix3URkGWY2P1oIVH8mHISzW0WqhSry
FA03SIwQSCV8WPB3oaSK0lEHadsdsJjZGrZI4TZllKmJCD/UHz3uX1bL+YEPOrnMpunXEfLMuyfi
pKDcuovZ2eNIScC1VyQOFe1bgtB+6JiHDJEPU3JsVW9KoTBCXgOhycGykTnNW1C3xAaTQqC+xb9N
w24zTlQmUPpoMy2ujZ/F6rktxi5DWSznS1lbeoD9FDDCtG72XZC+lOw/3j+A4uxrio4ObV56noR9
Z/5jKvRIZvTo1bwHvBDAV+re7FMO//U3R/+TTZctpL3gCuOnrEQmosyEhYnEKdEixkB2VgSP2ckn
E6eINmVDqmT4b4710wzCka9sHTg6wGMd6x9LLf6brem/I6DrNKFsMefeHh8DiotrqNniaS/Pl3C1
zoj/z9i0S4G+RnFP/cOU8CFe9mcFN5JycJWDPmB/XB8ZPEYYo8dMN/8gGyspdH3Tdy+0cj0A0NFQ
k6PKoh7BW4c7YW6GoaKSV/FAOzbM847ixgbWX7PJoDnV86OJ22u6sdnuyowVTmECXX36XkA6Ygaf
clcpOPrTs28HrZVZQZdC064dXh/nEy+dNXgRdONz9Rdl1W74ZGg/6FuY0NMByqO9ddh5wxBQqMKF
i6cNkQkaMmq2h5OHVbnjTVzSmTunDLsL8egXisryd1PoYQPOP+8/r6o6b9h0C2hD0GatWQiVh/Kb
0aDWLibbq5S2GeQFHsByxf1A5XP1Ek+qTzpHoXG1AH1+p5/CITJwgEosdjrAKsc1L5uQBvPSDCjP
JwhjY8eqcYC+mVfptnSM+75hv7FYpiKAyMahBCa4glExl71zfCRolkwxR8egOZRdQXLxbYU18laf
ldlEErpwCYwBntQUyR+qrawBEGkcVija38yH5Gn4dpUM2YuZzb1H/Q2ADWJgdwt3pp42GE1DcMSW
CE6HPHcQEJnNA2kx3NMbheki695NodvANU9Gy+5w9NUuWcN5NAjhGsKUsy69rks9RJgTh9f1Vxss
V5o1XTro6eFN3tXOBKJVETs5+PznHkHjLQ/pnstU0dtJLtzZVfKVg/74u8ZxLFulC4vblmmUyFAG
d33X9qTZDMJ11qY4JE+7oNKnajxhQ+aIxUuvELzUvpGiTAvOR9DIVLXmpp5B8w2iJAc3HMZ+Ispz
ov/VurHixyUTrh/8J0Exc0O1XsLk/Jwvqyp25UA+5RYTHYaJMJlZFBb5r9L3au8BClWryfnwldp+
p8PLWmldFH/0EPPCob3BWjGipumYsJQOjKBkhfc9eu+7yC+QOgC6eQkco1GrHq0a4EM5zTCs/sb4
TD3HCUlka55uxPKe3w7yEDiExxP+oCyKFx2rJcQGrE0dEZpBm0bj6Btu37FmPl3G9fSZ0qKkgU9c
CVE/8As2goTCCattqjug+ZZciAQoGz59YGPxUsuOFD8IRhbU8FDeKBKjnj3CV+tgUwjLrwFYKyaP
45CprpZ6xxn4GOjw+2OS9JL3K8lscEbtRaGyXxL+OZtWNLPn4b3m1d3xAlrehOOqxwG7VwpR0qd0
nfuO3JmnNLlFFPbWCaa3eyqy5HVVK/VKmnIs8t7/7s5gnzWJaI/DVRXvgJARqUzqBbPZFm8zZkfr
uKI7u0558NiNGz9/m8Uf6P86Yw+loPHZM/Y+HIQEVMX20aJ5ucREsif7ET074S/+K2BWb5GkCHft
pMSvGNJEXnncGINGwtBA5NNLMZbjurqie5Y/tfKNNng8IpZJrt0DwSuxdtpdMUo7HPIZAPQfPbfS
nCmJaJFxMhJgDExFsae6ikGgxo/dYaqTUIc+Q6z9hlZEN1u4Qs7ZcRYRsdOX8hjtA0ue2fuuDEwo
JgyFl9CfzJENaonC2aoqRfJrWMVnQo+K8E5dGdCTzK5vHOCTFuO2yev5nuF6bX9Bw3HZT9BUlc93
HTp8vLHj0IpD3lITwQQd/2UbcLIeKPLOhLBcDYZqtp3TGbspRMoNJWEShGFPdAG2x5zCmXjEpNu1
c+LE/we8A9I/kxplrNCuqapUHJ+uGMSIFL1a9GFSKvvhTCPpwnZ8hq/tvKj1d9UYMxB3kEO2v4zu
s/u1ugvct/r89JWq4NCN/1TrNAczdU2Jk+X3uaokypVs6C/C58daZMxejXdSMMfCPq9bwgh3o8na
sqgCdzdUclNYFZV81y2QZSN2tWbOcnCiim+wfuuZMnCo1D9HMxs4hvs17zYlLqvFLEj3GzZIMDlx
wpk7PSAtlXLt87wK7+36Gr864RMpuuPbkWiyD9/JTj45bxrH3fKil0yVCcYV9swayaMtZofoJ4Bd
1gYSrC5ttnxIE/3wWnRBYCp1wnq6ZtfkFHobRZUXVWB4wP2Oo+5VbiBmAYG7vnIzlgSPaNm8lC6+
+b9gMe0K2/JJHMrpHZzhzaZ1c+8hAjvOFPNbcG4uyNiUKa1ALWPghJc4phkpBB7tUYgtE80fkF6Q
RuDHaaENZGG5CCqNVmSH59754z0DJEiKzYnnDWNlErw44maWcdCHoPhWrE3rsYbvY3S2+88gptrQ
Vdy966rEG6deQ41Dwq+fCkx6vsb6SweS4R7iQvraJ2SLUtm6NiNFWdIKAaxk3Fi5joy6njY4w6d9
4EqGQEsdAd0rCkUpQwQb/QK+cqN704jMZBm8qh6vyrpyk6DpDsqE5NJK7leBv6Yy/p/oWS3/l2v5
74zT4TEGzZdxu02rtX/chxPsxMt6bQX9YLsPNILO1s2j34J9qkjRyRlxoHpYhDWm6o+5MO5TTLHx
rtodEabORuu4x+B533SJ86XnQ4ewRowuHlEm5IqtrH5fMYf92ClXgGIWOpc4uc6Z6qi8Wm/9Ap5U
hLiEZ6l8Xk0QzYW3GJB8ibJEuryCQu0CWl/SKt98YU5+KiUYh3Ex1DP/Oco9ph/+fIlYq+vIKRjU
TKKkgSqGpg6bm5VjaNuttx4LZUnhVeslkvbxYcNXbya/R4QqErig6rOT2oIRgJDv+DbmJ6w0NkiF
lG/H2c640BqtLCMvs3H6GyJdXkDIid73wRJTdONBhxaaa3tplnFtD128GJXLzOjm0+Kv9EzDqjUw
bjcdzvXBhj8EYcduQPaBC1fC0Jujb218h3jL/VrNXQNldzXNMghE2H7Fu/FQNGCv4SM/FlyBMUxE
sUbfz1oECmy38oqjhaRpYdR1LCsuZs/UVzQOycTviG2g/5SaNpwQeCzDllPbMjgoQfP93He/hZWe
0XRQV+jCRwatKnntB4pVx6kPj07dOJotQWCltU0//jqUPQNV/yUjhj55CqKI68TVAb7TSDEWdW1S
LJYe2AyGllctO1q6yt8f4Wz9ONevb8GaijEkcWBtaD0W5dP51lqyOCzmA6RBiOK7n4s0myNsURuh
0yDX8e6pXJe9RXLKloqtOlTpwGeLMHnD8+/LWojrKkSv7yJVKly/ZMf/Vjt1uhiUws+IahoF/deb
X72065zM2GHzQ+8zoa57SHIdBMwneQmBwsH3WeMyENcmC9nvu32frAMx3cH/+yvYniHQf7vembEl
D6X6/hGC8avMBLDJdn73SP8m1Z/Upd91NMAfPnRCxwcLVPW5SQ/Hv4dAT25qTsDSnaHdcKP3Uiq3
Ciy7YNBLTfu28Ev+X42Ejcmkh5jaR03hyt5LiPIZq9IeEm9B+ET0zchtKVeXlxpnVIEkRlv9GuXj
xETrKk+UwM2UA12MTcsL24xFYl+vTq0tTYskUvXRI7Y5DGLOhJ2OmpBSJqsNKNVm/i84iTgmaso8
pP+CLI0MQzeUpaLQSOc9noJF+tkhwiVSv8KaGk85lF3R3XGZfDgLoYKytfrLsIoDSaD14aYSdiNC
1+x4WGYqY6oAcNLW2RqTvVttsW+5cpJo3BkHib2Un+b8U5rgeXE7Tg3FBs9+zmX5K4mXCWu1uGAT
u2OX0o7jyOhIYZURt2+sGHucsoE6PnjXtW8lMNFCw+ZyilXLQ5aUq2crkXvzh5eciIFMQ5Oom1hZ
eVdfLfCe/ysg7NIvvwkKK0dS0Ss2bYeznbdAqDhVTWXnOohTEWFH1eQg2hG8yupTnjiKbEj331vo
DYUbAzemAevLDYONHf1lDrkmBvvMojR+UVVblxRh4r8XGWzW2QUDwR/Hj6NDst7yLBzHYhHaX02d
U0U//K8fOm6fAr2fUtqno3hHvspqBxJ8Sfmc2p7md9DnwVOQj+WoF3QS//1rS+knaHx8MQIDQrOO
RB7Tp+5FJmVoLsgQwwqbJWLeqVTgCC7K8IYvDL0gmudqh6zSWBN21CqkzDcyU0zLKOFBci8lltpM
50EbjIbCFUlTOseSxotLGkQ94VwyY3EdT+mlPMmdzO/E5/CdhxJ1VEkkloa0WZJOzWNht5QRltf1
7RGPk6g6tF9XCOtYVI2J5REylu6VUO8P1tccB9E+xiZmknqdXICrS1PjEcXqjogcD9Ff0iUi1CGx
TqStfSE7wQV5ItfiCbD8JVdAQVrnq0z7PK0nzlSLAWwjQ2tgo11tI4cLetUSv5LH4V0T6glNd4Tw
nn2vp0yKqztsDWl07k4Q6GUPgfYJDXIb+ozCdnDmEILqaOlGEDY7Au9wSRbJOIXglwJHFgnkPsBU
AbrMthwFDhkbfjefFpCVMOSD3rqVfZgdxgLXJ0a2nVY7+jn+xNClTyRGey3Q9PkAnDFLkI/tAca1
LSGQ+7K/gbaj5wJt/3DegcP0YWAQsi1d6D/JoC41l2OhnNcrbKh0lBqE9g85AhKguFgtnOsgOhs7
z+mGgNfBx0/Bn9pTFKAbAVDkI0KYzoerwgYLntQEbaAyofA76CtpNefOAIMpCqNTkIiPDt8zDsFe
RwJs+o1V8T1VWrKmrlgglP90+Yu3q00uhgiCz6OETH0SwIdpFO4eZXrLhjpcqIMyeAGlpXX3M32c
5zeA2uczq8Dbbql5ObfSh1k3J1pSgWolUjU8Mag5gQqJxwlEFIBEkhnk8HRhCUALjW9uGZ1XScns
xq7b8kQakTRYTJk/7qRmjHSDFnkG0nbAqmOscN+QfxeW5Mwfu6bmHz/dvl/icyO4GXNboLesIDTE
o0+/RfrQWvr+cOjCcR+Ww+g3sJPFNGDBzutLychgtNYFroW2KfvHlD+Y8oT4KAkW5Or2Ehc/bIXd
QfsnOl5IIPYaTYq+VK7/4WjOn1GwpgoXTZpITHQkuGTSYjQXZuDQNOdXRz2ORkeLe7H5pa/LkQZn
6TmTXT2MEhZHld/2xtu7N2pJPvbqVy35pl4mZnAiJUvr29uT1bayacWIbcSLTiHaihrJyolXrznC
oZnbZwafuJ+oNNb+35KYEOB5gP+s1/o69uf+MQEuK/fC+Vs9jPQS1ttkuEg8/8eTrlno+9zxd9M0
CjRBSjD/yTBF6m8gJvSBLXsaMwqL1C1xVQmRmJAmudLww9zWur1Anwz3OllN0sh7+NbaHx3FX8SI
pHp/4h9inQIissuc7ptLwdZN+MgTKZA3lkz+8jAJSpIX6+yuwSqXjCNHtoo0cjwv0KYH4khMTyQf
h0SJb5wgHGJT/djMQqVSZtaCyJvYOppqfaaSxh5xqDvmOZARfLv3obWG60F+Utc/EG3tk9F9mYBz
2+uIsgwl1qOpufkw1E7qr7qcGhzmkVpz1cGXIZwoauEg1jQxTewWFoIkrhev2nmpC6zy/zmDWuLM
bgKagNDDTgfd/yUfa9ZbTUqyvW6I+GF2APLT3DGxuap/FSQLr0+IgDCnC23k+RfMUGL0GTrpQF2K
8u1Pctk/cEoBssuFr3bEhHC1vYQ6PTJKXpMmqCVucoM3AEbN8tJUqfBmcDxdd4U3zA9E+bBSOwed
O4h4mzu5xuuKD8ysyVZsuNoa+snbcPxba1oaRN7ZvHC63FXBN8OoKNlL4KqeeGWZQZfRG1gGOBtT
oWKGgHPspUgazRuXKUILnz3HxifvEEn7CqvGcNqX5AXVXEu2ykxhq9i5h6/kCmz++tp1U0QmMR9o
CMA8DBB/3SDAjlC7lbCCMQJE1teXQsq7WQxwpXKztiCGvRg63maK1xNJvfSQgIfjt7oOmbYtb7up
03IYYHMFoTdU4Xy9N15/Dg1BdfdzuWJ5BmrSu3wZCOgQ6tKMd0f9Gv8gcIUGWsljLY+LxiSyR/p2
ILDJybnOeaexp/YoIxbOheyM0xg0AvFc3S5MvUNGRlCe7m6SJkRxSr/1X/gBe/Lra7+d2PD1u6tQ
A0gUvZbolNRBcNr/34/aOS5R1dne48uXWnmwCt0rhP/JaBjZQgkr4GU/B1FcQccyhvmStmEn5aSh
yie7qHYNxulQ19x4Cr5GT68t0fhqHuu4SzNc1ujFslG8CjiTBV4h29uHlxCMHejTGwQMtWLST22k
dG3MfPE7X8rYssA9AbPjqfvM5H2zX9jklm4xBivDWIQxHXWBZNVMpXbwp2IE2iknh6dDKMqEWUvp
k80uz9tDoPp8TZrVBxREhlTKVP01LRHBH+VrSuKw2DG50vuV5Xpao9gm9w3n1xL0leuaVG07sll4
aGXKZ9frnJ5RcfLYORiWy8tTYIXCrZ/zYZV2dyQvAuaZCdhL0Nf99LJebgx9xnTkV9IUrHX/WCke
/T7bGtcI6G3PC9CWnhoodcwIw51+KYRIXdfmw3s0kyl6hSnTYMWmQzD86uG/r5hCb7owa0K0Kx9U
YKeGkT5SqOPv2seHC54V8uBZ8zyzz6uUQALrAgDk7tsUaUHuKJiMDyL24wO0xV0rU2MTIZTzlHLn
w1Z+ELUE0XjP5JGhIDhFykG0koXU7OiovHk2Fvk3eAuy3pbTceE/Io6UMDHcgpytrb7fBH5KNJNM
Bk0ThiJJNi6dVd1zVYsrinL6RZjhH2dWl3bYxxOLpQi5yHC2d2PE7BCUJEoQjp2yI6G+QJNHIaxB
DYncNq8keicvzhIvIXsz8BKoRwbFsm4hGve6DsdKmkl9Z2ndXPkHkozgRQuA936GFDPHpkxLwrkg
8caUavG2m+RxgkYoPpnelwGnk6ZwJNSYxYepiWwIf+czkwizbYJM5Hyzueq0JnW7CqpCHGCrIpBp
2IhxGs+7jDoXqAvYsvP5nKKnxq2WkPPMCPDH723Vh1PHGgFQ8RVqpSlaP2QC7wxancePtOA8tDtf
yPO3oPe/H4Iio10o85VHBQg8N1BfNrf9rGyCRg9M93DEgZPW8LAW+UP3fBx4UwcLK9d4DvgopnwV
t0qY2MIjgUYD6B2VBK5b+NpN+/VuUwdtVfJJUDsMZKkPkCQTVzxRwT9xDBLLGZ5gXY1T0yF/PIpE
DAWtuRMpml+hnZqZDlkWjb8iEPRQrrxURrH3n9EpqJB/fTcTz3A5Z/UDc1ognR3Ny6zb/YDg/KTi
/+zmGzB45uNuZlotzcYFHmUbFCRcHPqAR/vvopWosYReTn9ERxlb52dp8tz7lXvCeEtAIRy8xrKF
gn5KMwSEkGbWX4Eqpn1OQPoxptOrlx9Omkm5W9AyvAUcwUIyAwq72H+fiIP4gcmyFLd9AOeJs/of
+ISTsbsWZXQQKZUSZZnpoEHG/hzFePqm388YUDNaaztQdEA5LVU9oiI6aM7CCTYdXlTN6RuqNxpg
2J6Rx44cUmSAEJvs1a0TC2iXDSMLrsqUAsQ7Owq2d2+MgO4H7xoVbfamghKd228KHX52XxQy3C2K
KieBTuF1feeeMO3g12XhCU7htTj0kH+8ZIZq+DHgBDtvvWDMzVQDsAX5BdBkFE9MpStjbIDkfKdi
bh1hF+bSuhhqD3lYSmHSz/Vgc2xDhkM0MDFkCFuiH8cf9fEkhxpHEqR1XMkrlAKSBzgJgcFbx4en
7NnVO7SGT+s1HZ2uxjsvbRNRNpKLO3/RUGMI6sF1spqcqq7o3JfJ7TtHQuQdKdbgdKsjlGLU58qY
zHY/tW1n90kz2Tdg2bVhOsUyDhid8hJrpqvMSv/fEMv0+FVKnKjzEx9C3CWvgz54/GHm+IfGkUnx
APJMQj3YDVerP5pBl6njR769d1CCfBrFCYru7YkIxnQtofx49ZIauxM8ZJ6oIeL11oPvAiDuUjFb
DTtprE4D3GEUDEyWsjyFN+dsq3stCJbb6GaR/x7k0QlLePrIs1yaYf/DRAeAFJPi9inqzcNeLRWX
HUnXRhmA+eWbEYmWL6BMvFgUVB+Wk8D4jxl3/z/oxR/GICPRv6HzJVxMYEGBvnrkGJ3HKk9S5LvF
eXkrFQ1TcVqONlVOGUXlUpYIsBH5DFs4Hv2VDbh23D3b4Eze0mk6DL8S8UO4EPwJZPnJAHBqa6gU
rAy5fQHnM4wpR9grPON69fIi+0Y9dlhU2D71G5HD7uCxy7RJFlqcKsB5cml6uCeroaSu7qxxFzVN
35HJMo2TIcaSwI3ADLXIJGnvHKW02YNxhG+p2Hx0inKKLtGmPOtezt1vyW0oR9onkqXEslz9mvPR
O3GZ8TZav2CDZeyvgcUQBP+RI6RjzUZ/03Z1a0RuSXc8IB5FE2axVJKlYO79CD0dh1cQ/shaASty
fqzBkujAR3iHT9FanbthSgcL+FrNnwKwZn92rJ0bcNXduz49sPOpcX2qLEwXtFIWlttnNE2OSWgQ
9b5f3WZph3rxYNenA4zIjrMNp5meAAVYbavuKdYrySaVSIOsHUVrEi1gbLTncDVLyMoXcPjkk7IZ
biDsmn4ZzeLYU7Ly2KcYRBX13Hm8u/F5GwgmiWeV/1RTYycTLrnbcCujKH7XbqZPIn/xO3sJKGSM
4+Ovc6ZB3bmVOyDF8KPPzCWVgbDxNO73nHkglZLNoTt5N/NN+e9G7SxXUOX4UoenRvoqPZevezak
rgHJM5N/p89O1Ser2Thzi8OojXWDShUrMQXWDaIedONcYFa9jCgTbYoFxhQhskSf6v6dNSKZfnJ6
0HnF6niiFhQIUnulVjY72iSka0hfI6rFyhAhecYoKjrqtQKLWph7fF19ElkYrT+ocqqvZMCDrm1a
4L5j0abwotTh7bm1pnHSEz2Dgk2KqmsbUbzZA95FQ2QX2Kiz+V7t675Q2WZIyMgmatSrEI8nDlNR
1IplXzMXcEMiXf/hYZJDIyzQOOgyVkvmvy2v0zR9uZ9qonum3zfYos5Kr5+BXlS2Tg79wBNUq2wZ
dtyRVlmwTgtoQwQxHFtRnsDjwZ5XKvl4TE7MZiYZRrVfAo8SsL7W7gdoHa4mLCdd8B0Ln4bPylxe
GhoKus2uiOMhjwJfZtCEHE8txvBh/wA1wvhZjC/hqXlxW7GgklhTtTOQIGag0BoR6ojfE0r5CIzL
BRqSXze9+M1OwNHuNwLkW8ukd3TEiAhLZYJiu0SJRrYTeQsBHDroNoEKRaGAF23eR4ZCeybpI/kq
VTMHlZ5OoW5jk5SNNCq0TfNMoo8muKek+4EadwU/a5owTd0U7yDYhOTY+h0HaYyXhsbyIDo+bwRb
o1TbPPeRt2pbQNRhe0zFcXDpSgTUzxYJS0EzQjQQlB1saC4PE6CEqtw3yg5OkVCkkI1sWpm4u6dU
9FawVD9of+W4/DrOqcq32ovwlVBRlZ9ouF244pyyubC6fGO++oExst3u2mRoUW1QaZlLoA6kFoU1
IsPOyS1cqLEY1RA/NG82V4nRPILFoHph8750lnR9uW812y636+RIlXiXR49ibuezJ1gShQPXlnTh
tECWlEMRyfYaOuULtXx6pKQke8zX1BuhQ/6lSszWgrxJ/bt26y1Uan7TxY7ph4Py/9hNAEQ1VPO5
2kDPNMlkyoZuaTIeFPZL69HXSuoi3Ihw6qsJZaUvB3Hq2Jel6gqvO93RKkHUraV924742GBLXVV8
yxN6Gv2Z/ZLJR6c8j+LH3SXHqUE1E6YJHTe2RldhnsQjpW4L35HdDAqejlqota/Ey8d6CQfJKO2k
oYsb8553mnpvlF7QZqhyD8nXfvgyCYVf/fIBAuFVdkMpuqQG+CeIJz8W9hB9D5Dg9l8hIlf7bQYO
hUmaDHWJ+usuF7OD0Bn1Nm2CaDfXga/biIq/Ohxqwp7Hklxdfx0ihqFnQ8hYWydLIE/nz3vnjd56
hpCGH8VGFcDb070+DdH3Xji4JUol7qElyPjuEbfh48BlCE3OLQb9iBLzQ1PXk3Gd5xRw8lstgcrf
0m7slicuXNvmg4t9szKtL6uDU2J5NtWzjs+tkN45fgZsT1AEZyDhwSDXoMRl5xS/FsF+tdZw2B1Q
hyDqzwhjJ9gxABKr/nb7MThb+eQoZCdZdGBxY67O8rBNtvpPJKEZJkojFfq65NAGVLONmcFNpMwq
3+NJ6NJPMw8a+H/tJGqRqdUmtmJyr5i/0nGxhF8X5EHCIkN/B6Bu6N9PKcmoud/3b/F1bhHYka68
Hym/tZs798KhupAb7vht78fqeBFy6CT6HZ0ZyIy1owZlsBRTICi5SXHs+3zS5x+Tjk17LPm5VfUb
g355chXuyzbofVMfN9WdxlUwYX1K2y75RYOSVEj4QZVLRZx7VqvvFzNDOS+FRA+VTPYyr7NXHejg
SS5WuWWU8QeARizTPnebj6cylOxnXAtp4wy7/m1yio4QF++mVN4UqevbVCixleIfW5AdoZ66oa3T
sW7ZOJeLo+Gx+fyAgTnjXEPJrQqR0NCDKwGRazu9S2yoLQX8YFwkZRx6STdQTzcBLiEumNj5j56E
Af7oZpiy5Y5+u50t9CQ3R3MMPEoCkJGZW3weF2ANOy6GhZsBCUv8ZQNyIeEgE6mASXthQidCbn4o
6odBiwenGkEzRPowQ3EbHYtyCfGlsD9jqyeeoIvHVcsHUb7PPq+23q0zg1s9P+AnUmmJpIah3FCv
B58/bdCkeGd5lLrAxJEnxCZgyvUxJ48wo7cFTGbNu8YZFMSpme205g9995jpcMht3IqZk+jj6MOg
f4y/AOeaD7MggQWn5KbTcfQavPS7mDwRVjyFADvlgIQcDJqXBYUw0Q+tcMga6Pb0vEA3dzTHX7Lr
8inIJOGqxFmFs+YZajVMQ6jWsPorCspxUHHavramjHKz3jlWS2PNRT87pgQRkJGO30oqg8L/GAgT
Nnp9K54Vq+WAWHTyn09Yogd5IyDiKRZvA0qzqg5hrLxBurIZKRtGESLkTMYd+pLNJik3HYbcaZqV
au3VdZbIauavbep9ZCctXqiTJCmQpWE9NMJjHUf0CCgX240DcpSU3baexSgLDWY4ix59OkEajwNH
O4whPqn6tThGc6JQPV6WwYFlo/c5L2oJKhsHEv9H9TROi1hZpNAzOi7sIzy8JnU1lEvtcaLT2sZQ
Bp0laAGpMWvrvb/v1mkPc/pdmLwHi1TLd9rFb22nzZ9Xj0riY9bW34AjOFehhGkruAbQ3VsPV2fA
dIgUmFGmM+C50cQnmfOKfEgscXWohjJA1yBfh21kluQJrG7SAjDwgMqpkJB+5RX8Vrd5vZTM3wve
7KO4rLsr+QBHBq2JM/NKC3EnJpFeUatDlblC20KFxwcoOEQ2pz31R7QNhm4l7KY0+ygFXffRor1K
bYQYfQ3CBNuzWL/BlMtzJKUGfU97gPUKo8i7FYpXcf3mjVoEfbvmcIYFxlKlMRido4Lg8MZ5jrei
QPxwm38nPh+XrqQKZA4oogiGXcUdLdG6dR9ECjG348cPUrSypHI/AEPMkT4Az51elJ6bTVGDUXlb
qf5w7u4IVlM9VLDzcoZcx+ci2DOoISOTotK3pKTMQnZatLr09QIwXXefPgkcfl75umiDoOqden0m
GBLPjTPnevj6hweJqEtlwYGlA93062VKsedXGYaIx9UC7Pfn7HH/1YjmeKJW7E7ErfV2ZDJG1FK7
3sw75/kF/7F5Wgf7xgvez2B/dDJABQvrLhefSWo068EVLKLc86dZlFKWZL7wPd0lODJMSU9TVwo9
exaIajdUm772oNdqsSJDZ8TjPBelClIxRc0mYdEvV60x4fPADlYkAcW9zUJSlOob60dfvM+vQrFI
92CWCCZBuOUIeSn3BWR//0MDxHfWgvW3B+P4eNhsBwfOI6fmEc763XpH70xZqgxcwC8KiRWzAx7e
teJgob6uEEQ3rqmcA249vwr99DwwKzAa0LvyhbvwlSICiFimoxIFjwm1b8UXqaNCB/pSPTvLt1FP
KsTfclT2f4xxHb+rRKmC/gJ9Gg8IVhleeu4lgkzanlKnvTO3HWS174V/RQoCLqhCCGJeDgxBsM2a
2ej7Ks9TYqYir/dnuuYsCQnTAXa88g1J3abwODTXmU7EoTho3WNU9SOVH6YCx+2tASCsH4+p8/jQ
n7BCFGrWjWZCTOe47oUzun0G2qj2BD4/vi970gxgX7L1xyRX3LiuQ8SXSsTNXhI5KUojacF7HZ7A
BDsAvaAFskonWJmrrcQvHaoJFNfUiH7Dl8yuwxrWi+R5mnhfUY8fA6Kowq6c7u2jpjanNpUd01UY
AzzFsCzhOZc4vlGQ7QxQUzsA0LFw8SeXKGwwmSSS9KG3/iTl8dbRo0v2ns5LhQ2n4ghgUqdl7Vte
TUe77XvgHthTXt95lKgpfE3C2M9AMKeSkFQq17muweClj0aH2QEmYy0D900lTQjHm64RjQq5CVM8
QL42Lxht8kXXFGh3nODn/qy7R0PiAk1qb2+1MCHYy26qpFazZ1q9sK0jWeAtvneGtig0LtiyIlpo
QFvOLEKFlIta8E2crBF0cw32raeupSBOUsl6mu5ae+91ve6bpEiD7iQKfkVkYbhp+NAHhja96aQ6
CyZr7BPWl0oThQmrWclTrZpaa8wQbbZplPVy2mpkw8e2hZvBJtUvyIrZ/USVpjm8rop99UliH6he
iwZN4JUiDY175Yn9g3jjPtyKXDuJtZslID2Aeio3IPedGGCgfQeml4BFLswuL7hK/xTWTGpCHHoy
9+1aQft9YFJqSx8uTilTcmXzaey62dOSggwJZhDBHvtRbxftA58TxkVPC04cBhs7HdXl+QQvrgnG
CDGDUHeDH+txxO+YdC46LPu14CUkXnaNKyXVw1CGAPDQUSYD87mUgp/6EIFiLGykowzeBli0OiJy
ZwSIU88a+Xs+tYeEn/pWPaU3qOkU2KEj3UAuvtSz/6KsKyfpsXTcqsVALV48tU2INAFTaqTpnYP7
LA7YcjVmuoNhGYYE444TUY90RcS4aJe8BRwuBK6QOvc6aaJeXPcBop4XWwFyZcF0dK1CQVQk84G+
Z0Kz7wEhDp1RXeOno3mbw5d0CJQvd95KHtfKMNK3NjWSQgalhAs4QQ7MRgf5hG6sEXBTAMOILQWN
Io/pFeT5WlKCcl9UQWm5ZFY72q/FCAjqjCHVduDlVBHDMLxW06dEvXTsi0JSIRwr/CKMvNrnv/ug
nT8AdEkILESjBm1jy3Fqi4i9wP/3/Y8RZTY0NfE+UQQGr8BpgoZW3ohbGDGjfzIhbAjw6B87xKQz
bT1aSSDGvdzMjFSmTsvkp14ROiGrcoxpFD2DQHW5Dz2lSUzBoqwmrhD2B4W++Mj2CKrZen4z5EbQ
jVPbsor2BC++IEO3uIYqVkROZLKh0mHp93gZ5lZL1DFPjp9o5AEOwi1FkF/wKy/tBZRflQEOOoQw
nZQuF6Xir2WdlVbQa1LFquTOnyk3+mwnI60oyf9vr9U+taTJPJqUkC7Sn/vZXh4c9ytYAoAl+pNN
LXjLQS5yxTZmeWiBMiwMJJSgtwqyiacjDACWvXsgQJg8ZY5MrnuQZ301CM57QISI3qa8TMOfsF6S
MKArJzIZAoQBeW051Foo6MjPcnmvGKmM9c4t+tmOEOfbQfwwxylA+2D41LsObTXzT4wrnLw6snHf
Eu/8mf9GYqLUwfyvxc20C7T+DMzi6dFghExe78vppzalU2x3W1ukUiJ2ws4qx1ETVvt8nnE0kwvG
gGSmH68NVBrfySYcFByNMh/XGhRlZjBFmfP0tlgGTYlnUkWQWuUfnR0uSDNrletTQVwCbcCc6x7f
dC4r4nDWAFbCVKHBNZYpKtXsAfHL/7atMT6ZlWJx9i5KI5GSZd8Smy0vw5+XXxB0UPB6Fv2k2QGs
rLh2QJmC/eVZFiPKomknQN6v5bxpxG4zhSqmsKmGhDSCxWbHomtWe3c7zTrVn+okq04f4DHflQVa
/NMGyeWBeJJhVajiUlCnrzJydsh7CjumQ7tUL2mcVe2N6MyydFyij3DPu1d3Y5N65Tcnyy4DNku4
BmH2VhSgJ4CSHdL0smrpM4rOr/D2ldv7Ms3aM1o/g3A3c/uRU6iC4z0BYdQpuGY/4rnyK/ulwhPr
xlrVseuobiV3U6h/r0vYWrOLg/foLpcntTVLNDHbCuGnbhBY1GE5A3w2s47mD2DEFTsUap/pyc9R
nNkuVTBkOmgT9x9oleqOiGvrmTsFWAUMznR7okwEY2WBxJF5xcnUlqtGd+y9qeDxt1uN1P6x1aBD
G0hTGzhRIHD2EO1/VT3X1GrFK/OqbV2a9uXrLu8c1flJg5TJT3nsEA2OXsrurBaQsOetU4PvjCTi
cC7ej90BJH/TaQ2xKrx8j5VP4vAGhLqQeYMIMQ+zTQ/VCGtEo+qWe+Q3Myw+z7PqseTzhH2TY6Rm
GthlQQA1EW9BSmcliBrJCRH9imAmtOT1YSJxtcAI0MtN7AKgihNaM34rHOhP1XDemrp7/0+rqDf2
kAfiW3GNXfWICq2xgdyjO4z3e9xWmrBH5DU/CVjAr+99fh+VHsOhJscrlKXaMht5aDs41y/se3f4
fcRryVicSbqqhc1MtM9NF96RUeYDFxq3rkU7Zlf7HF/9MU0qSVJNB991atmjsGC0N7n/MW6CC9fj
nnyKsZTMXdH2o1ToKTBedfigQPoH17i1B3S0/9Yjw1x+vVspCJ887fdQ5TZ0DODPqRV7ksNmNm8w
QVhL6mhFLpdUVNmAFbprxoJLqE3dPfMTal6z7D8TCCFwQk3N6//2Gqivbcwb1IFhI8v3M5ujMHlr
PBPGbi8zsmo/B5hnambdGF6nqvkhHpjer9LBojtVSkirZrPuFhRdapbI+Vn7Yt1QvR3mwy1boQtS
O40uhs2WCQ5LP7j1+h0BS/0HutEp5NRQLsaDgcHhv42kyWTiJFje0Y8UndQVFHRI3+NKsX7HCzWw
7QTbjH5iCS8aUt0MsBjnKOuavxeOzv9dUFt15P7hAqcPyqLo2yz08DWceYimdGL3iQIq85oPfxni
Q3/iH9h66Sipm6QiRndwA0E9GD6GmRV25LkDlYbN1k4d6P8QSCedVNod95LlUr5KOYndg0ESLee0
GyCo651HNWbktv4IVmkhftwxS3lO0HtPUdhfu8N1bYT+HEhVBEO+R2ysr0JQcHkO4cKQMl3FhCUs
GrQfjRVWL+vFK8ntlGtjUXW2UM9ikS0WVulEiMgnRMAD5RpaV+6+ffYDFdy2MXZwLQrKXRyWRTPw
/v+V8FfXeT2M0pK9uENfq7X8CI017p2/E1bbYKNnbPM+aDtvmipd4woRtU654/KrZSRAUc9k/NfD
tsIiqtAFYf9p/aIicFjtf+1IkL6gNLC17KOg+jy2TpTiiCDhKzY57gEpQelUS0NXsbhbsJhLUNI+
qYgEfD+E48AXymqmdeHpyWNIWDIVJ8uykHNgIvOmCp/ExQD93fon6bIRHXbMtWFiGHNbJVqRtMoR
szZI/cgwOOSeDDaaD31o62HxzLU/iwjsqdHn10GXkPg+4U03qJTATEDNmw5rUhjCRhjSH+NbQZCc
xF9dP0qEmYD+/nBWWouuRcxwG9JqYrwJXfdWwcxkykxRS1eurucCEY47/T3BEduNsYbv7tB13MA7
cCxXoJJeJosj+rBzZVuCISpuXQT7kIC/0IVN+KMjk8S98qyob/vV1tnAwg5uZfYAvvARLx40ES4P
MYMbA7LjaEXVUn9a44geSC3i20QOY1ul93zEaBTxWkWWBlHRbaZ+xYK0tvRzHrf0JR74DjrlMDBR
76NU64i7LrT/lK2dzViSn7thky9avsYUbxfXkr047YnwoCsdpgtb02mtpP97IBPBmtaXHrcgkDme
YvjdKPdQ609aD49U1qy2UZ7AYdHIBwFEf8mXMvDtHo9VhTzk6MXIhJiPI9Yskder0pkNWfRbvaKw
3PKjwOGvdq90oy+CCbDsFIWNCA9hEuFVEFdpJgf33mAf66Ekht/OULC8pO3ForMO4z8TS/JevAk/
vuwYkdmb+CzZQx+T1sSkB7UIsVAODePGLrn/r64WtSKaRKO9AmDchiil0oYcS/Ge0kV0p16rWBbE
trx5tc4TnlxtxQhfVbj5IuX4C4+GymBh2QVxM8Je+eHXV+56RWr2iK7DCtlcMRl2TDSkiLd/RQie
uge7QvK1l+0HRBGX4bRC1Mmq7LtEmkAU7I/26UI5wQWi9gZwlx58BceDlF0X9UaNAdWofd9qEwgO
9GS2FfrgvF7WoLGxUU7JhqE6MJI4vPZQMQOYoEmu/4SVPeXT/a9BfD9sbQhIvEQNICNttdyRMYb0
oPFyG743uNx98z3XJj7b9dFdbziX3hJHD1dCNwrXdvSI1I7MS4jJ2nBzf2hvhUAjcYHbUPx+9BX3
vZneDAsooFAe0Lr6XU2KsNYiMBxX2W8QXgTmnIfdUV6c4AxqmCUkHLxxrUKaz+EC5DCAtssPxNpt
VbcBqhW5VsYzZbEkrOaN/Yd0XOQNi/FMHMOkTtes3/GtVNFw2RJwt9Ug5EU8NgNoDUdB/hdesLHJ
CUozmic9NtiFsp1nHvRVZZzYUv9vUoFEaZ/onG33EeyBFzXIF5Y7UeITsiRUUTJaVSssMj6+Fy3N
QNGkwEtQIn8PDwt2VoJPu6Pw5RzggaEcDdrj5B8bkcwyc2z+n7ole2Z/lH5zBaYapmHia+GDgiUg
C+REWrjwC0QdQ/FqOW+UZA0i7B8KMKMdxZUBTGhJmtsHUvAylZN9YHolio4SUagH68J/0amNdIh8
FVmxzlWOh6jqWdPWzZrj1Hv5KiYbkdua5tRN4NYkyVqIdWKEAYgLf7KNzv8LymwFn5h3eAumjwI2
x6Fx2Q7M1T2GngzGhwz3runBhFh+w1Lu71SAgki0B5G3dk6PDTZK05pOYk/hxSnGANpEo6opzDT3
cKk8fScFp0i+0uC+XpSosVmGelsov4dlv8RB8b/b2gHmgX7VSAVZh9tzjSn+Ucwj32K4kZb1yvIe
/Qh6A0hBKLPiGfxB5I/IrFmeguAamkObXa+cbBjfXd00Xt3wSUQqCJdLQQ0/9AVQWzkMRW+M936t
zJIkG6wgffuPNyh+nJ7c5+uqXCbI2oJDsIbDZfaFVDQO6m4/hzbeYtTTlyUlkItWvOhDezINZgZ0
OvzN5vQcfMuNj9m6+gyMlHkbPTfk/fF8pHCU762nic2d4kZk20RYmeobdkGYI5eytbkp+MsdPnVN
Fbq0aEZrkknx9pEK0YgzsHhiTFNhCPWBfSpLEthMSnVW+m1qCgL+vOPxS2vrZ6zgMN5EFxz+x6Cl
zGxpOaKpGZ4XherqIJV6P4//wLkF1D7NMSk8PQoXqJdtXGjgmMUqZkKghke165ehqJXW+j+/0kcE
b+u5c9i+jTzkbNW7CKiHkRMVJWlrcfcvwNcJtrvfhVPHNZK+t8vkVnVGWA15WZOYLLiPDR73ToKd
IOYcfh6I76t3c63rN/Ep8PwX1GyFwM6ESXFewzdj/nZlnCzXOXEa1cNChksB1cwQGfWbtwD4E61C
1uizJumkx6IN4oge3woAAXDjFq5Z3TBJHY9+PJXLlmsyI21+5IMZYI75ThcG+HqZYijwzSDtBqUB
KJWsD0ZHVinIrZBeZhyr8hIKPsHQy6lqWpRO9ASxjQiOaK1HSSgdtJL+9FxLp/Ve2K4i6pj5muKn
uSzcY9BwpVCMd8kU7R+iPu2MCnxaB656BDH6e7xcOi+GQD1rPDqaFqrZ3h6+bXHYUaExOsb6bBfi
wLIxosRJthjx7x5I7UxNWoYqaanG2HNmY9KoEgGT/e7K9F6FjcfUHle3qwln2tOUN1loz4y12Z/R
txffHof0+fDFeP2iUJ8Dn5/BnpbXH/QTLK1aNqQnR1PFb0W4seNNtF1FK+KoPshkEOSrsYGC6bG8
MWlRrBHcBfT+Mwj1krWwyyLORaDJ4KxERbTn40+EpeQFfksv8n3/kdRkCzOtX9pWXNXzW38XHGqr
1lU9S5d+cmLZD/A/+fb1Ag20JJTErGrah2/0lhUCwz02rwUE4AK2esUramPNo7rAgrs7EifApYl2
TSckOOsklps08FeX+wRxljBRu1RE1RkuaqS+jbTPcZp3q4T9CjvbdLXMciu2iBjbxwCGYi98ufPR
nEq0UXpkEDIXJaaHQ8UE1Fd4aCIR37WdgY9b+WIcicUOcyOvlLWvWkC2ojQ/6OCRyLnP8dT4o5QE
0uhepz1FTxUMQZVve7IRnblRi1AcxyHHJfY9qzOcQySo3tRKR06yTbsskyTCi4r6y1TA5LN1bWGO
4As6bOwDO4Umtpr9ugSXT3BN1pps/rMSHbJdOeks6WPCXtGZVK1bzXjmT2aD08uJSIwYNjmy1tVd
fZny1sfem+gMsaXi2UPa6XsqWvwNrnA2GBZH9rdvNKmWPvXvgz7MzATPoLKj66xpXDojc+lopQB8
wutOKFlx0Bu7BKk6RfQiqksG8Atq2TDDtORRFpwgYJQOaH6zx047lyFyJpQH/xt1O3tcqFlG3WY0
Vu9eEt6pYTuTNbuNonwtJBf9xOlY+Pltnt0r3OKXPHCUEHduQg0AuLqQiTutRlyS9GK25zmH8e6g
tE9t7vFU4ya23pjgUicSEnmXA+pGRo+8+y8Yzpfg8i4c+B+2RIWje4taMJbROFvI0AxAKOqkznLJ
d9G1kGXkBHhXC+OA6JjrogQg7QLmb4uS3VZyybWatAoPaQw1t6wFZwvBH0Zdj1H7XiuURiPbGMya
jsfjLfX0WHgd+kSlhtQYjIH2RTL5QFhWu4hR1eK50Vh8awGoU87sX5cK/gI1rZDX0DyYrbvsRBvM
gTnEtLpsY0fGtOKnQr+TVgZ62tytXv5+YQ51DQlGGQMAyH3Yntg1AFKU/2UsGPgC2kfcP9qFsIdA
ZmWRs+mHqIpwhjquORRiRaO5LY+f2FBG0P0xVavg/LaHnWFsczTd5Evrx0z+VrSqxGQKjA+J3qDz
EhojHu+yz4z/E8inpxfn/mooRrNOv4qjR0CYwOyHGuKx4SxoyTb6CM8h8/ePIBB1DbUQ9fwNPap/
YtvVY2Z6gbIq7G4dFK4i/iNufZyKjLqHp0wlAyZScUKeXFWOhABUh3PKZBHm+2AxuOoXNO6ZwB+h
PopOkI6s4Z/kpQndo3cKfF68MrFsfEkzXvb5/qF1riEWp8PrT90SAmRR/f0ISxcR+FZV3KeZ6t5Z
oV/bhsxl20VK8bserLlMNBPg1SI9LNpATJjM7OHKLAwu5jy81erf3MJP9Na6hdA6yf1kb1RzPX/F
5gongIAjfAfowaQN4K6eMlpHyd6ntBoMYk3oyOGZPSMRnp1Y6ADDvA1VYJqjEuCz/nrceqLQayNA
IRObrBv3ndIYoMfnS9CxfVFmjpjnhMMwmjS8GmlglGtvF/WqdHoZ7SEhdQVRe/+6Ul/uLw1n+76A
gwHqRvjj3rpaAiZda5O/eg2rVKeRdGTInkZbm4pkKY9nxtm2U4Uxu6dxumNx8rOchUgCzYXZ0VTQ
FeE+uspo5ZylApYuldBdM2nD+ePGbJ3bzOberpfmPruiTFbbf5Hcvm0l8Ei64+f40RFYwQ3ooUff
jxLvbr5WE+A3klU8vYhPERfzpqDcpDyQ1ImzmGT8MfjKUWhJl0/IzH62hbtAL+W8MXHwl7A5ewLg
/m5Seh2e7pJKv7iOzu9mLjLfKlEUTm4d7uhUbZHdbQosZng/AqyCX/SkFTj2XyuRJdl1x5pZ7MVa
vvpu0aAnbRXtl/dfr1vi1Ak+V4MVPAL8SnYDSWHJqoyWyOKBNJ2qgVvc20MgGvLh5InwvuBxaMNb
r0FNwpgAfwrfhVPAkL9xcfLTBwgzySy8PzyFzA+mKzZWfHvb79AimVhyLa7EbzT4kvdx67C4EMGX
42I6qCd+37ZkCHNCDgdTs3rKOB32G48fom5ao2bQ06l105MBQQ+xO2FayQ8AqAF4PmFSh0F82iTG
ihqUyrPRtp2Hku6BR0toyie7w0PTQdUu4AdKVkqCYbjCIUubcSTiSyqWNzswbsxpcVRaPXUWrYFS
awSf24i0S64zLuF/HhhYY1ywBtBijyJRlfHoSNZoqJ/JfmDtiPHY6Yi2IDEAMTPbFiUmIOTxnRKx
3ieV2cU5JJFbWahXUX6aUEO+3HVoyJghNCiFq5kY9BrD2aE074CEGzp9mVG3xKDyZIBD61gcTT5X
3Ce8nY4GUtvGqycWczLM7lsiAkQrcvgo59DGB4W3RPbxIRtP34Ib+73601enVh8Yt+/WuZnd4Kpb
1rN2j9RK6rvEr8cRapTTG5Zah/WjQVgxJrNGLoz4Qc0dLfnmn11YSzOzxyjU6/oCLjJa9qK+Wtgs
uID2J3WwHNKeDsLTXCdpWWnnS+3kUJbYYMCg+7lWt2ct03fto3qWiLPqCChEXJ0IAi7HLP/AX0f2
ssSlWQ87eGWwhRCjeEOyIJWcnLEI7CahZdPJjp9P+a3dtLEPThx0dnc+6yzpAB0AjtxXJUAkpbRI
G9djx+3zlrLSgWK5g01P7MW4LUGqyafvmEfl/nKZ4dSsYUDWg5u4L+aLclovF2w6+ytL6jc9Allt
ymT02GnLZJRaTr/qNVLkxEenURuXBhjRiZCYIKHd8ZZyOQcXPOPAnWwPnTmQTSGKAB6f18Da+3eM
Usnr49JcnSFKIlj3J/aCt6wPUg3ZmN59dpfwtw1IBTjW1CkM6kCVBdqUxdAPQ0xXlZqiIGDH5G0B
hI26/T7WzYjqEH48NJNeN5Ld08ZyZfX3wVa4ZogJ+8mzFhfWtmhAJtzF1KSFIcabAYiNPkb3L+HI
vJZmBk+ldhPTAkykuGzYpTZO9pFhefMFRaKmLppibFBHrVyceAxNw8N/By95IGZgAWBYXPAFTNLG
JbtA20XE9iOTW+aGoNYNTAnKZRPtQ8zAbMaPzV2zuYmoZKnhxYxadQscsVW7UNo/F3K/uCnUaxFj
rjEI9+iBqJN7wBlLN2U96KqOq+JDbSorK0QhSmgtzM9iEiFWzGNb7EFNU6CVYbhjB+McDuBVTBQ5
zWmPNWthDXm9RdIoRkaX0mJKxkwM6zFlXS/RQVAyrn6VB8iMYzfjbcupmvhgnz42G5vZdnuAEAeO
l0QPVCvRcF1NCNOfhel2kNY3kgiz4E7b/Lf15m75WSqp9xWxH0jPd/zjk/mgejDEttHO+h0t1v9c
i2KjUWQ1AzVvj+mZbm7F2vGCzuQMCdZNZhe0Jbgdv3O5dOjtXC5+W12a0Bj86Bn2igLjOKVnRR/P
pWRSqnrRqWSPkXagubbo3drGZRUEFDNIk5DcMJ85YrqgBeqpl3arUQgs+mHE64+LI1HUstUgi0np
tXcp1Jxo1bnxMGqztFLxuiUwLl1fuAUMGDoZoYZQ2+QKyf6ATGVfv5Z8zlKovA3YBNf4qs7aH0gz
rjNrxCvUHc3876sTUxkqzIFRcGXdJyTbG9+nMWaxYoDdKAXkXvx8oCfmX/s/1gqLUu4Qks+yaGQT
4Mkwi54A3f3ETdhFvZjaXW4NReOicWSPWyWUu17CkqBZGd+C/KDg/JBmZqLuY1Xmph9pH/Wd5qi4
DF5dHm8JFQG6phbPft3xfzZ/bTfMAcYgNp4tZ0U9HwmdLKmJ9L+glV8HEJ+ptgxN7uFWQqMCjtuV
h5Im+Rz5aiI/OuZ9FgJnDwkQ3qz1dDuBJGc7mMrc4V9bPH/FoCVC2HxuOf6oghpEfzNMAFswCoJw
qNuxTiabN/M3LHWqaoen2F8bTIJ9CYQC1jQxZHl7RMg29Xk0pcYgNZNCeSAJKIttYUwGt0u1G2A7
bX5a4P9CXseVSOIGm4xnqZKTjuQDcxJgIhwJ6yrI149dPvcb86upJkGjHqrb63WJE8RidZZbQQlq
q+b9ALheEIZIvbGcz2el3ip5lpnm/qcyAm4/qMB0NHP261NzMAq/DdNirNTjZn0zM0/OCblb0Ejw
rhQahBAjkaGO8cTOoWAt/h3HJ5BwegSXvvLckMD7C39gQiKYJLNnc6LQ1mCIuy7LfkOos5/lEpQW
Rp6WzF37b85urqRXhI2tJ8ua2erJ/AGF4caoehxzvR1peGZ9u4ceRZHZz3wnJGK93N/jAGBuYLWS
rBCXQZhXRf7hjXhkhguWNoECE0dGmWSk5v1Ef5wQGixYyfkxvADJydnzg/rzJdhJ9XZiFgTV5j0t
iCg7lMZ+wmweGaZQKpx6GDgS3akdVLE1H8U4xPfqK7DK+SELIqWfM8KfRJ6NVbG/X+BHIwWUaohF
ao9ka079zXvtw/YZUFWPXoCDGyLhXWJZsjz4FN4RDO4h3nokMs4TW6bCcBQg6VrpfkP+9sDGhVCO
L4mbAHHsdhllFmm5YecP3unuEeHfwLpdNk05pFTdsOXO21SGMlP24YGg/AOg8EROdykYHjSlXDmx
+6LZwmio9HzcrfawmUHxngegvkNqoTTcxfUoG/5kwR/Ie64MHRy49IhkPoDlvH8nrq1ACSFgg47X
T7a/7c+6AJDhV25RqV8IpVtEXLpC5Af6SDWldvefBlHyETj5SIfzGh+xnhTdDaZgIx6cAP1q33Y9
63VFZoqlkwufcn/F5N/0+0t7E3s5P1D6SSfX/rPS4W+3A4VN+cZzrlU9NIkwhpp3UMlFxf08TR7Q
q8i9ypAhmkubKr38SmpjqJw49I/BhJ6IYQcic7bBY4QiyIzOG8cjyNXe7kl03WxDymcuE95Juo0e
GhibD5O8bUlQ8p/1IVpt9H6b1HImEDvPn1pvWqsQnZDlAaI4fVi6xdRNFdZhSf1JRUH9BeoffWW/
fv7lW0D6cIqSmJEEKYWg2T9BqNi04iygB0vl2+7PH01dAD0aBiqJVBAyPkxADYMnpRjqU2vo0/Kk
OQ4nabHx7P0v9+stnMjITyth0mS2fq75OlcEA1gYCA+URAX+PayGFa+T3H4UtHHTl8GWhzbeEXOn
SFZCNYTnJjD6MlQm6vI9DsjxyLbmqIfWCUQieRGJheGk8yBrT+6KpDgFkLl79xa75BbpDPG3m6DQ
s5cnihjuBQqcAcCnDe+cxSkhvT5oD24RdXTbq1CvVmme1YZmDwYfMXRduKbRVjmFAEVV5XHupH6O
B/wXHaC6Vya5HWHMFxoIUyNf6fI9D94WqyJvjFohBcV89lM+gx0kP+0NikM2wRM/yHJVecoNvkt4
siRuwGj7M4BN8SOk2Sef8Js57WdvuL4bjJGrUJx6UKyJMZDbL92fAHUjrCe6Ao+ONmMFiiKSJEyV
/goTwhi1ZrQewFd1J7zRSurCBd4M1hAyXGT4Gr9ZpTGLPBsXEUoIEF1quZedSm+1LJ3c9ptu8obE
ZqeKyB+IVd7cvRipbq0cFqFPANYoa4dU41t3OLal4YT6GydnIxXIfrc/lqlAoT8acAOOLZ+u/hoV
PaH4WdtDumn4KesuQ75iK/f3hhoIjtH+orrWo6ADgQDwO2aMSOgIH84FdD4Ia+2Wj7Kit6Q0+tHw
UzIRCeysE32edIwXQsY9vffw+BmeWC1wSBRKWROS50Z3Q/Sfe+3Wd4QadpCFpB+pggBZrV3B5rdB
IE0jDCwMe1qOUBoluSHNJk4mE0lQ5mRhftWTIyzrZ+p6agJklTRbjucXCzJRO0OaqBEjTFifNOyF
iqTr10n9dG6IvYglA2YdCuNRrUSp8/48uYOCMTBX0HqSqd1KETL0rZJbteLUu44Op7+gXcHvL7+Q
vd/b95JMV9ggJUvB4CwdbTak28emfQnvegSj0KeW7hanXGh6JTS9OS2VhaIsbZunZHr7/UkT7442
uXCrCO1M9Dyuc7s6BHwHq5BrsDRqEmo6sggfuAdKa4/uBmlnQBIUApPnibif4vlVxBnVe1CM+DJP
8AhJxKGaZOyXF/UYYKQaWHmiDkugtCywI2KDqxGBB4k1uTaEHb7vHcdXcgiRj6NIEko7h2DkOrzP
BqbwcWttQM/WkPyH3X9DfTCuGoxzGH+aIb70FDsEAMZ5+tXjQSf7Mni21pOouUpa++JOLtb/T1/W
XtYetpWpsAYHkNJn/DrEsSjaudMFCQye8XYbQtA7Cdjn4B1yD3Jl5LF8ZXMzUN5ggEgNXaRH6tEZ
IJFrpohdwxqDr+LnnBxxaJP7LYRTSBri5ctdzZ9ecU7Vm3n4v0g/b9nlaPH+I6/PFuoOMEwKm0ms
DPqp6WxMNCWyOECX/LTCZs8MrvKNIiJ7f1ABZGolqDSDBR7W3n1FHCp1+PPNTIHbmWp/y8yOUSOF
fQMg3N6ppexKZ37h/qCU7Qm9Wst/DUQfLMK5Cu3Jvjpn4At9+AMwyN8PK1SH4Rv464f18ayyj9H7
gv6BZS5noZBZSUnbDonOaHuQ860e3q+f1nky7OkI5smnL3k=
`protect end_protected

