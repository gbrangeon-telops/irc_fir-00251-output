

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
VQBfeXA4hP5orKlsy+AFFAe2QBxKheQVMjP9iwMw/NM3O4tSdVMF5nSpUCi2zqd6Xl/0+S5YrDyH
MbW21sN7bw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
NYnVtYYKs1fo/NxKyeagmW8datCnZRNIFQJ52Ut8vKAvoM6z9G59Louyi6BpOXJlK7hkOA0EyUcq
xnrhn5QTbG+/jjVXTRQq5boOLx13BVtwMvklEuJLJaUCJSI1mkPVMU1Tw6P0C7fzMTIVY1MXBSgF
huHBAAQ6j+Ca7SHEJMc=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
UdRiCUwOSibQJYHOoWlsqKR136XIPiU7//1vC9LO+s6bwL8gocVodj06NRrITDP0xKYK2ZTek7T4
6OlwV+xWr4k2Xf/sx0trTcVrHoE3bps3QkJHk441qMX8BKjF5fCXU+yOMX1xkQlvuWSD8+NvN82l
uzCDbBA0KjOv/IsJg1WHwqG44dahfC4qa2RHQtygQ4MsVR/PxcN8lnUdpguLi+YyGmh9q+fLgQBq
cNHly9YC9ZC1urY1hg8yqWcJm8AuonE47dIMtl55BTxzCygZ9uoRy68FfVsLU7NHg3O2kl94A2uq
uulT+/Y74MIANEyVFkVes/FR1hhgCPd7uNhwkQ==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
tQM9oFLCOLGigsR+dGte9FyrpKbOg0a2HEe24uc9a4zzPMiWT4Zq+VUMyysv3hVDjsM6Rhdx2y1P
MMtJydYUSv3+V7JQyYwaG874Tc20f583mvfsydp9rtOQQwZoTUUdaw84/pibQ9geh55pxtJYjyzk
ltK5Hf2dDqQ0W2qoU2o=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
D9jeI9qTFJwFpVSxwOhVsb671/UONJ+BqwlU4oe+K/dJiOTSOoWnMaaYQ9Sgy96AbPfvmkY1YYgF
jNHbjBYJx/eNgXJH2lhqUlU4xX7po7K9tZYQraj2oMsohZUwz/eLwj91c7VL5ZRmCXaHh3hDU0yM
tta+u+KG7UfDjSpBDQDdNd7gt/bWHfns3Zj0BeTNOQ2o2kTzIQxImWuXKku154pI5L0sF72lK31n
Ls7v+PzriYFrSA6JTTtqAnDF5uCY0O6Lpa8FB2AoeQSutIiakkT+T39fToTawon3SeQIsthaDWDT
WAem4lxQFA8q64KvDBTwguerI8Z6/8BM0gLy/A==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 20752)
`protect data_block
9rMNsXUkL3IcAjyTdafDc38cMf/0L04Wc751LsfHuA9Yy9xbpiutU3zzIXrs/LY0RDQoU2xzBl9g
ffF8lOHEzRhrHERQx104HMrmTOxEPv6/vycevMBCu/JnL13xJMlwTd7iT8gkQUPHgWUPIOTciWu0
W3w56c7zRQGmHjJeLBh+rsnkSj88EHMwl2Dy40Y/y7i9w79B2z/5uuTshT6t7ByRektcXtFuXbqU
J/gayIPLg05ZodF8CwegrdSvIcKTNhZCmS4EkvNSSnOS12kR3KDoqbta39yIhkQdOpCpeM+3UK/M
egFZt/4aROsqEGlN/kv0lL1Rqi3Ho0/My4XbG3+UcExcnDtOvy8hPO6GyDzcN/GbHY630SD9bqw+
lz/mEQlapMoDgU/E1GKgQH1WA/TE+aq9n2pSSxuFit3Gg4f5Ev0kEXUYAzKJR1sFRXVWAg1Fbgmo
b8ZDcIyZQ7UWen8BVtV7O8DxCk9sQvr9G2bYaMRRgORtfxmVgOvrQ5AunMBqLfIPbBkOfWfhXJ0l
ssInRXFMdl8OYu7Yyu4GEOgCo+2OBOm2rqT+x96wUUUpeH71NmIfc2//pT7yH3mNyef76YYECHmF
90PmHSb+QJ8EgEnhU+9TFjA7Ghl0sPmnlWyUSCx9jdF9SSHmJI/7HoMXXdNNa8jHDjlgHxZV0xdd
Vm6Msb7aF4WIevx4o4rW6ows4mG+U6Z3udfn+4QVMGRCioXZjvS9x5nKM35v0cAh6agMOQ4d+B3j
ZQQSvLFOgRL2Q1BsbwWUmWmhzjOwPfsQMZXAUcxyYuCoKmUguZHa3fdnRnyCX142UZFFRgSNdZz1
hVon8twE0DXqUBWq//FfmhGD2x+O1I6sKo+GaZdD58ZZYCxeUJVV1SCBB34qUoYwPML/j6OJZ1OH
vtjJO/lcbumIAO4MqrzfIH+yNxhSOl6kS/2B2eRf5u5/M+WkwBIgdBpV8PBa1d8l1i5cFvPcPs4g
mSDwlu/Uuzkoudblmj2aRIQBwm6zpw3hIVXKPNggJ7ZGrc9mCiV7Tr+wBjt9txOQaBhhBn3BCcH0
yz//SWYghjphK2lI4vNOr/YP+wa1HYfV4Z6mp4DTnQeXB6cvPk8ust6VzlSGfj1eEmuFMSXPKEGA
HBHfuxkIFytwA2mws0vzR/BMwavvWWEKhpk0SFwjtO9d8nKV6EDD4jTWhNOq3rGLvqNvfiyZeGK3
GN6NG6Hbn+Iv7kbrgYR0Xly4ZjxmfikpF1YHZQoRXSREXCVVPoZEhvWVtdYarcwCdGxHF7O7UcEl
vW9hHp3t5wG/9w2bAFFviL/U4jNRSz0ErN/Ex4D3Zf5LoLMfsMsr0wRNajyEhZJCWvuL6yaIVgCZ
tH69pnMWIYP2lzWYYiVk/lR5PHbsrIcQxnwITD6iHCFlsnEEdl7UbwAuZ/MjE7xc0EapGWZdi1Mx
asrK/jnqXan7F+MXJhYMrZdZyrhrq92EzA7LpTKNmGiVbaKev5Vt8L1Tqsr9DYxV7tAKBOy7WjC9
2UAmV82hd8FXqiwJoj5Oh5fnFYQ36y/8VsLDLMkwSqF5vnTk/0fekAyJkGqRhNT5JWRbY4ev3xID
HqTdCtZLyMmP1XX31Awmk6VOJsxRVmS0paYhyB8SbjDQgZBodxvqg3jjFm5zCT+PECOItJYZo/RG
dursW55Rbr6Nkp5h9BDLpy1b6KMah3/sKTNHrhn3lwgNLVATmiGQmHWaQl3+6aZ96hdj5DjFiJZR
fd6KLfSTYFUCDw3A6RsH3z84IRGKe8fd68fcQN2VnxivFHlg1UiSw8xZSM1/g2TlKjDt+7DSZO0c
XjRk0xrGIEQN07xLhM3a2TyS7XxOMM3Y4wjUiGp0sz25UgYdvz9CJSW9HWH6GG+POCy5A3NlLAFx
UZBAwXSI6dAKHLnK3nyDLTc9faS3+y+xnwRbnZ7rELOdFXjor9mwSDXx8uClymI5arVX7kPsUy0L
xjzeMmeve9RkBkMGY+Z8vVyGyBcy6JSBmIJSoN0rgn5BDxE7OnhBYOsbTppPAO/OJLUffXJKMlkW
pRNViIsKfJ8OxFw18H25HtByoNJIN8TAKwpKR27xRoum/icOKTu4ugDpCw0MXaPd8RqlHpbqKhjd
iCm+d8U+WqGTrKvLe4U0VnZ0Vj4YxYci+QUCEXJB4p1QkyqqGftxsVp/bMmzd7KPRpQwpLHlaTRW
p0NNkuZLNfk4pYowGG8N7x/fwmvwcUO2w1hieLJE9jPQFsvbToX845zwgZ6v70nAiKI23D7gWZMB
drjYY8HUlah07q3rcrDPsI/yR4mlXUU4ewRKopq4B0xc9/Co4HvxGzPnjrreZqrQjOqxaFjhBoHG
9Ok/cpuXtn8eDMgYrh8cfzR0tgZF3O34qhCNg4SxvGBW3K+wnv9guNhAml5WkH/rGI5KT+l2o5+f
ShCiv95skFWpk13iJFy1Qp+XvEdrDGbwHF2CL6fYCFgvB+02rXd1LVhVHkyTbHMc01In4y3S/Ltv
db6HsNvX0o0Ht+Zt7pyMIMyki7sWGwV2OP/NhUTJm5d0ODrG1JNRMod1ykG5xkZZxH63OP+dHNRX
fni5s5RyAiel3untaHscOfcctmR5vwmPVkJxPSUuR6DOG2FB+gIN+ozl1SnGQWMHb2bwWPCnj+Fk
N+D0ksVXnZPX8tJdGaTXA6qyRG5M6bIsDTFCjwMYoBaulXadBbo1C7o0t/rb0M19vk37JKXk2FeK
fnptJsZDsKBISSyz1o6QvKgyYKHHN7zlfv4V31VkRcCobOpHch1B1LSXXT9Ae2GXT3tv0F0Vb/ld
rbPwc12c363uBk4PRiTehoEKDNGpWrvfUAcar2vAOGVKZREA1/5ruUMYERu81cQLOQyfdWqQDfhe
T8XiZ6QWoztQc5lqEjst32OehlZPcjhkd1UOhcd5qLtLO1QGSsgaIN3mwxj6Ev8e2vDtCEfjwjyg
uQh3Q8oDvA3hkfqavvZLjlR0r1LDgQyH+LB8bRQ++KRXDClcNNqdahwr53ey9CXc9ftYT1pnuHN9
gKNQQR9PT3Z/yL8iWiQOUiXdnyipipGFQr93aKn7rrGyCkoDylmOHu5D8IwJVLuZ7WnODhP684gq
dme+XroTX91GevKEtlGYHBZAAShkCDzFqr7EqKRz2Atrn3EAQzXMz9CYdPz7VfUknPymnxemNsWO
LR5/INYegTiLfp90RM109ly4etknV1x59hhluDxVpEKjnsYhOqTJ0C4QoGMoDDGbCE7qHZNsgJnN
91AYULljuq7TpDM9SrKev2OuGBHYDO0bhrG+I4Crj8/SvyFxr6v+ky/A//RQ9kRBYFRTejbDPf5c
byJ2TDoamZPvWppwBqlNlsDpQKKNHPkRzsNFUH6Q2/zlFBRcnleGASAaumGu+AFaOWSEJP677KbO
HSDJ7ShFq7W4vTjjpy0gKlgz5qnBpvLMuqhjY+0G7z9VXUjWZd/ils6zNjqx/uLFigdn7jmWZx8t
om4XeFep0Q1xut2pUyREOXEqK2856tI3zSSMHV6CazlMrLiWOcbLzESj3fFaonyljZUrDmxcV2II
8vebqO6caxjnwjmSDJyNxg8R+YEI99k9qRwbdNwLXlTlBTLoryl2ZcLyRlcKS+EXxpfuPTgoVly0
iV7cl1ixxrByH4OwnQls8Gh1CP3ngQyHveNovvmKNnVyIr9PvVIod4e+DYzONmj7Zs7UZD0tJror
Jc8xaIr6+sKNuMzFv+Iwry1ySBslptTuRYChBCPQHwUQBpeDr6T6Ujgywd8agTQuZHf4GUmB3lB9
0TLZo2gYYt/RPQ0XjTLi2k27Kovx91gijgoV8eCUDRedaIQ9ch0z4oiVdUYwUiA4S31xkUuQYSVN
+qy9pimTjsJcpH1/p0x5/2jn6RdzWf9iW6r6igDnTjHNKVQAQCcpo+zSZhH1D20Hq2ptVV6hCBTm
nKUqfcolNdvrEPp0O9KHePfBeooLOz/i4Fl4SiTcEZ71xcpK6uzYXyVjbAwqPZRkHv6i4yiKC4/q
/hCnHOraFdNLZIf4d32KxQNLNBjBpkUxPjzgFZhw5LYIdkwY/Fog4h/iIHuSIEodU/y3DW+Hflo7
/IY4Nxg2TKfbXOexiBAWCkfbTAd4np4hnmY3PwGKsa9Wjv870AG7w4tCAoeVx5viJsoLKn3mASOp
wMlBMII4cQaaLiuAZbO43/WF9If3x2qKxwJGwO2GzTg2gNij3QlJR7JAjxKh1xgBAZPOfTbU/5q5
VwrQzouXCmWNZPSMaCLutTEtmrXUlyp/dOQbhsDJRa7CqzMqul31KKuTAS6sbrWMlYb8XCB+tHgu
4PMScHwvWvql7Hbrj6+IhSa5P5lTurXzyiDGmiK1AU2gpYutEh6rcTIdHmsiWCgje/t9D52EuLAQ
dnq3UxS80OsDZCt3NneDKL/MDUY7vTrfuJcOLChBa9iDnZC9YT4MtHjTBFpdDVRkaKZhezOuQv7z
kReRycEv2N0tLxbHyGo/VtmikAA5VpXlVkzL34iFcRUd2ai+eXnc1V/K+kfzMfSfDUJRKEHQH6c1
hrMb25J6SRjfG/NhRCVX/906wLAnegztZMPfTDbd/3H7FGymg6vgsmg3mW6doDwK3faoaVVebOOB
ITs+iVPWddgudFFI7DzPUZI1kts3Bf+EWRp9A+oKcYhC+pGF4nxQc5oDzHCg5i2/RhwQZPztWOOi
WdMVaoGZzdUIRzMF245klsgrXTzJHC/RfAWv2psyuVwR59F6LcfwCeb9EzSbA0thTUhfusTUU86T
QVjG+P/npV/Hl15t+CpfINtN48idugwGV9LcAeA6RbbKDv5M5EamyyYRXExjTyXbY0Pt9rxB8oAN
8HFHjfZribTSh9J0PO9UoFtCF5LTlwzJW6z+UpKcDOgdIi2ggTh5i91zR9Pyn/PlrcgD5dEXRucP
0xTTjMAaIcQvl7hxcON2XLN0qWq3Lr3qmJzeTj3AEl9sEukcsJAOVCUE+dDzVRnH+hI9DDgZiHgy
gnPjm17odDISUzSeoTSE4MEOAdTtGy04WWzVNhkhPjekND9kxtgnCVxDc3Cn6hpEkdVbZGbBcYwj
S9hGfTCnOg538QuPL97RrC5VfmhuxuQ/I/FnGxx00wZxEm3TpKyyZT31sBGekV7ZVf+Xs3av+MGH
BFToqksv+i7/GrVR2jR69bA/1vfNh3T4zJ4tFzTdAf5Gqq/NEQxQlYWbB9p/SH05v0eR+F48pLmS
Uw1gI7Z8pCLMY7oNQA/ay7S1bNJpW/rg7wuTHmivPes4bHv9G09EzlqCu1f1LrstsVInGlZILiAI
jW5S//teBnIqBA1nuSLTxEePQFx+UNl6UjFhYZJ/pe866l/7k8JbKXqSyBokDHDP+Ax9pp+KUSHy
79mpY4K1kj7AROEEoDd/boos5V70G/mLAXwb3PzFd4ahbmFht7+w6c/Ct4VPnMygr9+sFdfNwlFM
9rUF1WGP/ogQDylAamxDkoWbBR8XfmoO8IDqMQQbMTRRRp0zGJmtTRQXCt80cuRTPllggqkNfi9j
6Ft/UVYazMMhPmh+jcF6GcYbgXDhXQWXRbIn9khs0VnqDqAP6ueTNEuZL1EZUbmqaXLdtqpgQABn
mj9DhUVitwC8EN5RDKUXKLEccpUG+syHqgDgvOfMDafJukrjPNWvWCzCYr3SorCZseO/5EkR2dsN
mgDkp8pS50TuQYkHasUTFgHnLF9mTPbpZFb0oGCkdZdljPECv/k1f5KknE1GaHaN6aIfFv32zAtL
dko2B4WQS7C2jmc4Z9TemObuBuRAUZE5WuoGzxZBmECOn/h1Qe1sEUqnTBE/t8v6ibBJ0T24EGvS
CGszYlzV15RKJm4aTYEPvnHRNxSjlMLqSimA0bUu2yYtzl4Kmm1REfOgGqZnA5iDcBClWTt22uVJ
IqC7KRdMrQeLejdtEGFpHlCIw+9zxKaaundtZ1aL1kveNhffEFarrKyzVyiPiSyUgjFZqBXU0lQR
DXwDfG9OxSMAwt8WNP0x7YzKIK9BkbhkVqNB9qockZiI2Pr/o9pFrW31leKI1g1+sdSlIqLHfTT8
6mZUdzBjvS40F8ifVGATLQT0ufBLrDuO1CJbyrDZk0kPr7rn9xSaZ3tboEQrS2XYFzNe7WsFOWsa
hSddxpvaGMMVGyAPEBGgHET8Oq63kydzGqkVjBWdiDm5XfuvfrVyJS/0nhJ/qY9qcwYWBW+oY/XV
KngfP7Y4RxqnuN32xRFTR+Jblk9aWIAn7W++22iZcVp077mmD4vus1887oCz9g3j0Q9zpyCSVJuO
fe0XT5Ydei0Z0XRoakvqcu2pTI4Reiun9030jvw/NkSOyheBF7htJsOUtz5MdhRcygBK9erRBOQW
5EwlcZqVm7MUmL5zH1wNJt/uTb1EJTYU6Y4HSXqFtbQwENkQLSz2IDVXfLGBHwqKtDhqs1k88klc
KbjfDf3PVhF4zRXO5o5NLySSHvyO7FjefAC0QWyyZf/psTzH8sD4VivG9haSnv83ds0Ctv0+EGAX
Db23CKDM5fpmgQhqKSA9aOvEnct/1cN5Mc8NmqY9FmCxUzKc7QIe8OGfNUYq7oVdW9Q7rtgw6wvW
EInqXAvmtK7379oZL9+znF1ljk7mMELxiTBNWTzkef0dqsQP6UGxoZIKXUgEbsXvV5fmWYq7/afv
GPolOH2pT2iA+fce9oxnetF3FbkVW8BZe7ChkuvuFWOR1WTn+jMFDplMwHhNe9doG3K4BLy+z6EC
cBNkStCOHRjPfhxPYC/u5AmTJ5WLPy4QHOW1sfyX9Vcel3e1b5K4mV8FkWruaa1awLVKl54zFxRX
cCErI2XRRYeJVPo03z9sXtlfHxmTVqcxEzk2DcRYKmATeUPZtVLym+h5k+awDwGPO/cRQM29Tz+Z
BH3nRgE2FyUOCVBl6hfsyWK0rZtlP9vfsZjbiiENCDS7j/YtLFCgFg1dvJ0uLObOeqWFelKwrvZv
Got0bK2l5TpYb+v5ocuVJ/77DqGNxCW7LP871STnE8/AqxpyX1v29DvuN9NAJ0d2qtxfOo2lCq5U
eGTKLE7i8SoS1u3+iHxaHXaFzXIGiMzZ04pRHrv/3tpGUO6ciyQ5oyB66zdwLvX50ESCfLLeEjMX
usQV90qVI6D/3ZNoNU88UOn41UwYKP7jKbDukFV+lATN0f8p8rGItOqFTwlgn5sZCG3eo9qQZFgv
KFxE1nOPAh6T/OCQcQgVdQBWA+J0Bnxk1RdrbxMIfPpHvclQNtYmfj/52hEN7rYGzQ1QN85n8xJv
LCcSUYAn7rZwSx3bm7+89K4IH4mh/6ZStIp0V8J8t81MM/isT3BTyxiWriK46gLu+edq1o7NlRLZ
m29rv0lU+eN9NgbBmRY9QWsIYj3QY4icJ7mKko7JJmN2eZdzxPfsyrT+xaq7V5OfTuliAL0bWxSH
lRWO0fvSChvn8zEBuFM4zo6gjz7bR5aA0UWv9T/7qZTiHvnqejfzkQFJyn2lSfBwrEdjgmTS9cPS
PTuzVo7qCdLByyUUGWIBsoB70AKKHL0Vql7gb4C4UWf9HUygoVgaZgpBwxvdKDAWM1qPb6BWuIaT
hEzliSK+Ailjf+uMuickrD6F++scfDw40jcprm7K1fY+ZIQRHJmPUIaykD9R5WvvfHL1eWvY1Lat
OLWYSG3JmfQOYCB7z1PqCKvnKR1BpwdAkc9+DxwhWaLiYMW6JxzAEXHPSHXa3bJCTG/1YXri/A5F
6A/07FhJhnrZnHSlMR2+w6KkWztCd3qsKvgEHN+Br/9Ha4YCFq8AAuwxGkZIlHxXpNwFbtLOb279
SFnzyOdHV+5LmoJCc7Z3lpRQ0A26cfr0f2R+RG3wZFBSKLtgHUz6tpqhLhNnv9TFcfC/1fAJoZHQ
VpumwgN2FMOl84sbM6dtttE9zJIZQd7KFqIa993T9iOsW2kNbYUc2bGouuyRx+Jn15PMiFnDqyOs
RMemHqSeEq11AMQA8SAGr9Hl/Bsm0jmwZP6Mbb0QTpmQyT7P38HKYvcfsB5FdIscyJwQVg16ulR4
9A7InGL4V66RDi13EFowPl+UM6EPa/HzsOzbXhewNNHJ5AhlS+lISsocohbW+d7Iwf9bjdnM1xyI
3GP9bT97cUqnaAbPwl7/XZWsmW9Gd26YfQSiE27GHu8AcC1rAJ+UitUU3Gai2UIQUcmOG46qMw4z
qyozFjpVfXL10UPnorWr8nJuW3QI9SL1DSj1RAL1b+JztePMXxFqpaW15SVSaDC5FUgwaHdo1d9o
qvzL3Xuca9n8viLwrtiR41CaiTHrQN+kMoZZ4oVQ7GDgqPOzQzL4jl7QI7QpPMEUKR2qpIul/KaR
EmAPeAlwZBS9TdPNtceE5IN+3o69dX8QShKCY8ZDnX83QGwloa+LkQvRPknydcG4ak4PRhpoPLHz
XpsBcVQ/CyF+FHNCmlxv1aZMcEX83vUk36XSrkkk48FPrRxVz7YURfk9S2VLxA2+LsMN5vzCZU2V
6bXwl9qWMIZEqezougdiX9+4dSSL62UzJMnkaUuJinL3o0II4fyynuzqePeM+L1UYfcTJBduKITe
7OIUXAw7XiOX44XHv633n3kE3/w3t0tXF/OGaCX0iMUc7i5lkbu74CsAUZSolocAZo/FGLft3W0v
ePAjsgcDc6cpe17QsaswYHWNwYrrbWT7W7Dk+FyfumNrHWQhkqAifep+pgUlc5amCV84EPyXujKw
84OEwjRxVOl88c1Xc33NZlm/QtX0LOLKd9HQPQSfxBaPAQKkpNsqAFHotgXsqCF4F1MqHmacAf30
uOTjuFOT0Nn1dy+Qcl2U3BN4Y5hGK1HRChsVTbwFTYXt8XuIQK1e0+Veaa3esEWSxHf2q/1GXnHu
5JNeAGdso4qFkUHCO41Q6Ve9uis5V1V7aHClxvmMs0BnAPw2x8GYsQS7OQu8novS8XFJRgiNO4ha
hCEPPp3Ov59pkMa8k2pLF5P8WQz6ZXP38XhguocKZz4sfoW7o4/Yx0e09clPGKu3scQCl9yunOKk
8KwyOf4Kf8uV4QIPLusq4UApKG08KLk5ifq5nWhxQNeBHZl8ejA1FutyJ+/1cAyOI0n+3sQdf0h6
n1C8aJx590s9n/xqf3o1n4xNX74Q7KK5pNYgt+A57v9eNdRnfcwS9oSSeb1kdKsi6gJPM+Q2KOeI
elvoW5N53vLacfrYggcJoPFj2JsLT2dhjs5v0wGnFDpJVCpVfaFQ6LeY67aU99xwgZkf1NqTS02Y
v/PzeVSpzZ0VSGrZUb2Vgfl1hmfLDylpaoRUetVIJGBVhuqQfcpMxT2OhzF1N4gKZ3j/18uRAV1v
AcbQBJl9YvLzzTTvooN3BAFCPgrxEB7Q+fNQ9CtL1lE64RWHdmHOjdOgEo9BfUSDKjNRy1/zlsBt
FXzUpkNvJZ+qdK6cT1pnbCmZ1YwPz9lXraO4+FKc29XigatFbHNkLqIalYpDGT1CD2EViHQc1uT+
aTrGukZEyWnNYeXRR34DlqXYgaABgGzb9lU96A468GgvYOkW1hdJxRrV/vMOgL/pyRpsfXDF3xMD
bXxkYFkQXXkLR59TagGyWLad9xFgbSsE5cGz0KV90rjZ9ytGJt2hM8k02fFSxnjuSVw2ZfT0rXq4
H4rUG2PJFaifqySojBNF8cPBUnOVYge6GAKgCNYqeXlSBOWIoikjtHdmeYB1wnDzg/QANdk7/aDk
C3l5GoYXbKng7fj4YtIH7+dnbbuis44yYieEOGFBgHQ3UQarE2NHiBkNYn62Br5suRgtjBHI1lGE
bpvD7egbeyHSc/J777p4IRj4kIgO65DK5wRgNMDnNtlUsncbvKxXL9pFH5PI4LOXxdAxLvrDX1/q
Uk4Ih1WTTJkg/rKPVEpvqUISln4AYcc84PNe6ytRNLYTOWYmMnLqsRMMjuATtPlxYmm6FX+IGwj9
HcQSyILa7ZRBxHhp6h14TbsUOOnhPxzPUVd9b0y2jSCh0ESxUt36Qmj+z7Wyx19Qr4uOu4ydWRM8
YpBqluxhrj+xs3YI2gkzubkoEUCEMyQEaJSVezt7VK9BNWy1jD2t/AftePzMSjJH8PpwH4DB7U8F
0iCqv9EvkAzA6zZYbM0md0rm6L9rBvnCqgTnpn12JuL1DhIKuUq1hcbQ4HVkG0hxsJVi0B0Zd1SQ
nStZom+X23q4Nz3UjaX6koZqbjGTw55x1yjDAK4Qk9xz3uRldygUwsDpYwd7W24CFXJf4Rg04ICr
NoMqtC9L+aPy7N3MF1yV4zs+ymM6gUUxyk12iEn9Rq8oilPYfTTrWvaiXPxCGchnLPHDyfS5mejK
lAppOYIsa8OSXpBskLuOFvMycwKCq0Zlglgiefid30toV/xMBqk3BzygnsaaS9MZCc8Ebnttw2Wl
LwjU4EsRsGpUYpduz5UVRgjj41+DFDUgYDLPGijOjDm4tpnwgP2B7szvN9knRYIRQvwd5/fSgfPm
tS/SD8bB0SSwGyCLKtAZ7ExEzpcBAr9nzvRnPGzSxTf8sZcTk1Vky+Cmwdk5B55ItFs/Pm1hq5B9
eiUHP8gAvKdXG91YmGbCFV6spdEz+ROxP5i9U7ZSIM+XaD8bH0hhMm2go2/EpCGjfIZgxfvw1YFb
VQBecgpmYykq96V53kVBnQFpwkZY89kEdvKRLZCgE0aOkdGp1G72oLEeIakqXWSTLasSwV/nSW+5
mokaTkWWRNG/+HLjk2uaTq05mLPF9pqUxiUVLXj7S85yEbXARC3a2gth73mCTb9zW5TOUSOccWOP
OoLxi1RYTzsGKob6K+NIxAgBUfx2I/WFUuGuIeH1pjqgwWM+Fw7wymuunhd7HOC/GXuUxxcVmA/h
AKw3L1oLEBNhQQOueSk+ejoOJ+JVmZgQLi+jy8HP87NQ2L3EOAkWlqm1qzAQ+Tpmltp8VcVhG9jN
DSY+1NzTvTRughnkuOyL8BCsRwUGRlsOGyturx/0tzEh/u7VRsyn4bsvEto52Wb+yqa/LuRE8Weu
FzniPhcgtyVFiizxHDAj8HewyisLRIGwGRyBAuLsm17kcSZESOnYGLROaiQnU7XLEr564mRM9hb6
lmhiQ3TOjIY6Ljt9O27MLUp78bNdCV0Q9p0LNrKuJlZa5zDUoEZnJpzhg9sgSbl4kjpMANO2KFaB
uaaad/1AYPQSrrU0Q9jDfJb+Fz1uRQwu/uAfbxDsLay5OSPeW2nsCXqplRCmavjeQk8vnSB9jyHz
TTp3834XIfXS67I2UgA7BVXIG7rEf5e/V33+sW0F+tZAUXH59CX1qeROAjkqbl0tXa6Zs3qWshTw
O1wCOzpf/AT0/Ext0togm7qrBuj+mPdJp5+yEPmnlj3QbzqlhRVeBfi+z/a+4GfCn/QznPvuUdCR
LF/xP7ESCqysOkvwZfSQXzbM6PjgHmJR4Jr9fz3be1IimnkZlQlBsBP+AhFQ+v98ooFMB8/9wtxo
7q8ykAekkqRYe3hfgMQZGUFVu2OMMyjHrIxHLCyhKc0vgh/BMOK6GKcVsrCQDw9GWA+TZl9eCNPm
ZndYXeVZk3ZPXs4fMpFYlowQzpXNoxIaYL5+IWxIrUciWtUG3+Md0JqiF2aUt2+cR+IT2BZlSKge
5TxzWAxOuko96U/NM/XAh9dFPQsVk90KHzqQMpERlkjrTX3xp3tzj3UNS4vN634sGco8XSOFjHYV
/VphUA/Tcia2eO0HhfUUp3FfTMY7KRlqydXig1BNiCESssUQ86nhLU282ODsVLSSwO/G5XH46Xd9
QUyJllcxHglTUToqlEcHlDw1+qLk+AJ1FpJK/C9gVc+KHl7jN/e2vhRiBBLQuJciSaRgAwfO1L0H
dphAIXQoX2T3137/8LeCuFeHvtzHct3GnY4Mu431NA4NIRcd4rlXV8Tf/eAWsxUGDRT2xlCKdWqr
reXhEM/ovvO04RAJSwPImbJrRt250OAODO2H/Af6d3lDJrXN8GD2ZPAx3R8QKOJMjidePozsLkQS
cVD5qCZ9jAw1dY9ELNgM5g6oviDbYzZz2mrXK68EHdBkN+xE67of4t7/XOlqQwWcfcwbJaU/xzcE
zy+OitM1Y0ZW8lN2GgNhhyulyulyEsTFO4MEani81m8Ps1ulo7iXlvR4QO9usZ5uU4s7WeozccSd
3qc1B51HAd/b1MAa3QOaY1x6DQt0BcDnkuA4p88JXRFGP8BkF9emrGeWMHEULcOIeEVmv/O0e3az
rXuAYcDt+A4jZ/2vilLNPOydLCs9n2MGx0WZZRzU9cYLfXIcS/pXVOSJyyJ8PPsIOO69UNjHXBZv
Q+etkpzMofHc8awlBmGL1Qtbsp/Fp8sk1teJC0wyDTrF7Quca5Tb1PwDI6w8UvBTag65xFKtAkMD
yHmhDhQAPE4ApJmOJXu5GpVugGG58oCeijljfxyUPw06qfJQvMOgt8Ss6CNV86mHySKhgu4w57cc
6WB3fup5OSnk/GHwIZMnxlkn38I5/jFNcjkau0ndUBFHWubfxRcw8fJKc/K8RBhvizWYGlnGr9rc
uuZ3X29Bz51EkchAeH0qw92x0WOeesQYqy8Xq4Zy4gw7TqhAuhuLz5K3YWpwi5eKVwNOYEOJQEWt
fA6FsR46v4ntJOU/gybxOIqHL2wkXNDx+s8c2kPVNpGF3nQHjZRNMDm1vWWSdIekBODJ7Z50pHRf
OZGRgmZ8EkwzQil2nz2/dnxwbiF3KqdyX13OhJpOBmPINbEN6ue81GcjiU7yumrhlyOD77frodlY
Z1TRTif5CK5uJB9cnSVttzDoFxsAiS5QCRL1gqrHor2PFf1IMezMwX/G1hYv3vsS5yShpbJoFBzw
nywHrgX7zCbrmMChbz4EwwZPS/mChkVPjMynwUgvNjulrVH+DDURNNcOqYOJLITFAuBbqmoZvtxX
CywM7TDUG7oaZxYaCJLk0+aTOKl3pnwmA+zlMzRXHXxJlyBgMZGM4waZ4juwWBKygKBKbOuW3ZBz
7nJvrWJfdmTy6NVNdFliOUSoatrC+ZQJA5zp6yYtVzkog8QSqihAM0fp/d2Aq1zrtObpe0igPxDn
Jb6tUR1LLw8ELMhnTn/OoqzfILJF3VCf0wsMD0xuaRaBjvehufnWKbWuW5D/6J4pnoLteC5/vfAQ
t8HmCp1dOjYEhFtxoEg5pCtroMir/GRx3fF81ivYqUJZdoIL0aLBSBUOKmnWGR35IlmLQt+lXSco
Ykn9TlvxbWKZ2H2SLZUUgKO9rBD1nsTTXQ0irw1FJulyVeKvKSATPPaoAFOE0ansWaivCqrUI1C4
SdJje8/5Y4OFCRD8yrjCnheMN2p9xNC9nzV919vgCGEY6T3OV96VkMESSCV4ccPfBoIUdmYJqESs
NKsYGtR49c3+rVeVnSGCslLxbcjSu0PYo1nvCNGKxFgC5DpzniwhAf2hKdYwM9Wq/yNlBWKugLzw
bABgfa80h6FyML1c2zzMxWScpTzLbkAIv4VEhlX31NARb4TZ8/atB6dDbTifCj47X6ajDfF0SJKl
/g7u2xOGO9Mq8eoz4CzAraLWUsfWFbbLGfbCsqSP+kTzx/ZHHki3MSd+JAxDN4jEZ37JdOrD9X9O
jpbx575BCHHI+RiyLuxF0z+VPA3k8hbt9iUct4zWMffwsYV/LBP6iqLzmihj8x6z11qHgRYCAqFf
bP9rWg/5Uk34XOIKjgZC3RkjlZ3JDluBz8DOFDiXbHe4mnKgMQL+e9KIK83347gkV4nZn0N1LrQ8
NUMBYkMz1psBJTQr0Ul/AGh2e3zzv5l2Lers+cTi1DVNjP5J8+XZge9o36nPDgP7/bM5yVDG+g6r
BM1WISdRlAGOF29XEb+CPw/Wa2hRLkSP9wT6p+NmO6e2O9u6wS1flNi5WGeJmMbfXcPy/a/FmqmG
uyOX8wQdYuteonbGPv0m7bK96Q0vFvEfSvuXQ8qMMXJVwrMK2pk09ZjMIIkvQCHhPz+CfxLg3f5H
hYXcpOFT2StCvEwsRcP7MV21MoXNrR9+5It1FUtM6pNZlz4xfPkPbfJUcb+pgP6km4VWtwosY+BN
yRvpo/H5nEDzeK/6TF1J0h/XridqazZ0KA0XRhOk0DVhwxgief4wxAmN23KGomVQtiwct4RVgEAR
eQSe8GsOph3SLYZSN8Ar23DumPo8xyhRlC1B9hMGielpTxsYNlvsVR7s7DsjdEZ3uj1g+UoK0v/y
cb17uKbrB3pFTttaDWdf9nqk7qK4OBJRxzI6EAOLIzent/lZeBhF+0Ggs40RmNUwIkOpYIxIbLun
qwHqKK1tIO6DAhTvrwdZ4UKf6LK1QaXWrqraFptzMAdABAb6kUHHax4+KnFOhGslwUXHLuTqMs6f
/ImxHuAgEEZulVUIB7Mcih4jGk+rMCPjLiZvK8sysluRQwbFAzhoJ4q3SSBg6RWn5T3CPDuWEPq8
cud4v2nI7aljAY+0B0eKmwWawBx1pVdvE+bLk41As8sHLWaRA8k1VNohdNYoNXjN8SSKAdZihR5E
YPmF9YywvFgbQsSYWEym06phTIh8vXm9GNcasNm691tagVRGY2auPy1ZH0UAjvv8nPY6Atab9WLs
xPHkoxN7UoS9tEwS+J9jb18Oh/LAmgjEqb1xxdc0lUqROSxzXjYK6/1mnKB2YiW7+22G4FJzOmEm
JIL4pVMqJsU03H96FHBpb58wVj4Wmf+F9UpB+SCTvp4xc2M+O33S5wdWgw0Vh9CLl+b0Q52Ueci4
biKbyY7FFrnebwsgXI+rdYLjjTO1YuhmR+ldjzoBujEI4RSKhvV9FQiUvoSOS3SWcnsggHuPW+0h
Gpd0BH/fDE38cjO5rFfq0DbxMplRqIsivPnQrb5cMtks4PLT6UNPjzfz2phacdALKBL+YlmXsLtC
HVlmQ0AyKvakrThlBOfqbL5urlRv39xy7yZw/gkL+dNgKw7cjUHNOPp4/ev2VFSVIhxrMgL95rNT
UGh0SxxggBuUKcT9TrzIhVmAnJk0eCNbXzZRcNmzf3dVojHY2qLSYtnW9nxJQN3bjr2yYBII2wf9
o9/n3W4jdt0KKyRhEj394uDFp1enKWfmMzK7Y1RlI40TCN0Vx9MrQMThaNJwq3mnOAA69DPuKU44
6zOHCKrAGWZskcbngxJ49CwOXIDKDsJlXjMturn1+ZNXn1QBBpRGkXP8/UGevO36TekeZjBxJjOP
PmYBxuWmxITabRNSgKhh3Rl0a5UkPqKs1u9OAPeRmXpnL24wHYVlKzRfytUUENFwMAqDgO5++CdJ
U60VV14ODWiYMhrFQK3mK8vj1Y/S/GxsMAhVCpXqZ6KLN+1renKDhtJYWctatr6zPp12HkFctx4h
y+Sezn9FrOw28a/9dMeKZb/zdHbdVWP1kbiJsnjW+2T92ALE5MHqzHujQEGf0UV0S43kJfhA+vXm
ttXzkWR//vSPXqqiIjos1GJHlhVaFonyRcCls+Z5pogE0aNz19/88Ou+CMQNCsLXVACWf6qtBfxh
9lpkc+nxE+rLL0dzOu3XpqDU9D44FFtQYkxNUjgVT6e1CgMzdVJDyNffEEsiN3XHLRyh+JaglUOi
BM7QxZRmx9V0JDXyDxF8zl+x1NqYsRYM/7j+wvOPl3YfZo1jPOK55ZWNy5tU0MfA/ARvtoRnARXC
PQPV03Gs16b+C9W6DvNpuJw9P2Ukl31T0UyDlvOR7WcjfRBuIBASX5hQ2/SXN2ueSrUYvn8FADb+
z14EC7dmfA2g282+0BIeWiboKgg6fJYL6TnmIc3yoQ8aOlzL+r8ntx9s/L1dwIMPQqU6zrNBor0t
tJDiq7sHlnuLh0+5OwC2YdgzlS4P/eCFb3g8LvbsmqzT2GaBddin7mPnhU3qvNBGx0doFVwI1KaG
LSXqcR8e4lmGrM6FdqAglpt0+BZhclhbgEHRO05ykTH5yzTVURRE9U8rUiPjAEdO936pUgSYsyiy
3mvmxwGZRBlmCCrk+tArix8iVcSf54vDWE3f5fx2x1GbRq4PiH4rgFPojgQ1UC1MM6Vw6MW7zr70
E5NNnkNHqIVzXZQc57jp+WIClj7YKxkq6jjT1Jp+yFeo0sd8EAMJin3HcJdIRiuEl28cBs0MGqrW
o42cV+P82KrC+9CbNo07CbzaDUQIFD6FKcZXwsJW2OETwDB4Z3VzANv3+MwAvwxaRyC8FMgkaHpR
pgN50uMmXUXYVJrIOLSJhc3/2urz7F7ggzyjpvUm8DLlE7qWVOwamCQiNgpF82PJE4ZB0dQPbEJ1
OrC/pAVTP8o7CZbYBBRouQ/XAX2/0pMA/EapT7HOuj9kFfVDdvmP+0moF2Ntaj5EuNXxeqoaTGQO
f5yeN/zewiFiHVMnkDLFi4tirbMpVDB3HfShl8kjTxAm1O9x+i+igBIS26HczuH2smVliHcAY/7X
oRd9HmQrznPAEZTLKzj1QHiKn+FO+Hcuz9vE8NP5LEnv2QrkLuxTz4fYpy7kDBNY1FviyyJZi7hN
Wik6kIXzVb72uABMpTYxuKP2gLL2sxb7+GDZ05ee7pNwi8lgzUUL+SbAxO2IzDYIoQEFZwL8Br/M
ofcqKxhQt8xwYSI93iR/3iAdIYn1BPZMghkMFcvzZAXWmHykr8nN5Tzv8Xmt7njomfZwPEB/VoDt
wc7PDx5/53x572tL2AEL92zRWh5j3eF07Z4W0PePwyqHmRcjQbZUCUywuxys0cVakajQqRkrjBN4
jXiSWzXu6TQjloVHYcz6gywLDjuhmNYoPCYt6/Gd4ZWTcCjWNdqmL9ZM3S+6QkQ3nNxyhlX5xn7Y
6BBRPZTivkAIoeAL9QYYuW9r7tnPw32m7+Uk0mkfcOGeb+N3OuYQEdKJRhzrM9/P/Nrd8S60LyOV
PhOWTWbpD7EF9kvCSMzknsgouUt5GWYq6XMpdAaKn37ZOMbif3jrOisI03VtN37SUEGKYCs6Rp1T
ywTsrbQjTCFiOnA6s6vQ0SqlN66ZIZNZdoXSfQhJAFfbysIHm5DB8/NhS7D9Yzg/FYAIn3y0GFUK
PnGdw9DV1yC7vxCviFwCDt2VDH0qyKh+UAU8s5hHRnYoVB6kBYeTJmRnFc04+CWOK1pjAJ757jzV
XE+HAdv5iK3ege5IPdw+Bpqf7xLnIHCsHN/61AKnTxZ6rR20jkR6lzulDInh7az+uDWH3/8OokC3
1QBwvdPzZXeX7qmkoKkvJIbzGToplhmVBGEU0L2rvfswW+mti3Aglfr5hxq6NSrBpA3dlWrUDuiV
HG3DmkR9u5IbXQ+E2Qc0Pwt6TuiG9FF/+GxBYz8Pw4q0YKehCINX4XTB5jrqCQ2/Egwp6Nf7fA/Q
50yHpOgPxaB1lWYeYWo8/RCG9d0YLfIdtOOmxr2XFZ5DjIsgVJBOO0c9ihMCP83KKAFc9RBtswgm
+majdivSaen/nnCYnIATD20Y+DiVhDPU5V8wKLzYAGEIpQnRqWEn679zaKOi5CdWBkqqh6hxWBCw
xs8vs+2cSJVw3tbrj4tOQDM3YmXtm9InGoQLeSCEB3M28VllN2oHq6qOcMHrI5yBkv6+LYL4hHWO
DTW/Q/18vw6pTpVsGVhse40bAIyMHXpXzsr1PM8VuIksVFUX20nJVNIkBWXLZUU+HIvhCDHiplRl
biq8nYG8YxrY/b6wyr/HCh+qz9ywsvm6RwSwLwOFwMR/wxqsmXpBD5F2FREPt7zNt5rGRDe7MH/5
wvuKTyEj0lL35R/c1zXjDYLI7bBuyCi/djq9gpPGQVC0J63Q7wP3mV8gsbiw0ikmyLxY1J1BmnZi
gm/hR0m+9AJI+CsQAyp0vKvTWemy+o32ryXho3vuHfWF0Xg82b/b0Q3I1tej0wszbEKcHi+Vzt3z
t8e0IlFq/PoeWZFVMSl7zUWJnL6sQiHAZ5eCgANGm106PYJZzA9y2q3QngDehPdauFgrqdky7+o3
0+ABPmAOJQ7k9c1zqd169mQgZRj9MTMGXj2SCs3YpJ+QNaRKI433j2s7zSBCffGrtcQUbd9sb2JH
byaeRkDUd1QeQGhmi/BY4COagSB/6MpwGCwRQGA7KMXTPggKSnEAVvc7ExHvmbPIvzeXD/T9+/B4
1SN6PPR6R6apt+mvzyvgMYNA/a/80LNWuuhn2hynfZjatUGQycbdbFXMybgG1SjMX9ACq6JOSDTd
V1H9Q+POvNTAJ25Jo4D/qG9wlbAKT5iiq5DJLUlQhx3eodlPBF3hRc/XERfTCsmxfbZy/r6TClin
Qgg8ImeUNbtKZcMdRjKdsrnrrpwJyPi0YHc3rOawcvyMQ9UdgFzKVCWw5ee7xU2MWV1VuAMPmCXr
gHEEVatyVgMdaTcfcOX0cZbBFHDdGCItNPtNKmUt2ZQ48CjcS4gXMavMkf4+6uF+9Wdfa+blCtjO
PwkO0it7mPBupUgpW5Th3Ca7KKkBg/lrrNVlFvGqITKXeqRcGmfDnK+8vMZTYE/xRtQfrijv57Da
Js8TjInuhCm9j04VrOuz/+Z920nBQlhp1YI+Rh0cv9MfosFvDlnFLa/2W1QRx17Ql+O6Hyfh5hrK
kIt6hZuHzKHgehlbCbDs/Dk6aMYvXF6VW6gFUTq8OcrhE4o2e7iRw/E/3qyrjcpV3P8F7fIZJ4fG
zgKi3DAZiYRjZVlwVqNRWhujp9Vrd78O02TdWaCh8liO/gpmZwL78UXqPVRil/Iss7MRY2sWBUaq
eR0qVJ4PN8RJliIWnO/twi0+/bURWG+hSesj1ADoS85qsRjFdOmGmXYp6/pdlbKFi8gSUHo5F9tZ
yCUx+2xmWmeEZaGCqL5ZWa10utVF73vZMblomOPkG5CCR7/rvuKjiQ0YoDCsMhrccy6mOGD/grWs
byJ2OlgMLm8O5vFvmDSvuX3TD/PEXo57oVIsVl56dR2mxkPBwPZHYp3Ec739kEdugFEAU3TQHyFP
1Ui0wt4VFd6eMFpYeaTPdRoAH/C47+uixhoAszhVaXNwuLcoHlBn8vnMiLe1KjR6eHu796bVEtfr
vFgR+kvojyl+oTi7sQPs5Y7yqIT/dUD2y+CZX17+luEunYsphchrvxk+nzzvK+nEhOk1E5q3ob01
hMeoxNyhikVht2hz7mX2YnbjogO//Sj3jiOvS1+i0XDK1SIRJWHVd+IKPN1xgOlYZ3tjg/DQg+D1
4stW+mLzRD3U0R+hHS7Px4GG5LeLznc5CuGY4FjzikaneMNl2hfwAswGwWTRbP5JOUlbkYbt9LtY
q2Z4Yzn+lW+oznKYbpv7kIUuekI5MJ9Fbu2ibY2MrV/kVcQKmpGxlqS8y6BHOihTf0me2wWv1wL2
rRFGpFXE9OTyva4GOYG1rzMvigEnZT+S+2OFyovKxNPwlGjzpb+tEO09NhRz70RNaInB5V0bCZ/s
nJIvke4HmFsTL1HgIzX63iketRNYhZCIhDwG4zYQCTtnO8Ew9+mOtwCr9ufcgVbNXljBBDvtJCuA
cj1SAYo1ofo8SacUaTqIi1x1rnJD1voiRawmJcFxJXQ0gqyBLmPFS+FC5z1Wfm4C1kvgz/ceXUi3
QNXLI5ZgHQRDEvAo9ojFAAu9ujQfCmOeIud17Gew/jy83sjU2w9bjYLvv7aznz2MZHxJtWHrJiFu
6MXqVJPpad++LN8PiwkA6JNqgqg6slx/JOhgvYou+fTRW6FEu9TlyOkE0KTLtv48wofazdY8Uxun
Iy/xvfkRxmR/STpv75seDa3rpNNzDObJtlJ/f4FSuwEEI7XXfczsFS4iTOuW+0J99ZIBW4VeTVdc
qqxDR2C2bRbEyCh/uQDkaAAYFPuNoVFLA7zagw0kr/MamTU/jHJCR9tVbLoi/L/6I4yB6QSdJ9sv
uUwhb6RSlwLvPpFyhgEzAwG06EbIVfe3nPwu11VvKDfnH+nKMFD+N4SaBS6F7XFKeUX9KYnazL2X
2wJShY10I0jeR+t3gpnQUeNiboAJGHtylFnJuX4GuQ2UW9sCv5pQ3zOEB1wgMeVnIcOq3DRXdyk4
LMKKEFY8fkMB9HQhjKjIfIBwUjVJBq5gX7LjKTfNtSHGFNeloPNEl6YRomKz6lJyosCaqLecbY6+
XbaK14UyJf7Ur9sG+ukSbxHzQWPEk/qZb911PKj3MUA9wPUD8m5z+2qEjaJikP/qX1D0X//ho71w
iFIXld5wXiUSKz/gGFFwncOVf6T6hhnh5LBW0nsJIbyRVVS5JvyRuu3I4YIbi6Vl8OXMW603pfbL
oXo66B6wHhZeALM9Yk0ND4mJj1YmN4JCkA8Bi7iwmoTAQ2CngevvxsZPSZ2Kx+86pGdwFKUaeYiD
WcH3+DPc7cSzwXFs5GXtO34d5a5m0PnSFurHK+AfsQGobnFtlrzh1i/sbC8zeS2sXxKR8xwOM69i
eFmrAwh4AO+UEDO77YukDqrAi3VqaT6vh6BMwqUUdI1OJ82fG6pkWBXAt7Vq96HuSUb1u5eKSdmT
Qq3KJJ8B9VzLGb8fmA4X93/qHvwFQYRWW9w4FIOoo4KpFwv4ery7AVoTSE9BdNNGZL0rmQgbeJIH
7lX8HHzFTuiOynh7JoOYHm32fehhYiXDM4PIzWboJmuyF6GrOSxBrRISwKuZIgBir3PiDjydW8jh
C8CGZ62/9pL75/Xhxslc6sTCCSsIVvPbLseZFMCMbU+lJ16rYRfHlWeDYY9lIOsRNs2qhgj8+/mQ
HiQ6YpEGBdLF1Vl9tk/k4lzP3Hp1nknNIzFaKfS0JHs5hLHDP0fkqPxeu4nah17UeG1xlIvnQ1Hy
GybHWyLXs9hMG4tlgAlU9fKCtOQGkbDtDH0EGOusuNK20/f+/z53pDOr1BAkfGBa7C9DWWuPNF4j
cwZh0ChkKh+h5hlgfgM5XWfXT0PkPEwOArbzp1QHEo/sGX6pxOdq5VVYxuNxYCRXLu9a3bk1NL4x
uVfP8dsEYgPgt3xpPbdl1/m1UZaWGROdMhMLhar7e43fa54Mde8I9IaI6UqYCKj17xD5Qfk/yUde
S/4geh8Z1QRqcYsSFQ/a9HfV4wcFd2L+P+kFxeQK9QcflOHI8spK4polrWlGXbYZpm1Pfpzmg3u2
UIvh3SIUWSYtuGDd/l0WGPBVgKwn6lTFt2M5qege+VJAGJLmvMslRyJHPZhx1DZKAT/2Rt2q61vV
M84RXe9v2CAMnXYQZ3znY4TTJxeIZozgz0QGl/0b01+Hoopx80rhL3HbD7wgqMEWLheIYIxocKO8
5Mj6MO9hTn7I7c+Kt7iftVB/ds23ZEgWuTkn5qQSc1OJBnu84qZpyQJgSfYPm2RwdOOzfhIIEMc4
nJLztqTGA/d5YHrLozpVuSAHt9nr/DboLJqFWA9vSaxaFVd10l6Wp2L59nm/DNjR2tw1GBs1rYLj
N0U2IlU32vRFL4jYuE4nIZtyrkn7FwveFlyY/a/zvjet3LSDH7dQsVIcqF/ODKIRi22eauDEEPlU
UTAhxt5Q/WcELspECjLNfmiuzx/Brqwhk/HdEglb1sLWcsfXI0N7npa54uyQIT+UT1TC5/azCWmQ
MKi3S+TcMTflqwOLKsbzVFBqBbsDpdM5L0326uIVDAwqNhdigrIabzpVn0lmgoI8CI6GM2Er33mH
pzvgKCQ6j+/CsLdUv1eSIp3fZVkq/F1BeQkoEjh0y4Xp97rWr63gYVjAWXnC3FzMhIhW6v/kbXAM
AF0w9tYY4WsWbyWHNCBN5ufAZf9QE376mdsv2tQypgK/ZGtOxQNRBQ94x6IipzAjzWFoPyugVC5G
tlcG23ZXI60AAVVh8EQF90xFr4+Q6s1uZ9t1TV5SDEcp3IS7tYw1nlP3/iZVMrhfFNhVB59rA9hn
8lj3y+oecY+sk2+GzAMXVLDzztenTSQDm52k4JUashNi1kNkzEANvCKZYKzBaDgaC/+ONRAXifYU
knqFiTjeqEBq1NluGQ1KFtgjqOhRc6dGhPUHZHBiKCAn9K689rNCUVanyA/qOpUQJzRDy4eC4rHf
W7RUUOtbPbBwRUIg/GKr6tvXq6nsLCWy8rXmo7KBNDViUWjPvp460PK6kYy2Kl/ExnpCd4/9dZ28
59C8jRgApywx91CUTyM88XkGBDyk2Kxe7R3KiWyibz5feJcgSHwXAdgRcWT8L15/5wbZd7GooZHB
l2gSmSIFXTJhNsiaF2scUH/lcmCwZ0vMrZrtlvY2dKnKKX/xphC7Vs1A2e/Dp2JS+6RjmbZ/dJXr
l6hyLZf01bxIBi7PKZb38NQT1Mhb8STV/Vppg7G4y6UbnESQqxy+SJiPEJlEeHg2fFACPKjKeYYx
cSOvQOSoAYoycvUDoXtse5j6OMZGMaIF7VWhHUJrupFN+kP0PLRcD1r+Dv59vg/KxDs1KN/OQ0yh
9DLPFyqeZU2ogUI3R0qR9lqxm3DQf2Z7i+f+682uzjAmHEhUF2NvA9Hi+v2Gepfj/F3k2k/QsQcR
1JN2S980DkFeWSu9S5gNQe2xYGSaARX624DvL9WxtmyVNB9vlvRtM/ATHeFY8b5SWrJZxi3bFADr
IzFidIbsoqPZUmDA0DFS5iXqFHxTrePPmx8wlIz4ZfRTrn2IZFVfxv9BWs4LLjbPHkBE0zcOXhEv
0LYRFmhsafEJYHr6ScHooq4QgowpzIFMlLxpW2sGnQiaMpnE1yK/0A2rLKwujlQzq5zFXg182uBr
PK6LrU9dij+UnIkqZ3RLXwvzeoXxmn0vBm3nylRBaI/QveULqr2Xp8lzVJhuYCd20HFgbW0rUL3R
5Q8h7zU/bNDaRck/5tw77UwH/v1tRQWbTdxib+aW/BOM1SfEUdq4ROMuNU3tDJyDRBGb8boFSlrO
PG47k2R4Gw9gd9rDsVswNjgc+sxjRuw/6yftzauZLGdpyKVnvjWpU0Q28PoCML15723v15FmYc0M
XBxmTvC4tAHTaOv9JN4ngn+7hlZuS2va9r0wQbiWdJDGnwM2AO+XdBBL4tRSmp+vflJLGe7UYNET
djR7OISt8wjmIFTs4hddkb4JJ0ntNvegKB+o26/57uxdZt/JvDmK3xF+Rs+qTozly+UDtNAEiPaK
2vbF/nzTmmZBMZD2BNThu35hECEPfZIEPuenYIpVMTYNyMNG40VNvS4ILdsKuxAU3Rg3QI2CnANX
wCtt7htFi/JxHYg90N4KfjwWCa/Uc5BHaTCpgQBfUgqujVBHI0oRTRCMWbAQ24FYH7BxmEqfThcI
baCU3INKdXAanhaoGY/zYEctCMwY223EIjDkMcWjrA4E6jlaPuWUHQYXADnU73ya7Hb8yjNZTjAJ
LCiKfNEZ2V/A9zWOqW1rX6JR2gvHUbYF0yNbHob9pdsNv2abCYgAU5ySGliMDyHic/npxxJkdKjz
WfG2u+fB947wQv3u3kc64Omw0UE0xh04xAt2DyoS1rdV3sOTV67pAN3kbR4RFOH/ZCEhB37lbuiR
CHQ6rHK0xnXvk3Db+X0Co46RfHjx4kl9CgLWSC3KRFKKvNqFU5Ue1GGuCLHpy3cDBKx5A9I/NV1k
ghF8ooXcngruzUl72SlK2hGEv7pxKBY4Pk4EOidFRpAu8gecNCN2LdwdMcF3FPNY7zjcCYA5S6S6
wI2tJx1fwkR0frmA2KdYxTYpmppMCAXlVDDpYSNgYL7BszAb856lPnwhz8JLtUJd2oZ2kqmPaSuq
a0bLB44acUaKzvEYtLAmHOo/VsTnIikPgcjMMG2q2neQ2TNrmg4QLRlWXUOpdYengoUk9nJFvYXP
Q0cHs+xHpJYwW1DPEz5UzflNpAAsKwWoxdqG9a+oJLckDnkMSYV5kzKWOhXbVsYWk/er93v3ve1O
PILOpy8RUQmSrh7LoJfMGWgP37O9M2gMv+ETyhekvqjsCOmb1Y3xNtQ8aJiYaF3q4JEqIaOrGxbU
lyCjgkZ9RwMfkclJ1AV7JB913HJ1lcbmwM05kxVHjHRqxL1zF3G8JHDTi9OIK0suuQSmx+VlT/mD
r02Nc1QsoM6Hyl/WuRkroJCcozmXs7Bi0mHXeL3v9BCLo2rh7NmM+HwdLjRdKrAVO6zvBqrnPjoh
9+jGHTem1fSzNofeEEp+3I82WfV3vlVYJ4GxlAEPg1VIWz9MnqxA4Bvx4/WUn/wRp7REyzeISwQK
7FYvVVfJatYksgVwouyLTDTzQ284pz/SMFfAwxhzrgQ5PE0hTVWB8ssXlvgzD9bPHnyrlveZkOCq
XlFmvOHr5Quigp04JC6dqJZMnKLO2DHkkRKEBp5MXGkHDmKbERmch8CtLb23l3t+BiNLbjNML1Jr
mr0s0ssopm6U2WqhGBRD2JuWo7PJTp0S2TaouTK4u2C+9HxPpCxNIicuDDThl7Ao489P9nbA0Cxh
kjSJSVC/dWpen6jX6kXe+FQpTpt3G05K11X5J5/Sy8AhA0r/3XELKOFZcoA6JeugciIfiA0TdCKA
VnZOWIn1iBjMJixXGh7WFtBTdDP80SX+7wK4yG0j5OjPpAqkDFI5jmNoVDU4BgkCE4BVjD/S6PcR
vuPaDICwqFaxthVVLGMVrOnxZ88Ys/j/d08Jh6+EPJZ4DxQG+XM+xZtyBhmqSyV/hix75minxqkY
cAwXUfmjOXq+94kE3ubc1sykigMXsO3O2cAZdsMUsv39Zx9Sse+qLQkgkw12k5tQXbbw/+hkdSrM
VohsByGpvDVvpTYPUHrRCxMpLEQuzFkk3Y5de08K49msjGJ59C0EbhmXprqa7geBiGTuuAtxXxqC
10o7S6IWwA5faYnEKUiV9amDzJiHKKXocYzQ/l0vUcSqfsa0j+myG3eieWhD5iBcmLS+l7sXLjyy
T4i0XnFsvdaI0v15kRwvPHCeozEcAfXEU/85xvsus5g6CLvEe5KEZh3OrLkIpPPm52rjh0lFWzvI
EKsofwOKqS7HwSys3hKSuUupJk1FArvAcJ5rSFxi59RvKCF+lx+WHXf4+NVp45bpFZmwvNLn6o2Z
RNfV/cI0xOyP2CUa7XM52vqQJRwT8nA+bjl5CgBiOsXKJ3jMAjNG6WElY+M49S1XAm6Bfb4ztTrk
VnSQTQl/0jXA6Spu/VByN+CdjYPrzjh8ia/+A1UT8SVvpNJ8KEEdL1HkaD++WoV03b1Gk13hy5W/
dNml6YUOEFx/b9b2sUJGW1Vc3FUpWWxxJpQVAwaKfpw1omQ/5fvaIed1XQpteKBVe5zXE9q6OGdg
Jr8qsgUQoLeX1G8BP63Bwt7kjt6G5Km9wVMMXe0ekZHVtWQ76djHLCRcYb+vgA2qfe6qaIa1UjET
eVvpgYDIeqEwzQ6s2c0ydPiX/b/vj++k4oSBDZLBD05iSxd9iK+a3UjxmE3rJWtntE+vyV7vHnf0
u1R7Au0yhwYuzG7DOkI+qtnFsDfno/csX2jhdc4PVFJ27eUAiCQACWB0O1YAXCBziSrpDafkAv0M
+OnUJ8wNIY7DUiTmBPVcxi0fl5Zkk/BFNFov8bHe8lS/o1ntc+rgshhsmG8WW7eGzxIke2XKqsOv
ZrFNF1xpCkxbjxCJPc+WV8m4AMC5zgEbpcuOecxUP4UJEk6cHXA/ikASsShFR94ZkiAoD5iFbNJg
TSP9P0m6AmxMkMOXEKCh4d/4vzHBKLiwNrPRjfNQBDleYUxkBcWmXBXjnqOr9MhEUjTTR5FH1P2K
rGRnTd2D7gicfK5co5yp9WqviDNZW6P5FIPUfKExKMHF8DraG+3hMxd/ypXKDDB2p2xB0yNOvc0k
TcAS5YsW6mM71CkhTnBhP9fnb1wYnu+/wMdpj7uIs1bOjGDGTGRB+NjlXB+91MCWwXk7XhvdIG8Q
L8z9tiXI8SLfGTU76iztDeTr6gIDJukE9caIa7l36KpuS7z9hgMlLPYbYl19gvNZYAvNeW9DrHY1
m76vgKIoq4dX6LGed0Hve40/MJTtt8alme87U6jWbu5+7T+hFFPFO8To2CQyxKiuL2ljSciK2M4T
Ua490KDReywBn8s4Q6f/qYFVQPoXxck1qQukg/nFj9GhxJbjKk8aW1gWjuVaBw+FKYcukknHGAb1
BJr77fmMn8+rU3tMJDli7GXSAGTb9CJWEQ5NuAgAkPYmbdnKHQTMN7o37qsVmQWavPDDHWZIWncM
snJ3JREkvpriNaMtUjTjT9UiofYwpbaDnt4cuEp8CjgL1NiJ6lIJ2PjCbImx0L2Oo8g0u5FGuxU0
gDHdm1NjgPx4he3xrIHM/yp2McqQY1WRXm7/KGC9tpugdxrryVDLa4WqO+bFEtCOgH4R9D1Z21xJ
xZxg6/lCv9sMOFp0ERObnBA5ui4CbsnSZoBWhZSynvrYpuCRX1CDkfmSiGWQ2qt3GkB7hV4rR0fA
1SwPd+v6Jt4nOiBuAgQe1wCkRxv6GLLXrhjgkqvkFHXHjEdl5SjQEOImPYDRbzzfoRMmbaM4H0UI
YFXe4f93uf+CCKrvZzGqTvYun5ED+Y1FHLUuXpoJbM9BnKuKubU3EcDrq84E8prS5rRNF8Rez/JK
+Hvb8MUPMNoGPYYslWGkDXQCfBC5v//A22sC8gO+kdJ6C+3NV/IFhG+IQU0Yt3UcA6XRJwpfaIqH
ULBEohFWx2d9hXUEAUzF7FXsFqVSGB5UACzqxTe/z6qAJb1+SnQgKNpk/Ricehk/Nd8c0hLhLY/g
eP+VvU+ZK7tfpXBcbzdFZn4kyxQ6uw3/gQ+i0PNozDIF/KOgf1r8akUhPxde/1Pvxo3NQ9NiA8f5
E5gjVPsMlynVsX/4DX23pYXCQ15aLQyFxtWPhUIPZJECrPwAx6/BudxMuNVvalSW6GgjBVwQlpE+
p62nYGUn+ZX/I/SDevVVGQLYCxGNqUFT1EE7tZ0nFnLBBLDi27zrUry9UQ9JI8ojYYmj5gInLJBJ
X52TGRv45fOHPhr7uetuaSP4dxFAkM3zXIdQ7GMy6y/dzlpZ1nRLN/zIIUePnZT2+NgiOlXR6HTe
RW5o6DBqCTla2SOzZls7oTJ0SbU/J/2t5AnpnpHoUr6P2zI2TGhUUo9uskvfOennMaxCh4A5aDZx
zxOCDOlgtYk/j59/6gdxA4kLN1pxOouJDJvk2wOl/288e+/9SfoAHFEQPQGXLK4+kvtOOCi6Zr+N
Kw2wWoqHWSI3j1UvHQ7zvh8ZP4/E4x8GlTg0P9DArxFQFFFAw3OXhOM655g6fw6TNdl224IM6wV/
4ABEFeEvD8zNv2N5ObVtV1CSJbhknN3lwE7JLT5on4Ayfcihq5usVhExTsAPSeZG+wz1GmgJrl3I
BwOkY/Cn0VpQ5thzZSD5jPB48meju0NAb63fk6+aMlueT2whe+CLENwBkKmWeGkup6fsTWLT8QSD
h6HjgXLCgjIh22BSkRpQIbM+ftr/5WStT52brCBopUF8SU9Ov5tusVP5Ycb+sxsoJGAp+SVBcvrm
OjttikF/x5+9INdWpd/MeiioyEPLlfH8F7+gxuUjTqOxDUc7dvSEE/3oTtXnvY4KrK5t/THIaQpV
iemn+/z0/DnDOm8e0KZEuY7soe3ipMuxJr0tIrnSoBctFhOJxAQvNXES2JcSVZzRIHwzyljWSNhq
A1vfz7FyDJ0qQIm7UiQDb85MTNCZr7vsE9qxboVju95P/W6iV7q6XyFizDFVB2QD09yGe4BYsjkW
KR6cCYvuElg5Cz/3A/ACekFL8Xhrli142780ba4ZaIWgxPKUTVwmZFfYPoWHLoYwY9VTfmejTDCc
8DKp6w==
`protect end_protected

