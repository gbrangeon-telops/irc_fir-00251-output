

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
DiIoz1dwiCymBJ2I1DU3O4UDdOCD1IYbLUI0voLUvMCBbKM/4INC61S/TdKSOoUevx63V7g+6/mZ
lHiHKW9CUA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
o/flwcKffhg09UZzkz7gv/qZXGXaahpZlLeLvCPnGMHOV0tl8mkXW6lQBADTMwmBGUm7XZoObamg
kh0wsLz7sz0k84YCYY3YnDkU0s6XZ4yFdgj38M8k6+BTgeZETPuk8RfxBp2vQOv9zQhlLgklCWqU
H5aMJF7gqYDH9lzMxcc=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
3XDlc/RrM6J+fMEvhngyPf44nazd8NnlO+9fuAyN3g8+0X5quo1/68MLGc1czSBp+H9Wyu2aBKOJ
b7lFkbCJ13UBsZfTOKvBryDWOFa6KdkhYbTVSV9dfXRZ8PoouPNER1m+r+jF8e7EermzCIExWInF
5NIain6XV3z5eFAoF9+1wNHgh2DL91NQvcMqUhxodAC4EBuf80hcej88xks12032BecjB+B/gAMW
Fju2sqB0/mqHcdt7IfTqsGyFva1zLX5LMPhiF5YeiK1qj1zrDwFPgvhslJ9mmgozdcxNrfEp6yGo
skXdLgGuFnqjmzVIe1RLirf5OErXnL/7fcq65g==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
DYSqibotPAlt8I7+ZHxqG1W8t0MXnDrQyejnExd2/xGgdjHg+z1O251s8cO1MsyRynExFZebXN71
+rcOQqj1RiIoWzG/7+iJR/rcMh398jmqlJyWLU5IbIHCNoZyFsPrWxh/+WMiLYcvsaCPV1/bb8z+
2IY6rcDkaBrqk/EwYjE=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
otEsDJz/b2bcmmVLOLfSwi5yawHEPe/YwdeYC6bj4QnDnh7iDtRlCB8Vxsd5V0BfHeL/WYjoeQM4
255fcpmsdbIm804UqNFTD5E3bD+pXsp5hjDUkd5BI6UEMxrdFYZ33Vo2q6da9Kuh+R1oMK735BRX
27ixqS9zhC9yoKM5h3EFDD4lGv1ah7oo8vFXQVvAoHLV46fz+yTbcdnzjY0CBY6ZcHBHkW/tXesi
gSqE+UJ05pdgmjP4NMP/1EbWm0c/tA0kZtZOMcSt52FHS77tvDYPPfsmt8s4x48hzc87BHtAtJLb
p2k4Bl3eRbmVYlntF4Wojcy6kk0ClpBDQDcHyQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 32608)
`protect data_block
kFqfSueyR6NntGO8C3FFksFOMRY4Lax14nlSL6Uql/uBqKyw97vrQQ/4myp7xhqWyYwtkQqAIu+C
vpLkzbbZKeBpqYM5cBkJhxxWOYiUfV5b44f8rlMKKdtZ/KDmHIMYbn+xA/HsHFg4FSSXiMHtLthF
5n+6Fc+O2PYdqnTayL6RaysHDLqGcKPCHg+mXHDWkXEYRCH6TE0AsIx6lLLHFXq0KHbQ83xI6HxV
TnIwPZ6tdjZKLJxmE9WNzOkBi3d1oMjvS/6atye6zjIcfyU+38dV224z+lmhCtEVAGjt8KEihQjK
7u54+xIRmKgag1m8OqL1H/QkMfoXJmQOj5oYBza43RIWVAOeKIw+qJvrvW7R+/hLHXPadOhB67c5
XLnCE8GHUX0qxZy5o9VOtf1lYJH24mztOX2p/+/9MGDumhGC1GKvax8mDpimolpMVZErH+xWVdW1
Q+SjIzjBIVUborIHK3K/RTSFMZkdQbXp+8ftCKjkj9Rl+tLiLVgu2KUr0uUVN6B+SMUbeWYnb0Kq
0Mci418/0Levm66I2U8cX+KQ09aUN9Yg0v4+fvRNIZSyXM8g1EaGprJk1kUiGD5/FE0AdyLQzMEN
gct5fHV6VmpZ0SWc0kaChfXAkX/GbR6bHDU7NcsuyklHjn1SiTa9B/PWNPjOHrBqv+2QDMGSFgDZ
fCC7IPfenc+YTqt6QhFZ8C6cGgarNqbJIVF/4c9bnaV8OscaWan2s1+a3z28MEr6aJGHgV3IAeOq
Qj5XcqhU2Ukv3pWlelhlgFn0lwBdST5WlEb0tlmoAXaY3z67mpkkxkWBb2Hbb5ERW2PYmwXetERA
3sOzL7/+H5oZVNKN0RwL3B7gt0XN4wg0PDm6N5lu62hpz86Pc++s2zWn2jgIZE6U+ngTPpmRkEmi
2+suucQYIbHuO8tJd2Vc6sU5qbNpODlKVNT6iLfIG2Mq0ioq+8bLW15rF2XNr+snRkLeEKy2DT2q
eooeEJnfV5XRBm2Du5ZXfuRmrMcYeNMC5+q8JU4p15lYAifniLoTT3M17KTfZWsN7Igk282vESbR
FOGY4sswNE0OLmPmLku59UCCv2sVCTRFGS9YyBSLJVmxQ3bWxzQFXmm9o+/GOkOeHIpTC6o4iyjb
06QSbvZn9ZijwaPXDNMqO8LUNlinxn5OcHyVwuNwgbrgIEbDzqoXL5fLwMrB55jfwc18qcGMHmuj
bjyrJbstPy7aNHxszt10PeNq59emRmcQTzq5Z02EuMvvLRIEBAuc7/f/r3CH439Haxa2GdVA38am
GzLo5Zd51tfsuua7Zk430OKRNWlY9z4+ag6gQtMae/Cds259Elny61848B61UWfhnB+CC0R5sPDx
APe+etJN7qGDT723JV0YG5oAasHfj1msprhu7LIE54WjFLYRjTgge8COLnH/lmXXPefqx8a+hQsi
MtbckpZ7TGKTqZgzb/+CW8TRa7iBEAFPboyIJ7M2KQ6arEMbdIbZ7uSCMLHdB6mxSwwHQcyJb5Mz
cFScN9K3yXkPjAH3TB/6HDFzeBmQFWj085yrjdYLHnDkqoAsF6bVksg4zRXz2uvSEzw5dmoKHZDI
drTZlCne/yJ1Exn3837QXOYcftuYl1yY7es63OLyo6+wRRc+lSEPICF2i4QSh5r16WRUWBJmg9LU
Fzds+ZFQTG4M5XRcf9UHMjRvbJeKmGMVaX86J58aMkFEov2d3ikiOtH5Nil65y14GE3AwEzMgefD
zW4yjG22mztUOeQR8TcRBMx0+ywnJ3p1XfSRdELF8YNh442Tiwy4nh18XZ/ngY06wOkm7ME8ZElk
ls9MvvFnEGPTJ0vi0ZRp0s3Nnv82ChmKzXMgBMc8V4Azz5pyAN7cOeuEqYNVy6Zce7MyFO9MVP1e
7/p86cQlB7oGZLz7d8FPlBHaJ2CkncwW1QbBnTU89BFAPPucAwUcxGQMIaJhdMxOgfVYxZckXxoJ
+YvIp0f4QqyYYHF+PBQCCM40fONdQwmlczjgBrN55zYgof4kIVw8QwU6AITUub3GmnBkX0WQP8EL
IAS/UP0BtlNIjKClC2Ks/SZ1cchCVqsaiOkNnHa9Yn90FKm4lPvzhI7OqNS0iI8hjeDN34Pny0od
GoNc1SZH7ob9oOXCKX+gmV9mxCZPTlI6Rc10sopJUml8Th/eyYApURPDiVgfMRliuS9HcXfc6Dlu
iP/mWKkFvlUBlvu9BQXH283kpGMZ0i7igx2yEHQB0GTZbhxucgdw0OnwWyIrCbUEcK0jl6dO6JIN
crz0QGwTYhxU0/Q2ZYxD6NqBVXsJI4Vmq9elrCexPInZKoHBIsSO94KS2DB5VYLXw4lbQOPO3CXN
8PYNXi1D1YdCVfhKqu2ltqezoJybRYqZGpqubv9xGjhYSZhckkJFfqn/rbVvniKzPdUPKE1xXZZw
BgL+L40+Q9fPTGFM1RAy8iRhJBnjPJqErlmPaTLwkIeL0+wSliqzUai+jM5O1umw6tHegE+csGUW
okdxYImevof4YLIrg6mcKA1jEOkbu8Qq3caq17KSuPq4OyO1B8ptvg3t0ZYFnxhAWuWoL/x2+t4+
QazROUu38f17yKTnlyRc1DXAnRvugbYqllbDXGMTmAo+oph+S85MYMeMnZ5XF45s+qQEQ3pZJ5Ig
7pRcZOegYiijtajJH7FPTVsu2xZFZTt9eJ7pSMpncwSLukeeRIe0ZDVo/eWO/zYYn+JmqQJXumii
feh4e4F6ZibKR3dKSNSChXXcn+dp7v7FxKbRrlxrE8Q4c7laRQMtBZzKjVafmFobnreB/pbKPFXm
4u62GVEaDzFX39c9r58u1Ry7J/M/edEPYE651yG0Hez8zSYe0buMy7xOJ+64FyrbVC7HL5APZtZY
5bYvH+075ZBgm0NpMzs9yrkJnZHzc0bYCy3RFrjXaGsFhGGbHGnl2tyJD42EOGgOwIoJXjXy1zHd
jLFunQGPqcNRaa5TB8KAzctTsCidK5BO7BBJpwhAs799Vj7Y0hf0B+qo9rAR7zl4BJNCz9Wker66
hUtxDi1boEm5OY6KlR4u1s+lRNVqAmGmdncKC0uPhNCAyK6fFzL988aJHpYfpak5uwE26kcWJ96d
8CBDXbhHADg84OB3sEKHDvigtvwnh/kmoIZLcIBDpIOwOpFRCQ61VPmddz1ks+P1LbjKfAtiMnsB
hBR2pDONHibkmwrM6Q2U78mVF9n4PA4KvlIdKhe/y4OghFbGHUtwDjvtAWXKHGjfsL2fifBc6I8r
WMy9WqScYsVBaQTBIOo4re9mhSuRwrcW4NewrUYN2cgbgLYpfKLBaMaBRfr3GRlN3j7sR8p5AiJG
tr2ueUggBhP/SbiChKfeAkQD3XWdzHswvG04SRjml0D19On6wGQS6JSgmIb/joPKTIQ58rfWaao4
AFjy5uwgKGy+0dYijct/aTIO75SamSovYeIzRaZZmJrPvBOytCoQrxo3pHtImF8wYNh7sHydwLGN
yd0t9PIdt6fIXs7f6m+pOE3apuJuE5BEXvqyDAD6SDQdom5qt08VQusKpoJ8fkZGoDfuo4CD0Xne
zdjd5QCVA9VxFEJmIjZc7P/t9gsEhoTyliSwhTEA4wczocSQXZadRZT9yH+lGwXKmGIiF8nSLW3v
BVaEw0Qb5XyuLGV+ZfOzBF+U5l6D6DR98C8IgMpZPHTA53xs8H0whHObDB2t7TuQFZh9/HptE1ae
12NFJ90OIeV+7jwX7t1EvZUkMxQ+E+iNkyZt8Fo64mswMJrihKOd+RkzhifT/s5dvFrpMPF0lj9k
qhyz6feTulp2m5l0dngQ897ASvhkJhoXDBeJKhIhtfYz125Jp0qqwRyjWu3UIRpO6CGTqyYgSBkM
UsXApix12NFtJv/cQPqg5bheW//W0/p/EqEyasgeOf7yWzyC+eu6aUrliUyyP9YuhR2uW6kTinsZ
8WCMquL1m18dabsdb4olqQ+fzTXKpgmm8Kyf1JlhrTZ4CRc1lX0zttgSoEqI82vL87KGlNMON1Rt
o93U2zG9i0gI6KWbDy62SxnNXDNJd4FzXXN9NnE1tomRrCGTYf+GGIuYkzGtJhxLwzBuY8GFSBd5
ixxO6BYTyo3qv8t6Ztsv2RFtnsZ6wKPynPwuYmgd/d7XEtkJp00DXhiWwPzQmVdqTZLNW1+gx1pd
ajw448+jijY5zc7EizxVOhR7ZLL+kLdDUNFHj5IzTsgHlJGixiso1aXt26NCYH6N2VS5Fjch4W4O
PIujP/xP/47UCUwYckKFsWC+7xpygPo6dKNoczCxEphlvoLgzvGdQgRhqNrKNnzGxCUq9FIzXDjX
kYqMLZ71OjpUiOLUucNpjTqpu/+IepzGuMvdafHW7vNm5f81Dw7w9BTKAlPavH1FSKJl6uF49KQe
/xpNSrMg+yu1QX8VcCKn+l7u+ZQIuDdkJjg8erKudKoRTVKY3NlFCQONWUtyScJsd04LVzxwkyHT
8GHEhq5RbvqeQkIlo9KOpr+St1GhzVZgLxB6HBbJNC3xjRaKNet6wvMcqP5gQMK0oygGERFoj7Iz
l8y+0mWEKMTUz2s4l/SjBcbT+QjQs5qYh5zj7h43szwsMgCmvdUlo1TIaIGrDZi32k55kakETUt4
gUdlsXjVl2NDmhPoBmkkG3YpPprS8zQB2U4IdgwcxT1E2B1uBKzQmOH86IW6yGXrXflV4lbCqtNT
qeAY+dy4Ml/qUQ854w+X/G8SHVnxMFRXcuwpmp8gvTla0EjwPx2i1af56yAunIP71yqK0YtEpC61
t15oTp+KBdqYsNpBNUgEugDfA/se5f2yp2NF7m5FoPsaiaOXlY8EPJukjucVXt0DpYiR+O4rhGIB
XfQvOmYWqwn3WTCFfBQUQzy5nS+dUYAKkoqMFJokUBhmoAxzaKBnuo1HtH8CvGSVTPgiRq3hfQL6
GCBatFcI+H5Wn+fs2ZhZVeqwi3xmUqsNGgk08VBTJKt8cOyG188yi+ykjl+btDIizb9+ZZ6saN1Z
L1EMAILQVbe21Nmmg82LT5dxwfjT8HvchcMlygIwM4ZE4+5o2kcuRRAnqTiFK5eTACzs8SSGdYD3
OVhSf6x6MSUuVJf9l78VpYxi6I9LP8NZh5EGuDykRblPFAatNpFXiExNMI+Xorl1fJfZahl93J/g
XXBQ7D9u10D9s8WYVpPtq8w5d4ayL1oUnp1hZ91Hjq+skyKzn6+tKLY9umQZ7mvpobu54e49Ho6L
wwkOnfZW4qEz3yYkLRd3V/jTChBW51PxS90nWA+2e7lw2iSsp77ukAETMPA1whObKhonq2rpTxaB
zBxXn5CRhEV/D2gA6qQvcHbfEf13rthJMkTMkdNHq0e/ZZw41X9R3YyW3iTefu/DvALSXFFSjvjV
mlwbjKXdgmA/jFgYMK6IKXJyOOGSgp0VvPBogu0lyWeDsQb2yWPUkoGWg7vQ+fZ54AVpmfIKvSh3
xyqULbWmwyr2mOykpMYL8wFpFPs1Pn2wP7ZPKx7pL3TUCLMZMbVjzmOsXehCj0rIr/LW+qNXXP8d
0u8AbNFQcbihUn9Ce9I6yig0uYUduVLJeo1pO3kKO9vUhDzKcom3jwTPqACbuUsXN2ayxypJqy0r
SQsdJ/DzlHzvmJSKe9Nh5NiVHlcryA2lU1s7Wz/zv4zu1w56c9AAfKkG1c3D3ICLlOSLV83aksHY
3ECPMbjDenhPzdHmSbRSJrJWzHXClbC0RrrlZbVKfRK0Q0EVbtK5F5vcspbusmW476IKiYVGAjcB
eIaOF8J585AJOHr/yuzuIizKatEDx5L3MmACEUkVF8QyhY3F5WvQ0lrdkwbJSzs+uyPKxc992O15
ZsA9k35bqRRVhw8YMLp6+IDCxc+A7fro8oQ0VWTfX8N5Fob9xk3MSS6z5QajDkTTKFzrz3c9yPnM
iCNDbrgwEz2+pnxsPdnRl/LOGfpMg/Zy/yrNlO0iajAhUEQVD8F8vzeo8qmZ+TBjZjhJlNKFY9ax
k1GUd7cp9vTLKDjj5ECYgW1IG53Aom3Hjbfo3aCnGLYIzZKYZQLP0vK4UkrEiZYjvOh1/HzMcYPB
5bmh+u+DyomwATEwi8zbIM6+SCj+gyeLZN0rQQYRRuUxotnsQXl1Bw9C6ce1QxbugDcIyIyGrXgV
B5Cb0fD4+BKf0z/yMwBDQhFOpZTck+gg2KkAruLqrc03foM4DIZiDsTV8raL50JOVIonNpZ9ZZqp
VSHIt+6ffasHL6GBRuu4wmD22k5xzoFdvTeg8IWrU2Pjds2WzKSm7sTLTZJz4QHSds8b99nay72R
zzrj+6GQ4Tsngec4Iyy34+UkrYdAN6LIOQvzrtWvbU6Mjf1kXzmDq8TAojhSvWvzqvzF5aPptRYz
KHvS+5SNmq+6vGxgUc2BDFOqNE/sDrQbukqNeSS7kSOuqSgvneyRR5LIcCsIpa7C+4UjvppdTwKu
qbcOBaOjY/CTRG5Oe4mgRuq4kOZEqTe4aY/2o9Pi0EXcSkaI6g4MvnrOrgLCXRYVebrS/0YEJb/n
QH/CUMaCVY71wlFDocZdtaW45Ac41T8TYtZRh4m8wDunNdKQCuqKngr1uQbT2zKvqE5NIcREjdNh
9jLMxWT337qCMpG3CGAY63MZbtk/p1Nt0VtSLCFoSXD/TLRIzJromYDFHFUHqWZ0qO7QFLTTVWJK
t7y0FnpSB/GjK7/gancEcBSgB/tqbDqCtEJIR78Md2MoFeUF+R2Z6USx6LQ+2wPMnFiv48pjV/JZ
aZwPX5bMY47KS3xiw6Lt/vjsbN24cXsOx60Xl25/7LfaW8s2tb9idJLzs9YyRLwr19yjXnFfLMS5
wtw3gEhRsBvvchZ2xiIClSiv07/+FduAMbFtqc6M7xq4YJP0byMmd7lFMfcjE9AFpy30ANhcdV1o
Xrg89531VYEUe0fhZ6v0aa7VJTSl4BVtDz+18DAIuBwqofD3sh3kxvk6/FKMkWH4Fi1/5l7Nh7IK
W3dPZixfmQaDTkq+rVgqV7CwE8kEuuPUnoSfY4KeOsxlkVTT9HN1EiPRhls4xKOMsGlq6zAkqtI1
Xpyq+HH0SV/+DD6yuf7DOgJNHv9xlwA3eV1Nqfi4dqhHPUgZgdM3FMj35+qFXa6yhRrTEeXMEEXo
6DeFXGuKbDVpWQoqQKZ4QKs+oww2KvrruqzYjJryVzmpgX5/Hyfkpjsqn10LqjlYKd8d5r0UtYMY
wYSm37AHUzU+8iEFXSy9DNxUYjZjyPw6CGyeMLCZnnBWKuwoZikGxNycZSwnz0FaUZW5UZ5ne+MW
+8BqdW2n2ReqGhufHmR2pjCU1XFsSmv5EyQdedGuiusSVRZSfGaQiOpQ3Vqsl4wOr52yVpSiTWti
wGMO7TN/8yA2yYjfa5kGfiAVmkWPDSEUs5al6cGNEU5Ad+Tyed9Pz41qui/F0hNHLJaEU9gLpJyz
bX2A/9IKCZF+OB2ohLHk8y1AOOXDU7DrEX8K7YjZ6/x+1zf/UBfE7VwoFOPFW6JPHgDO9uaCPqDm
lzW84po+s/iVUTfHywZG6OVJ8D9odmHUPW53qAmEGgQbxQ8OuChb9sWCP12i0o+ilaieio1SabXe
SsFRjSRRJUGtehrCeO8qptljdc/sZFR8qk76tCnnlVyETATP4/nkvt79QvOk8wtnP1CH1q1c8eHx
9BMQQZY8Puw/UI6vueMU4fT3ISxS7DvQ4ZJl59fT+smgrvyaJ89xmQ+7sdxK1J6WGZmaC7R0/Gpa
k7FyP3whp+DnclUQzcQpl+tPHa8TYCRBp7qUlNW0AI+hUzGJK4QKDFAwn7LhWsSegus4NT0JC4t6
lgMxLSp6fmxdhRWKa+ALrh2k1O5euzRo7Fbztvyzqy5pEworfCPy1piFElVGcuqBn26svddhqlvC
7JNdS+aHu+hE5+qpIT0Zu5CP3cgro+9lojY7UVY+OpjJZxk9D6DqJCqu5FMq+fYz3ICpnTLCr435
daZX20+IjXAtcGLqyWX4kCVmAb3SlL+7BZOUNJ20zmo33t2UqbZ35YkpqIRDDytMZlM20pXTVxmR
t/kq9kL93VgCdwh68MzZ4VR8oXpxXf3ziT42mnwJXv/F4pUoejC3rVmgKqSRALCQrn46NFpDP4LC
XRwXsNlSIXIBY1Yf4X0Cygodpcp5WGiMHReUBdigob1zOTImBOREOz2v+TnteI92Me38nKXKBuMi
RIVLc9MGwaJ3LUel2b+OWLAk0VEb3KXPiRqeDvQTlBbf00HIj32I5JttB/k4YF6aBV19kZVvm1dd
tvpdBcocSkybME42VLCTNVOzonXufSp3ceZC7Cmhh6IBthYCrfaU7QUcFk1SvJP1D9DQYT5NwzWt
JwgbdMpOLDo80HIvSv4nGMcaBzJ9h7XfBRS5HOgMKJUuJ1cm15FGalbMF+2ei40xJwmF/Z/IrF8k
J0InQ5KwAmkP6M8D5Bhrbg/F2/JodYaSJVLl6B2mUVttD/g2rMxS45SLUT9NNMS916EZFutEoBuS
+yPod2COQuqzWRkIQnG+/AHCtSTwbYhqTPxr52qaVv5A6hZ0NImo4JM34Gy48VAwrK5sOccjKwJ2
AaYFEaQjaWlZv+9IsgT6yS3kbi786RFY1gWbhHk7dKuogFknR1yXWP/AS5j0P4AqBScjTGEMKHQa
ywLfJ03s3JD/wouY7hUR0npxi7Mn2F8nxk1wBxx1XIriGdgZbRn8N0VJxaG3aBPeEYQxdXtYOxj4
884w/y/ciGllhrJGPn6KJ+WXXfaFdbdskWgTIVlYVljQUAeRRmjuOUha5Iv2uMdghRXbPNv7PyUZ
ijaLuopqN/Je67HDxDaq27FlyK7bav5zz0z2oL2Sj4mTw/9UkqdgsPjcAWj17v8RXP1rs0j7H81k
5w0j/iOVgNAz6w85LritdH7f7rEcTAAZwlWolVJCpYbs12ARTh/hKB5IyQ+DWiNfJmzL2lye86X7
DixFSDpWY5GsVlVvf8mcXve77MjQoLwTIQMYNn2HiXDPcHx+f32SHNnpyzA9KftGfw4Fw1eR1hYM
/RltMqjKyaXHKeBTx+eRN29F/I2hF2vq5TuBO7IGVltjq2RXSYCTySlNvOBMQZBysMzO749CLfPA
497on4SfbR3N9GL6VI/bVJOVXghoZCfY4RCN2ZIIDHHcp2PLvIrn0XmJ+2DaQ26H/ejn1zGhC43s
b3btYqFGN2WNzDv5SFTqLrc05heoTrrAi8ju6p+vRqBsBCaMGKtsQQxHURMxkbjqZuM53lWun9Sa
h/8Mn1nwYL9tl9zvOyATmtt5VergThYD+Hx8z9jFe/+MGXKqncXMveKS33ZERxrNOgbvdSV79Rp9
Kp2GbQiQgR/TkQ1jGq2CL+XW1eUZUpVWrMWHUAIK4qfdWrXjaQCQU4ch1CcWK54NSyBQMkQEYsKY
d1WngN+BMjDf80bdbr83bVWcIWIvLb4ab06DETsTAqd3DwDqBPofgpkXI9VSAM62gr0U5yZw47OL
WQvWXyTkktrqTJJxp8Z5lRMgYP7EORgUW8NKkyUc0Y1DhakU5h8mnZiYIZPuBBHPDbmiTE0uKFfB
+IUpair9TmaJQMGrzyDn14MIHUujwTJxSEA5ccKaifrORXZRSUMvBtfHzjPkZQ8xtdo2wPRaocmQ
fV4s1cZNd888xeK/U747/DJp6e6Z27PZIQE/ksJYwSa1jk5WIqzxEjCC2SdykVY6g2OOMC8JHNmB
W5Y/WbQ+VH4MmZBqmbAik11Ci0aav53mHn+bTvmIon1ZQkAb4qP/dJE2unDZK/e23PQmuX/M6KWj
OsWBBD8o2ub8QqL6s8rBBzl99KCZJYFMGC+fwaX9bvHBOJxA6fgc9Og8zIBDd9l1zr1q9E6OjTUf
hlyhqAKeAL4eT5adLxRYz2UEPlTnFvaVcwtAF0SCxMIY3qE6JElEtr+XABDFbSw5Amouzr31Dgb0
pJeDMIDsXbxO8kbdZHwlxiWqqmtMzkZM+nArw+vAITBm0Xt6p/B5iSEsYwbLeoD8gSTsXGhPt4cK
rpdPzLda0SWNrOKa/DyxfLBZpbT8EvCO6lgznZvOraoygna7QDkYqRv/WqBOyP+LwfZduuUnQZFb
wBDgKiGl08x+UkvtFIq9iLY/6HACn8tf29Hw0yf3PElsILzlIkldgw3Nd5HqtZ3ZigTsGpSOLBlm
QfjO+2awsEnP3sFG8r8acnZtn5eveyBKwUeJD/oYXJK7rONHXQI3HnaoGZsQ3lU489nBSarpgQnV
X4HavZcuR8rhgNpWDQPOylc3mzdTtZYi2Le00NHq1gPiEUIhPjZfrTQN1esV5gcGlX00X9P9VxQb
rdQgJlgC0bUFygwD2XVvZfnp0iXdbipPBD5sT9x/9JsV3wsVZULs7+NkXW3sCzHIsREjeECcbkvX
x03j2G4A2CAcRt0UQLHuy6s0gioqDHRnrjFx0m1CkW025zcHlE0KmM7IIf2QRpAo5QGU+/lydxte
CLS0G/SElMXr4HcYHYgAAqZ4w6vmQFDOOljY5MqKtzQt/o76nneSA9HSf2Qbr10GPFMSiSv3r5q6
IR9SiRgBqYG02ag6grVdgwCtI5WH9yHWGNVS6HAHEX1XFV56D/VkFCMrc5gadVGT00q6qHGMGdo0
9o14n5gsWcOc3WvLKhyRH+TrY4+fYdZzL2y2eHO7PM0HcQVvCEqRQL1h37H9bOr4D+XEYjgd/Nne
6DFVBRsOL2BYbOw2BSHsRQWakdedIV1eoz/LEfJdylOY9WqVQmx4JUQ0PMO2e87HWLcuJjsI0KPc
iZLhG0OIq1VhKQ6q4W0VwH1hSETNQm7EkDNpkpLL4ZsbY1uNjBxDWqYSSmZZWfcK5Fd5DGpuYCIC
GJ2XMvL03VOOcLTAscmHh/q8wuehXkwTfdPUaGB4a3CuXhnMhZFuR2nrlB4tbvDG2IWTah2q8Wf+
in//ZpSaPx5n3zM/bPsLJ5EoxAm9e8UDxtvtdxBJ3sWlpj+mXQU2/NxE0K/oyPjdFRe7S2gtk/F4
FnMht4Hrr1AnWVkGhq2Vx9AlenT8SFGbUqVzx/kjlIYY2IIBcTnsIQchpmjK+wf8Bt4Sed9COAl2
CdxIepA0Ei2WoMRACMIy6zTedz+pn7iM/qzgfQCOtzpBoiLE+f+WndaGbZT1e8BRzojkp+NiXJyE
gANMsSsv4PtCHn1Cwy9bLW5Mht5v/MEo6PfSO1NyEcrddcmyiHtzWOf5JVnkY65PoOsN+IsWc+25
tzwXYYpp1TVeqg9wkZwP1EV2g1UQOpXCqQvUzZGACQVOLIsVhwVbKMfuFaazyAqYoZ3V40BmzhWD
SaUPdI6J9nE5UtoR4dJTq7iuN9PyMq7v/safehMLXZtvSFWi5OkU88JYnP8/5cd9nsAnGjdz0r9s
+V8jSLK8GQ9e5B5l427xaTyiDP0dsJWvdmTcdcz9HiIGt9/pXkx4f9fceQ9nu2cgoZ6o8nX+osW5
t/5DoWvOYd+LHmzk3svVX4S3MNQoTKaZEYR5Cmapq5utogc5oais40ZLIuaZvqlMDKgM3jHUHTkC
PVwIWLNaeDvGktOkIN9CyCre5gaTJgSl+zOmeQAIrAGr9KXUe34SD4Qxm+dniHDzBMJeezAx24VG
dtPP/EDEQaY5t43OUyEz75Er0NxFogBMRqwpP6s09hxHM/v9LqYodUu8zrRnxsAIzh99PFu642YZ
64ZNDMFCX0TqRXZvSiLOsOyZYfIEHHW9eYE04gUMvU/skiWcmHIIFvtm0+RAalAMwCq7dbitzoAs
Z3PUqOz4c7aBH2vYSu0p0kPcIL/VvXcpkMDSh/gAqVDeRcLFqco/j6xPp/E8Xeo1cy/uXyDuQZaJ
ysZ5u5+LtqiumVZw5kjWa1B2xP5yjf77fW+0FXLeQ65lCSeC6FTq9AZ2IJ62gW2fH+1I9nJulaMi
jtdi0RcB5/hFcBkPvWC6o+yKD9lqUJurgi3cUGRY+O8/vhtp4xf63Ziskz1kCFx7APjwf8qH5Yjt
W/Y2Z0bLYJNhfFMsGqQmIeKp+eQhMd/BJy/mvh+jXUKFrGOrWnSztBIypwMDFhP6yBT0/hL7yc/n
bIdUxvay2mOtfwwS7UbaeDLEysXq0pNneEn3mgHFYIt5Cj8R68tynfzKc7Ec0gAwP8SANzgNRXMM
KvZFIh3CQ3KjB+eAnB/wjKV0UY7khzuHnvgmBneM9bgRDmG2J6xFRZy3B8N/dVQStibn44C0tDLu
ltOp6wYV4Mcnf21fI2i6O4+l660Uzikek9z7ezYHWZPoL/+vKcUPEMR+3LbOFy2l8wo3u/NTcxIe
Dp6VQfH/jkOGGCsLJYbiSUIgLAEtdPSA8fIi+2hX0vt+cuOm97J4mv5nLypwkcFYJrrArhPXQBE6
uiquVAd0qgyirR6Jy8RJdPo9Ba6uoUwx8txkSNcVq9hbXgIzqHwyKPY/OQY9Ml49NmD9TvCARZ5Y
YJo/5H/QhsxlPWEXqzwtc+LzvNs2xb+dlrovYdt62+A5Txi9YKI+9vb3K0L5ujg6jaRlAE8mTdF3
0Ou+ISghrAqr08pV0YA0BIWMOLzA4WAnU8xbub71RFrLzh3wwwWBPi+bgbWHsXeLKmicpXfYWc2s
hPM3h85sgnNjpfuzv9wVWBb0r1HyHkoCho0ymmIMTs5UTAQxpDySg7ilo2dizwAd+ASVCSybQF7+
FRjMs3m2vKuCDdgBcEpYnTMNH4ZRl1YNCrkxi3jZO9wTa9D69IFsTAxHhaUaBcyoYdXZrj1j5fXs
YcNk3XpHwlCMPwpH7p5qWHmfnHkgoHvAHjzCSttLKEe7og8OdAcXRuNYGAhuiSHUyMb1jZOkvxFd
32xjmHz7MgWVX6qedAE7d13GUlyk3VwF/tx96csmnFkgetUaSabnQSRy9C5t54OvjGDEDzWsaaN4
+g6K7aX8t8x7p8r5VS0ujvIIz9BzrdNDCybH7SrntSgpRDzphMVxVULuQWyqvV9oHRonIDk9Ly37
PVLSUulqub9CuOKbb92B72YOR17//130glGwAIcfON5uwtINO7RjIOcmULpSTCMfosPzAoZggBBp
uikG4eMti1vPYQQ2q/mGnCPcCUG/BLLQnZO2+krgsOC5Ufcoq5fEtM3HiCTp9kg90yOaDv71tMPi
mArzkMl9GRPJdnQKwcsZNgUjL0kMxoH7GCA1y5dwCKrMCA7YF4dDyiRfxgf20cGK4hS27+LELqcX
1p6eHvjmSf+WTDfIDG2UAZr8HIL3k2U6ATmwEXdpC6n89mIORSjMq3PWxh+RTJtNRtWi/Bte0BRY
0Gcv48ZXjSLp4wE1v2HdBkvjh7HRPlDnoeKMHUB7RHei+mo/0LlqEOHFOROA/zRgsm1BvM6DCi1t
4Fu6o7dFEjVr6CLZbimS3CRdrz3LI8S7LGX0zYWPice9Aywjff2YNoHs0fW8T1WGwi5dK/Snj/mo
XkCYXqFo6Ffkk8M7Z1DD4zH46eV/XDiidWWQFE83290CCHnMklSkZbN4jJHrKoufdLO0prHxbvLI
ceZVN75QQMwPozyNHdCxb9b1OoOdVIb1LWn4HuBE34JEzY1X1LsqU2Q5nh+ffvubr1mBe0sfe0A4
QvVfZvqvYBfZccADZKOB6vpa+UPyZs9A50FmLSgxv6QZM79uMsbXNnXco9hCo8cY4fGEdGZVjNoR
7ceUEmOf0bCGkGBiIKhfKDy53axR8125tt9E8caZEvpvpEfgEwlRcGvK20e4W+z0h5mnyjcdYXHg
pBSRDDH2uX2JrPyxOMTaX+Nyp/7lZ4whr4GMYFlEFvbtOlvugyFUhOoE89J6RWaC4AtWBtKKPcsK
/RQX2AQzsb5Vlyhe0d5ZS96jmsrrSen+ZqGw5biqeaxm+obDKNatOyCxzLwrWDTVnEVTueOq1VzW
QlcvINnZVWxnNGqupg656iJtGO97CvzM8z9l1XLcKi8/FXiccRX6+RB7fRUASrGAuJ6iBS8Na7DK
xgj0YO+2yJzuZEGWBcLQrjTPm1B/vPJKdu7ut5VdYI6xltH+fCogs5J+gSBp73So7OCo+m1paFHB
vHWNTHZvblbLwJwEz5oy61xmH8xrsKh7lNjX+IZnkw5qs1Bd6A8bya9yGYQqE0WOqeUi8xEiY8bJ
OAJBEWyCqxULgjrG98tBX6/Io7HvAA/zcnrQpwcBB/vSSyQyCFfDu24SqZJIvpbxkB3T6/1ZSBf9
EacfMRle1Gwhk6/QdJjxHDREw3mMRoHXUJhaOBy+WEFwur9qceUPb0q/uLJ1kmIgfJwQZ8YR/Z6Y
MCS292dqhGj+7I54Ve1DlW6213fx7HxqgZgxXN4V6k7WynIJiTdgOKmlB/bJO3ogId2xWMQAClUQ
dmE9Yp3oYWYYZmHjhEToTCYxBXWO9BYdr6J54QK7/WSJVO5EfNLnyRZfIR7tc1s/3y9fMl9jJKp8
e95OPxQRXyxu8w+z9CE5D52YgXSVGbyrfJ1Wm1MCFtvSp8+cjSKewSlUGy7QzNVR399g1gROTk8W
TR70Z58+ZtGkfhpT1rqiY6RHpp/p2OhdQg7DRB+hGskbMeFqhV5rOAKYzP7BwWEY1l9UcbcY2frl
7WzPvBqwgjWzKlQRpaGa+vaFr1y9rCochkaMdb76y5AwrG0GBXCqg/XFhhNkuidJvK69BUlQNZs3
RWGtVrL7NKNXeVo5xy3INwuyrxjAtC2Vk0pZV85cHr5G3zS9ewrsv9gD4Db8RwHjQa4kzBgg0+SC
gx2zrVcc19EyQ6nUg2KcUZ095VKDqKpA7gIdntLK6DfjHJCF+plVw2YAG8Y/hxvI8aVvdG4z5I9x
Dwnby8dmt2F1YjtxFuhwwosfV0hmifN8ljecgRcRCEwZ46LzoRokuem1MCtr5tUViagjdqrcTaDw
2sXWkxMOh0lcn2DIwk6L6qdBU8QkVsl8+kwWkPIRi+tMzBTfz6ldVPy2Re9LsmAxvjJQ7Lbp5sjx
mQe+9O/D+BqBKxYK2+wERd5BEHleBoAXRFkOk9MlWitoiG+2qOLcbOwkHcFp/7hkz2Lw9kFSnUzW
PwMDoch+EftENnEP5qR/8mfE+plCV+Lfh7nhRrGoG5YnOILbvbR1899InAQI92q1zLN10gx9yQ90
LpSVsLJ77rVJBySqtLN2ZAfio/T1sYbRuM0GMcPqUYP2wuCmnJZjso+jQJgO7uOzxMiVoFjYDEBi
e6B2qOYi/U+mDwK4TvTi07zQO4pbB8VEzhOp+1lQO/YOmInVIi+5qP5H0dhRkO7Xb6vr7yb6YADm
lqfaUsBRcPPYlmnOQxiJpmvwdbmMG2V5zR2yGENuy8h8wzyj+x+B2SFiOxEAFtk0rOT9GXP1b5hp
P01WqoMVLKxZ5UcakTcystYuWT3mImgxuNzcySthgFC+GzYsgXw1jnz68QoM3f6Ll7Kpfzr8oA9E
7AlSNigtGVLyYm2C+TjMNROuvyySieSreRNCKvA8t5twT0EAi03kWwCHSN4Hn+vGVAhk65HfUu2Y
CsDruwAjOj79OS4ZZYbxhMvZDLvsDNp6FF+O6ttPZj71Q+MfSZgAuHgVtUF3cGj1fHkHoczVFXKi
RXILJkiBUje0pxZfLNMrKgttX+vCeyW7h3kKqCjkaIh1R3vX7sFzJI+HwEE4w7AGffbvkeeEqQqI
RHoDCrOpoqGBbU40Y+uE4ijXpbtQTwQLEtOpj2V6XZJ5+6kIerctCEjaSLNvkTDH7s+NPVFi2rp4
f+FsclrOZZwOhHKn6F8Dw5wqW8GXjenH4XAf84XU/GKviIh8IAKFikS7JYOOo3KdY9v6mM9IW7WR
AfMvA9J1QMM/H/QNpADhmduHonglGIrl7KXgdXBsW887FlsJsm7FPjYA2fZWD459hsweGjDMPFL3
lCzFrgbfPDPN1vy/YWOQJFI6a5nhlVoAgzJpKbic0MDOohDGs3wRMX+rPjokpuWpDWls8J7YStp7
t4Eu0VW23H5wVYotQ3r0Kc6X7iN2ln5jORVumkmiXeMNWd+hqcEObBLpMIjc3F/NMZTs9YGOP0KU
GcaVFPPP3NSzHg8KlfrfEeiwjuoKkfbEyRBYusXHBvrJvS4wLvAgZ50c3apkMJreHy+SC8tYuMBd
tfguLBAy0tOPGYZdYpkyA2DkVdX3vQ9oAHS0pH9K6RwM5o+wSFwKLOrlt7xV9gPiWsCcD64hjuQv
St2+ydkZNZSkMq2LFsiKqwujxMzXeTPK8CynYVxSNg25ZvLRztUMTKoOtX0T/fsMubaal5blVdbz
jS1UU/KF9F1F/Y3ow7Iv23dNvBKccHoiOavfsOMA9n/Sjd0It+KJqUtRjq4PXhdEIOxkxDuWdcpn
mdHpwQCHa/fJDDUQowexnwEz1oVqgoIoueZ6nNMrip4H9ydtjPK1YJH2drBKzCrR1IE2xetgQj19
6uoi+SzE0YNBdM6gcaGLT++G1bUFvdLUBL0KYHLjnrivmZKBaJlyw9uj+Ax877cy/LnDdpQE953l
idhjtN+F+XD3l5vtlN6eo1qMg3HOZ2ObKgGjd11P4YvTHChy3mrcwHMWwW0RQVUi+756iW2Bq2wv
SjkuC35b1zTTJReceHGzDaTm5ddpc1woQnFJZRvfTrE4ETuQ3CPLjB624q1ZWg282xm2I9O1/aik
dL2Y45bcFLpiMz44yu6MlvB62P4S2SFcQdBth8xl6jGN65RvQ/Xqzxa/Y5fpflmHDcUlk8X9Oqnh
D9PDhJnla3K6rJrGf+VVJXVAELwvtRZIkt8qzpQrqSyCogINosbiOAuUv7m6xVImpwt85xWRErCm
QZFvLkvHejSNXu4OAejBU2J5R5WXwy2R8BUTGSLB1qMGlEq4tlFjAupioI3yXfziPobELEeG2eyM
SUhBDSzG+oaJBF2HK6KI1LUlHAzdOjBRwQK9+jDoWtwMxfV00RkOtF+J1KoVJn7icFswMAG0z2un
3N4r4yYgrCsuuvyQ3sQ8asM3xB/4bRlFCY0ZM2FQ2eQpxKUfQLVfQ87KHisE+wUo0IZNhrrajQYz
iBsspjh/RX2zGopZybvaSnlS+sQCzuzY6x6f1LkDRarCBxpCSouSk6B0mJ0LSmGmUUiOpCfs0tIe
FvFC5W1zljuHQPUGSHrgtp7ahGGMcSH6jeaRVEIZDrG9Ab9biSvOjrhJNo4bycMIfQALGGIpwCSt
FTRdqtWFS0LOIN7Rv+GtaWCwO81FK8LbKNEz/ewI/zzIg1NlUMR/eaE0gIqIe88qvjhk683+qRe0
8b9GLhH9K967/r9JYAkonbH80akNo8eLD3BFcNFCpSa7dVAvmRxoAbMHROBJgJWNMeoscA65wPSx
L65SYTIOKLWATW0FkcDopbFgzOsf5cBuW2tECTxge6kjD0Hj9IoMInuqrc2pDl/YJ6elAUbnQHuW
/bXFbAXT2+8edOf5GqcjiinsJRd4NuLQ7i4nd+Oz0kGzputE68NRWyBooHIpod+rLXAI3fVQmJwI
IndOauJLYYFASy9WKoKqtWOHd/4N+cffWyWK78R+wtIK8CgnzB5DT6m+xnmiNyO2c8C/u1zOihx2
Knuumtw5hbEe+phYqJP6qZLfSqV9eSf6EbrwtGxUagQKUp0dUG7HPdvzgZZtpmLT2Taf8QawWmAi
hyvTDAhJUGjBvncuE+/ZW42h91vFN/QDvap9CcW47fxR1rJAghrRwkCI8PBT2VVL19qxsykZPWJx
LA2FivknInBbMNlYWw+Z5aNBCtOP4+MWh6W92hZFH2cEEVCs7h4ggSKOTzUyBzT8zr7VHgBphu9i
3MzsqgWGfk39EpoY+rgFolmqxJ/LQi9IAja/p00Xis0myuf5qFj9f3k7LzcF2KP63jk3+VX4aiVX
lcYQtpVrs7Pj5tS+qKKbnrSIonZxVMFQ5PaY8NHzqnloaRQrIPOgnbL5e47IDmiAURfMnVG6dDGq
AXGN13P4zI+As6fMWlSIVv++wW73zYcpQ+oXZahzzonDoUxaApO5SS1PGNGA2tCjnGZtaPsMbXwu
edugGFEhKFM0JSwXiekyOKosWRO6+rS3ZR87i6eVz95amfvpgLCGUoe648MoBgwosLVMJEN8fBY9
rBmr7HtZHccpXXepknfW98tHKlrECRwgq6+Yxldfx3wHG5rQ5jvLleRkXxU+UTCnMEI0Exy5bhmV
Ekwf8GFebFtmT3VRlZ3BIo9OVFxWhD7L0gI3MSgdCdEy9EXsR1s0PdqsiAN59ib2xPpPm9Fbe/rT
JFtkuAWQJlmPzlJSpj12GCAFo4gF+TEShj+wZg9KDXuVsh0E0s3Mm7mUK/3OBM/RSz5FtNrJrtGl
IZjsr6webY+ICSqEGIH22oAxYiFgzankT5NEnL3yMIzqd/SKFEehPtrDaZF3PorEcdZIiu60jqlV
YjTcDjm17q1Qe/K0xiTIYm57ODnJTivKHZnNg1BO3pjIr0Cm3b1s/s3C2TaV/zF6cVKdogpjVVNq
qlL+q8XrL4iEib21JpwMCbpaJ5pj6b3b4XT0YGrWq4Np0KdT2FJYPJMJtEsPy4SfRcT9mRmNwhgF
Gsx8ixlk8CtPz6AxQqvmvmKsziLmhDv5aWQagoHb8umB0xBesv4FdM5eczD41mSfcZo/ch+c1OC6
KtNvAEyMj8yfM9mO71X9FhHry0COomGKEVEO5/RvOAnAzHhstPmqCDMJRdI7GdDhTs5aUZfGgTcr
Awm59td/wh5es+zmFU6iY9/iOGo4R9tc3VYMAECn77c3hWS1sReQLJe6e7O5sybipny/0bWcHMmw
eBICnse9ijwBrLraZBzrg4c5dLXRSf1Cj/qQmo8kWCyCv8fA5p9TXrYkQuS3s1Optjz9Nwc7CFhf
V9Fwzk68/KsgQ8dyFmr9SL4csACVwZzwf4s5ggFcCPi/Ur+xkZCobyYalMBIg2A8ux2BXFwVxgmV
l2DCQBBupcnmPJMQZu9/H1x9yoMIgYPWBnwuGt6g3Gd4We4I/HIFCBG5joCGW72+HhcpzWgSCt6p
LckrEjiRh4n0EflgzHCn0iJJydR5sVZ30hUeddiPVbrG+o1rD4NDvyqJKtSfOlaX0onpiwHdrxN3
z9nTXTn/Wk9RhhSq0eABela1cdCu9d4GaqHs4nvIjOfZdbxWo0Vp97k6lUY4SrUO9pNXcH+ZECCV
DSkNkAUSPq34TNbFm+54amgCpzF9CCy+U3kZPGCN+kn/WU+QvOtAScNz+HSpWxmmaz3fmi3Fkyq/
f7fwfnpqJ6mwj9yyuI9uqy6lneiOJ3Sd+wuc/vh6x7PXrafsmykr3ofKLAiuk7vidMH8EyDalfIj
q4a0XcJi6ts8lR5TgHS4BE0ZNmqC2gy6BZAetPsHfLzYyJ7wLo6wY2xRBYJHzfxwi/273h8nZdwH
DJXgfE8hk1rAUvV/jcG9LxqI8XKeVnZOIXwVH2Q+6z2vrA5xGl02XSyQznGz/VAFpaMmfsLvR4p5
wxcwD2NyyhalrRLxHKDofH3F6ABnUE3LrEVRlrgpZx3p8dv6u/vzTGftUziNtHgWY63Q7gwkAg02
/SfE+AOBBotonE02LNoKCGUDIf1plZ4gCiMhqeezefr6DtRjiop3mgHvPppdKzlSRFOw/8U4YI9h
oFOOc+XNftHwOaYXoy70t9uI5Ysrost8ZOiSrW5WyjzXC+SvjgFegkXgYP8hXY1m4c3XPy/Ml+xE
eZGhPpjYiAjcIe3wq6GQj2f7PcC1Ynpw2lzQ9voCTfRFU529aCIae9SDaXjlIWP7Kiv87+h5ZgsR
1Mmyxf1gz73HtCmEeOBXsRd1hBZa3ajlKvuu+OEobZDkA/oA4+Yl5aexivFGch65n4DYf07xr3Iw
DG4hv+W5p2JNXhSa9MJneHI+ZNdDphukihHvj8rS5miBbK6pX1aoDAsX8xN82SsC24adM/QFqoWA
9C5L0ZcIDve3r5Rk5EEp9bUYmm+s8SpqO63IUdKa0aBk9csSM+VoCzNDR5OtQw6+WmwB69D0AaO4
0lo0UchPSg0YLauZ6c84ig7/NylzLrLW80ISxRWgt0QWUfsFr+P6TohS5rbz2G11yF9p0EWmf5ow
fQJ3BsCRWjt+zonkg3Px170FeqKOcWbA/JKiAYDp/rZi52aBwvoNBYmi8dbfwTaSUc3hG5N9mL4j
a6P/RG5dc/UujPyp3dhezqROF140jtn3nZ4DpxQ9vMFpIuhxTcCy9YTug5XlMbY861ll/y6X+D8K
1BbX/sHl8pDr9A1HjorEDgfhZfEavxqthsG7T48/72zbO2y/rliHHek65anA1ANALpAqgocA2AIV
8rt4OzSYHTSUxI9pbTApBzRa9tvPiNLLqZOGBqccj50wvAhM7pJe/W7r5eupVU1xGdlWODcYzngS
d/GC2jQfHsYl8sMbX6jlkLMrMyukMCWVd17ToyMQyXE9h5dsFF204YrU0GTX7EVz5yIKgWOZ9Ws9
paAkTIM+KFzNMR4w1/mJIa5ftmrf8w90BmRbWpvLPoQCQNk0w/wXBi2pAuFdUd7MFVHdoa4/izpC
uRszPl4CLiWi9Utom4x+iNxm+YMUySFQWm63IRmG/LphVjFiqezjpt3u1t2ReFrs4XYY3zYn9yWH
AVjhAm4jHbJJ3SP7NklN520R1he0YSzRFtRjEPavxn5WUtS1AuOsdxsJEIYmaM3lRQETe8G1yUrx
EmXcWFvtnArv7XVSEGe2H2Ql2or0EA+fj4B6nGFuGjLdlQp82yTEfIGleqkiC9q44EbnISz2pqqe
bzC7j4Apiiw0eOBLtSyrxF6++rhsk+x/dKmjDcPlXTBYkvMXSBcz7EzdF6y/EP/sohAK8bWIlKOY
kgMr5rqrtqmAw/wMwns0VmCNZOhKUnS1lklLY1d9L2AmeJNlWl0MvvVx4FQAUwDbR/DvkYKm8mes
HuGkiNJljBI3itbiLwyMQ5EHWoOAl1HJcCIScf0gd5pyFwXxvKq04ggEYEkIHpomrPIsxVrV4/Xd
i6lwxKXLdvJ9Sjh2IMFccnZY7ueTEAnnEw4s12LfqR6hBUfOEpoqmfXXTyUkke898fcK1ee3gevx
7x5FIrh9iXVsL6GhURmWYrHn3kupHFoXUCtg3Eu6rwu/BS+5mkKPQUKurQ5HFqENbZBhtARi9Suj
LItXaHjsx0sWidym4dF/AYS+odU6NLk8wH2y6hX7ckK7nHnLw/9yrNWhKHTRhtApnlSwrJY/uqNL
83ZQ2tXvzYndkfgJtO4ldp2E1glks8Vk9jx4fN8rMFJunc6+gMShiMuBSmo4NqHnMlMmkDw4xbod
p4NIbMXAisBw7wL557QMYJaeBJGgFRS9OvVAfC9s6zWgT4dAxcnszYP+XWDvvD3iZ8hEbAvWlNgI
e9IPELkSphbkALBNvjpF6dpYNdzlAvI+uEH+je71CaqVcOjfQBMcSeOEwgxjlky+5TDRZpSZOU2i
G4RJ7cVwdUDf2Q/nG9kDxMASAJuz6MzzMC77ky6wbJ3srljISgb0q+h5YriT1JSL+TF6GwKRKEC3
i4YYfAC67nK2vEb74oUMipHtVRX9ahIJw7taRdhcOqz/4M+Ug1i5XklUvVFTPypFfLtuSNR3hrpQ
srLR4XKXpdiz0p1E0EYfR6uB6zfvg2MUfx6EIp7IXldv0MpJY33fdsHOI4Vhf6W6ffndf9J45yg3
7GVI9bAsa+S6+PPUzquHc72sAkhlIqz6L6V9pRNf8MKFCaKNE+a7SxLb50/F9ikDoStlPGG7Y7QX
K5WKPW5ajQFVUIs8ITxxV+Wt4V0hxolLiqdN9Ychy3VY0CblV3e91h6j93nbfldC0JNi1k9rgwo+
6P4duS0Bl3NvLHmBV4OlqI98Y+0KHTAwHJB/0yllhKeJRQlTY6tQps7M4AV7DqZkGeCJeSvgZzML
PlBcQO4/F8GPdQ5irnvwrE9ieauhkE9hLXPpxl5OtM9zO6ww7luZMuIGk9IMTwdwGf9Bd7wl5hqC
jOPNm+/bM9fB9QksTt2bcOIbKumi3DVLs/wf+XNAoEOr+w5uvZyzo+iT4ExN3eK4dSOC3s6t2Xko
nV5nQDfDKKiCC6RJwB/S/4TSpndBMNTwUqrAgVGFdh9UDnBxmf8m/rImO/MC4aRGmz2s1oD7MdML
ibIRKrnGJwc5w7ZpzgRG1SDaisYErg+moY05+ZPS0eeZdU5hiJp1eeq0Q81Q74agbCMpIPRAeKJ8
6MyYPkmaJCyuJD90ddhjvJTqltGnaNlxsBfzw4vWVBkjgVXV23voAHcHkx90BJUwWxSP2kyQwPJJ
9H4rYjTM1bbuZ3rlPjXrxg6AtCh5b2fzyuB/opvW8hSkk1mTf2vq3jUsxMKnj+wL6zVIO6OBlCVP
qchCSEGGKD6g2sk9/uIZjmwReLkQBCmGJbWXU3XDQccas+/dB7Aoq2FSr5CIWj9IQxhY9HN33zDC
GpjduIP25mqRURyaNhp9z87izYcaJKDbTuJLR6ctWXyo/9JLDcvoHcUulZk4qNUaMQPSEPRp0PwR
RLAMq4aW1MjP8FZGfNpJYcybb7+ufF4kDeYEQ2RtkDSA2ASmQu5IYu4aT9gV1/9CRYzADfk+/+01
PeUsyjPcPwuz0dj7bBGLJRyWWBXto6X+cM6xy9Nj1rkMDT+pDHXFU6boD+8I6AA6e7yOnAaSkzFF
8MWa2IzBYrz2YCdBSUHinETblR9Vb8UVP4dgUyBDcgEeSB29cN9FLiXVEZ4pXk9w/NfNXwxr42F7
nd5rEULW1HhvvnE9yUN5//mZnIKMfTowWWcsdUx3M2fLUn3PYGg+0v91WbKkeG6qK8ZWcqUAtvzW
mhYDXTJeey++SR7dKmQpXl5qRMXCCyd0iG3nIof9vl0rzJ7fTJmD8z9P70zJIxINaD+2d/Qb03kL
Ng/i7YV0bRm63PdBxRO5hfejzFex8q9iexYADRpF9/DQN5Ey9tMDoQP/fqKi7ngoodeUNCApiJ+A
I8ay90TqTSdue+7a4x43k/FWtogl5Zzu9Q1qfdiD+G8Y+LafrCFH4l6DqLLgW/s6+6eMGyZaw+Ua
pdTUesVbfVwhltIOykrVjs6P3elpGrq+DTr39azcS7/iG6edJbzIlT8++G32cD3lQbPGZhNk/dJT
B4uyyCpd64GbdLpPjPetMyMyS2RYeKm6oa1NLT5+WinWlS59bL3neaI0p5Ls4E3SkZgOtCqgQp2F
EypHA5HcL0FP2BkIZ6+23wk0ufHxl2JzXyuSsIghfElofSuPXK1cjITtrQNy7zmuY+hL53tqy5sx
8jygROxj7X1in6UNS3QW+HyOxVMiFqwgzw18+WrHxzmNx3rTLzJA6wdTsSJIO96z1rW72l8nJ8JZ
9/XYhW0hwuKRl26ldWCXBLMIOdHLPZaVGDSvN0PR+TKw0/Zw0YIJ7HjZJB899XIF4ObhMJTQAjwW
EjXjRV/9rAw7HU04onkk+PIi+QPapKUUR48wElreJxFNzZWw/LWi+VIZZnfBAjfO2xZCFQ6dDuR+
ENGy2CWpSvKR/CIcF//ChMyOt5b4XIJIXambvlrO7gRQHODJ0Yhb1TFPI2t9Y4ezsXsJpOu+fGVW
lEfZkd4TjsQyHl2KEIvIdx4hiV55hf4Oo1tnA+INmP2cMSRKVUnijOVkr5jN4J0qCmT6nwPe9VTM
gjUvuyb3ohTtEoFC7A/AekeOGUGZBFcLN0zEfA0HakXBLevfRZSZLiqwR5G6t3qSyuAzxa8nHKId
FIxF6pXJI5OqobpuilDZCPhvZUPqylR+0vcDbtGcB5rT7+NVyCGm9eTJBQXWuIU7Vc6eSxTpr5q9
+acKyNYxed/CK+c6r+5xJuX63rRr3Y9mgKGoOy9azcAplARTvYNSEYGm2wdJXDMnl9poUsQsRAs7
3Uk57PCdo9iP/RY+JqaIgeZZkA/AN7DBK432cucpvjKIWTdRRWWGK2umN+bpLih5IZo7AlPfm4CY
gwWyxqKbaeNoeHdJgwfNvJaz5qhQP/hBRCGLKPvoUCjq6nI4WS3LPYysu+jtKfnVfKBr498pnp9E
LZjB7btTt3qUDKuQdXcYyz9LQjjqd/M8D1p5Ihv/YymoizPLKhFer6dUHbEPkFS+6FB8nqmeb0qP
+mD0GzFlapMe8ymSviOmVrUYxMp96D7tviJhoSFYnjZPSVg9Z9yrzNaIYrRyrT1E0C0C4aU30oS1
CcyoA1RPzkuG6rLFiU4xdnAtWF19Ww8D0ugK+hHQ/BMoSSonPukaNs1W++/9M+61GSWLzWDk3kdM
vMI5erZktwD/xnZL2vuJpwPE0agrcPdBk2Bx4tzIDkftpro6QTgC7gBT1B+0v8f7E7KC1x2ubVcq
JOTB6Wr3GGdb/o3xeroC0XH8/TTy0e8ac6PInRl+3EAPW/tb1ERHIZsLwzXa9fFsM6kbyvrs95Yu
p5o5tE337XCmacIYEuCWcTUUmjibeWMSKi8I2wmBCqn/OWzell02i4RniIszMKjWN5P/wZ4kANwi
nWBR6VAfwUVyO9cyaOGJsizP4+W9DR1SyDWFJSnY6FPe9u88Yqsvfq2YXRlfTLeIoCHl3GXxbwnn
g6Fqi8GK6DHDssKv46RAAUgXZK6KSInPjhX8/dcf4DHRBPC733ok6xh0aooEVXyoFVxkNNvNUfVT
gfcuDD2WL40visem+e8pwhHYUpwvbsK02uIe7IZ5nCbX9seXJvV76fqYondJcrzzrbbW6hdemtFw
aojo581NxiNyKJGDb2suTPCA9ue3J65fuPQ5J2Kv6fhwhXfvsXVlMHOMuNKe57SCPBQ75MKDzG2+
hXzu5ZaTbhRc74bCn287oUNCsP8+Xy8MSNdXI5/LI91PQA+iRgnbdQhnVZXjOb97rMw2mxwlhtRN
DiHwk2JEZZ3SN787zW5dDGWRtuoEVBl7YssgBkJDrYooOGGrViQ+sauneRByzQiJM0BhrHI2Me02
Nbz1usQJf5ReG+fo1XrxeSo1Xv4ihdRQtxJcTRlgAc8RO8Q0YfKz5UMZB9od7n/siJIwMtnVJLDS
+NJRjufMVdRhAEKMelkHuxKzZ/JrEIH9fFRL4A6y2vi3Mwey5N1gCQ6uLBqlexngcPX7iOprrcq7
gHxXz7cSzJ/75Ad40Y4ECpFuIRpTatrwiz1kOCrBK4cS6zjue+sT4I/cQaJ5amrKz77VqxrkByYs
T2pcI/+trvPuFoqkBABtNLQNkn7BzmeYe9jh/6qxV41DYtRhrfF2juynvzqm1Cuk89ludAhIm1ag
D0RLf4dVHag65rb0sWl39yDYltXb705/L9T6seQSPqIU5I8Xb2HqLVkur3NZX1tdqmvoHWQqb5gJ
474eQVUHzBtGmTWM2MzTJZJg6xPT5CNMmUlMUmqqBSq5KYI1vT8Ei3uZuRPQvZNSx3uzOQCSLWLa
zXaFR3Gd0xcu6+vG/42KKDBoeO6ax5FB3iY/I+9zDaOvAdbgMjS3zZWH98/QYfqBh/NofCaV5Mi/
4FGV5b5mXyu6LhuP8o1R3yzQvhnlUHLsQ6omULyhNMbTrTmEnR1xYcBf/+dqPbOnhJQR4zsyw+pD
jqgxe0NJa8jjR34WDWLqmqheQZLByAyBg9RtcNrY0O/CsD+lxSD/FUyBAk820W4AfXg82kn4n8C3
zRiEa6xSVVOyOerCMfxAi+3UxWQDjKQfEi4vubfg7Mk9jdXHJzsP8QxRivyB5K83NHM9eLtZXjiK
u0g6nwSwjtfX/BUOFHy3DU3elXTdDnQ9LXp+2In4L3GanIkCKRxdfJnUPCHeK1wOgeP5ZSL4h3MU
AsrpWdCIv97pRI6i3S/NHjncxBbTLyLz0KA10T4sjgUDUvR2rEs9vTn0A4HJDDFeiDkGG2vBirCM
4MZTFZ6zX+yxNR1m1hW5ILGN77kak8h0odMbj0mLbVUanuDjHwKYECda9OaSb31o/pA05+QSHO59
CZZzdkUgnBxZjifapECcDq8lQq8b9qoAfkJjWcNfrDPr6Cc2TDPyb5cJQyu4cH7vUMsfJOw+tLAM
5NO/Iia+J7lpyCZwfqNnYPUMvCaUdFMq7b7f+8s3wiN5PXu0PJ+WxTPYFR0jW7FiL/07LAaGZ1QS
3gPJUQ20uHUFMJbf324lWHb4Q7L6A7rN+nksz1CfDe/dzZJZDGYY+l0OKSuQKQLSoe2CnF3GlVth
Ey3ak24+P2L/fPd2lUUdXyCQ1drOEHS5qydh/ty9fO0o6k6CFd8LNV07vOU/NEyVJ6VDJph2EEuU
aDWeKtmoeGz0kinzN54UMPF/x3QTlU+jOVhL3DkHck/b/3I/2m2vPo7vTF4uI9tpitIKNRWTi97b
fj5MdiUNtR5+in9kfriMPqGy0+eYxi0TO3BRhila2R3PjBBJixhztnnMa27iHiChlFmH2ZqNGyoh
PVCtNegkIAq3waw8FleA2o3NsAlg10BzOreiFtpoBE+ucAwyjO89APwJMkiVYvEHD+uUGkw9tOum
J0/3mYO2NGRFDxTxtoZ+AOoWzCwISn2y7AbvH/4fprK3MIIA0Rq6C6sCwazmFwIg2d/0bJpwqtwD
UTZdDXhGOKEsCjJP5Q8UtK01ak4u7GLyytXWjoNjVGdvvKSa4mhZOO3UZcMI0YH2N5Wa0lGANock
nB3PFZCNjNa+173FcLE5GGZ82q6fFRa3YjAEsn0IuOoPhN6/UL73ls4N9OAvxcf/o//t3e3ncDX+
kRWljrXEdBQfxK87mJgHMnQvqRgf68/qcECUdUHiKQ1E25FUJZQ++3sNE1PVXhoPTm2/G47ir9bA
md0pdH+me2zbxgj/AkQuL8F4eCej/xuQyksHBV/zhIL86AoAOp3u6fG1gM4ZzSPcRYQy/T6TLmce
pO8dQS7ScdvMKbreGhMZoQQtWYGFQsztQui5qbOs/keFBPW/O01wOFPAfmcXwnnvkA5ZOzmPlMtY
ZTS4Qa4FDXNjMKhR5NPi5Xk5u+x7d+4s8Fu0/dEDbtL+HpCAsFP0tPnyCInbOZ09/Z1csUy4cKyZ
UQ1Q/3Pks0WJvdT/olrOpd39bezDIgr7TqMEB+nV3xWeu/aqe2i8mHYyV/9gpwmbzdD6lxuukBeN
oCRo4do380NDQ3l2YvZ6/AIS2KTQ8rvhMs/EZDgnPvZgKcegkKY2fORQLE9/zCDEGdVdyTCiPF+E
xFJyuC+L2W8NOrIk01wWzQ1qU1PnVJAbP2+foQq1y1vyaXE/+Um6CvCm0LJKbj4U9UcOXAEluN3i
VupguQg8yn6m9e5O4jQ0pW5+gwQyGMHmj0ERBlv2caui9sZeY+CZAIhiem2XiHh1KPKpuCn8I8g1
/gSycadnI0T/YCx0z/jbJZ44IaUEneR5uenyawLObubMXKDk8TyL3wpAzRqNboYkD+LPsFIUqtFe
3vgff3+TN3LSs91Pvz3TXHPwWqZJ/sg7jQkc/ZLgDWONrHp8z0bSZLHDzQZSMEmOXzRDCyBrNw6Z
N6DQyurWK09rDzC5Hofcg7YFWSlGmRAY0uCx1iQk0zioyZZigs7wYg91NVgcRHCWMJzZ/bctlUll
giGM39ZbdW3na9B2KvSBfs7i65gr6g4/t8OVSxDfOkfiiJYNheIZzWuhPrk8uA2Xw6lMJcGU256r
4nv+En99vlccsf3GeCvYcQM8GM4CzeGy86qK+LcmKepgrnQAQ9E54NEtH8SShqOQp/mG1XSC60fU
8YVLzaYb0fcwEBEFRHUpSSUnWv6JvvcG97tE7ZpqMuCa2nJAqsRL+IW3GXWeDkXuYDMsX+XCi5l0
7avYHIeaowfIQpIJTrNWnSNenrLt4wZOwTtECY0wMvXh7zrhiH2bSTwc29rMO0lYOLAXcQokI49+
PmKkejVnFigdnoA0RUFJjyQYn5COi3BACncisT4+EJm752w7QbqtImQQxXyNSLRck9YZ3rscoH9O
DixZgORzmGizDA0Q/AQ/f7wgs4AWBfT3ZGLA+ZVXaL0Zse0w/nj/8RrQRiZ9MXV3briLK/F20ATa
m9KAVliPyRKkB25XrJ36RfZ8bgT1rpiG8OTF0zWpBWyDp4AiCBC8yUJxskSy7yWStyJyX5DGZBTA
N6ZZxUpCJ0sS3kpgyMKpX5EljtAWY1l+ob5UYRE72f3MAHq6EwlNQBs+jD11yXf0D7g9ryfKE44/
2uA1fxH6SxvIesZ4f8ETCT/5vErKggnWL2HEOW9BBBkJWF+t8FCXcltCQrKsRg9s2wBlKaVfGUic
R1sP541vqjsAFU8ovssxZqEF+4ku9iS80iD2wpEU8dBr4INgWpYwg8WI1+WwMQpaRAEOByLr2Krz
DQww9Y+CK8jO5pKZOgkQK0vNdargeyLbh/qu31zMkf2G6S1/y/0MYBZolZ2o5sA+eS7YZLWbf2J0
S1JJN+nq3evs1c0CJQ+FHd55MfpzYVNfyEJ57LObE3Hcv8Ril3fZoTUtGQUKo4p+k7LNBAi/5OLf
tHwt4KxZwwYlu9r9imhQWrwpukidPsVWHbgNuMVwykIoe3KV6TETWCooZnCFia1NE04euyu2EtW3
p3EPtICzZa8veVm991JH279WchuU8GQO+qJ+UM5KMBTlZTxJ2m+R86sljIeormsldUYn4Xtkuw1Z
ZtoFy//Sx2l23iQ+buY9Acwta0Jbq0NLbG7pduyol5b/pxfhw4rjioaodk5betZPCtI6VwdKmvOo
GtM3Vx48qurbsspk0pN2L4sIUFRmZ4BURPpHXbKZlxtu49jHGHrEgK06Sin1t4QYNlCs1GwEf5lV
duFoQrjiIg9Z05tHanB7iGxVxqP4wJNh27RMd8XSGCGqpn0KGn0ykAizhmrHtdib+YqN9N2uPiai
Ji4ttmCj7SNmyL3zQ5SL7fw6y3NKBQcS9NWhb3KMTD6iA50MwqJt9tgOTAscBr4G9k55NoJiSj8Q
3dLhLgyi8QTu/qg/MkdIyLG7ZKYvPIyDOw0KM98qyv+qOIx3UcdXozWIf+IqlAt48QQxtg53oOwe
iOwH5+0sE+JSfL4crUSl2ibVm2jy6c5Y6YJ4yi0svgEsrO8LTFYObANKUFOyBXSJAH0+yfg7nP2l
sIbwhhbfp9v28WjTTbp7Y3ApTDV0Wc2b/r3mCy/LATC7A+14Op5DIvD7VZgjImDiuCBgBtlZNFmT
giIRxP5O15H0ETE0RaYEfqR2FvVSohaTRumSGM5Gvuhx1GMmXrU+f4mv6+jBw8T613dvyB3SGQKT
Fhjk6V52KNCixKujbk8FivlcaKhMYgbdsqz6ZygJBZX1nOYAIyKaK0ZNU9Au1zI1ls/OXLTk6Z+b
KbaTfU3dywi81zKt1gVdDymPETgvwl5Cm3hQMQ3tzIxLKduqp6dhKBFc1ao4kC59JKwheA+rZR4o
HYrNJ548UWnzv6S9ypqEWaQwwlfJrdiEu5uX5u3MtCmDq2ymroGEqm9tNjWqvvk4WGv3mJ7SUlSI
yqnoZgcmvJIUUk5plYBHAQKXd6UMsdNhUzZoRTK3NOUB8IU1VvwwNshnkuU/A6LHf0VCuLCrcWIz
YpskHtVcAah8GxeMh1IuRu6ma0HXUNDmapMwoNAz1pxDGA+jcSetkeQowtzbPu6bImr0yVPxUhTp
yRSrPkYvBs12zMiIm83xxvpFnHwVL+siL1Bm0mels4XpvRPtuE7V5ThDB0JLWBa8yAn/esd7HVFJ
61jhzzbr+MxGc+aC7/rnlIJI2S6seA0kYHHdQrADyQxO3QEyjZ/g+KU0RNFP6ePHj62lfjh4xbkd
VUAlarx28DGB83Nk7xGNcqIISlyNTJQLhgJGXi6/997101w5U1blMzJEzeNJjitqX4yJprGqyPFC
Rvt8Wh09o8zn+ATmo689kuHaYBpgICnJAaQ+TQ2LeTMa7RTVSmx84SN/Sg36ZmlVX5yciWL0ELfa
nlHFVJq0xgC0sqHl0SuDO1Ff0u5jcUTaeiLPHYPCKPm6RmHCHKmYVbXCef0NraYDv0M2Jp/9ptkF
GWO2iHUo7Vvg31IxaKyVaFH/bj6YgMUZGoO8m8ga6krv/Yw7JYlz1+YUFO20Amx+O13L53MnqM2O
IFP23/Kvmz5mkGQb145hGg4UDwHXM6/vWolcJfxua/79y4kqqMmK11GZqBQiQbcwzDcg80U3OOlv
WTlWWCiAR5kbp8zXxgKesmc2dbyf23zEoOst6rf9QSqsYlCtCA/BZS5gex3LfGW9Cd4wS7YTMf8F
vfyN2iiCG5gnIZswCm97mNFGirqgM8ciokNK01NH1GvFmtG0BISxlqdBCyI6BtcckK6k/RBUCrct
R8wyRm/tAT143zvYy27Bqp3ZxwqFNapzGlAdNK2u90fy+3Uds8WMX97z084g5FH1K+UEt99Djvsa
4jxwC+hIHu+bfAolfkm1fM6Z0U88KlCB/OFe4+RbfsMqItJnAQ/35DOY2SWSRHBsGXyz/ZfpZgSY
Epa+ttUcr/iarHHv9VVX86qFcnei6MTgZzazd/rJtrLOg2Jyj8fnLHZKiUyi3taO/r7VSyypNvRJ
BiA02OXi1UKfYWrT85zmJqvEfusifHj42uZsleNRsDpX1JXdNFXA8tF8AoONAP+j3s3ab4SJBLUz
v0tD86HiMhNGrb8Sdj35EvzIP1zk314UFHOHLRR/YlHvTDNW/AbCtPZzF0KTQhmqyujsPn2CBRk5
JZ8jAXZ7mhQcDlTnw6Kat/p1LeocK86XOmb/MElQfQrhR9js/XR8ZQsKMNTgsJ4JvgGrfZLEEyCG
dnm29owy8UWNgOKhcQBu5r63hGrUG66R8YJAO4jad+IHarBSpdn6oAVo46Qpg9RDhutMA/Ef5T+F
lGHhlWLG9Zb4gxTwblZVDdU5lL4g1k+7M4DsLHswua/fMsA83lio7TeqyKZduhjLbPGcaU7ORvCk
h29fqtVBQH0+VHn3K3UDJAbmfMFG6Uox2Ek6lGTOAzViGs6uaDeatC31Tia65lTOYPX0qjlCN8VR
Bsb1Zw+nHiYJ1xFsX25WMD5G+5g18sAIIISiG4qdHQgvq4aotLIm/BSWbfAI7nyan3020FWbil82
EsZ7eIGf0Hwj4ArEyeFXvfxitqfYhOsfX9g1Deh5sVHnrd9Ku2D5PyPxDDLF+GUq1LX10GrZRsi8
Tnb1hb5K+3kCUhth3js9nU7b75nGTOFrh3Wrjok3O6X7yRyP6OlfMwI/mndusivhJ0IXPxWvQp3b
Mn5VIKEXEOgBrttfFCYRD42Q2gvI1jc8WpHc3YpqL62JfmbJYxVyShj9oekWi7e4tzTaEjS31TZk
DjSjnbsYeJSCPpRXA8d+AXe8QTBw6wvyZyiXGBJXa6Is4Q/+uxroJOQRGpAOCu5LSV4V9ouVce9p
M3UkTsPdsEjK8MXNO5iS0L6LcISXYxa9E66mRN4dLfDrXBJJ3Ya42nOvsUPcRQMShWooRx3DRYvO
5N9zhi/J8FBRgE0pWWgDb3MVrOaMxCN+XrzVm5hrGLQakTEzoRFVHXHRr/8g3VPB6snG6hXln17x
+aIuP3FQ3F/HbVvw7kEDtGPdH9EDQ614cDTD6YP01TtcmAvQmLYtkupugw0taSvDNsS1hoydODPS
83VOiGOIzsvXag1Tw0UfF1GvVwyIvpmOmGkjek7dn31TT2RaoH6KTSh0MiZQ8CUezuiXfXIK3Y8s
dLH69qncz93E614vH1TbFqeGck4rL2FBC8b2iqeHGZ5siFb4LG469Y5/17XcY6uiTgD6Kj7GPogv
3rnH0nr/AspOqMrV5rADuVg8Y0ldl8Ergui57FmpStpehT2k6OJmxhyyduavZWExeobFkHgeEwC+
AAER9yIylKLlDcigUCyCVyD0s3N41+7TMWPMquulrg40pitdB5J8hwCrbDnrT+rioQ8IhfJ2hayT
kFrKmbSUqPUZIM4zwGr+fCxTbPjpIw/kC4UGgAiOX2pSotB+ZpY8+GcZJI9R84ImxGdMux/r8MpG
A1QNQj/OuT5j6jf9YdbQ7XT9hjDxYzgbwhpZY703ESp0SEMo8NNWi2NwcRHe1PpAR03AhDAqs3xy
P5IWWJ1XW7dk7MWVMcbvxgMaJMzCFsgW1HrFUlXgnXPnKR5NzAIPGx1yKrmyXdgRBVAB4ATThY7i
637j81pvdx1QUlxPZG/p88TUWwTvictwCeNJ4zkLwV6GySdG31KHwjsIrU0EYt3rxGSvF2kkmt8E
w1t2EWiS1q4sPFJqL3Nz0cd2FD4qtnhZzzPNoVFD/GjnE6jtsfSsYZhd1aMY6kkx3/cW5Fb4JHn8
ucmyIA6r1OntW4l9MiH0sQsVMFwbeAsBYlxYAdKnz88NSKoNSJcYxWc9zU/3JDXauDXdwNOicBF2
m4EWPHInjMl0vTp2NaHeDHAPZl30QNvOTkTRluIQbnBiSglI0/3UcapMcOzwmPzwByj8nE70acc8
m/MYp/R5pDDIQ3ddfNyQTKjGjiWtKH1RTUI+KxeiA+PakCrmFD6GpSYzz5YIfyy/Lh18IW8Qchh7
tX7Za/b7k67/nngwL6HYYTRwsnqqhiKKRVJWsEpuP+5ymtAj82q41uVW8RQivyPU7SX7yWr8FHq3
xhjVmxVZw7zJ8FMP9b6jEDmxS4EsYAzf9oQ0NENk3o+r+3sIM77IwUmL3EHLDBVB6gjXv8WpMnX/
oJlvSNnw8RZuOidRFUSlCK3hxpUemA0Xui+NTArEIJwAnRR0S+jSXjHz+LtejAiRKR3Sun8KslZm
6DxtGECib601XYyKbPv6jP7aIvR+Rp3KShM6vIEgJLY1Ve4QrEahjlqQKeDAvjoDuXsFPP5pmhDT
JFxgJ6mr+4IT3lJAZZsHW8gNKyNaipZDTcRtAPMCBZtwJmTI+M3v9qy1j/U7zyszhWSnwZD5ecD6
5QcNcsRlF1nlreTMWawGdksdPwiAEX9vXR0MGgsAzBz3L3CjB3gASktSQo+gchQrikpyJgNkNfj/
/2d23eKn4QOHmUQ2PL57Z4ULQzs3rzuXDGjtE2/+Fa6Ukfs7LUb5GTmMlw1O8xD0XYJZCawdWMfw
1hBncHTeOglx7CSZ3/y1VVFvRsbuWG8rgTEzJARaA0OUqZ7/Bv3EgSB/GdChz7acLJkUnN79Bk7s
MVmA/3WBSRsKHN/3OZziLJLyHiKBIwMqgwzmaoBY5JJ8mUn1qsmIu3BatxdFqv3c6XwRR6aLaPCF
VtxEI2BJ/fKoyDrDRxVXTNGgnI+qyijkNnOw1F9GTnGlzunMkkGBJo0Bmspgp0kw/xnG0HLEaHbP
bU4oZgciWsKgLvrwcJbUpJgVFG9c0bt3WLPC8su6QwKiel9nYeCiXsKllCJwPA9FZRYlABuZiAaR
e81NPUcH37+BeWXNKAjMcQPy/6eb5KXfZka/fv4KZG2ewZSO3Y0n+EtmYGlb0iprq4sDYK2i10c6
PMo7vJ4Z7uDzyoRwwWG7zNNOTo1UlQ/12CAUcZANKbPidsQJhxE7gJd+6I6C5q1mOa6Ihu41RPE0
OCJk3CPShiDpB/7gW5tZrJSYjLAjVns9C9cIqyH6DkeE5Eu5zIpLN2/MXG1+LUOcaD+2LUeC2VQr
BGibprwjGDMPaxc0co1rzx1T4awp0A24uQFs8SUsNP67/aARiNAA8YiPGRaAzUiUWorFeW+PKvTS
Jz9VuBlnWtCD0oqBiWV9mUJwgkYE8MCPxH7v3BnR0OByZi0WmLwKdwt4YZxAl8ZavFqohWjb9NR9
H4SeUFgn4AveZb7rpg4H3GKx+odug9i2VS2qyxpltbHnoCHN+bKNOd9P2v/hNI+otOT8NE1kD5xb
vw35k+1AMlIPZGdXoF/uLJPbZc+88jsjW6w5+EH2Q7rjTsh6uOrgRAnDJKrqZaoh7vJxQYVyokvh
U8eQZtfZ8zrEqQ6fIxmcgnD/DRTqwmQc5rp1ai1Os8jU88tDeF7tIu2Qcg2UaRVHybmkBO8lBBtP
LV41W3E2zJmO/3eJN8xB5fiNue9q6fCLs2RQpH92odFQJYhHHUwJ1uwA/xSxvET8V4EPh2TKPzB3
wVEbmVdEftKF+Z4salV16t2IeWcboNgiWy/jC8kxeHHZqLbsxNIbilT1Hjpr13v7nPAAt77FGegG
9JdkWow9vUhbbqXsVja/jxDDPDy2ZUHGw3iPGeyGOTGHE0Ah6qYIeWkhD5RsYygsQBpmC6cxdI2j
pu+DcEgsC4f+wz5BmUeDE3uEJ1OyqPFe1dPG5LZFaiWLvPQ7ZEAYwmVVqtOp3nFkkKeNnRHiNykD
jN+mNqDVL08f3zp+EaK+hWgib7yBjLggqrsrIw1GqcwmAHtOgODOn+LKzubNZKgvQ00Mtos1O/XU
/i4i65GVvytRsZ7DIocbrQ7U9i/oL70BZFVMmAH0uhjFAcmVjl3AyBhtFOwvGRq+7EixxpDf7vRn
iffX2NS8py+NGAOLXuh1hKuoCO+TD6mmOTacnfNZz7pzt7ALXxbH/QOwin8O5JwO2C31gw7o+cGl
DzspyWtew9sxqkg3b1/8A96msUOF6eJhvDgz1HJXnDpGGVc6eT7EFsuE7xAB8oyOa3gS/UKl5rqm
2sWEAoBundyLvR0VlklxHGFaICyGSqXNcZpVFLd/Q2jgOR1WLTqmvvJoWRtPwlJHU9VORq4wg16w
5nUtfx9xmtVlk+vnRvldyhRmxkgpM1DKo1P3/qsUSlx3kCS353km2Jhasnex9mZLFUgjJFMi+3RH
CgDZ86zwewPPXHSkklub8zDUnCm0oHpOsIzU1PWJCQRoDa11tesSno2CWqWdEcMYJxVmu/cXjKHz
bcPA/HXmyTzPsVlM9MS8XpQOaxJs7OSE6MO93+TXycKpTTEIJW9vVvY9XwtkETMvtUvC+rb3+Ng+
lrTMWr352sS0dPZZBNS0fXKMImkjgo2a/DWuDXMiM3a5429zEZBLrYt+hBSi67j7g/x4PSOMtw8Q
4mufd8cDiqkdNCT9iVQwdD5S8SjLR6mXFBafPkWtL4GOVS6RMBphylteY3a9pXyWw2ClG7nRtAds
+tS/5yd9lz80HnjenYEPdl98EX4Rt7LZNRAgOLYSsA0y/V8K5luGvmg3CcUlK8eh6POc9QNckSQ3
2bam3noBP4JL6Ky/mEVjan9E6oRhi4plCYnHBeUZnU0K6gklLfJcNomkM9C3iUUez1uUHKHz4Cv6
PGij6wfC3Gul34/T/yLDAdmjxMXvRvSnE2hsf4j3ksvDl5UCn2qJ7oKgaSZrIzCi8DBG6OWFdIQ4
J2/ofiM7zuF0GVvE4KsOSzN2JhgpWEjpNGB/O5jrDp+78M+ogW2dXImvmbph8EfCFID2Kr9MWPYw
77841vm8edOwCJbCs8AqdB3V3VaWOCN1HiwrQI/HxDp4pXOwxa9nUhPoYD/5G7apRhXmxscqgMIL
amJOuKenPJ4NCVwa71o4r6D5K25vC85XKd+LA28uri0L77hHgBIiv0RcMKPraz0IlHNNnI52xv+H
sCCBrR3OXTaeB1xXQDXOlRcrlYEq8qJgENiHrzlOjcJEX45c9l4p7xwx25BJ1vRr/uJ1KkeSYZ4b
OMvBm43ijpLzZKVb/ovtkwATdTW1j10Xzr336812wMnaeCyArApWPiqOqTTbWvOuCyealkgRBKvb
rPE52Zfe32yN69UTPweCGcpFVFJnNlzhYDZAXCcbjkP/GojrvsQsQiGWZ4CY8zMwJiTjJpQUoI+H
1uOk345CM3w8iUchWhvK2zTMInfz+Q5nla2KMx+/a1HqUgPiYSswt/5FYptaPvwFBRmFHUxoXvVv
s0AziPKWt4Cynsi9UbV28iOfKbjIYOc9Vr+dAJmQX+iAtsl06JgadAkxmi6/JkpveyrCo1+wMyAq
2TpQOZ+33e2XlVLWmwXe2x25UcH071kcOTCiB1MVmKmetlnkAQYljxZ5pMbmadXDVXc3hzZp/Lbp
IykHxtwF3TqBdmBF1rkaGwnbl8+9RPmH6rFK1kOZ8gDr12NVX5Yg9z4Kcl0+sH2NdVeBmafs2KAM
fuv3lNED3vAnvH/nAbJOzsGrYlow6tw60LXXSGzC0V/MELHa4yxEW4YERdy/7CZoMf8HCwhJNUH2
mHz9m9tNxo987ggNMbI8QnxNDn1VSbuBLT2ub8UQYsyCfQ9ong0mXM8pnenH/mh3iW99AUcyXtNM
18SfR/lv3SQIT5ro+4/qy4AcE4aMymZ5Y6NvoI3QypvDkLYVtgHxEpiQ5G0MK5SeTZS0za036pAd
tM+h3IBqcB6wYxWz8IBaYaQk0jFoQKTHui5s71xokbueIred/Dxrw+qUy1vkkUyXK78xcSCxcnKv
5l1w5VBSJsKYo7taioxAjTEI0M10ZKCXHMr4MpGMX7RP3AY7JDSHppkovSpbvd75/AEcehGi9lEJ
ld4kUcGx1CBUI2BEu8ogv69UA+GRqhvmosOgycfDbSg4oRSsd2xU0y5p/cCODWVTAN2xpjA5b9i1
R0IaBl+z2G/aO296hiMwkW+9CA9EWPIQmUaAspPOiEOs/dWsvYKCYR9C7kfBEBh9gbP4HFRkbMws
nVurawFQBsw3eHOOyvFW5+ycRxSyReMWDRn9siox8sm4Z188H6EVC0NcwIAWoPDS6zYwORD0KiEs
YAGSvZkXQz4QFfmemjlHzXLTDXOVD05QrURc1HjpnQdGhhZKRv6DATKngjvWI47Q/9kiH4RBZium
ISJTpvQJlUWj2khNqichtuFTGqWQnzFBSncwkrR3TT2hcrkbBH50bVefNr9XefvKAaeJjiwest0+
TKu+KWLoPjwemVoZrImxxQhcUSuyXqIUUyIp7Yx3qqbSehsCF3fgWWl3J0iWNAmrZcDOPEUjt8U5
BpLdEA3L1vPBRuNqAFLtvTdQzCxdq24cKQlJIYk8Qt5uAlAfcZWqpALqhAGR0bPC2BQx4qB/z0Kb
ELvlaJQD6KbbhlErNfLLkCEVREk8TFvT28ooMcZxZbrIQ4e3CdY4ZPVtvZLd5jRnfccThUHCaf+I
KE09INiRT74L7MnCDeuoElprDbhutC0ohUTGbD7a4XnEq1O2f/acbF9o3hVL+q+uad2/e6BR657v
NvXxZR5IhnTyrGqK0VemsVUbR17PDkZx9IX/IflsJGNqp3ZUYWnSIRopIZlS84PAXo03sQpvlhoC
gkVCQ42N5D+tFdg/Ip4+CPbv2p54ty+T47LUxtldlMj23mmxILSVEOXBjNFAEztTw8PVNmrDktp+
pjh1ES/Sg9XKeq8KEkw7QWownSZFwz5D7u9jSTnVncHwkZSai9xL2d2KfPlWeuAViDM+a7ogaziz
/DXjoc3X0+sVemmcvMMpzD8bzt2ihs92SWwvxxkpur8901CHHiq4Dmfh5C/F919dA73r2LPow4tC
8srzlORajczAP0NgdD96AtvkEgA5gDx+xideW5mHvhFhhRbgG5ZURzejutspXAHwhIlTumGT2b6h
Lz0UK8OSRbqZWmizFJPgjQbUAulVs8tvL6cvtEidzb0/d7xRnDugV+b2aY9Zn0RVKCLKWf9wVK2H
rUJ91pip028p/NHr0qAxpYWmL/Sy++L5Usw4L8a5+qxpk/pPq5C8DRxOGdRB3NsXXIqvIPznNXNh
VvL6UjWeBXaAZun+nHDO3Cj2jAtYRnahiFiR3B3JOjgnsAAV07DSSRJUki2bDA2Wo1fSiERIgC7l
fKpyL8AFaYUtNNlJCXrx2UGKSmD3KktH0couYQY593B//C1jkfhKG8S6HQ6qB4R6PceWwHFtE3C4
utMwWP0i8JK6/XRyMJyfyouAau2toK9pxglUzwDG0OF/0yd54u4tqGsqSS6adngQouHztwOkLSst
AVqi4dx6Fp8VsitmG6sVAcjJUitAU+eDVQDe8KbDwShe4ivp7XjssMo3nQOTgAkSlYVo7wK2M7T9
i9kX8ERVNUGe/RsfcvNljkJVJyKvtSrUmwPwOBDymmroCY5J5TuXmdsUNDnVzSp5gnge+GKghc9B
PnLUWLete0w6ehSmN58PttCxL+4a6nUxMWXq+RXyslVcPMeKT6JY1/f7DJKyLMauVAq0gjnWuZUJ
QV7HdhZy3UasPspa0mzc6Vs4HNHwYmdfiI73TRNUApxoGt4OzMmvBeIhAK+6VI4er4YyoDemrV3E
w11nZxRabpqL+vGYHJpXRbhGupo7LmFPhEdIpMYHz2fkQ2KJrzN1vIYBoMUgValKCK4dqKCR54MA
nTk3X1zQO1PHxrmIGKwML4FLxROzLOpsO4S7K7NlO+bmMbK/VhhgKZjKpI3liJcFWHaQHExGSw3Z
velgB4zPP0HC1TuZ1NaZtLEII2y2+qBvxfxxK2JGccoXYmfBldjpKTxZvMHMPEwIK7dcCtIxo8IX
hGa+5+K8BHNqbtOgGGm9eCe+YqLcWoIScJawjNShNLH2gsPPxVvzrHoHR8/TAEP/jzdv4an321eX
ehpjfo622MaYkvRgI0E5gwJdXXG/xZck4g/0XzUx18vI8gdZvnjqoeG5DWlj7xXmIHzprYp7a6an
7xRDjVtDRrsMfjzIk2Ds1tRyl9AQK34WOVI/megNx0yDGPcAiMPNZmGkZ66i15A8/PoLxDkFPi6w
dlllUBV49ecyFZpMu77JlPWJcub2ZdnOZMqQo4zoSsE6+O6BrFeJ00Api/XO7IFQGOGkF0Mabqe3
IMn+9hHaktRUMhLv3h/HQGKyxBTiyuxyJCVT7/SIL2h2othh3QAO1b3IKrlCyKISsgc9OJwDVe54
wY3U0L60irAK4+e9c2dw9DQ60otCOM+4l9kw+Gd+qixv3KmumEZw5CIQZ/FFYIr2DH6vUldEKKHh
weYJjqrVBMZIUl+kukmdynGM5OwO7JUFzRHj8iHgsSl5Ca11vuEKL2i+rnHH9fKoT5QmerV7SH4S
PSUx8eW/UfHuagI77nh7Y9D+WYFfsopDDGBnsKXpnvPCq0bAZKDuIdxzx7C4bh57stItKMTv2oF2
HT512e7532D1NGemZtY/vvFCetZxpnbEqeuusR97umo3jkVm85AHmUm7iRan0flTi5pVZQq219lc
eoBCTVJ0kKiVf8f1XwSn/Nz1QmrJpQh1Cq05ZR+a93DEAF2vVhJJhy7Kh9NlAw0aKcDHKaSkR2iR
dxdejMytzaqvT2oL2OgwaPMygH8RsM1gxCFRlhYV9eauyO4xkRtLXPAfn4F43mAkDpmcDbq6dEkw
YbsiILtc9bdksxbWfGWNOWJ+PW5xKb/Iu9J/fvVbicrFetbFrGj/AxXsXiEDcmFXBo4uh847AJF+
eKo24hAKckdtDjcU+docNuNdaAk30atqeLyBP7Afv41nJFl558OEGZeluqRxC/l/6M+YTv0M5koL
4+X2A/Lu4h4zTnGuO5SyVfZinPW+9JWLeqULboBddQXB16SJYetaNP6e7UtN8w+FgakwzzcaE2Lg
CVhir0OvTlKrrk85WxdFGAcAJNsKcrx9ZDamhi4VuqND8AV6h8TPUR6YIQ580m4+LDmcQo0vh54g
UEONn/BhLrLtGHhBoPF526JpXJ2ThS55Z6uIbZJnzH7v4ZxDaN8n6vval3sA3D9QRd+SZr8ZBEIs
Uy4rnVXCoI+P7ejR+2zogc+kKbIz9lQ0KNd4TYeCShiRtxV6QXpDyA6XwNbPHAvV3nb+RrwdADXo
NAexKdWOyJjZN/BDg8b14oG1WeYiFmdWCvNQMp/0NGgXm0BKnQRG0IVw+krCiD45AJ0p97zb+AH2
wnOBPM76po+rpJ0snjvzhAeLP4LWZeaBi6pntEZsRGPqWGm6kNd97XPvUVtzGv4Ko/rWS5Rm4uuP
Wg+s7z2PAW4/k4FpYyc22ldtQwPgokQBH3ggsRCJ6KFNhW9ga+GaMsKMJ/8WQGspjd8mImkkQhbV
Zyab8gwPsXHHQbCotXi2Zk0hiBOKCJ3NY8Zv7TPSCORURwOpkLUdh0L84V9ohA/NCHYdnfevgxTT
leOnpt9H3jsyDn467wIJlCdXpNss35qyTQJl9EExrdigv0vVeh9Ze9qBxLJ8lZUrQDCFx4UbWfkR
jK15OzJAwi2gre+FGKBt94k8JqtHlpnVdbaNPuT7DSbI6+1zrVFZD5AISPCNsT0GWbBmUiqKlOxG
/nF20mdytOYswYM0pussWtHPiIdnPFVe9qQsNTiMKrRa9f+NmSbOHSdp7V7CoSELs8kIkkCef+Tp
zytOcnKu6luOGmL8Z9R5aaiWTfAKYkHzZMytpaJ+QQwb/aauEKsD4lSdUrHHJnP3koHs0pM6b5Ut
tyOSzQo/7QaODXAdO0UyC7Lwcak1pimflEiPNDGj1JFpuBFDsiQAG67bJmzIUTUVzqP7QDkfEvp5
dFgu8j8cmOICXfiwtKy70Fo+bj8+A9LB9lcosUSMV9Yu5mARuskMRCWrEx1bVS7Nacrf/Hx5Pxnz
gCy4SetIxo8lOIrxTH+8WgH76lS2tp1dPRWHcZE9qlUjo3cv6QPSeN+GEbGmKoiMABeQ7k9X1GY0
i1kpAh+SNgtDdrUZ5sX1dBzvOSPL8RKvN6mZ+mVoeNo0MWuTbn5LAVAUwtMBhwgZoWqna5IPialO
Tet69PA0r+uITXVHTVs5iiF3TAKEf9Fso5Awz5uii7zRqdiycNHkHFUZWL4N3MIs3Vh8MnKJ3VB/
cMwA+Ad6sn8LJjR87IGcRF2ZIfs+WsfDs3RafJFDOfqXQX3KwiDwNWDhdQyeWXPw11ifmWfm1mgd
+bVAIYucDO9pYKyxaYgsLi/OKXrtDGMa6flHCMjPHpasd9HU/zAZBGroiVYPga4rsNEUS85dxDqK
g/EZ3Hukkw5cUw8JQ/Wc7eRmkkl7wkqZgK2U1JrEqXLFP40MwKj9hpWzgRG5bHPvQ1QIUx9KKFjr
MS4HNlFdpTfScd+7lvv+HnjsRtMM9VtJcaw2KN5bQJMRRBJC4lpI6hR/bfw2jKLBlOPywMpuhZm5
IxHnqhgMUzjA0RHw6ao9JDRCUO7thdoNUURnMEXXHUVRcqK2E+q8s3iyyiqiaPzBCnCzVW2wfQT5
QCl23V525+qCb+akBVE8fpFNmj9tBAAPhdY6gMi6L5D5oI633z09bHkdQMekKVsfevG7FAJn+W+r
izk3a94Vi8CT/RS0nZQKqcqp/sRX48opjpNOYfA3Obk4mopny3qAiKRa0y4ze8vDa1mMm0rACfuU
nG9JD+WxQap0a4fdVb7kOb6AcVZEpWy3og0uvINF88CoJs/Gj/1GmNO9A2bv+W0NKGMNfWeM1k2T
D6WfW2/x6f2Abqfffh4X2NU0P+svdChUukcvIhWnvcdvKbeXNqo/OvU43dz82u10jcbBvPB0DZJf
jeIUvoUmpQufVpusdeXit2Nl80DiYUuZcnKFTnhBY5l8VCxwSIU+EX6x0EN+Y4lWidcC5TORVfXL
QJMw83U+761P4qJQ+nvSSG7NRjqtqZwp7e5vpBe6Hsn8/oBqApr17Kv6CUTF7eG/Wv4OBo4poroG
HUeG6f+wIemHY222SZFIbH3iCOHSgAsUdxdlMJe0znxbRn25h4d0bfkTCyE/tnpR6R3JnLFoEcnu
APiQ7RsDdDqu3A+DyNMR1LL+LwVr0lopeNg3/eiWmkrxNRFQroWzYiGR+M9yYOJIUr0jibxnUkoT
z70MgTDJXXv505qKb1xnFZumaQIDPNKvMLaSzweqT1v0YQp65WnS10vABabCK8wKCqDkgDv8/agn
CfFpGa9Aa25s1TgdOcI8ypyFxbwwsVIpUuP5LNLqhp1IQcnEW7agZvbYdff4MCQbfGUhpZYtH6P2
GfCVhsL8Wx4VKh+PU7WUJH78i7MIaA8pFBs9ZD6aIS32r0LagAqld0nNuBVtl4LaFpkakahgh2F8
J2l40NXpL079mPx6OP1zRlZHsyoCcORySZfB8UmRi5eCgvHgxzHRFXsmFopcVnoeSkQXslNB/Q4r
aE2z2j1ISREiM5diBCbSQGHyxZEKTdKUAd3P/o5RIdYKU92inldpgfRUD71izjwkVlsePt8FJ+Us
hsrIJEep5RpFPq6dDoFQbzHU/R95Ka583t6eYut/EdNDV1Rz1SzJr9BG2sLRp5z+jkQgx5TTbyid
K9uEx1nA5OpGCBPfnFhVg0xFgS3Bs+/FYKtOQbF9sQWFT6Y1+k4/H3gXUuon3ruHJJnwpZjvjPnQ
aEcvQQn89PokxdEUjb6ngHxLG7eHSZyi2SK7b70Qc75QSwDNzIrOz+BsKJHxT2NDDhT9HZaQ0Vsy
6mGzVB1gqYHDhvv6WzbwzWEzI7VjjJ0IOXJ9oRe5rXu/iBGbwiwJNoUmzKc0zu3eIHTySYp6/GyX
ca6N2bqeU+Q5GxGn8CgwsdqLc1Jzxj0GZsJnVq86jCvvuPXxhDWGDkZTMHLE+QrU8+4rTJGO3vv2
tKq7twsyRtayW0fb6pKXi5yt5mru5OxRi4Av6ZBszr8+ChGGQyzlJRuuE/GtRDlWWEPmwR91bHas
bE0DDZoydvFnwPnAqm4t77ZSdcsjM9mA+PVuxbWKFrfEn7kuITzBPVGTYzjZbQ2ttsM5hLX7FxER
yRCT9YCsJDMGUY2inzC8Q+W8F2SsbJ2dqZWcqGIGx3XjqSXS1Vgkjr59S/8V+if8Jr0Piq7H+qlo
z4VqLy0vaseGafqgKv1KZ0no9/fJxxu9i0IHPNFGoYRTu/cqcr2aZsCZHpOJ6h4GezCYNi056x5G
TlB4U4RTFwpmr7D1Dii7pYLiPqSjvzE+7L6dI/NMmlcvLBMkwTCwVdpUhuTVr6mFaKEPOpAAj/wU
4ZiahrCkOEOLiEuF0CDdDt6aJxxRnfRKbSK0xx2M3y5EzF9+hUH56HHmyLl3HMPoz3xBLv13IVUX
igk7S0bAu9Etecd2RLEUT5R6QaFNmm58O913AMMhz8xkA24TQmcI51ruH6BIzh+GejRal/WTdtIT
ksVl/UDPwOzKRdNEGov8FRkh3lX7NgZvMPaTRSegnbEnwR4dakq5mBiJGfX/asZJHooiv0BLaDTc
CR8oY6jkWNUqkQKXEdjuhZWFPTYnCcxDAR3oCBDrSDpJeFuCnivGZXAwV+ZhhpF00XChGA6App25
ZIeWymQLoNji+TgNhZzuBkTJuSJ9u1yk+4kZWmamj641YGl9mIFnjqle/gM+5eiCs7Ju08clo9Y6
ur4Qy0C6R/MNC1aB4aJKvOwg7QbFHqISvLssll11VzPron9W3qO1niA2kE5XLU1PxgEpmx5Eqlt+
ePTI0utmtT6FLeIOZ1WOaBBqJ/Xp0uNvtuT1pVS/YXu+T3oi3obVFcVJ+ITXV+sJoegzFcwXZs92
5jy2ProtgO5c6XEGeuwHWW4nXi7yiFb3SDapotzxSLEVW9hg89lb1nK+KeorEH+QAOuhVMqsNyLy
3cadONL6Nhy9yqkWPMcE4bHEGBX/yyAATPclrsEGIXFwtpR3PG+udzrsbY2FOEBV4/Hb31alNJ/s
aCZY0DJMvHgEnstDJEBS7gkc557FGPQ2y1w6AyODznWbCXSA7NhX++IN+XgYNI20AWVEjaZSy9Tu
UGtK1g==
`protect end_protected

