

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
qYvaWTl2dVn1UYauUm5HneGLdmTNfKYL2CALcG7YBWzuKWoXlk0Id+l1oLffyjtPstUkcnB5XMcQ
6NZs7JK9Og==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
QYtaB7bKNbwxVddRWt78CWZ0keZknIQG6IQKSIZ5COH+hNdpgy+tCPVsEHq4IVZzTG1P1o7hP4Vk
F8E4xV3B+P4d4XumR2TMQt1O3p//18K5GFLVc+tXegTNm7nDlHWB2EseJW3Comce24tPY9JdBxY3
PqZ0pdNcJu1q3elLkyk=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
dcPEPRyvFmW4PpA4iDmUUiTH0W6w8Tp3x24VnlLzTcuDsG/S9IG3GcyE78eNrT/x0pAgwHhrMrSY
yZo9WE5CUIc2230lFJdjwqsu1GfylgdJvImjNnSRTPzlw78/vxcWd8GQIKrHyFhACpS0FlCWX80u
ir6wyey6yythPFMR7YL9alngEab5jqlcDLLq05xFb5xa60ZtUm6H8H/kSZM2WCTQ/2EYo9aRaoyP
YNJgznw4M4JlCmjNGCsEEMbnrUH5XC2MOkUpPSJ6HpAPhZTjHtmrQy0MjGpBzDrrGJZmxlIzL7x1
7fFFHCW51Ue16QvPlxZlJr0kCC3nTtDv9f7xsw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
zhiiGh6iqBtYa8uvzkWpAts7vZ/x1/EV8yeLKnAXP52susoGuPOfmWMYojIG7BJlvNdJsqMcu4aO
YgpCERsfm5E2WNcFxUppU1uIOa+cnCBSZ6N5aebRGghJrQL1tUzWpRnQ2slMJ8Q+gRbsoc3N0qtc
A+A1dAH+z+hdTGoZBRY=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
lbE1QAVb48OwhlUCQuKav8khO5ghQAvoWa4EGI1wknY/PAoHSz/mN+mHHLZytFcumXquM7gAj5vW
FkPYXzAy7xSUZBC0WEUc0yo4Xa33jDRDxY7cxGlzHmyb1RsXl0duhVMcX5rDmM/+KiXLbAmtS7n6
pXv5Z5tj4x3AoNn90rxrYgdqN+pxQ1GZhPZPFZggV3JHWj2LJUr0U/7aGlgZSQCcdWV2V8ktlt4l
b9BA5BfHfgn1UuvjTl44uqXII+j7cWg72Zy7D/yYZ92M5Y7nPBoBrEiv0PrxnHLMrIv8+jN76TPm
TMiyhLNg8NAb1xNexvBsDmGJWQnxf5cukp8uDw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 60368)
`protect data_block
InVzAV4vt+YnKM6WiJapm4KnRrTJeK+HQOtv84c/1uykbXvui8cxnj606vpVtGZkX7ckYn8M7F4j
1UybsXzW5pYPJ1lRu9O4iEcWDXoAbp7oSTb9ict1vBs6X3Tx1y3B9mzsrSordjKiPPoqPmkVE9JD
zw488UQSvA68JqclEQs4NZy1iHldkg3SjQ9Z8KpqfSsiUYql7uZKMIzsInZIQNEpa25538oRf9pv
hIsJvzXHN+fAA0hWBMSUpsUW6u6D2oDoX2AoQvtiSVonvFzDhJUWDulWrEnb/ZZzdiCNN4KjLWpx
xNrXiBlFI91dXhQF4wJQ8e8nIGX72dEw4VYeyxRcWZxQE5PjkalHIyRyYmAIelWb2O1q3gqa5KD+
ZWA/ONTyCpNqr/uPx/HTnaRH9ppYFAwjcgTal+VkXHv17igyq88msKsJ5y6zwO9Ii2pt712eSq0W
rlTnmTWlhEGysZTdRoptYNVthcqzB5bfEToWt60GyqN4fqQpvK+zFrqZQFVJvVeI3GG/JLxp9AMU
Z/2M0puJIfcVk/A1Yvc2klXg6r8XdBaFwEqCac9BA8eoxdGgQ55cT91UtBlQbluV2o5lONhTHQur
JVs43Z0r+kaJcEEl3VxapP3UedCl7H/xluJNSssSV6O9YtKvV75OdxT0TaUGpT0KWoShwaIIO6JK
kucvRASH6HcNEBh3KRT3QOeo3q7F8y8w9wfzo1SjxIUiTKuAsMNvP/vtcSUoQvM14bv97aUZ3ZMZ
EBdP+xI/oEwGvgKTweJs6gRidKVM0pxsCC3iWKgWWhA/Jp+woT5xbt8BWb3nXPVa9W/Z2sfaqlcE
rF/qDfzFpUIs5aJm+/+JySlpDBLHGpJaDPCNgjVkoYNQFtQqvperDKETB3NfI9p+899ita+DIBn7
wUd5kA2GnxE0ZJ5Wi3M0HLgy9LGwGScYFaz4POJCtahUF5POP66DHGIGqyUZfOQk1He8y7rRTNe+
B76TE//NDaOcxmyvGGp/yaP+amKy4oXEvSTBExODusE6KfYXaBZkpt/v8geDYTqr8NDfGtMtpGrQ
sBDvVLsGeFE8CIRydgE2LVpWTY+H/h9J05ma6AEvSKX04kWZHCD+rd08R73JvjIX8P8L0dsPpRVF
XN9OpcyNh/d6xdxcYgNk4maUXVa2wzyMPl18Na2yGxc49+ntNzFs9WI0sWmlBqHlJrggcXfC/FkL
QRzSkUElGjLB/0ppmllQMiGpJ4IPhcZWHVKenL6upuGw7Bqxx4eD/bVW+h/eroPTMLy31qalb8Sy
LG9kwkpLyOGufxhCdX5B46EjjSPup+e9a8+wTYACkpQaORA2+mzHltTVhz6Wwe+sypnyg7dETc3J
o4GRikVKYDhrE9qNr7D1S1Kf7eItbRtWj2EbgX+owk2CAFy/3Fda37SaYBWu3p9F2wd1V/1DwmHK
ZXwj+4xpQ02BWpN4n40JWab4yB9caXgx8dYJIrVFUKQvH8ii3ZlBWYUV4INf1CnE687/L1JQcv3L
gB/00CEQ7XPC6/6eH4RXMkHyIZKDpCNu4LVwccsmCe3fLFU9FboWcj1F+3PDKcMX0r/xhdgFo/JK
dPHW6PwbrVyDM7yNOjbioQhpqmhiYcsMXIECePqzzh6OdlTIqafLx+kQvb6B1ZC6Shyqq47aGXdc
ktfnguYPfU8rziW4KiiICZpLbLwHJ6JqHCma/r0cnsIjEl6N3unw9VOPbH9Xq2l4chKkcNwuSs3y
RQ3g0vy7c56p+cCMapESsI9Cp9QyfBhbwtKNNToIUg+puCGH9xAyWCP0DHQfHaOVF9f/F7eISYDz
7ZnNWifyiao/zBuThgZcxeeNfwNk3ZlT+5M+qucovFt3Ui6ZKrLRUiW/U8V6woVoEtYbtBoAPfsU
voTeX5RPAkIRfmEy1asi0J8wX6OXdFvC0+N17ELwfjK8SjCtFXhybkEF4Shtdqy9pz2aMokdnxlN
9pYjRSE6Yr/hKLXGsH0Fi2x+LbyvaqMdcpbLOQlAbGGkXjpbwoNo+RB+1om1qkolzH8ZK9e5lJca
333DZNaUVZ4kwLXgUjrBuQW6oaBKsdF42QfszzXImgrxtDWkCOQIq7Xa/6A7Qv5gav10GXACVMsj
AAlYYqPEffnCk2fO1kiCQ0VeVsFOE2iHQUmmwBzNOCvEuTNZwgJNn25R4uIEzJu353Uef/UbVde9
wxETkykbovMIk80w425GeP0s6OE98mJmF+xYBW6ykA1B7se/I+X4l7bUGa62qbwH2XQkFVPLWDpT
H4RcW6bRkXnqqaVpamGeOvKexQbBH589rd8zzxnvAS8yIzrXppu2Wb5ZJ5WMb9B4tt8nm6KklGQS
/90hO6mcBotgCXQxidEbS56qQD1UdzC5mmjr5GF7Tfi0mx8yVcYtNDcUfDAUCd4KYMAYt2L+AfJk
u2S6vIeAFSSaTODKNp8df0xo18DaKqKKR4Y2nYv+npCAIYlgbDwtY8Kqngk8OrK1aYrjQDshc2ig
1KcE0TTJYnqA5vBDAbb4XcTEdYBhZ6ZOSH5T2cTWM+7fCut5Odhs5xRWWeCpgjGdSShu+mU4plJT
51nNH9DyNawhbI7ptzAc2HnZQSZ5co2i5k7s/ky21HuUB3D83+CLq5c8U/a+cFOKMgeew5DfDY/A
iDZXKmdgr3jtk1Qqsmv/h6XlvtJRT2Mdm9a0ktKUCJcg+M3dqGQlythaIPQlsTFn0JvHQL2PNlpq
661HNUb8HbOyV1cQm64bvtFVo53RDlzZ9xzGVdq/LxWnGOnynqDdr1TJdr/JJ1I4zJWzVQPOcy1D
o47U6ndMSxBvOJNVLl4GrKh+qpdTEgcTQEwq6LN73hiuBvuF7GgTknuNAfjxaIk+BhgA7e4W1+l1
jw1kGmokvFX1UpA+lJBXisFs0MpaEhco1Ef61hDcibk02c6cEdtT1qKHEfk0GlRjB89nNVf/aWUL
CRN3vh3RRjSD/MQeH/h6Fn4ism4RrSs96A65j6nCgnyrPgyD1wS+g61f+VhLqcktLYcPvVjnMS7o
o7rQ5T8WVsVn/VzxNxLO56RdjLRfALhHAmyzO2q7/jZooGb1EWbio2TQTPuDuSGTc6MOIPv5nmjS
M6kEzhfRnPUN4a88oIkv+1UqHrNu/b3L7IkE//pngn86cF6XtrmupZ250h4hg9tIKCRM4hSjO0/C
VPuLLTxDrj9g7LUwVFJEk8cJKDLVjZEe7dQr9ju1PX5ZoLEjm5iwVBldmwZz2Aw4kwVnQutgAeyV
CaOQJHvAhyujT3WPp9FZc3pG/lx7A07RCSybmSQfHRcW/RPZGN2jdqqJ0SWbz6XPFZgMdy+GDDdz
KQreh+Ofqyoj1cqDDrEjkeRr6jNGsQX8rBN2xAfDPBq+dbiO35vK4/kaBgmwwbetL+FC1znQ847/
4TkKznoaEz+IpaRW2Pq84pTHLxF5BjMRKO7zEpE/Ma5dERHkAtDrgqHY4rozkXhrnpXjHq034DEM
SkpcO4VUPGzo5DmIpr/rBmsIqSxwX55CX6DMYBjGALT9VI+tMPPqIPbQRSe5mN/5lOmnx4pEmVGB
1ZgBfiKi8G0+d0qGGsDh+sjIBXg5FS6bSIGqW5MzG209X6ebViFsRNTHT9R7ctvVKUYrJuqSUkbC
vUEE7WQI3KABMVIyWNGGozx0WSaRfG3DLAGwtrByJFfNrXCSucjfv1QXRmlt3oNoqy/xztqpn3P6
sSLNQhfpPmKfqlLhoCNxiU1PboduEXXdOAavf8zIJx/yRN8Hxu/rBpnfrBN2WIc/Y28IGtvOaogY
36GfdvFPWLAiCjzpS/Pn7nzr6T6fJ7kKbqCAo4Dc///zwrtcA0SlGa/UxLLfedlzDfzp8IiydqL3
DH5bLvt8ZgCyRTiDSmlpva4RRJLHmZweZkeWmW0UF8HTAE6TKsweOm0WJi6Y6RqLudWCh1SDpCQn
d284W0iSE51rul4PH/YvQgByjccvWdMje5JUJ0CXLiKwQvcrbEA+OX48avPmJcwhECMviljuME+j
i7MB/tq8UNQzqBB1B4LeRSFw6HZSk/MNQUzw5aYOTtRDaUKX9LX8E0/tQYWJbg6AA9Itq79cgdFj
bmhT51jekn3ZQuq/4M62HIlJ7J8TMNO8cAs5NbVLczoNnotIgeIAK+90OmTlBCRLfXpnQf4C+Igz
JlZckv5gqMlTkTkdbj+iDmQR8Q/WVFBh48HKb1R1ElCnSQXpX+P3ZvEM2m1qOI0GkcnfLWkmf/a/
gNVQN1RuUKlv2CSmE/zxZEcgvRb4gGQUTvfG4x1J2z+RoxWI/BLpkPDx0AdsVjpYDET33FWt64yl
ubnQOlRtcHvFrwBfpGJBarxMcei6APR13+V6EGX/LYnmJ9IGMbc2vH4C7Jq3Ry18s/6VznG8GjRz
oDoIJqBPq1moUJ4X4gG1+h6eBdrhZj1o+sM1TdqdEci0h7w3utXcRPEPR/MyWrH0GXvOrgHkKExt
RZ/ouZdaPMNl54PVSWNJ3poab3l0lEiB2J8/wokSzpFPbuAhynsio60CWqi0Qfzc/mmOlm8RNaPq
H7gw8SDl/+IyaQLvJa2DacJ3dcMOymBugDVBcpxplmvQcsojkWnurHPLhT14cuEWM5lLlp38Xfvl
ut/s8GLIrdgEzGOIHgY0Wt53BA56aTyzTxVQHPz+NSvEq4YjOjYAE+M25ST3U8lgSwrMuQiP7z+j
YKl3GyHNDmcIx/DYefSBZ+M2jtXnvFeqTFih0EWnFkynxRewxFygVhIFqXHcJLKbIaxXwjd37QOU
ZBS3D5eSg+shAj6G8bf5NJdIEppPwxNeh8TgQinaEIdgPoRwf3OdP/Rccb+XTRh2p6/2qneSM0/v
grfkMCxeTJ4oB+cRpjwGwHGy4k0lrvB0ZzOSzLpIAC/rO0HhFXxOWxN2o6loW8TZSPJX6Vr/jo0F
HxGNiI8Io4r62i/8j9iCxHKu2QsXcoCiSFHJJbp8RCTYBhJQR0/FDBbX8+GXDGs4jGPVkH7foAcs
NQF2o82A9hghyPJo+QYpyUePeQpf1ZNyblbE3wKlH5LZgUG2MckrxiDHgqpteeK1m3fet+lGutAg
9FCntL4wdqlGD7bw9lEczxstYpzfgTmSivUkfKvgzKvNm8BdeRx2+n0XNcOvj9d4hjVGXnOYu6rs
vIqHX0q34kIxk5pZHm/gVvRQljn+qkpc77xT2LmUOHKHNhThhPG8qQWgvx1g2L5THoylcQ9fCG70
3n4GUP6LsfIzYMuTEyo9ayieRAaxget19OmnhIKjAF70bhApPjsaN/gYXJhXw33dQ9Eba59EvCKq
ExKU4qtNGp81NBk6F4ujKHnwJI1V97TGIfzVJAfQqPOvvn5Igb96KApiTSzgpXO+j5i5dMQ7Bp4/
ht2n9paZ6v+omSfxxiELX3YN1CuP1rQfdY/Qy+WfEjGbn9wXhd7lJGk654pJPtCzAx5SVkxTf5V4
rc19DKpSHe9YZcmDrdUuSpiyfso+BB50RRI3oDLtEHrbM28ZLK83fc/FgXvyWyX+K9T3Xs83sMvN
2gL8VM6mXOHSQGni5/nMYHs8ikietEb0W6xuBJHb1ZhgWgLcF9+2YwsiuA17VMyRo1VUufaBWV6z
YTkvP22oWcCdwUnSKWqTLa+++s/qEdXpmNSYbm+M4LHfB+XVljm6k5j5JBSYzt8s65xctnjfFaaA
DCIj3dUmecsfNCS+3P2gv15MntKOPbVptXC3dZL8mjC6NQHbIZeLh1Llw3mnG4hTdXLI3Nl3oloB
Yh7GydreadxhqTI5OmvMjCDE4XSwcoczdCl1QYnVbFgDzXYOR5szl2Jm/gl4Js0+EeUt3tWBYtne
CpPQeYif99ZCLDE8V4sE4xm0iXC5gd7/yattAO/PoCzFPeW0thgt9G5T4HypCNuhH4K42nGfwFYB
nJIjRF6FVjl/PA+Knn0j1QvlQE13CHFfq3lw/BoX7n0ii0Y0HYoPc/ZHmK92KTjjwrBTHnckS3r9
hs7QtfdKGUeX6/PeZ4sYG9FzJgjjMxjTpBdsWzuS9GM+z/FIGlQbkkez4wgL/Jq9ildPBieq+hd6
II3Tyh6qhxG5Dxhc67ZmAVO5keu8pDFf1by2P0J/cwQ93SO+j2N4cNvp7EEYDgDTx5xIR4Mpa6Wi
5GdyK3q0YhFsnnLj1EDmN19GWemMxGKi9LF3mIwSvkYW4z1seKJAstYcDYODyp8eyqk048AnlOn6
+xGAKNrCs+h6U5Trzp/csZqeed4sS61Z//wwIj2uKdIGZjrVYBvIA+EXgoJM2Xtfo9yhg50EYrRe
R+6lEnPZyANIxfr6QXAe3snwdkF+hLhGHKfPpY1HqIB+s1G1AUi6eNChF7evhCld9dnLP5qLT5et
6gLUIK2X0v1W+cOsBVcaZXYJX54N11PYYMg33unLUnfk2dBQ00+GcBZ0wY8WVRf0vFkMwMcw69v9
nwwvhVYOX2tL3wExlgMbY8lYUBcemLb5vMvHt/3nF30M4d7mMOJr8yKeKeFGF41yUlIzLl++w8vU
FY+9whUDKbVKCCre69ZkT8/w4G4wKfy0SxP/zeg+dxevS4y0PyL6oaw2KQq+Vxqp9f+eBM4BPqT0
WQIAswQqLM+XSAT0xck3DZdZYnvJ6xdEetI5Mr2a5p2wFu2Jip9Hermvo4WKakaym3CnInD1SXs2
gzEMdWNdRa7Jyls8rWlBj0j5rjlbCspJvEU53k0k+lf+iu7KLv3o6vyr66zr9dv5lYpqXCq9Phjn
YYsMkLBWRbDlZnVQYnBRkCCGI1tCEk55EU1dEGDKQlOCABNTCB21NDKTKz5bDh49OhnRAIOdsnfO
/mSwLdONDFshGkmbj5sypSsrQdilI+olMbmYMBlHTTDeCfPZ8K/y9uSH0N1M/OrLxQqU6+Es69zm
5GRXb47Gr/QAmRi9lxF2MmCIrpRXwMqTWFtyzuSuTL35ie95fUJzl/Gd5NHY+4CFw7vvjXw2KqH9
uAp2B94kLVkzS2Zikz+nqwc09n7K8sP1LXoKXQrrkuijPZWKKLmcINpky8m3GzFPpBXlhvOMrYqZ
oAgqWzNKdO2H09i+ms7PzW39ie7utXhO6W2lexlguiSo4P6PntjtXYCkpruLmqZExXMJ0HcErUBJ
R8hFBhd5ef7KVFYYGcx5NBWnOwo8XtzIYyotP0CTjMIZub/EDW0gYnq/gzhv/HxoPeKTX0yxhj54
UpbhOawcKYirfvQWB5Rj4RyLZrtfrQ8kM4liB6hYE8A/u0riTllRW0apCvbjFsQDtFxxzWaszo0l
jQt6paDtpLl77nsuyModCmnmPvvTq6X9KxjKcb+VAr6cfDentTdCc7jRABSWrVfFuNLWK66JIV9Z
M3Qd7XzYV430CSS3KmCsWpFYjOdP/fvx0dcbeEvGGUC/jftfqU9RU40jy2gjBr1T+jY82Bhv1eNk
/N2bHldQtKu+E+WfNg1mSl2ZQPkTdXpfpv5jW3pvIbxtEx5kuSxp4HFqtj4U+xGu+vUrRDmRbKvB
USMZgqTvtdRPq3X0vRobpdjZyhl4AqsKvNoFSBe5bLnZH5nEYFqflV0Y15LYb6PQd6wP0zCPbo4T
lXSAoYau8qWcHOZk6rrLoOk1YFCcMUQowy/MIhFBFez958bvHhbsKsONmoAUc4OuVGUdZMWKXwqw
pTmdK3PzUXzlngKZGZQg+wIjYq1cj/5DBQcVD89L/H6XbNPYKJyY8VU8LjfZ4b0Mc2MGeWYOiTbc
wJgkjAixRFmLVOdxDu42Ae9IUYg1IJJzgseIHabRbPdUK7Z2o2jlNzllqpa7J9Qxpxn9rVrcY+2W
V0kO4iTvqggvvdwnM3O7ohnMnKC2fBXtwGmJGxnPRFlmreD4aY/Y0Qa6HPeLzOwHBLo2YGJH/MDY
4sVbDTYNYg1qUzq6U04UVoopx5KdwhHj3NuUOpB7N7serm7dH5/57/GqreDGILkTjRk/HoP/tFjB
3zVBRTvPW4MuDK8j+beXi1NOFSpGta5xI1PF/Hx5orkGaZSAlCCYmO39NHRFnzVAbUGSZ9z0n+Jz
D+iSfMlVrVcJtfgTZQSPWk2sxJDScwmvUQgJ/VRJBZYFXCgV+tMW/bbjYq85KiCiaEM53Y5fZ4Sj
do6d4oGsujrHJSacvQSoZKHn32BzpcGnhxo66tw1DOE6RMYu/MZ+eUCZ4UTPuJ25f3A04dyNakOe
QMDgmh6Lv2pSAgdMoLhwf9pFGkUlXJTrX71Txj9+mXU3EE5seUsXJBipNV2a+qjLcPJB65b02Jq3
9GQIvZRF3TWBa0GYO0UnaPHmakD7gkbfCo7iGuW1VlDoPPrSl9przRdTY3VjSgJQdqQ+1nmSBbE7
/236KiOleWPF9jVI+R5U/yMCUC8Pg7bFt7BOKEC0VX21Iz4yHvEnNepXuDIThBvXBNK6recDwmc0
KQeSeSJXsfaJr5I/fZH7Ha7muVYIjachdcDGXJ5Sl2MZPnR7lBu1/fiz4pXXVWigNU0hPj1rT2LV
ryJJ8EElqTuuaKPCJzfiLfSdXMqnMj6GkSaBEsvb2Fqq7AoFwv+treVDHF4XcNLygL7vDTSKRvOQ
VodfmCefqYWoMN9lPsvKjcDX8+HiPdKmWWpHMB62Hov4424cJ29URkYyHznjPam+lE8i/F2tlEcY
XgLh5TupbX+GMjVXyf45ybdCu074cfiaiw9LVyPR1TyRjw3gheGo/jfw+VsU30kTTmmGN2TU21Mk
gHrwBdx8hwYTVQTnB7vWIk5HX+p95nuT9X/KYh4usom/w5Fsut+IQBiMkFGI5FjRLgDmdMFUrzEV
4YF2rwXp+4CpXT7Zui3ed/VeAzSFU6BgBAxD8MLUkhAN17pjbDu17w8KU/NgWW0JRTW3Z5Svp89A
7hhWsrnlKntwudF2GkpiKt0KzF1s8krb1TiZfR/p37t0PszuUH7SVr4PIaIL05R9cNTaIBrmh9xY
UzN7II9i/G9wLsfe/ioXu2zCVdTdpLHyhn3uKhioPpYb5YeBayx5FaALFvqBkJ9RJIp59tL62hLk
wevQ3mAM/rL9MGQdiDjzHsWJd3P4KrBrMtMB6T0FGXZ0F8gwBlRYi3TO7bBz3pnG26ctKmY8T58h
rmQxtPPS+2OgCxWW5qRzxIQHHFetFBR6LmydxzIb+MCQSY19SAIhUkEUThcGaeWEMz1EVoNQeYVP
ToH2GvlwCqRrCkZFmjShcNmau44i/K60E4WvtLjCdrSgKL30reCP9vkKbedF4B3wP5vJc8n9GDLI
tVd32UQcJO73DzpRNHccOBbm78FhGg3qD+TEE+d7P7uUv2xbUek6nOAu3zvRT37jxPk/iVSgNp02
fXaxqlbl/Fqk9Id2OkZS9m77OEZu1YJJ4Y1iO3Ax/MfBZfAXrySnRtMyIvWf/hWpCe7/6qWdTInh
041uObDbuf2SZMRCosVLBC17BIH0S/kkA+hKqADR70osKxZxUXxJgcMC/ltR5H9FPkqW8W/6OfBw
VDDSzfdxIUJT25V/65RCn+sW9uLJzvyrr1IG1MUt49CMGjIgnWFf0VdJqRLjoOqEq6Z+3PBOvepW
fvnAJ88jfu0eZPv74iBK7My6YOSUnIgBaD/fD2mbwc/1ZjUakUXe3bhvzYibRJcl7pMzT7aOa1/E
sT4dxkTDJi3VXTdDPer+GjkSHyIJD5U9ch7clHp0gIBXm+j+P22ZygoY9KPAfr12wxaE7lpFsqtt
OZLeExNbgqDcHo679RlUxFU5yr7UCbZj0uvYk8z9d26DctFZj+/IZWwFV94H4mKh30/PHn69g2JR
DB1Mj0kxgXB75MRBBRQrDfxkd307U3W+6Z+Iqi3eTNrUnAoN9IJ2SToPkqEuJug8WYPLsJeNLQ5e
cnVErqGdCzVqAe7Y4pDk1QHVHCQ28wokbduoS2MCbQViELMshG1StDFJ+P7NMSc3/Sxzx0+a6ynR
X8ewPvxAfASrmxZzg/Q1+ZUkw1e0gpNd+ACYUFa5vHEavNZO89L8hJlgeuW07ZhcpkiR8hSyjjPH
7ZHnvYZ5wexS+bhDvxc3NcCXmJVm9TLy00BO0FXQMgAIsMfB7Q6FjlvNvHe6f62Q1TIwuNmE1ddW
QzLxNdlVgRGDKeAFeOY4SgDujOgaoJ/zbbvGKc5JRNzjrbmHmSf1/bdaoz6bH7MjchDqlrOGJIpo
F/DLp8rOAc2Kqf07+Yko6RycEiHeRXZFUR/PTouX/wxdZ5/4HhGJL3ztoIAxIQjzq99aKelCjryx
HKQCPOof1Q99wd0TCAlwtT1eTj4GyzlhZ+NvSbH30kYWvnxYqTV3G/oyDtVUnwZj8x+kvZg0nFMX
vmkrd024Zls0xwVZ9WEAHNde4AAxmWIq2svN4dJGfXUbThaKWk8l9FEAUG7OKQZdD4CcPzd+R/EO
HPHW73eI7CQA4pFI2gns9tS4irYNuQhdF9ehJJx9Znj3p7iE27Cnq1l0xbFYIrAn4zDxEWutgIq0
SdM6ugyMrKZhsVtivHhx1LJh6n01+TNTIC1J28G23f1Ev86xiaAzKjWUJQvUjab0CqfHOeisw5A9
F+y1Oc3MIyDdyQLCCo5JzREdZGx6UXwA9VzzhDB1jlPtF55p7UFuLgGnK702gHqzM35PEiymSh/g
yzkob8vJCJuV6GM/LpC73KoBqfxqzGYs/s1qQnMKOALki2q/kI0HmkVnC05FEvgqaEf2NYxaKyv9
A6PYyvdShvVung7T7b0+j1dQpPoMwO8TLFNKxTmGcVa3xyfpy3+5bE0Ja2sqHP1J7zjX9BQHguVx
YP/sq4ieXXsg4hh5xZS9Ft9ib0naUqmgsoWz4YWJa7bDOc/YYdG2RjOcclfUW0fHAnMG6Tt2BbXk
xS1F6N9TdF3VL2uciVqwr/PwozoH61Jkm+GAFo33OiPVZamb+6yr1H25FLE/wYoJ7Rlq23LQNFt0
TTNWskSiz05u7pqi42wrxkwBARCDVWx+ac5XxqUA5IZFh7gad4TB26gvAP3tW659Frx4+GiRYEpU
uLzanpNkHQly2MZfgBqlYHta6RPrbZamNfC9x/pScquWsVnOgXRmwI1vkKZ+rg5uOKwg6P+m0MoA
Fp4z9IO2nf2J3C67ecaHYAAfwyGCDRsYxbvAhBUFvS4FRyJT4PhCgo2ZbMheUQKfMB+EAepFdS88
nKFV2WhwoAxIwebCZnEI3d6Sr/IIO886/riJcNLAsO6+iJd2ZKFwv5QQ2aSbPDeNOxOXkRcpx81r
H0/B9PaOuNerPI5kmCmuMUT0NcC0PnaCNEueAaxQKRiv4+BF8fabmu1lVZr5/MGX+RKZWVsRYagv
g9fGkl3GSOuTtiCmE0mKBLrm5s8Y0U+fKderlZGXOi/T1JK/0EqFSmiyoalZT6GNDh6mKd7t1hYe
ndb++0KjbcZfs6qYPtK0wwcuOuNKsK5gDFNYeBfnC2+0JmolpzHn4hrhpUZDokulUcO8+sRSiOgA
PE8Y7Oc4x3yDQhqPZiflaB77wUtxslBwSjL7oIvXQ5R5IZRdi/+JTRucxQh91gGj+4t0rwlDckN7
LjO9KdzdrXuH6VAlhqiqdkkJt5+S10qu4RJWXqwbHiBRokyjaiTj3jVw6Xay0ehJfX7vyvxQax1K
DGl9ui0Ds1XgePnx6T+EKmE8M1yHoQiv3hreDRvgJ+/yG6vIcUZBsZz5gmu1wd1bqYHPzNwN0Fmp
/czfvkxqOengPvVmJKlLU9GvIDr3jUMMkh4846Fi7rWG0/0dW0dhn67graOc7XL4mn3GdK2FwlMH
XA5K9MRPctL13z/ifwJfttrtkraeLyYvqGFHXZgvYt+6ktSgkiCvTLaRb9MrEju11KOmLo7FtdQr
ncjlDHc40wa+uTw0+J8L67DcUuRNOSstJ5rJeVj5QFiPkzSX9SAJL4kt4+RdQweaM6mbgn32c99T
iz2GfCKLyTfWqdMzNFrB/0LoCg/ne17Sy4ZE1+UfhRnx7Z5Q6Dd4LoDW4br8dcTpldUkkMph9n9p
7jwp2zLkGlKVPEp/JDu7fHlzDc1NsxaCpo4RgTkUt80lCtK7huuwgFN3/phUtTWX8r4VnmCEFIeo
aN7oq3dU9d5JRX67UHw1LwgtIpe40NDmSIv4BBAUA+OaJFLraNZYbGctpnUZZ7gcgR4EzLqDP+uP
6yfiIhfNTvl2jhRfgh9aEVEhigkotmj3D8PlBKMKfYerMrkKpiMdIsH34IgCRSzyQkWI9af3TbCm
WYxZ+xaNCZWeO60FqHlwyC/tSDwDL1BnhcOhvXXb9hQOnNcB7fposiv6cHuZN0rUDCrue3M2zbQb
yAOWFd1GL9ATHrrqsfAKGIHFZw7lsJBt5/rd7yKny9QX6fn7HqtFH2wOlZIQoqnfqRvC6Ysa17oq
TH2tmPuIti0ZPNg3wTktcFaB8rcX7azkkpxCPC7v87XBk9IxcG3zVLlb8yXYWXVZPwre12cLFIpK
4g2dxcakAdeK/b8LEWT29UQo29S7H3XGtp7fzt9BWNuSw2FXvDEf6nU5PecKPYtiTv9eSxtZbT/U
KjhpLBBTSOUwXaNC8xcOYZkLfCFUNUukhLsfFNKpIhNvdaMXWOMGjgtJ+FgwXYWsSznyIE7omfAb
DgWKnDdgpD+q8AZ1M/Q+Kcz6A6nDiPLIC5o9rLnoafwanxn6Xv33cizp3wZihzhSq40mLvo0DIoQ
HgOnJakdpVO076fFvZlIRXx6zlQ3SOIBT4tF+KXGVZW0O578GY5F6nth4iuSDU2CYc9PzRtbR21L
eorFVKo+DNlfm8J7dRD0KSzZl/NmvEC9yOF+fA+zLrJUyjxy3O1auNKIUU+nDrZLxB0rrUl6HxrY
daAbL7LYH3Oydt9oslwGgChJYYnDWH3MyBj0q6rrY7nAI9SbTTIl7uwImGEtc0um7tdi6S0N0MNr
q2taKztREffDKn01bih0DEuiNfGfCyIzX74CppjxylC9omHZeLRDNgJSDoICOcAVmyGDtYdx8HHN
vfYHh6iRwrUNAQ5AahztdnI5n/8ZXbV2pCK/UyH76UlS5ynxjR8RjDCy+qAQWLTV7puwuvFuHwv2
hlIP1/TK5vK3QMbkQRTFR9N0JsUdoCT0sRcl2X/+FSBviLxqNwP07eDQk1S4Y4wFsG/8V10kgXdv
/DhkG67G+4lzQ9x8L4pmBFNaGg5UZvFMjmoZZeP+cjtmlrRCM896GbkGC7FgjFRMOV8fBlvS7xNg
Vp+0AM+7hMbkohaq5yqPXwSw5lmm3fWrRisVzjd6M0xEsz8CYDdtucw0jaTW7N+hKDUvl3+7fYSa
agJTmMV79ew6qoj3k8gjr0vSWPPIUzzM4EV9BUcFcxTOOO+D0ukUR7VRbvo+FVKQN8fzaQC4Md44
67RiU7QdSwNPIW2nKo6jHjIYK8Azd7BPazn9IYWKnunkTdewk7cVGp8yDJR6SAj/dpdyiRi3uKEq
Q1JpRPBOcvQjKQ+4B2SvqXFJ7VVk3AIGPRtOxe/rxBqCoTa04NVXZp4jLWITDBZ1ICCegGVABAec
3zlFz9sVtq5pZ96aCxJenpWjd8eTeS5HwBXzrC4hnQvtAz12C/rbQ20+qTOmg1et/2ZN2map4F4V
gUvdy1WEGqqgRTFNlq1eE1eErOTHM9zO9XQcOYvVLajFHk/u0+kSfoRIchhY5+3KAmD8G1LVntFC
WEBBoQTpX5m7XzfWImxdagenn0H+WmGSH0zt6eED5xgMKiYxTbushMTME93RRiputb4Cis7edPpb
7if2i8Bh5u0EiItcC9WNpJ/EZiezrh2BvQq2bO28v7DoiH5yuo8CEDoOahq0Ycxxf/wzgTs6ciu5
3xjTipmEuGcgyK9MsNpe1H3MvfHZBybKozKgw0EPdwhxa7dco/8jDnROIafbWAY/leHcgdYIxSNv
ePCRIL2s2QRAREfcwlwNOVqnQkolf6fn9iLeU0rloyWRMlDdGdZ2tHLSO7o2Jy3zpejBF7XXLJBW
ppRfB8pWxxZeIKYzMAg4RFqUOVDIj48cI7VkeiyhkaiRpYVXsY47UpPx4tOW5j/9DkpLNM5YrcKy
/ygVeMeUSf4+TJveqOGjVZaffaOktgQk7zJOhSAZKLZpeFBr7tODqwTkznv7RtrRZg9/GEFxJq/3
uaMWGrZLT3NVrYX0iyE16wW7n1jCQmVif6xmlt9htfFvPYXdox2+bmeHYF8snywE80mFh5oqvyTp
RmS7HHDYlLuvQlMKrcFOXkPaAzZj9YwhhBjjPJVoLVPMpyJeMPBH7Uq9NA4aUiC7eH6Kv7B7gkLc
1WTl6wpp/VdaNidS5b4IxcDSRspbOOdO0b4tE9B2U2j7buZYQtJeFNA2g/ZwV6XKHBwuZS/9iZUw
8QROIFsFpEorKv2tk1eBqDIv99RYKoRgklg5CZ2kcABw6D+FOf/9qUQ8mMfD9jZqlNu+puB3GD++
lxJxOXI8NUgx+KFd8nadd99Wc61fXdBAsm2v1CbCZ2Go5Vm6PxXXALnfowhEyGRHsbK2Q/u+/sIw
3q/SWi1bIRZ3WDa/FoQGHTuqLkhZtP5ZIb9VPwMaW5JgvgCuECZtN6ie6L78E9lXKgdA3bE0EXRm
cKfrz/wg2IX7GtIJovIs8Dxy67i9gqodacAVKVLQJ0DtLF/jm7HvXlwlhhnsmv/MaVFXCUenfWB+
j9IlL6ahZXjGhl4hrrOyAunk2zrjCGeaclY3YtI4ksStfR1ngJrKVWuQ77oyrBgaYE/CjfqEgZuL
nInCNIOOCrfdWdMD3RXloxLEFC05A2cZZb+97aHFY+qFld6e0eRhDVXFrYwjwpX/HC64DpCtxrS2
kz4epVuQKJXeLakskzT8pFg7JQF9ECslOmg7UhTebx1Quao4m6pixJ/ZpNpcGYJzTKB0WsdncsFW
zYZ/P6ZauCBzZNsmbVFxbCh6Hr7JEbPomb6wjXFybbN2KXa0vmbjId6XUNZdUm2JCHbikcLyNb6w
dWLTXmyYatOw7VEjdY42V9zsVBcCkUVu/4C47q/uDaoryUqdGMYau5/Velo2ZKisr3Qd9hepdm88
w71Rj7JIwCAZuMFj6ktFS9EOq/Hw5hjVg93IbOy6+hZxMbfp8oWVVfiRk/Nh12zmtCuUnEOy06Z8
wkNiPnk2nMfH13t4o5j4iiPXrpbfVhqGwq6pByFLigFbPQW3t1GXYPxDDQxPkSXGYc47O+Qp+faM
D70tQBE4tnd5hBg5nzZZE85c9GjJhTmVjpagkXdkXjjXRaY/HOmfFI+TOWfqjcgZubbRhNg74qmJ
hp3/svNB7NrjqxdFQuxgthjx8XEdjGnFWeLESbVb15E5wADyIbqtQZoXtQNIL59h4A8085bpU39I
FxB+RO2SnPOUWRmICknES1cXTL/I7/e5CgvL7iPBGvXH9OiED1rkYMnEyOtDcb34Hphgh4EBI0/f
XfTFRN1zHJq/K8k5Nzf7wQ72blgEMEjgo6K/HOrcXJtMwxeDX4m1IZk3a/pIytOGzMq/k4v5RM/P
ARycIUoW0SkQ52pGOGuEiYnlEiSsCOQZoOqO0CxbHhTGhke/+gVhBFC92FWjM+wN1akPrvCS73y7
iDNX7ligMjBbCnvgcR08BuXAFZvUz2fvRy76YjIP1sT3100EgpW67FWzgO7QB+lHrciWbYgn5sXb
iXOF35jA/GDF8ZRtZE3bwSQN2Z7vxUxFncGaACdSDIs7sD/x6FyJfBRkOQh5R0d0ORUeOt5NB//X
/mHbpLC8U7IZJq2OeO5M4Ut5h1ng9gSMmD6WSkZGk+CH0EdOJc+TUzWipBxN3PAaJCLUvxKDJ7Qp
lj/4PwVzQm3REhySXk4WhbvdhxsCNr03ArxxwRHuJ9p06otuoFtqX19yy+SvqOTDyIxE8LSluWPq
AGEhyzyhqQTO7qckL5wyq6lp7PxUEYQlYAVYEvLKgA64PZzb5kszZFTf4+6U5cOxjEdCReVfwppa
9wFZHeAjr6cdZ2emBtvKCvE/OfemqJ8k+qY+QdempUmYuVWzdZCchzhrA82x6+fFi5SjTFUtDLeJ
kMqlBzOzIjfuZqVtJc5vqa9YBo1tVjiPw5/1WjVyAbs2XBoWl2oa830J4T9/yYiqOX0cDI/gUKBC
b+4t4J80L5I2pzL1LaBaZ6ccF421Y2s7EXXFYtO6QbiOzNEqK8c+fDsTehMcoQ+MgK+0e1h8Kj+v
KxDyAyKQDO+6gVhF/LMfv7wb5Mv4znK/hMRPKAAN8euTjX+GtEmqSDrBzgxon/F6eQQy+yU+YrvX
y66ISTWcWWsGUU0OYfPgAeU1GU04cZd5FQJkzT9a5sJJxAsDxj5USomC6r6COwm8s4rKhPYvkk29
Om+ZRqm63M0XCHwbkwUlXUIAiLX0RJTWfIWWxuQLb4Fw8PGfsnFujQLFuRCqpbex6gtTUbLh2b2L
o+zGillAYDmibFZX45FFJGBDEcSUhHiwTC/KMM1cz3cZ7ldn2bPANO/3rVr3t8zaTD9ElaXSnzG/
NGNmXWB/MMFdnz10wnxgyU6XoR1GXti5a3kolt2w8YtDB0iotrChdC6V5wjwp5qrGFkI+lpmJnU5
+I3ktkWUny/kQl1SeBOdkB765FnI5EEYRdbblM2uaWOC1Pw+bM1XlBwbv1KUvmUPaI+nBs2GHODD
hDrBt1UfjVEVQ+3KXNQQ5l6N5RzL3fGbWpQUUAchSANWgiXhJ1b0oXiSrXXSRJAGB0snusuB3O0q
VWG317mKV+757B2KemRyEr9MfgfPoYf400f1NggLbDyd31YdZ1lJFhZUcVOFRDtZiN+lf6b3OZCG
bvmAp4GsjxaUVwCp9PYZH3Ffq5ZrwZM5yp6j1OELrZrl28k3hdWvEHs8VATOC5U2WUyhmW3tF8S2
aS2QczUwTEFkNBrJvn9iXsu1Ze7MuuaewfxTFsVrIhoLIolz5kRVENucK9pM9cX4G7tF6/jApk50
bmHK6seQJEP7p29RcGbxTb61++X3KqaamZtRHRxmp9Y3Ao4ejPtsx4ng/dHFCGhH0ViELOlq1E0B
7d2CfwCWTl5LnkpkDUBNu9uWnOgFe9Ure764HS2SETXSZag1w2kep2bH+FIAg1ApgZ/+F6BgzkDa
Qo0nVtA/1qVlMMz530RiG/DJOfKPyZho/GjMo6rKRRUZBVHlxA5IocQvadSaus+LxfXXFM8/uxHh
nHU1m6SHz2qLwG5KPZhUhcMLVYWLAbJ2+czbkrB0v34fA51m5vtvqu8XhrMN15HfEPVzU+5rY7Il
JU+Nk9Iw9b20+HsDN7zC6veamZE1gavqkAkczcQSekftN/3riUdFDuLBfZLanUmr6/WpR2rymyBA
ZapT7TGjbCBv44yPZ5kH38U5G6CLpn0InYjfVbNi5Jiq5jINxtbJnj66vHlMIqBFETVe57hzg5KJ
qDUWShJkgHdbNLMlhs7ynfvvPF6wYKhogW46/vPJx4JH/banqXmN7OCi7Nwf8TkZSbm1r/6cPFC5
jF8tOXYCeO/QrBJcrlJD0EfT9XeacUu69PgcjFUFBk2wgufXjLEm17vrfHkWfsnfqlWyM91Nwcr2
Z1/dFisftoUGGDdn/2UTKaPOTCh/5gefIFN0o7HsKOBZiJvBqpcFeoHuF1uFRrlkguirNX6t61Ao
pvjG3+9ha3xxnDYKC3EMg5lPeQelIwzKuSx8T/MXeCUXtiDblvyGXD/ZzyBjQdQTO8Gc4zO7Wg7C
c60bDPzS5hvoiVCCi97WLT+/K2uGSejxzlE8DWGI3A5nsqxG1aTNP2iA61Bc1qJgRRu3wea68CWG
B+TwJctJ6VGP5dtYJUTafLCIfkb5bytsXYi/sg27Yr9GK2a+vbXyWXKdNqDCz+zGs/7A1vjIayZi
L1+e5ubzAKl+AXmZcFmweG9rgGa9f2MiBKdHcZI3zJmqT5tjgYhZIq69HUvxModX3pI8yUORJNdG
a6X0zks9YC7aEzLNh9We3BzL65AsnNDYvpwcj1JH53O3nNjYTVaDUm5C1xqPmr6WgBHTR4hKJod2
59xHo40HCZFOPA5j+Aavmr8lrZJvUxY/a8J8YKlaXBG0+c2MCz2GnvzSPUrx09rHzT74MtOcmqqF
fPd3sTtIkIz8cdHM/0t+l0HwyjZWyVjmgVvAJ9BHEF3c47JIr0fjneqsTmrsM1vY8FJ6CY3Xto1y
FoWUCcPkGW737jsp2n2Ct/n4Q9apJnvuceTznUKBGjq0tMgY7tyrpk3C6WNiErCj8JcjJ7iDarTl
P+mAvrk6jWeimmVbHAljBlwT7QEwpNpJv4eH1DHn74XWR1dZQf4bg5UdG0A7t+i2hd9joTgColHJ
WrnyG/TE+imvy+chOfMKTmeSCCa8iYbyF/zF0nosdDT0OsNis531WJUGCwgWiGmJBILPLuiwDDxw
uu6ySRAcyFWAAi7XEqO/Px2iwZjbXqzj+qHeBSgjJfefDtOqqUk+6BB7kMZzPYRLwxQOfyNZQBh/
S7alqrGXEAdeCuclVjiCYDvWuuOTz1Z+6Dlq0CLtgyw0bZxJH/Qt8VzWSmGAUWptEatydLjTMZlO
IgDpN/S4pOgaAt/i7FSRsrNk5rqVyFUksYVfKjAoaaehEpM0d29d5EyOJ6JQRhb2jwMBR1m+3r7K
EYJSqcIK1c3XX/JNRp2iDw6hPDBvz52HvT24xLR10Q6PlEGtcgXvw0CLPFiwt2IHW1GCRqEN2fjt
TRhf7XMOUJ8UFpWHnnS0Qbp2f9+ephWnAr7d+PY/AZcaicB0GforDYCiIbebHM1st4gERMB/Xrla
g5GmRDShIgqrL6yvDW6A3+5vraZIQd5NgSbw+hAxjut0pZ7DPMHDqLxFJ8OGw8BExM4AUiM2JXXR
4jU0RxF6TI3Ohb81NPecVAVEYrvE2Ia/q/P9gBbkaCnaNapI9Ha1yXLRr7K4tOQppc5bKWzoe8I4
StbTrDfLHwgQFm4iZfkILkusC7T1eoThUMeZQ3puvU1eKGvkAVarW92Ir7mxWTouRIERIQFXsRen
RJqnu90oKlLSMfo8CNo5UIurcQIL6VvFnY8sqaQlAb8ex/dsiLBV6bUZXaRjgBmaqoNx9C4xfLkT
rR+SYWCgTiVnOXsSK9YhiFh2ovvh+bWeg0zPd9piAwf0JSH352epyI/WMilasymx71/tHd0WDLXG
4unLCqMo/vZwDNB9OlARxVKGWFT2zEKjU/4ubW8jVOOXzV3d0WgARrstUkfAR19Rf2l6upS6U4c0
REKpTBLmvQd7/jdhuIr10T3CiW+U7LJcBErqtXpmBWAqgUxYDopyb4YNS+P1lfq8KQUt+nyfHIe9
cf46xCBXkFSkmSPqaD+OtrBOZwuJMLS8ZWxLJ8RdDcCI6h5oFe6Uyl/tsxXRYLRB3FmigZMAS/eP
IH8X6hAWd1m7cKLOIVhB0A9pG8qVa/fTxQlB0RsPUOrFoo5aoF1d6lMd1uaRIpmQIBM3A1nMusMO
suxlumN5WoN216hujaKoUtxskvWCRsTSIYwLnwvI30z/NvOXw09uBsTDqfZV4v5bMCtJxShvw5El
2DZjEWXvm3YHNgFvA6PV555JsQJZlI8IjEG4ZpHOHcOiPVii2scrX0QoN7jlfbYYu9M2RPfu5ycl
OrBTX0vkccqiQmkLFfGs5RZ9LtsJHbUoYmTLdcsg8mOgaNl0H9ekh4gA3k7AXh0X1tti322bQWzE
dgTnxLtMdQsHCuaA5yLgn1t9onJwmq3TPz+1BVZxoQqmiHx3VocfVBhmd2lWY7FKtpazpJtRMuNH
+aHjVVi/MYEqKrJl95z/XWyt3O0qFE4oOiu8VmVw5rCrU9hhHnEd2rzVDZVEdwREuta0m6Fy8hJT
V2d4fXbg5lSd8BPQlancni/WeDFutuZrM5TvAivkGFzHh/XGrljzHooFtS2+wZrzIgsytTKxtk5B
P9YwhF5D+SQ8w/giPKsKv3HBDljMDw+cbLIUy7MJIz2qYSC2bNV5n8jhMvdtqYDvyWLF2ZfzZP4c
dbqhLT9d9o6kwE8rWg4BQsFtqk/iXlHa+3OuCSYRcWBBypSwZaFPQUSdFpW4zsq7/pXec/ZFjb8y
wfPrgAgkW4E/qpG7P6pHamY/FFPYrHz60hoXFtu7j9ntotfPg4Q9SN8qFmIfXynogVy81fC5vLzy
OWnkH4i4Y7rlzdGuYu2EiXXJkoDd51z8noVj8pEfKMiZcWF1Yiy2VthqPNSo6Hj16UwYY2qyOKKd
3yHokeWEY/Jyy2XlQywlwl6Go2ez57vamdI4oZK8oDnYC1d/GpbRzguwtG+1qZUaCdjAmlidh6Xo
HriXcMhJNpux8T8mhT11yWXX3+DcRq8fdAHIc+Jhhq7x2dWgLiCa5ChmsCcITc68koLmwZaVZi+N
F8JY9LNr6+IK7dnU5DjhBMJ7pnTK9OEXEqQaifVxa1KWxJyXZJgeUQTtNXGkKvLSiChNb4hUz5Sr
jUZiYn9JuAmxfwzdd6+AysaHzsRZWT1x7LtnOd5GzhB1hBSDrk39+ZRhSFlgJQiAJ0yY/j0l4y7J
U2RL1O5bbCI30WJIsWdok91gJrfMipOV1KNLqUJCIzvLL/lpFxM48tfuUMDEAW3dK7m+jL9t/Yb9
b0V034ILQ1gFAcJ6JrAOWJsgfiIYOSsa9tmfsAaL2ZB87IioyuyhiNfyPezk97QBS6AfpCkdl+99
oij0794IuiVbpcKlDspsavdxkJgacLpbrrVK/bq3yx+XlQAenMLMTGmN0qcXfp6BqPMt0lGUVxZc
MnmV2aByWtluM2TA+OCmeOkR+SHiHQvkR22oktD3XGWIVma3C0EYfR1tf69wL3OgixtHDV1lJmNQ
5ee9xEi+wktix2kOcC10ioxdIPi52DSI6ZMIHEF6Gak1FDSKRm5BIcS/1FdRnfuB1lcKwhVrSGcw
v7QCh3jNvn1ru/bK/cUOdT4L2AgFoJuCu3Rk5U4EzpL4lKW+x259LmVJvKaOH5hJdOX3k8b0i9DX
JVg/kYUOz0HMvlmYpE9vcZxA0yiR30/+/qfxmNotQQPVowhyelJIeKcRj1JJFPvepUMgMCox18FT
p+ar34q5uVJraNQndpwd2R5mVxqyyeDKcc5j5sJTYWFtb5NKNUywxGLztnoHBp62fxgxEIsziA8Z
JMsmPELgwuvG8kyBrR4N239RUavLVRXizCSwlPYnGy5LqUMJ2UB583StFo6eVU6NO5y0+0BrN7LV
fpKBJpwAGkBK1/l705UNQS3RcQspxFLpNH8LIKJ6IXk8aTlFcVD5G9cPJDVWI1XH52er43o0/mdq
SnBQUmT011WVFjv6b/VmLXuKQENm1gu5J/WVCgCFZRVRwjTKbBq1liXdCfbP4+CTymHjwdyJewGE
d+LsR9F57K/aRz5hYSL/bmcTurIvrICYGaoTY6G592kvpiZ4LHb63FYvpD1I7uLY2AcM2wbbsGC6
ekvnpQHC6P34XA9F9YtXzDTlg4dlCCiOdv3RW3uImSh/EOKSkAwB5+CalLsCPWmhp5swrxgwix+d
5AN0m/xf7SBTg8C44O1idVf8IjUoTbdr1IutSltQVPobl5mxfYMiWVlirTaHFLaNdWBVQ39dy1f0
G0VBgbYz+q26CrR0HgK2zrq0/a1DRhqlsKXKQQq5KysRaaukydxZLrr6E+KozolDluDkQllAstQF
/IjApk6dYushMbkDGBg5wJVDYWJNZgzZW1vgNS0Bah+mCATziQxH12QT7OUi2a6cF4cjP215Wx91
MlVCgqACt/7w7xagn+i0NHaGgGCJrX2yiz7scFXnWAFda+NfAph67s3m5m/k/ZmEkhnPkHZxntul
3ZYRirJLy3gmq6Q5j6ccYtbodlFykgtMrwxvcXhFRP9EK5+DLBfoi79YmesADfnWYqEyNcKOuiRK
xH5FsGM34TSRDoZ4M+75DIYz9VNhraIx1J2wcM88U3cxhpzomm7c05jQa7cMbFFftDyeULv74Dd7
L3m7fV+BxxMcyw+Lwhio973tAN7ETZ/djLkNBrYGpzGfAwm3sn/k7pmEunK7gF8y5bE3BnhXxVcX
zjWa+J3M/M3pRIH7O/JQRcCs+/FiB4PNAR7jMTqnTJK9EOdXYKZfFPIEC3my/KFALn9EOBW27S4X
twgBumOp0eWSy77mcLT/NInIoyrBnAtoUhgu6548MncAwuRBoE6DBGIViT1pBb9ePSsRIaLkoKTF
VpZq11f2Uy52R1FYR6zduYCdr1TZPeEBk6P0ftqp3ENz1f2QO8D1wbTVYBoJ65kbqS7vHQbDkx4y
Gf3Xt2bV3VXUNsmPg0sZuNIv8NwWI5vZVmUakqgHyYpbUAC3jPHTwG7W5vuHHB1TrcGBqsCAcvaY
PCijeH50NzYm3H8cgA/S7y1ErPG6gi/scVvzNl5JRZa0dRPX0mkYra852d7X2ngwjnlqGrPxTmRo
AxWku44Gnpi5gAtYGf1zymWl2CJwKnPafP/Vs4cQfeXkB4N3GHRTwxzM29PFXR2LhXqogtGP19xI
GxmlTfP9Jp8bn0j2Gg1IVAg9q3SjB+tEDsejfYeavqOV9KmEnT9/kzz1G1U9LCGjbdNOujvLUfKH
zezdy60/+gqgY6TAJ9aqYBiH0E5FNpttJgMBgUc8tqHA3hegYu5Cw0jWmLX1ez+B5I4fqUjcTG3Y
kXsXGSyTDQfdbd3eSR5sG4/y60NyTfP3T5PemD9jz/vICi9EelNXiWoGG9+Rrm8LbtXvGnNl7huS
QumpLaQTb4Yjxa5yuP2NMPzNfEy6NFAxsBr1IDI8iuAby8aOjuW+j0nWntBLDmNyscbJGn7Y9HWJ
nlmhkNQlY6X/6dK1mUXvsbdwJyqGD2poxHUl02VDkkNtIv5TZ5vgaNZA6AAcMbJHaauaIFtmmeLd
6pRT5Iqbu+t3dT2qaDro9KIijAzty2VJyQ5beGoTwFOl7gHodpIt6RN2iQup4KbSwt9rls21Uhib
9V5v45ai63fR815vIlaWIjrO3az105hC5PXw+YvhzBX+Ngov16Lu/4KgSiH2Dd54pysHU5twm3Bx
goHrL7NLZW9DXDjP/OjKI2OYkdm4yfeeazJm4XeTElxVmBzmaoZG80s30AX32nbGZW6ALLQB6mzt
1kJr313SclMm+HDa+eX0DK38NQpEqO0vpU2Po9oW0ONJTVksE0OgQpWtSNRau8ob5BN7XC9PE0h8
vPkl8xB//gQ5q2VM7hh2/ydrte5kj8pw3ObBcQiUh4ht1kCKg8aqXlIbJhbh6GNX4R46q6nY813+
D/KRij1FjUPQW48aPZGpOE8Z3mDJDMVUC9EbQ7DXs7/OBv4BOGH2/EcFe+HGXP46rBcaOGR9aTmt
/UXNuTZeSyUUg9aXenpufPSwglxIP3nky0CRZHm4nlOKQPH9w0C8klcYX0pqZmkleQN1gKh5or4O
RDi4eLqZDsx9J8n9CsC1skZ7lkgCpYeVXmqLaHpsoJFF71xxTMYumOVCuLW8SSPA6FnMG5j4rh/1
6uJjBOAsScVvkpZMgXLk0Ohy3qIOiwAzriNe5KEyv2Yyme5UZKFixIFuKM0Xpd2NH+088oGo7Jpk
bgfyOVMDbXCb4R+YQaivu6SbdClpmZBtyfZDpLBFbIzFKK3crVh8wtc1m6HRG61N3Byf6EPOA4Y4
BMKmZi7H/ypnX9TQghVNT8PxlxrKc7tTDBkBZzWmm+FOzR/Q0Pg+/gBws6smN+/UqMM2rfoKbe0V
08KRsYmdIjvdI/Ps1TyDK2IP+IMpQMitMXUXdU2JDtlKU6bD2JPVnbSk6QuLF5rnqCLGoG0nzlrl
IaoTLdovIzORdvZOckf+uvhzDb/mGUt8X4kGdbw0dr0GtTAX2b7pDtFP3rRg8b+afIP6Vju9v3T8
iA3iuk3R/+0YpiLU05HuGlp650dwDunOLUjKjBdxtqxvb+ZMvr9bZIdMshm4lOAO0E1VIqopWY0d
bXRiLweMR4CYeziteG9wH18rr1Camld8dPdULPo02oF1HhKrtpuQxXRp0wHhzlph+7mNisVV1TH5
cVzrZPS4e5QdL1DzTdVd5eUDzh4KzxMVNMM65E2UgXlwPvAyYk7GiN3jAhDB0siGfoKPem65RRLY
uvQWx/znxP9ZeHnqtqMHZ7ZRBcengXjXKKZMkebMNEzTwdLEs0bYdBIGiu22wrIabVHWH8LmFxC6
d4Oy4MEQO9vb1LxY7ucPLrp7t9a5sCt4yQVRG51MX6LC4vRqzQa7aKDfyZN2kWz2M//le27/M3Qc
vp68dQAToCa8Q+rmvD33hi5f22bp4uJ2Sb6ykCKzgYvERPxGdcuWyypHeUETKcJpeWZ2sjaZSVCy
zMk4bxpVZ6p4O1uSmYUX/4EdycvoCsZxooDOLR0S6mVdO/DE9ZkCgDogo3kfB/8JNUTKB+LwxeIv
oA5MaGPq/48puLUdKbsGjsGiAUnUdNMY6TM1U0QYLtKSgGkF6RIlfU3WalXiIm7/NIy/H6E/4TWA
wPqgtyNHfZMb0yfZZAm5gK0PivzqPTEaMWclB3dupVOg/1fU7qkGYtPiWDCSV93hSP7h+0wsjUJa
3zv2ULDbqga/+DL5wTN8IrAza+32Q0AjbWgHTq/eOM+pdP68K8n1bsDnuq9BvI7R6+1kZ4my/oh4
b0q35wxz8QFS/ryK9R1xM6wSQwgQVpX/d9jtsARZEB4UZBAPnUkLHxLJcxRyy1Gu0tuTtaDWeYN2
s57Dn6MvL7ui0mhkGdrfGy389bigY4MbPTY35LB1tR4xvZG3ycVkUc2d+pqFb+zT4rC5c2uqY9R6
NYleuyfBym6mHTXlVes/mBnoOk4TMT3e7WECsq64BMUl+IoJAUzxwCyF3RV6jbIRAGFHKqo2ooPy
BQKcmNBStuRAar8hXuzVFwqINKmblKInNuTrHHMjxYF/YN/ZloZrdsVvfEku5BwE816+cMJ6pkVw
hcKSq0DRTUn0g6LMBRCoXdj5jevDMRrogkDCEWJ/MVEY60osTOpJBIf/GdLrN1cKxWCPJfbqY+Cc
pftAn2vUPzWI9BS4poH8KwxYHK45PEPRbK9mmPBrfvqXQ2G1+QloLZDw3zqtZ0IMxQa4D/mbf12C
LzeaPPFY4GuqGFVlO2vQb/qEyNTRysEh7jYcFfyKZURVVGS6SE1cWKuGSDxw5xMQlWiQ+Z81Cjdt
8Q8tygvtRocTzgDrdchEd8J+R4LgBnVmm2f1R1CzBTqe7bPrOy695NxRHHSLRg4tPo3vv3WQSTKD
BsETNfVR9X8Nw6a6lZqImP1luOvmh+0hPhM1woCrty/I+bgPZQ2q4R20pKjee2m+cUEE6vZ+EKTC
cI/HYTMWgzPhPlJlbXXTNCC87YD+vHpkkfNejB5PCnQgodTDZchc57AgcxC+f7LbaT8n0jsorWNV
27BRYEVzN6C4jmbjRev0aB3tnm+UV4LVv8SB+S7bNdfteaSKH+NtLk2yJPIlArKr95bXF+f60lnQ
lY4O2ZUWohHFHLn2lJbSLc3S0yB+C9S7jrKi/SDH0r1js4aQytais1gd76Y2WM4j3XXruhYID8po
mVklApES5VnbsNJBLRNhCIwvkmtuHC5QiKOAk0Dn7TRMxX4ogJddbz2X3hrCm6N9ZNy86G5m2ikK
PXb9GA/Jpayu0nOIYCLpP4gsl0jzm62kjcxnZUAoAZ9zGqvPvFFgNQgm+rF2nx+QmEVbPKP4Yq+O
vwdILhc+c7xks1MhggIlZUwnHG8libJSACuTn/zzCpKbafyQZupswkybzj0nqU9bXTQLd3IJOR4t
6LxybuFOfu8hduL5WZJh9LhLU8ngZyYCDdbShNs0M+zagQNrf5rYL/kIUWS9MQFHUSUYLPFcO5Pe
jlM7OhBrW0faFFx4bp7ODaoiM/Hr1kWeMfdK56+kKJB2jg20muTS+84PxJj0DojTXWSPDuh762tI
7tS82tz3EL6GU+YfzxQa5YGnINlA/2koe3hI4irslTcFOSAoN//8p00pOvV6frto4ji/MH7qhukU
nyUEty9Ss0OI1Q11ztJvcMS2Lx+XxCbbSrVl69unQbTgB4IOP8ltxKG4SsXI2Ot0gG95SGxBPtEJ
WThUoNt496cJ5gFNH9cKoi7kOtVH9emv9ROzwPU0imgik3BR0OJj4sW4WP78OmU0n+jo8t4HI/tL
j4/vVgVayFbcOcPw+S4ebYhBtWMmwCaBt4Qh0no9crWEC+XUOYFtIz7kFqqCgPVLUpz9FLtsWHoc
5mxYyZPVaw5uJ5HRIiG9LSqttPmuvNwbidF7imkV6xVyRx0rDnj/f5g121vjH4UXs0UQpFaBbVwo
vwcPR4t1V2mfKz9arvX+w3HxwSajBpoI4upqPzHdh7CFdhdQQSLIAKdzmwxYHH7GWj+Kn1lphghr
BzTmS6utdh+eBcilLdKBdKgjS1o7gg9ASifCRQEQnoW6s94i93GxduuaefKsnnJfFmAWFrW7Othd
8GzxAf2mp2DFl4ufEzimo4Qc4JykJKe42d1XkCCLJHgFOjoXlL01aRvo4MdAXg9tO25segTCfGl7
YObiDJYV7eJxXc5H+89vDk4+WnefBk6Fam2CLR7woTAt08jWHbByGVovCpNkvNGadHGOWCBlBcdF
FY7/fMq7PpDnz1kElsNkbPnM2okj0gsrUPbe9sZiKuPgNlfsVM1he59nIN9jIBlpTViDHhN5P/Zm
YOSC3FM4GTGhAGCYXnOFNLwbaAMySEE3CbM5/tadew0Qq3qvz/7VpfEsBHXULDOnN04qL7GCTNQ/
DeNKObseX6TYEenYnpmDmsdmX3cPm8l+cMApJPjfJNagtHHjzpD8JgBH4ExR9DGwkPkofaHe1t9+
nJI00iDMkReHJY3pFWL1dDQ/fD9CDfEm1utDcc29drsher4xsPGYLEfQbAAXKPQdOUnXHX3zlY7E
Vw/x9uxIf3ZSbDR8NSi+jEoZ+fB/1lkjZ+fzCKNtHIIFDq+uBzF1wWAlkfiNnW8Wdvr2svraTHtw
20Pnw5SR5pyMXVMImtcENStRSDeBNAfPOW3vdRI35QjglcFCW0OWRByNq93YdbBmiSERGIxll0A5
o0UC/euSGGbGhqeA5/s1GGPRc++c3nms/bPB9uVgNl5lSz6CoS0XncTjPVwlurTmxYyVamIkDz7U
TLF72iB2X4SpRQ0EPIDqop1tjJ4MQQaRCe5DPIEvz3sZQIegAIOyRjM0B0f10J/MMW2VO68QIxeu
RpMXPtosIgj0BqK6uJC9frxRPbG4X6YTpFSLbKSt1mrNA2Vv1ZcpmAvVv7wvIyrPO7bYEDCAJF+m
F14uOvo/ivKGQqvwSYk+favShaKh/vpA5CUbAcoeShfrmUxuWCMkHvK1wLjakGEm1qpLvKrZbkqa
wBYncw6OsItUdc3QEnQPjtzFUgOHmdIU8JTagXMlVd7qBEeOGo5PDukdGrJLDgljhbx9E17CyZfZ
ke9iiTC2TW/ERZq6d3VA8QBlUqXcBX4fQYa3Ya3e3hpdRUlXh7IOJywgktrnT3rDlAtXf3bK9VjJ
pFCx/dloz2CdFsFdQsFCc9s06TXVH1GwJICITefq3LoGa5PsEjMQ8xQMRkbaAHF2bCVw6S9rwkGL
JRmchGx1ncimoqDItenHO1kKrK52tLkPEE99gh3ocjpoqE6fHFrqOZpLkIS5kT9yxz6uQehXVhXK
xw6CGDoy0RTz+h9+XPPxMNPvlqZXAyzNKfhDqXyvzPgwY9Fpdjpg1r3ZqoX07MoABJXnyUsISPRa
cbj24j+sIHHRNU9ZEg67CWRZNwCfozxS0tw4aqTPT5naR4XKMhEV67pZoEbpbcjE01jTv1e1W1x6
wWq4xI53gVew8zaANlwM3DlqyBKLmXInS3GlqhPMllx6HkGvpVzgjumynclTJf1u9Ckd8gcMqUst
5Ry3DfwvOUL1qXL/5kZrb2dJNiHgRb6mN4ZR+uKw+Bs5gjS55gWlPS/lkbJj1anCzthj8/TEsWbt
j1DPB7TGpuMXhE93keTzI3vP55X/vEWc9gCX7AEFDgNB5IGj6mKPQy3WPtpj0/VIu7XxhnG8en1Q
HAWGWUhtJhWajgXKHvY3UX8gcc0HFgBlAqprlfywl+eiHmz8fY4EVFuC7d2Bn4ZJJ7rOGAuUl1VQ
m+RFjgNxTWeDzrcMsJIy22B/J72AKoeeD029Mxcudq87Dgrtr1aRvmhQxHTINpNayAs/cFwkZTqu
E2Hn79N+SFW7Me9uRolSQb6CDzVNwj3ELC8BiraZNU9e1sb7Kb1lQn3XZGCpenpdRHEJ+a1lXrYF
EdTXX3FUqBiusLhzpe3//yUpxYIQj84Yo1jzKWLW01pyp/dXGGFzW7Of9cS8KQOiGL0X+EtDoG+k
WZzlPInJlDmiXWnkaSRdblliPGFIPt+iOr5BkE+nriKnicNFVR0EuxSBe+LHbwrd5VMdjKUjpDuw
U6GLU0Lq9SiW6OeTPYmEH9GVacn4+TmYv/oZUm8zf+nKV3ZG3xLq8m9ckM5sGjl45NhHZsVe1Gzz
x+udG2jYh8N10/WEFF6ONKa7oEJWa2XStDAlnzho8XWZbWrzQNKYGRB0aZfFm1HLpg7PNW1FrZCz
56/roRTtXjgVVkCEJBNO0wblf/Qj5PytSW0SIptaaxDkRicdYUAUF9WtLN5o3YSKW+cYy3PbPM4F
EkMX7a27oN4kUdCT97dlrec0RvIzKLYW7mE3CjMTmuST60WGjnWDYEfQ8lJVD4JI4olG75CO8mpR
AkQshfvPW8mfYnX/XoUXY+1oWri6rHLeygq5qctEH/eWzqFy55CaYN+cWNcDDaN5+2PluVAdnwuA
OSsW+yszr6iBNVuA02M/QvBJJnB2aax4/1YOpBTlwo7HxBg3+wKmDykllCC9EgrexCI7R5om+0kz
T/zqMX3TWMlteLcMpIBQuDJKjcGpKfme8dRcagaIvIqu36gnjqTQGs51OyVpEM5rr7eiHYuzBkS9
PGW+QS6MAzjg0TdQL4nPX8p9xbzHxLxsr/xs+WrZR2mGpQ2e2eQoUvthrZCi85soGb6x/hAhjZef
+j7T4I/+Hf4gWZivSrtsQueSRKEABU4YSNphoi+N2Bxv0dHQPPdQFj1RzE9i04sV/YjIN03wufiL
XnbegJgHyIxrjwO6rVq8Pc+jXRnyVNFDkhRGSwf4bNIXa2o/odQoa/v1WJeeaAQ1JWvDGHf5iCQE
G5WCYnr6030LhpUY1HwHDMI0z74r8Kz5m1IMkguiTQ2wFPoyCK5T2wDRBuRMOBGdmk1RILSNaCTQ
ejLoKBM/dG0fI+USF3oFdFNsGsHy9i5bs4N9PltKuDf7xoJIa2dC2LsCFqTFiHFQVDjppFKpZmih
H9UEfQUhq11c22f6ShtDShmpoZ8iyxY/rkFBGVV7Lp+peKYM6oF54+UAN0OokFjRDFjX05F9G49o
I9iFjevJng3QWnmJBatwYGqxLB0A8+LH7b++rp5dRexDntJg34ZpEa7UL+RgsVnRIx/00lL76m4V
5ST+krHW28psI8yM5lwAmCqGy8DyezhtzG/Va3vDDVKGYIFsInlD9wEXz3m6bddWUuRlgDV2PNug
0oneg6J2NPZVaz0MlxBaV8AXRqeC22HNxWr1/omPsmDYNaV/yyvXpJWmlpoffPhDn/qNuw64I5ZR
7IkQ35yaw/3I+Y9VrAgaS+mgvgiAQvAG3+SFZ3B4qZbfLi7UnGbUkd44dZsS4V3atb3+DktiOeyU
dR54aZXWwk6CP+FS8PAAtAET+myQXK+xW1qmt3Ek5JIkXm8hsfsl0g1ipodR7VSJrXyIWFba3cuN
ziObOkewfmOboXNn1F93nHEjhWlAsv5/jAP1cdSBymDLuDigYXvoELNIlleKjGEsPBtH+31x4KJh
GWVtmR2xghWz6DE/NsklW0KxrKj5RTtuQBKB88tj9VT+E08bblK/ZeMKi08v7XU/fZ8yFprRH2JJ
3Jc2XOgU90b98PvG8xPYHL7vEiYXiOAYJ/sIBs5AoRtzR/ue8fsltkJk1Vc16ompxW97kF9RoLz0
7QuOOgicUqTq/YbaSq1kJmk+MXjV7Q9Z77Y19h7fWm1AZ4mDJHQJ0Yr2BBLsxRBlaORY5C6c0ldM
wBEddgnofuGWasJSHp2gXCWSG0Fw8dGajzXDk7f8kSe/glMctkEen7G2ZmAKJb0sDFcQXUVettiN
lAb1ulm69QLQLBQGqB6k7O5cIQ53V+fVZMgTlsD+Cbhie5OMMaxTBE7IjOUmQhVYFiSuZSblNBuO
OfJVkF7iy3Jp7XH08XXJig4KSUmiaOXhR5kgQQJvGEOJzRAjtkF2bnZsnl5byd/KntsAn4u1NgsU
ca0Pq2JX1XjPAr4SlKqvR/eHDxn44eKCbRTc5AyWAduw5Pp4mfr3GLzkPCI6rIfhTNBK7Wk3/Dpp
YZB43eM/4d2rPFY7w/3w6bPu8UXoJdKFvTuyAfxv+4ZwHsNlJV8UiB2EwhVa20acFlZl8HIfHkdk
kJJWuKcdFaWHzLUtnteiPFD+UHrhXwJ9/63AIkY4o/SSMfddvFbADByoHJJZp30E1duYwjgZwZxV
WxupJhdYn1xijQykkJErW7jlmy8fABKt7m6DY+Kuh+fSUfWIBS0UAeFv8pDtc484GKZ61w8Y2Wtx
OI2tJjqzQjjgRpbsTKtCuYY0xa7ZITyuORz5/LGaqqqMCwYjXhFzambi92OJfPi/pWiGE2TLfOSs
ZZ3inFG/ysna5K6xxvypdUg/6emh4JZw0g9Yl3Ai+KgCKRbGNPW2sFbrpPAj+V7oChBcfiocO3id
E6qPmaiRAQU/im1R5Q40+IjSOOcsVeaDPxepE7CDTBdPRDoa8y/DQaVB01u7h9vv/hvz4kTS+Q6Z
MECKmLilvpX+mlWtIIIVfMw3Sf/Rlt/goj3lTxch2e0Nx7qIObrQikIuURB2zJsmKY1zBcYN7uiO
TEmenxUT/mu2GSYOq7AMlceZTBFCsTl6CtZ3Qq5m1Fif1AeU3Cqz64U3J6EsbrDVuCbh6sKwHtiv
k95MR4trAN/QF1F+esJya7iNqyVu+2Alqa1N7J29dZWxPZLimCrUS5mO8V0esYCsgnipt3iMUw/O
JX4b3iwZmELm9WpnG1bmEebKSveomovcf51I67qChJuDY9HrnT9e+8SHYNGwmoC194zXZsPBSIpE
6l/BA+Z++GNWAnxzMHibVy2Y1LnduY3NOzndYETPeLniolkqpcg6ZwhwTxA6VFJV2xKlN/Z75xRl
sTaOcxEudfmAeBzEZdkwYOKmTZCYr070iTUtMC6egupOEwJzZZikRtBeGZaUH1bhfID6g+njvOEK
F/eUV0FmsAQtMqLuFF2/Cpk8UFgTGA1hn5H/hqWBHWkfAl2+Af3v7PQJ6KkPtge06jNFY9YMJMJV
Q/9d6ICTYxEUCjkCj9YJSOQItEtJhVBV++GMJNiOtyKgexecyUfVcbt/YLXSV8l19L5aYLDgzRbr
AaXhwscDFNpFvcFJ2L7EMBlf3a5ow+hG9tJQYkjyZRnnAo4lj7pe8wMvNW/fyKydQdvybO24G5I6
aBQLH8IZZu4zW9sGpl0CJzffZ6mbUDTet9RGff/rcfpYCp2DxxAFvEq+vBCdTZkeNWtKJeBPWlhu
v4F2MtVKMr98vKHr+jw9autsupweW9ss7tncolRM+GRxe3m2Bg0/WDgoOCoSWLadaheAoxd5KYRY
ahkZEiJute2h+aj0DnVg9WCI1t/TEdSuw8pbNkD672fP2zY5LVWl1g19DgAYMU7cxtZf2owsXW/V
jQWNwyGNBguXuduLRTJCObDzVrSoik5O92tN/658hBtvxojvMJPe8bqqEm+/TzfxYm+pdCTZMNu0
ht/cM7kTpuuXJq29xH3vicXSVVmmFq9fs8wnvYcAfShJDL8jbdUoo1WzyiJlOJASXTJLPfUtpU/q
yY/keO+fdpUtyttcURISNXc880RR4VRfx4uIpTwzeBOALeaA9jHMXGAuxuZVYr6YhV76mmUcY8j9
GQR8qyNjrIN40WrcHJa3BbxxpJJNxW4rRyaJIplBoqXR0TMoO6YOEIEPxkLBDGH57Vem6Dsm3ULt
GK52IV51ts8/yTAQclJSUUZYcgW8V5aVYotXenk6/L+AWLsadJ8HbZVykpHX4dnHpa96xwVygtPL
zMgjKNdXU/fpq541JaW4fyxo/6A479lHNIHu8Xmu2JJWOxbo/+KtJs0TT/qucr0WfzSYaKGxFoKD
uq1GEXLio3w7gbGpAxux+SGWW9T621b5Mqngi/l0PXtEr/Ms91OLYEY1AFwoY3WPX/bNUZC4NcLK
nN+gGbnMpPwyO1pDIxjU+Td4pdDvJ3wFOZuoeNw1N5l2beSrMkrgzHBN4Cn8v3qy2Ymn2xTWOMcg
J+Amajc7xJAUPt23ojZSZaJL3nf0Nigrc19OZmcujHha+EIThQOZ2p0j3V17FTw4vYkGc2uKflSk
TPo/ji0iXNRtxvdH3RT1mkCGBO+2xqnzgFOPBRShGxbknuWgoHBF47ndoMEN6oiOYb6c/8LL8nw+
NJWJigr+jHESDmEYck6eIMF8xC7diIEo4SBA1RYSPxZRa0Lamr0+u5KwhU+VzaKQGXKOS6l2fEHd
KxCYFjx2q8uvyzdxqDRVItry6Tv1IzN3ztxqLXIwy2S3IknYwEIx4AH5urobD6+4A8/1FeOToNVV
ZTR1QiRClTIGmoIlR9zAYTPMWiEHq/GooHAYleQYHQo4YjLnjPZoEDpA8MLVPFMTes/CfPYC8CvS
3xZsmPXC5ovTVwimAEAm5hxnUJaLs5+6qBiqKL74CkfRa+24QNtAFZjzuA7Dxzfna78cNRC9eG7+
PBXblpigXHgiLlccaTBy0q5U9V+fb+p3MdwzplVyvNbBLKETRDnR6Gni00h8KjbfAE4mKZQH7l1G
I3yeDAxK/xSpiBML6VLvzD0N24sJpnC+ykq27/xMfs2Ia4AYxKdydaP+JuFdaU6O93DSBq0ecnGj
2/7C7mwb38ENB/ALq4z4QZg3F/5KwQJFAwMWbx8LKmF5HAqMH83LxWbYTkTcu+3IWU9tKgvpuaGy
sGaJMp9v6BoKPBoynT0BtpIEVdTUJdLeg/GhAZU8fFPP/CuM9mfiw7hkgAWhOLBNiiPu8iNaW7zz
uHSbDWzIrdZpH9hWj5c2Z/79Hjd+Aq4L0GrtCI1tAsRSFvylBr14rhexvbtD0BSMSNfG/JElBcEj
xZV0mLJ7AGz96Q/AkqNqABylElt1LFLhp7uMIgV+bkwn6c4N9hMLep7mMQAH9erEgAcN4FbcNTmU
Wa39V89aCiDwamTmBUbNSRcBzp1em+VHebJXbsT+i7bCPILKPJBTc13XXCg723CmfTzjxtkk95pK
O80xb9CY2nafpn+CIIiHW4IwT7f7MK/9Kbfw+EZC1lVaIaLKS+2x/r4zB+OCuDQOeB1J0FDhrIzU
OhZWDtcMvCONDxY4r4jSSAAIJPo1+NEskThmx6f9G28r+kytXwhCdCXx75pB5qw2/GKKKruVMBu0
kWH6SdjEmYPp7pA8/FDVqfT2oZn+EcLCKGtdxLcXvGedc6G6s+7H/sFo7HryFQHPwJSp8tS4KyDO
Kjt+Wo4kGEYcBLWA17wID93MKds+/1loPNKM7klIYxuRufvCxDgdrIgi/jGF1Uoiwj19occLpn7y
RIrCSJ3r8JZa3VikYOHzENvJACoEja1jvR5O5kmfXC5oG4czqpuuumG4DMBcPHtnSgOmmPhoYqNl
lyitIntXj+b4MlDBYF2KnwwUoOLeKd67n4yXgYumED3RG+OEItRupGxAu7SSeiK+0xnbCpq1EM1o
YMA1g4TyCZ5V57Ex92S7Cktwy60pquoPpFum3GJulPp6gqsX4ZyY1BBT3zynMx5unKmm4bi99msR
DPSyeH4iEGTmvSkur0sKG4J8B/TtZ1LV+eaz3qAjvPFnzNkU0AUeoBC3atEXWvwHKuy2Hm4F2R3j
qfXqAiY/hIXCB5Pm3de1R5/wAw0+sPlHcXW659lhdMIXf4E8wSx1VK3kMxfD1gFVub9ngyR6j9gT
/1HiWQ1D3xjpuWAw+uGuj4N/0jMyKhBw8hm5OXhP1kJFqqnbaRRBvj4NEgmh1Ln2nziPBmIwHwwV
WInSj53+C7V7K52BmyRALRPx3CnsdbujtDYt9SWOd+3K/0hK+AUbJEizSTQAjuGQbi5oX+hDj5P7
BUiPx1/LLHRDFTP257v6AZ7BjpT7jxJ8Sj11h5X0RutWMMHILEzICU39lQpwjwX3WunbR+2x2CWT
5dOBm+Klnucn8BL9+XAW9MLTISrQYfx4oET+AExcbqXOj+zF1CB6ZVpmr68h/L1xdTuuxQPKgsQe
EYmRK0kFEub6Nq+KMx9aT/ntEUnm5hwLtVXdEXwlwxHdwEE0hH4+mq7zQNUlE+QMb8Fm1vMyE/2J
kVMx1SPyWAZno+5zd1cl7Bh0OTARLydR9xjUnnBzabu2tCnyQfFc9WNkMjRP2IBlbkMTrIHAc+wq
i+71x0iF26T2Q10FwjJussB2ajiAv61lcClOQs6UQ1D7DyPUCKnLTD8MfxTS6hHp7hCZMUcda1HC
1o0sUrhAf9vxCQEFOHi0njBmujJj74WB9hD65+nzyP7n7swnz0et7Ug1e3zxc2axyZRra0CKwQ/A
+4GqC+e00QEBSEf9wQ9GMTfyw/cyufJK/g6Nfg1Z/XBiCBIc1pXIJ23Hjsw8/ltfyDMkd1FM8dGm
aeIVKsy+mXACtjnWquAt82itOqB6lQo4V9x86kReoC9GMCUe3LY2zDMuYEN1Qb4eslNJfCaJbUzw
vzX40x99nHP3i8ZmhwIyvl3BNWmu1vTuAXR0TJfz+afdBMbqJCPD++LBt4282woIbcTO5se0j7jT
duD8vtXcTvmijacejcEJJ5jprts5qpKzw/BJ5eIMoNcEbHNI9ox6iJ86wXcR5q71FhGpzL7KMih7
pAJfpw8yUED2BEKM8117dxh16XY8/NCbSSp50l6Doj5/QRhKRp3+ys+hgwZo072m/rFs3djC5M6E
koFCfb2INUHcjMNVwV6bnXFHhv7d8OT5IiDcHXKAxtt5OxDwHRNJimiQ7q/cKV/CGrzspge0EYPw
9WlyciFxpbiMnEbwPHzYlL2ujTBNBiwTBg6lB45PEoT/F/K37SBpC9RtizILMogO4OZSgV2aLq67
SQwJC4yypB9ILIUHF6or/r87WZqz0Z0n20bAqh8UDLTq6CV872QGrxibZ7uE7FEDp7gybo2Dk2ci
Ym9HlDJR+fBiBsSCWtLyPZKtzoQJz72r6ktudzkl1dMpv4m1BaSs4cA7L44lhW4JEcabEJirba2z
3Nn1YqVN+nuAhnHWLbkTAdNmTGyr0IqRxY8T/CmDy8oifb+ZzYM9KzsAoZ6mI1xhPdcDI9W/9yPT
W89QBjXyjp1ernCmUEMUofqmuC5pbSPQ556JdWXlAdL7zwaIMLe52M0mlWpnxEoazkEOOJWmk968
QFW8kfrW83AiEjFnnCJbKeKSsp0PqRZ6kMv6+Bc/tY0eOqv9tfRqBDq/opjucs0nzDtbxJhNVLOP
9vEdOCNc8N14XuJu14CejA5k2Swan10Fv4mP/3pNLRGxbqKCXEura4tQvQwgRgKckS5bZg0lpgS7
5guaMkJjiDEPr+8GOEr431ZI9If7mCFBJRAy0Q4sl6qVfAjSYrzVLwG3RZmVA5NIG0Sy0uDzC87M
kBdfAnL+zpTcKKa2b1+SYIL139qeGwDUXp9e0rPiPeofRzb3TEH//RhTp+lLKWVGguYAVguzpbHZ
4SFYalmWh/6RsUIHBzdGv71PixAPYnLjLuhjXIogoDwmzpDblxUztV8wWcNBNMC59vSqDSD6+zbK
P5mvWDtkZiXf7QxICkhxFwdyN2etFqFbIfIUNWlbcvvcZaDU+tHXfPDnh3RU3q9C62Vv0IcD9NrI
6ndyea6chJMGvYDSr8JhQ6jxdJRaXyGoDUV4nJQ9razpDsjNTg6T+B9DFOkBRUolh0wOD5EINHQV
BnzYxOyZlKAkh1M+QYludCFyBiIuRysuSqoPxu1aCN9TUXYljxSFv9EMxK53NAf/OSv0RXAN02S8
tpIHy3n1oMaAy/o3jgamQ+bES5Ok/K9UnHa+HmyRdVdqq+7DqWeikT1e+6sG9JSX0ZmqbvZdqwiy
lR8iyn6TZanFlq1s4cKfcTlxS9/tp9yKJWFsPx2YLrJVLbcZyKrEW6Qr7ylCqgf5eJxw/tUdNE6q
FEyHQ2GlW3K/v5bnnO+MKnROVgZJuvYvlePTXUR/JEfNSSHqpIHCS+oYYNve9ZisDJzQqF741HfD
TyRcfmK20p4u84nTbGna8+1ugYSj3aKlHv5+YfjArFIEdPMTAWzZiCa8NnOH4wcDcKwuYm/gr2pD
99jn59fuCm4KLjfI3z/Zxg1M4T+6muuxCMbnvaSmoIIxDgeiw34nehAu8Art5zahV2RMiCAC0dpV
pQGQDpyEP/xoNeUhM/nc1vzo5sDNiDTnikUMY5NqcDSU2Ub3h6Vga9TnEQEuk9cv55pyfbuh14/G
UhMfJaU//MmyBnZd02ObGCqooQclDgjDj31fJwTaKGxm5fkehDP99o5RkeSd32dpG9XnAblZayna
7E+La/eA+ynGZ4HBUq7bl7MTHFV2/ods6vQYsAvsuIx5D4uDbT5HCRRoV4jH3kI0E2dD8lt3P1BR
17eD8RM4MgDywPrRPD9InXEJWSIAwx2J2AIhOATXna7i9tqiyb4wMIRBBrevmhah1KhJosTOg7Zt
s0FBy3ExbOE1FohZEu6L1/rGtf2GijoEYiIOxS0F2sufHTiMVI9wrVoWuGsQ/yeZf5j+AZF32gSL
4uuQMv9BozGKuqbCAFoey503Bx7QKTsqQ/G5AYLFe/mCMBxilFXH/k+fzYnJVpzxnjxpisRRsivB
+DgLcWLhXMXNVNfHgrDF+12rtikA1/Y9z+vUHsxp/+zXv48NX3meThnZThsiNlYc4UfApK14HN27
L3KkBmyx0ZP7lapBXxPJnSRDH5IeOfHUS9I90YCjKQqAp8x7QcfJGcFThfyNu45OxYNXL6pOBmKd
67nOULVZsDfD3DzdhEGm/ZTjwl52xxXu8ld8342FJX+Z6jKVnD2eRD5gfVGBhKbDRWdud+N+VNRk
VN0rKUWmC6tG2X3myYKmMkhFNEncj5IijBRKxr8byINYRk7MGS1sQguylh3aCUUVKCGDeBjOIHw6
dTEP9jlCFEkvHeySBZcoKnuU8Y9WtnKRf87mvY8M+wNgNksndJ+/nz/gqjW38YqSlmh2MlytrME5
HGyxEpUxtk5ui3GcuBcdT11O0bN7Flac97ExxiWi1GCZagAwpGGSZfEqsGbfjC2doA4bs2s7HjNp
hqDgh+JvNGAe0vQqxp8XAotZARWEZ264HmtyBHb7NM9HEq4wMMO/EWb0wykuMPsm6BCO5vwBhIwG
RoDFvKgGjcUXLtUQ/FyWXiT9vl72F+N69NsHifGyKb8CYiYEG69x4Rpt0MSceO66/3pac8HHkK9g
ZuTrd3b1b7BwqqiUzp8R0qIAhXEIZXIRcYFMY7ywkjly9MwUUEXVQW5kJQ2CFovavUB09z5834Ns
KDvMP9gImtGn0/Ub4x7q/bfh6nf8M6GDITdmhDsWS1FqOoCM2fD5UI/l9Q/pmQsvQDjEQ3SUwmZx
D6EelG15Ww9qwer0DonWsKhy80s7R2WbwdOcYIQqamAOO0GvsNMpWxHoCNSBLZ+3Zc7udqICf3C9
GSercU1TXARsUDQXrRGj0gDt6jphEUGGAXysQowi/xw9w6fYLQf4xU2AIuCkG7RSpKz0yBUTwh7l
dkGVp1zclYUfTOEXYvb/Kbq2QkE1iivYjUYGK/WnOkzjOHHR5jswVfiebBYF9ukcQj7UPHnE/PKE
j7Inxc6GqjahqvzNV3u9GtU9HKgLi5KB8B/YneV53hsiLQVoje6CHnHOxvXFtLlgNjsTQj69QvCf
Wp79549OOwbgjNR/wj7WpSFZgYYKIfDPTH9dh0/GGFw7ArrWWjnyuJPYFV+jjtmp7k3alwgzu1V6
DBbDMEklgYq1Dh0Q2OHoR9sNpnMZO0X3dsWWrgm2Ty+D9uxFhtz5vjuF7l4xTa4uADSDemQhKa0h
w9aEzNfosWSN1ka0cNZ918RBH/m91rSgqse6ygqqljKRU08RNccfU9fTbp4nq+Kc/czV2E5tteox
rDUgGbpRfN1eAXI4UAbZNyAkuEcpwsCPnJndmJr6DVn7bFDnrVrbORytcphqDcXTok7fERBXpcp3
1YgglNmyOLhVH5e0qYjejaeykuWfdnWgMpJ+AKYBDdcRIjlQlmrTmbYBQ2oXlyTi94eza+9/5xld
iSxnMnc4WfAKSRihtzOHBBrozY+hQgXD4s3gG976jFQ64/+cEvUE3wNeBUbYdxQe8Zx5XDnI4eLe
1GSXvAwLIALzutMb59X+C5AMAgxHxS0p8qJiDYIChRrkH5Aev9lE7mMMjOuzGW9i4ybx7Z2Hpo8y
lKXRPyTmetW0sLwmFEQCc9kx/RsclMCGkNAmEa047ykV9BjbFTQS/khWrR82fesz85El2jckiSGB
fOXQYOf/+MnvVqoW75WXPtsePUqp/mzcrM+9Y6FBqZzZiLSQb1+/jXdQwSZQwsJup8ox/LixwzP0
7YdOIbiRSNJbyDwRhnF9oWPYCU//tUPcNYGaJ5z1dY+Su9b+tBKvLA8/ugjAe0on+xJr4UZWFR//
XJmk2EK1dwd5hlm0Abn+1ocxhKakatd93uwpTazYtE2ESSxgiACJmUB1gFasRQrSr75HZv0VwfZm
IVpiCtZmWhFA22U0U03ILsnWehJld0XigGVMaqwFoJXdK7+wsQgWZyCog6S85VXq4WAyx12pYBvX
MsuuHLJRVjnu88npC4/iudYvO7+1Ib1H87tLwFa4gluQLshPeq/FGq3LrCftfUq57DNVHoMXBUOD
AgNDThOgExHSZenDTTs9WSbSwvB0z5opNr6LDZo9WYxOja2oatv9gRnVLLKKOGjY9MK6EpNpnRUi
/kngOCygkxn/ipsMqL4cySLjv61DBdOAgBZIE8eAkVQKM1wgfvNZUoY2qNL7tZQgpctnxDjILQNn
VZdH5d5JdpmpPwyIyqVvBCRdDJXSeaqcAh9g+NVdVZOtdQuMS02+u6k4kshNh7Kzminw8FCtiroi
AIby23OG10EdeOLQqU2w4PNStPLg3H4sLvi+QlfgoUYuEx+jJUyK2E7QM0iRkwHZAzMIdj76gU1l
AvEbR4AcYg00dVezXEBq7AvoRb85cccusJyvWLxkl7kZicBGPSYeBpIvzpIDDPE5MTHNAsJLVRdW
yxR2VpBbEkLXHHPn93qoBX9AlKhh8cbJyikYvI/fxvKUgfZ60GvLr185uVV/K3hyQQNOsDOLY0e2
jiIWF0EWxEoF09Q9lsjVOQoJ9MI8hzn2zyeH56RkAYVISzgoSikuZE9otCEewKQk4ZBqkcZ3WNC8
Sj0HJgtYe+fUq/PYC0/iOaFHn+wIvt7bj+UjIBU1xPQyWmOSoCJHqNlRA5lrHJt6ehx6UxtG4CLu
5uBb/Rckl/rpjlssGoASUVpWWcHMPoXQ8gdIqGUUl9XMjfDzY38FkZOa8+PMzcqYsvmMeTN3nkyE
g8nB5okZdpXmoTPGf/soe16gVQ7CT/mb5lXswFppK3r7pPDxHc0ea/WFf4JwbRdXLnE6rFOpOy5u
vB73HZVNjLcMDJdIuGMAxNplRmPD3tVJ0xHZXFoSkR7aadxyEk4oVGTBSbsrgvGULokUA8t7TeHf
+ukBk1cj8PfIZ+2/ovUJ5E8mVsNQdxUWz6+8PHmuCEVsuHlkqrI6codmighDRu/a8pRPSvmhfQfi
gE6r7hdBZjUL+W7yk2XQdl9yveYZM9QCtBOPF7ro3d66VDEwse6hiZGU4TNMruIFcbNXuPAc1RYF
pAWa4NSBBhLcAgGFpeDOLEyTllX7s94mboIgKayUUwtcncreCsdNaPW6hU3m81WGwXvqv+I4IACq
nZT/p+jQRQmPHwvr6m4vG9pf6y5hhPwGGErBZ8GntggTXWMJmYeCvsEwT5t+wwoWZFUJslsA7Na5
zoBxNobbnCxQkqDSboFTb69DY6/AoubmKH/iJkEV3H2OYHIdMlhtaeVOP/SWhgxrytYufrLaIhZt
do2401RKF4cfAlh/a73Sfx+ntvipXP/w4peeoORbkUsWlZ5zZRM4STQW4kTH3iPH46s3ivqoTmBx
GRdmX10SERWUSHOOIPkdLeQQzn7qGWggoVXa2/Rop8A52vaCpJ5Ti4flsp5LnR8BtuhyJ5VqG81f
KN/lsQ+OCU/adldS082u5JmiRbySKQOSkmJK8cJr6CfJDqaM2jhU7DhpZaEx2d4elJ1ujKTozM4H
TeuBJXOWPck+fX4rNQ4BESs2VFwJXr7QHXiK9XtyE6YCVVUyNHtfha+QDLGBmBlh4AMFMDKPPCH9
x33XUDqem3K6ad7bJMEPmv5nQRypf/CgcupOYYhzpQRP7D+S1JOiHPnv8A6K+eFXmbi/wV4cC0kD
S+A0lzdIPOAP7RZxB3igXt/goHAOVKjVUnV5fvM4EXtWb7Kc8ojT0i+FLByvh1waryGPD99kBYoU
NBYJYpShhirdfjIevwFQ3B0lOIak+aPAcxg5PvvUiRWZUgdjVewGucw/fj+bSuK1spgueFXEF/Vv
cp5rGjBkwQPT88RVrp6L8NKEdItBIh8gtfyaIaAkrjhyLEjUjbAzCki5mEaEMcXEX/1w8rsRKijQ
CN5esO4ZdgA+X4ockqyzRSy8pHHZREzJmFEL4WMZzop8PsyJ1WCBMyf/sRSrEQRCbUU4OMbgYPUu
WGpasPiMy3hk42c5AqYcf/Z8jKBsb7lbsFtyBRFLEKG7H72HkDqjqn3W7010dHyFdwlwmq2EM0eK
ErDHcUfwVFamkcP64Gau+hz0W07/Ysu8hyCoPeQETNEwgQymVrSKuzfRvYWnY7/J+WA/6UabZyTh
Vs/2AEgxzCNfWGcLvIL0yu2P8mo4EgRGZcH+1RVgFgZLnT9o3HeJkH1HjlESFDtWCTMNKhPB3xaP
lWV8YnLir9TMF0kbXEscIfyaHRQIbZUBR3JGLB+F5sVeCJoQQm6LpNTqugXv/4c9drfNA0gwFD43
SAtY6jGHapCYZkP45UCcQuFM5DwjNsXsfiwF4o88b7XtuoXSvuIloaPn1i+9DEY79sj4j9ZvemaD
cZM8PBur6bWv1nElUf3JN71mCFDzlxMFS9Lryxzo46dQEdhlQ9rZgtMv6gSmIHyF1ZAaLm0rbcIE
6xIXFDxqaRAfBBta2mRSAgapxgc0ziQABHiJxgqBvFgVVpCVH+p2zUCfxmpGbvEFsQQ4bcJhr3EO
sRD+I03NNPmitrQP9iI+qK/rhWnHVmA3fjF77k/0l3nn6vUllWfRU+4CWKLw9J4nw10/bDHAhL5H
S9dnhkeG06BSoTQcWQAc1UV/Ejtur79VIdMBcWYtc4KRTMj624gEWNt2l12QIv/rrGih9uVO7NR8
u0m0lWi9urvFMzdUUGMd89D0zm15gy/4n1GDx2ggdUGMrlOrtdP9QFZuNsHu5DJjAyj7a2gzU4Hy
kgXkeLVdVEJ6j+bAKngLHR2i8VopcsdG3pcCJzhi87g9pX7K7ly0LBbMqkH4NzvkgPkyfbIkl7ZF
hVqv4SiunhVXdT1ASdKreSCumD1vepN0Dg+4si234lP42II36FWt6OMQno5/fVh4HB9b/ApdmRU+
2a+Wy9BxSt7pyGNVS+N/pUKrwHVQR84zIkyuj/ARIgQslKazOJoBP+uHodk+fs6YeywyJYjFPkyk
zKByj9jCXMJUqKfGCMkY9biri8emDjlgoJfomxo96yoxtsuNKdRoQL7XP4kXnookLdM56BL3crSg
/jYNtssDEhDDyl1V8ryndVUOy935jnu5or5Z5tn0y9qwE2FmpRqkFKTzRJDQ4+9+YQjh6zOl/njQ
LJd9HWsK96S+q6bKP07fYb5h1SULTmqJFyomYJ44hmmiOf2sLVh8qHYrv0b6xfkoJibpM9IBUm7L
cyACrKYA5Cwp/aRe15GU2Qm5DCqVVJ57K4Hj9AFB9ny8yKsDN95j7YpjlCU/4MiHfVlaezhmJObS
cDJWwYwptarCKqMlY3j2zVHzfM1WJYBT+bLOdMlpRH3/Ec51jD8uQb0rbnDoRwDUGUItN5v/ZUiL
i4+pONCthmVTAssB8Cawd+4EXJgEmBIMhS7rlAAy3RWy9ou5V7/MS1neuMRIarAD/PdFhaljAYn2
xeeZHpP63GO1QqCQvlN7V6Kmtim3K3fl14HfXzfXNQ4rCodt+tJPbShqm657ySRXSJqU7VHXih5a
cJT68uAQI26VXA8qkjE3fJk9OhArlLYOYTDr10gLPNF7tmp2lxMYwm3UYDDJuEGCSjyFKeLLs2Xc
Ky8CAgvqA/gdbRbxJsFpxOh7yddT6gs5K2kjZgCQ9+hfG8cQ7U7O7P3BEUJH+LN1hUUWtSQCVVs8
ZXJdeapTtfpq1625YHU6qRPwGfCgODYY5sdyCqpgutLITKj1KDKShaQvW/t9Dn1UmrUE9ZkZdGpj
4z4y61IAbfMJSkzk7j3mQZW7m1g0B2R26SGzQgPHitfxZ2MIDyUwkIn+ES1mGj+0gqj+ckqsbL7t
V91nAG0070AzDcnncpD+AELt0vWidAWCo0yovdEkW1CXv86kLMU7SldSMjkrwWebcTPOj8tzyJPd
NIjMOlXakjAjU1apjnjbQN9aAQ6HHHmqtRNkZlN5VstVlDr2IMo83jMj39sqvw08SJ9NgzKhRXWk
0NnM7u61r+/FXwQf+M1n1DL8dUYcfJjHgZW9ourFJeOutkC4KaHFgxu5IdZKTc2+1iw7UFfoXZRZ
v3wUKFFjnJ2ZKlOdemtIx3j+feMIFhjAS3quW1cdsSeMz4GmA6nUx7oB+UJ5Jg5IHZp4eNrNRacx
VstP+kcsYwxXAzUhhN5yczhdv48mRkJHStfGexFeJBO33SWUVFpKpIQn/l4HgIc+NTMcgqTFnbVS
FbmtfqrK3mTmW44JEiAeguMxMDoqm9d3KFS6cijZtC8erIojUv22lQb5fLMPeykepipexmCr8Q0L
RiOhzKONMzQAGK3pQ6MQ7vLeJcGPRt6RM+pxacfNST6v9zJQizRg3HmELflThSrE3ALhqRg6mvsG
uXuPfB+8PljK4+LGKKIie/SODOUpdsOKu88i8sn97wHR3Zv6xmZXIa7bIgvwSRxEdm4WqYkDyJSO
T2M8GY2ADenycsd6URyLhCJ5jWaZYgF9WH3VkimM6KYstxemaQ3TexxBz7SukHXZE+TEU6J48rhh
307ghDgv/EJQBdZQM67uGdKapgQb+aKTtk0gN4IixG3SiCVfcaMdy+xj7ozkkUuRHOm16mXPJ7RI
qAdTks1O1l/aVdZfLUlFL7KVvWi8HvmGXc1w+hYcQvuyxSMlIqpJmxfBZAa2ALuaCakdEj180Hzk
xgex/83DSeEMRprp5335kFtcuJwQtf3M7TarvZ8t6ci59djl1JnKd6o4xu/Y73W1CDyp7hIyEgQK
seg2HrRDa7Cv11FvI16+9NNPzi9GbmhtlKR31Z+ds4CL/2vDfvi0ikGuvXkc9nWctxvZCfhnGozo
eFAXTm8TyIahRX59/i9483WEYwhq6cRPmtwAeEtv3IYMsm/gGJWKuOhtgi1VopySSB74NjO3Rt+8
nS/hM7JWgK/yLoA6L7xgtnaEHUump8Di36lvRfiW7eU7y83pJ2yYrciKhaiDbtuFn8onIj3u0n1O
OgpLDyDqwxR7Z/xKVerqIpU9P3TG6D2Ywtmp94iE15D7LvKMgiYmBgzzZyNTCDVIl3sqRhw2EH5f
lYtrZqgqlWZExjNDZ9EWtWbuENPwVNt67bHnG2RlFnAgUbqidpW3C5wBzlbsI5xIDGeVyLwiT36X
mWEdUnu6NMAlcdfPH18yPl2YWb3nOm3e5ODkDtXZ4ttK3fOpY0Sm7ri3xVOXa/xyubgPUaEDSZHS
N8eELg3H09SH0MD+bTtDthF8kGZ9DzWHI8UdkhKzq82Vw/jqB2J7Z+qNy9IsGrzODt3C9msXt0un
Sp/wsKvKlNd8HJUYhQGE/6wwxgONGprYuBXncGTa7q/OltvJELBzuEOXi6Y2XvYy6cYxtI9b0FmR
EYk9uIxilkB7Kpft6iW0Bvm40Y9Rkf89QOU3tWVb6fCH7W93cheAJKfsU+ZaztwjQNZnPOfuiY7F
Kvf1XrKcEkxBGP4PrF2Jd6c07TOdjyEgy5OeI8dyJvWidb8SB6tUK4wZS5VfvEKvgrYBxiTWcn2r
aA9y/lyjm2+ahDHvrJ/2NIqtMm4/iEjKR5yUdBW+Z8rDpB0O0M0NyojlzXFS0dbFb8n4hdCbUd+m
aLEmeyMI1VJ0DrbFks3lL4c52VMKnIGZT3Prw7hN5Jr3/wvaPquumHmpae/9tEEsS74rxmqUEtd1
ve3GDD0FfaJBlmAhUec7VX59DfHx2O+/0hoTBAf/CuMcom+/t0NS3I6zJLBNgwauWk3xHoAN1OuK
SBpVxQR5oBgBDltMt7lzxP0QX1OXifJJ8TIU3qfMDUTLZzRhbGLYrsvZNzA8drcVrCC6wqEnsz0y
jHLcRe7LMra1h5AT1Gc9kMgujlb+RcI+PC5v/1IEecsI0c7DSbHXtznasu887uBVIxFCyGuuLUgO
NlPKVe/Ij+EqERULrrl30o/7uewMKt29wcV89g/kvsut6SEvreZdRLRcjnEOpHzmy36hVD1CoAlA
J8lZqDlyVk704L1G7qV7wuJTRnFxTMY9SHuNxNgsOzW626EWjxU6G6fhSQQ3dvgh8srY2+0g4ikN
nL9PMgceJJPRkJkSZ7nNKzFyOLORuRDD0lh6OM6YjB5iyrMYBhd+nj7AxlI6K6G2UjfPi2YyxGyG
0f3I/e5POFY85x+h9L5NS4Gg6cUUV9/zDMooaZ4bjw0nhOdGqYWOXY4vF+ylneyEtFlEV/EZS8k7
spttLzp+O29+G1rhW8vVVgYpStGGCghWpaItjgBcrD4ZiZnfhx0Fm+qcWw4ZkVpTSFAWNdI1vxSj
CBjZlCpQSjQZkilsdMGcKVpRaVH89GtcwUF+t3jvvocQ24uxX2HP0gkRRDdy7SVAAAcagC21Z6D+
3O9Vi5Z3TeLg2PidLqv3VU0yTBa7pfz6Xj4/5YWCRfG/y/WpuZnhvuwGmxlU4/K+cds+VhuG/c5p
lS4RySwjH9q9xealsVaJTGNNB6bV/8ohdqLothFLEFhb4HTld+DlQlUJxTI55pC2QxYZTUs/dxxu
Hf9lvSRHuGzV7s4lW9meI9NYSHVI1k4+STHaMjliP9jFe9MOu0/bghVnJjMKEQY1AK4pEJG4mPcG
7j+01OwPQHQPPc8JAs3m4dDFwYUd1Urb85O3c7OzdqIDDSaEq7X37EIx/UWcaXjpK/T5g9WWeEup
IzhSvlBaZjm5NsniBAVPUxxxZ9DXz59H96bJoQkDaNfNaGuJJQqvdTAE1dKNwLX2kgzQ1eTkZoge
u1dQilVrILcD0wrYRPjzHlUuqhin8lEpT9VfcXv163OFaStCi3bqBzbIPsQ4DHJxs/amMF3BO2SD
iU9J/p6WW5CXHyvlV9qVWmYj78GT/13un7AXUPZxRM2drvF+43Tnr3GgB0XZ7RdPXEDd4ehC1LWm
5ef9q5Zs78HaAqsf5+MOlIzohlkac7M3Wo7FvFOZ7/6yf5zKM6auy8vfErJt7QAez4QH59Hj0IDO
k4eenTycYNdYQzvn37qaKSdTSYecQ45ch9bA/oSwVBWLBEnEcjirkZJ5oiTkst9Blwz3S9DLTJ92
rf4C2iuacp5g5vt4Vf3w9hj7ThT7wrYhkq6FCD0wTLMwdNjP+bDc5Qfq3xGMq99sCFjoI00cjDYd
IUBTTfAMcT8l7KexElkxCyVbLnD0V21L/dA3BpshNJRL63wHh7IHi6rAKjJPNI34BOfI2wCgdpiQ
Kx4IfH0IDBexEfxO15AATPTSPCDH1bv9AnqEaXO0uH9zYqlDCDmnVzmtt0fjNYqeZV3+RjhNdQGr
zB229nYjqcD1iw2omO4qHCarBrTdEnIMJlq3VRAfH2C7Gvxl4tUjW2YXOs+SKK4JG/kDAa2l/Bz8
xcLJnIPaKEahuVwK8zsUtQToAkJy69ezeb4mOKHUp58/rUoFSvgOQodKiu9WAlcXbhlMIh0Ze9b+
MR9jPbOPmtQZn46YkvgcgUd488P1bCmzknvfUU9+pHuB6WWaYb0GbwAKS2U0Q5UEUdOmEizQLlo2
xqagImDAan0KnDP/GHaiRiSeycgM3XZJdHJ0ID4JR3Z92PvPLK2UmOsmQpkg54+nVqthpi/l1ZtO
yt9CaAtO6Xh7CsBNLsbhcR4hzHl4Y4Jdgq+tqvb7Ca7apOWt7Ni78CUiDHANDw56sXoI3C+YWABa
0beYpFh4HGpzm74wWTkk/akIeDBocsynjsMUSm4K6ahrQJL3IpyrweCxJVimHS6R2J2a12cyQsrh
/KwO465o7t8aRGVJ/tozDRr3PvNxqEO3wEg93E67cdFZLGS90aPF7PatkZpEreeGU6PEcDuxxvw6
9qE9iNZej+LpOPQrJVSMijdpmNZAGDFbqMLKldvZPRNT2ZlHfZNrcxz7s8R8WC7xcbgYvhyj7RaZ
CujwMvPteuD8gbk2igYb0K8QzYsamGtX/pr7UUG8JXbm8AXLKOR77SEHMSsNJE3bh4ObBhiw3BOw
KOXmOloOEzi+TK6Up6K77wdaAAQV8Ms4HyeNA6LaHO8heDLT9p7pEGLsS6xM+4PNy5z9JHd9rXSP
bHZ2pFScLdRskvvsP6vdvMVgkWOUVzHjV1TLwUq8ckztfWHyKYB+ku+QpOAhKv8A5HI6Rh7YQHVk
XvaEMFR5RG+pQqYqjm4rwljT8M1+PM1vEQhKMftx4Sab6GjuWGQfA6YECaX6kERxg1YUsvgKRPPJ
50A8LR1d6huVkBVcPAfqbQesn5c78DFo8/3csj9KTmdKscCZQxdLweN0DneTMd1Y2uPzLCmj8Ot9
jRfXX/j5+83K4N2xcYzHjgJZhcikCyA5h0AEAQsBGkt5HWr/t5e7dk3hicl3B8c9U579EdPOhIo3
mScp0OO1eyVW4QLvyGqUxgXpw5wKyziwCp1eWRmqhMIhwN1njvzHWM0esSAYTFZysxPshZhxuooN
LKFXFWDDgwA41y+qGlYfKPq8R2efqggkp7J0ljw4+HVdfF3Jgrl/HgpQ3AGHuKeBeRfEousiWUkS
KsyIfbq5AXDBz9/DbYA00iPtRdUIw95smiFB1O2EPH2+vBKZHsF72uDFhZWzoc0OREvDSUOx303Y
+6nrJjSB3YFSZbsdNmQQ+L/4sZG3tQqbwZQu/6ajRVuBjTLBd37BppGZaFnCNFjhdDOqT6lSn3Oz
kL+LFccp1QqpUAKLPfSZ4CwQ5cd0XW4IBIYzT74r2nDQZ1GPo4goSD/rcjCAqmbeWp7ac5YbnjpN
4ILH7fm9nlgI0f3NCxpI9bamuvB3jSXOAQuRr0gwA8ZcyAlPMmXzpFf6vVkRNunGERSV9MRD8Vfd
p5jVq1vFrUl8URCFGNTxxCwN8yFAfHLRzXhQd9uXepy79b4Rw0QAnu63dclCPCXaziCazDIy62za
y2x185sFRSjTAEuaCqCC9yOedC/tjaXEU4DgHKW4vQB5e2Ix2tggg1250/cVUyeVxPIcPQ3ZE2qN
RAVddqboiPSZBs/dheItmypvVHqYs0gBquQ1V8Q1K8H/B0z78k03YCFlFBRTjnX11DxME3pfmK2q
NlXadJwaMas5w0g6ASBo0kWUuSmzyLrJz3ZbNhxIWDRWb87SUZnmPMuX+4jznYdlmO0qQ6ZvLs8x
GFqWzD8KNq6u3EfXJLwGeRVLr5PmikXqmJ2DL++UT3omprgbeXasxU8G7QiVsE8EJOsZ40MfYaKH
yM6HDtXQqQSoOKODFwCGLv99Op29mj3uyhX17hylqGKq8VMfRXPbyyHuiWszyerfaVRw1c86wcfG
QbId3TEVXx7H7vXmGsB6QIpPs0ws5PoQxTmhN3+UcvP/BoCQxGoE80tMaQvGMPq4s8yR/5pzdU3N
/kBAyCztiQldo/BzAZ8SIFrV6VUKS4U1Rr3KfloGPUxZQiqhUs5QC7G9mPS8GSOTbVJqkhdMi9l2
rwIDhGst7WdF2GlFQmepvkJKvPs/W//PX+fp9dpya1Zn1jQmjunFehXEK90jPQyeALGqW5dDwLj2
yzQpV1796JEbJYw8A1WIxQW3f2PjvuJmXmf4NQwM8MX5eD4qXf8tkQixjSrj3OE0K5lN6BEHS0ZK
dGtT4ayKcfuzrzsuabpdAROIEEUtURsCYSxmCamRwIl08J4qbo+iXJuDlEh6EFJfM/fjBdBzuuPl
Liot4WU+HCxtFIrGOuj8wSAykzOGoMAXKmh6yqXA0zAH9jbWPfiar7UZLbu92a94BoCEPQD96M6G
7t57E7567aTDf2SXtVrdHWEioSZWLJK0ryejH5mw4DZV++cMTYMKpJDOnbat6fsDE+bT+xj0Ia7T
d1AeDye7XuUFNXXPyJlMaKBI6vYPZKHXpyeIoVLiC29kIRf1Zj+CUPpMw7JwHtpXKqw3eDRvlTOo
9Ek5qKErDTGVXrrrJ32EEDloZOr6XsAjNo39XdEyUjgHv5cLQJJpQDbb+P+PaS/sJ4qzC5/wIDV9
3WxI6+VCvg3IuWlXjig/OtUszvg9DMVGiQTxNjxmvQMb7g9ZWFKPO2VTQHVzXZj31qKA2QIwCPRG
KOGFsWy2Z/EzqAno1TT5n6JhdoFSszb4svPnDsBBHJ+NMAffOrdES8rIa9pRdqKeE3Bykq7JNNLI
ooqVjFfSltlRvbAoLPLuGtCAiEnDCVVUGISFpJ0BMvFiFlowTzhKtlWyCDPc4RSB57vPjDiCPoTL
U9H+EuINODon7detsV915EBYlCWu1SzRSUJoPsdPuOhph2DIxRQ6L4SIoyFTdzRQYmHu6jxSnGDt
1OgSFWZQO31dft5CSIiFVMF/BkkbBsTMGgFLeBTUkwRxMjR2o0ghaGIkLHp7zb3kk2uH3gBTrwSm
01zVuRVxfp8ElGAN0iMwWrzjB2ucdl14SNiXXhKjefdQbATYaKat6nWcHhByhW++amL8a0PifuzW
Ls+OhEg0C37qJ/hqrV9vP+94DwjW0u0Xjm/s26Mel+A1tScprnqVs04kDWVEfrIY2nNAgHauCgCW
G5okCLf893oZFJ16/sRyMtME+VcyxePpFtmhYIcQBF13HQdsESmayP3zLc5dbQhUcG+VahZsFKMG
zWZmFOoHEFDG7UgTx3b/YKotHukwCEAOMk56smeIlWXn9aqbNpb5GFuTdOw7cIxtm0GD1CEH1gOG
grXxANDm7ZucNLue0UAoxKb52Md6sh/5eBdlnNoZHd2ruOUZHbfG4pyAEiWDP7Pgza8DKtPyUf2M
gGphSMKNqHohV4bYRsPL4+CvT24wi/L8S2oC3jRSdHZns5cr15/P9icA//DiYJ1oR88sYOWNxlYr
qU5ydqUieqcLZqT/xTGDTxRHlTa+591qySVHn11VRtzLrmu1H2HHpLuyI4bIyTz+xrS1ucpfmElg
BclA64SUzwrkdOBCSP99Ra8HujbiGtoPiGW8rT8+GMbMuOTAlJbDUi01gfMVA9fZl3HM7vMabdNN
kpKzPHT14M6KuZrGxxzL01AP6jFd/mGL4Umqbg4NClizEwCYyel2T45Ke+AB1t1+wmX4PDbzQbza
LrHN6c+xWk6qlDd6Watayl8G1epPTuMNMlvGlDelJU9sNZ56nudVSGKGI+ZPi/6E6XU/XDB62DJb
eaqZCAyqEuBghbjbV6MguEEnYVvY65wjCaF2NMXO7B+p6XhfVTjBN1yZ6SLT5XRrtcebpHRgj8ax
FCkJ5iPDApEJEjJYryzNLB7k4zUZFpSsof3wbMIunfsIhJZrWlI+bv1JIA8dpVgvU7RZtZc4kNQc
NZPUJku07+qzqaegEJglRJCP8Ndv/8nyhLQfrHrHp7qm/ojhfaCg7tVgVM5EjUAbIOSIyBDnFMPC
d1g7KsRQ149BSC0Q2nFcHnZ+3bed2ECZSzJB4aeEcWe5WnGvLtnMgEn7ciYuLOf22A2n5Vz4f6Uq
lpPOyRcq/6dBVSP4dN/X8aBeqMIkfzc0cxPvuBp88kMbJed/0OrjyISqijILPaIaKYChwRPUQOTJ
DUKjf56LK52Kh9zB99mlBMnBoRYXSHp1aRBqDvm++wBFKlpyA+htsP4X/Y6A08GWKbHnP7ZpluEN
fCl12XCdIUPL/PkCrHfRbarG7SWO7AmIkRs/xrGhl1s2v2dR9eJBzKg6p37Q8L2qs3ypDMJz1RWq
ntoIs5Gab2xvrYSLxG3WAut8d5jSlyTazIefzInZr8d8shCi/spmsUwCo9DGAnf1nbWaCJaO26Ut
rOTcYYK30EfBVQROnGPr1Sjfx5sibl2we08javuYxrO0mpqSswbQqZqhkPesEV2qvkyWyOfpmdai
OltnTFMVuiHSoqu4mTP4HTc+EPW1i19ZtUtX05/CnTyBxTHnz6C5CZ1ED8NbLmZQtXGePO8nsWi/
67cI3Q91pqZrmW63WP97FLdYYD9oxX9xYh2jO5/UNfxcenXZyMhnmL/soH16AxhfiBLwgflhiU3W
OGmdXiaX4MD2BQ1noGVHKJCX+pj/gHaG84vpbGvQxwm9p9qCH6CyoYAeMZxDhQLp6NzTH7a0qCZn
Ri5sm5jZfrNLffxkPwXPvd5288pNv1XWgOAonD0Tpo5K7BwZg4rsBJzkIfwK6x2/3W4vRb5pczF5
r5WMYpOrM356Pzsw8U/ulyCQwK+5e/S9e8LGVkGqTuptjyjaZruSINTfl7kFwGZFeoZrTG+BqQN8
ayyg1prROHpsT51IMku89dN+tVDUceDUtFcRBRISmolYoClz7WDVNzR2E3rBYewoQplmPGhCEVFl
c3GyJltqsr2F8IoXeEq4ZuWzzneSb+IndP5Tuf5s0d/uz3n1uMonfiKKFZEc9N/QKWC1fJr/JNrv
w1KXrV7C8KMlj5AW009UmJHHCR57IjWBK6LKbQAtNT1r2miT9p1boKCzqh7J3ZWbyc2TLMvAsIs3
1jFIgq/jumgxmYMbbfy0tta/548M6g/xN/7NbW/JPJJnCQiko/ievFmlcPfEYYGuIKHfq+CbqjQ1
i88ZaoPi0wd5cgWMfPyZ+zpeem3U0gSushx0QKseI7GB73nbcpvVFY0djSbNeHFbZqMy9dqziB2v
my20+skn277E1S2QUg5W3GZ6lof/6jjXgWNh9FeUhWSO7wnXi6T3C4KmufTkxTUTOLqcPnT5lDZg
G6fxGReWIG4XEM7NBIjN4Rxbhcaz8y5fjqhGnF/9cF/6WsA5B0Cl5WT+9zMDGkOLCqYMIGI6uuw7
QpMS8bHb6UASOmS/6mjC0ihW7kXp8787eEVngQCpfKKVGbCpHs8ljbJ76shzJY96zK2qZ3QkIiui
+cb57e5+gsYeOH6TNfljeMgkDj5teGx3/L59FLIWM12vqB/tKuiaVuyLZS7DTpLHMOmJRbIlr6NI
QqaEmVJRTpaEoMeGGqH5asnWijOBa3Ub2TjbbBUu9ejyEFuU5+rCwdZeMEXUWIwekUbPQhVBf7f5
c0NWh2kXdICJbnh4TvS82KLHsTCGHe+Cklt/eHwhWKY4piA+k/biUuiRyimjnARrR6bBiPFQ253Y
aRc+sy5JCrTvlxpxrOKcNg32RBkyT9JKdbBjs02feLQ+gyEZnRrMmVQgtFRaQINM+9lP/k+9PMPu
ySAP8aWkT8atZDJT19tP00nQ2IzF8W2QVjYICHpHsxg+3lLw1vw0ZH6JINd7MoLFuJKWezh8Nq5n
TE/rHg/c5ChsZfE+ng7/grU9s9G+WWEyNUzgFLzhi2q5HpenvAnJRoLe1rH70qH+ncHCKEJXF8bA
yUMIxyHn2Br1jLos7PxMeJPvk7/ZPeSq3vbHkCJYiNMLGGXkmD3puuzhBY84+GQg3M8ffUCCnn7y
/cZoESwMgtahxSndjahaA9U6U57gaQS+f61qz+ZLLWqYDpidjy2TklTaNhRoRAOy/MjduiGoFc1f
GgYkbN8Eg2yHS9FQw/cf/N6/TLsrI91ntTvOD1NzGNP8qr61yYyeXPjaZTXUigkjyDsKpqBOweF2
YbM18irmz0JV/nVlbvOC0VHZK2ywhcuoYoAN1dqvL8TTntQZ3BuE3Ry17awoD2yHNHVzcXuaCwIL
rJlyLShSYBp44pV2ONdQDTdHQMSoGGHOxr27qe3OxcG/o18jcBGRxbKAgrn52Ys2Cayu/XxNVUx5
xxs9dFbkPsbYFTfTjU/B3Ah7dm4eScjff0SlRPg0rxkdY5kDJVgc6FhB4RhKgA5Tz3Ff2LHZ2A59
a480kIm+k0A0szGRaqdtqSwl+HKH9Kj8j7qfPHEux9Qxyur1/O3EEwmC83aZN7+Rh7UMs11piXnm
iwn/nLsW3Kx4pgr2IrAnG1HhOKHd77qnokAjKuOlCNZd6A6iOGuKgx8BOq0KBhnKHWNQ7fX4bXHZ
dhEqwQIHgg6xUu+2L7/GbAnMmKwIVDZJAoRIjeieDeYPIUGnAqAt5qN3CfvEPCb6DyFjccNePsex
yy0N6Di3wRKZGqEuk0YPm0zdzaEw9Mk1SqQkF/MCXS+i6tXndpWpXlJec32atGmvVkT3wtf36e38
KGfeMukwl/Sf1Xh1inZpHWFxfgUkVNd7zLPHomh/3MEFsT9wXcqLDzHkzqNsYfcJ0QtkhR6qwo3I
HZSy0u+D6cK7TNkKNlnWsTkdlOjOxNIlBbT/+3Ra5WtifMPMiDfpnMql6YQoGSe3T4noe5t/iNtU
NA/axLjyhXHv+YqkXRl5Q4P1XkJyAUuFtMo8eKHTOYub/nNbgVw0fn8GWHZv2xHgwloq5FrPdg7z
UL17t5XogpMfoZ7D/sABkltAw7CupsH4JmjRBPj0VGwikFwHY0GeJgUOzVqYl+VYvFhkXJH8Mcar
JlIJYLVyLlWPVjvgasslTK+1uVmnzMbVRz0FDQuwl706/CR2GSjKf2/mWSu2InDKvDXY0mXH5ztu
xVQfCIYXfYCeD3e257oLoV8YNrpi34ItBP47ggUHAZkFMSh1sXGIXT9YZA0c1BloFpGzPzT3L/YH
pIGw6zSus5K4/boUG28NdQZxTAZL1PWOgaeGpd9tkWYtWa7VyMnWQpz1S/D4PzXkpf4Rye2ZZSdY
bfYs81tG8MO4CV2JwyiYX51NM54VumnaDJiyGGatQhw/MIZGoYcYp7DMojoiGXpRfS7qr7nsfXh5
KsuNxiOrBqG7O+/1Rt4bNYX/KVZZGk4jqqxqyRZacMImoL3ZigFJDSICn4S1r0FzmkIl8APhjzN/
eRUcxEokSDjm1MrzBT/wZDNNWPma0Elcer/8cdzAd80+S9albNb6U+UExn/TPC5QE5bacRZew1wC
aJSmHFWMaHy0b8WEqqYkEfioBHmA6nL0zHcV9YSyH0uKQmJlQtNh3M2O7p1c6UW+CYNcgBTwa+DL
JV2mlpvSAzXHZeIKSevgfxY0/bYsRwiBP+uaZHpeWv8/GtmgYe5avTMugxEgs/Zsfxlr7y/pI4b+
QCxz3h+WhXGAWhiJsJc0nW4L0vmvP5MNUzbkfksp5n8Gw9H5ZhiPOLvRCU81jEBPBblnb/v41CCF
EUZb/DW3WyX+XjrbpAJkMQRtLEIxDW/GX8YOHorHfOfMa5BzjQyGoLbjjCp8Y9PLVULTBiPYSKbY
mu3OJkrbzlMY4Ys4tEn3SxFzEugynlnmfgInspPYHVgdeuXLaA2AczCRaxZ/XsXfDWFgbD6ECMFk
cdH/CUCF6WVNNwMgu14Fwa10cgoXn5BBrcpqqs178SV3GetWEhqB3VQCVaEOcMmsnNPC71fUHhMF
FVxDJbuHwH9YZBy3EJr7HLQQeiYrOM0gC1kIb6AUS8qKMHo8MhV1rmRkaFZxUwQLZdo9vP41bVAp
Fei5i3wf1/pmW5tfQrtggEykZ54OBrMf7S+8w0BqzROTGRdVBM9yb56Yzhe9KuQgGY7eiQ8ekVU9
C0BuY5vVSgSa6++sWgnsNi7iHUJgwDaXTVbueOZOPeFEi0p7AcIvOs51175Qs6HEghpZJW4Hmwo9
S9pavFqFa5dI5//DInlTnplXtTkU2QblNBCwL0aZBPzLNZTgNQGUji7dgPGRNE7/B6udq05tSbsc
Zp98rxnr4OLlKD/8z2XdTeMHyA25hYMLZ7m4pJABBucbGsKUlNo9VVZqljolp0V3iZHv8lh3YsEG
bJXTuaPFSykpKeh/Ed9hGMlXJi5T3aS3Q61ADh8UkuCP3eMvpBpBGvoW2q1o/OaZaglyXXzii2Nr
YJhJF3UHDbGMA7RcHBiN/G3DNqZ1p4Nr6vs+Pushc03zJsnb5OM/1ZwMKXsf9PyoCwnFzdzSLybe
NwLNAdUXAW6yALTElS05gyhl4Guh+DE+O2qlDzJJPAyii0L/SDUIAM6W8M+38JSRlGwkWHVtjjgp
98XsO3CV/VSUlzQVESNak9gc2gx76ovamzCAuq2TmvOGpfGtVZhPaCXr9FfWZ0oiP5kz/E9BO0Rq
3TitHcB+Pwo2D8Jyxs178cae2UXUi+vj3OErm7tGZ5BkxuCxas+PlCHZp7liLLVPLxNjVGXBIzl8
4HirJlMFQuO6TWHuYQQYFRUxVGcVlsrbhHP5tufdC4Vx4152u+UvF/AWXMf9XiZ4Hy4sI5ymdQr4
c535LkGJ+MqRoIpxq+GJfGcTktoqSqrkiByV0O2+xWbAUHY0KlmCi6dxFCHci2emXb8TCw8VfNID
oHzfEHtz5K2zEoFowPUKciGlatwCGEOhqmEZV3YUInXhvBj2jCWCuL6nevghTt0J02BRHoe2htyN
BwgLfdK7awrAI54EqPLBDRpa9gOeCYHdq0BrepZZa9D48XGqBdNruvZdb6rMGBfaJeXwM3f0eHqr
svmdM+gkMJq4bXp5CmL9cm/7CAGCwrEXqnWKy2E01JWCmxHhWp8J9e1i8XZ7JfWMTurPbDQiN3Rl
PezHW+2Q66aSf8wfi2K/XRdDThUFyUJqdYa9RjnQQ0Yc+cJnUA4WGrRBa+s2a2TWG6uKi9e5mr9z
bphfDpdN9RuuzyIXUsK5Ix4s65yboSIvvK8bXQ3/i/JVqd4iIpfJq/a4g2UgvPbNDj0Ll/aJSiog
Lp7sfT2PxeCd0cu4tGflmzLTbI7lyPA0ETN2rYjmdvb8XDvZtyAHcBVFEIU9Mvs0gfKORJBQTSSK
tiot9eVEFI+6ei/C0gAPqd/prDjIANUW62k0bXf4mC+NVVjESbOYoly3o7XrP4Cf43LtlPC0MZkN
yf2Og0c6yEftIF6GrZFXeyN6OjDX0NX8RH7Tf7HDXWuZz9ZNPhqhKGI9HqChOB80Us9HPKGhoQ3N
GF7D1TQPOqqqhtfd3ATf/VcEMQufgasaxrGRvVJYQsieRYy7EKqzADS/mdzjoyKTQA29nRwn8pxS
NO18c+dRQ28Q/hD5ju71ERS4eSINMXZKGO75+KDY41P/o40eeVAir4gY6Krh6JUSNN/g2CdHXrQL
10iINHGIuQzIF//TIlseSuCFwchTUP+c/wq9n2D6FXDXFxln4Rr7uqVdNiJ5nswPa0n8Z/cW3cdz
EGkO/h6pdevWrGC3AuLy1w/v3CEnJAX16ndRyNDuqZYuEeG5+5MR3xupx6RHDIiC36lYE+vGag5C
LCpXiUJLEfA/3kAz/smT+FlzOZcsLFVSowEkAWVAYDNo/3JQZChXy9N9FSIUl/DnvF7QMJVhagYi
WNqkg+x7LT7KF6L4M5XijgQNkem891Ir21fltlKNp5asLIp7UL6xM+YwnyuJ5k7a2VB64EAwTCnb
73hTQQuxlBFBqtXaERJ1wzJ4hHsmRkPlCB1By9BUmfTcNROfUpfCcHr0Ptm/fHklAIsXp5aU2fD4
lPe9gSlCAsW/rEe+NGkj50zfX7yNB44Q9HP0Pcj8bxi3K+TwNEDDV2B1Mn2n7nvwgzSXtwQWJbh3
whLhJitHj3xx7xVnWHJvamvZUx3LxKaDjxubb4vkgqqJPEYGPXDv25+4Ep5oBwdDISX02Gcsbj8I
VRqnQm8Ho4Q/gw5x7Wf+/TZ6Y9hAP9sJfmMH6Yfl1I7zc0m3otHhSGDmh0nMsmWQcPDP/oR9Jra2
eEdys4G1//GLEZ9Phnk7Cvl2mBxDZ7+YiqQiBmYOB2PRbzDMpkWWpozpLRT3B9bvM15e5ps+XBgX
QzY+7dwJ2bBJ3xI8WMFmdvSHP89XsZxjPiyf+2jv/hc5Q3guDkbMifV8PmzRfRm5uYfMzZWR0Usz
Lw6Kg3zyb7OipXizsPIT6wG83kpuUX1XH7tynoxiPiJXLb0YdDKYmKH5AdshL7oJA2Ra9FEgoWdY
dxIJHucmHid5bTDGmf+A36hasgyXBzKmxItohtppHN20cIcoxTyVJqP924sMLCiU3PJ5ZbKN5M3H
QBmzEG7x3VMh1O5jzChzkGR3g+ipGO6eGw6NLPz87ayK685p+kqKzP6obxaCGojIkP0wZv8jW3hh
2u1BFkYWoijPvcLHIzuLbzKGBL5qPni9YPLj00PV5hjjHzw1yD6A9tzR3vZlIMivOR2/oGEodaVu
dt8tnpG+zMFSOCnmo90D15PKwzZrE50bUMcJb36jk6uqv5VkG9ZZrcUr43gR6w/09Na+1cL3VSWX
HT2N7JLbydKVMkoSF9WtLG/BjSxBqdFn8g8kxMFIylft4wJHbtA5Dj0vcjSr/dgqFK3V5+pEvx/z
I537tXwVDmLaxOIqO1H0RCC1I80Fn/GGF8QiIEo0aw0OZT6XYo3BXjQIIz4RnuUgUC7gbv7BnXO4
MxEDjWp7vnrpFQ+5VDgqr+LlZkFgZaqvKyhkWb5e1sQ+JZHjDjp4G0/Ebc7n/MkAbTRa2NgMaQVR
Nh6XQdd1/+yMALCE+78lkec1YYX6YOjDxTLvHGfVyPtvLQy2wT92Nt26ygxM6oUwCbVekbI9BzJl
IhtRFYBRrX3pbTt1AptirLmlxtI5/vs2XHPnS8wWetV2nrtPddflLysfYthwDJZTrgWKD+VsE4us
of/qZlHqueb0xb9VQmFMxNQDBXGvaWCn0hwNTXLPbvdcnbCdUpn/lPwU5pAcYwmazjVmJF0cje1v
1KrgdYlgQ7LkCAJe940ggqfzyu0lKOZ2WFDuWUMXCRVZ75rLyEm4c2HPUHAEZ294lHyfH5dfwVr8
RxB+yxkq2k6BED9uekJ4lVmubicgMQF5RVhBpeqf7IZHu4Av1DIYwb2xvrX8FXHqTcL9awj5At4m
RXUTTrKqwxF9EWEOqXXhqzatihR3HecmQpY+SL157p1fnTfrix3GG7XAzZiwqJ/2OL36TQ+6hK+k
/HIRIQBrrqO7RDz/ZEnvp11Pd7hWj/Wm9TFEsxYhHx6h03eP3GXfqWmlTB+YC1sDeLyXJ54I7hmX
5i8N7EJmmOoBjgDGivx60kUTEseAh5glCGzLkLxNUf1vNif2xMcaTReL8ksVD1QzS3lm5sKuUlf2
1Ktkw4ASbyErOVfdzbtCTGpvYfh7M8A43O7vTgpwpXjuY9V4A6t5GqsQ6GVtDFmHpp3YOZwSpYzn
5I7pJnjn4D9paCO/K+wlu8Lg2KZm85BHR73S5Exr9UytelY2UPoRDVDLl4HTD7+fw44glHrmPH+1
Ec4JXGAbHu2nc58VkaQ3tpob5DOIhn82YaeJxDNc5rktus5RhNms8PvtqqnZQ4dfV3Hp8jwGezWU
DGo2262jeaQledk/cNxRTcS/ZP+5HRolGF7bCfQdEL8nOfyWmrsVeRS7htJwRcLHx+O4Vv1Fn1dI
rBrU/VHuyxU8TSJuB24AyTTSeToWp3uIDUTx52aYtn2ZJAYBY9rayRsMBZUVAbbE0lY54WuroRE6
TExn0cqUboOquehAA4sH+QyzbZ3oLCtP9QRSqU1bWfp8JGBfzMMLOBMS5uyHOc/cwniQB9tg+G2x
APDXH4Xg6bLg1lybT7getGh4sH9wTuuBmJcYTMbpA8vTZiXulNmBWtF1VH/BSSZ4wyfTfMWDE59X
rNy+uxeLbm+g2fGdL6pAPXXUHpL92gNnqKnL/znJ7kz8/YnKx5xBcsOJQ22Vx7dxIPbW/yDQ6cEp
rwFSGiHS1GKE2swlledfPSeg/BVCU124kQ4kmTT8oyFBNLE2BskJq8mh4f3jaLJLH4v7qOxRSsT9
JzgUmJvipgZUnyjPiB9CIRuzjr/UFbm2yq8s/0oY/zcH91TyPfFMm4AaJTM1SYVWtvliWrbSTea7
RixrCz3lxXKti8Gyn5FVAqGbHbJmJ5fvnE5uCfGV1S4zlYkZz16JZCQa9QcITgzk9+V0V53kv2Zl
Za8RwR+OLc0+mcwgiDWTnHOI5GOD2Juvm6baCa34GcpoupfNAGLOkH7tI5MUyqne78knmeLq3tCo
JMlbsJu0X+DS6i+4DaLxrd2UEq9hJ6igrchAauLbCR5JCHBtXZ+NYT+P/etkEXKDI8HNSGKMeLmc
7cZsJ1DlngSvQlY2aY0RlKCuJ9QNIr9qf9wPItr1rvW3dE0UaQWo07bQC5BnnKbAvpXT3yW/b4gZ
AKZRIaAJkoPBmj9rQbmK2EomUmAKru46cnGaEsPmIMkh/irNa1it4iWw9qc9CneJHMWxIOQqJwXR
va07IsGmFQO26aEN2zJVVPfe8RKGRbCfUyJPR0BBn0yNHnVjb/XAPqTj8mkB/9owU4xbZXXfxW4t
jtRClCw5hlQhQCCRy47v9Yy0aUwEACyTDJ5mNVNJAA50Kh9KwIkq7nQVCu8Se9eb+nm/RfGjjEdX
TgGR0Yyofm14x5xqUiHdduCPhQDSbJ0lRAtK5An/5kYMOGF10Hhs6okZAnPEvdxBnfgrF6s5I+qY
peeNFwW8EIgS0Tm0TcMk1lwZyaIQSi3BiHBy1jZ16Q6zlv85bGZBdGlKwxplSV/RpmZosUSmKBMO
bWulR9/xDkJlTBZG2zTm13tn6RFpGCwlv5jaK5heOKGhhaCEW30MHFkxDawf+MZnqWhAJrqx1XdF
TBJBsu2ffezMTxJF1/a5UkcG/hyNj76K6D75/IFABvMwUxcZeL99tB1IRoywvee1f//eQBeqYheX
SOomKZJHNINFThnzouGPgXBCkma+t0bCXlo3fQ6rkeHRFZPUEqRc0138zPvLN455WWH+KKNcL2iW
1a8voAmNqBmA+bOZKEt6alLV4+mTnFfyBqvVax+QfY2kzOad1smd1Ey9DYTdm5+gTaaY9nrqcOTe
CvM3wYBTwLfTCNfAQweuCBAQDbPmQgoiIRGjxwd8Dt+kIWmVUmQXLHyz0NGyk0+2PEspetNDTc0n
Lz67JxI2zJJCWzWoWPEF8rmAVI8yqSor1lqoNAhSqz0Ud9z/zJFQGaDu1BiI4tiHWEfZjaNq8A/y
Ru1Tb3opzvbamlaRj1y95eLLgZgVzLZF20AXBYhtk+rTRuyHFxTKWaXKE7DyNebwMrbQJRBsURFv
J2AoLc2SXWzYLsYQG80xHAPgam/4G3arwZw+gU8URY90fCuvl+mWTk/RV7XC73/rPdFkE7gbHiqF
OsxG/XwXSd1FWhHyNQIbG+KMY5g0yqDn2S2OMA+mWRSWSMq7Aoj3YMBwnH9tKU7xT8k8znnKN6QX
C5/hyczxUFkBjaZ9f90GD8acGKI5HH0gfsYkok1CViVacDONH26OzQRPRpcReA5SSfZMRGUiZLdF
oWfh7/gH5R5ENJwNZIJ7wvBvoi+fo1WoqWNTAcI8PAg9D5t7HEMI8CENCcpoTfTmAvMtWK+wt5qf
7KWmofChyVAW0OIqdKPNmkQTx8n63GiCb+JrmfWvwylfjr/jFr71GBZTnpUdmciOi/y99R9Bd00/
sTjsqV1dF9Nr7cor+Os1KMw7GIwT7K/huLECxkw/JUiaQL4MDMeiOYclyu2cYFULdFnDXJ15mrJX
RPxcjeBt9gDiLxhgyaYNotjCxNUA5BGFuznL33IGpjcyddYWA2vHSkr+SSC7m7dVb62YZv12W2vp
VAV5jBtH8fBgSZ4/xsWZoF0/fK1s3Whgb5HRlyqHXmBpCTQkN2pmmNSsaXZ/qr/ZuKvq/XxWaRgV
x2OTpQfw6j2/DAkOnKWh5oN1H6y98Y9BLX6ZH38QJp09sKIQ36Lb8ZJZbyqSDMW6SMqRg+q2i5a4
7RE1UoeTqTyyw9F7FEPEmGl1DYavuFK7oOKnZ+UPfvCUeA4QPdSQmtjVBU/QZ2Q5KofffJmlZ+Y2
A+0xRfXmsRACtfau/qtDl+TKnFCUCrKav9/iU8VoQutqnN9mKAwdvjlLq9iO4PC9fBzRY+wTrEWZ
wMU8G0uBw4kU7o2AJ13rsFXF0gToc+V8iWFty2mWfBLb7qGFdU8sxa0KrUAMzXP5H64aaHVT3BnO
Ni2nLmJtSERit/iq8WDeUxtuLMrz/ZpcMvBWNXCOptZwGpaf47KY1CVZFjlYTM0mKeJWvxRS1T3A
1heC1Jnk3lb5qUzMtcwWoZg3eaKp7b2D/jvf9jWKNwiICIFvlvl30x8MUkzssW7lOkDAo1jejxGE
2uIFZ6XFH+lwikou2rkhCcbdMH2cwNjZgHXnV35rJ98rQAgfrPLI3umgG8NIqgNXW8SUrhsV1oF/
4B2Tf7giWiAlkCYR/r/uNOT4nx2aA1m1roRyH8OvQz1Ky+H2Yx9+xA3T952KssPm0EcSnApjbA22
7m8SrP7eMxAnGlJ02l5k79u7UA7x+0LjGodHDe7xY3pUcWEB41Is1yV/6QW0gQgwe9ikEFQvLj3a
kWPthuNjSqWQ1+zmKXlqUiEDa7Of0IeXODBOb7Zspe+aC6/UGvcTv/9CMD/u9vyfduZqqiY5c9x/
bq2HG080RNfnbtKIHUPVaMyo+AeykbY8hyGBupZH2o9lWSOmglYK+KIrZqXN3FQlpKCFYO1TedE3
d3L7vProecsZ97NHv/5XGf+kXcjze+sfOmQOIbu43INLa/lzoG1izdnMJ3rHoOrN70ZiadJXGDu2
yrqDEK9r3JNB+TtAMnYZ/FjIfNg/k9xzZdLAiSf9Q5CrXTaFTdo+0N3rDmxFuWGIWJWd5kd+LCiv
/8IJ9thzgEX5o2C3ZJGQTN4kMQRCg0dRJKKW+O/WyR2kDXGYegL5Ge4KHo0RqqmeXRuIUl9Dng92
/9wd22FPP4tWLm/DYoCPOE2s3D+YqnW9GPgoTu57Tu5q/Tf92RVoGOrrkCFzwLYhGSdh2cUS/hZy
qG1IF8hsRAGICrALvUgp5xEsG75DUeT4F/GHtfiIAC47egJeB+grznQQNsXUdyIEBStE0CNYviWG
VjEZJfhvYXR12UAJFiokgXFpFZTdj9FNSSUuu/QkHWI513lq+ctc1bRJaV3kt03MNUC4A6HHn/D5
EfUOm9OmEdfWK7ua1nvoIF3duZdq5s/BKrMG5ewcvZol2+Wr+rkOTAriLZXyhWgC3sAIK3ahwMfP
ewtbDbF4fsVa3ilu1bczwOui7UzOXpFTb9oldNCgEveih/DB9X4NghkcZ9CsDfDLD9OJnSTCzLZf
amgVt8IVm0v8r2Ze3pRsniRP1J9xfKRZJ4r7LNIjzfAtfuyoANTLYtcN2jCqw4ANryGD5ARmAX7j
sP0RIU1k7xIrk4TJWkYWcnaaSCTifkNMU0FUvaiF5bLKP7V9MfAu74tH29eZIcCj7YMJ5HkqOOPc
X/ZFI8yK6Ll2C2yWVTUUpwIrneOxOraoZX/BPVNwc8rA1YqEjihKL6gj1GxFGUkw1QTTbkZyLI9v
ikJSGkinlQ+GygQBb4FI9iBaof80b3W0T1z/gQqjuz+70F5mrZErINk49UsSMGzfc0nxFm2PQcdC
f02te/QPRIbL6OdXdzKYYX7LxDHmeZknwOa6hSI/gX0FQ/KOTThKHuEXFMGo8cKdf73WepDIz7Ph
un0yAssy7TjPbYnuHnCHLxpPC5cjkXF9laahPihjQGB+BxgiwaFjexP+eMBCnQbdQzZb3spN5HLb
YoJGO0XOAG/y40+SqueQg0F9WFo1HtiojIy/M5VKD5dgmYIsh8WKqg0TR93+EYW423NiJ+aoORln
MblCVqVnbC9eaIv04vp/uX2HO1isE5QKZ3mxvO0DOTisIxfbD+g8xau0i7SobSMpa9EiZcBIW/WC
KEXAl8iQYcSRCynkp8vTAHsmBKWg+8uVZspjW9ChJqad0dPTFe/Yxz6HBLSMNi3dotSFX3t1yH6l
t0DjROXSIAfLHMbOjFCFe7rN4NhpXAhaA6anRVLvAfGoOBjhPfvh1FdmYf2Id+Enqspl7i2nw+0T
xFKXfV/efGtgp6JNRHs8YX4Rg5sAt1cUwLbn08r+vk4Cl9yvldgkQ/TMyLUMrxC4cJV/lDmlMVes
7HBmi0MKnZw5zHx/gYkJhgeLpvBglfAIYfmzL4sLMRey6WCQc1BCdjioLVVFNCk7C43ruiOrIYgn
3+kUbolgmJfT/I6xFvRXtONMU78h5naTAJEH+KsYpp4D0OJttUGJLFrysrJ6KQeplaWOOPmxPcYA
8LKLbuGpT0rKmqtwpKtFg7SjnyLuVaJA0aSfK06T8yaJ0ggOiud236BFxyQLBdMUji54WFPRxi/5
yS2MmsRBpHIJJlUH+MT3Jk8/J4tFYGhCrV40t4zweVFUkKK7R9EQptqKNiIvS06nMCI+DQrPHbqE
Vkfs9kT0lKPkqew6rswIPhjNJCAsSLJTsWGwmTazP2gKgvmITpFm+9h4W7iFFyNTI4sriJ5etXHS
3EZI+x0OdZ3Y9lRvor8ABx1eLWOEdQFO2aFYsqCXkqPB4n3oKJ/Vtvifa+MTs1aWCIX3hkzxPnur
uiSV0ZBmG1DezLSkX8/x15HNPqoF8+MjDr1nTbK2TBkmx2xkeAPwoM4k9c8c6PJ3jDqbqE0BG6rg
Wp5Asy6gzGlyEIcgj6xKn6F0xs2RezIJQTVa8c/KENXDr0iuMdTzgRB+Ks6tADQG1e6IaExn1TS5
vEvlK6XLQw/IFJNfO8k3ZgHf/Zy6qFa52P8lOvzWTIkE5pv6J9GHrU/9GMXKfEqzjSVCv3fItsyy
gAXY9YlBtz6CS2GUNuJ/cyUYU/7TpRV2zZtU+Scus9oLu/RlNVuqy+1NPqzJK5r1baSN+QgO/fpO
O2pb1DenZ/RXc8kEf2aRdNGeN3Fw4ygHyb2cFPTqgppWum36qzbCSbd3onParWfINnDt78JKitkx
JfsmWVCOVDwbCcd5QkyFp8jdCjFpaydEcpIDCgx9jIJbGnF3rPchnExZR/6ZeX3WvoILX/gFgxng
tfwCVsX/U+EiKL8XnwCMKIgLQ92L7OkxF9LTEAIuayPmbqZ4/EQ3xYuEbF7EyPXintfN4aXeFUUk
O+ArduK24rvIqowsP3TmYqXGpzPecd2fkNnYhPAL2MRX1oUVwa5ZqEl65b7bHQJYOM0rt2jc+dsf
JDT1P72Z1rnjPVl6ppif69ooj8WrcgZnB+WvSZhKshuIxY+/CqNy23/uKFDoA4xhLo9PuPyAEvRd
NvwfLQC73kSZHUkFrpOnbnkzGMLSdPTTqv7qulih/VlMV7ArrqTEbwbaOp/57JANwBCEJbBEUJSw
eYzdZn4u5IpAjjw71Hkqqu5jgEAYTpEgcf0ZqGOR2ogZgKl96/nwZRBV131eBipOztkUOkd5SMZt
9z2KOtnC5E6MR3Hs/rWfI6WM7USwtAqvk43T+UlglAq5IIvYKAydP52D/g2XD995PeD2WfcI1Yzx
q5aK+wqBD0TdOtX3axLvZJ7rkwkxsOJjfrmbpbed0viVrCyDP07xsufBq0fF5YfNoHI6ins8dGAM
JLRTx3ExoAD/+xcFVRbMRXc1h1zzGh84fRfm/ppUdE02zyYL+97FaaFgYZNAXGdFLunEqX/slgRt
0Pzh2yhZFHWYkZxqeAGbxAqVufSsY92LE0JxVpEWQhL9ZEkD1rXuisf0WRVyuVKYFZHAW9nx6OKH
2OeJ+qg34QjiugMvBpanCMbbnk+7gVpyf3GbXbCTsOf7X+O19CCTvh/rthBFPiOZh41ENtXnCDzT
x0LgzPYKSx+7XKP9QV0ahQd1kQNFEwZ+PqnWkp4K4GqFaQ1P5A4GMlu9sAfh4ikMqysTfxxQNNik
laxBqCfyFw1bdBVaUOzPWYGU2AMGoTFIm7KYB/O9LpG3IBwk4larG+2h4yonFR56AtcitcQ9Khxu
W3FDb0rrrTD91jLOGxx6LbPzwd9VQrEqNEmPOATSpaBNHJV/6o7V2E18xVpAEQ96XdTfQu1MhVHU
WUJXiL+BRIgPiTiNc3n5FS2T1BpqiH/DbLI5ZM1ytklf3aedlMsWEJufOkd926uR48wOPo0B1+hA
9BxZXLcU4etlwytATDsLEUshvqyxwcB1zGFC7+kcEJ+WfCAHSJI2Jdtlqk75rjSUo5n25OLEJvTG
rnT7KkbDRK+TqsWUJo/3oVBRu5PFK+dCnShVnvx+W7b99V1CyZgyoVUgWKw+cR5Ay0Ua6IeXGHRQ
6CRrU0tdzH4qREBf359McC9dj1KaOGayGhpPCm54cJREai0CMh8pHTTHH0DDVUqaRpAw7SHtA7x3
9+nh5+BY7aAzrN/Dc5+kLT7BcF+MxnpQ1Vzjtex3pRH12U3mmCBYqy2onXUuIhYorTRa2EDlqyya
PG6edgN5e7KQg4VqSoT0ivAf26Mnk3YHVhTbgPPPGCohdsWRYURJXX5m018WnwGSN/as90D5AzIv
kgNx0+CAdVxZ7QP0dI+Yz8M0Ed2jRRHgeFxSgtbz40U184Xk+bzfYZZVxSryEu2/Ut+MIaOD3HBv
2VspndaIvMDEtIV0V6r8HNyraDqZehYxq+qAbcM5elDf5oAlB7Y8K0rGBtqcnuDU1/jTfB2o1yg4
6Cr8Urpyo3F0xRBslLWGqyp5gftA/INwkY2OGQ2gDc1bS2hA6x+zKNXJdiOFeBc0uzYa+HxO8Y+1
r3nnw/hVoTOTr78xz0UM2lVBTuaVgpHMPzNNQrmsZyKMI04XL86lXxFjdcRoUXH5COs9B4sFMYTZ
kHX78Yrk+tE4lofcpw2Sss1RUdTWu/Tw8gW7ze89uJVT3FCkx59OxzxuBJ2yEeZr2cSSewb0ub/Z
roRNcEfgC/Et1GsAECZvrQDxPS2vd8nEQIlDsJnUzvPyJzp5sORBDtgkIjCHkrLytc8EzuJPOPNn
Gn9szqaPa0rdwsVAzsDaTETpunS3/xkjeT6tvniWxGMyUztIzwZqQYFogdkvw1Rc+39U/4GXoKhH
Rok8WICvaROdrCHCNCAgzCaDAP6QrjqpVZOrIUrBMZUZeE1zjJ3YTPGbKwYXIakawsvGoCPIWlB6
Zau6iwM6wKBltpzKCCoXosgqLPiHqHiWwO5JF++iBujR7fi9MzA/UTvd2pRhQbCunQ2LJpFdo4CI
1NMOi+szbQxVBho0iTHu5lEZ/jPoBRn07+wfgAdME3ki4gp0cKURBe/YOq1z7ZKv1ehSJIcrlfD+
aT40SS8kQqChhqyhxEhludt8gdJAG0lODKbAMhyzmY2lX3h5Uupm4Vz6ScHLwDNZcvjuMAs2xxVC
2sqbtrl6/247diucqxr4NZQYOOppLpQjzNARE9XJYX7h1BDn8i+6J0V2lXZTwltoQU0yCM+UQJE5
w7Fq7oVP4g2ZxLNveZobQIECah5xuMSAo93c9RHnxXBwkYqLlpWmn4ZJitVRHVkMcmnjNyd3J6CV
aE+HiVZREiqGW9vKvUDPRWiV6el+7Ac1NjKhev+i+e+xGeaDCJI759LKRRWr7wC6SNItwixlGH3q
hD7d9Wrn2v+vA20Te+jQssMw5YFbOB2KLnl8CBfcHwdLQ9Eis/XYQcchPhKjco/XRkUgeHno4nKE
R2RXfTmmlzwHiRHK9I0XqsL2uBvFbFBwn4gMLdtoHcoABrcz6sZFHD7MEztVAP/Oxb/dPNuVUKRb
js61Rg/rMy2bwdqFnPdXjvEKx6mUHkH/CeLFt6WPmZD/SqLMI981m3NWT9VfkT5QCC6GL13OmaKf
69uRNL7nZBJ9JCrLN3vS8PTdCdvdncg9GznGNBJwQZrgOxWqa7AEXWR95DZOl8tok0TKjbRPgtSr
d/3GNEwE7ESslgRHPHtF7W/tkGFM7GEnOZK2Ad64F+tyuIeUBEru1qSKck0GBUa0KVoX1ojhryml
DGMv1RsSE5ljwfIO/9NpfDI/ssYt1/Bg+lTpKmtVkY1CCLD653HZF8LeJ8PjRF2u3hgi6q1598zM
PauSlSTapHoYNawl4akousY6CuLUuTBewWdbU6vmHvyhxx6iiLXmNMnZ6g6R1kuaSD/gQgawxi3W
gvzdcO1+WenIcm6mVH+Cok71qiUUJjsXJk0UOgZr5OxHwpJTL9Bm1hGIDRRdH8YRz1gyfpa4nCZU
+ygRnNAlVmBliW876+TYlmyGsEXoH/VUr5oYYZuinhxqSCYnjchnEWhrRDAujaCfB14AkAtq9w9l
5V8sQirseLIXqR333BA0gEYITv//lXgcnD92NIOQxIYHzKeUCmT1WSmX6lZ64LWK0hQHDKS89y3i
1XCVYvJkS3VCdIHOMKfWSPz6jm9KNGlCL2Dnb6t/Jit7h42alkW5LYajb7MMSpODplQhY7TC57vR
qZ0isC4jtdXtjqmCKaTCydDdk5iYkim7fsjJjRhzqGdXx1bryy1GUPa3Scmw9P0WH7AcG+27zTA+
xxpPlcFWSJ3ge5WCgPhrAovWIrq7TKMyyz02amGbE+khXkBt6+kzO1+4lE8IZaNb7TPhEFjlgLJZ
+ISVRIx0B1Rtxkp2sq9O8/NKbRnZENTNDURwSnNgB2QaBXHwRZvBiv1LEjUlIVxlYXBzyz2lskQr
oWsyy0gs3a3q+t+/Gyk4Q/oc9XCRrpbBiYkYG1LqICcd7eFCUgVeaRwPcDRbTcv4jQ3u4Z9a/uoS
BnOEsFbBVHzpvO9eaBRnmeHYo8bAa0D+1JVAt+wo/hK5aTArwFPIgKITbsC3GgN9wCTwMdChV7M+
XyvShV29oN/7qY8HIVNeizkjqX3qVtRUlEU3+ZxVwhapWlMqev6QHRlXP+gkxq37iaPy9JYJM/Rc
rAHQRedmo34w2cxPwv5Xljhlug9oiPaDF0pASTPwA0z+Tz3SToEENUCiFF+n77NlFKBBxscg7EAb
d/TjBfqYWgj7Quk27P+tbUbAsp9grs+SowYkCmKbWZ4432WuXqSlWQegAXbq5UN0jGEmlNo95SoA
dORAzqzFDV/W38hKl9V2vRZtUGd+v94cbBHVncWZzrw3iv2JoKThprG9QKOtK+ROUNlFwIr/1FbE
ZrqpU53hroc2e+XL/ob8ZroF3cc75NH1S3mhN9ADPWG2T8nTS9eMy03BAQkalS2zLkABkKP+FUOf
iUBFqsLRdt/DT7E+pUfng2vyiTgK0weemTwHCihyzDCJ7MDWC1KGBguIq6xT0fL0XgWeO0gcNWVK
OnDtKlhfhr1/L9BMxQFK+JP9ERu04SjcULvzMQucvk8VXTm4YmM5UqUek7efWwnSuVpeMNgwwwce
9lCTpw6VobsPx5jhNwnkEXENHH0DtiNgGFXy7r7biOENni6XASLsjoiHESNq4BuGEbk+HBTLVfTw
KUKK2CaA6h3SnCLfOuMppAnyXCEj50Zk6nJpnm7Rxmd43NM3Sf2CAMiTp83hO8tjXjMxk6RSgZe7
NJF7WnApLybSQsxnHNIzhxdT5csJ8RuHm4ZcvNzxXOehZmTJ6qZO4A3DNCpiUUhK987RLB/DZko0
lc6gPvxnk03MVC/AJ+xvpjFsUzQmrAvA7SzFbIrvK068E2BTAPssocp4mrmeCAT0Z3Enp5dVjTmt
Cni44UqBn4RylcBvYXEcMa/a9BBTyG65mGhu4/3oTv6daLWThTRFvVUtp3aXKIm5d4deJAOmZXXh
bMB4sIbSCcdeotDz841bdzturU/xzJCSQoa9Pe6XyXWMKUeKoax2Qkkc3Nu7Hm1EsFmoTPudyAoV
/Lw9Lx4wxL4rOi1zYs0glldluLSvli6XdxWhLI880Jph7lTYxrHWQuiqwf6ZIcu+hQkYOAwSLQpU
/0fCOO3gv7/P425cBoWX08D7Kvh74KZJ9VommVyt0gj5JXQwnG5tHGDPYpMy1xHAiD6oO2juqcji
d53zjHkAyU8+hr8dNu7RM55MsycCFqO5Uaxl4BVjmsD2JSSmC3WFFFyNbj7LyPS+CVbbVkugoGe4
y988t3ewuc380NMlBc7pMzoKAME7SBMmFG9bE3tjTVFg/hgw9Mtluux+dNTrhfQYQHxmPHwxQT19
qEuUwug+R1wkTgHlaOWmDGf6Ixp27CRVY3MVVIDJtBF5gLal6hCiu0FcP1q799W+3FyjiBKrkai/
34xcX6rlbFYerxj8mdasN+7FvV21nsbu8x1TLQyVOuUOQWnazxjV0t84CJXF+em8zF190t/Up12+
Cmp5kJvlMGUlzP2TRz4iiKRU12pRW0d8BJZ3qW14EhIxjbfFy+gckz3NxSOoFVsi0uoUqg1b/9bW
Kj3IFHbgMcDrJCW+L/20CsGnyI11blWst4sGqVsJv/S+en17TAfEbpjrcSvT33Fd+BGxtScS8S0z
Th1ANe2KMgOqTLBN0tjSB3tsnX6uau48z1MysDGVEIGf9RSRXw7hlJ7ji8XSueqvvbVypoc6gdEm
MvnP5QhdGB+CAjiLhIGkseXstEpBn6pbCURFxKETlkWsb99pqCcCowxMaGhxXDkgmSxmchFPHz4i
rk63exgBIBiEs3ugprY857ehKmbEsILMhKSWn8TvclkcJyUGtswWS2T28/URA0pKYVdJkNyoypHC
PIznpY+KkDNel9+248lzKTKPswKGRA5ePy+gt7wXvm4p7XSwrn6LKuiWtxu8/xzNPg/VBFPyqIeS
jgl9um3q7mFuQam3XsbiwAjMc4jJIjr4H0NQ15/9kkSljM7jYfVVEaa6Yngp7lTYF0vRFQ6whAl7
Je1NUVh2CtnEe+CB4/zZRkQk+vJD05N76TeTqQq9NjBJmVc+AStuoqWF/OtPyZZOFvhHABnIGkDx
L0p1x1ceMdYQxYp6URUtiK6ng6s6YkvHKANlHA5NzxIbu6uwLX1nIdGRwNxtzlRGpMxvSVL3nA4M
9uCUSz6ASTx1drLbj1zok5zYI3qMR8s0dMX2hc2A5/p47jtd9Be1Kd3meIQgUZcqTLppcgS9Ih2u
d3xEF5FLpbg/AUik5rSEOsKA0fYQhmipBiI//1s5o8BfGBBJB45xv3CgQ8xwl0E6yLK6bRJqopy3
Ukp3d/mBCDFPunLkbkuAHUAjN8GoU3SdeGe0LglDHNHtCmxVjAoSv6OTNAbv34qG5dp3uyEp5GCZ
G9cciu6nw7Lr3uoyD3MafIXYt5CXbwkG7otUCqrJR+jGfWFrkgMvuRCwt48QthIFcTwGUlMnYHX7
2ARDc6kSDxQFzP804V+3bzMM7Y1W5TpK0dAIB3Urdga5nfyCjA/i7D0mBgxigusMgmPp6PPzAJrb
zCPXwok5BORAzN3z+bjFc775JDad7SYcegC8TbuIQaArPN4h/h1Ttf+KPLdB6a+OVfk85iiSf/sY
LD7iCbFNHRzpvtat7NtdfKG3nNrbX+3ivBH6xYxF0UNeWhvec65ZQXY/eXzknFGucdWIZ9IhY3I9
g+U9/fHttwqxCkIhVoPMj5jgaCPo7jOSRlS5xp7VBpEhtl8pMfvN5ATyJv+B6MzOblK7z7QvnjRt
wC0P/a2lysnPnGkxUi4Ix/+SVB2Ezt0q2eJVZtOds3sm9Kni0jlU+saz/XU1yIqDlnfsB2h/H2fh
PtcT1Q4ufH01e+kD89sc44hWmxli9GKPkF7AeivFcT/LdTdQc08H0Sdzbhjn90XBPNwg4b6pijkj
tca9NVSaVAWXPA/kbwStrWCpCsMtXG8L+WMOxJ+zpSwLCs/kVX/H1UbPdTxO5484qLFLcPspQr9S
dMBMGki+dDKaUwEcfTpQWjaoBVIzHbq74zVdwv8jjd7HHOQthvQmDd+wdNd5yYuhiogdJnDpDot6
Fk6APRy1w7hJu1HuF0RZjgbCWTpiL3lPuQP2fnSBaHlboqwCspKO3mWSZ1PK2RCVZtON5IILSQjs
Ko8YQ4lw16uzZe5BolIY0tKYBdG/enCP2+jx/00cXMpFVD7ROFFhwT9WLGjfCRw+NlLKbUDI3sfV
6zqxpCeorM8T5OpZ3z9nxbdBrhaKuIsHBwbVbazaqadJZt4ZI+cMB8HXA+zdktvFVUXnrizzdjfQ
7/8Bj+f9bHSVvt1FyXKzImaXI7mP6cK/WJqxEIGgnw3wW2jeeL0CJgk/euKPzTdZhHnHiVZh+VyB
zVsZ5w7WDzCBCozKbyYU6/+/PIJ6L5aXDLlgK+3iprKqMe47TBRYoj1lD65pk3BzahW65zCWb6F/
JbqGt5qPcAU7tOb8/mQVstdoKpN+Hyp1b+ohu9vYkI8XwFKe6Vwude1MyQNaMYB0F+jfpTTMGq2k
xjJxwIkMZllnBC68Lg0HwSPrgFHzKJenYJsaCh4Hm2ZzTME1YoKTwqOd4KJQvD/j8dyriXx61RvY
pl5CltCSxGknFUD4k7maVPxNa30jIoXueGQ26OWg0OPA6FrYvb31C8O6AlY8A9QbkZFRr97z3TFz
J69+E92sYuhUd345/+kW8eGx+djoxm3fCBNIdnOoWIt0tmDeikEtLSf1K9dwcaieCDf303VSwcY5
ZfnhVgKGsNuMBonxqqwrA4Qx5QeFH5GXzHET2dzX5eDAwZDhmBzPknymc+O2LvMh5aJkt5py/lyA
22Pgmzfz8FmH7iNJ90TYZzP0E6A0OPbHDIAgXvGFGA6RiMvymHF1++37VghGulfaah7WDlb183uw
Qhp1/0e0b5csVDYD519h1MEyNVVcDF/aPOHVR1l1v09EYL0Ymt3DX3m7fJdsEzAxn7EGsoPqkrTy
JNWvnGShC54Zb+sTGJndQx1hMchj2BcoCGuGHyJymMd9MhSz/d1g0ASPvS31xmHYtFz4POGGlyo5
WKVAKKCbswiRjYTgn0ajIYH0VoIbO3Lwu0f9GcKlEMKSygAsb2S5C9MPqSxCAD0EZB/hDNvKLFFG
2HK+hm2YxmZ5A2YHKfWm/FDsDmXgtmjPw8lKQfLAYugOEHqrZkgKHw+81ZgRMTldPQs7AiPDkJ2w
3xHBHbAKHRzesssRSwfzhM543NnOsBDcJIKUrHykH3V4DWQiGWD2DM33zFdPP2jJWg7gm7CLOOqz
tTc7or4MAxECyiYRT21k9QWumkq/WnBXGD2eMCc8+Vg2HPdSAC8Q2P9DjZ1K97UdAOUYbDrHdvN9
7vFz7rFpUzsBbFUK0z0A6G6/qrY1TuamgX52cooLWgx0wI4SOHTdfZ/YvlSC/nvmEQUOqk2J9x2H
xwgscyK6e8uypoUJXJfmf1suG4CMEgRe1kZo4o93VNai7xEFp7GfhfIx4WlCR67hNKFKko2nOIl4
MkMOfATzXJ8yqozNHZyj1JfE6FqpaZvCLLk6kGHGsohWkDH6mNX859lQhU2xM1QeAz26pwgYFh0q
/FIhlULInjyC63g0/CA7xOpZpmQiFgyDxM4pbiWdLy9b1GYyd27wWfjCpaW/D+h8DzJerqm0Gu/q
pQQfxM77coueeOtxHcFmKht0sQ8EPx+gIcIunGDIVwFSaPYlHb7cfQjfW1V3Bkvv8JdXf2A6rHdo
TeFWmWCn+koiooVjd8NTl4x7NDX+fEv3a7P5WLGYvLTKYH8zfk/fsNQetgrzookd3J1VmvHtwOQ2
1owwC/ntKxaiOld0PiDJsYXQ1RGk+fEvPxI8Hc9+A3qXVeydFOngpk5BNnwDGYvEXs0fCcB2yo2G
Z7IBxLc8Wqr+PHyE7aSI7dypKMuOn31KVU8U0nvUwOlPzKFwKivoNEGESH2z0JoadcV/LYgr2tIK
NddqV8SuSCJOq6i6ipKi3UPCit0LU1S291EXDogI8wU3f4wvSNUnRdtppASHWGVq/V4rcsx/j3J8
/gD/N47QRBWVFZyyMPbblrCGnsNP9InMi5rAxgz41jtOzr3t7WQRvD23A39OzDHUu35xMLmMZRPH
PM6YQzRR7OqKgG67EfxsENtin58Fs9RsUgZkeU5I0ktEz9Vikxc7aoZ3Z0tDfVfXkTpMtkA4TAG0
hCXPVlD+xKjakCxdL1pKRW2/Xgy0U5J2jeO3SoQKy3mCuSxQt9fmfTx4ErH/dnHhxLvgKXFwREUa
zb+a6lznK8UMq94LluRq0BIAZ/TNLabPBwCrWFhNVVTsX/xtJCJiI9E2faLek1s9Zfb1kts8PHi5
wqFIP5651eHYq4mWJ99GV4aGkB9coUFXhjMLwB8cG3voS/okRcOhQpe5arlatg97Ie7C8oqS8Lsz
cMU4vXHbNWy8oQjA0opw/KRQ+ZwGO7T8NUKijOMaiITm3kZzlfleyXZHFfMVJ7GHphCaYk+1OWLt
qWlfV4yMK6BglWaA5JEQwLGxcskGM4ULTQUHQxosmBUdJGDgWwnFPSj5QFEF7Y6znUwE6sRfrmMT
vCq52f/b+7ClkELJOLfjlSVHh1MpumOzjTYSfAuZZjettCeE0r1fHcHPwtyI0QlgMaC0sJJtDcd9
6SExlQ15lqV2p3cqkxp6Tebr6fLrydAeONxq0DtvG6MqOI2Py665PpASuA2UVvk6VqQCcMSOgB2G
Qhn2hayPNCckKKwF/53ka1t590l8gG4ofg1q6U3uEAqd+s4PJjyuRirYodS9KyHOAo4FM+xGVm4N
VgbGdC01TA4P7PzauK9fedHJc68NQlqsbLVsQ5iW33RbJeikpKJhug3TssHAiikvpgitHlltJaSj
URbuqwzCaHmEL29GfjmSx2NdlBwF5JRS+bUn73JD3fyR/WtMKqL0GHU9ajERnopj+rB/xQh9GWox
hD2ei5gX4kSwQdgtKXo8cU0kXv1bTJLXxN7p4fSYPRQg8j6SMWQFBEAfz2HLuYd9ler6NW79yEQD
TawyRYMUVQtgjp4kZJ8UmRFJD0VlI3DqKl95tLrWIOd+Ofp+PMRuPBh2CS56QdVC19sm816LX+m2
LXmYQUCSYumVq+XqV55vPma19Pya1NGRLAHLCHnW/z1jNugtxkIWowmXclAcoTkLyhbs8bVYrokI
5WLVRYjR0ejMFVsLg8MVvejaTLNJ07PnNVA9/GVmsQecnyInXr4NqZMiwhOHKHtofHZ8+DWAWu3v
hom3a8ZOY7OpxZje1eq6ycoNMVrfFwQyqxmyvFDA3wKxW9i9vjTQSXfeY08BJjmMSlUCZFKZQLDM
cbyks6Rwy91suJzDFHtnvCGZwEd1TcJfYqBOQp5mUTfrW4JkdGhSt5qXfJFw4jiqrflOp+NXFjY+
E4hAiHwAJiT+Nc4Dcmga9QCssTJwT/mA7zqhsRTZYMUV7u8fVBG1zU9z59+wAKf08sJBYyOju7IQ
wH71FBfi6sMNQdBZCGgj/durXOioCWl9KQAUln4pa4jjDhGBGt0pyvqynv6D3oyHmdR26n8Ysjn1
0penZdcVdWntSRURSZIVrB4XZIk4dhsSM4LxcUI8PslJuh5GERMJEprgLcgFybGx2TtdEv8hhQUi
vBmjRNjRMa6vWCk/6r+uK3o7IAXknzLHlW1wSKdRhGvaPQHSVj+qrGXfD5gB7q6YIuaFxdhuUNbE
ieEgI2bwXawGY8OVDNhLn+T1RWq2WEEZJzDHMb7xcE4kSk04P1WWYZTMi33UNTel+lgEl6BJhqbP
XX9auaLmCVpQhiqDY4Xy42IErHcKUTb3tKYHHip3PuJSvJR+ehm/cw/A1up0DP42Fhe+DhEyrfF1
j78owE83SYi+p54PBhETrSNwm4kNukClY0pRYLBjCJ0xe8Pmx9MF9IevzYKBiSSfajJTTV+g0YRW
+4G8VZRYZMCHw9KzTYhrn6uIJyqGPHPfmGTxvcIydLcDc5HY+y9BfwZZAide82Gl4YPjfbGbYUg2
L8goQGSUxFal+Wqr1sjBZcS24Tvq/BwhSfE+I9el4Er7Y/LxAWOqTV8/d7kD88sP3lVdsr7MXmK2
YirLzUyxqjhelNamIvAuuTu88f5jGmGeUzcWGb046JLigMGFjihoivdB3a2WrQiAHdL7Fnl/0fso
I8z6/ef+CHKcdcYl+UxVy4kBKdDnH6KSnBo56SQRy9hpDZT2o0gFPCmXCV/hITlVqTn6fGXouH0J
v9yGF2q05TZXKHFyuZxiMCVf9QqoqX6Pz/BjAaqrDIGsWZDJwvyKM6RhZKjPJUkIPLeMGeW+Bvrc
LgMM/E6snUIYWB/aLIGHlfG7PA2/PDHWmFji78tcYB0O3VGHLUEkrKpY6144FLl2vH44vY297MqC
Py+rUPWtxwFfqtel52PYGrMrp2WyWiemi7go34uQNelil4ztmF0EIsyCtbcOf7/1RL7+xghq/Ufg
3m+osNXKdUMkkPKyoFcOMigpxpDyFfGSJ0Exp4ssJfebHO5ET0up1EaOCc6gaCBRNSm/YRfX/lmI
DyLRfYO0kXNClyePYn0NMlEILol78ywM/7vpWpWN1nfHFvfIDomyeFY3XxS+rspcAVCOBamKNIdj
LO6P3b0/ENG6fzoYnvTsJ0CoTro27I6K8GRCzXs+UQtwhFTALs7bqXrSw1+VoplN6apkG3riDS6d
O2iL3ROepZG4GvLcQWlbcvWJjLu02l+/mLlBXtlXHObCpkW5/f1KtxXkpnPYghJhNq9sYtg9kd50
81tYq+9UGPLsROjHmKSpbDLhsMHsYb7bJv6g+3+6CkeDtBqT3yFQoqSwmP+ERwjJK18OLoj352vY
SdesZvOL0hJa7pLS7LqIRYtRpMe8ylejw7pUDVVh7DYLJV1lyLRgj0Mmd2J9J9wppRWdZXRBzKol
ttRU47eZyc5vmjT+7xV7lPKpT/noD1cxDsUXuEq6slI2oukZxd43kgzMZDZmR6mwCtTH1x1azZ9A
iywn3Prr1wTFPfldPwk0vhR7jwiaAx2I6vKatI95JK1yoogNcpe6mZkY8qnI8dNRZBN0DQ1MyCv+
L+fOjumg0tKzrtr+Y5ojKqZ6ZXF62oWtk8PVoHtvutGDr5CXei6g9rjfgxvJRVLJupsQwH4bSFTg
eUdGzJtPX5S/avwQfHPBaqG0mAC8U1H+cH2742gCHw9U2dT+OpB8VEApQWe0c8fF0fg0C7agRdyY
SmWzg5qechNYvRlUwaObhlkAq9EBvWbU5IfP1A5TNTa1y2Ij26laYt96KmEZmXXmgiGJd2OdoVgL
7X8tED/jkHrZQM03jampuHInooum6fy9+oalTIZJKd9pXfaJWTiPp8i7hZgnFfZ60VW0rool0zQ1
EJoY72DFPb7t9suuabuqQ1qhdgGZY0KOF61FSEmsGd4h6wyz6AS4waFoQ0p4C3y2x2nurMC0RBcl
9/CGwvwAcAf8IgjZwuw88GX9SsH1sk0yLYqE6FrU2PpNcC2IXvdbtSkvA/rr8xwIZUghfwrsgMxR
d0ScvlS7kE56idoXU/jlFFx7xmscDDisjK3i8TumgBeH6e/IHRwwiwqz9qUNFOECg9Mz5G6/o6al
30MtHzFnJXlSmuhbT3VMHnIb0TKU8QMZ1zw0YgMN0vQpf9DQg84tGgQxk2ubGk7j/nmvuwMAnmYJ
igSMVOv8Zsdjg41ZiU+xXCYDdQXPIXL3cGVsKI6HIdTTcWXeAXwyF5onDX/ypDFZ86oipNKCuRQj
8+P9V/hXsaBOSDBHzH9NBrki/VluvYwHHo+zI8YJ/wpuVB0OLWw6bloWUpq9Ii6z1oIxvRGFrF/G
/VblWUIdk0iSep2ow0cqxmTRUw1yDq8yEpuyScKj5gebC+K9I8RrdkcuYL/bQ2yVFqtm+4ckhBhr
4Qau9CeeFnqyQXCDnuX9IXmu73ojOJl/PdCa+UCc6uW4wMki3Vnf/39WQz0cLDm3i0XKcZpsFdm+
Q1mz4PlNPVmtfKeT8GLASz/J5s6+lRFU/1rr498sfLVgRxxxHhX5WhTn96YadycKPdenisI6VJIG
qB9rE6h2BkpdMAVl1nvId+W6Okk/AP1g8w2h8kERiwH0PYooEr5DgTy/MpT8CEfbaSdpWp3pxytk
uTc88AXL8wadG9yvIshMJhdFiAfrGrIwBd6KJeCsVr3LKmzQ0oSQgItvSXdQdmBY3EdgwaDy79aJ
FNzY51kSup0P6js+zVdhrMEwcXPVkRvVvul3INkN2KhvCJODM1X83CqBH2PAZKsI12Poct7zgf7S
V+4XMnvmceZiM0qi1JGC+ObZKeaMUOaEsqq9sF1X67xASa11jIlUfPZmDKNqMDxaRvV8Smg1PS52
4bjUz9l8MaNJum01HEy+jupVjCTsMoqW0XHkqY5+59jSOHRVNuvHHR/SnmieYn36WyvOZTDeI/8i
NSUwvTTmp4bGAXcWli589vfhdo1i/YfdMEtDPeGv0NXlQmotNRN3IGsTyrgspiKsmqkEEK6F0Hzw
EnsGtnYnaX51p3UdbiBrDQ/QPipwQQdGSLEnflVaUK2wKWgSm/37b8OpxzQ73CWUJssxIzoGW7up
jvCguLUpDGr3JfrnCsBZPUAibLhh35XHy4G0qjPkS/z7lbWqZfLw3c/FUqA/agequaZiEOp2VPMj
ONJ12Xq+59Tm1BU3ktSxkJaOta/LIV51orKfuYLafJafu/cG2m8EY+pCPls7NbpyZZ5oIAftpK3M
QIhPa3GKWUjK+gQzoa4fgqx6AsSLxIj7oOeLnB5rLpoBLAKaSXqZsogyjZ/dggiq5Y61CY6MUJGe
28hT2x6be/BMYP3+W+8av6IWZGDpUf4K67q7KCLzL53B9Xcm/Uf3oVjIoO1aO8XNtiBj4hnJ99oq
Ruihx5tEz+NcTGGp89O+/ZFYk7uTmbel/UycjG3di8fQOk3RIuhxNcaOMZuIaFIYl4yPOmghNeBV
k4IdFaVWLBdI8ucUo7xyU1gnb5oLmlF1enKRoyzL9NPn2oUZj6n1PaWaxSJxx+o1wEYgvCgzLWKD
VVQHMCB3FWjdWOfQ3lnoTFIwuhZmFIrAkwWDfI6jrRD4qdOAtE1iyCCOj7Wx5SOhU7mwV2Lo3zdX
460LAWSaZ9Iwslx4B4nUiPkcEXBO8soIPlLZKMTlMsmAg+oEi+ddvy5WVBZFyYDPTJNt+l/XtRfd
QviL+lkt3O/1HtvtxCmp26paTuvKsoiWzLSlfaYgfNuT177mbELzzR68QTk2W7F/04MGCKnE7uvC
EpjLQVYNStEpBwCZ5pwmQ6J9ba5swOTRrDvQSx7j4gvOxsA8HG7xErlAAd/LPXpMivEmIF5/JNVa
QtDvTeZvx+605kgsGLEa32cnUg5eJOPu2A10rhzAqtIbZq7G0EU2xXOu6Fwx+nT7l9CvspentnIy
5pTIbc0MSsYE+bpfCmQS3vLCl0aZgCVh/SrKQ5ZBpnAJqbOYYvatn3mERuB0qVJEYXGy0UiUlYEZ
e3i6h9imIpM8+8tcf9L6C+ZVeyjhVZX3ghaRF/kw1/SMzQ19U4o8Xm+TNE4B4BqlX884QkDn6Gie
ivQbyFOIrGlWX4gtuduOAvZdEalWDeTEzi1jdMJYEMvfVAgI5d4SejKBtVwEbFtcBkwNB0CgvGU2
c9quJta9WRwJpXUDpl7KpifsegHJg7wZkhaYckvM4ZcXUkwuou2ecinm66c4huftk/5cdfLOy59m
9mHQPcrW9AWcocHb4ULh7XsEBEJasN2/rmBXKkp7XlhUKarG6sMyFJ7ehvBV8fHstY7tvToUeY27
olGCBsw/q9eoOxlp2Uu5Hvvb0c37FEFRAeZ64g7gJgOdfL5ZX8bml3rAbPxuOtEz/C4bxMxYUkC0
aMGBqV1RRJkAtW2/o3swW+/Jv8v0GXJA6IA6jX2mp8DUv5rkPgrEojGn2gF+hfkh/zyKPCx7ptYF
Vy3QfztvzpD/wskPVBcqZFoA1KxMEI5KCYdmiQu1YM+MsFRmJBRO+SqgZnh/OEdEHvX3IZ5lK3xN
fOt+MNSZb9GiIzR+6Q6BmJKrG4LKBb9QnVwJQ0lG/HXD9y74jj2Ek8BeSRopCsZ9zFry9oLGKBrd
1smLIXu02Rsnm5xe+vKpY3Q7Jy4Vzes259dRGwi0CD6QBtdofpyGTSHHUIBl1t1r0NzdIVjv0dWn
2iFQO8Dj9k27JnGaJxwuGMko+CCeaopqcyGE3vr0a7htjtHH6xrAVw3AOB5FWZU2i3vjWibk0Khx
Bs4xm85+xlUiHYDi4O/JejKC5PlZQSr9XjdJwjVJXFxbqGR+rgL9gt7dS12It24HDPaCStNT+K3j
EFa8rgJUnz4dp5Uh5Z+BPXKfiQAWvoEZczTzkawgVko9GLPtp1P5s1bmgdRD2jsBsMUq7n2d11vO
uxm3udZpNFLqO2OpUO1psBGCN17uh8FC0xq8xXLxicVMow/MARZo/nxOLt54kLednzKFUcU3ReRq
szIK5LjlUHO9oFoITRsQ5K6V6ucDq1T2mO7hRW/x6zh2kuR8jLvfIlgTRKEZYEiVGcxXQtBhEKdB
hpRu7NRLqm7J8zmjIdHQTia798/norsISYbzmLZPCvpKKnRtMxVqH8t3F/NeL+g6GjGolPWzdgcD
Va0c7ryJ1GLflNAkQeffpeWr1eULu+KRpOQfNiV26XxRj0puPm0ewvBtuNtfupZWGhtJXIghegDP
sW49pQrHsWZ6HvjM8ekfnAjWJqDaAC5tLjqTWz+rQHuIw+7OWLoGaGwJTFF0gtD5xEu3+6UxyPiZ
r131RNPENYF1+xmYzzTvX/ZUPaLA2MZobxokbv6cGgf9U72DjAXjEgDMVof3p3Oxg7XKxRFNMi3G
t4U8xszgEU/nqvUFxgH+82DrOXjGELGPNU1OgxKjS0GioQEmIYPAW7Cz9svJxS5nd7PdiwtYRBGs
DxG0CWNBgRdi+CRxwUoqaEMUr0B+PK1gGA8F+kQhsMuKoZo2RwBqYaO3zp9oXauuMzmsJJ0l2Ypv
UVDeBt4BMdD0Kkz0XBZyjVnkpY0oPsj+wT3+TNXgS9BJeuqkZbYH4pL+LoP5iIjsKuov3ND2osuK
7RMeOjes2hrMHpjfbz7VXt4eH5avTZVyhL4Ro4jeDN9frweHvAeauRSZdfmkgRjgk4X/f5etn8a8
UUPCLPkYXUQBgwz8lxhLkGrXxnwlfRb02lAYwcJ8H1X4HFKJK6OWFA6dCZ8dCWIdaQUwoGdrw2zE
TVbMcimN/1YrLoioOu/Pf9+U0DcqJ3JXwzJQdjMlM5z2ieiQ1tqkB4RKuYxKDRArtRpR4L6bcE8K
qPnDXgOCwXOTb6amf6OqJIg7V6XmbUjvdwEbkyscU5X9SHg/5lPIFmoJKbZMd/diLM0hLgxrBYSH
Ha3WyIeDzNa1J0GOtb5qQY9mBg8zdBB5t3lJRJ9/X94+NIz+JMPAXbUR+oOfdxeSwrxqUjQc7txg
F24GTLJlfcsKVbzI8H3MUl7pPgS15WtDg+Hoat/tYc+KMJcoa3vgZNC34Zopt62t6oHm+acEIsT3
q8e4pTayWHc979g1Hlr3K132TzF3iMA7YnzKlMEZmKU5kIS4hYbYZc+QI3rccGVrsLHFqVTCaobs
gnZQqGtwR6xpnA3NKhrigdF5ycksJccveubfWW8ByVQWW0H1HRtuiQDBjzw2csmh/3/uFMPNczDT
aoJ3cx4TiPuvkqCpFy2Gmbs3NkaoA+Rpa7Ey0SLMKU+l67IBeM6kPX4iPWvcnrf1E+NBLpcf5CED
8Uc/Vh7nsa04q46H2sfLz8V9xteVGFXVNEhmXXmGF+sDb5dbLRaqn4SGgrLvPuisJFZAX1GSz5CM
KtIgUYOHZnD7y0sz3KV/3VNq5SKwYiqEHY4AjIKgoUPMPbs22Jdtm6ZdJJpq/d8aFmRsmeGnhXn+
6N7WDGofTDnxrAW/DR/6t8qTSwQkuj72jeFVl1xo1egAgIdIICC1VPkD3BsnWLo8TgHwn2T+b3wK
kzm9taPgbrENTAnNsDHUQPmQKaJF8omZWTbfkbybhKiKVqa6efHHwcjgsdThzViUukLA5wEXANJj
qANpZSox7fFZYzezuiPcSDY2/5lsNADMCeOCyVZx7qAI0dOJZ0E2r0Mnfq5PTD+DzgOeV8SarGu1
urm6Ra06lRmhQgDwD3dzPsnvS3hM/aW1Nyif8lUmQqm54cyOGLQsrE542LGb4LTpm7Y4Rwjcllzc
oZgbXGPYv/3y2hOYFxwBoUKlZwAKa1RFEquDir4J3gDpHvOEe9ZLng63lguLZDBdA85zdKzCwTyw
EP5vZv0=
`protect end_protected

