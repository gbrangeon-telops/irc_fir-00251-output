

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Syf21YU5JnKptD7LOLtaHZM+q1VIhUFTxsmS2r0ofwQ3ushsF40KxXOCQsGAnXjGfc9kVb3Bn0ME
1qO92hlu9w==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
dY69aEX8OSz52Pib+7B1y1Wvr7162ZPVuHYqEcMQ/oCfJJrpwF+oy+zQI55NVyz5aWKsTxE6uM7J
HbTWuphJFeGo7mzwyRD7dy/8IFTp8OHV9aN/fKWepd3R1nKJ/+bdmSsliOOw+inM7pfx0a3YODTn
FRAbVAMQuwe+OVuT0dQ=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Q+4W/1zvXVAi9QMds0GLwNMATdnR+yvz4Aqge4tYro137XvQ9NhFGdF/mXOn40o0ijOuTLANSGZq
Y1fe5IvAhv/BzIqGLvvBSGadUyLWCe23JTco14xHGh+EcGpkQzSMsD+MtFlsKB5Lh4Pk7Fki+zjY
CYS3IH1yrExDySGaxaJ/xIpVmbcDUIB29ts6Ape06rDNuWSEZkqi5ATlUPCMrVpXs0LgVRBipzor
Mr/lCisQJrroeVDmbpQGOxCT0USTTIePtqKzCRURmGOM39JzikVR3QvCxX3V9zs6LEiHJnsAr/WX
JYHo8e0tsbF+S86/2TJe/j8LJK3VvghHADCdOg==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
jFetHSEk8pl36rsszcvK1lxgvI24/D3eeWIqqx4SgMWK5zMch2RGKDJVjZdo+SXrQZtG4vIfoNJ/
M9NL/crW7IJ+pa4Cb2wH+GD2pA66Yo3aRE1Ld7EknU3x42o8aAXlhcPIjcxq9tmSO5RxnhMKlfjh
dMPsoD+Mezyol/EwGPo=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Jgq62sziWqkTYcR9/y/ZRFUy8fWL8zR/UZTwiK9JRpmOKe++dsuUuVffmjjAGJoOkGM1fnXZqKj9
LDnUvlqAYGJAQrwT7QRdCNBN9eBMyr6WJUCOkpNRo5aWbRqVpwZihLgqtvesSbzoaKe4eDRdiEe1
xKR9vPyfNmAnPN1pwf+2YDUftVl5x4CmlqRUCO2c3iETzT+xwYzxqYKolk4Qa8DTTYe9PvjYqn2/
dj/jpAwnTcOKUqpa/3FaAU1zgLKWphnnTU+MOfKNP/ow3ZLVrmyiraKTGZlBmdJF18AzYgHb4rrc
8Z8DuRLa762hnT0qbzjf0vtKn06WBHgWqansQw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 19248)
`protect data_block
S0eUOz0l355zDEfNvwjnzPml0juIpac7KiJ6cjvumwJmikvri/3JwMfPZyRK42ljfJ2p8SSG9dp4
jxep30qi1wlW/ZBXGSKpvOMPNs4OkxIcECoEAz23OdQrtmGS/WVQL6vL6rVSc3OlTI0fiQzstpT6
gAGSDakBkTajVdZx8ZS8hSSy/DBNl8oiQk55M7tFZpgtZ+sM7/PFBuVl4tKU9LV4VQM8XkXIjujY
Qib0a+tr7Ncoa3jF44dYIbPcht/PT+JPakFtmZSrDCTT9O9ZBtvZX4OEZrn/Tu024wn9Ptfkmg5H
Pvq97Xg0H+UpatLWZSfRaz/HATnbPsLDqOE/tkEdjukqtaOBds77gjiOixys9TJski/hkXorLvZW
lHH5R8ANc8S7gauJZJupNnTAFFeBMOp5/unMuiNg+210X077iP4aff6nGtWVkOn3xnn4uYv8apmG
HTfU4bB4bDfGVfui31mPL5AKYC6mga/3pxKIU+Rv9EM1b5+btA4utzVznNhJdfh0st4SRiKrCc9X
sLuYu/QvEJ3bvwX5iX7ewhxQIMvK0SvbOWtceDc5c5gbKQXPreJCW7a3XayG0tvs6HocWdV4ulae
t5AEOREIXCGdSOKLUHpJpxqmR4Bzxc1AR1isXDgWahaNpxbl24KGJIRWbHYAQcOK6YNk7jPiV4nU
G++QsAL8CNkTsb7h85RMr2iiVozlKyIQhlRGiaLCiz4MY88DjmebdXyFV77fWGsfK6UecL9q75Fq
eYj/u225gkzRIrAe3/X50rxChFUfhvePymYBwwbvPAzbr3aY+fLpSR8WBrj9eWD9T4wD77Ergzyz
vtu1qXuaobWPefKNl3L2eaRLmbAus4TzDcj6hnEF2FcZ5DFtJIwnrRsj2KNZxB7qRj3BXj7mp2Xm
dmhPbr7smDGLDLVzkDaW2qsiHLjhHWLLlAS/RWue+aaDRd9AX1c+QhB5Jn9ftHZBKwKuB7r5ORla
XZtfW+PffT3kzckgzXzs66DcmkTff4AsixTkvm3ut6eLsA76pzfOdTWpCounA/ciuEpq8jwrCLJs
k2vuOdGZfcCOFcsGp/V6bqc9bIILBkji3WTwSBTXFBtOh9KSJXFjAI1S2E3aHW2YX6rjj9V4fSBe
+2PIwacj9p9TweXeJuF2479/lbm5qVeQn74ZcRl1I7SXEX+bpK7S97exGgyOxaymYni+rPTkMv7a
oM5xuUg4N1QiHwYUqabYcIKgt/bXv4PBcB085H7Gzta9tVqTb6nSKe7PfwPt9Q5TG6SnrlUeWbr+
4MjsDmcXWm6Pi52OYB3LssgugNqOoq7Pmf3deKCa2Dq+JYRa4nHEE2aJja2+NGZfG8o4c+n/+H++
1G08xqw4+cWuleRaO5lu9qukb6UiuHcxDVSrDIo40w9RFDB7IY222d94BzivruCi+q5Jv+lQNgZi
I8f6l72/ceEuHntAlZiZvbBUZq2vtb4pEKYRsz2TSmQfkWxmWu/xq79s2W4633XgyAqO+8/5uPRU
Okvn1FbKjPUJYPYxaFQYPBw3fSjO68SDWmyUJs5m18AGtJPj7bfqaKhlRdhWV3hmII/7UAuCBUpQ
mj0I3hLtDuifiLYhlq8dFfkJKvaUECgKF69MThFRNqliAAhdq3gxYvjSr4ErNK4mDB+b5bnAX3jz
U2uXQozXVKfo9EB3pG2xFMliXEnzj1Bxcket5vBSIWcD4l7ftUyXLpH4SBM3I1izTW7FWjXco3LE
CuyskYQ352bSDL1bKqWaYy1rZAUWhtaC3Iv3hKrRiSxnkFZ2UMIhNyFVFG/wyJMDYfeb6Rh1NAwU
9yCkyJRNU2FBS7EKgMq8kGf+RU9RhapNj2yPOQSHvC46n+E2/ADut/fGmX8gZSRRxZUTmGvRAot+
hlTffGPIb46CZHBZrd9EDj4VS5hK2tVY+YZKO0snN+raaAE4UquQkRxnoi6cwBdzAlq+R8dEazIU
MzdLiljnHaTxkUelgQ08taJ16zEN1iaLL4eUFX5hGG/nC7zI/ser6ZH/ioKPGbiaKrR99hbBuenA
heBRr+3VXOhVfOt5ux8biTsYPkKOo92Q4r+88sbhvL0cezqqHQhAefG93LhEoUkTJrrAC8qqzpQw
eIjneo5yShuB7cCm8ZdfZGnMMy+fgGn4NpN1TnT4F+40Uv/AIqm0aD/Q/tXRwCdQj95uXpbR2yvf
obXmHSDyXa4Z8xqLO2QNImgJiMT5MvmkNn55duYgbZW6h/rkCxJT1beLmz4PBb/g1R/gpvQO9pER
MaUL/ihLwHv3xTS7YbAmVcOV/fbAc+Xwco4tNlJB8gAVBlnp9IhGtYjpGW9Nye0+PdM5bw7e1wMe
1DVhagFG4XAPl9bVJjdAFej793c8u0SnZqYlUvit5Q357X4/xwaR8M8gTga53TGs0n7HCWBeS1vt
tFhN/fK+JUjvQK77uwgNp8cwaT6/+BbCs4olWMWx2vFhAmjJ4ZkIDPHSq31ewBv9i14AZGGAr5p0
cTAITQbl9lVAAZT3dDgcZ2o4W7Ity5u4OdCkI9jBlG3/TxZK34GuMzAgVg2+Y7U9rH7bCpwS5VUo
9O0wzcffDqvJ0x3312sWSLqFCopXDJXF0eGXePs4NwXAf0WwuytfEWce8tgWV4vFkTgScRVJDNGL
d++9WUrU1dhpV757wPdwAkvBKCBN8SOcVAz2zjiAEEtpi3ZmaVJjVy8UOLwMlMGCQAzd7o77xlgu
0XYXOufYN8kS3p2WAUsxHoCRo7bIO45O8qNLfj0vye4CWoQX5N1z4I4esND7I5WeVFfXKtwsPh92
ICrCEJe0SssyohtRlr+GCqOUlxjWsoXsuJe09eEXzDa1uKlvihXoMEPAxY85v1m0/ngPevq0rY8N
zefkILlE9+On8wKJ7m/SoKVAR3/fvViJdtnVkC2KIOmcP9FzYN34wmryLjXXKsyRC/3T3fkCPiGa
DJ5d35Tk2wWUuvM7dcC+0womkayqB1bm0c2q7glq/2VTYhnB82mivQqdkU0W+JO4/Ppfri9TCHJk
vhIw8blVrkGexdRTZ9Z1rjceB66drSNyGX8xE4Mz+hlYS20FGeMix5kjCSFbL4T/9BJnKS2GBA0/
aLnuX8i6PiFYtrGKqu4G4AGLw9wmdwM7xfDVgck6xrc+eDTa8bPVrmDls7LLmAgc1e0+HTK3vdJu
90ch1f9ygbm6nF8s+gwd+DXZGiEoLQA5z1uLqqlltpELceah7nOJ6M7HKIrsM2egI6jh/PgPC4/t
5q0IfHJvj+Vb5qRn3W8FRNUyfw7Aw7gRsLzMrZ7aKJLxQun3xTyJ8Xgt3l/AlFxM6Yfz/bTWxmPA
iabmWjbiQ9sp8YyEy226M+HWbvfSQOjFGTErLxOc/DXnZJYUFO0pEVaX0PUgoPp7ZF70vVUKKcRR
XhlOf80jfQMXlQOvkU4Vmg4e8uxJwRFcQyVg1lRvhGURiC+puYHZXxydTu92p9kLlFUAgEVpkAH9
My88fXNDIcPVsK8/nNN/Ux6RvDRoNhiZr/JWh+zY/IOJamCOtoIKUYlczaDMD5wKMsPMPnVtfLV2
vSX9meBdG6fIVA7KkLA/mIOcz2cXrU2GdhgsuYgfOn1v+lXkQgdFmyVAIKAoRa43QEm7AIm3HBhq
QYTFGo0DsrNYI3bSTYezaI083RVgwasJgPLQC46nrj+ZFqll53mliin7pd1RKnMj5RrNFFL028EX
FdtMh9dTMmntfXpzONAon/gJifcohozamGhbz5XUPBxQAEDaQ5usltlqIPnQ/Q2T8iv2J7NlX2me
RmH2pq6YqaCsGxcRtzbVZfmeOxIJWMzzDzH8Ng/GdjmySKByrtqsEtrahTrVi066+ciyT12IEXKn
Ssvm5nProRaR+K6lLkzqKUUqiMkVQ7qNB8sArQCPLJvMAsv2Iah3hHVIBOW+o8/GF3MOigP24LoA
G/YQq8K1ltzs2yZJ+v2XV+YuOhzpLpCNlj0a53qAx+Jy05TYDqbWNAHaz3By+To2Z55U/rWtVjX1
4L7DfYEMo1g3O7VM8CMQhRDuGcuCL4pMeOxWflSIx+0PGFhD8MRvg2Kz8ozA8Q2CTEOdBQbcj5um
JB3LJVwnneXJyUmweSUF5s3y9TaQZ6eOs7kaAyvssAVFnf3yvd7P1O3eZkquo1ANSMrHdezoig/A
itgqSM3NbM57IDmtUMnfslO5uPLJ9EPCCloP+vt1pzXkW9t91Xqi7rTje0zAe+zEYHVUnSEJy7sh
l71pPVZIWCrUCQIJNoMzkULwrPN3nmo+TpI9oek2zAcUwek9fWiERNrGhbgA6eECYRWPim7oFTun
C4ZMHqiJEHGp7PfGoNofNvUdGz72omuCpC/XzOdmvzqVjA6jQdgq+pI8Zs5O+tJpHAKEsUPHQKYI
n6B7xGsjcedeJNHdtQGIQ8XqWxWvxDIDnEAY8PcqrY4/w1Pnhd5CZJRTp0hc5OrEX7KPt87kgecU
7ySof0E5gKabVxjyvZrNj3/pAtkTcohK6INQA9+PorZM+7RQLCPt2MVYjZI2d/I+ImaV6VWuk1Jo
nnsUlUQy0lgvO2LxUVOcvInQSbRRImLHfTT4ApWOrQMcXgENHO8HRX2I660LR82oYtpIsdQ3OoVK
Opek9fUKhPfyszc6TGNUvXjgvvsuuUTUzLFCpVTLT8gUc4Kg0LUhsXhR+WLAOEtC0o2AlDlfWh8H
U7v3cHtFogeTkRywyKPj2wvTYDjb7cfpj9nexwwzfCq7eASm4ctbt4rcAhfZRqjxeL6iVMuC5Ltp
zBL39b8VkD/7UPQR/DHCYnYsHXvjIrIo2My2r2Za3jp587gWfiYQlB29vVag+k3vaXgMDSXyFHlp
QtNPPKwTLrr+V5eSeDhnQkdQsosTc4eqmf70OphGcC6Kx4cfeH3xx8zT3/wKM7+uJSBlcG2i8dYG
QHA/c3dO3y642QWLjvwRMkS30HbkhTuN4hscLpMO4EkKxxI/cxbNu0xhSRe/kOfoFUbMh+0mFmOI
XFeKQBUvgr5/xhVUOcHFYuNZvuSRiAFetGj9R8NgoM78ak2Ebn7BQvl+tcEbIhKh9YdXEwDN1RUH
g3qPxRiO3nTIEOfIBLzrH+UnmlXiGVD6Wk8qm40KMyhamZbgjxhgKZjssdqJqWDjZv2wioQVXHGb
eXVYhaZ+X9jzBoCK1b75mHEP0a6QzOpZz2NueS/+i/hmoegzThDOCtYVDmRmVgtg/n8VwbpiK0vX
Q1xkqImZ60O/UWQ0x0z8Gt6NblS6ELq/F6X8Fz3xHDUkNObAK++zVaTXcHjCju9BPRCnEG4wK6ht
0e2x4x5YbzVovfjmKt9uVLIyQuXJ2mT1WUVxD8/PsDkeAdnfzU5Mhun+avRPxRzuK4eCaYZOrouN
Ai3mBMcnjW+JwwHXFj93YtHqEraX7u1Y6SlmFrjBnezdu/kw/RuUPwQDwnjQgNGJwYtcaSwkMOHK
On2nHs5Cc9t/WfgAbM3c9hKAesati3tE2zeHTwgruBMRlKmVNgz2hCdhC2mz1BkJ8LZlvNbMstxT
cLBo1Ql/Nzw4stOhLshMbt3wtleMMaMKt2SHlE5iMgS1dyRnoSR8Gm0sUFCs5/mIzwoRm8Y2QHkj
B14R/BqVMJAtL5bEhwp+iMyXj292pH1WfNCSP/+mXPT6g5qWkIrc6uO9DrGn8KTTL9/xow867AaQ
GSe43nSjBMZsnFlPO0v9XGQYvNN3EIQqJPi/RjIZJlQ2fjMxZeVXB/ZytlKU3AMpEbhPLi8wADX8
u/PnaFV7nMZwnXL0o71EI9pXk9c1ba96jD9H7SCutebp3aKlpFqTMQ9CcUALYGV+f8Es4Gy5boCO
S/QAbvWsWNPDQ67eepUVjLeidouanhDMyBr2v2OQJ6n5bjhvsfxrzukfhqjt41Wi85waZXblWXDO
ZdizzQxoau0Vq6Ssx0ICsXgjoXorSIY4B0niHWVpqswE2IeYQ+2PVFI+eDkiU1XtnWcSsCiEZJKp
28wsaAC1mw5wst5hrz2VCY7rqRyhFRISqoQ9mmg3KVe6461UiN1Jp5yKWPLF6HSWT1kQqSQ/TDlT
Fp2cNlRmoOrMd1vMWWRjGuSvFrkmuXq/1/HUTgirY2I70x6UJ5R664KFWFO2tiaolnD4rQllYE7P
kBP3x72zqmL1W8GtaAJ2foE5C5Itwo6Wu1kzf3UlEC5fChkDeQHabrpwUL2fhyO6eXxvVg7vwIri
/uzlUSbagrXiL41xBOog3fZp9l0q8ILcKBhfZZLjOoI+DzSihRuMOzXUHlJm4srLqbd21iy130lU
wlnDyWMUUGeRy8F7iBkn8lkxo2VXOMx6NPZcoS5uNPwPBwwRoC9nxOD4byYrmal3Dj9USZFROGxV
5l0NTDMTqkXkbdPtGrYiPYtj9euLT8yIJL3PL/hRMJZ1JRpOPOo7R/2v+LOtw9PowhCwotj8Lc/q
sOUVG9fUGCbzQ0pTpwnI46jjdkn6i1aDTmyq/wvNihj6NeZbOGL1f3QdlCVlFybfcyNcPY9RYjRB
J4PYhtm3MWIxXLGwcSRIfaKlF1HAo+Z3jqFYGDpP0M0vivIOHYm+NI7g14mLQ0FzMTewfF8UacQ+
p6lWte4nJrw1lTXDGteRkQ8yXzoipywPNgIgwJUHCUAZRTagU8Ur4n5foIkczGKbZYrJebtQXifT
9dzT1oG8bHohocHRe/T6zoiompmc1dDdHT/z7e77s4ToJ/twP+L/f0Wzkf0UIg/IBJL8SiS+dvSG
VVBZ3wJJQwshrTDSPY7Dt69yvLSG++flllvE4IRdXisSLsYyWW6Hd2lSWFOFphbCRx8ejGwWbKAK
wC9Kk789Ton0yptuzFl99CD/sovVfk4L4HkV6IHhFQmkdeU1KExyG71/E4ju5I0EiPIK6JuMOIV8
HNfJqMT0wMa4uHPnPFf+KYW17HAD1Xg5k5hmLFBt+xhlvyrjeLxfg5eeMSuc/IKXemeOZPTq2dn3
YUq4PfMWvkVISQKI31Xr46w05tvB1TDX+SDmmf6EzcarUbK70VHcid6Yeias06z+gUPnXGLAGaEn
v2y5/sKIdIEGcSgK9e3CQ/HK8KTzRA3GnEIbnnPXgfnbBPxo+ErHU5lBubkeQmWuh2N5jGahBSZI
n4CUNeAZ2WhfUyHc2cgH/SfOlY4xWMhWHff4uz4uivhnTJFm45pFg+g9lGB/BLzlaLdXELFC5Vyw
OwhACxwljtMiFH95pva+1dGAZfmvH9cYJrnWbGlSOoWNWhat26UUFUkHvwPmaDJFXTV1nA6z6hNR
DlpSWo9erV88Eh+fGeT4+oYyo+RtQVxCV5YLAhGVEBjBKwDdzBqstU8KG/ME6fv0ZwnUmoGhlU6m
ntXU0JvIjO8OZmRwZ0QLc/C07IZWcMnRv3zy0GUtbuNJj7gGJ/4lQ8VEads8eRQq/mtEZOU5BYF5
J3ZPktXkjn/uRdsYgii6mZ82dQqsq6hmrYX4l/pNI9EUrPZtcRcDXWfq7aY48wQ/+BeFaKE2wor3
VTeUjqXMQsO1WfFrkNRCuLBJwu9c8O/51vngxqKaBO3MVTJuNxteJTSyNFGlknP79EwMvvU0KfLQ
GU3f6396owebe5+v0YF3bfeDMowU3+PRS6ftbgCxgwwoqsqiBK0b3JMx47ixkMuOzYb2MU9wbifo
hCU8lKJZ+Va51aLYK991w31AVRq7Xs3jT0cAKi7hn2A7MyGD/rfFa0dH2+sggBRnN2JR0zqJU8Tv
mwymCWiANSEYDhvleYi/bl6QG+sF6TPukLubRkqnFkE3gRTjN7iUttJCOrw4RsR5flYokcyWsDbZ
PDQUmgCMqPrqXp1UD3w5xntIcibfZw9I/l+xj6D4GGJjgfq4S/dSo5HlDiswp0m8IuB14SyTbb3V
DJLLuAL3/JNOfDzMjEmfbLEJxdR0gNVb7cYUky/mu1rlsASy3jB07joWXEFUbtszQyarc8RWE5bb
HJLaHC9UNoYCBlKJHx6D85SzbeG4coyzZ4793LdsSUY/n453IFKzbTQmhb3Jae2cU9UgxAllQRlQ
wS75j43M0we0aGJ8WaLq/N+NA37JiaAGFrLab/r5AoCK6t0PmjUQK+GUbTX0DkoL9ChxQtvKShqO
vnaMUcn0CQW2YQSKljqRUKcRveKlRaoMYxB05hKhlGSsSYq/nLnstU4Bcb52JI5/5Bh/UWRY9QGk
qlRtap8oNCnbsBI66Hb5uWs9u2AO/yrObyUVp1Y61AmyxSvxKR7EMGcySmdjxH5TzhEDwR9B0Rkd
+H/PsAMSHFK7has6F2A0OmC93wyF7WdUSbaz19wVnXpKFRk6FqONHerBVb7DfC8zA2sKP2TBdTIQ
SvujkczsfbOngukeegjypkEaq7uN9x4Hg4x/wMVJkjbcX9h88TI5SlxtXx4TFEI5vnDKuQ8D7s9q
jAXPvzhW6woJkNFHgMdr+lZkR8FWjNnb00Z1sjdaV5REp549W62NFP/laGktZYVOPMUOQm2fHF/h
A+vQiO9iqib5kPaQsejWzU5eCckWkhaQy66j15OUXIB/mpdmD07Zk0FejGOU1BwRnQyBPOkMyNC/
ixlPaN/NRYqBJAIUsIn3dZC0Xl/c+H7RU45StrK2Qyd2J2ekJPceFh6IQEunspmoWscsSQeXxz/s
S5qkDHGIST2S7NMkWd8yFMySu4q44vobrb0k52xzSXd805DseIgMPjC/co+wdFzJGma7DRp0zU8T
AZqMqLgygV7fQYng0BsNVXtAHxWwTg8gdqO6tMUtooPrakUpUJyJh3NpCf21vY/4aNog2Q1eCD/j
+rSvuE8BgFs85Rj9doyilzX95XDbPwm9em6Tzzx7J5Lg2/qUl+64PlNPnFs7w/okZh1f1T7j1tAf
abyntCzUcIOQiB3dJPez+5shoIQWmRrpebe3Gt+pnwP5rFv9s6xvlvbGww0EB00HW+3tR0XkKMqQ
/5MrR4tCc1e/YiaBFZYBOrIpFt0+ev1LG97kgZHQluYLY7cy+LCQi+jl62GbThWkiuR+fKusjRM9
C70piO3S7GHrjr0j980T8Kdv4Atc1D5G+m5EbgngkMXXSw95mWbe1ZESkgK96HfyTPgj5tlJjBVk
UJEGnN2VZp7YP6bFlY69f57KrHYw2wyokXohEF7bKuZ2g6Gi8uQGPRqWXGWTTK3kmTw/unFBqrUA
a4oP3ukwlUEc9drcQWVuTdcK33N3RCowQpwdjrqMVnq6SFtgMvy1uR+sSPdP/yKjKGe3QG004xB4
8U6pQD/zkQ/bTTCs0BdQyE/O2ye6Aznivxk1wpdAQhBp5E8XQIoAziyuGP/i0lc2SSjyEhI0NK/L
DGi7FW0aJrNj9M0rj3ZvdWsXTYqeUkX5J4Aj6xS1r198SPetS3UD8n79KekvfP2G5bsPRKJAdhcP
DtYPBYHIMyU0cBdS7gGWuDUr2KSiwk/pUr97lszDj1mUcdmQhr5zFrjOMYjQJGPTGMg+qDnfZzWs
fRbjc9y5vAwVs9QOVFLj7hNlT+LF2TFm84e0zEFyZOmYyw6Z/JMPlRCAmu34CmO5Lw2gb9B2VhWW
AExG23Xk8Ymicl2VWqIWgu6tMFIecT1BChrP1mPW9nDErJjQAWMDB30li9BCQYJ+L22BTm/RcOiO
tRdXXcLhLwtf8i03mIsr7y0TuV4I3kjYhw+hSAdlGN+yuoNjCS5YJU/j15gUDEJ24zaYeofeKxtL
eHFRt1H0osJwmC32dHSF0ftaUzrJwOrRvQ5SxmrKhDM9Hf8rFXDaKaxPhJS1A3UH6TZDOPjyDnho
++pi9f2iwrsb68I9MZzIh7nIFGcZytI4ZzhWCNonuGaPJuCQd6A9yvRtsjFmNvsyp+/ZlfcRfWcw
D6/jxMR5AaWl36ACWeQOacc2lwHHJAaE07DOdI3S4auiAIPo8I108qfqjiOWhIdbsZ91DAO611xF
dnbfcGaR8FpMrUhl1RIVTVj3oAfKgcFF/moRGkKn8qgg48Ngxcx4+/J3jLLHZlpl2vryHv27bF9f
Ke2W0IRMDvJa1j3uSbWW0NBwncYZF/5Pch0+fSUGVm4+FeeqCzY2rKgJfUnD2F88SlNSsed8BKF0
kI0KXU/778SpL+M7wtt2XeyFTxJ13X7RCe1B6HIxEpq7DicIAIwKqNyLxcZvfbe8exi8421GYbr7
xNRlg0uoUe4rwMVjwaxM0rUtcetp3LkL9z9DWjvaGVJk+w3kQOiq4OKozNTJiMD3KY4ybqJRIOo1
dFBXB0Cvu9SrGAQQeZRmvtGUR2NilUf9GO05JmeU76W1LMiE8ql2YLbqdyVfzQi1e4KZZgWWo8Ji
/viVfKXvnzsdRp2EyYyH4O8P4it5iV3CNfz8hJO2HD5M4OXzwSmy+NQYp80XdqgBLEvsScyKvEeY
bQXbNg/uYR7OxsW6/O3vkh1SwReF1tgCybzCjzyU2s3xiOr4bR8BW2E/E2GHW0Tpb5/Hj20DpEHM
gFj20ZAEQY3U286eqIQ6wLLuC+J1PwNBNybe44tAffgN2jbivFfGd72KEJ5zsOAzQ2AZS6EVPhB+
upgsKx8tMETLnGthzFEjqKXSXtyadQAeQHljMj0PHOkolILlKm3qdxVUNMGtwP6BNhb0+s14I+KN
K/JbcC0cbpQv+Ol37GyvT2WwRoUpWwODGElYXdHIszlOg8RoRz9wiJBwUCdUb3aMO7x5uRTYde/P
cKlDZjf1O/sYea7Yn5tNC5pHHvZXzq5mQ0g8ON3FcbRF9IgS/vCA3eZdPpOt/6wcndBAjB/xBOJs
kNGggY8g10E7DrJWzurKHir+bleoq7bY8mzA4gZCUPrI73BE7ILAMWwni/BR5mpsftXzPrxOlpEW
BLmx/mN6FzKm3MD7Bg4gBNheVDytUXE3kINwuDcWoKykcTYScAywkbHf0v61uCDW6x7+/coQ28aQ
11RtyCbnfGjvb8jYpLpF2MfXvL7H+mKOnLfXIXyR2WdC+z5V+FVRpA2t6b5y0VDceN54yJ7qA9h7
IBFPTWvOYor/hjnwjHEu2w+snj3tvblyudgr9+DwFjb5g8AyzSAgeYjrVyU2qeXb/7FKmdumriWx
q7YgUPSWPXpNIpio/qv6e/Hwpy3Wg6z48CDYeF1fZshtpTX1zT49vyOfGBqkAWVjURKgq2h3XmXD
mrB1T06+S03HPcYsawlSrcdVBMk3CVX2iMHvRl5hAZb5jE+dTsfOLATNvEQ8nc6ptGKQyzYLw/Qv
kkVPXatvqopInbldU5t0pKG9Aj+t/INwFDGz7tiAqeCnUHI9xGU+8i3+e5BVea7XjvST4TqY7SCS
SVMaHVsEp2xtvsys6vJl5oiyEhhL1GRaMhwjzctn32NgaGavlN/B2kWjE7URO8SoAdwhJkTboLDm
gMVBa8H9bnKLW+PowYhs2biOZBJKPCvqnBK080bpmB0Hpb44psyXJaZRFNPgCDV24wHZ+sZRCNAX
d+AutVrvgMnAc6A7TulBFAzjH8D80bhIKNQsqafQY8AMrtl/hgo1gYim5t4YnHYu1IvxjHMa8VML
fbk5MRb41r9CAd1Qj8aapcgxS6FRS4Hsg/NNQ4lJYgUVyvT8xNLayvYiHKcp416xQTVmE3iaOaeb
BD2UoJyFIF68o2dYozstsN1/RA67meaQG0xvjDet+fu6d4iG/7Z7rp4lPXNIjKE9nqG77RgCHlmr
CJcgS/9nJqEgLp4fm5E6hIwCixkyGSX6juJlQiCOc3mTIHslmdn6IKQDj0O93c33Wvmk6jMiIFTZ
/nm04nlVhIBt9rDR5GQhkbtJkyuYc8hiZm51csjyBP6DT+v4ROucWjfR5WoqLhTzgeTXqb/FOB7b
G0owX4CFg6xgYXbWu4jG+aakPx6POCEImliUfooFwteTD0lhMDEDxyQeiFzFTRn5IVyQaiWsOxJ4
WFGktafOlyAx/2wSQlgRiiig8/vQiRKKIuEt65bX0FYEvoEcSmjnAkFJC6srW2phEWMO56LDGBRu
N9TK8JfrWT32TvlPFeCKhpbpm1QvZiqY7YlhdMmv5nHAGl4iLcEFvgMuvg8YVTFUR4unHJbpwdP+
sms761rR2nZ4vc6XHNV1jO4RtES6S/xN0l4PUz7RIudN3I9b5pjKe4k78RqQLdFUeHfmpPjox1BZ
7mu+sVZEmkUq2rVCLscU3pWG1cZFdZNlFSqo7cNKKVcrKdp2yxE+tlcOqFAvLQNB744hmZrGXGn8
dX4NkXmRws9LpjYRdzEuKGk/q61MFkSDkfgf5YYNFu1iZbwxKnGJ45kwRchuUTnk7GuuMsVMuaJ6
hOxLUIe7poIoPh+7qYrjvgiY4bqexW0vVpjKDsUFg/3vN4VTMJQdXeQOAAwS1Wht9L0psmKxtk9b
OkkOHjV0h1OCSVDwKoUuCSbzVu7uCec/+N8eWLh1xZJZmi3ZZwFtAYGCwB5gOgdewUVQVrJEqwFp
ohDadkcrC/M2T7YP+p0pL1OiVhT44jpzmBYhsCT32W4A0Kiz8zT7xhDplPJpdi2Illefm7W9YyLx
1hV0RnTesvLTFA0pyIy57U0m159LI9ut4EHFtuDscUnF9VJTPWmMyKtYfZtRwzkb7NMElbcmj95E
HmIfMHExF6SeoXEEiSVPWq4qTSEnwVHjY3Y/4Fh+HP36GvvehT1NYaudUHXsyeW8M4BRSZaISa9Y
J28xZD+oFdLEi0NF2cATSzsRsQOI+I19zLxRwOqLaSCI/gDVU9ssLJIs+v5MPOBNLxj/EpB5Sk7w
O54roF6ho1A/zwVtWhH1OYmjWvpcyS1sonNnZa/jguCkJ/t7QgpAe8XiRJVlQ9QliXq0th4xK4Bk
clpKnbZDB6hTp7C+f1NSFcsog4xeId92N84T52MzpDq45W2QKIqv03q1ZrPqh5EY2a1OXkOhrhbS
qSxd9cO69EQesB660CF6lVmoEkMJpUprRBJ/gEGtKuaTBSR4xI5fAXLepmisyP0GGwgt0CPOBuKe
/UMGdrs1uSlB0DjocE+nj3QBI2JzhKoxxgZJ8o0loQXlREXHjAeQ03m7CC3fcDAgbcuY0eg7P5CI
q3IVvvAX9gud/ZtRgzyykpxANNfSQGxbbd+ujkQacIIwYDVXWD+BjE8BZ+yyKQ4zAQBcxUahu6lu
rUR2DnD1v9rEbLJOO1SKgq7tsZIpv74ckBi/2PDzNK9xyfC2hwVO50czQQ0DLoaHNZHMWj5hBtbQ
vAlLoBmKVLP+T+LGDQrHZAPydU9S5b9NovIc2c64kSu2dftppN62uV+bdir20eauFZVubOZEdJtx
LQ7WKKnihsEFPyOh6U/iFcmcbt5jzJA+xvj3o275hJUoZ8BtUYrByq7L1dJVbs9MmTEG6GUxgdKi
Ha6s+Ms0IsyPAwkC4ZpqfjNNw/g3M3RB1MhzF1m686+jgL4twgUxhjQCzBtC1JDy5r/fkg5LQVUL
8yTlgKn2dW5JRmeJJyG8+pmMyl2Cf9wMY+jFyIE2oBKA2QBif5LPohh6o6NIzAtn+b7YfFPXFa0d
EaX2ZOzvsA/PhC1r1nek5qvYZL77madAMNVYbc88MZ/0vmeYxXvKrnKxw0rfaU4FXrKyStmEFzZh
bvUbP0LYp1aJJL4/vx2zbktQeSesydoeJIuBW45cCVa6LUgyDZ/I/LTBkfML1lvugr+uVL8JBUOV
2AYSeyplkt/Dgi2Mh371IGZglf14OYP0pNDYvsu2ffgVbw/RkmADxg8PeIw/ZHIgP3/UMtQhmxT8
ENnbJjKj5omTnK7uGW1AaLyymFwt8Roht01wk3c5VEMxiPJjh5B7I2YS68JAczBgW8wkZ00Qh03p
6dJzuk7uFDm92b8TLNpcuSuxdieWBqtd3JaZOzdf2lhPv+NjE6vBENd5cfYVfkpxix4/OaameawA
43qE2NqOVCRQix2rmpMXE392CgnXhpuPOiCF4lxSnxbMVBMsIV8/A/xcgjQsW4KE0hxQ7rdngwkl
j9TGx0rWcbHWP+F/E/Mgo3I7B34jnggtdIdho36fT/YH4BwfkJGZOwugy2+2yXkJzrwlq4FaoNMW
Z/S4kIqjmpHmHtzIlk/pxcjEKMntGXZ3QLPW5oeJi4rSN9zPUHUhR6h54E+FvTgH1q9YfvRiDolS
9zJWanImi5RTHd6JVzCtmIoG9BjgfqalijDS0avRsTiZ8fK48qU5uTon3LMUfL/0bp6Lw1K10rUr
d38yVi022QOIN3txm8OvHQW8uwEZwVdx4B1uGN2dlzjS3c1ntjNSjZ+wS1SB8l9pb+QpvdhivFhV
SjtM2hn+5sMTAKfX5WegYbq1aNTYl3yJXoSEce52cy/mrq2GbNyKqipM0h7Vxq0MSjOgSelCKbQQ
B7xIAJdnTc8v/KIxUoNrL94ed1B2d8XDexO0jWuK8geIFDqbD0VueV1QAUoVwJooSPhZMHmr6NeT
UUjJq0HoKuOkVXk523QUAG+VBxwJXnvVruR4aF2uSuthqK3e2pb/rlKCJAbbZWBd4rgoMs8MeyFt
amFOUSgdVaR9/D5RPRi6Rk/Abo93T/z4ohTXp2Kjf97knV3jvwBjifADhWQKPY3TnHPccwRilTHD
iPDX0DFdtQTnw389oPr9YHiifLGF+yBjDZfZRiXWLNjBFUJi3TQFvBrTjzZjtYxP0iqqjz+cVxe1
gtJP9guRn0mUx/rVRK1apoQRtnFGcjrz6noiICY39qzxP+j0p6ynXO1cvTsbRyTWzmJoRK34EMEn
nsn/+3yFqv+GGH+DWOphLpq1JQZrw0C5fglSCoE/jGtGL1iicMYcv9CZjf18eT4ggN4Vde5vSFUi
e4LN9ntG5Sev6VYR7bJs7SrqPZZOH/cErlv7GWHqf40Nld3ns/O0HC54pRBF82dlKQvmhPFlsirm
NYpowQBii8KNDWl0Xfqgr5viI2WlrobBO85mEYh+6NECWynNyMP9BUNnoDa/yJZqTSf+Njc2Ygqz
v4VwQDe2OsYy4mSCALerzCoycCujQ9AEB/XvnACoKACGm1AAfHMP5Wg9SECLA8tLgMVMm65BLlkd
bYS76P1v3URzoKGoy6JE4ug2Byq6r/uUUf6Lc8bLuIRj5X1rg7nyK+n9jbVwuVMKKodVjYI88CjO
Izdz1p3iQmDDRlXyW75hFZsKnAWI6i4av+qc8WHAaynSCWV5d9htKUxyFcsz0moV6IR23r/QMYTz
sW+jxiPnfwgmPjCSVEulA42rIcXLv93NdHiUVSeBK9xfXqkhGP6kpDXDXWlqOfANMlwLFApLD25g
or/G7UkViXVg2NNYpJww0TvN78My5oiGU9f5YJDyrYqm1cTuUy7wyb4FOD+/vNbl0EuaMskhiEpB
m8xkn+Ixp8eLS6YcBDqM0WZqzghaHlCrwPBBiSA1mQmuMWqm1UrYOtu88NKKhn0QjSSX+9dcl/fW
naVyNhVxeFIlmF9yRlE1/jFp62tMn9SdRCBwEgU9jYshwsmyIeBqvXE20rAPTYHwZPa8AkalM9Q4
+VwXDbsILZYcTaQKdVZRkVVFHC4wmRrqEZ3/8QUytMW7zFgPNkPjNoT6roGvySSARiNz1X9qsmj9
9OlMT1ld7wdvsB+ao/h47F0EblDq2pnIh7ARpqaa5j6QKKZygROsW8DH384jPBxfSsfqHlIWeEiu
lKwrWIucUG/J1wlANQGIwue/AV8vJVoPmpJD/4GFGkt8cyZ+dwdNoqxuLGswecMRLbjl/PyFQA6A
2g4xlO7+UdFs8bl4K2Ha5hdaKAlW9nmG2TNznPieovMuP2LnBg5Qa43SYDRxDOtbHkDC+vm0GqIP
dvLBuCehezYFui2YJd36Tv5DwTsS509QUCOzG7bt4/PNeKb2E7T7hm1vi0oIZY2T25Tsx04uHNXH
/7W3yV4ovjrTETY1Fi7ndJa8NuvDQHGC7nJSzsuXn38Mf6vQ5RloyTsPUlDtUwS22qf0pdqBycYC
8zr9Db0awCIDbxKQqucrQJ5ty4y49FbK1zoS5o1iGH6bsZXT4zGvRjD/oqJA2QQyohOM1GtgpDJ/
MgNggg7HVASqRRu3O7+atgNF25VxpeQPQoKMkKJlsCFGKEGmh9ttOZ8HHkxHq5NkI5ItNvw9uat9
Uz20LCuM7+x7Ie5hgolZX/lv5P1cbwmqzpkgRMbMxKVr1EVXbIzMEr0MY8m57wMJODkEThFtrNLr
YKmQBu8eQehj5lgZtN28jmJ5uXnq7CCBxf4gwJPPXJ3qTrVCTI1d3LpDp3rH6xJaxopL1JjKRB6V
G9RRMeoExs6c22ZFr3RFf92hvwUDN2FJBtXLqo1fRMlwiGOvdnNnxFLFYOkei9POFRlLsIHUuRSa
cdN3joqrxV5+okwjKScjHvSXfWSMUmQ+JPHX8CCqXVxbFG2/uKHNa7wU9C86mxzIuUfgxxsDWW4D
KRJkpgx3NZRfKA9vntD3FDM4gDYlaclTkE9YDynJRtGF5VDxRrTOaEutcC5V9KTHodnqUv98tosy
H/BCjS5GMFYMQ9JV6DgkZKH/5vvDOcUX1KcpQUxrCkl8LvjFH/Q6xm6A455TwhQvjfWXq4mbQ0rq
7bDtXbdnp7tNFiYYSaRziSFMFqcXLpgr5J68yh21DQlVjOaXONhcrxfE+FqfzdMmoRnB0E7N6NtQ
eMnfRQtK5c/l1aVmkFtQI+u9ftYQIrV0jozKt/zW5e4An6VHvL8QagSFmW2f/m0YlS/6EJvhfc3R
cx6dJ02dDcouibb3T03zl9mPp8rZ1bF6E0HeDTZSzlqx5i4f4OgivrKxuuYkRVrBJsUOvosVMqPA
4W7eSZS1KvsBw3EJFSAf13LZAD73YeJLrDjlAqI+rvXANsALS2t37a9YdxulpP0sGAWEAkIhzGJT
Yhq1pJpvnhl0x6AZRJYrxfH8OUIOnvSlVki7UdGFWOlJ/Z9R28bMiys41ZLBVP6a/VDPqFI0S7tU
M7jyTmFWv1u2GqjxMFuSzI636cjBJf8COvEUXli4d0fnb3LF27HeCdeq4NChnU7YDsdo9P+IIO32
dmt3dnKFiETnKY+TKHrazqz2oJN1Shw0du+rKD7HaUi8S+cbB9K/MPROt8pnH2SOgWj/e6ZSKFix
CIqfG5asMnBCv5ygHFn9ypo3NGj2POi6LHo0l37h2k+6AzLfb/xb1R9jyHbQUpvoz//IIwyvQCXY
9eOumVJ0yA3ykA8L9XP3936CN50yz/HuhvOxyAulHRLKJz3f332vhuYDe9D05bY5hOPneMqSzBmh
8dymwZv6Ysc1FSJr8lcH7L7Ueqcc2CBXRTKB9kRRfS5/IXqsaNQ5WlWAPSAx24Qev6Alq++W7kUd
J2b4yzfKSAbJvqmThvdZXvaOQ6ZVBFxHm8XyvW7BqBUO7mDlOjNoG2NVEIwKLpjxVYU6gftnMNQX
KQbxgcoNxTJxUxYDCa7c696SzKraNifxq5yS6ivcDzLlvy4EAxxh2dzRc//ayBRi0zuPsyH9oKmJ
wzPOu35r/xYKDqD2pThmbJY7Fs7YcUFBXXiEhNSw1i+qRSqsgJR1ioA7rJ6YictTqcwnnmFLSmI4
OFe+BCaWHwUEW81zE8SL5mlNnCNNyfqX7cNj+MlQLDrM9vW15f64OmHKZWioQUq00JZdirj0HvWY
6wzBKnYZc1u0LRkkyqDMLooyivRe3EPCriw6bQBieYihKp6KdV2gSr6I4tjMbHZJ3wpCo7t4VXiG
K6LQu8Ubmebo5FCk6oLDSaEYEICGsMhBmve4FAmZZBCdmIMNUnWHPRzcBbvUPgZST8zsVkXNvgk0
UrHYRFqGgvEm94WLrQz16CrHemhnHpBBYAK+YiQkYUqtzV50ub56m2UltymrtYj+N7LPZex9cLIA
UXfX+qR2nSEu8mOobKatjTf1egVrlKjIYeG/NxDcCBI3xLJvI9qqS8yVzd2GgPplub24oeJMafGM
ZaBetvFlNK+Q8jD9RosOV04IcoXWjHuxwE7kJZ4Ylf48Wbq7/+AFzM822aXh+p4rmXC2LbsBDip9
YLxRycZ6gf3Ux+0ITn1tbiFHKAziQrVNdM2Tk833+2OWslw616XsQJrMClTTxgon9RJF1jRlZjxg
4mRJvY/zXc/8Zg2Fva76sxzsakHyrjEgsUxhzlBiS95mVM1fh/eZW4lk6yIT+C0OcS3vJT9XAsJ3
h1bn7QdXRVWh/+q5H7RtXv2ZOBPf303mthkNtImhSPviYYqP8ZVQt43TdHxFm7sAB96+7JbZBhQJ
VxGugbbDKXlch89otUdWNOtIZM4PxCSNIp4i6Bave6flgid6ZUoX9XKUOuJJzCozr/G+/dI3Fdm5
6KzfhsAUnyx5p1GZoHzk41c2ewKDXIWY1H2/3QUibIN47n+BY8tNKGe9efBlsU+zU13ODdkBEmcb
I5mTQLkuVfmLOGl1WTsYXl92qx62yGtevnvjxnvqYl8fipN93c5uGP3SraNBm0dzvjh/EFssP6RM
Nigv6b0wEYq+TeyGKPD98L/hd7AYD77NEqM8D838dVVMypMGiMBIvcsDdvpqaloraCxTZF2+xusQ
/x9Ddk5AMIsB3pMoau3jD87znzGooLDgBUXcTR0wOZp7E/9rN4Qtj/NGkdHQFrRoDDoxTz5vMWx9
mY+vU4YPPJmJS1QeVF4oWwooAvAyo9oaCyF1aHhbE5aAzK9jQEY7Y4wgYQivm1m8wYDZ3KcQX40b
TJ6IIOdRkR1VrdFumkqe2uOgIQxFZB2xLAOw48eXMJe54ngDkOZ1n3SR/TNYEJoZFWa69wwypNSo
U8CAPK9JLfrjiiTsg+6ABV+H8W0d6/gZiePES3axKo8x756jM/FeHjINE2weIoG87bXJF7oycaZ9
e/dxAhdDa6blq3IkNTNQBZGaHVFrHlP1Ip8gLBUhwOWXIKOKAZTxrkXHIF7efSTgorNsxB/lROUq
0+W1elt6+Zk6ru7SKLLU1mxEEXKqyDtA8lHz1ors+/sEmlA+gaFWZTTTBDrQynSTQQR+pvJiJ9E5
6bsWMJMIgJNXb7I+CJGNVuAL0uYDha9SD8A/3cbxFTYanWAaaPmKMlU2saH1iUzuAlhX6MQRGUsq
mocjBc9aau/4Y97smy42BmoyWnoFXBTYH+x+jzpwZI7oEAZ4U2KmVcDsxMZ/eYEsj0uBGMEmaPf3
gzlChERRvumXmndl4uA6tFYaNT/bgQyu/NnKoaH8qseL9pVuZDkj0ailYmNjtf8Pka4R3v/XLExe
avLfO5fubglbgcI2SCTU9ZzSE9CoUqfyFJenE+6+2VtOsu7WKZSutrs/sBhcjvxe2KO5PMdrzlIk
USjU6cZNfNTLTJIwJO/U6faQtytQdI+VtVekt1BzxjkMz4qwHqyPGSG9SvynmVSRUSfBHoMVkBMj
qPuAy97hC9MT0RqMvukJCG5eNYDxTTJxgmGeQmg5E3gCrchCqOfjWf5CMi6LWkhIQ+uKmyZEBUh/
0qcEbY4rKzFbXnpakOXbwwqbnC3wbz+wCOX3akmMHfWlmj+sH8uQURIMIvkPFx0xKoQuxjGb6Dsx
wGS3pEQEQdwM0W4YVLQSfphF1aRyTzjZ4Vm0RiNZtd+yvDF9h6BUjIinhmYT/5V/jIRqaknftxIc
sY41kuUmMIEGXDRIV54ZNdLH3lRUPnkO7E6Y6dbQgiSkmzlisKueMN0XDEpgQHYSb2r1XrCvHsiQ
jg/lCeawLKzfnaJWU5hfNwA7pliUaYs3jodDhHcx/f0d31MjQS3qnWi104NIIPjBWYsG+6zVxMzV
YGpPP/cuGrm7yQYMGLOp/jINzXca4XkAi4v/Bhi311oyjzCR5i4iALHNL/ZPNQm5HdqkVxFqP9S2
xay70YPrCUWrvVzqTWx1D9iM4qFTGRpTftKx9jYEPIeT1AOHDJTP4PKxFdb2PT5h9CyF3HnDLAKP
yqfcDANZS0o5wtSfqoGQAm98pdLYzo5DIEs5XOL2Hf4qLVuky+/s0JmdP9uQzfdIGs+wMDVndjwU
LCtWAS9v4I+TI1++OIf+8WarxB2MnYhvaTwJhjuzJFtuNc2fF+Pf5AVZHwmy7C3dWuF6vRdokOYc
DVsizs4SH2rK8IuyZHllyNiDbaD8GOOvnSKLStO6UZNEXZlpqZMi5xqiO17ClruubkZP0I4GtzcQ
20wE+4RqkJJ7Hob+cTEzivzQOxrGCf5Vqd5cJ+2OAyZQT6Kjm24eJFUgrkxoOSgZeaYGUZIQAgr1
ko4j6f2o1pc2EDGzRj2HbdySXDNbB1lUnYiEPImswkGIlcH/Kz9FgHZgH6A0i/CwNwFOBdes/f5c
yumYejxtNrpuMkSh0g58hzayXZIi8PZ+NYDMEFpIyYH81VDpoaPtVRUAqqrQRXkjN0Q6s+hXu8CL
jxtrj6MJyWctdV3yYHj0exdMFlnvBnunlEb/cE2yZCJDNm/rJwzr54Q3JzZ3yP3kmk4u8sXrLeyc
RhvUX5I+or+Je0zZ//qiX+Rfla/EJZg+s8+QQY12Z8FN1/14zcbnbYdxCRXiW1iEac7QtL409OAr
0wQvwEbwQZu+Vd7WSq8lLnZxK2jC+BL0szSdKQELfS6gDjmm0YPGJlD3dHwTvFGVsfH10dNY2W69
zG4cRvwkO/YnlRVb3dGo+S7rs09f2K0kxv3FMupy91Eb44XEwduL92KrXZB3aYNSZNmVbf2VqFq+
i3inPenhIdGoQ99CeH5JVPoxEocvkI3jCh6KjaeiZ7X4BeZiILWwyn0P6v4VMjpOMoQIKcSYHl5h
8p5owH7FAXLKZXYNNIf78Wv7DRXk31vuF9jwXW9qHRUQb2kVFxSeSIqfrUzEN3stL4FkXyeqDDl1
jhl3C/X0+uo07xcnAFeAn+ayAHj2JzAsRk6XANVSjPNuywZIHAgnTjyQY6bK9va0smN5S74Kt2Cs
ruv3Pn4FF2CnwSSbTskdWGk3wOk1tOnxfeCPXfyx5GzgqyrhUeRWxU/kAbzkQcK1fEnRqSqLRBc8
NmgoFcdZ5Ez4J8tDCA6d2nRlyW692BQ8Fi8a8NmDUxx0jsC+rT3nsL5qB3a7aVZwp/wsqznqI3HT
UalGKtngyf2uVePHmvzQTivNRcoBvg1Z/l2HStuj26qO30WaxZ5x7UEyjBLAzu9yBIl3fEBJylh1
2QpvehMUsKS3WUgXUWLcLFKfxNGbzlUiKGxjgrOieEEhVJvkSsxwCWoeFtctoXPzIaFhhjjBBqGo
/k2D0YOPS8Fp/CRYiuV1v54FQQ8a+dE67AfVSxa7xo7dQQJQRPrI/4wI+EE96Emrh6PORk0cM8JT
AUSFBUSRuVkZYwfyTKH0IhViKBZDBXbG4cv+CmWKHoqvMSLyUGEar44SOA4SNREIVeowo2wio8cL
JC9NTjTtLhkSVPDgFh4L4pXVzuQCf9dlNUgpXPjxIkF0iyzIVApEj1wJkY83YlRl4RiEBt+Piwrx
8CTBVB7BgejaDkx8dT/qDu8pkHaRrU/sWVoo3e7LiqeicXmFViWdAuecoLv5C9M8aVNtNTCzuXwn
zQa5Hu/dhLgApYtIBPSvWOZNS4+hBh3UgYk9QoHwuFQQ9wlvaae+xPGASYC9hE4oTs+ztBlcUtzj
TM28dbNRN6AcCAKmI6pjkRqtN6Yr2L3pkExDctZ/8Az1e6HDejZCyuX0pFzA8CkcSbGOeD/CmXrq
QxOZX2mOg/tlrL077uvTZOQlWU4Z5qVog2EfKcomOakgyGiZVhT2haocRoP9GNntxyL1B09CdlcE
/gfjr0yYAOLvfSzvp/YdXXpdJePR16rjUX6eEcboqAEioaDKEE4/0Rq0XqMDtphwQVmEKMR4E0+g
hHTOn0s47PxdVwNbXeRNKn0UkXnbGz6+utsRfK2scQHAq4ZP5XOdiqTj9eGAKJ8tHJ+GKXtqQAZh
9GVC2FY+ILomOuTzR4N3EQPt0XO+WmxPD42cibTrpTLfm7KljVfDnhbkXEezV/bmiOdB5uAEUJ+M
cf103oXeOJkn1s9yc+On9I5Z9Gn46JoQolQyiLCYmjW6wgK4jz7JViI+HayjDQ+gjtEgQxmYufSk
jqGEM1EnmMYifwOAxL4wZ62OXwCjORkIOhCjmn1z2NdwOaygMuCSe4vWVO8OiKOuU3b0Q+bGxaNj
5b6+PutKOKwV64DTP0nmsfsJq0kidm8WhRX2Ohw7L4K2K+6Mya0KiW/SM16R6twp9tWwVqp3LGkf
YqiA3HHfZWEdR2qrZydCK+zX1NUjnORAIXzHTRcv39Dni05gUEZoTl4xnFjPIXwaBgzaySE74/Pg
WE+KasqjNkV0oBXQQOb1KztfPT5Gu3+Uqu2EZqKW76s+o53ydcZqU5K/fdC4oaVqs6bXoH1dPBIP
AFPvOMmW5Ogi49AWJGxEa7d1QhV4nAhPC+egOCuPb9F8k3SiugQ7P1Lq5RzyO64eVhYFNwdvua5U
K34nfJNFINLdLuIqxxKZ+IG5DdAkjh4k7I21sgusN8xH2F/ORbyW9L2LGD7fLxD/YqYA8X7an0V8
aG5T1+ZlGNJdzlC9AYWsc1iGNkoCeqJLvVvccdAHsRKWSHizynmv8Yt2q/TABAGSCySajxkrV/mp
T5k+5p9xUAWoUjdVqGED75heTk9XZ3QYwYh9XwLdZ8/m7in/oQjsf8Lr9GdjJt1Qi7SxTKKQa7gR
H9lnDVM8NMHg+2bL+/zo7wXtmNpT6gZ50tYxYMGqpRvnlx0WITqXrXcjqmdxQ49CEPVA5r1NaeQ2
DWiSF/OAwsBYhsf4XvAuNXRldP3GLnjZw3PuVp6boLKc12k8PNqtIqJ/BzDvtc42ImxEY1OXQfw2
MyzxiGSLUpMX9pi+wXyUtjRYFVBQ6wufLnHUDabtl9GWWWJmjWIFfPmdHwnS1xAfKJPcf1dNKHXf
eDUjUd6TkElPWA+CuT0wOWspvLSD01jxEXU520ygfBLm2R4OrMPRPFDGiDSOoroWQz8kDf1kAPnY
xUwiCXn+OzU9sys6vpzf4uvEcQXlJ/BXt+3MKxS/LMeO2YEbzt8I4oPxatUz35LCfZE28qPkHGKa
jx0pcNu2PYqqyQHA8hJlx6hno/7Sm58tsFcTefIrJQJpGCurIsFoLMM05KXFLW+sXzLo8Czkfc4C
5wi3Tw52KheThxHiWR8Z18ptXGQVmeqgXTnIieDMVbWM0jI71b3E8AEqdpa+HCaWU1pgW7963beM
xQbDVSkVXld+ulX5ORrDh2gAsjbaNepVcILOf9E9aNm15vxTyEAF+I+RrwELy15ItyK88Jj803Q+
jOWXQOO0MScgxwrLPgIPjTH1EQQxNEEgWmd+3cT/i7Q25w7sTUsaWHS9WjtRHMgaH4yqXiXmXMhj
ovORlsMXZzMgvdpCszrRw+avO/fxl6q5Chs5RWzOJE6zi2BG9BkfPE247zyjvv/jNn0gn8NTdqXi
W8KJ+7C/ujxFuCoYlyedGEOHfumXPImlqxbC6BkrGARPD6efsdi1v82Xy9XvtNNEVL4aBnX6cTab
NBK1kqxU8DEyWbMTsX54MJg7XBm4+q61JbX9xem5iF3DPGYcyx9gc3GnDI4IetC3A45HG5LveIk8
fSckzuy0/PeD/oeEvLTHDck/PyjQ4jBCWXtKk4apWGM5ffEqImFsKb53TMT/lKlv1nvAEdnbCzoM
cSDXNcSWn3rMx8JC5L7u8MIxbbK9xvlFqvMqaIlMko00Bv7zIEJ5wfQ4BmpvX0kfQIcOAu+o+/4W
tRUCUFWFXVDN0tCVVq4SiUrQfyJrNIF2Yue6UQiFa7lncA5xd8yVpo+mFLIRj829ZCQPSatKJSQF
iZt1B2V38CsBGWNBl06fTdU+EfqgFrsLjIb6SJHKjfoq+ihBK9DAK12ooeqEMopIalNOxPdrusD8
Ri5NSM+xOnPe0tkr5YrNdewiKs6WQ8NZkEuloJWw3q94C4ESkgqrXJ6IEV2LwIqmXO566Wh6bkk7
Gs3dmh/VSWH8h2Q1M8hSMyo/9zLky68VJgcZRQ4oMcZK2S5Ii3zG9k0VonhCUWhGRz+oVHHGvTGH
E7dAFs3ejsMVFggI3FeiIuiJWRzz7/U14rEbAwXKzH23gQt8HsT8nKmRMaiQFZy1Gv/0Wfxjpxmr
55Qixanx9XSS9x8C8lRUu1hTeYPUquFjPP1hz612r1RF3SPohj2GZ6utCMEe6yiKZq5eIZQzfqxi
tcB9q251xzXOr/64REXlV7jRfbxDxD4dRgWyoVqfVw+HVKGdr/8jLAIUruBXzAgcrKHgSrkmSYr5
Vfpmp4EUEAxGuhpwnNvqlLzZfuZoTNSFh6nz0Ki40t9s8M1/i/IhT9hh/gFFRcumeKhgQOMhQog3
hJmSD94D5msf/JThDnP3oYfXVw9RpGe07Ciu/ZTF9RG7w1qbFfWpjcero83LDu7HJK5ekBjArA/Y
UjOu5mgm7vpXIcKqHwWNJ2jtXAjRutIGq/88J0rLfvd4lOLzYtqS/P5/GnuqITeVHCj5xzzCkXnc
IhFfkPsnOpumANSUsLv9DyuhV+klqs32RdxW9Ru7A/pNCud30hzCde6lnAew8CPoQnYnXkSazfpn
Do7No8ZvIma3peRecJPkRqCeWHKtsMEDCf3CG1lC6YHA4kCntJpDAWCVBI4yoLn+SWlUmsJ4Jx/L
GQWANuFYY6WArqyus2me97yS0rYCVWp/MbXkA6LOsa1gRyZOGcHh17ZNeU4ASUlWlpHITT2I76EX
cWDli1mf1ttkTFSwCz/sSlGqZjCtoiytvteOU1c1WWVy1v/wvVwFdv6l9B87lUGd4c0DFmnTzAH4
Vg3ywjEDYHXk/EC1VEZxpY61rQ995VnNpvOEQKKxjyFTV78X1gR79Nlkgz1WoKXaifClgGhDc0C0
k5+RY7jxNTkrfMPzfU9WQIPFzbZLs2doRISPmXBy6QenGEwhBdt/yEYx2945z6ZO/AN4H4jw3vBY
mLKvn6rI2no/rqVAY1OfOxg77X/TMT85JrRikmh7a2zOXY+P8bmZ+C13P5IKP3MS/dQILJCYPa7K
3NOwJfGCuPSNvKNDqhbgQsdu6+vuA8zpRmPToc539Gulcj3gZdV2aVco8he6wkAohVweYCzZYmnT
l6HJ5PCeqeDJWQJzoPYmaQWbVSxCKxscxEYko1jTO4l+EZOM7u9JnFxwqr3DUK6/Y5z18VZ7riuf
QHyxbQVAW/8ZxxI7r1h2j66ET1uXGVcao7q8cth8T7QfnAPCJdM3G2Ow5Xw70xE+7P1kgBQVKhqp
cCxW6w89ZZ8RY3/fso1f/4OJiypfgCqDrH0yQ9FnRwJqSzacEhX6EFmIy9LxgM/5rrNoslBN5aNW
sLOZ53TiGonTqvzotlMc4MLzgfN50SlrFMqrXy8VMrKtgLSfYREg+i09gP5m4qXn6YwWQ5mhhmgd
BPuweOnWigU8TbqUoDpeMH9mSnhnH5es68dJYWn+f2I8ECzLw0IydJkmgrhPrntr0Ea7Es02vxSs
wDVNmKAZDjr4mGsYM4WjNEXHIAs6z22BtSB4fo/o3cU4BnZ4JXN4ew172J6Qk9e89tat7V8h8Zzp
SLeKLvgaIwKI8ZwAo4Yhge7o0ZHwwhp6mUhBbv11eJZYMa9yCOT+0vmsLJ3AJHL+BH4WARCO1zrU
FV476MZ2tVSKWdpFJUBPuDABJV8Q6rPVNgip23hkV+WirrdXfmV5
`protect end_protected

