

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
kNSODHF2BA8phv8L5aZNyOOK56HCcQ5lgKBxF8hcTzwkWRF6WnOKZaH0cAk+oZsvi02J9SlLLySq
oKFSyBG2Dw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
df+BuhfNWqGLyuHwX48C4kdWet0FAm6osy35ZO6nvLm9LeYvgiC7d+QWQpEp/leK8jaqvimQleVB
qNUNsNTBZzVm+VZnT/+N9fzr+Kn5brl7DACKZQsJ/J0EK++GrIymGQB1+7LWFg6RjvqxHctXSERU
pIxXjKUtzcqAwrR0kd8=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
j4klfuw/RrSoDKuTiN/Si4GPF3r+1zWV61wAeT879HAyso4ajbQGVJETjBzL4XBayVtdsViewbVc
n3EWjppKn7DU95ziVUsafFQrG5PCVJ8TPZUJisZwRf1u8N8ojLSjd7Gi7vpDvGySyTXx9aoOQ69U
XzJmTqPAeaivz/FLFyjHWzMuc078i+06EYa3j0uxrNsDH6/IL5syM3QcJV3812LlPGSBhRN9Wynk
J5AcITSvkzy/dqcKICGyxp5ubBr16BEoG7l6F/VEXvTJm/kJnHW75YZ8OAQ3I6icKjHkLZysnDlK
KEU2K5X/pkwYnpID2ogdwsEuEQr/xxo42oEmKw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
AG9C2Ti5ZMi5neBsWpJ1qwXbrUaWpaRO8Qn1fL70JVZk4SiqmPlFkL5Hz8GrFfE4eBlngUFZoung
TTZ2IeyMWjxhdHHDVda6+BqJtPiX+FBQnaCzRd4VBLDnB8KUn52eheU5F9XtqqkHq+oJV3U19TRZ
Rq+NhUtknFhYrHlVXfM=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
TuUXpu2xk+duDJnZONHfYiEzeCuzIA9y6Ut5Y0LAE72Cfiq+aIEHs4lmSaypPxj5+E8SKfd42Iqd
iKQPBy7GWczcAr4hdHMLEortigKfhxQvyiAB00CsQyuj949i0l26Eh+7iirhYh907kSXNLc4JeDy
uXkHZzsX9mKBsIZLMO2TtO0R4ECsHQbqo/hSpi0B8kY4ucdqtZfLpEsAJ7G3XH1L+CD4o7on7UAz
BPPpoVV+VIZR6heT9EgSZTHhg3uYl38G0Ezv8g8s1cbXnSuowx0B9mx89vkctBzRxFOLnzsFdBr8
DIKQCrHZfdOhrNHz4ZkgOrKjCDpwEkMA4ATVfA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 26464)
`protect data_block
aA92h/dMfiiPKloj6tjH1dY72+/1DtULyEX0PsM4rDUA2CzAOchNwtXBL3++qjEIy6YGUHsgJ3QF
xFQzN3kJ/HoWh7EYmvvpkx/ANvME9V7CewzTMYUa2X6XpeW79ZdLf1LFKTEDRnMNeAb3+L+rUDVK
Rdwyq29QhWsgW/xUksCrjhuGwfv1LfKCHNqAqnzo0hCQ9BtODnyMTOEj1Rujj26pP8cS5MXpd8kW
R4CYdelX9kOirWzPAEnba0EzuiD43H+7nT+3GyHfwHsRbchsROyCKf98ux9xnfDWOsff1wZRCsRn
OUaWfuG2x7+VwOA8fiPyVydd5ht82TKZHNcARdtJZ7RnM9cmgHO1ec6CCaLIfvCaC5PyDJkBTELz
K7WBd0+Sb7Pz5uoOlE5rhey3V31iLebBkF96ws19ww8ondB9IkPFHzG6vugqvOjHs8x5NRSEYR7Y
zKsw7d7zCeHB4NB4SsUBKUno0GOBdlAVhQVnOeDg+xKPEEaLjCWsMcK5U9kgjZKdn1s5x0Io8t7B
4YBN7op+2A2nteW+A9bj3oteWVgBHrCfdm7Zd4mTHsacps/xzEI+2RCL3x9y38UkdRk2+O1d6xrF
npnBI1ML8KZmrBjYKfcQ4ZSrqndy7/ZmhDYa4LcsZkEwCkgaMkN6H5aG3QF8HCDPyqlw9mmFP82a
FvU9BPuveKJnqXswQQ6FjCvpTVo4+jHfg8OBpApF8hc++IaBpB4xwJF3GziKZ4M3j2tq0KWu/Kbw
ERrWACIEAPD2IULNZev/6CDCnHNnha/IhdA09XZ3FJbJZCC/jAs0ATuiZb76nv3cgxPx4+5nlA5P
CW6HMPHi5LCtRd8BsOAagM/Wn34D0d86Q50LfpqguUE5j+AVv/9VzmO/0J87FHaSh0WGjCaH+UQB
TDlTDVK2k9dt4LH8BYiEymJEXcZck22AZKwHz6tKOxQXx+erDh+U/2Aex5xcNKW/4c47M9PpSpuY
qDtcp3+WhDhC6e+KI7EUBJB+Fp47KYuERw30K/V7rQvmE/+DqK2l0RSc2Q0W2Z1GVmgb+DNyUTF7
T8C7AXSlaRFE57SWWc/zHY+wzdqPwiFirvEns/ygBTBViNJRXTKKZBg0RTh32H3RTj8j1sIWA1Yx
DKk+H4uHXmfr8AURgcVem2RXdzn1xtpcYihh0cYSyTLthIlQkn9bQzV1dH6wWnCdcM7pQBEEvzh1
C0Elsvhmc4kPZdoz9a+6m6k9/GCbgY7fMnAClhHFqVBU/8Zy0aU6m9zGfIvvBdMB8EfyN28gC91e
20PThS14ygGTVt1IERp8LzqplBsYhgfFch3qzRanpQduUM95IEanBWl2OzRPo/sPhNQ2Wa4JEups
N1Fm1E+ARU8ZD3zlLSbRr7zNhxJSKVybErn8c4oQ4avgt/VqK6zv7FaXtsuC9Lr5qXAeggoG1dKF
3PUu4E5+efY7YPhUSgQgfKtK6+BHIW25uiAlJSEJ1U7ElUBVhrUHK1ZxF3o8UOBps+nPsBJzOjkA
89pcGR31HsTm9K8o1nsw67q2KrU5CjoKVXL0QYPUhvKhhyvPOb3v19KKUMrz9AoJgDjZKSiPSiS9
r+PL/dzKIbGv4U8Qan2Q5w1kzV6nL6q/trTC/Y22ix3sGX2MuZcg9oH1TTWKJH1EpDeUH8FXnw/F
FtTBVBOVkxfo6ffhhxzhNIKIuUp8VGKJ9i3IoJwxw3roMAFusSxMFnUSV35VzMjGcaO2uORZecRy
TNmHkBrHlBNaAW6sfuVY0qpdzObymlWQVeVNioMxjSO4UDhysxgc2PJrydE9GX1oFM0iMtfhOUcI
mjRrp/44OB2urIaw5hJNQvVGKBWuU8YkruUnSJ9dIlCIJTX1JqPMkHQxnNDppEbYIPirxGJLVsgh
G1RGnphxDE0ikiENBHBfhaebUFAdZP+W7Hm/DDnfJ+NAwAX0+Hp/IOd+AZW0hl4tjhq3JBbN6clw
8Kj4C6beV96tSzgyUhi+cDirR9yzbL/QhdDf6WK9HKyDJpqJxcrg3yqx1crjzM13iG+WeDpvKhB6
rIj0e2SsG1LLDPHfqt5Ps7kQK/3Sjabxp/c2Ua6/hFLhwvNFpZhAdAGbggE61vsQ036sZhwmgH1J
xbLPeXJsgGAKXx1t9UK+7I58oTiFSnBsJpJC081nNuhur4ROi9wu302Rjbly9vkDSMtAi+ABdF2/
LWf5CmCtTbBFA04Rs+2ptmQS4nU59NZBVMUX+CrITifH43e4Gw04Lycn8qWFuurCd5PkZvgNGiCZ
YZjqNCKK6iyD4oriGJJ0il752aBGmah6oRJ1j0boGzPMxd317/AT2NHlALQnzRMd4/2qvyapwISc
t2bcjpYn9vXoiVt68Sn0+gEg0ige2PlLUaikWRFowJ2U8IV9T22YWxoICWCsCKLOlBzKxq34GFgm
BGlMfphuQarIZYVTcDHmhlTnnFkaxHyz/uG2Uwl1gtjN6fq9qH2Q+EL08ycjBsS6skM5uKrlTgEl
VfazNnZVjL67Fiw8fci9sB7VwnyBj9DF6fVtljMUJp5HMtI3uotF+fOChNZkqVG1o8prT3mX23g1
oaRRSxF5UQkK5iDykIDMi935QMFQWEN7Sps31MlqCnv7MHVtHc2yWvQV9nwNUkse6Gj70ENPy0gd
r4B1JxFMdh+vCKdf3uWhbQZhNAFiLuJqSUSVX+0qdESF4fH1TffvI62SDJajVaeYpQ4AI7qYLxEj
r+eAKz23CjS9D2bByZ/s8h0tud6GIcmO8D+2Nwsl0tiTgNvjOYHO2b2OvNKcKyWVQ5axFXdRx24P
uryAWVb7FMviKC3sqChRyXL9qNSu7vVq9XS/5jhyUpX/xWf+QwKz2qt08Hc5H0tfQiq6jvX9zxpZ
HQh0XdfgN5qvOoWyEVpSin4p335noVf1UXhB0WYq6pGUcR+sNdzpIvnz0bx5ngZxnmx9bZ5cPuXp
aB4InLPIB/BdgFzRKW6LpcTE6Jxx76m56CuslGvHmwou0Q8a3bm7Tt3CJf+xfBCkFW75HBwCu/yy
0tiYGpkw3+EC+haUvb9KmvHsSyEu/fNso+WzDHSGN+m7a4e3tLI5nPMOubBJtrjsrW1PhBHD+waA
3iqliEmU9fcrcfKQvKpPSHm1tBV0dpUY4dxxuf1gdfjGp81LQa5dXVPh+OpifaY+Acc4NI1+0sf1
6penLKbPjPE/aeaBPCisrCnaJju37gHiASlgrLlidyag0yt2B5gc3fC40s/RQWZets/jEXSq1WQe
BT7wK7OQvaNXrRQVERpnx81q+A4t0VMZ3MFK3EIc3Ce+j88EXwQSgHLT1YPRzf0zQacP5eSryYch
eL2gfmzgPdoQLdJa4jTOfBTtIDplSlfHSDfmhuhNhZqP015gdR9igPOnmdpAlecKWCoVAvU7DgtY
9l0dVXTCO2EN/RokbpiQM52m7/r9Df2bACQqS+4RoUnk2A9I665S+u+CphfsjzeZ53KF2O+5nTVb
LWwSrRXwnWblafW0DSiIVBv6FDmoHyDnJzs99XdJ22iogGk57QTta0xMipp+tOAUNyrzwqvkqqXW
YUzUlYN6mCFFs/z47xyMduftYs+Tt8C/e5Ts+82lMZpgf4fna1xDujEb1ka+7fvf2wAYC+l8Ia0g
8NauLBMcIew+dvYa3dAPN5VfbKqXtPT8w1vRUgDauDEoL4zmuynhikXRzeNuvBlNDDhO7IpSci3S
CdbAjW72C9E8sG60drvT5ekw/DxoLofMh27ILMJDVsWKVGNvv1tP7rFvpscEE+pOnqIY8J3FQXpo
cHCbX7rFDqyCjf/xr+jPFVPycTWfttrvn80PmvOZJtVpRyoC1HsCT0JuDPIGWevUS7UylwYeJ8Cs
KbhagJxMuCqVH4U/7NXYl3ZdtIuC8NUMXWxrKI9dQmW4hjQx3OHUgUulUvB+T02WQPM93i4N3ihX
uTK+j0J8Z1M/NADEqdcQfuRA6pSJtvFvpYtKudA0EVtrRVQ0t4V7aDbFD8R/rll2HqVu8YyrcdJK
UzcKeNMWOglUU8kx//4wAZuzYU0nQTy4wT2hpVjr00fL+Fw9wlCT9pmY+Fns3neyPSrQKvOav+pw
aMEePzCK/nTevA9mE2qmZMIQnmhxArV4cW+9K4jO8XWq7G2vfNonZj0anZkIfPl3fTgvNHCwCL4X
1MAfcn4Cznc7UGLLLFNR1ZTejcCVqH1jEvOnZPx0lrFSQyBMNAHftf6hx8k9VlkUtURGrTNmPXvS
J9vjeKlEtH7lrQ2H+JbijHGftsQTjdrP6HQHAH91bzifgN5D6h3aLIQ9GU9bZJ2K4JKTJRL84lPJ
1l2s/BOKo2V8vb9jNawspHei1oNRn7Vc4O8jCSFdlPXMtfqLyC5wdQeHjLqQq6prIbk+mxifqHs3
5+bCuQ9nk/kckXDsYHU9bnIX6K9RHodYE/fMCt2EBexdXOdRdX9Z6q+fuKRORZiuAHnZZG5qx+RI
Fsz6IvAeHyEhWSticsmFjTCrJdfhutv/gb3XdY5A4sBRRvuSmO3jmMglE9DC6fX/He4In9lBp1Rm
tFHgClxGm2DD70fMHsv+dwukrzqjHSGo70aqZO/LyPFkgBMyXymCemLMqRfGN57hQrrOtXZfdbeq
QX/+NL/wGSwaRBF7pqPnv291D3HrQuQuIu8Sp3FIlUhsL6TldZgUvDH4Xhj5vRtPxeF2B27T72yL
5y7OnZzaY5c7O2i3mgI6+Wphs9j1NQR3hXJfioCzNFa9jcS5U5vjoyAlOJm8coQLTAYzA9PS9+PD
fqZvdhfIo/YyR5NVlfVEDbVtP6QVbA8jYLsC7ZGGVeOzGkqQM1t3XYQ6rbcNbTf6i98A8yvdNSxm
8EB8DdVpp0I9m09rHPk2R8xccyVYcnhAxqRboawanGQwJjYvZmXhAkhabtY9njT3vlk8x5b1QkZH
RsEWwkADzONP830v+o0aa8BRlI1byjNJbIfEQLAcuVYFqoEKsn9h7w8MdUCsQIb4pVQVRvcfACDo
LqlFV29p05eYty+zHWC9UXdOaM9fc/U5oHNPiRP+aW34Y/WOFaj9CNySbfxxr57F0EA5eqzOaeum
hbfKwfiluPPfYsjujET3du2d5ZHe+/RxsNM5oBwFi8+50+WFiQT6224AzsAFDajrIFeBYlunTJzh
88etc1X1whTjefKtCzvbEXy764fFZIiWsVzyEF8YOz9CWrEt25pcm4+rrXB60H47dOpTzZfAYuoc
FHUtwWlAJ8A2Go/6sUZUmb+c/nxJFOq36oy+N3Dbfp+ppZIcgnrm2qCWheRb7/LFEuLfOxpMCMkn
1WMv1IwLi/lyC/TzcXFtXmzTcJWEk/kVtLuXXPyFKXVqFfxGpUueSesnhoYBzc1kYNE2pXLmVndQ
MumCe6StNXY1+xCmQG9fh8cOmugrp9SmE8CessgpXgy5/vir07pQsqDnEajTIVWih36MOklM0gim
1AEj04NWlXSm7xbcz34bOGavPnpzg/CMq87MPsgdLK0nizTFCd5i/dDKVlnasg1ANgOZk46O5e5e
pU41LXGoSP8/H+Q18cB1mC7oDsmaNCvlOEoPLD+7Anmq2MylZ08DI0FCb7g3vYMu06NZUhmf0tEe
Kl6ED+h/TlhyMZ+8VUQrbv13R1LBhRxLqijFefR8Kz106OkS5Jn9gwlZfYDwxeFMl+k3njMeT4tu
lgyTVJuMphw5bk5zR1Km6dG2rXsAXY72e1C4ZBenx6C4Fm0wLaBVDS/NgiWcs4EiHh/3qc0h+tDJ
RpRKKXzzrt1IgHUcSNf3/m7ipB9+H/YsOaw2JdxhS91SkyOAs6mxGgqRTrvkDvDxLZrVRLetVGLO
U5GagerjrvK+AH6wMdBeZ4f1W7kf6xeTOBhiaU+MNqV3xfqLMMzJ+dgM+0IwZzksz8gzJth/C05S
Tu0FJlldTSpOnIeDpgO3GTR0FKxeB0rtcaRlgOpeseNHwm5DH7KarFGT8QTx5pymkXR9ugrRKWE4
jRuoiHzqUzkSwoksLUSjmeYZshaCS4VMlCzyn6SADMx5oGfVPUf5/ZrgB+wxyt4wdRj0YnTMtEzS
LGlAUb8ngW2/5RWIsQhRY8BU5KwMLQoedQ+5Ot1EMQmbEtxCGGLnfQbksXCHyYNC9OHPYpV7XyLR
kB42ViuEwOpqrre9jLsMVXWrc4FgSeNXaN+iklaEgjYJeM545PqjS7ivysWDO8uP+DC76pSUsfMo
kZ35naIjEDQqo3+Bb7AGgT2htlMlcwTO7Fp6nMzdxNDcVise7f1Txj2DQ0QjMxj5JV4CQj37RIki
q9u2mP/TBiav0b8pkI6KmhvsTc/97IVJJrGpReUgIe/CVhza80D8CQ7IUR4xAn5+zVSbF4M/hmDv
U5i781pbreUOraJ9I8lI5xO78Xb2Kb/xsUt3Vqz0NmScZH3ngBw0QmWilBs1BEG+6K7BZkWhuHzd
dsAJHmKMyQvj4brMl9AewOjNHHoNG31KLygivP0lwM2vGJpQffcV0fs7WOaPpcfgh2mlid4dWX3k
faPtsuqYR5JD8J97GPD6zCIco2r+lI6Jp99sdFTTSuidKxnBFHmg5KY/VnGBnpiBE8eSnf9FXMHV
AM3CodeMmCNblaHRsWei/Z1un4FYfww32FjozD2u3o+TO3iVrohN9Hr91FQTuL9LqdB2uV64Gm8M
rYUrBL/x3hbdg+3a8xH7vGC81L2esn79/WgsKnkGr6gAUYYHQ2hoVgudB9xFUYJC/LK72gRZsMJn
zefIkuXozzVyVrAWL0JQ3tpSYgYp6f7cXg8YzuOKhe9ykoUFRC/vfRjF+wwcpoqI4t65n+4k9hy9
JH9SJdZwIlO4lqR578qz6b3aweJaZhFi+0Q2ArQhnJFSshtCx+KaGX6duZnoiIxfYcSTb0TcAaAC
G7HIbKvQ9mAjWYWtH3b+SXkuCzRFVLpMz5wwJNApVIB7dOUtgoeSvzc3/rtXnoYImwjgafxbnman
/4nWPoLj2VKNRHdlBNnr/iEDNN0W2Z2kuGVZqYz1XIa+raBhBz62Fpiwc+U/pJUoy86RmCUnvH1/
QpxcNKmoEMYUTCh53OQHH3175SNGFzRtslGl9saG/aJlMyOkddKIvV1udyNW4A2aL7Lyt0xl2mUL
+yTpNPY9JyIClbZv/hg2oLw3zSAF37l8KnctDKhQWYzQudCadf3f6fRksCgpcsJkuJODeCZBhQwE
4uGTHaI7zogqJ29FTFqrWACByVDajMiMnlVv2eMSb/Ceq4y6fDGwEO2/QOWmeOTooytd5f9J6Xpt
esO3B3ETRaHHwSeC2hQj/dXNF/Pp4tWiyRW9rm+GnZEf7S184Zn9rJ0QWkOgOVdMJKYqeQBVCzBL
6lPfDHqd7WZJ1vc+2goWZGq5rHtOJRxFEFOeCBrQP+sLF1JofRg5jAoVCG8ARqZftm44ctho99w6
xqCD4y6wST0PeVbH72J8gepkVEtb7gpymYMKRS/L/XLDPcgUOtkzp7wjU/WnfUOx1Bgb2s/okFGX
iPyxmr5MWc61vk9hxxJNaKXgJItPJAdH+9+QawiSgHbkknQ2INdaps+2qXmWvv1QuG96KMmCqDKf
1DgcPhq6vB9ucXOHi5h7O5q8iLcYD/vvrkiIBJZ2jM0d+aoKdEmr55Nqjdhzn3HqMd8n0dEeqeSo
nKdK6kzLyKBxg+JKynldkkdOgNPoPhLVeIQ6zpCqBphtPikPvuVlpWqRQ7jm4pDn/uJqrKVp8qjA
1d7kvmZ9wKxW+3hh0+ArluQQMbhglZC/bNk5hCS4LfMPhle4bijcJtbT/9gw4ptbtizZKcD1k6cM
y5C3aTkZrVCRkMfxps77xU5Wh+Ov2YegqsE6zEh9wf0yOtPB0vnENqgDAMYbYSFeNguhYgyXWwnz
fKsKHw/hAn1tvoYxUEEguC8QgMrtCqhjM2Umaxvb5cPuwFfG1KX+HfI4HFvQR4ReU/zPIPQudDwc
/+O6pWG0P+4NxTAsoCYZ4WTISgdvZFW+w9ojohfkJfzaT7rJMgJCnjRhycsu9o6g3XrDhTu8mE1l
z4QPuUacsrfJx59AfQ1kkgcQ2AgjDYkr9c6F/wTTAw5ZFl79q91FZutWZYXjlSdfn2oE4cJNDlxp
xE+5Rz6O3nWrbwocc6qgOafQcMeyUSd1WdM3GPunYmnKY/nozIxeK7m4R4guMirNhsDoL0UKYQK9
JnguuLb1L+OKrqVoYQRL0fZwpyaYsXG0fZPeE94U+D4PUEDBVeUX2fmsg4DsTsZ/BPTEVKKyNZia
Hkg8ziBBNeSo4fbgmbzkzIYQBos1G+OApWLFs/luMO6nFIHIdxCYjCQLLz68B2a1J/n4CMQP+T4c
v88r7TpRXneE42c+8Ro9KbWGJvRPzvD8t/QA2v+UOHWjBOd9UJ35/ydoU90AUHzLkuu8eDXLzKnK
6C5Q7TN6tN8Ex4Ghdr94ksiMVzLd1WX9cQR7QQWVYV2E/+XRagRSp9J809sTKzKzk56okixl9xUO
BQEkx378GD7N4tPa4X8huTMDmIlu8r0F/JtBFkzxzJA7HXfBCS9C+xdQ+bbXe62BPCFCVBfzikFs
/QGsFyD2Ekbpo8KF8K8ehriiOLSX5/7ZwiRVfraueIF6XmGjHaD7CWCei57UzGnYgH6A3PKZx84F
WCVNVlEVL0v4UTMLDQqfwuCM/qLx4STu6/BpQP6qAGXxXE7bzBQHIIXZUazdmpLigpC48Elu65kQ
i8fLv2e4WPyhU8g8SZz6hqPA4c86g7tRTaLsgq9R5z4zvheEnYTgG8UztON/4XStAwTviMvpXnae
hYs4VUd4TxxNN6U3QirsrVDsJqCwFTUXQqsdcMz/RklVvrjBOBNwaZ+tkFdCFDS0PamNL1EPCgBx
p67kXAKxbQLiT3Fw/k0W0HcitVDiZod+a7B1WTjzSge+ebmvRUMxT5JOFYbTg4oJ5WAMbKt/+/Z/
2IeHCTYJoGQ9z5HRqQrJQWX6Fx6F8EOo2LXT68/LoRax2BdvNa1eJzVBTgPdFtVPz7Wb6sTn+C7e
B5NyrChvBBgRPFslfjoeP2od155OQjSBmZ1NHnOFQioJ2ul8YFSQ/iBe8vf0nUUBFzwV40WgNflG
ReL9Vu5K1VRwmL5izzNRHOp9SRHWO+md9v+hfhhVxAT8GHAc/LYvnUxtU3bh7jakIXivbprrSrsP
F64axoQFdlysL89aIJPhwnF/g2LdUpWeLntbPYHsQvQqXAiYGdAOxTjLltBsVyl/izdGMq/i4GO6
S/K/1L/9GHNWXJYa9SVPjkpI5wXzAltyVd23+X0Y4iQFMnKF7MrFoSsvtssEgwdkDzcv2Hl6EYUm
2v8egf9y39BKG+Ol69avk9BSwM3842wHRpfRLkYg0Iol5ZOAb0naqvduDubAwHbzHZZHmpT0KVAb
dXZfG8b0OuX+/Byc0tXLQYaLFue7WHlfD0KArZQYsFHK3s4y+kHSV5ZSSK8Gx56f+PCmcoHQujQp
X+YFvWZvkqyMVz/OcFPB4GjP1qs4NTYu5OCi/KAAPB26+c5MHZxVCqMoeq0G2evBa1Ms7FOsWQ0O
Nu+pXAcG9IlV17Frs5R7UjjL1nBkS7krTEVyLskKy/X9/Wu+lGJTVOSOdPL3FCJTOP201i+li+yL
A2430h1F4dkMUGcgY0z+W5z7XYaLyfGhqQrKGgkckgwvo1TQMm1d+JhFgxOIBtL1Zx8IaIxRETCH
HBa08oQVHR3eJmkrPvXFHYoCtdt/GHZfF/kyr/vLe/fO4KwiZ8fOO2WwUk/OGWHCXwJ7vfJokrtJ
pzemuTNGvg4wTrfKzFprWTz5hP7qH8sBkLU31MSmBLxpdWX7Yi9/Gufm63Wzow24Rd2qpouSd0OD
DB+hrvNavx8WqnZe3B1TMUiKMxLormUkFSuiddAfSkaYJzDXmkJk71S19GwYkrwHT4X+VMc8K8ma
zqh23I89uzypqs7lerYbw4NHKREl78esacZ6wrqGiy0V+CYU0TWQPZRR9YV8UyyFl0AeBprueEdA
K0EpxN7JvfpXmi/xW5aHPaxFolSxzRrm0O1jBFLSsV3QAGxwEXpLO7IbCPwNpNq6sQ8KkqiknR1r
b/08TpQhfygNxlJ+64tsN/K2aSoBNIPrahkkvPKbM+rj6KOPlZhfBpc+TJGzvjiyuiVUXfoF+JA4
PoLOVO52eo8H3FaNd/YPcq+dyu9HxQHtQZ5OXIInHwp72IvHH+5V/nMZcx1Gk/Xce8xmlVwKpAur
B0z+a/1kVLzaeaoNaxSyxBJQrqnr6Tr/3BRrO31bccC2x1pr/vRICSyI/L3pUfV0LN/gZN4sxUbP
DKaWrfHgJsZpx7r+dndra+ZmvuboOXCfjJTzqUlAYGSuXBYszdDZGmmXk9VgG0WwdQmA4I4tY8bg
I/9SPrZWavB/tN3BFd+yWOMSaiOZUMNrq8Br8uqnXSxWBaUDPLChAk9hhPhhmDmRQk8+gF/jKYJi
NKv9QtcQDBVvwDIkHX0d5y1GaeEw4c035XxUnRP/d/ofkqPHlJqMFEnGB6DTmZaExykGz+xLKvZk
6sJcfsqiP6i1zwGWiE3R3kXa2CPD7akedEWujs4Epv7XHvR+Z1UUQCc8/qvynMxR3JE/vibbP5VL
s4tHJ1ev9Wwdi3y55rkF3+vcQmFsIl8fMaHzN0NhhKnFE1+iYwV74SyNqE0mWMDlflvy/I5F2mKI
zQAd73uEZtAtupFN371Z7QvCqIIsYvImn0ivwc0BNHEmhPBb/2zO6OdFL2zojZFMnDZj4Kjh4Fj5
DcROPBYcAQlrkux3M0x9ZwPd7wYigaJbqc+DM5ijvJkAs5YZ0l1H42pUIlcxhsPmBePVota9EdNx
thY/IODW63d6O2REUk3Cq50Akg9K+bX+BJ7ibXNvmSpz7+cnj0xaSHkOfROJ2k0d/K1rXwrwF9WL
/6FnVxwt3GS6fnTZcnKSCsJ5iJDwgBJDBQPJkXaTlnf9UH0mXMH1P+FGW2Q+pQGt4JWfCpc98lez
faMU6LZiE1ZYhgmS3V7KPF6xclvvxHAARTkjqWTCAzATLUCwyAnPkiLLOmfnuDwlH8h0pXZ7Ktj8
u5j+5T7ZI0Czb+WAdOT9h23DP2LvLZzl7QUXMdIoBKcGmgD5zaHHyOAifYV43PSCyATf+5qcSikQ
IOpXEeawrgw9P04UGei5cKA2TvmEMgffUG6GQPAHgqtNeID4ml84kwYmVV4SuoazcYgmT+iSNIP7
tJAidxE2It0FwyQkYnrjQnobZvB9wj62Stg/L5FvJjcaQN/4VK/wpQA6F68tm3eQ1ckvdR0oLqDd
4G4uz8tkWHwP/x5aNeVNtcCZvonpzV3othYtVHX8b5hD4BOq+TC5QmRR2Lt7dh9CN7hPFJpX7AKS
qkFcsaoLgsEReUvRsBcPiVDZrd4NhcUDV/eusoiizz7rdJ1Tf9vfhSwrKzu7lVkKG/VkKlnX0iNI
EtKM9NSv3gLcKZ3RZSMpUYQxb860yzmQSiKKNBdnUw7kJh0oudCuZZDDiAW8DTILZOPN9NkFzCf3
pT8PKO2pKL1YTebbAevJvgJBHmdSl5/kYGqZ8F0zq/DBvcAxN1pL4FcF5SSkOMmNzP8xLGoeMyfE
8Nexl2cggDvZwwN+wnVb3VSv0g8Ljv4Ef8bWdG+tU+0LhHIiJUyOANPE5y+muuzxdjt/p6W2oxwY
OuQYc5FZjwQQ+4Ji1paHFm72wWc18lfwJg2Ek9EI/zCTRbkeiiPkUcT0h2eV6VqDeMzeQqZC9XbM
HFYweDo+/qgdqIHfHDPeWVp2qUu/Sk3HTGfLz2zlHCMQET/9UvIqSz3xin5EtVmfIMQ+T1LYHsu2
pRoF5NseDCt1REkSkPIC5pQsWv0GevABCtiSEkIpYD+2krbGL/DH6AMEAX8iD9yFpstK17RrRA8m
CCoDYmi0HJTLxm+ybSeXHNfJYtX049Y+AnYQ6v8tc26GRKpaCUvi9c7O22Eayy93d4ObVJiumxpY
Cvka7hnN2n8lSDui0Xmldz8wFpB5pQsKWm4GIpzUtQ5ncWNT6cMc0biwx0T5ZDBceH+xEhX5k2Lx
2tFxtWBhhQ5ipR7qw4Emx7pFKeH1dANPOdV43mhfYLXhzYRK/uadY68FYDIwtzgWC4heP+m255bO
K+UnxsIITezGHvMmlDqX33VS+X4gxFDZQS9Bchco7C/JUflA/ZTz8MENHzjqvdBXSDwkITg2q7nH
ix0u6E58aUqpKnZl6mBBgGcOPcKyqjdgib5m935vNkR59kfOChjJeVu5gghYbYcVvMvn8dPoBRBF
U144ybOvYWJHNHcM2bY8UA1UtoSNbCetHDK3LcLDVmM1pGP/w/NG6EVs2UL0sQRCOOLC4DnFwEM+
r8R3/vIcGp75KjK13KG/z3vrNhBH6liB6ACQVftAxtXYzlxOIQXBkDdPxBOf3iJ6vuTAOZfWhCfH
zIn0sxZUnQHfL1Zlrb0bdrYlvN847TJDMnFhcUrrgBQnI86xUGkSBELf/fbgiva8whUMTZTfvsyn
OOryTB5Fjzj0rMH4wzWlexyOtD5GuLC4k0lioa+FKBKTq7s8QM245a2yZirzJGazls3jR5ccCht3
ydR5XwkYy4IoirO3ilZt/ErmsJwCuZYRj7FV6uuCneq6yBd3Y8kwAh4EeEaafdBDiWZsyBpv+Jy8
U0K+nWIyaDXLRS4RYmLrKstw1rzniPGBdju7tjTYsuRHE3ZVC4MGCt84ey9F2Y7/X9Nh1qEv6gZh
Aqr2WvvcK8d+3ms8ndshEgWgVTpejF52TQ9qmb2PVq9t0XFM5693XdlEdBg7uK9JTrfbBSgkGZhO
24PZfk8Wt8LZS/1+uzLa7AJOq+1Ke5KkUcAJmjrWhnA05amRC5kcbIbANFXgZ7lDU9hEdlgYnV31
8ubOQXIpSL0p5cZr+Pt8Z0fDNIzRhBmA66ZpU0bQ70R40xoXx6j/39yx9wZ6KK+Fc/QCer71zp+W
FSUVGvKDRQKO5BwQt6sJ+o/e081SpBgwHSiUeqNqQAYdAX60A4Mw27xGeqEO7XNsXkAHA+EuyUh7
4FZWLUE0+YnmXV6WLrsvE1WGR++swpRcGUKkRfmsFRN7Voom4w0Rf02KjEwOgfXx8WJzufF2IpWQ
Ruy8ElrIzQwowx3vX3ZWEgFqrupVtLLbmVUayITAYJTIhddCM+JNIjzKZCqx296n+UJjfQaiVK5q
6aJ/qQKmW2Cu3q9TNs2bB8X1SRwLk92S9CLqGoIPTrHkKQbZDbOblVDnNTtfJb1mcmEm6oJAx31J
AXOGlto+zr2IMWArZIaan/eD+VN9j5cu0SVhp4AhLNBHNekYp6DfdSLTFWTWQ1yXc6GUwJka5/qd
in9YttZtpT7JKdTjko9FthDd6Jk0Mjy+MCrIc5Q28EWmt/4RgV2KXKskVaJix0tDv3jNJC77OJKl
G1Of51K9V1BFGjaceKB5BAdcPFx/IIjsl32TWWoJjwzVffmQTLJBJWoGHEkBnaoV2zKUg98wnvXQ
Bwl2zreKHjIwp/bTkwcJ9Bsc7PLY7gphpGCEdleIWyzJUxtgFd/xOHqlJ3q+X2WjnWAbDzvHEe+U
GDEBea59gZvh2jN+ZCW6DBXyci1tRNUDGxFgnJG1M0vxYWhgsM2jJO8NrCoa2vKq29IdIJbaL497
wiecmSVeNvyfDE5KJYWRHcaBHweo9pihSeLBm1MCkn3OvZrdC1+DEDhqzT+OVQ1CXTOGR1gcAWGC
07DQLjQ8UVn5QQagXLnKSx5QKG9Eyt7sKiua2X/fVwFkgt9hxoHjbDhv8cTi4Sc4h3ZFu+Rte2Kp
1YGdx/GnzgdcnFSTEscfyMuoKopkULeT7iPrB8f3Oto6lXgoLPXltVDh+aegZ9Nh4PT/u2Wotktz
6VdfUcu3kklgEnk2W3wrZVUnUHYhI+8Y7TSn3jvWhvAgG4OG6JX7quTpNJ4mGfFlZXU0tfhnvad3
Phq83i2Y0DbaQW93K235T2Z2Cw/0QVxEX8f25E/5Cg0WPerZ5S+onRp2BNy+7ASiyVKMj9vNddfR
6KyVpRbKDjkJW2saRlk+2kFtMCcIODGZSIgvOCON4hnwOlkQY4cT+nh9YMA8A9GQkfYdJa6SJb1F
JCjcd9qI4357+lbIPsIGAC5DD9b+4ks7Zws9v19GAXTuIlvPhjOuf6SGBiSjJCzI3P8Ki9a49e09
yqD5X9BbnZDGkGauNT6jlJacZCCIaOC3Hh15hUbO9FKs55UjYLhJ+iof0G6i/p6sYTPNSbRonhZL
BmY6Qbw3ZvybPVtXuJC7AJ3WudL6RBB6TKTQ6gdcTFvyXJ4aJVEreTBrA/UeGuT7CV0RhtoZyG7R
DWNsF7OsVNKZbsNgDQeJVoWt668wnBu9askHA2F43I3+6o+wwmCQEItUlRJM/OYmDIioQXwvpGCV
HEBK+Q1sH6Db4r2uEA+KBPYdVBddkeeZzHnWV8Tq+tD0e/n6sRzLkbGzYy3qF4WKzBrqKr7n3RRX
Ej/rm0bEt6AmhyBH/vFwmE/hQt3pgaXFsKnkukgt3h1LX7R5exbu8HGaXiXKS6vdlvOUWvAkxpSf
SMq0/negoHS10lY2uwm3L50cVc7Le5dG8UYDKZ/k7idEZY81ZSfjoXidw+6fdUcnfpSHFiX8Hf86
/9zMbShm+AorgSUX1zSVWHMlHBlUruL6zPX7yxh0hqlzDfDdH9sL7Tw30g+1jAcv3JsMz5L9oIiz
NiMpp+8qFS+sJHuXT8pW8mCh6xLU25Y6sZNOHvq203bW2O+6hN323beBH9oimbe7oF64ZY0rOanI
qv8e3FYWJhq4AlZXcnB9B7j2SEwxYmj2MDc/jYS5AxsnY9yVjTKyVVTuOli5HtePofeLk4nwaW4B
pkK43CLkS1uifytfEF2xuN2QB0jWtSyqZLvwX924UMYv97HK9GoJ2Fb0KoUnXy2YRllluXgjch1c
BfwO7r9qDounzCwCa5uezAelU9N2Imw9YprHwmaxsqqoChajgVEVNg7cUPDEs31bz2MMGmjR3iYE
cXWIvRh/pDk1t2eFB9mPRnMI1R5wQAXKs577772T66cqmvZFfhxUTo4kp5aophtB+FAkTCVt8F+4
xIn0Njz9FXmfdpYt16L9mnjDlBP2MXjNp5bUbtP+/StqtzteHVwu7Ny82Ef0+WByNBQWgJVund/h
BHedKZTGkAPY7Mp6cHlVdydApPUhJbV09nsvU7vA1SIiKw3a+lnFOvagas71qBV4oDGLD79rGvPB
oVoSEaYPxB0ssbmAy4rGJQf6qEm6bFKtRi8X5lCX/px1AHfT45bRzi6JaqFcckcf3oB5Fno7sVRU
sWCgg8D5WKxR92ib/JFm97ZATzpvUA5imBR8RShDqsiCq70JhwZgqr45xFAd8hWQw41S1/PfN7Ht
vdgi3Br/onvd0yPjtdfwhzB6QPnqOY0h5jYWaWI/b3suiyEHRTsw9XFFEzIako/kDbhfh1RsNrBe
v5LagMc85N1rwHArExY3n9YTrQH3ISmoVkVbrO+UNsQ2epcp4Zf7n+h4+7DStk4VUSYqmJM5/qIA
uWjTeKUM2zLUfU0aR639bHaf0XcQAv28yvKtdLtfR4hBL2Kf7iW+LQ9gtMB0Kvs4v94Bbf0+cKmG
WowKzdDqGt4wSvtaju/jqo3qz0wRBBuUilKX0ch2Rzwdx2BGmGe1YCFjBqZKrVSsdTg7zfeT9+Uv
WLC1zsyWHRCcQeZr3D9UTitqI6NgDO7lojRvaBomcq/haWUSKJbFJxBxJy4VHc4p2q1IzxTaDTz7
kEKSIpWMZwrQpmzLWUBQaODepK9diYbr3lq864xV3Qkx9ICPKifLssdLGiZ4RLSQp+CVAI4tIWLq
XCDGcUR1Kp28Y/cOegtlsuvA08mY0HIBK9eT8Q8Zv9U7pjDDctDssK67SLbAGyObhkqpzlcejwE0
us0ss+KDrrGSxK8f6tXy0W9129bkb5hVTEe8nwhvvlOZLzUrtwc8DNR+G71myZtIZqaBynP0UjIl
GrdhGKi4xi9OjDm+BgWs+bv2BcvzXAt+4hJDb9xmI7+WyKn0BteglmE4i0b4Yw66h7dSCF7Z44vG
dm0MKTp9Y8X+khXjj8L8e4OgeLHJE0uoLsc60w03qqtIMDYooP9/jRiFOui2xkgG2ZAYYpLJu5wV
lAcl4khdOnm6ZJSIcxdsWt4fS3s+Lwr+DUKYICyld5upTOgoeOBBO4d+vNnK9zjl9Qx5Lt0KLj7O
zFB+gkYtMJEKs2M7ASO3OhMlvnzSwBndBdpvje9GxdbC3xBaBrg+E0NwIyQGpifmJIDcc1/RWdkh
cdvnEtvC4bwa7uYWQJ4JmGj6IpBTrsa9ga173VwZad9kc+Jwg4RgCoTEr+6cwa5hNaIdVEkcHvI3
sZRcipNze7kjNXenDEyLGMtGo6I0NKiV6l01erIifSG2gSEfxekydQvXf6tMIN0iLkUkBFgedQyW
UWj6AZv2CL0kjIQCnJXFXc7gtSmYdm8qNSL7Syp7IDo0W+z840okT/iZiBE4kVkrV+UliLgienTD
o+lEIJFNlhA7tm15/+/jXyXAqK4dYoCYyWbPE1k0Qjhv3dXfwtxGSM24KTDTC5OWVKQoVEvfL0qD
Jgi8yu86ln8F4HE72O7HG3xADriBgVmGZ4cz/kwg4FB9xMORc0eDha/Qu3ZHfu52+6URQwW0FPLT
LxWQXFP+Zd+2VMCgr3kPgSVztSjI8cLDEbYoQO6YyJeBOpkym736V5nwVUR+q853BLOp/B9NR1gt
2PALbZJJYxnJNz2nVcOsQ+dvGY/Lw+3X5XvQiU3fpZALvUAqRiwYhu8HyuRKiRf08SY4jbvCy7nY
FjyQfv/pTncQVl0oiSXVeaneKEh/a2ZKZqALLpfykiDiVDxflxr7tNKxInxnYsyHASV4bzxAqYr+
eFcJBUVL+pDVz22WzkAV+6s8lzaw0aDM92UVUUfzT7PoO3JHOrhio2MsYF9KpOIs8M22P4p2mwwk
pLe45ymztAqBXcdNHPvBRvHFs3Cao4V+8ihzcRLwTNfVynrZpyY0tTk6HFV+J2l2/VVUtH4rSUIo
JlE2sGvi89lEpnGJRBS/9msy/2mmdbE64YsUqyBoPtETqVA1K3Z9ifeEYFcBASkLx8spruOXbKvg
v9ehSsCtfZIZlwJacyet4ukG0flfY1j2VcSolG620yM1lBqn1HbRB1kvQLjam+QkNSkRFkPjXOYP
5u5VbAgga/4RRkBSyotAblYvea/Ec4hII7ZqFyvmFXLOuIWTJD3tNYu/DSw1y2sQwtMJMdKRfLdM
AZpw1u7WpLvEIP12pcgm8t3MIt4jyq/PjBPmqKLS3QtZEe38p0hrBkNkYUxjyYvucjPSr6Cluxvt
+nOBf7MiHjbRXf9vK7AVUI+x7ZUjg5HdFasioiHJMer7F2j7Z7aUVJzLF8NYQ29TpWWXcL+tBmLA
2kfjhvirPXw98GzS6fkTzbsAfX1BlBr4xr7VMDkYhQ9BaoHSztqPPMC2ppLdWQjcJrRjVQ/V0iaH
oVPzGFDjF1AoIe9x6dHIHuRNsa+JiovufXY/yhr8ceTt+m42SQeWDb7UY4quYNxhF2na6g0CVS6o
W5m/Ybdnzs0uKuplj+7DXtbt8D7KC+O9ilXHuGmcIgG5qsi/iLHa+3e79oBh2KsVegAX7NJPdKav
f0IfGzDY9n+MTnNGobNiEsgkE+Q9QIsV5ZQiPymf13wHte+iVmQsU/1UPFsuJRlJn8hUHmiYsPxm
QntUt0A8fageUqVbEtatI2ajZibzWm/TrjAl1A6Ohu3m/leu5/QiOnJnf96MK/V0s/Nzr9HOCU53
BVyU2yJnBOOO9YyZyDKBvsQL6uDgD0rxyTF5KLSvYlsrv5wsJFX7XHmy3bp2bG9TlsJSz076kan/
gr4vmAcjobAvzSMmuvQRtKU/YaySM0wJD9RCaQPYaUhDJlOId6v1+srmWaJqoLEInWmrXQCQGNlv
DUOkc6kTpGyIMiOiceeyO/xetk3F8QWfCEtU/n57pVuZEIFGeTHelMojcr/MBi057FbhpYdq2stP
CoUi0A33v0lRCp50ezi4OWJa2x9GT+ajwRKyO/fipL1ERg1VP8QsG3zkLBMgG+EKsQ+Nt+sTOfjV
lIJiVzLHq1hlvIhb7sHo46r/doDLiBJaPo0gMVKSwrdFkXQwkXXZ/jYTb4AJ8ElKdmPKH7NOUGAW
4VDYFVBdKDlAWYpJ3ckn12jmxC0tim+dFzQ0vWsf5Ra16A9D96YYCAfi06Y+z3prL6pBBgGhDfI7
Fwr2a4Pc8sMDDE25N8iqt2kwN10JUOwqUfjNWeDj/yn0u/koPQ3rXXDcsVvCMOg1D2eNe/nIJweX
pMFI7PIy+aKD2Wx+8UeD+XkWi4OQ0MBRi9r5g0uptGtrO113GWBrUOq/XI5CQVPGdA4RXs/9HCLk
pfqGrZQx86fmYWQhY4vlQmIeqVfhFM3gPk4F+jmfydZdwB96foYfmkEepnWK2vR8ks63JmRPYViN
SHnp20se+O9grtJARfpw+ZCBnC0WdRxu/uI44Zo3eA8aNKacscc+Uwg61S3I3/aCJroVKL1zWYqe
+aThzIDliud5KIMOPqav3+eDKLG8/1XA4u8rGi7wgZIa5rTHKZViV2cKHgfZmMxOTRDLdlEdcAue
1D3xtnLDB/fG4zCQOfYwgodOpl98A0Hfn/LTqOpS0OlUmKf1Y9VvSnhkIFk3vMobRYePqTkj/TA5
AayTRAKK6a5F5WXTZBac+mOin9OK1/p6TsDDkrZXKHA9hg4gS5lg6+0btAvizUeuvvDU8Mhr/7ZZ
L9iJ24edP5uOVsMN5+6sZ+RpzOwtcfbAlJr3Axm6qEk9j1wfzTMPHXDyYDuc3nFEa6ZlZzLBQMhe
B2kkc6q6bZJ76E1t/5xXpeCBqNKQFORVrDn1uwe07ZZCsElKQvlPBWZVlfoFwRM/EZRGnNtEWcEZ
OI/kPgJanVTZ8tvobfJgj+6NF4chKSnfOcHEETQvZEXkANpQRf1iJSwlnQG4GCKdHSLwecsFoqpN
HZa83QT0JSRNmi4hd0MUyAZGOlQf2LGI8dc/x4SHdqF9N3mp67F73YHpqa++AuCHqiDgD7T2FzfC
XYPmvPPun1V0piFXLrE0W7xar13EDzYvlaQDpJbPuiVN1LeKMuU40hR3ic4lTbQ33Gss/akEOpdz
DY/rfXKew3/8F4IXytTX22H3vCmZjkGiKHAy/6437hgMGlPNj6k/WCHxaPY4jN8kg9extarvpnUQ
/J/LvbpaBqNYMyrBzAGWdeq8lJtro2e9nzg8UqG0C6SXdbFNXHHJT5lNFrMgmANQWCw+6kvAU/Of
8kTY/7Pu5oUco2kgVWGk3aBJxlHj6Pbokhg/D312JWcBqwuMuArAplc2Patz43dL4p/tfxsv5HB1
OVi41U/NBzvzAz//7ljHp0kwDGoHhol1BXMd5Urz4OzPwFxH/gGVIsKh2IlSwMDqJTM1ltpJZxlX
lRa1iIYEXEAQZAZSOHxDkdRmDMfcl2R85qerL8cBcCiiKjB7FFuAURC4pQngbTRd/GQHNjkOv/Jg
B9n0UxU8JsKmuhmLQ18Vzb6Y2hGjtn4r+aOtJjJa8VYNbU5hnd6/lhMzB5Z9Y8mQSTc64wJY0ops
1daff5lRRMYbxbAp8BYKy6X0tsayijPl6VzPy/27fer9LuFBCdQytFfqh8sdRBpY6zP18E1jgeGE
uAhI7WwRtx11XNtqflHgJvko5PoPUtNnDpu2hvya1HTjeypRhjnwIgBcuov9vhuRyzHfNLEHi+V+
gtMVBorxxMEsf9qNi9TTBzVymHQG3JKn0H7K6r+3qU+wmgzJ+GehSbc558XPzLOg09TwIDgsnEyU
tFRIPFwFJA4aRr4GYMWlaP2t31iTL8r/75ciWCETUKOCwDgG4GxupPoheYsQjTK3XI+ABZsWrVj+
vskWWuEXe9hCKtDyVg0bjgASl3zsjXlMd7RUwMpLgxGA8YwBVkv1+gq4sA6TBJgzfqacwuKGn/f1
nB//Z6m+uDQZN/UNozS+v1xzdrJBlE5JJC/q/mYZVuXgpfVXiWg4O82kitzGGLwzBVz7Utt7VVnd
/DtN42SwKU2TzbzbdZrnOt9z4kByAFkMCQJU7ARjpUvtm177dKJkGrV6yPImzxZlHuWM1AngRfds
UAwc6PZ3w1tuzu7ifAFb5YiL2jyfY9qIylSb3c4Dld/x9m0fmLpuCnO6oVO28GD0PVQmwllJECog
T0N8yXR7hyWjwwWn3YbRXMVe+4NdOcX5i/8LLfL5nJMEBKowM5nM4+wHvIUBIMYON3eou242CSyL
mn+FjxbHe+jH1xCHniXoD7g+IogZ0ijripkQp3lGQzLPzFS9/mqCeibrzYv+28+7+iib5g+3YFY2
J1jRlxAo8LUAPOqgfVXN3y1NiTcMXqRnj4LwnrEpoZqFqAgyWMkQScZdbHekR3YqFbh3zcQLsn5C
jzZUUWPw2Y/BSsnEv69kklxOQ0dyAt4Y6DSME2mRwTCY0A+2vm9QiYKVEXAejODM/OKf/fJ4CFti
AGwVVq1Pf8dmjUb7RM0x4sscwkCxeGEMev2d4AwYTmpC3Kkan9V2/RyJKUmM9QIdNgBVfMv6zvL9
U5FrIgdbSKY5wNttf2UVQ80VD0HomkVB9Ri0kBrBb4S1pit0rONrCNOKVAymbPepirFsuuTlLtqX
jkN903GRmzY5l+JezrnImVkOQdUHrHJsAF+mlxrfgHqMTtxzCEUCI2z64rZO/81uD8aW4VMQipYj
m9okQJP1Y8Vy0NlxPw2BkQo1CayLT4tas7VYun28yl6fZ2cV9hcUEsbHR5bkKkCzMEYL7+a5aYAl
h2e6NeVhcBDGaLPGu+MkY0WXuMqq2aZCYxIDbr1H+UaXqY0pOOVnXQyWGvXeBA8xglEoX7Kv6jmh
Y3ASxtyoRzIpqLs4E6JIcSx6bwUFgWqid6124CqTM3u7MAqobdBytLcY4zbaYzjIbbcD34/9EenB
iuhoDp1QEI+EbIBRZqnrr7eXjSvj1qcGJmRfiBuozN107w3PInhrsIRkcyq1t4QadeqdXEhHfy9O
qOpmAvGWgT3BB4kLqN4NxpyTfxvMf6Gnl7mpqfvG5nN+tPXMzYZ7P/PzaqWzUW04SYJSoXqCXmEz
hmVMQEh5AvGIkWEUp+ppMH8cN6fo8Hm21p09agaL3e+rzmZdgtu12GUqH8AoZjA7kLj4Z2mFAmyz
49MzaF76YJMK+bIXcwJkJE6QXs7PXP2fFKSEUcz0gcNAwTFrc03AM5+fXkTRB0+ue0beYBmKDtRS
y24tlXrmlg2O/dGfx24V1gHsl16QokONtIYQq5GlEYZgC1cEdTmyNjmvBQQ3XTnmV3aagPXe0s+B
jY2MdIpNFU0Yh07YgxoKBO9olcYwla2SnxqPmRiEpLJ4Pj6ndxITv9gdH3bYzNNkbqdBnrLmaHE3
VC8AWHY1aQHW21HoFnS6N08rul8RXZ6M2AEPP1XS7Qe+2HKmd62YW/IH2ICB0+yYD7ey9FkHKjOz
asdBOkXPTcJWUwHTMIhGPGP5BiuB/c2vK2AyS73z43/NrJpUnu1+lOxiGbQD6AhZgdLgP3sLIUn3
TiyAJ3URjv8Dw7uS4rYGgPymOd+Fss5IgyEWLT+Qf6vpWxYtM8nSMzuBvVBBDtMziv+j+1ERz/aD
IO1SGvwZbJxkMB05GI55qKtnYf8Mbl6XijxXP2jGVOgo9TW0Ghmwuab/VCgATheNl3WxIEnFQzfk
YjWTvbd3zgOdTlLZb3jIIAo4ZqKVv/R0kQi5LiB3XzM541qw9HXsiiyf+9tF+XChfYWAc8fgPpwQ
YCQs1pDjk17nFI43iLOGuAduW6PlgIHMEVrQLyMGabiP6ih2wR/8i48wCe7LfCh1RR+zjiljRAWT
biM5yvlG8RdperkBpycPizKhEHr1iUG+wlIQLatIixjIXzVaMfBTwXJ5Y38+m8svmMxPJgTPZhmY
umt7JdEDmB0i/W65N/nDd86FWcKefB4CplPh2t+yedG2loYbhdlS7TlUJ3btw3QqBBxCKzF4vyxi
+BWxCrhFPbMyWToBhPhyunAGwEo7yT3cxGk/pPyJtS/6PccWutPNZznawkQ89qpq8W8sagglN2ja
6QMCYd++FtYcNiIt3lTzhn0L89qiQSYmbyUSbk9SmXU3Y8yKf90CoNOodmEUln9Hde2ecfMlkwP3
S2gm3uU32QJQ2uKWzY4vdDHRfCmIPl7qN/VAHAhxbxVPfNrIubL+YVc6WoAL9pMAVmlvyiqxMthD
lJJSXPU/BFJTFOz4cIZf87yVCdtF3iYspKmHoOhvMM2p02WtUh3EQzAPczxdQwJlqhM5Cx6iTP4q
X0EwxOTpwHpr2UYrv6jxcS61Y8lZKVM0UmXt9LuiX8bhzfnmNoumXLpVeGaptvs4DkZNNSDTYhY0
RVp5jW0HlTpYAtSsMlYD6yaqdxHYV0hhpqSPNiuXkh/HJOO7aovcuIGldmH7v3SlnxluTqTQVIWW
XAE3kMUPrJK8UCn0kCX56I+40+SK+97xY3F0WgrK0UY9ti6iopKtVJhHnR7BzA+k0cRI/qpCx6MX
zgBzkMRex8/rRJmMDJ+mOouU23oljlw2ZzbYXu7FwNNTUcebxH1qrZszvTrJitLx362OQyYSONph
qq8arrhRNwOIC82jGNsTj5Dk25jwiW9Sme55GrszGcRngEhKSMicvrOb36yzW6qj7TBOKHhroDV1
Q+0KgXPygkKXzJroWcQnIv7JMNL2D3kPVFhZDmfeuMOrmoE4hgHw+LE+W9+uPwLnXAtmJXGt2Q+S
hWb+klPwxqwrwCBvG/reQPBsX3HH/njrqi2UuQbvU2UL99BscgvSxhlrPz9ox0ypPiBArS9IIoVS
XbMvuWw4YS8oNfA0R36yNq06vognfniNSQO8m1eBsazsMIl86SuW2LCmPJgw3hA5oSQjtxnsXhOT
Ib+jyBB/8TTspAfvqzVHti+bDGnrbiKp5rN+pLXIqRSnMnpU4UwDGMZz1C1EEwWMc//lgc2Kpv9a
ZkVyiI9bdNK7J5jWjsGzVKMMKtWMvU0Dq+0eSoDbHIBIUQ4Bxb4n3jY7C8xCjI2JcOwYNc1Teqhc
sbOwGgotdWcnHubQKKoM2UBknlba8DJfre++HawUuagOVr70C5Jj7Pm2CQtXYc/k3rrea+4qhI8M
2/facdctP2uyaBkRsZKfvMD5UFfVYzlkAul4hfZV9G5yos1t9tXp7j4LXn6vvwTNB7dO+Cfjfd+S
AabxOdJrsHRf7/zcVX5uEYJpX5qyATuDi18Bd5xHecxQBVg+3au6bWBtgCY5/9dKtsBVQpGVDJF/
6GH8AcGeuPFJB8+GKaVR25sA9lozwWuTpxVLPWE1Gdv/gN3NEZUvEuLX5zUSD8R5CXhG7RmoXu2X
2fe1frTRyBnrnTvfE9Fet9tstbH+od2UPy0dBHdhqN5Her+WENO0KkZNvdxOSgMCzLVdfnfIZG+x
X4V7EKrVo/ZyLhjh8lV4qLXhHqLDGm+ZNRjHEA6ekvWzkC4H/oruDKHu/plVmBnW+vdZc5PMkyuK
bYbZ+0AV0aiCIEaUY6gVaYmws3J3M04MhjpciA9+i7i/f9MXgobPLtTSD0ePkWaLMAgc6Jo0/Dvw
tv83IaCvcHxe3AmRLIAWs80g70NDh8CsGr8dDGjwP483/RXhANw2ymbSzrENnHsocqgfQcH8A2l3
QcrvXhKODdKLf0zxuLZXPjx5FMR3RO0WLwqhxH3Vy7+BwWmViuPMDcPWhWn1mFIyBVWl+zhB87+3
o2oTCaUyswuY34pXf9+m9REOuj8KYqeZOM9L1pHdfou38JKoELQTtxg8fYUsNWCgG7+EinejfnP6
5mo+Nksd1hpoGHZ2/dDwkQSJAeLqu3/p1aLIdPOWRgFZBxIRoukyauj8+g4X8Tt6OTC1TKlBrSYh
BRjE9XwurNf4Vi6XyLCJVddqCSIeXdBDd6NZkJCTB5Q7vDRoHlaYNXtkp81etkRcbOEy8MMZj8y7
V2hxTVou+P/4KKVnKz1d8ylYuGdOBNqb/q1JKxSF2QKuxijW0/dU/dwUuhe3/DkWz7ESOj1olk6Y
/p+XFfPfdmcBcoW2crzvDS2ymDdvE9Z9ax7z3BSmJ8ivnkMTx+/BxmYl7XrPjgAb7j/vEpHSA5Uo
aOVlRzXjybyqMtGfo1KmPaYDvzarIDwfjWnKAYLpPyPUbYRgwpMEXfOISrurAR+DAgM5/s4d7Amd
YKoaZIxT/iwIDv6ktjOJejrJ+NVPAP0nIFgRzUcG9g2jm9BxeEGGj1MKAlD+ok/jlNTFtVfkShSs
sIR+MeByVlYkgY1fGk5NrXUE/tXioBC0BEW80MHJXapzc8tht4GhVXGBilJXb1nlupB0v3j23Qvd
ikXjFogR9FOSGd6IS8oU9/mtD9oKb29C4sQb6Aiv/jTtUEYrskPeCnDtKW7iFXOyzsJ0CrMaBr8j
m9SqGWSc6DfeLWewVpB0P/MsNDoDhEVldCLFrM76xM0NJY7GlOwXasa70LF51Ro96c13YiHfnKui
DGRc9gA3Fwt3ECssTYdohDs6JSBLvbLiYmZ7P10/zURqn+ap2ST1SVk4sstFugX+SL+4UGDip7wz
2DienKCKDBVU1cJmZ4jPHRIRBvUoYxgyG3JAHzx1YZxFy/4oFVFG+FGaaltzEBvdZriwKkZ5axq7
TC5CNm32k9aRAKBNzQlpvyVDIyNdYiH5oOfRpa4FRa8CnkEfZRFQIod3wu5dknAAaYGn5RTItmRm
wouU1DCFh1YGhDbsgzFupXui5801YlaH3ux+bPH+Jccx31nsmqwEkw7sWOHpAlayf95fWpj6IasE
qAlZ/N1UYm7t67zjIo6r+SqqzC3IFpMbKNzsCGw2HlyJg6DJAwNibh/mqn7EjK9JyISIMXwzw4uv
I19wTSDbtuUNnpTuAOCoX8YBUbh+WEI9dh8OYoP+gqix+gQRHOSrAEkK0fnXO/v+/mkEalamiYdb
1D8mMVmqf0PNq1btMdev+7kUwi0cgEdusaOwJuaqW5GWV9jIvdUD1SiDukdNfXqMGntPVJLYB2nN
s6TeUf3nGSnfJxXXc1EY+Fg/OITP1TqyHXRp0h5yv5JcdetiQuJrIvwYAi/9dYMfn5t+PG/8oNIX
bf4ExZ8DGzjhgL9gEuqlpQsfhyZXiw0aLtK3tqtDtJJUEfLpdVL2wF3xM5j13qEtDjPccAbjHLo/
AddsvP3JFXgPxwzSUPwZa6gi1u8WH3f3ijCLimwki/V/DyfRE8/JNiaak7MuZ4bzF6gXYt45T6pE
RbiYmtDFFbkT/6axvFbQdxi64K+uSuNu1Zlyb/18zfwknO+qbIZSi251g71Qr3eGQp9fU/lQk24W
UBpyCmGE6VmgaH38CaBzcE+RCrXE3jtvY44a4EQWffETK9RC7oIP67BvgdrC1YHudbezRRKIpFph
e+sqCAXCdHJazQNR4ns4JybxJ8nALlyiMMe2VAFsLVwHj4VTPd0XLxKZKO6HIXSio3ckul/qSncf
3iJMqgOLvj3YAdMOwfYusnkL8r5dgJrkRQmQliKfvIxAAMGfLQycpFKSYjq5de9b4fHjBd98wOoI
wAE20VWz34pHKFk7q41+1tb9Mo1ENUW/rNhKB2ej5X4J4ncsYheYMItoRecdlKrHahDMHTTRvUHs
NVeZQE7ubec7iNZV6ft1Ud/duLlxdGAKWu8nmmDRaAijLxIcRv7hu9iCx3c1Lif0QeCFTnvcyJFW
10PyWb7lNYu1xKz7HJu76MJpV5PHxWbRoxOH8bV2S3nIL2OCkbrMY56lpiZcOFtBL1r5rptjkgLd
YDVk1HtQ5ejNHGJ5qjQSidaCqdrZyOkbvDxWnKI4GFg0B0NqcqgOMzr69lhCUie8iwsdz+r+rnlR
Vqk6gCRwF04HPeBrTGhKb4y2XV3CrJjngyMYHRxBbHKP8cXj4YyXggia+XekT32eqTFBpzFe5YcJ
qxk5z151UU03bYq7qmoHRY206R2RZaZQL+XhU3MTQqx35UKTcHrDg7Wtltk2Cz8KDVPigS20N8XE
x0oxf4TvnW3AZPXB1tTQFDRdU4oZhMQ/DEO9UpEXfJhjgm7t18mVb1KvDnFQJbYpDDOWis7Mi96u
OSCo8yA7UNY0vwfifKSydAH/MHhOvSH3kK00jeU9L1twREda9MHhJkXoewk/OKFmBdhGPqQecCrs
tJraepxAElhLJctZ+A1UmYCKCrnfClVYiyP3CAuA1UjiZNUXE0aC8qKGqFMgGTezbeBMZHeyatIx
1v7fmmFKS/4Kmo3HexPncvEjM8Wb/OMDLcibd9juUpW3OFLsIVPx/9y0xFnYjbb0tX5zbJLA3bVi
4LVdzZ69co46FjUhI90/dgSw9L4lcHHRNxVxe3fiKtdbMQe2aRReZ3zMvPhUYU63KjG/M1Q/BObK
tFVsnvrjTm+OIQ6CzEchGnPgkwvhGbBZ6wOOmSSmnbD+x2yMBkAqvjLcxx/KSRcFRC9fIgsWaJcq
6n2qci2RAAajoaTg7yaxcGNHuB25Vwlc5SjKgBmCI0jOfWPOcj+wz9Gd0kGDEdvgSjRful8DWGEy
uuynQDhwnC+eaQwrjKWy+Rxfn/66Ketl5F9CuS9OyBrtb0ZrN/NJFWXfNvGvhMk8LvOwc9B9g5SY
hqzvE5uGgW1QCdelqcg1JU85Y1Fc5+ynygakqCz88AgQEZBUZuDgMIjhxnsZAt2JwFvZFkITrbFc
m84tArHqCXIK+yN+Ix+6ppFQTIvEwIqHO/5d+b/HottA5LOgCAW0IXg/TRcRz+EKoVPoEyYo6SWK
Ajn9YDG61h2zCBCZbi7xFDsDmiGHae84Z/M56N+DKQmX/RJLAZkgd5DqGBiatSgraXmj3WJq2R27
aWTUfcvqZT0u0i+8dimWTwfykXgPNCaYY3AYNiNTv3sJtTGY7ZR2jcMV//GpXJgJsRbxJkyG0/Ct
ftLeJjV6oesMvTsQQ7rPhmQu1g/MCjNLVp7ZcTikP7/VpDt0T8a8mUbEnpkY2pCHHyDsGcE97zLA
JuHseFQlNHHGtqcqF9Hh1mRNWWxie+oXVYIKQ5asGQaN1D+3zcevZHX3AM+mK2B6WU1+cYgCJzMV
HVO5BGYklR31cH269ZbrW0vLAgfHnG17Hx9DTzr87/KXFBlZ+wSSXnjYgUwlMxZO8xY/D00GDLCE
OhF3Jxtd3y28vI/Mhjcqoaw+rVWML6l9Ar54meKeD3qJAtnE/OZzo/ywL1mjPWLMuShm5HPSJHPJ
nP8hz41ekVYg58N7kYeU7mHBglPARTFB+YaUTvrX2xo/SvQXSlmBdPgA0rbDP6TrlY9haqUH1rhb
Pk9S17kjFvGwkG2VUMcSjC+epT2yJJRMqTKAUHC7w/YSxHVDUuaueG/85MvuC4xZ405Ze7U1f25K
SZxh81LyXHsJ15arY0wzruTYhxJkdKvWybyBDc/V0W0dbnqSQ/eGFM2sJnfaVZg0rWp7RfBLZ3i0
BNNc5VF825o6VvR9MwZ2PaEFzfx8vVcdLJ9n2y81UHGCoCSRZ7uG9obrHAacb0rXpTB+2ZXM0+fZ
4n4aD/iaqyy+yku1oqckamn8lVeDQkCiks275KAmmKrtDCBtmumgM83mb96XuwnWBSUNT06i/giB
8fwdT7DxBN+y4lwDAR967KTq4xSzQNnvqfKkV2gxkSrG2ThXx7GTmvpHm0LN2o35eSdL60L5kh/p
VF8EkR4ozsIXfBSUWkV/ODVqwWddUrXxKsepw63vqzakGWSu+gVulBazF35RjmL/E7Hgs0h9ZVel
vfIfVcn83wV/UygF2eI+U16O6hvtF8YsuOImt8E3eKNFEn2G5E3aAMHN4fs6wmnje3CDlUk9W9m+
H7yE6IUV7CAW9+PxB56QzTjpmyBcJGi82XW6OV1n75uRHaPpP4s6GuSJeVLAYDOM8KVAKE8woOJu
OBBHuHSikqa1ypkLPWd7+ItS8sWJBMd0z5B8+d5KBbehlPzF7whTVjVTFdwPS2t6ByhKkFftVY4i
UORQq/Y0jr0q8MQsEibM5ksubS8que6XpDDqiKsEZ5C+J+q5ky3jpAhe403vZDUnunXdP2MLOe+i
Zzb/MNxKcHwuvZtERriHC+7CibLMogmhYZzJe390VVYB5aK4xBkX/CPFWhRurXpVnH1eRgCQppOB
BzMfhUkwIGjEu507XhESARUe2QjBuw9/I0RbmWvQ7oG/DC7Nr26YbmG8fmGgLcXu7sNt0kTjtxch
0bEexrs7fs9DvLVCneckCEEGN68crpEZlrT4O7cz3bdsaMAtIJzuw4NqJ8JSad8namQzj3v2AJmd
UX7e+EvTl1bfiPnJUGeWNg4bvRdgqo2W5ucl0bg4JKE7yMgSzT6x6tHKpWMaNpQCtJ6Ziyn4fhO5
kaNjbXXsOhqcBEwDaNg/Ya7mFBD2tzYtKs45kgEnhkVWHp9nJWYaUIGsLFP1ltT0Wh6s+22iYGMR
hBN2Y5s2VsHa/00sHzGxpGH7vH3bkZdd9Jyw0wRBRqmKnQQ4mhfw85KELEBw05ANAqgEwqO3AFn7
LQncyxjeYcjZukatRNipgLEwlK+fkmsN+iyNn1rwWHv0oDHfdlRf9pdppiragx/zN09udYzTr6jH
mamab4RGMYDX+9kkkzu3gfSeLSGu5fq4e58BEw4m7OC3R9lsx1feDYsThkAtL352q/ICnYWMQy0L
M0Snbrj/x/yjRyHv6nvXskbub+gyGYOna3Ra48LF4DsiR0QUmshmg2kAyl0xq8SMc4ny3dWK+AR4
UeJcBLfqpCa2GDE8wiaKlLK4c8Rx3QB4ue1kHffG+kMRh1WCTPPpl+BqEl4Y4/bjLb4/KuzmfqiJ
y7TZfw8W/AztZiR/DxFhLIX0H5cJmdGiNs55zkcbNtyWBDklB0+22+NvsUW3Xh9KXI4NWUvGKwf7
71U76EVEZAgW726b1v+CZAYuBhxpGj/VmraFpC0jtDtLIgkh1yVus0/BVMoLBz1Le5rDyAhmpyFk
Ib4cbqBdajkBm40D70bKpbhvcXHj+8VIGNM/04459Yq40vMlvlISAwPuyHdAqmsWBiX5ojNtK68W
iOao5a/ydZTnJDMSHI7YOx23F6RZDe0k0uUFd4ggsterwDKF7VyBBlg61bYQQTZQqYij+ywut8Zm
zUYjuZ1oZBAvpAqhhnUv2TsbNim5qkhw6810jIuWlOAWH/uY9asDHpzcGR8+XstDdqgs3bazCyW/
cg3hjV7VCIUqWW3fsp4LUVOh8hWE0d0ceiZDBnhLj2jqClolIqsF+MzBLwypTW0zR2d5YuDHoxGt
s6jiCwsnww5eVSR2GVTF4PwQr9nEgEIEu3VVvoRKoHzhtCGKkDTk/g4bNjMn5ubl0igGdTVtD2hj
H4ADyUEC10O18BWx9Zp6gTangAKhwO1j/gpQtxJ7KhBDr/AkbUaqZrcONyhaqeYBaLuK87d4B7vL
XhleMVZ/Jom365e5FtKOsE8YP8wujGAl0cbtqz9KoAV1bV7w1MKQqnh/z7TM3mY0+PFG+mPtOCPN
u/wPuPm1P0srlgq5fnqQ7mOI2Dp4wE9hje2uc/IYJl8nl1Gv93HHbqQ7hwkQyiv45AkuK/O2RSNT
Zyrd0gkPCsSeAJtoqhpNeY18YpSS8FNVewi1WySSH7kEGxJd5F2N0eaWXUue8nmAzW1+Gsm0+Sz8
McqOsTQeEH7x2KC94aRVNW5wLoTtqWZgIwmq3kLbaUj8WZg9WhHCl5IpMYBv3y5GoGoGCy1Ghtbf
7/lnn67wx8S+YXoYms4M3DA83kZXgCNaK1HNcyDP5EmSLZD/1qrd+Eo82a5isVw2+tCbtlTWNZjO
7gb3eOFLJE27aJyIBuKlFJW3mu4ilnOeGeGEAVuemejJ+Mc5NzYaAw282jxbB9fRjQRlyzTBYWlA
bJcSodd/U9oaVIJMlIWHFkwrF9RP+y0daP/nmBxbJep6zLDDr7pyYOQNSdcrp+gzIQpJ4ivfMoMe
z/TTu0tCht5ZmsPbfZPRAW2nWd1z1G3voT+o8/NBsTyRi1R7AEDKYmhrp3dFgL6bLLnPxLGAquoi
G1drDwiXgivvltCQZ4mdJ4ApgDwJIVv9AOrnki8OtNQBEyi7G9wikXXpgdfnq0MSbgGLgHRn8Uao
coF5qyPeKKT+kziuu6S1morj7qvuTsAzCaIuJis7GnW4gm3riYo87oPwPt9Wkfqpe/a5ya+UaY2l
Y+4bD+kpWJOCjWPFIuK8B6DUVfkpzVsbraqJvGJl/tZVr3/2XbdR2l2C0CqN09ICKw3shDfld0wn
ObGZi/M1WSqMNfMHB6AaGQoxL1SsWHZ1yKcgZhcBhrUV/K0huF8Jk5JwO20WSxJ8GXj6cypbh6aa
xnhU48YUy2IzQnioCWWkAEFO8KfRGMI6uURPSufHPTsUFmn2DbFVB9B8jHj3mkuLQbS9VU1EKsfY
7+s/cOQXJSmm/9HcFJksoPamEqbD/GYJ5lXzTbd+GnRvdUyI92cXIg4YEPjV8sPZV8csn03KC7DW
APIbCr/o5B6I0IRzqPMFmreSJKKfs4MmmHEJTplHGmCZ+OETCeTEIkMP85CRgdumQoP711YnnkeD
4AzMUahKkw0XSc24KHSoh0SoKOzlo48cZs7y8LgzgvOs6ZJvs4hUv4r25kpdUDvYIYyIBw/ywxFy
JNaa/CsYsm8d9AChgGcWqAVbrBjNcn1+tbanzsLxsurOyhRh6boUt7EzHRRNNMoclnvK6l0sJDcS
j5MeAmjxkLhvT1TkOjJeSiZbTuwXKQE6sKRUmD8NtmnnIybJbuN1qpd8P9ioP4Q4CMehSLHma56g
OlUoliAkcuW1QPzjzkexE6QX6/HdgmexQk3jtMeW4TWWG+4pOMjHvOrV4PZrV4InBl52p6yzM4PT
N2bfT6MmbXF5afHskiBnv0s7BB9oyIl4hKbygU8gObysBt87LUPMflB20cvauNnDX55WS2q0dL3d
jGWAiyO9tnCa8ZKYvn3XtRCK4a30+Nx99DL5K6jrDMvceEujxQ3ZdhK5U+oTwzkJVdTAmN7UAE4v
9KvvMYs7BO5HFLp/QcWGtw+FGN/qiaDGScBZCOaYuDEezSlVFeT+IqfO6DkG74yPyPFO+gk3f2kC
O4Mm39Z+UiYcgunU6TjY3t2ITz9aINrL3YsNgyo649uOmI9TnQHwNAuKCsYik4swrMtk78O57I9r
fRJosqd85ZYjrb7FYBTic2HTJfBxPw+b116F0Y8m4LgNbJLYhPKscBVxSSzFrr2eytE1kogDuxKR
A6ou2ty1FTEJv2u6SRWHutv1uaUiy1K4HuIt+E1xzhA/yKwi+IBqMDTh6csYm4yMEHgVuOZ3xeu1
wcyuX0EdCt1XwmfxFQTD5820t7cckS0xTtV482RUXIKySpZoNYksrFFH9BUPBy3/YgY1G17iro4c
2mOigOsDMBoUrt2qVpwG5iUlKHcqHlTmqeiGdaCLcHS5bRLzuXx6HpIQ0diyBd9Xl84hCjPgDfvg
wd2obZ3o1cUOYExS8nMTih/q7CUdbPIE6mcbSTOSSC7ylpbwsakV5HR9xnQnl+wjDjE4fXMYd8Il
qAh/zlkfqn+CLlSZAtQnpMAExqppPS4inv5I2TC5TwUgHLEtjoZLKqH/VqGIXML0SsGQAJ62Hnb/
AIi0TooLL7nGcqepsOLzzQnVoLr/guStY8mwus03AJhdZ5EZoXRISC/mJZixjFonmr2ZXkCd5cVD
Ua2H47eICRJVPpAba0vYHHaKOhp4hS81ONKrApUc4rrd5d6xdN+cF8xPCw/6mrmOPb4xz12gQ902
IcA5RvZlLbMnYrZV12/3CsVSBB+jfvpWszwSAN5psdTD3Pek7BxMk3pxRxU2U0f9y1OcUtmk3rEo
bzQMIKPFXZ4gWqW8qXYB1qJ8D0fTB+gBPJ6X8htreVNpDHzzg7ChVjADSEozD5ixvO7oYTES5vjH
LZJRxWAR7is2WrBy1XQwnfDY8K8Z4zt1EVSS9IlpeNQRYe7HrXqprBLMKMSQbR2m4Vh4xdJaoRVn
v8FWDZNmKRlAO77oVgOVsG+OOwUHkXvasmmUC4R4pZU2jhXQPldO8YHnkmrmmLmLR4TZ1+kGH3bv
Q15IyXA74X7we2YET3ZNZ0t2rs+SgL3QUdIfgJJQ328YmtFlVRhO2RP8emKFlgLBnzLAYKz/qLMl
9XiYwHJnd93JZVyDe9vckBj/zfPmUmvrSF65V88bvCEYG4mkusdBOf+zCutYFIxuP6ppQMqMAas3
5H7aLByxxxZTIbTMid+QlkZuuVdyM+aKROmbnmbMWphq7/zvEU0JSaRCdgPzsrrk+e3h7UqkPf+Z
uBOUnbjh71ADVRsBdwCZFPtW8yQtrBYvkfqrzumwIywwICU+IbwI8sKgSBYqXnUkT3iFd3ORsN42
gMuuxXtbcFEdA0wl9vF9jUR7Fuabh8p/B5HxR3SFk9/NPE0lqoJij+LU3bDAImESFzIY/JoobpGR
B6vP6fYF9OzNR9JlMXofLxf7WrQKe5AedNGeA8hlfcR8odwR/qZqQuiDI4j6d3hSeQ8nr+y2x/ae
dELJvJiQltH1DWACjHdUdrJKUnaVru3M58yJXNMh7iHonuhDV/M9A/WhUhADhEqp1jlrhS1Cr3LA
Lt744ACP691kKvdmCk6qCDCb0C4UUnXsaL1KXV89BVYOIW82fefZG1Z5YcdZppvXS+6TWDsg1HV0
ZbzTwxSHyjWIDrA2/j9EpwmEbbo0QES7gdhUkwrqAp0FcXxmNK6+uHg30Q/GRoBqi2FTbClZW/Cw
SWqEJlf14Inm9a09MNBx3+0+/Mp0MS/DoKOHexeZzj8WO8q/PtUa+Gj9uZAWqXKcTV4U/o1BSjTi
ylX97HZvGcrOsaofSSwQHpA91eRcLSaZxAuw7k+z0afYRC8RVGuyyNfzRRW4gihqpoFVqi/EDyxA
Kl+j44X5Ayyt/uR2GAfn3lEJIk5igJ924d5PzuM6yN3ZtQeObaJI9InpMlX6hveJvvF6Off9m6RN
t8uc57EOaVmSqSgWte7Bluw87NBz/P0q89HZDqSs/1ogxuZfmcsB/mPLJZ9+VmeWnCFvcqIX0+Wv
IrCTwqWeHyeXV9pegU2PwdLPKviQgIDuEEXJWcKt+JLhDJcqjXSubPrApDjMKYsprNNN88oNZG4W
vXLmcN1NE7gcIdIL5y0Xy2GRiOGEqDlPk2wXrqjaha29KYyIExmuz3aaOeUNguRyfyLxslM4Lbru
0VkvCIYVSUIgc3YhrVQjAJ6Oj19KeePqM0pRCV7UVqcr7YC8dAWs/o6thqW7LYCnqL5qENRc7ExL
nVUkyEOT53ovDMR0fczJJhihKQ3ht96HankKCOBJFBA/Pug+BxkuO2xegARvngzu5+Uc1mZbQdJD
AUk1mqJsM/6HBhzAu/4Fc2zQ3Mlio1qaNaHP8/WKQhLLV9SZ2cEWvBT0GlTU1hlI/Ccv8EXqsb5z
DfWRO6d7+S/RE/NtWEa1CMnq6J+fqdUVcrXa/DFfMuIIzrcxdKB1VOad8xOBOLg12C5sFFgdffFh
GUaUDrxCnrUcORqy4Fdlfrvuo2ZliE/vBy0D3MS6yox3P6OsnDq4yJXXtKVnx+Zho42OQRK0kLRo
BkbZDS0TB3Oe0Et0xaKt4bSutY0sYSNkmDWRlz36SizfaQ/SYf+10SiYJx1PW5zHn2U1iM+CUhVI
1ev3CpEW2aTrAZjfT/Suumgf1XBSTvht24+rpXizeyIm9yf8OaqHCckGk+MdqHMj7cPkQeKAVrtQ
WkpzL8srWTcIJMT8SvNvYOVYnfn1nLm5qnZwMdR/oDEXvPAqu9YkwAOWJasUOobsvUFeinrgYMxd
eoPvpsyu41SGxZjE1j+xiKdz4s+N1xpBOQp0h5EFI222JOXgm1oFArsQS0KlSOxA2RBkrsn8xvbE
CgzuQR8X+UKwbGSYqWTMeP4yOVaKiBCqoIEDvSwWOLex9ZJ/xJCDmyjbfs46z41hhhuj1mmCOr2j
9ioW7ORwKJSHILsIKqtAyJ2vdmIjh/+RA2ehb5R5xFE2jAsH0HPVj3/ZJsG/gaUN8WyTH4sOstg+
JmCEKKkuT4VmJhirS/X6FasijTexqnJfTt/Mi3eY3W1BLEylVmp81u2PC6E1xmu8Tv0kzb3t4Vyb
DHOSVniMPlcJqE6uc+Q1B4TjlYnLoFW7WvonTpe1NzDANZY/AdkvrCjdH01ir1Mi16NoXi0ts4gs
anFckilFH0HYRsJDP26DHXIELJkju+U/db5DXu24QoL2K4wJQomlVR5JDj9RDKtzZywd5WgPpvBV
2+swCy4W/FEHwPmPHJJ167AQxlF80hlb4Chv3mDfRO05nNaK3FsdfnZzxJSgQi7VrH5Pvj7dNAyd
qm6i9Lxi9ESNHH2do2XkdmsS08ELhnWj/H847XCm3IxYAL8/h2pVJbDCXPsm6HC2+26hH4QCcngT
mYl+EJF/ewLIP2CkWryc9DD0NiD1Ivf98Yh7iqhVwmY0/CUbQgqFgvnGu9Lvm+QwFtWBriAbPUKv
isI3k2f7prO8hdsnYXeDGTDOqsVrHJRitjtxJVnJ7gTZIUShSxc2PXHjwgOEwI6IXgPECwhe2N0b
bR3sUBh5jL9llAqXI0ZS9IpowkwJy1AZun6j+/ezQwSn01p5hBAIPsbjJ/mkAupE0+cCA2pxv1uT
ipLiGBWC2klLrQ9iHx/DnZFn1kiDJW/XNVRW2gU33uNGZ3wpuR5hmDgSnQ1K/AbtffGwJ+s4vMdH
O+R8S8GOyvqwyk2qzAMLlVVvHR7CYfw8LA402RmpM4zDVQOMlfhlitRf2bX4PJQlazrZXZZKwhi8
HdG01smMMVJ8AObLFdwullTGhgbom3Fe9y6SjIsOnwIhu0mpuBnWBfsay2c9WjQShsg5OKAer3/F
NDjPNVPpySlplhhgrkCQ+uGSs4DeEjxbPZ1xFj53sSNUPwsN/xi76TrZzn30QcBf0Gpx88Zbh0M+
9Y7HWcjkyz72cbDDHykJW4mgaAzb7gxbjbzLdLcorpg6lBtmbt4yqkqCsziGE8bM41+pnDGMgv5q
DdbxeV24Thv5oixLpzMBFv9HxlSEKsU7vu4iibvXReyr1psqKsVU2eWrSjzZIBvA5eg2A3b5QJNu
9lOe+W6fHQe5cIKByFpM2A==
`protect end_protected

