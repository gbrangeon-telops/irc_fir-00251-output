

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
CmScm1EG7+yOvSHJHM5cOhdqnLzZOcepWxY9DkMOyN4kLbgbdLuAH/l5P4gSPyg81gBN3kT+DB4u
PBXNo4263w==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
fwqNpFcMm3h5oYp0iLLBA7jw3Gfbtf9OYXqaNYQK5M/u6ozJ7zqm8z/7Gi9eaTLXS/9fpHpwK0LS
QxC2diEfybnFW6aKTP/iU4AM0T8Jfwg1fYYXa19VRgeHNuXnOnQbGrbwOzyL+M1AE6VgNshYAcke
HFUgdv42HBSaLBuVCGQ=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
D3xIUFHSYN/tuU6xykyZi+w6uytCi8PG1RRIohuMCP7mdmezS82HpITZGe26wOIBAYGliyfJF+bm
//Xu42+HAg7awD4lB8/Gfse7Vws0SwmUepHhRYxtuQx+Hau6aq1uL1eE+GMEUXgxZ2vOXH0ipYrS
hLEg3TtjTbccTVimoRhbMQB8xVTXKgd1xaluMo7+0fNF3EBfFdhrX7VNbbmxpV636ALP/wC6VRmP
XNe5xXQjiv3FP3uE/Bt2VYm+z78C9QX2joRNZHnjI1wlv+JUs+OBnQx0uieg97dZpGTJDWS/ROJD
yUMDQnx8oeo5Aftp86QvBAbfaqE5X6J2q/lamw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
WD1VRz/pLvBXDYk7fWsqqk9E+EKCxbcP63KaJV1ph2old7nkwo7SBQkXHtT+4KqXUeTJT6DxPa8j
tS5RCAcDnWldx37xHa9SUujjT7DruuKAJejsjhxtSfv6A/nEW4C6nOkCH10rAuqtBTv7SUZEElTR
EXiyr/yJfBZig+juuEc=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
TO3nxTWXykAydBE8oLE1lWHpTk01Db/e9HeGVQPfEOiTpRxWensjccZLTO1P6wLTocrobkWdnzeG
BxBt7prIiPwnDDfhHMe/xea/ckp4CqeBr0GVOckjbocHEF60X3dEzewbdNfFWYT0uATcWRkKB+5o
X3VNEsL1+rzFW3yXd3oxwxLZl2hrAEzHGv2AAZZgDP43u0eLOoQsuloFBUh5XzvTCc38IZkfTB7l
fBrAnLiMxoJyYNeps3ny9evx3MIX3RbK+6dmn9Aviq++SNxcoN8Y4/1btHsL6F9ez079jTeANSEU
ZvBBfKlGq2n/FXU3NGHAnGxirPn//Y4kyfC2Kg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 10960)
`protect data_block
9ToTLhba2yaS6DUGetuZn84H7BoRj2ZtgkPfHjH/un8ujin3dWMPu58Y3mpPtx6Z5+C/iVd1ivSN
iNkAfzk9EKNLemH2pqQcy4zcdSJpGUx5ccoXt7Kels5Jvj6HXkw94/Epx+T+xtIATBk64J1AXU1y
3HmQjLofuiVBBgf7Roy0gPEk1LQAZclieEt30dgbUdB0+R4cHgjbdxXkx6qmyBKquOti6Xtmqkfw
rZjVs7oswhZDH3jnYVCjRsyHzfE225UeEWG2XBstUFf4SoADEkb2KDlauEMonbtleJsZaIRU9JYD
sCK/v1+67/hFzaEyAwgY6PrwmelpIvHJD6BVLpqnaQuPpD8qp/9SjcRBD2MKNVnWImwF0V9jeeXn
hBDMMyZpbvhzGCGOA1tfYvPmXGmnC7Ee2mysKOpHUXms2VrHbb75gKwV0Dpx1v75+MZH9BAOyCzg
HAqoBVL929axT89mticHT3ywoMubwHHjF+8DI1m1nAYK/FWVg7xpXdhgg+Vn2eg2/QeVBmbVQyb7
22Vhyw9abPd/E39uuftKXpsb2XiWALdXCRmG/8+z19poBw90P3/czX9qpB69yUFbSgTmD79x43ie
G/75r/bWtnCmQOqKGE2d/4mkNrm3p4umwlmWkjZ92Dn6hPrUct8TzquAGjS8udsikpELvRmrA0rV
Pe7u/A4bStnayivc6xCrx355BRQQ7x+MR2YkTkAGp6Bgi/Yhx43yXArwSWJXxy6Ea05SDELzh9L2
YcnX0XBngfb+heuYcE/w1kcYyC4L76EwdoclRsIfeH4F+OCeUtMJTYf35FbSShLlq94aUhNzQ/KT
twTVJxKjqg/nWVhqML9NmSdu6jVz5st4UGfWztCDVp31CiwEQ1aMudsdYbnsrVLZdxnabXKz0bxQ
p5jtJM6as/wp/A6QcMojwNLMMQDGCqH1rY68i7N2lT+oDEJfriVgR/oHZr76FrBX23J6y8+4ChA4
He15ziyDznKTAfutFpmGMA3p2/o+ZGm+yJgg+X/KMNqpGKZBYg0wjeMONvk5jzt2zqCAaXil1UuG
n4bJ5SilCJvMVqRp6F0dvppbJOakeCjvge32MCwuPwkxVpIGZDXYWJJxHaryR83MLwpdsnFv1YPP
qYoslnoJNVHAGu1+JKISWoAwLKKjigLm/THsmdniSglihFpH0Rp1mOViJcx/GUoeGQoyqoHnULf3
MhokPwfrrnqVAIhK8z8gpF+PpbPg0eGLZALygczE0qEcVSt7uBwgpdRTarhTpXTLate9x0ybVzKW
dFum0EzB1heNtlJA+dbm8smFruTzm2+X/2VgMEESEmzv1M7dJ84LpJ6VxkUdMMi8LiIkaH0+RQq3
d93vu+HU7ZRP+zFW/4wGj2+s9cewYsDf6Jbc+5wTtztn9OWMe7/dsLxjEMq/C0sToYoVujqCbE54
wjtAJzAClAMiGDqQTK/vwkzmuP4TigEl1/vFUauwCYhXpyuLau0Cxc1C522GycOVnsyA2mO6wuy7
8bt76I8h+k1/HwplASgQMa6b6JEFQoLFYKCvRAuwr4x5bclxZI1Q4063lcouw+rTMsQVrwoZRrxZ
PsGoSpoln6nfQ4+fPMtjYfo7c7Wx3ObOvy8mfpFUZiqMrQXQvOKL+2/UOxvAnBUjxrrNVpL7GK+3
2oxbrXws+6VPHC4P6+CL4dIZ3qCXXjckgpsf7u4ko1ryeeSHlWvhZAmtu8duMYOS3KJTb6Ah1Wia
BVF0S33Zv/y59exB4D3hntZQD8gEzLyhKi+Amj4eHG6H34fsEaitoSer57TKWZjOUKrmc84PPgiE
YqmmcQ1GnfZDr6ETwQ8CUzZgfm+q0B8LhLCjCX7FEx7+gfkuuoZMM2jJRIOYIXz+BXd1QQoRBHJK
m+Srp7aDsEqG9POCz3aqvzw81RpBSLEzHq6l7GuKH3LiWYzR//O4q1EAbZQqod+IOtqM2nhR/9pk
sxJaIVd0QOAEgAEdcpdQ72YsFFG6/L7r+7xAOjr0gtV4K74ZhdYOJMkCj9mxEJ3IZYReMKLkUptj
gfr7OAxN9HplMaZBhCtd79PxUbcMu3DY2ZBiVsSLILx4CocKtLtB729IlP1aHJBxjzIosr8KSNmj
yrslG+ABIdbf0JpAhVzxkMpVcsrYmZY7i9LT7gWZZi83wJstMILerAJ9+1HJ7p7jeWi6+m4MVWx1
1oMFVgRWR/irBPYvKkkAh29JupGU5iMe5qio+BNY9RgbjCYTnqMP7ZbHRMApOEfvSzcrnkRtks26
ZgX3yVi1S8wlWiDOyXDaacCW+TnXJU0slVjLju+RBiw063pb8erpUPmjqxvbaBXWxBhlgKWTogfS
Us5U9egJJySTc8/LuwUrevDV8AMfwgyg19LBp5vBPq9LC4rQ1aMzFCXU/XjUAHl1S7CWp6RIZKhZ
C5yzjdZKLhkKhOqhSmrCbU+1ApeLmOMxWnlPHMSFxbVyqZoUk+HNIxdsMr5jCKsFrRwfB0mY87kb
LTJfRHJHeTV2lPX0xu5JUYae7ACDmGPBrEZgPNR9GdWfxkNYPq0BTccS+Ef25HBdO57JrPptwNnv
zju8D0/dxBfTjUDo9QhZ20SFo7OaxUBFT8IZqIdvhg3dDCLfC1HYLbE/c/ha2vJerCStXCsmsxA2
BtcFq83QI+vh4es+G1za4yprSUVlZpp2aIM/qQSZZldrWm/k5u+OzaU0mBZoKaP4TKj51P8wX9fe
a7c0YvkkcwCmelbrtpzYeVZ6qsHjG38kB7pMuqofdMrpwddZuFTMRxCvJu86FK1DJOcKtkvKU/XF
rb3Kndok+em4eps0l9mdH6O99djM7f0qpPhnS2IWKvIK/xthyTUKprFl0mv16aZL1t2J8WTg3rIe
M/BOn2vmxWBxcRZ2s7/tbzAp2OpITQTxWeFWRQ0WUk2/NLv6jv1vaBay5td79+GD147nKIVgQQmC
TBf8lsNKW/n2p1RLZL0kn4k9gcBfnP2raW1ww3JD66pjNWmk5Cc0XBZz5MKVhAsFprhWGLnSbaW/
zhTGLcdKEtHE7dOfOaV/5RH8JJ5WQjd8PFibwPgwc8BuKHQoRtrJUP9f9DKDfWomoRmRIeJv35T6
oJQUse1wX3B7fKaz3UWsJtPT53QvfWmMadLi0u5ZLRm+sTynUm+CSRJObrkl9NU65wzQztbpgK5i
cN8g4WVwTvIM+MSAEgfoai1yJhpDgXyMRbKxGmFbMagejB6bOzueAofpuvRRcDyDXdqBpoml5Fl/
8FeqcujwY5hA4x3d6YE6WgnMcQDI9f7odGCaVUNxJ0shV/ufCir7oc8/pdQFYTHfXyApHhoYSIi6
2PfGVOJ2MPw7SpMSnYUqsNBZmSo62xIjyqGQP5RSUS29EF3NctWGien/w3NZfPmawmXRQtCQHugT
bjZENGR5vR9ZhVpQifQWM3m298DM5UyHElgx2FHYmQvreOFxfEV5bXfPQK+/DPCgNgdFCwFNE7l2
2PuG/jJLMI0XtEVA8XC97xEkVowmUb+r/p0kxwA5YS8UAeDNXDsRJasDpM0l4shV0lyzBG48Gx34
fBg90mQZjeIGgbSIAB5bFlFwpqa41d2bUA0EmnBxaH3WhjsylCvn4vfl2+u7Zzp9ZRVKEj5We/oq
Bz1dSndLtmK60vwU/sox8XBr2Fp1GuHqlrCCUgD3apvHupjN4SujCzu2u6tR1yT3dkokPUQYCTgj
XtSI5xGaHU86HW7UV7FoXNK/gYEFo0FCGKta7MV0tlxB+7oplgd0+X+BQZU0pvJXalQh5QzEQRUp
9osllbngNaa0hrm0/XLv9pclEGRWEzQFD8ZF9d5F0IWfTVW2CmRWd7bGpO3Q4LgO8PAVgDlGTgxW
YXHK5xvncK7i8upim5qlXxkOt83ReH6juwZjIcJFbFKEJSDnr4RdT2toere1CTUxjYU0zEBjhEqz
RoeTsrw4wggYI8fHGhEZVNcf1GjnAhwsuJ+tniaEgSwhS+icH+Dt1W/769lUnubbFpRT4/LV687X
hcxyvTIqhRnIVgVmfLkt+nJY1PeZClE8jZgdMI6tpLOuWMf7h9OfJ6A0xIKX0J7OYPFQ7KvwTiSX
arCrD/LWDd9kTMBnPANYDql45o/M0ZACJeBAfimqczBuCZSFL+zY++Cl+CucWRCOSupJoXHi+hV8
AKAbD7EQ66hTKryeetY06akmjkIhMfDnCx609ie2bOnlPtEuHIu4P/njSZN4ZQAF4OAIstrrQ1Cc
UwIniCBsLxudvYT8cEtZGLRK8FqRDmjKicSlGFk/NDAB4dhoNM7cGbOsOb+aCwfmQx8Q2PC72InJ
TqodNDYkBtgaDMjE6/k3yYqIHo4l4VGJoK/SNP5x6+U3pt3UL4vlN85XwLbEftuEhg3iH8YWMADe
kFPVP65rczszFXG5I3DdJlBIXDoQ2ojLGcJiHxEGJ/W5QRpGxvBATm+RgLflIpHwgHOCIFdHO63/
C8rFe2/miNdyTGU/svRh22V2g0wyTV1LsqArjaDXPa0iDPVQg2ufxQPnrEtxlxps1/xAjlEPI9Xi
/eYUmtuW+it4zBmNvBSGPUHAO3qYCHsyXodsUN8iSg2jeXYFkRP3gVjyXgc9HD8ZLiXaERakkN1E
VBKvgNQDIZEik7qx7y15WWmvxEnUT7SBif7yrvmwaQzWdIqFgDGFcS7pvds63l2ZItaSr0obclqM
oAyZs8PdCiOd58Q3LsvM52wQoexBffycrnyr/ufR6bHdpG02msGalQzf/xBgAjp9QqxtdFYxChgE
NO777xmFBkRQwzboD1mytx+EKYMWLlZ+NB2y8Z6dLRfjBSexemPMWnW4jf8eT3IPGwoUcsf764nN
g//5DLg6uMSwL8BCdlLHOWLqNDyCkEKUz7L6fNS5kI56xZcNsp0tdgTAZ7VQD5xa8UUKSKboH2t6
9ANMzYIUOx6WhAZDMkVo+FsEJGaxMsWqRG08/PllcPNDfH+9Q0toI+Wor2nAkrqe9bkB0qKfyQ5e
5hzWDH4amcST0DH9ob782bWtfBa5vNDXnKFLf84SN6tqz8ZMU669aMi2pYVTk2+09H5Yif20sP6q
DUVwXdC7Otl44oaiZh8Q8vMv1TeqZOZATcdpuSdxCSC3Y157p6VuxxoJ7xjIyFG68VZjkQ980Lpv
pHAkcgRhf/Hs2/DsSr1S4QDXG44YvBztVWpX0qTZWRIe7WoLMqI3U2R07r2skyPRXzhYSmi8SHlD
86/wDkvjj7l21PTYXDe1ZicIvqCI7QcGjrY+U6MalRTRKRW7fTN/x8iZQBbSKV1ogYXw+2A4161D
gbNko6Nj+tzm1WDWLHq8r5OLNsJugKJ/Jc87YFeo33GDTW0iYvwmJPNdcMo7cckBbzAC24wvIGnD
O/HmlVJbl77X1jvYLk0HvF/mysMOu9NKk+xFTf3dpZm06VS887todJwYzzXNXmm5LtT8KilaZyq+
5Q3lazMO7GZWjKNVLYvSlhJ3vlDzpFRHVFZq82A7+GG6J8IwclRT+CClVpLBknTTBTYPYjxKuIGG
+dqmB1A/Qb957RB5QnGuHPSg28Pjv5ZxFIhxf91bXmYKNF04rS6vNssheYICLlkq8+MVUgPMhQhe
csJJLWW8qulhbi1ISineXORynl22H3FId3e3OE61qZG3K+6naZ4HVA/4etKtkM0xUyBc/4z++Id6
yttsDYhozxi8Dogf80lRKyhApbQhcspiHcqEoRWfql9W9i1MLsVZJ9aHeQQonyNLGVTHDqm98sL3
LCYlZqwgRI8ZwsasuOYfjKhq6S4jei5NzunKfXb1gurLXN2TrERTNU0R1He/5xILetv38zkO3IIG
uO2+FO+qlqnp+85QaXkqL42nc09L/2oJgO13HlBwU+BIfSVEF0z0mrCgahHJglKP7UvfQ6RH1Z9H
4EyCDR5tmnUVZZDCoQjznGD5toIebC1uCBbYB94a2FycY5O8T4E0EdEzkwQnQD+KkwoDJzbmQRad
1DyOUPaJ2eXcPUQFPiK8TS6FNpBfDI80T+h2nuUPsEyrBjpXJG18MkpjfLNpOpa7jueDjdkxfd7c
POquuP4q6eFG1MX9l7PUeMK0c97RMNA0M8DGdkumu70WdztZiB3nMNuW0hIcQo6eGzqjcHTE+L66
AS/7u2aZowMksRnG2/LHowWwmVZgax5dW900emzQxgTqgu7KQ3D66DvkunL2zcbj4/lf5HEmdXm5
ey0jrjUcdmLZcvQxQ3ygPCGalRK5yEKql0bW2GBe9E4GyBnxiD+rWkJ4UoH3WcEdM8t4O+kRtUbU
z5MeJWibf68mH3zw/DFJZdAQaFA3jmfnYnnC+fQBXMH7YzrxW7ht9GNMTbPobecG8z0FmaBO4u3m
B8eZm0sWn5qKMP1FEKgGRzZkHy+feETU8Fk/sJqGEzBxM1n0DF32DmTx/3MyM4JupepPcQfCW6uu
kZfdVWxsM87VS5gMHk+nlJzruG28pFRStkbG4SXsLIF2dxhOKQlVemeN3vaE2SRx/JfOattTr3YV
L97iTSSwv0fSymBbkF6shRwr+McN/5dDOCZTEpj0x2C31yxdEt1K24KBpgIY0HTL/Se2oMZOVZba
2beUyRocPbSn0imo/851Y7WnKwz/ZWm5Ii8TWAF5oFT0Gm+OISf79Q+u5U0KuqpMXkiozNDCOmti
A6CaMBgZws87mx2RNmy/Rm8F0Brcm/Lek1JDnLgWmLJbYR37DZulzUbcAruJVEVL95bvHfHCthrH
DLNndiJP1InmdKDWH/v138weVtSlRkvVBMLOKr52oka1BH4PaGlNc8DSwgLMzhSWOvs/1TjSnhoG
a9Io8IU+9Gt3LtkArk8n/OEooQTHhVUS0wSka5jrxI4Z70qCUJo2ynILHyMGbtE/Df1u7YjrkNah
HQN8pBShHvLC8n++XljxQgPbSIEz2zJwFFxpC/jS/pRKZwQC/GMtodQyozXPA4RXgtHQilNxIdfr
Q5tMBUsLiT57bu/C9vLpV9eRXVDj7jm9em5/uj/3wvzi+Ref0pdGTDYAAKFldD43QUeCoksTZcDx
NcV5bVaqvQcaxfs5RT9R03KyO0GAW5Ofnm/pBX1ymlP9i8t8ObJZpAICuepD05z4UTIWrIhvPf2V
T2nyh/rccAd2+kZY3diXU1DJicYS7ECdPCJEtZEczJvkPnC4DmCnuvjIzZaxim9oZj7SmAo46zG4
hgbZK3op0x8KAp7LTq/EZzoDLihhnIbqLOAfI0AWmdei8ENi1lqTNfZYqMhU3JR+rNUf16Q8Py9U
HWawec5cB+SXkgoC7FozyC7I4Sq6irmSXBF37jY0zRfSzYlCFZ+1xqHxfabUW95zAvoC8+fETKxd
CpnqtWd/39Z1zshVKvy9ZiWzq4IkBYb54/hIdBOw22ZwnJpq2g4JffhTL3WVIIDsUfTGKvRPtquG
8LaJLUQ7nmZ08pt+pFhjxgASftS/Cf0V8sAUeHUP61isHI8XfjwqQt42jhhdQnod/JDXmljb8Hga
h42o2IKA6pQIEZrEG+3geLAJ/IOp4QtoR6Wb2sdet0DcFN3intFev+UikUbyAOVd1w4fpzbJKHDI
FKqrqHhYZW/cyQyC9iVwByc4aLamMPQf+1sFgl1JhUvu8tB0ZK0fB05N9toPrZatAeVwn2ibE+wO
qZcHKtvLYUi8ECYv5f8TqmlK4AznUIEVFEU68Eu1zlnhqsAIu6f0ClDYy9esvDngdutEWCQoi+KF
nenBMUKTa6u91NQ87y9rH0s8RmlTdh7bwHAT8P2KqOttgFWJiAvp4kd45xgfrT9xHB3qyA3KgV9G
fJQ3f2Fz7BQ8Iq37r3CZJXMVgIjqFW+0bOWvS1ukgNx5f7R02aT3E0aApMOheBWxvYM6CmTOHAD9
z4bI8TXrbiZ1UJ/oMvev2/eas51dSNESHM9X6klziE2Ks789Mn1Tjrf2eKBM3zkD/a9UXF6j/Kkr
0Iv0gvbRVakoadQq6JpQY5atzfRxft6zrC7csS3NrQp0UlfGSyWggijB5CK7bXGZl+ktEoqscCsJ
52zFggetOlXodiQ5G9kpNCGXSOlRZYkzW8Qx9/R/UjzzJv+HrpQScYHGdejcEVN9kFLz8YWx/x6o
5NE8RcSbFl+1PNQ2iedUwluPPZyexci8b8hz/dYlU4oB1+3ezLfzTd+tWU/vC0j8rvhTUiPxluyE
IMIbAl9QezWdf1wrvioixdIEUdNXEeRCSpHWGyKgYwfgh2I10J3FVu5GkWzYK8hxFHu6Won6yfB+
6AKIlv1VIkrDnJjy3MxMrmPib5Vx2Y89v/BH6dwP3wpVM08rgFFW5G2k3jZSws0woSBUbeUDSbUe
LPFb4A1N6IXmUr6AOVBgfkizu/o3TcOyt49XX8o2H3tWKg3sDhkKG6D9y3seUirOsewS+v80YWFJ
o17ocBpZZoW61LefRLtJcfiyYyGIZUYxHaisMSXIHi4YnZJwJwyfmozIFVffrLy0kxTO47DvVazl
yeyrzT1YTMo71jCoaUp00ox6AaOzYs4tB2VE0e+EsV7pM7jj0ucWDfQ2KfE3KP20yC3SKRNJopyE
18mojS8/0SepkQaUtL9+T9pxmtqjC+yqVnbvqb95P0bFlIEP9uh1gcSee+p0eWMwn5nTCnyQL/3S
jLoZDlRniaQQCtoaI9oaCI0mAaz1+b4daNGi6A1XpXDphIHcbUwcApvTDmyxtSBaCtkgqNL+LMCD
BSvnRDzw8LrhrMsFAXniI288+PCC2i1H4vYnbmu+/Z7AV4KT3Ey012zZ2zZ9c++dll81xHGXM91o
yxVHJnv2fUTym7AAeb7biEw3LQ4R1EN+VW8GC2T75OE1g5TsaxjhW514oO7dzOB6M2AsMrTx1TDE
XyKG5OPvyUXlDIwsYLcDyJ+1rDxJDioZv1Tnm+3CV9VgsblSgkwD5oUX1xEYAD+zNEhWXJC+9Dnn
mPI3sZXqmETGTdMdmqzIvKWE+WYVdtpSDFXKcXWk6gaHDwdxkolFUVBGwc8EW1MJ9IawtwwYivUU
YsFHZvO2VDJIe8pllAJXgEQzvJu3qwRLpg7mD9yd9zef7ZWs8qKem4e2E9tjOa1E47FJdt+ngG9T
jnIDQlGcn1CH2Z0KKm5EshvBM1SUOjqPtYFkEaLdwbnsTm3pkRR2oJp6NJFBSxWbe9b4SDkS8aEs
DvMNSJES69thX0cfU2nIRw1dyNGEqt6nMVvNWAOYoE+ElS74l0Lfd1QtXmBWxE8NWCToS/3yqffs
dzw+RSPs88DpHoE1n8ggI71VCi4N3BR8XdOcLAwes6BP1P1ZcFKzsmdbOgEh8viJ5Y6d0qEln0QE
F6ozNWNZsVK92cnt/U2zwjz+GjY6oEdSaKFw4gzKBUKdwqHlmdDtKsN6pOq0yEoDDyE1j+H/ZMPS
cqfaSGpLoN+f4YYtafvvfcxSO85k3JLW2xrziwWUA4tTKmNYb+Ih5pClIcT8NJIzmYlf/q0U01r9
nlwCTarGQc40zOvdyzXiz/d/Wi1tPTQqKeNul93+7+OH2qVv1bSiKDy+RT1Q/Eo7tXF3PHxzvJkT
Pwtf2GsHREu6HrwsarZrnsaNbTKVn1J3aTZRwYhfCHvH4aAKG7cXiEZXy0L1m8/PFseKYRofwdce
Soet078jd3bx5si23xRVQR0GG4n+uOOJYU5bLUjPQ+QJdWz0EEBZGX8R1eFz1rp2zV1edohKpvN0
OUtnZNGOLC8bXzfMcnE9eDhi/xBYJ8I6cLTUGrsDpYkGGz570AfxEYuETLGk4i7JFDiM5D7WEB4w
QV7qQ7pl/VrAfal/hFH6+4YeyIN0buZymYF/f/qf284k6xTAFmLrwJ9jCU/5MTKdBeeaoNKjnIwS
Ki/Vp37AOEjSNsuQuQ725NfRir3dkUkqW3KPQr9jhIwW+NFCyIa1reyISeeYG2DTQIuNBydpIEVC
2KDKyJT/nlPiTWhhXDda16kqwqNF6k5o8sP+SjU0stZNRaTgA84dQ7dLhJCfkwqZKCL0fiTqxiVa
E07enKWjh2eF5bUhfiUXTEvlDV0uxXJGFCfVC3KlSu1Dig/E/JtBrS7ezGoqgeJ4WE/4GP07VEzJ
LsC0uxSRsV1s2n+skieNvMePiO+vVfS+5JfmNaRrTIKd/ubs9mJZcD7xk3v3otQ0V4VpPkepGM+k
QAs1EeunjS1eu8dfQ27yHOA9G55SP5/c2VA8ka/t9dZXWEOngGwolZEcjQmadHC93jjNP0CB5Hkc
WyvbGtZmNIRIupuY307g3eyfztPXDK+lwDZ63oeSeXHbvK2D7YFKTHWrF4GMsY8WvEDmaEl54NOe
xW3tQmZAjgcz7DVgZ6n4x+nEYYT/5VRhzIWhUpAf0f8t9LsDpq1NzZ5vFYeOG6fsYWDYW93be09U
MjMEK1CjljaTA/2teeQooC1YNBKewNUmuRr0da3o6akpUcNuO6x7cEIUxeQm7yGKyMmZn/NMIBhM
vjCtJJTRhMYTLjB51dNzLOEFMMNuF7DOB6reIWygGencVit0EjUZiAsFIS19D3mdXyn6Jm7blGyf
SdtpiWQ8uEnnBixoUuie3Oi7uZomgb5re46d/QBCZZJ45uspvt1o5T9AjwNgsOSqp4Hy/zmwZa+P
+1moVcC3A0OEtNUNcYdpT6ExZAJWuf3HNmXHHiZQCLTeYPtFYvqlZefCKKFfnhatNEEqcZhy7gz4
k8m9fsdlnNC3JnVdjUvTibBWleSZef6E5yFqld5I4I1+iV8xJTBbRs1g8SweC28ZVxd6H3PmAYXf
TIVKcz5TRv5aqKiTwXWzo794b30xu/Na76Hewyu4W/l4ogX5Plq16tEPVPbmSnytGCkqw8S6esCL
nNoRgMGEQa1ONdtc5y0RS1c0NhWliq7HAjkvf4mrv919ne9SLPjz61aazjG2xrOeZn7z+ZLsYGUl
m4MFnMdBNjL7xR716Fm124GdER2cxUt8JT7/RedfCNHhy579gDRSaIC8hmA77BuuL8+21YlOYhWq
/X6dkyymid5ZOlNkCvgQWdc5CURk87YfrvyBofNr8rRXsK3oe3SXxd+BVVYHAYQAMGHVCNK+hVCe
g9K+q3RvnZhXVcSyYOtLPbEYb2ISpsR/SaqyiLbudPRr0euPNplAqMey5QheVb+mZBtAX4VX5vxj
BvXuQeKcDSFnvBzN6eT5zPhy6HJVikimhYIrfOlJ8qUr+NnIcofU+YBNAf4VHbbAKKzwJajf5+vc
X5VFcw4Gs9lCOCxG6mOgmutC68K40wKPIeByfEPFHMHwJfqM3g9Pd77LsAj/+dz2dhmWMy+WiZ7o
2Vtn3nQAzejozneLer0dnqzaCen4QQGZnFh12qhmW4KHnzgwWLZO9ZiX2fT2yzM/YEF1UgcQzQQe
Fuf3V2RC1yBp6bPZiDHM+2oEvXYnhEfSlRPRQYLOGrQZcAZxs22vwgWRRDeIEL/QZ+F3SXkvX8+Z
MeLXygtpsU4WX71YoI0Ki1DaTaou9LM8Vx4blKGAjbiSxVSyWs6APbVAFvjeBCMP7CwrbmxjBGVw
77V8NXmPJhj6zRHWDvSDT8LMDhMn8AcQhwkFS9mhQpdVVO171aLYXLld10F10I4SqVpomHxR9CN8
N6AIuJe55pIznQ7UfGSf8DIgMkc68BRIGUjmPXx3Qr2axifiga02edqsfO7IHTPxAOOQCBM9x8c5
wjWfFOPHVHMjk6XCwNAkSYTMM634MsIJqbxAxTbjD8pt3pmwq644+jRi+kz2jzAWZHR7urp6L1f3
vf73k9enp+7y5iApKET1SuJyDAn1XK9Kldo21YG6cV8Loep9TqWHM0OSIx8h5fFWUgc5WpXCFjyv
ZJ+4us4HZdinGdE2cqnO2LITz3yD/szKtyP2Qm2c0qBj8ADZkRHqkSxmp/aXKjmQALRww1Pjllez
wr3rRR9lb28WLFM/mWlaSJb00fblZZM0BToshBMrDZZNMIGgeUjL019j1jEBkvZ5rrUBZ5GH29NZ
9TbeeiU4QiIapGrLJNwANQ5g2c41Om5lnTaA+SLWOBq/pRCRR46dn0FT3aG5Lq4u3wFlXRSngIVi
Xi+Hg5PkZRCmtNr/shNPNav5UwkMunmv1wcETViZ2Y6rflc+yc9qN5285IxXHdy3OOvpP/HBPz5v
chug7najOpyCE6/LMJ4MR+Mc/UDNemBNrcQbYrJ6mEilu6oVZM+LN1kPPXt33DpT82jrr/5JkG0I
ODyiabxYjSMer/HyjrLsz2wbqOId5BVxtqvZgmykccQuj3jk33AoXmJjg1nwIEzh81odc6kJ2yeU
B5xcz9nKcR/1IoD5aNtC5dtpvtFpcyYRZShHi0UFXQz20FcsPqPVGP7tt3cPMDgC+A5rXZbmxiDU
aYoysDPJruRwrklBMUiV6oyLDEE8NJjdqj/lMChO0TTisZrN+j0XgUM4mkcBtZde4nqxvtclFCRx
lcdNfGxAIOzDjz9L0AoYUhfiSiCKb+FfnWqdx+X1vd/ZadlYytSlw51YLU0ZYyLmc70ETf5imU61
6z3MB0lTs4wIJLDhutta8mhX7kWQDoEE0OsskS6KqYCJEBTNr2Az3lKvfL7KmauDQI5BOzNfgeYA
BP+Ab5OwZu9HGadlB6+GXBNm3CZlzYReN2Vo0mBX3B0EDhn5YldxHl4+BK3nOpdwBGUVX7wOlnxS
fp5HdEWVl18F5zbKqLMum1eaT57a3+BfNtUPP2kuRFK0SFEIaaeGNgoDcGwm7S/+lEgNP23reIct
wdRDjA4MFhpvAqNdOddnKNDOXdQcfJohyIRJpkZhC0R/pXIcUF4CgacCa4ULBc4U7+wfnCYofnyh
WFJbHxR6gkJmLw0fhizsey5lTEyK6R1I6KmWgoC5RPm7jqgAuEdFWxp0pQsez0UqH6/ZSyrUG8gm
ChPJMJOP82Ze232d6Dvftxh1XXgU+XDC4Q3xhPrCEqYgpVoQly0NvfkY0AhmRwDJ92z6tP9DWFgn
/Ag2t5colEvailLZvhqyhT9pw+LpgJqJRoe6bxxLecQn8inhrwlPuv0tQZMTUBA7oxG1MpeOnwaL
cHGJbHphGkjjpMyB2b6xrqOw/AIs5bN2XGOs+KQVQP6X4fdv4QYkEnTlDQfoMRrKPoOo7AgagMrT
tzan7HwdI9HmPphKO88HuldL2w8QdXe9mRjniLRMJNl44cTHETk5RCPu/EtACGnekjXVZIMHgtfn
idPDVHhhMXHElwXurPWWHDYD0ua1bgum0mHd3sTFFPkD0qZJjPL/a3HUjH1m8cY9Yb8g7gTySMcs
JCl6np6+a3Q3QhCB3VRSkZ6vP/rJsyowGZf1ldMjc2qCDUkBGOg3wuE7YHpY1gICBRLc9LUU60FJ
OtsHeM3uEeqMzjuL11KdbJ3V588fatK/BY9b5dYfO+cM4yVOOI6We8zgOHlJj8K+qX/XyIC3PIHx
+M6h1ak0evkzF/WkTaWknHG3aIu4hguqcF0gcGgrwYeRUBc6O4uNfc9DWNw+BqpwgfX6sbLGupTp
zbkOkveFCaGfJNP28L+kKOr5jwCMab7M/D0HoBybPWdQTg3sahYul7W29KKv4LvjFo0jJZj7mVPm
62VPvnoWtGa4Fx1cxmLQeA/pP2WMZjvx70j4Un8CwPxpPfG0aJijy9ARG8NsoGeuBjCDHjGIQhKo
t1U66jOfRBDeo998FTQCWOU6o5khpSqEAwKBUxHcbq8dGp6Tovpnkn4okhBSl2floFCSI+XqLaeS
HgVctBQlwtUE1cuwkKNcfPji3l8V5+OetChFyw46+sI8Bu5nwvzD36nzucM4QFnVVfT6Zt0ldomV
GGxqnsKXUTjN67gkbLtLkLYl1w4uT9ZLK44SNL63opWOPGESdKzJNtpATHUlfKw3BPrqyZrs+UhP
JS4hd3gQ9rL9dTcCo1npfp/rWajuRW+yvYzxBRA1eTx0NWX3Rw5Mdbzxc0Vc5g/xmVAj+vU1Hkyi
DpDw6OXzPQk4l5mt16J1HlQU6w/g2FkHlqa7S4jivUj2DkBlTWpcqNJeWhjoYI7PYu6sRZmn9+/0
4IBsHUaWbNZc0QTtVGNyI73jUf0m5VwKT4ZxZyFQYnwIMk89nZLqZ+WAhFF8cngWhWGyZJ7NPhUI
OjTK23+PrVN9t9NFF+vSP696HwIcm1vsXbSnC6QWIA2bDO/9yy+MBx27iwFzs2+pHgn59pyKfS7M
WuGl/7yvxZLwu4OaDvC40clBTbjgi5Duv2iLXxu+R1QpHrYSplPBuwUqSpkPNm5ATeyw7YtLG0Mc
wa/wTZuJU7SFU5zbY/r70OK7o0Nce8yqkkJ44ChkuioYnUh0SeDiSi8wvrdqpdAtYfDwDps5XoSi
voaUtT+oqTncuyr9upkU8uhlpl+ciRV4VgjZt3P8rvInK4PuRANwNklD2KJ2YZwy2jlJBP3kxqKE
nnHAR2tNqGwUr+Dq/u6XC+uzq5+X8UBPD3QGUj2z8e/YHfEvpr5fglRpITlFVqA92Ip1SzbstFnC
sDljEfhR9JFlofi1g6Eynmf0pVvsOz9fW08R9sFx8zY/i3WOXJIg8lJeYdZ32ANZmgX02LANUJ3V
FEW+BwBvcEboHzWNBjPYbw==
`protect end_protected

