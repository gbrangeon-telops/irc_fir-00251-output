

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
b5iEwcuh/jbBlgyw+948d3lvWBbFsOTNVYtA4pJb/+7lAHor6DKhd4akfRWg+MPGWaTgwtrV3Hjr
bBdLdBNTBw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
VtyA/tLK0cCJJRwkcmojHVnJYFSH/hY10K0O1xHrVFcESK6dXqpZL9jghTqU0K8Rgfgyj2mbpSmS
d3OjaMJOT/0rjwEIwUBTQhpYCQbUdyb5e+tsu6Jle32rY2EO1nN6daySTSkOW0tup2zZBsIOCr3t
+ejm/NK+miEBBu1xCLg=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Sf+0xczGTqZZx6dcqp2GTylMp6ojNl/Es91rC3p2Qk7Z8FK5U8FSMHtByvmeihj5pitp5aOxAIcO
cjVP1mZpqkA9QTc6UkTBmHGnHSpwqkUrzOtsT2ws44zFj3ryr3hssigeWwtnVK13YgLrM+5chsUj
26gA0jBZIt1YnLsbFPdAg3CFuuIkHWQ39NEQDeG2BTbW5KtUVyDTnpctdLn+1GQ9lYJeC7lVtfwI
4B4xEL5dhZYik7uaLaobO+7jlipeHv29o8EQsg6BnOj1c1kxrXtTLsKozU5mRUSyPYYAw5cgAAvI
P9ELz58Fq2bFhjjPjC0ULrxEE7cl3R3lE+lEcg==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Qzj1t+dWRPGHMv8nVaAMZRu2BQPWmF3UL/i0LvBgsHGjHy3fNoKTLAs04wnbPCVtn8n3ytCSqZ9j
YDEGkJeQd/ctkBALil+9bfKGzVPGZiyWs36ilhf0nuaehXbM+Zt3Nfkh/wd1LKqVrJhOB/A/iGYL
jRkozXf4ccRU53dhQZE=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
eo3jj49OyneaHUaTvAS2/lR4/3L9GHwLzRAoxweYog0SBxlqFd2rrO0OlKoc3GfXgogda87o4tmz
l/UHxih0uJyK1snlhQ6A1EHKpMBpfD++gCN+S5IJFV1QgpWejKXt+0a0zp/A429l2cS7KMD2pUZc
B0C4VRE2SAMGJhfx1GIRczPJREH6ZIkDU1qmMs04rSp0PaGn6eV7+euaxeQcoqowg8QlRFnxfvHh
5JrqhxNCP2z579eEXYXH3AWOzWM/EnKEFUTbEaxMGP4W7RzgRCZvuM41apmXDWTVjEj3gQq6xKn9
0OWO8TXN0ID1dcJmFJe2x6yA91duGkuqWQQaEA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 43760)
`protect data_block
5MDxRUFrN47Y40TtQHsILMtYnJDRxVIaMnrZ8JR0k5DXniPHHYP4/AcfNHZQkA+QkGAZvnzP4wzl
jrd5CDiVectrVUQgIFabsiy3Rhu34wBdktTB2rxyqhlj+TKyb7091MR0n6gxUpge9AlsF+AZMTi8
vcx6PUa2MLZLXdLrP8hjKl+AWFTp+YM2a+DtgBlgicy5uDT3bE6abQw+zk5msXyvEqbJ1hox4j1g
dPsaYbCvhKMvyg/QbI51BtUg/2WI6Wp6nhihhE8u0TbfKoqKNfZGdF7dM/lBVLYnGogtq+aCB8dp
gDv1H++jDqq6jIJOuoJ3Fk9ymoTEvBa05osPRc9AfNEifAmaxx70tegwmArX118JVt+7hkIFFdd5
/MXI82WI/0mmFpHwXvA9gX5JvGAR+xiPbLCI+XoDsCaFehErC0ebMnxzDreOZITy7bviZSGkNl8/
81CzdaAXrdf6shqnIocpcf+8A85mmApvertNsC+F2ohOaa/hYw+HPYtC29ujchkTWmcz+abErRFp
J/EMS/p+LzP1YxDiuNbGeNOJEY8VhYjYY1503yJ7dnY2PYy9byQ5Ri7Be9W7uwQd7XqCT2ube///
aBAm/iamIG++Hj6uc2qZR8gqeIjlx2HqqPSUAaEsdxHyIBd0jQZjGoino+jPxnZgJnsTixaM7bVV
XSD8b7yIqhTg4VdlSikAYsYIlrGObU8GAo3OzKxgjbQIesFkXm/uRlEESEOGH3Ro8FmbGqhuefAs
O+1DJ3jeuiiMQlylNBuObXZ/Q+PAlYr4E5cChsIH2ev1a63JYcFF+wqw9hNo3EIJYXdEJJNUf3Kj
DsG2OMf1Cr+YZDfxZKzVLr5fEX7uYwAOBSWH02Gb6q2d0Bv6U9WIm8ZUOp9S6PlUoBrWU4ugw8FO
kSehkW49hI4feE3tUMbBcKiVy1xuIzRqBJbnqIjb4KegleNUQ3HH46Er7aIyIreCNrhbb094ca1r
kWZCLXFcZU3iJGaTjZSQed9YwGKNv4T2Wey0KChs91CHeu8ThMY/lD9nv/Snq/Nsl0tIMzX+xsaK
d2OnnY64+i+Db7t1QpRFm/L6+WEHTivmy/UoOoKBSJelzJlX3rOaCINAAUAjAuZD+hOSsOA3VelJ
+zuHaPDV/g0quB6YXMy86JiRDKXlMFCpD7AJFQu6AgQyiR++TxGmUqX8iDNYwoALp3p4RhZ4dOq6
M4YTV5pMvOrtTwIMswuETiDxvz+38OpOcFmKZoc/uqgK3dXs+uzx4UxrCT3Uqa8Ouep9n1emKl5w
TghnyedlkZL6pzmv2lYuARt4E3+do9n26pwpcYzo7pIOZ0yBV4TGiKmBDxyqdzkRMeaIOBHDkeEZ
AtxHM/oAyd3eeXXY+YulM8vYUr62a4Agln1a2w4bKZE6p2DzzO5HIt6Gp646sJ/cJvlaeXQZHip5
q5WG1cxPvskMgn/JjukQ68gQ2wnjIvuM2oVQk7qwvmi6tzi1d6fhTeuOhgjWPS8OulP3zkBfTjKS
DD7+6HGz8LktfTSWMvhhH7GSBS5Ehpa5d+O8L5vyyu+bI2ytTxGO60WwDQRnw0q0O7HMOocQ6HC2
FdvD9c6qFLeKuv+pZ4IyU8Pz88bEJA1xamp4l+WXG8NxKha5HdgRR7BRSLSDUex5mpKPXcctnsAT
xB8AtoXPdeakTMJSbbzfP4w2nlZrSlGpHZ0UbozhwCNGL7DNBZjheOZoVZDrS4T3tHTLTz0dlJDF
WBPYV7YeqMxqD4aAxQfWO/gSH+RoNNtYqu3NsS7H2Bcs7AXN4b7UtcN8cOpctvc2nDOL1ywoyWIq
6jNCL4c84PZ0AZcZK+Ez+YBGWIsweNl+UlCxxKbSpKOFb15gjDhGDI0h7TCqsrBKm981CaXLSt1+
/9TRri5jPkpNEDIYywgLmtGrUSRyK0VlSm/ZiTZQmkBjLOatoaufMdqv9Qt/U7jdDpCF5AtUyyaE
vWK4da1meltqqbfjak+kawUS7Ypt742oTFJgv3ath/Wk1Jo9aez2v0gwecq11ZJiIiD4MxBncqeb
xB5z8zKisHG0CjFcUhNMxjxibMwZXldcfnheI7g/uazMDLSMKAfUQsrpFQ4q4EdmtVHrkHYnpk2/
ehKZcGufboqn3FA8nfQjgi5u/i2pB/aaVk0Ok85qUC+GHTJbZ/HTPA7/bR4mkxZ+ADvVU4vjUzdU
d1vK20fmkTX2RrkxPFcFKyTcOMMAcScyCULVQdnyhGzn3QyqYgX1433T72IJZhRs7p7WKIObIieu
SVY0fCtYQd4sfQm4fsXw/hKzVftXkwnW5lOiWe98YHWk3cDPM0uEfc19LDOVJcu78pVwqsjzptmh
mejyNDZWru3K3vM/knEQpIfwQKP+nRokezXft6jGUXUaKgowo46PVHf68zI2gZy0bl4bWZj5trBn
jEFBkYceO7GZZWlzlKsLPtNx/OxK6uBGL4qSb+hrSWF1H5uxT5jOrA0Zyte0yd9yufV2geb19GZc
g66I4kjHBkb0FPEjvZLjG0u0nwpXGmw8SSSXWzUv70YWartVToNY3kdlXf/fbfOhxDJ1TK0f/ODH
WK0NsgsBJvRWTpidEPAMUXJOeJPzBub7QCFfQx+L8fo8TO6xKMAgBNraYhD+m5ACJROFP0j0DCJV
vI3fSNKf3ISTd4FOJAYrQjAoeUPxD9Vh+i6h74gxUwO8bcs8KpidJ/RG7y9Sq4uWopXQteGF6zxj
ECjvhPWewm9RpmRKLJqs5AxkV5t2q7qmK54dKgOj6kH4QQM5Fe53V+1M2WKOAi3Wmggw1X09iQUZ
0vZy5rstiGU9+PeSd0aZ4Zj6vkgjbWgwvU0PLKjBPPTQRTAlkJMf4vSc1vnWEesVyL2v8dCKOh/q
7XXg9jioORX5O0mb8OqadrzI2dZFxeHiTN/d302cKSZnbtXAVsK9EqyCi9wQugXP06TbS9p4jUBm
D8kjlPAXHa0GyKlNMJn0X+30a6zIEsnYam0UX8O8vBtSCXRjez+Kk2O3IBjK/gwW8Htj32a2CfVK
+8nWmaiqubm0Yaend9YgTnAaSauV4zaMQZO7UxZUSUN2/4DXAMacFYW4j0FYAShkrnF8NecUpYVX
6dbNx5f7DE7wO2T6Kk5BGliMqW3kUHRNB2myHb3ohAJACdiwKnlGxzQEQ4YlHBSsH5A1VeFF4SxB
FcUWiOQrF7RClMCjN3nwEaUrKOpmQLn5yF8veR2+mgPpbbA3qxhG7lY3UOWuilzxspsor31pbFDL
WajbzqpNSQaFTtZqOjm5G/Yn78Eoyt7JdGW1mDCP3mMh9YEObJH4rSsgyGpdqfKoEST0QdfBJT7j
TtLkWynxFNhcc/fEOhyO4ZOW/li5T2QG+sLqheEiBrLm8c79Se7mr3uyVT7WYwkhWIwJQMkYRqKq
lYOLuzp5aUHL/Y28ld0hM1awJipzsSgYWGw6luVvzjSLCJcZOWmQlQ3Dw2QplmCaoN1mZrHGVRmO
87dk6ql7I2eitSbg2Hu3eBTPfJwyMKMwE4IMWCbXbt5D3koMHcRC8INe3oS7jfIv8ZI6w8B//wH6
Vr62uxNQd4tc5InZ1AVNu/eNGTUcMJCb7LbvrA9mI2ciJ+F4g6sEtdu1D6oiXIDTWIIO900NwYe1
EPvYImMmE9TznwvF8MlNOgavpGBHUYzohhbWC53EFkgb2/WIJ7MRNIhmhqfvJQplMG/qw9y8+CLV
7Y5X6eXY3jHKBuXRmXdbuguTA5WdF6prUF2Iyww0wSxzWDya9oWdAOFrud0SUKdLbHjt+laWXiDY
4gYtI/axJr9eXrTwdNE9zbpd1BbxTSkhwlmQ5W5vvzPuO6LCtOjExrXmoqRgvn4y8WWOxXvOj9qo
saaC8bWlY7S7Mkfp7sW4wZm0wrTIF2RddaC7QI05BiD9RGhaRhH7aGDhhfz/SP8pxC6MhXwdRzIn
gA4pIJuc4ZcBwHdHRyGsBsLeSIRvaO2oz1TTRpulEyZb2CteYxc/1eNnHrQvX7EP4fMqys/gytPd
Qa69eYX/gdvEXw7ZGihJzTGe0Vt7TQ/nVX+aXUqGyLeYPno6cWmzYD5M5l0rCVZdHUtv9o4bcsZ0
LhRf1UxYNimDN3IXPCciOsPQ+4ST4pyCUvXbnaPWxVVpC7JdDmpslWHgrIS5Bpxq+rkcV66kf2dv
D+7THkj5htXhvBKj0L8k9zktK1AjVZfskaQoBIwe7uvW4VtW98Hp1y/81bC39P+QvltNp0uXgnKP
/eBGqQYd2EuCJlVM5d82yqVF6ZqRJW8aK7ufklOSDEuB3l8Qd4FS9sz2bI8wblJirakk3ianc7XP
nlqhyFiPOsW11Es539tHXCNajmTNsjlaA8tRk2+1+ttZDgKtvK6OP9HC8C89Q6u618Ubxyg2Nfpi
rj1Jk7xiEis96XgVVvTmxQyx5LXrnpsoSRXS+RVogvQzIOMKeoAM+s0zD9nrt9ylh0AepNdhyGR8
FWq/JPNbeb1fth2FI5+FvCWvUu2YsQCNBKI5E55//r8jWPyxFnMiyUi4QCz0mabYaYYblXBbVX+b
gXffXbiXXCdorJuib28TbVyTUErFLlIrouQ8nqIxej+DOAdiUrvQcfreUZjarLGSTMH6g3adPL/+
CqAg/u59KZHmCPuou5mFuw3URZCzjYfqyUHmzwLOuSv5D4FhGW2LSGOGe7CE8T57lkxRAIXgy8yx
+Gcq2HUcVMfEgHhWDHLyxL+lA+ujjgc9+h8ZosXgBkGmbeJd31IlEQtQPDl+85PWgrJlTAhU/XsW
3SAV/e5xDRfpEiWpZjRBB0KDLNuMYEgkONB6w4FatP+W9YE9+qpA90UkgiB+IKhqk9PyhoQQFsdy
ttWlLPZNkU3mfYv9lclx8/+KYLD8HPNJrlF04KPUV5Go1UPzn3cLs23yuyR0Yvz8+r7on8jiGHZM
07BujumqjghtfJO1L86ysWTEtP7MvbF4HxN6oYetMn86J6VWWsVHO1w3vRv86LsytL/3RUCHwqtO
ymCHkFovyrepIpZwXzM3USEeJbXScuDSVLQJQi5p+i5EX5QUkulhyxOa8RfKpDUuww9sK8BHSgg/
ISiuu/Ricm0K7gFZeRidDi7QVyRCzNsapSgCrk5zMyuxg+bQ0SV67nzWIvsBImryW0QgLNTHUCx5
TrazUhaGnnOuCEF4F1Flpw83putbtDwq7mj2KrxwG9qZlhcXSkrQk49trWIxKFul9lrpypsASipg
WB3GKI0QLoyc9oogXuNMgWvqayyzT8lV5kZaSm6kPbeL41/gx6yar/DeV8rvbsTzoq6kxAlaMmp3
XWojlVHoB57pbjHhdnrx0n8qwCRODh43NCnCFy9O0jGjKIKkPbaZSKJv4E8uE/2IlC5ebRBShLOo
PXuybS33OWucSDOPE2a+kVtLjxnDwSgQ76N2eZR8IjUF11B8x39hXLEwW9cuIewCI6gPoick1dId
0Hy8m3CCAFXgLj1euhqZJP75i/Wjm48w5bGAeKpzSYnX2taTg8rEHqRiDmALW4biS7mC6jCWGlp6
WWGmJpKejl9xZ8g3f7rlAvSc19tTTeI4X8MiN3zsBrnJJily4U9xyyj0yLPU06zlKuuM2lYTQtXe
FHb5cIwAa4dY0ZOm61aMZ2Hh039724A+bk9+i4hKWixJ1lyYQgrf0++f4yfILCZSElJsFhPvdh2I
7qGRoTEmKKqSg+yQsZ3UOObR9r9O28FDl6iq0QI4zTNrzzGH2CqkbSpGAXCs4c40Bt/Inpv5qKYb
R8MLyD5qWoeyE8IWE/mJPSXlsj/t2acE0QLSHmrY3FCrCpRj7C5A8PnQiAFWQomvA+mPIFlie/TC
zEeavirVGS7yvXIS0oWvoGTd65Yzuy2H72Jw0gts78sxzt0khyqr78Wzg238vJcRAj61T5Hyuzv9
a9T3FBqGxx04FiWmiE95Haa3beeNbusF89HweNV8iZ0Pju4EzXQUj/MIAryuli2mH+npTud3JiQi
7IAYzmtzvautl88oavTe1M0i7lBb5h2KCisKs15XdgdersYnRJKhBhbTCRnRMXTQqCpVSUPZw9xJ
rmXk6XgcT4OPsMbhDLk3feWnby5dgKQmUbDDKb2O0aonULdmEeELhGkSvLG5pm3hbHgNnCWeGVjU
bIW+QzqqsvbWDPnUM3y6jDNkNTqPywfVbU543EFFv5TaJWH55XY7rBbaMcIbnZq0XFeNQr6Kr2I9
g43qyQ/qnJSzARpKCEyUkvsyC29Sw9QUaFz2pxw1M5612OLAIrqYr95d0rWIisNBycS9QXfuOGKP
iqw60WF6NEFTvi+GECOz+4mzcr4yYSaJyC5NFJJmE59UGcHzsh2hyo1T1a4Ir21cyC5FBb5iFv97
oiNjJ0zOqgf9WhCYk4J37zbziGlviMX7OhwKbnCI7oRsiRxuG9jzlxd5PkNtwhwmaTb8aHmap/kz
wUVd1lN8WAOxnX9Nenjkq3tKa5iRTqqIfhPV9rQRifXK29Ss14I7r34BCwAC5txfYnyz6CV7FLL8
ESASjPqDKkKbYk9Sg+zNCQGdf2wgGTekiKOkl9cpIKDHPUGyL8jD3D3mXyJyPhVw4se4Pt1xEA3v
nsrkm4Fole8YK+xr58/IMov92XDsUSKaJGUdg30efxSBfIYxUWjWonZAIO4HJp2KeCeh4E5/c2Fc
DStGO53T7SHr2w5U/aUglnx+LvoQD71kcMfOwVncy/G1Mx5gJ/6ib90xkWdpg3t/13awpufB5EQU
fSJ4u8Vh1feX3KDlymej1VtrbalRuutp36NV+PDU8geTogY2x5iHUiP/dxF3aKGZIBRHCLd9gZno
rRnkkMkcfpQ7lh+veE4HjvKcSS3VZvecMAhp4dawItfe3be8z7ku9DwEpc9XzW6jHg//tM9Tew+Q
I5tZNHTvVtupehzHs2R/T0BKYA0339OtB+KpmpEkqbv+RjR6gOpfLbKIrIsKYExdlbvcHRA+kwof
LjhRpPP9eps/ULQnf7YxfWq74RiNTKzCdI7FMpZ7P9AvIzDniOi9Dh3+4STR/HHudbsVzWPy2mZj
7b6XBYACkBsF3YTpeIRqt2pPDlfMZklyb6p0YbhDPMFm++/65NuU/08/tTiquYbJmiDiQD0++RCw
NYo9/1qEqdDvvpCl81YgzaiBg/9GC1w3gh7J01HezFzTNbEsUkA2Jk7lZ1k/4tTlSj/S0CjfvcCl
0WQ3cxAqH55uj2JsuCdq7nGM556llA57FkH9Akm56B7bPuPp1g1+42tEeS3leGOSDSVE3cz7kaSC
/+H16Zp+/pBraiBZXnKosLO3xD8kSDUUoUQNIqj2UIR/tVG02pnakFtbrB9+8uFNm4T4VcR9KvsZ
4ohVr7BGI20ALsml3JKS3HJunyn3xXdsQtLjQI26AH89kwKJhD2V0/D/pR0RKteUSCnCJPy8dBjk
vEr2mwJCxnAT5NmpSQpx2fFKitH1GRa5TTkDwFhIvONyt3fOpuQisIULCH3Zt3Sq8yBzxoNa0Ylz
zeRooXsWX9pUwwX5SQctMVYdOa0kJpQV09S6lWZeWXiaqnvSm5i6XNTy9E81e1gXxSlMBT/jfYGk
Q/kMKaSbT31dB5b68VAwxushSaf5qZwUOumx27ZWBetDMZLLUPBq3/bewW/7iI0DuaDlub9lOJqF
gJka/zafUITchzeQPP0hTZ+y/L2/ED5LoR2kx+vN6gHOy6YS4mHL38KzbtYCv5iuRs5E0DVC0lk0
ptBzXF8/Qx4MtRfOQ3NYjtQglzHc5aTyZNPmLaHdFqA+7JvJZWwOq8mzoi7N4GQxiNcccBC9wDYM
IipEToucPRZRuYaDsqaXDUEWE4XPXqVGqxqL2kW8fo3iDDzjGIeK7mw6QEMr9nuABfRRKLsD0jjr
qmNW8A3WCwe8BvnF9XwBidxdYOh6zRSH1GQkT9T73ErG6eTWVnsciHjhKN8R2vxqkh8363/Ly/g8
Z6KAIrDzD+iydmgwxTdpHjxM/BmFzSeCDr3bbJiWJp/0h8W2dC1H9mShWshfYPvLP9Q4IMicctX0
lIGz6SkKMo6yqZEKE9LCERv+OfSnJoxnVrr2KO8lr2wajW7RBRQtNGO6at9v4ZUDsq3BqYBaezrB
4kIhIA5yKUb8+qiyVYhXygSdESMWRlyG7TAbQn6kvdbW+GkEHiiVPVO6LbzzB3a3ywBM0FIHwPtk
82oyv/0WeiW9xNMSaU0ewFV8ouH7MI8xuLVdDlHcyAMfrcVpJz87W2WoPfHZ8NTnXstyycwMtyzB
crJRJZL2XA8l2DURaPRJ889l96oTVX9sKPiU4DULwP2rNnq987E3bZKZEg7+bf+dbWTE7pXArpi5
7Jrh4+J5ua2HHMR47dXUefBQCq1ZjyZAo56d7qbCEeEesZ/RhHrC1mH5yX/LprF5zVmfEZyG2OYI
ptqWL4nzYPSNBkMTZQ44vjSTo+07B0uQE0ZftWvPowAIn0uBG/d+9z/tyQbfnVgyHr+On5CPkxQo
L7FhRtcHaXLF8Yut1e93vJ3oAwdo9dPPRc3ig+tChTKoi7TYL73WmAC2GC9Wlnps6ho1bthXkA0B
B3loWVGBmVcerfXWOZ0ITvMD4KIkKuj05CzPgmFJKjW7xnpDkBfOZ6z3D6Lbs9nN7mZ0xmiHbpSM
40LXjgn63VWCA4gkfzNMqAes8uN+uaRKzvyuQMgdty7UZjLs7jBMqYbRsKigWHNdHZO5Oq3ZvDs/
qTN02UTKx8Igge8ld8Fk/O8lYAiRreOmvVg0fxvrdA/pKVMBkaLHU65WPEhAcQjRGLmQG0yQr9cm
uG9HjbZguzENQnCXoWH6HJ82QHDhKax4sVQDKgNXSpAIZQboFP55ZKL0UVrsm0wG2WGtbC1kEEGS
LnCd4zmxOGFuZWOK7t1KkQWb43dhJqR/oJNsERaalVr1yx9I2lvs7ETGG/0iEXs2y05XWlKWZ4Cf
seQz3BLLlr0IRgmXzRAP+xYMpMaok10q03O+bMupfOOl/IwJdqZ4OYY61ljQZmMy0gwpzqU7nVOP
TLT9VDDgSIyFsa/QI1fMCrjBwNJ5JTnFRJ1YdyPR4qCXQrwXgXHZ42rCAPqbFQ1M/8+KCFTooI0X
z8t3IOnD3ehte1RkwlvNJ+bIinUKglDBUvMrkx6U+ticMm9iNO09gKM5FsUJ4cjpDVM7S0NPOz9e
9AMCw54RyiD/M6bjrJHa5cD+E1TajmfT3ntFDL77jLBFB9oQLoEoPtHa8/N8yu2YoYiNNe+3q+Wu
uHQ4HWrLtWJX6ngLM3Pi3g3M7Mum60DY508OpTJXvdCowEXYaThgS3R+6gI/1nbWK/V0+nKTiuNi
IRctzu6qT5+kN+8RcTC6H63SCwy3LXv6IEXOO/jvzP7p8a88naEfm/SatP7Wx7avE5cdGidLkfm+
WLsKUU9SsRtIAAlvU45E5xJL+lXcPL6BMYz2zWloa0mheZDEMnXIoi2HKJgNMy+8cvC69Sbj11Ub
JM/1JmGL5RIO3QT0ZLb7oXXxnkYAa/n0CpkGbG9d1ujLkJsQwXR+ugst3+V/7rZgODy2H9+mjLmK
QDHtBdr7+Se8NqfKz0S1Ga+HjKps4+kU+bo8dluk4CW+gI8OdYD/KdDeaR3btxoeZdonmhO+9zYp
js5NVTTybzAff917Bwv0vas/pi3OYuA7B1KtGi7WGKOW0AnZ3mleRlAkNRY5W1r/IPH+W1rAuAmi
8qqJA/HqNqzuvr1uI0RROpxOu0PzLPQFnDMP5+2ovPfSSBwhbwQlmphgP7eF3aw+FnV8KxxfffWF
uYgRne2WeuXrLwm17a7hvd6g3QnVVV98ZBsRc3Tv5khCAiRgDMB8wP+k++yM4oYVL8p0qxnKA6DD
2jeUgAlcMyNONf5NUUqYOgfdtnDDvcAw2eZI5VvbTtf4HL4N2VntvOY8iOsnL9xdGt3QkoZKsR/w
MRKBulrZS/uqE4a26zPYP7hl5ZwSHJlr4pL9YI2ECLTdDzKCR/9PNYwoD8sPHn8FQXV8J6qnAt1j
wKuZTnP05MhbJqsEUeC/yY/EW8Ia4x7llTnGAxc9ODD0rNpekj4z6T8Yl9kipMynxAxnpPpnQnuR
LeRKQqVnFKJOcdLWqORqqHPm5AR2zhFOpcWjwSr1yRCrUEMpGz4OFwoNFa7sahZAjTYozDQ2prp6
rG5RT1qf282QnpX9IN7ow1MPOkDJYPgNk80ueF3Piw5L2sD8U0XsQGlDPyVnRHFlYBRee6FDhHo2
eCLEz+Rg7DeVG7hgmgpfGQD6N2TjF9K9sdBedy74ObJzyrvpiEJrysjuldow3wv1dndbFzAxZbLa
GDpV9hTrfyDjeEDKXTfyT6ml3g4GGlXT+bfyE3cwe3PpLzLqk9PxHVsl7FJ4lZ7L8wLxMIBNv3M7
yBKx17UxTyauNGSKLVA9Sshp9Lr3ysySw+2EzO+kFZzYHUgloICTTiDmf601IVhezeLNGeV7D0w6
Ryr0pPZq6tEv7zGLSk7Uz8+QZ8WUjP++Jd5EArLz4Bqy10GlQz3GL+WmcswT0Es05cRYU4C7fWDY
Iu8YmBQ2ISwV6KeCS7FQR66a0HwsGRRt+iEzdLXdKTJKSD8Whx1mUqI9ahFynU9A+MXoX+7Ob7w3
PmpZ+Nxd27F18MijT2F/VQ0UDPROcGpNCpMhlr9xgycjUhxhxSNcpincBt0E0g02k8pV9q7q2904
j8Dv8/GwivRY1L27bC3dLLRaoRmFFgptdUtCRYV4dxCIWQV41OLhqx3XO0BKXMNGq8tk0H4aLV/Z
XE1+Boyo/N+f/cuBY86pV1OxTuWPnnEirbLPRvvsz6sEcmCcHZ2Qg6IfFSJeVmfrxE1lDQwm7y6m
uZr8vHHHsHNPn6xRJbcIV9rrAsNk8lExmo1d9IsEAhnlHnWKf2zePADj430IycB2IWAQuWHMQCT+
d/acDnZylBZs7qOopsLaFUixRcwQyEUsU/qm9hBMQmM3JiPngbiDB4U2CaJyQjcFHljaVXQntB8e
6WQihKD8hqVCFm+UPPBexlKmyoZZIxqUVKel5bskDVEnBri5b7cdbDXoIbipZckvEJAUGt/xPpQM
orphRd/ZVV/WhV76sn5u6cENfrrRppdzqkqrK18y2N/Z/3CCf09TUCeZOmwBLXde8T39ZEOCAZsi
WgCBnaJ9bkBL+XGKp3VoY7Dffn88EUDfeD9A/UO1YXbJicXKIZTtPMT/5oM5MvhBlu3haYEBgzOC
4dYAkLTJpQJFtQS8Fu4OQ9TGNzf5o8ninMoqfqSXfjbudWRp1wzTq9n0blh5+obR6kNdSlVmOr+A
vk3ybReToKpnFGZ+rEsAJLJ7hGa6+q/N9zyxc735euhrW+7fl7RFLB4R4und8ijUwSuYJ5zPnDu8
1J02NL9wU7aGLri9dPDHzPXH08ZqsCjlUYydxG/EGtWRC6023NTLVAdhVfvhKd6QENJ+3hVIk9zX
8SKkrgozrmCsiWpzDlnnkHvXGHQjovwShZq2WjanZUZBhskeZzMclbw9hE4v0MENnWGTOnZw9409
cE9Gs3T6YOe2J1kvquaHnv7s1mqCU3fBl6KZUK0RIPgmLYmfIa9r93Kroy35nG1Au5Rmkv/1mOrt
U9JkhnarMKrpUsBRBEpmfkJz9gXcG/Uf+Uwp3vj9UKrGglQgltkz17CrioZoHUEJP/rXAQEfWFHk
vpcNRQoyMtMz5T+iWLKW4WtIvkU6EbzM1rp7p22RW19t8gzDsqi/bzKJKpMPYRjh4og8GCYlZFCG
54X3+1ch2MS18vRUlbNx37UOpq5Knsk+PxzsNUwnq9Qrml/QnrKpwqozw0jZ9/6NYfhtlapDbfcJ
bcHtdIQzlRmpq6Z9GXOrLYwW//sN47v4Dt2YStO1raI5fU3mGHHlo/KCDMoK1PHt+n8KDe4VySju
Bwp0sJAg9vthj0zqTCoXeffPx/rXYVqDvfqM+xyd17M9Rz4IgrVjzchThoARkNRebE7ifcUP8F66
7gdwkmd3KbZAaDhld+YpTDe4XGAoGOAq6z6Nm9ML/MYXbbnNnsWADW2Xf6UQTGGS1hTb6p34ZctU
6J0fvazVFFqDpfIcFX51Oiwt5PBBRgsU8W1mhyCxw3mZHEePmXrmPUFW7MF1wfXAg+zWaBYAfEGA
umxPirofv68qyyLBFGOmk6/0YRQveFuc0CLjbYCb9qxv1iPyAmYGtMttVWunG/X+6q5VnmxfIdSp
cClvWuXHSTajYN+RB39DmoNveVynA30MBT482Ka4QILiChkjB6jnh1tZQ3Pchv3K4l/kyl3z8l9u
w/YXG4NktzQXxgT9zroXx1wE4R7NGRsz+iuQ8wnP4+r6d7oeiKRP5OcBROSlxp82h3cCvmVMt7SA
oHgo3mMR+cbC+CFJoUjYsSUGNUs/VpJavFZhLILcDZhtN2y1lBrebjXbz+hYa7WnLqUHtaPyoBoQ
gj6IUhRRVr+zuOYfw/IXkVJRkuYXxXe2g4WdebzF3I2biwOGt8LK8J+CqX+6ffavnS9mlSLLC2sx
m0HOALKGAOUXGDUPqgb6jZglBavFmJPbhhcpDSaVluySBvc4yglpHb/Ym+h6sXTz7Avm6dH8CeCp
uhz449ab9y+UprP/aitCoa8NfzmRZNwbxUjhK5gFBQxdewniR/ruCl2EYZ+Xr+p1xeZfByYtRMWN
DCsYF7n9NDkB8GMZcsKS2lopJNZ0Y4YHTOiPnzWWYrl97kDE4ZvUafLqoYssSIyUi7a9B4btRINc
bPhCk46qraLCl9HGKiM/5DdclPtQ9JBCrO9giOHequBqMOfwD2JbL67/0RH/QN0EbbS6XTQYpR+x
DO5QdtUTtGriHTGuUUVHpfms/R+ZdP/yNSRnNh/0CgxsQHKFmDfbgMGbeJzrHIe3x/FUhPOA+igj
ympPVK2UIH87G1XzkS4A0ZbvLGd7t79Hk5v/givgRjMXnNYNpYuTvyBTZ8y2yPdEFDIVGGwxHrEB
NkhDulFwxjbLJoChjL8PJKSEYVm6mTwsXiR7N6YAclnzztf5+9zXt2L0s/2XWDq8XOoM0Cq4QtJM
Iukpp5RLHffcG0kaI4G0It7P51rhFJjr+HV8MSb6jh0NAatfVlE9gK/5UtE0HqzgfwncP4bLw97t
mJVbzwshyP9dEUycBSDZwecC5J3Eb+H8zWF9SbmvWPh8E1Ll6d2bObNVX/dOQoSlvd9lbHIG9Ja5
vdTd0Bc/KyDMTNqkhBDuu5rJ1eOAqRzQDTS3ukOewzYHZ96WAQTIdAZCSn3n9bov7A51jDlGT+QC
DfwYK5U/dqQucRi7JjBRBkdCM/Y5rD76e/nSH3yZYTFPzuHZu7Rs8cPw69xmSM9L+ThYppjxxQA0
qhAV6oCU8TDCL0U2uyyFI6yzubHtK8y8cre70tZIyC743o0QKxbjsWb32n9CkxZblQ2XuAXwRMAt
skzrmSWFDXUWRGtSCp3VHfnde6DKcbuJq/oOxFFDY8BRHEwW+w+ahhyg5v9ER7RCLv11ltXnZD3H
rwD1wVuMYpHQBgva0SRcGyTa9sWjnBv7fctbIKwEkfIg1uuGAHf8PQbFzPqHNGoJRBpRgB7GK74m
d56kwVPz17mz6iITE3I2AC93DssU9LdFsN0FW+s23B3oq0sKvlL27fu1XA/jsHShuwcoRkiAZMVp
BrXEsH+mUecsEsO2bJOkfTE30qeHeMo8/bDwE/r7GefK3jMUqCcirz3h030ge9gkfc5bX9BdaYKQ
TizXrk9vhpl/UYHWjMSf6B5lTQEobZk8YuM+EVfFVL4PM1ilrsNlv/sa5wPvbkg/399Ez9Juwrtl
XwlC/2qlGRAYWUmAZ9b+or0X/IXymo4U365eYJ1Qml/Rneqp31wr8ZjETs/77XEYMlwVPs5kGMKJ
J6k4Jxr1ucoTIy+6B0p46Jx6BDSb/ZXE5fulzvo9bl7i+Z9EwzAMGEuvMqPpT8DXUCPIoI+lw6es
GmXx4/k1Id9WyezNeVQ1juXEV1nY2pHqOCp1nSUmX55yfQa2GSwCDt8YvjlFIs6/4+h0KRPbskwe
kxgHFjiM0b+jFh/lIAshZXDnPBDTiqI36OW2M2WK/A0vLekwGKkbzdkVjJZvNKM8FrVoKq/KS7j4
quQ5nhAS7iq1QNv5vionugFUqMnFKLartFWPgzABCUcbMODV5cT2NEXh6y3muWtmP5f3pxNkK/WT
CecsHXCT0iTIJxRugPBmq+ijkERTRbB+/6JYE1LRpX3UnYbG9UnDtOzP+531MiUvsg1+DxepPMnu
I/E2LtBy5bgTlxHL0mgiyZ14hMB+rFMEyi4/63eSSsmFikcjMaafUvXPmpbTV1pLvBSnNGssFKca
X2kcjbNqpvSKND6hv07JPtqDXRfr/SYM/816W/Jp1VxsQZ0XSMUCun2IpulCn6vnkL9IsKouexxq
Si70MHoipKfxNxdKQ9GfPgYGfGRO+30dp6i+q6nYWi42ta/140MysNrGDU9k/9nDk9q9QT6wkyE/
Je/hr4rlTp8wAMJkF2pJnQ8izY7nwK/Ptun6gXTMZOgeugGwS40fG1xQJTNQ3RLBXjtKP3wDJQVq
RBXNqVDZHHj3NBuktQE5zcjDQ5ti+d1LxHrxJISXO+WXdKhkkxKfIiteoma5fPFnQnWi5wJhGiLG
mcd0s+/BhdIHsKdbOOI0xe8e1N9HxzK6pKPiATRbScIYezWZ6H+2be5O/rDUT2Wwoj4pOFkKL+f/
UXO3a34ta48GYdsQkDnpzWCwjqoNxyr867GyrGGy/9T3Avt9VWGlWuqpqFuYdtHNKX4hugf80ZeE
2iKXoyvZv+qOhOOlWG/ypGM1H5/tLxx2IvK7BTslI/uvOwLo/yX3LVbCQG7ieCdBZd+ApSJ1to/2
0xIHLgTGMezSjrI2aLmzOAbYnrF/kJblIIfianTR3TRKFjrqYU7Yi56WXXPPsYN3S+4W4ZxKJOtZ
uqnz9g2uMoJazu8fFKOoV+TTnm0zQHVc//2ft++W6mlHkHKz8skLDXoi7ZNN5mqBJ+bK8+9F+EFW
TTBNx8kOHp3gHqWfxuiNJNb4RdhGD2OKxYIFWuzOuhwAcjAevIvzPP8lClgqEuvj36nKbzS/4f1J
AWdWDAtSSLhGC/Gc9XJPU5fUe/gMu3WFF/Ynqk+G+DKSCl0y9jaOm4K1hCxl2jMG5L6z1Lu4qVtb
l84EUkDYMRHoJTJqFawcZuEiujaR+LUeSuWyNZf+OQWuZkfXvOJz4VcXPhNwwvAuYAkkxmTI2PxR
EmmQ2WIydbbxL4+Jh0DdLOdRKkXdmcEKW83rHGPL8TvBWoqyPL7usi12UwOh+awvhOBMIwr3p19d
FXXbhfFsu68bEf4r7N2as4vC2LSdSx4iCTY9xnEU5VqSAu2+Aap4lVvmAAez+XlX/U0M9KtA9/5M
D0E8aH0Rvr8n6PEHhL9bncBWRPziwXxQe0O6PK6c/uuVq2KmRD/DaibxxVN1r+ZVw3bpiI+rNbid
m5WQI168izslajPY74YblxC3rxC8FtgekGxCc+13je8iBRT/Y+CU6wbvs60maSL1fJkY9Q7OdR0b
zUqv+5II674S8+Cm+LRC/06zIYVMRfN8hZHbORlYRqzSfETDYcFkw+nHIRkdjIsZWB8BVPPB+znI
3eXPCIT+LY72DeHe1EADMp7OnTgp4PeLLBGbknQd9zI4C5No3QysDB8ItdcGLs6ByZgj9y44Qy0e
xlfkyTvy6Bp5ouMGg4+hx2U0eMVp9aJy3GxEEb0PGdDsbNAb3s0LQEd5fzUX4B46w2vLFFOrHvz6
tKbi2Wm+pWF7unlZk1pWl0Qzqicy9L/57Hi3UIwCeAtjqC/iUEVp4FpZMzlYnVGTBVnrYdueBtoP
yU3eBjO2bLmuUDdqIg3cwdvEeXca08DIcy79JU4YShlwCCIi3KfjXxz32ajUgS95WhYt83FPMw1e
bFZts9fUTWH8Dk8M1rbm+oQkwMot/qYS8HnWn5A53YlrX/KWx6fuIMAG0KsOVlq8VnKVLCduYo/s
VKXY8ARBoAhgEgyP4dqQJeu6pGdKJUA1B/H/2roeHmVM2Hi743+4xEDRrv+C3ecJZNqFRP/wwKNN
SJG+QP3k2Zy78CiXOLCuTEmt9nB024ymAeZ93oj8D4/X8MslFMYrvlvf3Krp34qUMPKFnYVTty54
DXWkIOsAqZQaICDjhiulr0mPKEl5ekRNMwXtVahyWmW67HHK54EzY5ASFzj0Sjqnf6XATXsvP4hH
PSafkGSIyNDbLLwEnsc6+lfc/oxG3gzZ9MGZi0jMy1629FgS4/iUgEusq/5DPo5qPAgoOVuuQzRH
nrR1eFlpGRpZal3ezkEnwFq2BP0WEubbxRc+sqSzFGo+4BF8aYRXK+pMi9mhg60/E+8x6heHsaQV
dT7uJY0e7J3puccpMoomWnqmy2mjY4qOwakbOj85Lr0hT/yCBUvDgGQY4Z8uqFhg5gwPD1FMkBWn
kM6lUUGwLLW62XWE/5M+sVBZ4j5NdrHdaiepSIEaMwc+BEqlm7RbdetRrVF/hlueX40QG2JEx188
iyj3Kz5fv/xCOOfRz6Ucd8Uyh9D1pXcjJPcF92dLrNyq07Yg98NKR2yaVbQFuhFuzkY2MxTaOFxy
D0Eqx6DvOn+x+FYYuHJkEDRwcBYXffftmXQdvXSygtAWvcaDSrfK3Cqq36KpAQ/7iC7SsoLPlzQX
QGO2EQCGebKL7cW6vkpFiSzBrRgkEb66VtR2+Q06H+uZF2TSge4FpQgfs57L1Gms4nt42TIkOMbw
YZTvvfyXXgtFiAZwneKGGbSAR2B2WF6F97j7nw9E38kfuusoy0HrPOW+OQFxDSMKGFQkvN5ER8KA
K44F6fw20YxW39n5t3LoFAnKGM2idZiI5jbawNjTLMYhTWXsH9DbtorHtVlsco7m+TXYX0GDxHQO
890nByOYJfULCPkkTBnh7tpRHOGo98YpuJznPMUS7oCl/yj0ZnlkwnOQ7a3JhigW+Nl28iNoPyzI
je4W8hSuFdiRZvQJXDoE/IKdze22CTk+j6ufF529p1TYDb62+cL2CMhIOl0tVIq9UjbAHCrmO7VN
l675RHK/7D+6nmZyOXKhN42NgMcACsVCY6cF1tqB3xYSQOdgFj3D0jTXMs6iePYsLTI7w3k99thZ
0RY4TsWIaFcwGRmRg7aOqPnrvyfA7idvLZwJAUOyEHkXrliwcn05CAcsfcXSC6iLuHDtKxAfIFNZ
YAyJkcVZJ3zM+OKKiFjh5iX+XgcdOwLL48HALPbYz+rwrUultk8hsMIzFN5nu1EbEzmDsJYK/xXJ
J3qqLtK4CtoDzVuEOLEKDnL1C1LK4kpupM1YwrsBj7PwboCgBdf/NvWs8JQ0b0TCkeDy0RzxJvcn
5+TmnPTbRWeXt6qFWjdl6F+B1orp7mSMlqQVFJphIWRTrLQQBU8KD2QsvOet6hRsCETvNixJxEer
/cWNjTPYsWUsHF2bmAEBXxmJd/J5Tq4AzXd+ML/nYzqGuNNAOHp/V5kmX7R4NjPPP4r6MHEmK7+p
kDQuvlJraVGVyhxod+PwGwU+zfjhfUGuk5IfDDXsyIlxxCuOnHx1yo+PtMhZnr+iobgF0sb3pLUp
BSHJTQJWswrP98JuzUhKzsx3ftyoF9fbKq2BL6PSi1BDhL0JPbuK9zANDUNNcmmrDjbqI+eoQey9
nomryOzgNRKdSwJqVZ2dvHtSLSpqxL2MPpxxyt6DHziZjt/y1l6/wbOORCAbv9tDIVY55vNLG1FG
jJC8JoZiUnnG5/bX4+RArHvmebGxL7j5Lw8o16of2Xpnlotf4SPLRg0XdsmbqCt4xA1BrTTvLxym
gdxCx/BE6VhhToKFxCQpwew3prdpbA9GUtIbEoXu+R7OaQwLa6zGL6ps7HEE24ssWpcwLNxHzX/p
4vVuxEiLe+nt7nb7KvAlefMsQ/5GSHOwovJ+YGL9enUmFYoFro4slUfZxOmRNA/jKExF0ScbmqZG
udZn3a1vw1RANTWoDbItbugROay9MZt31et16JAJvwqvV0en1odG4Mmzo0F6OfONn/YfxnjAXKjP
axWBcY4GgAxyqpNRHLK6m0ABWxFen+paOkBPAI+V4B5lGF1lEl5YJPkHRsB44rlK74G+vYIpdxW/
GB6Ij82Yv8Ig3fLUVv57hZ50XYv9my8mhu0MxIQ40F0Qj7UYxjRCEPnioLEytEpI9YDf6eb1L97Q
lVtQRZr0bDrhQ8YR7l7GHiepP2SKTq4yEbp1PKxutgGN+5Yy5EccoCKj8wriGaw3qF6PCfKo7F+g
jqJ7L4I+gbfP7ByQ20uk1kwH18sV5oA+qETCVBuWJm9abvIR5lzUSTWV8ltAliiUezt1spPv6Vrx
F+JvNc0vTRVJ4nqnshSdAUY6cQ+PSN1vNM+f9ss4qAEEUEOxoLdxiY0VRpvNzLTzET5Ym1g73HBP
MUTCXpKsXfIb0NPCJ0UV9331k22p0dYyNTG+dR6At/TQ7iAHCwIpOidCmwie0JmIJpJigW15X0bq
sbncWngl4bbCyuc8W3srPd6A2XbzAAALFXK2kS81flk0TVGw6502us3oKu6FPtM8i5VIjkhPx8pD
6jL+fbyiti+nJkEH7lHBXi5Yv16Lh+WRXY/D4GXBeDwyrOjq2oIc4SLpY2YzGQuJcHAjomTHCz+s
swMofNxElb+YNfQaowF9D2ST85R/mBkbX1zPy79CCuL0lSL25bVNKvMYl+A/94WFBnyCFb9fbRxm
t3zuc5sa6lLRfU3wHpajhlLeBN+jOGOzoskQzPx7m0JjAWFvgiSbtdzJjrI6HaUyrHpE2IbOEUv5
NvM7BtOCcPAOMli3icfzfPlNiqLEctUxAh/PCCqiF3XfC2A/ERjkI5uyVkO6Xz+2Jl7+bV8GffOA
pC6cCgkW9pERtcI3ElWf6OziZbCXH5Zo9XuFdr/oA1J9kO8JwDxadpBBwu+s4qw6cnX6T7lEfXFC
2lXApoWyOJHRF+O2it11nam+ObMx2N29R9196rwEfIdvN9McDSaJAAWOvBdhDfRojq16DLAd15b4
GbgW439ku5B30le6zcoNiWioP2nVl64C0ojEiakGOp52S+awpKhLRhotecTUnY6OS8uR620wznYz
ClkwZxL0DYnvRPR9jGsFyVUFMf7ABYnWpRJw2v/wSvdvWhMeSH+4AMpmSaMDaK30fNhk6jWW6DoI
3LzGbMxXnDDAYpz8jLP0ZMffUlhZpjozFOeTa1eUpE2HQ5bsI1nsKZUM7YxJnLjScXwdOaZcaCX4
da4joUWUnRFzmx5vMETU8pe+JVtdeTgiUXDEaL1BE0oH5qx7ZWrwCfLhu2yxoO8H5ubTbzspdptM
Z11NDnPgZ6qBKOetT32hz2YD/17JfSlM2+D0wFJjp1AQU77KWhayWdpjt1h93oHMX/XbtNpXI+9D
HahJFrcKHw0ZmlTPJyissvZWxJ4Suk0W7E71Tb0UbrDQ7YQfNSPnYT4FmDsc+XU9dOQC2HmEB6kH
xnb8xOQzuoRUCWCNC4DtwYMf+ReC8XUMyvXPMBh8t+/dVwXQF5QMWx/mEztZvzBq486lmhaO31Lf
Y+ybr8TloavJYOxdMmGMkq/aiYMFJzK/RWk64L0nM4g41jxHP2TWYX7joxv/faPCAmPxR59mHXow
4tTvUZFTnruQoOeO7oPyyE0yoHpifV35mI0yc4LI8WXcRg2OqjEwXHG6WXxAM7RiMmKis65jOXla
tDnmywTqOG2hYqf9oiYIqCpj/5Nmn6IlHxiG+panOoZwEiRaoHUq47F4lxtCMt/LHBUcsAoj+TMX
KFUaQB8oihpbV1z/98UbfaUz25EG4FTsbsYP3HT42EL5rjWJRvQo82liutY9Xg0xdWyoTVSbDQSv
VTeASyChIB7gOKlblHuSPdeBOirVX8r/9bQCUxtAnqrVQl++O01P+oBzBYuI7Ud98Q430PajO3C1
pyUhw++aM9ffe5dpubE0g4+y/Kde/yvg8Rc4aTvqZdP1SzTk9iDIx/7b5Z4rIJRV5CcBApsMpB1H
be5RUHKVbRve98sPvthMoBOviTW2kRUGTCao/T5gYmvbfFSIldLrUS72/5g6opi6qHSOC4CaIKKr
eNLXNBMxIoz9YvO53tl6c7f2cwZt+qA3x3W/W0YO70ESuGL9JseSvkfqUnLQoMEu9RWRbFuRvxzh
McWO1AQJp/y7c6fsf0JYf9eTNxYP+rWvjY1tx2XZq/php8T2lcd7Nbw0+Rreo+rX96jJ66BIHhaG
wf9uXmWIdtr/2UNIskfsXPRBPU6EBmwIO8RMEIGYvcbfiY3+OE8vKOnsEf0K7L+oY2XXGQCLhYDm
DigmeKzg5TCVuYvIckuGESJo/OUhT+8Ce7eQq9/AN07fQLM5uiBiOyLprfSIKylHywGc57a/G46L
1KlQ6KTzIsLXGyyofM5PicYYehotPXkBMQUzgVx0I7SITLSiOHUSgkvoK+tNeKuIUO6SsGEPKvek
i5tn4Z6BuLHFtRTkjMSe4/PEkUR+y40lloMsDkwtoYcI2sC55v/8BSaHUQrKBDoNu+2Z03VIymUa
fpXfiHeBr7Ig5Ou6lXxEM5suQs6XLEnerEgrmtqBqcnRhEDtto574zmMVv1wgSFzhTAOVoeoz3MK
yT0VQSkJgmS6uoo11+7QVM5yMkVOIwKQsYmf6qWvpG/t5Y1bYqdpVp1qj+oR3VaujAOsZc8r5Xt0
1prjWn0wEpCDqkDntuxneZdfgXv5S+Ll4RpSkwWddd9qulNUMRZScdFA1ONOlfFRBJ2LcFkwG8wL
1H1V1mS74mj4Vlx/5WfBCZy8WNGja3OnFQVaeJmiHAP7YqBSCmZdu4VmrtLTeRTu9e0VgMvbtUiC
Ie306LGnGcCMSmeH1cqFLE7YHSqRuZQl8hQSJ+JJp9p9wPmIf3aBcHzhh8eJNxLiPbli/XbTnLPy
ycgcFEbPkvzggZ52k6MX71n01ZP46NxpwanNrTICvbS0rbgSurOU8IzKWlFBt2e10UkuRjCCecpq
bCKrK0lzBlMC5SS0HBsJPjM3lJNzS4CgCHCtttdADk/t7UtXjoAfOlt0oF8z/wi0swAsaX6sdbeJ
0YNRv10pZPhI2EXkOWEG4BLSmp5ff4LZkRHTMBHWw48lGbiUeyfFwHYoM3/k7eIR0kJeJS1p1i71
Sh3PEFJCaIMMaDZT5jNCcRbuuDsUzZeq8sim+VR7pvF58CrLjrrQk72tEXF4/7NQarQGYfi2GMys
l4eqVd5l2Sj20y3NczU9CXzbFX5/Sg9E6YOzUH6OuSbDTa/SlJwMad9/lAToSneviaAzvESl3Vju
Ug171xBxrq1RcGXAD5hMA2dRTbY6EgyOzUIW6P8NLYwTF5w3BYJd/L+4g7urfUI4gm+5GqOTt2LC
t3IRaM9szm4N5NmKmLhHNLS7nL5q37KW6qR9eb7iC1OXQy9sM+3hclCZ1phXuo+69WKpwl/eODdM
rjE1ePDGwA0xpwogalGJ3wo9OXKK0tBIZY5RWXUAau5eUxYAC3WXYA+Yg88JIfJLff/m4IStVDzh
XGMVxeet2UoyGfqd61SSrJphp5ujB9N7+cGZLPjv9gpAnPik0rG28fA8bv+VVHqmjvViIBhSZREu
zjx9/GwbLnKSXDEVNl1BRbUO4l3hS5j0rir0VBnMkvUzX8NoihCof///uHsney/BqC9DW+PXvmcu
A3TVi6wO9cNdXjG2z6OpKOlx5c1DYo9sQ04VRHuoScetaU3ZbaUAuKIiGaW6AehqF1hW4NXFy9dR
HBopUda3zedCSTRWkIj5rI8tmLB4J3LKNCiG6bGf7AqhTz+Yi0WAiFp8s56zEfTCEirKGOlhEjNz
Z3/RLTrWrtPMU9+It4e12qpktYwC0YQdLtOckQs0xIr8heIEBWMmGx4T0l9Icpuh0eqIKsEzmKR+
XOakMvOj+hn5TEtCEFnbCaCohBYmgQcA4i92dzEYzQ+5/VqZGnNytEmvaS85JvlRfDD5BgfOMFO9
C74Kd1+REwe7tAsdGqbFpTgRcmXz7BOD2WlE8Uf0W38ItWWrFX4g9D8W+bQGVrFF7SrERgijFJlJ
Ur1SbLelyBarw7FPp7pBFzDs5K8y1OdAxWfrPzWO5pRkPFK58M+bp4wjT84H+QH29WtsvQfkTR0B
wATD55OBqc+mFsmekVwG9lYk96k2xHMuIgZTq+7GGbAGFLU4W5jJjXHO1fqj67neAftq+3HmRuQn
DhMw7nVzC4lnvjxtbFuwPDCPXt02KOVygiGG6C1zSlT/FiHcmh9fwJoXCTFpLcLTgKww4exEnJwz
RRkYJuv1w7QSoaHvg695g/iiRM6BB1xdkSF78w5b/FT6rmVJ07EzM2Y/ezdy8jPxRF31E3ijVJYq
WoIEiO6yxQtMwZUq19Dr1nDZS17q7qCOze9s6wa0Du3Vennxazbc6FpBdMZl41Lz6oFvPCNd4RTY
z9nZPfIZTmNNibIICItJF9jc5gYnbTgumnTxEN03W5V5Umhyq4S+M1v85Ve6xhzZPt3wda/Oex2q
vHhX34wHX79B6l+p83brYsQBBhlVYwnXCepN8mqlFEa3bDR1jXno/ntuecZb7VyyMNST+cj1vJPi
CBcfwYLhDTYqmE/FweOIsRCRVaSZY09EIVm3SoGaFdhPgki2oiXxGBaALzWduW+m8VWDJV/BFrYx
Ew9KIN3bDmO5zWt6u3+mNaF1qBNu9wyjQj/e+psrldMzyXaxpXe9Fey2V1TsT1GJSMUotFbyMf2f
qBtPpv4PO8A7shANiDIkyC3Qsp33jtGgQRlCWz61yZ9gHlWSaDBbsQiCDdelM3pc8HtVzhuvawe6
tSjTZIhyFUDvWDql2GikmGEQrRvsC7najif+e6RSDGwCfBE7sHGZycDZ2BynNAk6iyyFdhUOzOMz
Bvgh9SOqBA3PDqD43WbowGGkqGcyKJZIMHWZ0uQKGSYTdiXrGxf6CPk9vUfcuAzS6ft6fliPkn1N
2/xablYb2i6IS9QbOoItdSkqYV6xjL+1wkWiJAvOkt3F8pk2iOzZhLviPhgSWAVXOGRFGu9OSGtg
y0IpqjkQoDBo7CxB81TV7WuRjVWf/3Xg41c9dr8qEybSOZd4hjRv49mJr9uAjnXG+kMVa5hRnO5F
nwwwxeTdaAj5x9ClngwIMAkXgJnVwHcYhZM+h96dl/Cg5ov5pMf1F2bxczWxxzwoAeJ+uzBRwgUs
GFObW6HorbC//AbzZDNBOIf8QNdF0KiZ9iA+m5GABQX010KNwgNts7fVuujSKTrvLi9FzLFe2PLc
6rd3mywqV6ElNBob9Cj7xlk+HHRHVoF7aSZSzurDd7iTG1aHnypZbPxsVRNq2Ko033k0VnRJEC9V
f/JEPC6OSOIQmvRDH0RRqlVE3LSuuzNMfqeM2yE5/5zN0AWhfjuJhEpCfjz1mo2/aF3q2IfM8zIu
jLeWaS6UReZADSNeSvPWpqCVSZRcWIgV/dR4mN3EDltw13yNZFh3oIwkgr9FaoyzuHN22QEKI1fn
nPRqy/Hhz0tcO5WzCrYt2V62QH+leWAyRxap1J285n4O/H8L/rq8m+TMX8GRYII4qszDk5fVTKE9
GMiNq3znGcV61XXQ4hIKxuN98XoOXFXHpcmEKpc2v1ukSypaHCty0e7v2B1+qQDJyNFUIS+RH2P4
dcwl65tBPkTuTABWMtEHSx9j4XEleo8YZqsjNuiYteudkouGX+ltM08PfIa9nVSb7etmN2iCdCH2
DQnuLswozYPtXLohE82pcrciMEGXPGjwIXC1tet2v/cP42wzSt/1BRIR020YtN3HZAtDVBqzQ6Wr
27p+JsT+zK3evePzqZVimHS4gc0KhIQu5HKjxNrMkuCUJut7MQmYlhOacHTYOpcAsq6+dUVvv876
shm6kvjT4bidLlPQ8YCwzzUACcO1iNEMnC30j4V4X/sONxonpVhIy6onyR3OmQg3KeT9EkjxJ2sR
mU+TydT8FhC7OPgrtSV+YpEKgG0QpPRMqKftZAlVtuO96+CTd4EFlNBKTu6cRLANoGRgeWx3nFlO
gZncOeYvnRaS5nSvpwjj39pYLgypTq/WvPB7bCRYUVegYltyFfmekP3vhS3DKllBYsUgESSW/16G
APTuYD9dK9HcTJAKzALbVcJCiF1MJeJ6xvrYyIOvxTY/4eu833sFHjd9yUiq/fdjBLcYGyRyk+mE
yexIp1QVyU5WFVQLb+wZ9siuuWH5BLL+eK73pi0ciHKfIrH0lNsnxU4tm427j/XVsreIyrM0SgtY
g8Rl0hptzC58QbLJJxFzDqLpL4+X6J7H7OHWC6kG1JHlUmYVyH/KSKfAv24dX+LfQIRzCAORiWMe
qkI6IE8hWjS4pvlQeJCii9FeczAw8zSJTLAyUvQ9PnJ4n86EBJqJhPAE5GAFI2gMFpWTJCQ2z9lr
71p2IGc1YgI0ZEXJSskAZkaGUR+fwxuyt7XiH7RWy57LftCfeshcUGOO0juEr5CgztYRwuzRkLLH
QrFlsHyRR+dfDlLRgDvMNQ4/vmmAFzsPY15Z8HCIcHD6lGWjyjEKfcwL7C89gSbmmwKjr6JuS/Kj
tFJpapnXjGggdB2GK0hfxqSfjzAa0dI5qyNcc+qv0Hv0T/wIst1TJ7AK2Zxwm6+KRnM1Hojx9Ouj
p5RFKMVRAkJAKxz36I7b4cf+mtb9e0ZBvLC0lpA1CvVKO6eJDXWwVYC3hz2M00d8R0+lyJ9SWIgw
eVpmLlQ2wqSP4gkFTSOPaQWdBdlhAZg5V3u21WMfje+2IQS6CKfCn7CWjseDz7Gs+T0XvuQKSn1x
ntdXjMw2RJM06ntvaH6kJnz0j7CB8LlUHW7ZOlGcOhyQxU6SqODNNSW8/iyFGUfXK9EYrN0di9Yr
dzCQNN0g50Xc7SB7OckwQ+b574iCUKiwwW8n7exT4xufK0i8QtgT6wKGdaxAVpwA2P/wCUPUltgD
pXjrZizsoCnjy2MdLheMMMUfZ5LnaM5pcHODqovuAQvx13vju+O4czcq8gma2QtzfaVe+HdEv43O
sZK5Pv6OW7ztkSCYRV00FOsVW/lO5rqFPVPzCjdm0pdPOalZQDz5G9LUc/IXw1v0KeyH7/Iv3b4+
y5TqxKta4CdD4WRaiL9jzv1atKGwTSz04N6nmIvzOxO8uj0+SgVVDmqzDEPEBZ0u9iT9OlCuytco
qWLVO20YTwYh0G2BkpHUQKBzZxaIHGI6yqmXDlHTwnj/bmZJHHw5xiQbOir6cKRVXL9ZOVgjK2F2
B2KS1o5EGpGQJShhAT7+ybBFzwYPQamWYbHgy6YDd0gz8Vj5gUGI5G/MFMEOw/pycMQTtlnytrqI
QvbVMcdt/F3TvK/VXLicM0R4r7fndLlfJVt8nAKca1yZTBfmVU7oCO2COnODqm2So0D1r0c7ZxsK
oQvugrlcZCGd+s+69+UWAW3qlZ5PuGJR8dqKrDn9iV/wHQ8L0ZLlOEYjs1uVe+ynWI/SixIxeBTC
PlJmnKcoT9OBby8jI0gpJ03h9xkkyaYe3+kpjkFTHNaV2CBFjn+6pUjOaKZkS/64ZXIIyfj4uXgX
pKZ3EnfuYE8t8uVKI3tdy7/ww8JU/bMZqRLQSImfOs9/xUIWegHGWvS7tcnnahv3AtKq73VaHo1l
CV5mhL7mvdS3j7MTRHscmvWDbX3TEexWOnDCOn38g/vBLnXrAWgdOju1f5cKU9dj12KS7i/j8oAm
tnNg/0/+RUkB+3KgBZhDMu3QSi7DbdxGzHrkYoHZqdNAwdyxeBVBs9rtsPsPk9D2lUQ2ooVD/Ura
+L3zhmYZgbWy4ZfsCdfxGK1gYYTfaoG0FHuA2Vsd7hKs6MRr7kaMkHcJ8yx0vyw0SGa3tJI+WJBa
05rCIRxmqAxUWlDXF9Tks09J8sTryX1A/JyqqSlOTU65+9Zdv59mJ6zbSCdIUjOvQl3nECmeSB+A
DnbYYSv0D+CChDk0FKMh9zNqcOwptFUKgCfVn+D7qRCTGju1ticptmWm97hQQ7uejYPaS3DlyT11
CH7ADBmbcj17+ktYOWroI0VInyWaUbf7s8OgXQ8ZRdcQ5ZXUPwNZrfNB7Q65wteH95hI+k8nQ+nd
8bGGt6/26uA4PANlULmVu1SsRREgHbxHMQMcwKnfRzgO2/9aeO50IEOEmi0unzZZkkl+LpNZt0Ri
Rev/7JkcICRDALWk7bkNSsglvNQJzs7/w2WfbqhIpD3O079KOxFSzMyUPlWmzDhV8XdHqluEehRc
B2Y2duJZLmZPWsTxUtfoiiDMxAuUvtaCE4NIxtKMC0AKTHEUiUG/6EJVy2XTau5d8BLx8poPyOuc
H795qiIX2Np3PE/xB6CMh5fL9xV2mbokQ2L7V9epAJjWBdGKsk1wRPaW2AeyJsrB5QIdjXqyVK4f
3npqSoDvOK5CkoT63Bz3fRID9NEnDdmjz+i7lLhBifNek1FdtAAava2YwOKOUx/A3NG0YiBr//SY
KE8to4tBWTZaTWWasJ71JfvdteOHKriwLk5K7cjJNZ9fxNdqzfdm/TLn9307mNxdmCxFqOWECFGx
gUzEv9We5Ahbzqd+vF2te6ttXGIEosfbSu5L7eTvtn+31G0jgqK233AKmbhozT3N8bekKT9z7X1q
D+sAXX5MQifDEJ4xGAgMJWTw1epVXi3qCznD1uEAgfHgdpoQ3wZ5XRA8u4oZxKOB8hZ5uwE1ZVPk
woj1QiJAkBX8O/eHwfcnDnbGhJLpnSvnmusXJRytxlzL+BW5WOH5NGuuyvirQ9rP3SHnMThyfzVg
nB5hy29mBs1gVn6GBElfY9N3rTPRmmaYPApPLW9mYlypa2WEVo98QCSrAQlupI7KcRRbg8qI0qRJ
rdqqMn1fpKnVTCZdu6NoCU27lm8Yv3c4PXeI2vcNiw37ON7M8p+/kXrfwSQ+vmwpOwrlzKlNkx7W
fJ5Z/HmJ1+4L8liChK1+jOYwcfBlhv5kb6YE98dYuZVuhIU5NjW4dK4OZR2KIKVcvhvetzlcwTDt
AGXer+ORDZyrJ0FKzVlwOWlldPiDrjGLuoo2aBfFcZqnWlrptx2k5mmgwU5aR8PQmT4uA20DsvRl
ToEF/PbplZ1QlW4IXoQ3RBg1LxS4lOsnij6YRtUNe3V2X+OCkOkdcSBkH8VADMnXSHsxOEq+dx3V
UrQIY9f9KknzHW0FsLz3OEtuC/EVgfp2wVzJxjsCTTtyTkwzHAB86J/TG7frrvk1i+x31qyrAc9c
IQ5zZClnqup6q9fRSPZ44E5AW22m6kG5TT1P45E69+wgLtCYdlSXmg0Eq2sHmDeKMXamHMkfqZGR
f6TucANfclRg9SLOtlTrjVIkMPrOND/hiQ9BVJyl031cq8FOuTIaf9s3c/bS/jeHWfzcrbdlf+Zq
WWvh+8W5iHrRNYjcAc+JR9tiefvJZ8A+jpzwVxWNeYgDLjFmkKUt9PrKix6y0H0/FWeY8WMbIpuq
r4yroB+x0UwQmBd4zmfJ/IIVhjBWINeaNoD2ZjeXm8nfceS75hWX91tx1lLTM2gnGaOu8j2jn661
CaOuWHBG1+6R3TB2ZzQf+/wiPHCUXP/m53hi4BLUVzkVXz4NPXPy6Wgrdk26qHInnG4u9WISNuoo
fwiCx1l8SBeSon3uLlHCgBGPOxxcxyEKWYWnJkVrm3QwvCcSZHC1qtmopoqEdtWgufmph0kRCVG+
e/lLneFUr4u/BZL6i/W12kjtzxNb60erP000oinj1pTZJWmS68wy7VqocesKHW3Im/C+I2KOiO6t
rSjkfvPLkxHK/0foU7ODe0TwxzrAaHKNIcVTFZlEfuY8w1L5+ziMb+iw+BW7gRmmQvySlcpBVSri
dHNfnwHwoc2aqGZRFWbMdwgzfOpxKzrMlgYjoYscxGNYq40CDSMTMisiqy8fj64ZPi7fMuIbWc/c
UkD6DjMP7C36osGRlYXzelxUk4KpXYNiqbJ9oKefY6/VFgR3R8CL65NnN+Nlj8j86N3H8H+hcbeB
aD1U71jBWeGvqYLr03WrU1q+jRB/OU/NpGGPtO4FHRJUaOjAIHwv/ZbiDlJ7TK8LbyOcFuiUpw7t
TDfJ9uaPTz8RnTNye5KnU4r1IeeA0XQvU+f5DUewQdXcF9ULxNa9sONSGWpJbVXvRxUMhtX97wLC
zse2CWa/2WqijTXRf/U7R8ubATjnuJYVDnDhWbuxj6dvCGJDZBo+kgYPVRtbadh31XbFBAeiz4lw
RTKf7aOPc7ylmMuFveIlAvJ9JpPBdnToW3IFRggRbKdDVJwZ2LBZOAVJSM4GxT3pAbklBrI9xRg+
7rcZF9rEe3jMYSr4JEmxErNBvS5GLmtq0KWnHov5iQtjOIRzx6xnqg2Q3mD8gsD5vb+9OIXuF9Ih
uNR8UWDBepxrjolZBZ+yIUsaZE0AwoPxme+/M/ww2hUIku4sFzfwZhNmOS4KHLoJkU9I9J5TwU1I
OqPsb5g2ewzrWGgefIXWPow7P8W+CCUpnWqflaylAVAvK+fjDOnId8ZnlaG2cPC0BTVzwCeqo88W
xDfjBQ1wm8zLNHO754k9Es8V92bSBWMvmdNVWLAaVcoy1n/9T0UxS02nyXuZgWoqS5ytqY+hpJGr
fhjux82OktzoDKof6+abHCR4OzrE4g9az3urBersDHEYrDNllTW/8rIQ27TIE7aTls3Alz9NMuI0
s5We/w9DNw38/AiARcsqFKx+ZI5B4dC0vD5Lyn9ZnxAfcpDcooFF1JlPOe8CvnmOD3SKnzlRxo5B
PBZBTkEw5Aic07kIzU2tfQMYZ7UECD7uC9GNDjrmYPW2uZQZy3ZTb2jj2MpxfbazoUH7EjahlSxk
sjxRBrBm5xx5o6Cdi5V/GYeCY/e0SgeCOPxxZvIUKSLtIHIlovvKFoH/X39tiLpHI/MHndFX6JMh
LI5i0fUpVV5yAwF2qtKV8+OgwjYf0EXnJS8GG6GZin/k+zsYv8RR3exa3me8cuLTHxi/Cm67EB5E
YAxBTIdWulrpNbTp3qbDW+bbDrKG7ZLneujZeOMEHVjGSV4QWktP9+3nr4e0MS6S7SfT2zrO7wXt
1z/wcLD9310DuP2tze+4FKbG43yb8bIMV9rPjM/Zba3CGEmdhyFMK9I1LRBczVPPIQW5AEse61YL
T2sOuUHq6j+lF1w5MOlApSHlr5jdxBs8aAwM59CihwU+Wkr7yMDMRGxBCwnCGnJ5zdwHHZKmkfwN
JT3ENYPBE3ALNAFjpWZDx96QAlcy5BB0pKpw7LRpxO0mkh0sGTCDOp0SsNsuJ0g/dJo3ZozvmFUE
8FKpBHNBqvRoLyZeFuZcQzirKaozkH0VFdGHHBMWiue2YMvHiRcaFtcXxFMLBoCw87YoJKT5zY3R
nHbyoHYputwp670FvoPr8Gxz+OGBnPOFtXIzn7vOLyUSeRMOXZxDvdA8z6jW5/DNkyrVetYurzfd
sZklYJY/atCOAvctPqAAryJA5QCQqb8lH611K69c9fYmLdqzw5hlrM4/QCdjfn25EBsGcPI1gqgm
+0ICgE/lrWAYr5tUgRztG2IhOZ1l4+C7q0MHIQ/xDcjG5xqPIGD0uVfZKybDzyqiPErc26erz2VR
3fyu7MsfNM4WLf12G9jjwIMyvqstZ0fmbIbvqd+uXGKHlMitM6SBIoyMPmAs1cLcIgc+KWPF9IA5
tcMT6hx/n0/k5eQXpWjSCXWiNmNgYVcUKEJQi5GJsm+eRERD20owW3OwHbDKZ3lZWgkW5nKBPuLP
HJXgYdRtcFiwiyk9IEvStvylwymyhMFFhgRCZQRJvzjHsavwy5SMpmOMzxxYDELqZWKM//YLhhUR
oeHDsX50DIWefLNPhXrhZiojA1i9sor/MDzGh4CdBaaqplkcRieGusodRFukVdKh95Q+JlYg3lM0
bEYJPnMUJPAiZuClHBMKs6HRUYEsDQuzEMFeGkBVD7R0Sy1j6BbV2/Cx7Hd9l8NvTMensuHGu0vP
ePJjeUIkyv1H/bizAHq6TUDf0CHwKib82oF4g+ojlahDK/yL7QcEUdW8/5IamyD8jwJoqHxzhcNW
rCNFAQWmYEuwSlmyTeAo+m7btKyasTKSTV0cxfrMyPND2hBYzYtWCx7H2Y0V9yDfl6x8u0GcaTb8
62XqCUCfz1CXzTPqtrmCD5mDnW3F3J67/IEs9su7p9072XOsfjYp8e8eMF1oUYP6q+atACHm4c5w
4bR/41S9r5MSk/sqlvH6FwaqDMdYqNU+QzeyzYiNsaznawcrk2xqQJN/ixetDK3zEilpkXVhm57e
9bnD13smV6VI47q/GJuHBtXXeX/lxDEN/rRnpKxDdkIGjKq4yF5jY5c6zAFyL92kfeI7QOPoAR9S
YknlM0Y2LazfdaQ34jMx7rEkDGK+kEUAQeSIqdTRU4VwdxX/Kp9HZRlEh3YojVFeWQcHiZ+SFOz0
xor/ROClazi/Em1lkHWs2CYBg75LM4e1AZJUKgWGDxXwcNK4CFlCWUgCfkZ3FQUjTpX1uK7sui7L
1tm+gFJwklLcdNoK0rUMjzhx5wvXOoahQPvSqRiYimeQOp7dDziE0RSep6HyXmNXzuDV1HpuBq6O
EmQoEnC6oN2x90nlW7pDItjHjkgwrdemgKkzH3hnMTfVt8I0YtWIddtFp9jVPruKgeOdIJcs4ShY
rYWjevfTo6tzfEqhtPNcQ/J0/YGA+Q/2ntzptrormu50OA8zEdT9DEHHdTXfM/fkc4n3ogo38y5k
EdXUOffs2Hk4Dr3I6icVuvhddYnJyj105yut+e7XO6TrJqYpGBc2N1W6xDbj2t0PO5uhoZlxgaeS
5tXNs8tXK9p4c4kGnVwR1KOgz9rYEELU2qHnsrk9/tIkl9468Uc6R1M+59wgP96pt99WstWo0IGK
JSoOGWBh9fbcXXDUfD9Uu0/49UkSYRJIzqH6anM0DhUk1YoBiBDIfLXUM4t5YzyEXXrS7GS/2LeS
LuuAArDEa7AH5hrznNVQOnrQ0+nenYseSg7uBfQrcY+zgXUdXk9YjK+/xlTdpfYr7YEfbDs9fxpd
7VvarcgUnhhYITa6CYjMHIWSpaC353ljEuBTd8bFmsSxlCFDODb2nV6qr1EEF5IoVABnA16SIAN0
ID7ieCxK6QzdGJrTLaVIus1Wx4/jI7o/Er2cMgdoWMyg8lVONL5tTnxekFdg3D1ebQhqJUblPOaN
2uj4PBK+9FuJq8wta1N9LQYzRlvGvFJqalaKPkRCYiJctcCq2SFCngEipByZaBabDl9Mcekw8YKp
CgNe6hvwh3OSoXxbD1v7SM/D7cks19CJV2EjoEnQ9+HrCOsSmaUmVN3sa9+rGK+AVLdEg0r/E/Zu
VEJhEzcgzeAyq2DAEWUvVUXekjM8qtbH0Rdgfqffc68smY2KlTLOGjhWUHnErCbSPEnwiDH2gtsm
y7nOYavkfGGSfI1acPPJ/mKaXr0fhLe8JD3seCn3a1ku4uUw62YI+oThfIwqJVtGnKIn9s0Wf4Y1
wS5z0lW8ogXFLIxad5SOglZnGmnb02bROaLE0fdHfhZ3pVRxjG+D4wmaJQ9NhKXtE6CtIM25MoS4
gvoxg6x3hjvTFCmAgSE4GTEjhfBaQAFiGUGHpGtuc02/rafJ5018zFy5g49Gnd5LuXIEQ4+FFRWK
vMb3xWWrjJKj1j7oNUhBwktzPAYAr1iIprULIW9+bEmQTdOpBW4m0vz6yFqqbY8PCZUv+kIzUV/2
SWOq59sLFxh8PrnuCL/osSxAWxDkENzwEs9+5DlsCjTtN3JiHKlQopfwBbewUAyu3QMsHP1ZMkfr
8Xl5oUu0uytg33On3biCEdAWG7zVpG9FAI2FnuQztSBz0X8446obWHejSOve+x82Oi911oZ9M/UX
IO2glMCDILe2fRkYEOC5vVvwhzzlqiamBNZaO90nXMtZBF7OcGqnxcO0MurfVj1Nb1iSwbsD/kk+
3PTbWYRzVg62JbQSjnWXBncvDsVpUrDATbTw98d/KjW9GYtHGLYdCZGmZ8YkRtsBEcDglglW8lW6
SWo06bN+M1U203Abaei2T29UPXTTuKu9dOT0SeVc+j8gw3zVqN/CYX3UwZTVn3qJhMUP3pKisYjH
TkUOuhLb8zOU+GGCYGThjoZPLUvjDvwm98am9Me+g7+YM8EqM1Jl6i4b4yWI6dMiuvZx/ZIzg86F
jkx1Ex2+/hj49z8scffzjJ7yDYfxgMAjC/4VU8ID+4tUQFd1uPoVbpEp+2vL7ORYOx28BA3RNkX3
9yNWtbY166kTj5igD0GyoTdvd0RyeUx6nq/6JCOmUB6vPhHPXfNCzlpca2r+NowVEf6Gd4F2yjPh
Bul8yrril9HKp7xKjYxW7l4pQKR9Mi9LHGOPNGw+eiI9IDvb92spHASKtoocmg8zifP3ha91BZDi
MeV2vBq7wuCRdZIepRCYUvp4Yfp+GCtWrFLub/290NFFw8jgzTjURa0Pn6eGlP2vf5phfmLIPNaj
E95P9RS8FItArwC80v35AkLMf/eKnadZdtsvGXcU+ZAeUjbXv6bmMx9/BUQ8ebXupkftPOgfaVWz
shDRdAFjbzrdsxTe+/iDjPorrJt+jNV2DYjEW5Lwm9xm5hi2f74fsMqJQNH8PO96DFoVnMl5itf4
b44tIpEHCITcqdEyOxYCXFeNdBLmZ4Aa3XVLNjpvgWqdLRJCPsx9r1h4t0u3bDdHS1cAUOfzQ+pH
7OVxhtnWk7Au4qpnlHofDhuomkSltDRSHF1Q7rRgrpwHrQ24xZTnwC5Z59ob9THDp9g5O6ktIdl5
MpfUf4xhsJhB9rMPd+gOKdY9gOl2YxhYnCKPu6n7NxlkXJUp9+1szo2K2I558IoCbInau05rSp6u
5ji1Zih5lhVezNpT034MpHpT5ndKMzJGuixNTSR1EAebM9WhDRRKNadTvAbi+0Fj9PKwN/9tEXIV
8iYmhgIyS1QIEhibzsEEurEMXaGI437UcxLbNnpYxtzU4VA33p/ATR85PFsVicWbTg8kJ+5M25qw
6/Ario+3NCPb85XNDuGkzOODGoBnREAiuI0jyYilz18bQ76o6iP3DFUdXSOpt5hQkUT8Y3DarQ4x
P0NkJvVDgqor69tx8L5gv6MRpsqjM94hp1tOPMut88ZOQjaLubGH+doiUPgMOiSMm2mRhssUhukz
FIOfg0wjNIHbfTYrW3lMqZgFsgx3k3Kb75IevWnAdQi2xoCQUMawNsDRMbMMapdSu9WZ48OX0LOt
VoldTNKm53yMCsqx7rHesNc6kfQlYAw8UJXTS74AkJly/jwa26+c1PqhnTUDsRwhvHtnwg4f2zcp
RwfH4vTX4jsBfs2YPETdmScQfp6+gWT7pSosB6rzlZe5aTQb3sZ72AGiiKK2Z8nqyJRXG8+twkjw
Jby0KqgdJ670GuLiTfH2wrHTEWeTUE7Y2XIbCVJ/8BgebTpanM1yDsjmsv/c5up9kqu1rrMyRfJJ
Om0oXQRlukyivxny8phDpkGAlWBjxSVCHps696ydMy10H5NStjG1M/Wg9nrcMS/evFVAEgcRolLA
4HjYYPsWmBOFx9sWlZudhxKvtgfLEQOX9Y9E/K/hnWzDzxlcJbzYqqXTdl2ie0Too3nVptpfTkHQ
qviWdNwLSi6N5tgNRIOXMrBGKGQQ/Twde+fhpKhj6tiFAgdZ7LlcN+HuPRQMSheolyPslprXLxM7
g6tXOpUD/etZg4H55rbXT6fhjVhx2ZRrEku56fNw7LekxXQuLVpcdJYI2+pZv92H+IAFM4A92hxd
ZDEKU/GfpqzjueHtiGNmAlyU8V1x4oesgme9JXZY1PNpDFqrBYTTY1ds89p7SKnkPV6YpK+kBYTX
KSjj0+KzEB+7Ll3tDkZPuuehHvE8W8rTvHa9xv37Wm8UYjHynKuCq3kTGMOYUP940eAvsAI6tmax
W0AQSjZktzlFhu7sf9VAWJQwN9iNgK+AXDDS0g8H3b/R1F/OjBAHhSS1bf2hPCQqnq3QV1QlVDxx
AgQp2YdO5B3zYgajklE205JBl0iDqZeSZPeyQIShJ1zV3wi5oXckL1xIVvZJvqgbTWKJMscQbhxk
opK2o0qFBubkKGlgwRvBCH7GigsU5rt4zCPDFK4K/IlfwxmGy3udzSO7EbjSaLmivatWzl0lwCW9
yK148/FLjKYMNn/QZt3kY5GTm3errxPdCBsJMc4RpsLIG6yH0wRl/7xraxC0F4JrkAOCuAG4oWJz
seiWOuQNXOpf53RLlIie6PRw7hcxrTXs9MdBmbFXosEbblVM4gkZDVo4DjJQ3mMyleVvr89boVn4
e54VAzsjFK7NyXcgPSi7idh/xSnKwym1S6+h5WXOA4HzVm/VjxTjCpOCVu7dnas/3YV1+7bga87r
PN0/fR3QHnGcdGlvUtnyPcOOfwAz/wVhMcJ6ZBFhGRbXwDf8sV1iOqyRjMhn9YC21xFgZxEFQUMh
4GY4BRFYz3Oke2rYOyu3LOs44Xfp91CNklrwsofG+e4em1LIq9AHVvFF0G78c71qwksNjLJYuUcY
v5RsgGdwUTNV772x1mvXCzEo4SlGEq6t70sPoAGjiNZsREWSct8HnsJ9S4su9lnWSNWmadB/vBq+
Mg0Nkkljhex6ApYZL3EZcYjDi8hHs5tNwQ1U3kORM73xBqyJ/6Ad7LeTOetJrR0Mf2VTelN5/dTa
GBxHrLmPJhvcHHxKzqk6o6mStPgUF8H5DyC9RniOCQiXEQd4Pbnao2oX3BoQJ1KQya4F/wjjRD7T
381k7MYemLMFMx8be5dARisMNuF1nYepiUZuY7e6zhw1uXBIy8z+9hdnpTn+/DgQOF0l5goE8YX6
8Mul+OpdGTyyd7LCPaxTk+/8Q4OUQXILO0L8u45kYn+m2WNAYp4H0JtGfFarpdiVOkQo9bHzrm0B
3eMkK4wVZzLec73gzqI2qIBnU/9d1OT9lMCqUAEPkIqh8piFFmy/ZHbb3B7Z3haeU/UoWkChZv01
VyLZuuODD32IFp5CK/Ws/Gs4/p2Zl+7YxDpZ3xfc9KMBX8pxAylTpYl/DRjrjhv2trhj+x/DJsHu
aVSj9lLxF6bLD0ERCF3LmlPO5iz0wPc8FRhVpG//+7HRoxcvk6sGfnOZAvh+0hmIOWWroN3r4ur/
JPUhBbApiHaDFDXj9LTjhJCTD0mIOeL0yrRov15QxIhxtnQT75ejePqCsof24pwWrKn0WdpNUC1w
yYVxs89R3CIe9T0kXt6oOBQgErPziYrwcLBQleFoWct3ag9SSJrm7NaetXvctSYAFemQK7YCsNzk
dCfuuOqz5/s3gw/GlR7Ih/+NlT2SkNKTfZxhTdtGuIFfHN+ZFa4AlJobFTltrXj1ZLPqWmwxxmnQ
eQgFVbO7IAyAcf70KJ34EcpZMYEWrk4/H7ezM5LPZWGWcG13MyjmN7YWRFrPPoM81nULtbpmZ3Ja
eFKOQEFx75D/gRUnWRIHbMWM+p6U4jvnXySLp9DBJQHSE19jy90n4Q88SL43pxIu55iDF+F+spo6
HWTq96m4M6jxbk3yfvkYnKCf0sEPcDdF1VPb9P6Ey0Mlef4qt3C/uwjw4xNhURN7vy7TpHcWh7Ra
ZYt5UmOfaP8lLR/8/jq//jd02j1/BVFOGQlqvcYJq0+R3LaMc+vlB1P1sgYauJNv1pnHa6DLqzd+
tssrInZTW8isN7p5crZSezIpxGzbQX2Zr+hzLrrHflsbeErK2canUWEN4yi99rYLKW5B7y8Myid0
fp//B6c36pBOrp1M3u8Rl23NbOAv5DasTETkeU71FW2rpudqPbaL1r27IDlkatkaEqLjJPDUVx3S
VhE7zeWdO3n4T/8xQFycmNq2u6x3GRW9DqthIxDEncSUPnVhrQC7HW+iNja8U7mU7uDv2kJd+aIO
ITRVLPmqnUYhCoMoh+ZGIbAqqhDAtD9Fo6iW/wYsUxINxRE1ffV51UrdJ2KUbY1/b/dIL3cu3QON
26NyyM6LqJZYYteYk6Se6uo4uoCqx9ZoNWZ9eXMpkdroLWvFhNg8BIS7ZFGKqNv7Bm1uK5ZClMwl
Lc7CzYkpryLqrC12QXu7Fa2sBkiq3mY44Z6twl8CIPkzGEYDNrKmLzlJqpV/HzjX9YoK3puUcZ46
2ykoewxPFeD1GmoFWAJGKoinXXa/r8366N8v0VFeKmzcrNS3DUfduURKOMrMDq0sM+cIybgOSuUe
DBJRgJirc7sxv0bMFCkp+TsZ3tj8RXNdCwdyonYNgr7XO7foSdBP6hQJ36majyrDIPH2cwoj1ISC
0gqSxtAJ+0TeJcXAn4cQEKYrjhe/VlzewgTCOe1yAdr4CQT4Cc0F7PepVnBDvVTovj6o1Z1Ur1yc
cvZ1zywMPuS+ls/QWF2e0oEh8UEzPXjVQ76X4okucwABLpf0g1CnddBvhUXRYPJDoz/mWNcjsL38
Igf5tqJ3WcFxuY6n1qoMY8yaRm8GUKsCxY1qGwjecyhYkeQeqljRSMju/YO0IG1AurqBiXBebuvE
x/YCDNTPumLlo3SOQVwCyrIUe6coAlmhc38yGMeoBygslKoYiq8SUwJ76RKGpZl1VqMXetWXDEVr
AFd904frpoSmSNs9EW3c0HeDrQiiXxhparkVg+Jw5u5Iw2fDUBw55tVLH8XZQJhl7RlE7xUbQx/P
sEW5pqgRIk+kRgm1+mnSFKGN3NrHJnMq4r2BsvmmUo8myUJt1uPdCeIz+0TQBdToTOh+wlYM/KXh
e1UClhpTOq7ialxC98/rWRtk0qfV9Dp8GHjE/2afwD5zkLJKFcS3cExzZRFnVuORrhARVq38kMKH
z6JLIoZ++h81/BUx94ThHkMqjsQ3hb20Cg0FyDGA+LbQUODcA9/7IX1sOBZNu3WcPlFX4+Y7KK9G
aOVpDGZj618PmN00oIe3EIuUEXatxeOurTitxr7q8kvhTyZ5nSfVuBMHkonTwFOyOGq5PyuLbwwP
MKynmVIM98pV65eyZ98EqWBQftDl2B/uY+6Ub8Y1DXvC880/y/C3eAufUxeY2FAECjh/eevKGcoj
be4IOyLGJjBrU980ehOUbEGP5kbp9Ot6z8p4BrB2MqrE5eYVs/68h2fVts/pgfgSoFSIz+Tox9dN
JbWSILdMzyIgjz0WKc4s1pqcoR/AY32ifHcnatX8iDlk3CsxwWfG9jqwcuvh4uxpYOLc5jgnwDxN
zd6RIjjTl4bPak6doCvypq4H4P6zT11SdEUyo8CAkbuGfE0i+d/MMw6TD5HfO9xteSEMwC48uVli
WcpDu0b9CsBbCZca2Nq5dzMSqnX2OHQXfGW5sBg/822iphgzpQ5s5WefS4z+H3EqR4L8ZD8JF73W
H9vdugONMGHHcrmI6XdRhlDAezPA3BIUevAUzn1jS1qYnH/QntO1bcp4X4aqJfHQpjl3Z22XvVf1
kv2iCz+0gIY1J+qwlnH6tkdpxpb0fWCzR2bpMIJsdXFbqDi2iPwxXxPikOWsLHM+xmv/bq5hefUY
ovGehGOyENdlX4l6Fn8Uya06EHtVwzgufHa0BN77Yea1XedKxIQYhJ6ZFt7Ub0J+N0nZg9n+lJPN
G9/Jbwg0IcEwm9qUYy1L2IWIDQs3z0Xr4gAZQpfiT91fW9CdqHyPbivmcguAUfZTJvqvutd21yQT
XqROFcqaiKUYrEkB4HRkFIwjnnLeGHLag7WuZJPclq9ey/UCAzUOHcORYmU7CmUEtkKI9S5c054C
VSZ4jcHc0isqRUH7xt4A1uQp2HkMww9tyMi4caMxlbh+rXlW/uqAnx9oXOtrQAa8iIsY7n3PH94Q
r1SooQFvUpBfCLoVoCBsDiylRlhbGDTCWctn2E9rJkQQ/VFlZOwTAubvYBS5Jaofo+bdGYtsYMhK
6+Fhgd3mkB3Kf6cqDCX2XrYPH+MxmgJadoVvZP+E3utA3CzVXLjJzzTf+H4yLAHrt+C+QAOhULfF
lcgBgy1ItkkFVJR3MfK/PI92T8BVvLkJqwDR+bGMGk/LGrx24vE0SJqTJLaBNWV5NepbKsHMNKEX
QSvKXdNyS5SBR38WC76/X+xBhcXvAcV2yQ2bEqUsguqZA+lgQ7kod/0kL9W0rWi2F3Sz/ES5Eo3L
NoAnbzMH/zAjRuMg77oTXZdFIF7Dcke7Cb4hb2yiCL26gIBmQ/CWc06VNbjw4iPce5wN4LlsDqbw
yVod5fQqNqUQorJlYhWIBQmdI5HLWnilTe3VEuEy2JRd6vB/mbTzeK0kPVmk6ifJGwi0z1Kng9AC
xVz0Eq9YKFaL6jDsNUoWcJX9balmkm7jDJ4ccG9P22box9pkZI+/Bnc85h5KihofrDRLQgMzAtzD
DoCoGodRqo//WB/+G15KmjVnFs9GuLjM8emfNPJsXj6A99AeKM6hCSakTLa9ut7Oj3l59NwlCqlJ
HshYFNb1wY0/WzcivNGYXtn4mPJW85QYg3A9XOCa81T4mzb3xvLp3qwFd6GVehcCPR3yGmnsnqI8
NoiYLgwCLuA1HvfFMXZkk+iXP5xooAQBZoMhJIQmaksasOXOiQxHHfMgisgoNLHdHMq7dc92Iamn
jS7dohIen/0yT1zz7RT7I+P1Zds98MmaBYQTvgqw2h+Yzuex6sojYCAuc3KrA+zdHwqNK8vntw+7
l1xHahRsWF+PeB3rNfGXRruA4QBGwgP46TubOQCjCfaxIXlIbScvv3IgZaqviLRMSZku7dyPWTYr
wQYoFA1gLhyyN5upOH0AID+fZEeQUAtPiOTpI6/+qfdy9JPGum7fL709e0gSTsiEF5Qhyb22Pfn0
7QW3j8RYlCMdJWh/ejfa8z2oJhO7WxwtKflUwlD+o3TkdSFwdCmV/T2ONmEQBF84kxjzWWzkagJv
4lGHO+IL7UX9Oe9/yc1+fnPUw0dgyd4D0SCrhSCYUZRvRwQ8ivRz9VExp6hCsSrtn+Honkfz5MkU
KYPpXJnkzad4xyjzY0rbn10kPP9QH+tBT4o5THCUDzVOcPRiWHP4nkV9y1dyTmXabHkvSOfv13Y4
2GZQc1+xwjkCMih/9LFreQ9ompMdqHRbmo5IHsWNNOjZsO+Udf1gc7xaQgqoa2V2DgHCeCHD/1nI
A2NNvdAg096DO99Uz3PbC7Kwh43cG2E4LETmlATOAfMK5cWBeYxJIpUCWGxDoBFv5A3PcGB1eQrG
1DOT+s9RxxVGMcd7DuVIPY3nUmMQG3DlpNzlxPDNbtlrpN/EVLemY5zXpuDp+hBvExXLVT4c07oE
ZpDy4evtyo1doGIlLjxwZRXO1I90dU/8LWXsM3+d9ljGLVjk3+pmJat4o0h0fZ+rM6LGXHjL7mdc
MApScytDQfs0PpBXb196Eov1uv4WRZhA2vGxHkYS1kqhfyJAf9UZv9fE1mIibJOboArpc8txxNVK
NAVkHhtrZESAgfgaWxFGuu+mEU5Ck5usNojAt5cioJ4tWlIYXhWo/uJ0jV30PvRSXvk7dS1MRn8g
YFvRAwSnhM0h7eOkral4tRHaBDwGgmyX66hZumSFDarFymOSjWreqL3lbAD94u0OqTbIo2w6E8Km
tAEI4MgxdjuRr1MV92jPd5oBr7MELYjxkXf77yShZB/FPWGMD4bCq+LLXj+FI5JUhQE1slXHIa5g
eQ6GSnzQMD6hstQdvXcTLWLBOPwM9A2omZfjpYoZ+TtJlgC88qIItyHayUj6EFcHxYKvUljyFB9o
Arpicnepn5BxHEs7fpIQxKtHIS9jZTYT7Vaa0S+j982Xds4eTgMQ0P4ZENog/VMd67s7nalNUaek
r9aG2sqG1AL3o1x4Jcx07a5DpMvgjQz1P6RZYuPqITLn7NCutKQG1jFCxPNmqdpIhV6oPciRoDTG
hz53FP08gUb7YO9iheS7orjDMv6cQryvMuiAAsk0XtTuoGZ99H5+pzdAMJOGHwL20GHKJmViSiXf
AJbio6r/KK0UsEe3xacUKEEoGR0cD2hvAS1UR3uf5w9Ddy6yQ3DDZwxSjsYLB2+v9DvJvOSQbcx4
EEdnEKHVl4qqwdeyYMtF/p0lcPLwcnXtu1k8liCppJXt6vFq74bq4QL4IommXoOT/8DbBqqBLt9B
yPVc2mdG3/u3DsUhjTYOJ3tSrOo8N8xpMrYoY+5uV2xXIN4+lSSjNLVIDyaQHeZAVspxI+T1VK+j
F+ARJDRhEaTQHh9H8yUWtcpWFpHRAjbh18I2R4b9TDmGD9bBPJY2m8BnQ2qJVBUj4JQyGjsctK7K
Su4bnp23QAx+WE09bDaIX3to4jbt7BOxZjTkvG70FusKQV55ZV3oQf4Nccm1oe2uMcnKtQK3zQ4l
6S03qECsR3+j8pvWwp5NNJjXvmIwQwicMuFeayAAt5ePfPuPJN4Swl9IW9uyR33qjd8EMrrR62CA
dysu+9FRlyf3vXlvbGGwQajy23rlmuTMahKE75NZJONyrQXbpGro5OWltOcjqHClfJmqpV9V1lXc
S5EhUOS80uJogF+KI3R42Cxl76pCHS9Uek3uNxJnrkR1Mp+1JkSegm0YbPAAd6rbiyyQPL/tweeV
44AhI2eFQNatQTdENKYgrY4N4F1PQemJpS+e2wgZOD6vjDWv/Nbw/Cy8IT7gQli9HGsLTfGAPACP
sbVLIj/mssRG3wZFB6wBxCBKHtyhqlvyTqV5PSjkvTeP7M6dHofBYJMFG1w86NkbEa5IupMY6d+4
V2hIsZTxeIzqesM6w9IdTmaV0wevytIOiZ0YguGpH3JB9sO94mUqavLbrjOOo43ANgdSiKTH3Ctf
Bma8bj7BDNq7Fn7aMc23a2xd6aOUxO3+TO0of4mvvMYi0leD9aoNSW8BqqjU/e6aZND0r2i3Nd/4
a5vp88zL54iz/K2UUgSgb+iS1j3zTo3wupdfeqQKjN09k1nlLre8bnb7X6xQhlmty26ZeF48WQAr
LUdka9fs/iJNf9tWS9z0XXiMBrm24PiILmHfKYCdxqMuu+I+gyxSZMrQt/nduuMwLNCv+jlAhaKX
Euk19jBKtC+s9Py9vI2uw75Y004ChXFwBMucSNm2b4r4RWWs6c73NJocx7ObzmuZUMl2nUSndFnI
woymaYrdz6KkUzhXcoSjlzcKSv9ZE6rLKxgT3mHEVkEhOlRSQi3IBtvvmDzPoi/wrHMaIVGCji7+
2ZrBhfxjBKwC6BQNW2BuzK2reI8HXLzi2GSWVsJljUnbDksIa3laSbERtqP/caxrMpENsvX3IOOX
VWba3/qbBX2rhm7IC7WJAsZle6N0gqr3uk/QJCJDOgAkmvm+UNu/kMOxnH32TSHE4eIjEi4HtlDc
odTRJSSH8mMT/4ZTjxhjbUd8nFaEVnAUDw0tAaJc4iVnETkLqiVdxT5cvfKXYzvYSfwT35Uy4VDF
+CQXSB0CSc501NEV0lrcAqu+XipVfOaAF4AsWdBBiMxXaTIgc4X67F/kEAnWG4pzLlh0wL1gPhQ9
+Kj2uNZRXge7Izg7Nu4+6v8ePgixjOEw3zmLO9bBQVVg7A/HYAt4bpwKnRBBM/IQqJyn8V4H0D3O
6NhHWhVTEO5LliDMWQrgjC1ZoRV7TVpEP2twy9run2Cj0jm0uJJIL4cuyKfKSkVKWGpMmN7uw2Af
iJEv8yrw3TPFL5/r9LBVNrXCmELj0EcVEpMf62RtHkZ89k49eGjVaO8JnuM1k3XK5l765EmRQeJJ
uDCxyx+AHV8WvwztvmAhZLNwswAX5GzShwqcut/+VdoBVQg42jH8JZLH1gzcxmaMkmtT5QkYItLr
XauVO7kTcBB0K69XORe6q9ulV7UAxe1qY7TPVd4njuI1QuaHI+2rZTCEUxQAYW1r9ar9pMdjaWfe
LOtCC9zdYd0YRR6tjxG9RBKGkwGUfSRCvVt2E0sXQe3j8jJCJlb7SOERz+XVtVu/uuvg7UuwFaGE
Dh2y32MzlLy5TiWyiSDVTzAFsm1UokW0CcnUIbbKbxpMiiTc48k7XiRsxQNzHjDvzJm6Kwkw6760
RafrhW6rQQGRhAikFEzHmki6Aox1ZR431riCUk0zcWaYCK5e+rijEvbQtQ6qaIh0Y6bNPOL6s0Hu
COOX1Hx67ZFoEVSEOa8LHc5CU3AQqe6iCpjah2cAoXRxP4naVgBFZ5Wg/QZfyXjBikC9SxOqCnAA
h0bcUTvbm16wGYIOoq+NqRmzE0Bgs7ovW684OdRRoPAe2OZCrcKMUVopETHc2hOWqGGAGJjz6n/g
FF35JG1BrBsL4rkNXxLeu/3O7JCrS3Qt3ICUcxPfqY8mcphTEBzbKSRrVNa0kyUDNQhhZ1J3cJB9
+fORc+Egqk2I9d6aoHPUpqzi/+Th9B8DyQq40hNrzSDfMHSTjBPoxHaGNmvIW4nPzc7E8a3tZQsR
NK/Mtd1lplPUdIaxYrH7aWFYRGH65z6hMsqfBhzGCTwpCSQSlMNinBZvpRWGT4hYGHRUVQjowtKh
Aq/YS8W2TORAhmP2oDGaci37+DUaBcoiAkUHWH97c41BoZX+5ZEyUkvqlyiDA8uUtkg0OEsyTFHe
yAEZR8dROC/zIV4byF+LtJMg3aqQC/yI9aAdVTUXVVJW+ggEaBYIOFBcfQpx/4soaXzARI3Zg3p1
elqT4aPKwW/7mNb2vo6V76pmGDRFJQLLQdyCpX91HZHh3XdCBVgz5Z8lYGYjyqdS4Su0YPrOPce6
R9iBJdjMFSiZRsm1sKK3pEdyUSrzhN7AGqTTtQ8n6yxIoDSO64Vk9UGsLlYrvHuaG7u00kwoRUSg
j3KC8YuZIozm3wjSgmBincIZSXoewAOmOjS4bq17yBCrY1A4g2MVmepcF0hgNUeeqUu8nxZ/UraJ
PA5GfWxolureMKl6vfLJvBiCN22T0kkdCPZwjUJibbi8Mv8cYfcrfsHarQt6pP1uBuDT4nUctNvq
pSW/EYIYL6RPMWdwpiQs1HekvRy3R44WwxY99v92P8ui5v+kevu32s2k4jk4OauOD1ErjbNIRm5q
MdfTs1h1K7A9a6PybK53omh7b+8Wj1CjMRbIRshWAyDorAaG09AYI+BbIqcPMHUvMbzKZc2+ajI4
Qmgtg8zaFQFLDmoUz1jLskBb02C6r8QCYgs5TkSMpYINkK9LBayJK0U/eot4x2vmkXhjDNfg+YJo
PIi/dFBh9P6UnSCmvJ81kEchojtfXolwCsJmuhoYUqYf9B8Halyq5MsM/NxTG8kA7Q+IulTs/L3G
AWcLblysNUF+AHNfvIZ6qaXpa0vnY72fhpWJvlGDiCwumXlgkOr2eloXW6TPtJZaXc/hzQ/+R4tI
3H9XQhtX9YP0KH/Own7XDtTCYSNSn/jmH9+q3b29Q8Yd6ogHwpX0lVlCUDoAkrvqYU7MC70ocxFG
9VWmraHY40BMFt8XQ0v9iv/lMmuPqo9HEQEOgxsZDpQ+k3U+K022prq/SgI2kkfqrr70KJemYVNk
6A79akuHp9xucuQ5O+2ZyrmKdYbR6vI9Jlh7VpBe6uWHh5oXme7Jhi3qITJNMkCKb4Lt5zwlMlCF
qPpjALAh01k8URQQBZsLlFRtPRELRbf8leVJgpxabV0uABJ+Yhadv0p5yvkBZM4lHPctnxj4+uHQ
1VS8vMNq4fO8/mMCeE4mygacQQf+FhuotYSxWNq2rdz0kr+7ufus6MgGTw9IcQgftSS9PFomBsNp
gEWj0rU5AsTnwpJvb+UM7zPMhWWHdWN0rK2eEUppFqMvDuugn7GDJGU2Pg4IG50T6rnS2b/95PEf
fgMMeZ4zfYkPg1SH1eJDO+5fzQ0LDUvTklOSduu/X4vWJ9ljAkf+THqalXLhWGl3WKxb0fqRLg94
KVZ8yf/YQqQWMlsDwV2BPw+0Xtlpgb3UaZ4WLNifLmlqiZwEN92lFOXveDdPsGSKq7X+dwWgO5Kv
miS/P8qz2l4kLvq+KQlqNgJFfN+24cpeKQLUjjxBwfXRR4MEy27maD8vuQVU1vBah4BgaSBMgCSE
GBYzC5uxil9Rmzt0XDvPQSVOLUh1ogRuqZ3I03F0c5haH4iVFuFCeoNWA72rbhxhVEN+Slr3mz60
jWElmvPU8S9PVQYZlthatAfn8gWl+iaz3UVvDM1mEnyS9CCj/QTt+iFc+YFOXGa63TRkxANTPvMv
QHeJ4nHcc0AJYkDL9qhMySjKLvSFZKq/N5atlt7o7HKV51N/kISKgDM1p+eYN+9A//JuGP8h5MfX
6tjEiE8PLqxIJoEYCbnc1c/361Ld7gcQOUI9jQ1kaBRO4+TnqrnDxpNf46gpjc7BveV13D118USX
0uP0iwXOISrHdaWCx+UlXwan53u4JMoRtWT/UMOlXfM0G+G83YgKPPVNJoRDf2fsvw6AF5l0M/u8
npS++PBThpms3+rCYQIHQFrySGEUwT7GCRV2jE/a94IQHXXB2J7xrCF+sutCNyAjHmMzbKOikf3L
4tFv+X9q/K7hv28pMBFk3X/jWU2VqEKmDyYg8LK8u2tXDtymevS3KkcLXA1TKZSR4GVd0kDF2pZt
3Psh5k+R/cUKUU096fY39GZ/F3wy0hGr3AxaHKAj+22GxbFix6XfE9zYzv3wsMxGEzEjhsu7VVR0
PYRkN7Q2Lqn3iqRO4ZoE2lf5ERHtmu14co3ppqxIzIt2cLTCKUBmMQf5qBG2CUZEZjSlfFxwgW+4
04PPRJOyDYAgWMbxmGubRIP8RmYpImtIOHBHpKh7PrfZvbDb0LywzijGGhaOnMmdhiAubhMDCJHi
c9UIAe/BycV4OY18EU7Dlaf2htta1ENh+QBArK4CnNbxisHSluKfp95gGREs4GiDUzG855c3r/LB
DzGF1QO8259PgYyVCvK9eR05sZV2RwnPPv+P59TMWQwyW0xGefpYx5O26bPJD1KtnuwF8uTTFcR3
nrfM4nve6u0OB1DkDpBOCwqUjxV/nImzpTjLzWVjOcKU8qTvXSU9WZ69u3Kw+NGDdpCiRz1Ybdei
LInRg0tuGXEvZtscdvRjxPzb6ryE5E1p1dSfBxWGtk2qNUObVf0zfNHQC+omvIbs6YiiTsh5I1xw
Gg4az9k5cznlfZ821W0DpQmUvEMs/q7gTf4vyTDZhctJ/JnAKLbK35qEZOUTwC6ZexWwZMFCDIs4
bmU6LP0Zekr+ZHvU069nGNP1FJZtQh82EbEAgb64uelzByui6jgjjNOIznYEFOutEUAtfYtaaE+7
sw643KZZVmW1uQZIWj2LTZC+orlvb5cO8wYRj8SrLRRfDXkVvTebUauK5cbhgSEiyM0SIg5RCp5d
7MxxRqcxfM159FUx0rwJ0tEUHUTHXFzkeb/nGfXChZ100WINOVUL/a0bz4k5A2yuZq8EHAfGCNI7
YDGwnYEwBJm5HZh1tZKJyEplOfvSJbQClGRYXP9lg5CAs+rhzT1vkXnNArl+b8Zgpvkaqo+CjyLi
vXEHCg8ddbNXJaXeQ7X5I4yL5zCGtLoZ6inYFiFgXZVHfJkfPgJw9chQde3AHY5ZYBnxDgTPuMVG
5uifE26SzflA4s8ODO6yRwiAYLj1LxN7AitRR+0HeFaw4k1a42SdMuac/lBYud9NRLb4IO1Iwgqb
aT6FAI24jdKIw5SXfCcg6BlsYLu94YocpIIywENDlGd64xNyq2lCIFvntJMm9Je0Eni/v4aEpzkI
WC59dcWJk64nsIwYPWKVlVyIJqjWywfGX65rWooa9P4JlyaBVEdAALQdkzE8JZNBAOsOlPpkhMO7
iQosg/I8GROAfIwVZVPiIx8xD2CxAISBsd35rhFiYn4yegb6o/abB1H6TPeFuVQbBU27QL6cImJi
k3ShZjvr5SRdZJ1F28O6yUqYquJzJ2Rs1EJQeILFOnyo2PTdgVANnQ/ca35ufMmUZKAgDIQIH1Ci
zgSluHqes9IGU8naNbtiyZoa+j362v5/lzLrfsakt4rT7Brj42XH7aRQrp/wrwvoWrJRaNishNE1
whtJXZZhqVMZ8BQaJtxyNS5LVwqq6McbcBD5fee/U/fF/mlu7R3nJQ06sujPsaGGtQJT2HImFf75
jwyrCJ70fFN7Wobe3gfk2IfxmL1NJ3SKalUfhRp1+oPFp+EEo8S5eSMV03l3L8tvHDvpfyG0tyXK
/vH5JOk+s1LU4Jl8yW/PAeX/Ro/NO1akc3e8K11g8PbPbPP0aJI+RkHAMGI3PXhAw5mPyuhfla+g
tfWaJW7RfhbbPtPBbwUlPIj5VAtfI76J1RGPIA+oUHSbKaPdkwkFISeEB51G12B0XHHlv2CdjxzJ
cBYCU81r+O5FIIpFI0aKip2JkJWqRqI9pPcqFRM3dgW3CuDcMq0BbOwbLDGkhMUUwJsW5ZM0DUw8
7e23fKoUOO+wBR3oA3iUF0eVgjQP9aPCBiHlzCY56p9itkRk1xbjlj63YBVCoCRwSmNIEOlsmtjm
BAuz8DlvoRsSj8TYNcFy5B7AFNW35XqYVZ+xgiMvH8e4OyimU2880AfbNPDA3imQ8YC7Ae9pbrx/
Ms2cGr4kd+0tbyEhmj2fMr1Oxbd81KVxOvRsRJJn9Mh3JwseIRiSvyIdH9TeXa7cS9sl19B+gDkZ
u0pObSArrrPPyf2v+5BlY59CH/5qmSaVfk+NrFMrxvpcPu6yQJgRQPYJxSscZLCUsLdSOKtCc3Ef
7chBOuQMNMaLxWjmd5m13kuRaU2kuequ+WPm66aMIiw6NCFo4uMUMOyoGJyx2HYH+Hg/4QaGtWyf
jy/YPF7RQNbvbQknE00zr+43PMGXLAfuM4zbfMk/KjL6Ul8Yh/oP7PKujFrgo/CFUo4LqJkop2p+
tRgdgpd1T+z1BvZ1ZSNE4BLFCkfsym0Y5i3fzQ+w6xAj4qgw7hrPSqO2sU/AgPdoQ+HvDurbVa0Z
uqlcrNNigc9BE/QUrpKIStZPC/HhgJ4DHo5V4yGNVTjbm09bNWhRLP069PJxvTDtBkqVVJ/jzriL
yu1rLv6VohqSQgjEy8H8bl7abJxOtlRfTq45iLsX4puGD2B4JhQrchCv6XEi3wd7UgPlGeJwAVPp
bT31pH2XQ2dgqg3VbhSdR57zY8imFC92qW3C+nNR3MKBbn9isNcFCOatBe4r27T1PbIOsSGGxidR
B1i5vgc8UAdFcQpg53MEraxEBhVROn6cpbN/RsgJBvsJW2nynxkMM3CGSozuMV7mCVLb3wFgDfNI
ktX+YXyj6N+T4/M1Pxlfddn1ttbptJgg2Dp8Xi4lE2Zj5jWRaKsNHwQCkNemf54Qjtm0WX4xoD+V
8+8SeF+zEBIOsppEUZ9NzoePU/wHe/dZG7pMKRiSSWyYtC4QTIONKU2f4NQjKNG7jPgOzdw/zMUw
KsL36smYi3AQu7L4lUD71hcIrXEQAJqvJROkEAEAYOmWOXeYAEDyZcXjO4flA0eBdIqH3IYBd4Lc
4C1ZOe9ze/dm+ZkToBpYDTMRmb4oZKjCGsOenpH0f8/1NiON8lt7Ec9aP71miWePSIcRMLEAvmvF
mAWagtyUxpq3krzvKBIlWPpPqUMZ3IfnuTKmvApHyEsk3yQtavbN3WlmCm/rfxTOmhmgeG3LS5U2
+lBPrQ/63dccOA+XsGkhX5qnGrYl6f//Xek4gcr5rrzruSOJxv0fATN9s+BaZI9PvJXCKcga5xE/
NyAUvGZUFaFSkKxF1cIX4vUM2kDnis4qiLHluKAPA+7Y9rodVICl4C++LVxogeGK2fcMn0Ff8CT8
ICPUKZkj1FeLOzb9YWgU4PNwT4fU7E3NStgjKLFLsiwAfMtb6Uf1jnt73AnIymhhD1+CnPHfjhzy
2fNQKMdrmuSUBOZB0cr5EdtC5jaUBMZRqmWuUl68+Bpd4wFvBS1+/rc5WMWG5MAmuUQg4KevwXqi
dgIESXZl2+ujJbEBMhG0fm32hqsiniJwEoL8sA0IBLoPQVsyPgclZpcL90xSk3p7dswCLeZav+LS
tbt9l7bUywHz11lqvV2ZO2sXbtNu7Pi6L0BAOF+KMS7OIJINLgYhC3A+YywDOEXbcK2WCSOUitnn
NkVKj/BB+DklDfXKSS9K+wEfwJjA5/FoFCzYu0k8lsHl5kZKX2zeL7WbdYDY0nRbNTiMO9iYNSOU
QR+Em8SZ8zgjv92zhG0icyGhKUYezZd5YAC8+GFYRNVwO5XrTLBDM4QZ7656mMX/cDjzsEe9QaJP
jCJJcu7EQCTUReAXcLpxnzkRnN4kgEAj3ghF9YByOM7ZbeIKr0++dhQmWX59RQOaEQNdl+PDlvCd
5k9BOQtWVaLKSNTBYXTE1FZmk0Q73bRtag50j/9qsheq3DzgNmGfO3xTplBK3BqgnrLW3BIJ6b1a
ImzY2a3b9/+qBjls0FpH8Fv8DJjJoYVv4luApI7a77sa/HTHqIffRwXWD+gDd2CJe/ghMzXgsl1n
7V6hLWhXDIT8OkZbnH3tkCmzLveMch/AxEZmofvre/wWYXjnSxQ2EGNuUNj5bu1hfHcuhBB+8AD7
EUVIAij7s6F3OaWMI1nmS/ujkgJdMF0KNhO3sWDxhWtdzb+Q1eDx0UCdSSZgKtckCRaDIHYlKxAU
yo+fK/SEaadJ1c7nZ2WyKbHvqyO90bw8kmZxvFwJja4ZxGnKfi/TJn4GsHVG//bFUer0Vy9LBSlU
GOJZzmhN4fKM24OqPz4Dhk4DutgScewPAFrAUc9J/CQGqJUmmvaDO9KRVAsvCBdKbELmt1R6oAcl
F8BRn6NNinvEUGfR6/NZJKQB08YYu5us6ygNGXZNof65b2ujRg8Hw3+EZJkxWx1jGa3GhV33VTuJ
kiJFMHBMWzUfB8Kuj1MKeBr9fyX49NmgR1i4LCeQkWiUHoxSeFOyd+ceGbwqnTglwSbvSpCdb7s5
RAMU77USIIXaIAvcBDwUyo1VHIHEkQMqi5dfCqZoYiFZ1y0i+KR/+8Dj7/3xoeAj4FmK/MPN48QD
0GEjD1m6lifNhJYI6rUTbF9/CuFajYBCRy3UVk9+XWAUOWjQIB72KqjPRPTJNIo9EEAon++XfLpy
f4WThUNt6qGE4xV+G1DIHUijLG2H7z0eL2b8wINBzZvNpNVkqP23gafqrdNpLYP0lET77tzKchNb
EyUP5fMYn4lRjRpbOiEy8Z6mKnsvHk5mUqz3dcmeRll164HudU1AOYoE2Vx4emL3qU2f+NNZLZuW
Um1EDkL2desH0u/K7ZerhgfO/w9+uDBUNRFyle+cyoG2JFmxmcte8SevnVSFKaDXS/amzmFlGNQW
0VGwIQWcnxQH0CWwG6zV+kXk5CNgKpYTreW9ukGsMAfTOTthK3uU/qs0CrF8JCEnj07epaUKoo+3
aE7HymVhgpamuh8gYW45oCRZJsrSNAWN/UgdPWJsWmTNifcsM+PbS6s0qS5YCk1zUWwo8ovIL+Oe
BP0BLDBpXJVWu2fiSuyHrjDTtYfaWmjJ9Y8H/NqfYaD26ktROuhFT4CmGC4wyCSxWUmr3/EYJsdZ
FzoWl0qUYaDT0UCZlHizzJybqWYYnX4F36FZZNYIXUGTA2NvvYOq5FFLAa9lq2t1PeGgOMZGYmzF
Hkaw4sk1nIm10FQEBsSafT0oXkMBdrSR10qfGQ0wGdNhTQo87rQEcoc8d8Wl88ccYo18qs9Fqa8v
Po7C1LfzLUmbCvhUAwmTknsl5jL8/wg1TzUrP4yuVRe1U+3yvJXqg/tYbl94QxXv9bzQ8PyONNer
8revsNvBFmjgNP5IYFyTVgBN6IHWSeBMhGZFunspRWTF7Tn8n4+G4RdLyRx84k72kDzUmDy3ApwE
SQbMTE5FdBBg3jQIPGi/CaxgzYR9yxfN6GWLiB7DFwBApd0YP9ESwhcHeSE3rGslpVYfGEyYtspH
ijjZ3mljlQW3rSam1rwxupFOABDJydpi9Rndh6vtkWjTo2LncHFViyVK6yObNuMN/hqtahx9j4Ar
+2fh2LZ5bdiy5a6JW0/bt4knfz/eZTBKCXL52yuMxJGnjOtTH9FIZ6LBxQwb10c83XGAeX6odeQd
mtADSapfuoaTw+VaQl4EtUETRT0zIC3O78+YcV/U74S6HyI1TUJGsEGoGAMP6WbiYfjxQ25QRlky
FPhSI2DfjHxStfRE3c+gGEVf2Twdr0VONDfYvVa5SruQr7PH2k85uVuRBP4XH9hfm0yeDvD7vJ2S
Voz7dro2hxYs+uuXUoMvACcAlf8R6CSnwjDFVBV3IsuHNuDJD58Mt7tjSCgtGgLKn5j24m5PlIkY
eIkNHVhuj102dzruv+6CZ7aVwjEOuO7UPAOtzW4FnBL0dafigBOaDhXkePQ9JXNXgq4TEm4q7OOE
hLh59aDn6O1dzvdPs6nNN3fNsBNSXMqd+YrOl13MP0QW46FScXUWl8J31N6HiCkOu6wXVAdRFnTx
erP+0jtl3wo2muhgdiRh0z+ain9qwHiysUXN4NyjBo7WcRKV/7nXRViHqyufqTk2QDAJyb6giEAc
Zds+DxLVyfUqtF8fF2xtEYDJxqeb47bbGoodSvPi7zxVyJWm0qc7sv71j7HwjZhkhttchWeJNGjp
HZGiE22R9lavH6RJDk//XJERTtMPK40527v2q0hGikCqXT72Sj7d8RcTwON+FQNByeGa58dhlNew
D+Vvuwqb9URvdLKz4Lv8EAw9mLDOKIcrcz46d3Syi2Jdo5RerVmU/PJLDny9LFqNq+m2u343o1i/
HliD27iC28eeqpKWc+ETya6BaR/bjGBEZdiRBRDelNPWnXpAwQv6R23ouyban2bsrTkRkMrVkZ8y
48Hjjakh5iunqxIjKJvRfGOzDa8/Izy0JNMbIVod8LBQO4Pfonj5mK5rtREXjbxcsGpFvoo/IazF
f0YXG3hbfyUe7vA/qpYKESWgecZP++324lzYkZHrLqbZ/e6i6lesXaYdVfxwK7bxkA26HNc3Pr99
SIF2GpZpRltOcLwr+wHBYxgD168mhfD6uDeCSExz4o4sWtKigX0ElCiAvMS/QAoaz8+glo+c98b0
TQ9huQue3CuxGf75qGPHgSDOXPPmOecvvC5p4k7J92sewb750ghkqaW/XrRyBe1XB6k/Vmv1GF1+
yGwLJ7LvE7Xebupyn5vaksgdXRFMlPhQI9QOuw4wW8knr6nEQrF3SA9LtD8w5zaLnkS6Grms1GDj
hLfn18UhLj6/0UQt+NbDeaU+bdEfhfRgEWQW+HJ0TyGs3BGF33pDoMEYqYgw3f+ydehu18QKnIeS
Of/SMsE9dkFdcXGGQNRqXcm9kGgKLU5WBt5Tc3LjQufkkycdrXZAN1MsV2prmg3uMBfHF+z5VhGB
haGnMm7JcYYGwCSBT9mxx/BNsC4pIfSL0Eeylemh8WLJ99K5NI6ga+eCTw8g+puJIDYFQWcdC055
pzv02Zv+jHowyFnqM8s4AegGThPvU2LqWxU3BexBYcwv9tlMYOpZgV1u9s4mknFYRkg6uDUcvoB2
Z0k7QGwYuSL+rSNEhdqHMv0Yg8iidarLNvOMijovMUoKyvz3+nk7XHZp0iEV8Yhf1D48vBicG7xY
lM9c5gK81NmkNNpQ/5ez1QcddpppN9sorg2+oWcJKWUHN0Y+6F+CYxWRou9IHGzCfRp3RMTpsbsz
Fj9GH90zHBpsgTC3ZLWhQsZwurQu+gl1RnjMVggEk8QN+9CTRUkKMHr8tzVC93PizLYziShPKi02
xiuQ/Itg+A6CfjeCFqhV7XyMnFBX16rdy50uujcAH6WEMLPFOInqlvNCUCon5L/sTXShPyXdaorQ
riypVj2EzWTm8t/Jg7rSacULA32C9dGGbzOm4eiSGx65TATubgtsO4tFGtHg9O4psE8qQ8EJnCpf
J2N/Yi4aEaag5i1JpphVIxzVwnFA1Q94iPD9M/75MmwVf7Q8HFgha/58rJxT/5hZ7LJG7csV31TZ
D2aW3RN48gYKY9HbTJoXDx9UJOeZhe/Ls4ykH/VL4JPuTHGGKkTwybjbiC6PXL2unZzctPdmBoaQ
b68OIs9CVeb4/TzWSUT4YlePv7k8kuLKJALWKCZVADfttDLNI0hXZordejPk5+SAVCxvCdBj2lUN
TtK+HKQ3UKrmAJ0mX8mN6upBhNlgv7QBx4qqUVx4+2hWIqn7ZxHFvV5/zSXFUleYlNquGdk7M6Yi
IKyqPhZOaP2Jn9wqJsiS6dLps6NQKz5Bm7OFHPffEb259Jb/dZDuJj/eg8CjMwANBewxAs1RIBOw
VVhhSpQsNrZp72+J9X3pcqFkO1AKEgh1RUku3p8Rc+qANQRCnTWd49yOuoQb+EotlSRy0SBLHVmU
b20zAdK/f/8vr/iY9jTpKWMAPIJp1j6OI/XS5pqgeM7iDiioc46DqetnBjfaLW+mxHQRd/llCLKK
pUUHrE45VS2pdGo4pKo4kkpcNGKeTXinm3v/2ANpMEA3uyiQZig6Ib1+Z55jgUrnk/1EqcBOetg5
BRy9H/IlKKO+5WVNd4RXS1dNyvRMG56UhF1EujKlZyYJndk0le1dWPjRukRnrxTMpShC5Zj+PKJF
9JcRAesW2Ky3/DS6gGheHjrUE5342wLkE+C8mT+gNTH1F3y86a0NwoY9gTsDY1Uikvg3BOm/oax9
UCyTGOCu9EuksJBrNlJGBnjKqlcjWNSYJWUIbfpRxKp+v1CasI0uAkpwmYQ/H5WPVGzQ04Q3K4AX
nkS4yIYFnHZ7hkRwcRAn8VPjlDaOlUzQ2AxcvwXfEFZOqwadUx3RAfse0QrjeMfvlql94qWIkgAl
XWS4rCtZLnDQTNdcCAwWxl/QIbPBFoi/E7ukBdP2OJNqtZltF5iwmxxojlDnIzkGzqg8RqF06yrS
UcfWsyPOeZE81nC20tMy4skEuzKjDatq0yQWI34EWrjWBXlRlHeqg1BGp4Jc/zZF7NbPota0sv5D
LYXKV9P3Z1dNLrHYMR53OA40a7MDMvBBhPkepWSxv8tXDwwXJaerGeUigwJjR0DDbD9hU9xYHW9A
kXfBtOBvZGibhaz8K+UmacxNhMhDdEnztTs+P1YScqYFr/sYDpE1A4T5gWqYQtF2oard+K4RoSl6
thGe0pzpIDVYF9knKlCVTKGDzXm8o5yhzWCKsyTV43KZqSJMkVDD196humzZzTWuTDS+HpJ8Uvaq
zERUN3ChDZNUrVUDutTyQGrxkBlHQvsfBBPlvJl7HXuwhC4/W5XamfgUxF+EHz3Hs7FwBf8O1J2I
dMy0Z6bunscm3NYg26MzSZcQ0LDJPJy0z3/wApzY3eRTSrV+3RP9vVJA4C23/MyO9Hi3goOJ/7Gq
huq+blvLGdJsljiPoEuRykQ5LKkFJ1V+oevb57rXXrn9h6apLBND5rk0VsCA2Z3vMkTBmyUDXuDZ
0UA8es0ck0RmzpKNg4Q+dPXL/4PzCXRNb7OjIhyhgwh0isHJ5NgBBsgBhpBi2ZqihkMMbqfEQWTg
rJtMeLdS38rm6ao0POqdz1n9yooCoNGd3rn0CgNvwRyO1A4gPziYHsWOZjWaQrhJRrdshqzx4Kq1
80Ex3dTFkR7vwvrkU6DGWSfl8Z4efIYlD5SkST55B6ZvPDDTHNRgd6wJAsCbs5zXd0nwLcl3HB0D
yURstwr09Ubw3fVNHWC0vGkQ07zWjb46B9n4GiFBEy3pAQ+8p396xNx2HuBy0ZU1LW5ow5KcBWHM
E9P8Rf6rgzo9Ow1v+70SUMjTsGQIvgajtnRTRku8kVxg+6U6mGCbrc2jAOgIcWsirB1KcxrBGLQI
rgEdd1dhVpOB4nPK2520/98iRuFud30UpOiiC2IdBBbQTz9wfJavir478eWG4t6DZoBr3thFsOGM
P+F9EEC7rNJC4lAkMjK/fcxnDlO0HvXRyY9rxAd1KKtlSHt/qqQw8dHV2DLmOYFZOby1uN7JAczJ
wHuAD8ud63Ricbjz2VNqY4FNN2A142NUFvL4cMexogiLY58yw0kqR1401YjMRjdAVQ5ey4Efv2Za
0YlX+8u3p+swwFsMnwwPr0anW9KURiJdU4RxYFyPKqq599xQ+HrSLsPpT7tg5xZ0ZFNw+eOAkS2X
D1uo+ByKA4bSqV0fB3hj5bEjvjm3yjEEfAn+YZunraaB3NsZCvVSGCMWejxr8xJMoM65DS2UMTqc
Ipg3eWgBZVsHkrboZnJbZgvsBlAERYoTGQI6XSbFr5pmvPpPBemrluNYpoKNJVtkwCywTI4kybYx
OwEgbJA8g/Nkh6yzqoPZ0t2WnK7TGEp2JkYtpjbBk1NdX5Uclpnd13xn0KjD+XvM99c9opYwNkIh
0XQbgs0270u+1ABUGKZFeZevYbFLM455DQtpwVriodjh92lXqixDp5TwR8FtGBRlZ6/BhRI06Eic
hMFRcAkhaacf+DsNmGPxRie37Q6D+JhdCrnzu0k2F26NNlwuZVUa7Bgaiw0dzTjMc9tw/5t3vJbi
JZjj9hsm+mLdpnbkgxH6bG+ftsoWetsIHefxvPfYOEqkynDDadr39u+18YIflinezdf3qf3+49yX
1QoupsVsfPGiJhOPUxrezzG16aqO7i3+ZHzOD5yIlFVgjF2J0S4WXPuOGwNlhf7iqMKiZl/2lBQp
S+FX3dc21ZWjWRm+eA8A5BpXwtDAUWfmUJRfg8v05K+wH8+qNTdkkSl2mdXuWWodwg1BpqIpWr5u
Xs88+mQua5yNCNv3ttMCzwXN9Yc4+l4jvSYqtYn3RZr5AAYTKvqBlHLJlFXjBFW6s8qiFfoL0DNf
ai/TZR+kInN/wRCayxBpfPeKCi9/6ysVrn3VHfldoD6hzUjnHg8PqpTEfb0PBeN5sCU9L40nCipY
2PAWugltljcfc3Q/ZGqM8m8PGOL0/kWibshs9o4WY6E7ZDUUXk0nqB5D/r9XyAcuoso8W1j7pfMW
9MwzNSgENm6QFaoKkTHy+rKkfLzFTcD0xpvqQ83PhNir0vl0fWbrl6x2VEcMf8dCrmYDB/MtGfC+
82oxgQkGcxi7EH4PzuwsglJVdkGIfnrJYJ09f0EkcTtol/FiNyE0pVDA2niVoST1jOdzF2LRm7fq
FngMBrZKSc//DbBTvpzsSJIRVcVid9d4PEJ6yGStSVbJIX4g5WcAqakDYLGAlBR9EM+WI8Hkhv/o
U2/JeIfndtSKnSOaUB5H8+rxq5KRMdBjsafLS86ajdpL27LdTU6L2yiOGWwmEdy6CxX69UAkQS1I
iUIBodk0VT+l9m/o3mmT6xjUKVSLAYcY2HTpJrzG/0LP4hG/3Ettqiw+3aVUs4+SX71nq5PuS++t
vM3Oj2ps8O1twRfylvnArt+t/C62Kl86mi1NJDjuNOwATDGAtAtKBh7oS+qn/ZmIWNzZzVmKgtIX
Ss/C6jmuxstbYtj11ipx6Xc4X4KQZkhOZBGPtnA1dN/Bw8u8TCcr893yshxo++py/i8vG5berMOM
R2fKoWxDFkd4s2f60elIaol34ZV4eojNrLf4nCi86L6hOcuYDM5JJ/xuo7rZ5G9SO8jpVOIQkFSG
3+xR0Gsot9k/FLsweybRZ42QWog19KdGe7fGFQo89p3ZRrMjTr2yrdUd9fcE3+Uf7tOSkX1du75z
sTxozvb0P1/9solUdVsoSGrLO6HFQiUOgZLXusdvfpHewqXHJS9XskWo+Twvve2UnBl8+o8KhtHL
/F1Te/4XxvWU3RHMvwNhGgM4dCMTMQzyZCV+lPvmQBJn4fhDAyS3WQ/8gLyCxMiLl4n1K+fVGz8r
KYtLT1fI/c6SiZbC3cmDrpFrZeJ9Cmz8noZZxndGkcZXdC1dVjKvTVomcepQ9IYEN5+5CwgswS16
5GwYIa3Sfn74Mig8P4G/bUfDzn8wb2iOHKDDOb+2rskP9G54H03lSyEJMUTgE4xrzRx3yJ15tmdO
q967jyaxYwwRyEkT8lUuIXz1vMYKazQ2gEj2GdwiFzyz6zvydyfEaKDdcOFL7xQo0VS4cI32Lxi4
ntXNn9oNqT32aotrdCqeqCWSoZdxx906VJOTqrsh3+nwf8QslCkGFd80/SFW7SRc3rU7cbphxlEU
MprVcCE/8dVMg7xw3Wr01QXk/Ui9JNyD6Jn/Ve+ORQRbRxrJOxe9fh6/sGdjLnu6rVWZOlW8NP2E
mrIkntgegC1WR9zNp4Fjln1i3gvo2ppPKQT2x7wDbz0w8RnLDz1DApPTzPJ+wZvpbXu8TOoo4AQ9
B2GI/kEsmY2bn94YXNnAtGnb1uYMB1SBdZFObHHzo5A7NF4v1r1I6tsFOYs+h+3B22V1UKBzgVvD
UVRRdVhwyVCXM1P40KNGZtYqX129hLCIcEb/U5GGges1ibakHk9j1ije2o3s6IfvsZuXME44szcH
iL/HXUyIQGN9O1CxuoY6nolZ3Dvik9QHUGcbgzbTbfhbbcj9YQWWiOIIjZhKW1q7zTQ7CsI+hwA1
RjfG2tW6/YYVS/VpjhP3tVhcUaGb8v+km1PslVrSEWKW3eV1giLxhVsEy6uZrAp5X5c3qvPY8DjS
UC4ccF7DI2kQUIvdaXT/65GaiW8qFvTBO8EmTruAHHxLydEfyAMPX1jrTQJcsV3Iu96rjoGox3Zh
7N7wvJSLFoUuaQz42svGd9VJJXfYAH54DToAuSLflSKKjFOGXPejK9+tpA5Fyeiuu4IMTEK6aJpt
iyboBg3t6mFXYg0rU4oPcpxt5l5YVvTsHhVxL4h2s15IdVD/3ptD7FcDeCCBq0+w+rxvAIvcYwU7
Ygm97fvoO3pvrYI7Cc6weZ/I+QuAwoObIJuhOAz2fze0yVZxjS+CW0jl270ROeOc0CyDP+gbRLdw
3GhspvVw4cg4/+hNtQmf1Tw+7clOseb9RWl+WxMiTYtKY3uQDvwSw6vQbb0OK2e+xElUVL57isXL
mawr/NPWiVPXV2lXNgBXHp7qMBIhxBJFp/KDp3pfDYvQl15JtuMNlQbWm4Jn8o2XijqT81H+MgC5
c6WPO84hbhztdwZDUrBHh9d8Yr7CvoVkHXIwyTeMiyWFHpaFC91FvlaCyap0Oa2ZEjT0rSHkk1Ie
kAjuqiEcOZnUAtNmxY3S5NKk96ykAA5gyrGfvLeW0KjJo9pAsTXXronyKj04aNLFUfLz+o8Fx/js
IiTrgZyAlzEkw5AGaYZWPETmdEBCpEwAWO09rV3LJZN7zzCtQpHbPRdQE7pBRVKXVyVD5E2oVDi/
LraD6YxPjzNBkiyox+xlDzKo1ez14YWAqQ4R+/vdx0E1N+0oODu+aSr3AXWX6lB8PJDGcSxCONhq
6cfYoxhwkJEDFqURrR+hgITpSoBIuB0GPZ0JTE/MpYFJgy3y4YlCCPxgbTTFvI3dynuSyoMWaJ8u
ubgJlCYej4pKPFTrrnawKOVo22S1p4pxkzTR8nFY+30bPTQc3CO9cqUMAzWDl/GqaA9cUqgPklKT
X0LDhmQkgQHz6WM+Bt2BorYYPWGhR2xEnwMHpTdUmaz9ORTEgQManQYBVnJ2Xw4zYygh5+0puBZV
qvQQvwftiQyF/iDHvRwQ1u0cICsrH6gPgLzR+iyQOo1454OHcUVRe5JufZI4z0LJIFX4NtlGlQKa
FchfJnFMHsMHYAIxu0QsZJnKL3OjO5a2Rx7cjXhor9Zd5RNITZCpE/687FhsaWihloBaEED1CLVu
I1ec5shagK753OyuOfPFHSuSIm68f8colJq3QSgQkqGgnEt+dAtOKgQVtYSIgOqRf7VbKheHVEbY
19qheRl1R/a/36ufuwA30RNMO0dWuWdzbgMN4N7xbBG3s9ONAuybFchB0K2w3ECmitH3Neo32cdI
i9Y2BHQW1NIw92c4JDNwEBBqXiLrcRFi5yVdvtMORDRc8lCn5ArwUdsA0MOXHx12wXat3k9Nmqip
75nYCCEQTca6f4rXFzzUEJZdvhCeVkWhAK/G1wzyUxvB8NcpzzenYUoHacn9+tcHIYlrVXqb1CCu
a5v71DmlHKhD57105APG15Ik3dsxhA0VERH+S0eyGDRKML3qUb6el6e14CZzPCqZw8G6nNw01wpO
UFmjS2QEkzE9B+0kzN7Ch25KzhX4o3Voof7vsNUO0D7DSa54nl8xstO3XRAETm/2cCyDm8UBf8yf
C6P9bJ41ga6Yoiq5VR2L/lPJey/b+DgK2jPUH0iTt4tNqooh5PaVNFxfEpNwA/4k4Gl+Q+Dvem5r
8xXKM+O/kJBSwoFmCvdo8IEKmK1bB3BrfzrjWX85iIWvwuzrVrLNhPb50bdnF2BUcWyboKXalYu6
5J/ATKctNe4hY5aqDIJNF3YNZ3RKjk6BQAnJH+tqGZpxutRB0A93qWmIFMDwful5hZznKYNOBWwg
Lw7NLOEA9WNlZoz2RGhzf8CwQR4OfVp9AfCh0ECZv5PP5zv1D1C5E4c=
`protect end_protected

