

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
CZom0vHERP+sM9B2H0IfoDUsJRy9riNTVWFr3BZpkrcd8N+2GrPBLGYjWv5bwWNFs2qiaRKQWIBH
5SL3Ros2Jw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
RCliXKg9Iz0QVLqI8b9GfxxBU1GhNUODWipyNqGvNd7T9Syer0VoYCIXvffp6DiDgM+PWpXEJgNC
ZPrITDndrkqwjZ0UurJqd8Mlj+O4jokuol/hbGtnMKDg7LMTP/mcm9YRpJxuqv5WE2ZWUtD1WAlU
7OzpzsPnbliZhM0CcXY=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Kq4rQuO4iRu44woH6WSrRyNcsAgSUJbnevjDngvc9cypuoYRq4je1NTd7KtIptAfdlUTFMhOQTcF
fyvMO0ctzr5YXTPO+6ZCPBMymjnbHRykXwGANIGORUKHiAy8zVrLHGA2Tn1n2komEaNoM+u8Q25L
d17PGNi2LYc1A9ZX79yuNo063Qy3QX5dSU2poXOWXHho+u/vL1PlOKA9tvs+dS7HzKYxYNEywyjD
k9FyesJcGgO1rBPy+iEmTMF3cKMWOg5VxnjbUI6qOTjL5ZYgIsb5KR7Wy+RP+kUhXE6TZP6qsxFC
3QU0aGkYLyynNyIHyyLl9cVQHtYz+x8w0KmAqA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
3w3EGD6E+efCt4Fs6HRylWTDMnbDGksrBmK2LrIuuDQNpphsT/R3PC062rFGmzFuJg/bLf5Iafea
N+aHJBb97H7ueY9YF/kPUqJvkNizbPUPQpBP/2fJ5zOg61lddHncYUooATB8NAF2hcSBgU35x68X
0+ZIEJC/w3FOSQwJ1Hc=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
sL/FJO3bDIPRCCsg2DyY6eC+YEqAvN4pdWi2+bTJiJBIOsoCbIwvgrvycADXfLHet65F7sNM/rTn
YIBRQ62HHXK4AhEPCYJ16a+GWujel0mLrgVipEjZe/PIBzOTjqR8RXDwI8IW2xOJhTKtdJhHoHnZ
fRLpK84QgF3/ft41vG+L+M5INzunmmeduLlvL3yJO7PaDzNzZxm4Yb6qxrxT22OrC7GODv7eJYeF
/B+o0KrZLuu0VxgdWTSijA2jO6/yo3BIW6TSbvbn1C7fQYmUfGWF6ssH9kJPORZ7fLwb67UH+6Wy
MDlUpxP5xevODOWeiaWV5Hs+S3v9MGrU5a5myA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 18352)
`protect data_block
vDNEbR29/4FTNp0NVWC0LOhkUhHosP6TZQdSSFTNqA1O4OINOC7kK7OVUhh1iQiqty+rC8cJk9zO
EzgeTN09hBy2cLlwhvdeQbgk2fI/jml+1Yxkw9+3O0HHKkwkyBGz/j0hp+w4aE1ratqaX3jbMD2J
JXy/xanB6wHU1GwPZDqf5llE8RBKSZexyqf2uz435NjqFZrLijULD6s6OnrjsI8cOjAFQTu1bBFf
8xMjwiOcT6AZAuGAG+CuHssasf7kRbSWMp7WQDJf3ygWdIrJoQQT8K97kzgKzZoq9GDn3tAh3Vj7
EoqZ5xufMvTeVOjDwA4Aw2DdLOky5wh7eXx/gi3NygNAABS7WEmo//pRlLKv93mW0H3CcBVe1cZV
UegoMoG2O2eL9veVCUhsDePDH+6QltDkDNrAWvd2o4Ybb+rheKjnVlEjusuv+1quzV8KpA8yhs1O
qympmPU5y83qcPLVJ4S9OwyeoVjp7s5X5IUTPE7aGbhQdcywAjv3qr/UdN/LJ25NuTQ2IZDYE8OC
z5diWpGiy4TaSASR6bJIfGHOMvPJWDdyJ8Jf4R0puCQKQ/6FMfrPWMt0gFWOtD3U1XEppG+Y8yc4
xdKFXyWXsaW95+ZosvOH8CpOe5ed9PgNe7w/U/DrC48SJqI+OIfzPmx9Uzawn8/JJvoFGbmtZdnn
vDcoiHFvZd1VBAHqvkgbktibUuZ95jdFTPRd79vL2MvAHE1lH0dycWbl7WFASznCMisr16ZPAJaZ
aSnOLrdXrYO7fXY3vfmgV3Fv6V+ZanoPczKnLZV4HkWiocFMYW0V3Q6CqMQzTgyfRDKxc3wiqJqv
KijKfB8IJ8CElgJNg6ZLNB3Z4xpAUC4z3Ixr+UR/W52nCObIeYO+ok/ZA99mNi+HDT0GPA9pU3D3
imlmaIr2wriF3TX9G/FLfHAESiNWl0cKmxl0/3wVTUGdNWL/ywmVF8DqWYQ+380JBKQjUX9pjYAU
XlLlxy7MHmBIjKhba1LZdv9Jik2LTcmXNNEaJju+vTCpNe38XsjRZ9i+znnP1Ch2s6XKQd5IsJkH
0OULvuW1nHC7DTy0kwlDiRJ0bh781++VieK3ELNpx5nxGi388SDbZ7GudRFCnKiatxqXXb2Np+jk
x94gnN2DicLkJd5D7wge6pqr44rkCUWej5WxMOf5fhGpjy1KygqgL6Sba4L/90ShWXCZEJMxVUB6
zifFQHRhqByrmV65F2XvLpEw1DjJh5FEc3NBsMZm70cTSyFlgGU9unsFG0TqOIviA7W2IGoIujLg
UXb1XUhoIZ5j7XBMtyVgTs33CQdLMhRrGCE/excfJuyizp5oVrTFSJBmqiEISqqz2kop8PDiZjai
vs9QaSv3TB7IKcSG2x6ARgGNXJZXthdGv620T+CgN+MLxd++iK+px2ImWb8SEsTXRA6/5bvUfpv5
97N+aeV3Ax/whe4q2tbiBl+WeG/5tsWhGbDpu4o1PkgKLKqVoNyALZvGDH/Cj6C0ekoc/nbJkXrV
uuB66FliGYx0nCbhYXq1MRE4YfbCgJJLuc/MPe0yW/Twxjvm3nhF/4b5PjBXjRZHtQFf/tUT5G6N
Rj71LiZnVfpAg3giy4KSRYo5KE5tXghRQBy8X7l/Qi4N92LmayIdMguxayal3P81XY5RFC8xOjbR
HiULxCJ8J2dJK+erVFRIsRZA9DNEOe8yy2DrTg9fjKKOHFZBhp+96zofTiOSwDpqX9rapzzdEUeN
PtBJPR1SEqTqZfjM4WcjXmlj09LLsmXN6XvUUEeEFEZ2MKm3MUFkzE8iVYDd8SvvfqfaxUaop//m
7JSb6fRw+uNDKkIyNjiOG2XSwMLYw7V9KwEaGgglck2jI223NdhllO82GGmhv1oHA6Drm2JTPoG8
FPMdS2OMAo3y8QTnRCSe9XLdDyhFWzIUuqQ4b1T+kSsFfrt40D5ExbUuF6w6SyZIWSxDtVUOXI9o
Pim3bggc1GigaoEH3IZkoSnP/hmzxF3ZQ0vM7L3gLGnMhIMsYAQO7EmUt95MQszWUc3U20auiA9a
GOj0srRKp0n5UKwlWSEibxJmt9oydYkEk03W4sgVCVeDKCHPDB2XXeWIEeiuJyW8WrEuJ3Kd3m1l
vPH+Ezs7RlgLnsx86/uZOl1Gsr3mSVqlgU5nydQsdH4TvgIshVb3fvaFeT15qK59Liq0XULfjpPI
v4vT9Z8FMH4SkLOC4BmV0pCm58fM/GcRJIrbYVuIrw59plwmoIIRdO820VvuBL1ZoKPUmTOJRP4i
9F3uqwJPQM8iEIAgFupCHWUuJkLm5Ixc7Wba0f0X0J1Vu7EjM5EnjWY2O/7AXenf7QuHfx47RehC
eVIkwr87/rmCE3Su36yPLDmqtZqZXzxAX+5EjXcLEu8N3ttfJ3YLApg7IvNizFLF3fT5RAZFyINw
j++ng3vqj9kGXEEN1X/zYSWgvRTiEEFx10T7pRrMjazQD49JoxPTCJ6lR21ix84KHiM0ExvWvWJU
1bxDGndlDQpJy0JVt/4i69rU4yj+XUhEf90rzLc2dafDwKbBgNy/FAW30aPfXaiP8AfPo+OoZ6Tx
CqRuvth4kUsRQDs/9jw7r7d2ZECCM7nCl2ZSkNyrfkXo3izstgdW5NO2Z6gfbworUgcfFFr4tMtP
zREVkApOKhL2aGg/3WHiwkhyjq2bog/taqhX7WcUnKYkI5Xl95YMa1GWj6ILFTycoDl355s+oUhg
SJN4AWVhSEEU7+lVoho9Ql9Mjzh1HEq7ThGUoRWaUaw/OBY0/qKMzBU0m/2brURv1+G0fIXzU38p
AL+qA089ZmtFoPySGm3gELyPdKesUjM/1fkoa1Px5MjKDY59K2fcsSPpRxKhsl59M/vjYBh8m5Yo
mXs6qXhn+gHanPbv+KigcKGMDz812Ln9NYbNyVFZxvMQtUHFTGwkz64qOouVw0URBrseBhIN34hQ
EYOVPopv5+Y5MZs+/Tl2h0NsdIHq3Kh2CRUT0wCk11YaIqe9/OTmatNOWNBEP5ty2b88xRO+W8Fu
3iMFIGsWdN+y/Zvlg5DvPKqER24muvZGw3P/oKElgQz88MskCAQmds+F4czpWIx5EG9qaFNN38iT
feq7+vtfgn7NIqupT+Yia1a29jquUpcZ4fBdRmVR9UUzYUgWGqQTFFB66f1/u3aNOFcj4xadB5V+
QZzXq8SY4m4LEWDX3QJI3TcQV/+PPsmi1oPKa2AkuELCJQ77ut7t/t5hLCYv/KzYxO4MfL1G9Gmd
oHT+V9eAIoQ42DPNCL3ipGmuROl4DAnTcq1qqEOakMhS6KD0KKzMfRJ4PxYkLjpFT2zkn7PQSjvr
jvG+gyA84Q+it5h/91RNulspqRC20cGcV1jyRKLgnXxNeOwsZV9GcWpNAIE3DLB4Csr9oR9jQkew
Um2Iqtb3+kfQRG7YGEbMoYGr1HXbdDbNFz/Iej0ULipwtMYAAp+GJG+FGqVyGZYF6IqeVen4BXWg
0WrXdjN0nRRAeo1BhgUFLTba+OESxcDtOm+jePe5lsFcsdJopfjWqLWVBi1Nbn/KJF/dH/NmseLq
g6m9ycdqc5yLjjrDWE1UMYeqKOLLMp9z7EpbOo5jnH0f/Ls2srFlFao0sojXhH4BMYVS48F6OFBY
7gVTZbzMJkf0drZdnm+vDQhJ07BMkiIRzqTdlA6CfDxzdXzG+vQ2gA22et1KSqtHawhJ68U0lj8y
FvRMrm6NTrFDzNM206I0nefik/Y3l5GfE3ov41++4BtLNjgz4hVLF2bQ4B2NSnHtKd67Lx7RZ9Ul
erxZfqHu3wSHuZ9pzMO9FHeKHsprOmeAygG3Cpd6Bkgs9EKslXKeZ4hEXthuuD0bM6B4z9Br4lXy
mDqM8ZoS4C5DbTtaOD9zAte9bZSYB91oKSxH+U0IGdRiaHWCVlppnFo+mtz8r6mf5wwhZdEo7TD0
+eRhy+/eluo1plu+eSuR+zOAvwK8+Ak88Fsz5IvkEpUai8xzceA2y//9apTEmimylvpOjm21XIQz
C0lzRUJuR2bb8JD6IwK/tgOS8zMsYzkKAL6eKN10je8Q9/5vKrEJziRFXQMXtugGfgGawYeA5p8q
cOkMtjVOIkgC754hLOnJmGIMsH7Nu5cebKZAl9+KYhALQV2K3RvyFNgmA9z5wluYrueQxrUvnm1J
BhfC/OL7UFgFfMN1/O/UblcHMmfrbG0lIOzSlUMFjlhiNUrFsGWaq2dAI35loTIrpgWgLFGIKgiK
wUbRs2wNtYRL8+KDW4mOZARyIwtGO/Z9q8JHvKegLgt0KJaRvBm8oPYyCRxVNLE41KUR3lnMEVYX
ielwtAYanXfIesKLgR84/1lKf4ZcuMGLcEKPryci9ZMrojjArD0E81jnULq2c2XrqchQZkZhWhB3
C2jEkoQmQu/YHHVSrK1irS34Z3x3xMJpuLc4bzGZEczv97MF9krtJlTpYGdtJIST7wi6I68Hahyj
uMsODIMRGvydkb2KTbjHccw1JwF9ub2t6IrTTd3dGo2DCOEq7Crg8ClVA74z/14GbMMqA1PNLPZy
JZiy3j/UY5gKXJRdKyihZuxyHXXPYa0jBDd7I7mmRQPb5FxnHARjrc4X6Sz83zC9TRPuBRuf2jLh
R0NDG2xfvHhiFesd/iSyOCJ2Are+/XLjbKs2M28Qp0uJTfaj4YUP+76t245EeP8+DI0+2gN/487G
nElOsBLeZx3h/nP+EkA+qqDLFSB4AarrRFyZeTrHfPE3j6bzag6ydaElCvz0Md31My4ITZCBE5um
471dLbpdc8FK072sm8nylT5btwnYZQemqXGca0aUpkn9Uuec2+L00MnTNC22+zF/KxrhMJWqbt2D
uyzgXl1wh2f+ndHRkEv97DIGuGqKgoCEh0Y5gfHJ1TWUkZ67UGf4TtEfyjFguDrX61HiHLnrClck
lyGEYGFKEuAtEPLDmN0RoIMRpLKG54ytQiiVaH83UIyCX7U9gWS6fzIKO1CeG6OakWQouyZV7R8M
WwJnduwv2TkVk5yNr8XOQXbt7pY9rUX+zO8tQB8O6JX2eZd5qWWIG7hecA40/RxPWUQLLJxHv0aq
BcbHLrESlH20zJOFsO8szbkUs+4H1IuXDeb+sZgEM3NY5nzTqdAgXnAF2mzQL8cJf1uPzPi9zfOK
c02ROzEz+GNJU4QqzEgq2hUZRcgAcpKX5vByS7iU0URZhRYXt5/GhqiAzM9hiIVBwWUKkBYbKM8s
DTXvsseLo7uUZaX4VnKrSwpRRrBQqI9xFGf5Qp3XfZZVFtN4DEjrVhnyC3TbHQCHMiTVoT/93bhZ
4mRekxducS4z74qNhi9UB28NgJf2T7uQMk11+NMf8jX9Sw2tzb/7EqFzq+SEmB9UfW2MvgCwgvyD
3wDQWqJZcm5Ld41P0X3x74Vk4SFH0HdK+3HrckaHuN3hSRg/MCFC/uM23Tk9muR124vjOBqMmS2E
PmksPELC/zVWFLAQCSSaC22dVxroJLMsaFimPbnLel0AxiGpRiGz9GrU1lXjWP9mi37EZFJjSA73
Jh22sah1rPVo04aJFKqDyM1kuFsCH48fhbJZ3xA1py5G0nCgqovuWP9JnYbwRugH418TBP7rNAr9
+Qaal3XcDOrbGai+VP3Zw/FDJA/6BX1NdF8ynJLnHS3PG60aaepYKJsj+cMaA6pfL0QXs96d9LiN
nK7bK+PiOy3PEPeWeuCbm5zUIp3JSMHw+2NEfp4Qm2YDmtmxQ4AJCJKqDktwuY7/xKTLvMd4bmhu
hY9wumhowCbyqyezZJ1fZuarjM7PN0fGcMoxa7Zv/Nnsy/424fejkPhLCyLkVo58xhLb5rGMcxMu
i3vyar22sWSjtaY8wrCC3jlYWtSdeF368d7EHxxidJIbC/5M6N29inDxmT/WwqRq4YCaxeNHLztX
RR4Zm0F5WF+kW2XHFZg4y86y9mW1O8dDo1AGesL2VlkKn5b6EGcKo/s7e9k7NPU8CatCuWXs+kUl
O30Yqy2b/njRwwZo/tME4mhBgZUQFEpyQGM+H2S8SXe+MtPmWLNW95dPVrI+HKlX/KdcyrUMPi7p
JghWZS0mIAuUnqENjEXHg+uTP/wIjJ5/+g371AgZxxLJ5TClUDBRDznw8sfSsQXNNxrFvpXPa9j5
33R5DiMqcNDxFyMibmqI1Gj2/DQI0KE/mXxEq5+cB72ga4TfI2J4uXgBs5iKCBnYEhRvAo0TsMP3
aef7BNTZU1y/OGpWJfsptnABVNFESStWVG+VoGWBIEkVoRxmTdjoD4bWUNJ3psAv0o5cjkKH1ZId
Aze7q1A5MzseOWXDOkcdu0xVXwvHnZGKhloHs+dq9bGyzdeQHJ+/7192r7p+W1ytPecUvBDbGpg/
wEkTlL2Ppj6HoRrx6ruHwo/i8XurNXQ9+6Zr9kSgB4czVzl/I/7eqCVqXaLqTJ+hXy9XECTg5NKY
bXtOd+XTjMPzwOmZsAAlnTZJ0wTRkByXoJ0YNFwdc9bd6pyt/jrLTZI+lGvksA2L+obfZzYmzWyi
gMYyoPZLhQzGCseabhmPozFaV7y+or3xH9aI+WZTyRY3rf17xwviSwZr8pq5obHgN8GiZpA+B883
nGAtUPw+e2nEWOqBcOO76p3wc+o23mQiaemYNSGgyswYZDnnJaYscUc4DsNNztzbgkZST2KhObWP
31MRAQjjtIMkiqwJopDPXDmwedcjf7gO/eI3zVos8oWKj/+V/dANC6rdnHi/dFgA3dGAF/CMrUmO
9j9WHhQSXyjkKDn+iIrddQ9WSSrVfK7MKVU/N9scVTqIwMXI5HcAgEKPfNKD4paaGVsz4yEnjtXN
VOkxcIijL8u07X4lj0mIVslZiya840wr/ezz0l6hdqjxA+iINY/zho9OIxDvdO3JeupYUP/bpnOj
qhytsrDExNmwxgMPVcUgwbWkKtmvWzm5BdSEmFY9GPV+wHkZSQ22pe9W7e0GUiNYhKHPcEB2AfW4
D6WNOwV3x8/6Yhp0lrT79QdnQwco8Dzjb6gnH4KKrOwk07g/tlEupbY5lfBFlOu7bLV0GN9BJDix
rSHWAuPsoyC2nIUGtEHGuiXmzqc1O4A1cZM1H7y/x3XLMW3+ZkU7J5ZEkru6lR32PAWm0VDye3w/
Wd7gmDn/tQGPoH1AHinSgTXmYkTN3oVdYP7aCmT2VpQHWE8GjymMzxw8EmetxDoDQ9xH1GYXYkYi
nltsBt9Yt/8/uMTxuJFZwwf9aE58PPk/NyD+V5MgqdlxENebfGGaJxbV57O6pY8GMVwHhFpFgxcY
J3tkHjiYRRvnef7QxTms5gkYOeD+yxpNNaHAt2cpM5kRDUJZ3BSgdv5lWvxyO7+0+Z7NbKcQm0jg
fM9NqJoFLHgmKr8poonIxgq48NMIYbd57+QGElnA/bVru60Zew6nATG+g6ZB8Pvjx/Nfo+qVTYKK
ZLE1RkhF4ROgDzk1sLlQnBn2ps3RNcr1VXS87i2uVUNn5aL+NPyvYjwD5e2T3jQtihpnWcWVhbRM
Cs3efeYwXP+uZ4Pqq0BalxwvohDyyCpc/vpELTTtn2cpA4b7GzyI8j+ElMMuyG8WX6ZO5GWyHp+F
67AjyJqIZrCGfckYVS0/dt2weUXs/psLcDqE0q8w5xtekohj/HzcwqWeNjLLxh0b2UBR+5iKF1s0
OjSx9Xc0mkNyjpxTdA79siz3gLyqm6+kgCF4UADFopTaYZXz7rabCV5IN6ls/0gJzcMsAkKj6DkU
v8RY8HCfahbp33bUAeTJie019b9Y4EudeAUQllROrAiLlRqG4Maw7ZAQ77qEo3SBpi4d5cryLkGk
jmSVtNM2zqjtmlY0YxvtWbNExCxYOMtxP7W4WvxBECua/sH/wVgzjR1S1n0a8JGld5F9afNB4L8Q
leR8QRvRfOBg6Vy0Fafvg3kIUnVqVnDIk0eie7lf5rsYDpTBa2F1Y9Nkx7JnFbHbO0/XXiMUAHaB
nedKakZC4mWnsVFuobb3vrcVuh7okRpLKMlOO4iyFGcCFgVPP5U3ZiK5LTApPj+Om3hZYG8YGmL8
p2RePUZPEx1ayPqI1ZpqdloJY1J2J3Vhlvf492oCZBTJLJl15RmjZS/WOdW3hLqE/2SkwC35GkIJ
SPsAdazRoGswVWyHErsPGhvsJQPc4Jc1YeuhIiCMBFfmaj8M2IdSBEqE17B1Nl7RASrvvkJHlNmk
SnlntaoBrCuKLftcUjzpsWe6p2drjaVZ0idsHSp7/v5wMw/C1qt5rN6kWVGXR/CRNuNdoF3BfKaX
GBcvmwMcYpCeJV7olhtK5hMGGkxStCEyX6oocm7XvizlAC7/BXdyKZ9G4KtT9hmRl59Hf+cB/Zol
LNy+sqjQPQNvDN6qy2gHL94r3dmNRLhq/dSRvu8pmLq0JuUEU8W8JaYjp7aw7t9GkBZLBnHFtyX4
4j9fyP/p4qPA0Mq04iI6/4ZwOt3p8KahuTQa1GNX5/nfZ5I8bWK2L+vh3mPheVTox26cJE9kFwmi
f28i9QbhqK+dahXetPL7dShWN8PrpIn7Sd6nf/NxkaU7aBED1SYdeK/ZKkSqWMs/mu3yX2mvsmqP
RiZxJsWjEBULz5UdcDSO2oUga6ZfJlyNLD6H3y9HXFgSS9/CD+GtsazZTsPyK67LwBdIHWiPmCU6
hpVwdNQ3qKtHMPwUniM8JrBm+uG4hvqbN+tI0J3kGGOFrgHSukICiph+YkLDVAvEGYDUmkplRdvq
AEsKOH5VQo2bgrmNrIyp6xSXhh8sdps7EOVu363KgSnsOu0nb1JYYekSsZShJOwjeP97PVZCTULh
rcZPaSCLxJsdDSR4ERUK8AcxVT9rHCYDkLQuT4Eg7QqiY0f14yXST0cJfSXc1wIIRvZSNGqsDIR+
41uXCVEkLhpOW0RU9sczFyF8DJrKLQtpF1JfI1Q6vyuJw+UaSG7GrhpiUDfk8ORqJRRAjv3Hbj8S
OQqqPlg0xQgKlLeZ3XTqQOco0t0u4+iGx0eKblDNjMpaSzdUeniYE01RttmVhVIvzzqHBYsBKvWq
bd+VKKfTpj//MBjiOhc4KREUSyHL8mFycs0lTQMnOkevjmz/sSIUCRocyr/ds0qFEq8GY5LcWfTO
8endiUeZdCV134gLonForGd1gdlpFcxfvckJFxgWcFUo2mrKvxrlC/IBAslO+hfXCxs5sO+ZaaMz
Gm29N89k1O7RV5N3/1zHzh6LTzr83y2ub6CdV5xs+vKIFsPabs3M1ip9lJYlgbhf0hN7TJFDneMi
12Ajj57B55dBINpdjY7cvUApuNgiOpWYnUvt7cvwB0sYwuXQ0CVOHgfaHziZPKbKsiniZqhx1hlz
DKBlBqDo+JQmJ6dvEB73qclQYNwCgEP5jkW0FLYfhg5QI/7jFXvToZ92fMfKeABIu/Q3S1FQdycW
AS/t6Ipk/l3RKocxmIIqIzXw+A3e8Nm0ZSKIhfoPhZ2HZOzcfyWUcaZ7gieKKt+icbPdbaQgxnMI
rgTKrFi5WRIg98C94XKf0Ks7HHxt19v0FICy6qzhi16mZWnQJROUavskz6DOlneRK5P15yb6ReYi
gPLeoZDzsVesTJbNuyVe1E6tfCpHlvxvsqz6XVIU82cnhWqxixZm227ZOMqsqr7AbMW4extAoSaR
4SlN1q7JPgFmPK1aZXwqp8FZ+GKOohjKq/jPQMxErmVGkJObtnq+IcyQPCoYy04qJalK1NVJ+Oap
+VEvboWL8xc8oSm6EkODaJgWUDYIdaL5bksvMGTWUHI9D3S8H9rnvGgbXPE4PFTtwz7mWxSj2FRz
zNPM6l95Wg6lwhxvJKQhYNRWaZvuYxHfNv5IBvw5qAX1i0IWQLs/mTiFw+y7GAiWlj2jE4K5zkNj
XixM0YpMRs7MgtGoplvH3KOe+NEsoSU5h7TwUorxQO2FbU8YbJser2qou6ky1iTXHXBJvz7vbkEB
a1tQxE9ciTpqWQ5p/Yjw40nYyRFHpE0ANUef07VkQSSVq47BYE2suF2wxlIkqmHkapCvDqvg9gMd
TtHg3h+yp71hp0DHOAsCf3jDxJ6SEq/UtmyzSBQOFHzcOGPM1PINLxh/GTSF6MWEzi3Ax2cOYdqL
DUGEVeKiEhRWjBI4AhvrYH/+nKfZ/qQxOGr04yomjNdfssU/XZh61wecmcmPqwF+EJirD7yGME7r
Etgc7N16UKWINkMI8C9zYNGAAo6SX9llLjIYxvME5kwHV2DlxPeE79L4Yqn5ZG12AIywFEXqWpzy
/IgWfCZ+jbfFA2yexPmpeHUT9lmTuX8j3XllhkvqwbRVWQU50SayaVkJW9wCdtpFP94k2dLFZPeM
J9kMgSLiqjApT5/Wf9tm2y/QIGl+kXiIiyacGCANr3d9A5igE0IRr1d4T6w67nAmOjayEK1XtK+V
qrNssX/cDeYwl07iAtiVR+YyQcZWgkQSG+hxJOylPcEu1ek81F+FirEJiiii+ebtEScjn6KKtQ30
ESpCbVFBY3tqaAfXCzLQGFApU8HTWDg/t9cDQwrZw5SzgUb0Crv+jSj4ndCT6DcSu7jRLwutNYmG
ytsf++p+RcXCKXsKZqywQ5ahcpQDxLdoN/Uylys0zQ8fImPT+uf85Dcmf8nG4HUO1dwyB0WPBiOP
acrZM9bbTaQUxi0mMRMo02wuc00hwj5EGs8nINPp5KAg6WiJoPHoyupclYXjizBX0fM04ygU9nVb
K5De7pqz9z4sSu6serUQPo716Klas8N1psL9+YzgC0i3x3WCA8lSivGeuUOm4GKi9qceOJqyX0c7
LFV9Jk9OAEWa8fSKsiXI0TKGYjGiePpvrBopzMAXDdBLV1o7DcGo1ZipugTUIiSwOGz0vdSQbXZP
Ix8TEkOLHbrTFofdTd/liNM6/jfzhtxZm1a4mF9l2+bjfrBiE90qVrjYHeTzuXJ+vZeFuAFcK3vi
ZswQfzHl2dsidVZSA44yvjPoU5Rx4TXuDDbcye5m06IgQn/JRqzzi8KTBlsuqZy9hCHyT8KXUO7P
h5oxzqg3ZSOaHchqh3YFFRfYquKV6AcY1pkGNfJpLhsKR6IsMDQbEOgDsX6V1iCekMR0yh40i9Ed
OoXN8SnxseizvzT+m5SlAA91oGq+59Dw8NTPfkBgCNnATZQfQptff7f+iICBlQ6yrLzeETMtpygL
Dy4+iff2m26JL0UiiDH6+5+5PLOi9l7JY+wYPnbBvoVMCb3VVt0kig6kWcSZkArNh8i5iGkYb1GS
w/WnFA51skyKSPysuMzWpVasK3ldYBa/Nc4skcNNNmPDH7qByrgyts2C5ZxzjxiTl2KW/KA9h+7/
jfoqyFKRA7s45+Y/ZO0Eoq+hq5MyfOEADNwzveTo7G8c1GuFJOHvZvnaAQj8adUHsqFqCX1WK4yV
RIejw4r/P7zOVcQ5bt2u4Hs0x86d7tDzdTheMnjsMMBg2BknxOejuthSKn+xsaeZbksGyl8XWUba
ekdk/NE/5JCVbu9OsRWRLT7V4s2G1uof5qrWA96lkMVgbjfxDl1mjG6+fqB8Ekle5Q2882Qpt0tF
+6t5JOrgHw5DHIp9owCg979BUynixo5W+zE7ejnrVEurTx3w+8HKA86QQc2MmRfCbuVq1a8abxmj
n/h0DWozvSCDzcxp7oYXFlnB0q305zG9pwSERnMp78AF2/5Fvjy0qSPeqX2upvRYZMDdKadGomq8
KxrVFkiEHdCwGLA1tQByVIic5EN4O7hv2tU0yZ0IdSXwW8g6Z/GWsX9v7mAjkJLJ0kTF60nEeV3J
Q+jegwpn25jKmtG2PyRo/CqvIs3j7vSUvivTVXlqw45xSuhhhEG+k8xgu0wSwmoepmLSlj10FM9b
uTTiXoiRCd1VSt/Zmsae5w/iFgIQQjesCWzTgdTOrSMtlyCvIM6yCJ4yopQ1o/cs8rSam+7Dv3Zt
gLFDo2t29gf2pqWaYLC4loRZ9zMpuJAWvcwTuz8Y67SCR72CHPHmwGI0ZNG0NNf3U5+xdlrSAQJO
32VaAuog9877s1rbvPPutOnSN9ZZkXR8fIk76d6CgeFXb9+s/J/r3votpkgwagi85EO3tCWoZbAL
n3YMGhaZTS/HKBP7PGNSC6O5G9gwq9CmG9lg4b9QF+FDZ0VIlD5pmIwaeJge+PYyN4pdTZzAsrHp
ZvS6DbzY//nITCL212i4Q3j1ZQ8Wp1bTMv8BmlnJ6rD3YnvbT6DrJRGaMQzJsYR+cFITidk3wrY8
02dhrXxz6KcYHRJl4xHpJS0QUj092QS8s4pxMDY2w8+JWveFM+vrtbU+5t7gptgyJvWVXmwcfkR5
uyApAVOpKvizTWvGR9I82C96sCqjuhkmk+T9uRAD4tfaMdNz4845mUFgdeBfq+2JFlSqQGD+cjZ4
f19/XnV6roItXFq/+B+WD9LQ8+EjFND9aLgJ9WhVMJkS/UDfNDmu2l3pbbe8DIwPdg3bxOEJ7ZRT
8MP0sSM62apV3JlY42IByggmK9jwYMvVkJO0jaCH/8eNj2TtHU2N+Tfz+y7qDaLRtdAaRuaVmdVu
Z2pJ/9mRFs1+RpspedZI6SDE3+KeRaPkChyb9lM+KsrVly21HhUCFh3xvMMP4L3LwVMzps4lQBUZ
jqDGBFR2suGf4GAGUZIYRJ2r972YBNpWSJaPYwDBeuaSqWK02BnDc9JgDB/1n+lBTBBveGH+h/vo
H+Vyonn6jwzE5DW8GAGn/YGTR8DX20+lUYr5djbkaJVupODt5Df8rlPJpruv5bF2bVIe9jEKcxyy
J5n6MbGiq+eU7IlzN2yWo6m1s/WzZRXjhg+WDgpxHfJH7/peg3eFdc7ts9+jaM3LwtZcx9gJ6A1h
kuOQ1sQfIwaj1j1Br2ItT49cmQmWicVrXHOii2V29qhQAw/NJUQAnVIimqIXNyP0/W8GLBR2TMbI
srvtOdXiJEdVliZrDZzo23IPFKte9tdqYAy0u1FShuREDNWqjBAYCWtclYzbExtlCC0MuewPH5N/
/aNLkJo1nwyBDmmJBow0x1+dUf3BNChK84AAlGnD5l1CLCkG0Z0o+fKl3CJImWuccHWYoI/Aab95
7m4SlbxgQEk59+rL6JdiStgUCPaBWqiUZFIQAB1uwCkbBHnToZevBHeHSW7Dka1FepDAYMSLGRMy
87fqY+3TrpzBUNhGmnhRoYk3prRn3IwTkc04uz0nCGPWNs83XjrjuSxyJJBKMPP62tjw7t2ajpSR
/BKKXZKC9CNNVkBn8w05bNnY6S6YD6HivdYNjoOGdq/QJriupx/n5+xdcF4YmcZAvEe1XraGo2VG
9bMH6U288qdREcbWl4XddQ3YSxnEB84EIzBH68p3uUs/GXU1OY8a3XcGUTBq+ls3Uq3cU8uqCeUq
lvE9Is7wD3aRR5WSAWgSbB5qrOEcKW6gzUI+nvib/fogWFXr0V3ulR5zD/3cxGQn4GrcKn/Tn6VW
6kEJFA2EuezgoGd9e9AaUKxXVJ3f1KHDAwbqsGwdKE4ozyeotlGkc47giZ4hY19QQVc+pTfUPZYV
ufzVC4NJy5kp1XF5UQ6aNTQKD8pAX5dba2xrUb2H/QleJftmK2n3kKxkkecbSgbHcb754JUxaKK/
NLCrJhMDCusjS7+X8X4lt7X9TVIeF8rFUJTkG5KbF56Z30K4nTg8RZzfOGRdQvXPCKEULUTIQgi7
wDOmn8cCsTe7Qce4Hm5mYp6CXeK3QBj9dr6TEnjREw/dWDGkN4CMaPzGGxqLCg2LOCtRQozTtfZt
gezlh35kYKWRFb8KzXOgRbY7L8KKb+t0NepwvsYOQpVpccl7EkSSJK0+Y2ccV53fOF1Af9JnhOlq
0KylAGOEqQRk7+m55OGB23kLDQy2ZfDapWFa3aUHaU4G1QI/tnRvjL+KggNBZQEspHaotDeK1v65
G7XHce+hxuSLxbBxgCTD5aSMloXi4mlOfOV1Qon8fMsyC9xkKl0TFqJc6aLdGcr1Vx9VzoyZ/KTS
khv8KEzIQwq2xgODZWKc9EdxmZGVaWHzoJCHorMWci5S1lHxK9vTmlYwJnhe30TQV7/h1PCERTdc
cE5tp8Q4mcXCcffec1D77qxtPTC1OIrJJgJ/6n6yVoZ+bGOcore4Myk1TtsXFmnzQEVIcp9I+T67
ZxHEMBJz8t6aVCONUiSqyX8aP7kqwW0LBUOdfugqpyiRUvszH8DXBv7DQxo0Qz+774WGzoHA6Mdc
qpvWR1uPFkKmRC0mBtkZ9MEuyuC9OLtvKrrk4y5bF9kR4EdDeKt5CBNi58Mk5qKyPKNUNNgIqPP5
LB+EQOU/Xu2s6ZA5iU0+6q4uFqjPhKtPwqq7QRpNoqLk/FomtGJMABDkS6U3F57v989x3d43R+e9
Y2djgGwYDFM4gTE2cXuWNa4YliJ5wq06O7XPLGyTG/7JBaQ01Wm09eBXgktLotqSQ+nd8Jw+C7R+
/S+uL4FePepF5m2cf4cBhyK0m2xw++r3/vAzD7taN3sDYi+uS2PtDluZ6bLA0w4C+QcWjFVvkKmb
1434wS9f1/qNTh1nYe23KdRYwPHLRsE1l2ymZBHT2HRaEcbY69X348IPSBrdulJL2Aw26jKPfLPc
AWqE4bgkX/salkB6J3T3sVnhJmsQOu6+C4l8k3fgGpNhRDcz2C5Aaw/bWl6P/M2AWvKgvS4sOVQ5
Q8M67NFdyhgnVvKnGe64ocqx7HYL+Dzj+ueExNtN7xLoofv4w46/Ysie/6ynBX7xnRAcc4AuZWfS
lQsSAKsouoTSgLDP+BtHmvjwgrFNsrK4HB2qGFCxWuT1Ikt0xv3dmI1rXNJ0xMsJY/VTMyVqHFpd
quHkDeTyPu2r+tgQbE85Ln4fKa6rmMyMHHlSSnXkO1N8jx3l7VOKGx4ex7LREef06zV/dn4YvUa2
KRD9537dBEca3MdnhSaJsqIaYTqG/HjbWjRJ1DpD66HFlO23Z6EsMnYzJzeJjDq4XwIkN2UMtqkU
9WZnfLfALfRlDId0/s/DQfAnIkMT17n1ikCvSVz4IlgRKVXdp4LAiMvj3e2LgiYSq1lQCiVuT2vV
Jin8d4mh/cxnu/wLY49SevPmfTDDRLtGlWATOGaE3UeEww8Tb0fI3H6uRM2VsQ759w/9j1sC+1QG
Fe21nWw7+yNiUl+BX1XGb19P0XGtyphYLfzV5Z4A83noLlc30mtebmOdgUwT+DX8nq9qFTXMragH
mfcSwvWAzV4zejcktZvWBkaYepDJD1x2V0fKZQTg2dOI4DS4uWAoB2ctN0nIGG1eiEIRE6wWGgHy
qgnr8EhbgfqGEI6Bd0sFkEeoFMPVom3i/METB8ohTCFtOo8vTuKcyP+b6PcBk9EESTMLWS6Mc0Xv
rczx5u8TCueWxLwPd8x1EPUXDcISfIJ8LQQcEEmznrjB2eHgVguSgd7rlm0grDEYj7tHdHwjI8Bt
5Zey5t7U/oi7yTCq3XEPGQJCNE2xDrRAqpbaDeXPgbesWURT3/6U4rCiIr6BEH2YzChJkMMiqtXW
LBgQQ8HprCzDaK4Dz1Tu73xBdBSWGosjRtM8mClinY/LJF8bT/qkRKpa2NtsP/hlJDud8WgJjJfw
Nf4L/do7Jm5zRQKcuVQYzpXaikRMjUkBu8RJZL/4SUqh3SJ5dpYJrNxfvYWP5sRrSCgh8EYl7sds
aVEIwzlRlnreNXLHaNart5poUMnqhVTD2nudIgVE/Gz5NBdbpGFHiUOCsz9vTW8RUXyRbJBBvno0
uEFJnAhukMP6AfKGZwdtqd9pYAFqHMw0mAVzDSMT7ZnGG0O2bJPvreCWirRSdHSUAK6T+vBEU//0
vxoR0V/TfTIJhk2W1wX3MWJb/t8JBBTdbuZMPyfd362gGwg6mobygyVV7LeZX600AuzyZe0rjiUL
eH+OHpSAUbE0yF+yU5RlsdTeG7kGBhANMzhKQYpb5VllL3pt+qQDypYcTMl1v9qbQGK/rZmD6N6j
JKS2dUODlcVzXjbwxivnHLxQpBe6Hed+aRUdsUyIB/9TkCl0eBfpjRKSt5YbK6RmX/hCT/3DAf23
jZ8VrtdzR4BqGEBItUVpVcIe5cvvgVjVUd9UFUsEu4LvwMt/Brf6PDXpaKz13LOmxOaVOfQ6G1kY
y/8kofjFZwDLbZJJOpzEhoR1wohuXodmof2xTgBAJ0mqO1+mFFMG/3PQGnxOIbcOBF3cuzKnpPgj
uItN2LCPEnkLCv5oRx4bqOfA/sGE0II0EA62fATRKl0PZFOiYVOFw0E3R6FmdEiJJyB3jID92ffN
8NK/0GI/fbJ999oW3pDla+PMB/YESRAA88G4JEdQ+slhMp1ZWsRqofhg/xRCzYDwJp5l4CpIXwJh
sFwh7Aw/zOaEjqY+guyZZUBgrS0z5EKpnToASXYxV24OaAA/hMs516u/E4Uehap7IAvBn1P2DVV7
XoQ5FIKtNfTeewPIQywXfXhz4TElXrHfQj6SQyHQAxTVutb/d5NRi099ApbYnaU90JLpll7xSVzC
XZ+yFuk2zTe21O9Ph68mgGr8KEjAx7JAjLaYSKK15QHPKMgYeB9gEy8rnTf0ypYtuMb8PSH11VcU
8o/hxO2zjRiREJ3fJBQYMAOdcgy0QLaSvQ1BzqUHqGpeLI02YD4bxcsP3PkFQDowlwfgR3tc/Uxp
yjC7RHtfLE4onSiynglVw5MOnIH5L6zEazOcdMlXqsV9AA9glrJmUcqbxvAjycRdrDAuXjlVOH4V
qeoMijXETSyx0HlXiOw9H9c/QU80Mze7E0uA2+2isINtXvJmnS3srFvMUSRC4I2YAZeUQxWYVUgd
/QPZqjQZb7M1X9h9Q2LOMrTFmBQZFHVLWXrm2gxipcDerf5zesgPHm9fM6xkwxuxGznOpmLNgyM3
PUUYBUC0t7PBrtl5wl1LozrvTbchd5B0DZgYzXpNHTa4hdYeNXuWvNqon9HR3TQ5HB5JqjAy5/oR
fjM/m2BP9H42yE67e9RUwY3hpZfUlXqnljbTBJVyVGri9FZrb1Vvt0qCRXzpVsV+YIKZkVod1KBn
v4GizLiP9fd5eMLXZlZu4CTTycJc8ilp53k2y8CxMWT6/SH5gFNPtoaRmWz6PAwshTe+HIh9DDha
BMiNHES1ERDo5jQKlpypyBzZr0BHvQ9AV1H3Yz3GJKNMYC+7mHAV7/JgEoNjisNDpO+vcBbJs1fG
R2+2UTNtVLWaFZugjLm2IkxPtLrwiUMVSaKtWUaGoxpCnYLA+ex70vi0xQfX6yrectYvE6qSps+e
wjO1Uu4g9Vaj0lmPHOOpDQV/qoOTVdaTj77dvnM8AWmFqKEob3uTdmZv3enqboKUcrFQn4hvLMGk
IdunnjHYp7lyxfLB+3Ee4tRFdemKPpBCx6TVmh5hu8M1dm5pegjwkg+Ooq8hSM2UybX+is/UAnoS
XkgP0y3NLR3wJ3ugHSqbbpsm9SReMhJk13QBLCrBIK2pdqvYn6IdGYK/+P30MTWr221SMLisi2Uw
tiAvCoVHVK0bgekUzP+qpBRdmFU2NK73uZx8VHhGSTYLgJrjCXFzi/TnlJdSBp15MFfZoL3zspVO
cACytk7ykO977YzxKIgZZFgQGso2LxbGMz/co/zYTmp4q4aH16oPY7GNMKQvyE5aUzVZS8oKKXSN
tz230EThoZuX4AIeopEOHxLxB8KDeRGhR8GIck3Q3aK4BTwd2iZCw/V1j3f3Ugba9D4tw6OIlI+g
UQD5mAWNdJ5PLQTXw2HnNIgmpevOeADUGRh8nTJsjqhnirkRTiWZYE6G53BV5Y+F9wneg1iBtBnh
i3n38JSiUP8UhWi+9W7ISs2HewLOdfUKHWoY/d3SY82VgynxZ/ZYUKrxoVbenmyQF1zybeuMiFjL
pFM//sWqCWKce8grqa71j9ILmsGisLOAm7rwMuXsyGokSfT+QzE5GqelDes8fntOVk4KMiv6QbuR
hJKlnh+kfyXYdofoEsqpTrzA5BuN4RbBN8uIvNe/pGIarxy4MQvKeMgZk61jROf1rsxF56ipd+B7
pIWxjYLcI6C0wGv5PzFLf7ai0TNTMnkS/pBYi7lqo6axYCGTJoIyB/a5hPJzh4axo45XBUfgc3qr
haBMYrzPBmgCkEpzcE6G+zCC4QfVvGm+Zeei3Cz3wVidgV2tTAX0NW3DxV7yA7/oSnnt4d1p/V6U
mCvStOKPJyDCYuF4v71KnXvDEaDeVZ0blvVn69PvQYPAkJWS6aHg/5HgjaFnR1ax/TQWLgXut64L
jYEeQeq5t/HAIrvKjmJcjoJnm4MwtO1F245PSYcYLHbnGQ8yIjN+KdExMLftaeR2faexZuoqxfue
fRT5eI69Smkcj+p2v4QT+eA39gQfhbHXIayKCeLluQFq4k6s/hFRq6Ezgw4rlZqKUHwnFF4wNZIb
JGkfqURavvpbDbJ4r/B5+E4FBZ+AJmrU2Qy6Yu22SEuUWjyuyvneSMUsyJxFsTBsNEhaLh9OD0la
U2RaqSkopuzjUDCh5GlCOpIYk0AYlfDM3l4zuuHDEWDk1k8z7hSYfYIUomPscfa1RTMaVGr/tomQ
dprJpXeQ9E/sVBFEIlvgFbQ+wXeBIdGlerBJU1oZDcudRkRDK0hBzxWtDARoi+oQBfy2H6agksib
i3EBjh11PprPRJ6SYxes8szXcqvxb4K5vo2mDzndDCweQ4Eg0UmRZyy1JQ0Ew+Gtw3WPjmSNO9PU
UjLm8G8x0ZnIb1Q2EeFXLRZUnA0yeLNQojxaINydEgC/wZjDOWY/bwWHn+e03B6CdY769jv7hGfr
JSS8ppHzMpESJMRu3ify2MnVx7DnK5CMrfjf9+qketpw3pcBuaPfL0/H+TjGZUTRGIlb+nnx4Ci/
eoj9yeerlD5v1obxyVn7d+2JhfjZC9jetMLb0+2p4sRmz2Qq+N5TXWMLljmB0iKzePsBwYBD4d3Y
bGYFY8YVtdcyd2uylBRYYzEDPqWBs568Jc4+RgN0o5cWabxU1omL3xFj+yagX1knbB2WjWlzRvUq
kMgaMnvgWVe0UBT60Ra4pkM/OzxJAPTqPNuHFqKv5aRTcLn9IjAuLCniY2M+I/urqcrPkL/wR5g9
y54fQHQmjEOomSj5i4bmrYYprhpoGFBBu+rpZRH+f127cGLIi05LfmXZoK9P/0a7iy50u7ZRS4jm
rflFxymKoI+FB/1FT2T2Mtbj1d4nLd8qaoFTJIor4ChF0f5PqgFiemdQyUHE1DRDZ1JQQHZIJccz
xfv/FEXfQJ1pSdJwjyNmLexeYHG/QueIQct61rwWJCAdFY9YPpq//Sj64brQO8tmQsU/EqgGslKF
Qi2jXxQtKDcAY4kLJKfhf5+3YTsYfkKMJdorX2F3K2UXhWHJrkzTZ2iqBa7tZTvB9EXlMeQ5oMMj
CSASldwXBF8RPc7tLxm7tKci255HatBWmMY6SgG/dftsx64Ppg3b9UKV/yOhYTxmYHHTI+03IYac
2p0dZm5NR3I1UaSG4vhyZUflyT5po3H6EQjGLqo/F8aBKBKeHbwsWRXMsDjpYpezDnRlWzOQDhMK
FRreJDOMFZdQFiQZcGLT4fxP3G3lystrMp8djvNBaFmb/POdqGm3uEGgWpqFvbl64pxMzB5WVMJe
ciScB4n3zK25lKQiNdKh4zwvX1NO0Frx+vnAoq0QQ7Ni7WswYkLu2QjRfiNkz/lAKNSt6m5aMghs
HqHS4tQ2FPmXGk5Q+mIa13yPvawalI1iYvk+tx2gPU2hyE3nm9ULcM5ywV1gTTRMnTxhWs+ZA2d4
7zjeeVyznpI2PHs75VBIvDGiAotx96yzcBHSKTTn7TkgcxiADblo0k92T/nUbXBuOu5wAuk6kWVm
6fbFPNJE6Ij6iaDoYLdWHc2jyPSxsWJz9sDWo9ILWurY/k7i7ljDMBZUGivHUd++480ODJjke1WJ
45GmlStGMwxkGp8X/jmAHv6x881iwxpSU0UZtXcYkxUCAs2jMDQBJTjKScyG6oD6cWAiP69KcWg8
z7MQ8IcL575ZksZD2W6BXLuLHO1jyheBJHlHoBHSoPH5hRBS5fq7aH3QW+BffcpArHWMCgLXGGkp
/Q0idmhwEgz3KdTXtmJ4iIAyO4+GiGUn3f9/52HNl95++IdKEa6bgxtJoSAMBLcL7dftW3aUAzzQ
0RkmCYG15JfX2bVe4eHx0FAGwnnpkfZs4Q0PfjG1J6dSm43xqwcg9SmTIfKgPcfDyIx41JorFfh1
NLyf9+egUNg0qfunBzG7s166MwDJj8ibuWwDsCINcN+N0XBe73oFBp8NHSM9wcN5YitaRViAKbqG
J98FAkoJjBbaVi+U07w77VQU+h/4ydJO8F+PL5maHJsXI3YrOisf5PDvfdD5WwTMok5w8sZL6Y3L
azo52hautmf/0Ly4iHaiIoZ7QWNeKwkRpzkLpqvRUZEsSz+wYXVAwGCJoi1s7l5TQtXcbjnfJY69
a0hIKecHRhiF0uuMBMSbLqM3+9GzLZZY3XWlbBKB0i3fHWPv8JmmmmFusgbVSCJLh/A1wkvYQrWs
itocKVen9TZ8gAuUNQsg8oiiQujlNLnZtOgNNZXlu6KwxyjN8kXXnZZ7lJUA3yZFzltyibF4kfzo
6chhnjnFcRw0cDsf+g1RcTAakqgpHyk0YnHbmJAwXCoU8dRlPPmam1xFVnNmXaeNEZtVwWKaBxjf
Pa0FF9n+kJfG5YQq88nPk9G+eP6a18HgurpkNGmXQsW7Tg1g/u+0K7y7/9Uc7Av2TpQpBnX2RxZ8
T5rGd7V6G5PN3wF+pG29/rxBAGbUXxkGpsGUTzYFIjy53KdcTqPtKWy8jjcChYNIBt9M871uWUVp
vOcZOI0NBl9GfSWuPIfx1gFnlwDGnP0nP/NFJS61DyYJKlU+E3Rl1Kk9NrvLpc6cQfELQhdktbHp
MRfi/tzfcKf5a9lB9WyheqbCZM1XiLN9qdfPuLVrSnVcGS9bhg2jKib7N8AsORm5VoYawi/pqtt2
x6Oi/zm6aE0LgN2FcErv2QpUVnYTdGpaRzGvnPe6Lx4hj40k4FWAiLahiVuPhTSo5ShUStMa/1PT
R8InKWnbe1JJHspMDpozqVo9OfeAl8qVl48g0cjYrGI2VaAbzM/wH05/W0VkL4R5oIND9MmpSIqK
wgLnJdkg4qFc9oOpntY5cWJp1XszqGkS9g3rarcqeIobBG5fvzUoAM5K38iQMfKhz6Ya7MQNbilL
JM9BJGwXNUU0LmZrFCrZ2WrcOhA1TUhlTK08dNVEzBGgKCmUWmCbIsSbZ65Q8yw0O51YXtT9HXKD
WpbhV9pfKzJpFGFcCaFTa7IzFLFYOpKk5OepER2HT7pVmbT2WoluHVlzgcI2n3qR1sUlfS/8dpuD
inFlnBPh/wCzkXRY+wZvc3G89EZ5XuqISBbuO35VemfG17ERaPLvIwzSIcEmdcUZ77/nku8WNKuj
IT3g0N1Pge4EP5BTL2wxHVhtg0jNFh/APSdRPXHoJZ69j/F5u5Wof9NiOM5o8BfybjZ5WiLuFmEi
j9C+zDm7v6xztVIzRt6jEJnVg3RWFocHHK17v8/z2NGVhmElPQqs3yVvpJ36iL/uNIeKhGvxNVpA
97aT894k/i9tj5Sb5hmCqb82E1JSdnZjLRVfi16aNAUBm458R0za5ibp9jpoYOX+QWrHm4bN3rX/
VQWXs0DkGLyWtJGci+K0hZ4mtM1KHJH8Y7uI0HxP/J+eSgjFkkXBsj7meo4ONHesTKT/oyrlARkM
tq+lm+KuJsp4o/P91YJmE/TlqQXIINDxJfO47uq4vzfpLhjki/USMTp70JsGtsLW3Qgqkq1BU4oq
cbpzFRONbNOKk+dS31+SwodymeAl3fM2DE67YSqHTlJ/5kpsCidFhe+KcUenyi98rylCf1Wl3S8m
QUlSpN6hq3uOyBffZ0kvKJDuyiRFvaJJGmVO5WED/Z/07XdkvuKfgQpyVqXKcaGLW5IyfoaI3jsx
0M1W0VEOW6PiXltEaEt0cFiLl4pQNXuoWiduMl5KL7oVIfTDgioGa4hroDIUxFZzwDVBy2S+Ig6r
CbBcrLftwc+h8NnLwcC9tPXkbd99YjrYj5PyfSjYI0ktOA0Ubdb/CsitZn1RSpXBHGYG7qSLmxYK
nPN2Nt/ktjnqlnAphPIizR1tvj9EY4VPWtQ5DTx1ggj0PNvVFVmQj1ruvmvuQzhshx+PG8CT1ThV
WEVjcBkrqmpr3wdzRxSKUgnj7eUz/w3C9MzyMpwpP6ef7LI/glSR4tChMXrl95Xenv7moWOlMxDT
gnZVRUsbWvR/GKdX4zBmvWGu3rzrd/ThLSPil8DabZVNPvViDTSF3W1RkBNDSIZBwOH7Z6HxoUjZ
5EQuhPCOJDpn+i7Gb+f8oibSpzy0hd9OUJradQ95zMgQ0LW3bIg87xyxmYYchGkLUPRYR6xWBU80
utQfcI3ShdB+5ez0AmdoWY4RevhwmeHFAvcV519Tm7j3aMxw4lgMuqAC/alL9TDHpOxsh4c59RQ0
Sr4wdw7U9kO7GH87tN/hsSV0ARTTugAHCYSccxZDtqWS4KskEVcM7lMexsz1t7XDLywykK3WE9XA
lRCzGtT1WbaZzXADHXOgIhUxsMFT4QfhNNua7BMFHIMk911jtmTh5X1cpvx/CamPdaI8WS4A3ETl
Nx2LSZqEnWQdIxVy8vw6+QAFG/jWMsubWPsdXYbo/x16PdXXE9W3BmjG5p0OUrWPPOoznNX9SO64
6rVovwf1s5DyTbHl6vmJKdLQOJnNIpvao7rS0sfprjksDwQE0oTH5mVYiUeTZLKwNIdid3D52Bhi
pL7qQsjt0vCbA1NJLsg3EAD099tEx40dQfV3ECapQZCQ6K6TVFZz+0qr+iPiIhHatMGwbF2R9LH3
+ZuhhIerFNEZhEVJRT6PU9pkMXzq7urZcbfOVirmbFfyW9sOwntDKklkyxHmHbtUC1478YEKTu64
dosKP1pdO2uNYRJS5WqC9IDXSisgLtnkT123WLudPVaPg0GQSDNN9rjKaBlk/suMl6QGQtI+prEY
af/WaO3+qKl1LSacLDH4kRn2scR4TYvMyrZmPuorpNWFdjUr+WEK802OHixqXnqrIhn7ZwwLU/SP
Ch7Xm7GQlMr6w/5BzKadgvEURnwJzhROfgjkLC3VnpyuFDKaqHGvGUz55YRRH1r6mfv0pvBHSR+G
UY4kPn7TNY4I4N9ynQDSZ5B393KukFlBZFmIj3SXIIn1ZXIEnxU7m4NeAeIX2uoQgerRv3t7pI+b
1tb8lJL45ryYXe7pIPRTVu/wAgNgrGjY7M9Kcd8c6TTNpcnHPaiIQUmq3y79fI1pzp04bQ5ljNCe
8Ve/t9xvgZpvqMJe7HlcQVohJrNA7NXlSH9osV2H/6SEuQLEiB5x//b5SwRZGLRwwb02lxM6YXoM
VyD/2LR9seWXOspKp1CdfXlAEF/ms7WxYfTJM9aHyzv8nye64E3dUz+jmXjybksTCL1YvIt1/WfR
ivyPUTv3Qv5BylAX2J3O7Z5+mdNQB0wYBCu5iDN4gB8JNyKfzhyjVfU7lPbWgsuuxXt6K3zANHe1
9aiBeug3s+zYWFucT5kfNfTTHIp+X9a3RqTWeY1zlnXhwdVyyN/j6aE52KG57/KSQ8YtdfDZXRbR
ygepzzuj1PhwMskwXeDzyeDeCSnFDj5NV3DWGmi4oqPdEtiDlsuSwZqsuzDsG2xhUQTKScktRSVf
2u4DY8XktLx74vcsHe8qJOQhlgbC9xcZ0yBj2hfrqQVatGusAmZ8/u/SfoslHFjm506oe/keb5sa
CkiebtE5DkWaDZmMB7AhFF8/lbyNWtX/Ja133UqMtkMq7pwBUc0gDKxCpdFBiDUfGLSCxU97NXOs
aC4YHvPRMX3djpFYTGCYWo3k9W5F2/nm47zTXtae2UTiw4FG+trHhmGtGaUoufYLbqKo2/XSkrh7
M11Q+3Jtxb51Sn/1ULVRJ7nneLT3Dx/I4M1xpT8v578qgC4KXMbqyX/yVNdultp/WqfwWUfQH7qy
hs3ZNF/dq7O+Wu1y3BYbYXTXTE/PNZWL+qXWen/RlughflnCNIIQuP9QSoJScqoF0pZHsfcFT3C7
P9vhq6e3VYwjJA2abptFwno++IMac1qOsU4sBTLx+xyAWA2wAl9AIOW2n+dlHhUyRz0sbr/nvxRS
WqciYyUxR+CEWHJHsGnS+Fznd5+QJzK3olRC7tYpt7+CVICJKMYSRhMWrvTyo9oRMs3Uuq4D5NJc
O7CgXcEP/raMJwdlXy027wOLs71HYLljVQ9u1ENNZ3NbRLX919kjF175SpdtmYqmR/CVRM0enRTc
sKgYMORfpl9JahrALbZ/zhG3n+ZL64FZWDt4unMQ4RBCf/v5SiL83CAwY/lNrNtMDcMKRXVPtGhC
OuzWdl/EcU6N9zfUQRZYk07xU6weRHfdWdN5Ahc0x5N/HWbhrjNH22zXCTaYvCedFRd81D+Thg==
`protect end_protected

