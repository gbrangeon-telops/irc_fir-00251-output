

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
g2RN5TBir43ECxFrT/y2GRXX5NGDYpjq+n5gxNTYWsuzDCjF5YeYUisYseKLr1ryeyQynd8Epzt1
V06LipLPYg==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
eJKP4nowQhkS+sdlDJ3aF081jbTFWdzdlOBNNOlq8qkrol2Z2K32WIgnl06Lqx6yc1xJY0X0kmV8
eOkRE5vog2ePPioAy86OAcMONOPoHTqykW2qaaCPwvHqEP73jf7t4R18PaTf0PZeg4kzgW5BQXqF
THWJ0viu+pagUeVYQuI=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
MDIZ/fTOzwhXm05ObJ3zkVB2FpJAN9o34cB0jHfFprFQZmUeUQ3tZW60svZwBPLmTXGm6NjoSEnE
d1b16jr2OvP7e61sGc1GOIzSD5lAxq6KYGFDCFGlb2HKuXZP87xm86ePu57tT4ld2oGvDNavbknR
LLxhx9ZyBV7SuzGo3PKuxBA2tnF6vIEJkp4n2dqwXnKJw+xgySn5xCMvJuNm4ghYOfBAsNQGJ39j
9OlCVz84SN0I+ZhsnI7KhLpJBWOyFN5hfdsD0RVsTRLOBu1rLKX6200sXAdAwmaB9xg+3o0vilh4
pIPe6hkIVYlfHVKU7Znj0kURPqGkJtm2RI+CaA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
RvD4A+WtjqxHYEUrji4gUWEBsLfMuiFWzgBi0pzOF5kWQsF7tHiiAC+dbiIZv5TBKh6/SeRqqj5f
up1ybf94wq9EXJ/d1afld/HRqNac4VRPTUzPBHt4z5dEncFPVDK4ucOaLAd/3B1aieNd9xn+mBS/
wR5gmSxp/s9f+zaVsS0=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
NS2iEv8S/DLjr8oIhLcaUy30De4W+2t5q2cf287k87h3kSCMEoBnjvcyRcG6CE1IFz2i6ewnJ0mb
4oesPU8Xde+4KmwGSKnw2OpNx1aFtJHy7C5xPLKHuYCmY+9zM9y9RMguGvxUNsPvXEO9G/4BQZtJ
xHf97YW4qiiYtbOsAO8R0m9UHVOYT94pj/6x0Itkq5yeU0YXuubMwNfZ5ZRnrVKNyxQ5Ilm1kGqH
N2bcD8eyFlVJydABBBV388JKwKrfOh5ZHUd8//7U9+6XMFYO4OGZzTYmAvyyO7iRRKEjPElnyW25
UoL5ziiALbB2biJ+eBPz4dgChqDQ9nB8HsYg8A==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 16672)
`protect data_block
s5ZxkCsQaP1dt25n95Ohsag0oVSB6zp1PYYhvufm42jIi0bm7D6CjmFi0A1tx9nZxZenZahrtQ6i
rjYaTlht3ThH/9WePIsCUhD5Mu4nE5WeGFz7spDcb6epDvs/tvUzZWlOwbrmtZdv/h4+NHKFjS/i
DDINZKL5094tgPFBStWecxh3MlIqNp7r3gIHB2oSbikrvq3BCMbGjskJc7d0MGu6ZIiLRoB8a6HA
vkQAwx88/LL2wK3qLNdBLDvsztw4DXphT/oxQwBqnwdqky206Wb+lMo3Weu4kmwKAvKNeBG1wTsf
pL2wxcx0vCTZVoue9MHNrIMoHhmmKgwIgAVPslAsKeTPCtvmebRSSaD6Mh86xBkpGIzlOh+OA1lX
eHnErxcMV1vOmPl0T+7YPQ9LBFn7vcLsfcXPhVlfmPT3Ig4I8OJFDIz4tiAzsL/ChQcCeIMuRE/m
YsydAFTvAVx+nZKkx1VFT9icb7jRxREI+dJ3iMcj6kgdGnIks6f0SQmNpWV6bSr79bh4YaF3+WSg
vUv1ZbeRj2VHVqLhFY4/sXUGYO5OcGxNYKVT708+US+t4fhvFj+VgOTIkUiyqAyOZesmcoK3yBnk
2Rf/q9IcCylbyGL395HcXbP0y0o+g+vAsNSxlxmPjbhZzRi+glhTHrYofjmhiy0b1VmehHj79P9K
4dSOl5GlyB8z4POiWE5m60Pr2OBNCsM3eikG8IlULVY7uLdPstakQCLuW9caz0n9/o8jcppx+yS4
qKIHugY6gH5KfHrmYwsozuM36tv6R0vRPBBkERM2kowUXAFFTk1KXKHAoJyDNMZZFGXVTTvFbhul
KioJHiV0WtCvTjofS6bwX3sp6RNegG0iPk70b/bhGxMEjO5zY6vGd3dWopLg1/6ap7HoUm31KX6C
2zes1N9VoSZWXT4y9fPm2Nv24taXjyVXZdNIjC47CIiD2pqrBA+xE9Vq6r5fCJjfX+1/cStOZSVF
uHsZN4nAS8NjUB8rrjG+m8rPXuPdc1aZqENKzDpUikpC0JcUb0l/mgaFUe8vXv1zhxHGk4+cTHxN
k/DEn7tkyRl6WC2zg/HaD+I3WtYJWUBgywIwn8msCHSyvKeKxmhHieE/18nfXXAbCHUYamT8rt26
I/4cE3ha5Kx2WcBkIPI9sQV8vGgNesIq4Bjhs2vfSmY1lAoEW5fEm4gX6qyHvcKO0NwPO246BGfX
+ILBGMctfdx3Xw6i8ic3Ak8TQdlrPzPkry9KjuHfU6jLeX03ub09NDl83JI1eMu3mhCwGpXGplaz
i1+Zmo5VpZP1Z47y9gA0erRCqI2JtFRyJFuXYwnSY2TXPWZA2jW3h9PCWHgI7yV9sk7U+l7p7mqd
LQQNjAWrJ4bsQSLff9Avx9fM4n0BiXD1N93Tyv1sGL2HxM6k5W+hKy1n9WRFdNHkPXBK4f48cJwb
kK1fnyP+WKmO8QgibESTW4S2kO+ncGlaOstMF9BUb1BcQpICIB7m4Ri3I8mNpfZlYDiDvLmFgqs7
wUdAuHKyG+6lCaUUXUlOWW9vgACiFG0ir9BvzAaEm11kn6fHvhd95tZ8RnOk5vqRXA0XhnSY3ipg
ctZAQjdrmg64LxyZ9XvKN5V8mQhcc64mJEROTTHGYNZm5Mb6MLMvRu3+8D+Oem/i5xKw7JeA1qKY
M7UOvxmpk1VHKgCUhL/cE8AhMbRT5d1lf024OJCLUMhbvLh5UnEvgRk0+tk4cB22HekmVMLtCc50
AWbOuxyJou/nDe3u3/1jmxVZIBxf6ZdM8FNmAkAsT7cwDivLznb1QmnuJ3nw/MKPwSzohb4njP51
96tHz4KM4vXoCX/XhgXdH8h6fhYxfecLtcrpr4kiyl8Eel1qnSmTiy7PoM29bUE3rAl/CnsgeT9u
l+HveQAVr3FD7pewXgADuz/7HpRviCScNDR2G8uRLcLPh7VrjFlHAOzqBV0wmzAGobSd2y323T+q
6vVpHXP+aSZYoglCt/gUxQEaTeNQ7DO+yHFdeQeyxNUGpO8b4o7/z+jHtvq9QJt1LHT0ZbAz2Cvv
JQtOum/Ek8ztXDPYvC0OfZqPnCX/TcJxCH8mGE1LUx83uxFA0LqDYGybZoqVxdD+7pd9tvfPZtlP
9d9glkg9VIm8xktlWSIvOvQ3oLuCqjDEArt9NWiGCgo55S21/E+BAFUbrcQ7Lp06iF5JPbAmbaZy
t/VG0pWlTB4WbpKFeFUKngOwLdGILhGFPZpG2C8dUkDhZrk7oCskiqTfwFB6McEf5DxgYdcU5i0D
UzaBuBWjU2BOQpAY0CmnGk0WPom5EFQ2HvzyGp/UJEuYLBeUU7opJkWcLyTof/Vbja0Zr8Z7V2OI
qsEIhDB/0w9c9XZAkI6Um6KdMyuyvG5THh72Rj7Fyt/ILoH9nGDhdDXI33XYLAeiKzrDF5W2RkbA
7w6yhDE0DVJRjaWsBmq9S/DZppWcgAG2vEutVW+XhHCHtOLgvXtyWJ5Pb1wUH0UWidGSvFr3Zk9r
NtyW1Vsv8dcAGq1kNbIYAJEOxHlr135BFg7m1IikJTxbEzfpFUEaXF6sSeYoxpN2LhazyyWq56Sf
YYi0Xea8SnP9AgfmxPoz3kU61gKiBmQm+iah1foksZXQycCGZzjUBqrADNQe9BTSJsq0H0z3VBXx
sBURwnT6iha/Fo4BAosvaGzrcDb2vq08QYP/h7mDrF1Um0RKxMRq9/zYw+AQ9VU+yUgODZr5BKPy
O0aE4lb0NarjqnXwAvlC59GMYJcVKSNLo0jKwUyutYeeTawf7hajNBFFsoiRdsfuU+QT7pmCKa4s
mGazbvJQI24XoGAIg71c+Wpcs1VPwRAOAsqDYaGG/mqguu5WR1AfxNfwy9MptRy/mnAcCs4oCL3g
XSNI5remC1hZh75kw0D+o0BUUWK9II8vWAbrfiBwAH26XdT4+Mgp/C7FElE9TjL5GSnU27f1VRsM
6NukbvmVTf7FLksQZnGZeyAPQBO11R/GsCsMsu7TyeUACdzxhbey3IZWRMwK+mauwbYgz98SB5Ow
Spl2ZyXzgFC1a7APOZKqHVJRdROPmiL5AcOP5bZ1DQTGkwrfSmicoUnZ8Wt6cFwAm7i/DgZd+VYc
RKB5lV2h3hBpvJOeRd9QZh2v7ay+H/lQTAROkcJHwtSSs53F0U0UHJNYeL4JJx0ObdpMTMt4x/ll
da3+roK+BgP2qhV1xVd2f/DewUWggu20petXjbADMe3cpcAm8DH/Z6XdKz4kh5dcxtbg4rO8gxBx
VKz+7anVPiWxzGLMulQMwasxsb7J0M9qm/rok1uxmvFEImYqQM31F7k670UMIamcTwEVLAVOObXf
8J7WG7mxdq5V6UzBG/r1E4MILYgnQiCN93pF8bcbuAkCkcdPJbvHX8Xu1L2MqQyEcK7i6+NiaTjG
PZG0OgGXuLKAGgK+nAbhJkT2OcUJBmMX54cNNdRLczBGsT2B3p7xYA+OIQlarDBy/PDsJlloegLp
MjpzZPl4WCQJ2xwmf2g+VYkopvCaZaoFB5Zq3ZUu53Xya/UChF0emF0CsOpswmO1JvP8eS7s/dX9
QbMWaDmUuNFQkCAF2+or69bhRLH6MFBO7inv4tUprupjI38OSRCwpS/nGOJau9YLqqXsHARf10dc
k7KWtO7l2IfXfsdhL9dnMNotcCUYtmY33n0qLQnuaUTuKzRkF0N+vwfmNyGlQek+elxLww+HEhv/
1mE0O0mMQ10RQ4nQ4zUz8gsg6Q/76q0CKy83cczaYJU1YZMC2LPsU3EWcp1+kOTGeZXndMM9h92C
oHAtoGT1RG0BE0xugfoH1ECAjLX5caUx13cHFBxohG0VPzXqs/W303sNmhyv7Vlq9/eXLkL5T76Z
pMt2nQWs0wA2buGmE6XqBxU9N2rnnGgUaJraWi/nOkCMzlpqlLe2cTtfs9/KiqGao4HcyFhq5vKU
Lqk1oYJWJzgxFzis5Nw+8H7q2qeGD0EnTbPGk7ZfdK8VYTS+SliSmbTfPhh9t9z9J1uumApuDda0
5hpwK5FmQdRdVHMZD1A/jxVmv8G+GQuBgBWE303s4w/oDsmGqCZj6T4/YeM0D6JduVCQNQvJOf+w
zlejN1bQhzinI9h9f4O8U5jVdeKpZMwPL2IYGJy+K2qz20Z2EoDt14rz3HWLmsz4+HmwyXiwtyed
EzL7+OwvEtB4bBxYXPaaOdqGULsrU5ASuLBUkFY4QnmuKgCmFXvI9c5wCPkQbE8DwZAA1u4xAl36
sWqSyllLXsvkPhodzGm7ReHPjFl/7bsHMyQ/LvIUR1FGApeX0jkEOSOl/q88ADNg1mmkahSEJm7B
NMnCq5Tw6pktNjhCIDPjTLLaRp1FCwsf8qX6kfmp/T3401bC3JRwBVpz0LWY2TcYfYg47xLZJ4cq
yaEMm91A2QVA1B+zaGbwWaoBhKXOCSrT8PJ2f3hdCwBUvHyxpu1YJlhUlc9JqpYLG9EMR1EX8f6o
rNMEq6yyVpzLSCtX84t6XYOSLs1brViuFrRiTqfmaAketxIdySgfS9lD7G3xtjhWDspDJDT3oQ8Y
MRK6RfzhvSEkYPa8UpISPq0pVtsVmXy8N+IRH+yKPdrFitn71h7SsMgDiR562so92uZCVEPV+Y7i
6bcE33sqLZyVUcm5J2lbwo9F7bQlQ+D6NG9qwsjbeOj/Ej7fdtIg0hK4nzDUhMYVORI744mekb/R
9tFR2XYX8FqPLr2rttG69Aa0ViVLF/wvl00XZdqaC9dqSUtjXWa6OdUl+trnLNh9/fHMrPu8l0NW
eV0+2rOBctOHIBTvoFCjoWaCrSwFAH/UNnQkqI2F2ETx1UuWdgqwSz67f2/Yx5hVAqOt0EOyCyA/
n0xsISE8VDm+fzxevU5wr9Mu0OXn+abThKgpsVR7kcL5iGFu5UQ7sW20Qif+7HaWfN3vT7P64Bhl
HA/PPd72/hV90B9LKR62wjynb8r8Ew+/c4wdtn7YzZS/UFkjPSAYH8fyT00ffMrM1jS6ZGnM0j6M
mNUCeIttppfTP7sUSF3x1IFizNugiZIlJ3Lrjx9f9BBqs8GZA8UY+UjtO6CU802ygyZ3IOTWpV6A
dh8pX0hHPRA70HRqGU9IcSc3Mq/lVcG92OsddC7mqE7jus9x7z/kKuoc0ACZ1nmhxyma/AtlfBjB
mtqQ+v2h6IUXTUafSTghKYPbV5FqpoCKsQ+yZ8FYX4Zkqjm5vt/mk1JXq5vYUDzS/TNwn/BpR0HP
Bfki3Qr9Vnb6UWjeTCJgDuLt/63TcqP28jCm31Iw5W1KjFYhx8qbYgQDrHq0YWmhpJiaCmn4m3nu
ZkYqJfLkcyFfD4k7JonG1mSXnSNWRNTm1H/y9E09b/H+w+z9nJKiV0jko+olOjtUQf28ajAh6mzZ
hQMOEu6W8vqKGdjjOKIKugytUXjkgxfOhiEE6J7Pa02tNq5RgnE9JgdfG3qAgu8Ny5g2wa9c6snd
jw/pISOGuMmJ6svqgUzZ+nrAq2nGFo0mFmg9vUTt8VE9R//E/RpcXBYndEj5YEOZNCq2jtQoXrtL
5v6MY8zfCKiA6fg6KJx1+e9Q3Yy82mo3D856VOyUEF9Nt1N1Hjl2JYhWVAdmUR7fz/ktNCioA2M+
Y0rOkPcP01T2LzNAZFidadw3n28rP+OPf2m71Pd1Wx7IZ95qJA8mMxkUG15OWL6LQm2fhkuz9cDO
On7Fc/sUFhHE7yxLfj8avM6KeTPqqLjw/B2s4BwVD97omFJWSNfPkr/GgdyOlR48yxNBsCO8xqg3
3Y0UF4SdV3cOQfnrL5D2nciUYRexVn82Df++OWXQyoB0zF+jPo5FMfVKCUu3ogmsxndmU7ZFbwSJ
nqVZRqQ+8vCccV5od0MHgadT6jCRdL+OjE1FIzhizAbmHA+8Nt2vAVtdQcVwe7GomD3Qjgq4LIoO
rATa1OH4Z7sOo9occwnqpXCTFlMKJ7mi5L2qgwpdTZkd++axBUtbr2nizp6aPvO6JahW0sIbBmA4
j6ejUOGyPK1WHmfZv3+3HEJw90tuMaYxeo9vPFxjEDmtRsoj5P799ZdZARB5Up9oD+h0PTkqLMW9
vPsoAzu6SJz3PE9yjNd105B0mo5EzPxlb+finrLogGg+GaoZlqU78WNONRJ5ZJoQE/FwyquX5UWj
Ll0hbv8RCVK7w19p5DJ9QbrROfCdpKCKxTaOHGkRAtuS5PFwyEsFEtuoohaQblsQu4UEOYRSGhNZ
usNSLpMeV3HwkkDDM1ujTrIHIR23NzVmUpJDy5szNz/ilI86jIx09dNv2sHTw+bB8mFi5Vu56a0X
7gynUBshIpRMUILSin4FjIS1+zDzxf5/6Wsxt4kMVD6vWi6d09xfWhRYVDrkp4/J/cahRzRzWJ6M
a6AoVDHr3q38nypmBza0TIJSgiRz05TsF9jeqNEf52EXtmOWz3Ul1IR803errkZrqz8CK8iTGT5T
fNEU3fstzJmrFxPYBdKJSNa1JJqeyofaoULVjnj3iyorl9hPsJKT9wzSY8PKc7+pcjZJUtYF3WQX
nJ4hYhR4PIbf0fX/tchn2TfjKJKzc79IFoiptaJXTWvTpmBP5tW6AFmaYQolnR8d8I1+1joytVdB
3smId6YeLm2fm5NNiVKJSXA30d218TQdxB6a3JZebrzLZsPJ/AL+BpJZksiOuCDGs3QlQm64+nLX
c6fTyB7VZeAZ5tQysZFj68AIX625FoxssQHkhGAC2beqKbrhKTql8YaLiit8nZN6OjkX3yHyRkJe
7iBM13SM0nzE3AmNhcQONECilDVtoph32+ILafg2Um51j3pBg1KU4EO1GN3HAEg5gq1MgD+q582u
V+un2b6eVmgNvT2jXrsdJns2rsY1nu+ZZWHfJDZ7f7FdyYKc77UKG5Wzv9bbUiXAacoqfxsztkIH
v0yVvKgQMq2H4YQJXVnlQgAfcg5+yLmv/x9ztI+ZaqOIjkjRu5wc0kTp1F5SF3tU3J1LVmKyIC6g
joiuOLxHIx+yo6pMsNBy/R/zd67ltKlRfkI9NgcrpCpjuVv8htb/dixjyZmIUi56Z6fVWNEOLC2o
4UvG7HvqNXpHfFSNhDxTY/BB2v1ymRhGCFPdIHhPIIzLf+3G0BYdluH8bMJxmu0WM11NEXUr84Am
50/9Wypuq7DFEAkKfJiUTcJVgiRWuZToBac0CxJ51MHk264hfsHU9CuqHaZqOqUzNRj0VqWvAjXZ
HuloxsOC/WDPzVz708stAmQAK4zyX1Vj2/Q9kwFhKMYkdLAjJlIy5xJCEtVZaE0SbnRaNdowuGZZ
5PUnxu06BB/iEXsFb11o/CQiUHQTfRXPsybdtldXhQOojuvEPuNKDlIbZtjum49ZhjuVAYFRBigK
AJMQMiQEhqP6QGa+01VitWx1E1OSZR7QaEo9WRVoxl4ZuFl4tAVXr5H+u7r6QSKJjNaKxUqMCjC2
8T6MqRuMJbPFMSF14CQFPrS/AhBf4ftRb6hcJXuRsWzwkYpi9ZT02VKQUhivyI0cqkVdLWifBDRa
98hcH5RmG+yA+RYy/4FxsnpkXMUM4wiI0v4seUcNTnEpzpKrVH+P3Ad9lTwJGj61xp32PkpIGbt4
mdPSeqp40CNz98vWfwRtfB/zH4HiZQYEnJCrczFdgcoxEB69dq7rC8vv1+m+q/OkpPl3kmJlWrMR
xdt73TjD2mwGaa7a+5bVdJic79cSePZ/kPMLRCX8fr7IVPHU5XnGo2AeLC2I7LJStcNrB/5Rzcz0
eLvZ3oR+gxY66tbl+HKToGuthrD1pJ/u/vz2mOrhEvSvvdnlEjpIYmlVBcY4NNpPsSfE3XVr10CM
549ZqFvCP1hyTvfCideraO4QRJUxaUTAPrTXof/0F0bAytSzBaDpioIDAYHSOh7NXTkNe7VL9tAV
7hIqtuJD9/JKnKzmy35uNnCsN4KhDbSu2A/s4JNIWkfcPh1aNVjtp0IiY+qA1Hdi+Qt0qZoDZ4JT
jxDuVDPzpPYM1VbEatX6MD/bLCKlYRJk2fl+zCYrsWd08aqfw4TBlRNgz5ULROHDYKZYVYLHsrLL
wv9/RAeyc+ag7gcv4ldefiQBMDZYmKyzMKKX1DMFocexrk/O8888VkmWSHhMFUUEddJtkfYkIimo
6x82ooMNZWlOSQFBC0/nDt45lah7yUiBpzyndQsCV/Gvx6hz7Li38ru7Y4ePzBoxTgJlkcF9BhiY
XQoAqCllyPxcM1aahEQmcG8DyUTtrvttmDQ6IZYnLs5YazOGnyoSa64TmHfIa1f6oQPUnV/2rcU7
67JBHczvQ4tdrpu0tl7uRTSKH0WwRk8arrnvW8NbAQIGohKz9a9vDv7BSuYcylw5vruNjRHxtVDQ
H8t8zdDULNPIZh3LgWWNIbdj1E1wuMk0bqTqFgHfuRuKX3I0wRHyK1zqeiyYbCv04+1o4mNaL3is
wgTkQTrSA3MZlbo/4bb5X4IhvFs+h0OnFDldEyIxLhd93dqJNZa0GG5PHa1w7trefrtVOoJwVxN0
BYCKBvi4rJHaQyXB9Y8jsr6fb6DFRv0Ejo4/BpDmafABbqUicUIm5TtAk7bzWPsRwWQZlDIwDIUU
pQKKsgmgNi2VZrz1TGaQovIbMi5cbF77ZJKyMABauDfuucQSW3iLhQQVHcD18qsYxQjsqongZ7t3
71vR40zaMBB0Y6Hu7c5UiAfA832JDPCvUPKbm0bp6fdHwEFTlrmU18/EXQ8odDgpSRuiwtLlgwXC
yyrxnuCu6lhKDpqD4ktKW2lseMo+UT6YnVqmCwJB+vQE/yaEcgPGdpxC/4G/eKkieeClYdgN6LV3
omgzykg2wQg5IRr6g/rk2diih4730PoXj96tlIJfGo7S8JL7Gd3OPZ26naLbCmrRXd7XlflRruZg
H0tj5hDABa7HWPnOP1RUlg+FBbubt+KNRnbu5knAUPjKONIHbkfF0lBQqIiftjTrdCgdSv9oa/Co
ywRdOmPmpeooX57FWAiCO/jp2eNjLeuz2j2ZVpjWzGwoWlxYIYz11YhNvv8mSuHk1EoDh/3/F2RF
rCii8UUPOR3SIgHDgs6tvsHePL4yxt2qoela3hLKR4wVYyeWp1i/06LEAYZE5Hc0NrX6aN573u7W
jbpD4EuOWpHmGGbHyPtIeYq01+PdK5lQ859cMViXjCSTjLkb1Hu6B7UnxxGVcgdqERCqfzaipgbC
HFYbyZFe3IkZF7L+8xxJso8/CZe5yUwPkbUtFFgozwtZUyZgABN1gUg4YRoLagEkKZn8dE8rY/rr
AM69G8PI0R5P+xBW0zVSA6UouCZSP5pMLl3xoK32Q1w6R08Oo6pB4nUvRZ9WHcSYdP1sr+n31I+Q
kqmlx+EzNwsqcL9kXYIhgql7KjJY7C6TnCcpo/daMsbGOMlFt85AtuEi7gKOOkBaLt+sv7BmA65o
sxOqW3qBd176YY+zTZlK8QKd7dNGhG11Lzaa+dxCCzOpQ2IGr5px8gwPWn3psj8723hxxNL5RVHm
9jlgrbGFPUYwV8CgqvKNbyQWY2zI19iLOf0ZeCr25jrF/I0RDy8dJQ7vSk9IZ4ksg6v109HVQpK8
bGNZc7/3leud61MWSosa4TlvDz99K3+bRufUePyPoE0AqONQl8xq9TKG+yESFVXSCPmpMsLK2Jad
FJXeW70ZsnfdiZSJAMJhV5B0AONurx6E7+ThDkdyAHuObzer1Wb9dXtv/IuoJCFYv63RUb8HYJQF
WREjyiA4Hyy7Rc0PC0xre2t5YdzWLmbUofcZ1jep3XkjlyTy8FF2qpthl+H3ZzvnMARkJQwjwG+l
dbza8DiF3Jnl3Tv6jpJCIqfwePRAukUDKJ+tMNXdf9x06bMQXNQPL5imm/4VyOCs01BG1V4mJXUr
Z0LNON0bqIjfvx7Q1p87f3QUxygYwlp5705cSedCwNNx38J8DecT9Z3D8us43bg4aq6vspwpFEtq
bm0yaL2KSwArEBDIfHYS+VwEyN0cP2uPyDZD+WRcCvAPT6dUL5XAgsuCVycePffJz2gMaUaqVZBe
XxIWa9c8s4isGT7a21C/MOlKgKDEp3ogfh2yArI26jbrFrClc6k7TCQmOLKDdF8vFvqfoGMCwTbl
8EMe7IyDTVN3FjtIitfeqNdV0gRjHytyJNRL2o6PKmIFVhU5Z45vRxkHLTOBFx6YKPdbypdefw77
tei4LTfv0Yjn8jHkSxdyv8kWYdxCeRh0R+czxo62SVkoQjv4y87DimU3I0dPZNOvoys2odPOCr46
zANOoG19txWTIEMldS6ZJjUX+lG/jQ9tz8t+D3WMAQU8WU+FbrX4CGWP6zD9v0a1aTeiwcaCXdQH
TGisRDGwqgST+SoAJXfuPyZcw4WYwIpkbPa+n/Bbp72TebSiECN4B+ksDMHQHS9NPVKqtscD0duZ
rZTGgV0Wt8eSeaFrPyc8oLwcN1MTRAy9dc9Y2tBVKrrDJED0DutFGM0K0LChkREMZcsO9HD/oGX6
3yhqwPRyIxHnxhJMMui5/2H3CGUf04K3/tluzccD8eclg18IYmwlwmmZnU9ovxNRP7WERSVaHZfG
8/hTNE+vD/Myu1hA2gyOBTZf1SiCttx98Ygkd78vzALclYU6ZHvniFkeb0rgpvBbBums37kWJCNc
QZT01QiISW4YF3s/hJ/lN+65ZcpoSm40b2RndiE7WIQ42AgZs7FNLcPve6xAWHYXsfAcxDo1AdiW
2dE1Oux47NvLbwvFDR2GXeoOCDPq0jVPAofRQkPkOvhCcvS9M1HX6AHSB/z5viF7IxaL2IpxKSUI
yOT5r32rzMzoG4HpEk7escgfLnYtEWJFYf0zc8I9fNxGhg18lYoch1zzVB7jljl+7oW5mf3qPjRA
vk3enJnbFSh7gl5Xj0C2zpwhldzjrkLoyE2Kpz/OE+butJjFWcbXd+kiIE0nSZeP7xH193QP2098
NmDAPpSuECQkz6O4uthIdF+mOBJB6OWK7tiilpwZeiCajFos9XV2GN2q8ix/YP8ve1eOzt5Q6eyj
+pqJCpWDZdeTXHdwW0xQLhiJUn+vJB16vBszZ+19h/1qZZXrhkampRkwV7IE+vHWogakEgKuaEfs
CGf+CfKVyZHpErVYbnEphDITjYZ17jMeJDL5VkUrGoz18CIfcjm7n2oegZWJpf6XGuX+XvdKzHsP
vpKAMAzQcGJQ3ayhGD+pf4iq2LNOwDF4X7hYZLf79caJ1IIitbMLl0/T22hMy7rbr+/IUamzFxSS
KJycfN6vThkHcGveBFZhx+eaKOYCZqS6oBed3YjGDd4i5Z6Gawr/1f0DU5WCpEDh9eqipFCiujrp
qKHaQdmoTqV4Hikjyutwz1TC8pmvWM7+DCHztkD1y4FlYoMMq0NVx5mkqeKuwF2lvosdmtxTminV
Rc/pAe1UqqvntcY4a99vl6rU3fDxMImPJ6vHJPMsbl7IGTNz9kgWv2qkml2A1+1oZ8oLh6O+/odE
D19WkKNQzcxAvoBQbPaOgYz5lQNwSa9ZPMahFS7MpzKPfrrzBNiZmZx0qJgX7VV6gRgEyIzNTWvo
Ggn7bPRF5S20C2BKNe3h0CTzlLoYB99KAqzkcBRMb1w0mW6YVOmoM3xa+7ZsWZy201G74+jjf6F/
Yl1RNl/oa6b8AbRSpd9Q5vTWFXQSbqumIWICyJ/N+crF4KAQyMC8lUOavnPvsSFhpRJ639nKUXKQ
cPURbyjNm7AH2i6MsKn5nH9dZkrVYYnyGDkPzJt0hFl7iXW+ZpRI44cWlTgnqcpIAZTyzG9DlPFY
lzVp6q8rgSVNuCRdqNDnD15Gr9UbtX+zYF2eHnHuDsPkC5M5tBOG+mUIi0kvsNci1+9bn8aF9bgV
BIoSFZa52suXNZ4ChDU/Ua/VP9SVHRwGv3dUj6lkAfeIJqXf+TuUpq5jLTgtYfG4YOG+MAVTbJse
I3vsaBHmssdH/gEcDa7caz1AC106yTUjEirGzyBMGK5dHhhkMb83pogVi1ghFEN+8Rf8P4zAIdW2
TTXaNb7TphSKNT12KOgYilt7TUZExDELCYcD7MnfValfsA9idGzUkH5OqJq4EIqG4iIrglsY0AKk
nmRbSxKZ1r5fjSuAzCOx5s1rvyG8jg62umfFgvmPbZJBuSipPVzoKV8FTDGWtgiwIsDxkKCZ/pnM
B9mwP5Kmk3tHm22wrwdwRQCeklcHyBQKQDks97esSbryrRQ/SrcAETMcasyasvzYPeW3inRZZLRi
h04zrzIHhf7HIOUFzphR7jj5sxUnU5pa5vxgY6tvkyk2b5ft7s+nt9P8LvXYDJK2xLI0VVL305l4
dBYDiU8k1RWDECFQ7eOjP3JvdyjZHgVa1pNvcl9aaCy++dhB8BtXaJi294lDC7IWXOmyFbQ7nF3i
jDyu4t14ehtqAxoKz3p4DS2Z/2RUZxB0E1fBdBeANQ7Ih/aVMHMEmRZD+6nHP8PJhjRD/BONpkMc
byQ4GgBdE5+wHwSCX9iq3hPIqQEEaLf6TUEgMButsnAsSz4u1Hg8rxm+8icaFmAP7tC5dfT2pJPF
I586ZUhj/8x3/KycSL04y9Dpa+9Dw7xbTeq2HO7cGy6CPbIptWELxGTyhgWkG4lFtbcNvXJfBy4b
EVrwCsSyAnmCYt8AGMH3GS+7vCdCzH4xios58DMLv2/0t3wf+dRNFkP+NC2zRz+2eobhM6Ox/grO
Izoqz5Lv+rs2FTApHvM2aJDECpTreBWKnfUaCRddohUtyVFMEmuSnV0iDdBOUS236vjJR8VxuKvH
QWIZtoT0XtrdInpZbTX0kT6anTDv7n+0aVZ65+REC4qzZkU1sKB/QKP+kdvD0gUJhOfj6is7Hytk
/Bzfa3s81kDHDNOd2+dHqGvOqpdoK4AS/aAWNSyt+0YlMqMb7yg6wJL9vSyLDi9ahTTFXlrJM9f/
NURgV3cHovHXPcUMzUiI9sOkhNh5980x928bsZ9UwV9n8qkov2mq3rCg2SkJdm+BtalvzzmnK+3Q
5m05UYYpfpje3djYa58oDKWXxE+kFRc2Cd+IbcuQsdIvssmX60SlVOwrbtCjidWzqNjRZ6F4bDNI
k/uVtUAmxoT/iM0OY7tYI73h8pklloOJbv24suYbjqjDBcr7S3Sbpdyh8e7qTOhyQ+/t8Su3Wj/W
S7YQ/Oc7VuA+C9i0YNbRwFoZPkKXFFJeNtQAJwkVQZQoMnV9lVqwHJnWmAo+hBSoiQWabVILn7Iy
7zAnJ/WlwZr6AYBBHL7rSathWMuOrv4pdhlsALUTJkgVKrOyoPJZQxdw28hiVM/RueSh1Uaj8Gfk
gTLYczGNb2Jkvfa69CjTlgsTXDmcOkUf07YBSm6dUV0kMsDSmRQeZV13OchmHNaKhg8VCVRdD+Zd
lkIX6Pe4rq2dmES8e6iekb6oAjqyEVf3hm32IA+STRmTlMKNKY6eLiM3JCTgY82NWmBLNRCr3bXp
321KYi1twLBrkYVHO6FIuRP/+4ktWQU+mQJspzwl4MYus1EN7wOjX+NKVX5ErSu+LSy/QpPXZtTq
EW5w1AaMsPN8nfyWTXjxSHX3mIR34cd7SaEGl96Oha4msdlP6C3U9MzTWMFBkNN5OTvSS9j4y6rp
/VbAPQ+4YFJC9ZQ5amw5yxnsmn2XFDAFMNMan3oTnqeO73eEH2B/Wc0Of1/dRMWk0WZ2WgEqsCz8
cqpyVQI+Y0AXdiE8VycnUDOMZqRchXzSkhv0nBxQcftCLIlGco1YAKxE/i2TusXzVGXakTHtegdI
lg4FccUBcu3LgDqeeBJHPLgjsnp0QLjTRHyOBSzgg0WAtrjERjX3TYXdJ4z8shZzRmEzlN3D8CJY
kFkbHfD70nSXOO/NmRhJGhcFrnDzPzS37G1to7fT+Wjl6gUCKkao9HYnZ3E6d7lLFU3y6GWaxIdn
1BtAf1Aax52jmbSaSgEI/ZriobDvG5+znxev7RJ25IXeFxstfIADZrKYtyD3jPpANCWg0eDVvzNB
KF8pOKMqvJjGYTS13d5GApCcl64S8zEjU7j7IT134ryP+vHO+pMuOYi1TZK3OS1jPdLBBHAJ/sHc
L5vMTgdNxhJh/JFCeak7HsSeW4FcmC7bSdqmMzm6QYrq9ypkO45HmAhd6iZR24diq+lnWPiI9hGg
b0I57jUbMU5rXY9nSZlfd9xACV9p7U3ao8Opvy55qdbYvGUwAL6LpjQwa2EfqFmzYUc1ppYdsrtf
2TJLN9scui5XjyZK2UhY2Pr2E1oxSvjiBQHPhC/5bBNV3zDMndN0DjEb/NDj9KplXQmqHqw+unww
APkUwoKIMODRdJdi+Gr86qsiAMkh+92SEuQX0Ovogdvv0lwXk8+LkrjBfkh8sSYPYHts0kqnIYAw
N7cJcrlL8NbxZUJ+ofqTwEjWvW1oQN6lqcPUWQQV+5R7ieBjNQ+75SsvCQO3QWPNmVzp+w5zwg7w
f98pQ/b9YOOGeA9dN9sBQt02CvQ/kW4LKy+i87JTg5LqHZ8OxmurYi83SO1pfA3rfiZvrToWuij6
6EaOMbTeimXVW6wQZznN/IcxsJUenpidIbU/Q6PA0Cx5cSfygzma7vPZmSF00W/gy7k3pLCaMmXj
ZFwNrjIxgG0z9ThMU8C6k2OvllvNvVYPVu/MYCFcEzsGHq5OKi62+49MTFa0PofN0fnp9eHdSefi
merd7LEbok5FvUAjRbGeGydn7SRgGBxPvDqZJ2/+FmB+82qnxpYNb0D8SitazK/57ZaNiQT0Nlth
Sv2995Ib6Ic8UmpE9lpY+yc3eR4KuGQ3SV2Y8+CRnWiqpXa4jZJXEojCOwa+5IswwCSbIDS5mIP4
Y4e4aeBnkR2HBFBjYNMw3u/yAMkCwfUfR5QRiT/3J07mzohUey4RTGBW88wayVONJ46HrUt4soQF
AQSO3Ghn+UkWzmN0wW51iIgu5vv1CqGO3sCXSHtZbgOzZgbzxglR8Yt72QX91wM50yQTk2fh/s6r
jbIwYywoo4W0DrG7iczYvUyVBpq+GDLhyqSHvDjpQ/P/zsCUg/CukscmW1QodKj1ULkwWqcZPNyx
HDI490UYzOO5Bd42jNAFy4Dy2lzkjPbvfPlwJlkr7WEICyjNCDvRX8efF/YB1mb/THHym1x96ZYp
0OufOg+u7eUYLCIqaD99C44+BAc6i7JRxpxR5z1rZxUjpSLuoaZiDbzEWT/ZO60tKNJNOG4XYt1K
dy6lGoOhbuvqtNey3/MHmVEyrtH6jk+msEd+ie6taBiEq3QwKUByBSW2KaNHXa0RoFZaetiKnwLB
6VTmLB9KKD2bGaEh5Rk7lBSoaxnTM9xdRYsEj6BbwHmNPyqQ/zsViKJXA8CNv+e9wjNIepYF0Rxt
12n3yOAwMok90d6PIZRyJE9J8QvAmRtKKjAku+lQZPYRyAiuGxPXb+qyw4Bf5zKareR73jMGKiAi
9OoeQCLPB5LmxfKPmtbe/r6+I40hagBEGDJ3hPYRDjJjUru5h13cMrw17RQ3wxx9mcaLr9K6a/od
fe8G6h4ieQ2PgcEQ6yE/ChSXW9FJqDz6lHGCUNOxq6A5F7EoELPecFUshwDLmM4hh7dBdQheBK8u
Jo2gx1ECcgMipyMRhPSPUN3B2I9zE0KwXgMJ/6hdCawhGBJpdGhhW9GTTBGZlvFQCtfSuOIBS77M
+N/4UlMhKhGbeWBCLCPz2QmBhdSGPN64Gg7va0znE9/c7R9VLSkoCrKPvZzopSivk4oFIfkKcY42
noEDanPCMKyEFKeZB/It25lv9VPu2u6ShmOiBsxVF0ovB10KsK3J06jD7P3yGUGZi6QPuu02VxiW
YL2FlFR8ig0O9ajAUcudf1C5qVC4+YK9pN+n1f4nCxywNUq3iMvKfCdT/emr9oqxWuFIvYGRxB+Q
p60YijuU63ExyoJliLGtkKWWBr8GlUuH4IjrEtMQoFFlwUCGW7AC7k0NvGGcloOI+1/vqgFXtT9G
jkgH6ZGan9yvwmG0IS9t/EmMRwfk3lHRWzlRvk1H+ho3+hLGBLzbVDhtpT6KFQItkdO3Oi7cj6dZ
yUVpEzhFqPa4t0r+zIAhkfclCGfP2n2Ar71juaQwl9m1JI362VatM0CojDbc0tDlnpwjmJmpXyxS
d4c6pwAPOF9ftW9Okj9oSmBIzTCIn4lqvwx8ZkKyC0abE6/urKsI4O802I7Qj1nodLLusza1VrIs
mGn/sOeeQU7tBUY1J3+8gTma9kFTuJff/8NI/+MHxm7QKOj9vkHT+H7AAr8bG2sLdGqlw9aGXRBX
IcKSvX1aAinvujLRhJUspzx5kRJI2dSpDrJpk02oSaKr/JcQ8fNQnXfV90qK7+lcERpQYxWlsgry
QwT4mpwpXlHPhvJOoju9hTKSiHIHgbKuXpgD2zdgsxTGeFlStb9du6aUUD7i6kCM8+DrCLrhlEfZ
Ol65BkPVz7N89WPyhHWJdr0x3u4jEfsrRfpTw/mooZ+VITzj2OG5n5GKshWzq3WGm5+Lgvgmt7Tb
y13+qWlg/ajRg2LgDp5n7G/wJtkbU61hY98wQ09rzPYCsA/ADAwkIarcgiyLaezdlTj5A9KXc+qn
B3ha+rKamIB5emV8o2HDCuD8e6+M9R8g/YNNxphV4mChPjiUM4HaoxMqp50LWy0rGoRQ2jIoL3Nv
maqdwPveNp6dJ8A6GY74iVXjPWDaugXp8CQb5PW04V1IYP16XEyDQ8swgGpAraQxEiUL2BFVZtxY
u1Q+kqXwqqwCrKvGjFit5EsVaf0eKxebDUI3kA1qRNMwbWggOGUJAgCtANP8tuOOWEU88zzEfC28
dAyqWHMRl9PFVpfZKXC1nDwoITQgMJMGGXbwzZ1RB97LQjgD7/bnPfd3qBmfZ5s7oHyZDf8kyRM9
Y91lBgDAMd+GJXUHKWLiwoUenjcUJlET821+BbHA0F88R6au0P/E9z/tNQXjliBWiZ7wDy7AR+VV
UdKjX6kPaIXf3MU5rt6aNKdiv/wAWS9c7/X3F/YHlaF7B8T/JsrxnV11WX+TXFaOc0mk+qIFJf5N
k68P1ansIP5cP+T+GmAkIwtm4/XQLNbQ/V1AKu9pRs8U9nEMYWcyGtFuLAaaJMaYnJeRhoUkB0tZ
g3/QDQrmbidfOE6xAM7q6/czMqborXo4VjI83s40hrS3YqBHDsKxIcv7P49YI5+haANxf88I2iZz
D54tGzZOUnqFYNJjwUPIc+5wSpbnITgPBFWlYDk2dhlNZouVZkhYVhIHvj0jNpkDBkQp0wgcrpQy
Q09SErRgdq7tETbQCmuBCKP2MKcUdReMJ+6+6eNu3tQm4XQPsFs1bI8cXZBr9RLJ58eu2EORCRsw
Q7byZuJg1LLeL6PiSAgLk0Mj0BbMpCMhRlUH8AeI2ahgpF1sJrCdN+x0/BEd8JHfNGFVQgtFesXW
6nS3tfJRuY4zFP/t856K5RY8Pv2EzRuVECVC0Lfl345uqpS/m7ZzfSm722LsKur/ZRYUmOL+rOzP
l3N0dCDbcQvTy0bLQ95bIy2nnBukQn1dN/Ur3githA6kzgIrWwdZpnbagccaFOJOzCisB11huBNx
mu5KomI8R2DJtoljwEP16Z5kyGLglBD9xGpHQ20pT6mNrbF+IglDlIbKwZhoYzI5Av9nZUxIrg/H
+nk6OT0mLKZOiTOHFrQfxRyisqiKsoevfXndDB+YDwPrV5lqMFMaKSlvGyX0oUNaMlrGvwrSmjKH
MhQfrPtONMdBW66JwcS7reKb55GoSDrBI2dr2bEi6NT6FSCmCwnlVPiSfbdbcvBizDCu6dI4MEvM
HzMVYsas8sdFzg+P2qstEEMLZDhuaNM4E3ynF5NONwLj6viceiM48rSnXlkcwUg+GDteri3iviTX
3UMrGZL0e8JZKWWRNFTjZw+/sW782sG8iM1g2e6HY+uJ7H2QJRT9gXvYBYt33OneuGwdI031j9oN
04nc3BwsNokzZusRboJFDncM7C/1KEq3p9fTPCc4O0nzdt1uEy4iODYWevngYlRMsI70Qpr+qZ7r
UDVJy0O+u/kO7Yv0JLrGZUvL6MgukBFR7iNjWSsnGHuQYSRQbo8Xznlp8hVJA+nsN54uZDG4y03p
/Mmj8kfUgP/WKyNkkgdFqSN4QVEa7ClP2XVOHzcKJY6RBeBj8Bx71zcSrdIH5jc4IHYwMDxKhmBP
b5aV9Kdaq+XGut0PuD4HD1JUOpjrcmUh8p6b9jYOnVo55Xqy+j6Wxfv2wXBHftA1n4zqUsvcFAF0
kfuJIMWKVyxfULidfxcJeY3x+eui6FCKwi2PdjYEfgksMYlTTt8fyfI9/6vlLVsLe2/TTO4xscPO
Snmc1G3biYk9sm/sYCv5uj0gtONHv+sxDwyo+2AFrH2f2dCArYpMXkHamPU6qScx+goy1mdzrfFD
TR7hpobAD244lJPLZRK0nLkCH/rjwRSgk9vkCutskE629IZjiDc37NZXyh7c5UL22rg/aIAIZBQF
7slnIdUtL9pBkHdubjW7Dz3AEOJaRb8qo2BqLgBAqrmxFJE4ott1dacH/7UWOYdBNKbNIFwTLszX
2up4OxXepW9JViXQ0oAZDcayhyXRynE3nd80+LZ9Tc0ySLWqK7ULeWJRvMrR4mjDjSUxM9gR7bqe
Vmnl+oxW+WcMRXeCCakj/PYPN1w/EomCQIPhhGoeWU9RBAfmbTkZQlPq/FCbKZB6YgX7C2D9w2I6
a5WPnoBxKNqKfCcyAu1hYTDBGt6tPcgy5EfCJrKFvUsZHmPmVHXV4fqbL7/83t9+bthg4n6VieR5
hkpf5Y+i0Me6uNm7D6t4AQWF62odAHYl+T9Q0T0D0zJx9cuNCqjtsiOxFy/ccbauMP8OBveSNlqp
w0hO+kWHBlZW1yh7bLBm+yWfNjwP5V4kRZxEIRYedO+Yo7oIQ33atjN+wvJ1VOMDG6VbC+LJ7o89
5fct7R6bm4dkTZrhM5EmbisZuFztvCtt7iu9WLkiMH6i4JbvbFC24YWapKrEZOyoIoTz3VlsdBIX
VJ7Rwm1X24h4S7xTETI8QdWheJUeafcWw2kQvcDsa295wpkQ62kBMPbMMP2X/ggD8VWRsUL99df1
NDhxDaxtAlUQD7G/PdeqMnOCwoLczD8YMxuQuC4IxXjfU7RZCKRcqFLpz99oYO9gAf0OjH5xVKwH
XtRHj/CQp9hR6t3I5rMxOFunf/aMYKZSwThywZYvFgapM5G8FmEMBEUK01bZAwa2rXEH8nHEN2bv
7rAVtHqRKS8KYEs8u0sHI4lEJ9AECHJjVDiNHFvgI/ZAppGggGqYkw5T9y73hO6uTAGgZG1vCATq
89qye6E9J+ta59js4/wJsqAAx/pkXjIiF1Q5bVN6Gl29sC2RxKEQfAiVA+YU42Cm8kQKyZMygTiF
7giWrig73QlDjck7oXw8cnHErVovepoM6jnHEqHIFsbsm9bUVR8mnpFc/w045/amb8FDPmVpiwNH
tvjuRt8NxQNZJvCVHZyRbHpHph836Vqz+7C9Y2Pv+0ejbN30c4Aud71GV+k+F9YrzWuj6gOli8bz
buuZeF+1otHHNnBUZk3Kv0jmXedsPJKU9wC4Zs35hqjMG8RskUubpoHfkB987X+WKHYdRs+aSNtQ
PjUQyXASQRD4AX9M1kej3jPRo28mC1jJN0XRH9tk+FN1CRAmh3H+2rSHaFI6/UQKTjJrcJOZjFtD
Nw7fxFtJMJfcpZIaN+eb3ca0s+4yZ92MbeKLRIFf5Mr8eFugnoJXpSR7maWj1+E+6/Zro1UegxQ/
nWgNcwIqHqBYEShabx+1TJIdSOhUg0J88f8Vi2YSQzaIEyPpDZVDH3h6cOsmAuA0Q4mxZpeb+HBo
Dnopa3W5EUCcp1f84Oop20DZckoIS4Wwh8mDOEKVdT9mK9ztZlOnesef8GMYWWgBKXxjUMosPR+9
bK371eSCQb0aDAX/m/t6hIVMjkXbA4+pwat34WUxAQ4YHwRzykxSdb8mHn9De/KcYRIVrAnGrBh+
ljZo8tgDf5XkR+IV4yDdDDmMeVGXJ4u/Dmfuq9L/gCmCTC4QhSTR3yPYbo4mHhgmIYNdO6V8BDgI
B1LCdm0N5d6dMM0pv9ZqlVSVCkhCLxyUF1JpmyMww6oBwkoQCGT2yknXF82ooZj6k3qifdH1BKUZ
6lRGy1X2xgM1PU5Lm/9kBk3j+XU63atnWGOKeQWrDcKnTJCajwNXRzKhSyLgyVYAeLmf0RkQ86X3
ettHQ6GeDwl5zr1d6e79KmCQBuLWbvcRnNZgBh80sEGXmCEDmH8v83ixv3Yo/goUX3SbLyU/TJJs
70d8F8qoul1nMVYpt+DJiQ/4a02aN+pn6OlErwQ6tAea3VE7mIzTVpb9Hc+5s4p3dOw2GIRaV4Kd
qWRUKsfgl1lwLwnx362R1myQy0g1Zn0MetfMKDhrf1uN40Ix3Auzu2mWJAY/qmtdsmHh8uloSymv
ahFma+JY17TF/e4GqNTpP5aTrYjqDgeedutfBxJf6rXQtMmUktlTLTz71dpQo+i/VZMaMjP0oYln
JJzpo7uhf7dmKsj073ZcUyQR2JpNiCOLWv3u8lVMR6yGBE8xUpz0ncJbUD/A5CA7QVMFWiVdrnxY
YCDGMA+dCBck5hi1Nxe1okjUSTYdXpnh9Ddardgj7djws3ix6w5x0dqlkuk6Q4Yk/y5clMjnrKoj
uejwIKUb5GlsOjJmEhwLVujL7OJMQGbtvtqat3I8WWlIeGsxkUukEbLz70AmHB/sEqpew9nE9fVs
PH1p+VS4BM4v7iZXfstIOgpJt1hihkM1iiFYb2/+pvq6wTNJYaVJBiHYg4bX/e5RVJ1/A6NI3P7m
2a7hzpXebbZ9a6rNYHnqZjMikWldd4tWMVESnqMl4vGEP+weghUKFyHhkV8MwnbspuLTymwL73WW
XBftjVxD4ubIB2ANBqKMVzjGkIYAkJwvbzucPYA6+g0O7RYZJ5mqOdihUVc5TA3yJF+J0KeuZJAz
LktpArJGbJ4esG1eyiHIjK5P7TfI46zurl9usQtJV2xFYtVETU7kKNRtxI4dGjNSSndaq95MZvc5
7KH6aA9J5C9AHpkaa3BPnp2JjYZ4/1WnbKBSQf2rswUFLs3gSxg9g7YFLeqJgY/6VVEz4TPGpXoK
3DYiHwJ6pF2D+7+jAzIWfxMtjCiWdjBL9N4Q2tWxRvfRMk0TPTv4D8hI75svZsKxGa+dcfs178VS
kzoA+4p55JKM5+YQl9smB0FzNXq5NZoqd2ONEJapUv02QB8V/qCJ6gIJNHnkuRlybUOsd7Q4vDHb
vS3CDPMlkc81JHo3dpVDWRDIQMzNfS7cxojwvBnRuvsKlFLg5PYbIyIsh5/MlmPzRjMURK6BBIIo
HUSPgcjcFgCCvXDXnG14lcWsWnO9yDOn4xqg3qqSI2dEHnh+omSsPPVsMe30daAmosq4ax1CLmBX
8QDtG/PfTJ5XVLopvMaSZ7Mx9S1Vaglo3ywLE7x8+PsIMyTkoUpHgY4hJkAC5p6/bd7XjR7ABTOF
+sg7cOL5DPzwwob6El9DltD1A+Mu2A+6NhoutpSJnueXbOb2l7PvNNqKLwquSahiRRAdPD0qrPiu
PgRE3/e5kx+C8eIvF5NEZWNP0rNcbsGDlWoM2atvYF9rRhPUSobSmWN7818Pl/jMjsJWGjcgX4RX
HD3jsnk347AR2JhKLa9p6tca5svOLDiPX2db1oFNCRJeAM577vrv2BEvl2G96I5G52k1gvo4Xlsb
ixtKBHGZa1pkQaexcY04+JoLtekDh3a/jDxDLxQHjpedvbOoFRvGdRtxj2N98lbT7AZYwN0LwhoX
X9xODhYYY590vX8LodiDIZp2+g5EOTXLfDqjO6J49yqpcS9eoj0K3BjsurlHeqn/ezgZhq3fi/eR
NnU5/xLOksVwbHU49c/PXRXZ3I0xlxSD9Iafu1V2F24oV8RiRsAAMWXU20zGkkRMLQ+STsLwfED6
7yVzcFZYJBfMg7vb0S3NX6VypdJQg4ZF5VoqV4WKMOqUiRD75RMcrMon/DyaXyNZy9WhXqVLQtP4
PlxRry1LmoVoPJ4Qq/kuMGnrkSHpoOubiqjzWtPo/6KcL410XldZutXiE2GGq2sTuj3eq+4ZsOsv
NQQAQtww3GABR3PwpqcY2ztFFCBIq+PuATRt5+hTPOxnff49R9cOEgl01lKQJZLE3ZLjyQGOSUt4
WnIMCecH+ussyNz35yoSxkBt3wSMK837T0Bp8A==
`protect end_protected

