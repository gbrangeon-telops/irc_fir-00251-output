

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
lHZAv/MVAAt3F19GG6CyO2D9ozHTHXUyHUqVqPhHJ9Up8V3v4BMtL2rZCdPHvvrLl9m3lxdPLeMd
yZjuwpNKug==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
V11pDh2GdTX922gInHRdE4PGQC5LocLJP7s9hbeXjPbTiX/dPLHGusbEN2B0toY0K8U4vuWNSniM
1aH2SNR2JV5BnhJYTc5D8l2e07TnA0V6ktY1z+NOBfbsIHPai5FO4rlYQdX0gfNxjRiE4WpTGufJ
+8B9yaPmasK5qJ0hmyc=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
0akrUk3wQb4EqzKkib7F59nSOOeoy+q3qc0fQDYykXO49Ll/FgY0ewL69TWySlFx1Cac/+BCy6vf
iumuPLpTjOS55mFm1JTMxYzM9NsagXEQHLi1lEkcr65/dw7cjFH/RPICXrv18S5beJM408VyZvsr
NCAeZ9gbVAaeGzkHq6VNPIh/P5GGGWEK3241GOn4p1v1t2GkteaDbOSjGK7wX7a4kTfRzrAH+xYH
86BcPdOp3oyEseFdQgL0BZboHxt4zJr0bXL7Ln+oOm7kGCKk4PXPdudDDSsXKQUPtDHqr2MHJwZk
LDVjKe6pX7e2DnCF/lojAxyhWqtc4aJmRRvYWw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
P2FMFi4MUNbCcmQEmOw8kkGKpCf5liEfyrVflbrNDPfCQyQhrfO1z3elwJF/eYuRk4Q8ng49IhJM
QbJUTOajY+rTGsCSJpmNj13e1oNpCtCwEA2TBzHdzEyAxDwQ0hUh3ZqnFSNQ0MMnavo9wEIKRylK
MAHL5TjDsmLJG1Zi4ZQ=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
GFuz3jjDcNus13vZfabnTsKTQz9Q9tOYpUUTv0v99miJHiWg9X4Bm37tDSsBPgge2ZWYV/fIZNhM
o9RFowO2ZPIK8CdMOp5y1r9QlxbgxiEVYj1tH56LRgvbv2A1ghGFDDY3Qvyz5G2dmEuSZ/58uAtK
A8Mm1zy2Ln16qChURWHrjkDuCcIOuGQ1GysEn2sqg3E/XWxojTbAmy+LaQrAOqIwoDTGFZ/Ek5fe
49U6fyDbugt8sjMOq32EEkOAQwWmc5uVOZWv3KIDCD6tRxPMIg8J9cwcCTEoanlasaaRs9KqN5go
7g24OWiCSjQz8Pf4KXR9USnCWt9Xh2mPsrZAPg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 20576)
`protect data_block
0QvQ7gCr5NwY8JHUWY8uFaHjiW2ODdDVup8xDtVrXfWCpjqEpaC3pv/BSq5+K8U1QXIWI4xbjrbA
45BZiD+3We0Vm+zRsTXiMxwiUjTqq/l3aXEygAbHR1OZlRP816pAu3CtDjot49Vm71SVX/KY2FoN
Xzu1gOJN406mueeAwswiHHV6aPIx3mtsbqgVWpCY1jUH2rLg+ImjRww/IoX8xPswlwNx1GJtVSdH
xlH35yeKxidI1L5v0UsTMh9UtDbRAaUYPEvvb2vOb0ZDwNDDhBLHFF+0FZ+/aYqFcZ75XdFBwsgm
60L76p8lXCuMrQKzSjVGjFg+DKKikPZhoZbMpqqEBdnkTjlOPk5chHfPWN7Ivq/zzI4jO4rL74ae
fNSV28MdJ9qzzZTPU7CO5kaGPnxy0fh4WQI1al0tIaEsK50OIjI6vCPJ9tobxyXx6qvcPkBtBTtr
6fiply6lv/EbZYL/HIdHjD1M2DrymXJsaLxXcxd9GQcItB+0c06N//NtPNF0HM/Lw4zLJp32eS//
ym8Fv9SYoMPmyOzopLBWb8JCf1FDdf0qV1SYQJ5lyNEeiDkfpP9jaV+LNChKCsKU2rDPe5h29YFU
yJc9mutbUPMXsRVBLBF2Ek7ql7JqDpT8A+UMuEcLVXqqp04GJrbMuGaf+6O3YTLcCf9l81FHJFk6
7a/pVoPEnpCQW677XOIAYxtuCiLAfJDiJ/6lFyhalggvZwcnQkC6TObVDDH9XARc/RXtRgbfiL69
4Clvf6qf/8klIFoF/wE8IQiFDqov7IvBu3sKI2QbEMang1rwDO32HDOOHpMZedClFJt0lYmOC4Fu
oQ6dhFXV87OJ3x1BGkt49Yxoj6p+dLsHBC6Mp/f/DSWnKXXF7hForWgkt4qUXjYcNPEo8Dxys/QK
z4Fj3UXGavcKTae39uVQ0U2jmU5KOrmHgEkd2ufejE8b0NF3ArE1ULaR6W05YLzPqdnY/xYSGGQW
qfFTmEQrPBXnE0X+v2ynKEHPuNhgOlxCm3CF81Y/JHy7RSU+qFsRxeXIO5Kw87EKcSH6gxYEvUKH
GvLg7bKCFGfVOj8yJOYxRUQB2w3Bzct55v0Gzz8AWU8IUC8K3A4pzmjPyHycML4V1/od55P6n5aD
hiGe3iGRXXkwle4gDKOcEx2jN0OBCapjHO9HDw86uQM+aVduYMtXrzm+vbzgnWWRdZ470FBEC1zq
zXJPvrgtDiiCdsUy3u+mNz8RHyL2ZseFyYMUTrLgdOpvjyqt3bZfNpbgjnzMZbd9zs9wMOQG0XTc
OxF3maQf8iIZWNREBedOd7Eoi0ZQYe6JwVkzwHujbxOSkJgd7Qa4vPUeJUAS833mqQevQtkqy8DD
s2IFcbneJkLoe1gyc4zhE4rOjYh739KXzdK46/6dvVu3bXHFxlYc6XGLG3QLdpRjnryVVo/QFRmR
kY1hkU2AYb/Q9B97Nw3SYzA/lD2Zzn/D65j6OUxmz+PcT/y2ChmLcjSdqAxXxP7ToIDxLhqMQK0L
Wv8rLYxh06f4Hv+Pwy7LPsopMivf0606toUQTGRk3uXzWsCvUiz2GiDvYEDayodYDc9vg2JaBH8z
QAHCoLCKY0CIWHPOpy9YChcxghdZu/Z5st9zW8U3BM0PFEIh7n12QQSJzRr6U8dqITLKRAERwtC5
VRlI6e7iQZRdiuOFHFvJptRgM8vq18gG0c9XAFo3DX/RWnI/Vipq1Rxq2/K3iNiVJp6L1IRgN61q
i2AlP2FZ8SMVflvvPTpWaNBWi3kIaeByCqRxyDmw66kYmYg22331DVaqavP3YlNGDgIW5reLjcgv
CtyvFnzWaxgfFD+eTQLwn5FG6HaRMb/EXkBpTkdpExnWZWzWvgul/2jutoNH2cLL0TGRviCUZeTq
dd+mjmuVMNFuZjV/Ingn96RKGxZxs5cYCSd1C4L8ksO8GVPTbQ09dUmA0h2kiLdqIj3eoNy7OwqA
JE3imEQXthS2T+RfrrI6dizVnAy5CrMj7HeveLSK6zOLYvQWoB2TJrVLxwrxrAgdE/p3jBz5oAme
Or/XUBkozsu24+NXpNf8tnFcT84Qby1P+Gxcska2RyNV3RrHXZXxqg+E6a497dbmNLV24vjJp9cd
jlAdeWvxsvZ+GZm7499Y57k1S3kgtOW3KESdXIkobM7URbl99adeNkb7ietGFe1hEyueNXff8Sml
HpR3IUP98taN7oqz0DzWe56njitH0oPOjL7F6HY1j8/E5lhM5qfGVcrF+z/PBt9vTw+FiD19l/1s
GH21jXJKfN96zPI1/djNA4Y2S+goD8cShW77PI6KL2vofX9kUyNrme1hHhlbjP56hmN7j4Xsb3gF
1gzS4ZZ96/4X9VIcYtx3JobJZBxQ01NbiUGhUQBaJGq4voGAMvcd/u9BvrQjZRfR32RXKx7uTvHO
uKijQcTT2j8qaXFwpghMJ6p9PBsiV5rGpjlG+wxk2KV6uaf+EZAcR/qg9KaOR0cdwmXxtT6en96l
k3GeQCn4If9T4cr1j9aLCSMYe6FE70/Syejs18HzxOWfBjvI8ahOgwB+xfFLY1aTDEF0QhHt0Uxy
DhZS6T9da8BDEyQo4Owmn+r4rVdEYty2e3OkyVEjhz3fmruw6H2CIx6DYeSqZXLPg01mGYmJ5CD5
rLGARcW6XBkddm6OU20YRyMeFFMu0zL/oj0nDMXDmExMjZIiaKufYHommmo+tWOOfh+O+QbaS4iJ
jWX0E+znxe2mBuTv4LoPN820MKRdYWIONpUe+62hM0LD2ZBShLfMpmATVCxCii5ZKuj2w71/p9Ny
Mo5iVvu7XZQ6fLQt+lUiiU1lDewlyY+rxh7wlLhc9t2dWVA3O7bd1p6jpgUwCfLlAGX661KaAJrt
l5ONdHnh5imK+5j4wkr//SaX2MkPjpIdHfzDlGNCXyKSVxaxXD6eCRqK6XEpbVIcVmKYScbReiCz
ThcJrmNQmeAR+ZyD4cai7h9sBOTEV+0tc3MMIynpcxloVh1X0hftOQNvEwKKaRAyRhP5bOiR7KQJ
sQXbmptnxWajpfRdkV8VTSUvBv4NqWColdWfCU2PKutuxTYMDPH1JNduj8KZn3rxMBTfj073PPI/
q8ecNqoDoXJJQEoX3rY9i4eMXv/FBOdpJ+jH2VEQL4wOfZITQjCass6sHW4EILXKA6ldep4H54i8
dG0Ol/mqdQoMUkiFBDFdTFFt3Gvn01CfHDdC2ZGkjiCscHCKGBPT/FAYKsK5caMu7Uhg8T7UppTK
TyxPoJytMQdMnCNz8jj3MXJeF0+3PT4lL2Gxz6ujDgPnLpiHHSqnSGprx9P4dDiTkf+ezi2V2Q+I
0qE+ahCspHCovT5GRCjAcTvTjYvYVEQ/W4bF99aMHpJABpPG9jzFN0NgisGEqeAEN5Mw2F2JxXUe
RTk3gTdv28zv8NJMfK5fSMXfaxVJcwDlHiOedNC6R2D4Hus9SDPTw/mBzYeFUjn8yMYdaTXHfHOR
/5cIvZ6vjnvohI6uTVU29LXyDlEeCd40z6p6+uSoDd50/XukD7Sgqh+Jq5TsgrJNRSkEpKCin1Ze
TMlBf4nhR1EzlX95Wa9pHTNQc4ha2mRMugKHo66j4gNE7rCCmCMqUzgQWLnyomJ5vS7Qo9Hc9I7z
SnIYpbRgDl8GLnihtJ+iuw4j4fuKMd6j7FgJ/iWjPqDGOEzsqx93bs7dYw1Oux9NMXVyDvItzcHx
otd14Lhd3TA2U0pCBGjP7CRNDPdwCzCc+KUEGSRlVb1xOgs1s/liQwFW0kyp+kMob6ckXN8wjC6Q
wpeBRNNwuh4AsijwxKOpEv5d0hlmGxhv+bm1A3ohWFP/8s8zn+udZRyl+CsToM7ccXd6Lkew6EZv
HC+cBIZfMj9WL/hAgv9i3yC4gnO/ILR/E7nH3fO0PozVzzsptuiGwFkkoUsPEqo1/PoSrVJbH75Q
gozVXve4C3BhQX3r16KKLOnr6qB5PCDvLjzN/jzE5c7Wwq9mF5tKFWy607wgOBGj/uQ6Zgh4UNSV
dw0tAzaQK2Sdq+mlOKa6k9b9qdrds+twAXHBFS8W/vwCXniWONymCGvFheWNcA/3JvRa5ozosKKl
+y9UkEJ4R5X2jebIWWstTRBXDuIxCLfUbY2QB4ruDj5TetmzovW8z6CpMM1tZJhF51rFOCtbL5RN
1LnfNumm0HyBX0vzepzXHvXzVEvznHc9ZP0HwWx0tBeLiLH6DZ27p70Z2A6NRVpKS/7h/d5YMZNN
Lzuw0PLmOJIDbT/A7tn/26ULplxGUOLK7EMNzQ5wVXSuphjmuiRjD+NRlzvf0kZfB4TD427OHPOG
dNGqCmFVjwkEJgpDkdk1ZsLPGS7kEtZK5ug/vzA7lX1fgjQgajajswZpT3hsf/IuYdha9zF091SY
+Ul77Xy/J7Du/F9YA8e5uZclKTH9gQPx36ofhF+N1gfuNeV9H3Kp8gXZywp6c2cPfk3KEQtaPV4E
e2SCyPza+wwnGV721TojAFq9kfg4pAx/RHsRaVvZeNzKMz4B7OkERkD7/FDyV4+/qTFZvGCXFT84
VoSbGEGDLTYOMUlNuvzAI8kS5AKXrkKjUQMfsoDnDNFezCIUKMosKqR2psowabURTSTTm9qVre+l
76tu1+uuQnzqVKim+sRb1w8IppmSbmY/APtZiRemA7kkf1jRUYMRcv5O69nLDW5yNW2aNTOKXW0x
/aI6aD2hkLhAsrEksPXZGl0cmhlKOBY9e98oMcRIH0jYWiqDzail8JgKfqPWuPxw3Ocw44WIooEt
4ZFyjMUNUPR2EPbSA510yBcEr6faoJrvf0fcn0Ardkr/+Kv82C3r9Gs5u/4wzwFvp67OT4VIRzoD
PC8cW3RmVqOQeB49FTNSetyNNLTZ21pHEOp4IaXaeKD5t5LyNX4EtvVSpA0VK3c50w3AfKWaEmjz
uxOl0JVtI1OulOjriIlMVWqqibkJZzk6lkoDKbNhjbyicdgbCsvoWo/ffH5OHwZJarGdRjM1D4eC
9ftSPQbhEBS12GW6QBEDuQJogNqOgnLtXwqciNYAMywyBOOH5Ra9/Dbq8iAayDVbBIF/BIf8vzjl
fU3dItl+cg/LB6c+OlVscGuI75qmptSjpVLqlp8hMpRmdGTE4oQdl17v3fUfkh+vR7OfUrvibQqZ
EgLitNBqLieYxkfmEdjm3+GVjpuHkHMvJ/0aLC6KHOIYAp5CdzAIrMw1/z1GuOkkjWOpvNwamCQ/
C4OPVBDumTSeyPajn3Q2j9D/4VshxauipKgDGs59ByEZTLw38dpyPcALhBBI4jZdP3bxgzZFyWE4
YjtF3FTwF/E/TGblKXJjn7VoEdLly2eRKrSYXaS3vNUgBsxLnbKMaccZvbWD4VtaM1sN87TRp3E3
YiAm2lxbBHkp66lHWRuVn3UWptYIUbIBB2jx9WUmCiaDDck52fu83hY9bo7kCvLoEnkTLgyCLg2X
WkFpqTBq36Q95lGDJVFl+wCrIvDKhmIoAg5ISvyqAT0azDgMyur3voXxrqlnxRKKiCB3unFnX7jV
QVqRCkGbcQWbdkjoGgPCw/pdUTgNj5wTBbBicjmo2KVdWx3Ptt5AH5xSDzY1rN6Je5sS4k+HOvOT
PDNP6srAf5ZrATLv4ZcOQ1ngLkLCVhTIfx9N6qTOqEswPu+vj/TIjboO5DcFpt1ZuqgIndHGDR2k
T+A9aCjIJca8WF40Q5kyiPYhAWjCETVdVEIikH13j/U9ahgEAcwXCvh/x2rswETRHNqGje5Tok/J
e64glEMzjWm5mi/eq8hEf6M33uxoAXJbJRbhWJh5QG5H0/H1IFamJWjp4CfxzQvR2tNjqWiM7HFN
fqKMAX8WAu7iiCjp8ntxJZ81ryptCOoJgQ390G4gkvn94J/W/8YA57Bp9UNS4aplJ/RaMg1PMEuo
ELQ1e9jTx6odlZMV3PW2NaXfrEqSmVUhzf0ePsJ0Wm/n566JRipdcbGRA82WZyzodmGJuNj5D2yo
LIdSbXg41dU06QGYvtiXN/rCLTow6HELRVVsYwUvaHkiUIU9wLKZEW2wm3H2ntNtqJRnFcBYYBUl
3gpWlPDNy9ZIKsfG58tV7t6ktj7FZ6Gm0CHFOz+uAjrr80HBsBAPWXcEJ8mfuD6xV/jEpJ6/c/VQ
HonUqMvRdBuKikBsE88PkoTVZJzTetYKe27pP93707aJGiUCFwuYTy80koOkFMkAto15gAAukw1I
nrNwkOaQ0eWaDOrIUJPxfWhH8CEUezp71mq5dh+Ou/zWTUgoB7vBm6HXbBs1vQ+BpqsXBBFwiTzd
Y983Iey0mWgRYUZJHG/fKB25BP8k1MJswC6ShOyKu8s80RXsRJ7GMvFX0Pmma+YyvkesSMy6Qrzf
PzCNc/kjTAutiRSJ41ddYsRoj3DBmQcPtbA95HO47SZifCKW9Dws7UxFy9znVOuyDtg4TTQTsZIW
N8fRZ7S01R4mH+u6uVOx7OLHhCxWfF/XgX7zu5s3+p8kPs7nkSVXVjzcxrF4HGmc+CHTxulxDzWo
y3IpqNpGSyBAMa4nSGXSSnYJU1ApVy9bVPBsSjhh9ww+cU21z9nfA/dDhiFs1BGgrasvzGOfpkjL
gtDy1m9YtyjCcgqYvv3QgTvAbjZrGj4aERuTCpgWrFKhD+OwyxTaDOjWVBtuEzVqr4nmi8gxmuop
MO/JSGOgH8Uc0YtXUKvBTT1q9U74PPUXcQFZsNFBg8gfB1y+rN/k2ZXkPvdXYh/rwu3Lys0/52eF
jT74aOpdSfx5hoeLVIgi3rQZHuD3UzVpLs+3LDELDQTOae4ru35iSeEUZEp5Rvp+ChPvKr4fX4tN
HkVNpd8O+LzbUw9kovLNIOV5ZQjvVdrpulkyZr8ZTqh/GdH7YCYd7W2Xd1s1KJ2hFpSrIAP+5PzB
VZ7Dorj7M5V2wGNyopvpH1Fi5yRoCiF6vddMQauOlGJNoY/j4BWdJt6bdynbqaE7S92Jthx1IiyW
4DqhKJubUMu3nQSETqkYJk5TRDmLLjR9+j5ZySBC8YypKzlto9FiGpTux6S4rHS5jOpuFOQK/6gP
SCRlCGIsndS3JvNFpWX9mYAnUtlWIfjc/CEE1oWbbc9NUla6daA2p19oiPIIDEB14fbNK/s3UCCn
FEN5P/ciYwbTb7e0HHtu+KEc1kL6GCiTkuE/+xiwHD/ZMhp9wswZBUxONx1A69h66W+IR5/M9lAJ
21XFC1MhN3v9I3SIW6C4r6EiR6ZI9uR2pu0pMW4ZLsuODN5fGDbkk/PJ1uhu6ZSbjj8AN6QuP/Nx
4DlWvxau+DfOLbF9pWg4fKRDtSy8KsCQZJONN7ms/jQdo74J/KYj0NOc12rZ6OopqtjkTmpCdGGS
Aetjppg6o5ZncVRwwvqMrmCj2xlVb6912Nz8osdY2/JpfSXNt+bXfCD+/wFJtTG0THvIQlPt0JrU
u7PXkOClrwjJ0s4C7xdeDbO1Xb22L5k2S9nmVQpLYbKPF88W113iulBWtQfhTXJCDo2XF11my1dW
QHIbijvVoQ4OE/S6uPSj+avi6j0F22P33sGVA7+Kovfmixbu/sCUxLibb+oXi914A3o1tHKA0NX3
AEaxH/cH1Ro6jIVvppyVN2FvH0qSrPFH+bS4K+zy0CV6Lkx3LxCXvTxgjf6I6bXSx1mtYjvzLycm
0AdbsA7WLG6/B94FlDCq2O96UKjvu11Z8XJCTcwZpjBhLP4gFzvaSD+ogZUfuftYT/Y2F7oPJmin
aFh7iQeI80cU3LRoyK/emxC1BP9iv2a3sOY2w3u9h8H7HzqXcj1YQP7VAbAc7P93r8ja429X5INl
RENcIxNH0oWLFzgRXPGho9sSK2c+4A4tBEaeA0zClPJtlm2DvHIij9IpN2skKiX5+nLwNGIOdlHF
Ll4oJo+cP5z3xAA/KOv2htktkdImdhratqNsc3rLolkVcHvk5zN3lsnzO4BouiCrE4ZPULVvI4L/
fNHW3gvb8YYHRsnDzq7V2B15myFZ0f3ICzu/PGhZ68VXCYvSy7JOxzv0d/AEmcaaiGpXGgokZmXK
042U9P/uctZ+gjinqLq+6JGx/639U2U5GsDKcHDHJo4Q+se3Z83oZOj4GrwYRRwrWvMWRV6KRw0B
bPtGU7hkb3geAp/aoc1i1heW9Z6nvg5xaFYNyD/g31d6woRZ1gX9hpGOIHP/wSM5ZWpU56yWNxHs
WpqPzLvOUv/wXTtJ5oYTv8fq3Ohtg0HkIjzjE2+CAZIPZzOHPc5nAQePzmlmFhDhv1n8+frDOZmF
fLUoNodMGk5hLcEGQ8RKwy0gw1MG8a8fK4ZvrbOQeAuRYXEiSwYy29mpYWQgV5N+Kf13SvAOEjzk
bc2VFUhMawGnLaOmw9Uhrj1aaVysQjUZVe41QMyZgnfhLVi0m9RKUXljVomcqRbL1qOwxjViTn4U
IVigXjUtj4s0UZ6FbVKMJxXlkaF/5xhPoFHaJoKKScUCIdNQihTO5ClUV6zoZzAthWYvYDBi3e8t
aYVy61FCTXeL/mWqiABdIZ/bFxWhEdc9ljQcPZovrFlz+yaAuSJ5ibUjlf3nLPEHF1S3A0KSd4jX
s/3uGzl1ohq754AtbM003OM6e8FNgiNrVmWw3kIouc7lzUg7y3XZzrGuTfq+CyhIkNFMIAeWjI0J
mX+Lena+tJs1D6oy0xZbW9TCdrcIlOid0Y3PGlhn0OYeRQ2xR0yd66zdDf77Z/SxZCuk0o5hf/kQ
/0dHNL0p20m3rO2eqs8B47hhRVWZYJGPygqHsw4aARZOp+6O4agQYn2j1LzieZihhHFDPT+ettfA
6D6hPBbsjLuV5QQQ8Bos7FJn4DiuZmSrs2nTsyvE1cp+XKTj/RqXaX/9epzOer8f/TUJqkVakDZS
lpMFPZPDy/gh3fJu/ognu9bmpPrCuYrVJe5exhsCQbzo8lRFODUofaRWHIGrcfcFyRN7iMG8NEVG
o/TzotLvxcoCjMyoaflaqI3D1+P34hk3mKZjfPJqSWgrZXZSxiRW/KoqgCqMqN7JplyorWnGH8bI
dKaPUnej3POCApJ1kuOxiAiNwC0JaEfg4B7nlfIHaiiQua1T8oA/mxCCQ+v4e+5zXFuzihdLRxCE
AJpnMT5WRn/L3EAS+mS+7uz/hoX5CuYM1fnHsvg8lmzzKPISH6P8YkGdnWDmjkfscvSOnqHAnh2G
lhCqC9oe6G50iI88TKd/ZD2IrYGz0b91sceBmjKJ1tp3UHnJidL8YhGa/qQOW3XBsdIXThBmfJq7
hF/JZoKkUUU+v+g5kVxUAW195cBglhheqH6VIGVum2qKtmofZWrKj9RO39iMoBeP2yMtPPj+oIYo
u3xk1FyAjNZY5lWHDJ9fUYoUQgQLTzXmUca+qAPJ5I5FofFZWVkhgJY7QSet4EuZV9/L5pY5r64o
2IMXyfZx8o8N+gGep4qOnMk/5+mpQoBMcbGeqSB5tvcjKAS/mbZQzXGuWr5tqpADldH5RBtbHfYB
nHQEmS/fTN2xYSFJRuaWsCRpnt9vPfr3d43sHtQ2OUCwjL2UXQJZz13Cd3534saemjIaUkik2Orz
wX+fOo0Dk/bbfVbK56IA80k3EsuKkIcbVv5Wx6BmMdWAHQ38B9NO9ZQdzRn6xca+mfj7phTVhRf8
rQgAGULVlbN9jzuwCaEGnsFq1GlRvh7N0v3BVyPEOLc4evLm5f7MHff6oDwCsAYg3ESSw0wj6BCy
npaPCe/snbJaOfl23RVR1tSpRxgN3Np74F8PgJBFm58QBIIkxTLhvTg6syJGPic5bXt/6hh+tBB+
WmoQ4NByAMn5M7rpM1xqpf8OXX5ALU5e1VYbLe9iJmNFMfSFps6QzsbozKXZSuKqS8xGdEPcJyM4
XF7h58Vbvojs0V18l+i+vnJM6yRJwD5RzFC6iks1wTD+FLWUAlSFF+g67pIfOgeW8dbtZpN5vPch
avFHpuSAGbZ9n6MzCzqx7Bmc2/wvtdIywJxzTkDceHbx+kQ6dT1MUL/YDCJIr+5I6OJusRWA0HmO
fTUpiYW4EwKaRMPqsK55Eiztx8hw4VjomDHCN1CkU/Jfq0nD/XfqvkuLwkDFkFderOMSqX3NhmG2
ijykwRJ009/8u98G9k8qW+ygqVfnXCKkR6sW+bL9PqhSSLrXOvhxQx1F/v32tPnmG0hHVesuvxYD
c1ZyZVI7447tLNB12WQ3NPx+5ybcfOiZFhmhUrKU6k5APgVfv55XT7OueDYRJa1GLLwwzgNUgT+T
QMd1gew31hlj2TEdGXn+2BNpt1mR7kloOeujSvRQgbqylyDBAekK06Z59QTCkGwZFul4V9dBf/RG
tPtpGMRDRb4jR56dQnoH7QSr9B83XkBEiVb1OndUL3+rzhHbdaBGFFztkM4jkVqPDxs7q+baFZeG
khFY9GzUWaOr9tY9fFExpSG1aj9BcWjMxS65L/GSxAPQ6PXfQpLJ/hIH9OWiz2ksJpF1quLZVcmO
CAw62AYEWtaLu2Y93KHCq18J/Ug8YY+NWY8xwVRj32V8f2L9JIuZb8BEKyLDVrAiKHcRDbw0tOs1
FzLvwlrO2TXUh4HWYbH1tYETk9dyRlBEvd1ZWmRKTXVexEYGAmiOK7TRVcE00Bavk8myRgbDqqFm
y+raOfoJF/vCdmwxX50rXI4aQEVWsGMmfiitaSGS35aQHRn51+mJ8I6GdWFGtgk2Iyqz5QElXgGb
ma8nJ8AczAr1Fi+364531fN83SrdVJ3lt+J/3jfi1GoMieLMzsA/rTVf5bihmVGCreyO+8B4UO/g
zcFZEPkfBcF2BPjLo/zAwYIqJdNUx3elw0tSC/kUxRA1jsVDj2A+vHdvFxpK5TqUq7e11hB70h4s
YB5Zmhbde046Ontg+y8tKHl2RBjyWCJ5M3EcUXsO68RaVVm8EPjyhgHH1llV3d9nqwbGbhpA59A5
f3XVoBPxcxKNJnTpIsWiqQ8KMT3w15hSaS6quLspjwAqKDxyXEKT1sQv1hPQ54ZJQ0dER0eEbir2
xDS0t7YWTyCUDRAv++zEj3oN4QjMcDv6zpePQ4J7kYnQYs9I1eyVaGFcAAmUJZiFiemrYhQbrZdY
pUBwFhvw+YqNvuyFP9g77I1Ze8eBm8SQQP8PPmrMHL/qgAEJdchFeAgZDs8XENoCAsnkTVt8Ew41
F9Uzxr19RAZhcgOMNkkOEqA3y4UqoZl/UKB3dFRogDmK4zewPSy/I9iCYpNzY0VrKmXJUgJPV2/q
C2zylPwVmjW7d5KTDQs5r7FMhPmXD7jNNbHqW7IpMcZwzuOjoVB0fEJTyRGTMiQvchSfALeMYc7z
pVw4wK0hvPqxUw3EilUmUlbsdSZrXTSxjkWu1P7/YsT30duu1WrT7CR3Z2+vdy5kkvidrN0jbsbw
LXLS2KnbPFeNXKEJ2VLi839V7AzFXhrXsgFtg7YUCvAibyqH0COJhs4d3Gi5aFDANL+6EjrENaOm
u+4VBrfa8Ql57UUDE5nIjXXaEC7PIozvXSAcEVTmWj4jYsi+RUQCVtO1B7bD2ttC3Dj3tQ9WyrE1
MS2sMyekgMf2iUVpBgi9fQVg4nUm2Y1HuqN2ALDUE2Gg0HsDPg0R+TtiBnJopApxxY7nzcK9owzn
vDTLDhIeOg14RT4T5lgPFijmBztQK4thD8Q0ybwqHAfhwZTWE1qfGBspbOyEwwvRg4yYjb3fhFmc
DDWrYVZHh/MaxcATdPva3NkVCB1S17Pu8TxlFnTaJ/9Gv75FG8UPyPP/wnX/iE5jRsSIEged/H8j
f0O/b/P+x39iVHLhmAYHtQBAasuiVXbej6vDvAY7x/zS28H9JDyw3KvLlIMQvEmf/QkWLaELnDZQ
wEYNSh8zVxS0ClRqb5C4rTLCySysAQQh1Upsn8flNlUxnEICemWS3k+BXkt6cwXKPNLBk1KUMHx7
7F9y7YoO4C/3jS76XgHHKlsVJs6+EfS4ykOT2cPQWLzLMky7Tuj+VVJKfK34YedZbG4HOep+q49G
iXkDBofEWqyJvLDTP3qpzGT4y0Vj14pvr+rIOd7K9/ULcPtJTJ0Jl+bFkdc0zi6w7zmQJT/myOgY
vXTzSPGAbMdg9n+irorxEf2u+kMrUZnrJ/b1+D02IP0X86NRec1w429ApbrNhRKPWvAwYsTGT9TL
o6lqjBiO9lXqLirquDd2Tg1EYaCS+DoH7WzT+kRTslvukskp4Gymru5D5hvV3yrTSXkMRqNQQS/I
3NH0ArqN6o2KxTCX5sakXUSQ2P5EHF+71tlOrxZVJ0T2eYdfV60HbAaLqkkbkjbH0lo1nVCpp1we
3LRmHFjQdIuSrSJ/2qaskjFskRMQY/cTpnjj28ig9ti6ZSW91YfwKD8WQYus1UoJSAb6t68ZV3C+
4mBdKssOB4ojAB7Z/F3rxw42DbEV3Xx5aUO8fKBDRQuNyOjIfvbqb5DSu7yuySJCq18Vp7H0HbSS
OQvKESfjYLHKEDulT9qVlxrruXyISgOlBjSjyoF4JOsh5o9ZSa2G95YOYTb12ouYZZYgu2cWaTqh
wbgmajrXc/O1hiVhWu4me78tp0fWh/WzyrCO95WqemNujQjr/KwB6eX581TQKWnuRZ05gJYtiJXY
pniR9o28UiFYrO8+Mg54Rxbgi8/JyvPYeGrECAsPZthrQ8JZmKPlFJS+Y/Yc7v1pmzcQgsdSoEdG
YubogO6f46LN8B+BJnIIVh/2XZeoU0F8LcACNnyklZ/M2YQlbIa3GMSo6USts6MKbYeVgWbIIVYE
5DsCeVT7EDcI25M07G81b6UjFHkllylf6bHokhb6bGJDFLJEbrm0OhVvyXEkUo4q+BzH0g/e/5yg
9sCJu3f1cKWBOXV6UKKpRQpdVW2yiTc1Jy3U3YCTU8W8RNHwi/x9PZgmy0js2K2hbLBmPiGPqs2t
Ct0eBf2fCva032FTiRLy2cLvTFmF9fPm95NmROHAsl02VefsLeJD/Lc/n/hW/8cvFYkbVkqSsnav
tSPhkO31trYB9vu0ggGd37CbODi3xDVyhmuexwO+98COvjXaSfuoRoFG0xY3VhMMF018jhsfzvWI
Zm00qY+VeEYmMSDD/UupseA2PPaMWtbjmjyhcFh6qk36pdF06O4rhQG7H9W/bUVh1IBpg1iudpND
n3JOqrO19PblFj2Bs/u0C8eeuswjkLWQ9g0RIm86mUSqZNVN5r0dLhTeptAd0WjL+YS8+h0D3GjY
yJRXa5oR7YdKs2baPJfI/llNxVj/dpuxBmdeTnhXC3YwyvuQyS1ComWygZ5Ik8EmyHa4ItJCWl3s
v3HfFTtUl+W93zhZxMepnVBdbi+nR2qpvBNaXNiSBjbu0UOfPS7wo4SEYPhWyZuqiDY2VuhBSmGG
14YAxr3nKVLWsb8q0K64iSbCF306xUCKe2XLujFiLGslxwHokf33B9E8zvKbrFvDeHt3jqg1tOKK
KzVzikBY+7YpKbl7Mn5MU50ZRuJuc5+yyiI6iitHd5NZ1LYCvMvceiEJadQIFuOvQKaQ4MG/+NSJ
O4y96dBDbMJqR7AAxqS5+Haodi597SUuYC/d0SoKWqN0Lypt0/HynJsVUliCf5UxNaJSNKVgf+j/
TmRT7rZsPpb/AtQREtPOE85MSNrgZFL/5DLkLKaz0Oira7ZePEq5Ud2sjP6HlXVmIOjCmCVvz4mu
5hV7wqWhk72XATG+zGQmUUriuthIBEIp472WxM4iN42QV66JQB18RnGKFM42DQJq2QG1Cc2/PFDf
d2P/aopsZ4G5AfsYB14FW5+J3M9gUe154TNhJYQ9cYGKN8cfaE8js2WRwDA6EUVOisEmZUCKRdzI
6yOpN+VlANTnOAnfHoIQWDWnwNoe6bqThhR3S0ycR2l46Rl4gM2p6FR43D8c45g5WcgOSTNASq+m
zzQX0fx3TKABBlbXjhzS5K5Ho0bA3T+vjNyskuRwH87ufmzmxTc4bDWZtAeHTaxHgXFLp3t2C/FD
6mtJAti5edGebzhKC11LDn+IS15H8/XwSjP+LFYkToau2ec0EdiPaO/NLad0qYc2gbIJAvQpqnrl
You+fqVp0F86UhipgWLc5zvf17BwxL2iO66dIEkY6XFKAm6EQEb6lR9Ymk3XSfhWy5bRQ8grLjN0
c6nha6zXVvMoaC7Ppj0ekvj+FrmUIx9FVkBMCZFD+154bDaCemLF2Auoek3PnXfLAEJpRO3JRETt
bGdGFBkuh9lAnuMCVDrTODraEcnXBdnWgqlQyZiJyLeT2TO2iq11yQQ8+RPm9uX/QqeMy6uMeBqW
3GwnjBkP16YNRELJ1F2ykl9bnJ8SRbhPp+3qE0+hIetvsRHYezjCVQV8b3MZKjcRVF4uORWYjdu+
FurNzShACtZyLRfNt+5dOUMupWPhLlzPV4HwofqU7lMSeFYqNne3R4IFooJAfHMg+se04hChW5nk
eCcDXefIt1adg5WI2XB9gS2jOfTttL8iqxul5qGLR1quI53U8ToknKL7RSAcQmL7r4fTYtrTeqvy
B3ZOr6a897nnHeQ9I2gdckMDCP2hSWZ0Wt98Eb3xtomazn74UfyR2zYZH3qYVGSZ8/E/n2waLq1S
meEbl7a/ZryERw90e20Cp4M2Tx3w2chKb1M72dSFAwTPZwjPhJZ7ilGIoocZNFJAIfDypmpCGk1H
gFJ6px+9Ttc9uR8mI2+bO/RYLM0AlMBj39nRSM+wLypEqWHpB9okNUWqGk9kZQ+/wq/TLdDJRdOj
oKqxXE1friJSPsgRApC4cXY0CaM3XZEZ1HwzET95vEWAqWHCR2V1ynfk6sjjQy6iDfiVg/sLuFNO
c/7fqYW6VcTJYD4hTpNn/+QHaXqxLVRgVj+1AuQBPmMa/7jQYNd2By6YAlngXXa9w5qPuCz/i+po
E0gCEmsaFMlo7eeRf9Vyzxtz0fGO186NuINp1QzvK5LDn2M3kKvz6pbl6BjWVR2XMXCpeXreGuPf
ehpsyIPjUQ1EdR/9F7Zy64xOpwLZKTNHCt/tmGG4GvIlnTTTG14/+LZdPR+xeWJHthFCP/TK7Mhj
v+K9nywcsFX12K4I1F8NuwW3QOTi3MIP3V74tC1Vkg5P6mk5g6/TWtYIWfgwzLNpXWuo8Oq9VuTW
RhYlk8uT0vScjakLgfkK9BciWaRxjmj7nvlxmgS5/Jt4RcwTOlLUOYaC+Y0rROpKAXHpx0P5QbbM
nos2L9uL2/wVU6lkXCrIEuD5XQ297IJvs9XmrBfJxMgtrBSEvjuJHgVn+MT6IvfhpVh+ToJ84zHZ
+2Th+3n52UoW/GbNK0wmujAqVz4msVwv+b6xCXNJe/fyfvXk9LqvSUT0oENrDjQ74Zko0HV5km2G
gjCGopF/UvrYegea5tRun2mozBv/1k8pZvPT5BxfI5QLAOTsqOP/LtGSP9f3RnKnpwbf6Pc+3yF9
m7CFQxAg1uWKnvIHwhwznVhb9XeyuWFP/PeE9i16cj5ZxgcRDVV2ZqHwQn8LELRoUn1cY1WOudRu
IrP+xOT2A46vvtYsb2AskNIUA4VYeqGseXgV7Ot+ahM0CiS09l7Eo5/s2jVgVFUCHivr64KF/+D5
Mm0FvEnWpnqbzAtvMmZoOlgz18WoExYKJeGOapp2ai4lIvQW+6jCO8sD8l1mEnTuLJwm+yydQ0xE
Gf+JYXERqYYPe+uXkiKNe+vRxpSK0e1MdeikSMcWnCQXEfonsi2gsnxJnSKlBzQC73xPizifJXK4
KjfI4+CrJPs88XYctBZaz5O7YFKIwImkpcFnM18RKvowQCvM4BMfYNpL6lGlokYoE16cRAN97UME
TXvBmKwPvxBhqhwjXsn5nhVP/39Jk8SNE/ZrZfTDnDBNWC+R5WTjyl7vjEmxC8gQw7WZSCzZJSvg
6wosNURc1i5qnClgSS74q9QKGwQOcroR4REHhHcg96UMIjjlYD+LhKl0qHaBcFiAITrwTPdFVlyS
vKWQ/WtHRLSJA1fhYCExVvVjPcg+cW1wRM5uqlPLYdLFaCcYO0Ziqe5IMW+HQ1aMu8GTlg2EeHnV
UvbK9LSu3W5fJsnc+azLqg7rjXDUGniKT6EMd4baTELCyW72cLzBvZodqBurIJGlh8N6pOgQbWKt
6vC9QhAdH/8TP9e7hGRMKBn3JKtV1hlOoPc9MzXl3LWLnmeoBp4072RkNqd9lnBOjVax2y9A+uQz
CSjs09kiclY+JuchuCaGVLiXEsHJA1A9IY/4bp0/DvHYfdD2hHDwb+D7L3eMGF3y2dTwE50zoXcf
cDmB1NTwZ2b6mgKPyIkdAvBDRxuFEZ8P5HLtx9/ywLq6L0V9KNtfAGQIsKc+56qouyLmVCxhX2En
Ka6deMTon9FabD/Mi7lHZFJ9pN8CQjOQ6oqbX1lYKquDAHw7pinbtTIScQwTyFXlJSUy+20JUQRb
hM0d1ErbgiQHYESXvO/JuAUjEGwYx/UUSKtCxWhJbXpxYv9vfmVazuHN8k6L9eLjy8KAYlvV4khW
5FnXLxqxKS8mz9G5D8bv7z/S+4EB46WX4Y0bMowlpWemK/pGM8RJYnmXywoPwWdcQbegICdfo+r5
yeydQBmhoZyMe7LcbbL7jAl0sUr3niaG9BiFBqQPSbp5Dq7FpU4lb3XJuHDwYZlewV9m9aB6npfP
3EREOrGpARPV88nIEf68KHbt2iNDj2+VZ3u0QQk1Q7xdbpWpd4m+XbUKUQIddxuqHZzlWiD1wjtw
c+O2/BHtgFIfWFQDSTcVJhkDpWMR0NLBVbj8rM64Do1G9aA1zVMkrtshG3skUihsJJHcNy5k22aW
w7fRcn7wGfrQNF4HCY+rR+wAzfHHbjBFWJLsU69dXL2Pe6OSPKbboLIMXBB+7ESaULzuFwMlcOeU
Gsk9INWFKrtT4jjbKHwcbvTNaGyj195wbD5DuJHcPIETHzvUWylx5fS97gnRtu58NBo0HurdfaSf
Q7Vhy9IGxwO3P8rdBvgHTOc2Ju7BuBLwqrHdUz15joTDaZuDiC7j4muzsgcWp/ZtViFKn8BKJQMF
T7yQy3MlqsVMpTpD+4pBT2qzIslaX+BGlagd9h0U9QP8BNjwZOr17sYf+KfhwDdo34IxTuFmqoHr
qjj6b8VpNhhfqmybvbz0yq1SiR1mBP+c/IVqmwHxY8Cf7bFeF2NqrVLiNR/Jr6j99Xeo4GaFJCVc
LSQwuLo6j6FHebPUB3wVUs16Itfwz9yJalYqVuJl2ECuau5qXmk2KXReoJffapXmuUUmWobO53oO
b7GelG/Cipt1F/x3kgOxpc12QQr0+taEW5ArCaDVpu+E5eapvWunafC32KdsOXy/UYziVdHjpSbo
vh0RLuQMt1aw9eD7yoJ1k938B1LlwoEXsPSb3IOT1HLD3G2I18iUj8erqF55ciCATaT90/lMPQ6g
VB4YIkE7oj40/wr23f+OmuGrVOgDMDXzouCtOChMEwUuV2nLN3lM0k4u6jhu/ULNQzendBQXczls
5WVsvlPPXqoAmotSUAxdqOBAWlXGK1vvgIIAJ5eiOyx07ohWqwrscNqGKWln7ETj+vLx98HqwgcO
MhX+M1Jb/hHuVoGbtQ+UvlFx6ZJpUyHTFUiEXe712Ei3fQh8scpDvae/fv8Z5OoYubRCVtWSSNNM
coHzcLXH3KiuuoJznKxuprRIMu7mfXq0Ul2D8m0Y54wLydYQbl++Fe6PzPeRyKHnF0c2jAkrwwFL
92OcAHdVIOwLG/fRS0fKrbLOXriCZjoaBCZ8jMyvuH/lfS87J9rC3QAG+21fgad2ADx+uEyFXZMn
4DqATbAPw3kQtqV3tEvzjvJK84xBGQq8jkEfeVXovRjfB21li5oR8aRb3QGJtEEGvti26UVaO6uz
7ERo+RLFJ907tddop+EZ/zFDMH17h5tpdcwX8owfs9A81QvW2cwb63mIa4cfmxNE7KF4ePztpXP6
JpmOezSglbEfUc/S2nuQGEx0bEF45s5oLZUcDESWwcLeSDvBGpFPdPW8Jr+1KLsFUMYK13kV6L/h
7HMKKAIlItdeVDVRYFpUQwivLFismzd9hAJtNaN2CK+B6pmZd3kQ73fL+Dt62cYajvw13LCB55aX
6NaXMGBoi0yOzqySy6NVBrJekwfe3HZy1znOfa6t5/wtjAoiUAhF2hhnzDiuX0cPXCLp2zikR1Um
T/YdYfzuAPKXprr8DTlY40sElwfS5M5L/OQy00ErtPBngLuFfVesxBW57/KY1vP5nrlxFGSyRz9A
g5FPzt8QFcvBsVrUiHLe0/havCz2kGySiY6i2ZQ4Y1a/MOJyPw723zW+xFzasWPm6tpMyu0lZm01
v3LkWwNvnB885I9EJ8QroLv+cfGsHe1nq9rWVc02qbRUN4Dnuz7cU+ic0Hw9UgTA5SGa8jYbKlJH
RA+BX7RbZdyTFL0bK1tVJc5IZMozdUQF/emInZVrlcjsL8XzXAFJfvC0hPM9rU8wVk0irR7an7Xv
raPu6LXI3KHV9IrRGt3eRpKNG8p8KhzvymF3FZpYYer4OSHnJMrNmbQdzCw7EMnouARlB7Zv+2Qd
7GIpkxfldGEQ1SsmJL3WL2dS+N0uInwSrsEEH7Oa9OIUKOjsCao4kpRv7e+M05yV26DE4sY2qMjt
mgMbEzZFVN7bwn+sdmFgWH2h1WM3s0j63wmmoxBdf2D+3ue3ppDgyqowDLaDOz9d3Pxe/WvZ+z/R
f7yOe60KhrSQlGhZu0SttEPFKr+OPOGdZdg9BaArCqIvbRWHkcdO92PAg1hiZs64vpZIJ2mIYq7q
idz6rowbxh9HQBjsYEbT4VCnds8eCggVWmyePbEDDi85wSdvuSEaVOnphBdWxGMA6NomfjhWwYkk
Zpe4+4jkivHavs/5v8PvxucWpoqfiaLbRvS4j+3Vz76IJvg+EfG79SXdXRYyLdhdHYS97nObFBWI
lmnt6WQNfFum7/McfCxSBeAfKuttMcN3H+O7eS0tf7nrY9jEU5pMLI5ulFY8LSLnDP8rC3DD8vfG
2kl2rrw6iq3cHw5Z6Vfr6TMrEh0RoW6EbnYAY246YxJjzgS7k1BDNUV5edbr4uK7RrTayBcjbaHO
2xQtpRDVtFIDWwcYng31lmfxsyOY9LBCIrbMCl5PbsF7FCbN8v41qaK4MUAI3OvYj/a8vnz095xw
LLFh9oEP4DPoSq6hm0PqlcCl3punWiz3aRL84VC9xyTQs8BCEg1Xsd5KF82OMiYh4MHXHuCXVJRo
jPjCeVaWDTQzRzYUDp7x7MyvQLFSjNPZXG5hMk+A0MY2yI+4rrrR8eWX4XTMLu8x1BHvsG/JCtqm
Ffdps1q4mcA0NZh/bdfzxQ+nbzrfYPpHrL26qRUzvfw0g1GZPmMITELeTL5F31A+DvSoNAmeFUGR
qEGytMF1XtDNnWmAMhGDJIGw9Co1ISZlvH4TyOWjZ2uw7bK4i//plBR1SsjMG+HFT0V9MVYzP8WX
6B8+9WSJSXlA3JkjnTRM7ClHRHp/NNdiigU/1l9dhLZFL6Qz+LXL3eUI2RX+KNpe9zDoURaDASm4
z+sWQCQFYtdznWHkvR5KFXbjeT+Qltm5SMrNcaVTh20hlXsVw63jeKfWjtgzLfMD2eEafQSHhUZ7
HJ9bYgdFInJpJBL6t9ijcumZ8VYlqS/DQpWgH5pDSO+8UrOXQjtP4dtgkkZ34jTf8vMFmBQ0AGBX
p59Bj5Pofnmzn2d1LThvxlwV4tO+vLsYA+Q2uJUqSvp3/aaXQ5zBeJP74XWDict8W7KXXmVw9754
RPMqh1dl7bi52FrUS3R7qPX/SCDqqIgQtAEI63zKEiwJzNOLMo3IcUBogs/MUb5+XbeI7LM53htV
93VdTExNfss91osGQIpOfErdTbgvcWZ30uHKrr4k/mY9ppsYxM9KYTy14C4vwLq4nUl+O37bneVX
VVuiS4xNRFkMSt8JyV7pnW0Qp2WMRS/Fp3v6jfVTqyFj/YXNfBR03CWVflhCM/Pea3PSl9rnne//
NOgCkek7UDzGrh6JkrdM1GbORtBmY3MFWYgd52/SC7s0Ohb0IeM7iWhOyef7wSFvu1EpgiV+cb/q
xZwsVOJijV/G5NWSYILMDoINtLuq5vaBQTQ9oZuueXCTfPkMAF1dcR/YcxuMKjKxKZmKouONY6Co
JZiBk+PL3yR7YMKw0n9y7hS/qBJclfUKIL+fPUx3ZN+O/uxAtz5nPpALXZY5dEnUkHTXEbc3qKUp
DMBelxec7Y32tX6AYPDkaZw+MOCEr0IlcCLkmyzTSh+Pn8dqwonZrvEzf2nEWzzFkKY1mxe1xWJH
GDOd18zXzdgc2w2pQVbroBJRf58RjbO1AeGw3plil+BOI6yIOaeCEK4yNfoljryEp7bZU34pUTIq
hYYdVkQI9bqWaLQAUIhwe5cYZ0GbXt9y3EnFYP+uabd5gvRfxCYD76ezy+RUXEkfdZ/HOwx2XIxJ
iuHp0lUBwcmWBHCKPD/QI6fqWuHpC63rHTSmIJoDZ7291J5MiqRiTp44M4dksx8I7YBXNbZzBT4z
v8kxvZI+dX7PP0JrY8L4+TrdGVwjVVz4Mg5OGkERPzfPMREn3CCEQNy18+npopOhOJDRs7LqSwSD
/lXSin5zQ91a6DHbMNhqpCk5I4i4ayZqgE1JLcQlLb5B3moDMTx0zl4AviUGbK2lY4Fo7sqRd7Vi
UPemBIT3PDSxxM1Edp789tq7sdkvfBC3QGYX6L7Hj1wl/2bR1Pn9lxQS4zYP17VNgv9ytygzRNlu
AHhQ+pByujHkk+FaXPpcx+rBGRNGlVf++Q6LYDbbcfMfu0S5n+NcGiiWXr/OsEXbAZTtWmrDz/RW
LyvgC4cq6DyBiWObMZSBU8114akyRf0LkklHpvYixSRUDpyYXf6oNAqHv+8cTubZCy1/MHeBQp3/
ZJNRFKMndkYWEra92PoH0s1YpcrVP2yzRrgU2UR47kwWLKj/Hobv0kJZrN5JixCdj3gCSj8xKdN7
Bzp0vTNgBHQLyrI1lIi7AKJAMGpw7QvhVWQ+TpSMOOrfi2ziwsqHN6K2c+VlmhuQr85yBZvodRlu
OUjJPbZRgGl5b0tDR6Qm6dKLYZiP/OhGimJl+nA8PQ6agVsx569+DVgn9913r0axxwcI8ipn8Un+
c+yNHL92r2NMjJb8EUxQEPpwxnMC51VSBgqeV1g9E27ejUhWxIv+1nq8asFiLphH52ARB/VzDLZH
L4TR4Juxs8dfa70MMxhFAjS5AkXeG1bGsv69YAnXbC7IffKY9ZUg6GHslw7Ji6uvi9o9AwKrioL8
0khPCUhGipdH5B88X1AcnhjWzE20uSaO/Y7J74ul9BgFfKxy7j2dYw6I0VULh2qECf1ACN/CMhQ1
ueoahGV/nFRuL6bXlu6WjC36m91SDFLsCFFXyK+ehVBDhOiVOOfhXg3EFt/yEyWMtHquH8n//7rb
5kMQnG/zc0VNyhq7gh1ATEnwlTg/SMKRGLWmWRK8eLJu2K6lImvEIBVOQQdHhZLchcih6HrUdkhv
AFTnAhyE6vTbyLztkAnsrGJbMn9NohobnA+B1xOtZtyGc3kLz8CZPcjdnE3oKn4DP86ZhmLa+179
c5NV5cwN4DxQ/SUa2uPWkSQ3JCRVPmgizc/9C0SkOBgSpiwEe+GantOroAesbHTzvzX9ulPDZjyN
60uKIVPzAumCP1RkbXcEYSKaYf3VSfFIfh0iiGASQ5NM1MF/ub+8D/mxS4YKUw02i5Ho4MCa7Mua
mRbzYHcQM7iSXrlVaeh8f4OxDlUZRaOJeVYgQ9VsG4zYr3sqUAqeRb0Zt1F4vpLAWPcLY9sg/ivD
NtnapZ4aktpAe11bW20CRpcpxH4ZtbAsuHE7lGHWpSYpo0F5wlmZuiuriSk2eNNLk4yNJs9Hp++a
CWMlxbg+uj6g7/mXZqhBFYRz9eG6G5l9Tq6Fe2MKnrBfveFj+DX8gPgI0hVV+U3UR7kQX+mJnp+K
UhO0S6xbpp64Nz8/cs8S1+Zvs4BHceMfoMNf+boo0xbS1baBITwCxrT/MAk1sKb8zmqfEfknDQK9
gJqFImaqrkyvxVLVlfkUFyh6nJK5IAGH3zm9IS8Rpt5TYhR+pNEblHnhpoHUdQ08K48ejmxYjhKm
O8dgfrZOt5gXXB6fuMvgtAlO6+y068mN+3KI8O82SrVD9BZ38dkcMl7bf1tN/XotU8wxH68wBucK
ZooKXiY1yyNZMmg0bIoVVZKlKXHPNG7dXHk1m5qNeMzcFSawWw1yFyyDn/Lve8q145xkalCwx3X5
tnnaXBIlTaFEz35N1yEkXs8UU+IU79CKx8ag1ywJkRZfQXwIAF1vui1+daDVp/AsZU//SFbcDHdj
h/POppHqgEDoPgI6LCBfG1pdwFu7H6nEE6WLO+unCs0WnWGPFEtgzjSXcEsHUz+5TsmQ+eH/rYFR
qkTrRm0Zxqmu2JQFSLnVRFwjicoe4RUkq8lIV+pLFxA5SUdL5j6QthQIKFnS0oc/5WuWSgVbeyXz
l9JToimAPn7x1cO5uMe5ZMQj5kF05yj+wNui6Mzi7MhQ8DV8wkI1vmTxzKa2E4h/Jc/qs1xrkgeB
a7XuexLLjMvjiAGHRIojVenzzp3sG3vGHB5Lgy4zG9MgCG09f28biFdgUCPzBmdHMStVmjUbZ7VT
QTdwFEo57qAJ5yUvxqFeSTif2zj+PUzRbr1x1Xdhfp50ZgOw0oE1MU7by8uzh8wtDz8kBKLyBfBQ
lC9M2ePAzW2Du6bi7Fo4+4wy4ni8tgM4IV2zVO0hny3vbKB1puClhkenMyV7vgJZ5oCuPg5LSIWR
QApofMnUWXWGLfbuimtnLYmG5OQzvaMMM65egAlXcJzxB1MkRY9ObVm+9FJ7/KxJ5jUba1V3GFoc
TxsBR1HekBhNWZVAb+uOtay+FaO8+8VTPXXkNN8S/aVwr41ZooTaEZpdQ3b1hBKxWCmg4ekyKln9
R3w2hEpaPY4ygimVx1M0vi6R4zh0qOH34aVHBZ+gTyMOzaKGrMdECs1ROOI58zXc3KuSSbpExcXq
FB11HGtq/BNhSk82Qowt5frJKpr/n40Xuzo5SXoI2ZlIOmWdvW3mP1NODMFdgqmn+eeyxU7an6PT
1Tj/Se5S1sRKQOqH/NxdPk9Bbba9RcxCRLWXmYwNn1+ZdT7Ug6qJPrTE8EufVReIZIsNUl8wh079
mSx1uZeXmPWLLv6rpV64Oj2co+qLX+iCNXN8DUIELpg54zfr0K60p6XbMD1yvEn9MYYoLMp+VJw7
ZQh9EJpBCYQdT6pCVh+qnYTHOYMK57hT8eLXgReZ9M+OJwK8bEAnxPUsMEAgcvcBkKq02Ex3Ii7s
Xba6wyuI3GjBeI36JnNuUd0XOzHg4jewNvhCcIqgbo9yFDIfQUU9N+2bjieMemr2s/tK06oAy6RI
UWi+8KQCfbSpqjU0z3nZgtJF+1w0geL3sjKx75TM3k+jQDYYGx7K4b8z9r43bUotXdzA3B2pNvGQ
BM4XK2LqNm32wZUwFbkP45kC2bO6KMfy3FFIsaZ/C5SFAB2PN4PtYmtsihZ/lpqeL0kogNsOO1iY
sFvl5+ENTO9WL9nYJ/UhBEBz77m+xx4UNXicLEjb+9MGLlkVnM03rMMOw82bl3WZvgwsMvKYZFkz
Ajd6/3sgHhLqXiTsp7YXU0jVTfu8Ut8iXqVU5uGJwlSaQcQMHahoUrdO6yw+uI2fsWtpqSUwvIzY
reM6RAmih5Tq6VSsVsZCoATNfw/WgaeiKtsjeyONwpCkEZkTFuobuQHxJj4cLm6zeJPVSxok3PHQ
vSXvwg/XwWf3JKkD08ocs3bw+ymGoXvUA9jX5zUGWHk9IOIoKW+GSZ3jiYWRr5F2mB4SgvdOEE20
y2UG2qomUSd2BqMlsUW/a7Ub3YJOBY182yrf4KCrYrnoGSXdYelQ0f5/T7lLYrp2+S/2DWaJLkP5
kwO01n01QVQ6ACG1DCpo60GUsAFjmE8D+cFSbEIWXPh2vWT+hpPfk1h0y56m/L5EOFA4Gll18iZm
Q5Vy8qDw1rxAA9/UPgPrtkjpJpzR50HvBei5ZTmKLwnb66kpzX4R0e5VKJIodBizlzgfJEBuAZZV
ISD+mD3tac4W46UU3VcpnIH8vXIMv3nCMbhD9t/0JqlqabfOscNfgn8yTaJYzQNnJJQDyQDlODrG
4hH4CseE+ADSpQ0+SHDU+jPRkW+oQ0WNAdCsWWrC2aV0FxlwQhfD7wazxjzbyj3CIf1pfSwUTflA
uQRd/1dI20W5EHJGDdxEw6JGiKKCgv9MWDjtk1V10JLE0Lx+Jyt20HGUUs3qpVp/WAbpwrPvahKi
c+5eQRd8RLcZG+omchzFy+AGOTJj5d2CThKczgS6Z4lLnLVnJmgki8NJXQSgAmDpnPhXJflY/6aZ
O25xz4DpNomlTuJrEGAq3CpfQgW3zWq6Y7xdWuHRMDAONPk9YDrUGGJznr4RFxrs3pnxJlEZXIOB
iPAi7dXk+/yBnEd5+W94CjOqnhlk8wPjMu+zJb3TUiPVcBTV2zmxTy3EK4MWBlP+iayP00iTUmg5
Pxeitmig+y827dGKLrDjQ83TQpyoOJwQAImggBMMdOG5S5edEhyAf9ERgVF59qp9DGMAV1bRcLmM
iz3M4mUcPQCciOFphjq89S63PqDMtqij3OjAFd82tQ10ujLxXrAZRdqh8XayF2kiOzWBXavscBqI
i/1ccPrHq3TymbFRI3vjQvwNGLZsUQ5o6OVtusrcJMi01QKDn7jfj0Z9XmAK/bfHg7ArAVONnGKh
ex8FTyITxcn7HRc3rRCnvx8n08664mz5ZyjhQkx3Zm+NGXneJpiNT+U7JJ+OM2vLc3B+7IzJ4rQk
YZ30jTj2SzxZjhAVbfMVLABm4yUF6jRMuh2AKroeEHb2+qeQJpVVVQ2hMXY/tiJgUjp9DAO7uiEz
7D3Y/TxEu+bYPkYoORiHJDaxXwi0Se6eS58v1bUYgBazKSmuDuDvjc/e7K3j5yrMH8uR6c/paZyB
NdtIeDkQ5ge8JoDU1h/dSEiLUdYi+5AAeGvwbVXB+k8T5HyOIZbBVn9Ft7r3kU7FCFDFArpg8K0n
caslcV1iV+1yNkXMITCfOzix87DM4D9WZ5Y+HHU1j/xsxX2mxNn8Xn5XxTRa451quwSndAbXfu1q
MTTprzr9+hK2dhYz6gjqoZ4GZY7hdjig7ifMLOOEDArmvXDCnUD3T4srzj2/JwQ1sA+W1Jf29RBF
krLE/qLB5gExBkfZeNPGCesw/In+BUShretFreFhu7SrpsAE34YwmfvEqlrZtmMmdmSPXSBTgK10
cTQ3IV/I4BEUPsplujOUfepMxWQ4nJDVfr3m5wTnP/ssOvsZIePfUTohv9iTNbwYwVTrEZVUP1fP
B6/GpwT82gLTGI23Ic00dumj1lZWk9fMeEqOos3bJbfP6C7v9MUMsOq9XPoDeOXUPQ6XPm2HHa14
wDfynhs+dGOMkNiK2kANmMawdnsZqq8D10Y6nU9DagX1nHXgcr4TWbjKKDPeRcfg6Hdsx6qhfyfL
fiGyMtjbl02UsGJBYgALvT+SEMD1p+MeHox5oGL020IdoOD/gzIzIks6/ke5siLr7LyWA5nqifPd
UHnHRu2OoSv2BNTKMjfZ+FyqW6Ujbia0Bp3kUrlcL5U0d+hTK4JriA3sSNW8ilTDLVi9UlpiOowl
k/MerTCXIn3uFK75dnz2S0cB/xCtfNIn34erWoIa+z5NzVESWfdstGck7hGTu7rBCqU3YC8JqESV
DRAbSLjsZCNOr8FSN9VN8XunVf070L32wHZP5TbAqgVoqwlpyhT8VC7uw9Ed+JYTjiAOGb0z8o0i
mrw7u8g9jhdw7QEhUYgcPA1tTWSbC51pbIxAEmS5XfNatTgueamWzpcCF5MwHXPCHCJZWM0LZWxm
NSIi3O34ZPkAJFVxHU+iesyK+dYJRISgQBmP7OPxPjoa/+YYOvWYfeksecm/8Ljj5KqM09T88pmD
QIaBQR301yn9xW4fqORyTQzklm9hC5MVDVtC/mQN7+psPQlkeOpxRRZPZPNG7pQWrdLfCSA8AmMZ
Yo1WvlGJBgn1PHYxl3MtNC7Q+eZWaanWntkfOkfv54c6fTHEDmD1FVifrZhBf+llgX+zoOEeY58F
Hhz/NtMaWO2i1KFFj3aCoPSJGuyJP8VqEdtoWzeDNDeY5J3T9Rzicz1fnWFubuxN2pSh07C/36sa
QMgeLiRKhFf8IDw8SkvMDOFQBB/nzd82P8lo8ItCbTK3wUaHPpXr54i1O5lQnH1rK5OKl8tU7oou
cF0b7RBo1rdm0aDJ1VIqCp0rGNlDm0A/+lHFZn5Rs5tnFQJ+lcGwViib+Dv7GPXaBl5mdzRRt8dj
YFfUJ8Ngo5FycdWt9b/SX+Vktpe1tc65U3bkCxU/ekAZ8tt0WCUfiTB5S7NsRj8aGwCQwRhF9X/t
s5XEBf7I/icsgoshoEZVzE/wJKdiYyLLj6LrD2zo2cfnV6JfzWegz9AI9DN2j6vWuKREstVwF6sX
HyFdh6wRQ/wjl/weG6jwoGMkzQsws5TzGovd0cg5pVdgsbkSwSt6X5yp4V2pMTdFgFRDnqVRedXX
tVAZwNMUFaLaJF5QdZBauiM1nkJXCTCGUSyGnbP/X1iY0k5wOUc+nGwygXCbYRtI/kAHygW6YGFn
9BVkvAdEpL9x8iNW+lNvJGAPMQ487yd3OkWi+lIS3rqCGTW5Nq5IUpVcdLIdb2mmyj+I0ahbMvZG
AldK87LFZ9PC2cjKKMykPYNjVhGu76NMDjg6gqvfFVWXDK27Kko+uuVEZ2o2gLtXSjdPRLvqJZoU
HLDpYhzpC1vJ03lufcdjpVMJZ5ePmGUVIUG1izWmF66oMHClH+wVA2oF8aWwn8PFxoyZS5yxGpCp
g/h1Ugr/0OO9pZ5uTaCKiBi+hO2m0lm+eKh1j14G7AwJeOD8snzQ6QGWYM9lNPSjoy71ego8jre8
w/7XutzXy4yosOvn6HifaFDz3Cv9B6i5iSym6Ah+EQxWKFD6VInYc84My/oAiH00eFDwak15f5Ur
KYfe6suXGWDJdExrearsFtskj6QwyrVS+vbB0NslPYeRiiw1mekw/PZjLj/S5RrZQ2EDSfYj6l4T
vM3AKsSAPqkreURYoE9XcwbdgHTH0DMiwEfEVJPJ1siWVd6IMV9V4uGmZx953vtgUnIuSY6b2xdH
ls13mfbEVm6GulKuysrwUjs10wGBHAONv7TxQXaGoUVDNteruXNOmuHhmc9pVrT1CWDc2HmK/uhz
I9zZlLhnlZJSb7AQGqM1j7v/b0ot1/4OKquM5cWdwf3wzR7eHUuuan1fmv+FsfjZMPm9WihnPel4
xQvAY2CmZjucgxmWBG81iXZby/r5jKQUmoVpGQ92boBg+cMAcguOxA9ucSrbEjhIaTiqjexl18Q=
`protect end_protected

