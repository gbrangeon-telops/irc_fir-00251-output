

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
SQUyeNX8cyskpzvvW2T3ssUGj6xZX5vHX5fJU9Ms0M+rWpNjMO6za6Zgr1K2FMwHi+buwP0Gw29j
IKEYpdzZOw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
hoBaDPgZL0nmY18FE8yzpnxIEfx7SKisNM4FVo3Ao91EGtVywU0Wb7yA1enrW6Xd+oLWYcrMdoDX
JTxy8JdlM3o+jyjU7UKGIkB+vX642Q6fBAuo3SZKPKM/RE7lQknQIOi2Y5V60nbw/AM6mvYDKdTS
wiPRLcQIZpvU4dn9GkQ=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
o9OFQKQt0GaB68TjFqZyGwbFj1TRgCs2FzlOtaWTgxoDRMFT9IEssmRwHo9pwJ5Tn3OigUlzbBbd
XTy7vthduMEKESguEgGeFDAlZPJdvm6/cpwtG3omF99Y9vBxA2K/3YI0+jDh2eyUvsHMcDbQ/C2p
zFKW1hcipARgm3A9Ys4mkgzXMVKYnvnQiSsmezjrXPsPy8jbFYPXFd6vFSGi/ZwrKMMLLNZt/Boe
k/Pl01HBEt/KNoY9VFx6N+e2ufES+vAz0H+DJSGPch6YdjmhkZUj2llujVX2dT6EzXeB2X9+1Sar
qYaNJFQdqXN7nDqoQMCiwqUZBJaHNrPJdzAMcw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
gMFEdGC+ckR/NJmX/aszkYoB651qUCnYvXxq63Zrpc98jREIyboMJaogrhiyZ1kntx31alD51ug4
ZAed1vud+wZB4IN9oJ1STjbhb+Zj5u4I029j7Gy2lllPl+1O8Em+DnBFlaNak9VTW5oxld5AFJs/
EstFEKIMT8MSbegVIEQ=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
I2MWBDnGcReW7SMjRXdvt63Rjoo/gu+NQcstRp+eRPxV1cdY3BaChhCXefqNXs4HwrSwjy6eXoRH
K9pkdKW/MmeSQuCCGBXm3SZnri7VuXOoNwZoR7yYcuzRHYCe4OVzWrXYc7CJVdShI1TzYNVzTc69
N+748OjVGLm080Ri6+7tnRVNASpwPZfo8iBz5hClukZRieQCUQgdHIAZx2RjUyVQaoW7cJ/urtOZ
zr2GA2iDsweYcuo/xtEmVehzY9Jjyk+XsH/W+/8SFJEIN/wAiWoW84/gDLItkUU21xaixyhQCl/Y
sHoICo/iHc8aTOV1SPHo9yWYmV0UZ8KJqveuUA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 6304)
`protect data_block
ht8jBCSPufCe9GPP1t7HMN7rB8UYrgM5seylw1j0cYzoyuv+5EkAM4D0DyjM4tRIy/0c72OjyYVX
FkA07Y5lUlcRCoIIGDeRWGgHkPtlPgW28J+BsT5Q53j2jMIVqoAsSQp3EOfxhxAWgh0JHGmbqZk6
/bV/+/ML3NHmTUtwGzviZNva1UIq29DVepnuPJfk5Qnm8I957pjfK/j/OOr8WIQ7+KB4DeZivfe5
6W8xg2V45ApSIt+wbRyzZd8hDTCuInO00liMQK+JJhaRFMKYNgqmrUJZV8N2o5wil40YgWQWdwOh
s1Sx+nwJDmxITaD7N0+5xZ1dAPXlLQ1EoABbfC8u9FPCZDnpzbsAnncLJD/0xAfgX1VD5tubjgE2
k6r4Vm8xwHMeUDrEjgPFyOVBR9SWQb1SbMYy10vCnhf05loi+boBwQ38SQ0eSV8YzCG4m/0tM2YS
wu1beju5uwkmFqoUPnf0kvimYsyG9N8u2utakwXPI88pBRVOWKo6LZ+FbKfPIvQtHwOJhwvoMzF6
Dc1LUk2cp9AuoIDNdIphL8BygXDuMzWdEridmypprx8MVMysx3MnCfuhGo8mx8y2aq9QlW3QH1L/
hCXZq4HRnLFAXsen98UazMAtm13j92GYmkD5L9/WuRHZmc3rLQ1CBfQ51DdUAcTfBDx39ZXB7M8h
uZnxiN16MUy/EIFReZqcqIuiR7sjMaKMXGky7y2M/GOn5kO+yMm8sOnQpTF4pCpOpdEi2HGv9Goi
X5gPT/7GL5AVo9Vjv0mxEsx/CckrVT6nTKPRrq9alM2dW9NmDtE7/NbYs6H7+h31aUIrP6GBl9is
kUlzBlrze4KZeGJC2GAwRDAXPFyCUPqvCBIPQfabx2Jjeqjpx0VftoQkMoVsG485OLF6PQqmcUGn
75cSOf83f8rcb0HtmwAc9OwYRSfy4NoCAw37U4dPKOYPywtH6oAAYVN8eC6UGCSCR/nX0mUvtQmC
QJUjECTsp+jO0v0hGt9CLI7aBRhztIQAJ71AacQAjbzf+dl8RZevZSWsyrsea8jcIn1hjWWwwnIz
ZOk7mJivg5SCThhWgSeg9PEFMQqwgAZVr4xHhm2+BcuCWaqYaPkUq3hzwUeQwGIXgfcEg0YbWuE9
O1DOPINceww0gzJ8zztxNjcndZYHvCs0R3eoRY75ty8Cez5WSLl4g7wrFccOJF+OIStmZ+47iXMJ
eZgQOw5QLVoEXTOx0VwRYYw9NT3RBrNclIiqme4kw3/OMBqpdPv3Cf/Ab8lpHIlcSHmfHh8Bb7ki
EkL0PWsyRdgAJ91vaHx8fMS8wlxyqTMVyF6eFAzmKFvcg9jZssbyo9HunUuPWyvjOBsu08R7H4Ki
u3ymgNySNmKprbEYJO4NIjBrxFN29tWjXSUeBkxGYICZS2akP9PaZ1Gff1m7yqDg5AxMdWB6qEX5
+mlpLRQdvA2cWxpUvvg/KeTO97yIjCr6wNLnD0U8YtVNkh5l7Tdhb9kSImFwWYgDryq1zKXhMU8L
kqNeH9IVswxCFVaz+A7jXcuWTveAv5G+e71rypcgdRDC8j9WGvUXSAZVS7mMgx0qVcBXXgQnPG7O
MoZknSMhpvYA+lvOv1oaSRP9aA3JynS4n7iQd5M2f2Hwpx8f2foVGwFnpI3uUvUDv2HcaSLfrh/E
ONz8xOq1/GKzTC/2gbRn7K6kUlqygr5hAx0z9vVZT/JkECnMWTE5UIuTGFANsHIANmutOZYCyP+k
km+0zmtY9SRLYDuo/bLbj6cduagAJtoY49FsFDCWbi6dOlC9WPVR+cy+MC90wjLwjZwGOqrV6zOY
afHZ9WMSwaCYQUZ0hWaB7vPkgeHkts7n5DVtf0nyx+CpAZEfLzM5PyOYvAI0XY6EGUH/iQi+2Suj
mjDEmiLSK7pRVXxWQnuAWdpvYv+QOg3t8dUShfIZZ3sSI5GhuD8SWGjSFnfrSy8ZnisyzfZY0l8l
hf89HLniD+EOf/+5wvw9U72xtQjPze6AQP6XN/bMIC7TCT1AXA3IcJVG7E/pP/tk68103bJ7jFSh
Dsuih0HzGUliLJyIFQl4XFrV/hNf0yGByOXz/1Q6jwwynDwLbtG6TV1SlLAoBGM0ihznKmXSfZV2
O60EOlHiN4snHQHKtDXCgpaP7mpq9Sf3V25h24lU7yz6vb2tCLldKNhGM40qtZX0tmcG+Sgopi2Q
k4ZB53DyImY7dvdXv8ou6h4VBryxyUPswTqxuhtyO9e+TskkxvDkSwPU9q+7HERDrsUgjNiVKpVp
g/vYOz1vy02GRQWq2iF1ZQiM2EFmkJXFNRqwsPA0WrlwS83/53FatieXS9dmXHqnAzm6Eew8GxsC
IzpLfp5bIwG+A/1LoWNdfn+LW8A1U3kCXmxzoghcLfAvyxbrmX+YBERMBs9IsmYqKrKdDxSraiIQ
YKo17jscVt7ZFh6vFTWM+W3vmWR7EvvU+G5taW/d2ZkCag6UAtGXclsRCJ+SQPH+r7kTwmSaQhFI
bUj2xAHQjL6IBlLqteOgjGElthi0COT6p4JpWUGEiRrn9GiCPnrlr/GhzIB2eYkiN4V+bELIAtK6
YtFipCTQdwh03zHXVX83t9T2umKtulkA5K2f/6ZDB2K8eSSLCD0z8nqvYf3XyUq4mP3t/afjcT8U
yIP5k4hbVqMqDx1DZl8Bnto+NRUB0dc4E6OdNDg+PbLhFeffX4QjTGRtwrX4ZBoB+QLB4mJLXf8J
kIQJkGEnLwVbIWkI5wvGfxtQ/yMu1RD5YBlY2R3L59RvqCDatIL9ZbOJQEk8vEKiNjT2VWgaPPN6
coeALSsgntqpdXMceLt2qxRNsNI/UKqHiAJBOqdNeKYyCFZqKH5fvU0g9LBGdldTjdP65/cGmndG
T1mVvTwXh6GIVdmLcaeyGuPRxuVAFYyBQelisCkpKqyQt1I9Xft75Xx9kftzQ8UHHuOuJvqeln6E
pCvuzdH29VchHirsNdLwidO0YQQoL9BkwBu2Q7lgkA9aFMRxqPiHyf8F2d7BHklYj/ufYonCNfh2
O6s6rwdqCfke5Y0JqvmJednChcR4KvnpU4/NIUM1ggn5bMNLQqDk4F6ahtdRdEDCohAIJ/j/vS9R
PnTlogW6MRZzaagEggqdS39GTzU6NrXUM3slYEJe16GiPOXGsGjdr9A9aO0ozVnj7MAB1iNihV/q
pBUyvvdRISvaT5z4eZA9wh3+5eKmC/X3RCmzeL9RfEXRoDYuKE6j7OUfgm37FTB9nkY33kOCLUk/
8VXRPBkMFn9qYUnmaivHmFDLMkZdD4k4IOzW1A8OyCKhLf9esAxpaxz+tHhPgtdBuglI7QLVsP8k
e3JfxB1ptPSAp5tOfCsYqchaXVcfrlaueJVUT7rUC9DWzUCpAsx1pJsGzlbIL4xhE3moaWcz1lRN
zDvXACkvCUQJ0Qb3tSg323SXkVAsSFSc8ub4JzSJjKMYCAEI62ifSC4ButPsUK1gbUoDZHSxk6wU
BP4is5Dere3rSfxkYUYksYuqX+W7A1/wHGSE2LbRpWC3wrqd+/FTMgHTZUtdqyKEpmDZHQXZN0LU
Ky82EwEdWD7bK9ounPJL0b6X0ERgs/5VO1HBIh1WQroaIqrfMGXJEoGkW74GgsPwYRRopWkRf0td
5UG8MO7NyFwQK2tyuLcDfqwpBfqTzKILaBYHKJlAR03+/Q9QBOfdDkRcNAlo3mzp2xf1KttzdbMr
TH/YsoUoLxVG3NYovO4igMw9ulrso9XwzucktMXwgO1XOD0iTpdE1ND/5s1dDTaiqRPfWpYZl9D8
rtWV5I7aq1sTUX+5jKhmPXKibN+GKz1dtdoBQv1DVdbakJgVA1L2kkeGW7CoS3AYjKajQ3vQWH1R
rNaM3ogOUVDw97tV/avEttOYgUwAfzDRNSjdUvo97Q9zjwwaL1MmRdvooIJsH2348st4sFXLfcfs
E7uN2qagleJkFhhEMRdYCqQPrQi721pAHvT4jfmGo/wEpBh3Ph9awBCVnzTuQ6zqEedlxWCDgAip
yHsm9rZzQy0iHEswIeS74pC4mvdAxAA3SWZoga8pSs4Myi+4qKsLHL+IuHKxZmU0TSqmtC1sOLvn
0jsl0lb9cM3Q8QEU0pRhVSUZzo0Cw+8YkA06a5b8lr4qolbfvfyKzRAi+hses1WqtY+BHUh7t2Gj
3Pj8z02Sz51A3OTvrwdarS8+2w/Z1qdZss9xTUnnqTiiSt0E5DKs3DRx7s2sIi4POC4qbvmQkaUM
7z7qEpD6d/l4Z+hP2XydbME5eVBP8l4cUOBpvko5aganCIxqNm+/GGmiXpWiTq3eRrgqmvtolgle
Tr0ebn9Of9XN+DTa1WAveXZaNr8PfdLN+qFpvRpRTINgSUzUJKDg8vM8rDtfdOCgvBzRF94/asHm
OtNPnhn8YnAZajRBTsdauyHKRlZ8rR0PyFOiwJ66RBfwfGxnudIc9AXbNqMOuzoh5hEzpw3OCYny
dDOGVbkRWTh27KOKZwlD3VIog13yjQ8RhziX532hWS6BjqcucEJR6Tn4A8+533aRhHjTerUUIca1
PYN5BazHVbclslE1GeE4Fz5EGrBGckPqYYewJESouTvGndSNtkG0J407qXSB9i7J9/ghADW7EA0v
4b8GYNMCfmkaC3O1/+4WZWm1WTTCtKXb8hdToRu4HoCHP6vtZ352JQp+hEAZiVIJq7VRFc/W3m0C
cJCk3SBAHRkWdo2CudP43bXl5YpMNXzOtSa+pExbdsxQyhcVllrE9zqj5VjGKUzHEfX33u/FfcjX
7sHrsRnGTKlmfakRcYZ5nN5azDpetPInCAR2O9MdB0gGF5bSGPMrEzVPXkhuWG0PnGDIVh2njQ4G
Er/0J+OMTtRKtp3sDu5yBDLrjXuIgtc4+6CLuDJtTKdAzwh/ED2scje7u/het7nXY09qaQcppW/N
3cTDyAa24+TnWO07iuBf+z2HdXcuY909uE5cjn0/qSrbCWKdxSUVcEYt8edth69lg7RGLd4lzVuD
0KjPWwze0us+Qf8n36QSw8WvnmDFC6ah7hZXWEtBEyNmT/n0K8msWFJtBUIc9rSm8yUdtcUzXUbj
NEr+ol0vqvZD549ZwoI3TYHTX2w5A8QkauDnoIMByWjL0J/Pn983DcgABrEgf7Ga/FvhC7Zo8z8h
fF3kzLMGA1OEWndgHoi4VhHUFLCqwXiDhU+if5Eu1pP2sjLeya6Nz6J4hxZ09Z+CNcM8Z6TgTKxi
KZYi/NOh8RGDxIDbRQRv8F2NyhQGrJEmVT60iajq1ZcnwcA3k+FVIODFD9YOpFFAMetKCIlyqZKk
nEGA+srUF4VJd9fptl/b8ZbX+MGFiNRQg0HwOiKzFC8X9eINjcAXnq2SKiOjF++6Gck1bHr/yUEB
8T5+dNtm8Nrmg4GY3uCWjAXu1QW36cSy8af99oL0IVlHARj13U3dk2bIaMiodTL9+QFyzKqTjs7l
CcFkhyeInwD2afZctHvu985XpzHQnYG+cNpAUaY49Y3IoJehUQap6Vj5iq7FkSRKtOf8K705nZFu
tcz2hwKQ+K1Fvrd1NRSosNqG/N3oWa4LMQBghqmGYTPq9aQmfgIzIsTfsCbv37ZLWMRRezzZ6APS
LYH3lQG0uuq5XbOR7K5i23wMRFKxSmUE4RJJfVjmNbUC7vVkpY6Rj+ok3d3NlfmRsbySCw3oM8rR
B625qWd7Ml8TRMtnjRsvKwnJH90fLbWXKVby7aqrlAGGN14L28oURnPhghaxH79fj/1j1tziOtAF
g5A1Bnm4PmjUsfDYAJtoblYz1ZvZI54T11+Nx9XsuUgVfATXFlGzwAHPz+APJiH1PKHOC27ZeIzq
rcVlNiXXMXBQtY7CJE8Fd7NnbKIJpzeAAwqmvvMGCCgjecicH5kVUMDP7HdjyoH5f3vsVstnGMl5
Y0HzqOM/Yv60EjXPvk963mfmvlc0sp4WIjEpTJJupzMhBEBXMKBC6x+aeV6SLi04rKbhW6CmGgSP
C/qeOGUYGjBJ0vnWOtVup2MvRj8Sn27qy8E50WbKbNRjjythZPnYiBcTe26SjnCj+WA22vFfCjoe
zSEcYKAlpTC5HlmTSW9qlNY1c/KkSRmXA63+IOi9BfA4eG1ZGYFgR45T8xZE+6ec84s6cJ1gB45O
hoj1/EZnuOCLU9QYYFBA9f/+r48lJ05BbRcUteSr8+MqhrG4sVaJ8yaEq2Ac/UttlvkCo3fAaaex
gIlsIMhG70Gf2HSPbYI7BTYV5ZVRVuB7uzlcpNY48Ph+eNS0d3lDO4cY/9hp0F+hGQb/Jyce0AC6
VTHHyNRJHWUiXqVwu3Vv3Sok05gJozOeCIt76viojOSPYAb7w43zBv/N4rUrYh+fKFBCh6vpda38
NS1Nh8+eRTQBnlMGju8ou8LAAqH/8JCnCfkpssKOtP+iYe4F+SPRkACcjahnMD/U2NSuGoiIewhv
P/sXba03/4oE+aCfxwuk8fy5BSskMSUNhetjeyOTAy077TMmHRAnIxsvYVFmWBy/JJ9A22RWu6sy
QU6LSR6ncU9ugYVyzX9DlVB3xQf0mcbepwaGDi7EXh9uIMAraaOGvIDId30EPgkiW5HvPRSvCoII
erufecc3Hy2Bdxo8O6OTwjSBk+U0nZu185IY/k2Vdnkk18KhiYBkGBpehcvi+IbNOPuLp4CJfCoX
z6Pdt3LbI6MYbu+gexzlHrLY+xbJIFIHUF9weuSaJG8IZW0OFsd+O3KB04jM6S3hmgLNKwzpw48v
mUoIFJfzL/YrQZErrR7reEHM1RIMVeuhtkd3E4nW2IVqAFRCK0qoq0vz5O3NU86RybcyTWmOywZV
Jxceor0WV9wmMOWZSKlGkLtmWWP7nF0TqEhuRpfieZfk9QLlTcnhBQB6HwI/K/zHGahkfQZDwJQ2
5SvOukirTxcKhQT32NSX0stwgDAgRHSc5FtpbjDj8uwCZ0Z9nF2ufvXYTDCRqurqPPZ/X3fyIzu0
kOKYteFfkw4vMBLyxkkY6UXzzlAHk/LD6ZQ1b+PCqOntRxWbqFyhSJY5qT/BO6rWO1jF+WunD2in
b73NCqO7jPcHIg/gTSWmSbpSjU98Kj26fk6ZBSddhzRBxVm1k8k+mvuh931sXvoWtwTqeFF9A7t5
mRxBKITu15hvjc2Ax/2XE26pDqWW9t+I0JIPJBxwTbJ3QDe0yaVnBDccHW2g0S7ZKRR6KJNR4ZF0
XIfS44qI7jCRDrEJmJYjwdD9SfqB3KeXDZNTqr7j7VANxOh6t/g4+64we5/Fb4HHTHuoU8MtP6If
UKOHRHtz+7KDjb0E3Wwutima7khVnRUMhY3O03sCEZN8AAwbdefrTweIcK0VOZbdsig/kvAsDvv5
/INjJJLcPa8U/sG4I2Za8ylBMS3nbZ0bzlhH60fWB4lKCnFtGBzeNcap32rjbvdXdiumyDwX5NI3
frsJrGHOGCYjvSr3jCU5pMEt35cc19tyMmfhwnWOa+05bHBsB5c1ErS04z1Rdw9WMmvu6ZqQ3cat
1Lz8RKbfMsIf6N/sA4wonZ4dDxmB/1HirzC0AXUjn9Esl5Yv6eBLZvpsuhElLln1mLhf6FzP49CS
dPUaO7FfJoIBDSOngrJ7y0EEQUc8X6vtVu+W/p7I025MlnH9ZQsEo+UA6GhbNNIA35y+YfS+qjVY
7h3JVfgdVGhGbyEeq2zkeVEKt8S2bjUcO+6utVZgv/PqZP3K+ktLrFjvukPVgnJfManzaM8HB0fp
EZAeNzgzxmBoyLVc/8i/ybqV7AP2b47rWD6cXPcoqvtjm8FRk+nKt96ur2aUGfS0rti5pMqMMxGL
0UfX0nZaLSW4bLIXR4ofb0to9JvNmZaUjV6pJuoEgoyecY1nEkm3Ltqpue4vRlCfbwVxPlxI0S9s
lHC2IXj2GnTBSno0gxHL7mRRCdi2zKV3mRqOwrdt7JCvPxQJylGhbTmRBInoT/XqyNkTzSgZxa14
Rx5nAbkvO4CS5rdigcupDSlyf4AjlBjZVu7WII6iieizxRDR1212p0T8jgqzAyxlZvaRaCs/cG0j
UnswtI+5Dser4AC+XYilHhqjGK/Zfxp88aqnncDEUXyYKjTS3McxL+asnERyYMJWZL5iJHyfZagv
mi8Vp6lsFyMsyCczdqYUMvpp/OjNcLWivaWfPLL73vjwj7ufvYvKlVCY91WTb+9qbnQX9mzcjXJs
l1ygyc51AnDurRqQhAD1B48jHWpGG8ioGrgq04EYQ03252ThySenIvjw7X/wXfNxExY9FTqADJUB
2YcNCu1JE8/YTe/lUqRmA8aN3ApdZGzkkarfJEsZG5xx4U8TxPVMbxgCL0QOcp0tJK6KA785Wy+G
EdGBd5s9NlfG2NW6xLWMnDU3E4Zfl3AdDEKljq6pPMk9mw==
`protect end_protected

