

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
UXXDHK9d3YtwspCksVg3cn1OQkWFk3QQ1bnN8kcpv130B5dMgVD8+qx+9EwjTR0JFb8FYrcL/7dg
lIwdmlKGHQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
lGlirTrah5ntgtsTqcFN8kWYeCxRHbehSLZqyiEvescJE+ORKShYIOu42/ExCc8hSawNVl9qCirT
UlThiM+Fc1evKMQYzaFIzbKiio/Xw8rjRfhTJKjaxdK3T87LnrHcsuSrci+tl+anpBCM3X47tPxD
oNmgZzATBY/NVtZsbvA=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
UAOAU0ylQuQrszr15mLZsCg4shnqFlxQBAKcqwUoJfM+lTESkAcOosPqKsRH4IbbLlaKiP2HCFU1
aKEFZccPWIgd9WlvneNU3oFbpPCOyV9eZTCX4e5jNTf/7OwRRATKc0mjpd4lxBL9xFrSwNaUKgs1
3vjH77tdesEDAIn5GZ1C/7l3wjwnB4tAiaRNqLY90lB834tlc4mPcP6x8L3rhv5EXfqU4jyJC8B1
4zsO/vH5+VVa1595cRZ3xWXEGVMvmWhY+6TDUJCMhztjp+p4kbQ87UqJz9ddvZWB4hRfjo99Os6I
PqyD9P7zikHIa7jafFMtZu0Vj7u4HDelVYnPyw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
qRFhWXCy25iIpt8SG9Mt+xW3HRp/MFye1jJpn72azeuP+g/A4uHCFxvcKVhzcuE8lYDqFZ9IBM4P
ZjcyPOhURivBaWk0KosUyfzbkORd8yS5XcayTSj5/d+90PPk5PXVCLjTrcMbg0+NO3tiyKtPpLQJ
f+Ih38e2az80fHBgiqo=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
tjh0p4bhQQ++Enuq/zxHJnIk+bY5nNzFWlWKnTVXUtnLIlVGko6ShpeQRaCrGzeMC58aHThmj0Rv
eUmPmT2uqc307TRbbuUeFDYMANj1kcC6Ygs+bdXnSkWnOQFu5reSEq5SE7OMIvzdCIaR/FDvSj26
cuj56WGV7WVTg7EZvTcQQsjBPGe7MBQPj6gVbjkHGUTFOQ09cS9h1BaC9UWWfJNQjyJE48PH9w0J
tqmbE8H5AkyiSVZzE1dyYA/E3WjYX0ib/4FRIxCW96Qs02ypuSbfnvJpIyeRwyQL7ko2qezd2p0h
VgIw3omrmALcnzzjpdcOgkkF7sgouCeIApSqBQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 51440)
`protect data_block
eArT0ITHLv7/yuQMXdD6DuLj+QCd1HcpRz4DkST1XI12N/LEZ1PyavR5IVID7YRl5hnz+fsX/OH1
5CqkrIq4yS5yQWppmwmtZlvLuo0b2RFlslZR0xRnE1sfp7zUt2rt7X8z2VcI08Dcv4bFraqi5Ohd
tayBFIXWuqF6YV0YvLnv/hOUNdPowLLhqvWXPFrYI79acQ4C0QEibQCm61PgK1amyNu1jeSMmQtF
PL4tMyBljjGmOmubfw/AcixJkQamPNViBkjrSecsahprEuIjxKBwLj1wBKlSOHu50M85MZclo5uW
vQy3+y72EM29iTM1vvSNV1Z2PBNmonp+7AoI1FJqp5Jy4S/cSnW1UTyi5A/dWsRCHKDbAsLLvHo/
oqV82ZBep1BSozQ0AU7rPhteEFJ6xT180wkka2FHPkHYSdEZciQDMonGweFxurzLJ9t/mxt93AmC
TpxuhFHWDFX+deMdbmx1+rvmYpdWA/XxVpn+xaOM9JFlyYZEVBDTGC5O41wqXpwyZpis6gZXVbWG
+lzzxDL0nFVHVyk26vUCZPtjFluThoP6LA/MoLCQjL0nI+TGthmJvhWV8pjxyVi/PHE28qLBImBh
8BJCo4W/TTtSJ3t0u/eAEwc5F2nysZo+SvP3vvhqgyGEK21a1SpqzjJey+PHi1wXOQlWkZ/GM6GJ
HUEomtj0j8CWxhKdMWIhNs8UlUqRNDOE1kFYEn3sZe2hPCWwuvqSQvFYnnLuQ7Ion3J+DILcJEao
unO+fIbW0uNYI/NVIKXn/T/v3IfUCCqJpKXxBPk5n2rL24pZpneVAfMdnGIF0JWtwMH7h4PH0JBi
pR3hYn01dlEf3A5AJ4rgD48ZkaqakQfP91DUNvJKo1FF6BR7lCsHNW+L6y3hd3wUC9QXhDV2SOt7
GBtL9q6xHkwSqEdeZpUSopnqLfs7j/u6huCDgKfag+K0HUqkWl77y0W4QojYEtEuxRvhwWs/hAm+
bOYQC7OYpJfgI7gyVmgax/CbtPdZdL9/jRQ/pigjRHI+OlGXDJr9Sq6PrSwtwapUt4XFs5q5i4mc
TCUmbq45LbSuvzh1RyzOzhc6zrdIkx4N5W4FimcqlZ8BZsvQ0u0bLqIkIHwuAmiM8UwLBfquDtir
+8eRBeO5D0pwy5ieYuSF/TOZIkKn7hsKRkUjdfmhy8tW1urNC0NB47aazGhxTeN93mNw22cn6i0l
JO3Xo5W2Ew0tkM+HwQnM6hBkLVt0BmjEdAAwDziUTnPGWlJmzWOBDv8Ck3leN9HQMECa+zDI1jtC
UDgWbbpu4IEQjAjjuVk2/HOdIKdzhlJHnBa7dms3mumC3BqkKfinltH6P+WFH/7qmbq8aPVjAcTg
fmd5Abym0ysY+Zvw6QOdVwhqgjDb5r8msR6XesACvDldJkRwUJGxi4ju26cDAF3INfO1n6cgS2Dy
p1sLjgwhpus3l2GtqfJb69cNK4sWn3TFbErHT4tFtYtvtpuYA0K1bDe3PedcPlelrzXAegKsQ0M5
3u+crxrJnSnk/SDIzBSLii4/QBuUd8549/Vql84qgSBynKxdM0PpBszVU+ME/CkMjPd4Ox8C2hIc
6tUs9jXV68lDX77CKFOhj3nQktYaPsQ0Yc9PCobvRGYB5NFcRYLSCXCm/cFfcBTpQMUF1xepg9hL
60ZBj1QzCpZxyIQkJFzyzEwTrrDXvfrnD4ZfrNuH4xbbdu7PSrYQ23492YXzGu2CICkuCBxaqg4b
nu8s53/4RB2E4G22gOvlmlkKGLfKKu0pRh2Zp+OsALrzNftfHfzPc1hYkeqqcvfqFXBsDcryNyeI
Ud7VemECqoCtM37SnWPBWMZbhzTPGW89ivEPYXuUXMUpNmp8HRMOvc74PriehEuciLWsPNRfMFHS
agdffnrFr3bLak93S8HqT3gwQDwXojKvlstHAOuDWU4ARBPcl9ZU64fNWwj1vO7B+1TIcxbNjZU5
BtLnwyV6qbEnTQMh4AONgJED2W3ydHxKdfrrOxKs3sGQE6SFvXprNvPDtUOaK25cecTM7aqGzPRe
qW/8IoDCtdoxbH2+PXl9sL6Di3hrxe8v9KL8GCjFuxOzvM296me5+nM26Y7bvSxJOF6yjI++I8zp
m1qSf2G0cawM1EIeLTJudS7l1vAGrTcWtkh1fn2GqpCJzR8SSaWekI0/6MhTnmUcjJLP328YSpd0
S/ziN+fh4EFCBG/eQdHySbdktNPcmEy5aurKACv8yMmKtibVsQ6t5AzWYYrfYK4FcZhfVMrzMaqr
igI3Fv2uwDShoa7VBJ/nkF1JVGcJeU60vsuE1wRN0AYFH6s14h2jCVC+QhkaSTxSqIID8vMpRcrz
PYPe2aHSiO3EuLPULKnq8UIWZv6L6c3Tw7NdInLJdYzl5IMlZsxociQw8qfNc3600yHp2mEIZAK8
qJhTr7k+bFuIr5ct0ZSCb17aumFj/1+f5KBdcJ0IFbzt9OV6bHRpoWmTdE8/MhW7BrP0U/RDt90+
Y43Bu0Cumvp2MwD9YYJsWcFHpMpUOQbOoH2pDIcW4K9gNzbjLk1Vv95orDWWYH/Mu57EqxxMD1eX
RLZn4uTrkMiBf2hK722jFLhVVQ0UluXU6uYJJaJmfcNShxxuUh1gsh73RhlryNB9VrA2ntIscpKp
sMIGWgZm3gTOdGpUQM5aaUjjic+FIlNV8c2FxqguGG/pV6c0crYrxl9evQ5ah7M1lR5hYUwnua96
50w/+H701faFfLEa/588o9bTdMAkrw7LlOdjLYGaCldBt3Lgjt472Mq3NLLdVX9SRglwmJWncPE4
+PDcWWlr7YroBep7ciCZWZBhRIRMN0ZHnYjo7dACDunqYO+SHNisuH8liJNvh4VPLmvw2vd6bfeb
OsDlV0jjicmE00rQbgIxlL3Ff++sMb+tdMT60S8dXNt8g7XKZInwdVFUNGol4MVei+6v69V3Dn1J
B/3x80Zu0UJzHk3hsbf/MQ6Tl0d0fUvIMiLRNiuKa6j+aoJgAKiNSx2VUGG1fSRderhhBDMajV3j
ivXhuSb07DVwntYbsVWfltzgx/Q68KqwkFWs0h9rukTFJo78JvkDftTQF+0oqbU7wyKy8Ixbf7t0
DrNC6b/xpx7k4efhbDB8/McNSw8obGB8Bp1yTBGcfCDk8G3znXz62hsyixwUGqemt/SrazcZsdbK
j4cI1ALNgjOK2dQVISmFYqElTpL2Q0yIo6I/s8smStzarp4BB77qq9hprqFf8fOuYqm9PY/6hITE
/qoEPanFZmNO/OumDYpSwiuOwSM15hsoHXIz8Yt0MQY7JkhQyFs0wiLF9VsycsEtDLkNImdUiSWy
sO8DWl0b9V+DCcRjkrMOJbpouSKYPodDNnEwCkNM0ncqARaA6W13mt6e1IiKhSB18c4ggXSoxllf
BPPvim0tT3HflyYdvQKNWSlc/mJP/S/+HYCI0Ube80++8Gx8DE58nx//tFCYctatvIy+hvm6Gs4g
AL+Z716zCWPeFsPUkNNerFTIEDScEPhjOv5nbUKd6SbGjWkbmtsydUQeCaA85HAbDa6q+2cxk4ea
PXIsYrVbx9rkNFEu2d6+qXcs4khpdkxO40S+saj4jQd99w8akC+Vumlf0n5EQ5spDwJOdiM477bs
IkPzyO38cX3cDnNDL5whJsxousIbCm0BaBIpvLMxoqF3liplWvcGPlL1daZqevNDyNHIVTO11EPs
madN1xA6YZPKqFa68U9URYaoBRw9W9WQhJPiv3ITmlosUTQXiVmVOd85kZzUYjXKC7l8ppHg4/5b
MzAaUXFlV2M249ayGdgU+GgKNLjQVxGENeMk1AXxG33qTcuXPm9uoRZa0JxcM4gHdZQFyBv7jNnp
U1UsTZY13y/vK7bVBLETT7ONNLWE4RTHuFLa1Qjw22/x4tHakikIdxONXUpz6KYbDJDIuBauiCgy
jy4yf9SMcpbPtdZCqL+YVKOT02AgcEYo71wFWEsfiMY/TOlMLuUp5WxUX/GLRHQXHFj2BFw08LLs
+ZfCnuFTNKAI9whAm3u+H+TrdU/sYWxWOI7arQpMGknrWKjwN9g2BA8j73omNl7IQFJorN6h2JJR
f87grzXEcKtdwJk1MQL9+tLNHG6lrc+Lx2YMGxums5WTd2iZCSnr6vb1fmqdFtANgNlIYoQFphgP
UIWFEm7fVHshINRospYMeDEYEDAb+LcbZ/Ax/loMW40RQuX3dugxn5TwUDi33XPUTtR9D7xvR2f5
FAynBACzejZr95DNVPRcw4+83uY1/98cjz0Le7oJZstNL0LfH0ki+EG5dPlS3x3j99xIYiDc2w9C
8bjjpKVzpLEcrZsbAxT8gVUy75L1MJ0vJSRxL/vjn59YiwHFuIvAwJH3TNnxMxxDPJAj+d7hTrjI
gNf6NCA2CdVt5WYbp+eonn84nYhCotV5N7iiA/ayaFCjpm3ndjQozwow9CadWAAoGw2bBle43QdW
2NT5hBZxnnMk9+KQ0M7A8QNw0bzkwLaNWHsc0Hv2kuYpNZShG/yM4DGKqrZRNjGUaTQMAQpvA5ux
58Ulge3AIyV/b82qumds5ecyLUTYgUbCpiJfT9h9Pvq4v4GZnHgSXbZFdMRrsYHDfIecluh1440s
yzmTulzDNgufjtQjBW73bTq+PCZaKBLx/gx3n+fpRJvBCqH0PWUqCCx4o/QfXp0ws69dRl/nzOh6
JsVYPqhWMqCBWoYOycj/2IW6jheAFAYAl6BlFFwjL3e4F8dwDqRYlX/2vKvN0c8c65h4ZUSFAZck
ncJdjvhiSwK9YxKkxaBNwcITdqrz7tFzooQiwjvk3zI972adUvfRIWX9g/VYTpYHXhdYnrd732gE
ixAyeLwSUiy6TxLjsTeJ4HEs7QjELydLa225jx3uoulHxSmAJr2QHoiDfUwj85bSp5vHHTHLlxJF
qQphdy56na5Xkg81V3iIpDvGo9R71l1Mcp//pbivHgbXmIIJFCm/Ywf0v1qbVwqlLDmfOI5mhskZ
KULfAPoxTGP5Yv943jZCDz/n4C7FCmCDQN1PolF4cooYr4lQr7SUV/fuDfebmwhMHgfQlzrEIoX3
U4DlbkRp20hun8SPm15ZuQcj1EF5PPvW11Zi+rGKADGypG3XebP0ItRYblBT9mbdC2sD1qVA3msi
HseSTaPMR4YFUs3hfpgLqm91m0Yg4ONd5P+b5vy75X/r6HtqqLx8k0vT9J9hIDdCwLYwq0Czr+ar
wJjtV29Tt2gYVFdB8rc8ILMI9/CxRGAlOi44kz91tLlBuTwf6l2RNw16yTEPHykAp/D7NkDg/t4C
V3PFcVyi04MrACOM84znQrYWBoSuADr8L/zWh8sxp0BzIGyKYAzbGsoorT85Icoxg6RLFByNaQ+D
Q450dXt5SKUaTrKUrtmnzbNcIUmTR/ZtL2hgXNDQhAAEACH4oi6zc6BvDcjLr5urqifsUg4nBLHP
ZM13HOu83rzmBSGyNIl2zA0sZ6nNLtQ/wxybPK0TR+8wZ35HS3CClcphhsX5WhgBWCj6SNC868bk
FrXEh5Lp26EV9W6BQ3LU1KyU14qoi0t4g6AyvWdYTtwox7ua6pI6UVQAMhnv8CRyburcUp7PrxEl
vRn3p4jGjl8oAUCQcQCLWcArC/fo3th84UhanlsSRrypGzdHLtvLJyiA+4VPKE/NRwC2oYPUlOuf
EYjy2fJ0dA0cQgJlpnQDGx53wQgV3egDBWpoLTKdF0NmQym6FblccONHeXuXV39AMq3q88EgHMe8
JPgpYnvHK0Aauni1oAw3BlKxSocypayBX+adu/sln17oBbY1WfMsGzsNp35WCirMgKF/vOMrmvYj
s2UdFTZPEAVEYfaI6IOZ37rKYLm/vI5QsLFjNYSlQLb8WKmZIiPfg3TD2E4OWWWxntil5+IWjgLH
9BkuRDr8gah82dRFyMKe2MozgyLGZrGzWTntXHbEeY1K1VYW8VWbJsTmldy7SeP5Csh8R3J4qzIU
wH0x4X3CwsbyuEARgZ7FVW8HEMznAmmzeWoIf5JIqVuWOlJ5YAra3qwUiwzdL66/EOwxnqzbtDUF
37+53LjZZXzKZHWhzeBL1xNreH2kSg5oHQl+rw8VfPiToH112ZvhlzZDWLGONDs8hoK5k2uE00pt
JcZdm/mMY4gBbBN2L87ZuZjMpf2h+UWKfxn+Ph6Th0P78DlIV1U1np5g8WiOnrUof3MAd4vk9Qcu
JlVADbOdbNWGDb9JdeQAWWrA/jAX9YaX2Gre/XOC/nTVQfRpNyjfofG63mqAdUN165au87nHYGEG
DW4ggwTVjX2HVmenfY6lO9/Y0o3vmJnktfjphrSkPpeqKkoDH08D2l0EnXfmTRhPLKiuzu1SoIWX
J98Yo3Rbn7iLTaHHFZwxNC7yyqMOpm9LqfW2YT8e+YA8iOl//3RIrkNgyE6RPfmL4T7V3JppYJBC
RfLYxloM9ZH/Yl7Exl9hPc0nhVCmbekOcgXe8BnJDmN6pK4v9EqwAMJ4Goy+xCsCwRh+7nnd6iSK
nSu97KwXfxW9Jy2rbqA4OmhwKwfyQM3qbkwRnuXm11tufKV7PqvKYU9raiwfBG3uICq24QRQDTRS
I2br1akCIItLR1+hyKK1q1Kne1Evthvp6qdOODY9Ovzo4WQwhwYUUbciyGRNpiE07ePtlSev+FQW
3Y9AI/6CP4qsLOCPgjzS6bvOr9gSDffWU8xu6DbVk2qeef2Qel9U72KGxV0HCQXIwo+ujWj6QJiz
UtMzBzcc5JGALR3CNs08pBel2pt9wkVoLLl828rNO6vnzGncmpE8B5xyHQlwhTkxhOenR8pu6KuR
6GpM6aKjtoURoCX/E1PGSu9k0k7hTRkWpGtU5P9W+257nryZ4raYkZVnaXdNNqY1jbnsTqbJ6MKB
xhUskbd7lpbeLCSDwN1KjBFd/uF/fnSW9QgSCuHnqlHtF88ZAbZA5zk1UAHACU00BlpOLYW+26c5
k9vcpZ0ZK8ugcBY9C+bXQsunqwYQz1VGyNS63xkkhM6N4T0CROghIn5F0eXdQu4076AUbS6s+k/u
t/QJJ2C+T6dsZt9cQaXiy1ak5dj4ftSj9fKgn8bxKkQrPH0/gubVVwapNhRBxW63pJYu93NthRus
1CuiR0J9P3MAusRnUOpvMbESyyDLpgGQDrLeoDesT73o2EUD7nYRKYa5roZStiZrZZ0khtyKx8ei
fdmM1oFGQBG1xef5GpVGsqA8QOAgFgGc0UuNrmyems3dkW3tJ6LTnUqLtUm76F41TIlRhxcHUTBy
u7eHDHJx870ARvKS2m3p0j4auUVtHZnFM1/QEbV22qdbtuU6B0JfYOEtcWgWeW3yBQ8cjY2Oj7Ab
jntuJCBwJGeiEamecm/xSQuxaoacuZ2F3T5HztiUf4TTESyk3hbOfao7zNwyTeVQvTNaUbUn1G22
VyCTKxbTGVpJSM/aMkAclhA7xja5Q8RM/gKIeYmZn8jo+l6T8c8B0XyBnEmj8YGXHsX6MtR6/tyS
il7VOIj3rw8xJp5dFZGuqqmktYFCl8rbE3u5SSAJDbHPlORHjEtwgDguKokC7muIFf+7NhZupecD
IgymyqZH27ajTvPMGIx3CGwjPFkSjct0VoFlJoQgLA8yYZAbJ6wkDG36rRUDVdHP0kckh3zhZD5P
AhFBpwIWDYEPPyE37F9DcTKagNG7OxdnIFYzvzyA8P/Keau2ys0TgbR/7ItMpjDx4coxFJmwij3R
2v/pVKFako4av9DWTVWItZxfpJpGvFrrEAf2CY6a0OBg6cyp3d7jOJLCEyu4kZvWapQ9zFMMd3VU
XWN5AKIXqNOGqSjmy26QgbCZDuDBcaEzpqv6tf9U/7T//Ua9VWcXDqu6WX1+5rA+hClF1IMiJclz
fOVcVOHHUQYifQszmeXhs2AWunhyo2ayC1xxyIHM6Khtwc1q9+yBngqrY7NJmziN+CifaoKmYJZY
GEWJtrUVdVmrnpaumDh7JZNyg+SRw8BnkLCz5g04glGwybXUi4B8XU9rAGr2fujoD8cuC0s2o1eC
3Xn7G3FEs5Wn3fvGbFU0wBOu4kOdz/0Ti+dge9/pT97xa6CRQrvScG/agWVX5GjeLxIjPN2aeY0D
0/O9altrhdsqTsDzpT0E/izao5Yvtr6HnGJ9Drulus5ARgHopIL4Zb+dR1/+UmEEmMa9WA8PeR5N
yTot+MzsuZeoy2M0TqGvmGsAd0NTDvwJeJwSy3VpopIRy3sNnXHcIPup4kKbI7JEwF3kXhTeFWsn
int8HRfKXrYundHtr4BAxUXCJH9zMeukuCGbFTndummR1x747Ouz9KuSDBAniZCmHZ6hQqhXAyvQ
ixe/v7fYKy4ZUgnPUCzok1gz5qnagQSbJ/BgcfrmBx93/P83g3YqRLLrGLP+BHzUWVEgK8Td74QE
ZTyLb5hzvAiIvkujM+W7OaT0F3h/GXQa/OI8rShIQKCR8DLeZiCTb2VpE3yrXjMJBOYgKdoOzwUv
4EInl+dtwmzGfLZMOitgyuseSU+aAczEnjK4hrcjy0joVlwSTRqfkhf0bCgKLBUqh6bbtXkeIc19
AT6Qj9TA1i243m36BIHOZHiSD7oCuJ2W1L6pFtlS8aSRFWhUluC7m2i4WSK5IzoM6JlWdKZ8gBQn
mCH56RP85oyP8BhIB8yfsgzz29XHHdCSDytSeiQtptjoxuMsFA+oYdV1hQJYE+I5Ad+0SJn01KJO
+NzZMoss55Dc84ZlLZft2MeBrOXzqQSgs4CU+vYEuPJkA0VEVXDRJgmgyReu/Cogg532IfL8x87C
zlol0vczJApsn0itvxo69EMXvKyfj55JlwlSf+Hd95iCQEClSMqCwPeft9wgLqcsstY8TotGTaZn
4wAOMfqAdLsbNohIgEHDXWPz2NLk9Fvd3lhq0Ekoj1FefimMSh4DLffoCS4FCgNC2t1kd2fXImpm
dcHnKPkvwGDeYq3/v5iAWglVun4BxVPboPIo4lRbInDataWUU1FSOscr4Az19nbhWvQY9neBObMu
T7bG3ByGoVfqX/FVLqpnWgw9vnnDHC+rhfirFuMIqT1Uoax9CUN8DsmMFi1Mg+X9UpVL5ily9IXK
D7gsDhMBWMIYNBDezlX2RUzRnVnRqKbA2nDqdZ++xe0p1d7sxJ3Qtj7JN9iI6TVoqhzrYsKuJjbu
voGAUF2SwBpH9axlvNVokPYrTT29urxHObgZ5zFClss/+uNVjo6YwneNl+Nl0bU+GIiYXvMajthP
iedzNxAMvBO4D659w6WOY2tK1KVw3Tp6pPBheq0QCzUCvShZlIYXLbnwIz91cZinzCVPd/EedYLL
oOPHWsDrOEqob0uOT3nReDtqoaHPz5SlSU8vGSvscfVMLgiBdXDTRaKXi+nsw5ZoEfX2qbeuojsk
l0ZC21jE/+VqK9HcFjyi9z3/NLaPlVWigK+sg2pu4/Ej+gUmsmhHeCama3MZX0/zH2TVmrWMxDjD
R38GWRjJ+3yfVu7Lyr3peAAxyMlGIC4KjLKsvCQ6506F5omG74kq/xHAMaOpXjQkxTMtIeSlp7Ly
3NFTyAy39wxa+HA8a5KgeCWYsJAMVElVOm3hsCNOWNLPM6LH4CafOFEniatj9VVohk4LcHaRQ4SE
k77qr/85Q6oh2UWFdYb6gd2K2h1McN36Y1KzE+Npx6Cj1wosInutsQ6d1h17upipmfFLct8ZV0pJ
GL6iiUL+icpCEg350dA/AUDafhkf3jUlvT3NwmRbRH2VD9glj+vHVglCe/H2j6o1t90mTeJJcC7V
Ec0r9lWDNltdNHocqzMQFSOK3+4XemwWbxZKdM5R+11KX+rCmqGYFMHqDEKjt5Uy14DKO62Vjz5P
R70lJbI0JXpywVC+6AYAffVOKu1Vgi7ujf1r0rTloJZ+iHohzebnOtlx++jXtJbeGsVWjyFLpz4Y
lJmnx2Zr+dZRfxq6yzuCCv4sAkGX+v2ywtM8v8aNJRlrq1NeDFM1bZgN8yvtYdhj/QoM9dDpkMVB
dCZxb0ix7htWcMIsIm99pwGPomGBCR8xd9HE5kDfioWa22TViayJthYqVBw1I9y0bnXSQwi8bPHK
QTeWohuZayp2HJf1ZoM6uouoZryu7RHVDgWbxf0biDB6L21RBAA5jE1ljAPvfqekN8ja+6IDCpQR
AXECVk0Xh8cfJWYUyYWhijcXdLdmmtZuvieXQBsQZNAhOe25r2DwJpaxfs3EiS/Xuqx82CKUcRgs
xdP/8j5AgxYIqq3gEF8VPtlKVq+Iy9lfHr9fgk1DP2LEKw4IEfbh/ySEdWkTjLKXXwj/mB0b4lOX
vBpjBqm5re69uaetX7KSE2Bg84y5Yn711hc237iwM4cz4wIrBnphJ3NCEqRzqmfKkLreCi2yU2po
/+rCdrAr4WO8EjOYS68HXtAM4tgNW4wRUjXL63vHBCvIbjCn3ze5vUlmmHVPZHwa2ArgvtEjIAQh
uziV2KEO2Qn+K0tMGW6vdi7yE3s8j5SpFtxI9H4uKyUKAcIQ+THKnzB3XdiGE0JcR12eJyuH1VdZ
FO9RLssRP4D4bHiacQccEr5yzWCXaibumBmt6ALh6Y9xZ0TNIb//Ok4KHVask5lcs4zHYAgRUhRK
z2nCUWyHfE98YqOxgI6QNoVgtJYg9VZ8e3jZdOAZtzROTVVPw7J0cmkXj7IvuXJ4FrqtWXMwN+Cg
JArbOl6D4J1tf8lTGhw/x4VoRYcaP4nJ8FdRg0FKrZ3Tf6zZysNNblpWau6j6WYGI52+i6gmnAzT
zyZ6Eo7l4AgCGntmop8Oa5/ejlhV5neEGdswmJf2ZYcROuM3sHEVUfm+Y7KCTTQ7q5iZk/LHoBt4
LVv9T5J+0TyKv/P55g8j6GmmD2qhxWK9qZCx0KLR108+xwR7mbS51iSvLjASzwEf+fxhZGHEwPNm
C9p7bDb/Ly0GHDBWTYAUNDcOwJomLO19oAak0wf1Oh2cK5VUHbJf/+T63bNPcN0pv5UNjtqdbEki
hyOEiSdqN0AwsIRwucUbIFZC+DuTp7mu2EUz4Z4gJ4+fjLzju5B+npZN6K+Q+q5Gy7sbfGsiWIYT
SVhXZoxQMcd0sBErMXXTB9zJaOaQ0Ir5N5vDDTSTsinMQjGbdGJMteJPMtVEumbeRh7f80brPRtF
S76ytXmIZJRP5qAYyLv3yNOvO3wcKTxoVr5ejkJT2sc8AAdA/E63v5R8EGc9AfJS9ZE//yuGYtOC
c7rO7dhdWJAKJ7AvpmLCiQNvb4NWEpJ2vp8QUB+Xs5jGj6AneMe0ROvs1AOVzJl8tTr974fiSoKH
AtKfaudWq3moDGsnayDxmTrrCzu1DyUVXlXVGqES+FJh6ge1EXimXjC9A3PalDKJFr/N6itmm8x3
fBInCgiQA0q3zswsfpLccuXnreAtcyBPsK/vv09gcd0GEG1pjGfSevR6Z9XW+m8OI8cMUzg/AglG
uavFP9wKwluThYII9OvESCbDv1nxjLPqkmX28jb1S/lgbPBGiS2tkR37itAa9Y3y4XfesIhyfMQ2
7JciFI1K+SF+oE7n8jOY03ltlgjZHFgJnj30RnsA/TLXEdqUx/rIwH8d8PyLjlUTGeUlUgvJVOEv
2FfKo8GjyMZv0VwLIeCd6sjlHURZcsUlOFzLWLThMF5F/s5sJqu41J5GTvAvOsnQa5DBprKM0x8X
WSfSqnkYYYO5sVEbFCGmxqP370pTO14f2/rpamkw1Y1zftTJsKvUukM4iOpmCYMwD18iaWFYEKuj
FQQyi1OpqmdSRiM5ALlFdKxd/BKCRe4YsIgpfODovwdAg1h0vAelm5JzQRG1oxbVHAgMUzz+jh2m
7Om9X4KeULiCQe4YxV6eGNbC/vL2W//H95u4SQPXbC3qii3qW1fqS2aX65rJEhElwub0jT9X5P+0
VbMaxjjaZ22vzkelM2JJ0iY+VARaqlaNmxQEnygPNJHCmW3ndO9REfENGj67RG5Ia6U1c1Rv6x0/
a/nGSYDBOkKgA9YCBpJtu8dxE5QWayjb/HsW/rSRfIa5FB4qVOajE3DW/OBJ0IQKjfWPRdVUI6HY
oC+IUrLS24go8oQ2zqqpAyctDeG+aOq0VBmmIxjV5hLCaiQzlb6yLIzCrRvpJdowjoEYWKBgUfuT
GVgUvgUzrxYFGpMtARXT9lp10lJHoBUxBD0m6eiwzK0pGOuit66ky2Mx8biLm1o2ydfIWiWge7qe
esD+FmOXAEn1bhzFaJn5pVDk9IU9DW3+nw1GvOYTdbrcrAXKYafqPdJT8fR+3ZH2gB6pqIcjr2rv
QKTXc3BAaKNW7XnywFB8BCtEzxHcn6u99wjTjaHf9HtE2U3DUDr/Of8Ml5KoMCp80KuVmT8nsu+3
qgSUl4tD3KRkEwLyYsXOh+D0cLzbh06N0PCYbpxMsDgKzBVRBs3C+iffB1+rkMcMairW+vvUA2ek
sRL7MnwtI1moyF1++uNkOJOebbbV/FM8ivf1eKqfb07Ahp6Vqlk4Z8g3jmEMpREV7oc1P+BpqN/X
HP2np2c5JiBYS697ruQlKLBVlKvhzZ3qXOhzHxPTw0gq4H+cZKwTHRZBZBIj7IC7jHxjLDLR9ARk
Q99fpXpnWqJVtfrFFm0bgScditTrzNdCMbDDGatIBUGuuRJOHhfnRNEH5L0efj6H0bdhgpqJHW5P
wsABuDZGBsMQrB2i4G5Yx11GsPMcZc+b6q4cERlDUsW+p0qf87J+7RVkYxMYzp56I2iOwVDkUwAa
4Iy2tOZ2aDmpy9txkz4/WiqsAJNojZwiGJiDPGza3Xs4J6EZwwDmfHCNRUGxQCUPsWxMDoZGqEBC
FbV7RE1ec6Vamwo8kPiYjVpGxBP5RK0CZTtiCVdYLUcST/lOxDcOq5BiMfRe0Sow7nj55sUOil9k
CrIRQheeuy1SAvq1FbvqfthkjNZnPwqfowSYqKa7JB+1d1iszWSLr6ebBssnLnnVDXyPf+mL+SZS
hGBYnNniQhQjS4pVAqj2ORpWbaBDhGdPaNlxXcRwE8akzgsBgyuI+tSxkI90UbDcCx2UZHayHN1o
48LsrrJpiaGX5WfiaTH5PemIa/sPujYalmZaOntCu4rUebHuZDlNW5wKg+JINGjRSkJofUBPzChD
VXPssHfzOGxS393zG0f/iF+k68PNWWPc2dLN9Uwkdac2BQb7tg5EP9FboWG2vpESZOy9T7gH3MC+
BVq202aHphPf7Gxfx20KhGGu9bhCeg0+2tXuVzbfEM7FEwMuomW83dP03qqKjX+94ZySJeHo054U
XMnksEoCCTUB5+ZaEXR/TSxUHKbs/9mcBfXaabmh4of2XdttI4mtrd4FS2KaY5e6L6SbvDQG2Win
e5VPY8w2X3x4EutvD5zKWnlDUsytyOVXIHWTcK1mKf8f3kXXaiVy2yvB8ZoLL78u5ce0FFABg2uJ
xfE/Xlkl5QnRgxl6oiWApwfIo1E3AVXmlfG1qVdM/RGc5DfHrcgi+d43HaIUhDz3BdlnhxwX9g7d
1r+n3xDJEGE/uR/D0nlgspY99f+EEwzNiBaIEpRET2zLYPfqPhRxIIIOavLxBG9Lnp97BNeQEuBL
nnr59X39WdBZekO+W2fqtDabrJxZddy9N1QspyujYd6lBGl4UpRbS8n0OAR0zca0uegbRDN2TvC/
SjaluuxBeI5eTCZ+qHki+fVDXAr+HF7RGMceasJ90lphBHUXZEDbI/RyXEu8Ph0pw6s/EmUgysWA
AiQd+6a1foupz5FB3PrM5z0HHSe+Xo1rvCUv6mcyCAVPKIwDzT6qC2ElVNfDaSueufzYBFUAgfng
7Ko7XVzUY5mx7s2AK7NpbRuQnaUKc5n3e3R9XNGUdjqvZx69DUJh8CSvJmPPUS2WLFafu2dZxLrk
/q00/spqx5ovcT8tpcbGK1+z63zYO22tyQ+GCvNAuPVYKMFmSjqMt4Mwl1lxYDwwXIiityu+pj3I
VW5xZ+7WUEwhcWlB34rennq9k44UbqARaV+IcVDfego72/Vlr2nJUl1doaMl46woRXjICkdK4+/N
psS376nRVhHieJ8wjX9YaoDmb220ilQ48Ipzc8J4acKghJI+TjcfU4t1pW/Vfnhp5JSgByz0MRSl
7/rOqNZwUD/6bhC0KLiswfF7CiniRTalkh+RsX5PgPbeNZpTR3pGKs9nslUlKFczAGlgx0OiHxDd
2Vb4uECVSDx7e6dk+NYo0rpnqlI/RfpiDUsdF99IyDF8kgXO4x+swJ4vN1Mxivem5tGp0V8nBa5F
5i9mx5QdcOPokse73Qs5rVxyT3AU6diz4aK+xCeWVicV8YR/+oauqqtKALVb7mMba4j9mbEYS1Jb
tec78hR15QQ2P/eUO2gcsSnkBmR2IxSItzzA/aKt9e8YbXmViuidvn8J1fAvxq9ZjjNDdc3xT9xT
oVZnyFQyQA7104b4aDnHDumu7G+drZRDqrmmye46IxMc53CNSYFtxLMpKd1TH6/Ol9T4pfX/iR9t
5wES35k5VQYLRSiVSPpkNBPAquUfSe1f9/NQWPDsdDoarE8B3u9jeRSBJHTCDhCka+FKnK20thTo
1XmfeOAgXgBAssnGQ/7klXSAGyXcCXaeLUz0PlD+KUq10ukVu7M+wXvZGPPLT5YwSSfOV/QcRrij
95Kv+aNlZ/rr5pExwEnbPc3rfJErsD6lNFEday90DKYoLxdE77FaNwt6HQcIw/ROXCJu1d0YjIgj
FXoZaJffgVId+lq2Q56kC84N9xkXCspsrKKMhnKawHl4z8QE3JSr9AZEfKI6rx5adNgx18LyLpBI
J1YYsEdUEOvoiBVurvD47GkB2RTRQ8XWMcRCZSylrtXwFpvI+KKVODbeZha7Uab/IUIczdi6Xn2t
xyVH4egjRPvzGAkIFmi1Rxa5rmi5R30278xe3c+Dc8IJokIGLF4WR0qrmIISK55PU9AKi90V7BSe
WoH4MgTEiApFueEeT7752eSmKgxigX9YdXxjSP8Vrcr9XetKCJuCiIuqoVQMyuzpoW1tvbUMt+tP
ZvQYv8A8PHVGYaj9sCpQR5MtQOr4/ItKzny5TIR416na+Oq+NyVTbnasEkBGA/pS5jpB00KJHQvv
9DYYXBkg+lCljBiCw9g7U149jA0Eo45/RWnirEd84NBqnq64qd+TW1A1/tQzczfA6q4DesDp6646
eBN3PTwk04vs66a1bbE4tcmS0IuPF4MHOea2bi7BA+l1+WUcGcrWIWHPQgm1cvYxC+TKdsaZe/W8
sd/VOf1a9fiIxG8lJLCOTwBo9nB6Hq9+L5IRbyWT722ZvaeLDpJcUvk4HXMU34x6g7c7XTcl5NX9
fK48uAzdcvbwujUoQ8SFmYfB7lpeLIdM2xV5Jau08BNc7aDo9A7vhE9WASkCmz2yZP49oW0IOEPH
BTISpTcC2EBY1SYMUX/9dlAQRSEA0/1LJfZzBVi/XqtkTchJoQ8qM3sjyST1ltiqV6hChyrNRP9K
ay1kiCuBvRK1yJLbesas+byIaohYzafedxV8rvr+0v8i96N6JVpR+PGGB5IcP0pqL0mnrObxjCYC
azSDrtljcOK7IuBjoTZT+Li1XOpzXhdCq90KXiT6FcfYN+gbo9i/kfIo6kLod+rcW00wPh0DbSRI
aa16409fnIw56TDntQ1DjGxB7/lcW6Bt6SAMAqCYgte7YZXeI9HHvmqChX/mLIkqAuEril/Z4Ra+
hIut3WDmiuhCCd+MxIKadqUl6r3n+23qv7bj/32REPZ4KzamXNeuaP12kBEIYEkcZuKtyLCk6zP5
/EsHlmnXMtJKoNNZbrp+/Z3m8bdjQivUl2MMjnZKzSvoWmuYoRiYOHVFe4L4T7tQlSupmooh/d58
gcZ8+ek1IF+ikfG2N9CHRb6HQ61xfBO1bI7ss9aCfx6yzUg+Y2vUaA7mSBLcwPNyL//3LDVTTh6n
bxGaGjndBoZX9dp62YNSYpRelZNAm6tcw6hVuIJNxI3P128bRDqcsc08nB/U3/l5XO7EAyjefSUM
QtjHkZ9JNytRXohISwIK0ypWslSHkXI466ifoOz4N1ZEyUkMgaxxvBG+C4a8L9N9/IQN7AjmFqGa
VFgciqEc55v/oqmpnk/lZ/Fuzkeqpec19RoQOHbzm1xoBp/j908KQSfZzkMwzmBGgaug478fCDMK
pWwTpIFt/P8bUjOaNpfz6MlHD4s31apFp05LN2dh4hbwj9noGB822JJ0vq1Bv0RHhaHND/On7bXg
fRltu091qLowD6k0NySzBkKHrRif8IxDmWWEOAvaU2QK6yev64fCPRZ8fBDzaYezfSotaSLFvPlg
UqHXa6l5EjiCLtLCcmgoS5EGs8T3pMP+hX7iPHMDn+ZHqwyIamuZ2NJmpH3SDH9uqIj5brWxApva
9X7keT31pb12g5RVJB3O4vyIDQFKyule6qB+soyLmbE464V9k6+JoL3Efl/RIF28uUXlN3nV6rrc
nr2lML+oALgDZTx4WvvF6BDzfUV39XhQiCjzraPKmjSrV968uqqQH+zQ3yfmwbi6ksdt+R5AFqAe
togpA34h7a5ExoIk/rV80pUcaXuFGZh5CBJa+nt8xdiEgA/bnT16XvKwWDpBT1oY08XJKP6lk0Jr
2+SLbyg2mMm4Mhz2FxXVHr2P9rBtzxsQEmJG+h5JlIritV0Dud/VkVctFhGq3jr5mRl3wL71SFt8
tM4zJE/lKj1qPCzY57An8Es620OKsASQAIKTA7HnM8yltuknM1kBSSM4J7ZbcO8XVvZu5tO6Hys3
HX9HmhIePs/p6xGPMIiHhZrlB2ZnlIRUt5Or/RpwRIwQ425z4/oMZrMvUexw9iVgUB2UbPZVx4QH
uuiyWKtL8QEoNcuFLeOEQ6n3prvaO54Rsc+FVIq90ZqaHf5i8oOLp5DHfljE/PJyprCYNNAgJvdI
Q8tHt1zzXpTMXnnjFSCTuhrSDQUIKA7kZYfY00CpCXiDk0uIDz/XkblQO6QCxy6RX3lj1dck3F6H
NMqBaws9fTe6JWB6FTOeTHzyzzjplUsZ70ZrXQib2E5Pc792Cr7wBCr2wzaBdj1Og6bwpludhsFl
7/p3T4dwRVbaSNxO//vJnGmr/GZuSzPt1A/sOpUTPKByiGqhLnh4Ynr4u0o3bAEo1FHrkZu/FXmp
ALjh6hcFEqZpNLdM0nmSi94uvNmOFZah7hLigqGPifdDbTb4z5rgB08vhnMzgnv90KqDqs+anzQv
X+NHRWXP44SlQp5V6lZeW1wbhwEOgv7s8jOioLx70GWjihPtyzzss9r9eDvIAxJD8F1s6jHwj9ne
gWrqjWAl+af4MTlFUPbmkyR82zyEjG2vX4Tt6zrjkhILIcijhVrFGd2zCyiFiYgskExJ0x3kkY/p
jrCZMhM75LbFwMXR5RvlsMH/NM+SODJATPnHZkhQvGvNYA/3NlJ9qhIzQf0nTf5rZ66jkr+vRIqJ
tsJwrl6HoK6EI7x3HLKapQvhPbqqh4IMJjRCBMF9pB6KwODVYVFgpG8ZFKPzJZH+C0pFHXFBhuOw
JltXCALtFC0xObrJNWHV48YsMs1MDsQ+/gB+Al32h1zMcONe4oR//FPR8BGDopovH/4OvRF+ih4c
rSnSQ/ql36leJcJFIZ8zwGfl0oABFkzrdTI9+Li1Lcp4l30oV3j7D3VZ020K1YJEQr+ri/a1XnUy
vswgwdh6StWnkYFaGEk736+HVpduf/1xke6GHZQJXMCTr9AAC+xsnppLCtJVYzO9UwXBAU23Zui+
613lopMGdB33hIeB796Yd16lKqBuXFCqT3tqKpj4cvII3RC9x/tVD07VotcvLNgaWNl9eDMLZbOu
Bb9sMbeGxI6ujX5ektH+22mneTzBksmYK0oAXAkT5J88Ifri5jMWGJbFZcgppVZea513c6Y6ftFf
JsXzni+RKM0a36blLptW93W//EfJ8TWzvzJXiCdr8bKeaRszWr7o/ZaSsFmMHNDGSi+5KxHIpSul
L1/CMBX04qPBvFvWNBuVWYZ7JcA+K5yPYl1F87/PWgQHQPj78rtpUtVklPLvHi2LnYzFzOyvmGgx
qb30dLDEkJLY63rKw9K2s9m6DdQy5CEFLVMoZh9VjEFYXV+EKitIaUEP2Zbll3QFeX9uEL4306v0
A6g9IpT+/n6HHCxRRpZ2UeVPND42MLskP7PHQHC75LEzblW2TtSLv8ljts5J/Rhy7OI9KTJYcrr0
cpxN5W44cqrEkK+dbPeieH4X1DdenZ5rTho9er071A0AQD5V1TBXzLV3TNXkiivET3d1Or4scfvp
XAkYIN/9u/fia/pOdPlBBK6v6ZMxsNNu705/L/DYo4LgvYC6nP7AaCfqYrT0tDpgENPfSbq2mBJK
XX3CxqKkA6j4/oVS/01FjqmoYXoPVYu0ajOedvevTpqaaClwJ5XamdOzHSQ21jRWrM7QZEdO6W/+
ovjs9kz+hySAZu7nEQQTQsKAKQO02AlPlZ3yxgmQFwqlSX+oPrsZefMb+79elxFr4gyvyjB4tH71
OslBmJZFXltWRX0KsuHIHbdV/a0d0epAm7gFpRt+Yi8N7Y9g7N17Bc7vqF4fZlIkaHd9FyZeyO9K
764FWuhcjzHBiyHa4AYnRs4+GVSACSbl+/jftNWkDau3/ybaorgFfmhgLB/rdkNUYEkDim2qS9uN
pfxC/vnUlZTR5iyNbWRh8J8iWl+gTGEgtkBWYWFWkk7aTobx0Xx/rhHB08rAu4HcujR1HdoHbLOq
O0ZOaV0EC/n/MuyiK/rnkQVLZzQbMqNZ90IkSJUJLjTInlUIPVdPBj/7vNvNjUnFHY2x1I3cmu4X
ABPEBPPouNSLP/W1+zAvSkxthnU9q3YpZ3GWtY9VqOjXh52frIuMqVgVFq/LPLeTPF4tlHWoGMlW
djc9ri9lqpxnp/BlsAIuU3Uku5w/jvexKox7OPFSFayL1y/khU9xzUHlxwff/gYCYn0LrwZVxhbB
KbYng3Ud1XyGQ//ATp34rmmZv+vylD2tfjudnyucIyrWhsjRHDW1PqMoo/FeYU0JcUQbLzXcZpfr
+1WZA5EqRlaaCBgrargfpPbNWJE1pmfJ/M+63hOx1YQfbzvnbd+ruNvN/jania5fARCUCZ1H4gGJ
JfQ2E+sW5GW+shD6rLMf5CgE/8Y3DHGbe1BU7Ughzzf9/cd7aV9sGaYThTEFD1+YH/xy/LsZQ0+k
L2x7xowdwqlzLdRacMTk/upDzPv/T0slHcETYDmaZMecz/yyiybi7eKpKL6zifeAVu/HT8spC+z1
0f1rpVATQJuRMecD1CynlUxkkmU7on7pk44j+M/DidLTcMVmFK3jAeEBLKh+UsLx2pm0Uvv03SHz
gGABDaKD/IPHnxcm04iSWF7fDYuRTpIXivsKE6/le66wm/XiOCY+OA3qABfJNthRrQQraPoZ+9oB
kjN81j/cH0ZH3KRE88MG6GZQN/wA0KQ2/LGTZn1y4yeE0m5mtk0rN4b6CDrgI2d/NrQxqhH/xA7S
3RP9nw0aH5QnVceKPZrSTsEhB984bYxQz5+39CRIUme5CeP5hhPlls7JoHnBynDz1l0x4zGVnCoC
eXdIR3vHJnTzeaUNGr49NkKhdI+AVRURwrbNmZIWxqkhHg7FCH/6v1MS/8hX9b8odS/UYCqGxJzE
ywNcy0IR9TCS2WV0uYDbUvlzR56tx9dNv42Nivg6P/np2pOieE+I/KFM+zaiO+keJTBiLruLeXws
NbF0IDJhDZ/z+svs82pLOz4u7Ur2y0wDA9R0SCDi7t4hH20A1WRak4Em4Y4Kmz6VQC8bYUS6qkZL
Xb2V3UBGw83c/vFONvgrQD2B6k3tK6cfwlcvvWhBZsmTIc3E0ZyZJoc1uEsI7wSW3p5NS+KM+c/i
GD/10cEVom8n4E/RrsxO3QKXWwjwV94iNR2bssDzhd+CzD5TiTTKYYnTQ3Zw92d2EDQvCBGDNZmA
UDuFbkLN1pA+Wun7dcIs8aIq2fZ8YPJrS24Zym0E/oaWf8FfmGoOTQsOL8Y9o5n956nmtlZkRzfc
d2hRZ6sp3Mw9vVBDfWaIVrajH7CzG6Pes0ZV4eIHTRBKj2LoE0HpJ6jxkNsDkJov+O9it5pffVuc
OAdI7ea3LRWN4tI3wWra8XQHTLo4gsn45fmnqHyilwwjdEpIw3wbCISeg0aScjMHVH1+ew/XKIlX
WLANZb9Csv5Qi1Ne6BmrUquXedcjGDcyUQoKD8ji1ut82Y1HcF+gPSqVXgfMpQ5RnYU9A6bWUbEt
952Tps0xRik3LlHAhXY7AVWR5gnDMyu0qrQyWH4h1rh4tdEmTyGrYy9ea20azrp1dfIRfQoYDOph
ZSY66cX+VChbJIriJzw1vBbAC0fPcYDX/xFbbfBw4WfN7cAB7w/GKLR+knMBJpYIoQMEb4HF2aTb
m6zN/XoF5OwJdvdelbwNhT5laq8l2wWv7tKCpDjTMRb5pzCTpMg1oIPZLXlKAGJw3gTdOt9IAaYj
vN8QjOhZMKwjc+EsM0mxi5F/OO8Lz2kDbgqjE6REbmiSutChUvj6e3PKnFi4XborXKIRtvg1n9N0
MAUQg5lOxFo30x4cQZ73nFQcYsc4tMqsp9nGnRJSZXRcQmm6HOSD2aVIeq7hhTX8Mc0PWdEZ9Y6o
lr2dzWZwNtvdtzl4pr8ebq3JX+LPT72yd1PiWvdKiBizGPVF1fICaO737DnjO8Y1t+YmioyfijSg
UofpYJwzu4HNT38o1dhDqHQYRqE3dpZHfAxB4+jEpiMnFp6jMqs66xLmIFupI4ZnTiVFM5/VmydU
eF48GRCfy9IvftyWgmOlUP8JCYKwoV/x0LJaBhnqy/8BLAmTEXeBtltonbnT+yqdPNFrY1w98H/i
tozdwAr23EIWzWEMN7koIbLx7iUH81vw5/lIL3j+CF3B+p8mHI7WcVIkkYzv/nPpPmU+vsZYSoUr
SnI9mxa4eDgDuabsU0jvtM3QIGFZBQwrdp3nr7mXLSHVhfcaInClpjeTTSBBy3VkNa5J1GaE/IoL
2/O3bmZJhDn/b2UiGZIIZyAYY3P9/LsSxQWXBp87LnAMpFQf4/wdRywkaODNdwl9SkBIDP6CVlNA
oG91KO+IoEobKTi3T2qO195kjjlTnpo923JhJpaXvY5AooTRC6ImPqPst0+k7HIMtSUdri1/Zebn
MBXawNBxorKjwM4z0RdvJBVYCOuchQ/3P6CfPEfi4xaQsc4dNhjOXZoSkrLiNKRhnqf2f4BkEHbY
1rU8/RXc2UAbriokEeFLV6vakcpivwTq/at4E2m/Pb3/6/GxoOF98+XNl21M9rDZhT5rLo1TJUN0
IrmK09LKKgYKqZHC3BMztWWwrO+sN58OEmhfKFbGp0vGQX17Op1QDqs6Z6MMUebaZzuKFjqvVbAb
Yc52dVumg5P7ZnsnwXr6SDtbsh5LK6nvXRWjyvoOYP/XQftQ9or74l6Ltl7HlyY+jr07E48gdYNA
Djfyydq12SWv+T9VWPN3CvISYP5Gnt/0uOgh7SNYN7ypm07U/Tmj04Uxosc0ZXLF7lbYtDBVUhr7
wptuELoFQAcNKcPWbt48kIzS33n89u13nkiNvOHWQjDKgYDpVRoNXjX1khh+IvT75DmkXbxEssrj
THQE2iGVe83uzy7QVGJo6cPAt5Qv1G+ldaX5k4/2/8IcfxCHbkAwmNF25DcG4EsnfeCNAj2Oigmh
ja65wKnkiBJQ/13kpO4mk4QIabswiGNIhHdQV2sd4Kub20Ap0vwg+mgo4zRiZ7Pex0ybz/WSGkGR
LXZfWeVBNbOdRf0HvCVbAYHndyX/IeDnSmptk8D5jzFuGPl5bdPlYEmNN4O0SU079AnCJyu4BiCy
k7TLSYU9kWmVsi3sfnR03WdqsiFfGhIKfxrT3c38hM8udpqL+lfxNbjt8ZOEVHEk9HtHttxubCGz
N6WZCeOJxSRDErj5D6YDi40jDABgJGeTRVSwOizIBvfOWUV9Lr8mAGBdjNH4yXNBs/+xIsAw2qE3
TpGJP+foLp0rGqPQnaBQWPOJ+ifu7JTJrQFUDCQ6nO3PU9SHL4wLVTurEQGFg4rFeNY8pdY3j4nv
K6+y8MzBsDZuGtbrsqnAS1uj7gV9OMa5DPIssCH2w8cwlEqLgq3LP4GelN3GvVitGagQFBahNuVq
bt8/9Kx1ngTYn30n3dkUqypEQdrAn/1MPHGAZIUjKMznjt/jUiV6ovUuwbaVv+4sicMV53qp5HGi
9BI9UItQJTO34HceuSrW3N13Vnmq6qnJOlWg5vhvbQUyGy55SCafxZCroU4w8j2+vbHqwUTcSmfq
/bXWocNtHQDFPBTpH/5xsS/f+89NPlo7ZUCc17Nvh3J91uxuTdmI0C4dOKnrNyT3pf9VtDamWYUN
VIAn1QSA4Hy0vVvobqc6ts/Yz2QnGCnQVcRziEA7vsQcAfKKda+DUy6nuuVP95T6kfiNBjk//W57
8aCnCp/wYSmg1kqjd5GAZtTDPT8kQ9cdA1vZ9MSPDRPi2/ucBju9WDuXJBDUF+pt6gfmfr1XWwjL
ydnxAL3IxD09XP3Sx8LRFzygXGxWUSc/kRPmO8ahJCl8VCfjZScft4lf905bk3HhgDBvAWaLneaV
ZJvyauKHRioGauXbihnC4S0YcBzVzi35mSwsGLHjudkqJRl4F7lnQ74W1PIdPRHzhSM7IuKpF7+X
hwD+S702sOWVLEqkffgkgkSwqqkGixNdimLY2AMjxjiOKwciNW4Mwxe71S5zQqgn3u/O5SzSQGSR
eQd0hKzAl7ORMi4o5te21SzgNXB2civU81QSoUbX/OyRl1JocXPGy/tg/iwPPL+a34RMP/h19Swp
nGGj2jKY4h1It5lFHc/lasURLIdy47cBoQi2vSzuv1kwlrt4hKm9H5VH+KTDC2L04pJvPiuF77/P
6fVJyd92RcKlM4QGLDx83oEbv9aeNOzGeAoPr/abgRJCG44vBqxVL8NT0JCwOuXi2ycOsM1oESeE
eZPqemcpYY0vH8I/dioz+pnN7tv+DV+Y3f0JHgwi3dUVr4q2ji1G+Yo0SZ4vX0WDtQt5DPMBIDhJ
MWfHgS/CzePPe+04upFBETxPMDW5iIwuEc7QUdfVsSYdC9Lb8KkeBRsBCGFTsTz1GjSsaafECzHc
4uPXWSzdY41AqIA16zFCyIb8H5mdpEKN2L+0fYvaIEKuGgPZTafbLaxihJ8IlLdM+S1jQsGnRaoO
oGvpdDLeZ1q5SnbSqf17sV8V4+4AJ9N5hB9JgTu9Fhhws8BsD1Ecp1ahTxc2roXvscg/MnIYYqcm
ARValFicFLT+eNWYtCPBP8adQIB4QHiFlNZ1O4ILT3NXjmJNy+dz4DonllajBgHxlJ+3eLxBOcHW
874vIzMaSBcQDXTkiAbTV6UYK2qEedO34DrdXDVLLfPJ7iQYHis4cqFLFXAAio3Q3fMCywT07jJf
2nxJD9BCl02jAsO4XpWNyxsWgZ1fFXKoUNFw1ydks+4BGPH+Uhj9Vz/o6w80QOjWC7dDqNbzRu7D
PSCKpXZ/eZbYYEHmao2Aw+LpHJ6LKlmHUMbIS0k/mXxIbO3HRVw1mYGzxUItfU/QxDu0UqBpvNvN
xsP/XKtbIi055JyVeqEo/mHwA66OL4tWSqMDNCtZDd58LdjpP1u/OGC0eNVCMKW2mLYmWqg9HBxC
M+avscklIeQKv9ZT9n0V+Vbi/Za4eKVekkDGkSI/G77dDa07uRp4nohyrSYE6CIhSyXsNLecz7fl
eo5UzC7w1d9mO82hQQUx2IvddYfEwQKwJbxKxdVIX9qLLqS3XeK7ZFrXbP3ZA2kckTB9+521srNC
hQ/e7PFhDkD+b3aTFKQns3taDZySzrYhIyAYnkr0Ay1DinwkvERgHrwk534m7lTm+ws8raSuhrbH
iI/7+Q8KVJ+NYeuFKzvZ8G+ek1BUjAAHMlm/GU4pSvR2gyI21enTaL79pJuKaqMuoBOHjOs6jeKa
AKNg8e1dTCS+KrCepejz9kIAeGjtFk6WflUeFZBrsAXKh4QstSvpObX4eKpOunrGAT4uhTpOni8w
QmBulx9IjIRRkr6tR4VOvVzTJl/x+87XeeTR0bNnMa0znkwGjlsiXjmr/BsweiO1l1r/jSOC801r
DlE/ZJvG27alUlbukHpMxR9ps3tgvFsyIOUdLqGeO8FtBFXVSZbWdpGu73FF9yV/01n17zAUcPDR
yWnQh0w4m0Fmb9S8h3twE9DwMeRA4RPL5rvIfCpldMQbzqq8r6cFVn1YRmq6BqwWXWoJHMoFBX0z
Ht37phOWhBonFhUMSrk0Z24yk3sGOSttS3+i3BfMeZv0gawbpoRDYtf+JsISwWTkyHO2YyiGm0TM
G/Im4f63mdiP3pd4nBSjGvWwTAQdFcuq8swxPhCA/EjFl43jBoIQZO3luo3e7PdB0X2sodxP0YGe
jf+VHvmdV1aLDR4GBf+GbHlsCRdbDFCiZ4dB84qWl7r0qFKvV6aBZzr05Ip65tU8wr1Wi6VLHmmg
8lKrzIirhdbgpO0wvw3MKDPYHUb5eXp1HtAnCRp3qyuWB7RgPi0YsE3VcgPPB8oFfdLQYgR5t83o
Ri9J8JLyt67S0qh9ogLexdiU44r1s4gJeWrvoPwqpHvHjVtyJo1zchgU4PADZaSTGgQv8MTpuyHK
9NR1uIuygrqUdUp1cG2SK8JL+tKR4H5iGD2yh+3Rc/I9S1wREGPA0RAlHaEajXUrFWmw8le03N+0
GOQC0ozA4mgdDkKkExvAwKMsqoRDAQszOrtbm6rbyqDI8oR1NJEotaJHM1IJp6KPvVZjOolwx81Z
NxFnnRLf3eT/U0PvwXEbxXrA7TgI2g5fG145ib59CX3Wl69NnPjrU2o8IyASlfgw/L3jOx092ap3
Plg2qSx5J3htGLKTEuZtjodfmNMW2+0M2X05gvkoiw0uI/L33ePbGlVTCuJXpuVD4dd5IXDxhMUg
bj5d4MRpzvK8qJSGDZsyrd/0Em/JSPOW3L0U/GGVcJM6fDfl0++9PI4lnSo2ZZq52QJaAib1aYMG
n9cM0pjGEfTdY5HzkTosT0G64Of8lqHFvlBm3w5HSeh5D2WHVdpdImTOO8cZCMxkIKLqpSoDr12g
pmcljxAlbXAvFvzT+7JrRPFCBITjBbLXS10CtlftCBlZ+5SsKWFwt1nDF7Aej1QzSTnI9ASFcMEO
oDLPr90p8+joBM6DXDg+Nl2l3Gv7Zo+eyxjOTtRTWxPOIFXbQfZlsPytYjlN2d3UFxHMXIJ28kJ0
qspqpw2/gqUhsZLM0a6PXAVpnaxItIRjFe4zmlDMfHbIuWp63hiql3YBLi9OWDSEDRkT/NvC5xB8
M35lZOiQQixB1I+yOWeAwLK4WleAgM5dZ/8GjcyfSDcpeAQQ5CSjPSHV04qbMc5pRJ0awsRkmIys
PPeRDuelnL0Ubhe+wb7szHglADHOLJlXwGFncPtNCnwF0tE04cGXEY4D0X4qTacx5ubVP1fwYwuF
RexeWQaX3hOokFWfgvK487TOm5FL9j6uFx4NKE0W7OKK7lcOexdC3aS1gU/UxZ7TQ0yu8em0cJtb
DP99LnUzP7+FQ4sqGNkx+U/MqFF+LRI9ZsnoaWBrnfuBDgnV/cr6hkCiOBcc7bSgBqOshrviGO+p
Nx+8ALqz9cM/YvjPSi5s3uU0NxnvWPgIPzIsMbhWAtwqKch2MnUNuLEIRFsoMcqJ6XVStUmDdAo2
yyOqszkd0/HKAAPQ2zmRoBsWaIL7otQsujQQKoUjDdYsPqWu88xfS+TNesL+CDbPwykY5RdFVwg9
mafb/5ZlhAM3GC4Ra4PsPosGbNdCmMrY5crZSDLMSzWk5xKnXGqYCti14bcFP4q1vgTPngGBWb4c
qyt9KM2zjLqDTMgk13rBxEviDesHOtS4Y1i2vBhK+AEUIcjB4I9muV+U7x0qew4zdMUqplBnEvoI
Lx948ywV6nVQfqGsxTSWy2youErPt558Dcrrm4QSfUvrAVDyS++Bvx48qJMJSqzB0xKH31tyU1KF
TL946GBe1eOUCGL8axAHu7sEEzXT7LlEmpkIefocI/s/N6Ww0uXg1cop5iCyTuFcCreSv9FXD2ll
nQnSPpixQVDi04POXojbapU0Ckal1XYEz10l5G0RxBcPtmOJ9X8I5kvytfJd6rH6MUig+1jyoltX
Av/25jh3gAz6PpfopPJI4LUasoFb3waFynDaghrXEOxXigxgLO2qLWCYgjo5NdjHf3xiyho5CY0M
wx5UlcVWf5mUpTRpr1DYcmHATOmuKz8tLlmVjQ9NdSneVFwBbTFDCtqhLp5CU8+55c9pSz/lVUhe
o0njeurL+Dbmr8JS1pexJ/XbsuTT+apVcDUBxVwb4AdHSL9lrxD7LKPx+iXdQzWjpI+HE1rhm9vX
Ua76PGTd0xAWBmaSY1wPjdLD1hpc9RCKMHoGV2uHa+iOpYXtWKYFWYC3HXIBjf44duVOfpQFBN/v
dzhAoM3DMMzG9Xon6ZOZpt3A/KtiB6cgZ4wTRMORpAAmR6AVZ3A1+dj3VltSwXPxHVsS+hg2z4Vj
U2xcSBv9N0x3pLJtXHw1zdOvyppl3Si/Sg/HDFsHc3xahmeGR9ss68H60tS33W2i3apgRIZl9Fif
s0BhDtGJ3akdj3MtNr7s+AIYN821crJe30h79hhmwfnWBcn+waZ4aSq6qnzlsGotz736PtQ23fdz
69C0BJPaubCgfwz4zRKVXfK8wQgf6H0ZVJCXHUrLQJR41xiU5/6IBUfFDFd6myYTD95FnRKNi15Z
jxBTs+FWqcGSNeM8jO3mrfz2tjFvC5CgIOZxFRlY56879vwsER6AT4Je5F+WIWOtyrN70Qrna8bB
f4wUFZKVw5EO9DxGxHa15r35LPXolXrOLl22/z7B7lXTC0+6EPA6ThuCve0CyiRlu1DGy6XzFX0y
L5XNd2hA9qEwPBarDdyxyHbPscLcrBRgLEFmCjZtcSfO/iKxhJSih2KJMz6ObS5pM0CfBULVmGtd
7KFOU3VHIqGNMuFIJzwV9UIIOHGXJeG3AaLTwhL0XEOY+1+rIGkinMYOz+fxht7xjPKlYfMRAm06
2qZs6Z66BDhqngrsb1J6BwieqfnTwr/+46sii9CvBNzrgffTZt9z45vJI2p3a8Sw/YLTAzap+/jf
lEZrNSwiIa1brI8/d+GgnJ4HN8NWqzwqZo4lAORu8rqncpkJtkQDnXJW476PMvyJnbkUZrVIGVxE
dEMmUH8JJgmMwldD5+UBxqW9EsDdB1I0FvHFXC7uZW1o2xFfuCi9Y2yQNJ+hlmE/5WvijDONTQcH
UnhbwvbPNMjS7bC8zeyDGF5ojmKDZeSfdhh7e4aHRmLnLIC4pc0+vPJr+AV0qik1r/UNCnFrsnan
yBsGbKoWY1GiZBGmIuV8um2UXBOKEns0B1NNIpNzir4bmddkL5IG86HvI/jUsqAxExwEuGpNBjSn
MwWYhdHcevtXrPUESJ34V31da7nnK+6hoeQky65GCTvIeGknzJRU9jg9Vj3DCSB5wwfxqjE2ZCOT
EvuefRG5bYZvfNRZndWgm1fZSnMNF+vGO5JXlxLNTUPKVbvNiXZTEreJpkQEt/NKJsnzOMcO6Lq5
3c4hIMAMgFjVLmu1rFNvC3oxrpFSQfX71SV0u5Wh0+FLsz8/1rwUIQxE7G/9pfB3b84cXgdH6Chh
Ca2ITdMBhk7hPIiEiGNPswy5R8+fgkgL4d0n6A05z9APR3v23x2c8MzZCHtCLgSI7KgtXq1LqGnl
luWbO5p5scrE2rj4sdRgfhwPsbahegym101kSyrhz60ruUjFOxVZ9gu3RKUhU7eitUHPn2TzC4r6
3kvddbceT7l6SEnJTOCJ+x4e4uNCG4cNc66Hdd/rvlNqdUYE17qm8uwsc/hIJzvgbDFBnJVAr4sL
Mdt1NQyUI7rf5XgCREPIL22MJQtOQnXcepdcy/j97u43JPM7FX7HRNmrp7ZpbkGEZafgzIFCNXGi
A9TkRGo03YXjzVWbF8vWc4FtyWdX7Zi29qrpMYoNqwszgKY9fG+Y+dPpE5zzo2wimM7kJR8go2qj
2kWUoUzh/WdgbkvM+K/BJ80JmV7cnVfv4kUvYpjwSeMV2CUm7mQXlujCGSsLg9VQDtrZQPGZGbTx
C8OXZnYEW9Ms7bdgi9Ax891NACJ5wNUIppDPRFOcD9zuGXyUQWIxr+0vvUcUsL3iWPJ2zKkGl+2G
OFkFEvsFrbpD6T7XBOrHAStL3kXTCW5y6tFGm9+k7Tphutoc5F56Ofrzmxiz930IyzI3Z+AAogn8
I5wKfv5HE8H/ecJ/P7wUHOetkxw8ZMIj5HsCR7ai8GbWnB3mcVuxs+xglMI/iSElMedcFJU6vR5z
zXAQ+ZFHeLTTdDd82faY8r+ZGrkLq7x8KncK6tcdbgVXigvzwhqceru2QsrTUB7EIJZy+CCHwnoY
zV+PMGX8wjvsGgnFGPIKTUJrPcvqnBvGPp7YbM9L8fEGYPmLyddehTRJEN13dVwgCtKn9xax9yx0
ekl5BJH5vMzNooYDEqPoP18cqReahIw+aeGOxk9k7ajKydYGe6mRFc/eN2P8IHLd/P2EQkOpr0R2
3MrDBZUQTpiuohOY5xe6Ibqz09Sz22zQQInx+3mxR4xcp/g8IsuIf+7Sq7W+irFJM5G+Zw1eWZGr
DTtDC4W1CsVAz754UPcZhppTGiAl5Fe73HXYzlX+gFw8aPL3a7b0Wf++AnnbJiwB4on22zzNuFHS
alVnZ0zMOiHjtEx2YCpmOtFWI72HFxihIvmfuPJ3EDefzgBJw/BVIqWyG5+Q+1AFe13R8Dw5QlvP
4sKz8FP6F1tzxn8a376RZinfKHKARzyxWiM5xvo0z/Yb9hLc5OEseVo4Ej1IaTjbgumiuFpY8+NH
hObO1Dmq1cqMqVzLFedD7UmJYB8gxAdsNrljVybkKzfHqqfBRPPrUOJa+e4roPIX6OsariCuaACD
0gGwI2Wxtz2BiNSW7HC0iu1sQ5L5YXGN6aW0U/AN29b3A/duXEjMOj+miOUXwhSR4ec0B90hFcGc
F/yRQFKoOznaI9i99JV/s9GQgcoNz4Fh7QcOW2qpCYLNOJrkz4y48smh/e2FQ2997TWgmJbZrbxb
xiIvEh0EGNgd6NxImY/CdWu4aMAGL6+ji2E41ZL6x9O8aLpmX1hmNC1uBNtvioKbTNzkrjhqtWQO
xIfPq5ar0x9GxNjcHOUx4n+JNgwpGM4uWIJ1vR/6faorqmbwfRYeQ7Fql5CpCJ6LOfFk/Sf4G4x2
Qc+Njh7nUgluA++L6UcDrqFEpRE8IE0k71QXHma6bGHNtxbvFtE1zX2R9qTO9R++XYSsS3aTUJY9
RNKBcwa7hVk+BrVsLFO1P7OcmKYFQM+FXTnjDIs5PGQf8q8hXEISO8+eIty6yjHrJiUphUOe+aN3
w/xfqwPkLgsxt/as0C41McV5V3Ve+lO7Nftvb6G8j+WAUb6eF2WtCRtIk1qxfoIFqGytvvoOLlQA
6X6fag10XkbGYCc4j0XpYi+2hb81FiwWQY9PO5xsM0bL4kqN69Mzixbzb4GkN7mENaBBw5I6AFE2
4YSs9SxlIgGTHh26+9F0F/cHISdLFM6wDxiwp4Px/mYb7+6i1xBEbpoZ+GBjhjNevSEMH/Sfrcyi
vrP0O915RMcEYLCJJNnnl3aHVo4gDORqcC1RFJLWdkxdVKWhPcYJEPvkXzdapjED3GX5bBAUtGje
MDhjXuK7G+oFOpNauZ0oP6v/q7RKpKn08FFhTrEunw/RNjF4ygm0i8poq60izini2mplVXwKHf8I
Prl4iYrUbJiyTXaYOrEZxKDPR0aN/809aGVqw+lISHbVAFCucaFbCh5VnE6evC4Qt2OGSKE1+xdA
AENfOjf4pl4idBx0AjnOO2bKzNb7g2qobk1+8PA5iggVPLM4bwcHHT80Kpp0Y3n3j+sjlRP2ylbL
vwAAVTQcLsDYmQEvDxbLhKtSQTGr45FAloe5uUmEYADMSvoc3TsWLNCmvp64H1gZwv8srgWZJPDQ
zo5bgpCixNLkQK3TgyXF5DL6baBWUAYKt/jypl4tM2p4LW5Qhxne8rmVvjVHkZvBPwx7FwVAOGDx
icgOmk5jI9eTeX1F3g1UYbE6Q8EXtRCLxMY5hX84Du+oXuTwqdzedxEez6gmV1vLLl6+9DzNBtM+
TWCCVbf7CReeMMvjOkdM+27zYwrTbWy1AmQJ6vTNulTzNN9y3m59lZStcWv3zy4SinVJjmZujAyZ
iuqm4NO3ey/tVnSvvyBRR8fMr07VuOdHO+Kq//5PUao3FQ/IoapICqDCTzHQMNEr/H1VPrH7556w
YpCr4OUR8kX/QsoTraj3fAJlvF6UXwakHEhWv7sHNnZMVMCzWXbtC+QIRQINCDGfbPXGGNDD1gxL
ajNAvMd6pv3JjQNLSm5njInaO3jcdcxz0pMcC93RW6x2xfA8YwHnnldGZpc6Tf1JvUgDOiAIkrCZ
e0nafey9IDgcEP+WSetpUox2YXoj4EjSm5qT9ejxNLDEcozCeelJmkpkTLfFa1ex63nvkaNFP4JE
ZeQ9txrkMTOQadZHTaoqX+WWmsNa+o0j2PnlCFwRW/7IKy38JzAtv8zzgfYnZMT0+2AzDwd903la
TSs5+T4u7pSaB1F1bCxZjddWYjAN63ec3YzOr7g52ajHepNxT3Ir1/R30YwLr1CMJ13hGdi6QRWC
rWONWkJlIWJkEKsZNmSIGLvD58uCW+JmYS9rKfevG8ueu620+P5YmxMcfFVN108YTZAYW4egoEkv
3IRn1n7fkthSnERL3lvMGvrCV0wHtCUr5JFR2TLFFPB7QtIW1T1VXKaPDFrwOOAaAFtYGMUYvujY
5dxFRpNPNrIsD2mtPTH6cBFpBksZE9RwhbNlRY7bBfE9gsNW9OxjsOvCQsFzmwc/oecp3AnDEjc3
+BUcDzzc1RdmNn3/TXiGnYwVI75TB53pdLxLz1EVxTxZ6oJzgn/ZJwrqsb9HR1CwNtVw9VAqgbM0
B3h4jpruKIYpc+YhMHJAVbqu9ZcyOUGk/sylth9lJtI8GaDP7Wkmw/wlAfiqZvMpMmg3kGtDDy2y
6/bbfa6Y6eafW3sXfurrPfghtu02M2ACn1O5wP4JfVovMDGBJKnAh+/99eh6UMXFFCWEeQwzwbj8
25Tmnh4eJ0QS8LxHbPU82+ATWOQ8Ad8OM+OWpYSGX64sneyWdJMBZ6PcuOB1PaEMyFg5/hr4dag+
4jUdK4BzYvhWc6SvWUf9Lg5uX18f+JPrn06n+Sqj/tw9nzjSprGhXJnaOfj8ISAFWqspmy/yNc1X
Y6ridd+2Q+/mWMVw1g8zierjrqZiOjsyXM8W4LgrIqa0BJ46KyAo8f2u7thfiwdJB27VXLz30t/k
9omtUyS/GPxXDl5CDcCaSO2zuaM1CkzunDb23kNb3fHdYLL4ddUaIWI2SgXDFC76IQgUo9flFphC
4m/R6NcuTyov12JrLmsBgJYKEOwyfVl35oPKor5+IRn0HPOIcaiFc1gXBbdg7zmg31ePX0nkTmLe
sA4pn3q+8kquxBS15jR3BvLFL9ORpLNBC0jK2DI6cKKFrlHD/8vqYK0idoOuX6gXB5CNVBauEGWS
RtOlCDtUGE+zz7rewlPn1Y4+aNNcye3hqxR1yUcOwfWv/bHaQmoNbuNvyAYOWNWa2+ngB21MbVSy
YlJ0yqPj/XZzTInwZjb9FJa5BfHYeQDRQEO+OirkysyEE7kSpRqtORg+nWnjzOFbgVC77IH6N5Fb
KJsOrwzV5vJqtJO/gWgS617sx+WjUKILyDAYuM6bX1OVSZNYJv+rJheBFsQgVWNB6Y0g3mNYvqAM
qff0kZIgMKYfS8ZuXi0DrKWlqHoSnzbF/gNi4Hq+F+dnwOKGE+W0HKx/aajd+yahOVbNbKXRcxrm
rcWUETb8oHlo11k9oBkFtiMyrP+pPC5XBsMeKLXqWEOZSlcW/B6bMgVxVVG73XILWPdVYA5REa6O
32JlCCJW6BC/wL1Dxbxoog0DdcrVwoFsCFWqcOqgSDeUF1Ns1LERrB79uqvWShe+mQQwj8FBUTI5
DyxmKodblgQDBtwHqEwQKuTqhMMcOpgCGqMFZmgBudQcUd1gKQCg7wgkXgW1GT8eWhbpIJnhcFC6
JlrGIcYQQijlpgX5oPUXYLJl/alat9FTJafO1pniciX6Dmu+UFpZtvuOj4RIY17J/MOgKRFAVHR5
shR8QLe0DyhYYhj5JB/oDW1ffmkPO4r+mrQNUsPl4YHnY1sHfg9VgRJNUZx4l+8ffDwKHIXjxI3T
Gobe3AKdAPKrgkx/9d/AdI5qjyVtPENcdmXBPgIlVgis05w+68Cd96ikmylZAHV1vDoxHgs9Pnl+
nMuJKkRbu1Ci/X9AsdJZ7/rQq1TWvWuBttcrL0ui9t0fq9JenbwB8eWJU1qlIyGnzGhmGKR58CfL
WoTJvG9vqdO+7dwiwgBMnnoIlTS3eKDD2vNuMv5QX9I+uvQQoUKtrMoLj/ybnd59uAGAP1STsPYr
bYy/WxTj+TCJy0ZOn3nd/q2zBqCosq24invuB6U9MiP0AF5jcdw1OXSTFYIs+mtmjpyoPiBy1+uk
dHa6baVb8bQwUltsSPVZkZT9BV11pXZ/L0gSmyXR7hbPGsHoViw5NQz2A/Lo89T8DReIJM++JnHX
YUO6Fod+aO6PP3F9rzHG2ybMBZYIJd4paUqeoIzckIfDoUq9XUcDek9UZk8ynHPNfCaIUYrDuJku
EtJ8GeH4tXa2ncYF8J/EIU51tqubz/za7lc4ID0wcWpU1OtnhuM7NEb9YxZJsgCNI61jgOtZVJLp
o1NWslv16Mi/gMeH1x0aahqNviFhML24+Gbzltnyds8cAJ2enFUGRiMAG3j6OR7/DpQ5s7zrh2MN
wTqtSBW3Rgl03SnDEXotG8zPCygAeJpasBJJWgVmzqsCfX4d5TuO8P5w7j0q52VakVjjHOdiFXaE
BZJ2AynKD0j94CCkbzifounA0ikNvarrQEbgMe2RvdHW4uPbFEM5Iwzs5TzRcmlppFAurHXnFa0z
mv1CTuDfLcSXGYwYSSmjO4scjTmLbbxh19VekvKUdylNZ5bKNxkU3yTgf6RNNPDgBsIg64KF55U3
IeuCQ/n10p2E2bGnOOElco//jYgJeiBVn0RmO9TbMim6dTZ2gyuBPK6HSuZlDmXYF5/C9Yy+gQnE
lTX9SaI9B9p+DS+zUY3/dDySXqaovhdxtqFgs6HCOVHV0G2YT+VL0lT5hlkb+JkC1D1CKNF9gPGO
6G+9euGRDKETgUKPbXzcbWX2L0Ab/QxVw+u5jdC7fMsI5RohilmOIP3i5tcuHHE7QlFdoQi7b46K
Py/trIaHjrtSg6LWeYMMwEZsxXGk7xAclQH1fQCHNVzy7ZPorZt1r0lMetQpN90r723jLg8ss06+
ArGQtNaG4Eixl9CbfZx2eCqVCSlDbgES+j8gWgeRBDP1tWylTkL/JPHbs6bonSEVzrtTPkc4xPPT
+/O1njOPKTqUBGigg4x2iF9gKYsas5wbj2gJy8nWgaQ4Ay0oKS02PXWy+byhlA9Ha8u4+UZqD0X5
vWdVKAMzkfSm6daz3xj7UCxeYmIoyHYyO30t7h23OSfi8So7ngoIF2GTywjmDJFUngZAilkeWE8+
MMvDinAA/Wk7hIjt3a18X4RtrHDFCDdDAgYChkGg4/vD13PA6BOY9NtBnehDc6UfU4gynlhpFyDL
C0ASG3f7IvcSiLuZf6enJAhbLpCXvyjz/yLl9FXScaLiUUw8z6394+VphZBySsl9BqPL9LORlc6B
ojiBdJieWUS84vTvNzOJAl4I0tj1BG4liHhzWE0sfXNER8ZMN/GKBh5n3+PD23uCO36eab3hGaCf
Xf50h1uWm3ueY/EUjUHYW+JNHX1dyVDtC7xt61l4g+SvmtB2GysY2ftuFC5XHcu/xMtajdK5fCmd
MHlj7QytC1xF47v5XqXLmq/q/LJYXRVsqOH0YleA+rHQ0x6L6+vYjdvkS9YIbR2BrA/K8pU+LGTX
EZhKGGLcAA+WMV+zd04GcMxrKCVtYuASQzKZPxrsSpbesIakXVRM7m3tAEj0aUFBp8hYgWTnT9Mv
tGy8L/AvTSczfJIeAquiAus93/9PMOdEp4ZEO4P+dWM0D2+zXiKAk2SNo9vZT30r8RcnSFKU2kck
qMwE7a9yPPht1mk0hV0Y7Ba3sdb2XBRqiccZsWvkk+5tHWPTR/cu1MXKYPzufmpSGWUNvaFRoXXJ
qSaJoMON0MR13cQm+qZpU+p9DE9j4PYVejjn/YovOFKaJSD7VqxBRXTlUvUKGD0KyBYtX1EUfcEj
J365hxExpq6yOMtXT681Po7WgWxm2Vk+DxI7HEfq6aEpcZEbOY8uAFY17Ya2Tx4HmGfvrizxIT1u
rpnyL+igzF4sBSRTnL9eu+bhRASvf88b0KqjnMfD3de+K+1de4DWSo94E6GwH/RohBr7ruSTUPFQ
evLAq2vACcDUsvPLbOMPGQWRFrxrnd7gndqlaTxKzRvf/NDTS8ylpbhdehPfiY1MvRMDY88PesTc
nBvyCWXAVK5VAmIYSNhLSpUFzd5xlcAvEGREDec7avCJxzKDAa56Y13PIH6piAgi2rOL1kU+mmhm
QcBILXMJBgfXO+n8AbL7ksCnuzbH+HEn/48F/qX6QyNP4PNaqmIOv/MuiIFyb8hEcgB8W3M0cMqj
A7aBdm8Fs6zpT8NxG5clsYlZ7hRbMn+umW97Iu1DxpgRY7VBtiFdU5wTQZqrRWXZ9ZI03ccEAVQk
dLha39+E/iWIKunc3hCQInKYqHKRpY79TVELSBjCn0MxpcWUnLRz7FxZTPS5Hs4YfjhI/113thUf
dtM1yWagqMop9jtwYTi1Al7lj4OOYOBSMmLkdhr7Ki5znm1nEt8BkCeSLCFY2L9wBdH0GAGC2eVZ
e1t0y3k9PZL0epu5AYYMHHjUKP8MV0xnstZXLv5ErUhGNZYos4SSfhjilH9GL0XyN4mKaDmEWVH2
3h7Cp/3fcTx2OP111cWyQjLGS9UM7xFUFCYeNlM2zfRGM4125jt3jyQ7mYXScsUrz25d8Y+ObH70
CiX12f0+sCyVZcvxX0HqeFDRNQUr5LVclrvJb32gzMTvcUwHYM2AHGGAWYW9P7GzO4h2pfN9t/hq
v/z9skNibi/0YPRNTmE24jN0K4jUzati4nm4yBHHHoZ8Z8VR6cJVv9RrQvCNuB1oEFHB0naGqMdM
YURV5NUtE8muUL4fyG+EbKNXN5jMEGeq0Of6SKy4d6ElsJXKbR1Ygaonq9if7VsvsF2EPkWpT0Ac
kjE8vHKsOWqjRMglgTOX8AndJi1W4Iq+omdQ5JlHF78N8l8CLFu0ZtAo7aT5JuKlp87Wzx5/40Xy
t1K9hre1V+E5qNHpLzXKYtGyKTmG3QYAbk4Xn/kU8ZitkAyVTt7vp4vTmaD5tvvj7Ix5kXrA/k04
XRIGKqVhq5TrBzu/xzgbeAxG2kpOSjkxrvBIvo9n/RBdHMCC+EMnsI4DIXlc56njwc3ognvDziyL
m/TpYclHMvFNCTvKmxWu8GUBZFmygrNt5CKuIECDfT/XV1AaWTHVLwg8M66pjcEqBigjmy9GjYKM
0tPaP2//z8CxCMWcroLvoI4e7eQhKhotiV421fUyaAaTaFZKDkvhh6YcbWzJFddyL+Q9elhhWm1H
wQl6e2E3E8x5bK/GCBhrMA2o0yp/Y9Jvz1JbSLSziTYUc7Dgck2dq/YzBA+pIQV/yVV0ZORtIH5G
1pzMqDgIVpoiC7dpcfYA9xWbktDHV5LHD6VChzr/7c/cRMo+ay96RuiqNI607sbJ4RssO4GvGeOo
Tacg5p6fDPiwE0Oe3VJhxhIBPKTV+b7G1gYE1DnzCzo+ye4rVuDaDr5Yoef3arnuICoZ6vBQ94CH
7lKA99r0xIUv+AwJXqVNgCE76TR6V88+Lpd8fMlL7aAfx7fxlzhFf7iSBNiuL5y4Sn0Sk0nNSb2u
QRtC7Cm+rxEYku8ii1z4bRzONhp8g8pOnNhR5loyFoIp33yciL5vwB1BLzBCddKm93G1eZJI8JZY
nLVfmhLvbga55+syX1UckkHudIR+nDHVGPC5ERnWfo36QDTG9RaOUyk3KzJfMK42Jl+gJjHWxaAH
m1FXEy4PE8puJkIrfmd+WxC6KYIPAzOME8ushLq6+oBPyex/6nQT5kqNcgfzhhgahHbdaUGElNgl
JJKj64s2XgiDxOKjjQxQta6X1UnkA5VUQxMA9De1aBfdzqh0wXFbZqLhrM93/6e4j6vNA1ZS6ier
ykw+RtaK5xw0TzeJdk/URUKip48PXPTtBmhlkVBr2ER6R0OVxwbkVom5dkKvmT6CrlhT7V8G7gax
esvTHnWtZBfnRY4dhmMj08BZcqeEyETMg180Qelv9u3bCNYbdGi2taB1tbS9hyIvzoa0wiJYkBrp
Q6ScOGJB/kEpm4Unkta82nlxYwTZB/8Yr6kwQl7bC/zHboiscGmygrILET/s4GoiDQcJJZLvuQYl
nmcBndM/bzgYwPmY90jaQsV9Y9EufAL6IyYGjFq3kfNZOd+Xbuw1obJndGVV98p1fXztTMYmk5dT
ICAfOzSgdYJxVC8W5o8cPN8XjbMFB3QUESB3Sjs5qE56V7Re2rLQPAgtye+0dXyrkNsKZkPpjst1
a2PslQHD4qUKbxu6HN7s+f6W3qXGd4n4tmweQ3xZM5eIg/pBXWaC5TDiQ4tQYxWmUUh4YiPtjJDk
NTBbz+DGW1Th/jEzHbF8kHZFgWciIRWV0qcpi7BA7dBUJQqeeGUEuiKKSqfypt0VDHb49dZ8xfWq
Xrt74mUn3PQNkXvl0iB987hlHzZclzyMtyNQaev9FuapUShBGGyWe3AMsI+sezMMQi+d8QoxXz9A
RusrOB2ESz4Kfqzpi6svntaRLVUaBX9yJf4IGM4zlmIV2U5ubNo3CRGj3ep3oh2OpHVmFKJA55KZ
bE+n08L+2PoRK8YihqqOJxL1XCY9v/INaYcW7nh1Kzj1is4yD59ttDoEunnEJ3nfjObtvhagHSiS
EqSWjLPCnqD+Wm3XXBAd9tR/5XBlwJNXkCy+ZlOz7XSzqtchIjVxHSVvAtDLjIwcM7ULsbcSXGAG
aTsuAstOg6KrNlqn7hvhMPlOIiM0vs/seDwoChsk29VfDIvAVOQYlUGfO9/esd1gYzh31cAQV804
W/aGSqmsJDAyW+HJ+sHiCA6pd3MWLr42ZGigwHlZNARRsiTiDBU4jYDaBNuMHa8roLS9I9RUVV+j
QyOOhXSgJlF9itv+M60U6UsDccATcSzGw5boUOGaMbC7mqzDoD3BEQ6yMFQBKTaH2bh1K7PttBwU
akVYhFjA/Kwut49M9wwwMvCLEKouF6mCuaipDisyWGIJ2L2r251zvoWRUMmFhYTlQCyGgvrK2Kun
IQz0s0Ve2RIx2yJNOuIGzT2OVSWgPDcuoJKcG3thsiyIy6QQo4wpYEKc8S7OM5ycnNVqwX87j74r
X1iLK++ZzlTrPPvffYiWRHXpCf/tus1VdGXoRszrfvQUAUtwvZrHEW/KY9CRkxABoDbXs01vwyJ4
jkqO8EMrVcct8/xXDlvAOfjYJMniB3eLjZ1SH71U0aaJFzYN3cSP8AqLaraZ/lAMFLVmGlfta7BI
1BGbCFkubGhxmeaX/VsaQvxq/IP5UAkMw4Q/xEjuT6SCszjv+OXDz69ZlqvrnQNSiNoqkgg4hFJn
yCzkIGR1Ewh37wiADeNvz1uVeQK+Rw1ldwNjPvjHayYlf0+RkG3kTYk4ty3JO/CNoxEdbBNfFRFk
Wu7CCRUIvRvQ3M+p/Yqs9NXShOst8MeVs0f09a8pxuHrD0ZmqCLl8gkrSaX8vjc0vZnhGKtSAIaE
DEllrjRuijTJgQUHn1w0JiXwEXLNdAe/wmYqrFOW/8BDXmgw5WpS8IR3ZRVjeVns0E30wBhpX+6X
uGyvNytV+00DJ0Na6DC5W5c/dJ3+nGRwrKNS4XJ47cuTf3EJJU379aziaY/hRMaCLIz0wPMxehpx
pAG0I0UP8xlrgXmEeYi67slfp7jMs1wy3rD+dAhjNrkVMZNatKd+G9hUDCvx07aRmDFMCryj+wVh
4mjdZBn65/REd1Ps3C43RofpHKbKxU9nR5PrerAGvA1zbQHOe70ClsPZ02riAT3LyeSFhEoVcQRY
okBvOljd6F21HLDBg3U7uPa5bcczt2+94LBg1jz4Ghg40XFVBK0o03KXyhrYTpIJ9IefrrAesFEm
kEV2vNLkGclrIGffEVCTKHFiJwc3OnAs41D63zDQ7NqlVYWoWbNHWX9aqxSV6NDv9rQSKLfY5XDz
zoQFjXqNYnepwNgo5y1cwc/OEoo7nf86xgUTgdvBuggfdiQI07FENMQcLI4Cv9IEQdk14FbJX1iW
QKnng3kU9WuHbV+QadqB80qA3lKVhKmLV8KQhlXaxmBNRHmmK2aCGI2KCHwOoCisgGWOBFv/3r01
NoSMYgzCa9aEa+6gitVMYgfuiDDTqzLVyicKayRGsy+uzWNb7qkFwWwh8krmbrF2D97rPTizWfBE
+h5bX0Ifd89U0xzdkPTBfpJrSHJqnww86jrXfEnmLRdkBBWDaJ5stgBpWfdmd2dE9wwGEtEpF7OB
oEJ6j3Xe9wWIWq/sYBYCOBNzoNIXRtisEzEkNdTHBoHhzFYNjxwL+LaVDZTyUdeaIzHmHpTbmOHT
UzVCpXyiYrW8isra9zlUkCqJ6vUZ7j7m/URlY+5wjMrudS4S8P35js+MYFuxbHemGQeUktIcExTX
Xdb8sLzGdCRqPh2+J6vVi1Xmaif+vzryFq0N5zxXTPVEvYO6jKFGfKU1OfHmFEk20vCA5Ze4RVuz
Yt5yJ5mIJUa1VSiLi3N8r0fnpOeoeZ3wBruP0PVVzdR/cL4e6Fh+o5Aws1Qh/yQOhoxoYpJEkSZi
uE4MJ3JkeAFZXS8k8UXVEwURdMP9fwy53fiOKKGVX9CCrA0WFV00FpgPgspKMqbY2kgaqCHNrczv
Cowt7txCtjtZ4kMy4fbuqV3XLABIhfP0Et2b/4/ki3qdNdMlq/ShQAzfY2zUNkc5iyyTND/aZ5WX
WGrfLB66e9ofDJjBwJ+6XRxMZt8fO4UQg52KzKxcXzSls1tGcmlZFCyhVHgJo6R7tLbe60IkYpq1
8Ep/EJXAJaqhPBhyAyLIlidV8xUlDBN/yucYOSWludAtXlHGaqadzKbC6uDt8EGz5vfczwLGGxjO
1AUOVINX969mPagRVt0SRN4vyBHlokpZiphfTUzMQAXX62+C//TgKz4iNTAg5tzeOXYrXwbOLjf7
slIry3c+nviwHKG0AaEyemslOY4kZbfxHT5+PABRSZtzcRGsM8Rs5jAMDCihej1JIsagggM+NDqK
ZPG5qrUIhmEKYqEQwYjklSqN9EFXxRdoWsRP3mjcT47w6epTu5guRYChmvmy9OIZoFTVJZXHyB/x
9zPlbhipTvFku4p+ZXyVX+liBlsW2fOGoC7xXPVmCD7ftJsmNcz0X5nlXkFph/kG3JOxaSzrkywT
n16j9ee0D4mTEpfPCDpk7oVd6q51fiCyyCMOr2bgTVBDaqhUBwmSfq1TZzAKeT4XFFQqZgVDZLc1
wAwNZFkx5cpDRrxPdFNr6Ei0IY4yzxiiG9RJRSqf77bfU6QZyv6jP3qsK18VcsEMP+HncNPZY5wL
Nn4aVKyxiRC2QX2kQrER9mu9+8QMD/Nqs39nRurC2Q5QScbKVYb9FJZ69DVY00ToNh30YJvbVR6G
aPE+NTDGaH6cn8hi59TGFscm8eiadtCTDL3Qf2TjXV4GqubbJZIpXKTu7E3jGgfdc/awl1EnpQsB
xlSHxQ/9nUSzI+NDLYvMdyIoJ2zvPSIPfU/2DbJik2TIewN5MQSPjdUIy6fXgCWHQER3jKUjLKdS
hk5hACoCaNNsBvhQa5Y6C6lTM+PK4CIg5GAtMKc+vzmwb1SRI8HplANjTZDT3/KCy3o8wbbPimA7
qty5h9bjqatvTFW/9Drbp2VCEb6cvNqEIQLSqCoUgsVgOmzS4OISbRcUWeFcYTSmByUj0SHJhC81
rCXvGYxnSiiGz4ma0Yqf862UrTw33k+Yp+hGMN4KXhaud5CF71k7HckLSnc3xQXG5vBADOM8WYST
YwWr6qeZ/s07qm/E0hxJ2RKVN/FACjwgIiih+6ksxMdpccq3JDCFC+CSv9oEYSUugVOu5O4YHae1
ItNU4oYNI2igtrYUSGL5HOJPxv4CdXmCjGF76AtHaBwQvg2eB4H+6/XSwsxO9aWbB30vUYWpbmlG
iD5DT2RyjMaDcR6TiF9qRlyBpyzG5qvaxxmh9+1SfTvkJ/f9KtQ+leDYeZyziFtBMjpSAxsN1CdE
4maDNTQkzjvnZN9UUpkkZFyA9EB2N2qdKbq1xg0Ez5miAs1frsoap7UMztObRdqDj8zqS3WlswCZ
CnjWJFOa+a92bWXL+OmW8pMen2hYb21b2Xv84i+DnHLz75Koh0TiVsF2uqu6xvsNfnbWvUw4BjSz
K1w5tLj/S2sJwOp209oPlAwCdFkUaMURlTligjX3D2Ho5ENvOI8OO+Lzb/0DmYYd/CT2jvYlNlS5
zNdiJHB2+LPgiYJUjy9v2Py9X/udJvYOaNeaYyHyZQq7q46kmHSV+ED6itdklQFw27EGI+M9Be6R
7oRTkH+7sRpjfGCUfzQGj6XsDkYy2eyYn9sMfUnrdgH02A179HqixV2ox5woo1/k16u8Hvs7Foz5
FP9eIYROyMVXvJTf2H8k/WSa0CU6tr1FDp8te+TyXcAz/Tl6noMCd4zm8NXI/yutne4kxfMfAfEg
JyIiA3YmLRv1d0pGbBiizmenaGwSenAsXBd8wEWF9li13mFivvMKw84G+RRwLBa3Sv19K5Din1zA
ULc4S4VnzGaJrsjvCoh3smlW0+Tz17ztVLnOwpxuRBkBM9Md1+Tn70cb0UZyFapZAkK8IXh0saOk
O2bQ2Whuri+prn1dKP47PKIW5lD7HzuLSp2HYi7pO7rFiNGsSmY1B+E7GZ9gz+1pDyCxKHbDoXqx
Bs1QbgQbwVNbD3LJ4QOkBluEuvH569Hmdg4WO5DSpzC0B6m6p+PsdnvFSnABqp4S4m8mIUip/dH1
c/27HMImmDxQwJzaoYdiRIab//RMcC2lKfNCA5cZjeYQNOHS0hJCVe8DMCsqUrbQYSHeC9YVls8n
0czVnCFTkFXQuBQR1IytwofeUXnkExfXFVzOFsHyiyvaHJ20qZNbpJ6pXxfJAxSYvXv0rFQQ/Quz
BbMpiqExBwhzI2+KSxhvWqbzEiIDvW/KiQdbjQalfXjDQAdCrHvxAiliakJcw+kfAwxu57kHBJQj
TPXlwSjDLJ+cXa6kihA6X6LG/6S8D5Kn4AHq+DSnUY78GKXB/5fEfnVqh9gv74IrPtKJrDj5LgUU
6UcoxU3Vj9XXuKo6HeA+oDllljOxlTWrDw3ulWjjcKilwXE6KvyGrJYdkfZO0O1BIrGxP9iSxLwF
BKU1zUa5lyQXF7J4CYnSvrwIdobxkcRFf0DgX8euB9j8QcJtnuh9kPhK7S8e0ttaIrKcdp0L3sqq
046uwhwRsmPGazpGaRZppZK6WNI+tkP31Ys6kFEyaJTYjw916Wo1Ltu+qpKXbs3vQSv7lTzjvJlg
STA+qzKjvFXVBCFZmNX3GGmCwn3gENmYHv/NRFH5Lu9ikmSdwX7HdUT8Ljt6bZxmrtOv6KnQWIUt
K2UlQaKqXc8luoMxB3KAb+s4ptNv5vAdLDaVA+GqWrKQaZ9jp2zq8T/Q+DBiv7LhX6yhpntyD9Cc
ZkQLRUop+rbXZ9B414BK8naD5GP45H6qo6fRW5sp46mZCkdAQgFsQneAvZyBal1zXG6W4++oBWgP
44gWfQL3MpyXzFEux4yQLFRMotggm3Lv5NVSt8gnJy3fA5+mNuuOlBpMIy349G4ZuHQ9EsSfRjtW
chj0D+QosMLCTzNGshqq+FWCTj6zLH2JnBRYMA0B0kPAjo6omQUvWP7vILHUkthzpUw+xxI9txR4
JzXChdzgFNyWQdGqnW+/LUOiQOrd7G4KRCTRrvQ2t8OCQStaOUZfHsxvajiB27wiHxAd3wsEvc9l
+2hN/xFE4vXdqQm37gjFR2QjiiaPH5mo82seZolp+cGJTffDInYWAAhi0wfXxIX1jN7UIL+MGgXU
eXRk9iQi6jYgU3uKfGAdvoC4wn1CqilyUSF4Rw7VYoMJQEI45fmuB8GjoYYbHUB2fvl7akYxOkUG
CvDaVgsAfl/by4MzUEPytzBH9SbRbJiaAewyn3TpRkQkaSk1BUOnMRiB6Oub8fmmXCOyAqZoSkPA
6PGsaGUVudIXo1Yco8ZBMKjEN8HTKyrt0NOQJdQaz/6F4xcyKQFC1m/BAbVlmgO/N4ZqiH/FhqEk
6N3u4S3I6XAKkZiA1EEmnDF8Xx/HY6pNx2gTqxMtI/C/DsqYMpnQ3nTVoDPi7HDPkT6eGWHoPq9O
cYB5BPwTjX7tkOCAZf+KbPaUJiX/2XQpmt36/K0qeivUWT7c6D3slEn6IIue4A23dFSi5c/QQPag
GxlKi74FrtSLBO/8jdqAtgYzpvmBSnlvkUuSJ3dGsAuABUKSLNHHLp81f9qIfO/kIlQ7ttc45L+q
fr6iqMw/F2vA2tvwE9hJcbaziLUjqX2pt0QZvQDATe4zy4egfGkQXC+8kgeQWTRdNQll6fnmrAcM
MUY9wBJ3tn2B2Tv/Om4s4OOIVtSCxlwCE+Wrkk+B+7xJBhpaupaUcr1DIY60X4z7wPTbueo4yiEg
vWZShiNJxOCpsWHA7d1T0CcUpKe6kMisHGQ2ukapgXRwW3veykaxMYv9bOVKW4WlB/8djyu3nyPy
iSsr73r6i+flntc69kVPX05rm6FOvoI4nV7Fh8qmSWA1dnhzeWCaCqehQyForZ41KH3g1ae/9fqq
wixICaDT6LHiG6hKHqZ07JIPyN/hUUPbGOiUKJ38rVYZcr/bx/XtpeoJjVLHBM3iUrvqrwALC8OQ
kNHxescJRYcpGMpl9r1LyM6xam4LIVYQ1rtJx67pUPL8Rj1WW5xJvADoQygzR+zyV4NqALPaM09w
bco74M5zCM0nwMZihHXvuo6zVh+iXx4DP1uAklLhZZMN3we1YRbZ7GUlHKVAxuOOO/M/c3yTkcot
O7e4mUKzbyDGJ1ajBsBh7XJF5W7igGsJ097HErDYmXOPRG7eYCR4AUEGj2oz0Yz76tENj85cN9RK
zy6ydDKS5zuDewu31rYNs79BpFEtoxY4jYfEk0Uvq3XY4O/lB+dYVs7Af35CVg+sE79gu4Hb/WIJ
JuS7cqZ0pVqUCD8WFj+mWbd/uAcDTH+Agodqb0CmFESyiJnF+oCRguCJ0tIwwzHwzbQ5RN8ALtEQ
mA4rW+shsMxAYPNPFXlxGSBT4IF9Rf/UPEMGMvqdzp5qjZqre0q+ddZKLM2YiCRK836V9UdulZDF
9YiZAcQw1ptjDWDwiqsRPlCUO4Uq0JZg1/sQ615Wc+qWERlMBcB0QlotrTNKdoX1hg2vgjJye4I0
yfq7H8H6Opn9J15AGFqhuGmcKVDY8SHQpC+rWtVStehdlfUmXuwF04tgmtkPkraNn26DkgX72jnE
S1In4yXFuV6GAOnE8AHnqmX9o007rG8wiZA5OfJO8hQNKQZgGvRN5V9/7C4FgM1Quo4DtTvdDgSH
S2unkVNKgaaDEtPoOTKT8aZOFxy1LgiOzdngcpxN0EpnOQQDBCz1D8ErUNMu0Hj/V5inuB7tJNFI
a7Emp2OWBRvBLt8YYPE6txi7eQVdLXLddZFsL1/fVmlDeFMGA72U8VliDnDl12uOcaPbM6mT2xY2
C+nQppssoHj+TA62u2rygg/h64vqAm49dA2js0HLBdoToD04X3r6ooR9ApYhNLwtqaLujdBXs0PX
QTnipddrOXb42KaGIBaXa0locyMLXLuZMhnRMN0M/fsWWvrLFxwFZtiNZBAyRGE+J3+f0ohmfFyy
fCO059/vTi2+SOp7OOcROzdiutNjpak7JpdLkCLhG9Th3IOujfv6mO+FnHkqx1+M3/1KybSzM78g
HLoHPpbUX0xNtOXKSDiazxp/AJBEVnIJus2v2n6iXRIvfkvO6md/G5HdtONBw8hjolv0a/lMnd6B
xK0rSkCCIVLdNokj8Vpl7BPFcRAixrt2JEqRpnMah53LLagu48hmQmGc5gAGcj12yga5t3NYuvOC
B/hHpHFWIjyIkhUQpBhdl3vZUUPJyNAo0TdQrFo2sSxlhE/Q82eFiCsD7vlooIoTzUozFK9p+0DJ
iFqPyKzmNn31YmNx1l9AATFmZXM49vFBWNPfCU0jelC9XmqdcYJ2KQtlxqn0AexykgGPuX2QPMMO
GCyNX4d+L0KOKe5lre2NS/UFsAExToSHbZDpQ5NNJOqkihliGzgBeYbkXfypCKEDTbDnx3dXOJbY
QYt/9xZuj0RxaNndhUHEciMQCeQvzv96lMC04cOGG4hV/Dr83hrjx7/dvgfn+MgIsis9ORdBB5uo
83uzTuo1j3vj9MShu5vnRkg4axNd1QxnGgXRi4UufkRjnYRe9/bJMg59G1jpevG3fHHcPlnIiur4
s9Av6tps2FR3rUJidVvORLTJmUIuG58Afx5HYGamcnzu7mvfC1PH/doNt+SWRAPy6gYN/6A+uKoX
wAqOfq7emViJRecuQiHw4C/2trJjmRXdJ9+4ohLXJJ1peD57i2/gj8kRiZG0xPRaTkxxfP80egnP
2VoqELoDk4rIEa9YOcpFsGk+aLcJIAv+1LlYkO29vFRJ/mScEPVZeEfTeglGWAEbPlmZnuOk3P60
U4Zqn3ywkmC6UIG4hcfXxx/3fzHzoOjEaeYuwqKLXk6oPJYj3kfWDkai3ULKu4K0ZvA8rQZsTwC2
pUiOC5P5cmjH9v+R0XLv+zX2eVyV6VDU6eyrk3kXUzogs6Vr0YT11ZPHtiwXiKxGQg7ctoUrZzXy
L87t8DOvGEMKyyVF3goNxrds7G0xHJiVI8zpiMQmzXdWIL8R1zLb38BMiVx+D9yUAyo/9/u/+3RM
Vo+4efwgqqnUFcV9/aRFEJ8g+i7beZVq/R4FzR3RKk4YLVyBs5flGtXQNFOc75iRfke1fkHIFzzy
xd0A3mPfy9el7OWUKXoNLAu0PwnjQIeZxxXLxhh4NYGSWgiC2rZZ5gXbj/R5uhehxw96DVllsX8R
SW8oJHwhqFt8WISuEo2rDaO5AyoDzesBgCKgc0XBUh/Q1MWbtadMPcmp1bbRaoSEq91E08PGohEh
sMByQ+J9WwUYnBxsVEmuwAVeocOiLVn1mf/0/p3rJA7uMM7Bb3f3CsdWUFz39qXmsisRSF3MNjZL
aTX+QJqUfGIRtmQCnigzhDGgxiEDFHL0QPw1G4VjUXc7cO25qCNpIc924nyQqwU0uUHQj53ALpTl
Qz0WtgsfhKtahRGdEZtdKhmVT43a9UZZMKnH6N4djpE8jpNjcTPAcX9eJnAKjxDLL6gYYqOVLrkH
M2n3LDJr5hzHVsoNNZYnHFonNua+1zmgLqeIWpj1+tWi8Y9hlXsZ3Cf6Hd8GLXP1C/H8jpYkDQXJ
naHL4o5GMy2/fvb8be4gQ+F5ZnCsnD1hQ8VUos0lFxGCu5ovxHJDkXh7ODLjrKXMoZwc++VSjd0M
WqqzbA+DJIYDBAFS03wZG2HjlvObh7rK1jGkBxFXzgWiYLNvSu2EGGm7o3JkYTcMN6AAazNDmk6d
df6ezWOm1ZfSADUnm4BwxmaQyyx/bZ1eSOQdClER3czEkMsYSd/MPInBF4EymCp1pzkpWVe98+bf
sL4yQ76mEsO+2iG/HBqPkxTyYC7vifFou32/0Fqux3E3KtQkI72QC2exihVQupCkKDzzZL+HBuvI
wXxJvbYLtAS7TW7wVuY7R0afI1xEXGFEU/oPMgrTB9Jo0Ds/on201ScnlazQKpHhtfGXONtlRYMy
APd1fUcH6HhtOKtzdKVIvSK+2OfLljEh1e00TOSZ3n4SYPHkM246Wd3xbQb896/Z/ecWPelYjkp5
ifraaEWO7de3FvuUfBJBNlA0mKWNVQ+O/7W3J7w/QY3GytzyS/1AWYVo6jDfnNiX8h8EH06/Kig6
n360HiLzDdDiUfIU8rGXNsh608LYb7p/zCCCJVaXtJkZ8LflKI3Ifw+Ij+dLjJU6+A0MeLxVz6G8
bQXxEKJzWw3TQ0SRLeksDDg796wU90WLV4qhzE8ye8G4IzPeVzwR77KeAUmmZJnUKWWr/8bKvWW4
3/nWf/fEljBTw2SpGE6DfmzOfOohXddC7NmE9kqXg6crogcYKL/USW7OrNqClZD+pWoqyVKqmKbh
yLZL0q6ApFHVFUiAtifXNsxrXIkDyPbXQl/+dua0RYJn0CQXQJAyeH8Tljx9PkVCuoDL0gYY5owf
osqO/qOfjW5jdnbXaUc28qRGAT9VZAhy28MJh86dCBt9bxPFcIgNcwvqDG6lXTq/X76LYUIUqc9Q
syDOLNhA3q0K4xIfyvSAODlDdLrhGWvMyNKwl2IlxIYfxvwhhNSLSxb/IKLTsOJ2k6ncYecfz3/z
MLmAhLOocC0uM17+iFA+Ws82E5s9Ik5QIKDfZlgrXpOjxwjGcAuM+hpobpjYc7FJPpwPTs41Ja+B
vIBRiIrC2/n2yy2TcGM1Ib5guAwiAS7IOUUdyYnRh/KaMElUXILdp0I9zcytQt1+f1xcTUEVgurK
XUoIteK9t3cd367cQHyLXYeZVmdXn6BAL941VcCbIlc72tOM6UUsAF392v6P2mpkXiucBaWa1r6F
QvqCzWg+Uk43Bc+x3CrU95hY8yZDyO1jA1gEB1XoSeYt0zKgQZ5Wqx/0q35NShWhebECtV3EfdQ7
PQWUeK5Ara+K7FS0DIwx3rUVSWbS+ZHMnL/8WPbZXhB/GzlmMqfG3MMcDo4ER8W4vu+dIG4ooTNG
wuFv5b83IWCp4z+aam75Z1P5cq7aut6nx6bn2RaFgcMOmRpq4Xbocc+E2QiO+ZGhfvIYW38z7Cc6
X83kSpgJWb5Dt9khe4hNQjkqYiZf7Hsn7/vkCGHdseGXwqH2tlNYwsOzRkc6QRCIAd+rVW7b9iNK
/3z7Jiqovqd6eXP0I6qzxcMvtCFtCwYj+pObC1AcNChTp3m4NHwVGnSmUvGPhSbPOwDJ56JquOA7
Cz9bMXA8SgNpgl8yLwmBiKFfO8wT2i1cwZXBKqV61izTllROItKAsUukiiOsOHSCV2hlUJCPoVzG
NoydeIqVfoYHyi5o5GxwpC0F9FA3+LcXBc0bEcO0Bn+n8/Ojmv+KnH6F/YlD5akzQ9LF38vxEr8V
kr2DVr+4phRXpSMFctDMC+7LTFAy9m9AHaZSDt2s18c/2ShxwMBu/1HqLUCZW83ksEWBPVUaljxE
37/HDuyFkRxXO5BRlzA0vlmiIzLio5PQ1YX+Z7pa8g4TPVTqeZD01kYWCyPLDg/rhfYPVQVETj01
VB9INkjG5BU+RIWvAZ02WPVG505spiCGP8PPwvQJwg84m0W5omNcjaHiK1jfCRUGyEFuAGZSLW1n
WGMfHj2HIfo3SoZSkZ1ODdgUaSPqIrh/jhlMkwa972GR0HD4iaTq8Swo1AK8mD74z63Av/jdo5Zm
4YZ7SJo0jxci/gU6cEEEbDzKVf79I1LfdXKj4RMiDqHBbxTP1EeaDwdbt73AKQLaIU2YcCRkM94H
2kR1rWpkbcpoJ5ndLBFlGU8T5iT3Qvy5BLMn5z/39QhbzWXBdm5XlpRrxcjQUzJ4XpvgZTgvL1+O
q+4oUK+YUIwfLrpms8u5OlahjYlLCn6D1VtKRIOF38djmzdenkiDOByq6K5S3z6eI1f5OZug5sZt
gcuQ/GIvFUkGcfYK50Y5uxsn+P/JOXgashXnOxC3dQ5fBOxsDVe8rb9U7jAdr89N8qYjr19FQzoQ
U9nF8cDFGqjnEMrd6GQQnPiiDI5qUQpT9/a3kHDzWmQrKAdhk7k7+7v5TeGSwtPVH8UYcOoCY+rD
0K+gw3mS3BVpH/0h2fSRqvbIBNkqUZnQM/wlH7Z8N3Xc8s0E+iHtNQzv8L1hF4SVfMI8cueMTnV7
9Si/8BnMfqE0lQYVdyES7pjWx6PzwLX6XonEtxqgZsHEFU4esnKvzOhpaUPIaBTmEdXGS3edg8kn
QoFN4R35vS80RZs1CWIddeBjtpnLMwkZy9Uhha5IhA4U+zgSo6Y3lSQvNRtKkY1ypK7a8D9CdMp+
CSYxMyFLDW17Nh6Ip2DhlPmXSHVN0cOnxpdiS1yKgwOf0KUiU9liHXT5Jo0fY+K0IptZGaGZZZjT
VwLS894S3MzPhUup5G+LiPQMapCt5Ac2l5h6sd+FyalTyFYYDQGkW3PyNOOrd4r8prUH9OBlGcpj
oBmlhyilq0XCDfYWP07VVoPxt8EJuExi7/vF2VL9Ta7vMONuiEf2ydGyV1ayohe0RBkGvw2mVx2C
Ctykc4zAPGhuHqw6pjuAn4A0DLrf1sZ1t6asmzWuQWeQht9Kq2GG27nYNdhnb9px8rSyVNBmw0dC
dOCqnQD4C/IkspjIwDExLV2i6N2oZl30O/wnVs+5oaHzDLzu4B+oZjUlTNSsqIvvnamVcQ1yC1ek
ktY8RV90VHKWA1Q+W4nOxgYovTm/NbHkQoTatl5gZUlSBqLLO0QiPTpucQ/8fB9cCS+OVeNS0xMS
13b9NDYW7nGtsoQB6iHNsl+qlB2QBAt5FTwfyISSYxOidG17o58AEdmouk9/uv7vFMfB8RqsIjsR
BY4K99Y5TpwIR7H7FdJlqm5Xmm/S8naVkifekBvjLpm1y8pjkTS+oEtgVc99JkyN+KCZiBWKLYxX
2nbFBF2AgrGlLmhnY4biyyyrbJ8MLjEaKECcpAZ2EqMXJxNIC7ehg6GMzEx6U1bgkxbcag8qeP40
fizJHpFnYxrR3ge1daSYpHQmGnTaaMlnd30sT6QqaQiL2EH+41a/WYE2PL84vjwZVcj8NiUFEIzh
iO+BsT25uBgWfHykkOOVkiV8R9KPJbDS8069f7yk+bdAaFrgGqrKdMahh1tFUwRBpPCssG6nRhYR
IKGSokIIMfS2PmKKMru5qxt82iWKrkcCUy6UKQpaqqmIY57zvwMIY7H5LmF1FaMs6SVk+onn1Bna
Gfxh3qXQ/43bZtfzP6lwa7uBdf52LB5qnY4ecNFwbzwW8V2rcIe2SFQoYEm5Fvm2wUA6ngj8xWtS
ipkvkbiDmjukBvqQ+HU3hBwW+hGvJluCALb+bd4kcuNpA2Ce5Q1O/mhmOFxRQ6ArSM8RUbZKuLu7
HKBlyvtuiARPRbInctCAj+wMFMax2ZUNsO1yLrB/5JJtHfiSyKfH/GIf0aq9xYxpMVGvdV0nd6Ak
MCV/4LMLn5SHGgi/cuc1iql7/fgo15iFRHgz2Qk1+5m8ULUpZA7pLkhFYNhst5TnQId4sTLX+LW/
mZsp1aJ2uqJNaErt5krz7nKzs5u/IXD8SHhWbj6sajL3xd0ilV2xpUEYjcSXUx4yn1BuiDWeKwtx
SmZPCre1je1mZk5ziuAXNYso7brbR/DmMf6ydpi48IWlI59dTa/IARaHluxx+MyPeYaLt/1f9AR0
FadPaPlna0kuGYvMEKuBoM/dQvvyF0uTqjfvwK0xwAYVuegiLAa2j6dJDk5ZH/Dj9L0galMZJNmd
3x8aGpAGvBNLf9o131E5esZ4fegpW4ZtMVNHBDYZZL2ERxuuX0ooZdfVfBVaDrWeeWfEKSbEKMt5
bfD3BmkwAIuy5iH3m8F01oMzOIudjY8BiiHaMlK0r/rsXAwd4IHOX7ZX6Y0QTwnSKavJrOfWz/nk
b9CQjyaTGosOBmy4doRKv8vUPkauiIsAXowzxpnZ9fR2ZJ/njyM1+0sWwbCHdZKG0IHGikW3UccG
144RPcOe1rfpzEE5T/iKCbDhzn4u4XqDOCk55BozOc0hLjf230P7PnSWKW4v7QO8YMtOi/qgKAaK
TvIEpHZY3BObDKLenwHBQMeKy2JUulFyyoq6gRGmQ921lMtAFhVTGgazpdEvTj2ilaywmI630qXV
fJmMTOjcssS94YUMxTVsCT600bwdsiNsGhOnRdZysV8Mmzusk2w3YrjKvr0Wyc26LEIZCR65KqEV
G+nFV8yCyxqnxn05y+yWSdUEb4MihqZyoDK1f5F3RJv1Mv/v/s2/FkR09gypphlHovci+08H3nUt
H1p/DkTXgwg7+BncoTVoCzouaJTxpf8csoJx16h4AqSwSk7midKmWVbpfIgEMjPJ1IuZ/nkHSRav
IxWM9CIcTWkyfSYCVO80JkyXElSm62zSh56sq42LUkW9AQb+y1e2vxkQeiNcDL6GTA0w0YtQgEXw
qGiiZQ2Y2ZUjJYLM0rTYSgmBuQEikchckRCEio91sgC8RQGMimQI2gMV3Vt4OfiZW0ElATr0gyfk
Djc/M1r4yQXdFOHe8HX8/D4MIhUOQ0TqvJfXHKRPHxvvFi9P/NihWKH0JR0tQIDhy20il5lyibKH
E2U0KrEWAKMXXBU359x+IY6y82AsE5wSDTW78M/+rk82b0DGimq6XFAqkeqTJ4RkmWjGKq3RoYCK
z35Ga5nzH6C/dv6hF0Z5H6nuECFuikLEN4RFkpZE+hsh5UW8kW2IkwczZcmRoHmnp9f6Tj8PGZq2
Jl6H4/4TJds1LG3+tZhOJR5ZtI7Aoq3dChYdCpuFRuTCCGT4Q/wyDUY5Ygm89jNLw76QSMsy2FoA
wEa3tc48xC8FDC7aWbBgCMiYQ4FfG721wxZ594NkbeFBDSnCp8Zhb8YspSYpi4eqVZ+zSAndztfG
2uDMyBVQy60PDWqhvIxfPkXYvx+d7SEHWkJb4Lu8pSQTxGrjJPdKStOpxPeESgaEv6IwZ3hlZCpU
JjseL98HgCup3Cu1AkpkaybGDRfl74wOqlLCbfubeJFHoQ2P+c2iMfEJNbQQf52N75MjTbDv6At3
VczUZ8uYfqviGXq72STun/iUQYG4+8kE0l4082u69WjA4fNuVGDclv+l1fYjDzAspqFnsqdBXZoT
qRQbASXCQoe4mNBrPaENMPawMB6s0NQl05e5BY+QMHxBqx1a6GkxG2KVXlIHKZnfMZcVXE/0aNgJ
F0mWNe79aIwqbXIsoq4fkGQ+kbAelJnnFyViLeAPrcKpVbtdggrcmo47SOkHt5bmHuRflXFJGvLr
tM0rkzcloNeL3rkfzQaUdhz07uPwHX9ESu3jEsK0jMIOGz5SGhLnDU+pElSQqi8jUfYzvZ5dmNBi
85krp9tuk1as1ZpEtLhyjude0ftGmrVtuW8tqZzkeSjparliiJ+CgK1WwlG8GKqweoh+ziH00IbD
XPOHAUtFpoa5I53paht2FQPvAhgVqO8gttTNG3HxFOma+lXlsH028hhQ0xAJS/EEXX/RkzzlxRGZ
paKXr8AKC9dU4BdntNxPHK4K7xLNOyTLBAd+TZQ/Hh9tj2i/t2FTYE6GCckjhx2OFJ+jDdH8udC/
Nb4kQxE/DPbTl4SphIaCG9AkH53AMd94kLIqMcefxhqPehwNDh3J5OL474xldNjWqhfBo+C367UT
hsGHEr/PQi+e/Hrq9RloTBlJJmft4B4mFxTuLq0G1ZK/LiFqh1Btl0FFlW02OnBvejwHa+PxvUoU
+DpGTCxTaDFYU6U1ASwEZRkzBAUWXqZ5j0DeWh40PyFxGP3Ml5bgY+VAhnWRNPbJdm/x+e1+6P0g
ew1zwVzta69ShHItsdxaW3KDwMpCCi9xKYwCzn+90rbMUtHof+dx4dl4Mq/lycBFSUWyT4tyBkk4
1hwyDMCa5nzk8Tdmi4pD9Ebn5Im180u0mFHIIuRQqgbqDpWt/JMTZghAkO4pGq2FUS/DP2aePZtc
3x2hlriAwv3hMaaXool1oAH0BH1DcL79eE4by5PTnakIBaXsELT1fugGJbUb5iJX9d3y9pVVmSQk
SYjhwWXLi6pY1T/dHblLy2fXr8S6h6CsOe01VoxRFRZo2Ks6KspReescg34fwM4U68RK8NGLAFGt
69+4YhbSEjn6z43MMdhRw6W5B5cKsYFkyRoKFYqv3wX5lYCJP8CIKeneeDYLMeRxqOwopH7kZ6/g
/UVCES7wJk/U74VEj6nA2qwTa2qiI5OvWgWDCzDgwgBroNtmDAPGUA9rVnLKlKn1ijel6soNsyY7
x3AW09g0QHyxdFbFz4XYXgXa7Smy9sf4bxMFl7lsCdADaIs7ztbJMUPMnZGT8RvFn03FXjlhXhQu
xn/WAX08QalELIgYKFclVclRq08C8Zi4K6amyCyhj6aQjt80X/5fwJrxK0eZXIdgrzRi6B++vKtY
kji/NX6M5ZdKt4ZVdUZGeWzpAVGT4CdCXBwbWdLGmXYI+OHg1Z4yDEb8HFKgi09vrUzAR9zoDshr
bqyNv0VSRVoo+PUb2mnm7KQb6TMApN/+SUdFawQT/EYq2gkQ+JTt5QeYmCGKyGD3LEXu8gyAYspO
bneJpgyTqs327DPicHhtZHadzbtDBeMzSrk5Jc2kQteXyQPx8Y1rkyoQ9srk+cPaxmMD1FrW2WQN
LorXLvBcaaq4CJuU/q8Zhh2+dACtyfWVWJi/6VFXfI6zhgiDoxctJp6Wg+rWJtz0fIR69W2kL2yV
sQoWR32Jsn4LIuhSiwaUmNLU3NLS4KtQS4lUmi5Ssi56CakoDQMEZbrwTyWGX8pfmVgddZKBahoq
vQvGvGwRphaMr0wkbu/Vy/AamBSX91BijhsiBqNBFRFI3wwzXGFODjNGdfSjKoUkANZ9r+nK+KXH
pK72ooqnXb0nTj976cuRJkHBGRwqh5+CCBLuicKRo8j8Om2EVvwTaD0Lo5MPjE3UlXEKEk5491zA
v35c7boeNeDneWfeQ/b1zOfArBYYjnF3GiaJsrjrv3x7cc4Fc+HSdaKgDbsZe6AX4rgwgPW4LyF+
cmj0fELgiY07ws8pNg3vl4ftR1bxLaxfF3/ZAV/yfq/SgpA39Be5CDMlFr8OeIA2trVGsluItH8f
myhP4Z1qmcIsOnzSexTC0Q3Afb6sEy5QCRFwLgKU8kU3JfSZMJ0eQ2nowXMTmhKeItJ/jPwQJ5xL
Hvcd2In1kOC8E4QLAQJMNUnb30LWlodPVm5Tym9WuPjuI7JftiQ67LOwrz25+k7aWcRFSdoEloGV
Rc9OcpPpB7F+gp9mTd364TNrCaQZzSjIiYYAqi1oru6iR14t4L6qq8w2hk2rlH9Gz+VVigGo2eIC
dGitNNjbGZ9r0RRFJ/OPqX6sTFKW5zmgYe9sM4TEXHTvAc8gHzJP7bav8yGzac6+b9+qZ+ByULLA
phpN/kh/XcHZRm5dQxgV229YtCE90VUmTiBiBo7dZvFEABXQ4xsjKIJiZf97xzP/07mIVx0mwnOa
4v+CabFEL5BLc+SrmNFK2WEgVvSdIVsb3ylgHfeP4ez59/ZFB89VfDUJl6ichQ9R8hU4xeSYwhIj
S6AzMBauoHYyY3dGGHcv2CIzGukYtPvObppeIUxZ8cnnAnCg9NC9Gzto390zdqmeMYHxgA4wSu8x
G6BIdbnPQE9g5CScDVKo3CXpXZvC8g2400aIaqnetVaHuNJiEoxbUTTuzOA54GTarL15nfRZNwSX
VhWhwPzFrtH0pYAio5HjX3lmYia3XmSpbOVsTM2VKaY69lp3E8qTPXf3jTZoV8fOOQ1rNfV9k37Q
oqMCIhpwQtajAF/ku6ShaH179lQ9aUTyOwO1H3Khjo4XrXNxZ4x7yoL9IB+xiGb2+ZjAy/mLpeOJ
ZzMoBdvS9h9yXrpcXd/bjtazct7Yj2uad4VpnOBqyvKvikS/XldWPnRHlfOpEym089C3/XiVKNhW
tbU7OWNXHvzM0MjP7gxlZsI+LpP9xuQNDlXX+GgsKQbplnveaW4ruEgttsg1AjnQEsHvUMPIkht7
6XwKdl+DibQZgBBt0VCkUvrgHVg0/FZjUIFz1LzcI/FLNtXTKKxRfzumASlDjDavP+udWyNjjllA
c1zGl+MAJakg4Wov/ALpQg/kpsJlC+HWwOi7n4n3U4oRiUJivD7V4RTXxnEYb2bvQLA3RR9zmE8m
inhUu3Bi0S/kAhEA9VyAsq2ES4Yip70zTeMbWSmzqvkHclq/KEc3lkSVQe6Pjw5g1brEtLJG91vy
aZffEw5+sIN4e7qSGGVs0hgqam4KLsnkT7/eYhvCcf3tiBjbgsyTsOPOTRXdMwra/y92itJkwNTE
/1ebMJoiDqbQ/CI3ZHLq/wyHDT4SRFhThJmOuSkRRVliU2XMbbDbfpo8ybEWoUl9JHbJOyR/4eAT
BYIeynRVvCZOqZukzcJ6NgmSDFTY4QutjNbKqDMprIVsm2xu4+iT1prNPBP/0CXqL1ejK9ThVtZo
O4hSF2WB2AjRkmG7k3TkY3qlMi6yqEWqXnqeKyI6LNAFf8yXCNi10seQsiMAF6VOar12XR/rQUnC
84Q91GFJJZyDcipJpXOBITCEQiEc5l39deQLPAzM03RsLmfKx4f61EjYtRL5GDhtH3VZjO71jJUT
jwYCoFu+vYla+G/DgRq5qDEb9qhXBVxNki7FgS/x65TbFRK0kcBzybie3K8szw28lvv/9jobqA+L
DCXZKi3qqS5J6xY7FE82dN2SXn5eCcVNu/LfYQPe4kCsVlJoQoe/oVA4eCDSI6D96naJd18sf4Nw
mswekwyWk2GkBa8N+qdLrib0up+jZKuxo5fsdmzKtwQLEB4w4y0cWlUrO0Mc30yrnMukqD7a8B+D
o6HJLEqEOfzH1l9V672HHM3Kz8BgrIh7p3JuMNpO2UVHrYkCvUUTCQX3P51+/OxD8IOPIsMe803y
JZWSV7yO9tBrAOub34sTsAHCN7zbcCBScLzUe5qnhGOdpb++FZ9ZizmZ0pUT6V7Ghg4ttIqBqeEB
y3FR1PgivZJVVm2Epx011h+Y28pRiUUSKsIO3JsMnIYenGTrXjbOAZb3G4sWW9GdkxiXkGoKC+sk
0yt3ASDQ7MfTY4/n0GV/DKLa9jUuti4DCmB8YkJNksR336WDOQQ0thkk/HyTJu+3fHVzN9mCGAiw
tPskgQepd6rtPNoH+p+JoYVCKQKXbdZSL6Mv9qS5/NNy4fjOeXbpLq2C5CwjikfT7e97EgQz2CdB
9u8rv1fGuxEfxCa0TZ4+LG8eXgV3/oAKNDV45UaLfEZ+Q3LOSTTEtSlDIXTniJT7VHixZEXqKCjT
IlWHnF4Ak+S/6bH5Zq67L1bOfl/hAZovbzs73aQUo6z/WBmhTm0+m9al5rmRzsnIUNm7RcHYp9xA
3AtJUwH6PCZ6BHIUdAnvxHSajtTosfDARdxMSuIPjsyoBamgU/yPtaSKpjS3oLyCW/WLUfAhkGuC
/eOcdXJE+Yj5wcsbNj2uK6Uq7aZx/Pl7V/ZLUh8Z880TXk2EbjqppDzo9X5CXfJavyGQ5iFa5emj
WSh2DA7hkBakv7BMpb7qUpvDl125k/tfSzgMMTsheLHGwTlYBVi8XLlt2wiKvzPP4IWiHySs3GU+
AuWXLJeWFdsNDuBQDGnSDsJuPRTTc6nwTDaEdf7h+qSbSfdOyWj5k4bRJDX8cw9GZ/ef2bFVYG9o
RMRkSP9G8tYEE8TJpTxYUNFwLXd90HEleIMwuQGutLUmPN/Zz22EgdSQ6KFcXjHBCqQ62C0CobES
MMnzOrgmNYZz6A/t1f/5mb/qqcFhdp63GGJI9Eoqj8G2BJeih06OytMxqr4cc2WjQw8yuhSTP4gH
2oJUSLVeHeswZiQTh/CKZzSvrrhxWq+2VRZ6qmHHeytOeFMpqLE0NxDMFYiVcDTYB48V4E1hh4FE
puL2YQg22d5JJ7qhYDQMrTqyLK4dGoCmcreICjN5wO+1vIkWWWtCw1mjK5BNc4uVMTlE7NwIWAPa
2ddwutX5TJ0mX1TN9kTk7TOThTa2fUw/lnIUedZ0GmjxLMVOVoVAbCtu/l+HaBxcaVagVh3ktpHg
9JBkeMraekmMfK9XJCaLqLdtWrO+ibw1oXVwrqMDZaENpUlCqD49oVwXCKScR4aKbEsRcGYp+OPF
TdHKDCyPIn+bUuPRJsCvXNRhfZ4pV+9SHq7HoIGTDxLO8huhyNbAnSefVLTtyALAyL/rQ43lDKZz
nB6gvvauK8YYGcWra5kfDnQfNZMOaZ5wNa9ZAwJ6S+kZotBTCff1hTW9+bZ2LovkrGfUB935/eZJ
RSZDDBEDoDF+iGKiXCNlsVSOKCl65PnW81hpQCYEVl0To6uudJfphfCcgxtHk0TK6S4Gzs15cLsV
dh83LtIxPCsBy0O9JrSAnVswZlaWVnGWLJCaQGKeKUYi9c84AQ4PwW1u5K3PoRNZubYEiRyKHaAk
Uok+KYWlsdz5adCfbZ6g8LptU1+WX7lYibRbfZvBceWu3DI/TfrFa8ESwxMTmE4uXMNGhIf5/H2f
bff0lXofx9MglFdvqYnQTkcIoUQ/jL/6oEolY39aYevOfhmLyzV7S6txe6nfCjfEaI6ex8rbdP9J
tsf1JgOF7KYN7R6A+TsP1X/AOsMOxAt0mg+1i+tU4H9kv1AsfGxm7TyMayCRkzG8jRtIvFqUaesp
0EssScfJwSe8w9jITXKhSR54BLZ0UQGk3yCnbKo2wSHRE959spN3Curyr2vEgyb7YltsatoXerBd
xTmQPDOoPpTMgh0SpkHwz22QqYD2/HzEcQeUplOCaS5ro0p06NFzEm7YaEPP7Dx+6pgwVVc8Ka6S
vE+KA9C77cPmTQ9p4EWe953Om91JXjPDSeLV6yuRT9ZtY8obmmNakFnZP1J0Iqtfr8UPS3Lrl6xI
CF2dhMYXLFEQV1sPjRdMlYlCBSGX/QlUEP24hxPitJeeD5n0BR9965cmNnC3l/Rhg0kAYsdxPq86
N9RrsjUFmY5gPvXPhFn9u2ni8ETS247Fi8MHDMWjPqhV91mAWxucaZGgP0jQ5z+bfqS48n+6G+Tv
6hznOeSrWfFreKe5dWvXCtD39L7cRewYJK0fveX50ZYxTm2D8HnD0GtR8E1d/xtT99peVlbSUoJx
Xyx05GRZhMSRaU8AB5dHW9sLkO/AbCioQ4OMhPe7nrQcO0n4/Lz4bSxYgxa8yRL647m+KSZ38x7G
fUOKd3wCF9zhMNyQmL/G7YcHgn0S6yZKQ6Ckv7wVbYUGSkK8fEXu3IpYkKejrSgi2OIC8Ss8pLCJ
BBKvLGK6mTK+RM0L2pN/z6vz7vplS4rVWLk0w5/BZbTz+moa4+ynia7U0cIFbltlea8pakF+fifp
qK0/ijAyWUUFUIhRVlpbzha4XYYCW9jD/xX+Vqrg5brBUu7zTYj08T0Bpe1y78T6e7taOFO7K6x2
pfD/V1b/HSOoK0X8VHsEi1X4odJuuwXULhSU85o3QHdQmNHxAw/yEuS/OuKHPM5rVfFpmVc8TAMw
q4bdrvgTmDn7SeQhu06VMuJkIePs9IS5hJU/TVvXlXntLkLMY/+uhBLPwP2XZ/BZL1h0jCL5S/Sq
hyP//iETspJvCUIxwhn9XaEluMh0XF0Y8qbTGHjocTkefTsdSQ5IEp8eT/wx59THTZZJQbtiFNAL
jnEB1AfOiRW3vw2HnqlyMynJRRWDypLuzDjwElgHLjFag1Pi8Rwg33rRRP/q8B7YU+AZ1FKkWj9S
EtSKRyPeyAvi7PGCfipP78EovIaKTjbXdwWTSi0teox2W5DMGcDB3Pw9qOgIb9SD/MhGOl7oU9Ky
PmNcZcG21tlcyVsKa6Bj+wLZ/H+2GNUFozia+WKlfr/aqeVo8xbJHb6x1ZGsejE6/q0KmWC5e8Cd
fHSxSEaOHyHcIkVMXlfIldUzz25Fm+Zs20KKCw+0yQbfzCHmkcGMKpo4ttXae/bfUeCcJnm6P9zt
SoLrh1DcbEGgShbZPuzKGs5rq0iAoe5BtXeiDcnIJWoF4PN44Fqr3dvMJzBVb0W2C0llmZdaUhqj
5XfOcAnsTzSYAzPmxL3VgWFBlFIzYOz/cJB6Tfw9dJknri6wAemLaq2UZTMqdmQXjEtvasEC0VoI
/pBF0OoZmt/y/HcN/v9Yb6u2KmBxCsiQ6EofdMcfkgBM/9nRFlrSiC4aUVfH8xsh0dQB79DYI7u1
Uqq6HEab4c32zrwpKEFHyUj0LGl0jVBs0FwbCLtHvnIIqHji6YiBM68W8zUXAGc2njdJmIShg3Wp
9zAuYO3m4kZJMsGxOHsP9VyNWqXP4+8kLtFQdLA75rAXpnb/myaAG/DRAhmP621cNqVDyZfQUkNR
jhfK9qKhjOuL+BBlqihVoonHPaQ2p2U4/beH48jgpjXmwmOKnaIGgJMqS3/p7wcRCUJQ5gfA9iuv
nctwTmCxHpwq3E5s/8HZhgpr/51jbP39bIxm9gmC/RlkQzqp9whPGyQWgrTE4l2pzvpDBliv5IDw
qxv6LRmTQ0Fn+j54Nj8CEekNiTRlnByOMx2nNInExLueGreA2crQZvp9AEm7UWZ4THKcWc/Ig0/h
/AB/gOzAZIPeEqAzXngUq+KJ1mCGo5stL3wpftic40hnGpemeA43JHaMc63XWxTtLZtzI2wW05wq
vDNr8XnmO8m4GU28P0kILEiGzCzdoYb1AkBVvSWRsn/3+FHGkHdQc2yukqeZNHqGLPadMOTydGkh
r0BIAjaKSvex4UttPd49dsJbviIvUJraL1PRXhYsqsNvdvifyco7fWwFS9kUETpVhlEedjJW/FHb
ybLK/PrFHubF564lDVHWyzkVoVlgMEwnhSGnn2YmNWcValwF60ikLU9kNmjj4ZD+q4KfAr52FY+J
KVJc/qtzUgjBzjF+lHoeBWHi+HDoXL/TKmjSb+T0l8cBpNxwq6tgG/WVyOfIO9roLZLCH5tsXnhG
dtU7B+jkqfClefeEcLgl5Sl0+izeFCaRwHwc1jhd6v3PLn2APzk++3s4fv34pvH1ohROGD35UlTJ
OVhj/n5H4IuNCzxB1WFwR/cHBNBblpkZWDzhiCJ9DaE9Cm2coan1dn0Zlpk2i2doULWR6WVeZgjm
K8AmSp34F1MSpedkPjCCffbDPUI3EIeSttJjRXCxZNDmj/3ozjSA/PPPbsPuxbxvtwIqj0QInlW/
Fr/ykrcUGU5xzUHwR2gSvTfb/5q6VJEAikL0cBjgJxJXRaiY41qSYHSQWccaZop5sHLsxWoy/ysS
8tNo8N5dCsLHYJh0J8WDRY57UjDV2A1JEbf3NZWF+OwEAHEovqdeEx2XMe6dzDyZskHfz9STu2l6
AidsXRfo0PJ8I2FmDepOtg4Eb7rjyoUjCvTgSh0xcX/YHrEgzzLmG0796/Yj52xFk5k1WgPlGtcB
GAP+aSP7R0NDUaAQRJgWOiFzOCORx9iifylpeYviBr3nELuQRE2+eFWM0pede28iUB3Ot0vpAIxN
ghcDtPMTU55vTYoRgERKjyz567kQPfkzr2f1+K189nioSZRkb/6FJ45J5bWMmCZ8DUhQSQrviNFp
XUWdTtSL4u4smpgBaakqBWI635JdehKTLKiwlkbM3YOfg6WJwOVwHLE4PvDgsSo5duWztEc5jKZ8
yWIf1lFzQX17OzW9eQfh9Wqt8qcjxp06Qq1Pupp8b7IvJIfRB4+pPNM75hb95c2qzgPMRNxjO3v8
LGBJyZdHNdsIJf9sh2v1iE7ETaiWKyTt0CdyudtYWLaN5g23TNULYTVeKGeF3TdIPMtHGzLkqffO
f+B1rhG+/ATPGZJ9GcFlxaVTWqWUsXhJhmCP0+extVdE1T+AiZpLltPp9jfxAXXLqDC27d5s2lCT
FlirHahABctZE8nIRlHewRVUF9JBKTVcTn22Tx0zzIaAUqPNmelhsM/MfLlIwWlf1Dd6nWIQ1WpZ
AA38179Yw+Fr7tEptpjFcmbZsiWjGdFKUqv1npimgX3+Ca0+pETz6lNKMj3fyuK5cLM58Ix+cNDc
xaUjEE0Me7qYCwo91eqjGKdJFoJSlW/5szkqlTvYSuFQPYEtsOEMG/STrjFMkWBB0FwrTwDYsZz8
QMiFxZcNyz8dXyin53dLjZeIQ9JQkaqEW1inMtes//8bjmnZb3GJjon/kUYHL6+R+GQOub1E3PQa
E8Gbk5PjMXNdx8Xb6pkxiz6DUkaJbZ5QP4vOK72F0LuluWaQ5swVKRF7jK8ckqOFJdefBzRUK456
lFnHcq3GzuATh0nmPSIK/fi/JvGrsXsbiT++Kbe553eXhLsJf4x7hKZSuCe67MTjIbhIUpz+tY1u
F/4F9pwsqldEn9NDBqrjSSsY+S28i3ZyW2Bsw924t4gPLLc4IysrrUSXFe8PF37MMDuGTw+LEnWk
0YBIEFcqVPgGPQoEZj5RZblJbAvLQq+wEGf9/Xg/XJAZE/UGfIUQr70OVU+CuRNILVbzsjDHDCM1
3DQodpYll2fxjPVixmb9/6yytZepeAD/Y1zrKXmyY5/3BgSJHYncsGKrysyrEsxl+4G08UTuoZMm
MajFh/lFdqu6wjqLimzutYAOKqmAdALUe/15qDlveCzlCv6l6w9hS2ayLFMMEHoViy2Zd5HZre44
Mu9IVT+Ob2mYPru1Z0U7qrmdc12bfkzkC8L0Pk09Ae8YNW1qyA40WkWJUIrTdKuG/WU7uRf+IhuG
vlW1biPPaUNHOhTEo8DLp9UKhQFjr69EvOLIdWGkLqAT3YXyKXsopQqsKKEup7fOfe4LzQE5W3pc
GsV5VUOs2k9ZPqyObLcO3wVRLzWYCMi6BUkNPVc+n9YHZB3ByS4kiaTHwVLajwdvG7WLW1s+XQAw
wYCWm3Aeq6yC5p5NJh40NYfC+Rm1z0bPLUDyUpsRHqrNWxkVs63pCGxBJYWfsAzkl9nI+oDV9el7
HBNfuuPzrkI50PDYpHwh06MhzK5OVkWm7YwoXgtVJMM0/JQ83Fd+o5iTH/9kjNa2OTsA9Cyeequy
OZU4DfOzpgGPtQc3XBmng9CiC3mOxRcXD0Z293NgO4g8NORJcSo6JuQoqCi2qXAUkCYtQSV8kl9h
Nq5ST+Q7XjDj9MomfFXTimu39qzq7eQVX2vkzACPvpWh/5lSgT0GzrNZgYMmYK+6Hi3CrLS051di
my5vnEWNdr6HJ2tIjNGQjRUQehPxsW2DDbaPee41j/JrlQ0/J9X1mUkdkN2gu7bk1R7P/AYexlPo
KDVTwq6wTHKeVPLD737c37LAGSLjYXXRxfw+kdLIoT9CJR1FHs0muBfpBKWqQzr7gny6CP473GkG
62leS7ly3BKJ25Osi3OTNCbzMzgFd60zP5K9C+mTXOcBOdOq1Hvfj/EtSaP0y++Rd/dvObwkgwo6
kBQSQvx55zbe16wYDYen6rgAk9RNU2Pba/j3M2Hx/EOhlRig7zc4p5UinWk8VS9zu7NljxTzcd3Q
7ONJlCPR5T6VGB3VvjGJN0bNxRWTsdd1lY/6fyI5ru/Q8rHg8VKHmvLv4u+QXfxYqNwpjuO/MJDl
uoHLtwYjoablafLQI9Ts44iw1O+UVmD3gtPHz6W4CwZ/4miDWuBonhf1oIkWmu+86+Z5WJpnenBY
qbsccgzA+ik2hQfhJa9XpMg2a7Y2hjfTqQYCz7J5fGERzNPFmLzOh/yi0+NnBYMZwWZgyu7Dxc4H
DUag42o2hHgidVwXNsM0CFjH1l5E3sIPiVFw1LCXMgC78xed7OBp+1tw4w50J2vwz4J2QXSpb3AB
GIkYY7bEAEK1uh9/aFc94EYvm4/0k69sT08V0G5vHosCqt3Z3RlNUdyK2At6J6h6/is07bXEZI5T
nJmcsgYoxX5IbXDltS5dmmByrdv0on7OQUYZhdYiXLhRCYjJ6PYWzzHDIUeqkzEdlMZyTt+UNVTt
06HsWTfP8PkpiqIrvjjNzlDTPcExMQj2VI8oQ5EAa7PBhO62JUl7Fy9ps6nrCfz8M1C1AsLLnEXn
ApBsCzLiDc7K6Ppus3wpLWXQ3AnsQZ/eTfcwHleMpoCZAMym0xhmG2crEhpYPQXNzxZKAH69hF7E
ljiHbZdfRJsTNAYHc4AMYDMY2SzxdyJUFm5Vr8ekOkgGPj5Y+oTVHldSCVpXbBuuQBlgS1bLwrJe
llPe5iFH0UI1GzmLyVDykbpVyn/5GL/Vg9G5mYDS4ORbx+MRudRnDy1zNsGjzS9bOZxt4O9UewYb
fOBzFywWdb4LmvyLCkcBACnV4JIZ1iiU+tQFhSHkh+b+6soDSQM2RJOpjIXPkM/rIP6WuwZgVDsu
233JJq4ugGCZbcRrIH2yRnFPM4eCQm7neAeDsszxKcMLPPHRLjeBVvxexuQcZ2x4+kka7xmVdB+f
yJbb+GL4CqhZXeJH2CCjdRgzYq6MSqqSgsJkPiIpSkJv6R1baKYSXmXEI/CpmztLDSuTftnlN9FA
zOD5sSPletvHX48wk+FDDuJ0c8ZOyR/NIkUHLRgAmsmJSfPVy4rZMEAfzB9Z4MX41b77+ZBJYfYZ
fMe9P4srBE9es9Z73Wc4a+w9bvae8UgnOO6memkZasuVomUBoktwlS+sjEvLbwGnDBIPyB+Sx2M2
B1C2LNlhV7dRUrPTbWxV2aKxH+CB+xfjBt9BJmCagd0XoXs8iduD0Lb3lVZNx8WGVRFEk+saBaFH
ZD+/nHAjy8TW7mm8ADdufQwnOjWw19QB89mQ7kyrMqiW7izJ9KxqYmNMAu1D79Mse8OtkSGX/XcV
3gDKUYXr9m0CpcKzDHZLcHhEWbuNFrSvPOrsnnWehTbngGw3U1mPt/EX91+vKi7y3yybiKomwMt9
1t2TYJM1rKwFe1ZOqevOD0Eb5Qe3K0vHfeF6RwfzEo0saFPJH/7+TW2d0C4pIcYmzQ9sjlaGSR9e
GYrLZXzKQBoSbDDZMjpNYIYxk7z1CXDhrlj//QS0JakLAqCDsbDCUhyfPnD8lVrYertNp4OgVgIZ
sTQ2lBQVuPfnBrsLUZBkdp3+Umn3j122R85P18T3+WE30JNwdoYdKlEAHRL49Aayo+2A9S4tDFxv
nSN+YkjWAs4HAubrXISpq6dZ69fCim+sn4UIXLv6qZ2V2oagTih6kYrVQ6khFGxz1h0bGrScMjvo
dqEbU5gqAHMdAvrPyq+9/7d+zf/0UnLBdM47PQ0v5dZ6cTyGZhVuJbDEZLDdSKS9YwnF4N9eLYnO
JYyikI3ot4OVZpKwk+Z7CFqqdYDujdKrcJIZnwCN5FSEgEPt4ma2c8kDXHIJ+lmpZ24UC5jGFNF3
rrELLZWV3LTUiARiRW8H5Cz9yj/jdElq3lSW3jmlR9+46a6bGdPGb4f+pD0kmfHJ3SllTOtGh2LJ
PSCgKLNru5DRaP8VZjuZ+jjLMG5SxGgUz9Wr7xTw4sTLw42vNNL793zDscf8dbVGFJrrYvy8ctbB
qz8YCFOiwf9oPA/tcL5iURc1licsWiISeZPDF4lLSLUoGIYc4qIeEHqKUiGoZ6em4fg6od8wk+EI
fsA0ff+0XNHOnxNUT2scXQVU/Ywq60GfsEXtqfO6FuqEwgIKlT6yj7Nzs9H7Id7/YAT25I8CkKlb
SltDSqqP0/S3ndVkdP4umdQMGzcv7epVtUNxYSBA2JrfDB79wzNGgOdz/IdSMWu9trkGrSIzSwqH
zA9rE3FOOcUJuxr212qNn+9TeEJuiEVr8qUtq2hBltm0q5nFILEhKILH4hVYlzOtr+mFfYeF/yZl
3WjsATghdSMcR0/bUcSAcErozSYEPEeLwUVEM10w6FamOrSwc/Q12Uvij8rp3bXCtu38BI4I1r1x
b6KgtATyIK2F3h+o4I9eaRNrsAd0mLCeRX+/5ldMSCvXQndyDMD3dccZMbRXBEvEFRX4j2y1bRMD
JvoZ00vkUGAxmGxLkGhuWBa4duG4r6GvuMEldXkKPVf7Li6I/tgvMVqJZdvlWx7tcv7lC/S7842t
t8BfFSLiLflLR3/AvjZdp4p2kTuBQhZvH9Pv/oTfO1MEkSZMwz048nb84ijNMafKRfDIfwGonhB8
H370FHdBjOTTnfYsg65hiNDgIY9Ly8RbJZ6n0yOogyiCC0BGsCX5GaL/XELw5NZCigBDtEnokzU0
oWeDBUh9v7D+iG60A75w6KFWZ9LwD+fn4Jsrbo869xbfIUQYqgdCDuFz5Zgm+uQzJGQkFfaiezV5
abhXsaXQYW6w0cFdDa7Q5t3jG5Y/Amd0yr4Iyq73mXzAUYdE2wQh9NIxGNVGt0WyGqbg6+0unTsm
UbJW4Mnw5z/fGTVUX4YZ1n+2hjCg7RwX4t2+qYsuIkQLiaVICklTVfmntAHLwg2DbP4OEz2gXQou
4TAp6vbTw9S7gDPrZ2urmfIEAgZHIB6f3djFsKiZnxqpVpJH7wE7XYIyoHU/Q2jOh41DslFnQl5v
r70zqm6ialDiQQ/vyTZJ6T6I3uFys8QeqYl+REvIg1JF0jCIZ6alXAv5RH2BvEyct5hB8DbO135b
lUagw9o6Msf8ku+zkGlOE3cmfiyF0LXK9Kc0JFD3qTi0dBZV0JkemidjH++W06FMfngKbscTYYJv
0SG4cF2LHoU67Eg2/YYyLIxBvLijpRiJ9SZHXtUTHduJeHDIygNG8nBsPCIUYDKpmSpps9ESpDKj
qutbHvw+pz3DV52ESehdP5uO1LUwkfsGeN4fR8tiY/MNLJrEtyOpZG1Yvd8F3eF3ybF2Ace5twh9
+DlQcwziDIHvjcZQ4MPBdf3gzuU4sdDdSghnSiJ5DIjeExlsmCPBO0fSwpbDmV9rmcCjNzRWM2yf
0yAQeWQh3VqJ0Ibey1spKa/LaZEHRTWcfcO/FaEnGoXny7gKXavM8MHFGKVSQMbsD4HyIq0dPQ9+
MG7Jb/nHRF6sDOvUWrEoLkFo9PgvemlKAw3CUIQoB0zD+bswj+kG6vn0to2W9eiC1u7gSxVdexMB
40b6TrTLN5Xo/EabtS7pL0tZcuR05uRK0PqhWiKDLx9ytOn0gVdmktAcCbadxyZMDaGlSQXLLqQv
opZVzd25P6KpOinUenhxnLdjfXjDQVuQ5k/9VzUbA9mqvnum4XNu1CHwCfLB0FLpsMP5nhw/U7TW
Rt4hTmggVGg3osFyWVoAti7cZwKw9N1ACebZZfn1Yx8afGbss7FM8D4gyl5s6BsFOJdaET92Vw9L
XipcgquVAMoNa2Bt2PPRWa4Ceu+EBkmbr3uz2/xu5GWNzJu6u2gqojoTzBg5VeYM3FIT/GWUe4gc
MNs/N2RThqQDuq1D/XLl867LEhNjrGCrAUtWUTIq3eABIfr53NGPeM8hRF5qP11ugkpPzf3Z8hR1
6dPBPXB/uPWAKE3XrqJQgqOVyKXGAhlB7/GS5MqN+yyJFOcTVezPuK/+A1GUK6ZmTf5bnvUh53Pe
o88O+9MmW7s+6jbC7DjaCGDFpdXIHmX7j8nh1ErnKIPfd/d5MfFcf+HK3QzZhqakBgYM9ZSbhvXB
7ZhkXlxbu0WgYWfYDMVfqgfbAjGMC4XI8OlD+XO6BBfyxdgeh4kQx7EfvvxzyWzX7/OM8Ay87Lej
uYI3+shGTH5x/B0cG/OCE4srfdYZ+8ScaOLUTSv/P9NgqWFjT5tZFo6n9LtmjsTmXLgAkvvBp34w
pQ6/3JIv6314RUwJ8i/P06SD7QbAv8UCdFxT/Ms0CDbG+Q++/VUwgMNpw0KMHxQFyDIMJRMo5wnC
uczVn+56RM8zr4Un71OjGvQfBaCcQ7AGTHeBmYf/j1Jfk+sIzQDjOmrIAsKh20SW+ebHZGWjkjFa
NJN0ka7dQDbqSFf0QWuQqvz80IaBhSxq1PlouiEERPBabs7yGkOG3vyGw1a43s5dpS98Zx0taXlc
X1vPx6d297xBJ0DMI17V7PMZlDMtA9YXNCeFnTxvZ6zhz8z5kkOdqsTSCKzsxAlLkisaEKd2f8Vq
rskuBQXRXtxxejcQVJwn4znDsfr59ho5Wy8qsX6ius/Dn5dmaAhL1Bh8KeMlBcqRFqEvAZJFv7M0
i8KvnMdLEfSPTy7358X8wOwwL39EJmMy8BtkKWo/gb+9XVaRmTzJO03a5Ay62gbK5y9IdwseQ3Dn
Q574rBWfSZZG7BhczkWylTqSHQ9oWEKPZr8m30WHRWd0Llf4hZZwtZDc7tfyLkhI2WOU6y6l6y5b
lFjijT2Ax+cUkeZpxWUzsq1PqnKkr/v1Q30dmPlwQVklM9rFGxoXwj2mX3kRIEvXU8fWcZClPiLi
pATR/FRBQVH+W6Weua1OAtzQA/61ZaQKBzZMQM7MnxUpCqn4M8HZHoP+lGpGySwhv1v17p6yPFgw
Rwng7TwCl8nJt4a5iJDQa6LTq6iaZySUtwJRip3qIexDyExDFyLKE4qf03fcK+SNxyec3qJglzvH
TlDmh9IS+019AvmqW/z4Hj13gcJLXx2imN2guBfDnV3oTVIkJo110HLyb1xs5cP18+HUfFzKXk4L
B9yIHHx0VoIdE3CQDaIMP5mmQXH48SyqNjCwmkFMxXdQQHyurdv1B6YP9TgrHUM4ZBA1SzG2aq2h
OMSuLjb57icxQ1u9BjR824MoD3KaxozT6eFzM5d+ZiYdSpA5IkpMsNtiNmRCB/86peXJJ7BoCUUu
NKEe+40wLazZTRrLtxKiafucItgE3yNBuYTaii/087eULfO5/lyN5AbFUYoMMmYXI4KlpL1W9WTh
IqMXxgF84tzDQGJvhxuiM6kcfkWgaZ+208pezs/CGrcVQy5exg+VxMbAzYtG8e1nMCpCHpW755zb
3jkc3OV07lQClgK0DGvH5qaWBF8/dr0BqeafYUaWr4njEuF12Zn7flCrdKSJmMiwsade0NM0fgiY
+reZlmwL2k8RDhSDMQkEEvEXbbUDTVx1nN3/wjEWvVffzIjR9WFOoiXjkg9RK/nFe27Fd8zRGlJt
bNfqrL7O45QjRxRBUxw3j2CnRPEeoZa5R67gSgRR19wiD6xO/UdAkeCvk8FJBnDvQtZh/5mR8Y2y
00BYLLxXwOuI76UkRrYdeklbvTqEgoZAJHiO1s7Q2zN5JFi2WB+htQpP22hL3VMZK2meUSCrlYpw
AWvO0YDFS9e+THeq4EFf8gWu3DgSSCwkOWHDDGWFEESeLVOg5IkrZF8HgN8uTGzeJ6Lj6ZHs+Rc1
2PpR0jlpc4safWyr6XiwfBmzWLCuZ9Du2eDEXmcr2NG/tb90X9xAkWkUfzsjLw2LysiK9i80l417
2TXy7Y1vpsSvR2pbIzIrhlnEfL0f3vuIzMXT/KtinIXasN+b5I56dZ4jaT8DTDgzf4qgWN8KwGUu
v21FGNOlCzKTxVTNnve3LvWHP32TWFXO1RO24V1mTsBOj3dOdE6dlahL0tu4nZaLb63VtKlTpo2e
Lr2Jla7088E+fgLUeAT4NZ7lMiiuLsomttSuAL5OjHMpNsS0pAe30cL0ccthfIczk0p+3Ss0WnBB
fLL9qojBws7Gb36zuUhO9yfN0s2W8+vfPsbew3lKmt8TzbKBWh7+rJxb9bIzSFpjX8QlqXs6PB8o
2xDrl55MPOys3RNFzNS5TUWNsIpJhZJ3mbdDIaLZZPwj6TF4lXWGXOR91xx/DQLISfnX19sWybvw
2myFJsbAK3K1XWUwrEOhEwUbi9LZn+qTn49sO/5+vIitg3cf1zWzZ7esPp96jm2idskXB3jPJva3
KSkaFYn+sBv+egrSCkHss8IaT2yZMmWs/r2RbqQ4cc5yPCeOZcyHkQCUZ96oLY5hOnc1M/jmezKE
Q4BmxcUQu+q0RBLN8WTuACEqOvbdzYhFnpdnp2dsK2T6lAEccq8LYFXwt42NZ+0By4muLdYHJPDn
c94May9l7kfYmUEoiXtr9Homqxa1Qr9bVGdUwOWlZDEgbbyPxTk+dkfAXOpkFo3JKMks5KgxIFWV
ivhYyBXQlsFWGvMu64zKkEphqx1+BGksIZgkm0qZZz/bpAZXQkbZdvjE4qypf2GVCPw80Jyn4BeV
AQ27z1/5L7qQ0HSk4XNzK4kmZO2gWlmoZ73pjj1V1FvQfC9N6EtmMN+uxed+AK+cDDjxJaEtdcr9
10GC2BMZ6mDit0piKgvGk4Y60s2ex+5t25geuYYbL7sYGVDuTwUDnPHvOHPo4smriTAyVOUjcDrw
f5w+zUaCo513TAgoOzDAElPUJWYGdrTgi2y0eGKC/wFtQDLgEsnUXubmVDTphdRGmD4p1qntAxDC
bhm3SmNB0W2TURFFU+VqUACQ/WSDRjDjHbtfr/1rXREDbBIsY9sY3LLpj7jnaP7ax5knAzasKc/U
3QUrGn4arTWDXdSqFd1qnCMKq4hir980XaVYhFE8ffFKjKqK681RxVnpIVaT3ke3d1lZudLu4Pks
gi2ZqVCCd00pL99vVSaGmOnESWb6TG7Udh/SThqWzaMC26dgb1R2rOEHCmgZsYGyrkZcuePs12j/
OFVLl8BTWI288PM3oJNl831oXUbrcXUgOfc=
`protect end_protected

