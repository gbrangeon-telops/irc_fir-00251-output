

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Hz4PNZqDQYlRQ+ken68CUlKtwl5bD3KVcGYwK7pLDyYBwi6Th9L/PQr7ts5tJoXAIQRYcIzRxOvE
bOvIjO60PA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
GP7r+Hw/Nq0CwA10fCvNkrkcgK45iHUPRmPqoCkPDKd3ozfduaGFS4NbQcQDFEPry0eRmQ2gSn3i
AGkmBiS/ZMkSitJxD/EIgYbO/fqPeNo/xyESKAW2O+T1ZwGwXyv6qMAp2gFqycRAbj6T5U/FUq52
EYpn3NB0sMc8yOEFyQo=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
le8HFUmlytAxiraEF0H5rT3qqsng3b8xZZHcvlli3mx0SdV7s39NBBuklCsi2z+U5UKSzgnk8WIo
w7XOgbkBH4I5bMmtC280eEWQOIcj1GSezKn8Kq725OUTUl7WIOM9hdaAEgsyYV4aegR9ufM3pfv5
jM49vFUeG7XEd7xqdKUxYcrZmsZ8CqQuOZKMv7+xnku0k9eaKv42hAQ7cL1uIXuIFvzDlZHyC8MD
e2+jTkJtzyJMk7U2Hncf7jaM/O2gSIFGoRR2sNNwVB0ATLYzGBnoP+wY1MWKJdSoIbDQ5r0792eb
YO5yRbe6PhUe2+UdG6sNzgiR0viGJQ6R/9i02A==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
tSJEOPsqlnARL2Dz0wpm4XWyg0nGSs+Wnp+fpstkJG7juRdPH6snLi4H3YFLGcOIteaUd6+0+nV0
HNDEDrgudSIwom4ffSyyotXElk+U/5goIr091+0B19LyBlVHPMfovruJJsH5yPOjkIUbE3z//OG/
9D90RTj2hDW4+5DRikw=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Y2U+pnaPqDjEYN9Ag4nM7UfxJ44UWPvMFi6W/IpytPtcFc+Gta7bvyNellM8zINHBtaT4/XvwpGs
zz9LduYm/i37u/eaLh4notjKL1KlEzSl/RQQCOAWEkJvBF59EPqbeUalx4NMTEi6gApYczcwU5ry
jjndsvqks3Obkc3R6uXlQHIzKbPFQM2kj8SV74srGUscAjTY98txOVHFhIk/okWPW2x7ScPBZlnH
/p6enNTFgNVy7YICPLQQ9SjExe9hKly0/QrbtcXPdI2+m7HVD28iWrn6JNqPDPmkYTv4lqGhGruw
jT2AigpLW8vV0cP+HITHbLQV7l7eN+9WNmGRNA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 126368)
`protect data_block
/y6HVwbfVC1fGOEVEYXRlgY41rqBwBhAbpVaaCUI6pkuUrGqdAjDYsL+UDLrYibjyX25uJwXuWjz
YB1+hniS2Ns4ertsCKH3LqJ++xgD2eq2/KbSQuqt4yQIWmSCbstIpKT2QVbGBIUbiOIA+wMT42pJ
PkzDl2CeYksfNh6i29iFOpctCPvDLYK0/DOqNwGX2RXxOIdeb2/h0T2De3K0ZgGKAb0RUVWQ/dWS
ePkNAb2u+0ppRm/nnUwYUQzRylaCGg+GTnDrinqGBXStMvqAvpvN5FMj7zsL7XB2I4FJ32FxVvcC
1Zo0EQg+dkLoPbIeTW5wjvaARfkaZdD6yalPBtoyxGlY4gS954dMX5mAx2m4m5pdoJjyKR0taYpE
ZopdAsCuOArQw6Cn6ma57Ej4F7wz+TVGD91/MrygAzWFmo4nk19Mj7/LrYNmtu6vXuy1hGv6AeQo
RZAB0Mmg1PYJ7krfTIxYFvJSiz0Y+xesdh354CnZFb/hOD90v0cdAahzDlaaNlg0IiVCasTeskTi
TyS0tyYDDBizK+l/EekqES0HrajS5qvOMxftCFDaPq0NhLvXfGov8UebYACM9NEMUle5L0YWmPXI
O+S1T66zZF6EZ6A00Xr9FRo33jGwHdnoVf81uE+0QDPctvdD5HAGotteXlTRK6kC46UR6UOGXDVw
4P6HsUzkbSyAo0LkIiGKHXJAeYft5yTWHfoRLMrFnUoBjz7xvA4QgZVhhe0AiW6mYXj5i1NYBxBg
5uZclsQfPLN/Y3mOAWc339g94ll9B0pfxPuVVqzVivsB3uqkZDrmm5bzCtnCXrdbIR0PVz2N3cBn
sL1YTrMwSsCPuHKuHv4dyGCLIiSrG531BSta5HvfnckJ7eE8XhT/W81blfkyDGzDFiHhBT6FMNlu
hsjF7uWZ9tpVE3tZXVSLmYGs/0xoS6QvXbjvLNOgNMU0fOfunslXJfunfRfHEMrSshhm20J/Ljdu
v0pKaD0R/c2AQ3HsLKupp504334gyOgWxPXpnFTf+kCjw22DPtCeYWTxZ9Ofo0y5EcixXL1c1Brf
Mx1c1/UtDB6rS6nHXzu5JCU9SE1QsDrKK7vOJ1shNcRKdkow7iAZ4k4hjRWWCfOZI6eATPE11VOP
mw4IbaZ+oeQbjM8UTAKkpQMYxx/80MAAibTeM89OC2jz2qVakm/6Byo6aoyOlFWRPKK2WvfBDK4W
9xQo+WQKEBMKIOG4SymI85w7spbwe9HTvSOlYmB8z5AhpfL6YKiZqpz31t+AyRpfq9qP1hvMfId1
f3/TGnqIa+EcaVxSfzHk80qjHct7betcXddgsQNwBiVlgQem0ORpIzUMdH6jfbFO2W4Wa0XbC/W8
oH/HEViVPv7QexEWdBpcc57ONtFqreap3Qp9jjythcEv4V2jOUJy2gx+3m0JIlA6crszvL0BEAsq
/rSgDT7bOgg9gBbXJ0qg+gq5NY81BiQrtWpvcgE30M8vmdIyCIzxav22qIVXmjJ1Oct1YvEaYNLF
SkJlLuKs81kqaE+WhyNvTaQXnG+WmnVpit2LOpqrlus+HUkTkbEf91t8f13ZQ+qdsHBrFEzJOPsK
vc/R4d4QC1keunCMemsDtFtdFX3BzYW88rnWPbWwoeB5hT8KfwRiuAwaiWoB8maCP9SivbIgR6H0
dwZL5+glZCgGz6jsD5nCbOMelpjldxYFK/6OyFPLkvcfEEEQOi54Fe16aisS4jwPD9MD606LIrx8
tVAfGGkYbnl/DSV7vGYJBeO+DLMhbMfOyI/oTVeaZU3n2/J8EO//zAorvmdqB8GcTmxZJXY2HC6K
aohH6VHUi7y7O7TcPrduP6A7FTnXLb/QdCQk5ruafrFiQEmgvY9bXNpRIITAS5Buf/42jowOoSQH
QtxnsST3rixlHUM3tSs04JXOzrRZAlqUWjGSh3I7iCI/TKA3AbzNtWdhL7Cb+qeEBAky+KASgw1r
PnXC3WWcr+m+r5YNQo3gBcp/VQRaORK6glXha6ZH6LkcNgs2uD+xFvQ9pDhoiFm6qKp96TA6ieWP
EN8NyV6xt24/bJj5K27aVvlzMozZVstWKvn5ftM/yQrRGc9LwucCYHpCkVS7Ww3NUrPkJ2CMMNig
NFDh/Bedoa1r1GeTw44evHFYETOpOMTPjM1E6f1FfTKhoEAZqqt0I2cRVmAQUcoV8eZrSqSBy/Jk
qlGwqjzC9oIU4ohkvsrgqzfOV83ZJGMTHuWUO/rk3CML1bwFvPCjUGYICX3E74JjyU3LHtAB0c2i
9NY1rIw+K5UPBkxmJZOGBwQZScMx2e8Ocgfi0KmfyI8UH7VGajYv4EFKsXCSykdZE+2DzXmpddQb
ojEKmZqxMat8R7uLgdEv0+V3SjsjKu+MQH5XEJTm1kSlWidfXUnBfM0QxvECBUqi3pcVbN29wIRh
e923Fqqh0Y3EihV8vr8jdBmLdZu+R/DYY/1P5h9imucYxV+SwWY++Y5NvrZPHcjstwKb6ibGeHaD
wKPuCh4RG5KsFs5+5L9bzyfElAx5XwN3SMymmeZDux8lT/kypMbdzhMpUnzVBZhfqcffHKw+f7PP
DwyuLY4GaxLHaqTfY6CtEMSIoEeikXBXbfJHMnbMIvlkytm9lr5hkaawJi6DnffTNWznlE0v3tw3
betNqcZrLzZ67GATYEM0NBrMxJo7b+oaDMDYSkkLfU9KKdI/mfBUJyL+P+ScNN8leAjVzk93Qto7
urxhjwpKL92L14X/yl8KFoxyOYXeO8lVrV0xQoVaKhjKYrVwSVvfQe7wIRtTbjptIoW/C4uazSKc
/7SwFMqhJtrRRLJswjqtu/F7hJ3jILsWFFnnrf1lS3N17NYvTC/S5mvXpNUwhMGmN9LchQRPPVkO
72l22J6KLLNSr47AceGkb3kwFBzlo1eWj0HBhmmeIycP+Bi6QUacg9F49qSnUY8CF3J78lMSbnm/
sWq2ZH8EX7n2x7raRh9tgAwEs0owSqPZX8UQKGBOeU1yOAWPLwPp3WpNcImCyhNbxt7eyCMbIxoc
l4qSGp/nE/LCo7iW/RrXQsu68lPkGYBKWehLaA1jN1xuAqzY3QKBarf9+SUJm7Tv7TaBa7OL3RgY
igrzP32D1hUuafskvLWVdj/NiFuojHbDqOtRcn1DMZH1Yzj3IfhlwkUKLtsc1w7JrX14KEybxaqW
VNGVVpBbn4NCFPOgPI+3gg4Jji+omLSge1gbXR3JIdsfFAFRYCzFvQu1Xhmt/7xDvCVJ+1OrnbnH
VPtutlwW8QHKTDFx5O9ZmCAo2JZ0vlUafec2KQEvjQt4VtFvGSwCrpFu6NBUDcyOyaGPACfMdy5X
mLxV8j9ShHTmI0pnlroVeduiSPdo90ASq2jK1h1rDXMH7qOFfGuRaB6+r56TPsWH1ZAwbr2nT4zn
LkKUB0V8qsOQ9jWQFWP4nzx2uQusemP0UYQPF/f/qjwk9Flet4+2Xsq1PE4+JP96S6t/gHdgukV9
+u5ozvFKhl02DQ80QuunGq3HQdPsoy1NuSRcnt0wnJ8TOCoSxrqPwUgjQoZIYGFdcAeggpT8XHm+
gbF6ojAyCrzhXV8yWP/G/lFnf1YPny3UI7DpV9eFOOQKlqR5WmG7POY+YFNHPRxRvP3omhgxWy9H
j31eaU/9mujKa933VnVd2YXlpXKml+9+bTW7aJKUwKgApBVDFbdkmH8BIGQxyhB+lkzzuge4rOHi
Ioye0pVdywbGvWJ+U6pYXabqBNT1X7EqzGgGVVpBJNhbEyKFoiSXMM5sj5qNBhomX9zANPS84/+x
ef+aumTm5t1rf4igZl8BVNIM/i1J2AoPkl4rstVslnkRVySDlxLXWH2+/Unb0jLq+XtYNmgW31AV
ORi7kHrTC98Jg0HBW2JbK1SHpxMHwRJCZrhsfW1p0r/8S2zrYtSLLFIDLJ2NC3YXdTdMdHtkcsZA
md3/YSvS/JHwpXLEsAK87frzp0ji8q31p7gvsZ5Ga3UY2WJcrUvMOCf8uUps5TkNbhv47/Uw8acC
yLfLcLeGTwFh+y2byi8BIbG63K1sHFyvVOtd2dYc+Q7xmzKJgiWlz3xiqnVqtaz49oq1qGb0jVV8
yA0o6GgrxQ0JNfvFmI9AAoaPlpJOqlDCVLSqJPg7ly/ydnYybsAtU8J+ngSKEc61xgxMt6YwjT0X
an5XUwwqq2+0yqxaUHdLFAkZXOiRZTjL/+x738adgUI/ZUbUpkR9q41c6K+9O86MuUz3EGIOYUG+
wW0vP91zzo0eKDhAArHYzhoDm9QCfALdEezphEsAjd6ZhY530FaGcDwyLgP9uzLC89+qJBDaXwKI
9vRQha4oWCQIjO6RqQxewtrVQvU9GX9Lfkxkt41D0AP3xl8+0KlQksuX1mARQD9V9J0i2c+8RX+t
0MEbQFeH+lEB4C8ikBu8vsU9wSP6j/vBzn8frnezrW84rVYfHtbe+Npbilm/swLRNe+bPw0wUSKM
zClwZ7vagw6oD0y7DzGAbdnRATmXrqIqVEaSdBGHbSDI1fPW4akHXPoE9NC+VSL+rZTbKF+1m+g9
87KWsaFV5YpM7MOdd+XTRDNP8ZjvtLQ13K2jI9E79cJg8S+AXGvQ7lzPiMgnqUtDh+NQ9OF7qLhM
AONLbhHyC06/UvPDC0NRNcuQ7Tb+bU49+e+mZKWQ9gNn+PiyaiWFcyxr0q4zxIm/hv3RwNqtn5Kh
4tHiuivupRPbYlgetgf9InPlFazXezMDoRQga27YizcOug+NMTSRbS3KS/2ZhVd/LZ5A272OA7qF
fJKdFJWG56sKhEDPDNDFfF8cV061FcxIXMUYx6lu8uoZBwx8FLa35nxfXS0/lCkswXoAe7eaoItx
6uGmhzPUNXjoY65gbyXfHTDvU1A3xxoHtlgeA85w4Y5S2qaGL7xo/9vzHB3Uk2HrAmNWxB4XfYSM
H2wrshnLSmNXJLiicP9vGmSuRUq+0mYlQVKWeAv74wM8LEfS1WbElQTb72Fb3TqBNurWsmWgRETU
7EbCmemBcmQO8yVijQdZm0rqHY+4tc5GKENA6rkfHI0R91SVdD4gX4x/RGJQHEgE/5cOCdSQfh39
iSoX0hHjfr9IsJE3MC5jC/tcEWiIJudJ6xNW7BCfzcU4ndb0iJqbZxgs5KIfA5oGbRTjzeQVrzrW
5aM6CQiAjDMOTKPoJvcWaWzIVETg1ClmsArUQ7kn303oJalaXCeZr6ahhZB3OlkBnw1XFeNVT1Yv
vbOr7FTXOpKctjnq8bZ04s7OSKf6PsA3CuOozAHcHaXPCxFZG3DUYmWWlrWmZHSmcS+ONXERqEFI
wHGDawnVj2aLJbnSAgZZzAKJW7hgsmx2YAtnk9zA2vNgxECvhieDXFoV0bGhLT0XJAbWSuVsSJRz
QuBj1FogvjffVnais+iWmJDJEU66v9N/EtN9CGM6jMICKOfoUTd+M/xQAsipoCVuaK3FjcYZnRPI
CmdnRmwfqQVhaxPYTKxlF/wlEtksbyk+BXrcMYrxLLnVp3J+CJn/ZgpgZkCvNtmb4/6PWmQaQdfl
bkvTZMXV8BJquc+DpKWOYMFx5BcLZqq9HNfGgFNAGjuPzL1w+txYm5W/Q2jvQBexMkM9U0QvS6Yq
6VbB0KoJlmoN/HrrlKChcvV8LwZzU9XmI32L1YmKwBuCmAn1rp+XhPIZ0cwEz0TT67SB0z0DQnjQ
uPXeAYMxqqMWNv0eUQZX41MHTdmYh4XPFb0YRPc2j1zPxHyBVNU1Nef0Ac9bnIXE1IZtHN5/iau7
/RpOYLkmYG7Pp4ewxBAzsYoCZEx3g3ItWBgqpwOWvAaZ07/BO6agWjqhUeyOyNzevS2eJMIsv6Ks
v0d2vO/BSRD7hv0+eDFFCiHS4eb5nHo0wviD2Xq/j8gyzOtFq3hkEJCbdk9KpttvO9TGHL0+p8eF
sNZxG1By1a/Bq6mTiTedlZnBnZl+TZANXpKEnyyeD9GyWEKCgajn3dEqDjD11+BwaGYiqkBrpxjK
1LrKpdDxP10wWbHCi9bBOnjVN06uv1x/tEZGZoB7l8dYnWG0Ii8n21dHFMBHK+GidI0a5xUkdiEz
4/+tJZ65YwgePKdKygd2AnX7keFK95JDaFU8ILdFTjLhgjPWvj+TQrvTCdpeYFU/jrtcTcef42An
SQ/jMm76SZnn2HiQZk//s0C/C0pJO2Jj2HDBosvqF3upOI6A3CgVrIbSS7Mrb1PnYxou3B4q/2yE
H7+T8N3KoelELYMNiFa/nzLpyPttBw1U9w907+ikEmqundVRJujxpAlGnXMU8kBwCQjLd20xI34f
KHw9ehE9m3EaDmd4dKjejjxiaHaGO0AEfkX7GNP8HTLeeXPlJgxxTHpURvvRxK0+wBkPb2nFFoOo
f0acIVjLVu4xRFQNEFfJLXVYaoRrc9rVaZtu+N/OwMkGxd3plFvR/uz/qNwjzFrb562v/pIpFGXY
io5zxQwie4q/XbqCGDePv8NNGIa4q/X1/AzsSHSirqROBSFueLJoksyEwFxn5gVlyGOWyZkh6du/
VqOMoRjYEt8uu7oo1HspEMAvJ2j0XMrcTfNRdXj4h1FSl9gIdg3qLPjWSaK3QOVwY5nElNSmrJbO
/kmTAleLkdLpnC61ld6BH2iS2dPbIsnCx/JQ38y7yWg0XPdtPL00Z8UnblXlEFseHyziDmnkgKBV
UiZuwDh9DS09gRSGeARuvDqQswk4fTMN0+6s75XXvTKUS66dwJGaT/jRzk2bILJo7uY4o5X5iOkJ
+zMCbVK0fZmr2v6j+gvwpSECMf9OCZmRqMsjiXhFwBsBAuHZj5UatLAhn5+uGi2452CiZ7AAH3Vh
dKEjbm/S/MN1W3obOER/v0Mj6GbJSIBmb9oEQRfGqJfaIz86s1Ac6yj14vT5WHq5IqTFnS6PoQxy
jcs0YUc44U8fWcuxSGuYJJsF8LkKFhBPamWw10E/ae0XP68aveSr9dhFj1oN7WQ6K/NoPsuAejOU
W3aBSSA1IOLmWWX4eVCuf7A2pI7xvuQe6XD7PU6VKIwo7xlkNnLedZ89XWZEJy1N5QajRYyiYGnB
Ef32vk6bpNfKPVZVOeuSaPn/4MPAZrgnx7ZVVncdhwUpQ7gdWvDtor/BvksRjqjSW+U3LSupGSuQ
sY0rTky1ScKC0/M3zaRN/eEGNLGL8e/6scFDRj4d388Nl6cooo/9Px7AmLjo3feCRCL2WIPJLs/M
ixUCFTAWKfte52lNaCt+uJJRWAi59jm7eww42GH15Dt0eBIoG3D2sCyvcqV91JoF2VfusBERGlcN
QVkqQvhni6Yfw6ogoZ/nKPSrH4VG6gEeayxcq2c9aolhicJe/GXNpj5ZXI5sIHzxbQwP9lq7xBmp
D9FVEnU563tNxb6j8t/ikvbPggxmYXWNLHU4HTiG8ggSgBattLG2XfB0nr3lKV/HHH3IngTHVy9X
eg1VacgeYDV26t+oBxZC/qMQP3dFludeItXQFuU5qaFICD+bsHA5nF0WfNiSW60CK/m1NgUNDWrG
3dxc9x8DZoqm7NmHjKiGiRUYGgkd4W/9YjF3QsBgUz9ueQtrwTvg5X7FNP65D0uLw1bcJezcYPnk
WEAc7MNGSSW7BdqbrqeQxYyVJNAUP2QlF44CFGK2qNM53875tKmv/TnEZeE9qrmz7SkRN1l79f/Y
ONePiE4P1f09vW07zI6xXndCpGVKrOexpRQRVFKmy3nx5prkUC+VVDUQgoYJhdMbyy90rFUHW8mf
3c/Tad2FZpzPJQ0+02kMPGwjGtk3LehbaGPZuNAWtyxDljC1M280/WSsiGaXZ+by0HhU/RLoSi/V
gk2NEIDhRpkQJJzpHFSR9GueEec5kgP/LwxE+1xz/e+igfSMhTedInE+HT4jQGpcKNmtyzLIm77y
PIMLc+B0r5y4YpTnqfG9rkpO7m69hYO3LBREsgDtDR7B2IIh3U3UpPjU1K8w7rUopAJq9AxJVazI
YDIDZeS4rpnwGfdwfyNSfak/6OpXaveSLEHzaGAIgO8/KTMLwwH6DXT0qr9xuTzze1+qzE1bRpdD
oMyhQfwNnmKYqekXdgkUZ8Hzt0dzuAnilbTGwsT5vQjBNiLO4uo+3yaY+vX10QCRhIVpIQ0ooFqU
91YD4ko0Z9ZggnY1qC789oBg62mYw37fQSvgP8DYXZE4Ju/U3NX9EOd5e7mDxoGbhzhH/xW+p9qd
HHybeC4kgtDW3tHf2s3LTxM6nRvNUbzUh3TKo5NVzLXJnZvctPhIkADzj3SwfHlghEnDzsK1zFhZ
Ly8192hTk65dkB7lufqU5QMKPCpeZfqSW76+KgjGgH+01Oq0dbLgcbEZPoYLqE5Rp+TOTUqmdpcj
VVeiWt3ZMji4MHeqW1rePaPMlZ09K0VhG861yZ7EEKtzADoYfXI4HLJyjTAUiv6cs+O3YcPm6Es2
T8md3ZNIzIRPHLs7XMEej/Z1jvaanaLwTxFfTslNxMNHflKaDwogbo7AaVIFZau6MDsWyT4j9pZm
dxJe8I6X9P3sF2S9aF3KNBqdqq6YNdXqmKs2WaqconGu+t+CEuNZGZn+DEaU0fsafbkJPJt5T4qr
MKfPDKlIU7oj1fH5GnnQ+vEp4SlZN3iH9r8cH4ibDWpp4HjnLIJ3Xab31g+FhGN/O3v29mKtu8vo
2Mg+71nMWYIyi3kHaAMnwInjGTV/uBvHUOE0AG5VjmzUs7/BBuiOlXcQzIFwr5W7FRTud1wVYLN+
JRNU/hqi6T7xZGYNf2X3c2D+U8jJXqAF1Tsg7EhJWcOXvCZUrNl1cM9wk8BNjCiTdGI9qDYCV9SE
/D1ujnaoCEJYkYKdec8Za0UR6jyWBOrCQbvUg0PR0RxEKJSIaZ4Y8MGBZ6jjukiJx6CAy/Iy6sl+
xSGCJ5yEBuLIK6Q3qK25rTR9PL2vdfk77nQrYZxEit31wDUQrT0EbBjrGfJLpAGVWwXhAqdfCCIJ
k5gPY6uHflIyRmJprU5WGC+xf3BENQ9uIMOoUVmfXuL+ratzG5a9DVtqwy055fwUa2TVPgWFW87G
dsv28pbmKW4nocTvk7Ph2VF9GvppEQZr5lrVr3tiiZXrbxZQ8k+SQO/q6WcC46vg6XJ8QX5t4MRI
SV1PHL4W/4hz0Xu/a5HTi6PVCY7wXFryTD9Ev3YzgJc8TF8SIU04LeDB43Jo7zUUWdKSS2jmSLaX
DlpkWw1Ef5C504RA5O32QOYzSQoDyDHC9aw9r6sKk5l3G1f1dV0SzIjMNcyZ/8KqDBZ9oHTi1ebh
vPb9if7ll+C6jFTgMV0rfBlVI//NlrvehuzOtUDyn9Cd0/7XG2C6qgSEctF3a/DkJ6FaHcjPbxH9
Ld5n8ACPLDyxw3VDhbE+k4eA9mPrEbA+tiG47ACnD9NRKw54fqANlGNeb4l4qGYu8KRL+YJmJV1g
wx0vVfZuiEA0KqU17TybUsWliQI1+ASSGFsNRPi1hp8p7vfl18/y6dt3Tsm5hl5aDQ3U407Tgg3s
/BMGRxlm+QSQEqzocVPRZ9fqqCm6GYfd47k6z2DzCeay+vEA0KDK5u28fb6eZAdjm5Efs6Oi5MIj
2qFCCF2WrLp/+FzqAABSYENomD2AB/bJNx9bspuR8txtNAVR8OGHlD8sJvqPOyb+wRbQqxBH+o+g
sJgMNVhdgva/2KUg1ety+fOd/JAwn5Hf8xKKS78u4egO0Q6eti1VoQ8VVVS0HTl2JodkTOVCIrIP
ugsZ+1WRc109gGkuw77Ow4ZZnMxA1KpBujhN9Mg0QmyscOUg9D3mEWSFuPeBPAobgvgYUE/JyZLE
BWS/lRVU2jbtiqbBNG8iKfaRZiSWM9Zf3D1JqW6ze508LJRVfIbaP5uUHxigUAZQIQlrT+S8AKP1
zuJnboo/mKRK+Fa4notH44XeK+BcuM+GK9hkLv9aUH62boQU0n7tiMO8ss8LQC78vu/gRD8o/RNe
lsqGL2lyV+WOTcWe0AV1KomMpgivQUDlJYVEtwt8e7upC9Qe8SMPMerhIKwFIrenDL2JBDt1+C+l
3Xn9rhnarNXK41Pteg4DATN2cTVptyRgqHCLCnL/UzxsLJJdYGeJrYUK6WbXXxQoE1mj1Z6Dvkih
tyy+XjWUlZGOine7+Sa801G6AqBX6GOun+t2o+n1EV0UChgpSNgxr9DNDITBro8v94WaXCvPNPCy
ZwWHzTFnSXY+ndL4ArPWyKPT4w4UEORgTNR4ilGOZB+yerpvpfqprJSCcaPUJxYivkwyV5hotgB+
fiYmb1EGGFhWJtRC9spedOdUd+CHp7AdnjQmvAxv4U3KoubJWJpIQGRn7Q7ifXPk1KOLD6GqPOq8
OzwzWQxg33yGnwkFdVaaEZNnJsLFt9xkq1mWGoHT5JKqJf0of8bmetw6lbm9rJxdkFbZMk5w2rJe
sIt6dxPFpT+/8YdOEl+Pg9F/OEMUm0oniDxkVVrefBCt+kS0PLQaYmzumBTNNF7wDMXooeUxGY+H
xmXEVtutFk2tmpdT7inX8iOgo6ksoFt2pV+WtPJMgb7ahamFklEW99ZX8E47MWhQTCcQ5qEvpGew
EK3cWL+UEqv6G5LFhuPBRqRcHdGIDKQYqdw7I2pDLDrJlncXFuh0pIenFp2F48hpMdCo1QR9XlHP
AfRQhT2Ally7zdXjuWh8TFi5EpaAs3ty/Zrbtsac8nspsbEUjk0sl/1vAtF1I0rlANMeZU78s+z5
5QqFuFuNF9haxCeOKUs0uQP7rdRBYXH7IVS5IMbnyXOgYtGZayw+DjPnCscSFaCZaCj1PJJ4TS82
mREmhViqUevJfos32dhQUrNykGxdO8kj/DB8jKjBpB6RoBM4Li7zSfkBH/pKGfw5/rzbhhC8l11t
LMTlJVbrkH57fE7U+9O6gzG2XRzANf9jTVJoZlJOApkPA6HwH9OCpIbFoj918d3PZ60XYaVMKun5
fC6JKbtLYgsWyMMXElrnLQ/kDMTUWHmYvxHu23iXKZ6HvisyIax4o5fktOuBiIaocamLm309nagK
SH4C2aX9MmzA4ZTW2Kt1V9sp2rDOVqN2pruQkzbgmqleEGDTIRLTg7vHw533pdDwAP3+cKojbG+4
FlZPE39aM2E15XXAwliC6vgBbRPFC45312oM2LDgbb/kWNdQWngBMMltRmwu9dZ4qRPEOvcj/3/c
RpOUFrBZQu/jiAx8eOpRKPFfx0KMiQTGL1g9L1FvRZsZs2y/TgzYAN8lY7A1H1Es4NZrB6bO9+VP
l93uDiF4eXc0VBjJz+iDikVITBdKelrzDDsVH9H/DR5CYLPlknueP0PwMX/RrQYjZBYTzA877b3G
NuHmhdtlIerQw3T17BbMWjwohaYavFQdXxRYjxJnf4xhBNnenBqEtCYHVYSXhJDon+eiQT7mnFCK
RCtYkvllFHoo/e1LRLUnL+x51+6MwYHmIry8/RbUtdAuERUunczmSF04OB5dpIujwAhyLIhUX9F+
aMKhDasvpOZmVZtkKSip4Hm1SlzVnisevJgwepaO3GG93sm6omMpIQV2ppQNeDDXQIVCV8GVaz1h
QBS2l0dfPXi1IN9/RbDIE115+vP36HaDtqqeD8iYEtglxyAYbLNXPn2KwJTIaUHLFq9svS/TYYXx
HLyqqQ3QskYdCDOkdhe3x+de6COHQpux14QHBqjOmRJr4NZJfYV/OA/5nciELjXmwAm7ttvZKOj8
WRCpA9YnNXB0cfQKGWtrtyXt0RIC4u/OLX4V89RiwwlenPIuVBHSJivktZrf35v6sVOZVJUFbA5R
KmdfE7wkwv931DqaaoU/xmg2W9tFnodEByPTaMBtesyQkb4K2mpiYs1E27uJm4im0B6HKy/qdCpr
tF0wVNFndLYMncqV2U67hAu5B1jLVgCNrbNx87yvPNr5UiuOgWjO4nyz05qkI+VPSx3cUNoe56jP
FD9dTwb+MhKMu9toVr3a2U9r5XOiXT0HRMFA4sV491fBVXZOf3ythe/e8c2zm01u6HV+lcwbzFC/
gwmN7r6iQwugFElBRMJQMp9WmUv60VX+RwjQbfjj2XqPdAaMwbOabiP0beGYC4YT2d6hf0keO1oP
QJ7zBdtjD9LHFcksjfXND//vC/6/YAkpGMUBSnkIeLnX81eDs8++OfTP0+nZs+ym1jDtuHGtKHHl
/IlxibG/23i22YoN2aZdmY68MU176OQyg3RtkMB3z1STVFLf7o97+bO6GiUBbvFZG+KH3ecyh6Qh
U+nZ/SMPBpFio0yfQPu68r4rO7XcGqbPJnUD6K5+M01BCJqeX37IzPloPTESAPKDqEvfqbO3DVZb
c4hhv8MKemeFesTGyMNOiSIfCKuTev0Cgtsn/W+IuylkCAkOHTkMPW7kfVUKLAOXDNAQA/Lnb4Fa
6gj4DSksTrExFfoaOMlbsNPrBVcdwVBIsOzQ+nWMt1Tp1SH7aUCGZ94kYMZCWFaMEI00HXMke2dT
NJvnZQHctskcnOaOxRmL1zPYc1hM5P1VOaZ4yo0trrjQIMyxH+Na60b4a2I+4CjjbNFbBek0qKNI
uovRuvdKGm8IMgPzNcjQbsa/lJaXU3Y8kpBsSN77DqA2P0oo1lEwNwb6UjpkaNyExtVWhAgzfEOa
Msdsreeo73ayJjA/8CyvDZjlxU+bhmaCXg9rxJUiRcixsTxqp+/LpmjShQMJu3ZuMjeJwPB+obrU
xHrcbgP2ubg97Zg3EP7t4UxMG6pxkOqJAFcSahUg9FXvNlM59zNuTjCKf3wkxD51QYKSeyFy47MK
Sfe0f1X0bJncbYdhO6BqErVBdJ+bHszhV/bRVBbwnwfsOsz/7b9qzBHEFFJMrR3+2CqOdyHmg0H6
M6jX0qT/1RzOUI3aKVkqV4EmAAKdrZhyKEGbRstFxZSQe0crCSBRiaYHg6rAOJ3pCWn4KqgHVI0f
mfKePhWohBRJ90TEG1Aw1Fo8GrNqoJyiWhs6DHrcsfW3G9du+KNbIs/W4iSzDg+YJnT4UoNd9a3O
EYepDEfeRq7A5ShxzPjrZwJzUtRcbMtmp4aU04r00GmuwM3C4XMe3/hfv7fARIWxSBIZt9r+FK+v
WmtUr3/iyqxHD5wepRgwEZbcIBcBITTkWt5mqp+Lc/wd7oS9bDThBpEh1t5dSbXOUCFkEQJxXR+H
1t1IzBI9a/kBGrhS7x6h18G3B95WpuYD+2tRY7olS00pbhEhNLIslEKt+0BDcQG6D8mk+RWutl2J
glebDTVghgNz+VYwl8BF/r+gMLb53nfDTqPfJKZXGqU8GWTgoICTpTrI5kujSwmF6pdlj89J96n2
i/FCkVOZ9FnjzaXE7cWdfKgnXH7fuzh7xwm7Vt0fi/1l8ch3fCmx1w+6ZcXIFESD3anf+2pagGRD
OT0x9hPUo3yBAJa+TFpBnacx3rteYmn7vKGVFymqtPDGSfU0x6H8sZq15NdRoO/7cvpjMIJ1Mvlb
I0fpA5on3qCPz16pTy+2zuvoMYEVcOLHeHvOPfPRF7WEUq/r4MPhjy+9tUYZyhzarT10/ki3qb3O
/TDyO3Uyqg6s5wqeiYeE/iJxovEjORblyw+bM4D58DEXiUCsPoYtqCvGYbsGEZYdE1ZbUKo21xdb
6j3B+6tPOuxOgO65t7bUWEaHOLtI+4Kdrz6k7O2mfugK9zTXXb4DjYsThtHuLhn8cmOCzVEUfeEL
4fT6gECEGJolRgi/ap+m0+ngtp0LSUSIQkA6dNDqyVe/KCFBjBOWZzntnkVjIUvqaaWc7vvV4nO9
Gd5itxF524txi3tu9bsLcVoga9tyHM/zdzAAt5gVj1w1dshPVJnVDsk8BKxhu5NN2Pvc5WoMajas
UasLYwHMwapTTaaSeRVbelZxRNOyb9Odr7VKok+u4JL6Trv/ssKrdAAEyM4iksbxchlMQIxGpC2g
wbVpqcQX6nh4Jyq5bTkMc15nv0Rk/Plpg3aHzSNLNW9IlOxC2O6LnNxDe/s+0CM8Cz16O2KM37+X
u6xYwcP97HFw94HEOnFowJxWH6F38Sx40+Mp4DrQRpF2HCqn3+n6yClmtzx84pS46+zKNWQYRlSy
lNo7JMBNV1nqRpl/Zy1JdDi/lhpSDcVr+arl1g81Yh1VRdBsQKA0wUv7vr+cxmB75iRlExW1+fqy
fQYpxY3IvWtWjq9TIyPZdkLNmlIioIAI9Gf5uVktXYAWSe4JArgdyACCCMfVckqlNPOQYQR8Dq6u
D2ZLLYEPSpMPN3Eak6cctHYyKg/uD4ly43abDfdsav3VrWU8ENLpZ7nXSMnW4XYiuJDazcJdO7/7
AugRToFuMts66Vde42uxvNgQ5UagHYq7OpgVXMFoaiSDLmrNTni/zNoiA1bUTXb1ySu+bLdG+Zgs
CC6CunB5Ltp7J14l4dYmxwNwXxa24tc7zfo6kaej16WTlAdAq1cU6cODhx3wzCsfLQAJSA5vwKkM
vvF8J/ebAJy4nFQ6eR3ioKVttSNlJCoKXjBcfvsdVV1kC1PsTDK2DALtZGtSHNQW/JAgDeSZ3hA5
Wte4KMr69sWUJxd3PrGuq+7NBwypYXY1Ya4Zgp1/aoe19pQ+QboAMGAtCZDt2JNtRHdgH1CErVx0
3sI/TFELIyFLIcBeKZ5GF2k2iEc96bWvRRnooZxnZmlGsR/VP3wVZfq1qwMMApwfo9q1xmYrHrDd
qlS7cXm2ku9ZrgJvNUe6QP1XZMC9s5/4RJEdRaFfXr/1fmFGlGUs1mAr7WlEHZdZjZnkJYT7KHO/
GeK1xLO7JJ5mHOnkkMVFmr0uHoxLxm9jCPKRGQZxrQBWhlWpgVkIsWhg8sLNU1XhiZzkR1dBDVcV
vAQzBgN0tB2PTBILsqAmuU1nN3RSCAiZTa9Mvb8CUABSmg2N62RyL7LrKYqrM579CFr+hIbwuVyX
QqjQhN9WHHWt6zMoPqDwlCNLfvkyjo1iMyaG9UhRTsmhz1fbNhyNn6YFPVvRLS/VTiKQGeVkfyl/
akN2g1gOjm1oTPTg3Ds6Ln3TpefD7pN50Kp2eh0T/9tuQFo2a+SfnSCsStRRkl8mjtq8waQ3c/0l
MfwNGHL9PS7wX9vMW6Cic/IAYtaSG+sBPzV4EGcjEgQTDknQxaAPXsMesoxbptBDTgDJdZQisMLN
hz2sTDGpxTC2UpIluxC5XxvoixZkMLEewjlKI+lIUbULKAEOrvBKqSPn/OcLYYrXpLu776z/yDx5
Ss4k7wWiXB6+dqJWwDbTtqi3rofvUgjYcBbAW98hJCe01RGrlqDN6eZiYPR4vICLrSmqc+QBhW/S
mtfVuoDgJnqaohsznARZPiuEGdXHUaaXIfgpwmuoZFsHkULdQs1uZcxnfVCEUcl7Ql/LB+H0OL6o
evnXnF1ZCusNcW11bKo0EP0aztZZZLpVVS4gMvNu/X5UbFQ51+4RCrZG7GMlY7aO/tOsIwPIi2gQ
2GM7Id02dVW6HJVxoWG4x5z/wrhH+B+u0DIfDTl+O2cfseCGlfAqUSbkhntbT+IEBZqk6JMrFeQN
oyaqiOCuRfI+Xtf00y7Y1Xafm8rnqGhADdKGbJNTEzycyZrCJ1VWdzmgrkGciG6qpQXRhXSeMQAU
waRlGCHVyxfzvfisBC/GJ4MLvnN5LuhQoVbsQCkKt1FYtJ+Ux9nfkuWw9+hLM3JdmnV4biMV9M92
Qv3E2qDzWF9S9LMo5/YBUzMssDLNxSsluWmOTLxR03h68KxQFoTOr/ramKcOOOq7bTO7fJwYyGT5
nyh2au7Bosti5Vrmm+98OJ7FhQCrNHRzsCyo5u2CWoeWv3EPDeKg6fDO5RXY7mHXkZnj7tC2siBH
Irs7qn9bNKoia0QFakz4TdzWhTWusjcxSYrKMJtIqMWBFcPB/EbPhgoqR5PJn0eUqC0PRN7AvPmT
lOw056AQqu8Sk47xH0FxYkZNoAdyZLQa2GSC3AieBkU37PYqtKdGUY3pwu1ghdAZ1La2zHIuCRxK
SAdCQsPh3OEHWC5iijJmLeuuzI6HR2KerYvvm6921TSfP1oY+7BcOf2NhbupxGEyueknwlOX+rDA
aQfrb/DPSDJOp45S6Epg9Ah/e0Ux6fIRxoaZRC1FuCp3FLM5nk2JOpJX2FrOmAZoyiUxndeLR4i9
gltfke0EYI1xoxkE0mv5knQWtPpIC7PWxHI6ljD0XXtoFGyqBwL3wP7bA5/tQsyi0pcUmggjfQUv
CGS5kiXWdgFQEL4cOk+CyKeKCOCR5rT9YRa+S2Ot70yUCK7CsxqyQ3QLSfL07mKYdwZmFkoiYNuH
FAMUMNysdnl/UdfOoiFR+91cp3fzW0wm8PYtqPFwXy5sFyReDCeqNlupbQMkdp93lIyNwXh42+uW
KLt/W+FllzDRLpvLeDruKcV+TItBhRs35tW2NYH8S0ZZAgxddCYqJHLdpGeC17HL0Tou0mdORc2A
DJnAoKyDyjPoRpNsjzzMx6wZ2KwrxHMd6o7IAtBPC49cvG9xuLZSvu8/g1PbDPIEMtinvAekKO0s
RZIGZ7xjG+2crm8HHiuwisTHj7+joJ2YcNUMMLGFS9QOP/qvj3SzE0QF/ZnAETcUu6id1TkQteCH
qd2ahV2Ccv9sVTXPOs4DwPGbM8VRStBbX8BDeTv2V7AoZq3cHQRpuoV0t4igh0QzhI+ryftopGJj
NxEq5v7hRjqHJ5phHdN5ZzN4ifi3DiLamTkYgwScnqaTmm/Rhyi2HsxihxowEyGJa3bqBNPX+5Vz
DTmYRC0ISo+l+jzg5jSFVE2FdrxFICVn+JVFw84NVxPaXJ8K0P4yfuGuEnVNYE+c6LBM/T7TxEgq
dFZW7MuCiwrOkknjHOZMZ7CAjiMuG2WNNlggeX5ASelw5VeBvnwtijAC8yV6VsDebdMRPjoBNZgT
y7J1ra53aNaoshgnwEFdbhmBpNVvBfc+27qGgdbE3CxG5BygLzHyrkQ0abfBjQDy+m9tVOt4ZYa5
3kBBLa4atxXBRTe/6rrX1wtO5pzAyV7D4RsNjSVq4+oDTCyMjPZOXfWMx5UQgn+ucprDxeX5gWA3
ni+me/5EyxxfiWTSTAd7r3+Xen0kjBm3aRQF7NamAmAKydzuTvaw+Dc95mKe3a/9/Q4KEpGV09N0
4q+BB2NvZYhTry5E52qIiYzmVrs6OOzOv5syQ3wVvcX7H4HDYEXxuIDdpiEtiTilKUiIE8JlA3Qk
bGBjjHi62xwqd5NFuuXJGc09pA9D9S5OJAqMSF3S55ROqFgK4Bel7TbLrrxIuzG+dJehHHmIbfqI
KtY3lfnbzlTlqeg9yPjdUA8x0laUGEUVBXjhoWpRbYBYXn93ss4ZEITI5KFtNI+kQWKtOEezIWqu
J322980Sw9NdUoX7Cno3FzgdRtJ8ZK2vOzzo+14v/2juuVbT5cn4V5DRz0sbIN8GPF1JJRaxaWo2
Xz7k8Tkp2BYJfGGt1pP4lV3vwS3bBR/qOSPDGVKFUODoYfO6gpEedH19Pxda1eUrACNM58jn6k+s
el6nepZP0fWtnYlmC/MUqF7Yj0TAcJT/NiHc7HTW7L9cAOxU5H3ggx6bvdQ6bU502F6pHkvOL38h
Ur/b3s/M4ARb+r+RaIfw4ak3rYK424anxwt8TbdwVrSjJzmHO7+I46g7h2/MuilfCwlQop189jaD
9V0vn9lM0HDxRCeSv+CYem0CFQ81wU1N6VZycBCcpNQmko+Md7F035mCr24rGFYsHhgoDN+/6/zB
EnLWrFlOT0KLVXT5Eb7snnF3xMexhROs4/rVgPI8jLfOnswtyHCau/BmB+alXdO1/68tLJAFHcqZ
PTVqghFzMx+///BlsgPeYnvgu8kb4TVimdzM9eAk9THySveONk/OnL/T3lALFGty6yHsxXi3iZY/
kSRGP1OvwGf3r7vSBMnmBV0TN8lXVmBl25SYJo36hK1rAppaWIzHYHlDk9Z284QaqtC81ETC1T+X
1R40AueafSFndfbHOSGikBo+2thrFsimZaeTIp9yIRx9Af8rDIFX375+QMGlQZzYSvYgBlkKM634
WdahjipLCxeEPB+L30vMwF7uBzyXDHs3SDnzDRRnM3kZbDERNZAq2JIKVwKmAaJYzURGBpO9OfM4
s8heDqyDHEV+Zh30MAzcu/cTPy0Fp1rj14WUU0jFWSg7C1wiunU4cuMbwW/ScWh+sfkPZGpZTnzY
rtJfCQR3/NqZYz5kaunpBaZ4QVGzsIdN7D6JAGIDRZfPf063N9QECAYdnXwXoVYzhJF4UVKIL+XH
pTd1TxfeVL6NxKPIkLDjWUtQGevpZGWjd2ddw5NuDuftEYV49Dl+qOgn1TQNeDmv1Sk+yEfzQCi3
MnRZDGo/0n5qSGKEElVweYaVSivTeQirZe9ZQQjbJ5yS++DWcraF0W7U7Ue7vbx3KM8cLgwlQeNw
hswtAURnL7FtW/4rbeaabrlvywCo6T+Ry3trTu7i3m4X/eCl9JBijPo+iUTKn16umwz+8bi+zkXB
2GD7Q4M9mJM9oTJW/7HTzsCdc/kq9NFr33tXEzmvOETywvQCMYE+6kLriq5+6KEZ5nlk1WPnVKe7
9Xwcy9nbVbiOvWCwFBQ+nUT9+VX0hgr7IbaX7F0en50ifC+NzcLtBKg+aiHCw2/Q9zSVrcyLjmI8
t1WUyXld0fFKcIs8s9IDfP5R+qPvbI0/a5rloYqJ/68IkoASd32OE+uPQmV4btKlD85zi/CpurL9
hTqK6mEMAJKjWezId213sAAVdbs6rm5ieNsTDBknp8Z7CRDpK3lhHgefime+tdrI3Nf8kgC+Btij
fbtCiZk+fpHyPHoI4xxclfktdbUzNAYPmxVX78Dd+/I1EsVs5bpIisgE4q+sSUaf7wJzEnB/i73o
18x9pORrIGAtFOwUmm/OB6FW675alPjxFdXFEER5cw1CtU062J4TakVfwxicwR3GAkKfK6Kfiw7d
tMfOXRIlLkU1UQpIkU0hlBcxj3MqQV8FIhxpWwtq2gWYvtRaZM+gUt7dK0Y7rQb88OmnhUiTUJn1
DsDkKcRBrSXrAChXoF0/hTBIm3Z8tdgEpKo6m5bWyQAmoNYfCIWtX4AJJId+n/WOehHnicOozahz
BnFOuA4gze9zbQ29lIlIbMD9kovLzTDXpgzUVD7CdU6BY6MGGOZrZVXkUuHkGkOl972IATrX3FGr
5upFHAn2nPrkq7DVvz4IHADAq+0XVyrSG38OnnRVHu7s2lBNfL/Y95up5ag6KuzBzZEKmQWSgJpi
TEz/XIfj1artNEMc6QTNqsQb0hMEydRC7Xx3q/aYBN98S+lZFN/CejbHcowV3aJSZKynzeBqyZP/
wnTsuZguUWsIRGF9JU+oN3y+ESEmK7E9UWx8T0J7cPbExaAoz2TEmuCKpmRmcHmIHNVrh73oL/K6
qkdk1W9Xy8HcFOe3ngstxVVJm8z134dpFhW1ECRbDHzTW1vWaGLDEx0x/I24FVB2VW3pOlyAi83O
iwCBth/iCJT1o0mINjr4Zmb00cW9HjkLJl3ekL/GBWBGmrEuTvuK1vG8P5K6ywkqHZiOHUmhpcj1
tSSeLVNN0XgKLd8Nxm1trkH5+KFWZ+T2LlwbNl06DZFFo/MaG4+DxqnnzsKnvBFlgvJplc+lAZa5
LEiHJrqMBSwY2iE72W4Oj8iZ/T98NBi8dlDizHTrEr1eP5fmTYuiHOqYeEy1IiVW3Xz+25a1Zafa
I0uAADAum5LdSjQN2LdvCCIWOE0MFM7xQYsX1DCGYaiKBj2XDXfLK7JnWEeOjJSfZnF7XdTKrtsl
memHwYrp8p5+OozGLDtj6m+5VUrc2LRbl+aqRL9uCWp9p9kej2YnyJ0pDatTjy8qbFoC6Zwpj2UP
sLRxYbA6c5g4OPXtAYFTUeQq497oOhj3drzE128Bbhfa7o5V3bfrJBWMH1HZ38/jBVQI9CEZ/e8N
BN4BQAWA5OLC6mT/dK9qu2JvEiFvVPfTNwO9BgT2bzMbvbmbi4yr8X0iD8IQKP7OvK8ub2IZB/Ue
PlvkNh2a3g+tVm1O3BUh6DnAezo27zSs61XoofqSedzWMD1qzBWmgyeDluZZcA1NXv2N2QYBvOwG
YWTGVfyWtel8R55tlPsfwaOxTh1+7F6L3JBw7hYE/Ggg81wdgk00cDIxugOViZinsviyPj5qfb3B
wET0xKwGfsfAMZ2pBSAc9NG83+FYgE4a/D3oQGYiNiqIPlMclFQdHDVaatUVczbUVg/v8X4EH/ne
HeTVCrHGCM8NNDR3zyYC+4gH2jvrtgsPiNkdspZn8NIjesoYASsBp+ftinhErxtnFM+0UGFx6hnn
p01kptakMWKxcpffy17sy7cG+1Ipyl4FaFuJrk5oHQ5nptHX196KnSlyDwNWFh/5wSZtLZ5kYxv1
M0lJ+/yvJeonbMTOVoYJyFvgR5SBakBQWTBZTlliarmF+w0Hvow39xV6rdPKJEW4RQgp7bH/l117
VCGkbVOBL5hgYK9XH1IMzeu3MxpahjgNuYpUEe9Tq8lbIDNiIK0qdJ+lGN6FYxFxFO2Vpikk9+bv
eciRDepSu/orgU1k1AUvgHaerEBNi40bzt2SMGdPB66c1Gy/S9jqIa5XFDdUtgDVPwnYPkQN6kod
QXZcN0oIpA3j7NORtNTgrO/GviqIY2hqcGokmyOcm4kEIhY8MMKPdU0we39Bf6RvBMTFbo4ah9U3
uPtOJu5j1B7FhgEVnwsDPdgGKp1Vtl5q8w3Xj1qieIPjrypPHp+ydvVegfBc1UFDAblNReYIPY2N
xaRxHQISik4/5QMX/DEHC81ygfHcZY1Rsx5C2ZmM1Rfpi6yFs20IToVTWsCJiOmcKlZE62ZLMWXi
ES063uUXLxUsujEByVNDBH5P9V8oPZ8oS7fPlEvUzQ0dABh35UnXP4XwfyXq75wRIt6AiBCjv+Z8
a6iP7o+Ap8yjArbjLgxRlB5dE3eac61cs8arOvyz3vErxw/hSD3tKJ+QqmuVY3j9ab9okVZQ5i9a
vRAYXXlDiujP/nYdeRQXB0q5MdSTSRrgrwkwDwwWnNdXbJo6gbJs5ne045Ztf+FW+9YBw4/nijBu
emulaTSsubEjiAb+1iT3XX7LbEthk+kLj0pcJYAswvGW0P5vIJ1eKXbUyFgrEqtlhfmUXj+fvU8K
Rl4xWIuGtx6ssQh3vAH4pEsEGhkB19TOGEnBQkpITNMjvxQkZBkEZDyoH9LZ227Ry3yHm8HOBupP
SspGartzGm+PPPD2Kt7sI2/BhMM+ZllWf/82Y/HjyyVBlKkI3EmH89NuT+fE3F1CY1x4FC3eegBW
C6JWlhB1F1K1wjJ6zh38KMUjMWapr7dVVBj+lhg5QibUf8VwYUqS7YGupfSDnbZJgPL91ngSUQHb
xE4z/qRb+o6mkOKsFwXfeBeUIOhHKkjjJl5Yfln4pB8+8SBXGK73MOIOpRbTlVXLt7MwdlKXE/D7
G7z7cybr6PvggEgQa7F/5T1rGwS/unXBh/4yv0EatE7Wf4x3Bse4N3NBQPOVml8c9OGBCzoraHvr
GZyTtOc7N709IVqHWr4qpIyDgciPIvR4hRWXeRL4Z/oj/upI7GJ1+5IX3Xs2+uI6KQ3MWUt2/jxf
rmid/0f6lA/42UhYeblj5MJSeeL/MvpODaoTEs1Ir/GvSZ3JxF8nevtVG5ZvBd6haLhssYy4g2qX
gowBgdNJ0CdGqO/ucXG7K9jTVLfeQgwRH5gRTsl6YlQ6vbqbeiJNfzkB2HxpD0/HmBebNXCZYkth
jasSu80PR0xGddyC2fqUxTEgHL6TymB3O/qWYIOFQ9q7n7Md2hJqgEiw6EPsXVqDL8NHIZ+S6rD0
SBBCuwshlnQAAyyr0NrGUbQgKqjKcM4WfAVvo6J/Jag4QSeRGAKaXnOlymdzqmwiLo+UHjOp0mzU
p09DGbN73iElFGl9wQ1Rf4yPTcMdMTK3Eh7G+lF3g8wxYRsTlWzqs7EarhwpyoYC7Mff4wEZBsTJ
4tsFrkgXv4f2+/tJshdK4mD1q0RDRLaVEg/fN4veecQvTd10FOSg1r+5FmDIZA6r+q/5ZCRE10e9
mypAxgwDj2zLMIOAKRBtNP/JYKzLNUTF5PucPEAoUITdpBQsr2g0plGVClotPWTECsPFzxltH9yr
lfI89+8YVxTEPGJPneLi46fTtgZ2M2BWqYlkU6AHTs1jj5oq2mKdHFoOgPr+T0mi/y0pAADq/1hJ
t5uoLnY/Zxd5sy6GACU4o++qckbYLPK2NmphhYwt8I9nLdhbF7KANUsf4HVBuiZ+RLT7j5qCxOAh
A6hV5LuC+BDjuyZ06yGbg9GvMTMINk07h9gjDB6NqYHiFIc5T0N/oydB3ZR3yr4r3gqZNdEKc3U1
NZKrvjTZcwLXiWX9KAERsoV2LPUtCR1bAxtHOeKVtyKSQPi7cgegeS2Y+LIDVTDmhL8gXZZdbhnL
U8pv0DNVAJd+g5OOqgNuWE7VMZvwdaMIFI2MCQAW7E6gJa3FfhZkL6RbK2cVSnAE5C7YGpI1Ge/8
hBJsV4moPzCgESez0s7yWsGYJsdByDb1M3eeZ5WxsMnYigN3GnNrz9LPZOzir4pCiwRZaL3cwhmt
YsFoLzLwzpzXho8XifpTaGvlj02fs6QoqHyawbu0KQp4HMCrcG36wqyaMZvAsRmCijb/iPTU+lzj
FFE6vN8mUF/genQxl57FFz/JuJqBmGCDuu9laVfuASWrze4m3AIPuY5woZ0otQdkRHCIYcacfV06
pSdEYWA1g0nBCZfPh4+47pBMhJEO90oBZnCkoGRacnSbgGHWvPvqkCtAJRb97Jk4iNudxRENoQmn
zQuSUMyiSXDxtxrZr+RXnnZaJpAXbqK2UW0evhLYjs4ki0ONW7MQUw8SDYlwiMJTcRm43dm1WJmy
G/JZinoPfZnBrIpzgdshXJCf/Tdv0R9ILwhxVGpkSskoxeBejmwFdl8b/O5s9eU7mDslXdFRhnWx
DrQNQNziMxF5udlSyHrzbM/NIFZCT+HkB3c4751f3A0MifU305lNAlhmj6jeXisSRIGX4rv+b6te
bVn/qfSRoH2iMvOhJcN6SAehpkFs/iVEDXOA6AeVnH0u4mERe/od77wUMUjV18HGelwqJQ6JC6oL
qSML38XsnWxER1pEEP5u1qYl9axSUBfw9U0sQoCHfOTiyrn318z0TohVVZUXWl95mwh0guCkr0pW
WkjXf/4kvG49c8MkJf/B1/q0dW0gIyUu/8UZcZ7IJkfcOmOpLlLE3Df510Co5E/g81iqzWGiKEZ4
mIrPn0jXsu9RxJS2ruwipVFi83HCQMyM1PyO6s3YXY6rvMhFaJu2u4ZofeXSbKoY5ztRnEhvSp1M
hdZLYwvxJi2XyOUOJQ3XDJIvqEQJRESb9pFiTzo7N5DluxFkT3t0HsPedqI4wdwWBBNUWBS08wlA
ayJ22sfQ3va59o2d44hDaxotZHgO1MEGXWTH5cMAdfvHRZenHFvj4QevkrEXOR/5vq36dGpSakVf
WYfqOoXINX8rfziUQYmbV6cdKszR6sdN7QydXp9vL6qbb1kfOfZOx+0J+0W0dqtn5m3UQerJNgp4
fHaGFjjkmTC+0KrSc396806BsS9MG5vkdcFZLTsvFToWhSlIYB84j2zqpxSgsPPjl6/QHqPt4aRK
kTrJxfAzm+RrgjSum+ru2lF8dGgJFOTJP4sqJ8AWhxlRMgFdOQoYuYS8SKh5Pm5JhqFbauuqaO+k
l/tyis++QHloGbPbrN4Xac5/1dY71q3gpEfaOSB5NMisGpKwSdRmo5DEzyrUR7ZctRCQ5cwO8Uzh
RUUSLLV4BbNylsxBllq047hjFJ7b5hs4hV+Dnn9GeGj1QrgpZ5Nh+P4XpHvuIP3PBzdKmzihxbkK
1Ygjz0HWycnsN9XGqD4x/7QE9UuFmg+DS+iB+RWa3sSQ/n98c++TCuKzymhaL9+RC89EfC+qpqWB
9rhat9p3py9e67iX1TYvcn7J+rnl8qBx7GyDxciI7amQi0NkPd3RlYxrR+0CUlFMJmPaSUU4LMYy
IinkCIwAQkWx9I0AGrfZOFFhsxGQyXhPv4WH1O/FoQeUDYyXns3iouzNONTrgOhM+l8oD2dnM1CE
Ybd1L2tTB/606DDHtAOvvtcXTJXgsds8uaGL5xohEwsrAlGFk0B2pvQZIka0BJih/VzZBVsS0Uu1
19cP5Ih3657ntYY6oa5Rp3ypxtVO+S1FPIlZkDi0C8901Jz7mkuez2a3wXb0jxj9kul7REhSEBqY
PjAc2DOUo9Fg16uFte9L9vFEvTR23qxdIfG81sTmp55AZLcvTAxcCh0Qv24zSQLA6XMhh+Ukdhe8
kqTNkB5adS+FxmqqmW/0EqPombrnMM8x/hIE9mzNadlAuSvRlOIp7J2ao6cxOcg7FHU9dx42Gjwk
V0ibJky5VOSK6KjIl3choET3j6Rge2/wqHdgskZng+sgpo4ivs8zlycG6EhV6hCtpEyTISIvTP32
5Gw8kn2Zs9Nj7f6Z2HTmBofHvYMghKMl5HQsB0+T5iW2VBIACK7Ft5J2/RzzWGiBLGaIc6E/+NSN
mQERF+IwJ7l118FfjUqXr65JnoQDAUCQ85XrPhTC8ygdg1/2+h+szZg54NXlC0Ujsh2IfXN0F7D9
yA8nqyldcm/UdvGKDsSaPSUCuHPlo0YC2RvKCGq+sJIty/u3AnlX0av3C0+pUOJnjbpt155M8BpD
9LZQlKk8QQb89Y1VuvmXcqMQm82bkodRE5xJQ1gfpgnUkdIK4VX19BiTm+wr5sAFI287XnccBmId
eAkXxnumLeT0/gB97BVF+fa71oR6BhfelKKaDKbeYIhgqGAIsuytfLzRXEoP/L2M5b9eO8y0VwTy
lXijAdIYnPZ7CJh4Wo7ypfVMxRSde0NTAkAzRyK/kAamRzBQgrTEB4Uuf6xwbhY3JOoUuMpLm01i
zP7yKlzf+8jdCaJ7YV7Lb6Xjxb5n9IRpYQgkOL9AIhCR9MLVF4Mk7kS2POyeqBbAnGPKJUbMaUzV
JhWxs7cHJ6jthSNG/S46aNeaeOKW84Ym+pjrb2R6g02sZmQuvp+teuA74ecCLAip2LBGLL/lzfFP
sEk+P6a7Zby0HcfiQ3QcBv2YllNCJzjJ05Wt4lTXFDNelLG1H+r962rbctvCa5WjhGffmZTRvoCy
Phuc6ddy8DU4H1ExI0odaDIUuaQe8eJEg2/FMsLoESli4bNojpWFguFVAT527H17RpvfrqGDt/y+
W7QoM/+NMixS44qddzOZc/JzqqLO6+FKNI2OvHH9scIJHLaH/630Si+DxsgWFtlwbJoyy1wG4Yzb
HGQq0vG3SzMef2DXkRHQ0GCHZc2yrUWOEfo7ebNGcr7LRloPjMFGUANV1kaYJfFENjTPoRsjsIRn
MHgMeHlT9+EZ5fU7X3H/tsH6+BgGWsPQZ+QJLHhSI6BTXNIM6wmcR8eTFV6YDgHVD2gM4AkJHcCY
Wl8TRwHa2WsK4dhHN2nFGyTakObpafiqWAJSxZ+LKqUO+cjGgcElzaWc02pgDmnuWxxxhHaFGSqd
L8HTHvDit8rSvMMHrEPbQvGbOwJKc0rt3179/iJzriCL/og8Jeu4fIP+m1hymwCr/C8Gw8CFJwdR
RrnYlEPJ8zp2QvhxyW/HQbUnn2P6S46gd0EZl/WjcRrwRB2I3O2hFmcZMbrGJII4Pve2p/ggnyxC
rMCJp0xfqddGUyILqOl0g+a0BMTUXG61L3bbUxiPAG0iZBEjFeOCbYWS1wm+dKR3Z1Hakt9AG1yQ
5qfA7Lsx3MlYZEWrNnHWq8r/Sx8MOiJgK6ZcbtaU6yZJxXXLANoDFHZgWEAhYvTMuXNITMhTxiZZ
oE4fWoCdx3MOtWE+Kd2+qj+i65CWfjZBnTkzhcwQFnvs4sfhVJrSD+mJS5HSedm6+LSeVXzXkAzJ
e/FIylnGP4wlYgofE3EK5lbZcHzVA2ZrFTY5SN7pw0b9CRv38YzVPWy1OjcgHmH7/XS05ql+zaic
cbz/1Chhie8pVZhf6agIAlm37c9wwEKFROMF0uESrJO66aPE4erchDGyK+KvRUJqJFSjZkeD5Zb9
+Bl/w/kPcpPySpc1VzRqefcVjsncG+z3BtE5WU09A7jW4xoVaud3HVNjvJ+aeZFD1dxXyetgTOVy
w1nAX+9t2CU+XSilAUd6dQsS5m2c5mEtqxrmq1MRtwfty9ZRvOKILizaWkc/Bk9yTa9BRuf6NVQM
CdSUjxXGfTmJvsXb53HsSP21ttvfFZaEjLddHzWkr88Wor4ldf/ZUvpReXNSbG0p850Q6f1VUZM2
1RbkpnJV+HEj1lBoVcqrsREdMgBU83voWpnbuV6b1f6OcgF1h3m5onksDTbUNoy6BVMPqWOB6PU5
ndOzPD/gF5roR3Luy/xJFYxF6NusFNi4NGyBGFdfkfEz6RhvvCyB/LyzggYu7T/Oq5wK+R+IEESZ
4CrbWxOCPepZSkbItokeZTs0XUul1iU/VYRjNB2k1zC9QwcDASj+nE47HTUvw365lzhtMBPqSZHm
YYnyX3sUZVLMonQbWflmdsIDZJoJ5AtAMrK8bsC8a4Arx8V/UEIIZiNrwogkjppJ9y0Yr1ujLlSq
vnnYCR0JYI2rc85yI3pK8eoylHRRiQgQkkrW1OGJ5hKbWaOGY3IaAkqUxZTpAo24roKDwBgvBaXx
TZ81HzlZa/x4L2BBSZgA5hCd30LrAZ0gNUDllD3C11hLPLkilGNjCrm8cL6iin3X5VRHXPrPcPtV
VhgPw5jQFoVhOmo2/gwyQvZ2uOqsu/JR3jS30xFA7Sh5Fa4rYNzmZkgZ597UHMjZDitFfA+k+LjK
R/rIHdpitBI1Dqi75KVIWye8Obdy5jVTpFa6nmH0LD1Kg6rzYj1S4yMWj79ayMqjEbw1O3NbP+dh
2KC+XECUClPUZoslHWeFyovpl7PD+IjDq+zDthF0GsMiO/L9DiZ7BR1/HhHILNF7ptRwqmNxf51D
HfwCfGrMfQMK5IDIJ5rA2NuLXSStm2aseDlUZLw9lgyZ05JR/jlgTrDUEgj9jznN14uPwg3aDpRT
YsHjaHoFABOko3hzO43+JrH4vo7eTXCv/14cKzxEdjYBhZBCud5sFhHsC41uggEONUxFdkZiVcPf
g1TLlI9ZJ+XwOqqsHoyaIEdmcGzy0YW/d0fn686Ig+fInpMRFyvlZt+786DYy1hekWXjl98yOxbS
MbniGtC+iYtotKS8WYIIjpWcklerDCJXc8XZo/0pw3cpPgo232vbVQmD4Xk7ReQBFz5mNj8ZHlb6
xta9/eRQAwmoZI4wqH4Gx3PQXBgq0lGSCu4F7EWP26t4ih4V5Xs4A4Ray0W4HaoFLlzRCob/o5Ev
5wj8h59BAykhzsseaNjpO7Dfe7f0yLDg2CdlmwLI8BV0TjQkWovn5Y8rclwtjPy3dbH8S0bEJuWv
Tpo/jfM3Wy8iO4Z7Ks1H6l7XaUvw1gtiU+w8uWRVVvujRPo9FRhBw8ORPoBBFLDZJOK2649Jvozx
x4VYpD/gJecu2qhqOYE79UyPzzPi+uRFVzWLSi5n/MSeb2eBDHEtO5MnV/2yFcEhn+RFrB5stKmh
ifXYl9TX/hWQbgYmFtnvHrHSlQHs4ojK5l03MwjfU3iTBxafdHnuvHyewRn8NFheKTJCb0/hIBiC
vZynLPDXmNOGqo5Ctk0rxE/nvMSvIobdwZ5Sg2ZT7ZVTNm37EOpWn01O6dpAPEDJpWeHmbXBYn8x
yVHHvCvrID+sTFIn8A/+8ej4rTK6mdJRC/c9WCPunhzEFVxzBdnSpCrecqCe00N3Nr1685STTr9F
uOJlVfi5Sg9gjOP8JqKmZ2YLJH2GCROpwrMBhmhRTu8zZZReP7KhWgrDyADJfbM9LmCLEHWTemaZ
DOMr8v/zE6W8K5shLOqJ1Q6e2LbyB6QlJDSzi8879naLqF//iMTIxEYK6SDKDivAWPoRZAg9WOrU
cK6rw3Rsi24QsZTsPuWaBjvKV5yIo7cHtYc1fDb+XQ4KmFcOsiTFP00K/BbQcqB/Hq9DOM59OAS0
BJb9XJLA/e+/o7qlBiprKZEqkOtUmQC/S+EYOolnwj6qsPFHDFnCzyIEcCIpcSAlaS85yxXqG8aH
cW20CLG3UNoMi5/ixxgGGm3rGDlkIJGO1gEeT0JKlXQsKDUMEDwsipYjSNPkRwGHZF5US3Mk5nHe
tLPOuRTEFDGwmEnZRCVqjFZeSVp8HJgY2G5r+iUMXk+X8FlVUmp8ycTVSCJhqYqR6FQ6Xlj5HbGn
dJyMYnozVGuDudXzewHI19+zTnVhfdoiYQMjG4OeJ9LJlA62fKOpbU56amL8g68O/qq1j5/P7ze9
aQ0wUK9tlBeQRtkHi80O+N9bZMaFYJt7LsMxJJss6XkjuCbOLWipz/rbPY31a6+ztTrSVMRpBRnh
xnxaLzu7ze03xbx1+BMb/59WI/fhen9ba+EbS+qC12lODlESak4F2km3fz9ArKLVOT6xRzj5iiWn
IEBbTKYqo9GoA3pH90SZfQZNIA06WXc5Z+fV3alCdAyR+0isQgejTTxeKQUKNstIiRiIjYHMDqxP
NWXJyfWQ+V0TMZOwVsAWzfamolmzhdst8kqUaCG315aAYd5Exc/WNUbYRynyolfttEXWug07fQKB
JB0NxATZMsblpId4D4TwGcmy28UR80HKlBfyG+ScpsOBIOC0kNkHgXwc8BQlyh6E+r6PyJt0X4Pe
yb+8tvaLxWkXCg7z0ooiGMEfb3J1xT5YTI+wZyQRsR/C4/S9YFes5ebav4XWpPntiKEbdGfbQth4
m0tG7ZCKFw7+7CQskddikqEjhDhpWJjQEQMalD11uCf5Cf/zJI4c4FrdUHU+jsVLXd6noqRy7cS3
S4mxKe2abPTwUhvdijSgTnc6H7+HYxj1KF99DsM0hw2HhP5BYgbWo3imFB59L1Wkvw2bGov+TAWc
B6cnScPJPhTWzwVtFiHsQgAVyKGXCy4v00HjxAJz4xTvN+CjYwSg7FLC2NBy+43xXjv68/y5iZCd
Yx243fkhjErItjLBR0LCp7K/uPA4k0Ct2hT/Vv9rkXu0QuNEK0gjhvMGT/hYQhjJSi6GMnn0Ct9/
JwxIzP/kagfW/m/yaMk15Vx3XUQX091vuyNqEQCrT6Xux5+JcbCuOe1FVMIT9ScFtbWf6JsF4t4v
wC4hYzYQA3/q4uQHM738H5d3zMkc5z5Fy3gXzt8ne7V980zxraAVLzspYML5kHroK4RPg9aEjoEn
8C4umLdSj9b2rksWA8UUkuXCJml2F5souSdJVPSQXt7jarcjKkBHOHWYVSG72+hjrsjl/CkFDBZ6
JC3/Y9PEeBUqeIJfe2AXsoCg1rreaukMnbz+KEtj1dSKcQlFZpYim+iKP39Ot1DkeB/5UxKI8FOE
MDin5SGe+38mxWbIep9mHl2KZZ+I2/RESZAjEWuTZgFaZxH5gXk8OgtLMDXqpGJPCuFvnAe0n96l
5bCf4V0ilFZLSe10LgvexE47cE4ycBg8p03NTy27gFjy0dPZwmE8Uct6UfQY2FkqnbjZaXC/Q4pa
Jak5dYnvml4h8Mr0mLePHxmd2KMrSuqAj/fFJQiAmV+4d4vJaGQn4+eCWu6IedBG/KphXYXvt/xa
FsekuzLyzpyf5JNMUIR5hjSaH934bdbRYLg3C0iA8Y7iTtXFL/voL6a6fbKtPZ95/qy0QvzYN3uZ
YPc1uTeyb66+kRygeqiW/XoHsYGK2jCZ81E7OUhIdOWBF09jf2iMRoE86YuyT7Gmie5ETZuveFQ3
kIQq85y/WZHwo7OpcqApVUJFPSlriNtHus1yKq6KugHAbD68rSOCUcdHS0RDabWx8EO5tdtXTW/8
Gzn4j/1qYoAWpG2EFa28AtQJ5JBD1bbJyxMa0OCPDXe96t/Ic2tdE8mOjnFtnmPYtDVZ+X+P/RhQ
OanvFkfhj9DDh8yemjmyKXYCp3c/m1LQL/Tkxqnk2ZuzyaRig+6gXYHz7Z636tbJpAwb9tuNMMfr
JWqi86TvIq14wdH/88q0r+8que3vlXxlFsQGguzuBGP4Z5zgsrnp8lRnN/HeSi6+P29xxshphNKb
OquPFh+ilgUMXhd4JhS4/LmVq+UQYQg+mYtOWViZL8B+XSaMz9UQiPKzMHUdEfrIQca6AA7gqkS+
9sE7ohVEwdS7MFecR8eCumi0ObZB8iUeykm7fxR44rpTimoTU13OpuK+Wp7GReRlWY2NB0zRWiF9
gvY43EEQKcm/mJES5sF6ojKouVZ4hwCJqarMeLhbP9Z5JPQ7sZWiDfoC5G6k1FIIeYSi2qam1Jk/
fWKpuFTitn/yoB7ERGYSLHRa9jLhIieQfPERroIWIO2tV+jm2GUCP4hvgZXuiU6Rugjz1dOG6S6P
uBY8Xml6qDEStHpK0199bG1d7b5bfoJwd0yRsETiQowSYYZF7mlnGDPTbsfSNKKsE/DF3DBJDafg
QH8NOFs2QFyVL0jnfoqC2uMjfNTrCRUtWYxNVa27WdHO+5NtrvY3yHi69wARaScyWPv7QpwL3yFW
HMYquxTuJfwol19dfCZVE+bZhKhjdZsDEagg/UjMvg3PVQbZ7QeW3aRy+AUo2vlbUdsX20TyZyzV
5eRvQuaPF4LEI1Wp011g3b+U17u9J5qHGxo318p+i/nFMPB0L2hwD7Zvl+uDiWbv7Bw6yAzOHvoc
+8EeiL2WRzMDjLJ0cZKozzevSDvnd8P6Pl9bO7UwseLENL9sZ5yhnjfPDetweTMVhtqwqHXiHqa/
pFjQ2JQID8L70buv2ee5JwBMC1iFethkzKJT8Hd4IKIymL8yNQ/0Jh4XxdA78nPfiqehpLkl2qdT
OjtESnY4DLh6VIXWsqKu1PFJbe6XbXYtp6q/wim6OsHVbiEzeJm0Og5VG8S7xP2b+YyME6+0fHOI
mza+Yg4OGjH+RKngzGjwgySoxQAmPwZ/BdOaZC7404ZTlg2C52ybD7RXR5r9I2BI7eq4Ry/IoacN
UvUTbMTSPhXIA7VtPoHbMyIvIJzTuEfQKm2F6MEZ5a+LyvZD54fw9AOr3KP+5maXpzJZdTMuSCVj
94SMRxWU4oCOndqJRaeTLfJySFQFJ6iI3j7tZBw/jUx3PWi7+i4jJqDYO520hXBdioFXNc0qaBiJ
fHMfMY2YmUO2wJy6xRYZc31Tt23Hf6CzhmRegE/w9KTCo/PE+tOXt1oe2URoeYsUhfHkmgCu+Q+5
r9utBJOM6pwwT+HUNgdeD834BhYXGNxFLwHIYNkAPOyKLS69rlcrW9EY2SS9hhsn9W/VekUCDwPw
RkEwUIVDmkB86pKU0VyVrIP+GWLRURg+s65i76Iy25osniPOAQ/eNU8JT3idHrjUOlDYlO5paF2W
jU4neJDgtstufdPL5Rs4REVSUB9enUvJ2xsi8NE4J/jWFJFDXdCNRuSmw1HfhEAKLlonvUMLYR9j
WaULsSnV9PuMX2chu5jOfj899J5Oojqt5hhLWQ+9j0tIhdguFq8cdLTCgFOEDRtYV49Z7SQEbs8f
2z5TTsiivqjD3sECv7lw21xRVufDKE6itkuolsiWkZ7u4BAL0HxBN/ns/AVfOQtplWnCG/Im3Zbf
qFQVgr2vz3HfG8siPfStgAJeS2+LFtmfbxdUhmBGtA6HOnaT/6p8jdk5e9EvzdV7Ht7VzvYOaEjm
ER3fyrsleS/ASq+0u8Kco25r0AZ2fY6gupoLFUowICPlCA/rgB/kFfl19byHBu+U98m7tAt3YaH1
kZDVy9EixOGE05n8MrNG4H/mE+BugE4aKTOSFgDQd81qQ3XbXBBlW4P+DaBQy4rOiv4yQE0Mrob7
zIke5mQidJRouj16074JX8SQuZ/nO5QTdx3KYRnhzOEHzG4yny4BNq/MMpRorFtK8RKr7EbrmYz1
C4TNKEJuhV9Cpv1TH0bPqlCpBNx8x27Upcr4SdYAicQtf37sRwYveZNefDEJL3zr+XZa/O20xxoG
Lky92K9icFaCWvZLU+t/GwFYF5C7wBwjP5fWwZ08YRXGzw0DfWhrLYN5RzRS//UZWqsJVKJGykde
U2DX58s+4aJEi60+MPYLPPHzEf8v5O5alE4bgqDNK6gZUKwptgcecOsL++kusx7ZhS3P1WyAeWl4
IMCjWaATjicgS5zHTmDrd8QEWjJAhq0SAOHJm8hTWsr4B+0e8jJywSQ4siOPJaQ/AmLUFhqph2b2
FidfVlwkwrD44A/lP4v0M7Fn1aCNgKw+0BRMk4tbOiIWMN6fkyOqnTXEu5vV8P9XLxMnT84pZLdl
o80Cpqnwp9gDuXvpN7oudu8vZahpyk0DHGrvUbE6yjqLIhGECZSugCXl93ZLkqCYBw/lnQK96UmO
hkqePxh8cU88wa4yUWbRr43w2JcSeVaq3kiN+5lAWo7TWwz/Z+FUu0shOsi9letENJ5Ny15VQX0N
/LSPVAQl2aAOJy6di9CyQNfkNR3Zl/nlYliJX2n8IgSsDI+lWj3RxSQwVwRgldp6mDXbhRhWWDM5
IHWzxEDv6WRaAydfE78ZKbNlpZiUs+zs27OcIZSbHen3aiLNw8VypTQT+TwrSkFtH90EWE5wnl9N
VRu2B4rRgrYTqUPmZ8sCIKoIdcAMbY/RJy39KTqlnecnXhVMGH0PKp+QUxwlAX9ccfJa5/L3TKU7
IOqpF3Auc32D5M6pofRic7ViW4we9zxMCgochsFLOGoDcLcyFHE+6YwkyO0AOfGvRQENT1CrGSOG
25O50CI9/w1TZkTFkjsJ535Q1pyj6m5wdTanHdwtmXKn4X38QjQUjU5Cn3PNvcZkJIi40mK6GGXL
GnD9V4+NcNQpvAyupcrUgOM5w5AhOu6eWque1SQESHVML1tkDs5iv+sI8xqAeofAO03vnpOckIBR
YF3A2Kpd+aIUpHROV+4KY6iBsHKrHo2BPix5MaWwP54JIFK1r7N9uCOh9LhvM1bVofs7R0miNBji
+p9xIPyfjWatkrf0Cclv2tqOwSM4s1WWVKrCPTLgUmkzBSU5trys6qi8ljsbMVqlY94/IJ7Cl5nz
TepHqKETVeHDmvxD+bXx7MjwSgl0++bk1WsVG3hdD4LazE/HqKT/KVfKj4rIW1JAFBGGQFjfdt3p
VDfpuwOkASXCpkD/pBTX/Xco6VooLYOt47GVNTn1AQ8xUymuPl/xp7oNbYkdId9Zvx4jfif0e/RW
nFvyAIJ4EQtKxlabBMQ1rAN20IyoZwV4zy3lfBySwxMUgleNpI213x0F654YSlWQaK4b49FJNUcd
gXst6+qB8uuHRFx1db+dtcG2GqqCRC9pdBLb40eDF3M+yX9YoBszu4LFxnMjwd9rzWdHysejBDyr
AhXmVF8y5VvNAS9oKhJVsvPEhRdO+uDls4p336LbL8Bqfo6keHXDH7/B7t0A1nGEsgbKF7V3oPOt
y+kDLsA6f9dwl1OMHByHdxnjYIiIDWArfSOt22dy/L358PfwjLGZqgqBztuNPYvlg/U4kEpWtJ8b
mrM9z+qsrLnqFVRsOR0faOjmmtxjrWoz6n/NIKgnVt18TaVQgNv99mX8LIesU6RMlc0xM7+2zIgB
R0IrJ60ipU3GW7jrr9cUCXGDUV+A/VoI7g5Z+OBPPww/L0CffiYr38UskJiqV2Gu0L9rKHkWqlks
NNEbCTCEEjfuC4FFEShS7GETaEE0Oh1VSmhS41HgOoXA+w87kxdAnbe+IveV8HKE9HREcTsEunIy
lPZdJrxl5oOHFXWUMEXikbYrvzDhjp+/xsoal47+ldXSFyBLv4YgEAc5hABsq9NFWFrshNJ6YTUy
5VqC3Zt/p4QIt/i1OIve9YwHQw/eGv8jj0AIsRXD06DV23HgweRa0pmJkyHWDXSu+zpQ0awtxmK2
ukeIFSDz9KRl147FY6pvz8ZtFU3i13tikl4Gmx4pD02XHAVZhqD6HRRccUQxdFhNUYTTqPQe7CXY
kni+qCf96nZpst8MPkQ7QAAXfhwVDm3qordYd0cGVfON2ne4TsgzGZp9+SYXC6dwn9RPgF7DvZg+
BgGYI30Q6GILQ93WU6H+QMFWFlKae+LWFOKVJJlXQXylmCe17/1qC/lvf0tfbZb/Dth9Yr7/bk8X
pSAS0+gtwnDo2LxXP+lxXH8LJuD98xxocy7vWyMyTPMCvkXQG7IapEM/Hhzt+T3HPqfwPo5KUCNC
KTntUeRGHo9RaOUvgXe2la7K7Ue9zVGdQn0JJmQxbhT0JK/GvbMrHgzuXGisp6alsol4kOmfUrX6
OYI190yOABKJi0F29qMAM5+Z1d+HxvMzq4JeULt2ZXhGtgDeYlQhIuuC+weOaD+NqV4zKnUCS3D3
/Aqm48mie8tWvgdy3WD2t9cyQxDhQ2pyQJriDoWEKg5rPx6gU1i+lMj54i5cROT+4z2deglyzrQd
sCVNecDgEQBkPtASgqTdoD2P8/hE1rJyYOKI71h/F1j2bDSmVf4y3Yjpa+Bx0zkK376ggzWKupcu
e0g1n/fJDi+B8pSmecwhwVCpaH3QSMYth36R5ebm3EW+/EUhW7BSvjOBGXKs6yFbECtqc6KlxXOx
Woe0hlN+wcQoZlF8ma0pGXOQSj9RMNEjk4B1yFgGMXQpUt2rzy5aGnfMBRwywChJRSlccvdYlTKu
CmfhL7vYs1q8GUTtG/kCbE6W7hlkAp75QpcLZAnX+ykF4ZuhB0izCs/BLtKz3QhjcDE5px6xh+cc
f+CBeTEtiVeaqaPYxO96PxOdtNjDuSyhXxXm4ejbZEFd1QvX+bWxdpekanXH/JWFh3VlyEQNNzPs
pv1cdcCXSmk40VvpEzQGfWV+XUoYMrATg65gS/uN+RGJ1opQ8bGYs5NTXv2BBDYXcMxyIz4mKNHk
Jl0zn97zDVWscaOnJAFNax/GTapNz5p48u9IqxkVGs2n2wouGq+edDr7UK6+COzcDAUpX6YGQ6Vc
IZU+ElqC41zVG+DkSfhKQb/lWd0sxYzvat5oxUNnlEM8mB7/AOhbL83yjo/pCcK5oHPiUQyirZBu
pdDzrwsLB4Hszah/ofJkkyd075Qvjt7mEfr2jDybp0qhOHeGrweYc0jSbkEjQ76h2U4iERWkOCq/
x5z+16MoqmajEoqHX4hQcP1w74xm1ExRmJbQP9rytbQ99O87WpsJUiXcjGkOj47ipd/fx6pw1s6L
Q0cPLOV3T8w75rhiCFtnfzXk31JRu2FCs5Dp+JCe3eCar4t5gML/ENn1LFZ1j3FAfNIa1SjrOvUg
zp8TkwuEgLXBsvBOaOkYjUWPdT8TKbcC80J0TIobJNc8q5j06VQEQaI8Rfq3zy8VBv5bJBdwIdTk
QJQ5VzNcgvMqh/VrOwJz5ZHeI+vRYXveNeMzsc6uJNaQz66sXcSGIlUbKvC0DO4TDaY3kPWPTLfE
4IZeTp4lmv5cdqf2BVeeuq5sceEixrE3+lIIUxUtefaudWiZHqBaTJX6h4IrLyI60SnkHo49KxjJ
GqFbzz6yXwu4ncDwWf1DVX7KtwJJ2eg6J/LA+ke89xtWQUkjeV8KxlIAWCJPJYcef/e8S2RXrBVT
grv5vcO8wGqfjwy6LZ9ZMKacGze9/uhwchjQ95C2CPedEoWqfAkEp3T32sIQkUkheSbx91vMjWj2
R2nhHw0U/Z6xOgusz+i3L7dSEL4vvij0ZXmCGL6C36Xl3/fFSstVPWA01Gtihpxjllsa3V6BaUWt
+UKAjdH4j2kT2TZg6WbU9oYZq6+++A12ysZR54Jw3mSSwc0qdc/VDqX2c6gOdYpDjcy+BvudaFCs
eGlpzSYD7N1hvTIpMFipYjKe1J4PueB/vuqj2fCZ6mEi2uE+juPQAnJyU35VIY40h/0BKhrg0+IZ
j7wO8q/6QJmzeb1NQBR17ybv5CqBK/nX+LylIvUzsf+TsS53lPCgDS1zMQDX3GUmffBC5AGDGG3t
3wMc/Fcfc4iS6UVcQK5sIwsxktxC26Uo4I/1aw3mAjOQqt8YRKsDZJrdlTNwFpRVnvPNqmipMuR1
Wpp+FRAFxJB+vLeMc130MUUk3/4CSmXnryUTCvCrfwaZ0FjzwKoGslxmlI6Gdm0bX+f58XOhpcmX
WvKa2c2qkZHbTOEIkcA4+hsHfxmU8lXiJ1myG/aQQvjjPyeRb87NaOTZfgq4EsbUS4bPjxVex8w3
GDRsT3fagGul3VqwpHOuLmGLEoI572TLI2+InSk6QCZ+d5/nRk4BUuqsoX/M2mxqjpDPkvkuunLw
n1DkU84vMkutflxkt+ShGRa6I2oVmtGhOZK+ZA8kxV+RB+U6gGwmQjCWjVz+Rg/EcbCAUPhOGWBO
PRce88woz9t7QDVfPjOcXyksctqi5AqFLHMP9rZCsWe5oy7f8S9dh1oBjZasvHijVpgLGDUVrgB5
BCYUlRXmzuikuNjwvxWb4mMLUAmhRuAODkHIjmuQYXiLeY5PqELaLjtS97BTkgm1dz0HYY2c27Pa
mTqm2BzQiaiclSOnnm5v19p7iQ21hZEIJuicb6HXpEpbKFikf0+9pyvGN9k2A8QGWRArX/C40/xp
cNTv6Q6hc+wp7I86/DDxnhAIyxhuGuaeAbpqr4RerDweHK+CYIxrRQNBBFOD882lZfAEzSsO1ozo
d/9/qlqqD/hbKKeV0PP61j16QcxfROiW5zyJRtETHW3OefFjLflf+Qx+adG4E1sF9rrTI98MYWYI
YuILoVCTQrb3TAZ5ZGSRTu78X8q2xel0g4je+cgL9AOUxzBziopLUMK2w2L32S49sdJw836cw8r8
tg6TNhnllNlINgKVbON+5qCtU6XOXT5spee8oEn/LkHoYu2XTe/E4bqOFGuVYyZ6avhJjPGdn7Sa
D/p/gvtCSER2iWJWeyhxVCB6q8XB1oBrtRg1Wu4axAnVCbR+F1gQrysrhfE3PEJzW3khLK5Mmljn
3CqqkT2EUNz0QqzPSR72c7OcMQIMGAZHuQCTKHVqifuMuTtlPphEbQ4nWXnfAvMdaQe0QqYkTLuC
yDrN621zPRpVtVIbTFdd0lnVNZtr1C1NEUA0ZRvZeIrM+PjWWunl6v6T5voaSxglMP98VO2SA24l
+YsyH/VfYMrbGScAkZ1wmnzqR4d3o0zJSPdvNc62XXnI0FHBoKctH4rHYq8ObuWtQW13glDdcWr4
Exg5vJtGSXPSr57uaX9eWOKXYYSFoTgZQZ5AjEOto/JW9SgI9naJlSN6G8QeqDlt7ZFuZLvQnEKf
L6THK88CnvW1UgFKOwjJvyjKIJmiq21tWIOlhyHITmW/Z6hdP+QvMU4jnw7vreXvLHuaf1rTK4pi
iGda9fZWmdvNtI8l6yflKC3DoVBZgQWmZrzqDuotwq9aea0oU1tj0ItXrQ/1cEZ6T5tZ8t1uqrc/
WOmGI0XoLOkdQJ+pO5D+qk2KEiWXahSWaY8gVY8ILWq0ES9UeHbdtm/Cxey69Tc/67d6sYps9JrH
+Jm5jgOWtQR42/nOQoooMhu7A8ObswP9qOWYejVCXAasUn+GR9xMfynitWrExgX359KDYXAR4LPA
eHMqFsm2gKGer9oXWphza4lq/z8sMfkX71/Hp684jA+cQ0dyRcZXG9BQ5bI/VGW6tu9Bty6Mtdp2
YAFeBnSyJPQK0PRBht7A1o6xRmpkuRESZn850TvZEQE7zeXIasFaWtxoxeD72SH7Ci7fpeI3Hz+t
Dk2/TO1d0hTWQpzfbsqSABnfWTBlqA17TTjurSU+RRnGxa9lcyiJ2tcHOK7lnIdwhxrbnpuZjxKE
2sPStAlPqErAJX+tyN5LtqcCoaUXOzNsO5hkwAjVmvd4Y1S77v7uTL1wSVePAUyYpQ4BxkXSr8Cf
n9pQmEd3eGOJhv5fJDcV8cXEiLF5lf22REhApV97dnbykUwnrau1cIMRmY41gjK9V3cvDqHpCJaC
fsZD9E5S0/HDyibyP/upGPBwszpppojreU2ipcsViiAieN8Nzz0/Wq65zsW356+PzCyIzF/gGUKc
F1ChVDBNnK9rbbfwklUELoIkLh3rCrmtZubyAG+t/ans/nYvDXOn1dxCZulnqPC6PYa2tssxlLZU
UQs8J4IbSlYbWg9GEgI5WKw5o8kjrBtMTFBF0zs3GFzXS+vcwd7q74Fqqu5pjPl4tDojSK+3HWQo
ldmw7GhN3dgwfMduXKXbD7dP8fGKLM/j1NrelxVHsRFejTgfgB1E3SyTepqXKlwKPl8XSPipZY4c
LXJ3jQfw20Yr2ObsPXKUa2WnAWTpDOj7UwPH6y29EAl0LXbSEj5wMvfgD5tWbrHoGp3JCez4jlfs
UH3H1h7K7che2POnXtFQUnlZRM2TLTY1+E7Q5CogMcUkkvz9H1Gm6/eDMkLxyR/z+Pivtq8iYNt3
M2i981lLgh7LebULX1fPjh6ff+k9GEQimwzfTQpUxe5yCP+2i7fajfSXClou8K9jHDrTaXf0ZR04
GyGgyt6lsnljVRvtRUCivla+7c23Cd2a5Eo2asBS1gnseHLPAl2Ab0HepmjPCXXYEk4YJv1JyAhP
KpcqgdccjTFQIJkvkE7MIvGtJ7vZ08Pa1jt4yFJmYo4+LxoDoEhy6k9tGvcXlXKeFNGNjCQIqYGw
ZQJitact+l9BmGk4TbqbJxj3OzjlFWw2YIePO9TfG+c0r43We47p1dv7BoTPZv09K6j7A/ghPTZd
ws/JC+W3zzpZxugOEdUdofRILKmW6/1r2P7fh9iziucQ5WHy8cM2dsPYPgokBOuQIjWYbf7AFTwX
WuKKinul6aQEhv7BdDUN9oYUSOoPSTsx8mWA5EMP3+nOojTTjaQhOQML5gLYh/rbT1kUYQwDdrR2
LTKeZBiKTNxUzMhEusKO9IhRMhA3QdVvOWKqNuP4f/oiwTy+k60penmA+HpS7SPkl/tmX5Ju3k6K
z0wsL5HlCeVzWKbJhZuWugq9nFU/SpoIyV5pxEJvc31yoDkb6ldBO2K/fgrvvAU5I1i+6fBvnytf
a+VniidKlGQXhNj6eA6ETkgMtZe9JC4JKV7PboiCW2YNlZXSOMXFeVZx0T+5Wdz5Y8OEejma3y9W
5TUeLIhyjB9nL7hsSxSj0wtZazYpKo5sFUfhBNcYBFLxE30NuRlCIIfND0TJYrODigtkiyg0oB58
PMnXohIqoWV2QNnIpnDIsUK+prUtEOtRZjtQgOos2nX1IEayZSVIXkU8oX6L0QbXZXC/Y7Wp7+VK
Z4RRMYeQYpR5bMSBpp1erf2OU0RuufpXGxpSPbbxN96ONcAiWugD+U++d7hKZMOuV1eCgeobmr1c
+mkqR1K6TCoGHDsUEq97O49laBziX4FR2/JhwXf4crg27aZ8G1ZzTir9qtbnodvXTm9cLCdMEAo7
OML1tq9zOG/Vw4WNI8FJBgOMhigeV/9+wUiuxV0Ci+AvLnh9XtLdOObVbGRY66TBuSMN+E22tKO+
6LeGRUlZVDjN6/hR/1LTfYLfvFXnFhfxc38lomWNGcnBX+sPgj8JUWK2zEZGQvucWqsfExoiR6hC
175KNsQlTnY1uXZQWtYAp0efYjtQsgxj5T+lUuGAbZ/Q9L8oa+15vdzUPeaaBLirWtV6TybaVKm1
0P/Iw1Y0i64NaPyTYZZ7RU1pg5f+wQLK36FU7lb4z5EAMVmrNqjqyGAYIDqTUg2mugWz+7iJ3d7j
lNs75m9VI8O2jrzLPEhTFi4dJDBRVP+5L0tlC8Lt0x97AtSzEchF/sMTa5qSiTJ7P4LJADilInSx
PuGjSdKYHWbio/lGcUPPW+cISzXQNQQgfyJxPsPuraAhpRThjmvSZJvLg1g57GsePWfXTXCIy0dE
52Sgo/xVCVIRKeQcTS0kjtHYzi61uRAajpvV/+B6BcaZCWF4Bx/ezDR4PBA+i5SEdt6ns1z7BeHX
jJuT9oaJKi0lXR8K/GU7X3w9MRR2eYb3KyDj1sntZZw4+heG9XpI33zDTln08/TSoHKNv5kKYu2z
Trt+jpiXTw0bbwBWROV1MMvb/49Y7MnUzXek1XikAA+Ex7BYLEaL0RhP5z5TiI7+2259pLPl+5bV
immbsM+RNT2m8MScTnDW5BVGs27MtNEa4/BnZYKG5bydOrzDz3gL230iRMvo+g7WqRU7D5Q3ng/v
sFEfsyLtjTNXB0ZA4lSNJcpWuPfkyJJ/CKvW0xPrlLbOBKmuB20IlX9NTwp+fcq0chjhjdBgnxEZ
SaFLpf3Bwu3pWQg3MsOEwwpPrtttQ5dJOfeSXz1CqNzjS2+OORKocjaZtzHXkRla9pckNRuVRp5K
Nzav1+T+C22+UXwNA1gs7FleuxUZjABYlGFIMwpTWWuytHJEu+q38SylrLFf3kyrwnt7oW1XGq17
CsHqQErATjlJNaMNG2Y8nUjD5IR0po/eay76VWavIiEjAJHxscXn0u4+I5pdB9YXKr/x1C+YHSiK
W2NGAsGJOxFdYFJPYuMvHAsqFHfHNqTxP+Z4IDpXCiBTGAB+T1cPWYrzwtgB2X0r2YyIu0zOIIuo
cpTfK7r/w6Ej/tTYKjraVoXaQwTSV/1ocrXmy6trUBoceqz9pNFpGNaebrH6zQtyTmvz9z9i5BU/
RU+tlm0UDZrXJSuSVu/mgUagemUYXSZptTFH3pej08ZVOY1vXS4IqMtyca85sCaCQB07NNq7XYpl
/F60GbWQaJsm9KpSklTFKXJ8cwQHDLk2TKDvTHbAG1bDPT31QnFkReek3dNwPmBfqlzoVsWZO644
psuOHw975Q8n+8OFPAxSGo7Upmw3okaSByxZD+/M5VhOm8cYNQGA5HrzCSfgn9kfeJa2SDyDuUr6
Dw5viEi+aUqmiQXA0rjKu6wyFSOmkDcVh4GLtw6uvxIXTEF1RH1jcGqfjuCAlmqWYB+jriURqXMo
FOpXggd4UHIKwk0loDv+VbnhdKJeIG07nt+gU4Ov7meER07VMIezu945f48mqvj786nKHc71754Y
RwKCe1HElEIW8Of0cDRJquNInEdv9nlc0CULYjMUI+H1Ex1X9jlGOjIZedAH3ZMr0/CEsxkJ8kwC
nfOKQf4N/J8N/ZnZnvPeHI1D/55/jc77nD/u6xvI3+rJddjJoNB3jA8dpkj4NPFJxyPgmeAG59rB
EWlJp73HwGjKqhTVpthTgKZ1hQUla7n0RAZQNNuPvcEC9uKXKwCKLXvc6FeLl0ckDJCCDzy/3RvM
uu0ioSPgOocIc9SQkk41+3DQYPHX04yAAkmW/7rjbyZ9p54bh35akmYegFUIoH22LWcT0XxmxNFH
zflsxuKhH3htCjGSZ75SU4ai1x+SAf58yJevLCO+0OJOjIIuyBbE3MM17I7+l3ziiyIUdK1ujn40
uwFJDH2yWPY5MnqEpzpzcphqfShhFywS2BP6ntq5i41T6pjrckJ336ODHyfj9i6VU52yb3Nxd9rt
XpsXn+kihcP3yYqxoLs1wEsQvB7CNH6ImDffqrK82LciqxHLWsj+stfIKTRYN8eEY/OOB59XGa6o
e4V0v4987msVcbVzgpFExrSst2Bl4Ok/lBuFtdzJjkkPflYFjK167IFAes3S2w3jhuX9mtEABzNc
5LL2Lyp23SDTWFkh3AVaaoN/FwO8lvoJtSw20CHF/fxoqBEpA9UxK7SsjHcY/tNPvdbDOUM5b3BH
FOV0ZOu9+cozFl9Uk6QmEfsldJGUaYodZ8PXyNOLJOuI1EglHdFFEDlUbos93aUQ/wv/SD73K5Si
9yBbnWLWI+fIxqfdgcGxOpcGFvAp8PxwLgKHnSJZhd8S37VYD7+TdUJrtT/l899Oo3RGPSDO7Xov
spp49FyY2fUodl6ALcEJZ1/I+j/l3VjO5yMCHUpsU5/hoaNzszX+00ovz3ZZDA8K6BB1b5YgL1As
mQ4BisjT7hO6Q+PPO66od7gyRFuEK7hTdg8hjpeZLKBqY8s2HDp5t8fWVCaAVNUN/9k+Y+j1Mv9T
B+sOFIsN/E+7vQr3uwG7CGgJdlQPbyXHGEy3EN3BmXXE+8T4OWvUE5fzxwvZSPajNiCGYZt2vu6x
rftBQa6pVwInKKNRqIZ7K2wvN5Emgn3sk8uAcR1yH+ZEfHGukpACERimkhMYIbqSS9259t28KU5w
CCpZH94aRR/8DpsjzK84qGtO1VWpAuTkLo3PDSybzL2IXn7ow3yVfR6X8weLhM5AABkmg7CXwpmv
2lu7l6H0hq0DBDevB5Nibn5+JXQxH1KeQI6sUg1q6ziLq/8m0uOrJGAadG3QXPSaCP3xNJ72qD/U
krDjYVa4TBjaVnX92wMbblHBzkwN8y9S9nsPuyS6D2fJLmMTZaTs9TkN+nqJ4R5kbP/x6HqDph12
XGCSkSIFLdbU6GILKZvjIqjWW/ntGctVvSpUfg0QEs6TGnoltcWS5PVmnkAWTwN9oU5Oofa0uSax
hiNPAIRsEPl0F5tAIvAkf1xHf1tyeHUsxA2J0VjkZhi9YeiCpOg42R47OPF5Tx1/9cK9E/kaLv13
hUsrjUAwqXTivis0pycdnNWhSARip3Q7fcn1x1H7YJrJ28pzD8Hfk7AfumFxEAOLce7nklHabgld
KkCnMKSJIAqEtDDIzanzdPwJZz0yiNk7wkIl+aZuZ0mCml/1YL61D9X+uefyr+wAzRDh15oEKgCY
Lin2AFnB+PROhF98B1Fw/CD63xoQk8zi6Cb6X1hcu5qyKa5u7Wv5ojFnip+MQWbfwcCVa8ebkrRO
LRGhczBV4Nr206wNZNbYzujVgDYSsUfKyos5UtnqdROXt21chRb/1dqfbmciUp6ou/i7CD0nIulm
8ha0gaMmdcuHlU6ahYncCP7qmDYiTKxiWmgMLryg+3hSSdDwZ9Q7HPdJWQh19GBWrMNGRAUGmVDL
OgdF491f7JyCpzgGbM0/wvNITXVibOhx0j3/EF6XtdZ9DSRF7O2j7SxDQ9US2lC/Yc8CzSFIELQ8
YnvbM2atgJGNdliqiv4irEapIfw2G/tfjL0rAx7ct3XK3T2d00Ssum4xUNf3fQAaeZ8EaRQba4qK
qeJ8wyEWJU+WDtVHyF+TYRB9WKTjZ4Ik3lXhS0PujDtMvBwYbt2iiWzQh2i8O+6YBeazF1BgXV6o
xvNsYAqCey8o2ee7B/bzJTeMCrhgi4D9+DHkY7uYJEHQABUgG6ozpHlRQv6wf0vMkDbKP3nYVWQ1
6O2U0/Gb6lGlbkptn1NdMOXu9WoqYXCpwpRN2kJTJ7c1jwpw6p0vuYHO4TANUo88ScWuWnXQ1pvM
zMTd6u4YmFwWmrA9p7sHNnf20YwNflz4WARL44YuTDxIYh3lhZIbhSZcFf5TBgqDqoCKU6EBiKe1
HOWmmkN+3igegTfMEufVvTOAheaVgetlfDIdLOsAh9xzmbw7iz8B3WkS7wgSzwUhqFsmaXp7Ee8l
FXDQRHKBlApqj+gb065N+lsBXwTiod6ZIp58Ez0H9QtlP5qhWddV7ECBAtAiRI4HhbQ+KT+z1lEp
vhbDlVf/RO2StBJ9h4v3BFHrcvkTC+Wf0Tth3HxCVZC6GJz0q3OoYJJWpz1QIBnH21O4lD1B+lrI
4DgROZOLKq0hYejQYA678dZRYd0TQdxjQdhstSXeDuNf8yWEWHRFIMuX2YJYxNrNGMDgN0QJ5mcB
1G5t9ZpZ3ioIXD9jwJxP9XNjNbzFJF7k9SkLUTVtyLmuNbRV6OjeNpMNIFhoAYVusN+4BjpCy8wN
gTbsXeNPisKgCBlauVXqQlKoDfXVejMlRlVFeIcdaHQDzY1cnoLDDUqnfnO8uGMC/X7x2hyWlrzi
f373hN1KohoWfLTclF4qF7yU5I+txdwzLcxjPthJPUDLcr1gvmYYk85eAgDiE59kWIBoWr12ddt4
4gg7gqMYB1Ml2zxxB1qBhnB+O3RkBWNcskwkSR3Rh7ga9QE6eFLOfKN/+05aKvXk7VJ3+0S8H/jy
MEo3K+KMjECp8fjfLmiGMohREVBNbHpwSu7WjtFTT11+qAxHuvpdhFscHHqR+Le9B32pHfHDu4Fs
/q1pwYhLFJ3fDKaTMMhpWByA6uneP5xZdbC8RETTZfGruRTCIQqi8rX8f6RFUzbJjFK40vNlwEHD
f6rJohyhoj6Fxtz8l4XVNoIa5NqEa9BU5v8lQrxyzkMeje/RnspzqiFsnr3/hiPj0IHwVxKgfXWy
NhAJaoaZhhYweLj78e0QB7nJ3TYVx3KXP7aVrqyblrsnXZwEwNeAsKfvDri+cf7Jxl/cW6uIWhB5
Sh1jqn4I2tJrSgU0at0sVwcQabBxo4fkxFIP3jR5KLvjCdgNQSwgFTqpJkZcDKnVSDVGQPAn2Zm5
awkpsoNxDnfVDUjAM4QLHFp7iaGHHwGoYKOdU3oFCGux6bbl1sutdOkIZz6v/3JKd8RPoMI/eX3v
CWaQz9LLkSkx++flC9oRY28/rnvioOdjL48Rklivxlm5D8ptCVdm+qj4/MrYNTy/rw1Su99ArIIp
Zgr13Ek3iOTtZ0A+Gt2ozbs3oaOIg3vX/gD5nqH302+EdWY16AxAYUZC66N3pMJttIDw5W3g0fkq
Yu6SzXhNpHc+Ikkqnj4x92/FnDcb0Xv1AJrEPgrhFKGnUXmAI4dw7FN6eOJHsCz9nL5NEHPvpu2g
+hGO+6YrK2a7iQ/STH2tdqSgrZkfQ5pwOJLW1OolR4Rq7578dIlu0GuOQxDIIqzIY1UfJ6ghnyZ4
jsk2hOyNtpNR7isvDe7ecw5Dwc12e5MCY5th3NFcWW6SFW+w173bGsPQdRo1TvUChUFiD+robBnP
RnGqI+5ej8AoCsRo6Ue7oflV9oqRcd3xGvgW92qPH/8cDtWJgynaCtK+bMHetSt9FeGpHlVk3sua
rIE6VfFx6jmh+lxogPPTWbEw/yeSYRulA8voUaHI+A2QtjtxVJPydZrNhftic6ActP0kCB9rZ1DR
aYicbiNpqEiF7nH58bAE71tlhV3sddDhQ2BGALXrip4sgxgCyVTJW8tWARvdwkHyZC/DWLUc99wx
6fSXZTUu5E+Ij6+kDcvELoGu1E4ZU6Wd6RyfSUN1u71UEQ00r4SoSLTyToHZrh2rkv6W6MbuLqUG
Qe6pl6SUGkyDLPOzH1PRlirPiI3dghn6EcFugW8CrQi0Uf0Lgan6fyq1Px2UMzStfyjRxa3Fd263
UBbnBxsoqwN1oXQ4NmGxkfZi0kWYTfmcQkMtpWUoZJ3p/z9/Rerd1qBYIBKqEY6eEFRF1OHsX35M
KdRmil4XAagZEFbevMvb1XSKfq3ah7kupRGm+VEp19Z6/XlMkBW173V+9+mUDSD7e1PeRg2NhCoP
vm0Wz1/b2z8ciGzs+7A+ftsS6/b2DYK5UAtHjfW5MFQmgGw4K/c0MYkd0CqDi7SPtTlljJgP4UHK
1zpJ6w8KN5QKDXjInMCrIh5krsZ6yVNIMKCd0ndn7juric6pwPqZVMAJf4cYI2UvyCLVjFs0EdP5
zeRzg5P34XgKiF85qLemhLNnEKEjCOmFK9rJMI3ZVFJeW3kc2PEUrdQ5BdAoUJBwnwR0fGta+7E0
q/MwMVxout+uy+vpUr0Qvf6bu7zrvLYMTqNSvPl6r1pZrtyknu4UdXpO7ODL2X4fzimwj1UdYsDX
ef24RLwgvDDcR3M8qkvogl2/eXlps/d8R/w/bzQVNmkeWOrgZ+K3kZmewVVu73j4THmnflnLwOM7
IahHp1qTQBYYK/UcSiLtMLulWCdEgZ0Ei6I3wBe96OLxDkf9mT3UpdamMc0el7+pcj1IBHH67aqR
DiXKBp43/1Yyoj0g2/FKTcXCgUszvvBf+jiCC5Vdqx0ZmmcywYnT1hJuZBgg2DUyRn5fByKWw6+S
BM4Nn8+EAbxHrwAPdHfDu8ud4W+dH3MJxuMU9arePD9D+hefY87ZDbDufYpGd/j66wAbxP7QbDpa
z1FBR25Q15yI774tUr5py0q/ew2/TkYfeD/WauRMHbdVuQ7W3Fhf0OlKibcm+QjHblPYjddLO8XL
Yy52nK3zCRuNHvX7qi+nyvx1JTUD72UK8bfjb5V4VdGu4k1FEQl4ZesLBI2R+2BJJFrgKgRGPLJr
JVn+9TRIRXVS1Nz4aCNZnfNIaauAY8ILJ1OoceW129+WvpN+lHoh6zZkSLTSYJAOFEOQUBNmzahZ
kRJ+sKzRrRdJu5Chp6nntXd1dPzhOcQOo9MGvMbsY+Q4w+0vqWeuf5X+QCkKV+jf6+RsG9x0tgUp
ZIKyiIq/ShCQ1F2cGvVdsWGJpTrsLFTPu4wuFGgzk8vdVisGOePPXgxg9LMul4O3Bjod8h1CTE7x
08Zm9jXHxhmmRVxVEQx4vFdgcPCfSlEXr+J/M50S+iCJCrwuZRRj0ZGJjIUfKlO+pyA7LROgrPJG
SYvpfSrhJhIqVsbG7qi23hKkx3cKjVFXoUP/zA8uLYDGxNJGhDTG+ZKX6haarpJVIXZto8egB5Du
ZhqNd8Y4TMlLGGsW9jOPZ4z55mUDkRXQH01gAQEFx9VImv1HVTCv+xUR0Ifr2yLIoUfB9OacmjYc
SoIZGJcvoNVMW8EC57zdVGdaF9b8wHEOKqMZG91/rtRl0xvq8LDBoDmtRPnJvM2v2BFxT5N6TQPC
JJ4AFAZ7+bAGqHRKUzNeGGt1LNOEGBWLND5iL0ZW3c9L+6CVBEKpV+elT4xRFEKsE+Jqx3j7ReYh
L+5f41lfHMSfRfroA/Z7cOoZ/Zw+fcyKu9vlQNOP8J2Ulj1C5F+IQPR72STmMhlSab1RjXxU69bL
fWuYzM7p/oUtbVoSj5kRWIohBWXz7pKi+OJKBcFp1EeK1mhuaOOf7Fs/fYTxfgmbRUVZ1XXEKmg7
HZPYWL+KwV9npezCvQKCeyfBlkvAqSIuESS+VdLHiDgcyCZxBsjDCsWTlnNukd2wAFE5VohDzNkw
tSk3Cj9BMy1tEW6kNeFjrsg2OJ6Nxi/XbWsJ6O2MZhWArNDGkW2vjmFa86l5DhfM7V4hqvUp5Heo
zzbYpQlCxVVBBroWBGpPctoyo/Ql5aN3EYZ5JoKUwfE/ITpIpxgWxhUk2vIg65FhtfxLm1Z9BGuJ
D76ekkUdoJZWh1BEFVY9X7mLTNNj9wG/ea9edlTFI5eZA4ddmwX0P7jdWMeZ/KeCgxhUWUvpcbQm
2k3dPjlLDTdKMB8/SQflzFFjGFBuo69FB0DDlTxcjFRkUra7iUdyNITEeZ3zLzskt9zGA5YaPZSu
BmRBoG6N+jWI7yLY4ZcUDmOKLOa/mDq42McCwH2pXED9iFTYuPvGoQKTqRAUjt9xdJq6GTaiDyEo
3zPqHYFrIEgV7ary4MOmveA6Zi+bi0JFkm8UdegeYDiLDsc8Nx0kn3Ne0j0yLAbKnPfeR15CeVeN
zZnzu1T+ZIJ5ZKsF24UUyZRlbsp4CIHqstzVe/EEiIOrYsgrAWJ7F4KIY9wZJrBCW2hXIIVrzXWl
A+QdVP8/sM3CuCBUYhdhVXBeNLmGjlUmAXnmCFy7ogAtllUnjaAi5eacYOQ4rt2IkQ+8QUqmgUFB
sDA0xiRJsYKFgakh4e5A0XRvKtZWlpUTIZ3w4tUN52S98vHeWXRsr0Aiy9yOvnOtU1IqMoc+0/t7
pXn2O+nGhvHb43WegcGM1UC51rvjupYp3+MsEYvpecsnOVa5wOzkn8nTJaAmWYGr8zlmh/6GWROC
vPaFTHUYnuSOIyb66kQjW5eYjgT9NxX4M6eCDMYEGWqOgUINr6CQDbMY9uIWNj7QavojK5QrDjnd
kkg5YhJdUvZVChxhRcNqCzM3zyPbZfidco+0gWfXxjtCluZK6gmRMeaUDduZV0izJb6k5vqAjqdX
gpkTvmuVXKl0k5S2jQXfffHlZm/dpyJzrC9BjlScmvS+ZxZroUsGujD5Ir0eI/6gz7bpzi6kKWww
mOS/ZYBx6smTz25X6MZkWh1kB907tYOGFN+TajXFRO09TwxqRxgg0jnyq2ze9gwMWRVZlXHLalzm
PcylOy54zhVZ1IrlC+CFtj4w8P1/lQJZUOG+dO+O6pI0QuJMOUrs7BgLETEgDs73OJ/5UU3U2AdV
JqcbLbwDCWsbzCeT/uMW+eC1LV2Tg/10FDqLOUqc7tOdozrfB113ig7kbYJ04w69NdlUq0C4k7J1
FKYPE1bOrjWPGnf3agN5BDSP2qREagKcewdPL0rexMzaHAAZdyWFi80MTbRQdbtGEjlXZ8RsxrdX
IOnElmfzLjnr+sNy8NGf//azqLDBUU2cEHfs6VZ7lRpl/Jh5c7SWc3s/w61P+qg7dTkzZdFLz4os
Dfll7eCXpNJYQdOpg/jHqOBB5lLXnlc019mqJ4kRAT9wR8Gz4u8oijxPDKDjzUD+A3+0lY9gcIer
N3ZZTijVmOBYxrE7KIHc0LgMu23tFYHAg/scE4Vc8LJYBWPlM3IIPHTaneSFWsUpG3w3+wxHA0uS
BxkNaU9/qJ677P7QHlG+lc/aJLl1eZOx3BR+6ABIxqZenE+2RSIzYrtyOLDY/D4hba9SWrvn1cxQ
tigmgHpokjRqn38VMolekaPzWTrat2M3vguE88saLzsNFpIaj1LwRGod9ESFhDNfZldu1fipNUEU
O/zXroiJCWYIcwm88T2PJ1fLrD6iDrh/lAcnOj625XtK+2TjUv0kKvPO2wZoMq29tR1sg6hNvVb/
q0I/rKY6pU3VtvCwYHGU0vIWcrPdDlY7iCbxU8RggqVetdInxEDWVZG2qZksx5uHpueSUWi72re+
CtGqm2AqfxTDTjjAf5qWaQYUXTC1GKXaIMQkfuxPvXMazGX/qgodTaMLcTJFpWuy43eU3taDyQ9A
fotzmul45dhn/BqptcMR8L50sd2RkeTeEVXWBN1i+mOxgnpF6ERSmfNYayipAzb3o4T1fo1RNanE
icr70smuxZbDHl3eUKHue2hU9DaHwq1h542lYk58Mhv7QmxkDDUq6/PyrkwWoSQnFFHU1urX/9rZ
f8T9dJFEzDdPEkcxSTIkKBK7kuohocn8ddq92xRo3rNiIfD8auveNZXHn11NLyAlngL9dU5oSYuS
Wp0vQLwtCsro7LDJBDejCXYIijUvHhVK45q7eorfgFJgogL0O6yNvdD+b3oFhIOH0GUnSHUmh4hm
L9G2jZpzHNWMCc0XSUhV4DNadzi+FWAtJkoBnvwDg8at3H+uhI2qeJZJD341C6CbOVyhA5dW0sAU
pNyXBupg3BSSe1/48ndjv9M8cpkHRC0VTHb/Yfw5vWubHdhMHX3aYrttfgCzL8cW9B9GIY48eL2p
trYVwaVPwv8+QvVsj2VtC32p3iI2s0Iav3Yy7unZUv8L5u2AtqYTxgB7NzeB1do8yToubXR23iSN
+QEILNCE1zOh15g9uIhWlzSLofJ2ljwDeCmtgwwSQfwh80nNhC1euD0SzlEdWpQ6V/kKEMT09KxL
v08FkXRJIyy+H4zJ+DmKn5gnGX+qwR5ZN7UlLfK5R4PAN7kQIV+tPYGrQSC+nrOgOXyb8m+aD3UF
H6OzaMP/pZMbrIZiR7g4Q92IzcFAIKRcU0XymTpt4I4EE/zFPfVmzBP0f/J5+u9ej6iknGxc1qcU
1zWmc2EcPNWCwSiKeroNeERYHpNQ51TmZPlDEeidwkLbesMy3X6PjoJIJ4TqZSTxSblhotcFruSp
RWu8XlTSTBRZV9dgLe12PcpvMOnadmuLCBkJfA/evCwoAKRhInEiIEFhezA5pj5NpXGEilP03N9y
VP0Tb4lA1LTSKNPRbYmfS/lIKztUdFbhykJeADhHWNxru/pbiGvPcg5wDZwOPNFgSqMYStAsBWV0
g0miqy5EKWS5HmPCUKM5IeWsk4z1fEXap+XIJbSHoGIycPYZCxvOjj1xZfqoeBcMxRP0bA0tuMrG
N05Phgpqjme3LsVEp8Y5KXDlt8BMpaZig6sHvJAzQkkmTfsB9w5wNiHUtRcrYEod804y+gJt5zyD
S0dzeA2B/gs3Aa56QTKnjw8o4E/yKR4joxmhIr1rNXRe2MZdPVRPF0TnYoEHW/sAqHH86tCzBwoC
La1myNFsjc4Xr/tgTCsBGmMSl1Vfl91cd4dqtcQg4LGGTe3CXLsD24Xe/tRFNRKIPkm91Tj3fMIB
3t+KDdREWl+PeyDSe0Cir97Tan7myxX0BeCTTDvuHkY78T/8mX6NAVFa8XGZoPM0xpVn2i7Qp2BV
ugfgNqkS1Chbuu6M66CCT0f6AoVP5NlG+i9W+gUKUw3xYrKv+t+cbCP42EWb2gxD8kgJOZqSFGLC
3rTUt8l4q8zKoia0TliLp0JNu47w08f7S7QAIxEEx17HqkuQeVa/V2CEekVD2cwyU4qCe+eKk/fn
8bbu+6fbjmlKLZCdPYkZo0oTiZ8PSo1JhOPwpsWjvmj2kKrSv/HmAPhiuPPXAwyyjVx3ma9Ez1pp
znop7IBuoXSvFHLUlDpVai0/D2vDGQ7Q0UxJT494tCI9Ki86Sxw8tqC5Csg0lSCTQ7Hoo+eLGsLg
EYHW2iRDdb8HzuaHfvQhrzPWOkRhX4bkZ4EzOKtiPfSFxC7/LaTHvaG/pmJ4gwIo4ARNeck6ESiQ
Zwt/gBzraZExhB3vu0/Quz2KT1kFhnD0ESmJbLe/vcLVFSYi+poISI+df+ZsZe0e982Rl9SGcGYA
y9C3TcEwQ0gn61k8SzHFQ7w2NJCw0mB6U1McOz1hOVbqr4tNl7K3uN2QJlVVHkWaZ7jvxIPE+sUM
lOWWMPZeEkWrFAETY81Y51SWSITN0rQjnojA2Ca5w+S5lvIp85SxUAmnm7tiD/di4+FfPx1gshtd
6xkX4c0I6x4TFJt5XNmzwWSbWi6jwQMkFZRe1ioAoxTt4hTAFDTtp63d8Ct2iMvdzPD26iTgYhKD
JfpGzqi/eC1MzOda5VnacJjw5nJkP7omONLYqhyek2trx2q/h5K4KJhzrZgNWnODJUpZxuVZx/Ig
zQi5dwSkSyn6S++HdKe5e269N8z6gMLbnH+pAiFhcFQcvdBwbaDyVByWS4ZqRBRBe9csdDCTeMeK
bYrAkVbnhYXEGhzExlu9wr6MIuzgmIdOYA1AHqHrJzJV+LHe/iHYQqXtV8mfSXwmzdKvcoi2N62i
4oyHqIAgNVq3+HaZybwumKjHVt0Pfy+GTk+g+T5Ek96CJQzlizjLx12HjhtUczGYYiwKaxQ/d9+d
UzpfSRe16bTe7D1idN/BzfcuZYeBN12+bEe3p/cvjnW4d4lRWULp+ld4iEvfr3FvGU53oZkmjvOX
WhKOfD6zvm5GfjMjHPj/GNmbvEGVaHcLynTWLnsxkz9FcVHhlG3ktxIrUuMCDaBh2bMseMYl5RWK
eGqFQUJnummVnZCIF1rI/x+MfPPd13AXdSD4qagDSaX7hd/mQkVn9hp9TaUqrLiIUYrWdfLFRl0H
s3KelhAVT6sNbU8bwKHLeU9Izd8x4nfi6Az3v2ebUR1Qtho95zTrvQfdoWSEln0F7XTIfhE8pIRg
NNM6s3smqewOgyUtw0pfXLH78ILuNVZ709iDEW/7fZdW6NjpjoAzi02IxjIMHD6F/T7f+3tiPrjY
/AtV1SNfeQHJQzBIDNasQRfUpedfKSBbkts2748FoxTnfAGLFr6wg6CrTWOMRjSaubVhiADpkmAl
2OTzHNbi9dlhRUSPEoPtIXGcHpkk3k4TItnY/w2OXIBpL2jgf1FOuCt+4tP3nrBJqtzrPi3UXYdO
yjNIVHpV7Sm6nGYNMPzM0SgsUM1x1cVsJ5qXiU07ibUQAPawWjOMKhfqO1jpwaZLO1cil8l193Ls
xqTU6DB3r6YiTBOFMEvVLrXgwaZT00trw59+jvnxFiztRQX7YsKRjDC10ibnZFPUE24Sz2KwxL98
9N7m6dzrgQ+u5rvx3UlCAn5I/kTatXIlMFPg+HwQBxzlkZkRReFn4WjOBrLhKgpx3g0g0jG2iD6l
s6VCnSf+gqHaZjsu8ig8TKUIhuKEn18VyyWGuB7OszbpnfRlvitTQeMrfHnuK1QWePl/62hX6yH8
ueSTJ3qmlI/qDE8fWrE/P+9z80Ufx+A8m71Va9BahrMQkNRRe5Ni4bmubk64/e+M5sFelhHUfK16
Vzk8tJ7DmqsomfBaipDxht5f5ZYYEQbSLSg8TDYnESG8ZBy25MnCpX9/LhNh/Gr5d49DXio0/ogF
bkdxwOYedelsqPw/1N1zG8blITsdc5FYL+wXM+/74JzELh7s9t2WdqNx/ao8djGbokPRsAOaVtq3
h0n3i1p30vkCwrXbs/ou7Cr3/anCB38cnKEM1o8A1euqPvLc/75mFMQEoLK3seE4ds+Fnypw5wtK
2sxdtznfr4Djklm3qaiR3fIofSG9TGAU39USvnAEQvSv7xJoFOl2cnSER7kSAAr3IC2HKIL/B8vI
1kPwMCeXreLeZ1ZAzv0bUjw4sVcAs2W5qlAtr2vIvRXjLiHs5A63JXlrkhR6v0uKESiFxhAmf75T
VwkYj3LYZ8iAAgCIXvIVWsv9WsG+5S5SZeFw5oai7uS8DYDFySVwYoX+GnUB1KrmCS6EIasV5/zE
qz925lHnSR+fMeA5UKZxpyLY2UarywxYDEPkmtAqRuJJyE+9uEHQiWP2Zcy3ZBjLuLQAI0wdWQD7
Yj+72vPvNkV/CGeYoZcUVZGwypuT61p2V3vI7vC0xhW2v4CFqGFBJwOPNlsQeQMfjOi9KO+KKLhx
VouEImqf9RZL3nZBMhg3tTsirOc8iha5j5PzqWCjPPIqjvwljkIbb44nWFeCytOlJpIahJp9EtBp
TCO0JvELO1dqq06T9DntSiYu+i4wHc3fXZDw0UYvTY+0JF2U1g8s0veZ7tPpAf7XTqPl4uXfW6RK
YRgF1iJ3EiCtyvpPzE/UUbmlmKmxhyohf3PVCJAeJFsnby1hbnU4sd09lY88R9B9WbD2ADd3gp7j
dDH3FXdmbMn1r5xaLNOG5qFRnNEGEmv4NsN+VJBduWmejCBNwcejchk+Z0gI3q5zohvC7dReztNN
+biYKULEUWpoR/hPj8TXKAvEqD4VONXda5bK8+cHEo8X4tAdfbgjbiMNxxr7QpaJGllVtLk263+/
CsqCAlLALtRif8zx6jQ/1UpNj1o+AmLcn1N1pjDTR0gM4o+eteiDj5LTkpfM1ZsTVf5b11xOQmOc
CPaKlczNPc8pCdtKdhCMqqXVajJnzlIlR5vSQIlLnCLiwa1E8AQqzyNg6kpDPqSDNCFiRHVoxH0m
4q5P1BOOpvVlPVC+VESwtZnqCqT/MSC3jLTNIYq0ywBrnf7RNrI+amuP6v9rxB1xR6nSDtfHufNg
llvah44WzlEX9v7BRvHqyWaLtFqJCuTXSFQHwXMHaRxvgHmJp7pCL3cm4WhKlEFSHPHhuIwiV0tJ
B4GCbidJAHQriyTw/lEwvmpbhtLIlRkdFhegAeSWIrVKtY3NSTz6mKPEzfCD+VHfgN3jlMl8+HQX
bNv79G0v1JvN5kFxrHNzGa92xCdGQYVjiCPKH3tUFN49mCwHWaFGcjy864k91IV9GdV6RmE8llzu
m9avNr1+i1BSXOuQ2D4C02y85sEXmrL9tkmJHXiIXZeFNgAa6PZDZEihDqnBHDS7SJYl48EUpc7l
UB5T5s0wDWB3NENk+0Qmsu3q8UjqEJCLJsmQ4QXnYFYnwYommdyHdiFhHFWBLTdOX93X6i4CWwys
ZwRkrdaHG1bgms+zXr0h4BzNozZwJvOJGXfdVkZnaYU7tMLsh0d+r6ZEqtuqcHf0uVvAG4S2KiqH
tEzxt8EZUeeiuIKWRZabg2Q3Fo99+SyMk6VNCHx+CFiVJuUG5CzohedrR7Z07fQA2GX4gVs7a5PT
LV4K62hqs1YDu3YqQ2xN36BykyQxy8wlXQdQtQQMnxvk+UkGRBqjZFBl5T9gvB0jMiXrX0+OZztu
xmJCFW+6dWuVLhW5ocDa0E7wjS6gFqhy1XO5zDGcUwO8TqPk3b2GGOx0Qh0tuXOcGmHZqTghR/WP
YrBuIy+dlHR/tEh4V+iH2WAl/KPwmXCQCzpE/7GcBPWhgu/bf9I5zCPdD/AmaZkfjcnJZOSNL9jc
sATmw+c+zyHC9+t83wvnMfjyRymT2z5zXkNLl5AohuS8xG+FCQRUUhk39BtgY6sgZqaK7kNw6A9/
b6p2vuWZOuu617UQLQhnIFr0ynWY1kFPpsZzzgMNMmDQKkLkTEUH/xi0wsX2ONz4dsyYdDeveYXO
PPhvM9uWZwIzB9AYF+675w67QnZTlkuyVfk+b03v3KCanvYcUXegPZYHCivpYz7S6CdZeCi1ph+L
CkdBS27FGih5QBmtTH7jilAx0ITRuGIDsOHa6ZVHnyZfl4eryxB9IKotDmjyM/IpnsI5frviYua1
Q0g890ndJjF03SGXtvRTv7gmwXTBWX/jfvzs6nVF+AJ/JHKmOXdPl2dbYIHlD/XiYL5sIgb0U9Ul
7qHZJ0nDjlp8xpHtmb/Ji5q3lGKYIKyS1SlkCzvX43+InAcZQdfI36ZlLQejhCDRA5HXb/h/oldg
Vk8rPHsBCD/QJL1uVhITo+8iQUgyJim26t7/JPv+UY8wQn6D8ipZe8mkU5EMTk7c4UGSNiWRfDCO
u7MaJ8s6FiwBlP4aZQPWK8BYXutkSbEhHGjdq6Wfh0zdVWp2T6qvyPWV/P0GcKzN+loVyjxDOomq
KI8ZiafM/zw5kfOzr1cPmulSy5yB77McIpwbDl94sGK1KIZD7raDKx1eanUE1+nHGKwNDQuP5qWK
MhhfQKt8iRmRi8fooAoqzXBrJWtAw/X5CCh0ECcRG+PP15DzYJVrSbn8ZA7yfMz3NzQNiSY/PV10
o3AObIQ0EXq1Fedo5SCWMKiS/uQ6WoIkQ63zSNV8gyhkHetOY1Xh7V+smGK21ideH7orPi897yKN
oVEk8hiYLnnrwZC7NkaC/j1MbultbHWkPby0VF3F+PBcJmo+OZeElmIr5JIXBMFST2Fxfz11eYoN
CShL0hvGryYU763VtbJfJSEyPYiEeCKpCtQPhoJokJn37Z9kArS8DzonBGOBgfFH70Wt8lKwzkZg
ZVC26aKd5l/1Rg+4G3ZhIS2dRO622u0hoTSqSgQLP2soSceeFfGCn5AlMNbngYBqeu+Ez6jxT9HY
BsEV/f9eL5mW2Ga0nH6j0PDIW5SocOF35FG8MZuh4q/yIVl+YW8sVTV7T1jccq023ozJfUH2qU1s
3UF3JoWNsbLMqwiu+iSRg/lDqAJG2U/jEl80eyYSzB2zY/Qolt/7+o5svWETdHNX3DuBAeAe3nIr
1MnSxwuEhudPu4CPH9LcUrLbdD8mwVWkFR7aybJrHqAlwkGcgrN8Q99lpDttojpYtXV2pEC+YSDy
5ZXhHrXuH7fUf8+dGMtBUIrd3c2hE2xgp1tia1NupMgt032Z+IuEWmxznKYeY2dj+7SAg2baTGh+
kcwahZQZdXfesvWiqehOdBB8TKct2itmyheH5rrSK9zLNZrrDU2MX8nDSHCSTGHBWaD7zrbKRFiq
m4MkMsoT8PqG8FFZ5YsN0BvEY4y7RetZU5ksGbjTPE2j4NSNSAh4VV5Z8so5gqEY/Ws85His5yME
bm7VjhxRO6kC4nTSc9YUEJbOAzWt3SaPu5Mdn/LTNdbdG5KLtwHUSuMeZh0Wu2SiY4hzXaazmBFj
OQbJ+dE81x/K9XYIYR/0p+D9h4Ige8F96C2c+CRLvOCe5Sq6KznSiAHGWqGlwIoRJHp8QcVF4SbU
l3xu/3n1y+SmL1xWTd93naJ707B+6xTLqa+jeXeqiuHhB/INNWRGmle2WDnSb0AbcA/ntprLk3yZ
lRLDWc5i8bXlOb+D0rjgHLhy92ZdBwC2SDzvKXYKv7QQXnwcVu0FFDuXt7kP9PF4IpTGeFcJchFU
4m+GNTMiEaTuhXUmpoiAfhWOcp8ELh0rSaofY410NMBFw+yHnjf1nAzHkyawiQEj6MwsGq0lXe+R
edszT7Y9CxXq1BI1if1cP2/yn4DKpqSTsvsI4tD250M6YWF2STEulA6VlLr9Oc62E5o47fkf+XE4
n1CikxoSzLumpOOytzMZUZxQRTnlJn0Ro963GzHjIVaIUq/ia8+rhizDB65YIsBbcfnQ4AyH4wR1
1yQnDr3keD9+Mf7ky2eFjZUIoXAHCAN+5Ev4h4eDWWWouEfF+NYVRvxbxlnjpO97MKpNK9t8fE+5
ncOur9XYFp9YR4ax1Spw8pPapysf+CdvI29RyydQB61nSDdDLSKokVbluFjESoEOTZSBZ4BlgSc3
33ujdfNiQX94DbF3c/A4DyUenwgFvOpyDuQVjkMO9UOnHEWEbtqL3VkOfVw8s6ujqJ6zn0j398rT
zEgrw12czlbgb6SAl33bZdWXYbS0Ouq66Yd+s9dEF6HMVfOfq7G3VI27+iBgQnktUjKWn8L0cMyR
BLC4krjTJyP419h4JUoWG9oxo8Nk4x+7pXqE3MEFmXvzD2ZdY7b+kgD7+P2JRMNKwiyfXlMRbv87
Xr1sxYIrY23B6raa7B24+qFGW8zKXQhValtL4W9OnH5fwK/7fD4AB2by5MnK5geVctLwaL5jwN2Y
7eDfHqPYHu4d/7e1P30dCrfH9hbOG+Yt5ELQrFaYywKfPjofuRfP4QfRtau6kq1uGPQLPTnl3hYT
x5ipnevcq0sVfWcsNH6dPJEZz2JQ+TK6rR893qd8LpIrwl8J65UYepBM2dy94wIOTG/T1URypPuQ
mo3W5cyVCT0EOgQ6cTmlcNTJa0gXoHxXFTwlAD5tdCG1r9s2J3gBE9wf31mslVx9LwN1i9hSvpDI
29Py06jmkSZYBdDw0mC2yehXbll9qa4/wHnKTa7YSaUuSbwIFZBUwYa+0T3JmZ5m8RQJjxv9FipU
foBvEavQ0hUavWuDn4XTXvUazLuVXAYLoK7VoMHITfUe3hSHiyqDAjuqissb7SHC8DvVBv6Fdhts
hbADvN0/gy/UhASbG2SFCBbhEtoAZoJ5+yGUDPouUcULeaxDHuSQZmXT5C5BtNXwMd8I3P+2DBhs
8pD7fss4dRdoRd2KiPmNcQweV2i8Conbjym0XN9F5F1gkLi593nw1+MHJfPGI/YI2WQLEBVLeRfY
pyTt/i08Xu1lGjACXe2QmaHAjn0zmt4pdpdmKD2V0SwsqN1ODbuXEmSL6JEcFUA5eon90gYaK7m5
a2z2ITfDqFeUBIelGjExcmWYD9m7+6ZsehUiHmRtYp9kkcFY7oCYRIYlIWW1dDrzQfehORECfbfv
l8lIUcBoRsrW+Z06X/CPQLsr8lWY+RDapl6mQPrCs3zzIOezKrC9Nej72brOBuYaRgxjabVHMvfb
1h16V3TK3E9nfuSU/v02vc+b0qf8JCiuNI5fYJY+j/P8uG54VoAIOMoZCcPG89coorLj/176sVqx
2PNX+GxoX5Y4c5r0UE2k9E1dlCGFyJsDclq4Oa2fBNt84blD3H5KDIOAfzU4pcvXxIRmmSeKuGZc
gLis0/opOMQNPke3sj9xEJFYsK5Df/w2cgYtsKCSB5e/QrnbCFV0ysmJxUALXX9fsTP1lPR+0OcC
znZRjqiND1qETf5xeGxDqCSXF1MkyS9vXaj0tuMBBwGMiyrCbPBcy53HmBom/BzvS18QRyuNADx3
1kQ9j5Ck0kGWuXg47X+rDVW0A9gI4LIOtlGJZy01i4njjEoqDjUwnYgePAcw4iArYqrHkLg/XE4Q
4+RW5Wz5VcbVAgekYlDjDTYjRk9TX0TFvuq7nQ7tR1MyYzsd85MVeK/sHxBxKeEKFZ5d7OfM0PSm
UeUxLVS1eaF+oW9bym0Jf3YVlMWwtOhsCnJshIKa4t5i7KIHF0j70F1inhlF3Sxia4TlrroKNutS
RhMweXBcxdsyn1aX+ooI8RWyVw7L4gnNl1pPDKJb7Lg/XK1Q3c+7KvL0K84BTlWT7cn6coBZXSJo
SGiof18oi9fo5JaAqs0yzDqtJ4Fw1rcSeitCrJFjeXL2vXl9Pzsijtser/KJqysJwhBox48Zho7G
FEswS+d//rfCpz4A/DsuuyHCqskg4uWfsyVsycmIENIK1XWvCHcl3xxQ38YbZ/XTxdjrPQLtPDWA
sJYi2R9Zcin3ggTYHrHl4Pz1YpD4JRx37ZCuNq8ih7E+3IafCDmOy3KUkf/XCe+9AqXJyJRR4ml9
FfVFVglRQBnm6lJOMPXEDXHQdIv3ROBvmQkOMPA6QBtMPPqsS1b7AsoJbGjpbwG6ZDzJlMmh2oYJ
4gGmj+0fQ/SRwyy1dDMynm2UNsIbDtZ++4PnftSyTWV0C0pfJtRo+B5guKeNewRrZyihGk87V2fV
mW+FDq1kWgg46dTMRwseBX9JSHQJVr+DdsyEvaQyEj/kKF2VUQvIOJ7fuZ+n2/UplvOzFvREVgwe
mWFe73K2gQf+VrbX53X72c+VIhhWRYsO3M5WiKcnWCe/c8eGKkqWF6JxY4FlK0EDzW9yXamWwtM6
7LaUp82DnJrd4oP0bzQ40CAZrCb5YuUCfM656Itm/6rAtKolBomNhXtVAn8GeEODCAqwo72FyHfK
lzQN6GTfKym3CEsx1hcWh5zBZAWEJ/ANaOGGeHXYeCGgQj0k+EVVI+shGToR1hEuC7e7riIbe1o1
QCBkscp3nmXSwf3/jnJ2sHQBPzKIwc2kDJb9rGTTBdWWAw+DZ37a4u0gidyFw/P1habMHEq7tkJR
6h3H4G4KyBNdzeoXF47lOWLt+ZiYk3SKO7NCH/V61gs6syDBW6Dyaw8WAdMc/raY8WTzE+kO7SZ/
6f0wWP4jKoMSy9uh1xuM05IrL66fefVRVu+g33Ur1C1h6XDiOSVyvKmv7IftQwmsRkUARgD0Zprf
WpMIJqT3V7Ism7h7Xo13SDrMu8e5hqbvwy0bqC6VLlDpQO34mVxliYbPsEf5AZhPa9gjNfSy2XEt
8RIG+LyKN2eMaxk7IBxU1EpKT0XQwYuou/iYzYE9jq+e+KFNjCbHjwaBzuh8h4wTJYVdTNpwrEz0
8p0tZPGcm7rz74U+sCDNu1Wg913TWQ+yBQ/3XUyxf6Frwkitji/oqiHL/tXXvO8bOWVlNWduZa71
NLo9pFwH3hUDkYD9AoPf0wnsa4iqhBSqrKSHsYpeURKuce5uUEz6PC93YSfbnFTfpnoZOBy8q+NP
bL2yyfAyfs7gT486lXMlvlFdEGRbDALvDKQOU1Mur4fwmW0jzGOg4gysZ0+k8IpZMcyvl7+or+xq
T2gAOsHphZrNSU3aOTVYjQczSwLOAHcQIU0O+PjZrWGnB9a+SUsWxwfxwyfp1zl6PDmtR6ikds/a
h3uTi30eEE2BFwcrPqlzyV9Im++jV+umjPdXhHfJb6Dl2Yd2vLmCzrNkNFqbNwnDwiodI5TDSsjh
0kfpqjALH9UDTjqvnFPHWjALXZljKTZRs0js0dFBgUfwRYCDm5zYw10JilBXo649ROBkDMfQ+v9K
8DNien50+GR7KjkosfGTIPK88V6M54LffNYWVcr3gDJrWBb45M6fLDIZMlcbTT4bGqyiXnbD1IOX
6xaTA4lyXup0Do8fh9RPUxSzi5GJgJS4W417xzJvIqGnxsH1Jzt84MrdZH+g+agMxpQ25Dccibua
J7Y1na+lRWsR78LiLjmPJGVsomRyrQK4Uzn1by9106asm8uvQzlzfgttKrlbuiYPzfxh7xaKlens
nSMpBk1UA7DjRl9A6UjqRzemsKNKiB112Xz46mANtxK7Oh4oZHdzdOHzTnRYExXZCZR1R79qL612
hREyP2if/Md+C5Nnvw893jJGDs23Dwc5vgiBOManx36LQsZCxabKl0hA02hfBP0i1WPQxTyYbypx
pKWl1CoWlZbDacgXYdAmXwTODAiLoxN3AB7woX/1ZofmDyUEKP0gkcSAQKAln6Tv5hAcvot+s7Jl
+YsT04tap9ToSjDI+SYn4+JhG6x+DveaVqMnjLdk9vy8PpNjXiW9zWKOEXXMKSrj1a4vJr82Tnhy
HPRQeaTNx/SOwzckJMTHOsc1uS9CKg1GeQ1MIXDGJs03eKr3PYXw96w2Zg+AjXrUe4hrMt+Ohu5A
CmXgOHg5q7VtqnxLOokdONADho0hIhtJjnIsfnVLFjai5kkIB5J79mGydaXITOpcug6Sie1HDsjh
cvu0ArBPbKdKdlciA9lkt07jUSQRBUhR6KHYyCxpYH056RhuzbySHLQtKpUJR517m92R5BD9TDFI
OdACgFXKoSu8+j3vZN+74Odn/a45qjHZSSGFW4mRi5aOoY+GMV/hh/DysdesC29JipnS++MM+PPp
CBF7StpoQD4pJGJTkvNsLPvYuEUhLeLx+gYDf9iolM98jq2kX3oezqohonAQKDbroT+alLNQzBCl
r8eZOwYalxARjbViKNrqHRWUU9sl/wleC/vy/eH3L31Osc6fLMSxUi6YFJnXhab9G9BDaBVYlHkN
kmAYAhbxyg0+YVhAiaDyKdfCRkjyPNV9ZHSgqT2beuTGWjspna4luZ3u5XvbAEcfjaD28jV+5Fb1
P6+2S6CmId2Vdf8WfBD+nA9iCUaHPNL2Vu2eO8VYBUFhQQzxVSGQk5omiSc61QWc+lWznBAeNFRl
1o5GJwa6YyHEd1kJ+IlcYreF9OKVnoHQBg7md/PA18aJv8ecf8C37o3GjT6CkQx5tEsIFDaQVe7s
yg8t7Ugu4bfRXc0/UzV802cgp8anW5eTO+ylbYVOe2gvpfcqdt31EDNLqKcNRPmxp/KkyziF0Eeg
i3mVrnKsP7Le1mx/86IWZ9vTrSEMSTdcvMhSE42vhXYWMT9m6HRgA3I6pc0cwae5JexYaRreemUF
ZobE5gGaqxRLAY2IIpwqpnvhN24zX+hKN0TGFqCVbtDcULs5YdtZR8UhLDHzWp85UcR7e/z2GF1E
8/lN/kmudrpdEy4zMqjaSSmRjgLfCiKOPNUmTH6ECiXXvnMAl41DffcZJUlEioGn2k2VsCcMyd6A
bYASg7vxueDf6oplfVbBYtb4bQekXQTZXmGVN4gkN3WN+tkgwUe3YskvMNA+T9OrTowoutQromVK
ecQ4Jiwuli58XzDqJGBlsFE5OIuoU5kcaxd1x3JEUepn1rp5brKQgBZtALbH3u7UxlqFykbL1qid
aTJpQt3kGpnbWqVZ2Uo7cyLHXL2YLC1h5tssKFmIoYD1imOJ5wsihYnME9IkX9wVRt3gbixECEDU
2ahxV5aZsLAAW/NabC65hjm1Ny8gbPbMoiR8/kZj+mL8Jhqr9URGVbMRds3gnsQ+9Yv/ySXIB9oP
0+d8VYdwwfHy9OZp9FNB2SfJDFBs6pqMhVDQBz5MGPN0ViMADda8L5m8POcjoP73/QUDKszLWNQ9
3IB0oavxHo36qvTidbki83+ZknLXgbT5fFG1nWgPfu82tziUQXq5iJ+6A1vkNm+oNo0A+qHcqYKw
ITnxfATSUCqN4WEgGCyUtgjL9DjTDqiuAAa59EuT9Qi3p5/cvWkoPVHukZ5QP+EttoCOT5S/K1k8
IkNbi764DOyjkOpwKy3bbdpD9As6rW977A6xrYS22TBBTWbOCefqJShCUzXK0xgqQ8f9gQTCfDxC
bUoEww8FOPL8v0XCFZrPfCMirVq/9qO18NyfrtSTpkiGCs14TGoah2qxfIfhB10wAyRYHs6CgzBQ
fbJJ8RoJHq7nUfPhMouh9MtLLnzc61q0IuaScfNDRcvebDUdDtwBX255MQ0gBwueuC9k5s66iJck
Sq66DDE7pxxOzfha9KuEcoXoBuxEmF2G2sHy6t2kQTqa8g1f4xIViab9t5ePYdeh5n+sPhw0vOdJ
oXHWeufhKUPibYK/UKwSd8iSnzShIy3BeJoTNO0Ro+ky7XwpjbTn0jRmnMmN2PET1UqdTywPZxO7
QXuBf4PvJNWcVba2sJpiQ/tFkn8s7LWrHlILIRLFdYK5HKhMrOfNDH4js5xZ0yDsPhkiz7QnB/KK
wcoazZGVCc3tmROeGmyLUoViZMiFL/hkm1iF7uQsLlcfKZl4MgC/pUn8lKOlVYeauYu8NTh/FS9j
txo6/yGcgFg/eOy97aU7mnDbuDXq9qI2S4IOSWCXE6YVsuwYDYXaurVF6Ue6Q6slRQr+iEpP7AVv
vIQp7cU8Axv9S9AlBVsxQVlioAA3xbd95+1jbDhRd6sZaj4tzujLUr4XG76Z+aJ7C0B5EkB7wLXp
DpD5m093BFinOgKzz4/MqiAbBNsZhZws8kNWvNmhFi9YUqXy4/tujgRZ0N7IyIRqxU2vhJEV2tHZ
X4/Ad7H3dppEmA8FDGln1m8BZRH+JPrtS7/6WHbgDI5gWMaWTX242uCwqAeeaDZQRIzclNaUaOXi
oCW23Ca5/qoDZFRd+uiLI0TRlzAP2LXxwWb1cnsa/o6siIouAsNdd9+brvFCFvsPKcTgEVZ90CQZ
zVU4DHuxF3Yvy1ZkiIJJRR3ykXuTdS92HSsnebXlWhvapLPZP33priJoMQw0V4Q4NDYbu/2Ritnw
77Jru1/Y8Xnl13Hhruijo1QVT8+cB6yhBoiADqT9Un8R1BRfcnA9uJ93V0uxukXczlD+MMymH0rd
COdnQESI8+wuuTKdn2w+znOdPnD8SSvlznRrrsJRIDtVG7nenpz/m0UodVjdxDeWl5hlmx26f30S
WvVANoX0c5li4EnAsc0LNNaJX8p2GgPw5XexFtnVDe2k4RfQ/b0pXoRkHAnbonCm8hBWW+n4BYg0
BrvXT+CUcwARBg06xc4q57tjQBeQ4KuEIZ+n7Y+8uC4qKBxsMO9hezSoWdmCTixcP51AUiGPv3w9
RJEr9p14xHc30R8xTc7Yy/u8yqir5Z+EIrIOHDGxbBTVwAhIEFHRC/OdhI+7MrsB05onIjw5X5nN
2qXaCE74TyW2YCUSqL7OH7wUnvJn2KcsmmCxxtU8OZcCo/P3creuYZDuSz/ACjjtoeZ199BS39UU
B5vHIROEpjwWVq3pvzvt6RkmqQB5wbz/judI6TKi280yhWe0UHxZTzZQrnGqkZAoGrjzBKQn0uVd
F5ASRLcQIWgL2rw9ZlELbzFAQsGiKunEZuxihRc3HbZZNkSAQ9UDiwtyRrk09HMEX8gX0b06WVjs
W7y7cW6oFMLjA1pI7rUpN4QB2KMWY+PsAH9pM/uVdAKIM8shRRUZkC8P+y/3d35QIy+Fv8RbX74y
9zslRyv0tH8YT/usk0ZGQDVgcVCx0btDQadTol4MT5zPcs7fIBqxkUX4AwwB610r5+2Mk3xk4VJi
x7pEpaASNqjCA1W6mUtghkJNcv4flm6yfXvqxu9CnXOLlTT/3Hcjp0kT+G+/VWNj5ywVBMxfyL9/
+eOKw232A05N2Ed33Y27ZzTKMVvOytlUrEhHyu4Utd0HLYKwRXBzUs4W4LQVXsnc5OSc/hQEIVhr
iDF5LxeQHGeoqUOiHoTvdCPGtttIa56Aa/e6CAFhhmqjVmuLyLUKX0Lc9nFGbqkMe2wN79xxpsJx
PAt7mX2caXI920+B4rEpvFlMNbXTA8k2jpO2kKv7kS5ltCDxFUg/woEwSyJXnlQsFz8/2uCQHkH7
DBD267mazDVHKiJNvJrr2F9xBtRJWb67+fH5OjEb8I+aJuRjt3xGnbbPYTLpZMgeeaJ5mGLvYBNI
yphdOQfhTp+Ej9Fs+ZFMUrkE+c1MJq9rlQHlVIY61Vo4ChSqlhCANXa77zd6S7ZQEJ2VeKlOM2jd
6koV7rYzzOJcdld0ty62nrmoL9SYFjORlqVw2+HcQesfq+Dhx5tcSeXSLJTcU60BcI1li5tufdp+
1y5peedML/Pp9UdIQRbVgHG6Bd5uNWH9bmy39c02xGa8Ge4K+TzmZwBUFM13M7GUFJc1ybPD7ZGW
9ceARShr3pKE/AQllNM8xnCP/cP+L4ceLlFPkhWeNjpWK/3sFOTQb7QO1ArsX7nH+kOj+5UvCG8r
tXWJ5I/9Rf+dqMBjhbZ8Q/J9LPnhdwoyKqmaH+IQJWyfjX/iSswPskgZfWAU/7m6QIA5t+JysJrC
1/RgUHAvjT/UhLKkk+AklUaWXEBxdpeLakHF3+4Ftg23cIdgS1UgAylxbAXLdekuwYhp0Utxn776
M7QWWSGAAIkFlvJgNAB+ybMRydHyjwnEFamKkhvwllpTjLcT103uZ028EpARSt2+z06Sez4+hMph
5ttWuog83yjKxlElWcTsHTBMG9N1MmfZmdvi2O8/c1iPqEiLXKUjb3LE8J41NLoXXR6QJz11jqlf
0CkOssIrzYZGAJFVpYNPZuk1dFfiUsk1YRzI0uLqArIiHagmFBKTRXkSz9mJIuogT6rzHlRuGMhy
ruaCt4AZA0xHbKy9gMNg3aLzrIcpMLB2YUfpdi7rO2HWQ9VhQ1insnLPjYJOuvDEbis/h2xD+EPN
3e+mCSgqhdEhcxdbyMvz37f5+8knU+8Qp7nYeQTy/6g8fJJwLbNFkS7FRMG1tnacf3r+ND4DyoIi
Nss/SoaWTi45H0Kh2JPoSrpMuXIgjbR0/JAxqCEivQN4T7G3FWrgexs3HnWlin2XNEa18XyVOwuz
Dni4/F/UGaEOU2xXOqBz034xHAt9+ZZg5gOlew+wSfP20RXB5TWrhUrj1udtJgTNpezqBLbW0XJ/
vaeAuBdK19DuuLsataiqbfvdnHNimLdMEOtu8r4InH2PplPnnMxagDz/AEC88O1RpaFlEQy5wvv2
CrHR8FlZ6afePk6kCHiJdWj7p4xMHtlhlP0ICG7buKbUS/lHj18aJm+hB5iKnc31hoIerg2m/JHM
0QSCQTznzCoIckgCkD9KPPcg8zf95zz5WearjqM9+dC4QY6SjrUsugLARMb/ncr1TDVGTpQyGJWe
nYP0QBkBOuL2xbk3RgJlv1koUZ9N4EHZxxPdyXVPDKIn0Bq55dFuXr0fpOeyipAN3ISld5Y/yQKE
VOpk6ZXoedvsMBP4vByUDrfh4QPs+rQecYMv2SKqeVWm7oUId0A4i7yww8GNfDcdnLymMF9Cjkfc
tAzY3ssZ9fEQmlTrC6yelnontuMe9XzfcQEK0u0if3oCB/dBDwoIVS+8IjFV6w38Qfmo07S1o59i
bwTUY04rPHOoStf19wnXFdilRrcrCYNHQr3UP4qsLT97uKwoODJ8DYLykJEbfY8QywVy7YoRaMgR
7ZTnYkCMy0hLppyxXYK8Lj1wFR5SwvC8lLRaZeJ6IuiORON12LiuwhmI7MFT3I5gNjp7BJAR+uag
gh1MrDgUlrFZwrehPUORl1w1BuY9omWrX5pvCfVpqWT3gvSoDLjL1ff1Mbu3CcxCn5hqtLsIoQlv
IwMvxs25eVbuG724K/wEAy6XquKm3iNhSSOvc+H7SvM2WC6sLINbk2N6mFUHjlgcmpIJDLL5sOqz
4CEx1OjjI0VMCxzViu6PQ20xlZNdT+XrfTHi5bcLQyfuouSybK/Qs2g/T7NsOD20YspQqdAx2x1m
uL8hKfsOWxnpWLoJf/WnlBeeoRrn79Ckf+PP7/pUG76dk+JsVUevtRgLtFDXx8HbOBCan8NfgrA6
OmGMnr+khCZCJiL+CUSfSV942E3kI9wP0b9okXtx7XOQiRFcziIP4qNDNc1eQIVfR0k1ns2P0C4o
56DJt0EE3Ftf2JUzT38xbs54qxBzw5DNPxw22Mw6jrzhJmaOpT4OIMWFgbGmXAb88ICIfl7yuAd7
2z3ndcyBtrdjg94ELSjaDD7DjSwrrKhhfpi2MK5/cPkO3G98fE3E4bmpaAU/eU8QQzAbJVnZTMwE
Ndn8EDvx6WOL+4ewn/WyaU3cqKJHkat7p0TbyzO5QzKt61Ot3EYHdO+FAx/CKqmE+CEvlpbMc95j
n0MiVuLW/zA1yfPJLqLWvT8Xwue4O+Mz2ZzAaQbrYokkepoVb1U9y8DxcOoXF6K6oYkGzZ4tvGwC
fq7fLt8QfgBgpjqJcZW175MDysFeZ/BEuhj4klpe7wOipBUoW4tnWjbXjWoluUTTgEbmLJsbTZ4m
MRd6kIWt6rcsHl25G+6xdK8YWxRbsaLSvJ8ZgcPLaMY2oobGGaqRuNZDQ3yXDpa5ueQm36ETqDrM
G6sV/mAqgZ68h3wJpQAsKk4thyj663Eiqedcsi2aHtHZAqxoS2z1feWWD0T1vo4UJkWhg1fWVoNm
RWaUQG+JOfzfaYoammgzk6ow9yYXsVzeHFuCku/NMTSaVPUeaXxkzclmsT773xPijKK3osL3DR+B
LjDxVu9Fitk//XljLD/dLN1lGBhbM68OXVs4JnnjOzv+5nYqV7y804O62/6vsDjXFtJOvHh0Ud1V
KvTFsxxOuyajyIgk3l1A+zctbGnrXx7hnMmcDmytux6bSgetokV05Rcfc7Vqd5rE/Q76Bgd7Yt2+
uKoIoq49qs2cDhCdNyqtAKky77AZ49Dt8ZSGmd78ViaFX5cDR4M1dRXeQwFCAjny66xwHA7OD7Is
rajPufFK1XU13gctN9wlZoMBiO8T3xK9IL9J6ilyKaFdHgcBSctHt66GQDoRNYWrtnOHjzsSS4P/
TgjsrlKs27FP0Zn4cQnnmZAHxXhib1XekgrigJsYRTdXUITjODAiee30DBa8S3XXq+rt+cK8/Olj
teXAEbXTlEJbNHPjVoflhHi1jwbY1XkibHfKcjtxTnbr1U0aHkblv8nmTK0fPzfMtxNEQl0WdAF9
xvZ4zvgfmMhvRQ8pl3VxbBoWHq70/wo15L+pnLB1miEqmNwB0s1gWVvt/bjxSovuDLelWcEqo5Gy
ebQdDp9SPkln0HdEj/duq4x/9Xz3a3laqvsC/9SZqUUyVHriASKGkGirm5eC4i71Nt3PJVyp0GUg
Y0ZP3HiuED9goAO4dQ2h/GOgZSWOAjOzUbZvMuyNzfMjzdtBPjY5I2XYyO7hChz7Stp0wDX7rFIB
c/KE4nz6wrRd72lR0Tgow52UaDTnK59+CZ9gns54CX3e0FjnsBARmP4A8fWfQF6+bBMBtQ/mJmFI
jLo/H/TwJF/ueN4PTAUONTE1kiWUN9u+w+TWFAzYiPzm8Jy66efXKwQfGwbvSLyycJsZdSQgMsqe
mZ1+sUoLJlVlU8zkC8ArH7PiHmMpsTxc4IFa75RcFAO59KIaMArPcw68+QkAOubXiobInPbbX5dB
JP4L3/oiVP4Nby6k/eiudGoRzZvKdSka8rOA97qfGEwh4S4NqEPHYABckOzMF48i39qCe+pep6gI
rBBfutIv+nXyGsIcxD3b2hZ9+BdMjCBoRb+9eLItz4F/nKH3+rKDjZ3BBx/JY4QXMvM+XzR6JaDB
BSSiYGJNXIfNvROUThu30M+yMTn0Ngq6bxSCjHh2k5VbEudtXAIOlrfxr1OLKcKTtiN8Nh/v8f03
hTK0okXxpHvdPoHvD41l4469hQpJOv/U4CFYoe3JKL1WahdKb9gMtCrNOzhF+4ORiyHk0EI1gNbZ
M8P0y3tcjtvwqGHUbl4Hvg+zw6muOSIlKCb07jv9pm+oTJe4vq7GQBAGxwBZBLAKp/OhePWpdiIb
DHEa43VF5PHkpps5RgPI4kIVaQSR72AtdnXiGYQcw3Fcj8Zgaqy+te15AOqCqhmxF/MFx0EDRacv
dGQHi5uwqyzqxSXq93pGypy/JtasFYqOtQAs+dJTVHNHgzqR8cGUULLll44zaCllgaDxsNchM7FJ
mXqGBoijlIgc2f6g57ZQg930s8nLAIRV4EOVQKjBDUBar04oOobqidnunr3+bS+93AiMA2YPLkQv
Gb8pzYEifffUGq70Ez0H1jnK3gmbyrBBwo9CvporYwLBKwt1E28d/hFtfjeeOImBZBDhvH5tvD8t
abowS4IvZbHePbcYuISCOO34dJUiHUNbZQ48lggsfpqK8spvgWfFb88sGDSGoB5zKDejHfXS+XIr
5vqXdcyiWJYuwdgFI9puYMndJx5CqzRW7jcNIXoZcjrGHvvYQK9Rgi9pDLcXb5ZPJtCbWIxLSghQ
Ie5y8hMRkUPuCsJJCYF45msrJJaxIj5htsjfogw9lDZ9F5exb471Q/Ffb3NVnyNeYfhgMrcIlYTy
LxJHX/wmA0qojZTqqkJBSA0KXVlRRI/vBlYSKS8txZCy4YNODbOkOWH3tBr3A1kvPlp3wVzBZLfC
jbUoLI6fNTIz3SDRfjxWgWYGkHX49j7N3vhQndJbAb0hZf1SMJO0E1JqEoElbPYY+O7QhDoQVpH7
hKYWUQ6WVS7Z2qzEb1+4j2RD9Vl0mPcBccDlAwxPABSlhNQrs+32lVq3lXm2u2QN60yUtpRMuW1t
tCER2EBqWSxcER+je5T5jTQFWTr1PV66fVfnmgk4bgqD4hnix6XOLL3EGCzLp2UlkykS0zjdBNlO
n1RKabbrHsdK7LlKYQd/1goeilP8QjGVainN+An+mX8QHEkdCiyV3Rj0qyqe73brt+N8aXyVvwi9
hjSeznjrjobYXDzVISglmb2s6acwwPpzmAnvg6LuYaqF94gDJd2EiZY0nFbD4Q5JqFv2bVFCYp3G
ycoI59+SFIGuQ1vPKVcO9lATr9E5x0PHajaTKVYJY7hkO69eOxL8CGv8jLpc7IawfeDc4DrZrtjt
Us4/R57RP9fRn/xh70hyMUKlHdq2j+YJ7cxWhuuggp9JKFK08Qr67H+VrEFngTva/8kj1gNgmBTK
K2zi4wOu61b8IMtsuUWNSK697zR5Bn6wnI51RVtOvsErcDJaoz3S1GW8VVVs5QVHpO3uGaUTeqEw
wv7pEGVO/G2gejYbmnORV5RrZ3GKGN0yua9nExNMoorHwK6ri7YCMvIbFCh4qQnwQkGUKQP7vpqa
tdCyLD70bdFaFoXOcHo3SeMQF1+ORm/FmTYsZhiKH1dfZ7QjCyNZ7lUxVRzBORggCDOgGAtoJcSP
9M2UpqYmEM9g2unphqP2wrFlYfXvvjv9NeB85aOc7CWzFajoowZAoJr7BQC3G2v3MZs1BrkmxLt6
8pnAJ7sIhAAd7XeV8pYZG7pbgqN46zvS6eTG1ibI6yVfzWGGWVNJSHzmGMmyw8MQH9Qtjb+1ij0t
sEuZ1e/mhT0anPrGaHhHq0webpv296yfmDeD7aJs8vDyRaI8Mf/9EfNoeDy6QVFWIL+Z0wXYl5F5
D1t6fJOy0XqgcXrLkg1HPryUzmlAw/qVPZiyC8uL5r4+XfvgOmnc6ET0YFRaUH9/9WEL+a7lpIS7
ZTmxYayBvRL5H00YFo/vWORYMw8xFWLtNaZqhU4hDKq8VWbkpBvb96AwHt0v9t+ERask8NMLIO8L
dYGhOY8bPoQkudfFbQghpKyLUZtsFsIc0eKK+1w09KKkGz5kiJ6eOj6w24otw82t2w9URCk77gnH
sF2J8oSIwKg+EVg3BhPDIzb0ECnk6BFHdy7gRWlgIj2yVFBV2hvihkj/dWObpk+xHSl9TdA35Cy3
MI+VRsqOd+Nlo/Yp5Weyt7/4kq9hsKOLH/UM5xk6STtvLaAam91FbHWVS3ciy3wcnkvVw8o+tkLh
Wysm245vTQFNL43caeAgClnhacGQjyX/Lr5B+WQBMFUWaz+LRvl2xwaLDCNF2tUyKdYaT4f3ytjL
enkiNaHm53PfMeg3rl8sAlUA8RvKgTPc8eByJFukttBhDLn+vHj1R/wEzXnQsIQhfxl5XqTsgLvY
ncFlz/3MElQ7f+lYB4D5v9Q38P0bAlVeSnyJilN4a5ci2pie5MObrJH91TE+/lqrxw1I7kJZtKv/
Cirvf6qLIAuvUL0Ppmc02+Z02Xj8BZX4ssX005O03fotTcYKQMlzF0z/VtbtE0ddTP29+kG7EWHW
kNt83isggO6h8uCMxSmCBvSBDbZ4DlNvKcHYFsgwB4HrrCLGbJ9Yq+LZi5eXuxItx6iG3a3N1Qsy
8HMaTQkzT98QV0tgUmQZwjFujQi9hXwCCbQDToXSaNjPoS/mNAKAdfiYi5FPMB3e4h4RRppvYJdg
FCG4aUYCRZtBp6hTME0/s65OlKlyaqmHfU9kdm1ts0GAm3Y3FMMgZIeT+YSC7Xqgd857PkYGYYAd
epD41Qwnxon0FYIN6C80d3kWXkSUPOruYYPJBplBdVPyJCvC8n0jdCdxwOEyAPJVfxfKMGz9mdHH
dW7fHKXdjvu3Mg5veoPAezjE5SY68/efNqEjJfnJh8LwpSPyXmqhUI1/LTr3A0V76nAgSEo7K+RJ
IHgos22VudHf/LrPBRLTJEC86xuYbXJLTfZ00msUYioElr9LJX0mS+KGd1Lv6E5H1QpjrUkWwyrX
coJ5pga4dBVwu6RM+wv1s9Y/4nXdMO2B3Ohmi9QZEhnbhBUOgtOJ7eOsh3Djl71+RNllb1ceWC4A
AWJ2ZP7nHH3lABj44R+aWRVWOavingOR5F4lWmt+tl4Z8nOQThpKJbdVSYXFQNhiCMK8hSLxfBg9
zD2MJbTQpSCDB28muqMpkXS/SJJ1BKQZAy+wNGzEUqSI+F4Lh5eeJfLX1AsqEL0v4JStBnwDmaBh
bgBG96gyr7lsLiyxr7Jiun3QUG+mJh5pasKfRFxaY5S9ih5CpmGX+Fk7HqW0bESuiQk5MHB/hl4b
HompW/KsGZLeF0tnypH5UdRDYU/7zljjSP7oFR7wtTGg4neaK1MqQAmktj2lc//PZX+wZkenn8ow
G221GyCWoBovYVsC5LKA7Hb8RBciFfBaLahBeOVpI4b1CnNwCcSoCOspIzz3rZlVQ+DTUe/O3rOC
j4W7F2IlgWRzVRUlC2zsrmCFqTRnNTkqyW0aVuCjzxLs7XmMf1bxS+3wNMXrZuiPQ+EHfclqSAdV
OJWKEkCun8ArlLNH4rPY23nutLfR1cQGDRyWeCSdehkgFoSjS0j5qsI2e6tCTW+1NuJCNtRmzn7b
SsZN9FaXcOp26PYfAcGJzLZKQYF9aC5mbcbmK9TRdeiXtPdRkYlE4qadZT8RubyNkxhwEBjt2afb
XQU2F43HVIh9LsdPLBvoA7cbNaNdD6No93SS5pDQVLV0VLjg14ZjO6e9WYQGrrAL1Pth1Gk5Vf3O
FEgg7avorhn3uuVbfbEXZr0Kwrh7+w6l03/GQhx//OlgAA2w6cNqXgTUnzlQ2WWZbUVoddRAsCwt
5HlpmtJcwsIYZYNrY6LuDJc3hMK1SeV5M6lZpPmsskwvjhP037BGr9M7plIZBa1o9We651f6aDd1
bZtVs0TowCqMD/YHYah+Zzuep8Ma9QaK6Ze+hKXM+aqvyZPDWEZE1b+ZcUgbKHq74H6Gn2ybca4q
G9t8nTiuTJZCZBFaavBVc8nMXN2batBBYmv4i0blTZF5hvYg/YQKm45uqlxt22om+AMxTVwR8piK
cebzVYHvKcsOOy1XTjMWkpNQ/1KL4hlounC7zQEf2zk5tdlJzhUUcTxF9DjDXYED6UIGDb/XZGhT
Mr2Xdn0UTGkdbV5pRrKROF4h+kyJZvM7Iq/5s9fXVJjWg8W3FWucjZjyYkIgMGBHRZXg7Scu+hKy
LKc5+McydfZNmzY9YBDHd0OiyPnJF2FDQb47ew3I0JWI9rDIAE7GPrlCD2aEVdHKMgN+O0aX5Zo9
ZV8CSUM3CIzu6NRTNvvlEyLO++pXnQFyD7TD1pCcIfZ3z/91ahukFnhTQ8kEsmUSX+AFIUQrrpoS
jbLEEgTT2Ot4hT3IsLKgd0GeV9G/D+znvz6OKaYedZ0376avJsZDsG+VJ/+GY49EXiIXcN3f8N42
ACdRK1KLwmK+wkGJdrO00c/Fj+gPBViCAJ+Xo92SpH7VFvl6eOmW811zRBC0rQ7eHIeWKVjziZkg
njkdCanNERNvVXHdpAw0txCtl0AcM5vmJYljeARE3GevGD4+u2ztdvy1/lIE4T1Ls5uQnfxilOk5
P6qO6zkVshCwWGviXzoCN8cQuVWFvhlGhKuMTMYje8fiWxhCreHpmjABb4b78zgG7ansiNo7P+Sv
8/5TA2P+//Wn8JAJZC9rDjazkcCaZTGbB5sr9VAzJfqJuJDEd0yKhRzjXTQummqP06wnYAQ76cIE
uwBqIwkC/bOyR5U86Fl3aZQV9eMZRhRoLBch6/Osfqee2yiqqT8dicRVjsFHb5kzCqeFdzmGGAET
zJ15DrL3Xitj3lhbDDkbDxafZ/jmiFqihZ8FfQbVLhKFuGT9UGx32zD5bQnYcbcLUa0Fl1adPIf1
j4nNjERArUcD2B/OR49Wl6pWuGG3FTLNvkWfcaURooMB312sngjJv/CTvWoLjgmb9Xq+ScMoJOcU
sQLSbRK4MbAqSX6SJb0anspx+RceymdPnBbPyRBsDD+wJ5ka9RQY2Od7fD2WGa3HRyLSBwITsAx/
kWq+70vWI9hD8YbkdiGwnlkCu1fRR78mvaJy9UjNpyiPGy8r2lMqxR3Xt0qZ2gbam+KuutV04bMl
x+H1jUiBRiKY6H5O6g09Fp3+Auqd5H5yo1YZBLe/FClMXapnhGLahbsSh/FllMcRvXd/FqCENdja
a/J/7LAtfS21r+lh/hIZRpDF57AYxNu/P/KynPh92LK/HZaqDdeH17UXmDmv7vC34FtHIMK7Ba22
KYtD4/O5IQ8gokA9nH3NzA0gjrWcIBWCe3TUWGkMmcbFCRQqxzamaiFyvChsaMPXTMZEhzJhrvOJ
/96xXfvYHXW1ApgyaWgrY/Rrmmoo3G1Cx2TmQf45I6iit7nVIJIR7QCy33scRHU7/y/f9PgiBznl
hBcOBagkvWor4/X2i4QxpOed0J/agKN8jwftxrucmccS/GMoIzYRyJ/lwDuR1dbTHIy7xnJiJn1f
pIqGfV/a3pGrZc4qf4PErYKhYBKxYdCVVcarfHdEXR1wvsfppj/9PYvpvTi3CZ3Zf3ujmEGDsEfu
sSpGLsASbAPqpXD43CmM0EMLFD0ludEa5G4ypFnYi2aMT5hvIHpsmm2F/jh/5h1raraMOjyx5js0
9YKFSc55x7x+5NgcBEzqklYAO1VSmwVg+CjZG09l0ssqLEUug7j9IyYjWJA34/JmrJ1QnxBCLryu
8Gm1PmyopDvaraAimqpN9F8rcWUMM8EkEe+qgmaTlMQ/33ut9QVvV1WAf7DqjzlWzUnUubQHo/6q
NYrrYKF7KCER7cuv13iZIEd+NOYLQD8iB+LgIpvdgFtkRIYlZW6bo1xMxOl3GCwmJ5Kls0ZCsPzk
cxPPLwvD6hizYUjxIBpwzs62SAzkEdr86wt/rmcxUyZpLhzgv21gqZ/M5sPVe47qcpscs6GlwBWZ
/BN1V8Oyvqg2VJExXaGTszepDfgezIVyd7eGpE0g2TZbIjZw7CzYv9HiCY3nWd3hqfmiJZuWnfPF
1I8m2w8FTSvpbnSOJ1svu4VsUBZyLdXlfa+ImboRPFoiA2NrCTU5FOg79Kw5dIAYE12Me0wFM/Wq
a1+Gih7VtHR3LAUYyE7IzYfawmLRR+G6l9I/qQYKYS9PEUsoEGpfUSGsQF3Q8IQDOrF58Cr5BLi0
cT6OCaZRk6Rh9tyCkwBMtbuqHN2qZecrZXmGQF7H96TI1gnGPT2VLGELmFsAU0iG0QatWSPmPfIX
4v1wSB4RwKvhp75byG3iuXg6nTpbSem8exXXk3vGze7HlcbNFwkE1YkJzfNtq7cINUaFMR5xBWvz
2TrZlkWGsIOi5AEBxnBpf1tJufgs1qS25BbhLcdSQ2D1xux9PYi/7FUGFtmi/wnrkGNnqh8kKFe4
K+WtGSmbS/nMhtf6OWhSeJakKwz5c7o569p6rpaKaL+k6hDhPxRRiCzlx7GawBzHw8+dhyHuH8jx
iAGKXhuBAgc6RTgk6q0/YngLuPhKlYQ2M1hsROnYvThuNVJiFdPm2/zIWMK2c43J9Q6nwZxI7zU/
JqAJ+Nn2VuRZYCs3Ia+k1FKLFXr1Mjvjjrwx6A5y4uY/eW1BH9n8iJs+k5SXYdTnYYsoV81VYy2w
uYYw/WE1LdgLITqg66uPXGgEu/lwVMh+sTSUdaubMZoF+mzmKShQrggmGxoxgcGo8iAg+uDxNvSG
yZOQHMUO13U46iVPeM40oO6Os3CdQ61THsVggDHqLVF0mUHMUiuP5kiJY6dbfGNvgCYyK5OfLCFO
KDon3NruwJTdmTqK+ZglzAI03FNrWC7ert6k94opIVs/DMxyzkfZgoIEUZE5Eh6RV9sV3NIXNbNt
Ypd4H2efWtG5lYNcFmShs8DQT1RVdPjoGxsam6BecJE/CjKKshBaPxkRAyV27bUy8HXXyI+27lAJ
bcxKS2p3Uy0xLmgTL0TotUyt6fRISA5f4XjNw+iej241YxFTEVpx2fljCKUnv4OLajf+zc5ISC1x
v4mwO+7TKKctR7zwU2IWvMOBgD8nZ3eDuGytIHH2ooC61A8C2XFCLWy5r1XjOnp0Fs58ozBNB/MC
5+kLPrt5QOYDo+F4aU/ohGpwi8Z/bl9h7+Cxqq+PCgXN3hmHha4+S0rRNPxRhJ/Cn552LrldOuS/
kXD+W9adBX3BOeZgtuaNZ0qwUQ79WM51tH4Gvk6QHT6s8ZTpJQTfyHRJYowaRkrK68o5mxs4I1tC
932cohXmh51CiZF9cIBLI0Nnu0acqgFwMN4V807OeM+PUZPSTHq6SO83iuR/aY2krUrnSpNQ300v
VeLbccYmfT0tVgJAIuOKVJxep5rJNsX1yZZX+iavQYsCK6+K2zNKESv+5+V7oS1yrqS9HPjqThcP
k4+z7Jg2UrUJLV1EiSJPCezuyITe80qiSwK9NhbyfEYO99a4vGTupOEWi3quBujtyhGl7ru72fo6
hBcLOR05T+n8aFgM1QHbEL5aIDEVH0H8pCPfosyOqBuQ/rEful3yuofoszwGs3lvIBHxHWvf63Ax
lHTohWaFVbpGVuVfLbREjrodGdm9fWhtRiLJyaEZLez3MFM92qQbrrQr6zFp8B0HpBg1VhKKLSiM
10XAlJfbrTDriBHCBaJgDljZc1RHXkrCnE31SlaTzrR7y0uf2iY5HN28WQ2yhdKuEmlbGqK1tmDG
clAGjQbyzeGxngoBnAKyCQf0y+fyOiEX860LprOmwwBKQjndzGrKW+xVCArUP1nq2DJqXgHU0vWM
45i4wHUXsP8LLTZd1Q5mmlihXCQuCLhFncZ42gKPne63Tv91QrA8m7QRf3rd/Fv6NWAD8qsBFIaL
Rz0d8k7dRuHi6Vhh71ORq9YtSslZmelAlEXtbUe1iSpnnfGQYjB2LXTL9HontZiUJSvxobw6mZKn
iGhmrFX98h6LLMcaEUTATpCvbMA+htHhkJ+dJtvRDtD+8/RhaaZcsgCwlM+Cd1duCpXmzB3mhRNE
YGnY5GSwArm1ph9pHf5ux5wXwlXjdyGrEfHfMfC8A3x7WTsU/h7rVB54pBT/qkHSN3N0uGrpPgCA
mCLfv72eQxn/LwGt3JSxCfd23SfZzZByiE2pe7SXBiM6HZ+mdqB0R8p2IJMFsC1LFPLaYuY5vPrH
M6Iyu2Cl53wIdojscehoNONSRnwaHdkV/iQNjKKlbQObb8TNj6/5fzHdTof2TRasyvUUUHWpXhL+
zpIaxLV/51xtvCM1PoFjN47leKFz6S8X1iPFAaL0P6ZioV34CxcNwLx/ITX0L9DMCNxnjMc+Rtk+
voZ+aztSCmOpvGUFlktIWxFLb/v4ydy2vhJ2hK2vTvgTHseiUZ7sxslwADHdpuikUgyuTFkdjAL1
NTSHkXPS+rM3pvxBRasKEGl5PvIOtBVdKdbRyEeIvSTCYfe2h1z//eo3oFDhkh6AV4uIiYIzn8jW
HCFw5Sy5FxvxJ6uZJXW6aZV3UdGbhWWjsAYFnr3uLShFL198eMqSP6uubOnqqgVURagytxbPPDB2
QsWk0MofKJ5oPIScKPyZ99xG/ij0W6CiVxIWgTm5QAsdEgNbXQ2cVSK7C3AN6MLsrLLTJLqp9Nx0
plbnBSuS0K86EzqLuhM86fTo39Fw89CtCEe75r4f0REKxOlQFbQnCAJ8Jq84p/kGXk5jjo7r6m4V
FBl+kTXpojrFd+kPV3SMyaMfvdZ7nrNNiwaB2A7IEJ4HJi6/HQf+efeUTLjx7NpCnFAAMb4VU9eQ
1xI6efj/z2siQOvXbJli0rwxgcJ5Oh0zu+lAzuCYR7t4P+MdrX/MVEl2KfFy4PR71B2GHzETBmLe
QKx5njwJ7AnHwE3R4OZUi3jfWXLGOTuF1EqzO4URz1HGc6mUTQOUHepOYgsAZJei25p9l/WNcHDS
Ey68Lgco9cQWYwIOdg21133Y3/GgrFVpm1gygWLs4mcDvreZx9+rwVrlb2UdSbqFa3ad6j6cWsJM
CYqIjckNzJi1/rlkIFGfr6HYUUluuG8mKlmvv26q8IxB6+r8qqIgSxf55DHhAAoqmR4CQdwzVNUW
hZZdnJbSZNkD8r2Mp33hsRiRsLAXbR5p2xEquoXlmA2HxDIa8ObEx0Rm1s/5ewSPQGXtNycWx5UM
bH96G/nt7q61veffehPuGakxq6X86YF/KS33RSwFKUuCocO2vs+FiEgADPEomLkhBUwLMYHsfRdg
HlCYAebipz/it1zsVGZzEJheYTNG83apXTMf2SNcmtzg5PSIl7NmD92f5D5dzZji/ue2I/KEDcIL
A37T1X24BbWRJYWDTU8st/S07NeZoLcDh9CilOvaaLKM8KT6vUgO6IdTf+ob5dV0ug9o2dmqYHjH
oQetSFs9cJsb/2aX24y/SKXwsyeq5s6lXdZNFGWErEsAfnOpi7rLa0N0YQWIoOrzceWdKTC5sAvE
C0JvRMjKvZPxpecZQt1flCFdLc1BYhW9SwsYP/MjeQo27PmHDk32StLBSjVefsFZTUy4VCTh4BGM
8Ct+bmT+7Lq+l9b6z8CnxPSAa9sE+Ei8gbHfKoqJDekxFdCrYr03wO1KuqojKh30aBqvi8I16Aby
5XMMWKhVIbHuL0x8bw/l44qnqldoKB1qeTVexxC8UrrTf9I7nGt3GuvcPf5rf88MUA3vn0DxHxq4
KkfWhky/YMus0ousQSt/ixhVTdcIv0BlW/Oh0BEM/F7c83kY1xmw+qb327yH5LqoUsb8eCzbWVJf
z3QwWp/BoW5FgjMcHpfWq+3t8OUUbdLrpLomY2yVicYA2Sf8LZPCbDQSnBDv016ADOJtQBM6v/vO
XPX5htAcrHSNiwevGIoRxw8vNNcpIyWs1+r4j5+Q3qBVUFc5ZjtSjtp1WmuMUeWCmuy1mvWfQSMG
37KnsxvcvKxBlq677PeNLBKOlL4QEClWD67JcjD8843JBc/DVcgvpZjByr7x6Jl74NuaP0yc/bjv
nCzIvkCOH2K7ZqVHQLaT9ln9DNQVJVrwylVj0nb4izNplv6nUfmG59WMVjhshbeVguDlQMTcFgs9
gAOkpAc1mEa5AFaJRQU6B21ClBmipMs8hP3sJvzErNlRU/DAIcOnu5PzQ3pquUP0rpLD0tztxM+O
znLQnBe3UEBQzwrUYYLwZivqiMZht9l6u3t8gTFfzDcJfP2e4JhMzbIZI+J4fMF149yC5sz7T7dF
mPbuBb1ayznRuf9JU5ZtIRaATjL/GG/b/U72gBgoJFd+Rtf4F6/AdR7lbbx6W/oBYApg/v7MTnht
wEXZqFqA3xCtBMhFQRWa97jzfqi2x0hgfeadQGACQR7v4z+Yt6iRKXJZUvdeD9DYKaAsIJjkhenB
92DBhT9+dEN4Kl3SqA8j6YSPjAqddDqQT34Qa+N9c0aRHAsadTEBQBvLku2h4q/SBFjGkurZI31k
y2uD/PEAytZu1stxPBQKgJbz/b8o92uoi6yPs7Qprr5gfAogLxBvTv33AsP0Uy34LH0pYEZDkxHp
WXPZ5kwdkmOX5DB/KiB/9tFfxMZ71ClmAHySYMw4lcP5VUztNKHGD5hOiDuF7PLepTzGnFJkSCT7
Mj1YPi4/M2jsXEudqM4jmiiB8zOKJf21E7SE4yE2TAhRTX60D0nTrtI1go+2gzwgEvcdxSTFi1fD
4ezXtxUL5Mp9U/Rtkbjrei9jI9cLKsCmmUob2XO4oNkkBBifK1QoV5hxGXS7nOkfmMaM9OOjIEmy
4OWYOhvZT59wMK0s2SMPrUdgvEMgnU82yYKFlb93err0NlygrujPNK7AKF3dcJd7R8xDqZhRlXvP
agTyjnOoJLCt87l4QE/kFXLfAd835qap/ZktsxiMCi3eKlNkSOKEStkCbTDxjKl1J0on6YGlYAg6
JNb2px4We8chOVN+YaQCHqV1q4lQP254j259+0KT9Q3qj05WR/uvLwmY3aE02I6yVudgkMlWJhLj
lqnTJFpsdhhqaklrWCKuEbAZqN45LQN5ro54Re/b8aYAmPwPk2bIhLv78LuKWsF4LcNQJdpe7b97
isuqG+QefVPHdeiRtjsrNWdqajPWpcZF7BYQB3Io292StY44A4hU0QsuYdxWFy4/DPS32NRUBAyP
VlNQVfCWdlZ7eJY5XyZ67ubgsGpRzuDNDJ5pIMbdPZ/5u1pNbCNqRaI5D5djkgtltXQIlmHnYxa+
rBnqEfjQlroDyvVSYVJxTR2jdVxpBFOyb6IhNQ6/YR5zCwMewCx/Wne0369j1YhGXZTzSzdwUDAt
D2OtFyK3nB3Yy3d380vB1dspVxVkW92f4UVK1GfEgMonwzpxWv4/uZms5wbAA6eMf4nWB4dtuIZc
wleUqZ1w/87WDJAF75TSLvsVNt22dCcXdXjCln6ANOtjceGe7oIC/rlA+Ks/lT4AoCkhDwnOj+mc
SrfukRV3ehtBxQnfeHYVHAsIFTd7f2WPCKZC9OdzpaNGr9WsVU+EtVYdcLjI3+wO5fr8lDduTMWY
z2tU3U52qXVJQsTm+WhD2AYEFSR4AdBEUDzNBHuyPQqyLktGvAuGtkgx5K13RyY6bEDH2NMCnqAV
0EoUZ4l5AxingJCHJC5BqgZU13uYvYeqsNkejCUsyg4f3APg+o6KAofBwvvUIatotpaarO0t0rBx
dhr7t2SMwz3vI5EVuyLFU1WGmVP1GwG2cjfUjKudIjrIrO4aKTKMgW0n6KUSexgXV6X6QV9OyX2S
Q/fFgvgRdMjceF29+Nx3IWmQrlIT89FGvQ9eCk3GXv0jXVwXUD1afVryXFy1axicvnvMItnKlWiw
U5d8/tHVBwznFvE+XJzEeYszqRVAaM79mXXKI2nDe3DpSpU06galyl0i1DWyKL5vwkd41eHMf0Cp
caI4rtzrUIwM3dPqXTrC45gVSkpcEJxCBMKmNcDHRCQVjJ5wgUuZjlqoJEyBoGItBs/5C6Ccwthn
4Q7+jOVjp934pf1wmN2ep1mwcnvBbfX8kapc+m03BEkC9h3/wEN/XAazOWSfLsgwHHR7ztfcQaRB
5JEfOcwkiIe5WlcjNHjuB3u12BbirYBaYq4wbDsLJ6RLwzK1jiZuHiQiYKc98OzbmDZ6Ce4aIGqx
lkJyNhOw3svALT8acT3Dc1eIhNF9EyQVpvSxqT7W7GiWpAxdgL1nSwje4fXfDAvC0tnSb46NHFNK
9BbBDnT6saFHqr5UM1/NC39CG5NaBymaXWJ843arWueX21ARH9iHwHFcqn3pZVuLShxE2CabOgJE
/OMDwtWBHxL0OLWUtLmoAdJCvi1AfPISbhu6J61JMEtsJKwG+/e1BZOLDLhEZg4NDS5yTfTtGhlo
4lotoO/+0HH3v7t3YjrZVvqVzANRcpiWlij/rY0GoaLliUpS9n8AXN7c94yivHJWFuZ0TjseS7FH
BB0GPtA76GZGXCjPUpMLhjLFwqMZVEbuvMxJJkhijJOraj/6fWAySsULRv7e2SwMkpnTTy02ULTV
4g88K37BCFKN/auDSi4/Op90AWEC+o417C6kd5trya9v1Hxoyq1jQs4Qvspbye2eULfZrB5RgXEz
ESpQooB7tFS7tOlCpjFMjG+Nbjg5pnwErI9DmcbWQBQbw+Rvv5NA/ey7/X9VCXgOA69ObwJvuJcr
tGN1SKe869eTbaGS2YtyZIiFMQaW4XbCeYd0g3QDM/vzOz1f5Y7F/hF3EOoiKYx6wZzIGs1F5KxK
FyjPRHIWUDT0YoVP8vgOhfgViSafeZJHQMSCYawqKd8w/R33SqX/ytK7zoR39XJX0wSk2jID9efG
NS5LmiaLO5c5qiPyTv5Glu9ullWvSPtexsMHn5SWorv2FGvS0NgWFSpr2Z5IG4KpfbgnmfeQLLfs
uUcHa+2ZA9Q2rx/U2bFVuAoUHX/vJTwK2KB/P/ISoDcLsXSq7lBvcqwiF0msVA0JvpsbjwAR1/hb
Bzbq3ZqV9psGqwx3uf8zZqor84Cq+KSYHvbbzrayLdSM1Q4fip12O6Rk7oLVpY7as+WQHuPTywNl
jgQQ1b504yg7N8FqQgDv/IpzmXl0yOjC+JpowX081aEF4E2RJYQDIPnyRQmTueSzFiJjC/9gub+Q
miguxK1Nw12LTH/6ixRQ/SU1KJOmxqDnGrju3fdV4xwSnlX7QVJ8u7WECPHVFqHHrO5Ocw42kokZ
8oNafyS4hmLDzcb82dHAHgnRlFXG7tm6etExT+/UZ2cApk9UTeheRnjI7GYDcGQJwTfG/djl81jB
klDjEl3IeKYcyQPbsoEAvtcKzsi3YjGfVn34t4YAcMoJHC+7ITVlSkh3F12Hew68a9ObytL2tlaj
pxMD7KM9O/r4QfhQiDYBHRxd16KUNPULUdzmKh/O5z4tCfroTUtbtT10P5OoVETrU9ZK7xWfsyXa
GFcp4hpRo+Lwr91RTWATGiLTmoT9osRh1+ckEh+EXuK1iS13hxpnVLtzhMM5YU3txSvHpPAixXiK
dYjyXOq1dOeAukmsu8HxBNQzSHAFykfHOFolDbdEAhAW4sB6J2R5g9cVo11OKWcy1p01RyxlmWOC
9HIynCkRcuWlfgkiH0mS8CdD9vZZl7OoXS4fNOJ9Avz/DkUElzvI7W1U0fvjPbCXjsvy99rESEND
dj9l8Ko4vL+ucHja4HswkZfYI0MxXZUD5wBvT5bmgKyUCp1RWaD/au2vLD3yYlAUC3rXVPHm0MXI
zfO5V5DnqAuuVy2+3UbPcUSk18FCi6B5D7qPd3TVWMIsro8vAAsbFU7HFumIikIRPHfkd7kcPYLW
u3J5mqo4iAQ5LNgKPLYo+6vTv9CF5+5pw+OQWVwnTWD+FxNICb88kiPrIdKZzn/DA9+wE9M/9DmD
RuH/Befxfp5XTjufZLSJvtsuHZCr4vDBapjLbZIHwgI+BSXAg0FL/SzwLoRS1k1PW7LtTPLxseLk
3QKgPY2jw6U403SMcYS105pBevhscqhn+e3hvOBFt31DjsJgqr3mhzE4kzYe/KLiVPDQe4yq169S
2B5s0ArPkiiNMfa74whekt2IHWNiKBclQg4STaQXynvjDgyZUWC3BpE8ef+XfsF2Vmzb44FxckmJ
H6UUmVZPI7DSu1w9vvl9LL4fZMAcTM5/wupbOwNsB3ChsoQpNpMFeX9p0zaSOOrnEmvoNKz0EMYP
yb4hCNHAb8AyQs1MLS1cnGlyI493T8Zsnyw8/v+PoWEQMM8sicoTSCLnquOsTymUw4uEgYJMVUf3
RaWaRjSLb7WAu7arOGKz7MzzeK+XS2kQ6dO7JdxPOu1SHJNrzNvFZYIi378g4/ULV737DnsMQKj5
64nHRi545gNplzy6zwm7TrvsM3e429eBURXjqQW0npLGRbR21k996KEQNcE5IKLmBDOZ+pauvaVA
0hB0FeA3SgOjpROVqRPYCYhtAMqZO5FtzWnJB2cCyaO15T9ja+v6Zm3t6qSCf3+kHP0DA7NPl6q6
kWTBf787dd7zTX8BN1ZxrsASHz6+BplvG6L01d8YmZY9Cqiy1Gf/zqH5cBNhMSToqQ00LiZw7pLX
zVaNUDJS7MbUGHawFf4YHhR9WR+S+9RtqdfBFyM9qbKgp+B1PpgRtNktTalHE/gYFo8fPwTudNUJ
AdGe1lprHxxbmDBVILAjU/Nja8CLdw+1HrHn/gnAJJk+lrpKeUN0Gs5bbwA7CRYSZ9dMDn+dpj7O
Tq0G8HeVQ/GQ6n+ZYJBer62ex5iX+Uz9jwz4DMK7g9ClZPG3Mf8B09ADRL/QMkpxMsRLU/35EKs+
RKf2OLIvMZc10xQJDyxu1yGsMOj7C8012Nh35t96Kt+qp3egR1nB+0PMGx2nwIg3zvFE6RdluVcI
hr/E7VXgrXcacQaAIx7RksqXMK8xCFtjrpUvpMMOLlnZRP/9ASMEBgRUrG+IfwIEvK2Ehtz7hMFu
qhJOjzWo3AcT50yNXAedxyqAU5E/APqR/XvF6T/IgoVmtf4iPvZNaI8N35Uf8cqSvh+Ygz9klg4t
oCyzRfqexqa97q7GMS6oaKDtQc8YXSiNCowdY6wA5Ws0o5reI2Nj9mxTfI5C+es7BjqX8zWPtE1D
aVk31sTwnV4QQetX5nARaTts7bMFqLwBmyw9UoBlKanRsaY6HXMODwP1QEDIwbmxaB8i1TUuf3hi
jNS2GUlP38/j+edAan6x2ONNWcZItKdYByAbbLO+x5jthMsil+9HU3I0AIXxEgSItCueXMmLLAZe
q7izbJ79SdPgn6rapL700q5F6yFVnYn8AJEe4xPbLm/lQfu82GehZisAqQOQvimoSGMhBHy3wggo
9I7zWzCiGZOLl05ULvdmPO3SPWOtA8ClNkgEJIt12M2UqMhgpdOiC/74ON+38Zb7pwffKJlKtYC0
roCUlrF0V7qkPeTbmGOcK7S9nh49Fx2ssw8P+mmAe4XJdN/F1aPxcZxHa9B1iLy6S6GRLwN7KPEL
FPxYcEJwTMls7lW/UdMBbMgYOtiamxutEaPOv5ZaOIlm+UXFJPJO9RgIqoV5yzdUoTmVIL4XH9N3
xK5001YKz9tJOWJ4yc68WiWnYNsVJiaDT6SbvCFchosCdKz6eeITp2BdAJT+WYO4PK8oKq/eJ6td
skoBKCZG/XPXcQhoXAg2OxLypUuNyuht2CYs8iA0glt5C5skb3eTw57yx5x8RAMlyuTcGMgv0qrG
HNo/MhHKMpAs0OUhfgmWydOm8B+NV4899+3Sz1qiZOnNXveWbWT2EE/DkFm6rnHrQpDWCtu9XDbZ
tH+gUQwE11p9ovBc4czskRmNIm6S7hc4cj/SH3HGA6Xd+4zf5ZkhAoMrzg4Yd1lRMnwwm3gWVkm2
kJK2nze6Y8qxRoo0uxEjPrYDgowlGVmlsq+xPBCnmVpF/jzWCluQu2Alx+3efpukRl/bGK9pBkwX
ebjlwNNP2Q9zL5ToQ4rL1PgARX3t3DmrJuhffr4ut/X70EyeNbtj3Q42XmimkG+txWfnKN+Z9Hy4
uvIJUCjc8tb0ZX+lwhmlcW5TsDnElG7TX8l7h3uvDGMVPG6oCHVJOLSxvxLhcsdgSo2oN9J4sVfL
ijGd/HC7vlVC2vL0E/4YP8qRcBVGL9Tia9ggVN9ZXMpDdFO+kcedyOZGTuN46kHzqT5i3QNUmFsH
vHnnDeUmz2bhypnvwSJIm7AeEIs/JKtu05mgqqTY+yjZa7m+j+ds511VWcxtBiNaA0vEVZ1sBNDk
4XucJxwMg0QC8JQwPiFlW8CjP795VROYETNDk5HPPdtDnmO8nSUZqhGUwZJTjzH3c3e7NYmlQMg1
pwwelozJW0MoNtRVHuw3xsOy0Rse1HuhR1OmPVu+XbiRhFdg9DVJ1RgiUEZH1w4Vr8ifq079qrk0
yrtbFeEyePnsXeYgskr7iUsTPMTZou37yh5TcoWy6ieonU18nko4bs02O83EYarErC6VaBev3v+g
CRe/0QeSk4tdh0HudbQCeOJ1wio0hcfbK3F5DJl3Lun7BMuOuAFkIBv6dIcBi32t92mX987U9H1h
doxlaqOwr/2wkyXglIMMNp/Ibj8no7tuuc788uFldoTrs/az8FP4j7QlPsHtlorDFaHRPypIMsgN
LSKRpNQ+VQUEUCk9eQUrwT5VcNC2hxgVMBIAh6NGBN9tLAcnOAJTDcKaqzE42v4VC4zqGS5FVkLv
0NEiMIymy3AdK/XHtgSszhSXPou0XoT8wL4qVGVOR7Ha298tAclfzVZgo3eqVbCnGUbAdrVINwcf
ZarR6cd8wZSE4etNr4yHLa/61A2fT5tHbzO4phbnxstET9xorpefv2Smll1y3pB6EkSbYuUzIjmg
uf9DnvD05aFK+yuZCsBoDNKPP6/Z+7am/6onsWcZTBYonRRkj1zZMSvqZ4R5Q+BdyF6DWndKV7Ta
1C3WTJY6pS5jT9i1XakLoTUkUCBi5/X7AjVqOOcOuMIbn3b+IK2cqTyNRtCA2rh4DHdFY4kJYNm7
a6eqRn+Vdwho9adExqqPwdqW2NXWfBHCMSFlSyO+CKXKA/YUn0JVsNsDJTjotPxFoa8lfgza6lDq
Hn/UW7E8qtV+Mf7uz0noG+4YR7emaLfmieIQ8V/ou3S0E+/5ubLcyRO056Dvv+e9FpFWJEjwsTm+
P81i1UIrpxqVbb5LEBtRKffZWaQr0dGQ+iIemUXPiu58WDhmrenHZnIsdfq/DHvKQNhDdBu7wHRd
5fwWgPKkfkrorV0fouE8aRZNhyz+o5LGn4nFcpBYrCkaF1PjwMrvvNQG15dkoslZzWJVadpt2cdi
nYj3Lki3ttB2M+71xw64P3TXm/wh5yzkyQyGdXU/98babeWoYNAcZyJz8jbcDikw0y2DqQmISfNO
u9m/E89MjfFZ5tiNifSwQlp2Ce2CQHxH44C61gStUTfmfI2DHRCOHrxCUClMhGld/Z1JRVrhShMS
JflVbpevNSWF7WoxEfL6aoU2de4Z3ekVZ81bA+s8Cd78lktFohS6nFq5WPwYC74PZWx1kmcpcdyS
iK+3HY9g4++r3mqUtXGbHOaN/t/L2NKNuI1mhR5+ngKU19F8ZDLOaX/Vj60M4jUElyO1QhJLCzvK
I8S3nGmQZpIKv/8Xq+NydEbcJN/h5vlwMFeCB6RRZ0hsolho+vVAvTKiBec2pLMc42oR0vI0lPil
FCjYC42IQae1ytxewcukLye3d9669hfSKUWjwVsFRe/NSooQrmnHbF3CX3qxRu3T6sDZYW/Hx1n7
j+PQ0dXN49blZNzUi9AXxhorZUla8wdw/DgxLmroHV8W/heXwv/6LXEPLh23HzFoVa589RCwCDNz
KzlcWJEH5ijkk2aVPsCoMXbo7R7JNXZuTYbK91lXMsZlSVO2KRyK5rK1J9CgJS1W9vUiqpw9CMIM
G4k9nqCY9MCttY7+zkCC2iQDf2v7dxmw8ZFLlB9MsSFoZHJJQ87CNutpDKZl7ceFBKLtO2vsbQ9T
4RcSdkFF2wuqwxXTHBg2M75vSS39tT9nB4bNB4QC0WRpnP98p0JENgxMV8KNtaUFSMgkJF9MouC3
4+veDGO5uETHJa90O086rUKMV5miT3l0/1Erv0mxXssTDJO3rSEkvhsRXHCohs3GDeX3MIq/QGVC
Q3MH+IV7G/cwg1nbUk4ce2KiW9jbe/wduHrVd2EaiHTEB/JhE9Zca2Hb5O5mGA9ASx+SPp2V8+ia
QJiIPuMVHlPYA0i2a+oz7uo3HYSNDuLW/N/stWVmglJNTlata2Kk2w/pp8U/R9XCw4e1OlGkO7hK
5cT1l4GyVMutl5UVeCxEONIVkIJyoWkDHOHytCkaaNrY8DXDS64vk/zPrmiFMm/gdmJu1QHjaeeQ
KHrI2Q+gy40b+CZX43+qt7DG1mCxys1eB9u1WJHXGnXwlSzTJWlbDXy1spF5hgoX66yZV3wlVQnn
GLPYQ1bOsvuNBQf7bVxmbBBjP/QgfSsDoJ+e+6jLbccVdzC1/u91yXCP0xdYohTFECPB1nHgp3rU
VZ+Y7l8G/KdzR+jL+OiMr/jJftNASHTa+YgoOycvfVgWWroTGQ/vsqNOXlm3Gc/ioxs0SKAzfNHv
Sa/qqs5bjhrLcaJFDd6aNhy6J6IT8Ay+e7FA1D/8wT9S3QG+aPRPIRhDusIWtdPYiYWWgJf2XYQA
l8v0LJ5Prvg68p6STjC/pgHeF6N3RkTUCFuOvV7EoPHEFYwCwf9TJw3qZB+Jp86MWKdA8nNu2fY/
zUCvgW7ISHVOZ83tvhh6+X237nkOPu6Rn2XWxOHvYF5V/nldlOW0AOL0iv3ySmmyJRi776bEPRsv
c02oa2rmRhNXzpNGStdJ7Qnt6olxci+QPVbauzRVboyJqLFa6FYomWtvxj9HzfWSia6j7GDZKKzo
jXLMwo4BU1ghxLFMd/B9cOuGuYNPoRtD7Fv+yRL9JrSOdA2VjPjIvQyg8EK/rKDy5+IrpJPEO9bS
HvEDYs8jB4LRzm95N4ak7vE+Zj1OajXFgH8R+050tGtXcgbDQbr4fswM3/4s9yjpA26JfcRxTBGP
Xwe/iXL/Vyav84emDqjd5gQogpQCYpmdphTvp4FhGI+NSRK5oBTqnYAjZyXms4En1dbCDymETOvq
ZwRSdhcO9ol5BwaBPU03HENkOnnPz7+IC6yGhVGvBGMAq/2LFTSvJyonJa3EsUpVhEFIXqxoM3IZ
jMejcFWS66Xqu/4rd+Hlf/+t4wa14IN0zQLD4fU0265/4N8p9M78HsV8nPQZafJ+zy5S6JK2gKDb
DnXYaFNPx4gxjoF5h7r5PA+DV0DVujYLCQTAy4+DIjqmZ6mVLZXSC8a6EXP+uQAxUK/ry04X6wkX
yqB7bXW1jW9pD1gmmsVyJd9m5mya1pyKyTq0oATaGkg0SBrrlSjWYsNP/ByyiKhyLU5b0bddYBGE
1XPegr9L1lVnBUOA4HasdTe2oa2Xr+4wGDctEhsIP0YtqB1PrVCytv2CBxLWxlpdecFNKwmRpgNx
I9i44atX6BNeJRKeguPXI5xIlcH1Dy9HpCHBMraFsnwXRk/E1V8eUysa/RJYN0fgBlh/LPRS+b6D
OKQZ72XvEqjsH1qGL6lsDSF9w8ktYA2loQRVJKm+T7DLrX919adcDHSEHDzD4iivbQrOTf1bw0Jg
bhzxe7cQf+3GemOjyRYaQxyh7cBdyEdPrxGtbBzwtizguMh8rV/tJEVeHyX2tiKwFdaEQLQcbswn
3Dm0vgovQMTg/P4y237/cccM1OjdbI4UXB/6NYR2Dxvcopp1W6LuYBidrrWwHALFos+3eM7fNCU3
/y1aLXMbS+C0mk2GOMH/Wlii5QQvURhWEiwuacTTYEL6d4LSlj9IjJkCb8O00npeU81zn6UXdCr/
Qp8XvwvM1R8EsIBSVU3fpWZuSAO7xq15APsoCjrH3O+TyQ9dCRgDwvNfMtczpSvAwv82mwi+zwZA
DiyvymARBoOYOoXfbf9dBIEZLfIhlNu+942THlQ4xSaHBP56Hkyj+AngZPeizpny7x2r4cBEqT0I
gCBpF0HR9boGVSpEnA0UzsqSkCqhYBTOnHT0W+H1wjOCgCpOfwLWqm8K42Zr2ZcnAqOzAe9J/90D
B1RhGoxP8b+A4sGaOsCqHXkH/bgJ0jq4iYXcsElhQRtPQrGWIimkEPIR5JSqtGdLsaOxiYuVnFgM
RF7/MfOcYHn/Nr42vJk56lQDQPJCbR4UUYoVWHj+oy5eMQL95EyQL8ogOfY+AA3p0/8l3AOt9zNn
NDWHJWJtHD+IQzp3z7z7EjEUNTt2nUvazCelvvHa1nUP0fyvQ6lPk9vpnqW2OcgnnQYPQVNPmztk
cYyR18+2nCjG+cve7wlTcq1zEcaSWMn1OUq2XTIqhz8hElhNTEYKY5jO/Dd1DuTIQR1T9tynKr/2
wnj+ltMehJyeYb3nsrI3g2II/w/yS6hmuPpahL6av2+lUBvefUEcft6sw4IiCLwseGA1iqE57V6F
bboDCvOVZhnHam0uN4/qZH6oBSLhBOj/b+tM3u36SieqchELXiTv3KQsJQ/L7EPyQF1ASZ47iEVh
oi3ayK4glizaZAl3e/vy8tbp+LfLBazAj6ysDrvsv4Sq2QVIRMMnOi34J1A12ZvMb4DVs5yTBw8n
JAwvaWpIrKdbBv+5MB8p3wHVG/a4bxsaFUzctSXMoyBcF8YqR7A6TbMPLWin4DAIOuOu7Q9M69zr
/IRtTTEE/KJH9iJxcD6dR6KORgSayxtvVWNkyYlSIp0JUKyYQ3idwoIPQ1YSOvytSV48djmdYHzq
nR9PB5MH1DsET+l4Y1YWfqxQGxR5n0zECAerX766AS9evOC3Dsyzi1uC/iQ9paz4CJOm1bHVn8Vq
wpzy5tTbrVHiyoNEPUepv6maO3AETvYC3d53uxx3ZDSJSvCLnkzhH7bGyzSeIg5W740+w5lrXXr/
KN79k/pZUS32B4xm/UxoVbFSxEZKWGqsgv3bFlUwqgyMb034EQb+VSQpJVOSZ5qXELS1hrL0aiYP
FZfLGEqBF8hV7yyi2WzQBH5NYpTsJ769uZWbOL6Pj2uk/67/kOwsIBw2vFwHFvcigK8iqSFtxToo
z3j5Z+QJsOa0OH20WoZDYg4OpuEhT6WfFIC6PS2zunyzoHPqn7NSbUxNzB4e1XClCoJWDkql0I24
FZR0FKSqwYP5KbL01KeSNeauva79KqhxoglfUHKxFuWnZILex2aEcGCB5cB9a6TqbDJE1H/sxyB8
kzXjTm92RCSqBhe1xjyWBPCbrL/RADfZ/B42mO5Fp7ZkMED1uW6Hl9wIijfCd8RiRoiiVSW+CE35
RL+/ogQ9995ftyivNcMZPOOrPIGh0s41PLHJvYlG6PRX2DVRl3pHZOTdWjZWqaG4nY/9JVRBpr3f
aipLY5kp3zDvrmMudCggkRGx+goSyZccf1Idb1FlzcM4BQ+z/wndJC0h7yoRfFOh1QJ6lilcBvNq
SCc7KSOM5gQbozkO4IkO+HHCBbuKn047yLy6Bm2OMnxWqOj7n9Y+Z+GyMC7yj6nKVGhhZGurzBCj
zC5MF2SpUh2jwdgrvPBrFhZkSlfLrIiQMYMgZ5sGLwx1vGjYddeKkPdVOxg4O3VWJ1XA2GV7KbCG
LZuO5H5YMw5IojAmdXsEebtyiZUdtslYA8HvBOhgnY5kkA2tvWmpFQt1V82s2Ni6JRladG/2H0h0
TL2o7b+BnEiENQ1zo8UJ0RLMRhdbza8/QcuxNf24WyTaY9jAzWx1V/I4OKpeWnEpO4BcIxEPKNmz
p7sthPV4gXquL+4cBo72pI4g982VyHJJ/0En4MdLMOSz0iS1TezUsgTH4xx3/K13cX/hB8fS690c
t5BNCSdonDO2+MKBCsAsOwbV65ISnvBKb3C3wVSBqX9FBGoYCdJ3pYbPf0pm7eN9a5F4a6NYiGN/
JetNe1UxSI+QZLSRve5kVjYoHX0BCviM+jH0vg6Kucmgs0KK6n48aGTJeimz/a27gbNdE1PmWUOR
sZpeTxoZYW0cM3DxiZ4fmTXBANIXUrE+xP506GRTWN0PGsvtnInX/vfegzt0b7LB+hKOUPN6DIDE
bnTv5l840lJDtVPopcAG93axOOfitoInDTRxlLPhZ5TyZ6YqqmbpPRxvJvmwTATAbhcmdOE3Aqv/
k3XYYz0h12QlO9nq9yXgGiYYzHFdafh0nkhsIUUqTHmlhRbjd8R+lL+GO/lJ+cgGNlntKd+DluUQ
3V46WKo7oUkvo7h/9WfTX6F9e8epLLII5b6a7PVUp56ydPSHrU83sz9JR7kb38FdEkDuyyP37jAH
pIj9iVOEZjplUZ+/X0AYKHAgLUst/Yt7MApDnt0vKIbV5Odfnme1AjgN38yj+JCeD7FE/80oNX2N
be4qNz9LKILWhI3O5BO0kwV41BOEGvHgij1qtTj7gGtnNSPnco3OZl0jpfPsCgSNEStuf6hO9z17
LFfVpkpUa8ooHN0DJo6IJWrEhtQdgBvPcpM4/rrx9jxonk/1gEZoJCsYsZjfJZl2prMD/d/a3bem
73hhn5k6vaYhozGNXqIJPGJfIPhcmNzg34Dlvk8i94JkMB6ygFZMUH+mziKE9m+6SzL8OR2GkUy7
r/GWURfNA8dviu/UPRyUa91sJjeeQoYBnLaxMmcl9SGkoLMxOk3GQT2gdJkSUajYllqZEU7dIwm1
ThVAgvKmtu4SruBkt0G9EgSCmrqunXTfAJwXwIPqaillfqefU7rRO0I/vftHrgxtllZFYJKOcQeQ
Yzf6Q5YMA5RFkhmmPNx77jSUe7LRLQoVhZDZU0e7sARGg8pdUiw+InB8i8o9oZL8h2QTMyaLgrM0
QnSy5/X1Fr5PoYYkhdMuTDK33lo7LiPnTUgzFiH4QoV27xPSZFs/caF2Tb15YnWJZF052A4pbFFE
6Zgu0436F96AtrDMlGIk/2crsEEm+twwy6O8PkYqwOw9tS219Ry7lKV1YsisTTUN30+lo7SJ3tuP
mXNveYzj+jdRrRXhLUtbyYGUFeW3llMTtG0LBz/BKJANaZPEZbucYh0AE8GiY98zaShpBt/5jgle
bTbCoPbg3+Rs/ZNtvmw8UQWZf+cZgyod8+9aqCGx564v3/ohIeKAP5ZGYQDUinId3OqCO2c4WVxf
i1xW074Zq7lcbCxdW+7CEh5gGTIf5d7Lq1k8S7aIXiIyynoQ5FpzDqsuxd613lwNaFo26VfLHZTV
jl+TpnMCMHyZZ+SzkoE3zAoCjGk9LvqUWVD7POPQAfyFPHdr2U0YpyvHXGo/6xC51rIojdNzHptW
Ae6Y5/U5juYHY9ZLZBZBG6DU4pQEf2xYZA/nEqogGLMZXz61nxY1tdsnbE3EEazATSu7l2fTuUda
bjJf2XtPaulA4VSO31l2hAegaStV/hZzdP3qzlGpRD1eNKWvplGQImBPb1fchmWeLbkOWL1labfx
SpzPXBXnNEIdtlVVwirWp6g0Zd2gRMr+NRCYWg9DF70rHaTN7Zj6BtUdest4wQi6shmIMhDjOof0
8cYxkbacfOChOVXEoQmLYG5QBqxugqESdUS81Alov2WrFnLc5K3zVDTJWfv/0Lml8sseTwC/r0QU
wDDbvfS45gY12bdzvC1NbbJQmBTF1Ok6M0CLpd6EqaI/moDAZqDFnwaAr+R07xQqR7zMi2rGyRCP
enzFYZIf7NtsvuRRNoZ43rQl7rCVAEriANdTN0dpc7hsbTKfWw6FoQqlu+oUa27PX84jNS8u8OJe
OrLBbakOHNPtmQW5RQZZMggG8zSZCdIZ0zJP7424o1RuhWnAbkoKqv5NsZKwPvVX/GJDkwvAq8Gs
DCbXOkrI4HRtpNQhEt08DZkbZPlEw1zCpFfySJGLy0hJqgvllpA1zmhE9o6eysyinDX35vA3xVc7
PKo804yrAT08zS4QifJeHV4DRKLJm8/wk4hSG9Xmwv1nsVdWnwztMIHUMQKfl7aDo3RPDqJhLgE2
ebnQdzYfJW7I1uA3otWR5W3WokbVnuq+96qrwDQHXzivHMdibzGIUwhCK95OzRkkiRTeHqLdulFl
vPHPqliIPr5e4jh4DLLPE3m/nPVNj2f6yxvK8KaOsN4f1BQsGPZjI2mlpJdn+xPhqd8ovi2Jyod9
PZkd4SfLRur2JSypxEE+hIZcolYBECmBvY13kuCCB2J8FvQ3btk8hOoPHObiMNiba2MyIJGjNZ/L
fHc5YD7jDWZw5tS0+Hy7vin7fIKibiQeD1Ymdq+13yNFEIkxc8GyF5KgDqP8CAOY+3C/iH5ChJHs
9dUyHJHpP+y013FlMVxCuZhOixtPLzhbmHc5hbrE17HgX32guWjo2w+ed9v7/h/18Fs9lfsPuc8/
ZheUhEN35U//Ia/f3h39Xf/pXKYSLr9S1kJC8a9vCeF0mcNy8sBZ9HwHxMFWNHc58VqBZHWPpsO3
58O84cc0al2Fdsg2wMsV8jFHYXOoOKy7fALeoDB49znCgZ8lvxNllGyfZlLmbHAf5ExxT9vfv2N1
l+Bph2eALPXWoFtANreWsFS0QyI1RnsY6XfdZaepglohV+8qZ4OW/0kBCKUdcoiwjFL5C8l0Ukig
BfzV7ZMOOEfVPnUpZbxHwQ6B8HvJUFSl8sHHvH/ZlfeXj9pu8nCgn7tfwnDRPBYiPJEbw54G5Dse
aZeHqdUPSPsQCb6Ibv1wnP5kMMZqESv9VI1seF0K6qkRg8fbEB4AW/YRMo6/A3tfUDrpe+OYatou
b5f/mGS34znLRTfFDErw0h4kWG+f3T+hYRgsMRe174pRM2t5PVCVmgeuqCWHUlHtbrrYLRBN9yln
mTp2mgu+5t+52iUpt0jLEwDje0vRUYWFx8Z3XbUwkHRUwlAjhjkeQYAHjjOxjICJprL+V2K63VwB
gaEc5CgTNa2jtGAQO+LMjrvZGpoJUzjl8i/G+J2ReGYvMnUZDVN3wt0wRFrwhweE8oJaHhsp21kd
YUuliWKsdOHJZeD3/pF3meShcShgBB3jIIg/FRV/8HqENwIWl6rvwcfqW7uzgfHvFrGVto3PsOeO
Qvq5ZOMK/jOqGjD0jCILXLcd3HxdvQQ8ELJWPvthik9Bmsyy6LFPotBxrEttpdumCWVBl+tEtT/i
y83hx1C0IvOsrc5UXKaX5KRBrwuqsvAolZ1q1Hisa3/BcnGYrFbvrpq0H/wNNT0CL6o03mf2WAnW
SgfB0qkkTuRd5+An1S95PXNsWI4NtMVEHBaMRrciSE4G8tkRU0T+w7JZCEI0TiH/of9XIFO5rqP4
NvQ6RPulXXhr0A4XC7GY4RS8pkUmUYijTFKxwvZCse6cr3/YQLBwTi2shCsd1uI1yNGwkTEJpl/s
/vbOsCsEi8GI7xD8++pIqmNCJyGilijm/cI4be1Ke/v9B/hdUW1J721/s5Alo0gNrMhhU9VezdYH
ZuSHjNd03yWBNO8O5h983yNvc4qDSlsGSqKbYNvRsfqW4JjoDZm3KSNVJa5e6IYPGVdjNp1Eu/kC
dcG3hlBZcYGjOx3fjD1l1cYoxL+4UASb1z1a6yS8IC6JbB6fDRMCo8BIFtO16GAeFn4/ATliKecO
3IGkBn0Mx0FkMYVzN9tswZlY4H6o1LpvTeDhdhlj7XLUGIHvhcth1vw9uUTFN1OMY8I4rgKroqmo
K+7dM/ASLy+mfiFzv5mkGd4OusOnBPCuA8l8hMC7MW9WlWPkuVPOtg66/m2SPWFPaMy6bmF8O97D
1Gir3ERusNY8MFTGAQ+yZvdp4wkZ/cRoFcJK7mKuQ3MLp0AS7i4Hv/4IQjX6ybLtAQEVVGmEhaYn
A41fB0GAt9W1wbSm+bj6PRAYLBbj+pgCIwibMha7jkOBxJgaWP0EaOr8GAi6hbn4G2d0YPg4WJnq
SKApf05vT5EoLXs11FyWJktxtgoyY4d3nXfgUx8L2OchQ2/mhx72i2oFMfp9ltYW9J9rVbhwvzx/
YypT3oo72IIKmL2E1ce8wNQeCCC495bQW7nmn8NXfiMU5YeoRR0Sh7NGAsbsTNze9QVO5MSzjJtQ
jiT06zn9Hp3wwX3Jsmux9gxuW4iUNKmcVbd3rvLkHy9UvBtExFusVxYTPga/knNdh739GavIVMgo
VhaxRbUKUOU8NVwomnN9CfT8zcIfuplHo7Wf35Yuqt41ikZMGZAqWDsp+uYKtQZV+qu+k9pXDkX8
qnWjFc5MIQEGmMcRbG+U47jgoIiwW/MxEaiUk9uPDE/5Udvh2FiypErjnpRrySXQWZ63h27oC4WR
9T85Bca1uUVI569WSGUYogpJS57iy7VjJADUSkAvxTUfZvj3N+/h2qkldnbVeXmuAXu7DesijNvw
ymHhuQXMiYf2IT8oIAg7MmJAMT7zjIXpA49JnBxxYjMRRXARezIK3HUUjXZsTPKMtrgCL2+S2rTU
8dM8vyfqYvEnnFH0UjsJe6ii6LZ/fpyEWTcKA3llSOFAZtMtKK9Q9bIkxrBrfigVj46Lxz8b50ij
cet8lu1Xir++YjWO7iY76BnVXKBJCq/82iVikLTrQAUBt+6kB1vT6O/IK+U5EiSM5HfhQXcXP1aF
DVZAh2nQoWpyw7tyf66/E7o3UfdgLhiCeOKdaH4jLQHKBijjOjbAyWS/gWrUKt4Wn3kDHYofhSxy
HeHwcFIrXgxJWQFsKfvFFeM2EEPf9Ts2u/B96H/v+eUxYLEgmpxewmiCgwwAObxKC7NBWry9ry1L
Al62twI5jXaWJtgujVKL/0kiI/NxOvHPUVAQg7yeCiFSAwwJZ5YiS4DFG8cC61R++3z/j3AmHHeE
cg5bJAZN4vF0bS9yrNm3AtMzmTfF6Xd6Qwi9B3KQqKrODa7yATPvS8LhyTnDRvcWVSYUY42ratl7
FjDSrYzuXSWAzRPrUTm4OBnMrdKEh5rAN3KMHfsw8bt2KNB/1CBEeizUqP9kb7hIGGSDbj/AwY7C
+vX1CqnF0+Hgv/zgSRnGargtL4XJVHOdjKO6H5cBqWWz4za/OPGyQlTnLaEzYjU7QfHRY5sf2w+V
9ZfBKCENxzwGzCoYHlCXHqns7BXvLcwYxhBKu3CLEBIf6r3eTo8xir2cQ0b4Z9Rc+g3MXDrjkHk7
mrM+lMrrlr3K/3D2LD3ySzcf6zK2c1ATQ+N71MQ5HbSJlQJfEUvo6HNkvRPacJkQY4NZKLL8Nv+p
26E1IqtFd1wiwll49ZeZ1KVFvhXCI8Woh5oL8dPdptFcsF2NOOZNIuRaLEiKr+iryc7smtE4v2Te
07iKjGrfCIzXaJVSGn5612fiI1erbL+uZqXwYxnoFYzx9bI0Ts2YiOrEkQfDHtmFcGiRtCFBkTpg
LpoNVJ2OFGRyhTosgMLiYNz4Sf1DE7qsx9R5ANgSlYtAkbBiWiyjDZo0mEpF8TMwPcJ26wSmsQfx
02YeR5at+rh/bkmgbwQbKNfITK8PpdmsaBR5D27X+hJxl+x1bmk6JkebdZezZWxdAPq85f1exhwb
0A+skWvVDJJVUa84R2/dv2QVc1QoUQaRKf52carPsWQejV9QL8ZGJgH1+GADkW9rveC+KC51xpLe
MXQrJTlfmiqcVjXcDzD2iyXLBUv6X5VSekIaeu9T0XqkgaMBqWjkIjO+jddJMD7k46U94NneDjT0
mWGVM498uuUo6jg4cfNy8MBIW7YH1c60m/MQNm2lUE759Mi9vF2iM7J9r//OYJKhqnXjUuFPpxS4
HXkvjuJy8X9dxYRd27vNXLRPw49ByUovazlK7mR8hWWoDGxNvK/io1Gh/8NXeWawbSmQQ+mswTrc
0PbdijwCGpch47uVIeW7sgLuDfXnXwhs1fb9o6sjN2l/ibApWJM3Ewmf2BI7TUse+yX+FdWCbNum
088edCzfZjSKmC7MEiObFQVQ6l8M8e7G4QhdKjGO5OP+j7Ci2QxnewdOJmEs+DjCquAO4ttGGPEv
idL4WwmlDDnM5iHuXSpjs6XhYb6HbojXMhSujNg7zGejfr5Ms4n0Sb2+deYCnWKTL77trZU0U7q4
/1Ehtsh+sQyXcslMbw7DrOlyceqw87vSEGV0ZQVpmzC9v/irZXpXio2HdXR4Bw+WyyrMdBjU8KBA
08tfp1KC3f4wv57Wnu7Nj6aPEjMXTDT8OVRBlg5ui4TOSycgMJv4dScwjWlZXDahG7cri6eQXvKe
AWMy+Axtu5r22htNNaTw7eje3F7YThDhdKuBJvpVjD0751yY0eB6GYZw8vtkTHldY9V368x/smGK
oLW7FqxeyRVp9ocBlSZR4wJXzzDdGB4U8t3xNtrjyxuFj2uISuMHGirB06sx5KHVeOnp70nH0V5U
sPTh2suKpBtrdg+LDxl7bz2O8UeQ8WMTfMhUWCS4MXKeRXkpo8HNY9PNox9Zn8/QLSzsmLlBqZVM
FIJmM8B1MKYrBve1PRstj6KE0uSIQysPG2kofgEnvAI2FCFidGn+Gacj6tCdfTl+5b6GVa5kwizl
ijPwuQLPJSiLXdIhMVeMyiMJ7C0nORm4Tnir7H01XSkEWibhxkLOj0QzVd17CT/Z7jZ5jZ+gq+v6
mMj4wLHypmPH4nq5v8xw3tEAO7LSeqnokIO6DFpewORBlihSCNcVpYS59ssd1pVqN/GroDFQmXcY
v4b9SxqrGhT0NALWpDazK0aEPOTdlPLLZkqAmFKyAaEyEZU6WFeD0klku8oRy/N8aTe/AWnAKFe4
xyAFpiH1/tFljjPyqfZaszZg4h5MUS/twvKs0xW+IkpUrbrP2Te3E7KhTSr5zhxdBhfVHwf24WGb
hRz22xAVw3un01KH0jgs976hJ2OfEGN01DAw9QEmA7x6pbC3jfKNv+irwlrh0H9ZDPFIiZLVjN2c
1SHTEFeyYZ7k7HA2S0Q6xhTTOiNaDihjKj7lCgsOFGZUBeykmWDWBhDlR/iNx0Nwia7GqS5mG3Lv
OjF6EkZKJXnnZOLcLTuZOKn7Wrh14aA+tDd9pabml3lZXgtKd12mMfRTpDJAfOiUae/i71u+G7ys
3jCCflJOFb4GUI7Ls8pOWg8A9Gj4Hgw4tM5iFd5IbbhlU9SsLn48mekNv7FQy9yCVBw0aCirhVI9
0FNvxH/xiYNz4pg6cNlTxChpqhH/Z9z2EvRHonpXF1UqMthNvwDygWRuewI/phUTz0Nflm/fwF0u
0zg2FzliTRWPTZrAYqRtZ3RRTXCZ+sSrql69E9YaLhc7q3inBH1cicNn0XSXb6OVHlsZtO2iL7oR
qAWGynRtA9/V2FzY1CclzfQ3McuT7XIzSLSiBw/0r6o/q0lxexDYWCpUaM3hQoydCuSoCczEDcqU
w8/1q2j1tXSKniXQLWqp/8rLNk1XjgJnVzGcAvG4VbPMUhPN3XqLU0U4kpgnaNrQoRR5YFArMRem
vTnWK1j6pfBTj3Qgze1dpBeEhhVDqFHvVyv4b9dCduvHX4ZRCIJS55VSEBQ6/+AG+bcr9lnBwHCX
CjxiYDFYlfbNVGR4Q1ytSGDBhDXO87fqbuc4CiIwuIXC1+jGDnFiD+gP+km9td2PXJRpb3Cy/Xq6
vIWB1SJ8+brN4iRpPWeHEpjlliGz8yJst4+4tQ5eIEVxn6vlqVrGPynVoT5OVdfhwl3/pU/NocMO
XMHDzOsMDmoLmioAAasyn6Q77nU1vmPODble8BSobFuEgo4G/TdQHZegV8QXWEHzmr5L6ajxUQ/A
79HrZFCPQMl2EbGGP2UCukUergcn4rEr+Wo5O9a6xA9I3oTiCYZGIEhJFP2/V9PdNUGpeXIrp9By
0VYXYURc/6BxLRF5P2E51jc48iwNCg9tNHoqKUVVovGdCTxsgJHqH9xEeLNzqeYMY+6xyLY6qQQ2
+N4tomZ2aKz+9VA0Gcv7KIu0SFo1YsWafldh8qrf2zVPKyLrfQRjpvHd3ooH+9olM9pdGyfVKL2U
0sskairCG5sE3LzWBdeqWN+Qru8qS1MZLW8cuqYHvSFCUhaKDH8pFbWKPTk/S/wHviPhQ8hRzqFR
xn1kqfFLLFaUwaTBZZL+t2d4TmRFcwdGkNwdB//5Ygsdr9/2qVRxqw0jn5LEGj16/LtY0zgYg8LC
p1cUAZQk8CLoaTj9IIMhPNBy/IrGNiO7T/g46HzHb60AE0iA6E3cG8/mAHLH5vJfs1I8iBsAVpKy
LewDfpdWH3FAMznndjS+KMJuMMAuDXsdaxhSfQOr5OSLUA4Ke3+ZwEYDzE3aesOizOiaX+53kVfl
CGfReCm4YBfEvSi5Bd8Wih9en+hZktBwZH5gCBSYRYtpP9WfMwOi4KgFeqJml3CHd2LAVXlXCYFx
vzKhOYr8mGL41yB50UyDecblI5k6F+bJrqpegwEv7+Udj5BG/HS6LGp4pVgZvUR3h12D9AciofYg
POqXA5bJ7bz0p2DGNTwZRjf5dwHZQAq9Yz8luU2oliaoV5OrrhUdXOb2lVI9t4aaTh2vmxfbu8tj
QHR6Lr1x6iIWNIHr7MRAwO8yFTwFhywCdfcDhWUsrSxKN7XvL4dERdmQ25EEMgRzerNijQHd91KD
Aef49gErulkceXk2nMxKA67dmfkHw874wwCSzSNe/eHuaDo8wIjffDn8qh4fChMSb3ijm7wsUfrh
RNe8muSH76N4ZbZUO/0OAp1ma5VaP6md3YZXGi67oQRmW0QO82ywaWBaIMu7409KjeKQKN4Od5kE
KImCQeVPW5hnjAStTUdNNuRgEDLUM/vbHZZmDGkfOl2rqbrkW5TiOkbz7FK9ludq3oiek8IAs3vN
J9bv69Q/zFspSeqgvPTLLbpuMsnvnHKsmjVj7DikebLs7JSIazxZ1V1DmWYLfeiu1LZMJkQqNuZ0
/ABkyU5aWIqUAimjVO1VIV/mCuXCjA/vrOxqVN+r64GFmYF6veWuMOdV9jhTKEPgkExc4MmQf74D
BztgJwJdXizVMg15u7OtjDTn33LAAVLU1n2voXCmuEGQrjM4zDmE5ewOExA03HtE90AqEGTexnEM
vjAM5JPeoJoom3s3aVDWaLGRHOUQcwo9ZCLPobKyiIl8xuOJ1mT3P9XQDKTzRZYk/+3zhH4YOPk3
HW3cCcRHp3/7m3ev1LGBJmZM1+V2QVjF7BKPCwEjT+4rn+yVzwtSdRR3XuxrEHfy3N2JuVgPzVX+
KyEU0vowPTVFhPcsi9QZiu7hLZy9SdPTkom+VxvdH9noiysEXpuFlnHcPBDgk+LBIpQlaA/2Igod
bUWsuV+aNG8Rhxg9CT8PWpWjg8aRWcXxaxM0bp7S35TMz269eTFTFN1mQzRwmR6bl8qzsnoF8nCk
Ld99GujShRVIDBhgxi9WNYniJ1JET/OPvPULg0EyC6GP/rwJAPq030bHpZgTDgHdh/aUJl6RYhUf
T8is56D2/FuIbdBfnKEiiVxfP3ABzM34G8zR2XVBtlYYWPl1UZalpKNasKjujBF/efvKhCbBi+zY
BeuOFeKOqygb0s4viKWnpDz6owBqLBikxTbiaymHTBK023zUXj/6dyX+D5bY4lb0Jl0vi4Mgluep
BQC9BEvq8Y169Tao5HTYilJ1eEIDc/h3nSivyY0SCfhD/dTYjWxkOjCRVj0huBgqBXqJ46QATk3a
FpkPHwmnyLn16+ny5baN5zeczBNVttlSN/AxKjHAkmc34apbYRv0fT0k6vLwvXb/m5jpXJ+Sd7K2
REzRHWSusWdc5Nh8UZZlT2rcvMEccj0nYpedHEsJVhsY1SK/IftpCCPyB1l6M2Rgh67xqcXk2lwR
8aPrALD4E9ABmWAFOQ04jz6eGa3Qs7DbfNe2UiHkG0NBHo4xHqcQSIw6pPwRUI7mOSTKkWBiwptw
wMl45gNvT0qSNVikZNddSBBINQtyuquqVOSNHxonHCUAXY0XLpWYSgQQHvzcXk+zHxXOPVERsZs1
iZK56g6JhW1TZZfupTB8LneP/cCVZtdL+t2bYTFSoLEUrzf3qmuNSGsFPDJhjvWAX1+QU0E4K7D7
wD7xFZUw0tZAtsSxe9pdNXl+YmK78PJAKfLSgijwKiMyRxrY2EOCkxUvcYJ7V/y4O5qNJq+2qjDK
eYfy/2UHJSu7fHJkkNh+AkXtaheR/SMkKBou8LeSwP9w+BL/mpjzkgjMevJXeQeGb2cU90rHCTaQ
RZo1yFxln73RGMoJFjknOFlAZz0KvK1Y/4vH4aCZTUI8wYH5C2oPScWGYThp4jq+EFOI0niSaXJN
2M3l56luac5U8KUyqqVg8sbqDTZVeXrpV8NzkOk5oU25C5ASAfrdjIFnPzSdXPfX6tIIElvJWJrL
1Mvur3zHLI2iARiwp90qauwG7P5Bt9f3D9ZzACXrjPzbXs/wnLf+P+rBa7eNNa12V8y8ymvxZNOS
VTYkKEuBw2NlW21o/PMS+0m2MxJYOWqV1SwQoznKCB1QYXa/23V5xHy/hjRGhqcYSpkGSvjaYEUT
mntBVz09FLGw8VfNbxezqYyymI8CESxroiFecaiQcKL087Jt93FD3ZM+qnvE1KHtzS9bRTWSPsNA
vEzC0+DQrTyhZkV3+tL2iOOW6gYa3/coEKdrREEocNQkZDr9LglJyMlaFeYXx/1o0GQIKPKNHurV
1fE/TD8vMlMpnJ2HTLOOhsNzLyGv5jTZQAFYBpM+rRUeqp94LwOISnTStgXvSSfOWDxjOFwfZHY1
JSTwXeBx0LRO8JnRWwKkdkXfAbRjgRg9MsMv+RvqGPvasWFTtKLoRlPh5KuWYoubOHhJaE43VLlY
+NESCW5RV5zJ1/pC38EihAM4noXW8LTQlwOUR4n5ZzDiE/SwczEX+i2EItVSNBveFgYEaFyc4eEP
I9fQSsN4zU7U+zt82Eox48D/sfPhGtWlTqc7BR6xsg+BmiJZqY6VMP6m9ZedKYLunH7ooJn7TRFg
5LpnPIz6osynw/bI0MS8yyhqGc6crjWQviyptOlQn9j+NnlxMGILuldTL3DOTnps6jyY09s8RXxU
GwfGjiw4lw7jn8PbWKmOMLCda1VoebT/IwPeyavFUkOd42ixyavpgSjzCC4Vg0F6ZGO0lbEQxmpA
Ac51f0FDte1hpx0o//gtOtQkoTf0UrP+osc4zaUK/Ue1e71EMEnK6BSuPaYk9rmP2a4xOBI7Vj1e
F00tFgZtwUQEcTtRRIdWrRMwZkKUzmyVMTYNKm/PJxSKZcBXESLOB+c0HEtKgSKtDCgcRnYa/TWO
+QbX/X96mxHg/TuAM9j7iQnypHSGkDVvV5faCJYzpKaFqt6LZp9UteDOtZrM9iJNmucRIrE48TZz
+Xqho9fjDM+GUub2DC9Ggs6xdcn2qSlviS3AMRSY09aDPcAybox8celS67o4GzTckxROinl71WCJ
PCYhvahXH+PCSJVSCPV6RvuULezhxHMcdWVK+On50ayZgT4pECqe5DQwRNWwtSjXunEAGn4vdzGz
XjaatNYC2nigDTN3u92q3V6XgSRUZ4ztIjXJaa4kB2jNUJgKOtwDEebrud+Keya2YFMkUWhbp5fz
H5ljS7vxLOhH59EkDS09QS6UMKP7wv8W4KhUZuy46lLfCOjUDtBgB+MVthsqd4++fIXavVx+oCRA
vaa+oBegFTbJN3W5DWIjFM7doVouWyE7wHHkyC3qvtpB3cPa/XsSdP8nx2lgPRHdLbDYGhL/UMoe
SNelF3kSBReZeGR/uTDssQEYUkYaVuaFv/R1F/5fblPTMmOFHrEzSEXIgUh9jciN2+Q+Gevd9tWj
tcCjPN3Qs2dNqFqVlii0Yr1oMtz3O/BTJ7yCZlfLdeT+7YrNQNeOUuHNiZ+cAlE/aM6McxJCLNgO
CafIaxeUIFOcM+Y8MwtHRtNHMZBbt8MBoz+/CS9gGAIoPRKI3L0JLRsnfry5WTo2x1OB0cnu39T3
WHatLcEvjYlk2qlGxIyMDTbWqlo+FJZOI2ED/VlM89a/Sz6OFButU3Bv5o5shBEo+OtI/oorrVlI
CuBPQenmj9adTOJQbVDoJG5ZnboOALET14LXyZ8Jd1LbWcVF03nu5Hu4uvMEfVlo1NqVnmY86WIe
b6J0MzwqJnEAfK33ej9dFcxRWK808wNygRijzjDvpGJY0evK45V4Gh+UhdnsiVIBeqE9pRR4FHsx
2ltr4prATLZMykQTi7EdhkxnzG9nZYUEr6XfuoOK8mv7gcvynY/oSUxSSYLI5QENngGsQCG7KmKc
oOtbj5RkIKZgAWRu6ERHN/9JBlvoW0in1qwbN/J03gFkeUkn48p3YynAorPGmcXS6t/z/dhSEqR6
cXRrfQn/LoJCw2u1ej0IpUO7wXdy2BOHQrET2UapnI40q0n6PqBDvWrHVlo5VKP6URnXTOQ0wMmc
jueSapJB16g5x2gpkQ/gXYbbnoTVk168/h85LgcRIUXXf0oNdk235BNUgVHfYidiFDiYjcz+demG
TqU4VBjUlkkPqEZVI8pAo6GpOj7B01a+0kBdCz6IfNfvCYap9OckQN7d78D+FymM7/Yk7uwUkdM/
8iCq6w3TTdIJQRsADFh2Ru1Aqernb8jNnNyn2KhRmeX15q2MPcPqY/bYAez5FoXWcWhpHzBfhR2Y
l4uGvqZU3wlIwcBGAzyp2bT9bEIJZP/LvX7ZgVXOJ78YjlKciyP0ttXhwONqUDwcxnFO6ieCRac3
8axDYSrQrRAocIoLEo025bdEhteBDfF3OjJhj05+KXL2dHBhnX4CiXAWWADV7jvxjmvBexi5JL+h
f3rYe77giZt5Q2l3gxIvPIlfTtzWc71zDWPxHWL18caLMIrGfz6bNuAvxBtU5D0M7jppJFGiaOHx
1NfY2DX0r3czwrLbU4gHwUgmd158puQ5vPNpPi1Ok8AZPNxGsl0CtaqTAcm8FoJsvczL5zBbNcTu
Y/w+X9UpaHvvFP11LnQWlNB5Oj8fhobQBYmGNyqqugG0NtKxXV/UOv3BQpcHKeLBeBvVTwmDYWf+
zj84GGv442zsA5pK1AjiY36vzBFWXtppNFSIVpMGG5LWfLwYi1MTuOKbrdUjIHtFuHUZKrHug8CF
wWhlzDbrvFO2YoVDIv7xLwNLFOINKpHAACApNLmM6l37xgivuXHF4rr6tmTPXTVK9LD9cMKQGDcp
YVaE3VstdCFjAorVPRQkS8yv/zdfdU4IkW+Srh9E0yEBMTaYvHyUERQQ6eeq+kWtMM5kgkyWIHjW
HKON3qkBDW7ONCGzimdOKpEzIA4PhYXq/QW74SVnlrQgS3XLDSSiNaPtJ+ghTtFzDtAy/V55DpOb
nuTg6HALwznIjTPIyu/DvaS+jWYpXDjKwfTcqTXw0znQqg15Ap33uDZHgWaUgiE9o7VrgwzemhaX
fD82ZGGZRTNeZcR/rGfx1pE9ZCEE/VkjFkSqLAv8nuISx/d4qriJgn3OT4nMz9/3aC9mAyZUdZW5
cpmpI+pFMdWwg4C2vfrcRE0Bn1Ho56fANFYNbhsWi4mGQVEuZ+QFm/EGiG6xgg53m7kJZcrvW/NC
Id74kMpKYmDDmLDng4WoVtAwwOWbYV+DJvhaw7f4CMnKXIpzeybWQo90DpQZCkXC/bnGmC91lavw
QySTuseJmGazsy7jBn+9tLAHbs5DFNsD+qZfQU6L6iATzYPvugvIraZFnpf8JEAbh2zK6d3UOcHP
1kSQUTAVhYwKo1pQRnIMHrQIhnd4sVDnyNnJ1ibk/NpuoEpIOF4qfOlHHEMbQ7hkn1DfF+4xs1oi
QUlH4ewQrz55ECCopN+vZ7YB4ZeWfJD5r1nWODG3Uz+Ui5pS7rZU2ckE4U/NqB+bX4Z30Evko/dt
fsknoW/uXoNedGxGcAO54gkYHYH3kzyn6CzMo7PGQ+qgNUCsyl9QbanRCSLn+JMwyMHwGmqvApmX
UjBNTyoZqfI7o2VrqbGs5lSYH5K52EW9qeYYS1wjDAcSBCHLowLosxWfQUSDyhhurRS19DA4m+RK
MM2rai+k+dzSOaVKpmufDyV6fEMvOZtzcQRnTOOTp/6rricKeeHOTDNKKfiWluF0cBpkCKay47rl
ucsl/eNAf999zmB9EffPzELDc3sfkKtPxm0zgm7XwogbXtI2L2wid/5tHoLz+dFWrq8cRFvy23UP
P43xiQmPt49dN6HKXXfktHqHFjokoP9Wmx6hJ3HgzJDlw8fRGdSnodj5+DG7StwO074c14Rwl5ly
7/ag/Qo9sn7U7CLh16AfnrqNtuE5LryKbSquRfmL/ShuE4COq3qHR43Nnbo2hXLB466xj5pFY1aX
gbhEowSenBFzhbYGLAk3v3rENflqyS0VERx8ZGIfyoau/MHuxWKv/eqJftTmOwdaYC3teo4RorB/
OwF6C2MIh+wqH7enZz5bkW6fD4yGf6QmiUQifHS1AoUtArSqa1U9HdpgWc76MHezpLupM0vf+Vb6
NmM3BJMJjqFrLE8qLjnT/ga7uJCPtIorm0bkXwe/5TBdbqrretAjlWmJLa3aghB23Amoyk8bnfVR
PLkDJIlAnWHGMAzdx1YzC6VHLG1lSSGJbFpWGE08+xU7U3SRxuySoT99rLVKTvxAACu3tFSWMCSS
bJNARqsZ9no6lRNxTA9ak0CFBQB9bIelAr9oBAdWCvBClAt/bbVher/JvDNnKzqCTxwky2LWEYfX
hrXXAsiaCjSWupoB6Htbg5kymju5lE8UwMsuXgAg8qkd9LltQ+j6IULPnemea1dtDHgrl2lZGhOP
aaWrphYtkyEDxXVV0VWbx6rhEmrD8raoXJDbGC3Jl8ZM4x1eqsCv/hfK57UzIr4fI8rdyVJtvAfD
i1CuNawG8Jzbklt8l1uAPWBGv7kxQA4n05XFvg2ubnJnkSsO/GSvhAuxdQ1O5u4YWm3Ly6/av4jG
UgEGryDmrvDU/Nrq7vuOkrar+0iU6b+u1Zw8vM/1tXAfju5/c65cmUyqgpDnk54BTMB38Mxig3rU
ghaFlFhREoyqucx9cxstDqCJ4hsDq31NWoVoZ+6SDUT29ZzcPznPZbR1I+stm1NDpnB+yqmZsQY1
0MwBpbgi4WRhHEZZG5R5vdXoKibdvvkl62Xob/jk3kPINzBV+rFoPGZgvHqFMfH8j5KJFUWCFwq4
nXERNIrApjv4UHvX0Md0Fi8Neujh6u4OA/ZvXLcsUrcgQ5AD8BeDKj7xstdMa+iMyBgmFyYwg7Ft
8eJbriF1vmx4ZS2W7oQX6CGEyxR01h2nMcS9kjbrSLQ/Z0PYmh4eh72HXsPp35Fy7ULli9e3KMup
r1wr3mXKXygSk3YFAihfWhqRXjzOhtrJMJ6+z+fu1uLVkZO6Xo/+PTjU4hDMbOTbbbiC2haykYPG
YEf9Zqo4picYqJHfc6lZhEoHtk19BERxDNOBWNtx8fBjh7VqNbLxk0Vps3JsnPbxaGCYbDL3Xse2
H9dx3FIXaNhQ6sxF9H9Ll/62QcxigreAgAtkowMqQEWHNlFMXlT5gBtM0kgNJ0VXfw0Ffo7d49Vp
qMBCqAkR8kNJ6GBjfkAsrKwd6jjGFR3r+eMSHYpnLkqJ1/p7Rs2hyVaJIDGHhC7G5IfZ4gqGu5jB
sA7tv0h2qFHZGqjFqyQ7PF0RVoyes9Vj2TfD+n9bCEVDiCeH7FBaPbgzhCAuEYXOnOG1AYqeR+iY
eGp/H9pBTgqNFvfUhbFhU6r3NPvRTavY4JJNjTWUi59CShbBmnM2v5/IhK+StG+LKVxfFuR/IK20
zTPmFYno1f5ZzTC7q9EQ/OupQ6OxAb2GH+gc4rZUnNQfPmqFrf3+UJAGJVm2Tl9akwOl1ixcEBTK
bE56zWiXM+AQaQachPHm6RmQd3UDVcRpalOSdRRcpyuRYY+CG0eC9xulSaToHknjRZJT0m4JVZAA
8nuz1mwLtrbXxlmw6f7wkcMdYaEim10is+o9786K5kcVHgBYOKELZcMAdcEEvWlv+xHoF6zRKe5m
I6TE+V5+CvyzrtkEvePph3kuZ0KAzd3FosL6mY9MNFV9Xl5FIVcJfxVZsMw6XuVwSgoQWy/xmol5
f2BcvZpe6UuSmbW/1XYATrHVt77SUeQl30oS9L/AxWZAFJSTBueh/NY13GL5mpyROivDTc5jqO6p
oVIahLtBL7v5Sys0ImOdsd0Vo6xI3vu4CJBwjGK7JERjc5LlQk+SW6XrAq/GT5O4IDEJsggV/Hp9
4kLdmmByRDEMm4VjkIiadneoQt1B28fKACpJJ3raQ0J6XtYwfKBanG8owHDIaA2yHc9uH8nDfP9r
CAWGm/pudb6GJrGVk9812yryFzMzP4wn2V91msJRXeTqgZThFWP93pVk1NgO0CSSC1U0yBQznAoz
qHrqHOr+y3hCLKqsYVR56HH3IR+L8k4fuZxDjplWEmm4OO1yUP3tHSkF1as/ku1zYfnCtZxde50v
WWJWKiLMU6vaTgHq+QlrERJlmUk4QqMBvwlP/26raxTb0aBYB61rLj9tL776t+kq5ZSF6M06I11k
IW7d++0HMJnd6IP4ZC4ozrNlIy17EEVt0asbnO/J7RaajxHWvMkhL0GqrQUAv9KE/Hr2N4vTpUwR
jrFhVxP62JNwBb8uvUxsyaCnUGKKaIg+1FYcmDlhMOTFLTLgU+5EnQkBw4cIpdtGv+TElTd5Be/G
WDQS9FCjUiRbITDkOUmWp/MtCBXz+uRinXPVrB/duvt+6DKuYYgSMcaq9jjy3DjPY54GYTq+Ea4t
iZCn7LLIbJ6ic3nGVYnZOzxZkuPixq+K1axik44JzPEUfm8+EeHgi9PqoWKy+D9IppRrS0cOQ6Du
CZJWVc8Dl61BC6DDnISUlcf8BJJiC02pRvsK/ViNkQX29CApO7p2dpz2kWglsV/HsXnfPQm7f9Oa
pc1X+FuocH4yfGsWKH41rM8jbjhddx5dcKglcmPNz6dzCgV/0JV8oFocHJUARAEs4GAjxfnUr/Ou
DF35lJlyrrtqvH1g6W5VmYs7OaIUAByT6PUXHMjeWePOoZEzJ1kvO9BkygFFM+VaV0G8eXGqC0PN
X0+toub/ADg2uKaa5z1Z3BGdGU5cnMJVobOQzRGaHRqS3WuOsfQqP50fCpYbwvyPPu6fPBf+skWC
CFulxkVeVJeOfGWL6fo7uX+suKkgqtCR9fbSQFMGjyr2/ZPPWLtH+TQY8vuFEVxhaQSa75E45efM
TNhot8NDFoeXxuPkmROzM9NpDTdyNYNR4AYjnJS//rG8Thg3whd3PGgq2F+pmLKTeSPqCgiGFl8R
ysnW/ncvJNws2gX6Q7nattio98OpOUkT7JCDz0BJd9WL1yiXVqP8Lymz6pbbbUmnwajKAAXlKoyh
SneixNuJCEJqms9HcXtXSK/9LVJldU1pehYfrW2JJZPPOSWZFlSv+B+rqgI86yleBMdLmeCxEbwc
VQLVwAnlfELzqpR8r8ubbInT3ClmvMLsuGJvIJrwMUJkd255iYhamTcGKGgHwQ++Z7oc2OFge0MD
0aPmUkk/3uHqR2qKZdKpmZr5g9R9S4k84PM9iZ/soR8TRuN86k3o164oU5V84SdHYIj3ZZpRWi1j
z3iyOCL7lwH6ENWsmf5Nl0TaVBjcYkk6qwPYelwaXX4mmf5yQoocmxW7zsG6bhJXLGygDz//wtrF
gvfvYCPAeFBiSDUhNmOvwj/76KTFeTzwaAgiRDQNB+EajwrwKG1F5pAcb7JcgGFo0qC0751gINB/
RCWnfxJGLw5LcHuQEEoL5q52eQwsxG9s2mDt1yBWzfJPy46PfcJmNSl4swsCa2q3iaxFptxpgTp8
yNOVRdbUY3MMDR3qXWv/Ut0f6mmO58YijpwVYstGADotufL+6e/g9M6zfmyIYJ19CRfNjipjD99Y
k/W5Rz0ZPmpIzI20wcforXgChWjNnvdxyHR7GDPaDyk2bHqH4H3wy+48lruI2Hk/O6YSPjg27ZkQ
ZhbC/Cr+A81XgRP2H2ThZykqOe2E8Phe50g5b2xey2ZJH/Hvqeg4y7HnrH9JK4ORcFI+vRqOPdpv
YK2c/V/0th8o7Vn0wuuwhKWjQiZBjEINMsQ1RoIguqXDsF5J9eTouaTgDuHKO7BTDYyoG8FsNRrx
767ZxGVqau+gfStTfz73zLNJ8KOcD7Hfh3WebR6Q4XiNVoadpFTdxLXxTWrgP3X1rgsovTzimeuq
kC0P/12z6BqLgpHw/GCOAZNOWniBukoNr72QV4A/suVdaJfCgJXzwMSF7oWua1NFO+YpU7FGnxIu
zpIV0h2clC0lk4IZbtu9sNPeFSei2c7RkOwy1wBDlo+cBM3bu4kulb7wnyJDegDQKbm6mzHW40CQ
rPt5mJHVEkmEuXb93vrPxYWQxaTp1l3ndOaHrvaQhwlIOGkCjyPfJoqRj0g2IOkgfxnrBXRVCRSQ
EYVdhfaKSA/QOv/OFlzRoiwY7EkhKnYd86B+VBfBFywRBhnj6xW2tc8ShzrcpIxkuxMMrMO0eeIl
Ur55nGgIUBy2qIukTRCF5WavaF3OVwBK3Eyn5JxVfn+P4V2BQ1tynim9ZTiet1yAjjnOo8xPHHOf
L4uTqIS1orRKcFDl+TJagwWK0v7ZLBEcHe/QtASyB8CqnMAmVTGuV4PxL6P8+r51pAu2P1PVNdE7
fP1frnLAmBGHTa5SnIZqC4wRfAAljlMJiMCChQVkIH0BYOe0Qn07jXyialqykq9+v8TMpPpYu7Pd
9TXqEF3atvnDOMuF30mKiQwnsYxS4qg3NXX/+JpCMAfGM2turh6CP7zuHk6QLDAuk3mbVVs7NAhT
joeKpJQulxPmE3Lu2PtAsrGg+hA4K+U5eSIuM7iigcjUTLtQkRr490+wGhN1kGXyv8cbLohoIFmT
471/oEGBAqUzI2X2PJmrlp5qbPQ2NU/xPDGJCwMWszdZGY8lFGNC6SqYPgZTf8MQdtUwn8DnTmdB
12Ilcftahwagn/jL8K3iOySixKd6pFICx20c18/xDEbOfB/ftqU8zFxjHxudYo1rif80Zi4mtym5
S4o/QmzptTEH0C+0Bxi/tB9yoEj6KnlXmKDlxOElgDgAwbUgsUgbrDgj7+aG45F7qrxNnW9FJWvt
uzh9ETd98nVWpVF03GaUMDlJoDgqEXwt2KlohIb3GMtTpEt8il8c1LPzrLHL5peCnFP7o0p4cKRW
vdIr8CMU/35iiiyBZPQDRfVTyQXmYKDNZT2EeNrJXeulhhLYZKmv2ohfsEBgF1511+P4zcwUADNm
dd7NzzUbZD+L9VWhYbzAc1iWJFn/VkN2nJ0PJ9n4vWUeJg8sso+zbOagEzcI75Z0Q7dLTBvB2Ct6
qMmoJfoZIRwWoLNWIOAHJzS6AAy6OwbKdMS8bO1zBS5+8S5ks7U00fEVdygT1gPLGWjLLb7AP8dJ
VwufCDxEYUGtmiUar0eYyvVjGbgKrbnsfESfGHfvSiWVtTtZiqAyMJVjljk/RyHV2zPUNj8C4Gep
4JgIpcOad4suxmjXD7berf4UZzAjSOcegP7+nZUVRt1aG4eWcZoto6rTpYa9TVy15LCrOj9GP2Pk
sTK3B0WK3HllIz124fk+r0oidD8n9/K9PyZ5xqlQp8bR3qhj9BxyiRzU8rxHbjDZ95js2QgN0CNf
MHGEZChq4X4akjVVVv4iYBMF0XwgjO4GpcHp3HyxODZkFf92L3fbPDRDql1Sq2V4uDZLn4GT7Wwm
ikM5keqZz5KkSuTT+TI8A7BhrwfMPx6diyaLWSOj45Vh2EJ3Sz3Ab3IHXXq2Si2xxWOyZ6u3gH25
y/lcFnDJ9d4C+TmldE9Ugvb+lZRABEwh3xltEp6omKyuctMTDdP51f1FRhvUJbGDeworriEI3MsH
BmXfFuGGoWCf2BajbrZ4MOQay5eGrzQmY5nhTOTNy9pAavHPao5pnO7iCw1ePGnOII2OQEoooPI6
iIqFGo7VWy+/+ehUwK/81PaoAVMtM6XijJ6SHyY/VJFl0Fm5KD5CC/ZgyK/p5Gez3sWOaezIXPr6
t+Wsv2SnegZRd6BxyRYnXVcqtobit0oavlpYeELu6uCU6OPrbcckGfbqtLpNN1lk8MiHrNaQy4VN
CKHKp0nMB1hS2dtjVSvyqteoAsmdNsApPkTajfv5+aYGxfUBMzd0waRepOhUegnzz4dJXgl6aOa0
e28UsSn+pmZHixTG6KuL97UvqH/li1jm2a+WO0o0j3jby/NNLi70Q+tOSwOTM1zGgX1LsK0ZXq0A
vY+VVx2/tYM1cxkikzASSmmY7lMPfoXAjF3UoNlajmsJ6jbN/Cg35BZbs44TTrXqJZWXgL1Ke1eW
GbWHQhv8cNICQFaGlFm3vSEbWhIZ8kIcZwDz3PXLgLbj2Z0FPg5yVnDgWzcHIXXFnglbson4Hm3f
EJzVy6r4BpgC4MPexThsXpqGEsb1aplnbXX4hiRt5pZAVdyfhSTE2zaOMf5QbQ1EPl9g5tpUeaTr
zzuhk68QHWbxn8UXT/AvLKm3t7LGtDiElBGm44O/nHXZ9Uk2RH0stB4rJ8gofNNW7O5DJdfyxlLr
eH+ZoJQhHW2ecqG9DCzJkVlvjJDOlWAxDkPNRsVB4V1MZxUmeWcNRXgE1/UBN6B7PqoURWdlBsyk
dj5BIxWc/LUNYeF6EYt/sJgkeUgIOxZh68lhnSX15OyZJokkxqmmu4Kkf4PJUGBXt/wp27Ykif5A
/vaQMFhzsP1lwe3YPFN7o+xyHDUmDvzFrKQKrqjLMaVFFxmclLzT51JVxujNc7QbPA4fHmBkEIFL
forytb1MWZa9PhR6Eil+sQUKcjsRfO/unv+bv758mW0O0tIHVgyrCiKqE2iqgrq/zIzNaEWI26Um
6PBXySSfSdUp471/k6dkTgaSejGvyS48ktO1HCo8wHMlkYeVi+Y1DAy+2QprjJLr+JyoDL8LTXu4
akTWQTKs+KsRfdK2g/PhyZpARQmgV3kmXwT4IO3U7z/Co0F09wMeaQu/RTLHNvScyY3jqYxsh9qy
EQIvzhDFo23CzptmKqZoSc6stiklhuQvgZxBNuC1M4nJuxklCmd7ouoeKAriV5UhrRn4XgNw4G2e
q97AAO5v5yvv88c5L3zX41uGWmqJmzKlwfWyFEabDZZo8uW6S67ol5enBUIKYDY5+WYBN3E8loUD
a+XhZTB5gnQNkFOTXJD0sSvN+9rEHy0wmsi/g5j6TO8/kIQNINybJRT4GQA9hflz1LTwTlLycDvr
Z1LafpgYcBId7r6Le+NS8KNzLnQFucs+MjGpzEW7eU1hHluWsGH+Wth5wKgi5yBKNE2K2jNq7Okn
TOk2tL+TLjEcBbJeM1aZpqlFCMkIDkqoEY70CjRya7b3M9VwE5+o6XKK06qTZzRSSFVJLJBBRKx7
ekqR7bSwrIbqtGYUhV/v1vB3MbIL6vy8SFDjDf3igxYT9mWoLq4XF11+IOauy69xwMn4B+Rpqkj4
KCaAN+qc+I6Aj8KRfGzJEDnBJ+qR1APsHUE5mNZnmZmC5RdKy/fGbpngo0CZB3ENkL53Q3+0Uvo/
z8hQCeq4Yjrt05A3NgFEORevYtiimU19c51WveEXuYVQRZs9rV43v1xHT/+lM1dcKQYyaxJwLp4T
rHaBi+/DmXZTPFnfdYwqkIcG3Nt5VwT1aDs/U+fMxYsYh3OqTGMRKRjAbewF9c61svD51jYG0K83
7kVYS6zpDiT4Du8Tvfl98h+r5JTr2JFmLdEProfneuUfnZNQ/TxFE2c1Gg6V+XYLfPbtaHM5c/v6
IkPVQE2v2vcJldu6xEUnutdJrjpMzM72IUwoDORe5LkKOsz0SiOUueP+0gLeRsA3cfFhXT6ZNXcK
gU+S0C50GRs6HPUiFij6YYskgl41namwSQrRteoN1WV+lfEibNvSEnpJMyjYW2tAFl571nQ+1cu0
+3uGIQgkBvJvfpKzDv7MqDPlPjcOmAXg7KSxlX94MRpphuOJZODJp2jy47jeI1Q88H3ft8mZbHSg
wQg9UUnrstuH5n6AIeez4r6iAG9Rb8jfJPJAJWZVcP9CCiRapsvPerLUNz4Rn8Slco2vtkPzx94B
MztvXoONnHkR+IOSspN98ZBLr8E3009TH/2BhBqA+3uPSiK9d5iqaGT8n2VsL8lwQxiiocOZqk2e
RTt5DhVafyO504vOdpSLjtSSuFz5i9oflARGoN6uG8Las5SmKvGKa110IvaxahKKZ5tH/KvvOvbJ
jZJEkb5UPDVr62mKZ7dNOI2FWEmzBip85YK3E23UYLlgd/z5rIUjgtLwPQ3WO6ePwZtUCYVhOpo+
OmTGvv4ITpB6Kv1KIe8UWwmpYQFISbA0l9noN6y7W/bXGgA6LHeG9ZAV21prly0W3WkYp7qtktDb
fgvx5H7oZ5SgF/S0E1OzQwm9irxE+VEM/4JCIBTV+iLBG4cStjYjOGT7fvgaDEu9FWFiAXkbb0cS
hmPyGB6AnCsMy07VpZnrGZf3ImHrFQ+SIBo4O/IOZIsjF+wYLjsz/z0iXR5neHc2j5m6oMTtqEmd
zN9vXMBnIacl4j4r6vujdoT39WljW7zh+3gbFTVgQE2kYWk8+Is/UIg5eJvddCsd9jOKRvy1HSof
D3GW39EujhtTLemL0Z2vd+Ck/2zuRM3GTl5mAmI4AwwVqTGifgMwfno4qSyITDOWYDFLa72u8a8p
0DDXHtBY9OSrkhTORbxzRPO8idsL8TojST2S9yngd9ceCzNHt2NiOuA1qGFHWnQgL3NyeJY7T6M2
h4F4gHEk5uLvCxTE6auCrYkHIQIATDFCndb5rqEyzlJTId/Mi1VSuzXv+4EwY8Ws1v8QgTGRMYVt
taB7Z2FAoxztou3Ksx38MwK0+urCCkke2LeaKs9yOwU+cYrY9Dn7B/Fw9d8JmGbi5pQPyxIQVWcA
QxFC99Lv8dt3VaxzeNb39LY0KGmq8G2FZslJ7VIkARc1gB0RNt2k+VJQWNkJWCr9ngdYg3O2cLxB
rJ/aTswTH8YgXqvc6JBLc5rEdqwoZUzWnzu0xrz/GVpaOHfqQMbtT3Ce7t+CaC6tMKEFliia4A4N
zd0XiRVsGZ2VvqVlq1CDppdtJr7IQOAanpa8it2Fxc5FHK+M5EKbF0eeOjcOAes0dNZx8ivuIrZ5
01EwLwXQR0iHNRjAzjz7y6nrK3qumDygpXrRwWypIMwK+iWbcibpTiNR8qQnfUFSJ0blhtMddttC
Emp1beAQ1usc3lEY38ScpkHjt2RMybwmjxq8RG6Xq4Nw1h8rExN9qr3CE1ePi3eK6ot+pYWRJcT0
VQrxe31H2z0mh1zSfcem4Md//ZsxcLH8MWM/nRdDtneEOAfLSPIYvQFJ5m682ihUqI5TkqxL8VV5
KEI9ANPWoVT7UDQoOHlkQ3C+sFjXxU7brwr+FhUXflqgly7u1ywq0qtlqOl4jdPyFWmyGKulzpSv
rc+2/TkGvcW0hvxb1ISQBnOWTUvEYGoEi9AkXWAUQ0WtrWEa8DtCgZsNkb8rk9uJFL4WumfGQ/C2
Y0oqClFOev/LYIaCe2tjVSUIWnYIPYsNwgZBoZ+tzpb5IsQrAMiPw+bFHKCbLbFg/tuokotjN2yf
lRuuqLQLs8oPFWJ28If472fIK2xMC1ZP+fwlDvoAIRmR+NzKXhfTCDRd5Tjw7U/JJfjp06tEr9u6
1QnKAHdWq5blQMqepjU3MYm+74nBftvnNpFbYc0cSnZqN0HTOM/vSYdURSdLXKTQVtuxUil9G4Eh
qJGsage3XPdc76LowKTXb1Nk0xlr3wZ3PcHIly5Z6M0cs6HM4E8sK4JczthJkUccWETLcuTz8Brc
mzw6qlMqj7Bqv7T6c10EwmsG8zwfdW4h5lQmDUWnpGAkF4antECEh0rA6lnwOoWvv4NjJ2BjaWOv
nvSnkNtKPkXltsc68NP0k437ogsOQ+NzskSLM0G3xJK9y3LwvBnLKaFiVzbhNOFR+tWqBimxHOlp
+r+Dsj6BsU0HNufQ3VvfGT4GNlY7oa7inzB/ZL2HfYJCNjYEeqRGYUF6IxnY2IRRGAcqSeUWuFaz
m3njIUgMOYy1rGYwCjgB65Fr+JjgNfhebBLMa22r43YgDzGR2pKotgstcPXrwrzfxL10alTPaan9
Nz8mQZHydE0iqJc+lrbTQdWoWMmYoOj8tqoUCmF85a1xDlplZ1fQ8/jCG9eR89DcQiLg3ZdbJiR8
btt7lstt7BvkFgTI47cFrjIjlBXZR7h5gwrVIK5wKtfRbC/zGGeMTl2vCuOG/YWV62M0j+J2WVj7
yJQc/L/YmYTQsukXjUqLOqVhambGDu6H3dkXRaCEPlAvWOMnOecvdngYEW41iNDAyxnnO8poVxu+
8PUk69cZ1B6cOvm8XgY99vNGeQAfF0bMVty/HHNtrL47YFlEuh0VB4qrQbeUqGhWKtLfmlEHlhOD
Yjl6AIKIEPRzQpvrk4DSXIK98P2PJ5NAespeIPSidfjjNgTBdwj7oR6tM4pVEY7iBi1oU8J7Vgd3
17VHyvnRm2MO18XqDNi3bBDe8WZRqAoJT7hs6ZEV0qiwWyDj17RNg4XmYv0ZxF3IYxSbefaWHLwm
HN7/qztRyqtvCGl/tJ1wXOJtfB5ZXYj1GjKJEDM82+vEfFu5D6JCmLXpIKOXDNFZiG7iQScmY6Ly
fOrtNsyIOn6SmvzUXJOn4xmYrFlH3U1VAopcsY+QkhAj8aux2DVWdaVwMusjjRvXGHqHc7qt/Jhc
/+1I4JH9UAUoB7EkcBrXnJ+uqFrcbOEex/wH3WWgFdcEGPN01iM9POuFNUHkH8HiFqehlW2aNp02
W4O0gkLMkpzas8uvqwGX62dvFFJAj/n6e9grODptF7K59MforNgrnD0YOc/ilonaVKbSdxDj2eSA
3x30jurDFQra8jeyUMrS/bBu10A22z3z1jEsMeLbUtZDsB2D3PSvJTJBjCsiLx/Xszk+T0GgM8iT
zwTgLS4E8bSGszOiSTyBtRNY9/ftskS7TeGggz61US26QvVUZoXtrqBdzJY/+4UAy1ms+feLJfZT
E86R9vsuwkGwFISVc6NyHDMAgTyGCsHNqk4dHoY0djOPcGHiY2WV8IbajIY52E00NXAO6vHsU/db
RY3paJvGquvdMv6+MaIlclmQli0669uhfkvMYrKDk4ayc9Ldk17VP6yTq7B0jY75CS3XMGfZ1DKi
U7hovgwK01e0d4XclnXgVUJ3SppLa6h517tCqpQjMCBiqQvIjqvRXObK+V+nWzOSNKaEPWEo4qNh
hUkTpSifNNN44cuygEXW78V5ZfZXd2kgv5Xxrrvk3JcY9r4s53Iluj7aqSbKnxYcnm8xaEnekDEQ
NNEDoF5Y2ZA5eYS/rawC+q01QDNN5nxeoDn4lmN9ADF2GaX63nAsRUHVYOajRjWy4GfDOchcE5LT
IUElNGyUPWEe28UHb5UEE5z9/J7aOQe7QOtWjUXiEKp8wHEntYVxgqu2G9ZR0mWikjo7tfrcPc1m
W5r1rBB1Jw6wHZOrUmwkFGC0WDUW5OHISx7C4mfWLcAoQppTPVtohBvFNinn4je5+FDsBn/9pxIl
K5i+gC+3uyWx0yWdBeHlFIuPE+29EBLQXgDhKpLZsp4MxNv2/h6qckOvUQ++ID4K+Qm8SVR8htU7
jkMA7eqnEB0blrTZ/hlNUwm6gmZl+5e6Wb8yV2ApzPPvjyh0dhMkDA1G2LfV+p2o/el6/7jvsw5h
tckx3emYp7Pb0gVUsfkvz9vnNaDkx4Di4GvF/Aag+6phEbhTECNmTqgHKoHZpMC6wIora4b4ZVw/
9PujzRlx2bAC9H+Kiwnl4MPQJoThViQBSH4frE5HPXr6+v4DyZ8jPnaucHeublHA5XZfiyq6SJpY
0sh8vj01N1m4nUUIUlLQRv1qdL7gv1TxSsg9VbMZSRmje8QPvZvBooG0bld4hqNKJITmcKRH+zxp
6pMej9OmdXqXA3HktTqIBgr6mAHYcQGEkkzdiWG433IvEXiWLVrW2ufq4515U13iqi2GenzXseZx
Wz08CYXkbwkAoPVyl8U60lZC5Iw+J2pQmGl3sXv7Ed738CAwG/HB+IEqJFVP3IZ/rjtuRAN9XmeT
mLeiOdQ9Cx+mAl3IlzOkMnxIT5Jp7Tm9ssYiE9GhSDkfndjEK98dsBeJRsDelnBWghGSSKHG/XJm
/ZRsnL2/Z+5CLok6lBLXi3PCKH5r/bCuFNNayHDKJFEjfFbQ8trLsLAkC9gvxUBjU82FOIExyqTT
fBx7YeekTXzOIMNZ4xgBhRIsLMnjQeOyixXvPfEKoQddEWE0KD3MSgtN2uBy5nQSy8JkuynLveLX
pmjd/pv4F8m5mu93VweVk9T351UcngF7YZBni0mRhsTf2V9MusNZUJwJSwvRwE5WA/XUjiI3BGMf
nWo9V4HPN+ItdAWpUfIOfGMDS8UKqZSIpBGC6MRpRbIB89lSlBkQao2NaHL+Azx93pikyLB4ceb8
C732O/PFzKSsR/Y6cs2f1udYouyODWcTTvuoFxpV2+ZL22jufa1zVit3j7hrPAw6GkVIK+iyuXI6
sX+HlcTFlQuo8bGNFISkM9HwD3SHuuT1ujPUid7WizA1ZcBfwVJk63CU6MNcNsGAgsx+cZoSgDJm
B3A3derER7Tzdbiqb0idI3aJ570pEnmNk24mJGCjT3w8WRhI7FMzQpPzRGO6aynWRogPJgJLIaDR
n/xwlRUSmpUzW58ODvPCZg2xSEYx1sI2V1PGBj9y+DjCJlOm2kGCeDLVtVEvwxEI9uOc8AWvWQn4
RTbLCTXuDuiKe7lLzbQ0t98nC0Rj2NlmFKAdYYgHUudYCteLdjc5e/YlTocA4U+nHarc/3COTc8g
ImJkBB9ZLU8xpFPB6z5cHbzw1kRuXqw7QPlpb/VFNmi6Fqr0X6oLUAAT8vykAhMhC+SM5v6qqLcs
1TLKpoTz6VuFxFl/JXe94FfctQMdu2/uaGYRqqrhUrs1N+4BrcScTQuRoLbOqppF9SltpItVRDEe
6KGsLgrca/Lp5MiyrbHhfsUp7CImsTDw8oB3NqALD+/WSmIJDgceRz0MzFEO3j4C/Fsn8tT/P/rj
bFBqAZnby07YO3rC5IcXF8QEjSeytlzRLajc9a5dch+gwEGiIueXuJxvr3OWkC/gGfzuk4C81LkE
xC/DpbzOOUXH/+8EI3xsiQlNxMJR/VLKXyI42Rd6D7IlUi0q1S6sweaJetDDUwEfw0Rzwh2WYJ+q
J84O+YOZ2rCQsjISkd48vMkK7UeLec7iN9iidHA+YpNj5elpBFedwS3xj/8XAhcJ7zgDtllwyHCS
R2dgs5usxYkHLOo5oEX8/0akdPZ5xbearJJlHjyePNgt0c2xYx3ImaaiuH2x3CF0KlnJBlj7P0XY
vz23URxcCpm6K0SSeW1Yfi6Yxzua7hPcPcB8Rn1QMQzHpVBRyM+6UeZFcaMiagc4+maD2pSZ9BD2
j3fGWChhz4nB0gvjK7FE9PvysU6kAMxkh90XCNWrK43ymRHD6DGXXUSVXLdzGYV50TD94NR7Y5WX
dHJICjW5jSMjeqtjJSVayRuQtLug9e6KNmnBl7dC8M1kSx6wucP4wgkukyeevfEw3HvUUqq53iY6
8oG6Q2qJMguxWdeV7siy7sTAEobLueuwm+BFfNQncHijkfRMY0b1TiHV1hw6aCcf/MJLufpwrEaS
y+COLd3JTXrk6UZVqTX0XTqHt2mFfhCkViyBO4f0U7mvEfbzzMkpB+166ZLwCZ5L920fCN9V1o70
r0AlJ7HXRYAet5B0rz1NcqGJw3PLybDUzSgVca8AJEz8lZHCO7erdRcIxQv/xqbORXp8QF4I+/bR
/esKKNturbAzxzAZHRUWS49SQdT7NDMXbWMglN4Zp8iZcCK0FYacO8I+jx8bDgDvEhqHRZrgEXno
X8th64bwurX9j5jennaVc98mYnp862mG7XfO28rPKxjx1QyUy3PQXTaIlFkAFmL/WaA69da8FPqL
OlRnoSeH/h0SR4+RTvc3YQ5Th/eJPKE092fKCmkMsPT2s78Hx/YFg7weCpebiPpX7l7R5PFsZy0N
204Tw2LcTKClmbSWhTXtM83KfyHubeZnsMb/mdKX7XAbbsE6e84AoqRArrZS6VSaQwaas/Y5DUHd
/qvxUyB1Eo+jojIdKQIaLd0MP0zXKJgha4eCSOe1eo+FdtDPTtzyHnrISt2i1JK+Y0HY8f5vghuC
YbnEQ/Vy9eS502UvRxpDoIIdBs8IPZnGnGk4XBzVhcMLt4JDi+1e4s3b/L772wELnehgtWCXyppD
bRVXT/Ix7uPKkE6fo/RXD/ybKd5SaM57UdB8RN9rmXIqt+Apt0jcB0E+lbcNJwJRLb7MFvPscXMo
/iinl327jaovX8kalXNkIMAAdizlM7fBWyFzaPvTklbdTPHXLhkT3jV8ZUeWg9E9yG684XF1H9gO
3HOxfcDK/PfKHqg73VFkdm3eeQ5/8Bm8MaqgiKPZE/hNtnV5aqaTwQX7Tj/BrU1OkBNhXyucq7u7
/IeOpn6M0v4yNdsmgHT2CmLMBkY5E+Ej/c8EeCP9br7CoMUo7BiUxTU6s72lHmGMCz08OuSILQr/
inKzmpzIyqQB46k+LS2Nktj7VXD4a2YXMFR52uJ+YSF5ZQuVD5u81l7jw6wxZmgNiEgAN++hl2bz
NwkBgwcmYp1d/pIAsiNYVMEbhuQ/nrVEly3gpKhD+L+D4sHLurnU+Tdtx5ooj6Ldd1uBSVr3NYwJ
Sv6jbHoR1HFU4c65RoxclR0T4fxZsz9mErhuLfwHJJwuuEz1LMbaCeIeOpWADu0P1cka68SSW68l
mcP7fj2aemcH8KWAz9pN7+nj35N5W3qHaQLOmw9kv2x4XtXSS1H8d9Z5nef13gEtHMKUeZOA4C7u
WyFGK3duSoMAJIWzu76y3kQFWSqAkiSgLrxkBTXxi3XFO2WuUZOSaICD9zivzf44ulAn7pdNTyVV
rK17T/6c0BZbc6lur4RKb7/zpLaZ3tYsdDeG9He9IFdMVYX4+rUh38DNolvmozOlaxIK+vcfhcFY
fbFXmP/G4SPxMjcu7Y26lK/mrvpPULKC/bEDcpsXSunSNRGdlZ47FUbuas6R5yq9ThVO+kPGJIGj
LZdHQHqlYeexU4Q8Z+SuVKh/46cze2RjqAa1bVXLujyeq6FVA7zbHF/eT7jlE1mPAFTMkz4dLQr4
SPPkDosyZqxS1zSRuGIK0alaR60mrSiENF/E6suF3Jzs4EDG3VQbR40l9B6GwCu+BZsnTTybPtVT
xE9RjrGdIyMyaECAAHMGAArwLdC+PDvixQwbZ9xO8JBU6+sgoRN41dBmI7DW1NW0XqV1sLA2BdQ+
l+S62z1kZZk47t29rFsioUsQRjNZMIhDNETa2bsF5wI9IGGwAZy85iMBw5nnwm5YyWTxR6uApMZH
dCIIJ6L1XXq8PeC76S/fw25U0nIJ0wXgy6CfjSDf3ySOHjhpfJqxJqzNp+M2UMu/Lc/J3xkQ5moN
p9jx97VRnhjkqxbQhSVrNZgtq4G2oOFQAtUD0bBYHb6OukOQZJCPcxH852EnYRfX1e3k/tlA2A2C
gLAwFWwcIo+pX9etNj/OqGSa6s6lLYJUKliQhYQTHsYyb33kIBvzZBQuDRgsfHZ0J8Ny9wHvfiew
JdtgJXTiyKpR1vbg66H8gnyDyoKWMNDpzD+TAV4Y84SaIh37Tr9XY1XycydEr0NL+3F7NWo2k/pU
xeVc0aBOAPzfuv9qnxzsUb8yJucPX+n0Ww7GE6ncIUaPM5jVsp1G452AJ8qf3DNHV66fv+Dwsy4g
kEQ2QoGuIVUV1BBYuqH6yMxDxA/kN9kXEAERJbzaZNGbNLtsS6psF0dC8svMzVLJiBlUzfK0yJlw
2cc3aLd8ggXoxoSheNin/duMy4DuRm4CObOvj5bZTWvnDzFjCMeDXGDmtY3Ht6OFoNV6QstJ1HxK
53a3r8IffqSO54qhna0shB8u5hYghCE2DAxRFNVUbIIHxLjLNyJV9e871MR1j/AgzsE85qEhB8y3
aqp+j6a8Qz22Wwsukc4IWMipTxgsf7DzYG3mnyZCRAxQzkPsgQw+lzBQZJc7A572a03fb6wzETXI
qaq0KIzdD5K0Fb3jod3fH67zu90Q70PH/Bx2ng2+yvA4xEEvhhhJKM+v0bJI1KduShmrsY9iBmAR
0BBMMzLcP/nVy6tbQ3Y674IoeLgP/8V0m7jN0UFUkwZD/qX97C77QWdKtwc+n475YKU5nOlGBSFl
D0f/iWurfNkNcViuGItIzNlto5bvCoXvd4VFAsTP4tvFMZ2RBOZ2nH4GCHCgg/7I3eqNf9pZIJTr
VHbIT+goKD9SSrw7Ia+BP9sujCLTKKL5gC9sC/aFaAXS41h/44tM5sD0ugSOXjZvFE0GY3uk7ELs
3XGrkmW4luSanzrJIwvhBwA+RH5W5dAGo4oS7t13JtXKGldSF5BK5ONv+GepYCALvLc73C1FkiLE
rGR37QTF1BFUKBiUIeg+nRj15sFy/uuaLSJambbv97GxZSN0o75jxiXhErriXPnFlPHNnMlFptOE
paP5msboViPFNgnjBQwx97jhOc75bbFecbDiFgb1sCci3C43VDWh6wjQCF6V5K072GZnn1YF6237
uUeqz8Zwm6NOPDcscV9H6uC/z/d76rkAt2NBPeeo+7V9PSvBPPqTz64B/3U+gNeVUfCSHAXEXNeM
JoPizdGgXWnDv/+afDrbwWS2TDB/pVq/80Gcbah9OPPlCoBZloME3ubtUU7N/zFAfmQcvouPMzZz
+W5IB2p4KbGOWLMbmO2WOB3JkbgBxa3YZ4FObX99p2MIsJoV5WAM3mVRXzCmqouCilXuhA+G/Ihn
6kaBHNtkjFUEGn0E6OjVvEcBl5xllNXqCRIf8XRShrO0d1tzrWtkFQ8XagAozbauC6GccZsL21jk
jXz1QCiee0++skQE8OLJE6tD31VNduYrbkO+KRyb/lc2RgAj4M48uZwbnaERBakmlFqkpxpHvAlY
+OOl7cJvQeEuETFSx4Fd9FVWJ+8VHDDTRdK6le58aZGodwt7UB3GT2p7AgNdFjzuJUF54VVxG77X
J4gVYxbyIH+Z/z4aJ44xv/Qn0oYtNWjEyaRNFwwfwqXcsCIPHuEcHiVC4BcTGN3tzJGqw1Wck6or
/0fv2osA0w3QLFguavLB5P5Q0R9C+8gTAk9fCkkL7m7G7FX7HYMtCYCpFPb+mxPUnHt4YqgR+pkX
15D/Ob5py/XF/XIDcMGMGcLfUnnp7gfiuw8wfCr3UiHVEdZolTySNXV/aiK1+JA1VJnWpGNm79Se
ZofEt/6yxYwpvJas8ZmIX12/Fnneub+a/36W0RtHk2/RX072C8RCumWFm6g15wu8qUhTwkdC3qDv
ooE2ClHnTwh48dweTO7bTKenJr2x5JvSz6MSoU5DNM1pCO8fSIjXcfGFDVs/P33tc4E6OTMVGUYC
rlIJHhEC1vBre40aEHsZA0QoFqCKemEeFEiga6nh5sv11YeZENh7nI/DfSY66ko+UKoe1lkljTMo
7iQUKnpZQHJbNaFGpMYeDchWolnQjeeEjkZYBe++Pn8MotFKmxTAVSZ3VPiHUBNMCokvxoWsvSKS
lSXpIKpnrSpv8B09vDhlvGwHTWH3aA1Mgh5sGhZmpboQ1erPPIdXevWOWGVt2sx2KDI/rGjZyIh5
pwIPYxqO1OTe6Qe8Ssd/OdLSXrLXpizkyDPKUERkBWaBnsLlGxlh+ivBcIOrDN2H12sRVrFn4oDT
rKjjrFdLaUxBIw/BAzvqga01xerWKQ22SoPj/7LLa9W+ayI1QTMgiGfFbpwDhSVdA75B6c6gJTcn
9zJzMiNIPtMTCHTmTMchBHvNJDZQDGmu0rG+hq4aR+j8H+g8FiD2HKSemLtmFDXV8OcOpBBqFarX
IH/P/Ry0I8JzHKzGR8Mp9ScTy01Yo7G/rx0vYUTY/rd7iDKHOr/1E7rbNha7YLqhh2acqNd9XgbU
GqAKr1dTvC3wYQFxBE9PbyTLJPOW5KF39MdFW45tnVxvpyNztbibGhTeyI/rJr8026t0ucf6dijF
1gE0y/dJDpvBwljWmWjvzfzWOs2KGy4tnfuGRc20UBC/qoqYz9HZdwXeiguBtunllVHGH57u9GgJ
+lF/ejjnilm0cRO7amKCEQSc920qqdC+NDOrc23bPl21t4gYsO1EypzKQw+vqub/vB+4JnCq3Ax0
NFZK8nC73rbQQDj4G850dZQzclF6IJ+BXWfi/xDC2+7EZRfIPbhP3KVxsirlBIX3usCt7ihhX137
qe0t+qUJun0RisWobhPNVmyA/0facjKu2xIyQ0dBDHXZ2fqfzKQKjWQDuxIOGZWnsGwNMYDq7W4J
Cz7hIDpvw9CO0HBtJmHJU8HFHzPPV469ZLy2FMk9JGvqqkuXmXsm7b6Z6wus3AyfxZUvmw2kJPqv
26ZfzDGAeSHf8nVhobXIIAkolwnonMeBpqUZipcljIP1KZ3eekFgCbCH8PrEeVVKRRLi2mljKkPj
vBj+BnLUkJnZmXIglj2Ep9wcBHGOSpKbnHdPPBCrIOip7fKG9WtzJnOrDcqMFDy1QxSOhj+pZfcw
KULinQ1Fr/VP4eQvH2BxRA289tmkqBeCSErRNbTrdPNzia/1HTUBsXfneSo4DFhvm3xRZTcQzI93
/en1n9cqLwEl7VtBJyjL4CDhsqBTrzt+jQQCuSOi9tyHuIyiC7ly2XdBayi76IRN/QHOWXaISNo0
wlK42Cd3JvpPNqNAQn6CTz4oJFSEVxdhuT/lz/uVbLUfNrNcowQ7k74LQDl5g6iNJPhT30nSg0nZ
ksyKrWmADBm9FssfFc+XF3GuXqkbyLGMPQTCdHyKK/TapAMrynSoD2aYWDtDB3L5UDSb6mNq/sOo
Zt7G+96uMf8tH+yrlW2ylbQ/dUNAUT74vZn2ZY0LuFiAWLF0Zcg1j06CFOf5yiz42iZyX3fMYD0V
+pDt3xv4mJ2C27CjobDfAoCYkA0hQjc3oDANZXMy2r3/R0X/nTpQvwir/aSJQcVMQ+iKQo8ziHjT
WTIQXT0NiliRehTHQ4GaS0xXAO6Zp+Dewwymk6aAYn5nz6TVD+9scNlGphxkFLz9Wln3HkKt/dJd
erynQ10dYG9sDyjZ/PyLG1ZB3V+1dJTUbUb4WyWizjTNpYo2WFs2yKD2T+qcAsPiHEUt89bK1Acu
cxCty74EBa12gMsw7+0IQZXZSbcpX0roRsQkx67ewTQS6D+g3QJhwFvDIetx1s/Ti+a0KdkebF56
YCYKWiWyJC20gD4JJWUihwguXU6ZPCd5kf54cdgz8Eyyk5oveKRWpZsdPn5bP7ITqZn3k6/ZrmGj
c0ahAXEXuMY5LgF0vFHIsLJ/o8fR61pf/9qHyuoAabxtK8vp28cvhCtRLXar8D4TfjlefMrXiIMJ
BGp1rIDGkG7jWG48dMmp17eMpmX67q2d0bNB5JZ+zXaIg1qpW4agBtkrOFpsI14LrFAKLa3SUsYA
H68u9pem51hL4B6JSCN22ydVivbmzXZV2AaywUnzt6A/FsFky4JhcZZL/LI+AWs5l42Ylkru0o0r
dU+Tc1iXSRO0TW84v7HykaTUSCilta/c29CbSM7FQhkGNiaU176C1P44vrIcij01FjnmdQPkW+8D
KZrU2+EV5pT+9ezLKZylf+d+ztWjbvK7v+wXpmZOvEpak4vQoRedPjrS/bZIRvfnpuSnhAm7+I00
4UR5D1pRec8JgleXNnIH8otqRx+gbQgOCpTw2ZxdkEeTH9vZ5ax8OTTVdy8ap3zbVjqLOMAB8Bw3
eEwnFIZmQC46grp4fD9pIbukT/veI3msyi3k+qioipGsPY0Csovvup+a0n0DlWuWVNa969uMGscV
gWiNriEx56IYCFh7krbhuxzam/F+ciQZFzIlK11Pq96d8PdFjvM428AY50VS+wulnY8LCFA6uUpb
Ag/CZLWudXTNi/bl4TsilKsj0vw91P1wHUHGdl0jCq4q4NAJeM5Ri8w7OH16ElTZlOb8IcA+cVvJ
5LyJT+esSOOeyP9vIviDsnenD1hUr16yhbHvwSh0v6HRrlkIQmfnU6DyeF37EWjaTzs5Z1IZq+Yu
kxfAWqmkkIKzEfNj/DwfN5a5n5HJLldaeNFYc4/eSCmczCUX/KkpTFTmfs4vlxPQ1qzv8tBv82YN
1iMsfY14T4YNqt7im1y+ft7dSrZzoLT7q/RHIyLkylGjYOiOfp0zPzM+OH9LC4avOY5hXStLyA+W
+s+jP4Dv+Mn/PnggvgZmE83Y51P6Xhf1ghwPn296zpO6ptg9i+cMDYZKCZwid5cZ+/XWcmN46Iqs
7YRBbIPplEu3K4sT92WeYICX3ySATZjZlGU3cvjmlcUSXSAwyO0pZFbXWkfqZRO+SBSEh1WtHE4Z
kIcmWYq3II07pEK7GvS6+niU6/QYHY8ta5pTXN5v7/EWRVP3SYBxsNH7KjZkou4CtGUUluxraexq
j1IAeUPCcyr+UhN4lgXKGzQSgy8sz9li9TU0gjj4giflRRlNDe1IHPPFmz7l9KOnZLj6zanz7lG/
7ECuIOkY1SptMfUjUyNu2iUDBYI79ctbewo+Yu2x9vJCJGmIRfKZQG5cD5L3hS0vfzVh2HjRB5VM
ct02hLddigeqvsIP+ZgFtAtwU7l1EEdiaPJGYPxfhWHzgud/XEdpZR9ofoahqIFHA9Z18Ue9kaCs
w2GFnD2oiLzO5SwNE9LEJ5xXbl7BvTY4vfE04PQJxiUksDO4FsjSGR8Vp0d7CrYMADF5TnN+pTIn
cfnjn/QVJ/r62oGTU/aBOVddmst5L18gsw8Yd8Xw1RvKHi9HITgAEu2Fj9+i5AHtaitsZ17M13Om
0dUci+Rm5mzg5nC/X5OZCbq7lAEiuaKgfg1ysCfn/KxtNypWmOZo2xtxbB3rLX4q5vIlEZdnCoF+
+Jlh2aUv/9rEoJQe0CGreC8l1hhX6jFv9rE81w66BzsvmUGIXWLYJhOpGIENV6XrNZA9iJ+9zuuA
WgfyxFJ2+3Y7+9CFQxIE8LwOZOMEO4R0PrnWRSOjCYjt97pCf5fs9+B1rEWo/x919tSY/ZW3jf2S
jI91Is/3CEwy+NVorbt517+Go/2jkmWYjVdwEflxSj/LKp1styzVgSFEi7XnBXVRPD2vwPIukLFC
OtTdyWKpbtyIHS5HWBX/dANad64s0MZqULRhS/RsvXPUC8gIXmmX+8RbljQzoxKffLvbIrrrZ5ui
dckYSPTfD5fan+5tIGf5RJVOzhiSOSK1ekrKnHD65R1IVK2nJmL/dIInx7oyeAgB8xjDY2Tael/w
UyxluInqNIb+ehO1z57OH8HWwoaY9R2lmpmYB3y03ke+I5hx6d3uEZoctrhRtUR1Xs4eU0HWnKxd
2ATHC7Rc2L/dhP5p024PPwrymUgTzB/FEElwLznNhJXO6lqQlGGpHRhILc6YK87B9Sme1hAlCN4N
TyIapNK4bgEL7mHAiz7nYA2nS+TF01RRDFTo6nTUV9U0+jrM/FtVQ2/gsJG5YJH9SwIWhgyb/0Ub
FGJzV3QKvrEbaTQuAOqF749zzB3aXOfZ55DYWv0/CZY+xVzE05mHlt0fekJ/neVzFEuIASuCV3JF
CdPIzDuy8Aa7NlEV/tbY5AsegvOASvwdb3QUAtRbmKBk+eO7gCYG0XkkJLmnGVYMIuFEGQSVseP0
DQxVWRLt9beJPfGCeq/SsG5S2KvXY+Q9fsKxh0Vy39rqx4vkFs7DTaE+e3lXgPYVhUYP725N7gO+
BTwl11uVxNNIwGfZ+YRdSs/Y8xyLFHAdELAdGnq7X/DTZGdWsDeQLlu3snVO0jW2I8dgLZpom3vP
Srg1lqqdcSC+azAf+PfaIsLy7iM3RjutJl/wLJDGXtEydUMoPYh+ZYAjPPdOjjH4+mnXjhN66Plg
awT3rs0StZFF6jr71QzdxfAaLK9GG6zHhhNTMtHWpdYsCqwOdnsL8fUNeCI8wnGTlrndLe9sje1S
EzvqIaiNlK59RC0EkghLGFaDUwt3ygjomv4P2l+RxyMVLF3A1xkwpNoBWRgZ3trFk0x1v9K2zXOj
jTZGTNQkQZ6ZjGqDz5sI/lMENqtWWEo7/BEyteCILaYD0oxfTTMxpnnv5krfcm0AN0P8wIIcTTWI
kHyYYVkMZrhW+kGWcK8LV7KUUFljtonX05SpIGH9OgqisrMZvNTw3/B1+THsz/fmHyZFMyKtJHzZ
fyW5BRZRJLGpJXsgfUKAnmItEXC96TpuaZnPS6z2ralF/VIVjmZ5XeZFEtGOa6n2pVS67VFbHB7S
byYAdtpIXbNkO+Hfuo7UhElpyDHzNengvTaD8BwogVrkz0Y/GqB+4q9ym4J0AdB3xGezGnxwj0DF
ToWMLIE+cp/z3r8+N8//7ZZCLe6BTKRp6RGpv+UZwxyLFZ2waMQkxz0p5zPe0MqQAZ31D6DX5cHD
BzvlCQux8VJO0c4FmJ1Lm4zeRrc7R/X7FHKgxDgj+zO+4v1T7uWHn7NKjECirQauDcfhoJ4blHZz
sZGAMEUPM+6N5hPPYqGW76TnzQI61nA3M5i/sbGfwax4tmKuxhf0NTkaMcqkA0ry4sweX+qA/EOM
YqumVlNyeEiSu7xZo34YV1ScpsydsmUJOvLwFhnv+ptuva0QgV1PT8UvOFMgi/mVsOR36wDi9GbK
pV2JY+WCHvHEoGLgThOKOi7iZzmtdRd5RnsPcgV9cfdqgm8jyls71nKRVenRgFrG0k3MAn9BvFi8
Le6oPbTT3DVRWTBc9enHGFSRZO4wduRktxxeIyxF9tk8YILwpObYY9bZR2JJSb4HNOHH0luiimV5
SQhQWJ7fcyws8H4zcIppMY9KQyRLlmovSaYCfah4+I3fjXpnWbS+T6FVh4tVP3aynXm/IjF79XiC
jVygYNIiq4q0vN9I+nT3WGQkn5qsIAeFBjU2q6kt7JL8L9444SE5spWONcWbN2J2zygrP2panruO
rC6i6gTSMeP73tfESn1gpMjpa0pyLn1kLUuhjV4fcx2JPJMz6NQoeLNbJUsaSH+KrCOSQbpO1UP5
eP5oQN8aa4KU4okXdWf0unMocGPLNFkD6GTqtgW8TxPjdhU1+cCMs5b0ng/jye8MXCN8GRYYKQrB
pJxapTqzUfpBy0YPk9TahNmyRoejNvMkVN8OMpxu8etmvONS9HI7DuGyp8P2bP5RdCSES3zZbwIH
6ZpKGrkw9Wchhc5MenRkL5sgpASZGGsuV9tYurywQZ3vCtvnQ/TGwjF7xp8z3347nq43tTw/f6iJ
jV1CpMd11d8RedjimbnTFR3nbGIMIiMRDHMeLISP5lXyzT2AFE6tf1P71PTE5Xa9qNTAW9N60oF/
GQb7WiR4Lw/en9pg4mQPoM59g5B4M4xKU37y+RSkXWHr8yXqfjqCoOXfFJdcz++XwJP8n8aNOFDS
xTMv2Knngc3bhbBnFLos8Z3JPLJVs4Bgi3/nBDW+MOO7UGdvmZ3cepnqBlcj0N2WPeiK4FPXnbaG
UdX+BC4VoplYyQEJn3FrXUyPDFBmyy0UnM22EnqKBNQp5URKNrGsZLv7pun5qX+29f5XGNNoyTJZ
EFDVKbMOHcnNaB2tLpHRx7MVpIZXobN4z/KplC1zJwemZOd3s++Q65idbSBphNptO1hXmf0FQLqp
aozlo0K+95K2LKcZqBy2q2rFDheycQg12A/FVOWffNmIpuA5fFtUHbB9aq5qxw7HGKPtSHBAUD10
4PnYZMUxv6QldXHkGC/4k/r2am/wgSLKNqMUvq40D0mOrWoQTZL+ApOdqE5wNbaV3zKUNCznbtp5
jWjPigzpLXTrcTYNW0cTUx9pMdqwa1H22HP4yE/Sur26jikDz9kUNjk0EO++4rF1CNyG6vBN/1/i
xvVaVkwreUVt8dyasvKyX6KbwOn8+yGaq2LmBwe4R0ep6PmcOcevQ6mhfO/2fKdvnJk3O0yabx8o
jSnVfOllRQHtcvnx57n9o1GdkIMcOyD1tn+S9B3V04LzD5JPlRL1yg4ya6SddRxZbVahpkxEIZ9+
l/GlJeRXIaFwUX8Ink0c9KEBBBF9XHTdS2AmhAEZoC4YdcHrnZUcM9Gaw6YAI7+mNB6ftMvkLTL0
Dk36wGw2CRlZYdELv4hc4EC4sujmdS5pLu2mNnsahvehKNP26P1rWluu1PrF7V7NTSiYLrZreAH7
IrVAJrXipPWs01DVZshqcpNdtR/7ftco3/6c9KoDDqvjhIhXHaZrNqcHIh17gmCFeuHh6Qzz1sLY
gLEZOo84wnotwB+lxSiMRotIboi3WXDzqsRGewWhjmbd1PRv2kI5ojT+WrG1kwYuk4JQVWHvpQOM
yctBsBJG6y19GRB4satAvScAShPsBl8FLcY9cvkAD+M05GRGN5nJxZu6G2INmkAulVzoZ36HCuBv
Axtz/RibeaCtMtPdZj/w3Ebyo3lpDvgTCtuzlmGJLJVeOA4Wvq+Qe2l8wYx0MEs3SfQxZ2crHEXe
ENE4O3/rq+8FYsEwI6GaAFBrLK+QzB98UlHW81dI26zPqAe89nIhHZvtx4/FuOjcnvjfDztDmjy/
uupxK6g55Uu5V+NYD5nepIb2qMBgqGJYuVX4GHywOlHUdoSnm4GVDyWaGsgR7f2+5p3oLGdxUhs3
VTaG5DHE0O8aAdMzURBo3ZCbNaVE6ulaLZspq88DdjWDXfnDG5wLfwkIy8OVIK0QhKbv76oRgpMm
uzxqfLOdzzPekFyovrbtuLy7FvFWSKVZt39ixhvQ89c370Lp8OOMd9bbmFKg4+jUIwyuEjf+CudT
bgydxxfilZ4dDihwM1rgjwHRtaRn/QGe9ojr890qrOwLbmGkLAnzgzZ4yilJ4O9nsznYsnKYo0I6
oDIzk6QF//zylGVBSklALjRi8nf5xHJXcJYNN3ZXECJ2Q7cs4lHI2M1PSebXUtqiZb4qUV/9uf2+
SH6RvUGNPxv+wGXQQuT+50l0Flz259Qf1tnAFyQDO77rUcaoiDQn/ui0+IcWCpM6HFa8bKPMl6C1
zQY0thMXKZJA9B1GzZ2zWX9ZQlhflhGPY9M7iriBjIV0VtjlLWEdg0+xzvR0JyaGivNp51KqTpM+
UDlv0dM86MdzK+UU9yiTpgqJaI3CUbjO87Da6NRnI7j/zeEd05jT9XPalwrMGU8vD0jK7U+FnGzW
SmZc6bz4JNGLAtCXs19en82oOdF7+Vc3xMgSj7N71xct6uC2d49LS2xtCAO4jddeE5gF5Cj/AF99
nltdwbVk6Pd7L/XkwozZ9x8ShK38bllNQSKeC2A2TJJYHbJS7juxqwfP/RgsoHA2Q9GgMjgKBs4I
+VDFEISfF4Q/VwKn66VR4QVh6ZR9e0sRsadykHZdcInwlWZ0bOMDpZvlswu1ysGgFM1i2fZQqP9e
jXdal76mgZwGU7dgwKf2Ddm7GGRZuuztu2eDNaVtPeVwnff/DMZ9txE2E9ypBT3+DooW9pqyOyjK
ibxg4FKzFarpk0wi5Ec0ZpKlrIi0GNc58vH8UV5jOZH8yQ/6M7VuolRTELpTkZ0SidwqHPtNpBaK
ibgBfuh4gHbYZ9GX/Rtb8lNt8PBcEtb1xY0lIphA4Vlg0nxZohu8h6Spqg5hh+jiR5k+U7xByH91
NrV2N1k4SgiRmOF4nq7gx4CtzDtICZ1J7QG4jjLvGAO5gB6GwG+7z+jxxrbNO1ag4nAQ7WUbHhub
QWMnB8/T73t/aOObl9f+F3iog/tmyfRUsQaHLersfvqFEbGfdksPRwYxWJg/4cn6CiPKCaXG8wrZ
rMtaf0On7Kz0AzZI8YdJcjl4UIZUgw3moeuMx8sd9VbC6ihXzSIUcoVDY/6sGYCBc8M4kQHSRz+D
YS/3F1fIEG/ckCbvXsHjWvcQxO1/pKm/QErh1VkHPUd+Aj4yzFbqNQzSEEIar+qxVdpalTzPC5o5
igsgFHYtO513EJiqvf29H1AAvCJYztGsiGYFpemTuciXA5fNRE3v57szDaqq7eDLBozZ/3doVAB2
go4hTrlY64IXqoJuXdCM3emBYMO5//lbiQO6v3vL4zEpRzrBhHZF+p3RTlOt86Z1wPdSfrtjDepJ
NvGND8wmmX/iQMR3FyemJEpURNc8uUpM2frFIAstOh/BYms0M6c9oBYQbJooArOIOk7iwsuy1AAu
8fwImVc12KNv2e05ZQ+VQvulyANL0lYAEXYs6iQO7Fh+48LKJa+cq8it5Fqo9PKgw9snkggj07ZY
+vo7meNoDK3qvj2qqMYzJH7q9PkHMXBfRMqmhx89ecIzlgCfxqVLM/z/Q+rODZg9Sd+hel1pc+GK
yfEL3z8uZKk7JNhyu8FA8BeXEe5cFfT/CJ34klN1Y1Tk4E8oBIxzzdpezXtw4wFOuvxF3KBtSN7A
vHXHR30VCDZFzTn9Oqkt48NI1R0/nn1I1UbDpRrDRym2f/1Wwv3HhhB5pgCSJ+dRH3T2+N/wLWs2
Qg9Cu2IzgBmiDFiHZ+bGTSJ0gjDTCKmm6WJPNX48874S8moL7TILABcjv4sVBS+d++zB2RjXgSkJ
OfGStPJ6cToidrPtxAyszcH7rzHVO/ckT/scNrpqslPA231kv9U2f+G4W7pijuPc3JQ8DMseXYYi
Bwzmgp6K9TEEOY7R3hyiLuwtBB9pjPVv8cRheyr9UyVEgUACdCljgmFv+8Sl/F4bIpeLxpggYN9/
hVjf2azS7u8hZKEx//TZOgBy0gqwuAlWxMvweNGbV0qOihdUNA5gbU+8UcjPg6/6sjL1gQSu2oq/
7dPYre8ClDOjMM6vRRWUaWknil05BTzOlid4YHsjpZKkHY8GCZxX7FHeMudFewAYZ/rHzWSGbxi9
dBRSsi4a8OcOPdA0rKJEu58OybmcLtl+lLiNCC3o6JLOaUAck5z7ZWDuq373L0aK1qCppQMXu+Zk
DdyImnYqLg/WEIjZA9r9Z5KuuLBs7wgCTpMjslTOquF3djPdniG0vWoCar2PWQdFOCFNXaIEloPi
wurHq9IQQQ02dOGEIC9WbMxiS9KHMsTpqxvZzQjzso028p1rFcy2OYbSHEQmv5cK86e3gucmCJhx
37KaszleodDPTh42cXNoCcpZLA5PWb2zNzl7+iV6ZP9OGhZ9ZhtGMzZOlaoAtbi/gkKbH4v586en
aaVfubtPMOMbG/l1fNVaQM1ypCtNPslJuyzpOIfdYPeLoKaZYDfokYYOSuKSBxwc66P5qwBhtZdX
WGB/OQ8mA7vMtorzIX9Hbm+V0/w47xQz7E0W4+y6+mkCJoT+Y7fSAhPmWhlHeGaALThrmQ2DCLUq
vIECnlGC8xIXv92BhpOIg97agBDbNPh00Yr3tzqYRjKuEl2TozmAkaUvEf4LuEyEQtkont7LKd+t
Iq6zoWhbbPS666Tg69n+Uvob/fHMknfXWtBIKtVQthmt6sJDaClKbAzWj34+RNxB/c+ZQ1vUxNcB
VgzsHqAYs7hIF5tIRK993/AMRIE8s3Y9TvvQ6CMAD3V43DUTcpwuC3vWjhNAvDYdzkcG0Xcm8aht
qa6po+oYDJDWTpKhZgV4eY+issP7hNqK+97yb/nz6d8o1FHih6eoYWVtWYzBVK5T//JnJ9iu172c
TZXD1NR8FrXYaXGzHM3gq8f793PotaJHJOTed9OKSGMZKyFzCUphWQSLXEf1hOXoWbDqNblvAxQE
2o1XlzyNuoNqmdlljhgafH7Do5KuSrJXbO4ZBrWikFu0gD1jPpOfjAaFCuGFYmkcOXig6KcshW9y
Qghl00ChBpcVZ4S5vIVErnXLJ4Lv2BeJOcZv0sFDhvNMFSszPL0UclggVFtO2PAzZu1ca0b3KvUR
VENAmYj4ceh3hZWgw7922r7LuCNKs4r+2EiCrvZoiCIgSi1uxZZBUEJBGxY32Q2s65Wm9Z8yPvPl
X/i/5GXFrLiWOOLuVRJuLmBzhluPbMuwP4DyG87UKBk61sStQ2otwF+bPr3sWg4ydZnbt9568JYB
sKrj5Qu+sPVwI1RTGxCbeJqKBUKZVVr6H5H05DnE2jTUH70dm+tB6GxpDpRN1pzr5Y584lu28VaH
gRi/pt9sVJBbzu4ZIrTBrtEMavlrSjk/HUb9sQbs56u849SQSeO3IbeLcJyKy8fqxGbr6+noGDce
GJzZv6BqWx3vfeyOk51kjKUQ6look+3ukFzVw7KuedRuAZIEDxjR1tWjJjn280HnpAEdynK+DGck
I8rd+VwBUsBXejbkigccPIgf8hGsY85RG8UsgSh/eXLAKgUHMlm27YNipu3NNVsNavKMAD1b0u+z
tk87sQ+hTsTKoCYSWReszaWd+t3qvimizPFzv98v1yEWNzw39BaAPyV84wY4K24pL7NOPy8O4kVP
4wsv7txXzzSAP+X7Z8qYhFsEXHn4L6OPmCpKQ2uSctdxy8xgQ8qsXWn44UoXBqYR5HW9CyqBa+yD
SfvEPC4OHvo6hUq9yT8znxdKE73QMPJ2gz0eZpx+REH+l6+7HrYM9s+Vr8qjO3kQeh95D14lW02T
BiESdWoJYq6tYSeY3A2FBIk5KQWc4VOorHxom+vq9xL8Yqms7Ms2YgvSk7YqUwx+dZ9rXJ6+aG5m
gHPsixZnOL46w4EbOfpWP7RAugvvCx5o6QWn90pjFF108VDoksrsNXEYItgYk2+0AzBTSpBglAiQ
rUB8b5fS9F6+pt5TPxSAOvncE7RVUqbthAxu5N6lE6//vSJpswJV0gXAsdON9aHLHyr5xSKQGGo1
yzJwt4eGkwPrCdq9m0WA5c2OIXA9CCYmSAFG7rtkrPJ89dEFWaPF4VbJmXPZjY3+7OOD6RTajmkm
N1UIqCJYHuPHAimkXGQXiMaA0ITHKq+81JDDuyPok0lSVWSC8NzzAHYRPn8sWqNfpsL5suM8Q5BN
D5EVhm3dDLiCguXGIvQVDw9ecyC9siGzde8G3fv4waX6KfEg7Akqi0S64Uk2uLX771+O0v9O+R/7
pIjvN5LIE82yEM9IPVOEy9ETaud/jvagcKnKtE/vjb1VUeCoADcEdFqT5o/+gmfaOSqkQq02QFqJ
klgHxVD4rAXmhwN12fXhsBSpE+mmmBK2xcpejeFGMHU8DbVyiMKdkRr7VlbGuKtSizl2J3ZktyyV
Re5VlfrAePtAwmKI6usjCx20OGnMDAD5fMvR3XazNpQSEMJYfLWvbUt1BB6xqg8JUdVEu6+gdn0Z
7kQ/A63yhb1sHwvrJy/W1sK7QZvrVveBX7jsWBuVM+8q5YMwee+3GGjEc86K6BEow3YgM+zIGKRc
pnJ5xcJ92ymsO+78Cy1s6511eDxSTeXR4OTUTD7LQxT9l8lS1tZTZBaldX3TY6JjtWBxnKwQ3oY0
mhRuWtTtXRIijZlndfwbcVhT4vKLffK6P+XhXur1FsgVMfZgCQJxqHy1DQQwz9nF1hSQxHTJAzRW
Jg1datQDO2U9XHOMs+m0HdJvv4WfZOsxwrtTQ2qBSP3EI+rUuUdexLm7dLWuqxpv+7X2NICmDLCw
xJMYMsj3kzPz0a7KPpXIpNJjteYMrrBj4erXvj0S5IMt2CEesOo0IFAgzNrbEqhf1/JJXkejHQ5e
dv8zG1uxdpDYaqjYrowdnpHD0pB4xaOQwxCM424+tK1IJ/PBJom4QcPWYE/L1msFrECGhhi85k+U
Vp7a10S71j/p4XKFu8H3UR6YVHMLBGAOf3DMzE/JxRdIymaT0tyu4XCESwunURaA31O+I1pRDnHe
/UTXDzDkbDIjBhbOMbA5MkciciHGhmmOP3KD0KIGDiEIrq9A4yObAMchSZJOstM3H/Jv8eKNhoRI
RSpI2ebyqcQ2AIqUVIsaLoBW8YDLS0M/YHZ6Ot1TmMgTxyQ/KdGHRZsfTmEE3pdmKLCpuFFhxlRb
bcyZesSLbHqDUI76whOAsL6U4rFoLGwUo6rrl9Ykq8TrV87D288Sm9lP71HpwbVcUv+10ZMZetlx
LPJkRFas2mjvpV4wOQ6S9Nwcq1Dl8e7Gpbo0Yi4bY15/aKBGrjJAAhxKfm+Br/F+bqNXaL30ce4z
9IIq6G9sNi77NyfLJhm6dxRyTUekL87+lOA7P+KTX1Ka6bZuHOBbvw5v1hhLBINGb1awr6qJ9Drc
xL2+E9Df/hlqj1NFxGcAxh1LK61yZevVjq/oTJLDQre44V5h4NHpc9eB9dNj8r++YF10MRTPIoL3
gQfsFoWsIxS+OWnPg6dE+6yUwFWhatGPzM2Jk4r5w1tyufaef0AVf3BF1S3lei6hUlpfy48MnLtd
KMRASsWfMnR9lmB6U8DvPjbfdI0ejhLuG7G/G390EOmMPkmVusJ8ydD2h3yzxOp/GKxzuHBjcgBC
IPK7bSjG1r6AdPZ6PDIpGK+ysJOsDQO+5VUZBZXsltfrCgRWakfrxvHg2RasB6cQqgm/NPVHfcSf
YFcSdl0KBSnYo6vd7cGVK02/Q2VO5egrKkAjefeaYjCQwEeUHVJpTn2TohMpm1XKqoz7ZFFyBfo8
xxPLXUJokKz9D0v9VktG1d7rxcRi+3Y6UwR5w2YE/NXe11KOslXfwVoFaHcol4LCqKszcn7oGS1S
uy/+hKsnlY4nsvlTGCiyA8x+sLnJmNSN2KJHZFUGltBErzy0JtwUCq3nQF6vrydz3SijzpWFxoU2
TVMdF88i9vy4vCtR6RJbop9ly+NhXNEVwQr24HjX9dfHL+lJj208tkul+oNMnsYCk8rwARkNCw5p
iMTw7gmnzdCRnbijX8e6mGt7JfjQJbp6Kyiv7JBnkb4zTrxPOLiV8DJjCQN37+O+If10NOKRi0xq
+4T6boEMOxedZRnsZwRcANfebHJ/56azDyjuKVx7g199pvws3Fj+jJ3iUHWoCfdYd5SB3FSUg7Y1
X8Mk8gk+VhNWwJZaAxgeE9N9RmjwTUVLoFbKi0AjhxhzqGX/0+yLpNCnMQ4HUdG2CCvQJ3gu6pes
ZVmVnltlUXS4yrEUNB7TeZ+7994GqKypINisxL5NElyRrtMaVg7dsehXD3RWSgd5zA6lqrXRnQ4n
dzgYxBiQ/bedyWFfTSmZd0AfwrzZy6jXPSiBtk6Xf+Idy+rmcwcfJ6VrtAUe/yvubrdxwuJ6mVPw
d/ZQ8Q4MoTkvXdcRzqUOonp0Fh6dQ4Fiuys6j2XI5iuecwkgV8pJ8ML34nl/ID+8GNYW46MkkxHn
PyZzR3baaegk99CSDKK/I0PZbDQZmEC3ie4gRtzRaU3M7jZQ0FF4zFqn89HYZ8ldgwoydcl6n1cj
N7tjxJ27+Ol4S0lxoc4Zjwasc1pSb0CzK9yxghg9MV0pXZ2Jm/5RuG9ny+0stU9uhLcjCpOwbfzZ
pF4hOCRHchNIuVvHGgUD/WYgbIKp0BRJ7cmnHfDokLbcNQ7dkZwM5DgHIUuFFYuvjXtAdpmoBXmF
vtnmaLBXN6abfIknrZA8sUIUaoLLnbQJLxRc95HCIpLfVUrWgmHPKUP8cN/6AfryiPXxMQie+Set
JS1fwoVjxHSvq607gehnWaHh/RLqCUUdmdKUDh/HiNzwKqEPMJZBBnjetxGup7RBt0C5b/T7rMr3
DK4AqFrGQIOdxQUnf4ZuHRH6shhF/UZm2c37kIFKlFgNqYMl7dkc/vyqIbtM3XAu1xi6aeK/TJ0l
s0eHuAkosiUEwZl8dcIsqeUFT4xfruY/YXu3PqALfaTahUEaulUq9ehzxRBTK3n0xmdlbwzhaLLN
dQr4Mdf+a5gZdZr8AcD4PJQlLKS+spTZKfYdTjyZYl3kgzF+nocy1uiMGP07Qqa4ywxLD6EEEzDo
2DhoY/cFgBbUSEb3E+3TxIYznOhC3XTfCHd/dQokESG0dXMxYP0mn3D+w4jKxMvAZ7wRrcKOyy+4
sh8sQtSv/9dZymvpUtsfyO133zU68VBGODy6EKmh2WbRRbWrE/NJw2nvSa18wSqK+QWeQuAjKssC
4kSwr+fdH072tFGmcZqj5eh4wsd9UCjc36UHfszHK5QS/8Pvqp4gvfcRphPBKSwDhSzw/GH0vCgU
jkeI1N3ZZRIGfSOEPAROCLuLF9WbveRYTVdDTNeoPnLKWuj1V/UvKyYUaWJ6jZ8WpqCbAaqaKYG4
kWXaCqrIH9zHyv4bCPzs/dYarei/qH566FYIu99t/i/7GWqh6zMC0jXqf4kuAZtpBVlKWDeTk3pP
N6pfQfnDcfqfKxBoUe0m8b/vQ7Bm97ybcb0Zipz6rbf/WiQKao6tZXSjK/+Dwn64ItXgl+28TeL0
YAlmf5jPU7sZMmO6X2KqEbLEjLSxBqD1t13c9l6IA1VcV8wgmnuexzOiPmr5HwriCYKEToIyE0cs
B4HMZAK92JAcTFze1DA4Z6+3aqhBSmYs3uKy9Dz1jMStQNfd7ZeW670VpS9X4uDFLfm8d4YE9Tog
IYCmuuAnw0xXB7Eid+3eorW4Oj8vh6geenb2h12NXoKEn9J1PJ/Xu86XQTqMiGbuqGYKIja/ucuU
imxNWGADs25BAzPTCRt55u+9PIoqSCFSAQ3soEKWRHz2BJ10TTE7sG6tD8NWlnwAeYNk28CA9Qrp
GOVFyWzOFExAi9dnEvzS0yQtiCcfMfDe43QQhwBqQtSPID3OkVSZO2fqvOp628xDIa8/On09gDj+
nEAhlJY81Iewg11znmv+xGG1Jlk2C5gJbKhDboGkvSYCYsA/b29ecZr3HfCqLfiDtq1p8ZBkkgx6
OTrx5H2ZnmnJPgO9WHinV9xuN5jHIvG2RQV60OIxWKfVqxHbAynaAN1Bfj5dCy+RqqQKikL3mKyH
+EJZfgIfT+g54aeVxXdXsb/7lkJDr5+6U9oGQ/9bgX2uu6JVpZYr2B4oNBhiNghY8+PSseGG3bFD
u2nGkKemO7IriFWfYrU+i5cnetoQxuRHsucAiUNg78Lx8b/j04nrBxYJ5li126dXMr+U/jxk7j34
Y/N1mesJZELGkDSwVmYazAUSpXpSU0loh4HFrzEhd6OTWu9LZYZLBc0bOL9xSbRpiuUjagaSDbOQ
FICp6ma4TVEyffZnxB89CujfsvDBkVbudLabCoHI3Avz29KSK42buzM9zxSj8TEW+ZOtCCOYR/DJ
hl9oRVrG6qLaztG/4CUvn+u0bdZDL1yaxqZOy1V+EPfR/f/OaRMlqCMg2FvK/LRt2gQz1pnvthCY
7UMwwOLojC8Gz4ZDUVP4KmahZQORoKxyHwwwPJDkcuMTaVzC6VQTQEQeuYAdXbmYsyH57q9Pp+Yo
ykVjoF26N1r2/B0rh7K1wM+Z49CQmRYMvchr7wm20sGjqT9u34XTu2FxjtX8YSYoV+plwAbKgvvG
AlHhZadH4voCdOfJkLtq31/EdgRlwERsd5qKjbxAJJPoX6ua5V91VZtWkR/gy/RIaJMAHNlGRMSF
cwzOUjhGZV/S3aLX6tPKrtjfahMebBjZjnaNcEofBb7eEQyiX1yfR7Tn9pDffRJmz/LrsG3YqRD4
Bc5hdrvhl0iEAb+P43HnRI1ddzthpn9V6qwhPtGpf2SyB6r/h0teiuSBJYVQhz5bU0G0iSvPjZ2v
Cc1mHo23UF/UIdlmYIRXKvUzZoMYr3CpKCBdIhkt0SbJ5RrxDwmkpbjiYGEUJ+T5ruxT8ZH4fWur
/031oal5twASJPhm6LnHUuUvlUys4nkRyoJN/kTldxLYTgWFvTSqlSlydTZwvlgmvVk7LHZqnBOo
hDWx4g6uF171u9KkkRC6Dgf9pie0DXDb/w3z3BpZNjvNNpT4N93fJW7acyxtAmI/x7ulbzJddwtm
GOqul5n0TwLWc585A9QTu1Jh8ZcoEAbUGkGE7yD9k/cHF62dZUym7/NT/TbZWgHKyncNfVTbr9IH
Iqf/PsopQMDrTI/Ln6Fh0/JAuE61nSCrXzuXudBsWMefrksocQioaoL17VryzGM2vhcPgjCTbIMi
0arzlGrL4Uo4HbuFrVWLTb3SeYufXrkHxnw+xV+xPh1GJe5sPOJ2LepUQF60QgOLR4q4DX+iVGGL
XUuMbeiVY7KVR+0QfxZcmHmt2XVdYaYXF/Z8YpxkiJI7k74CGkSd5pnvX0BKIRhmBq+NckF5edvO
LRPhWMDNUGb0jnUoOklSuSZ66NL76K86RwlzXH9oF6GuCn67atVrtfcVv3QcFcA//wmie4fZQ+09
lMC2HsNbRlPDZ4uB2t2jhy2XPYL9UveksL4oVfivkAw6KCr5JtgHrA8UIjZdVIYREYRKeytdZg0H
gfbixwIh2PiAG9V8ifbztXfPCYkbPjXgRevKzAmlJbriXAMErmuJFo3oP60ndxhTtAkHmvLieZFB
koX9O1tydIX8MfkjlRzfI1MXkG/JCW/iHBdzAE8G6DI+dx6S397rLcyhKQfzQkuFILh7r6azv3kw
Q5wRIgcwyxl1s6Gtibr4jpjpKsc6d3SOPAdAEsPWKuc93zgXj+RVTaf4JTmo8v6OEP1XZuN0sp0i
QqlcJlBMvDi1+Zjc3FrR+LwdraS0Lt4HzLooXbL1wB4STbs24EmuFvdi/0TD1VIyKxHuARQULnWT
aKG9tW9FuZ22/u04f2jRkM//TFsX9cU1Y5B0RwZZC6uQrJXQpx30SlwEg7mi+ziNUXtRGii0F3zb
cK0DvWbiIpxUZwT7UxqzezUyJLcSmKotujlhsX5fM53ywZRjYmyou8J6qqtyF3orJnDQ90jEVJe5
BUIyy8XcsZifdXS6HL7IHs2d1KjVq7Q+X6ocKfdU4tB0QwZCj+z0dlhL1Gy7t2wWGLx2V1hqXeMS
fbw/pF4wnWXXzrUTx4IIw3BOvqiiQ2i5YK1Jckdm5BXxRGDQEFjBEiOm9giuOmwrzL71TWlUf15o
fRSWVecM44HPjxuPwXO+ZuV32+Muuns81unPiWMafqlU63/Nv4Fdp+sj4FvgMplleaQi/io4ZHma
o1VNagnkYZW1ptcsBIrm0udU3qAOAy2YeB4AKdRXdleV1akGWvFwlTnvnqJ7Hov91INRlHtisD0+
huYrrwe9UIMd+NhPEDuSERbbwD1OTBKMTcFXfsQE6p85wr488Fvj7q8CLeXfrZUNewoMmg2VRQcz
eRhUwWW4gMs2IAF/Buzkt8YRS/kjQp+d3X5eqQjxEWGWhVfrTU/A7qtwt4INMymKgi0BT3DGJWxf
RDuodawqnAMUEYS251C4rRWUsM5/h2Gg3PogLrfjQGfxOj6dtfTjL8Pm10McmcUQ+HAkpVEdpRgU
0I5RX8uDehPHaPxlhjabPle0dhN1iwF08XY0U7Gcn1rSISgwF4XhBigT5JJxgc75dr+ht9I/PPAV
9+39OhhGZWp3f1Yv9tw310ciomH6n5Pr1rGNplpeOSpq+MLRPgMRz1iouvLozAz88AGffm2BMtMc
1BfRzBCZwjPnib2CbnDf9qf4NEyT4Nf7PeXoWUNUzcHUrv+onFQ2K9xLLjw/cd0YdjeMk3j+5GiM
QjCKbaKKws9R8Cu+L9UT7aKLzuEXzRGAFqIz8Zq2OZeMjPI4RPXGwF69KcXAzR2bt1X5ZEhqDgPl
5KgMbGf33qizWIMl58jT/OQRSL0Re4qeLIJ43darj3dnn+hc+4aKsfJx/32mMfWSZh9QaNmkqlMP
94k98FlMZDvLqQ3faLo8mnQTBYposVdrsDeROImDKqm7FoTHQd7MnnDaTQxGD+LzDh2cxE3PnaqL
QQockUeWp/cHeGZcKs4Mj42TTaXLGA30TKKiaHzB71c1D3b7ZxfZzDFg4yLu7r7VwhTynHdSTxq3
IxDQMTGU9vN1JUPM3GxGLUr4Vzn0Cml18La/q8hrFY6xZJWAvL5nvj/q5WVC0XnULs8PTsYfgllt
+pBu8cNCSYVuZdSRMOJUdij48lSWm38O/XG5D1aqK7FCQ6B7LUHWHPh6KDE5vjd0FBC8riaF6/BI
C2yDbMf0rUpPq3xwTzJTa5JHewzjTm3XSgNA2uklFH3qiGSenimLASDRKHjeDVn2AvAK4g5QxEHt
sjFlPUHmafUvuK3ENx09FXYVC+PmJ9oFRqMAbIFjT490poepbx6tTcQ9hhGQyJIMj73HAgRDpw2Z
GpGr4bxkuaXsHoAgc33WLqVSqmhMvZM4QRlUe4A+Q98dAwsuzvTYEMiZHGRqtr2fixeKNpYNRzgu
sa37ugVY8Uh1ZpgS4JSx067z1iEHn9KLmYQpTUcGHjwob58bkiKqi3aHTQ+oaybNihVx8Gf7/V8q
Q7OAMrY7SRT4ry8JtULLCnugKbDrQU1EA669vXAMGWELpdhOoBqRDBXfbcoxXESO5BrCu8VFVQMt
yDShzyGSaIEntOHlryMWchrwgWkWsCvlhIjTrjNAWVfC/Dz2nmh7NYb7VrBINBRUj/a/da91owU6
dZ/wC9bmPdW3ND/lrENzAv8MG8bh8JmzvgNJvQCS7j6vUKQ+yjZxng2vUckmWCc4pB60nXCGJPzG
maHe8XolzJh2p3iq4loucuZRC1dd7CxZ/VuAWIScUHxfIdFZ2Ce3h8u96bLh8JH6GcEOOUvlhc/u
OqF0pRo+rxALOA7VI5T8evNgVJ9U8ZL0DYM+VNZRqDipgr3hE4LRu/38+ocvI4/O96KkTebpU/Pq
G7ypqVNJS0LBoVAx0J/TaBJlWnz0Z4GQdDL88ekSPCL2FudThulGp9PSWHYEOnQSzchC6JdROSUf
XnG0ZBcVM3ZejFhuexRnFrGfFl1y/RnKTimTkTUwh5Px/+Y6FG9zi9HB1NDJ6zqlbrW/HrdwVarc
ceCyQxFUXJcKhJgLCe8O5hQLcRm7GRQ8vxuANCoxJg/w0zVFzAz438UgCRxsuLf4rze5QtU6GfDC
FRJrbYihh2Po9Xgclx1On2eykKfl83jpf5T3QCale2mmsD2lOzoyA3i3AOutyCRtnXqqlhr7dg6G
R3Xh3VuC6T6gBnHCPnsDIIo/LeadO52WkS3yQSmOAKqMpaZqUY7tO7ET06afac+RL4qUCiKDLFwO
iF3O4uvhJCCtOHNkPjmcsy8kb/drF1FWPGg+UDeA17dSzvGxH1hXHuafe49D7RwFl059WXdeI4bn
kwyei4+0ps+1IJKvGNyAwgwo3Pjj85UQTO/GEHhbYlPV/fn3/iq3VskGvEqkjPBXr9YEtj0+Eu8g
uHuE3vkWwCVRlXRChTZP2JCRFNMzNpOvDGaRyfgQJtRT2gEK3HgindyIZwyC1aJX/fRLiPT9AqUD
09DF3aoSmWRvjkZ0nOzPcMs9W2iBNnHbHlMWHXe4fUZyyexa3L5qjgms7mY44QpwGnIEzikwU15A
XPfb1M04p9PbPWk8brxl5Dnru+FHsaRoMkorQCab/rw9KQLCvwfugYgYfQI2QHoRA6SFCXlW6njP
VTqN18p6WxWhJ4UDjKioICijD979Fnb0z359OsFe4oy/esf4YYJ84GFmv9a2eTfZV/4wjMQBEfsx
He5DYgn/w9176qY2Nw4QgBHR5LHbEC7k/Sv4Gtvdkv2Cza7QtSeqAEi4rz1xOvvmGuSH1mtHf0W2
NWrzekfIOwheBMzXbuUglRkuWKug9wkIdmeqbft4s1uyrNtthQxaVRxLGlZWWuJrY52T2FtW1aiP
m1lnCkWWYE/mInSRdOgKxMQFxPgOi0F17fxAsKCjqaAlQVezOUSTIazZaqdTPddZTaAuvJ4ZwsJo
jYLK/GcgqTnYcvGO3tqFVtgN1V+LXilLl2OhCXy2d53UZDVc7cPiY6IOaCC3jn08zqqEegKZ7b9t
uzOjX7dVLtc+uFJBvIP1rMHTG3NNmVYWaX6EwB+fXK28sEgs/GG/WT3HssE9Xijo4lGb8Khkx4sk
TlYKQnhzmpT9KGqdNWgpDdB4oLYnyNGHBYsjUgVCe/pnW3wKjFWLvs48duk4rqH/C9k9AuvAg+KD
UR5nCjlqGiwv+W9HKqkk0Lg1pEP/qhqdaRO5h+35YzwM6KOA2X8qpgvBmDTPNDLixTwub1OB+qJq
S3Q5eeQmYTrxgqL6/dPXFerHZ/hcuoA+Wu4zzB+V2FL0KAMDIUF9zdbJf+XUprY6F++u2QJ50VRd
G66YDokXBYWTIaWm335Bp5M8RX4Cu7y7l0mlvmEun5yn6LYoSE8xu7ngYd08zVjGqnh3oVsutLi0
ZgAJChAOf89t61SeE6e6G0cT4HRm2RdHSJ0DU/pQLiA1fjgwKoKzYPA82L1jGvzDdgkaI7n7AfzS
ASnCsZR1u6o7UHFLbfH+okm5LhpiazimKJWmUJihhVhuAtIm3uEc1+xTqXaH6MfreG90iC7ZuIki
xAWQJiCBbeIh92yfDAzCcWeK51HxDpIejG/u4n6+qhTwtwvioX2gV5Tn3aWSiq/TZLv3/ZZs5O4F
5E7YpKxlVoOAKNz0+m82YltTvvDlmp7e6ohRvxqb/TS6PwhJ7YWjo6V7FYFkd56zNLreDRlITyAl
YKv/Ohy7ZqHRSivJvqQCh1BZbyJnXkMuFfh254alFsNgxDlwW7hpoTqG3UFLIJugoYDP8avhiK7+
/RQRWppGa75upsY+up7UGlfj15snpLg4fw2xUuYKa/NqEZSBpB+8gSJXTp7OtuxnB09u/nxkwLb+
HRrGA52levIoBzLzpKgWVv+mUSzztmZReex1cnmpCovXfSdGYiZi695Pbse/xmiBkp0qPGEjH2TV
tGGRQ3ob8iie3ZIFXL6XGBul4vaAtaI9z6S53vTG3x17mOgRzorzFW8EBPB8JCqnseoxOSobhMAM
nX9HNApAXSVZjftxQuMvQeS9/zrK9x3CJ6Ub3vgWgwEo5SCLteM4Lu6eBskzJ1YKAWZIPcp9Ch6k
Al6JMPGA/PHBut9ebRS4ZHjaX/jLNDjO1zth/IxLFQSEGq/k940mOCEHzVYJZhjIooKdk8HQS5Sx
jR9czcZetDmVw7UHc59fHgCfxb24A0rJ0TImILy0u2qt8E7Z6ZOu8ZKsw6+x/lqxWVL6cW3gytN9
kTWFqwm7qJVz8+Gu/CUqKosXxXh8maP8t6mhWnl0hxwhuLtAjCvIA3Kn3APdicD5uoRKY+/yDynd
iS5oGUEedmhUqYChHo8siB1nMsPlJI5iDFjpDC279EDyDUUQh9JFPnktqYd32WrcIGhpAWKxKIs2
DR02RH/TfzM47R0ZDwhy7CcV16/JnTFVkarTEVow/cUYL/WC3Npzz2yPYyIEMaHUre73bgFLe7/B
Y9zgKkJN1n3x7FASA/qYMtGAFac2iO2Odz/dQ2y1QGHdEhFkSGHtiBGq69pCPP/9wvxNxsAX4OI6
ZIS/qoN7Ig+9cIh6dgdhtEdnu1pVcje0yaDUJV8qPi6/bItF5A6nQAFEK2Z714AKiz7TXmIOST18
e9xqhvv6jUyzueqQ0pxmq+gU9dRbMciimp80AGY/wMygwbBjuRf7XjPy1Pvl+tr9jKI3T+9HkVUD
rS8QBqFLDZgLXFIxdGFNbL0MdftjMX9VCKQNo9hrPmGYRXgvr7v3GHThBM9bB3AW9fFBcV8QSzH7
7SVXWcimGSodp9nsTxKeKXvq7sFrwKX/eCmnV+VdzCho6eFgwPrqHhbccBP/0K15gRbkLyn1g3xW
Pejsm6IvxbXhiQ+oNJwz3y95w4mAR0CI+U7F7/y5QmJwJ5Qc3yChoHn1B9LahXK2BMkSrfFvVyPN
pB3qwmaT8KAqWBPUVvY+IxTrFVmQAYmLUV75MgVMkxl4pe6i9X/gibaIPSEsgHr3a7wj66IQS4Bu
ITQ57vAYCM48vY4Mf9ZLYmP1nYQxZ3iCxG8pu0u2Y2AZqgHS66FeCFVZWoTzlkrTosuU9H7Bf5WD
J4w9KGfxxnwf+7xCjOZFGvzrjiL/UEulAnv8K2bcMCnHoEUi/f/or1OaDpd0Cj6QGDGcWhkoI+Jf
LkGmaOiqIq8mCJaIhDlHC9MSjjsHWV9VXnolYd/2eE8iqXnWfxn9sP6/SpogPSUgzaqdWaoZBRbB
keCR58yJrmz525ixt46a6Iry/+rgyKmQ5w2vaGP10DvkbtgXsgdL92uAV9v7BIubFHtt4j3hj/BO
Ztm0FI5Z6rfXTqzLdUcRnjnufENYNOwtWhPTZnRtTNp7MS2079hdHHK0aNFtuNxcQGx5N6/IginM
IvdrOy9uU+MLf9iLKnT7UXv2GKxp/s15maihYzeG1TYaAh1+zxsF1OWB6YqYlFX+vHlWRJjk5j+r
7Segsg0NkEO61BIC+uRKzTdDiNFSfxBWtIBXAX3U4X31jcJUoCNkU6ww/q8ZFTNiT2MzkM0HFdGg
R1cszr5r928Y35TCdGclwvfhnDKMil49rErXAPV3O7iz32qwrRU3ETAuTRyQT4+KXCV1xatX0ktx
Z8h7L/EgBT8QoG4bTrjlmJqnh2brmeaKlUEt91Axf92xPSU4ey2sdogMk8ch3ojIS4Omehzoaps2
9RmUfDSntmntgrRb/wTtrPzh9AzJqpTm0qzh5oXPsb34YXqcvCql1Q1jn8aGHS05Akmt7TI143yR
Ur/hYMpxWlkojCLh4QBwdgxrfeL7q6DZjOvsMf42XoOHqrKH9+evHB28Rs8vx8/JHCjZutMcfBTO
lf3bf/sLdTx7Ma1nVk8Nwm2utBz+VbbcHHOXsr4hUiEoM2CMMbc+Cq187fXz8UBiRhRMOTGLkc34
ePDtk+fStNxCaTSq5vD4kuK/0vFCSswwD4Y8GsnNirhHmYlhYnSHKOYPn1eVN8eZHFH3UeKs+6Sl
T3hJyast3SvgNAJ4yh/G6U5w5XV1pkpR4k8n0PTBxZ5c0qoQ0FTv3743o1UMAI/2yQSF4gqiaQDH
KjUC06lBM8Ddtv/W4qjW2eEp+mvRtixPN5qgy6aUQDrltN1/gS4LbRGrYZoOOaBCQx/LXF8JgwIL
OH5aVQTLpv4/zx1XBWuQWAVSLaLYIkm+3+KcmapMz785cdFB7CEN5OUAPcVzEKVyiLeZbd0PCyfI
k/evHiah9sJS8R04ltePJASu6Pge2ARsJe7CSjOIPo+MgjFROBYNpzbUzBKE0ugiM9XIebZWOAET
OaydzJt2KEdUk+uvLt7aLEspUftssrA90bGgeKK01girQAHGqLLnEWh3pBF1sJscYo313/4r2b+R
6+w/yuL7mzq7bYKohw6MZX4N7YKjgr/e70Zg9FcjtFBaq4TuSj0KMoAmcythoucIShmo1khHFgXf
zyRbZoaUjPj2iT7xX/koXBAPWgBz/FP38o3o5ynGGunJK+zrC8CQUzDRYDWt2Ezc1jj2fnjxqZm4
xRvWtP+1rjOlTPVtjWPDWna7xd2I1y332mTiUCW0pHEuHLFRE5+nbdcei4kjRXiv9rJYrhii+c4T
dWliSR/+e/TRoNOS/d1PNgyIA2qIq0GYZzJpnRFMgVAa8wyHmGcf3XlsgBFfJq5KJ3mPR1NVA8Br
TcvJgZV0IwhyrIpFejFwqdLPf1R96q67ti5zXUs9f8ll0uIKTVISfvVCu0VNk70cnS7pGcFRcOkb
xnUSXQ1e48akr1hm4SbW7R7cUwkS2mn9s/E7HtzHDjqvd1FhlkAPqr3T/aXlnpsoJL+XjMIn4qDr
bkaJ0AqfYgFvBDAOgRyfMR+uFc/Q77UgzXDrPv3NMkk06ZDW670tCCPetYW0KuG2iVSYrt6sdhMl
TKOM7yAh71xNYYIH2UTXaDHTCgegVbMm+NRS0mdC/ZL6bMvKTgrwecXB5wddUPFrAMy9BFrvlqFR
B/3MQw0JXAEjZX2ppRZCVoIeya6BT/gdKMwzVbDhO7eScK2heo8UUEszbgwHu3KhagK2LS228ac5
HApHFgBSDCDuZx3vQvssv9yptUnqRNVkP/fpWJNrfbegvZ/ZmfYqRFryakyjyH9jLV+0kMEYzayl
pZDBzP2Ked8TqmoN2h++s8xD74SbyzQ6nc/mFboXDIsm9o6ydtFW9mQIsnZ9/xK9WbPECdoCH60W
8U2qin6GtLPm/glVsKUpajLKBHvXM/5GnLLb3YE0/7Q5Zng5gs70gDyUZ8NRs5w5/suvlfojo1wR
vLTRIZ3UudhD2pmFUbXvICVrahTOS8yR6YtbpBgSpVJgJTd75qzIqZQCIbg361jncgmkkQ2h7Mx5
1noKW+Bf/ND84hE1vkwdJVjIhLPiQCHNiR8iISDFUgE8BAo+saLM5w5UEX3Im40pRvfzeFyG6hF8
lS/zjK+yqHgvbLajHurlrVBPG81vU3RYDqKSacN3E6hM+TLqtRRJp52QX7PeM9/TQ4MbmPc77OAI
nwX3PuzLZnOwHy246fU27V0lE2nzXjfwmSkmespciMBfsHELcwHuRAAOWmN5WAUv8n5F8Vaokk0W
wpm2XP/YELMSDfjQOWLfZh+mDQeD74ER9iMHme6Zafxzb1dVqBGdKtHWDElHH4/tTY+qTJCdvaie
BwuGCnDk7o6sYiGxNUsfCJXN/UjK6PByAf/6PATY11EZMqHQyHD1TlGswKzDG0K9A6krDWn69+RD
2fS50+7oSVIryxESnxPkgI4G8nhzZou+CGe4zQQa4iVE0G0TXuwtbPdq6s/5cBFeeW74KxU5fk3/
n2NyWIhmGQtCWrmoUcyuXBowl1LbHp9vDDO4yCwjBYcdIlEl77MPpjASH9mJrG77bDWw+1xqss+5
OSFTuSSsPk2kxWciAcOFd2YbEs3v8+pjqOIenEUz09hS9U4p4mlLJbv+9gzEWsXcaQWyhXcy35SO
d8imngeNpe954Hr66qLSvS8eNsAz68i1jzOFphSrVFxCbOy6YRymRsKPaJ3sona0tfhFo0kuBe64
ky/LBSSsPBJNBtAO7oYiVFbKwNcKWlqMu6O2N2I9Q4M0ezIEIYobjqcpUofB+Yms+YBInuZcZg0X
U1egoO/UZQUSsFgyUSy6xzioRf5bdUq7B8WhAFwKz/SD7uB1pu/HMgWomptxcQDGx5HY41TU12Go
OmHgA4IfXfuEk8IO1gc8ML5SdrDxqX3wc6K9y21N8G44Y39vTGm5A+43IaIInVVaVV/uA0j6WmVA
kS6zSK5NTLb7CJZbWJwI1bIKMh6yYXCStxMaSEPQdtnqlAihnvhwwcEZLP8yPlMRZHTv8WTpeIge
Sm0Ncogmow1vgFK2j4vSOD5QnOj8b5/NeYPtgGQIerGQZXOC+pH3PaKeyCsIKQeLalUa2zSA1YCv
ZwF4ptBFo/P7cLBCujK9f7Eu11JM73Zt2cH5AjdObCMNPnYuoWrzh5FR8N6eQaJ08bk8+YMHBOsw
Hsv0vx+xiQGURVTMAgv6QOiKFeJG1ngVA2zR4Y7bw/GmxzcyhRH2BiFyPkEoGZPleuTeeYeTdz5U
no8bwdqJV02w7XnxxT3oUcOxvUFEU1SrK115AmRs4lcH7PfTUDdFQzTE3D/Nfy4i4F5oBC7oVIMQ
DHeRbSr2Sn3darkYy7p3iNrJvlpigbByBdOMe6ce/WIdyZclBZaEUXjoHZhp9cdJAhryYc05HJHM
veoSgyGE2xKUWJD8EHEgoPZzDIzr/VcOyYej+wDt5bH21bZCmZm1Jo5Al63cIbV1fLaNw0ORpPPY
U6Lls16gSQ+f0uvK8L+BjfOnidHToIIE6On0H2itaZPD70hMRA3s6+B+j26MyVR6/7pcu2+mjOb9
60WUhi3BWkUyKZnbDAtLGJNxengBnOu7eu199UGo/teBt0k5KpXNJqomITHF+va+JFlBtNSGNffC
NnFS4tgQoPD4ESnHYJocLTjgYkTaxuPN1Ujef/uXvrHIT9OaCOal/0/u4BG3LgyU9BuMz4RBli+g
wz4vgupJ+2D7r1X8jyALnEEcQ20mUjs/IJgMbbLi38Eb/9a+fba4Ou1+PIfhST8MNE60rPZeGb1V
xSChrOydNbqpt4oGzyH85RTlJ6pjMNLGxTQY4Q/1OXkoGTvR9KAGHND0ZjIKboU9CFScbl4bnHnD
hHGzjOiDjqEyPf5jeiNlzwLv+JJKOx/i4zF3hjfLpFKXZ9mhuGJFX4g5rD+b1fju/mRKp2GO5ZjD
tLlCS48cqMPRh2nodozY8FpR7W0QvCVKtXjxg8dEbcl14p2plWuMaEAMK7D6itLxnriLQBRh8AJd
kKOaAB5pk1wbcy1u2V21Nru9OF/OOk4Ew+PHZiI7q1bdk/17xTqywZgPuufDyJeIxbc4GdpA/EqX
WsX4mHhle8phyQwTiK87rPzC7q8/8cTDzB+m4QxogrKiXI96IDsJwX7TUmSpQym0FbCbwuzoY1Ac
SE1aUBrwZRGeNd3lKC0b1Ia7SD5tr3SAhLiuQGf8aZEsz/ttGZmkdBWoN/JQCH1t3GP6dZviWk2Z
Y1r6trWUP1H1YmJkldvJOb5kyxt2kVAtZDqnXjhPSfMX+dkjpNyOc3+WQgzSt+zAPy5daY9WW7mO
oNUcllQPtklz1hr05Nc7WHBjsRr8RNppMn27xN4bF8QtiLbAzOKcdRR3RIZX2gI+qdUld1uXnB+4
rOH690PihhsKsayZye4cJXGYxCoJS19CEe7dGOr5XAODwDR9bDxYYmF866C2J/CIhX7idTIMR5EE
HYL6nna4vzLX9OkRAk5+SkELDqB/c7HwlKBqulCrr/S430HnRhsRBMzYxZsnwqqM5czuHN9J3RF4
XXLA3Dvw0f4rBXgOed4WjVpsdvsY1+v/TmYtaOFwgGqOfWJjoOggxXuKBdVKUzdroeGikmquEyo2
y9CTViFqWt0QdZnYXqJOYihnd5bLhHxBM8ywoelqMmZ5HYLbWBmiLLvsxD//KTfK07slxzSt88fp
di6wiM30N4Hwhz9IQiNnnTMebZssgte09JeKQDs1fySi5mMfwuJonYVC4OWmnF4fjqQr8/shy/VJ
b6SCuaPZFeBjdh1Pq6eq+3vGasOFZsJJ/m8FuLX+NjlDlV/kupqcRWfpBEkjK5MfzbWOQ5Y/suVj
AvKNVlRy6RBOHaj8lhF7yybrfJD7krbl1QGJTxVLNChEBFREy4HxiAtIB7S8oPwOV7Lg9phxIofa
KauMsFqYJAeN6WUJADmhRa9TbZAP5oYlxezVWkpFGrQJRaXLAzFtV+QNUZQvmvzvUfRcCijcRQGv
cHK7Disr2cYrryh3qNHoR4X8XFSuHMpUe5qOHOli5FVhrK1zv2DnSw+L9ag4nXVkELWMHXuoWajC
vZpPnDoXQqPce9atKKCgs1V5ABjkBqOQxYe+qTVaGpBrDhJxQsaTFcB7/POki+6Sm5GNyIuYbNCw
ikQVUn/hslzhk4FxnAJE1temZaLxkC1t6qp6wttH99Z0Rez4wzhMP1rVDHFSpqqc/IDTLlqKNJR7
LYFtr8wxsKhW2/NLOBiLVXCFZZxGZAQz95Y+/O6JnuO980xZ614ETl2EYqy2tkDeVoi67b4IRV4o
tjQQTiktRZ+CYmF1gsdAlcixrFcGqo9eCuUxxsJFA9Pnbaa8glpR4cWg0qpNApDylkrqg/G9OATC
I1Y3JyTDB6hUVPdtWjCxJWmaEbVYr/f/QE0ui/GX7hYmuYvThylyx8cpSnjKuwUUKbAQ9MONl78s
y2LmTx9Kf43VZHZSC1I39O56QkA2Y2pjNd+Yz3sJ5fctBDhcXkJ3uqqC3hI91Y85haha+ZJZKwbv
noBAQ4IJh2u8vyJ27BS4z2n1dgZasdbmz0RXcIgUmllZxSHzp03Zcsijrjeeca/ButV6JSYTX3zX
cbeKwk0npawkJF2fH8XPhiS+Ip6IMgmeCoXUvjXT8f2E3glDxpeUrQKZdt0U0U20VwJ0BRYj90lD
jmeen1ReBP1bsOoAnPISAmAaneB/MYYobwRYdXkAHWhmbQKwQyK+MbaFXJUahKT0hzpgQ0ggDM4B
JiX042CAOtcQalhLA+IUhm5Re+hwuSVIvnNP3ELuJRFYp/kM9QCs2BXtdMN2uq5YBikq468uB6YF
bYKpUjXXwhB1H3Xj9DQnUYw6usuBFyY7UIIIPOVVHLxpYibn7YGNwQTRW3nhhAMK5ZP2Tdtgbr60
uaF5JaUsoZkY6Q06xlvRhvMaYMWd/sVQay4tRaWE4PwctfV9bF9PYJB0qmjcwXM4ulIZcovZiq7A
nP31hPy5unm8lphqNQWnuR1JTXypsB9Ckup30aSr7USh8o/86HaB+PnZXuHjpPtIIak4ldtBUlXY
TbcEgEpk+0TLWOSeJ1P47fsZmdeibbM8vWz579wfuJNM1eslaThS3erh0NuUBQ2GxZt0ahTnAZXw
1kD6cZoxTY9HRsMLNE6k/aCwyqRuRnq7TJb460S11/qaDO0v7BcuETGhWh0O44pgIhdAnT0wF6TC
zTIJeMIksv8yarvskty3aRXfXxMEAlsx77XO8Cy9yE+5zqhIDgGRUPn+vQXXHPF985yBpaOBKZ1f
v3jsyYfhwwAaI4OLJksXv7qMgaSYSS70UnhQUMmAT/HQ/bPPpI/bMViS8kWkihSdXtkT8Xo9qLJx
R86WuJozzOV3P8gXOSC5wjKk27TmhKkBFcUwlj/wbQuC2t3gYXvFRbbMm+WZnAkqYPsC8AtAPA/h
vPx0LaN5Th6X67tOCOmapbBfy4jminnRC6v3FaDZwlPq4Tu4oBvUQFCOCvCRDgqprvpfpGF90h2B
pkMnSZt/YdKOwYr8j+0CigtKqPIuitSiogM2tlm15vNA0YcbwJHL95GCJBrYsxbbFazfQbCnKlVJ
Hz/vp9yxDsSghFVicKbjGCEWIduyRE3UXB4GbDhQ4dNZ7XwzeGicXqA2rwidl++8oPnbWetpfYUk
o7FgLSod6mACS8NtnqsuL/xplvsX66Lz+WiMDMCobnYwGq1gO/Wz+HyiEDC+XRh0Tpmva6z5E5b4
JPlsNEkNZcpDTCkjDHDWugX12rlntppftho77j4TDWuzDdBxMUGp/voD9O5+Del4PGJTJlFyqptd
d1pxfdb7YQ3Lwdp9UFEOCcUk11ic1VCtOzjVzOCS03EjLwk/p5CKtWzRPxfJFdHic7eK3qWxx740
glIy3XFbPM7RT0eBY177EkJtEflKZ01GFCvhxRwCQkESUJcxmFpKAE3/amFYoM8+iM4t6rfCGq01
AO18hMu8uEx4UCnKgZPHOeNW0Ax46oZMJ7y+eTsdVkAu09tMb6wVOM5PWFROt1uLlJCYxJrsvylj
Qof5cLNS8kxOYXvk8t6zOiLveEl1YzatvN9yU4iN7g9dp3S1zr9rjDzRDqpU2PhC/nZMbaulxQRn
XHXKHvsSKTVTPZI8T18Ca5yWeSiT+KhhhQPzmi2t11Vjm5jgQEYix0Qc2btE84Uo26QlxIbcKUIp
sINRmvIRycIRHJdtw2OkhiuXEHaK5w5ozqjy8svIZWfiT8HjThCTV0qN3uBDXdn7SgHLy+OlITI0
rYxcvXpUNQTvRWk+bmafgrmqX9iwDmAIAqf4BaVKc/NHR720WymVlPakS+DAqOg1u8a0Ci2gCpVu
EZOgzTEI2JXjjYanUvDj1ab23C747hNXLkKISR6n8OAKp0pLI7D7ECx9lj32X4w6I39NbV9IPBRV
vR/wrUS1RFLRTCaEVqKKar3xxO8ZgDDfiXsiH+R29NCdfesr51IPY5524Q8Zdz46kJWhtwyYuGAW
P2Kao7r29B1VKnU1V8Sj8gCKFShKv7knbj7+mIRAYNKj7ZdLFpm06S+isUI1DEt0qMjYKEnmtB9i
vcdDxH+bxU+sc7Q6ebkDn8TUWGd43QwNZ0M88TIoaY/S9bz/qH5KupBjzXaG433HeG8Rt+AE28cj
IgzThNN0joJCemvp5KZ99klBGVlm5Yh/mQlxo92SLxNuXBPjQk1SheivPFVYWZJSTpIftrr9rfB0
mWfP9j2H/cULjV2VrnSjueT95p/sUirvTQGoTXNcOg6VMpUqrKZRQsRTUXwg9NhI8Kwdo1UbRLQB
wTPOWYlmn4FR9hpl0a9fyjHP28QuC3Ay85bbwphbCO31iHflJSXgJLvkGKNpgzGURvYr92obc5vE
w1OLOdZkIMJcbX/PQpIHMWgK5XwDSBr6Rq76K4Zg+WBCoXMI7JEuca5FS3MStaLlH/BQY7GG6Lbr
/5qgGSE1Zz966p6qUjL8uVPkt25uwKfI801wtEcAEHr7R3HN9T12vY9v0eElA+urnGTfw2oBpJgv
zm1kOWfSybX3GkCnhotwM2mfHilkG2bAg/s2TidjiM4LLsk+o9rVpe9zkcUez6VYoUBY+B8SsAeB
Lc5DXwXK+lQ6zn9psD8SToiY/r8SGq5ofgcpucQGolgjcATlXPMQL6OAKQwz5cw+Swe8tsICm3HB
Zw53QzODV1gz3bN/VxK3BFKht7lGFpgKoMOpla426hS7LWXQO8NrI1xAYlKhAeWWWNCA+Ow+I2NQ
sEJbaQS6+dhHHJmhHUpWG061EbstEYtFKIUpYtC9IYCWd55Zq+dKFtUUhOk9VzjQAz1DT3ePYmrX
RMXjBqCvr9lhzGDK+oXwDwI+EArlRKcLjXWcvWhY0mqcfCGruUTZkJJOVM5L1UI4MhcfMopxkTBh
IpNvdYO4tUP3v8SwnOHLmdTXXSw45Obm9l22yebr1QAdihib6vOSZSdjw8MR3LsfNBT3IpSjjcfl
sGpJMDo1qYPfQ4k6v3b0cZqw0cAioJAXQORN1TexLg94KuLrgceUt8CvVtX/tMmHA0ipm/YCmXzn
cyPNaa82Z8Hr21hvFm4R+TCO9uW4Wq8d/3ClS3B2iqC8PMAjqTiCL5A6rvck7IU16JbjR4uNMQYP
D2QURui90AmGzReBeNSsK+fP7zoufLhVKcoosdutteehKZydmdDq7H5gUJihfh/bujirZfaT7lA9
EniIUCFmSl4BMAU3WjNdaNovaU6u5VGkXkGJa67NcPAGBX31vcg8GkJ4uGXEinen2HVXpVzV0AeM
X9rIFakvuHF4fBLojn9yS5K3VZmG1eWsSgxpP0CZ1yIfPwFftu2sWwZKxY8QWbbhlXRw0SHvhsgc
90avxVs8VUnLP5NQSfovc2qeUJp/giqQohOwW4Oq+BR7D/GEPXnRiHXqnUa39NnmsozU1+dbgZs3
x/g1HzhTTXYxjADarZFxZ5oRzuM143gVWONaH5cKBlWWUYpO09/JShrYHLNm4WtIzLB8fbhn2taA
nLosfrtym8xg8RnTYFg1x99/VvFb6PaPsNJ/F8ZR0EAmJO+xRun4YRJkxnMwLBCKl5sBxTwfW3pT
Lr3JuvngMCyzToxIuxWpHwazQC+0ZyNCvL2jmZnVV9r6UBVvLwlssNxx/L3RB0A9Y4lWx7CK0ygq
O7gxxhju2PwA+EeiGaY3Z8eepZfPzXeDIWv5WdmQ8IdmLgftAuq52jv5cFp0jfJOjnyoauisZF40
Ag+46kEHXFm/1ft5HXUhyFLh6+zRmhi6f/TiimHTsJttAt87haQu1MHasZ+RKPP4wBzyRn7oys5I
EvhRqzlGyjhS0O4wjEbbYiPJcC4IDNnurO5lUQoii7H+yO73/x9YRuZdP9gpEqMKGPf8L/rRpI1a
snxr3zHItq0ssuuBr28QverRZHXeZvdpeXAxjk/h61qqVVaWJvmatD3hdLPrXyyKk6HcoWeJkFMc
1G8GsQPekUf8mh5E1+lE9AdhH+UxlOeV1nX3fZCuQ5ZQrfEfxmuo9IVQcsA7W9yl3aN+Jc1tlOho
vaffIPBzLIKK7ZTfAVWVR6zhdJYaaz5liUDNcNNIqUzGqDPMYXua9akry9Eo7bzdxoTVVPHduVYO
DWyIp0oE4YCWsd4oKZYT4foVsAf3XGdeN2TdqFigEAZ+KruOME7pf9J0Opp4Pyu46Fdy5URX5RcJ
HTMNQhFAiV0Z0I514xYTAagAs7COjlDlhCeVzdDu8AdyvVLTXXNPX1qPzdn/+pc+meGapgee+1wk
vtl9cnYC+/jYCmmbjeW+ZZRPDtnWLZsxDToo77RaJ81MiMdPD9qzJ6Ow3T7Fqlu+zWdhSf/7jCGc
4dWZf/0HNTVvFgsgmaJIzdO4T1mEeYwlyhu5ZrNIaERYr78gdpvgO1ozKaP1lV2Cri2tUzcYoVBn
td0KGLBC+tCJGLp3rZegcTSK2FeUFojfl8qMD233hrll70LZ7lqCSyeeaIQP+tIZgICqSbwp8U+O
p1lRoFu7apLZmLcYYHUBSLkCCQ5mKEIMR6tZvDoSK3qLCWFEB2sNrfCZ8Ysuk3dnw2bRYbs40DvN
Yi7l6yo0DOb7B4Dfbzi7hHDVw/usbZReySb/7QjaAuk25P1SGJgqsaXm4a9Q45qLveEe9A7BkWTW
s7CusOQx7DJRRdRy4mcsYuwTyLtVivFcI1wWB+7kZnaSIGG6NnL3zT0pP0kxFssv2D/EozRyvzIc
IZqy4pOroVvDD+RxdGo9Mso0JkGXD1rVm15vd4idiSQcVd7jAD4pTCKWnS29aN2PznE2HRFQHC9A
jnT++TsXOByQ9zg9CVhf4gQKsDALU9hiB6vmqHXkktLVN5Ddw4Jn4ZP3EgwhFLtAyrg9vEwENY64
qHCA12GhUXo/4rDvnqySUlrt/IIe86oPZ6evU0oxUsMiUNDlErvNBE/uTnuwRc5tBigzQWKg96du
KTRuFb9Yh8uDisKpAmKrzid11hWEbogoGSP/T6OrWMTpdFG11uT6wUUEcbIZKFwyqBsImS9mwq7N
C087DgFpa3zINaDljjzFFEE3KY3Uufiv8sK2/tbGocY6gYJrWTDYeA0GyiOClkkkpqIzW9dKoVii
yOkQ02Kj/u33qKWK/JnPnnpf6O46PI6fESHZGhArnsWhAhllaLRbNREYJzNwDtWGiOIb8z1NRLwZ
Ib5iMeEi3KRHvEuSzaXPc3KdxAC/RJCbsPPpyfCPVHOKkSn6JXBkfsH5bwNHBs4UEkadJoMnwZqi
CTbpSeV+p5kGhhvEoe2Wjmy1Ks2jJMb5jVuK6Q65xBEB7YCDHpGeC/fxUBPliuaqdNVi/4d3WOOS
WDvfhczJG5MveUdlzZOyNFOpX80YHIW8vagkTCrvxiCs+Gm5jmiRRhAhvALHrrpBD34j4MHBmM50
wa16a1+5CFwL7JBYFmZ/blXxkMd5Jq9zz1TKqXAXVzCJZoZpE1g+sDpd0EN0jJnNSKrbx5HM/dGs
Ri3SB+rDVy/m83tFHGJSb6fe8YP8GEnaUUxQM7D9yPplhBAv0tLIuOG3yO5n6teLd9mgQTBSs60g
SnRpQU8j3SLXGsye5H7GPZelEI+udsrmXVxkv5ghz95qVP1G8DPWyo9PT9MV92tTjK38LRKNSRgK
rcLAEwZnr69i13DEgg3td5uGKERcn1ra3qhHBiSf0+aVMzJ+iRcM5VGt6ptry0P7m4H8QrchDSb8
3C+lyw2KqtHpKMKwtfcBL+3Tkqc+s4xME125h2dTj0APfllsBBG3jhzOWZD2iUUuTwuDEPmZiMSy
aPdE4312SgftL+Aoh2bJ9qheUSTA5HbH3I7myHm9m0SYyX3egTEdZCd7vJMdNUffgjgm34Xc41h+
qy/1KMygrXNMHyPsKb0EEiBG5LbKt7A2KJtD4vEcpQ/9DIqjjMv2mwQTY5ADjz4SSIcaKPzKD+Yv
jKwV94q4bK/UcMBLjUizpum5tkvavImHA+mov9bFSMXt0j1s1Gzct8ANnt4anSoGAO4mvX1TQjGb
9XNtaraa0yYhgc9jYFVqPN5wgRzw329YYhpmYh7vuL6dRIJTF+CZB3sLK8Dq8nwqr04U8g5fSimd
bEgWdmtVOCdxkxq3czgQsd9IhjhHUAtd1MUHDmOkqT0L5ocZ6Q0Gf+35cjfR14ZzDp9gpalcUrr0
OC8g7PVv8ANYlXE/m+fRSwjWT4wEqSi3odJEnbpF4vbu/o3TG7PtIY9N1BhY0B3Hr4r3luUOYpTE
NuYnAhkFnZAk7IRXg1CXSfbg/YhzAVYEB8HhbBbovwddCFEESVTx/KzmGSB4wBwd76lchM1pldtl
TrXn2mKDsRL3tmOd7f0HrCQ0OJ2vT5woMV+gyCgQpra9dHv/pF7QzKElzh4pVMuhmJG2d8C89eK9
DybaiKcOAMJ6HnNicuPsbnTViUvLaapEPiciBGn87/VgckitcjLhsN9IO0NmanA+RJV4KwvehA+f
TI2hHy24Dx5+wxXIMJ8r70TlOyI2zL4roDX2ahCkA/apoptfi6V2xvIE2e3W19rmoIeh6XesD7gj
GVh9FJ9zr/CoAsEK9UqvgeTep32kAFmfvId7bP2bw5JKcF5yESjQRB3ShlF/yZNw6LiKSY2U4rtO
ISyHn2Baz3UXMjMBt8BCel1yvfAR/KxowaMLfm5cEl9VNBUclUoh4jzsJsR10BpncZtF7O/5VUW7
d7TlmqmmO9Sy9uxWpNSLFD9ucICg8/WuxswPU8LRkKmifwGGNTKXk2eQIZ+HBCsSxaauCHjbL/Sv
YlzZUCWZmbOsSsQeun9pJUz1I1p8wXfn65nySHjwsCFisk31DH2Bihi1lyaxyM5h8kNTEfbPJgTh
5e41ffHSzpWJnAtX5m5IGZBAU/44jpgVbLauusZjXT/vpJGWk04OuY+2yoYWbz4SslGBEOwvuflH
6p66wVedKLXRQ+p9DZt8fmQB9aDl3je7lt4FbHqds7CtIP0+KZfWX/8bOWICpE71FvDZtoKLUd0E
OlnTqF2oAkFvK0Pce+EDBzh/Hwo5arGeGC24bd5joLiKziYQ3agZwYr6BMX0+l4rhod4QAcn6eip
sPENsABqHGnhUQq7CEYDm0yhz4BUtxOdZZwK15lmPpIWZEg8jSqd3lGfQev4HFqYR5JSyGTxM/yI
xRW11fTmO7fjk9Up0ioI3GrEku741ICxVFGMGz50DH+FXUfHWQv+P1OMPtPcK3CJxfBkUskAiely
Q3DRSgdNsakZUt1ss7bDFuRaVs1RKq8jobKzyaWtXc0ZJSJ7tVHxAittsuwhsWDQvB9bqjfV23Po
HiSBU8QraF243i5jCNgRLGalFYCNqSUrWcplrf4Nodqwdap+yQA9YuDifky4RS/kUSQFHxdouzIF
JbgCDhMGoje4gDpRMXDEL15FyDqvejkUe8EECJ3m8OOlLZj0ngidAeMkvO8Bv/AZGMbmsYfPSg97
/taw+LE8a6GscuF3jw9XaP1wMkvXZYzEHXLR2XjMlJ0kGreRFOioWH3/VSxjfbTboa17sfo/GJKL
luGVgj0KG8Nrp+n4vQKboOM7fT+FPXO7XVxJ3uPABGtleZcygTJUMOIySOGr7bNSEvPd6XoS3rV5
q1jiYz5H2uJmLRGo5jKFuUMXAXhI6odLU577aKgjz3pcJ6Qt45kAJklEVdQF9KarjONLdeMVVSLW
nZ/mbN+iipLCGN1gMdf9vmKXUO0puvk2lp8rqk8KseXi8JGRJDWzYfwnEvH9ZVRS6XQJKmgO+Tx/
Cx5gSMY+xaLBZF3rEo1sxoiqGBzNTVK724wvMroZmyTWmJiTnwCCh1Ovs79694BHcpehzxc+znW3
9VSuLTt8cBsfc+R1Q3NHfumv5G1uZeu7nW3D3lITazPIwQLFPRuOwqIDxTCrcXuxJND1kup/AXpx
Z9eCRHeljQQRi8ptljc5YtEY/5sTQIZLIkWlvUW3qRlyI/uKAgqANwWWMC4f59/1dR0KvOHPeA2b
Gb7nGjeAACuIfZGRueiQDTZZsFNjO6jBIiAPxcgt2Lqz5cMdMlvMdRt8ALbLzLSKpmKIhlNDFuJs
9OPSd2pldRdj9u5vdfDOl/4fZ8yLw4G++S4Lk8k8+QfmsG3IvgGL+d9v1RzpbseQCtGsi84tglnT
m8e58rOFMFu5iHMo9qAQg9VXYbN0GPQcrxYWrJ7pdO/9QfHbWv17lrv4+aMOjbF15rRgRLa8ICRR
Oy0HrOsaXZpHMvJBgyOBsynd7R0edrb0Ju1Vj/SJZrz5ak3HGOUC4SGqmZFhsomJtAHeJ9HZpvx+
CuG9GvHgrgb7HzVnkzprklKA6kCTZUX1hYDYLrv3Fj+DtUc+cKujOEYrvH+5ObIkPXCxH8Up/AvP
Ro/cl8579HSkhEjyAAf2duQcskaXwjH6v22MTrc9SEZkH0UJFe2hF0hFLBiafKkn05Qgi4VGXmE/
OdKyWXbJuz68X4ZJ1dCFGWH5gr4FHdeZ3NN15wAZdJJtOsfLz76JyawjBdMSF4JseW3RdX8F+Skl
CiLfpMuNkTpnOuQfup09rAVK7nVvr6+EtfYjxW7wM7ZLuLyz67+N7/dRHldhXOseG5ri9AVGpftB
rgSlZPcqGO3SEGZwQYa7bbtOTF+jj9rDSn27er0DNS6VpXfp6FFMGDWJt3oJXXZCwLxe2afKbKj7
SYvRmg9qL3rblM5u3eUouimzoloqcZF8/5lVAoqbkzcOM+SRYr5IyZR7p7N5uzjbgsVg1qXeKjU+
I69g2J32dZSlPD/LMyBBRzuBwVKSV15MTN7eismGr+ytyditIrDl5I74UTVoIJ4aJFcoaEsn6Ax1
SNN1hVLdmuNCyl/jWZJylLejNQ25OZIK2QXZQnkzx+oYR8Oqyng2skHVKUfZnZJuLOcr4dI/5doo
RUUz4hKaSkDJuIw9bYWyCT5IFvrOnsfahemrk+7s+NvwlHBv+bZ00tqzMw6KanT4U0w9uVgjbU4v
JUab0op181FQ2lc/GtFutR0/rfzE8iK5yXsaSGyPVY5GntUSbNbzBpyHyFIR06lVnb7qIG84D+HB
/V+E5tXg06A+6iMg52igk8oklNCtnSTJLWpnamMF2ZlXJ1Khsuey0xHlT9ne3yIgRv8/Jd8j3drg
u3HJ22uDxB/NhqbsVI9vvyQHG4jGQhyfwVUT3MVMgJra9+bGq99lwjx1bjBTZzKSSlAwnCSwNxJ6
1mD5+1kE89D9WV7ZSInjYrwMCjX3Du76hKCZket3qIWY+YErzQZMdlNgAwQ3LOMJa09IMIOZXrhd
Pv9FurVOA7zqbaPh7Bxw1SPtwBbTKWYOcm+SXLCNRCu+Pwuklhxauh2z1eXLOnuYVJ+SEXJ3KUA3
Rm3RRjKXmCN6UfUl9Iogh8wdio4wP1hXJzgDycU40iLTTyp+VW+uPaPEjjioKcL/mXBghw+0/xk0
EWJ7fLI5JLGMcwHmxYqZEcnzVdgkBjI/Pdd5gL9iphIfqmsNgXmenf7qJQFh/krNKArShKFev9GT
rRZdKwxcIRrdrHr4g2yRK7onNEzbDJkw5/yyw0egHxdVwfLhdWdDZnC1c5+mCHbbU6MA9v/n51dg
SUG90FTpSZu8JeTt4yBSNJb5a+RyzO9CoRqUiSic8f4G8SXRBl06SWSzSiOS3SeGaftxpwshaNjY
FvERD0l+mVru9/NBEAINyZzZzHTVOmyhupAA9B3M/cZTtFS1lp7cDYeO+yTGOjIMwVV8eC7E9bTC
hpQ3I3v7aQlda+MMDLHnnFG80N5NkPqpWz+MDxzqMFdvSTxBjoMWBoDUd6/djxiSnwhfgrTF+Kni
wnHrTbE/EMZXvxeQLzq+6wHBWFb2xNxz3wxYzlFitFCr9toONPm4W5xNtoyWCsnZlEjDqoBHq5T8
TseR6YoO06PBWCVVVwP3aPXfqIhReRWWY7FTCAz3pXo3aAih0P+WDXKFkSJujMsx+YQ4BowWChra
LnWZOpLIUFI/8CT3OtXeDXFVs7vqpYqoiezkZkCiE1cZPJn0ZqzKSx1ViLvK79uzgGXRuxAiNLxb
9eOn3lGANNbd+zwmXAQ5BljcNdxyDQS2MYkzTzLeghb2sNeNm2v9yXUEXuOIRi34Ux7WBUoxYoyD
DWmsEj6ecK0VetLkmZG2rvjgzmVIbTb3im/jRcgl2di0FRvCsFvLBWQyPuhmgwrfnph+IJPpaNnn
Ctl0qvy7WvH5sn0OuE2IE449l0diGWzxzeperhpDSVQ7R3cm/uimo0myHj1bwTLIQXs2ddDxLrIb
ZZ9wgDDQkIKPCNdfopOypSGUpOtCOyd2vfl5OP9Rv47kXG+qVImlqxLVXebVuKtRDXluhlfc5B2v
OoFzyyxcCj64D+DQbkN5ykXojRk6bRurEFC7+0Qete+r0mbkJyTKk/EiYFdGgzZQLNrFIiRPr3ZJ
2+jNXzWlLvSSZdZCz0lQKW2QHlOtvisRxGOIA0RWw90yGZPXngZsbM977h8KVCbztOJgyq1XArEZ
y2Kc8VEXf8gLyY6bNJtB1MYgDvf68KX6lxBf3hwHcv8v0NR7YaUFGLWGJPagum29jHu3TjOl1pkH
UEU3E1ByPex5v/z372EtXONhLJCDMHXRJBE98egypsUZAEvCEOCmnDGCc8d5P3w/nBfANn6kK/z7
8sgDev11It2QFegyo5Ti1fN+DjccOScmXP0UnAMb5lEUUmuFQ+2ATA3kFiE3ZCHuPAVWps77OLFd
/Sw/RXNEUBg/p0vh0a/HHvcFbR8m9qE0hiMsAjYVJcAkJMOZtxsA1AgChtvcHPVaSwn98ilPQ5H0
okysqMsqQLcXBnWfKTADvkdE6HcUpWLFxyG/CmqNo8ZH3+NIMwzshrjg0VcXwS1EzP0TYFAMWjjj
GfNU/ukcaz4i0ZKTSl0KvCcRT8Jqh+PhOz49Tm/4tPFYLHWJbehZeNtRyiu4stpCPLoHIHJm1bQZ
749WTZl6JbRL54FGJMeG1stAKdbV6z51tpj4bp+DOs91Uss72d8MLgVqbJvkra2RDWDpDhbLzClT
hdt+htHzFsi0sD+OKr3TR2eifs/ptToyeTsH1ler8+QFzhkNoTsslZoOVmihTX0NCszoe9QbzLtw
2lDLktywMCyepbRVYC6tVGIeU1e4mri1o+fL2cSeUUTiup3iDSbhhgXYQ80HfbWcXEcr+VOHdwt9
+pq0dlDTd9rxNsm4YsR/c3/+a+4vcdYs8etW407ekwfTYlGllZP9bZMkpLijWSeKu3Ox7eXh797p
uom6MgQqRFM5JiIV+0Gk7zEuIfZ4UbGAmteJXmrBLpDTn0fi2doDk7nMCpX69QYi9xHpvziOAb8Y
cTojDZ85xt5gT7HpEhCAdua5zDheMxAlDj3e2YPmrYI+CVCEWsYFNHpF2AGACAmDP1iwrexpcZFQ
gqMINluC+7mP2QOVuZHmS+z5NTqO/2awAL/Lg8l89sQAQZ0DhyHXaMKZts4kXx6pwC2ehdXEPD66
90ZzAvdNqbG7+d+eOyFXuQXd9a00d107iqlND89jjF40Lian0du5sksAt/Ivfw9vMa16TghtyFmq
H0Vz3mEO845o4/yzuyMRdw4JtWETCafJ7eORTn0n5ZoYg+vugnckc2Zf7rG+E6i3cox5g2p2pSlx
JbLJoRpAiPBJ2QqNAhVvp6sq9PkY4C1O98a6CwWaUcrGP55fF3O+bNVRiX9uHgnobDLCYGWJuVpH
8E85KQesiRnLoy2N+K5Gak7IHo1A8lhWJBFMpGr+Io8pvUeYq0LUixIhiSWc0xxa6B7pIAQUQeH5
U42IAsflZLPglvvjs5LyzNC1mVZS3+fxP05F0DIQ05s76uozye0YJFUSEGRVsJXYVRfSUJkI3seQ
XsPAY86+QASfyIm6z/r60ANKBnFIjpJXH3UbPBLNIgd2X5XbjyLS30bD4KQYdYvftRjqisd5wDZ3
cbcBGYPV+a5RGyTume5dwA9oH8QUYpNzRZu8G87KGvnZZgM1hykiehUHoKPWXA1EGa0t+iXUuVmB
gWAQVAjHW6yiYIjHpFaFSLWs2/oQltFohUIWVi0pMrbX/v1I7zUFPBr0xIYs/eC76HG5b+PEmgS4
7z7LpHbw2vLVynGXt+01efKaCJsZO4/7TR+Q+Ee55F+uVZL4ClrEfId7tXHlCzTst8UTiP6ah1Ml
nAVqObHuNZudlEwXV0L0JVXh4S54EKdmkm+/O94eXT9/laMH8dNHvVhwlV4ji23YFCWoNqhLJiRd
7MjiDTpSLRo9NKiK+kiZ35CxTtz/F8Roxf6x+v+dHz95M6vpjDXn0GWqDFfisNkEctX5eVzuI9T0
1hNNlFijUsqHDJKJB4b/vnrxiYDX/6dm0zG4NCaqSP27ykWM/CF019bMulSjrgxhhkvSHcmQOs/+
4ayIpLvLRO0/3W2wcm3FgIHQHBBCRP/yyud1j8pfT2gwv5ikrr2upLOemi87cdWgN9C/TU52hbyu
dOORSDKaq0ExUb0lxnDpjBFSFwvnZ+E8KDRdOQYd7Cjdde/qBNM7rc75TPcbNgkCp1TRvkBBfx/s
Lvfm9Mrpxh8bF2q/Oknlnh8iNeU8iklwwXM4kbZZvgwalX6DL3viAqn7FOtuAHjYeWbvxVUMYJse
KT4UaqncrFL8vWFsQqKe50kZVAxatltEIOKPdIF8YqUM+fZj9Mp/OrI3evqPVE91LqPI1FDSVZEf
bVwHr2ZcvFvmoYng7vLn9CUhvBaikLWKptWnQO5xBjVDLXUF42pJLQIv8oA/nWVSVuxzxjaKDm3S
I8pS6OCMUXT5zHz67ur5bwTrak1NHFtlbq+S8xw4T/nvwbTDS4uY9iEJwSYJ/goA0T9XryckV6co
oYFK4V6NiSYNp4OoL5jY7KS2qLfY65q4qcKeTViaeWlGjmCubbuU02lfKtdoV0Wph+p/1y4ko+w5
vuIkoXAhiYDYHS9r9/7nH4ykNI9Qep9/yfCMdWKXLNoKVgwr9TWEYy4MNagdTede6nRbRud6FAXe
2jaANayhbbt1dbm1eWdafXBoxKvLk2oO0j5jKjQhB0yg9B4a5B+3RxmyO0H8DCBNqnzMeYOC1Djq
LBgYlj3TvwCX9KPNYzS4N7bK0eeNAgfgUPbc1yWZBe8vir3yfbfOiMZkYVnOhTW2iFUSCd+PjePF
ZysUUNINpgx5hP9Reb+CpPL8ovbDMgxrgP+9vb0A32YSEgwp9Z8bAe6C2kCwKuSXPhrsJb6Opgrx
nJR2r2WzCTo0c1TZcMor6WPWHUmUNX1wNjxnyKx6z3VLjcNCqyRyi76KObdY25wWeRJWaGHwYuDV
O8XosH4+pQRNgGvCvXOvk4z+mglcZD7xZu7uUEBgrp6fsqqelSoTcjmJZd4hCoT65VOwTVB3zBX0
ob+rWtq38IK0y9ru/G7LVc/bebRbM4Qqh2v0ul1B7x6Slsa6ZK4ZrQMxEydrqH0MseeeJ8mx8Zu2
zkz/DFCBDH8KtabfiDpZ1Fm62NgWIohyqX5SCAQq7Boqun1zYK486Lx6i7p72uy1tuxTE/galUOU
YhPw/N8/8zl9I1XctcMaJo4GoErQ3Szz5HqQljz6d08Bhp503txQmk1jfA8q/cCC6FgX6GOS8fzy
B82UygWlWeDpvJWl7BthoBcC+PN4h6SSZHUi1zzB17iRFU33Bf4dA++xKWTPEsOCgM/HggT4EFsf
29knkK+GFCfismiUVjUF2vJTHvHAgCvtzMNWLUTxLfL01zoJJSCF+UNDaaLUEdgOxoHqhNy6s9pM
MpRQG80JRNoTew+IrMcIFEGDvhzmNrllmveTCtzY0o0qOVRPm4Go4n8kdttS7pIohy7REc6M+x4D
+J44lna5wtfoR7wcBVVbTRQeocefD7Tyc2UpggKi0/S7vYY5lYt0dxVXr1OnAsc9gE8moEsQZZSY
wpT0hUXLomqwnF+YduAbhwRqF2E1M666A5uKh8z/aoQtuC2vfW8T+qsQzaowNjdxaDppCdjyyq6r
y3YINwdSUEIpmoZ1Ok73BSE8Ehp11ECqn1+LoAe5Hnkd5dR6XMmh1YGFDhmI6EMQrnk1soO2fYD2
rj7zyVSEJLTiWMz+9BA9ZyOrQ1IDoOK48xe4sxi/Txw9P9i/uNdcHqshlsQzyR6q19QPEQiETaSG
5fGskgPKr2QLKv3UzLG4GEanJOFE4SjDBqgFm/AcKBFU/FUP3CCi2P6mECHKc9wAVH3qU+uogL2l
hmn3fjuIVkQnUPnMZ6vGxA23Gx6Ny837eq3DRCXA9lz8E8OQlVIFEsUAH2fjpXDuLRxTiSt/bAAm
HdHnzhraI+D5y3Csn7x/gbl1jkIKhBUzmbu+tlfuC7RgrqDHjUYgcyyzmFVTUpn7iWRLaYVlIH16
NxYHW40MgTjhMutTTLMBPxa+7Q8xuEdY8iQQx+p+hm88Zbw0lYc8tsqrmpdg9Qg79bjp+xcJKK9+
BXNW14BvnOZQh8Fk+EytU5wFQu1lqd+Zmh5rb9d2q95ZzdQngA1Hc31MyXB7NWGoQ4O0gPE9xmqx
LeVcz8QYEVB2F+Xy+aJ0S+YLj97xHeWuBEeEoKkMMKmqyNSwKDH2nNzcXzpRY92uXkd7jln0GDTD
Us/a8ic0XQJJhIRAYcDw5ASQuV9Qeewcs/Nvw/qDF81iXx/lxRy6+5xik9UwbjExtYMSDXOyW2Lb
OW04192UN7ddIgjhIM3woBYC5ZMu4lD1rxCNCAXrPblkb6/We3FhLiTIOXV1TY500wCG86oJPPfQ
UuLGBTi4mdwesF5mt9Hdg1PL0emmzeCbJNMCRaKzdWrW30D/8hWRyUF0FZl9tlNS4BvDEh0ys+gt
+22X77S642IB95GJlatncTGsB4GxJ39kXlQYthhbK2oPcWmQNrsCGi6hruKlMOx68zWbwALpwsld
h4LpNlDd23lxRLbgnSVNldi6Wf85oeh0y07TPq88GnTjXdoYmPV4GBWk1I3rQ3kLa1EFww33NfOY
bCFtsgwvS5Jy5r9BsKAnIEqSCQqhVBoNfFpKOHEhTY4+wl1L3dXIjx80oy0ytCNrI1p0UXBtrLWW
tb64H7SkTxCRUXSizXkQIu3O3Lz3vZBOyvEm91ammLPM1MTeDggiBfiroIKktvs5wf28G+UOewWb
oDfJTQ5ZHAmbwnwNjXJLVwwat1W+RnUMXSd0HLzDkkGqwiFWKmtbcRmtX/VpOYM0sC5WKLYG2ugR
SHOmJMhe/ubuYgy45DJuHMA1XMlO+jy9QE6tnVnFOOvOZpr974mYeQUV6pAryK9X4m846xTB3Pxv
AJrYtzgbsSlPfKyGkncFgBt6mbL8VL+Zg4y+QBGu4pvj3Q1crfTk8XMsSbassYFTJPlC7VQpk61R
iSLbhEruWWJgqb/qMujOCuiF9r7nXUlOkAYe6RNBoyvA4y4ohSRVchA3ufvSu16o+EWjBZL4vkcN
m1RpCknyhBSy+7nVb31ShbgpXoUGl2bO7o9WX2/6QSbX4vl2t14iFCqyP9JcNb5bU0KfNVuJfqdb
1tB2qtbEM1aOzCyd5gG1BdI6lnh2xtgAX5VbbmKSwak/4asYzzbPTxma9pQOcZ91G3pVFVZo47Vn
8ViKyaTtrtiaepXD2ypAgh+tfRuY9NcyGfh0jg8Okewn8osY3Hi+7CQfk995USabKmHjId4c44AS
Zhj7KPhv9vRAv3vviNXZFROS1JxupxvQHrHDzAoKOVZfhixb9r3LJobCOZSoMl8MOLvEt3YQvvod
wkXd6f+oHgo/ZfuLi1oJPhN501PG8view8a3KTO/y/KjMfYrXHhMfV/kHAD2/dX0NpOtt6pH3NBe
GwvqCx2zI1aSTmrtfJ/+11KTzrrqi/PN2dcZxu4S3tIqShsnH9RkSqnprXMglSnXQRsNZEsql6fN
opHdClV/vC3+zOHgRbJQQmVX+pZPZaCbfYzPvFgzw3AiMLLGOgr5YI4DziFlfRWD+T8vDPntoJ1j
xeScnYPjbcVbDSjR9h8RydBNtWDck5SzNbDD7Lye114bgbWEQfMwnmjUknBwNEJTyqYifpFFTv56
82CR0mUoDsOzV4xa2AOp+uX8ojMRzG7gQr0l0cbtew7U7tn1XChj0FIQMmEkc/XFqZICIlzIcWpp
9aswLDA2F+T7EIogm+geEw7csNrkv2KOAHTzaRrHggXb0bFIwTsC0sSb87ibO5BgfLGsezz4VMaI
YTyc+Az2DT8V0q9SR9FPueG2ljNalSfvuEDmAXDf0cu9W3AO0ZsPCGvhXey1fxtbXBeE36ruRxnW
zQy4181RruxWPu8JboXgYgFxKjUmRh8JbqOu5c62DOfGiQyJp0/xWjdlfUVS2CrNO0eRkokFnycB
mlB9l7RUWpLQP4dCKHa1tNtvLwzRDxrq5OhESwGtKKmnVPwQcm8ChKOPO359Y3ZiLZR3Rekwh3rn
Xmj2erfZ9ZCU+b1vvPbB4ejYe+CFqPnVhGt3ULSOpLDas6JrIxyjf/Gb7abDBUm80milNrUAkqvX
I9GnmB+Me+v68GlcvlQnq2Ztsn1iahLOMZbBimRQCoWtp5QZK5qdsQTq5i5h0tOtSlW6Aqbv16mE
cp5fe48yMw2ZJgqoayw2qbYjWo8+MgR3+4Ixa5l8ViknaogNZTcGVbvhFze1QtoOZWw9y0+kXjIS
zPZEJq/RZJVYAm1YwChQ3x7Ft8szY5AiR3KOK94OgB6YkpjTw1/zJU7JvpNPC8uN5ioV/c+Irnvb
/Jpubjc/2bWx3S6yCB/pPjRhJa3NiaH8GXhymIXt10pcSA+NNdlHt6/xFvd1Xm4C1Z6hK9DmZfIx
vcJnR2ctBKTlv2MYmD1ds/d61nXTmbQHeZ8qMqJX47wQmlgVch9ar8+v1833b29UOI09K/MRQ28G
b9UalvN00eSf1xGqmTpt1KyzWYvlsosP3v8/iU62hMe2xgC253Mlv7qirJsOsU1fwbHomzl1baX1
mS8ji4HRMSHw9yF2mKpdVcnMiifFadzomkuqTI6B7t+UFGyGnaIFgiaiH294O/J3+KjiSuiWCKH0
cb8upYy0XWn/fnqVLc98jjM59thpH01z7g43BhkZ2gpCKEzs44zgk1cNxHNKiE20fEtWT1uDdfpa
6n/l3EP6iRg3PUhD/r7Zhcs+vD75gJC+lBFnTbR0eu0gcngvelYggml7Q45JVYZxNEie/8FIAFO4
IZzczCorhdqQ7Nf8wFIm+adb7H2aArmCwJYFMZGxm7H+gQdd7c7JxbZhFX97hgVngQxbcLEGoyrJ
RE+lFVFPpOYueuHWlrAJ/6CytDzH4F1V+obDLWx9rCQ1AFaxmldeG2KpdzljVDOMFl1ASRkSRj/H
bziKItA9tNtsGxTccxbGhhvTuyyF00urZJ90qPqB+7+uOo/fUhLn8Hax9JFmR5tIi+WykUHHcCJb
tiAMqsX7WPqdPR9bjpz6PEGjXowV35o88Mfn3uExI12JxzciHZWWHLfRQ6Q5PngucwdEN9qFFp4n
AoCAfG2CsXl506l0pC7rIEkxp3idUQKq4amre0o9BwgwIRN/quy3bzRVpsxm6zAPn+2JvfZc6g3H
oFQwT0sWoqylZnEYjgY/jt/N2au4trjY3nbe5U6kdc+VN52M6L9Ob2aJgADcS+I+gDdRf30OAG4X
P2Ni5/4eLfVwA9B7V4j0E+Ado1Ckjp3jE6W/Gf4eBs9nJpK6WY+hRmgA5lhhhk3YNEjXRPIdJrkE
wvJsc5g9TUrZSZp7kdldTzvpHefVMqv6LHj9nuwW7M6HhXzv+MPtbUMj4qaBnOKMDg6i3bp6ITvs
/QzZx4BjXNO8ClLzk24yrYPVq/Klfboic9QmGKbyc/y2vhzvGS2X98jlZvCIvO5oDQ2AOAEr9n6l
Vlo5C6q8/033ASKpyHi54/zZaEmJ2k+aXtxuFlQy+qZUWzd/LrqnGYz/NTc4oyTF1Kc3xu9sKGAg
SOJnSovzkgrlt/0O+CkjInW4qXVHrC3+QMbJRtGv4gGglmWLVB0+RWE4DmENPohWsBKO30XNLUBX
S/R8ult8s2mWeb17ax0nXee1S00OXs4axkHsJEmZ03hs3lx6wk80v2KZuoP8Qs1uPlWRplun2uSe
qG3YNK7cFPNCVTCRGEMGhjP6RgfMMoiFrzJ1sdrZMEs5wmXLZinBH27STpwIs4oscX5nyVB2kq+D
9kTuqxeWkvdCDygX6M6GfbD5/NPTB/8RHLw6ISq8GgcQOjzGCA9WoysF1XwG9Ajb+n+sMCXp9YPy
NZtb4Fr8eMaCjYVlHO3C0FUGcdi8sWH34n72v4qYRdnSJElg1OrwzPw0Amo91d81DVTqkfRRG14N
WD7mIgABpfHu7XWR24pGswUyDaIF/WXZDui0WPWhmTo7C+plMnTs2qU2++UBUd+xEBTXBGPH1Qua
jlrjPfw4XTVqIDFncYl7fGoQ0pFM1wJSlNsIW/AEsjc/sC3CkAdwm77cahrAIk0I9hWBPzfvY9aB
0QKD527VhNi2vwrkrogvfBcKKFYDDQjCHjDpTV1l5zMvbds693HHGfN0SipV1QmkuS/uuPgm71P+
v+mcSxMVEeALCutgiyEILG/brvc2JpSvItrARfug/Q2au6xE0SLmh5uPTCibzcublBXz8/io+ELa
mFR9m434cHuwbpwSq6NyklPKOlROBVheEa9/F9S7Yl7yNP+5UKIryHrlp2EHtx2jwrJWrqHqKVEG
QOsgRXf+rayUWBFdVO4DZ8E49OPCeu1PIHcUtA9ks4s8IOniRsX4166HRagneclkSBMXsfls2y67
sU7iy278AVmTPZ6iI3LoNrP8ZWDlmocklG4MFGSqOqBlQ3/ctJorEu3gcq8YP6JJay1uDMVbVjmS
m1TiIzjbqQvmFVGoP30Z62NazoY+5nyqC0LN9Y3HgLore2OUfQusX8M/UfKERPpuRfKoBzQpCR0q
49q4Ngo5jXW5btHpBVsmQ0mvb30qF/t8l5h3MLOq1BOBJAF2UagHxNYlVQ706lFO6vSqt5w4Jw8E
t0uW2TiVAT6jZ3fCMr6UZuGMOXtLoEnNFJIuczzVyQ8Upb2T1V/piK0tfWP3MMcdKfMr9yodirrB
lri/tOGNRPt0nx7LorPAarm5BDfy+Slg/9Sm+LUBEX3w2ADhEWqvsKSvq55k+a4CyTfyChw8zIuf
cZWrOKl272RRbsFJwDS3IhMMO2pGGXYxPt2pVxpQdUCz1DOV1ql2JnN613jtaEJtCrieazWOlb96
7yxlztSQ3tCDOIYrAbf9WGC1Aa17lV2YL7aZp7dleHP1/nq1bKlx40GXlLejno5bDHo5/lFlhJH5
IZuGeZ+gd+DqYr0lqOOJ/R2c6aoevxU5gGw2oSwXVKw8iJM8l5uP7mZwRwhIhIA+gvFLZyO4igy5
mXMqVKSuKsscLdk0fNz+YKskWZAGHC2WwGaoPF8ojw3QVbpEYuBZbiZb0s7buDmVVcPXCMuPnjVL
drTxGpdvO0LKuA/8Z47ott+ZuGOub5TafSXZVE7p1qr5mOCZevX3NSQ5GMgzI1zzBCHr13ZTcuVW
svLOlwnBVO3uFTvjOq/53YPqG/jD3Y7MlB127wHdXWrCuDvsT1h7+Vchbtq13++rTIl1FrhRThcF
tCl0K4+VG1ly1D+Z6r6rCC7eaEpS2ZVFBPZGNJV/Gpdj3Us4hbCUd4gOrxx9tBC3TLKLMwl8x5oV
P+amLjkBCYPHcsreO5TPrLNy7Zb2JDUlTlZp5RBf9rdt3vNB0WEeh6U1rph3SOCL7hcMDd2k4io=
`protect end_protected

