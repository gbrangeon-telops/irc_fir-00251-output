

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
esuuckrrKLBFMMgSrVud2ZnB0pvEqrOMx6GkXz4dnPp4yshTD6+Y2glVVVlxat4oj6oLNAI0JrQK
DY/z82hivg==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
d/1Syr0Yfz0kK4aSXCIN7lq+kUu10RASco8trwm0ImfJURxtGkX5KSPC9Owus8m9ZNLVa+4W1mNi
DPA1z5v28araMT+WQkx+2smTTBb95QnM1r7IY8WLJwhz/4br130YtPfh6ALhwuPZLGS7lh5+ZNqa
WUkp+2aPy+o7nP5Neek=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
EghETPBi398ucn66loN/344Jtlwrx7OhFAMdZLO3Gvsf81gd+y/lO92JbZIwpE5sZICUxsNH54dw
q7y/XtZVcW81UXDzCet7Fnd81N7WGIqo0pJecDfSTWB8jEEqdLB/p9QS5cVBozkWw9ZXd157NWH2
fYI6wtb4DiMK+3xbswRz9tjt4QpCCW6pl02xp3h0AjoDyHQfQiHlsbTSjlklPmKa/t4Bvl+J2OsC
lbC5D/MuvEAoTUQ7SK30lNJDTITWXb0RGcdN8tf/1AbxeMFGNs+DvhkJcoBe11Q4yCS9vXGZYmJD
ooCuGIJ149GuhA9Ebc3S+zqtQIqgB+Ip/rSAVg==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
XB7G1kS71wIOs+JCFd2Cvu1TIPgCW+AVgVRokt3aIVEjyzOaNQpUv0JxfFRbYs7j+wNszYGSy/VO
ucUpEKb3V/Eh6Je+1SiQK8VPkEGyi6kMKodRtbbO1t51Edv2l3Df96scmfDCuwUmCLxAYCnMI34o
GJA4Te4oMZLzNzksU0M=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
mYbz74Wd6t4yNkXqEEqIyqTMYr1gDkxJuJW5Rg5GXWUomZKn1t4qMArQDnPwJx4y9XZOu6/MtCnL
fPfEaeJGNkk3xubUfcA48NrBjUlfoqpqaC5sVaDR10h1kTeB38B7pV1iwRz53qngpcQ/++tRqM1Q
t9nxWednDhGT13iznArEKq20RLCcpL20e+RRoIbTe3wwmYnDWI+ysKyhOx1k2FPgh9jb+4RZZgn7
7PDivXP/gbNxEf8PXBmODTX7OG6mMJYh9DN9gjuP32wcsw58ZKTKhK7ryO26lHYq65/5CZ6bVTRf
+77RaLVhpZ+Bo23bR+0rH2ulVAt4vAhPt51hRA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 26704)
`protect data_block
0YMnjLtWspbgqHB8Ab6jPPsqMytuUmefgVZU1RUWGtD/ZhyfnWQ+6duVP2DdoYSSwlGOfLhS41/9
3vWjdG7lTVvY/RdhB7bZebr+Yn1pw6zNhBwq/CfEGZMAtTjXODx/nERI3fyIXDHmpy+9C99PairQ
dqH1PGlz9q1uDMckCOno3qs6Mo/J0kCpkgg6ywqbG3KhrCRC/y4o4iFM73awsjOdksW79pVT+Mt5
1qxIbGcjHZc6zi8UePSyOtDwVfHzbchdgRh6BjTJLIagbCfqtl+5qLwKcQ+0n3I22pOhVThXQl5q
lCBM8uNpABy1aSJIcpHtOyJJkhePh0AV2Udjku8TzD+RIzWCVgTgZ46LsQsf7y236H0S3tKdaDLT
KRTh68sjMBeXxSnBMAEANhG7TYHY6YNlGDvPIW9j9kSktjzDWOnMPgYqC5Rtvo0hFe70bVlr4SOM
Dflb0VPGwYrl96pMBXHWOEdSdj9ZQ7VGeqMV7GifiJ0o9ZhbkVWD+sP9b5MMEQDn70h+kKAWi88g
iWmZz5t4jeSst6Z7J3/Bd2pLEs+Nm1eLHUdPJHNYbgpkfXEofGifeNjhWoUI0FymRdBQNaXRcCWh
n/H2hdqHehepd9+m9FinfjN3BSqktfyN4kWqiIebJfnWg7mT70UYshjKTVJriI1Q0grGqWV/UauN
p/edjPXbttDsjlkujw08FqJ9ipwaA8DxTmr5dHtA+UC7mM6a16x3tPFZ7d26GabLZkEImV0dEaJ0
KBrHpPjAbHCvlA0acCziwwMysPWavnFXJe8SRaX6SgP8Gx3WrfX5urMHUhIqVSIe1Ct5rjzhafXZ
EftROvZR8hy9ubKvAac3D73ZVM2C2y755PeVZE4/aYrp7jmSD2ZmvEdN+7kizSvrEYma9wZNNITo
unfJcc63MY9f1yjYIdgF0WS1lCpf2VORJbloycQfYOqgPNOj4EgEe200yoFCWU6UVr2SccENAARJ
Ik8LEv1P6msRw0WNk2MzLHX9Ezr5bgv/z73E2u3oHWgDVDL1yHGrculdToQqD0aWj/53SvnAtYYZ
NGXvuKqrMgsmi5av6Q2fkELODOw2oFWhN+mQamzhLd5adCnR537LXZFwhwhdXfV2aGvg8iEbUABv
V55WFSp3K3bxEV3bDONmd2ZhE7eRbGr0iimVicNcMTzJLbbcwH14RKZth/OrvRzgfDhEe0Q5CxTA
ftvwmKXtpOQM3ZtUyv8kYu+lXdTic4/kE/Qpuc9cCo6Ejptvt0e9JDf/8oSvkAdC84kbtzM+MHDd
z1iROdZiE6wSAQx3QoMrE3MFQu6QtZVHUOIQNb4kjVfiDDhrRdFSDAWO/iCtyJjoalWrZ5fC/pf2
Yto1jdQXEcQaLW9NKT71nDTVDaJsIEpM2TMxsa468Qc2exuMoVg3u92YUwsoLGhsLfCnRrdRtzoU
9VZDDneKQAkPODYCZqyXS3mQC/VaZfJrSB3cNGHMk+92VcupAoD0v2Y8rDGiRixgEqf8aaxomrB0
GIGmhzSubDal10yApkSDk2+cb8FNCMXYf6gF8rfusUIUFnE2KOGZBT4AEkrNt3h068t272ssM89Y
AUdAT2qUVUTTHXcHtWyfRT29NNQeGe0GvGQ3DekByG/iepnPaRCsPse4Bd/gq47EC8vJzYQYrnpI
DahCs943cXj0fuv9BJIjMy4vqG2/MwkGvv00Q4o87cp/i6PSOxHVgmdgHQ6VtML9vi20v5eWxUos
mFr6M7VNamCocunjZxm5XGrO4S+K82TQGI0N1bthVvu0snG0wohdPn/47HJBbRsPm6cRjs3eKltN
03FaeHNhjYr6dL0triV/uOUpWyH5POVszY5fPtXj/cdvl6/c1WnWOwGTlVF1ZecebADxXl9AoGle
nF1wnAZF43NLRecawFdrkl5b656DI2G+4KMV99bLFpcCdceBm6jU77tWba7NL3sM0F58s2WkU06Z
fV+KeCv9K0Q2qgXjZjzMEQcZhKDoJzeuTQsxLmeVboIFRyLUbk86mc+uRClVtai/A42vLEXC4WFy
729bxeayFxlJUn8PXARxgFXJTfem+nY527W/jqS1QVj7wnW132D32v08MVXXok2T1Ny6owJpcPMG
WGUnWktG7GQ5JWM6K3TyXwrzGt4RGttMgeqdac5NWqhJN15tYCveZiu4JnQwSjkr9AgylUgyN+6C
HKq4Mus0P/M+3I5qzJdcxpR/6CM3ObUw5zXSX5P/PD+V96xhkGOOuYyqef2/VsrVhF8duaVDZl6I
Q5mjBD8YKpZEZBv/eUCI8V+Qf8zSH7lQS2fDQfayd1jOvBvnsvZkucLhDlgrggdqDVhG6RJDkdZ6
i2k6hqlQA5WZ4bR9UK/bsiL4TpH9zPJujulg9e5FIqe64fwP+K8gSAI+eJTglIcWXuey0gvw7tNb
59p+jjGWc70fLlwWQ33Xitqrv/Nk70B8+gBKj8/oAFPGlo0ySOfZ9mAMqXZfTg095a1hN3fUf1BA
YfJ3WIMQtRXRnuOFB7cxrezadnzfXtrW8l/PZQrcsbBkASZpJnL6iwMmVqlrCfho5Oz3Ywsgd3OZ
VCbFdhCGwUxVWxT/MFBOFZNjrNbRl2nYzWED6jCkRZwhFpnGsgI0b0vEMv8x8XL+dVCai9GJpQBB
QzFSQoABfdGyDydV1ByOV2Zfshw4Q5+0niuUEiBje/flYD582l4hTKTvzzSa+4nLjP7tFxshbPki
NSF1jmHIe2vbeRQkfubrotZDZLOiv9VBs+nMoLJA0V5kC+ADhBO/D0ioGwTovDq40plmajbQn9I5
SBovNzW9hCeGM3jihrIvU8tySgzq0DYBwG2MPlx06HskTCWq+EIjtLknoex0XRk7QCD/xZa188kO
gaqDqcDU+WJ3Xvo4XhCfabv4k2XPPZLX/vq4kxctg9dOxAOUkoLVUtN9brB5KDiuTrirW4AIKZAs
4N6HwbtXmEBE7VD2Uyq4BPQZrdCwBpXw3ecHPOEImD/X7QNjEVMtubjvOwAdRNxBRt68qrCNMscp
RasTu8LJTWuwDUhUVZk181ncSyd60zCFZUfcx8O4A763eG6ietzhdl7tfArFZWR9rqwiC9pZ694B
UEKkblTV5K69e5le1SHm/8BMfqmRgJAFeDLxJrEjxuHgxFCVb4fIQQsDOsvz11tkUUtPSzSHORBt
NQV3la/xBYdtbcotbqVtmOcxF/uxacfoXdoxbAjaOXgpcKoFyT7A9VGxBP3Kaz/1SyXLxEJUBqMF
Izx7CwFizfFcq0mbca4WJBKjtBRmHMk9pulm13RgNfyj0CHBJQHV1k2pm1t8CpGoYIgGOThHM1Ba
HhhgqdnODsL2GLnWTuRMBLy0hVUjyCxBrJkPqBzIWhdNUxpcRWBCv0rTk8xD/sNsEpGceevkeI7J
EtEMpML6/dZQaO/bcoolEQwLRX8sr0RrVMd8Zxgmh9+gCfa+kFu/uxdhQryBkydsGB4VMEWFyRq2
JiZQmSLq1wwzxLSDg2N1mGpCqCIgUT++B71a9grfnOqLNVJb45B01Vb/lXW8p5qIJNfJgH9Dn/RZ
tqN+2RVYfUXPVR7qEdg1IFbmNA3sgBjMUbxND7cu8KuUqNz7tqY+2gqQY6K8drsb3RcFgx2YTdNl
VSAGc4Ts+krRaXwXj3IeM8++sU8itpsmV7TILHOL2KbVObETrdVhfXeTyVHxjcfH19xEZZ5V2uEw
YnYYOH4/kv15bJwK7NY+DNsAerAuxfKtiQpGZkKY4Ua84j6RgaFpg7y79qw032OlOyEthhOQkxzF
c0aCwRFCB6SC6usOshUJGaSqvvqtYOuwZtKvkJGX3LV23UmH5SIn5gZHEwphBa4JaGy3cLtqDrQd
I3P++mkK0I5E4vNMV7ly68EMm6gPDFibOOWQjUwnQ7B/T10dqXXn44G962aqE4zGqEAKHKmmCq+a
Thvn9OB9qja1VwOwgTzVjvcRAqqCphuMO6Pn84VkbyqOguUXgZbRb+hO1geXgsJptLNECTEpRa7D
XdaWuazVXDXGEUbIdsS/BXAhd26mUqalhXbnKpKu0Vw6LZhtxh+DrnGcwGGTZ9umwwfhi7GdbxFl
3ZFLRqPTBLKRzhslTirfNSipfSbS/EExRoXyUfwUUHIvBtvb7IdZgV2LqnlPLVawGaCalTBLnwds
x+6bkj2T09s0VKxtQhGfYkQd/Lqebi43VijJl28Lamxo1wIBCQfZG4d9SO2okIGnZbYTPc6Yifer
vlVB6PBx0iPCusFPJ0ir+79cq7xhvkjzq6jAOWeGPI25bglYFIiAhGHJsBR7gjh5O7IVbZH9drNg
px6StlY3qn1u/FKxRk/E0fcttBopkzvQCQcSD2T58rtHRBxMTep0A0JdVodmkBJlkG5ZkQIaGA5j
6nLaIeonc/XsxlnHbMne4Q7KgEF8u3tuESdsUXOWUxQw68rlvwqqFRp+xWuHu8bJ1yzA2UcooUgT
pTSvUqMDb4B2HbsYbZxv7ux5k5XAAAre+JZ0OUTCuXXp0Dk3RNIjzKx2+7YuQt56ZFdjgEN9DNgu
thcMw6QfwTsm37yqXnuvVjgMn7kwXqZzWjIo2B1gHhq0di6rQQ9knssxCLEU1um3zDamidM/rzFO
kZaQQjZAteCGjMe8jqOoePKQoTr1/nYZ8dnkeHwybGVMztj5F0xZko+u7ivo140cJ6czlGgFp0lu
i1MVsW2DTCAK/TzgWgtRpAYUvi88Omu9W8tD1UjmUVmkaySRUHDZUc9HQPtgXq2GFQjev0RObEfG
KRo36XzXc4WrpJxjUGeQvPCX/3tZ2NHuPHoOeU7aA+iCvk4F2zjlqCswoD61Un0D7fuj2rA7GcQ9
yBCy82ib/rRO1v9ZfpWF9NfNIEcdIQ2Hfcv0phV79PO1/WpZMjMlTKzzNfhS3xEQkgM1Tp1ZrMGD
fOVORZUXbLkf7dPJ8iGTaUNS1jthNbobCw5sr1ICO+zpJpZqZ44sFu9nCk42oGbZIkr5yPyQE2KW
izSsVRbiRj3wRdzW+OYp4gfqvBLYrlAhxQE8MQ5C2von+TJasZLryBqx2RhCRnQ8vUXfv0xmW8Ma
rbSY08eJ875ytAjPKAxex1t4zY0f8UmBPQ/+N4HR/sXihuQgdK22XM5lZCuoI/8UEk/BQpjt1M16
7hp7Un0OZWgQBwCNjt9mOczQah6Se2cuGlS8x0GqgLxSsFHX53PH5t/nPneVMOLzuFNsp4Glbnzj
njxQD8wSE3Y4EgvLNjQ8jmMIEsN7YZfjQTu3RvhmLw14C3ZTZNudiNsHZAlVTJTxbG6NUnE4ZQDf
RB0hB5Dsk7/fNC0P0/X/QEvZ0ymNA04vwFuz7vRQaPHLPLkU9EGjDSoHcdgDPwnsbvfmIEVfKh3y
9bxye9R0iXi1uyw4/M6yYDxOAOQL61EJNPmUM+ru5nkV467lofEgparrUmz3bz8FT1m1YG93TTBp
zXKzB0aZ0b05fh+ELpxfTq5zfkKyGp+G6+g/+EFKdZvgLjWmsnLZIINai/8brgz7803sl5ulu1RX
GMiLp8tqq07w1oXKPzesIgRP4qy8YftXW3MeWFFKsKbi75UlEEdKhQUNtuT9s+sYaKpTztw/beHl
qv2ZGpIV9U4VAXdlipvsaAyUfDt2Vm1YRE0kk2YntNAZ8u2/w0aUI5UktCpkaz6u6UGZt3qwTraf
shvx6BlmL9w1MqiLNwNLYCPNdstBF1e3OLTy/KsSeS080dXe1pI/kT3LYds8pfsul/sbILJ/c50Y
kRSsd5zPKeHU7ndKZEK6myciFWRvue2gZM5jBegCrAralAwf6FkpZTkr7dmtrlf3KMYGyIiZanJ4
b9bjSh2wouDKsSaoQaJ2fr7gcpCquE5RdcKGbwdNstS1i73G/gFfnq6z3jxL4ZbCEcvlb3gLV9rp
7SFAr2YHbqbeDTzH4E52f7M9NjAEWWrp2saO1io9K5ibGrZG2jxg7zZh2jB04IW6U7mJOyVMvgkU
DyRCSry3mto1+dbaDYH7lfpMy9fcVLTBc6rnHK7e70wGBA+oPVT4osMnHInpNKQzvxhnGqbPwefv
2qoWBwdLJtxt+bfhwSKvl84PVI4SZlEshqtnJvDEqOq1xpeTlW3KEeGP/NpmNFXsTOhobcXe/L+C
zVeHxj7yU/ZYxQce/T+qg9VHDjftOwgo+ARwYe/Lx/LuJWnggqqzQp0gJd2xRU20v05B6f6Reboh
bb6SFwYsvlMMOR063eMnrcwbXtZW0sMvPw8VmWDFc/RE4e3Ywy251ceFqODFE939w+xpmsL5c8q6
Dc7FAMeRqHuJyaYM3AVA+vAMp1EEqH/H6NSSfh3m+Zjf5sgKjZQN+od+YhtWKYQcnsQN1+iMz/jY
PUtFwXYUeRaKf3J0MqqoHpjm6s6x+eaLJRvMdiwdLrMG5YgRNjYH1Et6DF/4oYUAngPAolLVa6c/
Myt/CHlkpbSfmFTO2N/lJqjYSEIpC/inb6vkdxB9ebT7erqoAMO63S4gMWgtDP/zdq/vhEyVmB4/
Q3LUjB9Hjc62THiIEupc74e9cXTykW0t5H+UgwuH4qIhPoy0wGt0iP9eYdsQhlZAmkafTE5Vqs9k
rrVbf9dm6R0u3OQmBRuhYjreVt/cJRPvXrG+5G+0Jvp8CWhRZRQznZBAgcCJUP+Ebx0mWFU2JGNd
n9FJZXwNIV5EKHQifgzBieyoSvC1IWsMNI1/dXJ+zq+MNibve+eHxmB8BpAsx7O+vp1Ig3/LMJpU
fwPcDC2ynaZCfTU2nV8yYsehl5iY8+aUTrHoO3cjUgI4Zk/dfNYgK87y6sDSWJKrC3QtyHWbA/iv
s+alxiFAsfOeOjtiU6dK45mQjIlh2oMUmfKp/C4uZML3zFKd7jpijMrB2mx75O0SL+N5tDGWwXnR
HwlB9c0dgw4u7IPgJIbaJ7zdkLRQROq2ZqKP8487H0EXW1h5ncnUvJERt8jwrX1Tv4sbsYrNeoCZ
LS80U+5HrAbQxAKzbMOWsDLarGtWZD508TqIz4bcPL8k1TDsSD+ee3aYhStuEP27VRd+TlSQq5Vc
zFT7QdRqPm24N8bmJ1XMss3aiCZ9prbjc/0aeEC7AIpVJs3pMCOBaR0moiV3+OEV7hyBvkS8vyqV
PEm8vfBsJqsQ9NEbytDo9AIqlBODYW4TQxzMbiUDJZDs+E5YLUcGstujt73i7AEO988Mjdpl7I7i
h1VoQWiVX0l/u4FT7oDdArWvn9x0kKhg3cLUmZdhCKubvQqi7SjzGzlQij+xETOBUwqjQtyU8zM7
AJI1N0/gP9dRMcDKxm8xu8CclA/PwTnTPX/6nEbPYu5nwm/63DIzoYONRYmvrgHNgTaI4jtl2Ywb
M6xoo6su/RZP7Ev6gD83R8zwb7NgT/Nl60cU3oTLYfAB7+riKcmAFpDY4MEHE258OWpO2wFQPEZ+
yGQHRew4GfXg9+5f/mzV1SEzrSiqIhMiquGJqfDnn4M7bKXvfwhguRO3MlAn7ash+vuOlGQ3DJWb
AuqM5GlbNTuhRZWlnXGbNqAuLqSULvGmJAGgH3vJGVOn+Om6a2mOIbgM9LYpF/E78odc3EPKzIBk
3kvZBYW9xctCxFkX+FX45kS5Or9WeSutgJOOlmsJSuHQv6KXnpgWnsJKsVIy8/CakT8yk+wThn0U
h6LH1cCadyy3G2luj+qeyC2joGVpNlfyTBdHFKvcnB8s5f11hPumAUBfYb11O4UZpZNF7M3xUC/c
TjUfE8ArS3rGSZDaiMm+BJ2iFIcooKwBz9R92XQjtbr1FKjffnxIK04NBvzyXfLfGTpWC+5f49b+
gWtzfVt5j4TY8UstrN7Yoe8DXOG9yaWzW9v67Z2FxhtEQUYX+vz+1SxyurFpasm2QV/ZRs5BJAG7
c6WoMWMXx7lvIKfk8SQXKVZlQK26yXQztVPOISoF4Yy/fIkePoekCu5TEnM7mBN6LMidJsld1pC6
O5QQx5wLAR/31INfjxXtRmXoVlv3/cr5tAkzr06iH3FlWHvk666pehEQ2Ydmavs2H5N+KiK0/WpA
4moD0Fax1RjR1IPKfKpqEoTk/sLIP7zxPAjtvhn61kdjh5JUnTQHT6K1bd4DfKzw0LWABv48AmP+
jDtHN5zNnw1/TgtyrHrjf16ApzuTDDzQpPE+gK53VSpZRLcBANW6oZ36U6Xz7p5lk3ZYgvXgXBKS
WN0LpU2JjYemwCGbGWREp21NQXaOUhcLBQLwEL6ayi5qcmB+4LMo2KOXJPkFFAZ4q6xh+ljLhVWP
pR9Sg9LYsY+DswjusxyBk7upKdu5ZRt7H8zQEBbgv8U99dcWdprk8ZsBqHl+5Lx8bhPl/ejEcDYi
V1mDBtquoRXyj9aJmkeNWZuMcFbazNkCXQZgos8SHpLTjxLrngTbTW6rODI+A0BTCushFsD/37Yp
P3eoL8PHUPhN2oESliRevG5lHoM0j3DWBNWd1y8NQ/AlnOXhrIh8uu37fNjY3Ck8mqVbmODleKd8
Sjn+9o6sAcg7UurGSNCNA7+6ClM06nOLMR0H8w+RG09aXSxb7+bDH1nFChuOfPP3/1a/gMm4jFBl
UPdZImzMriXWlBk8+mpgAzNzpkD4Gu5xxeFiWRSRzXFTrS1+pgzd1aTrX2nnZE9p+jzd9JtCyrI6
F9iOcpGTgh1N6nyD+ht4mgbe1p9yHttHBD5AUDnaawduwFXt1yYkyvZFxPCUhuf5mTUsJPU0pPSJ
32zDhT7D4WsNpkRWoxCLC/G8CmBqXLvXdTunm6ax6W6p1PBCEF++115dqMlZ3sMWb6biBHl1xw3e
VAKUbsmAP3DUbNXG+tSx80eO15MMF/h0Gbq423LDJP+NgGAcYHRm24ypmM/hhZ0lBdGuDbVDwI9a
aAG9KmbQC8GPLwdbN2olP3NJ7BiWpyCqRWNn95AU6xG0HqOex3i6DxggZSrzqwV5RDM6olQSra+i
CDqbzy5nR5insn54lrisdxGxwy/ewMpsHy+1TVCX99IyUGpE3LSLAwkNHtmpa4J3nnYJPAeOGP+U
IcWDST12y6XLnSaGGpKq6PrlqQczYedJWk+6eXKKaLmnfgLiEbBudHy20BxG+TCK2E7XVNQYXUIH
Y6TwqaXkUqrXcSh/QOGYSOrm8IHPE39BoHZM3uyR8Hy5JNZja+4JaiimBShknZ/0nC+sG9VgbfJ8
GSv0SeE9jQAILvVzenT9WyOWNzTTenV7h6kceMynIxblnzgAQjC67ACSGnqzOX3QUtP6zshXcXNQ
LVcCTREj40D3GdfLRg4iMCC/T1NU8vP8Ixt6hE3Xbffi0l5XS5bFOxrbFn1H9+cBV0m8pd+dPzpo
2KyjWZIyG9jLha0iYImjqW1b7xb5NDZfCkoAXvGwjLbq2+5t9CshW/xalxfA/rPU5H6nEoN7uFJo
0w3rZ0SuII7LkVQX/yR897iZ7Vl8/vwKCAzKR420OEA7h1ph73rHxo4tDkPWDtltGky1JfKuikAB
Wopa6/H6FiirHHq/hkUMQQxVjqJXfejGblDjFtG/PYK4qAw/ywv1+o1Vol2Og2hYrJsiVfkFja0l
TtQxCwPmfUZapJL7dlrMtmi4NNwL9kdqs4vmOn99XRIky6E7NH9PCXW9oKB9+rkirDyIlzKg/Q22
XSZXm7FADX48dYqaA4PkolZeKpZICTqIH05xbfuD+RQOCzklKwjbB0F3sC79vN9TXz8MlNE8qP9L
7jjpOM0fDqH7ZmTi5OlqMMhQL3q1t8AmrjJIacZcG3hHzCjcOiH3v+A1VtmRSrFDM4a2OxqcbNfb
QLCk77e85TBn2D4c2ERb5S1MRaJB6LEMOOpJ0wEUbY5Y0vgLer8ZwNkJKxMhq1XQ77S98S6jtOeN
UPK6+GNHu1k0TlvIVH9vdoxa4sSbslQ6ArBHQ0Ls5YNeQjYRexVaQVBz8B1S7FzqO65VfeKuiJ1s
1a84dMnrFR8NXmflW3QaChoVNdSisjnmbBFlfvhBDn4kqjrlo9d7gzu2Bcv1X5ZLNObLXY/Pid0i
+vnIaHcchrf5TjPeeLUHiADTpN8sJQZ7Kaed0raPFbe+mJGPJ+C9RXypz7QJUpdYgzWsYrb4T0ks
KSN2u3/IWCVF7xaP3eBMmUPDQOEgQFjeNDSZ19SPFuR4OSDC/NNMtpcGLui1UQ8G6h6F1DswAOrg
4p6nElwKEGsyKh0/O/nxr/203Jm1rqaGbCUBbQT7NI+GZyVH0mC3VUUpLZBOyxXN+6ETRV6yB8uY
4kN7VGIqPGd0hggj3Q84Zs6Vph2yEGtN/678kMeg6ipcn0Q0pQlDv/d/jXMDz89he/1BRGP/SFfo
RucYgwSUeckl6LfcYqQEqtrKaxL0y1Ta92+jC4yfPqDyQpW1rd77o1phJRq1M9L8NFE5+kOxSYEs
Msxyj2Q66qX+DnExBFQpUUHtGJBmn9ZUTU2Bz/pONereBa+Uwu+1n24XoMaeEqeWbjHzpyVf7z4V
EejhH0spFvmmMu6/hm9RMAWlZXBwyp2f2OFz5icWslqh444isROHXuUh3LijXPG413TSyqkiMdTa
Ky27pwFuW/ngZoPoGVfRndhutXSBd4VPFWAz0k21K+2VOa+wF27/1TbCtpDaSMs+7FghcwAJNU0x
gJAvzUuaRkqAzd32jEm/FMrByI0hXeAzKOWfugZqF8xIiNa+lDZScynfXQnAxPF/forNaB17TjKO
eKpPO9OEpnZgsbupg64I71lJ9jW8RHgSVq3D7Ks9ps/U7aX9Uv4juRiXn0kbcn4Jny6Xz8y+xOk7
w8XmMiAizbZL3Qv0We25Xtu7sMfloVjjT1Bieiphf00tQa8S6se1+zidntw80fM4VDXxYjWuMVhR
NeRrl4vy4EWOYOWiX/IvdPsmizBW72j1dm+Gftmfu7WU56GGCgfTDf3Ng+vDyz4zFXd/PcxoNveN
kJSADXSNxhR00T0V7TxqL1NdUfDowymamHp3goeDMAuvqeZIN8NrsilWxcE6OIX+1oK3KmPLgv8V
3VRYXsGIOXDmCqLjOi1ckvSo/Xyhsag5tzZHDIn4I2PRX90HQ6GD2w5Nee9IxKJTjO+l2BZgZIaI
ebi/B/WVN5LiEQe1P46ZttJMl1clhRzhO2XH8plAtSNZWYBNS109Tp5VhyotSueWZ76oE9yZXXam
hKPgmYmqFStsu6DXXINvjCyTc9PF24qLhTk8qXSPAMpHo0p2vGT+jBZQic7wdAg4g7o9OXsRRyin
RI2P45FjEcqdbGKrVGsI64LDmzJO8F5qqRcPEBEqgTSAWWjQTUsb8KxDVUfdfX/Pa1MAjsoNUqiR
C5E5b+5xrM7eU+/LGmSrv3dxF8rDHtRDhc2wrV2rs96dAqgrGcMkhBIgLqawtgebiU8Wi9ACu7YO
gFS9dYBUzZp7e82OVlSlJ4ZHyyGG3nyEMduSCTx7OiLAdGeamApVXu63qz10ZyNtH9D0NzJAdErx
V5Bt7/b17Im2TFTRyZlaYfl2iCmttdn9XxQFy09+7N8QS0O1kurUHH3kIsYBrOV2wee6LSVsFZ8Z
j4QJjJCiyqGaSrXiAvF2oc4nbZiahpPJBnYk3FqvoFiqFyJu8Ruvg/k/2AcQrQNgoyUv8K2dYExM
tIzUNGTYtOxDcmFBlESRD92S8gL0Uqh+A8wVIAJqtfH1qfLZm6pGQQUm8m6tVy/SJm6c7NGh3bfG
PhfwaBfhoEyom366kIPqEE8tWFM+DOwqpAf1Y2WNYxONfQhmVy7bWXIaN51A/fL1f6pIyx8EZDxb
hnXlPUHOd6trFWs9IqWjF1sfVhQL9YWXFKOC5v2+LQNEFMJh9ciQD08NbEiy6D1b67GpHEiRpRu3
sz9nrzq27QBDjl7UsbJgCLNsnnEykPQr24yoON8wwD9oYb5iYQ8uHByIQTzzeycvfFS/AA82Wb2S
G0Ti+nNRcWM/3V/xVdfydD5Ue7g2cBkOLosEETIdWl9v1wf3mg20/pep6/oHi85ie7vfYP3snoMB
Qy6Pme6mm1z23nouDvOZ1w5PB0YEv3Qoukog89xJA6M9CN6moaJ7Gk2gc5h+6koeI3Nxbk85Vg2q
G8p1Qj8w2lOmZN15gN1fT0Ak6oW6NxdfHZqURE42wZEJjgbQSe1q0+Z1eLXo6em/Gsgj7LpWrLrr
PowbcHa6VGvOGIEDRVe9dsFRRVj4Dlu/KrQjJvEqPw5tLI8wHxb7gpH498CYOH0dTZHrBJe2J10v
Rv/OFibxrodIr9x+IYQ5V/nR3rElf+yuiWZ+Lau/WkVm1XaIqoZiAp8YhUpqvVBPF8mkTgBksPxB
4fhl2FXMA/+/rP2wz6i5TA0iC5kRZyh3cUnW0otjbBfI61Q+d+rKUVlB/l6jX/9Bab9do+1FFnTJ
YysmtIjfdhXMnA+YhVx9+MNVUBbIojYrNAxtzeYqevE6+inovNTOA8gODjwyAjLQ/RtEd1vn3lG+
Fvl+0rKqOKVukj+VbFqmMn20+Bd7QFcDwbsDOoKkpqhMY2Yhs9rtaDMoudz0KrROQtNMd03u+p7F
WpXvclEY6X4/Vj+20fmYGzOvG2Sq0QKYoSWv0cRsNtnlcAVvI74TuGuoKbpwmn+Ke8zzPPJ8GZVN
BW1/hHGnK/lgpFh4bsSKkApXaZwAoslO3uRjUCT+wnE2iYOrVyEl0ORw6H//SBGFF5MKPP3pIhtj
EaUgYu39VAwQ9fG8nuQPq0PWJ5EzXBr21txCX+GiMhLdZyBLWmxrd0UeRqxCRJ8SlDqvPvWG2mBq
ghw5bYwMcbrPqohIa09QMhDWPqibbPFmFDzcsVWz9MLzDYOHuVo6i72LxJ52WVebMfWoY9GDfmkO
5vskjJGskf/D6X8GVnRIBqpGazPSTFLie8tooWtcNZ0WBzQ8bee5eMnriCp/4R/0NzuYG1brCioJ
5EaA0IaVIGEC1WeJK4SGjJQ0uNTobiR0JVUNqW+MtLYtOISDeaIg5o9AJ2kJwodvlFkoD5a7FwzP
hW2s8GDQuguCz2t8PIjd9uv/Z7yjQE6Sm5Fn2fpQFAKji3E0OLAqisEhdyKjGF4ZNJKk7LY672vs
mnIXH1Sd2idhQ9uYpvxEopr1Zh6AOQjOZMDe7eNq1xObv/f4JZff++I4zLm98CCMSfdtMvu2IO3g
P7PY18z9oZAjdH8hSJYalQ3zTs8hnO70mqdK6gDBY6s5BDZv6ZnWa9IuavMms9RQ6wBPxSD/LXSD
HszUVeIKhnQqJ6fSP09dguIlLn/Mc+uTbsTu1bi4S7prADyQ2krNRA5PEKymR9DMfpPzo2k1A1tU
lJcJBi56gTUhm8SAEUIdKgqllt0v5+dDPYSkbpR51bhz0QvnKm7mRtfKIue9zRwrprwuh4a+SThX
aCT70fREpDy5Ym391Ehw5OX/qJ6vdIyGjCHxfzYxgIwq7+DfUFIDjv21TO2OzVekvQe2WaQx3xdk
sFOflsjwFwPl6kXOmIBIW4ZjNXMdO1XUJALTBcsEuz7o0QHGPtL1xTPeN38aJLAOGFUxPakCXKYw
QBEtsiWfDRSWwxDYUIBaTsOo7qi301NQfTNGIcB8PH+BhQFpvuJb4uI5ofAX+EAk3e2+sARqeAIu
Do9ZTg0ER8Fl6gg+7ZYNdmxsTX5pDoXzXxGQ5v9Baodp0VRG9e+2sMAtm+EeaYNyMYIfyEavrZp6
ssQuUdY8RAABpc/D4pGYthXRWlth6xS4pzlxokvB9SsFLo/4up1qK2HV7TDMOlGyf9BnaKRLD1OE
tKU3ez+4/UgZ17ggUbIoi730a/45548ilyR5kXVpm8n2Vy5BbznDzjld0efSxHI7onSEWAvdaRQt
aLexa9N+vG0ggkh3ViKBop50A4ZwLDBbBfZSvuZ/xnHLptAKQt7aXVOxpRu97SHRsWqbAtEzGiPl
6gd313VzWX5+jen9cA9lIazSiELWVQstqiLWhyr68uaQmIBn+85hdP9xWgzFq1yp4dH4sIXTT0+o
61cfLu9gykkjnvyPOCJ/nGGOFwA9oRcLF65RJ5c2qbonrOql2zHBBGN9QPF8uKVi6f3M4rqNAGCN
ucTGMT9VedPC6tms69NhPu9tYiauDVoiKYBfH34FgvLxdVPmA7o+NRRPdxWQkMGjE0bAGpcAiYE6
mBTTkS0Cw29Qy0GEH6fFadIMkKdNnWUn7EgSEh8Z54BG0uJh9yppgKWW2qy70INZCROHqSSEpAZw
bJFIVpK3PIdE5q3qINuJdEYrv4rtyQC/KGEXz5kI7ooRoFZs9/fAsnG6PFWQPq8usDzQNQuHEioh
wLmW7vBhaktyINIr2bPOEpGIAgsBijdZOTJUD7K/njOeoI3sP/y8w8TFS4X+Xqd3CZFjNxirAt0w
q0IDxMacXsMxm9TNylQeZwVZbC+rqThYfhddgkFqoDZKFXN2AbFZ4k1fEt5T2wnANvzhFIHCfpWd
0tM0qwFjUleXo5x/WmsWae+qPQMPycOYPXqTLagkSOO+UwAO9yzJehVNTdLGw+eLoPjpfk1WrS5s
zlTWfpdhtVEBYECpTD7LavsdywKt1HCfgDmwF4BZRcHJVkT+NAAlQ3g7icNATFp4Yz5xmdNLpV7s
BBOtoY0p1zTa2L9zCUE0ThjFTQgnuhlsyt9/d1erDNKWIOP/p8Z6IsX2tnUrXboEioOX9VXn5oxJ
804Rq4XYmoFggE6SAVzcWt1t/0GD1u06GDobT5W+xmBZ0bsw6ZoGaPYYx73bNkgL1JMBABxQWXmv
zCXvlMntBSd803Y16PK8lJ93EPcDENRVJfQmxM3TFQcI1Ta5gBGvUClwnKrgqCtGHIvmdTge2OCf
/xI1OeQcQFDMUjCm+QivJKIWOpiD3gFCxii7+LY1pfYFwv7WYlgeMMTUpWmhnLkNU/nZ1audDo7v
K0qx5UziULCfq2Hf1aj0/PUdpEXZQtUK9/ct0P8s9FR/rtjG4eXmtoFbVT597Z+dl7FdSsYDgV+5
aDSzduP7PNyRfY7dlQs2SI76/nO8DtMTpQ8XsUlTvdOSs336V/onIOQ3/9gIJdsy5b3zZVWQ8Cez
bYhtETa4O0HFjyeM85b3H4GYU4d1wL1hw3PmXxMVgEGP3uiqu5mvkc25VKiJYIpefw6NQL3BbZ/M
tDMrZTEVV/D5kMjoiWD8uNDYc8/L8xyWEa/7tRMTA+qTPQ5Z2qEU7wH9b+4zFQQsYNRjWoCDycd/
zvrAOKHSDIjmPNqLBfBdShYBYUUhxQWes1IF16x8AKQLr1NElkal4gV//bkDlgTsnCYQXIiHjd+Y
r2X6MFX11zzDn+2Eyk7ngl/1tVJrIw4O4DPGmChBrwugz3IumxpdEyd41L0VYJVfwvhdM+e1vnPP
zVXDV/z9xOLl7HvMvVsa4oel47bhsAR+F/H+hLmIu+ZoFo1x1R7XPzAUNRqF7ZrVmt8/cWD8RTCC
cB8TZvoolkOixNYbIts91H1W71DNrfH1/F597Hu/cBZPoeSc+r99++qpxBgkfyuZ8tTg04VDorht
4kDN7BKp/uOrQX/liiZJSj9XfjgF0k/NeX6Aegv/OE1GmZVOO6LWJX6qPQ5oPN4PmuhThJ0hjJc9
T4JhY84lRsTYBANejSRIFINIZQRFh/NVkE0Ow9AttB56kui63YFY+zPgpCaEcd8QWo6fUQMHYVdP
BZYgi3+AWVQto4qZWr/bSd4puQLh3mJwOYgAWFG3dvBXzoaYruZ+VfD6lVxEDMqqbLTVJIkdrWYm
w/Sk3YuF5I3W+1Uj3qZGxfcWPm4d+AoM6yDYQNPNKHx++MMdKZkzUMTEa8aLS3IoL802Jh4BjIzl
pY8KuCtW0EEbVJc8SrJK7MiTpKc7QourKyt+wGdqu3F5bCg3jYtDoZWY3c/L7oQN3Tqd2zmmG8EH
VGH28HemrkX69uCOcU4xhWplJrKpMUb7M5uLX5WqwNGPZux4okS1CZ4y5rZvIYMMmzVcLnkVR/34
fpLPp2yYRi0wWcSfnMicX4mAD86FI4nFEXzBVZsauVQTHAJpSRqOe7CgFOmUAeBVzvbFAR+9woEX
1GmmFbIRPBSi837S79/Y27ZRLnVBPoRTgHus4ov3EBM8egIK0GHIbJpwGXkzBfeRBT+jwRkXjLvf
z6n4m3zVSOUZaaKCDXYV0JVCZ51HhtCL3TqSh2Lqt82RtEDznAeEuFKyjDgc132F3ab63088eeLg
I0EdpfrS2VpAHXSd2D3VkK4mdwRe+5Nq5JqWxabQhprTwGvRo/u4P3Kz16dA4pX7JqMZOtDCGWKt
xhF08PEqhsiR58qA+/f/BUimXaBgEKUr2DxUsN8v4sQL/970E7ChWb0i7xrO+6fObAKOz3m+TM0I
sQZi3xV2j0O3czcU5Umv1NNqMHqTapR+kK5Nlot8dtNY0rATgNYq6YauGz+MQkSzMAU17Wlfz+ra
HhWPCOo94SDBlOr8j8/1UCWCGULM0fxBGJMY47bkyiTA5wSNerpE1yG2N3mYcSfUCBXUctpnVJuX
7LVJ12WChDBxpwbefiOp+IzsR1IgNYLSmbAIvtBMLtJJ1zdYQKWNgfudVfo1CLMAqGwETSIurhEa
K+EhT6axx7s4mZ26YtTsvmOEJhzwSI6gNBCTAAfyqa6qSM1TpZnrw0eTHfa1S48VigQWRYkBgkgx
nSIgLwkj8r+LQ4g+4iXSp/+UHxTG6jF1EBLy44Q3zl3wCzSp6iOSA6At4Dy3ZI+SJ2a3vE+NL/vk
8Dyjwp+E8KSrMF2kwoFEeXLijj8PUGHAKdiMYJ0Jcub1XnYPglUp5HEUWxLDjghyi6b509LdsRZi
RNswpEJS3HZzVbcRtZD8hJx1y3A3kjQxh1uZS9Mg18fPK2uLqF6MFBURzYeIydU+nkzigrycx0OJ
CCa3CEmhFt6PWuQfWTdVCY9/Gsp43AFr0Pn982j1eKBfLcuJ4Ucx6T8x1jC3kGeLxsHNXOSMsRq3
3gLe92bBgq/dnh1DkI9L6UJVsqUGYiVG1mnIVt+xTr80lGMk+zpTyD41+gqwW4lWQWpTpZAZLdiF
4S/zLGwv2decJrC7T91TfeHP7en4ioD1aJWVoua150mS9n1/USrQxgdMnthZN7cKqvmdQ6P+JkFI
FIv6uzDJ8ZFsNWhUw9d+pHDgMbym1ee8UpKDmyRSxGUu4XfrUND9WfoWj5Nu8nuMVZTPRWvKCbbE
UjBqffCg9UEhv/2BCldPeKtjChyyC4Kx4v5x4tzc9QZh+jCzXAS2NySJjhAcepMLbJeSMlpnA20j
+XOBT4ElXqEQ0XScrBFrRj0gZJ6VKBKpicItwNWJVWCr6j08Hs65+TDvdMlXW77CQsEhmhQoYpm2
E5DtU8L+VjRK481rmHCOQ+rsUvITT+b8eulEkLYvsdJ0KPgC9ybnAP2oVNatyG/Bafy79XBhbR1P
fRS/4posO2J+IPNgKJfJPmtYVPFBt+YpsRqJv7TKLD7otqn2OH8aK91HaV/Dxkb3wYGRIwbtl6Eq
dNcDcQZeOhBbKaJ3OUc7U1vTubTdInGzhwJBckfTuxDplgSruOQPZykpy805iKNgnFXSOXRDIASR
pS1knlgqnqqVuj0ezQ+e4Kxbra8Ky7d5l9Ypkva4BBVD88uJe36w81obExgT4j25RCUpxfDEUPvL
pNEO31qdUE3KPMWlqbYdwHLtv5cD5y9ZvyBSgdbhi/XbqL8Pwaox3+pKRZKdMp7iBDQFcMleHObm
d844t8KVio/FCgkLvAkaPMSGSzqxA+8NtvxjROH5/RE63tIBUn9TCyckKoQJv3Cr5IgzRnXBCEpO
t5iEXQhzCQvDcZW3psyVCEz55wwXkJUahYl54CfEltvzc8ThWzUWAIuO6m+qcxlEasIP7kf5rNHe
MgJA9HtB0nELHfro3Mjh3EU95XvFuZpBBlKjcwa7xkdDbIsf8eaSspQuHgho6/oqxsydE3dLa8wn
Y9MoabpwmfQx2SxQjWPmtngLn/l87aeCyHWIcWEeN+rbPwtdLXETrn+AY/CWDCKb6tu9CCsHeqyK
AXMDQqP+p312gmMotEsfdnL2eA4hVTV/vL6e3RKqpWzdvrTK8MELkCpLw1WtTSQGwMoyZp6OIiY1
KrK50OvDz26F7emXnvgSJPxB3Kg0+9MezyBbCFxRrDFAtpVvyOBJ5mitTvYiniW/2KH4R8w6wc8j
HhygowfCOXdOhV9GXlcspn815+GCrfwCyIBplSdgLPnnz/5FV/8nv6Q30oVBIPU6E04F+JB0PXeh
Q9TjuB9JQDZEoPiao8FRa9V81nINUrr7GuY5bVQTIeEnuRck7ahBeg0elYK+SY9OM35x0f0Tm6qq
cNfEkHzykNhzk9XuVMnkF5Bk4E7DNUbef5PaIKsbiCsDHhaZQcxlbokwx+5gST5lmwJYf/bRBka1
JlvLRmfWAN5j1TlTM6RJNLZkvyD+rrz5M7760v2aea9QLN69Hi+nyg5Kx+wyN0lFyXk4n9HdAmLK
VQ9RvjBSd+VVsyfcGuVPtY/B+ZHJjXfDnoy0Et5iXmhY9FDac55GuF6izmwUYp0mnUi2Wvyear5Z
Chr0Wrdj3m2B3lCIyCVOzEmGub5/Ww6GmZWqTKNtArMANaMjm2D+LVQhP80s3DdRxhnpVQoy3oLy
e3CqdWIPF2ede7AQ4fXZcbIK56fW6ZC36kkdAlce2v6RZWzHeF43TaIeb+fMXAXU8HEqclCidUpB
FyRUfyDX0L2jFbdob3O0eW29/IrtXezIBpEYPbDVNNqQ6riz0AZOJCiEXe4K32643RskcRINu/ka
aqHfGSMzFUiu5gLtYsbdzbW9yEOVONmSmadhZ3kl0QpaobeaSutAEqbnlygFww/W+F4RsBFeyI15
ZAuuoex4X7MVkExs3VuDlNHPYryWfP0W0dMcRP2iPn0MCxpQ11gGAUKxO+r18MROTb2Tf5Rmo68g
yRMLeDPPl0fkV/wldI3yg48GOBZ4KJFWE8eRH673d10qkH3ukx89VRhC8lsLCyXyNuuL/tlsvhjt
Z+VT69Yav+0I5rdpYVV0T5nmE7eZAez5VWRvTA/GpX7OGSazCPrJJXZADR7eVsWCZA5dPT3Vugum
U09QPhvlGssDigafZsfaUpInuQ06ofxYZy7rltFxt85TeEtdCGw+6dfZTYiMvF7WdmsrBsY5mqCq
vQ1myLYFAtc8gOzT1HVxX++FZJFv3E1LhtO7nQulLrLuY2eKg4zdlv4wZsUUHTAjlj1CmTpIQCIr
QXZU6Yn2HfVbjV/cVRxEuVTY4mVcRJ+rg6nx4TWeEz0dh1clE/BMDLs+eLa/MKBPIl41vyJcy2gH
BkD3L81NiEw2D5k0W0sm395jri95L937a49CHGl1XWlm+f3fgJJjkf3+F1dQTsX54Ug/aWQeyOLm
y0r3dxQ7wOBKNq/mHqE9MneKSOYe9UhWfV33liVVDEGnqt5XEfJQHaGm1dTiyPmMWRluBLEqooz0
bZKQohpoYFqP74sb3F4vyJScABlt7+/DW42pBmApe5xvL6YgVbIuIfCMOX9cDcqtAfcCbkQ5/wif
aQliVtv3n7nXVTUy7RxTwBWHWqRZBqp0vbCDLaOYd+DOy8+pFIg3VHwxFTPThocDV1qu5G4TmHzG
Jg9zUl43u7p2eXk6I+2Lx1h6QiVi+VLeTslH62HeuWXHZgxMWBVuYDLsSWL/YAR7H3K2eCm71Lxz
BZ0FqlF7owCNgVo4ngrR80YGY3Ay86Pj8h9Sz+lzQM5nDtl7Y+bZqSBU7TjfGd6cy7V/G+KFMICU
CFlGRsPxBxIUr37uHS0BCA1qZiilKaOHE2Y4LwO+sMzX8SRaeF/UcqVLA10D5sO3fByCF/P0niGa
29mcgoH2s8HRMlHVD4l02jugfls9HyKx2zcusUgHZfNQ3/C1Z9fcr9cVSRYxEQ4yexAB9kKsKmYn
QgDRKjrYtmz4NrwRm19BoB4b2vdG9wk6IJMSclSBtT1xRWitkKAEtScm1wy8AWWOgjcJOgQEHQv5
INUH7F7d3D6izEjWJWwyNa6+m+x3ySjJttiFFU3i3Ugpq+6qK9dhLuJaLVX0jqrHH3jOW9drN/w3
fHaT52JHW0n8hkkfbPMB3na5ojjLVX+Up7D7XQd0x4bLLbvRsH6WXB0IL8VDTTnhZO76RFjsA8jH
lU6lHOYb9hDIrKc7hIeaRgGTDCSYUBPjw2E5cJvUmQ5ZJ6EvmuW20LM1OAf4I5UecmdRfiXBMywL
m5w1dm92pqDX1lt9W8LckxRhrZAHnshlEo0hzTAXREwCBgIbB6IkNNV7eRDM4U8HI+rKqFRin8zm
Wrz9Jg6KOtkw3eXbmGwy6C2b/D7h94k2Mwff+2ZturFr11cRj41KTCcNiVsxhLoOxi2Kvy8baubX
BaKX8hCRSH1h4BWHXJbQO2pIFkgt1MSkSS2soOvRSnx9Dt2Mw/8YoY7M2yVTG9GNDd502zFMmoNm
ZgezELuq4tN1iPPC8EqxPS0/MfsGnIn1gsXM1LkA92gMRf4wUPu0ppYHHk8wBgMZr6KlY1xCmJSb
/ZpG4TFoA9KehhQfyjC+QzZxJewJv6g7eZO6wYIorIYQw8yDsbADo0zuKgubkIvQZdYoqVeCQMEs
Abw4FE1Ok0KnBRocV3vpjTepyc6nVMuF5gMcKmw8bMVzWYo9Qh+8xKeg7yV3C3f/N4p7pbLvQa/3
8RNKKwPFe+5TRCrHwFg/Bu6fARGpvnhmFiVgie2De7J0ZxMPHmdUlkQaFOPU7uRMZZOlDSTMd4sP
TXkvKhFoyC6GvEkAeUh0P9vypwAdl1prd226qLWHesKeSULlFes2JkJ2IpURWUzXa7n76jPQMUEd
y0cOnbvCdAgFW7/gkacziu+j//SVtVpSFq9fASp/wTq/wLn0TjNzt7P1IPRd4Bvdmc1T9sX5hMhz
uU/PMm6pAWMn+0XNkfIw+PNpGJR9aHz2Rb6COEfZGm+6SSAW18OmIC69rO37/t6fjbpfxPBuLdGF
k/hamzfl+mAFuuUTgBRLYjV5QuW7LNbhZiHRyiKISCKLsBgoHta/g2oRRnyKrqxnDfCMfxMP1YHW
6IayHY9H4reI6u7RQoj8IJf4z+t6wl1/s8NJUfCFF5gQahshDf+KzgjJ4UW4m1/7pfMX6LNT162A
A5YtUSgR96AR/uyAxDz0wc747wqbe7q+7LqVVWaFfU3GLZlXF5bvczqXHr8Lpq+ycEjYqHl/V0PB
IwbuhmqePf589UojoQK2aNRypk8yfoUd0KAm0nQW09Y4wfmK8tiHO1i+huTccic/eJ+xw0wgyMsq
dhEgPP7tU0BO1CcclqnMsbDkORu3GPMqAk7Q7EIs+pgfz5epRZiKxd5nP6do3rIQz1EkZgK47rAD
2mWkheC7zlJeL6T8gZc3EZ8JOVmcVd80GdjDKwkZBePFF0StxZobYfhUi+KdSdRvHYQbRqaOr4EZ
qpchNoikR4YIrfnhf+ncA8w9+TdEkHHvc5WRF7gMAOmzEVNALLQqfgFwTOJExy41jxHv5k+p8Tpj
MVWj+fk9rXVyaGLM9xiaQJwaZExZhW1YsegwmtU2v/zE3TWgFLAXRI1G6Ild6FxxZitP/8XpTsZo
MozKHfwkXDqa9CfPk4gxg4Lld5oeYZim6f7z8lgFqn6M8+QOpeKfDrGDFONyze+U1aUEsGfE7c/0
iJig+m1k4mf5r2mXbXPvdbx+E+04df5VU4gG+BSgQxbfxjQmIggh/3VopAfOVwGHQXvwYuPAE1i4
qLYHXi+xpLlKHA4/n/UF+xim4cNvfdgT/q/noA3H2/k0M6/6qbjydJ5tkMlyvfCF2nw4FX/gpM/r
qO19dgZkM8GuR9+60NftMKKvORhVNXKKbEKwSlbITXUwtSbJSr5mussgCra8+qUtZEXKM74ouKWL
BzMPFYd7jTiHYFXRT5NBlti5yo6NxtBsy6id7RwYt0U16EQkQwSg2EcZe8fzbn5OXDbfLOrTl7cb
wI2QvIKVhfYy1JyKdmO6pr0BD4QhuF73tRJhHG4Mj4nPquK2pbx3CB1dMa3ac9z4OV/htSt247rz
yJT+UzWF8YpTP0C7jb/h87u9PS6Rnw21JOTsLOc9W5G0/KHVJjICv51ERRVEonUMOm43yi3Bv210
4HVHoy5XFhtZnHYeSPxpjxLvfX5HShomm9tW9TWngM8RMpct+iKXiq9NhA/vHayqrb2S1GxjG0Dm
DeVmVNXTIBjFf24zPJXqhIAMDjo7ZZyC04+s+9MdUQcOrh3d27g2zgMXJfOgcyIl75Eg8KqnFo8D
m/xXpvtJEGTHsmGlw8KX3yWkVo6MTB0qOOhDaYIfVHfA3b2tMR+xxzGV9CkLZ/Xx1v3YCinxzt3G
xrmjmueC4rSEJO5z+bO7xMcHaJdjrcKBYD8w+GeNDs4watbWPntbgoKZKhMs/jpmFHu7yjttXE45
MCHy0IVq8dJhemKxmCieRjNF/nJY+ujSVfuZ9+mDB2NyxWiCXl83L0VLXq4JbbCelBfn46LGNKwH
gNBghs+yzX8aicjZ0pNiO0G5og9dGt8gKVSQQlCepl3zbhefGW3rR3o4B0ApBAwQDhtzKkZWKyEP
1ik6uOUfORWb8D+1s1SJJb5o9ZLo4Jv+bkhuzwgFGPQmlJg1L/DuRQy5LhZ7sNR2MIvwMA3LhN0p
A41qcSTQGhE6N9wuUBIqrcU2MeXAV8D3k4/uVCyMV5oIH443hOHn88c8TPNWHIH7zFkWcqbroXwY
AJe4+9iewjttG3tec0nTH2o4PZBss6ogFNln+ll9GmK5zEOj+zKZ2fLZGrwITss4F6sW0o/y4yMH
iAsJqMQierRvgN2qKOny2q8jgQ7tZTNqrXGSk8py+JgycDEUvaCm9KT7yiQo3Gbs1Q0KKlBkNPS3
Nm/1tRAmwn2SBjWP/vgaQps6WjKm2g0fAbTRVmomsiWjIxil65tBSTyMtFKm1n8jlfa5+G40E6IS
xD3u/wPeUsm6jqTBbIFMUPIohJ01l6K0gnd33eaEdCIm7zfyf+qY8y3AFcx1T3xaiWd3eSmgoUX7
dM8GhdKw8Yc4432uLFg/r71Uh5IUuyc2dy8S5YjsxgJto4GdeSWtOK3QN8BJoP71sMiguUxnZqpL
XNd/AqKYAQr4+/6w4v9C5bPxDRnpCz7urlERV26G2OkNkE0Prk2DC1tHfKeKMY+teufQSWK7DM/2
h6nAT0MIPtXZqDMgUuFrgCIyIZHWjnYdgBy7mULm8o9pqBxxVF0iwcYO1SffbmWsUsveCT2hNIxT
75syFdl3nINczMv+4KE34pxaIuUVEV0Vu9XTy8+DkJBiXlfRv+Ib2XBHy/f/d2jcYUzRHYIWd3F1
4lboISQGQplQL2nf3NcpCJpqgyblLeaZJ1EwNZ8uNpxXnlVOIylM5rEQ6219d/t6OwdRgXm2OBNx
3H/cb1YwWxJPe5inmh5BNoPGs7SMdLPMJrCpAWenoZkyAQn/yeJprn0vrPsMRDCHqr8KXZRFMNSz
fCwLmHFu5MEzMsfp9Tv0uNIKKrC2KvtaCCM1puYhzNes3IdBlUSazUC/v/fhq1URas26SZ8eAVx3
0HToy5kMW1xGfZ//XUQEwaUiGMMB65GvZ925DrHKkY9A7dElmMC8IpMbO5XiR62tnvvsxV3ScgCb
oktOx1goKwq+/9HjUH66PyPmRVxYcWB53iuG2c0peWSWKNNdZaPcyc6CuBXNzT4Oriy/51OoBM/u
IujhgttO267JGgGidpjEcyhZ3n1mvIQImIV3dnt3EBj5nbPZzAK+44e2M66J7ulD2jAWQydLEbuf
aKuKYe4w0BtOiE2WhrhAET0JQvYB0twzu8f2hLuxsq5KShU00cjtVPf4A8iXlbMLbT0uGdiyGHbb
9+yqBRntkASP5gU3ab6ecMI9KbI+4Mo/J9+u/s6ZfI5sAc8XLn8QPoUGrr0anlSsH0hgvdxJSa+V
IT33Ha5hTK/+ODzibhcfnhj5/77oE+v/b0e7UXAyytVAE57INNdETLxDhNQUJbBhV9khN8AX5tb1
hDBQdfWq7CbgA1n2LEOUIO0e4nwr4aSyBxyuol+AH8EhDdirSn2JZ1T6l9hg0tRSbrn8Y/FwjCke
5hOLtRGDha8XYCqAl9eJHOeiIESAy87a0CXbGuhBEQree4yfpVd5ZNjmKMwUUnU1b1O8HrvVTQxp
fiLOxCSNntimacFG/4aekUY7lAqCuOOPUj32PiLjYuckH6Mz2nUZfIyvTulwHmRtJMuGyUWdbci2
gh5cJ70p21Ata2+8s/ZhZF71sHhueXIWk9vNaB3wWPT6+qRgrsQ8VoWlA0fB3dqCfWPiW9X5t6Iu
VII9lbSZ1b+U6lMde3rpHQdCKpr+dNrPXgwFw+0DvzEcFEttsVhEpPZG2cXyr5qFC/n+UL8PRfBn
fg9n8VFp8P0Hm2oBqFAmqv3xUO1kzWjNH4DOiVYsIr1b+xdWEIcyZKJj6oUvqJ4Swx1OWug69U5I
e+3ZlAaNkdWpeRB4MMWZGJ0IgK+wBTnJO3hlF2I6LkfBYj3V12emOIqf7AoCdfczFVfg0pPRX4tb
IaJc6YHdZ3OsW0l9V8apso0g9CX//xLYqihe9vqZmb7y5f3+yPH7pA1kKpsZ1b58CvHYJ7CyGpnD
ynYRVqcsfQcYDAf2Fgb5hsdq//YTvqkoTeCAqzfUD9J5VWssGDbf6fCwKH+lC2Hr3yV6xILivJBa
qdz8ZHrGXcDq3TY0kJOmECea6/7+sHGXDbpjlh2hF/sFta9+FmdwDKmGi96KH6nXIjyLhXkJWkEg
T20pevFJ9rSjN3e3CVHD0zQP07iEiSrCGHfy1zQ55mw2mCtBdNWelDGcC8Sl3X9m580x2I+wg9xk
kcLzIoaUykGA3G0IatiA+u5+eMLf1XtuL3L94yc9j4DYTnPmGjsDc97j4LyLec7ij0/E5RwKnqgA
PpRD/4ZW/zQGfQqBWR5WHORXC7DX2pJbyTx5M0tqXjVfAOqNTGQhg6iJIgeKDzx0pXe+iNBxUfZQ
AXBCo73szz0+oZTuWUtXRTWslMiQ4D8lviXooOxB8HPPUtYC5gkZjcRBhWHQdX9G+EcD0QAfwkrj
xSSZoSPyeymnY7ovPl0shMDO/q87hbYf4xKv3uqptkqWkvhyyd7gyliY/CQ4KzPEnETEa5f7vM29
94+EAhO/IkZOJ8NCPbkvqJP71hXPGUBisErN3qLVgik18XPMk94fe/+o7tHNkzyMpEu0an5D8b4T
Sg+5Sd14I3l5D7Qx5ezCMbpR9AqO6uc1sTkrHCi6llv0qLD8Ba3q1kOz1caOjkBb8KKtdqRK+FpU
c1/8z4SiP9NXqvylVJvjq8KiJVeE8T5ktlV/SCAVbjbqRXkwoKtwLImo7ZYy19R3RCIFzSFfboEY
lH8k1ayEBEgscqKdSPsLT3OWiOAj/d0yzGGo1XkH4e35UxoSeQOCobJOngKY2YwcibdSPlL7pDtc
4ncduxR4lTUi6EZNMBxOwH3FOV6JI9QKQYSmCIwdMVPj7iInvXkrNUNKm7IP0yhumEBnquljO/+f
wCpA2JB96s0gwu5EC3NZwTL1pVOWcRgmUVMS3fm3dzrcHEjbCGEMsaQJzW05/kNYNWO613PmPed1
yIxMRufw7f+KvSkghzfpNweK2qPcA/PBcaPerbX/5QTxwcUWF4Av2/8RnskgWNwo/wThTZl9OVYe
veoGyqkpTKCMvkYnEny52QZ49kCYXPcOeDYgwXuJsBo56k5jkNsRO8w4hWFtBUXEjvIYCscBN6oM
n2aFCN8yXkH0VWVb798jQF3crXPxmQW8H9KhMcwwEqW4zf3+CNLztbpeWHq43k1iNSgA7yjgRP4O
9oWBdaduZrYSJlWKn0B2ghTRhbDjTrtKiXTQP4m4gCYZ3gPozkt7O99l1t8+cT2kAOA4q22BQFMW
1glilEvKUCd4SnC1yEfjdzZTyFsks6K+mGAsM1A4VMBPnzKB2u3uOPkKx1VqLsYaV4v3DPO6eX6N
ZI6RrjusCs0qjWrSCUtHF7AEkXejaHpi9QTw/RCsgjFA7c45a6gOC1PW3hiCuQFivEDxTOHjhMfj
ehZqISb01NOTipw257QjL5exOo+LaJih5OzhgRWGcP+vttABbYwMwMRfsXqQ0IsEehdWv4dqMdyB
u1nIEdDGTiJq3wEHStYWrN0eOSy/k/dUxm18aRaraHD32NtvQnx034Wt3u5CDFUEkH/xBVJMUYC9
l6Nx/7lVUO2qenpkXPjHCYkFBO3UUNAf2wMJfSCU/vxT5qc2Ju1hmlncHgih0LUL0W2hs5crxM3x
diKyH+UqSpHHF03pfnzgCH+BXMuCGjODCMIvNHx+zzTd5+F/tyDEM487o7Cin4KPmpa/BiWJFxPE
Ue8ufFXUeJIden5hasKHBjHw43FTCG24zGln/YOpfDpjRheDuVzFE8dYvWJ8UstlMsPrZJwMQs5s
Q03XYHq22cw184y17KOke3/eXf50QtKX0dAw53M1O6ajx55d1pxBRvtwLUU3vx8R+9+r2ss+hKPN
wXN/icnLaqX+JKMYdvqN3HXI4AxuHnWZkFhllQ9b8yCDn2BrhVssnQxJ0AeVtBHZegfB26F4+KCq
H17SFEsHs2HLJ6idQ5Aff5NCLqZemV6Ce6OHBLrTXQVN/F5ohno5dpQ1O2nebWU8WCyblQ/AlX+b
ezXxJM+40eYcf6vkZMzGZoJl/Dt30H6yJdzVEufJgNyYh1nWDkagupBsv9EGBMlkJR8VX5y2UsUy
gt21gO6zCIjWB4pl1eIHLdI9t7rNY7fqsayRl+9nEqj0zrF9aGJv1KQObrDFABnZuqohQFHnjjdn
EeSufqyLGUi7sJm8T0Id1dERhdicJOm2GMzOf5/PeY2IbKJyTUUNDGaK9x3JqnQpndZMh6Co0QnQ
kddVOtlvB3CeHvvUSvSjxmKbO5Ul9kr6NM6FgE1YcAMw8nxvAv+xyf6+qsjsmhimloTCnHncfoRY
duj8dRo6pByy7LoQmoZq6lfvRsGlsOqxw7NYQmUD9EwSqgAYIZC9HA8f5gGwgDwurNml9TaSjCOo
JOvG8nwdVMxgXy7fY2W/52flvQs0EvdwhpMVWf/G8ypW8FjXJdBzqY91E0ZqdbwDoM1Djmze3wsA
sW5pJJCOMzjsnbxqg57Ip5RccHTNN5ZlKEev4Rkt7qg34dJZtjRNERdsgFfQ7XinMTWrJ58yeJH9
gV3KzhGJ9JV1kSA5VPIN6GT44xG1ZOWFEvHFzKKOkXPeaP4gdXzh0fre2fPeXqTjhRzHlNLbYXj6
RFfQVLZwB5M9QzwGoHIC2eItwqmBeI9wvWsep2JeeF6gemrgtHZGwL4HCSbzHJ11/WdqMfj96Edd
uVK2D4wNZLfWDCHFrnOOHX1+V3mAOxws2ldvWlfmXe3rnNxsHCRU8Y5uiMyRBsxLV4Bw0382VuNd
d+yUdKMe8COmWnzGk+dVZ5BFeAKT09DA0+IFXH4ov9aPYyrIxx25zLN9New74myuCLUi7AWuzwXV
X/n3ifzZGSqoJoFR2LnQGYJ0uNruR7ju3/g9o1aCwgosL8+0DJL4DqunvK5g01ZFjWYSRzXyff+g
NEQMQ3IGVQYKpNiBOb9HIPyxCloSAObYw2kMGOlm+ZgfA4h+UzlLD1rLvrtyOf1j+51i+T6FwsvV
ShwCFuQUX+nR32aX9FItwVuuVkGDbQ4O1Kztus2N9xj9fH9wZ/gdGVzAEuSO6TAlIT9wuCClh8r/
SzXy8sThPo9P7pGE1wzwBskbQWw0hAmKPVKQ+jYWgV8Poyiayc70VhlPFvkZTOYC5CtNjO5Kwmwg
hMsJtVWzBWy/eIWfKCrRbxsRe3LrE8Jp8Ytn5m0UzN1GTMxs6gJNVGFRXHVfMnHQhGKKQY179ZGe
pcI03WC55osEA0+llOcSzYnNO6haWm2Da8rcLrrvpgkstfY4tQJ6tnyCOYUWBHD6937yfZHjlGWq
7HaACgJJqZUOvpEPeC97MlYCNpVzgUEKC9BWSoO4dCJ/FDlpV+EGVajdmUrxxGk0/qDMLnPgrQC5
TPpadwugQZuj6MuVxufHgUN9Qof2iZyRmLCL7FJAzf6ndc8oSKsBx2L1NCWDsomNddB4+8+/tLzf
sFr7xtDe3PHdEn7wbnGZLDtupWJPsyn7EGq7jiRtyDPkWPS+dxkxWRRJrSL6Y/+J8aW87/IoG+p6
0gHTrnm21tL2YMctUAkV5SwoGp4DfsZVMQfLeHMiCevCMcYDZx86IlFRlZysEi5kNulKtK2h/8Cf
UmTA4qxedj/LUq03Zi3G7xT2r9rETM3BB9KTTMOED3Ijjk4KrYr94TwpwTQnJJknDu9JpzvyEm4u
ocRIBbcL7Nv17S6KthV4KanemwE7dzj2yttg6RJGo1f90HfvYdP5m7LKGCoSC2UDxkhvPqrfOclD
Ri419payZcdyn343u07sCw95bIfclC4wRXCXnLgYklmulf7qoprrhnEQquwEE3XOTN1F2SAR7HLD
RmUGY4ncR+XuIxpqR1B+VITkBiVzluUf1s/KjzAHdKc6mCmffNTLYntUNNQf0NLAkE3eZxz7VIcU
4CznY7xSbsFOmTuUwyboTD4Zxy1Nz8V4nzIBitsaCwgad+6m8VLbcu7NdLWGUez+KX6rMOPmzW/I
2bHXCBwcuh6tcCJmsC5XtzAuZQdc2OnwobNu1uzf0vtVlD+3Wi0fcxtM/qulIQaNWoBBe9oNHhtw
3WHdaiE9C90+msH2h8MHlaKJRNS/WpTgg/Au7ltRvjXujz2GGqowlLIVRPLRq9roPx52XzEq+mbQ
211IyUnThG2HQlUvQYosgR0jW5FW5Lh2hGfQ00Gw1NxkO5QZrxKB5tslSHZLHQpbl6qymI6+6X66
1i9GQjxAiF9tLOeY+XsIxcaT+iyzATkwVfXSUfnsOguvInqGzZYlFSc4wdLhE++Tg3bSls0Z+gw6
+Xvti1Ry8qoxTVXtnll8C3sXG135Y1OHP2w4Z9A6myo6BaWZVINaSBdDCO8mM2V/yfcfeCcsry69
i1EMZTB1ib0pEMAKhWQZYu7zjGzxxYoGUWU5J/eJHb83yNoAVKXrJT4fqBsMSC+blRhxf+jgsNHK
2l9apGVoZqi+ei1FPx3u0Bk8s/IE3yKfuw3zdJQKoasGyS0uH/Dt4X1B0xfdKZ98S82Dw0kyIweN
hkC6GTjQqEu1Fv7VVI8kSq56d65Tb9pjU1tk+wTSGNDw1cTaHN5Bcgxli38VVM0HA/Npx0yVqx6/
z+P25euHN7h5TPQ9qOy0U9FKr2cRbRDNU6E3UGEGwlBK6/+n3NQEiPj37efgm6o+SsNPyJi9iNUv
WdVXg4msNAwdOBxTBJdLua19tRkyM0lXHjkGwmDiSeUFXq7Dk3RmhGOnXGVCnHZmOIR/Z5NXwUgj
Laqh8CnhJ+CWhOnR68ox4u3/bD9vRcUyxhfrj6WxeEXsipxCkOdxLNo0AIOKFCOLF8TUt+JT/10Q
I6BeWcTficRiKuK/hnLWqPCcm/ZchvVJ3mcLPWQieV1xXKdKBUJLME1+Chj4dz+t2DTG+Gvbu888
OnC8KiLfG2Rg2Tmz5OnIOAs1naeOtn9mpgdZO7V7rf9G2FpRhun3lUGgUmY3P8WiwT+e5/y1bUBH
Yy51OCHnm94BLQdLX8oOabQRLGfJ2UQFOGa3IucjW5cCYNgMBlTQERWNdW/C0ZChv/XV5JObsc2y
W5GF1+p8FShnbTqFS74i9ylkZrQFi8NjQaOarc18BPBBEiTbUlZC5cVrO5bwuYOEiQJ2E+zBU3sn
DFfCxqJs1wQpwcoyoAPpNk1fpzReRv3nMAxMbpGPiOs2k9DB0Php0xwiuwlahtAPKsZDxqnSaosa
6hojkWABd3aEtEjIe7NLucefvUnRxhYekSarqnYUmX1ta1IsbqrBzc538uTxzYHd/+Z2Qp5ER8XN
L+JemDF21wIaYsBKUWC1sDgUQokhOmbCaz05iPHpI7UpqxAi+IkWZV/EDHDttqXccxoYisytLzi8
+5Rm0LZgRuCTr9Epb4FvP/qGdwBEJmZr08k+YsPdsHl6JNuGeFBFHRVo9EVERpdJV/F72PmkbSuy
aiAyx2SQL21863TpOW80NbwBrJKwk3glArGX4uRYhIawPUA44U0X6EbBwhM4+FjjUm9CGTtsU+kd
cGAv+LB6HKbvzc3zT2mzxsQ6wgzUYqMD3KnDWXQUhiymgWTXWxIj1a8dWZWBDcvXsleTosBTA/Y9
91Hs2HfQJGCODk8Kmw8eZLZV3sOfyxjacx1buxCksyRdnONb5M56PSBXWl7gy4jgFZFaxWm6WxUG
vGQJ0OT3ha1FrkRh52ov638HOgww0HLZzpXrdGWsnNimsi72rhsECfYO93zm/ACbpqRp7a3NqLSM
71wzMqgCrv9jQ953MIpUCjIQSOGmXkqrb93Ejy0eold2By0qbJzTyEbTdqKvj+vIeSSWsW/LF0O5
rajZHZnjJKdt5MuebCKRr0pIzRJC2AuJgsEVYfTsKVhGKhft0Wpr8bWfySMtyZKgSoizPck1KrNg
8CZWmFijuzj6LVqYE4W712diiIbqrePRvlhSWb7vSRO/JNIbJjdcY2YxkM1wJ8mx1v1v3s3ZUIuF
7xak+5awc9vdv4IkWJ7ZLRzP9Dm4PvMcLjk3g34J8/gw1zTAEM8HLYMa55Edr4VxY8s5La/PBvCJ
JIfKPMNDMrOoNkUq4IW0PulfNb5WKdxfZ2r4jutQmydqBkY62l+lh527B2pYhec11U+yUh65Jl2c
k1/lBE+uRxtu22nuR0NOo2ZW9iFJ1JOVLBmx9MPa9Zajx6ucu6E58BAiyE1Yx9IKXal3LPFgRmC6
YcsoP1BweUbXZAcdgmeEVXnoZjy6oo5zvFbKUGE1HVLx1LnhnQnIckznfRzLz5NAjUcc5v4m/yHC
Uy45f6NwUOsB/jy5kT4/j7ubxp00AaiEYUCBR8D/WXVLhvW9HedcNQVWGm8iyNVGstt3aujCOAoC
SwIqaYPW/KQfGjn6QOMrBJuAxp78RH8wOOwwk6F0DUF8u9xKtl971K6g6H9F1fivyVeQnpS9QXid
bB3jRwmbqyHoeqeFdPTyH8UFw4Hf2agwgUbPDkPPvwfT66Rrmw0nS0zMXCJeEvTjttm+WbLxGU4r
B2kNAXuZNzWvKnB0sQTxVWQwd1bMCrZ4OWupLipsJru0kfQNkezWWNtUqou0BQuLbiGBqSO/LcrD
AOYtl/ckqd0YCVBGEKFPAxT1q+O0jfpeYIdvK/UDQXMa0/TZ9Em6xSPkTXk9XxCEz0lYM4NLcxmm
Zn5AAwZtFuuqQATcvBR+6jeVoTUtJgFMbvbhgHUS1fnw17qzUV2vYEGXMU7R1xxNKmO9sCHxxrHi
FStjlihO6cf5KsP7JAkB24S3/+tZiJy4I0zM3rRVnFMfgX7AJ628OCIoZCQ9RalmUrfQPfvvnQZE
vqmthe4wuM3gKYyJgAQvothwBh6FTKwPDKKmK7ChD0zzYFVe8mWx7c1fmvNjnYJ6T4saDe2FwXOf
Fo1LRPK5wAS2iGY1L1gOQXw268my5JMA/UKlkjsNtT72JGab2Q8ozrAY+y/73yf9EMD1fnQKKXJ/
h1Vrk1W+HXvmJ6lHozb488zS4KWkl2SKwVtGX98dZAY+az9xxNttGz/dKk5GaVNNDLn7fmT9E8VU
wqkUYGS6lk5VJ7YjhaCMdrWjSY3dJnKcTCG+oQteR9pwoKJbBqxekZFfVvzVPr6I04aMyqzhkviO
ZOo1hPCG2+ZkY1A84IGfN/C0tZLxbUtPSpqPJCvPP/QM8Iz7I4KnEjV9bJDACaY8zAdRcl6+sw5v
b/lTBHW1OrNzzdeGDNIposREvI+KDIWD1J/sEZK60vMEiyk5YK4IDUBsOnIxtro1X1SOpgJj4n+W
KGkzzwANhzaOM/ElgK3N8P0Ukgjva41E8v28M7gsqCD3xcklIQnC9bZg4C1zvlkjIdWEhfw6p/AV
59dCHZoeteMgDekR56GTapfDWikfvBF6K/pourf+b5lraK8S0GWs6jBuGtDOQQLN814QjUjrm5Yu
MdU9TZPlDY82S0gFQxLt340daBwxWeI4XQ8W8n6q9etTHoyQrza/OlKhaHnKzCfjUVrMKXxqwJfG
fOJiKeh5O2rqswt0VFPfuoW3218rx5rza5TYLjMAoNN5XvgKqVrgEPnsr5MrDUOFnbq9Zy/YGBO1
TiqNQ1CWAjaVLbNA388u0zViuE6nnGMWbx+v9XNS/wF4M+SaIVril3uMtqbXXmBtn1/UMcEFChpX
NVSbj83GnH8pyYrfUZ9z+cYv2BfYXmFiVqVFxPj+HClzvXQATPpAp3mIqis5NQp8Ubyeef7Dafmo
3mEgAHOWpwZ/CYLL+5rVHU/sm/8ngou9Sv91Fyi1Z8gSGeO5F4jyK/NHnTuFBZTEleFmPeQehfQx
hfpJqrg8ACNXxgPAKEhJYSDiKOAx7S517D+71oqolpSyRLtWnhJTVV35qGzd4INwUp9ORGFRLSU/
Lfqljg1Eysx04eMzjdwunBAliLR3JtLNuS2ORmjxChvVggx2JNLNSCvPfENxhFCFHphSSF5GLboz
JJJR9q/liXqLDeXrwVIINses2lTIlGBapGW92lTaKlXOEPiruhqr/YZo/jMMNDQ7Kwb2C8EFe2kH
S/Tn7KhnGbdbzoS6/KBzO8T7HhphRteq74CKLqiP79nXWxqbsP4Gqw5eijm4siyqv/f9ioLYh5lS
xEl8PDXt3tBHLFb8+0BeUZ66rIvwFnqB23WquTB0fDB9L1sJARbH9Ise+hN274I7gmqnjtMi+Xwi
m/arfKoOM+grLCviQ9rAPQgWtJ/qe9czi/TyZf7doD1NphztdAP6it8oGSMQVqpzJFt/MVP8mkTr
wizv50dMyuiC1lH/DLsMkqcggr619fWs4Qt2LLX62zwWKUC5zRU0zY2OupTbfgACvJug9mb3g0oF
A5R8djoD4EdbqUUdV5+53+LDYp7EHYyP00Cy2DXbISL3dfXLBQWn10HffrDyWxSYfyfumaMb1N62
e935l+9asoC4r8eP8mjSU8X4BgayrKO4e9iassG8316SA5QZXPFVEwCrP/URRNLXInGhTQmasb3Y
R6ewaVxydD8taSdY3QBVWjQzsH5h1J/FcFObcMwNCKXiR+1ovQfmy7Gzp4RV7cjy3wLjSG3eq6L8
JEKabjYgVRiIBnuWXKu0549ToN8wm7UzKWYOqWFDTdklMD/Elg47g4Q3m0Jz+z6dqr51yryspPLw
uzTpBraJoOaHVzYeQ4m/mAW9Rc/18YbqIeacVu3/tTLHh7EwZcAJH9eCEW4Vaut7BukFdF9ayeKb
PmnhirvIYV390lrDgl56LtxpdWXan38SaiLXt2h8BXruKdxXGb5KEZsKppzCKwRz5gHQBsYx7doz
vye/plZ2o+BJM5b5ss6JmjnfLKgpldKXf8MFyA9lDUAksw7MtU2jFHlO+0cu4YYyFkEjN2TrHFo+
/EjdwSvCUUycM55T6yUBitZUFd3EFxgKAj+sRJyPG1z4koYaflr4GeJjuytb6mpfqNQf9nsbTXo9
yEhJVsMM0RTtUnrcrseUCyRoPWfkaEZiGtud+6ELg2aoMrTFm0BUyU3a44UJRwvDVK17Q4Ejpbec
cA4RjeSs46pupTehwIvkCulsUtqu+AO7f680u4Xt2qf7edm7713JdDKw+sPBdZamngAYxUZ1tB6G
8J/C/CL9lSrCuzuQcxu9PfFyuowxSIpTP/fMYVVveqLGdEnKdg54p4Dsobps5rVqQ+NihaLCGv0v
hKX/+y5Sm6Ndq1B8+q1RIdIqy6RDmk9pYoWJ7GysjbLwmMF3ew1a5nq0GRNQiDRbncgs7zi7o2Cf
0fx+aa5qET6Pd3YHw3pVf9b7N2QGanMjD1teGAxQAVBfQguiv6oYqWkYEbxhjS8tvACXpPleZ/Fn
6jWYK3uFsxr1jvp8ytP1Lq6K9uMbdMDmuu57r40MyEXseP/O95fbqnl13ngbfVpfqA0JeNR7bpDw
OuCokQCxYPejvtY8GvQHW9xqP/WELzU7+99HVLjR7b0hNYD6MI0wWL1vkA8ZkRGZVGd4zS58ylIG
hgkLmjzCDEeOWUzSN2XEqjfSNhWRDnJ5lWl/L8gif6BM3+oMZUze9AMI69P4d1Mv9ZTsjjgCFg55
ZKnvxX6L+Q0AsgeAUZlkEjV0A4GU6McBJOeIOez5Mai1bA8YlyYPzH599KSwyYKh/Is4oVOybSll
G/NCap5u3Zf5OnzLKSswWsIWYdTapTzSHQIUmCuoJ00gxwGw8aPQ/ENiJq9wvqPCxI4odTiZG3KI
CVCkMiTmr0XxDgxaZdLa+WGB7FEtdDNjX3XInuPEm+fGY1ezICi5jWsYdWnbZz2CwindONYppLlp
fBUB4V/0gNAYMB3ePqct/pKLIp9v7F/yOdkcKGyl9XyQbeJ+9rXwtVqAIo22jkS9hTTnip9Ubako
E4Z7TIruih8uGFh5fElHlWHSxk4aYMQY9OUn9b+2dK2ND7MHPoSU4O3v7nfdJOu51h4lJrvaED+m
vDmhmRA4RzckQU6FvJhmOxqzpTzoic66xhBS158yaR/hnMtsgSuzVQzAvaOOOenpX13K7rRi2gR+
EdLv4myzMLxzRrslcEXIshlGKrX6qhKIBllzWzh+r20vJwHdpwwoFgv/XPkbrfwaCovNa8KLQzsf
R6s9GtNIM3gp1kJAG/Epn4QADcxRBx58QXIVqcNrzeIfYlfloMWqgB6N0bXladj5rophLqirpQT1
bC8NPs32yq6VP1Ikhhn094l2GoepoHNTr9FAi8DgPh6a6G8ifSTe/DaD0QrpChsYSx527XtBgwXM
OeYE6AICUL1vmPVfb7cqAclOAPVub61cnhF25JPF6f4WUmGbsqi9XENNPkI30JOkaCb28UEfXTF2
+gETrGuMvZYTw0T1YdVAYCwJxgajv0WrvpQEvqfj8PY6tW8p75QjBJ4SY+m7OY+BYeC1Naafwf0M
tVgsOT1nU4od8vB5JjRjEWpoZIjLL3UpeHHC1nMYYK2yy5QZjeMSZ5Zvmyp8glNf4p4DnnfIP4oC
/3x9Z0S5Vgt8Gcdbovh/IZ94k+hnb7MauhJnWIhpGs0aMk8PUa8GJEIGS5stCsyVLhvdipzUET0X
P9kNndAFpM9FXlDEIVvwsL4/2s2/0H1utHTFtbw/zPnm2azW3839I09LEl4AgEtJadjfqKYrTFko
jcd4qZd4ZlgpGNUMeZlMJ3MGtiAqdBIyWa6eJVLEM77QChhOCVXI1uEzezBvjHPOvsHg//XkitJv
jIiHwXo2Sq/ibqxCqT9/riPlGZ642tRRcNlBzjAQyN/w7kZegBXzbRDLL6BKVOz7zwGBjLmiM3Yj
QMd0aNHgHmO8d17sAk6lcGyPnPrCJLXF8i19Wd9YVDmRKl8CYuBG3pVQ3VGG/cnbwzqa8vhlIsiZ
hkzgFUmi7lgHwl2om04lb0pvD3XIS2W6d+NQ4OXe1bsEyXKoGai8GZ2bGOA9D6KslR98D4Sz9HS+
GywHUAsWqmQMXpiVxaUv3oc/BqhrpI9DXbAL7w==
`protect end_protected

