

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
jmxpJaVr346lkZ1a+LoDVE1gRSFGUifNjtRZEnGV0oAexMx3qGrmrMofcjVsktZm1VmWfXDcztXM
2yFG9i0kgw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
dOSbcKbKyGmwastHjwhWcvg7mo0iC7nVbxSBuuKDePvzqRHFROAJKKkq6GTW/pekpDi7EYOWgoc3
vu3a7xd2BbB8KPxJrQPbDcHKKLsfi9Qu05pG8kNfZPTmVPdeph29tJwJuOY3Bue31aDGpBx9n97J
il8TNCf+vPPl3qN1O1Y=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
oj1u/InDUMUdQbb5KKzCbe7WKv0Q1mJ0hkD57NzdtON+OYFVa+iXuwhtetuyEkD/RFkOZub0bzay
EGz9mYS8JrDX4uhqviZ/lNeQvlGcy4m3aXFV0BaNm28dZ3yofXU/BObQHMb2AJcvSvAG3+NK2bRe
O1i9rDUCI7L9zpBAsqwfaKowW/ytJpmf9i24R0N1DPpd8Du0b8109OjIyuP0B6/WOaUz59+u6rpk
YBt+RO2we5Eynllzej7EOx457Zs2AfpyYb/scT1J2gg+ITQOiXue3l6rpuOlPDO2s8UVnv9AEDol
dBES1PgrY5H3iIxtkySbQdPn1RgrbUXGoP3Cyw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Nf7SNu0SV1jFULe1qPx1Us0aK2tBb+6HkavjcQAOW7vm2bkkBw9TTTcBYW2ZVktL2qtI4SdzYqok
Ur+7+BvPVL9Si1NxET/7Dtm+YCiSnZRDjVxRHT/nOJoMkCyfwzbKJ0c94Mhpx/IIVydS9opk1YOK
norD0fiQ9NScYfnzaaY=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
gGrec2cOqGtm9E1Oi+bdp4JmEjroHrWUud/ZaF+TGsozi+qUj2kRQyVPKMhdue0iIQELWZ+mxYUS
eLZifl90wtAXYuJxD08Z4LzdxHrYp8+GuCF0avDcKZR6UMS6GdOF0ZR2WdDmkxgQdaVnCHNmLABF
3DC4E9wBUl1YKYXSRH2xT5Tm/cD2sgS0Uobvp+lTtO/g/wUBgQClX1AYzm6JvXG56K4a0tlrJqsS
O19bJe8ailtvTRagvfU5lh5iVeppPrENq5fwhz7scUcyvohRe2r5jixGcPz5bVE78eEpH4EwzJTz
GDGFrWw8qJ6s5hJeVjOB9tgbpdnAFcvyrMEGaw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 16464)
`protect data_block
e1MNZfheJ1MNvU8RSVyab/YibUPFxfcqxmQ5nW4TiP3RICvW4W9Y7yXhqGOqaXtOwK9P0uQGbXFq
uOPAEfv4NwGlq51J4wxjj5HUrW2vSpFvCvgFPhW/yEIEpDSw3RSDC0DqO/Aikov9+eVS4PtbGH38
ChXNyN/0X+/IJidFefvtD+wi4rI2FvsXVXM42UCExVvTLZThCSMdZimWP3xivft0ExMAyLXg60VR
Z4hLK5wT+mOikQNNkq4yaXTmzFyVNaTjDjXG0sL0ADKrh3p6c5ALGhdxV0RDy2VbKuIJSVNfKNbd
n7h3AaMMRWTjE52/klD2xxnwu+nuWTGimiASr5OvL8W81FyH7FKU81pd6RCbRJHQAMJy8DwwjfLA
m2pDLjvD3rk0InNd6tv6EtBr5owLFfj5Qp/TohoXkoaV3K9kTIVO7xbqBk8ZPOzN0AVCvGRCMieD
2OV4szEHvlzzvHZiBFFe00SKkKlhnPFDV700N23vfqgy0k7F8ghtoY3kM0U+OXdX8186syUdoiBb
HJpcgNIdv9Nw1iNWYe9ls7wy6b/Sw3qukdy3I+xssGbr/S2dVbpMl8xlgmjaP9mMyx9MrvU8IfJN
gMBYgC6oe2PqkBqoDUp6GaejhQfDExZ/NPoGYwR6tpf4R733S0tCimmqYlpcSXTTuRiPm68u2oJM
exDdCx54nTfSuLnIUShQwAkjlPgmNkozx9ZXMS1pZ1y1EqedKQTAxypHo6h//oJwxYSteknv9nLE
Wj3aExEugK/4sq2//x2/gX1zMpCWC7gZ2q9ElwgcXZrVcHXmmvka0j4ybbKo10gaw7iGQTQyAex7
LlqdabPTs0TfT78Wf3fnfnQkhbs5/WXNqvrXYuLPzL8nUUCdmfttalEjTsPsqTBDzR6OjpzdW8qf
t1AKqSA47fp//pokAIp6Qr9EPnrXdGzICWv0oBIWyoRopzSv0AyUq/YGkURo/U0gm2UbwtBkc4eL
OBk876nipywQXfI2dbgUsAKe1cAQYY0eLLjqdBCSJ0gXZlaZEEtniFGcmHmucd5vPVrDFj9jO7GO
EnT/it0Q0Z9uqp5xivdNYYJak2/30jQSHliCfDNjdmYxEL5U1YWxpD4lk3lhtuZWYUUCbzbf1rcB
te/AjDXvUi6pw8sL74uD9HazgiMUGS/IbTnQEJfWX/j05lQkRf90vd5c+ILXKy3bzEqrZun7PNP9
WehyxcTXTyJXwurlUlqvxXAoQHdJLfzM8efuMTw359tW6IzO3YQkeVpllF1ch4lhJh4q05BkryYS
iD7FfnHv08PVxJ48gpU11uQNTIcOf2Iv2lpBpmmZUEqnC7OxN982toAVI6L5MZOTiZd64i0D5SuI
lJLg2J820WVhTclgotu1pN6Ky5YGBGim6bkocEE3WJIuxaJXb2y4o6GW2p+wMeL9zi0Hv75v0e4f
SFoJ5E/UvzAVFrtmYC7coTnNlvl4TckAYMkYGo6kRr5pW0TW+WHEwaiqLoQZHo1NWYq5vi3giaAv
DJGIQSUe/W7yzGRFo5uOlldqorBeHX6ZqlB7ygbKXZhJzcP97zuS7dcTtK5UnFuM7Shm+b4w//fJ
HH6OilPm6gmeR4/viUkjF5G+Pg5Wvozr9hHKcmLFn6zVo6kNLnZ7aAHPs4lkrWvA75UYeT4L7qT3
jFdnn9hfo5QTvGY2IoINV4T7jmJ8lWaHXkaBYFIsCJbCjwTxq7MNvWdJqIWy9HUIvGWGcwlYUfHr
lMxW37lwIxmEsFXbBcYKzXyTo7Kt4mPC5uR0UtluAxtXlA4927wmG9dihPygAEg0UGwhz0YGRjKb
Znos2qZQjfjIxpHvfeieh0zDFIQYLsUj2erlWbdwwJmOafwjuWSpH1mFBE1ISl46gEorzjH87Na1
XO6R60LYGZh+xLxRlq4pb6+Ovq1u2jI9033biABksg4zDt9sL1VmJuWZ4hhUvcQFV0ICiv3UrPTd
WsiMiJ3QAHAxdavsUc/oUr0S06TEPWujNmFQ779Ai998+flwfoRz+QCVb0gYpirJmtXaAPac470w
wlla/OFq5HBhYoCKr2JIjJzUv9Smx98UfGKqEYF0WIg7wlIwzGD3eIh/0fhKYHqYHhGybgHe479R
yJeJfSX5Lkpw6rUNEJAKBHwRUPgjnTBontv9pk4OHrmaWthYEaR6HxenRZm2UTsa7/vkKpzPeNy3
5ukm7E9uJi7mD9dyXHVZpsNI8Zkf3YZ7GH82Eiv7IrvX/ydQXI/8qjf9a2n5bur+/cKdCAKo8Rfg
Vdv3bhO755FtueUO09hyAfRU2C+45p0N3GLJKQsj8zS/ww/V20CQ12IQUYwRT56Jd0urk6VMQCvv
BgPeNoLLlXu4QtkCaUCuY8In6EDWeYLxvquz62h2nBHt69E6ysP34pde7+uLgHQe8wISO2RQkRys
EoklzdUSpMIw01Zveg64ZuMYXUr7/f4L9E+rQrj1KkLguYnXdMc7DHe/MMZx0YlcKn77fL9xcyc2
NAzmjxE0Yne6zYSfAOGp9vvYy6Iq8yCxYG8wE9JRAGNMzZk5lMUF+G/2Zvw+dFKxzc9JeahYAi2J
9RDUSvHpuHNBDv0Dfx74/GAfGWvLKYJYtuUKVAQYZSJgYuErICGjfuJegv4LA4vlvVUccF1Js0js
YRJeHgCtu7hcVXwl5A9mWy1hhU8ZoOIisk5FwDyfIKoZCj8OS/rQ6aga2H+jdZuSZSjUOk10+Ozx
rfxjE6xrxEO+CIkOQqMVWEZoKHPWUn1BCN3eIYlvjwXlgEAcaplvBMtld6lsHV5mgg0P1RLA2Lna
fdIzJLjdSTgFLFpSK85kIT3kKlsHWSIukxFn9EKE512YziKu18+AY5v2mBmCelU0QpYbErjmR/jL
zYSDF+gzoDEaiLIiCr24/SJN9ISqtptihaMW4PdrALZHXRysBPsYUW5IiTSGXbcrDokOVHRaJ0ae
gvqrKkXvdxivWYI+Lh5jGaJeGrxxDRUKmwvf/dK00hEvvaRcn/HMIwUKaAxycwFLHarEOQXW9uN5
la2BT+lVYC956+mEoTB7J/3eK7CiL83FBgYD37SGPGsbddLMK7k00hOQZElpBl5SDUy7FOz82eO8
fh68faft4xQcEqIW1WvJTpMCP/YL0wlCW0eJSq1KGGcK4gZOq/VCqTvFAXwCDNtFqH4PCIsnuQ7i
bGG4hgLZWCIm0fgUuM3kByxa70UnX4CnWlj7QnHNuFfsKGfYdVjlCn7GNMvIHH1vEbJarOnquS/q
1NqOQOYKh2x4QEBmUgy/7krNeXHe/TG+A2rF42Nl2Ga4mEg+cJxTAiuoC/qWXqzh+uj83rr1qD/b
n0ZZImr6gYErnUjvEUJMuLoA3lEsWcKuwNLVHOe4H5DxxGijfsLL5+GpCEIbY8UmPsu5nDHtjhqx
6pSa+xU1P44ygKSOVJ+ROri65GO2xxTD8l5maxage+jixYeukcoD3nwyO8g7Zo42swrBu+7DuWP1
MusuZ4mJvmSJm5P0QPb1IMS0EMTfn2QDjZzKgDvkVTVDwcA9KJZLGFyTO/FmBVL457rqcy7Nyhuz
M8yBq4yrPoPNqkINeEVHT3ncqZuXFYmC9NrmJRNd8R+h826MIIT0q4MHJ+B66/Iaj5NtdrvojL9e
9tnUT+DNcs5lnATZxhuY7Alvg3DSb8d1RGtFqm9TKGs7g4HHyj2JCOY20pyMclEpwBWYLehR4JDv
HAh9MjvjWVr9KFu/J1rlzAVM/OfuguWdGUrJtfEjMyXQFaNAPr0/PFR0xgxYeOAnu3ZZctUZPsp7
SDsj90lqkC7TSuGms/3Vf0I7awmxTX0fHs6r/s99uO6llhhwsLjYBhDvSY4NZ3wnJ7HJTsc+h60H
5izJKQEDvAOtEBRiAzQk9P7dN30Rhk+0nmpiX1ynBsKE4WLW03tMH6ez4DZTY34Q9L9HKTjx3gZR
JHEBT7atiwRyrERKP+J1Tx5wARl1gbJMkN1KlW6+e3DEvjKcM8CzL5bQXdYQnhJu17sQYcAsO4Jc
/tAgRrkjg0v7apOeccEwUKqAnefUldMVi/wdkrsBGJJewbfmsdRNSsQ84sNltnET0jaCxqcOUCf1
3tWmhYmzlabC4o1g3QsIO5lrBzQWU6dMIp/vZuGrnGnvdmRzhXTs/uxUXL2bx0WOfna7VDfwpuZ6
fR3LWN9mV0h91cehrfq6sIrxkxzzCY03tQ+JDNgtNGCBwMyj5Fqwwu00oKjJjqUEveVZpUg3jIls
GxfWP3PAq/fDZgp1gmovU+idzD3jwGDk1mdeTMf1ifUe8hi0Jh/SbvyetWzZtA07aphHAx/Mx+a8
YHY08SdmMBJ5dCnUPf5+BuMirKv3aKzdr5MohnL6kxPSDTY+010HAgtA/uWUaqBvd2FVXvk/w7m3
1hnxrgNGgXv0HGhL6W0QmVRBQCQCZf2xMTv2AvioP3cYrV+Lgu74SRLvX/y3IoaWXOZ83SG4J/RM
CrXMBVKJJKONA4yDRKOMVY0k2+NSx84kjIvU3qwlTbTDvjkHaOImkmO5N5dXVF+K3QpzQx3CyyaC
eFAPZZmavtOqQi0ZiuffBFILb/xQO0g45zVbNsoF6DMkvuMgwWYnJbv7xRXzztCJl1DcLQOJ/Mpq
qx2toETgYelXRfhYmjByMB9RtMHhuV8+RJSXFafXLbl3JDmKWL8B7WbcmZbO6AvU/3zUDYdbYhlM
usHab2xlSOYTyQsuJV0Zu8gOfcg1nPImx3rMoWY09EJsthnjtSuj1WcC26wUEe8dX8LKwgsdA3Ko
LY6O8MGsl0ZYE84GU+cCOJX3UFPOTEOxk5kwECP3BSSzkJmFQPMYw3nIyYgZTINop2K9cjSOWesg
UGVI1Mj8ErOx2YnDMmwNCq98d8G7C4QsKKBqWGMW3GCf771vVWVBHk4RpbIHh9uRmh+GUFfdMCTo
PQU1eeYqsT3FsfVzBm72MOX4X7wPA/eU31jlWOh06VM4KbS78jPgzByBy+1AF0/9CLzugL23IBHK
LUPgXSEMllfgEYG6tjBntUZKQxjg3PVGfSULBlbSRO8iWxO967voSjHNg+iQbmK0I0qILfsF80lN
Gog7Dt0e7bpPDnsvlq+41SULUw2tEtiY8AbvD9O+ZKI0tQS6NRFRYIvoxvv3W0rBQIUOg/xPR90l
IS64wekqHU0jaBIdHrNLUHICI+qIXGAyiaN3to/mo524ri3sGqcLoL5UwSzuX/NB9ITWjF+qmH0n
QRzFTtC7+lbDZNDA7XDu9kqAMN8fetoee24UF5Apoo8ehGn6TyxKsYK1DVfFAufmqA9pyjDTX+0k
4FDLhfHNDtVCHWWaah6W7Hsrm5g3a1uTPdSd0Zs6NysqCE3JM3CeQRRCzzpj02JstOcwsHYxHfiv
n1umqOFdrwJgiMG/1eDxY1n3Lrl0lX2F7LMp/tyIjDsbk9ysV4dNtZuAqS4Xfe7nVRoVhzSaZ4Cp
8dFIOanZG/Gwb41y98KYEuOXPPto4xC/bw7ZAmeYDgmmiz+hXbL0FF7ytMU3Mj4ung+buBni4hOd
0TUuw6jU5NNFvOboW9xuzJN8b+vimRp+DKmqkVBN1Di46ZEh+LaNa1Pqyx5l44rL3m7GYWFDbp0O
gz0yOiMY/YGZ6oyXylG3AZ3NvfOzZY4FGhpKg3XuT9hHvZ8TuACJdO8vALaV+Mm1JvJ75vnis7gv
IsXEWCIIUkrO66L8tLnt6SuZ8ODjZhcChPfMaMITDSfneE5vwH2mnSLlB33KVAgThdIqq9pciXEH
G54ZB/VEXfsw+P5QnvanQV4279AzLftWqXIoUNcl80C/2cNiYPv/OSNJngdryr/lTv5TJKAzUNju
g1X4RDknsKQfyglIPV14EO9dPhgj2PI054WXrg9Xly5RhU1ptb0Z0FAy+lxkJmh3/OJKz6b9qXN8
TWPXZ+ic5pbP427ohCAUxvAudUBSzc+WD0RCwE1MB1SKF3UrqKm6bJc1EOQ6qRlCuQuQTqlO1TfD
rbWV7qNmt0DVKbk4hLQHoZ2A9pkBBWxebGligiFkApbk2VKsrqcDaFNEu6JTVe9a1IeQ3tzkPMMj
iSlrvXtTg6PnDPB/lsh9y9JPyrMq34GQ3vo+AUaiFzKKOlGkVjxv/VMvxi5gzS2d/dCtR8/aR5Z3
2Yf/bzwfoXsEQkdL3w8/I7Y6CerqDiyp5NKuxUWp0EyTo2g7taSUrNGFY6kmrFfuSBvbyK4e8ezQ
DtR6cxQYRw78eRySGMB7VAwK5evXDq8L9irsuG3y1au8c6bcoOdBRSPgauSnBPV8EXJzS/Fq7mC5
PxqwmOeWcuDTrraIVfeWsgrRVSUz7lBNXxJDUv3YnWSJ+d8nMBatsx5bYZ4JpvQnhWtefHo6yNHG
VxdRX3rNOxYsyKeIassJ1GA7xAfzKW5M/lXoF0qj3NZo24QZwH0t+WaZsC1usDVh3ObHk0NNtxdY
I7BRYW5XHjWwYd+sVVM8LspqR9zNMa93sAFUfqC5M+Q6OOTL1enltGolRGscUO9yflcajP0Wvh/R
b0uLLJJHb/dCQl6evI0+lvV7uLV3C8fP/Kt+MmSauWp5REbsCKgNqedZ1KsUNa/YSD2N2Az9JmRG
0MfnKAgUTMRH6rysz/JK18vRP66qVO9KP3iUelp1gGIsPFVNmjDeGF8E/89itF+0d30Y/hNNLR/y
/p9xA7FxW4L3ZtgFDdyDzWDj3pv9YfFQGwIr6yv6XkDf/jUcY/1cayd+sG3QH5l+k4xukIvVE58T
lGL2k0fPYn2X9IN+r41tdvwzGc3pXrRZ+bFfmqqeuBDebRG1WIhngVWwvCuAO8X7qt1Vjd8/jneY
HRIXAtc/fvHqQ4QXk6IbzB3BxSzZqt/WlwCCRArD4yht2aCyaaZfkEAOX/x3NMrryoypeUkRCAk9
m6MVZrMI0uIMkBLQbBaVglm46V9p1SrGowCoPwR2paSe5DeNn7P6NwNaQJllwnXZhfNzxrzU2Qo/
0FmSA9vNKXhbAbfPiltZRxfWlDx12WmBksyIgMRcbpGMSp9Qh4lqsDV9f2RNLFElGxdr/5Do9vmA
dSeXfb56td6vssYGS/Crc/B5MfixzcSAfuRNm25sLO0vqhBd5WTKHHn2ITYeNaA2Nk37ozSRCJHa
KAHuvtxsbojdIsmrmlnIKcw/qOejtQkHP7RkKfN2/BsbaFieT7RoOY06GwhEWUL23IlYpIGybd8L
LVnDnEGB4hr2pohEX2bEpu/i44zkSlYOelP8OCZyAf6qmOoeG2PnxBBz3uKsOSLQsxdUQ6XyUIdQ
Lhp8zVbzTMjLZtX767vXNjW9v/iS5DRXTMQC8TqLInXBSJIFK1+MS9YfOLXUW2JBUN4YObHEi+q3
dKC7ktU/adOZjsqnVfAc87kLPC+7wfHnkKLCIf8IQwmet3a5pE8psQ5yreV6G0bwe4/3qEUnnKq+
wjuk0D/ol8qyzorjQ+FTJGS07/UuJp4QBLA0rdLwqCPGoOsKou9L06a1/v/W826YzfdrmGoCuYHV
X/cfZZDy2z2nl2/MFeEeMu+yVcxZjg7dVZXsMeXdBQMxr0mHqIjpClvm3LOlwxCm4b09FCZIdcek
9wAPDrfAUKqZZdlmcnXucS6xXDufJswl0rbozUIHvKEs3hnQmlVRDtut5cppLRtDAjUEgO6TbJXI
X/nH8lw1fKYdXkK079l9V3+edOpm6zPw0WBNAkVf7p4VNzdTlZ9IcV61/Not3r7UVqWP+MfIkfU4
oNH8byTW7/7ILVM22wxb8t4tBJlrtDbAZP2uOVOGF2mKCwbsq2ML4TJFmnfnR3QAOzCqGrND2PUX
MiCOLp3lU9/VWiyzzHcFuNVOD6zRvy6lCFTmRPjAqD3jnm9RmeLjOEwId5R742LQBnQQMWzqI3R0
Fv6XynFvqe0b2FSL1Is/Ul1lYtmTtJ7E5888JSPlOQymK9gSZKcUI0qiiuC1MsK5T3Qx36YXGDGQ
l5X5RSsVHbd1Tnm5wzn9kD8XTkKrb53UO9xSza6B+q5oPqmJjbygx3WJCqrA5Qm2snEGv+MpgTIy
SqOsH4rgSQVZAzTrj5UpnqVHIu8Rw3+3fjS4U5W3kvR4fn/zHLLTxbPWpdU3rcNbQGKpsZdFeCg4
SmmmW93tSUqX6Rt9ldVFVG/M1DhCOSzwI4j9/RPFtseutR8Ba5Knqwv5N/P3HAlN4YWYQvrg5wJw
9iGXvl9X8msWIUfZvVkMWSPTN/h9VJNusHFPXShz9jH46jbz/RR76AzmaiipG0eoTzf0CdoYx8SJ
fMWvQiCYG9RsSN4ibM9ctg3R0wDr2VLVhh+wU7GD38Nnl2POwSyD6zn+XKvU47lrvGoBw6IsJxiZ
O9raIRNoOdfD0RZS3I2alid6t2Opb+ps2JHUAsLfkMBv1sa/egp+aFZYKuTDw6OUnDVPwnFomO91
X9mpvMO36/z11xoS8DHeJfsXrL6lwe4rMBZU6XCWOcu11/NbtuylS615LTeAdcvg6eZJelHo11mB
akgPvbeGIGWEbzvcYNftjb7FEMAa+xSDKoR2eSH3/ovCYoAtPx2ViShlYuLQrK5gF2a8ps1tomtk
glUqUdXYlgumIlFXpRJUjNly2T5pO7ExN0PC5GfkocuUSG1zCDXW5qyVp9NAESj4p/8BC+73ee2r
XeLi3tvOJMgaw6wk8hp3knyXH5qRVg7y7XdYjiCYEFmZIaJo7Dl14uLnECWfDy3uGSWdsQ2GEehj
G4MW2iXkWwpy9qVjLnwR0Qf5ronuOdnmsDI3386nCH/p6VFyxI62sGWYP5/kggk+8GgPUQ395On+
APc4f3F+I8kwNOwD6NNZzW2hGDn+XW7QaZ7qJUYu1qvUSeON3y/ZCrgpIBe6/U7rtp+7aHyOb3YA
NqrUsimMXZ6ydLhetO5EagQCe4ry9E8T3wlKoYsNy8dlmwrkd5/pp+oAuz42mlldlYSghBZVP1mB
mh/rWn4WCgXrz4dc8kcYAcGqSOzNY7X1/lL9ef+dyaqHLpKeVoAqXtNsHHCkHSs9TXLoyj9IgY5c
j7v29T9OYrxVL62SV+x2HzGCixpjIg6bPHkooVdkobl8kE846F/J/cIPju7/hpoY3bjEs9OZ1yQb
EjiX7xJWuQw7F/fXKozzhuPNjRxb3b3pQfaqSI3OL9dnGQbrXRRXVTf6qJtE+gfpMXeUQU0Ushdm
9v7mZnrzA+ZpL8o8A4VQfdEaqeTg42vIDwvHTnfWZqLq0VmAn3TGFm8qOB/GMvs2Ir4fNiDbe+1S
IQkmLTVp6PbTC6vG9MffCmqywiswJptDKHrMyVg4Agphn5IxGYQogNO7Ay8hvB7p8qonn7BYQuun
BZiG3jDeJqUZdtcihs2F/+jQ5+lii8E3RY+avWViJnnCpefHBd8FsdQPL0PFc1N6fTETkpOg/dw/
qYZ7a03PvBj2FTeFwkpgcETUyudD63pzGB8Zp+rotQIZfvkTyTQaI2YehqtquiWaCngb/pSgaVoH
Zss29QLPSs3X1rg4nDO1VeTwEzKSXPCrm0SNg8elqeo4sDOIZoY/pslvEpKdm9dbuI7xWSo5D3vj
TfpOcf6TPRCSKuwhdWtgCvCMVe0potFAuoVvw4VDdUOw/F1MvjakX5rf71QitJN9n4CCfJnsVLyN
ILhoeuy5rfBWpP7++DWg2ddUyBcbkPB8HMO8z6CPhW9bAudpxvcVDW86X2uPma9atmS802PAvs/A
JifPCQYmXWyiJG20CNHjc/QAK6gTtKU2QRB7JmLqF6dNIprlE6uTwsbDHnMXc3yOQEK9LtLW15Vd
xOIjBfFJyYJvEZooZAAHvAZk4iP5KrciYC9QmuMe12GjbPCcLUqtL8YYn+VZ2DjuS3/QJAM7SCmG
Hn4iWe3U/2fzWXB6KToLUJ+PrG3QmGm/DiLTMlVE2XyU//wr8jEyo5DhD24xAqeH3FWVfmsQXKv0
UkO9fHX7O5joaRx5Q4uZHJqf6is1MFpyWIT3q29tnFik7WoQTtYSIuz9tId2gwYFuvA0+XHmbxqj
eYeWB0cblaY1Y6aD4C7VQY6Ya8nhr3v1NYTE1BlLpTd//Vwe+CW7Gik9H7kbxnkaJQm+F2qaMuxB
2aEET+TGttTgtPcbvNtRuWUeec0zmnaE1kw0Kevehlsg/hSxeUtomLCsgV8IhqsyMArnz1ANjbcz
RSAdSDqWt01N7ZPNJshhE3Ensbvvu03/ds1iy5EYLxDJBNrPr8hrurBUqVqbsDgb23wpnqXEtlms
1Jm5r1g7MzURSSJqcPejlQVLTscNlW0xSYJ/oDsV8Y6zPKW6AZSpSb798Qe1zrQhi7G+eYb6gyr5
YFJZGx8DKBy2OySQcvZCqbDWx6iWh+Q3RG0aW0rNrEWlRAgJ6qYEHXY6E8Mp5Sa65xB4y+MRCsXL
jOVWs/LPm/FiKquHJbwosM62xjhd1thdeEMfHnAVPv/nfOFBl+ES8QuPtyigLByt82QH17CZV6IA
JxYTozJDiMVbCAheUHM9NQYQ2mG1qq9kvqgAy58q6JKjI1XpAGSXRDNUdTPP3lz94Nvm7qEPE1Zm
r6FCxMX3a633nOE7r7uy3509tox33azPmxu0xcdMwn1UjJgoZ8AoQM6iEE5+Yt2IUzEdK1A50OeP
n/g/Lf8kDVfkA0aJsjMrmZsYrLQkDo+m6YBmsZEOKzIF52qMteUJ6dtpS4x0c2HW4bp5lEOlscyp
hv6W+6gOfk3u6fSOt0XW91Y0/aJ4eUX01We0Qt3rXlkYeGdnsO+7min2y3kFN90yBFZ4tF1ITs9f
KTXmbVZ1QShgm3sprJeJLRHHOsHQprZdEwTiV2U3H9WOp7hXTWIrl3TPPGNYDhgTIlsQ0J6p1J3e
2LCHMEf1GugdtHlj6iY9567QQDMoOmTJt+PGUDm1cG/0LccxHlim8c8o1hluny4+uddTZwdNarU+
nLpblHEM9L1QHkgt6/wKOfsLwabEWPP7Z2QCn//8ZVu7uwNlMWYrOI0K1QsX8XYSSPKV0NIkGIrL
mKtd0Ub7YExR1+8WGayL/qg2U5nLbvL4q9YPeIdIEa4Pn9VULUzn09EJGYRaFY2CMKqq0lU9f8aE
FoLUHj1U0rUndnJVlDi4jh7vIcznWPlFrrNFlXB5p+IpK1PVekW1xJas8QtvcD5PK8aT4h3rAybv
oZVe+JvCvCwnPfdLq8mK5oIPM7M/GxPDAWbu6UnsISjNkA2cGBuBiUn3k9SDKFwx7Nn5ndSNERzZ
2CfkOdNH2Pg5DyYUv+Ocn33vZefl+RDpN1U6LTmSASdehnYDIQraNA9NKypRBf5VtkBoOlg9cTwE
osMcbSe7e6ESN+S96almysM+Y7fMf/6NO1jgmyzj+vEUYqmInoHUXUL8zj33un4MgKxjyhe3+ceG
4Pa87OSazvWFYddKxWF7u2H+z9i2Nv8Sm0S+IB45tRByRzQr+8yx5Hh85jx7KT4+cWNnW4D1n3DN
QWs0jt1mQ86eDSnRNxxKKmcw/EdzEs4YUAyoivjslgRabVj1VxdXaOh7sg7Ms4j+lDanGwJDdtrF
ooZz/nFLl5IYMOJXOz+7l+pfnXOPuH3uXkklEM2hPH/5voA7mI3qiv7SmmCOKTiSG63xXJBlwFrX
b8f8Nt66NkLJR2BKOIJAC1qpE4jUT0BF4Qc5vPmlsZw48OD2/AwEnk73D8zWajQ3gr0CA2f9XuDJ
5lXygGQ1mmtejY4gM+Vyl8bP842r1n+brN7VG6AX2cED2YJHnY9hnnLp0mYy60KmhItUvvMd7ghq
6mjKnypd75GkYQlAfbVcMwUXb30Psn92Uy6kDGbUwnV3sBY5yJAGBjHboo8UEn/gcWcKDw3vDp1Q
q7V06aYzMMCGpEtXorCGGjFHDBnTuClGC4kcXVbw419PcdgRi3mj2H158xLcNWTwyh2pzeoytWy4
kQEdgSr5zKy+peBj0xKYz6YSbvL3471t+778EqY5x6xBUroRQAoB6X8/u4Hio5AHyIi7LzRltZsw
tp+cvBx+1wBK0V/1wKa7BB+XE6D+wWPfHlACRKfH4q7/bbFEdeAFkV2MKUQz6VkXoAIgfxtolzjC
Vf2aBAL9OH51+/QTQ/vLe3kaY5qBfi0nQE5rKRiJudgDcJyVzPurNyjQ5xUsixgkpJLTz9D51Nyu
ayHDGNpX5agsaS6shC3Cc5xhD/vSu1JcOU5qSdz9/Jy1qUlJAjbOpvQ6ZGl+eCXLAznlDrZzuSly
zjFQUOcuHgOLgPHBxuH8avUR4O23zOiFpNOhE23AO4OovdBauMbJ1tVY+ntVartnFZ6R8B7JXRur
LVxRRQhgodgJ6RZiyX3M4g6p1eGJo/nlz4zrkFtwNu3v2IGf4o8Cd6LUGYzXPB+wJHUhl1L0Fc1B
v1dz+0LOfEcvTSMFWFj3wfnrLMQFC51kIfX/QRhbj2s5z47wGPWeNCtWImed3B3cfXtwhYIfnUHa
PGRriqL3LAlk0PrP8i0blC6b5+nMCnm0exNg26HNb6KzGvYtHZ5kUELl2R50TY5K/GL+Do22OwQ9
xbOOL3AnAuiGdy13Uxil+XrSez/NGPJ4ERq6nUDAW8/Dmb3Q4aQQKkLH7GGWJZpab7PyaTLRMLyU
v03/0dY2dGl0hPUUE7wjtDek91InSWkMtktT5f0BPMCW80s1ff5Trtl7cP+mDw5QbJA4OCh7u8c2
LclRqat59xKBygdGltaMHXbrhPHwx3mFgjSnnUIv2u/LgKJC1ksxI5T2ehRMvKAMKrAdxKKywXrS
zWlZt+2iOcQCkdbKew7KLolXmKiRtkaH5Mu+nYX1M1jOmjPdN+QZauCIqljQZgoKxafDcFMHxPmx
CJzkADbxFWI2HyDy/EwDyUa3NJ2mYcJuVpF8UI6FuPo1Gn/aAq5LMMqBVx2NCocHlIhTU/2hYZDZ
hfTymVBcBh7hJ4sEV4ObM9kRbcj2vPCGyomxgb5jBxnQ9qr1J96U0ZOdE7zi9si6W8093s8OWl8a
U3Ajhyx4ruLuo/10Pn3Bo3zSc5P2OFpwB2+VNpYFKl1x1cQ5b2kHrN+aXsHca9HUtq9oG7jCGpXp
2NC1ehZjdlZW/9FHs2J0IZkVQud8jufEiy6dbVGvL8DRNJNoylfwqDSsUaGtXsFkj9rcfaRaVTTI
+qIbNgTcM2qvqbRz6YlbSwQIIZFn2Z+9tsHkcWCce78mHqlGvIlYiW9SqXIYUCGAWyzIUDII4qM/
4Ud3lQJd1nm2QWsNkod0y0UuGcV4tlStxq7eKUkb8Qmm0sTCq/g2IgWAtVrs3ek0oG9upaUWFlwK
wO1PtOE9FEaosn7ZlA5s3DTHsNuHFRUgUvwf+1SVu/Dxv0yig+fVFQAuti9Y90ix3g4+skUAvwzY
2yvjjHW6JixdK04m4cYhUJeH1VLDkoZTsCHYSZ9Hq3y/g+nqwhNLhWMVfmq8XSTMQoy0ASEbMDi2
ABdC/SwpvTL+eic2UYMlAcba1fulsk6OJOSlFOBD66mQrtN7lfGjLP/SwqEBWvV0DAW+lNmbymJ0
dZCK6+Qs+wWTIoOwprbcykPNqisu69qc9Z4UcXQ/BElXUgQBM3+Mgu1XDgR5W0uhDdQx3XhjCBZp
GN1QuRSlb4tlrkHRqRQn6gs6t6ZgXs6gaQ+Tl1rTom4W/wLbynaXq3IULeEv2p2zSuY+3NYVh1Ye
YFQODWl4JJJkwbp5lRzrKDaEMrZn91aRzX+cf2003vSVAHuezZBk6Qy5GFCpdVsQfbds81gIP6kZ
x0DtEIRJyWaEYhIOpqndgypdFfXwpIhBrOBE1dOxiU8LOaDzmStMMNZstUjCxGxz5SpJLGBdCgbi
gTBZntiY4uGpGSIDbDebdRJxx12PeipqC8NV7/LVpHJQxvT6246D8Q9Ru48LRtbFVAvxJ/WNOBmp
Im7nHCrtdNGKg44gY+CAveUOIYpUWIHNtN585zLId6XXa+BEq6Aras2kgDCcGvZjfgw5JLsG9iFI
O6X4VKOPuXDTm7k4jPjGW67JgZKm8OHKi2+DoIH6bejuq+Y9YWdUaQZYUpsv8zwiWYlkcjJwyVeZ
gCKSf/QLEmCLSmzn/Gv0iJEGefdfBiYq9Z2hL179OzXkzcT5mLSfxkNY+K+bd/l9L1LsQdub2bGC
nTKu00ivzxZAdCanblMx5cVhw9ZGVbBGwjCicM05kNEITZ7YoUrykPsngqUNLFIbXgmkvShzNHSN
VBeX6oJ3uu3P+TkZ9jsVkFZIpPUgiav03HH2apRF2zvkYqttvDOPUU1KGy51yWNzWDfMrNDZvqhm
Mxj5UyZFhN8pV+9AyArQdgiXE2AnpjMWuS64WIVj81cddeh5ZpjywOlCa+/+sfixoGdnm86Ifkd9
BkJttsJsCXXvKoPKzmFJHUjoBUcIB/z7cXvei/AJkvoI7nAqSFfHNHsZ15onsGNmTpdteH4M4Hbe
jr5cO0UXnx1LAhE0HRHyRrG1VZNsc2vn1r/AO4DE60jf2nIhYf6Ql1VoKoVv7CHPtw52nymP+d3q
iRVZXtLN54bL1I6EMULTXj66pj3MHB5Bcs50Q0MFl5WaCKuIrkv+AM3UziER9/x9ZDIgvoDdSmfo
FTglQ9H/jIF+A3fO+qlPaC8LzgOqZMIbcwNV6yx+YyMPxNzqilipCCEo0ojzNxHkN9HIBCrdHqU5
0937jo6dxEsJ/iabV4748wb2ZXm8wkEBoDeodrKhm1IGI16YGbD8MMBdxj/qkh2ejpiZsNBJdJZc
APnVx48miGHtLY3MewfP2qWnD/teHlJQlvqOYXLkXgOjC4utxaby63JlcIrnhmGHqMnO09XuQRQI
l2iDc7D0gcgoQK8EppjRGVJV5WHAjocerb2Yd4Lbl1ueXBabxkU1mV2hVyQ3HcE7YGWxOB5AZ6pp
N0g1nJhPCzEAAp5DolcDisWeHLKZWxDKWQ+a6C9N9qxL+8wyK1+pUXdTS+6NIJOIKpe/qhRDpsRO
7pVNMmDoNJnMuxzP51MYh8pwpIB9AYPqcBY11SS39xjGEbNCtx08zEVnDgK3AUBSZumCakOE7P7A
onzr1TeqGm2SVVmuYuW6JI1p4iCn+5miSHKVX3zeHOsTcbWS0lwDTMiaWnNobIpm5IYy7VMdRi9f
phmQZ4kBoKswAntoDwpwZuTks5+dgDBeReP9VdKDjHgg+74d42AXpyid32Vv/mtB/ZVY74I64Cdk
vd9fECUuTJKSX47YoMAk4KEo6/7BBfndmcm02gGtjTMAw2AS4K19pVx3eT+4wUzrxOxh/iL4vK6M
71bmK2MVhJ91E60ZYtoL2e8sya8FZO/+kYYRiJrHOxT3kdYi+q/rdr7yXwJVOidep7nuJJhNdUql
+X+uAwG47/7e4aXZ5Pay12H/XlXXje1H4sUpmr7hzLNGgkLqkXLE+K2efz5k2Rd+FANXP+TxWcW7
Cc1hcs7N1V8tVIO5cAq3c83NYeutSz1wiOFMFPA+pcibSAeZ6iBiDtBfM6u3ADJhXmpJ4o/QFf+P
6EZE4eACaq9WqxmhSQIwlDzGKHUok7WGGhpZulR+mMkJXO99Yr7ZACmii7nfZmPQcu3stity7mZQ
3GrRv3q4uZerzIINiU6UkXHAAhfjQDPNdxCEJ6p7Q9mTS/PCglULR73uVcng0HcQyUXrlYpxlDmW
caZxhT2ia1kvlpYcLMD1kU0Yx2l53VMBt5Dn5ZhO627MoXx5ucb1aXaU2U63KY+U5V0E/gtKui3+
c1OVBSl0YeJBED5LseXG7tT7Q96hw3sglJQ1VlplKDQXzXdh6IP1hyINFfgJK2fCj8fvu4RnmxYC
qVXTFCT+CGY1zoeuFFv6WMQMn2os3SE97LX0Ujzxe2nxOTvEaNv5ewEed7cCxNvwkEqqcJ8BBFPr
nnoP8HjNKvLDbt4+Nt2s2utv82ajrPS12XPQFMn2WRXcDrbPRqBVGCkt74HxUczGBeL0sgghh9Pv
WvmAfQluA2NqCPeY327IwuiWEdaddWr8v/CFRR08LS/y+zFzpQawp3y+DxnqqzdT008tXIZhVhTz
6Lh9w7BvloZ+/L9vkHxbYMKE5hDIRM5IPL4RObv37XhJ5XMx0d+QD1foJ/FY5hJ7mdaWwgUt6VMr
1ZYVSWlci7T1tOTwS8TetlY96DpfXJkA8PbkoYbK5OY6xBJs+pAMqW0JRklLHIsb72RXquzcaFYM
O47UD8CnqSb4N8fcd3dC/Gl1Q1rcWGEI6YcX5X6I51Rxf/72Cbw/sIAmZWy+n99cRkNlLnDEm3yQ
cN5/IRTQfG3xtvYFULu/fhIy5gw8YLP4VIFDNhIvdUtMiuKuDaSvSRfLccktPTprpFvO43bWa6wV
hNN7hwrF8Mk8iC2lWUE3J64vw0bLsTiIQIT+DRDGttJtUx0/VCkQ/XT/AvtS0P4apDx/gl5QS0vs
QEuVHyaCjNpJpMpU4vEEXVzehMBBCAjZ94Ey5DEKBcHwcdcSqxomm6LjgIhbvGHvt0wrBESKvM4m
HYDv91gitnINTwWr8053+Opksg+JTfXRfCgShfO7YK/cg/5UanNtQYSBEzOGncXb3KXjxeX+Q9WD
JuCfdZiuHnxFlZBa8dtNMhP2M1nw/pSEsZ59BZ4pY8kgdRoRxkQUdfCm85af6KdCWXerHQhlhmga
+XRAwvfZYbxtO5NIsys+VWBucYqqE5RJlvz5Y3P5vhso1tG+TuquQ5aeyOXJu/2p1h15xGL+RzWv
7OxPC8P9a3OAjI8/77as0lY2YlLBZxyqsTl7QraShmB/V9PESw1Pc7SyeX3cRs7Dgcg2T/ZH4e9w
LIdOO3jqCC1TPEGTq1vjxWuRJ+3QioBZODSkpsZq/ugnz6RBSvQ2OPYGYWkeBf1+utsSyrgj2KEL
NgmJdSZXQk2RU9oAIx5uKFa+JV21wcTGihXSyROvKm09ui/hcCwBmDLyxL+mnlbd+jO+4nGGtplo
qSoroIGe14YQhXGNO4p4VO4w0Lqr52O+23sUpX08KwnmNw402opikf+4AzeGDFdsZwBk9KVAEgOU
rBGACprK1i1vVuXu2uy7TscvBEiuSuqXUKel8bYmNiCgBnjpNU9X3jQuwimQ+xBc7v53YNNq7+Aw
118C4ABUtToOVk/sqVS3wSdE54EbBEaIpSBTfaAxyOFJYPI0z5zmlFQ0FuB58U/jqXdQgibJASLD
LC71D/msXYR/kwrAwa84C9FlbDfNg19EPBKVJJt5Hlh9FS+XoKLM1TLhptxJN0zcQIkWh2kzhL6M
nPiZ5ZclunLIA94xnLm03BVTlSo6HP+O4PnOBVRqrklkDLRSeo+EN2+6+NWMjbwaFMiqHmc+3PT8
2swDUyqHUhlSeB/EV8JB1BdL33x+aF0oa0ig5op+ns1bSKhGVxkNq4WCPfndWAMMgvmcqyUMorhH
IejJJsUoMEh/jYByq325RZa2Jj+MwUC7mxLYvk145MVWH2V9R2pgTM3X5DD4suR/1JF/nhqWEUrk
UylMZ1i5FXOZCqW7LcEuSiG/QRKssTDH2XNHnzGSLmsQhKEVrekqEm3m7aLdunJ+sK4eYidmsNfS
XAIFr/Ajn2FJJYlGHFIdy9gTU5t4JxrdrIs5f46PkoWqY+Ndn/3vR8tI12jwwKfsLieYBrZ69uaO
b+7OLa6hZYqUxUY9H7njBKzvd+Fei7AaqMMObpClycLIQjI6A7J/5XqWvRmHDHEMYSKmu2WpnvR0
9bWHBZokgI9tKDX0hNxsx9DKUc+Kl2wsNIs/j4aHYTvcTy8y8eIhP2V9RTc/J/5Lss5cfzKEavkA
t38gpkw9XkE+GfRxM7On2CMpBe38FqLfcagSASYmaMfDnYNQNpiAAFBP0Zsp5O+prWlXBAN3EWWy
RWVnBngHBjKcotjPOnELWJIvCE25aqAIFsCRECADDIVR0pJyRI/60R1xFuCeANPyttU6L3GSgER1
mTlwExlXdAw2/4dPm2EWANiN22PP9BbbnDhSt9rExshxqFswY/ZIjbCm7z1tQsbS5F7g0MIkGmjo
6SBRrSrrBQfH6a7Fp1MZHmTFU++uwUL+P7vVlH0rjS677JMYYZH8Y5HrFWEeKTp/Khluxok0136p
vJVHxjltl+zc1lPDcAEFWLzv4S47jnASOxbNxljPJ5Bc9hv4YcQ8+SLbbpJYrmoUIOmY/4apzhNv
FlBG15h3pWfSKtwnGRhbX8Ic08KYJaTdZqT0aU1JRaB9cQUCgVUDOLDrCR9fH3U1z/Fe7LoZ+cYf
ODa+0VOhcpBJZQ33SDxKou5xJQnLWSBs0KUxb0j9+gyu/rj0o8A232NHZFOpCKLVhGDaH4pJhvTH
BD+6dC2eIP28QzpELxpF4zQD0+Dm4CrSpBJw9L6AyocyeJxuJfZb2XQjUURaD2ywPEUCF8pb/ZZa
W6UVEeZBWXBjyX2E+sAxU3shPrj26h2UjZGFTniMQ1z34PxwJImYpFDph5w13rC68brSsfcDTJC3
r8DnlzAz9H4CTl+9vd4bO0luzsSX6HqJbbAMS6kZ+Jo8Cdko/+jCs3uF4GTrp7vKB0aGGmS3r+mw
aFD1Wvm0lYZJ1xaYuvz9Vbvcplx6LnD3KRepMPKxnpGlBeG0iKfGRRvhlyLvZTbnKB/BUEFB0SYW
zVnG1pUaRQnd+ghAqhclpn2OYpi6ViY1SkANQoSkxJt+te7apFKA/UUyDGR0ZbjldMyqLH/mVfP5
H0o3f69RP45tJFhoE6CYvXa/5ZB00gQrQwrQf8wBhIWh2N/OpPV1t5tAB1hxIyv9CyYfl9RA6wy4
Tb5eIhDWwl1MJgSVlRdecbwnQcn6knPsPoFYFTbXf2OAPUCquouCYGRTXVs5cXJHSKTxBDGTD789
5+zF1CgxghB0/xqnQTw79RyG4FaF36N/7V9AJwPBx+SnsAwjswCDdf8/0GDvdVv7xKJ7QJkRDZkH
3gs3sbnSV3BhgQkvE6Vl9H2s1RSKaXP/4JuZIhDA1511jzhJBsMLimc4Sci8t//ZubHkEEPhmUeL
i9jqTIxN8etFXb8lpylm9wwaNaGRuPoDt/szMcnPx1c4zkS+E+Xt6SsMkoKscvgD6jHFG4iaX2dA
32j+8KbDa8Xu+rNOsu8IIAwf8xkLgeVooEQJCsBtixJOVmwJO+xDgAq1awQf/NRb1XHGfN3eIT4q
/33tZ467VP9gRDTCMkJE6NS2H4HG8mfeUnnH8wpH4fvAN2Lgkw9sXGCtnlHb0SJBjCOGun64UYa1
MHLdRMjtW8Jet/uaoidUTMsUpBlsikUmsrp8rz5Nci8181dSGqKV4Zjc39+o9xVSwjEDA2AKO/HK
wAYXktxYZ4Racg9ciqeXNHEe8FK2QFNPLwWvBOyOrh4M0IGIi3iFp8DrYp+uEsumEcRJ903h2Olt
NORuphyaoA53/kRfAlcOjZmsvrnK+CM4tHLCdLyu0qthT8AZq5ensurKthEj9mdqouGslvFX45ec
QW31E/jMn3OSrrOU3PTs5G+xj4Zr6eBI1RmI3l6YhIAiQBSGNpWp1wR+bYlOxWcnsnak95vH5wo9
KoJMwNbSbglmFXOABenusujTWam2h52LckvQF1MmG6iKstTsf4m7JBWcppUXnuJmNni7IA+ZqId+
2vcejLP0n2wJ6hpXI9HAbVoB0EMpO/W8DJOlL4aJfNtJ7yIWwLZzRSh2ga4dyE5aNekjcrgnfwMj
AcWa1YXdTGXVAGMBtmuGI5M3nbT13uqdWF9MTRXcPU8TeP8Ee8dm+50sEOuXprRUa5P0aGkyAgoc
8QObNhhuTDfOgwwXkrBLXSa5qalKxEA3dtaTARdCJnGIjW8DqN370uJr5IjaqASHfpyUoG3XCMZv
GsYLbTPtmwqesLJlkPQSkJErv4hWf57CSZpSCouIc7YNbZCyzH/7RMJ7Odb7s7/JOqA4PlhDBykK
ZW4ChtWTkF/JL4hc/YFgLGw3zeRVN1opKEDPdKsCP37xsSqMd9xaHlo/QIy7CCkJyDsjeZ7ZBWX7
3DOAGYAPXXxVwdMuSSgy+QP3QcUKSu+OxFToTniJdzPCBRPzco/TYwFUTDFAEoJpGJwmfIF1HtWG
Wj6/vnJQlAd52pjPKG04fqVYAVzeNvkcqgU4/eJKfJil26jHIvq1y19E7yeHy4G+9mkLsG9uO6mN
fgGJb96ExvrEecgCZmnIaj909NuxsnwIdaZpl4GVoSEK6bzSxNnnpnSoyCPkvh3TqPD/vmLeaMnZ
y/JerMcb9ik7w8iO8/nqIbwk1wbuwowSJ68AEj070to9DAJ6xSo7o7+7ulCgRvuCtt2p3ND7LDoa
uH48fD6W9vvIhRm5nGGDZYTkrILgbawKZLwRQ+rZOyXAstOPtvy2N5Bih+zngSa21PSPy+WJifcC
Tr65JjlSMVcN+FUiuxjwGk/rF9HdH5eUg8x524RFxxkQdw4d4RRLgP6WveDxKtA/juF6MVtYPOox
mQEdr6MdpB8u8NlfDizLuIrYAWQBPSIXBTCP+JMD1Q7OE0Enf7HibFjd+D/FqaBzX0vx1Q8bUuik
afnVFMuS3BCHmdoMDq36+577sXvApQjY1su7GDU2H38iwVtVznZltVViw55r/DkMcp096nrYjKep
stwf25HzVp1Jd0w4wbCqt6BG3yAbIoT2aOMni5UCrKduJezgC1v33+DCvQ7mSCpKXipftaA/OF9I
mKOS8NRwkhT6RYsZKgNBOdMlb/SRRqGNdOfs2CHJh4ts/NMB7RZHlII/OdRvP16rdZrGO3bS0GJq
a6+UzRmweZMvI3AnXnmC0Ec47J5vLOX7NE0xq5O1yjy6nzzwYL+HMtXBDr7SsXioyAYYPKzjD2XV
c6Rs6UeqygHqC2CSW8t8wavMUX6cX85yzRwhOqyTgH36GIddS/CGhC6W0JwyIrcEbMaThXmtu/f9
Y6DORGfvisjBwnKN2o/Qa5OqFvusrui4BPBNNE6GxRF/UCWuevqpj29yg1g3y67hHeZQJk/SRKDk
Yr7VEPEip1g3Yrh1ucAUk0JisgJYG2aavl41rDQcU1DcP3TExgMFqoCVM7QZ1yI332NRAsC+osJz
wFcUIUbDH380gRE4JKfNPKaxoae5bZMgVDXQiKklO4x+UcuE3rfrMsZytFFSofDT8gNRytykvETk
QVzzfN802V3fLVR5Wjbk4w6xCjCQxvSOB1PuYKqCmbxnSTUv2BTd9+AitTahVSZRAMuDTJGlo0sh
g6+TXhB6dhDdnsZ2OqefbTffUaJSOHjdZPBVXYw2LsId8V8y7BathweAPDyW0VZJXAlbHQCz0VHG
s+z+eKTCFztbLquxpYerWyC4uETHlvDyKE8Vq2Y0VhKF9iuaMOO6XV8DmE2GAmFRiX7qoE2EJ03J
s2KNgx7viZfi/Cx8DMXMLe890Kb1y8h26N3lAOUDK6VNPZyxGcJgaCXGkW5F4568/yWUQJiEpQFa
e4XIhuArQaDgNcGUuT7mueTB1Eg0oqwO98mcVZXKbd5wrfm06t0QhrunLexe3yw2bBuHw2LAw8py
7ie6FlRaLJXbBl9TMU3YAQkessY72c29iIIrfhlupwW+z4F+xNoQJjBMtz8+jyEHnqnpGnMFMRuQ
h5dlFZOGOAPSsTYb+79+yaWUoiKwhoYLAWh9jd4SUdpdHQHqViWaJqVbHLSDw6lTFPE3FdbI5DCZ
S0Y70lpq6YzNhoRmh7xkiZUsqq3PLJJwgISvserggDFcOpdp63dRM/Dzn6EmuPTG57zsZ/np9Zkk
7ECnOIpcsY5iyC1ILn+sqcOrtAdutZpG9cXzIdRKOpuiCU4WVHg3b3QcqrOZtAgiBwcljMBRZ7wD
7+xXLFHoxdC/k7DHta6LCa59rQBcDETcvdj9wColtrEn45rIsWirZnWmHyQnnVNaoZ36GWbUEyhx
5KuaKdn7qwIvNwfTcwjVeCMkITcBVAaxLutZcbENEd9TyRmzpxUlzBnK26Mf+ufx
`protect end_protected

