

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
MxpeY9fwU4EddFSpExWohS5o9i8UPinR6kQv/f7rVpVjW9v1XPHFNv5NQBBqnxbGk/3GroOhKYHi
zeZXd9sb8Q==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
genV68U/jEyVif/FXdfTRcDdNLXMaB4JkzDnEPHISJLebDAxHBqab4xQb3vzSMzS4EZxJxM3czS7
l6/Pa+/lUNH4iHFgH3/d34ImoXy9UrVsNWI4O1k56f8CO5JZkX0ENM2JUr2+jZNnrmepHCpz3pyr
N2xknPLUPWomWT5p45Y=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
4dyOi6X0ND7jxJKLfQYpMzBQUnXRUvqhIlWd2qdz2OgGY9VUivCAp2239OkMu2rIWSpkdV3gd8Tn
4E+XnpveIi4nHAn1AdqR2yW6qJRqYI/CpvcG8E7ZhuUiWSAPiQ/jcxRmeyzLFdVhgEV4hed5vk+9
Qi0C1DUHqDNPvc06f+xZUSTzBSqXkxyUqGIa+j3ZmCrjq04hmRDILUEkjqmR0K0TOLNdsLd81gAl
LqIfeuzK3hLcVWnnJG54RzS/q6bahPN8UaYhtJREcAC9BD1S+QEdDXRxFczj2T1LQBL5rSryR8bI
LV6YqNl+85SCCMZmZV8Io9S7fDVIrhzNm4Kcmw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
PIdLn+S6alHzFt/ir7zZvMPdMeYQTL6BrWSuIGxsOazGugSdn7m2jtyII74LXXAGUQ0h11spxnUf
W/HpoHHxg6pfmAZclwmfvLsFiVi0w0hNMmIWoR8TGPdAC93Y5+aRfoAJNuDfUDfLzdBM4O7G2ZFx
YGYpvBcNhzcFFuSCCK4=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
KkGw0OOEdMUjhZKEmICwPPGTbEeQxk+K4HH0ah7Z5cm5dbbyDDJyn1CdBy6WY7ZD/SXDbXp0Ibi6
BH7Y9BzUsE3rhTUVWQo0OMHXc+hE0CnmrdIq6Yy3Wkf73IKl+pu+66Qo9W7SdJGNPpreGME4X4AM
zBwAv9xByRwGoY45EIIGTaE7VL15piKgLihjK8Y2Ee8q921qHsI62b9osdj+stH9M0nIgGIwpsIA
DiUOa8Naw0kRMS8QCXDqKr1fJ0jPj3cnclvP9Taz8J5tp8Sf8I6bs8irg+MGD1MgQIfeKkimA5VH
MerNz8gbn3+/Vz2X2+nKanM3LebAMLyCO8EBfA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 35024)
`protect data_block
K/Wj2WsLOmBkFcDpZsad4JnPAyhvLQWUIecCEmLvLJ9Y5OXun2WTIyTw6dmuUvkPvrt6vn+xMw8P
1jnxyfJSkSvxlmEBnvRJLhIa8Al7uUb4fbXigMkfkPE9XcTcLLo2yGjwy73fOb5e1BztOM04Azzb
Zx5dvBuhiznsmA27o6Qq/OooLNotCm5HvXRtj9Ke7UAnPMK8PIVpQZUcH5rM4EifpRCI3RgIlOir
8SvZ9VsnsAERoZxYDC9zDSHsVZo2ZadOsHOKOBc4YfyANZpcoFa726NL8h6nhR4/JZgOBvNfvSDt
+MEE5JERxli4QfRVS9+FNstB+8zl4KZDQZ6kia9iThDjaQuULV6h18eyzcyhICuXa7CdHRXCr0OQ
uTTuJxegNnB8UG1KyBrq0WgbUzW1wNDsfTF6I4d7S9zEJp5PZFIWSz7FBEfMH1gpDSO8njBNYaUv
YkJlpXgQNFm67MGUc+qIB2Lu+UHWV89bUvz+51UOoERagbBE8UlLMB7fontFymuyzL2zFUN1Fdmi
nqTENzI8RVaZqgYjjwm3GEQnurUjgQ5+PNyzJL/EWMsIvWqVacCO9N3dNE8365L5Ea8svVyT3rFn
xKbhpuHRseI2eBmPKESA0fgzEhLESjLcR9myqhURXwDk529sJlA3cY2sqFEmkfGmoNdypEVTKS40
mhkM9X6EIxb3/Grhtl+b4J8othk+BPzYx2k/ty0yQ22PovUfLl2e+3IYdFmX3h13lZRsoCR3m3nw
ku5KUmxsVlFw9hFRWpKiv5l3IaO56whj51G9vf1CqJO8vNvuNYgUcUyK+bRfcxFwnz28ktQv4tEp
G48rpCyMzuhKHdRsVKmXdJRQeOfeZgje6Sg7VrwGv1jHo0hYziiwEhP4Hy8z/xUNpgF0mtDCea2N
sDYih+EnVh1ddPrEmvPLtE28twn547Q3TpGOzuta8GIh7c+a4oa3Kri6Kyf1jMk1fkZhEZ8bd0AR
d45pMwbDcQxMyZA2xjNWD/a3hvcOFcz6+po9s2gKWLgDxqLu97bH+DWgHEx7UUm7u1c8rbHygBq2
WZlQ43614RE1NUEbWLnpAd1ouQDu0b6gpHZTrjrKgqJSzUnPDWefIYGsTdKUPFeNLIq42HCW5xuy
a5Ax6keY47uEzPjF6vekh0P5gsjM9JIJDGQ+w+T9LAUa5YLSGL+dp8HN5TmsdXEax7iB3e1tcXJI
w6KoFkT1o8y/yJZpnOgf0dTx+87z0T5Onlj0MXmT7bd/MjyxSDXgrNh8gpTV46npHI0vzkPXVz++
AJ0NaC+GEX6h4VS3txYeDdUWvtXqKWhcWiIwDXzi/WLw5gPvDV6rjto5daqedQI4MJDAc2Rocb+B
whIfrmCfV+Atez/CQy3NDXgy0fFbg6x7Kw12Gb4t7Ursf+yj8/3Xx+Zc7SkFf+ol27ESSdJjqK9G
UXbKWBJM3m0oXJr2woEcpA2VlHVLSAzwjxB8Q1qVBNvpW0lEUkbIntxbiPyN4QLxv5uGbxi2PZqc
LThJQM+vSWsMKzePUo2HEFpKurB1lnLqBGaqNlMZR4gLzEIOwJaTYz5AQccFuG4jPrwfeIbu37S+
WxLIXtKPZQ1Owe8T3Bor2nt5+UtNXjr/seVO/Nge3Fu6WYx9NCclCN6ArKmPbkGdEF/p8WJj2hFo
SC9YXAq6K2wXCyYC+2KUllXKcHVMnewr+jOMRuAxPqHSBeTKAOul40k6YrkpUtLagA/x8ax4/Lle
qDtD8bFARdKRyKJ0ch9zTBUWEvnLr6rRXJd4CRDW7AC0L0AxeidjRR+6Oty4CkYLB5t3U2FaFZ/K
yFuHbaVHqgyGP0u4SjFbutPVYKa8cpRCcMH76rel433CwziZ5tsNVJqfIexFBb24q8uO2rGbjuP6
sE7PMIlCz+Kc45otc9LTLa/7HZLcrvMvwlk/Yl66nCaQzbNHHfYfQpzLZrPpCPXFPlVVhxSu7lye
iSdCxaBJ7vfA1eYaiywm382NCVRRqvVXrc17FO5wqNyHPTTleWq60ogYsc0yNzqJe/wYpHH5Y/Wp
D+X+ovR361a23O/9ozDO9gxHfKjP+AKwPJQTESkEZLuFqtiAykLndHqocCb0bSmPIRGE78cKdCO2
K+J2mBQAc8mj7XXXpkzpM3hV2aShaozgDsFIAl2roMLNvG8Z2FAjkf6CGCwBQqRT14uvvRDWhWp6
bMYqQF2TYviYfbGrxhmfwNc2Ish7ZyX3lnYRWA3ihcjJ4ONpPZ7ry+aAGIShADsi7z5r/4PPCzwT
OTMM8q3mNHuSgA5FqAB+LI3JlIo2q5jJYqbSYtQ9CcDwJ8MI3mGLaZFwMTfU1V+3dEWynPRN9mnw
7FwuPFPgfaiqCBZu5sIYq6F3rS4A4XpmEbX5HZ3rx/xGqjXiwhhYXpH3VFq/3gQD9G4Um9k2M22A
ZFGkjvq5fVBjl+3JERFhtfePJYf6PXQWy52ZEpDjNuY+KFezAPir4pDaGivaiCZIZ3L2joIeEWje
ZWGoah5kwWHwq9undKhLkrcCHVsIC7WdWqrC2c4Yl8FqidLo5wGVK3BCPqdWgC1XC+L0oXi96cOr
nre6+UudLX6cr+FVP1ml8HUzYTY6jythAn/lwR29FL1DWCG4WVgGsZJf7JAi0TU7v3od5ZGFUTgV
3RyOzbSCwduvnNfeOICUH90NpDW/ifX/r2XL4R/Q9VD30Tk7hrWUp0uSpiyEGZWjUYFqwbpqR8rI
9ez4b2iNPfWjii3e2ZBKYSL3SYY+/y0cBJWydsyoMzSlGhKaj/DZjtZVRJaNpbjEZchrFysMJUR/
UJPej0938uhb43+45ULAqUey6ILHZURvmdZ/qxzAvhy9wBnt+t4asfrgBcthE1/03XEmL649Dd0D
u2w1yaD5KADXd9n22z808hTZzsQjYz5H+KNXxfknFm2BvBXvAoxRK8yvVaGUxx4uHmWlwqEtwbZe
LsKWQgT6slOkFdJYZGwqc9cOBBT2SPgUjasOXDgR1Qy4xt+0as0ujsoLxUV42X63pGPalWZLiqBl
gYYBXUTuORos4fVZodL3HAJaLMuKt5KCpVsaVqGr+RPB45OmBcL3pUM3wE98X7lWas+8QZZ9uLKZ
uNgWwhBaP1cR5YebLdlBwMKe/llWK9vCgtqNKRb7akg7y1B3M6y4wQGRgarOll64X6FJYLq6FL2Z
YQmyL1xxkeBBDpg2+/tikhedWsWnLebd9pwCSXVBBVoh6QRnxp+QN5VhI/uG+WeTIRy6hb0H76qk
p+Qsm2PJAad2DLa8CUJ+74uIEd904XuoHDWkl55ffwdTLDgf7XNzROWeN0T/WOzg1WX4b6J0hPuN
B817aosCm+UCcA/F0cIfv5C6bxrWpVMpDksqJKIEK613vaNoTcbqJV3toNQDmQo/csYhcNX1JNRJ
Na9SkLC/8u7k5ESVe2pIXOMqaI7uMPky66owv/ia+IYE7JbIEsoj3XKh7x6PkViCHL0gtxJdEayA
BVVnS5mcCkkOU00UWzlgbGLWK9JSW+xST1XnWEWHIy5D59bzZkq0r/GhikH3E7EgcZKgMvqs1s0D
KtL8eQ73aZDQor1ZDwlwT/syzEIfc3BrOXpE5L+0e/da5LE5kO8NiSHKRhKdguFpdklRSap8zodC
zYNwKO+jdvSUO10rkVvE/b7psPFrHiPjbaRc6PaCEMz+EMC1QDiwWV/FOrgUL4lxNd+ZNrO+lLHj
4HtcpJH33XS6ogYg/Jhu1azmY94bhKjL8SP+Edqqjvab5y9UlP9jm/p+TwjQFq7WbN9kTdxBpdQv
oPNzAcNzEJFbiHxBEUU5kjOWu37nybl969x/bVyT6kuEAyl90vLJPmS8kX2AKFpE9eTMXMloySqn
PekRaMpD50pyO+BgwrC02+OUC49/CMsfhuAj0m5yNhwptav3KG6Yz/ctgoxTogQ5gmEaorrLL0P+
zztDdKN1XM8tZJbjv5uTsy+rn/KZffnPPVheUjzSiGdPkc3GMfKUi+dAt0ObhIB+Em4lI6T6dJWE
uAwsLlB5cgF4SD7dl/48ttcC4wef5UL2i1rFq0tQrYCCwZ9TTQkbQDIin6SoeIlrNvCO5XMtSmLw
I0dTOlVNBY51ZTjnoWWGsSCMEnbqpGpjKQo0fDaS7Uw8xG+USHLI+UgoRQOeZUWFYcwjRDafaubV
i7ghUvc/oGQ13a/wOHd36P448hrIc8ibi6Ykvy4VLrWeOi++EbPYlgwNswe8u8aWKkyJ2iOCTTMK
HIyhC9Oi2cDNoaCCUVu8JpX2N+9/WAl3jT66F1Wgb+Pqzge0i6sq62xCSnhjPLAd5MASE5R6fJES
+Ja3nsdJwzLOIwY7j57OjFZRM+w8iFbDLkdG3om1i7jPvjcPrznmyqZuiCK5qwuxuSgELXlygG+v
V7SA+dz1kDFPOfXzqoz6oHN/sazDxI1Bon2UvdiCEeOxwv7AU6FTfqPAKPasQE6OQmQP1rkKLUQb
xPH5aDLuDj8UT9W0sun6gHQWu7XuCANCJipsqKH/oAkC+SVevZt8aSI0ScpVO4sxuS7jCRDRHrAB
ae/DB32bxZ3j56+R7Pp02AWZO8n2r3kSaY7c3QAeTMw0/jFFJ+/03/unl9oVcGuTAbpv/V4FQYyn
XxvTNVUHttCmA4oa50ubLqvD4jkxss/B8XrqbUeCogN+J2Yq2Vcp5FvjvfvDQan7W6Z7Q33R6Iio
IrHZJuHrgXhvC1lEU8u3TeUUVQBBGKrwoU6pJoIub1pmZGql3Xb9HzCcrFOxZMU1nni71tE8ML6s
IF9PT0S0NtIZ4x2lundXcElcIpnC5XL1jq9LvotJng9zed24ZpaPyaoTU4H6qiO3zHL9AUQupNK9
CyXpg3n40iu4KkskqDBfpuqy2NV7rpBcxe2roodlzFpbobMGTGahW3/mvS8iHplf18xaw7al5rU5
fu2BbpR8TX4vg57buOnN5+x6fjRnLDG/bNkXeIhSm9jzibHDA1TI6yAzMES3Ykm+vVrrII+G+VGb
OckSdPjRmI3OQVIaZVYNNWXwMRPTnAj6f2qjScbHV7xHxfiechSy6Ieuno0qDIfqKhvrWQ3XeEgm
4yqvefIE/oIVOzP9EiJhKM5L+bCvoP9256T3TRKKeZqrvnHWy603UxWAG55CtVXOzMNSzyQFKBzG
nvOEfnqrZNsMRyH5KtiDvnlQNi2VfrenLoDUOhttDeVwVpXNJQ+sT8BjBaxDSv+7injh1fiQNi08
sYeQ+QtTZOYd7ZVtRH6spcTzONHQUAmWHmwu0euYtaS+sNGbDRpEgNxU7mI79yBAJrV4qYUqKXU1
nNTvSCZFh0P0JxcOiBgBLxBOUDLyf1SU/TTQ+ep9OvFwQBvz7oxbds3x7RMS46REF02jHf0i7aoW
9hLe2m2ZKENydyFt+PFdwf07Hl8A+AfCLYBysAjiUIJtHANcl4ZcDswfRN+K8LBxmXfrIe3HOQdB
WJHCYq09uPGi3LllAo+zJIdAjzmVv15SOL70INlFYUHBNWNMsWdtabftvX3HQvZ3GtbdD1OwE46c
P2iFrqWO4wTu0JoQlWRYXerQH17QH1jh4vTEafn4d/sbxFu6mhk/YpluH8ZXpYJBl+BWpTkPQWYv
Sg3KbyqDGOiM7enW25OPKNLHrTB1qsGVDWxxkng5wPdr4+NZlJT0dclfEfanTCiG2sYN8A+4TzIS
QNj7WGQ1t4nVyyR8csBrJ8mr/G20jFCXY+cXyGgdo8pM2FIl0BD9TAWXr4nRwbZWwFuWsM2WxjdA
QBiQngckyc9STjeMQsy8k+ef6/e1aykHVUXQmRT5NtXWtCKt0SFzYOOT/eL9/96rtEbSpmxuGqsc
9n3ToEZYTztark+EZBf2fQeBvLxrKxtSF03zaKdE1i8tns7gpC9pQ0Y0MmJsDgaCvpQcHvQaQNpe
jqaVl8MDLkLfaRe2d7DFQ+5Ke6qUhzW5uKLZ6kD53u2fAc81b2loxflRpqbm/NPgHZ0uCaV5Lam0
nRrtZXIrJ6UllD+gFm4ibPlToNyieILBWHmMOUDthPoJzwQfqsQlsH8AI0taikW8SgksED/kymO9
8Pe2+I8n1ABSsY/bHhPchFtuvcPHpL5j4vObU97E+Icfzv0LvXcDixeK6P8FDOATMchNi84VPIFu
eE1xR95j14Lg41yFz1CFR6CpR0UcZXxFGRMaRvujsROTxT0Bjr82lpyUzby0stWgjfRX/ppQXJI8
PVajcwdp5Ilr9EtyzBascWWuTPATDomAL5Qx7ktXJhtOwbTWjQ/tfFmiwwSoWg+FyB0mcQoeQ43s
2z1Q8qCNLtNF8RGNkSmv76IK+sYF1qcfAyQ4ZJQdNOsViBiKLA0jyuwxWlh6spPVLKoo3saI4GUT
YbnysgqVGqwTknsxyf0nf6rJD9pHk8Ozgr6DMfHa7jQXk0gnmm/G/zl/f6AYb+WQg+DCoo+Uc3Je
2PMDZDcXcdrShZclAU3/vyVYPqZVzf98g6PVxQwj0Jd4VWTBJguHiob4puk5xDEbVifRMOMXBGxQ
CgDNKESPe3s8CH3AO6l5gD6m8YT2hdtB99RPLmxEu99XcGQ6rdVtg8eltJYM1AOfXL0C3nPUOd8Z
3T7GTm5ZvZLjx97FmPzvQLY02Vywvo0a/nGU/xCz8GVnylIZFjzfDhw9QrPCvDU1etx5kC+WmQUs
+AdPz8PvTw7H4VsOaf/2uALthY7/G43thYRAS3x56yojeJKxIfPnBIxSgcxwKUHpmYZzuRz69dJn
89qkVsdUbL6QhuvQHwqTIjAsfeTtl6VB4xtugriFEkcgcZxbPMRV2/iyJvWnO0GtEwTUslooJ/LP
yhcVOECO/qCmDE3+CTsnNQPQEoKjaKZudpfrW1kUgB/mUqXCnEtL3oFjEF3Y6l91/pprvS2VSG5D
Jci18kre7CBodexF5u/qF4wC0mLyo4SN4F4k4NGhKY+z2aJX8icMKmhw+J6cXmMDyVzfoSQFfnVA
z6UP0VjXLpMuE4MNp47BdGU95HDojW45qfxRIephq3nzQUywnE8s9p0eM8N+hk5odShuJnge2xuf
bv7xfPTmY/CCp5b/iM3FhrrT5GKbxbrKIXT9xlfdH+n6Yi5U+Lcifbpj4IADT/MHWYThu4ym0wh2
SHdtRVSZcIvupuzI74JiXbpRmu8qOlEyHXKm1Zll8rrBwZEXoCgBJZTVBDuItW0RPqnWsPiltNic
fl/kr0dyFUEFrW13xOzl0Tpy5Avu4layISe6t+u7YFLyGAPDtfO9RizTir6mOjQMu4N/M/2MXoZO
DqPjeVGm17pLgrNmVh4QvIdpLElOFZbpgz0JJOLHzfNgq86mcqnlgOZxNWV1SGcVKByCDuBVZXLW
XamCo2JwFnI1DgSejm9vrZGXHwKgFJXlyG5CksqDl/968fXUf0dfdw9BsUahXhg0iZWvfTnCbtrZ
Z/AxocqNrcO9kf8SX1jdJ6EVNoE/kezd0ZMcNotUR+oMlG+ZtSieB6TYNtRfTX123rjqg4bzYT3F
8QHrPFv2RnkbYqgKsQedIO6bPEGRZOQgpgTzfH/bAGpDFyBsnhsnEF3pBaxqsJr5tcIf+J4GHhzw
O/H37Kq+kwPu/QLmSN+v9kKS2fains8zYToUCrrK7f4NTgXPdN8qGU3Yu1eonP5ZmcFE4KCPW0UA
fQnOdSh8XI8KoYOyPurs9l1cbM2Gu1xZrcTfFdNCTQuYk5JjhdCBG4FPv3fR3GaRs1Tvw10Uq0gy
E2YhdDQ1ThxLIr63n8rmEAv/g9ozBGk+cptL3MdUZ4/iTxLghtQdtqx1eS54pOQMjaq3zJPURZs+
hnchYMoj/WBcuVv1O4iCIZdhf36f7b1mQ7RKEYv1icuqe/Gri/Ve1FySTYACMM2ZZszobgpBDS3C
mUYKn3j65W8vXFhaAhawR3H3zX6myvsPMFOSXBFbhNbwE8njbjBtKHZ6rXMM1aqtECWTf0X/ZPZi
8ukvJbCx/qN/r8HeAGKDcUb2vfo3vGg2E0Mm3i3d4FsaYvtSZV064J3wPON4+BqRJjGKNDRBqatP
7YmjRIsasnEAnfyUmT7erLYykjm+S2tMn9gKAUlY2/vSqiy81aReLg2rCdCFvw3k1UozGTkpe3ya
MLNNiJjiE4/0lNe4Wo2/4QbCM8eAg/YOdpH7gJB7Ulu974JakwJ77YsHvYNtpuCSrks4V/m3Qi+n
61gtiTvS+E7jArk4wQKRuoaEsRS+xVlIM6xJ7itXgz/BAyGckIP9ShxfuKvUG/W27H32kEI2MRzR
KuKKgdYk73714x6HB4ikfUeYOndJ7tE3U98vvTcOmE7DB7OTPEc2suOp/aCczGGs4PT06G8A0aKj
0sMGSi8TlJ9j1FE5D7nQIuTDHb2BP3WWeHKgdN7qSfCNhnN5xjKLvgakmLZixU4LY3660LiwOF2/
MmgLSlN1thK1V6PwvU07gOIWQFJXvIQvtSyfU15/lmuJaU4EP22yaFQ6mj5BgKBuIwONz2jink0I
WD6r0qXJMDGycmx83p47rIYaR6o19DdTr/lNSUnkuraMZ4ZhcbtKYl+vAPf0mGCUjTux+rV+e9wf
fobQBL8MWh/Nvgb0zIuMYqBCDQg1Jq4IVZ7hy7sT/xKC4kYRefz7MvQDZgWgUmQ4AJEsr+Kd5gRb
c3ygveK2Lg5X5Guhyj8T35q3DOK+7Z9DbpxDdbTdoUr2TDOcR+p8TmhsmSPlZE3npp2Cx73Mjigx
nGPwjzi/H69GANLSeO6hQsjSOpRHWezahN0CwFN2SY7szlNm3CvtUTbkUc0FkwyXQaV1dhJXRWCd
syAMuX7nRH9ytNhKM00wDHYOe/68DFwHcjw1I27i/xU+wMXLmT5ksZb/vo5Affvh4WyF0f6VGCXY
kAjnu9qzdFFIwoxxngkF3QrJGJBLYkh3Xp3L+48R0TF6ItiamItLBlXIcb/OGDMZEuZfmrUEA3PB
4RAVLQpdXiKTjlI8TI8Z6cS2rG6UapUQbv7IRCkUrh5ML9XrymM1f1a+4PMsRLkfwHw1H9BPFCvY
yrg71OEXs/749BOFSmkoXbIZEIAbiXd5fFmkjnco1qmoYQEN8zKQviKwqbZcPq4zk8nWaeJKlDU+
rn0A4fAs32hapPkJHhqlxMO4/bgtHALEeOM8Xpta9yIX6pEdR5yC4wbob+wLN2MWwyvzjrdLjWnC
SejwBf3FUGP8MtKrkwbgR2l4OVwHXZ8VXXjYWqR1kCZ6Jo/doQK4e02wLYuamz5pjl9NZRSgnv1U
5eMbIqdqKosZ+eILA3Q0Mm++LIhucpsiLtp6HtsIGYa2Yw4yScE22KQ5liDZ69uSRrAskdqWXa4+
RNAi9wVK9uWi12uW3HU34qse6oN3UkhjMK60TiqN2TZlGpzKUeUw+43JEY5RkxFr1irj4daefepn
8eW6Kw4yfpGi545zIU5qItKuI04eE/TL9PxCx1rEbfM7fKaEQ10bvTGf/VFDbNlv9sc/pVOlmmnf
kFah1TGm2mIcNPkL9mov93WE+g99EXCZgNQC75t15SyTuag5XbUNycyrBqDonZ3jDbgTeqXNojBh
cOowhA5TlgfZxtAsid+oy7qlrYLh977p9Vbj+hkazUA7PMQIplDT0pybpG2xSA/7Nn+u0ChYpPpP
zJEWJI9TUmtJ0FAT9sY1GBhINdflmwyzielt9KN+NRemHwLDBq+9A+zmBnpWFU/h3vW/Pg7+mC9p
qTY1RJYHeIHWdzkMd9mAAWUNW6Uaivgo7X3w70qZZTFewfqrcErINRnMYYOYH9Gqy4KvNeZx4kQJ
tUfiyiAgDkj2bVniScgFZXNUK0vTJ0+o7sBZ3gLqjz4JnZb2cQ0ay2MphBe/jg0ZdSTsSH1LQLdx
AcwlkQVxTt9FmRi1FLARwpdYI2N2AI+VFVh72jA95SdO+QIKD41CB/x4SxBptJGDCM8HGfRLLytE
nKwr0MEyoqleW+Io7ObJQA2kDUGpE5RktYg7meG/bJeEBKKVbuJVPp8tp+kvlRYLW6EBU9lyQePp
Nl+Oq094CPUNb0S2a35KhbwYPgL4N8lD3i+H3dfjktkLz5iSEa+M5O5EABV2lKL5ryvlINDkgiuz
12jFTop1Ds6D52rXB2NmdxCoNJRSqcdEz1EgDubaSqLZvf6jZwXyKCzEWFciPxXbYoXb4hRBV622
FPpIbqTuPQ9TRkkQQuWbf540tLVAcXa9lNJp/m3rXWLjJHrPWUW6ykEmTByGCdpCNVz2Kt11GlCZ
Zr9KRHUyNPALJaR4IDW697V0uPuB/iX6i4ycmlwfXBjP3cNd6NKid0tiT7YDpvl6PLqAYR9CDyDD
2lc2ea4ipnqbCUsqKsOHGavaKTRDIczT+KwZtz7e1RaA34WHtgZv2N4TXj3ZkPWLaxFHOGUo0xUv
t0H/MIYM+hE9SsFcD23yh5Vp7Vo5I0NjyB0zW9jxz/mP0fTTJuGtefQn3KX0Tm7JnIhdyjuoySB7
gY9SZiru6vvzO4UJFDDXkuZYoE2NX8it2mCHrilGHqA0DNxk9iwfrGlEwGbtVA+b5ybXsySP3J9Z
n/szX3TREbKN2r+mivhcoFwKh096DtIWJ6JcrTdawlz5VJKE8aLXRnWc85oauQ4XKqOUhi3p5Va6
D9oOmS5e47HZak1tCF/mJ5/oaCQXuVJlAcY1psE81P3hc2+iEANwN3CaPCKNoPs79L6h2N/+RkZh
KuoAkcaURU68ENshvb4Ikv+p3lTf8nakgIBotGXmb7LOyJGm8qE/RE05UFivSO++znbI4lETFLVB
V7MBNyGx/kK2dQWXcRz7ahwy7kaF/PrcwN6uAbSW+O40mxkcJPp8TLpxmhDEmWFV7xUERVvN+NCZ
/0Q3F/4y5+GEqKW/zO3detkTIJGuquHX/Kpv7VlfUtW00+H74jZfwE3paijNWGAenduuc6ZJkelZ
Uv6Yh08il6kkfSyWp0AGCrJTyYBczy2tnni8FbG959NjBMEnacxK4ZikDlcoMTBsCI5lB9lYMGS5
LhNMP2eKrsRghqkUOrNbPkmQEsNRiXxoULqJXoJNpgJWQBh6D2ySLBmP425KCGmcb3ZkhjZdaAJG
HgVbQsDUOa+QqZlFTDQBpyw0cFTW1xxAh38rRuSzog5e+MJejtJQqjS4DCidI0hHgAMop8G9w3rg
XLwFnRD86tICyB6e6VLRo9lF4FbNmiMgzj3rxnfkj+kynctEsUeIzHyC7VkbHXw6SwVV/IM62lhe
9jYxQ6xMD5hi9CzgckYC3EunQZ/AI0Dm0J0u9P4cH3gvYjXmyiSA5CP5OQyEX683lvlL/zFR9Mvz
c9elBjfatfHYYJN33OkGs0UUnYGe31NcZLYpuYSTlmOtX/5Ks8NSJi4FJimlJN4m73EguvrB8JiD
iRi9QrHoJUUJcstkP/saly3+9vRsYFlkaLzb+lNm7jDl7A9wyIbA+KDBIFBV+543CGqOPQ+09AEb
SizRliT4YRhsYdW7OsV49QMLc93kYv6lIp9TK/k4r1TwO5njdT0tppfQR5ZJ+QKEl6gBfEyczHIe
dTYcY4oedVjrsLt1gjwvDcZPWWgQmd0NcyccVa2b1tZm0uNlz4ZlIGO2Fggd2pBlyiZ0tjGrXj4Y
baJZFAQuBJ+Z75OdAqvjFEPywr7V9mT/ISrWxatJfunRs3KUQe5VD8cHsG2GnbBHlk8Y8JSN83cG
6Vh/3yIfNy9l1XnsBi5jeYjcseia4O0X79N8WTSoFqYNd5dT5X0kmqRQqdHfDuIbwYICNlGAW/wX
/ZY961FJCtxpzcOXxltQzzZZqWBQgWBc2QsSfAYbJb9wzDl5k45hRYiZwFP62Z2EWIxMruItBXWU
kI8bs3Ql9vrAZN29+h1fh5jX4nCdqR5TUpwrZpRkiSUIkJN2vobfTxfWIX5nOnZX5fHwrh8BleE3
GAk18xLelf3ivT2jLUaMs2tWzrGJGemzMR8aBgInAxwuedEHvYCv7v1rtK5tCobyctUBPt5Lugxb
aAirGEDBAQWUKyWhFIwsSCFc2vZSr4vwJSptxkBYv/bBNobTz18cqcXYDnR9W2YTAtnG6ulvG89K
rjVc65M7kDyJdaM+YraOFcHZl7eaokC4wGS+tj7Sv74ecdLrngdBTmfkVYgtj9bCJxVZ3iHtpRbI
aD/INwXd4Rw7+cwy6AH2nrBxr4fEFLifRuzYme4qVadomXwqOpF73UYcqeitBbh/DQIg5MvqEzHW
n5Hx0D/snM2z/1rjTrz7Tj3lrA87U2yyCq+3Y09yxZN8FNEgsYJAcwK8AeHOtgDAIzS97VWTErdc
EedqJnx+dgGhrS9pka5MygO8nYWzlzd1rnBQP3x1+WROfVLnUUxTEGApBkOR/n7lluetqgtcU/Xq
5vE6sCw/XWiD0BpI+uQtNVPoCaP2I+kqLjq6S9vUC07qkuJDKS75UI5csYZ+IfDhsH/d1VsM4aMV
9PD3xoQppvEN/9BBjOfSVLFk4WVOR920FNmM5sRpINlMWAIAup4zT/zGlGMNoP2VDUHyMf82rYMA
mzQYNuLTDKL6zqQh/MWpFZGbYC73OCU/7GtJ6aj4T8Wvo5Zb7LQIxmxB9mLCut0iMHV4JMpMiBVa
jeU9wuSf5h/nqqzeTez1uMoKJNME0/2hVmcTcFAMPduXViah73EPEJiCMsIEaWO8u2J4A08JvVDg
7o6ozqaqdCZedrSw9ztR6aIj2ZqdN9XrM/VIVsAtd/CrD7vLECspI1B0zFF9c2fJfgl/jj98gGkc
shHaJ9PiqJ7+pdNrquFGyvropiDi9XXS2YJhhevEopDtZ7E0Mir1qM0/kSrtB2EW0G+T6/ZlTi7z
pyiK8JP0CcME358Kj+vvbvQSf7lwHpwmXABW+a2i+IDAlHtfZCVwFLNxP1iJT7bnNkesKfLnH+Cr
OJbeKcqAeHJuTTv9bxVYUxnIgmY27VSB/W4QUo/ls8szzn5DegrN4iddqbX7yX2YjnI29KCPYbqf
3cNkAVOb4JJVM0EmlXpaC7L48DK+huy5J4r9F3jhYaIyrX851zIchqKAv/P9OS0AYYYHLkW9QI+Z
jCXozLbZhOk3QumkZOaFwXlyXUL9ykJeemT8oMapTb4kFv+o6GzI8OxXkpAtCDag7xmcebvkCWNj
KRTP0lQsIcllKLpEnAj5fTdZPPluDzySC1+R15TArLNZP6n6zsC6D5AoOkbU0mljkGRhCWqbB1zR
zZQL2ExIgvW4YcFwJK1wyjuIRZwQ3bJX01+WKXuEV+0kwNYGZHZgatv3CNGSJLR0lN9hDaREcQ3E
c185HyjTIP9TKXLPRrOhWDiYXzH3/AEXGAvoovQC232dkk1xXHjOmi4O3Y3XguLhz8sLLplTphrp
K0AQsAnh80Qg0Ua3RCVzHpdcHCg40qC285sDLfhKTkskzvSuWRFNOmo/qqjbEY989Hs++Q5KRNl2
h2stWveDMkAG2UyqhW6Ta73m76oJVITZ2JsGXyhgl1RCbQGKuxOnU7LN53fT5eUa4rQjvnV7MkBH
/4qEjpgWsjrQajJODGUDZwseKz3naDQleCYRj3PggpeA2NpTe/PMGTvEhJuyNTVrp89LJrNpXIGo
SAy08S3/4hs+7wNxnWFFQdVgzyqZSq9CvvZPSxZVzfLNnauFrAGmSTycZHfgX76dSv487+KcjYNS
HGxxcnnitrzg6VtNpLr4KVSYo8hFvGPKCU2CFT0jlAhF4Q7Fp0VeR/Fs/KPTvfeJrOMzR2+rUQsn
06Ycoft0qlp8zLDdQUXjpBJYkSIHoKkzhpbSMb9d8u0W9pEY6xLATQ0K218ELrslex60TLWXvdm5
z+s+etNTeDx7mmnLN0ZJiMqKtkgtP4ZuwaWPycFLg1Il+tJC41/hbu6/3QB4xpCKrpxtN+Eq95xP
PXC3JzY/pK2T4CPYglr/FwXfSdNEcMIfgjaXa2skwFu0l03YNeTk+ZIphyEnwhXHx2kpupNDe2Vv
QlHuoHxlYkpERx4ij5VW8Y4It7OREI7N0AsMVrHtjqkFHWyOdjTW19e/Ycovq+sbFulcpxpV9/gX
cxK641iTmJ7aUTLLNAEXr9tJForcxAF5hcmIeqJLbvtKuRDWbii0RW9wut/4Id0vbzXcXaYTyThg
Z0g16EnX+CFUI7Er0o4IfR3rE56/M53roNC+gXKeLFQMQQ+z+P9ylIWEt/wJBCAqf50Jn2iJvA8L
+bDuRbvJ2yvlqsAmHxcEDDYxXeMQcuwjl33JBungZsFqCR/wB89L5z19PFI85vQPuPTkGqiKFHAN
lRsTE3SaE+ctmyQz42a+5DPhgHQ+oLSXrqnbL/OLjdvV/NJxOZWWEEy32VtuH1qFMQdZHTiLdVNO
z4uzdaPUH6A/0hpbSiLQKFTj3yWJMYCLxYQ1T14TkNUkukfoDOZzmQJ7oFFoKKVv5TB+2oX2xcg8
A0M9eAq81JmRx4TWo73QUvTSxIUq4LNzYIl7XqpamLwXc3dvHHOTiIK/y+qCbxVBW2ukzpUjhOl1
+f4wf5vpsxSZaJWv6a3HS6clFojvZfeUcMh3+mbN3pY3hlad24DTPJUI0dDn/L0rfVCLoccInza4
jVlrOe6a5g9VvINWYThp84idxOSDX8ab8UwSi61rx3GchEO/R4Rvlw5/Xhy9m8z6LlqUeKK+Bq20
uvuZXyBbs6q7H2skjE7YWZFYVvnGSbSksVrFIRmWRoKgy3drh7B3m4Gh3xAjgY08LP+2C7UJNcJS
Ul8p57oyw6EoS68K4HnLPMOKPntVhHNjIsQAdFKK5AjVm5t4vSPJsSmxPSjzH1rDsL6zjvi1Cv9J
Xb/yktaTU0QfMOKIcpDlG5Bv5YLhyGwrs4RHHbWMyEIcEDBryAWOtomoltJCQznr7YxcTzdsTfOG
1wkeULGxFSSlvm7V+/0Ps/GhQzhKNMdsX1TE/8EmHcVIkXRnAgxLPOZarBOPTbQl/UVYEy83sxiq
H1xyv2fvCwhZu9oTPwtS0EnA42o8opw49GNlT6VvA35tg6MciWleI4SUEnFpf1ZqyvhJjf9loNqW
U9F8ZprRPq5ecRBpopZc8mM9i/UMeFvnOSRdgCLCutVtLcpX31MeU0YplSUC77CWGCznegugq5yq
EAuLjIVMSam2b3kmdWLDmo3gaXKSwojts+s2KocO0WwiUoG+bedL2P5VVkb7GXJGnq76vCHHJRi/
dlbTsfWi+YkB2vYG5L+HDihzNmLD3x566/MOoLOnPcdR0i5uNneZTwYTqmZm40wlheHoJZW6OZSl
ND/jKoLsrpHrS42nbCtpDHJv/hNxvYtx88fdK46pbjvsYyntPjfc8AZ+SyP7AwjIsL8gSOUBHQZP
UEPuKBt/uuHF8oK+5eWbkhadLmO7kom/5jq99dHT+ba8BBK0FQpP9plv021zD0fFgr3p6/zAJvt/
QbylhfzA/MnFdxsuobCEkmCLfxT2nyOTJzHWFuPvz+WBAgD3SmfBEa9MJmPWqCDasr+3cdU+39PX
NjRQqR9k5Muz4W0VnQ+uM12oEmNNjNz8oyLKVXE/fidapiLEw3mrNcdAGoBb9RdUI9QHhTDWR5iM
/yUHdbmW2ByrsAVBTejplmXCR9oEetYE0dh2FoIClU2M+bg2axbTTi98Wodg76qNTUZ0xKv8H5Ql
0A+cNno4w3j5bjaAwSygH+02Z9Ks8eLx7CDBGbfDWmSCpe/zkGrUlfFRk1vQdWND21gn2htiapho
aJsvS2eepduYDkIkQrojs8jSMNeWoOt4oaz2d9WhFsbImejgV41ln/98b87bNCUx4sLuLLXwVigf
bQZtAQ5PhC51Y2xNvhIwzK6qZBauOlbuNJ4Z1H7UKCu9nbbruNLpkOG8e/4i9WHYUeHWCJMxdYB3
0G7ELT9jU9aDGAKTer8s6eriK++U12hcvXctfaTb8mRE78wsLRYoB2GVR4iHKSxcN/1zbXMEItQf
u3CY31fAHRaefr5uKvXHX8JzH31aXD2zGgijh/z2AGFSwu/iTzsPDbZkNTJIE5W6yAmzfIfThg96
0ClFBn20frQFzVWZXU85aalpfHSB2MsS2LelOFHo9WUq1Slln9Ukws/et6YMA51xNVUdfWFZSjID
r1VKZZE4PkuuIV0X/V7YHS4f1cfevCMk+NZ6hY8in1DAsr/RlFwj6q50VtstV7IwZdKmJqeem55H
b/L/JIb/esuO4+ONzd1HcvMfyWbI3ortrPP8E2z4AInUg8wrWDHQsfxfCS90Xd2desVUeWpS3bZV
qWUfGM4sEHoI3PoN6nMSiZzeSHDsPqHq7XhHLqqWxBkVelXR3YfxUNZiK8wAS2NnpLdEqQnuBnKF
QIV58zKL9WHHmTw4Qjja4gfUKlTY6HkQaHq4mj+5csGDKy8B3lP2ETdmY5ULxBVNiomnqQUEQLBl
ENGgVfYHehhRtmCBX0HOnlMFYUT1CkfOURmGDM4Imv09ZENKLjh79VuYxFXIvwGhb5OM4gKbnZMc
lBPltxSOpRCS8/VvvV3H95kjprF9l+L74bwo1praX3yM759WKYu/SvwNAWOrSBBBltwG6wLUw9dt
hy4Bj+D7bD5BCs80+7mDmpgDybtcmCNjdNdjCxtS+qhbLBWnOHpUmbwhEfF5Jihej7UuuaSt6Uy/
qbimo2RF+h5z6kVdRqpKV+yfrQWawAWlMpXVFleVZ9srHPGYJ6b4d0xkufj/r7LyI6t4hsnDD5Nk
3v+Mp74LCv1amLdxeIuZ7mvP+iSpOQqyv/GFcBP/E0cQekT11z7rqtQctnOWvaZ7iKGhhfzIhvfn
cqxl857T9qic6vlxM4Bhgm4Bl6BYBRWkDZOxBwIqlLB6maJwLhJVUxXZ4nA+ONUbmKqb7mXryQ38
PHdMBdXmYKkcWE30KeD2VzvbGHvPwLJ8GWP/fkCiDZcHyL4+uLVTcG5hKH4eLneRsGRoIEyAfEBv
RyXW5pgCtfHiJhtIvnngkxygKGEDil3k7+YFNbzy4cSJit01pmIA01TbyF/6gX0/Q3Hw7sb1Sm/R
i+zOqtESvbHxCYyLCAbzSQKJoTikM1k/nrWF2U8YPsigf4+C6p/du05MtSnZEtWJPlC6BX9NgGsp
U9fYuqQnmLcwMyhmdOEOZ4qCvH7+s342MbyxhRlKGXvfBDcshQivdVe52G9leewn66Y/DnDi98t8
9jXCSzYbfxR8JC9KXgBDgT5r1wLNiLcwy+zbsNv0nSB2kSbkgQ2PGTRQTyZOByH8IbXEVLyNOqf9
kBDM1zVX8BT66OhF3JOScdZ5D02DpcoJH68L00yjoiUihy93rVG/Q4L2/6/cjX27KunPZRRTTl3t
GO1fu5VhP5AAZaC1OBs2Y/A0RvuiVi6YgXkJQqaUrAv9wkIe7SBGlio5VXw8GnzQYctf5xNRgKwA
QDjI27mZ2IsrajLVe2au0odRJnsBUirJEznuNQLzmcZQ67aSW17e7B5I9jgtAMX+LuocdyxFLCR4
7/Dy9xIfx/9MJ1zjxW1wW0Dx+j/+4pD1AI08HgRpKBWdUI+fY2wPSRHwLgNYBZ5yHvFGDkJ/HChk
QCKJaHl+vat8YCiOgQnyecFv5ClT8RcIa9n5G/BOd4z74SDBdCvk/UPB4PT6V86k5++XhZBwK18Y
HBz1sjJgLhk6m9qVueNlTJIxte0AB3dUF2usqct8A4+GOunhMthbXA06mH2rpD6Oarv4BV5U1/gA
EBVzGwA5YmGntw+c988BDqwJoSZRG+HUU+wJxanNR/NRrU/xXl7OT7ccNIgO3UnEoBaHg8ihZT+L
J0eCsshCSkzga4mjboQu3uIKSsgQo4Fb3aPfKnWd+5jd7zgrkY+5j5KYsqSZmbjTkxEndwW5nOnU
O+mRXUYI6NGuPr7vtQr1d6C+b9jCKHVbXto2Hi8A0xILheAgwJfNmUDn82/vMuFADmO8lTQNIXEM
r5Q6JzRKUWwgiFgwzDQO6Zo4IfVIpajaldCcHN+oJvgNoZ5eVUUf2yLHURWpNhqKPnb55OBDkKVt
JPeBEyUPAA2196NCZGaDuyAM6q2yPYpg6M74PU66viScb9uqBksN/g3r0G8eyXEHkLfY9qT3ga+H
ck4ugpl7rbQ4Q6g5yuu9UHxkKZ5dtKmhg2F2qqHuGUhRCUjszpfXvNyFMO4GJw6lD1PJLEV7Zqoh
WR02UCr26zE2gsO4sME8IWHjMtf4CawEsUFqt8F+slawTQhyPZqdCs3bzw98UsbzA+osIZfNbrUt
RNJ0TzuMKbs8QS4B0/8erPxUKVRCUs9AFHJf6zVp1mtYmtjT1wk2200qg/FpBVrSUip8BN+c9qSE
G+loalENc3yNdjXrcCS/RfTyAC3c2CkFabkxGm7vkIs88OPf04A4pXeBiSkzbDgn6W/oxEQn9t0o
MLhTsTPJYYBhjNlsrGDiTxQnpQn2LFK6sAD9iVlX47DHcOb+KYEAygLtj+AOB+zqaP2i3Cdv//gS
+gt1FfymN7zyBeULsqubmI8dvssBHU9uMGvt9rBduEDwdsbZ4CWFXsgJF4HuTL/Ws5BR8QQk4JU2
p8vgFlPwkVDK+SCQcuP3dj9bxx6GHhJ2jShwV13IlIvbe2qPkba/trLbuqfce7dYKiGb3vpCglTX
XXOgCaLNGFkr0zsuB6W80jOYtHoXvINIkLIe7IpGAj37hlrv76sTAHmBZFEI55j+UkfdQxu7jrEY
3r0kLdS10iq4005obYe0Ud+gsNgpHAORXX+ybXTsrEvBNtYZ58VaezJdwhMxW8LV1b+RNbu0zau8
1LDhpVOphcaigWSRm6RLZJcfhBk1Vm8R/ImKvDLFYB0SaJ926j5j31CFvrlWjhes9a+MJKZJ5h2s
XsrdUhAwjQzrHYTfjq2CZ72nUM/PgXL5qyRArcmq3L0407TPH7LCEDRS1N1c464X7Bx68MFuz5Ut
uRySarVI7jGuROYCvG1rS/S5GrbK0MZwKtD7hBZb2nL/4mEduYkbVVyySPaFSabHlvRMwz75e9Tq
lIH9d/mB7nQOZh4YZGphZArQSMq6VbqBcly6fA2qbRdj+YJD1bFqdZ+Y9Q4Dgr+l3OtxGPXC/A8c
WoanYFgXoxuFbuKiTd+FYLSQ7PryFRA/YM4YNf05LeO6vhMFbdYykU6I4EdTcALmIKGeT8TZvJ4f
bj9Ka0DU7Iy+kzgyferyeCmZC8t9CZiLgXYsdk4yP7i4KxQVI5O7YiqlginDTtFHDEwKvwCTqjdk
WhQTaFhxfXem/TuNJmF2m6rRFf/8OmXHhFR+rqH29y2AcAhIRMCI1jFjwNF8KNfeGIHpgBnJvpFJ
67+Sa4p8PXnkS7fWza3kWS2k61x6orCABkxwzIYFbITcDQ76r2nmYnTV1TuX9YQrgOjOXw3G9RCx
MfJpZZjbC3amN/Jf3IW1DkBgEjBYs3eiJWaF/Ua1SBVYQLX6rdDa/JYpTYRDcIYPAITuCAunPAd4
bE6YmsBfLz2YffmgzzxW7XbloqvBveL4lB4S40AD8bhYwBKY+CDOniMvblFYzzZWfYn+d9h6Gp7I
iobKm7cqwVnJfy3CHqeqK1CrH+3er6JS59zWkj/we3lmQlr44L7oDv+rzvDuowENgonmdxmAVThC
6rFUlf5PqQynkVojlYh3Eu+iNQ3lFHQHQCQhWze4tH3Zx2J13icCD4H6gp7qk0NZYywtxV/wIBG1
v+NzLRZ/Qi0onghx/xjMReREwZzcObTOzABaboJRGHasmBU1Eh9qZL/ezp3kJq1HZE3yBd0OWEen
rYpVlBqxbMWxg8Xg88Ch3b5CersqyIXWnbbLUymr/c3I86nvM08NYxIkqmrGWV12rxh4NxcIbAcp
8yJGU6fNaxjNGlsVW58h16W3BhC4Gnoq+P7VwrsnMKwuAiA18S6ORRQZl5WEGmXsnQ20OAhXEPON
ZzF1ICJ+pJEnQSoYosIPzo7W23eZNLzj8LyHzzXHMqNGx8QtBPC12+dPtiRapiHin/SfXKocr9Se
2NRZ55JhYmVoowJPmLhNA/qf2V/uXxXY56nHpI0gSXVT5Tt9vgSeQJMJLEqbkUFtPQbgE9W9Z+k7
qFKGF83+mlB6aJb88JNbIV2M/Gxg7w/4k98sWq6r3XnoDGn5uGaRGJboFPsAO4Gh2Nj+c9L/+Q9S
YTj2aBCSTL73sWhporQS74uH3x+YeN4Dvcrs2Zj5SgNvkvshdySPVyUxTlHtqEwkkHvRiQn0e/gK
tS/YEFTur32PKQtBCT1JymsLynm9GKcK8VrkIA8OTaf/OwSf91QDXU10Uvq7EFeA1FsKZkEXRsaC
ND7GCJ6ecjlYwxjXWXAP059ewYPwogSVXIB2seSJuQMl1y3W8banjf28X1NU5j3hZSY9jh1+96cK
2pN326GKDR16bqUmnj9trS+36jqR1UaHpZPg7V2to0kXvrN1pfmRv63H2IrHY4r44yojJPp39uFa
XXV8Q8JOlkXPMuDAolyx7TMPxCjWdox0i9Noj84ByDkdCsYF9Jt9TIYyaln1pUIkQvWUDZ0FcBMj
iYdDHjpS15rEUYkcGY3x0kIadJNnno0LB2zHgSNqGCmL6SkVVIkLiUjUio7YZTW10m4iZAbFz0lm
n3KCMg/C2Iv8y1UGykAi4dg+Q1HAeMhyDkxfmeSxD0GiriPulu5Xs44aaAoByFgkIR9pkV+gnKS3
47AMrMbrIBmpQxqM55kdkEWFf4N8WBk+t1WjtbTfPqv/cQKpMLJ7w6HAdjun0hdpNfrqinrRaUaQ
yu3QghO8phiw8IrB0YIE37RyICEpZROqMbwSipKEszLeeZlSPIUFOWhStpKAn5vgJQwoM/ok4mC/
aHl6UbwLSxkItvWaUe2A+jcqds0IMRAlTujBMshVcSM19ga9kSHpf0GYnX7Z9B30skzjWfzaIT+5
COqV2iyBHp8fsG/hvd5/mVcBIes8fezHskH2nBjVl/4ChRpMNNGmhnY21/r+yzSeAgYkyQt6RIeW
cm2MVhaeP0UvTUYvdTha/4fLt7Q6OeiQOMii8blnbbp5b70YOfV9jsSlbWS3vvEdvwz64C9EQuXd
RLPSUPX8YM6B7znV7s/KFD2dwPFPrWDzyeVAZvg100TsEUvy4NC9Cwvof5epjimZP9qkHWqV7/nB
y2AnXqoqIPrZvTdNqpr9U4IsnFYb/oIhxbdKzV/lnxHdTvJWVqip607cdi0PbFjZOR+JwKxGWfQs
4kvX6gVNbQ9RedXCluFzTqn2+QNG6lIv3rwCoYfbxJ229P1gtvuVUJTasK5XwAuQlxUG/Z2SA964
1OBaotm2mqCIIyzT6qbtHA+ZKX2lxL10LOh52FjXitnlQj+veKtpJbDZGtCbYXq6rPv7wClUOHjb
4DkEPrkN/loJLZXKM7RbkEcdnfpbvAPryhijdAdfCYyS1q4PpNReLoCBPccxEexwxtdTRx3r0kGv
JXXvZP46K+IA/w4tAdXKlBJ0Ecz229/H3HPUAqHB4rGwHB986LW8j8GBOxbXJRuUEVmzMa15R+jX
cGL6PX16UOzBpZ8UqXRGxAWe0wbz6ce08PGDJMz89SlouoNA2x4nX0YVp+v/42v2UGaXiOgsCTvZ
1s9vu11em4IfhlC94zqVdc9/Ex501mGVFjMJVPWnda9BPlFtTH71sEKVe1be66pIHrmiHah0txYq
YhqXmknencNLNtQEIoRgYcQRMro+GA8N9zoiTBGB9Ttxhb4oVEZJ0CQ3PFIq56eqqv4ryXm41x9b
tai5RCBHgbhxpfWUpn8rUBktpUdUVRsRRlxbRIWqI/QAzjajHd9gJ+ymz6Pafz3Hs9LDd1gsutfm
Jw7eztqoIYIBWxJj0zW6B5j31sPMHg5owVbJ+gtCGi5Pl5u76wYiCZ7TRZJ/zmN2pF8HwMdZSZZV
rgNtTTedidOgT7unsaCopN+n3HC+pFcQgIXutql0Ks0QyIE62S6d1cm4XWQ7IALljHLobjBO8xeo
vM/kowsCUOLScoZMWAYsBJpBWani1fvqXCxjcqym65mESnbsGSbJdr0WGTrNHR9TjWyrc0I1/Y2y
3P+NGJC7BHUBbwzMnxCVbZCrfd7Fmijawd1JCqrl4SVkppZHcIJo8PnIJOLXh3ytwP8djDEOdH3P
tqQ0AJLXpec/s6FqK5uuwHQ6pZnGnf3o+YJ09hSWQ6pscpbdJjgoL1/h7WvKBdwP3WEH34/kw1BS
+kZYKtxsV7IlY2bv4ABYCHHipBS8EZRqUDBhg9Vxmclp+vZattv0EPhD+kUB6hNVLZ/cUIkkQRU1
K91TqC3ZBKSLdDSK+CNTLcR9aFw4RlxnNLOcXZv+sxQr9VwAgyvQt40ryHPMGstUgq/sYqeFfEpS
AE0Q3db0q27DY7zpTkfnHH0ueT1oz/uFahoq6kKx2lnfcSfAkS70C7HbXaEG6LFZaNINd9BDScAP
4eSDwHooyhjPve8xl4ouqR6+ww7C02V9RFjq60Gr/X1G1Dv1jMW3C13AVUCqCXglGTEQt39wIxOG
WhELlUhbQNoko2KvtXyOtB2pQ5seKQBmlY8Sd+WtYcpv24jNCAjUKnB0pdsGqd5228K5oVxljKO5
FmlhgV9mMmnTTlgQCu4i9dueuZaWz5N1XbNQyRlzp4thoedLsfgnsyDywhfm5mdG/Dg+/1+uuPGd
GHuE+N92xPiuxWSxzWacB8NT/Twwkw44DkuQml8IoKpr5DhjrIUhzVMZVSUhtnoT/g+rQGTMugPC
qdB7TIJr13o9owDF450aJDoO5O44RQ1DIYPeHVcXbjlptimRrYjHDv/T4YeDAA8eX/s8pWhbVzRe
DZV/EmgvY9yoE5+/kxU7CZfTZ16y+vwcFgwy0mZ6wTovbwIIIhN0I+YnwYWuwd85Pk/Rj6V8S1qS
MgZIJH7ZJS0UYJNlu52EHqsuealGLEAukNEHFWajhlQ7AUKBl2BO5sH33sSD/Z8awH8710RDjyt0
om85gauAqq+8S1Y5gyNPhQeqmDNSFrmGFpft7kVa93scy30QvxjCV4tEyiUPQdObpAf/wu6ZsVmI
e3qHppKmteOCUbcIXb2IpbAL9OEPiZeRvCg6pwC1MJkmh79gwMho09BSDV9zO2vaSKEmQWcrdtQS
99b1kM6AKYspUqqSmVQDY2h+hfes8o7vLFJConSN0z7t3Fp7rszuxNOZAXTTGwzbDOPTmmSgvsWW
y5tEVApoDSSKtezChqUOnid+mhuzHnO0ZNcJpx7ws186imz+Xp4no1j4VgTXng/9AWW9bxv8tSFz
fHeGVOskYEncBQpWBKjGerUk8VYxmJlwb+PSXa6aXjfgCBQ+iWKpefJN2zo5xalzpGWQptkEYNDK
cpAyaMh6/r4UGigH7yCiApZCh37PwW67RN9+br4XMNFTzkHN0p6W4n5jBTkTCsRtzyJPBGD5JogY
8k2XAF/yhlqWrhz9DSBrQ1S4q74FT59vkwrOrD96xJzYNLi2Em1UFkFAeY04I+ZW39mUS30iC4qh
Asy//++jQt48+zmhZHstYQ8i4Q7UaYJFJl+HnlYYeb2/mkw0u1DH4VNNavsesm16Qfl5ISlurdev
gJbTcDA5pmmuEhw6WtUDnIsSrTbjp9RbeMYOdrFnuOa5JNhUTXjXUeKWLgRrY8nKzZDWgP4YawBF
S8Jal7zO9M+zgrwHe5WLGGe9uTwSlJ2NG+32rd0DL/gZALRvJvBlQetCiLTy/SYTDSqE3Y3GWYkr
pVFgsE1ejyYRCFi1tDOuRtlFsF1vutPC0WZn/5OuXmhCMGc+gGKhe4wj1tYEJ+wgFJbLqXNhVXGg
KYPjySPTVSGrrNFStQtoCWOJzdiLzh5dk5XTxchPZRwNkD5AWyTwRTAG01bmLi2tei6bxwBmyHWz
M7dMPAeCX018SSIIrn4oDzrHE4pMYVqPebWZafYfLiQxRqH1G6q52JBVTATWSyMbODHhO0/Qfg+2
xGfv8+XBhufdFAWF5/a6REEguKfslaOZ4KEx8fvk5L1LZzAFSBr2wNUPrUSH2eYFJwEZ24BMY1tU
8TjcR9bC957lzvkB173tI09lAfwSlc5iEfG61WU6PQ5LQAPmSGs4McXqnJ5p7EYZSD6r+v964k7H
AZlCydPGmtiQBd5f8kI5zzgC6hYoiGuVlt3yCVzPLM4dCNzYtxEZw/C7ilBpjYqMPJzb8a9z+5PQ
OphbLKTMWKxvJzy4tKcL1cuxvBKtHRh51RD2gkMBJLkbVW3nJ11kZ5flpaakw1BWlStkACBkwUnM
bJCfBPUPmxWIt7Fw8kb9AzbO37byEPQZP03gsJAktFVc8qUjDQ+SsUIHuQCSK9fJXyjt4XgH2Hyu
WEBFLKnW0ZV0ct+vplzV+SIr5FdtqeMcLs63t2R5EM5s5CR6gioifVtW08E8PgsxzUTQkj1SPGce
mQENd3vdxd68pcM748L1QYwsNltU3g+wnO0zgERdsA7p0mCcXkEGU4MY77sXqAUMe7FVtK13nVmA
vw9gbKVUMOSPl2jgu/XJLBOBP013l8D+z7B1lkOkOFkS+JwoFmZMHKuP7647gXwltohQDo68BYC/
YPTW5+4Sktcf5/sBqoomSfHA4ertBmnNr6LmdXJsYciqJEGAMXhLqPzpbRoeiF+AuL4RxDkG1Wlz
kx6ghnLTDjRbpBE/K3t6jUY95U1EKOIyRWwPil/vAS6DPmPZogT5ro1AAeuJmuyoqII91MzOP5eq
1Qu8y5YyBmGqfQEFWh8Px9IugETJ4upz/ljkGoIgcRx+sSsejAhOIv/XN4jQlai+CDoPEi8/NJj3
cfB+ZfO/ycknCfUvBww6icC883xzVNYSzY33B78h+3MZdmsnagnf7jbX1DYz6lAlJTApfAT2M9xL
I1CHpFR1wJZMHLNkWsgmkWv0M1VVCLNaeW9oAVefZOCRxLUqmtJ6c38TinJjm2ZcJQmfPDgBd7P9
h1Q+8Ic6vK+Jo2nMrJ/0fpLEzr4l7DSV03sGKC5+CQ8FqNzwxbiFqqPzfkC1ksY5iVoYTLriPNmi
aa4XEalgy5ijJWiRNJmDO/AJ6bJ5FYQ01KSCbW0L4uKyZZ3/N6SOJ6P76OkWZBPaPLAggK9yg0vv
GTk0CSxUeZExyxx+a3bax+5RUyfwMzvd+XGGAZBLutJCpeAhIVWbTbCOx9X3MoAWyS786Mx4SKWF
6yFTMicSvxrMf7y8gS4VZhGIDRwwmAmUMr65AnXoWYy3rCce3FjgCJwLxC5As7qoHdq9LhGTaPE0
qcXN8iJkqBwMIkiQOskEOCzfr27/1C+yRlUM1hKyC991OMe0nVZtQ5lEidNM3sL2pw/D8h95Nkdw
NCCuRi6Tzi5WrQWaB7FTZDHfkFU41hXgVWbVMxPs1+8meM+EIv2vih7cHq7ikBOXKEr0wew1Wa/X
IhdLzV+jcmLCsgNxW96i3+dn5Sf9x32GvYbohOxZs8qFJ0OSzHaYYY+/4ZcbIKDVGB+v+kkwefOm
oWwisoBr5UflhZugDGKNL2vTGP/gYdzvunLRL9i4MSQHzP7yWrsMVreOMnj+3Fl6QVGVgJEfi1Aq
hNzyQ2I4LFbhH7tSieG8a1DlsyooGOnUyajAq2iEhbeTfn1pxBtHXxRfzTfWs8e7KLAJ7dT3MHuw
B0+nhzXnwqgH0deXAthIPqcSPaY7IgPRUuyUcd6rTyZtb4bvjYl6NC8BLZEnESxwhObHYDoJinxk
1D3uS1Y4WLimE+VqW9owIYGG5SyTNggLyUBbxN8LrtQdSxjNDapxJe7afOF0f2ygHDjhRwhuYVrG
jQcB7JsuLU0Zy9/B3QkZ/Npa859wxNIGgO4gCS3HfwgQezrjHcdwLosUrh5p43q52HUa7dQuVFvn
lksIY5avLlWjIWq+HSLlmnTKMNcqtoKeAe/gKrtKMUEyjzMARxB4oLyL+8hZbsBurThYNJqjVQh4
XsGuP+4ZiTZ8BTngJyKpQAuHHtc6sGEx20mePLNABIq8qDY2UE3FSZw7BINuV/sz4s4hQ4kfV8la
yOLikUabIsw+CevuvgREmxXu1/du7Fgs0e7p+StSsVuLk4IM4QnDDBa9IlqVFyoQmJOqB+04rdc2
fqFiy0Z5E1WIWP7yI6lNJY2hDZvfoqqGBv6HDHjWVYKUY8QGTulah4iA4n/sDuRafdD58CPwli8A
L8UFP9EBfOiYa2377TXzSWy48Ngr1hjAu2sI0gUpHKYwy+UW7oILvfV6P24Y6ST11zTt8oYXDujo
xeiAiWnxfiMytPHhDfVygOlfE0atTBN1CCIXsUdGo2G0oYC2K0fc89eGpS/pEKSRqj5HA399UNoe
ZpC45Q5NNEDBLYs8p9BSHpYKOGEuQZ1N7jodlHvRXfxqTa/R3btXXCO0K9b9PVxt12qumcooJe75
OH4mYT5W68ALXmcq2u8u+sSXhjf7D97WnpLZdeXTcsrWdmpNawvlVGKb/JRes8FjW46weGGTfwif
Georeqo6D752QVXdiA4mJ3CojC5Hq9/MQzM60c5veAhw/SrB1lFI1MI2Wv6sN9Ik6A2vVkAkzTvm
CoMd9taGRzAbzcSl/NQDG/UyrsupUiJSfvC9WAbeO1UETZ+yq1r7FBiSpr2Rhk/bqkBT4XozA5D6
gzkiO/4GD7Pv0DC9ObDIrQfXQs6z0Rhz8VNfdQhVBmC9jSet04q/abY4bvxPVmY/B4SEwzOMcE0r
IqVwBtPcooEhyHmWHm5yFkN3oraMJsaZ9rENjJPETRFPyAIXQUdDNNW8A1tGGVuc5Cy8Zl618wGU
eGvpiqZH9I4suqx0VfdwVzbBA71MD9JAM0oncSJCk/w1SthC7ZCn3NICLIqaedhAj/hkyAtZX4CF
AIeBN9Nc2u7RPNMQM0vgE88D8nl4sUcear43lr2c368GAUw2DHj1XRXLAxW/KpyDA8Fw706eUByK
AUpMqARWQbhaQtdzcQ+VPBJNVy3/Cc4BAaPS7AjftT42goKgxKFckWq1QenRg9IUwBnqRjbouChS
4YsNiV6yCWJeBMaqVAuMlT4vOc+7ie8MYQzOyNtpCORlA4ZBbsjYoQORZUeWNgkhfoD2pPyDjRE8
E21oJyCplyaN2srqx63WCe6f6h+fMl6Yr7BHQwjqnmR8p8dWFzHfYqmybM0sX3H5EZlb9ZCPrnlH
euxZFZ97az4Vhozxn/YHKszOgN8y3/Uawlv0t30AW9KmSjX1hCR65oUMi1gndWKA7Cqv2sDFZHqa
YVmzSXIAlZXw1Hf1YLKKQkzUBsDpfQHv7CFj8W/dydpPvyjiKR3KzahRbzneqHZrTeZtwcQbdtFI
jzu4ACAe1cNSnH4TOLmmR42fCb67hVLNiP6dbQ0vHAiYIjQwuNbVPgcvotdms6JQUWXTjvGQTIYF
jVINNNP3LRfuCR8+wNMjy/Vc9RqPvxPxWoQiRZoeBRsvo3CYOfBBHbVuHDA152v0H9YxAA/SDzR7
OwJ3LrkWR149ANLQHqA36Dwa9V11MHAyEfRBMdeJezCGZMTWqkxh+RUz4B9NveVLcgNAj32kGdvL
aQymkb64GnPcoO+aR/kIgKaqj56YgCGiV8vEwgy9YeOhvI5/iS97J4MpYKuRJFjFT80Qs/lSsLdR
R8Yked86clv603mkj6rq22gFyqs1hDClmYgklWrKLRfj6fCHf3s2GU8XF+o1jIIersjg/VH79LVz
kQJJidxjEhcwFzl2elmJ3DolDOiYBkJ+zM3x6w/xO+2HwRQxmIHH2+W14JU/XzUV5W/g/vu47I9U
iZ80MSIBmgqrOGVjFM4cCmxH3388iwaDLYQH2XYT+W80uLZ/Mr+bdSgr871yOvHKHsVK/bW8GDvp
aRvfx5n5MUSXu11ZxlGRRT0nSLlBwXjCjrjTJNJHkUO2BDqtrcNS8eFV4Ubj4kwr7s/n4gHhHBt+
mcw9J8f1ank8+7M1Jz0jCPdWmcN4r6ATbSYM9rXWyOOt4OPgxQ0hZI2DsjEg00+j+Sax+piNTJyH
7kfpS68RZUw+UV4cJgbBuLn775C7rJuwwebwsXUYUfBoe8mZ9M86ibWKPJr+rsopgD0LIZGoRW1g
k7ncuQ6eAaviLxhNNBpzI/aey24QBUCa/F2fsMTep8dpaImcFu+9nuy2b67fCOU00OVJpBmSFPPr
0/iz11dDirM9atZS8OHizPLVB+p3/6J8l+hei++EGlobnay74akGVuCrUQa0zcW2nDqjdA8XLpzA
8P7Jj4coRrYymvRX0YDuLvahDLIAMd9WzxRZHTDjAglCKf4wZiTY8xTlnFgd1rH0opGmUyBEKMnZ
M6i9KAR3MmaO4SkYcErmDtNHYLwJlh2y5CynJQiLKSFquj1la5rvTE2Ggp5ryuCTbYR0TpH2LggF
tjM87nllFqEUrRje2pN1U4isc9RWeGspO6Ztm3idHZAxB7WEC+fptwm7agOz93iLUPpX0BpUXwaS
/UbXHug8vKckWKvoaMiOsJkaf2M0Xd/bXKGe9yUgDXJiIxFMnKrKaHx2MY6k7DshowlcDuvfYbQR
aQHIYYL1rWp8/aYq1Mukl0itxCYIbmiYvngYGYYZ1MxPg6a1K6VFlY06BBCuUDwS2O1op0grnmYL
PBwcE6RETIPsULe6JAlw75N6sWrYf7LOnTeNasuhFFi/Gogknde9gezrTjke0FhsX+QJpf2R7NTd
eqEAur3xPM1ZgXwptKZ8wi3E4VlMfWoa4/cERiozz92KRSRS8gDRS99EHH2mhKOqjCoMAPn2nlEQ
Fruu3e4WIQXfNT41n9wP7IGVLym5y4RErJ6i9cKM+tOHSIf1Hqy7SwR10xROUmG7P9sLk1Fz+9dp
IARmlHWWVaL0OMdz6fJwyXL3cIEgSIBfyUZIkzH/JkU1yLjGt3+Hpjay1gCNss5fLB0CU4B6yNgk
7jlKs+QEi5B0Bg7mjlCAYUHa1O/DKdmEOJmEsfXf3751KnS+cIFSpVNPSa9BDZGMleqxYoChc77q
4J4kAsBcGWFJ27FCnQ0BXDWqxILzvdBOQ3NZJk/U9mth/7XpmNuW0TTumUy77OKTjeQgBCiwHrqC
wOAv0pnzoN5iO6Qcn+N4KKJhlcYDgFJGHElsnX2buU4GP2I616ksJdc/42ahtg4hkimULxPTEavh
2SRiSP0Umn2GJcmRWnzRwONoNRXQ/BMimFlAoQg8wKywOM4z5/t1wBf+Zl5l/QlTe6zB1wXE8E7U
ckNRP9HcLsfN6DleLilgNr8w/SNFCCgNOyWLV/RMJvTLv49IeHuhKbIw9nyKZOlwkFI+Uebl3pry
iMLnX3Sm8k0Gq7DUO6QxIusZUFvSNdDC4+NoqzOdZm2ZQsDIrfNSjqRlgiUoeuBIRpnyE5Gd+Lwa
gIVTQEJCXpitXdI0ttYIQJdIak8A8g92lGmHrznAPGGk17z3caFs1NAmaxk7wwswtkHm92fF2pKo
HmEpFfBaMPXCLPRQC7DiI2i1QJw00i+8y1Z0ouXloZanHe+JNDIVBxxuB1CD1EVS+fG+5mTq4+nS
mORWdRrpi+ZISGlDw/rTRcSKa22hNuIIYDrEEYBZwpoNJ2MWtzInYvi4/mhqoZHi9w92ZLOLkqws
WjpJWUfpT6HU0IaBEsYH1PUwyDCl7M5hEiS90pI69neJ4HU714SO4d3buCPdfqYMMXwzFDLGqzL5
3H7DI6btjOpurvHMIzeIsvJc63I5/G/z7n55t7nvLCELki4/gO6NbrHXfssdYs1l/8Q7CxuazX/b
u/NamIh5kdMuiCaqqC9B3ix91eV+E94Zgbko7Sxes4FpJuru6D2oJ4GsixTh6JQgyZ0mNbtyzvn8
zjEu0WLMDMAMkW1PBDP6AV3X2Dd6K8NNHmyYKQFxNzFdItTUDL4vOb1Oskw4aroOauogA9RbOL1R
ea5jL0uGPWfnSxB4113HXzRkfrwgjflqFIwWYb9WEkKFr+az/IR2/QolHNhOis7GsAzqptCCMLFy
fzPkSn3LeCm4Ri3IWno9SCXmlHB6MFvDnMZSuwn/nX5eHR/xvsUEp+d3EE7DX+pAD1oMfQGHn9c7
OHJxYRWNQxfnQrRfKOokFS8phdgt5zK1jBt+qoOuaqCeOyKdLkZnmcqV1ZO1PA4t0N7uKvffREl1
hunGXaFV9OyxrDhadu1CakasBWK4/7PzDc2GSA6gdR5Eu44vVo8l4pMd3yk0cJ5Taa1fLI51KSJp
uRvYicn/NLslU6PkiWdUaKAAuVr+O0VKEQOJp2ylpnoiMw1F8AkSDoen0gnfKWSGxKXsT9kMHiFH
5yBakPAFy7ay/BhWfAJOftkqQYPykMasz42ZwVyOf8UDm9gb3ioK5S3UtMuVH0WYTK6WDwgeQ8kd
UDQ8srbWKD8jsYngG89+J2IrarwRVkYioISYwQ9AtxjNqtGIW2kpg85DwCs5T0bt16HZOvJQqTK5
OLHg5bWuENJQXUg7fL3m5rTzZfpWPBH+Riix/Czzb06RFvYFCx2E3mmhmmMer82MPzzajUkMrzB9
5lFu6CmTqtDQzj6InBKOW935atjIsNNvdPXm5B+IcUk6mRKDd+L7fqdEzjmA0DhNJ5X5KGYAKmnK
PE3ByV84nss/D/zKyG9g6GdQGtfm9h2WewAQ3g9LcX4wtPSp9pIRLSYDnD9nrY96UWV3v40TeUXC
k7iOZUKvhKc7aj6oXGJIzOEfG/syDo0MmQd55oZxNtbAQfD1LzkRnDWLUyu67LgF4R3X62VOisLx
dFUfLb4meZhPkDYCiRFG+oqjZoBpqIcMmXQRFpXP8NH7IEAacGS97sBUd7y1bFEtIFHkz4Wpc8aZ
I2T0SUIDzNM2psxMH4YjOQOSBP2+8FB1xmGPeChna3UFTo5qA+RyJxwIujtMFRo3w0imJduX8jig
xXPbSZBaBU5qMKGE9klHmmOcQHSXLwQ27rWdfVx+IhkA+rW7dt9SwC2nVZMKUKZvb3UD07p6eX8B
slvGk30htaz1sPGd7SD84P2OxzNeaiClupoSVcdKYgdK/zNojZjfZjrD/eG6QPYQsGOfkUV0Ej8q
bO4LR8q6DP+CS5vZwxHK9GglR2y3JZKidfiuQP0bHIrPZgpUMetxqyhiN3RVY8VD8QEuXOh0TM4o
WMDKrU7sb/Oivzc6lO5baYiivMDoH1eyEINKXaSl4OLFINiGTnBRsM8FKsQa3Ow/NsqhCuh0z/GD
RCMfzqEBaeysuhgPMatMS/5rnscqz03xJ1U74NRiTehtE4MQAAX2sGfsHdHuX/nDsd4R583HEmXM
OqCPgbskVPOTlcg/7zX5WOYbxKvRdTrQoUYMxPGuzZelE7vpJIl6+LX6Mjsn0w+nJIMJvQiwP+6Y
zWx7UjQ6aFR+Npo3GtwNwKCmiNKlir/1wCpeOmXQiIYvB72QLUfuKrlo6WtxqXwkHOwI98Fw8stS
YLeyPl3wzbN2Q/lycvUe2RpQOvW6A7aRlZIr9CLHLY+Q5yU7XGRcgZU3iFW0Z3D+Mi9tlRGAi2hj
hovV4NZXLWkzjYq+GCvMoKunQZq5hx8yQGjInsQ2Dx2lYreY1MDz+gydjXCdg8bXAIPkDE/yvdIh
sw1LzIg2kvq3gH80SQCQvM/Ybhbg/oLCDSrcc0ht7uhio5aldyrJLTUI/2thSWm7bYsK9Cfi6N9b
vV7DtGGSGNUjRCBzvuNooWT/t6/osnHVdm1zge7TmqhCDLX1YltVnk4RgjO64OQwaiMdavafP3C1
qo6g0j/mb/7bxY9xxLe4dxNObk9nyU4HsZVnyXoTt7b5KCVgwk59BHswEE10QG4dDmX0WyJzlW3q
5A7IEL9LYTvhY2iC7RpaESmWnmbXZ05Ajj1IPz1vzUjZaWK///kbVpLVRZ8N/0MQLczsYWjz79vs
k6okump58g44JsUZ0AEmHUJ7H7I1VbpyppvpRUE7m9iEMFVVWcSxDbJnweTJpQTxs8DuPFiGWvuB
V7aGwPaMSXjhhSTSHhCqlbaV5vruP7og290P/Qr6xejEUNkzAnpU1S2EEGEoDNhI6h+T8dCHE+EH
EZoZKM9RXU4vA6zcwVIjNyo5cXUujr86lRkWneORt3IZ6s4bkdD9LVRiHOjqBiXUESrM54Aj7z3W
PYzOmQp/JTBwoJ0nup8ttq96fmOj/IqPJut1ywwzcvAm9qeqDxi1f0aebCZIImjcrkDdBRIqvDNZ
AmAEnpXaCMZ7rFKH6oNUa1sqLo9TjhKp2gQmANpntwTbKctIpz/FOsYvf3tDPAIQBmY7iyRKZMui
hdZ+2Y75+WZXGPlHSbvAX/aWwDLvdQplHjBUKGRKmoU0N1GrAz6c1mu1mOdjgJGrGgFCp/yXfUf9
p+fIVhgbqvzo7wQyUtOkn99yykkRHZC68MDkrt4t3xNphob1RbOGGFmYIoE8ePQnVUpNmSPV3tIj
4kX35JBAtwKmhc/Sh4rPWewTSkWQslr4AapFveqA8xFQfc/q8oOXAk+xM1T+ksQ0LaO4znxFQuKt
epkRsfAIHwna9e9UduEzRrnyoAwP2Y6K5Rgs4S8EbOfF5rLt02+lukIY91J7vhM8Ds7oCk1dtPqA
qmV0tVGHoMLjwcKu3WupIumEs03Z/vIrCzc4D2fsUHvV0UT45RypUPbFKvXXrUTqoEEQIrExDBzV
+yVVPVDHecueod3Az/NNXuWHTYmFsvYbM2arZFRflwBHW7TGToE2GFWdNUk2EOMcdcIwXTDRZX0Y
xv82SXCzxZkVQzXqo0vU1jUMLxYR1nisCOHcINScueSz2udGDrztTc2tWgEdO9qWsgNrQG7vY/ZE
C2O2PPYpCzuNVqOU9t1GcjBLkptUFmLGMhn0b5O2whnYSLtw3vu7/dQL0iHD/b6sdhANWlvgAbGo
ufO5HgqVg1DgcjLhKiulWZJZbSUOIuYmXcuEKxueFGe3/tau6XBzpfSmiujgiPBF5hf4VaG+D6k1
3q30qsxht+pqLdzwG67tprm2JGd5Am0OAz2IzJCVchnlka3hjCojIg8ncA883VG5iDQlMb9TEnnB
U+cdxaEyVPcOU1cc8Lgjm20jIrslolaIYgX1L3AsasGaguscLQ7VORe4gxvM9pAUEN+anR6ZpSCn
UeKss4oWgG7T38mili1tyImkIJKtpuzjArL28vlSjrLcVCvfgGQ1mFkqYKwbyFzwy2OcHg5TIEDL
J1il/F6Bdlr4baSQKabaF9diknwYJsl2Kl39H53ub5nV8hEo+6c85VLtMtrDA2j7AyS7f6afL6Pb
Mv4KykAwBodxf7tw2rvT6td6qeycYFBIyAIlBzB9eYQ4DxaLCgc9PR4RiiOCJ6SlRYHTXoCPOp03
NiNJAkAlrAVBisqT7L0ypBax4c4dNepD2e5BjbEU7DaVxK+gp9o6ZzdRjREh+l0RmrsCmijelKtZ
Dp3fCMBfW62w37RrBv0QVe4WoVP51GVCpwferoRHUOWGuePalrYPZVYrZM+CetpWTdK6eBpakT/g
eDfBDiIjjriBGNlmDLf8CZEX6rjg6p6LdOyAWIWd2msYLAzH3wpYcokdWDbi4ESX0zA8Oh+YTUnO
Q0Qd5Xi/OxtVihhWoJ708IHoxml1hzT+g2rT4bGRLfeTQRBaIwRjd8etLQ3pZV1w0GY6L4d+QqQA
ACeWLQO80SVAFpuYQqz/hwdDIkSPOxHpw1c3EMjYFl1jmILrDvkpwt5zBiMlnyxMLNWHLZncbdi6
bfU+N36Y5dwZOS8bA+wfAWJF+tqII8LLx9/2IEOiEacxj0SP7qQn/cIyyicTLLfTVtYJZ384WoV3
O9WXI1Jz4o7uwMmfV4/y7Cj24xmbc8GeK3+/ZgyoHetRjH5vthEO+D2sIGpafh4eMoku2aSWNv9L
lmO/ikcKp5IC+Dpxz0m1hRIPlqT9XzvDHUQ93wfi3604wTnEGvpfQ2PL99Tk/b+oACmo7jUl1fqs
JR3Dlzt1bO9uhLIfeSOytxFvoZZBJhEI+omDmQ7DtKhPFgNiH3OuuRc6gAfSM3LAYJhZYVNuEp/N
nM4VCAqd9W+Ercpn0jMOTONnO6bD2OHUXpXUWqddb2EUHZiam/3TigGiL86mUe2yUWNF3004ssBu
oX22mRsGk2++PHp9Y5BvEJ1b5pa3JwE+ywFIJ5FJFvWTDexInJ66oL8G+GDUgNsNfkWtmgE4gMxQ
t3QoyNPh/qs9FxV0K/kyXDDUi8q/CFooI/fFyNOb2MZn9yqlw/IOzVbf+Mi5krX37Yy2Z4nqiTGt
UkB0t9rMCLl9zwi+N9BCB+3uhcafcbVy6+jDs0PxC3gDSHyPPOV624pC8K0WbAx1D8SHBZwwzWBS
/kakp63IKV9QUovhLly3rPfvlj9xR4b+hu5t44BSodq6/l2JRI7bEiGmLh8qcDYgvdIktFwX+lGK
f1DXyPla9p/Dd00QwcuTgEiQhqaMK7Yz6nh+oZrpf1mXbwwqGVUjLIdJzee6g4n5bHX77/isqdyF
E3nMyFIJBQlLev9qB3EG7pxfgH0bWShN3da6MmH+9c2PO0LeZY1ux2GiFmMOZ5rp8ZEePWv1xuW5
MEzs17Jn3yFrWDdC62ksJbhxk62/jJJMZcmXc+cAFhIsqyazlgGoGpQ/rCB1jVNM3SYyc/6fC1ss
iihkwJGBGj84RBLIX+zbwhY+5PJdaVRw7ghpVGwgl0fcmUHw4+vXPoysW+V9Js3iHdjUI/hP5LVS
Bq/5wpmC65NnI4B8vddZBX0vHTBW7qUBX2KdWSiOvdexocxnSomUrWH+qSOgKag8bCEkTehymhSL
6F5WMKVE6CvFdIYEdyFWVn1Yap7dlmKSw+Bd70ACFaeUk485Dbp5dtGOGUuY1py9fgZ8r3ftHnfU
4AccqQyHZVrtnNwDy3ZXerEVR7RTFZCy7/uLVjQrGJw+QwzJmmryTiVqoEH1FITu8Ml07f4aR9Oq
8QRnUiGl4rQMdb8TUrkQuVt52CC03sry8gJYW9YpToIrUQNyIv0vmuaGo/P7uK/9pa/pket5kWqr
PD3bGBbgTZllS+sJ9qrXk5GVc19CAmIKe0IKocDSM9w6qn/a011RbXAVPBpAoeQ6xOl42nk5sBTa
oHgI1NRAnbbAojGusHR1O0IdaR52SlwlNIPK47nAjNzu6khpZ9/I6XDytuITQybz2cQCVlyQ5oD0
P1sX+0eTnNU7dgOENHlZANxDJwzgQ87vJsb7ARxEcuCSDr0Z37+8cfIt0JRgvVjMxI7ddQKay1sL
Wj5i/CdFkDqvTH6hSsR6iyrL/hhFO2k6XULASgwocmnFCw6GhPzqNUfJtmjRiych2Th9PzRvxDM6
IKIsrXtK9jIjYLesSm6i55h+2X5SPfeSAqNpCJFQ7P42HzBsqdAlI7UghigGI0omj0DEbFouuibl
l8DJKxjQIsOG2JttUlsKuDYJ/p4pnavFsn3zwB0os7CQ4WA0H1ZsuKb21xPfgWRWpm7dSlypWkl0
cTqFzrLf+NhkUNKyb9NUxE2STTRoTPhOV7hsGfLnQgnhkYoPkjaUN6JQkJc6C9AEEMylRqMZ2ZXt
DziSXjKfOKLPhIvh/WZhhnpwggE/UpTYTFqR1smCBHJjJHttwHzeavwkZwUFJohCeYM/GVwT7yE1
Bm5zK2LauEZMZw4p+zQC0TG0fH39n0Wyvqi5ILJgHH5AfEcp3y4/skPJabhg4/4nUAbwOX4KTdjb
KeUb8FLgmocl0Co5/b+CcrvqB/zrEx5YD4vrQTqxMP5byandsDdKP8zvos3d2WVIEVXxMjzL/sqd
9/JzVfu9KM8imWWjpTLrBnQHWwqZc3/CFGohQzRgHUSaSxIbbYFsrD9t31dCZNIipruQ0Tvy46PI
zQfLe1WnONT4JYZdIZdGBO1zpDaIH6iBohEsMuzw3fvYVrM2Z2kvgWr717t+CBQCZD3KbOpJ02VC
e8ukIwRK1qC2LAeO1klxx9Xy/20wmu13C37n6aEJ4y35MObMaVzgpmv2DE0VV6DZWxbLvMq7lU/u
g8mrvYFIuXfrDH32T4rZWkkJcBMjeweIw9iEEjxwyuJ9ZgHplq6Z79M76/yAaopsr8rrgyOIFRNj
HsYBHsmLzOqFD1F5gzRyVwpx5dHUFcvaj+d3dtxqHvgzpt9Z1V4BU83qHg83DNvT2yZRKMruhay2
ovD3XHqShBZVsI1DhCQzqJG7Kijr/N3zRfMK8eguAiuxtydAwBW/xpkvbOlobQ3uij0racJ7u9VQ
GCK1ivIKAmjnLuy9kG5ZuuGfy1ZltnTu1H1xeUSkQPBfbJc0syKJnf9mQDVWr2smpPJnAFq+K2Fq
ZNknFk2Jwrk6c/Q+ybcOCzfNV3R8fzMo5mCMa6N7qofGXVAFKo6PYkctwkS/Lj9zz8P/Eyk2zi8O
E8HwxpXUVFJEA9MFACs8D+S2bb6QxfF8b4C4Z4ixPxy0xbde+/TFZS9ddmvanB50Q8n/wT6kn39O
vGR5LxNQNi4dOes0hVk/FHcm2oyZHMVXBtN1xKg2In9LpdQf2oOvBadFw9me4CnHkOmMIegwArWy
rVN2mZqrtLzYcAFy9PL6IyCFUKlMt6Oi4uRqaDUvXKTc6qv4LoThBsr0ReLQITz6zcFYdnWcv9AL
XcY/KLIrGtuhIj/ycNo0fIMuhxV52tOEnltpngZme5M3kBuLYkH3OvBbyo/7BbfegjJQEcl0jHo8
7dOnTQLO65fFITdhHnNd8terzn/ikhKcqv87My/dPjkOrlF8NrzR7zksdWgfvKYYqb4coNbY6QeP
nLbiiB6IWdWPCjqSRMl2bGPu596KwROB0v9ScfWhAaYqAYMbvU3URaWiNvxSRIHL2eIMBSddDWTT
diX2Q/LPz1qIUwRdOaAl2QX9zcGZMuIlYL8lVFWCR/uhZxnLp9AuqZtiaVIuQiwwJN8jre++HyAl
RxwFaPOcTDwWfZ9FXJa8jjEuUmVtgkIrJjZJfhrS8Ig2lliA7si6s2CI6iOvC+h46dUOdPDbn7Hf
E+iYTj5oc9IUUQZNs3zikli2yuzSztqyNROja+8R9HsYme1MVhnz31dQFEF/tDf7DfbqYBKJijT3
s0aSW60f6Jixqu8/Nh5ewUtZNEbjq2KTtfEs7khQWVT25sqjmyu1RPmnMgBRCOoodjNqKwmqq5HK
u0zlXPIUP72QV0Q0nzWHVwpSJY5xNYwQwEmHZ8k486pZKggmGBxUaqgl8OW6/OiJ768T6N8W1hTO
2zB7CcLdysBPL39VwMMe8asFLnzSatfT/t2h28n93Lls7Wo7JTncdwxSyWpyYKejY9tMNOPAxzBE
oOdV96fwD1cKoEow5if9Ty5dpP9XBlF9EeSnYT9Vr9zMg0mjrQGxW4Qo3vS5L0kFrp1iB2beUpbZ
36kQUc/PKDBAE2q9Nx8CW3vKLnh1y0+w7cWn0cLOZxpOnEJ4WKbhbQyAviBbZwCfxDoQFaKVLqg8
e9dvV/SNDvkFUuNyDajBOPNWeez3S1Lmk9nGX//zuDlAjLH7M4GoJViKENTkfa/3EqURCdtoYXXk
EQD8atDpyRHciuPbzCbQ0vQKriG2ThdxQPETsBDDaJ3cE8b9qNgbWWRNLzrLhLlgqAw/+rJnz+9w
3zTcWVfvVlWuBbNW5rtXNr184F3vHJV7F7kOQoEfSr5odFX8OiFvyKlXvXyMkeWY4x78Mec34L/W
9G5vYxQD42nq/X06Y5Ht7MvLTyB5dhtXWfMl8rd4d+yKa0OVtpnDSfGrYq43S4NXXMfiClshnXQk
5sjq92m5+o35RxgemSiKRrxQ8LcodcBUcsDXcqF9Xn7gCyCFSbs1VBIWT4Y+khT6yRbtcsk+skr4
Q5RI/jA8HzGxOFYX1168g6JxIk/oGG+r1cWgKi4Gdh+0Bw8/XQHE91YMWmn3/888AmHvqphHLrwY
lGyFa70q3dgqKR4SQ7iexMsqbxQcqxieWnJ8xcZz5HcZkKbTf9nRINPCBR4ghBMBxUU6keCAQIpu
F0S3gph/CP8kQvQUP7gYkoCzXkWI9kEI6q/GYvv+EKpd5ubGTj8x/X4eg73aEcvl/qOQFWMSdIHW
U8GhztOLdvyhfLdykV6/PLokx8Na0ApxiKY1AARImHpy/yDt42NmSCGunnL8KlEvk7MXdVuqXGDe
QIe3aCM9Pa9Qac4b0vp3UlfAdp1Hcn50VnOzXskYPh1Vv0hvETo0KKp0rNiki8Wufig4kZN0DcWB
tGIXo+Ra6N0Zb8ThToHqClsIzG+9Mb1Xq0Lw5iDSrZkp/IM5/LARe5S5DHpFKOvGYjuvhEUYq+HG
E8YOJNtH0tbT+6Of2LDeArLoOLKHcfN4EaO865DSxYN3AvBYP1zpllsVCOXWPIQB0J1RYDExLpA3
c5yGgQ3VDQCuvgJAty0iFzZqRyIPFphd13gI9EqYYTCyEGnD93ULtYJVeTLq8bKRszDZU57+zGcj
kVPyhlNf7yytNXnE9qWOp4x0ZmurAuzcAgLZO/CUj1Ufnz+KjJEcDgxDQU8H1SlJonohd0d3USJz
gihDtjkhWBg7iOM+cnK9auUbwQJwSum0tI4QkJ0wQ9sSx6+2uAr/IAdU/R3GZ8Zg8ipWRoSlgrBs
4EwbjjyX/vY1tPyozI/VHyOT0ZdbGDWxvfwzEuH+nefxyCmSG6bcl01sjw2702j3X1jm3B6gIUbn
rywRmQl4nrF3JWGDVHWWlhBxn8bH47wYn7vHwN/te7EYebHTEXcM2iwbhaJ16QUCqGWLymVwCw6+
0CXwxl9YKGa7fkUrSi/YVp0qfu0UufcUJeDANbbGezozj2X5SuudJq3gvHcEGtBNXqNFX4czFx/V
NgX39ZkJdyfEFrMbbewE5h/ydudqvrxEUEtMBauKopS58t83B0dDVxx1x5KvLTqWt84Pr4h3/KK5
IyiIpHlk80/6wb4TXgVJm611W6SgmSeWT13LMDyvQBn9BkngIwOpLv0Xv+JdPa7Kc8sH2BYPh4SG
ylvyEa5MMvvDUYxj+4SfB9l1avQXqCXee2oKn3OLntO6rX7QiaWt4/DbcM8dxw/UidlMjkosQKMm
0p+B4LYT8bLWtWUxzoXKO+Si+zIJHgus+uUtFa+myDQzaM/vWI8755810qN7L0JgitZefodDQ9hF
V6eyU4AmChmypmGCMaCdrCAv0y/EUE9l6Y+yU4Vx1I7nShtw7vuZjL9RH4uCIRqta8pXhRVgZNbe
16G5tlbv/9p3uJQqvvtq45+q5PmmJA0sPtWHlw2ftc6RmY6OKRlJN4wNijpdNtrPR6rTNOEVphPp
OGtifUStfWMhB13OGeKBXjBD1k5u9U86Wjt2QILLUi/MeE2ssRJflt0tAqRzG+pdi/Z2WizubXcw
WT7F3tO22Lf0eL20hSqVpHwTWy5lm/n1XYPn+OR5kBn/pxrDs1zZ9SZevqOYeCanzCLLtfbl37ZP
HyluVMFMYaRaDaOoPnXOnZwstA2PoEBOIFxMp8+IuatdjjtliOc33/Ix0lZnlXJTPvAX7U3+s8qh
rjNRVcN4baU6VfcfrU7MKEOP091wpyrRMM3eYIgLT9U5On/Zci/Vp0C1QmJHV+9tJJ6rH3reJNJ0
r7vJJCis6A3UjukJSsTnGzWtKK74Ml7XRmCgVxf6aYOeOSufHnPq+nlY3DtyKX+U49/QZ6Y1ws7i
BJtWg1sTjqz+CBvidFhDaUQY4Ijl7EAxGyHVAPOekx9ourpC8wMO3+Bsy4Jau8pM0KKZgPTS9sxb
R1oj6pynkj8XjsNeR8Twf3nDluRE72QfGVq9xbNwgPJaMPf1xHXwoQgJd6LGVXxctYAQ+nteRlq9
VAB5z2vks0fMrmGJIwvHSwjbOwtLcqmTTD4KctQNuV2dijtVW5fVHb6NMXtwb8fGBXGr8is4LVFO
L8PW/T857T2B4W8pmxCedqmR8SHEgGDCjvXwGi0iDsksG1x1/6oOc9C+d7g+pVHLUyucxcwiE6VO
ARcGH32yvkSdo/oOnMGP5IhvGLtm2aJtqPplYDeHmu1GJKnTmnMpbpbrDMChsj126wG1LYHKMTo/
CzcwDieMvtTxjjlp/ehSKphSENzWdVy7/AVG5FkGYRjQ8Qk2MR6WRBMaxKI0AWbWt+NtaO6zDkEd
H8cX3Ro1xr4I3AyMt3IWRieW3LiDzHw9W9r/VqraKz94z5CUf+ERrvC/Sm++Pi71/QurRUNl6rSU
xwAelJuT4aD4ctpF58cDKeyDKmYWCa+bqOC3X9Typv4SJNdkK7OYscDp1yL7lzmDFH86/S4ERAhs
gL4CJaj2jnS9eARvqLVbsVEw1ksjuy0DQmXhvXNujlS6mL1+gVWFaqA6S6SMWF860QnqYaqjVK9d
ewpr7TLHahxXsL1Tupg+sXpcMQ0hBQT5g0PUTxW1gUs/9+nlA1xuIKY132K1L24G7kpKL7YpFF11
sLsL5Pn27dgXqqBH+5IvMeRxwdyoTTTvmfAEyMz5KwGpilFxCkb+qNWwGl/TRhi5dBWbiW48XRKf
eDIzukphQcr9vQXL5yrXsnaMwx+buGLJ/N1K10q+ZzzxliL6KuDvSubvorS4Zd5+Xf4w8wfCEc2c
9joKYq0738nlffKlUOyGAQ+mL8h+5hGgKUqEOTZOhMJzQl81fsbPJLn6YdZHCe0xh6QGD3C/nIlk
2AZrU889Vk5DF2AhKplx7jCn2XSOZ9kEt4IIVTo4l3QgHFoNNtPBNVRYwAc6h2vhFSyI84DXjbZk
APoYHGs4zxr+OIarsIqd+UctIxBSQRfAJS0rzsEIHkdNdYHzZYFC9LfflIK9cS6xsRZepi/FT/Yg
g356MJc5AHSc70vYv6Bg+s51dYxrFgCpW2Eb3YNN+cMelra9/zCLzeE8IY4aNEX9/o+I2mWaPwzp
CAKMWaZXfOKBqQvmmXc/Nt0lH6JzBEEUnq7ilvzIshOab6VywWo0OZwVKlaxeYVwL1pbOKv1fq4a
1GWXt36sPbO11kDgyLZeNi6e70y4AnWFxstAowHKm3ipiU2jPtC+G/yBHpsz74cBlqCW3by4//qm
bM2pt9t9jMtZtoM6089WVsp+oZ32mpOgfCYV3g6nhJgtx7Nar9CYuWYp0sYHERQim7y270ntySOr
x/bmI26K7ISOpLXKCXH08/PDxuw9y//Hibd9r+7o/JykPAQkWWDGcrxMeFT6990Cv7og0awHfPls
88n7wWMUgpmYqUrbyronjuEDNF2/bv+Vja74jc0arXW/vQbM38Pu4FAvYYqfWxpMpNnvN7/HMyCB
n9+NmZu37f7rV6vuETBOmamK2ncAonSX8+Fm+T6jOxLoa17yCw9do3Czphn58tTfHjyTwL/YjzDB
XcKAsBHJoSWxU8KA/PB2YuwgG1r7UcMBwkW/QyyQYkbzEb9MPOybtjm3h7tiAGd/86y6xQ63WfU5
crsAXhGjAtXzX0R/Uo5zMNAJ/s1hMUcax7CEoDbp3TdCVUlF8pUVXkBFk/ahJoKG4PZbQjtVcHe6
2BFA6TszHrfGYO8NUF9Bk466kKdY6MwYyx2xqnqS2CIVm3du6hOsw2armBhy4LjJho7xLm64OpKk
CyQOUsW5pRN62wacXCmpdEKkkxcbihOjyMEjvhI15rxHAjbm85Za+3WEnAzZjGnJe5P+JjVKplyG
YjfEpEUpKEITg6MPwThpoRA21tjoAm/FwYoAEc1HgR0n4go8QXhU0TEE8uhabkdkLWAZpevD3icv
QKAivuiaQZuvJPNadsvXyicGYI1JniC3BbTMk9GNg8cnaob8RKHmFRts4GEz89hBBooRvFtp+HW5
pDr0ZQOLZtjXcK5SVCOFY1AYcg6mZN6JH0hwqqavN5slo9UtYFzQwFIM945lLMFdfyPvVTcT7fPC
PQoJft2X57aKGsV7LnqntPPqegdSmiX+ln8zAhnt/tn2p9T8VjMZVH+6tQUYsiyg70vHzlqNjPaK
bJIqZDFSBEiZqUE4oFZT3ygKsQnLP84HCJwwi5RVQknJrOGo8d0U70gBGzV/rSQPpBWOnujXgrXy
yy+S74z8hRMHU7B2VaXP3ONXZjwqVbe+OqSeDDbAAuzsujcey21pQHasrpwc2JjYTGzy4aOzo112
W3EV8/XzOONXehxH1HuXmHAf+cmrpV3dMvOCNxSCPlK6qGM58HlUQmAj49Fnj0ZdPMFjuYPctmMW
jfQ5GW0/e/UrRiXIkuuEKMvPt+577wCidBJ75N3fcsd+4fcZHL6RfOJxHHsKe0ymkb4v4H2ZIkVJ
AVKRS+AFuDpbKg3EeQ7BAH6hRkgTL9J8FRmrr/Wp7biBxwLu3yofwqcFumiBaR61VcOCFiaDCcTR
B1I5rDnaR94NwA7o6KPlTxXGDsUBk3h5w+AFwXevJT4NJexpkSOuMEFpv5SsYnbojbch+3tg6l/t
WQzzJzzdogHJCquww41D+EEgSPGISbr/leAWx/MZABHKwOn9iwkXdUntAoXRpLteSEmnLspZ2mmN
g7x084xOmP1Pi0K52URqbOHP2zGCDlU7yL2X6lBrs5yi5u6aPCXWFExLwZzya2xi5Z0/UnjVo0OS
gzNbFBhJCutMXTtH+3xuPB6Wn0UT4MEXx/X2JTXJ3jKrGYJVnh0QG/om1bm5TVtHGn93fiDmrWAV
BV0e43PYSxtagbuZ8Zs1GfHAJyfDsfn+cgjXRvObrc8JTN5SJnyVp3DPNlgG/eXdGYC5UpdOSQxX
esYEZAtLPKnoi68HKrWM/5fvOk9nAa6pKLvZFpTLKiipU9KC0YaQ2HN1FTFSiOp23I9higd1wUBL
yTDthxyOMoYYWkg0NIqm44FYZ2+IyKXhwoILjMUgZPbcbIXuifkt9lGliuXKVfFFHBhy1VsBQg2s
d3Kw1D+5+XS//LtAdjTiR7dhHmrXYnhmF2vOTGszsYCI7cQ7quFsx79HOaMgolCKgogtNNuCgG62
GIMarW+AvNvtaHl74wSJq0ovu94TCvdhoUL12tPYcTn6sWFAmwidHm9UsuBC6cAJbPx8u9NsSH6j
dkAs0O0/neFGUwr+GPyDSUyHd2oX1axPsYl+Q+JexlyqxZQFHUYsV//G9+6UQQxZNwuPEeDdnlG8
7+SGC97IQxvEcT3NtPLGo3H2hWbLLhkV6rnFdbuCfaAsNgoHnXEJiExluSvAGKypBk6PKQEGe/Hc
nStF8sOOsEBA4Fjfhxj6TzvYUZBlreWYQG5UdZChvnf7IrZALPDg1LjQ6MAsZRyYLXrdjDOsm629
8kqq9/oU5pFg4ratLI90+dtBnSv6SzOvfuidPL099xxmBc+K6m7Qcf3nUPEpLxQy5lxxIXQyFagc
iCrvSkD5oAe1vraWb9C5Y8doZ9W2DrfWZ43crigJ+8rdfJ7nyhJH4v7E9Z00NgMKDleHc2c1NI2B
1Sfn8u15yF78t2Y3SqxIqUC3PadHsQpVFtxKroQKxt5RRc0/nq8lBr8VST+Xk5cKf4xgU0S8nbJT
qpdjVRf2QOPdr0UINxQVUo323ahwYpD+kXKzCzHkVR2H6JAQIX51spRjXywxkMotuBFC/AMYmymV
XehLCuLVv5HPOk14GQ30+UV7mV9nVzBz9szA5bAFB7nJuur+YqRgteXk28TlGu1CALk8tXXFb9+z
qN9Wsjuso6KxCTpZUCJEXlSK+JjJGv19nLsWFSxs27E+RNsayWWBJ2Lcvhq+cKYgwZQh4Q8wKBa+
nGJ5U3JQvwaNe+6lq3uIt8PCbuCJaey5ozywuE6H5qxQ68LKJTmVWX5c05xEO6k42s5l08jaZlZ4
UrmcJJv39XMleJN0Z9Ky9Pj8QMkJiA8Kj/na7CecB0ysal7MyZjIvdwr9/eotFRg5eTQD44wWp5+
WTp7UXu5Xse2Ky79AuyksA+iqzrR142vZ1Huwm/n1iol7/3bb3MrniEYkUkPabbTUoZASFkum/2K
4kF0CyT1Sf+1KuU6F5gYX+kPw6h3leclpIcuKNk7Vb7GhxayBpmW3lmsxdwUPoT/zeps7vXk/7DN
qlkqlaxAi+SMuPAC/P9oV8YSeOPrshmpoAXOKhS+rQcOvviqRzCC4QXZyZipLY+Fhn70NFB3I29c
JPFR5Y+ubUP9+b4vDxUm6lnkcUdHnGO+dXE50cvJxM+uyi8XZPG1DBtWcfSNFGOSMSDECARcRxK5
e6Pp2uwYZkFsCI1++167rbAiaPv3roJfIftT5pJQ8Io687oM+MLMm0sAA0XhGwnCzVM9NugIymZY
C/q2CGHDl8VWWjp2bLn5Fu8Eq+kOlwrCiln931VExfqhzJlpLnI4/KkRFC1v8+4epo6SiH6qTxHW
Ct+j2ElZN3KzKlrdRuPdAgmg0hjfF9tJEEzA4wuPFprogjAdp2Kx4omx1eoE3cRUOE7lVldnY2Qv
Bf1dIARlebH9HCENmOvrxseFB17n106jA9CEN2EtP14lZk3PN4UMa2OOCHBtyV6ojrJetQ7+oQUc
uGMpt35VUL0Rocqqfcrc+nI9J21W3sVYyCz26C6YFgHBWUV3xs1o7QojSUf8ZvnnYSP43B5HZbaE
fEi0QKpVq4oc3et8xR6+5AM6TbsGBEkDWSa+9XUqMyf2nWe7DIoqmz218LQW7CJN9ieSUAI/yqyw
zJU/cU7TzPhsIKYzSOsdN0cR0vc9X1qgDvgCsmI8p4GDfEFY/pF/fks2EvIuOM6/ftx052jY2o52
aZ3NYmEyWwUx+RmTdAt3Szqt2q6tpr054pYQx9N40NM0wLUrtMD7jo21MhkUbjB3DET7gURAG3RQ
3hDBYA4RQfB0UbRl5htwARGtwHDUOUt/n2TMzUwmRX2gOwk5QNHM5osZ+CDxeNkr3Plu9ic7kb/Q
XCx5Ff6zaA9MiKShHxJ9Nt7TSW9f7zoP7Ksn8zuTabxujb6H7ZV1iqGIRH42dZ2+wLMeeUkadnMT
YmG6EkGXRml+euHCq88ekY3p9lSGmES5W8DcKbCnCZmauhU6ttwf3rb90ET0xU192oGmKoXKihfw
8+WstNDbZtvZFIcC3yMrMmNL0EEGQt/WpPGhCM6uxKVsuqru8kXcbsxnLzPqfgZ3+GMRRTjKsyl6
f61ONUYzaXatReO/x4B1QD7bEDgOkus+j2Fk218UuFA1EbTRzGP7IRtvj6NXegG6/amllREhxTGg
MlEfRgtqQLEWku86o1TqtGGv/wwoVSvFZV4DJq9P5lfjVdbegWEGnLNZy2jja0bLhpBUM4umSvpU
viQQ7otSlPn69zEAWlxBwFYmHwzmrk7YIb54jCN/qz1tx8cyQK9X3A+ydurw8HxWyPkfjZffc8mL
0a7C36wywFO9lpurou1oAas9ziU1HLmf9XtXoQpqjW+2eZ59UkvMO1ECciPByEr/fYSwmGlmvqY6
2D2JMabsw/e20JtVsn0Pgty2JegRBWpqr0XrLI+Up1YKU9zhNJCp2cJLv1a6ro1vE3zLtaDowWTZ
BiJCfw4TbMNPfB+npX2bU/lKE6lngjBPikOGceUC1rckL7s4W5zZit0QBgLTMao2VofWoyUbkFu3
IkjnZfyJim1ue6bSmZi7j336Km4BmldM9jhz5jT5zT/Axup0/WaPyqUx9YX71wDGuLFCn1En9tjH
mvNyoM24cVxo2hOxTGF9DUyQkQBVJsAZxLNfXiI8h7kp0eYkPW9rMcMa8iWYO08D5+JS4aLl5vsT
odMdABFrEEn82zLTPOHVu5la/QIrLwk3DY3dHp8pNPXSRnoIjZ7An277KLhByBXZk26cxVZWwqgH
28L/Skx2k694q8xAKpmsGevS52wOPW/p+3Ycr3zA07ZT24PC+Ezg+cjpIHobnVmiJsYwLV/yCGXZ
0XurlR2k4SF+/4kXech6B51g5WQu+No4d49WwV2esJE2ZY8RQwYDE5EGX4hD8Ah9kiYnJHpzqo3j
sx2x4hy68eUOD/Lz2/pUKhjt34gUYzuMS54DZWMLwC6OYBeNXEIi8gVi0HQSwCOwy5nZ28t8sGVn
AA8LC+LOuiHK1m6iC/Iz1zPhb08X2LVA1UKB/Jb8uLB3DOwU+nfH39vL3xqXyEHwZwksgFAqYEoT
gPIH/KG86MTaO6quy11yLWPaYpPGi4jREi6UHen8tWVC8/LKExVK8Oh1ZHcgErk12HJVzFRLFH2l
zoHbgUZkuFLyu64hXiD9lXByleqFEVfGIzz+AlcWII1O9YS3StGc931T5+qKWmoBIcfPKV1QTm2Z
+YWrqUFLqS0/wVEKViIqodHBKbjPUBlWdfUDJS8Lae0cd8GG0dZMIYf9jCuhGxvoWuhaFRY6CecD
HMnQuwdfoA7JeILycqMWufVctqC0C68TtVs9mi8AIg9ZtN83nxJgIHRtIA/NKpIvGUwTWlZm5IMa
yXw4Zv5vn+I8TWUDEmcQI0WAnhqrKDqoATqwS3zXuK6jVSoXejvanKIOaxK0bGWE/46XXZLRj71m
BZAVyVFziVxtLRgwPCYq1cm+3lLZ0KSqK7hWBK5qSqnH528O1ajP3zx2VrKOWA8GUMdZJLW+NIIy
koZkzrsu7HlMx+388QWyGd5LcxRvcIRAyJwbftsMycX5CZtib+qYtblk7JVwCFP2lMTVi1+s84Mw
A/t7nwNl1Yns5FpS3qTEhKpajDBK2F17JMawnC10BZbpNpvmzBCutj13kiM9E4a4u/yDGpDa1yGX
mqRKLd0PqmBg82uRaXlApbS4OgHOee1OsBp12R0pt7/0Myp0LqhdJ7QX8nw/5xo+xVjYRok0Eqdz
dK9opR70jnoeMHaGRLrVCS8ccM+SVvGGJbo=
`protect end_protected

