

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Cqo+FjfIOIw/0Kghh877RN5JtWmUPj/KfIaTRt94dXWp8zshF20HfBCWrK0/KjFcQ6xaC5bYfJZ4
kTgDE7VoLA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
P76DAxdsqqBm7Dhm+Xv4UBWtxeM3n7VV0uwUkGrQnJyruFJEvMXWtTIk68wS1svCurmxJblglPTM
AUuHl8lZTHelg/xsbfqIjFFpkYurRbfQPaEBBncWEUkGXitk2MsCEJd1XKoy7X9zf5gkivM+Dtc/
HmQtcrnx7yMmBEFf0wU=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
TS87/wLvg3wp8BEZbJFwjKct5crsKQKmGgle2kFCdS51Fi9lA3booRtYf7PKimLYtiDNKzFnNmDB
yS/M5Wwp3OXdwvzTqi7m8nPDGJzv9CPlgJYl97xwwfb/xlITgLx+mE3FLNjQYh1k2fW/YeWIYcJ6
dHaLGRiPpSzATplaiEnfWr4z9y5Zgw529sAAgbJqopXb1oauD9xMSn+2U51TKQlk6QzJOyaBGs0Z
cYN8i3mMrSJtz9+1CorRnx9v0S2lY1WHtTTmGGV3GXP4WDMI7lTnhoLYTdqSlyv31x9qhFidZzgn
WXAPS6oNxDavoZXEycPxfYnQwSx2gi0tzG/NZw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
NpAOviX6Xvaq+L0foSrleTOrW/NGnS56aJ5rqqn2Dmt6YUNEPYGn9LoXqfbnr2nu7OxEo+FueCzR
GTO3m2J9405e67h9qARcSi/hF0VUlC6bqx3PVbV+Lg35W+tGaz80NE2OUHws+A7UXDQk1Cp7m/EC
XxMS909JUlXKjJHNQPk=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
P7klUwNMTreRZK7TaA1WE7CMMEOTtEjomJfZ7pHl1XNp0UR69ZqgBrqFP7D39H55daou+YH1hnHn
RPI1HarNWCxtLMV4hOqf8NjoCFBgrnnB0U1fZ2Lr4Pjyi28WQhnjcgxXDHuFaQlXuyVOq9XUsvMJ
ssrZQdiUjtMyy3njm+Pnbmk63891Ob2bUkQGGCsGTzQYYho8qCUxVS8K3X2BjFQusmuscPspGR3O
NvboEcmhCLzlJh3n01BooLiI/MFAc4YbNKfLIovvQV4EihZ5noxjjP5wWP91DT3v8RKOECGo+vl0
XfgG1PKzgtiiXSw82pyP+WwelLF2xj1qh8+H/w==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 13728)
`protect data_block
CMGRPzHJ9vTJBzRYkmsN1wFwyh3pwd5Rs3WKcyEbBA5GsXj9nhT9Sj6hmgKKDz43hkyqUqs0clz8
CWowOToDegbbCot1k7SVWUKpdz43K/Dw9bcSVuJML+iy/vw+gZ9/suWVAYxTrjRQki7t6dFOiMR3
7u2gOu5o8lz1WeK0AteJjeizqfR9NUYiXhjEMFuU7gqCZt9H62JWiu8KBhhW44iwoNHkWfO1c+Ht
1X4aHqewSnWYjBQafPKBSi7ULUQLzNVTNix/V2BLZtCit892uG9LkyWAniCOxi95Rc7K8RabPAk1
37aosWfw6aHRb32wOj+N3XkWpyNDZvfPqG/pug0uz8rV6hecbseURar0t08qYdE1hoaaksw3jw0a
3/1KX6LFbIjF9K432s5MJw+yUnKE2rlENQq/qW6x5yJdQUOGkO4Gr91OUhTUMoEHYKMEZwkXZbQr
8+Lee1NKJk3WwDwwrNPBcfVQYV9WvFJGjWH+OzsCltzUFRS3OflQ36tg1iuhtYIb1F1htYAcu6r+
KV/FBQqKKDC47y+CUw8vElujBM+23ZB+9YGH1NeTd6LBcXQAbRILsLQEGWsUhPut5lK6PoQeSv4s
p8WKJjW1va2/TmULhEjs9MjWM+hlJg1/BmtpEu8nXcOp2SIBGrboELu0FNI8nc12nOkxILnattt4
9TpN0t6Sfp49G1J6VhkTuaTA7uPaKd/GKuflTKQhmxb4oTMOWnNGuo4WTGOb5L4I1XM13v2qt3Tn
aDxN/CFOaLJOwgM7w/QdfvL8S7KMlc1awkT8ZbOD7TQM+Xi1ZwDs6o0GdRShrEeIvLZEKQ6bPwsV
9jMHTZxgy/C2Za0uzFyWSSsBaashiTAbirOEJLHR2G78GaOw2DTBE/xFAbY7dhQNFv8HYD1iCrL/
XGBSmv4P4LBi8xR2cIOeYdsiv/6o4yJEUCNYRWIXJfoR+NVGiluS8yYGAkNBnfIKNvCT87grZ+uG
jeZJdhx1sXBxtK7EGleahGhlLy0V+MmcaBf5grnSjSV+crAnJQTAW0hG6t1UhGbvx/upRrJKYQKI
Gg6cP8VebdaM5tKuPlCLjFPPPiVGVylgq3q3TOtQshAIVzNpXLllLxF4oz0T1iAj96b/55JmWy8H
sQVuz2PUGZICtifunfD3wMqVIamf3VvOneuiIS6RE6fTOgOSv3FXbwdfdpKOLQ6fvQ2lDPrgy67H
lDBV4HKRhLYW0mP9dnxCseZH0emjaAjsOwoj9HNMT8UAnbXdTWXcaZOx7XJd41NJEu9J8G/wHqCL
QCWyHLOTo1cFX6agFhJZ0I/nbc8qOVASIY8Lk44r0i3xYyQzkaGdYC1+RNYufkXIoZWvG0FdmS1D
C6K72+fbx/SSpVxBM8lLmTKysQzMTMT0EOVbYpijxj2+fpFeMxYWz99F/13wMkfLwn8kUQ98v3G1
WwuM58v8yy//ZMTDmOqyeRtNf7rAo/3JVsBBA30Z+ZCbxc29cXkB1lnMSUn7970K5ZsHgZuq/bfe
9Ks3KwvirAHfXBXiabwRh7kjvPAPBKrPSFbDV76hz05l0oyFUtOctoK/crC1/zPuKPeoS8Y0iRe9
YRNkx1WP7f5acuOJ1kenL92IiEDXoOX0WiRxuLUn4H59J20x37dSyO2iBzewg7tJwGdzbRcfe5fa
6T57H8qE/J05CIfuK/apiiOf+UQwAuBp0Ov+qSmC/4yiWbDE17MnBX4jmavs9YnhjUNTKS0FF6wt
YZjRzqKfLo5ukVIKeE542FT8g8gyFR5vXp+jwPw2GHG0IxP8zHyeadNZ1lrqqgTGrIjjZAOn34v2
biwSosGtpAcx4Nu5p8GflQE0KfIqXnXAiPLWDDmEsWWgtQAjj//ya0GJmb2vD97YIgXsBiJDKmVp
t7qOYBszG5Qz5FSZbXBNHki4y62FuPPFgt6yUtJxwSXIT0Bg1mrfXwWK2dZWzXqGzVPHAezqWC5d
iS/euKOOD6HSOnJKUpPjomsy8DAdm+1tlbhko9DhimZkmETxJ21cnnz+P0KbdDQuWoilSYWZeU1k
KrFM1eCPNi174yGWpltR5rFF5j3EAQQHD3fX/+U9GdRIQnvHWJ4dQVUd8Z1z+aRNjyKXNrzzydNf
yM3Y7SBMMU4vDVkWGeU62Or2ucPVP5qiHCLU4dErtW62ABtLBTYXwFYrwG7sUUOKb8wpvFJ5hH/8
UyfeLRSF1Tsejyxh1U1KWwUE/IpwSLs1fSZIn+ldrVVBDB6djtZ1uxLQe7bmeHrmtq4xxId0y4O5
LAHvOlZAd/GSRzNbwmCPF8yev13H1YhkPnvKUjq8ODxy9pGCr3NDl77aHcd+ZvqJq2MmHV4YHTLF
FIu9qiEaFx9kUQwvbtqac2/DpaXHeo5wzQj0qu+g9flVpR/FdO0IV8EEhU99dQAZiv/boa8nqCyG
gHN2sopEAgXsUTfvvLGicN5/k/uOaDQvUc7qGYe/Z5ckgcMHmFto+V0XcUEXxydQE20DVS1Nb6wV
fIu0+lco/AM/W+Sqbr7BIjEOd1lPgWsO7TJTO/Gps8P3C1/HdBxLe6dQZm3ddkjJOLYclxYNImY9
Ma56D8dbk5xQIMiZ3sAFrIH3bJ1wCUUAm9uz3ijJqaF4VcHaa9v8vYj0tk47tBMbsayy5nYwHWNr
e+0zH8C32wBpEpy3M2yBvei1kknJkcDKX+B+VQSYrxVBfXfOQE7rR0Yojyvvac2i5utWg1QKeivo
IJgfXwbNhKFGw58bqnEXkckKjKbgqPs4CSYRj0OniCrI/vM1gReI4pFEsx1PdP5RyzEmqQxb1Q2c
BsiqDS0PjkuEmkC9MzlI6VtQMN/YEKT65QpR/7aWbH8egap35AVDteb1rQuh13IQ9FV2zVBUw/Vo
A4dfqx9nFe6x8VeH9Z/ZbX9Yxb8aHSbEyGV6eaZiuteIJYffeUQvPyr6e9/3kszONg4qKzdldej6
nnYlzkg+D3i4SeFuhUTesidPbt0s9Kglvx2J6MXgogCgkQKuSR+rYlJeeQ36C9rQXZwlLGTbjTCe
9maAEHTZXkqSTJsA3+VTjjQQpWMKQ1bGhoaNwfbuBdxQZWaNJF2BdxjGz0bzpQuR8Ec5YGJtBpLt
YBoxfC54fUeuqWuuFVuoiRoF+GTCXPaSFuba5O+m92LsUtcDmFSHwDpYTpA6grzj43LXGmuctOnP
MBWU/9uDZlTb4QWK/WqvnMmV4My/PoBdI3NplJgY8BKdceWScH2ICYJxjwWpr3tbU8EUAQZS5zUo
azxFg4kkYBnzOGJr4a/YdSJvEY2EUvYqPUL539T5HmRtLEDFvQxAA+Gc38sLrzZbPSc/evLwNogV
3DaMdPW4cE2Um0RtM4xze/qmoaOA9Gyz8CUn4sbtRSCJvt8Zl3qSAgazolxa2JlEMljYjnGSD+uT
VR0MLVUQwc9cgAZFdDhJ/3t8OAOOYZnMdhfKuMiaFiocu7ycRcRE9v3AJUn9GcWACN4hz2aygM3e
WlvOoz7ofcQdmyRm2jpsWPYZ7Kq1MKxoV8RGEu4wVLxEHdZK1hDL1rNfOA6P1hvGpJbeISTUybiU
qNywmB5TZdLCIbyt3lF53LwGgOvfnqLxR6iOTK3HWXfOS/FDTS+BllFTS2baEDVYWtkcoo9qxQPc
o5DwyoD0BusP2XVBBOy2SMQFPWLtw54o8raIHa48QDacLzbNqVzsksfsVV+Ik+muT/l4Z1BAa9jU
WOmyOYmze+6SHQWKsz+COp3rjutDcYa2JTApfx8qMknf9qe4MR02bQw+qJ/sszI9fOqrfkZ4lfuW
CdosZDlbLufH5TdhIeqzgw8QbotR2cl3HwdmGSdHQj4sMrdzX9ZaAB8bmF3quSfTRYJglW0ZRW6O
FC9K5VTD+IHHfQWoQlZJGAxHhS1VOqdetobMyO2Dh+X/NmYnHnKvoIDNc+u4+7ShkXzQzR3eU7SP
BCQVycd0x6RqJ3twY06pUMAQJj/AlXKdaKvQR5HH3HsRNFTPChmpU96mXuaVh+bh2/EURtvtBYZG
w1tWILNmuuEqPo7fi+iq/35pteS+zWYsuCs7RXulStBbLzwimIK44pyjILHuXoZ37jE4FPs6PDHY
D7Bora65FoAuBmSkjRFmxXIt9zbbE//4ZDRw3cZ/wlgy2aNy7e0qdFh+ndx9sDkg56Zh485mC504
/C5SvPwDlBnTUIbLiIQACYmBDg/WutJrZkt+9DMu/Pw2CWaWwWwKnO8hPr+ia6HmXNddN42fqIRE
UUbPb0i4Yc1WeymH/Bt6dddEUk5/A2247KyASbF9p5JoPjjh4S0p+aQORctYh4u/ErERXPbBg/sh
50j7XfTnmZo+NFgbSAB2y2IC90ku5Xfb94Ph8KYe+cu+dN9/ut+Q+XigVEiD8pZkA9SZuGoNBcXK
KfFxmUAizZKjUqEWM6U9ogPfGRXWY6WixdJQU4wQJDc27sk647++KJFPe+SETxYkCVMKVkuAuqI3
VBTMl6fU1r1TT/2ccyXjGDPT1P/5afVBi/qkm6oCCetxFO1ed6NHCjDGzcGV4EliYrp9H+wsG5qG
k9UCNqZ3Ud5MiuN3K77pb/yWSzzYXdrylptKZE57AqeeUs2W6YtTlmbdX053KckWAVdt3W1uom3G
suyw99VARVowzrC0UwSxNEw+CsSAyE04RAOK+6Q6MY8qrmQC+ekbERDD2DTKNhm+N8GdS4dpf84s
lDzJ8NUkrAmjlf7LtrCvAsaa++wmjCWasfY0xO2fniK0NO8ZQdoG629Mh7zt+DI3dNt3ztDP/SNC
xngz+xwK0c+pjmy+b7LF9bhv7TYYPTOmeM/Tz9yLqbWJZ0WOWIuzw+qOt6OkP9yKKWSbDLkLUeZF
TEPsX8liCSQaOBodbfkzsPdIN6ZqAtWX0LRAoCwgKMhhmcpZXRbA3SgXNPdC2oipGl6/L7o+aKdN
P0xhcninl6KAW79PfHHspLpoNs/0qT8mRQmfGH+lJ8RWqjJy8TAre6pQkdkkie+99NIvBxN/KDtz
8oUP6xlAPYoQo1x40Ujg0UiAsCNJs8eLmd1Dj8/FYeVaBD8NVhbL3zyPDJYG14INDcJipvY//f0d
vZnGSApBCWyVVVlZQa9zFkORbmLl7Ji27FaQaI2er8wG1hvUpl8Pd6QbXy0GXs+XZzBqofmWOC+W
3C/Bf9dk+S2Wqv/tDwJdSH9aO7Y9LI03QwtTgn25nLcVEGuGx1MqbW7KlIIuxCtvlkX5VCRAGOfw
VZul2270ur4YiTiXOV6wg+VX4nSp4RD6hjD/1yethcmkIA867jQkenbXKsaP1B89d7QSeG/Yn0f7
MEXiP7bYujSz5v5VFM+/7t7Ssy+bsocaBZai460vf2P1wyToIAaaMk2KXnFEDNDCuZSJuEaX5MZH
zvr3QfomItCF+jH1YD1QLG26C2sGDBIBOOsc/qhdhWVuJ9LpiPe4EshlK1qDK0JatBuOLZgFk6vJ
tycnRSFotpcJ+kUU1XNUdDyhmrLk+P3E7Jz5oR8RbiBRr7EGauK3t4BYZP72j+WtChMj/lG3J0ba
EzV2h4dGFh8vTsuwPoxPWjUtBbrtxCDqFMM6mcZJEurbviGP5zptLAdleBT2Mi/qAwHu6jIFy1Vr
aKijHj2YbpVeNhXAY0fwqkLj6nachmDnufFHacWldmnaESsHujiz2oJdm3+oXCnSedv5qCLJnStc
CNWPOQS9P3v13jKx3TG9xEIflmvS1tosKNBMMOjXinHyQ2Zyxb/cGg3eSd7RIcqwmVZByECOVXlF
KauHoA3h1ps9qozKK7XYMPFQXPh+rWaeqc6YDMTZFsPEerOPFTv7Z3nyK50Nt3bu3UMi2Xb8rfLW
DiBZIf5iyHAQ2Hu5ZB04H8lVck9NQu+cxJLYUx0sPGGrI8fD4QY1gOnPJhUqac+onICX+UAXeCbu
O6cmf1u0WTb4vSkpY8McCVE8lkwg2ceNQ95gj+dN+Eq0Wb3eiLUdUPCkyhc3tAcCgGQH396NpQhI
KBzw+oNY2VKplajmFcsltqOEQJxPgQmTUxjHeU3PNcn8ZRHYvM8xmalAR6EjALap6waa5zt3uWdf
QuTfYez0njBEIXLdsEIap8fhY8aeXCExVTHxlguwX+/aosrg9Ur+8rVgX52JBtI3NcRcvBKMiQzt
/HZ+T2ef+qHBNyOHkBZpeGsNwYKuMiqirQrY5bR2GwJ9G3XPzcGxhK2FETTbPRlSDLf24j3PbA25
B+FrQwFmVsmQJsNVMTz5ZJTDISvzqLdPBLhfItthoGXIzjqCw65WRQc1vWKyt6TIIOnXj4aGW+Nc
FcskdVjgeF2607xvmfVEYuPRgQExSdII3IP3LTGLjogfi9KaMM+4Bhv0eKOKN5pc12w04rmOwxda
I/nH2OwJ0FHeoQ26kGB5fdYZSmLA3rX0dFE0wHaZvjtU0S5dK+sP/0kjTGAYUdSepXTxwG5xM9jP
oUUNGvQu3mF6GKREWv2lCQMGDuwUEloQixZnn/Uhqqvxzp/VQ4MZmfTo9aGkw0Q5dQ450l3QTY4Q
erny9Y4/SvQW3FIkoEH1TKNk5e4vtxY1F0DK7oPjlSiuivT2iL9GKBwdDv7dQi84UiNc5tyLzOz7
AamWg2bXRxK/Cf43f7SJIWtvwNsXPeVnHMvoDFcgN8Kfk8sKPIBJyDlVtp+IRVUePJUADPk4VcAj
fpBi62mZjxreqZHtglgPhgfoqakKm/kHQhjA+hZbwvDWzVeq4LsjX0B70T4O33qvDEPS6lwIVBTX
3IFEwQn31CwB4Wx0wCjk9F2kgTrQ2HCUaKEc+PoOTLhcgtdc7zKdCHjWYqP13yxteBI/lWzapgFH
dnDDiguIEky3NwnLBiknTK1oAkTJ0MRGCW5F2cTcQYcsim3YWu+rsWNIwkKTYXvSd25eK0dHrR52
DouLJIO6EgBvaXOojkXGXzIQqCHDPKZQddJhajkUQnsiSoNmwVtuMb5iMq7NvigWwBj3xigJLk7X
rlTSyr5kuGE5j+HNPOVO1BUd3mx3xJWPslVClA4d8rb3LpsBRP7QzU3kh6sSS0Nm1HLfgxCQaf0H
zhiJsdg3DZKScq0p/4rps5xJ7MfahHCh8qqfdPOP6PN4igF1jmnMk+A0ifHNue/1heMQNFR2l+wl
1a7Ja2cJrYMnlUgQRwonPz6YL58GGLqw1wZNh3gZarnCwPGB37HjZSn8QTPfUtoH+4DSp/FgFEQD
rHSUvwcU5CoUbX6Z6mZK7vLYFPONArsFXqYVywDZ2CwaY4XmyvktBBkTe/mrnI9vDeMAnSRjaRoU
Pl3sx2DIqkFJIfwg23Lan2XU2F/oZ2eXj2nP1QmnvYOUqoEJUogBO+86h5FiMdRyZo436I/hY+xV
9X7HAsXXI1FyyoY75WLXZPOM1bohscim6SCNgzX/PsXpAD2+8NvkX0Zlumrqiffixd+kbSeV6N3b
2T2/pHSgVmazInihdLEedE3OVozgRnfg2GYYGpgLoohTAljc+/g1fDbpVkCSlt16vDMpNSORRSwD
F+fQRHjEheKz2yoiA8ygVHl+zDjjvir+w4x9nDh7n3O9ecSMDL5HSR9TnVR+H0caf/7BldagWL1s
mDk02j8sPZa0jX/HHr53J8thgo2Zy+VrXcts7FR11fwpgay0J0bJchI27mtJejk2dfaiFFhVbAyr
N8bjT0wl8Oes++cob6NOz4RD+egUQ0TwAO5ZpTnj4dQcXMAAKCwronPBESX5ycCPXq1Ts+TI1nW9
ih0FhHNrBMSXL6v9dJ7ehM6sPnT0SgPeikDnSsFpjYWNinsoHJh+bAFwybWDPT63GuLbLn2L7Xw7
A/QQLytEth0rBapMK9r1A8SXO5/eqx2CEIypkilXk8/FgUu4NBjRw+NfbEaek54woxGgagChApEq
D/VmosQPs4zZt5Iv/5XlZ/LatBIS1jfZ3FHrIOYAJbwG4vEEyd1wIFrfkKhAzBaDpmV2GHzwBLwa
ioM5ZERpYoJF3W7m8k3AMW2y7f+5RjeE5raXcGEN1SyDlrgVZwbFrHQYgrqjaZnohaA80Xt7FGaq
bf7GH5wSllvj/1cmdYnNGDBRZbEcm78BtA9xOrv7QnixcLTYLpcOa2mQFxo6ecO3AvQv8ETUKCnQ
lUSg+BSlNRN+7Zo40O9P121g4/wqYM0GVQzckzm0mQBJHJ4DyHR3I6ZLiKzv2jXjmye04fVgZQ4i
6lPxSYOeOZkXObMiZJfSkhXz3CBYBAbrAej8WuLQHrrtLFP1eqMYy9fh3xUngnLZS+L+RXsSkhWr
SbjttVLfonsY4dwChIgjy0Ln1jW+qXsWe+KHqOL451vMg/eNRhP1W6JxrrDADBI//cJ/87BeJkti
CfKMjk7qK+l4Lm9ItSpGMRHOV8WJVdiiHE06HqHPJvwjRfW1At14T/pzFiOirMnE/+AunM5d2MEt
KBYNBfFn0QPAb7D6YJ0RCVxOvgzPmwACUQYGCVhq3nNRiEMlDBocQOI5R96tSqg7gboJ9UJzdvGv
VyGs9fGvKrz+T7mlycVjmoYfAoJISNToEBaHnfRLvIbg7erCHA/xTez520Vzdj4y5KGgaCN+c51t
p6aXiK9a/c3kl3Q+r5y/RAH0SS0MiqoAm7RV2RHiACp6ofQRRoI21pwmQ/g8sAQ4mh7EvKbWAlV0
gsrF75VexH/Se8xH/CQPYSOdOdz6bEzsq7kMTprw+L8SeaTUHKTQRuiv0JS2LIK0Yve6dzlCzrpo
A98Xo1De70H5tpMqzGMF3+blSy0JfpH0HHH1BJjYJjU+XmJqhoBap8dK7Y/F913jwu5ib/EwcGV1
WQPmSibOvzo1TfSdFhjODNz1fk9iE4nKd4SXh4s/iuCfh31vlmvhdVh99KGCkAp8jVyLJkMYqR1E
jr6BRcCZMginMqokFGQ3Ww+avLPRAXMHZzUGyqMurYygh8nl1hbFtyKm9Arq40ETWGB+1d/VVgJl
/Xbu7ICWlb1z07iWVklSFZGPYTvyrNmAXXIwsME11LZMpMCTTwdIJJkZ6c3W2Ml07z6r08nQ1lHs
1ID9usf8grtTkRIHoZqKhcU0ei7TeAUT6oH0PzKA6mVp2uG6kPe/hFwgb0jv8LXawyoet+AOXQQE
P8MNnvg9EDQUEo0Pl9vFs7PY1XC0UfgOKhtWv7LnOlsiTQ6Gner+pRpidyIMwJ3EtBTAmu571fJN
13m2YAj/sJeMdTJ6eKcKXXPq/TNDraIW8+BSnPEsBZ9N9trAcAYw9UetMLD+7wpommlkDTtMNUMh
RcQ79utu8xOVBeItW0ssh/vo7pkLFAxxoC10qI99d2UJUDse57IY1p/o5nWOysLfLDMDSmu0oPT8
OKQYHINHv8L41ekBgKkZo5tscEN35sxHh34DU+/bVNcKXvB2WacK2dVfVpkXuk/EbcK1Q+XXdvRD
tMgFHO315YlzF21a/1uxvWFE5N6Nh5UDZXgDIhOIVYtGGosP7ySxuLV9dQewDy5n3/e/6iQ/r03F
KcEI6GzGO5RGD3P23GgjgQKMs1uOt9CsSXpWwGFWNmUFWVRVPTvFHzLOhicMayFrcU4wYhVYQjLf
7S7nJmPtmhv1ffjWV9W9f9HTMQ32H6KVFzphquAy+Ng6rxoO+3PTtnYOXwUitlA9EH8xVShGjJe+
NcePMqyBSfENfTaEBk8zi7185xps/wYWg+bljzsxg584hwA+guWRVA6zzSl9YS0vjcuOxbggJhwn
F9hz6FbHaM4NcQdX9xH1JA4+VpVtIO2g0EqEvuzU5y307GKZFb9EgPY/Z2qrZUgIRUw9cUTwpcfF
29cdWwnsUYTa2gvgF55bRsBHlKgvRXpTb1AOKTOyQamqukRNnwHQN+wgwcNGKDCJrOtwRrxMFoub
GPrdByAC10QHGKvB+k+PvjKTK1W7z0RWQMeW9KH50Z0WyKaDCYsJT1GF14icx1XNqU8vA8eXS4tf
utq5GzOeFwd3hbpNjl1saOCYNrixQdaPXpnz4swHPaNXgrrj5YsUby2618NlIBfBCfnfj9G3nzIx
3yayAoTRgcojpLSxfNiP7PInF3F7oAuq5xCbdoRYrytzLH0eZw+flLaBwzzsGa73Dhcy/g2Yyv/0
ba+8+QqtVEKf5gh12OBwP/rWmh40DOplMI92xOw3ox26qd0n08BmrX2eptgEhmJnuTnzWQzKiCGP
ZSiWI5L4UH4nQdIHtNTkI7aREhl2tfG/38g5r63sBkn/SoM3e/Wx35OtGwNSPPmjXuM1joiEfwnQ
dbIdCXr3vjhyGuAu4DoKTjxQqziYtKNlwrXiS7GQEqVOW41SfrzjageQFRbQ1atVJB8RiSkJZqcX
4g/KPXpedHxk3o7jkJ5OGVA47PUoct/ytahjR4Nv9iVEAB37Pu47fOEUSAnczpF6E6IvGrVYA1oB
Fc7dLl1rlj/LGermlNElpynLgn/p+MFNgHwQNE1yAbZ5fnSQ87GrBydZTxEEBFRVOGWqxm3n6fpo
4KO9EP2NjVeJ11k1rzjguvYT4RqlZVLTQx7AWGyNnKvifhUahtM5yn9rXhaRK7Sg7LrZei0S31rT
VTtWjAtI5W95WRV36nFibuPx6tn4Ry9slH3faqUzqQeXIbZRW5w43Bc0yTQU/65ZnW/AIcwoEujI
SH5ehOIpFmwa73N69LNvemON/HflQ+mHUVcFrFZ3w+LrBPlfvnHa5oaCphTLjTSnBiwXM03mQVtR
yTMNqRnprRFcnM1PaqwbkSQHt1/AWtWKl05y8cjoVqFzaQgUJw45gm8VGBikmicDo8QpGY6hvJu6
Y0TTrAIcSay3rsAXIUTCL9chqVg3i0WgeJ3F0b7z0Uo0fN0qtZqL3yFie2BZPg47C72tw6uI8oFi
+tQyLx3OmWbgND7CaejN7YzVAkEfnWboSicjgfPLtzk5A31lfp6GXxaQUxyQ/QswJl4pGu9Q0L2m
R5/m+9oudPW+jd7IOM8uTkF9jdoULJtxMQ/XU26NMsm+BNj4llTS8+pfXRKuKSkaH3srS78H9aZG
mJ5r05JbRFWm23406YWREJSGAgXxbZpbFeT4d2cU5xzqnqyP1ZDXoO4ipzQUYnkYOu7YKhBZqqGP
Iz8852HvLqbVMlwj6Pq1Y03oG6IXpRj4lbxtgCaVmGfpRvYJDmZjAo9lWVHOPNKKMK04lDNbZABJ
2PiyM3ofePUfOW3EHu28RLxvMq29C0woLP4BpfUutXpMDN54XyptCUACHioFeVYqS8s+gLJ+lvwv
4jKU2MOVjY6jMvfOeoQuwWOrqKDyoAbv5PXUFyCx/wSuE8Eootd4Pm0gKJ+3LNYR/2d7YjjZ4SuQ
+0wOktGw7vMplD8beIUqmrFMQXRy+0eHEXy6u1BW1A8LoaPOdk8I7kOuX3u6UJ7l0SyRn6TmxnMh
dy/gxc+WX55p+Oag6yuxZIzx7r17+Hj6oyYKbu75PVrBdJNjjdU6nVtskwb/2KoNxSn15suG2Dpp
hWuqrvKUkxYUaDZ6zPxADNQd1p1mTAxb/wWaO3ztWmZtSxbqZSBjzGg5vwRnfgu4Aj/D2qWUqJB5
QKiJC87k944iZz9h+TbsLH+hVSYjZ+P7s18bzAw4RICYB8cBLL0jlJ21RQ3zOORmZNDagplWy6JI
+qx8tLr08C6Cw6kyv+ImAjpvutIvwJf7Mbu4Z4bOuVKRPJI7tmR0eemEAkwMJXDGv88+NiUJPZC4
ESkcaYOOcS2h/tYylv35C6fNfrhvEG/SVMjuOHMlVMm4aNxc03zT9OgPVsyhqYiYeVDwaxstpe7/
VhwY/3HSk4ZtJ/C+XBVruKrDgGPjcQOp/2Mn7QOPUp05qiM6qZE1XWOyKgF9ZzCnzWmiFwNdaS0S
N3r8BXce5IIJIi2XmnlpXWg2hCLN7MOBVH8zTjfBGqK6r3aLURnoFAT3GAPGeCiXAJSjMZ86f8nN
IfBlWPbTGqqYu8b9oO0Koti0b0OdoKByeDI530Yzt68OjGZ2TI3vn8xdxdcx8qj1U/XQm2ukFNbP
tQ4Hs/yFMyJ6GDMwfv9TMin+tG+A2GGm0MRUaaDkQnuZziApkgh9hVmiIg6DzjvuNFcDZx2Gkygb
Hr8PzhYvdmKIAVIQ7J3xAVfCrKf6gfzeAVelFcmYAu7DU1P4CjYfp4fRgN5TvfsJoeWO3p/5Usng
jfCFMEsuznbVTh2h0a9Z496gUofs7DdUMVq6lUFWo0zZxjOgqV4uWzv8ta64cvZrzjwPbpt8Q2o8
MhoDOSz3X88Z2kzGh5uol/AtWGrDYbe475Aia2m6hhaYiCDuqNxFcHcLACrRs5GAAwNa0KqMozpM
ymBZjngy7yMYdFl2K72A7SpFIqD+SrK52kRifrovvNC0EtYZUPUdRVbhZ68nkfDfkj9cJEmOFeKA
pL5iBj1dhbFHL070IcYPi0MmqON0eKpRBC7nfNOUR2an8f2kBf8xtjRJxhtOm/Hlv4VeBZaasNwz
jz63EXyCINkkLQoB6Do24Y51WqJY7IxxuhG2gbS81tEVZ8hLtmPN3HpXybLNle8YHpIBpaEQLCP+
B8V9grazc1OXHCsZ6B0u4p5XRuc1Lc32qeQjsdGZ6fOB50ouuOqjDDTUnc1p96reUFS9KcFP3gZV
HWJU5tVgRQaUJLI6pDvX0tpEzAYUzs99c1saLFAezr9MjQWBZkEP/oo/ZjGPy2nH+t5NKntlZJh8
+nXsIgOaAwD3K/FFiL5NU4Iz5WsdzSGbqnqnTjYWbfZ2nuo8K33jaMtpzfTljnNgMAPFyeCfSf/I
nTCTBvIpQI0Ttn6V2Ps2GO/ZyG3jAkbUzlm0QRHx9w0o36sdyHygo+yYfivTm/Wnl6IOd45+XKS9
XV521SR7jgqhqY5d2mRO9Tsmk1SxvGbPrmfunmE1+4fa8i9tLS2xsu1WZcNBIqviDi8waiNIJO6J
Zmn/0w8AN4gxxneqaRvw9f9rsjb3nd8Vvlt1kvjNnVkuulBxqKu+TPWtGPerhYXB08k+PP3oSVEJ
71OJChGICiX7oMUdauC7tm8Hsg1aiTUGBsWzNaF87SB95UyInZc0ZDhXlYleG/ylNAocqp6q5r2x
Ht5Y0UopYl7GzCUEPYK9YxpPMTNxbveA7plK/VH6gi2AK8J5uM+CNUqRMuzUnzDaeenLEbszcn2G
0A0L7BGjFXCOmrKS2CuwK5BaMsMGNmuxFnV65PRN/YTc0wE5wf2FJiEarOZOzHtlacjl+kTOboZk
yCFOHaP83fI10om7zDs2oSCCXm6n24Dk7vm7x/t0uhTm6pXgbWIccR5A9/59fRwazopVaH4cNt52
0vnRmLp39XTGwZBFRpe2j8HZdGxzrUDXS95i3SgKTtmDXzA0Irj2rHLBQTnuZTL8gi7lWvF53y3m
UzTQB97oM/Hc/XM1qgNavwLvopue6mQ3flcUgmvLt1/kL5HzjuOqc630vfY5fP7yY9qts6sz9zpk
Zvgd0IHLLsZkqdwQu2eL1Y8TnhpDywa0i2UFlrakUAQIqkFyb6PySAPa2tUGHraCA8drmkbuLQz6
1SBdiz/MAhwUIz+5InlTx8R3aEn6fYbKzvMMcC0H5/WtrkXjp+zsIaS2i27VNJLguTvklFpEqAPq
AWXMfulTRfwg8URVzjDId5LZnZO9zkSfx8du/uS5vgk1ZjdpX/hy8yZAFbDnmJsLdCovp39WAZZF
HgaLTF0jlxBwnkX6k1sV3GWNoZCEBzjhGF+27A7V7k/2jMjMMDST+YWZRrJsHNYp9aVufkxDoQ0g
e8bYknOUqYKZkLOzIeEsYJlnVH+sZ9/6rPTbfeA5gkIZLdSJ6wQnReUWpytzNC2doxXbiV8aZtNH
2wC6ex7BXQUAgq8qmNTF1Uvo1mrosRYmerR8Qy/Jv4gE0dkg9QFDHsAj8EbDfGL7Zmt7lm3IlmyU
BIvQJKfWGCME9Pcgfr1YARRje/3u1/mUvr+8pBbMC/1/hYgXznjZZ/1KNO0bw+FdAnb2j5TWGmFx
d4cGR4iVpM64oqUE6bLjXya2qMUgl8/hms0Isri80NIWzJiPfSiKCyLDBYi4yAjHNlkxgaV4+Udf
XlsUZ5tqFzJlzszNV0aNlP9WJXMDLaRtkK+g9lJGKEPPlvL3eYglo4DnKUYSkcB4uQOl+78zV+2R
f7hcWm+jZOs0PeAkEzKqIQQswrSf6yrK5jUaqyNcjMO+f7SppG+I6dtxAw+xlFdQgTh6zshPIhzf
3DsznfBkl4MATcmH0FrpdMs3b2rmaGbLvAAZGIYgsX4muuIM6nz+rBUnQVqHpVnvvPsxjoCEAHoF
xXpYMZXOfwFzpJ8b771s/4etXuSvNnA592fqzxK326s841/8t/jZQ7j8Iiv+iIUsQ+ADY0hGkHHG
QmtlL8T30R6OL4kZRPYUf2XwTy02KuOoahNn2jRDuUy9jaU+/vkRNsM8lpQOMdhOqsYRI6sF5Xuw
P4Yz+PgzsAo8iljM92+ucknEAElFEtlhzrbWUB73fBLfnkyq+9JkXDnFr1o/392UnhKw7VI76Gw4
Jm+V+cajx0FfPcopD6LJTHdhQQHMHsUc03bm+DNebiMW/wfrimgTaW63x9w6hnx/ntQCokaZzPeH
rWBUX8J1W9GD9tj3ICuHcshS7BT6nbx3VpT+CS4qYlNw7RBOyJ+PbMXq0qtoMq7crUxu4koodnp3
bU66RTM0skkg8i55sOAEgPN59CYtapnTVopoq3Jo92lwyGqSIDpg/7F7aDit+ZY+hKqS+ozWeyU+
4q8ZfhNyUIR+HGDrq7D5DSLsrro8TNtUkg/WACNikvyrRBKohUAfOBMocF5vllQierpxPFpJFy8/
7zN6LYaMlo27DRuFODVozWdbgxGhdjmzYE8eprpyhfEnShCTss2a7xuf/u9XF7q22tJECbo7zbRn
XhhAjF5vtMwjjskmK4fA7C/QPpIKqTfQ03i60CtxH2HjMBy2BYhkISTEOFCuE50k3CyZa48P4LXg
U0othsbXW8eVf9mdlOgxWFGm5LOcsny5+czAeoD0rR20hMQZWPmgMmsVA0DePad8Yin4u2u/f/QU
fLxzqvzvIFfCBpOaaopCj1nI0RvLTzIYy6kI7nP0aHRhvp8RzhQZs8OZrl3wV6BtGAg95j7b8nPn
+f0n9w5DF0XIrrmY3LR9JxwYfOSe4IoY1RlcAejPb6AF+uDM5uRIQ81ONIxc5VsrUIyvSB6tSX5t
5uX550w31foh6WfUlfLjLhdhXpv2/bO4T4/X/GXoEbDnPgUs+sBXZXH3rddXrYFUP2OUlKfHdWdj
ODWPTeV9sVtP7mjcBZs2Hrh3W+QZemmKaX6k+lI7n2PmQQu2IS4zwgyJGjoY1DlgSxbD0PxTiV9i
PFzKFtZvQMTKz3iF9Pbc4o8r5lrhjq/OKMDXXRLcirh7+KawdaoiJseNHXSnv0T+bYRZXk2dGn3r
EyNH0sTZn2tGrVJ3QZwklheDT/qyOI8SvU94LnIsm2mdFcpAU6voGyrqQJpqr/VjQhj3GujcdA+k
uyVa5nmTLiDfnVlFlSM0HiW0iJEE/ELhI6M956q6bfzIgZ9jgMV8eRuec93kGIbidm/Z8fHosIZS
T9P2ck2CxsPFO5H20Zihelwu7AJmhEBw68EKk60UzRndCotOQtQ+e5DNKSelRmTH0sG5HGmB4kr2
dp04TBC/aIr6qO/E3qvOPqYGgFfsx7ke6g8UOgAIk5wLO+mjZ1GEyn1z7YOBTgKaF0EpjrXvaRkc
A2ulc3ZBjX79W6Y58+GPf7A5bDpn3cLJs/AIbGt+9I7jzGhUYe5Dvd4Z26DXoJWlCUSVXtiiujjE
Z2+zp9ZlWxAtI6gHkJJB+uUoHd6L+PGJa2UfeqZTCvI5nbPLF4Tsn3DoP35frzrLt/yOpqBefS2W
pQLupDkc0mGIMU6aihYNTXImjKzL21QaoVogVyFErf95OQMOiwSXFQJBi87pUh/9Bo3WY3wySu+T
4tpI8yHH3lXCvXfnv7+a/7px66X7EnHAe3KX/QzrZGtfY9/MxHwdmvrFkj5A4Oym5/U74mMLe6HQ
vQ1jWnx5B+a9sYZm69UKwXM3hcSNQQg/UmOw6VgUO77RdtZjFnp+6JFmDfaqL4uDpt2uY07NR+N9
ExnziQGriOn0QYuYFYUvyZYKgIwCRVRU4Sdehy4w4ox/HDyflRm5LPQTXo3yjOvOLUZqAFesRA3A
azKqDHw4q4JXFDhMjVL+xe3Khwfj9D8a9BYQwnVkCQFpYxNmt0dYRLqn1jicWvCI1xUKYMv6xtee
MgXoFbUJk9W3Pq8cwJKE2x90LKWOcZfMmmhja1TIuSagQq7XB5I6IXNyPE3PZbqPaor1UahCCSFt
NRO6fiYMGwLKGWHHs5jEMsNWvpgWyiO11NrtAfwoymxFe5Xs4xT03Vs/ykpuxzJTAh9wnfJuMff8
1hV+ZfztRWjsH3FFN66GKdbuxuw38z3uyuMe68wk0MfAvEKHs89vY/QfESCE4r1lhTEiqJOmna5H
xILvysNHSlypt3MbMwSBxsyeooj8Z4cxHrMWfPe35s+i99n1fcXuVO9Db7DOmGu0oIrez71yzS+E
AI7DYPM1zB12DGHtYwloW/WB4Kw0Tn3k8lMJR0nM9ocaU+LXhLCgNfOVHdLapoxvlNv/B7hCKZNZ
I38Bbc6eKoqn1akiuAn01GMNKnpqXBMA5Nw26BBJYl8i2/zhzPNwOkN01McFjb0cz+r3GJaA/9hs
bN6N51AEn7NCFQi6O6e7NjmkrSmNVFj3G3y+OBIbpBYJJCL/3u40g7EMXqOcatlXhwExilG/kgdH
6bZLS7uiQbnfdNm0QculSbGD1/AFu+d5NQmoE+2GlOBwPJHq3nSrZuxd8IPSqDgcWNwrmSZ1cRQV
FFYnwKk3adxrkVm8lEhEpy/3K4BaPzL1JjxDHmuH6InEiw8tKWKnjtB02NNiZKkYOFrAOlwCktqj
rbtemm0eHIQG3X47e2+pUjxyfLdkkcfMNL0OcrjPtyGkqM48CKvKAGuI5VtsaYiRFcT7bfDGsPRb
Afh8ik5J0jAZ8NHU2dC8ezzNB4rGN8Sz6ky9R1HH5Fl8lbvIwxDCyOhiyBfspEFzIDeGpgd+fpXu
t+IIea513lBrTRLIBU58lyOwx1kQEOtk0y+nb6sffBi6MD0YJRFmsmlVpy8ydyoGuyH5fihiuezw
Lc08kAqEgrskiWVdYGU4HwoiQPCqhxNRWyolNfB3RgAnYLIl8LSXfm95Ez8/uDAAqnPQ3IB12t8B
G7U5r0tX8jbRZAxhiSYvDRcg0L6hfnCUeHFsVMEMEmTbZi8MZII1gTrsjHpQok5QyuyZXy3jqpFD
/qLh42O7FT4GZIeh0SUYGV1QJvI7TxmCqm3z804LULinKEKDqFcI5sorwjtc7kqNU+ZgGbmYqwRa
7zQLfUL4g9KW0mpt9ZjtiICHNe27xSQoTeU0EuqKV6vtN/OgfKd5MqqMSXjAAUuQ/+9Zqy3ZSuQ2
vjkxmf5x8gS5A+kuDhCGxK9Sit22EQEtkmfL1YLiMFnqRAAcrZPOPAxjaILLJmL8SLFC2axWsl67
fqPeowcwpBHSVjNpwR/yxCDWzwn5GPOhB7TdyVDkf5ulfFvTh8YtYOgX0aOwolz7KRWbTZNM19dr
u/mttgVS9lDLYHfu9Dd0ITn2Q3/BejOZpttdlPUmn+DUo5/wMtVRYK0b/yUe+RNX+OOZnqLHm7Y3
aL6Cc07FErLIfFeTxjchlBg4Hc+3Y5NvfUlr2PAgr7pjJNj1zUEC2W26xhaKnkvI0Vtbja7HXVax
Wc06ec8g23AhikxOg2sSd3FXlM0p6c09NlCGi9JUwSSvzcWhTvAuDCKBaCysX29ZLzGZpRoC2LZB
7hy01uCqDKiBk3/EXkrb6u0GhLrVzbFLqr8EMnZ+gNsinCqN7n9ME+nVeHgi9p2+WsO7k2udsuY7
qidzcT8v53K0ZzJkBnFqLWdv/sln4o8O6zsh9O5AfobgCpB80IaVewO6s7FfECxjy5x99sGZvDNh
sogTmhzIH0ZWqHz13SuXHrZYOYN9RwLL6b0Ov7VEhV/xXEhEfjPvUoXYP+gVyyQJkaw630wIeGwT
cvFKuMpr+SmcN/b61E8OEGqU4uBPLUocZ3tmGd05nGVjbThij/k4K0F/Qe4aCle8icwdoCe/Kh9j
Hw2FGLjTHIIbuHJ3jBgPvgugk9CiLNzt9uMwoHl0UMmjwKSCMcuUGd0cEC0n/1j71puGvauMvN0X
KQmk5ndFyp/y1/cE3l3zvsMHP7W2/gCQS5mXhgCMa+Rq77216I5cK8vvsY27oZf7
`protect end_protected

