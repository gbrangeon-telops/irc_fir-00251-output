

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
JoMCOWeb5WJCBfHoFXpAeueDDgvCDiGp3AckCc481MQYfkwqbKzf91lDJ35VGRkR+lnFDdba8hVh
ebdPAvk8sQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
bZP6jV/nU5x88OLSeX17wUzGVM/1H7fFl1OvjJVlfPM0WRyEzOpDDBDAUuNgnxFvzLOKKYEuQdGX
W9Azus4jUwU+zlgsaiCb1S5W3YMjUJKtbRQ/PvNNulBlTlfZaMHLAox9gfCqP4OK4hzymuRCwSK9
PA7SK6I+FbKAacX9y/g=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
38Ya3DupjVbpSJ4i6CmxC3OEuL9qNwdAvGt4GnhSmvDhP9C+krqPc261IqfCwYzwzxzaeMibTDWx
/h5fHzYF2I5fsXilkoEoRxiVUecJo1YSbQfTJW8OEBtN5aYD4EfWNZxg7GXemsfNXYAT3IQ9OGaZ
Z3OnlMzYiNTbG4DNtpaaHWOF6C1ZcpZaMxg6JA0ZIcSPls5SVALLcDt5FUbDAqBNYpV4JoWo+qsc
FnhESB/fKp4TYpfMu8ZebNdGwLZE/v7NBBWsur4E5vgpE96o2V2PrhB/yUkeOaYd/sqFfOVAPPYH
mOxmomWznEckwZ7yWdfaca/+EES9Dh2xe5bnww==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
D5raxCdsBjNBeucgp+JNk0QydQuZbfT0hk9FPoXi6WfKMKGXanrHw+M0M2EvNOZMUencxzfv6CtL
nCmVqYCrBCTP3KURzHM5DqNYzQyp0kj6XGMA+Q1QHtCCtnTEsuFMkRdychCBXeOcnfn0sPqhPAb+
dDkLPxvSvOkSf8WjYwI=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
KE84+0MQOal9OYCn+WiAXywM19zQ4xYNV40iodnIlowR+vSp+kbADs/ClNTsY+01AbPMnO8ZTgZN
CGRjsRjKcpFcdHcCbRqcEDPJE7OK/v9PEqPDH9NFgGw1pSJUkP9IpUNC9/uKTepjTRYkaMQQIcwb
MA905J1RyQ1JTo8+T7ZjypavwIpWqfh9+/OtTNQBqe8xPN3IUu4u+7M4P7P5w0QOtT0XGFUOVu4C
5WyMVCFrGwdZoGJ0XcMR+keGC+lH3zgKGf7XDuZwC5nPj50Jr/CWT4G590JXwyjmGrh+LuEInmJ7
dRdHoyo/UrKvxi9s4oal4X1UmgumWAW7Jj7wfA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5824)
`protect data_block
DurdGfUTPG0uRIV7n3qylldi7xYuYAm+kDGTN7QJHJ4Rk5HjQ+bCJQO+jjpHsL8yqPo1E7zFTi4V
hkCSCOS14VImzp+6wEXHYnNAhhRSBlDMaX7yMh4LtlAsK3VxbRlCNsJefxRlS5b30pfoJJ004F4N
9dFs4mX4o9veEb2SxUj7E2U2Ll4PmLNX6ThowgC+0tfgPzcKuiHbZmtNmUuLPwEwKbOXi2BEOMND
s0hJ8u93DwXtTackpHVDL75SAtyl4gHHYTU/LsbDzxBlVNcy/6nRp6SMKUJ7M5hf7jgIdmyzKRiy
OH7ug2i5lrCouK7eq9KjIBe03WQpGSAYHHMXibIyLGcM2sXBx6Iznn3OlQir93j5qhcSwcXlzSnN
msii29Uj1JlDjqA3/Q6A6f6HnJT+AU/D2F6nOseDqi4EaC1kgDHqgUcalVUVTKkgk0GZE1wvFCM6
HcUXxZ2UVXqXhzMo/2MuTqQarAyX7hPQpUbKquDUMBUUOovje/1fx0nuzPpr+oAAsrtf+6gZCK9M
C2SafFdL3Bdr6pvuaYXIUf7Pg7jFPFqIdCZIQkouOjl8QujFqsahEqVxIHpTC3Odx1BCgNqHp0mW
dtK1+zXKY4pkUl+31KyHxs3FLg5MuAdTzuMU0XkGKtWzPb9qdp8LWB9khrN+/+Xbo9i2qJ7JLAhN
x0eUiC7g1fKS49ETlOExtHlYQD9oy/xXRtQMiyczbc4xk9FyFCHJU6AB+OPOFbALu7H4nBdbj7Ta
qfAAAndkLFcHuJlP2VauEK7C1XuyEKfppu3oXP6u/yqFlnr9MIiLDkyLqPBR4SROCHsukT0FkxeK
Rs7f9bC2RRAyX/5Bidx7qb7Tvj6rasB0Nhl18lx7t9j3wIQSl3uuPUIg2WR8iTxD4+YivtUfjnvG
PiEGJJXxN7uYD85xUpPn5rTUaRDMv6ohCG/7RSwtbkrX/tMvNXNGCrDFpqZePnGo3YpaoFhOOGuH
M59BTeu4l0uQoZ6ILHAoVqIsppyjt1SyAuPft+YvEaGWnTbqhcD/J7uac7z1TZRrmqat+KKlFKOi
QrYoa0W53itZj/rAdq1TkH8JIBVLwwOZUmu74ztuAjKWAtDSJ5e3HPGBSE+reK1GnIWxF1yBlF/n
HS9qgULI10RZvvKIA/G0ji4v817iHyUXqPWs2PBbHpmhEgSDHfL3lr6YXNX3oq9WCKp7/5DP1Oy0
P6PFf4s22v/88OxErz8qyG+Bj5nC9f0O1Q6gL4jNC1VUtesPu/h54vZdRnq1TB2jfNZC52RQh9PT
vxmPc4wO1aGX9QJhd5Jlt5/Dr4e805ny5955xtTCppFGwA/GnRREEfy4DmcsJ6q7OxQQAbuUjk1U
1MI2/30d03qqsibqxWHZlFnFfx8qLpXtrASJgQRZTXWlWyphLM2IvIVINNQo/688bR5Sh83T5RlS
QP1AdEGwmmKFn3zsPZgriaT618zdyWxkRh1F5jcGmaUaMaUvRBUq7ENWzbZWlwMct0DpPQr2aPIf
HfNUM83u/709sNCyRfWbfB++DPlsEo/O9KuUox71BHpZEBB6cN2lI6S+O0LDmsOC/bbohCWHFu4f
Nz63C+CHLMEuff6j8A809UWNtOZ5MCkPcWWRtZtQ2eeyjOFsXIxGQ8/9yDY4EfMstJDSs2+fvgkD
pFwp+AAKRV2A9ZMbqkK34aR9IONitdW9NY0sKmYL6s2iV6fc0bItNtMqVh4ASNA928zkfRPr3FtO
Vft3zjJn6IKGXoHElY+esyPuwKO0sVGH85t3DF2urJQqeKLn8DGX4znQRq7r7uCONIpgss/PvOla
ItEdRR6CNQW5PLOkDUIkVkKpqn6YLym5bd0+UqKECAIQzE6vATfX3z/Op7lvQkRiHRA4mR79q6Q0
4UmQmu2as/+b0rzmSRfz7l5kNlZbPb2Ae1GWywrp7vegNn+HbrZQBrpa6KhQ2r/rYpLXyOC7pwev
4CGc0NAZ05BzZCGHvyyaAQ2ApNLq8vLT2ctiVlk9PsLmP34kGZvk+Dgi6mcUwDFtQg1F1sEN0xzJ
56TdDWgvm06K0ofatIyoIPJkcwCk5t0itbr6Lvv3/s4BOjYFjTFkAAK2ZEFCJPf+uKtcVTG7RiLA
DbHxhwKmPwxWYy57OmTOFnVtjDElQkpwZTg577RB4p526kcHCXq5dEUV7w4WawB2D4w+itLlXXBO
grpGsaY0OtwY3+G98M/UY+qwKJ3Vwijm3pTtGAMUGgH1YVwuggOSaqa47ooQ0yNvkQ0FuH+HeG10
YfJRmG/KZYy7DAna8S9xSnQi9aJ0ZT55RECFuR+qO1TEb5AKO3aWqGJiwp276uSa6WCCCnk5YXYo
wm6WmkRSJebXUbRE/C/7GMNHZ3iv84Cj552uCBY2PZAS5phQvgUk7BGO0jkBFPkNc3opQEn1eKCh
2jUuQQNPuoLEnkeczWHyJw/YYwKVbTzsvg1Y3bw6Ypi7Fw9e+LaFOzkr1VgACz6uS9Oj90cUJooL
tr6gYtbilevC4ZerfyzP4ef/n+rPR3g3CQPs3FdMthqFc7T9geU2ytv8Q3FQvg0J5yFJcIOey7nS
IOOQVN66yl2oZsV3CKW3xSXR0cassrqFXJxKLn7bzzcvx5eVIBFqlVtU4OgNp1djAEBtUv13CKwA
ZOBJKr9zIWY265Ig0Dc083yBW1439ctPDoqXaKvNVQAcz6KVQGB4byqG06dBdA8zJWkS3ih0SiAY
+VQNCQhwrVRwGIxYpwN+cW7IFL/UQmqkVnctd4Y0OG9I6gHwEAIeup+OFB6aEI8h8c1iZkqWeG9S
M1LvBwPVE5r83eoCP+GpuCpvCWm8FGYrQGKr1PQkoPuh+NGcAQZmke+8uAwRTSUByzGsooloTcS3
4Jef3RtVrOXJFVglF4nNbbJ4QV22GXse8k3uawbwaoWJt+5bscuyYWxjwK/vLqV5pes2ZlVYymsI
0DEFyse6uU0nyez+yBUg6NbwtIopU2s6Kz2+aO3Mynh86BQ7VIagqVAeqa3uTE9A31GkHXs1cvCr
MUg0ACXSG68f1WDmVGvrm6CZ7wpCR1Wo3GDdlGK5JBQpQDawHvQe218tvSuQ5H2S6viJFOsLcfLq
tgWLDx9T1TFVXwZbmCKzUrooHM5VrN6n0fHcRQ/rYECmBIYmortvEfwIIcEseZ5tD7xPMR7vcMTQ
Pzl8l9oBqV1p3sS9h/wPdpurWz1PPgthTtAT8hlEmwaeWSM3Kr17Rz3jKx8STUcaSdudyTuQWeRd
/aNLVgaiKfn0JD5+viiF71OuZL2oLkoQN+wmiIHBorETemQn3AtGEGPakN3yzwDk99ZhtJOlXzJ/
WLapwbki2h+UYD7X15zNN+t4Hi2/fhBcbOVxG1duJRoLclo3uXi3omD+Kz0WL9K9g49+9jKxpBGS
u6Obc7Z5ZD7uXUtyfUYEJ7KxaIU+5Fj+w7LQhgnx7s8IstlorKERz1Gi80TEwaZbPRkkc1BkFPMN
QS032YvTkTC3v8WN0r/Q6JXxWOBsB0pR8hihJzsO2sUlI1PIK1074HHLbQ+Q5P49PwaNWoceh/XK
X4HQHF3oi/+0PhwLJA9Qo5ll+vhjJidh2b2SuI9LyVnxHix3u6lCfA1thaqy0+RhnFhKzLCct7fB
CjvyBN8DwmRFhiQ7LY56MQZ+xCydGSsNjIzonm9hKLbP2umktNhuYaGI8aLdoj9s0wJ21QpjH0Ph
ptWgeawRisxMbUVK1ZBZuDTaB75vrg3+B3QUYn856ExzzHPcExUlgj/cX0EOi8dlSqCpYaTyvlN8
L6PhSU233cEkdT+mLjmOVem0d4mL8/k5uiWLkJ1YJxZwUtOa5vbLxAL1xZS7nHq1Btt4Pe8N0ZpB
y6459znGGPdKDj2LgOXu2OOFvMpDHx9dr6pWnXaWNufpvtyev6acAhmGrnrItd+ypf/YVSJjShtS
lLeR2emahloUSojyPoFUvpaR45pCfYNhfQrYA495TuUkiDP5J/wKk09DUcUdX91BehVe8Z3N6OCz
T+OVID7C3abRq///BSUKlHAc8BKlLu0vNKMGYGy7NtR+3ojTlsSfN8e0yvKGfONFmQPpxOYdMF/D
5UpNXo0Ovka7v/gTex/aMotduUSCbgYwhCsMjFKnkNEoD2p5TVswV81xHc3oCZ2XkXV4Poc7EFeF
oAc7tN9TV8LuSNNWaU1BcyIUSyJg96teWWMOxvTznbFuUy9I42rXdeVvuaWYJGeIehNKtA+WVyeE
ODcPUDRqtzW/iReqGlRnKV4Hm3qrUrwJoxFrXgPzObAlfTcAW0Wc8O9Ic0K1xUJ8w4y/5wNmKksp
kMaxOd/HYgzqwaX4JhlcNz8M3V6Xwxy8zXdDb5ofEXo0peD7DB0ZaWQBUIUDYXo3X5dx5xCiffva
bq8hZyXKx1Ro5g2BY9b6jzXXt8x1YUJe6OvRLH+GDmuUc8YV/VZgp0rg1fXODbGP3sMBhJVbTsE4
fFjoNoyRlb8Kl92tMwadUCUi/pLUieG97pmx4WD8dPxAWG4fJ5yqw+vVV1cJaK2vFbfAwx31PCQO
K0bmuWEfom0m+rktTz4sObHrQqAQsPuulwbC3m40PE/pGPWjBIXFtKa2taiwhhO1ZdAR+7+nFrzF
qfQJ5Zz2leca+QMsn08GxBY1cVDx05gHYRv65H5/9qVFGaG0MZrUB/kdx1f7iYxnYg4d+iZIIj0q
TyHM2fmIPeF8JrH2crDmKaiLgSpzepDuyVQQIqux1XoD2dvutX+h0AVmysh6YVEiTA1VXw/NZpH/
gTIudqKOYbvPBpU16lO7MF1fNWZtRIRW6lOF7jXcXPhNXMaOzb1c53crNYqC6EVSPf/R2KWod6U+
RQejOW6HL3RKCH0iRPDsUzf2fXsI62++XD/zkw6Tp1pOa5Wm7Vf0YBE+KLo0gyv9GgFhylA9nCBy
pBX0NBamTOS5mVOtgUDLAX0j9JNc7c520z4NMm9NYwSit+/hh36xZ8VHG/hXz2m5y8FOani2HOcw
kVz8Qppe9VB6vwdYbNYae2X/1P8ucuh2hHcmyoyAPP+UjpVxLwsQBqtoGghnIMACLlAjEVzx0szj
7nCX3QGujThPbxFeUss0heeiGh9fpfGI10m9WM2KLXy7EN+5S/MD7DbiRcIUKNEUFvCXMVNyt69X
4Ms/ineHwX76S91IPfXVPAgvCqv6gX2RTpaL0VvZvI3lNIrknkLeXNfXK/jJhphu3DJ+E/bjqS4M
ERR3LP3tiPuBCGyCenPltfEWaS/QBYGFHJExwLASHkSL/22W6f0EjsDNxisXj15ymy5EwaLtn/ZH
1phAYC9SErHo9LdRcf4m0CKEX3dtSDcra1iqiW9NlPVv9uW5gSdjKChj+xMquhDlD7zQBz5nzB6u
et19JBGnT9mS5eMcnXZp1kxkBB9QalMFwy9Rb0nfFdJs/0tfyclHc7OyFb9URADWfM9Brw8b5b+/
NSuqqkdQihzY01Jyj2phDrHbnSDJo2+tzXBz3mVQZ3jW6hXbmgQQ6nLzp9yzzxitEAYkW9cG7o72
01v25H33a/9DZ1c7DV/ucPv+ofePT5DFJ+SNGc1AhxXCNyEvg2f1K0l8QOiLk6r24Rnig3qB1QW+
ZVw580t+g5CARgxjfzh5kLpjhqaFBaZXFG6ZQFySMcOE4S5s3/5LUvNiuM3fjnbPB7k44qYdVoq2
B9aU+p9TvpLSB/FoL+8Ny2uA2wdbLx1O5dHFKvqRXsf7fs8ERnevN9U153KKOBsL3elPVOiXWXmw
ULSAOzLs1ENtAmleJpl8qw3I6VDJKd/L2gL7LOmxtksqEOghOaf+H5rzHI3TVLaqmqnQdEyswvim
p8qoGky9s09Q96zsxiyPMRGkeVKxrAfMXlXJKCDfjJEwo/L6dbUZQ4Zp5EIRtv5Gku8Oi949prFR
57jo/yHwHGy6M54zzlBhljSQMrtkohcp7rOQcuIRxdxKXWi1AqktNPAj5UAy6cj2dqTOhrD8lj2U
o6ETs1HKIC2gfGwhW2WpKY9H/pKRfwVIAgt6BRUScPdzSbogf5j3eskXHUxF28I/nP/CIUtdpzXC
K445GOlrHRKJHlN2ohZy5h9IXoNiqTOZg7gSuSideAmzd23tosvAkWXfgZX8aQv1bImGSFGu9zyz
m7cK1HH+zgJ8lAxB8dfUbLrEccFnQjuxf5xD5LODVUiZLBvVDqzYJKHdKgIHGBweQHwOn/UIvp8Z
RFOdPSkQBhSe4uh+QR2il95+jn8JElMTpLYa3RK4loL/w2t9DLgSazGLJGLrvYL6ttl9TJTG021U
QNmWsN+ShXtDvK6qan+alBxsx08TdGccZvIho8Kud5GIv8pyxXjQLhQ5+MOYlDSeDonrkU6i5+2J
z0rCf/Du4cTxqBaEUYyfuOiOLRJSAJ6s9LaW0LZoOU0O3IEif0qep4JNrUoYSChZTvW0PpmOcquH
zhHt84M4AK6op+NXw2Qg6QU6uqZfeBynd8I/DWhljUBpwvwyhkA3NyoCNleXODNtAMhJ6f9Ppf2J
i+27QAfMe2F3RTyG5V1Cx9zsw9smOJrXuxrthN/Pc55z6Jlu3oAPOPy40JzrfJtuQfKg6qKru7zw
0rGpTKFWcDgKAltgsBlPVtwiC7+KfPZrGTYUrMKMnmbcDUOfBGEUB9kW0kphU76Atr5AHJ8Nevn6
4WPaySIDdmGIE6jRruWKZHa7m85qtWDew+1VR89VpjDXhubzgVjDTQbV6hklQ5iEV6tYAklGJbg1
SiaN0ASRdWhwD48YapNwG7PIz/YJ3Y32yPuS+AEGUsOmGt9lqAZ749J7T2XOwSP7/Q4i/ODc7r6v
3vOHyW7m4OiNO7YFYVUAfQireRrqib3Hiomp64GFXK21P2zqPBmc56/ZzrcweshP/w9mBZRoKci/
4Uk89NsWqsaGBH1Jq0nw3/UetAWfy5kxNsrG6Xo7T5ATmcu8x1dqYiDRo0zgoYXLOCiZpjLyWXFL
YUc8eg6GNMLUpuGUTT6p57QJvgolrcW6R8YcacQW3BgBTEr2GGfVKPXZ8jVwIirzJJUZUU/lo9i8
/71+q3OreN3iA9MOp8jX7VDMLE8pBjljC25OvJdDxcZS+HUbSknFO//ajXjoFWKNM0cKsDlIxawl
dWheBFTwSIiLsF/5Yb4w1Dy6Lg9zMS0PIlmZmacmLk20uAkSBCQmZeenNjIyZ19IKMrVFXJBjOqj
8wmBqz1+q97YebvcVhFMtJdToa2ntzqE439UT0b/7YKSBtSpuFJ04u+rADI+pQY00ZT1hktQ5LTY
PhH+aPqSh3XjhG6MPZY3gj5WPTpODOn2FUojlL5UDY0cbzU5NSseDvI0OnAq85dgiottpMLKfO2s
f1TyTqkz4Rv354q5e3YVPQDdr4WykYw/uS0cHcGtKSlAfwjRItULmf6VsPztP4eYIywsYmK0VAki
cTlJk6CLgcR1Vmz2ExWKw3a76JRxL57DdXMsa3Sjk28APmTuLSzpdJTfBO7klp6j8pKCFTydzsFc
sg2oH8oUXD3Nsi9a0iNYxPMy62z3Kw0QqpPwXlafv8A6yc5IMxHfDz0n2IK55fW1yg778dreq2/i
vFf2DlgwaU32bYbx4ZRhdVbqXXEICyy3h1Xb2HBTXtLNFSDgHcK3abhOJddRyLxxwRFX6906Evlm
WYSDYoI7fg+G7P04ZBF729OUIBcoNLsCNgqvNTIFKMz33tnByL0TrSOQcq1Su7eGtwEjbAp/Qv//
erHq54R4RHn3pw==
`protect end_protected

