

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
nqqBtmqfflVo0LfdOWD2OeylbTCJPLX6XaSqFQpCXkHX4TF1QAXZspyiDVaQlwRkat06cPZ5E411
bTzbr9/qZQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Q/X3qbnpTyRXgHhmurX8chlDRL2XjwnbHjo5m2aoqrTNSVAUPYEYGIGJVoJhRP1Bd27KZbGI0BFX
fZKfju5H4nz84jXPUC/rcsp76WTu945qoXwdo30XI0Qhi1w21P6EhLXccz1l4c9zfTwlHtVuYV2c
xkxHRh0F8KrrR61HDHc=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
jBFh6UBl2pQmyl/KNdwY4r9ld/Frb+RgwTVitzK9Y6Fp+6xDwrsib4d9Z9Trd2PuW5z5/ot40n86
vR7VZpJnONM8UmDjWgdiB8rXNXaI1rBfme4TQ3jj6RaF803c2cAi4cdZ4qM3X7V29W2B5HXbYsfA
+fn+v+caVjEUXZHZm4HMyIR7TNVnvmCWeeLj52d+u3MrD7UjjkqtqnRWdy0ckM9p4TE27eiu/nsz
awiAJoiVLZNTMmdaTdZ6vB/sS67SAe0JjX1nTwssfK86UYU1+n0NLZ+SLB4lkqxmhepGPNojfE8p
9hJaPKOTV3d/umJbTV97L90iPloNPMXpGK/m+A==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
cwUUX8orCEMoCaO4wbzIkA5h1G/QOLlup3/J46IxMYEEhFnVuE82RZ46tcCa958uxg+L9/l1SnQ1
1Qa6GFDzaEz3zEcSDS+t0jFMPNI7VUppaIgcalGdkOXBIX9fihrhASeWjqmTDrUSlTt7Vzyo+3TY
n3HFHRbTrCchXcVswqs=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Z1XHzIMnint6AvJuhSJyN/+kraiZwIT5ZFNyZxcRS4ee586ZcCrsBlqjvo3awgeNWb2yZNQKbtJY
UBJT2Ww9PtMdwpg4MPuZFMCTECdiBOLjqX7gX0K3iBdA+35RXRVkpnaon7ABi2dY8SU6a03iv3ph
ed9P79UVGmdGucbzSQNo8vkiW9pS6ZJElXKmEibSc0C9Vw6VmCNdLosnrss+vUEVkPDu65r8MqDO
9/2zcjIio0kfnpSLOaIDXqGefGNR89nRv/NxKymzLnDjvK13FSfKq6qNfA+cXOtnv8oRuf0tdkh7
e8F12j/LQajA5bXDfmPQ3bNX4Qv06vuQ9+MAAw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 89616)
`protect data_block
eq7yLJUDXAi5J/iIQnEnsCyLnhPB2mbibXgb4Bh7W/3cbv3W5ccZCFsZUJR+cyP/aqMthFrIRtFt
YijNjvaUayhMeqZjJsxKUapoXh+oxWaCAIsCIkmEa6O8omPsLMe5YRsmjtZA8mkQV1bPNbtxHFvg
tGfuQAwFdm+lkTcmDYyGtSkVPqBP9TGsmXCqH8O4x9XEnOPJpzNML/PNpKpz1xldXVEzIPt2SFv/
OYpI5Lz0W7DEpk5rr+zPTZKoqY9y+uzXooMyW1Wrb8ymK682XR9jwLf3OletLgL9CL5M2mf+vpU0
HpjAkFiR8+VyBkYmTMe8yznf8jFccE7REQVG7GhqZ9SNk+nKDmUhYECUt6pyXqSsNpYvJDT4Dpef
mdqxYgKhRSy347+I3Akw/SiYZ+Jxq8rAudQsvq2Dnm7+HlZyfmTj6rsEYb+oIuy/2ZiUTrNmwHz4
NyKmNTPmKmc0mfUDHyYkfgsOnOaBdNV8Af8cAgm0rSKws2wHg4Ok9ZSh/qzg+Tle0MZiWvAl5jxv
fBACdHN8EB20jfGzqzAWQjqRD5iCcmE7vFnu5ybd5Ir7q0uLSKdoNu16LTKWsxKmIvzYT7GyruMi
csNAIgac+RLCm2plomRBYbDk2SdJOZQ/qaXURsmew0g2uOZ8UA10ryKq/glfldPK/WTdmiCr5cRG
YSVgC53GuoFzkA67YxRZtW0znCeIkMcnt8LX94NhoIoeeCwfKxGA6ygqZqbPphhZapkzs7ApISug
X/wTVXduv1pXTslA2iEpiB+VbT31haRDrODndbyFU2N31tE+an52HNnpR7dnBTyXC+gfMytVLFBC
AS6mOC0efg0C7+5jgPuxSOFEAvAozDVLh1S8ug5rkT5+P/P99vHF8addXRXRooxTdwWm6pG3PSrT
FjGpCDW0YrSWWic4sBiQyHpa6T28l5/wp3oRYpgsXiQhvMkFbVpIKR6VwyQJWQahgeSLvSU7nJb/
7NifMXeNMvoMD1lnkZHRdaHAv95vkMu5FbKPTC/SP860G29Q0wIpREZ7VHtNTPJkvIGAG72QVnOF
jB1HkYmIFhXncM61HJafOKG6UeAGVOHeaaRmUqkrhTL8MDn0c5BBmQ8cRdKdFJWEHM5AYP2Lqs6H
aVK3Rs1MDdztZ5ORpUG9Y0EE6RCL+hbGkVNa6J8HB948wd4EOKsJEPDNwlv0l4pRqwipx6MPsoyP
0noeDn7bv0QVRrMQEmwUVoWuBOt4+Lt28/9YMYbj3qZGHzf9UH5rxJd56/C8EtT7yhI4dT59Shdj
Eh7dovBNSB67cMgWRXX+B/cS/zQaOOzA0bAD9dLhy94dCQ8J+i+0AsUCm14mCrFXBKP/4E+SDlVX
mhCBz2Idwud03sZxzaVVYQzsVThe27RRjeqmNaQr/kwYgEi6D3bH9AlwH82VFKrRNgjjS1dmxpVv
mcxSDLgKrRD8s/pV4FbuZplu5p55cZed3JpqtHOqMeZW903rEiYOHAaKmLngDtZ4YNaJs6OXhCed
rJIFAp26Ag0XXkNdQFTb3LmJtZI2/IJw91cO9p3UbAOHjRk8I/GA5SJreKzVmGz1G22te8gtLDPS
pY2e+0vbdHkLikQ9YwnDJIYXjBpBUXeJlGgyUqokYeve40phSYO82CSQVdZQZAcbZcNkNpg5o1qk
P4kaytASNqrNBEvRyoXkuS1A9xqumfMXvzPGQP8pujYFZpRxt0r3mMZ35fZc8VD52l4d/RDYtq95
gMHC69qt0y6Bm0he9f2GHN71c2HXCJUJi5alMrltc2l/W3rEQqYBwInpQ7LkrCh+kgzF0/KVk216
Gd/+q5Kwlbcj/KoCEyedGgsHPspdrUbMzFs9lYWINgJ3wfUCLq3GqsaHF/fbBkt9IhnIBj0YvlMm
1hpYBFclVTUHHrGjSGhsKdPt8Hty51XWNMkscKEtyUPwu+wTNtAA/TdlHb1SlAv7NvhF99YB0ZwB
CmVOw/PCpQMBVI8D9oCd8QFrg9hp9K63p/k2QAUPoP9hi1G6In6i5X+FXoeNb6OIc9H92hxXlGJe
FQNUR6xBleNqN50JgO+nwHhE0bSJYtfu0C/9hMLgTd9hUnVOQQd+G0gJ6bjqVrxbeCzpsOs9hM9e
AtjdjzrlNJA+AnSTpg0kioxXxmEWTAbo/tMSqcbgQNODOSqvGJR2a/zuPAnj7xwaoQUsZQc9Rqvf
LMpBkkA3Sl6dWVImHKYXU08T7yG7hRLTBIOig177SB2Q7sT9phZ7+ildbYUiBKWULYf06r/0uj2P
V4RBgGrfKXJt2WefnHRQeMaHn6s4Z/irgbQozM0Bqa3aR722qr8hMorEo2g5uYkWflXzq3F41cwE
LFYIUQQMJO1gYBH1BqrKN9TYksP4p4bE29j//alJ3Tj7MGA31jXNPe7DgH1QlZqobAWIPOi+aR38
0po5lX1vCAz+5NN69ACfQgLscdKRY8OPyrHGay8xYOD32Kf2BpIMnHh/D1rDgIvug/1m7F6bebKH
nif339CDNNekB3+ACWYTNWhrJR0jPd9LfED8OdsNhG2fA7AUkusmmydLwzZc0OsNYol75zv7OY6E
xOzdIQFiwHSj2zRClypYF7UbRJh/ldgsyWPC7mKsnKVYciZv0epRYfHIZOmD0RSW6PxsLTC0U6vj
MqsOefh9iMiXvOfIxRBa22y3fi2/KGAcSVyuTZuAZlQjzKUfTViXDlc6Iu9wvP/KWcc0cKs0bsqK
zCrQw601lN99ue2fcNRn4LhZJGXCVrvfI55cOr5eLnLlZyykS/P32f0TfQIh3+m5YxoRhZjq3vk3
lHABv5p8UyXcwDqhnYGmcDzLcrdfDC9duMZpkf4rZ+rsPeJrcZeaGMprYg8r/HU2PH5xC1KbyMFb
ZKWhpbuCt3LI8Wxt0TK8c3zKXK9iPSy85I+okUyTXI817UvEnqR79jhExcmKS9Jjn6enqUYqg/uY
a+y+gIL9RUAcKUFY0nF3Ek1diEdwLpM3heIJD8/ySntjgO5pDhdVe7y8/y8Wfb3aku3ng4ODUbmE
E0c5lXkflrcLFOjbdKUZoO/zLf/vDr7DMPDSK/PrWa6aub/eciV6AoAYhLl8P9U+zGlW3vy2HtcY
6TymMASdBFp+CZJ42yI3PwouvkKX3nDAIs8wHxF0d4AzhxF5M92zLXgAQ1vLAJrweUI7vq0dKEw7
jE+LVZetYKYp/kv2PhyOMXwqBdELbeIee3/ez2SD+plnryeiijQBrm0QTuexWT3s529zD7MGswIE
m0hOQ5AiQ5XhyBrFVdTFMQlVP4I28PR+rT0Jdbyg6E7/FOTX2THaEIEUnw5BGFD6TJzMj+qjDewu
wwhpwH24ZGxu9KrTGvsH5NJxQNwXB1hgeR/XHKaIKariIxN1udq8YQtkIRl7vdHTdl1vf9OjajYf
t9AEMqb6tXWXOz7cQu0Endma+Kf+vso3we/yNNupHBbqR81TZ7iAtPGW8liy8Bjc8LpStOqM6Bby
8eyW2WS0O2c4qLY4kq8BwvrVKs/wvyTWOk2PXF4HFThz1YX5gWI2jp/cdPtzmRn1tc5mO/S5DTKR
zZG+zoh11yC8Dy2ByrhPsY8SDrpUityd0U2VNILRNoOMRa7SqCtPeS07fG8H5gjb1yzSwUoQVtFp
ATFMHjkFJseb704xPKG6sfbdcRsaL0h0FxfGhY2AlwqKGag9M/58o0AkiN1kNb7F8VtVH0y9A8qw
ZR6B7C0sQLxmPMNIrshqadJZVzo68iOWPfKUGPsLO2Nyn/FKEL1aMS4y/hy1LeB8ctCsJhgsyLRb
h/FpZeudgXYKrmDg/iwZ3DIn0Lj1gT9s9U4WzAftxLeyNvuXDaTBq2WGjfsfU+GvOEVr0Xqrt2bi
u55oMH66kyr6B+Bd2ZohhTWQvWAZlqvUtExbGFy8q/BHomuUKhQ2fU7emSA+EsvKeLhtuob1x9bM
ptgu2bCBRcIfa+wAN3I4tPBBgTQ+1w+ehFwNLCJX0RRpVEeww2agvYpBotz0S1w1RSeA7svDpQUj
laAKgT3wqiULOOv6RkX3YLHfNKYbTIfeuzENyDtszvAVzunOXNjkhiIF7uxxJdzggg4UuFl3Y1E6
8X/m3GHNGkFHbYlQeb0hkkYEj7NBf+rJv6EPUgYBy65/ZDJZhRNbeFEOZrrpre6X9g87BNLFJTxH
OsYHydsW2gWTgPIDmeU0FpdoFxfU0qs0yAK3f1i+cjEU+hO+pQ21ASDqB0SrMyTrtgG+UysTKnV6
uouUMjxeqMuZqjCw26YS5MlPGk84mSw+E77qrUn1URnaxYwpeKcVL7AFjkr4anv1zQ9fTM7M/dSb
sdNJOEyi+P8eYRZjSJPqwJ9xx7u6D6wVEsLSdVNaGT5HxhH+R/iwTWEJIHzZ2khXIX9NtXzhcw/5
jaB1KO/uGBMeQKUuBKWYgo3oreetsmskD2+PmC9lwa+2EK0a7h9UIxi7c0aiH4Z+8r3x2U9io/8u
0zs85a27mB3CzTAGrT0QbWkEq6hLooelBW+3cazdx7MPnYWh0kIG8yQGj7umbRIQrpQjvhHRGUTV
s7Pu5zorg2FIBW/Ai3p5WJD0OWHMxbK/bA1HeV78FDeZ9ekQrTZ71OCiLVJuOcSCk+rClpbNfdP3
OJMSfb4TIEr3QJ1NXicuhXkExDjziV1YrBTZ2tnWZ30L4p9fiAj7m9ULRhHnRSOg/dMqxiw4qmtN
pWLyHPTmIO1v/M/g6S30wX7/OLklq0PVD1HCgE8alUVILpBw4PIcgn8cGglTaU6rLnEMtYdRQWOH
mq89UTaBcIa43N8Q/hEthDJVPtyFDLM0wuavChzSyMc4s1ubzMLzMMn1+/nm+OiB5s1I9CdzMj1C
Xc8m2kn9ZqRQjeAM6A7oNq95ceEjSEUpHF9YM+9m4C09mXwsdJAdDfCCG6eY1MVh2hKc9ged0Upj
IO42u9Y7t5DrgAebfllVzPFRgkt/Rw+Ov+atKvzBvkyQS0k+GmgWexhcw5SCUVVJgW1dH07ayC1h
zhEtXoB1V/g0yIpAW+tUE5D2CFsfb+kGdsgf8N3Hgav8QD6+2YhGRFW7fRKi+0yL2K0S3lS8Bsl9
SFZm6OKqL6SoL5rvUJNwTmoh9MlMeAKp1KTD4yTtIqD+TP2RK97CFoX93KspRAhCSIaKJaZ7EsnZ
GyDO9Cen1NfhN/mCFoSSh8s26rbw6aTMN947P2wOksJ5QPCWknAS2hcnxeFsroslKuRvdgPNs5UZ
swi4hUicWEZme8VdPlSnZbLoEKXZEq9QXwQdM6EpxRthUJH14CancJb17L+QRdisUAJvBC2QA1a3
mCW5P2frIbS93T60pxBQOK1HEjpiWMH76q+V/v9laqUhwJTdkItDnjZiDI5KB9PxQdlexjgTI4Xh
8epD6q4/AkVu/5KW4yriQwN2eS2gSslKMX42yHTcbhgFoZWm1rEdZ109WzFdULjrN8ppjkTgHt3H
LudZnz2zWA+x94aZIQvyo8iUx4Re4RvwCJ8zshAHBcd0gR6V2UneRAK+L2y0/BA+cAbGOB+Y6OHJ
Rt1m9kTZwN/WX6vcIRrJohcA6VoqHWL282IufUKgm2e8vdTty3ZyviCOcGF+ZZ5IFc3cpA/mt4CQ
SWBDbp74IDGYHQEDvFPgkAKrHCSRoRQzb5TGatMv1v+8qBhUBkKaaV2bo7AvOVy++gPgr4yV9XGE
by41KEn4YgqNowZg15G0y6XARmGim4sTo0a/TmbsBbC6Eyx391hgNqHnYqVdUfG702hTE/Wew5pL
vZKng5FPxT63YerW54XLYcWY/kzG2cCIUFbbWSMNWj9OhkDG/d9I0TKk5IBU0icWwI4LvZpZA2pf
HIXTlbncHw33wzf3pV2FlvifFttK5xvR0dLRsSx3KnBqVlaHsO1SyW5p8D7M5UH5ij7PL2stbbD2
YTiTz1l+xLjQuJOrS9Nj/gkEZ02H/ivgKLaJsl5DiyjXCwZf7lNBg9VElyoKU3rhAHdKE/iKSA3p
46E21zZFWT9z5gKHftxmwma5XR8Q9x7zsmn201MTTrL/SIw6CVTSemM/Sk5PnNn8Ta5pALFtnH0r
cARaA55q+4dMlXQvbneckzNYQOl5agPmf/muuoXt5G6eYAUAy9IjXuxW1n9qSDS8jjP5S+9xtatN
XTm4M8EAKT3Ypc17q/lFxtMEnOySE2MQvtTYr9JQrgJ3zsGKwjCtgpGsSsiAvkrfio74tJD5yQTw
tUCJfLW/2R0usHMffdSBHIk0Vl+3dp0TUQzhjWtEANOPOG2uOg12lh6WyMrgEmsrWtvq5tmmlkXb
mqtcwofzzLQBJT7F48MOOoxoK2+//0t6DTWZunpaHUTocdn4a2pqLKTJaA9TIOwe6LGf1rc/4vqb
slAKP7K5obETTcdxVZxMP6z2Mzn8AsrNLOLQL7CqKvIVkFddB4n1nCxyVFqTBBcr2LHov8CSfdR4
dV7FevtQmZKeKESGwrLXWvOnh90BzJbX4uoCmqKW2LMr0V4sZ72JjsEU8QFAG+Lp+i1EYogElkgU
YlobSy/f794fHgfZ+DofPlqO6jhhavAQPyIPbhdG0iPEpWH6zAPWtcqzoLaEcjcCgk+Z/VNkEj1M
EISLUpBrFWE90WKGXvE5t9yNK9UQJN7JO1M3X0BZM+KKdMxPXG4lOYeg+5liUH8ajC+oK08oWfAv
FAU0z0Gk3tNLkGbG6vtsFEX57rURnE6A1vDtGBg1D1OSr1SpzenR5XRh/0oKAhwy9q3/NuCUwzvb
dpsBOhM7tSk9PFCLoZCa2gVtyFJ9zDiXb1zeEDldZUniEjxRZ3v50jxRUuAtNXqWbqmHNLPSFrhd
DBkt1no8RQ6Ju6NcIjUR3INLKVpjbI5V2uUb4YdSCC43MChOdxnYQ+GkkaQKbPnXu36Ptyq0TPpS
Ddm4Nzl19TrUXuxXzdS6zwGlTfHW3UJWrR8pRxLQxZxdTrNx+kyqLMqzKqGv2Ndo2jIN5r/frQbr
UCKNr1p0Ofa+tuLvByHrEzIUmvzrHaBkkf1ZZCFYeEEoRknbGrsG0XZ2BtFjQ929QuJt3Khmojmi
vNnMmowO9XN5/497Tun1Yl+nrXOy+thLz2K8ZWAsDov+zRuGeOR+WJ0LbCOUCVb/Ko+S8Ma6X5hJ
5Izhjd5lWngvEXjtyxYU4LRYrz+mrSPORBxkSibnWIGuJvNBYG/MOjHZB/hJKQEFjpgxaxbSF/aU
/S+9lmUNAEGG+EcjEDA50+F+gcLFpdaw2d0vIa5A51IKJl9RZEr+8DmE4DUV27SdMdmCftJvmc7E
A40ZtDTS1tS/pa3U8L/sVNiriKpOK1zoDLDUPZNVA4raRrTEs2Jr2rG53nkdlFGprZJSI5f9N2jx
mul83kuR4ki5qVyr8sMLCvekc4ha5E9eLzh9s49Zc5GfMgNFf/FZ89ApT/+8OMpGaQZ9WPFbClob
VTWA0GX+FFKqyE6Ya7PnxfuT1iecLvX4Mn4vnDlrloD1XiaGYfQ79bp7ScbE+bXi4lKla9kwKFZa
Q7YDc/sqMF43zBAuVPFDwLgzOXp2dMSgfW/l0yt+a73Ls2Tmvw9JJdWQyFkzs129YRSu6dk60Vtu
/elAhAa9ZPUOq1tMpjmUQh2RPJdDlXV8jwiHI6PNfOGjoWuXhbAsdbQG1kdNP+n/2LdC8//8YmIC
JaCiQQM63sMZxPECCqNJ5i1W1SnyI7fIs96fc9TohRZQuc7pdp0HPy/X7BQdsR9KlzBi7E0sXtOE
Y6fQTD5HaWAV60agTtWNXMHRYB8NImfCLQVy8lmSjBJGGY3rwiPqpnd6nCza9nd+saRtMbo2lK2u
PlbfLAOlHdkwMCp9tPtVMUTrXyfkZjwTWxraiEBd12dP/8/9AZjxsy2CF1nQBl54cMSSwxRD6bNh
DhUaWs16oSDXLWQ5g150J6/SimbfH91+OcWa0Jasnd8YRn/cluPakhLR2XP4wYBGlZNVWxSX9XHu
vJqLAMPowienNNJhhRotWfqrT3v65+yoaU1Wsiy6mUy5Bhi5rAES6f7PCs6G4l++PcTzxq8NzGG0
UVekbuGyh4FyMhpyqv2WjkRbG25nNMGn47AqKBsmhA81HI/Al4PzkWzwa8vqeNHanGf7w58wwwhX
7Wnld06YDeyUY+VSYQdG6x9oMIwmNk4tD7wZrrVNMOZz+DmuW0Z7CEbBP/FqkfozPsFt6hzvCwqj
AUGadavvWZtYFXQLXsx/FX3uZF2MI2dD/EcOjowBI1kyxly7hnqY/zthUeC2Tv1blc/uFFKo5KrQ
lgJwOU58Zw391ILK0onbTiW5tm4swSxWLrR3JcJnn9M4g71qcWXkWweYnBvyKHJ2CGG+HDFyRBFy
h903CcFOL1kPZwRQBJ8Rhb78Kl3bnHvQTBoL+4NuVYzuev0eVppXncDqTwoUoSycJr1faLZIq3Yo
UtOtS9F062B8s47Tw2E0cjkj22O7HI1ep7mFvXqGckVsWGXIfyxmBq9gWwgHUVbANSVLeoSt5RIv
0vSfMKAjinktqJTT4JbpeBTklyguAxwDQO0bmCC0P+gS8/MT6xBDPzc9ooCvO4VxkGny85suV8E5
Bon/IjA81JROloYUE9JSyuseyZkCGMNGGOkqmBOtdgd2vTcAXwMAd5gVbsfgNKNJcHIQK2P9yw1y
hNACKIi08/XtOo4BxKv69IwdORniRNCD6Bu05xNDZb+8mGmgL4GUO6p1MlU2ltsGh0U3HInuNEuv
AR1Kb6oUI1JE51p0zwwMUiTNFwkWamZz5c+9XhHUjM0TpwrJy0zM4wg8lCJVGHecZYqVOgscj+F/
auaY1zJqOgyElJm7/NBK2ZAtUnj6bge2QiFtUkVQxG6yLLGRoM3o5U1H9y8Na1L9/uxSeJo7nSM8
hUKaR8Vzrb9+7S28e3q+8zDGqhCSd91RkSderQiqU7qp2rXZVfJMMZiL1tTur4L+QfC3ypBlOb6b
vmWxDv34Rj4HQ6RgUEHHD2tKdxj/UiS4YCPUXMKkkERGJkWDyKMpgDgV3jsgZ9xpjCWIq5WqOz3z
vbLrP27jqvdC3s8vE1RFjz4s1dCpmcrXZSCJv9QrnBsfmdd62Jykb3vSDp0wLxT1i/GEt8GGxz1U
x3TR99n15e7Z3xE990Tf1X/B1gGrjiJZpqwjIPUo3faiYT+aX7JfHgFoEj4eVKoYW+gd4zdaI02Z
wLrwYfWnKkTuZHIWwmqwNReCDr8MNdlTr5OuN4ldTk/Nih8TdGb8iC2y5OqGvP6slHRA+HzCsOxb
kJDzb3KVIuVPoWXw6c1x/5cG1QXz9xEkz6iIo/R/w6sUMnIvMQ1xnw8B0GK7Km+VKY3DRxuyX2v6
pDKke+atYjZIeJ7FSkC+uo6bMV1JfH8nFK6nh2NDjfwe7U6uYpCjkzL9pWPtabP5HsUjwlNE7by5
Zgh78y2SoA1wWUS2Cf3xbEFtmHNugM6HCr3EMG8OqJOfNg9M//iqqCIzJ6il9FZMChn7YWVBr0qi
EG2epvAYWQdOUbHL/SMh+U/5iD70CwNgX2Ik+SvvGFugZ8YalwYUBIjUGao+SCVa8IKMTQjYWTqd
/y2RZBk507rA1/golnbOYb+AC76iD0l2fgtFLDVn9EWZdYAP9rNt2HMcJZuje5iknrXPzG8+lNaJ
bUBl9OY3MYVlbZkhfVO7I9Zvd/DZ2+JKkKPVyd2f54uYGTbyIeEDIdepx98WFMoHQqDL106aOWoD
vWgRYks76U3jVOXJTRac/3FWdPssNpf7qMI6+eiKLBok5+0ZaUXk5FRvZLTkZSohrYNgzm7o2ofL
2Wae6OfDfI7HRkd94vXmWpekhuS76OPJ/eYHFg2b2k5msDkPYkYGClzTCkja+OLnqqRhq2ohtTHI
divA7AafHGY6/aC8Bu/pwVLfjjs8GakumXaXR2/1OKgRY/dygXvWyi6pkl/6XQmZ0K3vy51nnH67
DfmbUYEom+beThlfmmzP7NZHhacynNhNn4WdRm2y5plwOlolM5V3iLZpFnLmfXJibiRy0XmBVFF2
zC4D0dStaMmsB7W1Nug2hp1+L7phuze86Sx/OnlmyXgCvKYTvndfSkA18DlPikDdBjCKdbfN+zmQ
ItU1KsnVupMqdjpacvUFU4xYlwUaLBrFtyTSi/J7xQdUBjT+oDZHhvyuuK75Tm7lTiF2F4N9On4e
/TKuHAZ+exWVwaRCXaS5ovVO51xriUGbuQjx/AQFW2YsApVAHBN9ueVLV+daSghaTcpoTaNcDAxg
z5hOP3PAeQTv5Jjkx//J733FCYg273IB939mORbyYRu72lNSRZcKSfGg6UG54a92+y5au2EOm8g9
8kzEgA2bTz1Db2Jz3WT2nExOwW8TQdb1hIdw5chG3o7NWFNAO+6PCIzR55zgzmbiPEtWtSIXmQG2
w29nwqtJoyQ1l7Sdld01Vm7c26UgC4xDe87Afdls20bdzxV6i2jHC9xB0TS1Gw8Q+7f5t4t2DTpz
rPy4qU6iyMIN2lhxji9PWRrN25j48O6Wn0GNRq8pom3TYKbsy28uUW9P03DhTZS5WdJCu3atqMCD
9s5c+88n1Sd9zA9t2eSAxRnn8XdBhhxhfyMXg3SBXyiBHgzFaH7LkWjZGcNh8QD3wvDtAPCNVqEl
hSXqvz/Mdh8+greBgp+QKNbPbOZaibLYhYG9HnKsQ9+YZb0AohldvauFUr/k/Aqf+L957mfB50+K
cD8bKYJcxr03tl/YiReK9EfvutDfjRYjv8lR8LXWu+u1sp2fVcF0xC15sSyL3CCmtz1UtZciszZN
mE0dThESYiGVdVhLoiK7WtcWPBqlkPDGLNGuw1ZzSNLUNQZe8fTcqRVQcEoIQGijpya03UW2sGDW
8lf/JHQHzPgJ2s+J36MoQbkU3wIhaMpPBgBlLvYtgOTFnGrAt8XDkGAv0jCEzuRr/shbTO/36PNd
7UKa3QvLn8Rx1O7tNGTWqF55yQ8aRUMr9E+SV8PaJgEP1sSiLJHvkwVwYu2CyL7ySpjx9yI5lZC3
v0Di7JmBVSLK2yPS7BpWssUvoYQAIwiz0vWIjjlAOzgxEXQvheY0QI0HcxZvTOb5+Tma6X/mRyEj
LltIpYNlkV9rqivuMvEu5Xrsb0N6kTkOzU2QUrwZ4D0WREdRVOsNw+lmgRkGa64MKmfKwGYZl2s8
EAy2MJWyfhfj7ybd28czAr0T+mt5+IFv6IIVjQjxUWOmha6sqffxyqE1TRs3Kx09hwFmvK5UqICX
h+WkLcTZzLXZaZXdXYni7B7vbcoZ9UmQSHllxbACkZfl2cVdItIboIvo1VN76ND2/OZ4WxGhardz
hON2UcCdTXeaGMrU70lBfPn/xmss0ZpCj+JwK78qeq0WTC28Vxozcl7Sl5EA0n3FPT2Irn2Q3C/d
v1dyExuw/RDaAi6TfJ1mXG/hTRVLPKfmbymApfG/pNZXOCK4UZdHWr4I/SaraVul6hJ3T/KszOgi
g39pPjHn+mzHvIcVFjd7JZkqiipmbFfDez9dB8igSO6GO/CaLpoSUx1fIrcNNzf4XSguyj0O7ASc
NXxIIrXs+rf9D6IY+pQn7HCfp1rWWnb5BAn26TDgiaZr+/xh2sEb8Yn0Nq5YGvoJHv3qNPhwGjG+
dlOrU0xGDcglIq7ijc+LjXrTpSrlakUP1yZpBNmmS4V6tpOBT+ZbrS0AztfJolz/K0cMLXSRqcmB
QplBTH9VpIEWPR0EYpLSP7i8DDCjIOQ/vABmqeDRv/ilw53w+qeAjYDWa8ZzWJ21+oMyPVA13Wbk
ohb2rdb0v5a2vZ2Z/xQSSuvB3sFeOqjERZj5827otyA1HEumQWkcP6OMjyv1y3ulWqatzKf+ZT9C
5S1Og/g4DRychKFZjAbhBpyQtz1doYYimgqdDiiQG5dz8/lXuXQATItItdZo5xKyQ9aTZBWcnQa3
CznA4r6gjZut6Ism7ehAsxudvTw/lLLuQZh4loz1DFC3dgHd4MLWnvGQMGCJWCmILITdhOWqR7GB
4rF8an9jm4bfCWUaVgfrMt9OVrnGypga7D6cwylur9iNCvPwm4joY0rPpljawT2l40tRVKo9BsrU
V5hxFeJ9/Yq0YHlOyGSQNGgwMpb2+eRiViGpl6HPmSMGUN8wQhOsio9GBtv7AFABaRlCYMNaHn0f
4x0BdHYxV0Y5HtMgSMqPkA8i2ZADfPZhSsZSELFK8cPQm6tvIdanVgmRY154kzL/cYXWdELYJjjY
UDXKUIBuKRUVKpxBx0XcgB6mHUGVII87i3+z5T73L2By2op5aPYY8LONSc3vSF0EyOGQV9E012Cp
i7LeFPN61aGta5PSLAfw7ztHzcNnDdVCM/mFKntg6fFvFvMivQzWNabLn2nA+QVxEbQ53nCRXYFY
pTEs4RLbV9TGgr4rsIPF9FOPIjwh+5PqmzBsmy/zZuFkL9yu1GcjKGG016TLUHeLO+w2Ph4PsXza
j9ROYu+LkOjlI07ijc/JF9E2wy025ORkyq1B4jLZZ1+k5XQYMWq6MW12RG9sDUKVs9wXYLeusj3s
qye8FeBz/+MbDZIO4pkrboDsYmsmttUraPkxcciNYBOCGWjWY+dOpk5+50GXBGDihFqKn5krkQiy
QkvWd+tYNgE41mVyGX8L/NgCmipg5+0SPDWGCdclwdLLxtJdrTNrd6QM+ZseSZJJT5y6Y5kNzT93
KoBSeq+QULBC2x6pHTUS7tZqmR0KFLe3eMWFwdf0+l5kas2ZyX8/jTl8+c0CjWqj717V4AEP6Tf4
c7CmdGuXk34X3XlTy+FPJ8H/2l2TqIBUaHR9RvBI463XIIzBtxaoI8OnLIOzom8jxs6HUqPbTkas
fgFJwzCQPzGTDgaqdTyU/k9/9sfzIHVQBQdML60XiVBzetB1Y59quBj2VdLwxAPjFvSH56rIJfBB
K2tSAzH7KK7QorwKEI6oGm8vgaHTvprogIDL3biNyTut7+etr/hoJw+GT20R4qppUffrG+ISak+Y
xtoTrM1wZHNmSt3HNGBj6AmjRz9SbtiJ/fWOX6XlAznPB4UQchule1sCNL1im/0KCAQIiDC+Bi7t
/JC2Q8zA97V4x7C0ZLmdUAlsSh4oLZQX0B6MyWnPug82uPs5cmjwi43LDlcOQ+egwIJAwJ96wP6K
/eY+497xO9D/yjH94jI9v+8OnuIj83k3XTpziISizie69OKIMYiBxtCh8NfRVHKn4aSqe4Zft2ln
+RDeXacxcN3CohrbfwhdIWgjvjj2KG+AW11VxJBG2VWJ7WRAcVgwhdUekDZOfXd0gh7RLZFpyqKT
SJNmBUlHgk+cXRs3lJ7c7TrLg+2z4iThy8vkd0ubDCEoQ2g4KOVdJvvMBHXnid7gGHHuBPLlWhD1
Oqu/j0xhIjFlBiXDbTDZoa4/gJoQQAwFh0kAPANRmbWBihbwWKw4YNt4KVemkYJ7F18XZ2oro6Hj
M/JdZLm8HEgLVxUIzzXXKeMUUl5N/zWXjVVI64wc8xOEzVMLjRcZZ8N+tZYKbOyyPUpPhGfiEEw0
GPmDLiCKfkzfyd+aYyHtHyxYwKGyi4aDN6/XfNJ15C8iuVGU67io/ReD70gqUSPSF8oD7Jz3tNxi
Da27ohzCwgAZTJ9awjOoDkYWSyAwwaeBqW9UQyO2SoayNhfSQzL34y6ud7V8Gms/iNoVwUsYtSPD
Uv1+4+SlqvN3OFRR16/2O7GMNlWCB5jG1fXUugkpvMNs0QBqt8yXugnXR/Fdxg8fMFOHn8zWJDVA
jF18otI3FFoWirIa3hj5fXF75Eny4eTQxgUSh0nPrzliZrHTa42Qcpgrstmty/7b5SUF4vOJf4qk
Tt6tCz8PazSSKwZLHn0vjaEFF/f06Tpe9FyJEhFk10A1jsXgUk+ShmDXdJ6BrgKydSWWNjEzQchl
KvwI2i70oYO+3XASVLr4oSpYTKwnUcbtlicp/Y9/SYIuFlD46U46Dhq5dWC2i9zfAhPjhscLGn08
CamyYinIx/7V6I6FDg+fGvH0Fbt2/WZb3G5XrEdPWcSewNYCzJB1XfcV5zEiqGGv5+QFfL87My4c
rz8neHmhxqz7N2gy+E9karikSaRdUATHCFCQ6TK4sDJvT26IzYdJNvQEaulYWUgZlOlqSB+CC7kd
+66Yz5ukZyUgpXvQjzZ6j+zonHc5ZwmjvlaNsMR9yiFQ+P8M+2IKSuHqH1s+fCQPB4SnN14z0YrD
fL9+XChkkFlHih0ItjXfxyZHV05EL+AlAN7DziUbGcswkZg66PYcEgRfaZkjcFOw66bu/P4BfUmh
E1W0DSBo7Jlgke9IkTbnqScm5vPs9BmCRQJCzBu9fyW3fLssj2AxZixe9EE1TrO4t0JNs+Qm8i09
WMoh+EMJWXqeLw60utDxxpmv+cgA2QGrOuoVnw8TFMabzU8BgHuP2nqHXebsy4syVVBwgexXTpkT
6qHTat7Jes3tbdpJeDy6drRbVw57KXXoYMYrvDX69ouoQ/X4AZ98jctgtVNoxyAmHM9yd4JDRpj+
CXUPNl1jPvuBjVRop8cRd4AhzqBlv77WJzY5ZXhhXbc4J3nDmKGqjK54uVQusfshQNOJsY9yLA2o
ec2KhEJdRcoU4BC0broSq6ISQPXXlxCpY1VNv1ByVx/1+0yGSleCYQzf6fxiUPnrbNW1pjl9e+dx
ohpDkMoaPR3u4ftd3MTRm1fHsZi5ebXgFvhUX34O5zJuFLQv5L/b2UC8Yrd5AHZ7XXZrcotUxghS
MWs0u4603VWr40DuEKLp6L59K8azsDj0DrIki/oOXK68jZ2ZtZz96liF/2vjQCZiu+0IvSt/+oXa
/G9qxQfbcD467QszmNAHIhyxQzEtNTradzvx6DQZwqgDiWsNqw67PpJoRamz6w/+qwZIsuZQCAih
j0rfrX1GHuMZ7hJxQ56PAG+tWLFQFwhT+KfZmNvm3c+m4DN8qzs5Wc4+QBJuAa3P7iFUH19KOR3U
kJzbpOpMcb6xqdRollUgAxJ7wLPQkV9uPhlfk8S6NdK93Dt5qwupKipqk3X9GB8UVezOvA9ExL5H
b9GB5RFoGxHY+IysHI+NjL0Uo6DC0Zr/xwMixIb3hczc7WESvSmShyN6dqKdZIDfh6HzJgR1HUfY
o4vFFP8Kuak5AEPJEb8pz1sWH3yo2sGe+W7/4YprItS6P8uLcSTyT52DPNuY6g4nMXb4z1Ukma4s
UQyAElJsjboKe6rKyvnJGq8z3xzGmjGqaAWLTQz0Cnw1KF+FNrH5LFb4sKFDc3zbjY1Bwe8Mk4Xi
9ssq8wxWVB+Plifw59K2eil82HpoxftWFCL9wlaP9nCUFJJ51567C/R4AGTFTr6kAveCM4Db2R1B
MAN/2Iu4OcjoCPSeh51X0VaSsvz8HkuTqCYjeavqkawMQZUSH/QtYW7ISTNwUNgZZUDUvvOP46LG
CkmaEATYLnaXgejlTmvMVxKXuPEnNMY/9sDfbAgUWjd5J5/YFDkudWhHH6DLCK2IGbNtllKnKAzh
W4kEGJ83lSHhgPRhboNzn4gpStcOamGopZB5U8nVUPfN4XjYsB2iZWpvMsnbszFVW7nGjTE3qMLf
WILVoRiJ/IAQMAQNV9ZRwLIm1tScPpy2HdT0mOJZfX7PIstDO/2JIjb9gcaHhe8x+8A/iuL3Q7kg
YOkhMyZ5ZkGkPjDcnjhKv8x2PPZe/21q599MJPrrTNnIgJelnqbXia7iNRyYEXjgid8n2GB81jsb
WROwZCvEh0OFKBr3VJIKpYeev4MVekrEW4WNyM3vkuibhmoGRJWzUs02Cr3u4/rfpOJyXfUZVx31
Lxvlef0rvOEviNKSieEf/zQpscU5vqgtT+0NydW1xtlcRgEVF6voQ7eWromDZ1ZUeYHuBEyFCJ6z
q8BpQCAktUe7XUfXcLRJa6TZ6zNPbLiZDSCgtFLmYXWxm51PNoytRmUZEAQFn031v6rBJ7bsOX0J
RNxSuSYSlwFe2/KHhuWhJ9N1Wyd98r1YPYLQVViVO50Psbe6WiN5OVXcC56zwavhchYywi92LP3a
zlxzvRh1VhQ1XLPYR2BV+Ll0DFIOMhL0Cf4WFL29J0/NJBrThUZifD2nn0XvsBxLJcPt05or/ZCF
GgusIvf+voG/dnhu+0w4lbgZ2thIM9go4sKFYbWXN0oLEprfEdwyzR8PMAxK2OvshStiaKBocfum
r3dIWVbnhmd4/hbevAlYjJA7ogTXiUlpoUB0AXBdTcr0nASquLxdiOplodNeHsA0ZBPCOeCnS7Ns
farATPArsIMJ6u1MVmSuoZ13dy9RxjazZkWrPNKwmPiki2+ujlMHuQNWT+8AituP5gBa3uXE4svp
ABL0KtPlmGYYtCsFtzaHeS1JTfTDmj3+F/IsInEHo60gdzuETr+U+Mhj0lIEBR9VfpGzF7OyD+/I
/PR1sXn30iue+3mv3gM0+M0i3IkjQPYn9ch5C+RxFkxBfjVSllb2kEeKh0R8fgIhMTfZ8hmN1K+v
tbEKObkZhI79mSEZEwCz0bca9WbY3G/8OHbDFEt09zG29fbn9vDtTIYPXfiKFJyh4h7AVKp4NeJD
7G8WnhjW6A8yvN62UoR+GL7Xu8gTbnBOqYV5QswCHLWJWyqtmFkX71LVVU6T9+WpOxSmYR9k9Uxk
vPG86Dce2HrwC+/zN/+nn9mB0b/TEai8trx2RnLe+uqxRxH1l2a/2ecflC7uZF5VAFz+qH4BQQY0
DUZI4U0kIF8BkRptmWGT56gFL83RRJ8JSMBukFoJPmoP9elvQtIuWQE1rwBqjvw1stx043cKLV1w
2QxNEJprCx7jU/rwoSEQUJuBSAZYQ0LHO4gbXSZrndmWAcQqA15nQZ90jrZ+LA26gR+Hjf3Wo7Hp
swHUvwF7uEaVUaasK8qIMns13BeF2hPYgkGeVvYND3sw/Y79mZ4Yb1dyv5yhN97RRY2X+IWNCzHF
VSxPmg5S6W9J4xJUcAnNLDAXL7qbhfzXyO+cgoUb/SmHKt6TdmgVdXwXMB1Y9/kM+jXi6Un9qqVP
DYwA0AdFT1+pCdsFfSjyaDBJX5kl6DUdxhWtKfXHy4jRuKYzKAOmZ1u+k2dIxk//axuz1fdb1m7A
Gnw4oL9IT+v9xz06gCepNO137vf+LqxhrCag2m4gGVb6MAH5yFrsXv8qg65B+WfvnRkWZMBY3fXc
Yf3ImpiS162wqBZWlb9V5WguRcaFkXKQDXmxjjjIv31AlnB7x42SpOdIP6cG5duDONjhndGsNjOC
gm1ye/enUp0zf7dMNPtEWhbd4I3uBo+tfiAGljz7NwAqxBDzq0iNIRKuhftK5Hcv9rlqb/Nosse8
h3BPP/fxjrIiH57UvzuZb6h4Cpvk/n4wpowgX96PcJh483qH68FdYoh/goa/oMkbYMAY468TLAdU
B2oyTQnlvjNHS785Mn+KzCd8jsscXlkEaTIHggp5jogg/beazKVUrn6m9bwwOEc6+/SFtXH2yX1R
mR1zqjPWX2hRWcgLXP6CjidoRFJtVAQiWEAaEDKE9eFzCtrMmfwgs8p2w0OPXn+EwUT9G0mT41yt
dduozbfbeVNkQbPz/JCfHyLxJ7zeYr7SywJvn4Pgg7/g9vV90M2PFDimLCpAxJOMxI8NaOqpHA6+
rcA1rUvLAFj1ErGtRp+evx4a0m4NQiMF8qXZRfP1ELzITRIjdZV5fVcjvxdUVPh0pabkioAqKs5h
jB8OUnIIAzTlt93L0Owk2R2ApTInVED7137EPXzkMmLJp9syDiXaZU2yKZN/cE1YQnXbot6QAsGb
i1SrEJpwuvM6Y/uyYwKPcyzLg3Nh9babLbzmTibJNs8lupI76utmbELVhVYFJIWhhVaY+wQ2iUTs
rv34iN9tK08JcCjCnEqtSDOdOoAIHxOBY88IQyghT0Z3JOlBz5DIy+7scl8M484RpOhwvl2vqBvy
IvOMNxLR+i2c/gUwdptxLq50rj2sgvdUeDZ4yZCm4xUF2GGph6lNHMicBY15bkEdUIUPKgoP1XPa
Cs0gOSEnnr2SJJkZcp+U53BkxATnPeYDbyGeWngpogYYCDVBUXrmmcAkLP6Ysp/+LNeOKNzgskYD
ev6bYcEgwi7rWnPcOWWAgLsCFwsi9EQ4kfCut2vMElXptikUy2hAaBlJLqT6tw/SNEPWxkXyabYP
Zz/BjNIM1K61rMFsb6r6Pb/P5RAwhtIXFoWFLI5LwXcMzu6oyAFgPAOACbc8eBSKnLOpEKstdPPH
PXVJMCiy9mxWgm0+tPXoxWWIxBXjgLAaeLZ2x56H/HBnIXri4Fh7zW777wk4iLBfzLkjlNkGurNf
tgQ+T/ZmkbD9it+9/aTHtgfKu0SZs0J9Wp/CohL6eW9V8q1OLjUxi7IVbbrFZ/TWG0zHUjU+SRq8
sVTLgxXKRKfzyadRCBid+RMezIsBEUneVFRZyBnnbeSuzXqmq+OmjoWN8KT565kdQxEHJeqbPBVy
OE7r+9s+1iOA9yWszPBGM5WSj7Qx0Bifqd5JolAMBEI1wsVdUWNlDa4j9yTI0dbpKLy3XKzmORG7
45eoYsEZW8Us1nJqWnktQIpvVdEGzrSnegnuBweCzWjiFHyfK7G1y5kariqqV97w40WPXX7rSCMV
YYxEHDmWEA4d7caFq6+puQHWvJwxc0ab8DcHr1nvZAXdzB0L7FjJ0CsFFhW2u22YMvS3mIk1CSlZ
HFzoAskI4qcorfN3l6txhr/pc2M5m1v/hCSexyDCcpOpyEkbxj9xLd1hdFxGqNerwQG3EHxWtXHx
cmunrtgep/dvLcHMU0UOB6lZNRAzQ9qCwI65sHJnwsV9VWeDwq68FA98pn3Z1Eos4rZDEz313r6x
eRHTAFlsWj/QB9JwlrgKx1GOZu/ofTEN8KDC+5aECm1bsOBqsMCaRYJZHmP0as8TBS1fg1XnzKXb
B0qWEb10Jv2cbGSWoFVaoCawYdEnSiuOb/vxEf1dzyDp9ccHn2GPt2dcqaz41opLHqw+BUG9Tq9I
XBbWUas4DNjczRKKwMLybxTysCWjjq6PLG8j7x0m4d8KXJobSihkzPgwendrjO7mgcSdzWLmAC9U
yA28+bYtB8qsSGr+KxOF7VN/IZ0+iys5QCfUMgUv9nUYI5IdNvo1XnseKdQXePwFeKcVouSgeJSX
UQ84/Z62V64Ib/5DUe71TJYkcplsc8nXyNnZJQft2oWg0QY+mzY5nxR5H1DzC6vaUaaJdpyDqJ+E
jyb+NX1mYE9mzCqeZP96pgs/nQk5NwuRDlQG1x/LTsQITZ6VYA8OjXOMKDO8Qe+feWHLfMqsXxHZ
LgvREXPXuJY7p9g+lj8z6cfI6vB+K/te9ZggNiOYrFgPYWZOXQT4yNZi+hHP7MFII1Y0PlEXfWxW
OaKFc+7lJF0xDMxbXGO4UWANXf0O69KiY+BseJEk1CzBS/6YCgseufp97ueMgdikhXXEbQxFnwu6
vzI0nSaz8T0nk+8q98nxK3cMBhYT+93E8GS4aNNzmGl7D5FhmG8bylMTwBET9ElwNPFwyyLz0AR7
9/+h3lksCT9QIlfL5ovHI+ijLkP/sVx5Hhs2MfeT0FnRh0tZ09KDOPBqvpoEX8I9ThAfjzH318Ps
a5j9zTXCEOHZpfOclGX1yzZTsq+5ih6BWr4hSDh9i+PzvSlxHkHS6UXhbotPNmNQpGAS6nq1Dkyd
KPusEUShhKeqRdM+PbwD1g0FRp+3/vulMG8NDiAe/sFYzv37rbvrJZ/gnlYfnGUnb5hXw2KOSPSk
Qn33VXEVs2mwt1Z65rGZ8Y+R7RJ1rN0u3VcKjn4u4rEVDgfah+Np8I/nV4x3TIiV0Zs7l5/1EFnb
VBzNxMmsdkT0O7P4+tSPVNyZy6E0VfBgbl+bOwoN88FFE4BntcWGT7c0GVS0w+z4SgqOSPtcOh8Y
s76MlVO2dMr9h7o8Nu40HuddGDFF2oBIkSgRvrHcZZm5ZaqbkBJt4qjRybTkJp2Bl83EgcFjnRuU
LQFfoCpQXNToD0fB3t/aSR41S/H/8IN+yacE0IXaMop4th2zaYmeqOX1AayaU2jfCaWBzY+lqqKj
oCRZqRQElCPLJAeNUlUEe8Q/J3YhaOewaMj6JBLPMXqOeqEy2/JEel8SBHVBqxw6Vy9kTvym/WU5
WpnuJnBE0WZaGVGhcxx22xvfyFF8azXqraHLgAwQ+qcNqN64lu0NvYX4aHo0txOHg0FsmdSoU5Zb
3nMR2f0FjDu8rM0VMQMOx9pnAhKUCr/3xBE6q3SW6KgmezZ6LRHpXmIEDvRevlTnzBWC/d1B5NG+
77DubgErTgOf8mO3hWQV1Cb8uDIdbMe8SZPmMz12gugFTZLnxsHjwEw3gLrEtQPn13PRQ5edxZS8
p9w7ggrvjOMvCnPW8C+JiM7CmqiHJVnhZLhQauEbHzTrMWcSPm/Vn6BS52wBCYz7McZcs+A/AIrC
6dFJV66VVT/b4kI7hQ+w5VCTUmUYWsIZpPNhKRu155nxL72NotFqjp7R5LWR//7iw7ir2q8AaI9q
My5gmgPw+IAHrXkNPJPUVScwlvmOEpHep1tOibAo1aVQxbVdAEYfd8M4ArYwOd9BDW5+LPiLNrsA
zQTjKrQ8uGbvBDl8+zmXNuxBMKkeK2IgZSHhUIEBDlY9+BHJiU5S0RmU89G/YQ0TD/wOtG20ByLg
sjqGyPGhbTg6n2ECpnabou+uprt3oj0vUaZzceshrz+rFLYjGKQL3RCyQOZBtujh2xLUzAzHuDMd
+AI8aEkAk8vyiGVTHdV73NIoiiObgG72jYj5ddqD7Wyf/1Hdg/yEBy5aVe5jbNePZYROQJpe4+GJ
TqLBjVMVlsXnYq+vofo3xwsI5pDjCnGt7Dj1y++JNAuBGOkSVmHG5kM/0HTV1PgUBY3EoNfH4onW
65diX98podLvZovAPx0Jtj6Qz0xX3GsVEKllW56/9tmtLj6CkJDSWIhsuxqiz6DMxIhW1IfUqdok
TGPAmpFroh3Ugpm2HD3lM6kThbUd+3OMicJdmxcWt2DU3OHCWEh++U3jkyMFcLxKGQvUwErNcNPU
7R+dLGTQsXQj95T2cINPlzmFYSQx3C0jsTLL4+AGJV84NPcYhBh63ud5xZfeEZ7UZY2eIlJQzDbL
xpW/bX0TITOQdl3voHSFcspXOsqEEr+Pkd+ecRlXQiL00NFpm603Bkk2BH6kI9OBzk+/0acJykBJ
cAP5G2XzOoaLude5RlKLb3EaaKyW0oHPgRgXRzzaHJJ2lVGSLgg9FznuZUYf9THqdWkK+6b4d/O3
5jjZI9swAfV1XuhLfi4eCQ1lq4OqsD0FYzfa+36Po1n36lXkRTBghcfLNBNnHs5/QwDku5s75+s6
v3zWFlrjlkk2hsIfpy745tK0YhzUVpiqemEVfBugaPgRaU4mlF0tEE2nEH2Uk2qVtMtPALSkpkvk
bVyJ2/ZYSrbED+HQ3W1unUdn0R44NK2UNC8BDAtXDpR37hXXpf+/Qu2J6kf36xOVeYyQTrTjicK/
qd5dRwTwwMfwiatk2gtAgtOfA5LX9pmpr+DrPkISHMBxkqPig1HSJyuc6N8L4rvGO9n9I/08PMrW
AD8/z/jua618/WZ+KCmCHEsFLJbxleU1AQDp40DJQI+Cgl/1IE6+4Jl9GS5gEYFjPXDZICLhff+m
k0OD0uMdKYtJzhZ/rC5VkY7jAhCKNhGU+Pqty7piYufm5WxoqiRsrTMFjDgNUaWigiKfXzmEduqd
qs9wEbc8DaY/OM31utcK3gDGqxTX0lLjCHzuKOxE6AWaYAm/kaki1SCBHMcsm6U67reDwvwzavY+
6yoPEdvK8AyU/3MSfe6xZ1fblw0SlSNvbrExco3AfxTs/lY+XV0Uy8fZnOAfosFeRc1gB6d18SVe
JnpciOYwi6Z9mF1gXkFHBhx1rAP/Jv43lm/najVjtlvoiAS+495tx/EBMEl/4TbCuZlNlm4oOlcD
obaTgxOL9dCDRYD/oEvxwaSimRZu2+g3/fal8wIe4EJlY380LqBc9wIO1X7VtFVWSv2kVjayQG3r
paITXQVv3QlEJ+cZAVKw0xyJtno2fs3xkg0nMUHryLFItzWQMOBBG/LPvMu2MuaJHhx8CTwXLYzZ
7G8Td+C86DtliFIcw1Z/TcdZfS3rjN39mB9cT4uPw2XACm0Wxx0ynBheePvl/QbUYMAWhzM/NnU1
2I/WTCOpTGpsuEq1ck05TL/NhsugXDP53HBbT5REpJe+bqvDUz3Knzw1INnFfoJTx+fRR5JwM13M
LmTktq5m6O16d2jmH5VGa1pSjiMEK+k7ckuWQFDyrXp17iEr129pr+5R4dOtNWR8OipA9vWrVqwv
HwzL3VO7hg7doUpWbU9J8jLlE/cM0kMHPpPALTiPZKXa2m10Gobz0fWqhQ0S10nFAHAANviPlqrz
Wc8IY7VSY2hPWjN3HGOLjxU2OWvvlHuydCQzES5Tm8GYIM9tEf2cfoggW413P1/vLJPK1NWDZ6CO
VHsXsfaDLehzLAvk5h4TAhJ070Zj+2kWIBDYG7DdhQfiIE2Miot50ytCaeCd/28qUsqJPggbX3tv
anedDlGOwIYziu9YoCxjTgH2XHSAFcGs1pAqdQegAOUA38BZqa6DiGLweKfr3Mz9X1Bt/Hlc8W5z
DjGtsZxb0su4+8UKFu6ZpTIpYVoCrspBjXG6i3gTZl+YHGyvuU2nfTKs5dIQ6I+Y9DDruKYS3Ejh
I0TUpXYYl/YQQuzYUTB2Pw3KjntBJ9UJhhhYrEfRhrFpx1R3FgKPIxfaFOPnKdPT9I4zQmmrPp8T
QNGEZXbh3VJcMEzCLTAgOPgu6WNWims83kixbg2w320jvGRufqHnYqHci7eBmKoUbdBD5t/AXtCF
T2Rm0l/NWdAm4998K17Xshh/QIl50OXUtO7MuIP9sqUA+80LNUCFFHSSbY+5Uqac59fdGdvITQ0K
VLNKaBl1yjmqgO3H+3iNyh0JkexkYbjktV/o91w1RbkBm2jQhsiQTcBo4XxFAod+hanr6WK+pqfr
Pcm6oBHirM6f+vo6FxcJyhlnfUPkaYfbZu5G6jrZFzJeFqDS+p2CBq5V2kYdJlXrkjTLBNRYoF/9
EdaSM+OvB65fWTPwT5mm+svYQP0cR503DAeU12Jlz6GsZrFNDNsj746Io9hSMGL7NNKa4BQhQIMA
vWJ7z/HKslC2GFfTGvgBxrtSp0yWjHboFBJGHjYBBekdP0XCZOzH2frFgf6ALEBfASj6MgwvMYVS
04aMsLV8nH8Qnw6+/hqIZNOi5SqaeEzMb2qR/Lfn5HraQYUbfRDlGtmSVNXFew8ASJeY+dakS0hb
M8yLNKcC8xn/LiqlboWJXBhMJQi9pXjhqO/Ujjge5S+q17R1/UDzs3hry61Fkpte6aruOM6p/oUI
j/xdkDfJs2WasjnKsJ2mDUkBFhvn1aAdojYdii6RDbVOuSd/fryVPnx2tscHbmOBAopNiK87QNhe
lVaJ4P+H4tMlVzva/uEoZPRzoXbwP6yttq3vfnZPOy3K250G7ctXHPdZ3cqvOVVIpmOwJtzLgcn0
PFF6V+PEolCNJdvoL2TJDjAMwkfnY7w+7SuRMAyAUNMTeRdZJJ2yDZL0tHusKY/QaLehKZhq1iEN
FYNoNAhWV9w8jzxMfPFm8R9723OsFP+q9djgbeBWr22vpcLjI6pAwDu2oTn8ddgrwj4kjp3Mf19g
RCUsdwPNZJBbZQ9ZiqK00uMzBD2A5wT1VNDbzZvm9Z5+ib45QXtQKS0iNBhewzoe5PX5fBOuXUjw
hjNUo6iiCQW5VCjwDOsFBQvguubj1hBImkEmJqrC/FB+2WYpXaYcMMWclsfGJsF2VK9TK4VZ25g9
qXR7sgU+k7CIUoebToFJZWStVsB1ZHcoeKAi3aTAd3Cx9MPiHt+HZFlhKCYKt01hxN1NMhBZp2K8
Pbbz251G0riIV6DelA4Bh5gC4xB7m7Flm69eriXELhpHQVYLho4no3hDaIbZ1GybrwmdemO/kl8Z
NqPKZVi83GAJX7ZOcvyLvgP5Nq3WEaixXxFxaxDCHgHzgRITFn9imnT/6Pd0gSBmyHMjPOCYIKMX
3mAC2gqOo/sDwtrwzodNVw8V+MOiaW/au7CHq8ex7x1FZTE6Ud/fQTfDIZg2imdA6Q6g2OzM4fKg
AkhGDuU2G+6fsQCjjPKoRV6hMkE6z/8hlvdo67mARbv4j2SJWoGLYxxt9ijumhwSA0Js93Z1idGz
uiTaol3BbAppcZ1uQfW2WQc/Now6AL+TpOY/Jhhs7n2KQ8c8yYD/MIvBX8J1b5DJj/NAMV8fYyXf
c8K+aowwQYM6LOuixXqtbPoKDzUsE1TvqqENUzKZUMKteEzFqOXQ0X/5UG8qx1r6j7S1U74yMSaf
anIkGwL/IFRDiIe+CArqKf/h/+1h2u5fh56M37BEslqw8ZU3sitPo66tRktY58AVRZJqlywgCbmr
+TmAZ0ciBBceZmNiEICh713wAIzTygJB6hkbATtEv+iIJZ8zHdYOh3Q23lU9E8Z/lnO22cVM5B0y
VNnDMQ31glSl5wKCX3af3rn1U3LpsUm5qkxzTApEcZ1qvvUtgt+QC5ozdbHS8fSIX35maeExE9VT
TAsFszcayzSCvPCRbwwEsgYnRVjjnakZcnQVFI1ZGDBHHTqMnR3506tdEx98MMIwsPGnuh6Cu3Rj
DvhRmxGRGXUqAfbsgCxne5qDOilo4okdTtgwAQ4YjMry11pSaY5KQzk/VjmcYkdCfpPpAvQ5p9AE
bexgprdNcppkwt5U7EwRivedqasFvdzheaM6tiy3hPGMMuR0ltT9A/hVY6C/0FTR13cLgHu6IQcG
y4TR7qvjDCvAV+sy9uiSg5PwhEkRbT2sIAHvjHKjq1uQff9gkgDE9f+zSbRHNgXV0n/hmwVjL9TG
UQMAzYTa//IyRDyMVos5tWnCeqOki/dyFl1KxNmgf/Gt7B9iDwZOkEA6OB+sXLqQ1WHO9T1+5vZO
r70fLP53+4EFfnJDV7kdDdIUotLUt+1MZ8EFKrM1uVHI3vwDw9LuTvyd2Y49SAiypM1LoFylP+oA
hfXAeaeuKKHAa85pDYs2rB7rZlxbfD2yOiWkmEvL3PjRyp4J3uPeQFuyEK0b3wl3zcAvnVv/76tz
qxF+xc+P8jnDTZh2AQSCkRONOBSMfu5BSa+KdBz+TYcLRCsFm9fmxM/Q7k4+4FicPIE51sljzu5i
x4aS3PHFVSEyQWbqpxNzRUy8HDvBrpKEjCIDRVmoT+/d1eogEsaU3wQHIbBeR2FYBXKANMxL0U+T
6RVdTfpSkr8lXYstfULMSzdmiLID+HwZrfoAMHb5ROtTXYFm7F4SUoaCaGWnV6g2nyBCgl0X160Z
k3nZOTeCzn2/JlCW+r7VlW/MPboox23DWbLktMCy41fCMIm/p3xxX+CdAEqvmrpb7xMQXn630W2s
0ubRpbujxkXJ8gEbtdXzWYI74ju0QwNwK8O5+ilUNQ7YJVENwwE7zB6498DHOORx9lkNBalltrXP
GYckdGAa40neSao7O6/j277CsjpWRZO9XRqfcG5g2B+6/iXBcsxXMowbhvUpbStJSQmb8/iqjjg0
u6o2wfCE53Fh8E7SEfI2cJ5oxlLfXruTKex3H0lpbscL+XUSTSbmD5jTjA1ZPGoyruHlSb88z+vn
QOzRVqlHfSX3tfnvt1v+wDPu4hBPz6EoWAz5lAyedH1dgoHhCKu7coqzV5c3X+Ug8ApnoWu6lNiB
W2eweDDO/rEdmR4Rx5hKEejxaAsgwx8bFo7HL7AK0K65YNILVfLpQMZ9WO2oyRhiSkkICbgoRWT4
OIyUW+NDb18T9S7GoQ5jAi15brG4FEWEVjScyMGXxXZU+Pdm4sPR+/2itpNfqqUevpmRGg0d23Mv
DYgkiDj/a9I9L+IRwoFseh/sldkXxN/jAOKcrTNUnKnAnSXeL/X2Zzw6r+sC359P+GpDO+DWYtnu
PwgA4FFdjcJaEhFUtw0tvEXLBz5IWtKqZFna09UoAjGCqORX36LhlXUE5FrP9iiWa/7davK7dM8S
gs8WcCOxw64XYsoLfC/O/z+Kojo4bLHFXZWiqAcamB+cZy4zDgQIm5WVSbso3tvTgETOAIrBeP5/
hff87l/xkk6+6DxlglmKnAEq91cIXWSUX5AjpcBIiIu6PbfA5DWsaQ+4CWLieYi7Zc0YsVXJ4+r5
UIU8fUFYzYkpQs3NLZi7X9KC3cVwJtRUlcchATkpAsGshiQWgV1a15MqjfAAx5kz+hvusG5Oc7Bm
wkUCzlDJgsUvFiN4vzPmO60EExEy8L7TrBYm25nrU+GrzvK5PLE0ahGeoeWTTv/pcCSZMU9+Nrj3
K1nUH5XpdCsLZwHnMc/7JFUS/22W7T+75EPR5ksXDbyUFC69b83ZbdzQ9bbEKyWn5W69I1YdUx8J
pDbSKxHxCcoiC9d3jiptQMBKRBz+6LL3ZT54Ux7opvvtM6gbezoGc13poDDWClHqveVfwWfQVTm/
dbK/6qaQtIuizyW49Ba04VZFQN98hH5ofr/8bafv4/J3K/Mevgc08dDFi4jAAZDIIjg9kT05bOt7
NLAMG1j+OcsYDx/pXOarPUbi4rxRnm4tXN+V+czJprgNuGvi7PB8GkAD1IrlsVEOhCJvfvGG2gV6
ZpISopw6T7U5FpLQPPHc2BkkNAEm1tfRUx3Idu7O4UpNkxuvbygBxRbQ73AATOemRiJp1tqAKm3a
QvvUloScbroeppZ/RqRpky/sbMt+Iv2q+e9+Nt7XoApMUb0lKmtrQ0/HWfS23amlwDgsINjo2MqW
FmZkUS7/jPwVL11GbJRkHgPWEE1w9qggUz0lAehhB7FFkbhR8Bg5Pmd2WbRn+cwxRZZEOB3D+Ujp
U5WAH2KPlscpr/nW5nYOFUPsAaiIhlZoLHcodS5KawvjJ7cpsD7TIKsou/eehDaZ9ZPUUdGmqtbY
568xapfsxihPYP2kVQuzGrdqtdUjeZl4bMRVno34gf3MKgzeWU2f2Waah0Fby7nJ2WgFYS56MwnZ
M5CyPUzOGf27GEXb+JWzkJzUunNIRG6W8Qo35DwbfqXUGFVKKCiUYJrQymbPL03rcrpYgGY7POqA
5DptquZb6Uu8xGQla69YQtnnqzxlDUYdy0a0/th2qeIjyWbUZD0mTgmGagnn8b8Ajeiv2qmHRgnR
anAFla79DLEkhePtHBxdHu942m3HD4QFPUYb43V+p8t4+GQlnK3LPAEXguXxBBt0QRAxPJA4+yni
353/ABhdl+uk/zfAfQMQg8KoKErdmaQluhdgPjo5WaOEyXefpbnIf8ZGpQ7twfLafN6seF3mWvdq
MKxMAc4taET4bd8RCwmMvd6S6J1yIzM7PhuzJuzPCxSIKEVEcTt839lI91bgRQdO5+mWzdy1Tss7
dyY9zR+Dmlhgau4Tu/0dUki+rjE6ZdcuMtR5+Q91i02ng4LpGcM3XK6yyoji+se5XIEZlJqRmPlN
DN2FWtB8tVKAnxEgRJ211bRzyVIIBdUji+veRq0Ew2/Yc4CWn1uMSfFfyhdhJgtmi46fhUPkRZNI
Sna+3tI2zEU+NG297bVBJBCRt1Id2cqZSQxTbXWweWAyFJ8RS+oBHrtAVdWgGh87H+rUj6EbQUzI
UQtOAY3Mn7AE8/npV6AjV36hRzj8wZtOqatX56u+D/ztbm2Pk2WHMQ/FvX4I2UYmmyHmLipJ4b79
L8IA5XPcuvKKffRCFVTFV90fYOrb8kmjhYlLHCKZA5FgCS9B5glyr3BKvMX4Z5HRIhnMCfdYYG3p
AlvKyr99C8e28ZQdsiszysV6ay6Kp5EJI3BxzMv8C+IGy0qxWXVa3JHLTUYUCmpcHk0rBXvjzH/w
ClCf6elrIiiZWwFo3WkPF5ksQTxgIiGKvN+mJpk54xxl6b+RSAiUSRQpUh7AYsNi+7yu2dP5EZNx
b5Yj0Qw1nbKRk+7plyJiwQJQMrL9uRPGDpf6JMIo3i8leJHbi5pUuzO15vEKgRw1qLmDLQW+ssY7
FP1U8DwwMrj79j9DVTOiOcin8+tGRSh+DqnweNU1uuKLYZ0AQK6Kh7D7aNsnQMpQ5nEQbHVbz8qE
/u1AffnZdEfR9tPLmL8UpYXucy0K1oFg796mjse1+ujvx3wAVopIqbwJ2q3mWQ3QzBKF9dd3ANWD
qaAqrU/thIYQH/aKGFS+/0o8AXvkFBLUlXYv7AIlQL3AiS9RuZ3USxRjfl7qjLyz77TRlFDVSt/x
CX8SLX5F/MKgEWFYRbXG91FewK6ta5JrFdz2gTm8LTNkB6dpOJUS+x6FFFUUBwc+ZWNRjk0L0xD7
tsOVr6LnBAbecWzt79zkaLYm5XijJ3WEhRSMy///r0YUWUJxGs7aE/YvcoAeqHVwQ5wX0HZ8JgHD
cECr5T1jqhgxY8EpXSbBVFqdRlBXD7XnqFR3nlL1R/N89vc0icKawjO9pF4uvYiT0K3j6JocCXGl
SuwuBzD/hwVz/l/Fyn30cKXLm0/cb0HV9/nhy9e9wir8G4piDVg8QNFp0yquiPUIdUY1eQWxfF0X
5mrCPIy6ge6jAPKIczeL5WN0enONovborBgUb7SXAlJL2s+MxNyUltlTZMl03ANQBKWLIEzlkKIR
+84KVNCGs54zOrMaIbfpKrmfTJelLcAt1HTvrfrcny4tcbC372VRfadODjc3uGsEY5zF9A7jQulG
fhmHKaPG0kvcWfL7GZlyAeDy7Zk537WOzABZxLvmjnKyOcYBoVJyoNc3rKvIQnsvnxvSCUQ3piaq
0jiKY3NkSQB7b7ORBmc7Xd0WZfcdStJapDdW3esF1HuSSIq65gk2Shul312rP4CIC7hZORc9yPn8
Xv8qt0L8H5V90tLDxnBplUXqoyqRMnAQlgWjNpct+IDErVW9KLx6tkzmWRngzC/56EACDLQR7cCD
bfFtmkWYVO8t76T/gfBi0cgwC5NBjkVBx6M0pXlQmI2QAe22pC6p+8W8gq56xF4Q2VqvGPMFC+YR
Koy/XP8k3X0oIJ5+OwlK3jaRaj02kyj1KcMhtgK7duTIZDn5/79l+ugTdRX3WfBuX6kdLC5VPx81
y0ii07HSJO2tKssPlSF5Om+2riAonltVqLQroHQnA6BjjzaYslI2DxfCDWt0zQW/eJ88Om/MBWa9
nBdkGGj55jRT++8O8p+Bx8VvlTyLzoZobqXL7nN8mqIRp/0e1F7RVe19LUWny8CSdfOl7tkTyNAX
kidJTf9pfBEGa2i9WyAVCK8ysP1K+OdvBDVHIbkWxNBUOUF08aIq+e4UauBi5OlclTE95BdCD4pK
7JX7KaFdXkTn2nL3AOVs4bsjuu4VJD43GErSRhy+DU+2ZNKgrJc7YpjQe2hdLfM4bAbp0EJFDJ73
YfLH3hejcKRRU1KrnVtLefdjb6Do+WfWxhndV/OiVNiUMtfG126o+2t5omIsGxkgCAKyLA8VEGgA
ntQz6uAp1gE017UwknAp0qeMQklJ8QD7Q4aH4mdl7eFYCZdX36VdWzDiGuwW1dHzDT3C07daFto0
v5lW8xmdOYblwVELuxY8j6Hb25YyuuXNPstCVfYOlsiscl9K8I/AAijik2WfB1l9pCSJvZmQKFtC
wc1A3ykUxLOO9CNan9fQMI7Wp4bz0ZJvBBBIube0sG/cW9xXzcYakVm/CxXMv/LSiBDlr98h0J/H
29VCBCA7KD1MR8lQ2NF5cbTgybHIzLya06VMJtkKSTdrou8N7CUwRRLO6SBYYVSgLQgL0X6VZoFx
RHktYGoFTcrqoc/Z0xmiY3RSIqMP5JKPZ6Oh4qOrf7pLFwAx6CN4NBDxuz7kS1ZPGLhkxXT7jiON
gIDyr4FqM5Tv4KbxB2g3z5rd2S4KUkNp0/xLzN1ru4Xjl/rbN+N7d/njYYmHxV+jdUxAVp+jCD13
6Vqdg5nLfBYJEdf7GVq2+NzGs2mUiXIM2hg4nMHoIx0bO4MOyKowDiqIX6BqpVtpD3QupLiTOg/1
+pXd9X6ci7A/EPDJr8ou0u+5h94NikBElKkUu+U2RutIgWRKr7/TMCIo3YQrpglH3u0zPFZK3Fkw
ib8HbmLOgnDXvCnjOPCHTzavOmGko8FL9gmYnJmpXlh66lOmRZ7MGzdWY9iUOkBRe/nGFhmnmPHS
i6c3QDDhKgDRGTvhXNDPn/4nfIK440DmRzMC/yr3a3RR6wmnbX0wiKgBuS2ms3mFGQf5GW4Zbn/6
eCiCc9FBsYJdNN68CvmJKWF0OYp78tp3x4iIwh+uxkDP5t+gAYb1WSVnfB+OdD8VJDMpYgl/6rf7
pFHtl9nfaBSaw4JSdoQFYBPn1HX0w/n4ms812oatPTIl69LCk/vR6i9px32HKdeKqu4beX0kA+ub
S9iRcEOMN3LcLJ48P5khsjwQil163qtWMcJmI/upTKT4ADxkGkU79G2FVRPP6KgB9MFvr7oa6bwf
dnS5RPLAJv5YihPwOC6O7Hh2EVQyY1Roj+wUulZckxFXsxrhYSLyGmyyrgHxDDb2gQHn41nFlR3c
DfifIleVg9zXUvdjyB8/F6YoqUsSPrdInMwX7BwHQfXRT1LaidwTK91rea6/4XMPzRvYHMPdMwyt
MQvkROjMVCHhfeqAzRwxjyp0Kz4JzfIYY48rSD05lhZkvyIZCOVAH13s2aooV/+ZO64K1OgS0/I3
pBvyuA6CJOoWrqocQDZa/7ucY28Cp8UQW3wKW9fRE6axMnyjycbYITPyj8crOmm5q2p/MAj+o6GW
MPh5MHFltkQCmNYQCZJzU8bpC9nDdJ3k52MLDkmYoM1dshOzpVD3w77+Xy9Kj/FAImfeMe+sEHuX
5c1vpBv3GA+KYogHwuNrntdzc8dH7skMk+D+mfm+SBFY862eRiHNdwFpaX9d0WKiLf+KCoVjnJJ8
XHQ6lKHQxDnnXkQXwzGssg0Y5hKbbz8lxKkYszhftNrtcyqmLUVkcwxrGhsWxfwVoHcUeiiBkpyR
Ng7GdYX9uzKrocueiXohqk/q+fYz1Tvsmkt4xYgGWmNpC5E+gBgGnLkxtgClTwYkg8mqMNaw2s9e
UKdrxKWfXjqqnQ3xc2GLpDzARvcUEUCJFRkxGCidFQhMzMjEbou1+GMV+r2DA7GIoWea6OuhUX9V
QQuwJeVOX/M6OnaGznHbITOjwH4SZQvM4U9U551Ot2RasnV6Dg9ZNkLQ5cExbRACgxnz/yO49U9v
Gky6eqZVHWL/xPjRLCcAl6BToKr9X5ZTJlF1IOyB3s3Qb+XEC2TJ3jqmxnY6x9mPTX0FWCiYiuDJ
G54QT+KqrFD+SogcauZdD9J+IZ9lD8qJMpkNN6a4cJ0/tW7CDROg7QthAhnN6NHbi36VUmg2q6Rh
K5M5cihu1mQlKE+NZpB9ex4ekd2HCtHkY/w1kC9cpjEJ8OtAHrYCJaKDboy45aWdYbRokEb6EX5z
YOUipUjSHIQ7dLTLdvDlnnYhgEao1pi1YJSQpfKgbNFXFD4NwlOf1j5/HhpF06b8UAtWSYgrV+I2
cBx4MIPqylvr15QrhaM1k8DBcPSJBvk08rr4QMRHW10x4vNW37IJpMBWpoUszUnoXic/H3hcNuwf
F6RJsS65NliqhKLNu6nU9UYxX4EmqeJAo0GtEQiqEh4f3jrtY3wiud6ydvQRwN02tWxmj+lmIEhY
zbCqQ9OlwP4LT9Le6uMpCEqCQGGDyYTxZ89sA2yXhXcr/gnZjSrGrIPw3bp7LBW6y6MuyxWAVkp1
xN3e4tS8LoCKeU2KY1IuAsWeUKFqWggtfzr7vv83QEGjeDYMT5ujD1bD/RlVUn0bmtMgedYeqGv0
RLsxEDJW0oIn/7OdKFtWWhGU1YUhWOHdi8P23lH9DNjDXmyoWhLGzu2iq60O+f40T2hSfKFj2Mu7
6vhQ/Zt4oldCZUtIuVqOHeuzAPoq0CISulvgsnWaNqCgY4s5kWJNqR4tQLB2EwL5lx8BHoKkVP1O
qX9RB+WnIOp3iuFyE7p/9G1OKLraxaP0FANm9Q728g2o/oGWC2djgO778WIfoUfLJIliVr6aX49Z
hSfRL9Cr7nCePDuBTCzR0J6gW1ZWgfTVubTokLMA/jKYEYzpbXwCoUZ9yVhbksknfL+OYxhhJe5D
RLoZ3L4vlj+4AkCDHzUCZm9GI2rhqHW7QIOpY1nvxR+yVzUDMZKDZ+fNIGUJa2MkPIdlBDm8etKM
Bqnfww6Rf4Vq9vn6Dd81tlCBn+eNKHroks8wWVyaSXupeY4125LQ03qg7vkt4hB5FJtYCbi6ltZW
2usuqIDsbftfKw2gksCj2Y3syH3Ro13ES7YpwqcDlvc0n1ohbb1vNtIpHXNLZQ47Sm259/rkd9gu
J+mG4/mizD1yr6a94fetJFWk/Zd9F2jhiN22A/UWJLnTXuo5DYsIi4ztM/I0UnMEWLsDwNijIsq2
S0oeaYGoXryrs0UFQmturJya/LSZmDfw04A/HOSD69Rc/zPynG/nd+/iYFwnsJVGWW17SXh0echO
1sXKH95uoAlaf/iMaRYcNbiUx+WqYq8BfWMkceOzjYGjuW8nCVKcuizLPm6kez2aeEBO99pjVZ6e
ZGFr5uujUKNTP9KRA7qXfhAhakdH/5GPd7PsF5SPS8ESKoyieENIMkpxRm9cO5MuT1gsmkSGqXLC
Yp2plqm/p1TaP1CPy07oAcKnjw3S8YOxlnRKyOXL4SrTBvM6EO9qEKa0mA/tqGxIpBmWGjGPhedX
owCfoCbdCVcyXjASCyz1DFWNv9VCn4lExFMWSlG7RzATcIvlQfhQvei99+PAiMjYz2iJEkbKKSCu
7LMzvGpb6VSDk+2cDoCBYnHIOLmRZ1fxeVS6SDooK+plTR/G3IPw511fEP0b07Gb4JmwCwbjTQjS
tHb3BMuq1EFdRZGrLP/zqsnU3df2+jlLntUIgUhhK7oAXH+7T3MIKwfQCEpLb34Gu7AC+8GqQcHY
6R4Ues/1YSpaV4/VCVBLDBkSpXjjvbr2rgtE1dsdpDBlh5EjK83V4CH50nCobIaEm3tiPLz92PJg
hEd0+67MCl8PL+74IjQpQonsk1L+6H0sdv+89Ob/gHA36v9vju+M17ELSCml2EeNgq+l4wvIGQdI
2LfyR94HC0j8ck2VdL4A+R+Hg9R0/WG5VJ6LOPCOz7Deg8zSpfqeCGnM8fhh9Lvqvmwi8UO8Xo98
eGKmBqvsmEKuinDvUMZ+kcdEqgxDidfJAbdjRz7fwxhK81OyK2AKyW1Ssoe4a5j7zSikpN1iYcn0
BSBc+/iXxJzd+hDew7EHKDHqVV8gwCZyRuWjbT0V8l0NkQ8rcBjhfVnFysACo4pGPStWI1iH7bvy
YYEnwspuPLE6DWdKMFi3JhU5zmOMdlsRGv58t7ENMCiTua1jm47Q88wmHiQWUeN+mh2QruFN/tuK
Dpu4g/meUmASw2RjmAIfboMA/GlThuRaV8FZJ4Eq8sk9z7WFBVfK7rDYqohHBfGPrEfZJmQZo/kW
VBTvOL8L/DekyoTxaxVA0e+QlL3B5amN0IdsECdPgLb9vcEu+FSt7ZSGfhAz0Pj9WLThviY8pC/a
5s8McOIgbiELCqzlE6sLdj3yCIAV5aXB63ufV7z6SrgEph/hhrB+kiEkq1x6oQDMLbFNq5OA3VSO
91M5Ljs5xmvQIRucMU3cBmTodG10KTcknsLhtN3A33GMT7hFvOzYiZTKMmzoj9wX45P3aReGqopy
zL9cfgAZLGrKlJXctY7AM8ClDXEpvZNQA3pXrYcRnND+0T0Pxk12CyUo4S3shptFaqq9BiwKlGsm
JtgZpcctBCmnh0Ami6LrnE2jGfcnXCc2Y4mbF9sxnYha684spz1oWlPh7OcfiLV6SdnRSNmKmO7G
G7+Q6wavdDwyCFJeOAr0KTmSvd6fX520BjUSZPui90qXrNxtQCjtUnpGpwqEEskrqhTavttnH8wZ
uCp+SFcFx7nhO7Qan2XFy0q2loqbVMEyodojJ0KmTPRMl8OPBUVwcCkzgJs29Nzl07k6ehIHIFJW
zCeBvh/6+1ITi6Fs/bOdSIuOficfp7WaTguHm+gcmMvh6vJk0MfMhpcsptkNpAFmh8QbU4O4f2bk
eZEK/5RviWAWaXB4kPi4AfgBu1u53oR8IH4wrWimp658Bm2LCOIyIkgGzOAuuEPH51yYyt4r4SQs
ZlL/UPtpdlCGBqbtn6HFvI29Nk/A4VKaWlDEbrpg6o23bnBhn+e7r4n562Zh7qCRsIJCc7VJDUWE
kD3IloxOaHCWVDG+1ZT6lSybUiQh80SkBeGE+jaWtFjJWhms4O82/KLaW3cESc82OksjTCT/JcKC
myZd1EewqgTFRgzSbbAeftYRSsNl/gZecbAXdRnXc82C1icMHL8FuI3gwz8/DkhzkgsWcWe8IRGK
iLMOq3KJ0aRQlPamsEOYA1LaGHsxyDuhSNpKKH2uhfQhcQbg8/ZWr/I0iZDhIQn/F4h6bVDIczjD
ltqoX/Su4Y9U3sy7nnaXSHBggJcLxFHLdYP6ikqLwEiy3JJXzGLTgRWbLyPzaaJpj/IIa+OxrolA
jYy7JPUl9gClv7Xc/V3kNMn4uwLbE7BgpccZEbagSjwPgd143ijGNXnYB+mVWmGfnOgBpBgtj90G
XGiS4hh3mkIATqI/1oZM/XirzYasoYLaj0Vnla/7p+c7jZydn/un7CYhlYt7X5+zW63BSBVFOzcB
X4Uxwp56Z0A9PquZXLDUT4CbWY+m5qss0C5qTVGoRl+E/dedNIg608KOU8j8qw4bl0SxvtI4w841
MwyUSf4TWSJyvr+Qm54YIsTG/gvgsZHNTkV0c8ieaxSnFHQFZ14zsayvVpB7e32bwJBA14MX4WUq
xsCsh47FQjJsIkl0oMaZn38L5Q14KxUtHSyJ9iC/DR9iA51qX35T0c4PMsZkGbGCtMs+1UgHc1vF
8/XWV1UOEYvnJlE4gwM59N91unpybCvBDBtdk6fgRxgE0XjATGLYsmry0ncZcnJ/vLrKA5el98ui
1HtnnJAJg23Lpz5JWn94rJ561a0dm0uMDjTwuzkkkFyMc994DbIzLxmdpbtYZXk0paEqF0bVSO1h
RfPWNORhruhwK+hN4wJrWP6NQH6RBomvq+Jntmrxj1bPQ1b8sIieCw+mNB/2WbEeoFIKimQfr1mR
Sn6bZDbpeb4p0n9XSSHg6f0FHQJ0UXDvNXGpzpL0DKBQ6tnKsgRJOhX0F61Jbpd4XI0RBZ2EjJVT
wm6uW3AeYi2j3rxYdc0xCVS5dMvW7SK0hUXvdvClCSv1h4KCRfbrBH7VuvRm7N2yOJonO8jIcBf2
WHz82eOYYrSlzMrqqX2tJu02ujlUelqAY1w47CyUK8ecsNuqFFkHazRoUgUDPmxH69ZCsnH2oFsG
e0IhzemDj+TrP9a8t+/vLEDf6O6PTfVXNMLSul3pgfMBK4P3TZloSoiy/ntgpBLjlSYGiy8p+6sN
g78lVoWibm4uj5mKq6C24xH30iDVPHYn0xtV3tC0qZ1hW28e/+/l9UPvoY0m6JELY+Z5m29FgQlL
vShXLL/w7oDE8tKAf2FY7qO+xRgq/YyOtSC15uh6k4Ow3j8Ec5tD9b8WzhmHw0vKMkplxNp1RZHx
pFJK5j3FE9PSJ6zr+Qt6Y3eJMTwZ0nJGuufhSw0JQU80TMkHYP86iWhez06Rj8PCw5nrMfQfCReG
zdJiQKhp+d3KAqzCCOb9kS0LrsfRD0Nmrf2LLpW1iSLLc0IlAMzG4NxAGLGnj7hE7jdnrn4WdJfQ
6Wx/79Hy9GtBnrfaIOGxxxa0lkY62iKCneWSk36LwVGoG/a72VG3QQ8xzwggcHITobjlr9NEX0aU
3KkmWt2BREl2gOaG0zUNk9nbv9u7geEWujioCGwWylJGacgam02ik16EulK6T8pW53deilbehOXk
0SO3dLK29JPdUNiQUybzwRf9EZFccaWrxA5+VjDlzTzDZvFGWsY0GnVAFRP6CI4pX1JLTeGa3efj
DLQPh41AW9gPliRX0gBkdFf9HfFeStmdBs5PeoVERyP7PK1MWkuLtuO8D0K9tecex5L5SCFrR4dt
CLU7GwTzO0BkdVkdwgovelOL9YYHzedH3EkildMjpds3eYUlgtnl9pPLARb2xv2N0aM1pds/VrM5
P/UhauvnTZiZmaNqrCWbcqOcX//sTLuTjIHSSD/SHvF2rjie2oWM9UH626VoSWnK+uPq6gqC0AaN
q9VkfmA/1teuLiDzVYOTWvvkIQdj7s42GHHEm/NNNEeLhOW1w2Y8203TT809GNL2KZdjVIC5AsOu
bNzwH1SesCu3ex2uALpN1+ZYE5xyR3uYVI9AiqCJ4rxze9CJjJIfVtn++lVkHU8+BpvFuG11avy5
E9JqqRiACx6AvaBAmuKf+9GbGyZ+8mJTnRZ6fNvoDjGdzzEx8g5YhXqUKQsrF2S38fIxoh1s9U27
0D073NRH0/b3QLBmv7XEMqywY8WKYTZ+r7JcVh6Rc0r/AbJtlL31PiBYMtiA6Xwdnk49pIU9QGeF
ybjj2hbQFSPFzzGa1px+bs71Sri0s+o4TZO+DoP8zewEgmu6V5N6U7SJQZq8957X8TfmcHJVue2V
09FB12HYE9HrquXxQByYH/HcNvQxhc6hV6Q9s5BcuNSZ3u/CE/vAB0Rno3RjKa6bFQvROwgzCgNF
RWUaOloH/OObrTEYF0bSmGBf7cKdiAGsV832TlUxiKShu62+Puzo2U9JVl5dpHqznO+7BPHMekp1
5SHFyLBih0DqO2B95FBZLf2rYLN38FBkStpNXV6eoa9H5X0cLYiby+/jGlhqB/nYYSxwy4SJ1x9H
D4QMDvapLoMqdYR2URJSWpmAIbQ+Px1Pa6PCsnlaiBcmMrUHemxs+7eTkEJdQ9a1wPXLYU16OYcN
Uw5XDXaRGV39bLv/BvyZ/hsrfLlKt+bFizHpZ1hXRbK0bNkemPMu84d9mxfwyG/kTWHpvE554G8m
LQ49iC9uNzgkVTo39y0pqXzCsbtVUj5Z5+w980fOq4f4fyBb26Cpzd5t1+DVzdVRPAz8EN02YCDk
JPgNoOedsH3B7zIPXJIGxzQ0XtfeZX09ZpQKGDOkfYroLd7KvA/W59JQODQt1I/lPYIMPlPNbTvY
L6ML3jYgfFRF3vhE4WkDTslq6MjtCj3xSN5nNTHNeKGB5lxLGlYaK8lRS91QT59/1BBdEVzw8/yd
msVjEhV5xkRublqBbN/HowVHmUmW5SCvZjHxNPvlqAkbbG8euaUzko2XsQGCslF1tu/C2GW6q3BW
62v5jyolitM5mrg7/DoUTKu8WMvEx4bl4F3Uz29GkRKPaXhSxbyN8DS3OgOrOA6Q2hck9KDbuAw2
3/bROGifc6S+7fJ2blV7yMpwFcu9phk7ENd8HzjU+JfLrX4dwWe2ci+BRxAXewlpahM+ufPTrNJT
KldYPwjVxOHqTmGiHIJF1YTPVY/ZL3GUrdl5GOgJrbOX9aGn8XzMxtf6sXfI9HtiGtJOjbmCTnQu
OHYWEn+iHUhR9bhaul2ZtwzrIfefiKJcfDDUaa0S7EI7PIj7pFi/VSsmq5fidxmbIAYvhd/Mdu1h
DZ7KILA+JYDO45PtIN7bM7t3FuMDXMayb/iNMNyfq1t4Hf9kaAt4k6hpOjq9MPQVj4U8gyX6O3oY
pTdIQV6pw0uixGftJMKJDG1SWWO15S6UYECvvgOPuTCm/y5r0o3ToXouaNcfcJBKafMw/JK4oku+
e7qEt011iQeWTD2tvQ0NqxA6G1K2Qt3z7jRN0KvzTnSyfFAvjaL+9aZPERLbnbk/GS1vIGbMu79f
9j445N16dece32uMctLw4g/to3/yBzgXm1YPdRrOGMvTF5361VtqjNKoy/UcRxJCCBwJaxd017yO
wOeohcIe744ymKP69guWJmKKlVnRG+tk+1VP+lE0b5ICFqqMWC1Nj6JeDU7LQzNCVM6oy1x7XSQD
nXuRbxqa7ZdfCQTm4qVt57Ty5drsffh8jIdh0Lh3S01UHuELSD6VdCYji5yxYLuMni+u7gCMrdhc
fCTveCItkUmkqG62gOZp0ohz6q5OuNwqg2v1WRIOoiDRlMngz2I9fFVXOn7HHzdn+jZ+TRSKmrEO
TkprrzWLkynF9OC95CvbUcyir6Lxiq3kx2FVEqNK0RpHuJ7xXgseLqj+8kOKsDDXg6OlmRqjuVxF
d+HPuSBs74EDoFrV5xbUCZKHtcFGSNmWbmK4HrwxaLtUzrcxmTfv0b3Z7qSFz9TjMfDqoPFa03BT
q4+qwv5GJouzzTFPXXgEwjiajwhBYtncsI8xIGh1xf3ZIq0+BFSK38FN5f5rme0bkX6dU0c8SjEe
6/6vU5jrGNYc/nDtQhEDfzf4CNDuewz5olhg0bAphLXpr3Sm6nRKtH84SaBqmJY7JuFx3ECTJCqE
UZdu0YxOBQ3lVuNbwn7Y1UyeoOuf3ddGxcWc+8eyQ1ACS0dYFZVRbw7cBYCR+Vj2QDoPGBTD/p1q
vm14FRPLlZsVfvrcQ5bq2h6pKlsKdS4rVO+yQawIWGtgl2Ua6bWE6N7rOtiTIwKs+aTKCvfgqsf2
Ns36lxgcfCo6WxW2j9nvL60dlZfhgYkT9JbzwaC5VgvnRq6ImEokue1N7hXYnLW/mJxC2lm+rTiF
53vZ0WvirtO1I4hWJ9Y4+9pn1vckH6pVHhkxijqpxz8EqrhSLnABaywnLOALbKbZtrF1H1wgaFAp
XWyRlpidpi2OuzPFTnTC6JDwILzmmcYpHNxahFsfir81rJzM4XyE5QN2IhpPkoj44cvi79mXOCPt
HkGLH19h6x0mxqnrEOpgIrWWQswC9qrLX5kFTTwn6OOhJbphaqx9jkB2aRKw6S0JQwCerW6p9Jhz
bgfhyax/HRySV5i9zDZJZNENClsxIQXAM5g2uZI6lzcLi3s60yHpxDqIWSy8INPSuBOl4iwrwqsB
64IAiHKxJkSTuvxMlvn6OUhqR2XhewHTTBJT6Wk14lD+FKiOj8BuOEuI+HTxAFgyvjFSvTkWT04U
neo/GhVI8BVlLrNo3EscROXYQCsAWNhj1QJiVOTmV9VKhCm3LKsWsbji9PdBl94W2cYnoWfavOVJ
QDRO0eM4hqkrU4DN4HFJuWmg6FLAOEI7RkobJELsqeX1F68rX29mIQgfa1r1CgmdoAGuzvGTwmmK
DdPmg4UB4PAFLQfNOC+LIc7Fr0d5ft7/HWqErQthziBRJGtb0KkzVz4GHmUmJQuXPB1hTHjS4v3E
U0R/icJEa8bg4TZRHKnYgrjrRN/NZD1c5Kbc136JrYD3ERt9pqAhSbBqSsjeDmQXkSaNTXh95uus
J5P0X/WV1VN77lZFMAy21agIApnKLCmz1en6m7ty9G8ytfGt1ozfLtju49FxwycWYwDMxWSxBS+K
V4WveVFU9tRQ+SSoX1VcKBQnEQ55rYDHACSugTnj2mg+WmtzBnDab4T8NzQthRWB3tQHgXs+Qcic
bE4Zdl7DJgTvv/ATWck0i8H37QIXgc6DXIGCZmhdP2HkZtxA8N4IaZPyRpjlDQO+KGZP0/WYvOEo
76J9UxjS6UEvQ6hT3FDqrTX039pxlhOb1Iw+x4LjBwO3hA/7nKs3HVvUcSs+iQq7zv+MI/M/azAi
j35CiyWg5dbYS1PrwwgWL8+JeYLnkHJ/TPhtJ4gHBc/163VaWM8L8z2LyKuDQ1tL8Vs3Duwbopif
/n3phc/vYXHrBB5j8ntismiX4nD1Ih7gwBQvslNZWp3mvg8sR3YdLuAvEpWwAiD0C+tosqlFk/6A
asUc+tDAW0+zAn3nQA4nMKephJQR1NMkxc6qjZDlnZUMfmm103jkRIwxcH4L9SUNVM6V8pWhrObA
fNbtmtV3IK1BI0htEp7k8qoXvUz2deNUHt+oPyhYlUPZ2hNrYXbk9eHYv84ASzl3dalPFx/U02eT
t8VjdYe1wHI+7Z0iJ1YaqYFjQaC9HE4/5RVHs/6SInYq5IF2T14wXjX3apKblEZ2KNDDg1ti4gEm
CzqeoheW5STljTaeEx7/A4XbsuN5QKoMhNgpB612JhZTNnSKOa5wQ2mxto9EEYqfp/HBagMBcBnd
SyEYksoJJN/xEjNpwRBKi3oEJXJ534DGjbVIy7nX66ywzZZwCqDoKBYN9sU5cEuIT00HkI5FpczR
zM52WcNRHw2B6FlLcMkZTqPAc6jWHBJJ73Tnl76d3n/qoEiGNqFq12kvrI4pu/dZ6XyYGlpge56A
IsVFRRHE07FM4EhDYfrLz/TWIkd1J9Yyor2sl59Be8wtWn9Xtk2gqjbBDP4FvYQgyidjTbjMvCCe
f5jRH3Gokc1nCx6xLFBGPzJkUbrBP1NeMvOTy50LLIqQCBmdNZKb/OL9ebCZzAUXe+fMCTB9Msi+
4xyYamuoR3glItYJDt7Y6nozJSuV8fzpuMw6fzMsMHnMOQaiNI9bT8EkPd0HwuU8RlknHoaGebx3
RKnCH7o9p9ELn8km/+LFJTVwtwflElMrROwNjkXrUv4ZmgPfE8EYTEzMnYzJFbKyLWaKbSBwmmja
lyYFx7lLEnu2pvBfP7PKP5lrb0b5STk5UMYUlyrEfaJBS2Ba17q4qJsN1zliw8WMaBG4+5W8bL8l
/Rbg+2znHeQoXbcU2jyRGVDGZYEtpFCaoyVXKfVQRYSOSUnQvto7floF4LodvEw+iB6mQ4/r/BN6
DWFzgBoZ20XLDTdrNpPAuLjThyfKNYF/XudlbnR+hpVL99sSgug3vRlGBeUwJLpTmwtiiopheeQU
17apZUOx53e2WSWOb6wcodp62fyEzgRn4wGkT7dA/bjcichwTen4wKF1TjhjhpOpoyZiU/y3Sh9A
8ZTEVu0jnEXdmGxJqx/bwhUdUF7LrhRL1/HuJB2SbZM/U7V7Ze/6d0+4hH9fe/YMg0YQNuFWKbAY
kVC6c4jQxr1bohiSySUHxNqLvgjcyXsepzeBYsAvux7GHLVs7TKPNo9o6owxwcQU1fA1hzAGpkWa
8JKoZPSZ4xlyjpxPivV5imxSrK1MP0pAET21YfAKxaOvTp0OaebRuDptwBSaD+QQxW9qJx8bYmFl
04JE05dGmLrXwHDiax1N9l2xOiqOJ3XJi/hNvlrKZrR30WZrNb81ydN/U/Asg0aR2NSIo6SBVEmQ
gnqUizlVOseg7h90GgorCBJRFynCUcQDWoCTaknrc2TQKmT4oBqGoJ3o8gTB+v3qv6DRjPDR00SH
DqmJZ0A5RFJ7llqJj+4jrS3usLryfj0IxEpFq1lNoxjZaOLO1+DA9uLjqiduKGm92IoHg7yvoitz
wLlTJq1ydg5aNT14bTe+WwAYYUFqAEGCiJKOdWi6GoGgEGLG8EjGauo048NXkJqfAGDH9oLC3nHl
tQoerR8PdTrHYrzNb1tldMxEKrVfq9K2SXFm2jLBsdMiCN4dVhQzd+GRfglg8jZkqQQYLdbfOvLB
xW2JF06aUEmDNQr61e9aBGxZWLn3sCv1fnSiOjYmeS16+FBSr6kTnm7ydTSJET74hjCVrygwcrrO
tIVYcOsjZzDWEwyMLFQL7oN77Ptt7XebGez/aZl4rJPbU6YCnYXl4ByDtwuhcHRqcQIJlpf8LSxk
IUzuRjwZcP88iuRwYaHZmFAJvMFNSMSZuPNC4IX89/EtID1e406eRE0sANRw0+XjipB9+ZirJVgE
cksl9d3dA0JX7WNHCRy7DWdtc/wOOzTC9iZ7GI9ylzNveFp0HAiA6d9wUh4u16PmYVtf+q7purdx
nRnKDjKAcBYGr09PZV+165GCcMyJQmK8aN15iWAzmqaqSJ6SjfzjtC/QcfnGbYeYI2wEmClXMnI0
f7EYZmKbv/sNz7s+iG6emYu6XsAR40CPbczsQPu3/6SWeeWvdPtw/Q/IZCO0iw0oMlFeFk1GQjFH
R+vbf2V9AaQ1/O3kOVYEWy0JzHEOPRUaxek4EIKI8hnf+Hh8ErN0EeUtaDPNrKWY+tDH8H6Qh/Vs
WYw/dKTO4Kx+x+6Nq6AjI9rjslzrPJtU4yYhXTcHEZdA4khWQXX7tiz9gSouNAioBizOYn6mPiQA
HCvk3FTpTNOhIvxSaDY5rlANwGNZfmJl9YziNR0yvmUrAmrMHJhUFjz2Itw7p6MlE0LTOdjVBHgq
9/WgzZdgYxyYHc2WDFptqC4ocCrEpwAo96boLKlXHufAAeTT/VLj9Z2lYapITOC1IKVaZHyf5PMJ
FGHnKcf8sPM+k7y/pSQtZboOvigdj3dAKgJKaNLRN/bGoD+RPFpPEHzU4BOxViEBTg1oGJpIWzSw
ovJc+zZpJGj12DJeTGFdJ8OE//SM79czRsIPqOElYrdAPG+tENvoVslaWsvZX5rXExf88u4TMqqt
jv9m2rjG2JY627ScgT6ppXqn/tzLE1DGnGQ9GbsqLbeXOX270ISTnhkUutWRgbNZj++anwV4/43G
KUDcGb/++Z9j8iE/Ngz49PjfxQ2h0cmkJi1Z1dnH3WpvCOLCXw7VdfaLawYzZGN0h7YzSFcY+yH5
aybzlLadtVX1g1y5RGSsPUJon6Awulynl8DAADdKVTLgrnRG4azxho6n4cdvvTxXsbrGg16ygPp9
fz0RLa0K6EW7nwZTmSXXelQViqKqyWKp1DUAJkFGbmpxo7K1K5SdlaZmDPax9v1ide0jDWDh156I
Fejf4mBBkP57af5JhrxUhynrIIyGXeXGrG7jBxgGj4H0EYC57KSqp7T+OAqJ5tj+mZFiJyBhApr4
8cIvNToOvgr4te92zajG9sDll+yvGJYr1rAHYN4bFmKtGFALJOrTBbZRFI72VesoXX0G7ez82y5R
sIfh41CrR5lxM/OBoL/NbSjXLvDsNLVB214npdsqHYvBbMcB7paByyxv2l2oIPa2KN4lUSfI/3P8
yC02kHTEMKSvSSZHf+Xp/BUtKtb8PjFtg8f3jhltq4O4mKHvEtRbnwVZfBpL+7jgxyUzbXWzha6g
1HXtpXJY7sxYmDmuktkvnKOioEJ0tI6A3/3b2XSLXSnzZXAjZFtUryHd5Ai4lBMz1KCE6aOUTNGj
GIfUSnThM5laU6C9zzIsD3KVLzLUO4v0Q9XN2VOGHg9+wdkOLXtMwXl31wOWkKKUOqvMblWwlWVM
7eKSM84coO10Z+QJuIHi/jBq7YaINCFpYa40vhxgR1Gwpu7B6/4nnPxJtdHnu5FlqjlsVNju+bvn
4OWlF3vU6AIpSg0nrp6dq8S1hfEgqsKazIzF97ZikpSb57eT0Pbj6GMny1mI+y4mPMl0Vm17FkWD
AqghFSYtcnfjLzNqUZt0Pf3WzkDDBUQDAIJzh6E3eMVCb4Vxwu4WxbuSzdNcpzYiNQG0Uem2RrpW
5Dl2ZnfulmRCNqjQ/grSNPNqWQn4CIzNMBzaXKG20vKVi5xTvdiCc3fRGRsFpjUypp8B6trW/f0X
x+mWRyDH8hSNrlqRJHOx/ztiS/We6LxcD+KY9m1GGeLmRUkOPCTP/nkuR/cXvaW/prp0Fs9HYtmK
ke4PHFXad3jMt+dj6Dno+m8qWSvRCHsWjiS+3TxBeWnGnQuNgkRAqto1H7A3VxNzQ1/VzI5kJSUs
l78/ipl7bRldfjpbfrfGNB77zrqshwg4cZVOkBmu4/cwY0rArQqf41ssCkEMh5M0946OJyQQfFEW
7cWvs623DVrCRbFBCtwjWRi8W6gxwSDZw4w7ODD6f7mTJPLhXls//URAyEBn6xJ1ZHGd483ARPEe
Tpm++y+quV3M6Zs+CufHY3cjtzAeGdp2lWk2H7pdf7sK9nirhrnbfw9DuUiNtFIz4arTqWILjMsc
rcFoZkfvzgr/uqV+Vv32YpOBdioML6qoWiIpTuAuFy9AW4djd8CwWZiulzqIzCSDbBGR1zwkz7os
ggB825JmNbUQMTNLb81NvFCkqKf1/QwKYZxs1L1hG/U7YMCVQlJZV8Capfozw0MiOSEFK73t7hcy
gQoUKUFmGlGmohBjArk2G7iv2dYZLgmKiXk6jbhR3fV+rCha8tlU9tUHutwEL9/uygby+mX0fT7D
p0U2ocdkwwsvK1M5wahMtEAvWn8HydgPD5i38k9CXfOh1FnYc6BM3sHObA+EkERQZFl57EOBmIsD
bQFqVqee90uDjYYGdnjD7+PqiKINo2wN8nwsPO54qPIYCptfOA2ODqReWifhu9PxQDvi7ThwYhbm
tNk0HvUJ8x2jQfuh50df6FUczky8GPNEmA1yZKhcgBNWD9nMN3v4VJ6fTNMkWhtfA8etf7zMD6bV
BMf55aQ/ElF6wZkRkOnman+IT+k0Na4Xx5fwxlCmoXpYZIlDvuSO6kHq22hAZn4JxcPcls+NrFXk
5ifF3zpBq+kPZCnqXcLPQ9/5zGCC33h33RsMqCdde9uPNIrHcS9MAAWNtGXWD4VXyizt37j3dDMj
PHqknjC6hTdOxT6TtvbM5wcxg8Dd4WfcliqzAETQGzyKfR+vYPLkgaJ9yPhYWg4sxpVmJ6XW+y2f
JHOaOnJ+JLU3aF48dEQkup6LPkzndFllNJme2+X1GhQNKNDbI42qT6qnc5v/+brcJrDvLd6k7jcV
XdsqMlheC41KBZ5bX8AeZe5ZLh/qiaSo2hVdauxEzHxy7tFb8/LN/4UFEOoYWi0dRw0wcvukGhOQ
96WrQJDQuN57UUEwGzMJrdJjjRE6lxBQFhV0m8ljbd43RzHHJdrcVaXIcadH4rnfFI0CpNmUQ4zC
VA2DiiKQ2/v/YNk2iIfdnpz3n5srZbLqaGbfyNkqo6SZj/MkHjSpSVf3/w7hAjh0lAaPtaKgCW4z
Co6Vvx0U87IQlC3NP94d4hnhtYDYDC2AZWkPIsGODnkDe8xjD90JOzIOkzxy2bmtxx/ntF6lJ94u
y2g+ERDSSjTDEuYH5iG/wJ/otXL2I0cO1xI35mSL+lxmBXj5ZZc0jyztiSw8OPHPy3fo2oKl+X5g
Y4sG6RQGtLUDmxFT0EFThZIk+SpQwUJtY1b6CnL3QkCzV+aOulFkMpFqcmcKbXQpzsUZUh9iLZMW
1mWoVpTWVMfnOrdAI42K4TdIPuXdtK8jpgvTgc8aO/M87t6UnMx07ngoXd1a5bNhIVY+SUA/nhht
Iw1lpfW0gR5YIGTHsm9dvTTZeRYEcYi6IvSJeESWNr8ojHHMhRyMoja6QW++F3i8imuUF/5BuHBH
alzx7Uj8p2JIRDYB5xwrJUELXIJkZIURNWKCpvqdP+dfGAxizmUHboTgbmdrAAhmvcveT5kcrbbm
hDHV8lxpfTtsTlHhxyozqX+zJ+1fln7jhRIqA5jOurytJy+3j+Nu0rBYe2NnGtUy91Vfh7nkG14b
pXCsihs+AdOnRha3EJ4qZFq5Yb/6eP4T5zutchW+NLU27JttU9uA8s8B24YhWDpAnWlKlJQD9pvt
G4dzKFFf5hcIGg6f3I7UQnqpCWA965Ub/MIvoYm3gwTKTPuhH7GurGnpNqutwViKmoKZgF2almtL
JEP2jBmy4u0NtPOKRNIFv+DnXpDAA5iuHApGLEgfLziWUBMUWbF/wAiuiQTMllQV2cjBiaZQ8M1J
SXbBGjXpKtd8n1DQNSo4Fw9nikH+Vn8vR6toDcX7GP8CVKEikgbskzc3hd83gMC+O/76u5GhqPe5
vpuMH0w6ryC0gQbhty6m0QS1udtSDWDFO7E1C9ijrIz+F4TNY4ah5pQWLBi4yrnSDG6hoGnRj0c/
OfbLtGYWAe+qd4+hkAAQRMlg+SouhxOrERYn64m11Ht41eLmBeHcovjhutmLFeFF8dZ1krD7787n
+Pmzh3172FcWBkSEJL6ZbFyBgAQhACVsLrIrhLM2Yu/qgLObZyGjt1KlFqSg1WmA28WJvnc89ynW
G6Izcg9tsEhU7ichiILGuLDCxakmFRtMz+/Jp/I8Z4fgyyBqTsXzC9akYVqWq/xv1IHXR8k4Mq91
S0K8kIsk8Cgj+DV1g+8DfsWXF8WkNedvjKYcbsZCegnRD/SX7qIbIf1Zt4NHMuf2XLaLM6hCxqu6
61EbiTXMf7OEk+GAXemFsm6cG2DSVZcqudQlB6Riud1jaFnV+cxYcIY8rt6xIXor4X0iXRAMn0yg
Nc6Mr6GNBOnJP8+7KkaN7SdjrYVjbOMY9ZsylL2zfEN2TsTHmeGslu2/1K/1yYZ0bZIRDSYC/jK1
lII0VvEf15E8YGinYc++QtQJIA0bGB3g8PuJwa87OepE4qC48m+zZqkgChuEPeXNLIcQmPsIW5fw
DsgiFqM6eZ272daTcstqLtlP7wVWZXE74IaDPMLeRlGpL2yTRvb8yaZ3Ci6B6pYzColXKgN/gsCG
PT6OOM04sngtUjKPreLBCVbXPcdw1RJNcQX6BW0YbHIQDraeqN4SlDQXfY261+TiSJ40GG7t0tf2
ZWRa2IkXWTlRQN5234S+c3qXRNpL4LSxtR00dy8FcdCPWy7QPD+Tszr6Za1D3uivoblv5z6jx5qB
5D0t+/wdsLRQ5ox/qrZ0IQxBacxBmnjAKOKow9LvDEbJX0ht1/jGTBDINniVxRxib7SkAF5e8EPo
niS9oo2W2EHqm+BveroEXX5L3a3PAPwnJrah64fAe5g7hjGYz3c0fKisfXW/L/uHbVcc8KznV6ZY
LkRrP9+c1CDUV2tT0VNOrQFT786+HFg/3BxA3z76DF2irvhGlTpYE/fgoul/4DQlOQ+GwYb0VOaL
TEEuKIjtbfHNn2cvgqxj1y/KwIH3u9ZAUNrLleYftaZhLG9WMfS/7UjABwV+aDiQW3D6mcaQEvHE
JHfSI52Z4bmo4NShZku/KE5Nb9vfOq36v+gBR6E43ca27Nr71iz6CH+afrYzPS7XSaBHFncuZA8u
6F50f7+rawt1oCFxpXh0XQa0HOrC6LWJPV6kia3C/8jn3s1rp+xeTMroDvnO0+MnGFgl4gwp7vSx
F10jYZi0vvN3ksmAlEpNb+U8ZvnOFJiekNIfX4rnSAd6s/YtL8jI5q1Nhgt5w5hTDm7e9M2u1kDX
ycPAhvNBGgU2HC7SQ730cy7TKSmPkgPLovh7p+alLT5X558tOByw6N+FIfRO41y0DuH5nzBbVvpf
xTshs/YjxiY8UGhCFhe/6Lr6SyGW1E5ScakDpGg23kRT9oCKLe+JtqFLA6DEhl9ELghkBSMu+pJw
alNmUUYqgltmN0zv/vPVfUl7BAvq/TBWJYjQQIECZ8XoMAnM2zHd6aOB01QHjZtFlEnx2pKMoA6C
Kwt90DAJqkTYgIfYao7yOmuvBiim5yssSpff0nKWtzYU7AS+3aR25/cEQeT4XpPNQBGSAPGLj1vZ
KFzordY7nGTCR/I5njO0GdV5zEPM8QBbbpOfmo19rHmo5Uyv7sT7pEVlwav0IPax90a2qSsWw9PS
fH9vYS92UoEOtfOkH9kfV5taXe+/21hqheZ/vkXAQIbqdtFLacVELoeQlNXJdh6UmxaxLqWbDg6G
7mr6s7qJDRjaKYZk1SKSbkMiAM/e4QCLeceFig2/57nwklayV+1WpIYqI/9EPew8k5leXbJWVJoS
ZfYi/R7G0ugRfhTsoG1T1CbR0l3dBFmET/v2OGFF+DJc33cMAAeA06HdgmVkG0ngd12MRslvWX46
n6cEQ9C1+OxU73NLbLaaJe7/IWGkwqdbzydrXbEoYoLDTbUUrQNuU2LzSo9u8S45k902bsHjXekZ
2O26pc6+pXJ1EVWkIvaBaZiMqOUKeQJqMDsbKpwsZef32/QsovwwOINCjBUtBSqz/CO0RaoD2aaC
55FnSSti5IZKG3tNV46s/DrLXklFPWeD+l7dipHwPBrE8oB/O3wm5gs0wvYy9plg5xSRe4vezjuS
LRQ3FoWSNiWpHz2E/wE0wXAN/gHe7sWDRLZFKIiRM4ecXbQ/nWVQezSHBtjNGZU6FVk0ZtYtKIyG
ARJXJ1DJ87fnRMjrt11Y8OdzUxWnkA85hy4UIfNtloJfoizIS3FYid0xYT9pF9jd7Yk2JjrF9W/U
DPZOhUxvyXbFuJwRTg8VfmWu9cAfkBs3tveabsqX3Uz5rMKXoY2d/QKD3+nM+dr7EnXMQXq4Moq+
A4ylCeAvNAsl92AxlclD1QMM824DiyNXjC8dCF6YFc8g+5P/FBIMxDFXFvEc+v8q/8D1PrZ+Dn7d
wi0I5xh5JCYIT+MAUPq1q8NettvTgkRcDMHcL88yV3K7XrMrayp/I9Y3/98JGkKWDwjAXRjHhQCw
eH/ii5YZSd13ZiMLos6I1kqb78krRADYWOdg8qRlnfaowp0s+R/zVzNKdSWcAPzvBIotZUkm3yyh
en5nIMjq/C4lfSz55nQtNTTH6bnKrGTZf+SWw81BNgA2m+nvbnb/Clbb8HlPlpby4yzeR+YfiIWG
An/7IkxvBi/c7mDNKkuduNFVdYxO1bhi0JMU3gIW/MFqD5sgHHBN/DM48QZ+jNJSbVn+ZuUbj+Wh
qR5i/cbds1/9vXtFZuMzwK+2fdCK7raHbQyiaHX/7uL5Wu4oiIKUf48XhnHn9VvkV40mTnw/GG3b
ZjFJXU52Cu7Q4L0hn6963RLLC+M9x0f+jKI8M7myIb7qpiZlgAF9IpcB6dlt1O4qA88QylXP53Xo
td+8/dFsDu5T+6n2k240vfiZ+E3Njnp5drOmS+CWTuR5Dv/TkP6Kv7jQ5p7rfMoFWw2TWsviCzVs
HKWatCY6hgpr+PPgY+HQQxVaw7wxQB+ImzgF5Pcs4NzLWBL51hdlqT+nB3p0kH1D42NpIAo5Mqht
1oyE/clz0E1lttD6nuXYU9oZg2oI9q87osjWPHXDEQX0DMNZRx8s413bpjwwJLLe+eLW+OJSIVaH
OG0dYEkfwyEnw+gDGhXMK3QG5/7ZrAaC5JopfdFeTB9Z9MaXWcbNjbYUdMLis72USOhMCnsse7iO
5NWY86SUX/A5ppDvkCj/2aLhEZzwkfu6wueTveOnLo5Tr0BFpzUCZpetQkjWb4/swWDt3dzRtInC
rVDTwkiuVkvze7861IjplauaJQiTN0sc/ndSbi9WOhpE3K+zFyz21Ba/CbV+alDzEYwwBumvLPsE
Sp0weo5LRsBdij7IMtTHnEosJwCE5scHKOOcwGtICflDiDS13QsikOiVeUca32oubvdSSPAqw8OX
KGmtFtD0RsdWLxWhzevSXt72A2EwXOCnNiy14M+YVBcvYdJ0AtW5Q4QxGUZjP8GXrBiJ0yMpBnLi
t3cUmf/7UIShcGVrKJ7Sf70tcRGWoc0mAq6vSuNlv10B/tWPSijml15iKlt2TvnCtw70k3YsDTFS
Ubs0N//I9WP0VCSxnrGSzLLLMOpyqyXbi7LWdPjceWVrSZUGsopmAlUXKZRuDcBBv1zZTsAfHm2M
CJnqcUnjHckRTZScT7SkZ1cbbCv54gXEiIX7kw2wulK7la7OLInhZoQ+iLnznyyvKiz2Arip74Ic
I9hqU7yMcsTAN8g554VmNliVhCuEpnF9Pp+zR2L7S3oWV6qkM7+tbz+lsCEsAcZloop+WvHe/IrD
g5LpOjLCxSjpXqmmIKvhAjoxwlnFSPqqMHi5ssOaDSEv81evuKq/xJFhTu45vN7fxf3vKYywGTBp
N7yH9KhBwYPEgHgySmaP4OEyrz5V3hZLP0BY2zZDESVUc43vOSddCM1WCxGXgP+kKBOXBUlOWMvF
BUkyrCuQ+lfdpD6jkReWSdSA+qYQgxzL2udCE4i6ANhsTLn74YbpKjFCJPMgGvISCwzBIFw47lT+
hWSnUdN8c/QppPmiCd/1Nd7bv7xThA0bX7jcxfiaQWBT67OlT9fjVmf044CR+T/Jo8P76Bozu+vY
tB8blxFAfVdS+KMIZpd25xjR4xtM1eiY52eCUzbS5vEhp6o+8IdHDnoXycog0uVo9hk2IIMsT9Fj
ogatsCIe2lpsitVy45YpQ3OD5imj8oZSjky/Byd+cRDT7yjaN/LRsjwOMI08o+vp/0koAX1wY2Dj
pG3R4DkRKvwrkO3fybMT8mshmeemL2QkCnoP0lIGgk//LzIhZmFdRq/sjy3kdw4adlXCbE6uM8aS
qbTTIJBPBUyweDTM1WXJkWOZ3eBxOXn6uHejcHWwS9uTdJ6E5M7G8aMpYKvr60Utps11GRts+hUm
NiBoxK7UF5Jz5ivw8UKVO0UDJcLWJeOkcOLlz4SqEwCsRtZ4eNqpU4RhC7fDCjlGwX7fcencZL+g
Kp6jXBpgCag8Q+O0NJJDkGbubYZLAPt1O+mW8kN37a3ROiRS5P0ycYyf69AMNFye/Uv0b4AbE1wS
Iiu4XCX96Ziu6Abh+/2wMFmkqhW6T7a85PzS8mXFXpYg6idMEI74KHkgEHaTHPqnWOVQDDf8D6bu
4mlhIOtrlLxw1I88WcEfzDUmuHBcalFBXYIg6MAmVvai7+yQ8JWqcZUcbVy8mCDdZRnJF/pOXXdJ
6TdexfGdwEWYO7tR6ri/jiFo1H6tOcxRXSdJ6fZ4blmc2nedyYsHnxNIVbOuUJ9siQFseRycG74l
OAF2nO8SFShEAz+LMmaw/EoW8NCG14/Z22TkfqGScFGI2scunOhiF1LRMRnLrVaZhqHoG2/CsYt+
Yaj9RYScwE+YzZ5pJhAjZkASP3wwoTGgQAmwRj6mx+XLo2tTTZo+JZ24FiMoQaq4IKqOwlp76mtI
oxMMYqcdzwFd/b88z4pKaB8yyc0TzbjGfJjMgXALi1uZAKCOaWkf324x60iOSh21I+aH3pC8n6ri
+oj7dCSty3xItzSxd8AvKFIcfOT1Svl2zMRIoEPHRwUupj5XbptQNsJ4nUjG584WAmN7sczse7ZG
/0MxNPlpjEcZrcYrs0ohwIzcTNEaKjX2pKMY/qt2zapwUUSuI1zzHdTAxzWIx5+6y0jIBL2Ksa9W
ldYqNcrPj/pMr13RqkQ8JOB4PWYhjog3RWF7ADWjqyMxAMw5jUO6SiF52pnesV8XwcjydgAO2siu
xL7pRY81zLhDCBlIxKelT6OeUKzFgTsQORq5XyPlyCGKdYHoPdDUtv9iVj0cFN1QaUuOCIyu9+hT
BRn5IOfiZe/vWTVvf/re49QL4FiAvlCtyUuPqEW0OkGL5ePas60zF1489NXt9MAextHw0iD2TXZ8
DC7m94PMt2Co/vr6bsm7cCgu7J09108RBeq6lHHNrYV8J3Q4OVTl4m0lI98FHXIz07pIx16mkUNa
9+Ov4DSadSDMBQttMNhOeVXBC17myMsqc1DVy9zFN37iphdvPOmaY9cQM4A3rPqwvRyWdiD0bDfq
xAlElVyVVxP3X027YU+xNkJjHSlJ1AxKJaYzdy8QkBIg7qhvfgyD7dMYmc39qPYEj/d/forQOQJ5
giqocdSHQEFw8+E01s48+oF1Vq9IJ1Eu0EF2/kTFj4MxVQyy5kfg748XIhqdAXEcFSNl4eSip8WX
klyFegRXQw94SVz9DbQ1287OazIoWZgjMuk9ScEdlV/NfyJknavsCVW7OaduPqlSjnPqDbeymDOS
MDIyDphMK/SjsZO1LGthBoLhT/+mHk3hBbhZ3HdeOwB9QbjPK+2QkKWnnwQf5o6/xuvXPpgeUaN4
FWpGBc0cy9Wf3jY8NOmItCGmXRlkpuiKhGaXnfzqqfuSBjJ1KnQvOxCG7TDdMs4dugFy0Jlvwb2F
CM+MyJYnnA6euUid3fr49S8qhF4wj5xSC3gofotLQTAHsKNzhZhFs2RpNtCm0Amg6yUSpHuil2yY
f7m2MhQWq0LYodX/TT7RmbQfhjmBGZFQi4t50ZOxzHGuGXWfmvkZhpm6s7qPjiWgeawqe/cTnH6U
nDbgdBoFT/1DxOjP1KU2hJUIdfl9iaIe8XH03HYJD71slHV05jdfK+/zJrwBXh0xHfupACUFwtPq
gpzC6HCOE4NPyWfVJHnpWQ3DcNEpHXxgqnIf75Uq649MtJ+F0/Q7vHev/uxC5k6rwvx6ZXsbcRJ0
FUmstXeLFOu12WWFkioXmM8mLQK+95eeEK/RjfFBr5Momf/0uu4Aw0UL3V3yF9aYP0XvgleeV8Hy
WNr6iRpyc6r9EPz1x0zbGAMEgHGZHBMNUJjkd43Wb8AzqC713yb8uTbZVFQWrfqRtqrPR9o6KPiL
kbgPkZUjntVJwV8AwACvpULWlYm7m+QMpRQq0zxf5OM0hD+3I8Ys+nwjp0fxP8nuey7tgTsRRN1n
8k1bSH7uAUv2yZPKjuNdBHibcH4O2ieHftmBhFAdgBYjqZPYFGwBFdx6VAfvtTv3VxlwEuvb/k0m
xHDmvU7ogXARlQpIWYBt7tZMRffz6cU4OY7rs1Duet54dOKbfoDshaCGagYsu+vEn0GYJttyuSmI
oyA54TllS2yjS955HBB1j7e/1/3C0NYbn7BLyFcnC19ooLq2XY9Pb81pnI8yz0L2kjUMHNUL8fPK
r1b43vWgYymQ0VeoaoPZX7KYXgDEEsLvCPZVV1Z6oTtGGAYKzNkMAclRTkf2VA39poFdRbWT4gt+
wrE6lySN8lENWUsfXiIirVnZ/eUWwErlMu0VRQa7VP2UwSJBPyfMS1ZRtIxnf7lMVvG0Iww+ZqHl
sYhqVPNFCUENJ5RlgFn16V+2eg+BZ1ddvYVotajTQoliF3l1NknVBwbJ/Sq0O17tPNfDVAmXktwQ
a6TyCNAdSPsar1GeXgoZ2jDXuAaO3ZbPygXyzcOAWA+8lafcbd22a+YPh0pLZnYW+7QZOEZNe4fI
02kZFHUy0YGfpfr9s/4AZ3BHR+r6lld7grx5JvOAx4YVoM2169uSchVAlEJRriRlL2xkgsS+v4F0
KG0tsxfHMdCLM+TTBTaDaQ6Orxnof72wbjtQ/+FVmenZ+obe36ayw5IUxLQqtlT7O1707qM6jbKU
jtnORNO0Q+5FxBXa2qrv2xmVrNACiPCmeKYueoL96S1lDMgQqHoGSQCH7uJhr3QQd25vGFc9o9JH
HGnoolRd0/q+2APgCe5hIAl+G+EsAkaFHPC3/du4wb6XpEGSvS1CJ0rQre2GZ7zq83rhIdKbk7tx
rAknHhJh9MMnxpFvnQeFkujflHVdo9SOk7f5R9YZ1EuYJz3Sb61C1b+F1KWJxjnVh9gE1LOrKFdq
I+5DkMKGMV06GxhhvjRJi/h3WG+MrAPEhHvEVIfIcJ9q2zyoGObvXjWRi5+lbIP7F/CGYDxqUJkV
Hw0G7T297o5SW4shi+HnFdveA/d37N2w7P4d4B0zajvwTPdqSXEnhtBAprVn5tb5yK4cOFkxfP36
FYW2zSlZe0d+IGep5lpx+jZ2OyMNIxUudIhR7bjC3DdPl4kVulJKlk/xrNLnlVtNQYMUFlXO/Jzo
coRu9VbVHstU0MNb3PuiFVOVa437rOmYtQQKk42tp1Jkwl61efjyhDbi5416laPOiEC2Oh+P5joz
nRC9vIUaLWTwG7+amXS5wBQJWrBrrdV7z9LocAMiaekzm1R++AVOwGKOLN3pTDiPGJ7c5QVV8o+a
3p0FcuCcQfcjaDVSAzM/qDyTy0JIr2ixTEIGiro1d43UjsRJ/pkd2Vvw9d5XKROzEKwLT9OBlDzy
Q6dAbDNjP17M56ATW5wx0xALJ1AWwcW6Gr3bjN9tKqCQwc2dD4TFbD1WMBzoaTQdZNNvIOAG0bpW
Dk+FcHTlDSzawbFlzhgUqvMLXLGugYTmKcVFgxC6j9VowV5kLo1MfaVVyKJQWjsexl0Hzn+s5gWg
6KYFlpb1Rf4a56r4SgVd4RXK1Q7J2UyeLTnzT+4zgO1ZByMyb2FMkUhevZ8e30ND42BxODrkWRDK
awTn0ChUnSe8/REyhnKOehiJQVTpP5MTwcfOureCQOPCzoRYAyJ16q3pjWY9fcPoXLe4mOP4hEcI
KjZbeLk5Rmkoo3rwhG0yLZ6P7uWueh3tNkEJIJbyizvG541zxtysU3f1j4R35yXJjrGlk1MkV87R
1gb9rSrEDOZxA6MPiLij4ClPOA1nxwXlaUBxqHw5m3USxeIuiO0ShlbU8zFD/uxEKtA78ro4XSTm
5g1EJDlv1vG03yfTUprlCprBWcdMSVbpDAqY+HNI6em+Ympk/0EanK49MS29fY+XLfax8ODAqZB5
K7EwkOwdGt9rxwJTKELsoYpNKaH8F7bNlnI8VUAFCu2lejP9fnx6ADBnFrJANpnlrsIOA1NSy7x8
1zxPtbT5f8HzMs80s1mYcL7LntNRNTHHoamV4MOEylMU3X8lwi3zb7HDDua8hiYEt0tOe4MVMEcS
DMfEpr4eE8IvonLctkGGqk68oT9vi7smn0qr7Jl78t8pHEP4xMt2E/PYehmu17HRc1tg1uueO105
hKLw13kGxOA6VqJ9o4MWM0ATkEPBAB8VXlf5ypqGzLy5550uylJ6k6FcEInS875/gYPvZ2eUY4fk
1EbDxw12holDe447gzr0gEOeV36KcMIKHYfAe8qVFPirPmOsWe0qhQDQ5zCEiWUGq/Ncakq0/f0N
G2ngEouI7DiaX+AKPkxpbgRp/6moloM/ZZa69Zg/WZuNOcjYdslSmAtGcq66NG3A7IKI8+6jsvi0
8gR830vw4kGMYyQmOKVjDuTcEzSJCKu2cdK6Za2GfGeGj9GODGcpJQtG9wz3rlFBfEudCh8omofF
cHv+KGDome6J5jn/3T3z8NrMvbHznWAyddsHMV+UYHCQbXGE+7TRhyTfvpdXT8hjlz0b9ak8THRU
jyJgMj6dcdkkPnO1NAlg7zddtbvK/vYGKp0p++9t1wu+OXW+PkL0+1ClfBdD4UIrn8AIrE0r27Bw
3W/5NurX5R75AhHM49gaFD8sFX2g8yyqrlY8UaozHZARGCglrZuJpF/033Nxe2esyXRSv4HR1aU3
d2NMtT5uY+Ck4TtA3+eAj8bA7JJxByFfJEYA/Vwd+9nXpR33GEiGkvPDLrRXO4RaM9bk6Bzw5wve
S7SP4i9yRlg5oKa1InVlU2mLzv7lU2grlMZGvnsxlbGtRCDgXaLS4jPCBKRQG9KIsjto7FzC+TMw
1XH3ySOxmbWuc0/LVY4npnEFTKrI3AvENTONYaGQQK6Du9J0FsF0DVsAYN75XL7XmrYMMbOJ2JhZ
Vc0+/I8MvhjqCTuJ39ntWx49dsR17QfRnIxivWkID/AA/nn6uWVhO2IQwytB9jMhPYw7i4X7ofXt
i7qd23iPJ6tUeMvT3n6LexIBkM3F5BZvtBM+aQXHtxCgHgAOeBOwB4QCnma7o3caQwLK5ysrnhD9
UlIPl6wWCRgfqqIvesA4NlPs/4eMLisqrWPaiNqdTkJEVE37CAlt508wg78JHUUykV2qEXmZbBAm
Wdol4KLwp7fqw2c0Y+MMkS4POt7/CvP9Py7OOfwBE341E2WBm3wZNKHAS3oJ7hdTvtdgGEN5eJj5
drqTBlSY5M80MGVuqmsHKwZ0XSjFiTCjxSn+VC/8fSVbvghxFuYlYWuTPSyZIoyyQUICgUqgOUo0
blWxJqdJMecqxzUq+k8pNV1qu2I1S989lIqDVK/alEuOaOhELsLNYwyZmy8S/PgJPMhbuDRWuCoa
YY97quIHK04Xe0WiMteb3K8XoWnUHzlj6CfCPo2qJiiZSsaKHSckinHbBYhT/ed7i3FJjKdVx5aV
ZCm5ClSDCa1aKQyW4bx8Ii2Qjd8A1gre6r+gQMTzcMeD4/6qLIm0DMZcl5ONKYqbNSU6Q0svzvVT
uI7NK06x1QtumE5t19fmpdHO8CeWRtE0siswGTU6enlzuV35WK+2/biiTLW81nFpPkNKKH53Hwkv
+oC5aqYessetYAAM9Axh8AHxTq23unt7UzW2o/rbEfJ4tPn0IrDZXbg9PMcDJms/1Kr3M8wxU8dG
vh0jxpzjPrRgA410n1AXmy1bYrb6GAbLcXqVRoWG/adTTNd7IVLBvg+zNmtDUwtQtUXoEBE4nHmQ
+SR5ylwXm3EzgEMfu5R4c9+0YUBzRtDuClZHnKIQmrUcQY4A7EHjnNqMxvAocpa2ftLZIlVC25ru
jamSxSa8H6kkvl5itkciJMt6kZl/sNDimyebWMI8VR/riH+dQF9oeR+b2ZQCGhWYCrF7x3R5is74
EvEH47npDRxzMXyDxLTP11lSmKyEBTBz6tKhHaZn4rEl259wOJRTnf/qMPD8fu3OUU4oZYKZiTik
QwekmhU2EZlUI9ZxaAEnL+Ng8gjCypPJKhGPZ+w6iWf2XA4TFQL94+2NhMSV5Vbx0oV/4DJrvGJ3
B9FbEZN0fbQiFPsSXJKbpgkhDZwxe3Np9PzlUYemVcM19xhDaSBT0XSFk3z9qIqr8q20doqdvDPh
bnMSiXb1kXTsRDsxSJVy/K1NYAsV+Abf9mJKMpgMTNgBmZPnY4SFgHnDUAjgOHZydcFsfSDAAgKw
9KtF7LZ1m4UXno5VoYe9rtBSHUIdsd5tTt+NPvq9Zz5sgil5bhjhn5o1t/XsSWC3CdKQCBmzK2lX
AJSWBFq+d5l9rEV8px0wqOtW7hA2z/ULly4rR5zrlRC3at+VarR0ZQ9n+Mxin5a9JI5Sbuw12BN1
B03fntXgsh3K9mFt1+AxORdtEkvz/kRTNb0Boi6puW0IgLsEBlL1n98W2GyfWuGZo9k7ylAVIJht
1RUAanpuGyRCxtJVNIAXsWBk2HYhENZ0JVWSf56lj2xMhdbncZq0MqkO5UBtD1q7zxbFJLwcjY1+
az5fw5vlBh7kD7xq+xS4vIo7IhtvFwOrdmm5ad9weairfOboGxgsNWsmzfIUPTfu2TN7nkjksYNA
1k0ST34uFPbuwsMUIlXwVkueGm3DmxOt3Hd9HWuMySZieKgZ4tZMig/zhqGxA2UdrHHz/cMAB0cZ
yPZzVepS48VWAoQjsG4qYCGyNg/hlrPRMKJB8LkakySxndHrtIlhD+qi6H7PlX8/nUV5kwhJIwFb
qMnRP1V4bxcxdHeEOUPYfXiSZ7t4GFO1sNb2dp7KvckpwJGqSjNl0c5jLw/vPd7tbSpNWy2t10Z0
6sLtfGusRafEkR+tvyJknQhgOhrbZRF16Mx/efYoo9hgTd+/lfk0VchH3eH8lm/qIUl6S0SNTp6S
Q3UTnwTd1hhABGO7P9mZU7jQpmNLaZT/O0UEyy7igQMe0ISMb4btwIj5gYwq4GFCKAh6buiXJq2n
gQp0GkjS/ii0wMhAbeobHoo522/OWK1TZnHeTaPRoYKchCIwPbh48TN6iQpiilJt//QSvB7fdp8/
UQc13n00s5W11XpUV8lnlm4E/AoQjpM+JXVitK4TOWac6aDUV63uvcWZkG0nidvLC5ysC6fy5CUA
ujkiz34g+QuVa37jLAgah8xBg/DoLINEwmYaWKPEpABDUN3T3OI+JSM6YVo5J7BlLSBMmicEjIK/
jCXMCJmM/WYD4XAetAfuzlU45k/wzhiy9eLX/3gNC/mnXaNbdjWEHn7r7zpwc3/iTKfrNPJtzSxQ
fKYRWGsM7FuaNB7sPpcIcVqvbWZQsK0x7xz8Se/ejKjkVxK0CGxYqqdkJPbD0g6+L1qAeD+r/E8d
dhsB5XwJyHmYl+eQFFjYZT8M6JMQr+bILn/7eEcp/QSKDFvOgI2ad/zzVoJpgUYDb2LUmwT87w2Y
kOPdmIVHjqykseQ0W9MY6pvl6dnsbP7uxUUEnkHyhr5a7SVcRUk1B+lw0yjAaXmbRrt9OR1x4Oeg
aQKT8VjXGqZ7pdlIx+Xpqs/aTjDa3U4nZF76NHJZv1Nqejrby4WZcSrEv9Y+J+O8dMMV3dLjwHcm
XgvIMs/frSYEAJ19MbLutHSE/86L+YN/KO9sTf8WFLShv3DHtq7QAtXu2iRlFWEZrZ88YeZ4yZ73
szeTlTQ5weURzVnyPgFEsBa1agf5mXyafh6N8aabV86GX9UPyAz+hCP3wA1Q4oct/yU2s2koOu3k
kvcsS5sBUFno6HjnfqkkatZGglnrT2J3dHwyDA0SPk57OUc3Eumoa+KaIPY3oNDz6APaGwoUwH3G
LBY7oQ3AHzS2h9RQZXBOgOk6XPCIe1suURt/MwPOMGUagoZqzse0cfALxIR7iNoDT9HO19yyV0k6
WxobjUlt3T0Tbi3uIGkLuWMkfFO/4KxDMRDF1oLaYkTymFjEMYu35Si5dX5iNE/Y8GVDR3X5JLsD
YnYizFqvC1S9pfF6NdjRVvKORUn2CcZ1q3AsB8z3Y6YAgVb3hZ+rNwKWRWfX4rNUTou8S4HsWkHy
stxipD9LLvqxq0/LstvW5nYT1ZBTdOCZs/IE1OPArx8UDXh3BLLjXOpzIocM9txVxzmuyyVbRFr4
mMiUgnUWxYH16O7xjfM8pmlFky5jI2O0fWEOOneFZXTrHM7gHV6Mh4YY4EGb9I4iMZuiw3/yJWgy
xBLJNNIW/lAky48CU5MpoV0yF9DoEDCyqhdJo7l9EhyfF+MrFYRDjPdHNX7wSNFoI7UnyPl+cQJo
q3dMzrzlCU53XZf4jLWILzjc05fytF7yZDag5e9e5gwAC1lP2g9uAEpcPWskUnAv4T5bWlbW1b6N
aGFAo7S12+xNs8fiMnCNIhoZGMkL5/zySQq4rPtOV/IwYPQYvdWB1JdiH0u6UPyAQG3fJSBDE5Iq
os6Xa5I2y5hTW4CFHA85bXVWp7Z1uKhEgZsHwgXbrk5APx54sX/t7JF2soVVwJeImf00JN+O3fnh
vTbWv+ITmZx5oIwUkV7oSY+/QQMkHBqH3sQS1Z9Op9bFikh0BMuhfzRyXBBDwQi4/VdPVvNyRsUF
I2OP8m+Hk2cEnOjbFnWRBPtMqyY2qqd1zFDAgnVkyBRfF2BFOUnvG4gdeHCRQhaC6TgcfkiVLeaI
krElH0Rtoc1GxXb7ikSKXpNZQNc5jBnRZIYB44kH2msNKJkl8sLyf4zcoySIOLnvEq+/0f2PqIH+
OHVUDgs8R5qJSrl3ZCHMww0xO0+ixPSh2R5iY7tyxrH+5jo29qBrA9sqx/NqFChOZ81bOxCEuQXl
O+W/auqWQ07YjYHw+jGlO7kCR88vlj6qb1c3Afj5zzp7YLKLfXvZHJFbo9/2hdWP9Uz3mdSdRaAU
tFNA1WU4+TslAf2PXRFpmP6pQREOLoQl6sILs1EOupuxJZzi/9n5856Kfylbx5xXfeUuOFShbmVc
aiZYOUPowky/QyF1ee3eKIgkqtZqrwiLXTdIQlAjFnEHL5gumk7A7Zn+mAbw1kLnPbnTGgPQkAiH
GyVusM24DhDemnvrG1/CHsp1nOx0+Fynr5TpQ8lTefHXuhAi6ZpfS6E2XE2x2N8Sd2+S4zhx+0Dt
ArShk8jBZY0u5C+9I2+pWgcLaeqJwDnctmjkL5WjIr6vHnnekMwHC9cGBLYjgjCkeFRrnhEtBHgk
usE20tdhLIMde1xcIoClM5G+iR9b7e+0MnOpUHkBu9mitqeQz6OcmwKnLghQjcs3HUOiF3T6+bfc
t5GyPQdwzv4GxurTzTmxxFqsg3DYhubrgGzQ818ESp+RitGUIhuI48qrtU3KB/thAJKq61DIJVc2
sBW8OKLgBnRpr8N6SnmeJZmE+nQvqs50c6tod5666eHszwhJbmju4cogE00/EKYnIjvp6QpA+o6z
ViR8SWHAehFJIOJHMxI86yK7Tuww28VyWb7JrupNlL9gni0rFf8MZCJ9p3LkNtRYsiLHZzdN0YF3
P9Rc0nTx906QK+CqGFs9ZC24Koy1MQnwELmb3hDbnoXpyL3wFgma6ZUM2VRl6v8r9xm9t0zCj5Na
2ckA3kc2ZYCD6Ezv1s83n2v+nru5IPCy3CN38JjCEdenzfXuc0ZhgrCP7QHE0L5KJx1MWK0DtzoY
fAo8MAyJDVqRawqDG8eHzxj+g99u7SCa6hBgQQkBHwbP5V50dRIHzNgytbNznv21RyReVLqWAfSR
ONoyEJHxowNGwHiATqlz0SOoSiW3dKAm79GXNW1xxIutTz1xxsluxRYv6i0byeNDUwV4+IGBNOvS
mS+oIyg9tAnJdm5/b/ojnWggr4zRu33EdT1veitPUeL5MOldRkwUG22HUxFgpz82qoVJLUotnXve
uGEDFuz5ukU9qkj4Qk36hnqQViN37+1G3bVUkdGdPiNjNN2pY8hqJMUCvZh+eyKeaCCcDnutXtGs
/oSyI9S1fpVsm0ZYLv53IhjM8tXqLSO2b5sH3iPwTVAUdBlk0GncO0TgKTuE5mgdTatck/CvWzw/
6rfM0A8wTRQbgKMHYirTqCdeESavyyaUC20J0nv0LrDzMaEDgSxMCY4XY8nmDykqYr8oAXO+1OFL
r+PltS18thHt2zHWz3NQvSEG9IHazuivI+ampb/x81tes93Ih+GOy0Rj+VpomjR9nmwc6mRVkPNW
tIhTjvQOUxX8XJzt+Q6I1XsW/iPfYRmP1ksTq0wb4czDBZvCI41QSsslEznXLq6Cl+RS1LMPgSfF
DLaZkCAmouPPQoO21hHYXaJHQSCctHflXCVfTupA/aOrg7d3/21eGs7jwDaHYoDJMVSUCJIwWnLV
fFowWZiNKvn3RnoXRPKpZwdrL3KHBRJZNoXT5ZzdJbUhzLUODt7YLox0f+yu7zobDmW8VTcLfsD6
suOteBouPpZ8CR+SKCIvtVp98lGE+NctbArrr3FqEs2VhwuDk9dqwRdQlO5Apd2DYUURn1iJT8qh
JZDb60DgnMVSV+e2nWAz+rxdqkrSWypd+v/ewjllFadQ7GG+yknPr2WzoRS4IRYhinIMScVXlPbz
S0S7xQmW9HNMJxcPo+tGP4FIIhnqRRkMxPL/wXGSZmWvCe4vSnArQtQ5MCU0ZljAeiZDCJHpR8+v
P9MtRCvoz4+o5ACfk4ZBaJ1pj5dy95z20vDri/i05ZA6UytTNkEEWMcVCFun/I/Pp128L5n3m0oH
i8xnTEEWw5B57snlsLhPDu1MnJ2w1qbnjzOCEdDUuKrxnsY14bnIBi8puy8kkyY5lwUBTIULF5a+
SwkBgWgGVNpgh3L8ZMz3Cn0vx3NA6/+H8Nk4uGQt5F8IpBg4+Dijd+lWoXnJSfweJZE8uCPQs9sr
+h9aBTYetZrJXkoh05RdtwYlkdSFPwCEq8qERfMjMq2UoFmf+NSqJlgLMe/WXjIh+dgSEPB6Wy9y
CJbzlhJL+mV7wM1/BcPGMhd/JQp68pWdu4fUfKnn33zdbFcoKfAU67CHdS/SNKcDq9vlTDe8yRPl
OsuBa1Z/Z89zaNUzLmqHyd/agWEAq9s5r/g0lM13y1c9OUt03Gz0/7bNKkAU0aWP9IJMIyIOGTKT
bCKSNLe/Suc7D+P4Vf9DifNRKVXvfNDY5OfS9ovLXuUzmh9jfcvO0+L6KLM4d6oruVztCoQSnM/h
nlfbwWpCejxkf0vGvCRr+AyFNpCm92Og1fXg4lWRR0ri8WH7DMLy+lUCW/OcvM8kMJkXEyfxcv6p
0fVxg9oHRrtKQxv8Vj1otXXlVdpAczuK4GUmQ7gUphAafQNPCWqGCoXj3gSlkwCv0hTdBuOGY/rY
/GxOyhJBvQe7JIAVj83Dr6K6FsPE4Kc7uLjnmolhSaE/SErWZHU/cvkF/ynqLJsM98or7nIpO3hC
lVnwwegeJECkBWVq4PVRcO8qPwnkWrK+XXFyHUc8hUL4oYvlSd9kBAXUpvinIsNpR77efRp2zSys
j38x1NqVrC1bWLSPAMruMpq6hQuZjHNi2BiS2nqg1LsSmKSoeOFXhY4IcOaLOzGGN6klqV50Ym/M
EHQ1vEtPX5A55aKypL0U/7yv7jOZHLl5fZDCDxMNfM6J+yPjpJQ2ML3RWi/R8jWJPQbJE5gmxKQs
6H2N4A65hSmDMIG0+HqqN1rf8CJ94jzqEKb598dqRY7pjTE9HvlIAGzoriSguPk0V1JYZhQVX8bR
iXeBAv9m0nQR2oxS1Y34NG3YsBa7/Io+Nzay0wSlM+H6h61253VUayXg7OERLt5h/Yk+mpYnWbqm
H+8d2pcTFSZzwW3UmpJiG6NSKIwZ5d3JY/7vLbKcEUziyd8CkmpFpVXxPErPjXH9lPb98s/Gq6Bb
M1eVuvZ44tdxDmH1lhjcpnuLPKKQKNZHq4e0QafG2DJ/DzDUT8C992vS3S62TA8HmTsJ0qoiQPR+
hjOoYUZpdJxJz8OAMZLrcrGS3Zu1Z0CHSNbIg2OMcN1K999y6i+XRUV7dokvJ74iBJ5/QQufgTSp
DxvIUnomVS8zG4u+2QnLLt6XeCzrc4T/+HzcMI/tyPLEbFLqgy5LtW+WeiW47twgDyywOzLN3CLk
ypJx0c8DPb5mFF1gYCYIdplPGftSCkuFb66riz56Mi+t78Az+66wM+Bek78NlwhF/uPCi0yV1FYT
+k6uE7ABUUPknnwa001fSYv9kBgpZeE7loieEHYvs0DxrNgoaRr2OL5zerwVI921cMIBWVLTTLuT
sOZFu3JSC0uGqUTXVJAGNIjHN7EOaYJOcyRkqKTvbzxuQsZKqpk+krMBFwAnI2paCnAJ7ZzaDsva
yqVhuGfeXQWD7WNZqflF2KEis1oWt7RPj7zbZbDy4D4Vm5K7FykfrrGd6gTDKShbiJ2oKpNPGs29
MRmZ+aNxeOaI6Lz2KKNwOkYPFJkGdekMSQwtBRGDCuQ5F6W7V5+YwxUN2rehn9fpTjDU2nijkbIW
Wlb6br4jPJrYD+SAohLJtntEYalgWicXNaXzI1uaMo2ZaiMzpjyUJzI8AIf6sSmtvgy/hALNVwCA
x+EemQBEkf0x0OSnwTe4qVyOg/V52fTjKovQdJSZuJBBWmzvLdQ7bHIG5y5f+gP6+UHBcUntzc8n
5Dvq4JE03Md1RMmQgdBw/72aRjLvKtbuAxaDHYd9b+O+pf/M22K10C9wOONkXem08IpEOtsZtN45
GWuYYmE7YC+jB3fi80cnHfg5TaD9tuK3TEQGuWlFMjIbGNta948xwiLbTa1i5NixwI6ykwpC1Dpv
a0MwfPj63VDy+j8hVlwHtEMDWEUiy6hhLzId2cw9x3exSVfqbHMeNzAXADUALJo88Fxxm6bdRGc/
MMNWrn5VvJL7CkrapWXSFYvo1Spg7GSi9vmfJXGTCgIofq4PgwSrKFnhSOLsdS85tN7SRS+GmOCL
BzRL+cWt3bDkxbjvmD1IuD2/rGZTaXNIJbPdDNHNMMqn3uhmQtSpEB41CWuMY6AQ9zhbDRxHJ6xH
pJuYsmEDYuqQuSGgUzAcQdpJjh9YWEyYXmMzxvcEQ/RgXyl13er46A8sXhuRZ6qZHW7EpzC9lsv5
zyIMPQxx+PVejw38+y6PXQP5lVDsNt/0XLbPxHOfrRuWkqrfZ9jd/oQ/WTwDfTZcJ6FCODqSQiT3
6yN+oYjHnNy4eJOU5OOhloDq+HWartZsxsy1KulsfnYn705VnKfPsTXlN4Q/ZYCSoJfpm61IdK3n
020/U2Txlrvd57LiOtMOniUGZN/v2+1mzAkd4w5qQ+7I2mgxVAY7U8X6uVOSRfosdSKLh6RHaUqe
0ULmZ7m/BCBxV7v75s0NO5ps6SbE/+akjy0hciYJ9UJepKPFJ/SArRnKtnUQflT2rk54oy/X6soD
VsSsD/XN+RpFp7W+3cau6qlHpulwApDGOkLmvAX0ekRk/Dyn8n/IjLj1t+C08VBPcy+8sea6gqHn
2VkF9QwzG1UpjoR2aTN7LZm6f3a7FmRGxW4rLjjDt2vPPksSm6yNC+35fzxStv3/KV3ZssQgFJJ3
qp0VK+ryvQZqgyX/NN1UVywM1jJPQeVXKbUcGtwHI9XI+OjKf9HHraoRGzLOuw2KxwpR9EtrNbYD
5J2YXlGXmt/hmS9A6oJJVi7SBt6Rl4XRZRb2+RVxuCPqKQysR+dWpAqDDEfYaSFouhMTcYuAYEo3
93PHpFwyhxlUmNQjjlruXxV4UOsVfYxJAeX5yjjZ/0dgSF1RJ/pkbI40j+WZv/E2ZDSDfIzFN+Kq
nQO7yxMB93fd5oLNj9JTfwT7fjVEW90jSNJHqddUbpHp/S9NpSuTc0rd0q/AJR9ivyk7vLpvyham
TV6nG/5HE/WqHxT6Rx4gWUCUck0l9VVYWex5TxXQ+3NiqXMdcuY5ZrGzVKPZfLPRSsiOx9E4J8uk
YtMVIpJ/y6tPIAX+gbeJFsbw2C2LD0B2StD4ZH2BhAxsn/A1YgmJcaavpIIostprtD9oqPcKgKS2
IdvvNpKNcyGoWaSsMV4KOXAuLJ/Hg7h38O0iCuXrD2lfOcqNOoOP4PTUms5y2EhF+n/mdCIqPrFg
e0xK9HxxABx3fGlrn7gfezE68gqoVgY6K8MuUUjNsmSBhzY+wc0sEBc0CoVAG6TtfCaky9VAHO94
lm9shT3K3JUNwGkbS6HdwxtBPapQUgzeOiSVx7fHvOATK+qP3WUbWvcEFHDNrFh0YtsMlV9q+FUa
MRid7C+DeNz+z0aBHXCCh3isWqg1em2mmkNXujua+LC9ECeiclJeUkkSaVir4taaqLW4O1nwDyhF
0gsIjTIsDFaEDU2+wPo6MqOXn+iNWxEtDW0McLi4saYFGazhKMBDm/qj9Ug3at6Dx8014HHIwA6f
q+cBqD7jNN7sxrtuyVJPktzghHVbpBAelOOSYWnnlJpPbggkrOc71t9wVjCEADBnCF8tOgYHnKry
kGlqI6xbts6hjO4vQBYsbVPhpsxQiIRiz3CXfuXgPx3B6gGg/luN+cNTyTwE8/5thel8iKOh9PF3
7DBn87tSkrkushgIr7T6jjHntKhUw2s5ahcLL77AOgbuzw6qwDeGY9OUhDaaKooF1m25zw5yCSCQ
mfd3dmYd81rCdkUU7W+jYs7KZmnLKwctG6nI8P+5UoLa0XQ7kjMkWkfcAKMbG2a/zywdOO+WpZHE
zYgeijk90/RXqKqlZZtet2xgKJVPeL4vkrmYjSOHRCENxcEOMo4KrIiRM72Rx5irejIipK70aEbs
YHIxjD0vU8wDDceHtPXN0AsjDlbuOpYqqg6GKZYViW2pmd9iRS9kW90BfPZ87/TO27FWUEIScIpr
jpN5B7ZbfW/8lJL5fnKuNOZBl2sydzoaSQR7sCQnYYHJ2cZHcN3chfF4ejRhCQx4gE/as86XZENk
SFgtJVerT4bYlP97M5u+9I5vgdi/uZz1b2j3t88//ouu5Y5huQR9WVJeLU2wAKda+RyMmRZvoia7
lLeUEqORN+6PaQOa+cPpZTQB8de6+fhocekazowOsm30eDxXKo3lZB6R7minK1iiBfbyfbPSJj6w
fZSJlbkCv2/eWsRKJdBcB5a9EKTc7S8jfQ43VNlxE+IWzWP/iPnUUzciMf9XD1fK1jfXqMjfzW+C
TYFxsrvEqYS0j33esNT8kLrlUiISdfLrsaiSosQmr6ZiAxx/mIUvusVqRLqAO1pSq4Su9LCPnZEY
3pnT6rv6LHsCS7YduTtM3NdnA5l+A06fCExlLkhcUWcRUt0+4ltPeq+HePCM64mrgw1vm6an4dXv
MfNTfcgE+JiBdwKgn3ZyNM8qyV0vnFxKGZqTvW+teTLV51nbKa5sXsJwtTx+xgfz4P3WLXmHU3py
Aibe8dSv7IGxZaSLiOLt4mMG50+ERm7hHbTg5JeaB7UR2F2v2lk4lbq3Hc/MWH/dGR9qSmAWvSgL
fTkz8uDIo4iGRkgwofKHAgR/ymOT+avLrCY5z73s/krV2lpS4cQEBK5dCl3lRy0vvxtas05X/Ljk
DJ1PB4scwY/q4x1kDYRpE/MmPccFVkYtOf0p4FqEE4XxDi9AX2bTG2NV16TyFI0O7DL1M5ySSBrd
wVnIGHWsdE8zs8K94eFtrauFRFdVapqxfVf3CpS+LpAdqSg60Ru4pPa0KpKKEym4arKtO9JeTQiU
zdbUCprlx5/VheOh2l3GfmCVZ1qTJ2lGLY8bZObCpUVZiP/5FY3dD4EnlBvnuK4XkOMkr1qfpNf+
YMOB9gaHp17STFQGfCF532ITf9EsgUlZy7N/0rKV4J2kzPy1fciZaWil5uJEPxmmWrl4+hF44Gpf
HhC8HFT1sub+D3QrsySH98AzEDJEA23dyIWMriMdoGLKPB5H/os40NVJsZPHcNAB1D0I9uY31uYi
uHwUw1XpLWHK6rdmINc9br89EdTTVgh4Q7bm8drxlpubFKT7V3u2qU+A53Hw0G2f+FhW9YF9c2cb
yUEOfRWbXigpAXsslQg+/QwfIseCjFCClolxFVKfx9SHG8VwHe+PWi+A6C2WOxadxCqMMzOMhzcn
z/uVKDnZPEC0MF9/qbGeDPwysoRTJHU0uhj0YOedJmsgQEDKBZRmSYHa2Ohr89Thbl+EZ8/jlymg
E+ghq2tFvnjDPxcjHJnQohjRr5GCwCOS0N9HWuzvxxqBz5JeXGwHGxvFB8d8b/Vee7wyy9P00PtY
xIX/4YzYuznc7e+AMs96n4Ala+pvTD8klQ4CnOcFZmlfsichtNs36MGa8CO49CywP49LRSzLtRzD
Xn2E2K3f6oM9AntK4zP52ZXF8BZ52lSQWhdRDkHzQam+shIEEUFu2WLLnZYfzk6ilyzIuTbmCXJR
9p538iMNFOrqLI3khnVNkWwLJbGJ5ZNg9vV/zyoE1GJneXjjPyxNZWccdgE2UZ/+mP/0PbHca5vr
crOzxv6nslWDxNzvTybjZUt72rnIFzMuj612x1GF1ShzlIdRaVxJQO+d+X0TgjBE9USTY2AuPnnr
0kzrMhvOfqnIsSgCHY91wsJB70oaE0AXZm4WdATywmyAM0LKGrPedo81u8ipgeqZPEuPHoI37vSW
9H8556VOz0PNBcZ9QE1CObs9vHU1nA0iSFhg8D2g40s7U8j1rS3sRn1ZAYGEtrGx50JF35zyFfK4
uznwSOaDc0UfrUP2gPHGm5+S4suplIDcuHuTCfm9gIWWocMBaAIkwmJ7E7YYbaKX6DU0vArZywP3
6TbtX+jV4akDSDs28uex3ObAQ9qOZJqG6AP3+Zp5HSeHYNZSwcxsl7HMkzY3ePWA+R1/wWLrAVBQ
aWlVPjlW2VSBjuBvkvqNVS2VHl0CTUYIFUJpO7wcI3Rh6TxZprbPYcoPnsmeUnb2kARcf6+vsvdT
3rA1PZSHr9IK3JoOC/2vEHC2NUTDyb2Pc2ppmTXPd4poFHoeVdlgcQYEJ4FTOV+3TKB55/fwdHy4
CWgtK0OkePm5KW7HU+tP/7BIriw7SDNW83xvDZmMtPuOWv7FZrPuLVtinBOroIrqlC04iIq7tErO
lpInG8ykQV8pey8uIOsPKzDRdfY8gmIMKCfMNxCAdx6CRnBvsXCUVuET5NNqRK0E43gPBlKEarty
SvJGBC7oT4ICf8VhINVyg9rTNAlk5uGmzMewuZRJ2zaPhSLVYZhNKV2l8ck8JzuE/nN3qvdvGOZD
2Yhmg5BgHhKoTGQ7Z1GmWCqyPUXEg8oYzUR2JZfA+1J7AARQ2Gmi4zA42fZ8CyhvwZ65Q1svAGjE
9CBFXrM4n99EX/8Zd8Kan0XZ1PrnlZwulxK305S3Jmf0E3/S/xrIaTDn0snpVRQeAm/AZKTBBLUH
Br/ogwZzuzbwpYOiH7zXlfrfRIShmEqYDhMp3BthOf8LNB2ljMPuQGeget1Ax2ZUg5FvWONpCa3e
9ZLJpNjhtsOl2tX6NhdyYJ0GSB+dQDoHCEFfhlJg2n0GcAEzBYUcTxwPfd4SemJZTgyKIyMIk8tL
cpu/NeBpiJy/KRVPbTWHi3Tcf7C2ewP09rEsybP+cJqinlCv5VSyJFB+u8kQ6qUiClCdP5Grbpc8
koAqX0OWJ9e0Ptw9ZXv5MwXDXgwvhJq92EduGL7NXaJN/1sdSWbXh2aLVwjMiOmCixR7FWCi7Y/1
eIRkcCtHo7LccAsCVJSmy/cVQOmJOiQtu1hT13mhO8rQ4keTpAZQFH2WDv9kKQ/vGLZhvpfj84Qw
X8O5+6+fGDh7zMtiE+hTJ1T+G44qUU80qjIXq4TE5RP142T8Dr6yC7yf+QI6WX7/BzKHr0TYnd20
PpdeOJ0lPSmKyBZIhjeGn+BEQBg3bk8jDt4mSJo0OibFWuc0NrIjVNDys9GvrqED5gKeumInlOeF
dEy+Z6B/bX+r7FGsUcaX9TlzARGK0ciamrVASFwXW6f3Tb3Yrdz1u65V+J/6I6ZFvgM6G2lwz/Uz
7YUIihdvihA7pnHjm15OB/5ipN5u7KaQ2YUFVsXaXBEXJfalhotJdXNCL+yuKq1/Tirkgrtkdkfk
YKQIszOi4Swgo63KZpxEMGZXUMtfDaIbj8+tZ6r3J35Nhcax3XHAjKPG/FOcSHgsuW1hKa0tHXph
z6G5GSLaqQiySNUTrxGsU0cu0Qba/7PJukhjE06T5dt1ecJOAHNH4AU2p/35gsaYKf5wZWWCJX2D
cm+eHUhUofHjOIlzPEZvZT/3uhgl86KBlt9oIsE/Rb9ivlJIjTR5T1v3RkEj/XpXL9rkNyL4lVjz
BF3vzlrKAyeurqSgB7frmzpQNqJXpzw7oMXCJyquq3YVDlVq/GtaaeATJRRw+MmCSpLOI549PxfE
mraks45pS+tksTr1ifyOwGnp5Ox2wCxU1KQfzmk8YEvyGcOR3WaanYTxuVOTeAyhJOoNc4Cme7An
yaWiF7xdBSbOxy48/5mwkDfP7p9mf8yF2VQq7Bj7LlVrsBWV/JaiDZY5M5NmJfWhzEZeJ3audu6c
2tnDMM/49BF5dw35Vsb3u6+RXVU6wYc9j/LX7Cj2VHWjVSK8prjaYSIMLLOKiQNbExaeDQbo7D+5
bvZ5dBwbmgJcmW7tEFhdhLMFxV2AcFGxze47NdGj7mf2wPBLeDUj2K6LvneTSJstoNd5RJsuWpZT
EDv3HERtH314ovsmsPPvwStwC69Kfpdx/OAPkWk98nzsw0Az5mHD0O3j+GEMu3wuQZyFKeRcdWzT
mqmhECDPYEFY/NUcvtxGBPa7AYNpxk6aMrfZ6lfbVqW8Mqxc8OooemmgYxOGqGcYYY7vDza6QEma
bfnnHItaZhvWYVYjSMOXLv0+xPe9r0r6HmZ4ZDvEJSxy7Y7tD1xLV5yTIrPo9j8w08gYsQ1PnNxi
NEeBL/6Nrd5YM7HM1YGR8yE/lYZHI7u8Kd46WQgxAWxHH3Yui6+UyJg9KOE85OV1ieRvMClD94KH
5xczo5DC7vuMEOYaAtr8jCSC04xrIKXIIGzJcMEDRFosYwzMSnU1v6c7TDU1v/DR9bNCH/cb1EGL
YkAqvUh0h/fMnj0rddjCR1lXaTpaVbkXMO3fntqqg0FO/f3eJlZsInvmgnQq/TeCHlETTj81le+7
mdMY1Dex9QV1zfBdcLIj9i2SYaTx1EPFYw0nRpOz7IhzBvr3Q4eunnjECxI1tIwacQIn6Ugy9YCk
NwWUhbNji8WFDKTWcVZIr51n2dYtz7KpTEAwovXUsXQrcWl/lhP2b9qwPTNFed35Ns9B7juPx7J1
U8ljf138vnnZUJXtHpcblq7H6igqLmUk+MVDX6Lqt++9Zdi/4zqaN7ylsI6SQP8fCQVxLmBo9M+b
t8Q2cA2+KkYeHiGXnQfAhThI1qSdZP20AGiMI/JxlVtSk5ixCbu/sL48kXHxSNy/rDc/datve9O7
EpeotePMkaq/P2AeSKop7TP/VhIPzTf7hKn+3pfqKkzDntLSLKy18B/FBs4MjX0HWgHiwLHNeBFo
/tuMBnwUy3i//Yv4idSsPWGd2rrfRHkl9axb0sJ2nJPCxqdOZ4JySQkLjV3Fv2Sbv7ILu2XiZhQS
WdDJQtYa43s7F1EtJ56dsZbgw1pS+LdF29FWjOG7rt1sSAIV0Kbd3U2pTGROkQzZVH25KYJuJKpi
w5NFb9I/ZuwdS7HI1YbVWYaLR/jNLBtKkeJaXrpN7DC3vkcJmGzSmUlDeIYR5bpC4NX100x545UN
gyKeQgTiZOd/uzNtM3HeHjG18Bu7A2GkHr+0GjqizO4QgWPyMetNVtxAp/oGZ90sjB6gInuqFcHc
6lyfz7nfGfSYcNDN07t8JRXmsKkTsRDKFEWv49ip4S0tmZx66G5yO0v+655+N8RFzki4FZHAWjjP
YMOsdhpPtSfSalryOA7xvRZHw319YD3HG0HAREj/g7jFEdsniJX7bFb7kaPq2CSnEJBb7wU5Ne5Y
EjSfka29lxLOtTdPszJryltqzl9n44o8vpbKyPQKUHfNFbxdEzJ3QOYTiz4KkxdK7YhGJJzbkuaR
G2pKxzTbc5X6DCuVyq3us/VFtijE1qOMlFkRvn4tchI7Gei+3xP22cNw8xvFkG/Ui8dJQ2c/RUwQ
Xji75U2KomKIXtEl7yLAYAmT7enNXZyVfbJM1qea0ykNiOGCReiMaYfIz0SYBjCa5aNSl+og5WZX
xBvVQG6CYl4Qeo4/fBo9YVp391PvgqtaY2ncqwbopR9082Juypwaeq8sFeEpOyIlAt0nQLAAqgXg
bFlL7/kpnD7H7hhaUclyPONoPl1MZNpcgGcAdYHP/HejafIenr0K5V2wTO5AauZWZlQ/VokoZACX
i1IDpfN2N8XbOQHz4HvlKysiRi8ySIwctjB6qYvVqQ1PcQ5cWhqqQo8OWMMcrkxwm9QRMmy4+fgo
Zg1DYBojBcZuUY/wILIwhcmj0R21C/Kst4PFgNNl2RPu3YxfoQ3HxU84Zc18XFVDHC0nTo5RkkNg
0SHG4d3uLBp8x2iwhmvcLm3LhVBlNLuYSA6vHBU+SOFqL0xSRJmOBCBbFgZObyDtskUkKVnSbUvh
SuikzWxPp8DXtj4cfPS6ErzmtxjKpluKAeVGZqsWvP9wIe375l6pSePnTA80cG6pC5Yo6EUQ7Rgf
gFJ9NTAUg8ZX2iVglpWvujDOv2VsIaOII1yWmmlOtHKQCmDwRMmuPpb2ZyeHF8ULY9TCz4WcKWyt
XrxjSYBzXiwKsIlNp5YndnyqSGBXMEzuNvNuM1Wnwxexj8QI556PnlVNO0zNRfUjpdcyf3FUpWQ/
WfRNCfLyN9GXUXWAte7mY5QLkvztun0xHmhWGq4gnI0F9K02y7ZsfLXb33/h0gKLueV78tOTCv9X
/SWv9LXo7kIZ5BXHjVJsWjNBbx+ioOOVHRH9QoVmziFR9hN8SZj3sXPLZOmDBEKZG5XaoIceXCGn
y6rhnehE7n5QcOOSMoDckvCB+TF+13fTZxWXfKiMhbqf8YL514aekJPvaoZlxs8QSbBKaTl0KhL7
Dn3grmf+itMkAZJkV7OR4gvCY2VX5gErOKYJo6XUTH3Z5Mg8QPRPf9YvLs43FLAthKflzzJVdApS
n1CFFfDTo6fzcKHfrB+ujP5uaW7kIQeY0Eox5wJPfPIXsuYCIjhMl43ESgZOSq8y4bf907G+zt80
lI0tJWEohgTtLUZEK/aKzuD1oufCVIt6+Vbk2jWhJCfZnrtWvlXVP4VqLqaf0lWsBHhumMBZUI1l
1003o7H0rK6GO3qNHmfWFhbmj9eCIDReFWfAvZWQ50WQAYamDbu56CM2PMiDx/E2hmNDvtbA9o62
ysHwAi7qN9BkO0Md3ZdRneBV9lJLLJLDhgvJN5YC4Zy5tZQYiRAHxx3vwl0xNpAzvgZiLH8u6eiC
W8D7ZCA1QkySfw7+FSgVSEUQF+RmCGufmOpVZWxcT3Xz/+Hzf7+XzJH8cLkTFtbYPzqgZSBCU26T
8c1e1Eiw/9Z5COlYO2snwX0LwfpvcrPp75wL467A5mghhNxInproSz4LSG61cABx44ic4jevOvfE
JeoI+5AkfGkPkObQzltgODtr9KNR42kOetjVd6Dg/txP0isBaSnz9KKQdn7jgLyK56OGy5sNazuG
cvfONp+rE3IZ/kDnrqfQL6+Ogi55sM+KB4TptTBpVa4btyb69uhHhstCY42EoidqgGk7qLUHVjl5
Tv4WSbJhZmKMorkEiqgsTn7Hq714PgBglR92c8AypAaUrFbTkexpo9WnFZcqTjCQ9G9Jm+HYZnll
hioYaEf8O1Yf6z7WDbW/uVCxb9FzMJXiZWAQEU9XlZ0pRY1HgAaD5u4egXdRMa6Qr7aTaLASHJ3/
mdxmEMYWeNLTx+2iQ47sAZXhV/zh7taEOOWLPZDx+ZA+iM1FbBR/LWzm9CtebN6a2xtrl3IqRtTS
/L0T5P4BiNJamGPm0kxoh2zIAvmcF1WKyy8ZQmnR6w9+K7kE2I6D+pf0AgahjGVXsn3L4DKyTAc5
7uYTyflYA51pzBOgE+CudNz8Uf0lk7nbBhl4NFjkJRyljgy2sJIm5atVBinftNp2lJCMnqNpT1Pe
pQO03bUSGXV9u5fHW5jeYs42d2YI3NydEmC/3W2HyFZ3wanZKrINrOcRT/2cT7VF/61Rdjofj8Kn
ezfkrXTFt3E4tul+meuuF7KeVGGdY2X0HiueB3S59vfFuyJgVV5mS22yBqGt5kpQduCybjoScgUc
RXRBo+nROO07NTRtGioekC3cqngExmUBP2syu5Sl2iNdkSMMllzIz4I/CAFd96wAAN4AjIQMqWvx
p6tNJjhkOghVqmfegof+jQFxG1ZscMmppsdV1Kp/bEeJ0Tee4xE5mWmK6mHTN5xO+bliN9mWOVVw
Nxb3PV3dK/J02D98W0UQy1WxvisFgPa1i2Ad3fgHGER9t/Oe3FYaPbk7g8a10vPxDskWJCTfdWfy
nE+6aUXNkPc8FVLUFFAJNMHqLb+yTBSwtJ1FCCJWhXxY+QReaYTwzuRhQ+WFvd/UEuYa6SPK5tkN
kiOqy70Do9Ea+DBCxhNUYbtezzFOdpnofB25up9+mMyC94Pg/NXlsUxAhb3TTsxEql+pxuV3EEiY
5ZPj2FR7vq5k9SwNaLp2QKF8RL3V4tBK/V7zn3A+3hBfq0YCNw3cuOOtMXbd8TdJfpjk4/3ZztqU
JMXieJx/lgnTsa1mlCJrL2DX7K2cfj6IzUj5Nfop0W6h0tnahHuCdCrwjkVE3vh6RFnP2Be+hvj9
0V5zIA+PcH7iAPfjouP0+RIO3RGiDfYE6WwZXfaxvFELHDhnEEC3ZVY6mYWQ2We9+Dg3FkXRuWwK
hMB1vr+5FYRp6v/Qf+iLadUzWApWbql9yvtOTjOcge6vqTqKadfkTBlcOEtHln5QMLyd8BAxMrTf
sWO/AWYPicy6pADB8ZTSUpWr0RtAaTgFLdvcdQDPJ3XGiVDWsn8MmoTApMLUyrtKb3N5mtI7Yit9
sDzEpG1J2MGFVY4W82dWEAbu0Fw3kKXqHQAOrM8iGyVvDfZUT7Oob73CFYx5etYd5vhrqUhg6nir
Is8EdiViCilp/DuaJIkLXKe2ZdPApAREy0L5GD/SL+59dHZvqmqxphiXYw+xb0HzV8MHyr7bKEQJ
lS+A6GRc9DZCbmX9+/e1cl7TMZF5cEDpuWX/bEjRdX3Jhope690m7rQSJIm+tAQKGosH34urnlbq
G4HIsNkFzaKNcvdE9+TRA9AXbf9m7uo7owmVdJKFOYm2E85tIRGRH1VFBSPhC9MlWIczJAVL2+xS
WS6rEmhf8DrTOzgvDyvXKk+0FON25mXYf2lCHfzMOwUcrCBW4RfgsyyakYwjhcZhkWF6xzFmvMIl
IlVcHt6GRVO+WaB4ANSP5jgAk1J1UI/9LVGzswZfT2o6BPhS7al0+iNR6sYRoM1MJpfx+8CcVPyv
i0Q14VuYaDkXRgCEudcJXceA0uL7vMPM/sH61rzNsSmZooI3B5yRGgKyL0dLTH0Z72KlgAqdys/c
W0+CU3gwIgvxUvObsJ6RcGopq3sTRATMTbgNCle/CPCXSHr6pQ3uYF1h0BEI9ULILQguGVNH//j3
hVL555GpZuZX+Isqn2tLXephl2pvq0fp3AREsqkakG2bcIuqqky7/mESKjsDGPce3rmgqVTHKJRW
6s65KUy+Qlu/XA2JKjW+4WAjbA498lQixg8LwJLvJp2mrH9dxlGhSeKi8So6aO+7Sp9mSRoEbMoY
DmU1SLS+U8VJM6HDeMFye75YSoTX2FGjRHTylcVNzFUwT/l7DD9u73rOX6VkJfjj20C7jW9NyWzk
8qJHj32c3d2Xm1AbLUFH2zgn01wlG6a50P35vEXjXqvEnN/Kll5oEPjuhbc3yyje3VoWNWHtDw3n
5PbSw/I/9Z66Vfared7aF4VvyIgH0JY2Q6R88C2U2RCiH1r8dsp8PvgYB/Udd1uQii0COIic+NNk
sIPZAHQnpDWlMwBlL/S9xd82A4D/cP5NhHkNjv+SYs1PGRA2wsnrC0UStXS+B6BC9R0J+2cvXfaV
eebnuqt9r5+mdl2VFeSTbftxOV7TTzDp3ECj0fGecjcVNvTovBxID2YG/IxYP/BNiyofi/6oAUQ7
tvH1O3MthyIQ8AZ4PVtJwSf0sdaLL8hUic8wdt3Vb/ZDJU5OizG+Wg1p9XjxE6FDfwNVm6sUHe04
IvnnBPNKhHGCBr8UvRBJvnG7v6i7uDZUHmAkTbjmOMWstiqqnjZT/HWaBmrkRGVDB68RLJzoehQa
s2xc63u/rERoh1s3OtL5+/SR1+g8uvfA5t8FbGfizJioXsw9xj/ml1gq/sBPOcnDnSR+YcAPgQfX
QF6Ursk2BaJrD439Mwk70WafCDfbFgrMNYgyV+Sn7/IrMv5bUStGS5kaPE/A4RmNElG5RxJZplXA
7TgXfY1waAeCCn+u1IoRq3Dng85lko0UgTAyWjWgq4tGlXjvX0mQzeDTvk//+hZLbu6aXsZyeq4a
KEnIqi1QkZa9aFPPVFOOhvoEtFSvdkm7CZRXlMtbyDg2eTx2V42x5FoObjQxRhP9Fw1+yheLY8+a
W6u24O8YuUQ9sI51dOeOpO6nU0b1+XlUbEYm6lvY+DDejKmiqoDeOMa9cyMM/SBNoyi5kkGyyTcd
G/mzJqum3A3OmUCSJvoqB8NqNluZebffg9cK6kVC0UHL9YU+Le/IhA0p9Pjp+orYef+ChRaMLiL0
5dx6wUS9/4EpQ/12zxiNDtrIdgt+DlngQb2Wc9IdUyfAf/EhVZoWhme2Yg1hp1+IEIn8PjHfqKJ1
3+E8+bln0TVfS+g9b18eC/LnP5GrFn2iWpOllmqRpF9/d5ZFXO8l9kkL6Xyp/+neMBcFRKIAmmYD
A9+9qSP8OVhFaLazRhs42grjC0IY2LLfJhTsdLcpCcKFDqsj6ZHeZkxh7wBHlWuCgguJFvGJ5F0m
/uLxhEmIh4srEkDJHuncg/ovk86WQZvGgE9G2xUFtcFMbAsVCdykzQ6MkwT3efx+Ij4AVL90XUVk
ncze0SjQDdkSon6fZH7TRtybppXyhW+DbeKdi1wLWVt8u9KkKUSPdJVltJFZWkjmNnpoe9YWYqfF
139jvCKwQig8XZLVsPN+i4Mbh2j+VyxoJq1SIkAi+J2ox3yCdLqaigDGl60afJOjgfH6r+SNo09n
yW436p1z+J7BCEgVHEWQ3tYaAFI01rFAIlajidJxrknlF96V+xMH/RpluD1KUY1V6xczavbga1/x
4OBvov7ddaMFRzmu6CK2rQDbJME3n7DmHqDJi1fpSKq4fchvICCITBiC9Nxz7yoY2d8VtRDkNZtX
YoZ+NlP5hIJCWkptxejAiQnk++QlRbERXfKiAI5ZbejeZLADQCSpGLpmmolBGTXBlD94oZSeKOw9
ryukWP/WOB75CmbtRuXfCu7Sv1PzvSk90KnPo0M7b/57FS9HkkJfI+tCTEdcI2w1LD2RBgfgn8Sj
12DJJ+vHL0BwS7xxTI8FPqbFNGQs2SLRvlWElqpsyGcUoJPvRklNSe6aa65/Q1OMCqB8RbBjAAxo
EncnNWGf6KjVykh8gOXyiddbxewEutJZIAxqr5fG0IC9qi5T6kzgakkX1msDXKHiNtjHVxCiUoxr
Ug9mjxxjht9Qw+AtMGIHXKU3z6bWmi12mVe63P4ZRgtqjQWPHdDJAWPRv2JALy9WhH+yve1Zk2CP
1/K5gwwTTOySo5uCeYJ8TJmhGZlHbRRApqIwAiesFnaWFF2N+8pJUG3bcQmMkDONztgH+ldP537K
o88FPxvjCwoGWwKjXY2SnXts6779vT175PPrxREmMbjN7GAKdsyd62LOFWloIKb3co8wdxoq+5jG
JnG//teZDd2T6CZDA+B9HESiHRBLF1gHJ6C0XLmdxVBXj1u0MILI1iaIzKoOYUrmjc0DAsocZ9Zl
cumwwiiLMETyGiwQi1MdGceVb3tKNonhbDZlDo7XmGscBWZkn1Gx1kau8+50mosvsSumb6q5v2k7
g55qBmINLIxwlXk59BAHFLhJZ5JVrgVhXFPMgIdbXSjFaOYFGmaI0Hv7/4Gfdro8arF4LABTSoSh
wz8A5DSBXkDdXne/JKK9AgxOcaVUZGofUNnzcexTa15bP8N/tDVw7mANFk+pB8mPtsipLVXR4SWj
Dh5DdMlY18EbuUm3O5/kwYPIynafgnSr8hEFHdlKEhaRd0Hm/gE0Jb/5E4ZDfPIVzojhdmkxP3Sh
lSIG7TRO1Rw889O1JR79TVrkIW/WX+z73Yhz5u/8ANqlQL44AzBzv1xArL96w56c6jJFS7/vEsPV
9JXCLlzBdgHgvj4xgNaguzuUd1rGdyTZvFOexoTtJV2Y9GrX2BGvETClnDC77oU2CUdLF4Uf8dN5
X2jPph62pCL0DNvtPmEiWwu+v8etFSY20im/yNIlK5cqBDp1dtXeFgjw6I9XVxniWAVjRoGqQuqn
4EJ1I0D4uG/68PRIvS0kXBgQz1EX9FNdpgX8aytDJZ0Uy61SsH2n4ATzvKCZPC1tk2YXJx+zBBIq
O12IU7T7beJ9G0QF4LYSNRMBBOMKKfuMMg6yCtbiU/DuEdt8gHCsKpya4jYsiILphOyvZfeRKgZb
Iarrwi0qzA5Lgqaz3tc9OGXFFvI5g9ndNO6d5ohmVr2Xd0+x6kPRTKaCAQNiKUbqVwqDCf+TYWWx
9mNqZZ5bnWLIgdxLDaF5HHhKac74URGKsscYoMZjcWT4Yq2fBRTqq+wLHGqz3JGcrGi+UK8LK8hk
aPXP2K32BRl9KYSULwjBGxw7+iHhHsZotGQY5c6ozbOGe5LrH7oz2wk+QcHo94ju+fyk5ZhwMuoH
T6RkdLZlMiK+0MCkA7CUNPg9lLtlRAb4n+ALzg6e2N6iFAew582HBEy1fQePkJQkJ/zVc1azPhfi
bpcZpy2ZkaEldosY0LVs1HmCWORZgUjgZH2ZnfJ5B93m51OOB/y9vm800r8Dt9nY00wFvTHIP4RR
atvcMM9yfA1/KSbDa2TZdOd8SNyMxZF453PfWXMfVyKilxrx4In2scR9AH1Q/ugOgSqSoefZ2vlE
k+L6yuYQss74olHxcDGNNPHZh6Y0RAVJe8Ie5LOCNh40MvLiJULc7M8Apl4CGMC152OJEgOp1iGN
jm7x/aBSI6TaemW8bilzJShRb/WkfbE2h2Xw31l9LCHXbvg6Op44TR1Ykau2pLKuN12+EDQkzJvm
3TBTsucu1h4MHfLoKdd1Q+S405I0kzY9fVRJ/W6+Do+6K+Ro1ZJAlV6ajdXkHJSy9+i3v4FPkIlH
6TCm4FKbVA4vWMlHyZj/3i4mHyfksN95HmtFRztrLV4/jw1YisNMpEcVGFlYjvW+i4r7LKpoL5rU
CIjCzAcsINvkeIg6GtxUA/S/E5fSG7+bFNLEAcjDWCyKLCdfra4XztjJ3cm5vIY0DpOE1fATKPlR
oOrIefbWnV4OxMrw9bA0B5UzgAsPnKuYdj0eM5hjXlTVrH3RXzjRyrJxeYPOUiV7Gsd7xPy7OCv3
KOSVdV+hncv3NBm6dSnGX7lFJqrI6puVcn12bV4zUv/GvFwfi3Bh9brqP7aWGgt+CpeU6OCSb5Xu
/JOTv9jL+fCyYe0RPUTpIeyic9BWhdHGb+mB/OX+BW816A7IEiYLy9kJjM1ifea2TufT8p74IyAj
mtxmWFFgpCH1FKKg2jyd0Fo9u5y/jC/9DrzJ5bcpi32QmOZGh/ONjdLuxtb+gX08vmNJyAE65EEG
U2vRMeDuZIiuXC0LrV35QYKe+9d1d62XtTNQ45bh6fcJl1P04DEW5w90WPHkO45bSvng1PRXT3wD
61yOFgl/vcjmdv8CN+goGOm+i6E2Q6mvEjKUH3wMb/AMw0WDgUwNjQRIMmoK+9WDobMO9MZM06nn
59m01t36tWJRXkdjIPdYHORFQS2AigmLpaxmyTXCj0RtchXHtLD9060dyJ67MedGnlY4s2ymyLqy
I0Y65r/qGiIcIXzmI9r+yn3wKCzKVQqFzQOe63tsfrrqS88qkxIZ5P5v8JJJJUDqX9puPo8IQVXM
RjRmbaPkMlc4RATZvmUgW5gYMUX5ffs5fXDWAH+3Drz3go8w1fr7ajtk116aCcdhyj+DT2BTn9mH
b173aAkG9YWIAunSppT8nU8n14HYCDieGH3En4ztP3/aOUqAUTdfCo3UQM8uXs871rC91KJGkQJC
7Dw7mNCkO+lwLIcsuuRoH+TDzimZFyhPpazJ3rkZHOifVNIVlfMGHq2B9IovMm8zIDw5B4iJkoey
Ivx7DERyIv17zA4ejFVgcAe/eD3FNtETdKcvQ48gGRAggB3xnHAaqgcH0ltICRCbEfLkSnzslctv
J6w9K/QSzmpZIC6XeL4+b+waqtxcRcvvWa6UtjmOC0ztAKbSmnekEEb4Oh3hq0C2oucX21qadjcX
fWTTaGKhK+U9qVGnW7TH/ytL+3m3Kjc4C2hnHsylY8rJ/K3tp7yIFsxNFBiTz7Pi7RVFuAFXfbE+
r6oBLwAfTXShBRvYiKYvwnTt+/OUtSJdyyGOcLbp532T4q9LlDEtLTxQGjWIBFgeAvI0l9hye3MI
qsEt5AQ11eYHvbBBFjdCpFIp9jmnx+z+v2c9Ypg7XqGVJbt5mzWa1jtG0I+cPI+UF+irtSVZS4wd
/8axo6uyiR95er8isN8R1oaYiGbwleUVC0pxg05WwjLYnDHJzwq5nhM6X+zMsnJ0qdUDL9aSTQIa
HcNqyULiiMPiwnV/OQjEnfHISE0rEC1W8LIniCuC1rwtwLsBvh2ndNy4E9mCkBP4IHGBt+lDJGd3
1VCYKygHBXPzUFXc3Bpn26z2kqbPR1XrCTo+2x2sHofnHPt+IQlLO3OAnYa0DueELoHJjnwPf8wY
vrcyBk8x8bT3bxo359vX0i9JiM1fOgnGAEmrVjypn1rJpi7C9WAU+HaKxiTwOrwClHQSyGO6jDfg
DMrBqx4/i11BA4HX4X7haPX4X04RL0w7nhVdNJeEa9zKBVv7E5Y1rUj52C909ZGmcPGbDlMJOncf
GuHRv7OklOxbrhxROUBeSHjwwNdAJ14wn5BSzj6Io57QlMcI4FxDejYtQ8DC/Uqz7Gjik3scZKt7
spqInBUp8gPY03wcLzMM2wD9onQVz0uaSesjrcqLJazdgoV7SHFG0odg7biDfKdmWxXwxc2mu8IY
m/qskFg3a0ocIbGe6GrHuXDZOR+PoIcpjMg9l9buSaSipDPFB8IVgifB7HFh7OCEaYYl9kk8kFJx
5lI61XCk8wfuNFQfUHSoJhp/DpKFet5l5rIM3E5jEAWCsqMl/mbSPX4OVhdbkGrg6mBhqI3NhQ3c
+ZD5VpXqXXqIZl/2M3P141uC1+R+dX+8/fNbx+oDnpv17fz2AhiO+tMggpBK7ZRsnCHlgRFxHW1N
x2uWR8XrzgZwtxayebwCmOiGB3xPCHcgG/PxwPXFPXeQngB0QpJNzmNv+6ZfzyXE2Ltlst3UqaEQ
TyOiOuPz/5GGnDUk+HU3k8iBjJNgTs5TAQVW9KI6zUizYDFBu/wRwp7CYnM8a/ZxDpRUVDPF0vyQ
ih81Q0FpxaY3TyxDuGPkXPBmmX4lWyPO+fKq35aipC08c9c8seTKVFfX+aiCMSYoWt36IKDjXvbd
d6aumNhOz6WmRZzbiWSlfb/qE71NUp1L+Z58AvdZMIlHWnqAK21408zFlaJUwd0Aq9QL+mn2RO9e
AADHPbDueksCLcGkw0A+jEzh3ox6NXRTbh8kytEsXOH1ukoksXc97ZMkTmjLSZ9YkjdrUAqkA3Mc
OwkPWVomWHtvcZ9eLV9iXit2TGeYsN5gq2gSUSD7d1X6WVZP62bgOl0CUZj3WQbNE9otc/1BBDuS
5dwSG1kQ2Qy7PF7Ux3QZya2hHg6NwmhhJtk1B/bfjOutITw12rezA+GGe+F8VyazQUsuMMH1OTzq
yFDmeovtH8nKKXq3EZc1INRkIGfQOjkHm1TEOTUT+6GlitxZwniHvpz+klV1WhO/OK9j8esWv+t7
vX65q1cqAF5c2l/yvK9tDfJTDT9P4mCwIp9bIHgJZKe2Jh6izlfxLkR6HM19U2AU20LTVTcMghUR
8Rsc8Mh/XxfN7+IFohAIHxeyWclzB8l6sLW6KI259QJP498ve0fOxu+vJML7QYpM/MvLLRfeJQas
SSHLO0hJ9vMjc7PTfOG4pdvcemo9Cw18x/kkAhVjSFEQK3Gq/CQ7LNX7RzCBOHqI47QG0KPmQs1/
c3s4CRRixpNILogHeV2pwcEDEGq5UaAcVvnpwQSfEhcNZDl1MiWUFq477r5T3VB5gT2LrgA7/Xgw
u7z1BzHBKH3OIwuDS9g5NXSRKWK7Bp5Du8yh3WlTbT3Od5AZjYVxqbQTBnlnx8tcAHJHcJQJDx9e
y8hOS8AHWFJ1aMGUUSus3pl5nehe1SVJgJyWEhY84gOxTPOhQjqi1n94hBGh6wSmWxOLHeQx3AuE
yUSoaUxFOdHvndloSkh4S/mmZBybJXHsfPEmaQTPedXaM4Q1SicxSCBo8wTp2YH12Wc1MgGANx3r
5ABYkHS4Iam6IkC1vxBv9FD49na/ZS5ncwQuDMGJbEiAEs7c49grg3KWnjarReMujPR/Vt1c4Hdw
hNHmE5fJRRhn+eybs63KL8esBIaFLekyjyDz5itaDvAbHcUVTQZhVO91jRcLgo2yzJ2BHDSGNutu
Frv8cHvX1iyVeQzblu9trFzdDYGL29KdDLiesflErws9tuGYDFnfalZT+NesF+jT7Vc9I0IWsW8v
GOkX3cNZ1KGlBOUPQ9O/M6x7Ffis0zClk5wCa5b2OyzVE7h6oyCPakByVVhHRipyOg0Da/xANxjB
cAS49UWIw0shEzAheyxdIco8bwn5EYtsDJrZMBmvAWQDnovvznqAglxRwrgNQ7348ofbqBfi3Ilq
JIpmFs8PCCRQrEh1wR6il8ZDXkqqxvVcxrSg8SzTRIYzfnikEPVlMvy6I/gBbYp0Slmsg0rvOeYZ
i2Yic26s9mqKJTLMSeIcp8/tS3vkwFeKzl4GLeh/9MIW1VAO6MIFSbpX7UOH/zY5rusXKNrpopGh
4V60WJzlk7l+GLntk2QHkJKReOd5Tl/QkoSaCpFEWDmRXva6BBNtPJuTRINVGcvUnyknFCPagVdj
wxyYOgkhanwn4fxePZYbJyDt8sTr96vf1nS0lA0hVTAw+mbhZR0xWPxZ5CdXP0R4gTpx3lT5iHN9
W5z586Ao/s/Oz/bG6qggi/H4V/7aWhdLk+xMDuf92dUX39FE82Q+IRNML3xRGlDgBp7rFtZj+Vpm
kk/oz1fdlCdTAyr50O6D6R1gc29YrrQoJbBJd/T6oQlGTxnr9JG71XbQhrFKLhEAbCemGyWCrGjy
GwQ/3NQ0GQN7Ygt1GzzgOFti5hc4LdO6aG189vAM0vSdoZIOUypwN1sB56GhCmIc7Sos1spYzujd
MvgXTloz4q4jF+WwmNRkrU+74Bk8cgTiKDCFfjeh2gMoFLOK6tDl8MN1iB4UnZ3pxrRWcFbEbID3
OrUqtD/j6lNq5VFHcH+yCyizcqZNFsJ3YckdFF4GS7KWmHaPn5RexgEboly/BmDQWoLyp1HhyOQ+
iiovwZk45fXw+lo15wap9JlqVWc0Bkd2Ps02PP6Lf73HDBw40voYGONpMIa3D4sIidjQ+cDGdHqX
Cj0rEyxVg/0lBnGiYRBkdkARLjY6RZSyrlYBNiIPxGqCMti2YsexQT6xR1+YLJACZI2ARE/Bz+a6
tTkPdMaM0Q8MYhlb0eEiLUwLw91PLELz7gWacCSbuoWq5y6SuI48F0Mkco3qSLxqW8o2gKi+IyZk
gw67msk0JUOjy8VvHEljZKeICaUdU8QPm3ABa/4rTdDzTYMqAkNPONODbEW81D/8nj9P+8/02F/5
bPlw1S7uQaUFaax3yn2f8AYOlm6RXuf40JY89vN4Nnv2vyFLagEPKoVdsmxvFDVrG+MuhbWqBQuz
wKvc0O3x3r4BoQ8x8FI/PWffjIMqZtljEwezIcXazPzUkdoGVQxb9e+4KW1+hAkUum9x6ZXNOEPK
VeOywX/5Bj5xqoXM5KJgB2QFUNmug7OnTWGXKZJR9ILwCanE7Rjfqjv0Oxh+rgWvyNfMej0fIwxz
2vn7OWZSwEWSegQmwjE//w18Ol3zlSABIn7lUbjkQpMokRBUieT47squpyqIUgt4aFptgDjPBpvO
mOBb6Nvw6gr3nOgRmjTm94p82z/jazzSQwTv5IVeBOgYxqf/Hmw3hoW5D1cutym0W8jBs1S00C56
3gl5qOSX+WlD7Fw72Ivk9/YxEOu2C0ShIT3/JCpakjsAyaqUWfmH6PsC54QH6M3UmRHfMTtw81Gb
ZAXiGvTyhGG4KklmDbD4j+7/l/ssxbsA4G/SrwpeQCzhBM5XIAG2iqfy6nLB8sdR1A5FD7gzqkrJ
aYok+BsMTptnZ+oE9vRvtf9gRZnZ+IdFgLlwOPqrnZMagdUIUm7nJlStMMomR6JdipA20wg6JfqF
iS5Z+qr1k1U3ZqY0Ry+aYvQ1M1qwgkcecDda0lOYNo9oWBgRJx/SUYmlY5gVkjIsUmD4huuHhgfg
p5eDt2Xvxf4tjqGzZ7rZOZ9eWf06vR8Mz6BepNw+inVc/bW5KmixiMIst+r7neZFv/Fqg/263FdM
Sw6tLihcrD2S+uh8r2qqYV/BPG7kf6k9j2CQgO/5eUhKh7Abs13R0Zs/1TrYarLeYfwUR696uzCH
gEmBnEJMcoSrQ0Nua96LALv2FjwUFJY5yq6j8G2p5FAp5mhLmU7m2DG6Zy0jJR2H12aSE374R+FA
G3c6fHHNlEdv3e1Bk/UsFI9uBjfjOnRzlCC7b9zB3HEt8wXEjQhBjYzhAAZ3O0FL8EZRuMIwBauF
WR23Gw3XOf6Cq9pbCMJu+XVJhT9RVP/xwxCw3kRiyR/qUcJUxOJH1eCtwKsLx01Hn84dE3R6SNaf
egSnSQIwujwTGXv+lpN6wgyzef+hEsh2e1tu7wskklMQp2KX4g6M2Nn/KN6UsfoZowsa5uv6s5TZ
28CScydBovlioq2ZApe9DGBzrGRONKWqrrZH7B6Kcgre+z7xtxuRPCYNyU3eW32o+BhLOQLYe2n0
CAJHVbmTmoilgSG75uxuPCLz46kWtngPTTDtX38J3D5yzbOg//ABeHr7Mwh6Wkf/19+CZ19P1DpO
3zvaFbLkCVCneqkuoGdpzzJiiQwsCDb57fPMewm5ERIlNFZ68B/JOCjaz3p5CPqMj45+wpjjqvgk
xVT2R0YoenmKtmI3nmsrjrKknK9sYcvzu/N7C//960HRRS/Efs97OlE7eMjKCLQwt+aEtVcskiMD
DjX02fJLi7KwrNr1i03I/g74i/9W41Xh4TySdlVBZpfZ6GVdWDXCsrvTyEpo/q7mMNd1C1vI/ES5
dgkZEqnbjnGZkeuRellU7PkXROD78wStvDUJvWaIi+g3d6mo4V0mRLRWCNxgD+JH5gSHx/gcYUYt
zKeRd4qb2H40ovfbDXxprE1pA1X68evvAQmBdQ3FMbTIPRrYaG084Y3DvJLB8iAeb9xMgF5Tn/72
vsiLJ49o2xz2zx0aWBb8/k4wm6wCL54f7r80g5Mzs9FCVEa0vQCrOT+ufenLdwAZolPmdMHM2L/E
QSY+c6JReqYgymGmmGmqQ6Dlqp+tGhFhYknqj5TQk7yeQotXH3MzGaTAUxOiMdB1DC6uNgO98u/C
TK/xx41Sk0BpOyfFiGQ3tIj7qcfvwoKXMopA7YV8NYsIiSK9spV/WNvf8vfrbcMJ24MVR28o0Lgn
IYXWUzMvkrD63g98/0wJindyZzPH39tIY07fGKqPop8yFdUEiTIxRlaTlPs/CtrsL/UO0ggrX2/N
ref4elBJZ+bHAgeP3Exc/GodIqKJnohd4GbvEujenFQo7i5QlXnclFzWyuEQYprmFOndtqNVHG3f
u5FChU7Jj46mgF7sUKA6H9qSreC1dOGM5pPbhUXKu6EuOtjMACmzrTYNDegxx9aDmMXpfnPaZJyR
djJ1s+c8GfSCUynFov7A3Woye594H7k4a0k4d2quCTDHArNyVfG9I3Z4+8z4mJaD00bN4U/uL/Ac
2P4127t/aFnCiFmErsgV93GnuvF1ETP5OBAM/n8t8a6cdKD66DndLXf5wR62NxCvgj78bPim1Iy0
jASs/vCc+IdmnbQFZboCOAPjYcX40NLbJ66PAnN1owk5HdYI3iZ2FZnBCJAlVX1gtYTdDgTbLk5z
bMJIQ4N5b0uJgSGHBygBEMFdhIaAW2OK/CGlvWD7AhjJOmT1x9hZNAwqzp8DLLUFiKeOsaJt3omq
t5QZiQXgcGwTezxlP61Asz6Zaic4vr9mI4O7F1dKtYjZJ2A20ihqk6y6hbY0CxZXJ8/dpUTSZoW3
4cBb5A9oU8MoSCqP4WRcTu+XJfuyQmUhFjL0vbpcKws8Sxj8SpIT6vSJdm4wLYUyK9ET0bAzQHM6
nIb8hCqvrEywbZ0D7VuE6/1yIuTnbea9yPJLoobBqdsZVKLK+6MAcBLVLQFkV9L1XTm/r5Mfgq58
6T9TxQWwsKLhrmup/3IF+nhC5ifLoyxgCxVzZjjl3as5Rpj7QGHKMOysYrvct30fGhsNHnT7bj22
HIdX/dOHt49nk3hBT81QPao57ZRSt8NrikvGlbg73g4C/N+b/jQyxBx/9xGPWkMJGquK/f31Xbp2
VufCtoEQgSCHe1fxnQH/xRC/V/G7SPM4H9dqzBlyPEnEPwxv/VfH61FPxI8VKGfTxeOjARKEjvHl
EYFusEoDUtPj/8G0PJJtzmfaYrnPQBgL1Qjgs6p2SKpU17inNiKJ9Dg9frnjDYNXTGF7HTUX9FNK
5QAawEwhzBE+7uy/9rmTzMDGo3OpR/C75mJAIqXl4aujSA05VkFEBSdXV+jpaR6aHsme4jAceLvf
Dtjd7NGXIsqAq1aGZKmVYLrC719MbaYDmy6HZe4upFTXzHJEger8/0P4fIrgPMBgeTcratBP3hoy
prWQOhBRFaCBkrNLwjJ8DAEhw3hFM27GZWXjd4FoNEYp14VrCBpM8c9NehHUGZFMazfI8TJnaOFN
pqvv7Xbessm3Ro/rYs/irULlJN3l6CPLbWKRLCylF2xmQeVtRz/rvp9I41UCV81lcO1SOMMKygZh
j/T2USw7a5WysJ99pDniMdr2t0CJclmmeedlS0EmY/Jdj6Z3Yi9jhhOeOvtTLxZ2wNkQzFDVWBFF
b/1lX78x4mR7PF/aybXNTXKrzX8ypJUBN7PQjxin5gP3eyeCTEj40qzmSyhm7elQsH37otcceZaa
SEH/hOOsV2FkG6KYRLENtBGMx/EDkyloqh2GI4juxWSj55L5+xxwQuJedEBvet46pS+F+Nch46Tv
PKyj+VaUSBgRG9S+BL2t7+mMQsqHiLgCBBnig/jCt6I+cIypAQkOASEoN9kz+mFjs9vNMWkXJVVm
vBttj6WXlNrMnAZstNCKp88T93ftLbpehUq4AAK7T5iaAgA0RCTuTR7lLOlDkP4wkF0cce9kYOpa
JXweMcb35jkSW1dIVBVQIjpgavkHwXU3YT+vqR8T0SrBqJ3tH9I9pY/CcB2/XNizuNUrv+c2JUj2
ey1x5OhygbfP98qatXVF766AiKYIiWPMW9MXF9rCfkLz9AI8IPYyr0aeuuOm9ZSlJRhfwT2CEXNM
yI/5eeEP+wmGy5+i9HJuUd/lViXfwYUFyp6iv2qVy8yU0o4iskCdzMr/0VyS9v4YuQHbrLq3krF2
jMdUYQt51mUE9p0QCnr1dqpYV0OQjqWtzams/jhXVjlWAudmKX29xFLrd4gZhBln6ak3H6MVGFLv
hwrVVc8RXnC4zzLpt6rwa5IqqZoMnuX7HDKc2one0REeHSm6x9NSImyKek9KhWt1Dj7SX2+S9UIX
uKxHZftWex1fXElrL1hYWOq7DiJyhjQ1MIdF7LwRGG2hnyWBgxGL3maG1/5z458idIF+xcHB5HMd
sjVi7nqzkYDj8tQXZv//V+UzJiQYwcayLfO7x84Ju4rpnlJGHlSdRVzGWKxMbgmvIYZVxBP1XPIV
5+IivTWOHmQQHErJMHd8KRFKTYWjOApBTqKVckzgZfkZkpuLH/XBbZjTPYY0NMWt06ZfJKeH02CW
3Exy4O32c7wDVTMI0i7FnsZOkGIBbdaUx4AoqEsa3+wJ3606n/B1bjQCFMv/4UAieWQrrYgaWbWA
8vnC61oyY/KY7BFAiVPEXk4oK4pAd+6bkum0HO260GNmaSlhb+C11Ecv3r1+vl/qDj4E9DMjKyT8
3+Q+cigsaSksPUM7eA9BMrUA1YuQzZBsjCkMacfbeCyR5a5DM/zAdw9nqF6fd4hoH/egxMLlNsMZ
OoNGkYkOD2eJhZvUconCNwuYcl99htMu0/0QdvVmI0a1hT8xskonyzfIFRRi5Ni9fpxzt7CFoSdy
Hx1bF8PCNglrSTo3PvxiDXu+UWv2rJaWZFrNiclkU/YWQ178s1UXHbChTE/stDMQ3FkSYhqHJu5o
V20wfNTA+SuVFpIgocN/xIyM3TOH/rs2BXAynLS89+4b/17aw6d3xc6sdukvZhHokTSlnGemt5m4
8fCp6UhCd9fy9oUvaiJS96pCORxH38Vdo+cqlGgiS2gthyLuPct5nZ/bzj5g5BVgrrqIhj0wSLvU
Ym2pYZ8oROL4rTsCq1Iu4BjlD21Dq/EzAq/WomW8y47Fw0xNhT544bNYITc3jISoIO9g5TVeH/lM
d0dnK2SHaS5TFZKxdDWrbr+PRm0YcRdMi90fO7WOaq3T6OalgBmTFzndxxDHx6zIjY3FOK8CCtjF
Tf+CsshcaLSbLPtvenAacKKfJ2uqsOto56f5WeFMb++9aNiIGwgPctZWB7x/V4tCl/GSSU55XJFz
ljpeImuQXSiFrKEuMKfpJa2SqIaBLrqKdXrsA7CoXpr0WYnYPgqOUXz40K64MCTb3EFgPxSUNWVh
6OlOb8/XQ+CrMeuOOrPmMUB4ubZZ1jJ+paeXbOU2mYxCwywQdVNunmpnErWN9UyUf781ZicCEFa9
jFS2rdtPycCA9z17A+uSxHDbukcQRfzMH34exSaUYWJpkJta7vhVVCwfn5YnvrXCVeB90tSSChGm
wzoSwgJ53ShnzJO7qkMSt2dmNUnIsNk/bjobq5rAkzsOWhUXQ2PeoGQZZLU3o7pKOgchQ4exEBfR
GAkQ1+YzYk0lCvwu+wmMiah6hUODZ91afg5NhEYOuupDdmRN3z4BBODhDIYAM3nC8pGOYi7VuYMc
ozyqRc1J9pLu/rzzS8KWAPZiu6L+EiHmtujzDrdki4f5EWeEBMAPgtIb9F3W5ooQ4FCVu0Kpz2p+
3EWfRM5lpvnqWXnn4e5HrNwKfLWkmZmADzzNatM4U6N+GVU164s/w0682VZZU5GBxEwYCkYlq2y8
W/IMZ94m+fknOxMiQ/NogmAyH7NXurEq1EwZWZOuGPtjw4rIGfKNSgvvh5lDy0n8GklPoH9XD4Wj
+jJC8Z8a/oMBTUS0CvrdMhLCb5thOS2LpP9xcv1LyNF+KJMlbyXyAfJ3fLj9A3kHxCJF+XC6+qcn
KpK+r220s7jg0heAkFOirmkI5api91+K6U2SYA3PBX45FMVNct/F9N2aadSgnyRD6aqG2Y4rcYF/
ZmNptfAZCDpjhkWNVnB9TVQWu3eu7D3dfA1vYZNG+h2oRJhGe3l/rgqHVi2xgk/iCcO3EBJAWdQG
4dL+ju583dACtOlML/nQR5wdTrtzYrKnlGEMTP5CiL5h/N18/kNr9xBig1VrXTjaIHua5gJS5Num
EE4/Nd9/K5koFGj29MTwg8DAX76/Il1R2tu6GpxEOyufNXyGFfrFiGNm2C9+BTRDURI/2PXvPpnb
Ld6af7G1BXg0H345g0E0RNZBM4ZO+9H8/qPqMq0bHxZI6+1c6pYWnmx1ZysJMiA+2OG+1OkuodgE
ZVno+Jcx1PHBrvLcEfX8OFdzfE1NzJhItgpUHx/ypj3pJL/+TIUi+WAq4m2v69TMeeQHe2+9PFQ4
iRe57vxz1HGgNnAprxeAwBZqhpHJmveL53bgXGbOiEtlWiHuoG98q5Uh6y1JEjd9SoQo5oyBfsQB
prIchggrIJc/yP27pFevJ7nhtTmp7sm2+FLqEdYtV9IHMBB2/iS6NCG2f0PrES7U5apZEtlB6iMA
q17YUFpcBrA+z7Oz5FVyLT6vg0g+wzAtGNG8nGRmrsNFC9VEZHzen0t/U3xgD/zC82Q2jHD53HOK
IEhSTUj3RJb3DgTnp3i1lrojhoa3DWTkwAxjK+CEUba8+ZmssGuis9CIIT92M9uW9NIlItHfD3pt
dOyj+LpSKNNE9XIZkQ0NQuiSoW8aCVmrUhGcdaWUeR4kZvhvazAQra9nTeZ68YehExjvVefXtVPo
0BnIVf+LxJV68sIXkj3lbhRu/2Fvkev5DRCRHa77zgRPQCYe7ZfQC7PtH+UH0X7xG9zDihpRj89A
j3KdtRnIZSy3yQMBM/TZSXsNBWi95tikUBlFH4eMn42hJlR1xnIukjdxWjIEMQ+YcMiLv09yJ8G7
bczt0rFB38q8sqbwoe+3QrRJMbzpK1ncwwQJbupNKA2OoVEg14pcupNaVnZLdze8Grj0A9cRe+fE
nSTxkvowxJgaz76YmtaJ7UKcgl/AcsgGo+eExPdpdjmuxxEr4oK61vx1Hf5elOhVujYk1DzdYA5d
hPhhsCRT2dD17t3s9TH0NoAVEUj+wyj09R+FEJuN6ULaXiHaE5KxCgGsvx9eqgq+AFQ092dLLHOw
e4UEGYurOFn/ExUUDGb6MOrknlCtwC5mwUqs3is6FRaQCwYwdLvbHLer8sFUlsyJyTlO9KBe2RrV
a1H9sXuSNUuHZV+Cz4b7BsWM2w7tOA3Sb14xIL6myV7rqI5ewofL7/xWn2GRuGzHK8Vtik1OdXu/
0bR+Rz6euXe4Pg3Pg97z0hqZJd71uK1/IiRn7SkodjY6OIKOwIfLgdWmuWXb7St9VHLrsKa88Yv4
Fr8W8i/vPINt4wTID7H0V5W9tTqngtqoUcPGNYolDHoDG8UQRFuyhbhdjHYs5i088CbtnCsVq5qw
vZZ3OqTa/M4PDrrMFmYixVSMvGxMVKbWZl3fC/JS1rTA52EwhUaqqg81zXU8c2TEgbqujw0ZzH+D
CrdgDCl5PDGQY2sFm8+BS6ls4dC080kW5xGd+3wQgrTvznubUF3p/CrUbO0/WykkUSGF/j0U6t1Q
YcM76QA9JfFlKMMp9VbHc48/sF20e+OmQUCQRl24ttNlezvwO/1fP2BkQftxbxq4f+b5hPn78b9J
qvALvNXijayTvoMw94Xm00xVpNRK9d0SgoqoZJ+Jf2+Ea1MmxowNmekafwISu5XDFBtuAlipXeWB
i6QHnWtu4C/0BncEUW1e2UmjhY6nQ2KVoDYSmWauQC+Emw96tb+2SgGI2dS7ENFJJCsJosZVmw6a
wm5CnTJKggIFYT8WdyMOU2ik5rpBIXNWC4ShQulnvkSoz4Q2Ysfrf6yw0N+ih3a6ZuSQSr5kDf8o
FAdIIIvq8tB9erxSayhlYANbM3ai2F1BHgbVyiezEHHpRXBlHEJU6utxbtIN+dVVeF7hXC2nc2E8
7+62KFiyowAuDq2srmcqXidq8Xqfl5SnbdORhy+IgUZFk2AV/tYGCNi07zaGmdhXnrQ6ZDbIJFuf
iOxJX/Bggz2d5YUdIOj2cyV+eqIBX2QdeIvwky/BQ5goag7Jb5mh8yuchmSyuty/N4PELj4F1Yy7
KF9LXFge89ytXJsHe4rpYP2Lmmo/QkRiawGBGUS4cWecMTc9FCMwH2D0RDGc44SO9iYKdr6GyHs1
u1VBiu5BAC4Ok03xnZJGNqGkDEEIeIifEZOJpV+TYJNGJ+wv5Hkkw6kY0ThtrxwvFtzt+hjcMJns
BZ7GBdjO8zmxq3PrRLLlDtvkpZ7gvAv+s95jJcdyYEf6JDbop3M3OsbjQnKU0jucBk+KhJzS+j1W
UgjLbTLOMvJjFkaGh7lwtWQy2FgbN35edeTA7bz84V41pQ57ZnFQaVZQoisDKP8ty3yPUOSlMxix
IAabcCxjrEJX8FNcv5bsvgkONCCn7a3H1p/d0a4orP8tx1RJDjdHtbIA6kplFMzAUbjDxOmWMnHF
uEe0aCTKKhmfSFnRrBzbu32mAL0FerSVkW8GXO/xVsDKiywTA4zCXal97reR57l3OxhXsX+P79c+
hb3eD6rYuFpQl/+1R2NFf3JtrC+CK7Z4z8buwjtBo8/Agpm2AzDgKe9WUqt8ArfQJAQamMHdl87n
t7UXNM9lwxn6sZcMrjihs7o5gnndlPG4Lzp2/PMG85Yx+Yo+6dJCPqaXOSmqrTvhrempAOQrN9kj
amlwlTiuugeP5JtO0aphhxNzy4DFDYsmekrVNpILMxN2G1MALkBlWNtWDbfVIdBX090SMBfhqosX
ior/u/nOCNJnbMe0ZiTAZ1bLiQROeqBIuNDBd/5HhJrS/3G1YpTT7N6Uc2V+mQozgMGCZHwyqjjq
Y7sWT7xZcc08FhwYWA36vELXdbj8k/XcwD/eaRvufBY9yv0Tj4EO75pHmBLTwRz9+Qi5QRNBUsmn
yhE+ptb3Lb8N/UqgIx6IENOVXxGbpilPb16TseZKNTvxyg1EEfiHkZH63oNvpsXjfiP2S/+CAGPt
LYJVlXbXpJdZ7aEw15+Cw/JLbbWiSTy+oXeYE2ae+n8CGptxK34ZC0DLeb9TuWgGNhWWJ9pkNkuy
SMYz5HsJpKlE8nrTk9y9IgN54n8u5HcrA+fOAzds8i8T8TEWCkEGLEMmcx6S3Xk0/9gKBYBR2EdZ
1v4JOkswiOxC5m1UFLSlYPyNJaOF6UHFtkXveLIRfyQmRFhQfh6mO/tMdyHDDYxTw5yiY7vtm3pA
LFcNOTxb1txaelVsYQakbVBdirRJs+Vpm1CxrIZAXfHAmfjGYnnEB1s/MFca1HQLv1ea638odPBu
wTFdxXe/MNqU6yldqd6tyz01ZrB3yeWjMF9SLjaTJghcm5x6/F9x58cjFGxqr2S+7TBjQ+2zbpVA
+RtDHMbjgEHJUOQnDxZrmH6CP6bD29uDMRtjuhjpJD+k2DjbeMzNdtWPECAVL3gQfxUm5lkceKpY
NC+81jB8kX0e/ciD9G1molvy2qLk4XozajskNDOEqRHXWCOp/7wLMJbxqB4ThjDfmulaVs/SO3/L
ArFw+SSnoQgUkM7/NQH7x36bAsf/fHLpiYX4tGENQs5Abzzv2y665S5UOR7aqimtYvr1lm6RjzKr
SxX0C77p3XNe3DkcnK3jnl2rddi1AG8MrMR0c79lEMrUo2Pd3u6ALpqyhuroNmgyhaocKDzMvxJW
+lXHi74fdDkjCeLiEAq0YHpw6xAaclXKC9UqV3KEktgAUE2bJnbDaLvgwac9ilLs0Utbj4nNNr+3
kd2Ckr9x7VDuyAaKWqd3LdKd5o01mSdbN/tFGe/mJDhjzm+l+i2dE6soo30YseghUBHX/m5UwyUD
bcTGhi4BV1hcIX/Mvm+h2Ri4RpFRnkVOYbFdcUHjs1E4g1GDaYMwpX6fX47s2s+yT8fvxhxjzlHd
A77e8vx3tNAazDCFpLh3dFJkDjhyanYIv4MMOVw0HmgTlA8ii4rmX2DtKg9xGWWHDnZeWuXJl3iQ
5P+JlewCif99XitkTyYz0T4DqtWmHxzC40vWBH4qxZtx5hQIYYybS7ir982VWJOsidoUuMph6enk
R3/I9/hTUaWjxGjrYxceN914+HCiaMGyAzdvJo7b+FeGUTWKcigQhakQywfrZ4/lTQ1UgaWI2lvz
jus9ldIUOGEQF8m6rYpJETrKvPwKkO1rUHxCX/zAU4zdJVwoSURsH+baUxw8lSihOvajPYWwAmbY
YWOinTwEbF4ChyzHzBtml6YSqhcAHNhlFhQkxhxcyta3PDy0bIyYkQgJFQOfpq+mDUWTVlvYGCUN
KOaxZFBT5gPzrQAdA/IeaWmQ6b37o/1MlPHaBCdmlW1kaPDxpYtm1c4JFavqpXv6kylD906frXM4
43oBRTmL6YHxlUX1oS6CYiKL6TYG10lJt4rCSt8ostDzuo7eGKWkjRH56L/L7PpgueP09358CGg0
zZuCv5YSDtczSPsDxbqiLoTWvbkmrSVXkw1ej3Y1aoy/Vv604if4m14IRlTeY64WugiqtCHiOwxD
DygMgAg7yiRL6qj8VLoJ2npqlGm+LhK+5QnKtuA2yiYiWeDT8brkanfd9wLetanpQzdxsNrP9L/V
1eiZzYFULas5S/CiGaiZsICbEv30T9iey+hbZaYGpVPzZ/RroXOpodH+LSx8syiyEAvcs2mScRRv
+tIfrRxX2h+ygjczcxnYGLfKvFm+5odYDnpe36Txc/TuGbkUED5Ozgi5ecWcw9BSfMoW2AHWY4tP
81vskv3zL1lr175pcr1CI4e7NcbRAYsZlQz6x/Q76ttSylo/dGH43QvaoFkEaO6tiHle8UhxGkMm
dNztVnSfLVXlGhUXokBhr5IBsld6KD0tOxfIft7q1qI6QPpRtRTYS0bWZqdG4XPdFe9CU0LAumtq
+UBuCRb72w8V5hWi3WVW3U1LXC4gjEmixby4B9SvZkBG1Is+4vMLeHf12Os4EkTOcLmk72IWnnM8
jR/csA9DpW6ui0h5YRUpXyykzVusvWv1Ry+MkTwc2jvCx15NgItjhA/F+LepH84JymRK9gTTqlE3
ZTN88TkquiofqAwpO1ArOGeoy/agZE6ApSY775Iq7H4R3iMs74kQXF2AxNmOeGOgaGcvySChO43K
oyvOCLhSzBV/vz/K+A2csdJ6ff50tRTa7wjmNW3RIZZZFQrU3cD3uJdgyKwbWu7K76HA/piZmCcf
dtP2WfnxEcj9vWeJnWTBFGRX1LkF+jhtZ/vAt9HntIsGivcsEuhhnNF3150KX9SABG4esZPbVy3h
YqDIjN7RmfF/S2BY5y6hc0onvnv1Lyh3eRfjaL8q6nFcOTrJavwzoMj1eagLHSd+w8Ja73rYci6y
Oqsu8HY9PM0PR3DJNRahxxHI0fvRcJr+ukk6Od5lbjEM+YFGYUhpkV6Guh2Sqtu1us/j4cAShIs1
SOFfdAIlrKpnaCLIc1Hdy50KUHXKpCSVWQMAZ8fK+LZyG8/7xf0cN5RZekKN1cg2DNEINGZbSy05
6S2HXg9aHevLm1pSPYs5gAYeDfZhhkyJkTLkSXCMupXKihnS6UFs/fsehATbALWRDuFxXr/8CRxA
vC4VSTwhrGiCyjQ4AmwPd4uXi+ovGMiiKE61Yrdj3a0WrBdHIsVOx1KBDkhqbr8v7lUzxPK2UHQC
4PUcRjuXwxircPyymzgS6JlnGcVijtO9hHYYtcVW4eI3XYTh76pD/sdeRi3ZYmpLyxyYuAoGqYCh
2YyHHrh79YLhcMi6usBFKKvTLrcO6rGjup7dcf6O5bt2zMsPPs5P3UVGehulsEK8mMM+fEGhBv6L
4PEzNW4y/args9uhVBwyz/kwGJrEjuVe/+Oi9+haaA61InGadEAGIuKc3mq5MbHnNDQ+/EF7ZMvS
rDHexyFXm96kDwvS2bLV6Mjigzt4H8ra+elmmQ1biw9zKSuSAqPAactMFjMygxmnUOmpdezoGtij
jHoJUZ7NjRjLL1Wr92Y305lsfuZL8jJ0YQwM53x7JisVMfM92SImLTuGofOUKqkJP1qvM1yrr+9c
J2R425A8BwHZeEN3WqQffHn9j2gzadRWPpeqjOIJ6lgqKeipoZ3DEKvbwD5M8XXwdnq6T8cg1I0C
JoWcAXGgHsbBTXh1kpNxjWcMSeUm7qUJ7WZOvBdMKUMmFc35V+KpZqbhEG5j3qlF+iGwKZGCM3v1
J/IXTM6GltN1G8cZMSXveYbpkU95ktJblk4MT2n12p+RAyXlBZVKiVoHqBecc+9GtsdTRc4DokXd
08ClS+xTHfu5d7uQHedQQS0c38d8ZqEbwujQxaTQDIz/SGiONcQwx5zaKsYseYC73fXeW/InpkLY
yvvQ2qvOyaniWL0EuFyFpACZHBYjd0R8TU0OJ+13DvO1NWYh3nPSDHPFH8phQgFSzUwN021ITYav
AS9i+o6rwPT6XrVcQrDyZdU+HP4OyivpQyznl8rBUeAFQXTq2aO3dlIoVXs4a1X2XjIW8oIkOFTP
D/tGX+lvSE9XWLuD+/w9R0bLLUD0zmqLCR1tKz0HWUJRJ8Dkgcq8QGa2ny2kCszWTbq8H2g130/n
ImZcxGGkj8EcXTxBPFW+gQJ4GzQL+N53xs5u5chVsyKBytGWlnnAqGVSRVl2vmDbK46+RXYJ4V7V
9Qv0h0KAJMFkP4cHbJINU/l2wK18tpBVjrrtToiN0aJCRJGa1QMlRAGLJ7Vzs3cv69NOZ+emeuHy
Z2hU2m0LxkLN5jRa1EUXXNqYC+aOfxN4WdcYBnsLb9zk1wV7aYiRyjSKdssTVsUDCEUtB+6kIhGt
ABkY9jJV/EMvU3G7devlQumXIZoSGpGVNRmw526hWlhQei2vHrVV9Mnw7TlXavwJntwrkJOVQ4/O
dsEjk4T3QM44uSl1KLWmCvHYEuZs5iKYb2x4XVPvVQjDluY6J7ZrrnNqLp8aGFG9UHRwh8n4gpmo
bk9ef/AiyLlva9aDcBgeh4ZD71xMOuONMf7nfvFhnAmi6vSTeCSSd+bGtxpCEJ7ijva0Rlumdi4h
qya/f4QkDOCgYpIUIhRpVbKSKVWH6qWBr7G9/7OHGCHeWkVZjwOnlm8TAQV1kvmb4RC2O+DF1aY3
6iraVqWzsml6z3mLV2LaROTJDLBztLuQa2FjC1eK/mXAPAXRt0k1bvHor1YokmPNFYV6QmZahK6M
9nghOkvjfBKu1kWZfnAeuA770ISQQuha9xK5YUBXZ0rGCAp17bk+dCz86Iu874vfJVGbTxcR8aRD
9GCKInqvfzJ3KHJLcYHZ3Knkf/glxKj2U1ifYch3ixHlPiDqVtxXHtHyygdlty8pnRK/Va8rfrNM
Ib7Je8279fdXZiqEa+dhug6FZbSJsEE7TGks22AmfVoK0B0HhjTUOLn8MnJvnOhj1veibskxyrJi
7CWTD8kX/qiqmkK6YeA6ieLbLtzCsMg14+FtqLG07ZEaN/B3GhUwd4fQA8RYQLdecisdYuSgCCpK
LkWZXsEAiGOVzSYQn6fLfygSPTzXbB2bLBUCWOp64zbCXXN+xDTf6wbk1g2z0oFeY2PbPP66gSGX
AF95sVl7fb6qBoXoUrWWBNv8GeBT6vftIGuL4KOwtFSQI6fiLgn+R8BUZiHduJEI378mub1Gu+QQ
9J2dSpfOkxnh080sWle/rDQ/MyX6wKZuJHjkjuy4ge+O2RMcGw5e3IsWXaxDY6MSKcdu+v7w1ZdQ
NvniA8GXPkWo6uDyR/qSb+jQi+L8TUyvghcK/hO7DDs5N0WJGp4JYYs9M4vFxOEEK7R5Lr+Qos8s
LhqLXmb9t/FKRginv+KvfUejGPH540hUmvFSIt3oSQjnA6kzwGB8YqGoSETXqcvgKUFeK9YBILOu
/3W3q+8LHc2Td9nBTGKMACMKoQVnGEMFjurNVFLXBye5F7pX7Flm2Mfq+pM2KmaeyPI+l68lUmWY
B1Jh/GWd2zltltSWQkUE/GdMjxJ3XyRMM98vDxX9WYdcNkSeVjlUuP2Xz9QhpoCAYFYh4q+2jagw
x8kSJMkHHLOSHOh3D8iLCywB5khqNluY6Drw3EbjpC2fwjXPn93rImUrbXgWMZufhaEt3DqT6+t0
w6P3hm38MNd+rJE4gDmg+vl6Sh6TUPf0Zr5ZAiFG2cO+heWu2GvV+Be8HdYeGZOshBh4b1VQkITs
7tP1QAsrKgCAw2My1C7mx/eZtv7PYDDz426jHx6nEGUlobZodQtKRUaUbKMXREN1wGuhqF8JD5v7
/O2rGsuvTEpJ9Acx1acEk70qF46a32EylxHyjSlpr0l3HXjSwe9iqxFg5JzYahcu8amacbqibX7V
+SIG8aiukcEFPc4/hgJl7S4227LWoad517eD8aLM+ky6c4DeAK5BNVGlGbLGcj77e9nkp7v7APIM
Qp3IkJ02CJuT9KdLQP1f44/T+YQpcgdUJ+DRmMOhUGjeQVJATTQ44hX4qeI+lvLcTTIa6v1h0po6
xx8iwUFCHlXpjKoWpbn/VLkuHVAYHG+Rpm5EMGJ1YzmQ5RmW+CHF2fOBnzgmUlHEG/fDfiuQT9QU
9Ny9v5h6Ap59bO+DYDgl2R+KBjuetN3QHMEAEjjZuVlfUB0GwF+PGlWd6NdmPN9VO0T92icCT3Gs
c8tHD6Wk7im8tK9/WIqz5ntSOz16sEoAFzg5aG1qomQtb6nbm5DFzORfhom/flzLwLUUhShe7HP5
Og4I4miyV9FKj03OBie0R+TnzIEhKqiYOiq64EhS3VimIpvHWOoNoWnkx8kXi787I8nhTWbhVmQ9
rH/jlXLCZTuLhkVPqJcJ/+U47StgXultV56763KK4+q1ygXALMSEMKZTRuy0za+3NKAY7QZIxjlr
VrY6hJkzjEuHiS4tCOJpe6SST1//pSqX+MkwfSzI4ytY+0iDQca0NtWoxwKPkYMFSFACMl/3W7Q2
eQpqLP/zDo0RYzUibJJJB1jNpH6UbSZ39dgKBORLuYccUrvU6+RkeUYGDSrLfV9w8GV0/wr+KTE3
dVfM270owyLl+IQPiAq4v/IVNqmknilOKQ3S1obSpd424E7tFYeSm2s+ex5Kr77JT8p+xZSuyB26
exuclhxZDJDJlqNEpsBp4aiPmj9VGMidcIzXH45P13T3Lj26B0AYzFEsVOlGJkZpkwg+a38vyRrd
QBkASZ6mJYUb2hZDmcmYV6ie36xn5MALfCwKvCxyKDGNC9vXeKJWJ7e/HuKfx4TJMw5/Z8ae48cc
EEBFKPrhvJ+kxIPxCXrv0yQwIzQbtHdKty//Q058fD5JTdwhb+uWqGtLcR0hWpBigl2Uha39pI4O
25QSo3XlnZZKKcHxvUWsTuSmx24TsqHYv5PWeMDvzEzo9VbUFhlU5zumPD1oKIEjpNMmiz39IJ3G
VT11UJB/I7S8ff3R0CclodLvfLu4+c/QZNWojJcUU6MdkMm3bs5FXscFHvmpH69aUWaBhQ+Zk8hq
kMoisGZJxJYBQcWPg/bKRW3oDc3/xZQZWZkuUyrHIHMwHHm6vbJi+J6jkqDWOjs3Aj5HZXYtENgV
otuPtPtMPlhl62dyaG5S4oNF93ECcwgpRoVhtPCm10E8/qSMblmubDi0KLS7yZ5PElAQlLHknDDx
4SBr0nPaXqp1cv24ycLKDvu8Fja3iKzC9Tehsu+DEkMP4g+mk7UGCqLT/febgdcrJWB3FrNvdJAM
e+ZDwmUOzHyLtHlFgVmNP8YTOTnDrrkoUEdYH9ya3yaWdRsRFRqIxXq2fmcN3W+hSz3uIS81wFA6
W7mDXLnY9c7G0JOUdq/7oTQUs2l3SPd7z9PFCMbV0z5VQs5Hgl761oK+f0B0AE8AWcDByxv2Dvr0
ZPGgqeROsD2E9jjxnKsm0HY9gHt9VLeXANxRo+fqmDeUz1QP9Iq8ZZ7zdgD7DD7JvqgjEevUAQlm
lirO9p1Ijt1KoCW4Vywy0l3cQllVWAmuXIFFx7gwmsf8sL5P5pDSCF16C4Jk2uZTivUaZFN7vg7l
3APig3Qg1vIlZZeHvTB0rE66i0eFCSuKY2G/x3ahmEfXgO2Qv+diqYijRCiJQkKGkzw37QtYf4/X
NTJKV6SXeD/Ye13r5e8avUIARXOe/I2smSVDEnwltlT3qmI0QgZJNAoW42oy9qZzU3Zx9ZKlXGfG
ljZcdS0pdkhHAoHLoZWLxpL8e97RicXEg1AUFUIJql6dK9NstZGZOI4PwcmeiLzyUyKw2Yx/21FJ
4KTp60EQS2w3BhNS4iANtWmrc9BFD7vWU32paKfx32RMsZO+/Ojbm9XHHbnTltTcNQZS+7FLtc9I
iehEZg/cvUASJ2XTf9rsxbkHDU/fO86V6V283vFgDdx5ZrZhNs8BuU2I5UgfniIbSALE/aEkQRxH
4yh18uluQx8gAaXea4SsoenpaRmptOizzeMeOskuIAKNqxKT4qLVvsgfhP4QaxOsdYmti5CydHMy
4PxYnhLKV3nJDsTB3x128HWqDIbnPbwy4lb3qiCB/PuIIMBzl2UQNXJKwvDFEhTKpSibS5RbOqSM
SShto/q7rt2nvTL18l+ZYli3RV3Zq+441u6gYJ4YYh1wZoDdDYMN/LD6qxR4xIvgvz3C9LQlPArl
mdBFarGndJ/q1s6CgQTtKFEjy3TO2WiMcfh8WsHXz0uA5P1WTRhvflumV48PHzPN3vWrv2oLeQMH
q5iM/mmpWUMyqrOCPUKLjkX+AKSd+As8hmqLdqQx9ONrmK2rxpn10LUUkDYKLinTIZGd3KnaIFwy
LQvV+BX2EgvTTtlSod7Lf0MTH1tENvJwCUchCzEWa+8FhdvIbsRoS+96HA3puzHuBMDJKs8SKhG6
m7LrXnu4MRFOf+4fGZNukNwMFnUnDtc39Sm+ih2g7+fPQ+IamLbWLWFTd2NpV8qEI1ns2hLNt7t7
Yt1zVI78LXxCtbqdURfvBRjXzxEm7NXPtH+N0q1y2nBrlL0akMewY6yXpbSAXkRTwi9SzMLIw1zx
g1pSfUiwYjAliE0CmfBNJLUApn79z+NwesPqPVi+JUex4PLEW4vvsmWwY0lTIZ/zPPeEKv6WKQkt
P7qVo78wIKZD15zivKcppPt6JBWFlf2+rKURnXGlqoyWUgY+No8HB/Cpn9X9bqu9jQ6NAx2uLSKT
AcsKkiwJu/zy/cVs4PwldfU+k5Hnzv/1T20y6orRXJL9AKmdqmVkxKErttq5gYgk0pDdBl0J9P4X
NzdmiCZsSr9ygNchwVb1odBTh1EoH1NkR772jbHg1Q9OWVxHthYtJFwW+5TJCwHm2Dtu9XvotuTw
NUxT7awwultFFWmWacCd6PNb/ERB96o04WfOTPRUi3EyRwvMWbUuXBVxo+JQgwmuyLW0U+VCL9CD
31X+LcpAgPb7BLuWXMKmnPqEMTv7u2z0LNeIvR3w6DQqVtCRZY14CFQDkay4L2+gDyOKXbpsFc7X
BdKY+qD+HkRBzeYJd6IV8Yz2ViJYJrO8a/S3z9bDGLxQnWi6k0q0sx7Sbp1cQfBxPqXQl4Lg6AIA
d73TiFYbRBWG59ak9Vat91H2xoaHzYquAC4LxXl/Nb9I2+sA7hM8i1oEp6KsDXQxSX/ux6vpanWM
7MKOW2+CvNsMXL9nA4ZD7KFqy3j8QNSZgazb93HfjQugrXTkC78Omh8LG020ykuHmdZz9O+7Hn24
0lrDotrxV+6xdEV3e2zik1kAwbpG535QTpYrtHBljxJNhBGkx7mePeRTilRpjbENQGXVp7G7SUoq
gAbODYqEi+CMpsYaNhIGFWpBEgVIG6CS+QgeQ7lBKCpF0mYXvGLWaiJ8SgoOUEd2T+oMyLoSmNUJ
P0J4EyGYutgUcoVGSs2FmxvwMy9wJAXabTNY4IxqR+0yz/jPGZmqMiXdLUYBpxlQuNYyoZkEKwnZ
Cws2YuA2XnUnqVVDOhlCUTVP4bnBZI2lj2bIiFF9p2ZR7+69g0iXVJZo33aze/cgG9L9sydLhgsq
EimGSVbGleP4MvXS7h52Y8XLZ1Cn6Br5iZiFMyAbvYhBmVac1Mo6hVx4d17o62e2/fHxfiJB7EG1
pXvH74XtEGVNrDocEQpDqj3W9qucTBkBVWOlEp7wSL7rJ51OnCZvDbR2QKB0dqfCpBtYoo+PB7nJ
8IqsFHKoLUkXP8jSHPdN1nD0K38lNyqUd16EI5mR07YnyHz5UBoDivYaY3Y1FEgLyqlqTHqLYEiw
61pT5aCgf6DQBMarVuQBtx5zsg8gqWcIrms912RlrVcL3e8wTTjupD08orYbVU1AbtLZpZQUv66N
vFgvi9blqSV4HB7gIHae5rQWVy9Reqruv9y2c8LfWzLWhogRzELhyryLSISmDpq8ds2u23QKtcH/
XM3lQx69hR1AcO8WEx3ONbzn1gJOKbJeF25cBSIFUV1LiwwalwwK3h+Uj8QPBq20z+/zmu6ccyOP
gLVb703lj7KvK3DJj/RMnppqJoj8nnRMB6WuQMRgTG2VH8Mpzt+04R7+33ReP6vSw6g33XaosOlX
HHTDKOwZiasTHwFd3dtQa+zbYQeWd2x5qXYkFYVV+TXETAK5Q+iK8xNInEUup3MLW9s7WDANPG7L
MCmmWVTntdD9tpwn6cioad9hApFPU40yR6lZpn4ev6c9Cl3REAon+dkI8urdpaZUe1zS3CnfDVvv
SStSYHBbR8szLSmwoofQv2bot5mLGSNblZ9+RcQzn4j36n5xHW7CzVZNAOUd0hBM6zlt5mXRZXPu
gO7PEVvngm2DlQ5iWqOUCZS4HKbhpyMh+RA//tAFV2dCHA/L1n9HrRCICt4aBNYGAq1d3UZRhH8t
RBaQTQgtcPQfh7KQJod+Jqo0tTQYMzKJQT3WbwV8FlZCzjeiilmyTDNtz4A6PHhgue9ZzNHn0bqD
8Uu6M8VFN1IjiVq8aufT/plbnVXAnAhXnpAicgHUoMaZTjHC6eQz/HJhNM0bQNCU22xm6l2ESN0x
sjO1JbLy1NUEFJWekUDzEXHWv54RSr2LaSHdjqubHdy3RFKHNhGHSz/PtTOfVJhqGxwlDPlxbf/l
LyidL7A118Kcqr06jZaPXb0FJ5n0owgBifzpPoHtceQoKr+cIeEwRjB0LdqdrtBG5n/VxLmp4D4r
1qJCAURPizRkh63/E0LRTjYgi/r3C2UEysvtUCmX0C0sK8TWWx9iA1zh3J2Cxbwu7Xg41QlqzFNW
MNrAAzknEWNz4TquIjPlatv7hVz7lcAFTs9/FDfoKxw1paNcxYjpsCd0fWcOcG9qgp0jzmsgMI/T
dlmzlQuk5ruCEUUgcKtQqUpx1SDdmADvrx+xplHCxbNTvArHDrklD1iYmEU7ecumsvIP/c54j6hG
w1LjUh1UemWGJcdeZBnMU882qbRtgII8ftNSt/dnizvAXFhsuzElwsNL8xqpl8p3d0yHwBDEwOJM
+rQME+1z0mhuMwvf67W31IBGHGroAJCCJGVFTwstsacCY4Blg8USXu0eElRTBTj9j/rzAFK5Ug7O
DhlQdVnGC2OMmPh6wCJF9h1IZeE/nsFr5CYnasUjdXcJ9Wo6oXXTztkm8ddXggD+B3WgFHB5GjH7
ZO6+K+MPbs1DcrheVOcEiKO6oHBMPnVGmiquYv1ec5ZL2eOYYu2rR2YV36ecMdxtQe9iXZHvNi9J
YmP4dmVLlcbOIxNbHdW8tJkjIBt5oiSWEdLgHR0j05biYkYMqvKOMgxCHQ70J7MjOfZQZUM8UbCI
t8c6p50V3O9gaVe5sxoQAsjoKIcwzSXL8wCVCIe/h74fuAGB3TxvtWoQmA83Jbq4WuatT3j6YM8l
GeUh/QhLEZvRP4IrcHOTOeNp7xIR3G72TTnxf/ClDgK0PHHCF8XRbmsPtN+KhbbV8LoPlat+eAmM
R//h8J1x1ay6/65uDkefaXMzB7RcPkDMteaJSQoNc3e0H3YSSkEKFM3o9u0bguD6fXMKN3r05XUG
1i1fTtRTQ3RqMxIZMxOPvrHLJH03YZJTqYdzqbR9ykFL2jgGI3VeXhLVz8jGoPVV4X1KCczozm7U
GXfG/Kweg9VUeB4XWgdQh2H7rePIWUGM/j7tcA6CNeYlBe8ikmJ5/pbJC/lto9ioRc1cPmsAgV8X
emJkc/eTCex3FU2mxK72dC4sBtmISpEQfKL0hRWdBLeNzvwX8yMlibczzy5e6pnUBigrD9GenwJF
AJiGh9IUI7ACrLjVJyL07K1crPiegE1Sq3n/plQ9FQSS/9pX8IFo7zTbRnBEWPfyIngTvbjG17yD
lfX4FM4vH0OsCmZb7b4A9+fsX90m5x3kmj2s1051tO70FtVBfD5Rvh5x1sPVFV64dq3OV05U7oBc
R61g7mAOMloe4RTivx+ihWOWETEx23uh+wq7vBn0KgomWnqPTZ6u5SqJ3zjPtJENTGUm9I4EXDJH
Z873IlLuIdVKCb5G9c4x7n9Q2xPhrvsgE1axo8Q7ZufmYPDweMyqaprn3UgreixjhLx/Q3BZu5Sw
ixF5Tfeem4YlcuhdwIjqGe9UEjFC2DFQl2MCyNLNiw4k4nu1Spp+nnyL63qlWNB2X3JsqNmZtKku
a38ZpqxE7wR4Y3N4t3hxf3/wnE1oa6mDS6NrkspwTp+HxSoIBp91HrIQtiro5FjBEJttwhWLuIGY
zY5JGt+ciCckmEHMzFnoppqHr4KWrWbKVsi1/taWNu85jSq2OkFK5+HzTQ/N0zbgvztLavlI1TH/
9RHLhaK+DfmxY1zNOUPdJdUGrHmAQm5MrxcG85NY+bxzwLv6B24ARFbwsskjb4BvxlApLO2eJMW3
9OMWxtkeezrPZI1jgXdHsm5rg8/VKxKTGb0TzYRZjk/Ir6YCdodix9CyfdfwNaDwjEQLqkxDzrjV
8/6T83fFby3EQU/FFSF9Gjya+GLFRgPzNjLVHF5CxtTSGn+zjm2sDWCHCEN8V5aof7NEP9jrrlWk
TSUKm+JUTjfYqgou2lNhfkL4Qi3RVYkNJ0iEQ8ixfpJ299LyVJEfZWXsLk9D4aNQNeLC5AG815vK
bDdOeRodUZGkNUsUtjcJJbqy1jzYNHYT7AWV0Kbkn1hyMMtNpHpDZ1jt8MxghK0WZJooUM5Qh/jE
r11bpEXykrHHTW0GTvb6/QxxpgmfNZomi4uBXgqRCK39TJSQqVwb/oJ5/YTPDtvMRjCBJQlKSrxB
q2Cj1i1LAOL+AeJi1RCtVVQn/YwUIZ68UAHG7F7mb45JHNs+jDeiHvw0DYcmxaWo1/i7gHaSqGVG
VOvlN4nWWkIo+P5OrepThfOMSjX7TqCoVwkctJCVgmthwfkXuR3ImCNAgLB73bwMR+qpKOREN2yl
zj1/QFfv94BBls8isK2QiyPJuuLwuSp8ovv+590ij9zCx4OPYXerDrL0wUlXwfEhm5cO9SPwkc7k
kuFHqrfOLhh2IKjPlM4LOxG2R4RHSXPbNzvXivds6e9V+qV4gK2LyVXdGvwJVBqGASfXXPQzFGb8
9+G/NAEkTCtIdcQGp1NewdgliuVhDiD/XkrbDJTA/mOfKPERBHpMDW4ysCFNc6AyirnbrsB2SdmL
eF62piiCMce7iyOlQhRGaze6PLZKddboGD51WYgK/CyfqJFkEkGZCUk7TSxBFZjopsepO99xBNwP
t34ZE+vybHi4V87Dtr8KI+Liq6sbQVeEvXnyuEzw/4K0ZRHtzjCQ85T/s5dU0Rgaz/wnieFx+93I
ypf+CvI6vLiT+GH11fzZmi4dTfn+wc3K3C4hscb4vrh4eS/7XT/9mFufA8xbdfaFg5+HhV4vfxs+
RjvUl45SlnwQEjxHNm9tPGbl7qib8A/40b1cwt83ThHswgPkxhZanerj5fzAJnuUsfcBhDVNv0Kf
gq2eiecVBugokIWQbJjiR3Na+w/NkE9rDfiR1hUsJg0HrsF9x2VicE/09O+EBu1P6VokF/71BR1c
mIfy6sg6Hrf75BDE8iRb9FgeNuNh9DIpd3k6czKlbw4clXQ6sHPjfvHIg1GH4iLMeVaztTeumyTD
prcJ4IT4JM+m9TvHYjUvtnIT7V6rw5bEiEV4r0m7XW4ttdAyYnmAVE7Iv3m8/Vld0E0bm+VhHrMT
Pe6U8nXZ7r940DzII7Uy7EAMk5dITrTCT/52egjHPeqTlUSTRRhaoBv2BDn12+SFeVEGsYJnNjqs
v15/iNI0bR54T6RvG/9XbWhEmKWDJW679yIymhQG4kmwJyWlt2UPXZIe21aZZ4c9W2/Vc2w5zOOW
KzFdfvwJtWfGqSCPL5gYN8QW5ztde7vwBXWGJkmfGJC3X5V14KaV9npmfOglhXwhjJL/sCYR/MIU
8yOMbVNWmF8eBPUle/eM6ACaLdNMolJMsdRCKCyZoj5OW2SPf+LtIihe1mi+6Rpmx5e67iSuRvSs
ARCMK1xLFDtwnfWL8KxjP2s00/SyVXtBVUPZ24Ys4sYK18L2FZXQfRFGHF5X7vKNcfGmF8kHsNtI
M8aVnReVU3s3JdyHW+rDxEmh+gdNGRv713hafoFNPJ9g5XJVauR45hqiZhSDqQJ8t8YnDNZursWu
ZVK/NPRkUuc0vkObFmu86aY1fXEhdw8qeryyTjEd5V9Ts+n9U6UZDuu70mNcMRmMjnjZ1awqxLqH
33KGqJsCzAbSFAgz426WK6rQIi8sX17zAyncaEQzTkonmJK6YYdtQKlLn6qD+MKg8T3ay16PcAMb
eBd5GEEfe1UQocG98a3UIPE1s/Gkq4/qobceqqibmljUiuLYyslYoHbfYSMfs0qbPvBBwb76IdNn
LXb5Bc8N7LKVM/PSsgevP92oOsCHJIOV2qP/2q6fv/7Qpbi9xIUqJlUrwoHalnIracsyuwnnS1CC
Edm/uS2FgvBOH9EX4O3pqanFuL1SzqLGRIOWuRnpCI6kLasE6k4rWuqZMIWBDofdxRMz3hKMb0N5
DEJFVo9KZWLu6+dcv2cNkn3CEQsDj8wp06aNr/g/jp0P5a0koGOKhdpWRi8iwAneuasRa8Xpn/a+
VL8vuBpdqz8v/n/PVGwB2kiEF4wjavLW9571syBOpTa6a4xmbwS6gNYOw/nwNy/Oto4qAp9Tsmj3
epoB4fyyrwWUBRoyarA1m2kguKAaYGl09gmWnzGYfbWTKoLTnaK5zKZoydA67qAA7E0zzitC0oO3
MCu5l0t4Ndel18iKXPWEPTRDswCmxOFgOo1Nmh9VvjwLzqRBwm0Y2aiqCSimBuVdOGCfmNw6USLG
3B4ETY/q+1Cec7YTTLe3IJ36CxRCxg2FNmmtaL1w7oX3HYjmUhNdcddyVbQifoYZE2sf3QZaJze0
CMCF4F/RHLTZb5KNZp55g9yzu1D0R/BW5qOnMxChFCRAjWWNndPwMHYNZhu1fweCFbMRMATR9dgW
iQ7ChUw7QNZEjfc+yxQ5aV1OO7R7ZWxhV4e/gnOZfYgEnajJMZRG2Cbfd6HLWbbDmH2h/3u/MgWq
LHQ2hjR2RU4klGq5GS89UV5kUMxYAQO/Wo4BWhrCvjSFu1CUcUfXd7ZXD6OEe+JvkAZ61xfXnQC5
YwZrKg9p0WaKWSiHYPtc2YjA9F1ckTGjvmiV9cRVZS9cIUrK5PJqxdAgt8C8tDbgH1pNS1kfywg4
ScgisQaW/3Z0lHRZBFZekqRLjuXYXDLumUbajdmy2Zru+Z6MRtU54wGq7l3OK6ERsxKiVf8ovTF2
6QlFGio0LD4N9Ay3rEc0sdOWxt07guzviXEuqjsgLqxh7XftfwfwikreWDXN6aU7rPy6BnYUeNNn
TfGX8HKIU/1R23y6WuTodnsiU5HY3Xt5zmi7cU0ygtQ4JDJUAX+w96HbWORSJrngBC0taxUGqH7Q
TQU4wSyNVaGoJeWp9MYq/JlHZFbB0MfboQJZI9Ws5CP4QMZTRc/DPecwrVG44xjs2XrFsO34Gjq7
wkXZfREaMFHAFOwoIL9YKC1CDDFGwjKQomf6vPIIBjZ3b+NIUkgRchytElvJ2UBaw7q3c5r8VX8F
HfbFVUK4HuYTdZ3kQmPsIkw74i+AR+9d7rfXFefS7xnLlyyaPy5fds/n0VyFUOyFP1rOTaCVp4K9
hwHTyv+fYMwuKS5CQlCwjChBouhIohXwmmrDCvMJ85emdOi3428+qe/AMPlvyK1k00t4xgxpG6t3
omBblxbb3ybBJVOG/aneUEKohdXsWL6TdePMHh5zfzESIbKPp6Bc3pEt1oA7fxxGIPnc/YFFYh5t
rhYLrQzSXEUfOLpWiuRGmV9domdZNGqIyIALBczmyBA0AgLqxPjA8q1/XeQ0ubQzSrWSoffZlfNw
4NMxdmSHGicQCAxlMc3JlhKUZMG9WTMoZV74ct5RnqEG0Ih/Q+WPg2h8geIxIN/QAt4+Fgri10RS
Tb5kY3juKeQFzox8STSyp32PfmC/IQT/6OeqZSbv/n06sRPXLsP0Ga4dICACkHln0FN2EDaQJ32k
h6bo1NWs8b6TPr8cYw8DOOqlR296jIrZ0e7GUCjodx8aK35s6fKKIKlpBR5fBlq8uhsE8TND0HxD
9sHGRaagMDeSnzbNzoPmEuMguXeh7jOmcApk6jJ98rhYt8OP2qJQjcm8ZtP5MiNC8Ey5OyebUBr+
H06SPGciX7uCcUNZoNdwGujiTaEzwAF1OZKL1MrqV2NsjTUguSiKAeQzQHrKG25np6LperpsMEl+
ds0j5MR+pIv3SDUHnRdwpJ1UIyi2rDCa2KGhrKQf2B9tajpG0imUFjbLRlOLBMGFkLenkQcXFi9e
Foeey9EJe45/AXHNnNKgm9HUXTxcaD8XaQRvV2eQm+Wozam2BP6LPez6SDd6j3SI1yi309826OBg
w05GaWY+dEcXiw/eYBMmxVSvAp3eGm/8s23z+x5vKAfdZ/pUUlFXeQTiHfWAeuNp3Mc6jxZmdt8r
yGsEFYAmqoPTds3GgAnp+RlXuu0k07KD4gCtWBO5Ec5SavFxBDk7N88ZmJg9OMPIrGAAWmdtm+en
L/bQLeJhUVCs/d7VyrYVBvfcEwlSk0pEp9PeWCprxwCe5b/oDD0LWBH/RPWqpBaKLuBK5afzojsi
bIjAxOei072tmJOlpW0a4mZ9bnRqDrg4KEMNfpKDnqOyLA49Dje6GGxgildJm6KZwG7OmqFWQbOa
WR1ezJCeFjIdH0Y4+x+LrnnGxJWUMccKtwcIKiw38LGi+v+7nCSh0bAAgzBYzQeD5fbdiHjG5Hw3
RUL+8VpLSagZbCPzi6FsdihtS/aRlT9GKPALv2IuKPjw5LBr9RjtNz6t/VgPX1wgXhYXXko6Zhx5
3CCzgnLscwu2zZfJ+XY7BQwtO2l0ZXbf5xkBqqEMMmXlxv0BrFujOhp050WwUKoWcj0JMQwuKSZI
LplpLY9Bg4Gj6Kb621tpMitDhdiaHgqsMxqjfLCgcb3b/1WDhrfMAGiUSYBo8bJPltWc6zpq4qNw
KV4LXoH9WDTxBRKBdXHbGDouGhMlZW9Yz1adPuLMnjHVendK/gtkFHpipqhNM+eMU5KUjIkKSbJW
JBEXCWlvVrnWeHuDzWZLUc5R9wzDqLMnNpr03BNVlpRK5OiffoENxauhzBV5U2+PdXuQt7cECN8X
uIayQbOa+xIeXVJUqITgAgSmB9BumYwmow7XaHl+8pmxeNWzVcAfdFKGZ8PpcA80tRDRP4rHx0Ge
QA7mnX5Pr4Yr6whS7heP0VoTF2F1oB6aXdBRwxgP3Fi8P2zym5w+H9vVlyRm2QNBPGj46kW+uVbL
oQS8/JOC7edCda5RyN8pASMPZLHa4kRPHRmNrNGjgOdNG7hrNstaQaP9AW2eFIHrVRkrPA0H6tja
u1I9HXOHTcppLXtXSVSvswWjVaIPe2PDE79Hlbd/uwDONK6mRwiwviusE6OonMuulbxiuEyGMb2z
Y6AvCBH/qCydMDF6W0nt09DoxZqhwqxijgRVZZFoWOZusZ++cwJTi+01A8Ekp59afxXQpa/xKqHt
wjzAhE5Liy9g+EFoHMFe9ttggMHvvh2ai4TdnaJbEoL8LDeXkryLQWmZmJ0HkbEtRvxyqh7ifmvF
TN7x0UBipDRsDaBBFLQeZKWvMBw6DfiNeJeDNRyCnAnimCPSIO3AlUkpPNRvYRrDlPMY5OHJrzfS
/t12uBXoQkElrcLSsIpDBd87dsuAJeWRUcWwycsHMTiD8hNmfjuC70Wo/hhYbQJ96KEHaRDZe4E7
IyyCiqBe5rv5p6yGh7KUFeV333s8nluuA+aD+TNEVeu7TqWPD3U/8lCsbfnCDd2tIbcLvoUZoBdO
qDMuGbsEvnkZTXpoIafC3s0Dlbt9ksP/oJODjJ5NudT/58G1HxbMRPOgKb7wu0HBtKaJmOETbCc0
0dL3aPfAV5e4J2JEz8hPpzXkQcxT76csCwiyfwMNUQAmlieQ87s7xU+VB3teu4c6ozg9C2OjkYQ9
r+GBw2TVjnMJf+Oz2zHarako8+xLqRxHw62IipAOvy66SzzKM8jhm8U2SpmRyG5Q7Y/5TxRgVJ3S
hHqfetPcYJgc9FceM+9KlVR3vELp1z36y5jEoLULZ0vok5HExoHoQEvdK6HQp75HYThET+a7N54v
gq7Yj/vYBMi9jHv+bSia9c51PNC+vItyTgmGtX2JzNZJ+ovZWK/zwqM7O8xRjx4mf8Exc0/OML+6
lQEPx4nYTv8sp1tInMWvQzXQMY2FcxgHgXO3ZciwWCWHJ8VtF5810e767vaLw8bZkkRxgEp8TS3Z
VSIj8Osi5gJ7fhMWEnabcnViSVDFEgy5A1BeOsEWY2kssUmg/oKhiQfwqOiYuhae9RGh7AWjILeZ
3gvvbr/UiBZOLxzebgqIYptnnGhOS5zIhZHwUaFX8aw27i7p8Lq/kmdbXWS5Qssya3EjWUrScC/K
qfdZqKd8hcitQOdGj7dRudL8zA953g2ZN1uBuhU60+ijn9UgC+QQVG3yOUkgL2eTdvJCnCQ1/OrF
YOf/1u4/70pvRA++otuJ8typMoYjq7S3RtGxjjb+997aiGlbJ0cDZe6gNYMPKNyujxxINZs9Q5lS
Hr1Ux0ykOw7CvbFGnAqEGedFP20zaTTjNWXY9peJtnmpxFhfhfw1yx10vDTd7Zehivh3bdP4/gqb
smJpcYEC3iGxvITpmla+fWGpIeknhNuB95iBYZeNuNMA3XR6uX+gUrKbBvMMO/bp5PlR2ktHtkxe
+u55T1ubVG1V1Uv/E1MJZDe9cRXtIJAXivSBcNo+RewRcwwvuHMvhyaPZUaPm4KjdBo6WreYSTWZ
y/ILELSb0w0MX3SWWapS6ZLdVn6siIGQlTzhrwUvfgtGsLpjY/Pc4CLRZclT9yFNzrU06ZKXn/0K
GV+WBV5q3WxXfiZ/e34FUxwfoRxvsTt9usr142Lw5sFi2fB0TDm/lNuLDf0lH/dTaA3Ak40FyhcQ
8zpH5V7s2VHV1gxn5aq4XfpjYUbyGrsiqIWccL9dF8K3Jt6eXfB0aVfkGRWHjFKaEyeg/hL6CT66
hqoJM9wOfkjg5JE7l4TMkoTpeVCsjiiaYLjW7sZLBpBl9/ACmZfAtfU3GT5lqChH1VjJ9/Y3WvVE
Q+BaRCIScFBw6pha7Wb6HdCfizXjG75TfJCV/lPnuCD0G8cNmhzil5k5U2qY3Noam8l9iP7GNTzf
L1b1hQFL9BchoQRB66po6pjM9I0Eauv1Fe9pFJLQ8HjkKUOpJJQzdBXuzlVIuCIuxUxSYcR/7qj7
jhRi0QxTS7Yg+X07u9Ya/of65kvFbhe7CYYwIIiFcQyJu6ph3i0QFYzGLRVuQso6mcSRJ52C6fqR
J81qVP0xQJIdnrIUCD3pzhGiXClFcoeElRKEeMxsZJlMMKRmgYQTUMe5ES0XMkAa3DtZ/tvvFwTy
EgqFq/miNsx3oWOnZIr0LUlowl5rF2Yng28YSNFb8ch1cEPvWei/cqD4mcEmM3jEwx7A/SmkTM+G
B2fq4ONb4My9E6RIECCVqij/hfGHDduIfVGUTFxYzhCXMPgx7j4vcIEVG6GGQ727Yf7/zxodNT+g
5HZWy4nzzaxf0hoZkhpEOWmPF+6S5FkoHVYE59DqnMtbis35JYuQ/hdt5pMPuIJ7VvuFXrrhfPsH
hXIM/eTg79Xtqqfy2Eikf1+Erjc1Y3129GS+RP/Jb/dB0ETJVum5EaMiUmwIxYPLWakLnx3Ob7cy
UoHItAWxNoUttE61zbpSPFMAvq9WbH5R39af9d5Ik/veFdQGiUgeRnTwXIhFx184UGGlh0WiZyn0
HFbrdK9+CpE2CzPYYdfC6OxMnLzNgLFrj4X8jrVXYxz/poN+3X/QQ+a1geMnfNDgNiHsa4EJAkmP
oQytkOCMgILm306r39MytNQQ9NlhFCsYJ84oACcekirpqbEubtXLeFBsazRfs7CSZd9DtyCjnQXO
17P9XBrOE+Z3ITucD4I3kzcvp3y5tvz+vdWB1/to+HtrwQi7oRr72yCAeqtv45qhoa3obyrKL9ZM
gl6WLwXdETM23iH88ig3jOF7vGtky66nTrEN6u4oviMXFjJdihaW9/WRqlwCkEs4sD/5aWofTzf3
MyGKdLawMoYm2w9svREi47MmUAKtnmSBJ8CBnsPbEVCt5z7oxEHsY/FibWG8OqC/2n77eF1lR3AZ
j+AxXc1+4BoVWlHZVoXibE9slF+aRln/8OSY6nedqEuMjl19anjr3uNn41UqSdm7Eig2ZtJ4EZSl
IyykJuhFcFvqODYu0dDlfYQirEXPfawtCZBTaqGfQhRIUdJyZjfwLD7/JAItGFQtrAt9f2oIpnFP
onjkPBjlmvgaweYI5FQab2GhQcj1HKDswkjcpu5qAMBvxrRGxghxw9mceegKQJoXcrDco/QdwXV7
ySgqPYD5QWoQcQZ2NRz7y++3F7ZRRMfvuSr0nbGDkAoWWRuSWboHEIFclOgTZ4uxdBAl3rXBG7de
Xg/8+6vH05IpcdCBFuEMIyyZWOaPj1y6mrLVhs2zXVQjxJgMISAiRVR8SWFdd4Z8Vm46XO/MYUt7
uT8O2IFtTL7Onx6ARl07aLBYIaLB3Yu3mcL7dj+JV8/SCILTl3or0CVcJGdgRqeJZRL+kczXPjxM
wHlQrcEInrC+CnO1KNyxPCQdAOFlAYYuxgjIzOCjme0zDmPWJ/Q72RBAXr+1dirkFTQSlvItXRmY
8EMUrdeGQ1kyjO7aevEbf2Ff+hsuEbIKV5KdusCbRzg8WrBjI2U0prndP7kwN9Ybq0SQUx2Jt/HZ
RoecVIwwK5bVuwtZcNKktwin1+Za/+vuiBHM2ImI3T52T6iRG7CFMl8IC0Qcj/S4E0wKLp/X61Yo
5aVCF43Jkij0ymIVUk8SfEVyYqHTQcSRU+SQY37J8pPQNKOYo5sAFAKfgHavO7eSwC1NRRxeXL7+
VOOuOTwdp0hyzXtIchCPYTYCdB34QGy+wCTBuGrXF/HcQYOeYwcX34z/YXAz4f2NkEE+AH6BsVTN
vEDM2EPz8l3cStXlyv+4JKJehpgX8u+0lh3TuJaDp8r4qjrq/XB5E89RRUkFNtN4fnsYyiRQDa/l
fwmsr2u90K8gnhgySmhfNPFwX+jOFAd2PPlNgnS8vURdQE9zvcY2EXWA5VJnTcSzwla7Y52SiX2s
xlkLoCzG5c1PUdU3nCW2ytTCbDayMDiK/jnjaC7zdYIu1JUotAU5cyUC/aADIZy4h+YsHKoFVv9g
fLIlWia2QIDWcFWvHCYkE+iRe/KvPFuQs3Zs6Pp4RFUF+Ewv9mkqHg5YnF+yPFlBf1u659X4x+yV
XFcIQrVvQd/jbqV0RjeZGI5cqWhuzLjQfCGd9nbNc2RPU0GnrbykzTvOsv73nXRhkL5xVGnhWeZ8
cVSgmiXey7X4dioGlkKb2vdiNm9iLCyLo+GtrUG2ePINmByWHW6nAznmGWL14rt573ZixKOSrcUv
nn0fwEYA/n6i76SSzbUikr/evx/0RmCE/gPi4ZdJ9Y6r9RydK4PPos4yKlFGsHfatlFzJDTO4l5z
qVBn2Wc3241aB0VxTXkxZppYV4DiuyEknt8VH7fD4kLcXjWGCfJsm1fqFRr44hb/QOqblwhUqtqc
vj1kAvEcO2txKgQ8zqOXYWZkmLTl0VUyOnljBnJ/+a1HUsBMTk3pKkA1Gyz5O4Nqk1B+azF1Ftwo
TgzCmESksSfpWpUl/yiGu0BFsCJsz+isqUoEgg1ZvFYeZ/Xn0HjcTDKXKKryFhH/f4MbPd6yG/AK
VB6ykPX8Y+bK9XdmSC7HrQQBCR5E9QQuEMnibXkAA8FDYZXUCMqhphePkVZqjcbPqLQuuUmPXDI3
atnDdruXujye+DHHnJUwGHfjjx1PU0Tdf2saW+RJINYXjySa649+/+v4Mt4vr4LWpH2vZidhbcvy
+W9ux5AX8GApqK5qCMncldOqKNCznnQXutinHH3b2Ae4r82lOPwlzGvLvTGsIh6MyGMy+cXY4iQW
nzhw0lpsAeEN4bvxNJ9OWim5iY1ZQM+l7GMsxyJnEcLzu1lW2WE2rTDIXWMkwZzW1ArG2mNyea2s
vaLXG3R0NwJIzol4bfD/tD3RyLhjW9i4oaXKWcUl4eJnMAvGQ0gOcnOBItkTFsUNikO0O5Sw9U+y
JC0/82PmZRGBm3qIevcC7U9unveN8+Y0YA3Flr3J9Fa7fdnfEnEAr8qX6hIbavHArYmvqxBNRdge
PqehagHe5Acn5JBrqB6Dc6bdQ3dZJVwQ4SKOqH06Dbt9BAitr2M9f/LrFx8DTYQLQuoff5SNZRfk
I2ziySpsfv4CyyFePJKUYUyIvZq4W19iIGsJIjzSCE/kSMKzJQAvr+vOHt0ZEWAVpYo/BVnpXw4h
c3dqAKe4bT+zoT8T6SzTzuMcJIzHpzWa79HIjkGgJOn5wY1lJOh4VOVk+G+bYEOkWEaHRGV2aoVb
ZB+j/FOkircyTeoTTswwbn17TrQDNIZF7rlofiWIYB66nyj/QvVUj7ILXWGOrsLLyLDZAFAq7TDg
1cuf1702L2XsqnFYgTpNypbKWDavs8Hvo5g1ldj4NaNocMLVsRuBMPnKJD2RN/fgYcP2SVXIF1UO
HO+O0MTr3xijdOunxiZHtOpUGbd1wGla+Y4neoyzFWJ5OJKnuqi4keEl6UIxLWd5ELxNB3P2y0Fu
U8Dl0QRBke6OiVIo+3I1CWitGO54+V2KhZqKrh2bKp2uPjWd0t4Nv3/BjmkUo4N9AY/3K/KoB+tV
sCjyb7vcytlyOPXEES6HWs2lc78IOzmx1JTzDyAS0+Kfq713Tp58pL53xIY0hVioC8Y4dvrvH9NO
shtMSiDx/yroVzfoaJLfN4k+JClvWG4j3uhaGFW+63pIJZvHJQEGPbm9jZGPYzpfhrapJlts4r/W
x35oD+jjHothlR+iBLtZRRwPTAt5nRPMZulKEd7l/WYrnorP4coH9W73yU1CfSWHQLyO5K0SeUzO
jWLr+PQ0kTDj/WNyGgllDp+6+I6zuhnsqCAF4dhyuzA85sIZIYG8KimC3vFEmqLN14SmlWyPJB93
2mbJMauEg2FZAb24OehOglfu2WNK7O+kJ3olw4FAHTHzEUU+OoZq+JaveLq6+fmQuq/OYK4gkxjb
P7bJlC1qJnkQu8CTBsxmjy+tg+Fe3P88FKTXdoAxhnxVM/tilTmKXCTgpb8Bqsa/I3e4AiJKnMcH
Hc3Ib4KaGdlGmqdGWS5nGEcXB4IVEoXMVB81+NaDOQtEh5SLgiJYZENn7ebWGr0wSrHPw5MdsZvE
cacXiOtEpxGx9/MZwQyFuou2DpG4PJtV9moLd4XEQikZJNUnv9Tn76U3oYOsENGBxdIzCWJDjawY
xpJ3EHrZDhmXiIrr4Z6zEzz+G+jZpqoTvANmxPlfNYCe+OoYw5ELkG2/kLcNDxgMrQKqWiBFWcDU
ITkEDZGL/f+mePCNqrHLwwSaVStIk9J8Vhpdv7ydyBE1D6ZSZbgqCl6EcVS46fBYEA2SdR3XSJng
uYRbB/FwZsP3X/+85uMFM8RWuisZXcwRfl2atDf09H9sOTjQcsBUDGYdlI6Ul9OcvaEDLm7h4PUz
pP4z5lBmLwBRWRBTVt01AT/xXxL2GsAsAzFuJ3k+pZIFsxdTeBSRUzd8KNQ/lY/rCWXwEbTOVnLm
0n0+nYWyT2A6REPyU37LxRfSg4F4fRKhNkyiBF6oqBNV01XFwMwZLT7dHyN7zY0zcbiRkiqGKtnI
2YZZ5EwD19BfTSVL1HwG4aq6Y0dVKf1DaHTtpTviyKBis30lJIqR8goNxgZcIgRc96lkWzk/PiaV
aL4hjIKWDM5ytF35S6Trk0vAbIAU4HppBB2T8wXj3RGSvHgnJLWCGoX9dy7NcYN8lpYUxayZ34Mx
qpT0kvGJ4RGhZNiDMQw7HkxghVHBdiY5AAzyjZTG5Wo/wVfxoanf++hTROeTh1mxRiswM2SEqpXu
IIdlvLIRgyFDuIIUWbtbJiiTOI1EHg62p7/FGIQOUMcrXeD7WGIl+YZSiyqWku7X2KDd83JktJuJ
ICNIE1VcoAyXoMeZB1Kv3UN8BZRupxZDwMfLJGloO1Vof3a176w1iys4kilyIzmyvtDTKLyzv25/
8LXWGZm00L4L2MT0VlxZTscz/6o1Ny9Ba3knUUK6QKvNvu3L2es8f7iK4yMW0BipOYmqUt6TtQKF
1/9cx0okKDDMBmRupj5AMVYWz2Ni/jqdCsCuzgaKXSMhOfik5glP4e3CKRMqs/SMg+qUHvYNDkPK
J940GDavlzkUbX045bQlDu5TEdLK0d3vrlU6iDeAyQyXn0mSpLGjPF75qTfEUUnipDI5xpqaIupk
Bd6bgLeRBjMTZJoSMFZdNi1mXSP2BrvdlNi1XlSJDx/Gs2hynAuy5mgNako6jXoo2BIvDsCcTNGr
NBjRi62ZCYWpAGQP2UG+fnVa1f02twiJqVMOqucv9l3ZMDFCFHMtqMY+fqVJHUNurFKZpMSGSczN
KReI7M/yLGXh50iZu7efhChDQOdr0RIxE4YD5NB2N3XeqMYgNbghTze5aMZ5ttVmFOb9v0GfzbPS
+oHb/h7YK67VA5YuAFTUHv2IeYWNElf6qfpJXVXi/9HvjK2yCqSE5g4AKzOYA0V5I26SZNe9118b
yumKqLUHQ+EKvo2o6i6XErt+YOhyAKHdhgyS6h/OKpZKL+qsa3EZQ825/9KKrIpDapiGSc+e7GMJ
WTYzNKDOIcMeqaV+wysFPgeXyBEvuR6aZhvtbyQIVS6R1vo8RKqHHCuZkm0FJk3/oU18ixkQKoV7
+Z70YD3DsRnwffGW0zSUAThmeO5CTL6trVwvxeC6zdjkeSrRG4M+hZMcd8XW4P9+59IJOMy+rQXW
ail9Q+YMiIbMjeKcDnXhrPl0CWzIAeSGLI59IOxgHReHsDSTd6BHqd9FlGTB1vmR+UoULljUmhNu
JukfyIaIUz8JxSqYgYzdph3XJ583w+UwRJxJa/+FnY9uuDIOOT6TvW2Iv+w67jlT1+ifJL+i7WoD
87GpYo31pOGIbwz+5vJMGOF4+0yKI3zCYK8eRGhHYeJggXrnb43EnbIQ4zib5Ai+PL9zYDE/nhoU
ZvK0T8Vp69bvBwurgvsi4o8uihgxLjewIMv59e5g/5ILKPvgD/5aADEeX2VA41/mY2DuvFEbftJt
chMzIqFV1tMntdJL/dnZtjpTQq/RCVBu/QO8cIHMDG4bLsGs6u1YWd/3GmIG/Ht4vqOW2kB0FLav
/7JoQVnGwgjXhVLrkFT4tY2TJ1HAsB3doIG00YFJA2IbMQpgHpfNqOAu/cxY1lLxql0pFjQsX6Tq
Xr/0yHXs2tHUFZlMHbwDDcfMRJm7cAs8Avsg5IiornqFERMjHRKFUmoVxRIp9PwJc6oMSHkuUcQZ
zzKVexzy1KN/9T6fvVhnA4G6RmvUBvkgimmDSBr7DZ38RkObiVtV3EzhIwd1F3oriNDyTkAqcp5h
VjC5GpHoZrPh0jlWrexf98xyMMKbRZ2+TLX4/AdFB4q7r/t79KwTE6egQXnO6osM1RPzwXDRExv1
7wpV+rJBsV0hUgFumbXw9gtPgXcsvxr30rlujpng+j3WDmbdt4mUoR63sptQcVBnpDQpxUTsJfle
JBGwdMSHOmWuFlwnqdv94bTdgNrmzHQ25uK74svoIeH98vfCtmy7GUXWWkIZEwpFxoagS536/DB3
Z/eR4cNu4lWiYuvICTZNiMZuYiS9Aj4MxdS+LQOEgRgzqCmwvODg6hPkFhQb5TPal9DD49iUBqCe
XdEoJ/TTYJJCsvfS5kFev0YGp2IN0ZPzTsJ+/EWMPo02LR7S2f8X/QirBfBqVfel/7OqD+qEzwHx
x6yJXJ1QKR9m//oI1jgrio1XqbpCzHquQgJnPK0B9EOidQ1r0A5nPmDgKZ6GhnJpGD9Ha1SyocKc
Gp/eFHV/UAiavVn0GESY3V2yivYikWaWrG/rvGCmu+LxTcsh5QZZjUVisFazDAf/XKFn5MYyZops
Xf71dCuI8GaFT51f54CysapFMEvMI2Kgq26nqFp3fNXX0Zj/oRra+Xq2X7/BCtburGKJvQN6ajWh
owuCDomYnsUKKtcCbU5yhs1FDwteqkJPyx29x4g/4lf20tl2O9m+w2kWdheKbcsFNq/VQKpNabOU
CUTS9S6zgTd0Grt6LG6XfKnD9uKdLdpqXaZhvAafeLrm7GttB02OFsdK7uaudS1Hx/u1yPzyu5L+
rR4Hkc3aOnWMDoPoVA5uTlpQyR5Dgdsx3ziDaaXxtb1BynEhOqHewamK4vjYDaVHujiaf3tA83jq
zJXaoN2gEwSgAo5zEyllqYDdGtgr5eucXzSDcml9gH0tX8qgohuh12miJJWoluhTd2S4GNmZtl8T
JjHl054d9X8RhH52yAEp0lAGD9jPR7lgOQvZ9UZ4m5CZ0YoOg+5JbdPWIo87Bnlu5KnW985GfCPJ
7vbj0EtBb+cCqrNoNbjLzQGO54YRW5FexnrfvzhF+JmDtHo1SVubj02V9p77Y8YPeLO2fwiBH6Ps
zwdkuo7Ik9RvlDudbNJmaFMxjHrTqet812bYy5WZzmY1v/u1CoCk8gGMJf0rbmTYfkm5ppV46AEY
BvokMb/99PRWu01f8/V0yMGcmM5wnEbso/lFjAhz4tHpWGTmqQ4xtKE/9KndaXkdfgz8EooTMQbN
POGNcI+Af1WCG0nNuuqyIBhtMP6RyQHF5gGhlajvZ+IrcUrUauovcwiL3JEOy+07NHupP8gdkH4f
vv1zQskjHVStWfJ+je0HYHl/W6PWgGdHJL1mMR500/sQ9m+YHqaQoPi+M3fAZbHq+kH9EKMq6rXb
kaMl05WNChV47BV9k++kJdSslz6Kf5VkceBECt/NAfumA80axm+Nn9KwhzDb4rjQwdcowDhvf3j7
3AG9hd/h+SGl/aky+UJxmFE6XHcgtMVZMnEpxRplVmv99QENO/ErEL4+R6EhFVQAj8gS01Vkf3Hg
3t0Wy5VWw5tFWd8Lm9EOnea3ICTGQomeOjcx0L0GkOO7FAlIKiWolEhO3+Isax+I+KfA7c3SbydV
lf/NpDshFQESpjSfJVTB10cCJgW1ipbfhZ1qDPIZnsc04dtRKgi2AIiWw5dHGMSoGzjdZA5G5riQ
D+Rz7aM8Jc+B7wZmtUUaWREI5/H4yS6oOSNS8PfqTZoZa0yHTYT0rsRCnR0eiX4iJNf2h7ytDznL
VEslZs0+X4pa+26rHXZVcBCVu412wHu/ZzXxPLXINyCgb/lk6fLSZhJaGntyvqlrxwBShao6OLn4
zckXXNCOQEGP2C/zhBM5hrgt+NhYQnBHLskSZjiGM8YFQrYXqpltu2TYJ73+uUEeLUymvLILCCRE
RUxfczKIZySKhZKeklDHMnWQbTziqXH7UpVf6lPxFNa8ViVcV3sE+icqOx44NW4EK4TZt8LxLBql
is8BsE3HwaMlkr/uswLIalb6K7I84bZ8JZy9/IDDYZ8jlHJiqAE9M/ObtD4zwOEJVyM8/TGUMYRK
Ipg3bjXrfhfJKXwxKwGJ6r3u+7zTE4QL0Gwcpaeo3uyBj2v1uvic1xr5YKIsi10iCHHnKDqQ3JPE
5gCG9hq4fAoVCHWVWSgpW1tORQp4I+k2BhxQibLpbf1La0cCAw2yDE30OnwPUmj2b6fU9HGLjflS
FWqj9GrVG+cOlaNn8WPcv2a9UujMo7o0tZpc7Fp2hrxpLeXP3ufrttNbGU0Mj5xKbu0+4u/ARbpd
gFOrewEDe7A9Ij72F4Eq0jEkfAZkJH4SMMr3rYKhWm4pv027l5x/QyooO1Kq9cigK+zH4Jt2SDtR
s+hLswoxlmoUOKF2Fm6+8cTc8AgKPyXjroywMZ7ffUb56HQORgxoiXRE70ClacIo/HcOTM7hOVlb
hYxDWtI2NL3UDzYPuRx/JX0wQk1me3ekVNfTy1oRraIGXntSLFMeER/mHNWwQrN9Hcd1U5c0IZgj
5e+9sa24Sxyos+9/9mUo+QtRx7bfpNyYr1HCcoXOboIbavJV6sAWPoDdWMzaD2oV89WOdBs905g5
AXetpxmE84VxNVOUEhTXLQcrXIggKFbHSt+3jY0dzXqt8ceXJMBeW+wDese1gPDEZhoRsxBry2HE
x0APGUvr+GYFAiGVTPDf2NARXPLjJY2xfo/XXUrvw0hE7x6M6tsfmHn2t6rAYfJX3cxhNKN+uJc3
gkrA8tU+fo7wOjnAyDIYEBw5AOfdnlZVh+D4daTiWm5a3jcVVqMTQbf7NXKsE9D0KwyYJnlyVp0D
cDn9md6YoFIa+RyraIsIiRGMA5+bT/SM+QMkFSz1BrT6sBm8XWmZObLJZaCbbg3KRUeaJrmvFeIr
Sl1MPZf3REoTtwJHQEmYoWj/oGcukceGzloOF5DMm8DmzyDxvCG1y5tcJUNcS5sUs/ZNsTXQ1J6J
wnSysXZcODE0lPRcs55OXNBu4OATLq+/DN2XI4AoR/KgKqkt+8Jbrz5SKYPrIY2KXMelYYmUrz5z
kmpQOVoblV7LOYdfTU1pKY394ujzDhpf7Uqw4hmlsRW2DImt+RO06c99vfa1uixOLUh1D++N8Mu8
u7cgoSMKyY/Rm/lHf6HWqMbu4OPfsjLOcqABHB6jTtfb6BEHZY+t+0RjK+QyYXf12c61ougHWCcT
OjDpL4x/4ExVoXsyzlY3DcyM9GKNlPYHUAAdAwj+HLyjLdy32KwjQ/Osuov1qtHXLbNkMQnHAv57
BBaq6LJqTR1pGDykYILJfKQf4wMiQoTWNC1cLUwnHV15qcZPJdIDl2YKtSKbARcinGi2bZIxrcz4
AwVOp9mNsKq4dKghmO4vq1uj/7vgHApz21r9Qnv9dBOn8WvgomPE//T4e+unj6aaKQDmX/G6Uhaa
1I05lF/GEZgBmweXJJr8yxj6i9ZNKfro10VRbb68tO2iFhctk4xjmdTng2gnDmS6eB7MAtTdVpge
mDO4iFK0F6MMI4Ef491H6EqDIbDk/L/UVR0NaoXKglUe7BPizHOW1Nz9piyvB0dlZZqgh7UFYb9b
AKDZGwDe3LZvHE708OaYTnGdIAX9IkeCa31Fr78jC00pPkwKYj0sUFSQTO7Qux0N4nRqBwb39+7p
rEHi/Y93F76h3sEY
`protect end_protected

