

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
US2mB3ZU2xYMwSgf2KG3QONmAU5qxOR5gFmXyP3MzegSXblZ76jq0dw3DGi2XivflSREvQG+tGNr
93kJJN9RHg==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
cVCcDe3dO8A3aQlcacvtDrMlOeMM3iFulWP1GnL0AstVpxpdCCRRxU3UHiCxbevv+1Dnaf6o7WxT
G4MiJBrZR0NZpyZrN6elCTa1aex/x1et3mJ/kXtaSnXZDYRGWgFlsFwFLktb6kdkyrjtbx1rPCM3
CfbtCvTObEIGzIf/FJI=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ybpmXaWiA2h4ouUhToF83n5FZ6mSwY7i2SbAGhh214jlEV4EAw60pDdsC9S1DXRUJs2H5ijqRHjq
O6r3TnjNUgOULu96coukm/eTQWKkKJe9Aqdi1COsXCRXpY/qPst8iFpcYgvP7x9BLqj2FuOVCOp1
vBc1X163t+3g+Wnu5wdB02cYtsPg85Aym4KDvpdGC2+lcbTElJIi+JurCHNEVSPxn/s/byKj9Aee
BWqSso/XFdRP+TM7huy2D0efcTINLjUE/2qeG1Z2VdFBpyOvUXxDlOhNEr+qAiw/pCiqNyrHCapM
TfSbH498t2P5uuhd9n2zpj2CUOFq13OvODvHsg==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
o4nr3qLm7Rem+yVuZpGX2Dwzye61TgXXpiZsrYTQhxAIOttLQ5qy48oMqssSkd1Afuq4E1AgeeLD
pr9heGHoD5AjWxk13hv9r2YUI3BND7NaVLyrx7mIkF/pxjMjFTBF3rI5FZuYgxY00aftrEFjG/AI
XeOeb4w/KZQIUde+tJY=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
dHlANyrutuNgAtytsZMPMatpxiEBkM3u/gDZ64fIbSRqU16FBJ0WguNKCot1/TeXAq8CSJHQCt8x
3wxDlxfMsEEJdw5OF5Pn172rV07Ce6wZ30zB83ou1uUKjnNgy6pYqTworLe5Tj4SYl9VY0bcZ0g/
rN0niMih/6g+8XwbbPNRS7in3icwjpeqxdXwsRyEX3dbCrKVz4LXcfmP+ybNfKunFSp+imrzoFLt
cLJF8o/HdEoH/59p1whEdIyNin1+Ra+5d2hGnILLEgUP28LNS8Xr0dqjxGFNrkIDmtSmsmF2E1fl
JbLYu0fIIENjFn9nAJCzGQU523347ABwMPcyhA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5328)
`protect data_block
ChZP08MhNwY+u5cG+iROPNeE+PsKOuyjWeWjRYUUKkxd7W3ZzhmRf0gNLYcj3HH4qUMfxp0jv6bV
Ffp6RsLSXCdrJKvVcYRe77dDz6dUbORRQ1dIFapFHv13Fr7nxfFENvfJJkL00LXCqSXmHX5f60zn
5coBEFTGnZfbbssIT9QIoKEcMi0OqMbcvAIqff5SdVsKDfzR8ieevXly2H1qaSLSecrgePGv368s
26xStwS8RN2SN1TNYUZmKvccBNLSz6UVgYvzcemNlvh97Ru25moVK6652wwZydqdyoZro/6a5tM2
BChNNVXsH2LEPKgchza4EG8sMu0JT4UshDlZN1GsWwxoFzKqB4u0iYX1yxVBnPf4potad9tde2Al
osCkwqDyn1whnFc60GJUZhsfQLrycqhfT1G+hLOyaX9A3EuKohk9xTNQJ8P64/0MArloD8dtFMGo
ezurFEadBvSYP/MYF86IwExCuAtMFc6FRhXaQVyAXrI1hYfyFYsinhYbfRjSHb1nvSapfV2Zpl++
EXek4YWGyljfOq0Fz69LIvScCSmwlug7fb6avRxQS/BmUf235EPv3uA5ovHA8dC1sxHbuzREjdFa
Q164BgYcTv+Ea4L8OS3LSbT91fkEoZTtKi0ljebL5TU1RNGB0gkYTvEiKfT9zL9PIU2guUOzz9m9
5+I62np05RrDKaAcHfi1Wrw2+7QYhP0kCj88fhxAX9eaS2rdJuA0joAyJiA/mnjocZcivzwkSRs8
2hgTUZc2Nnm34td/QeMyi4cwP+Cp9IYrQEnNUMIlqe1VNtqskeXF05FY3iUcG1GRRKsi2mo5vXn4
kBB+ouNSF2i+gqEWLWlXaNSWYJJx3M7edLY7wpVmhm9Ws8eX1JQurEksQcd7vui/w4GlNdfVQLRu
ILQ6z7b+6xOA0EkPzB1c84ItzhkkJq5N/dE3NRP7pbY91wnq5YksABzmDt8xqhIiBDqvuxdRbM0k
edKFrbeFjhxoRec0sKA2rBYlFZs3xsybsnmttqy5gHhyb2Eru3yeBF8Wf9OqtexPDlx7xaUih3tn
BgmiNVTQ3cuiOg5/lKEIwBHaRnrf6cggv+vNpIC2Myzyp9vQ+FeXo6G0cLns2iwAHJI7twEenJGS
DGmzn+/ntVl02LpgIuj9NQB97zIoC3S8Zw1MIzvO8dIfHPoo+yyKTPRfIG9F1Dw+j1689RHyxbG6
n7CoEpBEdYssgyR3HFBk/0JVNbHNvu+osb93+X3bUTduI4dPTOphcsOKUFwLKRFhMAos4e0rh8cA
jKg2AlmtKk28kBRyIgBFJ+5Czkr0Lj7gbG8dd9rlesxisRIKZWDPD+Eh6Zq993of836JyiUGL2MM
77WiY4ItCjcBXFuMyShaS65Zzl2GA1jJH/jnj3w1l6SROedAGVqvEjiKnms55rC6kKCeVeHPOtQA
rgcWrNgCvFwZt5CucE91SRuxJRkrJ1Fff2ulWeXUOWugvev3LcgkqIfyO0Bs8+VWQuLMZEQQ0Quc
CxdJCRSe2PyKFiydWW5x5S/fMMg6grk0cRCjlWkhlGdMKM4M/2ntFY9TKJEqjI0DOPKMLsC0r0+g
sZayo3jWEK1krexGefKFIEjOJcnEQNq9MVOUwHQdP/FPF+QksPlCDgqNnjC5CYNfVQqCtnwUmq60
aG08exCFKh1H37x7aHkolquwsLgmMRFsgb4O3Fjr5ZHEIJ84OmvQn2cSNTKYjIfgScYgG3B7xSXS
uRpOAADVKI3N7AmeuDBp/D0n1x23++jEJVSAlvgHEEscyb24RO/jFG2srzHn0kVFNO/NKE8r27Bv
O1zLd3Q+UTL6XeNkb/lKwwAnj5KmogxZl0I/TVMWurJ3NLtD9+VIRBqqLMalb1UafAQQAWVlX2Qg
XapakRuoEc1PpR3zHw2DIjD4Gi3XlJgdb8pfSc/q+Z+5p3Pf4By13uFamaG+SKq4E+KE3VKNzYND
i6Crq+eVEUtpFjO3usBQ4cq1QaokL1d/dZyrC+OWbHKL30EUqr2u64T9eCHE5JKXjb9pGjCSOqbe
rExAN/gqAik0DaKJ1qpsS7BIP6ceUYo3B4m+6PeIulyxmkcMbge3AMtGN3vtb6SCK7B6pFs6BsT/
Yn1cosOKJVfrjnfZ5qnSeFZehrdTMfKfqgi99F16FtJ5IN71qRth+Bn34amjXfuu+aXC6CcNYIea
tywvoBJ0Eqjaso5Cvhup+oKkY3O9JIejETa99pyKWjtb2jjMkEg9SIkU6VSqF/XfkwK898yMJ6bX
RO74mB0m1ci1EBfyIeNXscrVOPTx0DglT1Mq80mqPII1Jr5dzhemj+RsX1Om//ELNGkf3AEWAoyd
Onkdh034EBLJuVxujrcjJiIVa/y8VXPDN1UGtoQhAGMGz+HqoRwl/E5Cjh3FWXFEOsXNnIogSz32
Wqh3Ka7IslqSTKdIraW4myd2o3x3X2NFe3u6VLFf6IxMVP9roG2d4tcvM1xhBeDNI1Wkk2TNRKes
2grY6O/dCuKJfo4cIHiD44x6CPhfq5FJq6RxSGki3mSBjdEb6KcAea5qkWQTDwbJ801Qmz+uzxQN
J1/QMyyuFBzdycAgo+KzkNDrHHfD6Pa4xvkXJ4Ase/wgPiLdHsARPT4nj+jxoOb7Q8QCadFiKo8m
gPcvumDZDuaM5O29kNw0PqTgVeEL0Dn3wWHq3AqlhNu/SXZCl4dT4BwmNGqnxgPVilUm7m2a5JvC
gZkhpvKrcLXCJW3Lriq5jF008YpLaeXBV7bq1Wzf+x7znFr9CMB20b1THAafffMPkO1N+BMJ0cZg
AcuH8kz3LA1m1arQH19lRWkfSF1J+XXF9sq6n5JsgN/nTz3v0eQHmyDVBH/tomtzrqzXiSVN31fO
yHdMuHb0YZ/gfzXKmx27y+eHRKnGw7TYVZy6jI3adta9OEptxiBAOmWVyZDUWBe7IteqY63/7vnk
fFT3cHAVKQf2Z/1n4YD2Um7u8H3vKXpbfx1fpr1bE+3qhC8AeHRuQPddR00MaDJz0olUCM7dOzBk
XyAMexbi6u6OKB8Zwfg+SNG4yYS0LBuGERZwtHa7Lpp4w0IMK50+8Gtqo/7o9I4TKZl7DsLVRfS9
nKTHtfsyEM66tmwWs0QBVGJJmSTYF28j+NDxnrlDr0QaGzDDxQTyuEO5GAYqqcpE3DRT8nX8d9Rb
jwsypYO+PbzO0lZB9ZBuXo7pifAtQ8q9bdDQw5R0INPqH2/Y85Yk9SOpcSSj0ah+ln4mvcULkOLb
/7SvNSqE/Ok6pOcDjjXvIsPWljbwncqC+vR7O0ROIjW6FoNzlaqCUuP7nLlZS7nwjQhT1IlhnaJk
gl50rloDeRunM2Q5cdE1UFF0seFmfqFVZZfUnjvX48Ys2gLG4iRsp+GgA0ccM4PC1Dpe7Zv7peaX
RvyceXzRPe9NLTMAWGEF8SsLOyHQADPWLE7t5BVt5AUUV1xRD06gRMs/r9ekVhcLOpJrB2zammbG
l5OGi3OG7ttgekCFhMAAFrDVjmyVJjnQ/gF7WoSKFh+Vhq8Fox4monNcTucchvxgs3EWCvG3pqLR
w+8WOagQMwQ5TQSPHU8N0F30O3IjXv5KUcYjrEw2GQx2FtmiymoI0G0klq1NGI43u1e0Ol29/xVR
bx83bidF5aQ5892QkuWTwLZg2qZFJwLRvwpGVsF1YNhi6O21oR2hz0kBVlCKjZKhEjRlxlZCj4pF
+2K666NltnwIteAuXMEeGOJgAb2eoWUpr4CDxDltaPFs3ZufnhDrByHi0MSQVQBrJNcdyoTPiu3K
0dlx0y7IcDy2co4hJo1ylwYYafoznQH59ZYtpeU1qX7kvFFGwy7qRk6cuCVKya9CQewQQoFo2e+l
9S+QeqiCyilalhaGl96Sl0Wicz6cklKQjFLE5D5CVahIcESWqANZR7N93V0CEsST9E5xymlZld5D
6aHLj0AH4yyQQD02XgnagtvJ38LholZko/RnJc1aBM60ZYn4DZlJmuz+TpzgqESed1h6mf+WgZvE
piP3/PlV1fGPN/Ko4wxiJhKTy9TyFVX5CPdutKbUhm8YCb+G3Tpjw47cH3bedkXxbvNdd/y5i8Qb
uGriIJQvuYBpr0HJ42ZOf15/cPoy8eU5H5v8XoaopYPclkVafzJQ5HQatElYQzZOixqTbV5a13gd
jLgvGxXqyjFGUNHKgb3IV4HVfb+LOxoreVFkyaVU9YaeQeUFiCp6VmXDD3RGDGxY88H9lQPgu5fS
0vAcejtKF/pte7xyKR+QwKReqMm6YXFrYsoAResPmDJTwI4uB61tFJa75OIdf844TC9QPwxUs3UI
3lDfGe7KqyIVjYXEkOiKENHCecb0emS0Hpb8pCyJsTxSLef/BQkN9La9GkjOOVeyiVHsDt1L9Oe9
OrgeIknnndqMmuISMHqCGFRryFWD7uE8wIrCULYo8YNs3RCRmSziPhulzpydvWrrYoir6Idq/Kvp
MnM+hobmKo+pGLh8frJd73DWMaZlfI9JHJCHjmfzTFs1iZaAfp+IOmzBhQkOvlNP9dVYy150wA7+
ELy2NrZYSwSzI0y7YVlOfRxXrkHw24ClzDgZxJfQB/13AUxd3f8ivtJ/DE8ZuMw7m7X4V9T4O2qF
feAvuoQUlupRxlkZ8YOeRPXvbHNBt5E+qxfEFhTtDvOrOky6plUopfelLxHye87W7LBN5s96yA9c
+OalKWW4iGmdtWOWcpkDWdBKUqLXJa5/5DwBck4JYI82WNYImidhJ8NoKK4GiHu5XcHjmPKJddbG
AZ7dWKAxYRwg99BbjuKz7j5iCbD/WBvLGPDfNAXQfAt13pj9T5sHxPGMqKfWCcWDBYT4SQUWFLLV
S5jGQSsMLClLDC8l2pe/c0HLuFkeyhU9HTcnwq7NI7IY+TS9za/38tudKZAJxyx9RgK+V8IqhE3L
BN0wZcy3+0mjDpPLYy6+upF+aWGwvwyIjDCjBPOYRP0CUDQ1JPCx8Ktu4/Syyr/9pnO1RuGGpU3j
bX4GKCckY44t2Eu0pu0lHkaUYixDbXzwGbc5BW/ikfPxCwwVSuNX9RKcCh/uPezycuIt+WICfgWl
ty7iT93A/tjxu+etVc7cIBnakCgcb8VHa9Liv22pKBPsgs5Q/WPaTe60WAVulqJExfjo/a7s+Fx4
Ygige116WFeunANxUafAlNyoYS8vmqVA4G8if9CpdMwUKKJiQBHLSf6C1zu+63iwlK+lniUDxopy
AfR75zjaIeFACj9l5w1bb9Yjx9jDKNRGCvo/Mo1FOc+EWz0ft36EwYMD34P+1Lt/6gJJ0VW01Ge/
sXyLExN7eKxeaSVINjFQujDyV/8LvUkq4/O0+Jth5cbt32g/30fguZbWHTberQOkYK3nPtWpHuG/
eljMg3edDkBkyQMD65hq2yPYVracewahddAiuOZvSLbjHiUw0oJjo2BpW4X+pkpz3kO2u03ji8r8
NstSUEt4wQxdawcY1Iwqpr/ZiGOzSaAuTJvEWFJatOv6ZzVMCLW5fjd4XKRuGgDc93/4e+LRypG2
y3q+pCKnqMz6lqx11cRWyejl41pEqbFqKXuvl2lphZFOFhY9eHOBHbnDe9V+rdmOMlSv0qJyIxJV
FwCrlXSWH6+BAvQ2qinrQDCyHyHXMgciU79K8f79ZSpiwVw0qrXzCtMWqbP2CYu/r1Et0a3GMW/G
ShWSNPac1Jlfco0TPJfC08ZbI8EqT6+O+YdsAirfttCm9wj7dAJHgoDP7/kIrAdV16jmfxz+IHJU
vSv2YiOuBpjsjrnhr+PbSzUEJ025Kuugjr5ovWhvnJa4gEQETHvZv0M5FQt4/lw4RMYji3yKjfkl
7wo0VPR4VGVyYnNo3mQwBhWOVAeB0JUOt+NAjnh8y7/fngHAI0O/1ahlq+yFpatpUT+iUfRVtvOX
BLfl83s7J/uXsVo4fQAETOa0G9eFa/UrBb4h+wEdYWcX2SyolLmIc0RZCyyo4ctxIkUhS/p+hgCO
TgydTkUzNQpEcdQ1UQWiOF2nYtQn4Kgke47uVdrnJEVMLj4fidv/SX1R0Qp662d3ZFgDF9X6QqAV
qpYLf0F8rDg412j62fsqQPQlk9xacG+RDGGJ6w9Fwr4tdOOLH0R7EsexbjzVT2y/s8tHC+NaIL+n
u7y3cc3fmSF6jrTkI9iRcaPJdLqy01BPcF+c1LDF23lPyMg48cf2CpfiHaW5Gb8NRaUdMmt9ljxi
Gf+ri30DMIp7cntpWAGHP7voXgu7vLNxigJUdV/0f8FsFjZoRXa7Wz3/LtVUOZFboouEr5KenIwv
AfPE/Chjyr20ue00HXT/k91T1fR6x+ODEObJ78vi9jf5/hY7kDMeZcVLmLnHCY6R9e76eigvfyjM
BlSawUnwiaz94nMVEWMqScC3SzJCnPm/4mEb5KQdlcDlHNSrV1lena2JQ2hiS0ek6BzfO7Xt7sJc
H16DNABP0axZMIOI2GlFUvFOpHGTCRDl4uKC29gFL733G3CulsYRWmDa6y2+acbJsPFAD7SbiO8W
ajBMZp3cUMHSsfpgwzIs0MUIAiSFpeMg/dKg95SFT0dKBzAn3UU3jltzFx2H0DBiTbCCPzb00E3m
glZdVt86mnXmkmCkP+LtheWEcvxhRXTy2harvdyAM3ULBXdVAeCBTlA3beRZETJIZwM5tlZspMao
KFP/aOHcqiHp1WiKd4z00nnBTGmpxnVZZoQRHI4WVi1ivENJDZ6UnhKxCyD8IwItd3QipCmD1DgC
LTsVGwuGvw8YAb1dg3H00CCtJxMhhMt0hXzWRGgpXteWyt/7h1DcdLuBlv+fPLVhmt5Ik3L1neNw
Czj+dMcF1ZmFyCcTX5+nZrxve68sQh2krWvY0AnGMEgKmMGSqVPmhgc/zlCvTT0DnYF/4iPod/G8
HQBm0sqHKVsAdVOUdtXlHE6JVg/+PUcLdoXNdN8Nkt2xjN5QLJGAnoE4Blnv+p+LZ1W3308fm1Ed
mO+MNkl5zyBkJeNQul7ixq0avS95lV/2rPghNYi8M9/j2aMQL9oncWfAEdZ03oapNa4Nj9/ufCHM
jJnTYfn034NIzdkVdgY+s14TN7ks8b1Ujlp2
`protect end_protected

