

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
VqgplFNkI2rH3rP35CdiLJAesBBzx3ahYCWVov2QY8pnSpbbPHZzKXALTXuf8Lg9RV/60SesvL5+
Tx0kf3Xi2A==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
YpVJ/AkbT/7j7nP1FpW0u/1drBu1Ym0xSQcZVVNR2BH9CeGHgikyUixQxXpCsKnhOEb3pzk2wV6b
2udOCqgzaZfDIjjaxTt9/C6XIY+oMyWDycOTnGwR4Bf/A6rFEzTLA91kxNt5/tS1PVy+wjb7FCsa
mgkYj9eNUdtmSsLezko=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
pSdvSF3+OBx+pmFIuKYX+lTRtc2CK1xqA/WmTxOA/9c1xuF8tv0giSEc/96tBGsFFqc25YHyYiXZ
gYsCabVJMk2jc2XaKW+XFrRUGrQYLd+QPrzsIggnGqpN1i2vEJ2/57QIQEt4pR4jX78IzCIP9B1I
Mief83M338G9aIgdzONBxsD1Z3XK2M1fqZBI+UT4b8E2guDKnWsCC9f6WqxH/+ijAu2o7kXfkz/w
wH4eaCjn38eBIq4U5maYpwbVxvzCRoB69hlCwEEVDievRmXHouMD407mzOTwKaIkf/tAbFyB6i0D
s5Boa+TiBtHShhLBGBRqGoq+2UpGEaVgj8o3hg==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
HVe+dxCY+VHrZ/rUbzyWsz5ix04KcDyyUrFaCcS4yZ4GTBKi9GYUFVfTsXMpSX8pxXieZIsbIrAR
8ATsmu7QwmViHDzOMuS6sHzr6e8dC4A3UKQC6xKKwbJdSWPz/il1AOb6t1CcrpGMLBXMZTBj00R6
KptQtwRx2C4sHo/bHEs=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
gr9tWfnRHlUz7X9jwun0huNacy2IvVfab84T3X/BBntsyGpCEQL6hR0/eLuvmgsVt+peH9UtRKIo
Mx38RlMVlftuoIDUnixeoGaAc4c+4+tb16q3/5V7og6YvplXdBH8LQEEDNM3+H5ouvTLLeMul2Yk
sNNMGtkGcvzxpzj7QTVn+eSHg5B5sba+LhJuLxq02/5r329tzFZy8dtsa4HltD5DQbMsj44UHU8g
J84rl4f5z2tzAq3mdpwIqfhK2vn+BHZu8UlcbrIJKEkQpY9EPDhgx0vX44IIfHNFCmG2MgNy3yn4
3WNmBdtLjzwOjBTyBBtqdvJWbuTYLVDhGJrWQQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4656)
`protect data_block
4fPgYLBi7ZHotS6FQqyxLw4hbf6kMyc5irbuzsLPfYkdT9dyrX36zJVYrYNQJKth+AfzV4bNTjX+
rADIdVfj2PxI3AfhiCeqQdP7BD/zsD1oAzzyFsipBJnGcCTaV8EFO46Yn+7nxNNAfq6o9+HZH+Cm
xFfOBuq6M4jPlPeFcE3fZ/YtO4+hDSVIqF1Q1lhCp337+W2ORiq3KyejdKIzCZDiwjZcDDkt+gCc
AylZdKDugdlLemUrcngUlCrpR972GAj7W1dZuL+/Yhz0bX2sz1WAt4gzwLeyoSx0uZx+oLMZxABi
b7UiLYoTGGWT9CwR09y0FLMLc5pT5WVmCW7S7QLWfdygQsb9jDtSMAonlFpsR0rEhHF8E2Hruu1X
SEp2ve3ySFECBbqnNBHx+ecC9gCJ4AEfZ2ulWwCSpz+ooiR/0KOZiq7VGcp9YHov3bwSSq4HxE/G
AT7wKoh9j8VRsS9QPYPaRVre+Z8gZiRK3sUZQ8ZpFlR3mni4ZjBnyonnznJp7e1Bxhy80l2ICI88
T6359emnEci3RkSY4rZYFBpDe9Q5pygLQyG3dESR1uW9ByCsIqjuDhD/q7hd88I8ziVBQrmF597n
iLSK9j0TVDLv9q656Wkgwh9b6Drx254fbL6ZrCM2kD5O9WIudO6vK8dcUjQqaruhFtoMdugg6ozb
nPSr15aFVRcFfAmZ56oSH4KS86XQrH6Arm2yAI/dY2LuI/HgjFOYBc5kkBLGcPSRRBrVEwOuj4na
5aVD4RJo2VNbDFvhm6ky31R2W6XZ4GXVS8eaAe+xJmrNK7b+MOLEXMultLan/RdgMywG9Zzg8lcu
ovEKpaSad2334ZwE77m1/4xwPF8xD0fAFwEFj/j5USSGZjEJVpoDcyVxebReEL/bxdA0njiNM1YS
Q1JIYqo3f7GN9Zi3Vu/ng0g8jMMqTo1c184jFYqR9jHde4uPtxg0Z1FL4w2NVpZS+B7Pd4fJP5Tl
ZXdKxJDY3tM89T//mWSispo1HcLeMpyI7PFi4VzeJJJQ+vJ9vHJzY57WlfaJxpvoqZUl6+5RKiB0
l6nm3SNFpLp2z17q/iKGzELixRWbZh4t8MEfAA+epWIeQyaVPhiQAboFhN14r9qEcTDzq8oxcAoA
HLEjIvf/wi2iKvCBU/eIN0mQEyhC2/dP6vF8eaZQbnXZzptCfquCRUWVKo5XKVLUuFgpT9AxWkqS
anWfky/7i31fx+o/SkxU7qBFb2dRvKOG/SkJzuIzZN9VWk5Rbl8a7uE6VF6CalG0gtuyIAnXDJVR
8Lr+FZS1vuw0xdD/UoLdU2yOaBCvHzvux8FMJHA8TsbHfXwudlK3gWpbLvugj/Nq7Hc8fNSAqe1E
vX7L0bEowOs6BDleyFd0lthUP/UEemo114/MAWNRdZFpz08xTcIh3Hd5a54x2GeIOjaRe8zKQaZe
NgncVm0COgxYQVt02TPA+GL4H/HA0gZqMjbxxrPXicqOEHd9sPcp97JgrO4o/T8hJZsv8KMCSTN/
dKwWnatOeBXOf3sxKzmoWqvE7sOlPU4v8BjLePn6NFKho7k5FlZl+T+whxeS+7a+z8Ndxap/8Gwe
04RBcJy7XrRt5LZ0xdEktYUiSn4LllALOYEwZBWPmqNrhMhk/3TWBdBSOQnUnPz+kUZ72d6xM/kE
KzLDLDtyzAVYCqanmnjMpbb7/4JVkT8JGZNZ6wDtyM/3nraG+AwwRtZ5I68vrUXn1nO8bBy90Wgl
K8w5pVKzUEiZnwDnPDubtfwIexB0t/KZnmVDfYZNpx4DErvbvdKFKoABrwmd80e7D5ddgFMk724f
1ZS8bibVZA7OJSdVAKCIhbrC0VFhr65SaMxaCjJ4JVROSe/l0FERXEG4mNF6Tqt33k/7RO5gLPGR
bY/qQBTnl/dxFTSG0CLPQncdQekjGFZUYxe74AlU8RqBFmuwD8t3xKKwPJj/sq9Bn7Dj77T8wZDY
1q4ic4PVGG7W1df8r+GaKVpHcbtbG31TkRbWOMcfhbct+5wte9kwfd8D0FEVo7Q1jTqs13B4UKWC
J0jAnuTMXTxmfq5rR84y9SN3STbZ+bZln5CBSVlXXZcPwHD51Ncv+Ff1j0LUJ1xQYaOb8vU5lf1N
/IxaaR3SeaZ2bpr08TbOKLPfAwfWaC0Hr6pKXfgTUphtGLPt6CiOJZUH8geC05VMj+DEH2NlT8vV
gkw3m2lyVGrbvolgUILySzgWeGhKVSnW+r3eH6Nqe6NJZHRQDsn3pEqbvGj+E8OzQD3xLTLqM4xK
6AihS6kE6iOpm359KAHByqcuL01wJFY4UbqLFpgFK0il5XcKUUHajFWhmq1WVS7NKXXQ2r+G3Dk1
URfpZNvgIjIO6FtS75g5dUVDvakk+JsgwF0RMQ1VpryRVdWe4cmdNRu6dt9U6x+R1R7dpsbVoonW
c2CUOqYcSfYyUjjx2RKovB7N0mzGGVfOZdxjiL7U6ER612iRh9agazg19GsjZe+5lznV87YjskA/
spNUyhKGH/ENSS6Dp4ooXLgM5PLgpke3QRecXE5qbLcBPeogqqaIfSthLWLAHTDg+EHLPnx52r4O
CnlG8w338Lxc+ZfAA1tHJI6NHLW6RDLviEJK8iCLxTsQxsxQ2kWifeJhZ7K3KoSCOfMB3MBCIOxI
456A9bcKzLmHF6nDUBs1QMr1tIg6P/5ERnM6tjRCVsUuFhfg/qApdZnKDYmZk+YDIAMAvaHfgkzh
Glex2QEbwJ3uInTd1I54XmkdpvYpGt/FTa1s2/TAZDutkmbANy59801mPGBjmnQE216GNEjCO0Hj
fnPbSesMCO6aL8tj0Ya6vzQsp+WsiKMBcQOqL4Ox50ozp4Z7GBSo751t7IOwre1wquJoMttQ9pOg
DDHwK3vDWSkxtBA6b3sB2luVmYRYSmPm054I84YXM4VjzbCdpjrEkZ6NEoWpCpBo8HxyNd+hYb2h
aws4EF3CknnfxCtKcLfcrQz4QhCiJBRRwluzunaa20Xnr1qz4PCnkP7v5aVnQMxe1UG6MzYK0i7x
x5sZrtTbYSHjg0Xri8oSIdNolCu1/EILyK9nSHoGE0G+G/3g365O5yihoedhN6L1iuCTX+TSD81g
XogvEJr7yLfV4zQcCPxzWBhQ6+N/r0V3n6gpE1x1fDrWNSaF3MtQh7BcspN/207H/ZnCMOTUtit/
BB2330YRi3slm8ZEHDh1xnJLNOgB9Pl1QrJT3BQWv1YdLtQSDLPWWHFC3QDA/P5YX/DPiuZ7YnFh
X2CjLSJa2w+Da1LLRyixYpWXJGrKfPdFywdlkvZ8hmX77eASKpJkT4YzVrme7ozYxpYpIH5tyECY
GQxauYpdDBqaUEMr+EsNzr3/Dg94ejeNtljTayZvT6dnts4chwMvhrahfPixAZPA5bFrNNk34loa
XYEQ/lvTgiarxW4QIrUMveV5pGVL3pVvLtxqfAmF644jALLhta+No/RXsU5yCQFrk+t0KcZod19E
jg78cT0UsxP3hoASUPBfxt9hsgLg2xwQRg+qvkunw4a0SOSm49f8lcWrpfoctV6EolYZnGVfdqC1
wO0pXZcNFtcYMhM0r9LvOci1S7pjkiTL3vOIhRCpahll4iO6Skc64eQjq5NUXjyGhNouZH9aYGan
eFF4DaYGAfZCxTHiTcC3Q61rtAo8yZiE/TKWTQCSNY4xXjiD6NBqhbamNnzGTo3/Fj5Lm5VFmcgx
bFJMgMP2hF+KrhO2pXZMcgSyR+jUIqtozzkIGFwx7fpts+uGqTrCozX+GQodkyeYQGqP54m6YCqj
Fm2kBHEgqrKkiodU6XF51Qo2ihavVASRMawSMFJO+4rBWXqx7Bgp5GPdh29zSrfs/+VtsDzPF1LO
neWpg4mRMYxUFkgX0GRj7lXz9CvZmBbxIF+HYTHO/BgifjdZuN9XL7AI7nF38o5x+YqLfo2utlGE
EQLIzDqp12XKoakPeOVQuFkW7lrDL4fhXX+zd/smxHV4Gdb8xiv/06gHKdfFwctd3pWVdshb96M1
grcMZAicwxF6B0pqDojEco/oxNiVCiaTXuVeMppMsPYCfEGsVyi7YlqaKGZyjfhSdEZFehBXUYDe
FSxd4xTfJiVUz337BGkguA2yFUo3ZnGBSOQicx2dKAKznem5khPa14rOS8h4jKliKowpwanQodbV
7ontvv5zds2NacsXKIt8NoixFQap2kKgu9k15DsIGBZZRkPk8rZRq+VG5TfvlYv0QJMTwZ6prSUA
OyixxjYVwWDf4g9J7XbQTWpANwuTmjizImSBi2MJCDdRcPbJ85gFdzJv1HTM7ancPVkNX0VwVtAn
u8uunSWkivVSG0FfiCxM50EhXD592Czr8xuCAOPE2OcYZ4k18gZz0stxoNT1D+csgwNIxMd5yE7I
9G7jsM32iMyoHl5veK0Xb42GSPkmu0icnh9u5bvaXQimr7wIn/8mvwKpvG2HsKg4Gl+1aCzHOzr3
2OHeTGPf50bZzeLdObRxpAs08/Nzkd3JrE4KQHDWfvwDOrjqoIGvk3PyPDQp7s1dxXOYgJiFeGZ4
94NLTiadKCSxmWNM5IBcqOnCVIHOPOTZ3tX5YvOGyGa6qNuvY68EJeN3sU418B2xc5HTfG6N2Q12
COHqH7kvrrbTf1CYs6AqsJT+uoe57bteL9dvzqcyLdmgMwEFRrPGTTSHtzjFis48KxTBo99J5AQI
flEf96WWBQu7SyBHGntlAb/zmYRj0xqXAZugOeUeOk2XI2FNyMs7/4na3Egb8sJ0ZTUpqwNg/ymQ
RuifV1nCrgqAWWKO4dZt2RS9vEx+JxdJHpsKie2xv5bY9fwAkB2aJgW/NosUWNpwRHuSB0JNBuGA
I/vSbeGihVN6jY6lU8voZa2OMfwgnW19Ozw2Q2bYlqO0jM37Iv3X5ANCefIwvzGZIClmt5GyhhtJ
XQ7/SMIDC0kPesO4qdxRaJbONfI7NuHe49S7ZIMxoDuoMQEM9V51S7zB9qcubtsn9iYLmQAJB8db
jj2dDaGgZMWR+It80DzkNIsqKdRIDA7OGjPMA+pLh+Njhi9mUtpiJGsOtmoKPuZkvzJC8zeWtR8p
82WzjjSxWhY+6wt4FmPO65G9SrlkeyPGGQxh/403QgRjcESaoVzQx+7XQNK5gEo9r23DfcPOphDA
8g63wPYsxVF87p58g+d93e4jT37FPm0VkQkNOfxTYs/iURvwwUC5czsnRwv29X10xKmLyLUwFcOb
TjuJWpbdN/gyfK1L3unFAZ2XDWFQc58LzBmyFHZ5GTA+ckQ8FArJAcCDK/XAEbFXpwsgwPMT3ylx
e2648qnC/FB2PnhbJeRwrKHCy7UKNNUZBswye8NOw8YAJQLmUAQl61QlkuLX5P6tFJ82Up+HJkSq
ggKAq9dAuMNwjdODqNz/gqrUPdTujfE1mQCrFQNBxRPt32BLit/mTmWPS+Wyoz0YRf6mlpWtboXY
iP8OHrL/pKRnZHnFz17iOPhp9v2Zqa2yAdazU+5FWhxnjhfWJfgXwz+Qo/5bmH1RumdRNryfhipA
V5afG3ItAQY6A+BuFXfJdBPZyMqHhkkS98hhkbPQW8TIppMbcYP/tsG4K6kS1Ms37ytU7uUDjAw9
zjUlqvigyH+eSmaQ3jsB1jApzkPnS2ODWOb3mCtm/DyZgJZbvsBv2Du44Yj3eVjHPKHFLzLIzA6F
ZqRriR08tQM/ZpujoIl6+0uTljKBlBEu6hsFZ8JKKdV9TavP3MfiP5mW+ViGF4bYsh5S1wAmj5hy
N+xxKrW950rX2UFSaGqe0v/7gGUQJDlTDlW1pNBlZj7InmA8iHt50lqwV7G3vl1GekoPPmlF3Ntz
BCqFyX7juq3L6tryWu0k1R6SpmMKQOzSJpeq4+BWS+lGdbpf+vLQVONilR6+vkuSzNzHIKyLo5bl
EfnsH7au+F+/uKBspRMuNfRviALnXdOSdek9OETGWb5IZIgyCQ52cNMXk3nignaEajXH2YZrdyn3
nqxIEBk3WGHrWvfx0VCVDHicuJemMCWUnXQFLe4Y3a2b6t8w+WtfQLihKBTf2JCNGOBI3BOmAqtS
4Wndi6ZIZnR+QaliUMfBKqjOMs2D3aAhsTNmcvxwCm5miDn9HKmuzkD1akZCYpJD8lHhvLBnXsLQ
7MYIC01dAX6KUuUxIIMoUQK0O9YoZzCNAcuYbNHTuiW9uDCjp874
`protect end_protected

