

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
pabZO1I/O5UlEfYaQEPwd4l9eUai0bqYoMxFZDUmBPXyS95K3GW98Ld97MzJKAXXnSlf1PewGW2v
0RIeWd32HQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
MnYS98CLv6GUlLtXXj0MDq/aXJWBamrEeFXZFkhzX7OjMU68I3JzEc2/1UN3CHInfTII6cQBis+f
MSPPkhHYfjWA/UnlZNCfIbUjCA7v4zzzEDOXLdUwHhey61M2PDbtjo4F0M+PSYsHQUE61FCJYZr6
+aBOwyo0CpKkCUVEbxg=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
qncW/Cwz6DQ02ZtEcvyp5WdAA4sItotGPpP0REUtLyqefQhCtJmFILcg4T0iyRUg7VuYEwIANO5+
QvHNNc39qIJv9lOesalgHBZQgvNRJnIdYWaRfS0GyacwI/2JQRwAkuAQstvDCp4RTc3l8lwP6/ls
9Kgq/wnF0FIDD2zIsqBFYPVau5gOg+E2Yv8daLhsLbgUNkGI+w4/OZjRbQGSUjwZLuzAjcC7dEzW
IiD8iCe2E3P5aTpTA2tXeuvseQy8KOwVCxJQuur+f/bmnE2QrPi5PPQMRcOyc4ok7k5U/64SCKlJ
oITfL/xIL/xwZa26tMPcLgkkx7p0G3RLvL/tVw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Dnf6vaqe/V3pNaiPDsCpL4mEkUhuRTF8jsptuAsYR5QlsF0hNdnCfK2+aKM5H69faCvd5mpbM0GP
Pqz+qhNmOYPHdckgaTUGR5o/7QyV8YKLvzwfyDMqTu2isTv6FP6Q6welH2CNBnmC1/h5T7i+fy/Q
rlaoXYJxfrB3B6n9clU=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
IMf8iBP4Q72XIQn7cHjsTbT2wNsnwrpqWy35OTpGthg9IgmIl2PQf4/c9imtaZPdkPVpIBywT+vW
p0seCgJeCim8uHSlCA4Yuvzi7NiJqnEZtjEX9xSzaDj4EflUudOJTsvuYMqv/3kxvUgkIK0AS+U7
CWRV3RwJIjyzXaV3SkeD5i2xf0d/bezTocOrvt7wO8hz1n7ziicW5bgdFMZpO18+84bLDi0MzKYQ
Ad5OLz8QJgoCqRTe+B2lLXuByvKd2+XBYArz50J0pDfy4RubYe7FYpZdW50ze6dgBWVP0HOw0tLX
Pt7eQrmsKxnIhjnIQBRBht+Bb5QLkHSbaJnGbg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 8352)
`protect data_block
m4niD/XRWzq2PN+dQQl1LhLz6sqFJ67buuGjhD3s3Plk6UifuhpqEgcJT0tIGtdwgNU2px7au7g7
tG6+EoPMVDWqC/iaA4YP3trkqSUxeSaJ33jTadBOvELjszCp0qaHY2iT665814btkwO/lIubPLM7
ZsKeT7ltJnMSSYU0ktfbr5FvQoIlCQ+rvpz4LCb+jqzRaCJm7frEsCqjw+ustRf4d9MIi7/KT8GH
22iFcgi/iH/BhyqK7m0Y+OZeYRGDnQmdac9TLV7h3OO9ZKXFYNjXi4PpQIZatKPVePCwRdSnxIF7
A0vl8Rzk23RP7tJ//UJ3kJVxyevQbQpPEbHfcBaOvsY70yPTDGNJedhI++tHaQGBd9WH+bWPOkFI
aYGSfrelYRMqN9GH+TuMA4J3FudrlrDX92pd9kcwsd1iG6ti+5sdUcTuU1w8rPTbxxKgIQ9lyRMW
EZRuS227XKA177Ja44ugxFy2oCTS6hNXDd5vZC/rPfzfILfPCq6XrLUxOaG6uOSvbA43v3oUtfKM
QDNmhxzaJSxR5btMRzbfuelGsmlZ95DJyvt45dgp4GdvYx5ZMiQWqAX2LRA9+VoIzGhiWqjy+tlF
sE/Gj4dC5BLWM1CltlGTRicjiYIXUykv0UzM0CDfegvN9B/L7S1+NZ2eGEyw34uaVOdcd6yfgMHs
ir9nZxswmmjUhU0Kd3WXPdsStyOUrJvBuBG4GNzATy/6GnhRgDy9QPVjUkmkuCAyYniBdn9GQ0wE
4mnteLcppG4+zmUqcgw5yKVlTYTW5SU6JWRrpfHCx/5g/Cf0OFJ7KxeLgkcQFADbCz9LEeTl5gXp
c9n9vm3h40tX2+0egfra0DrLRRMxppv5rfnalGD4g9bPK15fpaaqslIGKjGZVU5m7l9gqvkNt70f
zsHi/oICNqiUL5rebAZc/mWjFnyOiK34wmK+/1pubVzk23CNRa4xJQaPJLidhkJFCUVHD3ZRH0JO
scVRqLqfRZj2kyuHjyjDA8josmavqaWv/05QSFZEVUBrQWnI0noart/Y4mWFbH9qa2Iml4h4DWrL
vbrZGzkTvwBUjrzVl5xKvSbq06pmD3Tq70EehIJIFwocrXf3oT0gtEgBuG7eTdv6pjyMxH3a/AC8
Em0EiHfolMs1+tCZq+l7ATffiDS2HgtVH5eWtiV2PKLX9MGaZnj0LkWHKYXHq7DDbHIBfDszmgFL
wwIWX4REJHibY/yr84a931njs6spxSwh3/VTWyyMkqNEuB8gWPt6guWW3BMwGOoWPLgbDDdKBMD1
Ko6yhxC4II+ptLRYqGrYFDU9LDogJgYZ0iQKTIdUpEhE9bMqxSg7khKOFkkueoWPQmF/PVkInIm1
yx9VUHg0nvE3nFkgaqnZDb0E5NkL/l/WRbGluEP2AjJkBoUT+6voRW0aI5nqqUGio6tZCGb86jER
6GIvUGaSeZWroQ3RWEuxy8AnXrZ3r+3Pihw4tC6z9z9UK3euL8WI7nLZj6AncLCmcVpBYAvpch3k
joLgpGFxcjJ63xBKjM/b65xQ97v8fTNVL/7QnfkpA9s+4m8pngce6wKqwJWqSi+DiRaOhAEJHju9
YEY3QOGW9JflsjBB05zOOIfH2EN3QD6GUAq1UH3tQvxDtYwnmsASYked+cbUUqOdnB4XW+QVNyXL
mmceXCYpLQVHE5X3F2tCr6eXCHlOg9VMHZxzns+ni/c8X5j7H8pwM2Ctj5riW16eUcCKuxV3gmJi
6RYS/+Qk37bkqOuyQxZOJP7+e95PAOLsi5hI4Avs7YQQunlWh3BvpRj4wZGScxXOATJG1LUjom8k
7Th3T0tMcHDmd7xdJXfF1aCFHh6JQSI4xe6AbqeR3s+ojGtGC1vFzWseEYuyCjj3Q3PSPiKNo78y
OP5yylrBVSnqwtFUNxfm+nAUaJcm4+c/ct8tHW2uc/DQP/4u2vd7Xy2tvk3Nm9bawUL98WB6w9wm
fBkyEGZiECVkwPzmC8uKij4dvE1S1nNqCnEAjzfFJNwYqbniqCj9eA3E9j8Q5YQPSoYVZqkuRwhk
gWcupxfuTmzBWn3SqOD6I5a/4GkrRYjTN9uO9Y1UVfaFgwnKVucDZBvEsBHnB5D0WXa0ZYfp0ShK
yAmOk5L7GT/a1caSf2jhMdNfrUE3H0HlzN1Hvmy/+Pcw1Rcqq/TucxxfhTSRAgKDF/ECK2Gh7OdR
GBtKQKHrPtPGKofGb7aFkMPjZEacOBDvocdg4My2vLfRAQet7tCoiImVCyPPrQTU3EeXdY1Pd8Vh
qBqM1T4OsIAxj7QDVwdvH2j6ZbxQOx4l48LWiNY47sqw6fMiX5gZ8zr28gGsVYIkHH6iu9/NJHXp
bXrgxpxBESktVjCLXdElLXFh3lmCX8BmfIqW8R5Vy2/feH2gMOkVQMAIhv7BKSsDsIvlhb3L718t
oSRlHxNHPuHNlxwH32CUGMjpA/6bNU109Z35cXy1pg3J1ix6zMRTE6QDRkhxnuxFKLR1fr1b0e5E
3bptuwLxH53KwtUwxa69WvfR8c6cLLV5GyPUKJwubftPnuz13JGvOcNl9vnttzJJn7IEVPRNSvpb
Zi8ML+guC0GxS+cnyEPyW5J9ZLjceuZLsXiswza1pDKO9zmjI257Q7fkLBaX2QS/99C3DFcnZzeP
VvsdhryIsYo3Sf+4vx7TU5pyZsdAX5pvkKkd/Soliyjm6HhNgFtdyRAeWVR651OHQxEzO9nADGUC
L1QBaBiiEoonzQ16EDVeYZOJCIaY2lCkM+I2tgb/edCR1LzDp56+ZUuw6tbjqZTvAvNoaVqWVPXN
xZlzJP/Bqz86DpIoTVyIx45qvjRZU73o4G7h7MQsDL+KF16E9ZP5pnprJLDpmltSBPDzawhtvixA
9GhLYbntS+sxDP41UtBVxrEFQbgX0aquXrCxN0sovPE+uRSLtrQZAhCwI9JqqnrWn0vFtf7MkejA
cDnnPqMuNFB9tUocaOOiJu0lAEkV5QE4485zHY5MNN68Bh3XpI8JI+MK7OiSLBi/2IrkUluqZu3j
2uLpcUhdwUnKWZj1UYfoRkZmm8oB1FgtUegAOEJcNDsvWJDoFGJ06HSPO2Fg11VuuMnRlKiDeGot
NAOpm6bV+Q1z3+ThgFMeqD1VF/xXOHlmD2QKQO3DsR+XW0/DyhTaR+3w3GyonlBf/whwvTc/rHTR
9lGEzo6O5bvvgn463/LA91a2mhK7hyveMZT6xnSYxJoXplw4wBNj7srUsWF31/ZtiTHEMzpV7R1p
bswGnYnQt6pDoqfXnqOwePMxmVfSx6A2XZCanefb1pvTFQuf0hDKMC1G8NNy+2WAy5nzgCbqPUMX
yVXWHZkb+0r+Ybk68djNkxUvYnU4yPt8IXTPJxQnjR/pjT7to1GJqfDf6IqXHuqMZAFMJaHlt7BZ
KsGUOVNVS/CoHxHvskIzI3Md7Y3bVsKOBqD6/ylp7iKTzkQ5l/A8nJa0o7JXVUhgxvJDLhKElIlE
KS+9xCV0wzzUWqW5+/MziQE6VZ6ryBVWEOoMwaHUfqh2x1yNgIQtG9WysC3AdzU/jD9Xb9hP5Hif
w6Zd09b5oO68rQ4kCykPGm3IypNv2+Ozhm+CpJegSHCOOAs973tboBPYOdlUQJUX6P3XoCCgheml
hiBxC171RfVbQeBVpYeNZ3NGrwLimOzm1J0BH4lik0KvlqdJLguIpPi6HOea4cEzXWx0t3Gxb+Y0
U/VlHhl3KxiRolNB+3K3ILvREyrJbC1dotfiU9r/BTdCxuB19s2gf1pi0xT5k/h1Byo9Yg0oFavU
qh/D6hSvj71G4CoahPGPpS8HaUlvTNf64zmN4us0arFOhewV8ofknIxtt4AarIypR1zT/f37Mvx/
ZYJ/6SGOjDVriFNa2zmWL6nDUK9kjhhQ/SG28i8o/uSixTM/rz2H+kWF7awiRoz09E4Bohs4Kebx
6+SYqhB/czlGGlC2eRNCFD8ZOsvuUCLHkCaSJaf6SLU6+9wqS7u/B8sPnWW+L5jgbl2U6S07IfbQ
rhwnhanmCJYZYemFBSrOvy08SvWIz0g98YOhfifC+4haqVthC8CGz6lBjNQdFyWgixMNKu3+22ZX
d966uOvxJdAnjA7vN2iFoaFquSRZVC2IYrYMOGBDa43gNt5hK1ZMikNxBoPK8hQUrNdFUwEwQbRN
YwA1EhlLZg+PXpk+pHx2phkQ/uzaUlXNyUhwLlBUbE+ItQmslISabfaCShS5IYKeTMG3Yl3kW1/V
uWSaV/3VyeOz568R+f5Lo38INaAZ/UQQ8GlOuNH16xHbFUPPdCwoUmXqkbq05DqzE253sqP+KoJ9
B78D23KNWp4UNOy3PAUqjYmx1+Ppwu3seUKMUiLLItzXi9eyRf15rPAfskV8ErjvvzuIxuE6hejF
yAYWh4Lz10pAjnMWRrY6Ef1q0lAbY1wFoCaUkMO1eJNHRUGFQ/oLM9Ss/DMW9acMeuVpLW0IwvuG
OjJxr/mrg61S1vIWkg/ztBh0kc4FdbAaiJaf/NQ5lA2S9TFCGG67phyZJ9Bdgu3mkhZU+fqsr0yM
Extd+ztpMmHvN2cHV3CJaoK3Od9s3PxOEtTCnFpxKuOXfmTEF3SH8GZ13ALJN2slkXvvQ9uC2LVb
O1yeO+1pzceDO+j95rDILlPuBqypISlxTud9oKTH8NazaGcpUJrcGLdw8THRStsOK2Y+O27nmxcx
jSWLhLsZKZxuzr4yi+TohKWxFUtbZkAideMpNbL0rEafPLEmOBOqjmmg3H8dRE2OLnNJo/xtoV4W
UHdb8q3sqDUFoRXnYjDrsciS5yg+szksrC9BUH6rg0Umh0hoh5appR1XbASc84w6tlOlMaFLA/6H
H5cH2XT3KG+aYWzdZYebC9Mk0pY22tVSO2VicGl2AyTW3qFReUMoJvRzml8NzwyPSnG4VyxIes4i
2zhEfhA5VVvtWNnVYBsT7c2moBmwj991wXnj8s1QEhO4o9YAsKRXAqZtozDbKmmEkMCvi91gRDYo
lZdUeYKz4zFCwOitMYLsc3S0Mkq0/1Qn4NXuph4xYq+/Q/Tkhj8OUfMehBmvYjpgb/8At1jiEfgB
7bBQzeD6uozUQjmLit0ktR73kscKey2kOFUgqFVlL35VB9zTBSCNTnIwQUtXPWQ5Iy8JXe7a2S6b
bPTFYsYLtxGuNkuXL3WgUh4LvvBTQ2wBidSpYmxN61gO1/AVN3LWaYv0/lRs0T99i3jT5zxW9/Dx
/NbOOcYylhIst7eQgnkWmnsM+4OQyZ4Y5Yt8SlbCQGiDqjhVrJD0pArIopP6itddmp5S88aLvQnl
zHQXgg/gbd/DhTzjes9X8HYFUuvLs7fArSQ5UZkzt6ntU5iBUacQONG2CZzCH6QvePmTdASA5yvz
3ULQqzDnyIQg1Bsf30xw9kPZ4g/rWNBVJncr9VRWUp2WGOEjL7HggvOUIF+TSDq2FfQO0AwpyOeN
YVPJFrhjFEgGguOIsk3veHl6aeGAM8SQ0BqNUvZ0zVKFdj4vJO8fFNK/VXoBcLkwShEwgvMeRMv7
INK/Sj58QkeS1nS7VTWVMpPXgXY5Poyw6mIcRxATJC8VLj79y0EI8KS8mZ9HCLu7ciLwT30eDsBT
1y1GTI4qXo8SESMp7XRG6XHjTzbkGeLCk58nDEEv0A0L2CQDWFbQbYQruxgimVxBjSBysgnh/C16
zGkzMu8ZBwQJZnqdJgbe8iJcrQ0E8RTCGs9n85WA14ae9QU6rLeg6ko5IWUJS+9qHUd0SArW4gfh
xlsZG3pSVE/D46gotkTUObTPzuEgZOxdnmHd/8oMFAFX33XZAnGxDvkZ4n3psNVtlzKT+JqPAqff
iKorLEZldIEGVK7UIWPVioNVVwmjTvoyOZXu+YDavfcr8MqDArPLzl1peZnUIq+gIdIbyOetpmid
FOscIvxqExccfvfuPrq0rAm7xoymL3Mbgg+t0/cXkZel4WuGZtCuUjlu6Sz4MnKDw90jgaM9OdML
zswQfyx6qX5BmoTu60d9T5mVGn3K19gM9fGUIzYHTrL+HkwZ0cCeRcb5LA4Z3AEHuZREiv6wbKjS
JulDGN2o0JagS1YVLutT31jCwuwPpUsgshp7IvxVmiJ2YCEHj9OEDkc3TcTiyVMOwx1XzzqMQvEW
/DomRYyVcHm0ontULi26e7mVyGdytScPReCVLlzioGeoTRU9s9OyqW/6qLSK8VHmHkYPVNREuKez
th2WLFMHTEQZfkypusQFi6hI42NCi+Ymm/nQywDPjhWS53vTgL1U01rcjaf/CJD1m3qMVOHrzSqx
unZnNGgfXWVFuveFjPpmTuML8AMLFl+OW9SOyMT9NMz1MgL+xT3N6tS1LJwMHjrKRLkYGXh18j4E
XxnJJ26S/XcZKCch5hSTRLMDUUBCxJIH9blq29O7jjYPVa1KtWekwEDqm9rA9f3rKPIxbMAY2f2j
JaXDwdpFUbm9pJHnGRMQkBpRrukKWaXh7BWNiGZm8ACEgVUnFK3zfNV/s/pUMbK/fR+yRTmcpuM+
1QfKwwsMDnRw9JEtA/zpYeo7ot4Ta8nKTPnYVdI3G2JjGSBK6yd+rDYyRd6NKjoCO1JbPaJuH68P
YQcWIrNA62YlrL19r/REInVe4LlDsvCsfoLDTS4tKZxpTZeulE7wh0qUgIsJ4nK0FDkk+eUbJfpf
kubLJKuzFDUMW7nA7z6QM8VdcKq9DF/5His8yi3im7Ssdt+aNNoAhT/lNtrgXxY2HMCFBn8WVQgD
q4M0Ij9yMqDKjp1bbU0TPjpuKemDBW5tE7rKZBfC+rJocmewC0UOb8IAsfkLwcV5yKsGMZIf+RJi
PZXnmn9G0hYtwfuocY05wr7ShgWYMfwrTtVppmN1ZHjSNGjckQJ1buWLKqMvw7+kyv148VFtTSyT
GMlmnxNJ7i93Sw1J7quWZCbcYxhy5HanpWqJSo/7mi1VvQB3swr+f/4U0AKxKfVTFyAgCX+KqNbx
v4yodoOb4yv40n6jpVp8gUdTvKp46CUvYYvRSVn04PmVxf0N07T+Zqzpu0PKBNL+K0vnir6GPFns
9lyr2nSuFEdWBHcZrQ90T+KAF5jcROZijMBRiXrcCKLPmRHl4x8Ey9EJXYhkAwn7iHnR7/ipicDU
1B/4N2ZbRNKzCopQ6W4LwBjWHMChDodzj4arw5K0AFhbVQII58ZLD2jnujMAL0aJXkQLHkcRf+i2
/iFQ2uS18bnyfXJuqHL1/TCh24NLrWr2YqovuG5kCPHpESmUpaaPBZMVJ30KZisM/uKGOqbhLGro
pf6FfMQLdVlCs2i01TCzVL5vknYSUlWfsprC0qJBwWEGR7F4sLj92A9ZOInuCaBgDDX58bA2S8th
iBMQYIYqFNGdS3F/KduyPOYqq1QCqvFgvo528CuGvKepWNEK1s/7htzvhPI8zfJyctM+xbpAi+E9
WeH8tA83/cZQHAkH58K3NVpM/rCxS0dgs0VFoy6Z5Hrbz8ZEL7Dys2WmEq5/hBxUSflejLSPupyr
ki2n6z8S/9P0WeFAFE8hfW5bnO8HqA4WdgEKTssTjm5p7jZ66tqweyZKZCrGWMdNX4TD1P6iQdg/
OEoRMIDZrNYKfgy5S0EouwBjoUWPJHgmp82Vyuoet7+zqUzWTXLqnli26wawTq2+bjh3sOC5qQzG
UxIEkCQkshFAsBySQ9qLEwgdZoaF6i8LLTDEmaTf5NKv3Mg513Xe4I34hsdPcKX/6j+nPjP2x6x6
FoaSMVQCHlnM4H9uR477dOWFrCDu91sJJOFqkDT88zmCL7rU1F9KnKf7BIGHBca+XOUSAbLISeve
wtyBkVPekk3PGQ/MdPNvwbWLIQ6zWJNgDhMhNO0gCT8r+N7kVKpOQMzBWTC1JkoOhTn6KSkpg6jT
pxFAfBE66AkQeDS2e86Yo4dkUI5srTUQ1X8cfTIqZqUZ8FK86g8e8ui8U/TF3zGmuU2ptRD9djr6
YDFvvQTy551jjIXmS+1lqzqSg29OgLnGLzmnsjLdsl/1XSIZaG4nJITixJB8dnZGXMXhcqCEAK6C
WgPkAt/taeX3jUAC2ktxGVyd0FwLpo7Uqo7vVi+PDcgOiRfD6J9roYbttfBAA9DElO59Z8t6H42L
vYYIrpaeNgvb6JGErox8I07jE8y05IU8ZjvK7aqPmapExJclrQjt95WNv6XNDU1i+THqpOv+5i2H
zRrbp7HZyCF12dEHdz2BfuHmtwD/j+BPvSqJzg08v4wI3y64blS5zDGYIwvT25N6YEgSyZE8L45d
MKoPyMvfx8TzZ8WTkiVNVDWIKC6JczmmDbGteGq8qzjiB7dNDWMgw3lJ1SL6ME2bMmoY+SpBktHu
KEnxshMs8zeFH33sLY7Cg5Sq4yL2f2xKGiA2gVh+rqm+CV363fvaq0k6hQ+irCisTDoGLOleJLWG
9TNYYLmwgNpWAbiIckvKLEJT7y0nXTXRa3esF6YaoMkRbXuq+3e2PWSE/gEaKw6NveA3m8LOzmWX
Py+D16354gDplngYAAkZVUHGwoBIOkRc4aU6oJEbRtl6t+eV8HXYS8PXCraQuhul8BjqzpMzfJWz
XJE8UipRAUz1UjtIybu0v3zhHAL8cDlCMcvjP2QYRzPWB4hKFAbO+Di/7dBPhe3aDCbOqSvM2V16
NNnfOf82APzqrnClyxnkOEpRjy1v7pbNqq/VWjioRXqlICWCAsAOo+uZ1rrP9X10/S9sEjcAyjdb
8Rl7RUvuwJEL0tLPpkmdg9qiIxsfvHrtGY9N50rV1TkN7l3id7VYkOi76ERGKXZ/YvQJAE6QHcSU
eHqSjZHgInRc3QXWgs8Tg1FF1nEHyHxxgn9Cy6cMEzT9vA03rHp5yvHLnMr3QvhaGyXXdFi1zu+5
FpaeIXFcyxHjXMLf09EjIqkPiTo/f3z/g8ftoYuP1RM3ShxRFLFpnA3FqbiM4G4WwseW/UK69ai8
Zws4UfiNLDeUlxIsCSnIr6PnmqF7q4yqPO9OHZD1MPVPYSr+5QYqK3ZRvb7su0E9LWSIOi8DyEQG
Uz7wixZT0KV/TsMMQLcsA6rHRjTUZveucO8ry9BjLnoqpI7N2cY5E0AKcelzhosob7IAcmKasZJR
ml7zvibKdqEOclqTBmZ4o+DK1bUKyBQfjW8Kyg3ge8ywxn33jv0MmJCxb5ERDTSAVm+JNw7Jg5Ls
LuU8pp1QfFP1VnXA7nOAhLK6TYT+Fuu4lrfhWKzKoIaHdwtMLVFNqXSw9vcPuVIX6ZhOFNHszcjL
oQ9URy7UEFe/Bc7HRyFcPWSD/JTc/pUDsFwwlipsBsNhOv1WaWxAefIowD8vf+Uu/PzUdpVqfD1r
cAccJ5RQOabXbjdHkNf1Z1KP7M/gP0e5zWP1VdGXTyAhlSYFYinYNK+4TnPxc6XJZ+2ihvtZedc1
uKuoQsm48LJ2BvLQP6oyAJ5J03f/gC3QCAnfItK1GPL/IlwUrTTyGuId+T2VXUr2OBKUafgniHEd
3pxo4AaBOPuZ/mDyaymB0kPpV8uNXeJBLeGLhcnoEtloZGBYJcGOvWqkO02vEdqZo8QixWdd9Icz
4E2b6qWgARlaK8KT8IUyEeyv0hmwmFTwOwXqMlPjfMthT9M5xG60rU1aS9h9YSNECfEQ6X9P/NTz
yt53Vhk8dJj5dZGg1Dk4ioVIDBT8ZByIquQhZmPDkKZMpcgqGfKfbD+tR8CUP7OLZ07n4OOukxeM
d0fODNsPEkcETDaRGRksFUGwMewEQNinnyoGPRPQ8fUDHiEierNllMohuTnlHArL0un0gHdSNOm4
amzh/hsvrzkYpKt9bdoeHVTNm1i2cUEVkQBabiAJif74S9cgNjzv4EQPnMlhqM4JmDJ9qjYz044Y
cWkv+Pg+jvR7PWDEG/PXVGJAHkY4tbyFNcyV35hDtHbL8g1RDS4JOZhJ6qKQUqVVRij1RCKBxnBM
6mHImAa/+xGKUk0aYlpwhUtXbLf7WJCpy1tTnOA64q+OpwBOgEd8m8Ypkare/MK+TGHfTNDSaLwx
mcR5jNyfhf0gNqN3UlXOZQxU7/0ehnu12p1Y2S5atlqkIKLwE8H8imxsKZzvAckk60cX8W72eANG
AO0YJwI09gKd9+o7o0knHvP2JBDVF/ydmq8PvvILpDpMXLCykk0yW/t8yTSC0ij3/ZrL6rVCnGCU
VX7yTkwskXGj5de1o2h5fdp43Cqi9YRLEeTvBSXXLnw4S4yRjNdf5g41qnH+eVWuH+8BjvlFqFr4
EDCj29qeUbCLirzKmHfVVM2jKP3wH9TdzmjTkjx13Dj2caGbrQorj4IRBCoUuLsjGVvXQbKACJJZ
5OxjeS1ehWXqHrZ2Vna/QMWxOMIbiwF09hMfJY5sJ9e9NjQZPxDl44c8+gNSuvvc2ZjYjIkBkkv+
eJqaHoh5on4r+Z5EurJax7tZ7c81zPv0K0F2ba7EBYIvhC0AVtQmu7iDYZDL9NfRpcJBjmM0dFOM
4KsR5XWu0T+UhsBsi2DTjBOJEYQbdNB5A3IpqaxZgHcHC9Avca6QhHT8NZr5PydHpyEoZKXtuHRQ
vLsFFVKgQtHK7E7YQ8k1e1eRqSbJXMFGExqOE57mowbMCc1inFzLpMhqaOQozO4QMhzVQMC0d89E
Mz2Aaf6OroSiZGVWs9TXCGrhxr+OFI/c3YwFjCRr0+xp7I/XGPWiDnfgN/YrPQKgLEdAcZhBf2u1
usUQHdA1fJpR9VJzUZh70KX+xe/5bf6Lwzfc2M/97u9S/3nyKooVRnFiuuvSCz4pMSErLDyskP3f
o5HkyUyfvVD5vv7qGEQbzKq114VjQKqhBzQQYMDZLQ2+zLVforikT2FgUFu7C7jR8G/J3u7FtUgs
NnekMgzZuOmv9FsV6wt638vsP1FIAYuaSpwdals2enz0q9BD8JMI5G5E8emrM4LeYRYgYeLw+kmu
/gglTKFAFxqRDsOHt/77rDf3WB0sVt6hIgC+PvjWty3DfImx9QvUH12KSnFKqI0uHKQXt8DXt+/g
xIULM7uOxHplh2VpsdlKPJaM+3I/HqAFTQJNVlIRgjfziru9S4n0LmFReqC6Wz5qlXQDjy67YYbH
7mm33fOT5h4UrzbCIdxgSNstqSU4TJBa3JEtoAD0
`protect end_protected

