

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
XZtM4bLmkglBewlWavfkobXOIMkrnElgJo+k4jE78ykb7oIZp/SGV6Fmfr/ogrusY/kHxxmgAde8
wVKEHfi+cw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Qj5OXRmuDbyb7tXOe/IIP9hVzpHdYEdnGFMGPum5TPAz9WJzfNr2HnR7yYGe719tx6wYAvdRlfH7
1KYaZqML4WollrpclochLq72pgPwbtC9iEEWlamVuKdvYSw0+IzNRBHdKqTykxKbBvXaQ7+UOUjw
UnhOWIyi6vA2XCWBMhs=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
wc/9BtL9LkvfKqZJg7KOk8nPkSL5jxvAGfC0RV814LDUHBZcOVMBTQdouKf45+uYbzuqQuzhrFia
FyTrOU0b+Dpp/D8a4O6aOPezhZlqDF7SuDaIsbNJNkVeEPTzKN3+pib+HJ+07zD5sgOQyBLQtobI
4fQy7ggQ0o0bOrWPzlXO7kD45yraaLu2CaLqYlQzcDjqnvaWtdvg8Q6aRiloz0plB7OdNZ9a1tRM
Nl6v3ocdKRatScwi+YnBgJn5ewXMvGYuuBOXAkUmcc+AFWML9u7RnCLEmrft5oAR19N3inWP9hTR
9sdW8LGJ406SdzZiv/gZpUV5t/AFjTB8Nihgew==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
RuHNUBMTP+a4VfkYIP3nKug+Q6Ygohn4DcPwrCybnrM/u1NLZNct3nJM51Ftp2uYn4LtBCAEFd4j
J1ykZQnUjNHc8Om8TkpAk8Xoe4lNd9c07VFQ/PdNEPsRZobFbRhtaTn5kYtwFZszGT2+NVjW60i2
zzHWmeNAYn4vMcnLRnc=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
M1UhZ+OMYDjkT/STr81dVx9PmVVG5A+2IqAmn0405vupx6bbRZIy5mB6w+gLHolhJXN5SjXXAhWo
hTPhhYqRE6WXBSt+aNme9SGwhhYQCQHfdP7l6de6Oriyjp0GyOVTMXW7th225i4gd1/MFzrJY7uC
eTxBA69zF+OCz0UpsBa0iiqA6SmkbUtST66y3rCQ2iRlo3MqgxqTXadwVQPjyKh+YrZv8hSoGQfZ
859BObwRsVOuARh2h2mJuicqAywYo8mWCsE9MJAhCYkJvjGEbdjUCSpq6KjZZuBtdg5UMkBgdSnW
7odTSYiZWcCz00u/B4xtOP+tFTZhOrGrUTKipA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 81744)
`protect data_block
qs92lkZ2njw6Vnmw6MgggCoastwq7wJxSHQeTqE3MihQd4rlqLmTXjwRko2kYc2RQ22Cc6eNDCkW
yW5vK8T+IChOyes/w0x5VLMGELOCE2iw4WGqbUwHDCESXO2162eRPn8NZ5w380m7jAVVTNoOdnDG
HGS69JJkj52gRDhJTcoDD+ejeC1VwiXWNimVadwphWWgHeHBJpqBzyPBDhELKDNjcyyXmXq887Am
kJ6DuHxSMZbDOPMBEzzMoS+ZWW45PWcIK4WzDM4egVTdqEBheBjJ82tvud+ERlfBPuROcyiZpaqk
XiA22zUAywMnh7tLChsUcHrhyXhwXWmZsH+FwsfG3f/jIDtsn1akqzYCgoCh9eEHfQkZLOwWRj94
Hw0oMOqrjsXepbWOI+fu7vkGB9Ndy9nEUgksRd98sOyS0IrW4cs+KHckoOrCmjv8/rlUMl4wWviT
B4g52jE/Ml/bFMMnSg58aled2qkbegZ3Uq5Uw/thmFGIVqvI6aq2zqrLnkBXAhLYEZZfj+cTIVvm
TRad2fBOWGh2yGBNJHycHKMC0bn3/ls5lxrn27I3YEY4KY/IfJU1dR58snGL0NuDWgqf2LmGmDSz
sSxx6FtNUBpu6M19goNufHrDEtJPrn/UrqGSufd+TKaV7pE2dy1X4vs2YpRWCW1hgQBq2SbRXCNL
J98lW42Czp916Ggaa07tuXvo4Pk6VUXfLz3af03bBHBvrR2RESWnMdYtAhwfLT49LnOzR5OW20jG
UWBZRo3bv0R5GRoICzJBNh+TukgQVyUmgfl8xe6kcjjjrSjzLPbmHBonUD6pmpvHktTz0xvQfMV3
YXxIRGB5K5lfCCNj3YXlKn1SdSy4uRxHzhodt/W6HR2wm8s0h0to7xPwY58mJeCe70HntDE79qA5
yeIGMaJb00M/HQyF+F3vVOjfGEOSxYhiGLC4B35JARsGZ+4X9cu2rPbOHOk7dUW9SEKTjvNrxt1R
kkfA75C6KjMRBR20FqRICIhA5MKiShJfrCL4XGZbErxfMd5dlwRQsPnmvKt3qtGCh6ip1vFfGCQI
/PVUd6RyvJcP8Wd5TrQ5z4yViA1WHeWfLpuFberttlyrZnMN1XQK/Lq53SZ73qzBcOo7KDYNmEsz
4eQHyHzuy9ULkKqTKtiWKOToD7hEYgjH9BOOKFuwQ3XDYmaPbhCFFHqbN6ixUUhCW0qIB1W0/Or1
cq/E3djj3HJUi6EEqcOqecy4u9oT5+AP+Uedem/r7yj/hcW1oqcTFGM+yGlD9ZMQP9MfMtpvwEKO
cSxoUQMPK90l6uA9h/h9on914Cr49gpTbImqxBAqbJFlHCkFpLLG43bExh3kuzAU0tNflYa8aKKS
EZdI5ZaIRs0FuU1+/6evcnWyqOl+dB2ptgo4uRYDAacEjeX4tfhtO0j2JQS5lsPmwGJYzClmhJUI
Vi2l2a7rJeSOFuoq5qn2tyZiaG6XG/eI5rVV19VSzKItoGEGvfGerfGujdo6GYG17J2AxAk2o29u
99m5Mz2mwNgzaXt8aS/DqEgsI6xVYl+EqmZwZHJdNmdrHiv/g1nwIrqlBw8KAvP5j3gn372pNj0C
ou4USeOLw29Q7le5crujtvAyRlgznFr0H3ExE/G/IWkndGR3tUJqnQX4DBr+mR+ssLtLiwxtK5Af
zmCxqrh/7v48KRz17b7rkPLTp6iHgQRJd7s5r0q9yoo8t0WG1C6Ul8s2Iz6/bgthMBvmcGL7+5TO
o5E5QYHJfF/cUFgifZxud8+hABtyapbNFWpMyRCWoe6sOy3z24OIHx+afljex6xbUpyiJyBVbKgj
urULjgsEZAvHOg8PuvNga1MPKlVAaysmKpsfkgyumE40gZWAuab+j1SjOm+Uu01uCnGy69EaEZNU
TzzE1q9G6Ksjkat/wCQbfS9KsDTzSI90dLJeCh8FpW/+l2qTWpFOogQWCUYGHQwPVTZnMj7aJ6wP
GGeVu8hQfvAFpl7u6fe69TfS6e6fKRgn7llhhxmufvAKlroRLJjTrQO0qcgLjyJTlZGfa8iw9OGG
jj/YjOIHPNwRoqiE+zmOr1GHj/wzOR/48zWhT+OTvcF38kwfor4VB2KfoOmliD4XdhE+9E0YAMIi
2IRCggujHm7SnMpQx/QhSHTQrZYYNwesil4A+287rrPUUf22qWMqvZe0tER/pfvWd4ICRvsSn1sY
MnJbkG+P2Udcca9Sf2mkfwT5xGjXWjKdw6Ve8P8ZrhYEadDPusTebEgzlTDpwxu2fIanEKA7rXso
s9l1lTm/ZwJAq9O1n2//krdUYMnUmwoXEPkKiXCYecTWa75Obwg2S9Z6Iwq/vGwm07FE3MGPue4K
/AzTIP3SAx1eU83TuJE1uh+nXxHc1Soytyy9qWJusv0bevBQT/ICKGjhYoEdowuBMnzNNIQ6eOkg
esiGkCRcNWup/z01/BiASDxtesUC03nmnSSh5hrtGOMObD+4BZ9HuvPaVtdosPwxTnXL6LxztAu4
+jWF/tC+L0wih2Yv2+aQTzfQGs1EBBGU8PFR1C3evgP79RY6gmG45jaFk+g5hKf/zOqNoRyh6vfN
KGXJS00o0/GGAE9wF5PDO3HTUdGa7adxAledKUXaxbl9N4FU0ZJ5vCdCxCt4nP3XIW0U4HhU2T3x
0GFlBT7ULbRLf2rwNJ83xX9E9i6LaMokk32EbgLdDrU5eTXmFucl7vQX9DYr3xp6ZbXZnE5ou0D9
oVQVUBqDidOME2kay6KBUFkYywIhP0BHmm8Futr6Hd6hF9G60qmx1MOEYLmHLVMAPAtroeFE+/tE
jbZtPSGQGHfJWZG8F9CfGwm4DiMhKe/vFFlc4KmTfy5CVAj+ysx/lnDfknO8TuhYbZEuLtBxqqK2
fTY9BcIAfPEj59YekmCz7tpeQPx0vjTJq91kN4MtBa3ZbFV+U+wA5NXaV3q5+JZVcLCb1tg+h5SB
j/f03LIzB3JOJPJoFuInJrzExaVG3YWJvj9JaeU6qeE6h/v6Xpydi6jGAYmsEimJU9IO09wKFCwP
LX8lJZsqF6VPwXZgh+eHq1nKSuihFEvnMPclOoqEaQDvsrGASN59BFAjrcCKx3UshveSNRuoiRCd
bFPutFe/2GIJAH7ZuMfclmiG/8h5jqPr4WWkLXajFdeBp7tJ9EKKripwDnNm5jLhSR0lMp1a5177
Roaynwj4zg/RCMZX2ABP7AvjqcQaMKm8T5ZUHHiKmJcAtokMzKk0fMLBW8d69Z/4ZiTciaDWqC7I
an0vecXxZ3Cn4kpJlLHV7EMei6KT7Z1PuR+Lk5gagT51WbHpOAY5PYxenmdGu1/+FVLxrpp/xPUL
TscCUsPDPuEwaA/tN+jiuv+GYfF16825NK9UFtAYrR372FlPCCz7/AIL2VmGnEyM6pSA7YHdCEf0
XSktRchr21bTi4iLqnHFxIdJzwqDK59KQdVmJCLSDc0QhtgexyomANhhbsUzs86SQAzMJpWRgL8L
5DlyqsHa/9qew8XOVF0gUEPBSbwAND1ST8VxCY/sjzhjdVKsrO4xyflHJdveKYaYlgsiHXuUeHE8
bczo0ajOPlLJnItmwD5mpatSlkHcK9gRf7VUZc3e67p1gFs3hV4h/LGp8wzw5x2+p9Rkdz2zYxLd
kb9GzpHFWMLVZy5Ct0bv8h450kqlhSW5meAlJSVHZHxu2ya0wbjTSS6zlUIkRBRosy/TlKQVWqut
rdLEihcl5Fput2RtJH6MXQWKVLcumJIyLZV85N0V8lBE6g0uIzhPkvsxTArcLXD7k2iC50xa/Z7E
SHYSIUAf1IpwdrGYIH14acXXJgyNr1lgnjK8qk2FR7Dnl2wTyBbrswGAHW2s2w2JZ8ctVx9sTzHh
ZxhnW6USyupifH8FQo5Qii8isbHjgB9I6NjXXTVIY5x9SC6UTRhAzgBF8V1mRJM+afD1u0BnzjyE
zHpuBqBEfGHzlJMrc3MS5TD69iil4xNbck5tLZ8Tweb7LURSgIEWdD1vTy7g147PqjXCQ4pPp9Xg
brK/Dpf7VOPcF58EjX5BBBHvqTl6dasPY1bjFZ75tAf5EU5u1Wog0PYFyTxuyR+13djWlZYbV5rP
kUxY6IRRZIuEvZkH6Jr+1X/PFknV4Tnt25wZrqfASogKmu6uR3gE9RujrQg8UyauHgfPJYERtw0i
ewueQfBiw05ANIsSRtgcfXA/p5783qkm2W9nMw2bqCMYO0zJVwrWJZugMwKqVO2lSAj/Sly5PNGQ
gNbH5mnic8CLi9CCDJk0T4Vnw8e4uJ9t99ikDIVsNGmKLW1xsOMY47IEEXLcL7aD5SHLa0v3rX0K
5K4Yi11UIj9BUcrr90d0V3a2Nd9twKlde/CH5chsliw/RC94Z1hbaTEgHKxcJ8zKUZ6oiKcOGh4f
WhL1V0D/9YWlMR9hGqKjGQsw1BTaPmBsA4a6yPOfg+9VXClrd09FeEEoC+mmeuSupbgM4BadD6Hr
4Yi7W/0KKIjs+Ffnz9OgCbyrTYEQJFQZc933cpx4/w+BJMfPkVZZay3khbDya+9AI51zYUNWQuG5
fRrVlK1VKt9rShFr4CpHMJ6KQyhMpbkW/ySCK/XQGUXaDCojMWhFMC+dR7J2FDynEPSm61RG1HFz
v12FgvpC+jfL82U20sDCuuLjBFcoDouMxDZdHo+7BbfeS7h01uZdKAaGwzGyihkzqeUlbsK4gFyy
oBwE/q1zxYXq1jFKahPNkKIoj4+t5tgEOJ3v9zqGZuZLm2x/38K3G0iTaVU9WR/McufWQALwFQPg
gPzW5rwVUnnFGUoxbhPTAgdW0gkv+J5Xo+FNeIE0VKsmnAP2q7lSdnaw7t2LdyhNCrPg8YmYSxZp
OKRjtrfWiof0UcD3ypvRVn7jQ/1AE1gq9TbjST0pNuK6I+I5PR2WMasxlwsC4zW1lPuhLbrFgUWn
sAttcTJ6dYiGAwwqFLGpEM5MjXyg5jVfn9uGKpdor5h0+bQlSQKCWAL4pcAFJ5c6jIzaNqwlJIcC
VJSYYUTnPQMqzRAZrjy/fXhznCRBOkqmUp6IzJpcAgOi9pmeJ2F/QQkYXjd+vvg3cTc+JXJqOQti
kFx5J1rFPZmVS+ynQBCWTd6v8/JfUvw8XbbMBfAXi9wiGcfDuIMz06xS1AJRih85xyr1dfggoV5Q
hdbqCb+GGTe7b7x3d3eDRbM8NQjeamu5ahQIfcv9DYN9XcIP3AePw5dVc05D8tG04TCoImrrlbxc
T3hvLpBxYscy/idKx3UvAoUyfBlKfWArP9xPtK6ZZTJSkh/7bWS/wPUqg7cUSFGB93mPj2b4cBnE
ws6i3I2kPli9qyhyReRRg979xsIGWiT2Uv/Uzx5NgEC6qAmpSDX+J6Dwc4bn8oldAuX4YyfbvRXN
qVyRr4EEMwuqBCNp7QbS0GZVFkpJelQNdxT0ZypS2sam1GRwq8BTA4GH/+0m5uSZ4CcK5EKs9H7O
eI40Ogl9knWg6ySm22NU8tfM9M7Hu2RnsY3iR6esvq/YJtkgyWqZqAun/XPNIJUkC8omMeUAAekw
+BBDyim57Le4yXy/MHs/TAA0VFnBgaqJL4Ba1+2plsrqgp8ggMN9WbwYsVN0g7Ey3WYZ3FrdKgA2
iL4d2LBCtyhF4eVApazj7PohXXX94glnQlaRzJufNFCwbrxiwu0kbFFbdmh7HSxBupyvYmIxCy1w
PI0v/Lygl/wEbayApYsaiA/GE87tZbxDWK/GvEe5swhbHk1pRw/02cfx4aayVsm0BZI320+nGOxE
EpY6sBFhuKN3iFfMC6SR/q5rGBQ4gv7MgL3dV2UUCzTlaN/Kkqn/eYyWVavrbFoirrDngCSpXtZi
aHxGAyTpFMACe9y57DIyj6OSFS4zaGiuYuoNpw+ADHtM8aL5hdjiKZk9ZUCPaciKPmz6FZ/SlbEx
fnDCtUN/Dov+z2gufrNWFODDotCwYJAI2EX3TIFDQyHfUkb1b2u6aL1OqZkQ23qOgjaCN4jMGDnQ
K3Kv0GK+MFHsiCMeNcAWIyyVmDggKQ3Zp31Nj7GuCg3iSgIKV7VkawZ0gAGGLuAhKRMR7z0cDPvH
zHIz4/Fcg1p7wtSba8RGIPyxFZQODfWLbHHcoDJwoxIdYsra6CjM+7pQCd3+IijXpuNKPIpUh0lG
3fb6MaNpPJxW3KehZByHzkCh89JTOLpMzkKBGwAZMMH8Jkc1DI6UJvtRsffPaN3hDsK8brYNK0Y8
SU3tA5D2rVFMNEhzU0Iaib8JB0MlhtfoJqVzFlf+48BYgMkYRMlMowdaOaFRmQ1eenb/RSkP5lV+
dOtZEyldiOcBhgbG9FSHbpt4v8OXPLwZzuYt1AfugvE92oUkssy6PNBVd6OTk41YuzK3KUWiY+4P
4y72LcUM+onoSEemoGr04RUMwp3XGqYGtSXXO6Os7KNn/jpCrX+AekYMhH+5/ySlSYkfZvpYDYOz
jjXEqsDVjjNv5ovjj5pCvIQAl3xUawIOMrGSSGBwgEHnCmJR/OyMLg9LPB5z6yNFEP+fZDLkGiKf
YxaJdCqlwuavkV2gsklBWJivUuPUltJwVkwPTvGzxxeUVMTgqLZhL6yWmjpbqCnyp5D5bWtnRfxj
mu3uyQ0yamf/SN6WS65Z/WMZmxTb+PwkltUIdzaiBtOkUIDM4bbIA1aX8wQC+oFEyvPaMOz9bpt2
mydTiiAK3EWRIfaoALyunsRNsWH1cks0N3aHoAhXrGrkGa//4DGNjbcy94VVRsiw8HCnyoZKHqbe
ueh3dLGvAkfEvf+GZBoDIPntEsFnJsSKtlYYg8kwFI/AC/bHkN3Xek1Yhz/hl2sWdOj3wnwylM+4
8uKjBaZB12JGePoLM9a/d/JWL4TJ8s2KxnURne1coKhuonHurE4/vZNgHQapMSk/pO5PksDfzvxS
T2lA5ZhsBsmKGL54ouO8vEbMZ5A/mi+WdsUH95Ts8nmCRy/njoan3ONeb7EOGzEgw7mi9f25cc9s
iiH0War6IqNcAFtd14+6QnKqblVuSPA0fF/+PN58FDScZODSLBogkk4BUudNdfoHNT06InBwAKJZ
SRWRXrwWJaF5wt5ucU8NDe9MT4u205Z+rDMoXmrf19oaebHXD+D0YxFBGAZlheSLQRQabuR+C8NQ
OR1+r9zv8+pWAaFovA+vpHnSmmTzowsvXUeCZpkxdq17u11Xyy5rkS3hYcDgm7c64WbTm9pRSOtv
yztUlzmaTqc+dLmRNdkyOrcyJiXf5NSp5jVauJsXQSYaReNTsXO42Gn/2qtd74hTKLpm+XbEg5PC
ryfT3GDSEXGzMgAE6KbkyCBly7nTs3G8JJhc4Ggp1Jkpbthum04SxldNnznIa9PYI4HoI4ohAV3M
DlrM8DLJ3USsPvBsYtzNB6L6eXEzbQo8F/R6igVHC9aMRs0jn2vvDw909iaQtz/gqqIjo1PNCQeZ
3ZHof4MpKWXlIS4BEOD8SiF+rCvlv1UWEM2eNoX5SxiXSo1D1QivkwL/A4pc5GuFRjW9YPGwLO6q
JFOKK2xGGUL6WRrvCAfVy+bc3HQJqb7o28VwdSrthVjcXMRVpoydEHQUh5fCAhidtQBbFinRHgRP
aSqUsH65BEZbnAFaXIErCDzW33wYUcKTgh0n4hS4SBsqDEpXoek2kt51ewZZs8Is7lWY1f/zUANx
qp4AQvbqGLkHYSPGOn7x9kgC6qyEHiHohp3+6JyOh5Tzxja9pp8pmBf03vuQMPVuqqoSEU8JF8Cd
XUz2/CuyMIKzQdqvqWnYO3fsRZYn1+vbl8xCHOUtnor4UsmX6Hr11K4QXbNWoUEfncbmyoO0lTcQ
ufHw30inZGORpVIRLSVfeQC+n4BHlWxju51s0YmzzCNtr2r44zblLexXLEwOVOJiaX8HPUvCmMKV
R1l6VHIse76j6IrntVpa/qlSRabrRc9K2nwXFIER2R3QsbDnAzHwnuV62T068HyTzvQ07LZ/H9oq
Z7ieoChX/L+835WOxzJx0M5GfkcbfAtib1qbFo8qiKT6Bd/M+FQ5x9Gd0UJRdymNXcB3b4/8mzF1
ngngd9KFPK7fzsOHTsR9nGUV+FpArJ18BEkm7aWc2+9XQIUF42l9NU+3+XgQtA6TtWBbp0ovOAQ9
WvhsQV2k3HXbnKdf4+xheFYZLHi3ziyD+DMJKXRpP8LRndRra5zf3kJlfPod8FH2sYlmWLi7FIvN
Bwg+2lx97Lk5dj5k9PG7qFYek4ZyaB4aeEZm3SEjMkJeq+ZLw9QBAXRLQr/tnQFrGsOr5uEUxXfw
O3qRhcll5t9ZBwUTA8s4mVfSqbqmh3pVo758IFaDICl7oYRJQj1TQld29SV5jVT1RwNLcusj194n
5fdbPBC7ma+eP48aeR5jIXn9gKII4lLo0orhWtXshS8vea5jMufZj+VEPJIsv4wqT+EKDPquOnU0
3ltzR9IO8Y6jW3HXCkc76w1rU43vV/US9NHvpITUBHriGabEgK6wRwd6vqV86WmQgUHpHToN9oMB
uBqeYOtMkeyrLYLWzI9CQhIpRlEOk0NutnkrAkafGbd8v9Yn8ENfFhHn0Gansmu10fEMvibRKGle
PHiNT2QOTaO0eZCslAXftx1boC8HG5UFVvzzRXA/DbIVU2mtVNhn/kISByCNyTKI2POZoHhYk4fd
OG0Y7RB3CRvYcwLdRtJb5f9XjrRGPaOyuIW7LMzjutGrrsggG1h5JidFyc20HBrxidsNoASfPKFb
HMkaZLG6YxCaFCejB/pc32oxmIJXF2x8d+A3IX9AXV+C3JmUUFB/sGRYo3LJw+x74ntlw61e1tVz
7QD48QovSR1S06+Ao+UajhyWKPCWQH9vNHWbGX8v1Q7sFy44UtluhlGQKbIZ/BrU6GFw+FzRZJxW
0AFyZl/JJD2fLYlUZsxgU+IK2R+bGMzlc33P62V+10RJL8FWFOWBB0R3GxNx5w5BBfAXzSUxtK1D
9EojVLJdftyYFRIsiZA+08Ig400pVs5iuUjyqkkiyzDkTtbxkjz1xSG8IIjO12JCk82Id47UT56y
I08RNLQgscHLjUnCeK+4OxS9ERyEn30uNbQnNo1E2Npjf+zt4+Jr3GBtf108fXZjz96FRRojBT2d
FjWredS4kUwgUT/sUkgZ5RT5x5WBAn0eg1P9I1Dz7UYlVPVoEpxibftgnmbTiFZtMjlyNcWcKIA1
/S+BCOwy3gN7y88Yoz11zrnyig4iJcAi+F9xfidhDWOxuGCvXrJjpwy5H4inQ1KgyWd7WrVvihK1
bovzDc/kVevwtCipzS58B0VnlAsNde2zjJb6BDPvFAxLQefbgp/xB1aC3rOnYQRchxbAjicyKApE
8JY6UyS8xNb0Vlox8GeTWTgNS7drNEP5PBSZIxJX5nAgkIrBNkCggIwIeRrXe6TD11poQpAY92OW
TVivSkeGvSZYxMGsdq8G5ZtgeAY91L2387dh1d/RUoF5xFncU6pqrA1TnDkg+hJvkPYZdujwFMtt
Q4DxkBE/k+91l8sLZIE2Vgi5gMY+PYlwcH6vJiQXNaR/8X3jZXfP0k0r3SShnT96u3qIFwgLYnyi
+nJHhQ23kb7wK+/XNWb3hMKBglKusAff2eeOHB2iI9J6zUNUUU6TZ16cDmg3eRDPE/1SC7yYdB+p
zgvcpcL9qTlmpyr2wbEc5zGMK85OTziltG/NHUqlQwuOfIoi4JlXtxJhhgxyM0sQiV1R2YreKaIO
/NLrwRXXv7XA/dszTqGEUOQiemb6Ir8Mq8oUnbQXx4HM9qFoF3D1I5s3XKJpgHal5MWrfTC1xmnr
fSfoWOmhiyO4arjH8CAPlSJoeNuVGCFTlJcsDYyzGpTY1ewSB8jT5xhrc2lUjSJj5PWMs4iV30/E
ZcnN5kOrgOnMlNMTyZPPjdMKRadDGLur0M2U+zWFRcGAmqfP6YqnCq+SaNR0/F461iSdiaN3SOEJ
F0XswVfq3yau9jr9Y8ZAkVTah97u1bgoHwl/TYIL0zg9TvZ3vBKNLes0a+EYFZz6HjILsQijugRb
pt68lTIsm+2fMLTT8E1hyjC7G6FvgFQJ4rrC2DoOaFkT9PD3INqQBCw2gfpkqfRdVwwfGHwdMuUA
9POzpT62XK6F5WtKonr4EdEzNOhV3WNA/IiuLzKUVQS+jMkLziziY0xMpHdrQ4yX9oZROIICzJb8
wsVDteCsfkjXP0U+ilKUpPjapZR68/9zfPTjQ09/xgP1Y9YGr5y9NJzwBDJNFIXUhvwi6ykT408o
RVAOFMg1N1g9I2qjmqcRLFqAcKuUP6BSzmwLEIaRgm169BtkXjaYIzbBd/2hgn3rzVFkidZfchYu
j/AeQDaMuF2cX4LiapqM39RgvdHr/ZgSzJecwIUNCb5odlCO5G8ZsbC6afOTuPB9Gxe+IsVeTxYe
F/WJgr0ja9dB/EYKjyJjrAP+0VAWgK3Vc7mP5IuATmQ5NfcBpTTSj6E4ra2c6HuETo5sL09GYW2/
4Lh8Juj3zY++Sszf79SgMrhA4lKozAvu44euuUxLLPMOuG66po3X5wdmpfAU9rNAuyyPJPosWDjR
AYmTrU9GBG2Su/a4pB++j2SH6PjTb8NSv5CamjVcPYdp9gw3+PD7Owexkk7f/xzHOhzxq2t8syZ/
tmiy8bTtzXqNFn3q42ikS6Ugw9dHsEBz6NmbE8CMPnXQesX26csoDWQxSSZFWTP7TWahzF8r+Miy
yADMksW3rhMD+9WccqxdWXnnfAQ3sSaIP0lQkEm3DLkog5qrCBA1Vav2Dvk18gUCvUP3/4b2y366
y+fWxfV4rPCHf2LtjtOBlO2kv26yZTXGF8p5FRcbDYe6KRSrRq4jMcguBGCYKjsDY34YZINi0XIj
oLZgedsCGwmhm//XdwZFTz+1XSraP/cdCOhzngUB7oiuO2Omr8B3ziWIYzqWD9aFjrxeuK+11Pdy
ZYONyRwkllgVG6k45EhWGmOQcS8+Drt5mZMNoBY2bhXZgOjZLTtBbsh1sbQrWbXY56PkLswS7W5q
4uewwRV1MLXyovBLS646zEHltWDph23LL6iCRgQw6S2la12GZcaOfMjyIbpaWZJdbavscV231Pbh
f+veBEW/4u1cn19I3BNhbnN3NldGuxAg8C7C7XdjhjPIsBDM4EOLA64RWPZjBHL12VNs2aEtFzXr
6QKZ6BD9cbC/KX+xTKqdz4qv4Tr+NBdzG9ozS7Nr6//MOTKf1WuQCqXpbH5P6toFRjkEus7+1Nrg
vw060M90Ql9Ul4SmFx07J9YjgLG3Kr4UG2AOzhcOWdZ021uO8y7RXNuF+3ztqdeTJUqjALwTxsp2
kIQJH1HEitx+rFd/GZVtsMW6WdV+/78K0iK3wfMP48KfNnsElcJYnqhmchbrqNL5jNvkc4PI3th7
IsjsjjGn7gb0JNWAzQ9C9S3mnhIsY60z+kDMpmat5JuCWhd6gUHeWFF1nc0VvDnaCmaXcPgn/+W5
lRk1xAyx6BzNwPQtKdffvWFo4vy0Mvpg80wbjwvdUosa4wAtDKhodSxCAo6+9P2gus2OxN0SXJNW
idMQisue89IGhJEq8nfj8a/ezoXtX0+Zq+6Kyw9h5FNyH3cqdzUb/kvQArWtkmIy3g4xi6RrVAgd
KNxhrXGvxlXCSyaMj/hFtroy652aG1v+5eEurUEEVf/0tPXEhkQNix0byN39TUIR/UQXBwEGuuEV
Zz4599fEgpAR8GHTqBhN2cgFIwc/abbe/7qt/X4gOjpvOKlTff66ujiImPgWbj4PC0PKTHe3Lg1Z
ve2qkXkQEif+btF+BfAL6yRguIZPyKTXxY2aAh+fC059nh57RNsS4vSvMKVBgoJTZygJk89Fxshp
+01Ux8cECXKeNysCyrSbYv3dWnbpNDjAce66eIE4zCMExi0uEEzENBVzNfOIwta6P31tsgoEs7Ee
milEv7+refGisajtmtBMyWgrkO4e3Mf7nmgjqV0iPfNQ4di1k7KiXZ9C2GvbTiCaE0Ou40ju3aAY
Yp0sMk8xv7UA2Cbfs1ctzDqnhuuhl4ipoZ9idjvXPrGLxIJ3y1zEj8vb/0fBsOD4ltywBpgF3i4f
Wz0vZ0kMXo3JJXmv9BVt7K9C0Re1zrwFsHWAJdFkbXvdbKwl1xzDTlGiTh5YbkESnCTJq3W5UvWC
8jFqH9nUK6yL0MKCm+QKrkof3pI40zuOHN3N/rIg5EXG5vpZm6pzeRpUw5SeJ4ytapeRG/BCqtP0
hR3wd61XNmruXfqNo9Z6BUAaUYlCAnVUMVcnfQg9QV5JJIzL6cNdo5cBREgZno+8Wjg6z3eVJAgv
IgTWTwc8BpFH7FVEg9hffzXf2YI9ZFz2M/875pGX+opr5Xa6HnrrBqcCZ+VVEoQrBGbjAbjK0di2
jVZyQt3OFjnxTln05aIrR+q4WF3goS/DlHoXX2LPQ3cykfdGNJzJZGdT6Aj4CQ/MCVOf5b8CK6Fj
6EQ9c2OStSLYwPXu8Nr7gOIHZLvRvZi4KZohJc+zkYlAA1wL4g7wR7pDjt4KFQ1XdiEbfZKWlh0A
FFvVKmN60ZR1DkNBw0ZNsOd67D8xPiWC9v+9wWwdtW7SygyDu9LyetWPfmN+AL7ndt207P+155bG
tcjBebET7klX/n+tbTRPoKe2/UkXNADSSAVMcKGsFvtNik7xQJh3crAt+SR/l0uVS4GhG35PM0YV
xqOQFEm68krBgj5qX57TVRvdEVAutHTbU4i0r5RWVQxPEFZcS5RNn7DP68iANJLwwEzQdy3gqR+z
WHcfU12dtlNC5bwyB6p/3zIPnKmJE+VDpN/UoXI1hJIgmPBsDRlDXd8A382GPuH11WesO5CWxbHk
foo9G1NOSSwXdnfB1ZKXratjt5180TG33Udg9YRd0v7wPMzcCGxCBifkin91imKzEUaQGhJ3HSWU
0GqrMv/QV/R+Nnkz/sF5JBJr5UB41DpP0EtQv9riigpC0oRmShnGGPDaGd8apq1Qk4UEfEUxsUD3
b74/30l7ySQxh0trPOXM9jHkmp8ZxU8QMlFAecqYGGluUX18ekbAxBXQWBkEnhv8rKKdUU7otkrA
I26CeoE09Wu9I3XPQ2t1sRbsbePKj8IpSalFbQYJe5lOPyIdiG0XHnEhWh63gR0kR7vXb+WouBlo
ehGnCDdDPC3n5UuDl8vvvtnocT1TMbTNZBuljeWAVBAZnjhVdwnvkTBKq4UI0h5QYf+SbsA58MKw
ZJfcKfJcIlpk+tg/nraeoNZb+8rdHyObN/B4BOIg+nHH5VAbhvdGYR47Sp+iPxH9vomoYrZ3TDeU
drjWLNbl9c1alnQhDfBweVYL8t6cwudoMNg1hAc34O2q+9LdT1on5ITemXWjLYP6rmQe4/eTGTBb
5sGgqnXy5gCt5JfHxJSVJHRJ+xClG+xKnV3bfiIHxCTNviRqM5PhbdpxuW54ploZCCTr+pL8xQL2
u+d49EZrp4So5fQRlQqsh044zQKzpmvYE9zZecXt5g5jOG54R0EH3dwdzo3aGKsYrjgdTzaxBW8I
VEnF+JRbinuPqwJfkSx0YtY70J1OHzOnPaft5U8lAPNynnVzLf3eDznAlK37L4pe7tTxtp8clpR/
thEC3bM4l5nIwK3I+KskiIgWo5iFGctfKBz1IT9wzotxhGzd7c+HFmAzm0vXn1RcdXUTOFy2Khx5
HrQ1mWrOVR3UuGR52LwjrMO4obOOz9Gu3qX2H8dR+jzlJSPCxiIMgN8dj1FWWEbT3lFoTEst/A4C
0irMv2pZbwNf/3+ZCwo8wowAbPermcHa+1ZPSTISux2PqULC1TciWlgDdLLv2jrJ5KqUoRgs8FXm
EDe69j+Zz6MvqDh1DYNfpfec2bVTHl8HmswPTT6+APL5ZSGypClF9VIbAFbKXV7WuvBBLCIAsQHJ
9A9tVf7ulRxqdLAFHeAvY/VuNWCDCTgI4Bq9DLRcETENlMPsTcyegJ4INyosD8YDJ2JFTRelrO1W
MkDUOrFkmABHGoIpmyKnopK28A6O2cONine924BIOkaHL4gU/6SsiNDS+Ut4jnbznZ+tQeZDr4zv
WjFNxDjt/rsd/eoGjadKZOMaMDJrqjIGr9sMO8SYRrYlTHgp9iG/fAktRixO+VzqDgUce+ufK+yA
5nV7d5Bh9Veeho8Ia886MnZ7HtwzLMeTgNumL4+Ib5bmkWWb+9fH0DXa/+3mvYEBxR4P7KDL+ctQ
1aUor2hjUpX8ytTv/zYOuazbRVKmwuADnJeJqTPt+oAOcMsQTBPuEwP89b+pjTfypaIWxEiH7oiL
/rU+m3CwykypqUH4WksEwYwFmATBAT5Ae7VLd9D6l4QTXzE7fjVWTZc7973uchhq8ff0jejzgW+N
aWfDsMN1lZZiQT7YtOq6sH1IktfKbeoQDUOnWVLS+/uy6hZCDkEHzJ+QoYBOF5PBqZl1jXdz+ASE
ExZ3ZwT9co/iyrWIUJ0W60P6lK2DIZdhdcbBMtMeVfRLB5hqupgaPoyq62leUXRZRk9SDswGNZRI
TLOWGNkSUjDiBBxDDVORqwyMK62q6kbu8OFDOyONKDE11WKlBFrC44BQ7utLbZajiFTfp0uGIF4B
jLpu0uhXeOEZWqkQOAdtsmt9LGBagiI86uAdZXcAWn0JAmABGjXOwWtVetQX18s8iZlp21NKFr26
7PJ76xhwi8Z/oL6v6sIOghyvqxLz1AicEmjflwPiXVMVfbbC0U8d45PykTonM5S7hXsD8dRNEI2/
rp85XdI6HQ+piGQkW+dAatCg5HYI8Gc2x4VYSRwV7ht8uNSxidBhkrWd0zuK9/xONFUMPfQwoiUm
aCqyFUM5U9W+xPcsVL0S+JeEqTNz3N30v0iFQL3E9F08miRYOTdF1wT3co9yvRWg9bYMzVmSoyr1
AQzEN6xLHvJFRoxjJBVZXyHEWcApRD0oBDIu9GaXBuxOJ/RXXdc7ol6n2ozdFV4q18525HhamAvD
1M9LRDDWZnrZce4cWVD0dNs6Iwd/4zzsdALS8/vBmSUyQb3ZlYj1zh25JNcanAGRmo3NAOEtG3yw
jhMg8s8W9lGHjyEWdhfI/ao+3Am5EEjKMLt1FQRb88H7CWMZ4y+xpFr+Y+mjLCMWS0QG4GZrz/sV
drtkUqqvCapt1SjzOulM3cUYLnPnIp3sWL4P0mwwTrxpa3WlrJifro73Xs7ShUHMOIn19DmJrBfz
Wntq1autgJKtjiRV2M9C5YjzTu6LTJc22xRW+xf4hSxayFcP0ao8Ko26oIg3bocCWQuKgaVMhOX5
CKnJ0r6LP0s/2/WGR+yeUszpoqo5mwbZuNCL3mmrwTCnkRSe/2XBKSMaRYa3yoXj2hLGVCsE+43T
f+U+52ZjIu8VQVVE+zJ8czWbNOZ2Nh64qmuK2Qn1jPX4EOcEqHpwU5NZy4Eq27aV55bBJIWyVFiD
bGp1XW+HwEiZa/TAmp6Tq+Wg3vGezDuKxSqac15K+MmuTFhn/HTKFBBiQA07hEejzXiIu7rDKpzL
0i1goRG066G8oxHJ0tTNO1XjYDKYcS52CXUj3Fng24gsdS1ybhJuKlZwQ+ZNjSFPd+HBuZ8hAlgb
RC8HmTAjhuaqbNAQnpvX5V0+SRs5845/7LKW4fR1X7FK0tmkmC9zwWwZCw7NBLJ9DNNKZxFdvBbl
sPkl4OIeYRdtt/ekVhpPOuyHKfGOK1VZraa0YicBjLerWs0bWxeHeNFl+k6WMsWvTgwpnxt0qvUv
GoJe+YIuQ9oqhhl2OIxxDRWX6KJMP+Fv8Lgs7ffVtJXK4EcnWMJzU0RBcUVgde6GHSKWsVWdLSkO
v+LJt0zx3HUpX/rM9NVvDC0iVwUo5mNzNAJyw4AueLpQefqo1/AxGjp0Zd7LK7vJhfWHz5IbiunW
/9rWpdyGg0Xr5iTrTeQM52G5WcXM3ZYNbDoi4U/mVA4dxQP2niMINYVJD0S7QJLk56UuRZwMkKjF
8mjJkd/noIjkf46Oigbf+PMD2iBPTOVHBK2x78HOIwRZnK7WVGHUYT4Ur7uFXcl2YXoH5zBBigRJ
uHKcRCe4GU5PT8VSVSnOUkHcJ9TZ3kxirZ6KeoEpj8aSi584GftURST0Bi1JljbgZu6tD21+MJur
8SaEzTcbQ7nFIcBCiTaZiVfAnjvwY1MCF7g99wFVTgvQCUpfgsfMYw14YKSjHv90E9TlIvRWdpSr
emg+Bhn1d8FVAVUcoBNyXF7w1Ym0qY7mzgWOofKKzbcwhjR4V5Fx4jv8jOj59VpaY7dH5+oA1cJ6
rwaVo2BZV0RRm8+U1mPb4XPkmeC0U0PEBtzEEq9nUweFObPSBfM0DqtMZA0FJxFATqwGR/zXgtfk
/86TY/2INQ1SIPXI2/tXIkU/6eR0Gza+0K+EHyXfQjO2ImGc3YXIkfb9M6d0hHuslMDk63fwYjPF
RV1I7hpLRCDc/tRmRaAk8wnRbxDkIWpbsiG1RZaMYte9Ep/dBrAqzPjEn/QoFt3CvHLGXomTNoND
cnoUG/J299vZp0LiVJhAIqQoe/HBjSOXsas79OlH2Q1E9MggUpUac38Rt7iBe9Rvyq5Rb3l1tkjs
UxLPgrSoYciNKWe9HpUcEMPwmjVGLsK4b1xiRqncTh897/WRoJpC4QuBq7OdmrGAjK6+HcIQtfw/
Ho4wUEK+fd3DkzFI6EeMnw65qLbkjgGyN+56iMTlubHVzKBWiNVU4pNHoRNAbsOmYEWs9Uo9myI/
BQueyRCOunwk2CU3/3EKz8srv7wtBR3onTYGoq5kjxjZWvHaTHbaO0AMk7LyiXQcWL79npMqTHcU
EUzMfEHFZTA9unMNrDyyCrBv8yqisrSuSD/QU08u2jtPVMXjbWiGOKd6wzZmDX5uYiWrgZ2XvOxL
yDScphxv4Wxb7+EbcvnYsNGkzMAnhE4jpbGjR4UPPrmFP04HqFbixwLe7BJqkyG5JcMLUa75zxDX
FXiEnXqC3sVn1sLfwtZxpXqNYbt6bG9CN9lCcD8zbqPzULvyWxqMjDkJ1r0+AXegrmWnq14dJpuW
8aEINudVXdGHTYeTbSay+7hCrRHI6yaovsfneKPJBfdTUz9MW4o2SsbUG9tNqJNiexgcEWjAu2bz
aK1uCAoZfjlV843jESQwBZDsBt03YBWQiawo4JIMqysuCyFWzOSVgd0qBRad3fd7qV1ULuHBpDj6
VeLGUzh6PHIbbiTZKpjuQXcLX7JZg0mdf8NMc410xUDu/TmmDSMAEQQ9ftBBx1TfNPRpdo9kiTBb
+Z8anxgmsqnWhsuFUB88p4dmbK8U75MGao/0wSoTnTSiV4lKPyiLDcH66LC6Y2CATxJZBkIVThLM
pzpbllSb1M1+G8RI/Un+MOhdXF5hrdkRkUgzMZ0wpLiylK563VsYWPcEt61xP2BiZ4XB6Mlxo1Dz
32LPQTS0nXOQYfC/dBblKoCWhiEYG4tZW+i9C9AuHotDb2AFMkbhhMug5f7H44WHPfm025ojAy3W
2kBg3BeNrn/p82pUNN650Nu81L0iZOOnIDJ46MPsgMwERsDdycyCDqei4iBv+OJbMJf0ljvjwWU1
8eCu+F4EzVpxLL68gWvlSzQ/bLVUFwobF9XKz2EtxNFp6re7UFnUnuaIX9GawLLCx3yHEAMIP/ig
DEx/7Jk/BKJQbL0Nf8vqcCj7PxQPphyTrLX5viK5e/EwYVi5cjbnJ6j7s1HdeoAJlSHfVme4N0HC
ZWcUfd8h/s1/5wFDlyiXfhfvASKfKMtmaR0p9PsyMMzWv3NrvhIulTlBJfrIo+6zvs/vfhZmqyyY
7UuTPvzIXamsw5Xnrw3GQGUtntohcsN3dAg44Giw8DVnFTRUG9ecbM+rVh2xZLAqQvvi+lat0fLa
+lf3ye+RVYR1g5l5i/vmR1a610Jk1IiuOf6vQLAVyZe3ZL+BmLz6oKRZ18FXK1XL3C5Y1+NI0eSC
SW6ISQ0JM3LroFr5aaTKZfoKetOuwt2vWmt2sMIsXyXJ0cSM+8cvZuF98mDULrUnoS1WG4agUNVM
HF9JpC2+Rm40yC24VQMYygSWL1dxoG6Kytd1XmT/PvuPlMRT3Ar4IOnG3lw/PEPpSUwYK5qT7niU
Rj7FKPuXvbE4OBPszD6J0H1RQbDTUXa9TnIWPBdW1GEE832b0MxldO3olUTm6Juamwf1i+yQfyzB
2nB/uJ1mgdGcvypugT1JGu7tXQsrTsBZmrC+14dip9aV4s9YlxGrCAUwhH9JbHt6Fy3PoMlV8963
7qEKYSuyFO69t9DZyoIEZmmLTIApXcGH50o9k1AeJvJiZpn0z9z4Dg+ZQGepHnyuzddmxuNbt98E
MPhjf5PT+bdhAxTjSABneuA49N3tYKsW2jph3gaXaP81eJY0wVCVCyapDeNtPj5uaKsqfJwVfdwn
iG10xZ1gxIqNWmAMTlUaXCbOZV39AzF3z8XF3+RZphFvDUVXW6wp7MEOg3NZZFe95D2uaZRmobMa
FYSTkIWyv5CELlBf9++0s/vNSBKJtC1ydnr7OipBWVvsDnU9UvArW+MrgXI1xkkpf9nUMG45aWWT
ck8XnpTRx7BrK9RY9bqY6Ct5KjTT0Ioyr2rWntNxSzG9kPDW++YH8bKWYqWgB6Uucvy5/Z+WZpEO
NNJAlMCI3MJAKHKJcdOdkGvNKOdMLL9GuQ8KMPyg08udzUEXuu9bBC+C53l8QFmMLuvaiQeOCLIY
UNlWoi9ailujjoDmr4X+Jq2bynwbhNVsp5BXZh0xhIYknHPLYXy1cDuluffzPzpSCB/haM8AD93Y
Jeo4+dC5SjAkjGBiKzZDn3xh2NRrOGPDz7fzXX53pwZL1g3JT1XMcSoVhHqLXPhnE1873EKmNtaD
mG5ctRwXvjVHxod179Bx4BLiaAf9Yn+eavKeAgwti7qXlEIXeVz/qMOfPJSiN29k9BsKa7gLSod2
y5BQLOS9gv2lmIAYP8Eoon+VSA+L/EL1QTwsMosRVFcBB0nOF9EEI/ecrQ/nr+LpLVYXgJdf1ZE+
or6GQUspEFL0yNbMxp8W8YGupGhZePG7Ahq5P35TvNeoliuM+VztcWbazbpR30g0S5GC5L0K9+Jk
LECfvbjfkLj8JiicDU9kZF7r2mRH1sM3MwUNlkN5IKIHBsD+ekkwQNzIB+HOQ9KlE/EFR5S5sELU
6yXOH/WFz5HKIyw7r6AEthAbEDZhSOa55SVZyUvU2e1SI5wieUu1RfXMtifFPz18fTiDAWlWP5Bt
SMxcOkJ3WvmR3B71CujQia4Beqqvf93OJfD524oYF0GntfYSXmSUgKI3Qd4FWyh6tZ3ja45YOLWZ
AraIjVyCHEmsh5t6/TwQAYGJ5oglAi0V06rnfggWUXmTfq1a9TffvAU9/ld28aL1tjuqwBX8qvAX
eirZb4wXxT+zIrPMWZKSraZYFOUv89+FbD0i8qEfT5zihWtF0hX5NDtbrYyCBNnxF2Xu8WpkBct4
6j/MQpX/yjZQ1nIbkU0BccZ3r+RFxGdIwOgAoN/y9FiONEt9Yfe29p5gbTcj4a/iv/iSldKBYrJL
aEJZxeeRzfX5fRw8Ays8y6/bA4EEkxUw85cypa+gmoc6KVcuK4qeqHLZSN0q5Sll4xUqAyhkBbKP
KDdNHrYDm6c6z2/66b12I/ubOwUdvD1iPobYRm12yP9bBL6IT4Mh67XZvxqltss0ZoL0XqmOwetP
1qHqhTp9e6cP0CT275V2+3a1FPvT1JPi4txiDkPzNJuxnsW1RGgxFOKIz5vh768AMhyUztqDTQ+f
Dcnt2PiTavIq5OSpkCrdh/0/cg5RUthEJnT6Vt4o92zfoPcohW+1NiciHhyESddgWI+fjRuPfiD/
FA9jGxhYHB7XCzEplyOb6sI5rUsE2IMhSGl3R/DDgq7GzhCjQvMXiPqtKIz3AF0FzyysmQluhBk1
wvzV1oKClYv+rBDD+vT4EItYFFQVRTvNxgTGa4qLPl9UEF9Sn8m2RMozHEjA34kt3oL5X/+bkCOf
LonNwxC8xqj7RS2TLgaWseCw6E+Pk87PRDfb8IetdzLpWZKamy2aAuVl2J0bdkCABtXcr6kMN1JD
4JMR+k8cHRzo7FsJqgQtrI9ZSiC9gZ2RqCpW0fZbZa2Wwv0hw8336z9dq+Ef7nVjJ2H8cxhoStCz
Z/FoazLyu1433IUPI+f9lXYZStTHmSKGwkNNP0p/RGDq/bpKChwmUglyVcI0JkBaq2o8KE3cojFc
2XOBHXZWJnc6tItyx7tTyqo4ftz5RdxPwiJp2kz/3Gr8S5hw6SV2JI1GZmetq3SFpM+ydKxFIMaC
yZbrE6rKfHiOmIGfUjKpM3hy8h1lSvZkliQLV8Kaa27mOU61FOMwdUbHuWWCABc2jVxGgj9XfhPv
9BV/G/9iajXKOEuoVb3/c4hoa1DURV7NQerwc1IdbvqTTQnhlWQyaBIvjqMGBR2cL1hJ3xcZX5ZE
EwXkxymdf87QBadOL1KdF0HgyQjWvvZyulc4CxEITuJ/DX3VspgqQ9VKhpBwVPz7WibO/cVe8oRa
XLYj/AZvoBz8bDOxRRtWssBsVnABc7DaCfQ4vVugrQkIU1Hn2EiHZ9SETDGD9veM8jpfzo0O9qCK
516yag4PGlsdpE04Msc/c+57sF9YXGpvQnwrpMhg32vtarNZJlAoij3FUlEbfUflUjqOA/QXqsv7
XbIHxyG1ohp6Rk9RbhNp/+5uzc6MCCb6zMt4ZW1yfzx6EFX4mEh3zM7JXj2nB+AyKb7/pBw+wvlH
4F0IgDevulVOr0wTRr0tagc7y5pFreaBB4IqwgSzCIjD2Jm7d3XqiLWLy9ZeXordo39zsYqNjpJ8
J80zKW77b2lY2TQrwBdzedN5B7WxV7B+lJd8E4EZI5vXKrjqkMgaGjQJ2doPYAvve1JO73RWP3sH
skpbWxPB8/OAXq1LlMrB+HcbsXR29OdsBzry+oOFrnIg4MXihAu/bKFnWh32MyKacIFrGeh1z/mX
2YUz9iALIgbIPC7AofRCYMyg9isl1QDSzHfb0ykFUsesSLmRt1Zj/d7paX8+y4evjCvnjl4TaZVA
bXd/SR1GPxr62ubKK0a+v2ZgapL7yTuR7P7ASLczM5UGwrtHfdy6qo2MaHZUDe8TzOnG6BeQULvF
6iP2OcxeZvg0vr9ST+uwEknbBhKodTTs0G1SUl4/zTVEnDGcH33VdzSq2ZTUAccWyeBwApMS+GbQ
kLKQFixYJTJ8NutlLrFvUs5MCTeil06QMTT2qJsTxQqER4zUNtg/PypTXN+qU0gd5nToUHTconiT
4llKJ7cVGwi6HUf6vGKBOPcfCv9L/WAgwU6Rxh8I9c9Z4/7VKyNYmkulF2SpZnrnIXGdT2PkuvVQ
IJ6BhJ46pgYmxVp4AYdHAF1MDNIuOLLqRDuyrnjTO03snWJZorwU6Xpo3RHzhKNKwIeCQsrbWYkh
PFcSldEMLqUQ1RdEW9a7v8ayHvO/pXxoWdfiCloKI7Vajl9jtudQY0jgbKk1YjtL9GseWKJ8EhT+
KPLXzfAnyBkVGZUSFPdnQT63SXdCnhdXJ1NUeuQvXy3+PRkEtM3qvqQohCuAWTxBOUJvIhRn/glk
c53eD8cilmqEaLDZqCLEAlmH1lkf+Mp/yfiHMrXVSqM40oTvXV8OICgSrRlalUXEEjMHU8JZGaqB
TnSdoYaB4Nqc787C3B9JApz3tPlt1Qjxa0D6NG2JhUbEapDnsyHoDNEezwI0mXTzqH1Dx+AwDZaY
wiGIGIPkxVYXIS+MVvRiL9sv8r2y8ymfEJuGRS2yC1HxxSWolNalGtLt+GaUfR7wzZ591tpAYbqA
omEcvYwIpST1S3DCcSUwssLgC/BjkRAmZbO4mdU55ZHpoi8FlT2aVUuj9dh6jVn6UhW02rCWswiX
HduMyLJCMA5hjK4AwNGBgObzBwWIaovD2/yJVdAXCD+C+8OAjT4+xu2P6YBTp5s7h5yNnwcMr9T2
8NWM5HrS03VstQG/yxMvw6vy1NknPbisV8ZvTNKTl6H+AS5SEOgAk426ielfpXcQ/aVsLkSMwne7
pbILj0g+Nv9mTDfXv88CkfW4BDwKTxBZ40ZVgvwVUPhmUqDboYJZyoCnf/GNvQT0iBHFZfYSG6La
Mj4C8FUFBDjLdslqCgttTvGkOn9gk9uLSaFSVOFIjR/aJYPm4Y5/U4+79iJVp7yOKDdW2YuLBqoE
Urn11WYQW7TBGaP7b5aL+pxEtG8UmR0VwPtWLBlJvvvpgqVh0EDmB/3t4AXfmVuWRRuS4seNFY3m
fyfE2K4hRJlOFnldjFIO5w4uQ9kxC3oZjDSsfTUKkzGiN3wkQhMN/MOfVBRECryix78+7CC3tTjN
ZiIWGC/kl0FjYvaY+03SOynPEtIjcW13y+iOdkrvQFTcKK5ad5ueTvtkI3Wv1/lXuZIyTx8TwK9V
4KCZOpkBUslrswGAaehmiNqYSJil09TiFYVi5zCOl4RMnDvETO4ZBSpdNJPBThMvhfLZwnyfWWB1
Z+wXSwf3ELtSxhnPw3HNHcVEYYOY9dCgNZlqdwuOtncxi7yCOdEUimbaWFQFulTlzPsJuVZ6Fwus
979ZPQKP/dXBrnevwcoU2i9I44rg71iCvAsITKYwfD1+lsncalBW8+Z9myhlHwhKM8VubEUniajz
NDirRjxrl+GL1b9zDlueUu+ITjMW5Q39f44ZFF8+oNBk/8i/iHBBRMcnibUmLbrfgjAuhoy4cad6
8+zq5AFAZQ7HTJi+9NrfCLJsmi0nJF5v7RkyoANVgMgWDpQWmEsS1Lk5poNuIX+aZ/2KdVnUGUzT
WvdwUbFooQblYri/KCVAshjQn7dhy17PzMv5nPrh8102jedIUmJax/R2xETPdFlAT8mB0cIy1kDG
TWCvLOHdUn0oz3wdz38D/u9YiagrGGzw9hqT4L0XPyzKlVmFF6F/+TBpzpUDlenNPR4GEP2TQC08
WD1Pm5jf9Q4kWYEQCIDk+sFN1P1J/rrs6yyil5WXYXWEXPRlvtdvk7PZ+wF+CHsU14ieZJuuTh5U
ifZkpDACqn/xd55J+7hIZuA4akijF63uyGKODmWJgM6hjFRlZpFaH81mwXaZYlvEr8EqqDAAxBge
x4ABMnrk8oQ1ezy58P7hOVailESQGs9roNOJmCm34UlAy61petOOqrqiAddLCxXtZc6F6m2akQ4r
oERfLZLAaLtZwAd4VwiIpKgiERrmoo4DAyRlghuTmqSlWcY5h72nZ9OmAuD+V8QncKDrWacqM7rC
20ZYfsHtxvEz4kyGAKJnoLhWo37HJlo2zi+Oa6G2bQrdZ/jOhFz1IsuhI2KrmcuYEGpH9hT8hxps
uijEZz5y6sQVh9ElX1Bzb/bbbG+kdW/J05pgQM746RviDyj8w21d0I82N/MA/dxVY4eniZ4Wr3Di
kODv/EsOj0hTbaUtVQbaJltdYHNRsq2WKTBDAExCCFyJG/2brszg7CLG9+y2++VgcG76YBTmwZY0
X+Llldiv2YYciScjDp//DYcpIRjMu7C6gM2zW/VLt2Gu5bUifiSZmB79O1FmuYXLXqb9BsxGlqac
R8W3if3n278W/hzi5VEDwtKgkiPdc2vrGOGEnj1efgcI0G4Bomk3AlmUsSspFHfRFARodgjr99Iy
eIvIX9xt5XFyEqTtRW/S0dbY2WTRA1DLUlYHIL0/r23l6SeV9aTceIDJgNDHQsac6jA+pBB4mr9y
xe8bR7pYzT+cwt83FtfJyu5tZUOvyd+y1NexbLLjliYzU6+pUuqCtQLHZ1yghAnneatKiZkYkyy7
t5XCcQAJN+BMcMyv9D7r8I+Xkq1hWiR59huuJZHevY0gDuvfwNwxn+xLx2P8FgZ2JAr8JQx1MnAZ
8Zlr7pTeyCWaDAuqtuaxzv3lvpFuwLL4otUG6uW0Aas3HbXbiPoAAD938VQULrmokoN3nr4znIHZ
lPKGg7oCm2XW09loRdy6c7E7/0VHryiUAWfRH5Ttsw7SRqzkj6/CLtNUwCGoaNVhn12bnbaKcznW
pjTSksKEG2XgO66s3DnlklZcNuo7K5AK99mcIbFnPxORiCIXp1XJOm8ec2fs/C+kBNmVRwGc5JYk
ZOV4SpnY+ni9j2zA4C/LnvPPsbouMnU6FFCb77+mRFnYlfeMO7Z0uKeR14GQuZaSjZM9Z3u3rnYI
ecQftfnWag4qxUEbGsQ+E/WpVe4Me8iaFZlmoTZW7qLRKYtxTjxx8l6vSdRYuUkrGNw4iBugV9gH
uwoEn06H6/W0iAzSKPSiRrw8S+OuEo8IfhlBnTlYpC8++2xI1MfnM0m1RnErkKJkNeTYpuQeL97X
KCpK2U3OCnp1N0i/zyNA2nbWpmadjVjK8//lXmglboU2EQJjiTR7X7AedO+0tlztdhlKsPhWIoKd
aMy2cp2BVQjkI+aOdzilukwjD1SiDmv0au52iCuBd9XhKxgRPrzh1hiRnTCon6v86WXsUuiWQE5S
Bj2s4Efq7tAV1Mx+djEygKiceVE92EyjBuI0ghv12zRcSMM+m5oePNhtHpAIzESdVny/dkoFHwAt
ayqJ29h1xDYQ0uq4lYSYAtKZWLEaU8ZXvhMMkmHZRCwyvULlWyNMpFLest1j1yak4WMy2vRXqliy
oGM1iiVov9TasdBZqtMQ2DhwRGtXCpJUzalOzcFzxw+unRVRXKDPJocYefrngOPfT/L85kFpbdXU
Veo1Z0Ut9LPNjxstxKGaHzq+PeY8ys3+M1llf11oprZiAWLj7MP2WLRrx1InflOJaEw4MpAVswqG
rlMV7e+nlLzKL9BGAGh/YuLfzrAr9O052MJNlpDTz3LuVNXcPL6idm60EaS8o6rracKaekKcOtCE
pdFAmTyQMUeycMiQEdW9VdOjrOQbbpsz/oMlxM7N6CvgOPFrbEgaJuZtg8TaZiBmik5mAvoexSDY
eFWfyPJ+YtDCcleYADyJO4kt+HsWzffqkI1xMT3WXem1KK9nAP2z2wSOqRv3UWx7js68s2hA+K/A
ed+o1e5cbjIaf5YYHnsrVefYwq3OAYFvyn06C4FnXAySRNK1g2IJZCauZGvntFVonMnoYW8+mnAh
OT1QRGeCv8mHpvg9Uj9TF8T/i34FwWNQaZRkxV1r2Cjz5uCRyQRsPJEQAtLZHhcEi4tpjoGxe+OP
tWt1syQ8YYjA/2EeXpmuO6NdLyo/MXHfupxyouYE6TIoADggpZX9dyS1ryRjwkBUI9jqN0xyTk38
unrG9tt1Wc5aF9NVQCPyVA7DQZYkU1XQ01disgLEJFhEso9+96Gnss+8AigHMfQO7IMONwziRhG5
SXpDjrojtTUiEfNasucJaxuwbUxuKRqYM5eDois85VvoqJGOUBgoLz3Keh2LZUJ1wpn7FyYy4U8W
bUFOKH7pFLfsu8oW58X+zdpNuTKfM7FfSNh1wqhAPFLLb+BXe3Z1rudK7sDkSefkKbsinBpNuEaT
NN23uiGclk9PJcB7Gtl3vkWXIgcZfyPPx27VOOARI7r5Ii0VXteR+VVqIwlK8OQUvQ9NnvhQpsYV
o2cKroeA+2tGIs+LVmkg93Ci9b61zVihcGLOiC+kdmdQtU3g9rZy289GFjjEO01wMubUxmPbFlbq
iDct/s5gZ/Il+j/FVFWUcTAPn8p0hEAoa1v8S+wo4NU7yswRdd1XrFcdznNbuPezZ31uwa8X3TTJ
7S0ZAk1uSF6hBwvlFCt3dSvHbzIGG0ZX0f9yin+ZWboCfi3NaicaSZ7H3p7CCK9nDjYLTHvSMgFz
ir0DBQuVgRu+3U58Z83sDmj0gRBP2lYy4150Hw9GV80R/W2QiNzrDn4CvZWwYlDnQR+DSEiNvAY/
uulo0oNWvi3Cl8VRcgRGK0yDwO2dVODmNcuwpDJ9z7/TVRdwJ8Urn62KbCqYPxhPBD1HGG6XfZ8K
NBSNHLvGpF2q7M/4uwF6F8e+9CaVVsjdeERtjC942MKwDejA81uiN46MnYNQBl31navBOLPfPHvn
50ZAskOTH7UpxJECO51WG+M0wFDIIQercoXgCCR5G21otxKv6aHv9rR76A/DzALUuVIHywp7E7q7
Rlwkw0t7zA9TMNrLSrB+bweoN6d1qFrO3Ftu8jaBKIyuhn9wly7BYWHUqMlIXEKq/9vDab2rnSUR
U+2iCnHsORbeFQOs6JBLRdBca/hmuyd6N6wu9HAiOUX1cD3w5Su+JIPye+eE8RQvouIbJjBE6qa2
q/U+Z0cnHLrIKiTU/oEX1cctLHWPFc0jbQ2kIlmQBoMI0Orr5WEdsXr0xyDMVzpnGZl/n8DVEslX
Rliin6ry+aEZV7wHAWIxkIxwpwCFyrP8Yksn/6Qah0KTAFZZC2/gLC5yDciItdeCYeBxomXVwfkV
4j6+Wp+OwUxLnA7UjMv1eGsTKlGPfQ1W8leZxMT9LU3VxSjvkTCqX5oahl9YY+yLzKeaIY4dRUGy
NqzTfaGDN4AMjgpU29ibYm4gONwFZ7XoeZQ0r2EGgc1cL7zx6NznOai45QT/k4uBIA/0ezdjgDAA
S1opnfVNlQgfEVlPCf9jIVjwk/KXHgkyAYZ0rr+wvRPboo2f0TrhFXB7HqzKZWqHfwQy+04amnsp
CYPMOUH83pDEEweQ8kwKcqGvte7nxEldVfmCkG+xVYrJMYHd7DTd2q2fARI0f1c1zSjkm4jFzfzS
DeXby9SEAl+/Q8htyN2VBdCgemekbfCcyXkQ73ohHr+SJjMkZH1CCztjG/0h1bvHpagZ3WYNzA7V
W6/J+4l/fPOy4fuxZ+qpNJ02YMugd+TlL84BpzD8f6Uw+Us27uHv6fImzf4raJHuWMlrvuJ/LJ3N
RVXjN9994g5rB2auK5nT2Xjl8MtqEjPSkkhLWELAyEXJ9FyKRoWLmNRQReG5dJiS/BrLqp1XZI01
58hVNDycJe0srbdDCeMOXj6I+i29U2KNjKasvWvUpKxwqbxfgcFq2n4a6g69Dyeg90Qen+dgDru6
1CRN3Iuf9bNR8q1diM81M3Q8zQ+vRd5o/kJ+BD1Bngc5jK/RaFShi6FL0pvi9UMaQqvb7kMhplql
o6ElpCjDEHRQJ7wpZgFF/5ZpSaTACkDEGdpFYYxO69i0ewO0m7xy/+RVNR4cScWMCqJcWOMeDYXe
FXOWtz3qXgXWdIGqf6uPFW/9rHVLPsH9S+AAspM8OJOjyoXqSDygBn+aH/EPSISatyOZHxBFcR6k
fFTZd++/uLRQSSbmKMOGujzL0rhHg4C02/JZjiWFgYpTLE/1FAfHLVPs91P4QHG4/VHBut+qnrUS
vb9gTZUooPwM2P0RbsIFGkbywngGpfzJ1zpB7fG/iBozY9ooAfnkqjpPwy6LOv7jWqRb78kE0+IL
KMaxqAykLz36orBDR9/1/wKyDS6AumFpt1galXIUg1U+PUf6kKqll/c5b9zlXzvBWD+bwwqzkVGb
5thsgfZj9Kans13I0B2akYVw4GJSvwuqEliWl1ewY1m288DbnTiKqjDKcJdHb31HZXumhWAttTTi
pIzLx6/DkVkJ84kv8QwO2Lz71r/BzMBrGuxsPZmUCs/8uQxqIHDV0jfoyNt14as5Mt+8QJqzofNC
Jn+rvsgk1nLJ65tjTrLCDPYBs/Czer0cCRss0tAsvXJL+yXCF8M+XvV/6H0j2t69rgjXBQZ1KWPU
4fxhdUf3wkr7Q6GHoBmcRiWtRowly4m04LmD5U/qlBGJ7iF6BSH38kOFv0pIaqPbz2NilBvbnzp2
s1QFwG6MV/7fYT/JG+YPCy4ci9TYRkVDL2VZbjgmkcHxnvg+Wx5F6VIkJT4AXmK3LIieOBfdC8dK
u5a5n36Di28ODJ2i43FpTIQl7zihD6/x27Fu67u85ErMjCr6Z745YA1lpn4Wd4l84I51CmtNpEZl
IMth1/SR9crRcZGCngZdcLorV2pYPq7wznq7MpCQ3cQ5mMp/JnRrDxPGXqZCyzs2HljV8CvmW+TR
k6lMGD6BIxZCO4Kfoi4AdtA3ooF7hTvfP7+2/KRbprGTHA+11RBogTo6CKqjeSvC+UMiHfcjyKI4
/xtnaD+XAxC5wED25CL5GWDsy/L8Nou+8VsUqdTdcKFS7xgj8xl1V9yMksrA2K35yaG37hL3CB8s
U4Y1yAYOvNoxk4YPQVHMSEW3bMvdM2LB3vq26iXJkYuGmw/xEgWK0YpLsRjyRmjI9TVw70CXBq9d
D3USeHjJysqd/81HLiTUmSiiFGjp334SRCjJDW//dSot4h0e1o9C3ockJ7sFyEWkn/JkMuToCaV1
2F1ItDxlX/C9t3llWIXJ6PNT6jm7RQ/n6O6+yWLzKGjXaJ+s80MHgMceAOLCrnhaA4OA1t0yvFFG
Qc1IDkbPwvn6l1LRawvvk5Zszxz+lk6VN8sMhlTCE6r2yHxe8JRRk/2CP9OAb+LC3wXd1+M/t/FT
0H84P1iG0u8C+YR7u01QVtGoYPSxapWXPCNHAMUNKM6vs/F4RgUnOP+PEmlaWfGmyBbPwZFFH+Dc
kMNt36TgaDBKiG/ckoPYtqUGLeffvPfRxF7Wrm5J93H2ffJHkeZwK8Bnx/04Ce/HtOTw1hwnvAmt
wBAC9PA0icsBA5lUAlyaFgPDtSs5IYeNo+0UjCc5CJ5X9CIxmtaNOY3NLEEA97NVdt+qxRPO6kBg
0/geje8+QSC/zJHj1n/Q/nnkd8U/jtASbHtRTRlzOuN7M9Mcs0aNJpYHmFSPlzbnYNDfNyK1SJ/p
fGmE+GbgBh7TctHlxOu96TMqnZffHnfedW0oWUK6vu4QHOoXjqWvHEGoaoNlI8ZxuxB/sKG+6UCR
I77YmY9K9qCs/VQ9I89pS7ZrcOGKa9MG2UjC/0tO/q6be5tdfu1XuDgxFs5O58I7vvL03Tq2Exmi
DPIJj7jinlj8BHMWjmtDhQ94GoVkJmWBGK2xYWI2l58wl+5Rds+MhCdXNBctdER1v/PdA/m9sj2j
vP/5SEKTr3FbSoAURXf/1xb4S4MiwCjLxAmdHmpB20z+qLPtZTEKcNtSNP+ogxbu1z/rU9JmYOTR
Ki02HpjjmFyLHDzg/6lrTYofZNu1cQclaXTDEDppHitng3rGA63pAnGLrxbqxdVJU1KVAUvANe//
kJvhVVrCRznpp07n5lafrtLTg7ACCm628t3I68i8NxpcKr9ZmYVf2EtCkjfDuOhN5PXF/Wnb+I6N
TfTKvLef25bi9y+VuVA/CfX+VS3OGWFFeLX6lhh3AIT7s085WnGEfs52lWl5++4py959cNaizUiB
xtNvsOWh9g+bIQznb+g4sXpAehVLCFoCckapgbLTRC5tFDZuZKc+0/fSRrijP+Z4GMQ10QZfpEOK
pra49RGQnMzqtRXqLB/N6Ftz39B92g1Eqf8IWRv0FS+bpMcRnHtISuyukNRAGlb/f3Fa6YonKaDI
o4gxMo+Q1gfZ/Yn4VVwh6VzkoeX/Mh75WZ/sZWsIT/Sj7PYRBYyQ9XT8ZtKMXPhbilVsqUY8G65M
oJ7Ou0sa8YY6oXWo8q7lisiG1GPAQc4mBqa8mvVs2TwN6oQbXqtHZf0sTkpfkNV9WKp/UtOJRNTU
03Lj0o+2GwuZD7Cn+zbHoNMSBtjmPqpLkGTKaCyExaI7x2opXdLels1FMkthgUTwusnPaSA1meBh
UoREBmsUq7Jj4W5nqzAvgRA0sO7t0xsg8ZGGeIgYtIsTFG2HNFfsBcb+F63G7i08pD44AobSkp8Q
i7G54y+MnHHnq7Z+bD0RU3Ob92fRxMAdU+jmSyZJwJniZfEnEAW7rkxbgZEzZeqtRSmGasjwySO1
t3v0whuFVUxgnsfESZCiCpDk3cu5Dn0uk7aiII02rjqrKUJl43SAbfrBznVSwUcC25C+kEng3Wvn
CwZmPF1/sN48fej3BxfcRzMe1Fsz/IwnEANPRWYaKXaHKX69Wp83kdbn53kjl3I3Rfw/Nd7g63EL
baFqfxyMx2VbN3LxARsMrzkAnWfxEJcwQPhCbsXQ4L0ugUxBNQERVxNZu6MWJrVogs334daO89ng
1UUXNVTDK9AzNLm35HeJ5sPgUmZFjhEOIUEInS55PMYgHhgcCrww7gxS/1zi+ll91GTXE3UsEZfe
CFeNr56MuvzV9oqtDBVRPMWmm3dxu8J+LPXtXVpbfNgLBUXwmul9s4dr+6p2ujyS4iEgg2Sw6ySb
snj7hcnCRTa9AODeeQzCASEOzIjSMhtpaJVFyhsISRzIULH4mQQG17kmI5pNoj9RMhHhknXk5HSJ
RyGfJcd+1FfivmbE2Bc39grwEXTIBQgaSObFqTMfKoKTzok9vKTWJ2aQYObAbehFJ65dW5iOnZK/
Tw2GzbwjkeGN24nDW30Iohx8hSH3FXbXqWYiIAVcXBboir/aEorNmCoXg2qY+IfCzXYBp462KiZt
3XdOD33fhf6aqX0DMO53AlPj7ws3bx3QVFd5jANj2zx5D5L4kSCJUREj4CfzlKZdDq1qLeoArp0m
zAiz45BZMtJJyEfDITpP4GPwifirERFsPbnPVuX/RQCCQ+soyy3tIZawUrdez8kuBr9VoYe97PWo
bOritNGyA2e2h09cV2SLGaLegRRwOjby5G1GtwmIoAPosEfBkgBXHF7yymFC0+mjbropbOJc/iTy
dxRLWpn/7Tu01s2rN3vp4htrONPFRev7VNO0p2bfzcNfcTiSDOeoh1i+/eK9SZJ3246nAgD4UP7U
QzLz9AKZyiBWCjg4mHLJ59XSt0kJqfZ4GLUVAX/zGv8ybfY4CgoR9/pJKmtJhiQN7KKYz+KwEmYq
dgs8iRmwEtU204emerpo5BMH5g9VZRXZN8wrAjAj98rGc5ktd6In2nTcQdiAakRvn5lJ76NpALHc
8Wi+VER2s9uUg/JQm0mMzIX3silzA7uwmRSJI9Y6FWI8sMgNmj87Gmsgufizt98XvLv+urWV3kN3
N6peARxuSmBZsYD10aRHV1wbjdVtbkX680RWINfFm5mjSu/+HzCTKRrBl38gDN4bPiEFgmScmO0F
2gPVAVk/Rlyrb6nR7JOkYbIY36bUOocJ6FIuLnmL3BsZmx+ranTzN4RTysUI7nqskXMS8Wjd41Sp
e+3zE6UwzHHT2sm4PY7VDShdgmKSZJYgOvnusOeUh4uLzwPw2MxPC1HWr6MfglEZXQgvngJ6w3bZ
JDMLxtzdZXjhLJjdcPaRpovMdN08CVK8SA5C3GZgMGcJOX8C8n27OVYlmWUn/T9fqb76t1rrB8pC
kZuElw97IlLHeqjKpVxiFDam7Ab9mi+HU8yHTNhypbivnYZRExyKR8UZ7SG7cFU3LKjpI9LD69Qo
B5kMP6nmYt5brNpBtub6A3xDT2vBunGsB1RTwZ8nxbFpHUETOjwI0hVGHfUBxoHBObth7czRX/sL
hUZstgqvnVNIr++KCjVh0W82zvQSdqfqtALETOpCGcXITq0t7hL2e5HLoUCU06nI2c/c+y+dhNF9
C4B7Xtzu2kON+jlKeGXUOUYOYVZGfnfI9RNjfiunb6nwZYPH3rIyPe+/iPJnimSbKoBUtNAbHGyU
XRQqplnJJajMO7pPgR7hvSPqnYPgAGGcwEKc08cvU7TEmehc0EF9m2rwzzcEIazKlLLUtiAHnJRt
xT5XJTB+aMiXu66z3mrTsKjxjuZ2eqzroQOEFcriK+KIxFKLqh6M+nGn83Y3R+KXNDaFLYF3g280
lQZF8M+KhAUsMARh3lNnNZMNUH9yApmvLbU29ltY7ZovvskK5Jsksvul6XRpejiPpYBIJl4VgJDR
xXzbI9oSLcsKHLlW1HZaw28acCcjuxXOgWZhIfPKPgjGHJNlm2Ody7mcCMk80moaXNJmL+PDSMGx
SQRceKFVhzNdaUoEvMq33Mkm5J4WFeBIudm6SYelfa2a8U1NIjilc6J3Y5gwkR95kYGXl9KxM3ig
mUoeE1eJedyJYfPcLCH1/Bj2M7R70Bkfw3MB3J8MpaPZm3ERb09pSlXkhi7a9lGBV8LvrHrgn5QW
qAbgDqS+keOMonwMYNMIX6SsE20gHLLALzlL4exwkirS3v4dM89F/ye2uTr3yQv3PrfMjWGn4Oy9
0GFO+iOuII/k9ZbLJLpIsA4N2alnIIsrEKe7KBj9u9sCMN1QcNc4nyhnB2u04wTSTzHUaClT7+/7
k3U6CBFHHkfwXoU2iwqLUtXsojYW5GJiyIyrBgAL6MpRtYQzq7VKwS+Wpdpv34L/HELJcnh+G6so
yueeZrH6izbXzSUxtWFc8Jy9mvUcFeaaQf2yFXcitM1hYt24+GCY/a6hkTro1frRX7h+HwVZKVUY
9pYjDP51bNtOs3YKLWPPcADLq1ZyoZggyX7bhn0qgteBTOfx30pAT7mLRkaFeUfRxtabE0FMFE74
ZATzsV5y/vhG+sN2173KIaPkNx12gC/rOf5Vhvwj/05sMtoyoOc1CNIbQjr4pV1pfZGSRcKBegm+
CwPxw5rT5jRc1F21RgfSNrC4hTNPBaD50yH1ifNdyNrOUyPeZXQiZ/VD9axfjocBx3sl1SD7tpqt
mjJSSKrfsCLyLcnl8054/YJY+uwe3jDmcvFgp/8fAPEXi35kjcleXiK2bXZ10Vs5X1ySFW+asavG
WDFzDZ0rNGT6UiqI86C8Dt5/R4nQYdWcYQ7udgRKJuKfHKI/hw88b9vK2oHmy7tPuQHoQltvvDAF
pKUuTnehziFFpUtDP4bsN0GDg0ULzQAtMnq8n2rautp7qS70024bO2Em9EA9l+10hjLyTLh5WUfG
cDEI5NpQptpQRsjjjaReepoSpT3dmMDf11qhmfG8VCQbFs8WJFaE1IXXC6J8/+ItNyaTSmeFYCuH
Pf6e+MeusYzCded45o/MsldbLGP+f9Js9wdV98kwXdirEQv6x4Oh6+v1Oo3jWuMXZWoQkQXh+FgA
nHR6bwszdwwNCbcK8krY5apWDKhs/uW7lJeT3ljsBmhCxt67MBO9YjGPhxpX7sHCvBbEtHgU8DH8
oKfN19Ed3tjy8qPTii01pShajO5K5b2GUHF+ddOdooh6vnxaLigciuY98dxX3Oj8e+DNOJYMQw9M
vvwqR1VEkErEjd765JCWgZuc3LGB73yNorgLG2tyD6ieJkLmHucA1E4AE0PM/Kr4ykbUcZXKBEqO
mRkxwq/gjOyO1NzUMBWoJaEqQnWlJbUyFd4Tsi3nCaZplU/cMFGYGChvu5NfG4UG9L/tM7HzMwgu
Jt73jL4Z9OXEFXOylfmewnfW2Cd/AmDA/Amqvau2VrkdxFosNJlC9gczXSSKCU7HmPZAFepp8irs
tDyENF7dqQvMiKiT4BmDJj8Lg4ZO0bJUvOY6+E9Qfyc50nkZ1MQEW7LjVvqa7xEVj4YYj7bQoWHE
8u11o1Rlx15dSbJ4PD/xxBMzwJcMRiLSvdRNk5Ra79xMwkNQlSak1ycmOryaka1SAi+hSYc9iRsK
PCLII4G52buhe6cC/18ERb6/8XaZJcwWYq0WvbYUz9BeQiHN/sT9+h9oh5RAgzXIZdoHIu0lrnx7
e78uU3Jxs+b7ObJEoN3A3RX1thf6NqRpQpeMay9RHPAAgFr3x6G4Gse9F252sXucnRrkDJNHYetq
UjGkYDQAewC06uCKsYxH5t3EM7XiiAG2guFAJldjCJJLMnLj5ids635zt0WEnkgHZsh2TuAXSAiw
oaNupE+Bezy8ZX/2yWdaX4SBjz06KRo6OqpGqJT3OYG8bNk5c7PWLmN9AAie/mpYn7i7VLCjFOfZ
KhL+F8IhLPuz21F88mZx7mjqqiKk7emtrgKbjB6HLN1+quYBbf+AgSWkvq8WzKByPn8k6708mSrj
bNF5MYiQRQHriKIal6IbvEYInLCkzTQfnXnWIygh3S2sHLBm1fxK2yDzIwX11V6ls0Z8mjL39TkY
usu9udTZ46mjIedyfXXsWOAOqZKuMLcuPukDwcFpVzPJjnaW12n6RXZfl3/DYRGZoZ7VXOFcHho7
lfMEkbt+QMKB/7oCFY+W3oNzXU8njLfxFWl2q+cFABPxWGzka1EWTF6XQ508F40XSwvksY6bVHLw
iSgzJP09fiMFaU9PGpQsnKcHuWqqgVFkb71C3+7tp8LVVYtJiwUHqeIDQDVNEOy4i3LObYAINsBS
BC05Z1vgftzNHal6RSMVZ7tqlGI4E/O90063LUfw+uaImtDyaKrLC3c4TJ2M91wNe3QCdf15YQ52
PO27IEF4ZcPgwXaznzunXq36KvUgixxwgFfWxfiT47Ldj9iIMS1rvwhtZ8DbHUwfDOmrjaHmHPJL
QjVfWBRG64LBlnu38x450cetJORo5wkSzsyfGbURkoO6Fmws2tqqyfGM9QIB4JUn6aYY7lwrhXqu
BAXfwv91VxWI0Qor6e0j6u0HlxIgTYYh/6xQjaNzlj9aBnh7lQ4t2N2UkosnA7LPc5yiYk1st9hW
AZW2o15hsGZIPmWe0Q3PbcsD/4Mh51lJsHESXt5OtuVUcP96qsP8xseyY6tAnRXk99cn4a/SNpys
06DH/iVEnfnZithI84kHGucw6ZHO/wcqI2QWMLg6tZq8R9Ec/6Ft0e/ot7F2IZJCPgZyMuo1jZFZ
kOU/APPDPhzcbQaNKlx34jAMRKdddpRok2D6nr5zZ0fEvgPVfIX2u7CSIgSGFwtESsz/o4l8CX5m
XINbj/f0rkUYuAD0K8cwF1wPKSriiIW0hiHnimOnslNUyAtwkQT6MvMuBM7f5riQdA9rtlrEo5/M
um10LK0+WbrmAnquTQgRQQXwsyUfAYfhzyNLCacX+kyBI1j6iiEf3pGxFvONOlMLuH2uqFq2zIRI
NhzKD+gX6nlO3C8gYjbYFN14nowdw0c1Cl4mz6Sf9Pa7Kp9AK0OHA2MXWXaNHQR3qSwlhe8V4rp/
47Gdq8Gtv3HFfU9VTe7O4ipBFZ5wksL/fhTtTIMYEbzM8G3sVNrrBl0SKb4uQq+63jrWopIjPQNl
w5NEHtFYPGoB6ezErEEW6vrqhsU6xgBDtcAwJVfrbYeOnQQT/GbYmdg9Nig7s2i6LVpeIGvroFNn
4r8N6j87/AJRr1aP9JHxCh06aO/ORDobuTCOJRlqACcHdYT1CfeKRlIF1xxuyoyCzGl9Qr9zNn9M
9M29S7flODh6vdv0zlyzY3gfOcQND84u89s+Drg0vnP8rL2zgfp555KJgsa/qFE56CSraS3DQ58Z
bz0pWwIwQST2ZF/UYBlYusmwq2LkI7OjfNMt8ap+oz0RPDlZGXl9eaPhfVLqqxVZV7CFvWIHv8V/
atfTizBoEBCQdi1YuMlp3tToESUApQOqnONI0NcAiCk8UL6JTQkcGGNpsQVY7ZCA49f37eIgyxoV
b8KqIX/qhK+8yWnhsvcLP63Pl1uScJcHcVI97EoMy/thE3Y8mSgQ9RAZh/ZYLcOAOgEAfV22WOi1
MiaBa/yDbIWotOu/+SJcuqBlxj1UAdzmAMRavM6jYWkAS1ox0iO5OQQCPa/q0l+KEGvRxfDis/Cc
WXcSKe2KP25x+JOeGSiD9ihb+ICF/1c5YEMZgtfbU/fgpRY0/6S2qM807TSXDfq3tSs32o5mWBDU
mxRZgwWlqoJ2wG3jkbo2Y9i/e50YKsQTH/Cus6k/2e5zld3LQDqJ3vGCtBjB2HmDBFe4eltxIvZA
6o0VMYnQh8HR6/25fOwF1heFTMTqaxFkooGtY3JoJv6G9DbQF62OIfu4zhn5yoG18evGS68z71Jf
zoU+Vfw2XEfMp3STUpmRsNLXAgAwJicjEpsV19kTZVCElBgOjLXohdEorBRBrxbJbrQbor0hyEQY
eYh38uj+R4U4OIWoDjfAG0D5EHMmcFwB++jBK7AQLtUoz9I5CVinUAJotrMT6sfRw8d7ggdHxeHf
dVDYKa7HCCYGMBnkVA414BAGwhAYWDNRbmCcYRwgi3dVE1Eb+zL47qEtJDu83+tmECBgL3qYCPWw
tzSboJwPwb1J6UPm63RMCf/JmcysENy3Q6gFek803mdHPqNuBaYJhpDbE2wWlMQYzyIqw6ykt8Au
RsfYyMxS0a/t3kQpI6dE2C/+uIICi5BnlaEBFPdfJesCA104AIo+CPfuDjfhVkRwxkEEnfuElwTT
696MGmmBNoFWMkE1AijIRdxWvKzVTV2NVZMSv9gMnyvgoMuCcViD5cWH+bMekoe9jiCtYirrg8Zi
XAG2F0Ib2t0D7/sLNNOuxFtOMl7KliuMdFCuZ+ZVHAFtcoPUjh84NUe8vGnKdzcmZsCWGxS+zYkL
UUunU0WbX+fomXEW8vX9ILps+vVpwZ02eBCjtykXdn0ZVCB8mIuyLOKI5HN9Thk+V12bWgYONkJ3
GFBPg5OxbkYMjqHsXuB1xFFSJYW/IOVp+uLrWK3mMEcBfAklM5xp1KWZaJdOu9o5yk5phkrILeEZ
ZTP9Ea/KHMB+8+dBNOx9fx6uGV6klHul0ntvxKeF66lif0TkH5Sp9jqbqU4TDOqfw1BknMQ0w6iY
eGagw26ROxw4bz6JNRpjDuNMl/uL2k/cdz+/e0XOmNFe9eRUc0mcFbhD6mHvnD0KJMUTPgKhQ/v6
UTeU1KBHwoU5rLMEzArqU6xXx439O3hMID6QLl4ercBQnAXanbsJPB0AiNccHPvP9OmKoihGZVv3
4IqMzKTmo9GZn514WCrInLLMj19YcovvqLb/MzbiJX22TC7uZClEsTc7BsQ9SrLlZqvqPX4olcgv
vOiabDiBK6gXPvKeMlD+jQxq0nden0P393sZEb4Dc1jaMuGcN21nWBkbuO+xr7rB7IwxRe/ikEIP
RzLbGYtOY4ZOjb4YHqKvW4Tglpxf2bXbrQDTb3fFKecn6YYPCjK9idQiBl7ZRUL9qukClHlPXqat
c3jhD6tFLXG3JXZWYCNgKw8v02RDUjEDjTEk6xQlfZ6w/jKCA1TnjtOR1s8nWIltf1h5ksTeiiMO
4dHIW3MGjIP1C5JRUlrZKrLIeB7clDhj/tFKLVhcOlvdW+g9yTevbTSOH553Hd+B8xcGl+pBBZ2S
aeGpxhaQG9M3V5yNQwJe2AXvfHSgsHkeBqTSnzOUFUROV8dYmInbPxUNjxGmu9E0yqnlcLzb9Mda
3KAPDieHj2Cv5q6Z5dnUo/+a5Y3H4asHHWDedbRn8HxCfi/GqhcESS4blsZm88Zl8MybR/wncCbg
6PAXVQpDzwS6RzBskiIHj8PE9Q3uRycBNNZ0Hi4pSv4JITgszUFB/c9S/tmo2leSvEmLFHUkJlaU
6Rz2vwjlXEc8mtWUYCisqd0LdVbjwS0AD7BE0XSLjUk9AtNIPAiWkuoPb+HFbDEqXjnbNcIrUZFG
6HXbxH0I4KwrHz9KI73RoEQdMsrZUz5lfMvg6tbrXvSfElIn9rDIWgujBqmQ5ESM7i9o8pBWhHlz
fwSJh5lxGSOo2cmeH8EdL664qIeEbQI+9EAExNQe/dnb3zfNaDFJfmkAWc3hQ1urDRVsNh8iaDmb
FW/91qehQX+3qCiLTKTV5E3VdBFBJwOZWPr2S7yRkqv20iCBhvBUOlM9M87PVKUrCe9aRaBWxiak
E3ZBAjFqi8TWv8yN6rKQyJhC+wra2UAu7P2sVrzm1TZou7uDDaJh1Q8y9nYfk2Ou2Ea+3eApQ4l4
9wKAkGYVkeYjHwDHtxWvbc5M7R2CW/kgOmiapwnk5wXLnCDkj7avxovqaaq1qEx3UsuuGat0XcgL
+QC7Dbj0Dop7uLrqOvRWGU4GOCnDsttL3riJk+wVwORO9ZK2pi7pYXHFB+ZmWNDHBcAqyioAUybp
h3NvuZHZc95xtta9jv5+cvHz+RyJ6zWMbm93pfHnQFDCylzsEESH7whHFzc7EzEdk/jw05oQ6Q8i
gGgzJew6HSY6NIaY0W60z0sqj1VY7K52wzMASHeLThpxrf/NSlx36lkReEuYFbwA/sCzmXNuBmms
8jo/n9ozaR2uizcXVFaW/gtlevz3Te54ximLnLwq6H68H+FXjzOEDxtN6FI/kBCCksYF9dFZL1FJ
G/50hQHTPT6ikFET+IfZ55Xl34EYTPCyfZOwdsHPtGoA2U7EdFMIlO44hvFLaZjUmxPPiEj5DS5S
RtzUsrGyvTdHrNcrWS9w8AMcY2vFqvqNRAdia4BZY8xDl2XtCYCmeXrBORLUdN7zBcw8CBn0reLD
MyXPjWYaZd+u68eCaPhU0Nkbix7fWFiWF6HX/as03jHpKwcmiEyzhk91W3/Ep2nf57wziBTTs0nw
LCni4wHLYztHbCP7lLdPnU4kZcqgVNLQqWYQsB/0xBBGwqBn+jWLRnxQmqhF62qyqoz1DIv8fYsm
n/Cib+sRPi4Lcs5Ix99r7em9SEprhrKJ9pEIrptC2op7+IHc+0A0n9hlC/oLeywGdZJm0Y0vSKBF
V4h0O6p7oHS6/gFnmF3PU79tKKbVQrOCy8PFPxeing2mp+USNIoPjNNdiDgsGd9VQy1/zRquVWLU
8kZMx/OQDYd7Wg8HwjE5tfC8kItV6oPAeHK0pPbfHPnv9nQ53v5y6xAe3kJZG7MRb54m7gguwSeI
KfZE3v6GzQIsQcwC7ebPVp3LOM0OQgxkFdgklLsBkRi95MU1nCAZLXoOHoOma1/gFiUPSum8KBGD
9mJVZI25h6BvZ2J1P46UVlh7DVvulfVv+ScP5SWGu19lHiZy4LVlcQlOaNmE8d3tjd6OaEPaGF/0
3am9c0oAMn4Df0XWnKvXvS5idM6kESX4xGhkkMPIGIsiLV/zGbdtp3HHi0TsQuMS6gcomlME29U+
OrCT3ZQw2lf5baC+75yo9vs7eiDS7NWXpOxRSQKtzZkpBbFqGkuwt5oHdRpQCOYVWlYYwcnLPNm6
HhLnIzaBooLI4qY0iwYZxl+JqazrbIwh7lZiSOUobWZOXEuTkZgpvbps5V9DnPTHXdOHHnSzi4Wa
ZelCSDuOz+JfNi7MlZp8l77ZCa5IK7QHGvk8kw/tBb5ILEXoveZMLifgHEBY1n8JAlliBoBkJYFW
10JAbs8mOt/0u4HrTv6gLl5UeafzoI7LSTcWMG/tq/eIGy3PwTw5MryjJoxXj1H0tkml9syAP6/p
qQlhjFspaWuDNVSZHH/fe4yCLgBC442m5hICP3+Io3sc8D8S6FEmoHQqekK09KKu53yvI6Q2Oimw
KfLCrRpheZUX7+D1pAjdJzyz8e1MkOvm4N2vI9ZDIgO30xVJlYFwnTlA3Tl36a1wn6YDZFIsmmmv
8pMG5LO0TbiJb//5mMEU7cZABAGIGmi945dVMxd4Z/x/L1aZQpUjooj240LSaz9Q+HMqYWF9MPRx
AipbnoaB8YjT7b1Fl1ISVLPATCsGbfZrHWM3jKBrhdQjIlrpZ4LzRIKSN8NslZbLHpV2PWaVzzyT
OZTed4I996B69EQXdhwP9/o+xo0mu629KRcc1tufwd2PAevmlNo1dRAUbXmP729uqUVgwZmnuhx7
3Fj5oSVvxRtjK9Bc1+my0XLpxi49dx9Q6tUYN6D9SX4dwyUFJ2N+9idnD6sFc5sMJuh6uTB+aAfi
zq+MXTbORrRtACd/uWr+Q860VzCiSZ+/vAXV28+NeylDyFhWB+jl/mQKZaqhLwt9vTQrWf/qdvA8
FAK708IYI9/LLr+zhe60jNWiFYXlBZg5vcvPPDcXloDiYVcVXOGa+IbWwoL8yhXHVGTbDYUKp97Q
WVkZJaCggMHHgXiXpZopmtgnBsJ3YGqvXY5SXvg4MY7PdsYSPcE752yXcPqvAejir4DPFNv6FQOW
Po6USz1sliyh163PsMivW9nbUUu9JLEujKaPx/+9X0O2JUnvz38qqrjpkFOEbd7o1kf/UExQaFGj
dAiTonAh2FKYs5fN5ofs5Rpyn19ge0mHzxFqr31nCYcNHzn8TgEn+8zBO8V9jXB6xfFbdMrqDizV
Tu/aOZ4SUSjJEc7/gVlyKdYcoNwmIC1gCjntYM5uLCQdKjdk+R2Xy1/t5q8JM9CwR4GfeA3dZMEi
LcZITI0d4FH4nJpQ1HYxPbNunwbsbIFfHShaF7GpSPdP1fQYuBlXG7leSiqQQKQlACyn8df3yROD
Lq1EOIDj2C8RpuG4vF29lJoRN7iqORvu5Dh24Xq0twZeNJHzSkWSyfKuOLRDCweX+KUIi2h86zBY
NylzgY5DL/5OPn1Znpoje8GM6KklYPh9BzrkkBycUqtYtVeA5Jx8NfxjRqsksCCTWeK8JP3buY96
TL6BrdBAYNio/fR4HiJ3OjwQdV58TBa26ZkdsHKl5YA3pyuJr3U0wvehHB1M3rxnHXO/8qi91eeq
t56Fe11U2uHNVgFA3b3Q8aohr7BRlyZ7Ai+W4VBbjwbzAFzIkX6V9g6KclvEn047bpeJdnyUTBp5
nNcYVhEKDCvqVHGPZpQoIpVCNoXPjKmgzKevhYX0CcI1QSawuHrMOwSVasT7/WSoMEf0y70Qy5l0
bd7EbWhAui2Jc1J9u1jwmOwy37SZsgJ+n6gWFvqNcT+MiTL9b6kJOF4bGw0js64BbIKkiK4IXWCh
3o4Vx8XTmlkDu5p2GtZeekGcry+AJvh46AG62HpDu4+iKNKNXrRBcylARuhouq6NiOS2fapGq89Z
b52gXo31Eobc873rh7hYEkIYB6W357EPX+weHl45NZimPWf4douRwKqdhFCAilHO58oSNAVNMW7p
RyaG7Ui36exxp9Jb3F9Lddbsu7cYWVVt/PgLIt5ApZEmp7YuLpGv6+dsEOD3jQdHIXFOi/p8bmnJ
30huVJ68cfkR6IZ8/dLzG5+fW4aphIBaD+rKnQ9c7cP72iXRSozH6BqHGrjG3Cs12kPoeyYo3/JV
ahn1yiKQp+nyg0+UMmJXYF+VVvwUVvM8DKpv36hapAYlORD9qKS3eo5yEdW7lGBVmvds0NKezDoa
MmahO+C7emwS3kuCjZQ6/mT2aLNbLEmCEsF/W/VJV2GMwNztmQmf7vFKE0ijYXQFmW1GdWElbLKU
NAxmApyZEj1CLUOAdoGhNB5yEPUI72VpD9VDbjLj3faZNleP2oesi1Bm8pzvJoZ3xseZDnTcgBqD
8zl9hK0NoI5ay8ElZguqg14SeSgDcE8QygDk3SbaHxqy76MPJstsqZWiVmlBhLwFYn8/rx1o7xVj
dEM82c9d2hU0KDOmZBD0/W4nchWtvRZilp9GH5RRb0b4LURtYghk+Hq2o7LMXPmYDelK7v77bLZG
e+Ecnp37Gr4qLPMB+BjPsgBriXu1XyHbRXIpesNHwyax+zCANePHz9OQn+SB5R4/0vHhWVa9Yt2m
yUb+NgZ765/5UFM0LQ7KJ8gLIG5mC1hCBzxxnQFKihuhl0PtyhjTOPNf9608Jh2QfZqAl27/JrJZ
XKJ6spN+jzhRV55rNfFrbvLDsemZYnGqqzmxu6+yPBKH3XTXPXxgQUrJiada1lUdb29vh3RKmY2C
K75SSc5IGSXvJdCrotmqqS86HRAcT0CBOtBGYTGWBHRsPhIkgmmN4PQxrTvUhYWW2RO6a8bIFjB6
pT4JCsjjmW1WG17PJWXHRcQcqIBYcVduA/VZtjqpl4mBRpWq4aAKHOj/aKgtgDreTYwSDzeqaLVu
2WSDJUbwHYV6s9c4mMoDsdjKwt7lVzI1pioo97NggfLBjU+lRTBnoSd2odC056pBSiemizyJBlbz
QwLpjBRepaSinzY8oBurrWACt480hI4lEoGh/zexdXnCYIonauNt1KdOyYtsv7irrJNCB25/2SHW
2pmnPlyOlItsPeQP05UvMX1GDQw7u1hl+lp+uoAX1elj6Yu7hrrMg/gJ4DZMixJ3u/qvDIC4pkyR
uyqECrmSM3WszH0OdShz65G6Lv3myxJsUrSljA7fncWfvr1zy2bRj4KYo3q18zvgIqsxsts9jKB9
ARokmPU7ReJzbR7d5zZTWJfeqGN3uZ8wziUzbc/KtdAboaKHqGNiS7BUsOzMrbuYcuzhOfQ9Xl8/
5p/CotWtiLlSBRJwkiM0vGrtNjLydKl4RvaVUfiRAzXmXYZ03N4zl9ai1R8eInX7Z8GVQDfx1586
LtNlLdt5LuSaCBULXsXwpcjPXXmDsTWHgsHnr641M1RB1PQvcHk5LaJoWUb4OXtzEmVhVAE02SoL
esdWcfjMhopsHdXyVHZ6+ogapVTgWdfy2XhUrcXzYhb1k6sDBd35ykuVQxAr+gzGWtYkt3cNnI2U
x3wctTGMheWNWoOY3k52ezRK8MrBuBRqmPWx0DRq+RHBec1ijdaTXX3euGJ4nMQ4sZ3Y9nZgTSn1
DhRpeE5TrLi4hgkKnU7LPiwWaIbVC9ynO/Vbj9vuZukk0Xxy6JQGDxJzwkxjYXem4jLO0NiKnMn8
zvCNp76qhvM5GWe+0y3OLiXarTx2Rl01CUhd0f0hqbUP6Bmxe/77bfdZ72dwSCZG7U4jH/6gom7n
KJDJmzeLzWu4gYPi2eXdcsofFdyw0GNZkzaf8xTxt9umSTsn04H59mDhwNCwADUaoKFetQw54VKk
wh64YHriIh6cE0NtTt0AQQmO786NtD2KMw0cur/0WWpN/NZ8aiJcf0yo3UuWhYPh51Dn7nKYg2aO
+yfG898qVAO6MNL2uq64jV7Y34m1gUWT6Drh62mGlih99wosXgrHx4zGXVidN7Sx1xHN5Kh/qJxI
0V2z2/u0k3IF4ZUDlFf2v2EkQhqx8r2fGDjt/3ZV+ARR9cw/0I12RMC4AiZTKT4YJ/H2Cx+Anf/y
6PVryhgu/zJzIeVNKfU5H2GC1vz/hjVvDyXwxajnq4+HAp7svVZ2zOgbqXqOam4nRXFzh8u/XG7J
EDciWWGIoc9ZGnG+aEUJW0ohs/spW2Uw13nzz36q48CqeBG38MRXqI3shiHGJ4a9BjCzq0zAQQ9p
YoaGm0PutM6+3wZhHuHDNoOCFM+A24E4XPound6SiIEHZaXTqtpaBo7OabhxThU4CMfT/WtoOX8s
p485/YvwHsu7kvQUZ1qIp2kh+BKJU7zXh5T6f2HqkNGU6d3ed2PvkVy7lsiHs08kSRTwsoA1BXxB
/z8spDaMkMJfj933dFISMmxLCyRPoma8xt/0y9cDAheBIKoJr3GL3r4pBfmmzf6rjbSkduPu4XVt
jo/z6wjYbc9D+SP3js/vIal9sFYUmgXih9iDi6zWn9srgSqaok3mWzyBqEGwOWM8JfIbqEE2HQIp
av7uawS8je0d/q8tzte5KqRVOxKGQ659colyO9MYhiv6rZdppOw7zKJW5AbFi+IIFeB5nvL2UH+x
FVsTnR0KanWAJlnMONsukG75DbjRhFuP+UXDuZRl9ED5YQMSJB7xvAMeiNoLQg2A0eRYXWlrLcwX
/R7Mepe6zlgYe2aPchET1jw4ynsgbSZLy0pQYXce0Cz26bWEk9OnOCWOBb5jOPfKQtSIYI/tbzVX
NvrzPBjEYHvJQqljxrfjLWcWtcnVnYO0M5cboUOnv/aeYKfLOe66eAOKztHRcpiEmtguEuKb7Sgn
wUxy20mQcmKf0DripGJ21smy8NqtdawE+QuJmwm+PIkNlFwIb6cdo6myopKoKEcCJ/O7TUUVcgM7
1Ujzi9YlD3TAPmRJU8VmOGMju0j8PlvxH/U728morIvhF1M4s+O0bUmWlgAJiE7MiL7YCdlAviWJ
CDQAMB2+P9CTLck7gVVwE4gCV8M1BbM+rNyy09IuFbLc0OKcef3oS3/RpVYKP/0u/oZpEdvnB0y+
Ki/cBlLiJyqlSGvmg4s7Vc2EwejVf8+rb04LY6HFX+rZekPsGMicutw9yH/K+VamZRtGJ3IGg5us
mcFPudNpV4z8R1TV2ZFOE/BIpqpuBIVSq28/l00j9OWVKFOaXH6RBJWN3XuBIFFsOCKyUJmgqyX2
UexWOo6sOviK/XOTqHhnae6kkM/9C897/Qeu4dFk8Qmu/VU4QzYC3nciijjP+UtOXb3s5gUqwMQp
iNDF8VOyWArtxWt75L21zcOCJUdvZjFXn4bblExuy9L1djnQ/1Kn7qeAWYFC6nd0lpGpMbq4gLX8
f/U5w7hxpaYNLIyVKbYz8/zkAsJsvCsnTDjr326IbY7M5Gq4D5SVTLqvHi8RAWx8Qk/lU+FbD2Qy
jHNdznKayPXklCVQLFVaKtLOYy5YQGKHysByrFKihsy+jnTp/0gPE4yqyolhl244s3v8K+uc97Fy
Lq1+ygIfA7Py5wxM4e/w561eJDOQS1szUgalRU13NjY0gKD/vdQt4BoTo+qvRLae2HjjN6FTO+Jk
QgLsgfqK2pnhXBCvu8MZ5WNW9mK9XJaAjAM7nsTDWAluLuVpH/6rqvW6VvltQRA96SlM/qPvn+jf
XeYjpCLXoyU8HcgZOpCe4EldtjhZKfrjpOO5VZp/oT6i7OgNIb7ENywN8JVoOBMmu+TEqFb8lqA0
fbHWpjPMBixNwi8+6fGCUD35Wuk68tGMLax78Q9Y/A8nvKtV7z3K9yDq9LdoLQLSjrE1pPHWzMQ2
U2SxumRO2+5DvAWSozFKuO3oufxPJcF1JBjTaAe0blv+kGhaXA7aPAZbESsYtLt0NTTMgFp1Me0M
H/0iokkeD2Hs7JnpUcsR6wlItr3hlSe4tr9hC2o3RyzM2DSkIOP8a4XzSvOffYoVdKyZ3+cjTUSy
dTrGZgDb98bMcTe5UZTIh5OuXwBX9c+y02NsqNdPGkCoItrKO5WzPBUVoG1iGypxPXLn/eTq0iUz
GADZxsUo9N2mfQe0jNLKoBFI75CcqLhVKelcjkck4FdYzjCyH/uyWUEbbZEE2Hfwc+DmEnSkePjL
XIvJVQm4ApjJ1EBLkvSqLIrrllU7psIuPGJDSD8CX3M5FRVkcoNo6aa61WwMPb1yeUQTWU7aN9VG
DKD/fROQKz7T57q3o+rrMYULUILrifhREmXFGRDfn+klPuguDzu5IIqmZODCg/qcuqD0e5MyXJ+S
BMcUjFK1+HM9UDymgBuO26GqOqEU5qQ2iuprJ+88K6CLx/33HGWrZkLvFiSYyYprYXc12Yv5XqU7
HcZZxGGGhdEPadoGdAADiQoLaMl33zu1uo+qHnnD34huNVIcLyut3XHQE6njaT3bo9GbRvfqSa25
yZUT/fB9TW3deLUJF/NXgv1wHM+KaurdMgktjltfsJGfttjwU4+j1S5wxi3F4T2ltOutWax+JmOe
MkbiDXVZ4VQtKaQiETuU6majN37VzhhgJ5VGz801Wy/8YUvaBtxyxyYhXgbFi+KajhN0CWO4QoC9
xSCVMx//MB3TbEa1V7R8PKxhu2eN9+MLz5Bds4fVSgrKbbNg14UDJ49eSWWCFLw+TaUp3USHV1uA
qg22A+LpXIjAQMiDdJpFY8UEwbEnnqCQXgO2znHvv5PqmUdc3lmRstWUnjX18sX7DiU5YVNZ8yxQ
9WVOU6J3pJj7d3uAVnIo0KQOJRx0QMDmVWQAwSLePUUXbqqp2/0cxP87Ha7IwWALmVP3pjtRySxP
ncKKLUCz06g8ruY0nc02mJVKosqs23WZ36a6qJnNp/SfpmSZxwnZXcxCuinJzSeMoc0eZpnHrncj
uncQIAbdzEzb9R795LRE3qW6Ez0EcUG5H8lWw1Bx/dcJ9mBUrOQUdZ6WHSUmGEn6yPvbK267IPPH
2W+L9eJpIU4VGspKf5ro6CngQ0NLlvMw5keS+B8YPKudcks631LmPuXo+9yUJ/4b0cok/jb7W4+s
PDk99iHicu3J3HsdCChRA9yLLd8KZQ8BZp+u+q3+Kv5UKF0a0RII/o6XRw/nfnymsxUVjGxKAW9z
XW5/UyFOspCLWeb24owIjcuc3MTwReIeV/2+VuMmRrtKnr7wzqEuW+/dcn1trPWJI2V8Ja+crb7e
2uZ6lmUzz0atZv0Smfy8hRvnothLaMJePVfwcqIA9DBGM4yC31d75j4orBrGZTPPe2zzQyU0kSG1
j7ol8h3XXAbzKUDRBb/DlTscwfbTz7+GcX7YSRvDnAJr9t4PVakEgUQTRCm3tmbO/JP9hSwMJgfm
LUhHDmRA5XSrGzBGEiFbu7aCJxDw5VFp9bIf3wwQjkFnk21Ab5C++YWYtHJASqE8oeAuLAW1HWAt
/w/LGzJqqGL94qyBB1usiHf4SSaabpnpuy92X1ay+y9YYuFN6TjQKkjSe/b945nQmq9ScSb8WGPn
hyNHR5yPLX/fme7uakee5IwA9HK9fypIYZhcLhKdSRq1cKchRajoibHx3EF9dW3xXQI62r7f/N3q
1w4GWkudh2ctZqzABaXX5s4bb5oTRNN3PhoweD6tGPHYtL1G1J+1V0DHiP/MapbDUlYS24aoPVc1
VVwlklzOvJW7Pr4fw9hVyUQCr9NeZ9FL6MsfiXshGYW/QsdPCihrQLoMHkdhNrkCdGzPhWymV2WJ
5NDm3+/0ypbLDaV1QMCFTTYTWczRhRNHCphq/AW8SawAIFwd8QPd/X6c2Zt433pXfeU8mOMGyHKh
yVtj8wfLvsNMUh5mTZmcii++5El7qTiGWUHOst3vCqH1wRYSNCyFhgESACAtIDDc36tWIzC9s75h
beECpC0y11/aQivYZxojeAgzBwkfckW/V2aSjF7gsALqoaiJImiZzenyZUId9kbyRYPNzVKKmixP
q4K/cRozPwgt96ycHZdTeAV0DCdMfbcxznOb3Cz3VZGXiqc1ijGFbOGi6x6L4+eU9k+boKwoha7G
Sg2/6WYLpQace1Z3WF8aQJWUfu7RtU6DRAFrQJQBizWJ9WLY1WdvCf5uG0cQbkNama95V/3D/Ucn
k9C53itcM/AJ7Lp5XSKvjY86xeqilzRVS1MaPKaRiZ1LE6THye5A9VwKCERs9KJbm8P0+BPiFdHv
BhvEGOSsc6aLLeaAhlw7Cg9A66D/Zf8C3MspeFIi08+KJcdDmjf6UVKTH4aHztky2JgAnjONYFux
KaeesjnccWVSq5lJfqNkoTegI8aBxvSj+D0ocfgMyrtCSGQQqifcatryQmA+uzgs7a5x3LHlVAR3
x91SkHM1WnK9G724Ka65KrBzW7aKGQe7niEtO60mYZzq0x01bOnT0jUxukMGR+rzrBwhlSqw6fM9
VCT+275DQRV5g22MvZGgZR/vFyMe4sKWJ3m8cIqRMDPHNIhoItOvNfuOVPH9IL/a8faS5nrDgPMw
dLavkH7X1BJeSGtPriMiy8LWGU0yfp8AYL9M5u0Ur1Ys2DuGcssXLXDi39Myz2rmUvh6HmGeKOv6
JB3F7VN3ydGRNE7hzzkrDtti5mBmhbCgar2o2IcNHzS798W63ABLNxtCXKiShgIHvFKeVUSIZHDx
ahT00UJy1gLQjUG6tbhxQpXgiNIvlCEinl06l4vmc7dx5l/IQwYCxpuWlIG4QWeYdCcLZH+2cZAu
rRHf7gDJXx9HZSHpVr1Ez8CjmWEP+COia9LJ3nb7TC6TgNwoZTXbdM5/3Yi0cSOFWz005q7GTWp7
IDGt4Lx6DRpUnYJ4ggx485f52bUz3JUE8nDq5idEKXippqlI2r4lYqJsYEM1T2IO5ibMv5d5FxaQ
lacapEVt6lr+UNyqAewG6ysxHVotzypwGHzxJq5Vc4qsrLvffHdRN1KsuocBmx9SMlxU3vy5oI2F
p9j5j8HpKXsb+P+iNFrlle1WGiOExG828Xv5H567wntzBJOG4oNm9HRCCIgdtY/xLKCURf1QOnaU
DVGaLicz+skrQY1HO18V+BJz0Z0Iqrak3G6aUHV3ItciTqRJ4im6Y3L/VEpsxUrq1LFXTAeYi2yh
uRZ6TZ3U7nniCmY6K2aXJtYgbmlABk6E3nsiGJ0qURBZ97k5EYYucsiU7FtRbPYRZyKQWJwqBCrR
zgR0sOHNgQQVCWPFB6R3G/4vMYpgoxSHbWm2d5FvmVbY+BwmRR7FfrN6OuhQqgiLg+09nloQJ2+f
Zd/SkDLvW14cnEtjyKExVghSMzg0h6Q/f9//eu41lVuAGHrWpxSxzE/q0MZ3ABNlbb8HZa8DlfLw
ndXC54Py99XsvKsSMzWsVNs2N9BjH7a3LMEUihUC/BTYnRB5H5vBvkwNH5zCRAnGVbvqh/DdUXGw
p6wC4N6q4369RxOtPX0llELrsnduha5e/Bdf+tLGppgeRgp7ZxQ6YO1X7IfVnlgNkuE1uForGHlz
u98tGq84nRX0sgBxTfliWk2qJwVJWQWjacq5aRkqxSqtU/hXwpOhROsgscf+JzTej2FnWj3M+jDN
oxUcmq/re3V4k3ERXLOL5IWKLy5LfRmffgRAJNIZZBQnCLhZv6DdW07MZRxBPCvw2SPBDzHVYf51
DMsh7ZrVOw81r2gLjmtxCIFeXosc+46A7sEW1as7SPCoRpTm/QHuMzTZ7sA32+Q+lsG30niT4JE0
UkkXO163y+8V3oC2ubzmJl4v6/CoJvwDK4rbZ5qZdIlF4UB30VRczRDQZqh+o45ZRvV4yldSIxMj
kmCV2dTmMykekXVAJNFEqYPavnFl2k0pU6jV/dReZJA0cDa3yiJhZVEYRuwx3OPFWPnoZ9MZJ9gG
tvqYk4fCKvFRiKhhNL3GQznKQGac1DnRaVaU6Y/19u8R2IsrfUyu/IYGr46yB3mb/eMH0fMO9OIT
8RC5QqdFVjIJsjJ+eQj4ldG3n//2TzNl+ehDvJ7La1xODXC12SMg0i6A2rNTg82qnlHM4OI2X5o3
Qebf7lQEVw8XxFNAYFkwCNEDpXaQpqQSGGvNa5Jx4Wk+wIhNYfSvfVQ6eRWPAg2L9if+1JLaarrR
wRe7GMiS9XNmYISFT8/YInFYasoeoIXhpouscWfp5aIWFEQRYtuyCJVEk1PkP9J7OKzOrLNjQkp5
EKV08y7DJGRWaJ3USNCLOAvlAg+j2ltyeFmAYANbeFbK8f9t/dcOJ/DJT9XfDIWNZCCPUCOyFKHi
1yYJfmUrnP756rUfUDIbNMT7gGy4PUJXthOKvo4Ycr5CBSl+8huAr8MgfJBuLX+iwcs8j3IuyrkJ
KXLgw0yRjTfMwZxtq6OjYcV5bEDqUYaD0AYdOO2JuU3Ajk1ED6SD20TYep+pltn8CYv8BXVZSP1i
Mxt9jfPmq9rD3LeP2Fy1cvbVyDaoAB51leDqsbkpBiAkLTIFezQ9R8ZTEvS8qT93l5bZsh44HzUV
QPVvmamNUtCxRJIsaS5N6MB5OJ+zHClQuJXlDLkbf9c/Zocw3Rm6QEi12Y/ETwQ6uo4qzEPdVtLp
5rMF6VQeDKxqpVkA6WehWHmPawLb99URszOKKzoArUNdGm8rVlxc2aGzhT6BGav9vks8OhVMvD/E
/KbLMxylg2aXJpBaewsHr+rq2mHx58YwVZIlllgJSWrAXTNdHjte/cO/5WjhuG08Sug0VanwsPtw
DyZphiWiD/ApthEpMS1iCLHGqwKlmqmHr6vIW7Klh8dKsw56GW07uIcqVtUwk3uFnkuaRfN61uVD
hcIMppif82n7673d2dkTjCc7Fj6jJUdLDDEteE2NkN7NbXzrDsu67O4shmtOnlkVLC2AJHU7dT9w
3H4j6lcOX8DqSNv9xvcjmlky5n4bzFC9g7FB/p+9D6ul/UJwbw+YDFHxXA5r76FVXknNBtsk89g0
rsUlT6Qy78I1iHC+29X6CO5x6FLonrDZfGYDILEHPh+ZH/77a1bt66Tjj7DjT+VeaJOzXfAkQZRx
NCxg8Pq3ZBRcyJkuNoWW9sDNcI6YGZJNxxVQihWh1oLQtdFO98j5fArY1kF1Inj7rxmryEWg26wv
EXq07dl38ePTRH5RRg/7Lo5DzZtuWrkqFDVHgIEvG0CaLP6tKcLF1Th1wSS5kMlWF2brRxd7aXSd
0Qk8Psb0BdZj2AMvjYgN/R3apPfGk1C6I6ww7uj6edf6dNtJLHFWWKcU7CEQRc4reqzEEXl+abWw
EhiROozV7PaseXvsaM3rXCaQXB0AuIWGbHAHaeiJ0xHLDZCE4HsF1/BKV+8/5sz0EwGga1EAxGh8
vO1GYYoX3eFORUI+8DhO2TXALMs71kinEAEggppW4F57p/X7pXtrn/S/j1tkwvD3wDlinD6ZXadR
zFpfRl6nXEK9UlEZQ47okbMeXd4c/o1pZsmC89HWgnPZQBetj11u031aMOzirp8ofxe2nWUQZxjH
90uQSAMmG8GJczqgP3VIIFG6uRW850mmFUHaNDhxoCUYpgygwxGQALuhIJ0vOn2WGEr+PHiPzSmn
fI2qvlv+yyM1LDmxEgZM17HRZuibBF/dWLzC1NBvJ/lD8rVbce6EH738cZAbkcLXmFM/1PmQ3vji
17/9derYEonqEKtOZZ9xuwaEqceZeu/rVjy2JfdpqiYZ2RTZD24A70xI3D7v7OgkOzNCgGqQcTPJ
ACVixZBhro9P3FibxDxJIak9uFFNg35RsYRfG3Op7z/JluG/mzEZD6oCDdboL2Nig9HVxMMDArGM
zBCjZyWO7CMWwCIk7RCrtT71kT8LFmlFbu7AqcwYHWOhU+OGeaFmurbcZdoHVgR/xIM5CCKZebp9
nygTNXRMQY4nYSz2OZfSOLnQVnqIO9C2NRvEEr44PzzLHLw7fqSBTtQbYQaa5syD2yegVG+m+iVn
uDXB81TnSHtduNPFfwNEbeuOchtSzRnOvRN/6+lDCQN90HwAwhSKj563M+S2EYx8xPcjn1tFLeIa
rbFFabGZR8IrtUgo7ETKtdqCT9r0AJHO+iov3vLDqWIXEknc7OuMwJHYaWEWfbVGyGwPuW5EbL/J
U27JZuybBs2YcaVcwTCdxMMmMtsukP1FwiAZtXLVSaIySjwA8/QF4KTeo8jfYHCfhBZgMsxF1oOC
jIGv0jY+8e4qYJEppa/TlYRur7r/8NO0iXxfTAcBZ+djgr9vqNyMbRBCuwbKONcPkzzVKCbz5Hyk
XjeN23W1W5sSl72Jz7f79MlKo+YjQoLs0ccGlcR40+S4T2bxJ1mULIuS/BCZubcWnYwIHauIn2Tb
FXFaYiDQQHPI6cmj+B0y+QBqLfIW+tmB99DXYAIbfjfvqPQU/aAmWho5A8kfsXMVRcAtpIP7Ilko
B2UgzXQfV+j/vb9Ix3euPHZ9fGz4psTtomKwmqksAn4Y9j3nIP4MXRrpnlsR8yLbid834zlkEfYb
sI2O/NzMU9ZSyweF1v2rem0vFADUD64J/KqilS6GYGewA92sHBU8mN0p6+hnU5MUHaU3TXUENB1U
uWR2y64N3QwBP1ePr4UlFBAg5KCXO2wI2AAqNOrY4GcQXq4vP/gtEkvX0yBw7lqNAoV5Pw8IowJP
HW+F00MT1cp4RXCg5OH0xgKn+miNQ9AExlY3qjx/SH5chk7Ivfyzs/f/acEp2xLSi1YNks86d59U
caMGD473Xd59WjGRGZV7Wm9/QdUUgSiZcgeNCYkdcZAj3B0SwMwPKrUaNcfyZb2W6ARARUo4wcmv
3tUerT+xe9RDfAMTJQvGFCM+AabL6lXOD0s+aMLMkO9jNwP4nTZZR1RYzOxCouJ8Z+W+MTYFiYbR
SAxseuDeiZ3lwcG8xXgvCiRv86zdqIP8H7xJfCPRYcO0KLE46LbOWXRGUxq1V0Xl9SSgGuJPUuSz
2EVENIjPT3GO2ludOx5GtpbVFEQQOhrtej029jPunzsRYK5Yy2AO3Gb5vXln59CCcfVNmCw6ylSA
XjA8K6iipDlmNu3jKrZsi+Q/9ylEg0GNSn3E9Kso+DnremPKIOl4I1vj8m6lyBCAhJXtyyG0T7o2
H7Fzh/WJil328OzgEWKNyJ7hsfcJ0S2Q/a+ZLFuEwsoDe7YsVNA4NrQqd7lRShKh3ap4rB1JujQ9
4DjlndW4MFHEgtESK+5Q47BBv/OpMQrGiF5UmoKaSgRPJa/UIU+hJ+ru02jQVDpzpaQ1+zpm560e
MtgpnQaJYepiSwa7BOLf1ikITWyYcrcXfuauYJWYazr9w1hOY+krC1Tewp5tDOtpR8jGQddSqHIt
mJFsEMh3rFDb3ElOoTf8iosvcQVzsYM4xnheI08WidLjqBkWgvvhG2MTyvVuR1ADj9swvDL7XFto
aZbpGcq4AAGnmlS8hPMhJELxkTsLW9AfIRVsMPZxLbeYEQlVVmlW6IA1/o1MzR7Zt7Pwd8voBTsy
EHyRBI+zppxZ9Zf1jnSYOyKbCbCvL3Y13Agj/SNyWgemTZzx3S0NZSQDuayKkqoAEE5qaJ9qKrS1
CxvYhqloduvw9lGMv65DPi/S241bOaB2AfsUfZd7Hw0NtuqOvZg7I1ryl8m7zirRNGlt9YHagWEN
wIgUGgV8XSZFEyvLvddO62PGdiodaTX3rolfheL80QXtn31qv+EsBQdrjySewBCgy9pSKUhkHAvb
qSZpMoU98xHHYWIdAoF5pRT819OIBZWcdNp3ZtJ6Tga49p5pP6OIz8i7CgSuhYuocxWV7jkJ5ZZD
KR1PV2Woy3rziYYO/eTiLrdRYHLl10fQ39iR5eGkZDUclPzFd2akybfoTX4d3/UHMAKxw66LgfuZ
/41Ps9x3bTvGYvBvAovxo7y1xzuxe2PTD11N1tTAXFa23QryHoJ+iEncFEcvU8wAs435aRvxfgET
VIxqQIhzomj+NxRlb7Q4Yn+QS/ft0knJDVB6nK5myhLTJj59+4S7TrzNglZBj402bUvB78eHD3vP
djlAJ9yAbCoXKXS8GyPk8gZLaShB0mnnH9G3uA6FN59ziBYxTiAc/to58+XpjRSoW7UtzUu6Hde9
PoyGBpW056EjczrHwJz7H/gj1kbCbsYhQNPer9cJfOvd4gj/YqeiLJKZxVGO1rT1qCAcm8hxx17d
/JYmdCKxfmDQUdtCwF+FcpwTGoksncisXF6LR9Yp99Fbt5gp/++/x4TxcsxPvCsNIroeSSLz0AI1
2VuKLhQ0by9ie77t1BcpbZpLqBZ4gmcDyB6SBPNWaFA+U/DFvuOkLx08ths3r3Q1Ls8rHQhlQeUF
awVcmi9r9XCB1PIn4cTwT5GlyhexgNQn2PRtDKRXc7UDCUHgYguHY1nnACqUS1uSyUhGDQpCQ6aH
FQUi5pHGk3koqTawew/xs4YY1DGBAWluUJb8bMOZFgLoFkBUEadYD+chBia3aRytDqhBEbQ587uS
ztBT8mg5JNfNngWrl0V16Vus0cc99OWWBiSGD2a9/h1zC053h9miZK2hW0BbWxOmmvibV7cH0koN
VSVUgfWrb/vouVMcPT1cX9/lIt0sb8sq6qM/9Co//1CenP4ReX8+au+7oU3cB6w3NiAZ7XsCg8zu
eTa2YCazLZxUGLt8QMZ9qv/QlZ1nd44vGF3xJH5LuKrk2WzeDuz5z1p+oIBQTGdHhmejXygG/AKB
nrtYavUul98TmTm1q1QbESakVrY/3bdn5VGU9nOvCICqwVtOQ4m/zyyiA+9sY5KiW9cHDhFBNrgz
r5qZqDa3NlPQhyekquav5GAE2cmriT6hGOCuVowWiKr0UqCuQZARjmtPJsiRZNwH8a12MYcqw9tm
WlyO2pnj7A+VOzhWGbv1gg2liDAMk8Vzb+UhBANHYAzqEHmDz2bZCOrscrS7MNQIq1KydoEJFUv+
p7xqRqgyJ8GeYH3VimXO7kgUswqSK7PIX5TG28dRwkq9RCUp0bJIqo0eqZ37WZRqJ3Uy8dWAa4Ea
QhynOGFJQ5R7YjiEGLpOQDsG4Xu2FPaaJ4Ce/LvOGMkWpF1xj1cYl7CQkNVeDhzjZNd7WrojfP5i
BWiDvJZZuVLX3/YWK6VnY048829hYdqCmFIMDBVhpn6x+osGVDp0L0jnryZ9U9AFAXQPn5hc4IgA
4hlT6o4FT8qaSH8tjrvcRXdo6T8wH2MCS0NFMa8LqKKD5MgdqRjXvGq3GmfMvgC/Rpfqb+7NB3YM
MinQk/fw8MQeriACDZF4vBG/0FHj3ae8QeOdavZwQaCqDmSFTsxQVXEz0S2bRv8lQsmEIv6O1G5j
c7abeuhA9mOr0uR7OqBa8t7r+Gpj6/S1idDniLAZQL5PwidX5ZykS0ubEviJOVG5s1h6KZiOHFAo
kh6gnSsw/NcRuGmA3RMgjJUwHZJCKlcGQpAhDtLIiqjApz3ZxxG2iRnTWIYAVj7ydHWADcC4b8GI
jw5MU3rBC5WTtR4ajOq01u4lpBZ5PLk+SrC3KzGo0vSjF6GcmmgP154pgO5jmMuBRq8KarRY+NJQ
N2xL7Gj6YmIE3hVtAAvRZlq2VGjEm2yA2Z+fM7YJAwDwin1KFiMMKdsV1ANBM0xB1GDhDqOIxkfY
O1g+a8Ep8XmwDzJIXgKeAjBXedt/MtBLj9tRQ/YDHWcVgrZCX6NQ60z9Ji8B1SPDkzfdUILoat3t
c3Gab0tXfR4iDQnE9ziemW9wheGK+i2FQHD9+C8EfOjT7/QY/WJfm9N66QzHrmUeHXQNz+1MuF03
ghIGVSfQFKwzwFr14pIUQdutq+RWRf4Fza3pA3wa1SSc8+umRebM2NRjV3CjOJw10PlwUCEV5qJ9
vKzacNzggqFru4RQtyE7E/K+Dljn3hYRj3egOwdERGFCwqYGt8VbToGYAsUI5bXSy+Ph6qpebWp4
09peK9qowOyk03V2H464h2YjjUiRaaO1HKmco72jBWeBg7VDpq16AwDbTKHYLdVZoX5dgN1gG02h
XoS4r792IZ1moJzTfYA/5b+YEMCOxlV+m/4CjfLebAPTTesF4H3FOzpccUn2AItaG4gsiPJCjC1m
j4Xy/zoP9fAvLfjhHn9V8XQWtD5DHRXPoOeMGiakSssRjYsdXuTEjGL79T38yIZf4qIZiMcwvq7N
8L6atxcoa5DDk8FBZa/VZi5E50iKWXQ4a9sfM26MhO47bjKKFm7djuhjth2IuQPQSm7WZr7KfsDw
0IdblXvAjt7K9MROHiaUWPOjyObLa50ozZoDIixpq5hsb7w218fkw1F4nH5h60LoDKglWS1brwfL
q1n0zQ6+1tblk+hmVBCk0ABTf2hpp3rr03YELpBXETsQ4bQQqxLzTOVwAQhKTsir8kFJZXjq1TKF
l8RAHgEgtCSxGUqpnhe6AvV04h1OklmDSaSKiMOg4TEu52prIWVjee/FEDCWyAlQ29nKElrzBWM1
6XLmCimzodCOuCv2IueQxedwA/Zka39Eo7NujQMFKQvEJudII32ppQq+JjwvKJJleXdAJYyvtPmQ
gvRr82RJAR3uwD1S9QUCzPWFjoIDAROazyfZJm/Bt7VRdyzEYJfVRMglllEDECCR/vZyKqjTnCKt
RNwc0VUKQmOi+PMx+J/ptHY2l/KqMUHQxM622jDTvdKJ90v7ByPu5b3rKtpb0nGLvmgggolLBdln
uOLPAdxr3PrMufLJzANLIsaFmEz52nC2uDp83SSa1f/u8PcD9Mje8YDbHKZogKwiX/DryoSLFYmg
uWiuTeJm8G2GV+Oe3isV+Ka0JUItFCs0drYoe+W+hloHFhUmr6EbZT6LJV8/2lU200s+gzh8enyh
hcniNacg5QGeUuaUh1ztfbCn1utRG8DqqyRHosqEQuZWDROCE4reVHXy9xy7KVVUzaC9z2E1tnYs
oXqBGSGa0vOLo/fOnU91/WGF1qpoBFu5DGwSQM8+UZce3qi0UUSXq11Lb9+xtu5O45zECn0t8X+h
Dr2HfhOH5+uIBeKEnsiMwjASfcyscsXtJPZb+ThM9l7+w55lWkWZrIsOyjX3/l5n+0Kp/uMnu7RN
TghXh7XvKVTU5boQ5jcREU9QafZ+nil5JyBZs7icdIOvAxlSVSQrP3kl6Raz+lNwr/oKIKa/OTrq
b0CUt9SVlgKYSRR2BSqZ5AqTf1ZaBGbuo7tHDwPS7IcAhNSajsr04s70DGNYwEpTEQ49nILBjo6D
IldM94u7VbvOnehVmYIGESG/irOi4j45n4VxajF4oRZ7B/cqzkBCp0TtJgGCJDORdkQBmon5cWJt
vohjt30kmYdc/2HOhyISggNaFVeKLCkOCDmGpuM6lC43iWPt+gREmebtxLsgQb21zEgYS7hO9SAI
gD9+3LVwP/KhHgsy/f8En3omPnbqNMFjtLFPjWrAPv+oGHipXsu2XevDsWo3YWlH9+6bXhvbxPYp
vsJUmrU/dCBtbcDpCx4KHLg9H8L5WxFNgd/BEB0ss02OlwsNXThUgfDeXjnsX8ZyHMLvxsctssL4
+oVG98vEb2Zk9lMJaFGqiyErVZRoMlnlnbEfSm3/hxm0MwGV5wABjLXB4ZcJaGq6BwQUlJL8lCBa
4ua61zbQh8/+lAZ+pBKzdTXjH63U2sXdwr5WjsPe7KUoHyQ6Hfy2Miix7ESL81OOnCc7jsG/X+KT
YVrXgS/AsGuM9SRGRkFemOHhOgAbyT+7RxiyHadERrSDUW0eRDamAunG60R/g9oILzYTrtFZNaqi
6jqGBVM9leeyV2fPtfWI8lLlFNZ78xk5o5iNV8V5c3B2j5GKHCtA8abaEG9nw8b80EZko2m713Qb
f+9g7lNaG6muuzAGfWhBKQ+f/TJYJYWojED1/agCwapwEmW+x7SfBl95EBthmIsuLIMNwDa7Wmuu
3WI3HmdC/o7hc3LlUtOmbR83kj4omBqSI4O7hvyIhw86z3Y16PkFJbgqb6COmhWiphSm0CMI/v6Y
WpNrr0VcqgSidOKXNOHQd8vga3gpj8ugh6VKLKWoWpd+3SXY1pR/z0wdSPMJE6kLHGDLHQWYQ3Bx
bERAaS1Ds74Zlvkvou+xMTwY7FGSFimEZAJIQpOQY8zNbAqFSUmcz1s1w5D5QKCs4dVV1EyXfA49
rVxAt4HKQaoApuu0ZpdqFmdI9hQl/vSuLb79oEKTEZhsLZYTSqqTGubCFU5HXKMbF3ySd2rztJvD
R+yG4eEdz2xpuaYBVfU/JSD1O5vKWjrkCUBNFwhtCJbOs663Pfku8sNfP+aLWVQi4VRQKSA7QVf2
K2Jl6EKe+ty+fgbgqUHYhWGiYhfQBevoTBijaTvtlKDXS3T1loqKJld3zs8Das9u0xqV1zIuxKEE
3O0c33Qn+W62SEJTsYyBLdDRJYer0XhjPZtp1PLlKAa7NQMRDaHyYGy+c6r4wUsIf7qgzz0OtqsE
GQOjtAJ1V6hlONrTGfVUgeArWVkY/y+JwJM++/6tGwuocd39FYUJqnPdjzRhY4CUVvLGGwBfJXJv
Tlx+DWKSYRUhzhcCt4z7uJ6bRft/ED2yZRure52R1sE4KhtE++619nCBuV5Vzd0xq4Gl5AXfaXDd
h8s8OXFBZj0zvzjQ90H/S1CiXd0Eq/00T43YwftEpdRw1m97lYAVoRXYmOwKMg55Pxmc3KalOqhm
qppxd0aDSHxoPV3YhKm/xGBtm6XFiLdvNwBwGOB3BdJDWOhvPsuMww7eU+H1/cOZCCnNF8G/I48C
CRsncVjL08fMGMQpPAOGmNfGSfpeTsVrh2fp2OlPIe+K79xt2YWZzFLLFpRrJnx7ev7MnI3n4SgP
nFh7JGLHxWc5tZdZ6U8m4UvIIwV9mEZXQPKFlXPMJy0CzkxVJ1Kjw+9+gNls7KNIUjCiKkrn8lSd
ovYfmzV0D4qBl1a6l/DDBqgXilaLvXMLmbOmT2U7wX590Y9jfDk7Z0WL5tVkfPP1Wp/PCtZw/6ed
GmyBDT5F+hkqmUumb+i4Hupz3MnZub98aTDVb1zz/P1CvveSZfICwMNM2JsU6XvgUoNkg5IXM48L
NxduM6R2ClxffODPgOfLMVanRQi+NIOGY5FQXyEz0HjzpAnt8spCpjp/EkkWNHZioamfE0wkjc/b
2FcrahiaCICGAK/Aqx4tVJCWfGgiu2IGFiGR9u+MdWp6y0UF+481+gkO4qipcMOlxX22hBwPMrI+
3ZEdv8hHDJf/MmJpsLng3/n4sY1kmJPOl2Uk53GQSIVXUVs3SZ4VAjtzyj1DOU3fA5UvZIPdiz9H
CC+ERlAhmKo9zXRqBTUYcXBe4gzrM7ErjZE/4yVK4U5xPjbmevDqohXJAA+twU/vFbK+ylw2C9hr
6yavj9rlKnFkrHaN3mN4sHHh+FOkGGXHUE2YUX+NxGA/AC0F8hKNNI2nDP8uAOhFsXgv3RUpUH5H
Ftk6UlLUIk/tXWxOXHvighrWsMOpVrkCa/wX/kXCb3YgNKqCr36c8TtcXtLfa31sHTq0K+ny5RBS
NXh3JwzTibJMSYEK9MbO3aluskLa23e7uUMAgh9T6ISGOCm1EBZ4TEgJdZ2XHTrOvr/1MTV5IroA
NeSWIVVTLO9fWQGuWBJAv1yeMK4iLEmIlCbdkXMt0KuJZCgKb1vKm20icAXQrPahwFNlbP6OHaNC
l7nM70uXJqS8zRMC6yqz3O0z7SAygZXqjxdtBJhue/ZoHgaKnAo3xYrOU/dM7f85zEfUP+gdXwE+
HId6G7iy8bpsssg4LwWNvTkH5UtoETSUqxQBbKwYgPI/47/Rliqup788vywgTVOwqpwQyu2ON1DW
HIjs0gjjdeDrgLa4KeF1tUjHtHsiYCaNKweeGdcuw67FLVT2gznLYohBPghSsEWMLOrcFkiudpuf
ynHj5FrmlPnFutGCPAhKNe0W4Jo9mDwJUZlRKqWVcU7Hl6+jvmjXAFbe9L/XrWl0Mw+T6rWaVnXH
p6F3yoTuRq93M7tps2QX8M6Iy/VPSsDg70GcTlMhF3kToR76ellMyPDhhJp5WYtY1lXynKNnqCmd
WA80xuni2fbrhuRhjrfdvF85rPwsy6k1yot91rtEL2nAF3MciiwPWwju4DrVd5PhWlkcR6Y4S8fI
5y7YTN84uSQxxmUKNfFDDKgNONmWig0AS2/wdC8w3DpY9d4iF1ujPsqtUVpFYhlek4Xuiq9qzGhP
PL46nmK0nAXqzgd+iclakDEndAH+WRPkJFUHNllPkdAJeLuC9vE2y8dMZ5rnx5R0XYA4eMZIlOh4
v6BJpUZjQ4lohxDStiQZ0gZ/Ym38dN522aJLIGFtN09KtCOaxGfLv2xviJREC64p7c+gTRJGpuX+
WUeVgfNN+NyGkNI5yRRHLifbkJjUObbUmO6bT+TzLw+bzk9Gd5ajjcC3Ux3/VzKtRS7/2bJ8tKrJ
6QFz4r/IAVIy3exSSJdlJ6TL1ozxG2TY2axXtomnzQLyhLsNNgVz3K/CTVRVzfs84AAjT7zQ7Wy+
/FJcnvJdJCiDyhi3SFFcRYa8Eo6/KjLqRMAXCV4uFn2Y0SgPDQ7cfkbOjHfYiFKCVcMyCRPRhCOl
xQjkSJSn8E+zIVJ3ydfNjSrRFjx7IcyWviBd+dxwsQ9StKAHQ4Q/i8WPCdXzrArnXM8m5Ek5wLpu
uQZCKNqSf/+CG2ewnIiC3uE7x8hjzFkZ81KSYUiZNvd+8QxvD3snBowVj1ZeijyiX1B0UgFqySHs
iM2Z/r+rl3i4RWwVFta2ER3zvq83Ip1WnKLh4b3SCpOtjMjTBMpVHNG4rBTt/TQl66H+Ofd157/3
I319/qqOA8noSQQjPgIdRiaqfkLl/vnOsD+BcScbalulsUydekVp3utOpPjSF3KuTA0+9IXm8OxZ
GZzwOi2ic6NWNdBFw/f/S3odbfaYin1XSJ3JnbZ7MI0jLtH9clkkW+mvMFpz6hpSH5NrTdodJGQu
B+2KZnr+XvKkv1abbVsD40wWd3fBUNLy2NHhGR33xa/nPQ3ami7li7iMSnObw4zT4LeOqb5MqeC/
jU2yUK5TVtudn2kK7S2gr2nuHfm/js2/Ne7Evra0E9wYfmgWLEhCovLSGEP0fkhiz/aX1yFnGVa0
UZn31snCIdeIBTA5emapF2ENHgqcM3LJ8rEuWVU9s5+B8KpAjLSg2g0Qkz61GVfT362Pemc/voNN
as6xamiJ7S6zbWQGwEVzdLRkDjf8bG8fCECrcyzYr3HS5iY6CMuLTq/pMJpd90bBUJhPiqhkxOw0
hJbdCMHl+iZ8u6xGoluEu5JiE4zsncb2EsmYHDpckVsdbWsx0f4M2sTwsQVnnz8PUpdtkie3wP6n
eJFxz/e0MwLdsRFrL4lxkxLWSfwZ93tjBbn+2mJgfN2s7DXKwCc7M/7cSCGV0rdm+I59Fvu0vHHr
qsOm/TCaOSWPS8QW6lJhqfieZxAdvXbYu3H4qrM+MUTWLCF3SJFwWmBn6vMxOwIgrc/A/npTqdbj
/qWD/+Iwc2UF7pgMSMv8fN4BaN3jcKHRq2ByHO4FCcYn5z3ACXMJvqdycwr1KfNxDbJhIVhVii7H
svEjCeUOBB/tIhq8N2KLWsGLPjGgc0510P1zW1eIvMC4sRA5LiBgOnBWZLGDZ3BWmMCNxus8HZW9
ktfn8zozWaVJbfQgJCEBeYwlGOucmeBLcrrF+TOGTVzboOz3G4lnrbVZ1yOmiLEvV9RvmBh6zotE
ESmd/QSDVUNdPBfHpSv44TjoGMpdNd93qU0wCJhCe6TVcspk41U5/JAIfR1oo/NlMiHPOfkBkktM
Q3BbUx0gciDPYNRBVllXWguLbP2DWNxMdfGIZipqzNPn6HlIy6nTaNQ0RuzicAnkon+wFKvySAUt
zLIIIr00AAHh9gCIehV908LvwLaL5pFnHMKoGPpaD1ayo0oyCoEwUfrEQ8y7NUpCm2isesX2gPUa
T0DdDPs3Lu6edTC3CamO1Si/j2zg5gOtzFp6u71+Sz9YRzi4genr73IeRR7yNGIpTPhAW/jBulwq
ub927FLa01HbV+2cxUvVOCnjzcTTJ8frRBDEr6mb1mL0+8DeLBsfgfZE5GME6j8Fzk3ZJnd5cywV
DkmclQ13g8ePUmFjAgN7Dnvwqx9HKTqrt9twj1AfxWsxioCPSaheTrsKex8dsTyEoxtXohanmZeM
VgOnMs1cXD5IJZbaqynYIlEzELcM+zwXyyHSFk9qLJU3vwKigGfWsUC+yIwv3hnMBkMPP5PQy1ZG
a5r43hPBHoJc1hAetpkzj9PXQzcz6rcWnp5Rz/RzvzDxI7xX0US+bbzifw99bf0zWDZ2brz/3iQx
mAdbS7hA4yfloQlgT/27T3jSvZXKTagV2F9+s0TL6xHPrfZQolrVqFthKDXlV7n69GTkPh6vlMF0
QBz5niLDl4mf/1UpEdwqSRJ6eDSFN1q9jYEFJhmymkrD6jI3f0E+qk6RGhZAPzIW0kTvbm/X9R5U
gVsTxpK6FMmhVHH5lV9VHjRB+rW6vbqppnzI9/X+sXtXkTI8vIoe1inZfbtn7Z6vcqmndU1cUu76
oHCMb7UI825c3IuhOhkILM4WFL00tWP1/3ZAFD65jLII/zuY8KpMgwuOIxs8My/G6gxmbb1CKf0S
7C1f+mZOYNSLg8bDg9IORrnVVjpbwy4a1ELaxsGtgaPLPLGavg5WHqpVVIDNtiaYMbpf2LdvUmyp
QxTDo8B3+cO9p2hbCOOqWbRVtuXaU7l1ATbtAUAM2nEY4Ns584bMZ3uwBLxNiZ0koejN9gNEjOhi
f76n3/Wyql7h97iJ9Ci+ya79AVPWfmfYJ306GJ07yIFTS7lklbZg5enaDJybbt4iZzSkpKl3Jt3j
yty6mbUH3l3NiEEkpgwKVsj8HVMLSEhZMCG8e2tc0n7kluz3rB2gJe6Rq16OVBaqvYVZ57qiI+OW
/vNWYa6eWyEgFHvBOr/c9jl2Ju24+z9KeDS54e6EdYSrvYjcf/cB03BHbm5owXM2fdwXK0d6x08K
KH6/BrT3rdnjg7J4Dq7LCMRy4ZIJBucdp/KAG/FDPscZRH5Wf1Ox6/OtOzeMRMGfI4NGOoQSi1LC
r17XE95Zx/7C5A6vQmvixjpGw+XkcEZvw89QNq81Rg5xAA0tILPAmINJi79svixF+cGGuyOdV74z
5Th9t7SPAT3kU6Q7GAD2V1W6VA+f203p6wsOF8CGwkWXctutf+mXlTON+uulh7dIlrl55hioEtTd
HqDGnaBUiT10JP3mXU292V4cEgf+9uNlBO16EpojYMhsnv55LkwUWztR+ppl8FoF3BUQZUluk9Xf
FbatQ0D5bda9nD/zcNr/xujRMe47URYLsyih6HE2k1XWrnGPFiEJXIh+bxkfiTrKEn+lz4rwVgrR
u61gPjKkjUfwoZVrkDGL9ma1lXAobZf3CDdqKdgCu3dJqp+NKG7XFmrJrAfX/CCmsN9xf5DIwP7h
MlHegNVSX8ycqfNHtqCK1GJYAQEKqDMSprgoJ1+67ip89L0NAW5whN2xIsZeoEjyCzSshwf8TuvL
XHM5T7+VvPqjoIp0ZM7lMef3DgshmNlak09BhVCTuyU10BNKdK7R3s3r8AFWJuHMuuzLbi9crwpN
ccKUbQ9qdFoJnqfA7C12eRcyUUCCygCa8637LnuZv4Xd8L0FulfnPf81Eg40cZqUduXsBdu6gs3g
sSAX/Ri4Ui8EA87N6bmjSHnjSKdkT30a9NTLSGzmTLnTWKEDGLkLXPGlByoS9VpdfTOPvloglKji
phF6Bpgm+/dMqtkt6YC3VQdsheLCoOeBdA0y2GEyGWHNsCcZgdBlti7kxUeRweJuo57xkTjNSMFM
WRYjO6kp4VZnHxXxEVw68cjhe4teC14w2WFslIGugZTpxtXNFZAfrMvqHtnbSKpKOBTp7eki+Daa
AlX1kaMZDxGJBln2BWjXMBImMs8pYgRnv5mztOWaXLHQtja4RGvgzcJelzQWsdhDiWVHDo1QaqiS
RkXdlGUGvPCzZrsfFkHJR9aA1/elx8xlEVUXyEIBoiR8xpVX12QRL09aIc2CVHANUhxE6Tvv4iT7
PxfRuG91kL0h/hzSYgHYrRznBeWI6bNwY1lHzro5NzHG/+NB6DWAoXYyxSwHR+00W3AECSIO3Hzh
/n110btczYwrfgcImAQyRvd3e5INIlsEmP0xVNtP1Lnw9/S39e7B+OB3+IO8f0PJiBt0VPPjB2TG
LMpNc3r5B4qO7Am3yH899hh6E/iGjQIvcU+804d3KKNMATBCzf/BnAIBBEfdo1Eou+4ZQOU1b69T
WeG2fguL9/dZe5SdnzVWFpFoCeqKAlwtJ2dmhy2jAUHZQf9KjnXZfTu0kqFk89Mqg2owYwTNFAAK
sPixpHGIUZSWqnDkfptpNJcKAogx8+H2cIR2CjqEtONhSDyNBparwDarQkGlOvVYCXZH2kzO/3AS
EiLiN5895Lp/SFyJ+Q3qQJ9T0xurtNMCzysX61SGvWr6xUk2MaDJst5P6KXiwhA8UMWeq3f6sAn4
prsWcbvi++GzoR5kGIXNgpTv7hWmhdSQwxXOiC5uyjqBXXxv04ZKtqQpw51QCufMaLOFkUARlFFf
t5qc891N5KCntef7LK1lVN9vf6KgnTV+TDzX5RFTLrMqC4n7cF95dJ7NMa5F5qUCI+pYb2KusLbC
kK0clnmsmVMZvNh8H9LF0PkTR+zWpdszQDffFOgAzOkIw5eiN4nrRb+p+WCMlCDTwt8MB7qaAxCE
YGrhCE1qC2lYU5fjC9ujX5wYW1PBlM7mAg2YE3jLOmIUODz1lk5PDYYHjMLSqZUQ69cI/o7wnDE/
Exi9JC7GuHDdEZMEwSPUgLa8dAd0ojICCGYW1TkpyYgZB+R7IUxJSMLPCTCGOp2b42Yy+L4ZYL8+
rHn9XuSpM7kRSXKRAD+8DCG3WrRwY6p8bUPHomSblYwTEivoAF5gdiXnaJOMJtcdVMozP1pC9iHu
XclR9KAgvinUgUEROitZHw9jYXDYxJ8HIMF6z4Lg2dIMHKvo4dfo+CCaIW7TsF/sp+yQcz2UFOF3
JIdHptDUopva1mZFm57vetU0vAisuTp9qqeMPNI3OwARiHoBCiwfxMStLBTWfY7y/eSiPEPiCwt1
O9y9hdCjBSGujb/XRx9zPobqcRYxkS7rGRC8Kf5FqSud+0ZSza9bYzzJzTVCG6p4bNDGODs7VqIh
i8Opg7Pp++EOUgJwBawvnrtbjGmDW2E8TAbeyCwOj9xzcYod4yB0s0LbkBrqx/cAQE1MeHNJ3dMh
UG8gcshLzad0jX3cp5kQmaZrQARBZI6ZfLgY4vPntoKkDHDe3whsBDQ2VImiG2gJpVYa4Y7kcrX9
+32KUnyqeFvUSn778DT0lI4V2PGy6rOWY+WRxXKRxwAIpy9oPwhIvgdbV+GGOwS34Ke1N7il1VJw
3yYKZQZ7YAdYlEZzGaYeiwUCmdRiMBBe+egW14BPZp37IOdk59nO6XzU505W7TjKagyRtgm+mFSr
KAY1KyV/Ahp6EZUvUnUqqHFKK5BK5CifdAxFveGWJGlbPGL+DzvezLEQOhVXxO5EZO843IZTPCtL
1DHViTtmZo9lxZVJ0kPq+7DsS6awRp0WNw+w5SMJzfcz1bnHz4pEBJ7pqNV3T6kZ2dieDd0R2Z3R
CjeP7JrZemSOtPAw1EPYLCqb60t5BOxpZAOpaQ0jPZKkFXvv78rmSNNOh0lq7InyPvIeGDDt1VqM
7dv55a4+rioA5POUySWqqsw92KWg07/9i4jDP/nWdY6Ktf/BRcinJHSagPBSKV1UipkXp+MpyDPB
UD1k3vmNtpwtt9XN5Onswoo2KahqdNanAFoGn85FI+HDpxl9Ox2KzIH7MVhzVYsPqbCplMQWGZI0
uH3EjveZv2kKsfIrj/bdZED+jxw9iOOMlwkTV5ZVAhpRJAyMuXOTJt9NCPGwK4hZ+5fS0QP2q3FY
khqcY4pilDMBHP8QeSSUroTDuC8KCHMpoMbsdMk1YC+ySIOs+IHiZws5umkrq0AVZkyuSG+21g9d
XC4sJPlkOvFWzIrJ6Q3TcBBqQVYPkjjuZ3ZNXn7vI+4pZnB28Pe5wunPtX1+pRItcpJH69+JERPh
7Kiz/aud7Hw6XMzCLb5upwA8rfW5uqTxfRJqojHFgILlwBrXe/OZ3h0N3v+Mq3OGhhN1eiJY5WnZ
XiFdBC5qzFSnfyULW0L/U5+d0kiMv/ZsjeyOLkUEYfMzUy4NWWNaWTLz2eYM9rgzgKaGyrf04yww
Z5ahZrBA+p0wDVKU+QfieZFQI57PebNEPzqzPmrdy4c6euDYlPrU32sSYgiheHwJE8DR19MttzqZ
AeNrVvTU0m8tosOVH+PGF5y8Qp82ceGb0yrckjvmAWE9/S5TlTkWqPOYGuebxM3ZtWMfTffdSWgR
xX+lKnWhg/9dHZ8KEaQySuhrUgEswuc4d1uPoPo3Z8s8OFx9HPbL6w1Rspu70QZtfohz5Z5kdKnC
sSAUmUDdqbDwqggldxwlWzI26UEdG2H8Kqtajf9cHLc/u1xGpItL/reQCKG/OpkIQFoAGdvnlRgG
Cj9pPFPxhgBdIrDdY9a9fpf4IBlNUgVyLC6sVTZILsOcUbk98HsfhxOEFAHGbP0VIVrhjEukkHu9
qbYVMiSaDW99kxV0eXX8bHNxMgCMTb7L+oCJTVMsLljWpBOhx9OstbL1p2T7jVF34AGarUiJikvv
6F0i6V4xT8+YVBZaOUuwyoJuhybQoVjiKoD5SUbqkwmkgjc6f5Nacy6MFKtc4CTV3Qs8GOM/2Pju
vt4U0fU8QLe0xVwaSo984cf6EXUT9AUmt6HK1pPO02ZSEXHaaoemlyFdA/eLvCKh3KrYKHuSe0Qv
Nd/lJlevptnIH9UlgcOFcBts/JLnBLnGn1Mx5JIn1kMD7K7VH+nBvbELyvX+xJplJK9/dFjRTw8V
HnV+4erlc3ZQkiuvrHVyn0EltpDbPuFQPlEsQmOyhBCj7m8DZ4sme+vrwBrXOTymRhsLeDfjtM92
hB6vLlplcF2n7S1u9I8n4m0sceJN8UMtikCtx4eit/UED0VqwWjx6lIJ+EC1EgKXXFwzq5rujB6v
RiBULm+dUx+tdN/SF4Jh2BQm00dUApaTe3Bzfl8Jr+n7fR7/gSygyZwMfjLyTm8zmNOw6yaEIcmf
djZRb5q9UC4pO4aBS27Kw1vy8ZAImLkc5FFzbq9IqpvaMKO7Smlj/y0PprRCJ+/c1s4jh30hfZ+W
Ld1QPt4fiwjABLja5GV7Wm3BQKcfH5vwJRg0vJZcAI9t2NF2RnW+5j82wwnE9XvWvRAceZLYCTIM
9uGnC6eQJCJaAUTh1fDh0b5Pvm3PcCIZ7bCth2KPcKk0Mngne/QhT1aMq6VhS71nKu4McWQMZoeg
UmYcf6qpMGGo2J2vJka8giH14DNZNWEA5B8jSTh1RWDlndvPkmIGPnsOY/lyxaFxOVa2RQdRizLJ
0kdtF3Kk5+9moNsFGb/XREn2Z5kjHErY1CTbYdN53esk3XNOSxxnESKnz4EtZaE9bBniBIS+bo06
ug1k5ngFKH4HEiwpbfXLH/FjzA4obdxVrFnfD3yzmDYMseRnLrIxV6mU0R65InRMRT6EDXPbbX/D
K/b0rv2VKCX+dugvaUyFKsUQbMgWevTlMVFM+Yrcn10hdZwmBiF4J0/WqihWii7JulPfu20h3rnH
+DcA7LCfs2HfvX98v33NCCDZOBdbVHtzoOqHSGYaItkyIlJxHSTPijnJ08iNwNF3HHxg6FgTsFGj
nMcH6HHkzUdVpaETNfO98c7WMl7vcrRUJOOkn6Is5iQGUSrneANsB7wHq8ek3pGSo+3c/xBw21b2
xl+Zvxj6wKFvQk+93K4TT9sCxNCo/Z9orAnjyc0Ur10s764fTxfguGT2RpXoVltFVUjnPdqQjRN4
VDAq16YhoP2j2gTltzS9PfhPJMnaOKIMhPPOK40rxn5mWoonE935kg+M4abrO8F5F+TBxZZeXUpA
RgrIXEfYkIppMcwzJjJ236bPVqoXmQHHaq9QiQaPh1MwHqA/xgIGWdqIS8xIGqhca6++TMYVTNoA
+/z0/Iq2ful4DQSMePgpwnUraHJyyWxrwwW6wntXbOr+UJT6ieaTrRH8yRlv64niHcg5Jphx4IUh
Y55oBbNyzrqdDPfCIE3TMa6rhbnnnnAvDd2wnv8z17rBg6B6k15i0wXAjowuF5l6fYWAmRdX6p89
S3+hP5DwxvC/XTCPyVtbkRKrZROCvkV6UXCn50CJ0ZARJHk/Vb9HaKA/dZRdaNA/gpVwfYwp5i8e
IOtFxDhEWnNTPh8/wqRscos/kKf1p/IGsnowte37NTiiZ+t5rMr8bfyILSIDNoWBKDJgK7cXRBrR
/3TrTQFsJT2d27wR2D2N1ChrcXqfg4xcU/I/3GU0zkaqUVZWGCMm0WbiJGK9AaPWM2ZT6qPl9Y7l
UWgBsJOO8j4PfxL05S+G+wPpVUrWkjWk23s1cO0WJTHOST1acn9Zb4cJm4ZvvlL4WJWmD97sM1FP
g3XSyDil7Q7bqbEtzvI2M7fMlObJd132di5q8BHnAldlVboYzLYzrlQOOWKsP55+Cy9KMIqgd6Jd
bWopP6hUMop7VlpjVhWG+hDaAvXWB7KrCmNSfkAgMSM8kAW/iRLurbwEQbBOybflx/IinyNYqlmr
KuVwaGJ9o8AOf8R3/27qh4qCQfD6MUGbjukoku238sqlrp5FVKqkLWpmw7zMMmu/lKY7gR0yB6Ro
aVEyr2EMoKexip9kadLOsH/RTtzoxQwP0ivbUwUbSo0P8BnsXTErUxgXckfstM4t9LbLfIeG8J34
2CCQW2SeWJuLFx/KutI0v7xfxxrGgobwqTpRZ44IRvoEnzFarxncI1Jj7zcMlfwokr8q2oU23mYk
6sXTCWlVTOiSYKy9Zu3xzWL5EatFaiy+xnui6+R9FskkfgwjcJuEib+h02z/69Gpork7vkFgmzfx
Ir4mK+sv00INm2wX01cgQDu47b2wnFqmx9v6hu1XFEQQYhtoPVYYzRpL8BE/qzH7p9BxKlCyi/9+
8HxjwOAmt5VYsoXVNcMo1LDG6VInRg0pwe1dojk7VHfNf1KXLUhrkv0/huj0uxrdD+QSGMubwn1+
/vpkwqgSDmZ9V9hwi2UhRlkH/vjoho/Pnm+13xGPRpE4WnWFxAVyg/4kCkXzkXAVVyATm/FRD0fb
Ve79T6iLOgO9K2aCqMZIBQ6XSuuaDQD1XjX7jpDX0r5TuXsn+w7VYKxGUlxjZnrH8+e0BYo6kzqK
wByEn8Lh461eW2XTvSXn5/mFrnhJ7uvl2x45MquWwwBGKyvOBrR4cC8aoVqknivgWe3wPpPFiBN+
nFqyZOlGkBOFdrfXdoG3yQaI7hD7odNICeU9vY3hmCbNdPKl+lpQcIZzpkC1PeTjN4nF4vVpe85H
x8xNnetY6hOpSBtP1NNV+xQqIzJUKKJ57+UxTVFU9JMTSSv6GaB15SLnY4XTtPnsl3ukWJjOJa6o
KDp29OAPd2cSLI+aOiC33Gsm6e7+MyomlMf2jI1nGjWprvc4XM+MGXlxeeX6I+qZ7BGFJbaNf7ka
iJaMtIigr+GWo1PegKPTFO4NB02v410kOXuT9WCvQ/VKt+6Sg/U94PTPydFDsifHQ2RE4UEmWTmM
1jow3MVO/svJSmJtIDEK7NWk6BY9rru1cRn4EYRGefNM4dxM8TuP6sBhGhoELvuerjGlJCPz2Abe
Ky28GnHEzTGG3QzN7pNJGwz+OieXhY10EIkCARte70SUpCmMWuolxFcEbmfzhOJyWEAX19SxpOou
FJDeB2AoUt8Am4XWlLKaBwwDdOs49cEHkf/cddmvgCHKST/f3pxcBCk4Q9/4OEKv/Jqy+1i2GxRi
kH7zBZFpIpFjiLiELUWEVXKIP6CvxDcvNa/O/4fbKeuiD4lJpuFfX/7GBG/ACYC3E4RPzE0by3JZ
niY92CKVw+3PUUcYAlxT8yWjFSGDidGNMB1HCOHoKDO5+A4zqCSq8FFI1u0MQZXZv3XumvNYEUdg
9ddjPrXlWBrlRPwkigRDw8nQ5bDn9FvLNCsTaausY3Dl4xV++dTMOCgxUy/4BSjxLiCUaT5Cq4hA
uUAZM3FGGTj6bH+PQpHB0CJ+wnvkXieNGzOihLWPRRm7qhQ9i4zT+JpClwpSibzQng6KVaBOnqPp
zYgUxHtwNpMLSM6px7PLGbyN5wLgbCZzlKxkpcMTgvgKy+kn2eis96pLEMyPr9Rl/T0NaR43N+UA
+xG4kUNgRrfQ38fWUAN9cBFY3T4ix7uo5HeJp4966GSITuH39tuwi51Ga89jv8a0zMOZk42/ZdAi
RHlsGuirk4Xg4kybxv3Woxp8kGkrSB5Sz9OG1CVpobPLjZiiQeDmFUw44mgkCthxxDdjiu7s73VQ
u0Bno+Q1AIfS+UYOW59gUyS1NHDp/bGzL0D8/iEjk58c0xv6BBif8FRm0szeUazoMVWL9ljnryWd
k7/tzV4s/kDEkWfLAVH+d3ryor1WEvPO7TZi3jUY8C97tNhdqQvP0IS6WnD90u3JRgLnQd2beGX5
TZgbgamLc2puHeSIbJRqcwF+lw1FiqFXHybsdH6r2jyhQBN3MvNyxSgktjVl+uEi3In00ep+HmqP
aJ1pFkC1TmDzNvZ4mIi4I2aAbSb2gNPIIaE/zVL7tuX+pdHw5cKl5qiWFcYfmYuoo3mUV3LwkY5r
UbZ81bwk0yyyWjzkV7OhdiGztvgTYXt0VSQhGv6V4lAq4slb2LA7d+Lnk3AxLTG8IKRSVAWs/Dg2
3V9deZO+udpt+RQGIiOIb71bZz0rwytqozEoiG4LOLIAFo0TtLdKz/k4GQtHd/DS5Lf7zFzfrZwF
vxAw6MnHCoKojDGBhD9TcUhvVPfRXOhIJeH/VhPOKuG0MawxWPNKF5emeTSd/94PS99xPEws8blb
kqgXzGPmOY9Ycjx9sJhr9oLPIhBMS5kXAjRaw9iEUu6dnvC3sbDam3pBPgO6Ck9jUQg+TKOsiqou
Ecgw6emZ83gLIc+rUb9t48OxbvKLH+k2TVmbMGEa0jd7u+gSAzjZNQI3dzwUN8YmVR4cAk1j3krZ
/z669/5WKH3wyak5rMPM56eB7jhxcHbW24yuFTaMZIySRcu9HMJsX7mIiaDTaZtLUBy1iDn07J+Q
YCIAFjJIdL+9XQlS73C4qmHNsajZ/rvB/kaj3GRSinEDw9Pu7p1sTXDbHMjLGwq3DeSZoIQhKYWh
ndPAxPSxtIEYwc0Uz8RtHZTc0ByKlD2oahU1rvLkLD4fvW9zUgTvnadiFrKPKPmG2Uz/rdhcldY3
Re2Ayp6PgSsDYBtHwDYwkVozcvRa6qzQA1IU08P/PPl2CiPk4QHwQcWNZElfpYc/CTJ9S5VwKifA
v1ohBr76dvNxFyBIOR3jXvAKV9D0veAyb8EUTy4YSrVem8piRbipCX8AnJzQUiFzaarbZ5v7eY13
hyxIszA0bYIh80l71Cjmg+3WOib4xmeePnxqwO+iUyfwFBgHXfZeewSJbVHGuLX/rGuxC1y9d4nq
cnXf6GUPx6lGwUo+Nl3Fo8zhSLOStlpiT3V+J9LWpicVEfZaEJmF1T2RiWq0B8LP3DY2dai901Y/
fM6WP6gY+bH068KCEyOpmnQEtg3wmCl9hy+ft0Zm/vE+59ZaIzsd+f/a4pwHVIgD7fMldLzClLn9
jcKsz+STAb9u4LN1PNy6Jr5PNBo8Vf2EXuTlYz11ifJeKESICmBWVY+Gw71VQT09PDcbIp2Cdl+I
xXpR+ywfvgEk0+1+K/ztHTVb5dlFX3mettQ2rdrHSBd1sYbcPBPFJ45N5MgBAOqUUlLGje3ZJkTn
SJFC7IZYAJK7g8IyUZ6l/VzrmjdU+J6abECb1NJYTPXBoBUW0DyCmpBSjhOpcSyz4/p4URdnTbRy
GeqsqbevZCXIoYDU88JnTuFzFr8sjk9VT5u8NMNwPmNzBz5VTv2ZhGkeGag0xRZ+pwjbbQG3CTDJ
Jjf57gOWRwEGVYJ4eXOGTVMsZQCoycdi+G6ZHUYRhhcXDLDY/xY2iOH1wq7OTncZP8soV8duDKrD
V/LE5HfSbD556dqO9DXQ3LuotZKCn1UmuM1iUbe6jhQgxGb77UR8kTdpwJ9DkTYoKp7//0MXVuYe
J0R9R8VMPyO+1yCvuB8rx32jt+qplJmP6yhgRRfAA2eFScmAi1LIEwwcmznTWit394GJwPWqfwKU
IhFiVcOPIxem7WFNocACKBFdYryLjgo+gEnPBwKi91/o1fIxD+HRkBJhVvly6XpJ4GR4A/X+qMuS
iU/0BOQKPsVJGfOlx9SZ895BV1Hppq1GwnoKV0gC7geNKZsLToQbArEKTIFv5df4IEz9Xl0bZK5s
bF+xbTcTviWCsZkG3ql5JNC1JFaS7VJ4nG5RG/wU4SULvRMNOQpO2/8B0ZkVKibbmn3NB3DYt9YV
9QBwTwOQrYQ1B/4+Ps9AT1Wyj3F8t0ElCttVzETXBeOUsFT/MYkDEpsh0njQEVp2NVcxoU3+fNpJ
mdo69IRq4IMVtLa3HaVu2anzMzbmZZyWUOsT/EB0Yy9HMscNALRxJ/nyrUG0TQEDi9aoYUC7DVXY
ka5qY6wkvQOFYQp6pRusTR6Nm1oJdIeLIp2ih/8OpK00K8afMatXpL5hkETJ1DxyvEOeOcQoDrx8
7CdeP08xBzEJatBwz0ZordpT1dMp4AIqgrTK2bD2ZPBu/0/W/RXcy+cjvioIzvX9OlShO/cZd4EZ
BQhRa13Mmh2tjERSYlwt+Iho0jakd3p/h8OQgrhD4htx0gct2Snq9z6ntfXbWNDROOKYVr06JBAl
gamM16sw4zxa6OzEPHiPDC5u40vch6NmBuAzuiQb+wemKAGmxSSTFAmCMDDUagRvYlKzBd+wFVxk
gWFtidSFmOVEMvrSTHJ0z0WjQejmWvPVLzXdm6evEmjmIMuFAleQXOKhgJcK/NaJaP9+yxVQU2Ns
xD2YOeRWnjmINMLz5FyUYuY/0sZ6k3ruxiMchhGXVRHjl44usVXIUFKzVJ9Q2yrcw0++2H0SMrx7
qbMN5YWvPGQxHXyx5kuZrx/4f3dvcW9Trj0c3Uvu/EMjgDAXJ8WnjpHaEqSrEenerHUXut+GWi6e
zz/n7eV7WufAYE7N6nBthmJ+LOUqI+IWBZwdqC+V2r3BbO2J4JUB15v4V4HfQ6hrGb7/wxf928in
t2MtI6J97VLlmFrjKxEmLtXjZDZ0zLVnvThGptl8Tf4OIzcMTItvDv5zdEW6RFTm/YZC20fF3uLM
m/i+JLDO+icBk08O5aidVFAmJMIrw/R241Vrbc+zabyVYqTH9DlYEcUMV+sInvq+VM0LZmKv332j
iuuqmGR5Z2eSmd+7tHZsYMPP7fZ8dfEWOBxQ48nOOCEUsMZyyEmlrGUJf1wYqusfb0HKFMPsyzwY
qQSGWw7NdBtzAPrP2V45QLmLXYPJUJVsU8TbmiB11+fMlRH0RHBEIOiPMp2eA8fVtYqYT7E4KAUs
QrjkmZlvHASu8N5tYjBLx5UbQPgq01YgXjmuBdOplchITKhmV4tF3x+p2HllMhtiBMGRJsM0phcl
pbmPs9py9jjbyDCDsb9xaNRsj7FiDVSl3jYHn4k6MQYUwJ0h9iXFOP8F/LR0BSf5V6DFU7aMV8hW
oCFpAHa3rpRIpZ3bX4QGhREDb/gjy66btS8O4sk/0asAa80lA2F1qBFUImNT6wQA6bEmOz6rQ+Kx
X59M3GH7+IRbh/TIjLahsjHNni+4PwTka5yVrEyOl0Xh3rIZVQ/+/W4Ijxz5L4jjCBBuvVFH7f2L
7AF1dwzH3DcIaupshrKqGk9daxnCPMMRrW6lxKUiUWSZRPRS3LTrzH+d0r/dn534VkeDq7R2F79W
JdxsABhIK64NoPp7+RgCW3VN9bQODDxRAKByOCeog8G0cZvBpoTYwCtyLXbQcyFWIcnwS3Jdw8WZ
9wMlfc+uXr+4vXvVIJo1bcDjQOJ4YHPrwJ/taC1iN5fk35mm5OCoIT4vAXVL5RfDGxvxBbBBwh/8
s/Oe8V4qQJGRESEfzT10VEWJf/PVCzvWJ0BDxg8VgDqWsucTjNhIZLsJ4VjTV4iDxTjAMEkXWDB0
CCNwMh/Gcq1Mz9bgmim57CBR03Av4GagtEhntIzEqgGcExt+GyR49wPNoS6nokwNXkzAHPr+0eT0
ykJGFv2/lj+5+tg6znI0E6dIbRRMLpy+Qj0U/hvuKZcX2yZBfGk7n1gksEZ0FXeRp9YbhQtMujqt
ZW0NbZQ1bfxUcpikCzpcZnxibdoNq6dLu5B0/mgqrjxMtxmildMXCKIOlKRGNns4BkGA7sCQynm9
4W3N3ssw+dy5whWi+h4GWuF386kPbdLnzvptCJbZG1TNMJJh+bC+ul4OpKBsQtKYnBrdNKodHbBB
qIOPjGuf3jt2RzRWP5QfDCUit5aIYCT11WfFEABr+4+zpWMuZPl9OVuoho2asgtmhjSj+jJbAlvJ
XhmNSunfD7anOupZjNfb5Jrhg8gwFGjU9FR1wX1xwFfqGC0IyHzVwC0kCdXaXZcxRbiqkPRfijvm
0goTJ9So5GexpEqrr34VrT3HTTf4OYNGRXnD7LlZRhONI/oJZIj72cp+klOYQFpkQGqFS99rdVnU
V9F+SC2wsCmCwxy/5f0tuHNzrnmYV+Ej5QpSRiVZUcWVBLoZhhfx1Og2VYH0lPJC3iBlAfLcQ+23
GBCBx5lAqS+/aI4mBM1ZsD/oreKgdR2EaU3KHGkbQB1AQ47/hSEmOteBTiIzIbMuednDgeZeBKbu
vkD2JNPGAwU4D93juuBISB/w5OeXH64Tpy/z7Xuia7M/jNpTEXwkO5YWrJsvO2Y6ryegCuhsOn/v
JpcU489WY6gLz52djEHjHL8dtu5+LUqblRTWS6Pfcnej15EiGBNwtK4wtfxz9z47iGdeOhd3iXPN
Feq6XWywxf0xSw+Pb0fQkSDiywzl1ssDUnIZDjT2NjWHdXZYd01t61TQ14uoIqz96IKqaBc6hjo0
aVxn0G/FOW1N9jpSFPr/OdeBhGfOdzWx8a/duv6bwvlviQY/Ch2MeGpdS01qOLxI0keR0+32r8Za
cHIABGHdhrXW7ofeKcdLyNg71kFS317aNWjCILUkfQKqwIlwvDURRwxWVeTyTbjGA7UaKAuw7GPW
gzFLvThZ/gFC5xvkrx88ZxqrfHDSY0gDlCIVVttKJLYgCrgQPucmXPgS1TuA7iF9MSORSFiB/BAp
j0CDmijzpL5J02FaXl2TJGeFUQ0YQuYxk4GN9FnVO10oWAHZzDDo9ss9Pr6qRCyQqPeBoGEQsZnb
6uV17YC+vO8juuWpfKxvsbpn3hntSfS64JpI6F83TqlI12/1n3Pwp9SYK63WyTzqNrIiUoH9bsIz
GpK3Jr8Wbp1n10wG5rf5cKfeslE2xYPASA4U57aVK/mKZvP9pjqH4iWdAf9lLPLH89qTTgLuiHpk
oSIjY2CeuVr9n8bep3yi5AhE2AvDAUjtjQXL/chHpEuRAIRuGUt7Ao2BwhJr9glCiHhA3N4o6LEQ
vnwK4XBDKJhx//Y5U40b5AX59CotefeDIQxRclHJPo8wqqtXd9vVpxejIQFAJXHoo1WJYrd5t2B9
1cYroc9wZ1nyjl7evFoAcZeyk4QRz454EZ9C3Bvc15E3Fp4Hu7Y9Ue6MbkMo0FKg7fkkW67HJiw4
HvyLm2G8NVYfPvkgI/oTsC597KEE3qoKBOMwoLrRqMBFxR8eh/HXJ/ZYSCX2jD+cb08GbQHEF9rS
P1yPDXjIdhQoYEC7o7c1c7yfITlLO6BfbqW+yWMBRsZzrhZQXTY0i4wrfJGlDHUfJk1hycJ4uGKm
SfdA4o8o3ClevrTumpzA77iFrJEkuP7MjeifVwi+Xt2mZjXYRjl2cZK5fDKLxhPi1vhpanj70y1S
tt/TkYAyrh6LZGSVi6rKdpi+wCLfmR6UDW7BTP63n8rVdaM3yTNT2sRlXy4a55t1qVouyjF6glJf
Z963lRQBA2ghPCxMWp9eaAveby3DFTNzdXDeDOW7aE5fUpgw6PL7op3uCCe5gNNgG6rdJbUKCfIQ
KzJGQEw7WtGGVoryr/sdx0rxgSL09Wb2jLEXw2131Is9Jhfp4f2bQBHNvNnjuT1pevA0FLCW1W7D
jr8Cnh/l+K55aSz8lMPeYvpgkUVF5O/VGODA5Q1qgdtt4iIRDHScnKdY9b8nfVZVJxJboVADkR1J
jiMGMU9IAyRIBujqswCdpW1aLwJlo8nfENV7Oy8xduuXy976nVEQUlrNabfkFWPp5nFBOmKippSr
eZlZJUNhkhLyhfmLoWwM3beGtg+o2qER6MpozRrzWWa8gN7+oBhB9bDdcXeYO/Ltvfp46QpmhGgj
GrIeSiugYSJ8MQqfvD+4BBXo40eZiOkrsA1iETh9SoDMqn2iQ7HgpNoMBQi5hP+6esA0WmLlkYg1
8zXNBmqYxz260ZFEgiQP7lL1TkeiWpWa8bx5MptyzXb0vU2Zr8HLf2WWbHzfCluOZDTljlejIKij
irazSY0hTcHOQDC1SZSxN0V3NA3/yhKH5wK1cskYUYZBcJHfCObH8Sm+fNdIorQAuDJcawsGZYN5
vDE5scTgugk3PWOBkOQZrrVS4F3VS/SNxwfOgRy1tJiLhLjf5fLjW+xVmjty00c8dpUiaZBPOd6e
KboTm7bU0Nnh531YZliBv1GpLwsd94lKE9RgMtTPQ927p1zhtvZPlXNT2wgROdppLaQfwTGZ81dL
foltGFpLcCT6w8WxtTb0Rm7OrYtZHqCJ67eG2Xt8lwh+k+mtE4k0EfA93FxDYlgiCUImbP/SBD7c
jTfuafg0L5EXGBbZChc9bKZ+gqV1kCcaHQl2NFdhvBmeSB97K24wZH261+Abc17JkKNiuWXLuVF9
YwfZRJ1i17qusjdi8IUs7HL1vRZB8WBEZNzK0ynfTleRootyMS3fkZ1QJPBA0IwttSAkt1nBIrVL
p5NGvcWOKtY+dPYiR7i6Jt/Jn0tbuaC/U18MA9FZZ4gATKhFGDtQXvgijpRmN+R/RjJxvEdvIfIx
CqrvPLNUC9CQoOQoGsKHoiLZfowIrcUN0yKX9MSbP5WvhmGIw8rmMqbT0fZz2t8NgBGudrvZKMOP
yc9HzmYLpcTrMbCK1HEPpHn4q73ESTRI+er+Vkx0yvCOaa362a7JerKTWWRaJneqGKwm6cWdZAoa
M9M77tQ40ZAghPjiz6SJuAXO4zMGEu0snwylLfMy85w5gCQnrATbArKTZd6K/+RRtKRBMeglBdaj
mPL0jm3924MGo7ZDp3YKO1KY9PyUzwgzJtrIIYygPwid3kcteVsEMyn74nKWfAfS1Pa96jDzhysu
TPpc1bWrWeLp+BI+Dgdukyxx6pGAaj8dh+edTcFCxhAFWr9UsT80uK2aHeJj7JHufp9jZNgLH7N0
4t4TxT7Dc//y2mP2oE8QZGTXux27qsEB5Vm8PKXfr7Jo0o4Hrhqn8MyndPiWpNjTn6foAOiV4338
9xe0V+X01lYel12edTxDTQGRbghmqIftPU669DukYN/epO9yP6MtX3zX2LXHo9Po5guwI33937fo
Vqjkyop2wX4eNgKgDAKk82EkdbxfzSnRbDXS2TigezXgc2JZnvzbmwM1lqBYq3SOQ1i62rWvwO2R
FE+OhW+JTrDa9kxt+mZY5HhBX9aiZ7L33FEO4SHVXxg+1OI8HwCh8dharb6ParGnAalx7HXCZTBm
RDMFgZyUDBotW7Rq1ghNWVEcawASJuuFgMcxzckfYdpwNx6bOPxwuQHCZwnz0/CBWLxgKvj2mkW7
EY25DUOaBHQ4sC8NOTZvpV+oOo3nWFEzxYPghA9Z0umd6VcTc+TnxHXh69o/PMt8HcVUGbHCixb6
4ipeVfpyGqz7HAWW+ju6OIaXgo2Q/Zx1z6qvVFX+Ml4goJA/lTMRqvrwOYlz26DKwdm4RCo5fCBv
I46pFwwj0+wWKuVVLp4oHQtwXNnQ+OED43AueaIqTGNITVJw6eLzCsAVNrQ7kNO9foXdXPo9K4I2
ijcnGf/wxPirSFbZOxTvS7aybZes/HAYyDpFWpyCb33s7CEocUk587ADT6VAHKAtFVaRHzZ5N4zF
WdZgHKPwmw5mTuD0Tdh/iBK44C0c43r3KgB9XLRqS5zzOSQHQioCkhfEjohxBb6717+MqBIuiQvp
MEwRqgU2Za6mtyfeUpyWy6TiPqFJiUDXEbJfNkSS58nPS8anZwHGUM9n0byf8WidWvyuPeSA+8NP
wL8HKUajxD8TQKDcj9I5s+0gk4Bh5gttueSm4T+jXpyuZ+tFy1wa7bYCFeKubP3d5vcYv//q/82K
apROUeMwKFLYt2rcVBdyCxupnWiu7Xub3tYslAlOZ8hNEfPxOXKJKsVYSiupkphYyWkxhaaFAeGB
pJe2Kg9cm76o3vf7royCmkCHxjJEv2Ha5WJQYiUmzoQAuXHVnGOUrfFAwtP/JVBmsI14yj/pV7i+
QrIr8cNr7LwnO2md1Y2WNLM6TupCZXe0hAOmsQguyaHykklJszmTETM+9n3l0OhJs0iA1+Z+lzwG
MBq9DocgLmhrlqWdIxjIwtQupTz5kqz2z1OO59N7bxD+cD208BtU9NgcjfwiolnHbMkQhkCKYFAm
BGV0AbebOq94OENYlYiXU1oZQ/BwwspOblJgneDiKxjiceJ6nrFHGvNauMLCU1kKqlXbnuintmKy
qUCi8KcKyQcPHrQ59sWSHYEGnkpp4C8U2zVykOWuG9iMmIn1nvBI13sikD/JVaa4tsJYQH2fo4z2
9LUe/XcGp1AwYwQ/mzEiLGYIl0KKBKayXsBH7Y97acVolh8MJnjV2zIqa19sEB0JBgfDkeg3pZg5
nsAMe9WHRUshLO3UNld3rmLQav07zIskJguvv+WiSWGhHcG3lAm+A/P+NSYP7Z/MN9h6roW4eLqB
dtyQMfOWekML8usNZltG0vvmIoX7PCR2JQTm1MenTQw5w+UaTLOWCdSSrYLOFOCfEfkxdyGl5pxK
FQON5Jl+lkBWMacw52eZ8nbPZC2pRcszcaDRDqQmvmJoM2CgDEIwO5dXnghp9shbenz5Ui/vo+7b
EBp7Uf/BpN2lk8sPuELPgv38oCw/cpuo+U3e5/B4upGvYtG4SRgrg8zXKQpj0E97iVpos/ygEN4z
Cl/xZojlpGKI0Fd3DeG0VwWF1LKhq5xUBJ4DyNPGnu0LzJxFGsE9zUGSBy5gGIOSRBC1mPpROSlm
E3AkUYq74hh9ZcF7QwPZOoJtw5ZvMyTMl7Sx27Z7F/D3yuP6NIq9Mp4G61eU/+ZEGWO19+5NJ2f6
Q2cOpkNWk1SKzW9iliMi4eCKs+mUK+Y7aKLWlLjzAcnhZ3w+NjsKEQEHI9wuHnZhKjyf9kZ7ZWV2
nBSewAGADw6XMLRYvGmrwUICaoBfRQcpx/0GOZE1SdQ/jMZLslfOzcWiZ3UmtST1olQ992rT9TJA
FgLbxWDWfUE2TgvAQ0Av30xzfyNEep9i8N42gH+0JvwH48Vk7Ckxw2AoZwQM+hPpKTwLn2aHfMGz
/XDUG8lFjHVT0+tzG1VzENJGUwb/X36DPs3DpF20RwmBbgBZ5IJ8QGDUANOGv5UWdoV+k8TiDaTs
NYV+xlHasAPoPbvlSdfqyD/0ZdBLbtMsyM8x1GC+zexkJ4FNIAWtEqKHMG8P7y3CRIMkY6+vi4BD
AxXCIvO59nSQ2srEpQYGJzyVMh+MYighcQjL5CdctGsJpes/xgbs36hr0To189IqmXRNbXaaYKda
YMcfN/SNoax2A/4/dfbsyyD4Tw3uTSns1BjKZPrOCSv115YrQSTUFc5G8TYdEZt4QJCGHjg4Ym3H
kLOJcUe9M0VU/Il5zVkPhULVTXFK79UcTDZXFYQYN2O6T6CgwxZgHU/Yq1+xzG7Op2sf+2cPsZNA
39FF7b2b/K19P2tjT5Yh73Y0+FGSii+20QfTJs3WCN588PFnHE++6UklaKlRT5We/ojluFqwTcRa
NPPxEKfKp00p/42so6Qlx5NQifTdt4h8CdL8w+GpcENlgvEmn5lGZ+Zj79Pq93xlHq6DwmTuJTbY
qdTajIYWyQ6KbVMGHMm6pgvXoPBCsdP3KReFSDcwZE2TYcnf7BtAYhf53kwMjfqfPNSZ859zHgiX
ZDU+L05ZRafiWThpBeyVefQWBGtHZgVsihQD2y8lJjFBqU1SVCdKnSAKTCRSVyhEUDHkp45gnTT3
3SZJbfnp1TTjRZSSEU6Q5q9XWSsFMzi35XcnKGA/plzmLKwLorfQ6aByu84U6I6Bx/Buk8mC5I+6
0HPXsjHd7t/OUDO1SoYMeE48OCdY/5CyRylYMjsPFThJjlJu9LunNfxUz4CrjQiKhU3CRBXMFOkr
3msZnFqrh7UJVgWbLvx1iSYcBTHgh1JEFPRXx18MR1UpeWM3djVws95mjchQoRtmWfybmVdYtFPm
jMd/eHYMLyL7W6hEzefH0d8s+f+K1NYAwC82zUtfZaBcgvnJ6NwUvR6iOFPAmdVKQMjyZtKuRioT
SzsI9ytWsfAxTjWgd/pV4USUBU3A03SeqQyCi0+inV1Vp8AYHlQg7KjMRoZ/iITXQvkbAYVh11Ku
5lRnjJLyx9+BnUSTjrhyxhZ+7m/TR7aLVJi8sdYTedlE4j+GFxuKDg8q/OcHX7hh2CzOvSafOAzA
qnZ3uvv8nXOcWMVLS9TvIuNbhq7sVHfSS1GAsn3DAxEbWXT9bGS1rR2q7HTjcwch9JGhDm6w/sKl
YA9W/wrd0fzZnCssN3FdoKQCE+2/Y+9JAClt5VV43TKvO16Ngp79a1h82WhEuV+HCEkj/DsXhcsv
TL2Qkxw3QEFitlH2goUcDDjSACOtBq2RZ5wrydDicDmNHPSY/oplE6Z+PWl4J+dJt5+57vpQ4eWO
nynkKiNxc3Kb6miMeVt/XA+4ZxsCGPIQMmhd+L58D/1jcqiuvjcBZG7NcE0R4QEEL7h5NokhcRYO
q+2U1uT7vgbBiTZ06w8y3NL4cEb9CTvSKt873nGb5FNc2Fb964UQM9slQEcLnUoCRsIVrD4KhOHY
cDwBA6V+MDHRN4YklVUdReGLuNigUJ95U/ZrbIS/GWlWKexokftstfF5ueof2axKNkhB0pjpu6LQ
H1781sXscay5szXEti/QgTg+5GjrmDVdE7n/V3cS6w1RWjuXG7AZnQ4JtKD/Ssbmho6c9nsfT7AC
x4kgSnu8PiqRpi5QCHZkzcgFpEjc5AgmY7kKmgYKBxFVDQnZI/v9fO+erUgyw3XEm+TsvfVwIUAO
6tgVWvN4dNxd4vsFWl6u1cvrhn7QcYsOCmri4OCk2pRC/2bqhSVvpemDEVKdrNfqQL679fdu86E1
WeKGzBJERMqP2m4ZjVCY2VQeHsNm6kl7eXYGmjmxpiV2AfgNALolpAbs+wnici8gh+4LALL9Vk4y
uxssqICL8lVPNDLP1D5T6XFIL6GaIg9D9SBRiQOAhbxYJQEArJWWsXMhYDuTZayf4lLYljbfaLgv
LnC6NDTEY+l78LK6+fJ7A0OxruD8cBjbP7c9jS4W1daVwYXSybM+Ue20p70g35uvLgEhWYFC2W4L
2s7GiP1/n8S9HhC2Iyhh9o2L72nXKvrThw32z9w8ZjqoHgPP2OAt2emnry9jDtT/znWpjoqXVtCD
qZzQMhq8fm4Sux6tlRJ83tXDz3PcybzG0WcHTqDSEvUy15ym+pYKwNxdkIcxgPmsBEI2fYBZd3wz
n90fOOoEZJYcSQy1+LCtTRhDFLW/Wt8/NGoiJVI+QkK8apNhESoL8Ru319fTIkgT/4LNeKQD8S6d
0wkTEsGvTNZ9xPSgwjHz4z4hydxK8sZtd5BcAAQyj62xilwmZhZZ5fkY4CJqbdJVAOO405E8Ba3x
KuqT4ZU2vvukNY0Mee8q5GbXgHP29jNvfUfAp0U6LTzSfcpkX7XFmdlj6/EukxJwIu7geM8/cP2N
1gFxZ8j4UM5/i2s3oRJYCLDKnq9if6N6CPAKeTw1Y5Fb0t5/QMG/q3NJNHcBxl5heK4Neskd5x2J
3M0QtwqMP8YnaKNFO091Lo26MkymJxj90ZUxbekn4D7Pqw1O57mtLkrD3iwmCJzGduyAeYszJaX/
CINIda/uSeGVAoX4UihHh07GG7E/hgTGZIFNM4dOPmMNGir+MTu1q8Mvy/4trCCYuWKhcPnHBdQi
rWd/yIsI2i6rOrCpbT0MRgqBTLvtzIaEIwUlt1iaStxu2DI7SIW1aVPAa3SYT067kkbn/gC2Bt4B
f8It5WcfaoG1KHQQawTO3eZMqQeMEB+PcnO96mqnl9YouO/Q7aK8LMJ99LJNJ2QGnRRtjw1bYPde
ErdoJQhps9eMvnpF3xuphncSO0wI8JaUZey5YBK8rAHlLXWmGAQGmcxXKjwnIt3apDC+6q5hrDbE
iSUZUvf5Jk3MgHiY1v2pq8cQ468wItVrtt8Y9RXyQnYdRpSwKkRypArgjI9KAMSnhGSXMKUSboFv
V6Oi9nuW0DQXQPt9BM4Bu1jwL8mTzkWI2W0XZt32B4tLePJqTVpq130PBobvtUhroPWHMdzEmDvG
hK15MY9xVeMokrbZgwkZqiwjXsn9cRyTgKlfZ+uaJUWoFLt5O8iHg1vl8OfqJ8kWbU3cs55DejdV
iVqx1HDb7X8w3lkVVO2ZxCFHEIE5nu+iapJjpci4WAY0f/IozEUFWGxJkd2pu+8NJOd7af+JfA18
HxLXrkNRbmr0Rts/nU9A0XhsSIv5Lh3yB/Ew8Icq7lDWmvWHhIK6FuOp4ODrnAl5lkBiCjqTkQUb
ZoRxP5bP13khI3birpYoKGyl3l0Mp0gcngfDJgKDlkjyTgSjc3LOPF1T/V8UqmqAeYLhNvPzND0o
BF+75Ai85Eqw3GFJEap5kAi4e/Iny/l/aVwCIstRpDcaUh2dMXDBuCovVhswat7tfnT8NmXfOFZz
jNOc3CXux6D1zJZtanHUekP+zGrgHnZp7fTE8h7oKrs+roKYILTY68I43kk2hNpSeSHUByXxIHeA
TFkBUUe4gI+UOaxOnvL4TVdZ+FVJXVG1+x5vOYT35CdRTbRI/UpWerVmvlcfNmW2DlihlEd82UAJ
M6eX594xmJ92NpX84diJE3FgnztwiphExKyUIoSVhq5zlv07FvLWEX86xOxvhOm6y6GoMCHD7Dt1
Iy29CDOF5INq5sO0JT2iKWDmhNl88YaPm1xG9WuE0qyI049K8g0RI3pDQtKdTGL5IyACtyhu2J6o
cLsIne+sqlJ3VB00PF/PFo6jZxgAy+5qZVmW5b7UW96SBT64i1h6Qt1XyXeTxdR7Z8pPcNLxRqqZ
y1i3ztwFhvnQvdV9yXt7mW/dyBP1GpsrShPE84gvZaO04mtJyRNfuiHPjyVhhMhAqKmIJq6skpww
VfvHk2GUH0JwK5yTUTcLXepUuau/TOJGKlB/p/mwYfDWsWuJ+hVhYgnao7HLrLVUpd2/YS0IurSA
lDJ8kHzKVEsujIOHXIMt6NDx+lurVL4E//GRr9O/GFesxNQwG/4pTdb32uw2PuaNzEfvq+LwTJG+
Q9YtRCS4nA88Z4kGNpU8SBcJBFSbUKioGqDSjqBoRNtUi6J3p3RWjCAW/7UrQjozTNo/gONJAPJH
TNGhaHhtJcXoHChEPEWV7J8IkkheYUVuLofytw+UGwZoEQFosu/kXXPptrQSZgJZgIeBIyBCgJbK
97TXhCend2UVqEPgyX3fB8C2Q8j8FzUT0171uMzPQNYMRQeIVBvapL1DUYNl3uTJof6ukATzQTwK
iCsygNS3p96GVlgwMY2I2pUpN7MOSujsVqPDOG35txoyX/JujBy0+pFvx/XqVrbdVtuqV+rQ9bQV
a4Y2bOCMGiLFW235b9ci8b2mVjr9HGK6yLHTZYT8tayunxHkHAB//u4ydoJCKN0oOiXxGilK0GM8
C+z2X+lcGW97D66fS29pysyCDX8THWbBvUwFC3Hy49Hxx2OUyDzgBxPqq264kIvcL/6X4v7QB7Yx
hTG7s3NH3mxQJ/Q86KW7hsSQwuUJo8fLrkYmy6fHQjlDM3MmrsylEoqLsqNBTgo4tse6pd1M9xJc
AQu2PP+J5H3zdAUi7MPrwBH8Awq9lBszZhaoQxNGioaSwv4OmpGatU8kBkdK0I56/XIwgBhfyvHc
Xs2GDmZE5qNCnuByhsXq6gEyElJCvb+XHOLxOUoxvK+Uk9tP8QYmNqgiL/yhOXYv+ZFFt5Pkp7Gd
9q2oS2i2ugDD6mdTKqlHCPAvqV2xvIMXlnCc1ReeW5A5yNrWy8DWJgRZDeZZi/1Mp8Yv9Us6Isgn
2S++MMvMFnk+FQZmFpHtXMkm2TAjRHp0AictslZf1Rx4VhEzx9olD+bh4ke/2n50OfjLS4py2lKM
WFdqNTm9MV/nnIz03B4C+hjvCQwkOEDdf+2VXrXQUF40MijhE+jPr9bu62EN0NlvO3UNVv1+/QGe
1YAzwHWr8CfqK6QEwFubprmNNSdkREBxD0QGYCZccGAXou1kjaoH0jprlrtFaSWeDF5N7Uj4zcAx
QSCffeRoNWd78fAFJL1/pfz0Mlh6i3vw1VkYOBgX9jMBZG02eyX4hbmhf1gO/GImJIDsLWPmIQHL
Rw6pfoAqbf/OjjSNAyXuWx40DxY/HMlvb5LXoryCQyrdJ+tFEHjtKsaXDPn3y4ucpAdtlViHMBYG
GRv/sV3jO93jV0f9wCH74M7CDnOaMEZzGRWfiUha9+2ubPMrvUofgNWrYsUHcNlWGsL+tddT0g7N
wHB+/6SWzyhS/af3a5p0iz8kTZx3xkU8N1QQNOrszLrM0mzgyQWUBQm+E/7CM4+O1ZE62//QGljW
pgd4FjEVjtOPL0WXhra5rsluzlaMSggLX927PWCfH0ZoHgBnGEdVAv9FhnA5W9gbhrYYrWHK2vzI
tgYiNqxjlr4KCLnTef0BTiojxajgYasJUAvGfY84ph9ddjeynHvj6XvNDk/3XXEMELmfTL0WIosT
p7FercnmPjYUxquXOJ35jc6RDXM1vAZAGqEcoUHOJJjgkECxoXlPaxrVebXKq/YqC1AasleQ5eg2
MrPG0RrtBHIpAMHjAPoKEMjr+jVxx9L+ZwPDrgZp8ShqrdEINkRtvsVdoBC75q2uWW2n598NutYQ
Exc8I0w9+6jH/xqA1h4loSVmAmxc7DCJXaGaJllnV/H/aYEmsd+msVrRPYJzzJty5h+mNLzKbaSN
W/NKYiUR68Hm6WA5ew+2CpqU5OtkYyRjwwa7MnL8wCY8SucOccTsdVx39Arqsgmwkf/OxsfmUp9B
O3KaN2CSwI88P5w6SuID8CWrwYjAIru6k3NRgDS/27ooWGA/ZmXfWmxULuVBWhBYhyCXKXjA5Xif
zdRNpNLRCSLnP7p9ZUzlLlHdBI0CDEPVK2C6aajeAp3BoDnLZrkaCjwNFsAxoxbWnTuqhkDdVg/2
aVkJaDYf7mnWY1b0PpPYLxd6+OUgulm3rsG/1FgDL3PfYDT79p8h1wZ2p3E8VBIvilxDmueUBi9O
YeCRkfgjHHkZmEJIqKjjQa1BZy+DS6BAV5TJmmEuPO1RTljZ7hlJdpUvVEpzj63JwrMDH0yKZLnr
kTe0M/uwcAYkTEgDIqeeLK7x00IM8xnI43te0h1TZVfJB+7cjOVy8SNs0ng6B+tOA3sLFPGD9fdG
BQqNRFmhEBxWUvyWXWPbe7LHOloHjmZYwAeX915R0MemIiIi0Ke6lQ5ZiOupg2U0As0erS9SbAMe
vSl4YEkr+1Jr0368NU31gCe2Ho4QNOq2b2OWApn5Mk0K7iU9lbIdmdXYfjaRLJGlscnILcVlWnSV
fCxb6Beic7EOuv7tzlmRpa3xdlOueKir8vOLUsAyX9tjuPo1f82oNKFCBfzDpmW97l3eGfobqqMd
OBeO68wWsOmPZWZMtqPPOV6u3JKy+XQtvCSVnVjQ+FEyIbQoY917z/mhDxBBjmol0ovsaUYvNP3/
HSjqp0mPLT44AYPEbjxnBkw40ZQU2j2/0sM2xBgfurHDxtb5d5rYC9hZBwrwbatQifzUvbqVjFBO
NaYR20VlwJuO2w01PA2c+hpCLJtLqK8pn1Pt/exlOv6cVisl0H8UjvAdX3X/YIXVid0a4CT2N8Ee
IQVSEK+5I5I3NoQ9oUCVX2QGaFdi2CRlhJ+bAv4P0nR4FisGM+LzacA7jIfSmqYEpTabhdO5HS3J
yWtybjWI8Q4Unr45Bv2BvQLtWAQwIC7j4l0fQlQQeuSSYDjM+EmEDFEdiUGDbnxuZ/jtvemcWXyr
2w+ToGfa9SRczNkD6BgxJ2cdp06TjhQJNij3G7J57fgueVeBhudlS5vcLnFQgF/OZL+9Kzi5v6Da
547t4B+CbaJVFBMSxrqvEkUY2U1JnKCinusw3yRNqHBLmgMjebSloirAUHWK1KlnPIRk5MXmOcyk
AavdrRf7Dr++dd/2HSjI8yZFE42WG9dzOOZ77ldeyXUsUYR/ls1mwNBSJCusqwOgwINJc03keo/C
gkbC+TYngPBaskdDugqUApZStkFhseuqhCLxGML16Mh4MFhglWH0ZxIpyd/OaFCIbKW7EYs0MJHZ
cMdL6yevtQK32f+aCWL/lsEeFPK/ies36kDjTmwqf+AXV2ypfGStcte1nxfIt4tWi39hCg78GY1t
lhweM1u9Ihrh3bMiieIEs1f0SpJaJVihEsiyGEt/NJ5UXcq7P9C/Dk/CoXXcEqt8O1I6sh4tz0S6
gsMsjhsLfplA34+dwVDCmLc75SjVoIqGzM3Se5A5O3hRrIZSTDAhqz71LRe1D8qF0CY4fIbkPNrb
8oSDCsU9zpaQ0kNunCKsOMNRvw4quuv5z5TOSA1sutvcefnxIYCqOnObS6hR2mWWPWcDC8t+q37F
G8fOd+FM2t2VvhlRtI8RViiip0oOLlmHkvVryoj8K/uHVemBbwxtGjp7Z8FNR+JzTIuh8PkxrydP
I0oR/Xv/5GvRk8iArbeRHUQdtex7YMklIcoM/uq6oKWsyhKSEXe6yMgULC9J7GME2rTNUKQHyqHX
j7fBW4QhCQoDIGXrMb3vNICXzvWLwkbuglQ7XlqRviDycdo3DmfKxLtx3qYtPcP3IgpIuok2FvUB
KVmg3huBFqYD7kZn4O9bCVeYsywh7Iku/ltr0cyuMNinbt2UQOn5TmjmSHbKFIhY4Xg/MW014rFd
Ddxw67xaIUo/LizXpXu3WJ5a8MmMMwtNjO7jeSkni+yV1Fy1HWWL52yaTJiuXTE3Vb5EXvUDyEnX
R+4ctvPl6vU/HR9nkAjjZkcRiYxYEz4eQECxJUA9KO+Ot4bPwid8iZyM+YhBjY9fbWOTkvfkDqzt
6LUdmpVTqzJ0LWVGheJGt05o0EmX2Rf1Mk8/raK1prD4jgqBR7dju+KvEmPyXm7+yO4YaV/SeWIQ
lBb8Z7S2l3oiUVvtuSbzrmIeBLl3JRLI4FGAoN3cs1c49XpUjFYNXkmheb7SZvkHAvz6jFsasKnw
BEvF4P8ALZEWnmZEDdPyl9ypDMDBpC8pmCWrvWh81KEymrmfgYF2Y9mm6pjQBLbum45akRj+i2WL
+O5JaqvVS7zv96+rb52FlXK0uNc+VNQwA79NItSj6UGn0ILndXPiXPfRMTXSuZD0QXeLjtw0vzip
1+4ar5txN6mXmZ8badW7J5TAEtr3kboeETn5Ys/mBAeiLpiQ+GtIjk6pSf5VM+wtscbu7Sbb/J/b
Kt/Syd/YvgReE7Kfa7FFVTz1TVO+hfldZoV41dKGlYyjBFwC07WLGGoYCVQ4BFD8O+Rn8YmsHUsy
3SQLrztdzKmwewXF4576n3TH/UXkpJGD0KhMy6vLXRlhVymB8uyaP+NaVdbhm5DNxJT1a06dpoEB
P+rFc4VvDaJFo+I7dE6uAaPuYErjiRgiv6xur980dnEb7huB2bQvZK4D8nW55WxGlDX2OMUgyIyc
vV4llA9mbmtzRXAApFkg6AL3wX6987x2mDJrBoobwAKRqzQGhg+C6zjqxTLQcU6ZSvH1uXvQeM1S
WDK+D75DSLI4ZS6NvLda8/OCVg+4KDTKTN2MEcCvbMfk9epKgSJJQA1ZhABZiO8+VF4P5srtJRG8
sdkyCGJcPTs52Bwnw3nmlhqBhbiPAOE5GieZoe/oYrqqGYGB9Nn/4A9IWwl3If8Xy610IucgiQZc
aVZ90ynQ9h0jo04FjHFTfnkTW//XK2dJAe3S0yNm3CveJSebLMojux1l9hMrcydIDSfDaRYlB5mK
jwts7O65mYzUEKl5ag90suiQWHBXzvbcrsiWUvdU09F1RYm0dbNOOoq0IYVliomwotcUEuWQ7y10
GuZ/nS1t3/sIXvt4NAUgUMJcUTm+HKjS5OX3nKtIvCi6hNjlDtnKfPo8IT/KR6Jmptm0fEEK0jY+
UcsxtnIX8QD9Rwo06mSasjtnMSehzuvaZtSynCvmWcCCWlJoFiobsbjaYWZwT2aCtGorreLkDBlk
nMNS5ZoJjsFASlPpF3/D7Jbp2kQGj3q0KRaUbvLnH7b75u6+0U6TbRqoOOUtjbOWaAqG+zJidZ3u
O0hvn91CT6+vU4A3x9+e+EEJyK2TAp/3lnbaTNgviggzXjDgjq8yfmjM9yEBFAbS0LiJmtpmKdoI
XrXbE59h8UtENx9ykG/qjE6YXc/3Wa5uthQjlRr7HH7I0MvqPmAzlYAhnjBoRjODrtofTesnk74V
80hnvdYXmIxhduvN7djlxIKz6JoD4gXGVBSZBWXteblDuyyUtNKMEKcg3JrG1rFqFSM8ooZCR5Sj
7MFpbkms/q8QziK4N4Rkq0vNGQJltN4YvlGj8ejkxeOT9H81tU8fYX19I0jtVK1WN44I58j+EH48
+Rejv9GePwJSbcuMIfXuGYoMslp7+47NP3SgeZIN5JHm5WztZCM9v/CL6W2WkDtE0zufCGrtfPVY
IcYuPud3arNQocE40cImqwgYcPkc68SsrKu1v1plwx5+WkCRCbakrYj1WH64sdKPbU2EE+sOhE8m
taOFk8PwGuXKeMQcJBSWeoHLw3niliXvY4M810x3A7HJTDdTaEvpggKPyUV9XkzP0nDKImvDj5eI
mT6uigOTx51iLXVGh6WGsOMx0J9uc7g07ReC3ttdK1kdaZ1L1jxWnLThC6eIfDbLUuUuG7kHsHPy
1ml7SCNM5usEWEdSZG7Mo0LNaaKQNFZTstpXatgtI2TyQGT1bkkqik3a8DugHTN541yjFGqDPBJQ
DqCUwv0ZPFXuLT3uYvyG/xjNsjiTGJssjw6nSXxDJFfYjjI2ROVsEhI32vxv6vutJgj93hMOpkEK
9VyTPYa4zj/5yw231RzYBcTyX0/SJDwrg9whtN3Ymhu/FRquP0V2odkYYKr4VvsbB44I+kdCK0rz
0om+JBCRUn8HNROh6r2esZKb7mOU635oJ7Yfk3UISC6Ai9H1YHbyduOzXJ6jer9Rx+wwUlrpAuEh
VNv9/UzwrwWA0zsESqGCbFiCS39QP5e1fLBahi+h19R9tXQ3SZQJn8+hHURdeDyXGp4XXKHRhRJ0
nYE6jhdanASTBPmkd3fdK3aFd7sEOrpBEoDPqAgVMQFnIvpZd8gFzjpcJ/RM/DChvPxrQza7k4yy
a7Y5DEPYDbRKSS/PZrzGFE4FZic1AuE3FSvYhbVbfasEckW9x/guKB/z2TmD6uVgjF0ypk5M+DQR
pD9EprQOMy/GGXvRolszJ3AO+BqgmrZP4MEa2/l6kUbZqu5whJfj+clNNuXTwkedADUIAXnYVwkm
P4kVJ5vNCDYCC6tJwQ/ErsSeQXecnDKzBGe5djAAoJEcUcLLghbbr/EIBEwQi0sFQFWBAFCPyzNI
U7QjW4bh5K4v9+kLKgWeVph/eKjS9fBsBwlKF4zeFw4fqdmo56JxAAgAF7wXlB0Yxvb2u6DVpPK9
fy8miUuEuX7eiitbtyiPp6EWWPHnGF6PrEh4y4O6zWQfLA3G7Hd7u9w26eiEECqfXKryQBBazGTs
pDOGQIUTMjHG2Xp7AY8WMshQUjhfq3m+LtJtZrzTt9cwKNSn+j1fFLluM1FkERgiosNVCDgqd28w
91wKTF+M5yBo6tSU3R+1U6t/kCZae8++E/Hc7CMsxibKqQR3hjKQUojYk57GXDsBr1iwqAKjtw7O
zkpOvB/YOXhpsV6bs4B/Sk4UQF8/0afgIRzRqhrdgVF88GZEPwp6sfSPLYLRCOPUcQ7hhRlcD/lI
gPqQ/GCmMvU13V3Qt388LCtPJj1G879Ka5ao0mWI9dmTsg+z+xdM1xJXQi//2RvmK1th0ynu9AkV
KDE4/1OmV4300a7cfY0mS6Cfd6syVwy/jrEUbjTBA3fUSRN0xSH6N+AYh3F5uBd/C5advnBfBQQW
V8SPsbq80FsGj6W/SWwix3lwwEHL2hfHVqE5JYcQNCMd+oz0ONGNe/Kq9t8nLSMSflsnJyK1UoA+
Z6O/YAA7o4/ie+6DCvu7dBo+CBJ1fdjnlpFAW7rSjvT8Nf5A9SFVazAZZMlmKHDkRXc16zLJA3Fc
JiL0mnrEfZrrpcUsTU2aHjYpTQj+JaRcOsn3bvj00+43hjbshxoRI/VX5BeV0TK88WUNfpodosoy
J5i9+6mIacppJZvlIBXDIOQ+hO6tBcQ5qINXTQT7/Oj1SxoVL8z+4LYN8lODk6xRN7aMADW914L4
La2bFbzQPP8r+uGEmx609yxu/erKsBprw8Fq6QnR4RGfBLw37gXmNAk0pmHXqKSgDqcvNEFPEy2N
z7OiTaefcA7pu71m2nz9SOlm69HpbC30FHS80A7ctjDgtVHyTlmA25DvIGd54Bz9YJPVg/kE/02R
WBQeaxxTtm3bvrtnCNDy8sQ8hVIOdqgdMdYoWZCLEVkXFpvGlLs9rRhJrR5+hwhuI/YwifITrbaq
bCp8jkbSbGRwEpoZcLespP8GXEpeLYQTFapYZ8kaS7Du9EAQD0MYVLLcCVYOFm9TdqSrpCy0XS/9
NP65f74IDpbUvdifaNRZpYvZWzJ4XTn2QU3yInSARvbdUw0nLe+/CVps8McZ+tBNd1PdvtB+iHky
AfyutfTM7NzMI+RcIVNoptUqlOvKlkQi5nKoZ8IT05kYEsNzWVyHljKrn6j+CB6+DvA/k5JV9y9/
JsC00O+ehAYoxWKonmgoOaeR4FPAt8mQpN1h2nisLWlqp+PpiMDSQh70gXrDNqYFN+sZsIMmebpp
HSdUWq1EMlQ1o+MX0xT0W1ZodbFn7i3yBCwf5iyDV71aLlMm5mL6YTSu2wj0TrElUdfKNNgZ7sAN
JUXegNJ4zqWvHRruBCGH2R2m4gqpx/3Zo4G3dlH+R1awo0WSQ0SbVdhvAbKdZk6kQP9dtRNctvqq
RUjj5vhTp6fZUPThwDOgj34y9TVL7vkK/gIaux4T+Dbw7DE0m3LH/J4Wn7YxNlnUY9VkloFQ+6Fu
+1/BCpUR4J9zf09Ho/ClR/vajtxVUUWz4iLj8LROFIMnCR7ehH7sk+jnUqdv2T0DC8PmJEvMxsDW
RGgQZc26u92Cbkawc7kBI/dLkTp3EidzDR37Z+4bMV7gTG7iWviBpwPvi2RlpoLhK2k39XZ6O9Sq
ygJdfQeQjD1Ryqh78vs6JsNA7h5i5UKuqBJ9/AdhoYC83yX4Uc9Gz0iLIb3n1zvQmeMLOHmGzrrp
PvNeDtEjZBna8sg/YNF61IK8yoRFsU0z0r2etw2fCQbDlIDklIWaxUxr8wHfmZDcRvCXpk776iyH
5OLu3Ds13mSXkj1vECuiWpwv/OP8v6QcgbqdMimO3wZaxyy5WYtikw+/7RLndw77G/qJekYo72ey
pFYipugafp2/xos3RMzoAPNl3BgDQ8FDfdvDDViwAq5kphduR5BbFNhAuC6+iln4w3OeVOLDVnin
znUbbhfee3S9CRQksmIC1x05nxpHmSWvOhuztkRudEmI9jaLYxRhyX1dyXckAzouNw4jyhH6YCNX
rzI2o8UXB7t0Xa1xA6bG1x4Qk98gLkdWUIMMbXDUMT6T/Fnry1klcTV48853/gCSib6pGIBo/qIg
uDqbCmoGfmtmLrdlA3CGqgwtXRu7juNBTNf4bSK/Nq2kLTc6YBURrZv6eQAooXDBscKrVqpk904i
yD1WBQRIgFBhQYVrNDeyjjuw4MycBxmwafNoS68CU0Jqf5V46JNLtEoNUwew6QS0rDvSDFdF7WPt
ahRcsN/rUMTWBTizoSqZinUFqPXma7OmV/Ec0U1DHb9W+0yioOsmApte0rxI/AmYscsmJp/kJ+Ns
O2JraQOH2Hvam06O6iewg67++RMwg89pLckJlLEkzPRO5jDcXxIhoDxh8iza35RX/hTz1+qb4kRs
b363BtRDZRRj3eKROKBChrPJpVW83R6+tpRTxdj3RJV2EOtrxMKWaDu5DdxT+84Odk5JVFnbL4Tr
z7pwhUrhNisybeq7MLS3bfXSA4nfJIvPqbo3bVjyzoZXOkpD1+tizTduU2RfA+xWZsPG7sUWMXAQ
eNEZiTJqg2Bv/53LvN24fzs0v2PtvFi5g8cKCxVoMdkrn5Gdk8/PVthScyTzaxAvDsQcAeTFTk4m
TD6+/UZ+ZDuO26Zoe7B6dxhn/0uV0scT9B+r5Xc780XqpnbxylE6DXTR7els2XDS9Hi/otL7HdIG
42frIj9/Kw4BkVXc+8LkK8QVy+GajJz430b/jX+rOiI2+GzE3KaEtgvsBZ00pZV38gnormYWWwES
F/JAjRgoRWZX0L8KIX+rjUvyCiXNgH3mzNgKLjKD2FU6uM2AhyRBAzJnJspByRwtK1T4LQmNOkJw
ERdzAleGiMLP9OoraDxt/1PNkeIkNyQH6FbT/NeF09LYY/Ca3ipk/I3lX3959cLPymnPb3KevKxs
bKbej4v8gApHYHQdF+bR5GsFosg9GYduTY9jCyCEIRWGG9nYqI6zdz2VLcc+cJ/FHnSBIx6vJzmM
iu3UydGLAcP/cW4yvvQ6RsKjeVheCpi9mIzXnvWIpxV4ZzPptXgvdFgq4Ih7h2Mrv9lFi9ctdDK4
RWfuZmYTNvzF5iraTeEwoWKvArUNncn+UjvNk3vuzRzVdubggCQwjOa9CrGV9FUO24+p3k9ulxR4
Qa+BmQuOnUhBDPoQPJUkMZrjdKKEDZjQXaqtZdBULU85QjfTDyn+XxjLSRR6Np0eo/cSkEiML9Ff
dz5jMGXBS1FDfz6pscrUqpQKIfVM7rG7wGa1uzgnLMuCvnpfw/l7IdmbCCw6mC4TyXkqrojIQeQa
8uOH2W25nWxvNc7tmhi2U6aH2PMQfU0obfFQZnRXRFmjlpdVvdqIpdTL1sZ4W/8HJBAkCZLyWnac
yJeEn04g/LCGbF2Y3gpFgeBayfosgGkg1/PCQAUqqGYSBQu/2KmAqbyJlUO1ZZEMFJfN9gbqbn4U
SrzXs+8a27XN6hPXBD4cJgLhtSlZlUr/yXayUyPk+nhRUkpKGP4teCI0fIxQ3eLfyrMQOx+r+5Hk
bYjBXH7F7dmOivMm2JBdR/+uVKi2kl+FK0BdchEFYgrjG5TrjOQA+OxkeDGwsem8XpCx6MYbZLsS
yPtl9AoYPuqe5RjlvGO8hI3aObQnwVv7iLho1MonxvovVIXuw+JW3Y5EqfcOjfvS4wB6ZqS1sSpj
zM8oriYyug/yh56RqXXo/nt3859BYE648QdaJCtxZeLPoH1pHubyUswbbJcFn52lj7Ts8HY0FITR
t/UcjCWWCZO0qWuorF11drgIlGT8zAqU0ive5TtiWpRSIHYr/YEyDFoVIRogoCZExathHXpHJpJ/
Isxrdr1w186RKf6iR/ILuidhLNCLbO9AgO/U0Xd/S/Q40ksX2kbHXjjjdFhD7xeYHdQE0IKHePyS
4EbBLwYsOOF8RDyMwIgd/ujuy4Iv+ohFtMUDYqWdCU6VltSCH5X45PdgHbNSYXvRlxl2is3vXntb
caXUza5b8mhHSs/N2HI13KCYPfzF7R3eYhFUqCmhGs8/jMaNma6u3XNhvpFAU+7WK4nr7bq0IInz
5s5Zl+lWToEVj5DL7C1YzoiRhw+G5ZMMsI5puHUqksfdg53MJVKp7hX4z9/4UsQjDSPucmuP9sLP
rmXLOt5KcNWlp0UtpgpJwWL6f9qolNWLxmp5VphjNPdPMYdNkeMuPO8pP5YBzJgzzBw4oLGucWBi
LQdj/rJm9GZQTHMkh8lQFPH5hOaPblyv5zncZ91t5xPN9AjBoEBhw/9cztwK7B6rqn+FwVI/VkLj
dsQ6TtbHr1esK4tyDu2KYWhINIo+zhYmu5fr8r/M4U/dkhADWeHA3V/WXdSUX1WSciPiN/eIQki3
PqmJNH10bFgXVoyO+rtmCTmAdh7e3/rxDbaEr8MUj7J0WCq84m1Zns4IXbOOyapDIdqP3eIfNe5t
udBt0GIUvugFV+//KEzu1V//V6SHdVUT/UQ5rpaycf+NlpHyPy1Bw9H8KvD2oKGbAOvtzAPEiP1m
8SAFsRqOdKG6BxqWkFmXt0GGP68IQo22yr58E5fW8ED52nVmLjVSPs2fOtF4EL1AEErkYAlYn7qy
UJxafoGc8MVIsHxAOFUZhA2O9z1F9nQi89HsFe3ENMDuexdMqWIH920hCHDBbQWETcnrLS7lLjB3
TZ5ULIvwEKLSiSIbUvTzraPYWvZ2STezf2kpZtzAYxFLg7cOC82NMHPgKbNVK52E1ioCjXELolfo
YvY4H3sE58PQ9w09spRC2EiBD+Fwuo1sGAnOW1U070Ui1xX26GX8T/GLQxbDAHnYf3bfkxuAJEYw
TG0Z1VKprM1XgQnyS3R5snVCrXNWPwDBLUAQUV5WjM+SaxN9Vms0RFBqIZMeHQhHJYEB2mxKfMh7
hlMKyavqJHpv/YGenTxh8qwCcvOX3oNWd06ul3nCMd66G1zwP7F6fQ0U4CZfn+GHpwZocpXAlgHk
C7L6ZajtlsdevhAV2IqdXTW18KAQrtNcQuIGEQpx+YNKZuNqki9ZTJkO6Y5aKeUiIini2eIHDXmS
azFPshgsJFnL/EJNaWpsfvERXA0lqi3TGsmPO/ebLQVCVrQreOLdn7wHwpUJ4ysI+4ybLPby5Pbq
Aw0jUWEddNDX1qy9SwAqCazISgT0Q2o7b4k+eorlOnkMUDoqWjnurckfHZz/NKmdmPSwLXukFsFz
gXCnNTP/9lLza86Nq2xKqUJP9GOBtIlkN2LS8AMJbU39PhfXMWh4ecyzEriv5+KN88IE1YyuRzem
hESEogmusDG8hyx1YtZQvxtg+ZHeRKETpJeXP+xuAg80U/H/w8CgIpDqu0sGDYseQTttD//kRnHc
akIFqssrtnNfJ28cqRrLqhcchF56inNprs6cJg0Vt9Hh5s3Zt2FgEyxGPflRh1lwYHuHnEVEUb/J
EgUyVNXUR4Jow0C780eWyccEZD2F3fuUAO7DxjGAvDw9ApFC+UDFwGIVrtTgS8nH6DavOJ5aqFer
oGwVxybMyeMXfaYSaPf60AvlBkQTzHjODu9Qu3kJwk2XIgka3dmtl9Se7fdpwJn9PWrbirCgnrfk
taPhU8A3uDZiHrAGWpnjSA+1++xsC0akJ2wnTF3m+g2YplE4tl2WRZREEXVd26g6oiYJGlv9JpeE
isznjVinlKcWqCi0fZHwNhtQZ+TXyp11XxK8OHA0EKyZiQIqhx+8Sbj9ZNCyWxOFvMV6O7AhDbfx
0vFdhkNxcLv3Y/sZkHDPloOISQ9g/hWAl4taPrPwm515fBoAAQuPAm4MpA16yMU1KZc1syiJ4UfP
7gA5RbrHItM1bHI0cmocbsaMyO4BbFHyu9fYlj2tzEnWjvt4eb9aozLsDVA4OAuOm6oRXs6pbdJx
ozstjhpSJNXojLAqh5/V91/Dj/2BRWNhhnGd0apv+4Wrg2QARt+WnW5jcKx3+rgIbBx+t07Fhe0l
rvxuFp6c6JAWN2G6eMPBAE4ye29KUGmFSsv1Nf9BQog+JGLkxlndAk/3me4q6g8dqmWAyHRbmxvP
6hp8RSRh/fkg209Z+9HyBS2VDY3rriw43lASXap9NkL/VuFtVe13o/Vu20OoG8YDnO5cpPtOthbj
M2WYWb+stcwygwUeQ+/9DB7HsKdcg5QI3i14mB2C3BOOwJ4sOjQOZTDIHHOWV38esPLGXw1ddvKr
4AeIAD8XPR7qldrJP7gzcfa3Le9SJV6KN5OuImfOmRjWIcQ2HpMnBDLErxdMn9ZV1vr1zzjsyJMO
cunzl0LijDWr0mLqrjhS5Eokjg/q/R4RD6DHxJgugJTLnkw5gwfFZv8rUcmYgNFKlWvHmSStvcQw
e9oh4gvOlnrUsUjm3IPEM2PoosKtGHumYQGBHfBd4FpYP76ZtuvDJhE6i/6HF/2MopYTMXWRKv1P
G7e0zEK4m264k/ZoZj+K752/vBf9b25B3beKaj8R0sFEPT7NjY7rp98cYZZMRjcmT0Wr0Eem8CVz
iuSZfYgGhR8yjedRoRKD73yyt9RIbGjBLUwewoSYc098KyJoFQYiQu4ulViNWOisFB8ppVqTevro
lEEvNsKwfOCRT5zfPVhLLuFi03ePiyLQnxxjuFVWr6QwROYsDrNtJaEDLCzT5N5m33zBUuQ0OPW8
tRuEhSFOJq0mk/ZFYrXvqkLwKtnqMX1fbRKpsJwSM7CiKmAfNtlvCFmiDEmr4T9u68i2hzKOUUuw
tJF1DUDw8n6Lo7TrKbCd+zxCB05trmgQxBZnVbhyek8U+hffND8nJ/y6wclskH9RAERSyOblomVR
67X1UOVW02lS6+gOKn+kYnEAErRMzcYVoCpyGjWiimLDnv/e7dGbLXRaJI2SQ8NDHM4Rzy8NxTin
xd+OxfhjmAqv0mYYT1MKCHx2WRVA+Kpo4KbYZrCNHOsPIQKbbDApbkK2tKlv6qf/RVyeqCb0D5H0
gWWz0sy2XX1yfLJJB98irI9nsna4pIWp3ljbUcc3/rwPAxYvf1ZC+3IjGfOCqV0DKEo0j2ckVUuJ
wlHJEaqZx9jCTkG9CXhBtAQpQXaZYWN+tl/CH5pFcpGjbUB1kVBb6r1sXyFSxQlH8c2mYwxQb2vg
CCbcOtsgVlzkvmFKtsrO7zPm+xiT7d3bpT0LJK6d8VINTGFNpkZOn2OcoKNLUclKBydfK08qwPpi
U7ahdyTI58Lsm3YMX4vPQlg0xv9no4zjUmFsxZLJABu/IyJd2lIKSALzLzkcb7CiU83h5dEiPHPy
Gr2M8ZLAZCSlzfvZ2tkHxvAsd2slFC8e7sk+homImcnDTRvYmTnOV7w7ej6hXRvo5QYOkbiFzEnF
tc4FGrPE70BHO5H7nFqBWnBTOgBNS7oLO1zGige5MARvxcTHSToqSEiH4cXW33dYIFx5bVPPWa36
q3JEn6qyXn/KUE9MlTFDMKa1mnq2bRYaXG24+el2L8OwAs5RXZsO16g9k4/rVsUKJSbfXHciMROw
DI/XoHtMZekxfXWABB6hs58DuT452qiLJI0zka0OQmjTj9OSPjLpZQs97EDhLZfpgglL1Qh+LO2p
wo0Zy4/C+ayOUlqLNoZ9juml1ed5UOm7RLbGVhvqTl6ADvHWCbLgdVzKFwXTR37sPIOLoOQmPLXl
H3zyVvjJwZ+as05tU4M10YwLa6ZqYNNUB13kGzooIi2W18AEw0ApQcxNe9hDGBOIDRaF1HVy06Uw
WLqlttPJVjqKdlj24+vN6Mr+DCMC3mzrVaEWWhCksLxfEg0vrPm53mdqMVHYIkbfkl6BoMiQUJOl
iudPPI//IKegnpgHA9mQeAZAkV2mZKdEBIldVUexyB4wauliC34lQpiMXwyMRGgAp9n6Y66jhpZF
p8XlOT7HX7vOOoLbB6i8oex68DomgxTnCsSyLWA4E+cHD2VF3FEe/h1ZW5u1OSVG/crNQKd/xq9q
e1rpWU4pGTpPF02Zz6i+L2190hxpTS6iudM5o95QB5mRmVVIHBkDt99iOsh+Ch8wra9CywBvjYzy
PFINsRxMauVmfd9jl6to+D0ELKLwhjkR3cmqmejUsjYnvFxSt2cxsQkK7DZ6ffz2P911s7Vr33Jk
+6yACnAfvXt1YpM64IN9+n/dn6GeNUMTQwT4kNq8Z4jT6XBY2uC99z6/22/46jzLRmq9rJ66RPTJ
D6GOO6bZg8tY/KLSyCKHnr7Gw4e1Ibf+5oDI1kDAMp1Duktrzsr+p3uvMpaizb/Snkx59PZd1IKV
bLBI2Sdaa6tRVXms6MN05UtlqwVTmuZms5tOTpQpimFo4ZXx+U6rJ8SE3DUlahWpvRIOi1BlCLLl
Jeb9J5Lzu8hVkugmPCJlWUNRnO0hF129EhJZNrPNQa1riQ3S9UT6kl/mJesd3ifU9TaL8MBVgU4L
NU99TTMb3yY7EER05tAZMedfLpuJ7nCStfEKnrXa36FuyT05vp64F7aFneSTl98hRz9UIHRUpek5
TVvzDmqDXOPZ0Zh/JowOcZ5WCS8wUgr9ixAqb8Dn4y5iVc5k8Pxn4MXpMKbQ1uPnHJ/lkh5+TJit
5zxexKF22xH5Rw66QNHODdfD3wfHni/5RokfSI60nIbKKM6DjSBtN23hBjrm1PJr+AIqPe7tQ0vu
5/ZjWJyPhg+9NB2WF+iCUFDPFqPi1jcQgEuhu3o6GhKw49dHyFzK0ZkEhIWvEOOJKp9OwheQAzKA
wlmgimmhfH8ZcT8Ez+BUDhj5hv3tCgoz7kM7FcfLMs8O75P4Ywcb1njCXrTFIrMlz+yDqhhO6kAd
L5j0W+M+nn+xxmRX8N1UiCqpbD3QnmST+48hYKz9ToMI4xNPVwAdNj1Tl8m7E7e3DgWty3IahKsx
aQLWZ+lrvJvmluGJa1n4X52RbwJZTKRSB2V7a8dHQfu+3DpDrPS5rUDx86a5VyxpyHEVQCqDp+Ei
yNJqnYLEg7xv6mDYXix24ypBBXxxbvOGT/17ZtYIQtE6Ih6AE6a3E2bAEXgKQ0DgxORTafkpT34a
Xb0RbGoeacnmAGw+0f+zZzubuaajfSqu1SfMhrAhWGPuL4KQZK1EoCenaNBPDiZTF8cTly3n6j/5
+Jqfbgk5QYoDUnzjhPLCX6gk5lqY6vtPeO/Tr0FEsNY/TQa/SO61DEkYClx9Ebx18PP2kHpgT+nN
7tvROHERrksG40EI6N5e6cXhhwVESTu9gi89YIl8Pu54ty330QQlXzHZ9fZAWEmieSBboYo9bUxx
XjtpqaHMWv1ZQ/GuLl7GYR65wtMS8E8prFeUKxvH0fAaoXL1Y4zUH+sbGRNVnq3ieT+POndmF+VF
YlAYNmiK3tSb9xN0FvqTQR3dAF1qpq1ywt99PVgJPgk6lBDUjY536d0odBVfPLQ/F0arRhC8rM55
8+xqraaCQ7vhlSPVv5epInQaRs0eOnZC6nCi/nVGjhfTCwirnFCRjkqu6BFQb/AoEuYahN3LPY/J
0pIzmg14fOndxKZJAWgDYk8+w5cL7E1JC/gWYoBzskfqR3sv4RHdOI/Pu+6VJ5m9j5p3AOoviNYv
WzpQ5YassRQqBANrX0+k69mhDef93Vq3A0QFlkCJfm/O64TIVhlAm7YGJ624CcGQ4mR7pCrwIGKP
67s40c4nW3GKuXdnAfmrm0hl4JCfwW8RjDzN+d6Azdpsia7OycMkAc44aMgBskKagzOPCyiIouxJ
tlgb2ZksjX239pG7e+oVGYRrO+doXQoBqc23/srjYL9//VAditLl397LMdf7x6ZE+XDs5tAPgGwE
ShN594MZQ4drSYk9981naGsNs7yj9Ye4lLB0FvxSzU7ejbUeEYxHoWkOc6frWlexRiK7weQX2kAZ
PKrtW5QqBzU89MB0YYJZdeCMcmeyBeWDBQYEkK/I70wzYDOokkD0r1b1PQA6RKmsQBmgNLdg1+H0
bAZ8pfPZExY9n+zo5l3m1Kwpw0k7TCSGA7Xm2p4i4YldQhPiMTexfoZn9pVkfehUEpuhwjrlEQj4
67g3awG+y+hlmmOb1fVsE3rjQLn66UW1J1hsNLi0q6D6+Unoo2RUXOP+s7pa5BurtFjrKokuUW9X
UXzxQJQDAzPJ3Ck6aG0Nutxh/9bf+HEeqm9FY2Sl08UgmXx3htQbDegHlczU+J4Ojk911d2Evu0J
V9kBCQWF0Ztf4psAcRgaPm/gH6Am2qjE3epLuTLedkkhJNUGgVug9vcNEzOtOtlylJ7wRvhoTAIt
flvjm/tRJYAMqMWOiB/PY2bmtqysn8FZ5ha44vuB6e54IiV7LdxHE7ud3W6cctAj8+wdCWou6yvE
bVZ3gZhoUlkfGzu57Re2mBU2TtPgIKTKjjoSFrKw5PHMSF5u1xcrIzYGTUnMaMfXGcuuY60mc8B9
iFylwfncJifIyElk67VSa+Z+kOq33M108aKGnDzC6VS5mcoC1yKDK+Lpr/t9LfxZCjKzRdc/Yau7
aEFF0CNjWs8oxuvJBAZpAupOOHldmMkllqBvVFxZ87rwY9VvzSJ33t+r82r9wkvEAnDFj13VFvtN
s5fJjVrwR0JQBNYGJCsbazPRWIyHZWm52gIQhJZW7d5hcKjni//mwihttXckiyhlQQ1HihDSV+z8
IwY68kzempVXdQzfQjn+wekM5n0v3LxsypTmWXAJ+6L/f14tNc32FzquacusttTWiw133SI0yrnd
LDb/xyKI0BbT0Utv4yc2257M3LjL0hqQDa0aQpn2TC5vjtS+6+YQ9nw2DfNJw8QV55r4RjyRhMEs
R9coJP1bs+R5r3FWGi1HAfW9nuERSFzsE+JNYFn/qauG6wk9nSzPqWv7vEOkOQBUTAPnhKKKymrk
6/prlU0BKdvJ/TndzbqRmLtW6M1tE2cTs4BUeHnTjPmquAN1ba0KsjgMGUaQc6WChoA4PPCno7IW
coEEoeWnXJ79ggIPHyxeC598x20AyZsLvlZRdbFqSKda6BEnOx8W7J4z5ApXMwwQLGb+CgVEbbxS
rjc7/S4iLwuhwkC0CWBdwHh6D/5R3UNXkkPioS6ht6LC14ev2Sbahwd0ROb6j7eSKTshZ8ZmSjm+
BRf1sn0D+b/0rCBnKtdpluQhc5FrFRyY0LCG7W3KHhzjgIIX+jAY+vUvzji8d5TKyXX0ezd8Y+WI
oJUYdTzK2GUlZjVgke5P8f7+BBLDAA/WAd4z/ASTmgW9Sbt3r/SoxKxZpWP8Clsh3vPI6bq52zzG
uegxxsjjoBpVHxwCXTnePZuQMpyieVx8O42u+MNKpJ8CCLpvN/leAKSGCBWvNwmxTmyHKJeAZ/FA
nt29c5EOioM+iQkvYwgJxlvGqgCr6qQQK1CbAryC5yy40DCPB1VklW1ccygq81/MjV+huKh5V+9t
Q52xnYzy1Lv8338DMZKnVHA/KqkNn46qRyOaqslT0WdNH13O3ebaUBaXoxy3HQz9mEhHVSLP/R6b
G2C6bMXMhMS9ZV0xIPlOenUwhi9O+3cwXGCfINZ1KOA7AnycdivVtU6mg+6cQs1qlVwF/+rPuS9P
EqHoy2gG9GcJnoWfN9AzOXJG/mLd2xdKxaCJtwUv4Xe0GI0y/4hN8Mq/ljXyCoEn5FMEhpuVyTUG
oxCoL3N1qBJv4AiX/GrOImgbX76MMHGKdolmF3yNrlEaiSeaW5T8D6zguv3h7wLycQ1E9H/ff8xD
Y0pxErFCTYpPZ/AGQgoko17hNVNsAWa9cLAIW47slc/GCaSy4VzkK/PcZAdQB+QunDTNOwjhQbq3
MfR2c3f1GWVRXH5zW4UvzaX8lVBRz9vlPM5148rlCzNTOLTH77/an966/9qSjG6SlMydNgD8fkAc
sVybKc4HlAbzL49m/JRnwGbvovdbJ1OGqAON/EO1hnOQ3A7V/w1O1CuT/JPg6iuJti8QXVIgSwCV
1IIMoXUnDc8zC/RkDFuBBNO2NpEb0Jr9n+NlH2ixaRoRzTijQv91tHkI/D8a+R3EwZ8pRRBFLVWk
LHn0si5cRerwRA+2y8ZbA1IsW96qI6dfUNZUUSCeMB/FKZH+RN8p3ov3ug+dtFZVZkzOiGF+6kv7
buPmlmRHS+gIJpBQ84R8X3++XbG9NhGaHJrAcBW6/rLVAWzalBm0cYC94h9XEXV9mgZ9rW5F7E0G
+ESNjeEuEVlb6fkARDyyFQyxUKsXkV+34ljXjXt0xzaAmUjtlZRdif12HxXGi3lfqC+rdaWqLiAo
u0TYSU75iO6dPOZxRPfD+SXXq3RgW5QSHdt2KZuXpmxRcnroJPcA8z+Xx/YopwabAkeFmxmSXU6i
hY/jMEzQUrr8QCxiL3sylAVPmwidI4rB6Y/fAKEcWZTvVAYvvqFYR6DdBNEIjJEK/dqyns+wYotF
954enfgvFU3Gju2jUQqnoiMmOcbHABw72e08HDrB0Q3eoDdvkEfrDWgkiWXT5xvNKms/vty6LSdu
RYNsEMKM0+27UBhZ2OzsJJ/1ps+OuURDO/canT9p7BN/BjCxA4T/WPHeIki+ZldToTY38PO+bSCW
fAfA1HXHq0ocMnRHqjog0stwOcbVNAosbvgkfymEeIiasBdM9EK9/z8NmdIwAjhh5cGcGQ95MoA2
kJ+YtbVr4u7+En3qk4BeG6fc28bK6nD8HxbTjL/ExPamoPEPTUSOuNeDkV2LH5gILioTNhLfuQVs
4Dy27ctWuSCvSt5tdvpMWNJkHNyVv/s7yzuwrLumqmSNA+7oL+HknCSXVU/DfCjYISYV0aanD7SK
xWqXw3Bj9Ja68P2oFvMyf88hUTK0MapA8y/OneMh0OQudBL9MVKdp3yQ8lG3kfYhyZ7I7s/gmtjj
+faWPwh577ZliAAwByATns1IxT6i6K2gkcLlOoam18V4wZpGNOTGGAle/RRFwEeyD5y+jDAyoqGg
Z3NWp3cxtAbdOdwSpWZ5XWQSMGMBR1aFd95Humr/8LitL8dIi0Rrfok+MZY2T6aAGOWzpv2V0iLJ
/NIr+jT6NJBU5ELtFjYE/VVyGzHremKyDe9zdOljpD0axxKIPY9KzmNAfVi9k4rXUnVWgK/9aa+k
cIwfyWs9doZxEs5LTRK6vjb7agX3mLN3vpTnd5lS8L5RgkVidGv2q1Wp9kOTMY0m2I5P0ng8BYor
WvPOVG2dg33krQPsOIxtBcnUEp32IWaTWCmm1QLcZFQqkUc3D0HhHP9PjtLR8xdXbeenuBW8IZTR
tQU6IzAZI6LbavidXT8bHs77wi00PtQMqOt25ZUQdzrWrNq+Me0RFwAassEzO5fPOXrw21ht5uSY
kN66Pij7DkrmBJrsVix7NJTUG8mFTU+LnKQ2T0c9qTv0sN/tl8TBL/N9Frcw9q6n+9fYQL8MyKhz
8gfg3grtAdVKuZunVYgi5JrDNZGYY2nuSys8jDvAuAvfY5DZZUmi4VUxDrN5fDyfbR7xcUlfDB81
EeKpdTLaPo2zqkethrotqb3Mb7vdc61go/z7k5G9j0qPgDm77tJLNftYsnCsCbFY+1fizxtiCVd0
Lcd5/a5dIKAO/Qr22ABeMod95GCMZHnkZhzfPwG9Rut6YPhchycc5IoUTElCNdlbtyn4cJ4NXEQe
Y4HgDmTdNjp0LFWYSPYmlL74vuOfGxXuH2kY9aVnNzLv140/vWpGTy/2xK/66NYDA7/3lBMh5W8a
GTPn/vyBCtqzs/7qvXFZbENK9HvR2zsNST6zcwoWZI6eNHm/mYnq+qbz74B0xcB3A2g6tqsLOwKt
BCFnsc5p3WDN0fqyY1HTrCcxkXV6s5URDWWygjGw2avwEHH3Umxk+09vRIoXxVsocga9O27jrpRD
0mymUbrwCZzYe304f7+btqsJEbVxxnt2M1GXFgClJ+zuYLMOcwBYqbNCAibQ4bidIR7653WXhKMv
c+1aLkAw49euSP5a9YAW9p0I460AHrXnza8Wz+cBtzUrYQh6S0FVp3Cfb+BSF6ngrQaZrNsJZDNm
gIbN+lDdW00jwHc7NqbpMm7v51oKz+Q5VlpUD9NY8R9cygP1qaUiMcZM7ZgFsJmX7/z/tVn5X9nY
VnJRM1jz5a0c4AL5qAYVPb0S1m/iFgojCueR0bVrFkiI8Pti5yxyR/9LScCJwlX6gELsm4cXiPdd
q1gIpQduvbWWo0EXh9kelBCzxD1TyceZNpn1EiLLGP75kEDJ3JvVsC1sR2mLvduyEG1X7QV9D0o7
oCLa0k0g78H7uYmnfHmV48wpXjZVIHPbvsTFIpIyKCQ74DMdd1YFx1Ij8HLtdWREJl3h3nPi2rB4
xIEdxA4VeFxdOka577jgscfiYgzwcOoW0QQCuPwHUR1Sh1VIdAJdmK3JTY0L+tA7X77+LAfFY78P
stJU5ygQUeWPHXDCbrVELCqb4zSDTHMz7UxdCw5x1M43O8N4AGWHxX+y5mVtRtuZ3b+LC3VUjszG
2vXlKagkgD+of/dg0NWU2w72yXcnl3r5zS/yhiR9CLBZ+UlHjOqTybfaA0Z4r1Rmw81WUnZ0jDWO
T2gki1WxJd41iVOoLMXXux8Ae/+UbBLgnSsEsjZfqEIrtaH9Dz81FKcbQS03iiQUSwpQfR2B1bbl
UWbKIUeeaTq7NjvEqkikgZyd7zdd4r3rvHWYvuaKwUMrT4D4XnpveSuUxf8XeQH3D4ChGdgde5Fm
mD/E62yRwDW4oqjj+tZePXcgkOk3ZhB6cpiCI+XB2wMohhW1lVOlg9dTY7d5/kFZWHDCoX+Qiwo0
nQcc3PB6GWElUCEnpCSYDfn4rXBTvhELfIZ/zQP7b26t1sFYONYblpYbvpEiaJKZkYyqDKfgpy90
+iV7o6ruchcZb8a2ojYkL0ftK29VKuqTGmqCqMzpH2Pl9WQMFONpnqoJB9X9CPFrlLgCgqalFDZ9
ranWnt9BlajpIfKYx7NOVbJ1Ob9EbrpJx5MzHo8+QgU+ZkDXgsBIVB4y1xIpxrvmWO2J1lpJSzJd
l2Ll51Rq8OD5VmQvXN6A7d/u/ZgTu8/SEwSmiW1Ly74A5HVeuvxhJ3YqTm6pDFNDTzMkc3EPUaM7
ZMsWmVU+TBV8SSTA7bmkZpMQQSE6+wF/PaKnE+S0q1LEG2jabuekj21cyATWbVg8TZmdhlsBZjwA
kZiJv610WN+Z8YuFmvfL4oapAXEqJzGDKFlOtyft5NmzQMPoFSPckM0D800rXcwBfd6biR2V60bn
iLJg8RxK528VDJYQ4irubUCjtyjoGrOzUFgvJ5X4X6WGwG5Rt3KmULHo6Ri+w56t4AMAiJTRXLN9
M3MOlgDjwLxFE62/OpPXEEYUVr8Rv6v377XF+6/xJ+NIK2IKf3xsbEmH1Y0nOa5ymcImpC7zjcSE
pglKOCfPF4mY1qID++ikdzuvhB3jsplOj6+Cese6UEk69nVS6mBAKccFFZtyeLTppbRgYaMMNegZ
pNX2g5jOqfQ0nd8doND6uQG7WAlrCJ4l4VGvtA2AcUUqNRXGuDsPfsQY2KM4ZaRgumEsvbgD43cF
FfSpnNwfjIhtgrZTTRkMbLM9xxjkZ+O54lGnYrkmhyJEMW87nuqPn+9CbtpAi/yIGx5zLf2ovu7W
UMhVRbEjROl9hW73vSdf8bO7LX5M5SmToJU2WbgkY9sfK8TXuW//tbqzvZtuay4ecdwHAUwU/TzI
bVteyeEWRB0Nd7jg5nGjuXGVGU+U06DGdcJTjzIDjL18mnpjhp/Jw/MVyqjSRWM2TIBtkjsz0OaZ
CJ3OHROgFzSN8hkhNJee3YAgXv4Rh0XTTgCN3vqUxdHsaePwjfH9jLriM+n5WnGHiPqIJC+vD1Hf
LQuMTIP9vWLAea0/TwyQaAcq/YHUV/VGfwnmAygGNcedKGSfWkiuso6iTdL3mzZTZGjlF2TPTqAq
yFGOizQtbPyLS18BNPHFs0iwOqJFkGn0s1stwYFQSVmj+FSFxqhs77di6AgzqvQ7mtvjd4V/TKkj
dVlzkhFJS2WmF4O27l2u0pzsDLGu6JT6T88g7GwTYRC5wWlXbz1SJM4RuQmzYVEs2NgNqaE6iyem
0rXRe3ySY+BsEuLfVFfOxs+Lyb/dnWsvQH9rnREpAOXYL8pFnkqErlDVDHBNHVJxlIyp317RReqK
LuMa5FgDrtiV6tgNVAxbFSkda977V5gJg1T5wkfuh9z435VVjYiwZKMtfGs3f5pivEDI851VDbyP
svHMoRSYblfla++qVxdsCPFyIJWbLRbEXVKlIJMoiEEIeQfGeXD/Qcz0Fcmzx20B43PdYLu7axF7
wohj+tdZLIsy/7fS9XIxr0o/JMEW/NecLLDfW6B5+pZkgqaGEMMNmhJpaQpkgdgw9p6GythKkMlu
sCYI2JkXX3M8Il8HJjP067csnkDe/0P1tjVMBLKCw7wys22qmnl7hNJqMop+2+jVt+kBpiLkYP7M
oNEpD6CgPWYs+zy7HzNBWCW/tdBbYw+vErnBFL5qU0CrIh8dlOEhUiViTPEnwmh6rW7YNpUR82oZ
eOFI0gqGed5+OZ2+jx96uH90QSWlA0zeDtP8OpYXzlEOTPtEO8DTB7czhwQCH70YlnnWPOJUmQdX
J5lC1zOIgmFmSeN2zHSLlUirNaH8X8MHJ0H/L+SZ0e1hNhc6EUZtpW6uDD/qTgdzJk5tNg4lkYTe
pxSTH5CDgqo+Zfq7jCLxofzRJiFA564xK8ls2RHPYv/3AlQBqOiC1m72e6T0s6XjsEohGrJVF0YJ
NaJpeWAAgvez4JnrdZnUUZ5Q1YujsmOngVFPzVKB8ZwsyaQVSkc/jeMC4iF2Deex158+gtNvsL4o
HSw0X5Wz0Gy5+DrhJd5QPWTaJufuidZigvF7aLUcGVCcBBuWbWgYWiW2xQ7OmMXYnxCtsZazRXrz
jzifobeiCBLZQfrjT1tWWC0h/VfYPux3C3VLhbqR9ioayAgA2adDGzwr0NzKSyF1WlY4zbL4MOoE
LEYjbqG84jX+ijdrbkp5bekivyV4XJ2wZtjWQI2wGEypESFGj7q0vydKyQsVffGxHbPzHDYafTma
KO9msOTnHXHjmjfe7oTER/KZWPv0dIVnvRguhFWdekVystnrUKyFEvo/Vl9W+dYipnidyiN01Maa
UaaJZLS2mE2F6R9dekor/RNjRBN4xfz4NEycxh5ROeLSKJ+FNY44JxBK5fYbldVWhTQ0Qdxbian5
j3hjqujWk62bwSZvNZ3aJMVzreMC3QnYGcaFvnp2Sk0l2xxOpBg/xRe/Ji3NprH5TJ4KCFMhy8Rf
bIfPKr53AIasGLkwMqmuLH0a3ccZbNOvfhJkzGI0UiMwc9WvcLiAfU+PPek8pzrQb3iIQ2juGh30
bfmZpH0EeSD26j0gk47wduwEtVzBZxhOcAjmKOf75/4/JtCuXt4ufRs3ZWoKzOoEM1la8FcYmaEp
RhcxW+pqd/NM3EgZ9w7dEZQgM25uclOWJRpIayAjuEVMd6tvaHQLjf05J5wqHvfFb1YSjsO6O8K/
vC6wm404t8MKYIzsT+NIvsu9d/ZWp1jk3J89IgK3jnanxE4Hmfb3Y6ksPWRZMUks/l4RV3UQ4yRW
HPpNLHgQCbAimAz/QdZ4mZhXaCtDoj2ynjPXkre5mX7SBiUpsJLC5a+mVRRSpyfKaKqrUZeVlgkS
pEMw0pHnlzhaUj4xalJImGaHat3VCt5uQUdbgqyF4F26VXCZjLvoVaBTzLZlNkn5Ns2CJyKDLDrJ
I+TbOVam13pJ+wieUQBLvyeAFpDdpuWFDv8WqvAqVuRyBxZ4HqvftOcPJyDFS8tX05RAgFoMnkUp
dxs3onGysvjnobi3/FtyJKHPEBV4SHYezNFx+oG7MSHy3IZ+MSZo5/8yx2sWoezN3rjY2Oyq+alR
wG/8QkdKAgZ3FMB8CvS2CeN4zNNa/H2eqGZ4Zu6HGY+rDRlyeR30aly+xlkTQChmbitDIcXACKYI
lrHVQU/v2ndUMW7PqNtJJ7r6tw6Vyf7B5O7UwBokH20Npi+JpAP01Ob21XoM8EXK4vwPEUDb0RKI
RoKf5BKRwmMUadXqevyfUS4k26SQP9qR/q9Dbdv0Io4nrfmEI9qHcx6h3z9NnNKW/0mPKAnB2B0G
oUVEvgnoW9MMzr42Q63R8yadkXZs8NjG3090wHTfve3uH+xW9Emq/qyKlXMW50431BbxlCdi4Bx4
g43L9Yt+Vt/DK7f/rSttV+kHSoHIeRTiVFASw+501ayAtmTGO4li2dMMR62veX1GGvOJ7t9Qm7cb
5LyjsqYmheGJd6gfrYlw3D3y8Y8MzeBHOEm1QL1aS3AmYm0LHgBR6yhbqSJGtr/lZKuowlPOqpF2
k/a0iCOFEdlVx4B8GcnhYSVtyf46FKGPesnTDzxXsz8n84LBbAg9oXH3PAXvdx+O5PxsLIUXNWpI
ktgPY3Unn9rQX4W9eoWWbhTvoYQbHwxDRk3+Vu6YJqu7Vtbj31VXKnz3w52f1kc+iGhVlLC2sz1Y
NMZp2AV+vwnje1dKSF4cuKdk686LwqZLyPHZ9VbCQ5Og+icfreTPKakuAULypMnN2g5v+vdLmZbz
iesaQ5AKPqDFVfEjbjpd3VlSILtozBhM42daFXT34bpF5AV7AJVnPGN6uxv4s1RRwyXn1ZshTkjY
ue/YxF+pd7IfkCNQSy3A1Rd/ATXq/kOx/NHa7UiJGcyN0VAOHP6DSKteRCb9mRx+hyo9nxS65ep5
vgkxAvVIQZvBwN+BzLk+HDBeqoUM2u46EP1dRIiKAJRv2fEJRCrFR5NsyLBoM0KTUWiQYt1OPe9l
wuUOZvgM4noN+/oOdgGAdxJT2JvfSXAxoauZve20hMaDHAFDuSDjv4pTtKVplJLTX+scNG9tciu/
jOWKJnIWBsKhbXrPe9KlMY18EyHcElD5bgTt39oT1o9igluV1ABXCAwVyOE/1KIm0VrhXwJCgwft
b5Sj1Ktvdv2SVrC6O3w3IBxFuqqsWEs82yBVxNimBrgYTuBnCZjd2Jw9dK/oB0ZrH7LvbWnhb0WN
UJrCLQ+dkzyL8NUHHgKXsymmMxy8X0kpfNZw94IiCP6Y01qf+tGOwr07t4iVzTjciFKKMsE7Rr5L
hkIkJ415C6otRtQRnE+TswQLA58FeSQ7v4dNUzxY4tHm+x9VjFDnZxXtVJRUFM21NMMVyRyRCgD7
6M26pKciTtWbSDFI57M9ipdUF9drQphYlnviLfevBrDefyhLk4apcDIJmN8MbgTtOfpg5nckHeKm
yvoqIZqZyFiTzvjM0k0yM74ISOKV4bSBgsvHlb3YNTJLGMwN/Q3qba18XobvKZgQyeeHWorCa/3O
zBlOnEXBydGgsT2SCDfAPZpuUol4PBU+dN0EcRhZWJjlNPlo6xW4DuWf6rV8NKxw1xeBfOroRDNp
tbDGygyTNR6B7rT51OOIn8XXHl9k9Gwcq7uapQagMzLk6RmrfNy+o69pHdarTf1mAORzbbGeaUr2
5iJA120S68nI7MSYuU9hIJAToig0GffSCjOfH2VYlignqGIqg2aAwcqTiA6et3kW6yt6vjRwGbaf
uoPfkTqt1JuPCxpfcgi2Ap8hJZUJoz2pH/JSR7druZj9icyTdSANlYPIo1znr8PKuuxW1Rgw0Um1
/8tzifosy0yqo4/66yxzgHKy3pUdJZ6hT/jfbyCFJ9yMRjqCy2zclfUBRhDE+dWlP4kj9NB+lLYs
ACKoLtsvEhq6Uhwg713SlQEURQo8TlywpwhOAXm/AwJwBx5qftf7Ja8k7u6KvaBZ+vSS6KUsValZ
lTSwQKYRuvXfRthMZ731UgOZ1+IDMhlibe4kMtavx3AR0vvUR23PB55mfv3AaOiWVG2y19cKuC+B
xScbo4ZHyH9wiCjjmeDUGiHjfvO0qkHXMXkwSypa57jnIZ90TFk2NA5SuBCWFSnfvH6AjD7AhXqj
cPxY8dp1R548B98aIkNiSlB3DUET6u78NcKyinLlnKOZ3cvSfcRT9DZGj8uNVqSsKYolroBzPTT6
e0nRLrMmm+7LWrt4/X/YwcVfreN7cNZdM4VhI1pB598HQh0N6GVuN0oS22hiizjHUIbnJX7eDVwh
bxZqC5WUasFHuL9VtOwBYtxxOqmnCffgiclOdERVfRZBKZjnRyB7Ayv4u3iLEau7mFVEAiMbH0/j
l1LRqrQlRt7P5ElSdYTToU4P1PlByxnrJzPGiPxxc1t5ret+R4QHWB+HXozbsMJFjDBA1+tcQANA
hRtrkbGXXEuOq/uDwJnSx+XEkSG9Tzd6jmgu+5F07kz7nuoxkI7cCB//rjMP0IqrEfIWnHat4HZb
ya8JywDSLmVxqt0Vo7DDd32V3X7MlZqvgZlEXbEXFSJg0GYj7eeP/RgCDSjGwgR7D/s/D9a5xEIp
iMpJ/ZA/
`protect end_protected

