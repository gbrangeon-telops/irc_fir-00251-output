

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
e2VQd/JkHeEe4mr54dnWM16g2399v0mhU+1ZT8oWFJUJCdyMu4+q7oH8u3QZmAK8Rcnxp+2SrcpO
m9pYEpjU5g==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
e4k3IaAaNAlNFkvmIoO4qJK1gZoF/VExyr/L2EnpV2zV6AVGzYp83eEX/q7O167vsBLgWYGwRFsP
yi4sfYl5lIuJf2EmeuOEauZwESJuKd6uc1klxaADn7CdEBB8W/rBSaqjDoVCuWxTpK1As0yCX9BZ
RkI2Kfe6mL0Xs6sQpTo=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
IbtPpkhRONJmgAFUIssZ5lSlLGn92JCOk3a/5TU0b+nZGM9b2fJWwwoGbY/OL/gG3eCzPWC2mZ4Q
yQHVXagA0da67WaW3vnZMDAL5frakXXSrA2s87T1FAjqJLmQF7Unh7546PBsqL3OQpKa5tE2Qt9p
EVAvDXDTdLcKhvmEciakrtXwSTthowcA9uRLxUPk8f0EUO4CTfkvluf6ycg5PO6pxfumZFj/0WGs
vgTtbHeVNSCwdx/DPIPQrx/2AfRxSZujtPeD86jE5AaqkaHPmVodviYONlhtWin/aHIYEIBELmjP
OfgBpo4y7pdG2K9gwF+I76hLDXYgXkS1E3SJtA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
jYNHOo/XTSvo0oBfqkgIM6041mVNycidzkShFA7DjL3O3k+3PIOaz1gxN4XAJeVyBTFZGUu9UNpb
lLYIK0sXIcMhzqD/csYXqYD72yk+XSADEYXGdJxFpJfGamCnDtSyBZIo7PBWUINe2Do8h7OVRMiK
aS7bCOSSci8hvDiZE80=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ZHkoK3izETxxNJyR8GdmtFOEPHd8+4rIb//gPmmS/L1BfMiycMWs4JZ0IF56rYeBFqrbQeNtD9Va
BKnGrhYVPTrxcjX5+asuKlu46CBX/iIHEmzrKpr/LAUFIgJgUQFePcXNFNPZEAJsYZmhuSrzc2sY
05sJlmShgR0KVQTbBUWl7mt1DY93aBIhdhmiaHpULcmSxpAU6go9uAbU3jUM00ZMhYA25YYv6AEb
gg84k1+xXW4rmxbK8BWXOVrPImvNZoYgt8qi2fdGpgMvgaoBCq3Rxxbaiti+CXpWZdQ5NbjWArUp
y47h8RokwLA8qG0K8OF44wzHSSkCcalfq4pG0w==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 26336)
`protect data_block
2ypDCeFY3WpAbyUJKBCnTt0IMQgk8i5lhEx7GMe2djRAFZJZ0oT80hnpbnMGVWCd/PtJUlIeQPMW
DImo6DjIRyiOClSwn8sPLN8pRbic9pMGyqou7BrglmybNYXbi6SurdT2fKqjMzF7fFWSZXZ4nq55
ZHsUPW81LBTGeF7n55/nNfGdVYTqRSPQTGDPQG7EMkI3tDsB+0GCG8B2E1vBDY2IjDKzbVwbqa9v
IvnOvbbkc+HoOzLlcgBJTiKvhlnq8/aYnqeGCLUKFLrFwedaBbQIwtbLPG3khsI2HJ6kJCamA1rw
3bswkmQ5FdY9IcBb+8FLjOIvk5UjZUo5Nt5MLXF9MkU5/OVZb3TOuiM8Ma8uEP6lKcihS5HcD8ua
EnfcMHT3x88f96+mYdOnFh+tkMNtqy0HTbD2t5alS53Y0aDJu/zRcfPvrLCtWPi85GlbK6OG8kGo
gREphFmIh6+7cNWVikCnquIIMm7TmyUxV3diaUix4+zoWB8foW/BW48zGziuTrOLd9+VEfUc67OZ
qMB67vW8lLq6EAq4bYTROcL1HPfAeBIQFSJJKsM5oU/xWsD2ArZrXogGaoYThW5KaCMCoeNsPlGi
f2RrHlbrGxg5P8TuMpJMw12LJac7yksowfSoe2x2mFqoij3WYmnG21kd4/A407zhvlAkJTVKMJmT
XtbO9iF6kbGGvQeDKn0FLOQ0p154dp3GaidaUXvD4oLUmCeSId+BZUQCTkGfuEPShCnIv0/JKlqw
lNnpPeCoTrj2h5BhgdSBLB1+GXuiOsgJ/56RJoIBhRUUxqEW248FLvmiW5CU0ObUP7EkzcyPcbFh
TSXTyqqBMItYQNp9LtRFp14wfps40t3uh4SMKAJtl/4IL0hAbnXartT9B2FETMCEGVQYirPJONfv
GrO93VNmuKTNjRtcdRSLQAnxcjq0mUrvk9Ja5e61ImAflHohi4CUCsDE+EuD1icQrJV1YKrvyvwp
5E8/MF/8HcNVP1IjjxNSfmdWGX0V1RK2F2qoTv9pWYJjeVj6L1Q3/wdmTGjZLtSk1VFmy62hS8ND
29p0t7/62L/mYSsn5BQ5PCCVzqMct3FlxwaPdtL3mjMMiB8tJCv+yox31kli95e2EHRse5XLHwCf
xYzIb+yh5672ZyRqLQIU27N2AbkN7aCZwi00unitBAZX9naNx1cFtEj59WR/h2qK/jvUMG+M0oZY
LuQp3JrnbuC9iJ2JLEmx3KmfBdpuSOr9VCY/K27Mw6D0+BnI27ltgFimkBEmIaK4dcdnl6o4lXpW
VpYALiO9FhJyTsHctfUIElAiRF0fOmf0zjJSlWFE9ug5vN67prN8eKbR0ICZXpQ5S1CZ5XBMYe/j
QwhPUkZGweXSr+NqThW+zjAyC9US8hDAIdBefeSda0VxUeG8nWG+flh/MQVymaEGE+K1elr7KTTW
jC3FGHDRoFBo04exdF4hYJVWWRWOD5Bnn8htrHHkU9ocW1nw0CYJmLp2v/Qd4f7GSIFV01QXMd6O
GiChqQ6eeL2swZJO9PEjcGReQNn9rWmzIkPI2lAMl05Jb1EsMImHzZiJi2a8GIkbtwmuxlpm3WRD
OOLM5VOXeoQHHcHeUyHvJeb7e2HKKdM47rpr9LijjWPpDTie6UmX5r171RvtEuOoZFSkKgA69BUV
yPS8VMZ99PN1QP2WjslaH6GGFTf9I+amlfdPZJvMnGYkqIgGzmwMqf7Ba7PzsHSgjHvDFytlxezU
N9Ae7Q1/gKARycihfJlWGGWtnSREjIV57Qp5uwhl1a9bjoUdqbC8TLgCSss4S1avdERYtx+2rPRV
mqlFpnsfjWpLXfN2ia3ImR+IuSBgR+wDBcOwmi7XcDO0hJAznkEt25Ou68RGwvCVGkNXWoX4kSAd
9RgbLbIVLqzrp30RE6kpOOGsqwllZNC2fIiEUflYykt1WI38K4YDosOBxBlmm8m85aIN/eFv3h+7
56epV5jKptQY99T+2OgfAfrSi+A65A1jAvmB2tH6y6g2DPQJOHBsZgX0MnkDoVGGB3kGTJv4BGP/
AffQ6xVE+jetLHFczNaQzp1Pup0ojpDsWfU64zF8vr0XxCG3+U4d7bzrh9h7S07YpvZYzXHeo3hY
CXGWDQIpn13ddY5piMEQ/0c7kxKYiWlFrj1C+ARnq9nSu7oy4277VuKgXTL9uAB5o3m/EUlMKA7H
S94vhN0Q2C1bohILwoyP9CXjIvqDgli/pRNn5BIwQ0QUMKJ//+FU4ceEWiyJRWBiJYEYQYKkyhE3
u58jHXwOAROzssPbpkN6pckmd85LosmCvGF3TqfArz/qVAHXAEUKfwSNuRwcxkpIGmYBuXES1Wyp
ibtxl2GT9R/5mOaqjLwlaaqzgGsTSFomkOdvGZyJfLKMIHIHaSjrXeyQB6jlq9rahmWROMDSIssB
guKVgh+so5c6ISwXZMqT+WGYvSh0ggRji9HQ/g0b3NYeGpm2L9n69gqG4tqoYjQIg5ul4U1+o3ae
6tp23gzG99oMCMoe12LzwWff5AHfTnbNlbuUtaYgvaZ1bOvuee/B4QRK4u32d7BR8Z2wuKSs7j2F
vRhIGJZ1C4cCTPEvcBVh82iEyFUHEU/2NlaWTztmrnmwi8b0zFAiaE5XjuSc95MJeL5XD2Or85af
J15uJB3d+eTfG3I5B7JFR+6LcIDd9pcc8owk2f/XZlBwlzOJK7xW1o5v8ZJNUr16zU767fFmc6pL
ssa6ViohjTvdXzVaSlM02rLLLwTWQJYe2cNDj2xqbYqnBaxx26uRzLvJnJ6nHWAQq7i2ppzq58KW
TUkoiPmUs9VhBUTruOTM6gXeNXidEL+5On9pgsh63obWUj8JJfdogScwdk3Xe+AZNZBIIqFCgpw1
nXJ088OwNGT01Uib5ik/2VxDdCsCiKwqRkky0f8EP8kIcAmrg66I72q3o08e+EVz/sBgeNdFibDk
5RDNrlDRix8AACtkq4pw58qGJC5oI0vlJY+h0483hnRToirFo01UsT9suvJqUR07UZdJOXg8rJ2k
WgV07dh2cUy+KMRGpgVw9ijjNqG/VmzYRMk/gsZY036G/1mGfUqlbFsdvErVmREMi/aKCyuNAXo9
NZSogsqLiswrdxUFS6W27Iukr6qSxwnZWKhXWajnZNVgJH+WAywhZ0e/BbnKY5v5n+c7qfS1StLO
1HfUPI0Jtf0P3H255tz8ErGpV+1sFyg3RZ7yNFFXFoSBpUYIrmIBzhn8MdwcuyiMPtI2Jb29aPhA
ndNqseLBIEWKUD7Bgdzm8YGxFUtSxaYOqj1hgWiJotaYO6owxKZZL9pZZTcSrg36+3cmijFMN64u
LjMEab7v5nosTmyYA/mTYVfoiRfTj965Rmk9xzOcgwSRn6XbDlNKVTEn4Kbb5wU2jo5qF6cjCS/b
Q+YxguVI1TyW9/+D69qALMDgYl6MNaHdSCXbEQvYhbMedixy25OGW+1avIJtzXaF3Ywe6Y+O1d3o
aL5dw0OsYcntnXLqoTLOyBHvABRZI5bNRtskbVDT0PXE2CNB6ZE3RWUn56R0r9AXbROnj3xQBuUM
yIjCx+hQgpJrz7QlE0iw7L4ADTuN941iJUZAliavKnTyHvtqtNcmWAjf4K0Jhfh/94wgSlVGluVe
/gjfJZMHDLO4c4hgfvwP9zcrOECWuViK8hFHSpDcDsp0bT56h7w36Oib4rFf41OYPcNRu1vV80jo
DC2wZysa4LLbY2b2U0ZRHLAnZZv3+3Rg6GLNicLQAqn8ycxq3VGQ/GqTwuZupuv6xK9Z8ZEiBI+e
ZvHMw6dtv622Jtdmt/CDw1uxNv00Ewn8OI6jJujde2HRtWX7QMjaK5RVr7cgWeob/RFgIV6nPDlG
/0SsVNRwfpsNYg/pArnSf5sRwQGzGdSgPlMzJ95943fZBT/g1s4g0DxdqsX8/7FQZ6u92aQgGk40
G1ru+GIUR1S4WbFnIsnTdXItP4hBqKckwcdY9wPPmqZzBMYwI8Zf+XRfeVVPBE36/PQAaLRG0mbA
R5q6qx9MB47HhQxFijgxzZJOs6W5UO4uRCt3nJtISd6yywOLeJDoYJHXDFprhVHaJxm0kh9ykJmM
eFRA/IoX9hUExcEq3TMda8Nd7mOgByg7bPuyF55poFly6LzG/CCGQhoYSmhmnGROQ1BBPKdzyQXy
g4P4q5IM23R9mb1H6y9cWJFWAQD6xS9fre1grId8hrSDeOyc2HGYJynLpuP8UV0NullSfr3NiBTn
aQj8PP4yirlf64smMWBUX9EoKw9ZRvd8zi2b63KzFzD25HYY3mDTwBiR/qUNyoCn4o7vhypYJJa7
k3Ztl1UORDnQXRSB7m6uM3yHVb6Cn7swATn8edKSAnt8jGP07ujCy6TznmD0HCozhH8Lx5yuhJGE
Kzaf9skwe9W/WQ1Vn6BzQSLi1tsrvxrjAOloSc/PPsuJpax3Cu6LLaNnLisDtqUbNxvu5UsS8tE4
RvqN6UgRpMC38J1Xsgi3Vf1FH3MdIIRCaFKs2Z8e4mz8BUFLNeCXZKYERTFN7HaQSMwpkw9e5cQP
8/yQZ/ezHgUsjOlnJoltIhaVrcTsGXi7jAwD4sxe7i335nRRXXaCrjBJ9lMyicoPH65FJGrj0Hqq
rKn02ohvbjIsHZ8rHlvTbWg956HqVxZD5OmCfNCR1B1QEtAtC8BcOZPHGKZ7TczVa3+0t/q6GO81
2q7Bup38492LBqVND8ehYreJ+yqu8oec5gaCcc4XSldMoc5pdb3e1ZdYCnIzxlJG1urEWQ+Fu3DX
p/IyAMqa4C9IOVDyZsW/NyB39fFQ749EZ/6VisMciP9AAyOFzch1WO0Q/N1HGSAKRPpUjC19A57Q
IfzKwafR68RASyijGZ9agP8Tip2AJ8+A+JvXC/T7BVsPe8SOwA0H1mzLdWLhLSR5VMkAfljK23dN
56fKy09X+tLadFXEgi5PjzMuHzqzSnSU9kWS0AG2Ipoh8gLWtgQXviJVh9Jy24CMBuF8qXzD4UeL
BTp9CyTI7M+Jg5c81kI5p/Buv3HrblTi6t1/RXQln25OGtzLIAiCGbSkpqB33AX1x6OiE86AuMCV
jRjO1LFAS16J78WdT3bXUN/eojVNf2M8wG8Nt7yaMlr0B2Y+aC605w2KIecFvX6sWOc1IkpzJD3E
gYuKOMT/D4iZ25oPHYZVp4TQBt6s3JlFYVdBDRJecHPLNtJRIj3C9TWWZnlymh4eisfXyoeAAQVw
UPzJKW0xHtR/Orr6Bi91EXRAQtDTE+KXzksBn/D5yGvcTdG7UCY4TCxOqbYDX3FpgvDpJyAVMVh4
5qnSMEhZNNVod2+ivC2g7yq4vyd7ddqIAGExAirGn2mHF/vnYdgX9yh2AgjzjRB1kO25sk1JUxGl
ZY0l/XonaICLOeoqJJEMv1I7hgNu2lX2rXawsUvE9PtF8SEeCCc3C9cV+Iqkeyd/KLa2L7HtAtOe
KgUA/OF8tXoW3RsZU3Yis+4G0lwNsjCiuobaNrGMwgwkAvuevSidfmnypX9n7PHyEB2EO6kVIzPC
EdqLlOcvwQRUBkAfhJfqnWqSThDa0ClfKK557dD30LvzK1wRuWYH1gs5Y0IpsnM7bT+l6XhIa198
bVv3q7G9Xknc0C0zc5B8ouwTptu/JZY5X8pI8e/qTEm1nm1dgUiCsy7W01t/eKNsZIRN+QSX+xSY
WtSErI21cZIFuHkO/1uangw61npCy/IWiPpZwiePsDcDMpScNoQIHjFYPRQpJxqHxcwQurAK4vD0
O2R4X2PMAS8asq4/aCUYSPOP8rSH4XEEQm+wM7HB3MAVD3CcmLCs8hVdpRO+wF2koAkbU14fCkaZ
esrSUdNK7krJ32jvNGmn9ist9zvzZNYsiZlB4DeWC7d9+FaZLOK3dnctRcpAf1WBxK8O1NtAQmJ5
CbWWBajH3aD7zUvKnttE0+NAp86OKmBxtVYaihAiqRVZiDqI6/3RED6VTDFwigymneG3fPvRvvEf
nLwSnO4obGrnMwvVkhrTpxYO0PYHzOVhq4lqwFS2E4B4NvKjZkjGA9FNxqB/cLFEVPY95UyCbIIN
kAgsdKedjK2qwQ9VHOTWKD1xsxY+TJM2s4On4dTkmtmT27BS81sgZM1OMZJCSSIm7Um3/Z9if6P/
O0jJFQG01lrVr2TF7c7mKCR2vFPkt7QrNoF5+/4bd9APKRGh5uxN8G6XnXoF+L8RWJK6k05V06Mz
RoeWP5LkT3vKssUZQeIoeIHd260WVhYjob5p1U50kdOMEFr+Z76p0bXpcEsRIgKuBlRhq8Q4IiDQ
QzoJxObk06GMxigavVjv12fouAGKcM1NtMVW76j6HDuCMh1DLCA4VrLdwYl90/v2AzVHnkRt4jg2
GSrURyFEtoQNsPGgbzaqmXvHX/cdKePqni4PV/S3qLP3weC4jlXYRCkxLPXy4p+pR60EpMeQhDQI
Nc7uNrxOLVUNBOvchPnW0QM3s/BvTURTqjDIh06ZfNUIUZR0b7Jm/L1fJ8l+EjMCWAV1bkZoPtbA
eiV4uuCQ76seJUjObsp7YVJOfOynxsA+1d4GBTGEbZzqDw2b/PzSA7wJRd7mC9jXgqbi/oZLymFf
LQlVI6zg3Wasi5fdMUzJAEsPz9b2ZxZO/b7Av1hQr1pso7Sh1/PPoIcK31gUQZYZBvzNW1xPecf5
rYR/u6R0iA5UGzmwcjvm/YS+ORXqaWmKfrfs28mXLxuXsydNjsjr5IIU8Od4ntfNvdt/1Uzsei+P
clux2zWmpKKlWKfzdD97eXYnTmaVUoaE/0/kIxNHz/9NOjIf9hWw2TucMp8LbCtO6qNvEBSxsbUA
+p+/u070PsdRdxSqL43F6hpRy9twoWgqPsAzYn1WzyWV/i/0VNo+8ZhcCIym8By8sO6tWL3QVfxQ
r1ss0KTba9nlpSUvifRE4XCo2pzSVVBlS45MNc90ppEI38OupUDyIHgqIjBY3WcUjUQ5KbSjKBNj
7JVJ/xN04eU+gmsLGBahjUWXXSlcAQCriVEf/6I1NxHzlG809ublBEXadW62wmsMNKa9z37KUfYl
NYLhJD3LVMnsNEJ1aDHjyGFtuHRBEQ/HMjyuMCvKXec4wcFUSv6MdNu+gXUiyZORtsKScaZ3Dq45
Q0mKLAaviBy/xcsiSHLh2q84jDIdsI/qx/KH0S+IevEXitOaTp9aRlMTLaCjN9+PSYJzRSvV1lhe
0Wsj1bYuO18VIbzoV3UjjU4AT8qoaP9c7fajDT92UZupBLAYxp2t6SWnGFkPyeNZ6Hl71lOmZq19
9Td6Wsvdiiq6D9TcgAt/RXvpqSPEDHsaGs+OooZY4JL7izKfs/H/T50QyhJFbUHFQKPhi3nhZbx1
1e8eNRv/yPstZsJmniaQCeV1TaO9ZTk/TR7Z26Rhy93DA3X3MXNcC4x74gK+XvYoj7/r5btNyBMs
1M+jWeeM4rOTTf6m4Uweht68jEhknx3PrKrWzqhWXChKmn/WE8zuW9dMLuEmW+67l3yE/kBw2twz
HknGc5acyfEXOVjiV8dUWHfJM8VZmUrU7snr8xorUHVDCGqeN7JSYrTJXFL4xOItyUMeC2PwLtya
l7mUSQdIykct4QudFItRxmylxtydI3KvcABqJry1WYNzrxVjoFgW3j+FwTLqAsKcPmss5WnncBuP
++v+YGagxl+6uwCA4jKE2u7Qxr2L3sXBSkizsn5rZ7sF3XadRrh3u02FU6weIQSTy8QWbGatZMkb
tstsbbzdruubrsWWQ5fi73xs2xZO17FtJRP4cxsppGkpw3XXIUTpeLhXF4nvW+YYEXCf1eHi9sWE
qmI0Os56Y6ixVwDgUjcXPPm7bXzZ9j4Kl27IYoFQQAxZ+NA/7/9p3p9Cg50E3lR9FujNnknfIhxf
EuBJwF0GRrv0Aq7XcVh+puIVAzbR+KPpv9MBTjGOwL+n2H0rLsdfCMULHOGcRnuPsKHYbpLPDDSZ
OBd/ZaU8cFPvw2SwjbvpzhKfQaPLI6/nVo0RhUVuXLRYXwo3+6gE9oci9auZIqbxCcVHPK3KX+Dg
HgYLF1VgO6B0XsqLVeQrnZTKxqs0pcKdwMRabjA1miP/wh1+Grdx7xXGJxjMg2Ykbt9NML6M53GR
yyEsogwWUihaVFw8NtDqiRe33F63nUnCFbPmBGNdAbw2vsPKdZ4CRQ7F95aHnu6Wd9S6IT8NQN1y
2xZmwsh46Infxj8swc3/mZzwWcvcamkDPxxRCDaK2TE5Om1ogx7ZXVcx5oCKLnXIMB4pW2j9O4yw
Bja6dGtUtRfeC56U1KblhUnnz6qJmEF7NWPafbsOKcqUFPSA0iK+Ky+hrhVyuWERrew6mBVuChN1
wiXQgnoY6KdEhc44iGQFezQli/V+f7r8W6DO/6eBEsXEd+E4E8FpO0mV7eKNbt6r1rrlCT0K0dCV
mMJqHX88DnmGLi0/An5ydOkdYUfotwf3VpZl3nVUjznZjvBVrG61LoSt6J9kHKa6XaMX1lYym5l9
igDgcrXGvvRZgq7tlJjSWlB6m/TjZ4PSEAECdjYjcncuEIPq9LnkJ0XL0FgDV1O6HHc+YqKkLPvd
NK4OjAWH6SKJZBh1Zy/5dNfBaagQPaZ3zioAV79uSj6Qey+VcSdHo0X6ygRScosB1aVcjl1AVvJR
y+EcdLuGskLddIBXpCVB8uL8Sx3qiticogX0yOPro14hXFFbj1GSV1fBtgi5YZZYfQbLO6Swnbaw
acDF9WkIdYIpaQwYefMQ6m33vQF/W5lUx8loGCGym5lAD8w1yw8dbxWK34BcM2X+Dt50PXcG3Whw
0YAtrduvNhdbdkk7UEhZ8rKstsaOxg2F0q+SPxltVTePp4OR8njm/Nte4AHqvb1VUb5B/MFwig6i
TwHlzEqwtnWTA72i2PSUmSjrH7SbeyYdYaxLVbV4kUCiou0ZqGow3ZQptLO6wMQxmJTVKUNhdrFg
KRGgUmP5Jug62MVk8hDcfJk/m3zoNcq91ZIXXtCkQq2OEbqNXUKCmjHtOXTvF4zNHv9LCron3qrU
6eZY+YpBFB1S2ej2OYMsHiHB7V0EWajFbPqA0a/xJghRXFU1idvoCQGs8hHj4LW61CC3ohUuhUGQ
2XKyuGaUr6pEFFnVDVFCyvhIoZUtOMtkp6LhrnXeHT5Sit14NOy+y1Q3Zw/4xvjOsrcqLjkMV1j2
sC07NuMVAtv8dkpkPky4+NoTj2eeLw9MGYAf6wosPAhY/cgJzWPdJp2LDQm1uWA0bhSgkFhCglhY
IVBCXMFfIXw2ZOK3InDsAfglLT7vy3O/auJCkiosVjrd+5jbmc4cwQU1GODseQ24h1qLNBY1Lhhc
dnWg9YwrE2vM2Jf+XJPjjgia2J1LTuWimQxgDQyUH5ZiVJ0nDQZaQNEUqDvBgInpG7ipQnXCrzGV
aI2GtO216rXykaCQeqnII2NI5VD5wIKhkJjmSjmlSX1DHk961vG1X2Z4jX+49Mp7DHWY7MB9Ninl
pIeF1/ois862+3hecf1+gLDc3cQkfP2x4nGJu8DXPgAqC/w7Jcx4q2U2CAIhEkea7++s6EW0wm32
/Kc7lv2mhiiPE5GK4efYaIctDiPYC9RFhqkFJzLdWIQ8Q00vlGH728L3k6ibzonuUya2zj9UT6r4
ldwXLWQEWkUGTM3TT97j99RkscstGhtj9dxfj6hdWD1MJB6O9hts3mDF7+SDD1V+Yef6RE6ah/U8
M+9X3aRXdOv2xDi7/krrCbyHO1xvj8ESTVnv3BI4a39pboETRFg2Dd0RMZ5m7jzLZLHbRH/ZOnap
G1BPWNM8+gLlyPOkWuHKjyQ9UoA4ICtghFZm0/gVqrdqvqiDNL1vaDsEptn3WpHVY5GM3iBpNNNW
cA0VCenVu6LrBCC9B1/0GbtsrQweF3gEpvcg1RSi8LZEaw0aZMk38RKPMGGpMTlIQWOXVwXivWZp
4cripuvMt1qOfZ1gWeHW/JZvN9VXPP0AOp6VvtmkHWA04CW3I7xNlMUbVgkXH7dMYQzNbPoRalxi
5tLbz7Lg+UxeKQemnL2ObxZsf/1A2DY138XgdR4vkZbLs/ZGHHtXrCtIeiPlxOXvEr2vRI4Kaanx
Z+xNPStlRe7wKJo9y2sUH3grFG4HEjyzgeqAcC9xArPxxB0Jq/mgmP5tTy0cIqFQShMR94eOwmqE
Cha1g/n15XyOedn/W2ubQKdhpx8UgsGt2YBrlbqH2au7MtqoMcueUsKDiNkVIXr/AsdPtvhhCvyD
YEUfQU8ucha9u357cI0FaKrPJh9lD0oQaGtxRO589hTgrKx67hbpHNFaPUhGR4bfwM+RDbgrfCEh
HdzZiqcNcnPrDaT1hBPFolQRbZp0yR94AJ0BytIs8SSbNhuApqm+lFP6HwJeRI/J6gABAGwpur7W
0Ebw95SEI4dTEgehmEkcky0NIsGJ6DD/Fai14luKwaTSXSMeI4XM4kfJS4kBHOH3osXz4lqtgqfq
8xE8FJzxl+Ifx+iDNDDijfMXXWzP+tH7ADkiiVNwAwAa1pDwpcM9goclUDmOHGbO8RbbB4iM7Plx
gzc3DKu6twl3BWe4Fqbc8gr2b4ZKUOyiEfuK76+CHuQonCS8UVPkBzTh8fP6TnaNqSgAPQY4H0yA
9SY/qm0mRfFBQ8Kbm4y9Xe9cSUNSdMsnjb9WAKQjno0wcX0z/Jvrpe7WN8rop/hdcr7l7kjXZG7x
UBA75814PF7qwgczjLzTP95yPo1owY1kRkmbPEnrvMfuq2x9Te0YVensXI+QiOxRG9CKzU3a+uzg
pe/HGHyog8yF9GyXTkvseg77lsHMj69h58zbfV/AfPJ6VfJVbaE5+KcIiyxXYcFIr7xJQcRZJTSt
canLtygDmTyOFz0cwDu5mJQVn1fvFkuwmGeOzu5vG/tvQpIeJ1HfFsxcX5judSqYPQd2W55sQrPD
BLHxx8s3NvxwuN52AbpiJmKW791miWP9BI0qWc8V3FOE4qqKGZ+k6+zas8cZ3Z39WUsSBKQwJraW
bPbyPp7w4U/gYpKJ6/EA1tSlJ6BHi8oLGlZqXHujpoIhryubWQdg44KeqIFZs3VJJWWj6P0th9Ul
jwWr6r0TcK/2Z04KmPEEHDd+zjwAvsRHHmlOQAt32T98FLufHEnmz/B7laSNOJ+i+EXNpqKIxxRi
XapdUKXn1vV+oY2X2Pw0PI1gzfZj6xO9GIEGQuQoTCUSiqla1sbEB+EPa9ZCOuDNbTmfoKQfMR1j
GsDDVSau5jv7I0RXtPE2EIxr7ZyAgxe+4hCLyqOMRbQj0XnDTGOK3jgIdTvlX+Q6NjpJVYIZaAlb
fFx8sSBJM1Maqu/WOOUXmjibRxz6seIvtihpQBTjVR1alHGyb1a2HqUU2qS0e1P43oy6ef6RjhNb
xvQddkLTkgjoeLEyrKelVN73e73mk7vGF+2a2e3CsTz5aAM3o0myIw3JYpbCGsiVuP37AuJrcbiH
yC/0/J3aTd5wZ6sBoUsi+BEDNg/11XPOt0nPE6a5YqPUhC5pqUY4Tj01TRVFJ2mYBD1NBzY5UXQ/
Dfjap0OyZxpoiXTObzbnZ1+tNCH/HRbXtprG1Bbu6VpBjYlaKHQDpVkWKOvndRDWZuABkFc7kAVb
vhltk6fXVVN/V0yt1HiOQmpjAo/2Cf39oe5BqvgxLhff5EJAVxAyGCAyhNM5ZdQuysR/X+whaHnv
YcJ4bFY2mXsDhXAIllyJ8Slo9N7Z3e8JW9tIh+hWmDq54EPvHKuwh4vdWnf5yvNWBbFnxjOV00Mx
rhNTpM9fU6cJSzNBWo0Dj7Ch5hwNGIg/OzbjVyE57XLeqoUy00MtMIGpXEK/TEOnywWOK7aMKGIC
ODGm9yEbbLVGH/hxZF3p5C8qE0Muzk7jeYqGZ3RVS07m5afbQPSTdeVHNcv5p7kmLID9SAEUZpdn
7NH/G0SqFTL7A5FLc7fODWtAMFfNwln2ntRqj2fmfdgTn+QthZAO6moHwPWWLT3YCHxHq31fS9RX
jKsOE1et6zfnS4Da8MAZtujvyegOnTT2obX751+udSRExzZkD8xMmhAp8FY5Af0Ymb6nxAGeIEoU
2Kz4grqL3uOfkm0xk3tf2FLwgI+3CUjC+jv0rFzNWN2CMP+qCOdnqt9f4grbVuEzCXS3nN+UJbmV
4eESoNJki7sBz3411K3Z4StGowLWUuJ9njTT8vbWIrZsJpXzjCwYI/iTYSPqwIB8psPh1X8a3ncw
yfaHsYvShu3bimN7tSnafrSrGK627vNBhBNVOgF8DAQ4YZDdd7rA+Y8atLxpEIg+lovp8+hKQd94
CA/ouzfSMBjp+NEpjW6LvKisWEtPvisOBYmo3zvhszxkHZgVHPQ7kjEL0PkJbIDZEs0HTKiEV+p+
UvE/I08WkOl0MQwRsdWoCoGIDMR64jitYcfK4xt80KokQLW/p/5hQ4ROd3RsGExixDiRIY8YPGlm
EdKxC/KUFTFNGtDkVe/sd8kT8yoWWHxOzqeX93reiGZ6g2EscSup4ZHmxEjV5z2GmFWXNPZjRYMF
1an8wN91290cGMlVLab33+nm67wMbPqgDJNr/q71nP266WUOBh0f8RL3X0cRp1InEeveFWIqdhFN
9DpokVKrnEJozJBxg1/8qPmrCzXEVvAE4eMfViTpmalJhGS2dQ8t1DH2hoNX8N8iyXI4IxdVjxEV
L7/VWLiCH2frp3STKIQUD1DGTBYMRf3gyqbFtLXWAxeKqZHbqmDThT8SXu4xktQu6xHMZCURaGRH
RF1K3WyAqMYjmXV+hCRxRdOdVnOgontNthSgpGr55LvgrRYykQVn6OQRSW7+1x8gZsqr0GYVQzfN
5SY6eWhR/srGnDOvKXudJuq2oeHqiL3X5/YtC9+GhRX8vs/rh576FRirHgMlh6ZtaPENhG6im4Rj
Bq02rusZS5dagqnEiNArPcEbt+x67CKB6zH2c7fmPKskCvi47paphPGVG1LIVKVAfMN17I8vmMvE
c1LY1NwkWHK2TIiPRXRFGsReTHEzSCeyMcWPUfg3q2+GAbPdv0xx9U3t0q58a4xJWsAvsWicpnnI
9fz1gjm+iu3acgx6wv4H7JWmRxJHU5DwOOkfB7rcgGBrgEq5C6vYtuuvklg8tmr8/gpyyu8jOtsr
/bAWXjdpA0PfpimD0ZTFMBTzxD7frjjbJ5v0mj8s3fAW0+SR18sbHAH+WlsC3la+q3HTVGtRBLO2
Mvv62LENojRiti1RwGeu7LAqYia/gtqnpw0ZY7lrjsdymJLoQrDinapXL3RZ+FEkKv9T9t6hl5NM
MgG/pxGOwUQYLN8MHiSk2/6Lgd5Pa5CVLFu4s0pczszV38083gpoE3bNtTDqReQAxvsDLshHohzV
IfTKULzF+EnpaxoO4R0icKUUarwGYrrtK9/8O3PbGpBtT0h+x1UgBPvK5SPFGR19PF3m/+zawXyN
ylCC90Vm7jzOsUHrf7XzdNeVk5DwkXi8CA1Eb1zpqf+eKDqbQ0QI+mq2vOpn/MEM9IKh8pwG6m36
kkQOHidv+NVjVxB9GB1lcsVvTrAUJ+9DbV6uRE9U43Ku5INI3LQY9/Nd+D83MCuda617n18LchFY
hmYPkC+Wm2SWZHsIu8hQSKJJVkr4dChLrCA+A71D92ilTP5EcR+msH4xr8xFOJ+kghDAxCdaGD8d
xt4i4LYGD/5cYkKe6fauhS1Q7PWRwe0VGG8cH6ChFnwDAEgnvNb7JZ735dN6fHiQDmXLWT7xc1Gi
Z33TTS/A3V/c2CsxemkYy4W7FftzbrurpWsgRimBJikEc/26ROM14eiS5pBzC/8Do+JEIJCeNI4x
DwHvWPq9vy+SlgdRbehd/UAkaPu49YUMhGQnsELVW6vM0SjBsBD/dumuK3cZPPffOEgKNia5eaOH
6QkrLW/s+h67wT5jyXa/zLj8VnV3L6mnm27+JR68iwVq0f2VS7GtE31D4OvSxarAFdz0wqrGnF0n
WtzBMsGnibSLXdtmAJRJyXxxLx0fEfuS3diGW+EAmPXoXy2WIALMNtQirvBh/X4huqrJxX5w6Kzf
E9yfLUWjdhFkf1ZtpEckbvTAjNaUkBfSF20hnChj7TSRpLUl6CsVH7sU9wTHPDo6xrVZ52fa/Luz
BUrELfiAHKQrigG8Ug7ANKiKxLqqnbWB+Sfj6utxp8HWLXrEkOHXnljmcL8JxbNkSrs1Xg0TiDY6
GXdE3gGDkuZD6LpWyK9Yv1jvp7EnGen4dEWKe5k7lfknX8YXDjbyE4zHTM3yDx0gNszrhVq00H9Y
5EOZq3mBnlvpdwPi7F/V/RGG5LPvOH04ymsa6zukIUCkwRKo7OmQjXZRk9qZyNTmHJITDEvXD53b
bgiWkbWbDH9qAym5X9Pm+0zsYVy52qcryPcvmyJJHgGGKgyYVfNpZSiPSxfKCv29yam0wt1dZjEy
huHOfRPhZI+MGn/o7oj7LkqY5K9PQ9T9YFRCgTX5232Lh779raLe+/8Wsd2J+jPpXJtGvcwWl9Rz
2/aAbDSS02HMUyG2o2S3dtS6Ba1iRbm8C1wbjtFdQO9yq39ned2OgIHGvSqPCYnR7RUsOVPR2qQ9
yOzPtkKKTI3GTQTW2ldZa1iUOLLMmxAnRgI/NScR/qEK5hpCbTYSeEfleFnbBrx99HAYf/UBavGO
wssUVJ7dr7KzxcV4pXXwyBXTrBBGCxQEByJBucFvr3I0R18XhJ3CDxEmZDJejdqE4SI33mv7EJvY
g2FXlf0WIDkVV5rmDT95o7wHg47TE+c92uh5Y/CZg1eomc6RzNDHqoQFg1r64N+98GBEaSmRaw7s
oRy/+U8ajYzJcAskWpnzDa3jqtkM33uEY79UToFidpK+QohokIOV7hpD1tpjvsHOjmMeSbehn86b
MNXZk9ZBmEMAcyM1gsFVn//VHBoDcogiVMJcj6Sl/xofg1rH8x+iiGL6UyY0FkSK2MJFXq/9Ekin
10BpMIKX6h3KGKRjZw7glEQX9/8LZ6SDu1FmBVEB7Brd7CVOxSTCcgKgbGCOZDecw5FIL3mPZfuz
1m96CygsOLkdY4zBJg9N9hJsc8IqL0bgQq1UfgEKHCylQYqDOhK522DsZ+UUqYvAlyU3v85LldQS
NL3ZoXsYsKcIvHJZNPWOkSTMrNSkmBgemj94MdAQCJ/czDbfiwfvP1bSAmIaRzsZ5QJuuG94nJLP
tXtF17KMf6WW9yEr2l9w6ZFnnHtaI/PP40SaDqX60l+wirjFspkoUjy5l1Nph9zbd/DmzQSZ+f9L
8rDDuvfp2+RhSqAPHAs0FcWBMZEAul03484sfEdFAXbZJycuzuZpKLbMv7bCxVktd/lOvddsD96g
5NGf4pBioLNG2qHTGB51PGGQDVUeoJNKk4/EY3ewg2RQ6rTqMjVhe4g2CxRQDECNexi+Baoc9NJC
b3vfYz5HncEue5tfIpqlwOYGGMAmhdLBhJ+Sea8ZhGLSZW5whCkLQJ9cA0MzTHqQCijNw8dvtmBG
2Q6/OVEBzjT7cy7AHsZdWCzOQZnnT5E+/52tiXRAX8S6/z1seS2Dp9xbyIDQwDHSTsUtULe8fqv+
UwjhTH8fgeafw8s9VCkhOpXz8gg8VqDatT0r2QOWHVH9kTIe1aqg+y+EeuuVwcc3z/l5mJAahPhM
ck1l30cuDtKnisdmGCJ0COhPsH1LeHUVq2jKIsIiq2MN8SLERg1CFTYCFPlIMmutayx2Kdab8OyV
yHp/Bj5vyVV2cj6cqp42EVlJ6rYEtKRQrsIhEuMDjAm9jpRDnYUVLV+I5A+9NZ85z9bPWfFATG/V
mqsWLajcF2t10svm2n8qV2amF0daATmiR2S/ayhD3KkZxrl833u3yk9TaKiSNSZt73QJh28jjJMc
x90A/GgagncPCC40hEDKCJwzXCmJSDX5qJF1vfhGKpu0rCztqXtqSAXGBmTCECZTxSTFkkmb8wOY
PmqlFd5qPQZp50XT9RUYxoIwjwnQDU3hh/DnjG3jFH0ennnVFJvStwbN11iaoEx5kkbi3R/Y0QVJ
gtgKV3kgahqN2Fodi/TfxhiiIGSavblgvdw8IBkSF5OOcaPp3Rzzcq6PhqrimODtdObjJj5NXAfC
JUnCBhJbWRrDaTDsMWwmYkRobQ4xB2BD6Gwy7ITI7+4GWtfJuZbf2n5jhViRi7tf2FZv3gn3cLlb
fWatlym0INbFQczMyNHnxOFfHGINr4X/XwHxzH5iv8TO9QHdOw3NM7Ea4dD+d9dYhs+2h/aWe83g
EleAgTR+J33fH7qezHUFDbJjlvnGwi9heAGbha27SQiV2DFD0pUKbSMnXL6lo15aZmWWIeFvaU0g
wnsIY9mP5/xJZBXlBT9uWEg5Z2D14UiL7rEMgn4HZAAXngn9HI/69H/QeFEz2vRafN7HeMUgtMPh
whXCxUPELR+LVloC6cf9DLLMMyYAIMKCXjGDB4ThOv7pMyvc6G92jo1UzI1GKSAQaTIQmDW/UzkQ
NCHs1Uk6IOeEK/rH+upw6tLJP7TAVl+mazfU/s+ri5VAK3FLWemMJSW6mWtkVl8CtdiGD7ddf+0+
WW7SzSEmGiryPCibaGVLZwuMHL4uBYGo3nUynhuqVzlmvokuRdKv1QVbgPwtLPA2wIZCXF18GtBD
hFvKqGpzCnZcXThMBmP7KpccqZwb8lSh4AD/xOa1xOKriwqm7mrsNzTEYyjx1/YhydQM/gf4oTDj
hZTFmhWOuz6hDBJRBg6spf2xpFYzSS/PPjxXqeVqYQ+M3kSs1ygjoSHFaIJkdx0/YeN9QU5I1JbI
+YSyN2m8932pqlZL0EMWoZYyjVSiggTF6BuZBWdxFuNE9/fYPY3aK1SV9mDo37ccicBnXgPRVJfs
ONZnj0E4uNBUCfKBk2siUwH0IY8RkvG1KMCzk4zkpt6jtdfLs342JYiz/7YrrN+N2vNQXasYB8Xu
zqp0z1EBs3MvpGhqN5zkMbRBa1AMPR5bgiqx6oXTF3mMOr0fioKfN2PX0rIphH3yojPIcj8RKwEK
a6xexIaqCnWGDY9nRbJ3+CJ9dTSH6coUx1oh+GP3TJ5ci8b6ZQUiPAtoiR2/olXPWHwBNvyG7xEe
RBfo7r1BK+BxWiwyn8gIGR11vNrB5V8JR1xNJ2oKZotv2b/AyOO9MkcdWtBfxhpGHygXdaCrJ5qu
DWhu1zxKYnmRbIOPfc7s45Sa3DBFBxHuleBbWADeAYxobTPsvkhvhyECJClWYOJGzeGfyfM7qPWm
cXVSHPp0HMQk8xaK0RvEzXbyI8SPzZ20+pFiI1aAzcV4QERmGD988qQdCBudIJkmqC8Es6gvLK8r
aA0q+eFCPjT/HtPUTYnbqjsrqqG2o670+0reGyG4eDtS2mqlvpS4haDWc6dsRqfKG5NooOmu3fJk
lXsT+zs5dSjS6Z8jSkZfiWn5r4ySNacnFakyyq6GvpMMHx0oGFBy/EenYanGv9yCFdT/H5vJ5/jy
hoZxFuvcZ6m1Xnn/xA5lOgEgWyy2t99VFVygsiB/yx8KOpbDjGWR67/YS5HUN7AcgWRsT1nUf7pS
fOKFmu3qHaAihqx0eQt7YCLFJx5+jBc8jqM16+XAje//R3RSKWoV3hCey1lFCu27TQTcvuYvoqCR
7kF78H4biInB4lzliV2IFSvX06n7QmOhzuHvgBymVRCx7gOjxmxNXOkMfozsvjoz99kkgyf8aBY5
c/25C22CaPPLpx9eJaO5pqQg7xsh7+oEDcxnbU/Oo5leg82hC7r6846hfNYoRp7qQ4w6qqYw/cLj
PZd9rBkNXjZTcEs+NZILIRG2IE7re1iDrj13plcVe5Tbyy5TzjTgbzjd23FApBR5Gi3z1m47PBGf
1JfFuu4jco8XAfk5FyOSQKeuOBE3Htbz/pPY1CYroX26dORqUaJwjcdTGZ5iyjyP94PC3Nl8LCal
yZSoEn4SsFrAdaBV+j3mc3zqHWFPxv6m0CwqqoPFeR2tlSg3YgK/JU/tCIdOrkKpKdEKb8PpFRkL
wj2FSgAM/j8FdSoP0AaYjCls5whhjMfytg/DnY7qQiJTiBJzzCDY36q2yWxkrMz4aatUeI16yKWK
BhHUc8ylgO49h6qJn89MoD0ryQ/ZsZiusXZt+Aq8pVcEVSWPiUkhvAy2ipJ0tjLIe0w/atHvRu7q
EZa50hAry7GPZHvdcRVzLceH8cjGk7VSOLTxr3f+btN7v6oaf0Abv2A/3BRC4ACP8wtcXjYKCKW+
+AunSohThVnMazYsTiqR/Hj2MzcDESvlck3L9k4pz7nrj4+d+NWoBqqF5nn+EiozoA6qhq8YOw1D
ejqy3I2+OPOSW8m2E1MaojEqZ7QsjFSjkqIGS2zoohMRmD62y31cMnJp16vkCP2i4DTk8RZmUW2b
XLe7f8R+TIVrhNFH0o/wg++Z1BzCPMLmOACC21xka05NmnahVU0c99CWsWapi3LCgOt9XVId+xaP
YxMod3wNS6XFWSCAi/iF+DjG5XiTSREHmnK3FoTRCag1jN9Yjgz68uCst6b0UDhaujMa6TIUO5/j
onJnzdnM+a0U17R7st0RYVzNaI1+4jXbwGYkBsxzSyM/muoxWniZ9dk3aYgbZcayPzRj0rrtlZL4
OJIhGtf5jFmRUuxPvm5ZOl3DVtwQLn8IzmC5jfAopRcsqsAlmfQ7UCbHFe6fPMmZr4BtrSiO7cAD
wokqg60b7geWsFZ29cXVfjv9mObuyrvFW+DqxR+HPlPzBG4NsQzN4HNNV0/tgXX7p2/212enXZw6
uhbiWsa0rgOLY9ouKuXH9lJ7pLtprEKR0VkIisxHlMHmE5W9eYIRR9l5GWZughwC8YFsS9gddIXF
IYVITIkxMzg3vfoV7CTCO8w8E5yblI/7hDkD8QqY5FVZf2Jq8F5xlyHA5DMCf/hoaWsCOVrscgcA
DbVgoKXtoRbOIo60AZhfJmXuRfZVIojz1A+HBbEECpOc/1E7RpormHFGEIprYCs/aCixvk9n7mQi
80F1Z77gfId0ORZ6IHuu9MX00z0DiEr/AslLE8ICqZ+TD7zGYxopITLZ+d87G6OIwN99HHrGPovo
aoj5wJE+B9LlKJaOgz8t1zeIDliH4ngEZDyP4xWNL2tILRvkapyO47+C1+HcgoIXCoGFq4KRKwmc
ElHLi3WpHt8epBAwdPXKQ57zvDYnXOJK4VaHeO2zUqmtD75uTEzkb6O6nSZpZwLDJrY7LsI8MZtX
QjXvcjTg+Q9ghV3XXTSnpNbNKmkzCEF2ZAg6olgqEtUPFXps41KX6lAo1MIgB00qSsKUF8C8gyJL
adpDzRgIH2wn49ucLh5eTnwEL4uso/DQ1ftMNkAf0DRYYKS5IP40o03UwdXhqXidhyz+NqjR9lMu
bO8h0dqHDlbBTJmJA4YkhFQR+wxgUcwXHbbZ60g6UQC1+ykw/sWxpkClCSB4vcWjC8Sm/RLX9cVJ
kyFUKr3E9N7uVwQo2heHbNG8z3QB0YpVOUma8nO0eED0djYiwHk6jFFTRxv6+r5rGCcZorFKmUFW
Z4+FMmnjbT7ySX0vqRvA20Xz7r9mcYYgca6n7XNLEq+v1Kx4nGXTFi85nvyfEbTRPE0Q9U8meWTw
6UpQb4cce50CqBA0kZviajnw1n3KXy6YXAZ4U/mdiNYXnHX9ndKwJkFqT8xT2Wo77CGrAC5/Mfkl
cR+aLvafDbnnsWRm/bk4CDYwD6NJSRpN57qod68HdWrS7ZGT0OhO/tWwJqnbldewQEvnoOtT9xIR
BcWDT4yHrLhZwguakJigEkq+kYQi1DOFK2HvOw2fAIywaZN00x5N7N4nIE1Ge/QyHaFjXL7FcZbX
WU67l22aPXUft0w4ehIH0a2YItd9wf56FNkW3T2hu0rYTwEBNT7RGpqHk2lnwbkrkaCU6xVgLRsL
qyypbg72VlgZ48TqUkGyPoov5lzWvj+SpShSPvWTIi0vttCJq7ptFsRnvUPoFCH/omcln3oAnH8S
d164goYgDCBUi6Y/iirHpkjd9BoqFH7Wbe53s9pGecArFFVXuHxZUoMKqz2OIRmYZx8qEK55qHtw
KvzJXqsBLXK07FQmqy8NilgH+uRM2vLY61Ye8DUFN+Hoc/2n5/D7Kk0tCFUtE2cGcdnpARuDbg/a
65MdtXPSik5DVGJlnj4kHJZ6ejnPoQeMr2uGhAiJDNzzcAyOxMmZuG6VnkwyTJoa10VazRPeJCB8
fYPl7zBmIerHI4mDlYyCcEltJwOBgc+2ky9JBc6pvjd2mTo02/zMIdOddUsXnyLw13mKwPh1QMuX
UTU085bMr5AlD1n82sdE+A4dTIUWSZ3yQEB/KkxuNuMkzajHIAuS205R4WnFC7YqhIbLC5H41eSW
nb960mQcgeh475UTXtKsrQ/bEgXmZ4OdmRAunV1ZIbz8Cx4cqL8mzIS5g7DP86N6brL88TuA6reP
Y5lrI3O+01+Ibd1eMdS2+K702QKThY+kqzyrCiM5IWPVsiTaNoSVbiXXcn4tPiGNbRsO9BydISt0
loT7VnPE6X8jvjIMjEiN15LBs/oYpQvKBEEwxWglItLZoYeLr+8vh10PIIKgfXlC9UTamAqsLUEE
qNzKvljTyzdAP4jaQls5WEckVNK06jmNABq99FJGEZUKUcu2qF6KkEaVNppCt6y7tnBWGzPBLVV2
bQq2CTGGMxU6ax1s2cnlJ1SBk4DEFw8kImrEC5HwMPhGJKXj88gXjuvQJm+JCsDR01KcRrqCaU6X
ofTOt8aJyo1jdVUp76cQv6yzzuQ5UuQF+mrkJGLl8xWFd37kRz6lrEtmLO++ZPGQdn35xdDPLa+Q
g6bTu55FFkVG4EGhlFB5xN8Rqr+MNq8r/sqw+4a/1m2QPTbigL9wgzmF9yuZMDEdP6BM5B4J1q7U
E70bjQCzhcM8EfXY1eqdJouISfQgnPcqN2axODKhyVYyWjAOkfmaLVf1CmMfDuoDKM/p1B11Ka4V
0SjpXuuAyIU0Ru5kY1ZWJhYREaDNTqel/4AHUkaWnkbzcGBGYu5+Mqv6TZ8Pcy3+28vSwASmDrJ2
bzBX+Rtft8qc6frAPf3ahn2DKgrOCMFzxxhBvOqISMGFm6VeUEGh/XeptsAM/HZZJgbetm4n3HeR
AlF01inWd5/HNZcuN+QAuyGYsSAR2KGnKqlMkzXc5lzg0IlRQsYgxzr1dP5ovfuMDukCfPbJY2KL
5FRhnvpjTEe4mJ28g91/9KHOlazaQN8XpKOa8MbwrD+/+gnKwWk1lEn2OaDm4L/64M6aLI8+VQU4
Raoqj07wh0SpD+Gm1xBQvPpfXujZxE5CZZ0HmQ5DlieHvcNEeM7xkolF1rYpfJUpWiL4D+swRUgc
Yetk89hoy5knl9+jKBUDc4qCCQJBBqyA8SWVjlcjRpAsibuoiT2pThTwutI3f1wvv9rTLUt+KmLF
ISt4OJ0W+eSWod4LjolUcqMQpHrgs2BxkCaXkAQLYhALd3p5R/sEoCK5P+iwq6BQcow/Z8eD3iSy
Ltam9T0guhdi0EZKKYVrHgady35qJhVXmUNVzUHwdNDMoHKRbD6LgTblEZUjZvGIc2qMyQu/Vi6w
CGkuLdEXUmIv71yjQEZvtTyrbpDCpq0mtwoQa6X+crxhp9UFElH5rpTp9aNYjR+Zm1kKsY6T1lb7
trs686YShepaI2xy3FFA40CHlv51kGLXbOQTOYngTVAKTJ/t/u6cjSxJBW4io+EtX3F2tXCWhe2u
8q3iMVT4ao1Vx70PagVAU0uxvWNmLVFkronTgFxE4veEcYcz46JSQvUXE0jfyZTVq11iJ60D+CGx
IlQltfSBc4FZQ4XmNhCa4ZtZ3ZRHjteAncT2Mhv5LzL7uLx+eOBalJxYVMIiwix1rm/XJuLpOkQ7
Xv5Z9K9PQFH43fdMqVVM8XgpfIQkZ5jWV4zBYWDR3HPWbz2HfoG4r1QnHHCk7h7VwI6pcjEluaVl
tUCci1xMZeRq+StfHyEVuSMVWndY9koyBbso98Lc6k5Ngc6X3/sjQk0fmISIhW8ZqhwGaBA2PbAW
wyWlDbHNzzIQGPBPkmmt2lZL3Dgd7QtgZ4wkah5Oyci9OP7N5Pv3bG/B3z4Tr4Jb2+Is4XFeaZdO
ufyTfmMS0k8lrum5bArOhIBnEWEFAmYQR9Su+Vw/gqPriTA5cjqHMfIxnfD+9DfV5norq+ilr2uZ
fsRtTBZbPcG9xxV8VRgglU0BEoBJyZSDWb9h98QIinWofwMGRq2EotGoH2eeFkI1xfV5eKiqJkGX
cosOqaa2i+QHvG387Nroniv1JLhxfuHrdOuRhzYyIjubTxgcCogV3QSAOJzhPjQOnzC91FN5PP5T
Uya+Vxzw+HBJCHB97ztyJSbhfGwmIs1zSdRcWbCEmDPY4SVhBnvGYgfAnkFfvTOIHJ2h7Vgxs09o
t4ZrImDqwT6icgGSVgwb+y3iYufabPgrv02qcr3L2psxBiZ3i4s5kFHHJJb6iiItOAa1gftHzuvt
maHWr8QPEDucCuD5YTaEiSpdPiwb37QFaUAn8mn7EDFz2srNEUgWEr5Aa4TdIkd5yLiCVxmDVGIH
vxvi+uP3lTG6vMSJ0k8ctbuSm5otji7MF3TsgtSLbiroCs9gBm2FilSBD20oeqfYt8pOqe/DvkzB
bYJmwA2IRsePcS7AtHiY7VFWvtv5jjTNkedbvv77Lc4qMjoAqxDWEaTxpC2L25WJOPZRCJviP5ma
JFv4wE0sQDOvcEc8m6++j6xXu3ETVo5XawNCQUQZlrA1wIeDzx3mquJksAUBuv3iGQD6MPl95I+o
69FQz505tZ+N8G/LgElgAGDrwXaG9xtygNYQOygfo8M4OWZhtDXP3qh4LKbR487zDyTgF9mhyDFN
Tsw5cG09mOAIi6YufgI/eCeMJbvwK1dqp/umCsIiYP6KAh3/NpRj+vqJdLM4kvQlhc8v3ShXSV3f
1BmsWXIGKccEMOh2Yv4bLfybHTGvzuDOIn7vKQFdn6HrjV86wWOas2ltIZmBhkpPIr59dCT87MSA
Swaf+Zg17OJ6DcD9gyBw17bZ8OCaInoMIQDVBWODJitnREgVnlKS7BQFIEI0ReEv8gqjvvje3WH9
hiJqtedlln7eyfkYFpZKL41oNONZM1QEVlSqH6WaKJT0n93Xwk9fV/KYEFN95CrELGwsQPKLh6Be
YDWP6LgFQ7iD3XxchNfOwzxhbuQP+BS+3JKVKwYPpjPYi/xIAdqRuUpxbvf/kysu6G1Z7CQHFL0v
4A7SH/43VDYVFuc0rfntjqkVJi6QsUtg7rLLlbivqJJno5EMxstJAxQbo+MdzlkQQsivEEAVX9ME
KcFFAnesLV3idhrsG5eFt2eRYxBQwBjjv6CzCZTg3hOkmb/gdaoc1YxHAaB43PyHUX+b5riIj0J9
l0FLQNgoB9AOVOC00isBX5SIugDUTSBOieZctl5EdLN9TxjegEbqItyhAuHEkQVGvwVQxSw0aTIk
45F0B6MgDsxWkWz9uquD+VjP0cSkXFYPGdbaqMlJADhUQ7E156aVlKAyJtKzMOUt52noDQax3YJM
QPF/0S5JzIzHQTrZXeYODbLAUt3d5lfUVscoIlgcTB66kBjR6F6JPfH1zKxB6yEqmfVUWvf+ZVr3
QvPfHCZczozMW5DOUDqEaIycn+gJ0EyEjrQg0GuLp5uJkfB/TbEyeOsVFelVYZ8byto7I4KDqppA
bO+0sD/Cp7NaYHduai9Vd5Yom3vYE82OuVEpkNzbY7jsdB/KrAEyTW59UCg78BXg5hO3J99oSJbb
2QwiVWmYAlSkuAgvhQxcH2pbQasiKgcxYmJNugHz87hU1/WHnFT7K+kYBftaRaXOucnKQwdaVWxQ
FzjRqBP9fuZS4coEGlEDijo/BrN96oZeXk/D42rsTG7y5HLjw3np/7JXoHo6qxPTu0wqswJmMX/K
v/RLvIsysLcGn0PkdpXNm8oOSEB3jU53weK2c4lqNVrNwda40MUqcu4NSdh5gn0gQXm0ISDlMRa3
9E1p3lZh0TAS1dJpWyzgK22FI4BhNMSX4oNRTfiRo+CRJYH1yHtDTKYXweFeZLHQn4aJnWW0x8CR
rhqXgPHFjjloqv/9bsVm86kURKwYSQFEtTT/mEBNCukWBFscDAE6TFZFouLZcoLRO+rSdc4EhyGA
EV8tt2N3NZQbtWzyOHKbcIQQRgiGZZoz9CuGuOaAxdYYN1G2+KpwQb8iEovhp4AwVSDNw9lCMzJp
a3gplf2A3Ra/zZaLgDz++95vk8YKmf6DKpcTlxrNRPkxX+Zd/vEPzsnHqBEM8T6LTsng3onXzhGn
Bz7tQJMr3rujCw4kPJZadiZO5cp9R6wcGMA8Dm7moJIOZJdrOd1aaRpXarh9UkSu+lbZhBSZYqih
RalnSsJol5jdCQ2d898O5wqnUc3B70p4eH66IUFdkP/uy8nvvaQRhMu68KYscOUwwYbOrAjmn2ms
9dG+LQP01jlzK9aAnBgBk1t1z8oPKUtQKFGrjeYmSsV7XBKmGoSQXOMYFTQ8sDbIz5dS/DVFZHWB
NlS3zsI5ojNQgPgcZt3DxFMXFbwFY1wOtr4SX+KWgCL7a6LtuQz/7XyH6S/HBDpETdYpEWIULasw
gpXHz8AJjxJjzZasnQ9sRg0DOLVaOJ4XaXfjbnuxz8BQTQQ3NOGIdpSzidBxQblWJ6edl2sNR53A
W54NGaxBeM+H9OAk3uc6f1dlSgQbjE7q9jLc5he/QSmZiK7N0KFbDO+3ZqFHl1eWnOyaZCLolciC
WeVT4UgI98J4Yo0OFGGKGxnAjnJQbK1GinuYUpbX0GmQiMwrw+aMbjI4bUfRehnPAM003JSZjU8U
sJMJwzvcdMNMo975CDPEzgxOT0T8K9amnDEPgQKEwwnHIzJRLhexWU4VkvIPWDvr5yywbEX8CUwQ
kkwlYpPXidxhw6HJZIN0HnBGprlpw+hoNTJN1vqnNRNoX+iLNOSgfNIVAnY1xQ5vpM7rNaP3NZhE
b26jRGXMzo+YwrecQidZY9dHZXHxBGvVlAgbyLcfhPc4rNmwzMaNZPkkzN/tgQHffihHu6pTLybP
uRaMpxSwqaXGeb85xbqcMc0WishkVBTdl1s8lIZP5Vs9fx/RilMIBv+a5DCHkc1nzF97YinKoB1B
8Ryw8BzxjRcicQIQqDYpK44Mr5AvfLgdD8DNchN8Xqem2xO2OH/uqR9RMQ1mY3k08csooBAOKJch
WilnE0hQ7ibx19+kggKCLCvV8GAMMNzfZ77jjZAGQZK8Hv0k/VJJaU+LP04LN1fkFcPygP2mhVYn
+3VWl2uwjhTvmDI4eieMpzvGTaWZPmJYdfYD0wB9ZtqSqyyk17NByuqdBqqapv0OP8Ps3iVGK/BJ
3qya1ZnA45yQmhKL/DVzVqKKnp1IPns0XV4Q49qzqOCDxcWmcvTpr0Yuv6rtYZh1YfKA04oCmAwG
6fc64YVj3+IeYvRzaxa5CtGT5VKcUUP/c9z9NTLAumJKO0mj8xeY2X3YIwMHnKODG8KLBvwgrTJp
eej/9xZ6+PaUUmsNb1DdjODU9Zb4xDPOkta2OKLLscPjxZOdY3uftzKMjdURCiMNR93M1MyxVO7p
Xfc/Mocrak2y5alJHTR430ouxlDbtIxB9axvHM9T6uF9Hy1Sbpq63yNVhuTkX8XltGvzAv9vMCpK
MTD7ZQcOkhiyKWYDQEzU6BK6PN/lzWBpXDvKRpv8pnatFmFP8UjQOQt3S642xj0Mr1QzoAhzB+xA
KyHf0KbjBjyZeqkmuoR5580B7SEngtsC2lcGzjiXeGuweVwPGqQGQ5vO7SLViueK9MtJIYU9j9/K
PzQ3Jr+WdZryw4chCp9APh1GEA0jVUA4wIlbT+Vb6cDIR4gf8yleqnPv2qa2maCWGlHdioxBrxzx
ILsRXssXYxta0XpVYZJ4fO94Eu/RIuqLt8d/+N09fBykxhS4To49Nd6q7x6vEAS6qGkKh5csELHD
tKDgeKz/Gc8Ch+Cga/HdpQ4qChY2ly7xGSrdFV22SmBTAsKMYL9vcTLzNUwwf8IwghdKfjKkOnU6
xDqu0FqP6m4uGRwsD7m4/j4Y/DvD3UgnnKP9dXx3aC7sB9YUA7B8uCmEKenVOzcvKZ1v3cNYgqBY
C/kATNjWEjqkn6e8KfERM16nxFWefbrR87LESt7No9SfHCKh83Wnzf0fT5vQzYdexImE/DZm70Kb
rqh94EOybUBTGTRB30XrjwSNdPshevNXZ+5bQC7tCsD/BiliQduHadNiuLpx5tIDl+amnVbbOUpJ
eP0Ez1hUPEelVJcZOiTf8XRMZ77Rtaz4Sn+7uwm0TepR28l8RwVAGQ4ixDoeLEAyXYW/NQpTlT6I
eFlKXIR1Oa7VjZR6tEJpuQBSm4TEW4BXVBfp+hbjw2vP2hzM7+adn5IpdoLHJ42OdNnT6y4YtBTd
vBR0bQiE93nSZnrxbPIf7hIofRZge5wUJgsBN9XOmTNEbXCe7nucrUolhVZ9j9498XaQzzXZMC/E
ioysq6i7lpjEurr8h+Ce80Cud4G7m4XE0w0FxGrFGThrkx8760c71ORLq03Rqe6Qmf6Mj2Q2L2Kp
j+rPFvPramCE6KvyeoX0gOtLGqNiQwVzRH5BuINiyasLCxb08Q3H8SsZ/mjf0ZQlJ9bIhPGf6LlZ
VmCLrnM+pdUZHiF9VuimKM9XXi9LFKq/JnorzSbKfyIHFKSGAGrICfYMqLjkvsMn0BlRxgFDLH4f
a9yzT4vRIocSRQDK0H3RR1SzOMJe6G7PirnxdrO87YcUFizuIFCcgz85jOSQGlbSuCuZ1RXSH0CS
2qhx20bwFk0VENa17zNR2Mh7XdlmqVCSwCgzchgAvbWPb7dhkfx7SuGKXJezlYvtWy7wJlaUCuIM
uVUjJXuNjvoEhqbVGvmmBzW5a5zXiKmHaw540woivxehZWJudYIcFxPcdQSgBeK2PeCFd6ufLRVX
p/DCCq3LRkoqSZSmxIxzyjHov9dYFCwlecxtfkZpvP1ZnzOsjZJ9LQ+NtRe6jyZ+IooZ33+/23pB
RVY32Slv7XKv3BhaeYcx6pFMNjCqZ5vcDZ5rmnQTSCsDMpkHujTP56tuLrpnvpU6zw0o+n3upQ65
1JZyu8SzknnYSZakkXntOfD8JIgGcgDL5Tk2FDKOLaR4/rV/QkKJnuGDpoMEdXAyX2RwZAmVGT99
SgKThM2WlodYEPvEqVRyJDGh1O7p7vcz2/LCkSseRCKgAj8Hdm2esIl6icjqazZSLBFqXkDMmLYB
ixQ4cFdW8TwJFkrvH+o7FXLVpgA1uDh2BeRQOTMXPrjcWE1BWg+3XbhsYg0pwnQ6KC3FCQECvCe/
Eqb7X0gsPUtFvF0XjubvvXMk38gtz4PO+zFfLiEODtwPwGkiFi9djEKfyAPeZA4ebUD9SJjwReK6
frxrARCjpRCkutJiTr7Udm0BOITTCVU6gHNk/PBxJG0SkpI7hnF8beiJCZcaZ8UuFLuDBE5JzBtW
uBab1VU5IhloUwX47qywInJpQnDvfQ5gvWOK9V1MVYulc/m+CGS+9n/1CysPOrwLsHqMXP+S7RsP
YLVHGpKSKE/uwlry07EohIdCLPsvkBL9rBg3M2/aQBKWh5HEk1DVKATkf2rnFXI+YC6sKd4ibnvP
pxLmGsb6WL0+hjWzu6Zpcwa4GeZgpo2KJkQnVKOqAEcgWmwGnXgBzi/OHPC/drTqjCmPPAaX5Zou
ZlGWuvDC0cFui8iiXWqrQkWW1uIZdgzxc9H4oDCopfbg0vRTRmVP6jpDTg49NfUsrnUyZdHoM1Jz
kVvHejkMs94oZvaTsJpuxhh9GH/M17GCM3mU6dfvcGg++wAwGDvEIOHj5HhN975a94zaqhlamAen
w+f9aef9UrMPQi4c7M6Qzg8CsOaWGMVzaCNPWEp9837yAy1z+aSU4w79N5REAc4iwJCao0NOUHhJ
1gESLnMRdFNB8k3X2BX4PEYYj/ApLqHwdg6NYogH6BhIvFojryXU+e74QHeKMd09pq1NSBfdePjN
NkTMnS+7ebHRv3BUmX+E4mx0nJaJzO2zZ1M4A3dwWUEQEw1yzG8cqTjCtCgmzYECm+vfupUjiC/x
IGaVEup4nb/NbH4tvw2HnIM9dwkqzSPoM9Y4k5t+Q75EPc1rLcJdoHQhoGn7jRNiEfSliV1r5vKd
0rK69YBwPh+a1uwGN39bzF9d7MJ+ceESbs5XFx6TRE0lJg7Z41Gg/gDNkC5becQW/WksxjzSPXG4
C+75n6Jd/sqsjfQqzRo29P/Kn9d/72Ci4qAVbAb0tnEcNXJbMKoy9znIDy48XSxkFTdIUxMrFYTV
N7YGQ+k6YCqhnxIuhLBLiRZMVVMUD0l2Evr+FNwxzZj8Foya1s28SVG2r4TbizPt6TZu19U22Yh2
hTNZ7lm3xbT2DdmH8WfSEGfB4jL2P+zMRF32VjfNfzgoqmZ98jCU07lon1EcDjK6Kxharr9qNfCd
IvpiXhrYN1M/loMy+DxvwJMamjg/GhisGH203kcsK/QaKjAahRwJfBaM2kmOLTs1EKDYyrOpAA8o
swrgMo1DEHVCdOHCpPawgUfK9MfUdQqDlQUEOzhLFSsZPNFchFZ9+QLK4vM1rf4eh3izkaEgXBOm
eW/7hZpB4kVjnKymTSAsCAS9tBkeRHt06yFNA4avhS0VtEuxN62zd+UFt4NCogiSp+uhlVECiYVJ
glL8hC0KJ0MhfqY6By+D0R0rpoXAF8VaBikuTFxByeaiGRkOTRcyrbgF5oaIolZO9cXsuajSjfsl
Lbsa0F2xEL+RgHbDrdD6/CHq7Js6ri/vZGk/elalH/kduLuSvkqKXCNJZB/FV6lqPTeucCMsU4HD
u0SL73WUJQrGGjrcwUfYJyK4EDDSTSGMHD4Sga+IhHmgqWBigbPmIRI8GRfd+bJ1dk3/3ZORQ7l5
V9qvK6MwvD+DUWsuYgQzL51ZRb/GbRD3boMu6XJhsbFzOONQwm7LUXXDkIx1gaVNFCX5UzIhVWLD
QxoSVuGgCjpZUcUPVnWXqsidxAN/QCPk2jeUJcNE/j/e5/BumgB/co1LYyZRSz6K5MdQksYyutav
rI7PnCN34NmWNwXknj9aKjqtc6OUIrxeXxbAUAHFSbu47svepBgWwJB92Obbv2ECj+voV7kfXZPm
I+AcNBgqpBh6ForM12kJmBjh+ZjIhn+ijbM0n68bwdnS7LQMg2MNGYJyu3U+/r3aWiesbnEBWW2R
emTua5YJls5M8GAH76mj75Et7UoVGYzFjCZb+VC7IstR7gD6EYSCU1JfLXOLbzQ01qU6nx9eTObb
yHHZVUFh1lvll7yUCpgaxLV+BGyDGwpwlkOePoEMB+x+2iJQuxed1sl9OOs4GVqT61G/BTTsmBr2
K0uv7TYTp2VjaGn1mhvd8TNKakiDlDmsAGqZ6U0QqLPPFX35aGVtlyNYpfXEpseKxEsTSCbUrL4y
FZgD8gfKJOJ1MtpJjzOkZmWW1LqNBY8eNRLQN/l+owU2VlUGbGF5oF+u5pJEb6hvKCcVnZl7NlZI
NvNU1zW+qRsiDkQ9DGArXfJDrFSqq3LFVVwIj+9AilEwWH3+NjtZMfN0o1MorsKp/4LsQ+IKOCvc
DOpRpAh2c5lqevc652l+wUXQa6Ak5DWK1a9Y1QRFLfLs36GZQc0JlH2brRb5FFBhkRyOLXH4d2Jt
k7e7Px0ZnSoO4usjKK2f/INT5S+YC37cLn9vn/8EXHsOwJdngRrglZ3TsJ3pFYKU3Wwy65SsUHGH
Fpi7+KjIppToOPM18pbI74Emp4YrhHZ/4b6O13k0U0ki+RWPHV3vSl+ufmqBv6CJYFi5sZKexs51
9lfqwBOvGtLdtTPARm2LpEQuQCA4ju5XPS49hddq5XPJWXQyyx5Y28VCPsjxrbsiAUpvZsPLgUJ8
wlhMBNzf6pOd7vvDGJEg5CwXgo9TBnM0F1JVBQfNsxjZlf8x6SW80V5NHa8P8BQoJGjPokLUEyYA
o3lBQe2Yh8fdw+mRKaEgrmvTjeoTD5gozvWQp4dbAWymGcgjw28tu3P/6svE1+54gIDBATVGNSTR
0U0myDnDTXA5zi9qg5mhBcAL65QBebVtezDaO0oQy+FmddTc3cGf3pxxfSSdfmLA3Xu/AQvxQGnP
KLBrk2FpfhibA/IO7gI8O3VqxPgPf5UONs6X1sDOyi3J/3MxDgUaZCU6dynw2oSIaxG0v/3+HzBH
btsRXOWK+WH5jO0hTNtsHjZj/fa4Hp2JoN+s25cWH1SbI83rzptb+9uF0XfZkSH0mrWQvV3ec9bg
DP1/kksIfr0lHWTaUC5e5NeP/bG82BwEUO9ua53Qz94GEuMqSf5OBUh/5ww4ebPUUtKLpMckyj+H
WB5Uv/GF2e+jA9MUulGD/LbMG2dpwZl2YL67W3x8EmwysjMr5/Uv4IR+nvV0JmH9aJiH4771ZICS
PS3/7wEmIWBOiTPL6ncP6SrS9DCkJLzmHZpGBCWamcOc5ZuExopukL9zV+0ct0Tjkzyaz5aYdfHM
Jg8WRLLr2/dwwTMalmMYMsr1tAvXH2qzXTgEdvh+szT0v4B3iUIODR8fWBZsc6funasxgcP0KitA
j/bGY9pB9heIjLvJ9bxBmo3giP9dfvn2ji9yyRQoDI4j1TsuiS+MvOCPrXyFKttSuxVcp3zuK4he
gzUM6QsUUJOHntXjdsF+QlL758Xb7pMzVQzC8Zn2kGCDBdavlJE2wolbYUwpnN7zaFzlZfhed+/S
tLC09G6zgW0BnlmFbU7s97sdyr+MkJgsIyMUZtV9+sShvP1Q33vNqu2IG6xe/Jl+LDcH41VNGzPZ
W1D1sQqyEAoyme5iu4MbbI6VL3eL4k0s1mf/SKX5mJdkupvNgWb3q4zzYF3YYmoCNO5TV2EusAQ2
6pRLtmTjMPnn7SFKWY58sNSshkjfwGkNAYQ5pYXsQvR/fXGK+heqop9drjIqvgdakaP4ca9Bmv3g
1u5Z2x7/9aek+xWjYa0znjiXVbJxgIQ2SdchkIXo8VkeTTJ4GtW30YFgyCm9zY2XLWSrZR3nfSiC
VRpbPChKu3TmnCZ0EgV9yDrWJg1olBqM+EhdDbSKnPBDfJ/W4eerb/Rmb9kenp6v6x2VrtBnOb98
PylH4kce+VxEDwZjw/HnOjVHV/4lSbaClbT8HARkAXShXYnOzeaXdtoGwNswtS+zuly9/h8fCchS
OaAkkAUUdDVDkp8SwefBVVupGDT+evgE1MYQhDNGI+QS3fn5gycko6fyfVCSnKCcCDTjzN+Xi7mi
ghnkenk7AtGS/T928nvNYISrWsmoPdf730HiBP3b7gLke/OBuiyKcYtLKKI7MQvEXeY5G4Oe1MqG
rTYYQznYacNYRTiG/HzvsvQ60aeqphQ2kmQ9o9IyF0BbbYj3oSKwyr8Xy3PlV239Tm76at4X9ehB
74Hq0kpk84esx3mJ1Y2mCIO9iwlXBbBVzvKsdx7N9hl3G6XJKzK70X9wNp2ku+wMiLdKAsXjTpqj
4sYn3d/y0CdQ/vNeX9ZDPQphHj4220UPSuyQGtGzFuzHkK02hT6a+XZzGI0Az6m65tHH+Vz7iL2y
e9Cfkr/SD8ataOa8uJvlHQV+aT/HvlHQRRPmmVAH20HbopVKhxWf7VG2kWDOElgH3HveHBK9/Vbe
GiNQLv2gOteXbb2s68Ywl74eSKLkKhj1baRAdDPuzf1TY6qNE3t/y+ETcfR3FZOkOeX5SmFhf+gd
VA2h6Z9vLHAsjzqlwHj3MwsZATMm7yzsfU3f/xqlcnCIvRSBXaKhlT4hXP4th1Nmu033UtYnnz02
fgQS+Dpbv8CK3M9cNsEg5T/H2il626h1KZUgrI5OPFBz+A/YRfpS7Z1JIp31ElrRfN1UNwLfZ1u5
rjYrl1MuaTrl0gej4WPpYwlU4fkk/WlwzmCsFGOQ7aaj/YOXMpk2JNBlap9+udzxPfZ+8OYEmGZX
IQjtNDBooais8uD0kjuuX9EkRBAA41odbd2KMH9C1rtOdCgiQUBgksNHuAG/1v7DSXKHhjE+nXTn
18zxMEL3Kyj4Qr7qEoHJ6Apzkx1vSYerpyBgzjCqosUosOhipBLyyhgblnA4yUfV2upwQc+Zid6d
3E+qDWNvXTG8rZa5+C7VOPBHEC/CFutkk+l1LI0fWFnTPcgg6T5t5HE+O71IbK+gW7iX3eZ1qme3
7T35ip309kXeBaSv/0cmwYDCReMvdHreMTDN9mmnOAAIruvQP/gY8eRSyteZ1R/f8gW9GMPJkF4/
X/fRQHg2cEoE/RfmjNxBZBr81TaNpK1Rt9fS9/Hdzb1yuEhH3iqYkLE1rU2gDylHuGQWnQVR+vYc
h6U0TfpSnmA9ALWi8CXmSE3l3nGZ2ryMa+lMMEfMT871t7J/8LmJO+X4ielYXcal7ZtLDFUjgBYA
bj4f/WJ7MhHCIzD2AzqPtqVWTmixCkssuVcDrTtpM/yAn8LffUDNZBHmRrLSr4NMFNl7FCRBJtX3
Q9J0alc3kvB73axcLT3TR1asyr9FNlooLYcPhBNcRgaxfKb/3IklhYIQmIPYXl21NjHkGq1HNlM/
efr2phDwmOPHQPEOWTHy/qPrbUZ3ZCvb4GBZVUThkLpXzLcgo697ft4PYftbS+kR7ZPBFiYMSPeO
LFXAJhxlob5Zsm1krWKXNFvx9cMsfvCJrGsA4J271urYSJZ3Lq3DQlQmDq0OoS7ODJbj2oUSu6jY
fDKaIOTC/xu1KuKwhYUEmoPizO26r4Pe2l4BDPegSsu0JR6eCpjH+xr/8Nd8fOvGKvr2qvLuso5d
diERdjNGVFU7YOHk/XQKQws+6+tA43dC/Y8N4DE7JH4JNcrSw3I+tADZP0XAnLvsZr6vP4/1Cu6s
ZTiTFc2ZLHecWigV7YjTV63vpZDSbWTd6Nm6lCrZaDYXW8VsuVIdGQ4NSiJ8d6Q5NcdooDIE4G84
Mri+3LFORoI4/adFpr7SGPBLYXwNpVnV8cYakbAirPwmaYWAUjLuNvVkVu9/ZORMzyjrTkFAvMZo
H3kCgPbkWMWnV1fI8Wz5hTtatJKAfqV4jCkwRy8a8qviQGN1gr0qFYod+/3DbYMAcSF88zASGqWb
GCpGrsJiymDvr51EEjoQovvToQH+11iPqRItYeY+DCr9toIzqsdLAzembAQHKrUcPp1+v7sStjGz
NV65Qw+IsBY3JLdgXPdv/KgBwuUX4qBPeLGs+xyJc64+3FV/k3vB2WF/f2Z1CscZ46b+vUxPcH8s
97ZfRTVCkdS4lX5zuMBeNQGNe6KUG3oCOnrSECOENmbfOqrW8EULVjhqsPmur3oDb+oNeawELnIK
7SlkGjA91WSxKBOEZPX427fHEZMqDutUUy2GjqqKDsOmntc0OwooOzivVcgDJVQLT3EiVEZNRVqQ
pWRxKUwOqkFXJz2z/+tMqbMdJ9Kz38cP24FCFTKLrsozy9EsafycL5PrU85dPmnpzCaWZQEq8AV5
N8+WqjIBCTl71y6CMJEdKcO305kK3q8vnrnrKGUhxDXobyEzyOKzDu27WiJRxc7eb0Z0gUX6QsVs
dqQOGbUdWuZI8rz4yIn+yTBNd10XcA3ey+3R6ViDoVuvEg5+/RR6KpkdVmYurT009kwK7ejmrxg5
FZjMAo4yaxPXykp8uz57dt9C0b2CPEsv6jXNFrRBnLbjBi2au1MBFCg4c+dw4d2o2st2AbgWERmI
YPx0/CC4ZWFiCRxaPbNs+hKzYhtkcwwv4cj4eexY5IdIKQSg8Wts6MyvhFzGgbx6tZWMavpKgVqt
xR17S2WV56QQW7H6aJF5t5w4TlT+0nFul4cv4iC+o7hkIFDmF19sh4WccSTzO48LPacSUljS+bQe
Q3/TpB/yJVXip+jY0ALSa88L5GtrqesRGJ41scU5gSccF4czy14GU4PGDBZbMY0ZpR/fvCW4x4OX
WyY9QfjYmMJ0/XXhftRbTg5ISUuVQ+xsoGOUkyqguBNxrrc3kSmLxKozjnslnr708fxV73bUVoBw
L28lRiIcsDGUesTXaxAm8X+76th8owps93A46ip+u0d9vZCxQa9nP3NwmlG6KLa9sXUc2EcvBVmP
xYrbvOHrKi5tI/Xh3kMIFqEtLK296/11Rl/wCUwNjLLCnimisiYQF6Jz6rlnzVhLFmM8OHU1Xcrt
JU1ReSfQdF82nWmscKXlXS6PTBV19cvfltRUqY5739CMB05rijUf05Ipe9DBxubvW4KSjRzedFBN
FvQWa86KntgIoMVpfq2EP2CSJF7h1SMNdmpbjz9U9P24hEeHX+d2bP1qgBZWWGUqW/PO3OS3Dm11
oodxV3nuHaL9OPPbQ1YUGid22SWxtTNAAI8ppeMFZcnEOGzBO9hyffOGnXiVYDOIUpIA8lGKDZPM
OkQli/H2sJKDOez6Ml8cta0NqDxiFpmI7dre49xI+S/Ilac/SNPZjEvsVftp6jq+sOjfyzgkwsc4
P5zhqRCqDKhOUKMT80Q7j+Zz0rXGiBy6BH2K2CGQnz78cOFAYUEuD2EVwvvXckmL98N0faAQPLwH
ID+CVQepXMQrZES+9BxuVxB3J2xUISOpy+1F2VbgsxkIautKqsFBDBd0s5pw/NpIU9q14/Y4zTCy
R0+7douZt5N8qLAfvHDPXp0ETWmy48WbgP6wTqtE5uYODBEXAHXUblHXxs/q5fGkt/v9PIi45+WZ
YHyhUsQxZcjEIsbQBL8jRXW3Qg6t6t07jCtKNsp/Hd8yGE6l6X7ZHCzjRHIGB/FGf8DcVA2fShRd
ctRUyngOiT6L9Ki+eWamIhGeVwqsbJ2XFjAD5KM5oqm3TYLRwGuG3mABtFaSshkt0J6ETckOiI0T
Lw8sj9uvGxFhYh28HRBBmXZJ2nqufcybJ5l4t3OaTIxMmUA1Ss4ufXE0GoWm/BFzLkG8Kz6hdmXQ
A4LY4yZO1XmelCIahw7tkFXkhMe0VsRRLniviAi0whO1zsQCZMlia9sLnfXngyjyrkPrEdof0fOu
xzZbUdGSc+ztkRjC7T6zgIIoLYARd+b8WYEcHN/DdnSJjDlLEwkB5AbZJF6nEKyHpIVbbLMDAs9n
Bzs=
`protect end_protected

