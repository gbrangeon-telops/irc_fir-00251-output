

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
CWO2bSovBvQ2ByFi3vbGk64Kz9+OlU+ol4ZycfRhtc5mzW4spj2ZUNH57Z6TD/HWbssYOjRT+UqT
ip6xHZc7sA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
nB5KuhofnITTIpXOtfG8vxQ8BtQATMQkEP+DmIE09Znrcw3yJd8Ym9iSaEwPi49QFbQ4UCNnUF1p
Ci6v7CITkdmn7C29rKsxyl5fQwQ4Yg2Y9J8sH3IMncLyMWd/eC2FXu2c+nIyMZ2PxTUPVrUjVKNp
s7scT7Me3sAj5vk8vEk=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
MNNArzGZfZxohM+fQiY689sNLR2SVnrB6IH+/5sMb7hSfawQFJxphTI8Kro2JGGDqNxumEJLUYrG
7mZGSE03rCaVpdhD6Rm70zB4CVRXmxwbIpEK83cCm08nMbZ8k4fK0avkhJQjAW3CnUztsuq7IA0K
kdwznIXZSyXH6lPiqjIN2Skr4/LMpA0PrKFOFlQVuPkT5ZvNvxenTGhCq9p/EpzKYQA/Q64z1Pcv
8PTscPeWEIpmqBcuycpxO0kwVqiQNRqP/TotOuVFkjYLePFpvLupJo2vDdC4y5SiD3RT9wZvaSz2
Bb8UYdK03OxRsiXtjWytUX0MRrf53QlD+4mRvw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
JO39BJFIHsw8fi/kSg8TBE7CDuzx+VxY3tt2e34SSpwe1+CidGWrS2YpQSFw2o2o0JVA8lhp2pEl
VW+YDwewZ52gevHf/k4qIWqrG228k15Q2kpUAiHbcd1YG0RCacsRIqlWdSiw7wc/2b5Il9la2dZd
yyMNm5GMzs0PBGaInn8=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
DxfcLsCbVgOrlbX9FvTGJxwVAV0OB3tR+6ByNYT/Wivn1M9TCrq2dM/5FWlDqpdxHIYJfhQjjzlJ
F9cbuhfluBOxtIUuGdHg2uX5LqlRjgmnPZ6fbuzAGkBvSUoSqWJpXOKWx36bmV4iGY/0e23H2hgI
ZyfwOhBcKKufNk+Nq7xnSV7GWSBSiZWYhL47CEdCY+E8EYmyeXyXT8RcA9zqsfKsEZqdz1rU0vql
DdxwHxaE1OVS6MuW2h6qgK3l9I9LyDohZgyoP4VpBk/e9sTSLxcSmGiXwe6zlvuSw8MrBIn34Ezs
uAteiO0K8WEa+5P+7J56z0wy1dst9IfRzCpYUA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 45648)
`protect data_block
y59K9Vgk15TKReKLDfxjl/BS1Q+WoTfl0PEMre9yg9VRkuR9UlMpeFBPPgpDI4RHJBgblSfFrn+s
3ojeKeHqklduyJaR/fw/+Hu8U/J4ZtGLtmSHJ2dj8p520meFglAt09ibmo3WK0zyqY1GckLdUNXW
BTB4yDHSZg9jysGIdYC04meJUstxO4KGmuBi17VfXccW8UVwbLKCfxdW1uiFY1z13NR+spO10/U5
qBFaluqJvvQqD15hzGtWjcsYdzep71FlMBPkVEHROaaMQZv5aHRBCV7t2C+TkMUiRfeLz00eyUV9
vLfFi3nda6imZryMhiLJXQOlkBb6SM5ouW1OiuJTgPuKioDmZWBWME0kThFJhSk9DM7KsKJFVhij
Noj+ClCcXmW83EwF/dCXZoG6TnAcVJn0ZO022AAreiB21eKtJLXJyEPd8+CkKmP/LVphsvdk1Qyg
AYysgnmekK2Sh8WZEaY4ZM6N1gq6GsEmr68qGdCkIQLOybzNko9zbi78SgNO+eTqVVqf9XGvthUo
CIXPF8sr7a9ttVeVLlts3EXZoOU91jkeRNC2nTG3cXu13acD+GkqNN12vsacaCKM1Jt778w3a+JQ
tBHGhrEMm9JeMv65RywhTXEOwKWlh7L9k2zOQemxMCsVwhbJy9PjoYXPojJbDpZAwfiymOrlyOrW
prHSq0EfAaEy4r3rlEesA5ttSUVQ6zzAermMp0+8k//tWAsVXNdNvK5GapRbd2ygE1pzeFcdzt9T
a6bLlq62YIf1ZiH71UFQZZDBFQziqKOfpA+iRpYVnyVdtx4N5i028Du+XcS0TGbB2p7t191xBgcJ
2v9wO0KVhJ0sVPfiogzD/8yJHnrxnkL1X25OU6V93UXSrbiFFavr6oxtjeyD7pi7vsnPxzu5tHDN
gFU2AJlsetWKqr8wg5V2hAxNXiTwbmuNYtMQ5/1CWWzifbhVBxRk658vHt/ovGxPdKbQJRIYHqT9
AsVrpaU/A6jAeYK1oP++3s3KC++gAelfyDa5a6ia2io2VBhHhtQNjne83fsrZH+UQGHWMAaCXHPp
iIm0nkmwTo8LdLSxJMWu/CxQ7Abfak008peZ09rddH6aFe7EV8O1gCd7w9Bc+TzNhs9lcK2yGzCE
goYJ2ZEC8ZO8O7fytlthCKjITeyR01kgKwK/U0O+yBtSsRPL51XOWEr6iJGABnzTWUU9Ob0DSVYT
/07lJF2aR34U1Rx/Ybncdk12HxwlmXuy32ARgDHnl4WBf2LUErJIwUFzakDjsXhEWD6e8MXZeJ3z
1IdgB5qvUVkZ9hKv3SDlIbod/jqIQ/w3j7WtvIwwrXUKjnfAX9UVncQFdG/81wXHMetsupc55RPP
aG0YOURg1WLKxdACcENAS0ehEi5wFQsvfeNCn68KAgxg1JcUAvTd7Awvf/QhkNZ3Lj684eUfk0Eh
yUiMi2HUxe20NphuTpXe8OyoVSFHaX2kpPmcjraNNGc2ZA0RT/Qw+pXv1qXBS+iUcn6HYOin21tE
qxmG+JP4fJ8AHlmlUHZSn1AKuWRO89U8ZDh0iC53MfJGVGzHcnnhgCPuukXs/gc4yhzewqaCGCVq
ZXCzgPCtVy0iFJf7MbzuYfDuaGnlz6zbd8YAYr9ARwXdNHTSpT+MP/zubH1O8U5DwR76qOLw21ko
6IB746d7jIdtwHczRPcA4/VCkpJ+/mX3S5vDKyVL92xmfI7W6I4ehQa3CCSC87XTc18khzhEpnSP
/RM1nZDnu1fPvfkSEgLcvkAjGMfLcEz5wI006Sn49ikLFjlvzuxDVhhOjgrUrrYwbEH/zyWErcs1
B9+X2ue45RtbT3ewnHdwiUI+LR1yhJb8t8PaP7xgaVsduBdT1fWkAVnr3RShSevYCk5RNoDaQD31
RXRTrLInlyN7F39eij+MWljWfuMVaM73Vm5pPFk+W/iM193LnFkbtgcXwVrA8U1/qmSub83lz2x6
v2c2bKlfgPjUxU20IbFbOUfouhDQhf+o4ZTqb92Gx9v/AAxvWNFQ0xRxNDTIEU6LBRK94AFdnLVr
0bXRJASuzTRKgUw6oFY/leEwyI2hPJLJZcOygF8o/lLbpdofpu7PdDE3i6q1Axz3o0dNijwB5OCj
0u1w2BXOuxOcM8467Y8dqMzqBiRaC6vvtYPSzwH9PMZi2LVt9+j82z0fCOABz4poYJXAh+wGk9f8
wNlSWG4iE5k3T+UVXmxl3CeYxgZBPzsKl4NCIu2jMTmbfbFVMmD2kseYfFiibYZoCtykDFmi+rzN
M4JNe24x+a3lkLlmpOabG3YuG9DR+s5GaZmpEHJ1mFdT5XYpbhhGpDSX0saUw4nTtLZAMEdKt4tM
X60njCAes0YmR7p+ZVu70dk/QT/uuAFvkl3o0/oGmSYiHDf+nyCMCiqUy3QPF9RDqSNW0VAXzPDN
t9gxKXunTM/41nRgqDNwUqeG14IVM+TAU8Jdh1VgS77R/mKJ8Nf0Mp5lxR9/gAwOHmPawbBGKp4+
zIepJtnbU4srJbnM+K8gb7H6SNtBsNOYuhg593VXOZfrKBmZbqQ1BpTshkohLu14LpxLrMobnnaL
/hPrRKhmuX/Arjvfo+521MAM7pqtjrRK7ZuV06icAvUPg4+RKYXSvXRgTbXosvbZSiih6iMMUJ0h
PNG7tXYtaA64kB39gOcqTzAxRIdodMBYUuhmDOFYQClAdWfNZ+vVSYFyvp9uf8wRDN22UDUO63Yj
OVSFwPE4lfWd/7Sc7C+aSYv08s3qN1E0w1UDXd3B++jZNLU9o+ol2BY9yU6ehLNuzkjR+QFtKYfX
n7hhZCBF3youIf3DpTr9qy9+OgO/JuEUDON9OZZxiFd3C0ZK7W5WtJ2hktxi78oiV79MiFBQRENC
Z/MEX0QPOYZV2YNlIJmc9nP67iVL+XT4V+0SeRpoKfYRDrRiXtMEzBNiPwPw4btO7zxjXGi4TUCW
riZwg5Na/Mbj0w2mSPbfxUr8PhiwP6uVnRG1878wLqZOvvHQWsUC/fqfW8+4gNAjWaU7OO4lgHzH
jY/+YWwF9e+jYZfVPjYI7dhz3B+JRfNeFkLn0oDUD4ARnFMTibw9umE4Q2pyGs66tU7ZZxb2hiJk
gRyuz11xv3x7YbFbI7oAPsoHnq77QNgHaOO2sbZrJP0l+FL55p4DoLDWtmNShoMul8BytxPi4fBM
qdm94CQzMMp+FmaFIaWvaKsZ4UaVsP1eFhim0/KvLCRnm4UH6vhux9+ekwX9Fjg7hj+ZKe0fxwwb
dTayD9wF1AjwsuiXIGA1a4058MDBJ2XELZjTNjy1kitPa8ZrgfYgisiybVntqj269NQHXKi21mAp
kaE3W9RqtWddT4uV3kfNFuzKbHsRDhVqi6YbUplY9SBOrr6VBKG58oErf9EL+X5tR6yWEvusqEI8
CwUQd9V4RYL1mf9/gW4esqxxUypyBM2Xkz4NNEifrRoDUR3B3vRJggmlKAVMqfadRNtT8UFGra8J
QkWuJBoamblCs8RT6BAw2Jsmz9iYOiSSlrvMR5fu6dh1gs9iR+h7WoyOxSVdWE7kIrkLNJ91Xj09
obokJ+t7Nw+Ez5/gHhe6EQcCvKLeresc2dRsX5byon7jZEKtaax3FXkMmPfd62rxLQZ+Fucj7WLT
J1isftAB2wnyNmCXQXLBrLXIdFBYplyTAZ/E5nFNsISbAdHLnNQcQVHK+18Q3fxQQo22T+2NHJrK
2DXGUgWtICYyFv+d7R5pJfdAOkbK0hxdrduYYnGJKndCrMIAvSXfMAxDkwjjAzTWebK1AIbWW7kD
jQUxARTuPI6e0HDKv2d2cdTCL4Ns+n9bDLEtIDxHVq6JxUos+jEWl3maJQHd/pVdRHWLbPAi9x43
JWGfctdqnNa6GnjufMNWzDuKSKPNI1g2d8TtJ6iGW3JOCB9TvT36xz1zfV/q9o2fEgaOwYpgDPu7
RHhaB+iHe0D/8twh+TbXMz/jiTVRa3EH5T4G78ixcDvw0iaYANOk2Uqaw5fofCT7RCQVgZEP7KSt
Y68RY3+7a7sQ90nQ4qCsurIW9+kQCtAMHMPtF99PRDZkVqqXvQzz6UihEEVzOEkFzkgY0TlJTuSJ
/3Uc2WYsw1lY6O0XIAoqvzSwiilhwh+ClE62E2soX2VTmb11C6BNdE4iXlEktCztY/2qaTISLQyu
Dh5y4GRtW4EoL+qAFSjePDp9zKa2KmZJjRoqyhBVIufHGhvJKs9jYcqwle4htaNb6Bj4B+YTsmpD
tBwmMMKIzWppBZtzEbKKb2MaPW8+63C/cDQh56a6r5bCm3fOJXeQupRpGynM+NAkia/eA83DR6le
X7t1QTY31Gl6COLO5eFfasVjPLiIbDSH8/2eXeJ4T37gzXVtsDAKyc670df1dnYzPOxTqO3j4I1T
WONqN8vdaGAkaxgY1zQjjsBIosrfU1RuS1hGyJtIWK+vfBtZsEvqj4J0kSdVqTM9uNdDoo2sySn9
MrbND2CrdedqA1NIZ8xrL2tRFlV8k2MooV0oDXaT15WxCdch826ZOYzKeNVxEv+Qi9sRtSU/nZMX
hQFJcO1pLnlKcc2yBX1pOVXzf5b587E/DFFMC2rnS8T25oxI95Ro5kVwdkuKWNV0hGfwPYDRYbxF
dqg7V9Fehjov442UAwHymgwWmGzaNFYCn/PcLFCJ7/jHQfuK8FmMXtnCbObj6n4VZTle9JOrNS+z
/0164YCgNchhH22SW+sjGAP9aHdpC91Ru30mzRAhzCvS4fPQ/qseqj0VW3OAeV53ANOsSEietNgn
s4BoirA27pc9aTcCK18e023j7M/LT3vv6ZFCHMw4jZBxObod0rPiaPgnLbAtLbeOYNJcVU4CwuuU
13zbAdsaepucaI6RijqHmmtDXSYsL2h42mk87W0CXMyXo3Po5hcZD4FiDbyMBeBInsKrMFFCIQ1M
oUCQL/xAYknKM7ilpIqMmkUvv7FtOV40DZpebP6A1jtsTh82/IBk4nndD/ZOUpaUZwE/3lDN4e+0
xQ8361LzrK0Sr4utIEnioUKAZ3d2YiWH/70E/aqdopGnH78YWlOOZCiaCYWdjl7wwaJ8JkJPU7OA
86LLA6yJEyOxz7cenQutQltFTAgUCsC45BxLi/VIXs5cabpd+swcUDXnyEnxsoxzQ3MuCQJV2cTV
xUtbGVx0eassXy9vWXGWNzhbZ354GalXdLOzvQDl2aD+JXr3v29QuersxKJJ8G9PifOww00nuGc4
yK10Rg/t+kEeGjkghLdHUYA4rZo6Fadi5fm5/cNQJuI/QKE//lt8GBfuf+corph6Lv0TPY20I2k8
MFHaJOg9+x66JeFCkAXGuwJvg0oLtCiJkG/8Q4uOqw7WtPe1I9XBwQCa0p7awlZPw8kI247eg4YQ
rX3DIca8aps7YiEQEHqUi1OCD3a+MOaG56l0bSTNdyZikBip0wZrsv2wyeqE/47ZokUd31HWCDUw
JZPpfGAtpt1EZ21ZAaI3p0WRGiad7G508G/Xkt4LBeZGzF6kjK1DfwMzn2MP1YMgk0RF3MYE3nzi
+6JZVjdExOZioaI4EsBPYvlH9leLhvw6omnaE7sVjbQ1paYKJLmrp6R7dpHd1pfnWjlzEdSq2OAc
+WQfTuAU0eaVwAlGNy1dk+4BNqnak+fo+tzYGGW+e4aNFOlCofXvpy4IgcapGiYJyXhzGtHYJtqH
LyGXrb+Kf7wcz5TJK+tpXJUiZADUosoEsjB5CSsa4pc4C2fBzrM/mLemi4D51jITIVi1AkgXWkQA
z5nFU1GmtkQ0G/dZtUjEYVlt1Piux6N1oOd0IgSo+8EffJILEFb0FTywMzIHJc2vNN4pQZR7dZU2
HlUc8a12rOUBwL0hvPJX0Ku0D2y1ifGVGSPW6/7rWbu8TIHmDnLOoCO6lOxm3oWnxw7DA6jZCLQ8
AHFfSVCUCmH+jUwZFOEIp43LNG3LsEJ/Ga5w7jsC+VB24O+IJtxhdrwX8MBhghr3ql8Ou6TJM24u
TGOlIaD7Gl5b+kthNYok/KqX27QQ87uoS3NNATaDpceFANaH7f5p7LiH3QAP3L5MHzDY2mPSLVgy
sooaFbimA3wB9GwFKf2ZhL9unO0TMvV4zRg657q7NhOLzO14vpgcCppQ0apIvTFFShNME24NocGj
koJzT3lwT4vF49TvGiEOotxe+qAkdjaHtcr+ogIIzvxtXQ2OkI2XXDfWPdzLvR2kkyogR4GLBp9l
c3Whm1xIu70HqBIeaG36ffW4MaoZXdANdF0xUYE/5QKcDxmFhYOOMTWO/iV0+qMwdS6gewmxWCF+
H+2ITVdWVkudqXkl64YeMSh8dcDvWFLGR9pGawlgOd+3ma1bp9rGE2IpdEl91C4oTX0FCxLjHaWa
LAAT7gIZdT3JNDXPOfxgEkBTWm7UIdUwFHa9A5Iz4xwF5w+tmiWsvTv5w2VOz0g17l7HstW/3Aza
4hbs6uQnMHNDYniM1CZ/Mo+7eiY/TbEWEacqerNKeCuOGaq6RaZAhwz152hlbifV6oUaSUmyQxto
UcSBNhi62IOTlVXKbGDJmrnFnAIHYwtGP8vJisrWx1y2E8p5PQit+PdKSB4qcRpNp1QTKyNBzwC9
lx5tVChBeWgPL/GNNEKbHYD526y7Ir5fUYOxhU+QYoaLRYG/XCHZk1MTSq9Ew+CxXk/YL3MQyOzW
LMC+OPVAIpAgYQ9jVqtmQSmd/oXx8nFVY0hz+lSY8uzQcwuYFk4TDUHs2JUdbmS5ZqHZpDWE2Qr3
n5QL3wWiDOB+GGXwdTT+tIbNu15l9/4/1GWSO1WofcfQgj8N4by/ox9bwdww49bH98LEbBHaa7Cc
01sUiYmTMT72ibprSXnctvnLENMx7L//ZqB+QvzuzThlrBUp5JBAiuuBe1PXb/MTGc8G6OBKYHQh
zQ7v/vFLax58UlGcehvXQDI9WBd57xtGHK1v2zDLN8XbQIj0aAhA34YbiuS0Xxohtd+adSOzFx/O
GZ91AGZVoS+w+Yz3WDbxTCbUSGeIX3LYGVlSvkdm7cJh7eZDQTYi+g9F7VEynG8WYkRQ1ekZkNh3
ThtxooWuw484vU3y8sgkxLlnfiYFgWsw9SNaRkcTKCPHUIkCmHWTGqZqniBYfFQwz8LHKfC0RdK3
3wGpJdIzCCOYbuWWUWr7Uq9huI/upzwAxgplCCyddC6joSmU/qys1XM0bkABX8MJMBlxIPvahOdH
N1nZfWsz0KPCdFU2xUtN3SRKp7G8Fiybrh8TcK/0LykYTjH4WvW/BRm0uUyjZCLva6ELtuzD3hsM
Txzh+JZ+PumsY+tSxvukiWi4zs6R98wBtb21NsIomrt4IibctewwCxR9EV612ry7/wjFhneSwE7n
KdCADiVOpt0UmN9fRcVG5j4MQitbh2YzSq+/ADOM5u7MZ5c+EHdClUk6/Cp7aWR5GSo2OYKvgMI+
ZB9kYzARhUtBT3oQi9S8q4vWmaWUyYjpKdxclSNSpaHSTngU1sCLq8n57ApMwr2QeZwcWPCzgy/8
OWKDjgFJNqWoUjXg8qERblqrTY6uMm4FinUMm6pvScKnRsH6AgZZQCB5kX+CRwpV6c9t0HesShjV
AOQC7BmJeQGwgGGpN/y1QRXvSOvp8jBDkPHoqZmKFHD6wklFxgeGYbHAoTm3PrI7EM+VEqoV/iZ/
1+L6229W1GgUUbhH+tsFlavw0HG2g7QrZhvd7lSrQ26lFZEV7h5qH69Ju+ED1NS7HzLRD4DguQ5Z
hvMdpECIRSGt0rZWEjfk/DPa3uZmZHjExvrR3yqbDS3RUo0raEwRWSh8chNdGub3aRVbLFP+Mqiy
K+ku8DDj2v3zVvqtsLRm96QSdZLlytksOflyqmXvKCiTTRI9rQHBbO8eqh0fuAJ/pMA9+mzaMtW4
wLW8R2bUbGbU7g/SywzyHtF5C1AGm4W0ztwd/nh9XM0xw9MIzxHsXuP799XQB/2Qzf1Cw+iJ5ZjK
JRt977I0IOuhLqkfWMs10j5V8EFUVR96ynepp4Oii+zag4tGBGfVR/Y34yW1a82kE+lXpFLTLM7N
qOgJysXtn2NrIx7y5clgCPwmE8cpv4fFydSWXy3Rn25nSC05cOv7kwLSalAxYS0xFM8KhzYXzVZn
dfT5qQIyjEjgdF8qHNmdOWcp8CgCbW+d3bgp47My3DiggUYHLtzh8XVpo60VMnPP8I4Hjj1NMuhV
ir4dB7qyhmA634Ev3q9grs74iJQXzsHcSMBab4uRQd3QJeBH/kSSnRoQD+lw/XRMcV8YexCeKTHM
TXo3H3atwmCT1WHvql0zTZW9aWVR2v6pB2VENoQZ6WpaWT1jropqEGfuGqGS1NnAwpYL05qHY5JY
PPiWGRCMdfexK5goaaViksxBuniq6BFDYgsNQeuSDFQ29sVkG43xpj/Ngs3IojqT99/TKY0xVU5K
0JKx5WBEWQPN4rLEnrXuYtH7JbpBvclL+JZa2tWiVJEbmBIopFHTKZ57Uoxg2ZqP8DIkfM7Uy3bb
qIwX4y8ABt7aShoKiNos/46zV5ziDtT/DE0kHISS5PRPY9su7l4BzQBBCkwAFBpjO9k3KrlxJMgw
mFziTczi+jOVe5wUY8YPy3PX9c6BUSom6xXiARbZRi7/s5i5bdmT1vVfr8b+4rYAfLXVxAoOzRCH
HEdPJPc9YaGIKX3Khf/KIkrcvS2pck/OFwJ474rOQkqZ4faUDwmg4vjp3KmiVFPbZ/Keuc5obzOo
raGOvDd6NA/Kuz9FOGPF/RjSuK2P+jBHYhMlkz6j2oRjuOQBe8680dZkDMimGy+RB95yegqBukyL
CfXMe8xY1SRMZjNJuFF4AIPTyNS5L+COo4I9q9YMc00z504eEvG7PMYkDywR9XCF7Hg7mmfU9QoU
ECwh/CkuZdFC9Y3XsW8T2afeblKmkgcmqm+7gGGK9DJihlP+OzwQ/ZNTjsJvgHEvFolNcYq72qAl
3vyJ2RS5fjnrFjcjtgbmtUwmmymK+xJ89DQuIn8tmPQfcz3uF3B2La5E05kov8/qHDT2hCqGQz8C
NxPESzU3cFPm2uKDBprh3xq9Ay1a6tzYn6iETSIf5IQj8ANVSoM5M9aMJb6kRyoyLK5YsLDnBffj
bhZYXbDm3LXUr3IOkOQxI/sRVz1xRHBrbyGEgGX7reQs0hKr+F4/+hbNqibQprxfKGcmmOcQ4tsP
1ZgZhZAxXISDixjcDTHq8ccrsnO/hS5r7BeK6MxYDPObMsHtqLHr53kua5MrNmDbWwvxnq15Xlvg
KLAoMXReFdqE7RZfWeVQppxD2JaJacfIDV2vvKEgkabmy8+j2bW6s0CfCBt4+8bZFqiqmJbB1/1c
tn0AeGC4FBBN9KqhjR191kTsB485qj9/8J8aQ94upaJRn1EIUktwnpLx1YLG0PHb4ieVlN1oE/YH
Dcl+wjOvJGz5cN3qzhToZi0GinGm/Sax7rrjDYUPWLwoaRFlgSz1M1hAgAhpIztfIjgA6nTTw8Ol
8gm48dYhe8NsQiaCM5WZ8DKN9Q8SUMjqQJOIrNIZwsVwLcV1m05xGOvQnWFueX+R8+ekVvUClTv/
qJve7p+7q07VbOG/+3EUh92UbTRGr+hkgVlulbu8ALgfrqiOIc5AIUSwjdVWBGak/FOqZFNIZ6z9
mmOhfosgjBbvS/l2HhNk41reCM4sDZrFPTdZuyUgJP8W7kgf+dGSMXPKY5kY7niRPU0sWlqesGYa
COSjiklk20p174pt7mb1BvR8pWcAm/wpymeyojfjjQqjxkY9M7Ku0HZTA66Ivj3d5QWhazkNktRf
dHB6yngmEHKfJdhrh2atZNdG6wwiB0qqN4ll5SuKFKHqelaZD4bylhL+CBoshvCCyj2AcpLT59YO
mm5JKaXQ8pESfteaIzYRl5mrdfSMzLEC1Mtik1u7rJWuBc6t3OcpvzEBbZJ+ie+T4HK/yEbfkArY
US0Bbs4POya0M7oo+zNhBVuYFt2AOqCrNiHc+7duaUM+gzwusJc8IuqudzMxRe5We5BrUW7sXZGg
9qKz3QApipoG5KJD6+tzUu+9MGADCfMprZqCpypJq+B0x0USVRLVEa7taq3X9hy7Olt4n7pqlPef
v5Sn4srjdNXR3tV90aR3OlKGbujmm2ylQzncBibY3vJ33c3XTxTLUl1QX+EKVlN8f6MuomeBl9Yl
2Ecvejgj2jykiTOH96J6UBjp0AZcIPD//jpXY+coSfxocS3Y4OnKMgO42ZRLpp3ekGghEPBktDzD
uuh2j86cUTGi/sLEKK7dcghNvWvBw0kx1jKg96xmgwINQSwJB4VYuuC40pdehDUHzN4njSiOSHWT
OOt7aFjPJbOvQTXJNghPfyKx8Ho6a7bqnd5l6M7inOZ/ZSdhwR+TuiuGyY+mGpncGMBVX3Ni8AJ1
vyAIwt5+QtUCRZbcJNNJUl+qVucBP0o7iJe6xqOoSdy4Dw1wCXj+MPb8Elott6uY8vSLbyXAbGvQ
NeYGg8+aSqGZlImPBH/90pa1mQiZ0ty0/3HAYXzMDkECEsodPYsaHB61ImaAsaau+QxgHlQsnY9A
CNuONE2g5QmmL+Qd+XkMzJ0Dx3r2j5Tr3e0g1OzxqMWCBf/c6bIeu5WFR0NTQm0X9UziyKD0slSz
GefsqNzAVbe8JUon9FMuVFDpAJuqXwNsYBXAHE0UWZ0YulhvcXURdEAa9ub94qBs9FmaQFnDKRiv
HDLf/eok8FA6Qr0twLAh7GH+39WP4lEmccAwNm4Tw55cHrknO1Fa/NSutTqVrdBoXgEeAg8Sm4/S
fIGvGnY9EiQ5HxvxcN6d/TuxCPsbLPNpt/IOieIgDo4K2B9sfMMYO45WJef277p1Q8RSPIpG4Vwa
AolU9zWCndG+7zm3EOQHTXtyssJ2Enh5gvl+FDUePOfTRQc5ZTxh8bh+Vni99UHb5zwD2vJ2mHOl
urPe68GcK3S4Xmjk6UzSCp370Y90tfwFP7K//kuxcITd7IatbcKaCyrS6vc0K5S8Fm77J/KOtGYO
rH6HifbVl9Uh9SegohwPav0CtsIobtIqYViHzG3sJmrt6OyR6hVOtTCmHLwcSXEla7TVF+dF5HLA
yb70/jbfbkMwZg9m57m1EMoxViBQtrlxz26AAXl+VQq6AFZOkAwHs9EnfRD/n3mLpni0OuKV0yGS
67MlbDekej3lgWdsYomyVwb+YekSrL8se0BEAQs3xMFYHZlwNz4eg3OOcBjsl8o++1f7Pbb00qlQ
1vTl6nj3rtI3UguOh8dTnPjk7LcqHWFPGRDm4B0bM/pUUjuC0UtAbFgBuRpPsVW87jO5AawjuOSL
WbUUDHm/gwrbwY4yUK1iwvepzLgRb/uTwNjAv/yGsDGqnFvp9rP9yxtZC/1N34e61IEUQ03wXpwQ
vIVwCL24qShQ+YobA+MRbXacS7nA8oOAEbWDuToIiwABPEWBhEXgcOeElAXNTtLF5eramK6p4bGi
wiT4+gQfCe5Bqg4VTgm1Pol8mZ7rV2Pu9udJQzMtJQlBQYhC4LQ0f/pZ6EN/Jx7WEeHUAJAhvQhA
DqMhDTeBIUpVzsX4xAk8lP1Gax/DIYTaTfvFSU4HM/6EkljQkFEjJINDh1+3DtuutZIABFtGEDj+
S0JyQZvINnmqfQBWezIe+qmecTW/zSQtsdV9poFGkTdpUoKjbsR5LhDHIZV8jjOYCdCB0OosFRl/
v3PRpoas4gQsyjAIfgA5nPleYvl3/QaPCjcHWit4kHQM5yv3/Rb2w/cDzLhn6OV/kg6PysmAo52i
PaO2gkiqeLrCIJMViM/swffK5rt5hBkQIaZDSVtarYBfRU33RBNHBPm8PefOSvPe+mCWz8i6pAEg
pHnnhJ0A7wDjBeE9yB9s7wpEy+kGhtGuEMHGmOx+nupzqRGRdtpivbzts7l5xizHYerjVum7EdeV
XYjv9BjgoX0wEajtXOzHXzPCudS6L33sKfEsO9g0Bja7x7hi1x/8sOyQj0b/+j+W58B3uRoJ1aEQ
1N3kcfrYRcbQ39dyHat1Vm63PklmZKquso3MXKdz0wTLhhpicevxIPqzCS7Im3gZERqbRfgP3eRY
6+P2X4csdp16FHPRErSichGlJYcBOVlfPznRymu5LivRT+5eqSTEUB7qf+NshxzY6DPO4H/PL8cU
Gk1MjuX4WyGHcziJqK0o9gRobpHFgaQscOWboOq3Ig7DBqZvfVOpREY370QjTgNrXal1l41ZmHEG
RQ5fLyRgu2xvLG/8xB4GZsLP7+x1AeEY3FBYHAtWAZYwLxpflLFui44ucuEANVOGkW8kA5awfPj0
D6q1tBqJ8DB9zOa3Tplw0J1TjrSMDDEVujeIBIIMJ/0khxxgeDv4GKYW++bX84mzyiWnpd0JILMR
JrtXPVU8phMjiBzCZZdexYCVuPKCqnLKJ+gy0sbWTubmD83VGArzfQfGVKsnVcjamrs37DA0qRLS
H+WD2S9BgDu2S6Rs6EW6HYsh+PvUIlUkTC4MJNzCQHAgb2+QU6yNfiWrT4JGaIX23X5UrhD3Awts
5S+xK7PwmvaEqgaSpCO0cgtEoLYRd3TstC7dDmgiWW+F7mHZNgjtvWMXp9/r5q0j+ON1LIGlqE0Y
CklZC3X7M31QwK0W7WrabLC6PL9SY3fp5kgyRBxfRWHkUgmBaf43+iQyflrCibD+OOVLVHaHLMKt
1gMVVFuCIiLkbzEiAZma9csmri0ZHeoAijKZgK5B6PXWHlMsYNj16fb6k5qhPJ60MSb+i6aUFqxf
nYAoK4RbX2aoJyLtAjhyaneFx8jhZ+FFPQjx+R4LYLsWBak7RRmiXWxcf3Psg7tD9B7OYnWcq7de
iamO/83cJN+cnsXiueQXWLmuhlVQv4+KpNoeQVgcIf001wYkgpUL2S6cfzg4BD/7fR7SSmJzaXXK
Ns77Qeu0wiGxKXrwNEdhdGsRr/bRe2Z1wOdhmYxUL11WRrbUczEZLf+uwMRAADFi0ZkXmux+OC99
VtGOqSZOl4Oz7VWDXjq8D4cHSUDaZNV9f28y8SihR3eu96pmAdypXLzO0exEYoiACOgi2r+HQLNw
TKkkhlNdAonrcRrtLRnxMI2PIHRhcb+Xp0shiYnvGb+AAxmtC5wy0i2SIGO6l+XfYNnJZlvbtEX3
yxElGXlx60WVMyCXiQn+fDab5Uzi4RlKkx8i2fOwh9voYU8xJeviK0tGxLNXP/IU1ffntGrU9gdW
3N2DMyTcJTz957Da86V3xdr4TZCe/HnkxGmoIpa7mALpk24XWtBTptlt0TV7QdSUXoavVM0mVhmr
hosmWghJlX1Y7BSZ/M0pdlJk7eins18VzBi/wZTCL9ZkbdgZ/7oR3i9MDuESCYZnrsn0/lTbfuIV
MEXptjrQ2wZ/lJeldPEoUr+dHPbVuaikVPY5v7ZERMJZvfKemdzYqhkgJUhH0Nk9TilHRboYaepa
pH125f0l24JNdLJM1rOwDEm10gRItDezDTGK4czDBWrLvgs+TkSeWlRhaugoKBwVbQ6FFMivHeq7
sdobF6OiYMWqmC6ZbKxNVC81CwTFwhp5STLXyq/aCYjM/37gq5M5CrGtixXHJcQuYn9NdR3Vbky7
1pAuGUSwrwO62VwVyYWMKKxZYq9lwGqptOtoOCgiMyhVIN5hr8flzYJ/TL4WfXLP4ApZAWj40FBk
9QGxgORVYjOjasXrp7bYfOGvzum/ZrJsy3JCzh3YEApbRMDbhliXVzSTAMmYlcWHnqyB4H6FMZTf
X9XaD4FK3VBbaxUnzU5KiAVVEvBkJMVYZGHJ1TeBIcwlNFKhTtr9yn96DB1z5Np6U3D9TEl7llRK
Sqws7klWBTkbSfpyX7PhGodMEXI/9jz4JpHTv+5wkNVic7oQMtHIJZ3rViKt/FJB+SjNb6iL2VW/
P9TkWoB+13DQOResTgNrSnGqpLMxtMu98YmgNyuPJkjNZs5q7k8oexEGT8b4aIJZbWwb3g2fZmnG
q9k6jApUzZQBudO5novY2YPpE9erOhqkbZp+dKg66vWoCdGjzNL3kS5cj2vGUR6QbI3W235QjBqS
EGKLv60jwxdyqBi2fX4S7LSGmSncXVxNPknk6U+BvRKS3fy0TPi6JVERMgUERKeJjTX1xFDHvZAQ
DK9F5PZ3K5WuuUK93P27vuq+2C+Cerb9ub+JwFjQSwHsxubnmegXU9CxtoiCbEJCFgSCwvgT9Y/l
bE4/B/kfvgQRepQGxFk7CaMTQO3lBRj6cnhMk6nb16nPEY2LRvs8qYdQQCTdkgROTmArf0Ol5RTN
Ts3H0BRRtgLxP72h8dnye8+r0lbkNg/c4oycbfMXvmagYP2HEGSopeiO1eVDl6cu1RAQjvTSzF37
igsdtDOtDDZhoi2Tc8djYSTlSMswe1qgi+34vJw05+r/H8SFn+mW5eTBIcn1SSWO5x7laJi+AQOr
icepfMY8S1bPAUnmJ5eSqB7CO0IC8jBdIcxnDH0oUc1cJJ+EMhOpY11RJ+jPUb55W9q3ZmCfXlU1
BuBoqcf4rrxGSSgtf0BW+C6oIWcbKeYi+4ir2RYdDb1OqmXDe8BqTD+3Y2O9hQ853Fwg6B/04INb
d4dS+4MXR7vVqrdzEd1FZXUbYRV6g/yHJ4mYQ2V1G/n92MfL3JXCkXbSBdBPPdmlZTVpS3eRHqUW
cTsf8RCGTaToo9xvkM0EsPrZyauBrOYfGkUKo/NWomhv5cyn7oR9ON8MCbmSMOBRkUuzXADDXNtQ
hNudxDHL7Uhs74cXWBYF8ajNIYgORGJEXJROoXhd8FC110zhIjb8RULqZu90fkJZhQ0R1vNFikU5
F+9LbOpMH6fOYDLOdND8wntoldWSoxoXZ6eXs0RSDOuaAO/ikFbyUqD0gdlg4kLSbf6i3ybSmK/K
QiOeeZfaf87YM0nugarxjBLbmY4h6ujDOTMSwx5AThI/wLH/lSSuQx6XKb9mwkNGrplUnn9YBjjS
ko36pl8jgE7NgMD9XVSXoq3sbotEVbL7FRH25af4/qyD9UiWIl9VulVfGH+/j89L0+vz/6oy/Lne
4Rm4wQBDWCT76pQVHUuffuY7QtNfKZ4VTqBezwQ17Thq/hNIYPoaEPBgsXS8EdeXXVM8BJ3tR4/S
e0qB3MWNahkFN3LKxQmRZHFgncJ6YOGIh/nS9f6DCsTSFrHBRFbhSKhqn4noXaQL8logy1kXxhKZ
qa2BJMz2DiUhuYefD9aNtpg3Efyjx6apaX8qZjYi3NXdQ5tj8KzKb93O9rjElENlHKesgAvkL10N
txMmi2XolJD+ORtvRcWuCHyGNFPMr4onNBLZ3yHK3YdWGr/UefwTda5F141XA8ykVYjJQWP/OIaT
ldq4X2aM8wgeMJSeK5lneCJNhYU4EboRL4ygGYwSLXGzE1uehVkyga/lfILhEbh4U8Aoq4tCiWDl
mHZvqGUFyVW2h3GonO1ChAHN740lRhwHtkVx/naKHHmqj/0n6iDqEr0T/MpYMnaGR8UvP7fPu/aB
1u5Sje5+okzWMjs5HcD10E62pGIi4AmMg3dRDoICqNYpyBi+SJHSAi3hw7vBAtXaEaKE6onrN5AR
Aw9/tAETtxtmddYEzmIFaEmN1TqDoYFD7YIB7DHsXqEk/b3G62AXNqBQleb2Wkd3q5RXnjvL1Vfs
Z3OJIK1Z/w1Bjf5AxG1IDHRDuvuKzv0ZDQ5ZRiEy8NkPnRqlqHByAvNSucisV/xwao0Gn2RN+zBV
6Igm8mzAqDn++vUrxsx9qaD3FSdQdX+lhrKtg2vnHhcMGAmMHz3TT7Re3FRbJ6RTHKHJdHn5ZaP5
dMOJ4GmHIKm0e51LRbqLrtUpuIirCYO5Ehz220QstjGlNTdfbl9sfQUdNTaclYNDDtwcctmf/tCs
77771gxESTGUnx1BMVTTyWUtKgEADh9p/bOuGGxkB4UhvTEMf7vJ9jy59igJ29hxnZZ9PcYeiUb2
g9pWc9SNS6jHl394THazFcVqcl6sQtowNCq2oCArOxyLmYXauBx7JKQGuB/+ZG73VY0zazPR+4Wk
5zTss77Hc7ZRvzmQ3lBq9DBndlPsLEFu8Em8STrZvu60T/wF2N7wZDi/8I4raZlxVtaaKxjk9WTQ
f4H+fOBZoKZMjpgupi9jAMVc+f6PLCaK4an7w6vfhEGHHkLr0NJESfYjLytYsk5paATQ1lqq1SKC
GDiuZFoQNS5C0eDp8yCjVHo/HgfJTLAm6vPs6ScMTV37v8q/bEtqfylCHusNpUm71gS7LLeBBoF1
SUaagMb3Kixbk1bxNJGsNj8G+d8iQu4ye/zhsb0yvKmx1JRXIRthbZThfTOWDLYd+SWRW2gZLMpu
u1cnPLvglHz8vDhlfVb08OGmssKghiL0OJe6OqnCJ/GOiVaYojTu1C8GNrHiCvJoivPz2hjKkREr
DHOmUdZ7IUeZZktpv5V1S4wPtrAqNR6S6CJ9SjYxzNcm7PCBx+vTtjwXG2/VEC+7Refgw1zUH6eo
EeyKOQ8JFpzdJIwhIkKdKjdfVZei9dE+ncP9pOYHob8kqu3sDaNuhTp/nHSe6oyetbURdAo4QuoH
N6cSb6Bw/pMswz8ob1PC6+NUdgx0bi8D09+8m0hO3GikO4RqSgNIsVWOgG7VQRHB9kAMqt85tDeY
cBpwXYJ4A3VUrgzA45opJZCxjYWC7eUH4uLim8AMImL8DBuM+lfua7WQ9ZTMbSoMw+M/t/LiQJ5/
r+SsTDToRDnX0lkL9Q6u66a78LJcf0vBnWU8WNz2cIFPEaerYDtlDOji/Kh4YSBsV0AXGrU0+K9s
kwBI+b+9FkzeRUTqPCgATHe3IpIRJNFyDRmJJRaXevWsqX5cVme6X173s0LzHqPxAbJz8m2iSRQT
7dL+jUA3xi3iTMN9ilpw0YAgp1tWSjLvLbgfjWUzgpmfvyfX/lAWBr9eD4kxwGCxaw7wwEdMEuQ8
vLPi0ic9sJrl4S9SuP4Ngmpn4FfiGM2JgxXQ8gY/wXZiwPO8RguftR5aIuCa7jvMf935VDX+HZFL
9jtV0rGewvEM4gghWonbu664trZG6yT1fYgLTEqmvPXsEHpd59k9IwNa6nVbbpJWTAYLDZF0KOaV
f+Fw31B+oSBwr/U7QRVVH3SPlqxLCxnMl3tsBwHildcjlG47wuNqp1a5ccUi1CGwi+0oFeN6tVhS
GZ22hNPmw63FwqyJfjPULEAzD2NTDnisdnoa8mkHklR6lL33gBlM1g1N4YedRs9GqX+Q4b2K64Wh
Pdh1VbjsTqnw5YJa71hRkFvktmVQX7gMs7PgJXSiaonUEhkjZ5RoMSZOOlOJ3K1Y1z5pCqmjnBOA
bYpi5ZMtB/s0Zaz0a00+0J1Vs9Wt3GBADlPFbCtsbv5TpYJVUN9SHL8SSsQdbxf25bksKs5A7vuM
kKSF32xFtYUKOManpuu3jeQphbYg0gBMCrAX8HWF6ufm4iPlc8Fzg6EtYYTGwwK5a1VTs6DL11hu
WmJ0TtGztK1VGRJdPcylYK1MsBYZ3uRQWC9qXi6FKAY36dCnOangV97WzjKDYWYDVlKR4L4Um1xw
KaIf81DPVFi3YN7Qsl4x7HD4ick3PKLBY+xEWIym5/qg8oj8rhZGJzlnPX1IZLYWDDM04PSFvzWz
QGRtiLHmOOtdS70VByFB9ILZuXZ02OyL2Zl6VyIp5UziyrTKd8z22w3aeG7x8SyrTOC+DEQtgq1k
icBVjINK6xtf7QDfLhHKCiSlVIXpvMlGBWNHhxnpciShN9u5qiAb+2eInouJpFexCJtteMbGQB7Q
YWYuFfixSnHd8m3U0dt4qsw9yqbQT+17qkZ6HWfzMMBvvnz5ro6JS6Rhbyxdu5OKf7C4oWjsumZR
ouZrMH+73L9JNDqGW+wARW0P6kD0pv8XrhjHUuBPSLl+9ly+GGaXtyh8gM5oqqEqYNSFMs2DaVv0
7y5FYlGSoLykmUjy7Gep0vuB82VjlBnunK6VTB5aetx7+csDuI1ah65EQHM3F1PIYq9xoLTlVUyh
+l+L7c59ldW47S9CzTjlX5Gf0gxdgzoPxeN8bpetzeOv7Exd8h8HkhFHq6Pj3POnXb7NcjWGN5q3
lqsuAYvBdA8gClwCJ+vELT6j6kmfsy/nAJDbWtf9XId3MzryyqHiUYkFU1mEsokRkE+wen7EoDpZ
Ckmf0A9/9nZuvNAdLL5Ky8LEec4vA9nBC1ZaornRDiD//XQq6bJ70gsPN9FMasOAWvgJYSBoY09c
GbAYzs8UVkxEewds0TqC4FMYtqKt1EpTHlo40q1WxbkWIuFV6Bjfc1diZOZTAnNWaCluT4oBfZx5
4txVM/L/PTm/pVi1jXvqOviyi+qW++Ammino0ug7hpSE6Vz1VoC0VTPTboWrqsSwq38QxBMMJtVa
iBOeL5HMVGFUO5lyn/x/28+eZ38kokY6MTzDLC20z7IRNg+zWRHSkP7EWgenqCTbfDzH8WTUJTO3
9g/1ywTMvC6AyUss8s2DvalNYJPrDpdPCX/QiLKjpFp6+ZrXZiYr0wA5t5qdQezje05mM6j7JYXJ
asvFx/+EIiOZxadhF6RAjWjpSbgEU84rXWie452MEkz688aU/TzopwkWtdE7xl8EkJcnpIpqaaZf
DruhzkrGETabgZXsc1JoneL3/2/F7fGjxxra4ZQ0AeS1OXaOYJl/cQZFlUhVFYZdGMyPc6G2iRkA
ZtQK+fVpPa6t4vXktZAVizcNfVjc7C3DgG1I8WvRdQAAkXDFwIGfbvf6wShwVB68cc8cDsPyhiKv
7L1bOl+bW1mgbdya+dUZ963oVktTdJ4TF0CZWLYDVnljVhlWIvsgavRIn/VCoetsp30r6iPpp9b6
vmWKy6aeoheKzyNuLY8X+yzEJR0EIwr6N9y2GxU0AemXd0QS8aQxzfPzvQykCwb8b0wEDT7FxSs3
lCbFC5OWQXZxY+bPF+0/O6svRJM+y874lxMKuo5G3tT8QkdZdhHC/7Smb+5uwKZEPfebwG64cTHQ
HcZnSxdl9gaAFVqJNIhZBdecQ4CvimA6YzBdsa4izrMyzqsIJGYB6tCa2FqPHy3vwr1KYEQRZSTJ
RhFjPBqq6rBTZD3GRKSz77BTdDhcEouqVBKtVS+Wi7+tmLwyAqV7XFfnoMp1H4fFKhnb7L4pX+es
ZTGIpZkXMuYOP69eIVBcRt/OzkxAmXSQR6GK1IZl9r5zxLjGyWNU13viwVgQG90WvjpVesoGsU5T
fHGJ2E4tV/ReRtkpGhgAHT3qQgY6eidcVSuzNAwmaAgmmsXNZcAl5R1dfREW0LcjfjPj/7k+HQ8R
hYGi21UiONJHzFK5fedcM9W1U7PF0hl7jjJ0RXjpQ+/hnLf/t4gn1sfR6srFEehoWIzogxe7V1Pj
ImED7kSM0rmJoWNm2JQPDJtHVR+cEqXEVXiP1F5IrBBHh8G0YYvhqOodwXvo2szO4U4hchS2V8+F
Jvq2FXUgpDzt6MTIGezmCoStwxFl0N4MbT5T13C2qOBCLGBZT6HJfNVki0oTN+OE0YHbW8lJSRb3
V0mblUHaOn7WqLE+E6F0trLo9spI3chkuHTOQYSzcPPgscoAl0c/XpVGKd0hMg/2TblfgXhUMs5F
npaCx4szfoCpmFjMn+AwzJOczYiFsuo7ppAIYYkJrxUgh0+Z0t7XEfXd/S4N3WTztooun8T6KyVb
SdBKJSydte8UCEPW2zKa7aZdsVcVsxY6ulfr1Br3euy3GxGh5RBB6CMhTukyKzDCDB9+vrorJHiR
F2/EY9Vo16aRpHOgBvXYJBV7PVdW/rd9ohuhbZ4ZE2te/BHbn595uFEW5ocUQMKNX/2G/V3PWOsp
c5DOjflw/ymp+ld9LlNRa7Gwjzfr5wWRuCE02XJCJIVSd7Lm6DJW8ZMgGD8P348rZcD9d2XG00XD
SlWMc6potrJU3j/pANJoucx0fRJaE7rX3y0oa7DK0Skrkyyv+NixMyptRlaPQu6yXDvo85IejG/+
tmNmephO0iY75rAYKMge3ehHA+1bIL/h8DFtY3ZoobRFrtz3WgGxDXGMt22857gn+9avOSdsgnEe
+mpa7kDOcUpgqSQ9Fi14C1RRApJDFhdkvX6M2eF6xH8e8Z2pQAZmSFvANBR8d11GSN+Y0kUlZYQn
jaPgb25kxvUYsdPRib776YaZKlFOjZTvtld2s0h8iBF3XVFAsuyCzkprlwk7s5Exqre4Gz20kYmF
cQzXWGPzo6aqv+vWB0OTQ0l79CXyujzVJ4UiXJ6Hdgt143jQpLwRl5f2e1eFDLoG1gnMpZbK/McV
+aUc6x1YlXYjYxvh4KqlofD8Ai8sSzhaNc5AXOmma7dSbvXSR7OIvxx55wLXtyA0cKb6EEWwgc6e
YYF3khJm+ceH5MkKltt0ttff4+2+YQfPddA6/BN73L4wobirlhiiDGfRlpv5xRGZwyDgV431LKYC
MTB2tmhjSzE8KQr7wl8kVegBuSciaPOf6X6DTsDLGs0Y7lkTd8PE4OgxCt7ALduJ8a5Vu6/zCKed
UK/Bu+4PlHStvZumdCNSMzlG8LMNzsgmC+53ad/T6fRC/jQ6Y/NjxDYYEBczguWu52ehX06lB4t8
LCQqHn0/Q+IKPkqv/Su2MIWtP0b6/GvG5lR2Ag/aha86wpyL4O3nrcHW6sY5zQ9tS+jm0B9l9ECT
xYnG+0aq3XCluHjQvsLU7Yld6n+4WyOnVr6ym55H2woYd9ZQ8ZMteBD/12zxyiGWrI/4eeIA35nP
cHgBxIwq+SsTeHiLJUE+vDfV9D1pdmQVh5CJcHAo4X3sTY+dVsGm0loi9fTLYjWRC55fr58yHP+C
Q2ifIlDnF7x8Pnujc1pc/zz4vLAm4PvttegKTbDexweWXoT0J7O0ZN2l8cquT3e+Hqr32CzQ09Cf
rBM/J8+cGn3/yvl7pWXfljKVOuV9wUCwroiGFCSzjjKXm7KI0EGcxZGNgc1jP1F46m1gmZzZ/e8L
E9BJ3hNbi1AqaywGfwq+stsJacm/MGy/01fRy2sFx6qu1q8KCjbkxySZMUYPucGXa5rkFfSTRWq8
aZ0Sc5dhWx6AEKsdQ1Ug0yR3gOmupUgu94F/P6mcbG9PZHZiECBjH3r0Ab0DAei5aUCZZVIkK/Jy
9nUQ1+9zb6vfvZ7OWbPg+5bBXhdR9AD8nLbP5zhgspWUsX3L+0ULfFtXWB8QQTqof9rixbtIlxv9
lcq9PHLL7NIPN4sn8Z/NjmDNqAMMMmjm0JQ/e+BjOT2yeN/+MrBHCLtA+CQ1P4wND3ajG7384xR5
7HYE7XhJxJYunIRgSjS4wvqhtNuPRzCaAcRqGPAiFER9uxzmp+DFVE9p057IRYmd1bK0wze4MeQw
+bFrJFH1Atre0itAv99vYxEU72HylIncf24E9ToGMHBT39QJjM1xaSAsSideM2UkUrNJRYnzbzg5
XqeeTiQPHUf1LU0+zdimhkRMoi6qHkHCOVEHvNRdiHuitL5Hi/tlOiTMdRnHqti6sj8n+6CN+rzp
FkwPrU9gLsC8pK/kF6aF0w5Oa/7ssnWk6PAEudPMBZ7uqujxNu5YIxyPjqHMIicjEOyF+oVXnrpl
xqD4uX6vdvpttjARL/aamYfu0WRo8LR9rxy7g8/cA11fx2bdlMwPmHuvCKw8yHahiSvy3p3mRLJg
9WgODAXSl9qVvgpPN4ceVuRdxwEIZ/lMzPLzkWh5qZa+6D0O5riZ+GgreRabT5/fCWPUxPz0zwvo
l1gRrW8V8OKZ3guREOcYUe42vmfl1vqN+/ioTGrpiJNH6DKJoRR4Q3eLiNVsEq6gaF3TLrFa5rgm
fSgE9uVIBlKyAX+8zmbsWeo6gPeWcppY8yv6yKKzSoT1uJoT9NhxH2kwaFCKY9D3BkgpPVJZZyfi
REilMbGmIRTuigiFrqHrCL2c0WO9VXwi2hR83HjIfFk0m8mRHzNr44IP+mhTWgII3upJObaHnb+1
t67inAGN4W0zrZ4h+Xz298eHc/QGZs2ROj9Yt+FJTQniS0Od0S6J7YpJiSOeZRNugi854WsuLvXZ
3nKEiBaYl6l4YSdeBVq+DOBh7qWV8VdmyqQNRoE0zaT4LOowVCZ3tjLeAxZaWMdrbBFeJtK0d+Wl
rQX4uOuc9T2IiAumuicKRbyJpTK3JNrBxqZk2yrfw+aAwBVjyPKKrII9gVzi3gePFXC80yX8cTLu
/46/b8OEvY6Kc86wjhDhhiz5q39lDtcG54SpY2V633vYM03qzB/lz7sjRH2jVyhfhVE65KjF+7Il
w4uBDLHbpI6ohMdHIXE8XiB0SVaEqlSHQh17NnRQ7daDoeGQ2f7xfMo0/GMxeCNwlbDVi6wSCUcl
HjwbHTu4KX32M49TFIqZJYAuCmdK3gYjFccV85O0wZQ0hGvnSIu08J8uvrKZuIV6NOWB3qgnrtjB
3ueA1J5u9fcaieNO7QKsIaIsFHcb+ZTpXSNLwJsyCxuTEmnEGuF1G8RyMSOqvYF8LuvWM6SH6dpc
VT4woUMT//kQfz1AcQW0ylqrlwzpUnW7hWm9inuLt9BFsBlT7Pt5KrUcIw1wLnfAByhmBulVuoTt
2LUZNPYFfO7fBpz+eO6pC2hA3Ry+2eAFviqDbMcOHmhalUiVVq9yylWxkiluOnWmhT7Ue00W07fP
5yRYldX5hKkf5TkMdrGa1zFDTo67rtHfrrPvaoVfSk3k186FLRx8Hijb7c5GrUWxFlP8Iut1P2Pp
dR/OHuv+SfqFoAOHWgKioinog8ISZKTBwem80Nm9Qei5H6lZrYwm6SHCrS6ZTuR5HfipTQJYngju
BYcyMOOdsfMfElLnzze3BP5pJaY6Su4RM/nvx1gsmT0ZPNT6mGjyXjx5+w1CxZNATtMH+m3Bgpk4
ZfUz1ma95UUK3pQ0q92CU8qwEtHYEo+g9tLau4E4so/Hz6bAsSXi7dMmQ+5V3xWwbpFOU/7COOoi
XIRKIZpu6V5aulbbC8/LX9NMFuOG6q1cIsP0sYM+3vSstw0tJn9gLGQusPY+taMEhdg8jWlCBAQ+
JPERDZeRJRZ34NoVXeq6+30lzd38WkFO/RPvV9c/QQc6Sopzs1yaYAKaKgMVDucN2zKBKg154ekU
95gnaPqKneIl/ny1yaQbPVHRz7skaZOj25acO86NAZU+Dv87O6jIFlaZr3xWfxTmtG/X1tvkt6KW
5HzgerC1uBM1kzSbTYlvcCde4fBgxC9xNRux5d6nkqy65/kI+De6sc9AozitfImJ8vTVnRNDXTvI
wCNNpBKQA+rBPRSsEpkfl4tINjEXo++YWokPjMK7XsPOO81Yw8fw6+xZ0zyT2S6ewBrh2yCcAE9A
0ry495/FyNYyOoWZm+S9jKki6gQuo+6Hj4u36uavqbKajH/tIkW2xgA7XkDgHJqw0UDtMQ5xOHvW
dbQZnJTdG/1OkuIWrO5yZGINH/6UuBpwnpq9cAVZc9cyHwfBHFcbWwH2bxURLkFPRzNFd5T31qqF
2vnnL3I8RPiyc2lVWgEZpnFXrWU9ETxa4FQBcGTmCWEem+u3U031e4bkK4f9LwHRlgMRy3TVFEvB
Lwo/xUn0VJwDCoW2uWU8xqRpp+cRuHVeavFSoQT93+zBWN4Is8No+FxzQOfFPOCkxVJBGXTiBfSv
hCUwPxC6Bhs05TO9QNtxFOEQmUgQKv+AwZSL3ZixZZ+lq1loK834eCr8PoZ3d5hUZr+4qll84r8S
0nkHGzsgaysRx39Pf9bk+0XIg8Lv0FYEb4gcxxqbCwqtD952WbkiA+ZkxduxdxWOAUqx8zyMzf9K
rzMnEXlxb1N9rpDAttzGA1Qv6kbPrp8SWcMn5yJnDBQe4Zv5PLAgyJ0vzCmmgXLiD60kP47DdhmA
iPV+h4YotB8Hb4Dklv1z7+mi4Pw5X+ZCVF3x0HMZexnT9jojKL8flKWPJRFdJFPguJj47SOopH5A
jVgvERJdDPrtb2TBjJnMCSyM6REyXxQMmd6Kc1stiPYiGbOAHijiHnVYrcRJBN2LkUqOMypBM387
VvdD2aflrTkuTX81w1as4r9h1qEJac3HOvt++F0BIQDxEFlWZbm3uoF1gX9d464QG6aQIj3jjgOG
bhE8VdNCoyYeoGGT+B8GTCiV+U9/Tn7vEGi9bPyxP8qLHyVaQQOPZ4LCtk3xXPK5ZtwPTIMoLGPY
3Qrnd6ofkjdiButTjUFdfmJoiA+w8IXvWR94ymvZAcsqembeJ1IZB2t7eQx2AG+LvPA8tW/cPgNa
qf/OLEamfzGNrVXbK5e5+ayrKvwOmGeeVblcVp+091ilWkoQaanEx47FAHOi9mirtSLXHWOZ9HHP
g3D8PQkewgoK+kYd4cJH5iltVjOXMp/b7uaRfqU+7VRrQ5nj5/6NqccR1RT9gLVkqPjn64WuNmPi
fMppbUVAEyZxijtnQgP5FRk/3rpIDM1WzARhbvFPjPFv5aRmQN5cTbh8yLSBYeYIUwur+XmZBF6E
+KhJvokIKvvmd/JODw7UqxU54646I58XrL6zNVIMmt9sXCr6EYjFhUwSqY0Km5oelS2sC0RDm8Hc
qVqQ4FsVQRwNi+Rpm2/6CiFYCjoxBR2qXIx4uhF5JOMQof+uAXxhmy6mEJxgjVUFSIYR7ZNLRQfm
pdVXoBcoV4pjzWkjkb097ogV76cF1vucBP3f2rrRqQw2Lc6PpBFD/xnP/x16inWWkadZYZeIi9g8
7TgFOWaFFU/HcbQ4Km/RmU6SoxxBC8Evlp+TxpQhKZkjYaX+2Nq4palbVEQWmiT0xa5KdVW7HWCG
JFgvVL1oPKHlBrBVy0LXCy14E8bEIgDTd82K/zdyuCx2tg3Iv5tN9SO+DDviKNJiyP3YWn9/EB72
+ZqOuTUcNCnoOCqn8mhFtwq1lJEbEJilODLGM5pqZ9PYMVXsquBD0olm4g29K+A/OunpgzcOvyRK
wwoPhkaLThrFFWZExdefBU6leyLXnc4lJdp5RyV0Cd8PP+OnT7UIYfZIgxs68MgH45pQMjC92UIT
89C54csd0Ct7nHNMBDy2+4asdvHqQ506pF7G51GtG5x9goIwjx1DBJvdMeCCC8uDcyn6rKdaH0yg
t2O35LuWBff167AOEuwKLnlncS5IfJpdNSGdPdvZg7SAv+0+W7TKD3HoZruPOLSUlPEMEd/D9D8I
yTBRZLOVxy/PmQul8YqEBLFu5F4BzN1l+xg5tHVeMrhVXmHo6sBiWPHEfA2bFkO3N47wjcjgjAt4
rTkGi3YQpR3qA14L+rEa1kXwoSlzDaQsCrFA+osz01frLGwhsluL2T6O/NsIMPVwZX8GkqVZLNbD
OPwpKc2cki2WcoB11PNfM1gw0LEANtbwk/SYjLCyJbCMuqQdoEF9iipJy8KJbDUOeV4SXhbZnx2q
11NhnOuARCKFtmLPhBkkcbUYKZnbXndIYdNdPzU2HgTrE+rb1bpj8KQ8vxfdaRehJ7dV3XcaQJ87
Dj7+kIQiSbb4Hi7hhLtD0eMJVZwDbl3HJGUdYR4TjF4WFRcbXubyYe5D/FVyOFYBkUhcMR42rAh9
faUSZDLzxTQES+foJdEl5qank6Jqci+SB7PrNqpomjYKoCj0RwnPKuI5B5TB6CQgvlLnIrawF4h4
uI5GnPwWthJMXuHM37DQ7aBe6sBvCDw+TTvKJE0Sbrnrq2edjfgTRo6b7/9VlTDtExmKDJsuTKrg
wh12shvjU9fHytIWYHqDfiDmQW19Ks4Ty841gSQB+IcJZUEZiOvXaQk1tzE8av1NNgzSA9it8QKW
p9Afen84c27jJmlJIx2E1fO5v2ilD1is4zf0Np59cMyBoVWKw1OZiP1HuD/rjWzV9AUSIROWy50s
QvFWSnWu3XQUY1uBIaAqO5lbF+KcC6X92uq93YiSYzOEX1cbdX1It55ggr1eSvva6FsFdGaJPfYe
0OoFzQtEilO0TPy3O5cDz6xypf4BZ5gbt48IIXqCaRxH/r1/KHJoAVUeHDe1acxGCvXErnHPwrus
SuplY7dC+OQMvh1E5vhGaWz77rJ2lrHmaGfH7ii4FFR4vNOD9SYN9pPOwzxVrDOtlHVgRUG/6w57
qS6DZzpGFjowgHsk4pHF8A+7DhlGgq83f8UpEuO+5efl/pIvxKtaUBgQRNlr1yeWApSJd9hL1L/w
h4vbj7kbf+Q66mxGpK49KcEq+vFUkJEzgupeqRjY/KrT2Ft8zsqP1F9icHQ41t8+gHSwNktLbxlG
t2cKFfbbQJtHJj41WUDBv9RNOD5TehnO+XytnYGGFF3M1ofLhh1lUjuyVQM9Owl/XKa0hUXVq7Us
I0UKV74avCROVToKVTaXIQi1dY4Ox4zr+E6oIycuEVL6PicyQXs/hZyIFauFNPd4J3+EjL6VcAgE
Yv92cqsKAoBOf/gyjjsqEWvGYYvaJRLYkurpYL+Q/BEKIxzc/dKEVFVBuhRj0MtibCjW/drrAOZh
jPc1CtJd289Z12UreVbHBWKH8EWFr0nDYzyKkAFw8LXaj8XHGj4kBzpfEn4drgj+uxkYeDuBhHSh
/ZkZgzg/k4q/pjEkcT2g5Vfw0dFp5y3Tj7dJEsfw2ZonEge6OrcQ9m+WlRZa/XjaVEALC44Pb7U4
2jsbWNdPTjlyM0xnKRClqHymIZ1T2aqfzgZ+MlrO4EOyHww6Q0CTFs1pJ73X5VxJupzXoShe6cXX
JfvsQEaC6fzzflsm0r6WnArxtlZIOFEZgUVAQgZTxc9ivrf9nDF63kkTM81K1Q/zCrhkFt8U1FBe
BWIScMEzzHJ9DNdC0xUY+pzRbz9Oplq7CFQqxR8cZWG7MQbN/UuDRuKAsLcmjnf3UIz9pEq3Rocv
ZpSAcqdUk242QYy/8bs9yuLxNRpGr7jEkyN5xV7//T0JJBe4e1YniMx+nZv/yEj7YcViF5wfukRp
QfJoBYShcR43RS8fc05iGbfwNrUCgDX2KcRHHyZBUZvLChhazq6l7IyESp6tauixe1J2CMEq7weg
XAwmFQhbzwuQj/6r6UTYhKRQDXuL0+dbvv/VBoZrl/Glxf9C070bTzTVmwpku2wIU2r8gw058rHB
bK6nVyb68Sezndi3lmBCOyj3+uyMcO/KdBzPUqcIqYsgOmbTtbuRYTtfXNd66i4AEn522gEIh8It
y2OddpeoU7SSvEVTKdI+fhGKE8+UCcEfFteZJZHFVmDuJAo2O2bEJqFOriA7Bj30+tUWJJK+RvdN
VZe19Eq8GM7K0jLOF76oh2rKXYtMPnKECjD7j0Y1lbWonz8E9Nqnv5LFzXHPPTz+hFLCrLD/Wfeg
jnXQ+lMBv67flNENjNTDWjJsTobK6IGbviM4u+6ikOFyayW/IgQolzmyrRH7uLpDa+mGndspWiWz
s32wdGxEEu26wAVtAvieOrcWvq9G2pkUgBRV0A6YYiniiWsijYgZRYjLz58eMpBLq1/3yJi2vXYP
7qD0LJkiiKskQJQTLtpuak6Teg+RLOzeIzDAesCVUUx0h2nVXUEO585tD3nURlDPdLqW00q4tu4z
5P0fKMQu/WqF/GE+GA8KTW1cP8jDXshCD641cCulQe+ANFh5HTncm5bGwcRUX96P8dQ+a+GvE1zO
z62YbFe8ZXzwihTW4I28+FnIRqUMheV8eqWIDuSK72tohgiMigc9s4Mc3+dB1+kHPYLp7+TxYZgk
J17Lpm+kuIgNMjSoJIy2dqzlbQ1+YH4iHrrWjGqHSixpVUfKfg8bwXtpLgG//keNmogBGnJ5qTZh
NjJtKK99D0dT/LixazbyOwXaizsqeowewMA13mzFwQ7394mwSTaQ+PxmzomUj0z1w/7YjhJ89R13
V8K7Mi7uDgGRN9nAStlVmxhAUMNysWwiSoi9xEWsKgbEsQgG+KOfNjk8S+hlXmECwYwgbpNIgHOM
KtK8KR7KIotZfob58O0alOLy30BajxNuQzKCwAFDEQsMckEXCx6x9lkMIsPotbwYbKF4Cx7eANMG
Xl/WhfiqvLQp2Ywcag0a3m0HYjvUze80Ro/J57iDRI13FPyPnopubm2+4YOW5/b8z/JBQqz/wAx3
cO7itA4kxP5TV1Qj7GRBL8EB9O/sec2SblGmUgX8vZwLYxfIPAiyTvEbYBlj+J62i24zTX0T5DCm
mC2ynw2nmuPf3HHto4tZG0nT9GKyhR3/hmpu6IukCBZ0WTGsqQF0Xbp4h4jE+cbhuTL+MeYiAyGy
VzGzZq2eZHUJDyREgnBigoxzl4SW1D1H5tTcCmcB11wf8nUBlY3Ehwa+y+pPZvzFAMTrkG9koQMB
06mSWCWEeV5bkndb7lduPcX8/axqB81wMCM++uAkcW5BsMxt/P2sQUFosc9m8Lz6aDb1ccZ9x3eS
bZrPaGWUHQrkfd8exhh3jGSJVbAwUhrRBh9RuhtQVuuc2DEbo0iX1Lo0d9HqNaRzoaDgOeOg7ta0
iPx5eDyGJnORtyLvs5gOvu1OJSTuFnA0gZN2h24uOkr6WZlK/OeXrjccvZ1DUpvae4yJdxVqRbjJ
Xl8XRiZtJCqzpfxUHzKtofqyGodM/LxfZnBRheQgXtrf3byKRE2Bx49pyBwt0bjHzq95sYgWyuHC
sMNwcnZoy87hHxD1i2nRxf91QKHeeU4EGLxb3sKYG1JXBP1Axi8MhEbxuxnh1odtJPd/CyQGhNZh
uh7GAOn0CL0q+aTN0YCR0ppUzUtL6P6nPstmLhxqaPNp1qTO0MMnysbqjqLtje4xHYpyWs82VeW5
p5jLbfxJgB8kNSn901KWPOY5N+K8BxsBt7SxnKhSYO/11wU7Z0gG8VAh/hXf1ydpUHbFpreiOGNd
wz8V4c3hSW8uPkZlzKJyTsFh/wpivEKKjwAiMA8DrhFEPCxZ6aX9QcexcyrIqoJLKpjQT5M/sWEt
uUd87x8UFfnqPXrFWVraZm9mN0HHWGDJTgqFiPu7Cl8J+QTA6HanblCwShL2zTzjve2yWbscOn55
0m5BpWDR5EEFFq50DOcEYJ/wb2VGgdkO4aUdnIo/g0ixGsiYoTXRdwaEIcOgzsSnFRxQFphW8Ax1
GAE3aDI47Lu28r9Y0O92QhJh5+X5DRvsFRHpX1E5qvW2GUGSzadHJpYLgHlbA69tNHlmZhTXvW5L
rRE8kb82AukFydYXzPYeCXXW6T4X2zCn9qGXpBefhF0wacP5XvAg2xvniQVL0A1IdVaqq3oIYvMH
hq6a2Zn9AZGIsgj1m+u/K/C46cX8SOh0w8oJOzIwOa890ELo2LyKwqtiztB+SJK7bimWxN0s3sd6
aHG+Si3Of7YiG5j62iSl57+qHpM5kNC3T3Vrol6MzjdScB6jiu0takvY18vpegHi1FbZXMLGGbQq
CLcV7UEK+CymHLfo0d1a+akZNq2J3W9cEUwtvj0OQJqJ3PxRL3hNd820jDV6Qb4EXwI3mGrfSSx/
9y3Oabd48vOWsm6V/IsjZtHQ/3YzDjIsvPEAH52uBuMRvVQMPJksymBIbR1zev3F91MmlRVkuPTl
NWL6QOgnaobD6zSRgeqeIvubmxFw/ypdXswumDTM5ML4bnUzMlkmQNkP2uOo4aDegPgZqQ4oH+dK
2WwBgGvQZtCAvz0ySn1Dj8zyuvs6xQjO0h4StX1ZWTmn5u5CK/bWnzjOmy5RFvbNRR5mSCX40HlZ
+hkvtIwWGl6UTTku7yWgSSiUeuqt4sJtm7DBclW1RFLuPqm0khNpN6wdq9+Me7xMlhp2J0Y7QH2f
ffXDYU4CikT8TFO4oduBm973CbrZzYQrn8A+2xyXKKCwRicnB6Zmbd3ABMnBxyLSkJk6ykeUPvyP
V3d04RnXZD/Kok7ZNpbVWqH6jkREzLLxnFc7P/DJv+UYKT+1pFccfiLAEBeyIftbRIUaG+DV2KrP
5XhbsNcx+uXfm0K38aR2obwUDG4Q4J8UpgE+UnvO8B8T+EOKQKvDBkHSuo3XlJYP7SaHJlKEbJl0
UylzSHvPDNSgPcYwFYTHzRtmcMIOWjcAX0dFzf+vLKwdDnR05JsVIlN63z/qEgD8GdGmk6wUr+eK
+q4pWpGSj+jrEXNzxyej8sWIegmPaxnMHagW09oN42v87n8j3qwrocFcZQg16mwwc5Wx6iMgFPjH
kYHGiH/7AF4AoAzHkhKXfZ6wS5j98xwTNI38rPnK86Xcc+eZKbUw8Ep5HFHqcHQmRwlpBIsl2goX
ks2jIR/F9olP/xajI6Ac3vABrYBpiOwBJ7TpmCNY6kooy/zXaMZLasOQkhYgC4S9WIvY4kFhkfqs
FzyASPqsGV/sth+3tdk+vDiA1AShnSWRd91fe3Tq9y0zKwf3QP7JGevbXpQIUgvzSsugoMdeiGba
jCxr985izVsZJddmAyxPxjAgpTvooOK2JErYC8+TzF6l4Eudh24hyLSCfVS7MGqBNk5iiURHzeSt
fuunezrfTd77wrE0IeFJIdJczSbH6HaNiMFih6nOXLgOIBJ9xLX9JYCtgZWDKRu2jClnc0toDMz3
dkFIFiSIKie763J7dRAzQJsvoFHn1HdQCo4oWg5TNvp9Jz2vXSq9FFFGTYnIudeQ2NXnG/116mlW
kmbMdKj2e77tDOpVDQOTHQcu0Nv2r6SFKwZNGKltHunnolZq3Io9hR8NRmRdoWL9YKYkbR6Fbj2D
6+nkVlasOV9Nde0HngXw9h0lZvKsKIwCO9ynmSxnq/RRF9NDy0BJzEXtcjxgmUqbY5zdrLL4bbxX
X3xqMojlH6MGXNw85yDgKznWqP3MAFyblEF4HNF4az8vz3b33rAKCRIyCCBIenVJ6e3BZUDt0X63
8tuPz7le5BBnFt8+LUq5TLa7bywi+lAVWRnUOjPGRTC8zKvZfz2z+z/d+4NKcOa7O09kKlatQCJv
BCxH8p7mJoRZomf4Wz2OuxW8hqKuifjaZcZfPXlLNGlUCXw9g4t50BI2n1f24xdA19geFRTi1jf/
lkuJiHt7UZ0rX2g8MgPkIytxJ7SsZIC5mikmVYK+3sMo4Vzu9THUeW/Efj39oFQGoKQgq1DgGrCw
IPTNMwjoN4qOncSrbsxuqD7x29QgjWYP+xNErIR/XxjUwd9vRAeKtnVSmY0socwshVqNs8PpWcCS
HvHspns1YJdDgo6A8/E+9ZsuiilvSrYvdSDlrvKHSKmEEhC1/cpyiU1QgmheekpMEEAG1D96aD2l
TWq/Bf8jDjck99j+CBKbr4S5JU/Q3g7FuvdfQUpP/a6envGLSS0Y9JhkV1qX5qsiiEcMYLN+zZSO
Wl2ONlttBfkMamogHvCl54SrhB0aoXtdPNetTQWXv++TVP873MUSXCjDKykBg4GakIeUwzU8njap
wQsyktN+S2r5cOa59fuQ0iSJaVhxXCqsgxMMVYXDq2P1C0Qv0UU++Qzd53nhm+z/ZVixIyW3JZAd
fWgMByIoIG0ZYNFf5mb7nfpQtqxv3CLe28GpGNnKLjQXEmG+3sltdoUAAacWJMSlHavHnPRyVc7U
e4opnnxzkp4EnhYiVS0bMAfuFj+qF3c4lMQOadjACM0Yts/4QMeQonX+XEqYxVHrVs2eIRLroCdP
dYOFdVtm9eG5TQEs1458cIUa5RylNvQqvWZ/IxQRLYXiq0kEbtci/ZpguqUUTKSLmNJdWeSssoim
/AzXvg1Q/xldx7x/aXQOV8aVAKck+OJYeFzyc/Zg7MKgv3a5e9sR+NMhLcY9TbOtFbMI+HKIcBQo
H+h8eQU31PI48UwNJP0PkMqi7/tRR4nRbAXfgQSvY9751bNMfKV1OmbV0IiDVLjucn0oH6exuh0i
Q6x76K+0PYI2RQxN3EZfpggJ1PiqyFPuFnas8fW0piep0tSbFSHXBIrQha9/nhUDxchweJs5w4Dq
XSb+4Z0qAwGSV1Kw6A0G8PW0YEN9lvaYT/aNBBWdKJi63N5brQQSLT6T1jwIa0Kku118W5N310Pf
dfnu/J7MteILud4HdGYb3soY14bI3+XI4TFek8fpVjTS8Ma+hnPq9JiOj3EDK1X2Sn7XqV7+hUj7
7UVs4WSeiBKNha+Kn7PpC4nSuWRM3uH8Fza+YzWdXlhir3T46+S4dXhalwk4sTjxsMCU+DFZZ3iA
O4VF2nF/1qO9x8smK+11FryMFn7cDPYE5p+pErlDi+0JGcFkJ0TXgMK5wYnf6jmrqoYDDh4kQFlx
lBdw2JPAlcXcz1UFMmaVb3PliujNktOF1AJHf+lVafbdfVVONamq7ucmvV1SxxyFoNcN77tl1rzD
qsZKMxgOeAo+DOUiCPX+mROcDrw71274z5feNLNAt7j8MtV2yLny8IYmwZ/oHLt0ZQAIFtLW5Smt
6YOzKla12LdudzQDN38kta+g2kqxijfVENvKp93iRxlSmWHk0qavwCbMDJgm2gf+VRepBwMOVFWe
BI1BTY1DnV/15tYrr8c0iHY04BdR0owgfbnG19MMTwCHbjCGtL0yu6ezXlxiR2CRUjaEcVr0xO2O
k7tPdAtuQDYGz7imFaQTtUFMMQzZu721cVD86GgERX4c8HSOULAYEUGEBqrF1aESPXlFm7uBD60F
Xt9uuu7Wk9dYB38nmg8LNYdiIGGTc0NVyrd542/Ua/+rbhVWKzWz6hEjYvZsnaYv96oUmesgPHAg
wugV5OyEMxHB8Kz9JLiStitvd35faG5h/14R8mZZVTz2My+wsbqA67Z+qRkhRt5DJUnfriDaKdhu
mBmdsEbok3Iu+lAauggMo0gg2eUtaI5lWii06GuDUvvWg4XXZVjP6nAH+4rNb5ia8PrDqAhkQ9KI
0j9WA6sUpbI2B5YMNL3dyn7XX/SFtIKiQSuiysOPA8o92gLIWtk1wxzueeJTQ8Lo8ilRgHAGZ8uf
pqoyMCK4W94x4lzg4dUK0m0kXUwhwR1EsZ+AMi08zMyILNNlwnSX0UmQ8AFxOSVn446PJYJZaJH8
CoRvSrwyTFJvql5aRtZXFY8kg9947r5jqrQcc14vmlN1oVtVZErPi7TXJvBkzLHG5heBj3ntJXIT
x4OwZYYqggGTuBb0WJov4tydVwfnAyissUwHXWeb1dPCNdkgw4O++eJ75kY9PJ0bMgvo+U0u6koj
gM5o672zozPt8bT8od7d6nDrFt/OMDW+gye5CPdcNRdgIiT5z8Kpfp46+Gl/Vp1eg/ty7u/SuZgc
o+/ltgSvU2fRalu/PrF0ynfhHNgE66Pus0+kppDUlepL9+iKTIT684XqoiWzvzEnQihtpJLfkuwS
HWcQjEqCb0O4RacOw3gpxa383/SdciDAbTWVtug6z3qf4IWNl1UvByE4oR0+VPMeGII/VHus+6wl
JNbvfYAlfFaz5xsUf7gQ1mms3r2qIYOq9poj+O9rVCLkap/EIWw1YFwr52loFLnug1exxOawCpVG
qBAGFZAju9zarjjd3Ab1ZHrbf6JgM/HqRjduoA9n+GWdSlarFW3dxrCkshVRc3y+kQ7sQVbtCkzo
bTCNZ9IIdvQ2HHAiRGAu8n5rs8LLp4BXRe3RZu+TMQrwLIaNlC0whNBVCxzf+vyH7RWy6fHgtL+O
yEVeqzs1v333yHa0TDidjbGNKVYuGoyjxP1j8qgyWH4WasMfGXUpPunqU6GqDjSTPjpayYeXM5T1
5TxcJhaZFoOgWZVmMjVrBf2Go7ZNx4l5u5Y7vtVYk2BmLUaqxBzJ+VCyZMW/NbXXZBDjORneriK0
zkrg/PvqhG22sIOTiDosPVbmUC2VdOAosfp+PxQpfapf9Q1uTNOrKKyX80RyzOXxGQkp5gjHNLPX
+stfhdvMZDQ0J6iUOQJg5rJ3Pf9TgpyxIdFwgyI1g0hUQnTucbJugKrajvCN5F9FQMhO+TWkOdaN
c4V1/cDN6zwvMHNdLsb154q+SOmcQkDXmWh38b3xB3SwaEztdUdb6p5KKSQRvSLPLQ59yvDvtr/e
jDoYdfeH7kbGsJbePBn0Htarr/p+XgGAzOzVzFZJw+hDUc/1rPgqfO0p3veXoAFjtru3pmzSeKyn
wQYUOaCpA0Ufu5SWScQ4nJcTrI2MuOgMF6As43mQbaOlv4wvrNi17FHgbv1qL4ue/QSwLHdlO6Py
igxSa78drFT6QoQpkR77dnuVVmBA0rHtzcpaKc6e3TQxVYi0P++blm1MVgCizSTeMk9PKAkkqz0q
6zaZ0XOlRYg9FphJARaDyyVNavwISKpwTcN7XxaFbaMLeFFlTJDFuTdcG5JmDub1C+9E4WXt4xs5
NCYUL0Q3tGE2ytNgr1NH8/WIWNMOIonzfzm84inmQyqywoi0fG56eKJNczCNbNeVNfkR0GOB/Ud6
HFOFP29Tfs5vB/Fp60+K9Nxi764niDsrilU+Xk3ZgMNHdav1chL30Xwjn3FRcLHP+xpsH9D5ifd7
wia906jJN4f7aF9IVshmh6KXYpBZHWEmMkD0vg7kVhFSjQ7kwp1BVjA5erjv4ScHuOJArhQesDPr
k0SRs6Bc8tzdTZ1zRyCybfG9pCK5o2dXQ/8dT84i/0ppdv27g01hIPZE/fq9GKmHh/8JkcSqI4uf
w1TsY1yRo7jZ6dDCZYVjAHeBl0Q4OgLvaa4HjZn4u6/77NO4O2m117IoQ+dFsBltAXNu7yhZvBzI
0ZtIVcoVaT0DYCq9KPfyVHNLj8imk/N48fqZsDUGLTSwthOXhR8/uXDYWJQIS/ddxjLygpOZE5x+
McdT2C0iIq7TXe3fYRuKYglBw5HzqcNOSHLSSY4t+YNoB3w8M10JlIxQLt2Tk3OKKQudI4/CmLL8
+MzXRDU75RBBHnGhh0bAreMP+t8BZYGy1W63Qes1MYqH8r/pQ2N29TCrK7EOekfJgXrk3ZFGmsPb
ynC08WjLI7sRpzanmEON7pDvekunluBtHMgfoVCcPaXQ++67sNbzJIhjAuwqj+Zng99ZfoLWV0ED
VU46kPkggdLQ4KloMKHaguTQTXq0pnAnz6Cb7f8y/1Cu5wMoQQnFlhVKaJZDmY9TbA4MQRjXMvyf
PpqJMXgX+ZircrX4DbUREZZWDqI9eWNVHlh4OJIyY8whU8si2OpDGqeW1YvjWXulA00K7lxIpEW8
gfpqWLDtUltIf6W57QQdF6S49yafp8jFRHPoq+58U6n2kcx39WYmIyXIomBR1JUfxlLNH0IfyYjb
YBVHJKGKSdOcLwXdwoZFg8rc9+ysv0F/MIGtXb79g2bMD3NE4ratFRFRBdvkULYKzgd9HLxZDSPd
l6NMeUmJZ/jRAEalKD9psEdEwMrcD8Mi9+rBNH4ZP8ii58bNeouNxqJ/bSYwFo5i/9dfX0AiThL4
8rl8WwG7/VRjZd1aN/LU66NH2NNn2Xqij0lCZ4gBugC0M2lxrA5Ayv4NSCSGpo64M+lNeBlHomkv
8J7oiwaqBHXA2pTx1cXf54qMstDrxhJRRgGepsjkV16gThpc0GctkBN9mOrV0OlCLRg7PXrPXjvw
KDeMp007LQiTg4tG3rCx11FBJr4ZOIciALa7iirIcNudxC5EGCWQ9xwyJ916tgud7sxNTsqRYtQM
BhQI/eMlq5o+9DPXhqtEkBet3BinVyAWDUyY/DkQxj3iz9DHq9dK3Tmpv64MVKOukHXonKgw7uGb
3UQN5jm2kPc324wq6KfVKqdYcEwViyiJO9jiQ6eBY3mMSZRBxOBPOlH2N3LvHTIlcIseCX+VlkO4
9w+LVsfvOCLApm+WXqiy4PeZZLLaot0/dfYH+i6SBE/nIBETZEV0bQZF6u+yMjo94Hj8wzztRmup
KDa1a11zHUt0qnVyCoPtns4ZXMqxsiDjJeledJuyEjvZWPcSfm+DYnnfTeb1BcXgNvZyAZw5DDL2
kt2dzsAqhWSsVh1j826B6jNGjGbwpuHnHDiEqp5ZUK1cNrSQ6hyBEQBzxSckSPPN+hqG+JEeiOk4
sQTWETd68SAiEA14X65Qf9zWekvjs6Hi0sITtCfDky0TRozLbrp5lGDYK068XlQmhHIshO9m+WuX
3fAZxwSyXvGqYVJhDxe0A8li2M/6alACErxGZcWsUiHK5OUN6q6Uu1IGXRGkliJg84XOOUwVuiXM
VY8tVGOcG/JzJkzjHGFakJOdu8L4G3jI0Yw1ffmWdN4MjmJLz7B2VxLmfGOWCRcb0TQOMDg25qvG
JX1WQ5ua9uEZ4wrpJEJwSV9fiJ204wWuDyMeGIfp+ytsK4rB8ZhC9Wxb+5m2SMo5tEwabHUc2b+q
QHw+ZMCoMsryRU3lXa0QYNIEnZRVOu3eOCzOxlmiBHsKv46ImeK+XueRgZzYwYfVLRrf+ZGZ0Q2I
3O8CQmCW9Dhlm9aZuQHu6ednu/EBIblZK8JRkAEUn85GtZ7hzbHeTtPKPR6aXxJDUGCdTqMthcxH
WiVo0+k/c9+r6tptlT/gb0yeuTZ8LJ/TkVRPiQ03JYBxAWTrRhERJ3WYKPp1jI9SuYjEx/zeTyft
8Izij2Wc/v6dtGsJQfWdhJ7RmJFVN8VqHwFi1cRAPK72HE0lMg2n3XhTPz/wdRI09No7EsxUt1xO
iigFNYSb8Nr5f8f6WuGEP61j7gJ1wgdS3lZIWaR7nIUXdgIntmJ7sOmZkdg/F2IJtfikrngT1+yg
FLmR5nRsCZ3Kyocs+f+uXK5eaWiScHnyJg6N6puOx6gZvHjVsZFBgPU4fossnchgvn6RLfQ/o97Z
3Fcf6IZAJvYRpDykzC2lKB+//Sy7anPXhCvD+YEEysn+3tlZAdzrewpHZ/x3FEaHVx0bTVL29FIN
EKQgvkWAyLcu/eT0vtJsVijTc/3use+bgNXBRGWmK0lb9GteO/Sm91vSqJ5jSe61jy2I6IMbW5eG
GdMibTeyJyPDS8LxqbRi7wHkr5tTlZwYhNyjKWI1qxM2vMzRmsyfn88jJYEibymm8MoMNoNXDYzq
bpw0CaPowmkHPKWDry053hRxSiKdK93py5J7D2ScxqtoVyuB7bcY8k4Z7Ee3EETpL3RAOTYELt3u
E+58Y30Y61mhS8NuonYOITRNfiBlujtchFb6gxtgkcNBgyH52qcQ7CqtC7vYBDiovtjkWgO7U4sQ
JmWerdr5R5kBuXyVbmFx2QeKfGh/VW2sd970e+uOgG8y0LWwGdazKmcukCeQ76MeDeaxt+ek86hY
qMym8Sy2ffXKMShMnMEpkfhj/PnxHKMcP4Y3yTuT+z+SZMVzBCTfWYjGn5PCwYJ/Ds5NFPl34wxm
EacxwwG/QqR5ejPfOMqpQ64q+RFg/x5ceCz8XyigD1bH6eEJsxCWO7BuaimkiWAKHn8lnI5yuiQM
hsv1a2UrT115G2LOlhP2EK008LnZd1TC6kja9B5rlu/MSMCTIbzj2UYWggnwtU3Z1CDQfHsZxOMb
GWUOteCFTJ8bRX/46DUC4heAtWnruFxG9w5/wBV61kkegZm0YKzHPWJIi0bE08NxMvibPXanloj2
Ue4hUZpP/FVWfMtVjpbpid4zg5sEwjZwi2LIKWhfKA3l9+FECAIQ5/h7eDZ2S0krkJ9qswcvu4/b
iocv/sIVOWjeQ0FNMHe/gh4q8pQCqp7PK8frmu+rX9QnB9g5Se78g8FGyNednnWbYrG0EnrzVPjh
GUl7LpcJtoUb1PFYO+QZ/IBRWxmy3P0RbwqIxK4lEm8bgm46xV9yxfK9UUAMReDvusEcxGcz5kRa
WNs2zw7siYAaKNyKEdSaKDfRU2Yt4NFBqqvAx/+8/nMHnTDK6IG+NDspi0LNQ6a+XFciN/GnkzC8
8E1we4fNGeU2tB3FvmpPGvOnNOOChUrTYYhDDLqBMkORNb4cuoeCSPgP+4udQwV9Ti1o1ngWiqcD
35oOemb8XUjKOTL7j2G+avOGTRjzadVH0hBkpNf+OCGL9eE+P9RixXf5ygkKbKGS5dn/46CBTLpT
W/wdbfHKUP3bhVcu8sqnI7Gf6M8Fjex4FIMzxLlJ67Yc5+8Ti7L0uP6XbsI2/msI84H+HLVTNOQj
GEdtigSy+h+k2yncinjoKnFoZ++lL1EG+GfRBXgnxKMlhLFLxDj4/eetmvGF49+jMwKwejcCgxKk
/Vz2mAV3aW8/CqlDKqhK1IlB3t123tLttFpgy3a+3JKpLypSo5LtOEBl+zmGqLwMPY89huuDcSbE
3zLd4J35//4r+uYPDB0ZO3lhB22/0Ksdf3bpgGMQVR0ELaT/+wGxhsPCq5PkAGhxcnYL+AueZEUa
/CQz01aQ+A6lAOW1+lsNNOAaf6zmu9PaUwld7MlSsFWt4qxa73N1tW8sS95FHStputCs4tiG0iTI
Xdaa5Zprm94c7nukMAgzUNqWEAqdeb25KQEwR3rDPkzCudeeFgGNbqVmgn3BsS0qSoHmEVE04Ve1
6T1xk471tDAxygwJH6gN4CjCY9OD/uFBrtvU/T58ZMgk2Ew36kOPAKhQZqPiu0V/oKJlEsHDJkvj
PxUo5FZAUiZpm9lPqIyuvht5q5ec4a0aFBEb9s4Yj48VBbwKB935+GrbYIOKHj9dxItKlPhHla9U
B3XYbpWxiKBL9wa4PmlMN/91a3oSxboPiW5VLTkoHSb2Xkg9FXpI5cFI4/knOfMhBiN9wTrEW8a0
dBSvATLNNZzvtLZSeShz4i/QBIrRWOLOKYSwfk0x3EfeFq5XQnI/wfBU/dDYFbINv57yqW9Vd41a
NfmPnMfLfRDgDSq2/cBEAT5ZjAsnaJpa5ihTLAJ8wz0hLnmHmN6AY01Jv7gPkbX0gL+WrLLTSnvH
az6gK1GEHZiYah9RT2pwLQWWRanY7e3kK+qFwXQDYlvz4JYpLX9na/5NPiSQ79PnTHjPte6d2B7M
9yHKVpDf0Y6EjZr6uHMvLIEDXV8Pxvz3rlUJVtzuDbAAD0RmmZt0MU5aa6rtJQpku6kk0Nhk+0PU
hr1VeZW2hoAXVLER91io1rkKsq82WzuEIt9tr9Iyd7MCEcnxQ4DDneQJrCfYHYBVGgpzmmIQ1xMI
LvkOCW0Qiqiwkmypqc2scX6LXfL4k2nxlSdplws7P9eeFn9FPh27nWfN6UN8/QHf8n6vhWojNeeg
tPLvWDSsmtr1CLPPBswG1D7WgNpZIZboz92aKdkYEbewe70qbxz5dkkEwUY0LPKrelCaEfzFzFL/
MI2YZwVGb5+oH/D0bA6s/q38nXOpBQfOq4Gx4egwg9U+Z8Pnh8L68yk0uKv+RjdGnHjebRyPCc2S
YVHeIrAJUf1ogZ3Mv3lgML7ehlWZ4omgZxncToRDEnIP4asm3ozDQ3bWaVeeRF+Hd0XXu8/jl55W
m1LQUK3fxpMCMSabPZ7j4eoFz9xA08vx/ttz82jWd08Zi3RO12sqB3hY1vcQDvI0oe632WrYljQI
NZdW4zU9h6j2CHxzCaxdaTKoksuIBq0kw2lj7xI1/OK3FRWPgScuMoUwDSDsNAV4ZnY8Dt2fCYhU
tcnrH9OxilL+Eewa4E+oZhuKHN0MDS+ibArjoK7SmSj0y/sysrJuH1sp2mg32kKpZpfZgEq6GQZb
aXT4AEN1mAmMJjcBUczVd6MLqiq6f6uAGoFuwMu9CHQ5FeiCFEDVPGCKTXtBgyN6l56LqtzYaOVx
fR2UTSuyt7evXcLVkbUBVNUhNmdCdm1YBQ/JetQtzxnaTbFVYiDjaQFIMtu25CpjE274D/sMN/Yw
9y28yROz4kGd5fFrZKJe5WPbrxTQF+l1Yy64kpJ3MO9t6YqE0kSjlp1yK/P18KeIf5TkgHrnzQ3M
LPGsONsyO6OLwaEfn7GtUnfD5Wb1ewQ9FwB4GKcPKBDh3yaBf1MkJwMpsSypClzj9HVvbn1JmgJ/
qTEXG0PkgYtx2+8vGF7lBxcK1G6ZJEOlXSkPXarpECCn+KBUxhTy1kTY4iHksVoqMed1Fi8KxJdq
aYJGQ/F/qnaQdsZspqvRFdY1MRF6lQGaMSFo7fRJxKpRh+uR/zbrlo5YcwGmXivyq9bU8Tt3A5lm
Zdq/NX4aNStpVORCoM+94LBnM2+MawkTCLzmD0ivGV1FaC9SrNLdH/N39UotulB4xd/WnjKpG25o
tCgwPP+avSnXWhbb3Bf3CfqdmvEuMpV6jTu1ts/KP2CMWpdX15sdPSw++Tj2nn+r7wJPA1NiL++C
DCqNvcNWA4I7x0ewo27WWn4b9iIdekz4EuZk3OgMnEpnp1mz2tcpF3y8R7r92Hiby1mP5L049ngC
7DVWYFY+LIIirRbGGmzsy1XBp1IbFa9xGNTKLHjt7lusizRwy4S3GUtqETufVfewKPdJiITbMiRf
NHZOqHb9QEHXXtRPAWszCWcwb21NyF785chSoHM0WOFDpmU1x8at4yM6IDVerDeocIoVJ39NwJDa
EAIkDfRvXzfuCawMaLtdyoHWy2xYM0T5BtQPJ9FBp4wK5C+fllyO5nrgRtw0rTkevFtjNSVvSqWE
fzLN9XFn8ySwQkwP0ZnRCsXVQPZ1872Lo50RPQNovhJWDnGzCSyQIXFXa5aassQir+uf/RRLwMZ0
syI7HsZNeetgRbkMiKhSEIK4qWkSP+vCubC7EzDpMc+wb55X4WEOLIyj9iCXYhceUxR87Y8yuOp0
CM8W1+SgJruqVmVzyEQOzRImVnKZ7UQHDJyrcYXN96HZ7lKHoYkSrG6QUWjc43zOyXH+u1YCEROG
E0/00GrA2Yj8iQg0fDV2CFQKLuGoIb6ra54JFxm0OdYxUpJXhWHCpOm+bZBe2yItAbS7uQuVyRTn
aZTUxw59AI4QaM4c3gQKJUj3x/JPAiLuNLQXo4WP3m1YXyr9cTZH6l/J+oszcpNyUbyvsMoiWcy4
cTMykIT4l5TumgOKpArve8cmuh8vLC90prb9Z8UV86RmbCU+nwPYUa97tmyFCQTyYC3Y30ZgO/Dc
GA6YMESaUobglRaK8XkjYjKsgO7aqzqleavfyxs/Bm98vyaMo6tS2dESQnN3yVicmJf6s1mfhl3t
VVMifHkvo66/U4ATnpoox+dwxUcPKiVl8esT3QNKKVLr1vN1DWxiRKsrPgxVlISMEQ4y7407qOWl
MedCwFCW0EOMuORvjg9v0ab3RwbHs/Mru1m/T89FiA5S5lyf8POUFECdWuRm8996iO0jV/ivh0Yb
ZiwxtufXwt2Ld8Pr8lyt0M/9gfRlwu9BrG/fQCFh/IE+pvdX/hIaqbL0mQCplaC4kkwi23ihokj5
XqJVgCBi1tv5aC98WRHmpgnoYomh1S7UdAhv8Gf3SdhfnUhE5d3UAAjn3WGCzB3pGAbKwECtsKzO
rq+2shFZruM5UcdYcBTTjzwcGd0wM4mduwS5AUxGuAsZIPLwUfwHsxO1qVxrq5qzDmurR9CXcLrw
pDROJKGzMG7lJGKeFn7vL9ctudcvBijeGpY3tOcI6hTItS+mUsQp1wCbnULHI+pe3hJA1DHqvwlu
Z4UYr0+YBDA9OUJJeF3lOJUjbaH3bzVrmGO08JZcu6xeHFga0B7DPpBm4FidMEaXjmyrjqmv3VwM
PBsLT6MCgFtHN27erIsxHxP3ln4aKTNoFZDCMuUrgzkSgrlNl3p8yawEZ7f7n99vDAAarw07qOWy
5+KPSwxRNs5a1BzDrO7qtVMGRED+QUinQoKe01cQxwQlJgo7NWjd4PSC1xFlMe8VIFH26MbH14G/
lhLbtclkWDaalipVUuw/oBTNWjOvSl/v14edjF18GNEveaXNMl9vnwtLJ4+H1aowgIVb3e/leosk
t7wTICtVHi7uMBwdOxT7GYHdH+ufXIicRvBJhlj9YyCyRSH5TA5DsqSEojcIcH5RcygwTG24MsMo
aA0uuoL5WocmBwiHNyAcw2rJ/BKJ9mAC48806uHlfmi3U9N1SblvdSsuz5wRodqN0kIq+yIgId9F
1LBGyQ7P1VCvRf0QDCnc6Dff7uqeOOFIWFx9AeQ7ocvmhfxAz3usB7Njc8F9KsuRPisGs/3IRQhy
HrRMycfPm33lfTTUFCZpxqQYzf/nLcrC/xkkCwpe4/dj5PCJdPEZkIJ0IpDHjMhn3ZdoSvwrmkVj
ymh5aPAZXjFxgNWo+E5skTmuAZ8MHuvywjeIoHjCZ1CloyzRhRYrdtjcqY8ppifyxlmq1S6b1FDP
NuRCyXpSVbBcnEUPwlYvzCDu/0t8wVg/x2e0Es/r/7xXGWGROSTR2GoohNwm/r9DYdbUuxBhReuO
pRcDs26aLKnenn2Pd0GBcSu5LWMAYrJMbz3fqW0b9f7B41y+KtpeLaAv/i2WTliTB74w+ASaniWR
eXUnpe5IL0BFrV3nA0iFeIjnYOdKAcvpaHzS2LdoawxOibNNGRh+OHdncAHk4FY882GdLyJeMoJ5
MOjeZGfVRaQXkhKSc4/s68MC+0ZZD/qpWkKhd2rMuwk6SZ8rQGN/NsWv34wSE0jMR0d6nR4HI8/q
ZJMzVsvSVK2cWC3wrZqGETXvcBtr4QQ2kNx+edLE5xtl2fu5eKVZ9b2KYEsPb6JxTXgiJg9oviXH
x82vjQqenbq0r1p6RBqdJQ/OPCsuRB9sTeKCsvXuNPlmwqR1TI66mPgRh4tl60frINfcMfbnco2A
DJXWQRCBuFx4ZxN40bDLVbpAH9qHRaJAeQxPVM1IPX/H4FlONc7hxRcINWfAB0WJrKjei99Sh9Q9
QyO+OLxTfA6lXmk6LTyZLdYfiGDyFdwgtnznhccJqbBzAWfEAe34VAj6jyGJHAHFwL5yGzWamnnm
0uJ18mjn24yAZTk0ht3Iv9xWtXRtkiuzmPVyJtNTidVv7VrACUMwEZyp6QTJU47RSULz2fq7LA0/
NOKKYCjOfbtERSdVSMj/HjPAKX2wafjlipC+XHQuRHSwRZflBXVVtY4SlsHWvktlcb0G6V6FqQK5
ACW/lI3zq5af7WzBT8rj3i1qgebN8dOZE9pVWZMOMZfOq4S+DxGb4y7pOXrKqIygTrVWKlnZzekW
h3TvCDJOmWS2AE1B6J1mzUFvV26FBXU9M9MxgTS2VQbZ88U6Xcdh7Q9hEf3DrsL2gSJIiUmA1kTw
e2B3vduA3pTqoSPl94Orw4J4VKgxup5lzi9EQODQb6Dw3/fP7ZpgvGeUeqWlpwOuVMmUaufa07Cn
DBKBIo8Ly2jitcssXc0NtoZyCVCzIEtAKWyEWH1DM5g5lXJQZqJTjr8brELhHqEMJNbhj247aWcp
o7Eo0xqGaTbI84NaVTjdaEp9sXnk6qYqG2UrM1VNOEFMmyhzOj7k0I+b8XqghMZ3b66kDFCD8U3x
dGMEW2UjA7GpRJ15RmHv+5KaHU29fQzZutETvX6j0Uq42tFNhqeBQeebIB6fhvblIqpO16D4mCiO
ACU2qPJZv6LKy1MqJKqARYXRZrtxEQGJRtM3ewhJJF83Hah3djBIfq4VmhSRakDIT8mG2apIliSs
+cm903uk27LAG+Kqd7GNBy1D7Uy+KZxFTjEQwnkGQhZbWKwLbqWYfTPYgcbRqxeafZX28sRNt12o
Qxc1VCbvrar4I+fLmj9SnQrn2XFtt5m6wc8ngKrT72xiDt9hF1O8kp7npildcCZDYFYbm8eoeOir
Yu6lz4BBlJH5vdyT5/HZE29iSqRRGEZ6uCJiVJhqUbxIZuU2DeHQDElghtEJ3Ww0aWvnG0PkkBEC
vxpPeov/qUrRaEFrFBXrW9X3jW/HPN07KRvBJkFLqWGC3Hs8XOLOA1+M+Mgv8pn9kn3y6Efd5JZD
4ITmR6fhBxXtnOHBiPjGMngo9aPUeg8tH7K8YwNMjEj0OIYGH14MtJz1Dg38FEdxHCt4L4qMW7zG
3hWOcM5RT65j3AGjEBaKG1jdDSVocHTVov/UVRLyBei8Ht2W7MYGKVTRsccYjGyNsqYoyDIenLG7
xybKh9s8SFUYCA0twYntAnPYrVwyI1V6atG9wjFABjwjFGaLqwIcOZYwnu+c1zlzbf2EFbBC525z
YtMSv+c0lOjssAho+Zb7SvM0/E2Pu0TafVPOo6uhUgkM+1apGC7fMhyPxCd/cA8qdFLuQcS8n0AC
djSWqPk1AXTNZVa6WPb/azixZQsSjfZAecllTr6REEhLwziUya3KZeQX8oLof4CSmdJLjm37Dncs
mJaU8htEHDXsgGlXEP62G2D5yIoUA61wMQuLl0i2Ugxk90j7yJH3g+fU1vJqgmbEjz+nodtmbmb7
DEJp0t8TxFFRq6LlCD/ImffI0R87XDa5h4Uy0YdCukoeSaeOtp8W5VdJ0ZQh6TBpii/eBrEyhKFH
8tyhqIohLnvXo38RupdgmRQDQBCjAnXZbEe5hZmLMeDBO4dfTSsT5g1ln2ese6+BJ+ZZn0uMZV1W
9RB0Qqdz41Z1TfKZ15RMmXst/zErCdMbJfHy5A+cOiMhbTthP+Yyap+BqJfoS9OJEZlQlITLIjUI
K+QjBBNrTqLlRddZ0QfghVsau+bWydlQvcD6lawz8Ebv1qPX9Zc4h9u3vuPU/Kq0zj1i7JX2ZHAZ
iXmD5rwqAO67hM/4T0Q6lWUYP1OjLz26SSde51R4lv/0FZM0+Xc45EJzpAYd9G9/YU6YtXuCimVY
AKXAWxQ1cI/w2czlHpPB6t6QhL1pROk0g0Spw7/bR9ZOxtnlF1ChPiOPA+y2LnKvVojHTrhvN8g0
Y9M+3CfceHbzBVmVCpI3CGKgGQHdjsQoPiducDkcEV6aF/2VT4XNYosqSflbdz3NMAbDmvbNkqL8
b3qzPkJF3AbNNZ84YgiCMh3Qhsp99jmt46SNFKrJDP1cd/k+gspMR7HAcdvI+vV5sNaIE00kOpqM
0WgOacoYNi/G1DXGRxZy/nYOSXcyoDPupRALP2JQsQekLh4Bfbg+gMdxw6X/XyPdlnpZs13Spoqh
+jYBvaHxvjyyFDv+OstVh48x4cKksN0jOLIw9jr3jjXP3lMSwhm6cbTO38ByWSfBp+5BXdrtDcCt
VrNeSnCBaRJP8IrVjdFMY1bMDCHfg/9Do+ICYv5+SyIyO02tzEiJLVm/9SqgbChDddGVk00WjYjh
Zcdxy4pbX8fMrMf9stK3X8dRkMdPo5hLmJEkKla/tMKn8kiddbyaY3Ql/nilqMJYAnXp2gBmyuxB
j66EF3KHYzEBikZKqeAu10c9WWKl/Z2yOxhmgxn0PVgq8kvuZ2gj9ESrHWwPKf+/hTeVss65b6zV
28IKH9CidKUJ+NA0pCjkm0s+7Rd/trEl5bxdVSaqNAP6T57fCrwUsDshH7+7kcE5A8r12GR/NdM1
UerbMue9AYTfHaIJP+W3+B6NwIVMeRRaKR5Zi6//hDEOg+V0wdmA1jIfKzHj5HTUqKlJSEkkGvD3
rM717sjBaBdW12Ow9cUtoRMuF3WwGb14DQ7x6kea45rMQXsVAZoXYJWlSZ8l6fRq1qcE1cWBqvcv
Ol6ahLFfHG0kw4reSBOu6bEGZwpZESDl+9nlxu7CNyclyqUpF3WyURYBhl7VSc6sWQVMJrBjSvtl
Nuf/cyW9Ujp/eHFZPSSOMYizsE89bG0fDx+a0a4+guQMi2AT88t86AVgMI8GnQ4WG+180b82uJnL
DQbiCaJqWb9+7xH4vDl2bj2kuJhympAhnj2pbcljqHFyiqIyzSmoDAQ3itkuhr2pzhU85Haq1GM3
cNZes+w6zBW9GzAiDTjMb3nrjMWTX68BFgxjIVf5IgJVOlRDGbuRnrQ6hvrnE3TIK03wzU1qoITw
FEySjUXxpcFULXuS1n/XwvGGc5g9RAzh1te6qTlQWOaBzq8KKSmdkrbmFCfyZs6BTJDqPeCPUA8Z
G1PYvEfwZA2mdQoDokZDAQ4hmcHruWWv7uYytVDIH8xp/P8Scyb5dpk4RxsbPtPaZDn5GpWt7a+y
YcOkrGBdutQGrkce2lkS/mHrQ9qSlojYgLugDY6ak1ft2TXCRd6OXP6/N1Zxjwy2ncBecwkuBAoy
ny0tzpKMKNsj2QA9L641XdfWs86c+MDifpESfFhVJ2Hqk+sZHwQsRVTc43wtKEpUl5BmbddzO7ar
J4wZn/WoQ40+VMIKHeP2IL9DPBCuEmT96x3WPf4uDuaxx/7C0VqodFRNLmvJvkf20+KQEhYxYTbP
62UKwJ9tT//fYNJQ7Hj3H3QnYKSewGhooO1FGFlBvc5g90xMwGhU2oS/hJBYMxdNc1N3nf9kgaPF
3w0jDdCI8bxN/ilZZrtqawdZzzljAd4keT8KxBUrrl2LrcAMJ/1F6XbcX5KtdiczYG5uyBx13Zop
0grudpol6FYAnM7+H/XxhHKqsa0Nks1+ecbBzBm+lgKbx2lyq6vI20gIYrCP5+Jc15dc53cnONKc
IA6exTB/B3Stvck8vqd9cX1nkqT1Uh6gyX6qgsd7DWvsdyI/PoCZrgT2ULqeT+5svPphxCaq8wjI
cay76RPFl5VhkD1G5oWOSW9kch+A8DEzHgeOnuXgxq6f46obVspi2IOQbOaeHDEzz0ywFYfpN2k5
EvGUSWpTMIp2tzha1GQ1kMeH8yr05rrCRxYeKoeLRQR4jaWxW1anEFkIYouW4sAbL7v5dJIiXRy0
4DvsOdehTF3EzGiuoJYlO5bJb3lGmOZbQzaNuVs2hZp6kVjTP7XHZnfbl5ykWo3EPrpLfkn+3EyY
PwdHwPUisEVRGgiWf2FnfMLTmnyDtRcaGvpwA/nH6D+iTA5PzszlsWu6GNxN56EgLzj2iLC7HHY8
J0HHG8U6B8pl/uB/2s7EMLf0o/GZHnMt/o9gpq2ija7X2hsQa+IIOZGeTcn1N+RA9wITt1RQKbIx
Txc5k0RQRIxLO/eW3xUPRMoTw/48F4/BF8iKNRMzro4SzGy7ggSMW63t0fasLJSpnHViotiVxUWT
5+cATIsO6Oa5Ez+Gj7x5D2wnHNCoPMREwPT31joxV1Se23Gl5Ewl+KjPaOlJs3WjXqBoM7eHv1j+
4Oo+lNIV0o9aVAjxnzdCXaFkdF7M1M2p4VuoTPzLwqx9+0s5lDZRbAWcIkNBHEC+dEFVRWdi7RcB
smExtKGS0NwwNzHgF7VzDIsS4eftReQnHkatSvBR65rClodWWd/xs2NyTV5QZeuefS3hoj8/pmgP
VcivMKADmOChG+2Yofdhsi2/czNxF8nUSHBdMEMxFYwIJKAGTFWVJlSmK4j+3ewoDicagv0hPWjK
b6ezSx2wtIHlHaXJMxP7Ohnked+kKDAjXXu9lbDF0rCqN1qLDVqFpi8TncZQGaHk08gBx0J60XOH
EnghthZTZIi2m6Wc38tC/H2a0B7VvpKcjKmuHxECgtL/H4mUWnHYBKTSpepTpkoaiis/j7BMeKBX
1ptDa899yb4czYFrk7t1N2mZrOm+MS40zTjGboTFRRHVsDn3oW1oqqMkn1tmTCCDJtgrXBIp+MuC
dzMyOrz6IqnJ4btFIxoD+enRh0YEaxeUiJ09Bgru3h7IvU+WIkwqIrCrklWnaJgw1I+AR4OKabP6
7VKs+DUYRjDuEdiLtsbRKf3/1cH9SShQJxv59Q5xXYp/bTOJWOIAbbY0syyysGRYwHv7UJ6FxjNn
fEeMKOZcF2us+ApZbi1NV+eKPEKAWDtliO0piw3eIYzg0ieTussdCGtc3utZdgjSZ7ix+COnGh3u
Fh13GcTgSQHYy7sFoaZJjx/ZZh3Mx9z8OqoPjwdCjrlVxbIB+XHE7q0bnYDoCIEOkYrNfVhruqMf
XwplMf+eDZ8qPEWik0cDURvWo4WHuOb+GD/DbZDovCZCu6zO1lb42+fktsauvv+Na6xyrmLIMQ1i
61dySGkTV9eSLip0izjG2Wluaqe685HupYc3qk2vnzSbdVQPLcuYMm4ypMuilQm75cM75nMKeW1x
kydfYzBsfk1zTrfGhOtpxtSuEDpv4E0ikwSUcvitjwLPqJ5tLsKpYS2W208vpuhgKjImwm8Mx87r
lU43idBGNehqANBiNdnGjbjz0JC/Iai1VDquNPePHcC4zYcWAefJLpO73rhFIEIdTnrT/CyN08GG
vPTdBRU6n5QTgDgkMnvruD5YYP1LP7d/wr1yDS9YjmD49wkBY2hZhbjkP7ExMqgKoUoMrGcY7OiM
V/UJqSfsPbxrMVxV0m3x5Tvicirf6jxb2Eut1IYg/ueDYvUErhV89tw/69cnrIAUhBz6ZDVIic2X
3lpo/btlcNf6IV62Uz/nzVIXALuFnAXl9gXXpxoB2DjQCX/VzEW1a0xcS2mx42a08E56N9DZtFaU
maV45RSdpWWlH/iIM3gc/RFcpBuyTh0t2/iTONjoSmdO5iDCXTeVolMqDvHjQTD2Ikqqa9ReDH4K
5svfzXnDGbek8eZ55kkv843p+W8h08PTePs+CnRaxwyZnFy7pmRpWCGVTvDFi5NTCTE3h+lrWdCg
iAy8FPxcsk8UdVFX4JNbcrNrV0EzwqIon+BBmzS50DTdp3uBfAgO8Dd7RwegbJCcLoI9lF44k/PJ
9+utJx7//GPBsxNhOykk8dr1JQSbw6CXxfs2pXAIWKSLLU+lgZAx+E0Vghqu11w2MoS1rHNigJ94
5wknivThiuIKqsNXF0yJXSgBa3IAQFW7GUO7QkxQ15zs7rGlj0jIt8zOy5bJhB1AGT5iWUZatG9V
qFsx4rWg+X3oniVPUTUjt8OnRn2Y5OA19P/sAQgzGuuuuRd83IjszeZ9Da1OojIMS7F/M0eRmRqJ
casTITm/IYeMP7jvaTGWwSdZzvE9lnXnF0CqBAc6IvIKpUMOxF3Etw1HG4rsTd8LcjRFXxa+QKSH
77iHrE8aKBIQcYiex9bIpgvI9tH8Z7eiq6TBWF9p9FYwLGA/JlJvI8S9XxlkEEj/pH6vgJlQIpOh
MdyGoVEHPH5G3VRlztSC74npkPuQY+Wf9orInFxIB8rSbqXD8MUBPcNpo82QvcFrGgg/pFPPHJq9
fYtFei38tatDgR2YzCFJHc8Gct6ohP4ZjNqc5Xd/4WkZZVKQTE6hDdmK3n0VJTpcoe4n/Le8Mhpq
8+4mffKVgdi60OFGSX3h+M2Q2pVdpjFC7yJVwHOB3bOezPb+9YfFyWWYdC5mAT2+i+QJoxmUvODJ
ubbqQGnKe7dnYwRj7twj2COdBRklNd3BMI8UdElHeFCXWLgZdGFmutNZa13fFpmbWMttQ+YHMVHt
AKYpSIN2Cw8PZaLYdzkbP6FM0kLmJPq0+n72eOWH8Eb4TW/hwGJsmN/VzgL4L4BlODDzLcU+Xu69
A1m5OTxKMz2pdtDuZX7rRqxrxiI3qTE1XpYA6VdWKD5Sl2fH/Tt3QxsqcLgeWkNtpad7kAUFTFur
HICAc7vS0BN3JnVwEGYJKQ4dKBELhETJ9vaVqHvPmIg5urHfQdJMEIZoGqH0fb7LU0pqPuPKONRi
s2wWcLgorUJSss9aRmKWHG9wn9bdV6viX7nRs75K4hUhaKJRz/P9IkORyTWqWmo9f+UAVR3LrszQ
WGN1EbjZ38Iai4/Dvx5jOSNPwCB+CU2+5C175qet6F7QwjFelbGpbVs+gUR8k8TsDIhBtQfpjEqF
mc7bXvx5gcIbp3+DT4Oa56fxcDYyVIav5KcAWDz+V4YQ7HA9a5aFEeJpZc6iw3YljZv13UdXRlOu
dOe17ff2dovuNLRcsE7CtpwBcRAEJsPDgBRf3wzdbXB4WJoJnKxhShV73CSvTBW+LMUOX1OEtOKD
Hd0GOjE2INJJ6H4igWsxo/YETGcycmJWQopFuwdrzXheKU8fl/mOGXVpkIam0Tqg4pP8/St8PRmb
SxOfKIkp4veQpViKiJQkvoafvOnxrkts+L6hFrj4arxlbsRxQsBuJGimuLu3tEJ4F/82ScRoJQ/m
xB+6kswzUwcXeq5PLbas4f+E2cT4Zv+MtmEAeBXtCtl5fS776PpHzOQZdB6KQnGiEntyyPVmWL4V
pHPALb0ECzNwXiz+6WBOguee76HHcUja2iqIfvaoDVGHBAzMbnZn7cRvy12BM6E7GOTlmc6dxgA+
zwurZaKYEHh9U2XL3PH0y/r5hJdJjEQVuR8bZSecaH8jy42YOKG2rtSNTnnJm5C5SSZnIbvPnAu4
cEK6cUkIy9h3GspGncz9Y/TM+5GzdSUTjNmRd0bAObV14zdG/hXLdGVi70lODXVKfYQf4a2GxS4V
U5dq4JLjC8jERqToq1JAJCX9VSPsm8/MikytR40vdL4KT9QTfLIKQcV0RKZogyWaTgzFcNVTRKZP
d3Bxs6eedB90U6KebuhC4TP8Bu+/e7XP5whMnOLs43uWG+DNmEMssCyN6MmR7TqsJw6bCIMbMpou
I47KiAO4TWyPbQavEVZCA7Hle9sX02DzQG9wK5MhtsLeM2L1HrP37tsUq3XHo3u3meqmZmwsVjI9
lxvPbH60uac+SiSP/1PC7mCtoevuVnOvB7Iutqp0PbAa60dzU/Tt/aeWVpXxKBv3wd9kwb+jGb15
z5Mymz142KpPVv5Y7cjEFa6owErLnQyLU2yAkCNLu5jv8IcLyFi2WH+K9WfreBoniGJ37HRRmibJ
+MeXuApNELJvQfrveXvfMRVIs5Tm64dbwV6BfBTDrBuAAQhfZc4dAJOETT489u2B+UI9/VRhunmt
fUGb8urU+RY8Ifto6eJ3hofgvdclIMaT9nsCt6sxDRV4mCzWM70fQrkmqE9OUXmEJS+0OFK/ZiJD
1DIn2tksEI+z3GV/iBCynP1M6yyvU+ur4OdM1sOcZHXuZZ3r2IFMectN4PPrKxSYrJpbWngKJj4A
1FwgBC2IHg6BeEjuUAcKIf8YoXtPIgPhDCkbrl85aDfv9eA6k6ZoTDtTJNZJuISSrIoCgZLy5E2d
aF5Vrt6oyP+KTQh1aA0XSSrWqE17pWKg2O4fyhTKVOpHjOASTIZRjYLyCnqF9fRu9NhRg8Kbtw0k
mQiVhdIdHE+aZKlY0Y37KWTMB730GoGybviIcS8R/11PsZ0mEOG9gYmYBZ9M3av0qk7M5bcAqvQd
YckJJOBGc2pyxGFYl66S7ApaUomDYgfvEJjGHTeDW4HZXSrngW4qTPbRAgIstvKst6FS2uNeScIr
TqlwUXgtbZeNvr80PtSESb4eW0Uh1cqWPtbppGVXhSGco9EVvMH2xycExzmSkQ382UNAT1BaKB3x
z2Vd4cJxDrDtIzA/RgwId9823EwUpBT8AbLqxU7N8a+6W57OtgWKk+zmy5/ARoO78nRK9Ks59fm8
7AMchlq8Yn4Ix0O9moVbwQpWp36TrAuW2m/IwYTV5xUM0Q58j0rIz402osdzQtuMePzTip5QcKOP
WAgTdqkz5i/ajVPg0xs8tIsZAm7T4eeDPXVmW/rkoNvsIFHh7gOqtAjmCIifiyJUmHwVN9Vf+Rwu
w4kbCVsEGtdyl6vt7bxxdsqq9XSCyySczsSsKIaRV3wwu4lc4REyf678hbuW0M98kWz9PIdJXKb4
CdSHaS8hedEQXBdA3y5/tDWRawGfWBAKIkL1iGqu0S8U0fAX+D5oq+Pt/XutXjs78MIrWFIbQQqP
Y2wdYklRjCKzXGoEXm+Y8N479syIRCNDDCSRyfOm3huiADNbKUjcT19dreK/m/uTkoABReVee4Rg
Pjfrpyjlj5gnBFXNMWYg9IYni/tvc/N8J61lfP1mHS5v0QHNDwa3qH8AoKhN6ROq3ensf/x1HowR
9ldpuZRS9289Qn9eBVFq8LJV/ZTA2kjIuZpxEDEmKjQiu3c26tvWVt7XDiJz3nf2OyAjClUGycD9
9vnw2Rr263nwzJh6iYPNBYCsNw/YB1FTJlzCyWe22GNbuE2wRPkxnU7LFj7kJ4LFBU1l1sMO8Ngc
isLloXS5jzEzKq/FY981Yh6tG5c3JX4BmRLdPbp5sMfvNbmLnpOYHa/N6t0MPAf5lQ1sHzyy8HhF
R5zVjZ1GPcibOcX42CPQbS+WIZX4i0nZG4YudL4OOeNL+vyCMPQEhaAJvYpP9nG7H9mms6SGSxDx
IfZDcFui9faqjuzftMBKYzvHtg19bsP2TVJWA7XhZmjb7O4QJpgfBj/hAJcOGlwh3UXCrXVW/3cJ
xhmfndl2YWD48n59cWZhMMzrmwVQUok2MvDat3lzENwba9uSwREdc8mY+5ReagXGvfG2VVYUYrqk
CMSgWvo7V/Ioa80VkTJG7f92Fn/eNQfR3iwrn+jILEvAnN0nB+rVCHYTl+YEdbr2SEhqoI0Jf74A
HVqjRGEHCiAXeFYujf1DO+g0T5GxtctK7ael7Us33AZhpeKPgoaSCs1g4JLKgwlE5wan42vMrFzQ
MwQm1aqoLumQo5DTKFBed7whS8oHnGRucruaD1SodBr8QFQxl04mB8xxdCOR4a8Ob58SiQWWowEF
Ri36iUvqOr55E3SUIGEUr+ZW9DPjtqJn+lY8eIpQ2LTlDI6oa1Hysfw3PP9xvJ9w7Ycc/39W7/Io
ffkV1Pv+rSMlbNhROqZbWqZ3UVqQb5WkfHHDnwQ6F15maHWU/R6hY2i+aAEt2eAubM+PAehJkbZZ
YiUfkJn35Cpx7ZWzjMbPqV/5wzs5yDFP+mBTXqKn2aCiVD+v8E/hbSgMURj0TAJBn7DL8v2FvNVg
J6+0gPjksq68hUDNsZwjl7c25opMbuYg34Q5Kzbsj42Do2T89XPrluQDrX5yiQ4tGfFLGZsB1LUF
0eumSls9BkyQuG/3r98vQe5VG06ShDZEym1kRJEZz92Lsz9bmVV4t8MW0nb9h4jo0kkikoTJJ5Cv
IE5dpxq1lBsKwP/I1CLTYnw/qmcz5zz5rYQF+FCinTjnwhQjHtmOFAEfbmqdHdcsLjp3naYk2HED
j6pTbYuOiNsG9kKgKn5lkI17QAirIhMQo2swxFeRul1Zcw5ffYKCEns3ydEcXoIKkyqYoXAFFDML
E3f838u/M/2aZjjEiQotbFCvHvgNn9yskuG19o/L7gzof0Lx8efTFkmhWfTav8AC1/E19pWiFXdR
JU4XekoVeduYF8wQT4aP1Iulp0l5rJB4Xi9jMWRvY6qQ2oyN59kU2HXUVfwZZxhz4sAXn6hxtxCA
vXm20sDnqpxYpA6Oybjgma+v1+SZgbj13VdsD5ORpuwtEimX3KluM2uFpb/RaTq+CRoqimxRnrZ7
FTWgrAMKDDLIf8PE/6oZjQh/02f+Urmm2luDqPWgBMfacKxPpOXv0+4YpTC40ZGnAwB9j8gDmL+L
8/RL4qJgYcbE7GWROzz80HVxQBWhqEI5+5idERhh1WsyGbgVjsMjL40CjTc8m8IZCus0FsBXhUM6
HgRiuB6TiXTPM3QAs9p76yQ0IwAmc935fgwyVTd1e+1iYDOTdroXHvEDzAIYP2uvn3LqBM5jprl0
4z1eNBQFBEHpCBtyU6G7B86KL5XX9ybEGw4lu9YYIkZstYCNFS+wBZeRpat6nBYFljIkO95QDFPj
/Hp95eSvSPPSCJv1qhmaBaLytRXamlAVjfl68fbaoIIB8OZT4SqecQ37wLmno5V5mu1qAls2ecWM
OxrrOg32pPk3bO5vhU74iPwe3inev0hsqXvAMFYk8klvEKdylewsldUgx9So/OvvODHNAIzFYKR2
8GFC5lBoxWs7uY0fkw9/zQd+Etpekjaw4c5qs2X7Imn1buZt7Zx+ejCpUBE4Mh3+F3LYfUv3kisY
aK26e+6ykv5nBkVidiBZzfgLGG/crMwnGx5PY7lz9I1JLQqXo4xtzN9WKZQMGF0F8PtokeWY54h6
mAxlxgOG8hyKxfmCG6sdhJGlyCJeIJtddWPij7u6gs+w7O6C08jKkSgxILy4Gxl33I1IXFrqC+zt
MJrk0hHgmDnkUbqm+S2iL2ZP+PTTj0aFzocpRL6Nr2dzVpNv9EbtOJHNi8WGBTMx/oxzzDVg6iHm
f/ijJogaEotDYrhI0yViaJVOEZUe/V/r2bwfNfld5oyYEHS9MCpRDP58+ptRGKbuib6eXXlodpBi
jCHKOqiiimysCXHgcwAgn/zgTwPnA6vFDw5Q+E0G371QIGTmktP0H9g65JSycx4IoCigfEFhWzsf
plBngwVpOD6UZlDqlUUhuFgHvdCC2R6V3YtZxMLp3TVv+89d/tTO57R2feZ0vJqC0j+sDJDbKlUe
9wNyy87gRGLqV1wFhHWUeAkM7mxaMO0kgQVPaS9XtciMFQHYDzD3aKZAq21xQsDqdVNE4egv8CEH
5Y1+euDHbBsqlS6c4TpZfTEC1vsMHGYzBhe/6VqMjzOYT3DPFxzhdGnGUA/sq9vRnTvXNkpiYgNo
gJw1K8/joVcVXmo6Na5FSYVEysevtj5htoI/2Of2H33scFy9/q+YUQzlx4ACo94vc00DNhLIyux1
WVnnBbhpWDmJkFmuGbTuYGTBWljTIOfUUbqUrfLJeI7qmFFsBj02EifIjkxRjr3Nm8pY3ifqioMr
XNaWIh9qkDCIId87/WleUE256W3klXMJq+iZ5xvM4Fw1XCN54YZ6I+SP9yE+j65u1uXxmHm+rOta
XZ/QYmprp+seGj8V6lSaxAKJj91Ugqu/CDxKgICtm94sub+Z+FxdhtCltrv+v4k4t/V4QWmudIbW
uUYTd7lr6+wGawuxUhxi3CGVJbIEHZP/LMEyWYxh8M3saed32qnmyCPwYMoMHaA9Ka4oz5SFbH6T
HZ8UdhAjDxO3kTiu81c7Jty7Z3KVmjTfTS4nxM5oMz3+Os3Ckg5EbzM36gyhJ5+MG7yFWY0kTCpc
Z53Vii+MBwusyNi4/P7PV9qQIU7878is7cJqm8wQAVyRx6AOx0ms2DdyyhAoOMrLWxfunQWU3hha
L/EJAQUZXe36ZXS0FQaQX7USbas7AXXkqIBUOzQEFwtEFIvlwUoeBHibPTrNrGvtdp5BAkBCK1bz
A/P6ax97CAjkCLKQRCfE7KcEQ6jPnrq3EatgVeGnOdxaCfCp8siPebRfCGr7k84UpHnoQG96+3Li
fLSj2eJPSAyzT3gwdy6Bk7kFvqGBwfVUWVbsI5r6WU8J08Hd9l7arBXiQIpLgwbVb+rgvv4k4zuk
9z+9ntrGrRqABFKEctln0T3ynnTN447/hlMdrY2ATP7xlZl6xGJMLpqMNrpWUkVNCwccDn2hiDMq
guqQGJ1mbG2XCqwMXibCVKsmHUFrCLhjdT/BPcPovuN8BRejBuHD/p2Ga6ZCNLdcR2aJ2qLOjPrc
yioXOmSTjtJOTdk3eGyAJTixw2l3DuNYMrohNPP8TN76V9h3hnago+Cm39d24UmKQ7zx/V6LUxKY
H6WLy7KI3R2H/7gM1QJOCWloV/okMYOCCEH5Zsq/u3qoLxi+7sNC9i5nQL1db3jxSjb6mDyoz/Dt
QMlHhMjnj5NfLpOfEHQWwOGCnQJTh3kmyIcvz3DWs4pFQusSL7IWV/CSsXTkebw+0Qq7GgnXM3WV
cPkbfcYJhamR2PYp8mp/9+SLJB1HcFJN1vQEfw9ebDoaP0UtZDkOOxbkRAh4x43NhbXKpxvUE4cN
LlSb+io43UI9LZz6sJb/Yr2kwaIFLo0G91j7dkUesC8hJJ7uYVuZKIwPtnS76di6xFsDySL4Soqn
euU0F7HubqiRePPC3bjULS4XrKaliP7bJzFg01byio5mfU/HTLIXUzABbyuHLTYxtAX5C1jaReJ1
Yy8wUJgbY2Sf/kH3xhNi7H7/6jHsGv7uiUxqom8csrHiBxc6VXLRojVKsaahOnM8omJ/nif048k8
3/YMGLskjwL1Zb//nQvRqMBAvz5E1r5Izxn8OxVZ97anq59kDIRMvPwZOcNO3EopYlq+/NyHn6D6
DdAn/+VjqKDhYyeyja2SKx4nngER2lbg3bvuSw03E1kywuSFwTpR4Q0nDx/lF2883G3qzlthElR3
Q92M5XPx518BTok1GNOLMlm4g9PPEUj0QHAYIVZ4vIGn3Tg07s4yQLSENaCUs3+tCbVzp2g8kcZS
aBO4jbuWI+ciIaXsNsFt/b7jrYbhC2I/dXiCM3MTGDEeh1jQJX8fsggg5DZYUFmeRNSr1JbzdmpL
aN+v98D99GCI1I301zPMT6f2DFb8Y49zeI2oDD0q3hbjkDdoxAcs76/jAhUyxxTtU7ROqwpvj7Ni
hWFqzejnL9h0QKThRJCeWF0RAPacw5UGUpovoabFiSlL/AZQ5STBrfmPgV0yCc3qhsMPKeA2hGWl
4VTmFPjv3cOmhVA3xOZu/IW88b2xrowVez6FiS7Rocj4qT8OT49ZnFKPoF+TI5Z4y5u2ZExl/8Gn
wVSG0FdJCBrT7sVGUiowepPHbLpUQvNH/TrqiDQ70HiWSzrz6XAYl8C9XZG0iO+Refxa9H3nRzKB
Yqcw8uEkKzONCc44NUVYR1ffPLjte6gSX7HTYOLcuUr/FqsI7yO74A9YvS2bEbKFxCXUzJ1umWl8
4mAKPaIBuTEJ9OYP4xVOVvBsaDkgcs+N6eT/b/N0zff+A0cGQd8nvEyMe4J/HEqe5lCXzPMaKfxv
M3NgiHIIu5it3ypZJRoPlWN/2dCxbK8MkiuLeG0IEAm5BGkB5hsJkrB+Kiw+eZge+B1xLdIJJOK6
sUgL4gl+oQ1MtykX08Dhe3/o2n+Fkfj/6Jb+QTFoUFaMmB1jPl7TQggFK/zN3CVUctqbPX/wWiEd
jKm0o8n0c36r0iIcjrXomvBMDc+C3F3hml9VWWusHTex6qn7ObWES3TKcGaTTZbXn51/WSKJ7hl9
23BFABOMjcAxLWgK7j6kB0XnHBTcEIwsAiwXTkingD9y9ixNOTGK8L20zKJmu03DU6rGunS1qiE9
g//aBu+hlQLLSXHXXMVgOX90gNxtccCFYp30KRkxp+62r41meF4Od2tk2mrlj6PTe2zGVX1ptAo7
fPKR3BW/TJjeMBbNYhue04Pq5LyNMJucsRwn4WnUa2JY/IDJwL3Q0hyO7lDFGx0C4aCwlLlc9m1g
alcGwcFa34sbbP/ixJlwzMfRhxbf+aQi5Ny9iETnTSGwn2HbXouwcaKqoDx8/Snwllbs4kamhfx3
zgUz/s8+W4yNsDD3ebGFdfs84izn7LatQ5PDopR5P1dXVGPez2sLt2OWNBrwXB013Z9mzZchFlha
EZKPguxrP+6HXjbinBkMdG91RxGyny4KT5dROEHxWxzpzNNw/PJ1BMlUa456d6mKjw19AjLmvGEb
Zv72/l/nszkn8qDRrVJe3Bh+55HArU1qspK7IrwErq1mGrQMtO0ZuS9eBB6/Hi6ONEjKcxcPIy45
2LyouwJP1d6n2ZXQZnhO2DirD6OnSkBU9i6mkNAM923zuXqo287jMBX7C3mxW3kUscj0r+dxFHw/
odanNfTqAQglOzc4fhrAnZa9loj1RmkQ8PeGHmIN/dYCiB2FFJcI/nVbzAvVZlriLlP24QLnXLMu
ITHCCHZ1nFvpyrzT+WZrbTzG27PdAX/Tmx00AprqnhAYUYwXg4GS+vYyLQ/Ep8xTUZcMN4KUS3qw
DzUWoyMFhSisi04Sw5+HxvIsH087Tz7m/HAFSXrXwC4iKvE1wdUUN/og2iuVdzZpwBzwlMRKGzw4
B6REyoNTWOLEV2+euOMxNNj3sBx1sJi9VxXdfnZIIWNW3N9b1NK13lcw2L9sbxj3hE2b3JQkfyZA
6BCyNUxtH3w02es/pil8pPt/QaVQ8L9XP9BpbAO7jXQzgArT5VcG8IdRWEcOZJ+YGfmt4CNm4+XE
LKidyg24kcb8Ncbhb5d5v9SjlspziR90C1GJvU5V+skdyyFCbbEqQKwV5WJUDkwI4Q4Mlba4ymKZ
0NTLoaSHIO78HAvICgL73P9LdvYMEefv9cEA9Es1/PQfdaVMFSiML9nIZwjP3fUpJ3dHvfNKTdNb
KsCEd3/uMKj8Jx7XqeWKYTJf0dH1H91mbGUk7Lo3vMZgBbod/kOQgbawbOXq96qjrmamoigrP9pr
xuAxrpCMfr/Ev1TEEMbdDX+WfKrBFG7GBnteH5SlyJ7cY0OMWUnzD2+Aj2dMRfBoM5buKqLlVv7G
7895ZTT1p+YiggwZkCmLXY8Gj4Oye4T7NCrkD5zBzR5Z+unvBOgCfliJucEpfniGkQtrhDeXrFLg
BSaI2tIYT1GKxXXzwlpxYsqReGbLGBhHLkjPfCHI4runheZKtFEBvWLurC+/A8L7l+zKRk/9/wTK
UXt+5Vv7ELqwdwMdQ/XszsbIsbwtF79M2YE0maSYIsFiACBuodmFyQs/kofUUFImHE95PhlMJcR4
DGrWfb8/F4FpLHWBTku3XGMOSl5xdBOlR8K88LOYumJbHj/8CynVQKC23GqvsFX1gW/0JLSi1AMq
bCweH58T5YPh1xqgghvSjC6x8tLtFzLMiL7hw1rSsu9+4zyRom/ZlpCmuqZFJDmPalVmMMRRcsBr
8LbDutZ/b1sltQgn+U7SbbAZt2Gb/Jf/h9InHCLQfMvF/bVlWIQKZadv+YoKo3W9U0BW0J2r3Qd7
gdLCiK+bcyJBGgF/wNT7oremlxx4PHayGxjtirDFtVRGW24PTCCbwI1NWuiG0pvKNRs3CZdpfP6V
C7G+ajzra5rF10G/jAieNxwnvLgnrBjkGfJSd5G8Oh5YRcOyd0aJn0Vix+9jGg5jU8tEdSyt3GsN
7qOcABGr4ZFX7+kQ5W2GXWlaMJnWchOvAu5+sZPe8LacRtxEusP9gvuY8cNnuSp6OwBlMM4wtTJJ
bvjiiTJoU2GCNym5uBMNkU4Be/vg2j/4eigx2HgkuBgCxvTWVQygU4HZj5RarkytcYpa8nqHTnBT
GpRnlhIsJQDrzE4Q7uzM7BKqgV6f1rr8/zyA4085jU68flAgogoIO2D9ajKLc3b14XPI8AqSIzEY
vPtioKquIwv0wI9ugmAiwYbmnv6G+j7l+b5JmYP8fwdqs+l6gErbnYbd53EjFf0sviq5GUzYfxVt
HnB6VlbsMIp8/FAvDRLNo1vQn9SvzSdaVKl8dW1HQ+1w3PdtMliQncjOKemZqxf03DkxcCB/O2Uw
b7a9vw2AxYYEsXVkhD/EBxN+CLTbLa4ANVo93FtcNiPwIc0Zqh/WHxFnLXLaQvQ1W7kxb4RPvgMu
+UjJ9v9nvkzmvPVqg9gGdA8EDIkLSUZVeikadLldmlWXhmjne7uVdEA/MCEgSOt8VY1WjCa+d8Wh
/NBEgtPaaPZxFuEsHIXmY2WmCyflUUg3CAGiw0F9fu6I1cbsJdZH6Xto+CniEL+ufIRX3PKBBhmU
WGvz9n8iJFrKEKD5CbU/w5kyISPueRjd1GYfPvuTFzSbuuxrNF45DTZe8+69qAUSNltFtTEj968X
c8GDoYbKRF6GA+2lSBhxApyrfyWjekGsZSV8uL/GdpCV6+cEEJCW0+qyXkg2jW9BS9v8wpzzHcml
//X6xDrE8NFcEf7a/qh8xlqKdTL3h59xNASobM3LR2nXEh/r6UCn68kjNSdrC91gPHKj23sL6srR
kxotFX6vNu36z0T+B4TzBxd273x/HJQAk2YEGJXk+3yfPTtztICmbIMbS1nTeYqspaShPL+Zfq+9
HIvwvp3it2bniT6+ATEEMSj4Hg/QTlwV1sGZq8qG0dUEEdh1NQZvoIaM2Kthb9sbPTvnoC4+xkpN
gG5xCskVFdMMFBRvxiiZgufj+jvSIfRJAunIJayx2gWXNc7PEKRF9Yscbyk1uJjhKh4+g0FBQaC5
MJcqr6YlHpeiwjebGgVpTa1Opz6zGbjsE3bZlmTjvmXpK+bebD2ysnZ2vT6OfNIeBt8dhCoVXH4m
Ojce3DWwuBnq83F3JxnEX4Sc2g9984siZD+zQY2esO1FozaEMzAduwuEG1cZGIUF+T6C37CXs4Vh
URxc7s9grM6UrkVzaBznNwEMYnyzZiFMXuV6KuvXzsHR8IOSxNlfAKaVP9T5S1T6qX/ePMFNDdkq
LMEW+04pN3HtCyJQoTQS2NbMlZX6digeeM9GD64NPRPlrDtz5cAzU1KAAq5n39sLtuT5Ma72kprA
HE413Tg9Nj+A4g61oNthGdabAS4zxtGoD8/pzYs/UJlL0r5mNZXlYN3V/ymxNrshGdRylBq3Dx/d
C35NRs0B+A8FHdvyd7KaPVzqbtN2ecAlWUb6cWZI+nEkDEVhlbpYg/6jGnTW1VdOxAJ/xxxJHEHZ
qMlVweLhizMqB8ERllYRJSj6tR/Bzi3bCmqb2qFwqBJhph34q5ZI1h/nyqmydH3F6ZrrqFdSLRqY
0Iv511Yw7vR7AHRNkyFr2QO1XQ8knWNfpWdpcKUbWH/QVqPORV5xdD1D6m292fLiGoZShtWva0mt
35ZxPnQqz2a0e11ZKTGeVldA4cSZgFEy9TXzei/Fi8uK81w4ukIITu5CjqSKDOX+GJrFSTki8VPG
wnRAVJ7Jt3KDbV3BWd4qITGiid6L6Ei0U3NfYOySUj8Ck/d0ffe5d5A9gysHoBiCHtQyju7lDqDl
V16Dz83T3yrCCW4jVfT9D4WSy7EXYaTr/k3+wPpyY3ZtaVjRVbi+gAbgxm2JMm8yRLQ9V03P3goG
A9+15yqn5B9j+XXp42pPKniWjdN7psFil2MTfIBBheCp1f5F4PPqKW2M/Jx8mnwnk7POqIRDlxJ+
mgdTLKxIn0j4qkMDg57dPrpqyGihMrQcNLdTTT63/Uz6XVZoVMjwiApgjk2EPcPAwBixV7io/2fo
AJ7GOGALEunX6SAJwzAkvIpXX5SaPgvQkLuHCMtb4mIa9mG2hgk97RprzYbE0OFthd8srWA0ncHa
kJ1628BoxH1hrsKGJ2oaoCsfrGVXUtg6fWMa1WE1/6E7ofORgN0Guf4TeCXIjQCNQ418mVXq3vSO
f0cxtGwwTYlrdn8n44dTf9+yu3C4SCCpGqYseiOPa7lMZCMPlGEqgnSbJTj3dZ3+CORouUAZPb06
1N72k8mrmFQPqbnAEoDXCUB8whm0Y+cxgnY4jLMDRaE4yA/vfweCdBRvstMvaEmsD82v3sTj09/Y
vBzGkYQ9BY7Q0Rn831MvjyHGC6hsL16jGKwAvoOm6mLdzzz8EDA3SzsiAqoHGV/k
`protect end_protected

