

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
qm+ahCoXbtCT96FlU7osNjp8Kf3rDAFQ8vMBTpaKgTo3EvHN1CM/XiHNcIsmMQ17hbL+pWxo5SQe
TeNJ1GZN0w==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
KB+ek3mkpx3N+ihSLNljgKYzWfCbUQKXGho6dSjrHEWrzL9W93J5UQjcPdLkP/4r8XQ5AjiJVm8G
O0+WgdiO6dbDdWggVe0UZIQ5qp9jotaT15XQQVVkD2rcK5wquost1xsRm7MTsEsCbzkhqKPM6ASZ
mpW7GzuYQ2vDPmY/r9U=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
5IFnCgXf/KjXBNbWCJPfF+u/Xe3PWCvLt3/lqQEWvv6nS2jJ8qz3O+bSiUUxyt/rlAZZm5DvQ41j
Vn2wE7il4mdux1L3DFueP8Ob6UEbh6yobetr8hrEOpbRcnmnH7rXtvR+yuK3psDEpqbW7d8GyDcy
T6jGK5xIsUceYrUwudt7lxYx4bLnzP6q2c6uLhkxaoLJTWJGh28se0dzlAMX/BnMMfjK0HDKD6kp
1VwH2Gj4iT7DvyBkDmISaH7LPSlLhe+ZmQMkilflhi03bS9w9ABaqs6v4fufe3/pEUeBrvl3gRH/
oCU4QtUwSf8qfFsWdX+C6Nn7mzOb0WSGIH22+A==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
BAf2bWZTeSaPIqnT3j5aNO9C6t5/rcfC+/QtvmxOirWtcQ57aHowXlt817D+9PTxe4qEx5CjzmUg
9oMYSESB8IK4XXnHzrwWEKN1a7YOhI72J3KxmNssnP6jdEMx0znih/oPMXJaAdPPRUXzSczvXVqf
S7AhrmorMi/7B7tc1xI=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
dVk9aS2pcwcb0BrWR4Sm4FSW8QQWqHH7xHbqUaQTDLyPydXvHmrmxiDqUJWu8AAmbDSnHtBnMo/b
vhz6TIedlqcgp9o49Jh0CEli94frA6kGx65vbdl7q0c/R9+UB+XDf9B8tq4xwdSd4Twx0zVa9WGD
lmNliqJyvFk+OMbS2OJJyBNqK6eZPVzKMFkUG0UJu6TERfYV2nuxVMsugR94X7JoKx+W2jEprOdB
UQVXsqhudTLpaKEQiNqzDCaBK0P3FekkJJMtZNaV6veO7wX6Us6tTDs6pxGysSo4e6tLocXysaO7
1blW1S7foypb+e5LTkDXsQjIPmjtBTMz3Y2yyQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 47328)
`protect data_block
8CFrIRFTNVOf0UHFtrPdhHVT7UMAV/ny38Ala2y2oximOAZO3HWv72x9fRmBGIUoDHr3tb54Z9dS
IT7wtYKtTRcl4X69X2IrPACVs+WDmdgBwJDAE8jA41XhNPVEBOuVdZNzG42fs/TAl9quWphSIXd0
qEmp2ok6Nk4jpQ4tuAXWh3IhVZ1/aZazY/1kMckNBXNz9ZxiU/gqD2i7mA4bybWnWyIpuZluAOlo
D59qYPRPhUz9YVF8/bHM/UVv12xwhPHgCF7a/MRLVFtYmPMa+D9qUyC2lYQ00Vdqp7PbZvQgn/Pj
XrFKjcu5BmkFk595Owf+HayQ/GB/iTcVoFhakKV6aMjik8p8EApojSYS9/4NswEyHrUIDi8u5b8A
iRIP7NCCLphRpz7VQIgM35osJ9yOyKqwH47tsEZv70SdjNgK7unyKCQUyMztWyJvJLCwoWtFCQqb
qqfj3EwGPgTsd/TST6S3ShKOWHgR+U1ecTnY5K40mhrCi5FZD+aWUvlUNX4FpnAFl9NF+0dwWnVo
I/6uxyzy7tlMdvUAYMg2yrxwarHosh1p7cpRcA5fshaUSmg+VzUvvB+m0dlA/qfr45xYaKcDPkw4
F6u1FlLY9BPBRfYEEkN8zc6IbLn5tr8c6UrDN8I4taHX1mGReeLeatXan3kU7jXrdV+WQoLIgOSX
n8RP3QV6I6btraSYW9DEXwpXhJVHvsPcRvAAOjbzHx/6DC5hgwpymWf16g+VygseGBjEJY8pkYip
4LtOBGUs4BC24qVDzJUOF9Oji1S4jUueJymMUE9Id5JjGLidPT0atGmyzxWp02wh4iryI2dKwsCh
wJ8E7Ot/0AsJYVNYNiu/vARo4Ak8n/xTB07l1UG+wD6DAUNJWl0uBvxr/JMkMbuH1ffAkq/8GgYF
oXZFrzXZ1kw2SNqHPVzN1+9YbbuWbn8NU+MpDVkwdZaV69Vu/jLLCaAd2PQFeTeQsMt3gQROO9b3
6yQ1BRIfMmQ4gB1JWFEGR/v5bXmKXuAz2aUCYesPNN+1XTdNVfhIbIfDp0QtuEXxYELtj09LZTbc
S9hOzQG/S1xgQA2LZ+d7m127wClppmMJJ/WxqGWVpKlC3ecrlN9KTFGwjIzAEKZmlsDMLkb57bPH
ezFLwNraURmwLaBphBkkwirnk8C4XeQ/QfBDQMUWva9VSL33AUhuAGxyP9KpHkQD+LSiAO1ZhFAI
jiio1LcrWEdva2LsOH48qsyiCET76Q2TcOfBXbNfbUmxHma0vse1KMjMhnvwEH0KNESq4gfzsDuS
Nuy8plKy8dtFfbOdHvyRlehOfifYnhJoiQPNYyBLacoHEEaO9tHmf1r4iVcdVUvpBK6GjfjlIBSs
qCQFImf7GMFcGfOLvM6kG5BLeqHbuCLUsulvdp/h3OywzCVMxJdJ1AiFVzM6sevXj3f8ldmFKert
zrzk2fsQxiuL4UuhDct2HDlES8yyD1hnfpSaToHv+shvTyPmYDiQArslAojHaYRP7iFeR/pmNU1P
RzDYJPP6XX+Yfpih+knu8/8orAAiSMfMYo6RL4lKduQHK5B5IuWfoKMH/1oglVCgSdEKmZMhJYPI
nwDQHb2gu2InOu/usegq4f8SI25EenucjOEE3jJ1xhud0IUL1pErNNGQYFc4CmZFRP00Gf2wuFvW
p19ANQWsSJ3MHZL7tB8m5sNQzCkobaulIiIbod/u7AVrosoUg0qxcfMb+UFUQbPxVlHEG4HZbKKx
ERIXLxZaQ38CQnYdIbVgA2naR6J/S9lk5o4AnvwHRNASM9r0aonwSZ5wJZcBXvTSHqA49sEipkXX
xmxBgP8wA9UE51s75m5U9addNHFNSTwV/ifzvlnye1oPux0dPOU5yBZf+zkbPlKn5JP26Mrw7KQw
DzW9ve8Du82bQ8vHj+u1E5Pt1R3I7Js+Rlq8uY3GJEzTn2L4ua4sHSH84YGkjWXXnoZpEyczTfbe
nR9wc9lQcosV5bFSKIIR2DCVda8AiawaPs5O5TSuIbfQaAAzKcUB4fZDx6ETJF9+7m6tOs3jEoAs
8OyWjybrGxhMSI+QCc7lpKb0lfyeaxCa2x9zbIaQS06eoAZjzX5jPOwKP19ShssL6nZ3XnbzRjQS
/OozQWzi87GBwNTAiNXPYfauD2tZoP+LRotR1M+U0O/9jHd7/BSwWg12amv8djIyJxvFm+jCs+w5
IMC+kLlFQeSVpZHnuYEsnIMgFR0NdBMdxWoONXn6Kar6fi7Jmo9VqYODcGEs2wWHHqaov/E5Bje0
AZ5HikI9rdUdjQUnfHIpiTfcWeRQMwrbfo7N80PaxT+CyyTN5k6NNRgSus/9ajN7dFpytyZQlPeG
coNjMi02q70r5ixIRTuRcGa5y42jG/YY96zP8LHosVOTqRc/umuGR7L5fDPH2BCXbbgWYWUnVoqb
Ylm9orqPX2satCYYdsOQo9LvHjgZqKvCFzNM6XoTVS3eMlN+PMri1WMdQ/ZhcnbaMMNkhRBPo7lf
RxFpcOdAXccNZ6xzXYk7A8jLNQ+pIQS9pwr5tFsiKu5wTpANoQBB0FEBh1KwLW337pz8F3UEr4kr
zyD+49Tj08mIYb2ppWpYvDNBRoz5IcuyutEriI+Rluz8I/IgE96KFF3voJM5FRE/t/NM/O2rGZ/d
Ie86wxrTvfERGM5pvo1uQQFk0bA3SpQ+EfyIVD3UqM4qw4ag8DHXC8v/9A3sEQXKZGPIyFmh3yly
FA9X2aOdmIjjlWHPWZrTUE9VtXRrNoW7FmPum+DXiIii1LmkWbOr3GMZ14fRQ0aKn2ORKgZQyc8L
6aEhN/e6sOKsyBkth6Ne3sx28XXmA7cIZftJ8SPsuqS5n6dn3FYf9cJuJDVt5sJkFRP3vHtAolBF
V9/0g1P9fzkmv2eAThmf+mF9iLK2BVx7Ce+H3Af7loeVF2ir3Ez6mMvLPy46k9hN6AstIx7qt/rR
25bi/nQEQnyN+n8ZH7e8Tgpq1aYTjTgubS8GftwT2w13rQsDiBQT6PjSoCs5SomvlBikkRmSvql8
yofMF7Tg5JYaZp3ysDkOrHPGV/XVO9WjLfH82PgYP2V0ivfcajRY/3oy3X7TJVS8dRfDoPsshlwI
cboMhLeug8A4b2g8PRMXqcXVXXNJTr9RBMAb0mRajEq384K26vW3IqnMUmiqgVHkwRI3jLlNSVhk
dIy8hjcI4B3GjeeAeEUyYrjOdD8VEx3BPE2HtWusOe0GFj/fjwHc4dXZhX/VWMAri61sMo06ElND
l3S3Dfo/37wTBaNexgP1F388mDWux5pCRNbt1c0ctMXPQ35k+8z2AAPNboSgKsMhHis0ovbz8uKn
KgKY18NIBak75f8VFP0q5gP45dCuC7I9nFbWo/9a5a1p0xscKPAz44Pedhm97rzjtaK4OcG7ZGRC
A0/EwMcrJTAEDh1VGZdZbaH7YEbhpOb1FgWF1t2gdZkmKX86VPjFP8dE3TJona5J3AX9wvgjjlsw
/+Rgc58TDVnP1/h4rvW49Rxmy96L+V4akq0OqxFDdkVdsCuBfkaVRgK/ns8p9RI0SO+QO9KNoEit
NSbvGi0SnRIlE1alr1kxMiH5e+hG36LDuEWOFlSsdnWhb6/g1Rspp+etgz3p+q80Ig/GphYyIqz2
Ohl8OK+8ubfGvNitCAoCvbTS54L/KbQP7wUrOjmI0WsNXuqUHfwq2uCKlOLlIQ1WAOzaQUgt6qGM
prCqQ8vYr1vDiRQJ7DvnD9LMGyZxylLcan/R21ZRTUhiIAwSQjw6s0oXV5xLBNtnjSHr78VSbV5q
jhiKQPla1mpGvy3aKLWpSqNSftTt/sB0CvdayfIAYXP/3Z3jPV9EWOTMvE8ohbcHloazFBHL1S87
2MkmTp85IIqd1UAtKbZ5foqsM3k3etn8YGXKMN7nP8xE71lBsxi8L+Hsg6HPI+ZejfOkAJsFKwvQ
XLt5rTavG1gZD+sogUTu1aHxfKVraqvSeA7bVWOZAy0J4WZwH4brMu1ejGPMD2v75xsWLLGraQVK
nGInivxaapQzytPRszPo6IzOUZf5IIes8BLAsNTzkb/+wwswrbh9CLFVZaEXMeloh7EBr2xb5xDG
BjtiZNeHh1QuRNvyIdlmDc8ChT4MaQtar9dIS1w5a2xSJWhMqTgfHh0yXGqY7tnv9klRIgAFzrGg
Wlmyo6xn+qIgQO1OAPja5ubVi1vvYm7qb6ODKl3Y6lOVRYcV341qmt8JzGp65HwtspJE4JOByZ/M
9XqfhEj7zm3fF4i20mXtL9nbJLjHEBAzWBiPtjkAav+Zwj0fXOePcWOKyMTLYfq9Wz96lo5Tpmvz
W0DfhwcfX6ApXA0WmbIg3N5MXbx5tzVJEB40XVwVQPXYiGt5qtoASjwsWhblIzagigvesrcgoDK4
ndG9VOdeky+dD4SSpnTXD0ZoedTfJN23M/b2dpoD0XMsF5remWr2iwXl8zbO7VGI4GD1SyhVJRtQ
DDubFDl4qUnngsuTdFJhLv6E/6DU/OiXLcBnAWdXBq21X1Rp1oUwOFH6kfd+lC/VGlBLIob3VnjG
I9l0JZhdKDce+cvpWUJ6G50/id0kaiK2fO+OCLP4virLSXPfxnHtAKqNIquhFFcF20UElii7ny/n
LioHRIcDALuKMDXsZK3wG7mU/cOuPEYfxjzH+m4R1icPX0849ly+DMxqKgsVZOY4u/5jWD6dxxhM
bCj6inV3A9KYDtL9iX4Nm8zH+mzl/sY0S2N5OaZ+uqdDR1hr0VfSws3tkdDjO1N48715OybQQMDu
DUay1KqCl/xnXoFRy7LtZhUG7jvRdP2mz7wPV1QK6X/maX1r5Y8bQEZJ00fCJ+lWioe9yBkus1rq
xF6NogIzC/d6GuH0HLlxaF7OofuGTPK07yAY35dj4yhKKPKTlSctcX6Jhg3CA7XW5vglTagOgu3F
IZN5IhCfPu60EYcOJQniZk75rtQ862b5ScvoSmpVjA+SJTFS8/98wox1BM//A7fsNRMf4ZMIddfd
6a38hq5BxtMj+TgQ0cRtcnKi25oV5VxlAmIuKYggi4R+GwOm1zfSB2G4Qk0X+wGU5F4b+hvgmaPb
DvJMoAobSowuIU03X07IKLcoRPpAgowIjCDJjHmZcAiYEJ0BX6rcJlU6yJvh4EFEHzGNU++8Al8/
8eyHdsBHksgF9P4ZoI5o5DcwdFl6/kGrh0Y2lH/xbrJsBWI7s+T7HcmTtVo2SIqlCmvC9xOmqKd7
zcEtUxq5ZQgHQtYtwnL4Pbry43vnYmdv629GrcebaVht67fRclKBdyF7G953TVxaDFisGYNJpYr+
ZW5Jzx+dHAnSD8MdxhfVgvDeDRzveKvCgrLjfkQwlZpT9nvg69FQeWkKAtjrPJLklF/DWPtUc+9c
8tEPejWCHVBY7KAYE3USF61fLoLiwrhxQsS7bVGVXftIb8jBrWVjOTOdMNlEQv2ix1VQB0VqU9sE
tnXIXiwqYL8qeAsNi4TDpF/JodqyV3iaDcmWh95j3ZJpoiadNOvbcx9sEdqxDD9f4OvHWyNg6f0R
Oaxj9405qM5VlohYwd6+MY8q93y5mESciyS6knYvZHWu0mo1HcORCPNSJqJ+6zN6b7ToMkvxD3AS
nAbIBYZVWR6UUWf6iLeLsyY0Xd6Z+KHwQP32D5TzOWRRz4Z2TQjjcQ6+pXaesHNdR2PsW2Dd5pIZ
U1n4etk6EcBZayq7/0gsk0Bs2dhUNssFytWgY59hnzOjuYxkKyD0vZkHUmQUUYXIVUiiIXy4zMKs
UWV/JNK5QYyVP0w7Ib+1Pr2HF9dcN+VBIJLQ4KYIY/hkswP7lpYs1mWqnZLjPZF3BdmrWmzqVbUb
SoYjm0Rl6l94HU2uNqj2gOpn4LwP8DaPr3yhOe3HY9+vruRCo+lU2JGbCnD5Jp7VN6QzcKZ8nNMs
wxbij3mNxPFfjMPIytFa+98wmGa1A1XhTAKDYu47ICh5BR9U9lD6uu+RjVeNmqijpNxJqsKibhld
WEYFAXCvy48rYOjf1bIDwaSwsrkmhIY2Sq2isevFBQ58UElpVMnWbc1woDWcYhNJuzybMjZiuTB5
wg9pFA70StZNWsQyhs5ezNF5cm1WxF4MTboB1XCPr5l4YcJ7FSt7mKSe8Cz9iSRvxNrYgfD44JXV
Olhrig0jCBhAthuO6PZQGgY6B/UAB1nzZzRfj+N3/J8aGxbKfkU7V2ox9Bn/8ZLxSMaRoIPgxTR6
OZb6CXgrAhyaz08eW1SCiXBmA57C7AMgCAVNpYhlX2S8tCF2BdN0zYHwJnjqfk+Eo51ln2HDsCsw
27Mk7vbCmxIihCRRlce4iMT+0/2Zhe8k1r/QtqIuT57YQiEkdoVvjtjRpoIcKszAD8cNTC2yW3ge
0/N6JZNt/tNxcYAw5lKWG/DFylXt0XxT7VihBXpafhxy4d66ZlRKpK4bFPU7mpT5Oz/wTf6MXMIJ
y/KLxxVfByOjCq6TG5Uamf9iz+Egp/Zd0nt5bgWWWknFBcJPqzh2U/pOQfYwgzda+0PRTPwJ0aKd
kKg6qauiQUXUdbddPTBSGEhuy6tym6v/yMJHut2UfMwwmtweClLM65Ks0KsrdgF+usBikmsyJd9l
7h7naN6asXToocfo+63MfWaptarvrb5VSAQFrDVnhqyRYq9usfqRLPzzGUUEvn8jG1WVhkyTpa9r
e9cIyOyl0IDhfH1VBKFIo9+oX5/PKB6HtLfwXAF4P0SlYClL+sAtMv5S7ADXzJpf5b+F3FaXPA5+
8z1kPw2b0F4NyqcdOVSW0vgrGrGwhci0NzZfavHDSJvnm5cbZ92TPmw7LRcaH6ZOYYt9m/kZVpyj
e7kbpqqr15IjTcpSUx08kd4fMo8ROioK8EsRAmCFaFb5jJsiaE/02qGSf1BBL83eJY3DAWdthwE3
4M1C0KJWCa4E3mdSaQRM8UYbbWK4K7XiSkGMvwAXs+Cl7nkbfAPp3m3a1yyO+5+l04rdzukM4anR
Lt76nR19LdaXlbtJttgyRDiJ2UJDSLNuQdkXf50aC0DHqLyLTru4eta+89/Jyjq5WuF+oB7ah+T9
rTS9v+B9OzzXUj5ixvqVMa9Zp6OR8oNOskfPDL68TejOjnqi6EwDe8bZ761gpakcJYaGvbZudqvL
ELl1z8CHn4a/3GAwfnND5mbsj4DfxraV8U4LSSA1tQSERBQxtnr3ceaxA2Fzicw+mqJJOJAjCZEk
BOEKeEDzaziWA86nfZh/XyY6ZXyJGVywFDz5KROl+EN53KbwRmUKwLOU69uH5GbuzUxqdmxxxv+o
/4r1j+m3BtyBc71n/OEAznQFlDSha62Ks/U1g09k9Hi1mI0V3yfxA4FDUVjIoLy/DpN/uCUCYK3Z
4GLwYt8dZ1NRQSd926+mSjN0rEi7DMEWTfrFtdvJoQ32wYPh4QphbtnT+07eQNbA5Ws4GGhUJCOA
XfiN9trVfL4LxedrVtEuxxtS1wYXrfau2Xh7v0fwxo6MMVYl2suURp9LPRgc6Z0TzUkH5sUQjxfD
4aBmOjl1+Dv1EGQiJwfDimRr2wOk5yxOiWqWoJNDh1TAY3Wbj9OPDFJLovNPEb14/0NSdR3zVpHB
61puCjlM0k7bTF3JB7HOQJfaTJ5hMOUK/cw31r/Yaxx5LaO+LoFV+xCHhDOriQmTFigoU4L11xyo
mYHyzZecpnt4Z3i7YA22JyoUQKjsBlgJYYs4nw5BU6aZJa9+/oCNT95PhPCSJbXCM5wPFhsQxwd1
9/UfLf/89Q98LOjj1S7/oU1h2RHGaUOakRX0XP4cHeSJBrfBMtckbXHKY6cauyYIGSyQmD1GxiOv
3AhcJ2h/uxuFSGloldfCAdKdf5sNY3ZRzgxCfV60N9x3xVGra8cRSntaWuBs6Fv8mARv/WAY5IBs
FgjsVkdIsU9a8+xVyCrQUm9KkTHONbpHhF990soCL3xCGLFkgCYouo8OEN/knVt2zrZjYy7ih9/5
a8GwB2AgZKIngPf8HwwfXqVy7+/6CpJHWrttJMz3CahA58BhnSkAnXqJ1PUQ8s3qmKGSQoTIHQh8
BhYsXFwi8OgJE0iVyzK/zC2QaKyGOIiJjcs55T3BBsvA9X6F6DkMP+ICfeZxSkGT4F9aCCHq2SIQ
jTU7eDIcX9cR6nKQ1VsYex76u+Q6GyZbv2PYR1ue/AC0y0Lu0FK6uXORCMW1hW2lbywtSeh7Wp4F
s7syaFAm54dYCuo/+WNccENclenhstJwwE0VeMcBEkHysq0k1VvxwAC0AppKnRd3oBV6adJahn5r
cQxbvd0T0ADAWGt4xqjc6mB18jQ+ADFrGQBQHrmobRivsUkiekcIgebRe9uuaGCLguD9/z12Gr7I
IwtgTJexZ40I4e+R7zF3eVMvlISVED7u/SsdQ41abrvQSdSXG/+OgvFGl6pXLE4gpehytaPFEpwo
FVuPaCaK5zuFb+AfZAuFozfu5t6FgeeSG2JSzVNzC33uNPWwCYVJtu/WNsHgM1qhaiMgMda2bYjq
tDTKAnUF+QKQpMchEk5SHZ1MlYdHjJDzDABqDi7XglxrgzFwKbSlIaUuKnjraOW9PZ2oyf71RY4Y
rPhbRZ9MKHXAC+d8P2WiqsbkogXbd3B4oDgRVFAY07z65wo95pgE5HCD5DQ8e+STm/YrVKXggWQV
RLu7qrnoY8K8C4g75h1xs6Pct+JCgeVXNlo+D8zQVaBUSlXd4g58JBz6b0qs008K9s8VXc4zpNYc
I/9vsle1pR07NO5rfPw01dPBLKBjG6Dbf5STN6No8gA7SwwSNNuWKxHPt2HZ3by+ztMVtJanokIf
AlaVZHiEkgX2/4eHzrfA36HksoKgDXglteZ9b1xRr/WcFeQEup4uvi5oFgSkAwnfYynYQ7pSy4DI
S4yAnFXexjOsf8sHkYpw2XxautBO15onYNEURmXib0WfBh3GJhKekat6cxTgMm/czE9xhobgYNN6
8vbSjh4gKLEJUj3RGF3dE4F1lXUY1KA8W1dJ7G6xshcAATqn0QQ5z9xxr5Ii6wZlyJ8fXnU73eXC
kQqkjsAHyHFTIpbg+/8XsUU6iu4A5mwax3ZKv8U6qJedZ2/JPSaNaVauujFxmVZvhTQh98TR9TDD
1WNPWeHFZHHqFj/c2JzoN7cH4m0c/Fk58aiS5CLHZPYTsPspGig5Oo+1tYy+WtjefmtfSvutCbyu
YP3HyZwVUb8M31XpbMfPcW1xmySqDs2mSO3epNxHOK7mWOGmz5PCdAj1oU9K5bsr9kQ0D/JrFHMt
K8X4vdg+4/cK/u+jFCa9NLsC/JhL4zu2SIZwkZ4zVFo5egYOeYdDBCfElMZDez3Xug6N9WdHm4ix
ZQvIXOhRPYrsUsNZ9dD2KbZ2C+iv82BG/Lg+soKIeHsGyUov5u97Sp4kBD7lT1Vit4U116cUsMLw
nzXWKMtdnVg7IKRgGZWujnvVJlWJ4EnoP3ycLgPtMb/xTGYjWizCUrwPRvv4FeSYBLEta9ida4jC
vgIPEM36ewgq/aZYi+AueELN+dgDopcs3Ir1rb36LiCFGw4ubYNxawW7g4KYoB2rkk/vqlOb7x+U
N8o4LnFhs4Krct2KOoD5qUUqMtUyqtFwc5390ECn8RjCIVsILnGQ6FA3DK2GpdGfBL2noLYb4U/n
l2rCIiksqGiARG1syT4DvPsROsvYrm05KV5hNYFZV0Ww6+d1QIsigZzphnZOx3afFMX/l/RKdjZI
qoVNEw4GnzF66lb13nlJTbM5HWxUSlKE88NtUQxiWsxYYjhC/p+fgL7Tome3dArSXbo9iOMOMZjD
VGfQxzd2K44SktBZ5ghM3fGu6DHCDfas3s31HU8ovw1GvDR5vEr+0ftnL6SZH4P8KwFLnWF4bTEV
xrrZRlrc8kuljsAkbaz4LmLHrLbVXI9c7u8eanayWx3e18gVbdqDwcnkQUZNo/L4GL6tKzaUB4nF
t5y/s+7tKivXgCXrG3ANCXHMrSpYr4k+/LpNkCyvhVV20dmarkyZtb8ZiaYY8Mn2tVJdtguLWWs5
BURwXzq0mehHFB15iSykzXGTjKiZ/TZUrwuMQIqUisSv5CjJz8j9NOpP9lF0SJ9DSf+oVg6js0i7
pXa5KTw7GMcSgWz86DbT45b1/D4AQ1wUyZRA7czIM2U+18i9Pq2KNhaKIbzCWzq6LgSSs03mwcQ5
rg0f/xI1hnv3M9UCWsa5ZNmCGFUOBZcDc1ZrItUy+EjyK7g/eorzbpOfEbe53pYy54QzkiCeuL/r
SgST94COlFRfLR091bYajWLtko8c6Uq6rLi8Eeci4pv9ihfVnQVXFvPSWDQD0cQAqqRXHLu09T3l
D3cDJ4BScNExR9PLksEsjTEkdBnLfOAe9MataitBtCrG1flOUjTWq4pEtOc5y73lwbKAdAeKywDg
/iYj1QZPAaOna9jAvh+rNW1ooI3DVpLk8amrN9dEhzEtNdASgREVSc0KYUFY+ubNRW5vGFDTl3v0
zv2tu1UIYk98Qhe4nsZ04/kN1XUHrPWcryiuZRYfrNSOBqpLhk0zZHKGpZV69DI4Tl0OOyKsjc9D
wpPa07cr1TpjrvTcrAaERU1JRLfn7atPMJAsp62gAUBNxnUYavfrJ7kO4SbEYjBYZfjUeV/8uyNs
/3vc6Ojg3ItEYHIr0FOTzMSfsSXqMkSqA2pGnqF5hMqoLWdc6rJ3ZZ5miLylm/n1HXghAtirnKUR
4RnnocEYc2HwPA4P/wywUP1Vizxn/ZuKTPFU7IbVQqdTld6oJ3M6Y7q3i/7OGKCw/sVHjefOWRsA
PL2kyqrHndCcC3i5Vrde9BxzhOl6hJAA/b1yq93YJviW9c6axyHofnL5/p559FRnC+QzN0zSNwka
G91cRtpwYqNMVmZLd9fX1dBVZCG1Bt/vrEBeLs35zK1zsOlcNRVZFcOUTvz6a33NqgWQTn5O3OdA
bDmnF97ALtze9/7Y2n0NNC6xNj9bv1vs9hZ68Tpy/bfhHrCExbfkhv2r1xrEDB80ymObHuMYzlgm
QOEYDy4GXOo/MVz2lQFvmSHyo0w/INjQpFlm4QA8hqIsqdZOZ1VYUD9k+QoYpmdByUJjW0Y3YMru
JTSs1lXgq6gxeidjKAhWC6AOrYoP31WgTgFYg7P4PR5pYrxwi8Cy4BkM3SQQnmVYB22kju64CNmi
rk9eAu8tsv+UMPajvNAqMnj7Ubk/3in9Db+bHPcphb8YPX3/r5CxsS9PwvM1TXvnNGDNjGofT+Df
rxBn4Y5/E0FckjDzw0d21QSSDPmLus//K8OtPlLSk4bTA3w3v4hU1bS5MuPn+Ykmno6L1gCaqNwv
heaxK57Wvda4JFBuNuxI1HstJT0ZrCuHIxDjr3P4ig0dYBfmyZiFlnqjy6BXqjIRFVUbb8OF4Uyn
8QR6ZTI/q1aYRvpy6lA50/8PD0/F3jpF26rT7kFuf/QaZK1FvdMQWnYytzg+3/Q47X2NrUb0hHEF
777ozk1ONLxP0NY5S4+Ehkagfvmx2CmZzDh68ZYMx5kObemOjrjJKcPGVeRogQICeGwUns91c9Wv
5Bvj3vu6rS/P4W4bCkcdGfltjBRGEBah2aRUsK5nxfEFrRePK3YWdGYoa3i4F5YcOjhqsHNQR/FD
Hv5YRV/1eL8/7pzd3nUjtsRC46SIje1hXPqwnX0cTq/neGg2w8sORzmewsER/+mCOUhUtxQJ2Ac6
NTng0g93odj6gluusa+CqfY7zDU5TtYkv5QRPlQrikmQ6zPnXWW2nVTdh4iRef6fRlpgK/ebHT7c
8DVXcRH6sP5uB4wV9PNhNuhH4K5krUdnztCyaRE2uKaCMCl5eDIBzIshmpR/IgpMMJnE6VCHbp7r
sdh/aebQVsTl2EXXO9U3DT/ZpUStM9eq5fBIXcOvmVxeAckuy/ahITJVrDS+LV+Gt9Ry7KHGu03n
wAb6Mr7k3v5yqKilvBMrE5fgeUKV3EiU0BzM7JSg8Nv8xAnIJq7ARQDnIo21uqLsj/GHxKGcuvKp
WRxigINC/rS7BtskTg/WXRea9owyaXL2wFNm3CYmHUH/CmyMh89FxKzibp0cnuzD8M4pSBqEPHgE
IEe5vuoxinGL2KHPGATzwenmGArLexojuaoxcg8zxWB6VZBHwYyR00sX4tIU6U1bWafkRFOH98BX
qKD5R0t595v+qcU87GQQX3KL2JUuNx/wquszF5OJZpYhCu8fydrUB/KBgsVMvLrwclzF3JFdYjtX
cn0+bvpTGwZJQL2qiyM1xdxPhnwIdyH+QoNSxKsc6WCv6DfaLEfZ2RcsJn62i7Pfs24ICGOXAlcZ
+ayPsP7OhVyGjgUeaZY8q3DgrySMvq9drgV+UXEAfheX3RNaFt+pCF0nruBwg0Swpr0PZkQpz6p3
2+qIJ6jU34cFriG8W9tKRu+Azsg0qK71p9VcCwWyRJtNTBr2LKWIbyXDYXn2ItqMkAbcD/IMCOTm
MVh95eVVVk1UT/6FEpXqQZwXPFgrqYoWj0E7OXAm+M16YFLs/i1mL5UHFTxmJFpvxb6REr1zCm9H
mLXNEU4IPvXXm1aMZPQsogOZ268VPMVmPU/FrltDX/CLFpuYZtypYRwxhyybZs1kNvD0oGmosHcS
bKtlJTGWt0vlzOCI8Gyu+x4PhUifyqsORSLDCosf409HtZkEigWaDLrI9/YeZz9G/Pcp2TGIGZDZ
h9My1E6g5Lv5SRheTPylmap3tm9pdRQU8lTYAAtz8WroIxnwmeCTiYNtXIaU7PfHmhqPdPFjNt4o
vlMT/GcLEzBrEw7D69ovWtISXaZGVKHrFbzPkcGR0HHFpVjNRxFfwERLcLoeYUt+pe2CdHDRKLes
j2J1XESFqbxKI1IOUvZAHmvwDQr1XUjj2cD2WGsRHqzFfdsesroaJvNKuRK/eyjW1RGHNAd0xF3n
hZHmQ4MGvOnXNoMSSjNCWIvIJ47XfR6/XkM/s55+VnoVos1r3OF6k/9Db6/3LwodsZIFNU4pXaPr
UCdp/aQmtTXJ5GhsbQRVKj+8SMeCfvyYjkTIbDYgQ11H4vK1gWg2PWVSI40D3zTPyHiGVUfaOuke
Z+E36Adf/UGbGWCJ4hk0GAsgNXDc1V9w/LPX8one3rB1HkDMyOHRfnlvE0UHWVSPSabTbSxhhIXy
DoWORRwR4Klo781pgVA1m3mxTkiyMjX4Bh8c5FgHZ93tbJLn4xgFSyZOyJJUi1KP78JZlRy23B2o
cyqz0O/0N4ZJix7lIAog58nmumeWgJQPNnAWTUnoBiGFmlQP9NRKyVGuosVmxgc3MDo09s1FBxjZ
uT2z3kkhLUaZA+xQ7bP8Mus8w8Mxky9uSQs0yNYGpYqecMp3CNu99slTpNJauPNOAkbqsSnTqNVE
h+zNkptxpoq5tV/jR4kRQKehr+YMNmNWdFarn4AbRXV5UlFuJhvyAg2PzjQdGL57yeK+PkQAzTYN
Ulc9RWDMgTGoPMDZYkkRSNtnWLEeJhOKEF8u7P5VMbeiea99O7ef+R2jWrcOFgB43dftX2RWnW6l
hatnFNF97n1pMCOhFsMUtkhKaHuespnAILjCADmCYLWDGAcMihqO6kv1xH3u0/rUBy4ESOEy9hiB
OYp7h1QtbDPPzw5E1r0AMrW8Yn7nwM0w21OnFNbqRN4Babr5SPs0UcVgZfQRPp4xBSLOrYrj9I1M
EExh/tDQeMOH5QjSMcUIZjHG3azJb0p4o6G6ekobKqngXybI1ST02DKTBVzNMZwgYgePNCn+3DQc
YikU8Q4EPIEeiU4FGT6xDMCYz5tqyL6/5lxFPdisDG6s4cT1YAobCJ0sPSJ11nNY+/o2FRlEvlsI
qT0Uo4jIkkgauDRro4XeMneFrLxhK52oLX0qmvl5uy7oaw3TpOo6G5mbE5OXvwMb+utOZesgXDEX
DiNtyn+HiFc1q4hdCUpnR0/+weFhsaJ86eTAdiBLbt95ea9GuNxNCRNCJSeKSOO5N4O7Mlhe2Pf+
hiubJd2nuFpy7jyImssUVWlVSfi0jQE2dCcObpudNkgYrPdzCRx48dUsbhWfnMMIDOU0igdL/+6+
EK3BwTZvjOU0BvCLkMt+dAqtYeB8Nhh1IniLIT9cdcOK56KuhtlsTeUFmIoI4YFMAtNOMaUTmsrJ
rKMGX3Rtv8w7QWDORisUQVOpROfPgxsKNdHu43WnrTKxAILpep1Zrz9V6O6aTuIgW/viNdtP2mUG
EIDKNhIO2vLRMyPvYRmjzOeopOWdeYI6sfSZ0yTKswYrLHy5bU4qOoE5qeDtsYEIwjBSRfUw3I9y
lzPg1jwSy2oEs0SEaDDhsYBbe/zMjv+r86bP1QYe7CCEI/jfckuh80YBkyb5gz673OzyNK2e1w5W
7eOCO528JB5ndaGedJ/RyrVnhho3fhNLD3eGkd3oF9XmHWjyrZuwNCfNwT2ita8NR5P5D60X+WwZ
i40jchSYynDOAJU3I9yunDn0dblCz9kxkkHVPm49FEebWWgVsB/YEjKuTBrWXb9gOo0uCL9MaRpY
H+fNjMJVruBHGdAHeMl9wPZ3JZHq86vCJAk0r79u/PtQIKxtgO8HeplR383H340gPoAbkDdE2sBF
/aVbnFN1Vmi0vWuwkZQwZIxAxl6tIBRS2ccwqgZ8SRQYj2txqivIM4jPyr8WQ3ARafpGGbWEX9TT
isEZfRKl8sDql6syPyNOGAcaObztVsyDm2OHfa5SA2Nt4nFaNan6rKvtZBtj5PG+XMaqxZ8uV+rB
+U8ZE41wH9UXY2LkKFueHTVMdqO56fDM+J9DzTTU8CUClo/tBwZL/BHc0ZUpsWjRUm5oWkc48Uw5
8qCHkpvUcSQf8C9p6R68x2+/r+NC607c8z0bVsQ+AQiWg+7Xni1YHiJjVLJTFUGcm+l8LCYylsRw
LHCIx+FJwi4dMQZqZCXyvDn42VCSJYpV2bgsuKugbGdmNEbzZK5yDiv5raHAlF+5W6JiYmX1rIQo
JhdFOVZWWD3cO/V/jdYsCh1hhLL/wTqGFchsPzyaHsMjKDVEKM0M1gWSY2t3K8Utua08kjFKl40h
eLXPYVXSvazWyqYPFfoW66EV6iE8+ZGlcPX340uAwVulXcd+hLZVJqDLqU+ijCQ1pDkUSmtmHwd0
rVgj8TRRhZT48woo4/ZiM+v4aMzc3iV+ds0JBxoTYiQ8MF1UI/4r7czxoMcJOJ6XSZ3Ml81qBWKw
7n1LsEQe1kfNDl2ImivSfwY7V6wqJOIKxVU7jZ0KRRJ4DoWbhNOfZ4f6NO++hgTuuuzZzUF0btyk
2MruZPpI5KaxlaMdco/RLenfwOSXe0FcrwT839zJpEp0RVHlEGtN7u4LRFYOMPKbwXyPTwdL+7gD
I6YxZHLudSlS59u9yfbx4DU6ln9dfJQN2BBoDc4Mk4dWDBtrx1HD/dfpUta4SeLzvOnmGjroU9l0
2KomIbQ3DHsC7w/xN+iuYdvuNWDSLAWu520UTicbP0paUjxdzSMJFEcwLXTrqwPp+/0JAmIA/4jd
7P0tgluK5GjjN7Gro9dyKVwvN3xnu7lm9mT51zfazb4/JXKweE/SnBgsqzSKNh5ce8hd4OFxo3JF
2gFijx12NcPeqDw2uY06ORoo5/xc6M5QgdlWhtxB7KX5sOpiSFobjAJ78S+deiTWynmQFhsi6z19
SccLiHL+DV2/NrzdyNZLTemGdbMF60RWla1gUm8EsSNrxnfSer//SkMttFvMaSsK3KM+Qje+P72g
7PZEKAuIJhYXYx9HH88tS43jDXHkkgly/s9N7OmY42aXL5bWfR0FfSe9/C/7tfXfhqPU/IQm+Xb5
tMaVn/Uo1H/RKPaIN0xR/4y/sjKBzImnnZ+7lTMCCqXI6v3oVtYcEZ0pkyBq7HNQVbbBYEosP5D+
urEYyo5Pt2ioUtHB5G9T6ESlwcnupOS1021cro3JnPdX3KYZwFxz3U+QfMwDLlbE8+cZP9QM6+Ow
Wtgxm/WNZsePGuQ/H96lyD0FDcqtfhHPyQ5uOngO8lfAVa8vD2cu3hEmMBmm8f36esSYdi2lMbja
JBt9xAe+ZECUEXh+hd5YHNfLZSlm//B1VSNb7gL8SnDHNZq+PtIuZpZgzxuVSWb83xTOYsm/qXue
UdWxZwcB0XoCeZhORGTFM+kdWhJUWjFK8bHoPZ+AHzm/8qOf+gfLw6CA5RKUsoDAbCnkLGdm+84W
rXbZWMyzm2qMqtxlokL3gxDKRPMu7GlL6HECFGdY5oOFt7nGJI8pLhhstzYJJoicmy7u/BFLtVCN
gy7gGevJzS5pCtVebgkJrZ9X6bO3vadj7LUbb5vOxrgOHijGzRoSoRc4fdM0F2aHl0/IjE/29RWL
CzeSjOYDNpZ1D6WSeWYdA1c4Sd4WdpQYVej6M322GAHkM8U9vM+5St0YGBBEnJEjOESisLYqp/LN
Rj/23h5LjXddXTh3qC1OLBpea6WwlYsMsAgMHpVG+d/oXJ5B/1YzpC3Pr/jvfkvbk30XaB8Hr5TG
cMbnUgh+fozk3SExWJAQ9i5Kec6GgoBAqXVnQZH8fJiwt4fBVljrrPmkHja7EA8StZFpR4dSrsbu
8pMEku5xpQ0zMigIjhN6KfYCxdqamWaR8AH16k5kSXi6anc4Y3nAkh26WAHCjqaN03ajM5A73eSc
lgBn5UwJT5vI+odgepkbIMrVDQNW9sIVw0nxH0grkPI1Nku+9qt7rkdBHCpMtKwlETWMc+35USMb
CAs9RYZNfRsFJOx98UpFCxhU2PR6tHOOvfiPtQfR9ksc/6w5qJZFWXG1Dbay4FoiohozXVzh8s6Y
vwf35RMOYM6Jy7sdkfXyvgwACP3Ny5NRcot5n88cVMB/i8pNBuaB3d63LHDvoi4QX+N6Hm4xlfEt
Dwg51t4UWlSfqOLtMLIYQ4Oq5c1dn7FMKGoeLo23lSrvoLOS2XnbYEsjJReiSC4yyV0CllQn2PoO
mnw/V7aCvfegVkHBrwSkRloS7igSBdgX6tdMxuWiqER1AiqpvW8rG9b+j/QM3SgJcC0OB+4WvGaB
QOvoOrLQbmvr3RmJ6wF8Mcr/uWmPme8cwtuM+T6KIC2sSHD2640UibxOTGzQuM15yVdg1iUsqBCi
CmFfHsdi5JasU8M8P+7kyBlilE4IUOTdeC/hukkV3dv/kkU/kAQPegDBwmv/EYEfGZwudsfOepcb
F1yeQ1yLAZD1vuvhTvkp7JtOLtbnDZ+5NnJAutCMBSHpu7DuJ0x63CFz3YhEkTp9RxCuBymmXl19
O7fKVFu/Fno3FKwoSaACe9qEnhebK6dM/cEZZOBBoqOOedkclXcsVaeTYX+GjlDzwBLzbS41LY1M
vOux3zZ7RV1+cdUJfJYBM3utaCJE7qRTwdo2GYyKZ/eBQssLSg3BF6weQrfHQn9n3GhlJsLn3k8q
tu8WETIrGtoe5L9GUHdbPEcme5It3uOJRBE0x+29Upu0PA7q0sUp4PYHFGgkRZzZyRMJAsVKxuyw
AzYAA+5BhodUUdRWEo3lGUuMo6eFobJPjP24New7mx8De/CSHOckX8HDommOfv+OuDClR9zoM6St
NpX/l0TYNiX/K2PAlwE0CHs5tPSuQb2N1GKfb5cYzDBP+kOK0tN3e9p9F/6V+lxiujCyhGCzayYJ
GeQ/9gH0Jka4PqK/qkjIez1xvgIc1V3/osycUOPudlbfKBquNXf+ZvCmT/HShFicPYCEhFj0w7eC
RedvoausGS7E8jKhJJhL2LNOmbnaGTgyqn3LE7B+BkEJwspDcFwV36b+f+imjuqrHbMYmU2f85qZ
y9rzI/wMCRHeZ06wc9hRej8yfwcbipWtjKB4uK2U/UPezf73zZTlgxbNo15xJZ7y7wAkeSindx2n
5E9R4xmCbC+CogBjj1ZN67D+v8pJRLIOJdzQJmqDQZURkJjnLMnP/SrymgHM1BxRWAvx0YqRv02k
n5uYoadoFeSynEzQvimwUh0dgtb034Nn+aW20/avrDUrw/QCreZGxP60BF/GKEOY0bRZUGAxSWP/
4kjDdbaJRlL0ib0JJeSENgZvgywYbPh5C6R169umTPJ95MJrKYbzmuJQUpXvAZpooHAiHHPlBVq4
Syxtkmt9mGniNQNUWwk5e3GJeYgVxp0kKn/hnheZjEBh0zV08Z8G72i0bUz2csLqbDrSe2xAzqRl
lrLtFU1f6HOHWJFB6hjuX4C3N/ivH/DsytrAFQJ7zkMJquJX7Z+tKfJm0GmFNdwxmU0XTU1Ulg5t
EMUPBF1Qs7VKwid5/3WqyS4PGSPKhCbZ1zmfFnd0M2OF46s44/2UwZxZ64m0PosQaYMH1Aq2jExK
f/816w/ze3hDy5GU36eoPwlad4S3p4+LRtgksHG+Il+iiicjzomHIzeaOsnaOajw5HluiIvwg/VZ
ZTC33PDzhYL6LPdcTx4Od60VCx/TihOeMWAdO9CNGzub5qS78bJadOdRNjvCZ1fhqpwYCphEKZlv
adTeZ6m+bzsaQUml1dnca8CIDHA0VJuOwk7UVOF40jcE0fkjMgtY5sk8e0Clf+X5emf82WoUIY3f
z/M2Gqc272hAbfdi26RLjPj3ZkPlIr/N6hs+SfG8EpEYkrTNMIKK0f8S8NmF5waYDMYIvJUORp/F
iX8MDuSaFL0qmp4D74VB1pew5VlR4IePw6Heedz50BXB+R865IbZhwp0Asj78JpDyyeDgChPtZ2a
HZ8JTz5bJNhPVMNPVHn75+1YDwBTphsgNYyK8aeE/aXkKA62U+lHBzlE7ywlfPtCAO+VWs8p1LrI
E/sc4SiPHCseD1a0xCTk+9O2ufFBMuopEHmx4/vLyhGGNL4iyh7t5KNaR3I+jYRdbaq5+MBkT0li
ldUGS4L9jm/x3bdTtYRr6IdYFibExhZJ5YBw5XUfzGO9NrPt9BXyqW6DBtaWOUWzveDnt2HwcPTX
M8J5Fb1KZTKP4HtbhkHS9ArFg1hyEuko9sjigZnK2QPcPlK7rjEb52oDC8YL3C2f2jdhzc7ozxI0
crAurHUleoyR1gx0tm+rOp0mygLs0YiM0Ii5CPDbPU61zVSmu9fEMk4H5F5bnXCOj7ZF4txyi/Vt
Eb5JRM56Y1dmEmYByQ1qitCyu34jKQjHd+fP9+ZWiMMJQw+rC28AitW+vUjCD7YspbiCF6o1HlFM
+fD7NWbJeIgHUyhSHg/cn1ijtAwMvutoRXwDI4IW2zJWdzz5avACcjVuG6jV733GhlyeOZQfMsW4
LPcbTiVyxzBZcqamdIhH9K7Ii3f9pig1fsnYokzuj/Rx/afYC8hP6wR6W32HSIE2r+QjSXjzwa0v
py5NDT60JBZCnoIRARzU9gpQ98O5CHErUw2yF3gkIohFe2JTLvOu7uuN4l2GE/g3kQjz1xVZ/n6y
V2/oaLDhJZtdFVmQD4Anzwr3YGRDLzWiiJglBueNRdeSznXOmwQjjTb7OUKGeSeY8Hm8PN4+glBF
VyDTeo7/xeq21cSL8GpGq7xxkR7qXom/zsLOuemhwCoBzqZapStHhQ74Qr2DZE5m6hI5BoBW2SYF
98WKsytAr6y+U1ptWB+nHF6b9SN9e0As6jpw0t4YnIcQHaR4rL+jKGNHax90okhpS6oSdMqlZwNj
DHZ3fy0l0CnE0IcgrrWsb4mWJ4/lomhn9+K1MEB9Qi/ZuUHTSe45ueP2z4j69xdgjAfZ+sIXpnQA
ZpsRoog1+h3iYualxDq+jUUW3lpnj7fTPUE3A+At2leJJyIClk7nhLkt/O/i/gtpmhwxOpeaq6jZ
ro5Hfj6GEInhcUtvMr9OWg6A90HSRO4zDCZvXbIqlGO+U7fxu1iLuvy273TisQmmd8rvLjqbXJ45
Niwi+TBVl+X2AKSl9/E6YoOHhitNQxkK7DzQA0RhVXWK8KO9uiiCwHq7W95vD1D4Jup3eF51AXNa
25E4ghEXK+UwQJkK15Gzr1MH8TIr8IqA42fg/cTcEj5YNVA7sQOqyUdKkPtBkgOP5MFcfL1u/U3E
L++qm3/oc7NmvY76RzHXgXfAujxagfD6mDyEmBvcYo1LG5Ns/dlhwk/NnLGi6hA+43mdJgZQdBBj
3T0Q4k0phbvsK3ZTsjxc6ZGS7g74wqfPzJuFO1scNhf1jceyW8FcWUmNZU270o/gazSQm1Ivr+bH
Ho3EWLo7EVuneeaLvR5/BLqhQhyLmKm0dT2h4hFxltWksVYbtoZI7YHUoGt45M93qg2/Z8QlxKYe
vCKhW608AteiK1UGb2GwwSHFYw1UcECxoWNGQ0KV3gsBx0QMHuY7jP9V0e+mULDUo8ZjZjPWBP+9
BCqt9esGxht7Bo99a1TiDYI4GfZ2BRKldkHtWJKW0Xj5e1WFnwXhzvJvXV1m0e77+wJ6oGxRPK4J
3yXJYACEzyVJj6xSRzz3JmTbqz2IBb9kaC4dP/WnBQttX3Fy3adWEq8c1PNXhCia9WlA++b+37/O
Wr0tpAaq2VSZIAdr+zi4yTWdllLxzvxvmHgpSbwDnacOKbCWHVpYHaJ3naZI8BM36tk6QQK91YKM
57h5Tu8204oTxAd0qkepeo0Q2Lv246dZ4L5wSG6/NWWeEIcYay/59YNr2+G8ysv3WjK31berIKE+
zTwYnro3nD/IZyXdESn3HnqqXuXvfX2TEws0Pd+3FQnYzCOwg/D0qeWWEtrVfUawm4ZvoSmzEMO/
sAb81i8XysPXeXZJ11XAJUYAyGsTDdavAEb0yyu5g37XJ2ZNMHjWbcigBpZkritmsrp31IzVZcVC
3YmFHpEC8xdC1Pp/8R80PjiBR4t4PZV7BOh6c46LUtKdX6lh126nL5Q2af0zHsdtISMwpiCSb13g
dC0sGDLP1avdW9bte+e4wq9A5s8/osxJ9nmVLmWqwgA7VgrNwsHSekK5VP95zQKaDkif2ut6Oxi/
CheJPXXrnIUZXVN71EyacmrmZfpIMzk13zYeG64MjzUoknjtIxQYViV2WpFDRZG4c2ndY37QIiqv
SzikDuA7asxdHLe+pURkot5tqj4Z0gWkfAqrYXxXfZXEA9CBtgoAxXR2fkEVohCBjuTNS/fsr8qt
eGboVLfhqpAQfrHrn2JN6kM0MP7xCd1kSkrouDNqQUCK2AuFfEyKHD5mjK+rc+6eLbSPrzHW/DIr
In+KOJAQ/MH0kCZR//dHuu08oj1lDxYg7CQf+ffM0OS8QeiOkmP4UXMPuLm52ERXah40kOzYXdSM
smh2ohLIWTABRYyAT1SqBqytQZE9cVaJYPgnevrhKDTUbiOZnAZulPWDgyRc9XudgoVlF/TLcbIC
ecdGXNuZl+bg94Za1RLOyZ+EW2okKjbAvhtkPMccyInxnQyi3bCAWmFRZqydpXsH9tVpARuVqlLQ
F0la0b0ffklw0TgXzlVy3k1LmpuUIx5K9OA/E6/ZlGuSYabDLyNJY9l5KKdJfaCaVGgL+wXxbs3f
LsS2xNNiL8zgQCp+0zvdFyaulVk0qJJN27KMfebwKM14VSNXUkgW8Vh37hHPIwgvYfP6NjbeUOsF
BsupjddHSwPnR7dYJoqkCuPNZMgrJdNE++rFSxIlvh4QzQn7zGe102LqAIYKT3N2yU6gmHXqpUM8
rfXIedUznCf2H734itCcaDjhLivKAPZqCfA39mUOHDBUETj1UYIOlMIkySf5+zZTM1cQ9ojrbLib
scN0STuavxVFwVnnSsNfFpaJRTSxfEWu81yeqONQeJkUC9bf8BwKdmQ8wG1QSOpDSvBuAJeHdUJb
hqciPpH6BV8ApqLsdUuwvrusz/Ddv4TIX2xlEW4i2GaBC9R6MjqRfBwRKlzuYrmKqQ3UGS6YmwGu
xc7Z++M2Vssjp4TfhnNUPmwN6yS71e9xdQ4BEBpVdFZ6PfRhvQ2IBR/KebxUPfHzCSWNzrqmcN4D
SzEUjR0K10HwSeZee4MbDXuI5Vc7gHYzmj3N8YTyEsDF0PWyJn/CtRreo5N8bHB7BDDW96RXUgEd
U2AmflMqasu7rTl9IIEgO95xPfxdQnWPkuQUxUoaJkBSJMDp6njgFK5b2rFupPGAhiMw/6ZZcB7X
BUALZYr4fN5vtpSL7xHW/3lKIiWw5/HHNf3eo5a36dIcIi7JuaGjRGmw3BuKngkvxVyG0XJ6DbdM
NwGn8dEN4oXmcI7HkAW5cEeVUoGsPcZtjiZydwbx21GdV/e/eNavMuh98GaPl4XnjwFt/Id+iyoO
GOKc/nrBZZgfQT/QBJ4OgRRj3VbPuoW03Ci7bTq0/zEIzlh0G1aV/CtsqUfjxSUoXMx5Pi4KoJct
a0rPb3DgpKoKlfZ6B4q1oLUefOl01xeoVpv2KXib4AZqLcBG5gozGgJolmqUbYe3NVuG3v/UIjJa
PkasLyZ4vWLguE5eTuoGTUtW3w6dzJdKpgRasiWWtRSnmJbJTPtLZTNTvnI0AcnBkImCfCg9e5fd
Q15xAT5YUDTbT8ohgzQqAOeUgHrHV4MYg1JmsWgIDobMUl5T61kx+80UPho2MS8rpoqTg+pwKnw/
tx0e1DQ7b2ro34CaGsZ/dSpeD5Nv7laiHHzJgbWT1MvemG9AhBVfgq70sxNDpElzlHrnlJeqm+mv
SQEGMfLzChT/Z4cONJuJG4q7YU+J15TGQTlWitg4NasaNqlmj1z6rCO/EGRW4f4V5e+KfezpT7UV
FeFAqNXPMKOJOHnFmBTZ6zSHmYioWY5XIitf29IDhGej8eHnfXJrsG0/ScvfMGcjeh9gl4ncrrQC
Qr/g/ASlO593f/yMzQ+1nilEPaM+9yRA+Trjio93IuaZGi4WlyxcE5fCU+5CX4cRucsccGR2IYjh
U/L3v/jzpO36PsF36ZmJCNLRdM5mtIdv8sBvHAdhUDsmeiEaImqKtPPRV3rFTtAsisSOrPAkvrjZ
3xFj15BYM/9gAGZGa8Vfyt9VCcVnQUCCwEy2hYNQ/2bQfiRyy8R2vU8GISy0XTrJaLP44R450IPi
TgwZYcpkNWJi/dpKiToBRpVHn9GIYtu6Fjq3WBp/FohvwOn3pMSSDWXmDI7tFUi//eDWjwBr+nTi
k5kAwx+fXNE++gGAqwQcgFZvsmdY0bbmtYg75b6seWDicQh3oPEPmis9rKM/+eFFv6WlIsKGmEhG
swWfMmRsfLxAtqdLRJONnKIJY6DnUddOQpbtZ+b11c2M/s4v1oKh5rPnUJyS4vXeYXCecrHqXIfp
NzYDEhnfVzd7YBj4MncGb2Q7y/AocY04peBG3rFFg19o+QuAZWjqgD3pLcxsurd3n03IARJsCI8W
738gj69Fa2N/9V8SSojFec5PV4wIjUKHAm1RAJmaklSgoTzAu5AMsRQp4986zgfirQiMyDvI7e7b
L5OBKqlVlVUrOTRZAaoCJC/G6vuGzusRwY4WRSfnr8UUt6UykmKYgLPl2il4kRycl7Jwv++gT2yE
o19VWx8E+WurcjIsCkg3WG3cfyVVhreYcZhP9qcPBJEbmaMFVhP0WrSgafl/sXDr+Z5K7gPdIfbt
ZwH/IRn+oKRpWJ1Af+LVbkO+ZKuImJJtp822qD7oNybON5McmfmjKnR0jECGNEUa382O0Uw0K/ey
bKb/3+BoyKL4A03gE0XZJFeXrXWGW+YrRB9jKx5yf9ltK06IjE2u+f+dzNMwVXDAKi/0F9gi2fpP
voMZPniJH1hFihcgVQBOBE53ioK79ebsxnw8adifu2q9wwzdhD8siQCiuAubd0nS2xZxtAD35La7
O/PfaF1dcS7cynf23DHHIgf4kSACIVaCchMyRnhs6lyEIPDdoB4+n2m/7wTpGCJg3orDbtHZqBmo
bhz6vb0kyREVnVyR/JQuPTuWBo65AY/h72v/0oSgqrd69s6ZJOIlyIsxTwUCADPkh5CsyomRnq1K
/bd40lQ2qd4L8NYGIi47LTHtJ/bcWYHbeaij8gZwxhyp/fsi0UaDdEWa2CHtSGo1fKqbNvA3w7IM
fdQI3p0+7dP0mXpcVQKn6zKmpAKvDSxvYnrmEBwGI51kwyjkWcDvSyWWoZ0sMDDCLFVNImXNvGgf
vbsH85wrTzVUQhDQHL5raLD88AZE5nZPFC0UopCTmbuMU9mCIcua69gfG5AVPLB8dFnFM2ApZNwZ
2uYBe0sAhMUXTZkGKfzlm+i5yT2Ml6F20AipNcSxmOwnPnR+bqip0x12ZiFDsx1Uyi0UFFXaw0Aj
bSxto9ZzBxPTMKIUAAmvgGBQuCVbZQEHxCpIaRGNP2NKNbmXyo21MoWqzINVB13Yt10cO6e0fJfK
EWRP8WkUFGBCDmUxp8bXuhyjRWiZCN2ChDQim/LvyVcRP+deVCNMXwoFMctAPCXNI+BYLd4hVNg+
+xF0WVnRLAWGQWnHYyTTGGf0RJ1w1/noCYbP0xKrbBGqjqrxl+eJ6xnheJzyEdZty+fUxmmw362c
4YWVAW/swOXM0Dj8aFkd3scgtbSIaemAUAv8aOqVpqLPOxUVkZ2tnwK5mrvNOrjFFpfbnevWt7Dr
CuVekG3TLPpMjjhxKwTzfpBnpzkUN4V5ma0UGwUNiy4vlLMqYKrL+HpnOFD5/Pc8aDZ/zhh2npfR
elq7W0Tz+FiYh1aF9tzJ/L90gpouCbVREuoMhgaYUUpacgizzLfRs7LMNpZC0C5hct35xZJXtWnz
9+xHUKWWQ3x8wmLpCPsMmfXs4OtKh+KgFMpbl0VEVszCYXiS1WYBHhcVN28/mGocKLiHvPTjJRSE
yeQOp81VbhDckcpRf36v1Y62JqWruNJuoOz5RK3xXxxnOc/98H3uf/kcBWdYW+dakSnJflidVR+W
BNEHS0zXRBWMnfWJHcu9briXBUIhAiwv05qxz5WKQfGQmflLzYoYs99VyhwZN+JIPkCkIezdCtiL
lfsG4DWUfpscQcrp7APtdxSdCNvrXtJLf77Ez12X9MEc9h3j/sD/tq5Bh18Jz47AhfHXmywDpJb0
dXCrmc08vP7YTBMWG+EZ2NxHSUVKwxlRBXwR2Hpjm2cyPeyWuoCDInYmAjWYosWvasCYoFYS7bAg
7SBttrVHE3ypsgMx+wmfo/B7C/GjcSVLttYHIJEsV1sYtBVdKNVDnz/7vKe+rss8ZRtaftLvbqZC
JWuMOl77/QvMo9+p8Ghy2dwWQlK0uqTVka0SFQelsgInEHeJm+zbxlPHAuPk67pQFOyy3LTJY6nK
6iSxLy5kno7fDMD9eBh5kLP11DyItjNymeBvINvMPY3kX04dbFa3FKbT1BN9b1stmH8xxNJmEf7Y
DPoL7wKeUHgLDsciSnwkwkMJDvJoiyRXdTQZMhd7hQcQ8hak0ZmvIFmdIdXK5NWexRcDWF0P2riv
J212d1wYCnQW1CgXlnvwI61Pwj6/w+fXWCX10F7h3D5wuVIO9XkhXM8JtnJrkGaH46K1PvQa8UOM
IujyuBJ0PRqEe1HJZeqf54ACg7eSB6H1lMV+Fd8w/2KadqKrVDEQseSc94uY4GDtAVmTgGDir97y
IzapS7bpyoUENmNrp0F10jr7HLjXTe8QLYSWi3hU4QLADJjLICuC+JeS6oRSNDK0+SEBQDT/Pz+t
ly50EeQZXbFTwvUJw3hz7ZZFNdp1KsCKXhQCQf88+gbJ9I41Z3ZkidpGXyCr6lyc+lI0n72F4Nws
8+kdDjvKGfmT76GLlhNWNxeipgONRsj1TL7P+7G/vWsDuhKC0v+u/1XVUOvOpCibhzYpbFb5ybps
tHPuiE25MD8w1lVk75tVa1V08w86Y5CI4yuIiIE6tCLuHUlwsKbEcBpbdoj92/YtthnmDMAtHRiV
Mjm4LRW18e6N9d1pSSfI6I6dQM8PIjygxZ3kAYJiqxtJurFWzU9LdgVbMU2jF56yRuKXDIp3k6Q6
hCI7nIsKQMSdAET27imYo474Vr+poVb3cfh5li9pzR3cZ1fEa52qySGilVstczn7vDQCy5aaV5Cw
WmEOGiw6HnJBgaU6WXxDMZeJtrOz+LNVk2ogkVhty/67XROWyCX/UEJ+XikKd1xBUjOeDS60zFQB
oVeOSMtFQeViiVEzEhaqeWmEKlyzTulBkvOz+u+womt++i1zrFx0C87/xKNmJ0Zkbb2hWKzjJxsU
bmzNDcqnpnL4s/G6z2OEC04kBvVGuvVrAheFIORV7yyizOu2dG2rlb11IK43Uoc3kozfXQ4sHLmB
oEN6GEYGR53N7FgbYf2fFMwuYyi17xWaxHPQ7ABuhIVPT2b/xGjjVSwWDRhpZDT2ha02KAWOP+do
FdI0rmMARmsgjyw9tvpDwck3IAx8YKKj6lj8U4xcyq1h2dPjp22h7UaW9gdrqTZoRJQvqCx9tKSj
Dmvxe/EEQ2NznLjiJENOfg0p/hYxBNv8EndkBC88/WPS5Vl/5dPM8U4/f6aB9tBG7ugSEGwAjmya
8cEWgm39nF+yCYuYj5efm/jUvcXd70ycRT+6iBIDnfIQ1eTxCB4mxw4i6zzdGBOIWhopGZM4vghz
0wPPpfFl2YK6DuXN4Xfr+xh317x/lF0xagLIRAIJIK0AqLieHsyQuWpyk/g/R+fYGBmIX9dk1pMe
JtvXuloQC3BcnW/yPgZugXKN0mwh7YoCQttxMRL1rdsxKM3A2GdPObQOj75WP5JHDb+AIPZzAgnF
VkMqAsqwnuUrBRMGUknPBR9xadS25C+tlZB4ukAQgCYuNFLI37kJFHdZcSX3FY4nc8mt00qZiC8k
DGW1Qa6MyLxpxMtl+XKzuSi4322TRnmG5RwcZnuxGdluefweSMdCyX6FG3uC8d8MAZdr25SFBtFA
W0u4xTZ7R8DFdJFGnQzFcmKdi0dJTGJulsREsOLO5Yp4qwhR20Qc+aAfE1XEgXMxRIC5827K3AlK
Zz/FlOVSXKLtQ62k1LijR29veVbbVY/m0mJtbq2g7LD7yjYQcLE1blmjVjrkrPzsUUH9APdz8cmc
MY+zhKk1wtORaj9axMyNBRAfJ1rxzkA8bXpXt0BAiOVDEUop9uAanRZFn+kLnxHsyS13amO7DzTc
sC8Ehv2pzGxP0uELZaqmdSHe4bV+ux+VMg8GY4I/rgk32pYPY3Ht8XKU5sVWI6au4BIhzlAK8ewB
A5HX4HaCQyrCCj3S1532dphi71y3g6xltl3xYmIPV2vWF4wlcYaGKSxEWgW9j5TQ3qnKlK7v8fA6
/yNRltHyNfgBesxg2AY7YvQ8lao+cgf4/DrmnNz7MO1bhTmNuRk/fBQrp1D5NwYEuk3sG6iKvE/+
9x9j7GIIJ8vctGLVLJLiQigD5Oi6wli00ogQAB3n2v3ZaoYIgpBaCC31FMyLY0B94XQ4mNEwPieP
BAMkhN7247eVJgrHdS1is0hebfeW4EPzK/pgcanVMaOpLgTlJRXZ8OSv7lrcwMVekq+qH2FYWNyn
gWaf9KNxFDob+u9Ap+ch/zj6aI5+pLWsV4FMFSuE3A6GGjdtwiYr+bcoyyCitttYNczfKUH13ayn
uxo0a5cUs9iaj77WFYUBTJ8PnNAEAUD0URwqbJgRTUzTjuNc30z85KeNd9dTWvJ/0ms8vNSen4I7
cYiEOPbIM8LwPYvppXFjCwhDkb+arNxVucQ83g1P8hiaH0fLeMAmGzwg1XPW6Xfn2ukXXFVi26QU
PJOZ82ZMJGKYQKao3SNojqKx4ToDqGDJO1ZgkH2i/7t7Vjtojf6l6bAMOnTyBMpAmO7TWFEfhk6A
y4jyj/Inv1+CuxZIWmncQ3hk/a75KTB2HeYkEOGt3VP1o7cK9PoeRiraNuh5KNkzeH5FMJys3nMR
hU27WmseMQRF9lU+cqc2jZg2pSHuDBa+dBt5Y6J8LY0MbuYiIedbRXHrGUlblB/7apzxv+9q0sgt
G9+1L4Trh4RKECFa2P/OEzoobxsthqM4pyCJvXF1rWtZ3DAoYS6Ql3Wr0pQmrqQbxdy1kiK7ovLG
PqkEtLNWvHM5DjpPXW71yv5ZemY3r03KJscHCe7qtKWPQs6/mxRaqFKTAukDBKKFOo/7pEeDjTzr
u9uo1tFXtD2EiOVVXxPE4GAtB09THi0Orayk98alx2tYAxJfzPFaizoY+kECpljtrTuKzL04nRyK
SdAZxyQdr7Y5Z9Z8bXMANEmO1ddAQlblniac3m9q3GwLsAGlEeIxmWXzdYe4+ZsL1BUQYgG2U5Bu
+aw9W852Ne8XXWZQ+zo+x+7asI6j4/pzNBqzq9SDM+1Whh+GjqB4jzZYVc02x7x3HJtovVEo0ZpA
1npavcD8uBUWCNL5tmxZH8ekp+RIMY3oZPxnb/yKCQR2z/Vt32i/C6tbLssMKWsO6NottDTHOszg
7st1i8UI5llwLIgfcDpnqzNidAb4NOmuM2Hqg+j5wTBVhSdoLtEiDMjnH3TbByUhi+nlukADGUA5
AMjLJjcjZHc1xrHV0qB3UIqVqCtkTHzC2fZ5SB68VMwI7I1ZoCV0h6J7lB9aVIAs+6y96Nrp9qQR
ILTnWmnoxeQuD8kkSlyBaYAA1R945CeKfmOz0TiNJXf/aowiyront/s6s5aaT4JE6iwKMwyD0kpw
Y62jeTihObmr5Atxuvvq8J8vW8XmyRyWH14PlUWZ/xHVmD+mcnUAIowA1AEyR3q8G13Se5NTSszz
k2n9NlwZzbeucmVcJJLt+WODefF7cSLU2mM4YZC2WrybRmx7VwECImG4nLzw4yuY0IxuiHSyy711
pvJ8SqFaF2q15cRk4aHTx0uWl6IEwYBkbSOxHaeOkkHQMBGOLIOQ0iTp9RzH+gSfU09WSxgwG53w
BuMM7siHxV3b8K7UnW6UMyTzi+AzSES9CC2MsJw+I55s28Mv+LaxzLYS2Na+8jk4j6t/rYIPz9Zy
DjGz5rtd75Av+ZbTJJtMODJjjXZWRhp3j126ARDdwh3gzfcYYCc1PkEfXMu3KxuGf8QjtR6QJwx0
4JlgKGepmXUe/o0/eBUYKoEmXzUodt7bKOe6MVaw5lS237DYvlYFqm2GMCzSxGM2GjHVhs301z7/
JzgB1dTO3DvfeNWpIinXtMITGoyhx2Or2P10KLRGURQ8g1WmpEhWWGv4/9YYJ2+1eZwpTVtjCTfk
vZmg7+mRPTMyc96Kbs3T5Ac4PoEHLvL2qZiYkE1C0vObObT6aM+xvOZ3kD2xwomrZ1j5Ur9NBX9h
vxws9+T9ZpwdtAeqLOlelmjDnbCB3juGp5hP2OhuETmSeJrlkINHOhu4RA6PZAzhz8XbV42pGn7l
IHWzlnsaTqFrzGkZQxTt9V3/vmXk7qeCqQU3iZ97z9jXRv0xAP6UBxO0byMjw3Qn6VYCbLwO/xOv
LP0ad/CxvjSRq23MZ102teosb7+oGfdlF4kdPeqTQhyoHrj7XT213hocVGTs3CayoxeBB2ZXG572
11I7J5e806QTyp+gB0PD10D8ZwisF3XaZbHm1tXWoT2HJu32UosszUThXNEbuwgDA6JrhiBGZ6xm
HfigRcnmIt9Ztg6XWowT+Uiosf0wz6y/RDa4nEsNS5Qz36k+vrp5FUf8+6Lt1DzvfgqKb4bJX8Iv
idYDs89Xqmk2cE5cxTkADks+eKhdg2b5XGIEKceYAE4oV7/gYWlB49+kMw1ComIOqvbi2cMFs7uy
jzqi16Gib4kKoa+vGsSesJ5lJuLNNVdTf3NYuV3B6jaxCdd6VG+YWfD0fELV8gVePk5SFu2nJjn6
QeZrt4KlyF99Vsk4o4g4RM//9ckOLMqEdvnOyH6d4XChBe6JUho6+zHJEwV3TBmQJKIKRk/QHKaZ
+fRd9QX9xNlVa/l7f0tNzVedYqg8GuJ/1+GaPLRet1Hj1gm1yKVhoCq6IKhxkqP2Fr7QJ6PjVV1k
oGa+yPdZtSVpa4Cio0mfotV/Zn9J7grfH1tkrcETwqHJuXZDNNj2ErwxRFnr8x7ESaiwCmPoEWhy
Gdt+/fCaqIkF0ziBS+1gbhfD1znx4jdyucJatmdKVR6x/0ZRb5artcTvHG1MOtcmS8gJn9hcbVtd
GEPGi9dlzsSO/xpiDHT+Ps8dHeGLlFMmi0iUKLRhanL0zuNGyXqJ6DF6wDijayWj7JC3y4Chp2Vm
tjryCYp1sEHWt0D2bIJaONNjztxH/wlCiMrPPEDo2wYoh4zxE2chHc42lgIBX4dw7YOyzMF5DOQ+
yUsxbkafGUUsvYb68R3bweDa6ylCzVGV1DGTFgZ5eyLSUPuVre/Xjz9q6i2//Me29MsPgwGhz75c
rjaVAWj1Yegxmee4yXl55DsoD+pUe1hxXvUIGXq1Fjh8Ih2u7ZejLUC5RUF8IyK9WuG/1AnJBdhI
HfNZo0awXbyGgFnvmWN91kiFG1Vl6e8dw8VeWrF9Wk2fcn27MqKYTFlqyLcZz4Wv8g//hh4pgFek
2GSt3+pH0TNn34DiS+9CyB2r0Fv6gMRc3Ni5EkVPQoxm2n5Okjr8++o3fXpLlGRRYb1dmM+SZpVi
JuMGMqq2DsGbyqxE8AcWZI9XEpiQCKLwdRMy8Dx9wQ82XuA3I+AEiISWUPqOEQMDy/OlDDapFERN
YSa4dtiH3zHjhtSwu1+iQ2b/lFCLyYlafo0pVLB98xuFU7SCuLDmQUjTB2saVdUtE+SAOjOCOjHp
+JccdL2CwuFUi9Gw76xzL8G/JlXvFXmD9FjRj1QFbT62UdWEvAObAGLMoLG9TlPe5h7z/6VM4aYP
xhzT0OlREhQzT30Tsjw+wBuR1vtq6kcvpkY5W9itBTZNBpQ5xuTpYW7pT/BlOlI5e4Xot57y+Iki
5gl+S73NqRXqn25FFWLiy4TW3YY6xYhBY9OwfzcW1cac6sB2nytEDCEdz078LI661NfhKGFcZ7lU
PjlUh7w9w5yvcuBPMbVjtYcJpnoOULpa5l6lBsM+r7sInC3zVuxjrKMr4uF725mEOkiPrAadcz9H
OjLuq4Zm+QjvpD7jx+4S90yuVHcovlfMFWqON4AJrAXWJ7YwCTZDG/GlX4TlYskbLf80c37NATfo
2YH0+wndv3+eGTEb8I3I2DVtj5CVkbvse/IK1NDvUeQD4NfA235guwAdr5EcCOSf3y2JjA85p6C/
8d9wHH+VSZN4qeyNhvsMaV+jBHBbfJhJh+OokjeI8YbwZZIeqAy43G2Up6OrifrKKNhYX492UOoI
ZSMfT6JjnuklPs7uRAz4zOZlbXsPM5R1MlxbsifVJAqVUkmKrJUQGCTZXFItGa0KzkRLwur2FaRI
fdVPwkliRz2utHlUDTzpyG/xDN2SVtguTfaGfki/BJ5OFEkPahFWgVNdDhtV4f1j6xFFSXpSd2CY
6w4QAFNPgngqR2nAazu+aHuUZlxh3mDIGct+Fsne7riiFkrE2TE3SPyg3RayLA9oBOGxXs0fBldd
G28EzhyMehhFS1PJDmR3VGxmducSpQzrDRUB9Wab+aBlLADCRTzXVUtNPoR0Hr44sT/gJLXGid4A
ZqhDva18q7QjNETBRwQ4q44yIzrIMov5HhW7pMlW0bNoz6y+jaRmNuZaEwXtWo+YDTesDgbnof0i
3c9q1ibfS8m8CTH2u751XZ44mHwTQA+HXuLPoyq41c77EXoKuFk9h+1QmK3xfeFwe3aKkLOI/3zq
riPkc3dCwPv7zB90ZBBelzup181n7vWQPZqi1ExTodi+bfTKOkiop0kTSTxnd03TBydw9mdIjBJ8
ChCmNx7AaT/mzcDrjd+TE1VeIfDTe5aGBmmUbF0db1dIP/s/vZ16nm5wIKjc9USd5mRQA817mE2f
+pILgrqSmKks9GLQbgq2k6M+4EYBXy5OY/h6GKLLtjZgfC3aAjb4ahRI8q3BaY60bjwnVZP4r6cZ
xP1yCgK8Dak57nMqCTA6P+W/3Dl0i0RXIsbWCca3bG3bEiZ4tKqgUPE/V11HOHWQSYVO2bpMSrGg
9ONkROtk9NTjzoqtTSdCkY2VVM06TKi+yi4kq7Q6jqQMuqXPsHB4vtKMylp1FFNKX+C634mPYgDG
k/h1Q2YbkjHNZv/qhHOH3pKUkeXVcDlIZyfLk0Ns7kSrvkn5oLulSwUCNsr2h4jdFVpPKvjJGzmY
5QDxM4tzV9PRNQqM4PV90fudLqHQd91OsSzb+j8+OVXTIjd0MkHcWPYKM8TA1GfKrh1Jr7jNPYVU
p3/+N1PiONNXERsXnlL6Afum3G3bXvDGTE/19yzdRCMDyZKQnYseqtYRoYx66QvASJUrKV56CPVi
Rv/qURJwGQRar3zBIjcFoSsVa5SkLQoT1mIbrxi2ewoqwuGTf1t2XwFuRUT7LBYESD2OIRwDRRv0
vUyS0DNtd23IqUf6CObPhneXphT3XXuJETW29J75XxJ7qxK+c8OWxOmeX75ff5Ge+6dpKOXzWhS8
XBaFjwTyJZ1TtL6hkMr1ETJ4xfZ/UPKjDAkc9WDiqbzvCmLnhCwLB1KnJVNNleYU1prv6eJrutiD
JxoWMtCrI5oPzcHt86ejP6GqtNnJfb2eNhJmf3XUciYYhUf1ihruUvqTAcz2wyuHIjO3xx7apsZN
wmkdH37eUvj+CsavZZyhI5H3ya9j4ImnQ0q5JHs7UR4weyW/E9tKBP6OqRUvRcid3Ffnrg16/9Hj
ByWC58SYoeg1TFfHOqUXAnjj3q3ad1zURLT9ktlQ30tTT00UmNyqPyW5KrJQIVozAfgfkvnxnvgp
+deNZWRuwDiSSidyhju7qLERddUzJzMPLoHAh1+B3p3R9R1fm2PtmMRRMMBtJ+rPOxUknBVzn2ga
OHbHmsOm2f9JMTOKur8pWsoz+iKfrLrAljDbRpo7NuFt6Qh+VbD3bbeGUlDRe+aQguDp66I1y86r
at7/92xEEm/uCCc2qe7xvxOqom1+jPL3dA0pD2SOBhzV5KYiNqFs+QVkyjKW1Q6zcXiBJ/r2np3Q
AOj3D3EfNKijqMD+5zgvZggrGsr0Hs1Gi3Af6UeLeKUu81OdQ1AX3yi+b8gR7heSy+Abp8ZnLlk6
RFT0WX0TM3C+UYP9Mg87QMyg6ML0psjVmDP/9h+PzxFF3amQT0HAkYiizrxwjecj8BdMtYMfgpQt
ccUY29SqCTC0BmzwRiEt6RmtulcJVFogOmhjZZ4XSbOvj1qsGB6gLBKLK6W43gUt5Pb3Ym3ePdlD
EsSuPb9gEVRWBOjogyfnikXshPTYzk4GzdN5f+pmAresNSrla8fSfqmLnKW2xQejXwyQphBpRNqG
KkWE5uvwenvJ7qxQ6GhwKyT7h4uKZWAvpL4PTKqJh0Sfkp4Fi+JBFcth69MqKU3F6z7d7J4PsocT
HwmaHEUuvgjcljAg7tlw4GbQs+8ngicwsosGqiyRkd3iUVzB7cOANjTHQPg8M7i9nckZ8qzOswdy
fOBSwyxG7dd9nLXfuHFQL2ZgQ2tmxqlEe0ihE+Ovd5ZtPJAbYIHtjHRwh6t3XjfjnYgPwHlwKnQb
e8WMes8L9m+zTarL1p7ASOvSlkRCT0ocHaiZx22FsVv1euGtd8tV7WRKVFagLemOGvofoWoEi3A1
8VsVUj3oJnuyfYd7PvgWLnK8hfs66cWVaPv+KZksFPMqg/EFBG/lOEDqhIcRWfBHv3g06ReqS+DQ
2iT/vFJc4iWfvCQx2uCWzucHeE5KRMeKe5ZbWmjiw8pYcul1uvWfMkSNKv48Ku3Z+Nbk0PZNQU4N
iTkJ1pU8hiHfe6Ws+I7PYCXlN6KE7s7DSIW7i+ujMN1s4R89cFt7ikhlyzAUU86ltFx4HZTIieOh
9cNcbuptJ9VTXP8+7nLCzV4XlMESuBG7YaexV3xsrBkUEiTC9hJjVyprBj95aHO+4fxSoYXJ0Al4
8chk3b5EK+FowZSmeT+OI0/h+IksZhabTqE4voicBIbc7O2VaD4VOUx3ZJwiKsa9eWC4f458ZlU+
TwBeuV4vYOj15FFwIBQY7eRbu9Q7C7Fkwec8X3GCBxIvZ8E61IIu8L1g0bN5c1znZeYC/g+5gNJY
jMZkWc1ONlFYdDwGt3B/R2IAQuHUZqhxyaweaTb8qSx8paokXAN9Fq/DcxpOYYMNTy8/S31xpHTb
AiIYECv8QTjwv/xqMTK1JsQ2HNFVULhjixw2jbOsKe2/MF0bm4lgXTZU81GZLL4ex2ezncOH/jQP
FhPfwxkDizcIalbUem3n3bUKP9yVmOgbC+uIwJGZxzTy2KEHtERBIUvcuiG0L9VfbRmTXNmOlWsV
Q53mgHCVR9SbcLVazpR1DKS7N90SgEeQj/51Lmvoy8qLD5e1TTP9CZCIuytJdoekrF8P/PJAcDkx
ZWx62JYRsSsT4OOCGMtn19uYfLtE9rBGzMrH2PSPgtezYvt26PifVeIU1geNM+yfLpys5nswT3nh
gKu+c0Ktvsbzmo12ZsSpyUOLpktsJxouYXS0TnNwT/28YaBzl9zM51KY57fmc2QHONhQzTwrd3zG
lHu2WuVW+MHb3INlYF+IJc8w64FcbQQRkePIJj0r1fy0njevamTigghsetc4US4uWxX70WY4Bem1
vMoUw/jHWG3bL0ZjY+azKmm1VaqpDztz96QFiP0mQs8Qq4pv72AWArTTISHXdCkfxiXvpqXoBwSL
k4UyUWf/oo9GWmc4tdz8kGW7Or8VosB8PH6LaH+G80xp0QGOtwUH/Rf2+5sb9FbXkZt1It/4ZHyw
dtTn/0I47I+x9vpHsE3Sj7wp+IGUsEL8K85UG7H+wLNZBJH061K11bImfzY88ugFq94HqjyHQQKN
hEGiHFXlOeQYb+U+O/FxmN/Nb6MbMgWOJMU7zkIzNULXBrezkc1871n3PKFe2zbAvmu8dA5Nzc3Q
u/nsO5RcpKu/1runbz7f4vKNh844mEAG90wyPKQc3P2BDudBEUcy8BlDgT3BPtHC3T7BZVE1ZaRl
Hc4Nmwzj2ez4PxD5NRnh0ulP9pgjOkX2Qm34OZFdoekyZcXZ7aUDTtGAwiUPbeUtlnrpidLiIoiz
jBYLB7ybNrEHg6b+nRko0RXLgtEYLBZy0vw+AmjOEmmCqZhHiAN/HssIN4vpM2HKJV0IZfzYnj2f
jhoc1rAH6nYdzdnzxDOGhRhx+3jclmU5kBhkwMGDVfLs4AZWWfbOIWDgWPS1eSe1ZXlzNrKbFXxC
ltx3cAPYCfH+g5+ca5RkYkJYIBCiFV0ehcUZ1V6J9epSeTxHZzJJq3/AXKyARR1vmx01k6MMR/Wz
OsTRX3woYI2eLhjhb3HjVB32zL3Ri0jdHd73NMx/M8c+y8kM+wpGJ4V1YrOnTBEomDGoktJFhiRM
8m9baxj2lnc6kNRmyWWa2IX/XuycZGF+S3Dsue1uHc7l0Utp1ituvadP58A5Ih/CgCAyndQCMRfA
dmfSu1kkX+7RngK2i13XUz1seLnJGnfClWTfxoCG7JpJLhFn1D6o+H4hcJTZov79eDFLB2zQFXef
kMIz4jgtu193dpdmUKoPlXpOQSkaIK1A7M1lXC9syi1cbiUXlEkc2HSHkMzurdSDI+vYplKWao31
kxozovQciv+T6BWiVhZSQhNH0cHQ8DzrfbQq+fwZulQvKEjX4FfaLcse0OK6MiVt33wVaqhh1w8D
8p1s8jocLYK+ZPaSFaC9NS0qTblcCz9fnxJ2NJ6YNH2cnupjwNcNqMxbngdkZG2BLG77yNbAl9PK
69YvFx1CrQpyPQJPqBpVTIOXwt9m1Hah4wT/XxhmsVuNHEbZwmNA9hBD3fzxscMGBDNH+RCNI6Lm
0g1fRxdYX99KEPYpk3gKGRRo2Xb/ylF7YuWUpUucaH+AQAXVFMfXP+JlgClG0U23v1cPsEzVYLUa
5eaB5/Tkzn/UQJZ5/DqexpgxkDZgFZciYE9ELMikjzxXVp/VYYhWX/qHRgs6nHxeSzq/NuOIw7RM
iLIoBjgeWqUZhOYeWRxsqLUwRyl79yW/LHAsYcGfRs5CDtFmnVkrKJDniSb+hZe2SrqFC7tMxyvI
Yaig7/UNDOmKYv/GFWL4gcpfxr4chDzXxNmfnE75ULSZ7IgBJyvTB3pll58E55awnhEzOtLId/Mu
8J9Hnfbsc9s+NMPIkJfaYtX5l88+NyBxg8AmyCgKbe7XF6PoM8hKEJiOtNYSc0SCQZpY3ozvlEd+
O4NqU6h8mLNl1Sx+gpvXcr+A9KN59WRgdQoR5kAirQBQKMqyY1kLkuDVwmkIx+ZU3iqHrOjn3xC5
KXqlbiGYpWhZZd3H+zHSuRyLEEBXCo5vG1xNgIbm2JeELWS+m6H4e5nPGplcOwooqIsyH0R78XS6
GmCQhGnw9I7zxPoea586k8bLizCDqwv+KxpU0CiTIrOB4Zdp4NxgCzhCc2el05hjOkdLhUG5j+NA
7I2r+jdCcnVTlnZWMtYfv6mAirM/DZy/xOddd7CgwzVnVaq4DX4UFVtYo943nZ8plWPdlppWVXlz
5jRI85vCa1BBdVB41+VI3kliABSbSy6XBWJtjrLhRCpgDDrTOOP/xgDFwGYRev5mbeMNXW72Ayym
XSHIauWzPjcmcTFZufQFDtbh4nuy9E+V9TNE20qS/PAGuqEqOzIIbJTklSe3QgcXfXt6db0xhzMz
kxlXKhnKB3sWQ1nPNpK8lAiGcRRcxrppGvnjb0CDh78RWHXZg1D/lH1OE2p3CwCjPViRgxYTox9C
78M+ms+tdc89eocdhjOWlc1wckLw/CcSldpr32lq64ysqSGzmVrFjKi7NKAyEV70KWQfy/p1X2eD
PjhQpf09i7Cil6Zf2ImXxhGbbhLMd+y494UqPqrFJJlrNdcMvLBPceMByx0gHYZiyCQ4vxC86PWV
Sm5VAWddAh9sU5BLT8suLYw0ZndEiQN+mn6D3VGurT7lr3FHkk76PrdwzBUM97evUwHVGABGI3N7
lhkMd3CY0XYop3kPuFUz93MCy6ad1xnhityCAh3HuSlaaRNPAIHjEX2ombfMhMFBfNa1bINy/Kp+
tjAAMQ7CH5lx/01C+ZyZBiT/vpXwk/BCNxVyyjN/RVFyGm3shvFg7Z9BtGpimvsvPBsfT4hbhgv/
FbelxkezkpZbDQ3F04q5WmZ+x8YavIlKlq3jMW/fm7kg0W/b8NzVGwx44VYayDUbbbkdtgiJsECH
9XOJlAfV5r0tQNw7ekWfshNLlUhoz9AclFOC8mkWKUhjFAl9EgGRA3RVYsMOopIr249WFv3J9q9K
l7qhMWRdhR1S3AHTgO5jtevb+dROFVqreRvgEFO/oNYlqpAASxQjxR1zoTZLgoZBy11E2K/Oo4Ne
pmXaquP7xNAff0zK0AWYMDoh9TtZ1ohSJhV6MXnhLszNhQztQ6ovkGvLZa7kII7+QSZnsAW4AHwQ
+E+KlDbHy8lD1I22Xn2wk2CslVJGDo630LOghQVKiVQRY/qgIVU/m8TEhc8RGYwM8XF/zHm7z+Ye
qKWR6z6cg5f2t69PsjVgpyTCrXZsdqAr5IIhXjyPKVYBjPiG8YhDI9RQ26PBj0HLa5hELwltEUye
E85OZOLhk2c+ZhgQo+0+zdRGbA02XC4DBFzbOUQuVhbf9/J42FfWSA/6DW7D2tUk8AWgUTWglVg0
Zm43ZMcuyyCL1/5A2uSJiiPiIBCEZjhN4klhkczaMTKi3+WnkFAVIauPFSj+sgbB8K7ZRDrY+I/W
n9925+yMxryinfA9UnrdhRq0BZFmVRenPuxVoZf+zLGKd1XEPKlf3JSBHyRphcA5anNCIsYaeL3J
EXSFnoKseZ7c6NVey2wkel5Q37UvQaKvJeGS5yBvXLSmgDFiKv7KJ3k6KN/5yw5I9T0CBPul2dVo
iE6C2tkieEO4n1GnY2Dik4q9uOTB1tsJrVmbKLPhj69FLRiHOEqpf/M/5lAqX09L/693vuPYK8Xl
aBjmDXXrUfN7gKMO8lasK7Z5TdV3d8Wlpx1JOGmwiPM/GrbDPk8OCITlb82goCvyihWkb+pWIkBf
l3uajJ/7zuyg4+6We5UcK/7vH+x/+UVJhU74U/wUlF1Y/WnkIkws0eM2QR4hF0neQqNelfwKR29H
uMzsEe1qbDKSGdnnBt59YIDA69AItLyHRieO6lDa8oJThRmXVia89HKvJQXZwANbiKoMByA86QID
XuYJdfUaPha6HhdTRoN98j5kqvApql7QimHM/1f4RgHu8pdQApf3Fz7WPwDvnwFHJszy92XtNPW1
z/Z5gYvZmimCLrNtIPmNTWkahVLcVdR/sUaoVFkK/gpKvmPFffQBfzo8gdjeVG+MbKuIUEsFrEEV
FjZyYXgwBALXflS6rwEWTsgeybHUpI8nEJvMT+2YLOcyzwMP/Gb8nieh29XSZX+MphupOk8Rgntf
8UtLaglOQAxGDujTAo14o9nUlcWjQuQE/dZ45lb8rXvmWjC+zWP8EJUe3st4+T27u5Zc/LOU7RbQ
4Q8xIlmgZ0N9Tf6Lwuk7zMnxluvnmYayhquRXCrBT5D7svX/lKPuhyixl3XVkEqCbzxgIiJzhAVK
AMjFGiUdYvquZ/eaOvEpEX0kT3B8akOU9GyFr2FARofuE2kNDiFrkNwFaQ0H3RpiFCIwSvcvDCth
J0nWpOp8cR6AiIPkz0FNr54Xf8PVXlQFDINFifepc+upcdv4xaWY7fYSDr62/Rgdz/57dDQt76FE
TWTjTT7zTJiJq7A1NoC/s2b1hmWSsiFN67j3wXhw9sAg0V6bf4Z5dvg5zZl4XG/O53n/3QUZ4zlk
IEI65nDLvZAJOzC+tOCDckimAaIthY5ne3sz6zeyvsn8+xU1n4pJiWvsCY9Tqsqn21jYfnlbg+0h
OYjVsaE9/LsORnxYM/alQ2aTMOPK/38falnv/SMZOyO6OtVxHLcuLZXinnJFGrMGjZA6l3GaRVEz
NURdbkDWOiMSjirCFNcluWkAgBDwUwV95UgD0KPlWavZkp1RRz0QB73TAGiIa3Z7g05DMZn77S83
+mksE5yynLbxntUpdGLgcRqYfGlROMrAi1nVNxZR5B1WLzzPei+z0WtnDDUR+On/UKt4Ldvwkgb3
6bNRDnZj9WBsLyRbObw8XvYMi0GSnNnJ7budG2fok+ht0SgS74nG5ORCV5wAyJSCrWQhW1RKffSF
SDBBj+PIAHeYS56xh4eWXcCQ01wqGyaZz8rKQj0iEDsj2pKR9hMcZMFpOd6yHzYtAIaARWAD/VMH
6GlGxLY9arboV78kEAKijje+/2BSmN6PxLQw4UpDvNSvhpjgaUGzrDeNdPvd43Z6vrrlrE52hr27
Wk/PNR6Y2ltN9h2af1IouWFDvU+uieDQR53NHr+0mMBT5JqVHCvnIeAHTDv2pn+LlSKHMLyXNUpC
AiQgk/V8H1t3MkG699CrU5MlJwrxafW2thbWiF8ig2NLSQ2gID3sDyZYyAf46ssJFBy1JB2JdLCE
ANIpCC7VkpAjWsZWkrbFBW1SKH4yo6s7clD3ObwhFnhMJJ1bnIaubY2zThTIJnXc0BPTVvu74R5Z
QGo66qFTb8y0BvfqnfMfGW25eMusohIIwFoKAfc9iE3TynFI4KLU8gWbgNUUtHMKaYCYMHMylQOe
kGHiU2BUUAVu0H2f00uBc5u1y3j+uKxEItHVNUzaUZn9kZaqmgEncMGdLJCL5Ayc0+QH1/G0wye3
YrofafrKpBHcD8iXhbQFq+dQO2Y+uk5/chg9BVEb/mS0SqBkKeNgegTiOIghoXWz0vk7yCJx3hjm
sBtFEsMdQDeX9O/GRwRYDPEVdBoSrMbJo7+ggauDN1MjhfLjS2nFJbynallhU7R74WV4eQJEI1l5
tKVTLXPynFp8x0FsRLy7sjn95VDYl/mrRgXqrdvO4tKb+N68wAJEKdnwCiJZhMgxy+Ubwx/OPIWz
Fu7dXSHZS4iIPr0eWfHKR619PJBFQ2g1aS1nrZJSOxlvjIAF2vOkaSPvOy4ALXakDCBWQMA8XVAQ
Yxbawo6HMvFQgUOpyp9y/YR6vqKez341VNC2aCyuE+YSfcCrCUpBUVhj8sTDTgZRg4cmr9RtMju7
IhETXWtjS2AVXyrPGL+IOGGrHbVbpMVSjiAFsTjsZf0uYiKZUMLqQk8w11uUd+UtPvYdJq8iHVGP
EGT08Wbx+mO4bpapqzggjOatRjT2PDdedEHKoOQo+Yy1wct0GIX75z21KeVkcp+467j7/KgJg5EW
dFzeB9rsOxH7Xsbik6fsotBHSp32cKaqpldepp/QldXS97qUxs55gUTLrvtcsRqr00wSi83xH3mT
/ekk8/h87PAJZ2bwv6NzTMGxjdkw6cdOUZMPJPgZbXqsGsK5/TtmvX2UkPSHkcauPHCSn/O9d3rc
adn0vi1u9qGbqNoEqzp+hNXbt8ptvr49vbYiznbOPKDnYTfa9HrVOt7+cgXBTtk5c0QNL4sPPTW4
/3rka2SGUgqyVQxX4NiQrfnIJuzZhS1RydPultvVASpYACscKm8C8IRTzMEHYFQ2JAKQ/GBv8zgn
ZlLKe3r+C/rQp/G49+FH+H5e+E+wrUCxGKLVSbDN940KRqovTtqPvQ3jAGMLw+FctOv+00MHDp4m
2dtoqDNIaRBdIrRYwUHHJJAtrcAlm7YbsUOQCh1AfnNu5qUV84PjtgP5zmP2UwZekjvmnBAsNvAG
fRYkunID7zx1oMWDQHP2LUInp7/zCpuxdkEgaHc+OSbC3sqXytyRDEjfXnFPtn1Ry05q0DSAqXjP
N8mok3sC1x4cQBJMIWGbx3rXRW8RjekOWzMWGZnN5jZqIzCE1xGjdp68hM1nhHJ4Vmtlu7WADGYy
hgbmcVPQDCf/QMCqORTKo5zj+d/+fN9hkDeu2Xwmv0Up5PHksWbSSZ+jGGIAtkg5E9qvpQn6Fpf1
jO7YQOomcpc7gHbMYcew9Bzg0k0fZFt7q/dM79S4oG7L6wIvKezppczN7azvMFP4YZ7/WnjeYdTP
O6PqPWiI3wYip+ljoVoqXvopAJwJ3/8b2X0r84Jt68+9TBz7fCj2bNDiV2lxNJ0KTRRrI38pQqwo
/Qwymby92w+ermOILFu4OkaBmxgyGxIHyP75JH84amAQK1gSbVoyfng9MxwSqjsAFd+63Pb6W5N2
IJhwFTAM2AitMqbm7OKfU2tUaRiDQqx0ME/f5gaZniFEhzuB9tKZRecAS9q3aeZqrLEpkrGz+TBQ
Rht5qOmKOAvgxq+zbBpgpOrE4jNNX90WxghPW6H7smKrQRgyAg0cysR0WQiTbHxxGUCk/7pq/nhD
XcPe45moBi17h75H/lf+EzrMDiRP9fq8F1l7Bm5PoqCNMNdFK8c4W2RdQ14NsmNjCi6R0KD0aNe9
jJT9Egq4LyCH7DzzQntLHaWg2NPq9VFhmLL7RxP60y6FtOM2qmKZX4ds2N34wu88cxfS9ef57YIh
4RirXTbblPtHuG/rNA/un+3flr9SAQ4dZn6tu4KXN+NVYHmh7tc58VrhCn42Vs7deUHPcMK/+8oe
9D97O8bjIgppPDQeBxJ3z8gf9/E4nNk2s6ZxTC3O6m81BEgHKcMumFcB7bg0T+TmvvfRwkIc+Ik8
7jvpI04VlGJDXNcKAxDJZGlR0G2kTRrNwUwfxcBa90LjwgybI2lBTTipQGieayh8vFq2Ui5Dbtqr
mLBII38Ft8u2DxdwYNMbpJ4/XUiZUFt/KaJs55L9DPSlia3u3f1+4H15SYoFkGSavvv/2Qv8RUIP
oYItqHlcpcRDJM9jQh6sYH+dBkWMpJOzpG3bXVBTpa+hhrNzMdq70xGzFu7PCO2bFMY/BM+8jugU
4kNs8Cvheo3DJ6/x6ckhaAohgVHJR2QwuE26FKs7QxsGu4By1DtzrxddARgl3hkJWWxAtxluF6hE
IOFMiEtrLfMgL3TmN7hc53E1/VHTYmb4jAlsNUqIKJgghZhZTj3EuDz6du85YY0qB/+BBTordPnT
yXLd3tu3rCeOBDRJjXcocwhnwKBRCp5JfWc6kDRaqmueS1DQDH7yZM4YfTYh0rWD5YA/sA7jpfCB
N7YC8Cqf+v7o0xyoXAz2OyguVBoKGIz4lkWO1Lp833RfxGwL4W+seXs+NBLbStUom7f5vyCqAe/Z
yhPhsWEELpE4MtY+blvG74YiHivJ+McyOPJHMbYbn5YblPZPnM8KBtIzPlyvHN1YA/HYr+dk2PSD
lQPcv5SzZvW7U+EEVxH37E8CZZ0WwmCNOxsR1wIQ0dQ5/w8VmFdZLCSjSL4fXW3wHjoX0/gyfdpd
jXTwFLp8Xk1wTUtylX5KryslEWczkkYTeiYSIAii2XME9Ea63yVzfXqSJkQH4K3By5G6e+4RT4Bb
yjahZJsUQLj+5IH/FGYBlL9rbcqA4Ff15HzftsrjhL5Kxqgiu2Vx0gXtzC5x/2U58WucX7RmL4Eg
YxARo9h1dsuPgU3vtDdG2kP49XtST4BECfyeLyBFUzHpe/3IX6arHxL4nG6tpBk1kwqPt9B1yD/A
5VxNgn51ObcUw8645Kyg9Kg7gb42mImVsVlO81SfAhdwGb9iZlCfgoPcq1cuALxOb45Rq7n81ize
M+XpfzgPPld7Ah443uxWB50mutMyN43OydCOMOLJxe2dTL5bGz7yAT4dQXTiOEL/1Y1XOCwBUnF/
Og0gH1V+oW2BlggmV2VeBihrEzyBbEQWFlpYEjzg2eM2HwUkOsC0bnbk6CxiG0+BrjNLA6PBuRTQ
oDE6RhQ0JABvmFN5XytW2xO2K0qJhL0gd0xRMrobgneyc5VhWgTpgKMLY1Sr99dy9r3mNKuWvqTZ
go8PnITSBaZWAYHNwd014JBLdK9dZUDNw3dRz0qNZqCPQ9On1s6lGsnoJviR1aSIGv03Cl1/wO4k
DW+YDnAVdLVAs8SZVgwMp67rYRhv8Eur8WeIIi5+rL0WlkZx/lXT2Ymft9Z0X9Etojbm1W30ZRt8
t6dyrGpMgMfcxpzlRTF5w06DbSGkGZi9erWTTYj94xphXDqaWxkKV3iGI3xE7ILsaXJq8FR+7VMw
de8a+vzrKQcd3FlooA4Rf7HDnHgPsZMwN/mORu7SGxJdZB7xjpoEqJh2RFvH8/KM9s0WB09aIkNm
DmH9X3m/oyJWqQJZvLNNQP/EGxvMojrfHHoDaQsBSEMfNm4AsN+MysJYBttSk80z6/IV0yzdu5CQ
/WhU5vcohyopAPDGb1iiibMsZAXqsPNexzMlL5Q4J9wVrubl1/Voo9q+lsya69r63DknIOgwSgOa
rg/h/nT8SxfOXofw61D8ag82ll9AuJ0JFyZGQDx5R/FcMSuWmorfc2mIYRAu6MAHf3mxBlDZVBj/
W4eKxDhH8xPFmXajLPt7dktZPXEvlfgWY4QGdf0z4PWNej8Ek6sOSzGDOcPIg48plDU70aej0vDL
P/l5OAu4T+nqWnENguNNwu7xMV9Z7Usfw4ztJCxBJErNKhFUgUmCAycU3F9FJyOgzq2ovFzcWz4V
n7KH0gejQzjnKGol3EYX6t64DvmVfmAP4OzBeHX9nmgHBNRn8HlAjIJ+zMZlIxfrTq5I9aI/+owR
Isi5GV/iUYjoHcBo7q5Px7cU3gRFYclCsslc1I9Cend1XgILiO+RX/zlp6ut1oj4wOewXbTZHSwn
VVs0taj5nDpoEZb83fWiEyk4mi7xzDMQpUG5MT9lSvNvYtxAnQT3dNAO5Gt2aYzLaQxtUERfSNci
Gb6V921eB+j1/EVuT3JXgFWHNpOV4iZz222hlaurGRp/KTFAwUTSsGXOTg6gkM1ZBZnDapuGRpa3
R7R4YieHl54uNMc83qm78TOoFiwDT7SBV3cHN19sI4cPEgYFvv+2bGic/6qAn1BpMFjHOX+WeBG9
FH7ew+HLIWUtF1xN/hutnp4sUWZki2cxW+ZxaPYnUL+eMkkLzmBucc2dw7mUE07PLbPpvm6oDr+r
2dWCKqNA0JZN/PGE96KEO0st7su6pQAVHH4UvsPqaPxIvXARfGF9obT14zr+au5zy+NctScV/+E5
tLoyX9SmCPfSj+xwZtIJ0PhE1/UX6MM/VeKG5UWL0al6rb9ehGKbiAnNk2FINSMBwRkZHXR8YvK3
AlFLaiHfZGDo6lHyK6xof3RdU1cj50j05eJSPRwLxg8YqCTfynFmhfRIQt+ImO4mtkJwoGk863Z3
FQ6NqYamX/lbbfPLWxBuE1WOHwV4+9CB15LAlGluT2gGEwWde9U1n2S5yTJ17AQJH7HcCRe0pHef
Y8MChXNLGkornZbze1tJSc6gsyXIO1G6uwq9JYky70YyfMDUTcK/eD2HjF1RCg+v6GmOuN0TUD5C
Hm2HeYiD2bThtMq0ZSyWmomDdFkbHAcDxaGYs/9+U2crDhM6zEeyJuj9Hdv0cY8Ee/Hd1E3KUH0a
O2TXvJc9S2Tpu9yofSp2T1YrNEp2Ixnkw0l0n7yZ1wFmz/4OMtbOjZ9ubRfEJfW38d5ijNgZ1p8p
OHCzufr8Tb71qUTscdUN7RyJ4yLJ+UIF7PMvbvy12r0P6JLSlFMybfgWEUg1eM6opMf6L3qsYOO7
G+ry8Gip0EvP8hm3cyxJxZ/Yi96BxKdneKM5L1HY02BDHPChJfdkTx1ziXx6I9zYavIG6t0CJV7h
8V4X72/Vndjj3KvNh37uPEOxETkTt9mu4L4GSMHXUdNI7x4RJ4ysBf27VqAfibkWLCJ7z1HXwTNe
mWYd9hPMyOSvvo0/2lm5wgxOnpU2vKTBXYrP42m0wjCMwVEQojsB73o/exakS2eNzwcE31Xc4ADh
2jQCeHUeYeF4viCMYL2QJj+GUW2d5Sv/7OojE4gwFQcAZnttKhTGDh9T4yd+ToEhXxpzJ/iF2SdN
m9ZaW3n9a6UPjbIi3k13owI2WiuM82KZj1PK9VQ0ydciNGbwXMAT3TMWp7XZrFXSB0LA8ZwMx6fc
rtklt5bzbBLkk5YXmUYZ0d5KU6HpxtwsNRfb17j0cY2pYFoQTrDh5P3Y+sHVf/xdMMnqUNGQdJ+C
wbz7/8C+EWv/XWxbTqpGyZQiqMhXfUWJ8Ifk4RuAla4+V5Ww1pNBCAFS1cotVBlEiWEt++PfP6vx
Rzu674JsWZuINIs5LOUvnXL17StudrDQREwYMs92TGGRwQC7Lg6Jnav14H7VEG3F0+OUbDvAJrP1
PwpoGugpTLAXMnyRkMru8AeY8+F7yPAi/xLxtorPFL25LSUxSt0JVtgUTNC634YcN+SLa4YvEVEX
HVaZv7zR7Zv+fsyYgussGT/DPASRvlFbzFWB2t/vurwLzrg73emjgp/AALt8C0OftZe6EIbGJs0y
XauJSrJK+0koEyRY9x6vF5hjYMU4bpfpXY4KI2zhj3kKf7IyYhSu7emzVByqSZnpgoa6ltd46WvB
2c98EYIqKh7P/O1tlp2rEBAhxY7sKgQ2+FFTwoCGN7x0xRE4Pt8GEUP2aIH2L6gDKEHyWTENVtL5
8BsJXq3uyh8403fjibGyBDBZ07Aa/uTW30ZF3I14Q2cbAQmvTcGTWIY+/CR+67w1xmxsS+ZZEQtV
oKvfybYhRx2TUM1bFjHmBLlolTbA60t/yxk4dW+LL3HwBciUaJ9mKm8mYhFNZTzHOZQibEi/X35E
xGMbT5YMWnOcDhe8ILK9lZP68vmr2Q1zILhMM4VEuNHYmAQPjtt18Ki3eJgcSD/Hgi6moddPNkAn
xcQqmW2UQAscDq5MQyiY960QNt3gPzZjGoV9HwAepqHPJI+hw2JaL00iy2TPjM2S+S3Mn/jxm/1b
tsIs5uRmTWRoHLxx6NcMwhoKP9m7MX/AawbRpDjwfnD5zAUgoX6noOcWz2KwIE+a/qJObGyAKwkN
nHAqy0GZagrJP1bM1DV50rHyYS0etZ0R01+zVgZgKA3+oqab2kvACdQ9e/8mN0LNSYqFoFduOqBX
df7ScW8UHinDTl3kugkt/8nDhpQ3C72ekqy3VHj4lxmTGT9Ot5WXxnOAzUBx3kfAzwoUSw63WKKg
xacRlTYs2b0ZikHVtPnKODPOFJNm7D8sdgTiGUsrvv+r8glBvyUaoJIet0fkOpTBKGy2jzOU6Vn+
j0Uof9ArY1etKh1imE67AXMfmaVqbTavY+Zpv3j3qNWV1e7VPMvn8iPs4dYHvJH5GMJm5BpiJiPJ
5eGzpvMb00Kx/PQTIKChdl0fikL7QWk2h32df+e3RsEJLyUW7mVGgxKo5MzrfGobnpgOsoAQtNGe
43cbiPtzYoJNRdm3TO2DQEhlCjIRtNiTFTRjXQRr79vtn50eO/pIXVhKQ94oA/XwSWWtXEbtEWLh
haI2XzcaX2iDdeFeTYeIxik39Ys9V3f81RtL9NTQAGATj/91axzatU8cMlV/dN9LdSPhTuSHBmDU
kX7EOf2BvpjjdzfFMcyebhhM3abihm96RMxwlf/gSNcsnRIZpEQe2uEioSN6DtTjnEebsmLkS/0U
F/Tl4aaJSWv0qtWDbvziXyw4hB6AbjLO1kum+7NXby9HdX9ZDjEd/WwaCNkPcvAvyWt+lbqhT1+9
Y9zMnOsHj7ehZP4nwzqARUbRvOazkEApROqSkk1ugqarsOg7zhNoiOog6WOZ/iuC5pUwqlFEODEf
NNGtNWYW2yL9SJjuSzfz/4nRJ+SxhU/taQLmuj76+W0aLBR5mb0CdEipqF2NDbMFBsKI8x3CoM74
NHeey/QAUOqj1BrEz6tzHzaeBjOjhZRydKo+50D6OQQtONZZUKD35mH0vVlWDP8VjV3tnBTvP0PE
2Z7dOtijaPmwoGISsnihRyAi6CsHo+RvrAVwMGToRAQgoA7neFQZsYILm9yvpzcEW8od6JGQkJr4
CWAeuDudOItOnpoc7Wn7HaYUdd79ud0iffQquHPPY6MdFYxpSDyJKBtQMJy/FAyV9mk1gGprEJuJ
g3TfF7cs33tJOe0nhVySgkbMWNFazwE9UCt0H6zSLc6ZuwA0zhdjGnOpi2xZDaOojDGDONVVG9+B
U1ZoUQeyz0e2zKVEK+bN71W11ZG0NkpNnMp431L3I0XYB8nPVR58p3AniApul3SrRoQkxwe6Pwyz
XO6xOmfetcA8E0fbxpEI7khGjxBswZwGtR+IWqhihQXEt6wB81Z9i9T60KgAl8vvOBis1iqBTOac
HWvjYZ2m5QU/ckvSpHbUDA2Gb5Z85oIwxJC4i/lrHoZbRn4lL0qeoOME24/4VK0rAniPlh+ZzTvJ
vXxJ/BWimC6H52ZLa+f2ZSf+MMybCEKFU0NteuvWWv0zz1W0OyB6oD6Bxa0CGt9vm3ftHA/ZYWBR
lCMFO8Vzu52ZWF6Z4lm2jqw9IKGNJt1UzlCXh+PejdGaxXC5Ojv8L0yNfDmYs648THOpDv61GpV3
FpsfHJ7+JrdFocuVzPqr2haXopRoWlB4Y9t8yY3XDwN/PoG42hFEJSAxfixFaQAIT9HAwWGkPGWn
6aH+OQkmKREQcul06fZN5sMQiY0A185rSlggU3KwyoHa30A6EXMcPzzi1QoK8zpMvO/DO7moGWME
YNhDQcJXvPKzE6/L+5rNYJEn5sluxg4KLr2LdFR8Cp1ITD+6zyb0Oa5IJ9oKaEwJ7YjQbvGpRhN3
y8wHvaxL8ASbXtBYL6K14ywote6mCoBYEKPiBvajONU51n4tK1bOTCh11c3/9P5ShWDQFRrTx+Ps
CWUb07VL9uGYQiT4rjrdU7c14ZYxkpMsTu3nei4qSRDxzWSM4rAvt9cdLLPS9pck2ksbjXY3ogtQ
lrYwsznDGpGY26Cn6mGqfJK//CKPhNEKb0gxX6q/4FThYtkV3kp+lR9vC1O39dZU0oSZ4N/5d2u6
YasF2vwXTDnOfz86Iri/ZyAjFazcKig5EgzDN/9lDs2sSGJDCEcM6q5l9tYQoORT0lQn7vFhmovt
p36NebsCjhzNQ31dSsbby1/MymBGmyDCz1mx6UaAPBEPJpWYazKggBHF7Tr2sWl3DlbIVCscKAcE
YK2+mBHh0TVBb9m9pA2r0GwJEwgvVVWhze8h644pik7WvJ9if9MvfeUvsqiTcgawBxuGjuLTdEdQ
UloSm7lH+TM11MiSG0loisibwn5XWN7NNnMs3BN3gz5GZOQQ7zjEnAGD584EtePlgq9kFrzvQV2q
NATLPgxBtN+Qn+QorSAC96Hkud/HxkyaMezXWHcvriNrV2kLdp9CkZlFiivIdXMj0Al+mHwpC+nI
rpnjTo8NErafco54zZOz3dZfSqGMaYUTMqDAEk7KL7H/OYtyfviBanvCtBwiBARrDTOMaymlxrxS
XFIP+qygl47SdvXbn+d98aljyHx/33f7TV5Oh7KtDGK5gD6YpjXcLEHcBgLiipyAlJP4Op79ed62
Lrn1wEZm30Xq8lx7S1ZHNzxRq2Rb2yBd1Itcauz36AfMloZfgMglSDgUtWBhL22JGdLiWXWzCbPB
/HshBGCPbNglNglZ6JSGecwoqe/483S+42GxmZiZpAtQJI/4bBvgNgpJ+DxXv2noi4vovyN98MnF
6WOqSoe270NHKuDs1p9Mmt5SQoWfLwUX25dV0ULrFAvRqH4G5x1h/tm44rtvXVkExRhUDslTGfCX
8r66h0Ksm+2JyyYJfdEEqUZ8XSFcZCBzzrxQFU3wOvQpvGx62ljjmLDVOzJTP6y5BI5N49Vsu6JT
rDcgfJyoDhQhyn2aj6bZio0I+NqTLDkZk/+wXovKZWJz+kximd08ofRV2dkj3x/vV5XKB8NqCAFs
ySF63kXmPqF6N5ggY6/YHkUzKFXqtorN0CkbHjjDccK7z+Aj+lpBZK+Zoo9TQjwdjpW4RYdQsZZY
pR1kCuMPt0aR+6LYShxSoFpE3TRI/J7pkmgi8bafmUVrg372e4Kb3woixWWjxjXm6GSRTRpaTz+L
XA1iKyeAfAP0Rm6iWxUL74o5ZVEh8Q0KluZAZzYUc20oH7cA05PA+bYeoNSNocgIUbprqE4o0wU/
+4nl5JVibRXHdLnxTas+ptXbHAeSyaAt0tqU/w3CZ6BO6Sofc1PcdaTRhswXcO1QI+wVJajaV1p1
ArFLNooO4X4PvpBNB2TSjOYbXjGfY0vf0Ra4yeLA684McVvBeJHwgXkl0PxLWO5z26JLExxU8VmB
yqVas7j8N4T3mzx2gXzfGvMMlOEk55V/sJVlcKMTFEp1hhNFrwqJ+NuMA1QNlUG5syvtY9wHYklt
E0KjNC7vLIXdCVLsITLixsdQYbTtZ/7QcYSKfJVP7Dt2GpbhsudrlNwNLHYXK7qnFmbi7W4ncH/s
JrQ0WY60CcvxkW67L8zV09gw9Qn/+0kE1+w59XjTKlRylhCM8QDxiBpGLUOnJj+4F5EAaMpZQqos
Ck3q1IEtvrpaM2g1teTh0N2OBU3zyDnmSmyZFYuW42FJCAHyCPapsWdgnTBjsKMPq/1UK9yKPrTZ
pprUWPMSdn7d4fVA9wELzDTb7la6hSSz8FGcoLj8L4EjKP5gB7BTIpXfCmBsYq30587R1lmB1yt+
Z87uC8tvkFvuET4ZwFhMEn2mhPGTe/PdVgAfly/+S2jUro6RFFinpaUz9rnGrzR9EpFr0QRdKtgJ
XsRBYCofTHxM7W+Am6NA69N6JCAid0JUbjRi1hfL8MUEHKTtjSqR0xw3Z6rEWeiJO4lNiVNhCORL
80jGhxl9bmcwDq4U3hwnabU29dsGUpqgkrKdZWZIkdWHZn0//U8OfW2AntJrxSaDwNlnVyvHhuz2
fWE0U7IgYukzc0LVqrb9OrUlM9sRjPy7v2UDGY5FjLEthML8aMVIWBUqcevhVVNSy5CepIJWMAvi
N98JflDmKiA6XMAOr36hyigHWG7o2pvkViDLiywEMXpwp0vBL5vx+23YgPSGlOfZYVM/R1gIOljQ
8fvGu8xK4VgAOCcJFrZ24SV+ubfDSreutwLEkw+cexrh71WhHCb09kIDjC/733T9h3UiKahBl5p5
mmTGhAnd1o/E5QaFl9VGQLkefEfD1HzaAoOSlxCGidc+ywaI8dhzgJmObQuhzhO58GVdx9jIm7Tk
NXTZb+o4IzW+Wg+/FyH9XFCjby1tNLRgvF9qtrfWkXljuZJzFRblo35YyVzSkk2PiPkaQx2gXgEK
ASBCfwEsSGrfgJ4B1Z0VSgQp7wOurIHkDsayBj5Lbcfr637YgdGKugMQnazu4927R2hWgBzlZ4Jr
kOdE4/OODaV+NIdhBybDfOU+V5DgrWa/FGF+DZHSam+Encm8EMPeu3ebyNhJIX+NXeVZ5qgCM4+k
SVk6FxFXWO+RrYZgwN6VN+JCgyILHZ1dow318YLU6P5MznLYoQ5BFw2j74w04RaswkDOOasvnwfi
YRZ9YB6s3cRK8zg+E3SywvHIZBshV1gxq0mLIghV1uBISV+R63lGVlcmbAmzw6jgV5FcivD7M4al
GAilFZ/8ImdC3FV5RLRI+ZovQKiOJOt25rixhdOTIhbNLp91U8Lj5bz0v34YJ4h4tJ4DJdgBID61
UJ4IU/iZLGB0syx/x5Q9+Eoyjl9OGwIjeAk0Lw0Idue3gv2lJd7rJM6oViTcWuHPiNzLQjFNapOY
3LVyUqUNNXE63F5KIbBfnzU4Vwbhjyt6IeybjOmRY7oGDO2tQcaDkp+wclLNdsCDwAC15yqR6jDj
7jSEiDCB2Sfucb3VFUZCl9wNGa176V/NXTY+vgaAToKDacmIwoLN5u+/GWSdWdjT146iypjTnyyg
McYUdD0rXnYm1cAF5+k/zpxsKVCW1hp6zKxIXtUraS6tOhX8qAJ1VRXQcC0D12JYb0UvgKHLPAGj
iHSpi+yWMb7Ir6NIED3RnNAsFLCbenqxz/AqnktdibsEaeVziqUafKtLTv91oom9cez/xeBqkdNm
Pm6Zdv0WH+QumNAc5pxuAYvQGqdKLBsGqd4eFjXHeIkwVG+3LsSmVPGmFdCG0+OJt1GBXNrWbu90
PRLY4zUdImINdmQjgzjJ48IRY8fqY1462atu09QppIjMXQCXbbRWPLQOBWhZ2wuJ/x09bFB9lA/o
YYfl/ktHnTJHAGA7u3SUe7NBzKexAgy4aKxGCbCBNE8qKenrlqsLt6Vi4RGfSUJQprwXfbCgBEqz
KqqAVR2B85I/W5o2ESqKnzz436KTQY03G1ZvYIhHYmZX5czEFM+Iz5BigZ8iNg4r+2GU2ehgj/Ve
qIjqCxgmpaGkNmVoK4+TFm25epmo7Cx1UBwwUZxpulK11p1OXIvtzsybZHGecBRD+pOWn1g2sCtf
5p7AY4bwkVo9Z85HW4MZD3exvDZJkm2O4QnYWs4f2U3Ec5QJbYvp0faukLSeJGJ8ptunOqyEQjlP
Ex4ALWFfbmFacXJgR/B5Ybm+b8x4oWdwbxljkUobvmt2Was2Gg1m/m38mQVh23KpsSqyOc1P70Ws
/Hq1yoRE2dg2JXZR+rkS/tckQWQFuVWoidRUVOdLNkUuB2FIX3RJEZtrYKUIBuOJuzWUQXu3JTLh
2WoNuj+70uV5mJQhvBTwT5l/P2x3UYvcit6Kp2h1YlGekZfS3+ExjSF9s7V2J7lRNfHHAYCYd0uZ
llNK+tC1bMfbY9CviQ9Ob2IGaTOF1OyNKFagKfEyuTSEMA0GuLh6B8NkHCHW2KAvOs/3dHUSIxo8
/7mDfRYEcJuuljnwdJkxmSBYK9W7aI17oy5ddXEddzJCLGoqObVwFkll0cNeOMnWNV265PHfZ2+B
V33zl5OQfTZIO2vveX1WKjpOubcUVc7VaTlev7f86nzZA7ir/QMzgV1IbRt72dRM1OTtLfElx/dF
NSXm4JPNPkLCq0EE9tvNGy3PEjSeGhadFVOr67Q6C4DAVwdhc/6m04yXcRx6pqt773FAciTZdj8J
cA2h02qcJXEDzJ1Mh6TDs0swa1hZrEU8wqTCq4EVaWsfQbN1zKTUje29aiDyWBR/Gci3eyxy3xsk
4dVnrid+/OX/EnbSfnYrVSqAVcKHXL0oi9GLzRftuNNNnTbp/4ylbbjxcG39qPv6tCENssYaX+0A
oyyON8npcW4WqZxt8H5DpdX9/wtDWB2hJQEiJboo6TzAgWv+t8BRQVlNYGX6zo1cX6FyjStgEGcq
QRYJ/MEs0c88W4GqT9J+jC5vBENyw81pBfwxMQKAh4pfwQQi8FoaMbqTZvKI+7UE3Wya7C7AUNR7
fz1dR1c84fnbB1V+rVX0hpy9WO2gOAUDjJz1Ddc0bTNJTkyRJH+N50U2IEdv8T1IyBjJpmcwCLWx
fSSzbSZt7oM2jun7xOuEuoTm/w7BHZ5LPzO7U9P0w6YfrWT9Tti8AzgKpZ/1Y1cdiF944p55G+JV
wcS4FbnRJT1Nig4XAJzN4ZmzKJJip/UIdJ9hjxUICmC/6qFlJWKwF1RPqtIWggkL2NJGW86EhZBK
SkOV17SUeP6lSVbRzAq/mAf2Hfjo8m75YXuMUOEpHuEf50CjkazzcxSnF6Np654MteY+saKu1u+9
H7RsLgzH1HtNE75k6uFaum58ZhAs15QtS998sttmDwZyZqLDsh63NsjXuxVsZvflV62i61LDukCK
mEtHQIFnnm5eDBykMWBcqQWUTAIkNPJ6S6MbxLWLfzSyMAd3EcLIF7c0fGJvwMld6nIJMXF6d8T4
fo8jakR6EVpJcGrcAUiKjISJnDKJIfvSKGC2roPRT6vysBxqnmQ9bY95qBlaAOo7DNkDDQULS7Qs
Nxf39b75LA2l7mAQYwJMlH+r+AMRc1iSDoHkJbDBqm6dBjCYtuzJdXuATeETNjPgbIwaz1eKrwmP
WQGGouWiHMzOSWkrKwkAH9nbGZIOlGF+wOgeIShJF+0MnKF9U5tOHb4psQ4LjCMMZ9vxoVuZwe2u
UJuSZrlRPZidqPm819UGMarJ2eM+zWOMa4mUDf0gEz/2exHEVzmlFDCDZ+WYrb1Aoc8n5O9wne1U
+vq+UxGCqiTnO1gCeZ8YHg6QOTPpN9wleO5Y5OrFRkDbslve0cKJfY+sY/GXqGM2zMUHwRZf0b3n
Y6NdDzSBjtuOsZHIBX1gZk8/X6zyzRAdrb1VBx+riohQYqqUx+C1Kc9GeHC8z2s6vgqpRRid/yUv
IL5OM/kR8sMqCzm2VBlsA9HckdjqiBF6rQhquVRgm95oV7v4DcoEQPcZQuUTVUj4Eo8u0Wvf46Ot
MH9c40OFGJ24o42zi5opdp2Wx7365VT13hk2xd/IN4dJCECEIV9u54MmRtNWL7kuIfkFfMdbxgN8
nlify/exII7PfiUi5Chgwz2CgkZVCNFeOEzLPFbor+e3iFWD4fTBJr9iEGcL+qWCddIKNGI7Jn6s
dqYoAIAcl+3ll+md4HFI7gCELTFMMBQtKreZR0QJlW0qMsAqrypp9IxbrobmQS76OU8E+K6sS4qS
gBl6kVzYGbJkTkgyzwqDaVTqZDAWkoRFXzTpXD1CdKnNET65nb6d2rH3r+0/SUmi//AQwvSwV6Kn
hvODzEXMM9vHxaP9wMx3BgXS0fEj4ZpjrK6jS9wPnqMCva42NIUxVCQ9cIHkFiLgsHOw/yQXM4U+
YTraNS+XOaDnRf7ZOn/gFEgY6O9PGfZjuhWC8zZHGHDJ+XD21EGIt3IVyj3cz9kdtBkWfnrGTfOe
5lvHd4xwNcFyV4komiI6dRKKqjsCJuFxUBOridK44IUlC11F2CIw7KZyJlg9iCQUeK98ds9c2yKs
Qk9kFfAmMZgMNftqXexFOIcx7t9KREgtdU/ziQ4tN36auxm0X8AcWYsTLnFRscsIT08CyeTVNg36
0r6+V/Im+W/72eSygEKASa6FOd/vMiQPEVq1VIGi/x/JDmjl3HCFSoXLMqeS+5sMegFJapCRf8Aw
tTtxEwMnifmJxZT3j3uzSVqvUtREJaUXJ1mFpMHuD835NwdmjvwLUqAbie/ZPVw+0ZIrGMNl2Pdf
/70YLYmxsDw3iEAfEr0UpMn3XDbjiJyN1D+GU4Al1TCT7w/LJFityNrOWhoy6a91tY2QqSeslBEc
pDZ5D0hhgwkwA74aiMDouh7shkiFLClOvqVQ0sI6MKqT89O2CbbftEzh39w4mHIXmL0rrTXpFU4I
c6EgMWzK1rHjDVtOOXdhfYzstgbiDhAIUg8TR1tQm04dfsbKJzhXSEt39lvXRnuD4C4M87pUJUgV
ywqaqCkRR5U5xsvqgbZjN+m24E/Br50OmD8dMRnE1tv5wj3hguVstZpAvMT+KhD/5KVoV9jysTcG
El6WPe/JkYjPthNZnnLKOZTSqyABlIJ++FoqEEtj0aJeQJ9USEjxT4/puRGf/yGIXli3vcnJolb/
2xKJK+ywdWG8DtaLZnlrgifXKxwCBR+EPV2YUzABXn0eJ2kjkQEXHZOagjrcHvxm5oMrkSKy/t6Q
MQbIlTprpJsUkNHa9zUM/AJQQ7LmkuMq7WksrySTduGerTQJv6w/9Ey39VgMMoD3eDq+8tG4uDE1
whovRzbgkoIF92BLI41rDOnbU+Gz/gu2RntnFfBjiV+oJacsssNXLIrRSBwKf43eOIMPgkdg7cev
4TFtJrwCvnJUyIQvNsffPVPbhTz30/aWupRS39IC6t3e4k6NACuISxOhDbdcr+A4aALCpaO1B8TJ
zqNTLmfmsUmw3J5psrpzobg3sDFTvMd3un7FEPVYQlqacdREaPU7I9/ewpZWXu1k2l521Y3SCV9U
ZB3jCuV/9xNF2sgEJc1/Il4HaY3tUCSX2UDcEF9j60umHndbLPN9+UJzZMi7XeQmRq2MRAWFb9QR
0EVrs/Vdi0mPz1FmPuHrXC3L/7iEjEH6Fb7h1QO1ZXlYDe9NhkDdTKm7qtwLCm/JzcluWCBOebY5
s2+KfSSx7RsW+9RaJizvfqGmn1Pi4k+5yJ2WtHRN3KGkxZSiy10zi5kOsYNjGPLs7xLPgc3nU+mq
Y6muH3MfifX32Hvuee06L4OvOXAFAMbZTTOhBA00SuLvW6oAVlXG7MIo2ARGKI+HcHzA2MSPqfUl
K9q4LhQq1l5TzrrTIaP1GY8rXXAP6ZmZ/9NrvtWXceMv4wkFDvMwZP8ncnYA90TApgKBEEnqvUsJ
HnMzsyVz9szXHVll+1lvps9Fas3bI50V8GQx9TTyqcuSXF06rEGelWOpOGXPq2dvQQETMuX4n9de
hoo1chX/Dsy6WqI9wtQpwihYUNYlq3qi0KDNu08mNYJ8mIe/IAMpf1phUlEstAJK7Kp5QkJaWlFp
tXQlR1w+tT5cUFQPQb2F30zqXHKGecDfEyF2I5x+j20ThFTF9Ii++xanxYD7zGI5Otjs2b1b6xDW
Q7ns+norN9u9K+VY9ul/D71152cGNt2ERWWySYi0CbfsOJHAWS0p8o5UV2844qraVZZgZzZU3xG1
gb+dXdgQ6vunNYbCq8nI20egnaWq73vEO0oBBq4ZvGNGDpy1ZRx0vLyOxnF9C8p8AR8yX+dHuTJ5
M1/re7QT4YSU1w6FtkeV+YoN4MuzTdzEInZXFKX0/2NQxJj5cC4PG00WpgSu5XGxK9qDXr7iGRam
wnFV3cNc5EHzxDe4+y4NYNfgqy0bLZlME1ty7uAWADzjfuCs/13k7fVRJRAdeid9iUhs1IVQixVp
127h9GYOAC7EsyTl1KcSiT0U7VSJVVrWDxE9N/1ldEqUtVeV/LE9vl1L8FW1Vp7dSIgolZA99QPX
5Gia9Ok8Qkv8thRgRj9iaNE3YK4c26HC9DsBia96MAXD7gV35VmkDuKUlJZyCirNblpjIca9GUYC
RdKESMy+/TBENpGrd6Ncv9cDdj79R1cCFV1JtKB+AEeWWMf0M6gptyX6GHkLWhLD958aZa0oyV+k
pEe4kaaLmEFlUYiWNz7XYeEPDvI51wxfktSirCcsIvWDKkxqnrR4UTY8RSP0Ms0iYag9QXyi9OKA
sfjKemI+OP2zwaUMgox2SwpoYqYcemXP1pdzUPEMy8py6Jbgb26bAtoCiLP2LWJxG7M4sd5SQtIZ
kn7vdKUgN5ntfSibzHyRwtQOQXejQknOfGOU4jYq2NvP3YDdWZFnmx4z6CFCaKqFPyh8U6y9TrZC
Kc1yvmI4k0RVRZnGHYxnOmfQuWDPzxeURWe8EKRqIxLS/m2qFSiRjF0enxK68VBM1ncmftH3gmrI
RSYfQpfx9uiz+kvaPkwFfJ913ckWMeAEG7jGSfqNAVK6HaqU48heryBoFGKfinNeXUjOKcsSGePH
OrbUE97V62S0gkA8tFWRPYZsLpnU/g0Bz6WK1YEzEXlKnCiz3nuE1kiRrCBqQ4s9o6/N3qcQTl7t
CcDT4e1xdKj05DVJA421cLkX5rFU/DZ32t3iyfTVH3/SL7IUoXyKJ94tzkQHjex7qbWkMK7cL6rl
DuN++0om/X/XmPJSL8F/GpRnetOAaV2FtI0To3d4jp4NN3BIXw/AIEABlVtLjcRVBqNjQCuxuoR+
ETTpqFM31C604kW2716Ml1Hozyn51bPnaF73CySJyn0DM4fFB7C3aLkzNVLUsscD5+0QI3nS6juu
Qayigt4rMPulfFvxTOvQsWF6fxBr58DAgIZYlOI1/E5SVuDqacgNA9B1AS1kdp5S+oM5YplJETHs
1g8KgpGyYq3EssKc32JppJgb5h3/JED4pOyx6+qxIJYYFzraP0U3Arwa1KWC0ZyJDcCLUs2SKZks
Jf/ufzw1Z+yQivClvum3xJ82aW7sIkAC3XW9jJQ3v0MtS1e/GxiyFhn+APgSDBwX1cGkINCvoDzE
ME0dVEPva7Ga8JScBXvKLC9oYSVGO8IaZR8pF2bv7Xu2s3wYMM6BBQG4mHvtw30JRnbldXmtLo5A
okgVb6jIdztiFLrR0l5NAuth3Z4BLjA0ErXuFSpFJHE4lAn0AFqVWKmCGBIlDqFOmy2FOiDt3QHB
hlyErteukjhLkqwT5zDbQsnwacfxctF/LocarR40uF6sdyFc5rpKjfe0IyBM20T/QYVbd0YwgmvI
MommlX6RUpqOZmOzbVOnGFVV82nbCmDd3AdJ7RvwmERrcO85pYfVoPsf5xU2+UsLbd6Vp4q36DPL
tHycmKQJKAUZxoRI6Vmwjea8iKtWaPKKiTe/aklWlh5pWsfg7JGcMgTK5fLTs/yIB8XbNYzh0thQ
2cyhHzmZKBnVkVaZ3p2KxD/Tcz38PFxmJqw0w/TVoYj48Ua5nC1BtumvYP0nDtZo8qKlJEP5ikAt
F3wLOdgzUVX+8GoTsI70pb2dsu+Q7SfNBd7aqw68syLH7UNYoxmOBaZFcE/GBJ8S3bkVRQHSlUK9
WdP0nnsxeZ52x4C63J3tdtJWFB3arRnX2XfhZHMhBKW8fM4jB7qM4p6RLszNpnFzC7mvfVSwMsAr
icTYDP5+uDOpdXGCvfy14jSQjvc095GU1OSS4oPsjJxfvYwvTbGfb9Mt4bsTqde1Lw6wyMw2F5bI
MmwRakHuplbUIiY7olslM5i2Q9sHFyFed+hnozhg/ki/n5Qt7ibhCS7qFvpIHsAGMIoz1j/+H+l/
nMzZjO2MlOHGi2RcaOAdBGlcuT+jP31+jKGwc/MV4maBNCqhV7wobtf9GlIK7oTNoOATgRa76XLQ
X8cDmqt8lmE9/SorHi3m0ymzdgVe/gjJkuLoCbjSQIk5hGXTlTMINH1q5stP94CuMIEv0EuISFie
d0YZNXab6yA+lyAt9zgCgMK+WAzTHd4GSUhYXFtHUdQBbzx5xMhqJ8DJFsa6VgW0dJszyY3TfD5W
z3vNUkXBf0GQyrmN4tHiVmqYytcTSz+6BLviPhymGRX8mFgTEPjunUZQHbjbkmrGOSmHFWMGHcwi
9pGUvMoVzLNP6el+Iu9tpvCZWYJeEgrIKM+KHfWG8OKwuK9r52a8ydGVgC1kqL5L82frNnuLPheA
e0BAY0inu0OeyApmhVju5S9TzMXqO7IZ7dgKQ/vI6Ay94NMdzSTK8hckNMuBYas4tkjtRvm7uc69
3GLPMu3IWzhXnv5icuHZWCg9wIId1tjk+/vg8MTVftzrmPg872qceNMSvujVTu/ke4HeoOfdPl5i
BwePp8IC3KE3x2VtlknWbNyiDuWw6AOmGBvhozzuoTebZaRuzHGPGaY6/GyyqDv2crux9fZbO4OC
G6RW2tIS//0Ju4nu03Rm3x/w3f0Gt2sBqQEpElAv7RSbrSmE5Uu6+jL3XdskxFo9CN50QyajNtuz
lXnQtbx4CRB5ofw88SdTaU5c2Lyot6KUjn1Xfa1j/DRTNy3gZjjmZ7Cbl1pFYKwORoBca1j95a/+
qd27coxYyFrcEWIqXnB69tSpdfQqNA5RhLYDJHDysDgNSyBbZOTB2MeOHwDbkYROVnvTT4ZN0Z44
CT75AXpFIeUPFx+hHKsY8JIHcrsIOsk5vq47b231XteSxwzP5v+Xs/r2TMkS4+R/FwvvedXV48/1
MiCv7TtXRRXY8QFmPtTu01EFok3r7k0FHpq5RdnC4vxDblZ7s5poEv5ijVJlxb9nxeq+dRk33az+
fsHPRpWCkcZ6dLR2dzJgJ9cB86rWxL0gLDac4zE6BE/02+VDpGp6d3Woi8Pis3dWBe88ymE6txuk
inAp/uJrn4tkHnRi4HVo9NuS8dteCKU/IBGE2aoTqE9j36Cjsi8G+OE1Ue9Zk26GMz3rjeqt6ie0
MfhUlfoWMc4Q43Xxldb+BQzOkfSJpdUcpCLe25kVLFvzmcAIJzIfuwzABdiSBjdrFnuTtcPWNpNG
JUFHQmDvtDXLRrsYMz7Em4TYJeg3x7ClHWcLxG+TVrYsYKU1ZVtunoQU7YI4IiE9+3JF/IGyAA6s
dthlf50mFjcmatGUHIpBZt2l1v4r5At5W6jQQCSSEeAHHntDv4f1+MUTONs5jfoi3kyGc2gkCjuM
FCRpFhIOBhU5LKEneBinWXO1MXEj0b7VJ0M5DGP8AegGtrCUuW2CekFeq+zebnP3VF63lu0DEgaO
R0sws1baF56wDcMdmZyxacWrdjaKPSCMva0SIFDUcpsK4oTRZRFVgxTC732HQRp7U8cdApOzq+uY
2d2oEb9oUXq+nQNdKdVi4Ain73ksRdKSka2ZDzENBwG/7aQUTWjpYip4wq3H++48m/ceY/3grigs
HndspZNgnr69O6tnS8bya0hOFlp3/fUzijwtgug4tGb/6SVUVzvqOAMhb6wG4kb4JJnLmYI5MmPO
13Z8uMvfPEA4aK5ANJc6VXv+pKK2V8DU9p0uemEmXrUSKDgA26hvB6Nd+7urUjau5zkVYvYdTWZE
rm8Y2+FJhrfV0fRZ0XO7h6iW1oFd8m8c11nCK/D6xafA1GmerZSZFIuq7skKAvQdqBQsTF1h8TeH
BsdoFAvy0Y+XAgFTx6FE8gUMVR1mF1l0UbwvN/2woKaNxva0Py53Y9x04h8El2Lk4fInBSJvpSjY
hfbId4sLhIk9KtRCniSieG+X2wCtnMTXUQ7eTjWG/gLUkE1UO98bh4rVUkbU/OkQwO6HXMFWcn8k
sm6jFexz7R0ycOy6sC07kVBon5eNlkzuRdpzgIAGfJFCSAu41pixDrsNOwsQPLpGi/fNeMIXXAmB
FcjM3wT3Wr/1FyJPrC8+yFZbJYynV0LwqdXa5wIFvQGuG8V7KHlk07pE6wq4rzbuE461gHEWacKu
SyKkNT3KQxfy9GTIN3nvjhD1yQxpbQ+T4NxHJ9jMW6l4RB+A5agDX2xhlPz9vS5roKBzhV7K23IP
N5RL8JmL0NgNcyL2ftRahlHQDR/xY7eBxr8XrpdcNtf7yrEeHtMjD7Y+pcFtmBiGnDzakAcbJcCp
JmYun9krHfuqrIBRZxZmbTOvTM2Z/1Xr3qLT3n8cpalx9zGWfoyAb9UeN3kHchUJMw6STK0IHvW1
3ssQ2V2g8YcCrASnWM48FuF9Z3Nh9yJwFLadnHnrDwzlDx7IY5B8PevIk0ofz/DJsO+cu9Rpl1K+
PDX/He3ORXuIOh21w2ZSABOVRXpgKOy2gBYkc6dU3qhWGycxSG685iveoSaOa6RkwXh6h4lxo8/v
/6P++p5/UWKI0NoVhpqWvNlwXe00nfVn01iM08psD3qDzusRRfcKmEhd38JhTuCDVjzH+abFVvxI
LE4ukqaboyEi0eZ0RGRIt+d6ZkWmjvnoLDMbZb7NCJasG/n2PqTsaGlqcxRby7v/KaY4IXU1ScNT
ohfpxnEHhtXH3ipsXJfCkeGEa8eef0xZFrAH27ZOJmlq5xQy7ytESXB9cq1SM1U9grX0JKfIFP0k
SObVO7NTobdMEiPt8LatRliyEJ3SKw/yYQm5DhtnQks1tu+kvgK5gRdc3hTgmR8W/vJIx2lV4wkG
j8hl9tLjB4deVvx5kMkVauWRvO1zYvO3hTrn7uxz6TXtAe1dTULAmo82Lw64N0S/7VIClk6RcJJp
Bexccq3gtV94fiD1yXQtHzJrhP4HNN9O9ogPzK7H5XDNUT8tNfULVL4HUdQXKZquwUd4hPxY853A
+0Pe/Jd4EiOR/5tRYWzu7OMIXCrei+CaWGxR9k49hlGpvSM8xEo5imWjzv217iUZ96qtImTZD4rb
bh7znpTmp/Jb8WxTRBRgQ/Ru0rzHzjRtpI2RYrREYTmDCY4PKqv4KJ1T/CyNtXWOjkW/QJbS/7FH
R4w15iaGCIg/QEd3lOMNvip+uzY4p39tfRJWr3P3sH00TkSl0utLg0vKqnkXNGwgvAqdDf7yLNlx
tNsKkh5pQo/UsqERy6d0UOkw6A6kt968kPcZPpOYxNRrS6zHfzTZxtyVkeQjxRgtJZvtG6wrwbWd
+hYiKNiDtLha1CwCeeyy9lszxdfHxyqTRuTRwSPP+1/wWGoJTDXOU8iYiFzniW4ocR5u4J1WUUiY
X57SbsqwzvA4UL3ZS6RWULt/eMT/5vwDVpGr8tMbrrqVpUQigV/09JF4PH4eOF2oimRdshoFTh3h
nzAATEOeJ6V/8Jpwf84Z4p0hsqqnW/QLUGTrAEap2CCk+uynIFStTIbcCn7faYr4y1N/c2HG2JXr
cVMTJbldSaJnSa0K6DW/g2WRnrZ0EPwhGiuXZ7Bu3TJKZPbcsuXO349AuHh1JfQTyh/jvqzsifJW
TwlU4t/C022X4vKmbHHvV4WfJx3YEuSXbKwhPws7tpypNLS/AFs1eVpCOh/jpdZMrSqMtvScvSuC
wmvfdqb9ZO9aoqDlMqu3JtDBUvHg8WA+x7SL+/Zn3bxGYkldFASQ3Gb2njJ3qkTpJBF0NoNZxGt1
ozjmu3Otm1zTLO7ixSoVMr+piMwnySvI+3abc9264Byo5DFi2/SFVOYRCyaxmEyPvMYpCxvWMiqx
7rzya2Mvrfx1geM/20AjWocKDfnp9xsLpfPY1iSSetZZorPecSOSlmty7rY7CLzo+0UvujeS+LkP
Riu+gCmLu0fcAJ1XB4YoFFhVnJfKhTTdkEvu1zzLKGkufHJZ3dM48/fEv9/OnFgILJ5CuonmyAfo
i9K/wQ4ZtWK938hEMevlvFC9ww19JTRx2Hw1etryR4RoECl6McsucZJ3RGw0ii9JN6ucuk0FBlya
hI7p7nvyyp25ynFmHw7LvPTan1LaieHQXmpOvT8dJxlpz4VKWPlgaXBn0w9O6DbODi4gD/YhlYbq
cpBia/mpSHa9jN3LNrkJTYEfQaQ68ZMyX3twvMjCDzPU7VwFqxouTVHJf4ZmMUE61nH5WEuGlkI2
cDiQ8tnYn0wDUYkOBrgtEQyJZs0Ys8XALppNeLVjwfBQF7idfxlVMFoSFfm1DJAc2uEkgw+vWbJu
vM3y+GlOJOlSWFia/kxk30LWO2clHMG9cYhaxbQJL09KDzTG5csw7dlTuHUAthJvYhwFY4KVZUss
5Ew06E9jliVg43WuYDhiy1ewj3sHZlerJeoW1h+54N5VLnr03ALi8wux1/3rxJfaVe/gvp3pjezd
ly7yf+HT1mMnXtOHuvPUmOWIc2YfN8JMV31Ki4Q9Obht2ao/0xdcozN1GNu3umb+jnYue3X9z3hH
JQE4DVjn3HZClYgg61EF+9QFceMF/XB5+FxfQXTZby3PqFUSauw0t6IpIMhpHlgwMvsdo6X43Poj
9bENJDFffa0DnYLJCMAl9WGm2V5IYg6YxN1fypTAaG4R6tE7wOWvnyp3Lq0g9u/4rvT3OyeDhNYh
yXz6sf0MfwUJagSpWwZvBp8Vd/VCY9+6VCEAJLgLFoVaBeoZAV9egGJjjW/WsFeByEKi9/nwy/uO
JNQv7TJU7/6YG8MZSh9QhlDGjEHCUlVg8lq19ZgCqhjuhr43qz1JpwXU1cFcZHlO44PzPTjAIrF1
rI62cpsGdVIETZmlYs+GS9ERHJT8XmnuDgzQF16U4TC1+40iiibcq0QI8lzsKM0A+AUNASJD9K+0
CUnST0rfViJIREYWi9kGoUPlkJei3bPLB4JSTUVO27cw9JiTbDCle40tN+qOsMX/19Sfb2oPjoRB
3qfsLGpoDfuHoBQoz2WpyFQC4u5F3iF4tjnd+RvPLEUwedaDPMiY4ie9ckUkuDk2BWmYpNyuDBlR
PprlBI+gy0Ig1R37I3JEccU+iciipF77wioNRC8OS4T3lpADinO/JjggrKEJvSuip0qhGGOTL39d
idtNTqWZ6+ZayeAxImbDYwPbxxmk95I9kRPIxtqpf0pAOpVdRsCy4jCK7Tq0vlGj/V8F+k0+fsOP
QvteYaUMoCbooJJhWexj8MpOWud0o5dKiRYSlgS60vQH5gVUyKpFNyfxGgpqV7fy7GLvv3J7ZC5h
T2Ii7yie1NIAr+FaMf04Kh7tKI277pN/YT7GoOB4ySUXXD0mGxyF6ukRh/Vhh2kkoIJMWx3Qd2uS
P8tqyfS7GcFrxw+AsQubyB66osq6iETjzXz4zGOe2w99WIFQBWSy0VogiPxRrhtCv6ic1qTrW9BZ
ce814w/CeMhMp5bZGWA1sspUs9eKCR593GE6/JSLG1vj0XE+wsG1Q+zLCp+YmEuBLolh3tSoG6hY
Hxz/KBYVxJokppf07Q7cyokvkRSPEJvUXwG23UxzkWplumBq3l2eYQZLjMvzMfX9xs+G/V+tNNxN
AJyYL+WJrK1P+aQP+nacsUJuQmuuHCAd+YcUT83wQmRC67FWDOmNn5xF/mJJ3JcjR6nZdFVu3fze
D1nz3i9qR0okKg77OpG5fqsU+VTe647SKMzq18B7OOef90jZDUwUg4bAbPRifMjccqIWbZtTIkRn
avNQmOJwXoi+H4JIFirvRMIf6+SjUuQwqVWWwJaDWryzA6Rnuc8CyNThPKo9bhEFxdqH3XDzNn1z
z34PgChkIm6ktqQ6pCqSMrsW
`protect end_protected

