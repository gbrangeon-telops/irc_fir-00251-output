

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
bvOwtDo+u1XQuHmmirIW0G1Eep8h4q1lu6sagQVNOpqoo1dUL25zlZCKWpryXBrbavlsSVZj+/Kj
u5U6Rqq3pA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
R8VeuF45EN20zhkGmJksRGl35KTSV0YbXBmOJfN53AFOKNxf64co0R3kMl1KH48vuem/BXWPzNwW
17k9On+EP4ryAUZ6V1YvtlO9Er2xv4nZefuEO+pELxS67R6s3b0HhdPIKa2fxDF3e7AwjfjDxMiG
HOQbqK01rVOmqe+2yps=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
qqYTedtVydnDu0uy4wgVS9xnI5W4e3CBu2tom9I4ji9x6Du0u8YzLw4sHBXlBjTr0CIBWi+453uv
6i+HBaHUw6WLmgP+uD0PvRoMp9iMm4rcTjCZCtUo+5bxaKDQQyKy3VozWJN9cYsOEXUyn41sbHk0
MfnFQ231FTzHKrD8+sW8iXzJhrvAxVZSOCQNc8FKSuvFHDKgrQOZi/Dde7fskgmy7Y+pQzZQUv6h
7xsxzMyVpdCwJjhjdow/xj17Fc+yTtNKSxkHMIxVK6RXkbOidb7jBkIw+8aEzlqsG5f5vpboGqLH
6uQ8IqqBeKv3BDowwIwUDotWgCgTdyFmv35LwA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
xgoCG0tChkhv+ljdCxpV0I73D5nOgliZqF/G39R6pkQNEQixpt7jSEz4sP4s78dR6d8BiB9A3KNg
s8gNghB9SqKmhRG0Jvm/hSIBQCWAqWOwg26IvTnT3j3MalMVsj1r5WE9uyiqdJ+QCTo/Y58NBx8l
pM5ABblrTJM59LnIcqI=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
VTcA7V7opij8+vJ+tjjgJGiOJ+o6V1u444VHa/k01STvZB7T6/Ztq4KXHSVmD+driESiC+2EQRes
dfVcUifCMaPU4kNZrlpS+Cz6GGzKHuujVBDhNOZum+ncGM2VGmayYd6F9EbhwKFTOVOkQmEz/eFL
4IAryyIE59LghhLnEgKJ/yOFNS6XwipLZ1ztAAj7QDruS/h8wJcmBcjwC4vXftAO79YXKmVgRKly
SlrrXAPgfawAm5V0hj7SI23oHUFrT671NQiN+jfhZylivDC/aANQXHsoSuY7NkiKvHESuXKmJ3iX
cfk8aGjoqSspgWZUBuwV9vfaTHDt+AtBbt97TQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 174368)
`protect data_block
xm01eJIByOWVGUTkrA9Qm/guCRv6SLthlJtWkIb0ICjBJ25qm88gtc+SeEeehXgSQu5Vym3fJupQ
aiaANi/cChy60rga+3nsNr15rir+9XYy25KG+aSG0ivwk+csYPUOq69EtA2wMVAitEPHO5SoNqJN
S+czPrbe7ypMWnPWCEEiQlXAHURcFdb9WA59dswhv458wIXocuPqv/5XZd3RZXRE0LBIemfXw6Yk
X/H6yE172tWfQenji0ULd12Efg78xVM/8MLA5BwHjo7RINNBKHMaGg4mz/xpqYkYbRDK8Jxr2v1r
LFXvb/21Qrxj/jCBrd3AeJXE0Gll7kiqh90llaM3dbmatkCw95Pu+NR+3xASG0zCRpLuW71VLKDI
UPBmaZnrJT2rCXtXLYFZKoXGPtbraC3JIh/heNP+nM5pLcEXF1rmY4PSYOnDt0ocmW8v7efRGBue
zdCpzv7FjL3H10FlO7SFf2OLybnQE5ZiTVkH4pSc4Rof9aL1sB/j1777Z6jZQPwxzpiERRjQwnf9
3jjWifls6OFjgr0esrzIhAXv8m+J9CXATeHdNq42gxpoRXKYyco6bXHB6+lEzQrMdXbADzH15gZQ
8NnfKo1BX4rBPtPOUI3xoRXPWfC97LGh/TkZn8wrjYohYdUZL1WQHglr6Kb+3/qBLr8AOgiQ/b46
BtkhuNxcWeNjDTTf8keIc4ZL/6RHcoE2VwP6nbhfzpxVD0ZiSFp26q287wK6H8JMGNSKSRdZA7Dt
ihbpkiLLdc+BfKKxUbebrz65xbWxP/bByq70riYPlt0kEV13hQdicm7KCMyrX7cH8dnVxESAnMBS
ijNN9LUxQZLWeNhdTBpYlUlns/rNhUoRJcvVRk+1Z7udwhf5YerkeMwlBQ78g/v0McN9Omwkc5Ax
HpwGy7a2+amFID/eyA/04GifVwcdqEhX/QEj0aVL8Dm5jGxkH98BXrW+OK4i39uvXbhk0vm9kxxf
tDHwx4GSCnEd7c0oZOL3Y0Gl0rh5PLLNZ9l54H/nOIyyMR/A19WiNcwM6yWa6pBCScnM2qMFRG5w
lh3qv0/LNue2TSp+kAReIIlHJiYpwPNXKF/CcQgKb0/SdRfpHLdSOJgADqVohAe4kuOQRqwp7CgQ
IgR3c+iM0u7yuA9XmxHBWUvmciyDDjmd/Shdad4ftmEUBVXdxUv6a6v4fMWHmI+w2n14t95/stVl
TqKNJVJ3OSpnTMes41OYLdzNmtd43vbCyFShXGeZ08vHYRUC4HAeqHvCR13Dzs7n5XiVBeaakFG4
KyjZ1ez9aqjFxbAgLSruV/0MobbzesYiQvcoJ3Bgz8nkQkX5Dr2+mmN8+ldb2k1d7mbL/T8qDPVg
sE7GDXQub5p//GoEHxSLoulOZMRMEM5e3SRahG+ElfrdEe8phJAm9zYKQkKS/og9W1JuEd8N+uvc
xjG24Es8EJK16qEP7XnkiaeQpB6lZxOpozjoj5hu0YLsSIM0MWCoAB569XdbXwDoi3yAReR0IwzX
XsDkLaV8JkcRntwK6i+BJIyUVIuHur1zFQWYyF8UmcUbiuhCZzHrFMvZitWw3XrPcq8StTsjy0Sl
VXz+QyhFM1AeuJSy3J7JlpvCe6gjYqEI0mgZhEzSOT/qayzYBs4KNvTGAo+wqIqhNclsJ7D+1uQ1
TTgknhGSfomZV51E8yp6TuoMMHgUkdwUpOfqhpA6dk83H2bp5yiGy2uo3kN981D/hUb8oKMzme9C
xP9HvOzU/+99o+M8Q89guJNq7BD1TBd7fhye8z3Ox8O3Bptvh96dnyU1pJGQ0vwrsZKZXYHl4WXg
+I86cmAdyK3lflk/QtVHXRQNYWUR8tWXU7pkohSVU9aUoyZsLiWyx3CoAcT1bwE4bBJbhn0heAIp
vkMvyb9crpvcNGAUiRmQcWFZVjTDr1JsB6P4nbTSWT6a+mdUfS3cEcfpd7lqaCDsXOjTz/ViQK38
j++cwr9dZHu69Sf1fiNYjGQwE042Pu+8k285X2Po9WhGRibZY5aUDk9mFCxNPy2j/CNcCv+7wsNz
Cll6biv7n59Fenvpw35SkN411DLgzmj57UszGVufw4DdlSgvYA+G2OaE1BtpaceGAe5ZpKIGhEdL
unwqsxZ+VoCCPNjLh77MZgxBoE7Aefme/8Iu7th0ZI2S4Yt00JRuXjxjRhaDgGvExN4618j4Rakg
/vSY3/JYnpsrIL+MsWxQn6h/o0XgTFaULQztd3otZ0foWw1L+Jzo9nxT9lNNloSVFf9gMdboI0s+
TBhmswXDhE4DiB/jVULwzutmVRXoThSnqEAw5R9L6HzLXqKODE7nf7Dq56jBmEnAzUtd+XqTTqwD
4oc7N/TPaTYtnXhInIiuT8zzkpfLvd8i5PMavsaQdXx1HQZ8FucxsowalT1MR6A3mjQwY4GNmgYY
YAwpqot0oNdoOyCilUZ5/DgaCi6eqI002DN9AytEhukWYYp02QPnDG7MvpAgIFQvaPnS95zuIxiK
P0+X27hRYapb76sYFzrYxnpGasAmCEXefL/vMcdghLiBq4etjjFR5tR2eo+4mvlbCGAD94mGfWId
sZKRfs0Xdlb5q9qdFqfIQb+uevzNSdIb30ffMKd4R9o6FwLZW155lT+Fj/gqqkD1L0mDWAdGtbKr
I3nf8dcyMbzktmwwqK0I2ueW8Rzcujn7UMqg0hDxsXLZ8hcSAK9IxKFtyEVxUwjH24aZpfBnYtSp
V98oEp6da30vzcKKxtBtm3r60YgiTT/BUkR7DcLm9uopZbFnAzHS9kOQ9frnqtWHwdyjpBNhi/1W
ppj3zg8316448qk7nXZJVnb5O+ymbNWJDA5PVvYSKRXIObVevWhq1CsUN1dEWM9HtNVY4HEnNOqn
YkPAY0JJyzhvG8RrsdRd+3fqQvUtBOBvDUCnbDsv/jMmmyo0AOFtzbuQw8ZvHbz6H7A01q/41RM9
dJ44XJarugjTriff3iGnYpW3/Y8evUeb3G/7+4dtECZonojYEosOO6kxG+iX2DQA7VvXKYCpzkDG
Q4y7Zif/FtmB58Sime5wkd4p+6Pss6gpeKdn48MRhNWSxB8hdR/e2tQACyKwN7Pxn3ch9GQPNlrj
NIMm0FYTJfmJ7PDxgg81dVx55ZNbF1/akzSDzn83z49C7mg2bNtVF6USEzxb7q9OyFKQ1epL7hJR
3lFK0nnr15l2qaTIfKdzSCmNIqupLWz6E1xQVmD7SrHCBvWNiVw0hIna38CxK1b2UMda5x8nMgF+
uC97UpsnKaGWKm15te+dTAgzln4jJsnrwKjAVovD3LEXaQJudj2gzd+Pbqnruet94OVpEb7su19p
URVshphEKei8IeQr0VQCMlmxRMgKzLLSIjka8NyhOIK+7Q+ZAz8dxUoGQW+zBHxtNIjmfCPEgnwU
tJPmAM2Gpvi6llDoU4xDEDxbwk0htK/I+u4AKfb5M0b8t8EL86DNrn/yxf/5cgTETVYi2oOMZxWp
Vyb7F+21VMZ8YANsfXIdmk0CAXzp3GK3k8II3VzcZ6mAWPiT5W8RXNY7S9UeOJDr4rpGc/eF6y8/
Z/o/trGIjiOGlQo8Fn3poDQuaMS/rTombhr7M0M9qlGc7LEzDpmPBXbXdZ4J9dvHfTmNvIDmjvdX
iB5hm3oOfVckd3ognAqxe/t/GFAWwJ1wgSTmGZ9c/H0aAxFqGBlPjkM5vj6eTLkgttMsLBtv3abq
gOtX6UVs26V9/nF8JK1PkDexjr2Qkt/y0eKrqHfXEIvVPemO+6C8drG8QcaJ84HCTatJRts+4cIW
pjwCR56rPxkRjilojgyTMFkmsHPs6In4wS9GIeKXkv12P7fryO+9yPfDyol0RE+ZgkLakal+vXpu
bEONqOc2bnjehjkRSc7pJmNzLFLDmdyXF1ZcMpvi7uxs0UYSZF0F8Cpwcpq+psWmdgnbCQGK0ywM
UP+etgSXhbl5elojgV6mH0qR7DkAeNejKS81v1rxFx6xj+gGHPQ1bHGAPLJIvj3zCZvyjnDxXKLl
vlff7JVa7QxWhHJkWqIOiUhGsOA8uPzmyvVSG8X2f2ngr/NluA7Jcxo6pVqHA3QRngNqsG5VunW/
GilunRNOHfhTIgnvxFEBo85zspeJXhGC4rGUcUlpBDd+s95DQRpZjytJDf5za72OD/SeYTGuRYca
K4BPN+wlwV66lIYvcG+m0x8CA/2AfsOSjfLfzyACbryyZGpjht4FE9mEGGjRRW7ZjAyNBVUJXGNo
Q3b0I/Uy+oHfbjqbNzxl8m1vNW2ON4NhyxvnomnemO4tOyn37USg0HSWiiUS+IQLvlRGRsogpHGF
l+89ZTW4BM0X1ygrMKHYHHCszkL47qRBEvcm8DKaTny9/SCVSzkNxEVxVh9NYahEDlX6aNCvp+Iz
ZoFUmCoDxJxK4PmjwWiU02qJdYckPQUGOe8FipURK9RgilsOpjVBZK32slp+sJgO1o1qirwy3347
gYLD0HbxoQd+T+aqU8anSTuLtrBlwf9wAMS7YtFWKIFF9cBH2wenPzU5+BFhGKo5yvkUqqLPkOgN
YSHHw3Dr5zcCNBEONzJozAwDTOj8PzM5jQVMXkE7HJgkYNhIhusuhV4r4r2d/Lmv98hDjwkvo/YA
oAuTrp7tEseUP1hT0m5NvZjzgfRghqPTesG12tq5d1b3jsxUveZQ9Be7NYOMTTBkooolt79V0/Ju
VPIIYw1JSXhJb+hoU74zyCHDa4a39AdqfPyndt9qoTagMFlTUlhBGgZOo8C3wGNBpL/RrS9O7wZ7
bIgUirgVxkPs0ovDj0odxzDmmICJ4oKpomEApkb5Z59F5Si97OzAiVjTzYNRvdcYdRnDToR0n36U
465/wfIlkJWzqXM9mHiJYYTlSz8QIh97dTofoatexvYJjRHXBdYxYa3Wqu3jtgMOTL9caXMkhkzT
Jg4GO0p5qjCse8AVv/6foPzMCiIitEztxyTYTl0iZHjo/HbmpIf7Waj4TsW9iz/viOSrX4JhmDHt
kNItWJGVWsw0J2Ek6f6zc/X1g0XyePbasKFXKJ8/fANkSg6dn4q2hzLGc5jRdJLOQNpN6W1+JECJ
U2AxVHhvZYllWqFDC2Us5yY58b37SXnnfAnqxqqhqQ9XGn/As/VtvySFmNDsl2EiLRdaov8mSRtN
Tb60ZG338JXTDMhlqKG0imYm7L95/sLUqKaqsr2IxinHcSFqQzbT/BJOR3tRRBgU+RMj7kCY1CZZ
fckNjlkOVIX7kV6FEmY/WJv/U/Nd7vsHtdEXK1VGOObXW+z12rpyom5LI/gSvWovMPsYB99nlNk6
pyP07/x4JAA7WqtxwEw3CiS6f6CP3eyaJiXcMWydNZbDvHLRGggmwqXsLfpibtzNwhDS09Z2yVeo
X4LI0d9bOqSbAfSHe9vnbmQTDwalRvOkz3PrQdy/zc7ylvhcUKoqLJgxcvDF1lQkRTzZMWUnIM0Q
hiNGsVtTP0733DX3DDUhF7hH8AyTMoTXHTf+VuPpXySAHRNq0qKTFn+gNnHGJUA2JJ3dUgIf2CSz
8bCvsPjPm9LqVB4PoGL/J6jvC/W3HJcKC16AWFfPDfX6Qq+VICXVS2fZ+XIaw3L5dEMBWmJoP2Vw
/UhCdCNcdye5/EK6hfW87ePuTiJrVzZDm+i1JaAQk9NRobzsdkoH6BqCmd7ACux5M5jC6g3Y3LW1
M//rOqnGeGsqzRTdPc3ZnXpFIo1gUQ4q/Z3mLVUFp2Cp//OwOTcT1qzogvIlX40vXjBS9vsYkpM4
uCLcDrHNmN6XCRHBF6Z9rtuemLV0ayD8ZJqtOCC8l2MMRnJlHLmAU+cfvmoK5cqjP7hTCuXa+aJK
BySAqO95DzGqVlHdBtWgIAeefMiaCuEnCBaZqtVtSkUCYyA4i1A+7A5vcamyxUfWPyg4+mx4Dea1
7QNEAwUYJW72OalUndxwXTyRlcS5wwBkvKurSbXwUnhDcDUxmwpCHtRTFk3WJ1oblGGZVfdkq6Vs
GaO+xE0mN4w9RhpzTBi1LdrPy9mtzm6pT1Iruoo5IrXnxSGs3gT/8jFzUADDHePklXzoLetqzmhn
TfPSrQz28l/d1wOHtxNI4dorquhZuFfCNCGOSG3JsM7Pvz1QC8tH6kkq8cIWvhNcyUvBxMlkwcs/
4KgxXBhabOHBakWJMRpAP+BtodTo8ZcWL+EaSbpY/s+dHg0XXqPe4M4RnUwmtQocFChzKdGQus7S
uy6+Bj60nh7JbmQNYyVQqlqUypU6lRomAI9emtmDwFi0SsdxNao3Lt7DH2yLJIeakCgEJYC/uXM+
JlJb8K4/Ft1SRalj1uYceoUhMIKrVV1oqQyNjgzwLza0N37jrcVINEOlLxrON759CtPVQeM1GRx2
bJvlj6G367dXtrYi1/KyBzoiQedHlkH8Ob1R7Ywo0CTNtDDlhaEPkXNxpogmxiyCPtyrKsLeoVrI
e5lELMQ5jTRsOD1uCE2RowUTTScr9ntrHZ/EdEvbtHhR2DRf9j+ohh/zHZr4JpWDqsdZnIyLybkb
jMeYd4MxB3ERk9AYnFusMgraRO+06eRhVN+xLAHp7dvOb36r2TG9+FKUDBPE93tlFjn8acJ7I0Fu
KhjOZv1CenCJkcE+pubFDNnWOuPT8QmMzre82eXg+Z6daOSzz83SFrlP7o8xIyeE7E+JnUvhazzS
+582wm1cZTy22atE2BqmpbktAqNWSt4NwuNrA8ZQJyal5oTLinrKqy+xMwYPbS84OiqNAY1F/z6L
B9WTArwRwcHzP48RNQhniCjpG5HopWIXrZ4WXi8Fsj3fv3f7blcfv6lEZ2W765KbKP9swCmRaW7J
6CCsOoumuZn8HvoUwH1UE8amyQBPDIgpSuzF5kguki6eJygPo3n2q6RpP46JlnRDqB0CtK+xaBC1
sFtK7v7v+LZezDx8HcUs0QKZdk+MqZFiTPSpYnccpUysbKl0gweZBlRVV/+KOcOI9SM1eO9Zs5kB
2lgALalb3fnK9+OzRsLt0x/uVH36LvCgDiV/rO+L5PTuB3oTB7RzacGU8w6YgvepSg3Y1cDRnV8U
ruyWsJmyTlmy18P36+w5DLtmJZ8w0m76InToRaZTvAp2/mL7umsfcNwQvPTa35DkY5xRGjpbvjpe
Jxa4c7w1RR68GdzX/Vnu6mmSq164Y/4uHiMyEkLrBezcLZX31RKLmLaq3D//aYNcfbNOGSrnm/re
O+mysrg+NOuPqOJR/bE+eCB3cuJVSawq0YdWmyr+9YjoUnZlXCn2+l3giTVG5N7V243z7EuJmVjx
hV0NqDlo2t470ihMOcGECQb9njQuH87LXgaPH8V9QwOwp8HFWHFqRxRKv4xgdf/GjpTHqEsbTYxL
nIUmTueYG9KywUBNOZmXiKvg0pxvcvJLhdc7CqSovGBo05UvkXd/o+eHzzU55eZ2gXpMCAvXFwS/
WVcOmNq2QFSo5FzONDJXnpA/mUn3CUjkEYSfQeDqLsbMAv5UC0w7rEiWilqGUalYU9Yjv6K7biBf
aLBpofIj1aJ3opTUdV334vKWMecmou7KvTMAnoIkoZpbiSAi4lwQgtLFx/hElnQbbqFST7qifXVW
98UmLAQcDYo2Jo7oln/mvDoTt8lnoNjkkoNI9ae4i/2TepJaAp8rnv5MZEaNmoZBsryx9eLgjRAp
SjptHcpDXWoxcIbPfAMzj5DXdlOMYW+aPlLcsbun78MgEEIJ0vOk1yn3LpSmKKzxBsWiW2BHzNDB
ZEIbvkfOvqugu+cxuZaRp6xh5JNQDhu7SpvEr3hblB/czNNoIgjjftXTJB+iiImf/aK70k89T5V7
6DgbJ0XY0LOydfoVWxeRVVS8nCm1amslcPPx5QhJy5JEKDR52LctmH4VZT8AN80pK0ZdZz2bWxLM
M+NRAImoOxzTNzvb8NafeMJFJU/tAc8vXwz/RkC3cR4qNXPBDKk7x0VLVZoWmu8uROs/EFnS95Pb
9DhwS3/BiGVflTeS1OKh1iZCoNMgKZcjW5biMDukXLyXrEXHqjVj9F2zQHwThXgl39+hUi5QIUXi
6TBY6qVCZeGXKShS0lei3cfVlgWM5TEnR8FNZpsakzdfe+xCfwQXEG8Dfn/ZqgF3ZUoJY7IvPdfL
VcctmqFRMJ+zqUaN2MJGVlVE/9jM+w75sj/mXWr4zPYKh/waXuxD64zXvUYxtAQkVPqfNhZWgclD
BvmZHYy1TbczoBx0qBlXVcNpzPzru+l8g/K98L9E+cstc6AuHP84EY3ELFN25zgL4vEQLK3DPPrY
gcDLPCBMW16ZCnSDrMI+TPSzb0+jU3AfZRkubfJsAKp+CP+WtIqHZQ3twxuPeBKdKfJFpCqDuWcU
Hc6fAs0Z+2ZPNri+jDeNfj2Wla2YrhIoqAhHX8O4W03OaE46lE6OaKjPhD3VDqOFPm7AY+/SiXGT
FN71AROgGUBG/8NZGoy/luHccoDLy3Sg3TtggKA+h9EsLbuy314XRD6XubO4jiVeQZCY1PIv0CYs
Dg2YPF8hDFtuYqVrMNt5yCYcIor4FiY0Ph8qxX+/pmw/OKzt8FLVjK/MLjrXKoJ+JtY1rZEUjCRG
H9bGw7U5qsRIPIAPzK8Q8ptm8IvjlU1FZtSewkqQOzDTaXypZ43fr0cFmjrI0oLdllnvhw7vAhuS
euz0Pk/rS3kQn37mk0Ckytndnxo0vt5AnniCrCUUshzOCPHYPCKiWmFgzBcl03XhZiEJ0ifCcSRU
C4QOj2YZvNr4RpeCcQBjJh9oIqySTxsaBcysK8F04444+2MdGYm0A3O03EtB/Pd0S0BTxFUhFDzF
/VuoQhJWxpOYU7FlSnSghvD/DTMH1fiFPKSHF0TzOD9QYnUL1hayLgD7CZEOtjxyQ30L1zwpdN2T
ZWR213zxTDLpTdndxLXxvIxzpmZu85ALkRolbtpb2hi7x6uAjyzpMlXNkZnx1ZGGzzPfZFJkU8xF
Anq7q6XCpmCkqB3fScrIEsb8Kq5Mf7enV9rwCMutHAckyKO//wZfD80jhV47URMWWvHXE/TnDGMC
i5lc7iS2Fuv++13GAHUjnr/wiKX5l32+UuRWGw3vLob/K8Nydrgp556RKZuGtgYvIHPGCX/7Zodl
z9byFRKCTkDmX9fSft1VMYUA/BF83kcG225ew6z3omYTxGW3IBD9FhgQ1WAmU4qro2dwcYN05Sqv
wmVmZQXTkINvqrxTHJ/bCRBvKFfkhwZPE4emwBbQymEa+qWS93kpdwY4A24pbFOPprTvoMwvnpCD
a+ImOu8eUJuTePwqgLZySd99dNIwN/sX/JBWhbtftfMqmd6zFyI3X39D1VJomDpVOMYja4PhUZa5
xzp6sQuUxj/HcQTbZ6XHC7IJy/QAykQp3pjrdrYcmL2aJDqa87gPg6O4cyI/sbZC/YELMriD3P5t
dFlOlAVZ1sjngsQ8RnGIaDo72zGproiLhxAukgCrkQlh7Kc/q7JdFOy1J4nA01jQ1NWNtOWHLYpG
4PYhMpIE6Ial5Y5/6iCro0umGW1X++PSczHSu78Vi1g8T73oNHX98tz8ZrdNYfONbADROA8lFNgz
fhxfmEHQvYN+GV8camsY4VUcMJoqoKSlQ2237bExDtDN67GLbgj8eOl5Y2AY8D5OKFEnryFQ1Keg
zCt2ymZCRbMwZQWdPL9yiYB3G9y56zUWeMMIJNBPMnRbIKXTMvPqZW7v7zOf4Nsddtw2JduBeK4P
WqqaTDa5Di21FnwR81XV1Ej/cRfKvK8lIcQgGt49mpHGozqagRYE7OJhrum/by0kWYg5LKSPNjkq
5/MQw2it9IemQwuUOaIICkVO8o6B+/veLf3ca6nIoFvz08j/0Zn653g113fRQ53HCLQgXiDQ7cIv
nrmRRQ7AuEsQ7Cy2aogtVaq9CE9dGqYzMeIYLL2Yh1HMi6Nrxb0IKZqDLZJqVq7TwTbLYdstsnlG
jCZ8NzQCSlXOiyMzwe5pdJT0qJPk2k5eWAFdHuJSRr4PVAvm2/VlNTT7AtnF+cS/IctUR1Q/Bp/q
f18fIf9yfNKxzA+KDepI30J5x/5HBEHK1jd6bIZ/tJ0UNUi+QGGnpVrGd1RWU2DV5Lxj2cS84rUX
9yCdE4gJGBMYIF1ek+uqp889uqJ2OtReZBXoxXYsrHf9XG9O9MmpMX2kmKsxJ67gDFticiXv3r0M
XoKAOVSYy/68s8sJRasCjdsMym1o9T+UcIlqOSB8hKRo1GNEtKXaD+W+BMBliEDOht2BVxzDqfqV
AvpjPy7vJWBvKQmbacTs8bU6Q79mJmsKVFZr1TiyIJPQ5FhNDMi0jRV/o+gCgFOw0gQ0WhsSO0D/
iYt6EE7dmAmbu5Oa0NX8edQy4gQ2oVoGf2XJavtDGBt1RZ5b1WF/gPgdTmFKtvVdcuRVmWhz3yHQ
4u1af20mcg+XkUzWw0DtZt6Tns96TlFFQaGoE5BOvX6dgwc8uclO/8DAkLvIFEWi8vLeXlXhQSSK
0lZ3AEjSky0/C1Ht9u18JzxCs3FIbceuJcWLsih6NymIncb/KyP+ZdDC5RyPcclIE36OzzppWnyn
PFkGGGI+3vgP7YQOjrZGzGIy14JhcttI7MLA+dydyYxtulqNVE1Nf418MazKf0UwjWlUYj+Os+G3
1+c+c1nviCbYeb1sw04cRl91/28+KqqSfTQI7Ej212af+S66j570FzmZZMXZeZfNviw/Mz32OcXG
XVKxG7hZepRzGgtOwQaPuhPLaxk9UALxygYfnd1hQzK4JKyVPoPmyixNUcAus7ExA53b0dNXwmVO
hDznXf/y2qmFdbcVYLLf5h2ouPKLNsHJvzSbyXGD2jLmBmi5nu/U6XBsX8V95WeKZeha0CarruE/
DU5mdM/JrxltIwPKfuVC04lU6Qrk5HtZscW2zoUiMM27Lxd1QJn0LPFLNzb9Gfh9/i3lIRLjnxfn
w2jflmr6B8I5Wov6xKne8rITmQ+Yw2lyRhK/SkLTX6wvw18OjqysDwvrdDmT0CjvRVuKIYkMCc4N
5VMHXpJg0uH/r201QN4Ac1Krx1Gx69oawhyyXJ4miOT+5fijzA4bAzj4PzpTA3N0lWe/vwHwAi26
lw7sX9FQt3e5+7fLFTWZIGpN0Py0QYh+wBJZiu1VKWq+WToktSxnF7MarR8pK9aun8i55wtYfn6Z
6pMgzP5DQeau8Ct1QOqPpVHTXq5nBGorr8UjZdHZU4LX85VUZH/namOjksuDrSc5aTLB9wBMUlbm
bl16j4RU3ewclmK8iAbyXRTt6xx/jz46rfJMt8Qz/r+BIxHaBRnGNANdZuPuoVkscPEQRlqQ4giR
kAvZc3ThlHcpb6Xs5Dw3GEKgJOe7xJaKypFiMVKdDJ+OhIa3lbCIBYYj/FBbZYeAfSAAElqQQkkH
We5ZHtfYCngW1IjTgaPbFepeWz5dPESdd/LtWFmzescgZwMA9yn18LzNjXX5/r7Azq4AKdYLjtDM
cXC4Y44ZVGYTJnlwrpAeTd0XItjV33Q5+S9d5S2DKDCMpQ9ZXcYcJaKf72yKNLzvBQROCQ9N1oFk
8I1M/vLc7GQ8tejxaw70yGtyV+eV9IBYg5oKOU29xgGYqBmWe3USwHqviS7dmUfaHO/FF3CshU/C
XkaHjsJQBBZaMPxjotnVaX/N637TARhsU+t41ZUiTHETcVcEPWxILhqkp4KBSWa4PH1GAHk/V0V/
LqXWQqmMTNRFbTPok0g0ToGbU1otOPSMFIFBOjyfX9ClW0PgUUDzqS8lcsEdwKyup+6cn1xZsWEN
q0EPWO7eiGlLdRyb+P1+pVLN9cCW4URynSSa/xgI1122n6LoqCaXZCjDVcrL/r2zoh0F4AyhEjuw
Ch6z4lenMQfuf63lrpU01S8yJKRgW/WdMUe8ku3WaNh1vP3OjaTSlYoAFCmbwReRMOT1XF56WzUe
he5T5lvDK5A1CWxBxsCpjwY9TPO2nbzwISzEsGKYsyXsJ6grJyfik1RPIzeMv2heWAvbW0iliDtl
GU2Pd70FwjgyobHkvxDm5nTVsaYGxqLAoGWC7VrZZw1edKAhzl5/JT0d+IqjxcXSyt2MzXUVYlZD
zjCYLSlgK7tyA/l1GWnqm3S3onfmFZifsPhTDQSu+2KDv0pU71y4bC5/rO1Dn4QTNoa91NCYd0NK
Wv5CTEpNJC+pcw6T1nv9tDtUmGQ05H02blnhMaslQ668WRUx8JSCm2WoCbKpDXJXSWhh2L0vKfWl
RAqjsuSLXvUokDILpDJF5nphewWYK6k9ngi+l7/kthAfP6zmgpgyfBuN5Ss8gNwH+Dj8vWrcdTAY
9DdvZdBtatiPqt9C+255POnLl4NM791OFHsAm9th4pJwl1gxwRlOreTQsuKDhIpq2n7y5NCWZjbb
EHBvr7caVBn/F5iUxofIRJoGBl75zJlwN0fPQN5IsaAIP5uXPeehP6lZwFIoUnpIjm6VP4qWRkX9
29FMnLroxdTaIRAqaWhCzSA7NASO14WP7FJv84yI9Q+Q4YM04EhxwtZE2Sy7uf6ToxpL2hgcZafN
nrxHUDvLFk5K7qwsQDq3YD+DLWjlF0rf470/F/TkKsHCQ+KpL9Q1OCXfru8JZk1TKxPMDzLv5x4l
Ef766IxnEJcN1/okIiebfxMo6oIwq9D1JucJjsO1+/5dXUbUolLpmmtY9fsBJ29DBR8GLH12tLqu
JnuXoBx9KNLohvPNTol/+hzdNtOm3Vdugcm3hRIQVeR/6dgHwlZAZOyVFcadNZ/CLGwX3s14uHQ8
pDJ9Icne1AadITGDCFeLgo9GqfzzcAeCGeAhpNJaP84mYbHmpJlrdo3MErjHqu0+nfj4CrQAq0rg
ECO1mjANPupA91IS9pVnqletQIOkNIvgYOf+WJHSXiwscBxPIpd1Z2a5PaK1yOc1Jz9TyehnUaMr
Yd1IttrkUa7MVIfFW42nWJmTj9ci5EhulE2R0rNrQjqAAFX9rs6omzfejJuyXXqVzOJZBvdgAWZV
cOF65HhYhpKXFyITvgjJsRqZTC7cBRaKEYix/ybughX7fMmCyq4yAcrUWM6mIPUigMrIYfdrOc9+
0FsTcn6deXXkfaoCBcQ6l3diNAlGZEWkPw+n4TPbZmQVII4UzWCwyczFDTOKkJhpaiqIHWhkcL6q
RTZULVA3/RVtHq0ade1cdd+bGQolnzCPUMNgDHjIRQaEzwRsPAOwOVpDGUXqG6z766VmqAfYoiHa
brwVxm17L5ReWOadUELYRPQK9lo7mr97KMrGUbl0ILLwNudJ9Ik4/sttDyzqmomgEP/+/uCpBaIb
SpVS8j87VgohlB8GxynSqXE28lK1QurPAmdj5a3PGYdomJY2CI3jWhaXiRUXdUccIiBz1N6lct4e
9hNpmjJVdD+yWrWN5l1V2toca5Ox+o19XFWsCVrB23vI+SeEbiYJJ5i3RiWt2vCBUjl3JpfAPFry
3rOGMRJdzYBK+lHOhz4a0WTQvn3IbLnDLbbkN+0xoYNM5vbV7sRL+E0P/aRQUSkJ+NPzS1//4Rvs
W5B5r3qD2cU6M+7kgNvro12SIajdfVHRQXSct7xx526aNDbTboxBmIKczsBlJZJxgB0J1pxpgoSk
rgrUrCetjWMJQTmEjSca0y2GtGTOpvLTL6ce9WXv0rWMDfqAUsqYeoQ4XaMJRrT0Rku4//EeEn9e
qknrNxg+nnZzaveJUKUAjoiblYl7qaYxQAddVFtpOa+bScmGpaRL8oUx5f7xE+HuZUgaIG0WN8yI
vt8MSkW8mmxTxNYA5YXoygP6XHP0ll65w4p7lhrn11fUe8WOl+KgO+N+vFIE/0eRwNeEUIKi7uMg
Zp+fefsjb2isr/aurul02LPDtY+5ebR+aPvUb6D/w/dbPiZPHk+cRrp2BdbhRTLl/ufRhvWUj4Yh
RMFX9aSQPGnhVVDSA1JhIgs+K3lfljDvDpKgiQkI2LSDlroeUFEUj5cx8QMKSmxY9pO6sVOsdUKP
Q3mTc/4tSe+MrkeiF7bB2LVCd8Opju5eXchw0dmRfTDMpEdsqOxA76pCyTIG3OuUz9BUbfDcG11Z
dhZWxBpYQ2twj6j235VnHjsq6jGp2y/tq1brifJOrGDhhODwdKSt5fh5TcEwZlyRVHW3FqGEjYoM
nEEL+yYATE6RNiO4I4Acp9x4VUyWIqNWyWD+H07P9WeD+0OqsNQuQKbFSdX/6yDsXea9gXmnFT+z
wSRj4KITrYvSyzx5oy21RdCHfIPyKxcklB5Pz3N9aQ9bAif/HXriLWA8fbr2/5IGxiVvHGcxWkLh
6DN7B7zDyf+cFNggqG/iNzI5O48xYen2gWw2OKM8BjR9ifgnvnDiyHcmEa/1LK/quA/BbOalqsN3
gvc5Se+ITpl68f3HTHWI58aTtf5UWgM/iKg5Lxjc/ddpR7U0R7dyLxW2cGao4g5EiOU7ZPqD8vmP
F7OrI+GuDj7Ew4Tz6+hplKjJuX35cYNeByC+ydus5dJZsat91yVF59Q63zzctr0VXYbjv+DY61Wu
r/KpzbHDMZnBm3UjgRB6Q/MRshuKBofEtLJblv0M2YwzFC9EisBNkGdK4LE9flhaHlaOI/zTj+0F
/EL2R1AGf/8Vw0pG1V2+4zp3I5i43yXibSlnPTUo5cZ22H4VjzqclgQPwHcZGI3Igo1FWpqFhdgi
IX4KMWDuq3AJiTUHJVD1qptWEASF5HTbtPFkRivJsymWAkS3xDE+a4TVYhXGSxjdbc/7pxk+hTLV
S/MEms1O5cGnrDr8kOZHJBnjs6pm8Z5vmLWjGXKGQJKb+74Rl/AkyoL/Q+XyeMqnMLd0pso+p1gZ
FA5jasFUU8O2jeKXKRNgBIWEWcjm/n/66VKH6o3FVuFkfJP+dtgeAOHPnYlKhS6Xml8p3SKv50tr
z+Ft9sJuWDeAxjuQ1E7WmBdrBFwzHzQc8DIDv13ukzV+XNrCzeycJiQMplu5iTeay57P6pYr0tqq
5Wa4YYHbOvLaxkdsbPkJuOO8z5eIBciaugKVx++5y7D8wa50L4e41eAZ3gkh0Bcup1AiFN/vhxlL
KbCF3QuS14OaND0I6jxuCnttFRAbTnhR/ymBdlBxe8kVZNldagBaEfi4HAkTUbbYBZ3ZWFfakIwr
oRoF+gz+dA00bjgQm5AhXDCzoAuOTXtLnPTEJrq0tMT1b8BCvhhIdaxE/Agxn2crTNV1w7BpDqU7
o/40IHrFNv76rwDBJ2nm7mlgnxXMqAYeuT/1BGoY6YOOfTOROuDB88a5NU5SPhp+o8w6jfC2hFjM
riMi2q5uUFQ8Lj+xh32RgAFfWNrerTXhIK+WBx0xyX/qJrnPwKcaISPspbp3OUdkb5dCwbh+Bb/D
E2CWT5ZbQWLPQzQydtCxJeTGP4kHWDPGIjCagBVD6D789yghPUCk8fsWvYGjukGCK6wpno8Zjbrl
K8t8nCorfkz/axTqVh54n5L7lgo7Gs6UnL3VJ16+qnFmsd8kWZxuxCt8mwNgkjNgMf2clIwBq4bx
I/NgFD29Rd6GGxk99+ZchMEb9t4xCp8NmiUNtwg5MCT//LjH5fNLrF3wyrrhtO3o+R8RYRirMfE2
K0XrogtsH3SiypySM8R98LxZF7O9Awh1FsgJEm/oVyq/TX4OifjHG4jlt6NmlrY3YtH7MX7Y1pgb
FHGmlG1KD1mzpDg25r4FlNSzFlb3nHDK7Opzhms45TcRpQtvZveTuO3iJpaqcWd1gNiPkXNn7LZ+
+pyeliadT4APzyQfAwTSAdl3TyNLU+ty44SeO7eEF3pxjFKKKBMyJUs8QTuUX3KGpriSYiJdQtC+
srYtJBaStpviC2tmJUoS8P3zGZGiJXZlalGHil57OpeU4DB5scIWIVXiBpFJf6xfGHl7NtlMuj3l
l2UwhfRlhxKafWL0Vo01fvboxM9JkK8XyjqhFStfpA3yydJ6ao+xYeS7BLQQqUTgncmyYAbsXUzZ
0XQJtmQJJ4A9cn/wZuSX97gKqIifu0AMKTwGe+gHrNLzG9n71hbiGPx5leHTd4XMBYC03+Wv1AX7
/sFywkx+0b7SQsXjBH7+tKAG1CJz6qCpAQ+Azi3SYY9yONn+rQf6+PZ6ipi8EL4s2Km1o+jEbUG2
sRQXiPz1pkojOLdBydQtNiFbEXthsQpr6G4rEnWRfT/sDroa93c9jMR/+E88w62VSydzD58n5Fhl
7t3z9dW3oWvxqtt1QGCMBFbuxWHe4WVcWHnWvYQvnkr01Mx/C66N17ifCt9HUxLAUImqN+AIDkDd
4K66uqQ8+weO6AxJ7Ebf9ffF5iUFRto7T0qWc6PGhit0h0k9cRKzYEIF9lNZynlVfQvHf/2aMw/B
th5yNO+4SI4ALp7KrRKkj99H/+0I08gq1swvWVq5uYUYR2iNzXdp5r0eTQyZJQQhsKAu5K3qnZCI
wrbqPDTSGJSoHid5/6SOdwi/WBRIjJZCH2UTegqTUFvrGeuiQAJfw4gt71fKrWIsQDBAmkSqtzBc
/BaJiATKlrdt9+lwIP/qYoWoN7i5rn6ghWPDm8YMqO4nGud+Q9fzv6dqyAm8iFlMpr51XyAxRr3b
uoVgNRCUIiUr8NzRkRAw0kFnQnChW4R2mhrDPwkIAxPV5bmbxmFcCkaJmo6G/XsupvuXJFyDoBdA
I+9lQoJPLvVE4Rh4uu79tcWNLpBbFtBqFnnxWBrrg0V66dj+Bk+Pq3/1kQBanIvlim7Iagx1neYk
j7+J37HKUCKXs/Djxe1DxSJnxT7Z2dUn7HMUNfU7aOmbNSPMQUkJ5wa0pKDxWkRgJrQ3gMzKkFSe
A4Q6T5/lS2sqfFNw4l3G7QMLFn5v7rK6d9JcbcTlPMFnoVLVCt7Lb9Ltn8i74U/3mgk6qISjMyLf
gUf5kXXd2lD/ZEOWkm5nzOLAIiz4AJWWixMnNKrucA2cBfqPHfKQx9f0Rv063IBEnYRlmfR8U8I8
aoprornJSaLr3Cit1h0oLyNfwsvmCeg/mZJZDcTiJqyr4LAqM//3+YAtiwyip3dyMekcf3tmwSCw
x40cus7O0iCwWgF3BJnocwNz/apJDA7JF4CekpjWcYJJ0H9RKShVgVsjekLJO872Zuka9pOv9U8d
8j1TODxL7LJ0Z6+eHgbpIqmhLbmLlyRs4VAdvvlbM8Y3PoCGaw6GnbfEvGqz4zzCBXXIAqyprCHr
+b+uNbT0nknV4vOydyVfbTe952ezlprkHrlArIy2qb5W3nECOroZGju1pB1bYTnIso6A47vRvMzz
CtOyWXeIPY3a4fPfsJwH4mwpFG3gMcYqUbqyDtveGPreIcVq7UJqYB/nUo74R9LSd5Pfl8f0L0vo
sjD3dciAHaEFbXJqDUWWzHs86Kh+6MxaBXcm3LEcXODm3cN3CwaWgOca5dqmOd1HjXSEAKcVRsU1
VKmp3gtL4g+6wKgUbsPsnnuzbMOpfRQPJhW/0ziVxJfNsAdgPxC4L6xnSYsDDO7Oqxj0pITNPG4l
APX9IFwYhCSN/rmuAPaJskA/hCF329wUco2UoH9WEqmqmYsYqzFZLgffQw/W7n0rNq0WL4K+inCt
8XawgydgZk6Ssa+nYRNwBvjZjy6VuisjXQi+JMFCaH8FOj8Fh3Hm6O1XsXMvVcD6lssA0r9ju7QT
0xtvt6dMqYP0y3PMWfEuxFJ3O/NWrNLeC3708bB9QvR2gUlgBTpXTVk+MxN7snH0fwf464AqVLF8
R0byrAfoxsToUZx50JKEU5PnooCVvj/JqjkIcSaL8FD7TjiRKyn9y0iMgT+RTTNZrK1871IvtjH4
o8iSzIW/ATD7j2VB/UXxJivgU/ZLwMbOmbjI22ISS7w0O3On2j8XFrkp0YONqnGGFWSPFkxxGtSq
CMqlH65DJVNtjNX4P1F4DnrxOp2/H/ybFeKA1kspJhLPQW/FczNXvRig2jSQKGFljCD6HpVpMGYN
S2s9MkLdBEJ6gQSyLDvWvEl1jGnRcQHcbfVXxkskt/vB3ooXJ/gd26rl9M9XX6NOgnR+yszsPKkG
zk3YkOPzkcLVmGg4DjvE7/ZfiCC3x+I1Lc6nye65t1pb173S+abqBML5MmohgXXw3uxUpkii9n9o
Z0RCJF9JR85NLyX8Re7rNOkwMimEyGd2qj3+lcUGqPElE/NmvwRYeYbKb51f9eM3JcWTDQh0my6+
kc8YvehOJ5uc6SpAULDvcx+6f7VncMK7Vb/RslGBq89ALzzM++YgFTab/kBdPLmZ4hFIZ99fkFSS
GEvjvcMmBqKUexu7sPQUP0Ltp9c0WhRW1YDWEO6sYNkxU8RaYVvqfk1HH397r96sy0HcYDc5au89
bTZSxZlKOM/jFHSsuHobhHnam1y6tBy/1fOYYGF7Y88GPrJ10MBQjUyM202LdCZ2jZDxrsZ/gdgo
HRdkw+k8D4wSK8iH0MjPvFhYytPRy8jvIIIguySxMYEekAlKRJKgJ20xBl6fzL9Jdc9EEkgeqgja
YQ2EOi0EMi+N828DTjXOz0WnWRyFS2i4vxKmi9RRzLWZPzksJr4tmWdKeG6S0WQcGb2RDZNab8VH
vfp3pmasK0fCP64j7KA4/l5WxKQ0jaoo09x5u5NOTya4Cqhn17FQcIdaiyNpj6vuDPjvJrWZY5L5
e552E4SDDF7bx+S5YaOpwHinbJ6jPyYAaIKZmY/lUADWOd+JNpqTyovqYITt/KmYqsVTmUFlPtS5
d7ruFMB2PGrhVoBPVUfN1+SKb8cU/UQXN/fgz0VAQupoMukF62hV5bFQOM+3YeB1eb7SgTkhG7ae
HFLvEmieKIFzNBhV0Ld5knFNRhl88++ObHhhmiFKn5fvP0hC4os/CjTH5adw6OKHtw+N/EeUbDRM
hYok1gXW7PT5nkuBfpoxA9Zz/0bPQK9Wxh3dltNMy6/ttslG/J3dLpoUF7v/RkI6uVpmBIcv6NnM
YEMOBqVjWO3W3lc5WQSZIlcS5BAbTenQrYDW5tu3ZLrQ+mGI7iKb1UrzLEWrhc9+ZU0PIdiYDR5Q
hUzGlJtcNy3CLsQK95dhiWfKe3krybnqGQF8NCJMYqSDxwfckePgtpdDk4YYH8rsC5h3hxVu2EVy
slNLTTtXYoylasQWHYNVKT+8PZAJqy69Sia+ztQ8WLcBy6TH17tz15F0EclnFlhSWUouZibh4fkf
28RxxGq7A92NzblsOlDmpywTxfShh7hHlnef7uwSWop9kt5slFZxYxiK1ZrtLXhnyyAOgDU8BH+Q
w7KNutFWGQtpWfk+0v6jg9sIG4k/FBkU1ota1O3pebFEascrbRaxO1BdCJmJwSrjIkg51abAEf/e
+nYFhKSiCA8oxlcA11ThZlIauXfNbkrJpIFtqZ4cJFbbMCWjcsPsENuPS6w/+CPN4N+t9P10aw9Q
8jPvm8pL97wH/r380FbZ9KzzZnJOHSLrWFBH7nunWjQ7uDClD7VnuUJ//gCj/aQHq8TdjsuHsPvE
vvtJxLRPuSK9Rt+0LD4qFOF16OeV37rmiypJmfmpUP6zL3Xme2DkogxiBx2AdFk56mKVfNUeBc6g
gEAuKg1nTZzUNR1rV6cEx3OmxT0FYqtOcYxZACSQHIXzuOnEKDc8o6XwFxMnXBhg9gTyLeyHn9hx
GEbMKwx5JykYXo+yPIeAXj7dsuBQl3363ozJOyioCPrkpmKlEoiN/nwD50tgce8ZmOYRgUtYp4NC
GLQwj1P5PUuB3CEV2j0WXs1B7E9rudTOkUJD7Bgi7gwgDZnfeijg0bOPetoG2hobUFDfSi3ECcPQ
B6VaaTs2w/YkgxF7aHuWPNWWtLadyEXQNjtKeYE3JWrjoIdME71d8IjlyHy7j0lBn2u5n2+8Ogz4
WlQ5M6Azl0LzalStbfdKiXlfjn3J/acGTZS02/rE5sfjafn4wbNtj4V5bIZKfVAG/DEW6yn+Qv3z
3gG+wIk9SLe3ZpUliVkJUeXAbsCqSkhsCgmwL/1R9SyAv1fwHzC/+4hpy0yQ4IlAoaKkkqaa2/j6
PfFyrFVnzItirDmO7xM3j64bs6rfxkxD6vTV0Rbd/QZSBcxFpscXPy7tAmlXyws1dUOQXmyZ2UGC
AB4PTIpD3dXKG667WcRTO1azMtlINhj+KZ535pxLyrDAQZ15NoJK9uNQmiaShL4WhERP0aoi5eM3
UxXiobnvTGcERd+Tk2+0oIMS83nrwBKrAMSHqXprw51tuQSHJhYNcBr/zI8kHL9gl2a3R9okl7bi
M14dcGa4syNkiz3ZSbNCOxu9bsj10wxfN5kUNWUAfhVAO90H0nOoRST4CGI21tK/5e7WipkL7c84
SRDGj8XVj0uQ6fKFwA3oFzqKzi3bEGur6LJgpiAX/2NU3CaFW8+FFAzdOGtC9dAcBrYlXLeaoI6m
iSe3XSzi7333YJbAvKIvoA3cCE7HTO+zCkwXeLUYnbYlxi7/aswiGYbg31diUXonvxvwm9BOg7wB
yLZxw1ZVjGa0bOuqc6soRU4Vre3pH/XFHbnnGH4Fe1Vap2dGiU6GURwX3eqeWa9SUDJ1KEQb6kud
WdsGPCeP5bS5kwNFBTi40izxxxdNmxfkjE0jGZfT8JCKddPOz0R6Ty0IaTZ/1kZvCx8VUovySwJc
ccx0IJ01s9fMMbO4jqQ37fO15eVzfCenXKbDugPM1D270uPKhtfHrEEFsLT2NCt02IjAHWA6Fjpd
y5YIE6lOfIAs9wSfUyMboQShhJCctIJinpqNAvY6AS8no5q637pwR2MoegTZgqTvHmlpst7OyUsS
fjdW6OtyEFMVNlDdlc+fO1m1M8iwx1mDuLAnQNP08vD69SXapghmqsCInD2MnP91lTOlcvSQ0tcz
UsHuTvawFk3kX1HcG9ow3q5fGWAADX3KPN2in/2TtA/CeBDcOhhbCdFv4M+/lnmBSv+rKM6JCLzU
PYj5/s9LhvHXPuIi05qqcHXVOOfEWgU7owGonKbOsCMFwNXcwFCpkjXQEtw2HaNHIduVj06IH7pz
f3KpfaxuSuW6T+SSjucUs+q/n9GI64SUWqM1LiCRXqp9lkoCdMWb74IEbMmJFWwxYrIWoME1RghZ
O0R3EIMrp6HAT30mq8/WioTMbx4UMc8iaopk8rET5JREQo6BpPB6No52OigZAshX5/zo6Xo247YA
qkptR7ULRkt4kYaoncEVkKMutQ9gg1Zd5Ol5qIBiZXUY7u7NRO5qs7DQlYEk4ojrc7kg3yBpNvHp
+eqfXKgTWfBfo3i5Zx16dKUYZTNm1l+ndZCeg7XSqPz7VeiY5BpCOmDc/YA2ccCvCWzp2APk99UC
HmoOmVyYcNwJQOB74JJe6YA+HYbJiChyDjq+JvbrrGwrnhG1YtOJX1MoZybC/EfJnFMzlU6xb152
IhxTtFnTM9ScRaU1d5VbYLjjgqBRUt5om6VKDA+FaB6EeE+yR+MqwqNFphwnvpqex39huftleBhT
6VCtmYcz8j7KjKN3Mmy6Vx6PVGuKZqtsKveiaqI6OffKFH0wU1L9i34P2Mzz6aMisK9vN+hcMRYm
tjKjHuWjEe4v1DtippoPMjBujNhW4ljdqXHCKfJF7nShyiFN1bPp2Y0R7Q2iLIjwrW0nnobPoH/B
sm3QhFF9epJU/g5TNzE8Zy/TMxNzoncrGpwv2hfNi/6q4MrzOc3MEXrL670eAoAGG9FlsIqBGLfr
4nxqP66HE5soKu1ekNG3ofY6wI/gCwJp6JDuCRzmCxAD4maqJeFSiv4b42HD5TP9XkG1FyodO0U1
EneE4bZODP/gofEoXxd/5OokBSVaTXcmIzSCL1uPYbvtr3CGD9oOZtEYNrDjIwtD0MJ2qbhfLPdA
QSRGyVa/SnfW6/ucEomV21r/Q5pDvz7KIRBoKzKqb3lLrn/y3vJY12qu362M/gLMIAlQ268Jld+3
eBwJFkqkYTcJ7wH7uBOBjbw0kG8EpywNy0l3gSCaEaRWDlGXf8MYTUr0M6/JGS9Of1OEslz/42TL
+V4NV+ecFhqkWPS8JpwEGPgbfsHqyzfbjw9JmnVJgkgPSBqxg/MI4zWb3LlwR3x+ypHgtlCsYfXX
3W76TXCHZruMR6bG6RkMdxHZyzE+Aftsdd0Jj6TxEiQSvlbZV+u5V4St/ULVKn/+lc8vfwFjm782
r3bTadca0/5bvAMg3d301a/qT+3rpa30WzJjdCVXOY4cYqNTiR1ymLAiWwo4CQ4oi1co1Gl+gKWe
WE41Fe5pqVVAattL3wx+00OhEGztD2rycIQw1rBZ+jc+wTTkNbswgG4QuDup9cv4fWQyZvJlTBPv
nb5LieWQrUD+xUIy83m2tRPc0xhqIH1TBpFfJEWAPmV+1p6U1pWj2iGtwnxYlXlf/hiHsZiFE/dL
HOhkwfn3IX9O8G+A/7utmuf4VxZl9imrgOT9jD8Q0sISBYUzVcLfF0XMyPcKe+j++HOhgAPxZkmN
sHeMZiK8VGHHnyfmXmE9nOaY+1231SWxqPJU+WFIoTrdUX/rGGkOgHAPAnTstt5N5Z71adIRIRGT
meUPyHCOaoWl0TcUh82g1AQkVMD+2LlSPI3/sbrXYk9BhpDTJb2wVDgwoJCGa3//Sll6vw6Gz8a+
P2pkKD5maowYNUO/nGP3MloJsDt6t/3Mq7bzA/5uHNwcW/P7yCvwmDJrJVRl51AHt1en/3jMnwzU
jkSFQbjJJ94SByldCpkTD7po0OA06UxP2coIWj8WWmHlaSgc4V1ToNTy3ZBAcGC8jRZGtjL6IK0l
BxBtzACRkMv+65rkmuglGaRhCW1bLl6S2d3cXvg9meB9d/tAD1Hcc92ITV1prK846TOjW9SxIrVm
4KYdsKBYe8LHuX0V0y64AjbUo4n3HSCkqihw31FIneAhZK2lARFcRWpvzICIuGJyzwT8fnNuoMiw
uWIUw+e0/ZrF1zVGNT/Ohx2ZZSgUsPIKKUye8CeujfbVOw0W8/3Q4JY4Rx8m4DIQ8EU6cBrGmDA3
j7Hkydfkwg5w2sOQO1t8v6QX9XjEEfyD1tLwoehxM2AvAUbcN+8lfmqnUyZxeMsu/yFVjTaXIpo5
CEbrfGzW4HO76fiGsG2vnxkVLNJC3ZpPvHDcCQ7guMAeRf/dsyNd9bkDMgftaefqC5oAe4Z1jfwT
RU1gERWMlVYbV/CE4A7eE8weOuDZmlNjF3PZqijyW2Ke1rstMKLrSvHQlrnBbr3xTpLywjXbEgn1
vLp48I89VyZhkfGWji6VWqLirwu+AbI0WzdcBkvP2jJLlrgGtqMNGc3CbKVSde9mGB3+37Mjt5go
elLkTkfg8O7WZMsW2TIGdQtFiPNzhHQDTWmV5+Mv8tu3RxPr9G0Fz3iwR3tvavtyItWz22rIEhcA
iww1mPPhNpKe5dubJlEI1NqlplnjkzhwmWSE9xq+WSiAPCCUDyoGyYP6OJkb6QuvbtMrxgQhe17z
uyGQkpLwVxdBeMkPzzmWRcQPjJjvtjfLFduBIn4DpVGnQWDGaA9QIHTAI661RyoVog0+jd/XWngu
6IrlgWuzmhxBgZCdA0OyEa4IrgTPU/NbHVWO6gejhAaUOiFCZ8IEEujcQ+FGP+5FTvitW0+l32Kr
gjtvALHrQgM0hzTN4wqkApbyXfGi0ga4GQkqIosug/+dywinfiDUvaT7CcYG2SdvvrjzESAn+hMS
YsbW7dm25uumPbxU6X71NXV/bP2crvnORMUiOGUQ0acWrH6uj4dspAC5K3I3Cpfe/Q2pb5UlW2gR
9sTFV0n1xxK8/XFH4SmUaE2U6Zx20QBtUBdsSSKZ1iStZD7MJo/oEXi8VU/LAq+kK4iO/5kJTC4G
XXU/y5AUs1QCp9ZTZrIfvxKwCMDK9D02FfxMuY8QrJ2wTjcAGlc0AJgFHDO1UbFkE/1GDby0U69n
KtLtJD8aAxUiQ6ntZXs+zctF/rSpInCvkMIQ7ho/F4X+E2UmeyfQM+4FldFaNYEgxSZk/nkIwYU6
LciMUUJ95XjSABmPsFvuCeg3cNtPd9IoERirf4lQaGE168E+yfwCOcUh2zXZaZ1jRr6fBwVPHrE/
fNsynoE73sG+Sy6gka7r9WjPRwm0EF+NmCmu8HH3JWZKp9rzmzTIigNKrxRRKg6p5jnUuCaXQFc3
8+vr3zX0cfU16CeYGE3FQmhYHgNdaTX8IynPh+61QVTigVED2mkKZ10gRUR0dDPzIV2x8DsmjhLE
wm8KaV0H4fkKetMM6k5U9oAfuO///s1FsQhHL+mx8R1odOEKhXilStTJNt2GxZaKq3OKjGl0yNO3
c3ezewFhXBKmw5Rx5GepsgMJgVbkiBHaXLlXf6FyaQ1FWS6/4+jMdsWZrCoCBMSFB8GNmRyDVqe6
Q88P5AvwZc0GJ0GKoJQLTT1z6esk7bs2Uwr9gUhWFpEI/l39O8uGHUNFeUSabNO3p5SZuiADRVKs
GInl8DUv69WVaqa19XeKMUV/1Rbh5e3q6yC9qN6oOJ3rnX7rKCH4qLyoTuNORpyGip9TuFdJpCKu
utFJOe6NFxtfTygM1UilFxEslnm/n5bWWzmzbmKGJ8w5BPuT8K7O5fhHGbvsvIZUs4wNI1eoDbP4
w9pg67Dz1VZZTZf4wKkchqFWRwZPI4SIb+XjhHWYYVkRplmvizIJGG54phrqDUrTmaVO57qRmf7F
n7RkzkIJ/ax1MmpQHMWfOiuUV0Vkjvzx8FXt5IW9nBzegTe1b5ZpJLP7A9tZhwjji/e7+JVFwCny
kZyl11JZUQ4gFRf2a/AKOIjPx6cmkNPHA9a4lYvnzHinRQZjWr6aF+EO6CgjHvtpKpArhZSbU/Ya
u/xwsw8GNGWXiZesudXjzhxbYgwTU+eYgJbLo9Pt3N+HScU6aKWsB4KFLaFTlQbLvkKZRxQX7xaH
lZd+tOQQfZOgZlVEzwbt2AS8ENnsuV8/4rIYRyv5/pDizKfTlJStxx6EtZ+C0xdpAqALCokzoV+a
EF5DFsd8sRE4skP/+A3Umr0PvV778EzvySVX6YJJNp6V3K6PAU8+2YfibGnJXFxNOwQc6EMSv8Vc
AiK37qyzwVtD1uCled4erdGM36BM+kzb062nkY4wL3KGzhEoewABoVgQUe2Zekj1LU+7KTnWq7Mq
myt2xMNyB6vGwrsvG4zNU6j/CRAVeVmp/lQlXkFIhv1wvGjMaAZX7NNDevuu2Vpt5YbO68IX8042
3PtOU+ULxQdUP3Lom2gGBYV/wVYpNjw/2kgMYX0jAi6d1suM12QAe3CkJLf8DSnXSU5SPKrSgld2
q6pa7RARVTMV4JB04G4J+q1PCBjPkds9LjrLmKAgWsxRmVUzLZDxQ1MdhGUGxU/KX/FYAndJdHlC
fhOGX+enUWnk9bJa9IHTHezSQjqORBNEZOWbgAL9ckn5d2jvrgki+M3VKrQ5NAFM9ywgI1ohclej
GvmbFijwhZCVzFJFJjVwKxmBR4H1REEzRUM+7VhS50oXYN2AXhZ8T/zK84U7evnfqDb/Twmw51qc
P73p8QUEMoIqGu7YEz1ppPDv5p2AuKUdvgplhjba+JSGq921RDSVjLLVxr9fXruF4VaW86WNr4tn
lFltgQ4YKm1CuxLrEInMMK1NN6j7VyOm+lAld0HLdGPWSsAR2ApguBBiUWKdYqZN8u09KfKSxmDT
1/q/Qgs7usItq/QWM3t9L2sQyCgW0U7nY4TDvGtqpuUm711mMEK5D9X54hXrWTwhpffQt8ArXcnw
ThY8Xs+LwmDLEwpZwgj0bqp4bXLwfAqI6lRrx7U/uX5SFQD32SVZqeJHSNB4GoNxC76pOXg9uqgN
BMQruvTNrWMR29JHWlfM8wjWA8bbcHUmqdnhNE/Yq+p9PZInOpbmdAs+1wqcoCFHkJEs8GD8VuJS
CXpqzAyEWa+ombufFonzRBgMus2WEmDBBxvO7lS/4R3AoxY/lLeMhmhl9OIjwZDYaMqyhpRfmZiS
oN5YW6yyppL6OtW71ixEonwUTU6fIXtmiC5fDQaZYmX7KI4ihLHMS7ZwQVqmeKpu6PPrd22hRJ8p
iQqUT7VYRDYC22qzKbAcKsTgG3JSsyhI+o0zLY168x8MJDWA2yqTQTqdgKZ8liGYu54H+DUS8RJG
C5p7QkvlxpoKiBCO2PnCxXaqly84MPfckDF2CQHJ6YNs5LkdG0pgBAvpgmBKmyNuz6kVL9wqUFRv
5lY96IcJYqF8vG2kfdNcmxmMfHuHSlo7s60OdDciuL/wMGIhZdjCx26O/60wA9gW/mS+E5de0Fzm
A/f+jXF17mR6HmOUWihHPGffGYdZCZKU1QOIPHZmg3WEDmYCxa/GTzrfMG4AQl3s1xwKThTLx4dy
gA2EDj+cPZiI5/UANmPulnb2pIa7Ge3O7JqyoitxKa183mOXWoth5M6NP6S1XBhzeYu9o+qv+BUK
PMpQxXlHgZZ/CVLcz4OhclarKLWJySNnK/MuTKSD2yLoHXJXbeU+CTRWCoHw3wPtk8ALH+bByX1y
KS6TnivlgvcnffjnkSZUMM5b0LdPI+479QvbldHxPEPcOdpSHX3ZXAmwLNTOfk99qsaT8ypKD/b6
bVaBT5nKGpqN6zF+Y2k3NRtl4ipi5vF3iZwx7kxS47MZnwtWkWttrdV7UwTmS5wKBwDwv58A62Iu
VMwz7H09d30T0HTXEkxFn9I4tsopF865FaoSIWyxF38gNtK1QLkLWdUWH6UUx4DlX77vd5HbBmO0
ieD/We3ftCqtomPJl7me4hp6dpjr9gSaBr2zb01ZF/j6LlqiNMY2DafRen+gmmA+wYCvEt42iAU4
EasK5Xd0y6iEB3wjsDDTmDg02SLV6jf39p2EUJrWzaP2Yr07Z3O1gZdh0/uFFXtGCTcUfoo/nngo
OKfYJH0Ri/YWQBBLN7dC2uZeLHDPtlCM7yckuFfwIaA/REUx28m3AEjVhYG5O23qmaN3YmeAz/1K
DVLk/K5mMRJPmbeyqsmZtWsR3aux0zHAz1mUHkWNMkKk/1PiX5jQAZ+Ci7b8SYDUmenmwu/1FUep
AZvlmF8fY0A6zCR8hopVaGf1zIhWXhFfRBpv0b6Jlt9BfGTHt8EawamIJS2rh7Ftz9gDBINTnGZB
tDJJZX07ZSQQruJ5GKBG7mb39sHHE+rigLQBg8KqCnCYx+syaNae+VXqXKWk68ht5WLU6v7eC2DD
6/5qHFhuQlJtZWCJgHGV2xobQFAWfVNzIxr6TEwsr3KP5SoIQXofYRjQ5a/oSp1t9wpoOXEzuq1R
4MLAal23dHugbQ1JRxbXXh+Uvr8uvMeRYB9wiQI/bsbRFbZUX9FbHJ8ZH60T+lzicqCp4TqweBxH
M0q1lHP0BE95OxVNUoEsiD8vgvy+5wO7HulMoyH8hBfPWHdnYhPviArYwuG+e9PPFdJacTZwAS+O
huuWAGjFCDfeSpCZGBgyauFShuYJA4EAfSGDhYI3FHMTgVeCqzZYy07zMGRhG/qRqCCyQ1sCYB39
U4srUpyy7a5Yinr6xO165S9j9DvJdSfhwbavySeh3GS+dIp47YPgzAUj1YlLa/7GEp5uK8ZcUUub
O6xOuxsQwuo3l4wXupKb1aAnNKIcu+xyVfumWOq9aruwIzLToyCyiMJ5gMvPnl1E5qJM4ezgw8OP
F7eSfDpIBrGJ0QwstJA61YvIwptCZzQ262RrhGwjCGACTj3vdNLMGd2QVnLOx2xsVBhXLrDJ+5hf
2RTa4iVNX/w01SMFg61HJ8qz/sJNx2UpkXIprTaM/0iNLHMaRm4ImOiQhMSfkOkDWgS5WpE4Yh2H
tYL/fUJ+nw15CR9nztnwX5SRQZATdRHT02M8TuxmepQ2fRy6bB1E/CgpYb0nuCRn7Pm+nImvKwXz
6nlGJ8+Z9JAa5yRFb7mn7cHSPQR6e7VHpQ8Q04I8DCZaLunIg6G/wZYsXojNLgP/F0sXW7xIXgEd
f5j5Bh3afFbkp076XXy+e2fEY9dkB+DLLp+YrIQKRxpo3EwEVkH0X4SWyIEhPXg39ETHRDoZetef
kRYVdPcRFoPMu+E4FUrR0Yhb8jAzEOsTLSdy8IaeOyZ6VUdmZRqXKd01d9j0xxdOMgMV5UTJBX2P
b1YLeiQe2Yl2Z7bU00VfOfu/QWEK1ZyEuIk+yrW47GmUlLhOFj8Es6zvoCo2Cs7SzjZI8PrIPJhJ
S5OMRfUkg0v3qFnrxkEOHxdUbfe5oMn25jlXVXPXg2U+Zp2JY37mb/NJQZ4wfWrzfSW1qKRHfNqn
oYm79Fp7Z8UaBHqEFZ8rFNpiR32dFivvVVxqk214T2CXYN3n2f9MONrcvnDl8z/0eEDmGkhJ4yrY
hPc1vkDnaITaBacvwBBa6g00CnDkR8F/iMvc2cJD0b6k8XTU9Mollgy5vqC53NoYha52A2Cif3ki
QnL49k3hJWmi4ANe+zL5ynhvUv0Cv7NemfHYXH7r35QT1PmAr8Qnjt2NwcRaGCUBAicfZ2EG2yqZ
WQFVnoZan10vHLd6aPdi8CJpdLT98vF48HqtK+Fw5a75v9SwP8rQVSGM5SrHUX1ithAKHm5XOjp2
rhJi5DdGZD/Xkf3UYKtCMs19j0iP+2jqyDW742EvV9T6SYktj8r7YtcaL5rziisc2qMBq84rQYUq
Ujf4x0jJWLOED8iEpBI3q7dt61YVdgPKcIGlk9yfp93W+UzlxD9eWr03e6x7ABUwFRSANrv5D8u7
/2cBygAJCIXk72SHHxH79lKbnOL9Sdaifh50FotHBTJ/Y/BZXsfAsoJ0dzBPSGk1F6U1srp5RQvX
O76yZharN/AAr6qdom/qyS+AuCmGyLI8kTwQP84kxfVLIwjYebZcDHclYpz0v7JH0JzrQ9aQiO2j
bGicHBaM7T3O4Een84KZWvpz6KGeikFr8nRg563ATuiYm5WsbjPf+Gi3+1eh6EQ/zDcOx6LtjRo0
hY8LZB7UcfFzRkDZtx2qQgCHHvKenhTjpyxqnOkIxyCRAwxLlEvJpfGhWxLHeX12t+MOsMy2pttt
r8ldciYWDCrAbRhxEelZ1C9LxLNXr9UKYCx0AHi65KFN2c9DnuDyZ7i15Ncjne2yn4kaQ44nMA7n
AHxSD2zXEPt6tWwoImWULwyufCUFq2YnekjepN56kHKIUiCf7GstEeNHsTQR57kFemzRehjjAnx/
Q3+38gz2lxgPyvvpEvnj6bou94oVpKsKRlpMxJgfFbvCzsh3A0GUDncjGqylDPYmY94JuqLEbsCj
edUxqLtU3+lfjPVKOtGf4fHZWh0jUsblgFXXGwngKsvX4RN4bm6iq5WW0GR44w5yPwzXXNnyfPjI
+07f6tLXaF46KR7/9Dcq4ePRFGTHVv1lGAmaecNXWxyZw2k02rtdXJEdw6J5nRCVa33uMPiupPg8
wkqg4qkCyodLKOD5JN/4mQ7WsoWn/Euh5GnwL3pxi7FUkqSqLO2ELotPPpXs7beBmFM7je9y1nBG
ruFakrUd/Oa+mCiRaBJZHhAkyknTx0C9EIxfatauTBNyNgLlfWjo3a3kM/kIXvJajl7ah2LC46tQ
m4xiWG8lH6Zk4noHLpyjiam5RknhCegwf+a+8QoQK6DO7EJp0qC1Mu0ETA/3tI9J9JQsHbKCMJm1
pwVTfThJtPDCHq5EKSqrJhfXTLesUd+i3/v5+lOgw36Gi1RzfROe7quslkQc7DD35bs/Gm4XuCee
tS5KtsoAqB8FWB3h7Dlx6v+PoCnNatHtiNZy59lga+3t3vlxRFdi2Nn3I0nYyByYL0XHTwcsADrm
vhyb41gGnPJC08m7Y2cHD+uZVz0sIz2XURMwYld1FG0Wa42xFISCslDkx4fmcQdRY7tGSUYdbekK
r+PVoycplPP+TvcBH5x4P5aqprQEPTXOgqgeS4TYGRBDtEE7O4wLWKDtpqm6AjlUeIgvYb5spvBd
F/zzMGA1fLZDpnv+zC5C18zJcCSkip6dxvC2KDkeX2xhI4RSPPROSd5A0PtjlU/x4CzvQfZPKzj4
dINPgm1NzOiAACiTPKh1oCdJQRoVH0nwd+Ri4LKvUi2cnNLBYKSRDgBssIxvQ9HlvBxzj8TRjgUc
gP454Zr8DN/5W1nbT4h930NU+pyhQkholnbsLKCXoFh2ebUFIgG8xquXlLPObQoZyyD2RXg+IhDr
9RevOpfU0LBaj7OQpDEERqxHEeP6kQNDDwFWANmWqrbwq+KMr0uupeXUrtB9Aqo+Q6+OJ+Romu3q
nJa3iB23oP0KowgkTFBEP9B1IAWQXd/AQMeVY8vT3kgAN9855JXZf//X9YS2PuAh7kk24USLRKH1
n5+lZH34ytOWXVKZ3Iit4LrZzBNLFjHM3YaH7Nrx9Ra/QIfze3asmAaBRH3PPv9syzvrnOFtSKbd
dk6PKqvKKzsp8y0zbqsyHrNvofTbb00TVZq22AW5eP5zrhX5fik7Q/tKO9q8nSz7gfPFXZlnOY3Z
nlgCe1GYWbpLTh0tt3COZDjVcw3Ubd/hn32jrePtyxHI1wfHagT/zyCNDw7ymSwZ72+JhozuL6zM
zdcMq6WMkf8IaWopIwUJrdymbXOmhg1/mIo1fDW5QetVrAqnbny/jCTtYuJ2IALWPVbSdP0Oak3w
wWBolWOBryMPWyVDfB3qClvSipPt67vbR9ZOY2OyH5/Bm7ilS9kzDAnlvACCPxpcNJ53n2fXZ3Q/
v0o4GCc44z2CU+qGZqF1sXabvZ0nObgbEpZg7F0SR2emsdvyUbRFn7LxI4ynfrqSsaPfkHi5Nl4j
QPmnUBCQRzx0EVuQYz7eNS9US9tyTIpb68HEJdJAA6nI0L4QgMV0jXiQ1w1EG1ubsphGqmV39xp6
cFEQT9K5y7PWlEcgweUJgtTk+kuXfe3MFXWl9FeQt4egHzBBuDUrZmVwmI4s5x+b2hgqZgKECvZ3
Qs9DTUVUGp+XofPV/l9UDv0Aq2zFdL6XDkIJan2HcUwknqiybKqj4pMCqnPAWe5xNGpNhA6kN7qd
c+4B9fId2xJZwqJbV5monYsFRiCs+ySSfHFSbku/+Ebh4p0NYYiTjC1Y0VvIb7Lfe0Ne7GwIDs0N
qmQjeBwpdCvpKUvfxLQpxBP1wrqEznFLraRstNG+Omj+flU3HQ5GHa2zfnQDCsJoQ7yXgqrbhrvK
0L16w+5lfYFs85ZwhGVU4dVrxk153cah75y33y8+V2eE+yXrQDBpsc+GRlyMPkDrRqwEbYiBdU6c
inQ5kqBvDb809Mf1G/U06QO+cHvccsAyL2MQS//XnhTqJaNRZNk/VnopO4Fz+tWh9cOcOpPtwgIX
rbQ2F8Tc/to0KVWaDNHokGZ9pdvDPx+xjJI2szdcaJiDAnlg0eMLcmLk38VOYbk4ncSPuaCNKFpJ
Qk3+/jNAn7ZN+7K+lthVlraynGtKt7d2mz1+kkAr8zOdziOdLyYaSXJIcYf5NFf0f1ICtrDi06+/
a52XQr+w9grrSjAtRbpho8+vPZ48tzcRlBegQ5sEHHkL3SyHU/0XU8i2zTKtKZ+48sElxEEkDy6P
7TNWQPJBFkMzOfBhqXDsuOtNvchYln3lgLx27KyNQApX2T+K5r3UmZ5ud7xOo5QOjg4OiRyrwLuS
1OZPXj6iL/o2pnnpEVRWYxUCK35dmoe9euZs+5zDAQ/oLk52OK6J6UC7uPTDlS8prFukmloBNkrX
NqgY0qZChl4S8q71u7VMfb+Zv9Q8eoimO4o1XE30yjfEJY9KrYvvQ0OGQjcE6aEvvlIb/y+4Rf47
jjpL9sP1J/tI17UVsQx5mKJNK4sQbjggodfCxJlMCTStaHHNqrXSMqZ6d1xUr7cnpzpXDxhml0N8
+mA8COawtn50JdTxfVNHhy7HBAfNzHQfQlXJ43lLeWWI3x56awucAPhS0da1fhd7y1tyT8z7Cz6B
KWqAD/2JtPreFP22YolsuLL9kgN/2mCzhxfj5b4Knt/j4QxI/xvm6Sa9ZWJoL91IP8YpR399eFWc
9lc7iClvPdf+qWKt+M0UnqbKIxv5DOr/tRgarvTMk1Lb0DPJexFLo5OOqIQXolOfZWPfzM7RHo18
bh3mwSLXzYv15SU11yCtpVk974BsZp9fsdEDu5fW5N/H4CwedwOyqgjkxKQT9Uxo3POpi1++8ha7
4egx14thAVUVEhpNc2UHUJZYjfwjdh+vUKI9Goq7UQmoWbfq5GQdfW5HnAyqjhNvT4aFuyFTcVDT
J8yBX2oqSDLOu70USgdy+xTBMDcsneYzHsLzSSY20SetzEM3jZcy6MZaI6cvimh6ffr9xIrmyZ1I
FUNYrGEvgH1XDNu0DN1P5EErz4jY7xI2joOd/2KZd5HSkZVESSJsY/fLIVzwkto3zjnHUqXx1rZk
TpZnc7qsGd1W1B0oc7/2pBim3rZ04AOW7cg5bmXOOl4UTA5KNOYjUaRv/0cmZf8dIg/9bPs5te/E
p6xv5vTRsuldhFtgvOdM2ujGkEDhwQ0kA0Y/8CsMMi5L+dgJZxKkplHzgIyi4rpuN3+zv/vn+x/H
zfhRyv5cCiycxjV48I5hmXoLWZ8nVw2meOSbTsQFC4DzyOGtN7iH31F9vAosr02Gm3NxSjjcAfMD
hktFzPZLMj3s4F5h/A3ZlaiMxmy4WO9nRBAElwwBN2uXVG5FKlUlRsIZFVEXFWGNZutwKuQ5m6ly
6rJxI+cwR2s7n1RvHD6QkalqydiNVG9Ue4HXV+Geim8Rsb3klaGFsIK8meK6fMWHwVgvuMVOYCBm
1GFX5RfwOA9rg+pDCsuFpkppMR0oQ+SwM0QVzk+g7i8iRWsqxJlR8G+/BxpMjKhv44NbNVW4Wh6n
F5HmPtov1KwGjAPEJ0ReXMn98gctFKrEiEDEm2wLTfBUrBKUo+qSgItoVezMcHsdQhCHEmZD9AlP
/u105/HmIIgpqu+AP9E+9/nS4AsesED06POLUoH69MOEcxHPRSOitMs8XtTsxC2kW4ZVBI2QOoiy
7QetIGroulH4Sp1ljUTgiHM9sNMFDzzA2RzlLbwspwQQUgdzsZu38BjfaCSHVVH9TuCf7CPAKmdd
OuAk3db4+PwEY9Q4A96neV9AAwAccx8lo/HD4O5Asm17rc78kIGH8pT2VRr/kmHCRaCub3jn8sqy
UhjKm1lbn28rPjOymd7dXya2xGx+TNkAwuq7Qnt4fWCYxvZoOV44AGvybQRpmmwh0Y1u5EG1M4u+
VQlHksrOX+fWB8sQBq4Dw8RCpwN5ffI+xKD03pm3YkxleAJnbmtfXw0uSe8ndkEe+7eH9z6tY8+c
4wDmk2h8T4HHaRzlCSMFpp2uJRclK2oCDK/kIv5wUJq2SgOf+qrNjssFx8v0xHFpFXZa1Slry/uQ
xWOJYDmHuGD0eWXQyOcLvfp0/nhhuL5/S3Bbd/6pMC4V96ppiGk9cNe3pr7bXKrkVdPpwOHk1hzU
B0oo0825baX+oBLT4/sFG/VYVigRWJR8WyoqDeVMAipcMIU8ZTUSCpu871av7hP4gvmRydhX8K7G
7V8IBAHoAy5sxMG6zI4kc8M38NMAKq7vPHmJE6WIpgkRO2IBxHcjJJLETE1wZxmQwUb+djmXcjAV
zwL3qMDBaQH08CrShu1uBZnMXUNZklgfZlwxxkGaoZBXAO1iNQTDbf296TyNGh5bXl5FPirf4lOY
ntyuhT39BsXQWrVEqs+4KW8IMJXCUgYLMxS3UHyl9qQMWg+tR7IKeTr2TZE3Mf5kvh8xp7OHdqzG
0P95bsEhNYzEwpEdj9bRuXfmyF56UAiKRKfzDYnGy7kk/rygKbfSkurQTCR7A1ey6bKojRxhzKZ9
7St25ODvx3XMDqjhknZqZTaGBvIvoT3cb18UwnFUqnCPCEg2iYYIQ1awVx6nEbp1jI1sDFPVKJj2
Jlwc0L8hZbf0d8qDjMZLmAjYgQWTiarLk0q237vrs/xbTja9dJGl1wxvPTzrMlrocEEq4nLTBQ9P
b3hS0/5ddkInN6eXFRptcw2Ioe4hmEZPlWzuDw3a8bjPAO/dYAMaO4UQbDPKGYIWHIkIEM0fBJRo
9IC8afpVm3eDglsY3ELli1DxE5bG2T+aOMdVtgR2J746H2jbXZujJXwnI/tUIkXFwTX+I0oMO3qp
dmnvupV0B3jrhoFgg1R/al3MkHsXfHoUxmjenVzqH2EAklEuePRojD2mgU/5xGTVtWCMmD1nkVM4
/zzxlRS2+8EiD85KZA85f7D6ncgRHu0utivuPNIz6Ck0TBGHjA0Yp1vaGxt0im7ipLvQF87w9sWA
x1wVwuBWq0DBewM2ORxTxZbJ61bSR9NvwJt8YaTsqeJnkh4ab4kS3x3OIQBRrbrfrz1w9Q4Xsoab
q4OtkKbH7SI6uaP7RFppbaixCngouwILQj8xfb/vR1qYOo0ff4OhUf1qV51kKYfJkbiUFSwOlVQh
gSUqUKgEZaNIL6+UWCfTngmJLhZH1m8mnpT5uWIv5bija6oVnCLb6XT1NzxbbN+wP3dGDA9dFN/u
rDoyLg+DIQC/e+lZ8P7uH9VpMfySBVoO5aWF2eQhILqa5D/nQk2Io+J1rRkzwtYj70T8KAE6bQnQ
j2J1dFx5uEODrAoGgaewo3CEcVcWwsT3Mx/yOOHoN3TIJrvwXXRtPNR8mKpyeA533ZVcEafbxurK
Z0M0NpN+R75CBrYrKMcdhSAMsQ1IjBbFZVE7e0dm0DklZNxIaYP4Ec7zohFbqALUTD2zvLuVgnTN
eFkokOakWC2eOQV+GRrv7aK9GITOa85sNlDQHjw32U0xMkPYTUqvyP2W0w1rZ1a/wMXdpuKltS3Y
bpffAhmm1NJrcKZQm9zyrSi81B+ef0WCQey7LfgyH89ajrPuA0rYx739SK7qnHgly6uDtplKjOPx
zdSizx16F8nU+/Do+O/mDM69Yhq9Hquc5ms7xJPfvRL+a0UdY4qLxAzZp1UFtPyCElNHTERvNNkM
gLlumzNTuGEo0NmqhdtVoYiNKACChymw5s2J2qahQSk3B1260Dffl/bXuvLDd+vD/lOf0hhe/BzK
DNWl1ukUPXjPVbFjOJCqLx7cIk7++B+SwMm3ZgtKxBVaEZxRncAXzaa/LpvvM44mTi4cQ1NU0IKc
7ZBWmMxRzD5EmxjK5YjCduA6Qqzr2EWZ7MzyNNAcHtcZQrWzgp8ZZpvwo1Dr30trAY9E8wbBuvBE
D5ohxEviO6aqWn+/67NOndYDfJRsTWfH7qD7/p3KJDMPrljy1+caYoh+Hl7BfGUiLvTCxoudw1/E
givswzEpFxoSxqBzRhFzOpT0FkPCQ0NxjAAGHrBoJmYIqe2U5H59jfnkoT4al+GJHYAZg7X2hCe1
be/myoMxbZGcbFf6gnsxyCyawHca2OGIMA2PL8aPYk4bTpSVV8nag72SKrLgv631+0oo/DE7mzmY
hzE9skLfsefp/hf1xWTZ26Q8GlvA++bbEDPZ0svL2dpOy+F4zdmq+UdKx/UqcSx+PTKtq2nWdax5
nyi7Xk8UrwT/fYykJMG1TVaSXYhTkLgMrPSKzYMVBm9+rY29fNpDXqJUM7LeRR0BiWFZnCBF272l
TsbxI68Va/Ecpzz/NdV8N5LOFmwS5S3ZFxGyCVUhJANoC4uStdZ9OKXnNV4SPLN+B9VlGbimvWD4
SerHk1uaLVjZxJezGndFyuCiPvcY+mgtMAPiMyY6Q8Gccbz/3SIfrunQ56iuTu9e/Zp3dJc2KFbn
r30v9evKYyLgiG6bq/wDD408RfSqbzXecjygFd2R5RH7MgeTxzPmxos1q+TFFA1iBO5WvYvGNI22
JzcC+iuPgQWDMJjqcCSLbfosWUwEki0J0mkK1Z8KNovW2qm9mT6hT0K0V/cN2tH21GWmuv/gk2UG
5f+zYNxJ2tN2JjCr6qgeR1PBTlBPhPmK8HuozvllnBM/x7/UoAE5KiUax6gExD/18OqSi7mKIjO/
ipgX5mp8KqXhXwUPhpp8K9xGmnMw1rMZRj2LcP03Y9gi0fZYfs8TPaTDBdGOXs/qyN/4PeYCEfRf
LQ1OzHhIh1BFR6xNDhqjq1OFqCpvrNUYSSascNzvJVFBeWXIj8bmajCjLQa+AlZPd2XiHEkxJSNt
p+XYRFj/0rg9fPhfkC4HHoCTBvcLztNtqdgAomDOupTtPzweetWvgB9Wh1yLbeUhplRNev8uc3+w
yUTUvyp5bhLpZehaBUwlWZi3OW2gA8SGm70B/F/rEANLZk9MBIUK4yVMziXCX7HbHf9BHx0v5Trk
Pgqy3RFHBrkqRb+a1U/adihd4x5nwjQJebJCTeIwCRCSeSx678j50GVn5b2z+tw47Eqm2u6xnXKq
DE/il81MdpOHUrbWf+93QC6bTxIDhMh/cG8XdszoIxwEO+qP+c62afwfULrv7FlQ8FwHgnKh8Pq7
LxzDoNP0kz8bYCeqL3QebUOZGiEBB9559e6Dv/X8IKX5/qGiFiBmSKI6gwapo3XSUI2CA63JHPhr
tg8qGNF9lsabSqDEl918tjjLFfsNz95IakyCtOK4o8Ouc2cliZdT3U56q/z/ly/OPZUuozNsWunw
V650YvijgHOSdr/bT+KC9IgFyK4yzpvM3nng+72LPQWofSOA6eHyjTIBiVajqAzpZez36xeFkbLk
OqwFEhBY2CmJpsokT+W5Ih5I//kJdDtRVtjnPa6VS5YhjQEybrRaG+KW705QLPZqXDVxE/kCvbgl
PQ72np+9j3jCOWVEj/pWw90tSOjMAlmp2OEF/W6hGsjdoEBJasbYfBrR3K/br9PwO3Kg4anoPy3O
B2jjHXz2CG2xOuDkQVqlD0LJIm0YtDk+ElkW4ezJ50aBSFRiTF/RrhFBdzSOfPjaIy0l56C2Lgt4
L2GJWptPKLadKR61kI/X2mmH5E5Hr2M8hdLlRGomfLoD3AYLL8k00b7ePOf6vycrOHKyV47satfe
X0BEkvZ+ByVAkg+wQmzFtE4A4wFgC8gCBqGd+6dUvr7XZKjzeUkVx854vasM4X88hRUKWw4F5K+0
KlMeZM8hfVa+kmfWDlwceh0G4JFlNNc+1u1ml/4uf6qjhrN7OhSsHkcOZxjKdnVzlKTLJ8nM+yvv
s8v1T1motD/hBJxpOfHe2NBNSv775MvTGgVL/KqgMOFU2O4LPhxihMupZQ3/gyrd9kotzr5VK7a0
MXvutZlrme6yeBRYOrxkWWVlCBl17nAUtrx5QoLZPdc79wlzH5V30BV1LiLoncIC2u0IMj61Bkl1
qE5SfOLJ/G/nvdcWDv6NYxL61Tci74VqACpYa0mL6U8wEGgKug5u4Bu+rsVlM5wWetZNpvZTJa2u
7UOCYoPfkYeg5TX4wyduD4BbXFJt8FuvVTySX3VUUQtANGwNNWxK4vZ/g242VQUag7AbCheWp7gq
g1JI/GdYgQpqNrR4n1ZQrLA1AFC0JQM4kveHhsiDFj97DbpPkT4QyEjSiPGdxWxyW+8l0gJrC0Rk
veCvT1/8dU4LHYB3NmHn+0r51pZtzCmxf5J8K71QA3JqYTjFuHARkmIHCXn4VLPNSc0zX4ZZMl1B
HvFvOl9OyUs/vAxzXuMVjeMEqHAPNXNt2zaLULCGbRkhYB5/6dBspyHxKupIBM0zePb7Qej5Z9w1
W0RGYOmEUQxTcSiWa12v7RWh4sKfEQn6tkDpFlJefbo6fsxNZZOtpKj8ugcwrdwZ3XnNCSUOwiQy
vO9eTR8utA4TekcEAAVNjouCbBGP5SG4M3i2nHYg1WzyRAoFquYGpxJhuXsoRt6z1HkXUyGbahxX
F7+s3JVnjEkedFzQal/BX4jWy+bgHKVWOfSmTdTpgm+xZZ/GxItwqUHb6rwXo0p0RY5oEx5E9fmK
xu5wWqIkl1IIOrHTTdhIgrEAeZwNgYlzJS8eFk1b+Bg0citVC6GfPRSwG6a43n9YcottX3SXrL5O
GGGDBXNBEAffv1ydD+wxLsUpwBAsjSgMonm10MArYG9mRHfELYhcvrLfY9jcsJEOiQtTOqU2c6mh
cGUHlAdFV8CiV4cdlvkZ5fBtSGO733+mmDnc5o/RyGw90wIlpb6ZCd21kL6jnmkoR1WflTWkIfcv
AtxHAyvT+MOGgmDx4QkAw+67gobRXxhiY+WXWrlx+g1Zz1/wDQCz3ny9YFaN2/hZlf+0wDdw4oUi
0krEZjBYGfP6AkbEcVTg+KFaD8wjqKvYEGfuXJlmP+sFWyGjjcxeL4s7rE+1bpQgMDvM7ipinP0a
UCbCMOThhcpbaY8KnRv3s0lbBbigLSHoeCtDDb3/U5R1utr77qOrKzj74fs8mGfZjhIt9vmEQFUP
DjPxA++GswUon2lRsv/4hyi25Ff1zcmCRh5XmOvlxE0Orn15dze0joAVBJYjNzGCP6GG3jdG+Iuh
NPzHN089yZJluxEnrP5otaKde+wfRDrthR/cvg9C8TRD1wC9k2NcvyR4Z+uMUXJnWxnsK2ecudaJ
mO/Owa1OgNNsZRGooZSqTVULsYBSvLmsWq+9nedh7pyuYNOnr0Uok0s69vZU1qkLX55NZWsBN4Sb
WfVxvI2kg54D2TkcDqZpZs7DbqhH104JW3qAcPycdJnJUN7o2ACB8mkdyxekykJyasmkv/FV16Hr
W1TVpwCxqUN8NqsTwPNbeM4qI5HMonBxh0CXFhA/4CRFCRyV/mu3Z8Fok052AmL0JAcARlmxqgPo
/SvSKMn5/Dv4N5WnapHiWruRBJZ1sFzX9cYld6QGd99VdTqDFdCh64dJ5Z0cSllT2SqawIR1AnEl
7jGZoeHiNyEQXYv88EwqjdJ6bXPMsfWjNSpd3zotGLHXzKr6ZWMRdwUYPjSbz26+PVSIPWdqbm4a
5Dr0c1BGVp8AykxsIoIikt5D6XWm3TXcVLUPX+bU/VsLoUVyPi1msdhejOJEwXMv4aQ+k7JUU7yQ
VTshUAnrVrMvXsN8oG/67VojeDCiEa7hNEYhNRGCsVsgbJAEBhr/Suj2J47uTA9P6+aq20DVh2ep
0UsTF4hIhDvmMVwPx8g3rAV0ooHGdVFTD3OZj6JR6gTrAcVfzfSEcqzsz+bcgrt4QvoAuvrFQYTe
e+1UootxhIhau8awUIFFWWUNYfG4tXaPBrwqTgPZG7YwP2vecLNRO9te5wbMt9YRx/ACYSrXJFai
MPDjimtU7UwhXoCmQxX2q6QrLa/YwMPq72wwVx+TvMmXUdiZzVwq3JuECKFO0pn0y53HpHpqbbjf
ViN7+xIwY/5dOhGvTR2CDrDNtV2DBLl3YWtUGfkqLujofLGd+Fu7PnHXz/ksFqFu7VnzzB9csaAB
RSUKsPHslyflLaROsGh5Y5W0pgzlRNrCVcqZLUCeVYEG4jxamLmATyMWZGEv8fVxK6IuoIzXS8xD
e2g5Yn01HGpAAiZqaMn0K/a4KVLd/rNosCTyRIeSUviF1Nzab6i580/6uauGf1oaJe5ddgrhMfXc
Y9N8C3pZYhsDSEw/uROAE8qLgjAH9ucfimNEI5C9RQkxUWfZLOpcGHdu5PQ1VX9E4j7J6hjs/e1w
s0YmddJAglBFx9fvTq1zl/1uFXWC+T+VM9D9eUt+1GrqBA/Ekz7fmbTCHQWnZxuzZPtLaYCuIpF6
Z9BdwsPHJa7DiZG78PCNQaxgbxwX5md42beZzESK8AfzjMp1g/l+zXVruAzEA0Iy+LTkWQNT/zTk
Wf/dmLWgVFnN9rry8TSvZBdGCYorQ+/h/8DDx5Qt01WAYB1U/2rO/5xd+TCduRSdf5vF1Rtbdv9L
aeODzKp8ZV2CpNeAqcM6XmkAqIjIYuIeNQu6147HveWczOsQYEpEHlc8MtFfe+4aQnl9F/S4JCyX
Z0b++jsYN3AMiRO8g9xJL9//9YWKTwsAkEIFZFHAYVebUbSZbsip1N/Bpvv9/ht4+uzIf/9IFrI4
6MZ65LNd7b+HqnV9NgzhSzbogn9YA7/yHcVpvreT3sKHDcZ9WtQ+OTLrmF8aGb3roBipWhL500QD
Fuv3sQqeSjwoZaoQAcK98SbCeoUM0nDMOvfHUW2U3IcFAAHqkt439UZRt11MX/gVKOc9oD8NNi89
6ISsT7E5HM+TyjE2h7V4DFreWNiKV6pDnBEfDCn9nwZP2d/WO5HF1wxffRe1r5BsldOK4m+IW8sj
Y/2WmGsGrNpOXCgTAinv9+SR8QUz3pWpH4OhgQMnzpwDB+w956Bzr4JvwA23ElnEsX4w3S/QM0+W
k3MEm3CUSgnUaqalGYkMcBuuX+pYACfpu5WtHOMT/2xji9YMSoQ5KO7ZyYB1JKC8BcZYixRq5v8X
+BCKtodS2pLLHE1oMWhbvCaXd5a5ptvGwPw6IVk+yqlbH/227To3O0bazQ6dYjXyZxQkrMMeHVO3
Wn8ycwqclpXoxVGS7PF8EPpqP9jjVRXwXo22+czxNDYKKqmDszYqzX9EFcUMBFHTvvlqs6ITHOfV
V3WbWD39r9fXEhGPFYqG7/y0VO2PJSRS3Q0G2E3tFos4xUOEw68zBBszjhRwdPqL0X8u9uNWJEA1
k4QNbjlz9U19FN2N6N/E9vuxYuk+/ON3RvrLps0YSQGGnS3kufNUXpwUZW2DYh1z81jTyOtDxZGN
5u+3n+p+wQ3NUrVBOMLhPeHSm6t0IJvGQ7LOvbhJ57Yk3Oi/0x70VoiYvLIj9B80FSsaNxDpk6JA
4FvOlj94ucP7eTA55Q1V+Fn5J72m8R+ZNgH3SDMraHYsPU/3MgY5L2VCIbHYiT+YVAD8TUXHZ4C4
u/rR9xJ9s4DfynHhVrfi9yi/GmlMN2ojWw48a58ExaMDQ9UCXcKh9T+M+ISEM1e+q06hvx4CC1QZ
Sp+M/X+9oWjDf69PWewxNUliaEU/OWosI1FaDEDojMSbxXoTlq7LnM+KX26AuplyPO88Ivoiga22
cQg6yIcVHHed24iLfAo0FVJWpp+0QTyl58rE4cgYLPf9iNlg6QdnRD1vrUXkfreJ+EFRssCsNQa1
S0n9L3CUzQCID1ZooK9orvNTp+SBl98lTfrN27qU+8S3AmbuAgL9UXOasgbTj47I5DZvpxl6kBb8
9zjiFQkRWfugN4mCG6qBSj8E2ESRUyDOpWH9I5J0WLq1++48IOXgNQKF3zjwIcffFzv+xpG7ndRD
b/LICuLfoisMthg9uZvRITIBXXeJ1UsXNhJnIENLIGfVE7FHLRQ3BkoiNRNI4q3vlmb5ctprNf8D
48r8GVboTYq3VjOPcbiQXptSTcjjwbUEGFMOg1Fk1VhEk+/tTgUuYdfz6Z41hy5c8iIAhIo9QYcU
guUu598NOeqLR3Q3VU6pNU3NF2yRAWo+jImsLyirDZH20mi3Ac1QmLy1aAkUdFV0CtmjraJTmNtK
48n7ZX8o0Fv1qJmnBbsyHqz4NZ9nQ5I75Q/DP3xbYlgf6SJK6SiaIPQW/GhOYhIPj/U0GshzRDSl
USux9gnHEkg/Zb1IygnLsFMYeTIWWDSrUsMUbt4yHs9W/jPgkYPj0ocwNCthx+6CzE+6cIAEtoWn
Fm0hYX1qSm3FVG3iHudLD6bVDHf1gb3QYr2cLNwlXG1mO0Z+NuqlbmJ5p3cjR50BEde/0G7ndN1k
c74twHHro+kfckm+CBCvjexGiUMOcmTN/6closqtF4v9YHtiRxOkx1nbkxGbXfBtecmU5IrgJfVB
AVPk54KGWpwias5MD5Emv4AEP/4tQ9Ul36WccBSyGOaZlRkTpZjo+BEpkAB1ihBT2QM+1d7a5uIK
Q6rJb0akrXHlrVsv4k5nUvBY0h1nadXpoOAohKphixtNS0CeXT9tIMHHIpss1EKJ5yGvhAfqHyWc
8pwO794ZfSn76qjMSX7v04lUiHZH+CrxbHufTsazXQXd6MxQb6J5iImIM2OZjX52YPQgqM23l/zI
58g6ONauHxqbvLQP12p932CNB0J9m0vLjQgg5HtXWFlGUracOONneaXdJufsf9g4a8R1/1xeauC2
OTeqxlyfKa6hQN8agB6flBDFfenHe1WQTUsZZLXIJ2ML4kBh9vH2HBsyAS96Sg/XWafq/inP6U5N
FhKuadbThthlWwXe6on3ZJm54c3Sx1CA6EfBpNqs+9fkzLWCPih/iYEC8vOCnuqyzvnPPnIwf3sf
jm41sz5YFiLSZSxgvcLRVm3sUtbDNXe/lsMTiXozZrzs6CAUjPR2d/q8dlNueaD6Z+KOWmAh6WZl
HhW/MTweBoLDB/jGxjFKzCK3aCjGhh6r1BQslm+NqNysyCTf9O6EzPb5fPv0INcFH1B4aPVgBgHj
90D+a5MH110MHGbPnrfX50Ja16LGJBiV2aRDgzeiBg0kOxkUzIO+WUY8sxIGpO02yQASbKRXcvbU
vVb43zm0MMKTcf1GAHEPG8KUCkTd/qRs1RFxejzgpXp0K0r1FEYLB/Q97ON+xbkyURp3C/LMnYCO
lMV1KAr2fzTNVgIA8I3ctZOoPrby+p6hFTTPafCdt2yv7E9B9u0TeZap/zXtxZxp1l4wSIlIVu2p
SQewq3RCz5a4dPAxw9ScX7MkTNg3bXRxk0218/937cCv2QQTgZ9OEfsMt0zRoT2p5K0w9UYgfvX6
DvCl7FpCr5Gp/HnspXuqFDL0jPNfbuY5AzBMow+sQsFMw1d+xKfFvC0+mptCRCmDwyukMAhPtWGL
gkSXlfkqC68K1xIiMONEtDfd+AW4subqAdROse1+ixTcusd1kXY/cZdt2KKJGlB8Yhk76NRTKns9
pPaXXj0VBFaKpFX4ZfIqP6oz69rlez0WYz7KdZtnXrgLybretkTXOnNjvfHvHJtGv/v80eVNjGz/
wtC9dbbCEtA5YJBMxPnol20/sZuAwPnn4rgcechQniVDt//QMDvljIgPEqdrIhBnfihBsg9jBbsF
YWkk/j1SAX4guIjb1WS4qkPBDw+oKR+E2bMbwojFjcBmJdCo73ejTyK+XjpnUM4jeIbJ21C98X7u
biLRY0gkEa7HhF+xPPcWky79chYZqUYGF+76AtIbeU3UZ4iBRD/ftBRYfE4IgalgOd5j3+EfIyHo
/pgZlztTkjpvj57lHCSb+caeWxuAVS2iitmcKo2OVaUu3iPlv9Y96cXDT1s46AuwzmEuGsJIvYSQ
JVlUAnGdBwB6+UlYjq1+fMYBf2kHdDQjtY3zIHUR0OROqbVAkMGAYpDloHJlVJrRSt8jtQtgc9FR
/qrG3vHCWV4f/sqJWHQSOiotXJS7HWQsBpj9TKjsEaRx++cCuyvYQmrCfQ9Yp3P1jC2OuOsOUan2
IXLbQsKZCzLidBUCvmcJJPywG7gahWotWeVdzJ5xj2p9zpHTNbGJAXRMxs36Rk8+kI5yMKCNyFM/
zwmgJfpzHMfREn7OsgN1ebQ7GCqs0+quVDE3aAS9y8ygEjMPFLVIQ5QKntIwr5fiHSJLTcBNLpOt
2F3yWxJEYFGITK68bH1iVQS8v7Nt2gpyMyF1Uc5c2qbMzhvKPoxu3bbD3VGNIOcLmaAG98F1lLa7
FfQY3MhXQxsfYIKTn4EZuNJ2CUtk1D441qveBUC6rimAPsJLjc4FpVDqAWV3PEr2ne8qtvqr9mvh
WC2PCuvGeTvnXuEgwXmD0FYXdz3T+dyk3kk12mVtZGrSo7dBJTl4JVD+2xIWUbOdDm3CGPhONwvT
wkwR7SQx0aCBq+S13/1oWaDk3tuRbJcLKK3TFz6IvnU4aDA17BE8vXIzl+RrxcTYv2lpaRotxtts
k2uuAHbs/YXNMajydMOpZheXQhixS8+0bF3rSWuT0CF7h49stQ3PLEjRGeoreFBVGh6MEyUjwPec
Ppn3AaZwnZT8TmrVsbjQ+08XjNJOCjYyzjaU+3C5suY/vuzDmcJ5UxuepYbNhYg3+80QwmlvXmai
m9OMEODWf9sBq28/Z+ciSG+MWJGXoI5OGFhBNXju7Pkt7jeOmFL+KpdDFSz0XDIlMuF83b8KIqTs
Vyo+a7F5kuzj+Zt2A0Ec88hiCHBDEdouEG/bk0mlK9ag8qomUdK8udRVxMP22QNTEwSwgqrV8R5U
ZJfBH3M6L+wa9wTOupQgdDxzsUCBx8JnyFKTVysIAkCZFgbYfpwPYx3/lCRf2jGMkFDUQ359upuq
F4Pl9T9/WgvHQjqW/2cL1rrFOlaGyWBpVg3J575OkUrAHTzY62RnDjBmLtGxdUORTHxh8NmBZ6bx
QiUJn080jQHlMHL7IXPtC+pVEH8/v6W0DBDs7by2jNZ5zcrpMRXXDF3RlqU25SCkf5Rur/2YDzyM
71crJvOfo6ZXGRKOZr5jN6LlZd/To1ngZb+BAsB6JYFEi/W349RYeKnjGQHICyMx08ZCDQsC6KVC
qFCSjAg7hZT/XxTICuV813RPMDl6r0x5aayjqLae6q818+YO2dii/UoX0BhHZf0w+Clil6La9WGN
h9NshfkSQC2i39NOfAM44H8pwSUJQ0f5mXj2zzWdm8Hkstb698yauFmBaaddkA3WMm+uCfLQmkA+
ltg0KvxfKWkd3QyububsGaSWaoqqXb2APzmHRhq7O2hUkljT3AIzcY8lmRzrtQIwJ8am5Jox9NHS
lII0eEb+U1Y40fOpIsdFprjH2otBjWWBCKiq9rlJINbX/Oxen56Bshr+zL9vFJ8MhCOgH3qHW3tO
jPmvQVoNWO4C494AAWKiaKIrkgFS81glNPtuyJgvIcEVG3Wfnt9m9DcD++Q/uUQajjtZrouhhBkG
QcnANfxdbIwQqAjS5MaWnCCBfXvgBC9wJXKxIAlwaetwXNWEuIUXzPaOYJdEx54H98aJxYRDQNJP
PQHVYTHGj4DMCTTmngNMewMVLZ8rHkIz2XsFBJH/xCpy0zS81GWX2aEdJD61ZfDZN5A3rrdC7flf
MXRIQhH94ws+7OM8diK/k6Z9H/qo6ttqAVSG6S9xz7r8uS0izZkcVHOjDPuWzedrJMxxfcfD/+W1
ZZn21qNmivpKAKpMDOPuwKb/0MhPmXcWccwTetO9B7IjLzUpjjw2npscsYbBrWKa7vMueZZctFDl
4qW3yCWOSAJuZntuk+uSZE9GV1PbCTctE0uczY+xBuAGsC0//uw+vbPrcQTeUoVLo8StfRosnoSf
c+XQU/9v/QgycnAiMMRjT0VmQAC7L70Z0WFpU6Szm6GY1QMm03WcfmXjlmE84FiqS8pINEzHLwjl
O2ReQlsZWxEhPUn8locihIKcatpyIJmuchgwUpUkf9pejSLxg7o7vJ82QiEQP3uabVvp4f8q/zhy
sEVkQ3sKaRpr+3yUDat4wFIEpEqPqYUMg2xr9cts1RYofxDuQc2NTYRhrcJy7vQi7MJh7yV/8o7n
ScYLSZ37tLOhr3NXYtnR9EmSnVIf1iU3rKY5BeCaTgK5JB2CbnTJRF+rSPsrLnhF3yGd79HUmLcG
/HuXYr5T2jDgFR7Te/zcbK9eySu62p1vrIbJh6qK5e/qU79uX6TWAmmgOT9uEP/X+fE5mIwWeeyX
reoFJzfEduePOArgKA5xPB5YR53xanJtgXzrQNEPLO/UCJ4AVPzaOsPsTQZIWHyefCgHb7ta9bto
8eRtUZrUe/gsmVqZ66pEs2SwFrT+k48NnEzpK1IAcYCFKAwzdfxPVNByYL3FEvCiH7Xfl3PU9z1k
Uw3c0I9QlGsVI/wZywyA04rn+FAHNOfANIdqPsR+qpHs4jXIDkC7nWxdJNsK843DfdjkBlh+hJSY
AIkxU8fjIDTdZlrbJ8bQ2cApbhCgR8Vjwzk8uLghU8Z/1Has6fgloL+SkaN8JKPmy/rOoLCYyM7p
NSv2fRpnTbl9lELJ+D3LVCsbmDa9h6oJW0CeH6vEXSpcNRbCVNhNmvwnheB/N1R5QOZEOMvaofoM
QiqgCostDAro2ZFcxkcBQMnywRWSI8lWxWGsq0FacKaigLDc4UIDR2ddVlgRbmZastGeWgob+bXg
1wA39SJRWgb1tXbua7ip1xEALm+RXgBFHb0H7CNSiEYc9aLgLlmVZdghNxugZRvXRYO3TN7u9aow
riGkl7NFq82Cqp22gwpgltAkigE9337klASNWwQZN6Hw6BW9rArqmxzc8fZForOIAm+emTIa73SZ
9pztJYyY2Nk9km415BaTBGXu26QAOQIzACNHDusildrm3zhCU7YwpkZd6aKk9jjp+RYCtXiJutl8
iq4cUfB8J7juwnQA9iFYVeuqXELbWUk5r0oWSRq+gYBG3TtWp5Zui14J6yGBX0Oe+851S8plNmMq
vteWxe7hG+F5L7SGUEv7xCnOE3mgIXuyvaYLercZmB8iE3wcVCyF6grcR78Zn261L5uFQq4uaJgG
HjMkt88Kukr+H1iaZ46ju3eTKRiPEDKRqecvbFKTb9rTvBvNyG1c2ckz56jn/o7HitrvJvGYBs0K
n48J43EdNiTdaM+inJ+Bb5B5OI4u/539diApqJtjG6e+v2tH5TZwyjlqAhyAL4J+eY9OBDHAZgH9
IJFlwluYXxQLPFzgffZIi6DS/1OZqQ2MrrnnYLuUmA8IFQ0tZ6CY75Kxk/9rfk6ogbBsTHHTgTX5
+66pzk5ULH4lrCQlcnY4ZXaxali/KOM4q0UBHxe+zdmA3H4h6ccU6Qtvlgng7/WGud1GNbIeb9Cq
kWbqU9GFPPXy/IUVEdy3UDAPBU4Pih8nCxZK76UPytsYcWU+7U0k3JHc/S4wHcXxH9Q/HJNIBIej
Iv56fd6EkCtwyY0s+SbUYAZ9P1GwMp78u0vu+JH8bgTI1Z53CA9kZfW88k/G2T8YehUz6Ik1phiT
P4donvGIZok77i+R8lBnPcFS3hY8d0WnP7scboSbF7na9VB0zSyKZDa7enQRHJoXEYOnbW7HpMx4
S1uqhuaE2cKgsWsfQLWMJcqzwxGU5jPdhSSGLLumVh0Z9kMI095lVfuv1pnEj/ZSTVbmo0pPmz1Q
yEArcYLpRnCNiP2ZkqhOjbzvMDmC0KF29KYX1UxfpIQ0ZbIVSEGb7auuMUjbn2zqh7u7BfBSQghy
nEvCyygzvArnVJF/HzGNTvYxC2JvZAhfrspvUyhZm48hq+AqKPtuAS+SZb+U91UzWhdpj6kj1mcr
ivpoCbG8YAxUqpvWwWaMPWFbzDqT20vuY5wbTXh78qz4Odsxs5g09M2RCPTT0nEC/2e2/tVJJVKw
lq4G6T/fA+tP+BvJ1u+3Kl2FO6/b0fnY1bGn7sOrJvH03Pmcr79/eqaSPldfWGrELP5K1kAaOvwW
G7cGqC7UMhOVX1q2hpVDB8fRnZnIO1DZdn7T84IXnQEYz8N7yH/WPLYPeSSjGyrtpQkokRdr7qvZ
xGDAzMmlmdRFa869wUSnvOJd0S+QdsdsKnLw3fbiYJm3EalRBt1wRawE5eNa0iBiiC2549ri+kXw
YopljQBLohtrDCN3FU9KVB9M2gs/RZg7rGzguPYkZlSmP8yAqici2q8gCnS+6J+qpq1PvtLyOQy3
feUiI0TELZMcNAdhAlWL1mm6X5E7gBGHc6Ra8QM7vK6uY/3KbvwSLvsmrsgD3QE9kAZG/WT2awWE
NObcqsrD66dc3gXEgotGoGrmJBX1caok7BFPcBZiMrud9BM4ZKPoLKEoBPfKfbb/YK+B6MZSARi+
bmOjzFRnPvsX/KGEFqysR/G+2v1XG4ojppFzDxVG9fU49fjDwSuK2FZKliTSK2xbnR4Wnmulis8S
dIQeHY7kXWr+uLUJeyKlLhszCeOz8J0eSgnz5ihPq0iFsqgwTpaix7TIIY7mtUSCvm5IgB7d19rc
8Yis+jw2nL+O8SUH3Xhdso4YHGxuyi4mL4YgyQTF8lYapnQnxlyXHxmFXCggJQRzOYP0IBwWJd+T
Ev4n0nGjCKEV/nu6itOMz+oPxWM5K+UjIT6Z2NOP9HMR1IjaPy1Fd0rHvGbvNUCX8nUYNeSdWakm
g/+38saDlCKTc2Jf3OMpjAogBcGs/ZbCbt2tGjifl/gE7Q5t+ByEFZ0AX012BCAfZFa0BQJuXbIj
7XPmglggTy8PHFMTCs77lXB6N+195cM2+4rRn2KoaHnfkAjWBcfvES3EKvSSEU93vR8ZxkE3tunq
Lw633DlVqacNaCU/u62tZa2j87cXS5BVIva67w/VYZA08z5nSFlxRgLYZ+czUTlfRACHSwR0R7xt
l46G9KsQftsSd4YXa/0/6kLmDPUOmzd3mxN2TsJM1LGXHkGHfn3NFR3tDMGTKGQrC/BW9t6Efsk3
4KUoDGzcQwpNbBiN2Wi3aPaquYeX97wDKEqdUdIwJ9Kn1SRlkxBg5XUIkS9qFWRyB5UdtueSm+JF
8XIxPzot/mvZngDVEYKHs75srdgeUyXFhGE6nJrepSsmoeHmnP+byGsO9E/ljrk9XX8iz8lrrQcw
XPdrbVAsDwb3PlC43haOr2xzuvQXjmuoSHjZJ35Vdel3FV4X7n8j6WhsoopRPi2H6Y9FO53LOlTB
G/icXZE5wWA4pOB2H0Mqi2CJintjnanl1fgJUzjuS8686TovoT4mnJsODZ515fKvKz2trNqh8ZzG
LSTRKWBvJ0c1PNuy7Xri83oItQyPaDsW1ScvAD2LbHGhzPn3K8vCPJqgzncqsOIj1//x+pYldIpI
6c2BLJrp1Imz7r8v2pExMVAvNKrBUpMy3UGA6HOrxy0oKQKawrOkRdknlDgJmtEPvBMnkp8dkcIx
Dcw5UNoLh9YyO0+LWA122W7oj9C50xhWUqCKyVmZ2gOf6JqvFsTA6fi060lt+thUPZ01sLsikoA7
5yi6ZVBDA89FQ4c9zTuzq9njZanx2/S/ZGsSnwpdCgMSr5PCIJBzA2oHSStqdjoGryBwna249JNK
rf+mYjwDkDngwVskfcP2eHJXe3CMHTwSJBQxnrPI+H+qs60LVFW9Sr1YmUAsITUF1IoOL22Z/XR0
hfsKgjdGEt9vU3NcJqnefg4elFhZ77ms1Ud4loUMBR7PaxI1TqU154v3Qkn/KitegTl4RimV9S97
6EMx6C4YDZLvRKzLL5MD7m8TDPJYZtv/rrSE51jZcVd1+ED0isttw0lgHypESm2+9AD263qWVzTW
5pHgMnR8EGqCsGX6fWbZlhOC6jLsdHtXnE92KK8M04r475ZDneB4isIzOlGG+tRyeOBoeXLMsN6y
FZOwH3zvLTSqGB8Dr8cTqx0Itr/R4p2jnzFfgRZv8nN2tdHr63L5b1XuXPZwCPstK+u7hncMcjsC
KyTQN8sgZ11yxgh+II27H+laOFId7qaIstP38w6zuJWospaI5VWsRREk4C+bIvnNiHT9sk0qh5/d
gaqQBzzD8SwSNshAZ8BI9JflOe8qpqjyC+ekysReM+tti0iShlrHyMaeqBY46oRwuFIR3uy9mS46
Xi8pKe6wLqSg/Q5c+ypR5yv0OT3y7WRA2arA4ViJLV6ZsE0C5nOpzoKwzZgBXvRCnmC1Fxzzs1Ay
iutyclW0VRYM3iBkJs6hX/kH13UaLDIWnsNSDpJS+cG7rG24bY7KP5BOU6R20lUyLX8V1qiVZzhy
tRoKkVap40cPzLFptwNDwdPIDObi69Nm1sPUS+pUjyFf+DMv9GkWQhamv5z/Sj177BqDpR6mvjDx
ztZSsKJpd6iFldbreEO06kFXGA0yC+yKgp9PBvlWeh6Lgdshn0Pu1CO54xVZzcesJfwQDX5IAIsI
kQhWNl9EvX1mr+noEgzFtb1qQzM/EQrDlWO2T7XhVmP/aWeToiaT8rsnrfl5Ixl8duOPtNCR4FBr
D7iiqnbNDyrzviA25vV0W1T2KFHJRXV/NEfg3Ck+sOYjUKbvwrbPBM4Pd3Xs3ch1Gf6XuXCjYqYd
2ztJSh6te4uITKg/WB+lNXESwIomOKkOmqP17/DFerTjF1YaEcfNfgG9fRlyWimEqTgVCvTf2hs+
bB5J8dgg93j+edG4SzDid/RItneYQKhO5wyHcmhnRF7o2fixZP9wC+5L9ayOq5TysnpdHnmq9i7E
QFiYrMzbucBmWpWXvqFzxcq21blXzGbgvGdA5+CmtE7rWLsydrJn1LzrWJTUq0PxmxCX9D8QZVUA
B1IRNwsWRlibCJr8GlcqDEAgc+cqaE8FudUQ18C4yy7+rnWnS4pzzb8NYywn85zY606SD1gjCvo/
JND22BfMoF2x80BWEZn6PE8quEOHHQTeOo/Y4AAU/woJKsjtIKYXNszxQymqI6N5317F/QakTss8
S1jFYLNcYVryNSLwP9QEGVD/p83TccE7jmkZuY/1qULHYWup/8vp57eplZsD0ag37N6PiMurYN16
txi+pABqRql6kgVeKzbUPwbGWPd8nF9ldZp0qR89ApG24rbIneGAb41Vwdzr6w8vpf+j+KnN994d
RPYnvzsDBjYTU/OG32VT1sIddxNnTifEZSXcBqbgCgf4J5Gzawe8W6aFsduvqY0u+cgnjQAL00lj
LxSBobMzVJbOeeixyVHcKeA0ROeRMhAawcG5X2CliWMZBmawGJggJL1+EQulKAZcl7YARNgLm4G/
23bvU6ssCMKmElk6aF9dbNP6/rOyD/CRCNBSeOj5TIfcEbkKXeGiRV1XElK6S5HHv9vcRatzBfk/
OfBeoUY9yQ3PvSKtWdmLW+xB2VDdNRCTGVKEagfyqKsDQFwBfNmxidvxWkvUIlVlVV5Bp7wJfj49
N5ix0meT/Az03Vc2RNPvUA8rNWclNpc/SHXbZTZ8CT1/EPeRJzE6nzb2QrINCQouD2WDzz3smopp
rDl/aVWv+d1m//PdbEqPOH3Pk+Jvo3xt2aKiZHwGG97cXGGjrczCT9Vi6DZgPVnTdXhBUW1zempk
XUiddTnsgWBS79O4alMUuU7XQFroUiKms0DAZO31bo5y1gpSVvieds6jnUKF04Mh4zTyEgyvO/uL
U6mBn7PYOE7rOFXWR315CPFRKlaC5mhHa9HJ7Dlm2/kqurOH+jZ0xoRTnx2+tLeJknpq346qALJy
Tj44IvnYJPyPQ8u3qY0bNyLaQvI/RH1e4C6YNHlCWxrt7QmllXiBvlvPjHUAgpOK1js/RpeTNJs7
9OzJFOUsU3wORaRT7A34mHp0SbOtEFp24smqNE2KpRQnx2YtAUrnsBkMc4csnpUPnzssPtJp4y/I
hIXBGmTybpaCnlrMQ4UIdau6/U50Z4Y3Wtw7sIoO6NSw+NdChcLTWLKOhbdWB9P19fmwRRO5DAJx
QlVgljnCIYkL2NLYt6sc23Mua+zOlEZvjNBjn5D9xeXz/FuBoBnjLh2rgH+Rsl9Yy+7eEBtwLu/X
zgQirsd/2dZ/+ttE/ilVlm1Jdg0MerrGSZedbQsBgLu6w9OlBQroXg5U1C3NBeImxV8U4RsJI61h
E3z6fWJLczijIVpEuY7kAfjqQyghvkQb1AjhPz0dViHKngQyGa1hAJA+h2qi3dNZAnFe/f0/aFvz
cZcUSvKV/Vh+ZGgqyaWgTokTFiwFhjSF1GIXWNVgFwJELgffs8UEdH5B14S041qak+z0/+HFNTuL
Xdv9xmzmfaQwfY+nq6KKT10n5XZ4XGamvR5DFZ+x1tQLzt3A8jQGFu6E/GjFHJvgRD15xhqkShqt
omehg9VULFl1ETJMWxz0q4knA0Trw7j9Hk4i4jwz8U0uyAcL3fvpHVWVmPaIkLpWEx5ewWVutnK6
MbbFO7S9atwDZSjRVX3U0mN06jeFnhMwI0iXSZtfqyflxDLnKGCXbCwaeu16v8mf1FB/vuYUci6+
gsA7my3LAQbqV1Eyprz8m40ecW6dH1DXfEbaCgbJm0unVq9ars9qhDcqLMAcnYmT4PnN0o7Ks3qv
MYJaCeI9bUrrKqAyXyJq1E4o6DgJBAwjSaUM08XPmzMxbulHiXdyg5OSu8vAxS7TnWVqikvCCMl5
BEQ7a8jdaiDWHaHpKAHrbu692sluAeuRrdsqmK5thZ5ycHb1gKcgcGeNioQSSs1igoDiPnrtWXkB
NAfyzFAWCP25zhOyh827vqT4xLDOk6w+5vfmCeKH5hlevxq5LqCAjrCqywWW1zkAk+zlarJTP6Oo
Pz6IkyNPR3uV94YF3N57j4zazX69OTTkWFYojCMS8j3LSXGI141TAQ02GwMw2ELUI4tCR3pHzfgu
ylnqtS/Tt84KYEIUcUtMnaYi7Z0bIas59DrFdfFnBFTSJG6n5g2vjLyTlUQ7n7C8JS1Jqh8dRRQ2
mBzTowW0YIqH8Z5YE2H7kxoElMs4ehIT4/b8aX6F16SxEpowDNkAaumzEKBtFhz8zg2eUuiG/FnI
iEvcCpwyQ2Tpn7bXwcopNmWW+a/m95OXxvraYnZ4SJOmns6yxW/g7IDTXqIWIh/tcOCXcXj6vRBZ
91JY33gMdbZG1VTBsB/QwhLIkyQb03I6ZQ/jrN9kxKhGmaK6yDMrhrr+jpUDeHAID3KjmWfNQtWX
EnxTlsOanmMavwUXLJtQVeCRdSL/oHJ9KQXCJeM9ZuxQGCvijKnBdbczDHpmWtzaccV68Nb06pE9
dX1g03UP/7ui6XgUKtfE7JPRyVZ3Q3H83OgkJkMfzgKtRAkTpRErlAAN7DQ84Sy7sheHZx5vj+2w
WAVlF7+j1i4sCBm8MeY6RvOsJ9x21Ft/T4Eb/XkhTeabdFiWFsB0hz1YivlKseSo8eiFpkB8TrC5
CywnKTGmR6UCH+kDh/xLBzsx9uPrpdhsn2mifZVnBaru79BgGAh0EPjnyQwtA0538FT7o5sydYOy
vQPiwiBK4JjI53dQY5i2dM9+qTk3Frqw7W/k9PgLoCIljjD+m7N3fGV+i8r/ZjhPfeLnvueMLpSu
ehoEdKBvLN/cKtdppf/tvAGyIotN3d9gDtvJqp3jGkqy3TFVrW+A/eqXXf2PJZFKO8/v0/YX6Hp5
yr9JOV7zPDD4NiHk0bs1oUJbmN3FS6C1B1MDIatwWd8TvqkxgMy4WWC8RfbaAdtxC61M/rY48Jfw
1dm/HcGs8cKUWvhz5hfnHpQWymuuNACBHQghlhdHye4O9Y6hRMSxHnZgKxlRLzEHHX70iDr4pAOe
JZyi0+VaV2Ygq7JR9UmwlSADcMxbvFN5cDpK1YyU0ncaogBdUXqf5CBcDD1D74Bj/ieeB3BvmakC
lOwlhlgV6kxd5kHnkc2crXbhAyAgdrZWfU4xlvfAh6B6aG5j6rRnK9vu7/Eo3dQrAq9OkmbO/0Np
XzAAv4NrKYAkkjuOavUt+hEongba+xbRljIZyjG1lVwKoq5OPqGcspvWE26wEmAPRhhw3YWYnzIx
aEotchPMfapUij6qH8ggAtzdfBDTA6WCp9ryt09zQ/7XI+zYhAg1RnAtTc38p3lJ95zjEoVXqR1E
u4dZZ3mlfVhKFPSFtRK543n1Uo5RK3RNT9AHSPCeWhWP+w/ErBQOizxKaMmkCdcAGg9aZEF/O/Lm
fTMFlfCom8kV+EgfdXWprFAq1o0kUQBHu/NK7AkodPyjayLzrPVy3x/THOBwPsjV9utnfnW9nnb+
Esz91vWF+OfGoJjl4sJdwkO7WH3//aHncfwe8iQhDxu2jj8TZsyERkuTHPoJ5nObHR32qe7pIJ7z
6xrXN3HTfpZ5UhVIJKbE1K+sZALv61DyJZPnwr6Hc05/y6CWcCq8ApC6MI/JqCB81S2DvVJEbhz4
iYP0saK0TSwMdZY8GhIJqsuUEZmzZLSEt6eXel5hFMeOXgUiyFmXV50R0BgKv6CeDKW0F6wUqW5R
p5kxwUPkN9xz569TN2R3Hps81zcXupPPSycpVlbSPfxLC/KWIV8hlK1Q/9AWzxniVnm333idax+a
JhQ6kWTFxzSnNL46uO4Dj4BfZjMD+3GgAg+Cp6oDD0A5oxjnO8s/Gz+5nvjSLxXy6SiymmjzByG/
fSJI91ZHlJ3orJwAOqn1N5B8ysc0gsA0UWHVJ/Z3OWxwktDeDAGKUd9DZvuzxXXe609PcqRHgsSZ
kPskBZRIvE8vUMutXtiYJdSMyfnKQPZNLBSvmtPnioWGQIN+qH36QtSH5jbTlw5EjEl/N/hW7LXT
WZkKGbcPuO2tT0pqtEWXWpfxdIG32ohK75MeGFIpDHPT6HJBGwLHmkVVdBHFJlEMlCqnKWEYekxj
tqbIOEfCziYIYUkDVUHJjJz7SLonclLAWrM7iQquENP/Q/bO3IuUiLAQcq5sA2HX9apKGk9h2iGz
6Am+aGP3UyI5zJ4towNv0yHOnR83sTo343Qroe8U6gQgcvcmWhdOLl6pii3Oo7/XF1FBhmzFG/Go
fXb8iJpAPpx8v0IJDlrBqgzxp1tOgo+/qGSN34c7D/DsqYZ0EwsaKMafRAddiuzJdOu5J5VC2BoL
BuysxtRYFAF0cCt0IWIvU4HxZ+rr/4DV2KTVxJr5xDEx86gcAAwIWAI7aUThKlSUENbEk/pzyijh
xswVnH8ExiDvlQWLClWncBHfufS12DVnaDHqaVAFX09y0DpJds34uthA1aDj8dv6AENRdE+oWGR1
ULbUGY66iS+qSnsefKKMMuPOAov5AG3z7fp7MiKpVUwfaUhWk34W3Z3iwB82n6GP2u6bDODwQrlx
UeWWuky+x8hcO8BQJE292PWxJYONB5LS1jca7oYTluLU2DYrmMkQjOZM6U8gqBjh3wUhoR2PshnQ
vbB8MIaGZPEPPGl5uFldm3f2HCnMksXYM8e51Y8d4GUIHFEds0q/2JNDstzvGDqy6fNEO78cb2lF
wisXdoM5rzMGgq+FCISQqv4sQK9WIDkPcwKxzsuGdSO8B6Bo9Bpg6y5IYGJ6C0ZMxXwWokbcEqpL
h+1OOSaRXNHCzYuNGzBd5oPhnAWMEG3fCBMq+el0eaF3Hkrck2EyeLBs4pgBM3qPj3Lvlpi3CeNe
LPGTEKVrB+hseOaYSpyqJakGV+PYzcZxj8VjtXEhjCMfCS2ICnSUxZiA/Vrbal33uWHGtT91ftih
Q/1Om8ukbrEOqLSSLzj0obke29ZNlppjdqumGviDFw/ozRjW2LkNaSaaVuiAkKetBlB9rlwNVoAj
/3JjzYhnlpjvPBZUBN0qRUGCa05oK7+aJXcBvi6MlOSAluQNUsYMFaCKIP1H71hJMSI4jYq6fKGR
D6VFrLPBmRBSdwBtQynMQyqqG6bKKMmwR7Ye5kTAKSuBXJJN744vYW6TD5G0A0qHnbMb03OY9DlU
XOjCopUWWFb19vHVZBMMvXu+XnIO9jhHZivMqMnwypTNfo/4oTbbxIFM3cQJvJyjLMAVX6ZAXP3P
OnkZynVBMNIINTqr+ZVAgVU132pXOMwjOiPlD13iV2WcW2Oruq/ZDS1jX1GRjdmbx1iR5OpfsYhQ
+vBKr4I2yVp9vHmK1ybkVRHcKKvpsPuTh/dy+LmtQ4nVf93Y3cv7uY5UKdDbxlXzDpEKxGevtEF+
AaAdcX3twaglVip9Qqf9C1l7VLy8GmRDA8LFiout1i7UC5UamPdGrUWWpSP8/aa4yII250jUCet1
6HiYrJdtMo+pPZvt9OkZkS1D3hY9mSxFAQMXlcxcfB8QQGlsICDucSc+Kg38PcmCafqSrdloz4ww
oBkW8ac5wPp/NIcrrsxzDwTL8Z3VMWx+Q+mIZ5aDX4ZQM87V5JVSi0VpEWn3hFRe2yPwt01JL9Fn
4FgHC+6I61sXQaxI0BDIEZ9J9pt+t/BfaZfNsqujjM6r/b+E8YhaP/ovG1xIpTRpmUglJZk71AjX
35VG0RRLwhAPF+ee7m5v8MSjhRm+eWnO7HSPWQsT3jIoS1pr484QtVRipgFQfMkJF2NjP75lgaBj
K8xKj0W10ikX+2OVJEeYTie5ozyXwtbU3qJwPZviLdrMs1dt0T8Hicdoiz8AeEBgZlt5yFfvTeZu
1WPElQ9EddnhFdmuicKsCXUnFFCVRyab5yNiPP2Xwf8Hqj0PrG6Lp2idJ94mKNt4a5VCpObfcjUI
nSPtRVOZ33brHuNrpRPhBhCzts1YsxlUs0OA9t6D1dAI3KSzEhFYhI8K0GjZy0oz6BkTT70jj7dQ
buzcL2ClBjBHg3hg+V8TDvHJWXGruY0AGazvZ4ufCFi2h6XsTVOP2eZ5lALuzoUi6lDFmrO9vz/Y
nCj+OQPDdI4eTNMGP0Dz4pUCbDy4tVNf5q1MyVdTtVOD9jV/Ida8pyGqERjJrnXM0gZZzLE83PbL
A7a0bxrMjbbV5WKhBlF+YVC+n2kMuxnJS7HBTIAt2hwghi0XIhObiQdD3XC+zSs4Hzl4O28GooUF
2g7ckWPhA+utW49S1Ci5W6cGReDu/FQ1HLlX5g7+p//bDkVVERlUFUC14BFJ1RZtdsVOU/YUBOQw
zuOqSr7K+xYwK/5qFOBOmHZKEL6VD+ndFwF8Ek0MVBixIaPDFXQvd5gIMV0FTbOljPEvkzrMj4pA
08DcRzWS1sE7dIEJTf7gD+dUUvseHqPwZOerbYbPU2UTiNHecEM3A6galvAe4YbOfHvmTruuDZDF
iBB2jh9E3WnSDsaKkyyGB9wkZs8sT1HJuslVXPVjdSuVbW29olhUpjb7Gd7uxD7se0GRe8gZuPbf
XA4DBA+6O/SKxh8MiCKmyPrhMIn6sELT+7L8CaBmkC9lXMWbpm+ezswSynUUmyc4oiy9WrjAF5F6
viEzH7P8gLAg7tC6bqqxtwUrCU536bzotnnciYS24iX/MyMXwW3kg5rfqo62sNaPl4/bEbAXsrw7
sJ8lbg5I73oGsXVV78xwKnxgpwpX1B/6534RQr4c5lckYxMBlBSX9Gl2vHhkB6PNs3SZdW1ZhDsK
u7/5qQGfoxy8665JNbfdCPCqwH9HweJ7FfqnUwPCAMJrSUZcMdM78DF0htTOHW801MWJ6A8EncPf
0URfTZL9WPsJ6IOzB8a7vCLTkSS4dyWWdKm19fVxJU5mzwQgfmdiKK0JoOHSifYgzpuwIg0eazoQ
s27zytHw8r4iN42307B0q7NvvxVUyHhrDasnfT3qpDYHeTPvC4cbanmvVIpV6TctWB5f562Ee3vD
8aA/W2BIyyZosTKnNRjCHpOp6IjwUqbul6zK9w7lz7V6Spqr4Wx+dd3fq1Sf3dIR/sBdJnpmJTA6
UU5Svo5v4etqL2UJEVBCB7iwEsrAI3KjnJVTc6+4ZimBRO2WSXps+zFEhc/TzixrCGD7iBy6AxSc
3bn4l2dCh1eysgVlC5OqBT35UezByEsBmsAQAK4YcN2YCNRmDe2KloZW/3Y6NgNY4V8yf4IelTFn
i6ef/LtegL1abJ+SZQsR4Ii2bo1LBEsXABtx67aQqboMLXRlEwfFqjWhl2rGQJJaLWcDqIo/dy6f
MdLEpo6JxlS/ssd904wFWggryrTN+rZc0eJm3clHXKzf6+9INYTj8aDOTB5r7IVkT4J8Pxpqiysn
piXY2eSOfPi4pseM6kFVcaMK35kv8YZcLt0OdeYuSjEDICWHoh12qsM+V988AFzHi6jqF9Yg2XjI
55i6IlkcoaEKSSlhbWdWrKcQdN/eBRiETt/f0nNgfaeGlAtRYUwH+vrkPcZQbDFiuuBZwG5MWyzO
5nAHTwYSahTqh3kTjBo/vN6L7XuzNZyZIdTrAburCu92JtmyznwrhHl1w1V6FwwJ2Aq27w1U2sS/
pIlOuGRcldbLy6wtDiPYtnwYDu1dZeTpJCvuhto8yjA4YLTwYlCG0tv+AW0p6C3G9fSPZ1LiVK8d
UPz002r3xxK3iqfEoXi1n7ArlqcsA8c29TMGxID8rXAo+GCQBAmR1Fg2xMPXx10YA6HbaNoz9T0+
VqmvtGLeYVcGe954ZdVzGGeFUTODh88cbpo5joImMme04xDBOuIvIIL2tH/HwqDMNRuMuvLrItYs
SvtofXaFVG0X+lG5TNv0dU+dJ6QZGiL+edaTxiU8R693F22Vpv8yXJxaJXakhsTc7+ycm9MdMhhB
Uij8cfyxObbUJekxZR4Pa4ATDKuowImq6FxaHLJ2ok1KGvrKURfymaaNbIXYLoyOWhAkLcHqhyG1
A/3rPVEU/EPCV2svZ/+YNFLuYKgGd5EeMq3aTvASJJ4nE/zd8KJWYmBmcXfcSdf4LhXHEozvHehn
Fv45mutKlyw3c078tjHHoKkv1Nx7jHa/YQgtcTzqspGzxtjwKFWHjp76erdnzGf4lVzJoNWubAR3
I+XbJW2g51dbQ3Nv8qzMWMxT0OWOe0vQP+h51C4dJzG/SchUk51qXmF1xKPDuZz77vZ5X2Oec1Sm
E5LtNs+1niNvNVvghIOk1itvEIwU92nCZjTNy4kfygEsT378YQVApMQ2wGiutVkxeJq0bqswsvbe
Hm+qYKkMQjOxWBcnGoxLf0bU7zI5eFvqDSdY+T3IYteLu1OpqJOkRVEGGSJSqhow33xbrymjdzbN
liCgdBIw1dVB7uRZXhEHhL1nn1+OaPwroB9b9kyuqlb/+SOByhTfCt9LjbyWfH7687qofgznyweT
HaTjtqTIvUGFEJ4F60dE/VF2g4eELqZC6uhGSxzseSimCk283qSEFsGxMsggiRicskfk1wEUF37I
2b8Zw4iBvaxGziOb/c86WBgi6vdQ7lHIFLCAusDA4ihyITmgwQitn7pDnuBsmPISK9wtplw41ITD
wwzHe1J7OA5pET9ljJ4HtCGi3ONkRXcOUfkKzvXICPGqR28lx0vOz1T2sRow0d9k77JfYHw+WM9c
3t+rMvQVb8QzccF5qY831njqlPcb5iM8D3YEXtbHg+BTloCs5ylaA25OX335Oa1TYVkY3s+t3Rjm
vFNrzVKxrvDcSNXGLCi1dgtvWFMy3RkcHJ6/nbP6C8+4alAl4I9I5KlUyMcQY58yFMshhqHALYQV
ncjFZ4QD4lYiQO+lqvo6gN6pu9M4HxDYVjRbfSUXlev+cJogI8I/839zzgUKKvqZNSx0paeKcUUk
KtIGUbc5rvRSMGxj83HS1za7nQCwWP17mdc8M5PcD+la4xIHllWpTAgqw+C6pqh4fxcv1mx5Vvea
zNUl7UBedUDw9O8RZxCfOEmbyvz2SwrGoB/1HLnJ3qJBG9+o7hAsgWFEr7X+C997V0IXusJMq/Wi
A7DSn59ZEms1J6phskidR9gDH5zlLUa+cEN/x1NIgftNfP1ORwyv4PuaQ5SuSa/3Fgxd4vSNxKzE
TajraAVjX9U9NRIfVwKiQRizycaXbPDeL6BNtwHtbYE0aLNCZqqmNmyjjGoaO6vv9Oq2BEyi4u8j
TmUmcWAY34iOOLqT7M4DvKVyJhKl8d2CRFbh4apyyZVFVNWRimsk0SpZqPPyXTzd5dKFSpzZpVBN
u8IeCvZxdwkr73XunMYMsGmMeTEB0z+5n45QebsH/nFUL5/jvit4NUPrym11fPFbAJvy90ixHuCR
HskUyFkjdCBDH9ll4iiSWezfiEi1wa9Hz9MwcSOnfChTT3HJOrGHsiA98ozFo+/P3ls5dkQENNaf
ZWkJo506JC9yTT6aHkAJdn7RXLn+iY/nNv53IIK21sore7opG+TqXiXV/vsz9bBOEylx49d1UEM1
VK4VBhr8KSuqMmDdiKH27HNcEqz1CA85GBzD3y3ZL/QjUlFjfEu09ITi3Zs9Z3O0M0fcufkg+Wzk
JL/SUQWPSaJqnZD2zpFT/v7Ab94pG2JK406rga33KwRLjsg1j3imwDc7zBRVF/2vD9lvhw72TDZf
ElNaCYId4lVZoYI7HgPtFCHxjbiRLwRaQfw/nIfRqsBrdIKtPMMQbHIgd9Ag0/5EoaxDBVNJIzfM
pvSkWoLKog5kSbrCLJ6PbcjkZfZP4l4eha8ho8qU+H84099aL7y+MMINub811YbuuxRR/GXygu3Y
aXLVjLRs83054V6mK8hn5TlZ7STRSm8uiWjSURf45pZQS0TAZmkMH3aLf9wQA/cL/Bpk51A3OMYi
VNWHrWPnhsWMng+Yx8wGY7F0x2Js1G8RDjOrsCkHB2izAoMHUibNW5H2uyXbWpBOSSU/jdeT9NgF
6BRJCeKovcy+CPdX7J6cIEvIsddytB/nVhzzrj5qER32RZZIiWDFvm7unhehds3iSgeHNHeAIGbp
ExyBqElicCeQ83Q4x5EKWNGwmduvpK5nl2WlC5Di6iQfWthXWhSuKzq960ppnmpH/WrFkYisO0rO
mdX9J9L+ZjJSIcKK9VzOy4e5xhGcDW2WVMp5RHhgXw1lEh0YkzgPXRYNx9KzbLaB2wGGRBtYTP2E
AE6D550fzp97VOsmsKJ7utgfMlCEq4DWssoy/2ixYHgVDLj5XksscdmNMcYqUvhJ5nLw4xRQaaK7
tB7uVXeaqIvgK3Ar6+39m6jQ6s4IGmmODTnnez6Lygh1zrnyH4EKS49VofEfHeuk5dlgtzZZ56cN
bd2mO9Y2vWLNe/eKa8requACL8PbUM2dkUNjqlAkOmx83DD4cuKhFKALExvp3EeoBPI2f7vtQIKv
CCcI/SHtAge1iYfEPwQ7Yl2QLONeUy7tbSc/yfj9+xgDP5TNqvGJtjIMyusx9CMWJnm9Bo+5XXol
j0m2x3qpRUHPWGPIAPS9NSljMZNWhhcxL1MbLpDT4mTfcXTMHziYZlyKrIDLordry9fgY9IJIAHW
VvJ4EMmfQpVFKE0qFjcCwj6d4Di0pB10Se7OiuvnAU0djINPj+zTCB6uGBB6mVey7AxrlahqDzFg
Iaf1IGxrJzF6bIjkTU+Ct3nY/R6tfQuT/cIZYoHJA93O1+pTgOURgsNnfgrJ5IJA3EQxa+/i/SYM
0W0p3pvPXpZ+H/cWWu3mD3Vk8wMIp1tmeVCxln+dqPYeVqf1tyGWT8GWzj9IoSou6S0Ksuv2W7i7
YAeyqv9iAoStPjdXNGg4Dq4YLF+6EQoNA4kSsmFogqPQ8CaMnx69jR0QgF+KTA4j0ynFcWttg+5G
KT8Rlkqm1yz4sTze3SaFixOh3vSPhEntYJkpLA6rVp7v/aCyNZfVBwg5hzLIUyIX6PGOlngN7Cqn
qjC7nDTuGHAbPPFugC6zutGQh96GmJbYpCrv1TX8xcK4Q+qH+arakfpavXFgGITwujNL5VJrFLAz
KVSUvDLstOxeKOTayGMfALWwNQWnGT0/JkTLeqEBDara/P9+fKp99HGn71VX7MKm3gpKT4kVHvfZ
fl4hyqEWX/YRmGJeJyFmSdCYnXW3zg5Sykic/S/5J1L6m7bw/k4ouEYjIKn5zv+Ac+ELtPoPXPbM
TwmqLtF/keeXfonQuiEYf8NnRmeT4x6eDB/Z4WpSt3mjaeguMUV07nXjJfNp4f3wProO0eHqNozo
UZ3bIRwEysuspOBy6xpMnbBmsc3Xkx8N/ebUVeqZmKuBatLkHhL9JCWTh/4Rq3tdUge+CnvQNoqR
cHBO1qv4C0IGZlJT7tYf3sVV3JY9tDg9TB3kzAuY9U+apjtBqjL/trgugtHM6HMe1y2BsVL+5GXR
pT32Q7EZAFOcEIpJKbMVkpMaZKiludleQYIOpS3piesOVSj6vtfcOFX0clcXUeD3cep3z3STPRjr
GmnLNKXYpI/Q4vEdI7V5+KpcHF1xsSw/loeEvnkwkKYyQGKG2QgJDcL7819dyluMn9I+66EVKlbs
TagUDwt43arhFrBNi4HxlCHWO4rCAW1I2mwMIrnDmLKbl5Dn1slBv1w7znlhoBpNxxDEaGn5YulP
zUfOqtzf3BETZ8ytJkINuxP4lTfLvt8wBJx+QphI+7GDUYpj/K3qqT76I0JVjtVl4zPLKd3ybrxq
RKp0oVcM2y9L+6K9sEheGF1x2qUERTJxVfme4WiYImArKQKFhOGdZussWA8SUz0MHj2Ae1ub+w8f
ifby86FgKzhMhzIPzk3veKDnaj9mVvIzf8S6GWvVrg4tJWs4jp0yqUc9rOAhFsji/H7ZcWqCT4CU
toMDtbFupmtKvgctKcvU8aMSPS8T7hhSostxmAXY8+Ye47Ce8B0uhUm8KGMLmfPNtG6RaNuSqCV0
U5ukoV2Dy/GVqOwWTtwJQ5kKcvlY4ugos/MWLoIsMebxqC2zbQ1T5ptpzn2EvtQk5gMYkF+9VKjb
gZNWIhS+Y8L/UsfYL9+oGNUSdYzKOCyZ6wKWQW9gEIrQVMQ3H5WJeDK0HSslOobDNpEft2zKE/dW
QMzfOZoCPdmAKAPn7uOhtPtWTI15Z6XIVkS2tYaRWEPTfTm819gbRD4qXdD5NsNa3NqHPHWnN2Oj
5zAWoUASUs2ElQAml9kJhkzAfEvzPwrVhCSm/A6olkfx0PmYca0CjZEIInRpRVNgAkNSSCL8KpJJ
0yFq81OIAaGckoVoFlI9ZsjRxXT2J9qvg0hr/tg0e1i7hDDqVfEdVwlSYjFwxrQiEpWVmCm3pQ38
YP90l8lGoO7CqH9uktUGGXuywKolEXJzrX9Ya/o4yXtuSGczYG1rUkzXiERF1q3y+G8UUGca1C+U
iAqtYJbw5FwW2FvMhfeRQJVaIFVWXB8LjTOOR0GXtvYRN0dhraUsd8Wwvp1p+yDE8HEXxgr5V1Rv
MyJ/F7DRDcEiAuXqW6lcsGWuKlv6LD/LhjriqN/CRctapmzSSLTEcYH+Vg6rvxJ3JclFWaBMRoY1
a95Q+DwF2XhS1qTcMosbzipnKWOolJrT924Pyt7W885QBPKwKtQ24f8wfKyLTRzGQvQQboMKe51x
RAV4m8AxDFO2pG6+gZcBnoGj5/AN4+KZWNMXSVR3BN6Xmz+5R2B81vtrLrui4b0zjSITP+melQgt
EZqEaW1qocvtLpbjI2CvsQhKEu6Kn24QOFCQuGR/inzPDP2yHe7PhhcHiWo/BroxmVmTwBz1qdl6
PXE1bYByJqtoiyszm0HXiEIfM81ygeesSrBAwESpiwn2T39Vy6fxQctB1BCwOZZANNQlffsVkvV2
zxxyhIPR1un3VqEvexlx37vu8N1lOM8LrQmV1V7R1jyGDStKSwhcYb1FgG7FmIbkXIwiLUgU2OA7
paHyOZPN9vp4pI3vUCAZGHAnfKENXy6MV0TCNZeQdCQkCC3HEPrZf71YXCJZlnMNi72TTQdx+G7Q
JaSdavzai9ZqF8Ik5qPDkQZA0zPTHZTfX0cnEAXwXZmgZnx4B+8ovJMRn6wCDfRz9h4aCrtHwU//
fUF2s4T1oqe38AnImS4LA+I0xxJUT3N+WkjtaTp7Qq41mNt2Y5NUf8E5cibmh6gMgbnuQQG6VBtg
Mu70duNwaSSPBqzUr95fieo9P/QZLNfSIzl0E5Gz8zz2cF7d/WVCMQNhtrposFEDmtaXJnVj2hMA
xqDy6RUdDEUPfaOlNUy89BGlfjSbju5ckUmheRnCNOaPy5/rn6QHEj1DZLkd7G4fq3AhxceG6gp2
q3AxBQbvfPHpxEO9yDUvG8RjZacQkgUuQu6nkgEyujEA7QtqgVmao26PYpIaKHE3rklry5CiwkCJ
KoiEVf6c5yUR5IZp4e+k3mGzwUQKKiD7f9fdmvwUUNt3FKy90phzMcbSUuuSUGHhWzkwZs5gYjNO
L6OLfmT+wIA+pnVquC00p25ptWpCwgcVsm0yEZ5icMnj0DFXAwLNfLVNOfLEBpo9BoroZgd+LN/h
6CzaM7R/kOvWAqrRHUCjbLYtVVUP9LO+4zFeSQXGfja2BubySpYOBpcRT+OvEkFauuSnqWjKLOH9
BZtbiHkC+nFdk6P5QcLpkFGytpWHeypCbSph7W2r9Dk5mJk6MKvgX6mjhW4sw9GvYIjrbl0ZrVFB
fYogvpHKm6L0vYdZA4U6kVdhDpfj5rx5FMObRQLGXMCpVIhOgKKVfuTW1sKcIEsQmYZIJlF0/K31
ZIjltj1tZ+1P6YsyHTV7rr31TeeIt12ckVj0R3P8bbblFdcLRitfY/dkp6y9APcnLp7qi0CZiRxW
EH8oceVzKxo4yaWJ4mFCkRLSd31nD83AcqdAKmhDdN4nH2Pt60EF8RI1rH7Lo7C/xV/mwQ2lVhN/
3+PyhI7CaIh8tw25GbfZja1+4gZWU0W6khZ5Z/5FI+kDKqrfhxKHFl1BXFd3Uom8DqD5m/vw2y+3
gJ1Nr7l6tg6lGSxDb7bnxqLpXHGCQbwExqzWHUfOn8M6NwYS/x/At9oUd0QndTtsF1UzH3nefRRX
wJ3x0/4SsAb4KHOOEdotb/MMUXcve7w5O//pY2l8/sm+/grbpNv0CrSIz+yptcMQFoYdGw8gALWd
UucGc4XNLFN0Xu6TimraHCzdpUUMvB9OFX3R0WK0g+yZGQB5MydiKh0rpcuV6PtCy71+09rt+JvT
NqqOHKJwcK63S9j5IhGFH9MepAExOZkCY9B0ZqA2yFZ1Qe21wUe0Q4X346eF0fujmhkDKwQsdq3U
YrxI1GWYovCGeXHrQL4B8O3/z1avQpJ2EfvO0k54e0AynVOs9/2WDwh2IYvxqDIZHXeBGtnkj9qn
OuRJUqn5XuxCoASjb0eZS0mblIldLbpJ64LsmHTSXDERwrWm671Ckf9D36YGKvVCCmPs6i5yZlQ0
wecPfjYbHidCB8sitiWc4pLzY0a6FxvMAwnZtkV/J7Z/cuYk3ZzItJzb3a3s3V0BqV8Oq5Qc/rcp
FJCq59NuIxX8eFoQcUNAdd1IH32t4I0LOh4EVhN51swzzCLTm7VvQEwA49g5y4m9CtAEX0sUUdOh
xug51awln9/tfyVWoYlzcUp4SjN169EjPVUuLVFDOwxdd/ApiGQlr7qLvK3+ABPNBMLL3Ik4sgWq
z7RZmJS1EXWeMvYkGgpsJZKzhChNxtEKZI4BGlHjcnvRWH/keZVWZofh5nsHzFRhj1UI7/Jra6Ac
CK68Lx6wgQwR6mw8DEmLRnrFt7CvU6eceWdeXONy6Yk/XpYuBMgrxHYS6f7jcqr6KI5b2ev3zakz
DnetjB919RQ70Q9R/sjc7EiVoQRwfKTXn2wVfvXEk0MoP7hqoEXt2Co9Fh3i5WsrpIqPtUXgjGbm
w7WI3gOAoidcxZMd3S75a2/Kn4a0/uvXDK5YMnYo4qyb4WpkELT3/gk/SeZzccYJoH+z8em3oDBQ
LpYHwEEfjchdiEEbKQpi/eyrg7cYkeBkWZ7u06v73SxictunKcRCOLc9orpwsEtZclBsk47Pqity
/VcZRisOzMN+unSSZfNd2wf/uNf4qUoBRzjma2/pZuR/eA4FGE3CQi307mI2xRMtVKyUU4dhB8KP
TrZF59yaOCV5S0cv9R607HCwP6TtT6WdfmYR52jLkNLH5/thJK5PbRNaGiQxLgCFAAtsND9bLZ3l
oNdkmcDNLrEKnHtzBKC/ps9yuT/Q6IwGc9e6jlrauE0/JBDY8O1gFClC9Z2EH4ZEmEW52EWISpQZ
00fxeHwMYZJHrK/+avEZ/fDl+XaEiAMm0pKJeKI+q72vvd4cBJhz8fUG8Llr74x3DDmqWV4Gx8XE
F//SAMynb86MXz9BBJ+I8LmwQKlQng/RdoAWcvZ8iwmEn7hgI3FvNnBLDRKcDEhBpypIiCSSKaS/
rFPXk69VotVRKyLh9S/IDlfc6u/7yNB2scym/MamfS1WbstUVxJ0yRXQZW2qBqtZcQlQhLTLsaMh
shvCTRLC3H+JaQ7MdBMDAtrIW/rzKXyv8Qv9H+hFeUZMjn2w0jBEsN5+wEDJSn4+E8yKul1iWU08
V1LOfJUTSKvY9gqzdv1q6EtOTd16IW57uM37CB+N2oXzeTDkRZ21pJZw/8qjzzBvxJ0aHIAwc3/k
nV8LzsWDn4QU9VEx9JMU4lkb3k9O3fxTU7L6bpSqpgY40FH7YheC9cGh8/M4qT0bsLzYA8vI7I0N
gYsiAZfY3SiX5KzqWxoSyH6qmgfC3JXszJ/94wlYaHslKgbDevRO7M/9shd7OagfJThJhknnM6dt
2acRnjY/ClG/HrFN5RKrvC3e7UCY3klgbY+F9FnUWZ9gdfyCbuzCFgdOomf2Gpytp0HXVyFeaC7r
Gc46yZ7HBA5s3FJeV4mpRh4qP6Te6FqJJzi0km7aHO0IEezFERlFbzMaHAMv5LoQyq95p7PAYlx8
t6xK2/vgRhv7B3RswbdtSSAhqw/DoR/dtgnw1uSVb2JrK33K/KJM2hP6YWRpXjjIP0/i7C6Jzr/g
Vy1nLnn3ZnqqPKsN3MclwFgI7aA61kBRcUQQDMvSTV7Zvn3/1qzfV/cUZuTKFl9DhtJis/s3WMoG
86UBtS31CI5C9qBwBdscEWTP+8j2aNhPZwsG5dfgEG+m5bb1xfXjUJlbomtxXwZ+Eoz3uUsDGLo1
pNJz44UteZfryHRYLhMV/uETYuiXAqYxWHvDcNO/nvFZ+terMePacCDkdx3z5dLBwewD9JhZRVdW
gsIeEVEAVWvxYHP+8LiTrQsgIHVFbvYDUiCWV+WCAWQrq4G6ApL/U+3oCR49yyqHQYXqDb0bxbRq
CloncZNhtw/YRzX8VypWhekMDRIb9cBpddvak+2AS0Zncagd1uS2mLhd+L6lQuJZL1OY+TqsReTw
giIAsaQLkkfT2ZxigXxVg6Kk9ESEqBhMhvniTsKSPtNY/+Vb52jwvyf5cye1zb2R9JPUigSl8GYr
tDYB5cvKq2yJOIvDB0DhM9v6q9g2d+a9BMBCWiWWHRPuSdsk2kChxcS91T57D5aKGdKVkjlaangO
Yrp8C6y1iCpCCUatQkI6MJmn9dBnngNYnDBEH02hgidIx514k6rYfWiJWW/zmGYjbeaUa519rWlQ
1xO7rN17rgfYCy9SfC4qCC5xwyueo0envOIfN7WqIX8RXZERaqaCYzqYYCmq3EOXBulCKn3hekHP
s3IvN0R3BMr33asOIKYJ0xib6XjeJPuG2DBRNHOaHEGg+zCmg+YBdPw48HaIWqyo2jcJUSwBIWlg
cpFuEVhzOU4oFUUNc6MWldFOT3NWOK/odaw2V5BVg/q54/Zyn8gh5JCF4rdh6fBvMyAIyElLM7eM
Gb15m8c8owOUoeAcScTtZEoGaYO4zcDLIhFUSNzeC450jxqRb2qJDpoI3xe/Iw2HekYQnK9xQUlZ
rcMzdu/Ee6QYmQk0ms/i89kxRz29EAikdYzWQTjnQg+V+MkwPSx4xie9lEygezddkTLwmf5w6DyD
eW8OK2PkPbzXzbfsCI1aMMQgNk9Ma6z/lOD0ddsICf+VmqtkmA2YFtGRpRPKZSEPLk2YX6hDUxu6
bUfwRyAgBIcNUAbWeByEw4gWmjvNrZFqZgmkiIEQZJrFt7Hok0Xf7ciJ9eV6kBZqh92l9hTP2HsZ
XGqjSVqLHpv2IGToHqV0pseCMAHe7Bb02LgKMA71lgAC9tLnBVOgN47IJTPmQg6mYuLMf+PW6OHO
LeeY1C9Ug6HVuYu3SjdUF754obeNDXKSKqdWPBmPFoPK5XCBdse0h9NwyuDb92/tHXcDKfifAdJ4
dA8XfzOX90H0SqO5x2chQkUGpjCmVvKazXw5YclFpUe1OiMcApT0bVTmZMDHriDsUD57eJu+md44
f+Kpd3lSLFWxNSvP/22D9Qi25YJZit43S2D2+s3OzTj98Yx9oHtdyoCsdgPv9uj4TCRVhiRrUCNh
QTUxv1lLP0Rk42hw3U+SQ9Dwgnif5JG5qeGoQW04ltDhi6LRyAhxB3eBk045nQgimZJSax1vkmH8
KSyVn3AoZUvErK0XwQ94d9biHlQywTrsObGSndGeC/EX5DmhcfU3rfg77v851b2VRIKcIhoa0Jwt
CBRuAfqrFhBF2RnqkRTf0wdcsx2Qz5hWV2blpbqp79pc3giILV3stPD/Zb5zRcnDEmoj8NEXRszT
8wg9bqXpf5Ae9U5IGAtL0+CzN5kNB76H1k69MARM792bnk4OOObUfWvKsJHcf+9Bfm790RJzyLFZ
ks5/ws3aTS//sqpBFwI8rqGLuPqZmcwSI84cL2q8QbIZUupVAr3UZsWvS8owXUscbrlBG6aduqM1
MLe0RxIWa79Vvb7sReFLvJCn8gR5j7a18OYXxd/kuZ+CPXYQ1vh5o+I2anJRWcQ6FQA5F7+hdc1k
B23v2RmQME/8HTeMtB2RXcub/u/3pCtUHMURFevpJc4ZoExHYWnXteojGZNoNGW60gqT4hSOC3Jo
hKxVTTKHrnoJMltkD+16xQ5aLiYF4X6fbmOPv51TQ4o2T8Bh3wFldQMqEG10wz3wJBhKm1ZBQ2N9
WiDE5N1t9acCV0ohmgrWZA3KljCirXhUpj+twhBTPatEjRbWRmOG21JFQX8tKK92oCqi+E+IlTH2
ULE9ADRENfr7GisHfC2Hdd6FMpOSltEjN5f0Jvo0S7RC3rT2cU1AQTFcnAzMvbscDVHYLHUwubZA
by2Z2Q/l6D/UL3kt8l4A1wJA6rPh2p30USXpfuNLs7/t5ZXUPs/bh96UqZFEHCp4woP99fUe4tdy
qyG7/Y5H0P7s26nzfwuMFM9IacVnoCgZTL9rkPXsT/l5yKwNpnIlSCKeMvPFcW++td9J0U2lMhpt
VdZQKCrFnFjcIuYWoJd2nWpA94mdmIBdzbfMFs8neKNbRiDuhxyWtFfZ8Fc+AHCij+5s5ZfsC4lI
3xF45zERNFE9IE3tj4pJ92bzSf7CxNBmWZuXdgKw6qVLCsolbrj18UsRb/UnaItN3TPayIwtbnEM
fTS2fWcHAijZ7I7rglDMGa4U258P2VMREedROM0xGcuVnEPuukuumsxylPGX1os9dT0CAU+ZOk9S
o9yCqXzFX+hf1Qf40scy63l9IXjrzJcype7gLgHno3iAHNs8E5m3LmccqiDG/z6HHupfUJ5/SuvR
XD1GL0iMv3wi6oYE5Arl/uue6y8nfszahHivPhOGqB+kjiz9HktGPRcNnEZ2pyqT2yv+g6yXoRpe
GaSFUJL1wEiybXusBFAiMQsDCOh5xhO7DlUuR0CsY/4ZpZfGlTeFawUCe6bihNznvlcHzxhmL4pr
kJ4jDDKf3vL/SdKISNqd+5txrjYmkZaXLlVfaL9qDVqY0EXHcKsetpthZKvRuFDckygqrfYBVZKr
Ig2y6wGuQUSJXpQNNTSXzb48bQadPXZ0UNhFWpmmmHBVDhS+5afoSVAFGaKlJxp4YCxt/1SBd4RL
ZfwVEmZW7+zAmMrKKK2D+YHgaT3F8vx+EZ4Io90elBiaSJdQyMv7bW+mPbCai7MI34IIckq4gQ1N
836Sh/hSzz3LML/WEq0HHn0TUyRTfGdQK8x5vkL6thGXqOUXuFsrfggk4kj8bK5g7DYwyanmeJj/
cxmZbOi5EpxTr7j2+4Km+hUysIcZR//BePCU1elxy7DRXM+dzx90XOzD9W7wO07OBnyMsS6FUkRR
lIZhlpC7y4pG092XRLF9vgOdHjiKt3mSEPuYPJ3LJGUOpkTKcaukMnrKRpGWaKFbhZJt0zQBDoyJ
uqjyfgoIeNmaTLChTpdGyBkZrBm9W7WuPxV2ed3Zahppggsvz2z5Yl1JGxlpXpS0RurtLgwS3SDo
ukGE+drsfoPkVUP6F/y02gs4xv/8SRacXXY6SKSsvpfjh6g/NasYUlKiIZA12iFlMOFk2FB4py4b
Inwdr6kI/eGYjlJdGRxHF2EMHnPCRN0h3XgqCYHS8JjmmVrgqU7ULlUDyWurSDxyoHKX5FSiEkra
BhMmrBxnCi0J4QuebNK4VWRq5yR1dcoSFBrMzX9iC5j+yNyO3GswAH67k0OQ9izpKJ1jPCjNOMaR
fNYZ8vum5iDtn26Kf8yn8lYIOBYxqauZBGr/+pRkptm6OiKRlkzp2vNqgrbbgvps9yRgIVEz7eEy
d7kHahrvApuF/3dSWvC8+1runUapreDRrQ0qgpoF5Xg3XnCaljw6bls2qvHAzVzPdz1I0OFcgAWF
rE7syoA6Gm3wWMpEjEaJ9vRQmUhKINOgIQmYJr5SS0ucYNRtPgoqpyuClE46OVeEipRWi3yQ6izs
oVrnicKjDn8FoKblmc2bdSLc+0s39Lv0MxNsfC8zacErLSC81Sd3xamOZNAol/LLgoGgHAitWuIS
NFd5D9tioyNWihTjSjD+GsaGEQUidm8rXwTamcsGFETm2hqI32E4q8gr2TGGBloeDdqM0/HtH7vO
f17XjziN6wqmd5fjOoj5oTV1aDjoCPIwExMkUzbDYbjCNDGb2LZUuqi4rT2eI22xRGfuAZhMrIQp
zfdQTMcEP4uhpn5fE/bzaiQ3MG2vkg5xafdzNiT0WiIUjDO1/HcLSscR3uD2VUdmexapzvatWCJg
H1d0iORg9CFIPe/ttxuWrD0yTEeoo5YrUSWHLlxNOG/WqNd04lwupoa6nkLvsF1RtPcS5XVUTRfx
2cW8a55eZZqzgyOT674P2/xoKcPHqttG7Y+P448VDo4UYmHY/8JqxB86bMxC1XvP9bTXrMrz/Tmf
yzl+FVBkhdjG/ZGIH9FM5Nzu1pt5tY+nAdJaZMlqqUTKWJnUDp0QhOun9IfMSqg9bVz2QiDav1Df
HGdm6lBQZJq4B9E5tfolvGQl6ruVqFCRvtjlcPEPUgoUfmgex1MnGfNRzR2EOyhdA+WHOaIuQS6d
AiHQED++o9rSGJiWWKiRqON4zV3e1Ij69uASRIODPFDKGX5IP2yOPSUQzjXM9pJsW5qnBQB7psi7
3dCSNehYZimQpgluK0o6C8r4WL+brcgB3Ydwxa3XPV1jJnWaZc6Aqm/NQCCsn/oSRfhsfShXal5A
wCgXaM8bCmwaMnlPCezr+e6kQOPwSVx5E2nCzxmyUeCi9NLOwSNg2NBjIABjMDviMePREHKdlaNh
BkByWNaUc/gYPrcfBONcexIJz/m9Pyy4fHNh+LyXcqFSanKPaebmRan9ItNjU/n3hZ8tRKSp0C8N
ir8VdwG+vXK+wkMQaWsz6g+v2j6I1PqUD8VBaIaKnzzaTQV7zttQdC3uwa9gyABnGSRNlKSGPp1E
pSGMcXOzY9JQ7HXLU+thli4jVM6ggBmK8/5CEwndf1YAq6tVHVdrmaHTcB/5/RpO4oPC63cFekG5
MWofy4DwkAUY1gyFJXAdhW/3fPyDxzRHD2YdknsOq0gI2dhxU5fJGGV9zNS59D/X67f3wgVtLjYr
KEnQmJKWUCN3o2IkFXKxb/MymtlsfEuXC1GIRHceet5PLzidiK1jYVaonfppXnBN8UvWAGXSiTm0
2Eu7SrESTfpcYXl85GUDWqeMKwOtE0b02H0G8eLXFxKYTRimud8Mxpjit9ENTZx8oHoRZvkXAzvF
HgSN5MGBjgDw8dhNF1ulsiCdUGDX+Cpd3TLC/Ie7qPVucQaV7KJnsqIzAdtikE3hqn4nUlpMFpcf
d4ZlhAEK4DbfH9OE0LagRrpUxYv2/ZPA1ilUEbrePSmTqqik1agLt0sz/U1b1jxgVyBGoq8+x3R0
+OFHC+y+Nb/tRSWrjmpGFFAoVP6QVVonzuz9xGZUq4fAyTyFeJwF3M8Rrs5uOvYWF4yMMZrpr6D7
xFDOm8+mzw1Eo6A3otbSc9K1UIRWm8NE/kKraLhS2xGvIwxcu2mNrPp7GMA5ZBNGun4NC8zOoALn
oa3SO8zYpxjDnC8zCYEot45LlrGLx10GJN3oK6GmoUTrE0n0tA8H4gdWiK968yddre8fIaIBFIaL
5osxgJmVKLme6chs5Muykf0hjfr3zeH28+EI27zd7lKLVENvrursQf6l5FXKuxqS2ZNxGQmFWEG0
HIcGKlRHH8vX4Wn9rq/84BEGrPjHKiT1YaDRh+5zKUBeCXYwZ+BZrzOqMGTfDcVoFeyECrYXLDd6
QBdbeGICldZqvwE58fGTxQbsFwqSqbxR6t0n/58tr+2q5Dff276RJG9Pk0BZGb7CYyDpxG4NH/I8
yRKR+1VDT6iwAxp+LddtqerBjpTvl88N365bYr5+wMEptN9ptxg+mjnfcJVJawxDke7NHB/zNOn3
4LOyk0b5WrsDHWEXwu8+B7fR3EB/2uzHI+dDsed2bK15nCC2GanAUVXqUQZuPux1sZythBTW7D24
12opBt+/A2mtRddzBjDW6GoYCorisM/wY0zpiT/9KfELK03HbMl2gYhLka6NabsDi2wGhYKwaBNu
YgVW5TgIjWV6aBZ3LqXcQHCF25BrpBJ2dZZHHl2D2mep91IZEKP1MkCmZ3WxwMsaWjHCpSGvJiCy
Zh742d7Fx9nTjEbi4eJcVQde+j5m2lbT2c3zwWgxEmDVvXzSf4cfNHdlSS9vVIM09q6lDy39hAPA
IklK60oNX5kYzH2+CvKCOMDRrAyNvDXhrvWp45ZMdZMrwQZA2zEV9Y68HoLSa9Y1uujiimuU7xIQ
aGwn26N8IsxDswJ0FSRfHOTIXN8qe7tfx3B6wgN1XGA0HdxnaS2/qiOjZZN+1Qlbc1rSZuvz4jzx
U2c2uODmWnVV4bYQHjW+kjtGF6JGAVKhA1vtb/M87LRbBI9yjljTFeD90MtQmMjJcIMv07j9STzv
/DlLeqKw7IGlMzN1AnPHMqcbRJKEDhJaig8Ux9T+51OozraR4mlEQZ5CDELjq1qf++Bj/Z/FFxNE
zLkWjsr3f2sQ6viF9VgcAeLDtRvA5W1dZyhGhrF9Dhl8FHf4eNXkIkzgXzDvC648Krmx5VKKr18G
riNB5QwXQNlsk/QpoXRDBEywf9pSrynXLOCo961LOCZamqKQm5ExwRq2CvQUCjqwyc6kYSkYR+De
X4p1YjUMI/5vDPtYsZr+uC2njuUkz2D3OLzC47kt69y7sB7jEzApcqPdKvJ20W+YyE8KeTRvv+6z
EmGm0ql29RfnBg2ReSTdMpRqhuJdCqejQ67NbpNdE9MZamn8lDF04qcAOxuZpVe+iNNQrjqrm/HG
/6ZJRd87MDqfhqrw3c14YK7i3lk3XeU7se764vmKVj+rASdQjXUbwwaJzqEEMcjxdTltFcPGmWc1
4thVScavUC99DwEOk3W0pAOmMnfhMO/Z91R5TLVKQ/jNcbOb+f5xcFkSgfShzOtB02orKLhj32nk
q+u2gqaZu0mX9zMd/XTpLJkti2KzohGcZ6w7ZC27EJyXzU0fesfSekEQTqle0r/ai1uPHWciWqVS
55Vmanoc0e1Kyo0Kejt6vCfKYf9Vm4gSRPfVFk8GKpG1TwFjSEytMazQ4kpIo/LvErDmBLgVqBgg
aTn/nnuZXa90ttIwNAelghCb0LkC7npNG5gooLmKOZjGPGQvpXpwVEGrytLIDfqd2WAFF8xxXCK5
LZuuI0EUN8Qz1AQFSU+xqyehZGKPI3WQ6c5Fr2Sxa8LaS6Us1bPSrRPPJIWNjoSOyVeVUutbu3Vv
GD6Kfsr3B46UjUCMp6WgKUKX/rELvzhX/V0rO6VVV+QUdqh7PPQzhS09ZFjguZ3KvM7FMEzkmiEQ
a5K/Ki6Xl+2SzItb1r6iF0KcPHCh+Q7UrmTJCFZm3C47El9Xaq7S/NLjxFUD5nDHjjfKXKaZpumY
miHkEBF0GZPTcoMRsB1kECFTTbgGexzwg/Q/L3+3RpV1KHZfILTzWmib4+Cd92m4U4urC/FNHv7D
VLXIPXfpTwA5Szsvu6aDLcFDL5zswT1ub9onXRv08yrxFRHgskT39EbZIAkGSd+O2Zdvh75ZEAEH
0BmySG8y8FrakQJxgQiuG1jQ7rkqmPDDQrdgOAS3CTvf0tsRS18JDqUCj+EROdK0qv8k4bayAiQ3
Ub2umdopQMUqDI3hqxPVivuGxYM7MX+qS7v2f1XWi8ZOsKlRLmwz3VsLPcNH+YSpWLOk5f0lWqbH
QQdilvsbAIFQV5DY8DEKfFR4XjzpX4GMhwMkjOfNrhPzopnMtWP9Lq1+os8aPkeMiyvHhVc97Db3
aPKG955/Jy+akhiWSPSBV2F0fG5JSK6p4SX/ZWmqRrfHM0zUBEuJWkCzExpjhYWn0a9x6dLAVd0d
M0KydLUaGrS09KZ3EEaghukyKv8LkG1nRlBJaVSpZjilCy1R4O1I/YIZP6ELpWumnqPKHFDLqjrw
RuKmDQ5KMC1tgZRCrk2Ad4+njFkkohj3Y7QQfdou3Ks2GDfJF8rVo3vNqwkoGxyJrXKee7I40DIa
DqcOiDl+oB1JVniZyGA3NqTxihVL8lcmBJ5/gywQX2eKEF5GurqqFHVJzCEs7tsG1kb/EKbLAKOV
uJumVpQ75Ym5xASztsFHD29L/tWwNTh+24UGQmmfHM69en75onm5Tyt+iE9XYYstafyST7gawU0S
Kcw3rdJlm5LkALhpq844YY76NVRmC2MkwDh2m+gYwAKGocGuvF01HagUO2tdotQqHYs1lbe0EKAY
lCKRDiMDoAfUoODatyYzeg7D9+toBR8212EMgW+UJ5PK3pOUG+1TyMeR4DnXctB7bRJvl5Rt4C/V
OPX7V+ciQ29MAFys5/nhukk7rE0Yyigfh/Pm2/FO6o1PwGCrjx0VpFgWpqZJBWRF320OBxVd7JWA
zHl7WWzT3ij1tfkTKxiWhqkbk7if9HDy6fV/Jzb/Sa6Ksu+TQVRUO+axrjeHdf/xLKC1bt441WaS
rneHJp3HhLDQYgtuHVFEl+1ta/bTmnVstMDrL5W6jenOv9W7b50EgzemSsxXpko5uetXkiNnrkwj
4Y7Nr5Fsx4H/xNbacl03NkKISDG2xXcjCuw+GrfUputYLn3uGZPlVeX9y/W9mAyFdAoKXpeSUF/O
qUk41E0AESa4A0+iiul7lE260T0cjhA0nOjO2+r1WMsdIWLZeDsMzhgykji7BWa/2qi16FXs9Y9c
0UUC63q32hdct4n/Nj9v/yzdrIyuz8kyzX2p+Sv7ZUeyy3N3PFRvk/fZQWao8rq81SvEjDmEDEe4
B+5Sje+ivE/LkdjW4nSxnUozq22PxHJXVv2GrBWtTpU25SjAwn0OZtc1mjlQUXs9bhhuTN5vRl8T
WPTK4dZK4ENdF0ls1FyEBrK4caHTwpu+GuGfSpx23nHU9hFEuo3tZEbXwIjNUF/m62vbGDJNWVZR
o1NFcsGH0YaMwm2arnLWuasl2GGO4BKvmacNeTwDa0RV3nQUUJBrBvOIHmHzRwK25wpgahAuQlBN
53eifYfx5vna4DmsD06dLWnS4P6Nk5kv+xett3UNFjF78rmJ4SEP4CPUr7XCP2QEduxEsV2qvjD2
nWeiqk0xxpRvPLE5f22aM3Ip8c6voS4jBMP6QT3ujkFAUIP1TETMxeRXa8hte0symNldGKYtslQC
KayYJE9rYtOL65xs+9cwQR0+9QR2NFKolAQTXNXWU07L0jhRmqM3DRCht6GYQG5PPF/oRj3UpdMb
BgpqXqZhnPkV0mjYk3SN9St90URwYR9rXxGsBMycRe78Ik1AWqnaburaU64gCSPBdko9Bp5HPaSC
eONh45lYihy+zdLBrrCiEyBl1zQ+zYt5veaKZxu4IlUEwSPR8mW+cWayMSCnjRgnwkBE86tMfg97
cHNmzdzES6vpxGcakN3tcJjwdla8JOJBWJQAOBCglzcUlmJH2oW7b8vPF+a6zSg2hR9fbv+gB+wB
Usaag4k3Dj4Au1HJZ/Tl1RP8pvceNnf0nmWSYTszBJEYqZZaSjDruwVpNjd2iX39RE03sg0JlNju
OZA65XP8yJM5cin7j79bBt0k2VE9n55H69aOBi5eQ1XeOqysU+9SrdZ/rnQyHN1wXbJCurjoIUtJ
IRqm5vjkLoxu9tHXT5x1ZLZ/iPAgA+bh5ICONnW7Mms7Iroy1kchSh0fwYOIW/ai5gCKRdp3fK7O
AAuwTejIHhqXtru6xtgHHfinpFVjaR/jZgZIZIOFQfJmcoc9jHWklGuQ8OkircdMqCVMyny16YFv
/ekQ7aV/5Jmu4KMIU5IuW0TxC096ARfHjuVTgHOQ3l1hJSJemxvrx7lxMPfBgZtkD28zDs1pSi1p
cda5TafE5u65Sk76yps/cg9zOatjiTyHT780Ey0WTMAOxF1/AvL34Ua3ZZ3ec1WPyeh6MTQ7IdY8
WE/FD3Wo0QJSerDJ183MrVPdaTSKiNjfePP/F/k2XfZnqfIvumpgf4oHMRhmvoUicThaJzLcDS6o
xWpyec6THw32dxPaAANNB1U5QzvBwNIQ41HvrreHBfMKlMPTzs0UU4BWIKIzsMDckbzDzuF82pmA
uBiaBI7LP5ClrsL3slTYL9LbbLt8VeoH2gpMsi8mheBNsSckIP1bX/8Iqbnq/8MJdjFVGDu6sT/W
RMJwhIgXwgeL4wq4BE6+pyfdxdmkwkglkPCnvpejPescqXP8c3l4Jsjh5KYIN1ilNjG/t7Y/Gl+w
eUTmYr5vw4biZKHvdmlaHukCliLIQdTXBHo24GlZP8xJ0pZT+GgaWQa/2ktzpmbw6WqeIyA6b85Y
9tgeYNlOry9FvID5FpP7v2iUuSmFQhSCAzF9M8ktzZ+/N2LEin2QIyB1mlT1iMdsHKMWjSF+CEQF
y7YArprA+6GS466LI4MV8u3vNFU5SRzRyPzEobpiyJBYP/vUuclgYMfnOrL3eNiIE8PpZEFLSqsE
m6hbMZaUjswpHNGHS1PPyl7RBfQLJJgwTU1my+MqVUEgUe2za5OCVVehT+3cpLJXOi6lZepGYC7D
mnQWqeDTYgnaQSV4e3S3+ZO+Ii6kCNKjEuGjpEUceZ4VZR7hTNLmluuvwVgbXn0J4oP+90UHqmpi
LlisDrxNQy0o+ONTK8NeFu2s4dr9zhgqgOqVY0VSae5A8+yZ9Bz64YY0rQ/o/MUClqZMIOtq2LyB
15D/WBJoz967vOD2NK4JDE+X7DSMqrIavJQiSMhOGjeezy3ivKYQq6TRUq0B489728PPG1LncI3j
LYUk9Y4RefNBN4zff/3jyURUUru/bd8CCpkIIADuSP/OPbo3hrL6lvY/+xRwToB38WTa2hcJSyaV
FE5SdkFTImn6Pmvg9PiA4OF/k4cGF6hEX02MfZb6xI4yGHpQQPGsOAWaSlC/lqtBUmN9s8kK3Y43
7FEfJh8gtn3tqUc3lToZ/qNHO8GO61gUvvqYkwsGos+waf614WE6/4AybOMX/6X/S+32OjismELh
UWjoY8OSRSK9zchXschNP0Rus9ddRFGnUqdpsPPZa/OKFRBrQBE1KzmvBPhz5g7Il5NV8X4F334K
wtPrQd3L+cY0kuelfKXX3MYgeQkiOvea+oyt83oYltnvpcarvu6nCMbDpZjQ8d2Qb8FbGXYTOEMZ
Vee8nBe6Ck2d4zfimY7ja2QiH3mGblQbpdYyesmcRV+8tVYotwDiEz7VI7T0lLOC9u9FIwiwB7HP
o6Zb36iDsWRg5UxwInHACBSUEM1XT1HEciow2bnVnshx+zXkfZoem2jV0c7uJXni0Ca1IUf6Q1S/
Lq1zKUf2++zXPZkKngG9w2YawPUYPxQg+gb+yQnt0LD0GvUPFJe2M8N0s43O6y0m3w3hgJkPQYRe
ScEu527S0/p2MLtHmvxxc+jxLy/3ExnodXshIbegewGjoX7BPv90rt84gVfJZomk/YypmzGiY8LN
FBAKRK4lORUTaajUvNg/8qM5cVR6SIAmWFh3af/S2qJrA/pt5wpYBi4z+dG4lsc7izSxo/8oHQ9t
+f14PA4R9oV2hkKBXqV2hVNVkasnIl51PcYitc3c03CtoxYLE02T5B9QlGu+mNoWKzs+/2sR04Qd
fi5iBJw6DHXdAs75g/mHaRD0EINzKHbiRMJ51UN/tGEIkL+8oj0wpoI2B8valV5WECzqzd4GGIg3
HXjoiPrDX6JA1JsJ7OKgejQEvP3gNppO1pEEEYMvra9VVcELgrbirGtFNw1AwuL6rU8OJOtV7oBj
B4jNcSuTBF/vTSWOlQtyBA0WZ71ATZGWH94Emt2mquHDflJ+rKhi0FSe8HCd8XAIFOy8iSQmI31A
6tyzHKalFTjLBXIQ9gy7QStCmc0eLlitY003GOq+i9Q0KMIV+XYMJyi77vzzrcb1j8cEW3xsJsWz
oUFGedlFux/587425EwYbKM5QQQZbNPnomR3tUZ/QVX10VQ2BNRT+qLiRZKXFLDLE9tdalxHt1jc
VaH22EGG4Js4j9R8/mj+eGdXhHSsjnjxV+q0XW24pHrFfAuF3iPeaIqdkC/eHf+jh7Qgn1Xpr+TK
ez1wd7vaedJcej9/I7D3iwZ5eeAWEmkRSO2IhR+noOdGgMK6l0bsSm6v8aLNduugohG+GwkNOZUz
uqdtsri/qaRd5hV20zKb3mcUJKrXbInD0zMw7TwjpKbAdKSZcp3hX8rcXsr8i4wUJyPVb3KKfE2R
3uy6SJGkE3ib8O7ITr75VWlXlwui/O4gscKweBhRWjHJNTdDJG5xYkVfP9hqZsh5fnf98UA6U5Dc
33iY2D5O6dzJsXAILf6PIYTDcvGCJJdKFur0v3m22QOOFhpKMyb0j4ewQLhBMEIqOYL12TxuhA/Q
lD5Qmp3Zki3MKNTOwKpqCyiu0qIR8DhPZ//KhHWnySDO0xeoA14HDiXj3DHYwHm3nkFsNwZ6CYb0
sLZAFiVNZhPBwwdSwWo52hUA7npVub4BP+nsnsV3VJKvxtGfaw55Fy27SWqPPPTERPPh4rhaOibY
W+YM20DKA/FaVeDxSD0WRKOaqxjgQYF0G1plNAhOmykMv5I3LoCLMa4ridSeAHyJOzsZ6He0dlCD
laXlAY+27McMHkwR9bvgK8bHI868Wzl9Q8yNVHR1JMYVuZbIbgVbhd042j8tFjlI8YYIHBUEsGeT
hexcJaaKX/ucQcIkz3mxTObozlkxRFgJJlN5Ho2phkIf08UU+SO8JKZNGIuXLb4UCD53HpaUapxz
EvZq2ub1MgOrNQmJzO9DdMuwehFn317D44/MZ1+9JeA6l77BTPM2ZewQTDNiCRdQa9pnjdZS2Q8k
V8im4LxyS4eaW4BrF06fYlNzXSZZal1hGCtRX42gmH+IXWjXePYqvUJXyDCVE3OOtc4LTuxYpCpy
9WAUcN0CeTuY6zLm21CnC3qC4PSlhras2UxDUw0DpSDwQIAGqldrNF/PmcsQ+RsdodlF5sxv0JxR
7X8qfp4maY/KBYWpqgsv6BrF9xtJ7GIeDmN4WhakDKh9FprsAL45kIr0nf5v45DBzQRkrVYoYCi6
HjipmVfFahxhPgSNNJaTjdIb1DS5i769YK9skkDDsP5EHkyhsPwHE2bDdQpYs2o5PIapB20nk6JW
NPNSIl0+Co5IZKB38xYS5fALuQ+sWsfWl3Jwg7383n/14xeXD/bn5gzavxi9qQqFcgwaCHec3PAE
kM7ZZbsC9UXW+fsiI3WQ7YcqQaijfu4NQo+Vjo5RsfOxTrVmPz8p1rZ6A3Ta20uKbywzXd2Qu/6U
Xkl4TBVZSIFcNlopBWbMb5aHoA4u3R0O2hvJM/EoJnl8yL5oqupu4a7HN6VdZjVY3/+dS2V2ACXx
B85T7mV2OC8EVlUosKoEw0oJVxxNURUUV2ZzpiE50ccnaOXcncCqw9Pht5c97BpJBpIIcY+JJxFr
Q45cQNWsUlZE31qacsaGLmjb7UD1wPzABHBSAllGLPpK87IeL08npMuQgBnSvbIbskq9pahqUIU8
MV2b2B7Ee/qXbVGgZJUtMgLrudd7wnhJjNZ8dDirM9dsfZAE+pZgxYJwfIYLtH4W5MWMNexzjqMv
mRP4U29OEMmtTtAMNCqvxxhjmsJ0BzdjUNFsE9qhc4PtitOlszceKGHc2wJa6G5NcXKRs2h8ASrz
SyK/sWSrx/fOFgoOS32ZSkF5XYgtunvpU2K7ZpuYlpKo+lV8Refn24V273J5CTErNfKi4dRI8f+t
mHfvEHohO7611x9gtBsK6YVdOXFthHKLoJUw7fA43cHhxq+kOQCHGUKtDWLhJPuq1dbbQ23mCWJf
CIA6hhMEsmlXQ0zEeSc3KnthGdR5ktLXkOmep/xu+jWC0YTjfKDG11DdizfdioMAx+zxjJPkhVBP
iwIaWEmAyPXTgngOYzSlubczwir7yj89jzBf5OeK1E3K+LoYbwTD6NaXOD77ablzpusb9otc9AqB
zFPgJZgueZViMc9LnSHgy5827NUoRo9xZPtzAMotMW9l0KQdTivbKZF4yABZnyhbSDeMaGk6djZ6
fdnKVvcwQjiSNpul1kD+cAPkJ7mSt5beRifTiIG5IcIblRTVgVJJCzB8wS0vEiYXUrwXPOOyXdCi
tKKjcuegZiB8LAHNkDPap7v7LIoEe9mljcRdaYJV8Y3lo9hdi+km8F4azIEzo+jKVc6SvP42kNeu
R7yJONrX0hYQh4mKR9lZb11WA5SxZlaEfLSb/S37U66m6YK8DM3JbF7FWaZTKagqOR7b/pvAxBba
nO4hB0GuZzD3A7ilIBlSstDBh08Ey7XR6mDcsoHGAANmD4BTOPPo2l7gecBWrTG/TW5YEWNr91NR
LE4pRBE/73xnge1+rHsp0FX4J0P8Yro+KdmrDAdIuPwX3VtCGlcWVTZ9afFG6Wa+IcQTAZ8ewL+P
0tg7CPJNuOsE0TBZiLwd0e2c3i6Lt+cWjf110GGPdGkYK5CQOKk841EWq4EAOy7JzwdExxArF95H
hITb4naDxBSB4A91hkjwaXse7PfSrgr9NxVb7xQ+I0kSlQR6RZ8YUOyB/XzGEWTB+QTuf78bHuZC
UzIzzPSYNxZI2b/be/N7BMkPlejj4NGxEPbKqZgKBEK90tDVv6VUueZft2okOr+nLG0ExaE/7C95
L0g/zDOhkaEc6k6DP+i90jFaEqFSfNXp6ZCMDhgTU/kkmCAYxC9xyzYvpV0Oyex3N+5Y9cZYIw0O
3rco2abn8VSvTAtI6XsnfmOxPdjQS6f3C1tQrD+eA9tTJm919bk0YgVo0Q49KYEEn4tfeoB0f4+/
OqyScmtrYke0v7hpTD2A2keLyN/ixE08A8d3MVm171wPF5o2mgT1u4ewZ37xrYDB8+Cuh52NdB+J
e9yetsyQnTV5sKwtGwuBTb4FZEQysQDwojGR8nH3DDYqic+EQvm98eXvv8D2iHf7V7p3Y+qjCjbZ
SvBCdNAQEt9NY6VoEEQiwH0U2JkdKQeSqU/8+kTfVcDReBOk6mz0GtdvpCy9Hq8oGllSH3IRx+Wc
P39R8KTZsQSdp9d7GDQBq8REMMXfcJEhOAT4DkV4oaidHNjD7PERXDvpMVEitgo6t7ojkC+zPqMV
/VuoczW1YCITTYPjsAkd8AQZiUisPFUnmfPt3HHdVzMt2VQ/dLtGqnWzQbD1JzLGLP1yDz8MJklF
8XUfTqlJx0Dazrzyk58wfBQGRrHy/9AlEjh6y6EJBQIJpE5T1F/64FqI0TaCWP9Sm4ihzYFK+8Lt
b7/nwAHeyxjF/v/l5jxcped63zN1LzM3uZ1/0RFyWLTk8csmYSUcDreSyjYoe8WaDOOd6B8HZsmq
oxKXuVIbXmDb5WSP6UkTd7I9egOFbkT5tADb99uvAilbBWPiogE9rLnw2OaBtmkB7KiKIzKVtYrq
XvVYQtGnsqBVrgocDeiLdtfV6nj2KB/3haN0UQruluNASu/gfg0w6LvXrsttTq1FRX/2WW7TPb9b
DcF2y1dARXc9INbjYPl097muorlll/OR3ev6UoRCeEZ20nQRodxqBMXCMFHubWdus5efRk0nN/ni
p2sE7Nu6lS4kIgzhdS6gRle9OJql51sMNwYbYLpxS1+ievFW3RJL+ihF9S51fMpPvw3ZqA1ITr1U
dWWk2rDEccAWdPYdDJIWFlou9aIuZ8GQuPLQ8xMUADhaKORIwnDkLW5QKkcwLm2D9mOUNPD+BnHA
c0vKZVRf8WEqle+6uLfnr5Joff/oVhCCF064YZz7A39mLLS97PLePHFikQcqXEZ5pcMOPyD8buTA
tSZttGjNHZs+ClEoK+ummw0zl0DJsdaI0a9RUiM5Urf/MgG2Qb2CJbIJCQPB8mFH9GjjT6XgrUkl
VPijDAgiWDJBWgTwISxmDkFWC47bT8WzCtnyWgJeBl6fFHWTMerzMlpgGt8llibYEA7WGDxaW5Zz
wDD24TehIXDtBVnNvapa/mK4GRw44d6tCLpR6kkNvkySLL0/Yryx/dAdowNBILaw24WhosddTQNb
vJLeMtSDxCPH2rHb3uWDwujcOSZtKBTJr2FxQhkMtAu109cq9eh+e+odQogl1DcBGHpr/SD+OCdq
dP8vShLm1r/kxCcJ6Gr9zlTLg169Ly1BAdN6lEWwHDlro+GuCkkGByYbglBoc7bex1uX6EEpGScH
ciL7yIoh8XGbnWyNOQUwbSTlIfdEgs+zS4Wej4ZCz4kpqk1EyluBK3TNW7uMF7d95q+RA/7l2RkX
yDSSkzNze2lI/gcA8t0cYuvdDKn1xbnVBirGDYBKJnUfALM46V5jONUIBqK3HOA7gqx3XGryDPXk
xyrliQGbMPNFdJe44PoOT3jRWc0qZjRtPp1G9q1qTFX9p3DvbMbFElY0UD1pSbV5AOmhyeu1FUTx
lBgOm3qjidkQBfyPxaB4tkURbxcL4FuABWKvJVoXx95u0Xx31c4T+j3PnafpfGKZuiG67WmkM9ht
qqslGaXbxN9fsmzQ6cSIlqGMSBJ8C/8civJb9MLm3taaQ66gNYHXGdwT7KXp1Z3Ir1fmqOpw1FRX
2ap9Lbi4k86AGi1jbiP9MKc5JlGY77v2T2G4hSXki+q3eyxwX6+wIGiHS31N24G/Le0lcVMdGy8/
goqIoYOJzUhmsDkolrtl0yD6YXureybDRyilJzTyUW9LSxWjCvNcgyPGgY0ziRufELJuMaP7bxFU
MBSRxLgZnnuU7R3RlrbIbu0FV4D1ViLB0SwmqNA6vIGGtDHo22ucJWGZu5dnyfV1U0NG681TqdtR
fl0Ik5YA8+cOOIIU8MyplkJfggg/kO067GRI3uqEwV29pVKcL/Near7KvEgqA2OwIP+X0bJ6gZHw
Hf/CdC1D7V8yENj0Srar1rXuXqLE6onvBN9+x0/PwOX8Fr8IrDcTe77gwZdkaArw3qPBXAT3Ok2L
CMCRQFfCopca0kUkAaoAnGEpW3lWPNrNUQnjTwICHjOi33Ike8+A9bbvbPh2G8P6+YvMzsKHBnHh
fqznSX71IK3R5hftZ/qMrEOHTmQxEsnMZaE/Tf8t6OwyT1PtO1r1h4wxYmQ7votuIir5Oi2Y2gFN
WHA0lo5NDCAMMBxn6aUeztUoKXI0QqRRJL6as5bNm3BP69blZktS0rvRptSluSeMsuS96qLj6w2a
IE0i5rrC1dk+uw6hs3voT3WWF26diAAPjoO2+bcdOZygHtvo6SzHaSjlRnaPSPdhtUnAwMlh091M
Np2llz9pvfw+rY1pBpgfyhyWRyMjpbtYwKuvsYIJVbWSRqSwAU+C2NG3oW9OfNr2EolmnAgRNDdW
NTDRqt8n0v+R0E6O0VLcV+4xSba1m6N4BwmpndK7FG5aiBj+9UrKegj8wmrKiR5x5uCNaQZjI2ZR
JNXKlpt1R42kQUPvXxnYsSXl8T2O91MXY8qdiMlklgJuCVePgAEBIPIEKGSmlfqGAhSlfcB6WWJD
Kif1FHcuWjg5Ws+rc/JNf/k6D0hSNfWvyVwmWvwro1dAIWrUlVmSJG9fkLdXlizy5y2dcdVVePXU
+CBgGZHMYpFEtq9EjtYjSTPHThjT5a/23H+RU4HS/IreFeY9ah1x3cI0APWvmaXBa4dyyMtPrQAI
9MGtEZsJ7Er5Dpwsa7CF4z9+jyY9CkHNYQTZ/JdQ3UNL73aHs6EqMHIfR4HW7Jo+bg17XnbS7WCi
Dd6Mfm/UKypN+wvyQeXEINZD3zRZmhYH2NupSfr5n8TqHJBxoX8Cf0BH6+CXgRW5ENcsLMW1MgXC
6VyozKwR2LAZC0wbm8AeVKHdxsiPlS0ndLwZKZPGyiggCXCtqmz2A0S8WZVKmaVW+QCOW672sfOy
y0jSETmUPWM4a5nQHfTKsHFgK5At4hSGY68o4Ur5B0Sf3Op0t663o5A21wE1uIPBmQgw7NEbTg5u
VJCyXG4ijUpCM8m+j+L0m1u1h+kbI1F6GGAbx06SIFivfAl4+wa3bpe9hBkFD1Fgy3tEwmGGyaOv
2c2zKGCcRqB6nfnkriDpHShz8c06NSF6QGq5H2pi+c6nU2WnJxZMu8iG1yRR1UKefFi8PbtQI3qO
wF91Nbo8HEV/VvGkVvAFo5KrGEZ9zoyquQrs1rbJNvIac1WZSYaLOVEROubaxpH+6VVuo3OQgGcv
9rX4SmFodBnJ2Qnc0E2pW+Qul15eFUnyIIlxLmLWwXY3RKz5R0m+x722TwqhflaZfPqu7Yi+fGVE
/5Wjg6BL+dVzsGBr5YSQ2weEeh1Wvlep1rlFFhAJYj9FXULxNZy8Vit5Z0hz2gUagdUgmnsqJNaA
VQtJ4/5HsCbcJlvn2a8qRk6AR78z/Pr2onk9G3M1WGah8P/r9nFLyCSgE0QsIgfbLd7vJzpooC0Y
gp+cMSsruh6QapkpIfajw6jCQmo25haQEQzzgs1ShhQo1vgb5k45dRASTdMhwXXSlVUSq9Kkiec5
hrXUyaO+3BAuaUlSQUd5mBKzj1JKpqklm/9e2/StJUxuVhyEJ9GvvG326WQ54W4bhpZXCQjL+H+u
nLfftVQ/9ieQx7nUIjiyNg+FAwliYV0XYmbmooPl8Bj9WEIO7fQo/pLSsOHDa0PalGhxviex1kCI
yb1Pkua6bpaeG3zHORHrOBr0Unk+uJAVLjGrpjA5OrbmitAJKdd/yMFWH8lGXNkaZqy6Kku28/7G
nGNRCeg9T5k6z1JiRdEAWMzPuTrz8OMZie5oKviL6M8LaZunENw5bwozzfNk4ccuydv+TbE880TL
RcCiEKmEylvVptY0BpYKaA23RnCUxbxoGe8x1GbNSO0OFnwZUHlknCiPwQI/xteoVshrVpnJktoX
w9zBOUGJJuacsXjEN2I1xPVSMHZwvJXb9BE+bUm43kEEmn8omaQySxMsBkv2Y4Rd3iwi7FxQkyby
22QkfW4KS/Hh7//+ENFZ3EXJKny7VMe06JY7e2kfsa81vr3hGGNSLZk8SS74XNwwCZwTbxTfGWAX
gGr5c8vyRbsIL05LmWPwPxLiJG7pj7L9BThO1ZEG0MV/YNvcEPk7dO0HNUBYwyHKNO5MNMGIzOys
5p6jkrhP2CMYYVL34dbh6LIjsgif9agVw9wRUfF/p324TGy0cgAAxJcoZiNqMZQJIsEzXLS4OADQ
uvIol+uGXzCVVZ+HvDulNeI5xJM1mZxlqkWtv3aDwk6JWO0v1XTcP6b/TmnPGI8Ysn8Wrf9DiEDA
HCsg6nnz9VCIJkJSrkZkw+eM7t+73fw4X4LGEdmv+vSVTjt5jbXBbVDD9g/ycoKbevlhUYwE+XRJ
kEVhQfidlq9cO1erzCeSH5EAq5wIsodWMeQHrTA+bAVZc0bxLAXWpE+Fwib77srVYWd03GPFT2T3
3Bsg0LzAaacBWiYc0ypWcZyFiAPfFI6PkGPfVEF7UKnv40T1cv3GGhlOGECo1D7rUzrnRy27BaIp
xM0ZafSQK3B/2RsU4GyDS6iEMh7aStl+Mn9iAZJiNwaK9BYA2GbCbfQuaNJgx6gxBwDC7VoROYyn
3AFo1zJCw05ERxr+Pa+LhuKes9VprVeQYobGr2LAJQFUei+8jAjwTXaOEsHIYcL/l+RtKEJtOMYf
6kIB8TsQnqx02y+MPqsaRgML3mQvUxEzcBxGEfba25fuzMu/Cmk67lD2se1tMQUsyyakqwldK/W+
YlYcpH4jiUx/YMkQqldg4O+bvyhYEZVhBLNPksmtc1tnBnS/qrKXgkeY295n9Ua3nl8CTYlGdJgn
A6Yl6Uj0spf1y8WrylAwZN1V+LlXCo308WW+PSg8E6Q5jRKBrQEBl4sILOp6aTeJHEiGVQGzZcC3
fzME5Puckjq1vI22r3+sZqGq7WLW4LuNuy/i2m5dMHq5tNrDz3Ub87jGUgtNxUyorgooeDZ6uL5N
INSizmCazpsR2SkS1hByZumGW2te2BkVz/Ykz22AZ1/jkOcJMEne+M+4357FdMi9N24fPGAsGqUy
OanD5SSkPohoLdpPSWBL26bMFP6bFtkSL7XqGCaUdUz2Mq3IZHtV6WVonuRyZ5iuoa9kjLyz6Jhx
rwzwQ3qZLYzoyUAE5uWexp9+A5mUCXEgbyfTwTeO77ccb4tdIQgZJkRQI9bDIo5nisgeig7fFb4e
Snm9Ed0S/HOmw3VBWzFrXEeHEkRH+XT6w3KwHCaKqJNV/g9ZDwtAwoZV8QKpW8ztO2fl0UUv+qFg
3K9PZ6VXYki5+Ob/6F1fePmn7MryvyhxM9Xx99JdgFgoaIcytKiG8Dy19ReXiJFwE6WIt511XDJD
iC0msAYiDaMoce4AjsOSRmi0fZGl3eILMFbfYgQ4KLnsLpGkrUCAJ1Polnrg9KfqtoIOnEFdcTJp
dZfo4HF45Q8FTQ2RGzfo8E7APk+O8EsQhbXMFuVpbPWilEruoOK3yJxhs4htYet7JPrfRJemGgc2
vAxGulSDuhkBVrGh48wvuo65SbiZirFVCNtBxo7Likd7DzbzQ2M77YFGWP1Hljr2gfhZxVjgkFzM
DTiECHeTh/78F6/8k6uhs4uK6YIZ/plBe84h8q2qFT/Nz3TgKI2CxCMu4RwoUhVfidzX1WcZjCsu
x2cEFcWA5fkVoEGpN8QBM1BzyBsW6wByvzC3p62xLKNb0+U9BdxzTlXfrl24dsKQQ1JKrbslx1Fi
A88bo3wOW/aKMfIL6lPXCw3HsL06aRhLM+ty71AZbQ8M3hRMnNFjSZPsVhwwjuz5w8xOMbmdn0Py
1XSYi/EvHLMDPm2ibtavig2TbaxuXDL3/xG8L9qeRBeoeGT4kBxK0te7Q7M0+f2Wf3Mag9OEiE8j
inXz1icvMQYmDVaTSev3LhLMF7cQD7wle60h6MME828m+1E/nIC18wQ/2zaaIZxqdwTyQsO/REJT
bUMmMT0GYKecd0mcPyvhcCRK5fiEHDwQ4YJ9QP9P0E/ZnGvy236LJxdCI60jonQtnrKXz5rAk+3p
D45u/9Khwmvh1Spmx/emXLIVYh5dV8K4nwXc5Ag1xOBIdpLjTp8HDOP8Znowfz/aQCy1yLOcerr9
UBOQ5SzK3QNtBUjfzSzEqN4pKo5nwNDRHe+8ngxXOBlNnDtrjl5wuK6/yLJ+K/kN8Py4P1DmPxJs
xypq3EeqIZXTaIOStdvUpX9UeGS00JgZCFb9u6n2AfA6NE01Dt2CpTY+6jex6DWlFOkBOFzBkR06
9anORem9Vo5cQoFgY4AoL5cpu1OK8/d1JAY1ZuvuOGtu5/OMiA7a1T75Md6lv+GMetv8KtXNh6MF
PEGX0dPEqxoKyPXcl8X6fk9EAwdTt14RYlsMw8KIbNKeMcI1hd3xsHDKO4k86COKtwb7v/y7nqaQ
RH6v1G91TScfFvTGU5zMlq2HlcyRdU+PTKau87CpZWIc4ottpBZlDZfkJRcjzoPqZNWiabdddxGq
5pVo9Uk8G7yFvDu1Gkrbm/Bge5o/ZjivoKy9cNclymgWuonTI2l37V/902+qnx8PZzpqAq3E9lQn
E/LWPIVeE5cBLN8WYLNZehgsJwK+pjohP4ZftfEMM4uRcW2njd+0HJ1Do+ujwrLB671wsCd0s+KI
O8QlwRHRxpa1jNSlgR3hCsQdRqAeuo7tqcp+7TQq61gC86nDHchPA2Yr9OOT+0H0+to0Va/07ozq
OjJvFkXHHSZmZN7bRh8skuDROEgYZMjKbI0TsEyde8Fg4fYh94TM7T3fYPFg3A2uaVmJhBxWjKzR
pXFOWD6rqniiOXjS/XPuypaKVvP9066Ld/MTQOqSz/mEBNexNnUpuHbRoAxcTSucUkXIG86YkhHI
ztkUSt3LLcwJrENqvTNwvJmC0XQIG5fncFGs7mguIHpYe93PjS/gSAmizKTe/kzP3su9TEEnxk4A
yyCNzS2QdWgn0i5JKDy9O/c7y++ToHYOxqqq6IeJnJjkVnYbjvykBqBaznESQYjchHyNgbTfcUOy
uTq30CHQhY+77LjNy3Muz5aRFcV7VBrr1fpmBIceuqdBE3LAxUkl55ORIdjWYEpMowAZHqUzm++g
lFhiqKq9EPY/YxCXwysts0NBNjLrXT2/tWadYZCBeNAN01h4cdeAdmOctJaADzTn/5hLEwSk+luW
ruM9r1IhR9zmk+XOcXJHTCjnNLMsTTTeP43ibho/PHmZY+OQ8o0FcbutkmZj92Qnddh2kZDruyyt
N/+ULc5VKCxSCVJqAryevP0ka88u0Lbibvu8VGszwUXcWbENUg9S0g/pQa65yBVKYqrL8pF6T6xu
JKv1pZmr7+bf+sGOdKc5oD/UyIpmIkugQNkvXCGU4f66xkjdvPAWJIvh4Tgb3EPMS19y5b3PMv5T
1jjHnYtiJ+lHBcD1pcY680J+FNktXP7lo718BECkrYmcIHb00pmXDfClRqQA8UWIsCi9RSwQmoT+
RTHIQlNds9oBGHY4Bmf6SrFZNUdF1RdxahbY8A1BxOyJrQm2AjoZ8f9BhMe5ykfrKKw9UERlDWbm
TSWQ12dJBF5dxrbdihBR99kp/y+cW7MXNbl4UdQTSr9OBoaf4Tc3ckEXHinGOW/nj9pQg/bJtWIC
EWm6740n8WeABPf57yQwnVZ90OHSOsCcnzBNvO0WkITWNqiueUlKhyZx4P1A/tsd1jbcD8nDb1d2
wJoJEHgBbEAQQ7Fa36R86MXMYZFhCtk/0gBmaxJ+0kqZa8ErBbzEq4svq9u7WxpoIJMmpwqcSAwO
KymrRWS0pnytj3+2NjOBD2up0YxiMlXyxFU4a+nAl0uaFvzMMysj6ZbI01AUjEXZUxXC3ZYIMJcP
a7DDHXgrVyaRs2omYy3Eh7lkDvuicIhItT3v9jnZoZ0Sal+xCPacICs8GGx0jOHrITtNmNB8A+mB
/32pxjaOCJOZczMOrAGXKh+KcPoWxl8y03xKhDhBuezRwVyE/kQDWNbgEfjjoFCzqFhmd0bK1n/k
N6W+OOj0JpmXV67pPL1+7fNO1z2BH6TDJauHjs8H5d18PEqRluEqUtGgA/g9Ps3vrr3bbyuMflf2
OqVMsiHw3MCM3gZxQd2gjhSsVWyClDVqCCBAF19ThM/3aZYr+wDYBar8YCsq8O2KCV4mzoKpDyUZ
gxNnZudabqrfJViWNPl5VU+Fjy/AIAmX8B2uV/5c32k73f31lNbOYqKboVKK30VjUEEML9KPIZbt
QoTFs+0D0fttC0rNnYEh7Q9TA3QiwOutAkoom1h+S3Lkl5T2na9zAfyVLHKHYBXoE1qakjzXNbow
zi+d3aUxMYRJ/Nt3O75wN1wuguaH2sTNZR7g9qE5MfDCBl69f+Zr23UBvqKcvvojvivWermVx0AJ
4vsM6w78KAyRdJtK5QAjis3AYs3cnB4UonQ7UsKBrSGc19wqOzkBdgxm6MVwKneT4zMfn5BUir8/
gxqkljVroBrq0UPDpuMIgNLiaGo6AW/lzenaWoJpELbkBkejzAa9IEzNQVVh45t8AUXpA/JddEvO
xCJDSjEp9x9/qLzgriBZWNfPX9FXwzTh8Y9sws+LgGatHXD9e4GxmjS/zUFNpARL379FdQzem8RV
+m20TEQeprVOXuETOoA2PCtyMzPSr753MnechP37Lxp+hzOz+3oxDe8v5YpXTROrgaDRR0fJoKYN
cy3myRR6vpXVDK10aLWXJBikW2OK+/nnpDxh0Ot7EL0cJmxqTHlSwnUTqjgZOvCylzPUw8ddUgkZ
kXUZlOCLI8gFKt4Sfdjc5uXfdftT5Nyq5CGncOT//ydtouLgT+9UsuQHPrf5GUv33OL5laexEtOK
PPboHze87rdrbrZ6fKwYs41iBGduUpapnllBXsntrJWonwZxhbgx089kRhnbCtcnrlZTFadi0nWn
YpvN62yQEbQaJmeuzWsWaXgLQzzYr41DU1Pw+78wtBxH85S6TZalGF2GNKltxOnhBKukaP/CLF1f
0LGR3nkcIbctxuBXXdXTLNNbL55kpMkqAeK5SuLoW3z9sDop1hmpJKjsrShYJ9h+XbzZjZQZ/UL5
ygHkxLtEdddFqmZjjB/zd/V7mGKlVxMBcNN5xdei66Wx6U6155hAvFz/i71dME0TLUWt9igTIDk3
wYWn3mL0cuW3goSeWuCG4ltiLX/+3fH7X/YEErdqOPjf7bqmmufwAGlZu0WHSpyBkkzaLxKCiaIL
l9LXtz9LqBsOt8VCblz7ogRQX2K8/1QwZakB1h31XUObhfyjf75/eFASWAkjMEYrkzwhopm0+qAM
sDn5pZ5SKVTjposD7yqjo4MoRekY9jXKqa2XSByE/o9pcMxyO91v9tkCDmUSKiI9YbRLQsh+3b69
6bN4Ze0o3g5FgEgaKS1Bgp0ozsqjcm7QwwYqKc9MNFG09HroLUNUjuTeoxjeuzc/Gjy9+LbhJ5k6
e9SRXLQYdkOFw+UoWY3pF8ht9kiu4A/fOHwxjJc3AAWMJ4MXK+ZHXlo/DH2PO8ZWMclAfZjDoqIH
2asBmacieufkxZRLq3lEfm69XUEbOAhLcePSIrL40EGJ36VNU4z+uw5CobY8PEqMcZdVJiCNz0XL
oEB5KA7E5Z9tfkAYQ2w5+c+p0sgyOUD2B4ssBqaWcVYkGoK+R6kA+Ao4EIZQz6KN9NA+9L9lp35v
yaE4c8U8ltpykuHAGXxpl08nr089D/nkVYfr8tf/87SOYFghzGB7EAA0KavlzIoL7wuNERusnj2e
KLhqXO35reYmdCHh9o9aMHi2XZctesS+hwaFffmzcXsu9ec0SFinXwFeWqH2sPH/991D5LKQ18Vz
hOf+NfOliuc0AuAuhQajw9BBa3tHfH3E3s0uhJbYYnVMnS5tfU8mdmBqPf6WBfRRx2f1Z06Thp0O
kLC6lALKbtaorwSel9Cy2eiH9sy2WH1QgpynWnNSpYKbOGPgJ9sQOX79BzqFJ8lUg3gGRaWGOcxP
+xRgXS2SrjfLFSTKOjwOUFERTTiBe6rcI8tBDPrc4YnZxXdHsNig+svaeABOvn/3ZdG9gG52NNv9
kxDKCv6FexcoBYTrAw9lp8EdNcZMP1FPkFKjwuyG693X5fgAg5PoYpfIxq9vucu3t+Ap2C+f+vHf
vaSeVCMNbk86ElwYZYXIVg+GrlpnrxytSpHdxcW0GE52uhf7L2g4xN4FXK4P2WBJ9BcjyQ/6dqnj
ZQzZ2uQgHSm4xMzHnB3wRucxUlaCV7owjfXL5Aj5DduXP3Zdj09MiJwHIByKfrwVLKTLIVFT8xUW
FcgSotEwDtotYrKmwbQZW3nVyF7BSvxOEI45B2Wdy4uFE5uoWVilMkp7y2f2RBwFhLr4NTdjggtH
Wy9yNpxDJDda6xFw3Mk/GvSi5D3B87tppiVGglEz+gr9MFGv2r47lsBt2k6kZqznhqGlXah97YCs
t08iIxpUxDvGf8JFsZ3LmtnQl7bD/wRTBsV8uR6SSekCxHXbddXJg8lYRYxBBvpcJE2rT0OihUT1
R7wk0XoIjkkSNCDRAt2M90BQz4JulJximNdSzqyyZA42HYG94avpYNiCij9PEWqlMpH+vdTPdpQp
iCCVqYFTL7D45EREOxfv1bkxD7wPJTUJu4IMrBgn2p/JnuhzirTYY8pFI7lLF1Ta5PLZrPNbkswG
1xg4NrSNo822lKA0W8d/oJ1v16SC74PFfgAUJsiUJiyqnv52itH9nPH7vm7yTrGIawEn2fpkx/v8
fUoaDEONtIPtwtNEdoeyJDs0QfcRx88P+a0xi2JXvmKhKTwIa8NZ4dUtVryS5vydBawm8lbTscUc
zBenMcQJ5hTMEpZ1gLpNU/YHaj2uqAqbY4kXkwWsTAH9XBmrOxHN1AJKpq/LaOBowKksBoo3YrWk
KD6C+wRdol0Ume6h7sm6AUkVhBtSGBZmafzOMoqk2Fo//t9o32MnmM27kFyddcXkv9p4UUvCNE9j
N3/xedPi2Se+z7aCupFL5BwrSks0WOKgvUbAbe1u6LE3aoS4j8xysOeRe7YxC/XOflBrOT/qeU+6
+x/1YMz0vcaJsDXRqKf3Gbc/2rO2nnwZb199VZHsw8b8E99tZEcTBsDZqNIeq2z5SXQW28tub8YG
fqjFnYJLfDjPPKtEnRqOs8XMWdIV0Y0R+NlLU2MHCHMXwOyTy4wZLdgbc3cWdXD+mv6W3U2F+T3O
mvDFyk9b8uDLNyjDAMpvsyZB6V5ZIfABN4WD9hCPvE1NVYNozy+JfwIF2zm/RMUve2PUmhNjswrz
fS8Tf88SV3DO7Sss5U7u+CAojDeKpQJAUeEO1sYBSzg1TIYEGxlME+iaPrGuKDU9CtfjYCIH0Ztf
GXKUMQptYYLPDGO7cQE9aSYth7rUYw9+8xGApywhZSB8lfqmTt0ts+va2j9yh/HfagnkHaFMU0Ni
YO9eArhgX5g/SdGDRQDqSK/Y149ilxkbDhKs1ZtrFs8meDKo4aGIQlzGO/HtmXNPajh5D8dKtB9w
H4ZeITAvZADSaJZyp7iLH9WUNksoM8/1tCsPqMcAFdQo18ggR8EFqydqgPyW+dZqEGBBoFFBRdyW
F0wIRESRXJFPuMppO/tcRayRz4W3bDHCeTf7ibS7X1qoWmaTY9zKJE5eHz6INo+/pzlDNQdrIZEC
072buyire1Ls3sjhA/ks605D2Ph+I7N9hGi3UBiP4jSNllsN/BlLpQlpfDQCLmEA0umitbR+he7p
zpfObG/0Qf9CdfOvhxv0w+ZgGVBYyNqoFTztv58fdyu45kDw+bCjo707uLJlB377QID2PPfoNlud
YcJDScECTpC+xyC/La1t7TpbHdkHJcJsijZtj+NopglBSa01srG/2IBgO7ks7KO82glvUiehg7Ql
veVUArNJbyZwn1z6uZ1R2PLhGpb798do7LJRS6xBXEYlWIjIi+HJmQvv4YVpnxJDVfm5qUk3rvo7
hs5B+0ahMJTvvBcQjKik3vUpqDMMxImkOVhHR3safpSg5h9rLzJyBGtId4Zz3TWj+dgi4dIVIo5I
bJuWCQ8Q1sMpJwPC63i3Yrz3eX3wwgnQu5ys+Sxe6Rq7zJBqEnir3f71MPuVPmFlyZoaub5q7Aps
LRsNPDvfbtTf6oSRfGrPGmT0tRP20kb20fKh5JEmUdDEL1gkLQJ5SfvJDpMM5v+NEgQSX8zSmCFo
xCyztgZc2XwDxKeezgLaRea4+TDX7Zr1zCx020IuVtmI3srcxbJW8+MRduqIsXXkbpfW2SPTYlSs
kUuXtqangtNTLCPeKKR3E2QWfIPD7X0ju8ooNF0qiBvqEnDvZQ67BCUBRzraXOITq578F6xGrmg1
tb19c/QcBo7rih8Q+m15Xn7uHZXX3i8iilv9zJd9BwxR5fQivRwQdjufaeqN5RiBQ2zWtRBRwtJy
s6JJy8Znc786s4nKRzOTLlkMUmpH4XGpU2V9tyHx6TXOQV0JglemMqizc39uBHd3j55gJg75GVwu
gG0KiP2EEW/egVM12652ap5uNZyf1+llz/MDKqoG/yqpCi+QbQULELDRwxH7nm3BsWjgaX4trh92
0Fi/LOSXcHx8rgr+diNWa00BobDANNmZXTHDd8/Ls7Cc1CVUuD95dDnEY7y56clcwDzgtzS5pTRM
oNovNIplQ2W30yEt0bqbukBIsQr8my+zcmewPraIbqIu1/qhe4BxwBD4ZOCqwATaXtyFoln8lB8/
fgB9pK4xkepy1LqEeI/y000Kph9p1bT33oORL27kW5NKvhQhNsNVK7pe6lw/Ue9mJyMfahfLjKM3
3kuLQsYVZs2iKC8C0O9z4yb+CrcWnfsaKpqIQsknhXy2MxwenBrMm5GX9i6Aw2xKTdddE08kd8MF
UN7lxcWTnfW5MgaD7tDbnyJCL6HZAIqxcqlw2PU7RNQJy+cg8PVTOPvOOKSF1zOeN1tSvNMY/S3+
VXHLBTWerYkzDJ8but4boF/kYYsNvNA+TmjZQDRCHKMoZe01m2xoYkFj7SWOfv4+SeJLSz9oVBgt
pVNCEwjrzGqzwgN1kDuuZ0v2QdV0ehEXDHjaaq1ytNj9ZWl+6QqtLP4QHqFYjhsMboJKilLPPRjD
FWcFIkwswZ3Z0OsshJqRh6d6cm55u10oeQZxrzkKEtv/66XjA/8UtAPFspE+I6947zkfWLslDWJ0
IkZpdQWkwf2GspPEBLM1I/7YVaTmvxjf9pJxrU+wzTpyWm28uUc+pecVpcfQ6biLA1NmG1W0Khnj
Qio+LNczIi0uMVgqge/z40eNjoAu+AkrKIg1BlsiCIGxd2SGdmeFJ8N/HAPpWBSIYUIINHwCeq/s
2nZkzWYNiC+hnUZwp/isarOPJqNWqVzl2v97DAYQRA7BL9W8sNuFGt0EWyEAuTHYE5cHCvLxOH7z
GdvQmwfFSCEznADALxn+GCYSNhF3OLziuvf48aznEIzNDOar/UHJ/iEXYgVNjXL/xkY756qeTA7W
IPx82DHLtsOSUS99pJpAo0+lsYZvJK6eDGxlRAXU50UtO8fyM2/2JHXsKU48HgVZlWTMGTW9Nabo
AWUWT5iaNzm6GrZ9lC1FmXAUhVrd5968bp2Y6YtYeDULJAwGKWktVLw9GBxJi0WcT914yRonfuIe
79k6dg/zM9GPSNrgu2XQdK97uSN0Yce1Nkys00cFC5KT1XtUaMR8gtRIXfeZKSVpmoky8CrPl855
e0oDF64O2LBmWGf3fn7M3dhR0j7Lw71Xc5dZjXT9MyKIzrPjSTekY3sxzhT4/4DbZ7PdxaBhiNTI
Oob5yOCIStgpCfs6zmvfnUAo0Jdei4a2+Wh+sBlrEe7lzHBpxNSVUscjwOgda72V3AMAbqCtdZsb
2IzWub4cfMaHacykKdQZI+6MpIenH2embiiPxyWh8EUZAUGQXjqjDXj/glpkjARJ2yJC81Ob8Awu
adRXRN1vjRjD9q/Sdbn1egZj3uXKD37R/nqOxPCbhD57CI6s/IcuhQbY69BFQ3dYEuTVXD5ptRm2
d/ozM0cyc15iFkeV3ONDb7RRs7XQTfaW8jP6MIJoC/Rl46fStRXpvWxbR/ExXSTqP1iYf0uWGa04
KTPUzrUpZLI5CRnX2ZeZ4Oa180tYMevgxuqzVIt3x9NCOnPu/JykgWBJWkG2AqGSGSb+Ab9taPBl
vJkt5amdJbD1plizpWmSxILgY0sjAVlaCUoc8wSHdp0hnSFbPK45bLQZ27pd7ZoW5DaRg3TuAFX0
Mir9mN4qkIOlLlLg7UEWmh0oIIsuJ+yrc4Fjb2TYR2d4S88T/8aaD9vWUw6EWJrQE6Ohf15KJu5g
pS1X6wXVO/3pdVOV9pQlKQlO+yqEhp6Tz5eF8UsNxGkoTuyQ9rXa9i9ZDv37mLDqG5azqKRszpuG
ZyyW/iTwvcg2ZeOmg+qfzBYsXaBBVwlPCK5ALIdt9LCX0NUC1814Tms8JCyw6g3gB0JKV5iUPxZz
uD6bJyqkO4HBNsiOelmrH40TOUCU/xKWiZgGtpwcVFV+NU9ULTXr3iakvusx6GZjk7aPLuXWZxrh
wunORp6SCTC/wDYVSZozJrig0PMRaHWNlnBhu0b8rNd4AgL+kK5Ze7JdWoNndJKqARnzJkwZfPip
Xl/5Mda88vIrHud+5E+WqgJIuNPO8EYi37qBbbmGG6nutpFmjOontgPXZ8nxsqTct/7HAbq9kClM
GK2br22L225MXz9FbIGLcY8Lv7bUCtzN9jB/awDHqPhBSDw2Xin4ZmyduqJJIlye9DZFpR2tFYUj
fyDKMWVz0+dfQXI7fSPVHfXhXE75kp+Vo3fk+RmjAFt2Em1hhOPcf1/gmuDw1v0eZKa1rpezdZUw
FDkOdgyPaPxQJA6IjZfSyi0rcahmaJcadvb8IRVFCDWYBDIa1DBF/VDcFtynjyG2RgP7XgTYAZPN
3Vrso0pSkCG0179Fjs2rxtyGMt2IrSttPQN+4OTHOE1Il4aS86mk59LSolPqdCom/3z6yFRvBHyv
vzj1pXySMOjZNtlGioR5zncKOmIRWAm/2QqryyP8dKg4Zkrg3hqGg7Jdmz6FcTQKDM5QL2uTakK2
MMoPfNGs09IA9XaEKuv8emUGhDaqQCSBN4hBl8sJxbtSM0tBUr20aWScd8fyUCcGluqfIgFT2ohn
5Uy+SnA+7UBf3kF1v5i8ha+K0KPfqmckjLr1P0iKOQBXxZjlrmB3KuP53mrttSekf4o1BECjF7ws
mfufIQHEErUZJ9g+JSN6Qk+8x6bvozJIcaOZcOovJ5FSmQXf4ahrqeLjbU5E6C8d2UZTo2JsenoX
LCOOZijWYaCRAVhIf4yfxS72h6ZKKEVRqhV0c19BB7jd9tMQsTdJzJxm7tmax1u2RYDyOwGUAzkW
OWurFFZetVmBHcpm/eN1556aRnrPAedREqPNyAYDkUBVC9DYJgipmq0pXKb3/woYiB3iE5ipRyN0
ekfO9GE/rBWrwXZUSMyGl9aJXMZ2rmfqZJn/7wWMmvylbfhhStNFecOHXi/gf0FXyz/w36gezr6n
kdq8TNEVWpm1D6qhaeGFq2HqLdnnZhT2PNV/Rf8prM5nhVh7g+LqI1iQImJPTstz8eMU/3Sc+IkZ
PtSTRQoyMxLtKQ+akR0VnVlk/9WB7kn+QXTZa3MG/6q1OiZ4GQWKyiaw2UzkappZSi0Knho1h91U
tXLmE33TEAb645VcbYGCkEI7pcmlGFHisc2gnAVnzuIx+0wOYBYK3WRi4GPcnSxMzC0E6wdnaTb3
mozjKM6K45sOMhmEAgerPTeI1JKopUnJIR6E/NPc/AtJI/5YcNJwUkksh1gGUjVDFswE3EpHsTqV
oZG++yOAcpo6uDFcunj/zH8uauFU0ZWTD7LRZZK03TH1RseUPN3kbNegsec+X4riwkJ7BzpZrYiq
hYD7LTTLbEP9vfPKANaGoFjgzUUd3TrFfpUmof7MWj6i8RTyv5xsRJZTfgC8nMqB//YVuj64GFQR
r3UqYnSskGT+2a1WfZHrKegYdLGLLCEySGIeP+DI78YEP4quctA3AyMpTo8a5dQxxD59tHOBPg+U
Suv72awVTMYY0gdShMRg/JJmLUq9P8gkGSZPAgzPqnEZLnbwi3hyY+53wGb9N7XMp2IaAc7u/2Og
da0Oj3NSgfxY9KyJXWEoNXf7Hr4Y0KuBLtx37ReDLdRglzHrGw0MW7+yhmKmfHJHkUOHtfE/QeDy
MFC1D6JwjzA1eeUVEDCntBH+il11qUFimwHst2gNVu9VElPsf/Gt3WjAopzoFq+DhGJVlK+1gXPm
KlOIQhOg0nBL0u3iLhLCDEKrJTKw3fmxLJZ9kJqsNHNjg54S5TzS3WYizip88BfVlQIJXjm/dP+2
EYuQstHai0uyirrVxXZjO2cbduc7rOiWBazRyHq10e/NBxpj5yP4Gl4Qx2CXgrbSmfadP873THqt
pspgLdZJhBy7PNs2dTaDL6u+10Eg+Cp9biEGsAE1ztxhB8eIUiKBYGueBpYBWsJz6+G+t36x1O9I
UJ8L03QyT62leyXE3TUwF0gdkPFgHCK7tghN61eFwrZodBc5olwC8PkC5OXM85U7LFE0nwCmCq//
LF+FRt77eAblgIH2eIAYnmhGf2UJh1c5acq7NN8ZxRfPUetYIHQLsKvliXDub13t/4hVhXjsHA2f
5fNCoSj9vpL4iphFstBtOQQ7w1RtxcDuv++KV7mHnXyMwrjM0Gk7GUkC7X3YbFo/1SBZDczkHYCk
rRhaeozzwSiUO2kX6EVAsJgqTJVNFZ5Ca1qtwnuNoXCHOhNulXn/sH+lleo+r3j4w1V+gtS8HSrm
068WqRN6ioUkSXqvr1PMRdsoqlsYR5y1C8l7rQL08IAG+HNyD29No4GI+tCjBHEtOou/F/jn3YsQ
smsyKDPkuoYrz2mxAKI3vvQWhd23NDAin7K504J7O7+5QBTCIch6mZD2lvgiG4qK4VK9J+Ui7MFS
Tfl/HGiq0Eru/vCqhGAK+njNK7wMEXaL4ksv3N2uvnRpzvanQlBaTmZjrl+G0k2hQ+GE6exxtZHQ
4KdNlyYvMz0l/cFEiNGI2lv/7/CuzVK205cqegwmK684Ra9uMRCSMS6k/iR1PJg+8LrcdhmVW4sw
Dbz/cUFL21AtPwdmz25BO2yjt/sQbMWctsz8205yRI0oQotyJ3mMTC8fHPWNRpkBSeUunSQpHYxc
BJkuaNyDqAOl5T6sU9Exf/5P8o9w0VnMlwjOXLd9nfIQLHnXLR2CvwDGH7QTzWH2Fi8WbWRYvimQ
2qsrYrAfXkVNxXS/y0egdPb5QHUAZeW4+PvRL1WSeVpWFqlFtqdm4xzVTReHtdID6TbBVIIfk/HV
QOKDCwTcgKiY2Dhmm5xAO9dKPJIpZ3GVanNhpOGUAupiHop3wf2qLHVnJj3Q809zS9lhFTWCtRll
CTjjf+zmcVrrsPcvsqXLtzmTMvpjHA1Y4sl2Fo1phvJ8AIsRd2Bvk+ycwShuFZH2iy9dJgmXV6q6
qMXmQgEgkZg44f6s6JEPH+LTiNaPGBxQs7dvg9xbqot6GgG9G1hEdlSdkpJM2ga00/fDWqvSguPS
D8bAz0UmOvzFbhgNa4OsyQQ6Yrl7WHAuhvXzYlt0GvBx763/3Kr8UPTh/467ISlwwna55xzCnpoD
SY+B3nnNTqXtZhXmSWw47Y1EKyQoVlJaTex6yE+28z+0lpcE54/ysFW2t1vAh+mS9XOHxuqlzMOO
PkFxAkrw30ttCQa9l8pGP+MIFHmZk4vlDPNCe30TDbNLDQ2TErTsQC/kMjLmmOzO6SdWoVBlrowO
Skd5HgL+Bz3SZjRmur31ouVWJTTy0FD9/u2V2hbvTdGR97/4BYs4IerkVlsJymn4O+iGRJmmI+Fx
NWeSk9s/gvaou4SkKLDghUn2ojFoea7Bt1c2aUSYWWnDuWI3d8wNSChQLaaZSAMY9fyjisFLWer1
KlqmiL3i/7abUFzpbNZRTzXuoAi9hEs3iirJozuyss8RrwxswVCR0Bq72BZ5sGKOmGPRiLiOnDb4
1Rjxdyg+TXmxirRr+t3QScg8G9KBxL1ajTYri2cjhK+tanBLmwEaPIL1/03G/Oj7xbq9qiNhPl5p
0HoO3UbNjh+Ly/XFIrFKjszaf9WHI6MSHOIYyYCCBaIq9saNT3pqagLVshn0hY4XBMPVu0leZLJG
jDy8xq9QGmrIeWQRB2zWOahQ8L0sUXwUAM8Yfu5rv+DUdE+t7nLK1YxTDBYpdGm6wWoVM5J1DNBT
MHpw3P98k872a5mLVU/jVV2c1J0un3skNrHrryAFFwWUpOB2PvP4BIXzNcR7Rnv8Nz8SI1IDsNZi
uA3iDYOsDKYo1w/Y1mgvnm99Pwc54z/nVEpM+TNpW18C7pZgOPyejUfyl71p4o2Qg/08ID8dhkmg
2gn7yiemBRqabFUowYfPimjjZD8yDJfFlyj6gM4iHAjvEVKPM8Pd+2P80xNbyc7abmTLljzKKpmg
naqKyFfyVK5STk86Y/LP/o/+YpfyoSjbwkuOL9rQxZgvAcP+LjlwIrn+h0O6YLNeP4et2MB3/iRr
HShhe1TO1DryZ9hBmLvdFf5xngBzoitqwmPZTTMAtqkZy8pAskwEfU5xGwbRevDonKh2Wp0gijny
2ZHTI7M4PDoP+J5MbiMyrj7jN3+Fkgmy6RJUrn/W+tW1Hoqo6bmfz9I1VQnRQsHU0NbTUjv6ATvb
pjLgrkLlJ9H8VOLDFKXrHdywC4MectvEqKY8RaNolzrANz2ugdxmVMit3XNvRICkrXFkj6w3rpsR
zU74fbYemazSBmLM27P/PPpOYdKoUmYMIYOfxTkyYFGPhhylU1ERs6j1/QuC3wgqkU4GMKbf2UyU
8bDeKK9XDb58p7B8LY1D9V3OkkojN7Zq2jPMwAnzYOprYW91MOMtPV60TwU3XwuarnEwrKAUHSYH
sXj0Pu9hNHA7HZRXQB3mT9lkdjCQmnju6oF8a93QWEp4+h+RFSWf5iKskc7sxo+6aofRZVFeBG6B
jughDwAtEef6hFuSaL+wY32mnRcaRPC4s6e5nGcN+ZLeyiEM6xv/rYYAMt0KwkJpIS/oxmahGNjJ
kuiAeKoPtpSi4twg360Y9DD0MQcMqA1eryogB5YaJiFzYmGGRIuTGu8ak+jrc8KtDrYx9RaGGhaA
0/cDuXhscGgTPbeBP3rz65owghqG/xxFjn8sxppS0jx7rRyi1loMhf55nt+IAiBGz5vA7sbi/MIG
y5IrAanPUAe/Sr8rVJz5zg/4SEvCOLhGWh2xPKipyGKJjdU2SDWH1vM39lsNO5OUYkEU+HLGf/24
ZBFwGRwyDCEzRi4Hbhx4nbdULT0VDw5b1gVLW8BsONde3c0xf1XwfDIICrW4ZJR5iETa6j8iP6i+
lSfcLtt1eJfZ6jWi710cl+eZKHKx6ZOaDZsWUVI9JdotIb+n2K76Hp1j3MG/1Jx0dLlBVs4Hox9A
KJGTIto2u7uM8KUvAAk17pwY/R2aA3sYxlqV0Dyi5YM3bE466gnG3fQvvEwS5JaBLcawCMzjLf37
tksq4jKmwVCqKKxObOatXHQV/kk/puMKqagyM2VqGitguGLtRJ0yVBQeV0oxQH/uBOj4uHlWF7s1
QhhdrCyh5FcoNqwhJxW6JTBwuQZVeHQ2oYnlsm2HvJfG49GexGWk2qMyEtjGko8eLRE+AyAH8+um
7suNU1usRO61Yh1HLqAnoOMl+NTyNh7jImSb/kI0orpSpJ9oARgR/kvX504YI06jZt9w8Vnz7ivc
6scMnCIVO7RclYI9SdACPil640vSHDixaFDclZ8NmcBk3Id8TAqO/c53huuK98JsDZ7lAlAVK5XX
GIiRvOezcmSC1BFCF1xZzKNfFZ1wJvXNiMpZQ9K8UFZkC2NIMSqGeFkAF66F9czGvCgPY41aV/CL
dwXXpiVzfxeAsZYDDmxWGpxIylIk6JJVGzMT+GfmlkdDcFhCcwvNb4GPytJKHvRZxPOc+AOZr+Kx
132zVxP/oPu+tMTjbdpfagZamvkUjGIgim3Cukc/PUqYbpS6AoOXdkMFoyD6h6dltDVvvmeDReeG
F8NoRD/PW9bvPH2ff3DB7kmJgpLXGNCEIVQxewm0vAdat3bGh4bzLpEDJGm+LKDwtJOJxLpCPrR6
SeAxL4p/5k1+U76E4Nx3m9gHdHbTNQBPgLkXYc/DMuWXS4/ftvG/YME2h4zYeJ5p34HO56fDd2kb
OY/pWNeZHl3OwuLlVsuA7kWpco+J2QdKerz608oSQQ1zSOgSko4G4j19NMP1Vz5gNcXpnaTMV/It
DbKlP80wTCDT7AaFYW14u9RDtxbAd6PXRKoaoSjYGO/Gk3ObNd4c7E01jZl8TJ2qZhr8G3ITXO2A
mgQVR4SL4+AJ6VOdA7wpq5/g8hgNEAH2IcPN2LD+mR7wnc4VKhZEsG9XSm+fcSp5u0RMKgK/herX
17ixFsVgS6TFSuD8VrGregbS/T8fqHrg5fhr1t597dlfH+AxHKhfKkqbf5YOwQF8UWJ2iwgh25XZ
3XebRm10WpljOLJN4OQGMK77PP/FK7Zcv/DtOlGDzEWd8/+u/4+cOfox4URgtujcw9sKljRR4g2P
7TwM7ZJoltEaX7t6jWdglXyA7HbqWJ+49vvBoRS8wWPCKtHp+z8hN8CZOnT//DneTNDO3vxjTHw9
z9OF4C7jEItMt/DQQnljQHHuQRPnbYCwTS2K/V1aJ3AMaK88E3is6tC2aZIBBsAklC+8d6hX+OYj
kgdV+JblblTBq9xzXXZehrT9Q6MFNBcejUOeZjqcmgtT4gqJwgIPFTv6qb441RiJInVWhW3Ak3SG
gpknMGBJjqedlmh8EHHlzompoFzkx5OyU2/WnohaV8JLIAdfgABB+9PZkEijRZt07fazvLJUN9fB
aib5WPfpBRAukpKSajTdY3mDEG/5Gxdf3QEK41uhAI2KnNgqkU/GF4/8FUmC/IG1j19pKhTw7HX+
b9TK2LK4qrpVzDZloye1JsED+jOrnPIPFvloT9ykmGJUYToyIF0e0k7Tu7Bg8IF0B1BFHCPiEvnr
D5TDRuweWMrjJg+EQcRfIUAsGm3SDxGD+emZkV2LQlbg4YKDmKuj3CrCJeSMXPnC/XpTel8k7hIG
ONdXwKlddpXiFl894WALTSwKRkFUOQKz7iPROTOlpjk/LsYuEpjxbhzDoMHz0DZn054ug9c8gjd9
7dtzfr8pn5dUb+GQWdFizqSQCNKCCiVrY32nS4mJKX1V3NctGyZYVv2orxMogNrgjyfuAYY41ljI
f5Vhx22I4nsctNz41pkmXLHrYsZBbUSApsa193lRSxa+J91Iz9scmQUdvagSoO3gkOoeEm6i/rfR
iePy4M+gljCnQImu4mKzlCIYL95eyculTrpyrbcNzHr4+2+fZTSp2PdlUrfO7x6q2agcQvFvPGZz
N0VV4gEr8u7Efy2YgV8LMh/w35USDUMgBQz9usi+yXvcMDAHnRIBW0o1Ie48o8Y29mnqe0PHM8tX
woQsECtkm8Cw3CML2Xcp3io6EtzX8WYD7M8pB4mcyCEO5EfGNpIPIT5CM38y6sYz7UqlziA3D6R4
ea5BaYG7Z39N4YyPxXExPA61QjAbaGTxrCBMwJ49sIUD+mK2ipt4Zxg/VEobfT6NPBp8qFY2xtO3
4DPWV4MOnPBqgD+jgAfhGylC22OlGV+F8x7DiKLN3yOKkWHXcodYDvHEotib0B9//gpNTGTNjNhz
7lsgAv715zogDSh0kuA5ZW5qAz+QQPH12tWEqGCG0uo5R0qSEW04unHPGfjTKRcirLfBSYg2u89G
tTtsIlQFJqQEpFY4F4KUrakdMjGVjrraZIDHO1xzQRhUAKOZcUzzXQggyothyqzR6vg6cTSExLy3
zBW0OPSli3eCc9Y7OFsENeJNj5owmQBlc2i+1ARz8ux/bPNlvsES/LgWxfvZxhqFjABMLp3kYCFV
wmO3HOZRKV+CAa8Vg4si+C8uFUAM6796fV3QuawZwRQ543gYJBnkCTQ12vxZB+b/Tmg/WpSndYXy
ZU49pgk75AX2xsPke3glexzVJuKp6fhAxGrf+EKbMvIvkUzokLzVRIVfY/vEx9H3EMPOUchNxFz+
Htcp5gcc/uYUZC9BT+2iIXIOr30PLzqQsQcZ8NJ2MeAfpoVXSQk+823LxhpaYqQ+JvDGqfUajhpi
I8KUmbOIU1vZ1A90Wlvw/Ebd1fG4/9PftMPZXEPevtRLBBlIbl9BSgcl6smMPRsVW93GLgvPee+U
LlKZe3Qm7/+z1fh7YIPsb09IyrRU+PQpMyfiTPe4V7/RfUezMioqCDYLu1KFZO3IP5ATrv4S70kt
Ch4JJcRpGMysGXJLohex6BImr7Q7Nn05crBHXlGm+b5ptfZbnVfx499SzKhQBgvgsSX/qL4pZ6Ja
5G3uGllQUCE7qp39M3uduv3aEAirjJ5qwIAvWTfJVgXB2YffuwsMeuav31HalcEm8aez0QGknW5v
5sgjXhfbNADK27F7R+YwUUUV4dX9I4VnSeApERE827g7i7kxt+2OXLhNLPpEXIO4f+4oKq+H4V7G
tZ5+80iXvXsVW8ulo1t8Ox1iRhdonrP9BYnqU/Qq09D9ODZa+zCM29f8agQp54zLNKkTVQgxJyOM
3piaiAe4H353u6E6c6X/o2OszcRbBL+3ayuiDLfy5uZnLa+w6EgYhk64linPT6UYNh8+fBbgghV5
u2ULyhoinePRNyWrLZXFrzPQm5CUhqj3MYQ/zsDnB+f+AdxwZ706ocjm2agwWz0PTdrrw1dyikp+
fSxjiwvxILXAWSezKHTfphahNurA+kr3iMMSJ0lmalBzmTxYo680VLm+jjJeb8Dc0s+LzYjlBPr/
6oqDx7I5lEkaydkzAZbTQqpofaUdGYoM/sFntD8+6P+Eqhz4FjdCQK59rxC9KmoUtnmpXeY51bbA
Asii9plhfHIQYQcQQmkdRDME62KeChXC3INy9HThSwv3SLafzcYUDtCHwafuuivhA6PtsgVe2Ea3
n9BYDfs0JWe1UmiC8llbYRiR8oGr0gh66IWRzBKxXo8sZm8tBpAlpjQiN0ANlqZQH/pjGHgSMwIn
ocTkI/KrqSy9a8kg12qsSrah86ImzD97GM36HmhCUEHeii75zztSm37ZYoiHWNFzuJV8a8pmHPXm
YIb8/lLSxi2ReHJnEukSDSSMvk+uzoIPFUMvzmmprnN8y/FTRc4BbXIWx37xJXpChW3Qlku6ulds
CtJdbfKJaSPglLNCY2+PwP7ILPypdSFW5lDiPQCitqjttpY805uFmHQksZ9xYxQYUvJXMtkHGWcj
yNNKJxipHUMbnz5xFM+b9LMtVBhxcYaREwkA0IHIH2ofk0K8k1R+0EsP1w9za2nZHu6etbRlhJJj
apgD3dc7EqixvqXmVBmh8IJIcmlai7o5ZZKUwC/Eba8Tzb0R3q+2EpvhCmGmS61gAYoovklriohZ
K2epWJWB5BzxnkUu2XK+CvkOxRch09nV6cWQSxgUOw4a625N3KYrTux5SIkqWbbhObJiETWvNYaV
ew1t3AY/pX9kSX9bNK24GBlrQv3pjnz5JwFvCULT938IWSpDxXtIV7ObU+vqkWi4ss4bQPmVvyym
TRzLc2/n1kU39uUpYEmJeKHrbnY+IAhMsuAG4uVOrfkL9X/5FBo6lWUiOelM0qzG6ybSUx+89DLG
KDJlQ3ORwdAI7OEh4sCzdGls7LBd/JCxxIQDbTKfDIYopkisGdHPT+U+nwDnDuj4mM7cSOeYlHc+
woiHXqBiVYU0ryYMXiGcBLhwGVk+AOet+JI3C2cPC7S77BMYcIVcHTcoP9fFqeBTsqI/rozSipSn
Alf/C2B/nDrV6us+5laAduubMTH8hZbCQBj/6TMdN/W0owFSk2I5aBn8dawneTwGTprJGAvyEX31
z31aX/T1E8oaCHOVeBJqlMn1Z1UB5fpHDFemG5215q6WscYFXV4goq0gUqL7EC0SDZcLfMseTf4A
7UIg/XjZSx22OEMqbAV/2mqcSDWKh9x23BQHjrwNuVUm2bWrNkbaPTl0NaPAdFmgmGSWHJL9L8kX
WitNWv14lTJ34NGKodwbFRBSsRs9tp7jM2Rl/KN6505bHDzFpjc/gOeWHnblMAsM4uN5D1KhlxL0
39linQx6zCwVeEnyhYE0SSDTD5mOw29ZZyUkBC19W6CZD0WtHZ/kocJhiX34oW/WNPuKISdrbfq3
cqADNArJfH9L2ESBCuCJvox1NMTxraqvLtRK0nLTORJgcmz2y9/s0rQX6LbCT831ZszHOItyWoK1
NmdfN6D7153nqE9NcJINlkr3Fm8tA5epPFbzB+I8OL435iKPueSvGzDgLBZkRZqQ1agWbahw9d7A
hLzH/7poYnZPHdKX0B43XewKx2T2v7MU93rkSHKON5gcYEIWkm+LYcc9n7YzhGApxST0p8ZRCDKx
ED4h1u7LYp71k1K6tL5bZfLLg0XOgW4Oo8UQFT2om4W/jc8abjFU1pdMZ7k1p22V+Ai4t0n4x7uI
/WHoB/tm5MD3tRf6Jtxq9rsTGQMUm4+GldRckEw9AZCH4x3WzerbC0CyQ+rOQnHY/5phFyCa896G
g+NtOOwQyW6M3nixhzX/D059v1jqhG5EewDVceX2vQHlMiaaf1Pp7/y1NYnHWP5Vl6AqlA+gEZSM
bZGaV9zbs4w5Fqc5yhOyOiN2j2riWAaYyyAMQzbW2Mbj9FTtMfOU9VVas9nhpY9721CuS/Kr/52F
6CxOoyADw1lw/poac9ZbaHUCY+7IGc5YxB98kCgsO7qHxoxY9hSini9Wz8D3N18P9XGiuC88PF8R
NQCAyPF3do3k3RCHMU1e0WWv9jcRFcBkwyniwl1391i+jmGNOEXkjR1IR5F+1Dwtnf1uYwdWlrNS
cML4pKGcBQvdCIsa2vx7Fz2iELBkVMUhVsa3EXjZocnEX+BLmEH44zDzi04gqKmN6OOfa1b3P7Tl
qtVXKPYABRxlXHaBucmWVZoiHnYobcwPr1141MDUIG5THkkRD5jn5gQCuH/xbcaxxkD3cMa0aJpf
/U0UUdS1LE46JNU/fbpfi+uiyjqvJvKPDKbo9ayx9U/QEEzD6DgV+TdgdL2GSIna5tGQAp+V+UE9
PmqmwCQQO0bxGZiAr2jN03z2repPL2GUHoQ49y+879TJPi2O7vGO1KCAqbL+8XaBvnm3PeecxrDT
mwPXO/XKfVALUO2I4PZduyXK185/K7HYah1T8azBNGj8Pqp0CWLGlp/pl75mu2KJ4WYOoVZgsNwH
QfzpTjW+Gyt69Anr0c0lGrG0yaE9y64GSM+Zg7FmxveG/yJF6vIUr5Sd5YMbW+H1/pP1NPi1IT6B
um4AivxhyhJGQ5zdIhOEa1e09IeoARX8d9E2ll4mekmOBRSJ7lvqfBOfdR530VSgor5D397ozdA9
KJkegJJrF5IhZItlpcCVfR6vS279isPzjj2s9IBDCF/UAAOQ2lwfi86j+LZDLHydmv+SNxuLkgcG
mg6C47Q3+pl+rAasMOeXjFSi2J3TUx95Sd5mbfY7V+mM1W7WYxKUwhE28KkziyasSvenT5ai+UEH
cnmRu3Q2CXjnk+fXsVx58X0pL8z3puUFKllZ616JiX9Xjm4PaRSyyA2bTIP1mVJDmW7zJ4k5dEIY
FT5nRTlxHymReZRQZGx4CfNlGiO+qHhghfkYq+be7qlLj0HQJnLSAROpPMcYgGfL88ITTQ6uT/76
V7YExTLdz4u/QAT7r60JUW2cFT5f8fLVH/OYWhcCgMZifqGHCWjFATtFtIrtb6aSrgT4pT+BtErX
2C1XE1rZJibsBf84qfKdNRf1RktIoV/i8TLw07J139Sj+3W83c2Tg7HXQ7XM10TTp4T7NEdHrQDc
Ptkn+Q2nVLraA/bhAtNODhBUuQOG5hqxhdj8PPZ4svr4NFxQp2T1kQqb3mg3g9QPiWEWI7MdvFkw
TERbyVXZi3Adud9PRUMmYxOpxwa2wFtg8hFSV2gIO0NLKnzJBIffGKBZuXa5ELzjdLJzi8wm/U//
VR6zx1eB+hVPnw/Fe+NXLxh6vkRLjyz9ISpx3INBLEqB3UODyAchghrxNuNY248dbluUqMeNzUUQ
TfgTiUD5lf9M4pJ12kAcB8B0apInhc0bnoJZzZPRQf1Pa1D1wLDZfzyXgzayYbICbmq38chQbXBP
Wa69HqoUYQM0MTYvaSzYq1clMB7hZFRLaJPEoUYAs281BJlMXYN5T5YNOJobFzKDvNj2tx318bNT
6oEmkQ6fp6d0RAgV7nrpUeAvXC+mh65CYSuyC3RSHRsX5A2O3+e/XaVVC78r1d7y6riy7XXQ6aSt
vbVDGIxoAo7qVL0XuC8JLRmUv9BY20Eh7TmNDEal8ThgSjo7TBECOSeR4TdOVw3jb0bYdmX1hiq1
vb0DJbU/YA/YLzXwIWglUBVwSSeFlqCCuiczz18TcCQWPBcNTou3mN0YwyO25VrhwBV8vDls/PFc
G/o5dlpAfBsJEgNrbZkfRpfMVlsbkZoEcVWQXIxOOy3rgTLfmATwkxyO59dhmFUN5rZ8HpQPC0pT
okm++wxexgsVJe08FuavzH+pehpEUMLahUfatkepxdvBk51HKo0TLBXQLYvOZlPB9ubiRn2rwsOQ
s7+vMJs0UzSGvWOKJ5vQuI27POmk5AetzgWPb5F09Oq+KRGwoN7z2sW9noXa3+mXYD/pgTR6IWtM
1ey4SjmbHzAva+pEw4LISJH3HPs//hJduo3NOECRJTZyKMOx/euPHSxWyuCq/G468il5FT6Mxhez
f+nol3KRX3hxBkuvPMcie7jM4Yg5lYQpypej+BPj3yg01IKwUl4qgCW3HsrdhGZ6CwdU94I+TLDw
j4aiitH7cdeQIVuy1blI7Yk6yDkehZR2qHnoTnjofc4lFUlWIWJr6/LRP1gxUBZrREGrX2acqJ+1
sqDPgfyLbN86+7HeBp9Fi5D8fwP5Zdf5K3ew4oAna871jEXl2xf17XWnjPFF3uPo30UqObBoSsna
8qXtygfyV5JIehQZ+mUczb/uOBrsl2p0mOdlVtMfK+fAz9n6FJ0eDZVN3FNDUxsDiXklTIeH0cAX
9LCyd7EFwUpDsy4xVakUmrTU6kyJcETu2S8vds++IkIOcLRGYGPhbU9J4ReO8Pgmgv3CmFYfe+6N
k4NsFUwSqRVBYKAEDHcoz0h2pb+lOluddOejB+g8dbUE7y9gcLQrCi8iqxeOjU9TOJ8jK3U+Ayoh
kfZvlDvS1aiJHNMYECdssCaiS+vD9S2z2TbGOIoOnDN+KhxhV3bNj6qxYKCdewVwTWOMzIo9jqPz
e4rZclazD/2bcoeKvgCiKD/QWHJJIeC6DorhgbSRZ4tXMJYM7IxmUs7vMBSnY40GPX1kX+c+vak5
/YC/ZVgWS+dPNyH9D9gdGz4e2KrBqrJBF0HrgqJQi6jx+xriMOPpqRozwmJWHr+76KDtQk+9d9CF
cS8h3NPMCzfwr3ZQ84urKZKfpfNxiZr7fmRy5zhga7VkEXgD9J6ImGWkM44tWRP1g776Lr8zWh8c
VOksw+26It+YTHEby4voRiBM/fVIYvxnlbIjP8v7OGlEvLqaTgXEhm85X798O44vLD5v1mAI6Bfy
49j2hCaCfIlc7xxXeGwYiTpy5BdVE5WeSkefrJvSkE1s+IuRvsIGocfsJWniyZumTdAe4wJfsxCk
u2PvjntUfTcCBZSuNmQcqDPBCeYaILRC+73yiIw9GWFKGYY7J/OH3bg6MJqBxPdRFYwxmfaqGFgQ
CsCPd5ir14s8cjgx1Pv4QrJHd9yFTgxEpVqNRdlwa+3NqBotR01kRr4gMdCsphpjnIrKc4V4UbLA
sBjSls2YSH7lJ9e9/8pLRQP9HOyrzSYQGuVSt4qyDum28BVcVY7XZipKCV3wTm7pNFnCJshxke6z
nfrB2wk9IrboQ5mXRwE9LbNyQ+kp6LJhhCNHV3GG00BeFnpRL7Jj/h1x9YHYIb2ASpqbspFOZ8RD
nWw1+yfizVnCuV56grPy3hT4220sciC4L3Ps/00IWcf6LoDdOYkucFkRQ6eDvlDiKWr5l5c1v4/s
nbwLzUMssKYqYZzH9ZwPUVYEh1tyTa45JcPJhF81H1uDiIVqCa+mvaTx6tYlHIu7L7sAMPYP0Me1
8eB2fRZg5jCj8sYR97DhoanWwy2afH9VTlmJzv/MyNjI41z0o0nk7VJnwyG1hZPERIgzclqwXven
0j8JXBxrwSNpOTYcQreZ0c26RGEsatX9SzT8uXXoFJsSHqecc7P8PgDrz7teeHLcFJjdWO4eD7ZR
Xl/CQMUTbpX3wsRl5PYr00mCKy3I/bXpZtou6/OHhrBt8oIoSHksbV5Sf4WYkQVyUR+s3q3Z5rUr
SOoBpb/Iu0t/vipLl4bFXHKszmPmCn13cCyNqwd3Sw+zmSO5xsuqTI5Iob10NzmBUQtUcDBm+CC0
DIcoOm5MDFokve+BKF45TOcNGNgojCU/yLfMrfex9WoVhAyyuxB5WsGrYL3F9Nc6qdTVuGYj6mXT
i77WNMsueGoOZUQVQrNKFozb1kwG9/5MUcrsF9z9OjaxKnKMNQV8ekUSzpVrX7GXJsSftbIJso8q
9y+y0BROVgq+2i7B3KcYn8k8G0Om5nIg9mxx4avNFJ43idVQWpeeKTA5T6I5vHP90FIOcHosAZ94
Zr2CSYe7sE6fxoiU76ZIH3HBbxMeW/+r+z8LzHznInckCDy892Y5Psyl18a4E0T4h0HZnwaYG+uZ
IYyzhC5CiWaf7YX9gvNokAxfnZVr0+7hKy1LXfEF5dTQlUrzpZvHVIMRiQAmW3fj8lnB6pt0M7Om
LYqGsETfcoOgY5uqi0yfcRfm0hIlSAXII+u6h3XCqlnoikwx3Cb5czRqKMtQ2f85/srS+dz8i9Lc
kK85ubHFyaXNIDLS6GTPyYliy/4s0o3GcBF+U8lJpwU/vWwhqXSJ9ZTKsuhozv03u4vLdcsuV3sK
83CqLg0Rm90VBowQaof4zGtIA/nR4fP/Kyw405oh+mw3oSRRybwghSj7/LZoLlgm0QhSZZmnjh2f
JTsDT8ZhGyHNrGSfecZzkj7qBQqUNaNeNXJW9FrCiy7W8NyweRybOLMrLFbPaxUYObEUsGOzxCl2
S4FYtPxJ7L8bsmnMBwdPzHuA5qXnT1yKWg0hEFY9dwwjErQKQBc2HF53/Jl3qOK0NO4p+z03pIRG
vflV52zYyR3E0H1QMOYvp06idqmQ+mJbCmhVbpdOiTBi1SDj/Z2VGXZ2AzGsVMCeSU+DBrTVyQ58
mxzUX2dAQYR7OAtngBzclC55dF9K+rt+cfX+YqHOd0po/fRefYQTe13dUh3qy4NwwFtcpDq1EaHP
y4hdvlwx+MoJsHips/9Zagzp1bqR3AOSRDyLmQv6nZFKbe5ci/XckaiqUQGTR2WaMO3scrYmhCm9
LdnfzAQBDH+wGiXOfq4jluVdelnLoSPfkKObHRLDeOrVeaweSeTAvbBaNFXrw76hmTpUCEChYU6x
WIwIDJI+k6sbymshPLV1yeq7xfkuVvO7++qWmtBOIlZd0FyfLwiVovE1i3rqYSrgAtXkGdJoOyrR
HWqEQHVq+Dg3kfJHxypuNOFFxyI3EZEX5p0QHi4BNP3aWEm42Y/YBM+GaYVsJG3PNK9VNNU3L7Vz
GN+fSy0G0zyyso0x9JvmeoDAgZACJokICQ/o/Wrh1hDZLU0wEcjCZlInK+O3SHuHhRnpXMBB7DU/
RHZhKGgWZVfp0o6qBW54zZmUjTMYmUBOMEKsb7aQn4FnfFJXbOPlokP65xVrmDVWkB/HgjdM4cJV
qzjP7CoFt7uEhjfGlTzMhF+c1sd9FmPCeYV8hb6Bc3LTFy6CfDuvxl6xVQMew7LXU88zlrbUe5tF
oO1QRRuOZAD1kFpYMKbReZ1Jb8JLYga6wucU9VjaTQFFf+DQzl6mM0aNpKzmBa4tsc0nZzZRkKmh
MK5Mlh75rWwt90GF5/VnBgdhVa6bM7vAI/dSkvhBcYX+8WAWDaRpH1vG8T/DqhtBZRkdA4FX3dze
ufgmLGaZ5Q/q8hMR7A7meTfoqHPVRqGfSYJpXlTThWUmPalqCfGAglkxNgjeL+Z060ouzf2hfwdB
EIXgHlInKuVHJThcOm2r9Rwa0ZpxeRvR/Q3RagcDP3UboD+PSL4xuRU2VW1lknWxwWSG4//aCPyq
c9hpBOoGceuZBlaX4Hq3U3DWM5Yebb6dOlcazI04ZkEUsoZPfEot2aedOX1XKX7XbczGdMpUaFhC
YdIL8/Ye7d3pV4cKGfrAFiHEF4EX+09dg8t+8gZ5KJIT3z0pI9YS/FzD9+zt1nYv0PXxNtbFW48g
08AneGQk4Yn+7rHpuTDHq1S6qyh6+Tn0XCMqWT9yrf+KBXiXwDSuzfv5oeKkCQDjrERHpvO/aBip
lkpONVgAgbuPxxz10ehemRpPAuFtTonq5b15xY6ZXo+dFcYYTbROxxOJFAecfy+zkN10RLu3akJ3
eOS9icZcYtVCjCKyre6UMeHPH2BsTd5i5Yc0eVXkRoKT38r89qGacTHNYgcqxVAX4ex8Pb5352Po
x8d5ZhXV8rr1nwokpbdLeSptOhhYD0MTTgm9BXkYt9UGu5GLwSw8RzHunzqc6jNIYvxIhldtxMMB
zIO2QQucdHUMnv9Pl/+7RFHiIrucWWJ21g4bAr6khFAv3xCNDr+b2MlhlkqQoYfbeozvET9cVoB4
WVI9mdtkqIJg2ETkgIIkF4CIPPlcor25CQwGa6ldLQRoFJjpzBuCxnxhjcd4m/K0m0x59mixEx27
Z9Jwc/S2TUP39xInv1Xm+/GyMIa/bEa1vQ3CsKu1vpYMpSXOiJzXgHIiGbPSCAYs1jCy0OoZADqk
777Qbq2rnvzrROQYmCWNCVdPlVVyesrZ2bE4sns6seFliorqmRxzuS28or7pqjCY35AQV4fH7NyF
mzUbn53hnbWpNDyIQBOXrXEREab+M9ZWtzw/xMAFHeoc7AP3BCvdiMRCCWak+ONlby3PMbdMAOfi
xpIqcR2gK2D8QzqCx8iMz+amWaSr0nWtnqSFs4HGnXgYhrpxEmuWi7CaemiRqgAuzWPyRAPg0E3c
h/AacwxmM+BiCd2lB9LY2S6orxerv2n81txiysSkr2qFSOowCpQt0yx16IJYSpfkZGmy0d9dgXJR
rBLppaeWR9uaQoxgy8bH3vssRTu+JGPQiVfTeuBkVbECvF3zVmdK4xcGhH0qGDvqgFO50Wf2/3im
Al2+aYXH20V7VurJtHNb+8iUTLTIwOU5Lsh4KhrEZMqv9IRLlq85Cul14ih6GX2ap9e34sR0Jmg5
9HYZjIXg0TlNAzLQ3ioYtRLQDCMw3aU6MOoR/WUTdJhBHgNYjUQ9Wj6qIhGGyHsr0L2Jpqf5ypjB
4mgq/vFa0/4w/iGLOEhu5xV3/BTL3I+OyMQv+8CdICXh9LEVS5/aEbI051mOzuiKPdgDcN4OnYg3
uWPZI4HMhTCXiw/oDeaorINLj5M0tmyCwKqb9H3xmnDtBJqOCaWjWCWYI0lRIMzeTjR5mP6VaYV+
2uf2RJOjJ9egj4SbOMj/6m2clv4E0zqBS3afDxODi8if6pb03HiJ1KylWok7NijxE4FG+d4JPy8T
aK/CuxRFtn7O78N0mGsuM2u+zfcRqtipTfAEUkF3NFzgafNlx4oZ+yfj7mE4lQo3aXdKV2ouNl5h
D/pCzvmR2x5MLhjTgBtMhccxFvr4u6KAP+uA0Ae5dmydw0rLjN0dIqXJtzS25WmawvXJhPRsYsho
ioTFwJ+ncyx07q03FjmdqUF6DTqNb2gO+huXretGdlLqiP8auH6DhXyEgGBQsVFivHQutKdrTteS
UVXqEgnRrWuAEI8TvnkEf/OGigOifOw2fBz8hUMIo8TMiVQtzOM4SMvNgVU7OOJs1zrMs2vP8T/t
43taO9R4b8wa9nBQTG821R8h7YKZTffuHBTQPcKcyIMtczhkkAiPQAosRGf7GpjWbw0Gpwee3l3E
vVyayGJ+lvTHKCRvSl7uOL9Kaz6MyPMEqJehge59RPNqUn4Weut+roJeIn3+TJSVlkUM+cEvUj24
/08Idlj/S9QGdNa7Ntis/4qgWFA8F1bDJu/Ql+fWy/RI048ZAIPsX0NOLnib+5q/Pj/maBWy+faN
v0Qj9Hrp/J9luMaf+iH+nxAm203j/TF514Du0JniaBoPpfYCTEeVHEoLBZqfguo83fhrV4lOcpZ0
tAUCgEl+peXz3/luS0AV9BuiaBDaBRX/Qo//4bipVPmvUzE14mFBxYkhmz1HKomtQXcK8EYwMMFQ
I2QRLnYZ5XOU2lERQP3u3dLZ4JLw4kpB7C0jg3ASyoINd3JuuA3gHe+H4ruVa6pMY+feMadZyTyo
yPZgZjNQxCAop4wxSzaI+t3Rv1B4r2JOSQjvx/22JQ3IWyHVVlHNTKkUqH6epWSM1DTz0h6a3YHT
6OD3kxgOrpFtBjx08fXsbC+k19sWrRGWdG+b/rm8mO9qHBJ5y452WqSUBu6eNcKY4MHFRnz1ZN4g
JMcavI+Qow+prHQSa6uWnDw+fZVWXsuQAmhQobCDYvpD1FYNadZzogvv1Jf02UPGwKwejeqFwS84
GTVDQIKMpBzVVk/lbeJacGz/2mOw68Z95NjFiuRjKGbSW2ze5gmN6C79iVODsfKE3uIgGPVWmqVT
r4Lauw/57zUqd5POkOzrEJTRHLYJU+F15LbiizU/FtWYeJASNprHCc4MrQ+6e0yQz8lO+Ns9A6/R
B+m4lU+AQFBXUMWRc63bfHgZ8TkTPBVNFYWo1vW6PxAlEdaUZKMCdVv0qPVE0P/kGDGKdHh6DSHO
zTxF93wn+++RXvZc7dV5Ii9ALSX9w6kmfHnUr5P+tRhSPa+rzSHQZnlWBZLJ3Fd4dyN13k/EUlyq
6vEPQ6BLTXMi2DhCr4FPwCLqs+eDfmEadHZoAEz3q4C2Jd0qN4vyDn0IUfBupQliCIa5RvHniX/h
nGVH9JhfDhxMUfEscKiU1HEYp+B/1JEA9cdfqJmgoDuYrNmdm14/i82eUXjYyeU3cnW9dzCr4H5I
wwlB9lJRsLBc7faI28SK27a4PZG/YFHT+bjLNKG60SWLoS+g7aViBizEDRx+4TtSlCi1fMBLUir8
m7Atkp8OyVd+zFRNNn/M4oGQ3BV7ExsuvBUlj73TtaAqZl0EoTEnhJ5YJAL0ZtF8bxSvwD6lI2G7
y8Rb95loMspqZciNhkjSltVmShqz5kLOtLqJXXI2uP6wsDBuHXVBJOF39RGrt4Er6WMg8oIV8w2V
bvmQY+zDpHhq52ZnHQHPT/cClhzujPYg8rXfbJtShFIxtTtNkDZUVo7Dxvhij40KNJryAIPEwz0L
5UXO9WSpacNjfpD/16bQc7TBxVR4YYIHyEJcrPa1BkCju7nuwz1UzjlAJuRvLFrxXkq1YUHhDAlI
+GLF7WijHqbVU9hx5py41/JghsZEHsLXW7YaeQeFlkRDbNdp1SjqnPBTOzvPm5hDsnnSkhSBKKaC
fjw246UD5DG03aPgvke4mW6QIJrCHOf/0bwDeAAN86NMyHWQQaVfUDKaXbJYJAlpRYjr38fnUrN/
5N3UGoP6824Pkx8eUalUmtitY63VXWgBvEMdr2CLZUBWbFa8bLgiq5fBMR/GddgRAKSxx65N/IyL
j8/cdji8NSe/8yYEKanFs3cGzpkibjh55R5x9NW1d6HnAQg+4/DbzwAo2TD0Q2Q3t4VJjJbYN/zY
Xom7siU+jcY8m6NNPga+eT5wdewIdcQLAW0kc7ezfxh4NcaPIPH0mo6L1+rgTj7e4GxRlMPsS4Jt
MFiWEqfR+Pa9RE1NG3JNoA9yZDA4kK7Tf3YAh1Qy0Q8TT8bgT/L808QcDzW0aFJQiAYPf82JkLQQ
UvnqdGSBWpqCgmyTCqsoiSW3GYW9BfHAxmnV0bracJv32+tFKcLjkd2ZJ7a0pzr1BYmQmVrzxy9F
ouQHWtH+78kqRyHR/grWX2Znx+EA5hABYWcsKNhJc4QMdEOCEVeLbKatJGa7IV6TKlApSL0OaiDE
JwRC4faKvXg669NjTE4BvCiIEJ++66M+TL8iQg5Awzf7nYT69VBeIwP3NFrV4kEzatum/8zP5Rp8
tf6DZlC1tnDXwJRKoYRnhQedzj4UsjA53QDeofwav092KYqKqjY3AamurCuBSRtJJEwy3+gh50Ja
ROU/vQBmYEuxer4RR/jFC7dUBOGe55KiIZwY0tz+D9bKjufmpQMoNEwyGqkdw7A3K4iPadbXUohq
b/fxTinsna+cSYv3SxL7vV/iJJ0k+F3ZLtxEoSzmweOjZVlcCVw2EjUN3rkIhSqNrt7sGXIAnhTS
9waGHmFrunU1m0F+05rlcuR7nYjL8QWzgp4sMTQWV0aoAThgvoqNnOfcqEO1bIHt389AVSy8tnqP
i2U069O7kdEJDLR2rusfPkLcZO00UwajowwgWWBVhr1I9IGN2Lta0W9oaS+vVbJsOtcmOGCH5s13
K4nVVyGTSJ9BRyL17ReuYg962Rb+OhETr72TSao16ekaW5xfjLCgD6VSm4B/allnBB1KFlLlGUFN
e2+wElB7x+R1UhaWomx5d6xJ4l4nXlzr+z+IVTD38FDMWyCiXJOre23wneV30ngfFiTbu0GrCfFk
3HDZpEVhU369+PnUdd95ZAV7zWqLBNkEhJhDDepq14NNZbj9q3ur8ensygCwbHC6f3d9quMsguHY
W6uuFW1AjDafxT2bvvWMadHM4VgUrdLRKdSH4XOHuzRocQZ4PdhdAKEl4x/jcNYMWwkPSwYXo/Ro
3x3g3KeqVN8hpnRiJa/wn2iOtTW9+bTQiUYseXseqOUlfgEG7/756RTYMc4DZFgoApbCeyFe8C4b
5SyhWPJqgiO1lKG3LELedilUL2smv7qN5ejN4P049DybN4xWlDNMpY65xjnAz1kNUzgQ50PQGRxh
T5sYu5/Yt97IaxN8MHDolwTpyQngkYXY2bvmiLSmAgylykxJAOpcF66Ju0h+QpVvI1iicOpKnRDq
FxV14m/WvOaOtPgsCWVkXANVRbPQltzgyUQU0hR75pvBRZWZhiC2p4oUoeuAxc0QLTlrUlehb5y8
BwCIEkStmC7Eg21K1wZvsCmpjRnEeZSaS5nEuLxzrlSGLQbMmMiXRaxDxv56hkuT3QPfdnSintJM
PjMgyqAmvH7l5a7UZxPqOBWar9ILP5kNEFrDpD8EMyhwtu1LtwMNxZ8bBQ7eYCM8eH6sxRLTE27r
nMwTGS9xAsD2heKsSa3IFuMMxZrn+cizE/bWgyax89USoHUQ12gmaz71PuLhJL1WvRVU3e0ck35W
PE75oyPO6jI3NMdoL1kN3wqgwALKf4XaYYW8lO2XlvlFmw3jjoIQPvWqXXRliRGeApToULcWBNco
fL9ONpKHZBPW8XmIhR9t0Ci3W267NuEos1dXqDIPUF5OYUCTbTr/Q3kMq2/DxYTicYV3TtrVJNa0
XqKpC6xf1baNntM2SqOu88oZ3V4nLPtRqPEon0wztdmBIo8rKyYDKKDYymNIiI4saA0SLXtlVnHc
5lQhYiw8vtyaMikGqM6R7O8gV/4ptpXJs1Kk9Tad4YJl+xqvvpT47diIdUIwJ3fhE8S/J3efX8Pu
QTqr5F1jYwomB8bpBBFKJRYKYZ2Pbti8qqQXsTx7cghRQLYwtVFfsrpCYBQrIrcAMPwJtW7FXhyN
1fQhrIZgpt0h6Lb347rzFZlvYZao013Gf6CQVm9mepWiucGHt7EOZPknEepeZLtJfcMUWKCvnhDR
8RinXNa6Q20REYZlcSTwCasMCLVNrQnwAqLBAfmAcQTMW6Ft0eYXf1MXqfB5z4fhdaTpjYbjZX2r
rj/m2Dg2aLp73fq0y+V1ZXsqgoDw81eK7qxMJvn5DLgDzWdKISsAqUDcVyk6nY4etmrdWQcPfK15
9rrBYYRbZC8x3snKU5b+s2oNsnbBsQdDvmJco6z5nSI/GhRllscXamnpdBMf+bYSVSVaYEQlkmYA
CJTM8+O0TLH1Ww4y/ajXIEMito1UCdX5ABpmjP87SMvtBzquAhnymYlrK6G/roVz9M+91wEChtuz
9F166PSFgYqEI2OHeOjhAtzawMs0oAa0iaY+mwZ6bDd5CiD135jRoeDoeUt/toeG5+gbsJszHatq
2VuualUu/SqKo2bvv/dmPpcOzd3GmtdXdIrSB2iQiuICTqdtWWOJ3X1AW3f+vNDNAsYo4vrUMfBn
HPlHKZ2Nlygi6U0UOagktNIWPJOkM+8b6aKUhbRIN/iSQ8ks0EorXRsWZu0xYQNWQr7r73Ww6WR/
e2ZNrqBBb9uvC1sW2sE3hF0egreqjkAQydMkTyyILwnkWsvwIKY4SqXk3Hx+zXQs+txTzpyDiW2V
BXnMzFl6zxwWX1HAt1KXgY6UMpwrRCP1fFnEC8+MWluIQMT8Vf4KQnw+KhV5rA4zHL+nUDW8MWtx
f6k0lIoOrglkky+YBrTQl39M27tuT7dEjfQoCUw0QHbGFCjvr/y4hQ/yVRMH4xQqSQYN16JiypI8
d7x/KH7Mt9CAcjygQaY3XhMY0UFrqasmfVlTiv6ilw00fYrrWtbRPdzB1+eyzHyUOZjPszc1g4K8
sAs5U7Y39qjcu2Nvo8QS7tRHD34rAC7WvX9jsgQY5Ibo2OkP9MpgqkwbGiruWg56srEb6q5kp05T
RarGHD0EgxNqZtQlvrF+jDjQodNi3pR977rwsbaz0H/j/pl2FNKADmj9UZooIA3VDshWw8Oj5orK
lyUbfUR69Bku3zxyFMrYpe2b7+8xezeKhpWC1SCVsNQ+xyiOZyTF2muzXOODU9YryajteMkz71NS
aii0DDT4fc2Pp/JwzZy75Znj9xDYgxz8QIUH2SX3XNthZZkulSTh6jgff+GKXZXtPh8jdErvFQUp
XbaNKknSi/rejij77Rb9GHGFiYS4Vh/WZNczQGBTvZAMspaEc4zb3Y07S260ACCe/jPIMz5H9y6G
hYVa6U9anulz63xUB8fBhjaVRJKi6nf7s7cZDRXFgzx603CmdwksT5JyO4TXRO4OuyS6jp4C8jw8
bn4BQyu++iluQ5JKQtdAf+ho1ImYJRv4Op+5S7sr+no1m/2LAqo28oUBzqtDnUikyG9GY7i2P+YL
KOvbPymBdufkssB7lxTRVmOHLPYjDNKuJqleGOhAz2g/bZLvJXfRxHsCAO+SunElsQE5PnDYXqoU
Ns3Jrcuxy7hmzKAEVTZTDHJW9WMltbV6A2DLEVPeK3YvYR+Cce+IRwGXx15aREWLvaBuR1ILFm55
LNESkpVhhZeqjzyLB5/kt8JFPjhF/7mEFkS1t4qo55OpqK0dV+Tc31F7OZmZRAxwEbixdrlui5wy
IIBEhmh56npUq1g5rd/NLSQZ2i/iPakuN+/clxCm2JrTi40j2v7WadpLTVR2qKUIcljPaxo3o4G+
A4cGoZuTG0O4+VLa0M5A2DmwdjkvbMVtAB4VEiBja9bBwO0oVMwmJK+dlWMWfXJrx+L+hgadafpQ
ypRPYhUDYScXnVaI9IIOclzP80eYw8fraaNYhzQZOn1JvhUzgDHyHBS+zL6N6PsxNs9ynF9s3GrF
hL5PLZqMe2o5UFZkpuBRrRuhLzK9WTy9A6MYTNgnYNipqSk+b0nyYX6gh6ppY98WFqOmP1xfLK5j
RMwgiTO22FswTwlADAlZxaIQZyLZsiTgjuU6IEi+QbkbfsS9yJwwWHkY59KJbV9V1olW/p22XUzH
AaqBh3yFKyNN34iUC0jQ2LzKBBIeUVdpfn4pFn14WWA/PQuhogaoRX+Ww60Ed84NvrsJWMVf0DCU
AWvxUJuyQpnqdo6CClpGZ64RkD3T84+bbvqWts1TGXEu6pEityVyaI3aaH7nUgAX8KvdSj00jre9
pjLbgBsUm/WtZLKk7rAvnpF5P+cBLF0MSPm0IxYH8GaexZbLU0mRX4dt03LW/GBTtOMcEFHHSNqi
Y1zfHOpad+qcBgP6vqtlTPtc4fV72pgKm+Y/PNXfUUwmyWkLxKsapOzQPVYFI/pqxPgtKCH6cCs3
LoTDOtYpOlCmaaQUIjNL1Qt0cZ3jSFf2Qwkbw4nIXwueB1d8yPoazcqG5wwh+mFndBDonpGPwW3I
qoxXOPCXBeRHGEDvOj9GnGoOJ5u/wVn1hpf8A27sRmZOuiLi3/+0z6iqPR5nyseJbkuyizXWilWX
3g+JmjTlGjiqh7KTp7gJRhXIQ/2JWlflOcN+1p1bJv6RyYeNR4sWBaHK46QKrc3h1rR8ck18lChG
zCEkm7l+CNzhIYlr/zWyFonYsuBsXt7bwly6o2YwUuZuTgwpH8aG5jDLd4nQQl5NTPVHp4jH8Xxi
HTezk3Qnf/JZsQTZi2N7KrLKSvCGxc3zbIS+fxOco7xuSr1+mmQtdqSv+gKZy9EaPqHl93hIwC+C
8fBoWuUvrAy9kL24MAFC4tCxfqtUhVmof/IlPckjt5wI9pV9sdxn39WGO2rE4BaA+YBsmhdzDCRu
XF73nX1Z1nMmWWky9srxzaMKjahVjBeuvN/9sqPaOOYg7zac3rlLbq7f+jaoDBdhhwMhBkW6jnw4
lCmczjC//EydjIen0Fdb0Az41iTAT8wibiBuWx5MWuG9Qci4G2t6xQVyPvtLCxUfRO5DLZZqgS11
/u5/zhvQcvaAJVW4Nzh5lMJ3fS/6FFmN6U5+P6J1oG47q1VRE3JMWI6zwBKZk6UUKVn3ab4swXcb
0a3CDHQloHVz01KL5ioPG7Sraqht8pAU76GVjkz9E/bVp6oKfYMYneu/3Wu/MWLK9F/P3THGISGX
iCPlQGJi0R2ECWXvGI3ZAcPHmfnQ+l1gPONUey404rnACeDo56bg4kWTTFySjVYlsbitt2eZlZht
TzA4v8I2YtrPI0uXRuRYFxVrWr2kQ42+xOlMAMemHCDv1hBSn+rmFVK76tXut9gsSe7O66KEqDwc
KzDwqbiOdWyJOcq2ct4kNUdVqy3El5zsRObrLxnexKhzKu3YS6MjEcPP7dvVZCv3IBymwNjjFubW
3npvuu3E7P0FSrmAnKVNKFUbQooexAaWVKcuYpeKQoz/SVvGFwbmSM5t2L+amsNMPfR5ZhfN8S2V
N028Fmz8a0Wrs0eYdJfdMynRnamBSel1DhLWMCIXOrXlokfHlbCmDzBWyOf2s1vQ9yDCIAvOwcXw
7h8q/yDTlZ6cnlVjc+AExUQxckMdC94Q/lMHZB/09Y4nMyHRjzdVo/ZzGXF4NBmKsQqcCI/WPOiw
HfzQJjunqTdo3kcIafJAfnJM67ZbbFn72ZAfmQHoJ8a+YUpH5zgk82yaB9T0736pq/Aqo0cjRB6/
Rvm0lyZvgxcZoFhnvJZ+xxpEy8Mjm19iYTQ9biTygObdnb2DHFN4qba3KNFf8pgs4d9BdwKZl98r
rE9FpePmVCtegUgK8dSW0oEV/Mn172I33ItIIctrRfjRczct1seTm8FGQ5eUQORDJpZtEHxujmvb
PY9JI0j6nnc324Do3vgoIxsP0a9Xu14+jttXejupweaG1oCRsep8LsZMyJTjy47vrfSIBe3tsd4l
FvSlAfNYG2eiukProeQIIOC2WC4wG7Ub5WnZjHuexA2sva28YNLR5G7Q+y4+QcNIJ2eWeV586g1h
g9hZZmhtYn0FCU4w/xhsMcCIOLCyMgFj2ZlTWQpcrDgqX/DveDQ3UjbcBWVVVCO2QisU6o1s7Mje
3u8uVHAh+1Yef3zxIaNsLhXDVryvRUGt5od3Ut3FxrN2I8UV8HBBjaaPC1d5hbg4KPYOTAi9ViRp
7BxTlAj+t1FGOn9uCu0+bP4lg/qU2EkotVafTgS+bM75hMVGyqvh7iExDdtSJn5ymdEvr4HRPyT6
Qn1A5twcbJY1IlKbyGPTBTeR/AUeGq7Dy4LiEzo7+c6FYRc5lNxAoA0wjjXs0m578SkxNH3M3Il8
0AD3a/H0gGlQy84ef0pD6Rn3bobhFgKWaDWZEkdL3EAT42j4jl7Xamu7gZT8VvROwERmAbsWR1wt
wMP2XYHehFfa2RDRiaQ1/yZfMhNKzPdq0TB50w5fQF7xPPDDvt8JkXnX6iQGLY38vishzNh3VBJp
lWXOIkvqX8tluD2jdRq5D0CneFLMSC7y/3lehax2U5ROldkC1m74qzHHiwqFUuN2mHMD9B1daVIA
+INrHfWHTj6oIECRrfaqsrv6ZsuIB/UqyKYk1jxIKI/Xxv7AVD7PPMzdI3yBfvxhBCnrtL24xa4F
EPI9O35E0HYTM9xU5vp3fHvXWqcQ8BRB6otTb0S52ffRgtsx9MPTKglZ1g6pJiPa0jrHzUp/AmbG
2W0ZRktPJg3zxUGcqa631hSynMmQ1NeTUuT0hWXqZ3Ev7/ibQyM7wwIVY6YRyZuBL4CGJHBzAdeC
YnidrKUPIhhsNBrWtMgFsT/nwU1/LldpJ7ag4CgEVxuVtzkIs/sqRWT6uY6zkYvto3jFGUGpYGrY
CmTZq+aZWkkcsqWvRmANfq0RQVfXwKvu6/EDQ8YCFM4+MqvkR3UixKPm58ysTZWGpiFm7naipxhs
06MskKdBtFPm3Dr4k6M+llHTy9lrVLvPMsWuegWel3H69QVra+EDRAuNRTuS/dk9YtjyGpfRrLfo
Gm1GITLg/5yhZz5O4ZBdYuksA/5Svp9pKH6nhuazAghGLHguZ7d8egW+XhQAPrHolcONZvsc43TW
VfPiONMmmtQyksc8R9MC5TabpIB1yw4pu72dHRlqX1QELVAn8XSg8maFC6zc7jq7BqRkQ+7YHl68
pA5SJHl6oq50INDVQYx9CtftRuEkPWyaqDzmeLUfAcWOjYbOfS2YJAaBmi3kqdiPwVTnmTlJELp5
sLfwtBOOPJbNzDGpj6c3HwRdp9g6Na/KV7fnqOI3IP0noqD725Y5xtw6035U6Q1ElDzYyrCZkquM
O3OzZ9NDSkLWVcx3eRLinHQ4k2QCrUIi+hszBT2dNncewULwiAqcDLCoA75PdmDCdJY7azPpqa/9
7NXkl8TQtvjViL+WaCz3WVX4wxD+8qkG87F+Ftyw1cSRKFtfhvYmwvscoJo++SCLBxe+EbjFzWkR
HEV5LjzKfJOrvMTsIw1AIvPIksS35/HmIACW8lOq6iiszGfomCSmE/gsmQCMmIXuztU10u4xaX5n
FO/lx+xg9g3xGN7ETIfJpTEePVtJyHIC4o+mpLc/t7DiP8Negnm2YffjduTVie5qkF61yJrXiqHK
3z8AfvesiPCML4kr34Dp0CK+NRbDfpK2LrGR368lPDnQ5kXdWCaEyZ+PKuMCWKq4SeLqC8wEjSav
HxeduRjRAOdzWfa2mmsXtyM5Q/P/0eNk9tm09BLJL2Kl+PG9NrbdjkK98+N5gyxZ4KSseDB2chBX
+9aikHTQ9R8auyIcQ4vThtx9EScOgr7kF/nijxDIQwG4EXPOYIxIXD2H4kTJBJPVouKrdf1u9DlB
31NOWP/UYvZv6w+GPygtw4FIyYc7BzMkwF2ri3q9IVFpl9t/DJxjJ5KA9bDrzO3CI7ge8A0Dnz3U
6Sj99Y3RxjxELf4iWGk+OhT3RGJmhav7etlQIkuE3rEXaWPwD8nkpGAusUMSrXmQR2yOibRPK3Yq
AW+GzCR0CHQ2xV9JnR1I7qyY0oymU4hb/vZ1IM5WqGzPhBM+HWHAwLdAvjGXhhl11CsorG83jPLW
caYZUkyFsweXTvFxuOR0J7Vzfd65kDnsxWl4Vp6ydBTDXNOdFSWGndWyD6i3aiIVbLXFJBZgH6XE
Gcqm0Ij1aH55ZJu0aauawgXplaAqa6tD+2OwqrP1Tl1nr+pBTB/sHq6UvOUDWSx/wBr0ACECQpZW
hF08hlZEHQWjj+/WDX9/YvFJjmOau/P1F5iNVkXcGfBFfhvHRscn/5Z3k9ISf0+dA8H7gAybX17k
1G+KWn56ziHcglwAPaICcTSXznxe3uAgh7naGAKF7mkYt7+Cv6LcBPGR+I7hIvQHNuMpkeol+zcI
LYpDcuvs5UbAvbyOe4hBa909xqAlIB61MCgNZb1XT6ayMx7MbCpp7R7kW4BwkKvtvr1NorpKvMTj
4I53es/n9Z4o5KosSpQfBHZLQ/j6gW/hMNLI0/r4KhTyMKG76CPHqwMMr0UwO2NyUnVLQc3mzg8W
9mGKvgdpNJxGqDziSHOdIBqZ6c0F3p7gn8OBZaUVp5QriFFagiw9+kzR5bBPPcgyxwAUccISAX7j
VbQzU8QSV5ZjOXATjeY4PzrptP/h9Dq5Ya0++jOnvgU1F3oU/LOx/l4Ari6d7r6fSLzqbekxkdTD
eZwk3rmfzbHrH+2pjida1dUSSJpPPe/Y8a7ptKy+NZZXLkQgO4197nJnydL86FSnPrsf57umvyS6
nxiycXbs5ZBuNIjkXmb71nkJHkefPrcG2VHxugOSCX53sSM9/2vksGoBzucRqv9OgHV7H+13mdIw
BX/Dmurt286JVBk2TQy+ejbwRFygvcwLieCOmoJHxCM7SbektbTzMRgJ+sBvlccaK4UBijb9ovPk
tl3m1QpysAwb9Lm9Wa4uySXiG+TaeS/QER8NkwT1C3FtTY2LjlX18n+dJT3wxFQe/JOkZVV6XE7+
k1CIKitGl2Abe0wo4QIJAYtC/sPycLMGbZGYPaDf4ctOjPVB+IgBeJ5nLUBZehR6NResbuEpkXK2
ofIPiMeeJRCYyalgEWmYkUvdL1EnkEebnLShly9883KW7sCqYH82MSzJJKTLBU/vQSujXajo8Md6
aq/GXz4rb67y/uaHhviR9eWkVydg+igOZ5Qw/wezTn5TbDgXsCU7Hq0vDf88MtdXw59JEFLTNxSy
yHAUw4CL3HE+KUN8CZ/Fs1Xy2vU13Ip0ENEGZVRwDYnoJDVIG9Bb2Y3VpD8YHBfx/uhSNwbIGA1T
lXbCdgmicD161CvNHcfyclrPz62cufXEEL7WLj7JdJb+eTcRyhAHyb+u+J/cWKVlZB0gDCbpyfNL
OUT1Cadh6qAoRF+KFbXfISrRNXn5sgf2In43wzK3d6ReQpknZrVxBJxq30emuztZ3M+eh6Iqg45t
sbPuncyRLfij5KhwnXtV1zBPsjWRAAZpCwgt2q362q4GrGC3bFCc2UdY0ItqtTwl7VeAIplMHUbB
LQTezM5BCmSDTx+nblHE02+inAsEBfhTcpvn32fhJSZwYyi0GW/NLs3oOQ2fytljD7XjNMGwPA3u
SiFSZq9WfOlDHfqq1IX2B3d+hoE3gT8AsA91q0+cYJ7yocGme/C9rKWke6QWyYTV5ltZLVnNqMk5
rELCBeTV0jdPDjFPxvOQaajhF3DoIBRPO9yvTRnUEcv35a6foXQFHxr7BeatfLHYVCdPVORDcsiP
ZCfuKp61HQfeTBKNwO/yj6s5H3AZPcNZp8OgBOLchiEDZHqbF+QAoF1h/eEVc31KR0IAE+HE/aGg
+Pea0GBHbqdpAbGgGOq9YZaajBchyhVoRKib6aUprn08PZ0IJbL6vbHJsMu6kHvbVjJQOejazjqj
xo/Ry3Y7OBa+8aYNzE65b3ylBbmnyvGYUFVBYC8dbOfFJVFuw3ZNlil8inA8HQyKDuGSAlharH3D
NHaLaVoxxOE2zEVrdlm/Gbr/Rsp9VUXFhJYn+WVh/4mwksde03wJZR0iaYjXOmb6DYeLg0YSRcLj
O8wCsvDS/uzoRE3nd/nbD/UEKZfXaP4fZv7nAb+Jx0aOYx0SUNz+ZbIaCWpGl9F6E+1Ss1Pu4w2n
iLpLUqOxQVRWdOQvPk+JwgrfcQhqW9H6NgAQdJ8kkSG27ZLCyBwgBiCriKTWl6eLNlQi0wU1Uj0y
eWvNcnYUgt6yck9kX/YMoNe4REO4bCUUwipBH/pjk81SSP2GUU4mRk388XlKCPltDpbGH/4KZ7a1
HIdzH4c9P+hpHjrDYjbUapk1s6gqILXbw1cqqUuWN4SI3+6fCQjt4e/iXo4f7ksA987S8kfqz/Wy
GHey04J6TxgrQFTEnVqMHR5NFndJB3mif93/PB/gIWySa84MqQ37WpPGuPxrTSoOEtwfXP8tt9Vt
vCJAG/hoh7fqXyDAwkiNjpEsTSjYdy16fY7wTtwAupJjoJZjMawZmoi6HSTWmn0VGHGlAebfPjJK
wMOiGn+sV/zxiTbN++MTfGdVWZEcehVOrJEBO2C6YSyXVY6+/gYXjQA79oB38nmldnpXOTaWPMK9
peweQXVuFj4dhMPR5DO7B1dkpIQSGTz4o8Je4ndd8Z9qW7F/ZT2XUTqn3ljSnoFdDSYtMMcYlc68
newgpWC2vfRjjBqt+Hua7BIcWvg9LG2RPw/Lsc+Jt0H4q1mLQXre1HJ0r1RHTnMtZ5a53QgfbOTB
XuGwIPvLY86FvcpRZKNVimbnxh3oy18Gout6N+InPO/hXc25V6R3RBOZSgFjOMC6d+kR0EyyiiIw
wgGgh7Q6eG+GUda/N6sde7De2xNAyoOJCiI8SFDgHskaecOEPsSW+Owc9ssxaXH4L4YJsxFvRbLG
4c1PtpLLyiMM+1AxHRDB056X2OVmKt47ZYT9s+u/tYs4f3Ld9dr1H35Z/dX3eMEuWm1USYfmi16S
VaWt68fsfCgd73loNZfpRXRf60d1sAWtB98m1zTD8KQC/YKogDC++C2UwlDjDARALj/ezsphrnjv
kuwmG0FWRF+ogMD5iH+OuQYgMpafOUOANSmotcxExTQPCT6xaZ80fEEG1KuOFDEe2f3U6Wfgp8c6
QeMZFdsU5ogLkL9E9nOu9lqaOGTW0A1P1n4m7uH999yKYQr7V4KgZnMosOs/NkM4B5RTpdgu4YrD
G1axyqcQ6/vfKz/vke4A1IAKaT+qYv+C46ELeET7TvxthN96xesAhnEgAatvfuyhJ7CDC3YfvDnh
0zzLzfJJhPCdwcswAyOWVind0Sekumv+3FCfvcMQ0ZlufzO3M4Y+yUxzVDCTfJWMNv8/TjUSoI6U
H+g6CLGobA3AokprA3gE38IQFIO1ZfghRcF5nBoUgq7TVxY1wIynodFU4/Roa4T0CJJaFV3HZRH9
4BNMcyu4xEQiUEtPW1fXhFuh1iil4/Y+7pbo3rg+Y9Mpr7I1R2x4QMFyrAgbInT6ZmwxyLD4LzOS
uSsE7A7fFi0mvrZirb/3cRuYJ7Hp9S9ACE7NcHbr1tLREa/IioK6JI78eJCWoBuy0kKteWhV7IGw
XtbOMzElAonM6Z7Nu7/H8qT3ugWX+/dg6NX6r0LWLyEVoq2c1YlzX3zBUS1sYZk57AORo7VHuZ8+
VIxQ5DWMBGiBaCG6uhI1SEKdA5i/8x4rvlI+ZuKado8dK06KCP1XvX9P5XPfFlX/kVEuE5jmjJ/s
lPA4KDG4xACzWRU35hHZ7Dm8rYQY7rsT4FZLPHUiY3d/QozY9azTx0Sy7vq8xntSBnoSmmPUMctl
T68unWPvok7Hei2Z7ng21DF/lzvD41ZM9NQx3iX7Bf0Fpl71oRxKLmSWkMCMHIfol7v8Zee381PD
c2AKGdDcnCNC8DWTCxnCQiazumntZOo2aMyq+YZAjMs9zbpbXTuJkMXqGC/S8+m316RYc5cwo7NA
bTxN9DM+v4AyKmsEtoCoDG5RVauNqjv7R0nmjPYgW89uoX9Du3pUABlymjNiMZnVhEC00hNMELF5
/m2P4K64uKTEbIirve4FiMAm3tDb8LvFgPtSHN+MiI6L1nKkJy3NpQZf8WGHrZIMpw6laIeh95Vm
04D+nMFyYoOPtKZYgSJ60Mr947jpaZj5Vvraz8X31dX2p8pmBPLjYlsPRsKAX5s8iF9ZrsRQK1uU
kqa8CaWs+oCoVB8mHMUUid4+BezKfYq4hbPfKLWDs9kssMsHj7KtUtWTLxufUqTLPUyih0I/MSJw
lDuwYr0kG1gtEDkjuG5ZKOuqhiDtFmhpjMfzBSjUUfjlzTk2Q0lEsczGrTIDJJmIn3wahQBE/FqS
XSfyKoGrGi0aTEZZ9qfKf1AxUBhqzFLAQhRYDWWqnTUBELgrRgpOUYiqErfF0RKCTrMuP+9CSU6P
eM3ZO+Rp2bRrXOzdU7K7WE8Rsexebqtn/TY09TLRIt3/ZsnkuQvTAvVRhZsBon5bw/LMviIr5W03
Lj/34O1XKMuitYPpewaVcStsNQ49GKspbKbkVeXZBAmehNcR6BBRIbIfNg+oo95pY+PGchyNxCRB
u+soNWZ+0cwqhjkktaIPe4YfDUinDu/SkEpNem4PjUw7SrzpqMYvcLOJJAWu/6a5nfVFZliBxaIL
98MBNYpd3zCvIu1q9LWLyxNBGPpyMzMFV5kDsQvRCVs7StfO4YK3k5C5kbZKDtP0djy5qO8Jf1rl
2DK7FsZ8zBDG2HfpDMX4bFM2uqKkVEooqN8tBo9veXxx9Dtvjyqpb4zzJudmqJaACwMo0OoJXWek
bmzeYjXfptiCRW/d2BsDjLBBT6id4MrE8+aFBQCEqdcdGPs/ZE4NCNIB3jqiklMn26LgTrqChPZR
83yZpoy7d9H+n0IWl+BNwCUdQQRBsqYwLJnUIQqGuJjuMHW9fZK8vVD9h7a40ScVFBPlZIK4urFk
hhjnAtGwiTvqPMni04faYsiOdEvRHhbNJ86Uvc4yho7mJ3buvCRzM9++yd+J5u1BC/QANkh+N/RC
uzfQi5RL3Pi9rQVFPSMDtaa0yw830LjPqYYzKgX6iEeOP8BIkBAS0ORzrNuWeBp/xTKMy4FDu3u2
zCvBr2l6j1ubEUbI4wlDABX5zGaWTb4qzh23cT7Lvj508/elIl6NYK+7H2PIZH2ciYJ8quMXTwqS
W80vyvsrPJ0AMe9/lBrDL+cHQBWrW19Tlu7lg+q758uwNGA0Sar6kpQ0x+77Q21n+7iCqXP9JyRD
jdCHOxlQ4wASCplb2UDGIxlHVJP7VSUJ2MxRJBTQIOTFQ1p5uMWdqXiJ4CKh5VyEmKckP+NHNGyF
osm95/TEntLQjh/oe2d98WURiNd8CiYM29TPzTLztVD5GEl5tJUtyRviqwFLoBsUp6d0nvjwjAfQ
Zjp69hEoXINN6bLwFMzF+vIeuiOfqQJ23ZMValYaTUMcE0nxkwxTjFvCMZ9ZP48wcXDJrT2h2C/1
bR7JGHdxun3BuYvar2X4v65+jzXXphTGwDf0RmEcEVq3DAbJhKS74s++InoRNwbo5Eb3NykQxhiy
rnaelLC5uAV3DrRAvVDXTK8D8XLC0KtJd3XmMvHXPfazP0KJ34Q2dHcQsF5Yq6rGukGYdIJlK/uJ
TDhoY1Ub0rZ5G5hxY6bwM1xI47Wp4VS1CFnRHm1Z0Afyde5w6zeage9ZeUN6gjJvK9Z8kxNhov+a
XnFujVTecQKFV56CGYrfVDAZpKUdMEEc1Q5pO69yaaeOLNgIFYDeRaXNPRjxDy+q9s8UGoWepidP
R2MJ3y7dHtVAPbLWVFd6rj56Iq453uuSImfECIHyDByfnpCXFgSYxgkBMpVdhnzPxTPhr+gnV8bP
vh5GwGT1woqHj5wdgUHt0QEQykvT6aw7YzMcO5toIqDls7X18DvYowOZxBodL8Awbw+BkvOgFqVM
RM4ajUEUkiFDN/2zunqpWxmZo5JQa1+SgHuuhDL6XUV4F2K1TpGlkCsJ/AX/yoh8paXmTVAg+q//
HMss5vHTFe8NsRRQGUfd+Pa15oyni26fX+RE90VjVtCi1z1qoI5Sjudl6AUixgXoEu6sbxv8MnAQ
mEvTAlJd6DPq3IpB2TGnRkb7u+6aVT7n5svSlt32lUUwWpKKQYKRB3epTieEzreitLZjsZAPsJri
S0ut7+ul0HLXWCwtQMagB49O2Vu0R3VWwtxdCrDLtdbdM6dIbfaZhf+sbm56vTAVrI3k/ips67yT
pHAiTrCTLXnmAsN/MaVid7sEaGlynwKYsH65kr/U9Cqdj+L1yfpyQi0uKggN/EJBTKJU6PRdE7Q/
okarYNQarVcpbdOjscf5gA2zTrEK4T2x0Chuk6DXcgj3/Fbt2E01+WKOxvSNlM+58rjczfKlpODZ
EiLQKDCjdNPQASrbpx3UupL/ehvFp2BBrDoMNoSCu6R1HMuS6B3/ELxSfSJYj3798A+6JKJNDNDH
kV+RtaJ/bk6/utHtUKQw7Oh0zWCvZ8TrNuuSlzHe51LngdXtbVJRJMr0prvVs8ggIveyq6tiaYQ3
n4ujbQeKgUGEcDb4iO6QfvCK39+BqWszxKpooElUkJhyhN4PdsBdfF8+BJQgIhYNTHQfahEMZv9f
M90ZrVQhcvm4ZDKTAssiJL8wAHLkOEhXtxHNH7PdwY8/qjIBTy+PJ9tiVNnM4dnv8fZQ8IlAK8RV
79jXUwbth4HRMs7o+6zGTuIIJ+3xIbMIJvoXNz9ZuswAep6D/Zqz0/urEORnqe3lbteUXxTt9sK8
mOftRKkiq9/Nh+4z2djee0sQkLDvIk0T7JE3OhxUoNWXYq6iEJwjUH0p4a1+rWbjkdx+EKVFN5HJ
4XGK8BcYuxebgpbIzSG2/eAb688UDNaToWyRkvOedzluHeRQ+PQiCelgDGXV7XhyDdid9eaLMtHb
+c8rIOxTJozDsy4xKX+p1K7yd7d2slHfdufMRkAQinMgaYn2BK6AA1JngqVbdOG+NGye4EzQuFgl
wfx9xa1yLFeGpYqDBk64cZSFicWFxppbuPGhRmJ67Y0V5pEFQ4FwVYB2XOM6ZsDUhoOjb9wigs11
fg6HWazRP3uBbrjqNbE4RoZqsntGW8924o5RUd5d+35I9FKBhqWc3+yobfXcxV/yGOJAk42JPXS6
jYNprh2NS15EnuX99EICFwVAYD01kfwYQREP5V5VQHmkThwmtzOfiVHD7395F3B3qmfyM8PH/gMF
BfIbSccQsApedoYcoBoZycA6OcPoS2VrTHuZ2Vpx1Odu4H+PUBmo+ttlToMGeqw1Y0eMODF86yXz
gkEibPOZiUxB+9uYAGrJ4FzFWakvSAMiQ3h9oPtK08DO8NHIhVzrGsBpgQ1FVihxHUQX++psfJ16
uZd/0iaPzXed7zzro6m7Wd9bF/DE0+AlBgyp5svfMp1ilcW5PYejLUdnIp7u2r1Uu3FwPsTLOxEP
lFXzYGYCB7kJEb1Fh7VyS+8ytffkRJOJ8WT7qVUnswhEnPRLyp9GgeT9qmbD1zkdzzCGMS6rCmg9
J7eaNIVnu/NUUT8GphWP/FKR+TaUWaFMX/GggUBCzEVwwxP36BGsuawS49VCMu3jFqaOtmuNzYUM
xpbG5qTxzvP+LiBAzMmj6tgDk2BLm0vS8p1g18Z+NHIbvnGgio66yH6HmN1albALziBiXLFJsoPI
IrAqtTsK8+negR2yS3LX5mPldZ2qxl4yVh2kzD1eoQ7Pb3+HJx7ssSlUyBroLka7HO5slrH7Duse
kfNJRY8FKoAotcnWSEhf2GVw5otKBN2HBBLNFuFFQerhiKS1m/J8n4yRMR3IdLIbOEPeVlXnYwJu
eKHprKJKsJReozX/9xBln3mYig0Ny/Fp9Pb4dMp5jdkl+ZGLCLr3p1xmmAY42sOwlZ8hNyn3fCKq
E3rym1vQ0nbKffr2DYhcjU+ZPkTEd5cxnupWn6sktZAoLldR1w8UBDOdDC5q5dmpcXl1guDkXks+
YJgUyo5Tw/Y968TiYyXJYbQwEYad8lHbSBxbQ8kS/kSC2A6Gas6yhLzRXaZvsyi2J0DFAcxcwJJC
EczGQX2STL85kYhRqktZeU2ucw/HNT95OOBuNnJQvHWuYFLub5xgIFw8LBAaEA49SqC16MvanUFD
iboOt7Jn4EsQNYZ0Ae621s1gMnPtVz3G9PdINizPobq9v2teOelLzPCt5OKS9e2YD0jH8IDoJJTT
0NEN0dIFS2TT17+Ip6wCocN1bnEQmC30NDRy6hIo52je995Suu9iSODl5tIIeF017pEkx2p2Jipl
v1VybTzcZSPTLmGb0FGfg+dxXBi0OhytEYAT4phtUMK38ymfHWN3+R+SscrBH7iCjM+daHki7T4v
2fo3QgTdryeTF0WolfcEkpoKz0mpexgN7b/eIxrVmSIJk9ZzEUKknKHKciGXc73BdynMSARtCXJq
UjGmvlkje2QIqbQMlxXlcEI/J8P8IXSkHdcHtEjYQR8MPr+6j+I8hZoOsspr3FacHS+yTEnxBi4n
5TnTvUTZT3weSDwfsHLSsHS7Aa7v/lwPPsXNqbEfRLMI33e/ug7OLG6+818x8eZVshAn4xs+9O9H
BsbVQlwniCNgu5nftCW+I7tzQDkV4yrSNGJPKrEeQKf72IjU3h53Hqa+nozGaZnJrJtigZuPT97y
A8EeP+TsnUXgFYXJkWCDCLJ6Q7ayB6pHihqq2bsZHs7jkspyhyilmGAyAk1KiGVKQrRDLLb4grUC
FO9ttD3au0Bef1wTXsfxO5Rc5qp7DZMnxqaZ1AYc7IiEPlcoyjwuRrpOKD0rlzjxfQQvsOt3sqAL
EHNAHEAJlMs/m/rwjGKDz4CeDWv1d0T+UjFI6jMKvidY3H8sFDxvD4t+SspYHrlIpzWWqC9/0FX4
Rf11gsEtt9Pz5TijCbyWbjTPVa3ohSfPaKIhv3j5AFMIBCsCAvu64Ufa62zxmirPqQHUdFS3brFS
mEFjnqFOypJiKzBv3Zxk1lXTuvSFytogZ9vg8rYs6j6bUT3M35Swcp1vYbNflBiPge90ROu8WKlV
EfYDaLp0B8WFH/T6H5OngK7/xhtr8urO7BMvofw808r+Oo+ifxxGE4Tx3KZPt30Sasq0z+jixkgx
p2pVjRgAYXPfRoCUHt3s6vmCYFHcMF7usjGiV8cwBbDCEcGaQjPMIr60J6WKb5qGQcoYjqwfBIOY
QZR6qwGFhprCvQq8vsIR+41VPRUugwd+UG2cz+SXR7xT9SUcDl7+GWK4rubvz2MkAfj5kg8aSCib
b25DFZnYkM7gZ3S1tWMjwemtu9ZOXGzg5coA9NMccVHAoFKiKKyBzIW0MKE/pooAO+9Xre1vnBnI
xnGUTllxdfzvEnP0/kI50as1+X9B5CbGS8Cz1F4l98aGER64AOf1u9PsIFTCiG6odWvfXcOZLdAJ
2XgTLXmbC+pc7E78LrCknNS98nTisHbjhd5a+74aUP/2bT1lXNchbijd2eFir10nfDR68dJh4GgG
+LTJ8RzpCX/O0/XvOtxUmGlztsRFbeveL9fWhOS24f9jTzKqPMB6odTvX+t86Y7wwySnOYt9qx/k
gwm0ho2fRa1aEZlVZ9Dksx8ger6Ld5mAFWjDU38ZofLuykPESKIh9Q5OMBqGJ6sXfrJ9uV8CUpKL
IZChaM6TbkPnmzGUOiWwNHrC8omuzjsrQ4yabCjSiMx3uSXg4Budm08a0tprFkkPbr7PKUtygPiu
Ytu60nYq795SaMphxg2aXkVDoxj1n/yciNl2Wfw4j6XUWgTBcpB+35tZ1X06AjYtm2gRXctEghLR
9wrzO4u4vS6SaAEp3I+ZiJHchK2WFnoSzj1Ccm6Rl97OhGfNLRyNZ7+5M7oHZdVWFz5abQNzXoR9
WC5w/Tg94mf6o28WPnCStDiu5ePlsbSX32fRKwIECTbC508p0+JMB5ivsgBiuhl5KvTkvL0yOpY9
6seThTYU+4vgQ+wKiZEQR2PXJXhQGxBEjiA/WorD6qamZSCG0lQTylpRKcpvRrpA4jNPUpMHmChG
qHKY1x6J8NZftEW55HefaT1h76ajYa8ic7WHbhUgNyhjiUAWKK3onAC1uZfvVR4o/cD4sEbgX+sx
euKVsKEDgQ5bGuEGhcGGkwWnhf/yOJxxp2PC5xr2KcWviCoeiid4et44HMw6vdMyBSuaOFYnntni
Bb+ktQEWgSQs6UkVRI8JcQ1gd+x01aKamW2WCZtgMpQtWz8KEbkxKQ3S6PHnGsgK/LbEGsr8qX39
R9f/hcm7sbRryK1tnH20R+5Xy4UXt0A38LvLdLxenaC2jOT+zo0sac7wu5BZdO8arzA0OU3nXstP
dHW/7ofaGpC7BpxUBPKVKZGEGOorTdyXunjKPB4JoVPCf8hou0jrOZBx6ynif1Ha5VuVAq1eV/J0
Y5LdXbLG0yA+mfdRdZnQybD21zYIg91n+QT0hZfELtj0UaLfuvBxIfKW/QgnSzhIHjsx7umOUrQk
T7YngXlMX1gFPlRjdPyrTbJarZ2DGSDb3Ng4gH1b0OzA9OEjxZkUyzhcJKzTWzrmtU3q8egqWBZO
KrKbRmw22K2wUIw80bVR46HjuMw2EQonwgwxFj5oUHnsQY+3/6GTsYpoN3sLaKGEl01p0QESr3BZ
oXcSP5ZRANcN5Ebe+3Nb338PBiNUxKsbV8D9H+94j0APkNL0Et+s3dj6R8ijhzTwFOJrwAWrF/ZF
V5sYqf4pUluFiQlOkxtbRw1afedU+IQXGy1PpvJ2qWitus5neNKNtCnKV0+vOdYBbjyfPZDnjV7w
Y7suMPjehvYPNKGD7oBznBjUVtWx5rvTlqm1Wr3jY3FcAxPbSjsUBnTcQuR7vrPqOxSkIR1ste/h
5recsx5QUZQDZNtFpshznYbkaFu7s8kxEp2AAC4yRfLvogbCTflrNNbHawOEEJOvMOcNXdnmw18l
24pYl96Qh8MwWenPHzTrW/Ecovph0zZcrFvKH7nLG/cC3u0xScurckYZ8ETTPbDTEM73oOdiZAxv
kuW/Pkq+GrM5BFGjn6HEv1nzQL8z9vjlnk1L/wYT/o4sM/om+JxzbAbw61Up9mf8l+iSxX0KnLc3
YUoTxro2ZM89qj8YDD0lbo/f4oLBbkkwuW+ciSoEDaYZsnaA2D/Oln9F6j5MPemmJW1k3rtl9TZt
19eInbyLFfRWCWD0VGnXeu9fjcEHkfCgmnbdihC/QiS+/S4LcZWMzGSpI0Ivz6UhUgHAOsHo0bp2
jjFwmMTYAbfXQtQA5J0+QILbdM+LoXd3hWEdj/ntcAxp1BDrQvKfYoXU4sDmxKsKOWZ+jXQmv0D+
WOrwH4kCnPxRRcsYb3cTF3ndoXt6RwPyD/x5EKKRGrEQepBlX+96EUzaABqFW2UpZr6zz7NeYiMK
dC/zIld3YK3phdGhFQJCmJcv558Qq5wqi1VT2M6FU6W0k6GhmfBwEGGo2XmxqwMOHOhxSSoj5k1f
BphPJ5Gh7Dvy2MzO9ZtGocginik6tFd8vPl4ICSR7Hr4E7E1fy9nvnMPT4B5DE6EljgKGTgFj1Mq
KvxT0Blrq1VBYm3VH1wh9PfoYL1E1DO4YRavzuSmw9nLzHHwpF92e7FeWlsGK6+SfecyP1RHFMHK
0cGiNdmgQE5c8ruexdraSGT9gutVvWqwlA5jXzKEgNVLSJcuoumYaQgSD3eH259G+QOxhFc3gBPH
bG58eITXkeEHKFNh3eWWZooRdkZ/Jn9CBjJCd3Ptj3c18sAcUIMxeCOHhSlwFHg0wy9sNCkwZpuT
a985379WhxUfQxxaNdwzwSoFYHYsS7mIgwYGJLCDnv55ugARzNP/Qq+SE6j/okslCCjgBvvVOSQL
lahHxvj9HA8rSYPg1+fE8kvmDPocEXHO+7RzQjdzZfsB3YyoLPSbF/OZQv0zoDyytHDdGzKvVGQy
oIwN23G1hA6G7kneUP9fznU0ukDrVeaNkW2kkW7Y+jt/PmjYAvJ6SPEjULZ9QG9R0meHrhhj61as
LxQLvb0UYhdDpHm1jnmvnfFUHJl6UQbF6BTMJSNQhzMSv2FvyILRJJ1or5unt0tzvkUumEYfMCi9
jkWFNg3sHmW7kVpLBPxZBTK+xPH6FZPZkGforQrwxlKjgbecshVKx14CqFpaKtmMrs/oTrliHcfl
KJXKWDAr+x5+Xz5VzlpEWCa6sv5Wkt4zHrY0vxXATgRlu04ffAfPnUiqT4C+hFzzECOnhGCrk93X
zSPoZ5LTHLhDDUdxLpYyP6+Znk091bPv7HwQzAq5mL3Q0X7jNM/KRClfQj/ajinw3Ty277yC9aub
+yTyyN9V1LVn9xkfuUhrhDx0lZsTtF9H1JmHoENeV0COkwMskyA9og8EajctQyz7msEemlH03B5R
5UfTZ9+NmkAij2ohLQhFYcX/fXTn2cX+su7aUzeu+6xQMmm6wqD0ATnINM7VR3iQIoFyX21J7ilM
n9qIZklwMIGYqYgRZjivgZkwqyIzfj0s45btH5Qtjl3Jwi7ELBT/pO4dlz7KudnwTTc13OBjeTt2
jE6wpQS7TAM6BDvDoMOyVeO6C0AXFJ2yBHmRfjVMk2M4V43uoZDRpLsxqiuaD68QdSQsBec4xIc7
UVyZ+xJ67hG2XMQS4B1HAogBN6mEA7SGBp2fs8UIcU5p5dsIA5vK8FIp2bSC3q4X4FY5ujcXc9dq
GjUiNcd5A0O9qzBhAmO9G0NygGkyQFJSZLzXWtsXu9XT9MUyKwSj06o9reawtJ6Bp6H3XWuOWkzi
4I627ad3ut3knWFJNhCbhSrOPzcOJ4rMw4iQ/DeW7E/Az98JJ3UAjsyE11N9tlBLexv6yX+Uv5Bo
i/fZhn6O5NJnI22SAseemi5hCH25wNwqLcgdEXXnCuDz+HOZg+SYIYjHKYW4aTPFsFGR1zMFwf61
biMFdNL+3WrEHivzV9PItMDqZnCVg4NMqND8va2A/VPz2s2IO3NCWYoDUj/DyLHaLxYrwoYeoqgQ
hxO9eChsQEM15CrLBcijrkhm8ymWJ80wPYRWZvdUBfg1XKszVz1csX5WsdNUHQO5PJ2fc9mkTJN6
djlFF6FVv93CbbJ1Dc9UvMSMbIWn1yMnshDSmn3q6q/7k+cs2x58hNun9nMdWFsa7o81k5vz+RxC
2AJA5SydzIMJf1PLegzXo08lqalJJ/D4Tkc2HMSUJPNXiVihWTde/l7zXimMwUoq76Ej3VK+6gkk
f+jKXPdkBIRyb5u4TpEDgJNwPwC+ndqaYyr4VY5K8zrG6OFZGIb5MlbeYRbbk/6zpejjwrbDquHB
ThoZCLUzaen3/5OSdf/dUboz8jOUSkzWJmPSwKMsrIWFe1foANgEcs54rEMdo2Lqd9TMsmycAzzr
vi6OWrkyu9Eh+GaN274ZGpvH3A1yLJUS3OYucXZZuYdmdcPmFnbGzBGnKhxhDPLSmh+ujp7CB3Yk
DKPlGBQcHqxNvgl+/s8x/LnWN1fBYWlrm/64PAQGXc86UBHnFvcpGBlwHuP0Fv37XW/Y6zNTrOuH
+U1ctEwgehV9gB/kNQxp1vJdIibFnwYaqUNe1P70OIknrVMnFY0XHY9TiN/gwqw09KLwZnTP6xPw
2XL5RkM1Y3swhlqKjMSniIKUarGRbNXgXzTX5QboXzS3mR32A8ShKm3oV93gPRYSX+URG20Ywetz
TtqRfDMZ6I/hxEL/z7pswgoaJJRupTIeAv07ohf49NL2DYC4C/gf8rV9JJoPODrygf3oo6T7ZGg4
3Hc7RVK0AWKs4qPSLb5lusVr34Lus8Aza2Mgkm3DTEi9q4+lJ66/cGODibfArC8cctiz9VzuuBzU
ntwPy3/1n8YijWeHBdbPzJOKX8vUR8nAI4gIPmdqhgkwonNFAIIkOuoR3PAvk3W/ASu8UMVLolj/
36uUBh6HmsIUtVpgTKS/cG6xEARyIvri9ksF8Yo1MT1Zy1sQhC3QDSNkFnZFd0VDtddqZZQ24RE7
gpbJMmpwpwfIEhJrYHGMooceNP6qg+QUaXRxXUg1hJubAE8oCe9IZwjvEUjmUkqgs4a5SaMputU7
tPB7/BOxsPTIYxdGI9/b3rp97SQ2CwsANLcymPUxPkbXqwhMicG+HhGYaS/aKAWa2iNP8AJok+jQ
LAtufzv2VEPvAcDGejE5Knr7biaiw26QVJSPr5yv8iQ87AoT72Oyj3i/oKYHAOaz8ofSB8XcsK+X
6BmqF8y+7/m8AcGRVhpL42f0sZ+kyH5YNb1is9VTS2ItZPHxI37rIzSSppiitsdVZkP90d/vansW
q8GpkX7bucvGSIOaVta+clo/AF3DdbD4WRNE9P7kXckLAxcIX/yQWdoyTdrS58TmLXsylVwchtFi
u2LMfJG6YZPAnZ+DCFZ9DEDmhEdf29vg1wTryrQqwbDMAzm4/I3UNJQB/1dgdYW9r4h6rKgsO4C9
U7JOXQ9lU7asoliMJtSgdEs+CSDze9r2r0eeQiEx0wuoHuMgY2vrtvjDYaA5HlTGApFtnLZ3q47o
3nigueEVsaQQKBJKv32DBErUPfb5ZxBVdSFzwxkTuv+YTx2Vr2Il8mYaxxQvdV9CHDP68HHo9ObA
1TQKHTh5Ch3AKFxdKbqA2amKziuS7Fv65LYl/dp5Q4GAeMVRizdpPXf/eV7udn5VD3TGPPExZpYc
tsyejRyEWEENDfBnzQQCnA+0Hml4pL9IX6IO/0tmwt6vKUPIdz3C4jahz3tChaGH0ebrxf6avCIh
VjybCfmqo048RFQ7rB+T+iIx6lczFh9XoJaA6/VLDrbM544apqgPD3eGjd613zwyMyzOxSszLOmA
4VE6LTSMqLxFh88Gm3Cn/QRhOtwG9IXBJ/qW8wq6Wy+/mxJDEuo44phI4aOaF4gYanbW+vi3ylq3
ACIAa0ZdEdaLt5BSGw72+RX0hoW34YIBj6tPznbyXN5piVgxIw/7UrL0fyPu3hfLo+RNGkFnKfpB
C3D8Kf6tokaoGP6OKpSB2uM4d6suCtP9TTz42hKtpIe0SrKCwhRfYIgYFT9GBrW5RgEHPdx9Xp3O
NL4/qJYRzvrPP1D36FU5q0xQvaCC/g+YbkLaBs9Y/IGECToyf3bILzSWzCPQhGSXPPqwM0GDBWx0
kycGUKhBZIiuwHAy9IiBQVSIEYRwwumfxn2LE/tsXvknISVKU31YcuSnSgPoGymI9ece7/GsoPOC
Qsnf1vIi5+ukcVRUdMEIfI2EtgrkonXLz0Org6apf60Z9Nz+fMuLJcRUkNgQHrWL9y0VZ42dkOjw
IvEhNbiEYi4pla9SvjQHW3/zn0/jQ/uXTYWYeyB4ULE7fms7T9BcZSbxQ/o2suMP5dEcfihaocTO
Q9r3wlmVlyCZq47FYoPMBsFalZVVDDZNQV54n+Ohu6OYdyr7nRTU/V22rLFAGLyYGb7Fk2cbkaHl
1DkX9S+UWPvlZKYSBSvxbc57BiuzIiBtpqeoFGKAehG1DShfhgpUeuuLZY6AvZ8Lus0BgRIEYThu
nKcki5hSzh0E1cVMS5u5M79IbxVj61dCGlG0lOZMS8uv7E03jTeUkbqifEmXguVbUwwqxj4ZAirK
Um73ViSDyPcLxj/iL4qdaAiK4rCc0ANa6QpcE1X3dGBJnhaGfOiPOBQUlCdIN6rBh5yev61ZA61V
dfYvP2Q26FwnidnZ/RCNzer9SKiRZoFT3xJGMC5NDTkIF1UeNlU2WnriRvUxCtOpxjEgslN+WaKc
Y7wk1lQzFcgY70fa51BDc7gIkvrIJSd03fwvyFfm8QaRKE+V0gfm28WXRqbfIlTJNvVUoAEdXfqi
Neeg5I4lQWhntklAsFfZXXT6tOda3PzmoCI1aa7So9hhXJ13wSkZplSKr/1vUHIcY87ryo3482Fh
aIhujsPgD9DwDshE3se5cw2hO6B5Qzi7Q2NxR+joLx5rO08BfVnZJjjdQXixpn7TU+wNWEB6rHFc
1kee1OFIXHRTMGrxgPtCwIp5LkurkUYJjQEvwkeElaRRkp0K8rhaxQ5a/7RnwIMAQB4A5LhOtvkW
p51s3OPDpBDc9+XPSyZT6UK5ATBgx1RpWV3BxzMcLP1nv8OI8zztDL0chHdDNZJTs1v2OVFkp/de
HRnqftLd7QY/W7Quj6ILGMQedlh2juEX3LZZQ/WHSlguaqK3WaX/PQtvDFXUNL/4baxJS12lz8WA
Vkjn0ynElQUZHPUcWmARYBzgvN0/a2zT/U7nRYXBuo/TRlJbY+Oum6vwwPgzHql33o/y9Ju3S0a+
8uitdj44OKqeUFERjspjbFcP7evzja9L5WvUMe61G7DVSlaJNfodkE9mbvVgI5qEjiOdY6Dt/His
VkSo+9DhI4TnSQkSOONDDCIvUrmIwwpJg3mTkyAFz7e2mtDneVRm7KSwLOchdeQg1nZxqhgU+BdZ
zX3PIfnmww+a3TaJLZNeUo/HiiTFlFHH++da7pP9RBh//l/dPp1yYpTKxf1pZtn85hBCiFQyMdLz
7SCPCoDyTy4K8Q6cqYicDe0nsaeQda/6Ej+JKlIASQCyVgryExuJECnaNR+PFUhiUNGNnyJZJrfL
6VW/MqGhrGASYrKQ5D+ecDTLsWF6qPHnfczhz5QSQ++nWEa3Qc0EI6szxP4pNwJR3gYyIvscn2cu
VZlGUl4yhjLDX6LZnptBdc0reRyP+UqXSW965lXvKAnjvswYOOcONkS3nGWZtzcuYXD5UITfeuD2
+J80UtfreV1zqAkHd1CCpBQ2fVX11cx6pxnFNP7y7KHajGQXZrjABRmDzwP+3pjm2jQ2iZLy7VRs
n+t9jzp9K8Y5fOgnL82SW5Lk/25HPHcI5K1w9g5y3hkJhS5l9yz09NJVtgHdL3FK7iMuN7CslJBV
pNz5VprPr8vSeDrlNiWhqJBbWDtl13VYsVEpelzrtHr8gm1wVQPFIDbYtqhaP4xfW6DfA1QedCQ/
Ty/mloOzFxjyDbxhUfaYfioPhprXqhP7XNBl4zf8uFwiWnPio9pvfQXb7OA7TQnoZMaAliVHR8pW
Wp/SIt7zO6blWPRBFelboMv8vNovh0KJWvaXCXCF0aghLBVMylyzBUL2nK0dM/PtJ8abhYK5LkCZ
l3ZhmTzI+VGYglcGmgxJFUkp/6JcvenEx+PH+guQjWzStoZ87n6taHFrNm5Y1mEU3ZKNkiI5eiTG
owTgqNThSmHl3+0v+NC7AAI0z+W6sgg7vuwTj7BtT5DL3BQMmQdYhhHbBEkr+Vej3p+IYtx2XDGP
FynVi/VQquKDrF5LOrb3/oESlR7XxxOsaJwFWFjqT+VlUIrQR1jJQPOApY4LLdIsVnMr4TDp5eBJ
eW+JulR2TF/GgkI/r0cb2F92teETZ8SdJSzYNy29Mq9Oa39L9La5eBJmtT5uHKsAtgDiMxA965ix
qdYI5uJtIgYzIG8xOoFl83QUEhNQcFJi5VNjb0vTwpCgreaNQgjgcMsfDZuEBm9Vi7I4aDESKpVm
igowojNgOwIaxL7+iX69E2eJmMGc+UfRkOf49rba6h68UjI5wJADhTPymtgXETQs5HQmFYlSZv3G
uJPq5liFB9Mpy4Oow21BpUI2KUfdBE1qzINm/S5vDRCzlGgN5uO/8Je/+wngSAFoRmU1OvEu8JLh
1YOtOkwqCELdm2OyHLGoOCr5B7lqSiL9UMAGbFkmiPfsswPBApRGH1mdwOpkWqm6BrKJ+5obPVFf
lOXj1l6YUuUi6lVnG2+E8R6x1zFDNL1Y4X73TERpTA0wuGmcoYwDI5s+/mL7xBpRFJHPKieaDHpb
LVhCR8d1gnozYOfAVTIOZffsxntEzrF9JG1UsHmb5bc4KH9bjPXnGu1AdL4lpFDtKXrkJBpo5+sP
3abwIB6u1N3QoHTvcx/s++Xjccq0iC1rv/NByfytvRdKTSf0J6HhvvLZYA/sdQOVB74grfhURDEB
N5YBLk5dIBP2PA5yq6xtcxuoOCxiE9AZircvXkeh37b4ho1QXoO3t/Rxm8qjLE7iz29HN4EYsmho
9z232bDgAMB0QLWclpXcAJ8sGCSz9TfXw10xGgDWCWJOodDZ6B0FqNnQarMFOjU4KFen2j+7xM3D
FTCpB1DRvohOY6AzpnCkQyiEYmoqe2CJxL2xaXh+YPtTcoSg+HkNPJICP7sJvAaTeKFlMYMXGonM
r8AcPYyhbAHdAyWh7b0C6GKLhkx75kXfug+kSNbySgmsciVzyVbSgT3R1nRwUb9H7lp00CVtRaof
6yAg+BWwIH79ecMgab22RQV5QRmfNAG7FO4lUNepXV4ry5dDGltMbDe8kp4YKFmjZsJldGsKv7sy
sgFydP9DX3AMpQWQkaopWpbS9OMFE2Ec+sCg7y5a39JxjYb4Rk1mHcYCP4QpO0+KAl+lSn56h9P3
6FXV9I1nPM6xUO2r/RDJTC5JOt77J68C9ld7J60SbSIuUsprNdortvVHmmKiDIQuHdrzi+I1XgbX
MK+eVTca1rf1Oort0jUnz8escoxkhTkaLVY+xcKxPDXhkz7BQg1oZhpzeSSuv9us/ueJKPkt9pPA
Tp1anQOv7gPtnyFJhCn/0LnEx0fbOq0A1Y3+XyRZpfUqCIu5Unfb6C4zMsSrmCW+hRUnQmCJ3lO9
q7dsuROy7+mfcqUx1+P0DgC3sfbi0uLbOtX3FX+Aey8Wv2hzaYZJwiO7DQvxxWZKxmWMlxyhzwDd
L7QDJmNbrdI3PijhywyxmLx2uDaS1HxJhaLxFbVMoicHETiNkqwkDngAV6gJAbOrDEmNAqstaQLW
QxB9t2gNRNpELSPHHnTcETVMzIXNhVuAxMojaodQSmm92e0dkt288NABxCMruyR9bam/26uUc9GP
B5NBdbmFMdAxxHfGY+sNih0yAlgw74Y3OCwqialHtzJniIDYiTQV751Gco37I1OoRm0rEAq0pCfu
SHUvlhTI29vnUKdTl9xPwQA3t5QJfSqvW0uUtkSzplJyUzKgH1CjqfyskxP4QYsANPqdAIrN4HYr
1aD3+2lgbuFv0qzha7R7knsGCqUyGzhXdJ40PUpjlFMpjedHm0KIcb4vhvwOsZtGJV6uFY0lPxRS
cBfzE+yy4ycIfDqjEA7naShsu3pqvdl/BbsKy6wPmFGTcRcoAtTszBZfV9uebPffRZo07Rqt8Luj
OvwwdG5fwfxZLsh0p8PvnUeutdzCUiN+Nh3GebyfqEOE9zzDH8ZW4tx0o/iRRBwLSnIOo637ZWnj
cfAnCtgNlNAZDQ1mGTQVwe+IhXcQrA+Kb4EiJvXzbaTPCTzW3tgoMcyObwhb4ugmpRDMz0r2YZtG
dDfqttrr786aZZxNvXUFK+vaLJsf+9rjgFdOWxXAGs0mYwhDf+Zh0Q43jVPARvPugLIvYm2AlBQE
Y3d8yLAL3avSXiQ7oN2Jbb4bipKmE5soF97ZvWdJfaBUMezuuEJ1ENFFuWHmqtV+lrNqoZi5tFm3
6gaqx8GenlkU191d+IZWWKbu5+G1pSghLoH+m3TkhwWYs+h+UmQKNLERD2P/wqVEO841aqdadWyi
5LMfrn/z2E7UoG6N6EaPXzu/7oTrn32cmlwDuCodRzEpYOA4lqabgkaMf46ovgjdSjQTPVW0n9SX
iY77eA/0kODONOzk109oQXCS0LQcO+1tDtO2N+GueZZxEYlMdARs4XodZKonChJVdzJFVwRupm3R
kIHaTvPJLWUh1Nz3ZNzK4kPVwOu9T5/sbgshAbOQj1+tR+WyJ5Lj6LQhQMMEg5+s2Hzt1Mtaubal
z9N3kXwivoV2WJuR4N0Om6sYYmpKufrZIz+1afSi6r6KdVxCzQV2q1nQPlCl6WHqKA7E83vdrkYK
w9o06q6Bnq332qyoobERbFuC5i41PMEfeluYfmr9kEkgg4L7s5yhsRmPGBw7qLT7wUF/rrbJBDFX
x+PYSWAgSywjdNZzOKOT/UmPo8bFHU+NaRcrZ1Dp9/hpxpLtTD557Oumqow45XqiNi5azIhedEww
0A+6o/d54mIWl6Jq1XKWxBSfW5P5pR2Z4NaoPo4t9IWTWF4Vx3FXBylLxjxjl1Hjv3khcKWsJsVy
W9e0qf7nicjxZi8ULxPcJ6ytlIIZT5bgmrQnHD9Cd+e5BKOfH3wI0PcbwRYuMbzREZKarXI+Vdfd
I0tI8UBwzZzHzZhV2PMAaYkW7c1C5+VwsJ1kYw7NcIwLVF+VLonx4D8qq7/81aHDZvoeK/YsUwUA
JP+Jjlad8ESCFh601wK3Jb0bDK62mJ4+Y84osHbRNO5FofxfAqxptzMqDWXnxkS4n9OBpfdXTtRG
xBkj+9fpNIKHo4alFZ2AD7eMregTUfBZP7SUaj63PwTsgDC0SbcgJmOG2lMjg7sbcTI7jncGaFpY
K2opA9I2ukfhGUSUv4+UPtwkUuMAvlc39NCaYc8ZsX2kPHdPsdHOgWs+L3ktidlhsXqePudfdUi0
soPzLKcFW/zmhzI+pzW/i9L8ma0rp415RFYydBNz6eKPSsxVWbdM4TXSvsmDzXy+FfRYcB6dnh0w
kNVe1+xL1wMKL+lAxhiWcjc1Se/cbKjP7+6rjHz25l5rICBMRPAANpOOKl4jXaEr1BU2Nlpzjmzi
ng6DuYpiAwRJx1LX1yd0QGbhuStMe3XxLkcA/E1rf9Au+dasna6SrUb1yeAfsT+zbbNlY2DTODrH
nwMZYr2uIF5v2f1bijxfGvolS2dkdnMF6pXSVsd1SaduKm0JJy+FA8pPzbY8c6BeJ8eXKjR3lqRQ
ELPWJQ8F5Tp8GTsgwLSvwR/rbLA8xt2VTIkXl9+hWXSohbDy+Gi/zzucAbugMZossEw/42QRISKj
+x+yZUyigwcvFrNTGXOCtWXpF60//DymXpAaXr+3S9ua6Fg+/1cisCtwp6WDQIPJ20SCURrejgHq
PpcFN6sXNXzbeWkh2dfKHhkn4C467kWXjujsViI+7/x6r4O3Go+Wz0Lrt94LKUPilx9n+3H986Hb
W3WY4oSZaWjCCStuv+P+t5tlEJ8lXuD00ozBvjATp9Gb7QEmZl9q+47guJ9nQFcJB9oqQDqFcASK
jh95YJiNmKsat/JjXOSn0T+Vk1ABPn+cOYc7Kuid36Mbb/u4zrntqHIE0c/15QqQQP0/hllmEVn7
05vUYNEKlpO5vJ9+B7jbdM2GUJD+Kbjl3QUDfh2CPn6hD0tPw8NBdRc1A4Oio4CjjXWaoyRhLtP1
nOgCscvZZZ6V5QxoUgHCEmdm5qx8hLuwUiJGjH8bsu4J4Y3+2rzYQ7iBdYr/bcNjPWofUR8AMxIt
Fte63ejG20WqcKGuT9zXJ9VuEO3E8p4l4QjhoX0m7LdeNNeqm9yhgSnDGEvZnaFFBEZp4n1IsrKw
hzzIhagn/IZYc53J/UhUOJrXwXk4Y9gRRX603GRYYtRNP7Px9g1JylV97y6QdLW4QwEGmhSnszgc
VlDzsiPT03sn7yHtTC7s2f3rTYS9aHFc+hi6QdADQj9hbOpAALpU4dOD+/Q8Kh375z8pw6Gmz+hF
KN6lk/pad54zepuPcptXgVnMoHfA4OV9hgJ/aofheYD9IYlrIjU0TDZ4nnuGne8a364QZhCleGPi
arPvhTfWZsCTBHnYn2CTFZqQl51JBO8dOIt2/3FHipNzCffFNXZN4M7yWCkUahCHcLUWkU4a4Iz1
sOZWx/BUvdzuf4CCRU3f0fVljtdJ4WOBoiNsWuFIROGiYqrjWLOUCWcgGuKZeaK//+JPKA4umKYj
tLbIQpYG7j8coS8KqupP2QmbsLGyc5t9aSXFmoAWcfdIexG6VlJxuAQYooM2G5guR+b7T6cMmPsT
bEkHY9TKMNnlyhLUrJ6MHDHsJqBlFKf7ZBd47tnJ9OpLG1+07/gARQHpRtIvSOvT8kpullCqIklA
rxcMzCydJUGqCKIl4issZIcK3VHOm6IHC/0xikWct0cWt9vx6C2AjEgRsTW1IXAMCXbWe1rRgo0v
peDVgcLPG6+ldEwnKc+/uI+uxIPlehu79DmHwXVuNK3Tt3/l51hxFV+1Kbu5PeJeR9077HpWJr3J
DKuXUdm9hgFmkNJQLsowglavVp/o0M3lCANbyE0E6Xyu/mmrPsMp0kkGmvBMKHssAiAp+3ZBoE3E
MjtldQBTEQq6+uHATV9KkAaiT4t9n8h5oGFF2ZztUZL8WruqAVhYFE4OaWI0VtlRJDzHAc0YHoqL
COqBgHa0EG5u0goHGI01jwmGzPiDXZhr/ZZVo5PRR5yT6mOL+FwD8uCMAyRIKRM1pI0cg6nlfKTi
Onbd+RRVClBSzUk9nsN46xDM14yUIp4F122boEC25cWS67VOUABOmfgOyR+y8aMg6aGSNQERBy9y
pkGrHYWrJO4cqThYfxgonSdgC8tNevpeq2yW9iU5b3kJWTyI41i+3+zsBxypgLVLQuOX1qVq8MMU
kJfu/dLT1L2AA4uxF+MvS9EhNCs20Wu62nVx1T4iDr0Pd5vdeuiiPegVVrPq76fU6HpTWg6J/f76
XmsurQ3Jjw2TMtc3qPt4WRaIyCQHW1OUhOh7teFCxNtDr6OnKmpiqTvvxANo6PtGfX2zKWWukg8Q
HUI5meB/KT0L5qULyqQ8msY7OvMFo5h5jIlYhb84ymbF2QUuZ4dpVChlHxqRDSTYVzor4L04y/0k
q5TGBwn8AWReAuEG9XwtG280uMTDQ0NntmUU3c4o+iGxs/up3Zav4zWeckNcHNeonhV1gWVdJmdC
MvrnfG1H5GZM7aYieF3YnRvvovPmp9fbrKMjNPOy2uNccFJQ7G+N7x9LNTYQ7Ioyk2xP0IHYjsaM
ZeITh0mWOdl6fiUwW9MM6N3O9D454t84YVzrIdvxvRyU8yA6Wn1gT8ZSeDbhs8GxkUZNKu0zrDLG
ooyhcP2o8TFj2w8J1+jIpkjv4XTf5bfd7adAeImom4DFjEg7gqUJJSE3mMjQ8IaPzPrDwWJtGaIS
8+d5Mkly77gy6dornMI+icAZmw8n3FPpdfuiXXyei0Nl+LCkTdN55CqG6k1AiUl0HJVEMJsUqki8
UD4Och6WysRchQWiXYQ/zI9SgjCnLYC4HqpnHB68pMOdnZaXJviQCiifAZ4IZ/tZZ0kid7ihN0Be
e5O0KRlzWhSzcJTYgd+dsreG7HIgVgKxajBjMtOqyu0+m2FTJXrGzoiTDKaDEgrAxYfEpJqWDq1L
mtnEtdwTOB9xBV4Gqu9j8kxsO1t4kGW4jDpYONaYu/w858Kj0QqgPodZoB/bzpltqzbXRi7mDKBr
GVCh22mQgzHCHp6+XhOVSyh5SJQcku0MY8x4xADyATfEQhc3HmUDW7zIFrh+eIaFRD0DWxCvHkC8
qc2PZZszHPBgfzlOS1odRM/tIJbbcAutqiolZNVPxLOeIioMJE7Rw7NESBIkw+2TN5CRsQ7FhVbb
i2ghrV/9CFJAkw2RDhnX9WO30GsOBkuBCoy9zt7weGMloel+OWtM2FE/zO6qYF9Cu6MueJG6t0qt
lSpxcOYqp5GiLOVRAPfOXdexA2pIdEmBTl5mR7qaGdXWmtmiqZ7n5fNOEV1oL3cgnZCZfccuS06z
2qWFDcn9ChTvAKW8OiLd0RPliCjqpM+kh/84LL0PM0GGS7RLeGo7ladBfJapcAoAZRu6h4fpwsf9
4F/7NKGByk1SPJqTyKakw7PYRgAM/wuy07qANURGhsiRV/wrfYphJGR1gKGKiHAjTlhXYWL8O52P
NBn6PRPt0abRIYV7dJXXB0rMLvQtWNm8C7rwp/M7qyfv7LD5Y1/4O00Q8DlgMaJ3TEBqVZsGiBJJ
jRSMkKOdwUUkZWdSE/9ohrxXDakic7Wv/RPX24hN2GAoMgl8yGcQnht2sUnBBS5D1WslGS3GHyFh
1+f7PzBjiJFDUxSbTpDXZr6rF9HKcQ1eMEc/wIdTOYD3O4KUU0nAeJ36H0zRXsCPnPfswm4co6eE
BHzkPr0/p/56DXaJ5mKt/Lf+S8NuxgPOmxyFikQlKnHK8vOMUMy/i8uq6Cpqlkw/x7dMH4lSxkMN
9soOhBjhbzAJsKnIdSYaT/Rv0zgk/5VoFYVFvIRs9kLSRPvpMf9tK41PburDZ4hEpsuzkHf5dM6y
6rFmLtPtMxV2hOfOkwbTGqAhXF7oHZ7zdUpXZNaZM+ZtTRQASxFmHPX04Abp6gbCEMrwKfuIZ3fl
nhItSCZU2TwIk3JDfUcxMnnTZ1c+x7eJCCVQd6dvnouqcPs8ZQk8ElhJ27Q54Mexc809intwi61Z
m/xvkX7sdGhuUJZx8KjDcRbvh9ToIa3iaCdznr+OeZYnOt93nwydu6PFqmlXRYgBXAnMZiMwiVnv
bBn/Y7cOb+FTrWKvZSDBdy6FvtHrpUbgDRFmk/XRcjoRu5VvRf4dHwVf3tC6vKds3qaH2JgKe7Ol
8GgcHvwStX+NrRrEV45zzru5FCQ0cZyspmd2iq5Z7LErdkAiiq05FwTOHukWZ8pmtfbKxyqoFAj8
SHOErPdhl+quKYlMgHCa4eic/DzQL9IUTzL5I7qRbHmxi548OaaXDpN63eWMQzgIkjt9JqfAv31B
XahvUWkz7U8SiGF5D/456uEA9QvkeIjSfISxBNwQkGS+/r+Lx1TXS/KsBJm1pWyBVFPHbli3yu16
7fcuuN6I2SZnVMePAS/Tf5mkK3PcdPzTc/NjoVK5BFd2geUDrZYMAlWiwzzRAiDn4+2JrIpdZ3y2
uV+DTM6UvoRlCzRjCQ6mEEVwuby9OqinZE0oT+PJ4mhZmhpDTehyY6s0EqEOEeccegwxKDdlF+IF
AGIG+pBjUikQJwwuZt+Y6mt3X8EBqiHwQA+yAQ7vJ6l1Evaa7zzeKI5D7jfQZu1WyjaNpDf0rV6x
8TrvgS+0Cp3IJUJyZ35wEAiaY0xrzlGfve7w0NSvNiJWVepPOZ5A/K6TdpDom/4mfjg3Qx4DBmY9
uU5D/GLPVj5rs0AFFM9vHA/8mprvu86ZomWB0DEHeQcUpmXt/lIrseKUcjAVFAO7LJjps+yHVAXp
Il7fUqFMsqqj9d5jDldqsEuYykj6tsxFk9cCE91RZuOdf7AXk4xE+D86aCJ9cRIi+BuaIO7yiNAF
8v60rkC0caGpZi/VQyyRWJi11RChgi4I/UrAp0Bqbix3T8Hcqn4+cNQ7g+W/rTv7trrUDmZs0wkC
xUy7yiaBTHGYjp5EcBSml2ldkWTkAox1LjOISMh7/Mthl+Wf+bKIYM4lR8VihOeNPn19TGd7tRC5
HUt5UvKXl2zoAMLljDj991QBgoPLPsr2mN4N+Hu4V7MxtcIYEEXA3odrolFckWUvcKno0/CS8s2/
OiaJglJc+GqiFt71O/I4ITXzEQbHpYDE+6blBz06mNC3kHPKnoqVjuN6PnGwNyTK6njQg8v+jiv5
P7mJcfMywZRo+h699t0iP0hxsNJQjKvJOqMmV6ZKhyN97ZD62tXfw+hjUkHSlxzNZrqlGR+tIdzn
Rd2oaelBBClzWqBChzlwQxPj4+EAd3ESsVDKhJZKaJtEyg2vCdylXuVXcNQkelMmPdrxHlBMsjdM
4/ayTtB/wQuXSvb4ST7z8aehGcpvieJcAmjFrIWDj96Zj7/5uhXby86nGKZcbswV782biUAjTxtV
DD9dn1u5HV4fVUhr2i51Ju5IZ4Tk6eYinXJuKWCA7P80bagvKbVr+OoYpa1WhZC9gX8tbOsBUdGT
mqPQXuJj2hlW/tm18RAIL1aoCUuVXh81ZoYYhsDoc9YHCiaeZe1/RAU67DBGTQz3UklFiMfMRux4
6lPUGO86Ozo8Ghhz7RaHsHs7I1iONoy+xM/emcqNY0AoSLoUa3OhXvwZEX5RcA8M9GaB7MFydIKf
xJCi/lLFQRXbDjqkZb0BMGlxk07l4L9Xx605LLm3AoiMXG+z/HQns3orQ64O6WQTv63Cvv/BLfMA
uYoDqTw4S+tq4lI99LuzDZMd6ijNw5D+2OvSc/ukP7aXQLf7MSnDbuLUfMWI8mvXseBb7RyGbPQ+
YJ+VsMozqSgUnAUIrOn23QETLxYKbLMWcrVtFJOa55tkFREr5Uj5+/TnnZ458c9RHQPiJytlQAjy
STIJgAOxV2zZJqEHCKZCZXu7FO7tuf0BZcNuZ26fUWbadlY/Mzmi1HrD1s61RV+RyBs0rxtOZkfs
8kuLCMBaScEBqtSLNjx3bElT1YHni4DSY8H2cxeoj9C3icJmWtMMQoZ80N6m5/WT84ADUkOSJ0pw
jgKZyDJsJrF0k5H/1mYlkiJO5XEv6hymk8DM4hnNN8HwgUNbz8Rq5DKDR8Jj+uwMqHOvrggUzANX
5E+eNtCUH1+plt49lIx7l8qLq49rcHqh6qOW5/D5QFN7cl5Hhzh4QPS+WmY4FA+7NywPhtMciBt3
pdJfBwNgs8S5YCZHaNG1xDbRbwO7xNgUzon2W8OUELHfpnEq79b5pQtiNzkDGNHsXOswgvG2TESI
CQ8l9F94I0pXtuH/XFfs/tuS1z57niI1R+kNgpEwtzyljTkYYrgifDQL0pp7oA7QFM4iyMLw3KoI
MDN3OvwwsL4rrYnoaSg4eRpxsbsSn+eb8MjVo8jLMLrXiZmSxty9zY/dT5iLMKod4V9S9IPgZW77
pKCJAahjQnUho1AEDthpEKTbY571Sk0imtDOBMgUi88oSh4whIcdy6lTfu1E8NckQZ99LduOm/Hh
y5RPbImsAlXym2CVjHx+HQ9fQX3IeQv8eq+B6bA/lnCNymacISq27m2IYEUIBcWu6ZM+xwEZlhpk
V2g7xA7ultv+kEzOB8RnYfENJ9oyKEp3WQuv/Tr+kUOPPMN/mfWRqDHdAOBR33KBhmIxaRaFNQBc
rTCdjHcXSR6TAmTqyEGIInR6DgGM3ea1eNDHMFO+E7ojvfl8Wd5eaG+Tx65hIj37xCC5IorzP8yo
NLbf4AsSYDCmQ6o5NTZEdo2OuLcaZKLZhmr1GotX5tk2vvr7OSpkhiqcPXZbdypdDZR541D8y3gh
k10BJFO3oD/hkISxRaPehpu1JIxn4IABBZfMxiXa+YpJbd1I/fGLXBdh7b0vBE+ZiSxNkJ66HP68
r/HXF4Ylalh1gPy8CmQRd+SfDIkNSJYP10g8C82NsSkIEV9lWSA8MOlMffAjBGkW7UzaRhkPL7lY
s8RNqash02QGas1+lBDaBKKxqsbpsO2+vfOGL4I3XaDsedoEK/soSl6Y6a2KDcsP42oEO6vUOlUI
G/695dyDyvMZne/pYyMWD2lBVix8/+pIIpBf2XrhSEgWnpYu+Y1j9gMZklDXBl8HB+OiTaQUk3LQ
bbDzdGfwn2SuICW01kpW70zVGKfwB1q6JMG7FWo0gjZIRZ4gNkYccHlYxyvTyOjJXXBfKFcTkSwI
Btk/PJC4QHXVrmdqRlE7RPyqNbJDHPBcAagLtZFMNuEjI8/PSsuD+aaH2SBaM3MwxgiEkwWD1jvc
hKGeKdaNMu5gI/NnWOvxBjx/XsRn4yvmdwzgWp95FpNnNTi4O7AYyLEefpS+XmJAueEfd7LqsQAE
l9SSuFPIgyH7wllWlo1glUrcC+7iRPS3Vipqywlo3nSQTWT4Fh1mRiDoo675hA+RwNSHgueHv1cO
IfVqOhuzj0/6bbECrTWiYcwo0gXAflvv/f3Xpb3eZJWME39ys+ONu0Pax06s/AfD/DvoH5K4sA7t
RWSWSBx7ueK4C3qmTX46FfgNZN7bQteQ7gOZw+cgkJ431hoszf0LKmSO/uWzSLRw0F0Z0eeNvdUG
ijbGwrtaXU3aWYudOuPSVtmsYpIrz+Y4f9AVYuJNs3KIHB8oVHgthODP3TQq4WaFGdgWwjhb7Gl5
TwbMMmj3xCm5FCjZc3Dh2dWReoywcNgOYXeOjsyLSk7zFIUyFv683as61oYbU6YSCg2XQuI2L5ih
qLK4E4WF1nXhQUAywWhiEkzZwzjn/EotOEWxe3GVD3MzeShoUEPvup7Io9FZaIjEFDrlDcyBw7rl
rqWSrjC0raSzWDMlXVoD0iS+cClGVZMDHLyRg9XjKMe873uq9GqPBcUVPOCopFYQ7TG6cVYy3Ly6
gERnbUj1IQQtv8dbbRDor7lxpeum11K0qyiP9/IhrMq5M/1d7SkbHhMViWnEVt1+azjZdPMA8aHc
e2DFiyahqIPUNCHmA3lotUsvw5X2MuflDcH3vsspq3zQyEY8h8ANu8sxcyhcC5tgopUprsQ21V6c
1ycrqbQ4DOQxCQx+MjKgCkWEoMijAKFyL9ONKsEutvvEk5zHwSeM0cbjUVUzY1jXz6UGvaf7x27t
RO/fEmNvjY0iLpRaG9PuSSJbgcGplxd7kU4qLHBEh+xpgz1bfh3xTXz+zYm0beZJdNvQe2Pi8TJB
sD0GJafoJlekVO4lHhaWUfPF2j9hbtqhgQVUm3d3Hxo+PGoxOSIufQMT4XzV5xt+FopMlKtdUp12
atdrfNie+nyd3uzIwf3b7hQIGee4Yy/OzYTN8buYPuYQYn3NN/9Z7FfCwyfcdQYwNaIPi8mzLe+E
Flvp5tgzex/UKyjGVde7hfaueHJtMaoS+qi0TSiYYksbdOAqtOi4V9HLyYdxRXVPOy0FJc3Z887A
Uu/QYIsHmhVdXpKTkEwZSiYmRlU/tWDMdNAHVXH91ENmim6C0TGo+mOnB844bQzWJzp3h3dLlO9L
yQ3bJRN0DDj+eUWhUQb2Q5adQZcObV1Gg8MVtZww78WX8Gy8da7ZQeqRtivkrcI2xit6ju+z4kub
SQ1hyeUPtAhsmpObrbV5DHKyCKcdR+ErMlTO6lYV/ArN1tn9hGRIaIvhZNUB6ujEdqMRo0q7Xmk6
maJ/+m9KiUESPUHe5zV77tXY3E8XwiCXhgBbx9OsmVOkd1eVVIIMn9N2Khh/2XVZNKISUaEJiAv3
+9MEinNfE4S/e+DdMxGuEVzfxsykxPCy9JEwIDX7PdZjTfRsoNQ7kadVs3rNfUzRM8qM1LbDqDWj
RyLEbkct/iDKvgN3P+POYCcK3EohvRp3XOd4MG/YYfl2z4eNd0Zk9YrVOHQVDsaDB9VQwunsz8ka
L+7St1KtmLnJSjSK5QlFuwITosJqRyE7+1t42J5flUnPBOVnk/nOeCNVYsWlXsayfOdPTrcjUUAW
ki6zWRJsora9fk6wiT16+ggdCIcHovQWYgZxtpopP5WKIxbM9uFpEfsqejfTRgdtrUMmCT0aExYZ
rGEEdTXZSIKYEZaWUQE36RSMcxL5oiU+f2cHb1gn7S5a1l5U4DS2pfiwM3pxi2E/ade0VjW8l6j1
s/feqeW3OcSWx/+SXqV8NW2a53qbzrChkRyiBAxQl2rf7UpTwr7Za0HKyIe+G0++cmAY5V/az3r6
MhcB9qlTq/TEWfLVtDkCIq/laohjvgxS6P4sZV6oVwsWJ+o7bVqo6sEcBp0sEE/5OupPezai4ZrU
TeVxD+LGAEwgypzFFRX3ySJ5dzoY0EczzYc7jKNGGzY+rzoZi9dP4hMS4mj4fiMWdqGirqKd0yq3
8sxZDc13LrLaUm37fKGVTc0nTyJD8VUzk883kxItLYixD3Xy/uniC8orrxZVFBMXRXW7UV5jUAe5
9Bp4hiF2fJ42voHQ6gWnFi6a5sVMEXIJsqvyXS7MwrRKSAe9PQIPP/aneFgSYfHvtyC6zYAUqr2v
Rz4moOueDFKk2pVNuK6NwIB92Kn4QUHMBz84WdzRhmQG11WhXcbCk2cIdOHoMOXe/GgYiZrWliL5
vh55v2HdrDboJBhnH/VZuK3YQU1GTYq4YbGHBYoB4gB+qtSR+365OnLz+IUyEO0dVWbXqw6pbjmv
NLRWpxiSOJNT8EDIuzPBAcqwJgp3bEhLRgLBPRgo4PFRdqtNRtI7w4GbNk75Y9VJKcu8zUJ09Vu5
7cnY53d6mmzZlpYQ5X+JBs6IgicBZMB2Hlx2/bpedqI/kBPcamq/w7uX56NsJ5NXDSQO5b0KCVx5
EFwvlBKHIdZVKj+qHQQLZ/CFnEiNfpM/h5Kk0HHKkywXai82J0ct0ALwIXsA7GFHDNG3uvvXzcuF
oRN9L9RxfPaLqpsYkm5fI1Qe3TBJaMa38AIJiMQU2EyJ/YSfWyiywsCqtLC0AplOpkrXTU+N3gCX
Zj6keEuS+geJhna04UQWh5+s40PBA0RsHCQwjj1Ijjf0XfHp0v1eAyPQfqbdyuJM0YXVgv/nxbm1
2UFySdCvh7C5pbyplJeTGKmJrLFSZpY6zOoSziAhbivdNneIdsCMBevOLzTCb8ks99S4V1xPS23e
4rIlybvvXEMTutqecFgBhDng3hH+78Y4Co02MtHjnN8ZrraBLafdod4HpA3anPQEoELmyc+tah1r
TGKvV1ura/GaJUuuPwgL07gn4sAbR8gwX18aNW+KpQAQvT5pAsBqWHAHgZ3PXgDd2nUNtJCUiXmM
C0olVuLIWLuIK7Y+JaV4DJNMlO3OFlRJqedwOCaxM6f+Hoonx1qf0FQHcC14mn8iwYlwId3vFReY
ZLmpJmXmC8wyZIwrSC+R5/YDkTW8ULTqhtD2drbbpMJ4jGrSLi5dpezUmkKDr3/jxq9sAIxG902H
rDykhjahmYOs13m2WcNPVDrvC7obfwCw3mTPcD2RiXsopAhViqQb0derTRBw5B4lwezrwGB3kwWI
my9463agbvHODfd6rvRpEIxykKsYhjKDefx3WexmASRj1Od5X5uVUs8HCoQkQDgVoi8sR3mHuQoe
UqExsbCq8EFgWOm0RTMJZ0kut89+NFGuN1BS8WjygiX0+zOeydeq/WVeUoLkNxvgTpKcducbMhAL
buefroQd+yyCeXdF+9gafvSKF/AW3CY0GzPeap6rK29nSqDGPfoEkV/AnrZJzCBV7ca/4iWuCiXT
2Vg12bwKaTDKs+fPlKPXUAkDalhmD6yTk/Y1zMareATAV0k5hwbtyINDNYIaiIVX41sLZZzi7mVu
jMjKb1aQyuvZYrci2PYEFOh3/GhU7pR1SVHJ9ArV/L6FAFQraD7pLDKxFrEhZk2lBEFrE4Z8VTJh
XU5G35P4iczWkfPJVbiS2dHPbGm+q3JXdAxtmuo818S+fb/SuGFD9VXJvjyi9KKc9HUpRDZ/e8zk
q3FBbX5Gg8xk7uhKcd/lavZj3vlfUB0YzO/mVZkhfo+hkRwGTJYHJaS9b6FiFQjhSXNVb/hUMnfW
QvIdYwYN8wJ62r8n1yX6GBs3Cx6KTzUS0egUI3gGeL6qRm9vwi2VJVQKeWOT9SpWuuk6Z8oXp23D
0lroc0A0Odw1lUONE7fCfkFi8mDlRKmAtrb3Ku2qOUIBy5TFVoH5elJUUMkLXqurWOMlufVStwX5
6eYKeUTfWSQcS13CrGoTaeK3LCeUbYK4/CwtYHAegjLi71vOoliik8PV0VrCzMHrR0JJQw4w8igA
cME6AvG/PO40j5o3TcdonbhFeTiaAAfUMR99SB2XpKlksoADM7K8XqVGULdM3fMl3dJN48GYcdrf
tkHGJnXgmzn7SedK3cKx0761CtHoK7eNPX2NQhtdVR1BqtFFZXcY9QMfI1fTXusTQxuCVHSmcvxn
0ruNWhaAh+75BZsPrQH3zmNhNbz39h6vO4ouUcRBFLcOxZKMFwcotuE8N0aLdwImbOABDWcqrtbj
aL9XDXWF1/QOe6hrdu095mK6VqmOdtKw7xAPW4Uf8zCY953edRIYocebNQQefzRf1hL90xMzkPw2
qpfTzQJSUfhfyARwRbvMaBRb7MEQPf/1IWoqUVZMDqpdnnMtJ0iTd/cpmwY0CAm3MeTS1ggfWsqL
3Za/I9MasBVVP4caB0O3iTCNRTVLlcC3fh3aJP9BqY4XLHwYbnyGfe17QZ088kajzd0Bh5PskxN8
sysbm1oR88KUDQj6WpBZXj7/HyS8TanspMTRrKOf1Vm4SAnAXkfa9JH6JqbdksR8TSThgvKVghwi
FQZz0L2W7BVHHn7BvsJMfAeR6B57OQ2aDcYDi4/OrTLx5JeJeGnr1T01YwfnGuKQ20vXqk6aeyfz
dBxKVVuZDskuqzl03XSa4zRqICJfd9csDRNShfogxz9FOTs3wHo2iZ1XJokLb0defIHigTakR6uU
DS5JW6cha24ryiMIpvfrOfyyWtaNdw5fMPPwjMjp3V4rT7kdVqaAEvvgR4fek/9vdICi8y0Rtz/N
xZrO37fAqCqINDZuyO74bFYZEz7aMy8ZY7DZbA4siCpFBku7+MuR8KwikGuk+bQdjYbOqxNYh2sj
CQ6tsVi6DR1xvuKAwNncMTB/ZKLa0L83OagdnoM+5EWsjziNkuuO2Y9CZgck1No9ZGVhUizkOsAm
ODLIFDXdebHmEcgJsgd5QOOk9ZuyiG2rtf80MhBWhteKyTjzrqFBlmJ1tab4IGx63aC4cff0AlMm
Q0NCm3TB9GtpXMBOn74nmaIoinCdok/1rjn1DBRoYpUF8a3SGyWdBQ+dEDRJXzi+kpRyJsD21hDL
+go6ARfAjaE5S9zL04Izw7jTC87aQ2Chm+KDQf9uot1AwrC3RY2q7hCHFfc9F3Ul1iql+fYx4NzG
Zihe6kdFi/IHhd7byz7wWjmQbPZ/xPBMXMsX+O3fET3c8s2qzhAqV4Iga0EfEx+6bIRmqe7Eqllu
YQrePk4WCfpHlnjhKDUp4pHP8IcvQksymolEMrcjMtyi3mStgaHkmOQJh/ocsCQkuktNRNDt6Skd
RlXGVTqHHcIJFKy4L730bA5QjKjrPIgoUj337hNPwMOU1mrGVPilGZ4pf23BQA+l/XdJW3AX8zR3
7cUgGTe8jrOYWPEXiZt3P1oXFNu5zZNVtxk+jLWBn+4z122qCDgn4FkuvSBJ4do9ecAjwIbMStq6
ofyjJP9fsr2v+UhH6pmGkJ0ryOV1bBnUAv/iY4d/wBRpHIvyK2L6GJwEsYjOxMxiNLLT9LWgO/zq
crz/DKxx7ntWZixwIXTcycXLAF7qhoeiO6LSWvwGlc4CbiRZK6yy6shn2EVpKBRYKHzmvC0ZIeaP
rHfjeGfgPagSXffIXxN/NY2q+v+Wzrzxq0XW7SufTT9S6Z1MorpXTFoFsVg4oUiC/Cs1ORgMLyGK
r1YNPRV+dZzLDmccZ7JSobsfxKrr+7z9kGs8gYIgkhnEQ2B7l8sX137aQH57JmuxaYYcXJwL26Ba
0q1htyuNe6q1kfiiIxjRr7sHYsI1hQziEByfTnXroylA+N5cn53Hh3Vz3h/8K+cu/Qw7vxujtnIV
gzHOPfDZrjCYIfYLqu+CoEFhW6qYQe7gP4cq3RSj5fKjgIqIkiyHdtLmlitBtvRutPDhXZFQdmx2
C9sbAxC3CvOxCXo8WPxeWlvgW2h8tFfLZV0SCQdEwDXH1EvLJTE1SN8A81hcdVwOL8wb+kEL2Z5q
aVM5Xr7CDJtXVMKWtPorJfg/GNJCFUiVgmj5LePk04KIf1zFmETaNEhK1Ruk4ZjJo1GkRzJzGRO8
W4Nv4t3GM4r5nsyv0jOxr4FEcpG5KHy9QY146wzfDsN0NWJGf5wFoSjec4vBS/mTMWtC1PScBlfk
BuuumD/f0bWZPCKi+/oky8laKYqQJAVtQHOChZ+f0iP+rsVfY5WaHQmSfW5s47QBMyUEZ4rBAVCF
b2GUjUFNbfLnWkICJ4E7s0utFSAXMyN/MCWgQ8bPTFI7kqUmSPdFrOKS9S4L/EbsbNhmmq18i2Lf
acHCMRrztWQH3htFAZpKhE+Adr88sDHvtvLqmwJT34ErqjGeojExPx4QNBDT/ZrJoL9ge1jx9Y8N
9U98yhvFkckwyNcbysFliqZO25QHokH0xdg8F5/AV/wtOr3a17OQkOjCOKS8jby+19tzhG3pi+qp
If7RAQoDpJbLYBkNOdKgRPu4ieUrCd1X5JvOnUP0UnDV5uzaBGkINEiQ7L3pxgUSmMdiKHDg+tEa
KImEGZvjHMILx3Vf7jJiReTeBwdyIw8/L4Js7+1RXEE7clhoUGtR43o416UndJwn5N777fPghQ5g
GFsgE16OhUFp0ob9dhnIcgQLOU9BBuvZZpfiP3Gb/WaIAMJkwqTaBKIb7pRdqGYR1mlydBMgJR6g
ih0I8BgY+OZEeEFqZ6TKWuBSRMHGm/toIWMy1u4cpsIj2TPQcGX3k/Gtl+rC7zyeM5Dyb9+irTqf
/OWii8IvyvGe1lREeU3qlZfgh2XoC1eEaErIVEcTMSxeiok+4vbLcIACsBXkOClAii65Da5CwF8L
nz8hxUP+B73TOoPxPP3ClfezcaiGzWtsjSN3z6BtlIVJJZEHQAdUh7VFFyjoZ53SRXxAp2a0MCY6
/INmjUP78kmJRItUeNYsLVCC5yXDjLRvSfTGLyjxI/ew30c+eXoxctTv+W3AqwaHJfM+pKeo+bQJ
R2ftYzUeX5HmGbGts6n9AJAyCv1W+nwS2WN/iP9pe45W8qOy20OX0xnoTjpxvNZQdEVcGMgkeSrK
uRD76oVdj5osTPfCp4UZfJCimB3HMkq67PWVpBTliKo4+EvotuODSv5N+qC9SkgSF2UU9QDwUtZB
MJi2OmSnziIWW+pBFuyNgjTpgOoNZmN4VmflxblJZcplJ+btNA/xq/qq0uzENlHa+tpwkMXEuq24
bhyJDe5J7e/7i1FmrNyRed+3flFJnK+KOS+q82LtyZz+YGA5MWS+a0r8LtPNC3NDHpHP331W49Nd
fg/9jJPITaGV7ldmbZ1BHWzagvHRlHdWPhePIJo3Z5KV0YkG1OJb3ilTt2kEz0+ff/KWoPuAUlzu
ceS1oQ5Ajzqmkom7a//1BMCR5/N8S3j2ecS94IzVJ9OJgLP8Eo99kPEI56cxch4bkMOBwTCbPjjT
vxVw/C3dwgML7mAP26yfXhosP98mzoGlj9G6z/Xe5378UGh1CytV3ul+66cLMvtfZXZaB1SxVnKw
0NcOV5IoG7NZmac5ZJv+o71JjRqijR1MkKQkP8MsxpdKFKrv6S50vkep/NrB8MRCj5PTXqlqOqQ2
SSwXlVshFhDYMco251FLU+ZyiH8SN9NQ35YyH45XhSInCUoDooi/zTktw68mDr5/WL5Dr3fFkNyt
twNNDt6HPR136PJSqvlpTeGV5FiumktO0pct5nv77S8Wg41wu3Xd1XzXMYGIlhVRZFfVa6Je/2B/
LkvaCYZE8B/CyMejJR/ubeoQTILrt8OgyRR4ga5phSDptjPaQtM5dJU1dVtjeoer5TXKAtfkBAQN
OJ30kLYBrFPzpetcv3od7Igary5Oo+zymarDC8nMQXMy0OxRQdADwiOrIM6s+rViNIaxjkjNdVPc
2cgngh95Z1fZm5+yXf7PmAc0IgOG1GXdmOyE2ARLz00aMKg3NIWWh6Pflnsl9IExgBFMfXUL+1qQ
MDmhRyi9Wq1zhJ7bd+jbkxkiYaXxTTvgj2+rP8tE4GkpvBkpkoLEsGwXvquKHYOiu1DBnEn3X7GG
6kCNJVenl2FrhE9Y6/1jNydEXqZ7wcpCVIexx8ly2HCN6d73wufRhMb7sgTYa4+n7m+CelXASVi9
hbRS1e4XOZUdOJQUWAo72+oU/CKczXOI1SmvEuy9Lgdm3Jif9gYm72JGcmnkFR7pmprIas7tz63K
4xiwKC8WfHyWNp3psaqbth7c5usSbCfmr157vwpVQ2CizU6CN+GvD5ZS75R51IktVKtoPKYaHilg
Rn27Sa4IAbbUtU7bvNfZhMB0YGo+ZoIot9q1cvNhkKj4/7Gvw742dgVsW0+TgE1zIMahP3waxE38
fDyqOQyfFqkmF+TvROn1gaH+EE0MfVlWl6e+Djr30l30bm5AqzJSJ4ZJfMwe+RZ/jfVPPvs8Cq05
KECiU4KuvPLcN79pHHk2E32cpFsJ6/1iQJ+l/615ZyE6PLjlqB+6FRz37645UPJpH6393ZPdXg/O
cTMossZ1C9nS3Yw7juoS0peWmpzdn2Qemq06G5OlXJUg//wJG8GHTYhPFSXW+I6SWElBiaofkXha
77dNh87w+fIlTULS9z7jSXRK482y325FBpX4YZIztGAxVzfOuVrDTvl0hLjBcwqDkhVcqLtW+ocr
xm2hopUIAY3QGbfrx2evLOuOHUGtSsg9QaIsixdLNI7bfPW6OBboJK9l63TkVX7t2vqN9hGr8d81
WdIlDrqxD9/UJaFz/kh912YEy0l4wCraERGJneZhVo+nt48TBPWPszpVI3PYotmIdRkWS24NnwLK
gB0qbZrTesov+nB1IiGyves3ZjCWkDOaJ7DfImnW1Xx9mNMVXlF1nnI4yi4UeGJ0/0feB7VHqfPX
12yNMuDiuikq3Cn1gTkZRg9v0bZFcdl9euDD/JDEuBaexqch8VbHLyhUR/fO1mVsJSvS+Syjk/95
Dz3/Dyzrm9kKOAt45X2ehPeVepCmmOhpiSMFWHwRgeoPDpNbODaWP9b6LRMFppRNqrcatiql+dSP
+ojAoEDFxnijM+1FOXB4wNC52GHw7KMsBS2EZ/7QL5e0ZHu9I++ci/ggRp5UhuK6b/F6OiexgWzP
1bZ+b5GLeH95Z8BuNskscSPn0pB2tHMSmneIs3KtUBIdlFzlZpsWCn/jP0/9NFF9EbcRSu1Bv6LN
Kb8Xm4xD6g1Mrn9EQKQrkewKoWUjnLY2tj1c0s/mY4DcuzvZGGtB/Dn0aJcOTp7E1YjuPnu6dy/D
zJ4jnaBK3kNZG8kVJV4R2RnK5PSd92ueug6f09asnN5AMz9gaF3nf9w5KCCV88CueV5CbvgDGBP4
p6teCGtrEy+iK3/SuAUF1siHK8ztzOAa22h5Ra6ZcvicL/BabEbpGDuNpqgLa0EkejSg9Z63hIL2
wfJG3fexBZcRCA376W8ZIHvLkgrap8jVNb0firGzZDGSR4mfqGTfJ5ffBynbmBQMmxCl3jAtK2oL
HIw2yHDH0/EH6iUR7NK55Aol2HnddI4SIdblT/61etHAz/SrZgB/PXrxBfR4XYQwBUIaZyUHEVA4
89LTmnE3BloeWWNcYlrIk35tN+UShwZhrpftAt3C6fkl/9Tl/sFS/a85d/x94TvzWPXJBHCWnSKz
v+70+iZ4Faqr9+VFrePZ/OQExY7kdm47IkvGjo18a53eeHNk67iGUkOwUERc67mWBZH2LQICT0xz
jQ/5BAAPrN80t2Fe6zgybOmmTRvduLekFifRHV9t/6g4N5yM0jHZqYm3UkUMhxi5Gir8YmMzviTS
8VGh7FcjkERdRaZVRrb1G2lrAQdFsRCHzq2pxLzfo/2pmJt9mm6RVSzru2L9Kg73gEE9pKJaAkGN
BDqW2mRP9FqUDkKhzdhGjikZFVPZiv39UKNmnoPXx86Nfwq4bJhqH0RBRTm1xPq2ijIaJH7yTFJL
4PY0+gx+LZ67E3S9yXdjxTw2HVNE8KxRIU9trVF0fdhhOvcOfJwqoTEsCMZT/iflaCItSnuMMQUi
NBMWGO7lrG22XMnvRxf6hTfZTwUi/VApnPuuyylOCG9JGS1e1gt/SekFpPF33Q6P+zILSYyF8zm6
0fj638DDJg21iJHlFdYl/zWeRqG44WuV9ThNWeoA/etQSGDB2GQNK9YxvwvAQoaw2PVsJWl82t+t
Tb0wY1mq2vUTxTCdH29V29Je8QNmSSX0opUQAegAuCvhk00Peb362Ba2PMCg9kBLRjC9WiYAIiqx
POKN3o9oSdpoSxjASAcOIExJKBE2cd3qIQe4hzjP3goDpLGZ757c0bZXFjSgCBDza5WWlxuDqljZ
BUXXOmchch90WwOXI1WPR49djq4FoUR/utWzfI9PogN8i5rdgotBfzTdAB81NXs+FylMRZZdl+As
QjiX9odArRampCTA2E7SbfNx6ZS+bg1OBpGX+0ZxM6ii/MMyAE9KoKHq9zq4mFDcwgrLvsaGX4Ht
3GHxJ3rHBJudAv2d0H0iBBDksZlA6rTPKNyyjzjruJVNwnlcrGVsI3OeR9OX9xPAd/sdV8N2a89N
Rv8cPgNGjXZg2L4QnGag4/05/24qUoEYLUAoqprLS6rMMUrcYuDEfdC1YVC+olK0f+zVNXtTBVIu
06ujKIcBII2favqDDILXCijZ3pUIvS8P80l78VHiAmWFajF24oSnQl6RD5rIWIdOntLCtnxIjXE2
xEeCx/O7ks0NgUgu9fS3PCcj+K/DBlH7ZLKUE1G1rXGQD2a/kyJV6i6nnBo9WGKugi/FJpsOGqLs
3NUxcl7ga3GRkvlYzVmOyKUbmXMcW0mI3Dd7uJQh70mnkaU2iEnbaW6yy/k5x/Dmhy9Qim+vy5oQ
XWhdb9ysdHbBcThlyXJun+aJ2gUdCiP9pmupE/+sMpPW3werXnAgEjWmyR3jUghyNA3mT1iesQwj
gPOMULGmiBOjI8gGzNcVZPSAq0ufv6idnBBTylfj7YpO83asY+Nbe9lUleDDYB5KY78sylEfgLmz
q6Tg9ADttGT2McmeC8DRM56JKEVq3mwaeY/0kzZRGhvqbIiXhCqfwCFckJH4Kcw4kr+pa2H56EC6
qOM8KOfyAtv5vKE7aY2dUw6dxIG3CPnqv636NeruGgmwn/dBAsC23ghM0NwFrTAXK+HYo2Lpgrej
NYRHG4njg2M85Oczz9UXwnrjLyEpDjyXBwyc1LuO9bJusHfLiUP7WsfjfEpCJgS4L5iAyt+Iq61Y
sYpbsUpTnopDHcy2ltJu58SEmbYl+hzPanq09iEkgHcyBrdcpxWcUDCDI7voqh4Cg/dJNjOPUp/3
/kWSUiomWnrtpTQFIo2xdGfgIgIrh422zzRVGe5u+0aFHjB59GA5+KsmKE7J3g7+HYsXGE/ZgWlN
MnlXuNP3XaW4oVSZEPAIfmahrltDmPcm37wx/Lq3RK5IKkQANuH96IFYmzlBAvHiMzzv6OzQ1aL9
BCwIMBWqujpH24J4u20WRVeBpRcl1IJSj+Vg3764WbEpIMGPJmZcQ/pYynlUN3dy4J7YUu09+Ijd
EdKV5gpfgjNZ+GmxzMRvN2E/xJJzDmO2r/+ZVytn8zFyAnSRbZfJbVS4c7R2UoK4niKHg4MnbNOW
oVMjxKUo1xgCVqKagABtncjvZmq3pldW2wU3NTsSn8M/0TKFrw2qDhe3Fulhimhd1TGJQ3V0F1s1
dBtYhqI8sHA5FCwFPIIupzocdHwqS8ORoaW6xH2Stw6rP8tC9FR1tX21lpgj3Zlnxp8V0sNWhaGA
eDmFLGb8yRRo3bI47BFA3GzG1HQgkIDhLrnG68oR0Mk4ziGHFrnxK3IJyZCwfKOyP0AmF2f1zCMF
HijWpbi3GGZqnPiWtHWcE8y2EizSwBWTr0avYWjSikd0DR3vPZ4d679CTFQ8c+7BU1cJ0EqfmYK2
j0siAiQgx+Q8dWsQ7F6zXHpDHrrKi4pkihQmm2ltdCBhUxQJocWP8O15ZnqU80yshITADaNctmXT
HZRrZUsgQRHHL83Uhfb4Eoc7JdpvrqrTDzYx2UN4Ox7JYaLO4PNZ7ZIYs1s0ZW0C3JrFYZdM6oVz
rQ9n5jS65My30kiWUclWXvWwpNnspCNTzJRI7o3oRtXv0KaMGCjT/vtJo2Mu9sNL4LK+uVMFf8PN
AP6TiBDTjPm9LJSLJVU7vSRO2O4GyJN0irGWdNFQ9V1BwFHATQemTmTe91IxkLKdyLLmt7kxapZr
+j7VZRLuWdwnZ+NnsPLyDMShoj8aSKaTnD8vxN0J58AX0ngMAXZNCwiTWaXoU5wtSRw1ggcks0VT
Ko21kZNfLTvwDqRr27FlD36aYezE+lSY1vZyUIPPJCn3mZ3aR23uvIglQ/Ap2AoNHiPnZWPokQsU
HFzTe01BKvKUh904lgSYeMifohja0kOUgwGkouUoR1982rfOe5+4ZwVnS7kNDG8y2+LuXbuOTCSP
Ah44e0Of/ux7grfJ7ih1GCL+HvEuqlOm9MTJ24Xzl3YpqeJJtPGvlie6TSnupKxxXPvKTVIX78zc
Qi7U+6X4NOPQ4xxdf6HYcfuvW+r7/G7fWPhvkgvV4C4dAhEX9FwIJZ+ejymhDMMEWX45+E8V2AXS
yavT+4M4yup6nLFdYMs2AIAefuHy1uhfHIxJ7hTWdRiEnBAyIKBNRuIyn/bBHd3+fFrI9HFCelM3
7NCHB7FP6X9mPPpY5E0Q7DyySa+XLu8G/q0ux53ZHVd09PiWIcBDWrMxu/cfaF/e/PE0IFMCptoP
PrtYC1gZpxfUU60OvWhcXasOg5C8xH7lEXvrJC9TPhl/J3Pi0FLfr0VTUGwadjcRLrCwGMILL7qZ
1eMKn382IeSsZGuG5qz/DDOmCMesRXOCVpG+MzbhLb2SEjscH979S8kHRV41qpUE2C+pBdTmAdH2
SRPG2YDxyDtw3CGDZdp6VSd6LC/HSJfStiXGI10T6RBslVssZatwxhM+fZ36uGmxU0YxmWaY+Ott
LHf5Pr5CDZ6vHTr/GNGOaC232wf2cYGLjZU8vfU0il5NvykpX60ms82pm17xWWMP6OgSd51/0VQi
ci2l8DiIbnKizOhL6/FWFiRxg/fvT8Ypnesdco/d++vwiChKKp+S+FfAPk1eZlot/QVovKBzaA4n
JkoVxScBvr49jTuDh6IFkASCWlJqP0d3mBGGlT2+x3Xa1PEony+qR1duvEAG90KvtyUahoR4G7Is
lIrd+B7UAU7IzPYPlNq5admD0bghJhwgCHRIUejWTZKpqf45g/Zsy7ypgqJYHXTtEWXsrwgX+WsA
MhvwSU3VC0xQ15FVY0MnzG7N3N6T5uW2QuHB4j8HkQrUSltjCdbGBc0+G7RSQl7wW2/IybqFz828
r3vVnCFLdYdNcgV4lqyNdBsAfV46QhXvoT9NtG9V/rptgijtl5xwwiYe/J0yICJ/Zt5wW6GAvb0p
7uYrmuf6keHzahaV16GhUSKMcsNQUMQyQNuSHdVymiok3l7H35W5dZc3OIA41HLLafumOsjxgfB+
t+PH/JJSXAMB/wSJHn4stFj2GUVChUZtuRZt6Fh+uPmEVNep/qFoWSv49MToys1R4wKe46EagsFJ
LpMdNgKaxlN++ULfS0cIfey9q5gPm9hscTyo4wnT8IWTVCcug1IFdD3ilIVd1Hk2NbM5AdqVBAdS
7RS3ubvG6SAhfMPDLlHtknFtoUS4eeIaTkoGD6Sebv6VlN+v2HIgmjO8d4jdW52voW4JQ52hjWqJ
gHHBntAfLBH99RxAzUz6JNBYpSrpHQ8chuIE6HZdSqi4JHL6QLPWCxsa4G/5vOmIwmTnPN2T/gS5
Ef5sQ40anSxddICvJn4TGkPnXPtGyEGXMcrjF7WpjrnDrRb95klORyeVBBi1P0xDwJKnvT07fXDW
Qv7UJPSETJ4TdOqQxeOYQESuNKQKjdv+MUjpHboa2ZWTcvPPBF6feMHi0sobeynsIeSYIKdzCoQY
DerW96NMceUipuaL83j65ynwKEn5QUsgddXEzoVxdCLvjLKRP6ncKn7jUaYtCfEWUmVpnrTyH9Lm
X0oAXmXroR94hFcCZTBZzsqzttzl/TKIqBYI/9Uvvk/uEqn4ujol/N5v7W21rZbqQpqvlCyxQh5O
l/eDkeI4jG0SGAUQHPxA9ihwSF2pIYgDHaKKIgK/At2U6NVAL9Jtm+2KzTjVVNZ0DmmFKJ5q2QGV
rXJUCExhSEUxSNPSv9Bue+2pskz5cUWe9qOHvF8DfSkd3fVdm8rEgFPJ0z2MoUVvl6yEA/EZ/kvg
JIQpsCcBA4hVvLqgZWXOC6jxT9nvfAc/UD2T+K7bHbkO3zKgZ1YGdDai7jqbWfGhcpEnQZefF8Pz
NPl5EF7JvVg+h+0NdwKFDhlRRQJ2pfaDMcIQqm6+B3P5JZ0/Pjewb/BYWsOVket2W4LZVc2pWl+Y
pnXIYqoig9f6uN3z9gz2vllp5l2DCgC9uhRTO6g8BAH6HXTdXoa+GuthxsyYBOz9Z06ou5M3Zy2h
LewH3T9eJEcBAau8ftR7WsnTdRVbkIGgEjCcIuqEFdgni1qhvUzsyrprrH73fkMmSvF0oxulkQvh
f6NxZXKMw+b6YOcsADA18kvSq+uT7z4+tL1N6ECfulxZwzsO+9aNxKmtnwwQYFNE1sFWxP418/D3
gdfUkpJV04kqmmTk5Axo+8zzqeO1O+5EHuQ3/1s1Q3hqV1p5/1SLGfwxadRbBeY9bFopqrd34htT
Hh02HO4a6bXRAer1HWcKDNFLj5nyqeoaSR3wZ5khVv6Iep5WeHysXzLZcfBIC0Q6YahEcgI8ScVn
HkZbbCeUXp1tllRE86cMFyMY7X2dugXqYaE1IT8H7V34AjZbf2or1EhKYcTZZnaqdMjQIYIts79a
KszGxrfO+jP5ZtbOeaKebsOiBpYvqkZKqOKWa/7WjSpdeN111tSnBaUHVLNNqTITWK+enR0/opIO
dQL3G2tT1QaNU/w/1SlFsLdF5e1yoEsPhzFvj5g3EynaqJIHOuxu/8idaitdUNydsZdpAgDFQfKb
1zTIa709859zPIIrzzZHhco+F51BaQQkRW5d8nCHwvcA5yv6Ewrg1v1oBkkahbGjpBuIyGHH6dAN
YOgCHO1SsUNiZLhD33huby6ehxiT5bDcwWc/Uuc4MjvSXWO8ko2JTo/wYAfd/RR0MSlhIwBj6Cnr
mClgAI8t9pB0Ow0LFx3cfR8FIUmEEuARI/uDmVveC1KOqxaZFTVoU3brxfQ7m8I95ll3Y99aHXIY
uMps2sFYeWzgYNTira1is2xlIrWQShMW/sxFxLrE6g14q5ZM5z5YZg4/BrXvJEkC04PceOBy+3k1
mkofzMq3OgWEscC1N3hQvM+FqYLZWQdLHIEnvVLYN90iwpNcgqf/FK6X82c5gtTvbtq22QMfeswz
nZmaK422BYlWA4BKjSt1wUEx0P0gwFGzW556Plc5cdh3HxIOc99x0qB2uBH2JIZGvqQBhUz6g+n1
QJY4MhuCp3MH98IP3PusQ86XndET18uPmaVJAdoVL8ZkTmZoXmsSblYdI9GsHWU9P3MKQlwe2Vgd
LWPRHfSOLUEu6nKa6QPwnPF15fLewCjXOhbGgS2YIX3+54FmYl2pVj5lsQmkwxCpxxc/kjjNuPED
lU/KfVhyW1a63aP33FIuX8TymwMam8VM3eXJKgmGG2wuOrKVINq9eK4mGM9dCe1sfm6RfhAjzRDJ
6s0T4D6tPwq5wG/o18f4QNr3THQwPldh0sLqHItU7cRTFBmwhCKfLpZw9Gw8vpHvJmIY+44mwqrX
U+jX4vZdzX5NNGElUKEbihptjnt1BjM9JzBEofQFrTHye6WpVjdb8MIBu5U+pho6CgIfsGdMZQys
yBrK+HoOV3SomWZ4envDddmw90ZJHGBOdROtAcw6XIqx2a3CqPpfv92DgtQhUNHnr3lDnpTdVy8i
VACKjdxCqJVFqx0p5Mbpzp8k+2cEGrSjCcpTBsUe+hYDzE/rHdjC8Lt67uvVH/BYRUl07j9juCzg
jyhqdDmHC4ri9JHxNe9OnFBW7QjqVS+yMt08v/z3NWZLcNPvPhGrUrpsy3E+NmvVl4OfSbDk/aSm
BlIlHvcC9P0yVNYvkv3Y3NovOHb+tvaqzQKfwYKbwYJVHiPQyVgKVmTbtirIrsvpOsA3caYxQWsa
lnc3caGD5mjGXzKE2HVO0JTHAmDSRBT7dDmPJqoeizEtumjePHLr40DkEwFKxYZqVqiw4U/joa0y
cAwVItjlFaL6IeyqipkRdEJArhSu3G3JYEzA6RTYaxYkWYrYdZtOSd3OASJmNCmcQktF3/DsphE3
J96MlvUcWdTHLgCsTMb6vo+a4ifi/61IkDiuhuXiG+owyS6FP+7HqgVFf8J5JnYM4TKvPYEC0lTW
IDIbDYIm5BtQzAw4+RJkuxzfbv6PmVWoXbN9J9HjOXyvy+1KVf1Ea652xjRC3odxRd7V2pKU8N3k
i8PqsgzudLh+7Xo+uy9okrWUkV3ehHGV0YUFH5RRGjZldImi61j9oGRuaUzlD/BCRok7m0VO+4Ja
um3UaHsY+TU5dbkyUwNcTQDzOMZFfudMkQ/VqhS1WFstLplvwdMP8gmgbx/1bryAfOre8NmAxtM+
duF/VBmJqdX8rBhdkqoPJTGfZgv2rLMo/JfCYll1t+hvFpi62h0xatz6ZtSCTeKXMD5Z2qKzNUZq
gkWkLsqRRiKiIZgq4mfzLmurFHFF/b0v+9eOeSO4hz4WnnJnPK8bZnC2WEt4LXhj4Qh3aDDPklBT
7plVOEeYcPH6mPZAiSznEiTlbCFQRwTSz9McEivXDuurEoWsO8Z1kzWdA6qHi/Gkyzbpymap5pO0
ghhoMzHdbOLlQIIZdPmpJcqy/ptj5Elny3HIw5vXs8pAeUTLp3iaBWGBlFtgEieX7s8gHGlaGOQv
EFW5n4HsvFFfg35M0uOabrIW9DIbzp8ZcquAqX5Z+4J1OPgHDgd7+o7ZbVQNYhQkfaJLdfhd8dYr
ejto3C4Id868v5G01yoNebSnlBg3FEqKR2kyUSd7VJk4XN6BbV25oKW/U6GCID0jLOJIsT++xvHE
fX57QygVZd7k0izqUkthjts7/SxI8IXzKJOhS5jR2qJDH0EwAXzPH3naS5jMwVg026uUJjW/BEXp
rKaR91oSKJgT/p3LIu9gHkpc8yD1ctLJSxwbFfwnIEU5mtubmnOd9o7PpB+Fp1rdD7NzcLL0MyEy
/tCDM6UsZGzVPZ+xh5Rji/qvHWDnVFr4yIJBKhVxXjZrkfukDIjQSDruWqLeOp5ASU70x5cSuQn8
RaA5zpdJdGjA+Er/Zs7yrh6eh9MGhlRmbYvXPlFa2pUntg6CSMRk2B4WpNJOsfcEwIYpbXV26OxM
WRCEDMZFpFYw/4e7g1onNrGnFJSVAoycOHD3yzpWZa4nHMSOMnwbEFNU2lgnCKyU3lRyqbLHHPE0
C3o9SuyEFqkwtjT1EtRdIfvYpdWR+KV+fhYvsYm7URww6go4D53ap66Ivl+FukxOwGHI9Nbmp7xF
zeCk1OUicduI+MTPf3N8fX0Q76jgfPwvIvBOJfEz0kdu2+BbbXO4PhEYO+WtdHYZKdMmPYw+GBo3
E2p+5JG9j7UmywDz1DRAfFOOzCWvov7e+5jAW27oIc+SGHx7t+zIcmyBDvDv5pyLcBZ/aJkaH348
2MFE6OG0MzOPIGjuCPdMLKbrXbOtOCwxUJ28or08+4vmo+RmHvqiOjZxox96VDZvMthJuyJti9Hd
MpcIsmyFhJm854jewJYlCt5qHcR7U3NhEJywHFXweNzSCb4Fc4XHj9KMTyZ5WFC0XpdIA2Tacx+t
ZOXVmOwSsc962kxWvM3qctUY7mXu7IXFLC5d7s46PZnXSrrk33pbuYXyNV1WpbUDOBDC+lNywYAe
SDvHEfgPzCNO6ZnAHSxlv3rFBoK8qGPsvPvITojI7IWhN3yBj7mUywC2vDxOn+ExBo8Pd5+ixNXC
eq5IhUDuuZ0Qj04TdxQV4MwKapKlfah5iKpPP1gqdnk7uEeM5Vx+TTggBc73B5qa1JTGyO6xofRi
Q6UF+8Wib9UE6LPfmX/4NZGUgvoxnO5+gL+BzbkTFE426DjfJRyerJ6K4XiShpc6U4fxDylVzcgf
b2KpoVhD3ZTc2v8uV04imUciJkD1bn7vwboHYEKU2ChRWYuAYh9WW9Yq9pountAKuTkDpzTksCND
BcwwIPlR33e1GJjEbStmiQY8YsC7l+gFth1JNdRO6p29JhkZMRUrdXmD5MVKM2NdZocdJ4agnBk9
iiAKqdE15vgSrQ91G3tQpsK9m5vYbOnJGHfS41L6o5+aa/DAAugwYWXltzZ6AFIMzURgaYcTXqI2
wWwsnriJtnfKXfo9Gc1AvhTY2/oeC3wjOLsCXQld4ciKRZ1HDfv8ZP3g0g8zeP5XIdIs8+l/MY5k
Qq4VuTCFNKpoKxGCXDtEafOXqN5hjpL/SPNvw/kJuX84OxMA8m3mhMICRdx4EWl2janh+/r3WJWy
P0HDJOQo7pGnlv6RkzSz5LJQm+7RJvh7u/Jr9KQg4iwwXvkLGagcm8xg60TRLcL14ClJG0gKxuBT
YvL3GLEmuwdwKjtn46dKzVaK80QlthTh/FvGznaemnk7/Sw1WkcMWSq2mvvvk0G3L14b43PyLASX
QMjJ2YWj5IDoAGjK6DvC1HUty71PoyQ/yffZXwpCKPlztUMhw7b5wiK9BGWdUqp4NehHamOfDY85
QgQa1NaNVc1bmZHbj5zLzWROCzbvhb7DPa+a64zXkLFxlYWk2Scy716BDYC0duRc0xtqkXtN1h39
Pg2A+mXuwBQ7on9+11pcSN2RdoTQ0KZkwHGO7n8+sXM3HnNjqgYY8IsCMpmvDkXWdiA34bLhfLfy
JD1/eAf0Flc0nerWS0CIgL/xUE3GzDYNSpukZSY48T4xMzo3otix4gfDJcR6KkJwTRu2OOdS159D
b2eux0vLrsaOsuyyGN7IrNVmrQAHmY1jWsLH1NM3ugesXUC2YivC+uwKd37OuqSsYsYCqCJj0QFO
AJRE9BtEmACRGyaOeoFN3wXMIu8hhqPKbGORHuaEkS4mMIGlAftZjZs7QXzLRkINLxWZCnVg8CmB
wDyHn0XKha0Ai3b3sGHkTY44N48EupCq3aKutAOCvJTtVcb9vr+mR8nVzLTjpjtbB0WRSPvskCUU
K6s3383n5AZLP0GlWXirZ+URTHDwp+F7UxkdyIwxpoWKpbboo9q3FVPFhB9X45staZejbEosxktC
whpMiIDSrCXK6nkAPQf+eO2QOFgky2nLH2RozI6vNluxsel2a75hc6vDPFgBYiHiX0b/nc33mvQ4
lsuT5jCbe+6ZoH+PGFnPFDTAdnQGcPdw3eOEusYc7dXb7qxShT1XGR5yqrewmpa4T0+QaQr4VU9g
y2izM0nGSdKp0HY6HUh30UuPNzHJ1SGOBzR7U3qSS/nj1ILnJcizXL8BwKVSD5LB0qEGrD3f4G3Y
jHQxm1C/8qlKZl+S7VjQB2gXUNhxNTb/QF8JiU9CNKA+rh5LL6OCA0qkI+THa0hrPQ6PF89hE6TV
ybBUZ0xaj5rMLpHG8AhS+hOIWdqWN7waJZMo2xjaTx1iAZbd5ANWdXH860WawWC5X9W5WBhCyItb
55xtknA1jI7AIkipaMn08pHQzfT6Aco5T4sn202GPzeE5EyL6JA9TM+ndHfxug2ZJgw8XjIIhxGt
5hZ7XSyOKbfHOfTIrigJBd4MOE8pv/zJOmzaF4uhfrwr5NTglQqB1kiQgMtppJj9C/WCM7n9lCY1
AzVPxq1cGOAqRWxbe39f5ctEgXxpszkHMhumz6dL/szP5LpE5iXCsA5iTdw3aqV8xBc46/RBEleP
riqWxjw84GgiJnYRWhixrL8kWTVXSvnh424x2X/SAaCc1OvVHy4d4QKDJ4K6UCbVUkYOyWWN9h9L
5oHP9xuvqvXpsIKN+U7svLSaZ3TpaqcMYzWQyfqtC+77KM2w0BHwvD/JbVv7qK/9kuUYB8PLwDSF
GzjO+GAR7Gr9p5qFR6qHeO1r5QT9vlKJbekyHla7mwaYGJUHTNsGGwHD9A+v/T7B7hy+yLJNsop1
Bw0F+ftnMeq87YbrhLzzpx6CnCuowdcr9LDffACW8sExf+qRjy+ZW0+wfzSYuD3TNksiCiecLk5C
TLbNyMz6KSXiHqWWSFqKS+5010c1gGJ7jhVImj+LZbFdKelLJxufk9EOJXU7k0bUJLLenU5MVv10
Hq42SwV/N+FIUAsPdHGYoMaY1OFCGOtG9mtJL9eXnu9lLbTUpcq+PBEuQ8XKaKlZ/ZHnIbALJMvU
QuvYQWVONHyIqzzQBW5gKR0MaNloArT6lmtPMPkLGLrJQbGm+WzzMI1KvcIgLpa8BsCsfRj5U/aa
gar8tYlQYjpASQIRTNXaZI93dyDWV1RYmlPg5tb+q0Vd5cBc4JZqAw7nytzuZHUboiq846xenf/e
gFD6TNuoRn1CW4et07mMMoxFI6YJ/O5lWBuRbS/fJRIdUV+I7T63sa2EsmL4RPhkuBxEHCLfno2j
i3OCz1tBRuQfUu4XD0TJGV3yHeq7DfbOtGUfQkRc3p8ZSFklWtfN2Vck0zME0Octau0XX8xZhlyI
YsAlv3qYCXQ07+mmFLXxGfROgSKIa7IZtCv++/IpQgQydJhB62rfrjLkxNb/u4rAdHLBowLed5CU
Bv9pertNfCa1ew0JIl9g6bC0bp0n8EJaV11uePFnaDRRBsg3C+UidiOlyJkioxl1W557BzaIGAw/
X5Wjc7VVIp6HTbOUHapKF8hamOf6xqgfsK/KkNGXBxl9khqtY+d82otBuIVOKT0LJe2ft0y0QO6J
jD5Qk6GpPQEZEUarcv1I3xLSteLrLAWsz0Ni9ZdGvWGx4TZEzcORDkQdV22zs9/KsTMAWgQ0RBVJ
7/yF2L8wh/VKY/optisE3sCv7Hhe9sykFol+gdf/Kyh6MoaKkMQXnP6rDD3ka4tgWXoV6bDrakE9
ZhGrTfZVMccbdcu8ndMUuqo1AVl9Eos99N3TIKkHea4BWjry9U5iQ+qJqC412IGt6WwxDCdy2K0p
Lm/IwUMdb0zl1EVlQKcna9vWJt+1Dnk5Rf5T5ZBfNNcM9ZwubKKujZMYEuEs4cRLq28GxErVU6gn
WsoPfhqM00NsY6RPAAgNVn6VM6ukRJrh45JPm1t+cZi6HveHXKCv3mE1ePv6IP+9WNsbdCAfwppK
kOYU7iV2lRmS0X1DKcygH/mxDwnXlmWRACrSNERuMRaP8RX3fmuw87Ylna50hMP7F+cBTwVfwjBF
onGapjaDq9zSEMOY/gITqDhe3KO5bcNv9T25VWjsIICGuLMqLItfkfZT5lMzlOs+zoVMzYJKF9nr
UdNfWCZexO2zCnqN7UMO5Yb61mh9H2wApNnYbos0lBANy6Ckj9jGwBJIX3m1xgfyeSATxt/DX+Dm
6Q8VE2kRjxH+qACm7+IFlStglnskm9bTyMCK5blQoooTsdh/C0LkoF7RLuMSACf18yUfcY3pARTT
7aDvvLLPgUDjjSoiQf3p927IWdbTDJKwN011w4IFG2ebvySxB/fnX/gDlKVocYzvOyYEJ8ewtaao
20QgnyNIjZLdnGipn/qexbW87UR0z/4uwQ9buKFSD7KP+/Jsvuz35dY83BhrnM1mudd4URUExJu1
8SrsEh+N9pqV4FeWNcMCWQSAaSkmsxP9LYlXUNEug7QlHDyf2VzTNcSlV+eCqQgfhs8crm77IwVN
99w05jCG7a1r0Qm4U5IZ6SLh2IWfoD0tE57WmEhQZuyYUd8F1MaCBDa7XFUfy7+ngV0SVojP3/Hp
xtifuVAoUmRnsf4b0shsorOKrQ1u6G16HgGoN8tzhZfy8LOZeivW/3PWaUSSsJxlQXOAX+CJVPIh
HF5Rs8ZOd2hBeuM1a7UW0DJf7yWVKFaYTTOOIaSzabqjfvQ89gkSxfqmJ1ExELGhZ/EVzplSwcM4
Bz2pSvR/Sspzbn16Hdiq2CuOU7bkxCXm286WCLT1PW9IUYszO86xf6Ow7yiZOdQA52Va/c/1+AUa
LXl7obbZCfHEDcBcX0s1+28Tp/uev2CFXfYVXDxAaR+hIQ8BuPcZdEHQoB1D+72nLN4+PHWRMJGe
Ud4hBoCW0mI0sywOapQSNCr4QosMjqjoR2YsHYjR+FD99ZyWs8f74uLnAtN6qF92MLd1cy2JLRds
wbj+CIpKE7Ys8Vt4XooCp83lbugqnhUwTjc9kRUtPotGMUs387eqCQ74zYhePTZE9ychHydE3rD2
p3sJlyjZG8YEkhcKLrv6mucQcXVz3faQqQznNNNzr7BIjixnUMsBdXdu2awNiBzRCKLg54p74nll
V3cUfgAAEgCTu8KONAJEssogmsPqh9KCQ99zQKl81exEt+Wc+BJvbwx18l2wmMYcRk9mWXpDx7hn
BtaPBKCPvaoFp6K0/MbezW7tDVRSgFd5BRr3EfsM4rba/OkfD597m7mWOdih0Aj8NP1/UvsRzr8z
s4ixiJMeiHwhUGM6cxnBf6gX8hg228nbsazVZWacbbA4AxQHP0/C6g6Y7XfS+vsCxUFEiVmDTKzb
Tg/y8c7boSskNARVloBxI8VZspPlrEk7GraERZ5np2vduO5+BorlHLKGJ9m/YTG1nerZCYNqyYl3
piPQS9TnmVeu6FFo+Volv/Utwi983FzSlq9/m6l2ln/pXLt89WJGOBDZ+M6/1OGoaHVoTmn4LkJZ
3VpNcVJDmwYzv/rLh8oXgAat6tp4q7hPBXF8Z92LFfKSy1/zsmGgVfrr7Na7aKFneZphX6GFhyqo
9sPRE6ypx7m9wggCCvvOHh0pAJBz2RKBeSG/wHEOYcmdPgro+THF6nM2WJPMn3IPRuoXVNt9v0gU
N7FT7h/weIoNV7zhSB9nc0R+ndSdenjOH8CtBVPr3p1i7EsiwswgaHeHUpsOJJZURjKL0ZRHsO50
dWsh0M/rU+HwMog9bh9LKQtzd0VqCQP4XtZ5yUR3lYkDlyfIwBP/QUVMep+wfLhXQtsnEsahuqVM
e8Mw1262LyBzQ5tpVOlwVCNmb9pzsZYoIv40smGEcIF5dQ8o/2+rqAiTMvXKGu+J9JtvEsTsDuML
CF1//CBx27ZNcfiKrHR6gvPUuDZsQvDfkhsS3T7IxzFb8xIADtqFlRE6Z38IoZ/X4D8xfh15alAo
E00e2rPIMZ4VcPkYOyY0TUBtunXHjn/3ZkDR/ysYbpYI06uutzOLNUKPASnhDGnmueNiN1vUEEgl
dq6CQhNc3GhsLPhTNGuLXDodatTp3PKFT03LUTUqaysBNkmakM8P1KWOBrZUQKT6gpw0jidvGqR+
DWzpGExw8+FV0LGvAp9lzmVsd3vlrB54256iaYDoAOZDDgwTIM07hnvkoscEvVuBiI8t6ThA3Kxp
tAPTWN3oZX4cjdeWmwcNrl6TQkn/1PbWPLp4xkvGdVQ+2SCOqZHx4UPJpGu9skrqWXYx4x8NLEfD
iiSN7XH4SWxZchMahgyBPEWNTgpD1Xbt+RZQFQsCWcsQBLTnobbM1nXNnOIuyYb+97f3Ultxsdxc
CZhr4O6W8gLuF1KIRehsNJscbvY5vjJFaGuS+lgUwgxS4QhOjfMAZ5JjSop0V7RQHayRlknFB+z6
wSUnK5oRT5C8Udk80hu2uyNtaX3wkYHu0pRBJSowjKJ7EteqndkCZSS3njpxqwjpsZ2ZB7z8hVZ5
L+wkVqzVhtRbAEuOt3wSWq17HKUozpIitA+71OrdIY7+chNUYiUxR0Q93zCcKFpq+JAjBD7LJVTc
itHiITYn/fwQ8tQVLMue1/i4WZXdutR9BFXn+E7XY7jYcpVv6iWC4q4aHEHTbzGz4CEtrVHaJeyp
+hZSCQnS/McdxYl4EG+Wa8M9/+9QtrNaePN22VG7y2+pY3Nf8rFU9wCu634sRhwedixZEKzg4fPB
UlM38meb5g28icMMPenvvUh/qlIcypJDNPyyztfHGAOL0xkZmRn8HaAmsfx3dv9heveuBdVWr1DZ
qYIUdvF1/QWjp0cdVLD91RnLPLB5N2vqKQAyOxIduIhU/01OYrLBODGzoIicu/14IQhACkc19ltU
nRbYzDAK3I9errgSkGqFP3af9tW+y05YGFEh3u2zHBxO60V9V1nbpTH+e/3ChyEDhchzBzjH5h8B
7PHoNhkI7cEBIZFzgPiZ3aIm9RineJV9S0Uu8te6BpHp54chACLIPsSKyHUAxXf583CccY2ZCfnn
n3qYWipkEY7qrCXK42fji+2v7eAJZMk5DJImuRoDyqAdRzpfVM+OWvlvUUWFMDqEst3ursmz0MTX
b8i98hGQdTBr7TZ7dQ6ErvK9JqaFLgSQzqO34iO1+NOsqMHAAEveYBTc3I00eWPok20VdamgJrQJ
6b/xyy+hzD9zyAjmap6UaV+D6Hc1sGUnE76dqo4pp7loJK4thwu7LRGQaq8CLdPESzaOvI12dK0j
S5b7lbqE6gGbof6lBu4WW8cvgHmexRJaS6H35BTxSG8Hf+Z9RPkphCywsjqjFe+DAR9VT/ZrcWm0
hmuw/LX7o0ZFT145MTX45pvdGL57PplxG56Y8ckyzngqK9oRaQfANkt9k+A3sONpmZaAgnrYZfv4
prVtZ7ddNWyBwUlUyAiO29Icv6OO671w7V87Mgk6mWYMAUX/hC3tqW7v88GYc7bUd4ydWaFy8RmL
YzbaeU0ECNLmroNjdjTSzdcjwTAUJa62o0yvxKL8Nr7dfb60IxFfv4ta1G2fMUQYD38v+O4IDlL5
W9BJfFZ1ikoyKAsj0Dt+yl03FcVG3twIRrNS35762hEIrs5X6VnewYLM7NowiD+BqsCkAhSg8O/G
cOQQvd48wV8N6EPW6725zLBIwboA4qoBD3z+CtiVsXwzHVPRpUnioRajS85zUp32BI+aO185ydAy
v1TkTAcK5Vj2FtYaikpqmWaQWOgaJ/Pft7SkFzOPX+Ei/n00FZdrm6vq+7BFdIOqgZ/8ck88UmbA
LwPd/JE7AfknsiKiHHsh9wKYX3XfWEa9+Y5xDSPIGYcUXSf3KyxioCGyOO50omcn9pamckcwiZOp
ogQKCUn3rnieyMfTIG+boyKkNFIUqlyKeSIOW9oNryCPYJgVkOSYRhtatLQqf0bZdZW/74MoT+Xu
FFLRe3wH4Y69Dso6p974idUOPIWiDhrWOURiIjuZGxugWSeWa8MMve8NDRMPPGZdUX+Jlcv/jsxN
GN8Xw5CX79Lt4W3EdkLFrCG4LFzAuPDrwra/4TY5QlqTkefdaWy5IWxMBUYEi8bjixSlnYp4v/P3
DBUDdHwY5QOWsnywznGUTn6QaCjiOMYcyFDmQEL7hckU+L9+WxAP6/IXfFTEX0onCsP/7r2Hx8G0
iaWoFAy2N2GhUOyVVFrI/Pcxh0MH7GCR/siknk/eXw+6tvKiHWgXESE8aQEyyS0sbBucY3wIyJio
//yv8cA537B2IuofwA2EzagkBGl81HL+No2Nng6T2i7L2YYWfNnj+ULcm09PHfonnqYWxGfhuvAF
kjgwfGpMHNg6hSOksbYIwjadrmNwXzWTiEFJtFVuApHZCLVDP5lGU0YGJyQBE2z6jVZArpwtX7AX
PG5ykSYBm76J6NQD6ewtELBBJ74BZ3aAVZE30c0OEC6/YiTZ5Zb0eXeDu/jETv+jRjcyQGuCnQrs
8TV9jEJkVBDDMFyUk7/JKB710mNoRWpa03ROj3oTePYKqDgnp9yeXTRVSBCi7ApGRcP6koSOSmfF
FjYpfaxwVTZ7r0/8nxYbQd0o91cRyUMZmdi3jORhGpAzQH3TYXICHdMEd48HEbA4/IqUho+jAuGU
VNMr+opo1JWKZ0yH2o98bobuBInYdJXyCbBvozp9TEz8HdoKEj9oKGbzkPjdIYi8NtVDVZ/np/Cm
/Xyl8/an9daxlS0Wu0JllutC5enoBAdEMgtWvyRAMc9AgFgyB0f0JmtmvLfGNdrJqMYDyJoVWhcv
S5o3DgPpzxYKe+2oSB8T7PMfKBgp0ha0n/O5bsQunpuR0mvYU5/hzTIWuT7wGhWSox3S3j+IB6Ws
6Dw9ArCPUhlCCaW0Ks8r68o25RULA9rcISYlVD3IOmXzmavlR+EOmH1S+KQhyumFXZWX7jbFuCZh
1K9u8fLwDyj6Y/hW9pLojorHtd9EjtD/eZvQUZBCCXY0GhkZh6YMoV/4uLPFoSThVL0YPZ/OjQZ6
IjGUX8agmRJt/uH2bwf9EtQODtrrSazEiIShrMzIO7vqyty9a+fS06bhwZJJVO3JvssR5R6nRM5h
MaklxjOWnkY5Pyb5+euT0sPfPn2LUzfKuiqU7ZtoRsFs5oraRsJlnCKaaOJZuDoJJmZS9rUggGMp
F+J0+BC/hVS5uvrDxDgXYRCEXFcK8xI5Rcb2IRnom2yxJkCwFxlDwbZfZqJWQm4RU9ltcbsNqmv5
LqalqEtKxLyFfFXx2JIHCPQ6Qtp3FKTNqwbXHupVoZCj2YNEykXrSJzjU1DOK4oLOz1Ao7suJ21t
VHm9rPQwmTJnL9IK4TDCVmRAG9vOelErY6rTwvdikFLfGREHuoaQPGwa6WNGL6g0Mx0Uq7Wr8KeZ
c9uMnMCtvALRSdpftM+1WcI+p6chy54tBGKXLrQr6MOPrh09FURVW0Cj9GOEhw7A4yqTGwQFl+LN
TXai5xSDG4i/XRiXTZWhUydKYHRxmImld+Zq2qkKXVfcG4qX04GHjlSk40b/vaJy/dI5p5FBUhe6
NygII4r5HK1g6H2r8Bk7cR7R4YsOFfPlya7Mt34QYkci6v8tDR5MyFafKTbe29QKo22d1frCHz/j
YeoXiZqvAdwCC5kMP54uMUwmCNlWEA48u79y+yEDdWUlY5/hQnP4dX0eypJDWEBLdCM9ttmGfJES
I3ntYf28Aa4k9tJOPBELm5URNzZmAd1u5KPpVmxHsor44vgS3zegOilo5AS9qTxZEwYxSZ0kLeAx
8jfNxFodhk7Zs7nG040l47S8FF4KyBIXMpjW4LY0xTyf6G+sUqb5SNdlJMxSvoW8X4//9Cq+HiEP
cS6D9wr8pD3eMYK0ztnK1eiNLAOZkBHIDd6+nt3f0lZ4LByTOuqZou8zJG2im/c5q0VdYcDV4apZ
oh6CpFZKCghb2Sz6Smgz+p5lQtn8hOOC82Kr5q+qhNMtaeP1zVnbYO6kUD3q0l/azfm7uKQ19x/V
3AggflHszjUyy1lMb2V9wv81V1n1Ad2nrgyd9ySRUO0MCNC1lFs/9A1awKYw+9bnVrg/2ewWHN5H
hj0NRDtiP/gUtKdsA34JreUtHKqyxCx1xr6wD3fYNDNJWwMKs/fxVEGy7lb5x96g3ARdMVRrEn1B
FMTV+X6iH1t/sgvfX0t31pGpSC/KTcS8fey1hw9Ywu2A9r5zYRUW/S6POv9HpaTSSvv5aXPqOSVU
UWEJza22QPCHZTYDkhECUr1FnTSi7Oozfv3in9IyjjOrxQVtS5qAYgzBKwW2zPiMSr0FWqI1j2T9
6jH1rjvsGG135yVxJIJlqZ2JbNSVlJK+M985dx3HwfIGIJkwwWYjLc6CaLGka4TRj5xrRISFKQQz
RDWXTAN6VpMBvArKZvBt/fwj4CmnBb38OO4lehA0kfAUqb2Yv0xtEqFedu0BJVWxNxlW7RdCWwHb
49OBfM5Phv0GX6IDTjxH4cLTuTinuGK1LPbrQquH2mpkfgm7WSwGar4hEIyuUs2/ln8IWareOQyP
OKFdudtzCnaeY5vpn5fXI5/SsxZg0m1/rx91MXLu4IycxWdDE7woBtYMwecv1oCLY0hLqzmZzUHq
qsA0j+j4HpwDugk3CwzPcke/PAG7jyIQyM0pB7PhOfkH1FS4nDA34Z1ridkp/T4DsefKzTLtgNzs
HBskLv4cYj62IAYHefDNQJOCwGEUrF9m8AG1CzkHVPH3zrlCec90LINSdv2pdWlMziGN+vBg9wz9
F9rSbiZtq9QxfSscGzc+slJl5xixhqyvK+Ki/mKN9dB71r+UJYzm5IFZw2gB4C38qZ33b5YJQjaR
ubyMGHfQaZz0LnyUpPFNYNy0hY5wqccnHmXUt3U2fZFk91qAqYBJ3cfz6/zY2O8CtzBeNAWHP3iE
LAi4VEIsWL9vHtKHEk1AZebQ06rLbeKZf7LUDM4joOT6cI8w4IN4w5D1J1FtLuR/EsDDJ2DpoLQp
h0m746iA76geykODPzX7l7uJ7i10pCXmyg38fHtk6X0Hx0eEOm4/1SeIV1EDvlq8ng0SmIiVmBbb
OVu09QnpkK3Elsr2QcTmRpo7ibfThKIJL2/0G8ZT5HXPUKJVj+TOCyAHagvLY2xKKoilhjdsWuLu
gZ8Izfy4SAyrnxzQ0LjCwEf1ZA6z7aLF3ycV2/uB5szpEDwxaZ+TYFK0U6PiTN/W3YEcIC4w/pB6
lEnu/aLrevuNqsMqaZcPMEui4WHbua6/bBsohL5uR79Ftg3uEG/w+F2Wqo4Dgvf2XchTa5OuQkLk
kkeOGQzdPSWK2oRUuY2JZZDRsBg2T7Wdn+tJ/sQRTZramDRLVjPKJ4lEYvtA3mO1qYy1QlYQ0tHI
t3vKsB6P0BhbBzL6vOozM7FPFP7y88mzUHRJYI+t33iMTE1Jy36Mft/pEaFkmL90KCDbPgkOSjn7
+itp8ay7Piv6Mu+mwYaL7pp+F1Q9VeIVQRV+jGAwOnhfKsdPHCWc/1hEPS0xW8mFmvDXmq5H4gxt
zLLOTpzQCZajIBwm7f+eLeJcEyCvyGs3DL6gQwdCoEYHlhZVsvoiAqYL2eHczSDo8fpXjoucq9oQ
wNc0sRArHF9lx4nBog2gTUrwfJq8itsIy+vIvZ0okB74dWS2ZkRH8CJ8cr5HH8MeGeYP93u+XDAh
cFXqde32S8u7l2+clRCubqYSc610si2QVV9oKdsU6zOX/+F3d5bx6M8Vh8HYSryNKTgkMwCPG6XC
9whdgeAKBNR1z6BPSm+qN4bfK9aE1lBnmaHYV3tgHKyqrehO6bi3bGZB+FIUKEbN+5zQ9qmJVmZw
v6wwgwuH6p3ZNKAxKVbTVxGbgEjTTplcQ+25UjyrwEYxTk+S2uu/rlyfDwyEpMr47/hWbbjqK52W
DQjUPvBt1VXNCunHCj/NlQkDw+CT0qSm5OdZV/YKwxFajAnonOam2eV0OKVw82kzUUjCGSzv2dGU
PvaYy9b3UVTkRlT/YUL8+1z+RYtr2CpMp+gIxG1SPtE7YN0uD6DgF0k6SAWQtxIpDUDaZ506wMqv
mPz4ao/4iSU7JHFqJKqf2y6FUh1iG2lPbL6Gt4r5xVxE6Tf65yy1cTFOrvIeUWFV/U51mQVXVFD0
XqT42Is3UZk8wEGWUWUng8mYqz02HFi6xP6ewyc5y258CK+yyk7LB8hwa7JCxFaJERH8nlLhBLUa
b+siYqXVxwRR6dJBhHPxFfQjIgMmyt1M2MmunYmPncpMDnnu9hO/eEwUGAfVCdICNl5m/vfgSRJK
CZl6zIcHWnmG3ZelbBHORIn9t/PQBzvBkKBmOoVxB4RVqPI1ycQ5bhUaDfh/o2I5aRVWh2efxPGB
NyODmIHAHLpcrCke3ZKWKvx/Px+7bKVUtXqnl/qsPMx+HBrPO0JU0LEKV1c2REEcQhEqcKcxQ8VQ
IpMIIkkzgvjGKHUkBHoz9seX+MrjghHTc6sunElxlI8C9/PPxoXWuG532aGxtewu9SNrDckNS0c0
8qFhyBLbfm1FjWQ0MDwD0BCvBSXhavJ0/Y/0zXa016EKu8kZIBjz3Y6+G8OEhGSnJy5BkxGdmf8o
88PUutjY0VA6TGuk2ye1Ml5wgJ/OoLTWY0WhzLdpeCbUTNrZigEBFxkA4jTT9xGsLrUe3rfpKbqR
wpy8V1lxv2Kg8rqG1ZNJ9I46nMQbBm/4/BEHZwgrvjIQ/EGbRneHAQ2ceeEe7fZPR2LLizM6nCAg
UAo5q7ptcK5w7+bzCyNqGaR2YHzxOtxxJasVdmuaMVGUi5v7U+2qG/nxgw/42Nn6+De4KpNhcJDU
12e13jPZhguU2slt8mozql6uhHzvpBsXVU+PndbAV7ofle+BV0Bnq2WLb9rbvlzjHEB4IbaAxWLc
dGsG88se5FmTCSho6BDdN7l70bk5YuvwW/z9IqlCYUUep/5gJXCYeO/m4f/CtuibBAK+Rfb62K/w
ghlX0Ix9y7BSiAkfPLl1nivRdGTmtJNqBVP3WdpbII/alOKcE//9ds/KJf/4PJO+kCOR9+UsZMdE
T1nONDczJSHrd9aSS0IRacZUV1s3lnbjR4oM9pKyzdWOimD2iQF0S//lvJ1h6jIWgYnTZ0f0eWqa
X6Kqox/dJExj0k7e5KcgTj+JYE83Ydm9otwrIBRQyIkR0iS1fQ/LULnpQEbljg12MErvN6CvSqbw
PGiPyXEYGEFd5OgWIvYmQSXXW5jnY1eyiUsK443crqxSzmR2EGF/9aT3iiFqaGCbpSJev+ieae8Z
kqVRx7JBArWDY4obZkVklAlyLnp8wamtv+71NdbuBdQgzThBZWadlDzzJlwWXq5wtgLYma/Fc7fX
LOtXPDOGqL67fxcb1vEscjNn2BqcVwXuMS/otlmhm5JZ/6tfAYh6L4VJgLLFYydOYmnOhZItaY78
8/y/1a+FovLcnTNBMnbciCPxgHWFZXSG4xg/eQ68DGTS44ezKKR0dXwnrytQ+bzbiuE7U/8DSWnb
fVDa3u+sVo/ieXzNVCtORopBpGie2Yz3x5psMZSDwbr45ZudFrBvjEwLDdVIB16pPZT5e7dV8ocp
pwiUMa9pvBWyEGH90CtVGFFaB42YqQKyG+C3GE4dnQYmrSnShRYJCstjAuIdjdP2RKHbOMZWOf7j
fVv5nd3NaCRLkRu5f+p+W8kFc2PRToIgV3z16h0XvFHeGcWkldatKKiYVPhrFb5SvRxOUW0fs2b8
gkHqg/+DIpzx7Kew+eU7A0LUteqI49nyTvms2px2sJHGWt25/Fp7YyskSLyTgrUpm1cM4GwLawAA
Of1Aj6elhGnvpvgtGWOsZGTNUxl9p0WCKyFw84tPVoIZZlp0W/F8y+K3H+mGAN615gF6PRagjYlN
j0rpyIBPblaCVSQYvQnAbhkBpdnIomGF/ZNlUbwpndNOG/uSX+TwpPnZRxX4HecEFX4inpVEG7iG
dlZwvZWR6tJVnm9hn8loIJ03zD4Nt7y52r9aREICEiqxSJh7VloctRKS3Yn4z2qoSF63oDbiW5lJ
V6FL+VA6iy1TU9OsjI2O+RwCXExmxdLaLdhbhzcwprQwzqKnamOiFtI237zBxfgMHHrEa7SGFA4E
Itg8oc8DQhlxOOL++3b/Q0hewKGJhn2bkKnt8iLbFaRl6/2EA8qJ0DbFQJz89Au3WnATXnN880yF
gXSS+fratoIwY3x3ebbjX9CBR9A5hIFoWW2D/RKMYfLGUJuHAWEmCDk7E5Hqdgs3BRtUEnif2tyi
u8deHd25C3jlTMuQtg0GpUq76o+clV6c+z9PsZO8hnCDDFC3o4msQa8MflnWVY0ZXVSyN2z2FXh8
bt+rF6gMvi/uI35P5Vt1F6RPmyVzpLnNMXXwJLyAoUJbMZSbd21abg2nmuYo/jGKXGjqA3hVr7BJ
3DRXV0qDFM7mnJPS9Rj5Phx3PNqYJ1RemPsFNCpNhks4a0OZeEPITEwEV/RYOGuZXxkja0GK/fJI
tM5ekaKbHNBBAwuvkoCoKJuaFgZH6pgtmxm3eDYVXsF7ZL7ZxHwTQgSy9hr6+qvzdnpCJ4wo/77z
XgH0AzF/1JA/BrMErFmH80TI02uEYotj+VSntePGj2XLJeIVvQlh/aHxl+cy9J5UPs+ihYwunSTn
seqLJ3JeuYt5AKVs3qDRIJf3TCu8dcwcXhcm0cYD0yfClU9IopKGKaGSZoNIudl66YBYx6kq/8B/
9KX+jHbbkX545Ufb+sg69VRV1qoEO+Jdt6jda2bBVJ0gEceyy5kyH+mZ2n4xhVqGVRPpU33XloV6
tF+vGl135044/5kd7mAQUFfjehpWyc3Pi3J9YHPzBjXfgVOie1FNNd3zUfSowEYzgBISIfuXtQo0
peQ3EUMZS39f9xqfo63hlOqH4KYaVfY1cePvY0xEXzz9GNXoh7+Wm1iVaX49HNYMTff2QNghnYK/
14vZffA5gxZ21xaqD4LPPM1yO4zZGWy/5yn0s7+uq+coi9JRP+Sb5RpLbNHJL9gdG5yLgnP4KQXg
pdjIVaW/gudUgU3upUq/eHnd+miC0Wot3JcHancucwqWKWHktqhETG87tID00XUcLHvcfgIpDMU+
SApu5DPuS4hFpdnXJ9H9v/e9Xjy5CzykpIbKvf7wVob064IIxYsF9pukF7HCRe9iv6jEXmkH0+0N
h339VUyHcB6UOyNAFQGH2igOfTugUrw6E4ea9MujEAS/LWZ7f+WxQfXzj0VywdUmjxWbSDK07d3W
A3JwNVK0HqvJROZmXohWKPaCX8XTCkJLuvkjZQMc44NpN8/HzAGuUrQT9y99OAsW1wNIVRurMPY+
GM6WgHkwUTtAKZhlwmSRqYFBvyjufzN7nXA5GRtzRGDThj/TVcy4YtJql5z4hccHwoVgCgn3p7vM
L356gRsBjlSm4bcOhppnmn7dRPfbxpJH73r/tYMs2sF8io4zRP1yXVMf9/3u8ogm7AE5MBUN1nW9
ZyofVdoGJwlPdc6Ql6HBfa9EnUHo4D5+r9bAuFtJFkX/eEURev9OX6A6It4LseALMNVeLutcxSLL
79Yu6psRty2T/7nifcFvwhBJhI8KuSKmVCJcePxDouyHTiZKSE3f7eLmqfxlIwBT3q6YKCIFwZ0W
30U5cUbAZpDPQyTW5SZJVKrfb//Yb+gqWDxuH2fAxaX9Ouo+iLX68IOidhIvTwl/wB4Wf5ewFQcr
jd8cOAy97qGXbb7T9cdyeKZ9rtAAcetMd5bzoQlKe9zueQV3iwQ2G6TBSJA+w+MY+2giG3SnyZ0U
IwmkakziWp6+E20kfUVudsPkEMRvOUhtZ7N1X942P99Q+i6qXzMmSLcfxnC2U9x0YMDpqaniR6S8
erj2k4DvQ7jCQ+cPbocqUi5na/cUF/BdL0hdlSV0P2pIUOi+9HBRPgZ1xxEXkkWEvPjnFEnoqhs3
+4V3+wiv7YWSF7lnB1tT1/cpGk+tyVtHraN4SNkVy5URJvsCPvEtpWoL2+wr3unwVYRydHIm57i3
wed355dfh06gxn7thFH5tEnkCSsFcKD9lYgt7U12xfSkrnkVTTfU0ub57LjyrUpOg+kwDYfsVIwe
CYr+uSa0SpZ3JUsTPiJz+ELapA1ajhjZNveHsMkVAWr/JnNNMdM1iXZ3t66A3cdt7opplzZzlood
QdAAP2DnihT+y/4WIBPUQQ5MoeUKGzFNKbB1AHIhCU4W4mulktd+mNHvaig6ic0DlnHxslqZJNa8
UlbCwr+6pGQxALwwM1xXEeXzFwa6WLE9LCc4R0K1njLEjzr9eyDBiYeDtTeRq6pJ5IJ/2X6pqzcb
QcBhKy3mRYtxygXK8w2P9FDcc3+NB9qkXO7Qu183hFnLl0aZ1L9V4Fo3t+rO/gnXx/D+dEgKXqeI
tywVyTdSiH1p+9qug+kf1qrdnurKynrfxeDcfjNPFRAQ4AkaAvnI/sqTOrCyMZ2Nd/kgOqanqb2l
nrAgn62w59yIbqzHjnft0t3nNoOqF0BMWmv4DRPDyHo7Ei2yWCrWyKYhHB7C5PThehMQzsSBz8UU
1pKmIIgmxvukCotUBvljG6mE37YXYoBOeO4BkUEik4scZnOLjHycjSBrDGy3AbaHexN1HgZdhfNk
IcUN4xw6vmavvBSdZTNmv0U/tsxAyF8FED7whCGOZBM24pI74i2H6OSAf8XFlTf0DCLNcUFwrzb7
20o+OpJYcTi8yGRu9P09AlZpZDBN5v/3z/9rcNYpA29XVWTJIgqf6YWi3fESdl+QbcUvo70oNrUZ
h6qlVWyZfzhHK7o+L+5oa+9OjYEC0WE8DNvdvznmuJddLMugBLjOR5qplLCm+5ag/ozyuJ29KMlH
MBPdYz2yRxNkHRNKi+8Yu2UTH+LvZrJwFLFzc4C5uM/UjOIPeumeIs47h2hTlCvj6EhDrREnvg4m
zItyJ6slUr7d4nqz96NQotrPclxfdKZTDp0hZwzEb+jmDpX4mRqS2CNkc65NGAmYwyp0nLHiFtUC
B3728OHJ2jSrp9bKIfga6eDKE1QMcApqPFgSZbjQ3VD0Qeuxemix1mkDJSq31C1PgO8uG/1OroaT
d1/9ewXnh84BHeKxrZCDXZyk2X7jthxAItBFxLnhraaFTMhgb41rWWxRALoXxkmydstfnsFFZAIl
hTtOIP5xvUNgNC6vzmv2bK6VSHjZDOIqqBHRSkn8NDKHrqwG4ac4Ycu3btxEQkDxFCbSdoq2Eq3t
KuDYcuwXLdvl8I0H4nvtexlOWBWdnkXGWPsorJbORh0VS/AXofvuTjtVSUOeE4wxbisBilOZmXkO
SYhPm5bOQWfnr9QdLFHntDHmo+045thBSPwYAyMCTRkEVtgFNzoKPu5RZeB28e2zqRL2Pi7JQ4MK
MbL34JPX1xoaGVZcMjslBaVcOe34BL44q6GNCU7aLs9R1UDM7DIG0zBnyZY+l6Pg3zWx4ECh+tWy
fK6B2pjbTiTyAWj07V7J6JkxEM8uqPA24BS+sQmtvev/2kqQt+aXeentCwxYTYgY/bBQD2qn6DMf
1T5+pHd93HB0n6y0UJupotcEny6vpCuGqTPWYZaWvDlF+EN7DRutu+8JnxuIXuqEtqcqptx1yUJ9
GifItccAu7GG/Ogbl5wV+hKovfHIsPxmJFeOGdWb71rRfETb01pKwX0s/Qsuq91jCjXFLnIvGjub
duD4UpFX1M1qIjp8g5G+O7iihkqnUqPp8AZRSh0kOMNbCS6Z7I6X4ChWr0gJPfMyJQY2M2kZ7Dom
2oSh+999umQ93MCPU8zBUlnuN0MULgpsP/dEW/FXn/a6kO/Ti/nDLZfjP2KOPctmI+1koZmZmmBL
D2LhDUVGcEhGtdk6IIO1Kt+z+ynwvtbjtj23x95HB3zyEKyt5NJgKUj3BQXs544Mi9rIVV2ueuWI
qsGnYeE8w8VyC4YQ0J5o5VdoBqb6UP8ylUWIn4q5CBjViMtXxq9tVATcOpZHFUXvWVebC6AnHVqo
qqlUtyjQK14XysQaKxfTnY6FKXbrJmiGEAWDRHjueCVS90+pbAg7GC8XKRETuf9C/RBkWcyHmK3j
LzOcsWUX/DG6VBkF7Dv9NlATn+hN6UXgCQ5Vre735qV8QzFCoeohPYk1BMznBcgxmZpBbzybZps9
nogrbN6o+Rfq2s4IIeGnZbp+20Dyf/ZcdNROpbiqfl+nh1bnUFSFMOlxfanaAQSMGHllqh1tiueT
IOhSpeF380wNxXx9WLgCtLhd2W89hhHp35g1uzovm29/N/KD4n/jPQN2QM5i97GXsm0Pkwl8D3dY
9oe2P9CsZ6kZDBO3oz4lheEHUu3S6u4risdLjN2gdnMMWjo3jEiZSIvWJL0kwcLGHc7Op2MediZv
mLCedJUyr9cAywhM5lDKobcZJlOM4MO4pd2fB+8ZeZ40KfmXov7sh1Mmc2TZ0FGq7ndnovQ6op8L
ddSzWKfEy3QmMMotAl3JoVVNxsE3gDIoSHZiCE0n8J4wq966G3WsPuNVecN0oQTyxZL+VH9ztZIB
iHZPO8FX0+PZ3xIDjHzJHu/dM9dVxbnAkbUfCuP6Jr5K/ZMhcLnOFNtfW1viX6bYgLvpenVG79sS
p0hQWT2fZT7wkyzXzi6lDnBIcyRvaVGL2NV2rM7hWEkLcVXew6VfWahEkCzqSJoiWndQE8/HMdER
PEN9PnR3LQr0dLfdXwnqrnLOTFMdyygjS4awacvxwxo9hDCO7AGUimFYYLO35bvXbyoLDy+5BuhK
Ae6+nl5TKMa2DvKaQ1EVqKX0/8XAdVxgspFYujqlVKkEvqrXmd81KIedFUMeyyQRXY8mr+3o1Eq1
wnRRH3B9rU/MAur4CP1OOelk6acndO+STN3BHBKDCWgqZEDV15v2jhTHG6lLvMqPQbditeHt1wgp
WNHtgweAHvAhUjVP0V/Pg/rwajDk45vX12HyLAedngnDx8pL7AapRpXVgLvP1pN+ZnWhJvHl1sZR
RI0U3HdO0k4CUHtY9yQ/gzy3WVb8TtaHDHb9uN6JZb+2MI6EsfU0J5PFjMQpTSfH22i2PCTUYSzR
uKIfr4yP/kLReXAeECA+ZUk/XtKg58cOOkN4lf9BglomKd78vlcFaHfaHuWHLmchQ2RdcBx8OJvX
HLX275nyHm/arRTuamqvBLIUgLM8MZyCpePeyjxjqj87eB2RvAj4GfsIFaWQrvdemxpIhmaCngPj
MrjCnpmR2Gz9ImU+e2kjT9TVZo7bE3IHUU0BTyts4EO8meDhbNrJmlZOuQBi5e2Q1AK6LvNwW/9e
Bx0RSrvLXfIQtFga1bH5dfe/jNN9NxkIF37SPdpJRePHLffoEfbo1CnL7jXh+GDuKNOgli6nvbsJ
YNKwG7PpHXnqyb/9Y98mlImJLND9s8CLhtjWzfqPQoH+DJaqqFCkXG0HyH7ZL87Ndm1z9jEHGrcB
AhAsvHL91KZsljzQDs4+GwTtUudt7SvsP9JoDFPbHkC06MdvzZIklBED0K9eB/iT1dpLq6N8pq4e
hTFzrmVdDib6Ir/R69gbLHIdGx8FdvnZ3cYcQSaJSLyK9IgLlgkwGN4ISCaaacs/Ht/RYzSaz/qT
FN4F9lDj1VnTMR8V1OuewuANDTWJgifrvSnnIG/1PiznWzAyEAa3f0CBI4CRRnGD/PCaF2RArNSR
8DVF+A4h0WlJC8Hi2+SgZ75ypWoQNXIHJqPx8uPiGFxAwYciavxxHIwNLwb8ia+4oJ9DdgWRKBSL
Nks8sN31Xz9PJQhCqj2grxzQZBKBRugQ8l8ZJL+nbP/u4DwLxvE8zrkM5CXZqYRug5Q+0l6fYCAv
yG1/RdxhFkxCioj3yn6CzlNsIml724h4xxrpknJK8dt4W0Kin+juN1FNZnhciYQeoqXbPkUw9svh
rXoGyRRGqoCu5xCrWy3bisR6P5djuu+jADT6h9xoq0uhNpK6KmycUNF5GdgQvXlUBmN50M3HxlYt
RicUbcA1ZdKlYAGMIuo2TR02dK5lDqmhNZKUUVcpC04vkFqpFPYgdCKYtkqvQsDtTyI98a+1o+HO
FSInyMDWYhm+702dhQP1pV1DzRvQBBLW2tyzzCVJpT1vMJ2zNQazAxi9/kqRhmPnxnkyc17AynWf
/8IlIWy0XLHJtCRAv+QDUnF/3bPOveWI0kco0zht3T7552xlB2/u+hbHnMVRVizvp/9Sv3JRSW3F
63/Qolq+W+gNA1Y/fK+W0MTzaHYrvK6QiORnYiahQYsBfpmxSmYa7KzLpPbiHDpdxa/U5W0R0GDc
W4hMjALdPjkrm/JJqLHRE6DrZ9w+5vm1zaNBCFlM1KmXEM6Igd/alFh18Ouk0fpV1BnbsFea5gCb
GZmQqp1rXjIF3gJSOJAbTByi6BqpRopVdc7SA5v69QPzFSU0iZoTbIo7UEBfk6k+TMpU8plJ/Viv
lq4kQLk4gLQ8r6jN+2bq/1n1+YNVthfFQNvmGr3S4kjbcgzq+oaTn2CknTR3ORs9joFGS/lMqYRi
Ea0NxDdjtwwJGDX1WIh0daO7Cd4Mj7riejCsI73UMVfXS+PG9NWR6VApNpGQ90MV1JMioWG5BMbU
gBSh6ThvJiw0KTHz5BdwMbgJCrgSDal0GzCVJuM8lY3KEfp9isc+9M8I3n3gX/8XYEgO0+nJr1M0
CZM/WTywdP7afF2QUeVFGjZnVb+IDM5K718yASLLhCfPUCiUXoxtgyw+7jmD8p1ydqXvDC1PhNE5
zoH+GAObcQBORMIsrBVW0xyaWF7wAVPpdwrXjhErKaIW1nZ38TUxH9mH/7gQD+Ye62q409v8cowq
rO5SFOruYK/m1XuWUzQ16SoNM59eI2PT7vK+qsRcZhXAr1djGR4uUH9yvesvjNUsHo/X5ouKpzmO
gS3ir/OpV2toHM0AOeKbdzTl5mEh31+ahHkvak9Gvyr1m989AnnVIQb46j1p24MFr4do2HaxcmgQ
WDc4scYhtTu0ypxBzTrM/X67ucJo0OTACVjtWgOzuwjVQ0ohoP+mulHVWCMqDCXI5Hg88xLl+X/+
HgexTv6Uo297wMMcy/Hq2Y8abDWCdfNSAM831EefWgxBx182PDyMpeHHhwqqtYd7upQGIRQks4zo
08LTyL2N/k+35msnPPC7DuPTXtyEujPhlzL/Zi0pIr+8RpgAF4KX7BpA8GRvqusm00LUGuE+BU1n
L7X+GDvNV1flrsK/w2ijVHuTxiCxbTLiv10OBO/FetMufmcHUthg/FlQKTNMZnlf/c7tthuJNUAe
I4Lc+bN6cCoYIv7RLlL93xZz2BaRzR4hYGX59HeeLPM2PijRGyCtR0jjTmRtyje9CXQHazsAinFG
A25sehUJvfFQxCBbKuDBiKMAdb7b+MItC2QZTOvqzSvD5XzfNUEQJ6Rla+cNC08CHaP4awfesUNZ
Ko82QqU5RVXrWl2CS3qvw+2DMlWcalcmdar4g0N6zqw+SWdh8sOs1JzX/KaUNKJi4EppAaqf1cka
NMZTU5vm2wxkjNEOBjYUzFhquyiuxxbasL/WmubBLbZVM80/0myu/tdpGYUy9247IZatyambIszh
JQe2m54LWMWEXo61XBJwLUiQ4cg4bt4OYS7viNCXTpp0rAkueXjCpZO9muLjF85l0WmObkhV05MM
pixr7zpOVj7cgh1Sp5YfEOK4ts4K3t7t1vOAnmbAMepIBRBrNStAKJ50W3qqwTPQLISMMowGeSb6
JtTPdUnBNyzgJ449K+aMmpHaWf5c+Pt45/DTbLuSS/RadIEJi3odFoAXzFo05yg4ffe+HObqyImD
X7dz8JQskKb8o4xaL8VbGZ3EENhwqIZNUjTFjc1WyaYCPUg0QVyYA/E7oYiIixc2k46ivc8xYrtK
ISDScxKZfHofvABG12G6afXZyqORwqFX/L5JhFaIKeBD8zoKXgNz75ZOfCwVUQXdXD+adjPEwd/S
qIQc+iIgOTPETeYxbGPlfx4KZa5oHXLjNn/pb0mSriZrVKqh+aUrhCyP5CEAjoh6SU9g56yMLYty
dknbhdCHrtnqIkdjCPA8PHR7MdGYmWxNsjB4d6466Hsii1NHxOyWW4SpY8PBCIydsQPCVy9ToXJq
6zDRl83QQyKqqgEaLy9y6QYVqJMgk0EELB1y9emT971wif0qRu0LvJa+zC15bRj0Ub9DBE4rQWDI
MP71vmpOM5shrQl7lUazNf7EEZS0DDYas3q53ewNMj1md4bmvHvqFq7FLwPFv4coMfUevbo4HMaJ
L2ERXZIBZt0QdOeBygnxAtFDr2jFqPbWES3CassHewl0LmJR1cPtLnqa6YKVtViNTiOIsn7hCV2U
WYnHJPn6m1lL7xAtUStFnZTgOFAQ9MsJrMCV0PslybNhlLNHcYxLY4EMzNUd5HPIEq/Zi/NM/X4c
IsG4b6E9Jsyu9m3b97nA9SHPVd981m3Bm48F4fS2PbUpWbwQMDrasbXgMoYmeBTUfslj2OtvlmMs
GtzaPiXaLjw6zR5IWqv4vZ388EKC6c5WnCHjC8iHhNyAKS1NM74C9gkYPTNJ0N2qrAiETEsHD0gF
fApWPVwIyjB9lzmmIr8MmCRd1+MjVUH6L6yOhlLC3AmAK2LITrL9BeVEiKjtagvrefnc/P+Anfh+
MKwxuKC4l7QusxRKcE8v4AL3JgnKwIjiW9nSJPnTywyiCiJv5ipL3Xylw+JujnX/X7TkCPylMBA7
yZJRf6Zcp5txkaw4AdRHkW/0Trxspky6QvuENv1lN1koyzre1rGdSZsC6kEzmidFLDqol7Z+q/3T
5emjrFJQbU/EqC3Pbi8E9m/OJOvUymw9B55gLnmNJW07qVwv78cQI0ojmBtUDntM65FHIJozu7/l
27+q9rGbu1dMsffahkceV523SAy6OeZ6IevGAOP3qElniro8fmIQqpYnSgzCeqIAyIMqM4N0TJoE
nKtLvJwby6y8ep8JkQZyzc1QzWQw3k6ukKI824Q4qHp+T5kbGFRkRVvcMSxXFElGJU8m8Ofa0UAZ
QkpMVd32ld5XwETnQHPnHoweRRX/lmo0adW6fOBlSUBdkkWVHjHXco568QyP7f5yREHxx5sKgL5t
WCkxhWyMdIaj5ggTDa1Bm2pKOAiKj1FDE5/hVB0Fv+VYA7vev3JmLjyBk0KEPN7/UnG8l6G6nTT0
7VETre0UD3+x5gv8856m+EVt1CSTN7kbkOq1l49R4IWrBlPMoDV8YkVV+09pYQ2ce5uYPVDAfDbB
Q9NSLAkyGFuOVNQb1IBB6XtsvhOl8DdJXny8CAUh016fA75hGadVm+r5wEbPh7nCGN3mfkPsy2RR
TeG9GVqp1suhQ0r+a1OMGxcyuGEx1RFVjtLM9OwME6oxHq3kiLD3dMhjwDdZeugJpA85TPoTfa/o
U3QYxHzVNFrfAsliNPU/oXi6JUmEktd/fF/xLRMbNBCvw14I1passoAMt9h0pBWk+S5iYy3m6OM5
kA94G80e8SFas5PhHxKZpue9Xku+ppEIiFxT/muXML3Si4tKp9ynUdnjRnTuC8uMPr99/aVQpXMQ
cnlUeSir8cgd089w+xrluf4EjrJClIWMQ/656qZvufw6J8H+bBLSCMsQXXRdeZALIS6+tA3jcLu/
cM4oXUnHv7/Wan/yyQY1QmeOBCRKaLTNgkb0fBh+wMXSQE18MIgy8ejxV3ZWGIdTa9jUoVK/FG+c
p1Oazq5yumZUa2gJA1a8MGck7EtZ4MQw0Y/zDcM09OjQ7NEIqZY1TSHihW9c9n2Ds4fFLsUu98SB
m1wHAKnYmZ2PSuciXE6YXs1sxutPH6RsX2U4VfD0Q4nFBiBVCbjqmwcg+cg6lNNLO+vzXbNHzvbd
X+IRoieiXrTeg2zzKRjEMeLHWc7QeHuUzzDPhAWWG2axjA1+fgyHp4/UpnQ0tLKLx7IBaiVJg5pN
8Jmglm+gDdJlvQbPsz0I7Lk93BWDTc/biSSca13uMloZT/A1/e/80a5OeRDRDQq4R5GKN4N+8bcY
yPJfzvMNAYBqzLXWrWzuubnflRsepKeyoCY7Qcvw2i937yjBA1c+xnw26Qd5XSFIvFJQQ6/Swybn
jUOkq/TGFtg/zbeHdStiBUHcZnjvqNczOrVi7pju6d2/Bt4NS1mDjTy+7FYGb7IOn8PQCSAi0YKo
cf6BZnxftAuPblz8VgrYZP45XAIN0oNc0A2WLr7Um+A8ZvIWFV7CRUTPtNTZEBBMuA659YPTjYI+
n6RtVXnCt6PuATdITzchYLPYuT5ov9JdugdebQYn+2gzzBbm14ycz1Pz+hL+ZQ2RMzqKeEHccJ0c
vhL8LPDpuMBzUQqlpypKOF88IcDDVtIBCXdv4Fn7I9IQCiX78zNbh0BLlxu7VHHEVFb0DpCRinYD
zo9AjCv3Fxh7TyqnaiwIKqAdWZlKKh0dH3D5r7To6PNX4V+jyWUWmNAs+Hmj3Vsy7NFP+W+S+nJn
JR6QT4f0U8pqFQurAhklwZRoCqOOOlHe9cJqDLVX1rLL8mh9X8wL/m5REsJzH2g2P3yC36d2FQ4D
cWfsS7Ep5OldiMrb2C3giV8s5/4PI1irj330+FRXaiilSj1HL77lnRaz2Jwl2QUsjwVhraCJUMAr
tID4cpJwpTkwhfH8iZ+jfKueuoNuB1kvRRllQVDLUxO1y5YExugbTsljSYOIsXZMTP5LroPm7PxW
IAny8lApR9o+j0wAEwNxKZN7Bgt+RFio32/R0b0eBCWxGDJCVgxXSXNMABsk8qqE6I5hEithBiyx
sVZ/Ev6lBxN66tvzU4l2fDFEsoiTp2UWI56OcPvSRcYbjBSPV8weFIdMhQ/VpByQmjRYpZlVOwkJ
rfIeDB7JGXh8kOqtT/wgRz90o3NOLqBRJ+z9737mCZ0xpDhbk37lQ2RYiuoHFLSQv+hYz/ZCNZZO
Ea5ZXacJKxN9wtAeOOHeU7Q9nQvO5RdHH1Tew98I1WKwSRgza9ZJEqn3524Db7DRfclPBvNuZUmG
r74CXED/vChZw/0vrKjg0sOOWNpscZiNvvqMe1U1i51NgeAEgA6vUSkKjv0xQdHhubUuzmWyE1F8
ZpReB/WEHuqn2QFWa5GQW9RQITgAnmSt53/MDqt+kK93gulBsFMQUsHCrm4nV8zwi1zgL4SMaja0
0snH8RT0lpzLA2y+DqM73uDGhJEXrBcjhlxdENZ0tkWYM5VHxSAo4l5bCUFQSqv/buUn6zH2m5sX
pXLa5UURtVT3biKJBuIIVDjuXJ2Rd8Gnuuo1E8GGnYc8LX8L7vYsCniuFWv1eOCA5MN91Ivr9GPW
uODtdHEFD3cH/7n2RwNosso/YByGcmzeZs/Dd8girHnyhXPNM3ZOr15hxvAmgGBAbTcaSlO7pKLC
4SLzVaxmo4eQAi8gC/T/yr1w6H4nOhrTMSZp24qAjN7WVMmiAge6q/WYshmf0nZ2cUyNvf+x4VPB
lr4kYfLafNQtcxZ5N9xKv3mfexgmYb9rpAm9N4oQP9hJ+XHN0hFWZKnmWf1YEQlEDVBdMEOEvxZG
vNX/vOeKN2jIF6G6y8fjwRS0PItHfceotYUwVwKWgRFDtaOf40elt1K9JOe4a458+ap1Tvzcmet/
j2mRUsSvySvvzf8smy1wHYi5OL5HMFdS2EHuLZanwmPqcEPKnd3BJJS1uLfwo8TNkqR/j68vU/Sc
/FpHSnRJ+6WmRy/ODN+voRv5eE+euQkCd5qUyQyXoiznG6HUh76llIJ1T437ej/3TGwOAdmE7lUd
xhwX18mfP4Zxw41w/2H/NVZfn157FSxGR4zA2n6r9XqOUSvrEMIY84QsCIDs9XMbIcfObfhCeQEu
ykMEOo7JM3iRMvkTDDQ5yhDvEqZKPWbG8okcX0UFCgRzPwWImAMtfAV4vFary4Jw+veMWK81qLE5
fqn/nW6pU4C6LnHuraVhARzrZRkK845FNUW9jSc1ZbGmdhBjzCEduAqcDin0YpchKZ0dgld5NgrD
SUQwHt1j61u6mneo0aTpsrJMU/u7OoU0q5sbrNg5zXfQF6X2H2qvS7MXRNc91JzlMvOQvA5SgBcK
kRl22iOV8YYGhZsaY7TkPD9arPhy5AIe7SnvPw6FLLPPpRCTO3z0gXS/E/PHMi/TcZ+NsFB5exwm
I+HR8xINc7m49R01lLyXWTEt3PWFHDURnSJ6cHdBjH/cMwAjizPzcAmI8cUERP0XkTJLVPqVfsoa
CMfCDH1x+pkWgy7bvs2vNLb64el3XHkBsXa5doUYVpFMqK9fD/2P+pBGIi/nR97dDoY/UvH0JPFd
rnJcdzracVgjEVsJo8/dkhIRyBwSSj+VAoYq4njNJG8WGoMVLd4nd2GF5WFnPvCOyUv5H/g85orO
nkjlFBUZwIIY/j4Bdpak0IQ+JqY8V03OK6M+4nrp8Neh6oK3f4psv04jy4hhodZqZmm+PdDJg9KH
t+vFOGr6nrkR5HMpDf0m0nnakvG8xREozGpLNXNzYTN1Xwlys0FeDowid7CnrH49lweKXLaI5QtH
ahQ7vruGc1c+haqJHO+BHxUP+SDqgCvhaVyJIQ56hJ7buNCyhsXXeo9FZQJkOOmNFQUFcK/4hTQW
wGaFVMM7RtP+i10PKt47DstoD/iSocS4oYj/EIxSEAjBJdWMgw8rRVm81H9MW1ZRkZlLGoJAEKXn
oEWceLDkJgJH6o4efAzpzruEqoRH+X5rzQbJd21EQTUP2AU69Qa489aL/9JNg1HRCDJohINzBoA2
chZNCulbO0Nn3do1UhPzDOjQch2EJh2/YRhEGka/Mnn56n+oFUAlTIo0Uyi6Hxyky1k3GvKbuntR
V6pN3zHjEbWVDJUcmnCKn1E0qJDrI01ngbUCJKcalyGr+6fokXrPetbG4IHFg3bxoVKHAR+32d/f
z7OcuK2CtEBY+nwUeXgkOeroD1oGQj+1MfgqLt7A16Ye96zsQr0p9u+UJokkD0SdQ2ULSEc2XqKS
UbmIxzpbwuHl1CuWsA+JpcCnAkfpvDUGCj6OFDPppLpi5jqfRDSbSCo3jlKENLfnwHq6RL6bZ70D
zgogUK2gh63PiEZhn7JeR4plyQC9IbPd37hPXuqTS3m9PAwLmAsY4+hWHm5LjbSWfJTr5PimVeMA
+J8Y74+GIoXxcZYEFkcJCBPYOZWBBgZ2bKxDm/MKjmEJEo28Cx9+Uas2XtfdptM27quqxzaF17Et
Nv7/RqZDK+woQDjahLopNFqExX9S7VvOPHxCzIVBBMYWme0zf5ByYOcG3kw8QNDPzM7OXdclP2Jx
DCMC3KqcUaHxewQSnJ/qURStt+E+vOefkO3T4E0hXkv3NrNym0SUGTpIn3LBX/Gue7dlTs7VNyST
5NBhm5mUAaVeK7i1iJona2LETyNPRlnYIVCXGM4B2XM0LofOS3r2FWBvgXBev8/yp7x4TCYxcD2t
C4nKWytpPKm3M+6FcGl/wbc42DbsmW+iK6oprXcib8zOyAeufAsx2CcVilJNni8j6/uh1PeYtz8R
hsmid5waF7rQpdlD6XvLZqLO2rhe7gvRF8nDUk4v2huUkmzTLouZWhiRKg22H4ayeNrmIIOqRIP8
bZ5qkL9pwz1sJ8xMv3L9Ie5EUI/U8CzWN+1jFHwXxTwzBIg7AlzVpaU9/LgMy5nx67BzFn6AoVSE
dbL450Rc8nOFxziRxka3+JxuGSuZHtTkkAPYHpb/wiC23NhkV7TRAtNEjKKDxiydpHJ4JAbIJj/w
1Sb0j9TNCzZjFBlnQxZG7LhQ3JKGKSOKImL3BNPdJgsObFqLOYkO4e+On1LIh2fJOYhsnlcqTqyx
+c16Qpnu1B+EAzMsLYPXSJPV2Xmx2nQDXetkhvo2zmSpKGHDkVd7gR4yFEyl2nu53ZCYwm4PRfST
f+hntsk/DELHF2n75c32Oxbimkmdzr4CNrYENeYbavhEvo8ql2lDlnRfbvM2aUDliCb4jwpeTwJ3
T+I415xCkd3qVQLIiqEHmaJnjNFt5D4wXxhoAtzidMRZhBM+O5rFHBgKBhD0ypCjzAp8ou70Xf/+
GKGfJQclooPXOoy8QvbQLTyXPRUv285KjfTjCEaI7r4eHudrhjELUjU0gwipsu5Dh32QGSV+eaTH
9H995y5pKA5hTrXkEpHKJGVNTXyfJp1bJ6apzRz1mwel6mXknuBnA05ZYEMsXsAzigcT6yRkwcEK
vnqKl1YyZTw1falYThQ/8pHegvrjiL8fDxx6ErlozbzY9fiB4DolG5NqagSFyR8Aoe+/xh7woMPq
WvxItFBNoW32voBQ4kM9MEfZW8BFIkeFat3Qq/Mqqbyz46cbestkHrLT8xY9fbTm2SFdQcz3onpe
6bXelnqCtzf7hp3te7gHJU6JqpGQESkV2kAJqoreCzuvCVyeUTiJso4BcH30dQbV7kZDg2KibCZK
6GPWLMQya8De+c7OZlYezakWq2brYbv5rDhjH/LiB+7qQu0KVgYsqAvQM1z0Lmr5p7q8oBAcYNJ/
6EIEmMDtrb++bfvMxVRyqbCkmQhnK/i79jIyYJ4XS2J4yjJcNIYTC06cTMQD/shdf3SOl0iHp9ka
GP25xzN5t8Q4/81o18OjbtFtFZSbaNl0wHidsthUhcge+45cfNm1/vMNOftcIQ0mtLqWhsMFwvl9
pzys0NPDlNG/5EkcXoWJujLq7SW85Tzjje2TqbUqKPYMuNBqM5Aq5y2Ae1S0/n/dnPPiJqR7HT4/
s3Pw3nH+O35qoM2j5//h1Fihy+uk4Q4nXPQyponztp6USvITIbo2B+1SCgfNo/Fpdop0bKTGw3RW
lYk6hh6DKhNHZxs8U7hZVJA9OmirYqaX/riLgWTGz5EWQxeSgUAcqRHDl8niOEeSbM8wD9BIen4V
MGYiKM9+B2sXMSuHzOfZQuNg04gogRPZ5naz3dcaZM+2u2nELmMS3d/oDxEkmh2ao7zBbCWbFmn4
9IXvlz38hBRLffUb/8NHSOeU0NYPwI6drAZeM0E1cBEcbnVxYZQzdY4SusmkZ/zsmOg/7Z8pXojJ
ejWAQE0l7xXNHKqfcHcPoN9xaRvg1WkhMu7KHzsd1HRkXf5VwggOl9PT+4x3EUAVqGC9mK9CYjKU
zZyJKKQo+rl1DgoqQ6J76+gDl4U3N9Lr2zfQNUFw7Qg4PS9W0G6TeetCJBepf5GxUEHE7F16kKTz
ht2LeInSxdrbVMydRPCXcxsdV3GeCoVrdy308vyvWRArfDRLgxaAjUbRr/+HkBkk4Y4pXRe0QQJH
kI7qRlfk1Fg1kyxhGE2Fis0LjJdCoEudPcQusaqD36osP5seWwihddvBIlnn/Hw6+3QFcn77YVII
Fe+1KJgIBELsGl0deXJ/JOUBpIy2RhX+chhrZ7RMnB16eGJ6V3gqsmp792wnaGBKx/uDZ6SgKsoE
++CI9qlmzV7RBQ97psKqyX44Fi5X9WOyfU6FCBvLBFawwbe5h+LovVRDbXkztk9xzA4bXCMVx5aa
CYF1GIGTC6iC/jt6L7j3TQweJulpUXKT1/v2csM9wGS6rcqH/gU4nUScJ+LvowgghawNbSwWy2s1
juNuHR+J26vTiIbHhN6z5ykEJRl74lMKqHfebC67HHW7tWDsDZgK4OlW2wkdzWIb8KL5ww+I68aW
QjC9x7z9phY7C+fRqXZsRmzhpBm5BcuqF+YiCK9Fytnt2474kbky5HJVGjATzK7j6Zf5lKbIoW+N
MEjGNoaWWlITMtI6RpH1scRRjxoZ1JBd0vz0uMedm44/0toHy6+md54+xJJfLsZXtljk1o12HR98
sUJYDF5B11oWiSHTDg7CGGJh2Ti8502JQAmSoOcTtRFkRM85XOOeaKBX8/KAL0SedePlRHo5wSK/
0CQ7N7JJwPHv2GmbVwidEuAUs6/lg7NUvb9WcMr6uoTA7PIqRv72gNYUj91AMgnGe9sgpkV7H9Bw
JDF+imBqERdyXazW+kgTQy5670RJDE8fcbcDZAhMovp+U767kRjjKVibiUgzW9viPvjwzhmVzHdx
EZZUxc1OrXD8Cn6Yx4s9Mdn3k9f8ura+p7rlfoA5SoNhtRz8Dhetzw/p/QuK5dLfJnChoSGCraIM
BvJaGDsioExvPXITilXElDe/bIJyOMZdRvUP3zK9NaL2MiWRfZN4vrJ8zfH3doqp5i3JKBy+idWP
/n/rT1UuqD+gD9G74MslfKCgq3CVe9x3APHIKElSJ3xf3YpQ7O8NkMeKmhtvXUa7jvKR/i3aq+AW
eYeDTKCtJDreAAjWVCWvG1MvnR0AfbcHVoNIS6mm/APuuTZX/b4KxuXDcT/qr3gWfevlvr8466nY
2oPCec6uiNfuQ4n+5sv10k7pMrtATlz2W+nAHvT2vEieapjE2S1d7ndKOxt2eQlQu32ljMkSPE8d
Rvk8wvo42ayd9vBJs4sGHh2Vd3ccrx0a8LmUVWhKsBuq7hdI8mZNJPru2+VAN2pNOfhzEsbsbCBM
wFlmVT3ZFRWnvKGSNuH9jC3CsFcW7FMzoYZaYiwXQBLwC1KtU3lBKgh4WY9+BP0cAfX5xURLBtZa
ht45djd9LEe8iZS4U7Mgg2W5RaxkvDmegIGTokJBaynehJqZh5TzdRb0r4wZYfjX/BqZ3kn+wWql
49Ic2DPpy590kzBhkOHRFFRFBBEbWvOoeoWYA8UVNoZM47lCkzKfMPhS9gBzNME+PtNSAPaIME3D
MebgbKnkN+SuJdT+ejVhGhGzeZCoF4PyDq5ZvxYo1rPidN+i3h78nP96aZG05utRljuWFoSpXLGf
WUpGtO8DqM22lj/LU7npQ40X16bS+6ElvhmG/EfhMUj7pbQGVWB54bv4SoHoaF1jbozsOL79NUc9
gZOlf6dF3wO5akM0mjFJ3qcprLpqaSqL2GRgBdNt1laNkUXNe415J5SlZ01ahWynqvo8BzTpcXS7
GL8wsONCVB0REGu2lY8hJsYEqftXg5t0rdijFR/iyNpD+eVibuENVUhhvFo/zhzSc5irnzG7sfSH
DrVQadeTY3OG26geedttzfto+tJ8Xm2mRRcRZT4o1JZKhOqBDsBhCGSK4WT4VXFOKEOCMsLShP+1
ocGRl8Ph1jmP2b5lKzVMQncnCl1VLqiIGwR9LhYwwidVTAbyMvtI89BCHhplXKEZ4OJEZK6aJlFF
lHEg62b1UgnaVTItnhpjTikL7HvcSr0XK3QKHV14Q8iy8rVppW0fptfJKotego69rB5mHLaETSbS
0LnPsganW6uMrz9AEl9ywiUo6VxFZKVQOQePPbpiOlaSGZ2Rg03koqWAEMUWxDXZ2DDOPrbAlBIZ
RlWhdBkc+JQsfTMQfLxlqssOs9LUtfzWo78NkD+ueH5UBGb+BEEmf3JceUFpuKSJuf9+UILtZT6G
MxM7wDL0xhB3TgmrL4pivgrvHi1zmodYIi0LkMCuSAAQbH+3SFyPpNBo87CdPm+15coWddU21bZc
tFz2zI5AaV2MpqD1OtOHf6VJ0piWTrnk2TLd0JHEh/GNEwlsKQtV+NVlL+0Mhd2LOOx5+yk1BVei
C14Sp9z0oTCNK8Ke9vZ4IJ+Zk4IU9u71j+pDjIuGdP2kOLUJVVhwc4BK/ru3aXf9pb0csLRZfbD1
Ep2MccQl6s12W8j0afgFTWaeaBGyv2oHkn3MDVsMwQLG8eQSa1PeT6cLbQbQzxccaQIQlUw6Ahti
XwhhpqdEUgO7yLGlEbT13OLpMscgrZSXakEqt9bTuMbs71m3r/z+fuqysCGklTtm9X1xMsIuYchZ
DZf+n+hEg1sZ8+9/dmyUuOpqSnoHl5q1yk3yCUh6GVkHzgmrdEsu3eno9dm6DCxQN3nJfoDzN15a
CwS0CJTN/AyXD+i2s7r/VJg/yzXh9rcwc0kP5uezFgH3Oi5qMENvIB8t4GK03WAt/C7wkqPRkDk8
Lac5GXL1oMG89U5XWBHGwBEp/R95QWEQEm+/riphjIkg7epBcHKJmJ8heG1TEnZpqlQuWHQiIyUQ
HWKeCdaRejfszprxrJ1IDvFQOnVEd/ADxMO+l3DgG65bES6/HP9IajrX21Q9Dt6tVrzdDt2aXyaz
wpXXfhFjtJouQqwiMeDN3VfspWivhh9shd0IWnTe/9IUqPrNyogeWXI/DeQ/lRNiuutnaxvYmRhr
UwpXoHdbxVYPNvLvtA/ltLe46dbY6RAGbZyriGiMA5SkiD1SCKcA/IyVIqFLQaRXu+HzhaORJjKP
I3rmlAy3nBqvifzni2LJTwURfUTG0mDee7XqFORcWGi/vi1rNbzTucnSBI2CQPBrz12F7Yxz+Q48
Apc6vee61cfyHKLWLiF5PbB8QE9gLalstCEsWjIdFL1qCPsP7tFe/QwCn3QwkuSmz+DD2w619C6Z
91GtDIgpopR/6gt+VB8SYFesLQSLN+Bozczf92ByyjD71AewbjlESTy+Hfl6VxGz3cH8N4W4FsS+
jPj5SrjQYmmsjrD8k9aPJNpVpMA1aT975W0gYzg0At9/f03mXyZzjuSQRLp7J/ENvhdxcLep52Ww
HQ9hrxgPctkHYelOpJfrXknnRiDMAEeaGk16pjq2CaAAxk1B0q+QM7Bb2JN2xGUmIXweV4duybxO
8Slatj3keXtgKdJS1g+r1n7jhnNG7oiwCQ1nB743Cc3/11H3HmhJV/LU3n1uUo8xJidJj7WHot+c
LSnvEgjNl1e7Na8yidAE5Idx3W2g7lQY7woEJ2vL5mhV5RpvgjNYehojEWy88P1f5KMHMSUKElg6
FDQQoBT2VqPhhrN4pGhd48C/5ffcHlf6u8I7quq0SxzS4N4z92LXaSS2JqqH9p4fJtycf0YqZxPy
7TjAvxbq8L7Lf8muI5UjHqKIwxQylCM+kB7f1YjPIsY4chNvP/UkkrYcYXnQi6X362ZwPz83AvC7
H/BVnRLmUItKX6Cgjd5oL9RxrrJfYP0m/mLS9bmXG6c6WPXX7bex6Da2vchr4uTm3c5xSh8E8fLp
c7BCelBb7EoWX4k4309STA9/CqKozGunBbs455BSh8FyjLrj1V2Tx9z+pPfiYqU191bgiztegZYp
Z2TT0oX3PYu70j5h9mGEkrtnfIPJcR4jnCzOGk+mPuaSOev0umZ3IUS75y9dj8hFKatdEkjB/Oil
6yOCO395/+q3STWY3ufYvLa6BN75lBqQdv1QF9+nbNIhDwrYHH8tqjGpKPyeEHZcSTOGZHxPwjVQ
EmItq1IP8ARxYLJTLiFfaW4F/V3syLHfAo7tyKMwkjX4ihMWpiOIWMd+YjdVFx7GOcAUfB66hfwL
VGfnrMAL299GcAE+j1Eudtj94ReTXl5QZYvghwHdRljw4OtzltJ/s04vJNnBxDvFvV/E1hX9Dn39
hgF3FTCoT9aHZlyfp+gCEf9B23uzoCLEq13QAGAJaPtDOPn7Us2rI7BoeuQnOB0FEShyhbMiPJHo
mr1DZ/zFBzdGZ4LXBIIapd2IvWXOiphhirZH1i28xFPy0ka6V0kr17m+OFKFKMuRLjdT6CIlcF5a
Sox8RkYXtHso2Qt50i4+Ivcg8NmS1ImtOpFURskDoiCQluonmVU2bBcPBrWOWPc9c1jnL0jMqfoo
FJSeYlgorwMGgK4ZVR/Dyuf4WXxo9ma7DIdtgNRP6r/QGKg9ucaCEeAWyRRcJgg9MXinqq1igXtq
XBQfFKyE9ADJSg6tUCDt2/uEZNI9l7JescL/RDR8sHwRP7Breol2pLzPu3kYghUftN+9JYYMsqUA
rIlt+50/ZsVHLgyvTE0+keEnIP6C+7qtNjsymK2mR2qBEwTEvyYz6swbKevC23RlND2jNzMlPZOJ
8cSU/8Tpm3FHn7tBuOsN/XktTG6DKXmQHhoKdTqcpi6O3LmBDNPH0laXWcu8j0EeCC70uykaI+lr
uT0tlsPpbpKXwXMxUlSl0vuaCAvcp+oqu9EXFW9xJNuUvRWKMib2HMzfgfZI4I9s5TEGl7sp+DIR
pSCDdogaSKWz4jcZtl/JP4MxpY1ZvxW59CSTOfLd7LAm0oNejYh0jw2IXVs5QTF8whCzoNWm0INJ
VGGL9Ps+nMTiXmYiyVU/maf6rEpocsNhfwT2tHDBLYAtn0xI7dkp0711w9KDvq2maMKk16K8eqAd
qIW2wStPc0fnlX+hM8Qyr+nJ6vTyMIIHLIgRZne+xwJd2XzjHzs/0vlB+hjHVfas59S5t6/gWq1+
/4xiVG20E3RwJ+bqOIu/WAePNiEnx9CGpIhyXAaA+mxn9fDTLTcDUllwy8sXSBNSoClzXKF0/DkL
P4E5DlsnlN0mSJUYMRMvCROkzVQIzHl15Dm7p7KJxNIXM6jTt+SQvfzpSUEqKDGWu7JAAvyyR5mC
4alSWa04Svq74hFe0KrWNEEhuV96TJq/KRXIgDIJDwu6gSSEPWBymS4/k3fj/OA1mewcPxW5jgV9
gNUNnmwHVmT6FqzYrlhkiV81pKfch9ywHJRAXJrlp4V4XXr5HiLikZ5iDzhygx2isj0DDh1X30ea
uIWZ/Xb6DEKY4suKe/8rVi3dyMeoTVfJDggmR5LAjOSShEtFVYF4ZtaOzgqmM3lC82J1FvrA4ONd
bQx+8C3sRKhqa0+ibjIu1L8iFEfOmdAmbs8KT/qAQH4NzAixxwk2TruQT8atH7n1l1/2NlNuAfpb
aSYOAgIIdDeZYIf2TwPn0iNwmt4p+vc0hS/7l8GZRef5Y8azawhDYiv44QO3YBx8yaalZZPXT3oY
0Zar7g2QND/4kLBSl3j/Q3AxpiQBLDyCZl45U8SB8CqYcfuy36NLVbBovKs74NAo0zCoxnP5LLXS
V4BfexmwEYZQ50CrS9dnVVelnJxT1NMYAissihLsdtXAQAbUsvBmVc0OWkSMipfcaYd2nldEuWMg
Gs9CGFKTG9lzdCLJs4eISu7Hgl/D/Y4hTnfk1MdWBIErhsEaKzjh4JkOCgapZXRUXe3SzYWNJUSa
7AUnN6rorMEkj2VMdMbiAkBBMSD9+Mh97UU15JZ97aIJMT74VW1NMyW/LMN/Gi63GbBaYC0Mm1h8
Zv3YbPP2dIVlCzj60oCmB5h69rW0sHSlKgbf/Lsj1ZV9oGR2EGVCHSAMe0v8pZ+S+AqI+4mCJG3F
MSUNPqTxasZoE+Om6l1js9Q/YRfkI/a3G69HAdGwvOnQEXBGyTH9TxccGT1m7hse0bARzopW3ll1
naGgY1lMcfxsULmWWBafH+dpBlArOTnp5FJwQ8MNyB1sJjAx2Xw4+k1TLqsWR45nSC2YVkFTBjJQ
PkL1YD+2+QrAyeKdJkko2PQzwLI3mS4gOpWyFuqE7b7GENkwRafnClxlr5Tv0zchnnHsZnmAtO9z
OfBZKT9gWPrSCLCTxcn41JiqnQ+/jJmJ/qjznilWCipiKx/LOvEnRQgpfZk23twCz4VGhKLORQTB
5tiCWldfZVJvNXq8V8T0ONRu6gIyW7YcLiJEq84qQWRq3XgdseRfu1JZeoxGa9y2uBNv7VjcEeS3
Z0CulrQPJq9I5zA/zxmJALQvKCWVA2PhL185fR95G1DtP3fHSlw9dnPYce9E5nB5+oDmPLMM9eof
5mYzca+4I0bC0TTGTFXSi6CGeyjQLPNAc9aeRsU0L+o3dh7BO2tqiTj/QJafqVI1/eRLEEHmuwEZ
WnqjWgFKnsWflWUNrSU2bCGExFF3UwVir0uunGMnubGv5Jwm1rrQLdPeEAwl+Hb8G3aWua6qbWGO
mzym1QaREfdmrE78GIDcMhKwYRpyGMn9vH9FMcI+uACW+5hh8BaHiJWa0mW1Ul/KsT9I54MjbKeH
HLGoKwTLkHKK0lF7Xo+OX9z58L3waTlAFmf9KrxGw6LJI0nlHkwx2uKFlCGPMjJLWD886ZWd9+0M
z6GxOsLa3DUHyaZRkjDRdoYBkLkSb+ISrhBA8jsNRgSu+TEN019wjDPEfz15+8YxKg6na3qgBLEa
v0OcGhnFj5djv7hG4m7fddNAoG50AesG2Z7xvgmkb3Wl9joCBRPkA5AymWu6X1s2kMVLngXrMGJ+
HOqzlDHPI8cG3tEJrcUMs3bLYSy/QGn6lUpwFCHmCcHfDnSAw54scZ+Vjof3OqnKZFw7BIM6UYmZ
UiPjLuK3D5nBWDzzIWWxsPosVjKiI+0Vat6m2+pR/hNP2+BqSWrwa2b0yZJIeY1xkTSUaZyZVSxA
5c/8Bj21ftaNd8ccEKcaTatEsugYb+qymYx/oJQu5IbVcwbkX6iVpm2Yv4fPQ64Ht6y8numrOkXh
/mYBSpEDcYYFsMPnri+i47+oVnf1CXKnQ08HBypKCBvQouYIDnI6sVLBvmetJE4aEEK/yB9WnveP
2E8rCNHXugpqhHuQTAeCXO7b1HuZfDUZv5cXplu/nbBRaH1uXFyJJ3MOBKSjrah5fV4JUxn21CvW
7LobjFheyipVXdcDMVZsYBhvKHPFXT44lQCk4Je5HXmbLW3leQFJrUQFPNonOvj20Imi0yOBf8x/
aUxOUjiF0sqln2vL7ATib560RuKh85PB0HKsFQdR+HOTuQfiB8K9fhkthULcj2IDZvzJ9IjqLlBN
xNQLZc0c5VMoqmdQCMXxWLhziGRieeRq6WhWM+2qGZ2wo5h0fnQFfS8c+dfyFqSsD5x4H4jWgU8Z
1o0h7fY01WM3VlOtTuGGaL7G/5UpVQEmoQZMAOiwZ9Y8nmif2z9i8rXfIrrRXhDEwxdTmm84NU24
BXD/5ASrOxTHXSfr/gcGzjogdWqPeWg+zvTJwDkLDsgMDkuqoPeRyW55dhftTwSk/kNq/kAQBvBe
EfIQ3HcI95jn5xvODiQeAilysbwW0Q8D80qpnKndWm9eVm+W4+l+DQn4GUOkhdyTYPrT5d9+TkKC
rWRzPZeooidHppkZ/DcWmV2YAgDpfzPza8YdtDbCCvE0RwOgBj0XRnDJwAqc0/dS8Qn4xaqzcco9
8zOtizvjnjdCIjPREE9dzckw/UyQzjP2zZgJkHDLgh5obOa0RUfwJd6Kdvfr+RFauCBiBj6ubq9u
FHGaH+hgCyVLXoXOQQVs2s/jO3VwoE8ROmJyZgX1onPtI8kB9tMrxdyuc8nAvRRL895AI0N3Vccj
UUuSNWiUY5gndAlWbgOiTvmZBWHBxHTe2oujZKlvEmVw1kqcgiiokqtQ9hG5Wv82C6oGqCLTLlMt
tPOz3lvwJwgyANdRh7MYePYq9aeSDEwrLu0in2b4qth4D5nZmLFmqeT7uaO+A/68SVHqUMpMXESa
FoGPKbXueqBe3qVi44rT8BdJqM+4Igr8vmf1RdM8AT8ub4TyEXYBhJD+FAqC4Nb4GiOvuVCn1H7S
3K+Ct/4C3xBfvVz3zOokjQiwf7Gnrb7BPJ1ZBFJEhKpSwJsdwKRFeQnByU/ntxDOeS/OHHdauwlm
5d9lu2qTEQpI38GBMyJmzWQwxsScg/rU7lP+2jL1hrpXCbraOJUWsEZM14ize1y2awa4GieyKlFg
+dCqQLFHaHjJnk3TvA21EW8k5gJ5l9T+3cJ5yr3LZnXmn66iAI5h+8m6EXPx58TJzRViR7ggLZIV
qrtVNjQgRK1mNhsLI6g9HgKiRJnsMaX8wPImHLG9ZYPJlKrnYjIpY5c8gKyjYTFHThAfKE3EsGTE
jLQRQnUYa//XLnTbzGhltz4HQQu4RNtO9QTARLnM+AX+BQndx+J5UaGajREdJuanZtdFhNsGwUyc
cDy1QpXQkCHr/SmjHzgxD52iMZsDSaFgyqJgkztwC/vhRsyf/W1LbOShvu82JSgsVECULwYd8/iI
iQn+sgpYQ8iH+lYbVX9vPBHFhtPK8ur/Tl91/Ua5SVNFjcYqL5WiXo0Vmnm86N8BHdO+Tp+YHmo6
NkECqTMuyrWi8VRcotBB1g5qkVqbjefPuVez58XlNiV2lyFyY5iIn7UFt46wlEI7IWGU0MRhnUA7
miwiMnwcT4mjYRk1GoWq43yJGT+OW1mhkoV2URqvS3dVYCd65s77OT+zSV0OvkpTEathnIP9PWHX
tJ5C0HcPvbHo9LnoKmZfCJiw5J7CSSLc/pCo96Ga4p2nRlAx/8Fhn6ovQ/XX1NEyz1OOncKhGxZ6
YkXP4nA2A3wl6MxmkwWxYMBcW4+nlOaZuoOPKOkTiz7zQHWoTI6pEniJQ58N60QN7HTOUxE3+6oZ
Zgjrnpslwk/VEEJz7QJ4mI1cJNOyAqIF3iffWOUjUkmIzP53nlwHO0QmYeOqn7dZp+kCEJI1ghfK
yYolTgwFR3/qc7f7ZicmFwH0LwyIhXHK5l4RD8P54wgmzJplWI5QaG048otnuauA+8tuab1Ws5v9
BD9K/tqEuZWmk8o2ZsnnAmAZfbPwQTEF4njK2RJxA4Qzvat6z9b0yMySiWMw5vyyYIv3i/cGR95w
TpAmniMGchCr2MK+movN62hiQKpIXB0zzMDsFL2PJJZVAzg244a4+DZ1rIwfkSJpOTfszbOSyT0Y
FHGdTWzLj0EBrZbu2MxfyR4Bpi44HAZAq1A2E5RL/mO+COoL8r5nxvbmN3GB4/mXBOLWskmbyhxb
QdEQzH1S1LBvk67MPkc1sWO8HA2uMzllZCeT9816e0H/dN1M7P64JRAaJxRlaD/r29AifkyOWcK+
DjSLr/cZcSWowztWYgw8s0LbIADnLBh2J70n0rRie8CLB3OtHt048kT23ZbBPr/dLQ38v5wMVMtv
Kfo2EhMPG4dhRr6dACHY4AsJo3D9XEhJDgorsBf8EAoZrKNzCgysGFbGQQazzKA7OEoHjbZ4rzJT
Ifkzt9pCOaDEm7I1fZj9rQsfcUgYzhVpK/6dB+rgzP3qgp2izMZSfdR2jotpecDIbXGU14T26krm
Ut4kjNW4QoeexH2dzMMr1JqbIcf7WL0y1NCzsJDBDSDhdbGvjaGfCdxjBPnRXIhXlm2w0A71He2j
mJr19LWiPLCZOrjHi71QWoc/tAuq3veJxq/82WNd7zPsGS/IXtzLpzPE17enPikj0iy2WxR7O8C9
JfI5NIUQW0NoDe06qCzClDeKoNoissEkLDefvB0LRFyvxYjIxLKIlou8ZIMfudnHy/FdP6kekmtR
5IlPL8hJO0CpsrmqieoRGfejojkp7fKRku2462pyxil2En3ruNdunfcpyJMHBV/Vc3JeM7A9ewVc
o6Rlh0qxXMzKbFL9Vf+iP5dANYel9jdMJziJLZznRg6D4/1FWGk+hDOIDRH6ykZ7P7XXLlJ2omMY
GxnbH63SeL7ITc7u/B2Pddm72pzxxZ8YggJ9Qc6RM7lq3vvFygk+9097rL+xvoYUslycEbJuaOdL
n6C/ZEa87vNYZ21z+26wcxTXWsOCXHmAi3Egwfy7wbD5sVYs551U/7UXtcP/YHBgBjLXw3BDv6QO
kgaEHMQQj1qPNhYWp+MAQocxldTiU45Dgssgu+BLbe8CFGkRw715WHXDiFymh9ubI3shLKNj0qnW
eqwp011Kf9Jjg+bg0zUzbjq98W667qZwEsAArStaMvk+FzIko192NhvNx2XxkSX93zuvVCB08hDI
Kewv7iAlZI8X4pu1kUOU8ioUR++Kboe245THKeHu6e/5BOuBXCYZkK7TJd6pGWsvCQu32O9lrSIa
0Fbf2qTAb1atHCnZiwqePAjkvsGjlBAI5iJbWmx7Ev0URL5UUi1/KKn3nLpkSVtrcYNUIUzs5Aal
xNwfEAPbxg8wZxduMyOHsUXRDiWWSqFmZnc7YIW81SefxMspDhameb2JtD8QXYQw/1seXj51SVMq
Vvu1uEV5cElG9x3KGQKc87aThXeZfNehVu/h/SRpyEFhPo66z39rE1+x1TC/a8uEtMtaVMrGrbFk
KJqX/Bcs7UWP2nL4NhQkQ6CkPUEv1kyMFWRn2hQX8LHCh6itoH0tEnPo5+eiQMGZrONMXOmFLGAK
I26I0OORibYV7DSgGypgjal7QDJHHXR5IpMOg43txsv7gyg05I7+gOX1i4oL1KfoXQ1ISKNlOT5u
jqFTKt9bMapXFvgt3E4OtrXSJbRHBmGWds0aT7z9y1OutM1er0gPfz+aLNN+0oMP4/LNzvI/Hds0
A7mU8y2iVZlWdd1FmfReZA3J7i9Jm7nY+BrGPHOZBX81LExEVSJotYcvFpKa39uYIqDOn/ARkWDn
bddgtbkg8U3k6pa///hIQmZTLHxxtYIUHuYANqgTLRINB0T4VJH+gpkLX2tE2sqdgBesjrGfbhSc
2HAh+nUA4OpWTKAjcgOo5tp4tA05+2yj/Mv+Rce5xr/E2MzOrqtEF5DF6IdSIwyH/nze/arTd39X
ng9FvRwgOHkmoNrjinYOMwG4jMoCPQTo/xod4p5vr8uFm5HwydbLoek+UDLRHeQxK5B+CDqlEPFU
UOgUh1MuaJKANYiKQ17l/4hhOWiEuElfJanNTZDqsaQx3a+2LLvawhiHNowPgVTOHroF7tR021CJ
cVVFL21AzK8IgVrKutD4qgEfdp+WS5ZwZt/VFg4rj4sLhLiO1+58FtsvkIp4sSGpUujw/a9gNcQc
3wIbrlfEHEtQuDvk0sHk9F8/3UmPCrlYKdy1rIE92GbawcykvYS2EMTE/7XEYCOo81Q386HF5ffs
94Y+5nhNN5oBegRBrRpaWua5r8cN0c+bm5oHS05/bLE0k5z/CzUwpv2dcOpRQZWlb4a0ZWb9KAZX
Ouzkz4uoyRd0djv5Lv4OLEVa1ZTwhvQR2X7d3QS141+F5VqtUg1tpecr2f7geO0J4WPCd7WNIqcA
9Mbk3mq4M66rK027gG7sTkOdqnPVGtXeRWlG5Kwjfir4SK0wRzOqDKwpECdxTEiGxPwzGoMwon/e
PUhes+coOkPDYr/epX1ol5TC+RYNfV833bvjZYpCzs+jA9WX/iScmpPMDskoc0Bdtl5CDExHdZmI
C3dpqgukzqf7xTfn6z/aYKjzq7kS+849O39RsqP2NKy//NZY3WC35t0n3aJ1QSlumpoHHeOMDN2Y
n0W4SmWecgKwgPprSKukzK1v0mMi78sRoH1QCpV33AYXrPpjTd3M78uvTTqg4X45MZqmiCdRzMOG
fZpULRG4XC8OHOqGNfomSVPq8CUaFbbLVR0lYk8f8vIenBUKipy47BMFHTT+YexYv+kZG8DHyxWw
hF2QhntL4By9oJuGPvTIYajtCT4FezD/gPGFpK8AN70D5WzA8VpBZg8bGUU2PV6n0RvMQ7Ki5u7t
+i3tb3e082T6qlU+ZZFJe/y0Q7HGb6dnDjaz+yTrf/oJXEvay+hmBsOCdalkNlz+Skn3jXOaOdOs
eC7v8CKfSbNsDA4hzvKYzd+3YEM4mE7q8tM/Y62ajNehvWUn3l8xT67O4wqz5FyVEiOTkSvH5C3+
iT9eW39IuiH9mEmIOMa9h5wN4rFGwFXBy3P0DkjsYgUGar3NRGat/8wT4crA5uuAjU3XpGlOTkIZ
rjCaXPXHZJMmWS/4X5kwiPL1cYuxX524j5+q1rqUr30vHfm9Nk3KA+Gc3ZsHiSWhXdW+qzuT2PaT
eTJ2UXJoH3RYkRaNhxIlLI6Hrmgz3WU6VIWGs0GecbZ7yPRWuZ2kPgE36tthiUbPHI2sg68l5hqj
WqyRzALrDKgOYlObqQxAAXxHgFP6rwvu5poBTkACnC3+NYajV3XjzbCnRIU8kg5aY2X8VEwxHxlY
AgzjLHNi5B2BYqWBznWFbv1ZItkkr1dCLbz2EWf0mI2hEh5KwPYe+vDCW/D8/C6xbJvXp3g2jPfG
k0rzBUn3so72nGsTPcA7ZruuYGQEFkfZ0BBbZAuEXZRFnliSOQ6yN0qxhGP5e1oSXFVGsYifwze9
MOcwGkvmjhT7Ola5TUz7vSh4NXt+waP3zn9q41dBzlMygpxrgAE5rfgqoOXdEmgtSSLhw6ljLniQ
3UM1UgfNIRGPeFJ1pxfJR7HH0Od9Rl/sFkXvuz3ylLtEr+UevTUzNLuqms4eVuHIk6yyOUnkJtEW
nGrBZCgb7rteLV0031XLRDHRfK13h3BJOPYaLcAGUt+Hs0k67vQbu59IbTGySTAtDOvOGkDK7neQ
35j45/FrMVYVCtHx3OHR+2LsKicU/lac/euteV8+7O6lmE3AKRNOp6d7DCIychKOvVRSsLpTHhBg
MhJij7R4n4FLFvre6JTNPEPxyQxXW7zzLOwOzQIaIpSJPiYvNDkSVAH2/ee6PDiMNN/3HXahPR3b
uB9V1KOpUm293Sxc7S86qb4rCdEWxVugaJBYApZ8/3npXNX0oKo0aDkpxDwRahaZa1EDCyTPW4DI
UwrC+nAs4gS/TYbcKkLHLwuNgS3ruStddmwFqtOrWbt1/P21WkuudwpqASttAgQoMGtOSTPeKqZs
hiUWFti9+cGiZSUiLdn+iaD6R02kELl46/VPL+QJCxfSO9FdVqF5U8B2xCyau8Ubyy9px3tqjzPV
GtofcTU3YTUtL68S8zYKh71LaOO94geWDDdZ+FmGZ9rX1399vaTtnX9wvRTEcmCJob6Iu/ntYXH8
VJvsOLMJq/lQPeNBN5M5faXfxUJhrbsNTtUOdbpAIPrSiKntQQrd4g0JSZGOhDAIuwBEF9oJ9moq
rOonFNDpozA5TlJboP4cZE+hLcz3i5bdYTTdZ2DjlhXnv99W99D9+zg8RKWhZ61bIzyULQk/k//S
flouPK/Vu4b5e4dOU8OijrFbfgDIgbhLB3SZfMaZZtVscBGA6dI0P5eFO/Ft7oPPtlcX4OVbCs1m
+7mX8ixJg8+hYeFvokwBH1LNfvPPDNMxD/Haqjb8s4IKGAopB6noPFnFNYg5zaG76+7xISc0ZURD
wrxdyjNT0OqnVopYoFju4dTH+k0g1DyA4AV9l4MTxGrDEET5my3TTdnimUBmwQEhhwYVC3mAS/6/
H9j4LCuSvPFhA31oieW9gqOHYVSz9tHXOp1MYJh9tQ+9jTFx5xS1imDt5SanVG5LLBTn3Cxq+8EF
3yP9biS6LQLtmnmfGSDyB/HMFu0mQ17xj4Pb2RUulO1zaub52Srry+0jonWZZv0oSimDNmbwhNEG
cDSHhPe5j88tyg34ebNNIpNkNhcpWSlzmKMPRI279ggipy3jU7q0bsNzn+ZtkxnAczy3t8JV5p8t
tP8lSme8V44LC9ik+CjxMjyqos5giNWRA1jneLhZ4DmFPkXx4yDqmuQ8bA5BZxOwzdjS+S/v7ZUU
zW8pMqoIZEnyURxnI4eP/HXfWyNkdoYRCmj2dMQwNWU3Spf720kz3mOUzN1d6cqDYuxSK6ShH7bn
nlejw58QmENnO4/ijtXxqVO7sWbhURdt9+XgRFhS4EVKoWNeG9jK+ih0RtOzIjdDmnnLwZ9zYVQE
ouQdUNNAM+0tvIs5eUqQtJXXpKQMGgXiS7aOEwlaMDqObWLoMM1r5Am5mYYMAOLbi4/WeIApKuKk
luSoN9wwLAmI+r0/XWnSiAfD+iyZb2QHAZ7RkrY0m0RjHWcyy26ZBSKiGHt6qWSb+rPBZUJL5qSL
iUHVTwxXMwnYg7nBEe0P49gqVtjLzNZ26ISUIpn2MhTCmRWBIeg37QJTzy4Kq9LEWc+ahttp/T3K
d18lbh9o3YxpMrWbj6mRb7UIPlw6xLFs6ox6wjDEIfzH6u3VdBbRVUptqULW+ahgd5TGFTSuSdH9
/MS6FX9LRnOnm9Ca3hTsdsd+R9KosW9Zp8O2Xlkh07fyyKkGrgvq28DLgKtP45dUAArbBr410nC5
zIaLDAlrsbC8fJPmVocBReua2zzpTZ3fzOF0frOYCWB5m1hJLW97BwmGtcGkr1eQpz6n0Dkla4Rq
NK8WPti9GSbn+34W0dMC6B/G6MCJqrcw1PsZ4t5qrDQHyE6+mLx38x/8LTsW+C3cMDQ1GBLfXHzW
qKaEEAtYwtmi/g026NShYPKRuTZuraOUXHLHzFacS8HCMN2QzCOeDi1qgY5LyK9VaNHa3nXt6bjF
yBfm3ViuyyQR1Y3R3nG0gh1+C/ogaqxLKagm0/BwFMJ3UjTTCJow4yOFADlmP7OBZkXsTOwoYVkN
iiCCt5ySFBch5hQQ1FRJ4x+WFQBiI8FZGkw/ADgq55sbFk1W4VZiKMCsXTuoicjdkAjAevb4+EuK
aPxR24t1R+HxaClIxaijdFHPV7e70YuaH0XKyiab/pxCrDmMH+Rix/eRJz7gQYzeq1AZYv3+UgD6
an8LR700cMQI3qKn2Lo5HWLxACr0bi+8josP9VOLLknQFcDAGWOpAR/wYi4kI9E4baHO9G+CeCgy
11yJiI8MDIgbpilpZDN8AG5hqHuHstH4CmU33KxkDToz9riyNPuXJFQ0i7fKTNHP5fQ2cq6O6gBV
Xw5UYFkoB9VnOMxQYokhl6CGV6+/JeeFxvTFbDmDqkH94B0mJCNdb37RPKKh/YP3RMahK9VJzXf9
WikB/V4A+Pc3pQsq7TCKMVktehypoWwRoAsuXwL6DDOZWCuia2IZ0AdDFfHf565jNhTjpgAQrCOc
ed/yHfFKkYLA5z7YoA+y8HVVgwrPSDTvS6srLrnY++kVTEUJYsnEHSeWZNyFLXTWse1hTF8dR+ul
DquSOfHkMgZhksSgGu1qO9SHuiJNwAIcsHb08AYqE+UWolbmxRZ2wyxaBsNuZEcfcVEMXReLjMqI
R3PDer9UXeMlOrTXuzJbCkh5AG1otiF1KoFFcvry/z2CIiqJkG/wBSj3cTRJRUyrm/HP/YzAS/Sy
ZuLkKqIb4VkasCPHGM0cF9/p8kzKqvdWtzcnrhiLPXNCdd7CKwQKyVL6s4L9dVEUCIVNey0vPUEA
gIJt/9KaDDpD4RQp2soh40KY2DEQuP20PbKwtH62AsZvwk+FGpYNVs52aoHd6u75j+lsoeWwYYne
jUbEpGFsJqpa+kS7TyDbbIJ9E0OLaU+HYpZ+Lce2yFKVkQN/qwYcCtdw5W9pN1YuzjjHht2znTPM
n8pxwyVDGg4rn6QYrep555tUc6zByMTiXWopY4ZsAo8KeUW8vZWA/5O43ZWCFzpVktfvyOHGB20M
U3G6kFCYxxcsMl1ZZC9OhoiZT5CUjksdqJXF0dNVyiTry4OrebBUjv0oDQqosGjQ9uVtKKZo2C5q
gr/awBXBI7GqFiNnRC0SSaQF7krS8SUJ/I+Aonx7VrOmzy88LHMEu4QKsDY4ACwgPR04Ybs9XGcU
pluprR0ftK2eBjDV74vx/5DNRfgGMjWp0SoVKztkylB12OQb6NXzUQxGqkaxgZTrccWbNOxCI7Lu
e28Nqe2szzIzvBEbdxBr1GV7HzSL7NzCmf6p/JqczTVAVcxhE3jjnbpvTvQ5PmC+hyKZGCvyBMOD
fOQd+yjuUHQ3szDNyxT/p2CwmDO0emgc5oQs7nLnjBCw6XJ49EVP0/Hk1qs6PuyN+6yzdzs7jU37
F5nEfcXhF1H7NNAhi4JtdUW6SFRhRomANT53yRmAUR7ghr9dnF9Xq8HjNZYZIwgUZKScLTgr9IG1
1mmwXX1tSB26reoxoouzs98ZsqEZky2Clkl7fr/xLpfmM4mASlgKlsv9eKloq5gHodFYxSg9NasQ
ToQDVZLRfLVQMkECJYP5MP5XOxE4fPaKUP/qTdePLxWRAKRNe/mxX9EM0q/xrQYH7VmB8IT/0OWT
j3nhvY7qNX6QDFeUpOYmEYnepVC4jqP77/ohORc5U3CKfvCzS3nip/acdIgPB4jFv6YPRUpJF8bS
gWKItomlFJQ1Wmlfi1s2UKztlyA1gC7NTlSIF9/pRngscQjMKG1gb7RWY3eIfcb6FqRpPfK2AJ2D
h0KsaPKwBn+sEK03PII8dPR3GHmDUgZr5r9hOeCw/LURlGmcjccBIjcmgJdJ6vIyZaMzsinqViAP
QyzXXlVrfOAqLpus8FeMGHA37rXPz2dOcQ0DuUW1SmnxGEIGNsF/PCWXu22AaAmK7KuiiJvGr0iq
7Vu5SaHRitUspOXrE2ODkK124ckgnPStb722B+haZZwMUUcKVRNInCGBsYV70u5UpN2H2Y2C+/q1
Fbq8dGnZ9LZQeWCY+rVIjgH+7W/K2Z4OuOTEvWr/w8KK2Hg/APy3SjRS/sVEXidnJm+P/P1HteIa
Qh0aKfc2JUBvh9YcEC5lzJY7BcX7YKYtJStRmfT1lMnykAUjNh2OQsddPmK3GcWuZy0LRafAtcwK
7LRVlndCoVtx471A1thWqgPUz7GTUkRCmGwvygv01pH00GSaNotPuRgCbyLBdXmhyF04jy3eaWTz
lsNz4ljqkb1lgY7U37RquLjKud++ZArgvnq5LDMH9u9RNZqxoIx+FUgWZ0rl/m+Vqhxl2rZxmie0
pdhC3kprM4NARngMIaVH5/9Kkd9R2gy8IqoaBP7jyymrsmMjxix+v92x57Xk36yufozhFzp4t+/o
/4lla803Jt26VteGHKdApoJDPq2UfRriTUw2Nq60SO6Q4GxC9biykQjw9+Zf1eEgt+LZ0q3OmzZK
sCe/pQ8QbbeqR5nUYOR0oEMc6Yajcc6vNhefURB9W+2q5pqh2lx5ZE/EAlzmSZgM32Sve22ux+1r
iLPsSzVJarNdBO7IbRzUK/Gt8ha3IvkS4rYOmKh5vp4QTRK7DglPB+o/XoqeCyEKHixI6Hfm8sK9
GHVUvFrTJ/yUYiIHYT/6uzAnqfLXOnMNuWCxkDThfp0kOD8PuYs8UzjfaF8ZBDsoowu/dUO0UX+M
dotXHVEY2WdSTmdXs5Ki3B80+vXteT8RHycCLMf0eEi4OO4VMy/P2xEimB4mu9shRFiTwJhCHMQ7
RnzcL+P4sv13gzX/nCvhueLjsrXEoG/eWi513v2N9lUQ9Bj+8RrvKyhinF+u5A/7qZdEJXc4Ogxt
7yE1sMIw7X7Sma9v1wneBXYTAMXId1B0andPlECYg3JCyccovZX4lf9KZ61dpEKsWecQDOerV1PV
ENw7L/+xSuiPPW5BYpEBBam6Wgcs7AEQJxy/FaWGoBJflQOZuY+FsP+i1gfLK+d5HatfP3iEeHwW
1GkM/VQ2fqx8DUNA77dJElQ7tt+eVDEEaZkuh2b7iW3fwvpnSPVzMJNW44feIGewTkVzJE5wsa2V
f52y3hJNo64bm6VxWTdgrFudI5TFLdSnX4V7VCzQZrbE7GvWdm8fYcxXyHI9srR9toLH0WU1gmRx
goZqnGq+gaOMF1044CB+aGJjZk43hBczeOT9/mywuT4bD1NpayDAAhUr6K4khcdkpPcAz+zLm9ep
KNRnz+xxQ+zP4cGV7bDlZNVoLVJ67/zV6QxsCcCM3WoJwGN2WdCTPTQWGhHUWw8KK1ndgzGVHL77
sTyz2bnl8VYwThFRhb1ECt/HJVwMQ9Stcqa75CVOJud9AINSIt99wEMEptTm5Z9HgXYv/5oyW4qa
QE4zfo/8mGJbH0Mm/3PS8Bjb40dU/18oqNnPNLvfRS5dMT5f/JhQgUT/GIg/uWa/+YM2TTRP7ndK
ThkPmd99nhoYg3KhD+jBtC37JaEnEgXxDb3qBQeLMif5X3fBMJGs19Zrm3iOkZ96l+zELQP6mMU1
1gAJBxEHd1Q06syxnW7ghOJ8EK+t502jkZQ/yGQyST/IZcu98vYbRXy5eVLtZokkXjXI8XqAX/7n
MEdbZHN8+sFnMhUYaM3n6h4wVMOZbgV0HWN8X3FxKqm8+6F5gqLr3zcBRyYi+VqkWumr0sv4AQoT
yRGVhE1JwkgMZBXzx9Lpn3Ijs00b7xjv48GTYv71Mfd7EeyHWGiYghg7KycXOhUWSbJnAlPhwmfn
FBa4M1RTAAwtqLJWB1tAnRT/SySTUhaaDUykIkYGTGVFbAslJ6JIOzRRl/nPq2vF7T/LkF+oHskX
FF/I0fetowCXmf0iw/kFX0QO9xvX1+C50I5Xo7OUZYO7LKX5Xu0whYodFNdy3DL58TZQr3qbiI9x
x7oCPlSEX1rFrB6psZJ8jul184PeamTNkvYonK34X4R5Hw3W/dFxMsXRm7p1luE/YHlgZ9+4idy1
7M8h+tQWSAnzkYI+blj2D7hHn56PFgr36b1RI3r9wx+Th0ng4Khga6c2SYOTG7IEIB2pVGeWZSzY
z1jB3R/4qwqR0YTggV2gwJbWdg7QYALomkstGgaEJ4FJVBphZy30XrKKzpP7+VtTVSDz5ynrK8St
zpT48Xjnjj2Zd++9QggWE5+HqwpmyT4wr6dHEsDJXvf4+j9b3Wdm/pznCHPPyiHMwODSytzQf9DR
sIXgF51pJoqVePFtfOVkN0wOjFahhqp7xWI3E9sj0nakq+vjskvLMg0pdPLPPcnQQAVFOTghbsuB
FcM52yPKaP29FY94xchfIlXzXrfSZhgLCGn6CXgiG0muF9NvLNZPTIMUGlqT9g5Cu8USOxBfxecJ
bZd4kPmCqPfcUTfTtRHGnN/cF3CTUI5GgSOomzqpPXbRMqpFSCp6G5bWZBMXa5GG4rR8kv/SwxVo
z1XY/vT2igGPj6PSf9laTRN7l/+RpXy+iD+F9OplvchzKSUK27GR3JBehfEjeRIxE1CTtKhuyx19
wEiFfoXb7KHIL1tlbZTnc3pgv7TgeiOd8jbbZEmSvAQXykaSYyABo9Vn7fxE4MZRuzkJLA3+teIp
X3ubCOFlSR0M8qZ0wIbbe2Yh66aa32YzAmnNbXHjyP80eXslLB+Rnd56fcxp2U/bnlDJ0Y0zgof0
sp4cPcNvAsEzpvsCtddtrpp5fqNbhHSTTSxMflUAgX+2F1JOKkqp0ZPMghc9weDSDCfY+YosyRlm
eBDMOFhVz3HHVj+YB0RphFUgN00nY8nuTt9kItV1RO4l2i/Tob94eG1vBlPehTxYrgkttHFD4oFp
z1GhILhRzSjEUqWrxHwdD1nKCOOtsn1hGjKZNcQ8KPaZRPlge+3cDDHeMiKb+qQfUiiLWEFZmxNu
EQ4rZc6zx5BKbQeiTcdE36EZ1ClzyustAMDNINZ1pRvImB0FB8tDtyMFvNIvhIOMdDScv6Aumd4f
fbtc142cnYSkhh5DCcj06qWl2HroLs65J4wWuhxgKyHc3NCD+Y2PNS6HCdOryHyqLXw5fpUi4/hl
yhU240voaptCFSbVRiWrUcXThvdrbHEwDfdloRbRo0d/wzsNnab6aMezBinOZNPdwqZWZ+l14lB0
tgTy/TQM+nWviOoKyfc/5eDRBQiDfNDZhGOatfjcFaWMpAKw1A6DNxA7r8BWCt4IoDPfJTPTw6zb
1/JDZ0E3WDzikLBWBRpqK7XrS2597fzhAuwDVLQ5cvP90bS+6Cx+UPq3/6QojSNoOqAIfh5t/vkp
wpKkrtyItQXRp6RW0P7tKmGypt0M/D/K4v5WjH8c09VOnDJBNDz5T/dFTP0fFENpMUOJyHghZw9x
wCTHmw41R+bIcLoUAz8UMR1MkEyD8OQtgBk98K25fgZZ1t3kZVDuhmonhPl6lpuXhLIrKq+u7Kv7
cUfxbAIj4RjraBNyz2wTaPMsTB/V1iH7Ettrx9b6gP0JduTIKk3LFGrYyzHOA8grOnwNpt2a/xHi
s99Bzn1Qf8FXi82PmethHbN5GMB/tJ4K4bV6C7sA1i+lZ9Yn1tFXB9HLhEI6WdosfFCkM1OrJzsR
SOE6Y5TYG4OqjD0ETiCvPBDDnvpdZscCVk/bXzo7segg/Q+bfm0jQUtYFLtiWXFLnPASiM3SzP7t
KlR6H+sN28BkUT7MO5RAsUMSBJV32LfKT0PoTQx93wNtE62f8PsMEHnLCBBch9tQa3jhWB3Wjus6
j/jMmtfL0jHWIVTvn27O7C2oK8mjt8udn++CZBOiz5Kt8bEEzEEVS/dup4zkX7SYbWuw1cwa5xE+
vl3jZpECX/lAHSneKTWBTVvNyzNa7bO2+BovYm5Mo0a2Lu4zbmzp3oKz0fmLWccoWg6QXxs162a7
FH3lrqKGUWNfw+p222ADHs7gFRz4mXwIKrOUYziGrgG8cmt0fi/j81/r9qeHiOusX1XCuYpv1lPy
VhWyhDynxVhaLmqsoEYIbPtblegNFh+fVLKt9XNi+AS1RAFXZIcwVO3h+EljyhIOltyNcUytCB3Q
G/QY3ThvNnsDjCPh1VpY3dyjt5pQ26oZd9Cpi7fmVzI8FF9sngH+xPyP2DK34+DM1apwKG4DQ8zt
iP09yBYyOpodw1brYa4ZyF9nVvDHP3C+opISkSMayJ/Z9ZJ1zyp9tPV/A3OeJFVkpqZbm2EY9KzG
zNN3sWKUD2qaa9yV5pYUt9hOt6HD/XbQEoW1OEWvwLxwRyKpkZHbUx2PKgoZ9/zOzAeG/P8Uv3Wu
JQ7MT19g4F75A1P9ks6nqO7H/D7tjpFosW0o+bTFVTx1nwcMLFbYPoKuL9P2RsDTUTrLh4FMAO3V
a4loHCcn65Sq4fv5MQKO0o0dGLGXSFOf7sD4AyHAEMgY+3vfTczIe2bihb7Ss7RS70VtJVCSZLyT
RA87JMwDp2/h4ImqSYzmux1S35UvNhxEbIXanzDtFyZbBb7JFKMOdU+RWqx0mhjZzRKbjJ5SUKFM
gUR7yI4kuaiZ/R7seiEdzUl4FdLyv9HkRKhDVr01q6oBcJvAFFa2HrziYbl9TTtYRXoEGRsPGtBP
ShNgtiatOVryYtuTCzrJD6Grw67NDPhqU7VR4cn5osJKDqAic2cqEXGLi5AzQjpk5LzY9Wix45zv
7f/K4zSSFKrUTibKT/ITD8WDEOUSEpt+cbpWYR6Er1hAOpqY2S9eiJI4V9KAS1/wlsaXJUj4v7cM
1PAS+l0PcSteJiKMYzbR9/asILjw3/tFILMVQERMsS3252i0MpPWekfawbIKtfPOJp4iFB0J0YnI
eMQL6Kt5MW+a72TPQ0+z+lsgZ/+jPCm1z0oJV4jq5Z4Hl0sbAQrAh+myhBN7IE0Lh/HQDMrP6aRZ
dSnnkGfW228xbrz7s6ju8nTGlR3l31ZtBVzgoZVpejfhXGeiiD3yHTKcHMxXcrvhEhyZaHPwjdAN
ZdOFbHC+zacXct1m0FxbIshnNeZUQnm6Y8p6IGZ6v3D1KDFYk77h1lip/mMEXt6t+7I0Kaq7P8U9
7ZIfe1ozU2/9f+BMhJ1uSbH1xsSBRjwTUfJeNtOfHdkmyfnheAqBQcGTRLdKdK+c6Bx2m4N12z7A
DUwN/qxRQ1mquCrnZww2/5z0nPzyy7BzHUf0VJ4Mx4lE6/HjmfpdwxKSAXSyB8PiOGkZgIdNTp9i
FUS8nVCfFqBsO8gASNSLclEM3b7t6+TFDuZdKk5JQB6hYuBMomwCOF1lARmYA/ehpJFf8L0hwJUg
jDDkErr9dGBcnrf3+BQJNuTJ3wOYjle9hLEs88oSvmqssmNsS7OnR7kf+bT8BqeSnNlCg7+hJWl1
rKin2RzLCOhV6Umd98THpNvaBT64SLb0x9kOKvuEcI9zHcOQPLiTH/uOSVSH9KcUgJN722T5rSJS
MdR/HSnSUIRqO4FPuJSMDPjB9w3ZTkxxjrfxf0cp6b/OEvT8iR2qmj/HD10iU7jEomdDdbN2Y1P+
we0hY000u/uKIug2+eGzgyu+yPhMldXcbeUMK5Ox1ws2d2WtwTE2pdXYVbBHNwPvdk8KyUINUxRW
8XBAg75lVB15nRkODBlmk1wRcFlBLVbHQuajL8akUeZRAAyj7m53r3xLJro1hsYxh69SOf2y4/gt
+RBLzYrGjgPo4PD/lInRJhoKUcam2PZqn9vKJp29YBym4hxUG5T3ZCEqM+tpa5Bw+wOnHg2W7dej
WMazaZui1lWHvxhsZeKQjW1Sqg6h3h0f1LmNRKKo8miqp4lylReA9QSovH2Li8CFfdLK0Hbzy4QH
QLyFj4SqVjrtpf8g5It3DJ508GjrwG8jE/OVQWgnb9Q6nPzpBr67DNFXpZxNdgLNZL3cXeGBNO5d
NX8HKgu5TzgGs/6GjqaBxcQy8zLpNkErQHmrTtQh1gimB75plmRX5XWGCFNALoYUzJs6vADyxZDa
oHiEcNbUNPZY0hCvY3mGtGpbFcjaz+fel6i8dzusDhi0uE/QAZpZpF2g/hypv/bRo94MuC1k5ynS
v2oswt+ueR2T2jLvGMt+2ul5itM6+LH+GHM7iBmrqLrDGXQnMiA3R/btlZ5kNm6zdND/vz4bysW5
Zza1nrtHvYAnin4Yk4huw7m/yDIqtf17WVCxO8W8g20nUcbx8lwxNJmRZ9Frnm/IvoFXBqmnUXlX
Ng3VwdyBXYIfDotgZV5eXReidz1JnCr/+w+hMdRxzBZmNy+SAwFsXG3Atrf8QAhGEfrRNyOEZaPj
AlFOKZhjiGZxWzNJ37Sb8UcfOGlOEcydT+FZzShpr2Nx0KHfqm5NijH95UovHn+HaJgQxm/ZcwaE
UaUFgOuR6wFj/Ren9nSFluQ3lNF3S3vhf1shR1A6elXQlDeP2vpDNe986KxpBx2YqA0cU0lrMUx7
XNy84+mbkQ9MSEI9LiCIGymwnXJLx62NZ7nMLAIQGeg+VsNP/fW2mbHrkgJ+iTZI6F2jLHifgsDh
RkjbgN9FiR43SEtnVj6JJB4Tw2iIeJoHyR/cnZ0GLsa+bY5+1g1U4BCyG8OckVXeHO/chZ2d5f/I
odJYalYuatYlebUD+69heHzxcjCYwFX3y20GpPse3ZcLBMttiBLYRiNaq6IXOux74uJZsDj51X2M
4QRxcLNl/Hs9P9GkQ0t7Q6wha9iCgdFFGw+OTaBBzIJ6hnDijSpL22saRvFIUSiacdLq8kY8EBeR
7OuLkQU9db757W3/HScFj32qjN+QOwODpILLKcibWbjoYN2c9bX50MZimkYM4lYCA/oLyjbkEdCQ
GeJ6Bc4PKXVBWKbw82KDXJIX0Jd3w0aRl4pbGYR9iZi8IqjQBjCoMoXKVU/CrytkSJb/p0iEWViE
BhUeRXOgPQupbWFpA8H/YQFnz4o1ZWwPJD40EfRpFhip/Fxo4wVY6UuGEKqRc9BjkvdEJBc99r99
5/SWPV4y4dYxsLnDWoOq55uu482nmuNpGFqEWEVOQK3Txe2H+hySu7Yy4ysyY32divI+CGGM1Gfi
WSgfRhdUenj/Ue9xmJntLWpa+yFZNIIIGZzLpPencqnRMomB32kzPyEJ5vr5OKmdTH4yRfOpa7mT
baPzdCcn+a8tH3lFE5D9kyfjOTJAkARvAH/hDG6AEbjhdV8x9XF5utXBGP0sLRIWkiMkz9n6k/AD
Y4zDoC2zp3eIqsVX46tRJ6Ojcp/0s//sb4631X8uCpv9mjIbn68PSupedCtDUU8REt+YqxPTWpq0
1IJ4YzlVSELa1TKURpGHUyGqkGFF8KesMWe6skFzDYKXIwbOzU7tvWY1ncwaj12RthVzW3mC7LAO
ikf7urNEdzYdNeECx5KwBkgjEcovGxHmsmlFuGdHa01fph4OUucT+FX4M0orIrmPQeLJej2kJRKD
8maPHIbgMTzBinEi7nMbh+vNg5SKZ+2xqy2Bu9Dt+dvZD257ZfXpQM63x6r3bpJcvTIvOn0v3VbA
19yMEZVgES9vhHC4NWsqgWPALz68B69eWkFJE3SDYhIc6HjZ9l3NHSFYhdkylKHSBY9WnPjKyPFP
bUk56BMzNWdBlZ9qXey2F9LHDYMzC9vUs+6eqFV2YDLxpHzyKdBSQN3eDPrpj/cnFS2P0ACUsFTO
JwBikBv+ok2cxpLDNYenzdMpVzNo1IeNG8QbZahokFOP5gKq6zByuluqGO8ZVdYwXz05UBnLtNT8
Xaj3ComjdMjYd4zo70eEnTbQ7MEkpeGVB2ItnyxazEKXEU9joEApYmzZETCZ6nIzGllDjCbP4o66
mcHmmrs+a08/WuIiIgt6WM7Jkb7qUf8wMVCxFuCvkG8KRevUQttdL6+jtoOqSRq8Zqcc4KLtK1Qj
YeIoZnG5o8wP+2hm7ApOITgDLj1rHotP1VW7H4xML/UMP9vWQfrVbL5Y/B+1rYQtYE7eGIJeljIt
xxU3wmv9aLebvrRRWt9x4hNxPL7f2oxuVx3wTrHT7Ntm3NU/DYGgrT9PdvBjnNrHKcLtt1ybtLg3
Y7OzUHai3h6JQt0pZs6GZYu+CDZGi+T/B7zvUa7yveVB5Tbj/YAqUuWZCky5/oij5G/nfjzfKx4p
58CcvgxRF+NTltzb2Tzzsmz708qgJbOBO7UFCFnVhpS7y0j04ndbtgg59Df0GPj/zpfo2el25/rK
//RKIUrAP/zE+f1KTIOtQechGFURZFrHswpLdMq8ldOtY5zOoIxEmYze9G+WVvzJ6R4uUuoJ5TXs
UvmkMvr7TMS/GEAf5IG2r2aZkdRoNJso08KzkoYEn0ooXFUef1vbAtgz3LllrGXu/NiDbxArvU6G
0MwLcFA+T4n1XDCJ+sGQ51JGo8oHS6k4o17vDns20PkHTiheZJ8FQrBZaWYNKJkvN6E4S55oh6SY
VLs7k4UGPl/y7QIrLCXnD+PQiFZvknKfUQbOYWoJHmKAAaiMNPBzANUfRBtliIcOMWm+mU6KPLIW
/Lm9tLukswo4WTEi2HrT3bCnC1T63YcGf3m3gVbZ/TtvA2JgQFSmkhvDzFtvyLAb6tpb+lb1JZoV
Fy6TDUpWl6tfc+rfzPT5FyYjj31G9DwAmIqkb6qvKzW2W0rn+Ja1r1a3OFCg7bduHJy+WxRs4zpE
NT00dQi/oGOJ4nPH4zpn0LskelK35CRj8PKQvIaCfFnf0bAf813a00gIzexMowp4Lg6G7X+p5Era
vGP5CcBulwcTsyUFWullWjmrYn5/wy8uxAod5YbZQDoaaByh0D6G+74GX4sYrdrq3RzylKCbe5nU
xLHpnPiHMl8gHA2JgXLEgluWnvDnPv1FXgU2BGDgTCFb7M3PBl20dDzqlkXk0lHgRcI9VmEMuglX
WSoZ9/FbfG/2bRxf5GzZAjF4i+gIwrWwSYzKYFNF2liQckR63DdH5TCxEV8as6ZvLXCN2HkA36Qq
htKdYiO51jgateEy8JiZjcbdoYi0Ot31NE4SaV1N8KTXqHPzsJHs8SIeyx/9HwmQWShGHf055LCd
KSJLtYZLM1vm184e0KyRUzielm6JySgoPfjd0xyAkILFpNFvgju7wNGrVuWhCuXjLGEu6HabOLHL
x0YfbgimXhnux+E33qnKL+8We+1ec8NjodErSScMFIlHCM+01wL2WNnzUsVPy02Rug+vZY2zoYkK
ixRI8l94PxEJDiP2lXT9VGKJ5vC7vhyaBzPNfoGwEOdYJR/Ox9Jn50iOlu+kA9jwFz647agshfHL
FL1M4s/mrYb3yz0eVVPgFYlSrzyToKfFDLGlRrs7NbRjsiFv/2k/3GjL0rtpbpoBWVLxEkHK2/jV
GzeBWUhXUJR5B1Is45YpmalCCVElFSYJs1fxTTKp0k+kIz6G5qQEvENgc3WKL7pHU/v2FBxRdE1r
OCwH0w6C27SDASv7rujOB4e8yyZMijV4qIyd+LcvXfZpxjHqz0JFr/lob4gGqlckm4QhfSEjbJ0G
KHyzcoLnXXdIa+0CcGOoVy6Z+4i9zmXaWk2I9k1r2lHmuhGpTj+OXoD8V5D5H6Du3B1vGP33j8D+
38uUbVNYlY/cR8Wt/0ofe60Flifd9cJjNgf7jqRYr4lEq9LpdN21ifBrSzx8jjJxZT2zNs8hQKdt
I3oeMPX1WDy6H+KrzKHf4RotG7EBfXvMI961B9R5D8XTPVzA5/dCNhjAXXpqPUNommMeQ4UvcyZ0
PK/kgt5WKHIGO0B3eJTThadrCDjoWU1lQuf603y4WXP7PId2redxeXd/Qp9ErM63yFnPrxuhAw6c
AehmL9YiXRRcxNf05sFkI52/69DPbftFhGhp6h9sAuKRo0w1ySK6gvmaoOWukQI9NFzvMxb/wxlM
wlVP8HKNd3EF5TJx0w/oloJkmReJMOF79PuJ4PZeYAUdDGWQqoOO1yvqMukXDmJuqKePPMDbiJA5
/Mjfb94vZkR8ooblyMxbzS22RYN/nFWs/kxeVp18ppzlWvOcGiZLwRe7OZbO63D/Mmvv5jzDdvM3
v4eN2nsJ7w+v6E4u7yQXpU7EyeMI2TESa55gLaL4XXgfoBRCQQbZv5+kjPgzlc4q6dBWDM3cZ9Fj
JC0bE00UNLpQjgrQLMnQIHQqXq27tKTvnZMMwi8alGdlrsdgUFahUDFz6Y82Ctt5mHXfFUIHYCeB
foi5+7irL3KGfoPojIcMfk6eWUaN7UHzN8crDFZx9qztsoWUt8WF7tKxBuONMemVLcS2ZK5jqrkv
EwGqy5J7j7ilmtD1AfRG0y/YR9m7jwLDRXIeTyPo+bgafA/s6nI0qzYOdgmN3wD26jgzFQFoOKYE
6aPAKWLqp9krTB2B+nrhze1WheA6V2bsynuUWwdohsKG1OU5n2zH+Uja+4fNo1iyuZpKk7mIf4an
yLHfGMzHOG077bxN4NJ/D09+2C7MUpQB43UmrTXXjT1iLukOtm7iSbu5oJAiArC1LZrDr9MpdOVm
Uxy85kt/KIfBTeth6RAEiP2YmMlmgvpxrDIVoTqglPYtVYf/Xk8CpGDWFaH3d24mrvmxab98AnPf
5S4vYxnMdBQxXYl0ANZfz+AriPFgwBbOYMD8DlYjCxvwSiLGgLfLlK/mHlP4s2bz9+BYlfLTajlA
+4CTHgOkl8/tlV5aIf/HW/C1xzL2uZNLRIqHtCmB0B0URxU4GBug3VkS2EbWqqy3F9W1bz1rRgvS
iFkQweEgLxucBzZj7NTNvU58hyZwNPxDMCXIhUstnXjT42zb1GdRMbNZTrCGu1i5SjZ69gqhq5MU
wPAsARlj3XfLcrs8V4S3RIVoGbRmHJTe4WX5z9oFYqDIskW5hsvw8arQ5Oob6kAu6JffsjcvsxDG
ODeDDOZtNSCFtUZRsmBrwWAXUPvE8SHnIe6v019B2bS8rnkeB0516jiMdj33qgY6RV604+8c/yb2
yMngE6oPXfZyWRYcDEsiz+i1NTXaa7IunY0OfZM2svBi2v6dXgrP19hQOgSH4Y0U64Y17owx41J8
4PcBmpfZtQkn/Oz3s2PtRPFfcVOCG8rG9yUIh861Ox5FlgeOuT5QFNcjEShLHoVUI1bR+C1ln02V
HEKErooG2w4didSQREA6Uy/I3FnrlkQk3LZtgvsz3NlZ2DvtYB1dr5sZR8lXcPP1u5+Z0F4KbFSY
4cvR3mdfcQp3hrdIBhW7/Z2fBwJSe+61N7fyhRbigFY2SrAN9vD2PC/yHHGfA73KN1MiSqnE329i
WYRtCHBJhjNr8+k+9xPlWIMESN4YOzgcsc1Vl4uTxK75gt0za+YLw3n17dHo1pUrEo49OtxQcIpQ
3+RsfK6ps54swyWILVoV2e22IzwDUJgIpZ6/LV+aGBpjLZEfgqHuQrtHVPyJNrRZBZ++sSToixT7
rSEqxVL7cFLRWXN1B40VPx9c0suyxcey0wOb2OxCHAMRR9Hk2dTH91PhnHHUY1gF2+/2WNO57xuA
s95IXwc6M68Q4/v7ULLv0HT9wAEJu8pScBIWwFkE77KC1ODZCjA5t2synlVsJgry8XGGafldblVP
HAMCSGCA7dSbPXnDmXpFjexeN6M2P3WyiIoqHaMmqGNXr9YQegjB7FIw2vaUjYdPs0eypyyYGYZJ
+yxvdzcUhpuAjgVUQm4uX7OtqR34Qc1UNPl6oYMVa4pKyDesl9xvbsf9D28Tfjxr+miLPIoiwSzk
cjMBo/m0qux5H5oI+Fbjgu5SjPNaXl4x/HnBd+Zac7UGMYufJk4AtOZOWI3rDxCst5jQOV+7R+mz
rqzbxpUlwsognuXUpXAmwJQv+VfPVTWyhJclqF9ztMfMb7vlDIfFP50gkhj7Bs+aABuDpbR8hpma
BSqJzXl5PvfYG58+y/Ie7y5+5/itP+DycCiGFi5dyLwR5uPhg7GaCX1d6bxiDHDxO5s95JGnHxu4
LmECMuyG3Yj29PcKfL6kZJTqA/2rjkUvRrmBLdm+qtkU5bBeNLHfWzvhD6WogNHExwmKUTeHGX1L
LOFqo7JDPbZeHnaGaEt8t+ff9lSakFhrq1X7oKMaOy60C2KvIcH8S2Pa1Me1JePFh0GIclVxcYFI
kDMHTCgJg7QUZ+Hxd7jjBY1S/ANcgbao8RsX2x/qiAZyuC77/tlLc1K/RTcr5qJ4tnww9zgQ0U3r
w9lUhKkZIW/LNIZU1aCao5DEyAmozwb2OdQ57KUY66LMSmA90jYFn1SduNs+tmDal7Nt4Ts800t6
n35MwTvTIXecmF0EYYn3GIUetP796Nii2yiNYqgip8FkpAuorwzvQ4e8ovqrqQpUEibghpTr8qVb
S8CouYwyz5Emx1M/1mT1F+XL1fvlw+nzhBK1bsZhfUWMi8oJkYtanYSwKwa3EI6H6DR9IiDtwxPF
wvGkC+TGoz5J1LsXxZS3oiGIqE4w7krV4MMkVg9i5n2ulaAkyVz//SgE3b5KZV/F6czkVg4pvLJA
rM26Xl0BlsZaVZAfS/fV4Oun9CtTYY0JNcSqzg/AiHLu9DXEYTbioIGwphQBEvzEDItxCW7nRH54
Ocs4Wo+USSASH4N0v5NJwYRJYslegFlsD0d3rhUuy29sPByEfUBwi9VZpNTb3gVIw1P9oGgjByh6
gilreOmkK3hBnaxbb3zUpDfHWWGcNKX5nyH5QA/wXWw9ngmPAM6KyJxJdARfcazbW0buplyqUhnI
t2TJmug9m/mlz6xqRg77lqSeDw+1Re0K07/0YBgj7RefFvj46+l+/CWppZ7aThPDABmpNjPP/Y5j
H2L1A2JIdnsiIDL4wCBg8MmROXquuoBI7TqTnLpBs4sFm9kP11Fr7UjPvUMaz+8q30AK+m2ilIu2
tgBufTA7aqaJJ6E8TMTWXh2jleVXr+eLW6GbnmhyZM7V2Ke9zVpAjoSOdgzeo513b0Wy9AHGjJva
difuYeJwt5aBWNDoLmjpfJ1m0wyuFLm/T8CaR23dD/X6NBD+QCOIbRuciBR/8f5kdV1phQwe8z87
h8w1RRCwAeTFReIGEwKlha/N/HXFAI5cb9KXthgWmMZHyVN+6aL499PQs4CItc9mnHdjqIj1BPBh
j7/hzr5nv8GTk1lkF0ic/+f4jH/2EN7Zx7GjNajWF4+TCdT1XJtt9Ya+tUkDZewFeQ78hUalcBwd
/l3d3OahuChOqX2u649n9tAs3noo5mZo8NBn9w1IPkN/NrRlXgBwdHdNIZwwaf/deQvt/aCTrCNr
NfXBkU3k0wbrw3eh178+SrWGfp40uxLQF5RAkeQ41umk0vCKxqIiQ1881fXRlJ2k8vbogFhBmsAq
nQD7vJ2DrzzuREk39vfKgl5b8lYpgPNrU3WfG79Qf5wsg+v2m5/5vf66/pI5MhRKkNad4AYrcwHB
g0XIQ1argYRPuTec8hHYas6ann16E2x+9Nmk3NcudyGw/fA6+RMRK9VEML6/Onq5xBj2O4QbQ2/v
3xB2Rx8E8HXsnQpqR5HbHFIkJNkneAw/mk2oAQUsjDN0ihun/e8TRlQLJHNDiBiSH/Gi5AC+IrEr
DfYxV7Eg05mIeYOGNMesET/k1aVTUCGv4TQy0x+YvGl/J9bp8N4he+u7Oyoxh3gBsH7QuGMCsnNH
XmNrejYAR2C0OZs2zycMHOoiL+rKBy41Qw//sWIAFRornq2Y6x5US4xiG7AQn8Quq2/tMW61UvP7
GMx+0caTvqPyBxFA3LOmvk4+xtkw7Gw/sffmwcH5nzZNAp5EbnoHmXytt6PWi4TksqXd4bUnRdvj
3I1Pekb6l+Q4MXbi/eS70W+vMioFR3g7I7F32AM8uU8ccKDRtdW7e3Qk6p9ATICZ7Enqy5QYjTDz
QuLhkVKzV41HzUPI/tpnOGqAnU4NoOXkJuE4hojoW35gvj+9O82y0FZ7vtOmlgyebVaofsn+dRAa
E1iNjJMdKgtZyg2+6KVV6vU7baxmhmTleE4A2ZKkngxZcx15eTXdn2H36L4N1Ucib0h6WFQ6apHp
OH1IQs6ofOgNCtEWJxXNkjqarEk6+P4NCJFUeP6Bu0+aKJOfhkcugicfRWHFOm8Pm1H19kDHi59x
5HuDWYekROr0L2gA8ph0gS2QT6brwR0PuOhGKBbA+htRwocWQn1C3pl7Br3PJTpDujP1GxzOROYK
PCTSy70JOzR3ZL3H4IA5N9d4kWRfvdlNY4gc/jETizbp48gymBnfzaey0LJFcn09HE73lyEtqczH
qEPluRyFvxTb2mPFNS+FqRsFSjj0pBoLMZCQcaCAgsmDeToCT0lsDU7KmKIjKUrkFMdoOo5r3Cpz
2/Wph3wUDZh1snLoLYIyNIdSM2+M3zuhk+pq04ezoUSlj8rhZVBTC4yuHdA93QRx39XQoXas0+2V
k5Lbvbilo2IRCoJok/ohHaEIOF/67SRd027kcmE66k9Q8HkwLp/dGJg56KuZ2ryzqa2MQgXxCfiU
dUBix0N/5F7I7JAi4aljWIx8j5Sn839XsbZr/xsilmftDvMEfakNtf0l9JMyRJ0fsf/k8nHXs8oO
+QziNoyvTU0cKqPDhWGwFb6G3s/9tFhn8lHEciewA1razrQfeB6wSuU8xQ/AEucTaTgll+cpD8cH
IS/gCTgAVTd9IrNOUJazukzfnDOqQf68ll8g89BH3LoT8MCwOS34Njuc9zg/lcKsr7b+OMBHJ5Uk
JRGoF9kzrfj8E+waLCNegD4zcXeyUInO5FNBa667tTQOP/gZCLuDduVOD2qhIa9GghknT1OiwtKK
sFA7Y2dsFSMhyO8S2UtloMmLIKhDQFgvXTy4AhBLITgqZ6vDd75NpUwbPzeLKBK5JAonW2hllC7j
aUj+l8FRHFmXPUzHAS2uRFj3WFnzmSP+eY+bYUga974/C6dkO+i0CC31AdRU0hkAnvEtHP5RgCLG
oW9o+SmKwfsDu7ZV60OUdJEzZ03biR53Gz2SAcrdQ6vgPgvyCpD/m8RxssA0Ew99zWqlI8YLi/6H
PgJyvFtOuw8Fj5mRh19MKgBw6i3vDRdr0VHBRQAMbYCzXuPtSnPjKInKfxtXcgP+7gzWq1IABP4b
TPearbzX6vyBpbBBZg1eOi44Na8UQD0ClH1CQTYfYm2zuX8gfoihUgDjAdOjmmOn0M4nc7z6cTKu
MTOcJrd7Ta2nzdz0K1M99KmFwkgr+crC9BlYMn2gKYF365juBJBR1l2mFnuOwt2PvUYPKJMzl+9c
OcP8hcWdkgqGSvj0YK1hVxhqRd6NLxMbyVjU25PGRG2TgZ55MU16TLPZunGXJDzxpt7ZPgzfaEp0
emnFBYFQaUuq58C+f7z86GnPnqvxPC4pZvu4tu0PquwhNEL/ZUxRH/4G0hoKKnq76PE3IBbwP8HY
g2lG25jr4sEQ02Hr7hBPgiOOzoQuxYt2gE8ARNSBF9ErpufnCj46XxYP649jkAtLOXGiLdRqFi8w
LvYaE1zonNTxZGdGBH2ZvX/8zrMtig67AbKBbHwx+4U0PEt58UiPSFmqKF85cXWZE5GP+qod90io
fNLkXrrUzOiwrXxF2JAMw0hzm6sJtQ8I/Dqn0iEPQzKznX1YW8eG+ZwfMjw4juSJSxcXeF9gOuw1
JN9luKMUYuK7aLnqManceemob6NV4ZStEBkqAabrXohG9DNzupnPXddjKm9pfcVQNBcHpyArGNfC
8rcM95IZ2YMw4RfOUsoFZx2sb/XvJV7InNwc9jk4QS15c6Wo93xJX1lYs9TcEjpodZimJmM4baG/
hvf77++1PfzQ2cSWOOu1nBuBBFUOGIHofxxt8jBGGW6QfaY/z6ivFn649QRiw8Ev/p+fl+6fIuv2
i9LD0p6+hVPzAmboNJivXZCDIaSRwYKZiuTSJhhrXjFl/Yg3no3KCUM1EirxE2gCpx6HZn0Y++2R
OO1ib21ZjvynirnNDZpUORgHIFih3lrikqzBrERkT/098Za6xMc4YtQuwO4oOrGWTK0YfW5oQeez
q1po3Dw9mfduFMqo8WafyhadcKJ7df3Nd11mSu8dyCDYlUAm4K1PsCJFhaWhD7cXyU6GmraVedL5
cQS5yvBN+127jiSE7lpm7PmtThkl0XcJZO+PkWvKl+Z9cvI0+maWC/2cehdmdDT2E1t+Io2nxgMj
7tcPRip+0OetNVkHFSyArtNQP8aGTB6M+UKYpNthGqoIapJCD5Jj7EXf9kjSJF4rX6NkQFF4qMum
AF9YLaKfuDZ/JlRkhR1zu3lEN7nKshzsLBuu05eYZDZNBfk9MQ42F11E8QAxPZFspzqP2X5cWCN8
oH1g1LXWMzf9feieRr76o1bT0NP9moQ5wS/AWtEJ9fVjpeXbK9SEq2cEnx4vqwsIh4bchQtJxd+A
eK2e4cV+qCWduHdOaxM1Wr3T3RZvuhLwA1JELhV7YpTcxKYlAw7jweH5weepEi4+ADP0GZda6/S4
DV/RhEKBcDKQYV6BQQS8bslabApjbgG7TSKGajVAWTqCwy4pI8pl56frub5XjL1Z15/pw7xUkpEb
DOczPt/+2DVKTqgfjm6ajW+n1b7N7mNq5XWzjp41fAhPEePrhS4hpXBxbS3Pj8oWiscQ5+wejncx
VLguuYS0m4Ts0alPhwgo9XsV8X2094LLiVjTOYP4Y1qBF9Fwg9Pr5YWZ1HSKG3f5/uHvYPnm4c9Y
zS11nON4fV47ZfgXYQyOOioeA6JPmiPjoOwf3xDf+gHxgOpcZuf539tPJOS1kSa2M5ftmz8hLVzz
5gIVov2DGxuT8on1ay57LovIs/c3ilGZNFzYAcTY5bB//US2fzTmA/8EZQ1U82r/9I3KT7SBeT5J
XHgOyG1NGLeid8tokeQHl2J57Ks6acoRYEOUNA097d2KzW4UFNsDCx7bvIuPPk+FLZSRgxEH51aa
MzDyU+kDWsHzCwtSGiFgIx5y08ZS7a5qnyskkPBaWfnOo1ur//nSr1tP63xdIC/e/cYOHn7wv//K
p9yXyhO1rWYTkzcqymeTQPtjjqw4cKep1Ayyd4U51q7iudtq6+tCUhqyuWY1GmsdOcDWub8PvOi1
JgJhgBGt8SjRrbZhkRBcTFaXtLFMKz1YUzGwt9HZeZwkUMfESA9ifSvf0xYAF0IIYyr1MctgGFo/
Sa95K5mICLy+qU3kO8yBYDcRhHV33tc2d8Knl6YmesEE9mrWcNE6lU9gYA1PmhBw7SByuyngtJiF
OuSSisA81Y7wdAXMuQH1JRo6Deu3KxJZ0IS9X4FaVOWkHYJGRav1s9KTeoSYtYmlZXzU90hqCRvr
hMaWBGdEpZQRso/ZiQ5TxNDKp+vq5H4/QDgkq7g3h0DkByPdfFCBRXh90bbdxIe/f/I3+rW9x0sG
zP55AMCQcOQ7LZJysHAp5A3L7hXLK7N7SSf6uyECDT72Xjfu1XmX0bKy61UWiuVblCyMtFeRj6y3
eYo+BPptXbhTLru5sn93dTG6Jnh3srqVYr6fqoOb3X6zdN9MJ3mAFZtliy+MCD0M1Z9Y2WjYmnnA
mEGA1ProoF3NlBu5EIgS9z42thz86hS48fxwl/G1et89vVUSs7xXweXX+ewjDUovLCKBwwYzPZu6
DYdKBqPMZ+ztaTwj7Dar3GL6dUMsHnISG5mx521WTrgjSmqy2Gsz3vCFvqRKULSXvQ91d0Rj2MmW
Z4yK1pzAXqWSxfwwLgxN/lNUezF7XekPWltDqbuJBpzC2/G8l9lsw4/kYMc5g8yRf0lo5p9DvNjp
Isvo00k2VHTaqZXNjIw8uUXLcRXESNGEsRHmyYEymhi/dhbUVmhqOChhu6BuDHAVTzhau/LtGwYd
4++Rxo30rHKLFxWHP/WOe1Anhqruk1ClF5MiaA1vSuIpNKZCPAZjX6Pfmli+/4F1nibeiEspGS5q
TTpIw/VQUh/oSufSctvrovxXMyBwas7XY7oSbEjk2924F6DIfQNyeFCflRc1/ewjyzIX8zajCh0y
FYMknBBoqoaHfVBeTXGVA++NjJgAE6VIjyDduY9sl+DaONExckXiXiP/Nwc0fOBRwlyd3HVllKhQ
W6kAy3+Xe8P+sCCyYVxS4M8f8nRI4YOQ1Scc1tcTNKIlYiHYnvfwUTjSugi88UZRnwX8OifHFOOK
hPNtXtMEZBYaEJWjjDKfDJBIeJPENbNRwjH12CdX7jCnq0/DK83+TVWMoNBZXE8KGCkxPLu9IBJK
7/vBZnY49W/NVEs7gsLyUtz0wJisV6AhWxrwZZKxbhZ160G9RKW4wcIi4DoA0V9MTHn4l33Ps8jG
emSNodiWoNQr/91OlrCn0rr6Qxf8afpJkFXxdtYcSgSY4hpwAt005BJxbfoLtGdmc3W2+87l6gcf
QHDnxTHk05GQ7upsYePyR65SmASolK+SzATz0l8cobA25aUm7A1E8feH4YRjqmUhADB7jONU1Vyg
EyJ3NmemtK4EuypF1cBwoq6WxKdYhM7H7laK9dUUuU0KSJXQQtQTkXRO/ySVuwweYECQpLuA9gv8
Lps0MsgvD/omKuD5nJRGvS/41t9OZK6rcUaluiN9TXG4v/UKprzcy6TU1FAlSK5LKlnM/s+Ias5Y
RlbpRKwtuaSGHUb6i14lEo9uhfXpRduPmx0waavP6IEJU5ZG6ziu61uEtgEqSNJHKah3kH3LgHIM
y3a1NmpwOSEdR/HOU1rZl69wNIj7g1oFcFl9IiaEaSt9kXg40hHP2P/SQ46BVb5q5ujxmAi8FgeO
ULcQex5gnEfdf7MNp7A/TZmMgfGZ1LU/ShHo34MfDAYDgRL+sF5e2R6hSE4AMraiHpBULlZzXxIb
egQoaTGko2RALj34/rK2cCmLYs3o4nteRzxeOwXB7/duEIPQywl61I30KYJ2qTaWis2hP88S6Atd
3KrmJU0BEgO70Jx5Qk96hqsaCsFWTCcYh1GB8mdrcmbzD08rvqQnF8p0XFwVRjoYS9lizYcm6AvA
5VtKsduJQe5HKB0bqSC3SQdbsKzvAhk8tXSQ8SqjaCOmI4UUC+n228sr7VB4d+oV89tvyisl30CP
SM+ZsviRghSWDekvboYCpd2xtZaTA7VW9sfjYIhARmcL2RbG21nRpTriIR5Z4wRZpK3REykKoEAR
xPEXUQyD6sBZcu5vaaiXngbqVjwhMPFQ1rmQIUjgdJ8u0B7mZbfJ24ge/kWIl2TEEoBET6cm+9ri
ZPxzva4bFUcyj+SFT2xRuFl7xabnckJu1Kiufr4XzlqitxtI7JI7XW+QXarsqLhYqKrdYKAt5SUJ
IyAOmWRMrV+rhyyXWkD1Zxue7t8U1XlQT2PitIm79fIB8sy5iTfZsj426sk7C/GEWsGbQ3n6/4Um
QmP0LgPs2vftz+D9JanVW4/XiCCDzw9gHS1U7XkvD0aNS4H0bJvilO8faLdSdM+QtcIHZsoB4NGZ
i716ACtKUebmh8E8IqL3GbeonsSqbK2cowqPkZpA9PKAKBve2Qbr2PDq5NHPpdeW7LyXndK2YAq+
skMMJRc7DSNRr6G2BWRzzuverTjJLx7irfvy1rEKYyPRS9jg6ktkeuLUgdh8FBAP5OHoOhP6Rr1t
N7AcWBE=
`protect end_protected

