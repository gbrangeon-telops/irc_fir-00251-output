

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Ya253+37kdInKtzN3pd3f0ykMvIJsSTHE2tRr5TaFzMStJPqyqbq8G0/aCj9umOixPoTbod1oPEi
NM8lNQufqQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ZnAl3olUb+r5fzAKtbT+P9BDg9y9NfOiCUm1R2Jcpt91ydHcXeu+pZ8D0lxHNM0CXXGhs5RFFeCB
fQNmyCQv4qniT4fHHC3wrH5hPwmAH8kqSEyGt3c0SvSsHCYTeXhpF8Chp2XvC1WNZGYymRNjehFn
t70d4j3zNeEsu5WAW84=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
iKnL/TA899sfLGiFOsNtfsGv8lNgBNaSxC78jj2+skMz/TodvgTxrRQVQ/h/L38N/D5FIkKYR4II
+olODWgmPzea4VBkBMLQ7z2XenA/M8Uvin39meT5Qbx7/ksgG2EdpyOtsmAvmeXZQgf/A59DevU7
Mrm0rcVFwLpmjNvbnBOl5iGpGgx6v231GzIUzFEiOeCx1PkRai2IOZKE9lG2BMKHN7Bhsm6JH1NF
XhuV8OyupD6h/Fr6EDMMNZqriSBB1MM7btJKN6VC9jmTT/Bega2BSYjqAkfYdUTeyup0UqEM3znP
2BL1mUmUOgL1/UMAmExO5qz/A5ddH+Ai46kqhA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
bwfblhQfYU7J4v01pOh0vYth2hZJ6Xlf2qmEYdxkErcnbM5+VpJUpwU8+A/bDOJB4gUPbJHCeAw+
tmj2AabGe4D0Pf/UukkjTsO8eFOUvoPbwDwH6UV1AKQFszUSN+Z4NTgaKs8pxWumW0juNgJujhCL
2ChBu6ddPnHdB5HG8uQ=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
UTW+eKUNnZFWLDMo9paR505jK3kaKnyoN1JMPNm5SlY5iSmlguqsHIHMaqSHkHrYg25dIfFqsLa+
ygBhaN4bDhxyus3QZ9m0sw/aVS4ly/5bNlw+8ePaK1evrFFnRWDzqTt8U+H1O06G7NfpkTmeK+am
Q1esOyihSrmjwIiD3aw5SiSY1J84QcBDQl5D2DAd5uRtMADgrmEFzx9Y7yHel0j2iF6Z2vom7g5G
7K31eIbiTPvCntdYde5+aN/nl/kdiT8a+6o8fslm8ZFdkfMYbKE6CsL8CG+5F82TWbIzOMfxbILY
sXfUaKwgi3ZDGoeeudit9zXCRYxReIG0hfQ27Q==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64272)
`protect data_block
893idUBbBc+FJ9D5seJoc4ktPk3Zc6YHoQzltsDftdKHK3bRlSSswo4srwWbT5L7BXChK/BcAcNd
LtUx+78zxTGz8Q9bnTIo4b7egFEORJR39s4IZIB14PE7PEjPTg42VwlCyDHN6r21HBSzoFsfwpDG
P/wC8lypIPyP5E2FWFlJpwE3sOMupfw/FQiP7rM2A/JuF2WST5tFY7DLueESUm+oHebIMjRwPKES
OsX7Dg/ip7ScnI5Rdr8VhxEXctoeKmEYU5lXmTBJPMB90Z5Hrhhsvh67UtVOwOpXMPofx+JRrHlc
0e74+MEShT5j6BqS1H/Oza9mrCZpt2AKwwFcOF2OJ8D8R7lWI1uXZdqMWHraSb+4DHh9ToYZyge9
AiHy4yMMf5Di3cgW2sXGnj+hivhWao2Fse65mccvv8w+zVaaZoKA861Pv9Yz2nOKM4GXJPk8RXN0
DhCt6AU/uTCvo/m4vwViLcwAr/iIhO/ZfGiNEcs0SQqab9DKlQcMbydhD+q+lkZvnxrZiDhDw7KO
j2uBCIsY7DR8er+SSlhEwjphBNNRIpd49+pjChiBLXZom/V90i75VIpN1saLJ/WPNkvqhdRWrGRu
8ggJJyQkOU5sFwX8GlqyBBEocxww9OCAYaB4BU4B72kBQ2lyVtgioUfTF5N9zJZXEjKvWq+zgSZd
f8BcydLVTo4PdWFYLdrl2eB2a7CrTmXFPPU67IHQiWcOibyTGkce9lMdGxWb/q7N9/UuQ521K5gy
9OV5g3cYVGSXCoudJcCb/2rDYJNXwp9FtavCo/vN1sXaxoDnxBi7wrrHrJ0xPuEhSw4EcLZEvq8U
AVqxPHz3WyWKAeU4E/vz7d6P4kv0EdD2Tyx29ndqSsLSvcmx9y3lqqf/e4vaDUP/a4UcMOBCgfIu
TAzmLLANFnUYc2K/SQn3Md9vWhh2DIx+xk8j9fS50ipGWaspKM80wQisu/i3t0VImICmHpLOx6zp
uHm1zvHF4BLs0VmJnsCE9Ko58mG4pSXB9/g2oX5BQTNkcQhPTev4qBjGOatRtXEXp9gOhONBL8wY
IZ1kpnQF5yK9G4/y8s5WsgKzGe6prpymHzpJxU5HOOEC02dc4vo+aQIKQp9p8luLPnDUFkJ/d68v
MbcnmMD4IYq6YkhZZmAzQm0c5wQsnRjVsyBgiT92+N2jTnG5pCOTXcCRg5BEHIy+CHHQiJt1pyYw
JSjInmLjt3x+EGFhdrfaPqe6kdSuy6fKktKWr0bHkueVp95+LRztjiqyCPGQjqX/QEWXU9mgRO/E
YxkQymQ2TFU0YvxSqsftX5fwodRvGG0y74+ysVquWSCG/CtLY6KWw0lnKOSo8mxPRkSige/H+1mw
01GCIGcvn0PDT4wHC1mebFw0O2+4TZl4rJ0cXZB5O0vnaCKrB8bVFA3uCx87WaEQJTI/YQH3Ht9o
f13R8mxxYYlWH9QMBh/3/FbdckQr97rnm3iYAENR9r+4OUo5aHpeWAmhV0dtuamKlP7wmo1/esL4
b3xL4uhvmy21Hq3ysrlge7fhVvipWlXKVeXrIZdDAp1kSC1Pr070jdPaZa6wlXVxinf7SRLMEWvg
O0JJ3gdgHRikr4sFlm4gLSrgYvhn0O0rxjsev1/uSRAD2JZDk0pmXWUEpUFbi1/WbsPQCRtyCWqq
dl+AUfuRrtFEqpjhjayN9VGGkslI7PKCJ3xYIWCaqNTzwi40/mjXM8U3YhA04lYNtHHlZtNNeMwE
DTmT4htGR0PzEI1WD5OhR3ubfrBi1RzsBZWI7mD2TcbaCxDcgOEHTxNAazNdk8CLA1NkeX562u5t
dm9E25awhEXKvluYL2lq8pPoYiDQnYY/+CPKeUqnI/TcqdewREohHGTiJHE/2ap8YRIgSrjFSrLq
uhrZi2wzvjq3wocNVFBQsLiCz3Wn+VVv3bjuEjCprfBe3DjsgJFCCbK/4rFmKcl0FDFuOkxobpOK
Ql+7bv1U+0o6Oy5n+xp1fQjdnBsVT6Clewu0e95vSA1k+au0zkNfHOzd/XITlu6C6THilhgnlUTe
deKtu22o9M/OhocRXk7U93fLHhh9SFzDBpsdjuJg+HfGRq/G958HADkwaA8u8PIqnteHHPU3RHDW
C4ddJAdzdL9cEQLUdSJvh/kz0gF17LsSKxb5HzbmrEtNt6up3YAs6vBkjh7rcNg/x8JPUGZaFUPR
U/0LQTu6Vwr+pHEHQI0GyMPy4HwC4qgAgHZxWUk/ujK3Kw+6+QsF5NSuUMxxRzzed/x0CEWivz/T
jvDz5gyEAjvlpyUtCMQlHqVnKBWCecqBuhsk41i3L4iplcUTUjyJrwRjcoX7huxQcdMmv4h0A08O
0gEg6/jwlryXIEGEq9Y8BGVia+kRtFI8r3nQp7nPl+wfluVEOGF0248+fd3+KqOW2ew3xru6Y68M
OuHfyGhThiGqaGJDHEJHSVkq188Ko3pvTbZdLbCLN3uoK22NCzjx2yAFjIq04fNlwqXDrZPxa+bX
7DA7zN4zXAagNjp+sMJlthVL+4cY0V8BYYgPfx/+9l872lzc5Q3mSpOvO3jU9kh2CsQeKiM6chFr
u8oZy9ZEuWDZJt66sWaGd44O0Pc7el5IjqrRZ+/f5UTX3nUhKruy5u9dVpTFsh1bbpZEAaEmRKOO
xpUzbyBTDngfm1yCwha7Jl/IPfejcV9HbY2E4Uq3iqbtW+c9c3TrDnekGbsD0BZiVWIBio0+ZlQc
hVDyNs8T4tEVoQ/a5vlQdfW0fUWl0PvAy0CLeXx7Au1NKVAnYojBBMmkZLFKfn1sJwPUy3X4h7zF
VNGlRFJWFAkgbtHZlOo+7sd+mNseP+SAryMJispew4Z6sbWhht3MOHBycQUkZEFiqLguNoLNqNx2
L/Qg5rAXkq9tlgETf+AxQ6OHEhYtMg38Bi6u3CK5jtneptUXcwvdAvwQ/WaIGNT4KXEU3U8OzrTv
2Q9xED0EB3BCxjqyvYPWJA/MLMPOLHzzh8OfzwisPwRtmUtaYagbtwTEAacwQ95Ppfmh7lRtdxUo
QlP8H0JWR4zNcgDZn/rDk7u+QdpsThymeRKnobuMXP2kGS8EGfRV/kueGTnN9AXm9F5S7uu3nSVA
IQIT8ziSJ+6NydmGKtkxBirIRNZcwjgr/3QDBUbkT/8E9aqNClTOnYNtBejEvam8vU82WPGeCk4/
4/iLmP0RPQCWGOVfXIydX9/00PDWSyQXnp8nQyMZlqcnwWlDgJ6dfZxlIJYY9GcqrWm/uYn5l4rp
nulgxBALMPQDFtVAcoCc5vXAQE8d70dy/cED4y1b3WtId4jDDVoVp2nphBG9U6AbmADq5BfokxEJ
oj4egsvJq5b0uSFoLfXQRdPl8KkOaVpcQiEkWIcdxXx6ziBZg/0HBZpaDd17UE+DE01pHLHZtfoB
hxD8qQyJW+9GwfnXTjhwiYwyfRu0NO0Ce8RPVSUvIkPUfL+8S91NxjI6enLULGkYuPVkz36Nkht9
wZiX6NyeG32oc4JOa74p5a4ROVnhcSx1od7b/qKK/GKFVLL6sIgPfbZj5UCj8UJXlwaahXwUDtC2
nC/bmawfZO7sfJGCoIcCnoI3a9DguU149D0bFp7AKYq9JrVX930kyHXNsGFNlZR4At47zw0IEam+
Z7CB0zzreg1y/he8CdSxGDjIlTnmc4KF09HEkh3LjKn6GJwh1BSjJvuynzZI3DlUcL/yx1BZgHcM
XbVcA4WWx0FPfzXi54ob9WkbUXsHYNMB/uVlvRWNNDx5NTn4peXI9Y251v5m0ilavlayHbYniEX0
USO/IxwEAE7n71N4f9yJpnKmDIWzOJdkR/cDUG+IlyBRi915q6uln5LHsZ2Vt+/1wO43KJSvtVaM
8RMX+Jc/etTOtPUFcAe3wXxPuMQksqAlAWBB+yv1yWLRRDKbxx5T6uHGi1Sf78N23+P5C4Znbxo9
APOn7A+4de64cjjjAZ+sSxdq0dXTQI+apQKobLak2Rp7g4oWH4otYQBTxBzxK2aGiYv5LEdSPxV/
qyYvEpnfGtfwAM/qNkUp+C/D/EKaPcUJVxvyRSC1WXr036gYU5rqN5+1l5xlpcmaXMo9zgZPAmOq
khCE/9WnxEO1tGRTK6Y+U9HIKvctMHdUnv9fWsuE+HPG5kfUtKes9/tDSONPwiSh6Pt0jJtKumQH
CphgMZAE34SGfnEiPWMgkWq4ohE86OeI7RwtRgV/JUxptrJyApDpDl07LJLf59F7wPsfd4wNCCco
L8SmKSwXbS8C3wZHqMHq7TJXv34c7nFOtzlY7wfurKAoIlsEpXI+3e6nHi8I8vtUDQUB7DSc2Fve
8J7Y+Vebf6SISRcuAFxu2hZ0KM/qGTB60nDB7+sngxs8SMge/xHINJnAoUZK8kblHJvoqTChtz3y
123VLk8qixH41VBxVV6c0HRxaGcsDM3VV77wh0WmbZldh0flnzk9Jm5VeqEPg/kwRFtMNhBOKThO
fdJ4YidIKjl+FydTPKyF9qQPDdqSYD5BmoPtbrSGa9ExaV16aqTSybBdma3PQMOBrdOXjUbIB+/d
ns5eFlI7NXqpoEv3QGQwqfs6/Fl4/xz1dWh1SPIvW3HXSKDalGqTe3iJxst3ckV5QuE89RLvrxR/
cen3a/ducnTguXCbUTHu5AfiE/csIJvaqit0F80uxr37G6ESnG59pn+4HfJc/eeJEf/nJS0v7Hnj
Ql1pT5Kduoz+73Qiio/oU1ZrVxGUFdCZC+Ry7NrM9JteEOL4olHRen6HuTLxP2fZof7o5m0KgFQ4
gRUWlduQC1e0SxZ9y4tHH8itvqNTKgoUHpR+DKmohiVWpfiJACT7TbV2gE4oofoAOJj03R1PW0uf
IBUPeKQExZl6Q/W7Qloc/c/k1sFBL3Zu3P+rLSTa0FGay4v8Bskzea62ML4TQnzBPrScrmKKtZJ2
aO0mfld6EpHo3WSjLOeY6hWWOqARJhgE00krFfWmD3hkvNdZV8rorW8BeZCKesE6icR/4K5Lmk8v
OQwZmjvymscLqQb+eJOZtp4S5ro4mHjQkpUE5gGiElZKDmx0CUieKk+v+Wq9Nrw9/GybpdOgqAxM
n0l3Vc1UDMXuW6V6zxHnCDrz4Ojs897S1pEw+cQ+esXfJTOtsT6ba87L+dgwP+QvNhUBbLo5TaXc
rj0Prr5EX8r0kEs7DzizIOoOyThZTsV+iA6nou4qdUr84UYPapzJQTGAlXr2T2YYnREfIJhKEnKW
avTrrBSA4FKlbtheuLvw83Rxo7pZL4ptu52auQWQdmDmsNMle2w3VE02vbsT2shq2t79tO+O1Ubb
5kPKb68nZ9ORQRdaT8U2PAUNhQbnnChwF+jrfXr2j0IB79ZWjGgskzPSk3KBO8nQBCAAGqx6hIIb
uZZgE21N9RvyzXoaDTo4Mckw8ALFROdWcMp7ln0chWuUsSnoO28sJ9sZtUwi/P7/AebmXY5+9aZm
tQIBI0ynHPo/dXge+8LMnsFpkm+YdmAkT6GDh+A/rSoB3QL7KlCkWUGguaObqX8V3UAuiCA/00zd
k1OOsTj0Jdirlf3AAnhaiHa2PXAB8JebIHpy6Z6y62HyqnTLzkp4B2wIrPvVK/ECZLFmKc97ycye
NtG9AerwHe+mHG+VQvt0gInJ+JnYwIhqfRECum1UcGxfHp7kZFkY0ZbExfyzbaLPCZjWpdwbQlWx
kTAzlL22DG7WWCO42aKkdH960GIVvrX3bc+dI3IQyzeyyi0jrAbqwoAsMaDpE/L5/GwP8pMyA86+
JTp1vrXLI0IU8U9cwK6e2cD5GFCPHx27YEd9GF3ta4MK4BDj7mVuRjqFo4hR7Ek7TLrc51Qrw3ha
DLQF+bLTb4/nMKR6VdzjOYx3fIYwNYUCJpbX4CGKxLEVj35idje+TEreEda2qbqO5kmJE+OlnJxD
PKTnMZAaZX99kNxkgvy32mIB3/oyq1DwZPxkRwSqYYr9wzdRkzlY8olZkmJxC5Iv0D3kQYStsHvf
IQy6tpXQ8RvNX6D7u0Jf8L3/z8niJU9xuT8kgCqElLN8SlrM9k2VLhapfo+gJ6hv6/Za8jlZWeQI
GZSXAHjvaZMCC1iW0aglbzz40Hn+fqSdXgdrgiH0TmF9za8IIaWTMBYBBceUP+CkZY5aibnJmaM5
P0qO7MuVtUUactAjqAJzcQuT4NnihDjGEOcS//fnjuIAhjpzDOGqH+rtLWVUhsMRfsdsfGltLngo
pQ+4Llq0qv5UReMVy5EZT1meo+tx2ErYUZmQmlODA3fT5izIzzaz3wuW15VEDff/l3CBcMOnZSR5
qSjL0is2cZLyikHul+tSvY21hea0FXQHJXyvtXDEadCVFt8VV8vDW6RHb+wU4bemaFSII2AJG6w8
6pU4TzUTe9vG5ioFTapJXHjkkBH28ssBy3Cn1kBk7ya99fq87/pMFwsHR3jVFqbeuE0QL0ZUyt2r
2FNZw/czAck/f1Qy+XskG20QigxrMy0kgMzk0eMnVxaPxdzmDLPNKq8NCGNv6bkrbGaLfV0mAyEN
col7/2QLdItOeFdG33Tiaijkxz8SCksXw86nFWxqKdEn7KIEOcYO0IEnAf6Pwm8vCOXU6SW3CDzi
/vQZHK59PoEU9lBrbeKiYuvEUt0ts8DcER8H/OpKl4wxaX7xbSJEeptsEhspKScBoPJVlUm81+PN
7EgnA9udAEe5t+RFTmYS/qXd/aO5QLZPownOsGpQyqDRiD1M6zMewbS7K2DnExBbzFV/yhLK+RQa
R68vj2gdxIA+kDHoE1gTMmpabyPWnosL7UxDk9TuP8JFDMPoQLB1oa1QxLITFhCyo9AivctBV/4j
wU9J7GIwogdD2RXIEmR+1BB0BZmxij3zFf/72rd0/ZadryKsbnoXdaKvArM/XbdFgyGtbT1/5H4x
8OPRKCeZEibon97ATOIpqpcpq5eGS57Nsx32FrcmVMDsccaQbCXS/b9LZ4Gsp/eo3Khz67XpadkF
H1hWjtqTLGJ0OUvpXXpMFf0Ab/hJJIWIZgdCqir45qx051JsBWS58s2v7JsFGL1NXqyPPkolxFKC
dSgtj+7NiU5yTIvVc/cl1o+cPoOT7KqKed9Y68d8Cr5UysVkcZRsCynZtpQdpAVwENLDTvNgoj8n
0U/wJ8M/XqaW4bW8WhyuiWT+rw7F2V2SiMU6eEB5XyTnaglOkcIkeRInkTa8iKVHbyMhESo8VTnv
EBkiAW2N5Eo7uCpSCVflEY5H8m5Xj5EK2Bc1Vp68xXSXDBRTwUqohJ/fAujEhR4Q9G2MFqWtsA88
qN8i6hsFZv2zVT98ltBCA6x/z7jJElJECZGpIQcJIeGIg8gYr0/UMwKv+T1oj5SdanJXegDRhynC
0aWfxx80JZjMHHMN+69uwGx8n1fokrao1lp6ZL6f7CpAnrq4nnNExfePLYxGeNa05kzf/u62n9cC
FaoT+Ggd1EKZ6jbiIIh3fZE3CigSBxWI+kIal2P7NGJD8x/xnNNeo9dhkPdcQGOnp+OBgfwZKX5/
Oci5ZiUlEBf+c8WOil2ej+0yZdaIYXeF+BrYo7C3AUpxHdn4aTkjPDqNLU1pSWfYdIZBDmsrgbcH
uIfM0NzPxQP91a9BJjzaDGdK4pOTlogaIR70lIvsjkf5tI5fdbrNeeC2XkWdf4O8t0d5dR+G+muL
1U1VZx3HtsnIs4d5e+Lnk1d1/d7MVK5AaPD93aEMIdRXT+IydJNjitl4yy0ktsIXFNZN0fTeUXBF
UIhGhZM2KN+wNn4f6t1Qlh+1VdprxuIR0jiin9pmgiOmdYiYNt7cksso1yI9dE0lZLnXmXzIYOuq
8GA3tadw9WzGW+o2R83zJ6FaeZbwjstuEkFyYPSKGD0kzE2EMIajKlIvZa2shIb8qusA+b7eVa4Q
98DLV4nQjqaLBE3uyeJ7D6452nugtCq9XCkL9yq9Pp2jlFS9iL+yBQ7qrY1Z0dc6JcmpanbUB5Ql
uR427/6g4jyvhKPzi6LdQdhQkaoXnv2tMu4dBxWn90rWUkMp7/oWyZFZQXYhV2GKipBFyjseErJY
/KRDQkCZtht9KGcNQCSXQPYyEpDO/L3Kn64Z5rQWSEZgSoLLLmXnH9RdWJ4aoThZfXYoxZkMbXaR
e7HkXCkRdfp48TUlDB2VuZbqtPmIuZy7+V2h7wYsAQBQVEnoYi0NKSVx7DCxqFtMuJoAgjg/bqgq
mJEhQSLtM6WY/ACVwGax3pJfHXihTI6gbrVFXobEdCcwdqLtWu+mTXCubeSkZkoNR5MD8YVfRPxp
w8W2v2AJjDlnYn5j5NHeXqzDul2QWqFfUelp7J48k5/FK7RpSpeMsOvmEN6l3KvecdMwaI+d1JDv
IOgo9PQ7biHZTz9M3u3k2f+Nn+28dLjt0nWqQMzohpOokpuEQg1z2CpMm1jjYK3mGRO/Te5yw3wI
OQ/A5yWe3+vncoTBw9fxxUo5luRSNfIRLWRLdPoABJw/hb1OJ8dCsQyvp2RXr1c6e9A21KgPrV/c
G3D5/6jPwSmbBDrXfs1DFBKobXsED9kGsNGl9vjysDv/NSw2NSecClWgvpIgLpTJAdrbneGuxqs9
xXmL83n1lturcNd0beUPuF91J7xyCRDTdZ5juiv+r2bI1xziJWwyxhs4JGtj6MMAnZE+a5L2wh0e
W6T2hK5xXjnnEYS+zXE7QVg2N3F3SJ2ny/gj0oOwYVW/mNMrb+GBRDIlNSym13YR/ZTmqyNJTo53
z5yGJcPDcEcEbrp7HYiSnqo1Q7+CWLvPjPiWCt0QCGr+gMSiqG7HVgnBiXZeMy5H4cDVwcBMzKYb
Lk0kzEvG+b/XDuzgrzz0By9l0KiHead3Ksn/9vEjWpcXc9C6iqbBRACPovcnlBB0ea6aoghtAQzn
IMuPg714TlePdkQmzoTuGMrFfSGf9gmf1L6ppahhTgwYfi1rolTh6fV+yoPyf5Q0LTABi3S9pWKH
qd8dv1gXiqAhKl5BCp+pl960JvEwAtlFaMw0yr8lGDxYiCgb4i1kK0xDbkYWk9DV+YEJHhWoIZgx
ZJknCIZDEJml4xzEHWV/hwz/u1h7fUXRuF/XvZ6pI7hGSJf7tu+tjYYBL21TgczBKMj8UknEnS5H
LM9Bzf+qiKzEmXl/U63py5htA/NYYCY5Q+kAKcEXkBYUV61xwZQM9zgcVDyJtsdDM3g3VAd+Ywaf
VU62QR/Q7oXVr0q3E8kjBQI4AZbI9P4A0GxkGO5gX586BvhcDamu1Go+vH6GgveTPWxcFmw31roT
rv4JsPLkq98rFTmCXgzckWN9vnYaDCIjxgUtxmXkFb9nXk46BZUDNKsFSuk/iffSYSFmpPrB5Ee+
MGV1UnWgjCDB1WiaKMqEaeqJKrIynXxaiIJjVD5vFBFqOp4XvCzWpEcu9PYJu2kmk2GGqDAn2NNq
5m+5f9xpAtHv+mRTSiph+J52ZeZRcunjSErVn/bYQHN8jfbCIl/VpxvRDRJkJ85Mluh+uXPQACU2
23mp9rpnwOLiWbPXBvwsyx7nmzzzwDTNxcBcL49ASB0RSvoAj3lNUijeovNIsNDwM1jrXeaEDKaj
0MOql+EgVnhSuIsAKbQ6Em/BwLnptFv4F6nPSnK44Fn/UPV3x1V1gC1uJbXz8o0Rk4Qa7IdgqcY4
Tgd6ukzUNAjehBPF76L/QsDvnRi5WBiaU3tKy3jFf3F8OWMLwqLvP2bczCdMHe4ETKyPtzT308/d
n/H779j5Lc5wGVCDLai9zPLoUIumiUqrsYPewPpt9ZXQkzETnSsctpbpHT4+5BqHmvaJZIBLs8Dl
4peWGKXCCi32HVeAQqDig2Iz712a943A1C4+VD9DSXAnl+nDEfrEJ0HikNrWY4PiVkxUxGP84ADo
ifpNarF4ImusLwwaoj/gsjFGLqNaNEGDJXH1FjQ+RCLiQwLFF53rBZ7sKe9zN2sInJH2n28jJEsm
eDvAK6JIIOUZ/kYUKfgFhps5Q3XCMzmmYjHxQUIOPt8M4Wn5ANUsem2A8ncKeNUcJG66lw1/xLZK
iwrzGroZQAKIUegXcgrOZgs/Y2L5VN6rQR0aJJYI7b3zhIzWHWWrfzv9CTkTYcM9vID2sNmSwP1h
Iz4nfkD3YxwU1k+hfRpq//AujfAnHopd8wa5tSCRJ8ksCyas+tM3zetdI/tgxY0G6JhE/zcUQIhf
8tzTxfHnlX6VKZ6ArOlAd2HlS4XUZzSniTD9GZTeqtPVYtt0iEBC7PCRXPWa2sFOA7/xrAyLlIHn
YF60aORG4t6mroAHUItDn/fbFptEmrEvs/wHadkqofQzSTs78abyHrl66ZA0vmKPk8VBqxZmqD8f
HTQzkESagpQhpMbbecghjnUhqWvuuikVHRDt+7Y4o/5jbKWtNu4+DHJo43+Rc36oP6AqxKjtPIYw
gwxWTVhGBP1mi0ORXH8ZFjqlPn6lbxEbqcz3hMOQztxiWj7ebwnK0GoggreLhfcvHFUXj//YqYhr
QwP8TzpuTBrGnxBzyFvTqfet8cBuAw6Qhu2pxtb5jIW6b1faF4dW2580or565xPyjNOnwsPzmN/O
slzNiSGGySq7irE66q5yWiFhQQC5ma1s0cp4nWrcNKsV4kbf8HmoBaWJhiAlx37rpVBbM/xHrZnb
5vEmvitBXjsNwp6qFGZT0KL7nhVsHKSmnxzFTq024FYV3ehzCtwjQrDuLuKR/ZzBe9NdJDV8w/rX
2CcO/IwXuHqBsg4EFi05tBtvSVXIZZ+lpbVwzQeLNzWkNbooe4kw/vl5sEK/epPhnllrmWY5s8lP
mJCkPB4Olq8sAXvLhLOdFr2SC2mlqBgY6nMfk7lF0+OuJuTvv/133X6CcRbEEhyOE199KyU7/fx4
iwSfqsziBUv8xveg8pkvzMP7Y1V3kO1rDOUH8i53lFqvvvA7v+52DkjvKetzkDvEFKL74D9svyPH
bWTVhclKpi/8P94wbOajV1loafEDTzLufl8kUpHjBx8ub5BMKSfl0dZ3jEllTjV5gdkIF6WwSOie
tQgB+R3vtLck/5WEUKWqXQ5zFIUsGn+sZXL/VvqP19vKwLDMPfEy/41HBkPenWYO5h0MlIYi0Les
E8WleKzmEHDdGei24/Pb9WxukE9NhghAPHG+oNJz9NO/2S6AyuFSVYFJFpboZy+nkf5xyM7rysiQ
q7VBjQlM1Z+ef6o7wVtH04Lp7b1FLuUv3CcJwihqbRKHILVMxrLY9XICp5xaBF92KZS+cnmuVWoP
rucp6nvlVMsWCLRdpMF420gFgwshjDnN0kICenBYoLM44YLiruPMeXGGvbfz6ICbZcbL8IweQPU8
DYwJ8Ptce5phxawhP6IbEvFrDSJF4fXmYpQpZJs21Gq2idxDrXrUQ5MmLJikbtiQLKJvhPG63ADw
eSiug2np6qE72fcP+CrEK+mAJWo0BSguQeQDNvjYKyidhXEBCx8hRt9koYPLtuUvkQa2nYQtD6cw
oeDEnOXOgPubTXRSUh4ep12l2gxCs1q7SWtYIiN+YrR/qLdNcTNX3GVje4UuxDn3mAlR4M2H16SU
D1EaHZB+HPkVaxS+7ig73obUkFxCtjIoq/vmnUzD2S4pmEEAKvn3IHutS7w5voW4IRaTZ+H91LMz
7Vdo/F65fKYmSp/8QGaak0MUHrH1k+oqT259LgEzTrKSKVuvO2rOwASXoB5V24JzJKQ9xqTpMe/X
DsQ0l7ES7RjnUxtQG5uBrBUochJIW6jaeryc8ZGSPwkdL104lVlOIyR8BTWQfD89OCX6UW2hj+cV
LZZ0J5fI9dYut3LQtYjMSq7e3vQupfhQLvt4aXkUzayJ9flF/s2gpDaJ3JaeiNVIIL1MCKUkOIm1
whgMCkJX/jB6ltijFazFwfbPuwNj9m20c2bhyKCuEl+6CB8/w0cBE212ZAwbK1q2rTltvpY1SNHK
5QpfZB6RXqC07xNjMv+mNsDnJR9hAJEs26XyXQh3UvwOGOWwCAENjNHa2cfCAc3HUjQpvBfi3XJy
CerJdDfYvDOWDavczsSH8BfYkkSR7zjtZM12A//K/ubeqSuqGH2LDgcfFAWtvrTjzAE0f8BFt0+y
81ePWi6RtnH7qZci+hJ8ahqbaTqXeJzyod3XjDCvXDKtHneVOJ9DpHYDvRz9rFQabFGLKUVCAwPr
WYj7k8Owq5JZ4YehZsRq5As07rLu99oPRGsbkXCwdw6abJQBWBCq1per5STRQC+ihnraEhmW87yI
fvzRsTG6zjpjUi/63+14eXmR/1xNzmUie6gctDADpNo49h5TGjPfdZfOSGTN3je74zCZeMwyOWXv
qqGAoBXwawkXuYFi0jN4TcXumdf/r/FGTbjiOskDYKDNEMu4FVVB342fLQg4x5Ois5GZUjLiPVZ4
TL53bwMiIK5ZfRQKErhvUNAKPtjnInQ4gDonH5SIyIa0hkL2ZSZd3OF5zj8H95GQQxzP8q45sOWI
C5BthcnHyXAf6T0vlgKE0gcevQisXq/5CP/8rrhwjqqxfQ0ZV7UsfYyR+bAuxoYIW0EXhjsqYOhe
LaEeEYPYkwT0RuQAlAvFUfkxgbtFqjmiLIH5HRiRBQ1st43Z6zdtdeQ+1WmzPI+iqI7iGzGhiOZQ
/1rosFWgWlkg3P6Av0YbJDdXH64W4FRfisoIpyxHMFhfyAKm7+GX5NFM07Z55W7HSMqqEJMuknZx
d5A7lc+DvGdlZmDO1m5znNGulLsduHeoSSm90hBbw8cWyAAPyiMGe5OBLDEfLXVdnDe9cTiFJTwR
gzHEdKSVYw6ioOS3UhutfRAnZz/sJ+beIr02kfSsF0emsIGqFY648EeovuaW8suSxSo9qSbm4095
Nko/dooUXihbLHoW665tNh1atXCJlCKar6KaRoqr1tb52F8U76LfVcdgn8PrkoBSdUBWvb11bJya
2EAmP+lG5UzFRy+h/zsIJS/LvQKk12Xgz5EFoiKPNoNIfn9x9eP94E2+0FvYk0qDy88eUlAs9WWb
ZcXQ/O5ZofImFgYUR5M109fbbfPhPqJ+8WbrBsgbkA0yWwuPuDoaXnoxS4UOvepiYsI7w67HjOfX
vKT4c9aamESmIypVyjgkj9FA3YAl71mYwf4jmkJsvANL1XuY6SwosIvv5fxUGeAU8PWLdAqd+gQH
Jsl6Q0H1Pt8l4b5FEIf3AEzxz+2s2+AeDrKTVEvnvnkcoj38zlxg0wVTj+x2Sh91pdaCxd0oxVZG
cr09aow5nSiGLEIrCLA5UPCZdRG0vh8DQfy5+uCDWTZ9g90Gf7HpN+VN4n6EUtZ37K+RESFo+0Vh
+MrSANlcPnppACPgoGAZNDggBMG50y6dVRga1lP/VzcUPdzAQ6l7k6CiM6lKP99vfQuTPQ46rimz
/69+g1IrovPyzE1FBKvDWzszYS3seKsXReEnLN8cyrw5KQJL7MlOVbqRl2UnGV66aIJfOu0/C2dP
LqvGQ2zOxaj7Vmj3lJ6gWsbZ4mZarL2Jxm5ouJ8H6PYfegrrCLSp9OKNAiGrW7eiHewNXdcu6yK6
0P4Cv9YhRNMiIpiTxuXQwFhajpV3/k7VtFXAMtkAqxglZFgBlJy7OVp1Bl58ZZplCiGjjMmVComp
9Q1maPfPfDsyjs0Vylt9V5llxSWX9fDXZRgpkbOJD2GZBmEs7NapvQHd+lvDBUmhA9Ee+lBfW+k3
gTHJQt44+Upsb63PCaJvDm5+W4pfSIzCtHVmjofEB/tMfydFsF/+yZmwnCK2zsdXWfkHzEFhx8mf
Rq4rUfV2ZSN7rTj1DFErXHgLRdHm9h6mG4kFVx9Tbvqw5OfrVL9aW4CfMe9Yiy7GGKZWY4xR1eFd
UNWA5NewmBM3KQyVxvYiihaFsR+vDYJiTMBpIQwztXHRnk6zDJ27TMruzS0sfqvF6yMsyhf+yYWD
RudDKLBP85js8v+s9FlyjEQsuC0BLfnt3VAzo7o1jKLe0wAg67YihEMcoyUOgzjyEfnYfds9IFK1
ZaWEoCMa15hxRaLYzzrU8O1HHulfUc8i/dGITgQ0ymVrHhSnBvjGzQBcHpnYJ4m9iCuu0Qat3uxv
xgmxcHMZqpw1kukswCQVJ3p2CZ9XaVnWrPepnNTuxqBJEl+8nbbZlK8wyfUshpff7jggF59YtdF8
8hByx7+sIj9o/SLrN2dxzuPWLFubQL+ScKb4GzKghq4qHo4OL564yEnsxXg8pIYUJS8xKcUkyJ4N
5F239p0rF5UiEnrBcEM/RD5T3C4KM38HPdu6/317bgs984svcJBK4nQNans0usZ1ouIahC/61I6r
PjV8le9hUnsKICpwRqDLqZb/GMS9OeohZxsy+9w11AaL6h54EVDf4ySV1quMQjF12t7VCLs1nhmG
7g/57kWizJq+HtI/w8xE3ptPzVpEbx+RjJvkliyMFuyrA8sqdhAVl10TOlbY7jAPQsTYSc6LH3AN
wOhiIN7Inl5PhuQ2hhaQhWQMd5bzlNBLXmklxqHbtqVYkvxOzwZJKxI7tgPFeDUdWL85QJBUlxS8
ghT115fZl7SNRPlvD18UjqOhlQe+iTplWt3qF88PBtaXon5cjIu29hObOfPeFRw4wMaeOo/1c+NI
xZMmCwgt9/d6gndsXEW8RYkRqUyrC6AVinelnpql1ptC0Qt6WmGSpltRo/htBnRfgAiPAJM1EmFc
jDN49fvZuF6cxwJkt/VCBS8b0siLlUx2vZprj5miIxVRi855Fv062DnuLsTxIIfJsHSlV0xb6C1B
V91+Yah1ShfMXlQLQBo4xEHs61ZPW40vxhyrmaq0JE4XYXQLjK8cBYsVascFtJh5PeoITvxYGjGl
t3CgKkCDEilpYaDKMjgMYamrm5Kz4sheclQJecyJ2mUt+gdN8KM6mba3xHmyQlpPBkpmtP07M0g5
BkIVyy4MQoocLBKmuwvAKjcT+lNFTMZaLXAUihdAtUxOMvTHEIQpJSpqt/LFUqJf9MPKpyNt24ef
SPYM6BdUkPm2LZZDke1lMuWk9clD/wn7M3gYJTkL7VKz0j+OC6FtMuIq+S31TK15UNHkUx4s/ejd
jDafiM9BeSHz1hRftUWpCQ4Wi/K8gIciTlekuAIcFRnPRFwJdCKj4LNs07vPA3YPNtIqvv/PrTfo
reTYrTov9WsavOyVaTc/wyraWyF3tQG1YXyoRGjf0KVLTvNRfJJmnmv/6LA/HqqsXCZ+tYaYVZUJ
dum+s0tUcGHxqtZ+j1SiovBk4pVGWQbcr/B2PgKt4TWdnMeq9Q0m4ASTxaIk4LftwJQCiuZ1RyLO
T5bvVFhMGbEIRyXgqDOmtTU8qZBdaAc3qe4KnIgfjQf88O/fydPkm/EweVZSinmFfPs6RymJ77ub
02kgEjPSGQDDwDd+NiSCv71JNkYfGPt7fjBXADScg8iMg1e6lzgMcUFF/6IlA29672MAvtj0GTjl
2rpivjUzLt7mmOv5PopdhDIeLoimmyvrXjASnPwZibZSfu+p0jCXm1Bc0q7shOAOXR7LWM8XYp+W
uFv6l/ByIvErr+OsaHLwan+DhSEuahGVPIBMsMeeyl9bzE9bhFqce4AYNjB+TAtYkofREbAYGfRY
mRlswilQ8T9z37DZsgT5JSYaNxKeeyOyGDXPnAlYy6SBV+6BMAFq6IresibwJa9bzfrcv/ZZgEA8
k9sGuDef6Ds09x6u1cjYMouz1Pek4qh7DvoJjvWe4QiQk0XzvfHVkh6TNwXs4J8x3xAtuj0/nWk1
1H8oXNesbdBTruqgtX0vdHe1HWnlqfywqYXns/7J06uwu6DZVyl6Nlq4LexkgwXbR3DjUEU7Jf0b
wKJHG9xCnHQwSBzIm1Jyl8iVB+8eEmgK4nARPlHKmcfu8UoZuRB5vxef3oU/iieG4YJwAxVY3EI5
m9sFeRxL17wjZ2Knt2wU3xh51afODNVlXR5B0mYmVnJpS2mmLt2FfwOrQ4QiF96ugG0uP4yOwAJz
U/+AJ0Mw4gtXmyYOeGjzLP8PEwsHwmCHAuxf1DCs8ZDPoV0NPBBYW/L3GemVFp/Bmvp61kCJ/lGc
wKfGYAQm2uXIp3CJwQm737lpDkwqXoa4CBPXQB1vyfa6ezbkakmzGnUP8yDw7w1DG+sE9LalE+os
zv6mfwVN1knueL7kjp2zV14cklJ4CMhCdn2Y+E13uts8K0kCHjZM6ZuET5NgGucg8cftTNNuwhea
uTkBv7XEYtMp8Xh7JaZkG+AfeMJ/gxBG6zB35q6Ra4V5Lk6COaSggKqgCpBfE37J+Sj1CRvUMrdT
z3ONZjGQy7D9tmWhz+ju46SFhEvLxS6qs9Am70bcPgksofyPPnDAynmDIBswqSU/c26HW6ONKAhQ
easeA7Z2mJmE2fUM3OkWDYFGiiMV0fGtxd8/h812hWR33YOKyCBMwtl4AAMfBwsS8vte7ixP0V1x
brUEJkFd7Q+0xHOjL5o2FLNJo2ZMw+9pZp18xkuE4erkA2VVUCPOJp7BzCxPIAKEchHPo9xo8qpo
vAwQR95MKi3YQLdzQl38r1DkiWxxCd9+sBBzKUpZtygxngsKATCrI10my7cW0NceWRiumHgnF3Vp
MJQyVeu2URU5s5cKm9VDpXlQeNsWA96816o/5plAW5iQMSO3DkkHrYkkvflfLVzp69sViKbz6I3n
PtHe73Lk6Zhds+jOMEeN0N1Fmm0lBDL4MPN2HPMAMxsVHyzP5dYsqcUXTv8zOdtAbAj48IfLIHdb
pdm8bnjmJgX3Hp5k8sXn8ubJg2TX9dmw1gnyGFv+UMYKHyvxrDLyhmg6iZfXLXn8OLwvgGP5Ysax
E/L9QZ/VNM2pr6jwMBePdEWaZYHab/8FvrgtGQZ8Xb6SAneZuDoccWNKg+kXVDZFYlMEPooYbEO4
g2k4+o+x6tX0omwaT+eyRBXgRCsfSYrYa36y7TaBtJ9/EfNOSyO99EdycLOaIY/h9Dx3URtiCtsj
6kaPAHJo/+PH8MWIXH6WQZTqcupirUwVVVNcL6WhN5oTx9Is7UM2B8e39RaYuPjqOzP/bwZX7+g4
7x12BqIiEDRiDta8t/fKBs6x8x1qPcrESJyADw/fl1fMF9tqcS4OfJNvJ5YINeu2zQrRqlP9UiuE
Wj7VuITSfGAJCWbizKlijLOdfbj/TJtsYTGnpOE+I9Nsf+DEMARw5E5TsbrKdrsSN43L91TlgmKZ
Ld+fkRCvWW186f4FZ1hpquY4T74kBKZho7NUKT8DdAH2bDJR780aI/ySIuI5dmH/EEKnDcL8P81o
XzcFA50mcVV0mA3eZ5clJvG4v16EaWdsFWEfQgba6xgH0Vl1II6j2Cq5FRo+cquZjx4kMDHZlmLJ
1lJ2OBmR5VLFTj9apIRvl+bDlhLZw5F3nOcUy/uHv50WuPSsVD37ESKfRpzP3sszlf79Wrs+kaXf
GFLI1rZHbpUDBfsoQenTjSL0cU00g5tTIi/ZFKV0ThCtm6goPzqveknJ92NCxmB99dK3s0rl8w1o
gtKafIKKhoi9+LxpccpP9MUgDi1FAkFT6hCNq9Gxkn/OrJyOTznAMxDFYhg9qB1B6F97IFYQSE2o
l2ddaB1EB8yFcCtN8kE2iKAFWVJHbGCWbdwXz5eBZJzBx9Nms+Z3Y9yyl8qQgjracpQ2Z7wN0lpX
t0Ym2jKIfLUJjlv+a3AQGlmqFqJUlK/ACNS2gJBGUcIRo0Vjf8n1r5Rq0LlVX4pn7Mgym7tQo+t0
CkRYpERhbI6FIbPNLNyOfn6AvnM/N5y4SKu5ASQc1k1Go+OxYeumWEKOiiZVIgFqbQT9XWaaItDE
PXDEdXOdTHTenDLXwVI7GbwdHvB9Q4NNDTti0zMyBeMuYf6cGSMzKJhv5y42ZpzUCEBIkT1g9YQY
fzdmn8NbiwB5YSF20wkmW9Aja8UsmZsPbt2PsC6Qe3vmYfBk2ZVYVoYlXi40ZwABeKPfEXrKuxYL
93MZvZ1X4eXv4xLoQT7Hkcrj7e0QR/XSCiQziSqRsMXIMEHWE92kCLDMhV7V1Yf5I8St/KRULOwP
Lbt4eRaUmMGzM5vr/UByP5x08Hz9BPoXJNkEUYRKfg/WnhvNf1LeX24GBF/WZ55fDHhb/RIv+DlU
qIh/YMCx5Yhi1I+Ga30b83fpOmHs5etR9NsKd3bkfa6uizRdZofqzbuPfRbn8cIU4/ev8IQItTrB
p+sXXiLtv60NfM6m/F/7IsGOKblMsIX+/hZ1bVa1vT6SyOzQjJ6XHxr7d+p2rCWXVgPeHVfVExBu
XykcNeSheXBIP7pdP32ynNhA9ogIbNQCeoI5wXI8JmKh5R1rY7oyKjkH0bY8Qrzvrch6U463/M9+
oOGACJUmvup/6mc6nqGuqRqum42vpPh9TH8bRE73M+wl9cDMdiIPTF1OewFtvSb3iwui96RiWd08
NRt6tPWsLhN6CPlzwWm8J+6y/oCCMj+rNXp6Vmilad2lLpJQ6GPiU65faCiciOYCcTAtarZgBOdh
qHsjepswjdExLPRntpJ/9RFRFvt5oAvtzKDBg0HCzx/bBVS7UD87Yzt9cTZ9zDMPIA+UV0/TqbFL
Vr8OtwbEdAie0tfe4Ry6Z/7i4ISZTwuSZHmeLlZwZUkitxogRPDH0xoxURDcgzP9Thh4lhliN++G
zncAkNDpTu1sQPFkIVaVKwsBvGIgzh0rrSRUWufJgdkRikWM2UTpLNa69fPfINxbhCTQIk1kJYa7
97lqMNIiMquLb/HnFtIVTuQbbEBtRuflWM3CKNsX/X01PubDH6rEQgvcX2UI1fmyP8oBFd0WWg8r
xwR98sE8Xsuh9u/RCWttwbN9lBKxItK7t4YSj635IzBhZNII1FlNmTeUU+kyXump7aGSjtiCy+og
yNp5Pl9RCFuYQkrcZ5eUCy70jQQ1zGaZ0Q5u2T94uYh0r77hyWid5M40s+H9dJerEoec/J1GzPBW
ikl+k1cQ0SQWqoRzbsgtlXveoCE/hewc+w1yIUY3NstVv76HU9PPdxL2ifdQfbCBol6/r58TwSoN
ttaH1B4wlni9DeAyubDE8peqdKFbtcVAtZ8d+ZCFOfCf+xbKqKJ1BW9s19IWGBFYjF415o6coQMh
5BHtA6kJGQkkEFlaMJYZbflYUBMOmJ6hL2UtSWxvzQOUmCCTfoBvl72gGc23EQZb+HdK3Gmq2PEt
ispmX4DQPCGPH51n9iFiFK1C3CZH+KWUCR1LJ5mAcY9Qb/eyzF2S6EiAI/tszuhrEsqpqnxQtTjA
D+yBPxnagZXaT+3jK0LRfB4YKMeT+gc/n86INkcZ9nE3a5X1vwbcn0GE6X4hu72BC0afTrZu42Cc
iaJCX3skQeMPQvyoMAttYD79SYfyKmWl77C7OJX3BRnRr/z7oRgQ9urgw6T350PGSka97hK+34RD
OOD81l7pMYl2jiQoZvvs9zb/9xeDmdrim4HuWX74rRCusd4PjH3jQrxZ9m7Yos+WqqRRwgnY2Jpw
u9ueposfInU3llFM5AvHVkFQtmvfqAHY4fz84VyYzAn/6vjN8oQ00qWEEtV+cqrlGj+NK7tWb2Uu
Zus9/bhZQ759RmBEf6Lz0xbCltV4HVzU51Dnv+G9ROPocOABFEfJ+S5M2sP6ri9dDjdaUBsp4FJw
8IQdwWqaaSzYWsNps0m9/R+SzmFhgITGBYTLqVsWa6Ich8ntNB6EbBJQfeS8T6XtfUz3IVfWhBZQ
m/Lmor5emxiIhLatva/0W9WkBYBmd0QRGWYtfWG95Oxh9Iel57QQb/90GXJaS9CbEW0NBCD7slgK
4j7JV37CBsOjqhD3Lj9dBrs+QhVpsCiX9ljkKyDoTbpwHrXnVYrMnibhB9qOvc+FqrQeNw9D4SLI
I+Acbvf9ckPSkY88R8UyAejOEuHMuUxP42DqOvv57TGFV2FCROr+vpIlO1KI6msDMsCQknkG7/Nf
YwD+gwiwBR9C3lLjjtBeTmnx6MWhYIxf2FkO6ppDA3F6TTPrk0FaKLDAU5oSbky9VhCl5xSlxzV3
Txhq5Zf0PdC3scDChWGvw13DeI0nyyN0ayEHqxrm2aoPOmOsMfbRDGm61AZcIKapiipCtSBjJc0O
RN97ZsbfaeNikWRR/SOYM21YyxiX+tXYOLoOHmqza8FltRXrizYS2sz02+7aiWDe8BJ/ZLB6q6ZG
csSr/U3mJFarLknLTims8521akAXsTFaYv+jqsIpdgnsxMycqco1hevEHdZnarSkQQY33OyZ9BT9
AwzYDsv4AotAkIKQjWYWkQR1R+XyIaE68U6ZLsgG/gYvUCo5e//wMdPnnX2uu7qoWx4Kb0q/Hj/k
Hx9hqM31QsqqZfXaC+SN0KoJETWOvzLLkrtA2YpLgKdCjvWZFn043Ul7ImCJNChrPIV8d1vOJm7z
sDYLk3inOGnSDzuiFjGe6zDmrwMEzgdIQ0pOTVqZmPkB2O2fdD2PDgL5bdh3wutzNoyZgb7ubJxh
YEDGcHx6ZMzppLrZQgrR3xTO3pD3hKdpvEyzH5CQkz2yZqAzsOP9fYxIiEIEUFYiezs0X3V30p/+
zrC3Aj161WJQ0iJ76WBipunTbPiv70h64pjpKPZN8Qh9ilwkAmaV9IAAzelic/w91rFz3RrEBIsQ
8x8/9xfZuPwgPbwGoJNtutJHp9sWRo49+ExSpCt/CYpDXCahUmf3tmtFExzMn8646fzufuXMSU64
vvGfaohh3a5HExZ97Ahr7GEAjtaTTvoPRa5F9QpfV5floQiReEScSRmaKmYxfw2jbzAtWwf2XcPC
Q6FPDOdz66i+ksOlhw4KouH5X7ZZaiPDOt0y5WFKacm5Robt7jgtLO+fx/WqqdrbBsV0d3vsc8bZ
XYHeQtEWC4UlcrbntP44HigMcpe1p3KeeW26EZ6vJ/gsvnpWvow0OE3KHx5sCAMeZDxFhlgKCjNU
lLnzGtwVwGyNv21zzzLpgixEEx1+g54ffCtLZxtRRnVZsO/3CzaQuRE/uEZN6kkveJ6OrDEzukCz
xUivr5xMlJvE4rO6EIT9HkLviVpkfg3rGu/AI3+6A3LuKILTMDgLkGP8+kbB6YsSn/XKVFoSAFq7
I18OD3HXB8DAFQEbbt2SU8DY44tRvdoDwefxgL/JEFn4dd9rNREGfjGoV2GT6/G5wM8CNqKFgL+0
OQvj6xiW6g0/KaHe4AjOPQsaWhYcgaIVxz836KTGAuhHPBD7bqRJuJET/n5wuPwomIC42s38H80a
u+r+Vikd6tCsAgjpoltkS689IDZ3GFXq/RI7p36VkSO36N1fbDE0OK4mq4uCsDwLsC8axvjuyMsh
xlKm8LZoKJCCPl3CdAV4T/ZHtQS8zlfGH7DtGXvJ8kSup25UQ5fvRgUf+oOtYP2lqBiVskpcvBLk
9EoooJt0GUmVKJfNH8+wlHBXdZo4ngDP981DOYBLS62Xk3oeeDiWNRBTXruDrkB85bB1hFcXGPjc
JM17Du3IK+w+vHkVcoHqqnBQ0eo51EiZRrONSU6DBLfQNRu+uuMPhnfmftTLkCgTHHWx1MJbb8/R
2kCNDsGtJiajoTAhJn/9EYcuaKCUuSziaq6M395PEXREUNrBIFoL2IpuirazGe/PHbBzGng3WN64
cVDh0dLm7+ESZpwGHag95VIDOiOVrGgste0POm/BVKAvW4NghhfvZ7XGZn7zYe6yYbBX1HXbDZL+
SEc4puS28KrMRVcmwS/I9VuTzjRcNqgqi7AKKmc0qH79MdT6utwdk5pjVnVo/LoTbPmX4bXqA6Jx
UHhim3JJCNQDcPSspBQBKLggkv5+J0SzQ8LAk/DnccoVGvcTpLfuTcK76klW0E2VjHwvgV3F1yig
XcrPzVFrnrXRD/VrFajy2OgiV5lpYXfY6nQQGk+ailBoPlkqXI7qjV5X74OLKj6kDLwbCidECLbV
wqr2rBtkE7D8E8SMICJHhDmpsbWoJbsOFoNnuKWxgykXdc2nWYzJSsSuoOPmDHV+MXPqHmDD/xS8
Fm8pXIs3oZAcCmGxWvd9d2tDyLqSoIxQ9ZCWgVFOV3rAhIftSZQgJPoQKcQvJleb1kuKcr7tYOub
CCbI+nWyoY90jEE4W2wEklu6kSu2D+E2ZhCqae7CiOCNMBloJfGi3FnwEj3Q9Y9yJdKcthcDvBnF
oXrnsLfjb5xCPLB0NxmLlYHLx8w4YM4lI9LbCO3ubzb78T0SMH5+jPIfVUYBsXVIgPVymy43PAH/
3UTiZUZUDvXBHxk+U7rLJjTDACYDJZac1lWRv9PDAlj+/ANslfP73292zqP4moWlM/6FOQhFqlTG
wRSJTOwFDT+WJAsyhrpWpBF5K/1BwkKR0C3qcr4kXeG7K2/4zQSRfHIKAoxIu3Ps5uZHrDMsoDAE
I3C60obcDSZYr/epV+MR6csH+dyASS30Qi4DuhfVrUeOhx28DI0mJHYHhsHccKb4uKgJ85eRuqkb
xnCvlqHDTU0+/5u0LHxwBncJIM4BUSrXroZW6PzHbeQhPAPkfVrXFy4qBFiyV2sreCyLAHiEGmml
DM6hBza9ystV49pLFCjTnl+Jw+gqr4QssGE1U7fs94Ppg/r80YRyU5lRO7wqhM7AXdZO3vjH4nSB
LxjephvqTyr0dAvgHwweYkivxxIdZqjwTd8gs76B8XewrggOYijqZGgZhY19sY+tiXdybyzjnCyJ
pDGAocGMU9BgBMiy8pnTpZb1y5fTDXPhHd739Yfo+CZxUjNhWugfk8Q+nyN6ELY7IGHMuZXd3XZT
1ovtaCMYdMCpn2+G3QozDQelIi7qqAM1n0JXpNXc08WWZwSiP7OsPrLakDBlijZKmzVa2n6uFr0R
0wFmZDWq++y6cjeZPeiQMxxUov3Khv7Z1Edz4p7mWo2f3hqyZvuINtX8XKhU2OT2vjun8gfd1WAr
N6HUJD1WQmv1MreK9kZw1cPVaDlBy3uCm8JCSX98Ufwbq7KXqn153WK7EK+Lo43C/iWYTUoiFBx7
CzrLK82m2PazYE2f4pDGoFMcjEQjwqrTOCHY7G82OSJmPXJzVoDvDVuYTVMbe1+JQXsfKPBf0KGM
HNIefO6psOnf89TrI3lcI6+JHNcQI6z1TEDQXNhUrcTSUdTrLpka8OL4htb8wxHCMmdktVNKMSKx
79hnja/W8zYG+GKmXRDPv1MOGbUS1gRrsI2aL6AXKq3yjKcLyGN4PeLDbMBf9blgmMqo8moZRI/0
71xEHhwOPllNrdxt5LDrcOionU7CMMI+/ZBnP2FGtZd1mvk0xB04BUc1yfzbr73z3gqEiwpXdZhe
ncaDJvRZ2RaAiI4thvGMkTbdzttxnzZgD1gRJguwxWinCsZ4RBd9LdDz93GBTCcPZ+x1O9Yu+4gf
OCiZaF27eMvaHDtbnLesxxR9xfeTJdWpYUdgr/QT7U+9gztesXVZXmK7+9H9DbHparGlki4miDgX
j/0as16QXTD7JpwX78HekK5KT34LjzT2YNX/uCwpq39kYe/CGKtA67zcae27QCBX3w6FInfRqYcV
TmmZvvSah8gZOBTN55KUrEVyIriNHxBIGx+1e89ogHmhMNsx4nfHU9S1GaC5QgviVPUTd12FY1Y4
6bJvdw3OCLljYR1bp8yX30D0P7S1VWFaSa1KKlFPwD3m2OL4OLVvyN26fp082O1LzIFJXyZ/rYAv
Cj0OqFw5wIQ3oSCy4djeK/Zxq5vb8oyZAb8PnbErvfRm0XsvQQw2yxAEuaXOHJRglhWpMVOiU66m
vG7H1T9lCeYFc1sV5XdzMUzt34S0f0KIbq8cW+01iMjvCPS9UCJeg+5tP5TbKBfLHg+rKnwixeRe
zGUDCOBG+SFrKPLSEa43xqe8p6b2E0OmMavVH1UvKkuzCFJfyfx5RWInX52G6RlyYHAuFdHFqnGF
QXpALLn63zw74+HSi1KIaakN79cVxr8vJiJpksOYC83QzeBWd6SG1uWGqVuTq3We56b2M8PYIWyf
yvBN4gbqQRhxkLtJmk2ssMeiC08Iy2C3Xjq/G70jbqMlwitpTtYoAXazcWdr7WbiPBoDtds+Nc6s
JTgBcJBBobN/3pCVA9G6wOycJOs8v+2gVnIPkD2UddoKsotHejZKm43w/v+qJHi2GfnOoPouDkHB
+C13/Z1jKI4OwiNfKd1w5SByy3WO6wMRcSg8aIVXTu4Ww3RC51IQFhlDpSO2p77yYc667WU52imf
BDbOohhD4icVcBkzltFZp4K9t5MLnbu5Rm6r+HOZMNeTvcMFsV4NrhIFdiOXPwQUKIxHP6xB8IAg
Lm/Ed/dK5UhknNyMOG6HcsbTniRKGNlshNWJ8I9xzU6O7CLVG5E4MeGYqyS52qaRhJKLj7CNCwVf
a/Ajusug+hHdceFP3O0Pkurjxgo5J0AZn62GKiz00UUhcrR/8mvXfO1yTYqUYy78nVlVMEStskfi
qEWe6KAjNVx4X+MfikS6TPPlMo83EtZwI35WBtiy1FnLA/CDu1Rgn0IHk/j6vowvXz9n0AE0NT21
90KNfmuw/0zxA+m1c0uIQh6cBcbWCTZM3uw4S6BzErdnypDCxaVGMrGRZaXvqDQlVNgatasm1CpV
9jIgSnZ8k2K/WAhxC1mgKOu0mL2rDV6/f6stE69gSSNM2M483+3LdvxgmA+VWqfI68pBY7cjxMeN
87rgLoAMGjBK6LTql6fFpv/MzZfTDal/C6rLHQU1HKIMjjpltUgF1v+iIclU4VBDge5hRO9kZjeJ
0/nVYpZhttTuWbzswURQJHppO6+N5vWaxTnhPg/Hm+pdJj9+tIZh1UOftSbRcn8oqyDFJm2VZAHh
Z44yH2VBSjOAEj2A9/HkP9hsCvWNuTkHQv4pXBWus697QC+Fx4E2NVed0GNHJ5HXqC8/LRqQJiLB
HXnFbUuvP8ma113tU5lAVOgVGe50rI8gVSQfD9AYWTPJxblpS/zm8xG0JlUW36Ta6SvRlANx4Dki
4zkvisUHaf7AadPYO4CrJBM/l7tOrjF2EVPS2Cgzh7Lu6DgTD6d8g7bObx7tc/mZwoRO/WpVxOw/
GGCwGeulWstY+b0iMXHxEwNvBHjLGlJTB2QL/wQylbBAhiRGcs9ASA3LIhg3GmCsdA6aCAcvfZol
RZ2WX8DPEmeFg5F/w9NEPnkTYd8/tRrkUVbONrH0valtwdUEBZ71GuBTdhEAybJJc+cuxmxy/iiw
DFqPh9i5MgcwEYNeMBtQhRQMeRSu7y+3efKx0V3wArbXLFHU7xbfg1xYPKt//Me8ZHDgFlgjCwvP
HH39tj8nnapr6ZnLZZ52roHE8EqZMpalfk/S0tYwQjdJrnpgZgmxB4GM/JQiftbRcnW1vuMwx5Hc
1xECavKZl368KWMNpHJK0GvDiQyhZMPMJBlKks2Ua4YrMbVncrcJT3jxSWjO4R5E9aJQ5HybYQ+z
Yud34JZNK1kbxIFYNEQeQ2twQ5f1aNHGCDGunIZNtNVK2+j7e8w/TG/ISHUgPSX0UM2sVJfj4hoE
RvP9XPXOWKA11LX2jv0Qn8UfiSEe0RGxAykgqIXCsCs4TIwxJ29DK6zqNBOx3+Q6HPz0TDGQDpmr
qPgfqHlsjAuh5npmZw3aHxNbeXjOIDiLrnQ6Aiz2xPZdQDvhwcDSBRhHZnRf0/OvpAgzgo+A+T6p
ZXa6f3dyWgJ0a+lpiRlB6no4TdnIUkK1k9Z2Xlh4LetdR978aRLnTJ854PfRAHMxHrW60wwVjLa8
xcUCL33TULJCuU37SUCPFiVkmeVC2E4rQqNk3T2bNwPoQPJ1ZkRYj0mhNMWBYI+poKq3Fu2NbGEn
sWC0aaRTLNnXJ5R23Buakzlyf/xa5Xeky0riaE3bVRAC31jpCV76LZfF1b4UY0eDhG/Dw3SPlCSj
bPzd/LwT9LiGnoHuG7j/2DCWSJDgt2NbcMOYYtS/irx2Yi32pj9l4VFzdoLCwf7QZE3FxHEXH8xs
4Ehf/SXZfT8OvK95ib0QWqAbwhPvym96L7hs9uif48ulgTtnDWz0KWaHVFHYTPZWcXQtG+TynVQr
/JoIOxUrnCmKEmnXKZgvDRm+06o5L4sq4NDlJ0quF9/iX5kn5Glrc3a3j/pcVs0u5ZeUfDEk6VCb
iGeZSJIwd68wMoHMOaze4dvkal/YwsULOGkkGiiWImmM0fcItnhRC0QPDaFEaTXeoIDMm4T2CIZ7
JIbNZM4TTvN8CLDTfWNZ6HDq3/Y/tqCpFDiwCGzwdneZUmpCtQMrwnpvFpcop6WVgYwJpNAAmhKU
9NG/84HGjca5MdsdsEiapF1W3cXClg9pZLwuo9404nPiUxQm+vXukATm6LGTOcAHGabZtL73T17D
qYkl2Pk4oYwTd3tPwB3s+0MXbLiLZDKPveOZEKpoSRy/+TynzX49RX6ORRbzMmCm65XdIXl4+d/r
QGR0tXhlCPwY7f1H1tdK5aTvT3HWTRU4w5Bhud1H6xOhLCq8vOromSAGMj4pX/B5c+Tk9z+cvf5A
IWkWiYI880msTNER8jEVPI7KKuukUfkqgyV8NF5Wz4cjV65wwYFoYTBirJSy8mZ8wcbNTW9W6iNG
1g1vzIIKsxJnIpylncvpoeyTIW6/Obtt34fmfzb6XvoY05LEKL1IEIszNSpUyJ/6q86dfsEHn6D2
6ZkiWp+C2Z2Xd5ORhYXPDQvu6/l1kYSjfrRp1wqs8Q6Lt6AjDEyNRFsVlJRcNlZoaKUjHMdjcW60
DHA6jIj5LemcBJ+bj97EM/F+QmVdBHzdV1PXeTz7TF5nWjx7vVZTxKFl5hjE4NL2RBnW2G0/jWS8
fadaZMcCxvluNR8WXXNe/e3inBzm5+oXwYn93YgmwpFKUOHQ3D49CHVRzLuYhKTwNBH/CfbF6jHw
IisVAFbCyBVU2L46GUw8H6ihWFihWQLRYS6lRfjG2aVq81s93VAeuJMjEgQ8ehdvHXTn+1mxN2QC
Nau00QGA12KKcg4hmHk6tPzIk3QLHUntGjXIpriWPGW5NycDSNrGOx38nwWSHC1RuzL7NcGu8OBC
rMcT8Itjowf7DMF+ZROMk7AAkrqZh+3ZqjQPFNL34AKW6AdTZvmW4ViLnbLSWx6zX7NPPRpI9fls
OrmxzPNbOKllLls0/mXAxLJvhLxXrq06g2i5O19AmJ4RDnN24fZe3BYyKLuXOAqB1OnwKkFp6ovS
mrVuv1Vn65wizgepbggNjYxTGdtEZfByjUrl909WPkv3obwQtk1BXrvBqCjUrNdU5pBLIpVP1hxP
JUv/gB+SG8/Ov4uGH11Sw56JxkvyMaSS9upWnNm4d04fTVaJTake9ZjLHyPYh+HmESNFz9Uqcd+S
Mr1yOOxyAdg6R5j0+u5KAqIyVTBrfR2c/H/N0X7/a0CdlzDyD/eG1kFo3HtgyHvFt4VfG3BedYF0
/PwuoQOY+6YWSQSFXUXftJwhyGRue/r+iz6qZmVwuQzFIVBt4Vqaw5zKlOL1+j8+4HquxBYJscyW
NKoYwko1TXzhZAahDT1U+Cvg5ciTLUiB+G3UTGXp15U6DZ8sc06IRZhnYm5Ap5CsY7tSb+gv1TY0
cWe+pFlF0RGeIMlcxA1pRiooyuKPbyefd2+SrkS+riNXAj/xRQdDa5ThBV2v5pCaWRtGUGOAiWLb
QZD9d2qBRwYlR4DDxTtV1HYaQH0q/C53d4pNT0ecpQ5uoCAiW1uVF+pt46ikNYf2zb5OD3pVFGjl
sShbL7Z8+OAoBp9/gew0mS3V0YRx73H10musZEYPYoOHeI+4OhCZLcyKYpp2N6mTzS5McMjsByui
9X8zqtKvqwczflvDTL1/Upewt+RWBzUA3Jn4jnUakrRuWnOi02aqx0MC3eoZumirfpRh3PKjF0Sc
/JePW4a7Fzk+BhLRFrYuy0F6YvgyFlW+wuSQJdz6DCtiQtavZH8b2MFSBvGY25QwSu78lD3Pu8Ja
/CLdilN0UaSr2VfiCDUG1pMkjy7IdvU4vpvtBHQIlHdCJnY9J6PGw3YMTNqnuGV0OM6id0Ta6oWm
DRslJSZ+U3hwJdR4iVz1/9FD1XE+qD3zeLLEbWrMfW0vU+TO/Eu87Us2yeo9ae/T6qFCQruF3t04
Wh/PPsRMIDW4WD0LfxCc7Jlt7idFkNYOozaGICi+4Xx1ZOul3Ot7KCoHye3kBrbIV4jG0yInNeYl
y6fPejoLrsxKil4TujYUtxqtmNY5H3Clrkrbqc5ogLoVc9FSW+eV2tq6Zgf1gJdtK/RANZdwbQX4
ie8Xw1/UKYkZYa/nIqEWT90cD5etFLPmOO2rQqO30rL7gWBjhIpZi/SZRk7r5UupDmwCf7KCnKqQ
3sf5gffYho64OjyW8c9OmUMVyGXDY5Zwlt+rDTIbRssIrh2v7HidP427lROTWR6OAvjWAy47qb2J
PPs+8/6U989sAAXI1gdHRHrvG25uVXjF+oOZNs3UmkD6rNNFJ0CBA1dv0kUIjAhKKuVfe/T0y/P1
/vmwtx3kVi5myJAGBseD24u1X7THJ3HqRHugiB0Kf8md6+EuPpaqDNV/dvwAKvma1rNf48ViXB1P
kEExTtYpgdZ2pbBJiqdz6zXHV1KjjW8PWKLGvEIEa0S1knrEXcFY2Jl6O0UckpLarksTMn0SXyy8
uM7KYEJuHS5aEb1C9qnhGOR9+/g+XNeMLQ/1j1qYXg2eOJnTUY0mS4wjextB5doQijeHLoiXbLPu
XJuFgJqkv3x9lUlACxO8DqRyzEh2sIYyxBMtfqAUAhA2Cvn7ieCARnb4XD1LDQpjAbE1YYQsT0sC
XCVhElWlQgeN6jiLi02mtHrM6z4dVHufzLJ4XC85bPsnSKLVr+5aTGgtHxBglrjKNSRu7X8CG+sM
7c9guZVhp9DTJ/6jfI4NJoSy4siHuqRSlKmC8HGAh9yIo8yRnt4kZw9FWOXTUgAJKDwRVUr5f3Br
HF2ikYW1mwpSWYcCbR/HFsZxWAQjwjQmN3FVA9yELEIiHJEX92s33zxGMmUJq54YWC9rrBBEX1ii
4HcG3FXkNdiyyMr2BWu05EugK41gwlqdYL+5g09YKOH7jQwIKhuqDU9ax49XMBiYXeuRwj+uR8vi
HN/+1xvfFmMGIlKz3x0tRIWLzAH5mU1sL8MU4IsEZ3enBmrpcb5p38WMT5HkgJ+hgDToPWf4RACt
sOQXN/PGBzQY5TnqfZy4AsUOE/gQ+BwQJqCYjU32G4QdyujhZ3ykBmHayIMOxsvW3GSpFgHvOF/Y
OLVqvqG5SpJtu57rmrsAFrVf59pLWimOy2vCb9UruxCwOsuqrz7qeqhXAE4P1XGGispI23J+tgGO
m13SZv4kbk0tuBJsEhimQNOGFWNeINlXiaCD8Ag4VdxZzcGv7SRrXJdnl+7GF9yNoFEdjEkAW2nS
D01GEpSdnrxbn+P0yuiJg4JSxy3l8zTZs4d9H5bpOtOd0NNdt4kZaos4BW2DymsLzf6EpmyyJKE5
9yxIXehxqf/zhK/4hmSqKjsllGBSd5I0g/yPP9t5YGZktcGN39CrGVFM/AnIVouljGQ8fiA0b2th
cwjJEGhnabCocwk3vYg7i0EN8+JzjJD/3LhP2yg2Xoy2V0D0DeicMsagYpUG6NRVq8wfykGAbJpm
Y7oDHeDUUdprCMmBpwbQRu6apzthm4sGhJ1Ob9I+P//KTQaVHCzJUHo8IVrHqpnLMh0gn5AA17eo
DV2pDoPVkjjHHaxnbn8FNeJvI+T51pEsz1YcZUKFban8giSw3zGsldlNHDa+jWa8JUhE5WXSRFXz
21s/eBqb5Z096Jc7pO15kxbUI9kxKAg5+BkDyv40KIy6rEA7LVpJ5LEYa3eTc6gKzogIivJVIbBg
A1TTKVVBEhMnTPAa4Wlx73CqcEtzokw7VwGrPCV9JSkgWOk2Y9fNbJJKnQTgRZch0Na9wZMCLb4i
Mp+taCHq0ku6jjTllHzUbAIvDSm7j4R+h8/+2OLS1ZgHPLuY5GLMCt9EAK2p+cY3QvC9Qu3Hn157
Pknbes1k4Feb37viNh3LN3JoyY+fCezREnBZ7aEhb2RsehEW354/E4Vhp2t8QW+95XwzfbIlLaDi
QiVx7cFpYUfxWLiq6fjsJvHrcXkzOWeRjwjy79FlDeNm2yPfgnYd1odrlcdkYc2ntxKMkbyi3BYL
nOLFGtGmpZ4snNPM/j6oM6lV/1czyilaXN2aZN7EHJ0fsliurry8YATQhlucgTZgcC7k0mp2SXbZ
cSb1nnshFnna3zbzfaoznABxrb/VRLbt67HiNg/5rpW/QXXRTB76vbj7d8PPmQyxlCHLgUZg5e59
4gQlwMtPFkXGdWNN8msI1fdrXIxEms/mRBssjMwxG3Io2V3Vd3GeRKlDHsVTUgfisxMin4CbrXkt
tA3JfQMKGe+bnKrCMvQEDnB8mlHGcepZYJATN5Wfowt8t2k0AxOf8M8bLTDID62rd7GWVxAL3v+L
g4rZKDEC4/ubkf8rhRfCcwMciz3AprVBaIJTpk6XEP/fxmDTQDCTglln1xtgyDxi/org8aGT9snw
q1YUik1lI5pfX8JGP0KdyW54+W6MYKLV61SEx0RY+fFJGYiZB0xIrbf2hIQhTJRl83OU75xiwOFi
rqg1OamRvpupCtSzB6NZeryxxiGyUVNGcjS42fD6SLfQ8cH86SkVgjmJwwGRoWpkD5pKLCKhkbm8
JriRa+7HMbZ+P/VQJLh2QU1XJYYWXe3xSdVucmyvn4v6VbRAXM7bpLfHRL+Baxv6oJYthRKQt/iu
mdKldPqiwYv2dsY0GDmfj2XdN37n45ccjF3XRKY81XfR6Qzgf/uXVAhQ6bBCniSEsuZyCRT8LF41
thuO6vw2bNDcl3U5m8PKeHm+Bi2w5cJe91H4/ZJny4YLaOwUj/BkjyW7zepolp7dM5xP8POtkXT9
SB4NT3fidtXWpMuHHDdxZDaRTDjYQk/rpFKxy0z/phl1AKul4RotlJTtVXCJ3MRjJssfZiJdQOHk
LLx7zqLF843hJBq6IDKb+ABLkMyOR4koxI6xGQkX+dkNMs5raZHX/zv7bpFvIcQW+SN+xQCxOLa8
yK50HRLcdtS4sYiPIJi+kBM8XtaUEQovHQ14C9YNelfWNJ2DftuwMSsF+FnUlc9z9KSuA4HlPKwl
NjgrewxIjQT8NaQJsDJoRx73FjMaa9X3mQfpe5Xd6kj9ldsEZEPLRPG5DjP0f/avF8xTi5bmNci1
ecJHe6PQWp+mhsRGCTme4ScZZ+bnYBgzv8LSOozujQOEgMoWE/50VpzGwSG29e2ydE0oeAG+yZ9w
6vJwEdlD7/MaL0PYZWnft+rXxgnlkoMz8CwFpN1QJzbS2gzuHKULQ6zFNPsAn7girjox7exegg+0
Me3S70SYkyXZqdLJL5ADCvw5bIX6Kid92BhDeOF5A/gKnCBEE8LMiQ1m8Rj8dmKMvSRQzH3loQDV
Un+Rj/Auq0ry6kWpZ0oscyUs+Ac+i6TiUX48zUE2Abm1S9AEvhxEuKEBYYMEMVX4rEs/drnFZ4Xd
z7KHSTV0aUDGvlR1lSv2z27NzhIiKAHY3nmAQ7o4zP9otkv+9ciFD5swW/6Q04EEL9XoGpSpl1Jp
B+CGRZg5nmodEZ3++lsgbFq+qKaHJnxgqul/wpDjEJh+FHMYgXQUfwDVRsl24xitSITLf0O7qGXs
i6eUlJ1/jhIKUI5NjHPnHnVeIQH6123j6denI/kHuGAtrOj+CFVEDmFPytTSkU4xVUVOJ5BoFlaz
LitvBB0z0/FWIAuhyobRlX8GFhP5jdKcI60tZ4ko23Ey9i5lLQvI4hgdRCEzREHq6UruIlk2O67l
WiAPfoATGdOS+XYex1WaLyMbFSzZf14fU8iwG39uhZXkBND13vB4qtGH7vmqwU+OUziWvEqKXVen
cTgMXDJlA3XZzydwoqoAqedc9ynyDhQDd2cVJOj0C1GKG/eFQQZOn96o8sq7b1mlVnSxAPLE0x7v
2bbbYZngsPV14AdVCQG+d7K+YZfmauLlGhQ/vSI0iPt8OvITeEpG8fL3enu1uP6Rjw62TOLQIY6J
du+WY1vDvSJxqBBnlHT1cDGZQfSyzF9mgVJb5OXNEf+wy6ezderQHBwtjq6KwzCDVBcylwA8FWyn
BMiuC2zc77ZUhyohVECczv0HxNqRiJ/t2GcD7Mu2R6zzys8uXzNUnTxywFriNH+dOTNx+7T2zyMg
rlRu3kHSH3drBIEcxXQLio/fNO1ltbiuS+RFK2W+D8XRn9d2z0A1cqviOODY63G71UoWckOIZqN4
6/ZelxhWYQNC5mKFKvkfQuK9jJdk33X1h9KoDMacBN6ZuzmcLO8zshdQ/mvStEsPu/j2XyYfLLsb
z2FZtIwEUVCX4I7p4tXTR3oWIfATwJkZE8CpMJjnSQsHuY6mJ8YdE8B21xdY+B/RCuGkKE182txv
n0iF0xXifLdRBTdqgpzWeJMPnXa9zkM7m2HwFCEVlQLmz79CubH3JMFaYs9vKZpCx8DKCMnVDO/I
musy4AU9PZIH+oudFjyB6ftJE4hgEt9Kvzc4QK8CwFbB4GAhgbw6bdhN4zWmzNmXxVjTF0sj6Uy7
AJG/4Sb/EaqSUF/3TNY3JwM6b1Pj6sRCj7XF/ULHshYcgkBriy+xu+WrF/2rzeKTP2+EAg7hP7J7
xVuXNPfBuMWGVM5jWTk8fkgTlTT1opTRIssxUwsEfvap2AgTPo9HMpif6CrBqa1IMuMSAXhRBg3K
DSFTW9oy+3jQfRlr9hvoKQRZ+o6UbBoX4mVsvX8UfoDpgxIWymaE3pYA5E8RJqT1phJcN8RVIsav
KwFo4stu/jBHcC1+admn9jJq3qVfuodxpXrOaGiVb8rjzXNxd8LJqjEDd5OeO7aEJqR9MyEe77eh
f+9xArcIUjSCJ2YOXum5szuKEcAo/nxM3F4Z/ozn344N/+LGXNMgg8tXs+cLuChb4q3etT4W2RAn
c+zu1hy3B418A2uVuAdcMBUMd467w4WaWED8XxbtHVn9NRIWcUPonpL/S6q/UNrl4Txkk/vR3H3j
KwNy+71mEko4oGvE55eDcjWn6q+h4mq/iWJFDhKsqfTtCMwql1CvoFIpbjTaeEu5l/LiJKwcs3Eh
eEeuaCZENrGUE02YRyk1zYXYLlIzHMZFMgybPXT3n5D2nHsavEmQq+otEHJT5s4IqM+WemQpETW/
u5vT5D+un4jDnM8j1MZb+nb+Uwdc2+IH17qWFhlsX00gK9lJ+4mJ2QlWjcuecpNKDwlHcT+mePyq
h+7RDy+LVw99T+XciJR9yoItSFo2vX8adhSovOY2w9cZyIaq7kwR9QjlmcmpO5o6u0mduMXv658b
RGs38BuXKLEdcVLhdGaXfoXzJPC0oz/jnCS/beg20L6+xxBSVoD/M/ICc09XmlCXD7WRlr4LaKPJ
KOQDAWvqamajbshiunTdnu6BMq925lrDYeqwp+PPvew388bDavUATVtC9fqcmAU1TKQ/a5lvZAcg
vgvDXzo4m/jwWY4TYU/0fV0YqFkN2dy6ef2cxWMJ2n8xuEYwEjlc8w24vXtuWQZFhAhPWbkFrphY
DYITmRxAAiQGfpvo+WUJe6wpIJ7N2ChDEZmb5hfClRKNj+1N+sY5bAB81JN1F7btGjIY/8SZdYee
txDjibkTuowCAHrJwTc0w12PnCxZUpmv17u9OEmv8zwicSJVdkpaDzmzfieeZqzhgsyJc2/7jp0C
WsoNAvWC80O3+wg9VjVFx9/PTBwGTLqjecd70ndltbiG275kzaNL9ZASWQM8o4MojHIM5W37oUtz
IBHjsCHm24Bn9OUKXu9N/qVUJXdhKZkX6JOvjuQfBWMBp7s495Iua1Y6QaHjD8Y6Ypj4j7rkTkgo
RQABEUa3ZytP4n0dxPelzpQQzfniedJDwp39vbXoq1KPExbJeefOr0SQBaq5p8E1Sc1LWYtTSY8R
kfQxrXMKsHkBdkBG0PDdIZQbgds5PH7OFKLsqsnmN+BiGjxKxGfnsuBFMNemlF91mtFL2loQrs3f
99CDWSdrVGDSgbj917GfL0+qslWkU0x1fQOduJGhZm0p300OvN120xPt/shS2ISI9Em+ckLxyz6O
dRJa4kULv9OA1aj5+H2nHq0oh5Gs3n2JTVrtvwUlVt+tQ2XZ8Pz/LJ1+M7rgB38moFjdIhCubFm+
9UIDNZFq8FaD3/SW5mkKq3w4QsM09L9ggxtYIdB3khmD3ZZSXRZ1HId7MOIllHOEl1lvJBcTVdxk
2Tzg1IMdSjz5V+2s/i2RTNcAWY1fuqo66Fser4Z0WnXNHbu6LiOCMJG5iyDskm9YBusAOHbn9391
ZfPljwu+vgmhE+IoupciIRx4dThXZWvpXIPuHRrcuVEODalIlVnt9sFT/baFOLbWZ8HJaHiQmnzl
kbKXyiIQUSpDs3KgCRMhjOuH/V8JBVBmlkvRBYJCVqa0mJleLE2y1wYADuGd8XYSWBSbiBBp3Ca7
zhOV2G8OJdhgGcVFPEPSYgKSZ6/I7yTs6iqIfqugwGIhlZp3EoJMYV7pIHtmKXmQnFjZsd72HkX0
6SMnr75MIINphxC+nfk75OM+IwxAGhquyZnC28F1gF8tMDrQUIq+fUoe4OhoEvB8uzyZnhcs7/b1
c/nwYHzzg5gNht3ZTWNuCFJ23MvR3bJ+d7EF9zISFpj7JmrP8UfVnGThieLSF935rv6Zzn3k/ssg
AfSLcor7EkDV4rqqyiVR+LLxJAzFREyLV9+nY3aNEmu07SUCcFxMgZCSgAtr641kjJkH6cUNZIvo
X0u5VjNVETdp58pM2taPzraGZ9jSx5NpYPmUxiexzHYJEkxzQEUwTV78oP4JyP7GTVm3yL/kScEv
dvdCtaZIIdxFHFRpkqQD1pCy16qt736DCrFbGnjaWORzV37ah5bGpP8VDqtCqCj7mL5ou53xHUtQ
YZ3xG90Q11CSn00lQWBUBEoFRgjaR9NzybPX9cUdAiXOnEKxDYk3h6f4MbVv/jaqWQfErgU1ecBU
WDv2/zLCjopk4FF4HVJFLMLqMxKxDqjPBWeDwhFVNtZMfoUqwad/eLF/eBGWb56OhZOnoBhzxLeZ
EtBzkuBKL3XWWxafW05yQohhnj71sCnOKggArI9q2nJ+1YHlWiOvg4FsW6Tds0HL15F26CDyxDhy
Bu2qHozWvm4hGWs1G+gCRBTWhiFkn16Bah3rvuLbDbZbW/maEpBvkrlJuiGSkM12ScT23XoKRY4U
OkUo78JX79xgu7q/hs+nhz4N9uT8QMa3iWR6MTD7g3ReVwb9pD/ECb2dAnxzCcTOlokw43FmLGJL
MgjzfQ/hu6E6C/hGantGHg+Fv/AiQs/ghAt9B7WQh5xcMsG0sLuwc7fm1UFBVpLnb9tERZe1t7Oi
Qjc0WBQGNb7ZbsjtqgM3+bRz73Et/ubjyyTmZD2nSALrL7vQXT6ffb6H7omkLBKakDLuo0tU2TEr
a1PIUYef8ROlUCHPiURIvi7bG2IbuJH7eaITDns7wr5pf/RiM6flB5Un+mEYwsMhMM/7YmD91iYI
7GysmW3xrbdda2qaHW3zxxldhTFvyc7a3TDPItgdK0bppqCFhg35sPR0qS8Zaf83d8fH0rrbXBP0
FJ+PK4RAI+OQd1I6NlPxJtubSbltXx/8JJNh0IJDfUKPh7klEGVlWwS9h5NHEElN/CRzz9qw9MTT
/9URFjYPKeWOlrWqAQLkGl7SgvdPkcNF014DEv8pWN1FGFnOK99GrRKzsIKzLzL0N/r/d5ACXGXo
xX+iW2BUP5BBfATLfMfO4h72I7jhUYo7I8HpNm/Qj4vOuVkNPf4pAws9I9ZdtAUseClUU98lljfZ
PjY77z31PbhtE8uoHQrwiRwdeB0HDohBDpIyEGqIUrJGMCUdqSqBXD9rnPmz7q22QoGTKBsE7KlI
cezJ9dxfptJp+ZA63zgmy+aAy59JI88H+MCBV2yQbTf2wUbMDRBs+s5IStLxrxCCv5ITCN7/sQ0J
DEpMsEmes+Zip7+g66TTrA5gaukyZeJqqG5UB8orxRfJHTmq0wxTu6lpBdTsVKKp49jahinBhyx7
FVMryBcJYZW9P1jGDJyt81yvzROCXKdMc5OvImYzZBxX4oFj//sfzrTT2TJafZwVZxwJhCfwhVl1
I8v1gf068nOJoSt9BLA6vb9NzBJ2aD8DCSCY6SP2yCPj8P0Hqib3vpKeqsIkXBBXfNAL1gfnp3im
Ai9reDTD6wOJqIoP0tELbi6X+mGfaSCnt6AAg6ow3CzgSc1oLCkksYHpHO9oivrfFGsdEKvhmnxM
4LSliLJcjHSWQ9ibIyu3Kn4dE8OAgkVd8K1cVi4qT+ff57Fu23ONg7FiUtV9kOx/u6k7i8ofzdXM
/Tciww5d+v//ZaB6Vqzjx4IbNaA/AAokhMmusmIk1zMFSd3dcVlwu7859+eemGhdLHrIyo3caVWs
2Km5ASy3TWGJE47bOyrjzKCq2sXtPVQh4WX0tIQjZqAtjCtMQrdLqMFcS4BGYFQb2a8TR3sNveYH
WRckDKTvc46DWWAG9lAXwwVD1VJotIXWINWEyAGKgAWkPlD31jc0NeZmZqjqBeQtraFJJFnRc1W6
vLpBqs7PvgESxTcaFIDVrL+roX6LT7vuUL9aLgM3KtC5ObT0JTDtkRXXTIZQ6tKGc93twxtTFPb5
WJ2DDwsVYBHQJI7+FX6jrFTNS4j5VqtoyZH3CjjgXgCnva4ZoOTyqoc1038tuAd1M1jiXZcUsAot
O/sbMK7AXMZTsQTm6kVjnolbmkMOhsErjux0G1Vzmk7st/+di4ffT+MDHT1ockS60B7NM2kjavig
HTi7kk0mmnr44VogUsCb19eKmSLnw4WgoWNRVq/jlaqvyGksZdbl0yzj6vGXWm4n0aPRjtoKjXv9
0/f1hoqv5oUcIZWO98KBCu5rKbLqYWJIG9yzT0BqVddCVBS0DduIXehbvEE+3OKsPpR9xyVG5x7v
Bk343+6Q7Vi8hahsa9t/MpmWCqbJoonlG+t7TtdGnJQSG/d3JFkz6KrV/harI+9j3rwdLI3QXsKm
ijCuXyYT/Od/+V/RdiqYextksEAPTlVBIKsBkUQdxC7CVfvEfpKx+GcCI2x1PGRfZgkcFlqEEbUk
Kn7C+zWv1Vp2fIM6LKPSb7JscWH6pmjuNhvw8ghxEjbaww9Zldsetr4Q+f2cfqRc91FUN9RHg3+z
8XjtL2d16ie5ViFWa9VwPeSf+syn6YsSX9X7pWX23rD2sLxd7F3RKAgikXaqeQ/c1hJm9Mxbr6kt
q8o+vZqvgL0cDuco297jXlZlxtrljhd9Q4Vcj3HGty15aDa9iiYum9jhAljGnbUvcSIMu8WcSLor
OdOkXuJRaJNi8D7jOEZmlnhNSrAcWGs6idp8T4T9z1yCl49gwqyb3Y8g7LdjYlhqTVeR92CAKHlu
A7Xos55x1bzl3c85VfTK6v1gtxXcy5CwxhmS9vx+yKtQAZgvrF73TROgeNo1oflN65gD1F4rG4HP
9vATJKJuDKftf7Zk4C+s8bUUBduUzD7nnemVyAHbcb6l/lKJNG3NhlBqTZpMkx5erGVJI08f3K2A
zVGwj1+P550wZdExciG7oZtuUnsKzT3hcWAV4bZsnffFNGHWCPSne7qYigP+gKeAa09k6GqRPfl0
b6ggdP6kf2MBa9Oo3msv2vBtzsF0va1fN00PyoGE7fJLf6dZBHDMgR8pZVafigqIPCpvbDQdrdD2
WxdsVJfZxApPg4dU4WcFgyYSEEruCnrQaIXIozjRXHM8QQA6ThW3v8UUvJWyTVHyFG+EgLeSjVUg
FsIVk9p+J+5VHrEEkFhhtKbtUnTID66QJl29VVlsReothTxJOxVSS/4hCe/ki26UD++XRd6E+Tdo
z0gbu4YizQltokC1HCpeAqrBbEhqXrwFL+HgTnUL3E4jOjxCqJDhP2jB4wS5jDVCeH6FyE5UykPx
1E6D2SwWcMfwT6iwgTZaCZaAyc3g8UrEa6Vm84byDQECpny6Jot83I6hjVJ6buagY8O4cRYdtqkl
ZtTPeDLoJHwX7E40N2tATAxOOB+Hy+sbrYevrQ3sTPbKq8ZEg944GiQS3T8xLb5LG5QO9NqPyRNi
V2Sj6Fwzu0VLlKQZHplN0O5JpXUntx1aQGMW/mlh2ywerTlU8VxX9Whigt6RQ64ktsovu5bn/QDW
b7kth6KhAcji2TnAuPBYGJJzCBt6lhJu21h1J/Vdg98XgpLfb3P0HGYCyITS5VbdiKn38Kx2WQ7z
1eTfMNxs1UZzzuP/f6kceaKOSQjp26K/iKfFIdGyHJYNQwW39a54JCzut6IoblgbzsV/yCvAL/Ln
gy95c2Zr6vgw5WzJbcJT84+vNL5F6MqaD5MOL3JE293xztBX+JxzxDzJIj1CIBDyQYL8zv175NO9
SdRT2CzzuxfUhZrToMSkoPYkvFPv/8QLurTpvuzdLZdbEGgIo50z8N8RJ2bpkQKhzH1K7JbVyYoY
O7n1qmEww86QnZWqWCJvJg2gmC/Gl2TWzh5846ahWAdz2twuWsmCuLeZbeZC4MDBv0v7w2JMgwGo
NfHmdRJ2P9EZgnHVm0jAKrBLRpsNR08QshnhYM4j3OBcn8M2E769stiYD92I5VN/qMsZPVoGc9OK
GgcA1uj7tZamUnT9vCZJcmIKcv4vyVDSneGWUSfIkjp7qFir4LL8C5XPZqYoqN5skjfdvvsAPlmJ
6IwS7emHk2zjldonW+U5VTeSQnHxecAYBJMlMwX2ZS+BWVgTpm/hgpKjGen9/mVm1voujwDS4CbS
iAN9tms9TB/+EdctW+mNwdtu6MtrkriOMbVAkobL0NFKHL86IORTdODVtSPgDJISt7nHcd12aP9u
866v0ukUVDhnJGrR9Ikk1RsnGT/gKAwjJvuFXJpMlEfLRWN2GdSWCNxK+u9ZHMsSbhS2rP1RbyFi
Te1OmjUZ2NkIaHo1qjOtisl5cKFboxRQELwAxRlIihzTv8UYKtuBKHhtFZOOkTTX89og06gYvyUL
6R7zEYF0F0ac5NTFJAtJoEETsMo/4qWo7o1WYxXu/iLe/x5bEciVB4XkBy+tehZ5Wlm7zcr6/pyg
FT+w1YETa43KBsmB20TcioomOxUhITxcyZvaJ8Plo0FWeIAn94bkdJ7Ot8dwJArMbA/bn+K2xdyN
VybL0z4m+H967jTeTm/KrBSRseLt/1Vui7/y0Wv5iXGDJ8Jngj5taAABUsSC/C/XAyI6+evEk0Gz
bTgMmc+qn7D+RMIvYLIsJj4LtanQzes9sx1RWgAsmpPOEm3zqCcBvdICxueEkpqVMUpaWs/9j5xE
e7aYTNfuJDY1HMJOKqvVm7H8AKDItWXZM+wsxIvIHGGtXuSDwH9qqHS7czQLOz3bglUFDhhKOEgi
VtWuzLmWsA6E2wWGoXxHhwcvzTZnfjiBJ+/cUaUtnuoehcd2f1gi5Mzvh2P7CztVIticPOsQ/oDL
zk2xSqe4+nYrvdBpM0jjmbr+ENLfUMtmxhhHQCsA6pQ2+IwQw+m659P/bwnwjU5iFavNUzjfTnZc
aEDabF2jbvzAmTEnuy/NJUwJH/SNldBtFfarVRsPsan5b39OOS/rY1BLvqQRtZz6b2ek/LUuKDcT
GWiiw5T2qIIZiiOTRIEcXh7SJny9KpGwCfPyZD3TWtT3TDEWs8JOq7XtVc4G6p14vdl+wtMnWCSg
My3xOD9bPIH/beN8iMWTPPPIyhaKpNiNvar9lIuql+qK2Bn/AAzaOBSIhNZbLJXMkuotk6AlcmB+
8J8QrMWa0lk7oNhAnnOcId1YGgd6VDkGHLFnYKlG+uh5R5hcB7ykEMP9YE/phpqBsUrWNvn4jXxC
3I6FVLV0kWvJLrOTVvDF5x18Sx59XjOgdHNuAgOgrkapwFopVAu/9p44NKvO8kHzNUbzoTyVXHa/
vg2J1oaJQHW3+nhxj58hxutwjhc1avLmUMlhnnCAI+Ja5WFSgAyJ6nwgz2hnKOc4HWVFNZJC6GiC
prDz06tiIv6vL8cru6YLZ4/MdykRz2JzBIwHIyDyqIohhZi/G76px3sr8t4qIYJu9DYOnMsYioBz
ZUgaVaqqhOOWYcoBIlmxa3ZPhbBQOF4U33fA22NtNC7gzvfZH8wtzdXx49vmeLS0jJjsBWxKs3gp
75a9LZlHZonQKw8+zwc5D90t5nFonM4KD2OjJdEMb3KPz3IrHjbjDxYBTEa1joyfS5jrZ/F1Upf1
t23F2AeARuw8bqX6brMwZgpxSlQl4Sgq9uiwTv/aSW+ZcCkJVdL5u2wpEPbaXGI5cLGtbuklFib5
+J2crqfMtNKUwCa+utfFMyYMgNdHA+FWoM2k2YKB9APzwHyLh2IeQVBWt3gKyHzQFBT5iTAQ0Ody
DzcxJGLlr9ka+npqWgaj00SNfalgJ5+fJ6w4wOc3k5QCFH+iWIycFUMPmapMMQOqiIolQO12JcUZ
LKZEbTxhfbrKGDo3nAjI7mxmEhRtopYnYdM2+fdzyApOnCgt1MYXYpJuPf2hcwWEbWdxaRc74ZHh
2+qttiyQclsxdR34p4hPGsNCSsxgEoaSqdbluKYK4P94U5sh3aZcbbyUA1qgtkYeE6hQ4RmJ/8Y2
fQooVMmw/Xz3FhPrJyxCGOcxHeppSkt8sTsy5haW6ezwHZgTjNWQcT8QR8mTAoayfrrAFi1bmZdX
uhIYwC6jBEPdcsOiosSWGl8ALATF6uxVp0XShAz4XYIzuf4rG4ZWxpN3+vzZVDDWpVXHmhvuZI0y
cxdd4jt5Cmxa/6j7Urvcajr2N/i9BKRxPq1QRNlJluQxQDZ3h1ul00vr6yrcSoXsChb5TbCiGxFK
7S3Al0/mCq7IlRy+h32iALBNAqcW8aikGCrrbik/yLF6tcY28e3VWzjh3doeoHEjT/IZHPC2AUrp
PBfr+tBRIDDpMD2Wbo2PB0Ok0w8d83jdbnys+EF4CCiIGTpOWhFaQlLZfm1tgiZRChfwvxrS/8mc
Gcx+SJ+LOfBWuTqjUl8bAwTuczCz6wtNqiPFRr6do+oTSMPMwHZl967VoUXCjwtfXGZnJy6QUoKR
I67SjGGTUEdqSYeAwzVxyh/VzOMuJTeOoHWeortJb+wliKU+bGtGOGmIu7Kg/dqZIPi9vl8CaKMS
+L3977vT9LAw3yesDD5YSFSFv02oGt9/sF7N/YoK6sNZuNGx3dw9bMiCpiGpnznnLNshQI03ESuN
IcQycqWnGPTlzJ8gZNOidgON0lB+b/6aHOc+WSHmV6wKVCYYAqbtrOIcby3MLQ7LT9IL1TGkbz9W
6AcyjW+uT5FZ9wVbjuiM+BccUM7jckblhYnT4Mi/m4e5HLfbE8uAYNRX4WcCwTsoMtGMu2e6YfXw
L8pmJQ0k1+hckWwVKXJakrDN+Fw5uzC2YrlEjrTU7zbkhs7ynn9azo/o1V1hAPenEj5x84MZtWme
8MtOAVek6Hr7w6Ab9tCzHLkaQurr8dxlOiq28ZrV92Qy+xzdeXTbfRviPl/yXP/DbhysQlGzEzLP
ZzZEXcjCAq4okHTYQXFydPABs87Mnv9JhKBP55PzPfA4/zk0dHxs7qwJ7AzPNd/LzLvOHqKeYFtr
LDfi3ynHx5AC1rBpWMiV2QQPvAXC4LZkN/+N5blraLsyDUCcaT9vkfW/xjyrv8ziN3Y13vrAyU+r
zWnGbcfox5V9ZZCCkpGp4fxsKAUn/V/Crlm+KJD43TQI/p2+kSk/vuIOC/3s2FP5rkFVi4gDArIv
MM6DvJun3ozLIQNcF0X4+EB8s1dl4yoQZ7luWx6CuJl5KAWsu/Uc5NYtvzI/tEe9ztEHM5QJJqrb
e/9Bl7i0fYIeb16CbTLiI2szgiRuIvzkB9JBzfzP7rE7+TPKSzjf5OOnVTAXN8wW5dwnN/hWf/fJ
TDSF1psyxW0mGrWcGY2P/jepxniiqhKXapn7BweZWdtnsxIzkESGB5MqqEs0DkrAlb2FZZath+Tq
r/teBWt8HWQk2RZs77WH7nJfOKdZmsco5DmLP/JZPvkyOBkvwtSP7qyMkBUw0Ld48USqcq2Fg0aB
d+2UaoZ1g6cUkExJrYuKgk51iCIgbx+Iarm+M9iEoqYZehUYHFWigR34ikuMUuwsCOB240f1iMl9
Waiyk7zFI638r3+zGUFSsrUaKCHZ5APtTcf+9ZueKNYatjaBSpkVgAsI17sk+Irk/ODK8Fn4Hf1n
IM7UvASh00aRFW/05qUv0FZSTiK29C20Dz2FW1VipHZbixrnHOXthMVHuCO/8QOMkGtBnMkaf8cI
TNyXOrTYyQtMY1st+D1/q/EjyEDyAdKjcn2HIg0YlO30+0ADwqyrLZLAj2FvxkajGRBRVRR4JloC
sKOv2bN9TAz4zjCB5xpoMobJ0DPib0jYrP9/i+wd5UNEtglz9waLrhEgACXbSQ7ExuDyvT2EACcp
NdQ+ZZRyx7ilwRMk8ypNWNgmQ2R36yfrqIwXJlcXozj8rVWb2T40KGhYAdY6w7zF0vsj6JlGWzRn
IvcXxF2BnMg3bBEzAtLelLP6oWz7eoe+wd00N5r+qLPF4v1ExTfI5WY63pY8VPQjepwA0iAeQCEE
6CqA832ITKS/tANY9nXxdRTPb5JLWsfMF1tIHCGMkjmRUORNDIJrQUwvvenQymTRL0j05p8uVpIK
ldlgusIAj6g7rEeZuPoBG6fRNf1BX3V8Ye+JXCTBpMh0q5P9Zbdw/LRVC3zrrFp5Or2FFZ2uKaZy
NZlECKbn8kBa//5w0x5DK+oMHTbGzW2vWVuDee5Pqn+bf0HW6kz3oGeZwbheT5OqTjEIMqGJnj/A
Em5RcdCiqQwKaKi0Grq8KIHe9ES5PWV0/xjVPC0ykFPbcPZNylpmcJRYYgQJX1Tu+L4re3GeyrHP
pfXzEwmSGqeI6RquOthrrXA0FLj+Wc6Wwd81PVYD0VOw7glZqPWkcSpR+Kwz+GgkR9Ax2UDyJTRZ
aTB+8n2BIUs04FFXdqoD2/hYNX3yiuKKsUdOzmEvMAKf2OKxQTlHgAetm0BcuZhgRHjzHQf618QR
65QOEn9lBsyah833D16ZAWxonwCBQ4RDj1n0M5ORqrLWyf+6cVpxYNiY72pThD6LO/Jvll/GkUD7
S3zdhaQOZr/zZEzJ/rbeqs6XifILKbJhCxhQfldCzrktmbokAVYQmGxBTQUWLLaJVqNrsccgtlbI
pkAL+h4ChKF6RZh6E/pxo2qHqipUsryYXzb3hrzh6SqstYCJIg5EGFRZ6nsVRGB+wgo/bGXOnl14
xI4kZGaKnR7kCy5bG9bMJ2punj0lUtE6CL3eHMZw6y4jKJ1FO87XoG2ibE3TLjMuPt1u8PwjgQOq
HG4K8rUE/bADsuQyQ3n1eVaXbXilK/OB5Issid2NPOTrhbCj5bnAxjqCw0EkKd2L4WMhpG4uwrcN
YHxMjSAVtaVGJI1tz2Cqdw17+B6uuXmE/guql3n6UnZFCaEJf8/H06GsEf2cph3+NKiY0YNWwOkB
FdQHzy/v8orbe81L7spgElCkY6rf5A67sE+yOxpc8E4iZJER6XJ645gsetrO8r4DbvEBmq+Dk2cV
2P3BgES6a4v3qHUrULAbtq6OGAlobWn6BAHmS5rqct6C2Ps7hZJQviOmZgkUE8aEEN9kHW5vRIT/
+CtEeXpGBU+vtKKv74LHRjqmrFLLrOn+v6j/r9on0wNoeZWynQN9U5Hi7NCuTZufImE+W4HA6aji
CCdRa+GyMh1xHwQuex8E1ZyJB7Uv0eDztcCQ9IN0+7Z9DbQP4LdcGu10qO01K7sr3HSWW6QOtwXT
fxVtO65pBZKADpevxJ3t9DZByejt3xsvqA2AL2G2ZBcUJjItWrqkhy/AIqmhFIxtucYDN/dqIOD9
1dnYpRvSaQHxShmHrhGnB9VNVsKgDy8OH88avCR66Otz0XtartN9QmEmHYc8YlouPKBzi0/NNmao
ZKxsZ55nFrDNnPjWHS9F3pQB6kf4iUVj9YtCrf4uEDHsSKpEpatFf1emZu1sjT0YVk6kSXr1te9Z
0n7h8KkNTnJgWKFlRtuj0vyO0kpUWKyQtFII0LoP3+0YYOYvv2MCNmvZ8iM02LbrqOrdneAuwIaF
zYos+SMMVEF8+7Ayjdt/FcHmkFB/Px2QWONiDfnspvCXYzx8E3K9Zln7k38Xh09QXKAL6iOFrv3d
NAGSnoDKjlABzzLmssKmSDFry3UUetOgsaHpUr4xgF0unkdGZbiGomJpjS/hbb6BcqylLyHgTSME
fU4se3tzUXTNrU5s1iey8H3hDSAxgsHRiGVqmG9fe3HhRbGv69be9AuWV/4K5TPVkL+czpO0TUkC
xYchOswQkLoZkLE+svBCGUSiujywdA8KwTzngW/8r66eFgVx9fnvNU91SHp6U4sG0nui5rMy4Pyf
59BWhLM30QW6q2bF2PegGex2H6TV8QgaFv6WEDwzoST9ioIHnP300AR4oMYH54FHROJdvLVN6dgw
Ai/IFW53fojwnhlunLuvBWZvovrFQjQbywsA7jLNZWLNjJ2RY+WrKB0hc2l/6zOvitaH4Q0Mn8kh
3aZaziOTtB7jeV8HLu62pt+WB3PGiBzAmBe3QWeqUvM2Y52V1yEj8t0DZGmCI5XZCAF8416FAOrJ
VSioUnLFkWaUoM9B4M5JBWCHo8fFNS9GbpM8tvpBI80ytpFNT2reB+HIw68gaLThWGdecDd5pnVM
/8KfFBl5fEdYrFInrAuOoh+5gQeHdI5qUznOkbkfhMJHqXBq7jVCqWlfiiZA61s1GXTfJftHshTN
Af6NoRmMOJT3QLrWZwChvjoJSXwx3YJFQKRynQYS7lBtSrNP+AHgplBBeokZkWwgir/CJdiIW76F
hyzxjtaSLyggAdx+VXbRAtktJ0M5sZ3e9xUaK8bxm58Z5KB+2xFfNW35OetvT3BDTZab16rm+aBN
Bg00Z/PR71jnS3Jk7C3Wob77YEColc5/Icn0V8JehhBy4bgbm8buljMEb26ljRvXYZk/unl8UY7B
PtxoYELRlDjkZYlj/zcGNW5hFuoBtbjqOA3w28aHWpbZg4vR0Zm2Xaef0XLyN2Oru5db8920gQaa
a/6qDB3XPw63jTPL3QIEJh1uNnTshF47H59b9OEvMVNGNn1ykapDhhM5Y5Fp8pNZkwKsYphcCwOn
wc7kgv3BK0k/4M4yZIxZzCXvzjQRGOPfGt+aCYVbBseVm37d+0AQTcamUMO8ua7iM1jyii8JiLdd
sHlBgKmSV/Mz1J0uW1f+R9t45wV6UYYsIhxGnMMSatvaDSiKPzIwQdPqQB1LGwNYqpIkmnGgoVKJ
xO40TgWnglXEu1Ll4IppZFPmGLaK7AVFlmRwVFyfx6026WwqRM8en7Msp9ciQ5+mpcaFJcKDZY3R
9kQZ9FDco8CwKfaLMr+lCszCDxZ7YYMQnJ+H0n4g2Ekg6H/U53EsqAjwm8IcEtaAusZCYG6MCvsw
c12bGv0EzwaH9usUsXFSgAm7dVexK2ywu+5Lnt+bHvu1XdKPzfNP4St2s0JGp1CnRfrXoH5AreYT
zPeYY21BRH4Qpl5n7cjSAZc8449mmhCaW3IRuYms+BixPC5z9Kv1rVhVo+C0zzvB2ykRigiR3Rzf
DvB88mHoX70s7CURXzdrVhdzD3t6ALNZtebJILE9OSCigYERXOhixNHoDVOOPEZGZp9SZk1gCW5D
Ttoam80EHuy/JJSwelF4O7vbZnwi7H4EGV62KVMtB4AZl4EyMzsR0VpQ36wefHHrxWRyeRnq5gz5
qizLPvGoEorbqQZedch0rbjU1l6+Q+RbrgZ+LUb6ePg/KHCnU72yX08uwXrvu2nTjbH/FnFfWjr8
DkUg7dgocxI5ALqP8AtG6WymV3iT0Wsn9ndhYZ9D+8M2haxyfzBr8vcva0qnudZF5zBQrbN4z0DR
5ffoaw0Fu/8iS6EpeDS0eUudq15vhtmR3Dlmyqhz0JqcICZbRgZKeYSBjacib8pAtdfONdjFHmn4
it7HwZIiXzDFg4oqE5zHx3zNmbpc1IQWuGoBfwZFUwxkLZR+N9Ug/fVDFVorXFNKJh002ffF+UAP
F4v+7/oxRYLcDnLhXZ61zVvk8oqzkM+xPiCVPEc3CRGfFMmRZ2yWR/4qFMIxgijXwhwRl5BNxn60
k0GA9unGDDVJonW0Njw6m05pJAeGYZgFBuBquHy4+y0PqJXSMjXrWyRhzxcSS3buM6/1DYQM83Ds
VHKF7LwnlxykObW8BsbatL93Aoo2gA5EhpPuxG3Qbhwr/2MU1xbcXSW4IboqPm33P0m8rNBszHa/
T9gPZsin+qb5bxWyzsEQUxyUG+q5hEmCN4JliI4/ifneBw3vlPCqDdSLdsSBwHOuHgBtfGxMUFL+
bPvG8E8gjLSG0yE66iJT1qCp7nTumL+qBebb2DnY5lpozrBpa8KNWXbJR2yzmEmPvHo7mL9/TcbJ
sAk8i7AtFEZ9YkR7dqO7aQK5MoQsWlgCwebZLlbS37X3ZUlN5uvr652ruzC8C8xtpRX590NMF87I
25McCJeKMqphOoQkmyAvsGnz6kmmAIvv+ZW6L1iD+lgcFXhmma8wv03jVkvOnS6Pd8yv4/5EjzsT
TLkMuleNueJQQAQnuDTXaiqPv1K9rCo2QZkv/Ey7r6p/5l/3jn1cPOyJY/3rnHylJK7CMv7Fss0C
WX3JOuwqzJFE1DDTgurG9tIkdMk7uVxbwTMo1TFSWXSJp4YhyY6XM6yJxFGFySzjFkGN34ekHa/e
jurWxHC0NAQdciPxsxX+nLW2hIYHUWhjVKIYRM9UFr1Epw9Ea6Q0GpqstKnbfjlq5efPd+y7U6cF
K+ml8ite4c+kp5t7VWlqaMVaUH/moNcsygV2/4tdF7C94trgZ4GYRRXc299CdBtJe/BbXlBg2zVQ
m/+bMj8Pq7PETW+kJC0NbORjNoQNAnLdnZM8ZXzITLtMRRQAtllmJapWcQO8ZSHYCeQ/SiiAI/K3
gflbJ4goVdQwccFMuVewShu7jy7cy69EaTjzaOrPEIAtZw5569XupHdmL+J5NmpCne+yaBWjqYG2
D8NE0VJWftTMNVmBDmPZAxnAFEMRlo7ZYKyOtgCwFWOD2CjFtkiWkUSShpAdJaYbSFPphapJGt7P
WydD4l5sI0v3LQmI7VanKdav2JlovPgw7Va26w8RP/3kd21CaC3dBICgorpXSpjXesRf3Tz1jtgC
JHudB4v3pXsqy7GJwtjay1UZ8Uog3NVrjAKo/tXsed8fkgMVqamZjzbgI45mcIv+V7FmbiSDBQ8C
jlifcrpj5K2+84uIW4K2YPoEee9N4SjmPCgaVzIGioalg2N3RjuxCC/X5kbeoRxos2faM5wPWVK0
mqnzghHEGiRj3IHxpFbn72+T5mTbpdA3uk9rJTYxHeVd39wG9aWhN8UE6PYtkS+Q0CKwnYHtmngH
Tzk3pZHRlNUPvYKxwluYRemAwGxvFR3nq67TsUjdXXoBkk7ZVGKPTKcDmb5rrBu5d5vv4VltQR2S
tc8opxbKXv4zHjShvdiNsibgxezzIP1ZsrrNezjWeDids1vI6DWeGwTNT2GT3JANAwsrpeycIgvu
BTO5D2KopS0UHFeLLGcHqx1rrUrqkhwFyNNliDxHDB1sE7g1k3RSUXkQJAZ8jgbnzchYlVT6YIE4
2rGadjsa35HqmhyfybAu3kiAbhIFHoWUotzyTMhkomNpufNbiBOUYnqHjXS3pNJFVgUB0sBzel/A
cptUfiETxlbFn7CHIDOk9mqPw5QomLcIdGv+MmG7n/ftQIacvVtsYwRFGqLfOGuKbMqc6yeXWp+m
Fjkgl0TtwmL9Rfmw8sEibKqGXYvHeS8ruchmJ3J31OSzL7dlp/Df8yH0ncUHQURT3Ek+Rv1Oo0sf
GtcSYItg4Lh3COyGEFKMHXKDHk8p1pTL5t062jb5FxhJkaFPzlS9X9+B4qYSB5qQX8m2PFGJeqkQ
UTaeWyXzPFl+uL3PF963CkiqngQUuRvhp9fwkdChXIclHybCMM3XU7w85xNp0FIUO5mInuVkdOfD
iZGDUKNDoKpFnhGSemJi5+tC3tJUh3yLj5FBrah/FVxCklvr18slUHEKpbXKTaEDakY1zpWBPzep
l2CQ6Hd4v+A8yq4r8i/vYQ6iFNN9mKoIcQdoJM9sSkaYaiFt2f1O+LpDUtSEPMrK62qGI9VCl7Jl
Ysz1tilmcI0ihZLnwmYsGuWtJ75rXGj8jmmHoWrQm5zskjyWm4VESivRGOf7DVeqzjU1qt7c1DKI
u8tWH6KTToiRVGBBm6YXXbpjNoe+wRmxSqxxrQq94ZsZ1sy1z43VRUOdO0WIBqX/G8gPNmXABfot
03JVs38g/aRWEMuP2FvvfnmhuaRi3kqJqEv8C2Ym/fPY3aeAo9hJTnInWaAMeq16RUoC35lXrndE
oIoNkevQzoooOerpJijUZB8AZiaNr3iFlR5derZIVMkLJnX4Gfpa+zzFtJ1D6TwuPRsmZNPPR/E8
UWpN4yBLUyzYva6MwouRtSdMQzfin57jkDZdc1DnsHXGNVBBtUyJJOuBBXg05sgytzy+0TCK01HL
BQhDrYBwCOtQCgFvswweFh7iQDtbFI3S0uoh+V6ULpLsruEzBA2fx4VohA8Abnb2QWG2RVSwBJ1n
YQEa4+sHshOwgBoLZWa2A0KuEdj/y4bDCYjq4zeGf7dLXoMiCbXyGZZTOiRhCw+yGaY6t1gscrtl
AdsB1SfEMOfL+JXWkNRIN5q+80CrQAA3yHPyB72SNmboJ5tgIDwBS6l/z1vs89riqdt//rcRmpO3
AqaV1oE6sTwBkg54AeeBaTuWQOwwLhUAhjeVVEFu8fQ8EXo7eIA9DPlFM9oGOwsDrG6WnB3s4OMF
b43E1o97UiFQlQaG9QDLXu1RGthKrWKApf3G6Emc30/Jkk+9Xpw33FCYLRsFE6q54xo75Z3XL2mc
376iH5J/h8CyYWGM+mGTZJrcfMDsg6wHhXNNHi2VWzyL54X5AHOaV+ju3Y8FeXbiQdUM8UWy9gU9
7uEfsDgBQMPllngFrOl6bwlIZt1OIMsQ2Ogw6r1tPfDIpYMeUJdIrGNMl4+EtuJfffbO3tHzo6UN
745doVLcPRJ0Tut71xEGHlKDlLu2GL/PRjn1rdCILW/y0Hnn49fzDKMfi5qzJ3UyYlXTo7uHGEoA
Vvt/ZIygatVAS6tmW5aRInAnNmgaXDeDZ0LuKjvk4+XK9ZxXyBb9G4iBuCXMJsxE+p9a6y6+F2sq
0GXdNU5bYw95zeS/XMYifovFE/7mu9X8Ouqff0GcZlTiFqzh6jAkohY7EtftyqIQsLM7HS8wcD4a
d72R5TF9Ob08F2W3HpFvSI+X/GAfiS0AmPrhIEw4haJct2dpGIxS8xGuLxfDBBSe1YxAI4nr3DM1
QlvVNwDKaBMdgvWeyzDFwe4rUuUlBxMkf/X4SjqHIlhCbre5I3A/a3lMnr3WfsiqMRdjHcqV4lrI
fs/i+mEPx+i/gvpUpHTpts189kc1Fn9jW/CoVY1d4aZgqHaDV5akHXa49o9bVoeCXWaT3kckf7Bi
jCtEC1BHgkhhwNQykq/t4pb9OXr3hiB0zbUtSDLlfqYZ3TxD3zk4yRPMxK8Ma1M01yQkquzprFgj
KFvJbOLX37Lk26G7K4ewTr+OMp5kEEyWJIkM/RVp5sHWIBMfhPfDJETim1Uq3SieqQsn7HeDmA88
+VbLJ6TWeozOYhbcNLSr+W3a28gsYzFGgmoqwEYF6cmvocCfPxlK8MFJi6htqbg8x9JDHtyaVt1F
QUdkrsog6+k2Vr2+UoADIBSVrIp3Z7eGkHlQQfCOXLHCBCen2uiqspeRTgdsB1f9QGKQvLZaneNz
YO0zW7aKQ8C2WU8B8cWTLy7+kSviQmf4Fi2m3T+BhH5gn7do9kRBGl3PGm3DrDQY14b3PZsS8ngr
bjOGvWSozlvTcFTSSMjBdLPcB2WeTEtvXGLM/PHaaejiLzUs50GLXawMHXPfmulKBttAZBf+cto7
QE9c42w8r2bVb9yhUQQTN22dL4pE6iz8PtslYhFLuieBXdRREHF4goJM8Iv4UvV0m67zapf6iLek
4GZTlns6H5N/9qz/9GtQD2HLZoqLYyEMoaer4ixSzaCHSGmY+nTGAV6+hH+Kz5+hHEy1iAWnLoXb
Iosax7O+4O5YqzLOWCrmyzb/NkH67ZElY9CzzAWOrLfa3Z88u3z+zTvoX+40xgyvU49TVkGVqebl
YTlgzlkcQWoeNysm4DyCzDN/uDZkhE9c74azhirTuHgOrXJ3CS56RVtQhnjl2bPu2kYSKfijIgw1
SM/2xk+Flpmrw9bhcHpUjOkCV3Vl45luqgR5+OGUEKdYMU3RIZB8ezDw4naT2adwVpqG4qMXH9Zt
Ddp5MgzWWlLQMGYTKWcw1UMEATUj/4VrfFsaHUuswj8eLee4DQrHBqYssYrwgrg0mbP+BIwYZOCJ
NNhgWUeDLoNNLIFwcT71Z7+7j3FVT270yzqzdUcOTTwrelYZ9cpZgt890spYh9rh+y2QbYhkMYCv
OioxrpHm0IqE20vvoFkQC9BcOn+Wt2Ye+3pRCi1tSBviYEN3hgRuuNb6/x5wanVifhsvgxvxwScW
MGfir2BayDEjSFN7UKP5piy3pDVev+dZtF3DTDGWpH+/T/9oVw7UhU+V4M73ZlsJ7i++Zj9qe0L1
e19dxggeUcFmm4Ir/iC8Gzai+Hire7v4whFozMW5/W9t1fIAqrEUHanaPjwa9js50BueErO3M/hQ
Yj/x8dW8Q7N7bB3K8LfiLCkrEbGSj23qdEFg618ZcVrdh+XYvoemOvhjsEzDn2OAECXblsjRPQWB
cmkCld8E2Hd+7Xd70hDXfrtTGEKEfc5E/hnOlyZda+bjgyG3saM2LswXdubkXx7EoAGVCSg7r0c7
NM/gViXzhHGdrXOEQ0HWomjvpp/1y50kzf1wbiaXZZC8JyRPxRWSxB965ikA4gHaZDWusfnTaa50
owT4FhnKnIeIc1nhpa9CFsQ/1tM9Ppdz4PqmEP0voYZAwyx/zze65m1diCv0gEu5tYxEi3KdtpJo
HdvdrYAnkUUUOkcJ5ZVYDP0jHyWHJDjwIQvtw1pu8w4Ih45mtxwQy0HhbufhN7DWf4Rwy78JsLOQ
S8n/bIQq3OP81CvzQo5ReEZWsGUe+1e98KpNULEccUJ39byEWOdk/VhmW/TxwbM06W0642W3/4dN
IloRs2qcecKgWBk0A09QU44auQl8SbnrdVNpGzZff4TFqChvJ3jymC3Efdgd1TYTGail/C2F8f1s
3SU4HX5B8DYAciXbpowOLGgIzry4Y3buBn+6OR+4tuGrNu0XckB7JOE3529XIZMoWPFdCFgD08jP
9FIYkTe4GUX/7rsKwdUVSJH80AC6yEDSkfhk8srRkKgUoTDztO9DischiWC/nCaYesASV9kD9RGn
uvbYoTmaa465uGiPV1j/JwiaCNzq2pnCxL+UMqGy2lHQuZENkm42Ih86v8wCoMHCxpbr9SxLz2Gu
YNDmlu0rRTHID8mEdQV4SV6FWnh7jFNCCQEk4swjco5L7NijRzOavZwEUYlU9c+Q/VRSG24g+pN6
6w+zdvGXJk8NU8inRXs2Bm9fWzP2i/tIPezf4QopvxxvXO9Eyn3s60f9v8hOiu7agMMDTY5cPDQ7
lJN9X4dKZTaxL+dKXilefcl8xDvhiRBAvMCLzV9vi4ipmW0Ekau3jb5ospxbeKqonqYk7tAqUoDF
hldDjav+XtrD37Hk5xB8g2QYYvufhY2HLnqfzQ3Q0+hAAyLY8lKB6q2GPFcZm9q9N+1zjsYL++TW
WY3EjDrwBXKVjqPi8zbr4e4Yzo+jNbEeCyPbFzsA7aWo+JUrf8vNzFddFRGgTkoTLwLvlOpRTFX4
obsXWmVROzoofgUMv+m+BXVJF74huXrS5Z09O4ZoqTCxqtVjZs9Cn9NAwabd0/FNnL+reX7rX7MU
HbLw8FdYoqYhnyw7jT+jFb4vSHsqWquCXmWDVoI9djhiSevqvXZSDiCAutbTeITmd+prKObxTTf6
sNxHYP6xwUQk1qFHYJEu4CvFmjfQVkKiYansNKGecgjMciVWStvo6dMXquxtBjU3pwa3HtGfx21k
oIDBul5O87uqOkc/LAbiSF+ecC9PLcINtT4dHLzfMCKm/vhWaI6WQWifi3St1YJ2ST5egAyrjXDD
yCIprKGgk1cvnA5NsQiJtsuhyB8XAix/ujU8GvdWgh0jq+jmVVpHI63RFE/5hVCMaV+fZuEC3lz7
//EyS++OHvGR+immFE3z9uzHmdYk6gLqqGwBncikNVJsE9ZgWUQhvTqFRGXu/b98islbVY+cwQdG
mukKkfoTCixzMHWzN4xCiPPB/pX8P7C9Hwi7fzMqdGtPW5Ol1vDB0f5XUS6sYdq5ZkbU0c5KZ22h
sC3S2g8tmG79gJbHdOSd9Y1OQxGBluGoZl6LiufTizhBTm+A1XuipiD1/jbMku9VGl/chiN2yhYI
cZYXe/OVWJ6l6aisPYHpQioIANPR9zHansceO/GjAD3/+Hyrzn+bGILp70JlBmdHK7AZ/BDn4Tia
xn9Yh1Dkq+482hTVlivHJkYoxh4BpIh+NxD0HkSVR0EwfCzbYQX+2IKdlc2epZsSo0TbrkLCcJo4
f+pV9HI6doc7jPABKUZh7ALVEjzilC3+3PQwXiUSlrzscHIawkLjCso2p+VFgBZvISAKSxtxVAl2
z/c+Bjs7okzJygKTFM3ZsttpztoTjZjCnPpPdTxe+UC6OVYWkDfFodQ57J8QaCWKfqA+T+X0c6wS
wdlj5APZD+06F2caZBjTibEuKjDeS3OIUMqWEde88wKjbm7hfMGORjEKS0IPCn2ZZvYVygwQ8Jfa
Fn11f8QHhjRbDdy5HzQhOLLmBDmdVH8lO+tNmCy7M8J2ikDuS1gOw0tRn4RgLpA74HL8Aht1MKQo
bN7gWObo3tAAa6YxGBOJl9oFMumGGhatVcBGWl78YKfBhXMYyTRISeJTYrWTjiv1DiLBo9PIF+ED
gXrUqKBY2AsQdT1nQH2acLPEUsfVlGspMrqS4FEYnPDr2OeSXcaT+ttBxyPi24u+dHlGMAWSef65
NPb7FVGooszgA+ozQ7XlMROxgK52HtKq6Ja+Z8N/v2jgmE/LpXTSYr0fyn3k/KhFNxPz8oHaWYux
wRa2lSxO9fxVPyvh98z+O7gzrSd/yvMSZYNvuVERf8Eril90syUag8JcSxHLn/lXFZ3wKOdYJAbG
SeSz89/mops6GkJIz3ZOXp3d259ry+OCDmwA2Xb6Fms6p4m2peICg7GvH5WYQt4CadVIzhdQJooW
+p/RWZp35zOnZCtR+z6OZlAtTgypukUuq3/KODr0zXPfc/RlFymeyrRBPMG2WevHcZGjrwpCf0oV
Vn2uFPK9HFKy/y0g0N8HNfWo3+tqketcCR/J87PyXrKQw9gn8rZaxrzMdvdWRZzh62MIOtcghEjt
HryPeG/WoEQ0BUjI11qaXRVKErcpgG7mhKCcSNwXr0mngOp+Hc1Y0VHWItCCRFEqpjChRcrpWpto
sWqBeDDdOxoKd0p93pp8fogpp2qjXMBCUniT3ZsTA3DKXSyB4EiG5rIj7fwEkLG48M6aMckg2DYg
6OQxSdwE9O+qtWW3h+KHCrL2PODdM7b7N9wTjNz1epveweKdCgcHRAgEwPM0/QSSsHS9NkpqwXNy
3TnFf9nQtahV0nnRgI6cZUlQ24cigNoHyU1x/SUiroM1tYYpjFl4pczJBarkCD3voxxGTIV8kpuO
QWWC2mOYGX4mPwX/IKiGHTjNvnk8X5gECXjcyaKcZrEsppLqllhV+WlI6D4h25CwWe3bvPe3nLfK
khbRY82QSkDkfJux3IsO/AVB8j9tpU+MoQ2QJMwlOiD0+XUm9vYte+DV2qHkKc7JWMPtTYLboerl
FUN5Xe38CxKTDz/iE3NLflVaGx0I+PhR0PE/H20vPvuCgJiTQb1or+w8iz8SDfSsVFRGLCPwyYQT
mJhkz7L1mza+PpP8VLa8sdngVeP+2vvsV8P51UpMMqyuzBGI+80NavYGhdru54HcPmNocGAUyI8T
EwCrWRDcl79OCn2dFPbv8M90WVoBmMNdWirsKedToMPsxebUOVW1zo9a3Pcvpn7qNKUCwUczrHOp
cZ2HSO4zWruyeF5ZxPDmmawj11C7q5PwQGlYO8zwdW6vQJzXqv/QZyRH6IkzKGfCsd88ZWXpZqMq
dfO5i/D8ZsumWclL9LUbKRMSeumUAOG01Jlqa7hfWckVWA1Kpu5ueTEzN4Q+SBfm3gf9K5YmM87P
d3UQSZvfNVON9h4utRPHEdhkV+8x05H/C5NNbn1OGw4fFjbEwDIjE1cge+jFkKQNdpO+HYkDUf5I
Z6gRtTMy0MOdDl4CkBkxoAcgSEYRIuMfWnIaeqly32c4w+ylURvnSRXR9DkEgDKuqEUZoUWtoxDU
w4Zzis6tGspbUdq+sHhr390hYRJj7E9s8X2h7TfRGTA1KmRVi4n3vvrquVm8P/ADgod23WMQ0E3m
Cr2sgktyP2EXZ///f9sK2Us9GIVktRLx0/79XfYCgvSVTeAitr0TMNZh5H0OZW1/92aUFl2PMeRY
aGRw3TOKmivIKmmL5D7Oo49wkLDj36ck5ufFAvESV6GLbWjrcjNeOz72Eir+m9zhlfe8z3W4qFIB
JJAlBnzYdgXsr4q6MVTZgXPpq9WbvDHU+c3NCWLE4uQ+JoVLAZdYGMnrUbdNuevcL5JrGo9zQExU
DM6Ie747o4g3ffqu0YoSnG7UX81jXx9whfHMiWVmqh5b7sTrlP6+515y7+NxihEP0bhZ5WlDOqu+
qwBlfkNcaU0MZWs5zUPLlAvDFnBMSgqHi75I2G0L3LgAvYGtzQ5Fev013mJ+5OB3zKUN8AKh0Xoh
NuiW/NenFpXc4qfzRwfDYk4vw2jKwbD8AK3KIYKTcA801saHGk6uKFUjhth/CBNkmXuEalbuxksk
yZ5l9MurlLyV+kKfXZs9ZGpQGwFr9hi3G49V67xR6VsvOdz/YMk8NSnx+f+Cxx06kYw0v6jV0t7w
A8Lt376egSyp+GRlcasebSyiLar4SQXwbWYoZy8hzUitOU2LNpI3sUYN4lqgewimlx2jqK6vAzmw
7VQdYGj23gJR1KvKZyaC1KvkdgH25cwnaBsXwvRm2Z+8cBBEpBI0PjWBYW10AgdsdHe7DJggZx+u
OnLkndl4E5y7OFZ7MArJ57726NovtBq3UjuSRHNhdKqdVCI2HzTKnRERCjaZ3G0Te8sSCsWO1Akg
D32zlCCIoIXpMb9IjO9YrG+v5YmhTbvrQ6/UeX2f6xVTQkFgLGHemn0ShoVyv8AoUpqq4XiZF2vY
A1jvOjdhrvae1JyGONeOF6yR3rSIRQZwzm+mflWimBNSqWN0Ytpm9iU4GL4jjwc+qCrfmX9s+54u
xWCFI4tHrb/MlRrWBoZdCwwBf/WsMsPTuOg7ZEL7OxHHi0V4UF+M4dg7uTZ9CoQqe/arCibclSaL
0NI6fNOLfwESKLjgQSvXGHz2v2qFYmvtNw7a8GFUZH2qjSScf33jwKDfTYdGGzcKhL/ipPo4RbFw
bnjaYj4DleBYsGROVbzmVpJgB5bAs5wtiWT0WO2xfAGIVSBTpcvbYR+qJvdzuZASs/3fpZg3Em7D
GhBGOs68dTosMsRIyOS5aymM+22J3JPlOTsZTIc1p+E/kwHsFD8Bk77vbjb0lrBHZTl3cRhj9qCT
4NzhnKqg7AyXLIYq8LRTpK5vg6kAZ2Q9hWRxcJ/w+fUlIYDV1PUW4cHDfi6AI97FEI7Jgurs4LOs
nIA3fDYDYJ6aWeP97comEatOTnbIpDqIo9htYlDLtZwGmup3KjMY+WTjhADyaqcZhJ2o0LFoM/wu
X9BH0v0HE7U/u/fV0UHptsV2C0pLEdqPTYzLVE9QiGr6g0CNL1qarzrvMSVZeJx8Nz8q4q2RpnsV
MJ8I161HMd5Bl72Gz3aG8tzhfPcNEf8c1OIKdp4N7VFzWe1hjOCn9Rwm9FKX7wU6TktWauJAAA3I
RtNHd1+8NAt6ra3F+hRdbjTUg+lrXCvL8FdOnSt16CsszEhKs8QXRrAkVlv7KyRxqRuDisr6WH0X
mU+toR/J1wiFVkjYRNhE53a93IX+8EKypG4qXohyWXLkYYSlQblvWU/3ni/8M7DLYenhsZkj6UJ9
sbqV5RAoTjO0uluS3jo4iJ2axTRc1lM6g1KUBZABR1i7UAXhkLKDC87eZU7u380OYeMpfCH1H1Uy
lVAjCEi8zRwfLNbhyB6xjueWfuepHASaF94DMkLr/X2/je5on+Jjr7Gsbaov8stQgZOWHGwGAj//
A57U4yID/PibcTEdT7zNV3PEuNPWIDSqjE0rTEggo3WM1nIBp6iHVrKdY9UdYJrVr34Y1w+hRwrY
6IW2kdyhHqQoAkUViPd7bST4Hzb/8tsM/hAyuYSvGWiUfnL6tqoxbmf4nFtwWe7v132d3ldBpyqB
y06ftRFNCdSP7Vfai/9Gzr6qeTfrb6TW8Bs3EEYTlu6ICsiWxJAMByA5bsCNkyhZSxiPnYTT4jzc
fZXM3KMLv3a0wECSgf1Os6HBciuDNhtXRLfnVAkrL1z9cOqhM36GcQ1v+dPM/U6PhP9flu4u7waY
4Q7ASJhS9OVFILnqIlLOxLAf1MzgiYpomNAOyU6XSHd25d+6vDXA9bE0ZUV6ZIvLnVydux8UIdUu
TgqN9/KpuxIQ0+hhn7PLJ+J2AwzucB8PQVhBvY1kHFF6Mbq2f7yERfrFRGbdEtt8ts3LYXxFYrkQ
/pZaZ62kc8R+YHU4EYW7oBC7X5ulXTtS+KBYP2BpFEgLOIMtVkIXVWupkDSqeVxDnm8+U4BIR0jg
MdEiPFpwo3LfvCk64tdZFA8V8+y+0Vx07PfVPIZDy2S11diCyomSCFhPzaaF+R3g1prjtlqC1LyZ
XeUUH5UfDyUy4+xvUAvUda5Pe4dd8Xry6xl9cBMwlyUJYtMbvgyszvQalHbdcKfA25Lhc5yT9brx
ISDapWSVY/y+moCoaV+qHOlo8eFrxywFHItS6jqmsO2+U5zN6abj+b2uIh9vGZGWM7qz203+1NSB
i7MsSpT34SZslTci3AIRe9ZJvm4BCryo59TZ3VDyRoOxOe0EYG9yi4vxn9acHP14crz5FgLQ1NgW
6YzcDOEuq2+35ZE6+CIOzLSNkdi4eXTFuUap3P1j0wJ0Pmv3lFV2KSZFfKyS2HE1k8WHCOtEdoRC
G5+VaH8X07bhpM8ffiyDpTuxh6AqKXi5L1DA1FWyoeci+4KqYrTpsEd9b1fYHS+77LSgJ9Hkhn8g
dZGqaAkEnyb8AT0H20jAotnrpgd2Ev4b+Mv86rqZhz5SLM0lD33D9rtODdZZ2fE7GGoShTs5cjol
YQvSeooU/VYvqjWwIxDdKGyjT2aRiRjavS7cltlC4c5LzTYeGfVNNL+Gf9jPvqFPMTjDTAdZnih+
9voC9q9fFk92sEn3DYe5vJdwnVuE4hQcQATDYy3mEVg/Wqbi9nuOU8fdHoz8L0lbcUYHS5OtO+32
i7Ap8fG7NOHrLt1JyoTi8xSrlnV2N5G6WDbajszCGz36/6maR6E5Lyb+iWrJIP0PWsIC/YTkzZEe
FvP1QORljJENoCOq3v7WImB0xqAskNyWiGcUpUZ6464Geq5+bMr9hntuTtxeQ8Nj1xPtdlVcn32V
dt3Q+NVupctqczaTtXYcyvXFozHSjsSACQn3gYOz4rnMQ/H7ZD1+JrLtr8Myr8+Dnbss06BCxu2z
ovVt5QH791Ny2W7KNKASZcAhCtE5oFwjw4FbWDrT/MlQJOPYpbkrhCrAGKrHjYdfPUotQscrs5CE
QvVKM18WIavO/3apY0S0JMg1H+yWPJsvD/v8v22m0TjE/9tpi4NnFyYDXx9Rtxt27tpmpSx/T3f0
BOtGC5M3VBG1APP6MtbWkdFkwt9UKn6MiIfF/aHE0C9vRUbTsSvvNP8j+UDP7t1tVT6h4SnSIF5L
7IdwIM1hoIGronTe/r9aodW+X8IZa8BJSr8b9JHT93ARtR4A2UrpAEhVLdPruv8jHThwd2MimLy6
12RvaWPjcQ0nhppxob2oKzJVZ2nHNkulYAsH2kS+d6yO9jvDbtY0ZCe7n3EI7CTxp/MLqGe2ftbM
qGrRX8D57hyMH0RL/Ys5W1dXnfSzmwlI1VOIai3Avnuz+672pe3YCF3/QucRF38MDQsIX7X+rx2s
iq1deEJiV0QIjn6yZU4halvFqHxYB1mlj1k2CusPk9y8hmVAJ1xK1I1e9vNldkJF2xhCA/K4AASY
MmbBF3gTbWHq348+GpRneKrbsevtXqeQIzRPk3PPtMbOQpwjQ3ruGstRCkW12RTBFM9sk0dbsxpt
Oaf3PJDGMSCBHs2h5KpdRuKypvmwm866IFCUuXN+3fNlr7ccZ2vOV9wqxSNPFjCyAUgfDqVM+58W
0bBGudGH5kE0A+l3s3xzF4G8sQZZ68LNoahsTZ31NtoFV80tkHzQIc8Gmq7c3CnVORoGRWEUbQaa
MN/V1IiQqI0lILL7hbHwWb3+WVkG9PyLXCQbdmyqq9D34X3d3zwhEHkT1PyMKx1ThaQv9+hwzKJE
a9v4W/cmbxL67r80dtyZRFxAlBHRGP0lCTXCT9+E0+qMjfulje9vsrQ3Zc3/I06E8BevHBuWnGBo
hCaW2udJeouF4mRc5J7IBlQakh1Tw95FxbSFegg96WfMctmYqpF513ePAwlQ46ggKpXkZGGX9/J5
TILsgqFq+VH9sjMHeNE07/W67WdV5zWyKhJ0sUUf+1H9M7BENiBCe03xTX/CBFUg+TnKqtHw/La+
nz3bAvZywCFC8htFVyBsRbkpXdRJlE7X/524AOqcpUzwv4hRam3g3+2e3l9zFG9fHxLIYFxpt93L
l4ZhN0eV8XJO4h30ji9wjIfvbqjR6febHpicl1aNaw4kGjRzGpuzQjz9mLCE5BZwBZ3IoxyNuGQB
uJ8Cd1Zn/Qd3L6OZfRVJYodtQ0QuimGcMW+7uR2siacPvTjFCpAncPSflst/QWhMQlcTx49APP9o
fY0pE4tT/ZdlDrXmyritC+BD6NqvbF7RBff66mKlP85Zy80SouMZyP65JFEYGUXs2Ig0kGfAF4oe
2W/LTFBwlzyT7FdyVItBVNqRgve4dR3iXw6VLIf4BIx/LAgxDzU39VgOAR4bGLsxnN4TRC1iZP4l
wQoYAOxA4xcw4pn1Pe6lU49EfN+Dd+2r8js651RZWUrEddv4HmALQ38KT0wstEcTuTU530Cb1G2V
CkLAdYXlMnlVIVSS2Luu1KOJa69Pwc5+Hj+HMnj+tm/36uiDAbHm0FPnmLKnDZIIz5jw3ESVgQdQ
5K047qdIlUn05PQmS3v1yUXvfcBTVH1xZs8Y9FISn7h5gd4cUnFyWeycjH0NeCWnISDFT6eo1det
F/uFz9PTmDVWw+YKqXqzAEII/NzQJvIHvkP2z6nSQW7RRgPzN+Z7xim1v2LmAwqo+9iA0I5Y27Fp
7i3BGUknQuQQR2mYI3lQQ97hNYh2v0ODwAQNtN//VoXwzwTaWPUqTeXOaXPc5C7jkFjH9wwqN8//
B81w1cbhXzs+W0Xt2Gnthbn8bVfWFgOkCC9ijFYWLnBPn6SEyf8SRmUz57fwc5UrsBS1YRPs4hjd
Sjtob7PUkoiLvzQzufcvdsCmLUUUD5w25HzYI8bK7JcfhCci3xs43mV/5h3+/n0R3BW7ZgJM2ICH
x/H761XQy2HvKSnsrIK2Jj+EOgyYOoOjQ+HXb8KMVUIEPR7aJWKqkDvRjLlSG+rTVLbxhTiXB2w6
l7oWZqwXEsPNr8oJZdbM30Adl7pfua5VbZd62XDrYeT2lf96G/XwxclTH+yRWFjHSXDNNMuouKZd
wlXAAbzVlZtESp85s6HGgL7nGdC2pC/ZO+9EAVGABJJq3aOciw+BQtfRim1xwQOkGSoxla3gB5+p
J7QWSlqCYXdA1NmitFQITTWbp1xv2Y43P9bDDxoI7Q1C5eKgXjVuXuVs1Sbfq6jCI2FOrhBS5LE7
H4LZ2FyoZ99ka4Tx3e4ve9lrgqvMpwBjuiAFTLg067pJe6imVBeHO8vB2j8PS1ZebzlHfCfDg4fd
3C/CxmdD31fkLsBBXT6KyTf22V4yrvOHx7td4ZUp056ne9E1e3CQ6SOJqWKoMAd9EH000XzSemKo
0EDkQVzSTtRJbTJ6xN0lh9k9/Ihhj2ytIsr4XfXy/PFwIB1JQBDGZyKsNfvVJoTxGxT7ZG0JWa1j
xi1Bwdkn44O5NEjc+BFju/J1YK6BpBz9y6zqNNJp8Bhpr1+meGwgCflK018EPwlHRtknlRyAyaJp
HK3d4Oku1gDsxHMJvQka+CB8OAQaScbYp9g9MQlHrMyfUtYNEoN/twsWBK/D3zKfhRS8P9zlvMFi
f1g1oHo6kDS5Yc73wddz9yKmNZ+2fKCMptdNhxInshj87XbuMgmydXLpkdx6QaNKX6gaWJx3iUoj
63w5abPSnjmUhqwIM+dsNQzFM2DdByavINu5SNUwIs6jrG7zLxsBsypls0jO4BVLJAn81LH8aWn2
eX7AGkqb6lr3h9S0CyAB7TlxQ2RLHtcsoVTJ1m0u19pg3l80W+2p4w+HPVerhDS0TlVxNQxe7RtT
60ybynR1Aol4tzZxmRMVEieHZ3WEL4ouKt+3a9AS5Bwu0jcp9/FLngdmuTeJTxNs4Vwck0LDcTdF
b0Z6hweIYEhcsQChA0/lFzlUJICqrvzx2GPwoeZfRS+B1mlZ/dfkCH8UQof9z6zcfCoGqYxjSu7J
2hFnEHD9IJC67/RGf/00FAcyMIUcPJnKzbvBy+23bJjjjC7xw03tWYSDQrHF/7AoN5RKy9oq4Gce
G5a58mlUY1ASfcR57zPC2RASgbXHTVO9WJRKIJ1lIuBNPWXQoOYlWrBhT11k/gW7pDR76TUcj2lK
5EjC4sOxRUP9HkUNyxuiMfwd9Z2i1u+EoN3XdMJ3Q3Fdb5YJyHQvpjpbqdmUejuDixUFy8X+Rjx4
52eWyDXpdSQUy9lMipVP0ep5xqEQUFS6zAR9X94XMl5Rx1QxWMM9CXqLVNlWB3x/b6Lk6QHeJ8xE
vgG9w/IftPuxQ7ej+wYJtkIi5+cno5C+72KJ+ph3w3liZ7/CtVf00OfYRKecccPX+0cY40RFRg4x
25cIDHnQPaJsSKLCZrn99pcVRIVXFl7mWf+AY3mUe/toC+SEwbj0LXShGsynDe1Jkl/aOjo4X8VY
HEm9lJbLwVhoZdK/FaH/AXPMbgZvyiK05VtDVLUx0CrD4PvnsQm1ch/FFgf9rRry/r0mvtWnwSBT
6lBJt+rfpyTea1/xpikXcgHZxu+pwWR/0dmz3MAoGm65QMxWsaFgmrmpswreZPsagxhUh0B+QfZ+
+XOHn7y/RD8HD/idmo1EyR+h89prfoM6UfMurd5wPt1NFYHqKlR+KyB6DZWjFnR7Mkccb8siSLdD
BznDT1Lyx2QOnXAvzWOE3CBgLYhiu0+eYjM/8LbOCvCTN3RlSNgszUTqpbNemIMb3pAPB9Q88aPX
uloblGLmxGaBG3DkY+Jo0SaARfFSufRoxnFVEsQXZ0xhPr2jzH9KIhqGXcOWR4ExfSTpdN5fL+cY
Z5zR/RH0WwWq8hjTC3QDkKCq/iuqti5JZHbTS36ReA1sas9cziMkjTEw5PgokqvnfKx+gqCb9Njl
bKc72Orf9JXxOQhZz4exmHjw1bI2RXoUk7ZadraRIWaJ3o4E4fyHB9N7rCHJmK8VLI3zmVofOBa2
MhqHEdCNVMyvtZwp7i/WQsz6lHmlQVgu6T72VDasEkm9otx9ZKn5Z9AyhlzGaYc4tzcCSxHn0H9+
4lBQtrSTkD4LjHTE/sdDzReIXDrBStO4tW5bfwTBgPO/vTMNFTpZ0dJu+zELN8y6tJ9HS42fthXX
ZohrsTfPpF3U7BB2cwH7FVlZXuAJ0HQ8ElR0lI/5mfoLkC56AfiJIQjtsfwd9aCC/WoNRRVQQI5e
HuI1DYEIl2uwxAsjSMB6zEAR1Y50kw/zXTO6SnkEfidnl9E2tKDK1GrH/PEM84weRlADNy5UIABy
BTursRTBOqImd3MrCKPmf1nvJWjom+TCFSWUFCdCn9UMKn/ONJmUkG7+SdQ2UKa5exmF6FoPX5bd
OfhOaa69OSMcbxPCWpCXtCjKnrLhsxgXXS9icGwXgfuZiJ/fGQ/XZ5gF/5jheCz002XQXJHuF3an
C4CjtcVbkt+mq6Nj6CtUyjZbiyGviZe2kXlGPDIMh6V+0oR0mPtxbPrM7azaq9T+h0LHA6+n+78+
2wXP8CzcyWHk+AJfOyWur2+wq+Jsf44Y1W8ZdSpiVSylgLpJxHFLpVhZFzvMgS+lw1aP9GPvdyZw
0bdFaNligJGpLoIs6Gts2gi1qe2OfXJGe3R1WeipyUZowQ7GK/GG1xEnrwYf9k2ROqDkPkYByV9w
ttPEM3Bx7FHTaJFPVMZQQi94vm8oYPonlyrlrbwmf+Wk8w4qLafA9bvK2VoPH8YwOianqfoyi0nk
qLOX/AljZx5MY8z68RVgt/UJwJhEmd1IzzJbLVNf2WQ7rbnjSz5f2cPhxWP5oqJw36lxvk/BTZge
jWKQNycf6mxFY0UJmvieeIyZDNyJmKNtZg5V/qjbSpyJMyX+9ZyLfGdBGzYJQphlwTQV7w3crBEv
STVA2IT+NceBImx3F2oCME3QBRsQLqs7fyJlYR/m1b+TRmZIjeKNm7alNEkVwVSdV1GpQRdu9xdG
ubufRxBu+qYMX2rMSAz0sk2rImGDZxo7xVh0wpu87ECCGgR0vkWuKQPd1ozTC0S877knlcqGJzw1
8gI5H0Zw8nh0/H3qt+3mE5BkbLvbmj/EIUxszSDncD0P1fwZaR7tFtrAIroChUm1rxuoI2BH7dsK
xgJRlkaqdiemXHBUV1T9diYWaUnGJvsFqiNEiG9GHzPBnA/gDKLgsw66VKjcyqp8S50xbCmbW6Dd
UcjD83HDGd1CyoPsjYjGpdxTpweUTxGvZrrAx3LD49Lc4y0DM54nXjuUcvVMSsftRXXvRxHltHEx
8+r5BTAlGQycoVZuExHtbeY1qUrmahUwUVbJx7J1WS0G/81VqyroS4xyvktWFDg04RVnplTSsni9
O18xAPRV5/pHid5qNDXzdCLMpISCLs+j5A7E9O3ogjvlssahWFY/NBnQAC1mWFoun5iTZoaxQ+u5
Z7JzB3MkNc3vVpKd+abBcVXTQ1JEEzjZ+m2g+Li+Kb2mh49Kpu87CE+ajyCiK5b7BFXFdNwO2mlN
G6ToQlhxeE95EpSSQ4oJgdv9Pa4yn8+/b32h1hmiUtfjCEzr5swgjgmjG/ZcTue/FTJ054hrvscJ
9WQ9KJkwoy2G9IFWx+NxUBH6fIG/jF65ixBT3j63fulYgG4KUb4F0wi4dyNALml5UCH+KFB1oAyi
z/NRWfWTASFLbvo5iHKcovbfl/i+ouamHDlRZGiU1idjuXxG31zbHEygFQvjSqqQoYmuAgbIlG8S
zDtiAkwQS9i8FvQSu305blTJYzlcqAGy9M9SK+DIMDGgTmctNTr3ybONRcx1tQlQbUOGTMelCCsy
C2aUO6u90TJY0eT5kuxOcDcER5lqHBMWiOQjKHWogNUBAX+rx+hmA10pBWUgDwxUiRGFj8LhP4y7
6OxXshcRfVkmlNc/Gg/X3KMXDdHqcLD8nM50EmrENUp8zs1+v0v+KhC8fZCavNlPSUOiIExPsRrv
ZfG7F3j0jUnlrmVVODPHNQnan9YmmUmAXRy3l9jc2Eudi/XNaEI5IO20XjqTxiW1ZxleF5BmuNX5
wtf7hP4/uTwhsK35O+tIFp2rxC1RVpZIPidp4TGEPtP/iTZppHr58yHqqgdiRB3SPP147kC6qLKW
pq/I9PgOw61ap4l//xS6cEOspUADqo8TwZ7DQo3EG2zA/3v3uSO9N7thBhXMgCSvJM915DRMyGIZ
NQNtfieUrDCBKZB/CLshRNrVfPOCpW3BLXWhykLFilAUTmIoi7p4kzQxCPICD41ZxtvjGCUpFgWs
gI0avE1QcW30eOCp0TcYXu98m29bNrl7ZA6aWYvEeCOuejESPsoKtS9yu36jpUdwzKD9w5zulFKc
4EtjiGj0mRhp5OGd1Zr4TrG28+Vjqv9aLqzaB8PbGT9G/RdBOSagxD+Ua9ruRBaN9f4o0XG/cbpv
S8VkyDkj62S/+sh8ydknJ9+6oGyvuXEcX7E00qNqLFoTz9T7HENe6afY7r3QCYQO+8JGOfGqlqcH
HG7BmNAcDKVqJDjnsBp0LbjAl4H6aCcphmMzvx4ujrT3yIynF28onnHMrzYXHz1UxUJ0yD5ZjIip
dnVflUNElrXwQ4IFfjjauc6BRTa040yFd+Zehoi8/nvxHXULdlLr/Q4BcR+BIiRDL6qg2ABGZ7H8
yw84fJBLSbFGg2OIyG2TDB2ryqZiyCQUyNpn335FX6pJsuggeXTHZsLtKI2X7kiQ4zA/05dRgpek
7XlmSfgzfsp0Jql5i+iefe6BVxA2qTJDTSc8HUo0970UjSF8IIFmq7C27yJlbErHnPlvIw/cXWGl
MxNTKDaTxQy+APvB1DBCYBd8v7Vgr35Yl4RhiX922Uai18W12pTmv9VmF2NJhls9a+4Gom4qLq7F
uTQMi9u45qLsoXKSv+6CphQwcBmOdJGwOdTvnuLE6bH/9FewCCVPSH/TK8m8s0j2Y8C3+osviwQi
PTlgqz2WGUHzp27tQJofAHFkyC1Hn5vJ9FtYqHT7awraGVKMlTievgMb0Iai9r9dO+R/LzRS//9z
Z48xvVpKtkiHJRC8nfyX5WXY4wdDy3JpigqKG9JKV2/7pE9pnP41ny6n/XJd3lv1uIU/MH+nu2cS
2qOT2t4Qq8BwpBb3RwZGyHholNBoiQfM7WYBySS5RRthrC5RSARQwn8nAxLKyhyun3y+5X5WnU1U
+2q9N4iTTuwT45Tg/rSQmDok05KQss4HHUo60NIxTxAE818oB7NCgDAdRooZDqKV4vPiRKj2SILV
hsuO423uxUlRnpaBbQDmN6o2xBxUF1aYA7ejwv5B38j3vKzpECQixAXCMGN0L8i6fhqv+iiz+Orj
I7FGk9lgTBa3UZVfN8Xh/18BLWCxBMkaii7i8VbLcenlVhBwXsp9PhzTKJLMnFJ2MZ4tzrxbsq/P
xZ9HgmiDyOn9k/w3o+E+A23iA5k63Q0fTJRPyh/IGBQpqhVF0ehS8Tf90x4PbCsjt0bNj+3Td8cv
YHAfP0pMFmB+DY+eNbsw8EgCnhU0nb+KrBH9xkJzsAPV8h9KGB7ZYFFtlqhooeQ8CsP2K0w21MX7
9vPqPDc2gKG7Zgm8AsKQXIORoOI1kDHqLz7NXIqIXglqfDLAnAu/pjonzHlcS6vUxH8J+iBR2d6/
eKc2Rhpcjp2h8OblO3TMop7POm8u4SoZmaMYeHNfG3XUUeATMRW5Up0YSXss3kSfv+Awkq2EdrIV
QUIa3tOyAzkvGXtQkcKBOucw/zo/soKukcQ4h0ihcCgH5mup49I7aZ6J1PURu/TZfZ1yCSKP1Bh6
WOlVll+nYUS74CTPtjIdXzc3/CQljsi/XFl095QfkfQgk9RppAd/VSaTiXimM/kto5m1u09WdAp2
1ZUfVl7N58Da7k2c5OjOsR4FlFpkxcVQf2WmdSbbWS9klKJLUvIuYIg+3Z9x+pIPDGCzkJYT4XCB
2SxOXEmkHztb7ILc4zR7bfF9WYH1A/ubMamOlPhhD720EVe64c7J+IZbAgzQ+XZuh0L/SiHkIl+V
5FLTe5B1xhJOnzpOtbAg4dfPCDOu++5FEBqUtVz+dAOxvW9n86dhhblmU6Bd33u7S4RcR168tK+j
5fDhvWrbZDj0sQ00mOMVc/UMgRPzJ1q93PK5G5VBxBfbZsUSabfNZ0IZnhY7ej5cEqsa/SEjJoST
HZ42SCLUwTTai9RQ0ErMyqPubsp5M+KTKapU75JooKLD3pYl/f6uV4PMoiM0nraRVMnZaNdyHmgo
hB7weA7vXBxBDCIv9O5rYpyjG9dupVmBNjW7DtQWolJ5+7wYIZp+0N5iuJRfkCY/O0CGvbivLEwE
pzV1DzkEEdyEOTy/B3OzErkn+2umI7BD9+bhtcrcJb9CU3M6JTNvd3NTcqyaMZJJWF6VuGTHJy8Q
mZ/yJS6yuZxQf6jyQ76ICrIGpe1e+p5tdyb0rM54xBRGGmKjWV1zWISWHVWiBGGOGb8jW96asSJX
7ASNabCEAMiFYk6Pu1WdGHQUUIkOx13pmvI8KmJHKbKgDAAfUg4Ki0sA3VyELEOdZwXmbw3jhUe1
pDnmCqlaqrKQQBmNVl4OWTgKYC5MOoYdZnukI+WeblH/SaIKZHcN9ANuPk7PLm2qYlBABBU65GSs
a4A6MpioT8Wk/+3jsIUgC92aN0dzyc18r02qZN0UTtRWDUx35/wXxG/ovr+qk39NDLeOE2a9DHnY
w2cWvxnfLZtRohfRPD4eFgxkIdKZttjWh0PPATzUa7t+fYLR3fa8EzOmZZ/dRHkHpJdwNGunLsiK
nGNl2aJx8UcFb4fiYyDH6iG+FLQR/2Vqoc//anXmMwCrpZuuhbfHbu5nd+Qz75HbDFt8C/Mr5giE
7ggNTQYnxaLJeh/9iasZ4yupT+ZgB2BklH6JJheRUtGW8pI1H1HvGEeTaYh/485NyUqWg8yl+RUU
LlQ0UM/X9XSyHVrClqd7EViyyali/qsAQisWTChQ+BTqDFC0uJR8LN7SWNSsuMhmGKKA4obXotIh
0TiVvCNIQVVNHnbR9P7qm0n2TxPJwMICpsLl0uefKKB775MF5MYxMhxK2OCKnlOL7z5QTNxXBnGt
ExQF4Ye/qWfgiaiInMHxjxZ9Y8nqtvRY0WfXRw/1tGGE5TaVtRjakfzSPoLh0CBNZ+GRmW0OXhKL
0EhKhe3nquRnfnUBKcNTF4WRoV156z+b9bRy9a95gtucAyI8PO05eT/KdMPAFTf/NHP2gV1Zmd4S
Yr2A4A5ukR7sAIYbNWvdkkFCPAo2N4U9RJ7rK6vT7pnzLr6+CJcUF/knARvqosibTfd8I6UiEL8q
uRi0Nv6MOvjlMUy7VjOrjsXTtYRDZE76Ll4hKKXSeNG9uUImzLFrIy1TKp7st3hQccz09Klbmw4F
I+jnmkfejVOTSQEM65X2Pc0xrkz4xTCXmjtz69N4gEA3weJ9Fcgm5FXXFrOjVCI+Ir88nH0VYI/B
+lP18UxgpCjf34iPa8u+e9HXH8HgSyopU9XkOwqoy/G568yHozDAphnNHn7XFofhWhlZ5Ve001kT
Ev+IYWaWj5Bhyb1+UPp0lbndDeDG9LSLGfs3zgUifWgFvFbq6EePJDCLsSgQe8FTFhfVEIynBwcw
dA+oLBLlhnYVBYrQeoWiRhg9YWhDnNbnCBxIyjRs1g4/lnldeeSyRAuvZIfGQ8MrIyhhkvblVS6d
CfbvbuWrEVK4JTT6pYd38GdjfdqF9Rkw5iH/EKrV71BSb3eawHZZC4FP3y7oKxCLysP9hRHZpYAQ
HkVUb2E8eIHVXoZjEjHz2hD8LNwLAm8FyKf1r6yPhDPvZFFJkZs1rUKPenRw27QhuVo4VesiaHhQ
1i+Ji1Hah4/damZ2aGEWiAkZ7/49wDDUGOsRe7/U2sFfVE8itTDJ34bWt9xBd+NxbOcR3L6wyxbL
1Kkm/pA+7R6Nl0+w3ApYUPcjIwZOcS1etP84Qktr+JG4yhPkcSkYyARKPX+trsOJWwpPO33yFlZQ
Z0yw5ZYxjRBf+5r20piB8TV2uUfiLACy+UlJPi6JL462k1CXaFZeGWLRTYMWJZlMu5/ced58wYrH
cXfhCgH4xEq8W3T+0W57YR/qQdq133rxvYsH9pb01RVmB8MS/CIX5LZTVT+K+Oodfe9mZu9W0RVA
AckCRXdcwpXyuDqjBdQ2jJTwIbwElR5pAZeXxE10HphRmT9fduJYpi5kmyLIUyZ8/rf/lzYNLUqh
MBQ8PRLOpxkDYoAA1q+mSBVUoiyK/NqSpENm4EwCJxVIMunJBFbeRdy/8JkvF1WYcW60pm51GHwE
LM38UYW28QK+zS92fAKyYyJpnLUfGIDge2pgYymcFDVKZ7lYGiUfg2YKApjhN7uumvqgel2bJiPU
szMmOAmvf2fMiYdBx4ows8s8a2THqDY9rQHa6YJrOozx8/YmbLe7v2z1xp5qZC37CWKazTDpGCcC
TVzvZn/ygpD2KqcdgTTF7ghprriJoq3hEnYFzC2BijoQmJLd6khsf2O8Is9tgMo2A6nuEJcmaWDr
cbyMuB28VCRcca9FNs56ijY9wWYwumdOvJBnCI9fkL7oJN/vCJ1BqreA4JXkokRd/4EakmTb8rHk
oJmXI/uZ2c3saC/pu7NhzLDIUIz5r9IACo5MHG91t+GbWuNHYYVYVQ1vYkR+2o21ujK5bTbI2QVk
n2cxMGIbKW+gRUvofWU+J3ke0rSL2BhLk1D0zhMn6Uv34AboxJxzRFDt94C0RKMdi5ICX3CdUJm+
WPMhf6fGo0VnU9tSEhOPI5c7w03iZlTY4VSE1vJn6Jr7COpECOytnWuH413+kTYSfDGmPo4Ccfnc
PA6Bnh6spU3j4xL+UooAyvLjBzNj64FT6sMP8bDuZBUdeNLFdyzHYDTVzogGv+8alNxuMq6LwRA+
eQu/WF/Bve9SdMqukbbIzpe5olvsQTFuP4DJgyWB3s5c6nqq8N11oCUiYvc97jXURt3bbxl7zm/Q
UI68PM75NsIaBwHLmXu5esP0UoCx6WbyLzEeWhS+RKX4E+FnGhltr++YgEvZvab1SU7ILdQvsbVx
hqLCuqSfuLo2smP0H03vrNlxK/eo3cSyeqnOfbgdqn2vB/OUjC1CuzQgbAlZ2zskVW7+3Xtk+wMz
iqJ2n+6p3kD0rpERKLSePmTeufWGX2qyYZ8V5UkaAdn8eLrS9mfe8lK4oP6+M4SVx1G5g1ejUcEU
69gTxbuUI8IftTwGgKi4rJRMw4dAe6WSzeZefThVjq3mu/kyu8MDEDqk+u0Y1bVkb9zRVUW/GEQH
whhW0TK7ZbgUxLkO2fZxma+Cak5Sp51tq/dGVueFYBIHJuyCS5RXh9lY4FIb9+nt6OQm7srBeoZp
up/23yxPPCn6Hnm++yP8D1VCkRW9tQxzD4Fopj2/JCxNlh001TMMjjLBUDp8TRr/I2mkkCaOWz36
wF+3SrA1+z9wxtz0grG2qRRzAVkS94ieLfgvF0MmdkjupjZQMW9JQKXXdfUKNFR9cct8YNdAq+49
1yJ1rbh2WSzkSlqEDf82Ru6cA4jN5ilUk4lsPcZBxpCKRDbyom+UZhiS/YAAVRZaB/sPez7JtCNC
H1WSyETJSWxpetBdQ+VGDe0oLIBHoW4jnbGvHQxsAzlrIT9XEuV3j7pEjrAAuBZceJpKt7ZHdpCD
PnAcSnRRDGDe4XQCNcO8NnOgEQ9CcJBmvM7jUYDgK+uKBbv5MLwlBAMED5/5TObOzMAAcUhqjRq9
7tqbcOLO/RtCQwjH9msxStnOHqAnMrpL161Wi+jd2dK6KYGL2+TzopBkxpsFjUEKDtrpmP9kQSsk
oJqw4ldys2K1jrDDOjd8b8TzuWWEx3zKzrA/kP/CRKL5PeNuwNpES1BA47/WZOcU6nJqNTTjR5bY
OtnWuPZtPAxHk6FNE6LUi56rYIsEq+5WMJkkhqCcj+9JZ6s1OM1au0weYOMqBr+FYwwsV0n0vYE8
a/LUOS2vVWV+3vQfYp3LkzHnQS/8DFr3M5crCeMG01IouoU8UK1yCGEA7PiKyjX02L/cI0XKTjJj
5x240MDR6LebN2QiINvWeIMySXj4EP+C4CygGtOTeSa+Tgg2SwNc+AdiYvs4WhnJKeZuuPqpTSVi
PvmSqKxiLqtxSce9Fvw1Ur5ACkzZ6x/Mh4h81R3aUQnrSfqA1YPfc3GOnTdHuyehrzhKnS+1pxFb
ykzkzBT93nxpGpgNCThXqsbLFZYBYFuwVtM7KRwyroqncYxJeF4HzoAFMYMcukEAEz2OX9oak2gs
2PvUSc/NxlKQCcCR2mdUASsAv+N9sAcnmmKRTjAquczjH/sQ7P09m/2b8YIWjzVKKdJYA6ZX0/bL
yqNGhwUH3gh+ZZmNo7qzTpFh5ft0zAS2Ao4b2L8VgfJnoJA9uU6flI7vgFfhA2wHs+rIkMSHF0F2
7Oy3Dj/8zzT1YgHLO6dHyJEsyMh0O3XJ4SrfBlO5CDIOM1M8iQXuYKdAi3wwrQcIx8BX+QSZ0eS9
s11nxb/AhlOyhTZm4a6aDuwhdM5RqlH4SbKN0ZixuQwYoE7Gg9gGvcYAJErfuQz4R/WEwdgSGuIZ
bmGwal653adjeUHv6snxQh9yyd4SdQgjzZwub55SZAa/c/C7DYGwqzGvweq+2vb60snUQrayegmb
ahQ35IErGtUVrrfryWCMOcCpasKBaAh5kDoiUpPJPgz9D8V1r0C4I758QgbHbWZn8ABX/T6AcWB0
y2r71JCmgcJBhsHUNMWCb6fkNhP1i68aHi/pCeK7mCjiazOkBX1XULGapKIoYzbG9ybEysb1pg2l
s0bDbWtfNZ37EcoBdXz2EBFshcsixRnFJYeC5/vioC26LFH1CpmeZSe3afg8nCP27EZ5Akt6OSFB
JSWlSIrpJeevssmKuNCYC9t0Z7/Az5/5KSZwUQ7n6l/jtPihtUcONeVtrk3NYdooWDcEf5QPWxTz
yZy8mj5E0lSIYxZK98Dd/J+8MQyaorv2qecUBgmLzI8B4/Qc1luI2oWGHlx/YZbow1VwS7PFbcWq
Kw2riqOugqPT5xjYfAKKWhEEKe4L/Bieaorm37m+LaNNDI97Dpp8ONNKWAwB/o1T9F2yYXpbrJpU
Kl6Z3QLNeReiwzC2HBnzu/In4+xGbahsUwEPswBOSvwk0m/kKAmIGbA4psTM7kudjp3ZIvJ7Iwsy
BxeJ6gBsdzN41m1O+re1vwLW3awJ93a/iqln7lk9PYDX4Gg0S+TY1XENbmKA+YojqYBF+oGy8A+K
GegOAi6ADjnyzy/kTEkgXGhG5f/eD+vPqahS/RVkzrAdC/sh28vJLnK6M+nfPvattUhEP3dHVmHI
BHs9cg4YRRgUVkQmt8xrC4TY9P3QjGuIBaVGoGFFp7+2kwXEXEiSCQtmQif7gnVJqSGcOsFsZ9oZ
aHOJ1GK6IKu00ipFGROJNHBEapNM77RIncJundzW+kBnDml2m1UaTDUNpNR9bpcSDkytyZU710l9
bgVMeNSRzZmrgHPcxEYPRdYPEqpA4Rm5c/E7P7Yn/UBBXWKJ6/f9wiKkYu7mnppF9IRYbQfm4s7N
Y1WoUTdQ98AEtKk4KmIX07Rtb84YH7pOvU3Hoo7ZobWuCUgKlucxtTDWr6nEGoU70El4z3RLWCKm
3EclUI7nLlYkrUi+Lv+ZWsdnHdXO6NdcMJstvqqTUbHn47srS7mq1Mb+7icX0omkDlYQ8HXUh5CI
u2sfH/WIvnyc4WNfyzmK+/rLuntCEZ/fygdUgJKXCCzU4ZLpRk+TyZ7UGDZdfVvF2t8rmArCihAu
2HUW7x2Gf4JeocBn2xAFKTRaBWOgG26mAiV6N+T9Zs1df6RGoM8YLP0A6YwNAtVHqvdlLwy1wLXa
hEeGj7XfJJH6pXqzmxMlZs+ma27KDX/frsIxmsdhKtWSEPGl6YYlq72dylUpGrZIlTu1wwGgey4d
abz2heat/SYQgpbB8aw//bEnqql6hJ2T+HWUAjxBDxc5yNMynHaIpcykAQ3Dz9rD9mvr/V95nAZK
drBsnx+LZkSVva7Hl+FPRM4hmoSAIhvsZieyOvNOxoiljS+Z6+2z31qgQk4+6VIMOqhki5njxTho
AESIOkk4A2pcI7TIwM6TUylZRiIlNW8qZBTEn4E677XGgDp/DzXf3hR5MMVr3BdSA1D1rcyMuqME
czUVVV9drKN5WNMwb9Yt03l5ohw3ffYnY2AXfNu6tiTlqfvUvtTAcskFvVZ8w/N+C5YHRGHpSKnd
gW5DyU48Bu5c1O3zqHAo0xYnhWxPjlYi5LT8omDrvfWgKMxROGjaTEhnr8dvEjV0Uo94XQej1dbv
84xVkJoGMkZHHkc22mdE7a0b8UTAaQ90EpHZwnR8LZsQpyLbrENz2pGP1fXoOhvDVSzLI5b7/18p
sXu26NEiO+AEOSt+asizYSTs5eOavQ2c8yCbNclNecQHSyVf2w/3uX1i44eCl8elIxiashnxRuti
xAD8TDGULqUgdjpQo0NxwXPBEXzrA5iguyIzb1Gu2WyfQbh3wtNSa8cFnpcQf01mmmo5LvpeCQLe
/P2nXBGB3ozX5pIwgShu623gZQHuY5v53XpPEg+rV5mL2Jw7L4AMzVVoortpyRauVjFbHyKQsa01
31MubC7yHzYygY6bRors/bqA15RbhS+Kn//wEr7mpApqCTdZyWsQOgXRqkhJDalEdW6RBoWMbz6/
UIjsXBLb3GYqd7ZPBqm+O+WR0DyW6MsTed9f9h2d3fJkKFxVPFVS0HjJ5fqxghbOmXFJ5Yj8gKF6
wcERcQHrYifnWOuR+lghpA0sk06KjzpQrPLsDcVPnCS+leoLwsdX7w0vq0kAWV45gwL2QfXJXcMW
3IHAeFnON6aj9NsjzS9xb0pLx3qo5Ugf7JND7fKgatHv+o3n9TWHrcU5OZX2SVG4pYxqJw3pmxMa
qvVDSzQKJQkBzTiOBEq/APl2pYiLxkvW+v4auKF62143pu2qB9G021kw0uYjv1AiB1vd3ArsSt/3
ifr665IugTxwEdyB1IV3GnTIKcr8qlL9SeqKvmev/zUGbVT/m40deI9zmLwnOvct4SYDifHdr2fl
bIjrqShIKdf+nW+3CHXarwLGon2YmAAF3cAmA4GyK/2pFyss17Wcn+Qhfm5NDygk3W0T4iEBF0b+
yKU4FYrN4ONfFVQebqAkKSi/Oc4CA2j3GpPKy4pkRcLSqJln0bKrYGsi6fWuYnlWHMYpDhBdXCBy
O90K3oc8A6ZtMZLzls3PQGIBQx3GyvXepZUAXZRDH8D4zlSzqZEpAKUy8hjqU98I6GTGvmWUp3KX
st3IygrUjgAlgUC+QQNXWR/rIXkC+PrMCi4OESquWL7yX3aTzALQ6otaWH/CYXfsWJXNYzcP2EX+
dcJMXeM+PDA4AY/17Px5PdxZ7U6jWKg2hk9cOF3G1qYKj1oWF00fjXfW3DA6LBU2YTEhxkVY00n1
YA0qZxjx+bHnLDkTgfiN26yEUfUQoEmixVLO7L4bY8cnWmOTXlP0oFg2NoNaMgfXhWTjtM0pSp8w
BuLb4RggDry7GTDrBNXHYZynbTNeOK49WPRmkhdzBAZql5k9G1KPGViZM5yO+QWTB5A2fvqJ9rB3
GIV6JMw45TW4m4JzmXysYtSrwVIK1WVec4gkpDI05RbA4h7TSsS/Umo1C/PGZ27eLtiFaG842h9w
wshAUFCOqyFQig0q0I3aWkqS1zK1Abx7SpLac5gx76H1lP3K4u3SutNrvJKOY4MDAyGsWDY/7ZR3
W8lQtPMJbKkKaz33J18wSKoEO5e1Wy5GFxM1kLD9h2JpDHNbfO5EBZ2Ufye0a9lmKo4uIjjX/9r9
8SDhbJR3aMgugBZilneB+SWVnVLU4seCMAy24D3QdtoOILWfQP5q8YkrEn58Lg9Vl37QDqxCZhwF
deu+7AJQXT/c3a7kcxx2QM2bdgXicWUaXC+hACHjhxa+oglJQRTOExtgEUCChxYUzHb/9RWJi/Vs
+au2w8THlwt81nBtijaNKGjsgpUZV/VwYJxNS9yvxpXCoJSnlqwR6f/fpAxjCRBCzmNtGXZDtPdA
42y83qBrfuChIMbcb++92abKq9Zo2v8ixsHG87c2AfZukQ5O1QaUEyAst9GxxGTdjZx4zNw9jbN9
4lX0/BhbCPzoYtq6eJtuXhWe4RYgJ0/c7kZ+/1rzCdfGVBsyeSXfT+BMvd7lBvC4hoVS2xWi8YyQ
YHE4W6zhLca7SQQ7wrbgJ/7bWd8T0OY0Yfzo47bSDAzk3HX/NsRgwxhx5Qmb7oHtOUAoqgfX7CsF
N/1HLm68bF1uNFBwaoM3uBoffPDWbRnGIfVeINT1OB506oNQMDKEOgrp9TsnQHeC2UCZtYkdHGvp
i2boutm9Jc/pbbePpml0L82MJrjazBOWeRvqnot9lHE84Xa+wt0tW5iu3q8Cyte1HxDQYYtDbh5F
DNdpTLzVpqRxSghhkx6Nsn0U0L/3qfXx/GSWqB7Vz6XPMW/wX5Bt+3ZHtNLnKSUHqd7MR8/mtXiU
Q5IWJnDyEKOVVrEV/fbkMPIVM7UArAoFEKUCenAHBkjlQG0lgyByH/i/NwnKI8thLWyaXQzriL9r
cvF1a3E42tbO6nMpODP+FswxW0zB4Er50a/QgTFvxkWM830W75g729eS6Duibxay8zB9CRAT+LAW
ZlKqfYz7mSGfEgDVXacP5b4Lj2wegWKOFI/cNg/eXW8Z41QftfaMqb/XP5I0NfANP7F2YbShTliS
TicqJHh002UQqLxfddHYr6zf/pjdYaezHkH4vYiOviDr3gbXWm0madVeFY4BzhuMNt0nYIH450ot
crx/hAVyfmNK7nYX0LhcOMuuC+/WjgwPpqRv0y4/RQ/wPncHJeZDf5qoA76B8ilxcKfK8BtqkfZp
OzLDhGxAvTUrrd0r+0vxFHp0xChQ0pP9lcWGyuPphQx7dJK/Pl2VnlXhPHvM3wpyRFYnGJrNL1cc
cBz0ktyUL0twup6fWoj38tDh4OFeZc+4J0RzCimYwH0WrMkZahWOBj0VQnMe1Q8FYCP+ST1zMVTk
vSYCrABrsZlJFKNPYeNYkcSGpJZnPWuQaKQYlXtirmfY7oXxBdWUkwBrBreqcXmzKv+0gibrSfVe
3XOt5jMe98Kn4/n7Rd4467gHpg4eYOynoa0OwyYC4L5ONBcdGRcsVxx1o56CLRuyOCAmzbcoEKBC
Akgk3wlyVBSFxMP8A+Hjk2HAG6HifHJ7UOn5weoXgbppIEcGgfxWeGk+KoVm95tNWJHsjnP4eBz9
Y5okvfxJTKXcNhjJ6AVARvvAGuIa+QeHRCo6kaX7Nm8dXCKYQFFpj1gBjw+ME9GMIRDpUtEPkcB4
gBgvi/eKNdCmMNY8rdSddFvSL3GB2rolCKCC7eKuy72VluMuBiVUaE4rR34FUtxC81HFArxjn6QL
BrCjnbnt32Fsx7meO0jsfC6AsFWBG0mquJNRDSoBus52LnoMJhGtNxA77xZqLogE39WUJhSpEGFS
P/K8j/laDKvQPlbJ0KAOSUxEciRlNtYBhKXRe+fE2+hqbxG0x4rWhjjOQ/o4UebajXlBrXwYx+02
WN2K8ooAfXlsb+R3TpDc/SnexaAgznL6nD7mpO7L+AcVAQakFKAGOQQ0RPDND9pxxlML+IqtHw/X
KcUUMStLvt/4dOH48O3ZpHbHwwbai7JbpYtlkHrCJrrb2dpltdhPs2VZzjElTtEV2iOoYAAqMzeQ
X63W3TIkzcMv2NlWihcvsdIClFv1ipXogaVF5HtLRfl60s5rApDB8diolqR7fkQpknCYFyyNgXea
dD3NZzXzyoKJ6O3mW9ARrvJdkrQTNFZKrZn36Be/1dKa0GStAIK1NJPc0SEb/Ux4qdtIFtKZFr/z
BUQzD/fIdBaciynxEPwX7WAn+N6Lh2dOFPlhmkuw6XGaQfvi3aJtN8zRT12I+iWEVe4tAoGkoQPd
hDrfEQoq2zAcDnOzPSdalEmVbq8e7LrPezzpOa1aYaI2ZQs7CnScID+c9ypjtG961KgZypg5wERd
cOVWfEmmPhNN1ugDzgd/ukd+h0FXMqlKh7AWTPGWOGxke4RI1POIwcXDzZK5dO4nlyVG+kI34exX
lU1CLTu1vA9an2jRW1sHahWU/Cf1dDeeAM9gL/NjqpudEQuB67zoNYkYMx/has8rt71LTIf7NJzo
6ufqNDvBGcdVX3qbfCaJjL9iVo9+tAwYZPAC7Gin+UKtW4MrcnQkNr6nw3eKV0AYI/AWcclxBOTL
JjrNbNQIMtZCJHDIu8gxvspCCigkFujwuWkhPnYhbmV7Dk+K3Z6p6VsnLU/of9T4XazJqGkPOkRd
W5g6IHKsLeKxsj6p827ekoqMOK0ndCthWzdkq2pI7KyNk4AKBwRPr3w/jRPIAb3Bb7JzRewWSt3A
NMT3s3g8A+7aSMwKrlS3JSqRT5zFmCSd+xom2SZsCcun0YQ+DSQy7HWOL01OlvmOnw0lb4zzGge0
M3dfKOqUGMCLI9iI6AX+LRK3X6qj+HnuW+xKXmZLqGCLs47L1Kv4YDOfhvGritGJpj723Wf8/440
ghLZ0pMqg2crG8d9z9vTpIK9B/ZlRPfPUB1qciZAjCuo3fambfyLsBsxA+GDclF2oxwjtOJlJwg7
Ppx92tCr/SXkdhOlgXey9wrqpRb5vu2po0Jc4SOkD/+fkeel5pfu6OQZzFIqD552cZ1vsghouayD
c95M/DiTnGrtJy7mTdqwUNXWS4AxO2ScDOKHa+49fnd//p1+LIVUxtYNyfgDscESksq1+ItPu3KQ
aRyzTohMHDZccr7ONKL14pAYnSYiYDj/mo1Pc5rR6tY2N1k4Dt8qe0IwVg2tZWL5RwzD6U2FmkdL
ryalFFoFF2M4VMZr0nrdWSiKiz3rDDQLnTEqJxnZuD/8TbVZJqgyevxtPbPn1UWc4xMdTDY6b+yY
kGaMh3YnFmJZZJ9MjN36QTMUpePrV5jacmBC281phZAmhkQUHucWdIwOdLi2zJfuJZslrElnPJWd
XvxdcAmY3g9Hm5egEyF7cToTmEbcd6yJZnqM8SHNdk83fsyzs8P79OpbDnV63dQlGDNSiZbB+Oj5
lQBBOA0n8T1IjOrgkmKDguILwK2HruURVCT7M6U67GjDSdgdk46o/yDq34CsGW2NUS3MBs6artIg
IP8WnfyB/hQiBFNGBZ66L1lj21Seda1nz5yOkKs3SlSPmbGFCGx/ENyfgbHO3nCGriFiKL6s3wTJ
p2/DO2QtG54dnqA5HqdyXDDtmghHs6NL67w6C5D2gCO1ePNSc++tpRtJNHVegiEI6pect9PGq/1N
trRXpCKQdzWQGi02TEANH1+vHtQ8cz5NY+MNTsDrhp0bTNf4IITnnMoGyZbjfSuwewmcZI9Kzsvx
8k+pu796azp3TKjcwsU7hsHZpoaAxNmhxkhKTKt/OLBzHdtk5bk3rOA/I3VzsrlF1GMoJXFobFvM
RaUwNMSjg63uGtTWBh2zcanR14hYcd4Y04oiWq7jsOV7FjHV6nJRMvrA07WJnJXJp9dDlqorn6jt
cQ4qK50qnGyvIdXH2AfujVIpdPxI6zj05W+/YfPGdY9l00QzC483oH7GSg8yAW+4J4DVsnLuihN3
hrlkCnByWUZ3o4vj84tcXgHFjDEHhaoc5vYi5w9izNXJpXKhwdjhzezPpg+7bnPypZyNd7R/pp8g
JxVRexItT5hM3PfSxNCSLAe0MF0fePpVTcYpFTCh2zsuTw34o0vPZjPg1lzJJ0pwBiGN28J8fgJm
0ceDJqj46U8N6XBKwGD/Jm6XsOhDjlYUSV2JKByUS4bqUbLLSVGLF7TV4ZFQF/2dTvM/NgEG4NhY
HPZMDUhrIiBLINGin2o3fSVFVeP+nv/V4xZHLbbJ6yYMNNkzunI8e6DnJcoX8c+gad/Z8CEM0S85
CMA4QASge0quwObA/Ny6pO6C8XC56hcI/PDe6WLKnxq9Ykx4NxA1ov1EzKSnKdiT8YqHZrEgk/od
CtK1abU5Dr+dDYH5/tKV9Waz+NwKlzMfPpixvOgCEPaZf0CjFiR9cQnoDXJXQstobqAZ+EgwqUFw
381McVdmd1JW3Sln5vKJVZ8uxSz3zNAlg6d2MmyI1PAiuV4rf5nlb2kxiIHkQ9/f2boFZHicCc/w
5w9Ca8CJa/nFBElJf24IK1acO85+GqK3qUorasrjGbVp/d35c5HNxlJLLT2hzctmiF9bLBSqOxW7
FET68dscTPc4mq5yPCIq0eIS+Ir21dZHNKxFWDqdr+gLlLaGWtnms3jRS6L1uU8uSPKKNR+Rp6Ln
lZD8FZNVPnVbTFgq/2faRmFHrKyVBD/TSMLyZsnDHVdWLoo/0NjmPrOiI2fMaa1Ft3uji4LheOje
In+QBwg9PcbxtmuBVhqd1Fv1sVdnjwS1k8fbQfJpfjK6LNMyJJdsXjiZJVOdwoNR8Hk9tGsMvJeW
ycS6D3y/3fr+EWXO7bC0YZAWhebayHyi5fodpC+juzGPlFLFLq8wwagUlRjUPf/351Y+RTtPEnUf
IaLMsEoPVvlNyuttQjh7j2tGhSc7AKEHcVWDAlahfJQvB90e11Zj/4wbe51NWQaIkEMmN4f0uaz8
x1/UEduaP5/9MFXQ1/Oy4gZtyzkf+Fp2QKjnwf3S9IVb2I3HCgvV8Z2Df4jjIiNuR9Wx8CvB3O/H
UbCge1RLV4mhqxMi7SUz1kWTb8z+Rn7YPu/gx9Je5sPt6swWZY/7wmFbJ6zTivJTBxaTSlewtpkL
Suw4sG3epkgjNPF+fHQ0nQDzog+DLEa5eL+yOiAPTNJ3gb3ERGaE6X4OfKQhYpdp2FnhLo6SOxo7
c8dCPNsRxXQszAN0QDc4MQ4+5ysmAp+C6bksqi1sSUicuGmVy10Fj8JzrnObX4fW2X8dNGr1R+5R
CXcbauxb4lrL2U0/L7XBjdmdeE9go1QINUmH7rhz5ZRnAAsEqADsBcHKWh2kChoxGpaguEtS6vjB
tO4HXPziKhrdNR8raRU/LDVM4h/3msskEAajRAqfG7FmtcBQ3zqpQx65d3bpORwAHcEtOsEFI1nP
JPtUr5bXS7Mb712Iw0pCpVDeGwixbaIv81hoI4OuAr0ra9C22cohxgTGB0OAh3Owf1k63w2usQOz
P4MfKdWCm4qFRj2zb/dB7BPYk72K1KM0Ud/OSDrjKr+N1N1ejVx54r08H0/5fK4YTD5E7xcKu/ws
JoZCvDGUQxAdhK61uMqguZVThVRU+SOSD0Xt7A8G9cll7hMTA10/9eK1HT6AJAJkf3qzCbxcmeY2
7Ts5Q532NMV/SFR8pu09CS0QNcXmsxChkTdBN5kGdB+8zPAb3BE6CNHBeqo7tMzeQspA76ELoAAR
qP8bMdWZ8h4chr4xWvbB9pTTBdElOul2In7UwuOpGDQ9zt+1Qg7nKv0hEnermFa7Z2RdfJ3h7Otk
4dC9D+536lbHHZAZ2YuAJnXRrL/GW5Ccqmdl0jjl6Am+PcZKOWTFRJgxjJzB/fYa+DZDI23A8qYK
PY9ScHBS5CBE0O2Ujl3RweEyTRMLffrvRybvkgIBYmM5VJl+8/OVf1LbcdXAyGlQfVIgz6orERUA
9sMhXaj2Rh2jZxVIxZUaFaDKa716z0Z1G1fy1POwBRKAHQMYBvv9MWL69xf6g+Mrd8ZB9IfGhZIa
AWkLq6y6MzGSkbzeRwFP0aTKQnov4Vjj2GOnOV9Ff0+js3pFTPxJIOGMXYgPlzz0W24HVw2hZrtg
b+aQ99X2SKXfbcMkD/M32pntER+bKvjoU7b+4jvZe677TfwutcPmwj3I9w3c65P6y5+X3iwg7HEE
Ulohtc6saS4xd7Cx/oBEKK+QadrIuYt2NtuHV1OS05aEgJqbhjaOo6IA8jDUzfgqDwcZy1sCFupP
qEUdFNvXRwfsrzlugKfv7rkXIaxpIp6JXSEPLv/cvDeGy1BMv68VtbNRy4hp7Nd+nKynv1BDHlvJ
M8TtG/m6WayOMUgnDfuR+AB+Teahww0H4SlsAoJG9bB+/G4RVZxvZEQF+79iJMDwqnyCgbSaWy6Q
TUQSbYaThsCzSGke5wlRF/EZM8m59y964ExnRIEIkwj2DwMb7dOpNzAmKlFZgxH5W7ce7VE6/z+3
S/jQKj6Du3WjbkaAiEjQaNNn7UdMuCGGDClXViW+SSXVa9OhwewMmSwCAhnKY6u19ZcPyTnD1+Cb
CQL8hqOBSyFInns52icP6EusrLl6t32+BC+ieqBEDNnLQlbjRfjz469YeoI6fgYwCY3Zt6T0VgqY
m03RSEQ6bVTZ3Ivs/L2K4rTYm9PPZs4MdgKx9HrYGX4CClt5bzU+7LgmRdRpnfyoiOwrtZw8Ozhy
iMV7G7YSqEZBAPun4d8+P1In6Jt9Xkri7NLulh09ZvNvE166PvEljWyY/6ryP6tbfgijlN8wUc4X
oGUK1M0rT7lLjV2v0TK8ceV/gUfOsfuTS7ixd2SLh7cNxa1tyI6o1Kq0vCnikb8i6aOodz3/SDgo
dFX0GlAnmv/g7OIzoBoozCOrlM8QCnkDQMhAsz3sG8hogIRpQp4UFFGb+zPVG1K4l6KtuyJ/2tTc
dsCyb/R7ZSlmL//Stfms3N6nlkg7qNTmmoyGh6vJYj/QgU/lfeX0D//1NpiPbEE6WE9l/ZEItrUK
flMgn50fUOQOOv0mG5/rGPI4MpCjArkgDurtmp01NJzGV5gkN3dBajIkl5L9tBHBYs6+iiXcj57l
UmvkThz34yu8JYy2ZrLmsZYDwWWFny3Ke3ME9QgBHKVr7j7S0ds899iql0B6676sYqoUjc54r/h9
oFENRJH9lRuoqQJmciEu6oEweMuJN3Xc94JnEx9EREIQ5gL71j887gsO3P/kvE0zcmcPlG+A2krf
7OOqqA5jtysHX8Br3/PGCRN24MfhPjw80vfmpt5u8mwZyQQg3P74D9XO/haXAEd9cDBRVvcn3LtR
0Teh5K0j51V9r00+cM2+0kNp/3QiAhyOWVSXu2kQ+A9LjLnfrqy6LG4xa3D++DXmZDaabY/lHchP
hyWFFkNzBKfSI+ttqm5ZqtYi0CAD439THRECQ+ecwGL54/ekFvCBtQ2V7dKuuohUEFPDBR37bR4I
Z5Fbou6GdwojSzxB9z2uVYP3Qm7J3HSSunwthedzSHEx9JuN7rkwqjVvm4/giAZoJKFiJspmcYqa
f9nEXrjtyYNyQQFgcf/B3X+8La9RIwwMrt5Hna4Gbf7uVzXnbKr516/cGVi2Egigw1iRjTfbs4yM
J56ztlvIHIPPBkFiZE0zdBr9eZVPx6xFtVqeojZP/5dWcr97T5VWlFmX5+x62o2Jg2vn83fWeuT/
AJ+2Zqy8tJQkZWPwyWE2PrLLG+PLndaOLcrUolI3D36DnDxTSKclhqYSe2Ofkxl6b6vQK2pb7ig1
yiVlZee5f1B8PC00jYtfZBhmdR9IAITAwO4Xg27FUpUsFMC9ZoXfYOz1iTmugLik1ETsKqqnRKlJ
96ZMx/aIhRO85kU/0rvexMdBCOWeq/3SjnRC0dLn39pLdBJJjWLQ+FWzhrPxspXh4EvxL7xyEMcz
aB0vAi82A1h2Tyo9ltXYGbRq7sSWJ+jbI46wxOsvHcwUY8jeFBEA5EkOyS6PfBJ+syHzfRmecNti
qwVlM5yp4XmkhoHcT7Cyyw5G9pss6uLFXqP3+yUP8m45O8Pe2PY1Fn1CzJ2xlusOLnHvx6kc1cph
oejZAbK+RRS8RAP5JEoZTuaHHc4153/Rx8LjTU9Eotnlpc8HSOOKtGkiv9yT4ISn7lkexlduvL6C
Nxxb6Yu3fJksGbxtVHbIMqPFvDnWHBqwilCDQS+pzA+Lwq6NaH+/wjJuGwZ7N6dzpZ2CIC6XLA2J
S6i4dIFPD4sOvHTougb0iTDAE8xw4UezEuxqnNjK2AynMwyTibyHShkcsxXEk9Re5OaMYMfRXswu
vVFgkNNXg5I+bjfl3MYv+6AZ6r4Ji61d5uNnnsBD0fnlvGGSplB7umORrBkz5quQbHyLO2jm1Bij
wJ+PcjPttW+KTpJHsDOCbHlTdKty9WOlDdm/QwT4GN8diCGPkvwyNeB4H0+8IlrC6dk2x0A3dj5o
QUmvb60wSsHVRcM9jDd9TFNzTvEWEh8/0eVW1JgfWaUcoeaXoFkazkF/pZ81EeQ7kzalK/dUrd3u
0l6yGHGe9xtXbPlBt79CgEXrvVcipqHAHPgKSaU1pt6RPg7XBJaKdve82hcLeVeJ4p3C4DrT+gMj
VeM1abNB5YuGU7d3fZ/7xATCf29INnRtUVDQ/pN457iD9dhGyXX83NhFugWCRM3ZArHTeW9AiSdk
3oPEgXML8WCaXzrExxYCoJQSNI4n8zYEVfKksn9WxIik3xtpzSUaje+rH2JzR85qXeMAKr++qmAA
aDqMtREf69YdRwE2xOmohMwcP6hdGCPLhv2/t9lp11c8C7ukeDn9jLiYAlmu8eELx8OfxsxshgB6
ND0qBGX3hk7kxsJmvH3KwguzEU8UxyJMtt6OoWnRjYMOAueNUST9m8X38WTrZWSneC2VsT0iB2T6
tnc3mjfZVFFS1sCZDREC5jiUto10b45dr6Ux9BA2Gka5G/XvuRExC9z3nvvcLA5sP2NjnuSIpm0P
cHdrOh8kLaaB9IYTCgnixFrH6McqLVP4Yo+K/e9LgdzqljlcZElsabhptO8Ef8WZF4CNFWmRmOqs
PL6f1ME/roJUjjICdGDkzRrulomo1649Gszweng4iVN2U2gEWfYjCg9tsQWmXSw7s5UWqt3vAGmn
iJK0lVpS9yMGiMF8/s/H7JpM7J+qX+bO5QeTglOc/UsLJIjbWqUvB3HJVGchidbnyQGykXUAqtGA
zuBBRWKE8vKiFffF5b6heH9cKcL4yr5zjPPDMsA36weKSbK60Btccg+nTmablYvF7O7SmywMzsU4
EeE4gQOgo44a8EVJKiMbp0q4u1H9FpZAkqa3ppj07kEMS+YlImSxDYmQQ4F/QqvLVnCQ2DbWiREQ
C8dp5y8OwDYMxGFKfKoG7RS7USBFhS9ML7Ni2Pa93pI7tkC6ui/DO7/uYCWW3Nebq/1o4mCY8awg
d9cffnsarmi76e5jtkyx6TKRqLY3P1JAGKqboOFc9gm9AVlEkMbvFcTWfv3rZ6V1RG48i5bp0M7i
HZqZMctF7Qj2GaASVeE9ViL6LDIec/r2zxZiXOsW1Da6p2tLgBI3NsC/B0RrIWCL5BRGWEFbtJ48
tObiGaYp2JjZw8MlJ0f6TaN3L/x2DA6l0kM/zGDcRqkbWh1ydS0qvnLZgKTZ+6N8U3W3ebDmr1yJ
kCOETMM5rdeIHn4QjCzMNXNjsShUDRo9eAho8EQ7RXyo3Anh5h8FMafSU1tPl3032kQdzupnnXcs
WQI1vyR4EUNqlIVG8awZuX3Q6+OY9r1Q8vRtOYMUY8PvEuP4bpus5BhbN5Xu/KpIM3beRErJO1e8
6nSx6M4mAnBoEwnbnr7tvX371fyRldXRsu5MwRr5sFgUSfNEDq515yv+NRYPcV3ndbR4WkwXOqU0
PLSq4wWwOn99VU02KTxLUd/lc7JTvwYaEkPk+8IgL2ND07BqicMmg3ShqdyWZ/UFGRk+Gv1o0FdJ
W4U7K6lChzEz7DuNuz9QEeAOGKUKQLXXS+W0Y0vOI3Pp7LGMwZyvto0uFZBPSJnd2ABbpF7vmUUi
7K36My4RJ0vFDwbw38c4VYZwferQ+U93mmTnmx3swpArQI7/0u8xTMq2Pm2AZALDW5CWSQbhrTlR
TZDJBJZq/cfnZuVaMuk7X5A0pJJ1lpcCVmIJ8oj1cUnNZaxbITjDpWirq6qgUR4q2f/XcSZPe3Iy
rFC0n44ziJ8Pih/XeBw5fxOqcrIZT1u10n9Ni/ARuouPIYnRU9az1ha7EXShwdY000XrAQ9R32ZV
bPvUbxVOqDL5QPdTUln88GUw5WW5FnAp2nHuQlx+C8e8Irz9hVJ4W1gXzuT+hl0oXMEqVHgJApXe
XcmicArkcBLyRHkf7e9FHx/gxbNGtYfe0OJexnorP5YFJL9rkttlx89W8ypElAhyuN2j70eXnrrU
8iY/9neS0OMZvXnkg0/G4ZvdjYqGp7BIEBoQRgB2gETs5s/Fw74G55A42GYiyYjii7XCq6vfD+GB
ICkbJuasLuQCCjHyY6Ld/nHLfUqD2fPeIMxLGwqQ+8MBzKOIaAHIZCefL40mzP0fK+hWzdEU3v0w
nD+sI3/l5uym/wOuyfHlFITq42OKdype7WunLhIo7oHtFh/J4bwoCEoDEdeZ1sqUJJZBn0hhHvHn
uFxdhkdaAeKavH3xiF1zJAbZwd+E1RzUv3rovFkQEj3dLeNSUEzIx0P2HTP+FIDT58OAfM6aZ+Ar
QUq/8NEVPp7LCrz3GjynCsDOu3Xx8amjxFp9mg2dzgVXXGLLzz3Covnlzbehzb9NWHqmTwrSUBsF
emRc0jck4f+AJ+BrdDWSxnnPR2gMsdWQCZ0vW6DVsH/wwORoUbddMp/gOCae684FvS4lVX0vtmhK
ngvwZRYL1Bleol+CR9MPJpoxYp7QmszCIJDPG+cEh5arEOACiCsiKEFoQlMMz3EeC9ql6ocn8FUD
G9R5InoaNGEJLWOflkrNwQMkVKjQB1CCnVbNmQ8PaE6VynFleiKuAXmniOZByFIgHjw84f2d+kD3
oZcKqz2lIKVO7IyeUSnkDgB5hLpu2iJKh0LvFa4HtAWp0p3qPtkFhjt1kPY28EKhIx3HjX+lFgQn
jgEEZrNsD+jHYPmZMMxpzEinjcv1pIlD89unA1D/VJxqyBUdA6KQ4Z8YbkLmp2+JLPW5lcH81YE1
t50CKe4OGkqDgCSM+McePza2O4SjsLRM/6bmS+MmATvOJfhxgXPevL6F/o5wPmCkyxuXh2/tvn3+
I589gTmQ0VFr/DqVn3ln6i7EVBV1SdIeDS0kHy+Wkk6wYukywGFdYgsdBz0zF7pAwCmcfunU2vXe
rVzYtrB3OaLxlPzdWIySiP7ZcMAjM4GZmti1lyOYt4vAs63RuMbcHJpqoE9U/WrEHQuFAli1T9hY
HJSLWpWsSPMeFcUU9eJUnjahv5ocQOlTRgD/Bn3z9MlquRbF871Xn1mvnlv1jJNbFDBPHBpwrEPX
N3ouvTae7eoFDofvb7PBxC4CaFojX1/aJ1JQPHmXH8s50J1hvSMUC8hX1kxEjzhb7sIU5kE5Hh6Q
x+SZVGSLLFC5Q4QVkDNxd9ygoYmU79MO2/bwcgwexu3/lSGoFi5qIbMMpauam/LJnW+NbROAIr6v
0lN2OFvmJqvEr8gtEFx+y7mDgnAJaxjnsvg6qTERVXUNaKYQyLC/CX3OEn7wi+054DdQiUbSHwEl
HReWPkPp4hGQx/ryQdtEYoxE/2zkbSE2nfoD27618HC8jsUokmJQ11aRFu5JWgg1Cq1M5NUjfSE1
ZnCD+MM5kAk0MJj+lxogm3XcJDB1G7Gkt/oklo3hvIyMAo05DACEIx2+kouXeRHtjYF1IvFqoJ5X
l8DMitWkEJ+q1TLyfVsGMZ5Neb875cH8atkMWKw1IvPFDdYIITwJy9dX7O5e10vHNXJ00aD4GyiU
HfKrwsZYGl2yTWr0vzQUfJTv3AE797Fz7Wg7Tgx3PvBXUj/HdQQ/ozWLOfbFg4e1P90gWB4wbXem
re6CoZHwgNqMf66rWNPrN6XmMK/ZLglh/RR0hE/vsrW6le5UjZzRL7Txg7pVRVoamJ7914bi5eTE
X7Yhq2NnWn8HKHO2OczEJXOT2mp+yWgNwVrAv7samZEd
`protect end_protected

