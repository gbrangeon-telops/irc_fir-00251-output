

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
RZm5UrZFV7JOtGxR4Pzih7NQYLp7LmPE59R/6o+hZN+ZT+nCA+l5YH+/j+E+cmHHWo6IUrn/ULaG
ZkaGINks7Q==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
MRNQzUt4f7a/v9KMrin25EUCYvWi/twJzLlDdceTmDN2GCvOURSU7hHpsmsqqCb1xCeaV7xbvs0c
MXpZkAPeQc5Coi1irNf+9eKbc5uIh03B/PevhS9S+La97Aj9rjHplzcZDEBFN6fiyAdKvJgOrOyz
87nOO0u5LoaEOeyC6ao=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
L17wVQWzSUChaUkUbjAqDK1dFxRQ9orAmYas8htY5fjqeIDtBkS/PldQL1EGRGrFVbxZVbStDyiq
iWMlaMSfJiAW0codwFWqGkqnH6YMctbqpTZdQPbprA8qa73Xmy9S5tgWXo6y3vZys5HBTFHxXMXj
HSJZBGLfj5+GGMkAkDYYBZrgDs/jxx605zYzRg+wKonRxjx8C7c4r2cekqFXXjEfMC6t47HLGKZO
Wp8oqSV+SdxjNfsxTeAcFxqhiABG1hbduxwcNIQO/0mgU7awDWqjimqvnE1+KO7vQU/MVpl+J+Y9
bwvxkUUMkYnqQG/HGWvvQ7Zp0u8+rRyDh2dzOg==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
yJG5RZbV6QsAW4khC+YjJnbI2jNRxPOtee58pTXfgJVvj12BYVsRuhi1xiVJgak8Vy8V0UJ43Wc3
ydXie//gOHZIACOddgGz8WdlyWauaZ9sd1K4GlV+vX4K5HkoOyunq5QSLYwU2X/ZYYkTAGg7My6m
h1UvByaO98o6pNd+n1w=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
QjcZeibYm0SAHW7YliT2StC14hkmhpmI1+m8klXbQfAK/yXQ8NfNnDZicIHqHpAbgVQzoGSkcmXa
qhjmF7JhXI4I11rujpUqz61fAf/3PeUiYimqp9l0xnePLlrRBeItzqfetftMnQ8hBAuI+sARuLin
j4+kHDvo2V/A6kndknmKA6lyd7gI8Mgzy1xgvua2Bfq25TZ30r76kaSXXo5N6hFVjtfwPGqnYepq
02yTg3lN97x/f3REjUh0T05iK9mOISMgvqQkxFwl6hBnLhp8WW0zJBjFvAguLZDf4CMBuYBnnmGQ
axcOzl5DWDcYTgPm/DTciq3eoilijus/JUHuFA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 8000)
`protect data_block
rvj7Bq4AP3BjmTc8vzQiAU61nsxzJoQAior5I5Bq6tsbBDAzpzMjjtM0vh57seNNcGWmkLcWL2/Y
mB1WsXnruMzwkm5YPs+a91voqUUrP5X5j2ccsw6wxDbJEWUPrNJ4lAQiQXWkl68g/TWPZUngBlct
YKn4b8es467SyPtvM93MdTenRGVEhEgKsjtfE6nFSPYIoQkwmaE6JNdkK8IP1ptyHuWKe1iLg8UW
j0xEdfKU/v79uEBsctOSpGJ8eGn+0kkCs2poA4f6tj6nbuwxvl2+apNdo6SI3zk2Uk6zWBJck1Ny
fDs6+nm6+x4Cru3RJ8cyIwjhGt8+PLa3iCDqJ669jMErk23mCWc2wLZTa7OhOblzCoRbJ5pGROAn
Fl+UyquTvnMB+YxR6KaBsw6SsoQgKVH0IswmoF1Bl5wAAOEYBmlxUl6QjR2i0XhbRY1EPdP0dOKc
2w3bjh6Z8PJtpG0KNq1gCHVyaoVDhhS8hh/VvU74BvbjngunG1ToU5zu94ozkkNLqB7tyimUFAsT
8K+lWCO8CPIbj3UxCmCvRFoaRZyIDcpHBux6g6/ho9dtLMov0bUs+9eAT8IMHCjpiFX7+wUWYBio
VVh//c2WozXEerMXRZr5xjUTP+7VLau41JDK0/niXBeBqjkLs9ytXxFFN0BCQoczK+OMzq2/aYH1
3AIL+OFZlHABfo4FptzHMPFJkZciXIQvjFdATGmEdZAxJv8PuwnMnETH2QMb5TUYNjuRjmVJGAQX
3XGNllmcllAsmVjTX3yCLm+X+mAWdUsTCyBkY/4S98x352FNzEo4mvpAePMEvgS0ua6dcwFpVxZo
atWAmuZ+fZDLeJfvSF9w+1RpY69G8tzq7kaeWHAPKbeNp6aEk44ubZNQZ/n37lIl6idKFdqoZ48b
lI9Rj5gE+kiOe0i6R1BGt7d03S+5+3tztB0DUXx8M63ynWROWDcrOucJ1tA2vXQLfOoxOKbdRYuJ
DSMOxYPEV6mNR4o67ZcsCyfvtNSY2XJmaIF/4fwNJBBIB5KuZAto62X9TR59LyGvZIsn17I09o8x
6wpDZ+KhKEeyJonEo/Ac68qW2NeTKQobwvnIjyaWXCDJG9G6SymlNgt7RXsPfhhvAGF7tOpEd3F8
t7B2oIx26ziIyL+xh7RzBlWDqPKKzhap5gIdNMTfpjsaItw3sKh0sN/a3uFv5RAjp9KniAYAE0Qy
BJxMjCop+rQqlncRa1+HvzJCuBhFSBnQdj+hC3JLni51sz57PjYAQ5aYDcgJk3KyqtwWmFFQDUPC
FNnVZ15K51K3f/aczbzMC4vOmJ2ofIAFohT3ieu+dMkj2Ge17aBPb9Q0ESfGMhA6BjDvGz2NeHaE
w1kN8wXyH+E1kzhFEMcmvC44Vk1aJwbloY9yX7s/ZRfjPMEkHLrcxObkrZXfFE7xVtP1u4LwGFJL
13vxzl6FdJ46dzvV3rHOAFWJQi1O3HzqDI1ZL+UNmItlXaKWKY6ypTHeEeaB4ZccOQ6nyqJpuc/i
k2oHhu/6g4uafa/d3ShPQjsXOd24XVj24UH5ZMvKn5MtCK1g48pj7Cg3OLdtKitKnos0JqauDMCh
5yhBXskU+3l0hmWcHFweDVs9UvU9r3LJpWq84QCb0rR16Hol5hBomPSyIpB4ObJy/SHf2xRaGoGb
HL6rCaoU51RI2ugz4aHRFJC0GMwbLRusfy4BWQEjmfhcwamQn9yr5doIZ4j4j/41Ryjj0Jjd+D9M
TTM386cP5dtourrrbFPPNq3gW/dAQcMhiK4lBIaRIFR4bee6CZDx5xqG/k0OP5+35gLonLa3HscR
faFWtENpYbHg70c76k+9Jqrw4hRiK+An0iIbVKJ9Ksvh+ocj/ksUodFCxAarbsPBuHYzf8Z114vz
Y5AJb/sUQTqGbZ5uswmBBk01YcLxnmb54QI0TSECFwsrNQPgpyxepRYPiV3OW0ZXgj9YWfqZ6UZh
zRpE5FmEKk4cWpkEgaiKel7w8/qM8sorN2Y/FQGVDaQ9XTfAB790k0iTDNuCssGgNeB+xMtA+guB
kiqWMrgi37RoBVzm05sPnhsKm64+K66ew+8+cKPxhbW5I0Fxy0glStAuGsnCD/xC6tOY5FJlNmmR
hcqQDLPAY7pfweoSKLgxa1TZWEnwr4cylPsChEGasjBWSArPmlVb0hfvBxZpw6HiZUos2wOdLXqZ
VVDC22GCSQx7mdJU86Eurj5xjfwLKqvi26KirRw+hXkVGNiBlOIaAQuhWSOxYYUXXMp8Z206Wm12
TIAbBnC8fbx3R4twKfyqjvWVFM6qk+gd3NTTQd18QaEKcWlkz2dFm/lfzUpLDNvZoVUY2H7TnNJr
zalUs2w8l0HlNwXzlOvV06uOA61+Z+TEeY3naXcOnCeG5MnMO87Vkp/cOUTtMYqlsWug9PQZDjQj
Z3rXkhts8wdAapkIXgvF0VDaskCZjXh22H9KNlaB+RZ836v8tJ8khd7tqLCpfL5ddwkaz4Ofn+0k
0PqxAPJy8/sBvpNIsf0/+0XBRG8l7e62//8yMNi4dX98aG8UF3Pt+OudVIUM6cISMvXkHzbhwcU+
F3FAdXlvjdm5sD/UF9eK5jF9qk8uxmRUUsThmS7IytEAUAH/ZPS5M62bA+snQO/b3U3M3C3i/yop
2ICjqFrecUVEJyIWH8CuWWCQMX5cvBsoZWqzEx3uap3oC8XXtqexCscqioux+2fTFWziEabiXwwd
a+Xa0jHQNXu6vJ8o/kUzaCFJtn77CEFh67CIQLQyvDFztpsKbelLBd9Iyed6o0NirpUoEd5VyGpV
YeZ3pOt5gW8zvtJJGuxRWUvenGxcVFeLv95FF9xB4JAm3IdEaII14tWawPmo7ek39gGxSvje4jXE
WLdmQLXb3yCc/KejD9SDX/J5yO9lrNF4F7/uSc5lPSZ/QuS9TWhnjNjMCXdMcGvmuUW108k/T/1i
hO1i4V9kPE67ylEYu97fSn5sdM1FpmPaKJ1EK13cTGRsLw1G2h4pH+VoAU4hkz/C5NNiFeqMLZQv
tCVSbtfduBPDUzfxVWL0OxmNePAJMfo+VubEiXrx8L1yBjEuaVFyYH8/vgtASrr0iTYsdSKUeOEW
o+mxF+K98r3r/ebNCKW6fyFvQnp0VImi6vxv9aZ4jVhONORM75/F5Do46azojtjzYKiyTzrq3br/
m18Me4e3qcInlEVIPuwdMEQGGy0/071UguJo/7sKDgsyapN0DDJnfjcJGvEnc7cZeVBp4VvgZQXe
eqefH/A8zHJCMunQ/y1G7d1ickyf9+fEnR68H58vg7ee/mTq212IkZ3VPCDRYBUolaiQpFMJ6wom
pDxJYmr68Jw6pqD1Cn0GYxndhhMKBnO/WuuKS23yUOnG9YL8t9twKyF1kp8WEnn+p0AvF9WNnMZ+
yRMrfAUR9X/vocMOH9iSRJWm8l4hzePWzwRhphkQDpHsRWFQlN4pI3xMvY5j5vCXz6R/NCkBG724
gM+Mkn/QgYgRKCyCqHMJMoW7F0HQbl7Cb1wosA5WDox/UhsGs2FGCRxzvXUDrk3PdAaTQ5QrhcWC
6g++aNU8C8BOBsm+Tf+8KKMpPg5/nEfR+geLVlrKxiitc2gFrwADCLEo0kvFlslZ3Ey8rG1ME+96
QtV5uP+kfuVlmczy4ffBTVs0bPg9CadeMIgBzBFJV457k/JtXsvQxAQwrE4CeCAv02Pmi/YLpwGk
Ds5AbFhS5fcEvhHb/OjGX5MmNYSvZ+ZMkkQShoeD4ldzF/8e0YQqLHdqgAFauRcjrEMASot4qG0b
6Yg24x2Mtf8tm1CKatTrP9cA24amzWQw0jBo9GUWeM8GoZyGZndqyDwI9odkAOsvZOOnUInDhco0
4UYHJkLKJJpvYGoVB/q7UBLwKoYoVcJNRxI8SJEpS0geYspE+d+l3c8fU7BzXpnQv0qbYau/6JFn
VzZbW8qeGDaZRta4T0sFm3rDDdE/YiwidzbmyV2ELb5wiNExF9f+vLlHsbXQ7IYmkDZpSYw/OSrI
8wYLRjH+mbDJVmD3lgXtlecXhaMcUmxqjbNUcHXVY4hAzm+e6SjnRwgFRojqvpOClfGivBJxIM2O
513Mk6hyjrxr+LwiF54B7UfbOHh64oz4IfAShW5HZWAn5hmKSGrwpPlDV3J37ar0QdHIriXjRaWs
s2mWcLpFtuNO0FmoRUAUNcnNTEuU92wYDefvp0bpgPd3d2jANpoAyjz5+mHxZQShnGBm79hZfD8c
NtfnNXg5Atok6w4VAaNlQBxI1WEPtMvhnBgIHWt8zcW6sdDCN3pwyKqj8bSE7Umv0tzxIvQQTyDa
kBxq7QPJYYvU5KbwJwXfBD7aZ6ge7gNFbaMyEJdIVtldT1RGEJa4MGSUwLlNBIGrexCwKnZ5VHbP
jz13j6fWrljxrHwfQMoqT8qnwzANfX/3B9e5LqeUOZxLDKeQTRlq8tr10VFleqt4I7XTYDEsPktd
g5uTN5ranREgH51TSeLsuwCNPKmoEre6Ed7qKnKZoIi+m/LG6kX4uxnpfwTvRblq2Y5MrIeehPpp
vGsFQcW8bnwdYQcAuicV6b11AdVsvHElUmRup0GmQOWZi1zzvaHRkyiPzo9AEE3Rd+BI6dqqXek1
9ltbrik+VWoU3uzRRlIzQbmppkfKUZmsHTK8mHzgSFj2kTEeWfoT69XaKUceh3X0Rso4u3y0d+E6
vC3bOsgS/O8bJfb+r3ZbfDE4fyfJBI1DTz771ykpLbA74CWvf5p0Vh0Tt1cmbKu3Ivggj/8OT+gn
w2dV6FKkaFd93AYQH37QzejAgNORlLP6NKt2ri8Oc8LsOqsAYCKA52NEMMfoTvOwGbMbvchTDhq5
sQCqx/Vgwu/VX/Iy3tJAuYHkjt1teHHLrxU73R3ZS+ITzkpDb9V2kEd58hhwlhUao92iNYpL2M9g
UJbE/ALVK5BrTgYFphmhv0DAnMM83buZkmeNHL6gHJ/b7qC0A94SNDWc2PNMvZ4UtHhXp4HEZauJ
VpeCykxnwQGHfwdKszP3Cm9vYfbeBHRduyXRnO6SFmjTToWUJP6msq9y8DiUn3FpJVTkdO/w5nJ0
FUNPf9TLQ2zCX38VLbAQcpyDW7MXnENIqURcJXlNp45qmna5srHdqCXEbTB3nQcovoRzd3xnjDBA
X0MrYzktI0n6AjWLZwW2u+pq9OgMvePCF6lIO9dBLx5sgrHLZcacVWfq42rg4YcPUPFNQrhz0yfF
meCryw+pw+AafHcZyX1FLRlclRJxRRrGVrr9Bj0utBHSXCETYbvPWEadDGdFYDXWrrlYfl2VIrM3
R1KmXaaAyyqT38oW4JZyAIuU1DOks0UvsZ2gcQWSU5c5CrzbGcsa3vDckuDVOLkzm3KRb4PTFj60
/wUwFhLrrMQvMumthRaFNj4CFD2AtBFZO+xTDoGjsfVTJz1jPeLTPeUfm5MA+R2Xkjb0uYc4NF+q
ZAgCTuz4b7Sza5MbSnobGX3jBUTebGOyVrbK5zQv1/3DzcWSLbmSGKj6Zj3NAnFsNywdAmeI2PSU
//kN1V45JOtROoPDToR8TGm9vjX4ujFsObtwPXi3N28b9QeuVyAwl9z9giZkmw1U8MwRxPp22Vej
vCMAT23ik1wNAnjOckjhLYPGXkte95x8RPLbBRQdT1yveQDDO+rqe1cDUQcHtyMjS6w7vxQKM5eA
8cp/Vko91ENHvH9l/lisnD1w0vShlU0EsTNz76iemcyYU5szKQbgV3mcHGFG6ojV/QTblrGx9kE2
mCDhZMjpOTeze8hzZr8HETWeW5imT1BMzi2DruVo1/GbFouJsIXv/iMtPXPEMOX8LMrEqfqMRn4u
Py+1ksbnHoaVkQ3qli0nGtMJ/vDTj4yhJtm63B7bfh31vXD7NObHohWcWcjGg+/8T18hhjjA37S1
+3Dy1kAd1fsDGdWmtJJOIQzyxXSeaHr6CzWjmJ3Pa7z8OU2FKqMsZeCH+FjzyOZAl8gGhDY2w9LD
ZxXQdL3RMn4e6bG/cK/LdfvvZQMjVvSl7aN1VLa7kwXnOpvUUVURf6BHMCujI7Tgpok6oNLPZs2E
+2XBk/6bhNfbAsmU9VIIkXiCmQnm1BRLIqH9+gby28TIK3DcNKALp8GOvZ1xlykOsDeRA0DQKgX4
t+zMlzhmvdNg1WX7shTXZIwpMN4Afx54QFeF6MlzDBOpa1t+BTER6opGIr0cxd5NvYsHIgnP7t+i
XoorX5Oa57Sn1U8yo4Mcyf//UuFO1o5bCslty9mLX9GtfK4UdkKqyTuTXR41idcKK3xy5/LGQIf4
dLOHogHFEUCG2NddcA27TY/2YDizpIKJpd8aEcyibxyxM81ynrFqgikERtzC+UwePI7oxdEcGHDk
xFFBFt6pt056mJK1fU5y91cvDZnoWhda2H5Dr5R5Zc2R83+Onk7Wj9OdRJMtiuwuL5XFjJoGKryG
aPNRu5PVHjXYg20luEIefLTEV44dL6VniQyMn3V7Yg4j9kDFyrD4D7T8ZPIdF/VuQwhnVlFtjG4P
ysWE8MZo3YjN7wTbvuw25gpj9Y752viCm8uyDt0rZZMjjmf0MPWSPMGtDz+lUQljc60E+7DkxyaW
bWmfrr6FEZ7EDYeqqScpk16k6cq1UNuDPLiTlLqbwC2ZBwcTvI+b5Vvg1+ZBXSBKPSC/h0H7+BTl
pAnnyzr9mWNL7bG7xtEC2cmuvn6un6cEloVV3v1zELA707sGlTGoKgvAVGONSCE0awapMz22oi/z
g9w4Ga/2f6zwHtye3c+NBVA+t9qtOvC5BxDtLUrCh77R4H8PDxUMHtVrw5NSXGcG4qbvXEz2wShn
F5C+qvzM8SEyfy3ztzsCJ9NQ1HWd3QfmcpfXSlD71vfaKFY6J4xqaCVDUng1dxiew5yWNfrIsOYK
7mQK34PqGZ1JATBqdUOqbCuHLz3op4ZWzrl9jVaUV/v3riNJzafBezBuJcaJZ2/9tDLvYi9N575Z
t+/oe0s0qYaLBbjUc9eX45cz8LLhJ0eqXVxslHqs3HviePaAAJsHg4ja08NvHbvlKoVQkWaaILcj
sXQRnbWNEwZn72GUj/VuR/k9v8g+mazNYasyjba5XJaXVNP2M1VtoNCRaJ4yGnYJEKJo/mPg2omc
s7tXZl7eqsJCAHV0s7r1jCl8JANpFJFrTa6fGmk8Z6lJAl9kasPTcDsI+3WT4HkKHHc6DolWwflA
1X8RFMjZ/ENHyMvTyLmKbuMBIz5PxcU/kEPUGXnrEPufipR+QvFDxYuZQKraW/frGvneyje7rvj7
asIZmzfGYdDJCygNs1XB6aUd2RDrNNJtTOp25pwD7saiMgoWb9xqDfFv5Kk6u4o6b4T0tt3DNl/v
+8VpboD3jYrp+tltwCxSem/7cFmw877adgvOU6XFT6N3uH0WPWcqHj0wXJAamyRB2rGeLSu5nCvp
CrneYU0PKNQRQgnp7PW4f22OlAcHqjLlnNA/46zr5koH9/M0rKZeYiLkDFGbFU9hoasPeyMDvWVI
lydiu7QnQebJL+LNQOE1M94dl4twnBYrFHj08rvcveOviExVqKUdHsvNtzw0e5HDtDf5fP5ysY3F
7X6t4523aJ2QqJbJ4Ffth5I7Zn1urq/57FmYsoEWai8wN7Tm26HYnFoopm2hKnsYDc1iStCJSKqf
KN5z+/kFAOSXUNPBng2O5HUNPkvpXuIt+mw0XzQfI85zpytLg6wJE2njDbII2Ln0lI1zD45s2RfT
T3sq84LgE9aJ6xS2p+LkxWVT9coB4OSR7Ul2xLXtHS4CyiTWmWforbXdQ631EGKQ+mzuGSlMzayo
OVMJHdtB0czYi7mfAzVlF4SGyEri52aEvj1HFa2+SGYYvNc5lf8hiuJlesL0YmcxFhSGo6IU+BmG
HChbFTjDurNoD3UQrIjad+OjYYW+8oyYEo1tbUaJCbFtZLukJ1SJuKoK0vlzO3vu6CPzJzgrinX5
Z4NWhgtOBDyWiTnkd2fvDdyjZER3/4ndAx9U4PRp0hJhAOoPNwvFpRgvajDtugqwvN6RuLyt34yI
l4G3q72ZjzG6GvmFCOA7+xTFgmmXiydj8qgG0nXW+S5c5ISvxZJkMMIcCgvwe63oTaCqnJlpyxsl
BaWriDLtGMuqgIU3ADUbRcfIldeXKEq3HcfyJ0HrzZGU6VWo2RyilM4KHzA43LRU9b2h/kdm+p/p
BW4t6FUndsB9HO/Gzw94Al4Iaeai1zjxUloNxzDHb+qEjuDAjQcZUuY/v2elARQrxRXbVj9fG4zj
LQ86+q33HYPrbkbzKMhuWwr05nkaGscf/EyrDKXesb21XBMHURV9QhYQV0QlBxQ6rJ6ZSlSJ7CfS
SWex5Blezn+NIr0JWc7JzHk9MvThiQLKlFR93AX6hJqSAiukRH336lIoad7zi7Co24UDPqAz8WDm
UUmsHLMvvLhBDxKhdumEggYzRCqZhrAzEnHytvqVCu5wLJuJuYW5V3I2XNivex8WZeSB7oIFaH3E
MFiptilyy/t02jq9dw+eW5ruoLrgrhlTv0aHWq2K419rav7sVd7rhaxcUN3eEwqiclHnt84z6iuO
QH5a4nYaf2u60PFCUAWJfXtpDi7f1fJG2YhVcpEtKyuGC4p+j2iQABQmnAdO1+AMm45HsqbfO59a
D8M2uH5ALqzqJxkhp69sY8q+O0DPaAaOyvyXEwEfoz82Kd+lmb9C7xID6f3V2bzK1ujFDHaw1qBF
uX5RfIpZjhHMlpA8EtCRyhNs4L9z4bdv8F+m74RDrdTOMzlwOAvkP4oEK0h59UmRkEjWEta9LwwW
I+bss12zzB/wO7ayAOmvOkSGO+iCk50pxGs3PLcSWTqHa5dp+21F30gYtDDVeVlxxnrxXtTVnEnK
FzKdMMl78qO/ZE4CIds1gl0KdrMMz92fowNfIzmqYM4ZEHWypHa7CqZpKU7Iv4BGIZ2w5HT+wQxR
jaF2g1aZSJdm6r9gU9Q3cFzWJ5Beg9obYBISorgPI8Q6a23pCxbaGPOdv1h6/UNwCrj6edlF/hfS
h5TTKPVRKlTAe/dQY6MV7MAmOTFpHC4/y6HjFgQwiQKwTyXvPx+1TO1YUbyaYFaPi4RAX8w1wUVO
1XzyPWQQj1Ip9w7YtcKssi/FnzbQhIXKujb8QeExkWgEbady8frIrAh+sZmp9CLm4cw5D7y+iK56
NWknNUfuBdiZgSeJxmJdxR7Ox5LwQ0x23cxIFvuKh4+qyNIwe8uVTYHXnb7Bigwa/obGN7pJDFiw
Xq39ieCZ2KspiS5FpjCo/FVE0fmi4rjXkd6/G4UFMlvXhHFBpdpDNTHaA0XiSdklBgZKz0jNvo4i
ZNuabTaSwDOdLp/b9ATIwxhN7ShTf0E3HJ8RAiKot6Tnsp9xA/0UicwqhbA36lUpiV31R1zJatx9
SBIos3SPfstLm1iY2fCwZb/lr9FmLlPUIzvinw2wnaNj0Y+T7NcsQbpmKLzAfHf19l+5Ztz2yCp5
MmwFAQygT8sVzNNUgrTenSTmBBTeVyajpnbjQdKjWEBBxnYS8DOmmTCkfQe2TZS8hf0cz2on6J7q
IU9IA6qWMKhsPorAkjY4DkpZdv1xYhgnluxs7k4CiN4ccWaBZ8q7z6SO1KKwjpzVwJ2fYh64exdv
aNTSEdDZc22jbalaTuPsHEAATBZZxkaexOADZMH3NbVQhDwYZrZmLY3pB+zyl/uCQyIHc0di/cXZ
bVCZ+DrqbMCJK2AmXAmbdGctSatvz+KRbsW3UEzILY05quzMXQ0AqFRNhdI8buZVwRxS8Oih118L
cgAxu/60rn9jV53uYOb3dnhc9Ftz0/rMkHsL3qiKAb21N6mZbDW1Np1ORA7TlRS6Se4RAVtwrpgt
rOscSX7/4al5ADhCM9g669q2b1DkD/PpzFKcgIIe79rmSvyuqjcBHKbCrQJdjyi7pPx7l+svK86j
MjDMtHA+aGlWyFKU5UYCTcJspeDQvgVXRqRJFVZOVKq2N9MRCumBRbvUyK0DoN1U0NLZxq12ZEKu
Sn+goFJvsqcp7b1Cgy45D5yr7J0FsdsUxsW2uu8MSkBLnhTx5LvjpmAMqzbyzuxBgQXbdkKiZyM2
MeYJn026AfJry2P999SLHZrJmTXViKw7gNuzJcN+rOAdEESLA1qsznVcT0g84r2RDYTPf1gU+g0q
6a00oUoEMmMTuc8I1+6CFo1MegdDiSsUsZ1A9dY9JevVZs1lyermbTXGJRdKXjxas66yvkdmqjyY
ni0tj09m4vrqPkxObwErhZt2FaKRSe2MP4O4fcvss6fsZuhMgkMnSSgnXtgiICIzG9fCJ77KkKSF
77bu/u66cHPVIWSoqzetxBfNTOmreBVFfmyZWahn9AP55y7PW0a/AiJSaU3Aw+lZdROVlmfY/fTg
ebq8EpmE9rz6rIfapkH5ycgFV8kfTMwRozH/SGwC0bUrk73VK5OsZebeU5jxtV2r3sPQA4CAA7Cj
GLeM5HxWvEI7fLen/oz7KFug5C3zVXisggDGwJzGs7x6szUdXB3fsxISot2EWQoBrAscwKTQBVZa
YStp0G3ZqCdso3TUGL6z7Ynu2jD+bAM8wa+D3gFi91uIxl4n3Fl2cfuVSpvo/Bv/GKg1eeka/tGV
Ap3TyuH9deRwiHaQd9dne52NkaQ=
`protect end_protected

