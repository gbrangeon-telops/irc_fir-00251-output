

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
rMj+x3ocDbJ+0HvlMPtFLLYN4V3iOWmu0i3VYcvwPU8r9dUqilqv5BoOperD1z/j12cu4ait0bNC
TvgieQY6qg==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
LiFkBwHJvbvIRsrs7TuS9x+hbpgzWqPRKAN+86jD7W/DWOy2HiTI+Pr3kejl0F7PQ/wd2Tf3u0hB
l5PFI7Uciy5uXiQA7fDmYLdPcNoMNQWm9hohp6Q8wB4H3kSwMFgjlrwYcv97jBF9K/DD+f6kjMEJ
pjxxREwM6oJfyPhyhBI=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
mlNr/JQ7BAznEw9Lq2hOb9T0FUxDG5TxOJH6VJoPGS12EjdrVMK5Jwy/CrH7dSOtWY2eUHhpsxFO
HZJnPHkoY6pnOp56kFqNAyiHJP+z5BexlWOYCHMzTTDXl5ecpknkEs/jFqX2DjV6R1MuxPdeXOjM
JpDfpA+rd8xFCgAvhOcvKEKjw2lJmNukB/NqmGdLZU9Yd/iDC6mJcVuTrR2gzFDMoFjQUitH7TCG
r1krtYbVQjkm691WyHmxufh/qSc3KdzrpZqycBevqxjmEqCq0nMXCiMyQRHMFNk9XLymhnx09LIk
8Ck9EeU7sTUKIMhZ7oB9NRbr0Jmue7w3V7zoXw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
jcrZIuGwyVPSe4eEqA3CjxEN8wKBf64m71qLvmqrllZ8mLFeyFjj3f796U4fol5LeUOSCUITklpk
5B0LZiT34IugfACCFG6eSa/KnYkpqdaiyFEJag2zBthAbQTJIoKzv4hrVDSwoJffRhWS6ZAZmMOH
9HJ1Z4KODhrBj2PMMOQ=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
He/hsXsp9htM4v1ezeHFxTi8NbCInK4GRCTZh00v46syUmSwf+mXhIjhLm4sHKCSUqmWt1TLUp0m
CWcpoGxiawBF6wEpl5GgUNyVTq+T/CrlV9Oykyiw8ESh1/7hqCFXSES7D6yS14KOyEm1cr2UmC+u
X/NTzDDvOd9e5R6zaiks/z3Qdqxiq6f6jnMuQiSiMBsAMCHxpq5kEezVTATURKXvDebBjGkSTomU
Wve9JRKQPSiMHuUURnaiqzi8t62PeJzIwk64jI0DQYpuyHeGDNIZt8qQokGYPimAYp9IilmsSuGG
FM6CnM5XioVenoNWDUkk1F8M0K5I/5eHgYEnkw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 30400)
`protect data_block
bqam3pKRbgX7IdVaUcUR+Fj/n2+yZtn7EP7UcYWLMB6IyKdnNsPaLu6IlSHivr5CGUOS3oLczCJD
g5hFInSv3ra5zk1fQrlAJ+fN6A5rLv9wP+19GRyHp3fUF6xOl8YxE7J9Q2M9ERp7ntPoVMUEpa8v
VGiQVRlwp16oRzIhTTjB6oJeHmzxHplBjOyt35cllgNK3InyyXbh2BRSQZm3LA6ELnuuEm30HKz/
k/V8NjqsNz7eTxA1TOcnJUDtQG3XyOsgWKDMiB3pJbwbDdmZCa0h0qjNSN1/P7VRRNba/KPlIwKy
bnMGMUAUk6jj6kAnCazYI6Y2fUAuNAAKh/CDqRCRIbzfEhXYH6y3Z9WjAZfrFoAjmHajmoFk8ZU7
Op5+x0FDMI/gFY5QORSlL1ACD/fCpR20e30ydBBibtPmHQDP5FBdQOibhEWQkH8SJRMYIJ89XKyx
/h6C0Qs7IhZuknAX+onn9AO1zl5AA+9Ma20WZPA1yjAF+mOcZVxQoicVnfY/qaDtpEbtfLOGw6NS
uYVCWIc2niErs3T/wE/lFgpAIKKbJtYyGg6LdAe5qHasqWh1NvYnU8iFVXnVhss3jsofKNUpMUeY
COJwz4F298riBTSvetZhBs7UKNLsX19mEUhPbcG6r7LunqPSFCl/c/9MTDAdeldjVoWw81NrMFYe
UGzIEYR2nV0SgSs6E8FtfVBxHG1FpsivQXan7sPtmRN2j2MfGX+WifKfOAiS6mYhAfPe3ttLSfCA
p4LyZYpbX+ZFMylHCA9ntiQL36Mi5X3qISeCt47HOyNOyxpSSkri67yCO62xw2Y0hxM391jjqCpj
cLd/tpwM61pJFWXmgPlxr8nS8GFKkVNEsPTnSfTio6qzzQ6nOGAU5tHHVWN8S+00KAFIXo7ZUPj4
WEOVQRsXdJ4Ja/ijgSjP/NJgfb8vvmReWftdEbxtuFTsjGJiC4Da7p2fGYwD8g8m7NSP0mf9Jo2J
baFAVGz7yMGUYxF/fHWFxaBY1IDTZ8iNOdm2ShWJsSdw5wN+flKC3sIsw8wWo92mujn8zPRYdzq9
G9YYaKTRleD3Nw/tJHtGRyCQm5jR1gFlJNm/XbwgryOyrC4UBCGIe0moRIMRB7MXrJLbuQ7UApaL
Gz99vAeovVWHnL/DP/JZK6bGqv7gPFvMfSv0ymSt/5Fo+D2Ul4BKpG/L8YW+Acr7t6dGNy+ynvjx
KLPp8Y+nuYLVSSvG+NCvmv9X7Dzu9vjjsaG2EV32NI6pbMqIUul0CWyzBFRdBJhUbAsbPbPWjBSe
pCIf6YM9ds+rvcd3gw3FSSxituj3V13GFLj2mdQ6SZv9aQIyDsCX4g8USYP9Adehz4RcYoEqy0jF
r3HK/Q5Mr67Tp/ENWiRk/d3SIt0uR/NSrcWOwPA1DTOdilQiXBPmziER7qnX3pkfm81xuV0ULajV
HlzMNLl+ur/GPf15MzKHwGDe8YPeCF5mu2RiFYG9lRnihjtCiuLBW9awWK4H6TNwPWSSS2hbfD84
Vf/Tqoyi2pqh806TZTl2FuDnUGvfpBSDHOgxTWctolIBEiRdKhrkCqznrPWZy4BJUHDz3uQYNFlf
XnrRYwaC9YfKGYuaPKrTUBiSn4MrKn1USlfdPID0GmodN9l/Tf42XwIrg4C3ieKYbl6zfVNq5PeS
waM9gQqu19eBSzMf4Mfwsb47tL8zAJyVrJxJBS+uizdtd4Ts0ypFPprFCKMH+ye+z5mIMvtkHNJs
aU42Zp4VUbBdI4OZ2h5SadliylNPP8tUpG2O+dZKYDEWUmwmypfKVQuynL8nb+S9vL1/8uINE2Id
Ywi/k1O5CuM3snHIq4vpku7IdAszMsgwV5a8EoBM4clTFDSA8ewNpq0/lAKitJFf4Yg9ahVT5Eif
nMnXrqucvQgHj4mBKKpRYt9iUr/5jutWr8OuarGEAmJW2KQ0rNHRRAebIVvvOJ0ZJriZgklfeGA5
6zgFENOwhXYmsZiy9wYAVlts1sy1/3UWFgYhdnJTLPTMmQ8jv65yZ4n4rXGhv8aznOB7z0IsYXmw
cJt8aw+KkgepgN04KwH6n2E+rmxt+6JMwvbWQARW4/uOVAuSFJ9yit7N6poQ5TmKKK6l4XcRcLf4
l36Ema10l9EL1KaaTEr98pnySBEYMUDHzjNXm5IbXJ3/gMsefbhfUACskboq7NE/Qy4OxF3V5xz8
ivm2CxZNpPDj3eHxRX5/fQHwcGr1t6Untiq8herbvEzak0MNCtSamZ7OixPdJZcjqqtotPNL+sF4
pxFnYcXEBcu6tuKGyp6ViDc0iH3FXA5Dbyz5/Fu0tNdxqXYDQDYc4wB1QCsWdh2r3k1/VuG7xB5l
Ea4j0KgBYIeIWWWXb2VJ9whZzmV8z7Cp6PFhC+TO50iyttiom1yhOtjMR4xsz4HNwzkXIES4jiuS
QALE2ZcflsEiIkKnf2i0Zwgor+BADMkmT0EnEKHmogvcz68zY8VocHHD9His6drBrQx+eU98IiOt
chhiCGTt0msQB3yl/isfoX18ICSjG7sNZInmW0d/RHCTILE0PNxbVdrZdfatb/tCpJdb67dLfErE
MKwWwgPVgBdyrVtKrMHBtyK6UIU16j89Ppbxl09dlHUWpdNK3DcdW8zZSYf0q1gLu+5TZLcMJ0TY
/WVDCi8HS+CxwAg6Dw3Xga5sGnkefdv7q70pGJ52W5ZeKZctcoQnwAEbTIj7elW0LYQ31r3ZERq/
N6wtevWJ6DvlkOKFJjNv//lZEXwvlcuEByLm0EpZu/VJqLj0r0lUopZhU9LyGBNddlV23dFcXL+O
51cqXfOhYRPWodmgnhk6BWrIIRA9t7KNw8Jq5cAlY5s8M+QFJhrjyBW+Ar+ZRbmcqB6mgcvwVRxf
Sogh4My3mDy3ftGrCNgokXlNL0ISiQY5jaavUThP4gtF4UaG7THUfHGlJC6uN0LnT9+QZh3AkUNe
e/L1+Heur8vRBRui7Dj5Ge//fpT9LCFyc5OPdcK50CYu55VmEIccXq9NledC9zEVkexy2WtA/7cM
fw2+BnjkzUka4zOaPx2SgvSwC8xlPmFWDShnWb8W0Q4ueXULXr9uzA6pQ0KIYDl4mXWYLRo6Ll2b
0z+6X1kVRDC/GJavbTG3S+D9yhxj/+oWmc9FATfh6Q0knCm9JzqXhqF8+AlfSTeeIqzHg2zczcKa
kzaoUUuYvehatMUbNG0s0f11tqLOt7R7UFPdcaddjXSIieBeuWqXhTInuDv5qbFnH1c/tFIKP2pt
qocA5ZqMVkQDB/+Cf7L4tXstUjWMw3mYSKUBFNJw36VHzQaYmEMdlq9bH9Bhyq5poJEH+FgUB5JR
1kLkxXoujqOiTuOYNI4VD97NyaZAfR0XhORVYRSChGCB6i4Rcl5SYQ5TIcpC9Aw+zCqHEDy4KQb2
r1NmGEWI2ROpnJrVoHTJKAj1tvC1pUB6+CLgsgQAOF/H9AjdLAbjlmdaUAxyf6znYsDwPFpzr22y
PAE/i+0ZfvZsvYBZZWFI/F4yl+Rx8zUElg5P+uBs3SGJqeS7NUJsYuur9HAuGXpZLW8t5mlX+V2Y
JXBkPF0oR1jeZG1lw+Ubv5/eBiC3c2JIGlqDAXmaGIe2AYj4lR5VOt6LO0JG8RDuDuILn5/BaXft
jDREEeyOcmuX5wafm+0NrKpNHCGwxO/xBcqWKvopIX9LlmO7Tsp6FBeXONnUnWper3Apu0BLP30a
wNlVlawQLEC7Up1DdsaGxZYCwOB1IIYTedqp157NFBeI0ypbNlg0dXgtcHGS6JeJurwrYC5lLkRl
OuKlnO0FRwt1HfwTLdBlzq0GUbgqCZ6l8Lw7HjtbjSXiZ69ha/F2BlJ5gtMU04A4pEldLhmqqmOK
OqewxKRUNWC8ZbWZv16mC0srxwyIkqJQDTsQpM6UC0LIOf0ar1FuzZsT9dK3ybnZnNQWJvW21WX9
NOaOKR5I08s8fOdcTzxY3DAHs1HmPR3F/KpAxM2/t5LK/LSOiKTb5JtSmwihKgdEVZ6AxruhvqWf
Xdu6QWuQ1OHTSZZG4ZoDwnMy5P0Siwg3dgXk/jf/jPGPoBWs1QOQBI5jX5jc2qFGyUqw17NyeK/C
uqqjnA3YccZOm5gxc9I2JRJilBaZiATh8p94kU2cLGJXJuzHhzfkG2fkOz5UqilROafHockQKZH4
PyfO84ntSKi2TyaLt/N27oytrABL+SSD2r7h9LOyL/WA7iq9QoIEN18iPAqHjsBXCniq4FvWdCuT
0zb8jLZDLesTvnkN6Efz2SyBygegJ4HYrG6iSyvn4QtEMDVevJXmKbQu4cH8YbOw2nzSzNBiUQRp
78qnWh/ILTiQuBP5i3CL0mcbM0uieiT93ZgluL3n+tX6YzHtwf5oG83+wj6tzOcQ05jD8s+1EEUA
mdG3T8lZvV7ZKMbrryyXv+AersqEZY36Woj5H837R4r41xwJShuxSLDEZcgPsE5kdz3AnQEZH/gq
mS/gykUlv3f2h+/zzaC1xBLyjzPmYGcx32ub/C3rhwxBQeI1x9NIIoe3RYAuDz+PKgJDgb9NODzV
5ZDZoFefHdt8F5RZNd75Pj0l6IKeEGNfNqfsI612VCJPPlkOr+hMEChGPr0q2hQJKANC0JGjs+s6
olplOa3lG9sVRTNE4srBQ3wxyaijpfG/IHmLbRUd49EHqQBLnUcou9rAVR37Wke9/mHK22xeuLan
hWpcXd4vbyskF5v9LavDhjmGvQZtyrhuj0SBITSQ8eNC3GNH/Eyu83vTLdXuN6qmFfRryHUyyx2F
7/LWoieIVRkCQosclVnmS9iQa0r2qahkv3UBVHl24miNJrCXz1j9gpTFeNIgrrMsEKubjzWqyI5V
RzsqU5lSz7ioqVwjXnS92PklMfzNh+ndEDngVf410ogYbrGObMGhBOfoS/MWEFoPgE/W7Pc7lMoq
JvpZ+9yBlnp8qw0azpcCyQdAp1FCsks4qXae0FJeescRTZ2CMIqXJf06z5Zi3O8e1e9ElucwpnD6
73QwHKoxg8+zaB3ggsOpFWn3jrxIiviU1kt1FsXan+WBI3oEQaoHd0kIHPtumgiYMZqcZGnwlXja
UvfbkMRQEF+/X5iOAC1Voc6zBhhU0pIPt9RvIRg6VojIA5PzB25bP91CEXULUG8fYTmuNLeMn9KD
jc3Wm5RogJ6LflCAPimQeThCrolaqJVXx4Z+5s3aHF77yFOV/nJA7oIuZlmfS9ezqqaCFve/+k/1
KMnp4qBoaEBrrjx6V8tYiy5xFHBgiE+gWOcEbwQylzD0ogyIhKBDlincJhCQiZS7cFtCC/XTHAeJ
Z/+JQFldGvswY0ByTLzmQHrpYLohPqgbQ69Z0oTqIQvHTwzZvQKBtCQ26dA65tFBvsFdLa7fpX6s
cer7B1AAhZXMIUP+QSBuseH/dO7V2quUnIyMXR8FVxRKJ8+RrmLgGF1bPdQLjliWjqHCnahbkKQ+
PfIGQxKdKQHJVFLrR2O7+dWZeQ54oVm4i2Y2UOg4ISx+yXMJKwyUUTb+IBGAoh68P0czqnGQ8Pfb
ePHz2iv4V/6J2XeQsaXD6fwpOkPwFxTmQOAvVsOAsF7r5btdqhXy02pRngGHaF5YFSG9Pln7g5zr
358T++UA/u5LZ7reeCPNhVg54qBup7+hH5vdHknbgHXJ04+8bR4sUCKaGx9BopyWIO4JKl6k7EdN
38ZLsORb/3oJc/Q9fLB33Jk9r1+nUHvNu20G4jGXbXT4rui//uemWWxVUCzx7fgvifvKig0Dcy5Q
97tvTH2CkE1+xwVrrD4Bgs7vM+tLoG/KDxz/oo8+hgg2zn1EBnsohH2oVWhTTbKiFnfpczyQ/1Ny
wBO7pXuUVi0LVoAx7c078Ubx8x1lLWtcFmwxCNdzFCUk3hdLeMQx64WK1debl4vDOyPNJBiHjkCh
u1oYIaV0BgkZm9Dou1ezDPLMDTZsgb+iku8XZg9SWOwHSi5WgsmPOCCobdDcE6hA1q42ah2xk2ip
8Q1kT3sp2UPBFJNwOzUcxiN0qVeOKdhmVZEn/4oaV0UU0vJGcQCbEuo/+qUDiOPfwCd6DEs4ENGM
ohV2eRmshgqoUvfIHJ7xUQjj05kK9/TZ5SmLrgRjcSgEJOP+XQG4yEgzX8OkpG9O2FWxrZ7ScgEF
7FLo+4aEE2zkoDWXp2Mw5imXJcOvu8OP+AE2r877sC/8dPk0p1weudKdqrcPp9vWKUzMrNH9VJej
CAaoQM1ytnh+yMFsMBgp+v6h2+BDRrAjXU5AxtbkiY4KSvGvCwnELUTxBg71mL9/y76Z3ZyLQjeG
ZT4TBv1MwaqrtM12OJhN+igfOr3rKV86o5jAhJk5HqH85y5vj3AZdAlIZrOKrLxWF400I+1HoJrw
5QgEhcTqyx3rdQSgqo3JlnGONj1HEExVxySIpEKf1XGGjYoeGTepSYiRaJbrcSCwrfcdGZ7HrEga
FZ6YfPHDssxDfSjlsq+YJjBQjZNX+CrqJyl9Zkk/mGqwqBvHb5zO+vChWnXlOPJLC8hB8QvbXZgb
+a5rHYB6VniqGF2nzCsj/eOb4A98x+qT2lgggKgZGRA09Kpyl1QIShaWy2P/YoM/zCMXxfJNOb0f
kaQyyKCw4BKgCw1ErL59VnGHI6DUB63bR9R8/tZk5+kfCRSd4wdkg9gpvFkhBDFuLo4FDxk5uxT2
j7zQkC1g/Aya9SEqsyYpjHrpVIsWe7dB4XYTISOlS2BpB9JjmKpD2ejz6xGnCnMxonZQmhQcWqFS
Xm+5aCz2k5YbGrAGZCe1FWxED4ooybGo5JkSglSuJvxgolUqxIGAzVcub50iquHL24SqwtfaiUrE
eu8KL4jJShV/UrlL27BMI/tTaqxBgtIMHok/gz8bOqgmmjnnQ6fO4h3BG6FbMwcy/OMpg7gfDw3x
Y9bsGDNyOfJsLQ4+UxsnEETN7b9UHDvYLJHDZ6GRKxQYCD3r6X8eAFhUT+IBEQYnUfYj3atQNkpt
wpIGvawlcCJ0MbVuIQH4sGKg3ZX/czw0ZnPTQ1KeRP7UfGI4JCZPZprNyaRPmwMiRtefeOkl6Yrx
F+q5vgtqdmrGBI5pMwwMs3osFGkx3sTeuPbn37Vi22hVpNUlx5ECN98nmQ102MxcOjI/2setvMTR
/BVg+pDBJI6DSm69JGnzLJZ2QHdMqvFj70AJZbL9IMa7UFjjhANlMs92oXMl3SYtwXqTq63Cl3p1
+umuIncTza+jlQscJAa2bzEiAge2IR+DvZtltmT6wfoQVLZFFjIDE0xMRmbbQRdXhN6JAWLawzx2
AUdQ+UBaFKFg2YLhL8plhb5I6Z2PFYAQLHRYRpaKPcezHPl3X1FKuXrRTWv4I24XzbSJtAcAPUru
BvbsBYM74CRAiLGF9v3RgQy8TtCy4YVJqgNwQ/pj3QaWP944S0Ioad7kqsxfW3FbjByckHDk2nFz
5if9WO/TcDlhzL/uHbxpQrg/DLY9vQXMVDSJT3cJhLop2KvZYv1jnsD9WDAxQXM6e/uV1MtTOyXY
VWChgJpx2SLWXBzNFj60VOj58fddxV1ezfI1MAX3IStgdQhelrBTXOAIytDvPnCCgvPITnF0vSyx
4u2ctnOSiejVNIa+WNDokLi/EAoBBzSzuMsfc+yDUGltd0yFt/BwzBZUanIQV8WlvDCQYk2dNtXt
PrjiOkcqCwtWcpJCJWRXa1cVrdnNd+WoK7Zr/gzyfKv4GPNE8vENmdaOz2V2SgDsYtOKG9KtiC6q
ZfI3Z7LTapP4lXEpKFpFdrBFCb7eNExvaG9dmD677xK4FgUViFwS3JjIt9aeImZF7q7kZYgNAqr4
EwIbU8SffkVHv2XaFLQa7rsC7tqU9pn5kh4t6r4o2KDmaOf4LHXgZJvN71x1+fepEYHaQaGN3D1J
fMqKvevw6Ez8ruWdswKhAYVJYl41z1KcIknUV5GGizEKE8O4dgHt1RYukrNB6XGeZsCVh84wznST
uWF2dpjZJT4p4hjB/b31s4hairZj5quSMPvbHCxCN07rbPilu3YR/tuKPDlFBZPeOLFvi81Czm9R
DhxkOwKXIllcLc50PifNAMJdfhtU1Ur4eqYsuhylbvkXP0IqtLyeXlsJ2zWoMv+Os9Ovw8g+pNkZ
S2EVvQwOOZczoRU+wkHBqfqICHrfjHfrW50zoUTa9Drcqb0JnvlhILD8heCD24I+UiIvTA8dJqTH
CTi5/5cdX7wLNap5Be3e3e1A1yYhz9tN+IhGZekxWNuFCuXHpXoWheG2jx+RFT28YM3mfAYIHuHx
68ScVW82sy1h4Rs0cZ9RRCP/kNTiEJE3BU8fD7pTluAG+5xh2hDjxg/b/dEx0+pWViT2fhkx7kbr
d9IGz3Z5fPQrhmiEbW502iekDNNn9rgwG1vX8DoEhaRbMvHufyowvDb0uDKJ1p26E+WoMvCY3EMu
Wv9G3cu9zGO+nC6KF+/+H1ty20gkrna24/XDUVzDbHhskErhspHnLz9wVNiUBrQXT/UMGrty8RSh
7YDF7yEoVvdXCPa567iF+2+oUgtV2awfoB4bSi6QFGB+ZTIhF9n63N0MJQva2WLcOIxaEwFaSc9T
N+bY7Me9UZf2r5d08cFfibzgAnger3PvQBIPXojlWwCVr9WmQbLwIa1xJC8JnrdZJox2uDQGbIY9
1n9Tadl3KHsZIm2uGvN2EcC44/3NVf9AS/WJn8GYR2lzb8mmDQEFJKELq9Bl6q6WC9aqreDrNCeF
7dTyOSATC6f85+PNqoxJRxwNx/lClz/DHUo9gKGmJDI/B5idUGJNYA19lzq4wH/xlYWuv36cdj0J
yTrqJmKPQHtTsGFv4oZ+iClKAc3azyh/pk3xqWQ6ALNJTDaIXpIxqICTd+IS6cZpDO5ANNFS0cH8
/kbF5A+6hmMdpTN3JsO2pyNXsvomsGqcuUI/D1Oqy3RjpW7YbWuEVCK6rfkSTYhBoIpRgDDJG1MW
Vc22WqIZfvrmVJaehnES2NJGvz2oaODRX/XReWYLX2ditXRlVpxADta4pkm3qUXQmknXuHyPph2k
tSxn8sCUgIZouFFHUep1tTcc99VGu5jrcHoYK2sYudcDEuggPTR551GTyMG8lTeqJquQ5K2EoRSr
cGCmXsOanhfAeej5mC4omUIzyZLHIXeYEoPz1BqWFkuHep44BOCeCXbOtefaJFdDJaIldD/TrsRA
txnlEsG0uTnN0v3rfYAc251Rq3Z6tz+qoqEp21rhJrbkoWeFRPW95AbEXwe3BWpGr9Thc+n1q8G1
/tjmm0r9OSRacboW1EVwz+MJ0De3KCdsOZP5eSWupgBLUe91VbawJshvghVA1GKfSxRk01iSWKjr
/DJ/7XpnvdbEi6LpNlMCvIp9Ln1VdSFO1vaEX9mCVMMA5RBcb3HHpS+4xLBM0RMilVBPWqePve8V
80cakSbCAHgx6lNfQXnBbDK/xLCTOMGDjlqq8yVN9QvIib1qQOt9xPT4ZOuX5L+e4NuzH+F3yQYa
Be5qZPPuHzMn16HledjFK7mZuYdg8oMuNonbCXHPWxxayrXFAsgEnWfLjlsbEKTgLo9zphybHhJl
N4JEGQeOIR/6ZkhzsmV+Z8oM70FAtqp4Hlm78O64bAFmboOiZ98UpE9LpBPNqiFo1XiPej2puE58
+jLJ23GuFKdy9+L61WsykVLtpJtyv72AV45Llxkg7Sj3lsu+NU7D9PrNrEAWrEFhpeTKifTUSg1J
mBsul4nSjrgvV/2YuxOhPk1AURxxneLXJw8GezxuzoryExqgVGBSBtcHN+RDd/687Zo9oqaD6VAL
+Hz/G+P91QUlIKWhpQk5ItQuutyfiokdHFFjQDlejF+MPEYDFIWC5T67kOn57x3abA1ACf8u89Cm
RRbKraH9ayMmM9JbGzLNTUNsNQ6wXEnlWbAIEfeQ2HUtG15i2FVuShPKf8Y4ddWKvUWNW7UW7Aqa
S5seX6eS9Mjk/FESJkBlkZ7rw3ZVdSx1e7r6XpGVpxxl+BMH8/I52oLdzgZd6Y/bg+X2WYjwy9Kt
UYlMtU05zDl0sff3oE98tbVOAMkFPhxZFf0X2fVX8Ho83UwplCMG+9nEqguwKZRcdMduVH3p7wxG
4bxa7FxrLiH5JbjB+CzH0YAUec1NI/Mg4J6FG4mHiAsUN1UgDrl52cYBaCtX0OycruqO7RVWsvUg
k7HwclmJk9OeFKm9E+Ng7/NpgBVCoECs8BdKiKswG3xV8qIUfs0RcUwdKKWwhOIOVCC/hMZZSx5p
d9/yQR9p1wVqqF5j4Xvy7nfeKKw2pKxn/I2wQl34hptyd8RpnSk/8VE4pWzdUPNrTup14/Y9P93L
7eCLixYDB0PttHgIVKZwofRmWKUDulcizw/l+zeR+22x8Nw0G3UCMzv1IU/zbkUpq/ekOGVQKnpe
kWrZm+3MKJc9Nd7C4NIUv/7In2hHFcFBO3Kb0ZWbkfPQsw3BYIZCfZotQmp2wsOn9q9a0BLp1tx5
0rReDmBnMwnSzmB2thaPFRfekjwM1nTttjJQSsSZnuheLxVdeyWYdK/ez66MJm0mC843UnSmb5O7
zq4TuC5ooTFaB30yxk76HpPXR1KQNvVxnlP6X+vhb4JhA81C6pMKvUzokkINYv5cvqM3cLVNPE1o
0ehfALwzgqHNi+MLmbtf7FdQHVHZagGSJLje5AvLbCQGFpTpbDJFXMwHemCy8b9hGL7yen7TF6fS
ACfrH46hOl5sREY9MpIwte8E+vnwhUrK23CuLkpWpf+k9KR9gcKSYocjKLY9cC1Wd72LOmYJMS2w
JV4i61ELCcb8II9LFZvriVOLvr9C6dErq/hH7bxplqrvu7+mDvCX6o2d/wvb9d0WIXwfFyF4bkNu
qJ8f+IoLJNUBaG/vgODQhU2XgmMGgpMx1qhJtosOqZix46fuk6gcDiO83sMdDV+cEYXRdcM0po1E
ig2DSd1QaDnU7ieTYY//B13eJwLoP3MfLKvbUQeHpz4I8t9m4bpd1hq7D26RKYWQuQ8sg81sykot
Gi9+3YlIBMX3u9i94veJ6VUv5rsO2obxZ5vptbG0cnzTKqvkI9OQXlRDBT/JpwHIbpWXL2+PqU6R
dzqLU6ApERuFfL1XZl4yLpASrdUfat77hOrxcqcTWxrdSbZX6P50Cw4BtwZRBBajASTqRqSUqs8/
slvhsyIczh72lRHwTvFubj5kx6VWURPtjTMS1+uIhBcGQmCJI7tWbpND7D177FWRhOz3Vkvwv4A3
PYy41mJgo8swBqX5VtbK7S6bFFZ22frmETqlAkqJKzRuP+Z3OFfBAgMn/gS8kqmJX+OaZwBDonld
fZJGwpytkRVPJcy2DT/4tDcjlMGhdVvimAD9SEE5+DBYgNAYry9TIIPqotCIrWXw+96GepqtGhgE
8RgR7dJFxOraIhz8ajkb8/zY0VJBTV7LHYfw16GUtXEo+u55gUkqmyViC/dE7kOlN/Oeru4Z/uSh
XNI0p9lMAww703JOSOaodaGDLSWH1o79h2hJ6iJlC17C0W5873wDZ9bbChTsIPt04UiSHJaK5ZIX
LwDavXGe35n3OMrrwT7A3m5dE/gK7/Gu4hG6FIW6tXdunIbs1vDVQiGrSMNIHVjFELuIesZlsvjy
Oh23I/WDjyOAKVNG+FaaXTDYM/CHC1SS8aVUWM2UcU46RIoEQdWnBwHUoCkX0NybIFUIArRnhU3o
6QWVp3ACn6qQM6kZ51iSzJmIaiaskypQbGfpEaX/y8QXsLfmApa3otWzIUc+JDvtMsIdCRw3Cmly
qibOSuXh3dKSSU0wgkMgcmDSmWsgqk4M76pWcGv+7WLpYrPnvUR+GjfQ7wRoTu8yT64WWJAkxVrT
E1AkW6Ykbc+88NBpVSNoKESGevs4ljZGKb2Hd1PAKu7j5kVDlmwQkYJ/faNuh5DE2KD3GTcyPBx1
uUa35p3o7cdniWA2HtMYS4u7/tDJffLIgIhSzazN1Nl4aiJFJRTpLzUuODdKyG4A0elzPODSmhCi
MWF3Cw9egMv3+N+feytqp+UpM9pa0A9BTjpSaKcD4ipkbyFikwMxvNVGafuHPdkOlJxlUiC04Fbt
V9MNKPcU73K/a9sCNNA6o/gNg25uYlUbrH76D6XCB8smAavq1E/A9qMDN9UMohbT+uWmFx7DHFUe
clNn+vWT6xZHVmYs+bBR9imVlzqxfWSa0UUINKQbw4DqIu6pXLGK1LDK816sIhN/Ww8AlB8+D3zz
nxOTtlC3NMw8BNbh1Bg//ESDJZqEGGmFEiQ/J6AkqGcCD9nn8WW0xeWFJ/HsSfeaaOaxhBhba1am
l8aJe6LvQ6ui1cFV8lsMWhgyIv2fqaaMiKrobiaVpGS/2wApeoGcLozAh6g7uPPVH49jQRqwmTCc
sNf+2q3cjsMtYj717YnXMOy6EK6knXAkf7E07dKPZK4jzx/I8mPBTzrFyOYJpssHaoRUjtCCTKs0
NWD2s/UvXnPE83cSGsLd+6cRKV462GkL1vmDJdNHb5iyQDv5X+/mMiTGQevPrAfgMCkc2T8oDd9A
L6qD4sqKjCW+Q0BeuahO7jYzGEL62b2I6eciMPaB0hQveAVBwU1e7kFH/vUJTxnXjwp0zFj7nSLS
PSgMYE9TvZq5ddCn70gD9p07S1DSpYbG3K7HZA/KmrFALsym/1r330udF5WM7kHXfCX6Rt0/36Bl
VL2egW2eWl+3AW7zq9OWef1JBx2c1Euo8vl8nGg6YBNVwyR2TYy+wAalwZ38unZAjNQnKRvEZC7C
M5II62jmEbvOMmEYHr+d8/iYDvVYGULVCKvaf4nb3fpam+qS8gjyjWB9yccCXevseucA22lyhrl0
vVuVRMlLFYPp72HpTxFYtEzwGSlMNFRKYORWw5snrBQvLQfgyeehc0QzYkKHAnWfIumznk0TzTiZ
fJ4D3gvMjFyRjfup534RH88jEuvsudhtVt8m9K4cuiHvyXnO/mfIXQxxBx4PF3rPoBZmQiLblaDT
N6aDVol9UNLG4yzWzbNjKxGukfmSMv+sMBnzMskR9WAFtzU5gCW3266uxL8Wpuj7z7l854Z83WKs
ZnK/TYx3GeSni5mHigAxUdrfq/IiTAunoa2iq0Ahr6Cv2NtY957DrDT0jqdUz02phpPbgdl4tK7Q
V2cCHJFO7dFQg1OdjRXeiqofViQMEwyeGrBb/77pLU1PXTRlRWUbStejuFi61K4zJszMQ/QRjfMY
254NxRGW4Pc3GKnfrbV/dbgsBfb7g3e/QcMr0hleTHVQzxB2SsLyl3nV6v8RBMDwn8S8p2hME4r/
jifdlHGaOZJ9mHifC6WMw5H8w+t+02Xs5KdGL+tw5CMaVtAuTQzWKYG77V7T4sVMkn+nhn3dTuLN
q0dYXt/0HaYBHY7xPyOokSzPoBVPALqg7L8iZzWZ+b+9wZLPAtz5aPfCurjbW6PNuvbCD5tQC+dH
XuE9gYoOXInqmBe6DZncGzmz7g7zygxHKWZBoPJG9inwIkNUecGYfFsbdpZACsTDxojXnES69Dya
F/JBMDj2OkxF7lNoYs72eoe49eMVUcyHxGhvf1gp9TVrv9XEi2WMTnGT+bqa2VjjcwwEHBl06TFL
4gDA9F/aYAuVJ5TT82vPEjgxbBaMTGpoftaiLbz9sWI6Dw/tp2VZDR4U4X3rpdnZgtk7wjNB+OyE
f56Giq5cciUdPitQjAAsojn6TsgddJA/RA2DlEweC0JgRgnzLbBOBYeVIk0D7qblUVQUNwZMOJnU
rvy27ivRJhEM5aGSkIWnr9Vq25fdNz6hLKsT5jFcGttnJkaIMW3vaEYpfs9N1UUyx7q84/hsvdUD
klYidNBruJHyNeUd8QDM3ZKTc9DLGia0CeUeLZuBEHhWhtDfRH67zRxrAgUXYWrY5+yEK6bpy13/
jS9CNwiTQI1+fHQ4m2Pk9g+xonE6iz3onlsAPwnw4xjbXG3NLz0443UwCzoCuGbDMhm2MWJXp0ny
IE1oDcwQtn8U0OP8XN+8tNg0x4nyjKOszLKk+mB86tUnjvKAt1Z9mHplRR1j/R/l8pZi3kNLhHmA
zvygEsQ+yvNKhYcOLCuN3+KtdKejJG91nCMS0L53u9gsltzEG0NrinmMZtH3rA1wdXLDZQQh+skN
qcUEb4U6FhzNdEXUzAQtqXBCRE77Elt5lQ3TVyi/jT4/dpHMerR16y/OxdM/r2iwCYFhzAXPOMLC
BNsQDLN5/8cijPEsg9TYW3uJRXH1a50ml/REOYMsFgGOValeveKktzK0eXmfB5gbfcFuppu+//Rx
bC6k/7NKPuSar1oqDEYIqqY4EJD0LPGpB/lT/3cSXYgWQUykHI47irROnuyvVyFQF4yRnRgBeGKM
1vZMrSCBRw3sLPD/numFfBEA0C1D+RVFDgXA55qiECFXNP0Cn0KnJHnRcMbVChM5a+iu6cTZ61UZ
Pgbt+L4Mo7GlDNW0t6HXt0Xv4ynFGoKySXiaAADrzZBEO3ztHztumy/HQnLIC3yESqPj4RcbLfEE
JCXYht7fDZo7a5Sg5HJCkDLeHX5k0kR2/f+k5tdvzUrLsfUDb51yCYccHxMD/k1uAU/B/47D9NGr
0JcRPuH29sQiuve59H3dcC+JmXaH87n/D/+6GMkkxmUJbceKivoEQFZKQDyTqFHnC5T/jIDgaohG
wuTzGefEMcxQvKuru13DXeiA+5ZP4lCpX8hZJwp0w7UPlG0Ik6rraklYpIJng6FLgqY3Z6KlXcFA
CnvZYi9C0zLGn1PmiQjQ7jLxwuc2wFDOO0EeeezHJQEghNGcsyl1bPPbDlLjBB5g04YY8KStkeD/
nwRuYWFFQbQQCpLL+2MAbOFH1vqZ1OzHsMH4y0djXF+HPnPH/EjI/opZwRcaadN9oqv8WQMVlPhS
82W+JKEeoz3bEmz1WllJCxxHXWAaMmxTazsASsxbxQ1Wwp4+rusnLPISmp63cnz+YVnPAZrBpYeJ
j2oyp9VZRS3w0qUFXS6GpFEYFbrMkWFXyBY57LnxKCqjMAMssIGZBc5cJRLzmKFaiNm87y1Y7o8B
5yfwZ0YBf/iF94QfM2AwWX+FtyNMhYeiu4GRtPxx0L18IFGO+jrr6x8CVcgp/vPYTRjTMyx4yCg8
CXPPNOcD8QrIDZDGTjHZiL68osNaCVVDB04C8Ix8JT0a8iamZVDfGaNJ5Xru2xblsbOtcwtNOQo6
y/UsypTxjPEdYLOuFlx1DAT1t9o+s4O7veCScEkljbMVU9IaOP9ix164fQTYRzrM9TeHmlnf/hUE
YG3x5p48Rf875vt5pr2nhsEvgzsrY1ISBv5+/QcxYxBHhY7sqGUxHHUHV+xMpU3ZTZ9YiF2UmvU3
NBiroSgZZZsINsQLlYB06x/BHWFGPSNGpldnDq5Ma7qblPJCM3HnYhNPwkZvi8zzJZ6kDX2mSHo9
sUYDEYMF6/yWFjQsv9P5+RZNc1ZccEyNj8JTPbMs/EYZ4iaWMdnvNOCvZvdSCvb2Xit0kEsmIE/3
Xj8Mau9M6MdfwOPcaleQ4S3FTOv8k6AThkzP14+SJzQqk4VzxwDZlhHy88GY/IKqJyrz5VHathcQ
AO41OVZ+OiUyL3WtFn3+4oLUnY28JqGf+uGP2O5pNQu2bs+tZYZ/1YajZy8uc2mrS2A5WY07rzal
8EZAyqvEbpSDUCu3tKCzVCb5BCGycd2BauK9orB1dUWOzZwtf2tjdet1UqaPfcLeciRM+o7FnIqi
ruhlVKxxM65MsLogVWaD5mr7U5S+tb2w4XXQtMobLQ5Sglt73VAOvL7ZohD3suR/AAZfO9n12ke8
gEYITROmhCDto+H1ZIBXkuAuqJtFADqmfy3mjLPnVbFXjK52eCTBn+7YFwSa3jMCNOY9nrNzyh8J
HNZAxZry5kexQjkBmPkdpGbsdu9NZ3bOKNXWn2uryH9tOP4JKVYwJisgoLN0PKGHDW+CiYGV+UVT
U+F5L8i9jhuybi7voeJKUxR2gRv8ucBOeDb1rnKaEg89+XvieP0b3FSX9WtDCajYy1VRY55gEIeR
0Aw+QCEdf8gdCmS7QeQNDr6RZihRMEV+U2AVXoNKKeADEHotsAXWOb5RK0Gf4GBuIUSGjm4SagXB
H3hJRpj6bH+NnT8T5+gbkt1NfDa9d0KmDjj5hdL37A4ZSqkuJArX0EQsQAbSH1AoopFow7WMsMKO
tOrs0MzW08VHyzsQIIhIyfDgvpFsc3qMEW4P/h12hCO/fBs/545ziDZ6wQJLQpfYP+fczA2aU/KX
FeNfSwCDEb+hcBMJvt2sxKwT84+p1PlFsGM/vBh9Ac0Lh6BU8EzIjDIxbPah1iLkHC56fEtOsp6S
IoDO7gROESh0FWvdrOd/psk61xeNuNr4aNJizrqdggOEGLjqLUxYr+b3gVhwBrG/e0KFJqM8cWsM
Wz5NCYqkspYkle/Tjt48Y1M6zWGQ96YU4r4xzEUzdlNG3Lk0E+sJpZZFvIZgrE7Xuujd3hvH3LvK
RreFalEBA4OFCqWcdo9196yg0it6BOGEJZMHt7dzYY3m6VMM6c1+UUmPpAY7esMwD+BH/TuoooPT
zklDrZtT+JBzfcejz7HS9LA5X/KMSYuLOpPG4qI+pYBx0E1BAzwyvgyMOZUXJ7nO+o3AytML2nER
JIZGxVEDDeJzKSNVD1l03ad/Dsols0+EDSSHxfa2HXDpr7NbZ5qrY1mWbiyulL+KWJC3ZbKznwEX
JDSUZdXvR40ZcZfUcT+FJgfNVbFKzlM9h3/W37CHs8ABtYXSmy2idUDVXrM19kLH4omtXizj1tv7
0sSlJdSh2BbnljBkZFOjedks2unUsQwiSFNzZIilD8+M3aLpjPBVMyCCIFn3MwKeQWSESJlLdBBq
IEaQY4M9ScKqhv5p01bl1tm9zXdy4ssVftTwmvMmsZJFrazLixE/Zumb8mOfBSn2YmccJqxfV9cx
W+cXNV0ZiKWUNGY37X5lNWLdkVzWDme2lobj7u8XNKlz0+n1dEXQA1ur8yN+W8K+zshD8C7xmntF
p5DVzY7YAeITEhDHDyGNxg8MGg10P5B03YSLFIs8s9uES8QVz+y4BNWFnhPM15piOuF51IpJD+mK
Fa/g55V7jawVGqhN4UucToo36wd9wqQW3p6J6C/M2kjjRKsif4bzFkFoAV5+IpARYoldIW6WWx9s
BWSipBKoj/x5iB6z7MVm7x7TMjvYhPgBRoK3ih5Gib+IU21Jlo5/r0TGP1yw1sUwyzCn3W6fFxMt
2vK0xP3FItF7BIBLjJGN1M3IMExGlrNqwQwr/y28Z+ZyI+xh8oM6BRLiBVO3Xzl4ccDp8CB8dcWE
7I6zUYpi5F90EbG+uxTf1X7YAO6qTw+6I+IpC1cKPm73499J5ZLQkejiSjv3NGY33SuojhWTMYDq
WOluzQlcZWWtQB3tyXt1iru3JZqqQ19xmhF78OTnj72mlBdG8cebCfsCfRmki5RAqFOESlvBHque
pTVQMx8fjJkT6ejlLE8kZfEKZuQiAHvl31JSBhhIN67SbKL2sYtwHBHyPo0s+KLG5amU9Rk+kurS
S/2qZg6C01oEcEY/uwnqeNDit2E4lDi9OvKO3sEFI9dVoI/zo8dmshiAPnKy/KYS2/Z1O+y52Yg3
lrOJMu/VbjjU8L949KSqopYNpy+lMtJEPY3YFFHxvLuichSCUJwPoW57RKtTuUfKqi1pEePMzy2c
b/Vrnd2KyAgLJu2pXKiteV61SnTEZFqh6TqG54DZLw7G7ULQ5Wco+4kC++2di/qnu68FZZs9xi6C
ZcozGQaRQ0Ww9hbOP8mdUJ25b+G+AbJY2zfgIAC8yMCrqUDLHSlO0GYpB2Dv6rDQuc5/rVgUqnWB
+uCxu76D0gXGtUZRsfcidOeQCmpob1Q0VnI/TWjU++ME6na/3TMzDtQjf5RSFzn/YuLeLOGcjGi2
BxQZskiTtFv9PqqIWOHQeVb6/Nw2Gog0BaCtmaHmvOEV449I/nBP87FkFCXFLk/RST8itYntEXyq
4SeqQA16RzQcnhnkXEl5B6mvUprNxqTuxvds8eye0qZjNulfgxuCNFUdLsKJSIqv9VQSpWOOUj6I
hLWlb+PTIZueI+mUyK74KEx6/DeI1/PNy8PDdoDVxGhRikx5+nbQJKouMlOptkVUzqLL/tcWnoP2
UqDkBq0iqQ9mBIHTv+w3QUZJyNQol1B6wIhGFaSDP9wh88ZZgproAFRhjfucXkkxcPjKdo4jC8TX
9OQseBWobPm/pNvhQIgw24bki3LC7jOFfZu4l4B35l4VZsSY5QaJokMnyg0/wbnwgxNFIKgpELaR
WbEK/NaqW6TA7J+HLyAkW5b871gYHLK39ke0QCrfcJHX2GMMEKlnAlMN3D/9Mg0sX2M2UJ/GLusN
y8Rk/xrLHs6GTMjVzEhp891WH3CjRMiaoW6VqtHrwqjcRI+sCyVZzRcDtb36xi6fPLwYFwHR7GCu
CihtcbePP9jwZrjELfqRHmwDQbPBeDgkURIOC8w/PyDN870nlETEKb1z6M3DCNgKmtTr3U0c+GXP
I7v1nIRPCQ32y8BIxe4CSnUnqQ2js0M1IXXZyM0qvKFLwg/R4R06SeK2FkQnrexT9q/mLsFGpvp9
afyUonNgZLKFC4YytK6P9xvG6Z/YSsFKut1yktibganjTHZFCTo6o8xBeBuXns1wOaHpkhhN+TNf
HzusHOuNjdLNxcXqT0XARwJg2d5fIP0TSMXcA/wzce1Qs+xc1IJz3GcjSD7dCzFo0pHu68cM65oJ
zSqcuo1Y94oDFa7cJABiwPaX/Aasqg9vkfKeLK+jytt7Qrh1YHX0/qaJEtxaokb/IYjxzEYeTMdQ
3FdXae9ekcvyJfLsQd2k5ynzSnugw3qB+5ROLkN/NSQRJf5QkiutJazaKu19BjxzIvbHOk+5CO13
dYPaselgGLmSu65aDavy8bVTqS+y/gwAKU2N4+xFgV93vFT6ReIXhaUWgh7mcdTF1i3ipc/fL/09
/4IfUakeRhBKZzAwBm9RkyzUhkZZHTCsCF7iW5PDJlQhX/QU4Ck/eDGvEi/PEjr1RruY1jZnG8bE
ljTup7pOflS/5AklLIeoim8+9VnYqfZrRHTHzivOjVuw/7LkfLdNnFXiLD0L3eRjvOrLTxSHJhz8
cMFG8+dXnPHPZVoCU4vLaBQ3kQeSJ/O0seAUYM4HKRlKIU8UOp3T6U1kz9sXDP0t8WHSB+jBotpz
aj88VICjkmO6Nc97cZ+lB3HRo2b0PMTa5GYkQTo/uiNI7m9jB+jbbO5aaDfm82lZkeCLesWlZy/D
VBOd3lR/n3QE8OvCxfB2KfwF3Q5u8WEbeonavAzloWrZwAHrHrQOYf1Pencw2cbPGRNa9uv2sAAc
0h52Zxp6VT4f6hX5mhFHE7SWlJaQLO0h5JmsZYtj/wHt5bUZrc1WNNDghbRC7pIotI18OUX8Ec5K
wdSE7Xeayq4zg9DtL8S25zI2x5xAJn1al3ETyEp4sBMwtRqPXy+BM2XuzSFEvuhWUOva0lQMI71N
UkVhr9w/Ibs05AKhd10FNSgwe+fU0yJYzk+0TYwD5ItIbcjm7+pOhKJ+j7clarT7JC+6ceFh1flV
tG/aBTbyjPS2MwMfdcqfIcXsAlG/MFLytHtn5vBWPiOTy2pEc9pR/WRIf8q8tjjdgF1Men1Amglo
nb9//rC4/E99VzbGECe2rtRiP1LgS1J3/gSd/83fLiovq8TsPNLI9H4GJMzhyDS3jTEDbaKEL6oq
zlMMXbjL7eyv5zLJRSQSwXgpZMfeo4KgMmZDVbn7EBZjQWVjkcmO0V6vnU7ik1XPUQDuLJ9EdPv3
pQgCbyB6uv2J3jThnuqOpRsfkzj6Lsuc4VaR5/iXlbCZhv69mSfctWb1HXhYaV+GrOoHDXSvX/Jz
/pcVhbJklCzQ5YC4CNYqszmtrYSI8he4YMkWfirg10nFGJwP0Tm+vqeB9c7nAnkqCNKmEV8dvKdQ
89yltb7A/eu2iwbDVvHB09TrOx4r+vrXwyrW49GQAW4TrdPyEqFIbhGkm98i0CFYTcUCpu8vO2+X
wD7KSgHnCxYz8wJ4F/T1jsHS91MY3ztdg9WGg17eRktZB/QjxrrSQVQ9pGoF03JHDAiQ7rudPgKy
qS/g2RX1NQsN69t+QscTtDO66y7t68PAsj4Lt9CDMlRveOI618bEKmIMRGJqo4usIYybhmEWx5dG
t3zkeBMlcRYMXVmVFiA/f/Tq6VyC9CQBg2wphCDBG7AY8xHA9z4TS7oXnTk5leBqo7Bt93YAjjid
Ejr8li/cETb4wjDyuUJ5B8MRexNeWKpqAGaBu5Y9p4ov5akE2g8ZS9J/WBQevGc1LiFuuKJqcvh6
TlEuNg2WQTC4Z4FNPM9P49Xk4mWm6r/YwdREOV5kIv+PJCfq4lmM0Jh0Nrd/UUs/3U/2veb6ATst
j2owqhdl4fwe5i+BuNRfbPW/UVlvw2NNRcln26qq185EMzzWRy97ftpQsB8QPxDvskD6Meglfn/I
kUgCERK192TEs5is/GdnObGtOvA5pQql2NE3mZ/qagTm9gSggKu4OpdcT9KhuoZUIWWjnTSxvfGj
ce2jdoggIdHjCghcRk1nr3+lYWBIUlOvjiXJUXE3rVzfwL7Ap780IIWlvRB6PKRpdQMXiBEBbS9u
80/1a9tvtL8aPy08RG4CkEbReza74reV5HEJUmeDmC6Gr+MqMC7WTRssvCv0g+R5I1EoHqxDVVLa
KA2Vrbp3V/eYCwYvUY986q11RPcGhX2s4F/dziTW/WWgQSyk4pkY6i8WxHpJxkRjx3eC1PwnBW+v
MQBJOnmgNrT+zR+3KM25ewetWlE9/wY7V7w5CcLxcmmpGaFzgaMfmGtGLKWZX515KB2fgI30AOiw
GBDMWWC99/OnbnGq6u+6eEEY1IM0IvvjuAzoXIl4tghD2lEMTCO3pseyMaQ8lL1ljGWA6JyInD/T
4cyvDqzkH9mAWzfLWzz3U822H+jsqAziO/NXHI0wFRwI2P+f8b1pUdxPvJMcIF3t1kADT6P8y181
UPAATPJuusaSRC2FP58WI391CHH+rWy2cekSjDlnOlC7cbQm45MWk/1hx+JWprSrCHsvqKHkLr8E
LgG3itSgEOPpPlwmWV6VUeVsS3zxk6hgomaXKMFIXv1wORXwYAIodJBdv745YQs8tu1MJnPChn7J
AxXlvFwGhxHBFW8no8mrvH+PTHh6TNEMiKJl13eB4iDMz9Ezb1W3lQS07tAMVEQA1XslwmY4867X
msvsuWH6NYBWz622PewogMFfAU3lrT2Y7l3zySNdJxoiyiswwcr0oX8dRHlv/SUH+ErUvhgNFZvu
t20Oxuxk7nQeVOfl6JgEQ/N65QYaYhy3w2oEKp25H+lGmr7uFJjoxjNUjj6qCP9mHzECbUHwdC3S
+CqguGrSJ7gjRcZ84vtA9lux+Ozbuw27PRvd5bdwOn/77XkBXuC4Qc7dInGMJrINGgbyCBVPw+CI
ke/WOK9/GLxneqqg6mb0w34vLvm4ouN9hema8w4ZCprzy2kWRJBUYuf6w/HkfcA/ok9Y9grT6G/h
Ec0TmhJ4K7F6NE82wf46bjUK+4pWnXFfFtr5L4qi1Vv7VyBLPWKdC40Y4pNlBjhcsI/voStwAj2K
Ccjm4oOXvbYQeI5ylRXVSFnmwvP58JfgRYGYHwESbUox067+UCOO4Njx/6muWdvMMoOdS5DWTP1t
aoZprZDoPVhzBwpHK2ttaUh385f7XMaKhyyCPOhHi2danM1q9LDdPvQcggmoc/WA5dEkg2nKKk2H
h3Q6aeC158+cKhQCzTNdnzpGKOwLiTX6DeweOsMKzbqTcYNP7LAegLVW59y/6bV0VN1C3N19mIYD
kZOTyIjw9mzCuA5yB+dKKWOLEpD2/Vikhc+C5EeZtE5k3BIrtxZjJblqqHW/HUy3dVHnoLCePPbS
h2HwggVrFJ2g7obYhRHbz7OpjTL8poXmM/KxEyw1Wh9eEEJ4bekKmXglJ72tFsPSswzk/C8RxjMr
c+bAqKYjvNrWWXju2gyqU7ppXRp0uSUsvcOdFq21dWDHOneR016AH8MVlQFERnUcYP6uNX0Q5rBK
he9mgmOK8SzjgYDXX4crcDE0A30YQPKSSzJ6b0yAsktx6U9GEKEkXwc5KeNGJ1vfhvHU7M9q4Hrp
X6wsOd+yvnXIFBQbBploONS9X9RNZbi/ZlsaMq2KqAP/113oQfeweZBstx904AnQuPQcYJiUMLSw
6tIqPikH+GwKSlTpkTP/6zK2I1YHC8okxYf6McsA/bMzveGwauDC+gXHeT31D0U1hDjmm4coDBFn
OVKnsmPOZAJLXC27jfUTd8ux9f2ooNpGEbbRdWfHvnOfizjQfN//jPZ+MrGLv07LdjMi8Zg8Wk2h
1hZxYTkr5SbYhEftMokPo0ap0damHTWJ1SFDaOQg6q4gnxTlWjPRcDF0RFQy4wXtO8hWpDOZ1yWj
SYdij6BwOwT8F1kCdInU6NGVb+y4xqmPqyaaX5jDl2Syy7I0mzNN+zCARunrCGxdCH7faxBTmf0W
1s1ksExx7OpaG4GfPJWp8fI/lu/g48voVg4mEj2spxelcljueKLVrHG+Awrqqv79s0L8HIIC+YXb
OrqGHBdeu5ANq97g3QK1aA315wJAAHgWLWp0gyUQmo8VQSX8SOS8TnVy9LTJuzn7naO2gqmhUHd3
oFpLruMnvUwHy8jeOT2+rHCFIgSHTp/a3bmyiuv6JdzYqcAMzk7nnHyM0gNXwK92zdFX3ZNLcm3j
gBojuCIz3QFTs4QIIIa/sjm7kqTY7Zy5/FCHeX+N1iWMKlsn1xPzU8jwfWql5ptd9wWe/xwE+Kgz
R46GKTVG0092BNIl9awoZz0jPp/4NZoGacQLJvzgFitJclVj6nLmpiG0p9YiHqTDldDVJ7pP3gNh
WyEpihzBvYhmZN9x0WoxRQ3l5XdaUauy7j1OzLOr9SfFq//vufSbTBo+jR22nTvAZ15IjorwwUAz
hu0BLRuuRAxOG67pnmYERTjryVE8k3ukUzSwRn7F3XtFlJUHrjJ6cPtB8EbuPeDm3cJuju1uM5Pz
O5d1fp4nKUgL3a++alGgkh5saQdJXOF6YDGIIa9G9fqNrK0MxnYYDSMBOQcGH62Pff229cu92TXA
BaHlx+6xf4InRmRRG65tyqQyPflAeiuVFtVVBO2CKdKkN0nF9gxCicV3caZ0c3/9AbwFQ/qBNwTr
hYVn14Bcvfr77bfs2DC4PBGvYLEQn5RJXK38prauu0xWepU1LYet7w9Jxo/JYnlDKco2WydP5XKw
nvcWftOR2+9bM/6kcjGVWn4KrjV0GGFhSLhjSpnOzwnsOAe4MxTIgHM9mvT29RwsWnIVVTl1ftT6
jjVmpjvQSAmbIvg/GE1fMv0XCf4dUXgWrmoBOo8kheWjnJCzcYcPRrrb6jgAflIpx+Caq9/Bpni6
PDUIXk3tkUyffvrsUrfsIxoBgNl4uRMEwcyFkO5fj8N60zkaUDEwRsxmCyVtUVHHJ9tGM6e1+vwI
TsymfgvrLoNKubWNvQB4jSDqhetHtwT077Se9Me4xuj0w6rz5xdU1TeZk3ry/5BBP5YPpGnK0XBk
GMFWAiPgFwiNyPJPSiuZy3C9wgmN4NooX5e7pfFvwSt+NozPryJRVhRPw6gchurZYy41sRGPSr9V
5q8mUrzPEwZE12RRIUpSjwD9EElbiA+JQZmA7T3FTZR57lDIDexqR2MmxUziIdoruS7BrmuVj/FZ
dUorjklmOWFiT3wH1Q7/8WvpSd1VBugPaGTOJtCIX0Ql7S6aWIap4ZWrdnAMlpMxjS7lFjL1V/oo
BbUpYXRHCdn7XCjKeYi+DcUo/YHyMd+ePF7/gI++73tgXNW6nDFB3bla+j9XjNhze38Cipkn0UXc
96Ep7a79b8cxc3mtFAri0245f1LDlFxf8I62UAy3vUY6ZgIYrni3Xl2yGfeO3Uh+BmssvxuJFveY
tVIFS/TVgVIuRXVNMS2IM00F3O4dEXN1fUyEqg32D16+WQC3u3c/ELeWicT3lxtQ+pBzYiEUm5Rh
iDwSMp2QRG2yGDtM0SnayXL0zMovCdvm9gQp6B8gDqzIzt3JpOg7UgdgZMEZuHwiqaPKrbBNtSLk
3UAf/P+kZTxKwkINM50FkNp++1TZvoRNai31qPxsqOQViULSkad0GuNVyNqb49vdoYm8Z874+lma
1V9xs7fWERNMlAwF3YhXP13xZtKZa7YAsszwzylcwn2XeJBG5B3g+O/7HFd1bhjAwas9rWwjFfbN
Ot+8dvfUGZRuS1WDaNvsq3FBvQf9uPM8IVp3vCB2jF8SN3J1Y8mP3m/BxhoJNP68CcHQ1CCZyh0L
9wHF0jFya+diwK0ltOGKCA2/6z4WPnurB1/anYPDV36I71kaM72aLXZ0iHbYy9nlbWUWui6keUeD
ejRq+QAoeJLq4aYCqtX6I7VqRg/hpOigypooEAAbDvBZ5NeEVivzRWtyGKXO6Wgvez8uppVAzGss
NIBtNtgSU8VZLPM6V6Dd41m+hrmBSgHxQS03Za5Ct9N3QKp+I9+3Pe5hISAJLkMd7D2ZHkrFQIIG
XXfq698H4mTBfndvoYKCUkI0fTsokTuKv2xJqkQ1ixFd/zAKAG/9FRQVeNvcT6B/WckN8AajMBBI
WBrk58PebGj+byw3CMyjSoEw3CCSz3wsnf8JOL9F4iIshc+izQeXx4AMjsjAqrZJYqTN40nuwszi
CB+7MCs2Gb+34W3qsyJ7Le0x69x4RBbbMJt5TL3+A1jtXfjVGmBUV80BDz7E+eAUVU7H3XpkavEm
KX6cBevDPS1DriMiOispO54lFUMcbcPs6vHJafmr0KYD0ykADKVsEpU0LmBfjVNsc6QYXZhoPsEO
IGSSdmx0ZMfzZnp11khppuq4zXYPS61RBKsiPuJ/Iz1y08yV8SIu1skCl/IS9lfG7qckRFORO7Us
ffWlq8N2YCfH+wKCmHEroJJoSs30E9H9YHnQbAdSag1sP8cu7aGp8+0mM7jf33A2O87MX2MRrEHt
YgSFJqU4HDnhUXWG5CvKzp2SBNixIXy48qltTsTp2hKiaVqJmynkGTvnr1LpQRkOePDfaNYu3wnr
hYB8RgGAhGhQtIDPxUbj0dKRWt/pf5kbGWJv7GZA1tsmsDbnOeRMJmMpeQctLdAAJlbi0VgGtng5
T2FK9VVBSvb8B9YJ7DpIQqUt64i8AmmkNMKoBSqpSZrcIfPXZSGKOL7PYoJhTldiKS+8JMvQX9A/
2YuS6M2A8bS1v7/2JxuVudJNDKv27Rl03Z8sSyuPxvun63TjqSsMVYFTJmHew+hQMvLsyZNhspIb
LkHZsDrdV2NE/mQ79OxPVKNXWCFHsHful5EKQ3U0bQP7hOGxsU3sgrC/l33iyCzfG1ceCqD4jZtW
UaquqDav8TkGZ9dsjq8G8nj0+JeAMvsOQMfnQDKw61efdnzAPH2tGn0fkvh2iWyfaEwbG4NvEEir
YpId67hBkh5vQad+A1BpDwHBtqcKAOQbYhwpuvovCAFrXHyMWzhZJYWRz7/UNLgYM14M57pYsh1b
qGnOtncnG9fz0WQo7HHxh7EPQk1kzjGnnBvgNLxmqX01CyPdQYhWWRdF2zGRRU4QMurWBKvKvDDi
AvZu3FnHIiBFUgofuHNqML5RR9DmNc+1wqHnOZ2EC+3dkCwmjP7hiqWgtAziyQ2XdeMQdk2U1lon
aUL5JKFyRKBAYtiLrBbgUMMrP0z0/GChAxH/3DOFW8Q6ePzknzSYd3lrSqMgKJ2p6qfEiI7NTSNN
6VahVchfb+lq2MCbOHXG5HvykAijmCo9d6hW4g09AqZZIqQJWhXQ7gL2PO2cS1rN1uQsX/aPKYNE
SRWscntTX2KMNSXcy6pMJixA/5F/p/SNXlnzKOXczafeXX+2KFVRAQrXMejICfp4qQVM0smJsadA
16mtZtExMyd7/HNcSB8E7GACw2WkX0nCB6iq7ICtlYO8nuHSRHqmKqnQiW8FM9lqr6YU+aS8L0vP
ZF6GQ/GWlQXF9PKhQ07OkSOVjTy9wz+yFqxVlkTA976az5FJLHOGbwHqjMMIIyqrJvi5wRJcildI
0BM/Iu5D7XGBJ5Nb8JioMyfWV3wxVl4pj8/64A1H5e3h8uhWTJMZuIevfYyo7J96zleai4iE8XLz
hHK/sES2gtMgC4x6Gtjbq22WD/BWmLCzkTE1G28uwGPGz2nEZmN3SFLqEVCyEdjHfszP3sQPwTen
1YW+/nScHZ2UUCYFDZv/I3TRDAIZ6AxLBksFRicarXC3VL+tUXvO472tlMwAzU627OpGwU7J4Ny+
Annxv/zcM8UH5CWJ2BVI/XKmcAt7TqlyFXtsIKTWeFvwDUw72uY3RRFENNlH9ZiqxQRmfhZpEQ6F
XpLqIIAnL41ccR8lZjNMqXYMUxT6LlmymTCBRGT+BkIFazuyhwy9RURz3M6f2cSmUBVYNAaW8ArU
4UW3au+R8NZ5vS9LQH2OzkSUeKEpLAQIWO2Em4TZz7CvdHlgbR787hjWuoXW1SiNUgkz0nmDFpz0
EelBwiROxHcBEzAu5EK1Znr0jNY2L805dGExVujp1q/tDSoSAIzi7hiIvitUzoY+ozPV1EBfOOvV
E6hkG6rPheaKk6f128fhlnUzKrYUDBG7Hs+X+evJbluCHrcfx/S/PSkDr5jqD6MnWB+r5SKsMUFP
OKwyK+nBnjaKHwi8F/NBEq4ZQjvL1M1764oMhdjkhhtUCmaYMWg4v4yAOFbjh1G78ZRSvrDa84xe
EXhzZSzdG5K+sLsdNt9Y15IvIV2FIKEdESj17mWfaS/hpfJqnGcdCfPRqnxodiHTQEquGjDvTl9a
m2SzYNxA04orDdhmgHw85bO2UN7QCiMcKwAyesMpkzvq8vfBEF0gXa3TsdeGyUoUha1Zwv9Md/ap
zlrCMFx9d8FJRArEjos7NHexL3GfzGOqITgNneOLQ1h9dqhnqB/BLX7654dWAeZPXr/NrJBCIL0N
vlYm+fdBR9g63MGuzkpNIt//S2ebrqKcw/Lpl6XH2JpVVrSSQf4EdU4ytRbWOt31OPzOmTqfDTUA
HF5mgEvJm4gx4x2FF0zCRvFw30rNP8UDvbogDsEw+NbDrWdofXXKw8TFgblIcMMCqVQkfRHSh8cS
8g8uHdsFjnqpmNNcnrzvsYnfHyU6WJs9eLeqQDgvm8ZDWFiknhQ7UWGfb0DLx9ObEqkh5GwXOn0U
NM61N6tsyUwWUTo66dwKlDC3NtepHzHSuiBY6/C2+x4Vfkr170KCDArktEa37fgvluXdJ1Pbku0+
Jo9PSmW4QhpNqbVXoES41xkRFZ3eNYFiuaiNaRE3Y2tLFuM1ld2J1fmw93Q5tjuXuaOsQh0X+2Ag
DYlyQ77AeYLCqORV66Zdn78edy43jdrrV591GaJPFNWQXWCqJDpbc5bwsKwj8t3xGZjSlA5mvC/i
Tz73TQ/ZBaEoDRHOWFL+cn3lx2KFtzNujWGbe+QbMh+g+IjPmXQ78tDxFtmcd5ui3DeX8KxwIyMb
M6v+CZ4IKiWEb+y/7X2ScNHe1m9Csz+KymT3H1nK6aGGtSW5RBjxqQCwyq5Z9NkyrHgM4AnQpGk4
HX3anVJyySMUr4GaaMUPc8id4hofFfrJJ5mMKwzrL9XjUwN+LO1MkWr0Z5TrX91skv3GhPwK+78c
Iv7Y2z+u39NRxDfIY4omq18lgth7gMAt+a3eqEqWbKcVIgjRlmUnsyiaSYcUsinOF045bgIC/TxD
wVc5JcX8tdKWdy30eYpWfL9l8VRvFDKwQwi/MEc11PquN4PtuEEhv72iKELTnVyg744EdnSobARs
j+0T/+rF82t+KU4afMwcV9jldOvDjDbMUu6xOOxpH5tdpUYBLeq14YLz0jsQ/81Kg0jyIj1/jQr8
YH3FkcHEmTieHNsSHHDYTaJSx6n+rE6Mc+mTGexSW0tJsn7Y15DTHIG+M5ekxrFnPZYpw3TsBhWV
Zx4PB2hEQZyaw2At0sFWyGL/rUG6eZFxo7r2ZuEshz1L/8v5YKEzGCv5D8/lrfqhXnJlb64LDvsJ
OBLZizkTkTU6QIIvW8W0LlQ23Tzd4birLGRppiRE7jnMGqumDXZ4Nx7gIqtdSUKZqa0XRM0L8hZn
eL8EajL6aaVFgf5AzqqvB9YYbhxUxqSlWvotNg/T6W++iXELPGH1NhpnKXf4WPa9tZS2euw7qQ4W
0f6X0ZFHA1c3QWoFTn9DfKoxrsxIhEOtis72BxjwbZ52z0axqaxuylOb154cieS8sodh31YYNtDs
JcG8p65RHbkeBKTg11iXO3/4zjCDRwpr/gAoMq8iDxvwcQB10eMlkFgx95jGFPU3669BsGsXB5W/
8Oy5TfW88QnSn2Rxnj+EkY01+rSOPoOs70o2DwKNZvoIiQsTgRax0bGNmY15x3teHJEHoCUjBGHV
ESO6DEN6xmWQVD8MECp3y0qMaC55FB4Z1WuLLovpZUvuG9so5v6buP1M9o99hVlx8hwrIG/gVcBj
fQziBrCn9qyt0vg7p5VR2U7Ce/m/jBglTmHzX8haJ47kq8X0soEAh0BgHy+AoZ3MmbwRK+lHkEgO
wdtSwv1Fs3OHwZo+1C9QBFTtMPPYYeUlNz3n/O9HuoHRQPbuLs2AppOKTD/ZnkplmYk3XPrClnUi
WU8cLoMG00pIMlgY/G5JHqBqLL0daOC93cg0Tf+f8nbOQ2eWUvY63Y0r/gglPOFq3F4yRdnhbWW+
n4XcjlnFtIY26XfhEJ68CDPy+fQDvYpxe53Gq0vEu5MSs02L+zqvPxH+QaNWd7Pkozu63VySuHXb
vvHJF/056xK0iFD5Kd8MGijL8jmHmPdWmD3Ybh5bft8bpyKxps/rbtI8MZR0nxsyik4wzqohkVQ+
NybDd/tafOLK6xe9uyS+qyAYJct/WfHcw3oPpYZPuD4gtabfQI5ifDqzTML9IyAYACh1BeQUe9CS
44Yr7KYBWKeu+HtJ8Y+No9nfJqIoCACHK9epaWNZfpbiXKI3NbybbT4jXVJ2VUWgmHYfnncDoLn4
e4IO95YiOL5lLJT5ShXBV2KbFR0YWI7s/Pk8PgjeoVWiSW/N+YJseAabOyqV4J/IfuiPPUCqAL+z
PRmuwyuBNjzkNX/MH1wQNdHmyjW7fUVW5GPhwJkBzzd0s0rf7SGUl0gHHFjcD8Iugm7nV87VL6uL
9TRhqy9FWlCP3LpmxyU/wmwIYXYBW9pTyVchNM9ZVvHXE9GMLkfEKNV7PfT3CxI4Dt8HQk94l1/Z
tZ4nYLdQvvJzo7K4mKYVWSuAV+QcIAcM2W++jATvBlD+X6gf/ewCctzjSUzU4G7YUzYtoNq3KbTZ
R5rhI93asoH8EGySjhkBKaJB4Df8JysXCAWIwGfFpKfhJgI3rtz9VCRHNo7i6HzJmJvUXyvgPiJS
md2oxhGu8b7Uo9u8nJkt9WwxlHZUQ0cC/9w66hKg/3tYxb438ZjutiW+NRCemLfM7wOSe4yyyUzu
81o5V/gizy+C/KZRyTS38fehvDpo5sYyb6+OSfdx8zvoNPnjGRx8zkXlu9E9n69pyHni/Bsl558P
m8IkqqTyNLikPnObWgML2TvmjGwuTwvfxxHE9P06gahpGQOAppM58i7OcCYJ1PyAOEHb+A+qvWRH
1PUFc7vBMS687PRnxnBrzgRYyuA8AoMF3Bq4R+EWwEKe4S/AhTnl7dIpu+4+scOdCiuXeNilfdT6
7dzcZL0kZK4PmtwfikSNKJt8WNUD5W34+2P8u0ET69EqXpLtyr5zpLbbqYp7bLCe/GM6zWas5jEb
i+QtfqeS4u2g79xhGkPk8yXHtBALqEPDxwRIPPPN6D5KbLq0+S4r8pTyGkfUXBxiO88AVBwJKrVw
zz4hApF2BlPopsxrHGf4SyA/0xT2PVIsRnKkp2OrrOZHmm3JwCSvxLaVdYctrE1Q9bG/YCmwuuUj
Fb2f4jyfu9M2KdkWZA2Sl1qpoGL+cKx0ws0B81s7TJMRUltx2m9Nyo8bKlU/cTMabC5Y6gePLdMe
xeRGdvZkJfJhFCHHGj0UxZeFckAy8aOLb9+8ZWfcUEpsAmsMRBUyCpchv0TIThbb7FreAuKLvr5R
J2ZMvE8x2yAuh4etyWIp+ZCT6e45AYEogMzYMflrYSvdmeN5C6sphAFz9uc/p5YQX4wWXYojxGso
GQTLUo7IRlkCy+Zr5i/+dfmnDtPjDD9LbqxavSrz3s/hOLVe8XZGs1cYYf4WiSIAuIBJhSV5kEiC
KymFk72CasVmwMSZxv1fUKJrBIvN5GIgcFtiLTM8bfHxzAj8eSPJYoX3fAg/lrR3DO7qiVibuY2c
FrlafySo8A2eoEV6qM7GRFzkcQPcuZch6LPOK52BY8ZxIJXuRBK3EiOIVVSJhaaJUl3eRI/tI+Ii
3cd7wA3sJD6hsel6NW7xTIeyaPmWROxo1YX57YRcaWIxmVMMQlmnPxf8reqsOPzOmT+cfZy+Pz6G
p2/rGDNf3VMAZlNU6Q0aMx/S2kgYRbkwswFyjgKpiBilSvbSrqk90KBKyA0R4H4eZSN0T/TdJv3f
QZiXWy4QghAWFQ0uDKPZF18DmqjCxZ7B348zFhmI1BunWqS8S3wUWqobUqi8li6JEvaQCaCsSOac
fYeFS/HB1rBVj2rSRFRBNqyq8TnkBq3UwqpOP9A26LgHjrZwtKunhgzQbXfKRXwMuAcn6WMYBLem
JRajS2XflZGG/rZIamxpNve6pRUgROn2X9LDZeGM00lolV9UQYBkEFLKsR+GE5pIk9G8wxN8Fef2
ycIgX5DY9pxlI37DWIDEk6NnLeD90KoD9VEWB0y071d9rnbo3MaWu0qovOtz14nVGq+HkqJbBn+V
NmDqvf41nnrfgW6M5gDqw0Ybf8JxoKAarazMYCS4gsNUl5nLId2jsmaB9/orMlueMqRWoWVMUiLt
i/rdqDcTRRW/DfF56aBU0ZbCOBQ8SkPi0Swub8r6P7GFXrbSE+QVtnQpL5ZTz9+jP7IDlCU5f6nx
ldhFDIUXc8ZOMu9WRIQ2Q3ejzuoANHMriynZaEu2OIXeR2GXmfZFLjeg818yY5IQe2Epd4oEZM8L
7PFzHYh18WZOquK4EdOHCIhMqcx2p+WTVYSIM5FEigQJraivgQuykoW6nwpbDhzsoJAZFq+DzJrm
/+QmLSs9y7Q5X/fdEVglLXtZy1EPtscA1AhIjQTsvv8tidTZgnIIt7n5Q0XuKlIJthrImn2YCOGb
lYW1CF0CxoXgsLJHTfIX5GTffCW4ozXkFkTd8eaZnZgAripH2ffd8nsPUzjI+Pg2+hqJDk+7ockt
O/8yUJqxn2eB/pZsdlTVcY6VuRRZ8eup4UMBIwNMiNV1ftYKnwzhSM0hjXsImeos8YPySMgsWbL5
+hCtFFlXKHiBVf1/Zn3jRS0WU5yk8QGjD7V7rxTY06J8aorDEBfX1t30Xpa7BJNN8HV/1sVE3vAM
voGYBQ2ICtindp/JtIBe9rVgfmHnFaYyhX/KyU0jUTH2ZUtfRFD0noOULwOnLBzPc1lAx7RQ8KJD
QhasV66ZmMOQgZVW5Agy3NcYrcTZarQ/gR8GSTj8Pn2KriC6LcbW40FTR+/8tGxxFcI6RcZDF7+q
1zvqJAKw1uYuBG9qQgDSOo/Y4Q9aM0yDz2S4GPv0tTiIgtAiX5+5WDGA2ETxURV59cLwB3CNf8mB
nJizDapNvIDQ46N2tAiBNxA5h6kNOwKKeWu8yBuK4n85WIrHu9ch5RNGpRau02mYKe7GxbSeFvH9
tDlG5OdctJSzMRgko5ws+Ms5R84Jfa6tcb+4ofYsKB30es0F+WGI1OeLomHMjM4WRuLQJN3esvMe
WyuMmDI7+jEhl00vXhJFeBi1SArNXf8NykwvzqV1CLQ0n5OWcYAxEyTFCCutN96FSzXFI1nvZ9eT
vmnyOhIblBBLM/SYxTStgN3USbaKH+cRD4rLsmIs+KYz5NeElwwT38iXd29mwcGR4Tvzer4Yt5AU
5nG+J+4ibaWqeP8Ivs9qMcz1J+4eRWRN8NUcjIOyEq3HELWhM5jtJD/h0tcUQShjF72TkyxykW+C
KhIDmWUL4n87NP2nE4Bs/W2gvt6Vb3KTuYgiXxgYtaba3HhDuRgtc25bmTUT4JPAz9Sv/Mm15SiP
2SZpws5DZottbcgmt+rCTqi4TjZAJ/HAyBIf18GqlDASM0y077x3EOiKfMaxQUxJc1L/YXgum83P
HkrwbiKPrh3d/KE1mSQPDy/XsusjNFLeHYaUK9BaDj4s5OESi2r5D66T0yKcpObjRSn4N25zFyaq
2snyUybGAwajRniPqphtPU88wdwe58EEb7b8vdjH+/xeRIUgVw/EMF2ZlpKVRarYECD45ulq23nx
jfcnQD3ChmW/xJeB/Hjsy8IjTYSfkmp7TD2Fzw16uyHS1Xm3vpE/PiIDuThAMjN76k0qlFClkq/I
iAI46hVaJey/2Jgc29NlD3YR7/kzIThc3T+zpnFxA68u3zTWUJ28V3sJiElKVLGIVCnjKc3lv9RG
GG/7qZG+bDzwSx1nPY4cMJXIOqiTvoduu9om2meD8+VLa277CSQ9eigmErB/QoBfaxT8HDfla0mv
c2qGv+INTgFZPFQM+hFR99NdsRQ5YeSzP4pMrtP3TjfIwXDfbDmTeGMxKVD7G1VAcNYmIp4I8Hd2
1B9w7BO6twtLyv9oyF+dEU/pEu8B1C19PK1hgU5YyzcW/5cutT0QTUqg0JBVUHq3stEWNdfRmqhK
Jhh7fSL7aVFS6sP2TBB6Tc/HgNSQgcKc/qc61UQ52jXLZnG8s2qpXpNRcrmDV+Tbbl5bMzgyzl81
yocXEOOOm5BZXnX6hVDCV0FcveePcLdt7OjNlTWmwveOceOkIvWowJQGBo1/wNfNfedluIN/sK4d
BdF1IjSJ4uGdwKWqzmpsm0rB/4LeD4IjZPgGvBilKsS8abFdimlh0X/ITuBSrtHOTVj7w+yr9P5o
HmTeQ/ZkMWM9LgDai3gbaIqecMhSSgE6aRkmxoRh1en6GYzRqxgJSEz531JV85NWd7QXsjEA+ZGH
x8lVxp3M1uEex+wIs8swV84gdRLOVoXWxfGBl7mSEJ4hUI1Ckx+APKBQMmUoki9ixcloCKGJpQ+m
FRke7p3UaEEbRXBIQWuXv02SRv8OejMf9jmjZza0QYSLtBzUe5/JAo5HlvdAViS8OA5XPdm4WdN4
n9aHY/93NxaxvFGxKH2pIPZAPoiWzFCN7iJvUv0IJIpEy6WotBYkR1rAr5jjCDP372wlIWlseSzI
pB8RitgY74+jjdsvpJQtIdPN9K6DYncVClKUyd+2tP6+UlxwDkuou29OUcgj6donZmRMzVA6pvci
asRFmhxT5dLkjiCXvUvpN6LIlESn9Tf/8A18VLXSO9xnuofi8VYMMzyM4cSut0orQlgapubTdsk4
bTFkyXwxGT3TuQYVomCXpspg6B4lSKBZ0KPmtqXPBpmD8O8LsYAb5L4oO2b3StJcFyy9hsrLeIsG
IXg76sGbgxr+5l8QAdSIipexMwaxYyKV2dyP7dAezIFAv58jGBnA64qxMQMpol9KiUiWTXcx+xa3
73QN6aA8UeqxZkulJHn2n0fLEMrtP/DeMoMjJ4ZPUdpRAUR/dOfz05lGSQrPN2lL4gZzs/qCiqN/
GmUJ/8KmhIakPawABu5VYFAhxilYt51q8er50PJFJni6/hefa37CFHtb5+i84h/PmrPkEPiyNSSF
TUB0fBxk9X0gyoUZpFH6E5AuGUKqcRdqRb6MaVTH937k1gz2dCJiWnGsqAUElKstPOdsZpORxKpT
Aiq4onaTrogdzCC20UdTlmuWf6ctFoZs8yoYQ5o45Tmo8cHVRMpEtRoQXWpbzdZfmiK15nP3cXrX
3oZEbmSgzVCS4eahT2L9WvEyyZffTX7kk9cJ0tXTWaqDj9NlLB1oIXbug7IJDTk4SsnCkWNrW3xw
anfkuLk9I07ZTo+swY/SsCxY7kiZZYkkxyXZbQ66wVQYR01OUi3fRR34q6qV0ecR66+U5SyPzDD6
MzsKgmQLk1e8LcmLl3PcAaymvoKATRusJ3XeSkI3kI66BKtuJbZSA0xhaGJ39bHi8d4lHmE7EEmq
UVF4j9sFm9JrEOC59kg4qgTCX9HjVOFL0CHEDOfnjvXkDjM5lvo6MPvf2IKhuCO4a1jW8KVJmvJO
8w/AIj/JODS6Z9KA6/UUWWIvIXlP53fudRKtLpJLzKSwMLeD2Trn+yi73RLxkCkE79sGnUEI3wG4
PrOCkwPkX5ez6/9TMCxSJ2Pj0amdb6L/VgJaIYtidcVTXsGfwfdre+Vlr9AtkBiEocnPWiEBqMaJ
mdsdOnE+0MJY3n0hzRsfQM61YW1Ji3txp3gSgoH2iC7Jwvd3UUzKyMADc5hWryd5LwcC101szuth
0oBZksWpGYrEd1tGUiQ8ASeE6J4dWw6DxKNxQNEGQjxKUWEbmjLllASv/vfK/VzE2yvKiX57DwMC
XPv5OxmA9ml4BGNmRTAlxPsLvqE2BTs+W9orTaCyQzJ/tbLTt94QlJO34Y/0vLa8dBlS6uLUqb0f
QQDt1yvyNev/TSVeu6nidJQQXJS05ccqtSQGy4mw0i/2xIUrq9w1JTt1D3Ur+5ae+uU6YVrp+6UX
DnxSttDQcNYvJQWBVGPJosh2IHX7LOtKQXaJZ84xsfWcjJ4sQF+/MkIS+RNXE/7jOHXGcDTFHMul
8B3FBd8vIW4DciL4dITM8Z2su84CrHgHQ+q0bI/vhe6Db2aVNwn1y/cvjISK97T/Gsq2TwcC71GU
S7dDB8VTW82fwVJqeDCYU9FS3ieOUL0llxz8BAVsc/LTczLT4++odp7dcV8XkyWWXrG8Zp729U9G
QNLIkZD2/j6fiWXM7OMAK09+yuZ341yzm9vouC5vxjKUvRtfckVgYFTs6tmJy0j5Y8BRWfKPGu4w
ACq7w4MalpDifuZeahZivM8s/+rlErGseyIElPOU7trzDH98eA8j60a8rVk+fKn/j3ZoX9sB46L2
VO4iqu5wr9AMGWBCVQWp9KKDMfZvUhk7GsGjjRpmCivJm5Qz+eURZ6elaS0WtE8kvcoFkoifs/PH
1+qBLdezgoUMa6qXNzVTYj1x4Ah5XKHzAwX8yWdVaQKhSfoSScLL96kJ+KktKC59JPpNHgog/Er/
zVtDkdOJiCN3E1VyxXjuXIgrAqe9rZpYipum+OJSMSDHuP8hAQdRYFNk1qbOWTmF/s4p51CvpBRh
1O6hbCea+j7NNNDBROvPhaawaMKVjT9l6DAQR+ir2a0FJSSn38/N+FeOA6uvM1scKwGAzWi2P+wt
O9zmyCcLEpd+rPTSEMVn07Mmd3SqkQYhYy/cGsfJrk9MDnmN5g0mQ/75YlrbBNvccrvWfNpUO33a
vrP5ErN+sq+PYFozhAnPog1FXR7+BDkv6sqh/ov3VE7w9HWH8V2BT+Qowi4uQlAExz2RLhOD1kbz
a93MDmH/7umtdaFPA6XcdlQ+MXKcnZRbj3mzpFD8yJCO7327bkHmU3z1+0HSwfc5TdN5yhDsFeeV
dPNcZ1E8FACMFsfTziAPGwcqWXkOCrfeBi8yO+GcLeBOEzWAQ2XsBOr78vNQy4HIRhNg7rUIsNLm
2ZXXpYiknSfUVEaCYN25Q7TlAV6su1bBLwsEtT69SSUb0Ph5hsD9wsI0bM65jELMwpo8HzFP4rR7
5Vf3+ymSmGpskEenwcELmUZJwv0tdIP45s8SumA4jSHwyuM57nRbLR5OLbKyeUcNGRz9YDgBQrxB
CHDULy5uTjEGeyBDy7qt0CvYhGFSiRKsg8mqddQnlscgC2cUWReAFg8OjD7cZdCIqJNYnQviUhB0
7/lIb36ev+kCs3qB28JbAboi/RwMWpcTG4vYr8VWnknCYClOc73Sx+U+7R6UIMGWJ9pUnhpYQs0K
FedyqeIrG9Yax6Nd6bpYWdEgYe1iykq7WgPFOVlOZn8W9+WPkVoLLGdSw3ElKnS7MaNdHAtkf5wL
DNuf1qRSGXT8Ffu2ntw54NDrOFn9jG+GdTRvZYunKlYceVM6vVuN014WbbinwlXQ2GXm0riPmOp7
L9X2A4RrJ3tXO3zRKvBfAl6MW/HSmUYXUOHhIvWfkTyhR92Fib81GKsKPF1AlPsajR1v1oiEks5D
rdWai4VnDmSDVfPvRFSqHBocbvvxVfQ8WlcvS+gFrNgEJWuciEPxuPWHumOXrHOhum48p5dI2pln
apuAwAWYmRAeYDazk+39tY+3YMWlhAT1Nqnd2hju37x/Z5NCUl13AUYKW7mLQ0zF7H8DZOOXLGTE
9VzkFBT/kADaoKLY5cKIwhhtGQPthAGT8V9aq3I1sqEPNlSxH7k6T/sX5YJgIUQB8L4XNBj79vo8
F5hmE8GSD5R92Kh5LENQhpy0tTHFs14IbIG/hSbt60J+WAWuoXjraWNDUrNCABF9OVV+71LnsD7u
8XFQltY50Y3lewXf2p2olnmc/F4Kgqu9F1gvTtayXcAWnEcK3g0k/D1o3fB6HLAwuXJ1Q4k+CPd6
slQPY9vK25ziqpl/pJMQHCaxBDS2u9y1Vhrf9taOPNiSXZDacgV232az3tpZUD/25xESXlmAG+bZ
CZRVUWmNEy0aDFyB5Tk6z5qb/zZ5YJR9wV4SA3uxXqbv+5a9rXhivortx25cbzdEaYsSiKD6cbpO
jxJN8ZyFmAyg828SJkBCaanDCazhLLVfGaVFDLaz3K1yKMGW/AqhQmzzj8JhlbJmRfqzAUfCGSA4
uKgXHah/cV9dq9X/mm/9VGqXXq6fAGUE/gpPPw3bScumqnW32KavaDuKxDvcYvujjpro/ClNUYbo
HPGDSwvkx/R90QpQ+aTrZrDhpbCtf/4pX9ASeSJppjbUf07HFNPRtIiHVgJ43V5jbKZuCNBr0f2y
c1K+6bBOuuotECdOPnubwxegKrYB9TJKmVQDHhl30mu6wBYF069JQ702TutbWELEK19Cje2sZxWo
HldI6/IxhEcBA1uxn7CiOblPCTEe9dbTWgmHXWhLbh/iC+S8INPjs6G8Ji/UFm6hpaXKRIHvkS+N
MbyEu9AvKIBE+bCi4WrOeNzRW9nAz19zHDA13+GgSFO5g6WBVD8F6TghBa/Qn5J+dS8+5SU6Lr+D
G32tvhxxZn8gtka5zC7HPmf/9P/xKs4LtSgixSj/xSxiPOaSHhXg9gXaTAyWiIuOxgjumxq3AJGl
PLoj4vHE+ZnbHfVF4zP/hYuQjoTEU70qTd2cNVZb5huurfORfe7JJ/86kvqj/g29+0W+OHpKiXhA
ut40A6bBmyn55k1/sH2445lZSewmE1d0mM9vZMmZXlq7uKic+fbo+HWSCf/FqP3iLbtT9AK245Yk
tH+BIzXDOCxHDPrar5vSDByWYim0joFYBoLK3SJjsUvW4F9T7+pbFRvdlaKkEDB1Z0RZvbqrYevI
+mG1XhzpmRbLJjNP6U/yjvj9Kx8kc9xhbWViuS9/99UIGQvndEe3RKkMeFmnfilwpd2WDZNchJ+a
ByKAlrwGeVoYr5l0yWIMTOOEssMUVJWha4sUj7hsIk3Xkr5fWoU8IyYN1t6A/jeEeqrp36uJ1Z/e
OGUJPn9MkFd00My19G2nETM5Jn8mFSWNvFrDBSGpX7JBluhgVsaFENw9RJlUXoIW5u6UVyvXfcvE
wsRLsGw87oPE2al6F5yzCb1j5j+9oU1+EILIN6w20VSEb5+jEpeLvHha2NB1Ni4z7czqevczQTfa
Ik4bBpBOyCuO+3Ud1fAR+Rg2aVtd5UjwrZ0/DULh4Pnp2YrG7ABj1VqZglF4O3TyXxcqDxmaiPpm
uqJgI1eCeWPHvqGx71E8Z5Nf1uRO2N+UigroDTnTsukPI9xGAT5al6mivV32LqvnuGvdlIeG3LR6
3fXOVa7BeoNKfKZWP8jJJhE2mcZsUBbxm1ihj2mxlfMoiFtraMdRia0hU5gq/xhIUHVBqZ44yu1C
sn40h+qagf0QygCPk7faOZtySvjxmhQfPbDDj36tFHajvvwazp+Ygyt8NFMN6YrIOT/bvh3H0VeJ
UXicLF4dUngjxlR4QrcwQ9cgoIBtaC6ZdaoUqOG+Lmihvx1RvoV0enKWyI23z3+OMGoRsyC02Npy
JG4lDdjzZZh61jSBynrsD0SdDwzeNtddUv/teFbpHxQCAqaTNGYqLqKYblCOwePS796f90rS4h6T
qGwhkFKYMhYWQaLom9rIAKt1Igmt8ulE9Fa1pkJZEbX84XRARppsSoQ2T9P7XRAnZXY+LR/UAxZ3
noQfu3nGSPSBLYkX1HrlNP7Xbc1FeRG3i3WOifP/23vzhyiOrSt0BtzNJv8bwhKoze0JzWp5LhXd
AaLCKkyMyOaHU/JJu8S2pVl+Bp4TamNkbGB9fXQM/wiR0M15fFMepY76m3vtmJ8JkJaVNkUzARuX
zOlntTDFEVwStmAaiPbMhQ5OYhWqEvwlokHNVaaVf0whpWFWNcWxwtOGfAFNaLcCssslOd9Qix6k
GaiRM30546RRVh+YxZw0f9ZWChSNCG/sbnfUL7Zn7SxECnMR3aees0pGxCB8DIOe0mxKYdWBHCho
ZIVG30c63g9QmbZ7KPSrJiD5475ZzVJ3Ww/MEV2etU1o9O9yTERyo35fsDmz79RaQRG3ZmLDjdsh
EhOpcjGoJGf9o1wEsUkCaJaSiIkMFlquZ438w6giClSnHMkgrVoa2y6uzNEgZXaPk3hSFkHWHNOk
rdJaE8n3x353af4E3MtKGYfTSKKHysZEQMexbMdnfvQm2bpuPucgYQLWuZSywW/xJKrfL0bgT27q
0fPa24aNxNcUT7YG0cU+UDuG5HiEZu5GQLw5lmPfaBIWIm5rl7/Cwcs+RCEuqdlgVianiuVP08Em
4V3IwRDyecM7+Li/P/8V2dYTfZq2gYaqd5Gp6kfwPCPlCF3kUMKwOXwRrhSQ6q43tEERa+4Es2vc
MM14AqmNiEW5wnaNXpfGbsOOeFBChyRHU7yV3rrufzbC5JJjSRU2Ijuur/K/8YS6G6/59sVBTeFn
wTyO2WPDLLxlbUejdXymre3L+qdM98voAaD/Stb1PEJW2Pxg4iHZcR1X2gWR1yF3pzoVj2SCQ+Kv
2d01S92bexL6JWvaBTqHOl8B/8neAzpaePJ/mhdLs456iH465norscQwNp8EPNMMmL4aCD/prdXB
TlF5jL6cjb+1nxjYh2hges4Y7hHPcRiJpWj/31TNYac9LiSbHLwMeXyX9ur3eaZh8tme89VqLkcI
i4zkF+MI6yMSJpKlWkyLTkgGjbo2u60mZ0YZn04hpFC1oMlHxs2WLZTlaPdvHxh0l0srrzvdf1Ex
3sKTBBAExPvz0avEWZWggZzaWoOIMmSEfIbE4znWFHZjFW9QgfTZM5CXoJdB1mpK9NFzfgXlv+qJ
uXuaKT84Ld4MuYOB8GU0CdDPq4Vi64k5Lv76bR0kW91V4OZ5XF71vzyIFHUthx3Jk3C4F5hwBxfu
M7/2FCEceAvlPGFEO089rEeriXW1ptWrrOm2a1P6N3CG8MsuboskZXDdJBMLhGKwEyHTlynEtNqb
qTvN+xasN5Ae9PYaur1PYxROdZQ3OpBoBVoVw9x0XP/lWmG6MIJsiYek9vVL6vNZoFnUf+jN34Wu
SnJG+wkV8hgVoTYtxgJa41W/KHlrpm0L9Zlka+9aJ9FhtSEsJzDb1lRbKeWgJPngKgZCrXdbIu18
lqNaxXjyGNoE5ymqzGYzmlr/Up2LE2twMPvK1MoFDFz2O1qUdT9/6qMr2MVjpGKDkGkuWeaNvwDG
+xu4VUivPEpxGt7xm8L28Sz4t1FCArRe4wx6G0mqPrNemdmSPVVoI9DFZ8z+ANJlETXyqsTK+HGm
BnBCf11reEhNc9SMKjnuAxEF7amDfIzpbh/cQUhaMs3nB/b3ia0JlYEOIar0LstFSILKcmykAyFa
rN7Pr7DMHmoB6JhLxXJqV90TUVlqAiyTgqmNlKZI4BXX9MmJCa+2A8H3TkkRhbwk+WdAXOnSIy2I
usqQGPof0gyMGwKgKZaSAPIyWpHrrCe2B9VrKFzqqmwMUYcHLxWqId3CyHnC6evrJ96FVE197TS5
sJRHgcOYOlz7vXbHFjXoadVunIAnnM2r7g81X7S+NpyNly3KANmIYIDlmkmj5olTVH6j++iHY8pp
bIqSLUiqxWy2QWhCS6THL8v/We9nSq/GjKNARv1aZGmBOnNXDE5OkH/YWMTskcdgs/y/w6o7jnYK
ijz8pnUFEpUj4z0fvMv8Qz/pRXo6XgVvQsOPx4c4uVXmxnh060TReZu6yuDs3AASnkyOqcWkVEqf
vLHUbZn2XiEMk3qGrj7oev36bBdGT43ebrSjzCuBO5ghxzSX19+9smeceXt26KFuvje+vWo7Ndc7
0OHh03wqM7XMR9vDa5EE5yZCEg==
`protect end_protected

