

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
esuuckrrKLBFMMgSrVud2ZnB0pvEqrOMx6GkXz4dnPp4yshTD6+Y2glVVVlxat4oj6oLNAI0JrQK
DY/z82hivg==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
d/1Syr0Yfz0kK4aSXCIN7lq+kUu10RASco8trwm0ImfJURxtGkX5KSPC9Owus8m9ZNLVa+4W1mNi
DPA1z5v28araMT+WQkx+2smTTBb95QnM1r7IY8WLJwhz/4br130YtPfh6ALhwuPZLGS7lh5+ZNqa
WUkp+2aPy+o7nP5Neek=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
EghETPBi398ucn66loN/344Jtlwrx7OhFAMdZLO3Gvsf81gd+y/lO92JbZIwpE5sZICUxsNH54dw
q7y/XtZVcW81UXDzCet7Fnd81N7WGIqo0pJecDfSTWB8jEEqdLB/p9QS5cVBozkWw9ZXd157NWH2
fYI6wtb4DiMK+3xbswRz9tjt4QpCCW6pl02xp3h0AjoDyHQfQiHlsbTSjlklPmKa/t4Bvl+J2OsC
lbC5D/MuvEAoTUQ7SK30lNJDTITWXb0RGcdN8tf/1AbxeMFGNs+DvhkJcoBe11Q4yCS9vXGZYmJD
ooCuGIJ149GuhA9Ebc3S+zqtQIqgB+Ip/rSAVg==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
XB7G1kS71wIOs+JCFd2Cvu1TIPgCW+AVgVRokt3aIVEjyzOaNQpUv0JxfFRbYs7j+wNszYGSy/VO
ucUpEKb3V/Eh6Je+1SiQK8VPkEGyi6kMKodRtbbO1t51Edv2l3Df96scmfDCuwUmCLxAYCnMI34o
GJA4Te4oMZLzNzksU0M=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
mYbz74Wd6t4yNkXqEEqIyqTMYr1gDkxJuJW5Rg5GXWUomZKn1t4qMArQDnPwJx4y9XZOu6/MtCnL
fPfEaeJGNkk3xubUfcA48NrBjUlfoqpqaC5sVaDR10h1kTeB38B7pV1iwRz53qngpcQ/++tRqM1Q
t9nxWednDhGT13iznArEKq20RLCcpL20e+RRoIbTe3wwmYnDWI+ysKyhOx1k2FPgh9jb+4RZZgn7
7PDivXP/gbNxEf8PXBmODTX7OG6mMJYh9DN9gjuP32wcsw58ZKTKhK7ryO26lHYq65/5CZ6bVTRf
+77RaLVhpZ+Bo23bR+0rH2ulVAt4vAhPt51hRA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 26704)
`protect data_block
ywom79kuvapiyj03lybLoBXnsT/9JsKRHp6pGgEQD9v3VrWQPnn9GgU/3QdxRskoFPwVvbMhm5ty
twsEOkTdP6osFwurfLMEquupq9rZ6L7hYf4ALn9cWgNaSTB77CtXi5fnXsul0ts7Z6YkDhVCIocK
WCi+o/mgLje1DkDQ925WKIPZ+aR244S8wHQdxOnM39taBp6Owy4yPTOGoBzFArNstxUPSyaT3yGX
ndhpzGP2OJ9Na6ImPLTzlLueZftfwe0zKclki1w5y9G8qYoO2gTymYy3qtYGjTA1Bg9pG/CNN8Ch
jgMRNHjdGjD5fCcXkxOzzPfIHM0hMtgrTp8OAFhhjy5kCDfsAno/e/ALW319goxIGt2tIm7YjoCr
eC4y4Pv1r1Wzf0xkwpkJgKLJip12L5E7XcTIuLQUIMwNC+IDlvKDJEsYDIxWcgDTOOCgFIdoqsZn
n3EiCRE8F9vDnkgc00y+hCI6HMOVoRPt4Z0wxOMmdoeXfa5BTKMuS1xpLs3mytghxQX8wbqiMwN8
kyb3njCXmhg1gHpBifRDY6y0YAFYtDy5IvmDhvMR8HXn826FkHrS8V4kY1CHZCpdaonxy8ftU/h6
lJafry0mIC2uKoHCHzzB4byZj8X5Oq7UEJ3AcSuZZd/YCXPe1n6xE7RBuFqk2icppMRw+QtICl1R
5031N1rVBpIuq2hY6wAuxtHES6cEBubVzBpDJkroIPD0FIJkO6vyg09RzML0XFJ66ZVSyRL8Uch3
qSXctScOLa6GgbXxyofC51d+OMqIvtYp1sfk0FtOpDK/vUt6lMOtSgYIu3IHcdwoPgVI5JYrXkAG
LNyJxy7AlqXH4v4/j0prlnOi+KOBKd2m7HrRB1tfvIvmHVcUURkf8ZUl/eXlr/eHWqAV6sxV8QfV
KBJ3NBw0y6hJjfb5jRpNAgeuu3G7NYa4YU3OaGw5IoDtm7dg8JPIMYZ1D1UnCMpp+D8/9uqnEAvP
QbVYMi/p8tAkpw9Y94CSk7wvqSLCYmm/C42nTtG4PHCzIks87SXynHImwOfHwnDXM9qvfzRHxn0k
EGIY6SXZhkEDGI/8og4z3T270eArM/ZpNZmH+juxzyM9WAt2bHnqe5rbpS8bJYu6iOn62C7N2hnV
P71qy7jRyvE7mjFeJSSepX7n4d7tv2pnooK+2QGlf5VJHqTtHgTANswItebqMTMVBJv4eXmH+cx5
ILwglsD2YlfMuxyyn7SAcd1fQWMvtr5V4D0eGKCSMnq3cdw9HXrsyIvYegti0O4l+1im+lNLjd2d
siwsFjW0DE027XTeLaSMS5A38dWXPD1dDPgxmUTH2rPNYGv7RCkMOGguZJ5i0MpyWregVvooNrvE
NDUZVmlv/IGbLPTcUKn160z3PQ6JapdIdAZcs279X3Roc50Ks9oQJ4O95RKr1UIxIUvibn5vy1L5
44ZqoUVA47XkuC3NYrDSpBrvnp7i6hEWqEGzKOnsEFIMO1DdK1ROGsXVp+likedNcrG/h0Kavsvs
+dOsxHyw2XIcGiCmMVsDDjCqEgE7HmNK0aRYx2By+6aOaAOtH00mmsKaWcd/QCmiTwWAUfHMRO6e
H2JuHoqPNDKgW+yY9wNIIkYpEj9pcJxAZ+ekNV6zNLzwlfRdGzdpZ2/fFLriAMfwTe2r6Grz/fJW
Kz2uE7gJ48upuAusESVq1T6jtJhUtd8SRNGxJVprDq27rZNNHuwVF4jAYrXYbmzJmX0HKZFoYtH3
1vc8aXJn7mrdHywA4BO0/KnSNGNbLCRcKUyNbZ3pgZd88i6//q+1mSEdTKvt7twtgVqkKT2BMDJs
SguGEX6yIzKqcvDEJXnGZ8xX/wPYH1o4tVqLMhXNk9ee6Qk/s7vtFkuW9+CuqAUewFWELds8iJKo
R1tATXlSZH/D1+mGQtKlFLohSAQcaN65qJ8lElAZDyPF3Xn8bXMcxOBoKiKMSmiFbZqJl7dibchT
kOdFJKRnuWyjdHU0AC8RvRwsxecKwaDxlpGZ9OrzHbFbT5nMZyVRR3O22NM1k2yHmeN51lY76sYH
rxziQt9Gpps6+3f3qK+0VuffmtlfO2XM4hBLK7OEBItjaIwQEjlAT4XJX8Sdvt4S1xo3AYKvMuod
pqhs1a/NFxOmq4ZCV2nRwZnvQzGIpRn3MmsqN44Tz1V1grN6tMWXoaaIifNypn1QrJsgc6KlcraV
WD6t8nmplymFKgLVc00pcTDhosVbonbAZjDg2gHIkCN1lJmcp+RC1sE3uy3TOyFE6q/Iyoy+4YrA
SBaz6tvvK8hFZxUUkA1TSrjfqUNujSC/mO/Ct8aTQ067QcUXqNfsnYOkSRMqPSv6KFThX0lPG9Cv
+f88MduCUgnCyMIAdCfvlMkbfcdHVSGHuLMhZmAJYq20Ib/gkpVYqz/SnMPZ15aAyEsod1NwF2p3
frBQvAp87dzT7OWWKaSdIAwjlkBv3Qz34kYM9NnZooA1NJtkjGYmEDGZiGtMnRnxFpKWc9nQ6mLt
TcbmlWB0KfgVkxe+cpUeZ+04t99aQ8stti1qXUfQ2PJqYsu/FvmU0te16+M7gjELoEoEjRU9te9g
dU2gpol1u9FM2UY2LUmbRjgQHocsy8uRwUzBDNIqhGQQwRNKlVzHS4DLUTOdabxVdv3nsktS00LP
Q14V977j9oc4rPqoTB3UiEk+lewU2LBPQcALGFCRAmzq2DbRgA7Q/Jdwjjbyp5FniX71WTQjd4PU
ZeUqAzfc/WqBaEiNeKev+Zeu36pKQYNGT7KgyE3hURidkixTLFxnMgqMO+wQayAhUZvp8PEDq3fZ
zUYwzPvJyYbnC8XVrjnTXQ6PfChu3E29+SYxIic3mZuNLBPtztp5Y8ZpqHrJAkHsgjd6XZfSTDfC
OkE6omMzVJc6GdAlC4XYr1hi0Euv7bCvJNfYBdngBOE69vA8Hn4CYYzA7RkGCjkb8MfjM2zmlplJ
+TGBM+O1Rudb4KQPqMYWEcSgOnRlJYpD+O9XcMRr+sR1jVXcqm21hTfhHHD3qhA4xipCTqA2UUq5
VUywmIlBWVs3qHqiEAWZnKhJowDA/vDau4DMy5VGf0k7I7fIgz9yZs8sJbxvlcGa1VI1a0FhuhEe
hBwdUJN3Qr1PXMwIXv4+3Fc8Nn/hXkX219lzg6olaDlrHe0rPY5n8sOGGHi1mniQdJskjoSR6mQ8
xpFFIOBzoQrUVT7raFzgbjGFVFFtXim4y0V0696sp6M/gMUaDCo+0Gw1n4v+dTjb933Oqz7B0hSn
EuaL6bGjlPVV+AKbCLGzOeSYWZ4bOapA1WXi4SJcXlluZkkrntH/7Z86gwOeMw7GE9FgGIvkxZtx
r2b5hDuZKV1k/kG5npyRmilkrUEpTqO8K77MKdXTaEouwpWai24T2T6nctd0yf/bLMVc5QapRqDd
5qmKV73vrm0lVxDiIfz1D10Y32WWJkHGlMT/pyIQ0oCoIIDPYdk80PFSkTjMSDZ+9eLMFzhplPBk
oFLZZbu4jNk5Mk9TIgyhEo8zi+Nk3RuKbH7U7KRl9b1diqCBIQQTSrn/5ILoHlt0IZWbOnbyjHuu
xwSgAkyfBbKvbXPnwnYbdu/Q+Dk73PekaFhYJ0k5JqCELuHQ77fqbuK42U73xmGv82Y79BguLOPt
HQ2bT1oN9MrhFlg4/ysFc3CcIykI0eINmml2XmLJYz01eUTxZm75+dMU4YZ4XnZm92LiiyDfbyYL
/W7Ni8wAek0YPrfPdZiHUqWhXEydVXCxkU584BL9brbXmzjQVvApZQm9hAHN82vUB5jcPjj9UM35
Z3RxfDOLcYo6pWn3wW7uGDv2wKlynAjVBPcZtC9w45RTffnStOhclHS6ulGvwZPWUM74t8yubc+H
2vcYHo1ogXHd9SvTekQ7b1gIV0bom3qX+05ulNAjUPyW6hDVCgYsxcIbafJZKIS9RAKsF1TfVas7
99qHPZ9PHNrCrfY4itEDlb2PDOdH/2r+xoPawdnusYS9DRhnpaYsZf47zD7TVdv+zHPRg7x8gkgA
3VPPXBd8wmlnJoL+OP2QDvtvT49rwN3x+u2Nq8G/MGcTp+Qg29xnYmdurRhQgUmReyslAfFwv4YB
XgTJxkuvAyKD2BOMTfwXi3NaXVk2bM9D241xfH2k6vA1io/+JJ6OQGbHawV17frr+Fo5RIikFy4A
swsAa4XiERF58bdaoNgETIai34VpHFL5bKliw7K81Nr6fEg+lFdaoXBo1bC+VSXivPYLM7/QJ724
NCEmFnHRgErqHHJYPcji/y9bSNwzE/5L/00RZqFaac0xE+o7aWMO6H6bqZ10hJbpA2qNRLpZWT+p
9FGaWCSBRke5iUyx7Ysff3kKtpP6uMCpTz+5XRDuBjx6GuMhfytPLARPFpWofpHsrpcSdVoN8pYh
1HzRRhdYH++HjOlTS0xKGCF0gBgAQPBZdqmh6XmkwlmGVVQbo8nyD7vhv9gC46Kx9leebfpRbUWW
1nzlCy6S84wNpWsfJx0/Tgq5j/gDGm+wYm0edEoW/ExRzrMC5KB9jmCjyM6+Lq78dvJ30Nl30Of0
cbFGyXn/MwHxzPgmTq2BYaZzmZIy5IbW4QmL6n//u/G8sVX4L6AbW7/IPjGgOy/pEMIMK63JIkWd
wjOx0ZwdS5s1pZLulrYu7b7qrUK9uBdQWCGEMbjgw0vcxCZxMfWNYPTxmr2m81rAUKFZbO+KpzY/
FOEBpWSjMMpOWrBJyNZC6R5yKDpQvc9EeRqZ1LK17MbdAhWuuD57kL9nyQSvcOX1Nj9IODU3IpWC
OZlUQK70B1UGXiAhx4p6QI/hDOHJcaNc4hyhzx3HggiszI0quxIDk63+x1dgZtAwro0mhActFDcI
X7b8t6c0XzAcX1JDvYs0iXhCKzcha8DMU4qvkDISmAC8AuNyvGDSGEZZf2rJDYLHtOEGjYhsXUCj
L9wTnokCqGGjRmduj2BzjMPYgVU7YQxPK2oKmgxL25mwW2Y1sTTP+JRjNdaMW7RGZnSgSF5WsSec
RlRCs/1wExDbF/fjjylsWgHisTpmIF1pMyCGfiuBAqWBdd11cRJJz0j8/jam5GlQ6YpbXPcC206v
TlLblYDYkmnBdfr3P77AhZt8s8CR4B0tPM7/jq2f6/jxtiiKpq77EwU1zABuf1/7tozfY9Wqeu94
HuvhptluwEycRr0e7jOJfH80JMOArjmqaX+Ta/RSBR5o2Y1/0ThodSqOIAvP1c6XaGr/Yu037i1e
kqy2Ph7eWfF8qG8rsgXkXcpNJLPu3CRFme4aZPZq+W4Cf/Brtb4BpL6sbEx5zIm+OXVBaiDHHiFc
x15oPfVt6FtK1b8OWOZB8C5qS6IoF1sRiXZguJpmViTHH952A0+meV9To7FKzM59EKnVHgzX2uZo
S1sAK8vOMuBMtD2OfXuLpoKCXYO24QOPnQE6R+BtE6fLmUov5MwOFsomDBDhmQIP0lk5KDyGyd6X
w04TexOQ9ZBWP4oMCuURRlFi6cegeUwmvzg3fZd/euE9VhARqDnoNLKdesvHGD2cZMlZj9xMMZad
AerdXB3k0Ctwbvbb5FIdlVWLmKYihxAUSqSQb5oTBOF3MQWH0MJzwgMdLK5aSGe7Hy/D4fFCaSHP
iszgAZRj8cRxFsCp8Uth4W+3qxw8zLxm8JH7KOMq1VuN4c0wZLEDZ2kDqFL5qKitKdIJ5JEXgGP7
4hMbw7+fSU1iGA+GxYIpx6XB7+5MvBszZma8p6YwgAF1pZ/Lj/dgHzHa5PWGndL6Jb8rjfHXGVW2
Cytj8vXVI5sf27MQ9aQAiil+3/MiARlZC2F8Zpj7lgFPhzgpWIAtS3VpXwIHQ99uz9OfO6cTfz44
aKe91taTsP3C3B3sXLqEmjVmu8zh4z2LpEzevUrAxVzWye8uG20A+W9NIKirnpMiqx2eQgtLxy24
pZkSBD6ZB7vfuBGNmnXwuA3Zh4WNl4dYgCM/YsL7E7441Nosa1LP5OKlv9+PylIrEgoZfdr/XeOo
UBaRQgKKmPGsULZJ8nRa/yTGbPjcbLlKk+/LcuDLCJibgU5X5x7S3zKTTHFox5iHc5Y6ajkKtzzz
2kkxQIMqdtUwv4OerETade1r7GeeIO/EkcBfqaaL6Flm1pf5En2JuHmKOS/FqvjZm8jFEcTm7s1O
8+Krz9R8g9zLK1S1AvEoUBEOSCVDYhxzronkSRUzXNDSaKdf+DElMxKfLdrXoS1y0l+RRq6F2DQI
t+g1AcGy3XN9d2HNNTyOC6V05YkasZRaHMP+c3LI+qLvYdFfymzLeif8qu+BesWRYnywCAKUV3Tm
OayzexkEABa3GLWMJJ1zKpc/i4Z47O0/EF54APcp+JsyRYGGj+5206A82jbF5FuaGfRvNjDq02uC
n3V9J0M9ILlB88wFIYK71wI9FrXzO0tUMRVto82Rl7eXylRuuitwZlWVtucWPjcPyfuIFKbBYNyi
C4SL/tfrIe3mZp1KeOjfVowZk2NKXiSzi70WI+7V0YALdsf9BnX+tBaB61ajQ5QmeqjWT+y4DSj+
xaeEPZ4OR6LrqgeDzK39ZU2mNCjq+hMSUjZX3YG1VAU7M6KDjXVmwrwxfBm4bCFOAsA/ucNVmcOs
NCCrPt0U1eo7IqtoXnL7xu0baHXd2sfoa360DKnvFjvnWyFjT16AWgrhk2xd6AhSLmviyDubRmUA
ION7RhAeWxy4fuLAkWvR0oDMKxjA5er8hTc3rBI8QpPzLROgzsk8HkLgrdBtbdjcp8iTTJE/oKms
2EAy4ijZtX+xJloui028+9H2dEDr/evNqokcY5ptUQy8pCrnjZkXbXtuMwyn4FjJuB4BX3zt81Bh
UdsGw8FpjqRzBhHb43eIKjexp/x0voeLdEhkX8CgZw0ZSo68fXrTGfYNQJo0EcMJqXJbi3VrRmWw
n5z0iZN8siPcpZXgVqemiXCh1MNCUa+ONekIRpYsoVnfjjJfjTie/9FUDb/MO7UOZniBRzquEPjQ
zGVeEnnZ1Ob5hq8vbDVv3DqSFnZxNvQ02IYEnWB011kjV1vUQefLviqZ55pHjxdxEbnNb9eZi8nM
pFqXFvpQEGQM3yB8msdiS7U+1eMC1DZo5sFaLGPZy/w4mq1zN7aZO0ju0L9x3LCTvrKcKK/BfrAP
rzNrweHev0S9VoKCyYidboGwqcOCktluRCzj4f2x+tEpebBnhZZur96pC7JdVWa0/+SiwVl7wvAB
GeeDi9+e6L+BFimAFv6dGG8aFAu4sW/Z0TpJCgVh9BKwj0nrX8RzueEV4Ysf1GwduvtoPbOqLEeC
8bRao0beoj+8k529R8uXMmYctJ0dAa055bpWi3EItInIU7XGYL0SQK2g9OL9pd1+uZ2b3J4CR6DQ
/+UwALn72/d8Gk/kM0fOzpH9HntIOYco6e5qSCFDsBtUQaae+7rzLfm8ZcHxRpDq6J6HeeQiqMGH
N328h0HGDACYyA9LXintSzGCriFqIhnd3RMBQcuRWxYn/mf+YniJ4WUrxkEtPslJjKFX6GIQHbCy
sg4HSFweDyWZOPD3WkiadVDCBNfDiEBZTFGrNgqi314ayEcO0zPGK5TaTzkmL8yq0TAU5yeKnjFa
8tcYDs6+dBDM70UF9U/m9JKDlB7uLIt/H1FwnhxpGO+1Nbapzu37EPfLlxm4BerM0/HfSDKN5k9v
c2xRX46BhDDqEWdlZ2Npc1ceFzaSaG0F4zNlvYe6d6DB5k6WC27g4pLzH6t6zrBVGa0U/pfZi9WJ
SvzT8s5VOk5MX55cyJJMfiJxijCO21DkO5gs+UQEx2Qexbpt/OqG46XPD4wsleEQwtQ0KfkgfdOC
GAlrKmBcK4h2iOJaPdztftcyQ77Pm6UE8kCN2grO5g9RPV+1mxnBiF1NnU/ocYTJFPzsHB9E0rCI
85b+Lgvva3lPlav0G8+8C2tmJzPNt4nUKAZxU1BVYVUdB5mYlVS2yJ6ORYU6LjIYWgwqmf3ar6aY
VZZjWl95/CohML60yUICDfHDmjie5BNcFhe7qQ9IpwOHK22voJSOb+Xtj4N9HCwrJU0oTk/FXt3g
G4zWqb7crIy0kP1B8gPhP6Ct7A6MkBkfA+AGlc8Q1viCT+1smoqrMYYfaYiU4rS/RL9XRuwz7eo9
shdei0wvO84eXUDDD9j0p65hoN2YzJDR8KdXbXsVG76NH71S7LMDcfLpz10xzahveqZfhwgGL98A
JL3sFQDkhj8uInS0+zolBw5PDafCTnNS1OtAP9Ok1KYA4AFhBS2MBQ1l44Wp63WXHRt4z3bFg/bP
YlusczQQSQbmSRkRdcTFVOkxSYEpHVIjaaRf7DYGR4WRzUGe5mguJ0Bg9WDY3/z2DnifJMcxhx0v
5tntx5622yR+gvihiKGSyXk+MaAHsHbsYSZb0BXMmyJsHMguvadVAGpM//IhXDGr1c2HgLIN8xTj
1CJrrDQ4A7tuNYyL3iGCANNA0fnehpXP+24vG7rx7RaXsI2hm5wS0894bQTXQbfQOcAH14aLHN57
BoWNvuo6D4VGI14Cz+RNR59+IANkQYcqgkKsD+WZLx4PezYLcjk+td/Cb3qNgoBwWHqoGL31p/Nx
MI25islxJsD6mL8k+176zyQQbeGTh4QGBuVCTy05ZHaqhQrypsya2dtqKyfimuotpyldvsxu+6h5
SyujzytcPsL3Mfr1/H2+VUaTUo5M8WATMlIItRy97sSFrY9VNC8YVC0G5wHnxy+OzZqX0UxzVE0C
a2iTRZIj90jnde4CQGS0QKN+LnrnXXL/bjBC/TIJhABZIhymCdGY0t3ACVrPqlwznvDdmb1wdLHq
x9fRmY5br0kBrhdUBWGoc7x+7Jw8SWqYodXP5+0YnljbSOVnqpGVgJuM1FTWRRJL1ImRiQidSLUG
eNO6bWRjcsbgv3g7ha5pvujGpNxQTf6qUFj6+Tf4S4FOegjU2dM/9tRQib4jJx2JRO/iVnBtac+l
ppo1v+Py022D2/pP8mBb9TG/E3Q34dOKnLv1K4P0oVNC15/v/d8AVwpASi15u46ZzkWm58LaVGq3
P8LiWMx9esPR+iRO8jsnN81YbN/dwuzydFvto9JD+Vf0S7rk2fwETF1b7lBBUxpEInMAbgviKn4r
DCc56zRzsffNit5jEcwvHw5fb9zbjYioHdSfPD/tk16L47NSETzK6enXqvnPZR9T2QXnsEQ6+fL/
fKYSWgbyxkuWGqxWEAcqWlMNlzzVcYkQCrZRz0BnnKs4PVsiWqRYe/xjkq6p88XQno/2QUHXKwah
t5SwS4bfctR/yAj8BT7b6bbFExfcRdAEt/LUiLe0Spxtr7yqaLPsXf6W7dZ4llJcFtWgZurReZfG
btDWYgiwOpfbkTNyYvviYrjSdZ+/zqhhKmLOXr1X8HnQ8XL0plX12KQL8iAdzkcggrgVwpiFeaLH
KaeGOBL4XmMoYXNEk+y26hWlnuV8dl8A7K+Z3NNCD82IKpJWtEVYN3TEa7d6qoxBH0bn+rWb031G
kyYaGJgsAAq45BER8mhEln5rW70lUSNhwn4RS2r2kqhTByFYNS5NM51CtBCZwcVWHD6ukCYhZ3xy
fRXwGXFxglJb2HW8lLYefaj/fkgx5rZ1hd1/Zow8yzqW/Fzg8GlpUgLNsC6bC29Jz/Zofsxu8UAa
Fs3UQ3EjorlV9w45L84CIJiJX+Qhf4R1oY3ZEcbIUAWis0RFVP3Ryd9IbSz8Q8SWkLCCL47moHeK
tcNIKoPGKvI/b3o2Dj9WQbYsMXHX1qUtXJ0iBS7+ic2Llk8WdZR2/ngED69DPxbZvs9NR/X8sIXs
qHkzxv1Zfg3Qn59LUTO5t06UOuTy88jaozTihkmcs3U5o/w2PKHtMd5FdckKBZyHvrYl7eJL2icu
510EMdkOK5Vgj/hJer9AX0sdvUchoPZjKyAgZLGGDyrrhUPje4c3hWfUHevqKxb7LwaOaYeH7RP0
8aVZQX8eO74+pbaIdicsOu412OZOvR/d5cCItFPlWG76nmefesUjhtGAfRCYDX8e5cRTUVvh19vf
VvA2U1cRPDUYscGGgXAlbPmPyBIUcjNdBfu+QCBelbLRljdhlZxP9MeTBxFkn1Pr1+nN7M/5/UNb
yPWkqlbEyNApMWW+zfv3PA1tXV5mkpNGA8oGRBH6qmUZ8RmVN8b+BeFpeez85/ICO/LcgOm+Ihfg
SA1c+CVzS/a1CprvuPkA4JMjsaaxDEMgYbJm1EOVlL3vqP1UAhQdY1TLxHlZYPIrU0DWWoYGMmOr
uQv7kHw5UqHhxIACL85Kozv4Qkqon56QvrERE2GaFGo3H/ch7Kck/XMzs417GRDgADTq7j94ELEj
FCPyXN42Tc1slnEGIo1M8bgu54SzkBoG10jkcJtQM8wRK/4gdMTjhIXEsc6gAy8JN91PZKlkE0Pr
7CbpvpQMMazTI9gX7HX6eyptljsHG8xeiaoH7SeaRV3zpgokHHgasYjFfMjNn+bmG1aVvICLuBPg
cPw4U4Q3XvKKZKTWYeOrPvdZDV31vYelAY/lUjSK3lUgnBAnUhcIrozAdS+10sPlmIUcUuiF3SJZ
KfChw+zD3IWMszMYhZxNKJZEwEbdT3c9eDrQBDSJOvKr/IAO+WKgzde2UYXQ9DZB23Ux3p8oOFhC
UbYBSkPDK55hgz5Q43GR+rE39JtrOVFbnaUQ/ja7tcn0nxMSfdLWAMN/f5MJuo8jaNXkv9TPZotk
xLtsz3KAnWdN2jeszNB2Vhj7M992LaRT73g76CV6uQZF8oFQBjsJ8AUAJJJlxqiVIUu65aUmapim
uSU7019IX0F2SAkqGaPernfLSN4Pf6vhQFHtidvv2adALKEY1HQazA456NQKtokZ4uBKvsrr6e7V
xXmtcAQuNM7/T9iUgGuZeMzLeH6ubOAYY9ifjwzBfgVa3azzADUhQhs0IVPoG2+83Kl+IunqiQPo
huWqmaUFfq2Ktgwip+xzYbc8d5H0qhVN7mCvTu4bvs5/DXTKpCXRG+svcTPCY+rNzV1q6j9KStOk
INaCqpHc1tASq4cFCmHxBWV82QOtceHi+TnAXUVzPVEdyON0hMTAx+5dp3a9BHlYHVRb/izID+7a
9r1UMB0u3PP1wRGde3QHIesVul9kYLKpmFCRmIsmt+laQdeMzWGGrgqtH05JQOBT8Lu99OPjWq32
fidfn2/2+TPOpHUX+3aWMDpY+iIq3mAZZHKTfdTIc4o+MVHg5gENGo5yqH/QGmfLywCMNHcW3yZc
AAX/1JpAYorHV06TM64LASs3yCIbxPfDzk9aRdymjRoAaqbGWfJhQmzsrxA9nFk5Y3xj91ycsINl
NGbgiUyGKfjuOF7LT22LqC36RIZWOYViHsEV1bzMmKKiqNVz2DkaadvVmZIl8ZShUwhy/G6MApr2
B5nnqgmCQU8Q60KvSyBayrcca5aFh6q9JvxO9iYj8ae+yzD2n/fTEJU9xJLWrh+YtdqE279LLlZt
d7Wbxf70UzYIEfFZ+6mm2I15Zx5dCGEMjWb/IfVz+EGNiyezlEvRjnnRYU/TQZO5bjwU9KRQYwXU
oBPyxJH/LnEsMcLkQzM4NeIt058dHnKiFj+P9uSgV172vKkKDKqeY4u8QCsylNDJJnjs/oXNTqI8
W57Hw9vKW8M2oGHBRbWkeV+qgxos0AaGIYSX/UmTDhbvxUeL4eGBy+Pz/HDCqE2m9D3RruP78SUh
PhLGS26XghdiwM6AAiBQgDfYkDXZypVFHas5f36a3LHmq96d52TNhYCg1sG8Hu/tJ0cGRBgmdB4M
PvrxuqOfj3yalj7atltGNwV8E8iPCm9JYINNHQON6vVZFNWXHouyX5qMvfw0xMJ3gkxRcQgZwLh4
ZDBbEPfoS4b81ZbUufJWiPPLzrjgH0RiKvzNL8MmWehKwllqUf4n7MLr38xMQXRG6HtIVABVUwrs
hSnWHZoI/D2TWWBIhDG1lpBss/1U0WgzgI0aStXeIXL50UzcKVHNI26dpr0wjCPpuv55Edi73akj
ypjYJrvykV9dzskd3e0BD/BHp1X/lrJ27B9+QG4Z9CzJhAqhe6njt8n+HHiO88mYqm6Xjmrkph2o
O2B2eCBZ5WnVSwluktMpSyzh1CnLGebYswEcJRE5zzNH4laotE0js2maYzvAe5Y2RYf+cOpsWIxJ
dU0Gp8/Y1Lbdi0niKK3Objp0hhq+ErfcK6aTQ9QJZsqYxMW9qZ4GEMxRp9s7dzxvFc9Sr4zyeAHO
dlh44sMvg2ZbJTTcWYDEeMVx2FFxbwq4esX3b6cOshk3NBnWtquKP3EbuFqE4IQrFPzvOsL57jvf
4UIrzWHYVB7ou06BKok99Yzcka0sNRlL7Pp+ZnKcJcR+8Ho9J5Cw+zEncrsCOEeFVB+YuPN6diHf
2n9gQtAl22bl7xx0H+sbbQOFgC/9Dwpy8JqjIQdN15KeBj4EBioyBjrEn0C0U5iBtkID9Pix+7gt
IrG0tU6UDnQdFNTZf9iikErNKmgBev2vop8+YfE+JOLljzJhQMnz6SDuO79GMX3xgJkferO3jgZj
DG4KpgM6MU7d07O4mU9YaB1kzRfH/XHS/4PUv5uLp9R/IZ4Ajx0WqiOHz/kFoNUv1qp8Pwid93BN
4YBitVB3BmSpBRNieGKtbFgnmvtEdyCWX0eDCjvdK4PYh/SRM+jfBWcbF9gM92epfLzWn7oZ0pne
CnTHU32A64PVYcJzaLplGVmN/hwWWAAuJ4P2HWMnc4N4bdBxh1c5/HHjEbkfdL+JI6L4hQkM2xdZ
7FUT7+/iqdrcfa777yPpHp3cK9e/rLZkfdxR+u7hYajwv6+M5TAtOAK3OrXqsN5DwxqcqvRwejmy
xW6mb51sW8sdJWtzAi4jeKCz1laimRtF3jl+63IJnbb0dShStNsAQN09O23ZNMNpngPotww6btMZ
hab9fISjkHhsq2kM0TrpYlweLLHPD55LwqedfDuvL3htK1liXJjdvlVudb4Hn4FghjbsM0FtQPe0
WK6FjCJxnQHmXsGn6tRQKAu04jd7pI9aIGOQ9IfF0LuuQYy3544ONIREg+J6AENJoH197XQXExe8
P2E9DkivbPqjRNbDNvTnrhmVf8NEhRyjGOIlWKqqj9Sak/TPsSJMX5vDNskebD0sVcAIpNmM6d2Y
aHKQ7dlVvcPM8wPlvn1AkxDO4hN4cy4vaF7gK7Z9T4DcjIiNDeTEBrURifETwkJ9cu/x807AG9o/
tDPFv8U20Bs0p8WzRkvqd/MWNZR25BF19lJkiKcngCequ7brTFU7W2N883wm+ofC9lGGWXejDg2X
T2j3t2E16H7cx97EKPkchrIwCGg9kkalpmP+ofY3ru/kudzxocBe05tsto3RYjt8dSst5Fj4BC75
GqQjgAiFAKPAopvrqkYAwyMFGZhB4dIpta3wOdGRx7K06KS1T0hjym55MdPr4jH/KxpXMa6WrLHg
NSv9fE7jn9yZtCq1xUC1lkle1kID+Om6QwN2Qn0fnsA3lFGGRR6PNYX8ZNFtrLDY8SGbH8k9mw0U
eGpU8VO/NJFHPi5KYJAbiaELVRsk+2ZuAEBC6FpskP5Mng7jxAuS1RpL6Ze+WRyH/QskWyhDADTM
NnS3T88RlatJZ5y5J4YFGyA9VxhdQbQEUdfh20ohbjC2yQTDeM1Gvc8zlq01yKPq1M2Fh7CJxNgU
EEtClDthdsXuov0AYDSgQHPQHaknHtRE+/QCiH053JKwOpF4/3DAUcmyVBXoUngQ3LpnN4273c2K
kUdcBUQOR5AuTWa/WFn0yshyNnM0sos6G6WuWLbzHDMhqetPMyxu1t/jldwjm/HKug7b7qXdh+Bt
zttl616MVLm8ByKYohDcHIFvW/wU6O7Z5KNx+jWaCeMzUmOFfUD+JzKMiIJSU4Z/lSA7sKQK2w3C
DSw2+2ApNdTHX5AbXm5IvivuDEM1UYuJFpPtcPJ5QsAazPEMp5jM3FHbsXNGz4W2LjM1oGU3j4q+
LJz1UBhGkYRJ7uascWjc3t7iP1Smub0i1Naz1DP0mZkkpFd6hLK5SmmdXnzaGRyRqvuGvMkmqWdt
sM+QFJ1i6SX9v53YhOWT2kIvFfhN/g58qjL1lLIYZdYkqCwEthXxBTlHXCpa5Y2qnhvwfZNADxbh
mh4N1PHQjzlQXN2/xPHpLQR3gLSpCVJS6kUVaeXho73FTxtDcDKVuGZ6vL5vSXarMUcDd+0lsHps
NpzpG+1CfCkJYTUgRglMM+OEMAtpVEUrv2IchLO9fHhcmo5qALj85o53ndryiOS4c+QMsGW7vXOQ
rteFeREwevICX6pAL3G+mPIhn8otLZeobHFtCE6O/CV+rTVN0fSR9/n64Thu62yCRD2W7PxSXvKe
gl9rYTHLXOWhlGcsNvY0vCSHHvvf1WxfZFPaaM+IwalpnJCG0D8djh6g41QWxW+nS+8/jBxSiSqR
s1ayqohV5ZeXJCS0xpx29W79lgcmFTUEzHyV3/cCest8vEw+GnDF9irkw35B2EfN2/l/VGbs2MnA
14Cb2TqtwwNZIsC0Xxy3vmMXiLnyZmO7XtW9X/oRa6dCo+ouNDxG5YB4sfgc1zi3XftofAPj7mqJ
+AHaX0Le2TAzLsUrZOeWkdl66xfMhsRFTIkBwyxfIkgh+2kkGLUoiyxo7Qo39iyP931v3cjrjHCk
qB2tYL2i+1/ynsBb89Mdo3sgt9dm+f9EKXWf+47URf+YuRSev+rtt3EGSMDMON3er/1vX7fO0J7u
6YR+zR6/xOeTUZC0f5gILLkmOyWEf87wVPNFgbm8gwCi2/P+FNVMF0qe7NqCYNkBZBCag0YiE/5+
0cI9B+svWIfkuO8wS1X+Vode/ex3bo/Sf177gIb+8AJFkrtPQaKb/IKM7KH7qHkThSQgfmAGz7k0
+yumAcf/uNzkzkTBJf05M2PmQqsZ0Eoj7RCWnE4Mr7qXWKbb2xOQEiuWStdJJLDUmNEsfkxpZOoG
HUOeUkSUeQJkFrd1M42Gz+jr0HydgDSAktQ+Y7fSkTE8MpAFtVGr2XbVEVe20PVEEezejqV74zoD
6PbaarIMioZ+ntQI7heCGKPvM8TRfz4wDPrVY3ZiGdJA/Slp9B549xCRklxWJoIgTd7/Lu1DrLa7
skz46KStgzG059TaTM86oXQ3jhwraLzHbrBPa8GFvIeA2d965Pflw7YG3LWroW9AgtfblFWbeSNQ
sv7uwn4aL/wZ8Po83s4VSOZud+BdtkxzymIyec1u2p3KpNugMJ89M/aH2L0E4+l3M5LDotJc7reI
VBitqbYXurTyS3aGKvMtb50vmuCfWlxbqOJDRJvwSUXvTt9dvIK42Wf2ARRwBdY5NxmyKKXZTCnx
oDMH2tCIrQp+sF7z8ZNTCpXcZZaZLs0/IR05KLyvG4dfhCzTwH9xv+p2/V9zXxfR5ZDCjkNZ7OvZ
Tl0CVGR7oMelgeBXSKR4rEBFxtRn6rUwFTubfzq5oPeSiWfQFaxuHEf+O+y+/F+V8wkUe0sgVpIr
HjfmpE+BQ1YZBG8Mg09hyILiZzZL2bC07jvneSTjwXVK9gr2U80BtXzFQKJgFU7hn2hjH8pKGkeD
CUMZgDZi7iUGj6R7Ig11wXW2bt53QSSXp+H0dCnNM7lMi9fx4quhCFWB797SthPouQ7+rC6sObxg
811n++190n1kv7dV5SujyiBixNmvzIdhwOKTZ2xPTvgEhG4xOuBtdAXlaVFVgzT2O0S3Jja9IYsO
n20yIMUtF8mZlbrYgW30TCvskgKr3+VCjBKhp3vO9Wl9cF1U38ORvOwxFJIWc1dL1JRpaUPwqsDf
AYVSh6yqRXh6ifmUx4Baeuu2JWLlqZRBb1ptzbTvVFwPZwdHQTk4nO+PuJW0Yjy1c1Ikj1aNYxtA
Q9jyXWVu1+jorTVreCCOcjCs9zTkI0KHiRqjz+FDpuQnU/65S5pRxkXZHUYkbZ1uQREJtgSeRrdh
VCFlj+CkKlu0xSwMFH8k+8EI3JRZISlhFTKvzi8DD8xEjRljLiRQrDVcIwodUZNXOzDrwQCkykMv
pl14OyHDN+gzAyJAktC+lBTs+Vie3ipSTYBjVJhps10aUNPW4PoCY1C1e5044s6Dtg6oa9rcr/MW
3sOxF3qdjQQ5vGseddglxgopiOi7bLMJ2yUS7gh/o+7xL4L+LIAd6eI+wMG5IvZ237vo2zRycTzN
mbP4003n3U6CYC32a07QI55zjV1THu/yNdlSXMIkSfP4Xd4eHw7Aw9umXC5UPM88yn8K89KUFPS0
HuLW9PCHEI2BHEZ4n9KhG8zjivotAc8xnJRaSi2lg2KcNNTHOQ6K9xcVLS1MoHFhTl53s8QME/eh
ysK6fGDufymviJksDddk/IVI6JZxCTGNACryZ9e3PYa064yNuPisjr5oSiVBCCH02EEUcK9aMgEG
iAcMy/OqgpZfEiaoOVDgi6BBgaX2ywVEBS9FrS6/fRYpl3Li+DvCAAdXYdoXb80+eRiY0FiqTXIk
u3qApIl3SoBVaB6eJkniwKOzEjS0KzRKMXudgipHK43gNGucEFYjdxt400MMfVGMyhN6m+Qo5+XW
QsC9pA4HYP+gL6xymbKGe/cHQ1sos+FPtFBw/sICypkVqxSlvjA+qJsAyDm5+++EtYPZ68m+PVZD
KBx/T6+UQnX07NeU973VLPbYdTOzaxpV43+YG/P4gxC22p5xYAyqUa38nQbtvPgKI4kaQUd7n8qQ
xraEk8RIzyRUu7lrNuqwRdunkLdp4qEgxNXkeF0UyqZK8a4KQbG/Xwv3wXnE8Y9KDAZeiTcRBGm1
odomK+UqcmMmqW5i3FkiFpK9Eh5lpmfnVMiRTKtW7PooBTqujx7D6xWSuIlFZABjlEvu9ZKfBvWU
bIpq8RNy2nHjHcv3hrfwzfgRcp0F667TKnph7b7/j0+YIxcxSqh40axyah6eMPUFFwEBHL3V6fuV
zbQUnc6hNogexuqnjHv0dFYDCqr/1tzGxgO/ifB8silS9TfIy5CkJIseDV8SU5jgSMyZ1HsjhDdx
XrMzcYE6/viS/14RHx93f0r8pIIcE223SvpPg4TwE66TV0NZ9cMs/2JCZWZa439njoEZFcRLZ/yQ
AzgVAp0MD+euiXY3Jq9yc4QRiUAUl6gOzNEiapS8W3v3lUEbIKgGVmXqMVqcbI2W07r4QoOkLud+
hHBnPZA+9GfGHx4p7ViSdpXDd5fZN7l3YbxeaS+BN3dk0MuGfmfkptp/b8qcjMz7uJZ1sIY4M4dv
1ZVrDoLBd8ITMBtHqAs5OpgGz0HyuoVJcGJVywCm8/fsVDN8NWDZId1vnzr6YJ7KeaqIOqiFQPgH
Z2aBs+YJFGuUvhGytcO5WpJU5kSs+gOmFYKjZJ3IC80PBUxoAGLoN8xZ5+vEMmOCcjP3iMktpf4/
8uDJN3JC3aomT/JfnmYgzX2eAHiwgZ31COQTupJtLoY7z3NZVntDj0p6fyv1mlvSE430zNKZaPCw
3cqDwoOTGvstipBmP3nu24+qy/aujatM2tDt2VH1TFqqGlhGfIKLYYyfJ1+Ydi9UA4+TNDTubxmS
dKc6Srurs2NYZhOYkSDu9aErgT0C6P6nfc8Io8cDLKceCWO+MiNCwmN0DG5cqiLVAmnAS4x0eHgG
ZDFZPLnipOf8a7xhOp5UrkMmAmHOz9DyP+KsAhcHQ2l/epNn2qYo8husYDSbcPtTeXsk12/4+Mz8
Xk8F/NkuynLQ2XbbjwznG2Ud97eQSIlseKE6MBZMmDZn8hX5YeNexQcwCbbzKK2kP2xm3ygZ3lFW
myYAk96xlwT3oG/tNwX/T8lBeI5yQSZlV0b/rPGo1rDy5OW6BMysRL8QJXRX5VOme9QNRy6SO1C0
ikZkPnm6nr6Dg/mgc84tQ5uFlPlHmV/z3Ju8tnWdth7xOC43tFyJvp2+UEsKFNNDLf4N6OcNSQDs
2kvIkwCuJ9GH0uHOOlfiVuQqfCbB4YdlmJZO3Eql6TEatlIb9slXc6W2+6yxX2OrHsQ/rDSedA3o
mrcwW0EjlyYYx6wuRbsaBt3bl+9IWVncrEPVtGUYPrD5CaBUOxWdVf9q4d1Z8BiOuS3WIMWW2WsG
mon12mwB4znV8jeUHz33FWAS54uN+zTN+H+YMOxgZr1X5w1Ni7JZ5M2ofFOjJC0yjhWR2rhsyVwb
1kf3yhzNRpWE+5kRp9W8GB5JM+TgeNae8EvJ4g+AYluHQgZJnyNHikhcOc8uQr52lWJ4cWUH64FU
JWbUta+G0dAP7OwnM3/tY8zgiox1r+0uMgEWFv8gLjD3JQznc9J9JWKwmX8DehfITFBERxnv4Nuq
XT64FyGR3W2VinX85RpUlCaeoFrTv/BVjOYe2gMjBM66Kaw4hLA+q8CSa+w9Hh6LBa6gH606c4XE
wIRukYh5O2Pc5B0Ob/nds5cYsX9+8GvMtessTo1DZajbRrhzZCd+AxxzDvNg60arCGnvXjFhvu6X
Cejvroc+tB1Wc0wXiq05eBbg1FW8YYT2UqsQGr+vnV3fqvgWHeO3cyF1KgI2PZ2vRzD8D1KsMJnI
H5Ns7HoNyZjsFId76IrMlfhyAaHNqBoyi9zMLVu9Rpq7OVPCObdZlow2b2xl1R+vmJA1Ek/H1SCY
4X3VqEZPJkIOgu3OFKQteGWDckqcMMdbo/DfVJVhlOq3RqIgadPtbjURip4LYxYVQbw7R6RBsqKM
U+DG1NG5l7q/SXMNtDJqs2U8MCgdbenrWGazQtpfhWQrdrNvETxPw/TotXtkTrtycf1LmgNcAx6g
MZQCnIwR3wQyExmoFUytYazXX3SQ6LIN0AOIBeGQcQOAHFCioWqfQzO0ZFY6gPDlVB8LXlt3XWKE
8SUUN09MACwxQFLkzE+iNTi9Q0KCq0OSRjg/5bg4KkJdUqLU4HCByM9djGpIWowcS3EkcnK965Rq
kOxDY2KWy/RuLcZHGHomD2wkAHgC5KMMJr2FYpDH45Nix3TL50LCaCap5Kg+TQFILCJyMzshFfou
dcGIsO0QyUCcVsd5WFbsdwgO5KCjE+IORcMzDi3thsbSLO6Vi2TAcNgFtZ4CnstOHln1mWLJ5tkc
7vLvwW7CmM31ShYohAtkF7QwL3brD48Z83VpUaLzvoDN3HadzyrHudXdATas8ktFEtz64AwjKXGs
JMRK3fCWEwEWGvDc+HgnFKErON65NU6MDhSAtR1Sv6aGP+SRsJ8HwoUIHDYG24pLaLce/YlqiBWv
5xVJ4Nir6mfRz3kWaJ5TFNkyMGQdJ9zAu/bhW/NJtU0KAQaHahAAvOpkeTYCbg0Cc16+jaLeW9i0
gTty5sjvUxuGpXxUqr0fvbCN3JwDE5ZxLjywv0mu76HtZmUeW0FLaQMTGn5pmCP9dsW9oCpVj2f+
8sUdeZsxxJyjgkujjvfPygXYkEOqceNKTEBtM3MEa2oX/T0ynkdxsiU3YeDt16uSWLvzf1xd6yuZ
KbI9CGsOHM5UnPgE3zcDZ6Fk3xkeawgjPnZbvlzz6zNPziVb3KmM1jNoWP8H3JkULBTHv/vxOwId
wZK5SUh1ABifE4tOUXcpVZuVl2AYPsC5SkjRPxcjmBSUxnQ9aocdUQEqdwaYjmPQnn8G9wju4HQZ
7rG7myBdlbsttOkfP8qJGlNkLarH/DX6UPuKMOXUXS0RbR2RlvpaEAF0g2rCZkyoxQTA0lw9T3l6
UWJEBHtilVsGI4uacESNehfG0W959+UzhtEXL0ZEoXZAVWvtQousXGrC1+SWLIw//fb9Pv+7lCup
QJKqtgpI1x3eGzRKlr3/bZop5y4KKvPsV+mGTixMlnf6excv8k2Etrxpz+MJ4QREzYawWvY28E2j
sjNuMQncOSMIfN4QDPmwGc91J4R5lq2EbBVmBbQBmGvBj/KrUBC1MhUqQOUpTDIm5CwQeTCW7s5S
aS/6brukTS9wJhVR1JjNYB6AWYVYvxYpj+1olNumrTRtx9xSniMdTT3U3OlxTJZAEfRCxQ1stjF3
CqK/75dsFHbOQnxzNRBOdFxGZLyX9K0plse3QEhgVhCpXxIvalepSYajhkaLlKp08Kxnro7V+erc
/zTmakkO/LEK4HrKd/vObpYWSRfnRwobhhJfpbK2wJ8DdIIJ7k/3zF/pDiw3gB/RnWf86+n8GnyV
FIxdKMYrVBYVIHkwWrk4dsgCuffcBmSzbCnuyIGkJ+3v7yxocKARrRyTUEHmiRdqe/M0Q+WKHi7Y
eTEFf3UN8tNPBGW80iY1CY/kZKk/QplfMVhaeDQFkFac08UEQFJoQpPSVNVXUtG9GURRvldyYGhq
5pacs4B0KZlO5ItaFacWY9e2NVcghMsJ9Ja7WNJNg8mqeJXk49dR7/JdR72Oygrar+hw4oIPRtoR
iEVbT/Zwh6WO5mXyQZpDUmtEdzZJ9c21GJH+68QlQlYHzAPvCVz+2m0kV+Qh2ZJuJdtvfYMjUH86
TxZ3xxf5oRagDZvlYVMBnp4Zq7bimKM7SZ5Kn4NyHaNkM1/6LMjjNBO7INNPpoaE4BaiRklYu09g
+cftXSPksZ6XvoQC4pXeP97TmIVKWQlVjTFBp8S0rynGy8OOB0OVL9bglYecZn/WF2PTof8IQLVl
0Cj3+Xm/NNt8oWfAVeSMfgLV8HvPYO6/LQbHaX4Fs9pOzVgwXPXrRLXsMLOrJlrXE5peNLYkBD2c
lzkUY9o3BcEZnT/WUPfWqMiqT2cFhuciFD5K21FBstTk0lXsFiLTUqsNIPNpc6sfNlvE1p3PAROu
3jWgD3oRycoeg9/b3gWTaaIeO20VLJ/1JLf1RRgPxs36FLwtdIeMlNDVMqMsJ4c2KSljwGZYClIa
RtSrp2e0Fyc7whxpEojoTJrO9CkdBXXDq34CwVbc/tpYKYXNakaR+c0R1d/FAnWTObgBSkARGtEK
DEedvvEoENWEewUeTHh79bF+qawqbZOY1zJe4aOcwoYiBvKkW+UipbK6UJ1vQ8hpO9eJ06FoA3LF
wm0tV7r6k/pJ9cv1awKE+YKIMZuRmbGNEonHIJPxkrOnyXaXBclnMwrgIfYw+pb4KwgVpjjK11Zs
Ut4iRVrTk67WPJ5ESoZ8/cgmPzW/54FU2bLvCfJv/P9oB6LgE5Nb88eVxreH6EKz/nciypMUpo8N
qvIlI/J/Yx0Xjn7nNA3NTb2PN6HymkUOBmqFaUciS6iyxhq32L3/QtiJA3c/A8pimh9sNFjIHzM6
s0K/he3v48rdSoFVDcygkEAi2sohtPD47Qu8UXvnCoWNvingpNRk5Z+PvLiOZZ4m80RIlGYjS1Jp
AVctNmhaJLU0fAmZH/p5mLyGts80fU+MQiQNaY99+ywPw3VVCJ5esIOTzOOfmWOc346+aNvnCfkv
lqMKbFFFNOf+j9UW1aI9Jo6Oey+/FSaiHSipEv/OMeQvcLtQEIIy5DZtSjh3c4x/25BKNddWbTPp
T9gjlA8FJaggwTsEDh4i0u6Qliu+FPS8WT6MYv8lHKU3muPPqr2A3wPGMFBTPscRuRbjaJj+yKiA
1crHZfBJH+sIPNYjXr2bjm9Rhq7MYGnLW3haaZy0di6COICZdmQTShipoCTwTzWDf1hL9ERN0zy/
VGR+WKGxMR7QSviEJtLVLjRGqxYROW20kPrXtdwDx7EQ/Sz1MB57WjqVn+KbOmStk7E/BejcYy4x
ytxHaRu8oTVa2wiSYZ8KVrV4VLxebuIraNo36RqEmUxEwMa95044zQj8cCoLCh4FeK26PxBq1KHQ
oxShZt23Mla1VUyPa69yxjC7wpDjIa/Bcw+X29J6129VQxtIaUeLX2sAWKO0khDilkfJPsM/rB8a
kLtY88P61supdLWE78eL6P5v0O3tpqv/GjBaeOGB+A6LSDIA+nSzqcIl0Dyww6T0xptazZMCTQBu
qs5ZhvDdVv5c1yaAc20fAv+RhEuxsQgimzDQOS/s879uzqcbz3oG+k27byIxr7n7m13LgP7f0YPs
1GYkkJwwoV/nuQqU/5omxIn8pw2eKSBV/iZNf7hoQz+M8EGfiF5nOxH+32HuTwvfprkXtmOmCk/1
v33GCZXvhqxC9W5908rPb+j6BCgI+faG9ChPivo0y5nxOHPn61KNgwAla65Uww8rL+uRI5hixg2D
lf5ekIPHYlmZAjGfwFA2RrC3c5Xp9MvwiaQ7oq0RGWqlU6CZy6V9LcA5biQys5ADAPe5iLP4bV7l
Er0I0qknBEEiGm8j5e0mSfJwAsKJvCoOFeFNsL35w5ZlzN46bLfCZTJSsppN9jTcKvWE4UoTHCMB
TRRSiVYhai7HZw6urk/xoBLDFEkeVA3A5R7bg4wkF/IFfiLqlgF8wp/CJGg0KjJvBrx0wjHPJojx
t6cjAo3vgZXdriB2wD6zBSExQxhTFrN2sTvAcfB+hqKJ3iX5C5ieY35xni+BNtBCGsUpRwfI4sbi
vbEi31IayIh/3oALduVNZLPrsULTD1hHcoFJCW9L8UupeYoljopioD8kg5HGLflCq/FYtdvP22g7
PpMX6M9zuUBkDMIKEdiMDvL/NFE8JYT9vcC7025APo5JV3bWYxUF0JUBNWfVAJYNHeP7RYxdL2eu
HjO7dO1OoI2+EdKx9QULLiRwIEx26B6gwsCtSzvj47EaqIxhMAJ0uNmi4AMoX973RAwcZbjEAD3I
j+3uwhavwNCeO2/hoz2Z01X7mf/nq2HZnK4khIfY51UC91yrTP0fw9TXKkOAL+Nj8VHWvUh8eWcQ
9pAL+jBYb8+OB5+r1Z8egOyKcWc3j9s4urqbd+ngR4wOAtYTrdGCk+SMypt3+gPVJ6Z7KOAApGrL
XH6SQAtsOeJn65iCne1WvFb7Ey1UM5B7YuZEKy38Nh7JDen6aAweH1/kb4mX9IFMpRlmN+5oviOn
XUlv3FqGM15LamIQYIoW67r0clRHrareb52ggIBHtEkDp9JbP8BLs0Kp4wio4n0qSDH9/FGloAYO
X0GnD4uBjm6nKY1URmdUXlygX1RmeVHiEmwneF89H1Ia3QKK8vo3+L9VLmit668eJH6gzRaA44MK
ccqcH/8seN9s/xiVFthJrZTxOTUbRj6f4UO8OHhTEhvWApBay/d2pofw2mX1Wvu94sA7ztbSnAp0
zlXygyEIFz7PpOqUF/zuzxuAJgr1Q9KZo0ZPKjSgEhT6Hl8vTHkXBTEpi2cU/0eps5TDl3B5/of8
0CCOMb1OumPMEJtXnpP/ZjQf5I5WrKSSqdPEf3HIkfWGS1Uhy0gKphlW9Bs/C9oaO7ODQPebECsQ
2ckgQpmy/vvzun/DY3yhSxU8xeglZdgcNxqaVLJWY2c44pCfezX/YG6/xBpf4JWmxYGuhOjsKpFF
A6bieOs9NW0l65CBfPByvcr9QWb7fsFjeAKMlNyV77zHy2MN4LS6hXi815+VMJj8AFsglTF/9P4I
cUtWaMCDSKXgF632xitB/srmLVVE1ayNN0ACY4ajaTUNC1L51PtcgLxzbE6f3EKj5HASMAQ5hCNr
y5ENqIkfLGxyy4r4naOHwzaTGL3E+g9uMVITlrrOgVRyYYUVy/5vnCykqnKGLwusb+6d8dNeKmXl
/Sot3Y5woqDsyCq4lahDccA+69ghtlYCdkm21aRca1kg+AtO/G7j7ThXXbBNbH/EfzuInMOAM7JO
h6rp3nr+EHSRjdVc0jfLzm/7UbEvPPML86i5uaywWqz/TmQEIdTdCeUcTB+P2zaGdkIUzSNC+HO7
NCz/z2OUwIstHEUTtGOYaDAh8DPadYYWVRst/+nahJsOOy445OMIV6dd7+TTBjOtRbvQtVssEOoF
gO2QEgRuOKgT5s6Zp9WGegE4Q+fjXAZ0T+USEoHptQaort8ObsyANbKIoCFIwn/esBsZaORTHa+L
kkUB/EgFs5wTmbdrsoXgIwjYdrALQHU8t5KjkdvGNNnghSaCq7LbkmL8ishIsN+fNvUp/UTZAS78
qhH9cPbgvAV02wPEC4neLyHANEW8WzEZFmfhyvYGoXk31WIOjq5vR7z+7Qyjr8r7GtUnEp9b7YDf
/nsWwdzSuZbH3xy3J5t3cOydboF32qxfavdCab2Joktj3EF3uezAZHaFDx1QCp+ieq/OmeFvA5Mi
PbmsTKRRSVUnPUXHlrVgn9y0pnyq89Ax7xYl7Mc3I/PZn8exVcjQKlYxpUpcE5264W3sqjCpDMzc
GigG7nc9xXvyLJ0gvIdmSR9qGip/X2oxXsOr9YgUkCEnjjket/jj+OX43W6HH1PpO8GqzsKqwk5T
gigm3DEWcdb3yxAq+HZ0XJrITDmGcKxH5uCMb+HmMhWa0EjZIheAlEKKgtnocXyjqOxdUkiJ9Lxr
GCEGlAnkCEhuGdKwPs9Kj3+uxfqamWfixLV815fXZMgtkCRkyIo6QU8+PND0CPB1JLTGV2c1vgRY
5vUoYWOBw8dRXTkZ6jPysiR1gSrp1nInG1ZnP7z9YtYC7GRRlgpkq5gRP0BvTu60chfbLVr2IYPD
AuImk9ZTZQBY/HiQwx5OuB+JrBELxCDwr1dZq666q7s1u/Sw0eVn8kHUPvQbruUHv8/nsxXWalNJ
JS6gETvyZsZDk/mc3wtSxBJ2h52Now26XsImXlq0+9Wr57ylypddCUsSh/uXQMHdCCXm04k7cDVH
dZnywxnbnaIcPJRs5sEr9ytNjgSvmfnX4+94SKvaq4yESgKMg3bSL9I6flL/M+Mj2TStx/4lHGE3
u6MhdHdplcBse/RxxO62bz+rzQV14+C2cJ7CpSG1EXLvU1NT4nQybBda2+8nfmJX9xx06uEGCsIZ
4CZ4Ekc0WZYFMFk8baX0oYVnW9lj0Ttg6hxkh/oWjtS4+UkArTorlrkRDnjp7PPetwSQZHm+PzPw
R/pQ/zMZDlLC5CWD8GGYlk0yHIaOlQ5gNEKCzhhtznH+09O7y/v9RRvpibixzH9ZVCX9AHQXG4YI
au/lgEkkNxQkIBP9jumC1GSmyIQ6uarNzrmG9te83NQ1DvOfOPjVJXyhVGc2H4SdivLCaPdeIbws
fvZalyRZpD0Kia3lrljUX4f+agrB1bLNJqZlapCP74e1OA8jQiAWwgZf3jSDBNvdZLyWTXT3pH3h
sCRXdKtmR3+/A9AnRd1pE27cAL65UntMTpUfqBCMI1WNHRoMPLBgu1T1WIUlmjq/nTOyHUVoBRo7
nrue2nr5OSxVaHgRJ4J+7X6c/DetrfO54N2A89WYq3t/FOs2fuWK+EGW063pFtmPp03UtF0guj/F
JspBfyFpvYIlTO44aZwC4/so5o+iuisFByAszKOPY6P0239PHltEduNSFjMKX0WZtM9ZDVSB/sbq
wWPn4+/NbcjfCgFJaIBr0JIC2z98PwKjKlHPrA4hhrxk7ibCLyubqhgC7ss2i4zFtLPMvuLL10hL
wpGuoTuWzR0cmbnKmVRuz4bG677x9F96RPZpBCHnzgoilnLvAg5ppPguxeVpfJFD0aMcIvW8KKYk
S5fgck7ZzXd4yznwHhzygOEJJUm8juQAGCpyZawRtIdwByYw2yR4ci84aj5qrICZ2ACMkpuZkE2p
JF054W09SPN3vRdXZi9HFuSjwtbE3BCQXxslmdbdlzLlD2tjfh6JQGQH+R9MqroOqJJQ4XjhTf7r
uKIekUQHC6s/TDePKrmurJpXwx6HiTDZStjUi5m+1Y70ohQOwQ2SQpbmCCatwKCsPeTgJL0t/xnR
ZqqqdZ7XViI7pyfyoTlH/qi1+iB+XGKtNuQ9sAeww/E7Zk6jQRuHD6jkbiziAi8esCxFX4Rt34Hd
174JR3S88rMW62KgcMjPs468Q/5IdYt5017i3+ycjEgWvaaWur3v1qSSHp/bwy8erKkAQel9r9p3
V8IMWfYrSH5D4kyEQ2TYsDZtmCfiVKP+pOZz3hv5TiWTJu5wwVc13X8XQ7DlzHC0PrxrQitdA+ys
uh8xmNRtyyt2T6y9mi0YRC/6dFZhScanw7Nfw4S+qVRvIS5AjQdicPZV6z0kREbNyToGPSk1BYYF
YikWlKndfj1wLdqN7ONHAT12HIcGPgQbZwhnmEQrqLDDQDUQjb7NuGBkrA/NGWg6wEWLspIpGEEt
MUUM3BCPYWmECwObxKLN0PrCL/1QbtXxv0X2F7YCIiYr0IA6ulkuoCNyP4DsZpGWqM4dOkVrsEqZ
hlLrbIo/eSsfR8XSTfDq2w79XuyEhbuqgTaQ+gkYGz5eDimj4ADMHlDAAwLYdbd7erq6ricn2Hdu
QTxuuMtUZGGOtIVt6LUwFcJFhUiQh5kprDh60eQBHyL1pj+YAGvQCWoZ5z3kRCq8nNOeIiGT+XbB
cLn5Obkong38dOLxB/909UIdOn/+Ot8w2jIEjmsmhgsDc3/VpfRbAWmuTMFdS2VNJnduxg/L5CNX
OjxWIu26YKKT7nFdaKGc5LAq3CGAYM5m3v8l41Rc32Gva2NBrL2Js71mOXIaw2BDt8kPfIMQFLNt
oa3J9aXDVyRTFfztaOSr71CPG39IKbEmnhCUz/xZvF29xrjCi8q0NEmHss1a5wBu8YM8H6E4Jesw
wp/exYqVVX6RlSNrsn2q05TQlRjH1UfKXw6Vl+Lw1qwgCVDuG9oOWlxQ+aAJRM40ExqWxN9snor6
gHzqmA4xtp/3WQDkwqNQqofth3bHMXpKV/qd250jNWSwOfhFvyxuYjPbBisFEyiCieXfr2yYt1Pw
xUd8A/vWXQMnd2rt6qioDV+sPSIqFANinNudNeDRwg3tPvZCTz+DL7lp0aswZc5dlZwS4TIWRCSE
vCROe2gUN3k5Joigp5DVqugPM+vfI1R6L3gxbV+ll9ge8MTgiWybmUpRr/+V6PEZTGnmugvFMLZA
tm4Z9lP2t1jvY2hD4AA2+6LAGU5LCvC7NjC1iW9PYjCn845+xVZlJWbJ6JpMicz5LLxFGEZp+xxQ
LN4KllWCwk1wTap6aMYEHWHKO7gYnzp+IJUUdM/HKAOP5DD+tIbyGltsTKtG/x28qbWT1twuTud0
5GsVyK7+MISCDGF0zXMBfPPhjpxS3IgUnBVIe71ZKqAhszGu0Cp/oruxxohFyDrDTSvslVhZP2+a
sXu7V64kt7MypPB0dTRgyMc2DsrE6ZXtfRAp2r+p+MufgDAlozqvVnLVen0AOIGL2g4VgxdRy8ai
HoLhTw/zlfcnb5B79gOrMdgrFD960OGGf3PvD5r0+z2km4O7OyCPDp1tZ2GwWid3VFnPvGRNgFl6
K18rnSah+JLWuPkCvsN/D2zFU6MzDQhZzeuhJzwtwU0gcRaE+3f3AiUcQfe1G1X06tXQD8IEhHRO
ly5siOpd9UPTdKDDFbvKaadbGRiYpcu9mDIlXqKU4LP3EWREKoQlB5qZR5vttl0iwgkne4zwD/xn
+L5TIet+dEIiqqe2+o6CN+9gttiFWT7GEDZr7UvdNjC/hQhxmvVBQotL0IA1eRtSi2TOfYXttu5j
3nGbkr7nITvC9/iykVWdqTYMkdxYFs+x4sDmsAB/KSVYmBFVfcyIMjliZRipI1NHoe7mqp199XK+
Zmlr1oUSKyV7Bbz5b4sRzxP+YajGfyVNO7ypUeDFPYgxJ2HtcKx78zcylZCvcB3sJd4bpVUdrA0k
aAcLqSmUs0x3Bo2SezvKvDgoixHJDWoq2ZYFyMkfTr6vmiG2ot7j0W+eqazmREMJRitemYTOz3BA
CUrcl1xKNzdJavMhT8ODVz9cYnr/UYAHTMjREOPG92MkLs/mQv5QCGl4T04wb1YYcfs1x+/cvMDR
1Uox6Nv1qjD3csAy8mOiqhIm6tzCY/Cs2l7B1AThNsi/xeGXXFfujRVuJEj5iEK86rlMyWtsnfQb
2limsDE1dM7bpdc4BxH7QNKSEO4atBajr3zWOs8RQju0exP7w0X6aTypkiZEb1m3lOzDftXwacW2
gwTKTqscvlFEMmOywROUdj7HyNGloEu9j9jGOL9SnnbDENDe7wpZ+z/wNxToHcMmWW3bNlnqkyo/
RBKUH24KN6hgr4sn3P9hTMJc0aWcRvLOspLz6f4YBZG8hun/WKB3P6favSCrLjYu0aK9vq9PpBlN
eRb2ePN3IIcZaJ5N5ww/7TvB4SiEUL6n9uUS2U7r3J1pSDkq8v1zjdvgaPBTSw/qliIGNGugiUuu
1Z+L3CFUhp46JQ/2ZOhG5GQAaJ+jbz2ta8geCyqAkO6NKTE42VQOQQw9ovIqtoSXaTDQH5Bsqsk+
uKasGIKZvAUTK24gvTmZuKJ2WBjhHb+Wv+TKQmOLtCapGLL9vo0wgVVk/2r6nK0xrvUoBBh6jmYA
+W+TdRouwIxre40U9vwQxgOUFO01USrfelPPpxG6X7PjHduJNLlpoKF33/5xiqMV5urBEnhftkVy
1d0ws6/ve5f5bIPxrqgH1WfN60OFfCkaoufpqa5BqYaCTLFTtIjgpi2SZKy6+1xKaNAei6kKZpp1
tBQV/jljYPk6DIv4tqRoVQ7v9l0/lai/TdumQsndKL0z25IZrMovMhGNIvHiikQi7/0zMA/qmspu
PwCwP5KTFTBiawDrpfn202ZdXyhlLdYpyI+y9sPjIU1A0R1hhjSkEroexLNxaTWvn3pcAv2kDZRn
ewKJBNyZkq2ePRT6zVwNYdRRVWOmOtjybw9SP5IerwT04TxVJd5LCtlThBKbaKNV1OjHNkVB/Tzp
8dv/4QbuFe6Cf0N82ywq6yLQ2fg+Yiuw0ggSrjXFlGWQ3bNHeNlDlP3cYuMGvSlKE4dPD+oJJvzZ
BfG1fIC54VGAvB3Fm+s7cSU5vKAD6iuR2DddUVmY0gyyVkSphzk6+oypsxzmTEatsvNsL5V9/4lz
fSbRt4YrdfG6I0OFGYGAdVbeX9WPgchoyKCwKQNCmTlVbPXVwXDXfVhXuwdeUfxjSMKPExq/3e2Y
jhGy7WKDuWj2Q7gNahoNvIDD2DVo+571QNZtqo/oei9gzSYcUmkNGDUbvHPCxPKxWSW1uWZdwijK
F39TDSGxNlpbegiXRDHTjhwJTx84wDFPuN91/SNwhjSZGU912YgS1PFBbzqb0jfCo0Pd47LbdrTP
TXoDTjWBKwuOwhXGpb1/y9aG8TPQI24RaPHRZjPwNnDMDCPHSeWEHOOhK/LWsdN8Nco5zK8sgpF8
ELcld1ExB578UH/vUJ3nTXdGNwEY40F+qqDxgNY6L21wSJWb+OsX0fWTz/+BP1rhqUAe5PLBv+ja
+3t06noY6wBJTVIWw0c5W1NvTIZoEr0QdynClQIhlwpWHqcSPU3HdS+j4v4Xy6yvxxMSEf9rUtd9
I+DfO+SPwasNlMk4QPJ7pIIEoK6EFIYGKjUrxAElkJDnXQm3aKEH2YH0LCsN5rf7K9tDr2Pgzcwk
ULwqGV0uVxDG0dI1S4lqaRJ07nMXoKXc25xvmTtdTwc+Pu22CwYu2GcA4nYtMTpPXRmRq65UkrYa
sq4QpmbCmpH6rPnebhrLQcJMMLNkgbRHXSveyElWtAPoUUh+spAueh6USDmfxcKwa75vTXTI8J2L
DoVGC16Ca31P3dcdTiXYLyjE+E+CBg/HuCmDOtdOYss7uzq0UIuQ911utXhGPaWK/d+e6/aOtsbz
HwwqweJXA8JpunieblX1dc3aNXXmQVqvlK7qcFLEzNHUPH9+AjA3aryXu+sO9hYZ3Miutfxwmaie
7+c7Obmc9OiT8lJTMwvSeporAIb12ANLPGCplR4sv1iPsERbiLtrRQQUvfLRj7XaVgf8tS3gFctv
zTgboemnbOQ5sSD8VBlqyB5M4jpiBlg4bVZQ9pj3yn+seo+8qTJCFV1TEc4GzSb5Hyl0HUx48CQR
H68vhq3y76VbJZuq01JQUS3fAxMJ4dB9AEkngj4TbYhkrCc0F/zjaEP9ImEWgBMphTNT3nPzTFJ/
mTyxLiWRVVEjX1pM/4RRl46O/3eMS4Yn79woj6KiUcBC0TsERkWUDdTl0EfXAbjFhqWZjBHt3e8A
43RM+VHfcw3Tsy9gIeeXbyo36xmc3TXE9Coj11GmoV6zFWh5YNhFVm0A/V79rY+oIyrjBXzAKA7c
k7ju3j0gKBJPXMPpi6/GWlGbdwh8U9kEpXup/+I5eN6vXLu2hVWMhO0LI38ohO6kQ2eaIvrAG2AC
+1SGKxOhJr2DRFCsbUkvxCTxW+rk+j12oytnhMpGeX5jKuWCexELVSJUTa2EZptHEOVveURcm9It
DtdeBX/6CuzVo6aYsSEosbbbGqJukHBWtKeMXwUFgYldIJ7SKQ9QsWGnkJ8igrpyut4S4jt+RoFR
LqR32yd+wkkJASfZG9A+z3592WRkBNGR5C8J5IOx9Ahfz0zzq2NHuFr/EsjuiNdRtOvFaQLTkHBS
WsCkE71AyBWaR2xEHep80GNI1R5tHOqL5KrLdrsYln5+T7v55FCME3TyE9P1JdtC0bricp0IeUJ7
+U5CT1fz3eZ/C1LJoWZ7gCr65vJ2dl+ZOFeRPXZjLunIk5ptDrevA/Io4RxifJNaHnSR5P+0Nsff
iuwANNGXn5rFb07+cMFGQiwm8P9cEKP1SDfdMi+RB2MimfjMwuBAZpPNivFCLhcUjh5BMoKm1uz/
ER6WtiUhF4Ava7sm67UmNkFBO+pD+pQyJLEg63vJROocYZo3msj9RN87uTJyHApO57edffmCP5zz
W1nh2xu5Txjvzkd96oP3hlaipXjXoHB91zmq4DhyCpQNlrb+hIJWb5uCAplKvJ+IZr5+t2s1Vgm/
alu1xohMJ/mAXR3bKtCIeBh9cK8DWyopC+R6CxDfUO8ieeedPP+t6+B09RALWrLI1R9I1rAvfFYk
fxJqKomm3cUNSyJGqfx3hZfbqJIjKHDhaJpReGOHAqabrwD6/ylhNp5zv20JzDt/MRYdxfBlBoRV
UuK2wMdDc/8xsD4FDTvaeFwOj/PDkvrqB6gw0dlju6eJgp77n9l3ZKMlGHEIqxliE7DI6+ZZy4tH
q1Q2DRs65cXFtapdMVIq+tfyt710c1agg6vzfeLj7qXpSClsoKLRXybGQDOvZyvzzcBaad6ppjHG
7sBbQAKmOB/o28KYZ9UOTp3hMx1xJK3KuWtHY9/9V5zTWShz/sgC+zSZQzWaHXblXc1qWE8qSSDz
Ca4FMgANqV94Nqs8AHPkZGgk1Uxee/mexdPz8yGPY+skwSlhOdgBv9xZcNevASE9pVqhaY2+Favu
b08J3xkBfBiGxOO500TdbRGKWZrLNJx5QXRPWPHpsM3dCngsThyyldD3YhJKWorrfWpTrtbf9JpI
AA8KbW8Z4XmQ87U7Xw9mTb7avcoXLrSQqQtwdZhKZ37jqIVUHMnxjWsX/jSw+T6gFzHydDaihL/o
bMydnAaS8p0i0yowtPzXPgFBET8fT8VmtGg7gMkptJuuhYBa7oQwsATszm0GsQB2LQt/2MbSnrOc
PJFtr3tB61w+Atick/Q4/D0gpXOCHAgU696qKBvHGpBaHkkaiqqBsOj6Ta5zux78rRiuiMDkBNVz
WyGimipuJs0vO+ErUGrGKXkY+8qvWQtzbJABHVXfV/C/vjWXOECj/zG9KcDqxNogfvdIL0p6CzWr
hKphbTcmpOorEWwcWMa4fzRAQxq8zXT0TXt6JlVdRnHj9spN5sxokPsPCCu8iTenLpoQFrqi0Sfh
yVjGGWQd2j5gzVItBZFggiUP3wtXdHqrPidmcgvni1ItFX4s7xeyPW9hZX64HySOGb4lJksCbtQm
2pmBZSL952helQ7jy/8a+lVJXnBrNb00UO4oSiiwQpCnTmZrcpggz4LedjMt2phENjffBgkmAThp
sNAl917KhrJDyAh1L0j/RKkEWVwYGoGJ/OTHb8Tt7yzTAEfe6YUjy0xe6rLjjIgGyM/s3Sxzy7ol
KehHLnUOMrE9FnGXpEo4ttRnBZQNkFxhTQ4oDSSF+uEsrO2Qvjn02Fjw0caE/ac5rRGTavGDjPfo
5mbEzJJScwxt7AfO8K8jQq47NdbechhZUj92I4Ea3x3sXo0iiMPPNfZO+7RLRFxtRBemPJuaPoHE
Df95q/09QfZCuYYPqZimM4crFitULc5OPVDxclZ9Hpmzxomrac3uROwSY4Q9oOAuY5kJCT2yoXqz
cK/8hj/vlWMvHcPmNbClKwcsxVAIAVgY4NBokV9Hjd6tJ2leGp9YUFjWissV6mjjNcJIQA7KVOTe
6IzJgi3SXG2AIJxk8vVBJikX6ATXNHPElNWjTmTqoONsGGnyaIwpkp7dAjaTpINVbAOJVOlIUh6v
XREu3VNVnRYQGvr3aw2GEas3KJmEfFxjI121oYWPfxvgFn0udEcIVWjl/H5oExeqgHw7Fia81G7H
wgz6q0E1qyowtGbwOR4lSVIvW22IYHPm0rjvrgUOB8s/JWpqiXO+Mul7tZLYcqbUBEmACZbX5J5F
2MWEx6tTBn43C+tDViPMrWKegtFoNdlNHVpTlXJ7WJ7l4WSh+5Ehg9pWoohSuomuiNURT23XtYen
ELe3+7iuTOiypkCAJU7iMiCOf4pUn8oHPrxLWR0EXtHiLJKmirQ3EfVpFoiuRKRzNd1bnRhQoGgG
k2CvFj3jTnyobjCg1NYFgGA3R59eURNbZBqV0Wcaspeu/dfvkjEXaHYJKhaFqyIp7Bb5jFTwHsea
ufEJWmZsqgHZWMKvDfIwvcmyViCjg3rPWINcqduk7FFYOg6mRvKunD/+y7UgMd22bMAUT04nzN+X
5BbVWt34nQHpMwBIQABXsDNHPxyb82wgpOjsWjiagHDgZWzQGosDmKLul4gQ149EBv6G/ySwQHeJ
LLYT4tfGvnbZ8Zz4UHZE+M2G/NuzRwA/l1V5rSR1LFWCxtXaOnkPLwNr8XQwG9ihRdHbIcdtqYeW
tThVowvYkoI+UvBrlujBlv4q4WGHc2eFcPpnYaKfFdIo+koJSQ7FkiGqJSYQB8Cgf95/psVIUIrg
mQuUV/QY18uT7rTITflIyMmcmcsgc0zuNXhZy5ohbrFEhVk6Ajb9qZRAEW3V7mzsR+7tRCXpbEax
JCS5lnFba3gyy619pjWMSaTLsiYzzlrDTwFEhePG2RbtI6TnTqcW40JcR4R7uX60ZXeSScuChS1X
srSXroRHdhw8Ob7JsuS8OYTkzTZ2UAwaMXv8zPE9xr5DjD4SOWiZR51BHfXTyhwvkgSCsLPR2LIe
P26vEMyeTTtbaDKmx7TZ10M7i5NUFybwvxNeUWRWI6eC0GowGUnq94jd7CeEcUZULtHOhAvxrOHA
VDP34i9qdPH3eU0bK/Ym6lYQAJx7bx7lNzOnn4ZYPpYuSIJ6Yxi4FhNZ8D5QmFdtTRhQ3x1OX1LK
Y+bQFaQ1hQggRwZ2VtjAYQi13tF8tkLRYbW6dd8BqapzjxNJap5/k1I9EC3sg6a1NLzArPm795j5
MYHUvtxcyVz41GBg/BpR2dbHT9kbNV6hFL1wU3JBvkLjPWIooXp73B/AoX3RmN0JXXenNUuFv9WV
U/n4yMq+/Fp/fnfNmoaZ/72RgKsnGt35vEl4zjenAR3VgfFpOmyoGTROIP5obVeS+Lm9bbS6v5C4
RufJ1odIyuit+6S70MapjH6Be2ebfpgQWgn6RjYPBKS0Ujr8HICQjY49Yv9L8kC1AdQ0MBU8HUy7
2ciW0Qg4en5qUTw2mg90QlLcg/qz9RGkEiGuWTRGVHFllTTMi7U19Y+IuKXpHFHwwWAJ7rjgsJm/
pm+FCTsNKAO74Jli+qQ+vmEreMRMh5fqT3Fd2h+ypkasW/b3FsHgF0s6FjeaUVbh2MhZQ+p8W1Yg
Qxd6felSGLLLJCgcIbNs2HLAOr1OBp6S3jsOaNiBAZKLYKYf7l4RLKBQuc70APqKWB2SDSus2q3r
HW9UJIcijvb2lZn5SIeY/weWG1j6BkjAlteSktMYWtr4DtmgwuH63bro4iQArVkMNNJIhc6xKZ5t
Vz1dtsojDsJPnJ2oH1lXnDY+aW+9/TG0AhZmGqY8eTTsrIU6lAnyBlXDBG0kukU7RAzTXORzrivl
kuOMD+6kdHIFcReZstqvGPYUXVTb0r6Kt8ayrJKC7QWMCyQ2AZhaa41CRxEdQMVqopGDlshhhXFn
Vt+c0sqrO/E8jFJjAWZJwzHdSQdZOpq7+51p0qylscgnalxBoJwZlQZoIhh23b/DKGS8V/s3rRQT
qdf0K0bR8XJtN76V7kTF8zpDoO4OKBVNymcgpL2QIDxWb/m+/VRwNtYN+6BA+W/9jbwwqWhJUJeb
birK99qd2+NuuMoo07JFgRcsSGm4Tnwr/tkzQmCFc16GZHdX1psnwRZ0c+QMD9xxzMG9iOklkOqo
4dLKbwpHsRDFhva5J7MWhipb0fQwYuKGfbyUakEWSNQMXGyWymOizVrG5JDfRSli8PwfWVlMEAs4
RhbKZL9QIm3TJcLsiEB8RH7Nn4TYY46MGZznIfcAWuuGbZPSy/0j9edx7B+Of/BzDljW9Cy08vKT
5dhkm6cURTDqVgf6c40YUfXEyTi1hE6yL+SMeyrlckuB7LeqO0bw36q7A5O4vml+650v//0cjCJi
r1xFnkM90g2Z27uhc+7zBJRSTWnceSxcNGHl8hPNRfy0mq/vNkL1VvTbNAEk1PChOVt4iAb/JJHG
cNjB9S6irKZok4dTluqVO2AJBX4/TyjhMsruJ+izqXc8YiA3z0Zis4Hx196dcI4iQj3V1whd3vuy
niIR7lm16mexd/NlboDtJp2GKjYjJmLMUwAsVw3T3ae7zCw4tbKSbAM3yCtajUyMRr66635MZZhu
XxUmPChoTlCvmF83o2ppZQZHO+Oi59hyqXiQXo7T6ozaGLfDKjArxzm/rbAb8wqShKN/2oIL+AdN
QTp+UmcIIX7teRAuwsgaAOCf6p323BFonwIQi9fubAwe3bulG+iQqYsK1nxSQwLnZ0o96WR4yePJ
Yuirq8umhzR89fKLJeJDk9gKTbcG3Y3Xh3sBu867ikRGyNfajm/duMkuvb+5tGtgwSLtFx0W3yZb
PzwWuhhLyPEMPMqFv0Gch3Bc0J7M6V2V+Wvpe7qo6Ri0AQQvcJ+mUmZEKKq1TbPNyJtJqgaOYncM
awEksKNRC3jYYqHLuSvnjMWO8pFQ+soQfTSx20Y2O6HlzSMf3HDld1DG6CzeGFl7BkqVhSJiiVcz
AHtkulzRzhEa2Z7TDyPXlP9BVB6PcDe+IqMRf31Mc93vqLXz2erPb6r4ld+kzVCDPnu4uz08y708
Zgv63/qdKEq38DXMJoqBAg9ftM0uoR+SqIRDWyXLZaSTfyGcr7uliC9Vizwps7bI6rXLWrD9w9pr
RGACiqh99Y+8UzEWv3xD2p2V9sjcsMTN4NV6nNR5N3OX4ToCw3ec/K4XYktydKz5BVYarmcyKLSn
C0HUUEHtIfoAl+ARjxyQwx7CmyaUxlaJ57+0kaDdyzmXGAI5/ov0NN1O9Qj1pmSu4/sHKa+pTy0w
cCPZ6pFo8Bb5tVvH63GZWEWnzFw/xo3XamCf7ElBg/16l/yVvcU9Somjb5oB3rGe7PJjELUxByP3
wksXz1Y19s0Z+aecKEQn3Xx7mq+YFd0sPZs5Vrtk//jD9ihKMv51p71taqmtVWg+07EI/DlAFG3g
LjItS0tH34OzhewGUDnrIIcEwjiSx/u305dURQ==
`protect end_protected

