

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
VInMykl1cb/eyCcstyHEIOqfXLtsMYAK+iioa3bPNZdsHyKysw1sMYrwKEQhbdDvFZxexFV/BuR3
E2V10xNsGQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
cUXIMbq/fNZtj1t37ez/ki7n1ShEuWgIH8yPxJTOO6Au2Dmq6/c17dbZtzNOPZ13Y79JsIBKn47t
AJMl7N429e8DmdtbuhhwCbJ38cBiFdxfH1AfVZI7GGjMAdNcJoTCbcfH0JfWJ/S9l4OVfdRveiIb
dXW5fh7twSl61WcUJpk=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
WHbKIifiSnVyh9VOrHbsAOJaiYfa+g3aWjT672CoQFGtZoHYX7lHrwPeDjn9R48BpRkqqMyy5V1E
kZ30rvMKCifKQNzf0TevcVrl3t6QqBIPZj7dsFAaWjY+3fu0RTcnya994wdnAwJ92k/2t3MWJiFL
8UCO8DDPNY0Xt40qfK/53oP7zxzhOh1lPvsgCruLCaYCAr7BplNWzKtgMfwt5ZUX5jp0hTpI0y3m
TFH3zhFRvsKAbe3q2U7sLVIx7P0al79lRmHpf3nBQ8JKs1WigNl/h+LWFmAr0nyU052Sl4nQmc1V
27CTe4+On+Y4xMsv2u/myTqMuXN6bcLrIAsu0Q==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
xu9pS63o1o+cY63azBQM+vsKaznHACPUqoNT6W0vN2jhydQX/sdcqaY0W4LMPjU8g+1LDfLNYA4a
7f9gcYfJbb3zaKr5Y84jP97vWDuvkp0JSopB7FwosaQhgC9ZFFZSHrzYGBzwuhbZMni9A5RqvV2b
bQteOe3Z+NH5ROjD29Y=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
rwUkytz4o3nSG3lKXYNGBGGd6NQin1yD4vxAFncd1x1HAH4uRN/6Csj8O1eFBSdgBZrbzYpSigyS
irdheULjGWq2hoVKG79mqHugwoJaQ+RWNnILZnDjYUeFGEu0ddu39e4LQ3yMfBCfQxRQcGTVly4Y
EDooxEh83Mu9Wm4Uvi2+2y26u2oEwtbjgdJCVoicm+J7JrH1l744lVTCHFaZPWdZupXmaLsbDTF1
IZL005EF99uQ8TMXRMkzqTgTLlajCuwvHoYLTNcLy8P1f7qEEvcak6Aw3luT9m7/agpHKsss3X26
y4VegtaqqF/A90Z7VEb2715YgMpxzFEM2FzMyA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 15264)
`protect data_block
nIrbROxMnJd8IEGjzgtaxVG/hWsF9XD/owiKOl+Mo6dBBkGhZQ5uyXOoc5okIzVf9uQTXD53QjpP
tLZVFTGLSIm9K5XP1HcELVAuYIR2iCI9XFUeZ9ggdIwB44G+mHF/uJL90/fkRZmkS0g0+bqzfqHu
wCTk92KxrXcu8qMNiwvzxKCExvHqtUVY2P2otRegvWypID6vE8KV/35mFPfNJrO+MXjGzVBXpW//
+2hWwznyNkBiNqvfYPcd0bvmNuUmx2uHGg5W62dETafyJPxegM9kWKg1133pi5scq5fwbYMIkilL
wUf1R/Q9tm1gAsaN/8vLmJ5BSGfg7oIqTjRrqrLQ6bbEH80O6M1xqm5i/wSQpXH0kD9Y4upUDpg+
DGAKeKVB+D3NQUfiwsrjznzPbEtyXpQ1lCo+S7fazawc+KlnfILFTen2qW4XTywAH6MlaIRzg0cV
wHSJxavmYySlfSTiD7dpw+pnJTkykjOSS/i2C2DR2JV6aMJDhJk/RSAHS4uzkkEtMyUoq9YyNRyQ
785rVjx9qanZLZfExPpdXtnpWEflg8Sp1M/uQN2H03Bx84dtmSgm07v8h+yqrACtippPyk9TLSzW
xkTunZ46Ft84RBvroVRAl06NTRCk5tEC1mORQwVPuJBuVaVNVzvC/0/J+UUuoDvgmxXmUJLSVYY/
x22OnRthQ6aCR5DWPSdQhRkrGQ336+pJLJ9qOCUXrKYHbhkhVP4H+lIajwT0LR0jyE0e/AmhnFca
gc/w2Y5eqoXSzu9pyPB2/Py7G1l3lxmOdPpwAk2pWB3DDe2uFvCT6ZpO5v8JSOzC9m9chqyrja6a
qwqsAkwVUXtJQl15UfuqABGuvVdLh99iBYFv+yU9PinwjPI7ccGzDkO2e7IUyv0RlTkQGaZRIYrH
hOiAJjH8KDZm99PQkk+9h8uo8sYQkDN6b8U7NSVW+qnL5GlSOWdCmml4eK0jdppsRPMhnB9MzRbf
4MrmOYKr5B4hjtpCSiEnHvA8+4LKmnmgF2LjMa/7yMbwxh2eoh+kHoPc0eodYpAFlJBKMInqY6zY
nYLJ+e87IaVSfAsi/eoNitB/rCnheDPvbY9utxH2JCXsfdBHxL2jJM8D8x3oM2N1glLi3mEOeE9V
MqsStGoVXoQqT/y9RaA/cWKR/ToNnhwj1UCudICT8wZkPW/JoB00dRg/bRA5RDXx+uA+fRJSwvgj
VGzxeKnbSKNTdqUWWXPUh4Fyv8n3hYTMqudkPeJU4l74bNHGW0iQ8jDdiz4hgi0lu1ce4EkTSorH
JyGrHPLQXWFx3FioS6iJSsa3QQc6eHXgB3Z/p5bU8A9HOI/50WDL3C0pIDFPUxzPe8PY3qGHgL21
RPJ/X+20b2VkLFyD9j14TwpAIRgj4vxxjntHxykexYkKISmDY8omGYv2eECdKk8FHTt9uykYyGVo
KrC/5sHsQ8nj5S65ZfK/N05VCVBmgtqH3c7mgyNJpHRiatpDjouiPthiiyDu4fknP97frMn3CzV0
WzEvr4RPtVao5VRuWbJIPE6rXJunUvfLFETGmry1q2+2aJjt+moeaaw4mYpnbxuB/AVrpVS3ZAmA
bE39enGKWPsB/6Og3k+RA10xH3zuYVdduzF6KGmOliTjcDj8O3bwHY90dZ4e2f9XYZ1b1tRuRR+D
Zjn5/reFtmIkTp5PQIAy6nRmF3a+1wusPNuMl0YZ5Vmd5/WOe4vJkyA2lBWb2wsuGiVu41QOziGY
RRsf7bHvUVdBU326Oo2WiAz1T9bnWkt0SmhfnlZyFIGkcDZW0ClAk8HbNjJBXOSeGdv8yn6R4FYW
dCssEzRYTLBUCBXiWchsMvvCCHBuHdey5mIasQTuiJkuxk1VfqaPoeOzeBtEt6WPhX1EWv+2P6rW
FchdiQ/q0Fpnf2nGsaW26wk5k9wkC5isyG+ACc2AbPF9J8Rq1iyvnXvB3hot7oZYawex/9Rh7v9h
+fp8/qCL6vlBuvA4Dx7O3NBx2FNRmMJfjUkSUCdEcSQT3VJBqwVTQfhLRZ+xddaHfvUy4AJlYR2k
nimU8P030qc4/2KRGdU7TXUT+R6rVPtUvbNomLZTyLNxKz0FtiEt6EZlEuGHT2icRig27YcHslb1
wXyr2QKuRuZDO+1k0+QVendkCmIfY0HbY2esYNCwk9DCT7r/dRy3PFmXR1Q84r+d79ZcHuNlspmM
ezl4OaYayCephHP5EWJSv+GLSRUBlXTsLf86yEhjlxjD8XXTvlyKSplGCRQd/GYJCyX0QFkqQUoR
wvDWIXhFr2fCMVLcbVHULc4xJ5X4PBqBiZqHw/cC/VBRwsU0QTKRCWNNCWaYh1dB9nPJdd8pOd2Z
ac3LWuCvnb7qBTkFtSVHQyJDZg9tPiWe1aL5cDh4OABcPCsvAwVqi+30Zm5vMVS9goJlUaICb45O
E/aXa/2VNTSrZ2s/A/+Cvf2OiZxKN93m9X/Ozq36Es0xGEJ5ybvXnVM14VmVxwGLnXzuF4V/dTfx
8Bf8/2CfmfpFEjW/4KM26wgJ97kq4u7fvVq0xNi0GhZhTaxbJKrinfUKONBf+7uArfVuzshAtCr1
pQU2kz08dVJ36xJpC43ssSFNc83cFJzoCu7b9lYDm5UEE9LJ0F3uwf+L5tfdO529RpzR/AHVq197
vMLu4s1aVna/rf59EJxxoXRR2YrNvpd+wwx4+Y+AkGOziRxyAtiE8xBm3NUFPBYauCT3uUqXnwLP
iripBv5bW2OcrK+dVyhJ2n3tDdjd02G50PPmM+lrCOcMrHw2eHZDfy7D7kbnLkMuxvtUJwbLfLHz
c0mcF7h+MTNK6N5Ik4Y1TM/AkqyGzsFKyTks5qbGBg39Qs71Cb3Og7oNH9aiCwnNVBczITkunHsx
aQBsBeg7/xdKBE1KfyajP6UupCd18V3GdMXSr7WCjHppaa70EPrIKVJMeHWmHpHYwCBbRIjWtau6
h7/Bt9NFYG9fsi0QP5l92/TKDgjmV0CdKqQZd2XCFjHKFdPIOE1iUorBzm1SAIu+f5NlHjvWMD5c
OBVT0CWu6W1hrDc+dh8xdLvVgn7e2QSg1+GCOMLAfcYy6ERCHPj40XLFnNAHGEO/hR9QsuUrO9nq
WnUO9PX+e9EeGxtGB4R0hKSlVFM0lHYaSCnA4NaNS5JPUi/iic4uaeHoTZ7a75Ce9Bx/EE3FM03G
hjJBcttqWiVaqOlhBfCHcmJS5117TQyK1BugbVIt4sVLYSKpfOtEbC9bRhZgaysGWU/63WhT04AJ
cQv8DyqIf5duQVa6AyMfK/OnMSeFBjeip8o09LsGUD7nCBRDonJ8iLeX8Ny87bRaakeNVcFMP0Q+
CKUKvrlaJwEOuMBP/VBwQLn+1snnrE/IVTp+aNaBiLfJQt43nr6L82y1YZikFEl8CdgT/ADGJNTB
/I17BcvaSsroKhbUJq/YeqDhhTNPBAVSV7/5zED/p8GfLGN71Kh86o4U0GH2fs0ta+9hYBHUY0q8
VMUupv/GdkUvZVYWvP9x1RQOwqZ2//nw6VEEwIeDnnK6XDm70LDs9NHDZMTxyq+GdVLyPipOYfi4
IpYt4ILvgarwe0GHK41SlYvpdyVQCiTJGHPYFxPUnvx/lOs4IeOuY92g0ROoZNMzlKYVF7tpmApQ
a65hAfBZQWMH8aClZCmX1RLBpMtD3862Ug1wXyCoPxakFY7dsPiccNFrYApZVDZZIbmBiwamCIka
euSpJgmqAL7iAgmXIuya7M5K7JMYaxSO26sTtSACCxCnZc7Z7hxOlQAoUyjasEKMa5eS0QRvJOkc
T3Ci2FZQHKuscYsfM6XkkgAk/vfG5YAp1H8/DDjrrYnDzbOBaGwQtXN0a7wcgmzBpen5OLEkRSnO
16yLV9PXhptFBvnMnTv798v2WfTfIEiPNIVtMUs6FOgu/qiyaT6TMIV8lXi8TItFPB3o8H90Yf0n
g2qhaSTYDYe2JrEqoc8RHMFEAwcTQ0CGnbijtj8dGNC0aLMs2KtRTkKv5Du2KgkBSAfLF7nzu1Y2
pESB11bLo4v6hDixAtEc0+bQMoq/mFQYy0wMD2u7cvGQSuUSgQIgbEshVEnCrR300cA4x35HYxZy
Y3jRSqW+ZXVuybncobNBVf5vZvmcDEjhVBPlTXoAD0zxqtXp/GIg8nD2o3T0ZUvZEdOejy2hosNm
Yag3JhnUZK5ez9hIOCqi3ftpowBOj0sJGJbBA6Y0MfwTDTZ3xl0deZzsYDyY8CqTcO17ifDTyLdd
Nry2UKvnodDKQ0T8zKP836mK5pf9fUcyoQOLvUiSk0h8f8ZaSvlek3/1HnUFHt02bnUh+RgB8zKq
6Q4z2E0oAUMWG9u2y0jIZYBlHAiKr+fDMGFgtL9QA5I2J4i/lXjfNGeZ+uyMq3QKYWVlwslE6TvD
TBInUJkDZ7GuVyHbOEpW53+dwpExYgWfaKaI5ZruHXtswzroTMIvadIBxEHoN/VmmIAW5J3n5GY1
EtBFwcfO2HNwK39x3jJ+orJFlS7C2Gva99p9nEEUi0gdL80PJZNIsuV0M4GOURzEuvfO0eNHqFZ4
sOu0uKqqnxHDposoXSD2mejvN2gx6ZQCYaV68xvEwN+X+hgicYKQGOqEY1byClkIKBuJfsfbPwOu
iFX2rOQHAuOidBw27sEqlEz77LxC0vnSuBBpYBHsukoYlzF6evGYIWpdY2Zq0YCSoDJSrYLzwj7w
A2/41MJJzwF6rxhL49AcPV/XUXN87lUQMiSyZnwpmKUoeNs4j3ybqVgQd5xe7Vgs0A8IyIS58tkK
zLrv2gjJnbZzNLMBcXkrQSuec02neTGZC+lvHI6irEOpI7+l7FBpUTH2sjVzOCxGX501lqYviloV
SgrLw3HYvYGBBRyM2/OD6KUxhi1vkTzxGWTsdZJ8AYm183g/aoi8J9eyhNJaOtVUPOGHGRR4Kv1g
A4Ks1tJ4Aq4pUmaR0izlPBLYyfsxjRw8U9rrrW6XUxVhZZ9emvKFBWt2xh1ntCoFpLKh4Ra4/gvi
AxQcC4JRyMAcTfOffmfD5fcf/TQtKylQjbMGO1jN5qArcob7JkqFV355L4i5OWtCHGqlvSlGA6RS
XuVfonsOwKTyJll8/D9Jw8fQZ+D9lZ004Zn+HpfGLX6tDRDaLZc94a6ZZ+xM0fYH6BQ/XjLt0w9p
CkPsNUTB8pcDrMJCVqI97yY4z+mk/CX2CpB0JRVYFzIICuARvYJLS0dnEy72bDyBDandC7iDLWNs
MY0evENgsk7YGgRUJ553mx++q/e95K5omL4Zb/PbBFfCvI5hg8FU2RMbnaDD+mvXx3tjY+LRBZyh
MzCeN6bBRiQGaHIXRLiD9coiOgOkGH+PHlMhiqlCRFvmjHNKCmc4XczBeCKumpaupuGo3QtJEsGq
YAomupvgxnkVXdJXldZcCP/Pke1856/oT0vsqHi1F1QqwB9dKjtqWC9kICQbK1T+NgMekX2AWm3G
/Ng8OvvtWjn5VAihB41gzb/5Xeukwiul25Z/rmE+CxUwJw+nmnYW1FYav1JdOr48Sch/UDOFissV
v5+6y68WrOtsagITcc7fWya4mQyaNRxZJsma0cdDb0YZbMbz0fsHPryNHBqQklHctvzZCVJdP6am
XnQyvN44KqBSZu/mncQFAsgUptVRKLykvy8f1zG/a/Yvf2Pa5DCePTmUio8BF/mmnaCsnL+R7PnU
OeexPkNfqusQvBHrzqk06n044qtBJUNurTw8yPak36IuTOPlCmACQuwnCXFJDax3Q/XDIQZ3QoZH
PBTDCV43dom4apoUltXp7mqShdkhYqYpZyENB0iiHbPG7+KgzawF2wH3v6QbYpessBuz8SpPeoXs
QsyV0E0L/mCnBYckEJTIh7yPXgIGX/YyNWTGtDr/5oBOvAQprwf/jOa8gXDvTyDsLYxclJ6t/F3L
9uci1QGs0pePaAnrtjURD1RESLENyKfZTw5IDRZB+FvAEFyF6iicgwD2W3MczT1/DOYbXVykR6FL
Y61BaP4YAhpRFe/mo0L3XeZAniV82v08z596UYDjqM6s32SpaeDHe07Rq5TPohT2/eFDwLCJokpo
2/RL71hVl5KLcMA3px3a5XeQBjR6KWlIEObPPspPipQtAdvuWJD/VN4mMnfYLgEAv/HmidU2ujIB
h+hTx3Hef3HIMGigCyVeiSOY2g4BbOZBsTtESHJ1CGW+3GGg5ilrbaRhyNJJ6fMGcj0UP3ehCFJA
SKSxdZe1tC/xFBNedBhzsW4PqnGETqdOWY28QRu77YAhbklrq6NsBbA9/ZwI/cvtZTGjaExfCdQ5
tKiFHZnJ1XJqcrq8UvcoY42V3rjjFkABOK4d6S8jSlA5zZQoJpQ9KsIE378qA0lQXFRCETXTFl/4
t8oyeR0EFPu+8OR5jE5+g+XdIXNyDE80LS5Xae7ZuOK84UPEaI19k5ip+oJvDtz4pH/HC6038ncC
UR9xUiRwnpZT8M1k8RCpXiVc4s4/HKFa9UV0aGmKWva6gljaLkv79BTUrYheAt74jMF4HnWTW4BA
5dbOXqw5Gr++k803GENjGbGDn3tL9hq7slsW5finoaL1KAoJo5uhBbuI/Ku524IIY0qCD5teqcDL
qGYpQziwcdhMsvRwEfP5CTV5oKwoydSw9DzmQgWFKG/L3kzGRgEiZhqk2fza72wFiQXTCFYqz2Y9
AlLXN4EheJaQ35LNhH/gBHgWUppOaM6/TfLGHGsgj9rilSy+mX+54h18kG87Tc36oPtuWOQztE4A
4+B9loaLt2fGCUw/jBMJFo9lDlqjx2Yl9zLyTGiEbosLwCnydq3yPVEnv1UB+Rzo9BCNZD5hbahd
SCOC7A46MdMNzUPsOCwBb3YcDH847LSV34O2da+7dfqEaTJfGfHuAM9e5hZRI/yoJgLJTTMP39Xf
gN32h+eU8QWZD70tba6qB5jkrnbBZH0HbSn3cCn5CnQSWrJdkmj01nJLZriHozHKc5YsWwPHsKri
Hz7pfEJufDodI/CyfIAqPyWbXLMG8sLzfVP7BmkvVpwn8NP1Ks9AiuvAG+Hl2m90eWrjF7+fkfGq
tZ2ue1jVyBUTClQ9cT5+GXuT2GT2EvNGq7J98L6ZRBIL0YzQEsLJmtEdaMvOFdUEa1YLpRaCOyqa
kw7SteS3GO/2hkz7Gqz6kWsd5eobgUmgaZIJySE8s31KQAtFXwamyKRwXfx+g8jglwZ63PumdylA
BGhm63bYqxfso2RmyqkGfqs0yzxq5nwuidQf6AW680GDTBAFRaBB57/ZuCNXJuQNXT+ib/ErmTqF
1lRp9kficoLtrkcgvjAdrsPQ3k5etTkXhprZyPiAGR1CRqkKBKM+gDJ2c9nf5eIlUIyKLyAqjMha
JIHNdH+gpu5PMgvzLK3YGJl1rlfV3f2ZvZeSlJvxF4/ldp9qZI0o6S7K3QakqS+fkF+vOW9A6dev
he9HVk4XpJ78Np0HAYzZ5WPt6bPn4tGWoBkdsm+G01a9RmGTOZfV9hdyxSX+FG33TVWfZ/xK3LsS
YjE9d8RhZR/A0QqO/NjJMxvN2/Tv9tnmbzMhKmktQyGKXeoRq1jkhABifqqWejHzlAMxz4utkQlh
OOke/3jwP09PZxR/F2JgMwVT77strQHAHrfQhyHMw9F/g5JWqs5NktljLx7Rqi5Z0oJkYteOxrzS
dhzGG9z1hLMjEtdbN8J+DVJx5XcQa03Lx+fE4W/fTTHWWYa/YssGuG1d77Yn6RBaA0AHlj0lGbXx
1lLuMXGCXGSDi3USRV2CIgzjaSVSjPv6c6g8QfOK6XVIBTwqazBkE0T5eadB1JE5z8rOYd8+y//0
75PeFrWW7hB2NhiZFC2r+29vYsT8/zGsvM+XKTGqzjI1/Tri4a4RA9MQ1kyNGWCf3XHLNFRgoVQt
lk4PeK9Tl4Q1d5zWKH+kUTnNdA/fX/0zsTQ7X4cEE7nSv5mK1lvzbtbvgDE2G1MdEUqnHpgNHFT2
Pk8B5vdqlt25/YsRl/kij7aAQXzfwaIA06hof3FxGHtl2IzZn9fr/zy4HJoltL6kXeT2o2Gwg4v1
YwfPYMHG8ooyndhquUKU3sHdVE7bQ8Pd9wXWDWNVf5jWDkpLcdNtVlbVZKF5KX89doZb+D0dpnXm
TjfZOw5dYPM3YG5qm6Bt2E8ejmwvuBWUyE3whjEqT+cU8vG35bVmGjpd9sz1+LchVEZCqiXLxm2D
IVEqwjSORuH8vIgekue0mf7XshKPb1F/yrwcibL1VcewbKZHobRevYlD+5x1e3EGRzc8CZLzhGYW
1wadt4oc94R/L33PIpvIpnAd9/5JYpGkuJNSeFhbnh3zOzrp3drVWFRZaC70PrqmfxHGCvcu7f67
+d8vbNlsAVcGlUbBq8Ngu0s8s6WjFIVPH35tBHBK/C5vVgPPfHwK5W2cYgO1kH+x+DAxVJBFAsQe
ht/3hLF5ZLBa32NSHwOkkdHeCTStxGFOGR56NLpavchNKQ+43DLIEsmM2Gvh9NGKm2iM47Khozqf
769QPSEBVDaQlh359221tWZ795L/Ma9A3pG+jrbVspKLtFSMOzY3mXTB5qOAKC6CyX/U4exxAkz9
RHq4rt4HqkSUcNGt5AA2uoxA9Gx/jpyPUlV4tXbKp6WBG2P8up0jSdR4B2nwhkDLBCt+vCncj7S4
kuc69ByZNbfvE+nTuZj9p5ze2DHdFFEB3QKeucgIsrXdLok7PdznIK7ZBBd7k2Emya87fhac1VHt
PA8N43B9MtmNggPYH6U5xhaGneGUTm1DA2Bun/0yl9UJOc12xApD8Gm5bQYLw3x1/OzPJw5upUaA
Zyb4h37GDMjWfFVM7TLvxysVP1YaI6dpA5GebxhHtLJKZ4tRIwxh6OnpAnsndVQmn3Z9avBXgJaA
lRlNc11FhaOgqVn/WlU3/YD4I0T02oPdwtPc3PEaa79GdRWVpd+umLA21tQ0uUDcvsY4n6vJ640l
1wcf52o+JgPqJdgMv45/WumPVtmHyllbBmW4drj/Z9CIX8khpLSXz64ypurS1hLXJ0TA5BwdHjJ1
yDaQXSf74/sHUWCLsq55EglyJxBCbRETWQJIyQWvm89EYv8/uZzbuR4BWwa1jUkZ4YRM2uNgUcXg
hxJJRwOd2v/e4z8VAw71PJGEocBGmS3OjsfwUh437IFpwreMuIYnxwZS7wgvQuZTgKrqMuj63cd0
hsJFFj5M6v8GJ/EdDQjPVAYPjQTBXMmHttjZRpeaUkt9WneqdWZIUzYxWtMa8dXV5J/YqIrhmrRQ
OXY+TU/PnZBAUoVMcsarMfcp+DbtC8G2UDAOWCACYanLsjoJHoyXD6zLT6B9ZELnTTNPUzYV4lst
E/LJjhz3By+9iJ1KAhI8XpRQ9aqNy1LWSeJ42OCiapz6JNMyDghDd4oAmbzvH4zwbuYg6A/GHcgv
pQchbt7MVvlkGU0SRWapHaRisv1qKntK2FAWpVocoqBM5zjl0gtgNo8Fw6EV6KKjPktaXwQxEZts
UcZ2NPoWDTUpYtkq3QEIl8HTTNGo1/Cu0VYs+jcI/Ny2cNsMpmMgZdA10pw99kfP/M0ad0W0n/fq
3+6lezAQuYpFDHgmv0nsm+u8K3qS0Ql7B7aFUI0gRuQfKO1vTyC9XkwJFpZi/brwE7F7esXLgoyU
2TRwfDUmotzvCtR0b/8DHQIxJaLTl8gbhvNk+EBFe+AHehnU6yKTAbHd98e8YtV4r7cVAkqOKlo/
VJGJc4aH2P7ER6DwykaFGqSuaJ5hoGTTgmeZF4nh3AdDHRE/BiPx3dEUCwSVWjdWMC/5zmLaACyA
fyGTN5CsZOoYaBvPRVQEH3VrK81awhlovQWUDO7HaDBqR81BTaXLUj4/ieBdDFDdPErDI+cTa7YM
RwF6Y9ki/rFa+RcsCSOS78wDjYqolwdgcJEO49oy6/jw2arx56+lXfm0AeE1BcPSlQOSt915d9eK
9LiXyF6LodBr/4OZJc32uUefKYwhymlLJxG49bLvnRAM4PyDsCsA1CyZq+b2wEmdLv6BBIPWxWgR
6LvoyBEIlHVTa9MPforkWUC8soDwKpMdAwqEJ2pzhD7giU8bQrjyb+aLFtUDmXRsGz0y1e0GnGvv
iSYqaaT695rUYdykvKT18aH0sB8XxlTnF6mWm4NRKicx+myORNwXQ4DMBUonwBrtFSCZLAeBE4Zy
qIXka4KchHLwLFjHjt3o1qfjSwj8tuQTZRVJLqvxZs5DGvcEwtnFaFk4X9yyXZOYL+0nXA79bY4K
MAZ7qKnDyo8iGn5VH/g43oqKaaEK3srnGu/9VgjloQ/lo6ZLI5V0aP8pEK/bG1G2oo3q5nIIEzsn
O60d/yOpB50KyHUs3g+4/SNBQHa/Qja1BUyRrHZIgI/sGK4OXIzRk12PePKvv0iek+q6HjX8KfVa
yElQw+Onw5jvb2QBSqv/BNJCJvG2Qe+Es62i/5o6RKGBOCUgyjlc+GjTJSldfzSIh6xjqSIccEVA
iVgip4NMa91pDGAOievwEGC/8Sbtu22FAEM4/1KpC/VlFnDlHHhzzu0LqylP5pJx3UE1dqHnkhCy
j+D9QY7XYoAxyYgqfCqFqHtKcHeKLcN+Ucre+dYd8XNA/5Wv4wxL2cDioANjENEzNoJoRoBTYmuI
YlTG0F+Exh/+5ZYwXto5MyIo9ZUVhz8jxp+11g7u4SnEQPGo3f2tqO1fb01R2Qe5gTmEVRQLiJSW
Ble7tenBidVo1UNA/XyK2avWkIjepzveGQLN98eKahm+CaOGvuMdzImuXOwpMj1m2kdZtfxM8hHQ
b9o7BHJtv9aSVfGVpLzwHzAWynx4yI5wfzun4tJltvrBn5cbn/z8vqf0AvOO/qc7wahfUkPoYBtV
b35Dark79RyIcleNKeMS9567z/0T06ITjpQKrzAHmtfehmr9ye5Qum18c9xdynWYdUYRIVX7m5Jo
MiUpJyiq5I60w089lCK88DVePADPfVrj+k7rHVC3kn5wfjjKRTdI24/K7aTMaD9XjMQAGHa2uC44
NBjKVineNCEHEpAQVmdHjvxwQjZSsIwjZlN5C914xjCB0wU8AwGPGXEwcuMUwib82PDtoAEXEUFD
ziaq029RceHJqAiSYtxa8UqKiQGmsOWODr2YVOg8EogarbLEHhBBeUPv1IoXpP1zZR35HVMjGh2f
ZA119l/Nc0Tat0crod4VrmSet0HzTYgsyA8rBtsorTYzZZZKV3gxHf83Iaym+CdnNU0RFuY8rC+B
xrAGBK+GGObplaucjNqIe0Bvvh2UJTn7usQQBD8JmKf1rYgIWEvHb3ORgg4fCdC7jB7QKbgWE0/7
64pLCerULsn24iXSSjPY6rrmB/akirI8Jxm+Vc2II4xH8uO0C3ColOzKgq29GFVNJ6Jn1INetipP
qjg+bX4GRiLlBkShqBDqUNVzV48d/+sEeBmU+wyzjkNU8j98Qvou/c/APRB/XIDVuuZRp5LNhpdJ
Pb7YqWY+HZuRwVeMZBFk0PwqrRbTW0QyyvDuPxwmUKk4MZ1ZZa2leLM+wVa1FE9e9Hv34VbhG06c
ajjpUMpAHKWmfRg8mc9Tbw5rpbe5PvVtk+/nbGPfpXR/+m+IW2ROWqf7bOC45pDjKSMJdzedWldd
bKd/waMhAkVpO0PeQS1r49c4n5xoH0uxghSORjv1H5GDsGj6TXODLxmt7CZWHBOU3W7NUg/3kzeR
71V3CsKenx0CsmJyXtIgNrKdtix4mbium+WBf+knVUD/XE1T2KV0W9iXy620lq+kSAIXXpTsViqW
PHnEeBoHiOomqoVumZgINZp8mZfaqtQmtD8iIwgAhjBNXHuimal2yDHuzFCCnbtlkiZ9trA8VIot
EfjDp34/A+pzry9nLtpyVThAT7HcP8H3WqtQwjHdL4T0L/o9rlSfRSINxy07sXUxJ+A8sPC69U1s
BPTSiOEF2XU/0PTUYseHhbyr2OHR0dEP6niYtyKKmvDPyfXV3BSkQWpka1bhPz1/VDm+eNO0v+2K
aUeSc3UopIjjEQqnScYtTS4F9AZN0mWA2JiUH2tHnrdGkaEa+3wKALzpEiUFqX7RdQc4DVP+vu+V
xLH2pOw6vYp01mdXN5YR6wO2ly2rz2W4AlHe1RpVJdLQMBSBEnGzEoDiATwhQkpVpZKD9ynqYFRS
dxYYfKLgYCP601SEY6kJMaViA3lQZNEu3iH+O7cpb+QQU8j8tS0WteHTO8VkBwXCOjcYi/dqNud7
Tdidhas2AEZvb49ocZ9/3QYNnmKoYzKIacYrFFLKGncfmEU+v/GGaz/rgRRcefiueIG7AYp86Jxt
htDLQXf8ocMzMF7JctOI3ULR4eqK4dVBI9RTQV6xnfR4E42w+c/OzMTkaCUeCeDJLKPY5nfSPUHi
43Nqw+A7+LsmW4QP6ibtnhkeqASWvth+lBV4TS3uzeygKUvMVMtwGaWcGrffJ2ByK6W10hKHGROM
adWKxAgapGycpV0Y/4+uvcUDcpdVnzugWvbmeekaFPhEH11BJDlgjbgEEYafU2PgOCqIoYyyF+4o
SkoHnZ9WSlkr8FZW7tR19+CVlTowvfDIPZpAsP9kgPa/SbOtp/ZcgV0jDiDVewO7xs0jPZlJV88k
RvfpXhkz/E78dSPmPG2qyrXrLfDj7cs2ESOhYsDo+wZiGJJweSRAesnMo755w6Bcf0dz7Duc3xKa
nogzejzdHPkySywzFp9hqHBEW9XCErqz/rZO7zTIZyxkOc4thgGJxMfRlLdxx/vy2LlqgY0jMMSR
V7BRQQ69DqeO75lh8FUcmIIcw89VtqKsIWKWyw4oj1Ahh4MOdg1/gmPxL4W0raf5vaN8OYNoJG3E
QwPEBzdg5pneMMoxGGxzoZw+SGjQp/xr+yDc80BKuX5tcXrH0HN7xJulfh1P16GwIqfv0vqdZeqV
DGWvfvrcwiRHIX5hcGQzFJ71h562RTfq/1vHSagns6QbKpSkQVgEmjDh+F4D3uifZ6cGL1wIqh15
zMpl+28/SvBbYH6XJrTbo6RdZNhZ3tP2nptLVTkv/RuEKYgcg0DHnBW/NxeiSuddeoyd2QEunHcV
zn4LadXupqdciGOly2rafhKa0UyXsCiABs4mnFjaTZDJZAmK4c8bS3vM27z1lB8RFl3LefVIDYL0
3PutrR5BI0TK7PUZarVDrHmlq7Pz8nZ8Iwz7j3RukDUz/sOiu9O8X5WSvbFDm5KB7UK2XoiRlM91
Dtz5JtQ9xUKvelWufMGZTPH7O2sEsjQRQBffSJwzhd9HaISc9KVwkf5McBeycMS6YNqNTqFJBY6G
u77itrIXiZue1YKrrYMJMnKXdkdUJklE3XuPL3g7dE0CEu04XkzX8JJ9ObRD2humOUkVKSxPrAd9
BtPiRER4g4HzLamqpjQRO+/5QnO5rF2M3hZN/DJwZoqc5GjmGkDriP2o6+cveja8V93mZd/dt3G4
3Vesm+AL0zpxEyH9gEClYZRvA+uULQQPlqglCMrbUsELL0RJSbL/+TPIShqbx99NgHinI4jhl47X
vIoDjAjpRQQZ20kCOfX2ap2HefLUzqP0qxjReVSogWp1Uh+4w4vV79Sxq7fHdH4zW3HWuKtpTyyv
P5KkYvIERZBTbozDO9dMkEEcMsqLtuzYLduzBVhr4RkjTfCeQQhPR+16f2doTockiNwXKXQQQZu5
nC7eBGrtLKv2B0j/Z8nvlY2eeWWeKEHB1UhVKpKoGI0YhUpSKwuT/dDvB4IoR6CI2ekWD2g37k6Q
BwudlhuOku4Kgklk4wjQn7x8rSL9j/e5Qs3h6b1PwdVfS0qeTxYalkD29zMsRoHJM8H9vSRz2kRa
iRho8HjwJmysnkcl27lNf8gWfXqzMbXI8iGjf/KKZrDjajlL0yRdW6gGVputUyLR+GftNa0hBcPq
7ugTLjTsfo1AXrnQ9bfHpesDAkMFQL1HChEvDQ+sn6lhw3rjhztPU4/IA83nS+ROJSGcGtemSsi/
PXWHgjK1Eg1R+72h8w5ZkzkgMOHE89w56C5zQKUXrJTwoYXbJHn/B6ytkzVrzJenZTXf5maocy9W
rqqDjxtqqMgP1tUf4tV6yb/q1JKR/C6mxOpv96vLIKWNs2wL8tKqBDOIZhdxfF+mXZppuw3IS2RX
/OLbgTM1aBLnrOlBwDGZ4MyKQz70Gl+v3DV5/orZ6bSLP0pZjDH4VQeYw75ztYri/Vn/BB5kQys6
JpfoDqvSaOru2tTTinHPLO2b0pNcwS1MMjEcbPg4p9D46yzGGrzEcCydIkzcm69Gmyrq965Swk/o
Wi9coLA4eQ0qU3aypUQbCd1SiisURWG2cdCYLNvzzpgjXwKsvRc40+rSCBKrE5EgBNnjpVyX8HIu
1RnX4CQVVcRSJHgVgEpfNQZMN6ON8cZT12DUSqLgoj59N1FNLivJPSRNNzzoQv2x0xEy5mKM+6ca
gBnHGXu9iAYtNdeUjrSPq7ZkzCe47q7WvhcGQ26/kKKMzZh4glQgWnPSx152RJvrXPGaEkP40VVc
MvmAc/pWtuUS4+6Op4a24LdF0HGY6XScp8QVDtzmtzNX6uJnrgY9J29N2OvYeKUeLkLKUMBfxSxz
RtTvZUjP9IKnQRmUN7b2HDHI9Xdp0FpYHXtp2btILUo9JGhDULB1o476t4fB+HJMfLumyaqfuLDi
iXDU0Zv5KrkGM3oGwNjV88/HT01OwGl+T28Qd/i26vTBSBlW9Rhw+UdjsWeV2KBo+CSSyf9s5hWL
JhpegwmM2ZXqy0u7lUhBXruQn9I80JtopdUtGL7hs84WlGdxgYPIvB7+jm2NimWgkT0dUdz9l5CH
ERqdMVk62qoPf3XAwZt5frv6qKL3bAW9caHkmPkNRHKeY78+T53qTSpDDMm6qHwBt3ugEDNoOx1P
5ge52d+AW1+czraGwu5YzfHtJiUnGPpZicxMp/I945qyeVMRBUyywZ6LnZ8AZ5bGB2DPxqhMCLUj
CuLI3BJbWnPKm0vMtKtRRLAh/aU0tsmmE7dBgl0s+gYz8hIVzlpQDigtg7bxYBxW2AdndsBhSJ5E
GO7GjSf/qrLKPPb7Wv7ngAP7Q3I4gSV9w0Svs4376Lt8AKNoLiBCj+mSxNLf8JhHJFOo8oIqxv9g
p7PbnKqoCqncVD+G4v3/XWXQ8JVu91gACid8WekaxwtALHu4R3bsRxGY/1bssnk5ItDO1muyhKwH
PfDKzpypEIw1Y3JFSYlQVXvo/fl1qahaZ13m0ekr0gbGsR3AKLfgm5vrXYJrPtjwPzRbW2M4L1j2
lJWtrSEqI2Rq7JpY1goASgjaBMcrCGGH9kPRbxa4WSobpJrForsyB9tAOXJTvVq17xmY9X8eroKt
4CFU8xTnaL8nliLIMG338mEpD7oChc29GwrhvUBfVbZHPsKrFa9jEZAYvph8FWvMlJois8KercId
ynu5T3OVPi5/MWrrirZYaSzPEssd7FNQvOqiGgIQ80qUDdln+AG5LioHr2cl9qz3qUtYOW3bDi41
twhbCgCsKbJ0GbieYf3lAJwzhClWN8HZyk/eA1r7XwaswHTb8kfpMetaAv3NLMr4CcDOQ9VEN81H
eT86yVspretcIdA8H7dl04ORoEU63WkXcgB2ubYTTlRoiTizZw4PMcarvWgcyqemNqRnJT1de13N
yO4hOmH45vx9tcoTUDL0UPaYvQRj2u/55wBsnS905JHPtYWWeymgmr9T3QEFHaShHWpOVfjjOqSM
ykPa/re3EXUPT76tdwagg3DdO1pDNYl9CVn1uLFnF3GEoR+/yKNbKI1XYugyEwhkaT5peZy/SY3T
5XtZ99tkuvSbCTS2qTUJUJkmnunAjsN5MxR/fwz/NuPiKjoYvibfe6nkTEXSMVnXRFm1Pjh6jv1T
c2Yos2pa3QreHlVKdOCqfiREiDvHbDnziZwMbY+1BUg5I8wtVWOtIqVTRIxpO8dqJJ/d7/ueHFIh
BmGjXKsM+yhFpYlmOEAPZzoAVJFXq/eqecyEoNFgY5lZL43a3qZQOVqFU93UW/jh8na5xV+5yWI+
l+FDvumUS4WYcZTgwxoLlwvDdEZmOjBAnrMR6aXeB4ftLg4HszC2lsQEY9uD6D7M2GxxMwJyg4X7
bYCoGxEUJBt3Cbse71Pa8emy1dIXKW+0JVp+bNl2Xr9ipxAotVWUFiAdSCxefWmcbrL3XA27P2Qq
+eTY9GFc8k5EMCqBRvpQiIBfW7SorHqryBdj2POGgIJB6LOXTmFjgJkO9EzxiS9oQhrVgIxlE+/l
BFp9D3SijLRtwsHYHN/exayTuV4+WFOXOyALbnXYhRjjIze5eJePXyNV+0l4NYGjJuQ/fj1AaNxg
GBCRTX4dFNLcwroqACRM5u6u3V4MtDPCAAUjHb/vKlmBRbtScbO+0lg5Ty1e/bNzYFI+Ue8+1+C8
uDAw+s+swPoC0hBwK+ukcGzOFwGjVIpxaUyUMs0prypl6FoVQTTklH51KUl4r5sUmmAqSTbBO1eV
RoSqfBGjGELJsVme9u6HDgF79bl2XQct0lwxP/EyacS5uUVEvu/SkxbIJBUeYJmRlQ+6syGgyRkk
jjp/vdRF1ddh1Ooba0+urGHoV8V1PzLLGdj5oP6vsqdsmGz6Gi4kfe4h8wgGZtC2ifFhqOxikyPC
xLybwC+UjIsna7JqZsXVUtj+eCd/dw46ffb0pi10w1aurG5TVGrz1GbQplhe2vLyG3sDahNRsEjt
eUi+PpLJcZhvbC5EwR9s8liwRwEGkFNCVzCUJjMz9/z7AYbL0zNqwIeGEMFtWDr3Lv10ZUZvM95z
d0MLZkyis4R2Slg7Zqeg+h5Ec9Fx2ZEyyiXLiTNp+QmEF28nLxFmftA6mXbW0ChdPTert641lWes
NbDvp7Bxsa9TWgK1/689tyrq1XxdAsCRuQfjhn1T+MEfi3TR8YTrKvSnpNKpT2GjN0U1PJ43J3xv
L6OtJ7cjQpZs6Imqt6Brz2BetdKvpwpv3aWa1gAQcMB7T1MTiDkey6U9cwuuggL7+ZeiBxAs45xZ
SEGAjzkAiSdsela5cWqERyM1TmoykEu1tGcbyArm/6CaBE7qCgF34oWDkk6S3kx4yunp5lv19iQG
fC6co645J4IcFfy4gmnPnMWnrtvq4AwWEo+eti+b3pv6qAF3U+9zxQ7ZVwPihhKGOeBOx7PpRap7
n8d7b8NmwzPH0pVdNNZZ2GR7YJZj/LL5UCrvGildpzOxJKxoEEQ9DonugLV2tDGfoA0mjcJRlC+S
dKOHhNFGB7rTVBJgHEGfLZ/XGuJtkNPjcyuB9U9u8BQfQ1H1qqtHHp1fjCtpyS0IB2jqsaNXsFV1
3LjpIfHglv6LsuE753M/HAFK+WSyRVnTkibrybzuxk4G61GjW29BUTPOC07pa2QjLN79LqpK9T4I
neOeg0yi/tZt1+xHfIaeG1uvm5GPPn+CtGP9EgkRcEiaX6N2XCvK/kh+NEehCuF0KnS93aaUsy9/
5HqPIUzQt6DvV4FUa4hm578IL27G0rai0lXX3yLt+c36syU66xWl1Cx0qDfta8be75DRkfXpxxqn
spNXlaTNffqG58ATfx/TdILu4I4so8O4ra7nhWtVEHEO79wYK+lAWJzFxxSEnIfGKYHr+XjXJBlT
W7vna3St+pYFLXcjvy6/jVJ+hoK+HheWSvzwcXxNCBtHroO9k7eMDtP/vYfGeijidDcOYcmysjI+
1/Sm0bAIfNCYsZ1RUsyWcms6MPTJ17HiHlcgIOZAH99ycsN5YR6JGW3IJV8zP/mOqSMfxAFoUjYJ
gOE8Q+IeN39/Ug0zqd0/QYMb2sYXx8Wo/0BEyWptKknfF+k3LDwpuRrEntLSwphohQUBFQZSXCjA
cjn5LwR/IMIdhrzA/97BrHQECd3yv0hNb3lJvXf7t+/iMRbnWqqM4NSYC/byLnpq6nIO0MMyBRXr
WeF1WioPI2AQBgRkmdOtHip1r62+ffJx8R9GlkPawGtwROX+KMnZkoES1gYoUpAhD250T3MMX5dq
su7/4RGr6+ProeNYqRg/dFbKv6TGIU3of78Ou2t8QKZNJGzzfWkEs+nHQhEqUcom463iWwHN7+oV
dn6UNPX9imS76QP0DU8m87XVooMrud6tCO2/tYWTBjT8Fm358UQ4zP/P7SkCROjid09ZW799T0if
i68Dy75OE5W7NNoHYlanSffumLGCRIF/89+UWLm+hEqzGYQY8ZLDaurpqyweur0KJ7mFtdSnU5CI
fFbLCCiiZYgZ8AJPq5Dv9wB5+sood1AsbCuUk0+858nYvFJd5J3fyiUgujdyMx66+X2pXyh6oSQl
U/ZAlLWwoo3NdS2zsGU7luL96v4Q7gLPc1iOQr/nMBTqgpO8fRPlpKHSa5YPLFz/VufOSIsvDj98
NL4sciGIpa8BQmiprOAriLcp2RnPbrSxFgqn2XzqvNr3jbg5F+cOlDl4yedcti9chmnMHiY3PA+s
JAdVcOBaN/7Feq8dX5jawRJtTLZL8Mlg0XXzNujifFB1yzhW1a6I0wDriFzvEnZGVpZj0iKdM5v0
iY1K3CVP4z/oZUMFQ8cvesGnDtvj+nFN9XYobVwjgmxKBM1fMws56spQxaqWgiDehQT2rX/bEon8
P2bl9GpCzti2u5V24MdClXGsjmAg1xZALOFq9bwbrDDFnE17g1GJnznqWdAWik2BUK1FFW73MAVK
f7n6u4Pe+JE1o978G2nG1UqgXoCz/2kyx48WXy3+8ZXUPdW8/1Ihgl4C1kLJvH9KqRiO3Fg02QYZ
dx8tNl0uQC0hw6hVmJQ44iuNgqUBn+I2zzdjyekZNd3Hf/K0slIu6namuzJfMhlQN//LsW1MuVmQ
K9nh9VkWmpATyh+8W43NfpX3VrKTIm4dQ55AkOdvtg/uX00rNLZYyRX3ugOhEibwEE7GCEFYnxGk
dlkpjBnHnjLWaW3/upeSB6IzV7AzdI25zHQNQkErSMxhtQmpQIWo+kb62GVahNPlJlrsKHMjwatt
z+WvNmX38uiBthcLXan96nRIhghRkY7kMoR5J697Ao0uale7uBcaVMO5HJlHEDC3sn1Fiwa2WDsd
0lyOkdNh2TR6Nzjr/YcWjEn5H2Rt3G8qzYsOf1EGJMxZA/adSMYvRKDN8B22ExRwewm/CZru/kC0
OV3lCPgioRy8Tp4yY9p9rr7giaHUaDMOH+OgfUISHwPytOLYhsJgXADT/IIAuj29XNDZuyWlv/of
HNv/edY1Rua0kTbstqHAQOF4k9tXUnRmcfdrRvIOiOvJO0cvH3X23XJhaxNPHYfygi4Aa+GdM331
JCQa6m6mauX0Y+EqiYdP40qpZ0eor+cdyMF0j0cICm5Fl8hsPJVAu2fcL+Z5rdQwlPw3G1Sn4o/g
zhQpHc0vI4QMb6ixDEnpUJkLEEgN0yORDAfwZ8FjzPeBkEnk6d0GJYUKn12LUwd7xr+xKBGWtbfk
JvyNtF9qJx/ONQDfgwG3RnKZT2LfnJxHNN9XkgFt9MfRkBY9eFeMJ7esXZpz3cENyzpzJLpb1b+C
ouSML//lrE1bjJ1YMG8ekWGfqhx+WgqE06D7lpYiykpt1OONaBQ39FA89FXW7GQl4imQ2pAg/qfF
CbjbPsyLMf1W0cWyYgN4FMQJdW27nzDxv9fSYOg0G3PqzmpkTkB6htlAQOFcB1W9AHLKFVoAtOYK
3XaI4jqC4+K0VoBr3WdlxIONWC5dDd0rDKDDEyl4BSXv1yNrajjGxWBs9tLiXo+AjN7BsEYQkzXt
Oa5N1EQsE//ueUVIcu11PNHXcf83IkNoj/xXPawMJ1H/G+DKZ1k0L0QcWB/4mX5LvAljJaakSWRm
LEe1UBB2anxw6M7wbd73KE4jiG3O2r9Wlme5+stgOycIStXRMCmWFNyvc3n2P8GQVxhxF5VqwWGH
DL6dyzAMJjk/vLn5yF9X1QIgb8FNpIt/niw3FV4m5d1P8N71l1/SOxl2nmALVkHQ482xcIP3K9L2
6VFJR3APoR/0Y0bMCTQsqy27TKQojBkvTVy7pLRDnL/XqzWYIf1UnvxqY3jGmwEIFAwvlBEax3/I
sOsW/+N9ReCYkDkeRND1/gzfpcWi4xD9zzzZbWml5rPuuZ0iLUNSOtJl0FsnX6Rv9HDibmFIq6Bm
uuWBKqAEVYz0X4sHBJCH6qD/mlZp4c0jxhHx9/TgvEHVIhzxLREwFF8O/wThDffrp9kuvas8Fm27
mgzbC49rfLlKq2WWZThaKuaetLF0qicrSlK+aho3VGpz21/wy4sF5Sfuq5DHM5q29rUo4F0HDpW7
z5z+GsMbzG+KcewQImxmFOxtC6v85wwrJWZ6z6trfbc2zwrTlDFZFPtLfDgL
`protect end_protected

