type ROM_TABLE is array (0 to 255) of integer range 0 to 65535;
-- This table was generated with mat2rom.m
constant colormap_value : ROM_TABLE := (
16, 
17, 
18, 
19, 
19, 
20, 
21, 
22, 
23, 
24, 
25, 
25, 
26, 
27, 
28, 
29, 
30, 
31, 
31, 
32, 
33, 
34, 
35, 
36, 
37, 
37, 
38, 
39, 
40, 
41, 
42, 
43, 
43, 
43, 
45, 
46, 
47, 
47, 
49, 
50, 
50, 
50, 
52, 
53, 
54, 
54, 
56, 
56, 
57, 
57, 
59, 
60, 
61, 
61, 
62, 
63, 
64, 
64, 
66, 
67, 
68, 
68, 
69, 
70, 
71, 
72, 
72, 
74, 
74, 
75, 
76, 
77, 
78, 
79, 
79, 
80, 
81, 
82, 
83, 
84, 
85, 
86, 
86, 
87, 
88, 
89, 
90, 
91, 
92, 
92, 
92, 
94, 
95, 
96, 
97, 
98, 
98, 
99, 
99, 
101, 
102, 
103, 
104, 
104, 
105, 
106, 
106, 
108, 
109, 
110, 
110, 
111, 
112, 
113, 
113, 
115, 
116, 
117, 
117, 
118, 
119, 
120, 
120, 
122, 
123, 
123, 
124, 
125, 
126, 
127, 
128, 
129, 
129, 
130, 
131, 
132, 
133, 
134, 
135, 
135, 
136, 
137, 
138, 
139, 
140, 
141, 
141, 
142, 
142, 
144, 
145, 
146, 
147, 
147, 
148, 
149, 
150, 
151, 
152, 
153, 
153, 
154, 
155, 
156, 
156, 
158, 
159, 
159, 
160, 
161, 
162, 
163, 
164, 
165, 
165, 
166, 
167, 
168, 
169, 
170, 
170, 
171, 
172, 
173, 
174, 
175, 
176, 
177, 
177, 
178, 
179, 
180, 
181, 
182, 
183, 
184, 
184, 
185, 
186, 
187, 
188, 
189, 
190, 
190, 
191, 
192, 
193, 
194, 
195, 
196, 
196, 
197, 
197, 
199, 
200, 
201, 
202, 
202, 
203, 
204, 
205, 
206, 
207, 
208, 
208, 
209, 
210, 
211, 
211, 
213, 
214, 
214, 
215, 
216, 
217, 
218, 
219, 
220, 
220, 
221, 
222, 
223, 
224, 
225, 
225, 
226, 
227, 
228, 
229, 
230, 
231, 
232, 
232, 
233, 
234, 
235);

