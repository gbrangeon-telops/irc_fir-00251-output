

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
RZm5UrZFV7JOtGxR4Pzih7NQYLp7LmPE59R/6o+hZN+ZT+nCA+l5YH+/j+E+cmHHWo6IUrn/ULaG
ZkaGINks7Q==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
MRNQzUt4f7a/v9KMrin25EUCYvWi/twJzLlDdceTmDN2GCvOURSU7hHpsmsqqCb1xCeaV7xbvs0c
MXpZkAPeQc5Coi1irNf+9eKbc5uIh03B/PevhS9S+La97Aj9rjHplzcZDEBFN6fiyAdKvJgOrOyz
87nOO0u5LoaEOeyC6ao=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
L17wVQWzSUChaUkUbjAqDK1dFxRQ9orAmYas8htY5fjqeIDtBkS/PldQL1EGRGrFVbxZVbStDyiq
iWMlaMSfJiAW0codwFWqGkqnH6YMctbqpTZdQPbprA8qa73Xmy9S5tgWXo6y3vZys5HBTFHxXMXj
HSJZBGLfj5+GGMkAkDYYBZrgDs/jxx605zYzRg+wKonRxjx8C7c4r2cekqFXXjEfMC6t47HLGKZO
Wp8oqSV+SdxjNfsxTeAcFxqhiABG1hbduxwcNIQO/0mgU7awDWqjimqvnE1+KO7vQU/MVpl+J+Y9
bwvxkUUMkYnqQG/HGWvvQ7Zp0u8+rRyDh2dzOg==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
yJG5RZbV6QsAW4khC+YjJnbI2jNRxPOtee58pTXfgJVvj12BYVsRuhi1xiVJgak8Vy8V0UJ43Wc3
ydXie//gOHZIACOddgGz8WdlyWauaZ9sd1K4GlV+vX4K5HkoOyunq5QSLYwU2X/ZYYkTAGg7My6m
h1UvByaO98o6pNd+n1w=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
QjcZeibYm0SAHW7YliT2StC14hkmhpmI1+m8klXbQfAK/yXQ8NfNnDZicIHqHpAbgVQzoGSkcmXa
qhjmF7JhXI4I11rujpUqz61fAf/3PeUiYimqp9l0xnePLlrRBeItzqfetftMnQ8hBAuI+sARuLin
j4+kHDvo2V/A6kndknmKA6lyd7gI8Mgzy1xgvua2Bfq25TZ30r76kaSXXo5N6hFVjtfwPGqnYepq
02yTg3lN97x/f3REjUh0T05iK9mOISMgvqQkxFwl6hBnLhp8WW0zJBjFvAguLZDf4CMBuYBnnmGQ
axcOzl5DWDcYTgPm/DTciq3eoilijus/JUHuFA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 8000)
`protect data_block
vZPjbREj7Zs4UUN2Pqrwcnau4S/9a3wQLoOW5JvBdL6M5XWCYwlTPmaOwhVJO2nZ+qbKKHJMc9CN
zqYT1ROcoM9BgRbwFhZ06AWIch/rqjoA7FqcF3XYmvJhdGdilM+/cme/mtId05lG2MABxXgwVA24
RyR+CtnboTi5EYP3ONoviuvEsBRR4CqlFs2OWYYof/xKiSJM7VthUVDbzylnjQcutmJsXjNh2rAc
OVKLzees5X00klWLFMR/pcckljWULJr0NzBI4zx3AxdhWlALRkxNpqFFe0UhkB5782CdiMei4SPS
cqqZSnuGeUcDtQtB9rqbN+rBUgG7u2kNOW56l8Kr8tz9qSGP/3/H0s56qP7rwpcMmV5smMXpMVcy
TAA1Na3o+s9lW/ELDybE0R6I67KSElkNskKq7qnT8CkPHxjTm4LbupMm1aE+Gc9u+b1TzHkHNd2E
7uB8251/BsS1bHvH8/SjJKhlhfnixgFmwHSgOpNRhsPHDIG1LVmiyBIEK//hMfNdVAEP9ejC+z/x
uyGt/5k6zUsUTZph9A39ZbwVjNIT8DZOdDcwDIPswwsGqt2wv/WVuqbU7X2lqSm0WqULqInyfTVc
cbBkFl7kywSJUZU8PncM/xPeGEr4BlygKbQUBJgltOyhTxeJJnWDOevgexHVjpr8LO+aJ/fiSPEX
ufR4FkDJtNUiirxARexd/Qd7SmjH4xy3tMdpyZAtxTCsS2woV28tYNtc42lmJRYJh626pgS1QUTa
NR96/D/8UaT+4CcSC6orbuuZQqf/RcTcJseWt9dD1zLjUVWGBR+UwPWyzj2IRY/tME7kcbiFKKXK
ycO5S+CkJgswRWzKLad/SXEa6zTFXFxAx57X+Roqb8X8dwHfBXp4k4MnC0F3FQqJwJ4ZniK03JKN
baOzRVIDKPpgykQDLJmCzZt1+BZzW6CFTIb+v0uFxGVjiHJkImJrrRI55h7Gwv+SNTLMyn1e5xVe
XPIl8oYwZQpdGIcy0w8MfNy78QpV0BhxtR/Iwof2P1yYmK7upItX1lomvHgs3AfzI8QwEWmu8J/8
pfPsa7eNzDFH7v9nH95c2MC4DuiQWuf0CccyUdt30m+VqtjUQNqXyyM06HvHsMEhhY3QokwBUIO9
Wk2/YkcoxlnQqZCG4LroZPnfMci/GWfgptBCG1dsoUannj1/v8Y6oykU51hniryS+3hdkuCtINBH
PSPIkL2famAIfVO/QQnFJCwzohxLW+9g5PuOWhk+MgLzFxf2SSh49mUuuf/ZizJRawDr78Fot4s7
5i/E8gLmT9avkW5Wave0st25ssq86EI1156RacxWJqlKv3BmtoY4y2k78BRdqukSIWEd4wxa8+PX
UNC02KlFZkcKGpIKqpKoxFph7zEXzBZteKBNgCdZt+zvZdQgjTAjfopyXab/XhDeEFs3FW2xc7ui
8Oo4ZhUDr3w0OxM0jXwJC96roHp/iX4byr8K4fvxhr5PM9kEfnys7NMWLOlJc3P6NsLaGyDf8eSi
/f1f0bQr6FfIGbUJaMqqj/xLP5Z5/ej4/Xbb9tM5j5b2mu0sWjnDmQw47PaneOxSs0y4fQMEufRn
P9Btg+YFXS6ODEaazhiCkuHEnccaFVa40CSClOl8H6p23uEIS4TO93Mwuz8Bh6qZdhr53IbAk3sZ
QCx9nHCDeM7+UXlgHn48hHiMqf+47En6scKK6enT50QVvwv6BGE9RMFeg2J55n0bIybmGrwzrRaO
Sc5adOBQ2Rhjxbj6UtB3x9BkvkeydYYCOP11dH/2uXf3A0QplcpRnCIP3BVCD5n3tC2Ypyko9iCx
M/opQ5Jjz0DdjMC11Xfu3DQdGhl1myGVIEkVcC60rZo2m4INZaUFCuQsStH2vFmMWJFLVaAVZ1IZ
X1XUImi+Vdij0jPIjvN/iWYsCjRZn2kk6sqA9W+FA8qelIjdYi3Ejg5G8FknT10EUVjTAL+lofHp
RwtR9uEi5Dh3+3O/uk7fSLlIJT+nxHj166O0HoV5IClNejjcjvjKjDP11xXz/31Ed32uSow9miSW
i6wvklmElcP8A9iMr4ZJ9ydeV0fjiE05O+AfTmUtplQjLhGb/J+yJ7dgxAss9OwGDmSujmWvi6rg
U3B5p8wNBbiJAqCRS9CsVy9RcT4eW8TQgWeBAUjWlrVTTpfN/Aju+Jud7alcKDtmgWev1j3S7lQS
8RaHeax6g8FeGh3iwujf0UsIG0KIzGlLM9BaReOGrzaEvvu4n7NaBPOF4W5AKfr75zuXfrtckF7c
gQG18eMbF6FdYYgMG3Mt7JRtP1hY+0tvVlJtEIG884EcB5h4aJ7yEiEdhrxGJ1tSCAi1ocY1ayx+
d2DLb33tOuan9zLlX4cACy4JjjNR4kau5zAK1IauNdNB2m1M1p0nyytHpdYHAepz/+E6FGdOxCaE
3XOS35G+tM+QURway74Q7G0ScwOShhtrMlGgXglMw+bI9P2nUBcieecORHhNCeUne/0rrc1FcWM9
HSzWpmkO6uvGm10qQbrGF/4nwx5UY4bClGs/5x4CtqrivurLBezcMkC2zdvCdhDfYJaxqZNX4ZPR
6t5+q02/0T9kC5A7h4aw+dBTKLvHR4zcI1RJToWspqECHWah2Xaf8eKPNAeRJu/cjpA9mafdxDSi
/lZhUPvXBzuVOhxIJt6EBOuYnxPspB4rorSehBtynFjK2h+8pMM72C/2khGEIO76zgRvowym46rR
/ZCYG/Sj/Ve782+N4f/eKfNIk4sx2fgqt4TJIh4Sn8rkawKdHp3YX8lmvumZfedrX4SmkCbGFglx
M+hTdGKTOhSkMSVRZJXOwXdQEsHrAOmJ4QUKffvuQ0tg5J8tA26oELUvQmGCWUTdJttZbTxSiE0y
wJLDyTFftVNYNOoLAEzVo1x2XVdEOllejLNIY3fcpme6YWklNxFvA6OtHYXfBaeB1HgjdoVBZyxD
smSSNmOV0b16sp8klnPX5wXtuiyHKsEVUesn9/HNudKuxCKCEM4+Rt7Ow7XgqFzn9y/nCHpwjpNI
Yy2SiDSZYowkdayNZ9jwdohym9zcGBwGV9ukbRcWXLA0BPle/F5WcOtGIs9RQynSltxfvq79kIh2
x6vuHad/uMJiTI3GXaWUkaHEziyEnpfZyzX5klITLMgfp8WCzpZXf4GpM9nfevO5ol9ulVDW6glu
3BnBokh9VsHBDkVuq1md/ba9fQXiJRiqxQMxBxvutALoImUNKjMu/2bM3rXSLOcWvsRz/2vvL/kD
OBFOLINczYKQxqBETRB+dl+z9Y7Sj2YTxjRI6ve51LTpIucSiPyxI6la4PFo3N/LBkAqcvGGO9Wl
tHioO5q1JGFjq38ldXsBkXfkpL+DdjCQMKtR0SOECAxV2L0BD3TwRnnVnScVPvGDlIHR06hhKEQg
lpXrs3zBKoK7160B6sJ87KOyWu7Me4zQsDVLBYwN22+9bTt0hFMJVwvDek4bfN56BNsnYuroLUJv
0K2+XZQvpavPDfPjDjRQsfj4fJq/42BrOGqlLNGUDS0QjOM4BRoJSKQbchI9WOIgPPSp+ZHOE86y
VIN8UYHXPnBDjxciBUnRufzd0NjufRPkCeJuBtj31s7PXOA2iERN/V983yattbeA2pvtO58my+6D
bKNkv7ZPXHLoq3DukZxyt7HinB0HySl7P6DonD+YZ199nINvrlaNb6/CFbGVQLnjxyAsDbGq8OV/
3jYwqlDnqGAeM8bSpNajgtdd3pRk3ynsgTm6ifLP17Sds+YEQkR1WTAs98ortgugqNCjhs4olCVP
d57wpZxuW555bjsMYmzQBR4ejXpSbJRQs4DhJ3X496fBIfYgb82evtdxErd5GhFQ8jsO3f9/S7ge
JLxAHLSUCq8VdXZxPeGeCQuGSIjW6vpUxWVgUk6wL3ZEvTATOoJuI4macgQsJhSWxVRht68/BaRt
bAT4R3jwyuGtlLa9eYzv9fHnjNR8DpOjdk1uXX7BpAKaq03J/ZUEjb+jLfQpmH2RmE4puuld5gcA
7THS/3ZxnROnPsQl1sSvc9MdMrZIbcSEzYP968CuWCZAQTGrf6qS7MUZHIWTGgE/KdTxEvkvBDR9
9S2a+ILGFwCxzjMrU3M+IPWmmpkaHrVPGvdfjyrZaMZgSEGLNhte5QqhnWIk8/Cth0MLZsRip/gg
x0BHUjIQt+TTPt/U8YdjXhbmI+dISww9QciBbCGj9xQFeiUb1ShA3Yfjj+noWC6C1ZzI14kE2EdG
PKIQfr1xwfUp4h//YNAyZB5CO+FzJNpIdRqb0qM3/zm/7j6P6lEhANITqIPAp7PF5qEv48y0Abms
gH4rfaUBAaShXosGibu2IoLf4n0K4Oju0Fd+GcW8LcYbxzFaqN/D17CArMGP6YGvZzloH5wyeJiD
AXO4+V8wxQj1frCE/KgmyL9WVevTS0ShfjC705mM2sfHqy7rFajLZsL/7MkxN1Whx4gQq3+kiJG7
1jOvR2ABul68PWCGS0eu2Z84eF8nzsFgep1VD1L0wdZuxXLWSK5h7GpYNyYYWepERmWhwIIfdIrh
CYlJCPVuhSGRaJay9HLMy6aXKwIfXMylzDcXyo41RZ8U0ngPYX6eYDCtn2BDZzkd8GJ0GAd7snST
tNYAze+bAec+e7lWMDIGgULI5sp59eLmgeuT79sJ7woF9Ht8Gs1OPeUMxIMiz558koPsaeQV/szg
JTi2Wpag1jrdfFyo0j7IDJKJzJqAai9g6AsIF/VbNqbSQbfsBU2Pkje3SOQ0tyj6qJuZs4jnf8Ui
kA1zQP/deYZgumVKAf0rPI6nWTqDxid5Lvexoehp1ZCX3KBD/wkujCqxNtgDCG7hLwdA/p/9zGnv
+10CiDEG1l7B8O7n5TY2Yodp7KIXkYWgemgHrbPJoyKlvbTa+vejFrEVvXW59ljdmc0V7+y9eLjJ
zN01Im9Oa4RBbaWfsYLmr8dEFcJ6aVAnmJpqn6coSmHZG8z7ubxWxJAUZ8GuoEce2P4xsQlxakoZ
vsxhuSdLn6qup5A30NvcU/lJ34QMW9GugqNPKMFcYHLLPEiyaGDiwtaag0/6YijDb6QT1osumcix
/B0wIP4bYvLQB1QRHPs9TEDVlMGzkvTeA2Aeily0SANLQuR2kA4Uqk1k+2YwH7bhe7j7fNSb6Kbz
SQJLL2JznMQ2xe0lsYzsoMJ8iKHVKnWQ/6iXeX2jRo4h4R3nnNAC6u8YfTrzeRHZ80w44iUF9hcN
qgluyt1jZMN3oTt2ULD8rrb4CSk/5hvhgGkBLELa+PAUbVgqogHoRrIeqHhp6z9yNWw+NRkMixxo
CPhdZtL5h7/a/uKUYSx3SkCENfTyJ4EOV4302AsH/spExR1X9Kj2N5zDy/Qvg8emJAUMzSCE1tGN
VPPxS8o7MjQQmd2GfM7Nu5vk+4Bz1KedFQj1MuOs9Sarg0KyL1wK4pJMsikzPZcUvNBn0d8GP6uu
5DlvjEwcLoMmR4AKf6QqjXwSu6uyh52QZYDyzAQj08tQhWlsIL7AGNMiFy0b/lhqhPmNI53HmW5P
m/WiBPrSaPz0N8VCTSkDK/F9bfeHQma2j9kGtncM2SeW8KGoiujMo4EoYfmDznEXlR2fH2loqp79
ToY+NmkHWJuQOs8oqe/OkT8ndAZy254HNCX2e+KJ/C58SV3oI881dB/AMp6ae6QHc2+o/SbdlVAU
Vxg65rKTzQnYTmCREnZxIP7FCkH28WQEUmhfMeLBxqx0JRmQTyVI4wyQBTJTp2gDZwEOvOGrc7GC
9nEgr5fugyoKpGW/V9f0kqLdqQaF3WTX4bwbJ1HUXAreQBeBPFX2K23CKUZe5oJB30ZST7yJ8xIQ
+09eHWQCSTKcZbToNQq9rAcMLw/zeBlLP+SpezamWT1U+h0EhE8N5EwyvHmYqNwea+2ognKBy8F+
52MjTUsO5U02LiOjMsmtxgk/ZoNxH2dz2JwgNpK0munLdexhsQ/Vf+UWvXN6qz+qKAnVYJOR+qBZ
z6tF600kw8Vt+rEMuwYNGgryNBU0h5M1RNpyWiPldw3fwlK1Lilrh4txO2ebkeLtm+wp9KE4GLhi
MFTX6BPkUQuhh1IxTxN1qMWCFBoqKXM/je5TUJVQcjVzuETRoucP3AGq3yX4v8nnAX07IEzfJHnN
fDCy+43SfKVE69bbPtiaXpLThkatSmRWDvEHvw4jNL3yPFjIsQUwOw8tbDCnehuOKG8PxL84xPeD
oy1nsgCirfiAtxbquR/yqE6DpuODlz0PUC+BelcZ8WNyXbstB0PbprgJLrjq2fSPsE5OiCEStgSk
Q5DJVVTglCePmTKqaaZ8jMrn3ajObwGgc/sICeDf49N6KZZmq6tff0BztLMutivk8Qk19cKC9dHE
HaFY3LLGi1LYJLJDRWaXnts/KYc4BpNanJzlF38VXZyHRB3n1XXo4OAwEANxCoM7VAaeNzJgEdat
3mG7taFtJg9oaSAnEDEqq/MBqdUwaICKo3Ubg7o9vv6vYIjI2MfUum5LinzWcTMx3lmFznLTzRwL
N/MpVJyynLKQS8XKGXMHHG1r8AvyyubHsUsSuO5LiKtm3pGcu7nRxcPWFHbnjUaPzfX2Oih8odrN
khr1rFTmU7nd+UMUfx8B9aBFxmHBEsHCcPaKxR/KyZiTjmwE+0QBT7a2acSfliTCxGrcVUHvXpHL
LhtzaWcvLV+6DYaUK++FnFFYF/zlBg0WLBQ5NtyBgxdFDeHZJftGBaKmreroS1WiZgTtPv99a/Mc
toC6kAj3U46KaK3/cjexOSRru3DZJ00PTdJJq/zGlIjAdteR2vi18Wz/yUK8P2Re+jvmOdlLc1AG
0MsLFSoXZIsc8Cu9TKFQ3F4RG4eC0Oje9hKpwWNW2Y2DU7bcHNwkU3dfbZYzOi4ULXKIPu9ZfB+2
cHY0dz04icHAZwSK7T4XXcGuUi5iE+QhTQImmQxwLCYlUfrlboH1I8omrC23QhhGPunJBse9/GEg
T/KxudSRcZCMGrVfwHwxnX7tmAvflWsWtbmtWN4opvK+udN6KDS/BuKtCKBNuFP2Mkd3HmPv2ddp
W54jBCMYDx9hU322IuDq6uFvYno8sAP6/YX7+kZgTV1YDSCILTGiRUUvaIZWBSZe+DBmixzoVSIT
4YizHSlk1NunqaIjeC6GR6k7VzlIDbGLFPwtyNVOi+fXaCdhUG7SW+YMVaXdmfrJkNLum1bewu6U
oRBjJsJf7oF/m97sVrLtMFG5Sake5CkIMyqgokDvGk3pFcbTjZJTliYg1e5pG70Kn+98iDOZxHjD
DTfxRfoXKEMRkrrTtGix6eVmUUbOb4xZGQd1oAgvbKW+G5EZIro7xMlksSdk9jspqL/BaAIqoYeR
UjjyyxHHfHlms4I+a+nV+K4N9rzjk3O/EhB7y7u2+aF5M6URA0M6Lw1PcfwEvVyFeX1B7qEqgcw3
RhLqDbHMA2lTPUZs2R41tMAUHggIoMePKlr/NKM1V9UoR4inu+QMa4L/j53ZD378HlNxHACCAEm7
7HDH6FDIp9HmL6TW0nJmxIPLBQWLFqllm6/xXTsL68eMqFz4qNQF8EKeDsZBw+gkG74Bo4npCBKv
hkbfNHy+kovlN9GAmeRxzFH9c40ahihuwZTIOoc4MXc8hGpbqKjNT2CdHq9hvCUtNRiC/pSgLXmm
cPTQqaGIV7r31OV2rrzqVSYQ9J94ealCgymtEss1OwA2QckI3y7bjnT7QV8BB1uZis1CojGbp8IW
fcoNd8wgPGfH0tPGhL3ajFt0Ayv6LRnjbRlPEl1KJUoOsHhFp+J3scjhUD+wTPNbEpM+h1sJEQjL
UAwjHgozyd09P6YLZyWiBUhOflOnE3Ha9YdCYb58xeZjvvpiNRo2/4DfgRVtV7Gj85u0vE/w47uP
ZX8/jmY6c5nMN0dtkH+OSXv3v149wLf9j5/Aq6PohzadUfOqckCaV0pVLngUakVYX99UvLb+UUob
39pn/l1MqHRr3YqI76XI4TAEvQmd8TxVIJJoBNMEt3UFDxCb/UsY/6FtNufXu5oeCDfWGB7LmIqC
sYF3i0khYpNczTtb5f74Aac4iuu4yEmiRB6glU7n1iW0w5RmSZtomzheNJ56uutskPae8iSRZVFz
IapclJC55Tzk90REOr2xmXawNac9CT2ftBzJnin05kDYkn8njnXydEsIiLOWJf01J+hYeT2YnYwP
8kCHs9RjvDh2tajafuNAstHPKVSY+gMyRQiFtfzxMkj8KIzJLx3j473tFRrAA1IIx/e9ktADRmgh
HkNnGiHTnbxMrTVpDJAXYcy3givaOPp7CcY9ZQ7AOk3Ajjp4h1aFXoQPKqZ/Dx5IbcTmAh+36S+Q
w1f05JHLYOt5R4pysx1u5OWDnRWIqpL2owA4ueCOkLythm/i+DPTUSPEf4J31mSQkOT6e8pfas7e
Qf5HEDEH8CK9LvgFjcZTDAz3c27aYMWglO96ZpIufwT0A5A99BgTIZNwvaNLDbp1urE2fIw+qjTY
KAUmpANfDqFoIgUH5GOWuTwLVC/nSfncXu8YXso2VFIFqExuFOHCxe5SIU9C9D7ajiMFVvpFlqlF
Qzc9ToNRwGjCE15PV9ziMR0NZrBJ3ABgYySCU6EojBDQekvXBT/fKrU06TOPmlfgMk4l5g+Hh5Ot
Ft7bbi/n87qlLDdJ+hxjmRret95oDcSME3c0GPhBsRHjzos3a/ftKQTMNf7pHnZXNKkWuC4l6bsR
nNlSh8tDB0dB+c/swh4tk8lqlYJAMRPOFe8IEaQX4XzJiW0+NggqmNmBFRu6kUv7szLFCnfVkf4T
bxBlPzh/WqF07a/c74CZTIVvuE41GCo+eDOiPypx2jelW22I8CPg4caWu8r+teXDnSBRdLFXv8sP
Ja/ZuYLDzB7Nx5Wm1q9ps2WZUtw8ho/R7TWiQKH7FmbQoUivr0FY+mvQEn2Y8CBdqa0LW46KUbLE
F5B6NNulzNOjE8nwQ29sZcce+h3gs8fIV5v6ssO8E4aGS872QrR1N0OaaES8Mdg4BRHgJqQro3p9
LpOk2uJvkkQfyIekmhAVpbput1vXUxWi5j4BXFE7UgBcv56xH0pHB6kWcNC/hBLY5CxvJLpWBted
i9Bx+JzeCxcl8sS/0obaXpq7XrSTJkHrFNy0rfno+IQCz2e1BwnisPh+up84xi2VFD9fKbysDpw9
XNcdIkF0lpx9SZtZb9/5XdDYWIAH7hUSOi8EZ2tqgh1ICCfRRDAkpNN/dulx07G3rgWwY/otond7
Dz84RSdYX26GHSInsFcneFDPcmzLL9ZLcFnRNVeqspYEvY2sEVon13p8FE8dHfmpB4kHQnblCE6q
Nap1L27QHLOQgSKjY9m548vIn3d6PvToRpJH2kChcI3o2ztk+ZpLf9n41YA/voqtmik3g8R86FtU
L4whwja1R0TMRl3Z/F0hhhfikqBob7ckiiZEgVmNndNizooVdq68E3JdI3KGcN3N2iNUno9VxNiA
ctoV0PltzAKHE6YxjpJ/qbxRsCR58HixI4pBYel9LNTAJJ7txT6cGDVkrUTfCaj36shGG39ep6WI
q/GP5Do4BTf+5qUAdvhYMVkVSO8RKBt30evkqHWDK7eNfjE49eWnMs9LlAecSTAdvUOVusjz1SKJ
V1rvZTQgip9b8m1xUUhFTuk7rvs5Wq8fXqFmAANpUVBL7mXHJEVmEL+LxEWCRyHZNNXaEHlkaPlH
Ze7ig3zrTBvhgP90hjkwKe4nP26H/+Y2ddBcvpoZaJe9d0IrHpz1GYLifRAlIh+rYkZtkEWg6Jsx
0at4gaDk3ZUq1JHvn43sPppVPt2hx2Uyi/r7wLIPDZGY2NO5UX95hOKuryjh+MR/C+giS1jZKWSs
niqETOzOBo2yyoxqLvvcyWHpRqhogseBbKTJt8QmCYVuBsGMt+ymuqOfzCTbZ/wG7QwHYjy3byev
8wPVp35Eo6jiEbDuvr3bF50oYOiyEr5h9BsOzOziQKKuKe5bsp6cmVPD4zg286vCt+pjhqDRJndA
vG600LH4eabyVVIjqkn0BivueG61pOBinOFaguOgp6d1la5zzYZsO4s/7Tc8rkAz0+ldxYvzW5YM
mKKih7wu7Y7+In1Ej9oZ3f7VikEq9SzX6sBAYmLYonxov2goqD3pHlsm7auLXrQsQCIr6Qnj7vIt
PhtoAlvUhL2wL5/BifxcqMDTOkmnGL261ZxKfHAe8Q8e5Q/MZbbmD17cvNteuh/noB9EN+bZwRRs
MtzA4W1LofQKEdQMvGmaPAWd3QI6qq1+8RjZtAk52z/d3k/pvecxIjQ/P6xZeqTsBaw0x9xgB2HH
vKTxgJikAdlYu2FnT+4gsaIN1mL/VgrSshyyECBG+ALQCWIJAOR8i7wtUkKW+quMZT0MQo3bzmGj
U0yl2Prm7rVPkFRCFUuzCWdwfDXQzjpm5LACKRYBsyajDxw0kQ+a+mqmmmpkSewSakMEmgPPrDP5
ClOQBAIk/juu2WHX81KIzwvfs9CvoC9myN4LgOyPkMv1KTaEQl5xNeP0Jj9EBK9Qls5mr3/DKwXT
AEeYubrZfEh4BqFMxsBqQ3oBR+j1iL1Nxr9XWIm7PRgOBIymXLi2wHhMPJy2BDHaItmPlQirVAxR
ZbEVKoxnrz4YIunFY7VmK0VWNzs=
`protect end_protected

