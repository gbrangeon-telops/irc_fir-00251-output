

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
esuuckrrKLBFMMgSrVud2ZnB0pvEqrOMx6GkXz4dnPp4yshTD6+Y2glVVVlxat4oj6oLNAI0JrQK
DY/z82hivg==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
d/1Syr0Yfz0kK4aSXCIN7lq+kUu10RASco8trwm0ImfJURxtGkX5KSPC9Owus8m9ZNLVa+4W1mNi
DPA1z5v28araMT+WQkx+2smTTBb95QnM1r7IY8WLJwhz/4br130YtPfh6ALhwuPZLGS7lh5+ZNqa
WUkp+2aPy+o7nP5Neek=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
EghETPBi398ucn66loN/344Jtlwrx7OhFAMdZLO3Gvsf81gd+y/lO92JbZIwpE5sZICUxsNH54dw
q7y/XtZVcW81UXDzCet7Fnd81N7WGIqo0pJecDfSTWB8jEEqdLB/p9QS5cVBozkWw9ZXd157NWH2
fYI6wtb4DiMK+3xbswRz9tjt4QpCCW6pl02xp3h0AjoDyHQfQiHlsbTSjlklPmKa/t4Bvl+J2OsC
lbC5D/MuvEAoTUQ7SK30lNJDTITWXb0RGcdN8tf/1AbxeMFGNs+DvhkJcoBe11Q4yCS9vXGZYmJD
ooCuGIJ149GuhA9Ebc3S+zqtQIqgB+Ip/rSAVg==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
XB7G1kS71wIOs+JCFd2Cvu1TIPgCW+AVgVRokt3aIVEjyzOaNQpUv0JxfFRbYs7j+wNszYGSy/VO
ucUpEKb3V/Eh6Je+1SiQK8VPkEGyi6kMKodRtbbO1t51Edv2l3Df96scmfDCuwUmCLxAYCnMI34o
GJA4Te4oMZLzNzksU0M=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
mYbz74Wd6t4yNkXqEEqIyqTMYr1gDkxJuJW5Rg5GXWUomZKn1t4qMArQDnPwJx4y9XZOu6/MtCnL
fPfEaeJGNkk3xubUfcA48NrBjUlfoqpqaC5sVaDR10h1kTeB38B7pV1iwRz53qngpcQ/++tRqM1Q
t9nxWednDhGT13iznArEKq20RLCcpL20e+RRoIbTe3wwmYnDWI+ysKyhOx1k2FPgh9jb+4RZZgn7
7PDivXP/gbNxEf8PXBmODTX7OG6mMJYh9DN9gjuP32wcsw58ZKTKhK7ryO26lHYq65/5CZ6bVTRf
+77RaLVhpZ+Bo23bR+0rH2ulVAt4vAhPt51hRA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 26704)
`protect data_block
buun1/o11KhRnBZIcKEKdBnN4fVacx+wnurF971GnTp6yaufkhe9tintDbWkF8QFkvowVqDiFQbe
It6LMTGOcF2H5WRAjn13/RRSVpvZutdYAw3udshvnlrEfFMvu3o0g0qxRPX9guOs7Q5r5XBSXQd2
cKOYyCWoz1aECyR+9Bg8drH6tZxX2S+wmccqQr/5BRMY8clR6P/DpVDb60zEZYxESLfRJ1xVOtDV
CfiikbXwewUQrO/GFNGBkRcBcvvv0hn5K0bgbTo9cjri/yxp7gbJoSfIoLxvvmFjJxlU4ynq4HHN
nC2W1gsEKy4WlPRhPzas0GrZ2g7NL7gVQTKi91XAaz+1gZ3F7wNsFzVYSiBrFJJmpxeRqGGLt9dK
hFUAlHDWdUtWrhjlh7CeDSYXJVlewqzgzxTrPU9jvEv+T0OR3r1yRYHY9pzCc7cZTp/v5r0Zl8+4
W5F/oQwMwoBLoV6+/xapGaJ4T+5byiYod8myiSFn7/oCBGApXtuKFfTXdwCocTb5mMC1zRlnfQzb
kiP9H+mHrrJxotvdYzIQI5KWvLo5u/8IE12bXnSD20bNhwlK3nWfA2ggNCGvcmJIfZz/KfgMNsjD
xbWrtJ25of21iLYRI+LCAfQxqcab9JlUVsd4BklcIEO4yRq3AYZhzb22nAjYr4RdG3o+lmTkfDRy
XW/cDIDL+Zco8mUSOuJBX2xKiBZYiAHcvVF9SllvrFzkoD2/TEZBSMCTVAAdJAEUNcPJ4Id48dxt
iKXZ1eu9A7xlG1/ZWNUPVH/BSFpcnkhs3c58tcfyE/76Ru9gp7huwqpdNpi69gEFje4zqP+2kcLf
7jzikyw/WFgIS11zq3B2Tkr99nBIH0Cr1dxqM6G8ASzb8vzffQV0sQiA0enZ83D638YLhOf9S/CE
FqFLdT3P9EuuVL6OscC56ytxcUiiU5hvH6AvB0E1C8iqDeiJJQAGPpD/rQcKdymIbsu2npbn/hTn
Tg0O8jGKRQk2Yim/fwPyHie1jKpppxZ+Uc3GC4/wcVLNFrfWxphE1R3ppVgPyWJYeK1lVZ9DKv+p
ZkU1qVHIAGfXCYV0lwOR5FNY99NdA+u5W/XspgYFBrKV9UWCTLqj30Alg3RfwALHelpspAD0o07k
mVjsThCcCW/DIw0PBIBG7CEYwUvOjAJK7S4WcSgbowd5o4ROx7tZK6fM92aEOCC5xtP3Hk2qZ8ji
vnDXpY1YlJ/bSlNRxLRX/L+Nb0xCjlykOO2IJWmhGnYR+/BwjpqIpVqccbD+YTXJ0CC0PHHTQldY
Z55fM+iged0Jp/BZ11RIdIFMKYxTuO9diDrrWh2bfdXhTvamG7/dcupbS4GPKav+jd6dbg8RXGg9
oIJtaKUns+YFbmqN06X/5l1fnVg3iGs8Nr51pyALAASCHj/z6PzS1jD99YoYz2rFoniOMbVs7hZK
4vmfUSB72FBMQtWjj4FRdf19oAfXZF+P2bplyLwjZpYf6Uy+2WwImV6vNVkmZdfhNYPxXFbRGX+J
2SVOb9hEtTE1Tt3nWWQYp70zjYsaAwgybGdC0z8llK9wmaa/mSyXBmeLtBbOXWoVAgyO+C3qYlY0
cqh6OE5UQ7yEC7zBimw+4SbEUt1QrFz8Ysf0GzeZwYi5XXiiKrBPHXsmSkvXN6woXPAK0WJPQ5pb
tjGeII40xd3TSb2IWaJfi8Hy+fwWITViETG8tC4wuQSP6/HL/9oKSl5Hp71SopbhmgVrSRk0eSl+
Kbzsw1rewoCfXEYCa/I/P/qbQfhIVYsBfCLKw2SkSgxVCPyr2/ucaZD/yGw66FInRd9WfenDwJh5
BSwnGQ4yi+aThCzJNRFNv6yCS2Bhkw95UMG3YivXapvpF+eZGuab44svlO88el24hja8LeSN7jaQ
S7f/AYbxXZuCNT8RJVGC+vyoaAeIl3rswNzZyKY+sRm+qMZEi7kMXETDzNaco4MbX1nwuWNWIm6x
2WlULbs0G8x2fPjYUBLITFntj3Wojsb2FrBybxB4gWwd9/OX3dxQh6jl/+VYOzm1ftftPzd4DlRA
6m2n/Wsb6Q8cYWEhiAcVGSHT7PFhTuXfyDve806xrPNc9IRbIx/d/xgcivfdMwsrD6hX0JUm7dPS
O1073oLflMsfb+Fh/X/oJwGnIZsvVNRBvPgL2e1JERtuV+44VzgsiQNFFAtIK1Tma6tTswJcmVZ+
HO6/H1MzD213tLk3esqfZW3l94CHwkp53WV9kOsoSwakz69u/0H1CXaBLrTpAQyVFLOk4muo6UT+
kwkcMLECkFEXA8/QfaEE/s3Oz283h8SLKMgQJ6OWorknHa6sg/77ZDsOeQZJ4L+s/ueY7tvVSiVW
g6vLbghCz8wUsXFs0AE59wB9eCcflPAgJyi9Gme6rp65tZl0EKTsArpG+76BPw+yKFINNsHW2iaf
S3Dv7zxqt8XsW+BNElAV5gzo+K/ndKOpra+gncr+AZWeYtX1h8M7Cx0NaKHZWnifp4q7LG2yadZz
u0Kqx1HcBken0ZedAUbnDu1fDyB87Q1gM5Vu5WHvqC/3Ywj16c1m3U8glNvJHIYteHsp0BJohqjt
IAdCEAwYabwLnUUJf4ADipCSXHWYrA+GarDqNckwfvYNXrzx9Cv191gfsc2hQaEOb1rODJhTD+It
SQKuVis4X1L8dFSgelrBxKqTa8oGwpZPVqk9G/n+E0iJqggstV8PqpDty7p57VYT3Uj7JIUPIFHu
F+ZxNvL+8/eoKTnE7JP84YUD90cUNhWLcbKitSZ4SIedfnuy3z55V0WDLPu4r4vNK6HoZMOKVAFi
LoEYBAajH3btInOeW9uLfmtGl23xzGi+IosBtvb8mV2dej9Fy7jF3O8m+lR7NNwymmKFLHvpmDZV
6K525JbOPwimXc/RyIogzv8njqMtEaAYhnvrdvfIgh19zwuKT5d2B54syxZVE1+kXM5WhltWkK37
I0L7bRSyiLIzuIE8+ta+MxqCW2nuMkHYki1SDuazmHLE4OWagiG6BaAiT2rRSg6NVIYCq/JTSE1Y
9II5qWf6zpouWF6DZG3SBkNfGCkbnpaFBLtc2xZh/BlLbwtYbT8qP8jvs/AA7aXn1hJj8sb3STIt
jjvNZ8cHhI1+TwQlp9D3JVEyiI6qu9HEhkr0PV32/P2ifwzJjjdMUGvmRdQqtKI3eciAQxkWH0pw
4/6n2NYUWvdhrlATAuvgrp+56ncgUPh1/5y70c9mHosNypPpeGcL7SMF72BcmTXrLr4qRZRNEEid
UhQEJPAloq5vyvH9JZ3y36dbXHFyo8E3yiLAuH7FfppbnfI0/SJWjjwQTxfCsoQerEX9zt+kxNte
aMKpBP/Rqi03jR2x+bNDJkAqdYFVhMkevQsQUPnAEqFFRuNiA6Qf679MpyqZBO8gGpPF+q9ghZ1/
/py2fKxJW+k+2CTNAosMnfM6eyoPbmezu8ny2N3vZIlPzkGp5oydSDIO4X0FmlLGV15+gKW8Mz//
xC2LT6rV83tJTZAbmdTz/YEs8+FM7S/U7IbAJxjoXB5/M6JupZZVsjJrByu0KskK7U9k2RIw0UQB
euy9pY8CJ4Th7FOV4RbfInAwrvYR53h9U0j3hQ8x9NEL4iXXD6ri05jBeKcPZqzmnoc6mBohsqIp
jFGQZkF911cDPWJ4HLuZcT2FwtvwuqGoYz4d/00HDn66LCL4n7P1Gnub5L9Cu84xaOdonBltEmQg
FR7CmRnI7+P9gqOH5pEG7whxda6Y7uzTSNof1/g/EAcZH8CyVuQ41xNyIC82VgTHdlPmBRdN0Z0F
NDW62NqqiYO4UhAGjrYtgF9hbLTs6QbTsLlc/GMCVkqY2fGgNbCqidKMbfjLZ6xHBdZajSueM9Xu
RJfWQHALpFv4WoJuzxFL70osCXJ068mwzZgYfDJoFs+QurqYHqfPkLsajJ1KvWlZRs068RpGGZqR
HymUW4ZYVfhmOeXiSZQ36Yx6F68T6UT7pkqubfH0ylNgFwCO0doN/+4tdqVBSVJPb7qqH0eSSbov
Saba6eNS/bt+470IvThLy1Z2A2pqa67xLdE2SiB2ScPvQb0sfU9QLHYiUjwV7Vi6+ju4jXDzbT+h
CNPU0Dd9wVPLUtz6PZrOJZNtnoSj5rcIITzhnArRAvHJihlYCSji+x4OQOz5JMvLRMuqObIN3Wgb
02MUqI4tOtaxq911aSyIBUIlgQ6+fpXw7IHiEsaERz0O8TgXlKJY7WD/yg/Nr2cBSSijKRnzszoF
YIFhpUlMZ0JUVyPqPBg5SQIpopytFQkZMOM6+noWJKrIuA3q3jhTOC1oe3On4hYhHHuGnkboYHtP
L9tkxt5Vly60CmhXAOMVrJngBv/chdMA/TPevPauqAWOXW4yHDLG9w0y5hqwevzMnkmqvo3z4/Ic
hTw1xObK00NFjzZYrJbRiQeiewdei8YMbZPQfGYTKcRtNTp+MKSi2JbFY4YX1/Fwu/NldyxEJnUs
fXbOoB1PtIaiwdVISoFfITvaeXAjjODZW+m+jMj64tc4PMcmUcs/+w8+3jXEjUU6pFrXjdtWKy9N
GdLH4LMsv1VI4b5ilfU/ulaN7NzxEVieDc/2e9WHiE9UZNoBO6Ew8vFnObZTDXTDyzk+BWz+WVBE
mHqWEjEEAVnytjBy0jC/jbdeJWzPTM/P3YHIAd1C0QDMvzjKPk76CddYc8IaPivKWC4INTz1F48O
ggQHQxKVBpnSfgCtalzumLttpvOArF8KGt2gtyo3H7K4W6EQPzbkJA2Po73ow2cvPbnOt0MDMUcW
2i5lfLkeMNGg3c99Q8r9gu4ad3/M3g7/kGEIAU/P4otwi78QGAUfcABfPzGHZHJPVsOJuTDxXsn8
uGxV2oXJBiuGeXjitnfdn3uKX6+pkxdx/1PP10nVKXVSI3wzRN0saT/dGlpXXyhL98Jp0EOj0IaH
tKZmXOnXlfAU49ywb39IJrQlLWwGD+qfWyiOeYKhmzGM4ddh/C2SHLGj0A/QcQ9pzMC7hsNc8LG4
3dMV7VEF3UDGQJ0D4YnYGCnJSZdDONueMFDi+2Xm7qLqjrMt7m6G+gUrQeS2s7DKfMVH7r4qRamw
fm5Fd5wu618fEhhVBQd+Qh0iPbZNfUQQtXXoE3GhBtZ9AEvv30JG73n7dM0fRd4yukjhA6PNhp41
mkVCCIAs2fAsW0EsazPq1T71C4Y8t852xfKVFHSk85PEQk7a+Gaoz/+H8kCjpZCrEe8F1002Z3je
fgzricpPWzQE3nsOMnh6ZCA1QWphj5Yj5Yw2kyTdCtMJJChuUFb+aI7in+Z0iM+QP4sTvhqCTlrM
6542v042g/TfHc88azuOTgxiZqVr2jt4LW0lbRI3hXUWBc+QF14u55S1sSji9uq/T05TVlqX9gaX
ZFcivu4kdKH8KJIcGByDP32iPUvYiGYj+QMkm27UkFrGHZrPcJPntnLK4RyXBKDNQLZuVDC3fMJH
snJjhPlGZYFhaW/uvsnGBLrTjTo32F79KhW/f5LAMiMG3wMUj4UEIveH7NNnNsdtTg6FPkYGxkFI
5mmhiVFQ53YILCNSm84mnHc0nqhwL8jFnKcHZmDD8N034abwGYf+xkWp1XVg+affKYXy1aOgQa2Z
gRrb1a1Gru1EegGJrLLwD/NM+uNOtlL5p54qePBWtpOX6/ybo/D6xSEf9OzpFLFaIRsNXWNgca7U
LRqcS2RTuFumWukhMmfH/QmIn3MMeSq+JzNMHKrGYDsVjjGlp+osHV7jCUCLRqHbAW5EybBOQqNJ
9meMuGlezepv0dtn50kuALhGBgtgo+NDxgV88+EEF3rgHIeMd6FDJP3n4YAKn/Y3a9ZA8fIvuOek
cXH0DWqRXTnnw0LIM8+DybOsAmMPyfQWpvsQdLJ/oALJN6TTseN/w2swQKeEkhQrTXoISYi4fRQw
fmEs/larLg7bv8aqblJbmO+ehdJkaftGMCqDFcKSiBh0GkTiiDKfHIQAKvfLzrTyCaFHi7RusgAF
qimJfOUdkBfIp7E12xSbvKKedkkGX6QSTidvY5rZEXT7uGXBH4ml4eLfCy95KREodpxM2lq494A/
T6HQ9R2dOvgB6QoUDhe9OHeQsYjU6YUavW25GBDOSmsEub+uTdDL5jUWLD/OUuBwG9JHaAOxI23V
A9q318RZS5eI7ZgrsOZ4W78lTWUh0GimnVfzzT25Cb+8tjtNNTeTLbbjhfqnEOoa9TDUj7YFxOXy
tYIiyfLATpDHlGjJT6H5H7Rk9eSzp34sLhjLbcG2POVOr5ELq+Sex7hPbaCkXq4T50HDJFJNIKrd
Fh/2fxu51EvV3gP/b2qIEWfF+Slw3Ga9WloGRe37ZVecc93mroGfIzBl7IqefJW/h36p4lQPemwe
PqE+gKeEFr1nSWb6bP1k+hm+rCEPHw/iljuv8VAd3Bag20n7cz3bipO/ui0jIqgEL9iFyIEi8A26
m0z9Vsipi9fzTz6YNrjowvxziD/zLDw2r7/PhBMhorxdGojx5loijij4DvmkJddVSKT9aaAmCVKP
O7LFj27IwqVVbyTn6fi1h9fmbGItiZhNN8MAC+J/SnaZaB4r3oXRff3QJyruLJorv5loq5FpihsI
vr9aIH1YrUg2VkkVwlG6Lw71pJrFC7U6/LTZOsmPowToclse5oldH9DUpWUtrTLxi8IN11uiu00J
cBdj+1FQirWij9Wg/qS9QK/7GCbjNTtZGOIQhR+wu1KjSQ5Ruwn6s+Lat4CFOgxFCgBesAMQQNWd
AArN0JG9+z9rUzoQtryXKbfE4P9iGwRBrSTvXSFxoMRQd80YkjLerIf8FGnwMEwpYuJHgI7hzZ2S
fmRNR74+mGtlORn6VkwPuS5PxF56/ZniW6HpZi1uiRcOh7OTdjemPlN5yAC7JuyESoy6+svicnjp
rg5sIWg7HUhufUJNvQc6jGbVONt33FEIHPp9aVFE0/4PQoUr1vq5duPaOfK4yndYXoCzOnHgJRDV
qE93W92gDlk5yOegAmp5iujWbuIzWjiCm9eINkWSoHtbEdjvQ4f29akQc4ZUi4Igdmh2Y0In4+mC
yNNblMAhbVDyIjIYiedWgX+qf8McU9Pk51FAnVtGt7MQGsK1gO7PNbXr1DgY0Xy81aNPnDWfHJKw
dL8TazJeFVOgEvdi4oh5rJWk5JE+0mJdIUXiM/+HjnmjUqPR9AjgnBvyTj0NmtB7AgRoTekTfXdg
ct7VuUWKeF91Qj0JoSViAXEXIUEEvzEeUNLXPqPX2EsZrzQC4ZFTsIZEd9f3zPWdBa6T8j20dUri
X3lzmTCXJNfXfAyfF69kffwmMB3S2tQQVI9zS+ze4Ta1+CkWWpcrpr0r7vuaFGnfRHZMhQsVXPjB
lZgbpAo0hoKkEmpEA3O0TPp6vwyGlSz97aHA0fbA7juDeGSBjkNcbyOuNWVG3pgHuWkDLV3e8qkc
m/ijN4KP0nUEa/Vkc/pwGZq6AwKV6NkR9JEjBhkJWdlnzL4Z5WBQtrsw+V0nck8tBizzWzxZNghH
GVTL9t8g0i0Ek7r4kzWN5mFAUf//ak/TWs3+C9fPM+zF7Oypz+jBWrQ2GIclaZRJujhlPf4jTCTG
VZBBukO8oHh6hNngVQhe3YUmCSJksLKYTmBOeCyLnbVS5iKRhKq3j3OEtBy0egHDO+NX60D62Eo2
RQVEUmhNJ90Mys6PxjSKebV/HkcwPOnlX5lm3bAfP5jsZMppCn3/IMilTV5JWHdBjWUAx0XJoXUz
FiwJH/oz7ocD0BW6/iZau5O+/yaP+9ZH30oBDXDEbcH6WC69gjxbN9gLzkZQUTt8lX1xx4bwa/HR
jmqdRAN+B7UOOS35f8la/48Khvlm7dnen7PWPqQYV7MiyzlbQsUaKDIpwfK5mNN7eoVROs1v3+G2
hYCF3/vcMipEJvs55MBwQjEMuju0VRfFCDWnBI4FteSwHAn3W3uHKK47jEY7PKPkgeXQrTL2/uK1
vKj4RqlRn+KNtEnGgaXii7BQWAGcO6jxsXCUivvjCdyqicCmyGDB9T9kaXeDhdV8lsNZ2DNkzm5k
0W7DE3PSSbW+AEdeqnr0xqucWMqlCWbj9dIFMW45G8mX2Iy1sOn3FV7Htz+di457cFLynLtNSFtg
/9aLd1bqssEsqS3MbJfubvXdueNa1MuaFX5n9yiXleoL01MM99e/rN0BVpGUFwkXpCJEFg5zp5RE
i4JvrCuhVsroPowEiLKFX6r7TKp7cMHje0hQU9kxgxQuLPJgXxQiF0UqCkCu//WQlbvbBFfnd226
kd0wWoDxbYcWAUxcy19ys8wfibzbbL35ymfhAVEm0upNssnrGyEEUroWMVYDQ/iCvTCQXmzEj6Tj
3cCAC17Z/GKC6Si+8AUC7RMUg6150NMwfmQ5jbP7G+igvIq6IvHOo9jR/CwW43dTb4QtdEqUBjRD
ARdtIE0GOv2dIfafHi9JeBEl/V7hdP/VEL+fN0tYEPHGdAUSMBXg2z3rzmMHh+RSP4ikpD16Muwq
Y+uGvHr+J0dAPJa8S7uwmZWv5q1DAVnd/PfWKu/ZwiSfqy7ohemNKyT2PsN5rdC4Bbt0NUttHhda
Zwh92qKiFgX2LLQs9XpDSF7jJ4kJGRg8P5BeV3Zgd5/xXBH22n69k87keH5Ex3txiPQ1lOFf0tTW
qqdWUacFSrGo+PVTdwktzRYRfv9nEDpgfgLsWAL5kwVz1pU/xR/oCMob8p6Jp4e2VhYA0Pks9kUq
fzDmktnhrbt495uNyfZCrUG13CF+jRLdTi43Ij9rRKR099bZGEZ+UGm3bZtDupIXjdq43I6sTHtC
O5VRgMcCAfiBAeMqd1At7MSaX+4uOYr+blQUxp/C+vd/3z89SSPUmgNJgMBDGxD43IB00K9Tu4jF
REemIs9FRdgtqtO23EvGLFSNAi0f575vTzMy+tfXWbUlnseaITpm/H5lULqN/pVbLt6Dr5lVgN4d
1yzaObjWWv6f9Jb6PldouJnIQX/9NYRW1RiugJuc7qg67g29R5lqZ7AG/gUYDKgbgT/5sZMj7C7u
jqzX9B6Ah+ISfoYZUTy+nVWrZ+XeXpPXEBiFAfz3YwxRjW1Uvfai1rWxNExzWlnApdl7qvMTHq46
puxTzw8LmWnWWvq4wZy0EVk3b2bbTaRIXq9Z1hV51NhruKW3NKekeFweLoxme6fABqATnckYnIux
C3vVyqPcsGSpCvV1d3+LbFCiJz1uuEyADV8P6W7kern/ZfWisAeeuE37EcGzxFhXJIf59v7CKtr+
xcVUfPnXveWgf6BlrXSldZihRPIHWbYK4l6OC4QYxbyLz0f/6aXEQSKzeNz3znheBFIyW4LPGnJ7
vr6xamAfjQ/Y4Q/AeevtJXqsteH4ig+oeJW6a7VopGZcdRfAxBy5CMWRF/PJEu1Ugc2jlb9C5UQ3
+3V1BNmwju9DS2V6Bau7j2xl3mP6oPKBvojyq3b62nt6DApmJK6jVLQN/YhF1pfVgwJszSJfPKLj
AaKG9vGFuZptcMMn7DOax2zZ/CgywTiMa3nNw1DIbsUb6GhNQcHaf8ljf1A7mMZz6NcF/yJXWdkz
me5eFXdvXQTYd1znZXebYJvuLpP7aYqMZMWfaY/+6iETlRSWOTYn1HlPsX15ITs3DfwlIq90/6Mi
ZvHa6H1UN6WKZo6FwEECAxe+WqzQ6vswAS86xqQxIdqM7gT4dHM7eJIRgX7+KdLC/IWfgj44HPyT
PHXtDcgLQTCQvG1gdKXsHbAu7xOMcuWuaT/FOfTTm3u2pvXk7os1qMXlEdOfuIjnfV5MrT018vAM
RjfriH0VCe6bg8P1Z8vJ55cCnFW5tfUT8MgzU2K0hs5hEvEbqr1fO6lez6162WKjtnJSgV2dXu0f
w89BLkOAoSBOz0MHXAfJAV2QLCGQOz/LGB1AEpR3JPLki6Hb1xtmVhfY+6qH28n3Y1PjTgiwIib8
cqQMKT7oO37Gx7GoblTj/Ys6yTXBR865BNB44ZP791/Nx3VZ3uqQ1LqIneR1uw19nzPSOK7kuUvp
oE706/enZWDPUjBRNZUdl4TcP/QzyKuNbk4el1nZA4WwzAabr016ytdhRbBX5eoROsB5We3erOLM
6xQqkOySelzpsxpbvkSKfKHHNnDP/Dx0wCILMLxSfZMlVdcF6KAwq25AlIaxJKRDb8m/KuUd6KCw
F5yMeyUKnUgcnChT22FNuybm+ZlJmVtVMC+hqaauLqn60i+uHqZkdsVTaZXU+E6NbYPA1P58YA30
jsrsXhNla6sVgH5pmDCdYneEgfyuyJUJ31TKMMt2ESWR735+/eY3tUOPBWDY91KsVtBb30Vyy901
zjQfRM3o8PbqtydXwJmt967sfYgI9BTl2Z8nIYAuZvg8u/tsLjqKW95XmVU5zY4ORuAcH9fZdxkW
ahX2hdeE0QtaL8N25+aUKaojdukzpdPHkc2F5sIETLGfjfDoWYJfGrGzlh9KpopSW/AVN5MCf55w
GG4h/2+PsYxejbh0uiosDWmDewNbqG7bsGtDOGnYP2HYMr1kQ+DssFDG5LfKg7QxYso60me8phxG
eg4CVU7hRbp0XmQkiFumULIQbHXFiDFDt09fhegiIOnzYJvNWPXUc2YO4uYjgoCaaaStGIjpIRXn
RKuYiQ0iYO4ZqMJRSV8Yvwc4NUzoetavyP6SI+xcv/B9qdVriN/EQNI4aVrd+E7golo+eQq4aBIU
YkzV/0Xu8rQMWhaGJA2t8cgH/97wi2zAyGbjIVtqRFs7vfZ7m1A3Yn5WDPmbiZbPaOwvT+ZyY+eY
/OA7QjbtPknA7VygD6eO458WN7CLCJUg0e5vDTd2XpvnLB9M3mXLkoye4CGMDtZPsDiyjfeNAEbp
U22FqCsmcDTvk+hgMbOe9Y7Q7morlGVSxBXyCqlE3ictzeaBFL55htkY6qMniMWwZKgdjNOIknlm
nI2E+gNaYgVGSyQpDmbs6FKGLnz2Xvh3Z8xEREWItEks4Phjn3eWczSLItpB+j72GF/P4BKzx1qD
G9E2EEw8XFfboFFRIPnALZO6xNTVr8UCKoxqPisarkWyqHEbVJCjb4Yb04DJMM6Cr89X+AwPX06P
52zoPp/jdlS4DWJ6tufH3+GITR46iTGT8bUSDZutrJSh7WuyEh3BW3YGZQcs3OmF3yV6vsBo/aas
/zP8wWJQJJmDP5EePFmRDln2bLkalKGI30+pjwgsnnY6mdpLONFYk3NQvSmRWdd7p53lnVeEVJPJ
apL4jbYPSZSQtp/WyVp1COKV/TzrfZ1pPBWIWC367CYsCT+J6Ng3udeJCWfnyWY7Q+EEZY5BDK7S
kL46eqTth9rjiCtt2t4WPiGdHQgdehIW8+MNQAIWEvrmJYHNGwxDmFuuJbyn71Vjsx3WplTS9wpz
j0vTrG/wKdW2R9YoBxRvhFXwdMykDbtQSFhauTp8KsGKimo66RrhkDbUCBKFaNDdNmH4g00g8oAx
2aEV1qUTm3Rv0xErzq4G8jOprJgesFZ+3oaqgvvFjaHev4QDIrAk1597AIjRNTn2Q6YNb3QRelbA
/R4WD6vOHObwJILED3fkKHR2H+c2k+uPLVjRayKElwdeub+LWi600YKPRPi7ZGy/q0bcfmn4dvyC
9tbvsJ/l2uYj1OLhUlpixnJMAGAvO2cGgKNjT5a6FQbTidQh2vURER/TRafQy2EXJwD9+ck8jAWZ
BwjAVn8TH5O4m4eP62OSirxHdL/AfPeteTvJxXXUcJKAysbr+9tVvU5R10W8EM9RpuiE+kbMNmkE
biMxg+rimwHZvfDeilVWBCyOcvG2KJVtfG1HTVdRXUM2EDFZSEsVMyrO9kx6vw5eQPysEhsGKhUf
Tx5E6SXHGF84e7Mb7xpyqRHgwwTCmqj6xV5B8uAlc8F58XmnFLv35yMA9JjVG+s91qvlGWujCIkF
AbwOrB1v4iTWmdgh9CDgQNpL29zSepUDit2TcezJZgWbjVSkNRPixf5wTHMDOnHL9iRZTltpntn3
T65psSUxLw6DcAH5JbjHT28VjvhrB2ZXVa8Z4/+2+UxHepZe/FHKWX8/3feQBoK0xrcju2pDa7xh
Z+OJBryNg5efRJDUCw8Zu2q5GypW75jLcjWuDwOwX+cMS9pJ5bDOPm0dnPbgOf5e2Pftddotx5rI
IQnXP6qWLI0eB6Kbx01CPJmU5OszC9g9U9emEA0ZhmbO4U6aZ5APnmxNSSHdt63W6pZurgnVBQi5
S4rfJpr0pyhPMsTzSnBZSiNjRo67zv9qEHV+5WsWagcAXR1AOAMt1TqRTQsBqV0qPNPm9brvkmCa
1NF2Ynen87IYOzn1cJQF9VIoXndFiMhJ0feEUcBRllPqmOMNYRSR5kHxxbjrGUyAGKaS9czXwhMj
2iyQZF8t4AB42PPL9jaZYNJNilNjd+czj9cbkjATe9JZTDk+DG7H+Yr4Fpj43/kfU0J29/vflokD
IFDbHT6f95f8+4KIt2bhkcw0HAu5mMjRZ/UVJNaI3JSN6lmiHguTOZe8yIHJmF3ZYHxMY8IX1hwf
prK84Ny0p2lAH25Gv8TDqO4FmIZRGshxab6DoEubYrzsRhZwgiyb+kh13ONZ167glz+XKzFPWDs3
14f39vCyaXbxpefFN6YiCXZsYZPsLOrecByxSlBcZiLIzaq+J2lZxJS+jJlxcXQ3SozgCvDDAWrg
aWdST2sBv7Vlz11lcoucCw2ecvmq9Mne5Ng9YxoC9+uG3PiJ3aGrezpezBd+veOHNfJT6iVTrEgH
v8xCozrNYerdA9PIUvWs3fkBXL6oaTNqIkpunR7bnZ9/zNFt3OI612FnHIig3mxHTwKEn2sIZNVZ
1cmLr/Lu2I0Mhv4mh46O+0CP/s9aMLJtZJKKJrtkSAAOOdwsgCcFhmhfL+1WzfyKOL+Yb/v/6RMj
WwU6RZJPwrlj46Tqxp2KorKsAwbuue2OVaGb9GKXUgo0tW6OkTzYtbt7hxbhKB72iFR+DdcecEGC
G6GSmtqHKzi4+392gv853PaoZHfUGNQRaqsaEQOkXbL6OrLrfggnrDOfWeOQHqt2cNG0DPI2AWQy
X0oREDWxcMj22ycshg7IKhpzTjg6MDdNdwg6i3SAePF2PLA2NLXbPHtfXmOuf54vFBZ2w7LObklk
leXQMjh6hD82qUKB1C7ieh+f6vTS11j2Lub6flLHB8d078nCBnhXedSVc/9OpjLXpk7yw9hpaLiR
MLnSMPeUQ8nLQiRJVubTKZyzBUVsE41n/jsW/fpHQoh44dRDPOx6d/SMWcCOfKRQxLT4k6naVMEp
Rb1wawPpT9hH6BcjHtBuc+pRgau+mXT+LrXq6qMq16XuSNHuWAAVijmLfs6QrLeJn2BsUCrlYFms
EJBH3oJhNW+gcBfWnTZ57TtLTpfloKS8uY1h6OZPY3uEsNBGErmY4xqvxoKjziY46NTve4v+Y0wh
xuWX5tJqF9ehnBcrviOF2lSsKoT7DHOl6Jhzgg+qyORbhNjoAIr9qWZn6vJMk4YI5nGmMFAHsyhh
ZphR6V2FAksa/KNQM6MSHu/wTy4bmcsUDBtsKGWxv7csz+gSEX4adCE4f3wQS2KTwmoqmEk6MTBL
N884TQu9KrMs4Lkg0QJaQ/e+w7bh4Kx6S4ulLoeCXyPICJPr2R5sfYE6eIDVVJUi7IReBnCHifXT
5J8z8RLFuJaFSu5KWA+BEgXtuZSEeE9RpAFwkJdFT3GyFBVnzfZxikncswNr6j9sxziImQszYvgi
J5nsLuo/1w6KA8SrDCFBreWfr/WRx38LWjSxFszl0pSvoxa0Q/CyoHbKwVQIrDSyI2EZRFHZsm+I
uHddYeWUKdxAdb/zRqDoX3wWUMrR3SXnbaW1A4EQzQl0PqpY0Q5JeBWH+kTD98BzJa1TSSdEEpwa
2rP/1kglPYdDOh80MIIttujacwBvcpsWwuecmj27ocHZfhVTQHBowulQ++DoAnEH3JpvWyCK2R5P
RtWKuBnItSniyk/BAogFAeyre8XeKx8rtYte3jceL0wEvtJ+FwO4zm168wq3NSlzyzyzbUVCmzUk
MMN6PJZW7lCJYIsYmgkxiluvcW7cVVP6s5KLW4P/IxxcRUdAdQUleDf5/Y941cQ6bjTBuuDbDaLB
llph8cCEGDphFRcRn/WGs8lyQauJzd5rQN0vsxtJ5qM3Dnc5zoDCjEDCM1UWV9gR3wGde39tJkYb
JiXV2EbzASnseOnTpNKIGilx9kKsHqPMPlyi0UcoaB0uZmckPICeg9bL9gShuk7+N/HimsklxIwq
4ehleTt9vZUKamywCwzJPTprFQsPeHryOh4rstJeJ4tA6i1Di0Hic7ASRh6q6nEFqyF7k5R3nBS4
8HYr70bZT4zkfivymfZ4Jo2W9s60aXgqeIWnqQZDK5YowheR6GYbVCwaJcRQP+bnCxPGMT+xFf4t
UAkqx6yKs2ZcfKme5nViJ1/xeDYS+SC+Amqc0ZCTu6hiPlKoWtCIiTPbfrdNfz+uwuCaT6831rnM
FOjDYqP4C3W7dpf61aDmVfSeLeW9hwQmKgehb5f1lPE5ADWEsBCtctBabt0qmD+LGzeXXlzUQlcL
Bvf9hMyL/2QaeFX1jSnknMErVfH/RP14M0JOOrMgOQXkr5Y4IWjnAWzaP5fK+6flt8tuMRhHjphi
GtdDwBK1Fez65YCp9u+RF4YolKz/zcYEWyTw5lSv8rIL37AAAsYffjA5tET8C5LeNIjbcaH9hr2t
AGy+q6u6plnnPCWFNRSppZNmez9Oa8jiFX4icwpAVsgK7cpRLIMgblp47aDIhpE6+fUJJdNv4YB5
2MXASxgH3m6FOKIZaQTLm8UmVgKdMTtRZ6Opf2TgXAczjfGSzFiz/3CcYmnz664iNqI0BEj74+HI
ndvSY6BxwADNX/cEo6HzzL6qMmltwHFfT8SV4xYJXGhj1QnppMpyYaWCE2APyqSZOtKDfxf3gLmc
7/0gmU4p/4UhtXWuKHNdiRrEpotCBY94wVkqVl1PL9NJflSUcGbMuRAILjk+2k/++wI6ktI2plLr
3AJ5M/H6lE+Ec3G0/bCMhPY+5fzF3rKAt3vVmOyrBKMB4nttXwI53AOvF769mXb9u3o4PHpfrOBV
VxYY6u7EwSWZ9ckDP9xURYgdJGffm+ddcJaVXl0Sw6ShCSPSK9kJf3tZCX/Ba+ZXF7o54bvlvShJ
UWvKqQggTmfKADEPiDV/wycgHxYcLzCUSjqYEkrARd96BL+OG+mh4H96lGZDffJFJYZY4CjOGniH
gcLI9fpcfVD3IpJYYejO0yv7RHYHP+QfV1kLND9MHA1uLK8TO6MDxblAensjQK+mUlPZPzCQw8lT
SBkriScS7Tvz2ERMCMikX/M1EIOF0ENSniRGJ3aFeu1cguPN9KlW+CMzO6ko7XlS2V721UjXsr7i
sb/xtbeENpQnJE+SOio1DtxCOSsxf5KEbCCiXH877gy1SDMfzG5BP3BehSfJSvh/GJPzTf+vzWX5
W1xA1IQdtuV1K8PMVAXLAQt+AjOSlfxrsxs/tvjlx1xBitHMgZyiiUgNw9agRP1rXLljjZMWntY2
zdPCSr5LOk9nrvvdh8eU1sYy29kpunZ0c4fPMkAKAbNbB7w6xIaQew5A4xObpPpOk1tPG8ud7yjT
AJJEQVb7kVJg36pBPjTj3yJBlI8RhGufkx6NYMeRfpRmJmh5rXtZ0fIN0pZPCR6N9nEnfd7bscwK
dtoLe+A79KNc7HxSc9Qp6sxnxjnoDLEZrmH98nzynZMjKXf3+fU0h/qgcXw4GgEh5KqFqdXtG7pi
V0isb4B8bNbgFTsm/Azt7ubXBef8ygq34atUH5tN6O8RCvCPweZynWTiDgRP8693l5qB7+uQoAFI
9Ph3aidSxLmCcSe431xb+wJv2d84+0s77c1IS8iJdS8Jquraf3QOQB3gS2vBFcfKVCs6eGa+eiv1
42BQ/wqI4xUd1FuLD9uoAiZWySmDs/gJOjR5AJnuzhm5VJhpEosWCRFEAnGhp7LfnIXmk5BV8U/+
oCJDKvCHtSb9vJPYpxO1Vj6G49QJaEvMXWmCc2Jrjma8wJHGoz82pyA7+X7+2JsbyTwuYtOui5uS
bcn59rkNY4OvA/N9pcapY+H/okZ3zBNDlbjug/XvAHr5r+ySF0WGxIuUaTrLQi5E4v4xNcD+v6Lv
IhBwlCqcbwq0E/GLHtkxUV+ODFvpITqoMC/UncfqOlGlbeGL8ZaBSxi0ghwMmi1rfu/hUFI4Sq3p
YW+TWeY6Q7cHEQbGQO4iOrEbmOQMnAvPbGsIzstPJSinPMIwAt7S54cYFoB9Wm+urVOtUC/YR3iw
NeFOrmyktcFDZx//DKx1R+NCi0yEMQ3TtPlhfRycczDbDAmS2QsMXBw8xfzMrzCyIdL00Qjo8rCY
jyP9LwF7pfUbT1pXIsTwFQCLSZ82yShps2NdD0nXconQ/pL/fmyfBuQVbJLYt6b1X7MhwGJ8JxEh
y/Ga29jy0g1hkqHAgFJ4C9ClzIL2Qxn9dHmewqgDN9V/zGmBcSYQieXwOaUfMfQIKc+yy4YydxXl
1cFAc5urCCLvrhzAAh/U184hBGrx0rziBOiGfKhLG0HHehd6vbWeX+dgSNE/+2lU35gAVGRf5fGJ
HapLGJdycTzRQrYjb0YHPTNEOpRvM3o7zcBbEpigq5dXTC3Sdkv27kIzFzvQAeOizKNX4H2/WqA+
jWNYenUFvbvsfi3vXwqfmcmZPHHY5RQlA2CVpXrxwUWmB5EETV3ZywdU7i+10UyyK5pgj4GxjAAz
6F31KcORNHHGO9RRpRfMcPnP+/9C9VbwaUpWZR+bDhDq4lwn0gZiSa8TglD/VFTSLBno451UoZ8G
Exjc7JLiviX8XV4QT76PXNzzXD1+McPXAF4MWcgnt5AV/32BFwOWB2TyFjg77N+uEtb3A4dxKmrM
TYQ711kqRqHn1iWf1V6TsB84WHF1yg+3I/4WS7JHgCFt0UUOEXAZoYeM7OdCCj4FrD9yt3RjZ8zJ
VyB3pr+mt9joMR8asU+XKPh47uxNpVlVh2R9SJbv56jAm1kAjghQ/LfwWAKQ26Pc7jLK70hA6olb
3hT6y5lnC2jPK0/mHFk5D8zD22oE45ey/z5hH3Y2hMGqFtU9mgaxXK1CxNti36pRQMN9z7s1QsIE
9d4zQ3SVDbbfT7ywR6OlIhnSVhhbt9K2QyAExFwLvTwqOLSrsQzNPkkrn7mqRdMeCUJ5y/3bhnoV
1rOh6gll1K5OsJwf6pgA1JExVDa1Fxe5mnlc8IeRs2RMjKcbbEysAQcIkuXEXtwTtav+BGaLJRsk
rUgSneL6cVEOsBQVqTDWRMjQP3IHwtjqNa6jm36vbqRO5Q2FHHUx5nQMcsveq8wwz7Pxp+WMOTg4
a1WmSVPI39FPRrvy2S9MT9rZ/Q0AJkzrTRZQp6AlEuhZDJnl/pKi8kwfEOGsIFiGtI8qAJ1ta93m
oFweNdQeRZdHPFPDP1vhiagyQqJkeXCzfE0cdcoqawR30j1Cf3Yn6yFcly10p2+IB+f1KuBLwuhc
0xN6WRFedCxoOFJIF/TdOpQXRqpCe8e5G+U+iZ6bi+BnHrPTVP4H4lEQQNSG9mrYrsorhXTVKWuS
yWpA/Ch764BjbJnmz+qQJXulH5uYnbOdBbnUdwhoRudQ2Sg/0NZlbG8LTME3DM8dVJuVzkEkXOoR
bWWoucVxEWaIeMczGtmEHOOsSCBgzpREwV6GIuhmseE4yfhXA3GlQLKV96n8Q5CH83Yv2lDc4SKf
8iVEkCE05dHo2KrgOTlFJXhbfCOmd1NhYDuXbTn11en/gkWOthMeqUGlXqUzZNdV7JhqrFmbfqTM
LpaA374gez1XplCQDFXLkj6eM5fd89jlHPk/GMR1ShMaPp8/axq4VU+4G1CfQa1cRB6vqLoRO8G/
5q/Q3o7RFcAQUUvaXbbpT7t4nOUIN9gmTTH32sZ7tcgvVUL48HAPqs5BRQ9rw/knKP+t/i7AA/vp
cGS/tDLXL68CRsGdGzV3ZTLjg+svUW0DOTll7B5mWcRwgzu8XMvG24njIIZxMPm8VaRWwi9VuZJn
04pxUlnwha3CFHCYkKOR7Ff31ivPbix7NgK2nzpl2LlyBSFp6YShWizQqcr2MItAbV2ld7QSTL93
zP2BmXrlrE7msV2R302BVsgtfCPnWd8iGGqoXbQYVqxhZS1QMF/gLLB3mfIvoh/qm/Kuv11mUlHN
XxPg1pNjpZnMhSQSaNl0c2hpy2j0fVaczz4weK32IGrPQWTxjmoLrFKUc27Aw/Zmge+5wKvAmZQo
ICFmTRgXGM/CBBaIES6ajhUxwIYhQkBmHyQgh0vkIUsUQHxMEgtPGBGpJWI9tg7SdRQ0zc9h1aV8
O2d4lUHH15yDsS8IU3QhvyjDx9d5Hs2tsuj9bIiymKsW69bkfzEmRqN84LwwTBH0qGk+rp1EdX+F
c+daRwcOzUyWo6ml7mWPbOLxg+xw6Sv4WKF16F4HfZrVrIwJQ4rXKeyL69i1F+NnijWmBVVVF+ff
mi9ixOQ6AlJYSA0Zmlk2WCEyCGtUo6mqo9GvKV0NZlSY1tJp4tSrbgJBNSjMVBbCMy0PZ56XOViW
lC7kSDkA2yrwU8BCwh13em9hugD/bghnfhAhCBXXJQjdv9FaFGitYswzJIa9/EU1ifK/LFvBR3Zd
aRfXQdMhEsQbl7g5yevgaT68wAtNNE4bH2v1mnZhIs+lBqAuwANGKf/fLSyaj3WUWj54PibAIYEn
xwKlbdHSbbpWClT0KENMPW83omUH/SNKgdkZaj5H3BCnsHkXVS6HVBKXlfmU1/MODNTmENo1Rv+u
xXQ3UBq1v5esJlz2mo/+Ea4I9bd39FzTZj62n8rShbQKZf6R/LupftvDDeC3T7eKuD9lF5H78fPw
BCNeaj7V9PGOkoCxBNg/FL7tI8kJpAjorbC8CAJDl9/QJ1oE2QqmZ7pPH9SpTDvOIeem+/jlnREU
AIQW7DiWd4ECGYkGUuuv0U8lb/vjCL6q6Mr5JhCZy9aHX8Jn/q9+5W1wXomkyjc5vzJa/QCTTDno
i6ZPhmu+c060okZiuuixivUTW7u+kD7nRgyqO5h+BcZWCLi0G/f5SUi0UYcAPPXN7/yfgWp2t0kA
jCHrXghpHxiVABXut+45fwRP2A0W1I1CNoESgLak4rRSVxj7hr6u4Iw5BA4CowDn83l/ESAW+EiZ
2RScvUvo+R/olTy1CXu9LjDxXjyjb8ETGQZyRJ0vnjeRn9+k+np6IEFPjgCFnVT/dC9AabCMsTLs
yVsa7LQFJAv/xI0x8HJHET4SNImArF2AA7CW5mu9yuV/rUvH79bvCFmtKEB9a1CmB5Is8E6+pFlj
I1jA2tE3wjFXIAAe4hVhf6r/ugeGiLVm9hE8U+gmHYE34DRZZNUCRqENUhWFVrZ6ctd6/zKIaH8g
lHZtZThgRBlNSb8ZKdBMxRLXavnZ70o0cUARrmm2vrc2rWc8kD1bgdXBYHe1+snfd6+5OUBj3JRS
cDXbduUv7aPK7lzgsFlY2e6exWdOmkTNXLwavlwMF+0Uj49snlXMyXDV2aKc3c2gtxRP7Ecfgsy5
yX+cPIdElXLM2Q2KQg0a5AEcSkf20bUAiNnNhuu4SYbWHwjnna0gUiGLwds+U3HF+fGtRvABrdFH
483RRYEv+T0I7xj5M2BvyuG7WyCm2d12XQdgiqeVIusg1umbkz1czI8bGbn39nYqpYBTe3/a4DvL
M1YB/tShjGomvlISQ9r8AXoUy1rQ8+I6/210FUMBZz81Co3X49s6lCp+e2VccEiyddAJUhTZb+ih
v7hNxHZYh9rAizR/5fVE7M1HD0r0hJQMeOorE+LjHI3CqWCBLNy5rEJOACVTx538bZzPS+sOt0XO
/HBVsKwAvQWYbC5fU+8OT0dbv1mm5oOZrzEYKwDdrGWF9QAxL0g79iWAFzZpP3XjjXROQhMblWC2
YLjKAqNM2bdsEQp0twGdf57vVSHJtZ/iF16iUtU1S/tQAzmoR5mszucaVneHNF07ob3CC75pWcs2
V59jCl4Qa1Is/2qfZ6gd2VwnMsbfIkVl6SLU9MYTB9DWZhyRu2OGP3VhkfVJ58IJ+GG7xKKCtu1G
/4RD5jwZMA9X9gk/7Z0Y9xnCa0at51vvCYWc8NEMbvQUhcKp7AZ2mOUHCFl+ItyQmXvBeejmV3Dw
yptCcLA3otjwb4UXY/iZEBHuK5B0p+7sfVsg6qb8cW4L59No+enFnPpymWl/aLVqZUOGUSfG3ogh
PtEf5Ga26RuvhjXhbsTQpeJA0xTx4Vw1b7Q7nkfRdZCf4KyzdnrCqIunosUEcXfaF6zarpD2K7Uy
HZ0aBewLzKJK65VUAWrYuT5Xcp9E/Pg2K9YWjEpPV9UHsvWwxf2qBTwpFi9LT56NQudF9jorFbmC
/OsgDloAyutKOyg3/+KovBWpjb4NKwl7AO0kptKssZWsvg1aKGmxhgLaE7VQsIL6cQ/PqgSK+2nn
Gi3wBhV6d1WT4wbHStEmgGRrEnXFJ5zhP1jbip9hdYRcAwCCzKPgZiotKC0xVDRMhmL64rU5gIud
UjPT0Jf+wFBZk7k2QpepPtwmmdfAQkmL4vnQF1neWdXRNE1BRJpi1BSzGvgcjtjUgDx3VJpajekY
aWk+ApBVOGHuXF0zD/zkuFv9rlW9O2DB/M82EqKJOv1OA1tbohdgkwVIksjNK7tESlOVO2WF1B1x
4W0d1932SwLjyRTX+XQwJSHQbTaDo62n5lxUpmedexi8NXsMuJPqSj8KTbbLhzDRqKI84pe2/YES
HOWzwhmxkP6kVj9unbs4HhxJhU/etZylv8POYAzNHMX3MWWzx4NRpxgYKKFOm92iNqYcJ9cUNGgz
oKydqO4ec7N+jaPu1gp/xNVYq2zg3Cl2hd3eGi9jqZiNszlLV31PxCCEZwxy4B3QjTdu+ZmX5J7r
wcwelU60ZZDH5lgS8SKqofb5a4yJ8+F/INpuHr55x4Q8ujIGu5UE9VTEQCk65GjA23rmXNhcLNld
4Gd4AsrkjHfy/ZKDDsZdFNFrK7Gs80+4Lj1ybUON6y2W+zwXZKL6ybsR5No9nN6G/a6lPbuAjDJf
TBiul+XbGDI2WaUWn7whkYfB3fIToZVvk7/Q+iib9RjD2Hg1ObeYXpOeiFhakvH32M4Og2idaHkP
lbBDDYdgEodmozUCfGEs8xzy5SIU2WI2PKp0RBN/dBzFtBC/O5Gs+Z269+xNGUFkjyw5KxYFt37n
OBniQc2bVwRwVzdSaIKKCxEYsZU0FdkQiNDyibLKb6zVKCf/YiFUtLwg04wJ8StVJx+/mSmW+4Rr
PZ3LUDg+mWAWRTlzfj42Zd3n6w6iufd+CeUZ1LINy/IlJ3B9KtA83O/6M4GtdlizGECwMmrKmRqw
o0quDqu6yrQ9UEOsGMXsKJ/nt91XDuueIrv5W/MNS6tTK/EWXc7gDpr3llzDz1qA42kSbGYx1CUf
avSHgtOF/ijVeyih/HuKbgd2e6vMnjZtmSwHn/CG/otlCjECQkV2WWIVbmypMWJsyc4cKeyYFvR4
xdBzoWZuXXyS2x2InYK7ptZZnXtDXx2423S9PFHANsD/YEUl24O0qd0JnIU4iFrE1J00ojMJD03y
yLOGqJp+ZYCYiHa0XWSdl5zwGxPTfauQE593IRvZVSqKBqXuzR9mKqXaQOIySmMUnbTR91LWmN0d
2DaYYzdu5dwaQu8XJcVlm/qy1LIR8Pj25mkDoygq37y0ioKMXny4MJZFbVHILy3pPfzTd3d1uDJB
1srKTXVsue/zPOm4XvO9JReLFb2/Tawe61t/8oA5NII66mBzSJJEPju+53oFh8KHFYxSbZ7jv88u
Dyq5EDJE4RcMcfkYAHprG/DaBkig5A/d21Ea9fp9hg/L9Y6xITGy2SgKgQos/JoIjjoulsHokCvV
GzDvYlU+DxsYv5yhYuNBE+iW7Rqy89f6h8/5xR6KVqa52/2kBc41Q40vQT1LaVPC/FvJsQlhntVP
+aGZKZPckeD/HnqhNE4KCe/Cldgwveh+BOifzm2fAPJ0K/ykMAdFA2ogeZcGv+9mQwcGZUpnW7kZ
72jpedu4vAGqKzBUx5lZc3oLKxi2Kx4zSrZp0qs+D5oivMOWtShMqekr0F90YQamFOxR09OA4rI8
UYKzYT0v8l/SHKad71BDZlWeWIVyCrO+sZnlYrxQL+qsyJtHGwMeum7MMH/JvMaT1zYAcjzUN46l
NvZ9B6mNkB+RaemFJSC5jtccjiOITIbz5wIufEmHM4A/EN8udRohCe+5ePS+tpyD3UPnw2IUQwaL
mSYWhSJfO7bdazbt9hjAjeyd0MM9WghIY+dKdBaY0Mesx4TN1OmOnlcmS98pNYjNOx5L9Yy/5N7H
wfOnFtFUylqkcLeg2loDTbZN7BdPU1y/EbaQaha9PmU0SveHN7ZVaVrnE8MfAVEyxDIxZetoqNC5
2WPVEfqw5ugS3LAqrC+y+/zEliZq6M5BEO+J+8YlUN74cpLJnmBYddrOdlmi8WHx31nZxa0Nl6Vg
Am1h4oKlJcBkcgfYwVmqrJpa+LaTRpxUA7ypCGEyags08Pu/jaB6tc/Fr6EXEOWOugwW8jcL+Y1D
btQRgx4oW330vYPLtgwlSYdHh/PgEYvIs6Ix2In8+V0HqZ7h5JTAEfNAJA5cOMz4YavjsAkfBkbn
0Tm9RE8s7ApxHa8iSl59pPSZvVwicjrOWs5UZf/aTPBMfEYbFxqihKZhxHEK9ConzWumP98NvxHn
YvRlyT7xGra7mOPslV/Glb05mwEMkzfJhVh100QyDSr57rxIauJGzjvg0ybk37Op/HBsgPb7Huyy
kdCeVdq4kTupuInP57keDetTa2iV/GUla3a4glp1PD++tfcH5Vj01o8Sjw9brp1X1Vc5DGa46Kb0
nyrmi42PnYCXlWJ/HeI9oTe+bmqjquymmUYbf4cJUZm2pdt5yO9jtBxbx0nSa1GHRdJv2+YkSyvS
UV46ONeo7jM++9FLNzpkwbTnnxiXk3K3mPZAjeygxKkUM6I2bsLtxNXpzcb2Gb0l2nPf4yQUFDyY
3jMwB3SI+Zwy2mPYI8IRmQQmyM82tcLrLTgJxL4qwXgkGn5o6ih2CFNFDIUmVSe8FQzu28aszLKx
x6+9cgy7B9uM52D8GRmGQoULecpsNt1CxHMWGWDth/P5vsYZUTZH+dXhD9g2vuDPzJiiMUph7wRM
C76es4AufXYyRxTrbXJTTfJ13ptdJlyaqH7tsxzG7imbdYRW5aao1qAGkhettonVokVLk+eZlG1s
Y2Rj+Dg06v8z83BMigNDBbJlcMQedod5p6hx55FhbpYa1Xr1okWBArnNG2EZeLwKtrRkrgGNxjmA
lucLyfZVdqwNXoDpjXVsWVEW0Rb8YjogJu2qmSitg1y9kUA74HcClLJxdJvhOtRH9Bx/YhN3md7j
ZRYxvJqHev1995UFR0y3mb6lVgEn8pKvIeC6RzjUNBHd85J84ooAkmU6r7DSQ7iUrUNGE8YfdmAO
JKIDAwa/D/Q4KLZ7sFDGSdpf2dOVlb1aiO7ta/vRWoHBnjB7nsznN3Lz+Ag8xEZ5PaksZp+Fx4fP
0h2oQqgaSRVfBshSIhwr8WUuh5j7ULEQN5b8taYzQEAR7WdosFNkAc7mHzO6MilD1fTNm5ghHN7G
s+uO/cqM4CkKJRFqNSin7BA5ZYScJGcQfDiuH3k5qjMSNnNQDEN0kRBX5pFVcbT14ULggWVanAnb
Zc2AV2VqiQ+Chz4yTmfXDgeT40bpRK2oqhVxOqSjvII5H2I8IDzWqUxAqNgiiX9djsXt2FNkCZ+s
1R+p390VI01qLs7Wt+nJ+wB+uftBG5T96UR1xZa9CkKXlaqQJqJdIDOuJZ7JNFilx2uzfxQ5dH7k
V5x6xN5bvCxv3q8g2YK7f0bbvYBdvmZ4l7j8Qi4y85cvu7otRxsI575BCbvu428Fbt9Otq4ULYnS
qWat/5z0lbPx03QZi1zqQGUVc1jChYcnIxy4Ze2KkX+V8FDdsuTxP7nBkva3CkOyli2SMwG7HOdF
w1rpeT30MXNXc9JuWbGv+0xOa8b5/cKevuLQu4VaKZT8jr1sLfLXNx1NR4mJ90IAZgZ1dQv36t3r
rcvQf1Iu1wYK4LbxhZVQ+60f0q72sQPXHTOaZDiG9DGCoNW+G/A9r/RztkKGFS/Rsn+AF9dEj5yl
cYDo2d/zbFOoMJGvf6fv7DqE6XDG1NC97jbxG3WYRIoGdxuVx9u6tkM2VvS32bwjMBi8lyD2DCQI
7NPBFVu08LroXCwbz3VPonj+yLiLe4EiYXrqFTtrPZ9K94QiVwFEDBZEpOC0kwb40GjbeXXQoTKh
BlHkEGAnznfF2SdTNadThQWwtP+n1lkrxcCW9rSx3y35QdMELqNNY9PYwx6BsFh1xl2hB+FyaYZk
vCiZ/0biFUFyRk3d/a3mumGgw4FTS2Hwbrw81SRlAgmG9jEkwFiks8nAzJ5IZPy5ykgUu/m8pmd2
aiywhCHaDzmYdwHQTcrQ339jiGSRKq6HHepJHRaOAY/oqcDxPTO/PYaNfjDn9h++cZv/naWtH4l7
2IZySee6HZgsn/LuB5M7ySKlBCvq++uBz2rxnEboevQxynCclux7KJbqcv/G+Os69NBeo2j7oaRq
lVAJJWYWPqMS4Bk9zXcppXHJrJohPP/wqIUuwp6yqUrYo6iiJwl+yQI9Gg71zuQmsDjZryjFGDRQ
/R5T+1eEvDRmNS9T9GXzv94Pt7sG/CcSfcrsO3GFRU04NFER8DlV0SJTS2pNuN+UNnOpJKh7AJNb
T8AmwJjXhMu8cQ0IbRCpFYgmAWTMlViwbWUR0O3pUTVvFoK6jR8Bm+os5/5jvj/2CnUD3ukiAuHE
8SZmTpIpE95ch7AcvRSJydW+Gt/gyQJkZnI+bH+F+A0Gs34UFCC13Y/5nNF/SwuM7/zE7ho5iHGr
zqCgNTxs9ywCw6JSuriCKF1Q8bHG1vTOMCrdFMFNQ6ABo5mYuYGf9n/DSYehVIM34rV7yqxuEcGo
i0LvEIYuRlc4O37MYY3J8E3t0HCx9lNG4hYmBx+RYJp/ccYjQCTaXE3ML9fk6PJiyLVnR3iDEz/E
Qjy4ArXteJcFKRB5lx+KN3Ey61ef+wpLidq3QpoALFjQ+G7gRUr6rvSRlzImuMp7getC0aihd0mT
v4dp3qav0UzdtwOqmvG31dEaO+5USdrDXacyKb8C3w4pLBcmVL/jAiAeyB38YSMpfulN5duF4krl
q+Ee0/SAfBEuRXuBOWPcN7lQEIy+hM3hmXtETfR0LiBTut4sZlHt5+XXDgmP3bJC99Jk9yxx6FIB
9+E5CJ40nUNzmUKkk9o0Ch+5/tsQC/VVx05spQzUexfgmUrjavn8ImBAcvbC9GMvMaUfAmC9FliM
x8mhxPLKdDcClg/OtFcbT9b7VsgltxfZualZw5WJ5Xdv1sDAJts3Sd0s9xrJ512nUKZkNnD4uh/R
tyuEzRWroA/WdiStwurZtqlkw+GvngAfPsCGFwm2gGNO41jAlASfvYtdl9kJxYgvJ5nHnaE70Iws
+YvQBkbzSw68Yd+6aIALWh2Lj2A80CjRVhzuX0JuHwYAei9BFa6aTveDg3bl5gjDff3lR4/WwTYP
Gzj0pzzumTt/S02m15kqte8BhiMJ+No9DKep9HR9HWY2UGxqaOqZmcuuIqA8GfSxP7z6tjyQ9GnB
6dpS+ZQYw8341m47pEkjbDKfzTzEjzoIBm5uyqhUWjVnoi/xZDobXrmAhNJqKj2RO+aINIwmfiJC
bJ4U2MVX3lKkVmpQJs0nyKeLTH8SBe6HNzjDOz2aaRi5cmzHCTh9pSRYDatzNE+P5dguMy+qIsNZ
ugoI1i97yYK9Z48aTUQvLauef1HTBUM8KYefeG4Odkje19K7tKAdHJtjqIkpK+u0Y2jUhLr6Q05Y
E5c0aDhY/hgcYNDhI7/nfTWA+E1gF/FwicRi85S5kEloaI5DUkJt2FbKZ0huEwvLmhd8IVvREY67
zINL8MHIpH8RW0h5QhFKCjsL0LrxHtQKEHy6JFx6l/g8vUbnExt4udHqqm9bu1qhcjyuQRkVPWPZ
WQd5sQbmUHc+yiChQyOF5tohKWr3dJQHaLedC1bEwcxHsxOf7lqY3h3iRd7B0rqlZut31cps3HlI
yEKinOuCtMqvVv9+X5JlQ1HwTVxJ/xxnlmv6ufdh0xqyUP0bd7eaRcjFgEosJQCK9NXvuvmBIAmT
J2j5R57FH8a7FF2XkXgveZ8ZBef64kVYdJhEJMX4y6iqgY2gyhIFXdvl5xGGeXDqKFDzmKu8ZLZZ
V9TGCuQTr+hcYIFGjdcJpjuL/8lIzLtPB2qxbgtwkwSW1ngrbfiv0AKXoFCeegavCuexROt9Hhxq
q6zdtPRz65+AFBx27MhhD3nmiKpwILPR+IgK906rWQx6ek/OpL+z53u4L/9QKehS41RlZyCYUQYO
m9hb3mhu6/yLjxeBwFvjIS+Cg1P9PtQ/v3y+oTRCx0QfGfo6SifX8u59SKVmTrgbNv6MZwKCj9tL
Xue97/4lS7hf3AiA3KCc/DnGiKgSleO+W8ngHj//fY8tuAHgUFgrRRJyPYu5SFla7Kwjj/q3ZJve
+76vC/jyOZYxDw29CU2at/dUKOuSM17ZJ1/SnJggSohlQqJzaMbzYru2iiLoOf4oo4QDtoI3Ya58
hponhbSdTqnbbzUL7qdpr+ZyOCgryQqEZKk1aJCvuU8tBZ/cFLP07YPhyQOTvRP1QTnclbXCJvvi
RBlEIHyh+Kn9JWwgNSD2yENIb1J/y04zRhEdcZOr4phC9kjcethfb+gXSTvMABDSK7M4JBSSlNHG
9IzTdwv5u+e6JPEDi5Zr/UvB2fBIW8SGeOGsXx5uRwGQrfMXLCDQbY6O4SjZ+8tlpD8HqwC7j1K1
ZG8ES3omoFr2NKg/wmjeOuUSahNxp1kDpmQTOY9uZOZqAez7hPAyatJLe/OWPfyCsv/KLPVt+E/B
k2CWJkC0GFbxipcFOG7U+hdJzSRM1vp+DqyHu3vFdI4FJZsiwCRblj7oqTQ0pElErVYQe8lQaECr
joQdOVcoPjK6Cm95y/Hb9nRiZMgdbjQYgMpYmy7vPXWXAtmVLp9vLf+9G8AFNpu5tSInPgQkOBVO
HQk5lGdxQQr8ISJWJSHfxFuB3Czfc5rcDIrlbB6Tp9gguZwsai2rX344cIgy7q6CRbye9e/u2OUI
EN96JmvNtRfXcib34IUbErSogwC3Ev/FEthtaoTusvj89blfJjzLq7tglIiJxvKxt6Z0+KYtuwch
2yKn2XJj5igr2yX7cMFZoG/xCmlHgPamQIScxHZ2FqXbDujtAcKnP0HnbgtvXKHHkp6iLXKjmDGN
c9a6WXCZ3QXT+KuzFF00OJ04QHXskOXN2irPb9Q5XIx6paoKLpe3dwSUVEfXnTJ3gKCkibAlGBIE
06HZtcKXvvkx5iVU/jU90p89QLPYv5Eq6wvMN0FxWpU69kGxfSQIZ5OerDuLQs9UQGtQKMIQJyxa
Xc6tKggtJuO3VbWvMLtUTvS+QNOWA0x479tDWdEC2GOVofGubSqIrNzHLti/tIBHEPUmZG8iXvPa
TZGVRygTYu23XNkyCjl3wq6rBrJVad+slLxsWcvm+I3st1QrbPOQnfy4PU1ZS3P3h8R0tdI6RNOf
1b0bNznkMwxe7tIx68mmEQKjR4erP7hXvZldWIwsMbV69IsPJbkuPQJO8zYsb11k1h8XgAiLP/BB
J5AsIciDftBlbDhKeyIRZnt72uZGflJC2tnyqmggbwBa9Rs4Rj2oBNfqcos76NPsuvTsJVQN8g47
iqmIlhCSUpz5N1BcU5d2sY6LyojPgVJn9YtovcMH/CiFJCf2qC1TQNa69IqvcWvreTlIdlcGkrm9
xq/OpWdy2KKi3FqG0K9vcIwjnnxMxzvG2hFTCZH7E5DuSsem/9C/kKfx4z7pQE9yndIKk+IsDWQd
cxjwrZsI54mbh3iibC+uqtOjWzZwDn41yGW0FXvjIMKvdO0BJt3OLPsGjJi7O53PW4/Ldk+gZ4Ag
KptnE3LXKxHgz4rRrCSkoKpzsCav4K5WXAO5EZXxD0q/V2Nzja6rgqnC3VwuczeNOgsjc1Lkvnlm
fiPH5QDFJpMFyVrRYvRnxEslytCpou9V0+XmSmMKRz8xur3Edq/gfLYQuP5Hb8nLmLxZOmB5A+rn
qA518zVgkx2C2hK03G8CB37j96KD05pos8Ubmp77Avs+iCUiAsFf0Kw/V1YU+67ZrjEu0l82M91a
ud6zQwsr4S1hhPH1/b4Qx/X+PDWeN46OywRgE+T/DRW19TXk6s13resIPRkhjbKgdIPD0LQlt/Lo
S5EM5TLOZr1aQzvNwEtsJ5TXQcvjG/k06r+MXCOoiQWL9BuS3qYKRE+g7BLjPVWfiezlI6OZrTiC
UM4/gMmDPokqeKtceIkRFBCc0/PYXkVWuPwL68NdNHvuWRLsh6nN6RWUNfWe6Pshu5WJi7Ljo1wU
B2o2e0BTsns+sWssKjLBUtTHDAqYjAcvkxaSZTNTVUyKm7nmEmYF0no8LQMP2f6TSYlsfWzYl5iI
ZYFTCtm6LeEXNeoKGq55G9MY+VlKTpQD45Mupn3nXlfmEY+ZaN70DwJ+oYu0ajcktN4AQ2vKNAeK
QZ4m0KbNGI2P08sHguqfChnCgASYyn/vmaWHL/uhO+xbSob0ZhTMkcILL2HNYuMmISf69T/baXTJ
q0TvFzxRXgw+ffymnIv9x3xQtcYZLon6swxem/8UTXx7LdcRksYCGtEPFvofkEbNNRMNxbReg8/u
j8rqVvNnirAuuGdsQgXavxNphyCx8nPfoIRmzdIKHY5ua9GSzlzBgXLkaOh/l5k335lQdWHDShWy
fBgDpB1l4+Xzeh8zQiaDPLrKygN35bgpPu7fvJkHZpqvB5XJ/ip4SnyxAreanhd0Qx+RCnf/cydW
eXZcOoaSSDm/+8Xab66B69XSBTpNmSWFJjAoT8ymRyKSZeet5n7oaVKG9fZiIwzvKLj/dubWmU+b
wgemqPqTBIlKDgtgjvLT6PRtrESw+KKKCD3Tx1cqhQ1+5gHBBDo48hOmRKAsWM+1daa+vpVl3auv
sF0HAZraVFn2fx0hpyf0Dc/NTPwmCsF1+MQhqED+l94PBN6OVbYDy4FuanGeoKCOcpO1qQ13Rl5A
NKjipUOv5Fm+Y0rnhR+FiYzdgdxylv5xmchvrpIfXFpWUsjEzOOQjlujHPuBmKqi5+8x/95Mce4g
Dvpi4Wc6NR9nztQSmnVccIXcqiuGOquJ2NZauyJJLQu4HmVvxWOx2a2VY+wKbywzERTThrW11uHY
IgXnz1+gt1KF6X1gOhNfNBot/Qdvyz2+sflyOcVjHW84o2KCGZOqgPJaMuGKLYHD4HGwtt52Gcu/
RxaPLZDPBFfQp1ZtfdfMC3DZxoPpXHf1Zoi/iLaazq0Kw+RYRsLmM06Wf4jQWo1RJI/JOovSJk4G
+odhqBd+VkLqxTE8vq0qrDdN5xqa9dfersvrGiDS4VkIf9dUOBCIh+aIvqJxh/ejvo8dOLnSjNLE
R3xUdx+ikmPY3tzDuXweenZ97VPIhIMGyeIy7jOp0x+1mjB2maNFeTzaccUTpPoCSxcI1qkAvhDx
o5G2Nu1ki/m7deKMsvvojhMmIVOb29z89jQQBhsJcxekN4zQrROQ72DT3/LegmhOn6ZxDPWBjEPX
BMG1Ax9lkP6O/EJ9SCs8ZN4ZbuCF4kgfSmpjW2HEaE67myOAUk3Nvw8JbB4S7CeDUaJowt8bnyqI
AhO5+AhIxxLdDU0l5h+THzA/0TXKSuWgsqswJdSiUHaWxBp90WNXfqQ8OuONR9nXJ0nBYuxpxjat
4Aw5uF4Xa0qpYlBBI2MhkYqd/k7kwJQMg3mpYCOl9XtHeDP+WqX1p231XtKTILGRyEcOmNhEzWze
3qSKuCS8klZofk4v9vDitNLE9juqu14/Y+c+4hHD5o9SrYNYh84Xq4e3BULnwRqL89QGRuwB4Njo
SSIp4Cg4cXUf0KG4i7b3UFS0dzBLu6Lxakiy7GCwrfXpXf08jwoSmvIqPOjhpAS/VH3bMl/+4iQg
54zFjgBEWqud1HqFNad/qpp06Eeo9uwg7FfkR3iHd3nNhTV9heoNRsvG7RGv30jqQ1lBTPUw+t4H
OakGOrHH1q8CSghUFjOPgyvm9NeauW6VNSaJJg0aBKwK0SwYN9NPqQnIOOmqlbMh0h5Zyqy56+yH
AAc4MieFgiGr5QuVzoqnjj9Xh3tZaWTIcLmMgL6qDLM1gXycudl+wZQTDqLkYyHJ0VGof11pE5He
OlzgiDDAtPKj1GeL+8g9ELAXXq7JWG2TtH8YoTZxq0tQAT2fLMn+Bgnu5cjx/2vv2jvIMdFTwUby
wyQApfxey5//XDmIFFsmVUFLXhprXibYW/jl9wMFPyHwmraGJSXeKm9bGMTgmOfRexW/bbHsCxF7
LGl1T3ssx4Pu1B3RBiyIJfHDRe1i4vr+BFJq8XZwmMTNQR+ak5qTPV9/47plonND4O5nojQeqGEc
eFWY+aR2OQUVCkdOnNgTlLhnAX4z3V+wsZZ6vz9uASm+9pkIxhUOD48Go/fsrhMmPBtzszr/5Kvu
/755o+3UDIbNirur+IB1dn4RwSgh4cufSjCHxUyPs8yPhUo0nsZGGOX/CCJGk/rYgIjG+c6boY8Q
bvIMQ217peZxtJWBZaUtqxp6taZJPUiQt5Skh5EBIEYAScBbexkRvAHDxJ3w+zVLTbv6WrBtZmbi
y9q6GF4oR1kFSdJbRGj96iB16kCUH6lYlQ9unUCvyR9QDiSkKtGNNeBgRerRKDhxBKpOxDmXT5D4
r/32m9gYZYBXCRQs6lU3bQvZ1mDrQd5WUwBOvfzwGrc9als953EUtSyfT64+xwHOa3TMp0rF5N8P
WqRQX5v9aDAGumXeyfoVfGHto8ifCdzCjsVtCoxVqcbFjnWDu8+pTtvczRIcvD7lyX2BxxEKj8oW
rn7y/S96vXnb9oqXVYsOpBnXTJ3+PW3FcXee19pFCdGUC6wkofmWSEEIYr6ooV43/2qdOihY49O9
Ea9UVr5uVVX1iK7IDvZ8PfmAz6HoASg3Rjp5BZnHoTTxDfV/AuOBATyAUFbe4FzySeeI7LdfDkrV
7uK5clLGz3I60VPJ0j8vVI9ukrrDvreoiQooXU2HOwicpbFjnfKU9AbDjHR7xFzSZE3CduyVHhpX
jv3NXeCEkDctpnFVig2JtVkmC8b7FY/WIkpMzsVNyvwFXjGFTmQDk4rdn0BZhKqJ7Oy6O1aXC58P
wBQ3HMmCauL97uDSZyhA4CTgwiuiKp+40AVrAdMSLb0CvlfLHFHMZCJyrQnVNuugXNcLQ6C/KJaO
6YL5TD0ccoSkDwl6RYhX72cTWtNMYHSvo42quEMYK+3o7ZgiaDBam6nXITIEAp1cMZj2UC6zhGr3
Qv3oqhqdGIleVAvaGVO9Sa1c5IH1ufMH+Rn7Hqbq2C96akI0EMh58xvUr9C03YYPeJLl3dnGUuOL
zKBb4JCpBnE590Utyz2XwnqsncIrV7eKp60bsep2V8CFWXhAJMW0u5xP8/hsjXX0C4yTjVVCys/G
jiPZyP2LFEsIZiJckHDJyjo9PuFe3Y2CLcC/c6FvlAHEnz+7H7tlr9zRzdS8HAtVhVpXIkrm9vv/
Um6DrbItdVnuYEuBVLkAPIShEumE94dBignWTz2KDlTULUNj1+nGqHvBIZ8ZbclPVNqPbSEh5VQL
fUUFNZNd1GngrdUomOSaKmb0XhGUORL/e0LBVBMRStp+311BgVRRu2Hz4q/MkKtzyGkvZgjisUDV
lSCHDBiwBRgmiwzyyxIBKKgIYc/WuerBCFYZfcZedikbAjZe71+FcSZUJLpAVlNYgUyxc3KzjMTA
gGIK6Gsxr/pBWxBrv+TazVTtaJLS4XkvHeb+4faUWDRwNZYGSYT+luXfqQiOKeZVqNTqg9ziIynE
ppLxKRJ66V+q8maGsUXZUr+VVkC8EoVZ1VuoiWnjlPcVUSsMMut6xUKUZuAAWTPkdj05pNZFwP95
PxDEMPY65LxNJ9uGGxiKQcUf33DSARrLWxcxKpOrxRva9aXPaGk8j2OPmxzmjJEKDUVFnG8Ai08k
kcPLhS61UkfSP9fFrkp9G6/alhFEvC4zXkJxAGl4+svcrGnKBcQqFDscDMryQ1GyQnfYqmJ4THSZ
Orn+6wH8+e90wjmYMykOK5Psy8aGBiKBvesMQDUQPxEeJKPracZevvmSMwEDpMkdqW58Tt+VTnI/
8G+PGSCRzd5HDKNz9kB2qjDGA0iKluLMw8Np5wFC/nr1lvCEnN6cg2z0L/R5UEtBvdNeiwyYQHmV
nuUQHf18MGrXDpY5p0PIzck6yi8uYRu0YBpc72jfGglJv80tr00SIgN+POFPV8jTGPa954oO5sNZ
s4h7sWFWO8W/AnVi5AYwv9Sh3DnlFtSHO/dyK877msOowXz9t6dDwDKxUFVeWmzDH2+4iKy7ckl4
x5k4TwcIGiL4CDTMm3dxDqk3AM6ulQ620apWtwPNgVuHWQHSHCr4dfb6F7+kBvrkIvlByCXjiPWn
l+fcg+Ury8X2LtkT9qGcJCkxxk2Db2CqMM+2HOSBC3f6iufrH/6iGvSSOrYxts6zKehPogr2/D3X
aa70fjZN3IQBNOVWoRMNAN02iHj8nv+XrMDN+1yq32ylR7qCvWvpxeslNGGEugaps9ZDUhBd0yMU
GnLyflqHZq6TGBcXxFXBZQises3zRZ+a709KZIUpnOCkwNh15ZoPmzfziil57embTzh/2Leihd/P
C/Vztndz9E0nTP5/MRusdgAYbkpZdvToHTS02eDVVMl0cJGfbkHk7eZXjq3MoiuunS6Av3seHqqf
y/yC225sqaDGcWYrK5ixa6WLoY4w25HzFfkUuxEzO5TTMlKaqgvn574REjiZD/i/m+gUhKKYe7AH
MxQa0XRL4NZ7/SMOiwSQVJxOpqzcEui31BT+lyHH8aDnodsMdN6KjIY5WtCpw+mxTltkt0ef/oU+
lDNydVKsYgQj1mXRG9kcJPz9jNOxFs4i3AHwbSqUAPvYMpajHdu9dzT2uOmA7xt/am3wOyxuaN2F
nndlNJ5ne8PZY5/LorQ+KqMO6S9aC40VXa4lJ6qmOZ3uvONh2+wZ5wud2e0i0J7jT/seWMas9vol
7eB4KgwW1FRggThey0K3r516hOl3VgZlOkK5XxICTnrEhdnD4X8oTMdZjbHoFppT+bEAGL3BO3xY
txSgeUifKoWryNX/YhUNvAelnJOvc+mfVfTXMIyAR/KU2vkfhL3u0dLraEZuhUR8C319vw1vPMdZ
CIfvV7QazXOhLhS3h7ATRfdnX8A8zuOFMOzP0Z0WFqVzczP9b+jaD7HZh9JnRh41eDO1ydMRM5p/
4QOfd+GZztVK7LBDN7Bg5sKghC90KbWOE55vXPIJaa3DLQ9pq60sv5wfKQ56V8Eeyvl0jenC10jJ
JI+q6xyvoRNThBMExL+/zglXfmwfvF/I+rpbTpO0mo5I19exZ8gUqtImqpTfhxfH5vdUIQ/mqNHf
cKoYW9tzH28+sBu8dnLeJJm6MtWfFiXzEUsamRg7D+bogNUXaIuyt4x9VIduqPw8Rb6Qkvhw83fI
XcMS3UY0W2TMfNzqFFqfSXwSf3J1pv+jTqFbp0Qs/azPiCCRHSpa1UuEPoyidATNunlGBBoJs+TM
f5ovF9jq+gxxSKfNAfiGUdRiXo0/1tAvHmtwC8tk/oiIqHdMEnXLWuZagynat8Xw9i1+oOHbiPeS
9L4eL6JWB6kfDfhf4t6LTtwQsZjhyp+0Ol8jBvCcdXA5DyXmukeA9b4bTDjn61ncFfhKlGaWlDST
0J4mI8h1C98NalG3CUdNisS5XdU+2G2Fb+lLAArSHDhJd1V6xBW4++JBN/ECUlyzUg68eJ5xWbzh
B5vo+1DpgLlMPUwfsMXl+2RB1Cn2hUbMfiaPwPR4nfpWIJqfDSlpHCTtSUBCvprVL4tidgjl6dH0
iqVp6CCPI9vA6MCeyORnQ8gwGa9Vrxl2JxXM4xPXgxSOa2e7a8rInsu/SzikMqIy9Stx0AqMUAWx
krc3ikG+nPo1FAPF5tgzU9MyzNQUK+6ak6ajTUJ+J9457MJzdztpX//bV+wlGDlVmZpNr+OY2H27
aHtGnxurQJ4WhTxuAlp5RRuHWAiFYKKGXfSfNQ3uL49F4UeKdYgjqTraLWF/9B7k4JC7vxTej55o
VqKq5bT6Fhbxc6d+MJz29HD1tst9RYkMDvCRuaEvo7rgksKECbsQwcf6KTuFIeXn/5aksaTAas+1
9JZep6SXza9sYQmoTCBFG6kDYk7lSCYHX0ouaC8wYkphfLwpP+6d/AbfuzhIrokIgqXxRYUUMyuJ
L3TXKfFMudjXQxsRAKS+BxlvUmwLqwoxznoPf/kJP+FfAuzeedQ4iLJGP26Cdtmn56uQkSEvJIKa
83h9/eMF5JqjA2nn5vVPg7iUGi9wzeN+0RzrOKoEuK0iq+a3J1MEGhIER350rc4RGhMBynKI3xsR
i1DzDVyZV/ljyszjV+ze0LqvEoeF60qlRM6YXLrElInRB9goojlu8hxMazmsADXrASCSe9esjSOJ
oHCJqKv+PrpVwihWfXTjNAtFwnzer8ij78tHmFHBPNSNjcDJlhVkdXah7lZ9kpxJ8oX7B6qkiago
S7OiiZyEc4U4uohO/B74p+0ed6FuLrPoenux/LKjlQ7Q4FSpT/+mDMJGMjUbeDElHMplg8oMr4RF
Ehqbwp4sCDrUq2pruPghlS0pn3cfSLuuOQns1y4h/u2vWqrbepKYHIN5q4+F2sSNwEDUfU5/ALbt
jU6LcIIWXgdp2edoysGcapa486JrDkcsZmPgmBKHyJ7JDc+IergXT3jU0gJFqsAVs232ZfyXRsGf
nI2DrZYSdX+0zbs2er5wplvVIZmPNB1kyYl6vJOusm+NXpjwzQILFXbJEeyqJSzcTQTjyMdEsDsi
gh8yQXZEnVdl0pyHUOZVp+y5HSTdTa/FDcssmf/qno9VdKD4Ur1G35SAwJxOIyS7IL56k8vR0ucy
OM/IIXLjec+wKgve28Y37eOJ8pJl5lDNUOl/zmSYnpl1SmF6VL9veV5FDJNk6y8tV0SBOs+tmh8s
AqHjU9S5CWeov0PwG0U+emlwZ5CcppTbGw4X5+x0EPJ6Dymm+QjjUOvvJsbwbBQRBMtjkwn51U6f
YyWI5OJaLIv2dsQE9CCfMBIJbI7Tpl7iujNWKZMRYXdGH6XNOenP30gg37Ci3Xn7On0k3Km4hM7E
FnHv3B6uMG5l6EnmPi78xTXGCc7DAs9yEy52Py2jY5DRES2sr4dNTTcmYzNrz0zOQsrnkd1GqI2x
uLfwsJZZkUHKt1W5kMWYCguBJXfcp3CIK4jDjP92F+ICfX2fGgECEUc8WrJVSzJ7hSTgIbMq0EWg
CW2Ou2Y5SdIRXDV0K/9Mf8rogqEOqnDVWdHVkA==
`protect end_protected

