

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
T6wVkTPpNtKFC5HWYRGz1pDJeqROUhDmQQB0XOtYU+hhB43DLNvsfjC5KYqU6Qt1lGAhH0laXWbY
sFGsB/1X/A==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Bo87Ik/z3ZMfvsxWdQ0fNuP7YOCyp4j/ygqxg4KH1VshQEFmP82QDe0umsG5l9IQ7WJ1x44Z7hUv
b2TxMUXo+JqxKnlgUE5S7j3ulzSH7GuiH1ZZMyENkBX9PvYGPAoxkfBZKwYBwge7dC+ekfgtgSTi
JmblFBaQfl2z3igDjdI=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
OS69EpuOCXkwKDIJ7c3PBFNFMJbX4CiEZKRiPCWgGoIatev0sXIZ8vRiD53mj0pSkbBqScW3T3bf
nStSylNR1BolV0YoJstQyT1+2pFYhZ1LLXaZugJ/oBE6vqGV5u6J3W5eW2CILy6xHulOJT7cesIj
cRuZgsZzN/xmRcR/wqC0vFpdgeypXB6mda8Kpubf32Dxwqfu3L7BPiBg+o1IuskbZi2Weoc3I0l0
OeBzQzAzru491AqXGKlZ7sf8bs7SXbbzXRpVODRt7n1NjaKD5f39RasUxEkDN/Mf2io8pxFG53sn
wj8Vha0LEKNulGqvG45lCg9sffq+6YoB/PA6pA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
0V7+weIw8dZ+BPWec3DOIbteiwGwG6dN9psrs14jYpdIBALSrfKIpNuQOkhxmutTucD037ovCmPT
7tzlCJSh8b8Ydyh2TEeIpJfXn05PGHs6Bho7YXv+uAmzXPPeMsLwL0Zdj9PYL8wHeM9h3s3oFmE0
whlOV2wA/y6g8Y9g2X8=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
LrKyoRzDm4cxDmM9WZQaVOeA1DZCMC2sBI/JOp2hUeVDZFMUfjL+9ejUV+oaV3PC9kYwU9gS2N4x
T5QckNj/uBm/MDZii4ZX6FRa6E86JES6LqHqCKy4pn+VjDJ9xeobjj2ApHw2GympzRIfTHfg3BzS
Zkqs9Cmo3/2Uv3zdNyaGnk9f0Ojhxe+EEq2njDvi1AWk3nuKPvaX2PFiQqvWXWef/JYb4HJ0Tjlo
v5y52n4XeymzBXqfaj2Y0hccYVFZ6YVhMnGGV06K68vVbtdbUuaSPRKXNa9qJHwvtspPluLhH5Xd
ujRGgNTtTMlfDYr0Fh/3k9HYg9NPc+b+y85sOQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4096)
`protect data_block
UxFj7r5qDiV7p1nS/m6mSYZaGBODx8VuQDmXOkwAadHmlUWH8u0sCkCk2p2uDsnCTTM5CzNjoClj
+EZgvQ4C6eY32BqwlOTeffHGu2F24HbPz+NuJg+8OaPcdvwsUA/p4iXAakvXhpGnyCM/gT8b5m35
3YGKf//9b9375PErcyhAKws0f7mU+D1NDogkA4AqT3W+J+x3Onuxidx1t0dInFEMn7NlulZ1bgYh
avBhRMIGmhYQJ1NXBcYIp2c3Av98sy8azH/4leOiUva02LpG9hnCA45VWNL8JqIajzd0tWd3dl8g
sD5ga4dARccaCpBa30kmxETOSqZPRlrhCW3QMm6PAsFEGkpnyNiBgYRRux8vrQfg65DLxWygGH5i
2ZMVZ0hvYZ4Y7mEdwxvSbdpfOAi5f611TJZlPF82ifGtLtVTrj1qiqU51NUoP+fxPsglnSZ59IEw
f+HaCGGZ8gAsCsflM/x3aE6cYXCv2bWAIMmj9MRkgRVZnmN1iyUiE481dgMonql4r1FsSuw0sEeQ
Fw7BaKTJLg8dl2BIZiKON9E1Pv+iLjaG6oARo4q58G7DoJAsmwvol2z5RIz504V2ZuqEIn3Emw6Q
0x85JlTRTyKjG5R1lJSY94LrTvzOLzWCBVfZbQAiX2Oa0KKjcBBGVDaolz0Mp5mascnvp5C1VRew
i9D+KlCgB8o0gAzO2j8MHI9urutQhMC++0Wd9+uvyBctn5myvlpQRVKQ3K5WIAQLsl3CgDMME4IH
oSS3jNVSa1msTQ56rRj53KclfGhwa+eLc/QljrTgAa0qwyLRPNmVKhn2IkvwJU9+ivVOi0z/NFfE
KTw0LfOuZdMRdDJtvDm1gNzRERNoVTdaBaDCSlkjqCpcF800gF1tMGOmCToM5JjzHHjMHvdgYS4u
a3sc3Rdl3lTifW9yKWPAz/LmFrD01sKYydxmMA6ld5744+jZMBVLFPCOuogS7/8tjj0deQ/kNtQo
6GY71T2wWtiv8gaCfqVJtRXa/cW3e5R5Czkk8cbnhwNitcpRT2uADrogijWYCS9JXmC2eQjmBsXu
N9XIfGyYsS6JB9X6dRQmrWFsT+LcjVXF2DqB2w3ghTIV/hIGTgLMs23ha+I2AuzutzA+RFemHFMb
0+kDK15CYPTZD5A+o+LZ5XqqtPnr0HGhW0MRnXsoJVRmG2CrUVjYPmtM77cykBiBlfBn7BRpDCv2
95NkMxIHcrDaJOOp5bo1xtFQlJLs5/meLbr/QmuS/1DXqLQ0kFR7STtCXN2fhTpEvhGbLQTzRcaV
H5Ylrax1JIOgYfqPC0U6CJpbrF1kuBlbpn8ghF6olOHk3zxdtcufN8jLzXE9FZroRucCi6lodAeT
IH9eFjyqyJ83K6DH9QNCPrTZpD8UUUN+OtT4m9LP+H2Ip0niveWe9D+IPsEK4dj7mOSYsqRMQJD0
CYXw9b/HMge285fXnhGLCap6g0qUlRmy0V3+cYN0YPbl/QPmRNFsoIYTwD6JR+NljS6mu5dOyn4Q
7NGI9rrU1cFHbO1dMuzI2KPFQcDkBHCDPeE5rq0oIRKixlxdklfMinkIWnp1o+gY1br89srn4D+R
QUGvdQoYgBN7P4hvCumNxebOuzlUJWs2B1zNP1QQl2ojGWRjV0QT9WAsZWtUABJ8o76akepCpKtg
k8S2vrAe+oRhHKqGcWBNyc2MY8lpAuIf/NxdNDkj99DE5T9LrIq1QpHrw5gOeG4+HM67RNkZ7ewx
cnAIQm7TFA4mloPUDXpBOGYq3KahcrFS32WwIAWU4qVP57DyzcLHycv7E0azEf1cfNr33vTjGQX3
QNyja83GRw1ATvAycYd7g1Wbbrux4tTx8ENe7tCzxwoJJpXDz0tLT8nn1aEXF/iYVSRJiUCZ4MON
H5Qh9esy1wfxfPlnYCCwuO/9CAj2liIN/TSHPqRM+PhlQ93EMAdiSs5G5bM9C4eGdcucJAP8ymKJ
NWGEO/HmxRnhJ4jANlqABnf0wIf2R7K6mG9kJMYjfoE5u0NVbSGMeZAp3EV/6iZPQyXgk2OpoE8A
mKsYc0Ank+CNwicHrXyaLd5H9hTB5zM+RWM9uJjnWuu82ns/n9nlhA1AMwjtuKtY45MIzK/cM4s+
n2MWB/AxkuWGanJHjHjzzkxDkrSQfwag7fszrujvweEr1BmqSmh0bhL/p/fU5C0KYDMn1t5ZtUz7
sPDL+TvEiszwCdxSF96fB21GzGcmhKiFxBjtY76TdSnQQKpaOygmjGG/zfPQFZvVGGfQkLZehCNB
2tSXbVyh67sTeZeQUic2kF85HY/gO5DuG1WbvFn+uyUoCihcAHJaDqciEFfz3mXt0rLkmUbbU0xF
n7KZkw3nphOQriRwvaE92FLWghgk0d7luxM5SBQ0djK2NJGfLXYWo3nis20jodXwh37eI/yDuQ3s
Mjco7PNjYDms4IPp1jrxgMDHQfYYEdJ5y3hXCkUGTq5ZD+DMNuw1nFXZ9dBGe71QXQnV/MhXJ7E9
XL8eqS6Bi83452S9DX0wVaK73W+3Ldig6L4Qb3pxNzemMo2GjEH3Eb3e3/WJVFB8x0zfn8m2L4wJ
U1ZxWvR5SBGcjhpWqGS+WnmIXfACadMeaqjfZxAS/gtRYo0CGRPfwTduqgmZG37mouYNviONAluf
E2KEW9r8HWepdk/TCQQwus31jSct2ApvXiQohV2bprAQuXHbkusKC3p8lRi2JOXh29I2jIhxdZTS
mttt+Y/NGxjFJ6no3/ZUpnzpQCzawhh2fSrAdxd6rUau7GxS9aXdnKgx+cwomimNA9e7wZa/XRbK
oDhGPgquhiLL+A+AwbOMgKdbrMjrfO4gzyJF+FOpMJh+bfGz9u5JeA84iY15ZA1nTZMuF59eKNls
7c/o8HpBC6VgadM6YASUp66kOPBUG8x8Aj31Hs7L6gWLIF7sFQKYr78AN89o+f5ccfmTt1dTWzP1
eim95Sdr8K3ixKKUb5h+Fo9MxRylyz6zqriCGg4ua1HM3J2qKa1bTZyqt8mtpP+5Wb4a4kjUkgrm
+lrXnDw4rWRfKNz4mF937Qu959NN+nFmB/DFpvftRvCvS014jCiPv0z60tNrlmz5eDZ/pwrQiaYO
6pWDw3jvMA1YKiJNmyOoxXco+CKyPzVEKsHxigvMImg3YEJnbqMi3WlstfKoUNRBqDIhdF2V3voz
XRRrcVgnJIIwm+Aw9SRRfFMSQbOv0AA8ZhxYumrFcaut7jcm0ed9tB9U4RCBv3M4iZuM9j0PfI/D
0vipNqLgba8o0d05HCNdReTLIAzDKRNPyk6W3jspaAVaESN7r/g2ztT1Jzi59NU9djr6qnLJcV2/
QKW34UTLR/SwyQkO+KMqqvynMkc56JIcPz4nysCmfl7Lul/NHWdpvBlJdW3MdbQnNV6rTwLBytoq
i3f2eu2Mpt1aIluE0Uzi1Awr6dxe3xSlMWvFh3Urdc8SrGhB2Zbh89GxcdvwxLTeLIxko1s4g3eT
PB6pbLc95v0H7Y4rKOmoPQDRB3i/fW45+C11GhqNDRz6x0WQRyv37ESJhcbrdZQzbBwOmtCZCRP5
BLG4jw9hzLPr6/o2jHfzE/ln8/0OLVvOzctGN0p4NlNVmu9jrzBC6prtSURp1zKncu1G2Vc4xDkO
UA5rjqWad1JPf7yE9AJG4i1/c47uOtxC5Ue6DJHpvzAeJoZrBeU4JnGF7wU8EzQrFwhROeLpz0ZD
/OIIURmVmFIAAgsRF5zpXx9RxPBLjUwVJU4rYdKztgpqicu11woKLaY2n8LxWyLo5C+1gkaKZNMU
mKjogNTZKL+itlo4zdaYSvyB+7QQNfwJdSJ4pJ4rjUQ79qBMiPfX0iwoDqUMmdnhD/0Pv6btdSNJ
zYO+piTbqEQNu8ZMVCmUzEukKPfosGYbg7TOVBcU6O0pFHjSM+UGHmcszheGT3M2XFMYoYt6dbUn
zT8Xcy5uypDxRSXPSIiFSDeuCP6S+C7HxNidob+Cxu0e6EQoysnrUhCZ9gLYM+h+npurOGjS/1hD
PireToX5vrNhScnACk7EmWzfZdjX2pMYupnwpMjrshOmKxmGBkgyU8lP/ogLMh9j/lDXat1hJBMs
RC8KaVcJfVvuF/eh1dNovo2NnicfKT9Gs6tlpXfbDHORlSHpR00CnqTwAFKwdKGUsn7/nRHoDk+k
/bq9uVbAGosaXMPIWsDYGld/EFz8J7tNx3cvoLMg7Ucmhvi2rMotBNQulsUPf6HzXCTWCBkXb8Rn
bcmOYjPHNG69QTUX/TXA51hmMnpGl4hqG0PbtSKgjq5doKHJXBMkSwqNaS1krctjeesJD1oyfpMo
ADyd9l8D5WFSlUHNfa6p45BFzYorakTpBn/9Q/+89+qzJdgBKTsKDpSJgzR51YAJFP+yCU28zPGm
KGy0BHAL7Ow9OZ3hHb1DeFnqe7FyqzwvK7kQZfZnUFKsogG6AswwdG1pF73pqU3QkKM+jhoMPZwQ
CWdQWUaUT+46GA4OAoB3vuOVEscP1Z0JZr2lfmwV+0/37agHocz8zZycP1JXbjYty8j+LN+5JkiP
rsWF70kS3hMWnN2HtuolrSmAkF/YOG3QCf6BGpLA+eiKZM9yNgSxWtvChKCG1JncuqA2yWqv5SIR
AxVZy2YTx0+oeI4QEzuwNK9tM2r68sfQJeEiMAnyXb/5tq6lTKSvQreOD7WEqk1ntuNHvwSc998A
92rqZQSBMK2GDGz8bE4m5yh/OAP8mBcSEo+cU7VGWk0cmyKgiNLqHQGsAxWGQV9uLCh2OPmDF5FB
u1IMnE4LihPYTD5QYTi3PLiw0zOteOunvOh9DcViGi4cidmxwnezu4CZDB7r8HAJvNa4r/VKHVNV
1yzwfSabHCCR154QfsNXtxe6nUYfFuKOn0/axFybaX+c6xxp8TzddmTdcA/H8NrdWGB9176F+FK/
sf9+p4+TP3rs78pLB9BQjTdJvqS8F01KdsRPDoRJpXOR/CAawGMUoBVjE1xBovNp7gUuUJ5AWzuG
nS7lgkHM1xBmgL0S/b6yoJS9fv7TblCsqYpMwo6r/RBdfzGuw5/LaEYQQ+yfcLu8Qgs/nMUP5Kpl
DpsjUJp988NRNXz/wFizdN2gMkq0EHfvyJaH2QO7d/JyXvwKZ6WVQXuIZvVWFvFtNVb4fDdXwD/m
5JNb9BUr3fCaxTs8d8hNwdfKBt2DaWN4zuDD2qJo7RMcU5D1IbwkcVxcW2uqaqQu3if0drsTPCCB
cSdo+nfqL2IUidqXNInXSmrT9KOSbSb2QuRlux8Q6i5gXHIbP5DY26zq8AKTuHs9Yx6zH3+estE3
o2VmHK1tWfH0JPIJYayziN1/lYwb1Q1+vM5DjLJm9QX69cob7kp4JYknfIXL7Pi6GkbncRZYomK5
o/M2rQU2zzmJ0D7baAlIwm2XpKvmzxzz+6RvIjqDVvb6oETWBlcMzTxxV2zVM0SciQ==
`protect end_protected

