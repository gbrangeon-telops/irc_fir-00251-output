

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
dKfOe1Fgzj6faSFeL/IK/IGbXRIzt9OQ8DZnq2KAQwbAq1xs/txiDbhMB5jT5GTGOpfv1lX7K9mJ
mDVaIsrDmA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
cmnaZ+nYMcuVxuKDdMnuchBB9inZOxPR3/E/irYVdWCPhl0UM4JuWPFoKMQnAcsoQ3vgnwO/qltn
0x8JvlvddPokOTwabXK7+R741NBmTaawP5Y3zobRhI33jusePpwNTanCHaHjalZxzALXRseOguzG
AwGiKgpBkrzwT+frUqs=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
sUxQSwzYYe52m4+VJThnA3rSxL81p7y01A34NmBjYzEeDRUnhBCVE2EYcZxUZHf3SzWeAqe17qZn
+OUEYPsHFdXLy5QnKWkfeT6eelEedeGrqLjWta/XE+CwvggarDRC3yCpKHD1RObvSaidPkoLOQaz
Mr6i41kRIdL7xQbC4uLsdgEZKWh/fWAVQ0EsVnkKqE8EuxaCZ+UTjEptEyr1FyibFlRQuCcRV1zc
KGcqqHxwzSvE0/TqNDvaxlN4HZAny51ra9dxL1achi8jzJgZlO8wt9Agqbh7GQueaCXon2S1zoWz
ehgKeTmxlL7ytzeVDSpaRq2XKBPlYb/82fe70w==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
nlRZm6Q4mAeDfFS8oXcdcSIf6QMcM0qJWL/GpoNfKsPw7GwRrG7w5Fv9DZ3ev8dGDXi3ZhhDXcQa
Irin1hT7IkRZSupkXr6uysVtJeCdG/feYDkdTZzOR87EjbK5yer40aqraNg1lVIuObcgZ8AniYE5
0hMf7gQTkG+H4+tX0yk=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
HiHN8/USAozrVtx8xCHzL7SU/8fs0dpiHUe+Pxq1X1HHq6PWwlbojxR2di+cVlcr3m6I0F2zjyVW
WLu1kh2il765GldD+RCzgw8JhGbJOXcaDKXvV9p6bqICOBy5WCTf6gQ/vOVRu1kKDvf68tu0aJcM
5GW26Rwq/4L2jSNVHzuzVdgC87Mdq7eVgLL1qlhKwYslU6Eg0eOYTUfGfgCo2Z6Lcfi0atBesKpT
DSbchvClt7fyjz3I+qeNhclJOyfOLBdaqFIyBSFk+zxyw4U3h7toqFVwQu8Fc+NwLgyBezl0ZUBN
S4Kep7fupBYYGAqkU2vi+UvgcgkZQxj4+5jXGg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 14000)
`protect data_block
KotSLlU8AFBOyqMLP8RRvukEHVXo89Puv8q8bboqik0d3sD3sw0DzbsR6tKqc8rTt1gZkWlHNb2x
mDObj5dA3pdQpX8bw7gpMWnyEyFtc9OTddLQABgj24Kt/nG7/k8zuojcwHvusi1XyFsl/JpSUK6i
cabqvu6cWRC9mihaZr4jqqRv2b9NSOo/OS77cXKfc73GRPG5E7PbGClnn2UQeARiRpHpnesC8nCX
aoXUdAqtN3+PF81yP6EgLmfLHr3akJSE29eRwUSU5fNwaT+2SFcDV102KKbXD/DD6L38ZsyHGSqV
8OVh0wh7sQpOiUfAe/mlDcsKFQftGGN7fIU5vOFL6vK0vqL8oE+VSqI8yY/hskBtXTt6D+o5s+Fj
eUFDzMUvExP6BInlMR5Ul2K2sRplzxPWerIbGgvi3UsJF66Wwil5PT9akLZBkCGGRZQNLcdaQG+8
DGzdvkpHr+rw8N4pVUT4GPhnKszjEfGRufIupg0ZfPLxXJrEtsqQh/GDVlQ4tpvGHiMnvBuLm5gy
9dWpv8RBf7jhsaXbJeHTJpOOacLBgbjC5dd4ufHYJeXQpqjM/tETKKl9umQnJA3h2Gvc8o0wfq/d
CV1sL2PbjPkSebnQO93fbJjrliwlw89/+843xmTF1U45uCk2F7wtvP0V+828ChUdJ1uDxXFoEIoW
3qYjYQ2c8JETuMUdgfLXZ5Wfg5kaglkywaxYEylUCkJmKu11sZ/XBRjKytxRBClJdcq0qmBx2tZG
Mj1ZvAhpqia/eaca24DFeBshGr0SXvTG2lMLUEqmbaiTkkjLvNhIGvsV/yZZAdzXq/i+677Wi2Jj
GZPiCRvjwNhBjsGtSeiyaDM17xzMKNeBsOIimJOEPRj0CI5p08GgBT+L5wm35HIEHWvRN22QU9En
W9zm8XKpxKn4eZjwmG1F4x3cO2hlDlqaIznZ39v66v+bP/2oUZKIzJros6hdz8YGsgdHb+t3ipmp
y8M3lexmaKa6CEKCnKAROMc7GZdiWG0ONZP+7rzdpccMzu4lN7NunlSQOkXkfhMGNuhDHCl+ONy5
Cnz6lo1KLyf6LYlvsLY85BYufceHukA4q8YqL7/xQl/7oKkkS+diBG0BIDfBPzOl1EpDHouio+p5
ZCYy0DgjZMScHmHtKohxmC/GDDNt/zO7Du8msgBHkH7Ws5nYM53MnrRCVY27/OC4vO425nRjjujT
bdPzTC5GdL1HmYGFXJci7Km04OdwyM6ylaVaqlNvKXHlA4P1x5Rwcl4ru1kHeHzLOncT2NYkxnXw
+X570wgD+dhnBezbmj5iO/ND/0qvyttzp3MNjWP/g+I00HqQF4gQ8iF4oibN6C/wsANX0uWXDTqG
Y3z4y7jrH3y8SPLe0VIMuInP/qiwuNlOiBMhnqAv4nnrQl4WPvnlMQ5oIqib5SUdy6Vz5L19yoG+
EgOWZ0No4MDqyae4SqO2FjF7fVjB7lQvVQhZMbofDZG7zsrv5KzpivqbtYAn20N04gFOW+9RjGBJ
vUDOp2bm9S9rnsRb4pkiSTO5E1GLhDhToBCspCDwzofWSbKvYQOGAASFPNDI8NPLHw5WTyMJK6mA
QzRMf5U42epQA8hiPKVhm9e+GXvJwT06mgXFOPe45EWXFAgdhIZTqqxofGw2mjnYPr4O6o/fUnJF
rn9BXi+ffephtaTuOfrjuoFAOmXqJkZ2IrFdvgTEBJMpp+PDKctYsDazLhk7qG8TkXI87ebFrJWG
OqzE+fRCdCeMdDC8u/7QcW9Faz7iBy+na+fy3+EgpF2PYqlkomKi8m4WgGxxW2cdHZNapuKciQWX
Jub9WcS0SLDo8apEay1PcKwYZbRvPOAZJvg4RIcjplfL80OOMHv3hnXczwgO9zIpBi4WuroiFz/6
TVFRNtGA7fA6Zl5jftzuYuys7rBk8Be+osJ72DIkaUFkwrLh/LbLu/7bg6JCal6XDXdhhcmAQl6k
SGmYdILH7LQpQVtEfiFdwHHnxr5f2qUFf7vB8x8rBSb9VlIU0QHMOzW+H2C0Aq2JzInPcSRYIPDJ
BGwakjtxDvuh7UXBBPph4qqO0NjZ+1Z2Sko2JPIhpBr5bFBEAbfTWJe98mdY/+p4X1P+AKDubvZo
cPgJ//Xj1cGqd1hr4URsPrUDZt9X8jjTmReeIB2iTPRM+KnGgY+YUBxy2pf0laY1/YYHtnRLnix+
HulyBvUmR20T3lq6nXCtQIrbzmoXhJdyG8dO0nNn59N8NUo331Z4b16ZUJ5ut94UWwapDm9K+QCz
VfSKSGBcTa/beKJ8c5m3QWVTcpgM2XOvQCHurHvcVkTvrMRIa9LLIkQLCAqqLLV6v3Vdvi487n62
DUfhwFfmUF7Co4ax1Jaf0tAn0PsMvmOqMBJMuUgDPNR9+i5iwewmCXQfsK88MQ2b41gxJ2K+5S13
uvQWSndFirMuZl+yw1lBuDlkJBt//GHOGtTLA/wgkvHNopgdhRXL+oN+LPcenUeRuPl6MkueDflg
LEcLY50fjf4D0VEh6lGC4PbrYXn2RMPWg1lFlaxxOtDoZeaZrkUo2P7SLUlzDAKmzGSzOVlIFSCi
ssqBYs0liTD09Gl7xKG0O1mwkM5v1+iEdYF4ybQ3hKcDc9R9tjfEGr+7QHVNAmmnJuuDeSETxHJQ
YAS2+pZoMdZI+/dqYu89l3DMtIX+SsNV0EEmMNH7juACJRJMaJCw6LIuwWozP7slVfI8eZOETxVj
fW21sEH7/brp8ryjlsLO5YCS+JLIBFDHmgL4PDDsSTUunYajGNUwyA6JdU6Kd9P12a6DV7KCFrih
lm4JIVWhzmnUo4BVycfZ3UtCxYiz+WVIs5/Tl2gu7VrDnZ2L4osu083uz/eQxl0gO92obTjndZbx
FpSpcqEK/wGACKkJ8zFE3stBXy/uFsO8ZTJ+MBmHg63oksFp4jDRvhpbxsjaauqTx5QNYL+tUGIr
SpTTVIfx5ZqYAP4vUDnwa5cwcGEczayQ/ipVLmw2UFPhgiJYjOzgYeZLvhNZ3Pkq8seEojawc1I0
fkTfzSlxAkgIS6r88qFMxyJls8UmP2dQFUr5fhGnMtEfc5ClV9gtpI5pL8gGDum4nMK9cas410XC
Xwp1oHwUxionPZyK9xp70PThJRpLXp/vBL+KooILGHIBN8ups5A8CPm6Ms/bzd9U7egkRBNVptUB
fXnKsNkfUJdpy2bVpkvWQjNUaxHP16akiMPv67lWWCMjVoRHP3KEnUYyfWpNeli4am3OsJBvJ6AT
8OChHfz0KrmeHrVDCFdHaiAvg/O/+e7hlaxlB7BHwZZ2bLIH8+OPB8rE9OWX/kByUsbFsE27NOGA
QQ3uUnDh9RZ0ejxw0gsU1bzAgY+HzlLYA9uCJpn7bgkMJqL5CpxiYi3jmI/rn+KYPp6Y8gFqTC+3
DdtFk07M9seM8hRav3btVXxo+3POP2F8tXeWvt/iSIY9L0IVFkeSYpuA2wDy/OtKts//AvkCnH89
NKu743TaakM7WocpUmVFOXiBSNZJr1fr2+t7B+/dYjX4upCthpFM5vCeI2q1sk/ZA1Ad1RQX9FGA
nLHP4m+S6PWOosODyp4zVwizP1RUOV/spAbgQOsoUFI2BgyVOPBzysT7uQmEnhG4vbnyZyoR/l30
Yl3tEKJ/jnW87bDFb1bVQ7bK0qWbBt5mTzO4ZKPcMvUeHZnmFO3SYUrSo6a0UOm1hAWD3UBmIq1R
L7oPRWIiUrPisqz3bzxpdFRFersZDAJLfmnqa5HTbmoVQrdGksGoMLP9a8C2aTD7P4WjEAIMt3HN
8Z+UC0fy+/RfSZluYL5OgcYI69MMSvg+bmdJ1X6WkhXet83n8BHL6aPB2GVEmCN9WfuqtSMsc3V4
UCGgt9MIGTUPQv5EbUmIFNdBgKXMRkK2DCyIROgBIB5XtGAaNlj5xbOjehzJbDE7M3izhBwHlxpC
l7NwunTHsxP+nKXYCBtqftATr3QF1Nc4WCwx6wuEX/ngwKRLXCjO4oQOVYjvoOJHIh8xonfR13iC
3QYfZ+Yc5spqjC4hG39fxXUVVUoJNo27hZfyK8e3vQ1Vf6H6OCT7TuBrNtPfpavS5zZTpu5EFIvt
2GDleL0U1Un7ghtwc52WVkVGeOwOEPoSnH+XyRShLfHdUGyHppKs7JXHB4MGmFCxtjo0eHlivAkP
xNl0hRaQ1G5a5+szr3AlTJlhitIPTHFTkwYUn5EvGxiPfuUh6l7n2Rh9txX1KjRUbf9eUjvvN14c
ujD1Aa2EUqOw7hOrXvPi82W+PePb4bvYKv7EAxNFCMjC2Oy6ZyymaZOFO5N1Jy9eT0/13C0ZMnnC
64nx8mb7xpitVJSFaluoIHXE8izTPpUbuBX4Q3j04n2selhi2w0VNlDgBwjL9CQwZiG7GibkXBwd
z40HyBAsHKJGGr0D1VHsFU7xctlMbnzwf1+hGadRUPGa1kBgwnJa4vCeVhzdN/kaGIs/LvuBF7Ev
WEtMYGYM5mUzUVUCgFD/KjZ28ZZzIdTIMKHDLlzo8+imOXDKwmXcQpcs1TpqQaCSRwXbu2OQ04he
WIOZXkR4ygZPU6pfuHottu0mGzDJp1exASDtm7sj31ydJbkrLgtZM81dVljOubYxruq30xi0TtxN
p5NtSMLmUsu4QyX3iSIUKl+jNvYJV6BqymEjBHnv2mUx2H2hp17wIuRtq7WCD8L8yoXFymgNI5UX
2/97vDt8lnl3gnRUHteGJk3C6jFfdnShveQHSGT755THpTfcJeIbsm5UsqSzLPKGzmkDdfppHF5o
nulC8dICsZq9Ao6tvppqCXkPkv8IrNGHE+J8V6kpYqhxmqUfWi0UW/7G3b072Us+ej76f6i77Pnv
M3oW+mHl8FDmMSnXGpKuYicKQlHRWhJ24mMper58YnycFsKosS2YBm4GdDV9MlRPiyFK6n3+YsEf
l4etD/o/alLrm3XOY7xgnn6hL8fmmAnFWpDPb35lGxG0vjHbxBsHNRUxYS3Rm7qgV10Lf2OgwqEd
cTSRrPGGTuqI2miN7qLQsj1ZCTMwFYzpwLk0veE2OIaO56Al4T54HOadeJuKMSExGrMwpiYqfDnC
lxFGBfVd3Y66N7BjZIspDlTn7e4ykGBBMW0yjBLs5RlAyXyOX+xCV/QJQGx2SlaDszNiiuodoNCT
FidbUJATbQ0p8KfhCqqmCoUOJHYOeSqVVxJZSN2SBnOJMy6B6rbGbpogMYFYihodY+JKRZIngxWO
Got6MFMTmqpe/IkGpacYQ33skdlfSiT+xil28KPujAwqeSIDAYvsIkH/eILnSgN0mFfUbbf0aPJv
DA10FIb0FG5wa5uPp23DenEaF4LqeNPkVdN7H+0Jc+P9SVtvh3t6r/e3YgAPP5jxeONSsuVNH4ZX
DAIo2xpkEEMWud+wFucXmiR8SGBDfTfpJi3owRLlrUjOZeeG944rGS7b1e9xjScAW3/8TnpOAg1O
zyzBgRFJxzevhHUfXs8Fc1JVIf197mzK7/+ET3SIoHCqHexdYcqSDtY2VOO38fbGRQmEeMwQichG
B9DQwIWWYwi9tZNi+VdUhZbpPvdk3OmB1NrCqvdwaX2Zqr8LkcP7hZjAeN8/SS6ZXDvbbX94oki6
djdLUcOPeTGUGQywtY3j3vMHMXUxCF30yGG9WoAY+P6M7PF7Pqr0PkFUPXyK7kTS4Uh6p2+jGe4H
GHCTMuL0t8oxT8xtPNCRa2bRIo9XwosP0HMDDjLfDrwuljHQwxgRhzyIU/PgMDX7wMeosbdsXKYM
2kTjZHkEcfN3Fwbi6+f660fPoyVBT8krrBBzfxoCynUVc4DHdurqsjG7qtjqETv0nRCOWEQ+xw1t
Hl8+PQKl9Otlx1s7zdreFRyOqPeRov1N1L5gHzfWjCZkPSCoyhsadIWuO41WRkW3tzZO0lCio2HT
7PcET3EpDilUWTBSP+4xLPcWseQk40Yqfpog3oe5Vog+FuinGW/e3jjVI918W8F4LWzdGo5wd0ww
ZQn6Uf9pkc1jMeD+LKZ/F9QhaVLoIAi0TuuGV3gelkPX1bRRq6nVv5ibxn7c4dK7Ofu7YLur0WNR
85CED4fmc8GW1QcTfvZOrIcF7Qoq9s9DOBUVSg/w9Fa3Ay4KyM7FDexjF0IUjoRwyi9/TNuvdfiz
uWBHw+7AAs90MM41sDuypY4Lao35JtuGE066hzRKfKW9zrKcqxE4WJM6d3HZVbGS0fFQLmqQONq1
iiOTW+0BaE3HInBsOiQBF0x0ZldYc5IFGwOx6BmwultZVZIk7IEBmJW5NdB5Ubo+Xa979Ilnomb9
ScWVWp6C7SQqciBeuysdskVhozWc1RXjSHkh8LlNMyHRw38B9HQFjH8URUC9DzWi07PagwQQWc1q
OdUh6GuW9fCtc4vqUqX/diwAMulC5JpT9cprql8IhrGGHDF0qA3sna8ALou/6xSetw+B3FOT9eyh
UNqvTYNRxFQhnSkbj6kYTj2rj6zJZ6o0XASebnVIO8Q/m2bmVJ1hCzcnf8uWFvDURwt12kPKirtD
y68HfTkRS757biLkOovY+8iNNWdVC0anp8c/fjlB6SnPWeCfq9sNt/TQ+T9vMRVMLkZ5qrXB4NES
vwFcKBRs0XdfCuPTgaTt8IiuxDLTFERqZ8IXGW58rRNwbLOLY5M8tDNiwL2sy//jGQv7i4k/KTiU
RNsgUUOIacz9vg8m8Q2qWRbDWvDdwzObbfA1J8YmICCe/2a2nN8UJwGMprFiEyjTdHaI/0B8RD0F
qnkLmtMPNOyoWPDBFg/ZePG04WGEtvRdC6ZzpBhtgVmQzOjUEqHPPZH8xzO9tu9YhCUuKPV/QmSW
7F0QfhdZ4S7IfrpET3G10wt6X1NSV+pwoAAHcP0gzzjNuu74zootXxgkvVhcGSKzQkRThXpnt+Tv
JFemvypCBiO0gEykMcH4XZMNkIZd7pmcDO2tOOYaCSeWoS5n1yQrFxEMOYLUPdkbsJHDLch2z7Qt
MsPwDROyJ9dr/rrUXjGrkL4qzKks7mGKKOTpS6wEf8/JXemUloEER2bH2s1BW40yRWaOEOdD/m1f
mZRqFwndPXL8wBxQr/KcKeawCqa32szwLqeYAEON5eQTcgaZ32rwAipF0h/xSTi8Egjsp7gWAIWa
MDp0Ijek7pt7VuxobOPhVILW7tQoLrkjuYiEDwXG51Ym3GGRh3q1UVlwTAxbLwm0b7bedcNqj+45
Lv0Li9hebK9dKgZjkOEZBW1mrVHUWPTekESOKP7ieT/COVxs2EOJ8nEKbhXZP5bwhi5lzuNPcTF9
YKWEFWMy4w5HhI+s1LuhLfDokQGt7MW1aplB9pC8P/2O7GOzGoJolTpkI6JcBt1eEmy/txalsffW
m9FbuaIackDSRhmtN2/HY+Voqkx+XF/c0oPRmSa0CZ8oLnno5vLAJV1rxgwC4xRv1vs/slDN+leN
wA5LPNFz7AKxoubwzuPrTyiZcBvC6cHqv6OzH5FBRy1X8FGJLyayCXGB7NvbDNErhjTKrfKnXc4z
bK03z69jMCRzG2zKvjqorcpWDTf4sjZZAkSa4LfmpFBDTEkgsirSfWsJ5pU84DO9uNKE+9YQloik
kcrJ6Ce7uD4Aee7sBCVvOa2XtMLDzurmoJg/i0L9Cxga22nHEcO8pTxLuRcJwTmD/oxeOZaPqCp8
NNpAp5FlhsbDE7FoTOIJip0CrNm6U3leHGlR1HT7Ki2O6nRg6bemc1wGnSiVV+ydiPiwHmd7L8ho
ozsPbDXT0CYwre9G7NNJwOgkzUeDQrN/vEXDjCiyoAPSw+bNMU4YffXcXjcZJxRIk99Mc0W/ppGF
QcVp9BhZvgLaxQbaj/kG3rAVmW8mirRJFz0qjKPxxRKI4GZNTK2EnMdN67UOdehV7xsWD9gnSA1R
oqU9uInO7QwdyH36Z77sEFDtRWBmLGKoTCvdew5Z+RfdGZadl5UWpT8/WhWiLOAHhm1hfYDSK5oa
eC8xsrLNtPep8cX7ufDSEKY70y35ISshgxLH+xTbpgmIst/6Hb4YUbTR70yuvtqNJxA0lEb8clhE
DbHz1WSaloRksYPobnu9FCgt726/BWR4fpCKMKG9hJGU+KXj1uwHoAfp8udbogHVNWNOxd8dpGK+
oAYYfq0S8qLniebhO5+7nkIVpNodpYlS+en3+1JtDKuTI1X5l4NdZbkGra1OwHUW7FaEflME/ye8
VWLfk1CPQRftRtFBbussgZYaOqnthRvk1ASksVwJ4ssgngK+pzOD7+TIqKYEMzAEYCUzTSKcwAub
rVZC8AntDxZTG+zdO+2/Crfw9+gU8zjZGNPRtb7fruwTFFH9eePEOSqMM6ZMy+UDyPUj1Ee6Euir
2W9r4kGYYvr1PWlixNLPqYrr47UzhjZpn2zy0pSEzbKtPyOei461lSlnrPn0kxgqeeRC4b4xIMgd
1qv/GqgapmICzuGSs/X5bQYhsyQj1Au4QadZ7/OILOYivA7NFQp81CjATs+cFgplyWQsdcLC6GFi
TgIk7l30I55fUYlO0rGdgcpV90mLwT6nCOfMXKmh4gY8FFML6AEkDk9h7xLRJ9z8ySSi/qZlnp7W
qWcUN8iiHAnLDZhu4SRGI/eJRCr8f8Is+BLU8qWKJTs3dMk3xj6WOqSAl/jMuz5WAboqzxOyjzT7
kKH4S771auA6pFpIsfA+vjbeOHpN0egnW6MdGoDdjo2NZ1kXAmbxZEHAfeTq3Gs3zacOC4hIOzSm
jcPFBoJGB+IoXPhCJBoHASR7v69xeHobhyxvLWW8nPhQ6kZSNvRCEAkPF2E8TmxftbQ3e/oxm/Co
FTLcBEZ7NmjdD0LBADFlUJHrbf4kzgCNWpv4Rm+hkKsdrCWOI/0MRDCMcIt1LIrBV6Dj32kC+ym3
XhfbEEPDYLDz+77y1jBE3WgBAb7D3Lz9iv+nOWR9jjzK0IfPb4Hx3MQviBLvPzXASGgAfxPjUu/Z
hwEh59RpKBjLF2itpYkzgRpDmYKW0CDEJS/gG+4EDRVPKPLhPQDeL4siQ7mz6dlduVHRIzB0eqsg
lIn7UL2wet4ckHkYVJ5x4tturFJt1EAlAWS/DphRVyVq7uLu7KM3eVBDR2BkMLSTUvp8A+4RSxUc
3RmpD1AjAmvLewVjsIW3lSxH5DzN5GcCZstTkRInzi08K2H4x6ZEb1ctBMsNjkxohnJZpF0gCssH
OGlBVA3+5+s5XJyAuEpcs/WkOYrWXFEM2c7lEecPbYl14nTSP59XG0GqdMoGJmL+zmoFldng+wUT
c6TkCz6ygvcAay1FuFPjbMXfB23s/ftHg/2Tv6NELtBsM7yqEInV5vm9Ux1oRAquHzldLTwLHhJg
9a6N4cC/kMEgnZxSAJoK6zdFnnRJnTKxZeoAZqwkKIeqLINyzzsFL8jj6jpsHqrLMmrsVkbXIHmU
Ah7XsurNXN6d7fff4mgxzBYkTp+z7LITI5yRaP3f/I6HkWGN5+9uILB9eM2FwLMT9QcA0oUg2Wox
RK789kFeJJNv+WCp2BSSZwgOUocVbeJUD5Bd46p+/ukcJlOczdobBoT5zLraMfETCZFKpWXm9jsN
UltyPI1xF0iQYzzcYmOGNFLnaUdlP4rY4Ri3Trgfs1TLJDawtizYbGJFQ5/8OGRm/lTGn9xnhPcw
oxtHbd4sNGE5GKO9itPbI7DNyVomgbpReOKjFxOhBbHZYEPnsI9+Egf1cQCO29PSj9h7+SfeLff5
oAFOscy/D/ZUD8Z8PM8rY9F46RZb6z0fUhl4Bwco7+TIT5pYWqq8q9eKaBqnpjWrrLNUOFc7C89K
webcGzn0TrrviOmziMkt1qMr7Yn8+o0nzGCv+2WrbyvMDShkPHsqhXs1epsQACss1WMWmpE/TG7t
T1M48wY/C01a+lsXEc+vOhp8vnneoxAtlukKszAdO3IJg7q5XqcnholHkCgmIzoNgLNILz5NWOIp
Dp5p3FOMr7zvC+KQcKorIcCHO/hztiir+vfu/cxvS/K+PmNUlw8w6vjnS4jsUBdrkELywq0mNVVA
IwNKCGpt7eShzVcNAN6a3gMoJkhwa8Q/4fpcFd7re2HSq1XO45Rb+V9vyy5FDD7dUyG75cLV3st8
1BT+c2wNYi8qKCcHHa5SBh6H2t8Mjo/VmZR/MrdWY6yzcpxPRTB9hU9kpPCe27Z12rUVq2EOZTX3
phf5wM0UmGT8gEo8b7OKsUKAkXwd1ljZ3aW0FeET7D49LazS5CjCDQTM4XdzW0J+17Hp29KIZOic
RlY8QAMcUCQhPJtyFRBQRZzvZ1ShJ/oc14UbRIpbGpD00fLdEUKhmXqYjVpi817JSv4AYAfV2ThZ
R6c0xUJ/UztCIXje4WFpAMPUfvZfrxZi14SbwyUUSlVS4B6KOnQhDGCXgDoMgEutmJACqkhd53q3
xSp8+UK7R6ylSvlT+s+SI54AQipkXptBzNm0pgMFLlXXsGDqoUqpRvFxATJKtnIJl8U0XBY/wu0u
mX6xBaLFofLFLDpaxChF3+wh9/B69RegC43c0P2IZCk+kRng5vs6ikp1SZYAgYb2nNTT/M9V+Ty+
W4XLYwCsEi1KP97IJRtJQMu3O9Qns9aLBcw7PjOBEr4Yroi1h63bBoMm2I9GL0ghfYwtVGByT0ZR
hDaxhL8NS2KqeKb75WTHnfVE72f1PjEIvZxW25eF9vMDyEE6rw0Lxi9HcuJQca7KcDGzc8u+psRw
JKdrmjqImIEdwVOvIoLJX5EHkrJrMkJ5S8MU6njv90Fapk38+KxuYxl1fA/nfmo1FlUPZ1+g5yVa
9ep6XYs9koU/GmFvn13RITz6PAQ/fDceYxV9WimJpiyyhpSNj0l061qSXftD0AhHxIDSIFhNrqHT
ukyAlu2gMzhI12msKGlRcoKipwTdZLdJbXLEHYZoGHSWZPvGj/sQifJAWBPvZ7Z0zK9IsZ/I16sc
FyK/TsnMPzQ/fpv1FexhgOXqZQfYkTorizr3kpT5iUAInjhyjxwzzcTPkXpJduYkZjcEAkbuDG2l
CxNIZIj4x07toOczVpYCCtNbAfzHFr5bM5cqBwdCorp7ZbEgiyW8v/bXG1yGwRbIDFckPZAG75e+
+TMZ/iVGJgLJZfFNxeuVQeJoZedjiiSg32l/2sRb6AvT397BUCNZ1vGJ6jEjvlUk02kMuA9IaE71
oMcFsOoDwUyOZ5T6/P0/GTRgrNB2/rntSwEEbUt3MAxgLy8pHfcedeJccKtVWoAUNKuFdUh32cwJ
CFMvq2Mk73GMwdj6++xJqBFxmvwa+vrSzuRwyL5dZmn8NUDrx3kpb8U/bWvC919sA+Vp7MJEYDEa
rxggl79b5afhaHh9WCLHChlFkZRrT/dz+/S0z8hYRUhMtnqYH4SJpB+cVIBlaznOxpP9Tsw2MN2x
oTfuxYFQm6cCvCXpfN7FhFVh7jPZ7ZT+C++iX2oFlA2iVOEoknYTdJEnmYj4N6X3Yo9MHuK27wKV
6+dw0Yfv0GoqcLMSErY7llJduoCWkEOzMHUJorGQlOFkVr/bsp9vdB8axlThVbAbJLb6BdMDmkeV
S0+OD2p/spPjpq5JBuuAoXp237hALJjpqny41cfCDoyRaLQTX2kdwqHgQXMXGgX3cXryBhfDl41N
oVn+yc5cAuVjw3OCOZED60oZMIeXKzn9BMF5sbrcBOYvf3mh461aNkamUFSZi/xOyEgtilHh4Ocw
KmBUAGvZYUhOjvLYXk+nGmfUhikdty3cZPTa6Y5IsYs3UVK5PiIpwrIgEZjE09TD5GTfqtfocpW9
ZwvAYdjzb8GUrIR97Qh6HMzuugFAVKBWrI7eXwYSH5eN2OEe4D4Xpo7IlrwjHH9Vi/v3uGoy/Kxb
8jY7b/aDV9SIxu+6hqsyZ8sEup8hu8PSz0ZtpiZmPkBO2lxo+8TxAe0DUPxP3C0RWGxTCaaBJ2+Y
Se2EdDnGkB19gceWPzoRxO4tgOG5uNsVOfeCID1+XlcJzx24341a/z8VZIF4SgvAGnxWzTDukb++
yGlXWb51nhYWt/MLVR/tgNSAL/Bzd46U2gIAG+zvLLusRjl1H1zYsIcHdag6WMD0qtbY4d+S7pjM
P4hrR6SrZTsVJXTtgO/v7tyvzJUuoNXojUkww5owXDRGzQDdU6EvHN8ARVkCP/2B80u0x3XjnCG2
mzFbdkRvcKAzi+hhDFHX8diEz8uEjrw25aUxylmtNmBmZ0YWP7FxNRlEO9ixK2dFf5koIDaCbUfU
Vo292rT0aj5ZuU0r4kEU28GtecdJF/vWPkjkfl+udhag5+lmUiAr+z28FRY/212ZJZrkiZfZlpj2
Km8qGsrzoRwcAJH6Kgtces+njpRIc/43XN6GNh6i9ibyd8x/A2X5KqQrYLnoVs3rfTDFeG9zbm+R
Kccp2BiXtEYUWt9iFDhxGFdjYOrlkLo2aTeXfZdrUhHhNo89VE/9JSyg5c0VX1/EVkDdC3tvQbYu
lIkfcLXc4HdiBcrL/zGENt0N/F88EuKV58P7eGlTry5fb662vnESXM23DWGntKWg+wL+GG3F0ZKN
dE27aF7llrriWGsI3MPNRLkXJ6TZ3J8opu5W/DXRT+RE84kWci8Kupl1+LVW9fwAmbPcfF+fT4ay
f25stORyQqp/UjwLYZ4bvlIY2OSGtI/TmDQGm2940phzXolIHZ0mEPoyreY5I/kvZ0xkUPv9CCr5
vY2P3PB4qA17ayz5s1qQp79b1nS5dtx67MWzY4xOLtL8ZLYRzaBkHXd+5PZDJl6FdIuuQuizr+oX
yyDiaqqfZGoecEND28xfXYxABHDHtAfkd37WP4WGglFyfXtw3NVU8vfVWlcu0x03ZF8e4kNYG/yQ
0ojAe1j2gf6fN4fdznLD5hf1+Po8xLkPZdo1N7fbekYnP1UMlbFyBA37AM0TChbcor5l3O/6wJeD
BK+BYNCtvhVXjg0GWpDHhqcRClglHrVvnF4guRXvMAJo2RxNZm0UyYX7m8wxONbHITaLFdgI3lDk
/BW0lEgmVbtqhdvKGHHvtHkC8UwnhXDGQrvwnjlOi1kG5rAHHYRlhuZLCWlSISPxtakhnTBsW1Wn
bS/w6NPlEKvdiaNRAMNplpoF6aRR0TufYMSCV2YVQBS79Ss/Piwab5Tkd0bj7s8EcU+SVTp2AEYZ
yOt0tmyAtD0mw//oIpB9y5Vhh2vN0QSU9BHo6ZBsdsQ/mmnK68qr/c4qf6gIslebW2tTRQ4ctLMA
E83jFluSd5/1CHtUep3gzdSGJx2XnRXNwpG0dHlNQiN2WL/DYRTi5+/yu7E4MzyZxENNSs+BNzJr
zRQN/jlQPP/SWD1p7VGA34ZXE99Lz4XOh7HiQO/cBe/1XR0pN+oaHIHlmBbX4umb8PsFPfc2CGQo
AXk4vZ19EW7r/E8Gw8yIejtFwJpQtfs7BAX4cGIazC2DGq3rKazizadR16EQp/YO+L/UqbKYZtV3
uH1Au230BSnz4InPpFlR1DWzyL5PTeLtJbGYL33PGOTfknHEGYJzue2KmjMIqHaiwfLNxuaWPsjD
VfRHTxz/gZ7yIQsfYjw96DXYp9er4xZqw42LvST1ps5GLEwXiIZtb2Xm9B3XHSx8kGyQh+m807MF
mvO771NTdPU+kSGExHvSaj2RtFbZhSYGReWmtr3Y+pTEvdIKkMbcpSC4/GLmUEXvtsySeaMA9xop
oAfPfrTD/tSCJSnJhQBx7q9lIoMh5/t4IbzWGTGuiuw3QzIvVq9TcML6Kb0AT2geN0RRhvQRvAaE
WCmVl2ZMITqhO50bOlSkJTG+RKJHkr6yAExLf62VoBjDMSRM844m6z4n7HiTIwnPmKvhRZhqnwa5
NgzgO1mMgF+vtsllnf5OTjnieooItsnjd5GWAaSTQHT6fJJlX535qs4Ce8gwva86+oDGn4Knekaw
mYMLKYdmj8aNn0TBi+jWQPEB1aGYvPdzTf/MbIb6QV9pR31pYoq6BiHSUfT3MT5QnRWGMZI5QWmH
ZpxzHa/2EKf910DWngOpdcsRlQcMvtskv/33iAU1ZfyXAuzkvjE20hJJYYo/ZFc3K6IvdpZNITNU
u5w3WKObDeqBvgcqlbWYu+PuTiqLi9OZYwW29DX+5FaAtD2MlzHBcU8+UHGNxTZnNouIfSLNNtcg
lROFEROnpBXYPrKlLjmebzcRGb/4R9bSZMOcNdfZ7rBJfJwiq/JZ9hO9goMXVsbTIP1SLKVFNIvm
88/lie2448f8LWmGQyXUdFwLihuxGjpCS1yZ+KW6ZXgA3V3OrL9UE3AgnXbYpXL6ohNrkpyKdT9W
+KNptWqWUJH4R3iV+LLKiimFlFCMWd0ZuqLryD251ljtGFDw0AijS8VngpSPdGZwrRt6shXTN5M4
U5Luo/5KWqzarrT3qMGDp06Zi72bjCCs2xCJKswwY5PhzKbHonQcYBGhMzCk41xn65sD5jUwTuwZ
EaFsT0xRCopPCc+hK7Ss5ZiD6ziUl6yyTiPiYal6N6c/7gZsIaiMzLlk4TgIGMu4Ggagd1hzlfdV
KxTFmBaSv+XjPDTdyUXqkS9FY9UyQXUMmtXLMeP22Xv43i2DuXt4C1E7XaMfbFxyvgoh7ECQP3r2
5FnjCtVNGkmkIeABB7iK8h1TTdfoe4gl2BHSsHKlvM8eR8nGCU6mn+7nLzcsRp33a+MIeCXz7jq0
AJIul29PWftlBYyS5uziZYXi9cdZxs5z5BzECjyoIuMi2Wh4DBbJQ46UymH/gRBM4CEHH6TXdS0K
sD9kiqb3uDuah248OMs4Y0L5h/dxtd7AsutLJ7KfF6kJBc6qprq3tvu9+Et7WmNJHYv1owCmSdpl
kNf+K4WXLLIyu5mBIEe8YZ5MUrUBR6HT+yrLczGMGBS2aUrAsi6zXCUxyGErUsrAgSpoYttOWZiD
r+KP2xMkHZX/+V1NzGyDVqtM7FyMkbkPFJ4DakiHjJLKsR3EH2Hzdq0LxoMqZvlEW+dxsmuh2KK8
/UtDvNwSirNGzkVOtzsl0uBGWWM1ygPbSGLRW2RyG3cjHy6Xlq3KlCmemMUbn+iMLGLtWf6o+pjB
C333ZGM0AW01VzP7rAGN9tLrr4zmke3Xal+UEH+g1Vkh7w9n71lReluSi4zFIrZXB50b73ZhPWyx
VJ7V9ihpVgavkaLQG//qr5M3Ruf34O+w/8XqgUeDtzcgLZ90ZNM/3FBp2ltZgvT9htQjl+yufhFr
E/sVQR7hEpdLwpEUsaP4bS8aOUQNP7RT1OborJNZIV56A50/JiK34PGzTUN+1DilTyVDCKGux3D2
zkDTMleXIpqMQKBk8fNkem2SvpD58zutGZLaVB9+Cy4JrXsa+m0sdCZ4f/aLoqCuBHQTi0aO+/mp
w9rTRNF/X+fgDHBj3jQvQRq/zagPzfxXbQpYBPs/rYRRE8MGXcY/eBzdosYdXoNStgXp32tfu1Pz
tE9r4JivIAB5UWRWE0QBkbD4CF42khk27RIzmqestPeXpBgrurJNbhODdKMTjPaTRFmcAL2ZT4mH
on39qS83CO6Ue2xkL1ZsHmQh3R/UbCJh0EG+ZmM5PSufOJBfrZhT2hAIRwaCif0ZaaAD2jFoKjTJ
Y7uWuKgZoilZuaKxz9Dj8vwPUlFxIRQdrT1KwrOf9RE3eOhEaTkKE6CwxeIPV/XDRCZjyrRwuvCa
OuSfks5Cl7MgXjTDxDez8OQMU5az8sr+Vw/Oj6fr0ViAMDGQPMQmTST7nJGW/tftIjWDRwhdiWZN
Q4fCQ8SGgPEXzMfp4tCaDNsTet3dpJRv4DgIm/s6j6kpzOGPLuOr1TK9QPN9MHJ1TTAqW6+Q0ShA
3KJGNUnH0/aa62kHqDCDJ5lMaSMcV4flx1ShUeFmRdSC0KC0mTF1AiMzHye3blE2F+XCpJKUKmFg
Iuyj2DyxPV1+9aBrAVIHNfK6Xv1y4sQ+YdzF+MX4Gho1PzteJ3UK+RBdmunUloGy3HWtsG1yjUQy
0bssjytGXCm3mAtEfDpS43vNc4nAiKUQgz8J2xtbfjErX5fHx7tSddOv1YEL99pZinE8q0hHvsKZ
BKEg5TIJSWHxmV2zQt5TMMV1OIqzCiiL0+mKWWIl1AhOjfymdcETJA07ZWBeoT4kPOyM+x5XSzGc
Sj40fCcq8EhZnm3iMRR8dNAcpwyIqcIoWzKZqK61zi0+Zo2pudwTZazXPnIKW4EW6NozSh1ER7xm
zwON+JUND0R+9KEoWHuPrv6Ub93iqy2rynX6A7/6K9dOEKQWGdbgNV4TwMzkY2PsL5DtPz0jV8R1
r2TQgFy20WYr65ORZ0dPATN93sfr+s03q+7FHnGQM6S4UNI9y/kdXzW1gF1pmnHTejXUnAwRSwqF
rJdRaprulxwubxVCZ7uXjx9amqY+pW30xV4gEElz17llouWaYRbo6vYIme/iwMnLLcCZL989rmQ/
If3ChhDMG1MWt/4wGLofEHg9icmQnVN8STOePTz1F2EiONM4D96fthyxslIY+Ox9Ix6bZtXnN7DC
tVyZ75LqmzNm1tyqRileaIAaD4TrKxmcwAgx2fmm61uM+zCALGXLURVw0+ipT8Kwha0AjmRIocLF
ctq1S1E+FLa3+uyvGsFSMFyFfBxkPkDAqRqpMjJ5L2ay81yB1DLboVNHLQ68Yi97VVE6WTLKBFMO
po+GIPzNzCrO9SFjG9M9/XgHUi/tWb0N1AHDaLM5hkCChOTknOuUD4vrvGJGjV34foL/FwLw1O6n
8lxCsAto5ItyLUCBRw49NplAyunydvdrosZLblgAaBFmDzlMGL95LKuejBofNO4po0ISixvPCIYf
uWD4KERd2lzmkmRSXnbnAIbKjIqaxKjMM6fwAlLjJ+gKvZwzA2g80XX51hpY279QxO0UJH+NQKRh
EXpVK2wMpQ+KzyWcbGoL2jtkEExgPGdBj5dIqu1gxzY0GoXiBMQshqDBba5jPyt9DhAaiuOqYdWx
Bwp0kYYh65blsaKuCRb6OF/YT/HbknN90NOl9EiKIdoqQuZVzrxFbwuMqN88B9CXCHTc9CRyztJh
ERPBpVJE+Dy9cJQur19Vco/gG8GwurJgkpPXrJzXhPQXs9cq7aqaMJxFGAylEtigINa4Knsolj+I
PWZ5Tmzt8zLBrZp1rqntnzAh5m14QdfNyoj2rBwMthPdF+chTTzG/uHg3j6c7zGfr7Xn/FqOYF0p
2bTBc/Q9zn1Xw1S/0bg+6FBfmLk96h5YZD15YJd1HMfCho44PKBovXsJ1hZSEXqiUbz0N2GJdX4D
0d3tihpkYhBHGXrr37mBT8/GKaF1cqx31OiPS4+2N2XRc/qfLrMOKUblssGKO7DGwjgvfsoq7Hln
QM+0uwhaydWLC0dVfuIrkRaltU9xEaOjpKbx+Y264j5FnEdoPqcBpnrj2ZShizM0P+Bu1sJqZy60
cwZJt9W82crKMgkMiGZ7fEt7tsnctpZTA9MpjrhlyifPEBDcaCf2+MQiFrVnswlWWz+LiGw2wPNv
1Ee73eMyPFbMXpllSKeayMm2EhnFNyYyy7nTCBiCAF8/NQLemHwJ33bJtgRsLO8jCKWZjcQ0EjKl
58Vckfm6ZXDG0hojGBZRyO4dNVGxFPneiH8X+I3hawxnXCWZkAHtvc96nD3zrUpQJLKFX9JUPN/l
an62teNJl+tSYVJo1r+PUfmBvyxcnIPGw6pwL8C424YPzgHR45SyXJS6cmGqX5vG+wRNjpS8N+JZ
U568jj2EO5M8dWw55fmvpLTHdCx7R4zEd/EbHDQ2uqLyGZvxtto9WHjGSi0+6/yK9qkbnA3RcAoY
8eZhIptybuLKjK/+9bakPiQnwSQsmSGDSSrR53hddRwGWy65JURekCST8QdLvYCiK3WdL4fKKZky
3/a+wlQpZam1Ww58dPh+abRVk9ZJvDcGX15tJP5xmf9XMjp1Ry0VrGNJZ49NDO6r+HVcEtxtzAQM
9z9VgwCDcurWTTe2iXwE5Ufho4+u4P7ZJ1a7tB2Ya9XquuCTQBcyfJAlGOyo3dAN+XiW7+8eMFaK
GJlLB1OXgj/KxjNvAlIh7JtU14PnxPuCC1bZwEZR8q4tFj5f1w6Sn7yesoRser3MqN1rHILS8Wgq
v+reu/1j5UTMhno6uAcDtgzIMV3wpI0ZjFbidurpi6Qu5uAc4WmxZkTAw8jZWMDqS4+Y1krBbiLt
onLhyEahDryCaNntNcM3un4/oIw58ShUmzEalamlNHZxrY5c4835SXWJHP1cxglFFEF9cCVN9dcE
z+YssR0lTtKWFeJPaYuSahbEdJxi+qyQBp8IDPPi2pjxCGWXUtp7gbt4oQ3vIv3uac/ScdcbNV/t
XfdtHNqv86x0MhD6ItcqQn1l3NNhDZewo8WG6GVp2TSX1Yk42Wcgi2vq4wBAHeGxYleNszX2EOSX
fPibAse+fC8vF0QMonGFTR9dHnm6UNtMGiM2WUqJTe/fcMtaXqxWBZvOo67Ckp4dPvsYtJf7vcY7
S7ITsdS0Z9c7qEAnUsX6T2bKyiq8UbYRCK7YjfMLc8a9hUm+okT9E2cCKgnROWl84OQnPRS9KkSs
JJQdYgahE9/ODOyyPeZ4t9e3fge280n/1uLHpZaCOdx5Ql8UdopxoYitDbUA2vrDGHIHZR4J/Ip1
+UVXWxBYlP8PspgK8OWWLeRQjxx0P9D+2h2Vub9NIAfE5xg=
`protect end_protected

