

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Pb7E+qNVEP4sE5d3TkwQJMYKTR/FjAPrexB6qdDJcLdscPV5w27UvNCqw/kg86JgS2hNrfoEvTNF
uJ9eNTpy4Q==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Egq1eCtVuCp02bpffloqFi7UMw6fphk3UOZCcejhe9NQNeC0Z0b1+S1NY8yEfAVY74l4oz8pZ1vA
hbrAzplanZae/BDY57rCQ6UjD8G9keaOwYv6mG13f+m77D7Y1nVpXOE4Uujw3cZ1QgwXR1H4YfYp
ysjb+lxmo0pqYRikRIQ=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
KJqrZ5TKkbTlecBRrKRCsxKhAd1omWJvIin7DNafgTE5a5N2or7GsTSawdWWjYWHESLBvStvRGQE
jVUeK8m63dYVJN98fa8T9iAHTDt9yiBRki/VqfvAejvDOEI+l8row+LhhHMvCd29xmkCeQKiq4Qt
hsdsz+jNufnCYY4Y1CVO/4preMZeG5Ow85vRd/341CoWEOBji8o4pk0XyIttBBgjBzWO8JyhLpza
R+Z8LgFoZ5OTfgpyTJ4SjYRWp9IHP2HL9TShNo3PmM36nFNBvQSLoEjLgk4+rUr657++ugJH31/C
Y/QScvwJcbqMK15awb6twj42y2gxJSFzAPzSGg==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
KxmYEF19quU2lnDIx1hLVbiBV1iU7MlwBSbpQKNAVv6HLtZNpIjv2UPtz6sPs9Xac0T26s1Kjo2c
fAw+uaSeKdgWE1BMMV8ya3nIO40+wJlyaPYGp3qW9dt6kM+FZZl/3MCpgIMx24FXg4CPHrHNKu54
/3DZJ7o9x/QjyM8WSeM=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
n4InNydlMoO1IH7Kq1VdB5tuRxM6d++erhleefbfKU7rQGdfSjRtqcQ+h67LKfA/jQJYdDdZMjd3
Jp84+E2i9v4ovZP9CPOifgPGXKRtOz0XzimXarAjLF+OJp3As1WqoTrPJI1DspdbqtDWx5caLezn
hcZVfRSFpZUoLc9H0HW6DXtxAWvJT8e4ntjJYO6koEzzHlZPpMhXvbbH/rbArm4iRGWLOVN205Pq
oJcFHv1n/e24XGuCRksBqssUXd+D0UgsxKn8Hy5kQi4Q8xdFEXxEOVBI7ivvG+HKnJFOOr+UNhLY
+rNFOKSwlDtT8tPfpzjKS5GdaTuv7j2GVoF5Tw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 21824)
`protect data_block
AhnuBR0FRskpylgH1NnFAiZHjs3y0rVigpT9DaXaamgEVX2EwtGhJJ1gFkNHTCWw8PS1MgYksA/T
kxpV/Rn+HUlForvm3hyUsILYS2MrgKFJ3sAXuczmwucsoXTFVCYxRwoOHSG9TxZ0yDjjaNBjYgjm
uAmCKAATxuXs4Rr4dhKr9qjpLTPQD9dhQ3/PxOVFZx+TIjjXqJHV/8jB3Q1COcofGUWgzukRDHol
AzqtAvpSLHkRK1ItETWQCWHpyOvm2J/Kpuk4+oUbWB6dGUq3GlD4DPTzqlJ3VHhzYWW0kqSDeeWi
jLMpSFVrwe/d1VHpwC7jK5M73fqQgArn7DXlDlmaFQUJeQO+bfak+mDF4CDKYa4Cs0ILsDM3Q40N
uoo1gVL60PY3hA3pIPbGB6DvrxXYGj2pqGh7BTKzfmW4B45cPB9q2NU1HekhAOSsmwagfF01Z7HZ
GxBCd8D51wxXl5Sn78qXbnAX+yGCvBVjzfADoF28NXeh6CHsjt++rFmzLktHAQK60yGi/uCPPcMr
Dr1KneFv1LtfW0QCuPw8FijtQhPi48KMKql92v0zSlpGcBcP3v6ticS+IIZCPeyEM+H9lOtj92F0
nDShLDbN45vDHc1CbdtzeTEe4QnLdRNxgH8igco61SjEA8fmPW56OhVGAq8sBql0G6vfhqcYNCel
VEKxkyjkuUZZpN/N9mt/KTRqpgMVs7oZbaoCX/lmB2SmkN1yCVbjCxR17qBh9zwFgoxv9DC+nDRC
b33CZ/5hOuMGMIia1ylBFpcdGV4xuSTHdBUEDKK1/vc5ybsP/9QdNOOwVbbByOvs55X7BOyjvZV8
mDcBHSe1E+DOagtT0SreZWdoBxLiYsG0f04OcLJhVcf7bHI01H1CRvFNNj5t/YKrKDM6UWCvvMjQ
Jzy8E/6WwQnDMQxTOUOHTP2XCCu1WYjpY9uGPh6PhqmlUKVSfBSk0tL09ASo2g0RDOzE/98C3drf
IYAmNC1jRLmJJX9tn7UsmmYb5z2jXAsYUNUAEgaqNWoqgQevXawkwr8oRBKS0IsUNPONZGvpkcbD
NWLZ2BMRwM1wcSB+sLEi6V7piUdEOmwSgOcyr3rumOUJcFBlVmDyaAlEKw4JX4TOxtsoZHqlLeHs
IbSBz1VnDV2lJ6RgAaWql2fyagpFiA4iYkR2w3OBJST5uBiAE2DF0Brh7uKaj9L6I7BzNBHrp1/Z
puDJNr8SRGMjq9HGIUv9K9w6kqIY4LTG+kA50bk5tQRTrQu4FSKbpylJekQDMPsW0i1w4Za0x/BU
BU0dkZBe+JYC1/8w+g7k/KQmHVHGvz9Jf8qsDgX3vub4zkD9wjoRJ5N0oL4u5Dbek7WpuHaM4Aa3
T8r+yYtkyao+BHscb33maAuDzpyd8MKrWKxY03Pu9JeMm7FTaJ9Cbp1jF8yqKVceN70spYDsQGCh
tzn437xf1sEr8Uz9AAkB4N0JnIWZ6CfEIZccoX2z16waI2LJcgErAo3A7+CJus7tgzBUhFD6DaoK
o0Q2B9t0GpIBQWrw4zH52QMYMBjBY1+Yf1p4OZnScObkTbyi9EL0CWI4HP25Mvn7Ap51QmoCbdM9
8Jni869KoSf3rbEkYWPJInWMl0Bph78ZIYy9sid8t18bZDWPHQ9eQGaNygaj+92tpnktxhJJ7YdK
M+0Jmo/s9sJH3B+sGkGurBgk/1WkUqCy/dPliPaQghA6d9sKAJerP0a9anv3qY7GePH96i+wMXMG
IKuU5aWGqHU+MoI+5633T1jVZ6Vfyw9RpYGuRuR7wV8LdBcpXj9cwlQVMx7LjnTp7QIY57vmbIkf
nuIpjiAPPqo5I0akxmzirZYr5iDQQzGpHR0ea3Ngnpf/JkY65xuXaYyAyMZzbBHpC25R5WmSyA33
13zokCuDCEWg1p4mgeCM7LcxcYim4cRossicI2CTom462JCsttMhJH2Oj7KPzt2sU3pNE2nSus0m
IsUbyZfVdUoOJR0Bn3iVU4+DVeGKRYu28hbHOZEGIqp7GPzZPJ/JxOMgw8WGv+QLKP3nCfzJEVDN
AIFRpwXgdiWxjAwWXnL6PZ1lO6dFvLQCACJQgBZ5R41Ky0p2h5z9Us2v4TPWwRAgQJYbbj4GWt6z
yJ758BwmlurfamBE77ztfeJRG0ffDZ65dh6akO+WsAcQ62PRviNfQIu6yyRr3mmeXH6CC0jcLLXJ
Dv0alMKGLLSBx4+g+LD8+0A5ulEDbZhJ1pjJ216mAFsUJAG/1m/8C7jQnaEjWkbTGXSxK4WMiACM
tSCrpLuNAyfGIEsRMIpZ3ESQXUsmuvLMNtl64c44GYOTJiM44Ubz509VBKRphezkV4SQbmiVuOtd
frBXw9uO2EaBCbMezgRKTiQ6ynSsHnLjpnc42EW5RBE0zNmHxcOr1LT+GvdGsCfz8bi1owEKuax8
ta7cfdSPo5f9Tw+G29h/pY+lBJVdS/3ss4XqT+DFASWyc+X1AdlNfS2qlGF3mF//0EKXPxyOSsE8
X1JFpN7T6dw37MB2hT4oE/2O6g2Jbs14bQNxmlE+24drvyEr6W5tj3YVsdKmKlazBCaxGYRczFCi
yx+hZDvPMsaj3FbvMpyizHaUpyAI6k8RHn8B75q4vAQR6Dw1LS7hZ7E/TMCqMdVrEit6DJlkLTuH
HhWnnubVcmXtW/piLCsB92qtiemT2Znq6wUzjSWKxi/6KcdGsAcAVUsEXpzue2qAZYfNXj5FzbKT
GZnZ3BJpFGLkg7LJGpW0r39Y7j5tOzHHtoPssp9kQFrLWYdglRoq+f0hN5Zppm/QozaIJ+55S0uh
tYz6WUTYT6A6zb8YLyBhc2GGOeAbbIuZZ27CExBO199wegeBvd6/+p1EsqwmjGjyhzJiZqxQ+yBT
2nsavFaaMBMT46B1/HGTtNzcjnaWzXaOJGoHpa49/4GJnuek+O8prYNYREOHCO3P106NzABtgwlf
2ZYMcnC+O7xnwDFgHro2elIvhS512YdCRIxXj6zAZaiEZ0H67ADADlnjvGEWCCa9vLJ5uw/R10J9
crHUJb1QDX0nQEVWTPsztVVqe2DILY71PncOf4b6yA065SI1eb4koxpAshHaz2ot6oSuo3a1G4IC
NcHCoXGja/b9CBzfrGsSolBhXd7Be2/l5UI9UdvtIlFGCWUg8nSa+ibpwlSKvHD0OsPYToEsjYmf
tHkd60o99DLH/GugUvqCRtka7yrBPLu94oGtBzFXSViR5Uqkdf8e5LgSzRnF5nodu9rmb+Wxf5xy
C+io10CdJouODchRzZ91lzEmOWiuyNaTqSrSwph7TXF51//GneunCuWXUzOX6K+bKw5lavv6wWYX
se+zHy/XAfnaA7TTj4d9GPK2wXQlTOdFtb3DVrHVUqvUYuP8AOd1KQOmMxJpg0grBNjzF3Td5p0Q
CZ1QcevRe2Xh7GUcV/FYS6cXIIyRc7LW9Wh98gm3Qf9wGWOnbiOEd4ePwTlB7JyqAiZR7w9TcWoS
NQwD2k3KefMH0dSWENMb0mCnynIHGn12Si3KwnBhVHCtzYRh9/CCNu91fpGXJSL5bTqjtEdONRHs
OUOJIdMOVupH/6jRF4ldgbBbnv+G4/M0A1oePC7eQzkcvGkcPlxn/rlrMfLXeJZDqMrsITq4d+h/
NEaKM6OMcW+QtftIDwUzV1/ZInHomcVd6jH7ySd3UT5ETNALw/PNe5dt4VA6HYzjauVAgbozr3Eb
5roFrNavwytoDZjE7mpEGmWGzibv4fr/5dFv7Jye01+3K0jJ4EwhmLvHIg5JyiSDdsXca6wn7Fdp
6LL+dtMEjtopfL31KNYKrkCc13f19IpWDXAEZRmYvSEtWzKQF0ZjHd7dGT6kv+q34FBFxms6dCAG
noE6g3Voiqa/Ag4+3xURxPszAVOLritRMdSu/av8fyIHNZVPV6ZTlK7GgyGafLkOav4qwZSKlnYa
UbimxUtcpJ5lIPbosdvecEYA/FP+NONMlet4jrnZ+XRvJqXSP6n9ykbav/Zr2MbC7RZpWu/+ZLRf
tx4l1LhT21+d1zTIrnZxXb7tCmEmzAwRdSWLBsai6g9C7GpLzZX/p/jXslzqhmp671VjFLDVUUcx
az2qYWehogS/BHdIu0JmbzLppab7Arjf5PKCj3Z/50EWALacqokhpPFCSBaBVBbS3+N5gmN/OGIK
0Cq0nObKhd8mvzZ+W/edlnrjYwEbA6I+KF32v2yzn9wn4O8vATIuohnexRyfaP0MUDW2kU5OmKHI
Tt0/WLBNhytqoNKCpRflWQG1B7e6kv4tczDTjeQ7EqFZttANFlO3cHew8iNukyI12PNntLK5LUPS
02Z8df6GnXfsZefmikdAtuZ5v+CLlWF9KxxxRT2gdOMvguQIxShyzLZiQ0JkSvIbdpNX82+4pjOn
rjkKD2vZiaU6Kv/O+rWnOWvpX335L/mTDKIYP5iy8YoYfDKzMz1HHEmxYSneLk0CudZaq1wjRVet
NTuekthr/4OnCjkN6NIxVyRO6/3+ae3F2hFlGnQxBu0pAtLODH1iyTc4uEVyo609UasS9x0Rb2yc
ohb1yXcYCLdihTeZqlxrLcL2oFroF6upw9SuP+kt8RNBsRkFu0JeZe9+a5U7YE9FYuEWt4AhvMoF
DsIHnuV0zNy5wpFIHy7hWRjhnEs1qW2B8r5QCpDW8KtzvwJQyro5JZwpHEjNm0pjwpekBBmr1CWj
H5ts0Fitn3/r/3FUN42EbDV3k8eFYGmvVQQi92n3/L/CUxgTYGL0x1JIaSK0xinFyTt4MLv2FBkQ
s2RY/r2kajy3LX2kuFEch4qoUDQiuYeJyBEW0uVW7XHDjnC8YA5e8rnysv+djIiz/TSMGjkBMEcf
5Jv4NpuEQ4BejV2Ach/OOG4Yod4qiTCOyXzffDDlOxNkIapQ+4KWHmNRhTZcziEt/56aQMCrK8xZ
1Y0PJnFlqt2Tuv8Vmp6HVgPy37nbA7mkh1w96gHawfhx2pUZTj4JCKO4TkoPCGrGtnIna2pPN9bV
p7vupMakVn+daTsfuEGZnXAg7w7sv1dIJjRs4fNlI9zalD2xqpjz/22AYOiHJPT7/Rox6bsXikh1
P9pYB/HAGCheQw1x9jHBWzt9ZYol5bHehTOxj9b/MpEA8gkGOyRHBVkE+zl7Wi7QdUEJXRRqSNcL
LJucJBkwbnc7wzw+Y0J3emscJpisSiCjf2GAuKRqMOdQRejorCQ5GvwsS1kYSjlzv47M/0zl7eN/
8Yk/PbLHQXOK7QeB3U53+CftMoOo8aH5KlyxowQ7r+FBQhlxShcv8o3EOUDTRIBT53YBQW+mYfdb
0JYORyAeDCf/w4siKByvPP7xPiUSEr02WR4yKSIFPOq+WTcge20tNGT0rSxPYKtyA2zuJ/5j+RXn
9g8a+5ijXcqZC4mAg6PUaBnHkC7BluTXBJuACwM/le12axHz6m2je3MlsMBD3aVU8F4Bk9TCya/J
eKpucwD7asQaUiS0twWIIarMxJEmT7+6SSBAaxuHS3LSVN3xw3hbzNJtzEE3Pif71F3gHeRuUj/+
ECVKrCmYEWE66wfr4jpxjuEdmLl4PYtHGR5hiO8Z8wd+TMMltLdv2OZYo+0zrYxe4sSTDagQQHal
3H+r5AgUFE9y1NZtJ7GxWsO3KPdit3c7UROAVZtoXrZRPNcwy7ElxoM95QsE7Q4HgFVj9wvv0DMh
eEsdDGSpCHVBHTfVpZDrTj5U0eZBvW+cK+CBYQRHdf8U9tczJwRS3yrQJX+OwJAaZJv/qkxGv/2a
WON5pj/CiFR9uOgJ78d+ESBnk0BoHb1nvnlMpbMr09fQ8GhmNhX8NLf/IJ1SaCYehAy40U/eEuGQ
wQ+UnPqOP1wV7Wy1mq8vywcbM9lbsd3xm8g05O61DjQ3ZClDk73szBBskypauZnJ2OZAT1KVETTa
+Yi5WjYYZgCNlg08QnGQoZeox6RsMP8gkexYGvyHpsGa6eg+3hWum2eS1SFzp1KTVSHkAD2DDK6/
7eDlzweu5VmxbZZeTuI/T6LG4EQSXIt/sWDYz88FdfgywVHH+MxYCGQxB3I3VBoUNytvpov1g608
V/b4AYAgDnVj/euOcNtJhf93BLYVNhndlGlSZu9bAfpVmLIuzqVoAUwsllNN8MezJrvZYJm3hxYh
AQVlHQiiT4UaFhwiqtnPyyyA4UxXmu9uZvSJF8cAlCC6IEWc/yyNeSeiEGUSykT8eJu6nynQAj7h
XvMemBBC3cYyRD+bN0lRlgPgKPkOrBbnlfdHZJB0j6gwmGrIwSukmrLKfzzrv5sJfjwJQOwj67eL
dEdhAE5MqfllavtjuZGE/G5mVw/3+Zj7rSlwz8wEDLJjcnp/Yf7G1bXT6YDaXQDgWiorBeyZWRPZ
WQ/kEs7KYFiA9xYwqQF1W6IiGPZ0FO/SATMUstUe4pL/LRDGC1d4MxSvT1PoJc+cv8Zn8PYko8jZ
UMHNQ7bwLYRFJzfsVv/XIjDMmav2lt66j+4ORjPQTzX6PHBfH72kLEB/u48K/c+y0DmSDTNQxiOl
VHVEKKmxO2ZUdOOEF5X4M9u9JoVc7Mt6CCds0YSoZiedDc/YwcDsXvbtEw6hBDEwg6bcGypuHjcq
DHtry4LtKAOV35OE1v1ky8b7iVBSMH50tWmugOVsUUIM5lP9Jp2n+X3F2J2cKynzNNVJNfTb3Tiw
NwU49Ml6WAApPpAZ+moKItgIdgDfFbTxWT/ciQA8pUrFQaC62w2sUsUtBrv+ie74NmlGuJh1igXR
tKoj4dJlCYMhCV31D05mNGcDNFgq4U0+qJWBVHd5/++EhV/y7QSPUy+PQ795vmb8J/2O6JLe6ahn
7VTV3UEEM9fOVWyd6TF1tEdQZzG7cH652myn/hGb0fp+0zTtte5xwrfEl7tC+1ov8EOQAsf3Opce
DFNuqQk8AqCJDECOCfPsvHigJsPC0CqUeOE2x6dOfIYybw/EqLS96mDt2k/NqYHZbMq39geCzCdx
KpNPPK9o1ck2QgQw/25AcIyVA+WglmyfSavftrkfMT8I1RvkrsZxAb+TZyuiKAt1X5yJI9oMuVqz
gncqOyIHD/gspVo8kXZH1yVAwisorUmC9pzSgLZ5h36DDuYRc8kaeVjXdp+mAYrnH9l19CHSrsA8
jxSyNyxh4kKweAXkO2NZB3tnNzI2IA0uY+Nv+H1e8qxm5GIAPCXgXZigILva4Ceo6MsHbLZkcEA+
ipgf+z6+NMOGswI9rbEBnfCbqmSKlnrCpoLNFJ9uT4GUIMhg3OtPA9f0cNKQoI8PuHc6kGnsWQ2H
rPX3uIIZR0G1+UNDWvYxywdw7Xc04PEde1EuZIpKWxOifS+iUCKrH1bbL9TJx719v0eZ/yoAHoIC
i5KXfqnRZQXAIRqPrE0M5qVhypiGj6VU9p/Az0OVAAKHaZtXF2EnbPtRn8Nhr6E9j34La8vVISj/
88jcLNa8POZjto+YZJkXfMWnj/U2Cn6as/YZk7VUiXz+ileyAHmvcViTppXg2cAUEghDrpSGmZIA
crtK2sqK8V7U1FDlZK10RB1A+lmSrv+07z+5qCF2WUu9BQA+bCXq0He5JvVNeT9cx64YNQxEcYxW
AtGdUk0SaKoiDYDOHoD/AnUaS/GrpFH3zGC2IUqEZSCd/uyRSlmzilZJV0FysaTY5zI9PKRdx4s2
RqIZku26Ib5bmCrgWcmvEiTFeZbjWiqpAHbdek4odik43YbWOVqx1UKVI0DHo17HgPI3bfr4vzWj
HJS+9JoUia1EW4AXIoEiG5AdPEhCcTV8fDN14u8KpyWM454pJOD1FJYsHsyc1+U/4DDF6sm2sxYT
2jZJ+ERi929/Ltn1IzFyEY1mkxLYzzn7tM2tU3MOQMkaeMBmT7AoLDIXmI3VM9lqnC739LPcLrlu
hSTeBPbgqj5Dx7ahH1abBJIeS8OMbyhfTxRGdU80huSv8KQVSYjYvyNcz0HDMAYYJHI20RJC7Zcv
w42DniJgDJo033YhMnx4g16hbLnerMMZNFNxy8yAiZ/uABZ6wfEBw5PUsZgRiaIcDZXt1pUV1ia9
KHnYWBFkIme+0VBfl4lE39CoHziiSKu5OtKn2AT9rIfBGtKwuyVPhWxXZNceOYF0wcXR/28GWBDH
ktLiS2ecgAMeXfVsDc7I7qQf225RBY94fg3g/BqXmqPwC7NHxrm7E749rFe7q6mAwl70mP5qG+Yp
rpSBOxIA3abHtefg42G2BnmYmEOvFtB6hZaEHlYs+KLaPQPC0HhmWj+08wn6oyNN9fJFLcN+UL1T
8v/HXt7viptCA9NWo549uYzQEzHPY40GzPVrEBg3BozdNwE2ESwKv2h8SHkwor3SMk7BdlG0cZG9
VvlB70G0IIwNp7cP6ZEjuvihqW8c9rfqZ+VlE7XYsrXXa9zztkSs1hi/V/A60S53Y51P2zBDAPbd
l32SrqGMNtpi/IYP5kGnFdslzobARhJ3l95OobQXfmRYa3mZrpSSa/Q2OOheR1g2Y5U1WoA5kRMy
kwxm7RfeizjgyoytUeVxnpzlfbehMxgr23YnBxhPnyARBg94853sByqbXTrEwF03ywGn98CxlEvh
bRxB8puVQAs5t9KYcl7g5aRIIng5y/m+u80ePbM1wMHZ1fcKCmvbnYnK5oHVSpzhsV2Guw2DNYiq
ZDSA5xxeoc9YYdiZKhIuL81cVKZtuy7DgZVL+eUgA+Az+XyxpP6HL3JZVlGzlHNYImVcTGfY48ec
wcetoIS5SI1CdY9M79feYDO3v9UI9PKqkwE2xxiLA4FizmtPUCtcv7pV5shvn+SuirYC5kPO315O
cvIgUK9gxcMX7R9jiWcwmcb2qYG4Oq/+jA7SvnLpn3tycyocG9/ucBozmSlef1aOcvRFLu26LeMp
84+0EDAQMNAzeI5y79UkpI5WqiuBTQjc9TFNdGv9PeMHBfZhROyrYXqLjVAGlpbeUchB4KlGVvgw
4RK/0gojgOfxC1rAP9ETZsQ9QRnfD49PUDYIYNFhDVgzR7xv99EEdzZ7kMuCbXgUyoC33ZtVygow
/YfhNSc61LhTfL+XZzM/PmCNmA3bgODAmzuMLCLRSyg7nkWJD0LZwg0RGFWwz5WzrALePchPVWtx
uR3MD16MtdRNG0aN0XuHyx3LbctBqgyfa/HGSe2CnD2qvQd0sVydGhc8GYbxNxlUFOiCbDdfNePM
vGKtKrgmnCXC4zGS4QPSZX5edRSv/wLVDlN+WU5WCBGuxIpHldeMifmVJefsl36rOwSO2hkI6t9L
G31bklUrG15GY/j+z1oDGkzflnKGbC4JqyrO2XpoaWmcfxlekfOeOrDENY9hZ+038RTb8D5xvmf3
vJFjuxut6BO/c6Fz6EpqfAFwEqq+jeHnMn8wL7eJ4H6Ve7Re4/wFQ7Sn5CE64SfGFrYIhtJ0EPN0
m0Zva/JNZR/9KeZoKK+MlmCFUoIu4EEQ0FC5hlkJV+zun/+nmachBG9ckFbL1dNV/XMyb6i6k3pi
aDpZDIh+rnXMsjT98XxZt0WoOm5JEcYNst/cLh+0nIaQP5DLmkr0C0rKgIatQvwNN9BDXLhtLEse
5ZYB6yqqOmMO+dtd+H4NAePajiNAiJ9cBjZAlmx/T59TQ+tx6IbzUfo40JAk3ufHnMMK081/0kGS
vAwhMTTI/n4mv0C96WBq+NYEfTGfFUdH7NVAXPDTXEr7A1Wt4nx6q+vcLSzAbiZkalcY2HDls8jO
LVVpZ+Ht8TQkC+i6e3JIRv6MSztQyRunJegNrZ7mLpM750x72OR2khXS1IFUVMLp+qJJ0SRDFi/a
gHYBLRpOhapJx4MPXu4odSaoY7d0abRhGs6DOf41Ph0S4pGzwTvM4Ckv8gcIvKgeBaXEWahE1mzT
zdnTuvI5ySkFdEhQH684vLU/3YPjQS3UT9hEWPt3/6+V9UPO5rIw2eIv1PsdiTUqmYPqwNJy8142
XWdUfJZnK0Om2RX1IFsvGcw78ImUALpV6FGpsEf49KeLsfJ2WRrpAwmuJybNtTVGFXIkMcGlVDR+
PP5t2pd6CGbf+0Rt7FRcF5+GqRsRSBSQqKUIhvHx/GVHMPhexX0FqQ4ODFLkCxOOiTWO46gBgabl
Xfz1O8ezlwtgzpMoheocjmmre9rzlqK9Vq2oBSJUR6t6kRQyXVCYa1Gmz+dgI9Ym0tzPAoIDiQvC
XhV/J73mOWWr/o9pRRHsSc8miCfYdiWsQymZIl5q/U8SKeIU9uTy8LD31ERPTJ8n0p2itWBx7zSY
0Q8LiUFETIwFM4/qZ6a41bzn+O9mByxl4qY8Wo3ZPY4sguDx6kRBz3ocudVkDwDiokN8n5SpQh9l
uvgAyWDW9r8KWpN/SzpKYP0Vzpj7CuNFn2+FpbbPWnb1SgTDK4SeVGv7xmMrv8TC81GsZAoEHCJH
bgU+QsEI2QYxwIV28UYQ87PegZcPk402uQU8ymuPNDq2pjY+E3W06KI1AazegiSI7SueKApS7pxS
/qa3aPCQ35+Z3TDdEHOc3xtWfYCKSZd11i59KYpOYwep6AMX7eMGpcJmk+c9VMdU4wWGxHN+YVUX
EM5GIJ2dmzE4YaWDC5Lhw6+sEEr4bbYYVWxDRkhb4sdsdDv6RKAfcoxPUTzcRiYKFk2la7fKmG3k
UhtTHchRw9VGYUZhukOYoWXWRBSyy9HTP72fh/yCCIUj54VovPYVFEsd4juzhQq7zsLWgkC11pYE
zQKfFCAlhnXYl7hfb9NGWNSq68nktWvuILyV62PBWEedqRZOyQDFD6LloqNyE3E126kMS8aopEw6
PHImUNHB8c4W7eqYl64IrP9MydoYxXbdBxDKuohbesKPssxlLf3S6O5iDEr1leWoHTayERw5E4oM
hEvsVfvbbA3+hJeo30+9KQlUqdnKtRNUSTRP3OZgvkeaa4wnp1ZuuzHtWkefprc5YyrDtg0gsCSG
RK0Md3UZ2YxMHe8SZhDbt/51orxphZpxHYAJ/gLhj7e49MwNj/eYjnW5lKO983bCyA40Z6QT1Iui
JJAZPEIQ8opABaChGZRGiZ1BmaUskD+YUUNbDGtvWiMaW/HzPPmvJkTNAhAKSz+t711EFzTRVoex
ZepcoNO79pwgzyj8Cfuj7UGUOmm9ZOLbqCdLaWelQyQCTHR/1uviR1YosEOrPhMqpx93c1AwOcWP
USTICGRCbqbquYG86xpp3qrzxs2g6/4C6SPwJfEkmDWEdS7DwFJHIbLdO7GFvXEphYO0mwXMInZc
cr2RXGT3fKEzIUnz8R0Go5SRhQLS5sceRAlh8wafQsLvvhe6v1A9xrCz3V422qhJmhtKOvC0KTRe
UfqMVol8XBjMA7FFjsIn/nrS7cYYY7dfPPW1btwGDGcxK9PBAe2z2EnvUDwxToLEmWFDLNnipStl
HzNXk6E/iwrbvdXYAlhl5yuVIzgxRNzLrVQXH0AcKAlsbm2EY/ZxQKKuvOLAtmhYTm8F/+XckgUp
rIu0JQiO4A7AV/Pp8C42+q5wrc6FO/686p8MVz8LOvmj92SnPpdcwmqxSORBI2k25Q3T/WIJqDjG
duaNu+cmpQKA4n/Z9zlaiThGybJy3xyzwhv95+Litmh5Th4XJ5HjOM2vfHrIIjc7wgwMLIQQiQro
sUY3+LeqqhIstLYhqt3S0bc0YZjM8baOVHMeJjpqeOYPi5lCLESJKA0wPVU6fNHlozJPPK/21EOf
BLwEVXL+M8fwi+wR50YX+bi2NGZiz42dFA9TiPe9FjNPeLcLkHyyjuPyi1MwyYtmscVPZhIb/ACH
gTn/ClZalzrlQNrHL1A7rJZUfzRFw7+1QASE2QU0b+NJ0j+u0SF4UBQO1jmA9BMExplb/MIo/9Rg
UxApinTFZ6b6HfZ4p5vSLoPJ9kxGqdo7PV9h5P/FOojoRQmzS8z8k0mkIPfv01m+Fw38p58crEHv
cSoOfI2hUpJcNZj0MuipHCf25eWMnElHG79nitLB0yW5N1rhWkjhBiUF56ZQN3vH2eSe5KqfCWcZ
GJucC/RNRf0M9yXOGkDiRFIKNXEgz6/e5B84Su9Y3RSN33VE7A/zbWGmT7y0/z1evqmdodSi8mpi
NxzaliXzU69vUXQ/tqfS9z0Z/saig849821w4Pve/595HESo4dr0UuMOlTEQ5bV94hXzm4SBIUsq
gbtKVSj2Fv6eEPnt9r6bNXr1Fos9IOuM+6p8JoZaAPlMSX/E1fk/+6isnbS3qitxv+DgUauR6hr+
ogfvK2KutxfyqY7YL1DbqGU8iyceBj+oO4ZimtMSbESlwcZpUv3QIQbTVVxFQHqPqFUZCGvqNwVN
yUmSf7lUcYAPk+cDn5B6ycG5PhTUO4nbmoKV9SsYdiAc5dKaHYw5PsBJvmIJeeGeVlpW36Rb/k/2
ufE7m8d2cBvTloPRNyHtQ+4+ZLyVyJn5zO7oJn2TCJ1RXyqXZV/ktjtBZTYg/Ky4V7Pho1tjqC5s
VCS4wLhPt/kY2DOkS5VcUKL5kRnUzy6ZhoQWa1CnS8/KT9Po8TCX3pD2jj08rEftD+vJRJg/dVW5
tEuA9DJg3cEphw5LJ5944F34SeBS2xmtVbRyak0pjT9VUGNbdQXED7GLEtXotCBfCZWl3Uyb/tKF
KlVAQbZOPut9gEM9TGpzv3ftJZ9YfWbYZHObEMngwGfdzseMLvImCWNpygx6VCtOERhJdgU9/w8V
MskjzhrGPwnT+sxZl2kl7agFuqLoJGY5AxDu/qgjSgXTn0CDAEwX0xuDmmRckzmd5fJWOahrJZ5o
t1P642XZuufN3a+ykdaZDYW/+OqkgBn7Qb7lMbNmUvS8E0YtX8ORaRftbpZ/j/rUGyCtLvcrbkHg
yuSNx067LbqVk8snM0Gkt5T3+udXTGo87LTJ/jwU+ewz8ah73y34meW+rCj9fzp7J2f5zJXO5jgv
odJoyXDD1Q+eEGLGd6RWCCWj/LlA75FzYYqMa5fm5H4hqtVtpi+/sR4S4BLR9MQknBBzpsmaFja5
L+K0QceRKvDCzwDWTWcaaT9uRklnkx5s6bPOr77nMD2+0Hx0EkBlUeDL7Cyl4l8OkeKmd4aoeQgT
DeVkN5fEah/K01fu73dKS4MUJvnfKzASqE7+/xebqPBw/vYZXsOHhRpd+oh1vwwAEVebjclLNor9
0MIXa6PMPQTfxK3hoxDS0G/2hfAIDPcdNrpbFPEKJEtERApAc3cH20F50U4EEJZvIghVOleinIBS
BsAowX1uK5IvfXhX9rZIE2KislgKNKUZFLrlT41nA81CzP55J2AgiQz/OmdF9fEYm45ZwM4yMM3V
v6kFkPPKZHGeAngnHv1Uzk+9682ld+RyM69fwMeBEHPJsA2/JxgiFF3jNqePoZUxiq0jZboSKcde
h4DN4ptHWxIFbcY/a98cKjxTbrWaj1QnQ8Wz9XYnVwI80Bl5XCJk464LPsr4hdFrtto5GMQ0CarJ
gr/AaXBMHRiBqOwrpQsnWaXgj9jVZvrSOFgQhHOWkBZkDJoq7EMIZVwfyktt8pyF7z/Sogz+c+iu
hiWZ+5wSVqrmmJl5wJoC8HyOebjBt8+XTgiHyXwMP152p0KZybWID+N5/hfUxHoArJzuov2/Imwq
Dtf2lpAIKTMOwSZUuyvEiZXs0pwLonO4BIR+tdJIGRpT/0LSQW1L0E03sCwCeeqU8wzNcnqjZe8u
mP32Fgtoq+HPKLW61fDbcJyTWYkToSDQreyL8xGsr8MOTwEbX+InwCPxy2ftzLPu1QJxiypnocf/
HbzUq+O4N/qQT3OFylYcfr5gjWPBLxzdvOf3fIE3s5AtNS4O5tr+ISbuCH2QCTx363lzFSKrCjqt
zUL4/NnmeKMmHQ9u+6QTeci+nypOstX5PsLblvPwrZZHaUw8XAeqC0xt0pksh/X8YsPNm+K21Dhs
S/koplnxGLswOjFjrFd7UuorUTVboSExVYmymB8DK7dLgslxeimF1eDyxDh/781ePFX3C8p4RHyC
QC/wbjrKOeVY7Q4vvhgpsxJQ8innZnsMTI2eavEiG5h1JD5Oy0eYA3GzfLaMDKLTJtre20/QG9aY
FS4nlgbruP3x7CmmUBLKLcxLBHyithkdCs7PCbwDBqh9/kKydF4o164gHYLs920jdEYBTWUxj40/
qty8G7KjEaDo9iCYYg3nlmW7P7jYXQVdfsI/iQDKDNOFi15ResFqEo92iNWVBDz7hHPXjOMY3lBA
wrt/20klYvB6pIXfE4fKQLngcE5INREuG+6Bh8zTZidjebiH1f2vXD/sPNoAY3YY8cX5sUl7+sjq
kfqd/0z11qXEx7+RzFQF6SuSfmZfm8qtsoNiB+uXOJIwtwKVnkd5LHjb/j2RnGDICzNj+zxZgN6W
Z+xDf/Xy0JZ0nhRBWykUL/QHYxFVeAIwM/x6hEQx095LGj/pIm57r3OvT8FPxsw2EkwD0RlEuI4d
+HvJOT+F1f0YnA3tjH/0nhjMbeikiIQZXkDZjtOlebPmyC2FTH/gK86FS/aKBYMibm78JhDAb4pP
smBYPCnBqmfDZMi64zuYILsomXHlE/bfeAH4HhqiV8j/Cs3aPgyfI6lpleG+T86noLYIxPmkB7cm
PyHd0xUBxP22YmYmYkozzk7RdGfsl2NSvECTJKwRw63W+Q0i0V15BYmWzy9NLjfdqypDiEgcsqQK
+TrbM0BAhSR+K5jXFZYaakBpsN1ergScKkv4y5zWMhXSvtIKmKg+WLQG6ByvcHqPOrmHOw1U+z1g
kSlaG97c0XiNhR5YBQSUe3gsB2W9rTCK+QmdoXL5jFepx4PDPwVniHYTjTTby5O2j/7bRPcfOgsY
EfcdefCeuqHdepGE0fUeE0UgwCrtGn0wDij+GeVe7E5yZnqPKkr+KwRBrgITurYBxk+Vs1iJ8wlv
Zu0Spj6dIN6CAW1VJmVl+y3CMG37/M3gZQxnLwISDXNzIRolMfKskB2zM0ObpfhbuJdw48wAPbgc
BN8ijHriCLVfaPjFRkUXhwiMVTDj06+JM4JeK49yrVb2W0fn1jOWv0bfVe+9KTNWYBJUuDmvdMW1
nHNFG5c1Kau9YkCcwe3uEXpVGobM13VDZfWfoXIkVoHgetYKxvLdCfso11E3qA+8RPHs7F9QJ48h
wWaqzKZwXh1+KgvuXowVhxyE57Bz1FNc2O6/uySOh30wORfkXmJ8mSVeH+bWqiB1KFDGpq/K0uiO
JjFaVdUi1lSzOZbPtWEbE+OC8STBlp3yDmlXSSb6PtpyaBlOO0yVVjVsdwrpvBWoPWvU/rdlfD3v
/FQjWYDNsV77A1/P5hDJaTO41wY0iiANpaaTH4+Ynynpj8lglI6CUgT05y5t5eBCffA5aIHc969a
TSzyXfTdgdvi9HCk0q+ZJidHqZ2zTG04+8/kupM0jakMGt9BGpBiJTJqVbwm1BX+XeRlrADmRB7C
N/ArssbUUvSYBshG+4J5boZDqooEC0+RJ+LqH+wbIAY0OP1na5po6F3iCLcPecBZKxCTYD4LrgoK
oCbrm9jW3dGsT6Bq4bjQa9RZAZ0rgvV2buX6bKgJLsbG2emPWwnaCJQWmHa7JyDv5Vk/YiltgBbl
f848wtFxTwToF/c7MFtjcwvMlO3RwvWYCRFhgDlVr7O9dd2isltwdWELrZOsgzUt1v0zNj3escF1
6b66egAC0J7i5RDaCqi3noduf8H/eSRd8WNg99Xlpja9AuldCi0VtUZD9cMxzHvqfPsjOlGXp1tQ
3cM9/oxDbXaqRFfRtt78vl2e1JZBRO2dHXxrWKZzy4PZzfxu1Go3UY/fyUbuJgwHqbsFtnl3Ev/R
odPlNO7ddXnN8sp2JNNlbArFPfNlkdUHknM5+/t/aDvvSLNTPtjrwzkxdSF3jjbH1GaJCY2RM8AG
WfeAQYiNgV7JOvp+FqWqeGIpm56fFw/7FR/Ufq/QlJTyzbW7CI0ag4gocdmw8UMHwMwvJZSRlM/U
VMXKIttoFdT/JOr7HtNfUCGThVzzlNCaXC42cvBauiBZ07crJUa41e/0CoNgAtGY29e49xwZGx/s
vgS6EbzjXLEf2OTtIgUt5p1F+Ihrc5RMIdf5sERBmldwJYr1gv99shu0CZb7LdiMFAhD6MP/2eHz
E+70HcuMrImTV9A3YY81kpgtyBMmeOP6Q59tXGuoXQ5jR2yvevORTbCxzuHPa/+x815QemuJTxIE
ll6JHVjNI/3BR/b3rrYuZYZet+bQGE3LrsXS4F4aRhjrwW2vOVk8SuM/lQKLUwVOo4ETCkoTP/8x
FBmZ6eRavwShkHa1o7VQcXvC/Hi+5+jdPv7uFEscw+eo+k6VRYhAuoTDzy2LSiHWqBeq3j6MnG5R
WqbfGfnqHkRF0QFrBJwS+zzg844khHZhldLkiduaB3BdFfhEN/G7dqxKh8il5O58lGm7+eMhgzgG
wdd2zEZjZHXDAsJtT9jrf93zHFOrOAy469ZdI8W0jlMCYnXnLM/g9QbR9EeD2ty74APPkjbIihf9
HdX5zYXmx9eZoS1BxaIlxsvOZZmOlNcymu7X3cZmWhUrJ0BR54/57k85H+jqX61OWQMV3v0lAldV
nWGeuuflmj8imzIydNlcFL97cL/tcYNlqnnBTrRui2ltcRjWBZ3A/J4Kt9AiMhnSvz02rVfYhtZu
RnsRfP6nWkhG6R3whrxXmAg7vj7Y07dn7lgN/KUrJiyExYqcZFOGqi1v5cxQQUObXAHuOhhwtDJi
cIOKe44iAXIudByAK3dgfvthPNjCksp+BIaCHAnkpTLazoGFab4XLjuzDbHYbQOfGFe905cA3w/W
d8y6osW93Oe5LuobuMc9Zumbt0pDnpbTokqg6Af7xBWFGcOhka4n9J2I072/5mC8kj6CKkG88Swu
3/ymBUvivqVBeMxl8c+dMNMBx1kN96R3P2D0EUBIeuyZumflsj3fmwvZTy1J3T5pqsluCohxPLlL
fPojtxVdf7Uz0P6gVDwnVz6gXBmxCUluid9dj+n5omFO+7M5DLhKSFAVUib6gftRtkRdVUeUGRUe
fwyqyRKzxWmGJeMwWIf6lT752c1ooJIJa7hqX2sj3VfFBJTO/4Di/k+rzQRznOhytMw0CVjci4+C
035pE/xwk3BwsGbJkqhYWh3VZrhQjbbB1qeA0pk8WPFY5pJ2q3YaEADRWtD2GcrJhYOoKQ9V1tP2
cdPGJi9NjThzk2H1JaWNsiwFuLKCZ38xLKrw0i0y5+WL6AcZGvbl8+Y9lcNSZ7ArS6XmZ6GUR4zZ
HFcex+/0XOe3L/tq0gIVOWYZOXXBBxdAsiaOt5Gx+mQdUktwX5pntTdFvvrJGbzbv8oVv/jtqf9S
QZSY/OvNYwn0iJrZaQXgrj4p63N1/L0qre9ek0PiwJdjTZ9VvveFhguxmbf+sgBLm2/IblRjKUUj
8OcP7+1FH4SVaVllc5ESCfbHu3sOsAQF5WRokxFblRd/WS+AwRH/Fm6wzYy83s9P8LY0vNfZQFX/
ixLxBo3T78oS+yzK4f96nqvWyKnigzlWfc6gBoAcwOUETuy+zI7ZSOD8ppee3HYtrFWAoUM4SSrb
c6mVHdoW+jYaLIxW21ad5K9tGyWioeWYxzp7q2HRuyLfqrCbT8TAJelzJWGoXBdq96Q92DYuW7ep
rH6jQVGrwd145dXb+GSM01egOzgaa8tbS/74n/beB6HWQGbMa0mxWSg1w+LLryq7AkFsFE1FFot4
ARMhScdXjF6EVsNUNzHXF2m7hd8GefvXDEgAFoNwBBm80VeSGvvrPOSRj4Rp4bj0gNfyJA7CoOe0
JbsmTxRxgfVQ92XTFghZCEBsGrbs/frDQOpNYxMczf4hxjallQwR19ukWZId6K1MVh4uvDcp7JRF
9os5gVOaoPVbzGyk8z/LKl6S3FcLfXx5pbZOam69oxsPCtXPOeFRN5H+gVuf9nPEcfSXS25n93Is
oKwTngeRRMxP4VuMJEeDGwjDY6XE4F/o2LeF/6L7x8JxKoVnHa/pzIrbskYWoSkEZd6UNCvwsBeh
NALhqBk0pWWLA7MesOJw5l73ZseO24ZFVekXEuoqZhFBgoLA6XcqmOmzslFrI7eEtM2XHZlpJ1Kg
+df/ewtxCW6v0C4fdPeqUSH3CzF0RaPOF4kBU+3dnQXcTngodY2bkjejsoDOxTsn7EPk12OjTH5z
++CBhxoJ6zu3l9cNxLVcDh1yViLFMS4b9GvP49ZGO09kbduAiYxrcqBcPh4kUNwG4mlALBX1iM7i
cBL15NQYgXW9CiCkfJ5l2N9MC/YgpyECJALaWb0QUpxprvKPqYtolCc3t93F6Pd6ZYiU72j+Kji1
ADbVBQgCOpo8fA9o9DAt+V3z9OT2YQkax5ueHi/XWzepAX0EZIKt4Fh7HAhSJaZ6m1IvdmrJKgMf
j+alZ5ljFxgX0pJ5uxhfTi6QD8lqn9XKv5k2LPwCoVtR6hsE+SWHwzcbYOjms1sVXBvSk92NFwo8
koxQArencAJdz3JgYi/fSBI3LzxltReax9yplqQ7/sXIZidGHbmEHGueWt/W5eNPqRq5Eu5/asam
4iVAIM5Te8kZadKus7AT8O1MVGRNYuFwwe7tOcEgNpy17mx9GZzbPoI9uM3hXyJ9njIO5eMs2Crm
RenH8M0S7FUHW27OWZKH+VGCU26+gQpaocz2TCYAgLyZpQNVcICmCknfgWK1KtArxahv/sRdPLoC
NaZb1Yl8jmKHdiA/U6LGJ+3ndqYOxqS+IxX2ltwJhDZ0Oy/KhJG6CGBoEd3qukimLjgnFaWPxc7x
dgdlqzLZgf14C8CWWn0gEAatgB4/lm9YnZXcxDfbR8eGvzldEajLp34uevaaohNoiFKVo1Famm/V
YGb6t/cT86K4dJNZNPlYYHuHMDsEg9hjS8XomG4TlHorm2ldsTB8cb4ChGwRJrM2zXgYfTlxCMQF
REsdr/Of/HKOHNJQe7uQmoGVwPEP3FJLdsjnaa7qbXZWDpAApxFgrJ6132IurKXrspP5d/FagHb9
ndQPyA0iYU2foUn2HYkOgCz/i6aOrcD4L8PpQci094J6pNjbsRiwXupzfMypxsW+iw6htQun0pNI
8RSMyh0SNtZPQO6TEj9lZPRiuFaZEhNGCUx6HTTltYhZRi8JmiPYWKpJJpt96q09fwYqfYUllQC6
R+iZihCbgz43Sa88/gL5a3yHKRTiX63Y0doXOnWpipDGpnEWDJdfckCRIa5oponw5yDXuBzeZpTT
Iok6AhRFrPrHhs19mzX1ARgEuLY67CIDp+Dua9QiablBLjQnRCQ2P/a1amIM/Ee31mitZso4iX+k
zKPGBTBNLlfn8QfOjNlBo+0G0KbNb2Q5xaNLPHoDTxrquoanTe4MDN4FeHVKG2qCIHZ8g4auZsag
0vQBSyvvr6RmKWuAO5WeTp9my4/0ZiSj0ZU4eGLe9Y+zNlb1kyjQ4SbFBOYKSshBkBLeSnhwcV3o
Te/6qDmP//G0TTc3QiNzCXOEmoE5gmML2g1V5DpYeAquARlMVSf61A7ULEvB0N8hO7yxtJx0FS0y
fliWI3xJrDvAN8b6HMfsMnABIBduOw27vdfZQ+y7uKb8NHE5ZGS5I07Awwnt48CHcoZLJsKqPOdt
chOAnP0i7iWQRBO1nRihD0RCalZkcS0HjB3M3IwWjFuft3mzZFcitPxifpnlE8dTPFwK1e7Fikqg
T4BTpyG91CEdTZaVokFTbMmnoG8/Wji8XsSd4NQmAmB2yu0GKUQio0IazUFQ6LS/E6XIBVIYYpgf
FAKYM6f5KNqYHvGx95y5D3nyLkg46IcPEL3yWq5zAP8ca7vfHjMeEthbaodCMObUWLMBEQnT+NP3
mrCJog881IxliLmWdc7eE794ZCUdRNACF2O+12CZah81632w1dDmdeJIQ0Y7qxaAbVWBi/t2l+aY
Z1Mv2aOnuB3Ywe7uGEOnweG4dJkKgyw3JL2LKyKFWwar21G9HsIFB2mF+/rrpZYZ+3a5jnZMMpMr
5H4EuafGuzrdMuv0XwTPp5U+Iz9gcfM1IaU77qJMCmtVcFYcM5rCV2dHt4n1vqijY915DiU1YSjV
9yulG73Z93Gxu4X3POlN8Xwc0Uf5fqesvk6j+SO8qX7zP+IsQI4boddsf/KOCBmwtibQvyuzH4Il
W/J6iKHtqoxbcZvX7Vx8g1fZi1jfAdYQAMT7qnSS317Zcj6u6XIpZc4XNgbOOH6gODjnNUDw7z6/
Muf482K5hL8efApuodacne9+HGnjuKNXjzxHTQ4+ZZ0APSPkDE5Tw24JRL+DeT4usywzy7Joenfu
qYqT+z6oRT87NbkJwZFjVRkQvCbj9GAefMo0wtrf7ASmvNfnfBTLRtTS2FojvqYTvV190SiViCK3
wKbRvfoE3TgWhmNcJ3uH4hMvewv6c5f0T41boenE49/vizKM7nlEbpYEpV7zohXqqV5ZdCCGM+rD
ZXlwJMaK7PbXdsUdxt7q269g/uqCUkJAS9TfAFcC2FwlBsv7LdvSTekiMqm/wlGu0W+2rXjKf+ue
NBcs7oSm/9g94yiKJ8LhLsQIAGRMTczvpPAigtII0uzCObV+jc6GDx9ZmHucMibSxqLlamS5d/k1
0B7/9zkV+kluU/1Rc8rNSL/qeOxCPEtqMergtBc64TswVZPhijUtdZVX46FZve/IdvK3KYHsxm0F
8jayRRS7cxWuRoynzl0M/ItCOAlMHwcaFK1XE7dhkbvp+Ca2cIxXi5C4R6CuaW8wEAE2uhO5JXGL
PiazyXmYGHJM1oduQo3pWe1C+UzRmgLSM0VAaePu5B4sb4iQ3gs8vrO7/2wZWO7XUbMF3L23LQxP
GuV2D+eQY/tNI0XUZVvI2IA1FGZl2XO7iLOZshi/hpN6Ved5nXZD8CWIV4B7wI2R1M7zivXpUY43
NR6KKQMkWAedeQEatsjNOnz9xrooqWtI/AtrAlqn5L58LwasyphmPDDIG6DsyYNBJJKaosRgKDGk
rbrP4dbgOGEewWGuQMTpMGnmBAHxUMbv8jdDIi/rSzNQWPCP3PmsHwl7QgLM9QC4I4lwwl3gM8/7
AwVtBzzxxdZbktqY/NFdT5VeQ6HrHNdr+V3aGgddJSYgefk64/JYhyVlOeM6xXoH3UP4d2gvVM2D
cbjP54zTA+pbATFcWumJGnF7h0SO2yztIZYiAGslEgrz4y+woHbVqhlKPxC7QQGU52BTSq6iOBQ9
UXc7pOf1+jmOkeWbVQK+g+EvPM0U7WjBw+Lj8Om8B5+RVuWOojB0Ll8C2WbGRPd0a3e75cxyl+1j
jFF8p5SXcfkT15AU3p7dR7aXLBwioh8r2o42jXiGbV1LE+E2Y+Os0mwybJKPqPg8JxLHE6BY922B
b3g+OAo6JURNiS7SSCGYstj8XyJCrhjPpr23NU5fem95zCjsO/idDCM4WtX6hIrjaF/Pcb1BNEM0
GnKxNCZRF1Plkrs0tq7dNUINwid/1xKUnmMHMM/V3J9bViMWLJCNROxayGJ1UeasiMc6nVvzDkKp
tsECkwWu3yH1mdlgLNOf7w+N4GPr4t2A8KVdxyQuRkSkIigDLTA92e3GVgk3OKUzy37Rc/oULF+n
afSIJFGU4xE/Zbxq3Okm/GFRVRWt4S6HInsYVEtG7CA1+2QUXM//66AhInzS0L5ImOkWoE07zOOh
lg/K2NC1uO1LwYMhdbJ66kMB8EEcOUBnOlQEFSuDT3j1B3G+HcJGfS6rexAiKw3D7Jvh7JovCmW5
3QqzM8/mOxaAoqtSvL3sK7VcIzr8eOaHrIltDKj2Z5J6E2OoPk+0dta7naWUFvYvjkCILZO/LyJU
WylvLXHXvqg2Rstl2N00Oc2weJ3eAhpkgXzI1oZyV29fOSJV5wGcicY0hdZyxXU+gMlghXao3Wdz
S7W+hc3hHieyENJ5k/Ndw3x0vXzJBwtS0hWAteVOProGg2lj5qFGueUoGSY8k45IRMKBjKcDXbNy
Fmp0PSwAm+QOjKK5xwwGDcAutL+7iGPkbsRFW7HKmWDhFuwiFCJ8nTqsDnpkcUSEZOCGqwqCmm+/
uBrthgo8onVq/84C+Ha7Z+jjVaiK15+GQmVPkyq0n09se7UYhSzRZSLqV+9dw1NC/mmRLHxHn2tt
muyHOEGgYUQLkM+DcMW2peEfEUVkGZVMKJ7qDN0ntPib5opUx/M0OQ40/ZZIcg83H4mXTb/9AgwN
HXTXOIpkGnor2lukSkgZrNv3oShy2+mfQvZmB6XZIeifFsvC+OOHxueqD0+x9BwKULq9y+8vlqJc
dV/3MmeBTJEWa+c87Wrvl2XL9O6gm4ipkpEWl/0S7GpTGVumouRYKt1rKCtfNVmAZ+I4XtSI6yvn
ftqGDan+BM2dWRNcJ0aIsFnLqMF8f1CNwz2ZDDn0bq3oT01m/ZhHhSKwJEZUC1AmN//vSvr8uC8Z
U4Qpzi4xgM9Eb2Zs9/AQEJBOd3KRudejRY5v45xce4EzMbdADsozu9kd9w2LTKyExidFf5wLHkmN
7ZTotyBAgbfpDuxt0xw/hgjfyp6ZkxQXo9slEWu43ozZaNF5u+8kXow00OgAYF6V5SbXE8zW6psA
wPG4oHjKELG9fC/BxYfxlr0ijvwcpT+8Gjahx3ORS8tRAHjTrPslZ8pQjQgldpleSlFP63jGi0hE
CtkzOXHrXcDaurw6u6tQjBQK+cwlkLu7//GGVm04cGbb19PZFIksEXzCuk2SiqDdv2Wa6mlKOjbU
7x0q17rcXGC4m/edQqPQoSy42rH0y8AZ5dkuTdWdlYCTexU/iBLrfP9nnadG/ECQczZ8E1vTTHv1
2K3I0nLrRSZoeuGy0B2aWw1GpTVGBjdCJJrU8EZgJx2WBmfjaajDyiHPD7CyZCSUZn9JoK8hExDS
DNSPNivdkEu1xmGLAiD3ni1CjFqGu9VCsUUL/WThf7NYF0oifTHMBk4QxPtkQBV1kJxx/hMQb84l
V6xTYWqouMTkLlD0zAljOGfqdNWWKElIVtjzqLs/DIXvyyy5CJLoEKezWdYR98/mdl8y6Lry/HRW
drVa4fxVkF0Ca+W7K5W6xa8hLrf+b2+/hhh71m9Zo5sdZPBEZFj26camR/VQgFaFcfQU8E/0Xt2s
pdxCZ0WEvCafJlXzE7OlWyL8nLeIRJWU5f8TMgXdBxrAf9zpSW9npSFqEsU080z6Z1J7iCrct+A/
YkeZWLcjLAxwQTfYgqR90jz/0qN/wHmhRUJD5SF2EmMpCpDGZjbWWHeZvecl+mgIZI7rzIf+Z4eU
e+p+oFbRSHbxQXvRG3xWcH+A+nD81Fe22Q49sDg4b4dE5gv5yvo/gXtSHgtIdVseFat/NbmjKkbU
LJfCIQ3rLd4pJqFuvdPHrCyaKFffdpJgGZjJ2UbHsVhEG0uehsmsBIDGceEp+Pld5cs4svZ4/nEs
5fjfRR7FmiKUGLYDWIWEkKwUyA8OLHGexKaa3jhPeIM03X7R1YIDRFHkVFr4+iRdawHDimu8UGi5
EL+Sz8WPPdnOuAKWns/ay8r4oI9+MD7qw7LdUKCupNY0HF/Z3ErPXmoM4wk2+ajrXufBilNbQD9L
hcdaYyScjQi8JF0Lr6zluPyXeG+5Ag7kZFU5o/Un3oH2HjdbsEbWvXtPUJesw//7Seaq35ti0Sga
rKhkCfZdxVn5TeDKx2sEGJRsjuRfq6E09qVjabAn85ZWJDY0OdjR6FlG0Wj8MZtRM9B+R+unXr/j
ZZxVwqqqtiNc47waGKv6ncJc/pMqDJvicTB1iwSgyKlVe2G/488jc7D8JQz0G61x6oWypo8JvV+J
9OW38ScJCLIKBvjWzTwOgAMpDG9vd6tjuA04cm7nn3yqzH+gyefd6Ho2h+0u75kB6tOPa+RANUH4
G2LxFFViVB/Y10UhZWlBF6SHlXiTmZyktJyXDYMGKAmGifp3DwW3rSUByxLtRr2ECW1zXUOeZOUK
QmgHd0klSCYcbDjsZ3Ok1D8OZOCbsAUQhyfC5n+OmgLz0hsj3jQEerGVBk1xeGP+UZdwJ6Ns3tuf
9K7fNKmgyDdkY3pJIVM5rAtvsQtpHTWvswUiT96ZHdHkYGwJyt0q/QbnYKzUncyXRmUDivHVcFfu
o2k1LqxgW+bBcU2/BOdd3WUTOlRwHU3gt+EINv9Ty2sAUCkKFYdEpDOiMvf0ap3vbhT6H+YGRR6c
6SZYQA7EZq4R8mAaF35MSG4gSHDYIZurGwirJlzGrhXCrvk0pnxNVoHGlyq4MdAVH1jDbbBKZzWc
oq7+/BZp/273VMiDS7fcjdeXg0DUkUIyzDn1kuyhLazH4jhNsxjakOiKaq8vGan13YgRa+SjY8Am
ro7B1LqFVxTruCK3G+qq3VKHegc979TWv2WUpdEYNQKatLXeHTH2O++TlS7XRN3KEhqNlKBkUQ7M
r523rEFYjincsDQAgrJT7LUIjVH+vBizpVwtyrhwwCOR29xCeaCXiUVd08U4J2V4AkVijhO4dslw
7HRarBNxprnrE3tpxxM4QARKRbHfnMwlBelOrqpS9DEUnxs1CoSR1WSVgoh+j7Mtb5blvFuAWo/N
vtiK4HSm66bqSwQTIBLDM5zXZ4rM5kiLpMxx/JOa3ndEfRT9KXnO53lAiEMlWwvt/dHlm9ky0Y1z
TzCkJpYo9s3+gUheN5k4YY1w9x+SxIsTrN3lKC3fghCe5aTA/LWxMqgnun+ROi7qMGJtR5w81ftM
Ua2Vblt2hV6PBSH1WofJtJCihI1pcifBiveiEx/E3wkQL0D/GlOtNkDal0m88kX9bHFbXlNLyOMp
IV+7D5hoVBT0N/TZa4/l5tEfDw3OcHWbuoJVYn77n8hREtzhy60PVWmVCy602bpzb92xpG8Pix4z
EN9Qp1k/w/P779Sakr7elu9TV1dB0yOTo+eLZiiWf71s0TqQ1RZrMkKO8ur4kqnYjvQ6SbASBbZ1
ZdcboT2BDW8HmIwn7kCpll9e7+2soAqcJNGbLlLc6ZY0R3G8+fmO4EZlhCN5iJlS3mm5BPcXnSme
ADjZIbRf87wA7mf6hPs6WCTb9Otf/Tyo0GB3Objw+PE6692i78d1AiHh/rg73QmiYQuImlgO4PEn
LNLtoar4vIvLTPaAZbSWi50yKj+F+S6LRnjj6i406bq1J9/p/1lXH1oJ7t8HW3l1GUPNYwrvnk0I
N1NWT/xuhjww5yxDIUEZWuls06224LCKQ4ng3yIWY6Pk4cF+sOZGBV+wFnmOzYMvgBUnlUrSNNUy
rJr06lGEL8x4SHzjRauajEuCVcujanwIX1MtDJqECn149j221R4Id77Ns319hUnzRizr2OWkdTw0
Z7N4NKQCesNDx62/f2yQi4RbcSmObdA0Pf3wJHvQ2VxHpVvD2RVyffWnyscgZDKQjPbxBGsR3WxF
b9E4ZjPMe5CcuGpFjZUpasJFxzrG4J7Polh0NlwA6zHRpD3OHHrVGDpe3C7E7/CIbRb+MTJzwdp1
p3nv0lDtOhVi29eu9C4u8Ezmui4xJzb5yWNiKnR0j4GSIhWY+5XMcZJe0WpvKoboBbPW9zk6pF2M
Psf4zFJFVWRRRbhDpy+Cy2tZonk8WL7A5BhSH0FbHMm5hzkUPIImMEZilFCtAG8kJaGib3jFeAyK
BWhKk0nBGF6eseQrheh7UVsEfZkWgfw9c8LU003UKT4B3hNd9wG2WYJdvuurdCY3C8AQ9Xa8Bvoz
Yq0x102WsT/0zTwKBQu436Bm61rebyRYqt2FooJFN8I78ReT/osN+Y0BCbXHmQMz0FsItUJI++Xi
SvbBXtSzMFVsfxJwkv0UpqPNl0/iixO8zjkJIaN7FnqXOyh2UGTx4TMvHXagK4ctR6tT33vmbTfi
1Kzh73WdidBZNrueLjW7ippVhGdwowBrEJJOMa1AxKwo2SJs3PgdapE5FQOvNE72BQv+ulg1SWeG
42DPyca+JmFkiPdqYk6HrYN+xVJ2HCZVE/ygTu8G2083HiiZj2sQaq2BGM+r0N2yNNSxCu9RghV3
+Rqi/bvmWZ7/Qq5SeipZPDeuxz1++XhhKZ8UHYX903plyzMvQLOpZxyPusntLzvnC+agvRK5Iel4
brYqoZdgXqkAVn1/ocPYyI/yQ8Midl2a4oc+xf4u1yfVeKBZ/C95A6wMic8IW4VJU0GoljZPrZbV
81ezl8gFl0UG2u46BUINhImWmXqac/OFsNepB4wiwvthLcbIfLBX8anDYc3VzdxuIhemHvaGfED6
y+PgJdvyzNPwdR6cnWYf3EIw3HNuROtn65tRLc6gO0lyumu4/xKrQ4pzIde0vWmzJ9VQKwGSuRwu
ALP0d96LCRR4xIXKLsyI9DouAkalh5z52HVidIECHqSdsk3P6uSskuG+z06PdMz1p/nxRoAomAYo
309i3v3p92haRhp/gaEWNMmmsvQKG21B7l11hefLMhhlsxMhZqIKAwy2Tzmn2GDUVfz6qrAUm5C0
5r3mTdrsKoqV/vEhbADaJ8DyPNoo+vA0OemKdX9GrdpCNvlsBMWmC+o0CaU0bNtpRwk0tlwRyIFn
ZAUjuRprNkNYZSzbDxTRvlMGOzXwFisR35khfCYdWPODhovk/I4L/31Fv0tcJe8qcQqjdKSDoxsX
Kbm131QXn/bmqtY0ugduQMRZJ8D261zNtsTXo/InnBMMVcKjMCW00T1xusWliKcEVIx3JpcCr7rz
JH7KYp+gVC47HOaNMWPDJDwDbGPFSKoQMAB0eV8AQCerr/HpsTSIFdAqQyHnPzBkTMtGRQx+zJeR
Bw0rASJAGwJY8QPsCHWGRYfn8fbDRa6yDmYr82/S4Gs/yM9Yk59lreJSjkefueAXyaeaIeG/zaDd
V5vyDi3O7f934iXypAj2VmhiW6/QkCHD9ER1XN5nQuIS150tbJ9qI7MI9xGr/e0x02qitwVqSmW9
mkMWFtIuo5w5O61EDxPFFZRvl9rxPHOmt5WPNKLtgENV97KzA4hHA5wyBnetB/HI6dMyCpRHM2LW
GxJ+l7l30trONA50x42EDIqCiEVsdkUhBwgWpv9FzYzeq6+WmRrzQPZIMK3sWWySx5GrWj1Jnze/
0eMDEE+I6UFOv71UgEsR9Dw0khpEFwLD1Z8zNpfcTFjHRa1JFiYcQwugDl4+jOg6mOk8jfw9B2xw
2ugzgP9Uxtsv6L6X6UVULz8MjmQcIublgITZ10ftPlXZgxNEVyUl3J8MM16vCrRAjZk4zmSB4gCY
mF79jwaouVETmzF9PiUHHDk5605qq+E+mE2ewdy+hPbQ91+vX6xiPUqCtegc+p9KuTGNow2ynkqn
RTOGnGk+s4HuZMGY85yaKzObLLXsao5Np/VByVFM7sTm76FI0uvr4j/wvj2XfNESv+BDEykIEYQg
HeOcg26Owu1CNXdSwIEenmOX2oCSDsd2WM1ZxUiDgpw1vhPHdbzK2pTCd6+chwH/LTVBhXEM7beW
C9whqpBHdneMDfG8puRY48K+XKoLZxUiDq1bZxN/yT2bzW3+k8Ocmm5DFurNdM/Js3eamfAq0LYS
ngyRVEGt8Oo2SmhTMIFyA6uC6v7ZHQ0J+IiXZacPY2Hc8K8O0Peoj8BniAwUifjOC3kiZyRte1Zn
f7N3uvNEZ9ayKc77PceeqBrMwe436N4vukSjmcC7T2+bPJ2ixUUB4UQmjMzENRy4aTCZ60nEDZxJ
bajqwZlAok7f0I3t3EVnzTrvqPrHxTO58HqXrEvtbBYuKbU1vMLxC4dPAZDmEhV58HcmD2ZWokbP
n19dsc3HLeN0EMzneyb7DsLSQIAA1XZzQrMI19yPBMlCbhQiiPBon48cFINFWCa7oO4ohAxf5R2N
wZzzY1pZE5GeQo5yOfQM1NzbCiNteCmIZQcPiG9JF4wX6pqUzHjwwJiXdMzxoWWS2R2tQDVvNk8z
LrOcwA4fprxJnGZr5UFqa/nzROSEGmtFmezJ1lXR4QswyaVUno31DYllQhGFidj/gpg4dOuITPLH
vj3mG2sd4sZu4buu0G92s1B+ckc/hlJLYvvYMkTnilCUDKjY/RsdTKKXH7nsyJH4Wk7UbQqN5J9b
e5EBUkIUjyeAoUQ8y24YzATbqi9KN612jgWQTNkrvIeLFWzbfgxaIL+Rz7F8HcuMtUmmJedT0oFU
UvZoGBps6LjcrfRfmUVDHb9aI67g4ZsSPsCynKQhnWpM+YxcgV43mO6WB5jxdWvu9eJOZyzjnAr0
kn4hVtauPubtSeTDpY125SzXmUStGLT0pO4jHfoC5yNfDuixQQCm2DJoBe7ZtnLLUJGQex1HaJ70
FgD8spsaaNfTg7EAp4UhNpHLsos83V4eq04d8+MnaEbIWPuOE4PWkEcQAk7yBOuhT92VM7fTmVmC
WvZ+RXdUpNk7SexVLSfCS/DIzBcEEs17zPmHyMj3BINGs2yHo3HCyCHrIgngeLQ+wFbEagRRpmbz
QgHJ1/EwGbPGe9EMb+ttRHz07V3bOEPRK9szM/sAk6MWjx4XVvTBNHeRm4JP+WC0gBWpgjWPP86C
zRDd/AXqIb79wDbo+eK4GhpT47ZJC71VwQ3SGFtpiZ+JwyzAVut0FIZMgmZWxPtF99mAiPKHr7Ss
jPpH7y//cEvcqqE/doGNaEjcePrsMtfNP4oI9l7Yx8sIM21Ydh74DY41P5Y+a9TuPb/zLhvNJE7z
LIT3jlAGAFtouYgMKkE12lM0OBPyKrQFeJfm/oOlVvjQmiAqjiwS/xqdALzOezVYzw+hTW/IT8XT
qfDCz7qBv3UC9jKERCOeWv8kK7kxU/owPIBXWoJGEW+EWHYHQEFOHO+twKzJgNpZOT8igsA7EF+2
Q2rNk+tF2xyZ2OwDng0DWhhuuhjDpgg5K1Gk50dwUrVa+l4Sb1c31nzPYeh3wOWnGNUUsPzz2yeh
L4pi0xtgav3/WpzxhI9wdr3v8S8KtmmkQk6ZvU1Kpp7Tq5ZlKFw8UpvOVWn7hZe9RWz+xAyYZCDb
zvV2kd01rKtjEFphEKnm/5GoeZvZpAVYP1QVfzUIbA1RA9NM1V4j9JZ6uxoYr3v3fuLdovPhshHY
20tsOWw42hXQZGQDRSR7V1B/Asq1gl0ZBCLYx9uyyZt3RMxJILpYgmxzDZV6Cmtlvo8=
`protect end_protected

