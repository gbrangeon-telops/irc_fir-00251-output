

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
iEtOB5S3Q/0nxxj3yhZWc1e9CYVNx9kxE38Uvw9Q5GTpbeWA/PaP7MHi1hZ25jWcWTCQq2m6lqXe
j4/ejpW9UA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Xuau91ineWkILAnXNctj7ghjv8v9lVNvmGeO8/qKPRA098IIoEEWbPkQsDw9y8PN0Kc6j93b9RA3
24AkaGw7vS3twv084InDNHpEnlN63djkx5ZcyOiUohe4xecSmu6QA9TFBRDs0Woq2jQD5/qd0oJL
/BaRHEN9wihMkCnRmi4=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
DukDx60lt5tRoBa9fYOjxQXcMx39PTzSzi3mfBKPNtGRH42SBSoh47iSUDQLozXc9RVtQC3PW07a
TdEl+U9LI0QpSHNQLVojqhahZCfYOg99dtV1mWPojzxtpV99k2zYX2J3PXN/YbIzV8ZxTpLcq1Jp
CAIcrPJ/34KYVzvzXFRsvxEfk+CxS8lIGg/nVz9ZI/SFfi31TG5Gc9nsiydQV6NxDLfMTIZ9geQt
WjMt/ZdcVbixfIDM01Blr6PmvrTG06LX8uxL31TQuw5SZfsZBAh/PoXSzsMleljAYXIhMhdSUOnh
qfkHi0I/YHOxbZGvwoECi6yzPk1O8e4p+mbfJg==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
JfFouWl9C67kV59ngW+xbX0i0eu6h0roaptqFtm5oV4WYkqMJEDqBwmHay9e7sJ9CO+K40RDFIJe
/eeImbz2XS0Q6PwgmMgPAHRoOg4fHkGIAEugmb7hj+mXvk7iQo09CaB7HocKsvGcx4nu5U5a1pLQ
6UjYczksNjCCieDaJQc=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
RNy6OyrkxjF2nMK7NTVKf+mkYRQZVhnkvdhxFI69h+pJImlNAm3GMG9cNkr/rYPBFr0KpngtSqYa
zub6qdQpsLCoZ7qDFdEc1+wws1xQHHeB7VAyyByyPc8Chu9XZcfd6cEAYC55a9lNvtmKoAjppEfF
hj3OtTTwZQDicoWmteMIzi2n5YcjhwpDSzFHpmKq+NQje013CABovpP0/TVMHv74ZpkyX30HW4tb
0iH2SzLvUD7U/AR0ul2kht6wcMaLE9E6bQipSYn1DEnfUpMfQgGpPJCWjykHayljMFWfI9ucuNXK
1XTo7EI77uCstdWwv1uP3ZSQ8pFNDP7NXG8mpg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 9552)
`protect data_block
0Bz0qfDDU6RH1ap1sofOA4vgoomLxlaK4R7/WC7hP8V2VF4PQOpOGeFiJhpWt/szKsbxveRxLs6f
BBI3ZZzdAedUbEQOIvfDyDUCECAQETjRIDlPIui1F24VpF4drDxVGJ+9aAx/4HUnee5EE/wQncts
Sws0qf51BDXMUJ0nCKox+4thqtAifrQEip42oAqpRVCA+fC5QVkJgTqU1m9NkQmQqo3lL3Oe1w4M
SZd0BxWgdpVCbfMUCSjsSmOaVnv/mJgFMkkiMD/VZnyYT5Mvad6W7tGl3lenQOgVJ+jeLPXeRuz1
0mWIzHpbc8jQj99x09/cCxGY2mRlzhhA5uYdkai93n12dhh1ShXMY22O5UN+Z0JJc7Y1m/+Rxeoi
qtnUtCDqoSH/tPHDzXUAM2RlseiaS1P8v+5siWCwT8N3AmvcY79R52d9Tw2E3X6U/LaHTy4P0BJd
PWSFsuMS9Is2uahFPZ6f3tnLxYgTUzFmn6SeFisZcjGFAHi4n87OpNMe/0UCYOcdbb9wQFNWRcUS
JqnQq7L/ZOoinxRbISTk3ayZaHfC+itSwBl7qqaxRfhUykrbyQnaiHgyUtMl9MtU+EgrPvZDyDbz
7HFPO2Zm8sLyGHP4gghni3Nq7nZIBXS93KsSmTsCwtt8uAi9OPzHolljt82yqYeZTIRcViMhlH+v
7iKdpHrDVRcQ+4szpbWBAZhJKQ1vKL8FXyticxwfl3xZTzyB/6Xum0Qiv1FT3Pf0TC9wIFMU/13V
dTdDOdneO8Hp3vHZyugkM4oHtG2l8Z3P7GDgNt26wJ62UV6SwkNvxKGXUaytf1vZpCMGq+HLkD4w
Cvch7mx/ZND2c93gJecp5ru+hk6ZW6Xnhj7/sU9FsiTnmL71DOrT1tbTgIB6WWF3AGKDzSlak8Vr
me1KFVkf+F0rv06T2yL8tqmrk+455C85n0Gq9F+DxR59cG88N8JSnu2OLA+ebDN1FAPrYL20RGIf
WE7s2eQAUM4c+qkZOCNiokl22LwWiKx0kI256HUAg2aizdnMC9d6xsAMVKYynmTD4mCuFYzb9yIb
GqNNoxlOT3dRCSDn/7lyonkrbrkaG30hw05L0Nqs9dKSe+1pkUL905ZsRNZ6nNXbkVTHtt7e0sgG
0C49AWe7DT63gP/FohYxcz9VWG3+B5ZCSTI+MLy7uZS/3PoEKi1xBJ7c8vmhGFJ1DNQZSwFn2Igl
53kmIyNut3F+gEZ+eKe2vVTRlwMPy7W05ZoqeIRWF3KPOSoVqiki3tE9ptVEOBGQHvW96R2glOcj
Wm/tkX1Hg4kd3UijyxJJ9HdBq7ZFfre3yIE74pjK9+XKGR6g88KaKrTYSbebIZj/KfRTyrgCbtbu
0tjQ5/KZvirNvmpL+EIHOyowv8psf8Nav7z1lx1RocI1la0RtDZaVSvk8fNnqPfNBHuJwQo0S4Zt
awDNnBosfVfERIu4PUga/7e4rNOrzsGcAB/pLYKgBKEP07YNE4+54fbFKYgYd7YAhrxLBqujAGl/
CJCRthd2as6mLcgVtjq5hn/vklNahTeOiYl8EVSjkS6EBFyTfdiAKmZNNaFVfRspTOivypWxmB/X
/a26GkdSDnYvZIehgkQYscCWGxH6CqTjPDWxerGpeVX7IDj1gUppcGZBLSIMiTP4B+rH6YO+7/DG
ymlYs/UT9lCwdhxsFDA6n5KogZSL6eAll2Pq8S6XflI5p+WhrY/jDzePNg5bZJu3zvD4H/2TCXvI
YvWHt9z2YeiYMf2TaLsx6+dEETzgf+vc8obO1QNCYgE0pKHtMJVkurPXC/JnPqi/7oYzEmuGCVO/
Ss9THI6KSzTB79/jK7EuWPxoP57wYhNGLJl43NT3HMNi20aJeFaKZvIYad7pbh1Ri6yCo4+qXXcY
sNKI2rJ5EKdwp7jjPXmE8fs/gFWaA5tgsw4SJAwdHHSv8EasxUirLVY5uZVQ50o3kIyLZez2gWJk
YdNFTUrsQGsS4aIh8J20y04foiJaD5RldoYIHv9i3A1Z0nihXFJxxIFZW8DBiP5a0eRzm93eyd2i
BIR2+Q4ZwxtVyO6hkdfGniB/OP7r3gycns3U2L/5tLa3G0iKVPifPG1/Q/uNiXWlSMOAS0lOAywC
BQUaBbbcKE+XR7YTy6QszoeNsLsMkCZP/Xkf5QTNUJj7aXWCvX8Q8VV/rmKje68sV95MSw7yNcHB
+CGARt7FYAdPeeacl+Ynk0jGejIHON9GkbAE1GWWi3KDv6dDjDm+NL3+z874dUogp1mwCU4u1dMs
/gaD/JQ/XgNJ+ttykgs6ybWt9XjXM/OXBML4U3rXRU6Zp/kz1pNg2tvYnETbQMQA2RvRMZz+do8X
Z2G53dGzxZD1d9wkHZL8KlIkwMOEh3daKBsli2N/akiKt5Xx81cn85Ww2HyOvdKLb1ayET8Y/Cn6
swa2/iJyEfwtcaeofSfwUDLBorFEVsNKTQe2vnTlrPs4WurjTzSO0V9T5Ggg88JtSehXcJM46EkO
1F5dMIyhLSbys+0h6Ro/CdzJpZtRiHsviFOofvvKTjsaQ313N5/oImvLDYKc1e99lZS2YMLEAtt4
eoIgZVuvBlRgTRFrvqQDiM4QmKD+T6XzWY0ysONA8B9NIznk4Mt90WXBXKuKLVBEw5+gN1lmCsnV
jgTOXhG5V6UvV516Nn3dyYgVYmGw7dJIi1N29WoEuo7PFPczAmxCwfDWjZlwelHoco+bOw7WWsKw
Fg1Ey1ZxqM+cpdYU3tgsDwUGkYp1L8hx3Vc3MMo1X4/zBzpA7BfZubjVMHo0aZp/HUKhLY+r/ALG
HDUDuKvhRNsthMOX06MjNldT48OSFQCln1FikCnnUW5j406JVdjpZOJcfsQwZqIz0wxyLLysHuUj
+pEMmXzOzwq147kNnZ2T7gC3fyoJsMKv7KUwQdCaaTifUqNNNcYqnXUbhYS6eJbEVYBeKwYymIZv
X8+5H1KwXE38yVmxtD8iHMh9tIKzqJ7yStryu2Jcb/hFwM9u8afwgEasg99WE7ubO8ANGTVaRb1E
ySZ/SPNCo7y96IZ1dN4/wSk6UmsWddyExt9O1DrJyJFgXgdC01Q6WsX9TpkuNdQ2RJitQ1U/bb7n
EdKQRgP4ExfIgGiXISkP0/8GaZ38YepUNnSgBrby6JS/jFij4hUDGRj5Hsh5no/y2aU2azcaAOqK
UZVZX0BFzhFsxJxAYn7Te5WqJxo7vds3Mp6iXsOoc+Q6S775Zc3abezuve2P3aiUPKlK/m/Fm13g
IJ1umd/P2j2lwAA/48FhRsjzEbO3bHx4x90Y48wmy9Fwta8uWSxvc8M4lpO8LitjvO+xjLrGPDbo
bl+vPjC+cP6DU7yOhk/QQkBdn6KmU23GZtG2YECtZMZK5Zs7+QFzXptsMwP0X576y102uTyNt/4v
0E7DQr02JLXhi9lqI5cKs2K7+lilAbR2euoSieLUcSpq3Y8eapRb0EX62NZiKDhN1CKd1cbLtemV
5Scp2DEmCHOLYXsr4gsYIMHyJhHKVl4FotDFswIt4VurwzeA0x5BeOJ5dRiHVkG65KragPVI7dmD
kbGumFGbb7LQhCvCuzcwZNIk586lwVTNiaoGFlIdmwOTED/tHJL/U+H+ku06zJBn4ScX5rWmkpTd
1GJbWRd84WCAQuX0RK1prZQ4VDK8urR/Ju6nhlMifP6DtQPwrAHG7DfSt+bJGXk8QkUh6ync46Yj
qqaRF5ZnhBPCR97gU3UCvYSI6HIq9TKuonKhC+K7dPlioZD/iT4lkoBpOlb4n7ixopY9tU8Qahpm
vfBSiDk3v9OcEH3TLPb2sWTpaOqXifMW+IGYqfhaTIlk7yJ0+ae/En9zszhrddPR5oMw1vzIxEAK
lROVFCuVbTgrVURL7YVR6qQ4ab3NXf1JHY0DA2ILnqclvubECZ+v7vEG1FPnykaKqVUeHjkKs1vD
H1rUB8R1mIVWzWmSzpJUcDbGUrTd9Jpg/ZyJ7H3E5gA4SmMyB0mzcBTCPrrdL1PxI7JR1dMOiLJY
uW3I9CioflfhCnfAE9P4ofPUUgSu03IqnqyrLgjkDEihdGHzVxNdbfAfXubUQT236zefoE+4OZBC
33hHCqyeE2kv5oXf7QS0iep0q9w7yqPNdud6n49UkyOemyaa1h226oOfLp0doaKew/inESqjW5pd
lKk+TjycELEvnrIG1Y7ZRyRyO+aeYEdUW5kK86W7gKRHzLlXmkgfmsSrmLfgMNx3f7GkDI4OOL5v
BR4s17OK41a74eCxThvD1hAZlUjXUjhWhCMYd6T+lCTxjx+EUXOXL1w3qiHKMF6Y4ObJdd50wHYN
LzPzfaa1Dg5w69i2esS6tS4Js3XHSy0CIrUIkEW6pJQDEcQPqTVPfV4tqxLBMQ2wzGM8R+F7q3f5
GUD+7x2Cl9iy1Jhj1RrB5db3pN34Ifn2MOkMkS8TtE6IaZ5C7z5gQs2iw+16JUA/N8lFUS1H+q4h
4Ola4Yl2VUcLoNLFIpoi8j7ehm+a6nvrc+HQ+Vr90LUmLNKTJVDyuMwckev52rLN2+G7YUPKgt1h
ILlgt/2laePWpiNKw0RKdKXE+ysG7spcsgGV/gjeWuXxJDtRXjEVxAe68oxA8yiqFolg1ogSQXY/
G5mNNVX5OHqWcpKUlrQQdhGozypqIMjUCQ5bXTcIaaLLc5sufhEN0If/qzPBcIbqXgnKMjNwQp29
ZxRZAPkVBM9a5ZmGViWD+Hgtqx1pMhd7/71CX65MkB+oifi/krBAuG0j3/IjHba2PuO8nFrNUlqW
Z+v9pH0GdgtSONd+9YEMTYXDWW3F4A996ojpokyU9ghO9oeJSHnvcQDxN6AZbO8ecU4fMzj8R6UJ
7KVvQCewA9wSKEhBmt3QxsDdVTDDMC27FgelqPou4jUtCekHUvAihf72ijk6DC/LJ9qz0XYGQUFk
/Du78xZZdDxO4wwWnzt+oLenfPfP/Hzm8qcaImDsVW5U088HNEktOAGYPV7VDXZ9GpJ9I5c1fsa6
kL3ArmqYfv+b1kbJYje4SuI5Uajb6HEjQld/qZrMvA1w6Rks9+7E0A3/9Gp/EgaA4oy8Bdm8CMAk
/vxzT6f/qGxEME8pA9ky4D2CFWQGNC2h1T7I1dza4EPP2yPO88zImWQaFg0mZakP/vHn0gG/Xbr1
xLtRSteCetOdSu+3t6X/wkZ1RG5KKQnVB8WIK5zZec4DCiv21tdX10WakkSg/ptIITl+NCyfqH6S
g+YwpxaE2MXlY4uyQXtGbic6BlRtZ2QJqozQSYuhyLJkm3b48pUTR9ri2OIfSXXNpyljJ18DeTV3
K3XrZBB22nyhOOI/nU1TEB5bxFYWsj2mutfCYD0z8snuF8zHBdfqquwn4k5r7s7B2cIx0WqHVSqC
50IbCCgAVmgkvgGGXhjs3LzAk9PzWsvesuHd1dbN7x2yvMC7PKbo/FkHwXyRRAwJTC7JPApQq1yq
ghF5MDHo6NslDA9/8WHCSaWPPjDeEhtcegyb30H9CRaPlFL7zk5VoJIhfQ4oojqjMDWzaRy4X/7G
F8bjohvhROrgFEWEGg8sfEwa00OPOvVWmcak5F+uVuNLZzTTSrjDclVc6uk/eqT02DRUksZ4wbeK
eL98poDv0/9/opRH0wpxVdpchMescfcd9cZbT8kA5E5ffSnjFvxoemKuxuMzuESL9x8f6q4cFOXX
0S1JYExpeHmIFukdoM1+jULodPbNYWAhGrWHgx27Ze+Z5cJ7FedYiSgiISTP3qXVEzcu7FbjeCJG
nZ5zbU44hjwF9/J4ceRtIX39YehdWyMuLrlXuPOHHzKMcBYn9CHUmQXvZtBJtPOyySWI9FLu6MHo
JUrEQ8JNwDSHy0ERbDKtgi77kk1DOnewURnQvd9wDZAwVWfNRuYEcTeIB+DUUzAPBUF6zrFnuKio
Ek25PKfRDhjgagMlEvqHDwAQr/yo4GmtE0p9PAFU4SGhp71oyQ/dcjaa9Y3SUkEe7whE3be1LioF
lUalJubMDHeFbKuhdiMlXl8zypQhAV50/lKoOfQikNFGknfuNnA3zuXntOFYVVsZMK/p2Xxm6DF9
ltEIPk+zfJEm2xq9SBsjsZjKSsSF6bLZsMk8GtPkdJ3ANG76ZttTYAgclmJ97zS78FRS+qcIDcdk
y15eb6RdApMOkdYBW7zTPmmR2SFRgnK4aBVm5joKQ1yD5BYsLfFD3+VNPdc+p2DK6xH26drMFQrF
1E0yHAAl10BS6E+D/UVycAYPjwbDHMHEMGluJUUZYlo9yqxZw3DSAeN00tiQo8jXjDaphjQ7zmGu
VPQ0PWq2121V7hhfXqwVvk3lbFN0MKVJQyIN9yX2sfdq1PkjT0QTikyjrQfIo8Qa5YD5DISu//iA
T9lXHgi8Yd9QZ0aqnjNBMMgu1m8/SyZur6ORyJiR4lFk2ccKTyNmvBxyh/O39zb2gv04pwDm3tqm
BASnVhTK3NxFv0w5aIbimygZ6sQqXoRhD9H7oEFIoLJCiKvsOFhQhAWFx9rM/ON8qQSXniu7lLl8
bn7aBjIpWA6Tn04zT5x6r+7noGfNE7nDr0aAJUPppoYF1TPIPDhGDBUHosY0Lwk/3klGmbe6MkGX
H2cAIPtTG6nKXUXxp73C4JVPuLN6AU3HWdeWLySRX5NVjjjh/mKFLxjoIHybiL7QGm6/145aZf1Z
NMJPZ0AVCfEah+8XEAaI+5xTBNXPgRLi4Ne1Ib/zNfdSnaUZSbdfMKpYc7BA6IGXif5pxDWW4kpX
X5sE+MhEf84U3RwVWPpj6SjYnPf0hz7tkNZLRKlvCHCqcSjLLPXInU8ZnzgDF/N6v1QoP7BZbGZo
uMXOG69ONiz5Zs4LqpC74cJSSw2gIR7QzX1kTSnhl8tg1KWl9Kva/FMGcxEDvbXoUXs0qQc21cYE
ylYeDpyJDCJQzArtWnJRxTCuex7gqTXyL3So2ZonJQ6MHQbwoyvqQeCR3XnhaMXIL3HHFqOMt8/N
494SkqLfaum1DZaB/sJD24KcOfxcKyttCuNYNd2SdzCHQBooO9rPSRcltJJuOdYb7KH7bKYB1rVw
vK7UsgQRfG3cJUVJNO4hmDRWIyl4ZB4D4G3ee0pne3lKQN+uAQSJW5VUeOiGcEv41TqLN83PXNOZ
jLzL6WFAVzHlCXg0i1nG4QCyIPKV0g+g6SA1h/xtMf6TbnBcdUBBqSRIsxd6e+dcfB1xQmcT3EKU
OUZb7FlqXOwCeBdOOXPN7l66Tk4uhOUSd1TPlFX08ERs2fIdOVAlNxWaat4Y+q23QsHuaJBMtwhJ
VsbBMYNH1YnWz0TF2UHRaOgdSwh3Cm0UZMpBJn09FfGHjeA81HyQpw5tyCVbbvQPkIRpJE2oHwyx
FY283ULsV/ZI816M1tBpdrZwZsuEDtO7bAzLGUhHfzcVDXBBQCkHOrvocg5y+tsFx0LlECQH1WzQ
USlDwEo0KYcxkSCM4DC9sst4Ogjq5RalKB3r7o5GHIzKrshRbvXnm1U73Eo/PrTyF3WaRvTVa3Pl
1KAHbxoWwPSC4IaWUe89oKXykFiI/+IeR+gkWQfHAMvs7gNNe+He1KIdOe7u9CdwICVymDcVBJM9
qZpE81e7HtJstKfC2eHKKltGGuYEQHm4/O8uR4R88VbJBHp75IsrB9DygwkGDIs6tr1YtJ2A+SUL
BBoc6VfZcVrd9kMw7FOEB0B22bP22P1k78QYSGyYLSqygaNTF2Wf8UFNs5D3WqQ2VFozQabK6th0
/OyAxUIpn67WEqBjazlFfonJ/uydtksVMAxKyb+rdaVb/+WHAp/saxc1NnQ6Pp9B5TW8svAvEsIu
IWr9pVATHEcEXGuaUNxCtFNnrJaGnCkgyx9RPoFHCic04ShKpBlfShVnEPspTQfreCMw52Bz49Tk
LyepKcomfB78P8BEpq6QwbILAT7dhW679VeosPyQsfGRMbl5S3/IUzHTZ1SgShwfRUpmtjKw/LCf
VVi+4S7qKoJx2PGs/nWCkfkQcOMQM1c3mwzFnFtRr15nYX96GgOa/T+2BJSFs8rABQBbb2gOZtg1
FEsF7MnL0+QNKoTb6AqWRdFHIuKAKrd77xrLPU8reQ4n+Ek5wPYEhddDkWeI0d+RK7skUQkACHf+
96ARDijMR3AWHhc0xcITqlOeYFnkDvv7cmESR1/9t5cXAaWWQpsTwP5wzdIWJxqePZ0QhPx6hTTt
Tb/a9db86p7cSx/aOKFQ+9GCBZsFdd0HRUtVherH/oH0EdTVkZJiaQPfGasTFT8btKFuCmpomFdl
9xTIL7IVycuQQpKpiJQP8lZS8ytcrE64dfkovhLvZ53hrzAfZMQ623SoBhk4jsFBmjkqA2N/+cJJ
ALKCSP5BokOGEfmcHGV4RmSzFmScIxxHfc2nWlhufC3nZJECpzTCiwTJoFw9aSGldMlso5FRczQC
7YoDDT88bnQ3eOu+CLL66Vs18DpkY1YzlZu/NiOrlwIhgI1/FHOkRo8fcoE0QN/t5MbFraHKMVNt
cTf9gPtkxNHuvWCRqolLt7JKjkd3kIsG7eUj5vXWyn4y4eS1Tvijo2vAQ4QhNx2paHa13yIMn0lZ
u5p8ytgyejS6AgGP324Zjk4SOmIOokGKFAxlY792OtQPFbifeOrYjMTkmYViMuB36xUL2aD4MRbu
IJfJzwdDejc5DtdtF7ZsbWWRfzfHyjGeZfK0Mxjopdwp4KqYmoFmAhugIf4++QbA+AZhfJtohY8l
kGUmAclXYzWH7bcx61N0ccC6Zbx6f8LQouvIimwBLCr/vyQoVdS1/jjikmcdPaI5YJLkmozW6j2/
e52oCNexZUnWaRCwcc+r4Jdjtz7+7N9+putW8kCY3j4AHMzs3CqtxV6HE3yc0CqKho31E9EqjYi9
alu77MzZ28VL/DCr7ObVt5t8ZwiwWzF7mnyvm/vfMhouKFhXA7dPnMDv+jhq+MMaOWkTyROVcY0s
Uk9fd3aME1sUGq4e/3AucFYrxmOGVX2zRmbDAAXXi5NgUQzaNXOeJT9aHrKnET7stv9jkIxcJGCX
rFY8OyAqn010hvM7CdiQ6MbTlJhlrhdx4wHtrygyvIrO5XUQeGHHs1JaB8AawIafg4eSOHNWOYEX
zFRRKqf/dEiD0p5+JYkTNvOLyORhAVioDCdFLMEbN0llwmiKEDady+YVeTf1uT+HNZpno+NYt3Cs
Fb38DLsHlmwiw539AfFCZ+XPBtO1wrcewghdyVUDkzMQCqSOICQnUtpuQwbVNyz8dcpWaWoddww2
nsaSt6gnAn+wRKvfBqaaqWDlFN1k3erTbMSLzoADHuxFTN6rl+MrGzX7KsypRHXb6pyb5PVO4Fzc
mDM9wPXGsheVgKTAoXy2YxjioofGKXXPa3OrmMuy48jtijGJQCyCnCF+tVIzFzq6uRHVS+IRN3Qw
pOVh8TfG2aZNXedfL5tG2QDmedealBggi0pu2EV9UBVEwzZ1eq3yRPri9Y6SIMSgfDCUF2DvZ9rS
2x9bUd09KRjnqpBnxcnHqpSnyC7nlS0Fa2xwXncysHUtfJNpt4DYohYPA3hTJO51CHTviex5W+QE
8leQ/HVDuZgGNobOVXg34WL3xyzSO8f8JtSn53FvrsRb9cja4vwpPBwtJbuDN73vGNLPuFc7Fq/h
fiCvLCCHf4SWDUg/GWk030TaS/p4GSJXVF65gT0oWC2Cl5kkUALWVyz6UOiP7u3A/+i3diwXbe9k
PZv3LzuenxLCDL4oPIB9nzFmJMurT+dcJUYVlQO2SdOEsX8NnjwvgCAXu29De4cPUVJ8+Qhg5D9t
d+tQgn5p9YEx0Ky+VlLxAJf5CmTIIMNbPLS91W2TkD2DCDXamkBMnMK0TPNC+g0eagxx5u/gtzpR
gXoLXdQzejYsPMoIIdUfopIeBdyZfbxAe8Ll1BtpKxoXHrvx+QbS25P4LLFURvovZjspOzJ6Eswo
3zo6Suf+p9LArDhlZqpARLs41gVa8KSznmZlVT2Y/Un6yG4ojEHcWG175m2OgEJodxmj11d/535L
WBk+B6RSe0qJ+3IypjkP+CZ8wh3pm42k0DRVIN0esCZvI+r7galLjaSIfduwcU9lcxsP4094sjbu
gRz5x+/fH3p4lND2Vg0HbnG5V/YNXeISf70zcN1LeK24FJDRht3fNoo5dmwtDRPpTWxemzLSFF67
AOVveKv4evXesg1jYKs4PxohDqz6SYpx5McU5cpRanQMdaoyje6NiL2hWkSTWpt2e2d78wWPwrNq
fV9y5wRlKb8HJQHirJXAbW5NeDvHDHScBOaQrNI5frp/0sZ1m8JSmAVsLayF6uJYOHmx61nL0G9n
+GGNMVDdJ7F7NUuIg/3RooEJ1u2YQP33NkeElkw3rZYXg+NWB2bICCg1/vSUXhcT2KWFUVKdoxRx
vVJpRwlogiziAjP/UT5/rpuluBF0O9Sam7CjprwBusvyNoK1ltJttxwE/+prqG1oRUVVkpaQq+bQ
t7/O8346luJuPQuTCJHVfYTBhh5K/xspy58vpZFbvfwp82nb9ZKfMZJMYtNJ9HtBxYDW4tTfq3zY
8yUdBFRu79bN9w+uKk6q3DC8ijFOEzWWcMOMVBZqgEHJoqXz6AjeNq3H6n4TlOc04Yh4OSSM51X7
JXIgCL3GiPgfkXOR6+8vjVvc8k0g6pyjxnUcsYmIXBcaSZPtzUEMoCkbR81Zd77xrUYR+p2BrkjN
B/BNq3YSVLvURfn6lcPAathDYjDXlEP5M26fXLM7BGhTvJrdBHMvOwsQpfNa1b9+nKj9DVpys0z/
YPoZTKGXzoPh+rjzCDTwgdLIdQgbVvLDtNesa+pTBLRSk3pZ2D/oQkRt9yA/g+v4ckUxpKF6SPA9
Ye7OEcmxwVjn2QXei2aEtP8ioxJgM/erU4lmE0HZn1cKapxb+2N/vAdyrBsLEqIsLXXaOUmE0SY3
g5kJKP4jndJnY8hSTkF6h89a0noxmD05L0LFdrhEApFlfPnN1KEicTZYY+NZ7H5q0CydXkp6/x0W
Q4jb9MUrKCa9l+Oxy/vvrn1PfDT2svStZy+trcnZWAWQZ1tDb0F0MBlYq+NEYvDNlijXY2XTKt6W
urFdDo8JYF4dId2QQDIOVhFUPwq/N/DLoxbzKYIBzmCH3zSbhZefvaDG1y1VPtKoId28ZHAW7hiE
lCnmhG1Ya2GmCY3rBV/z0z87MtdNnXYmZ49+H3mU4zoMDEXARSAaOnx3300U2Zsx/0kgDjH1d+No
sX4XbTpKspqBxfNb5TLF6Q5sigbYLE3Z9EKbX9TSa+i4Z9a8oalWhC7sPEfXCaF1VXAUIQgmIVs1
Bc2ttS9ifCI31XNxt4d9UFRegn082TdwfIXHt533Y9h2Oi8OD4cUqt7ob4z1DawyZR4r2uPJzsvP
bgc9Zk+dPGD7F/EsBeyMxPZGuzWTCzvt0a02mRgZzzqhTIbHOgw6sWnmvBGD5/7GIjxdM3x+bdhd
bo0yBNK8gGQulC3NnROjRAoxFuvDj7ZhvEGXANgzORRanNojeUx++50N680E0d/YgOEBN5lg2ugW
UDHvSOQWsYERHRV1hPvmh6iQ4qEug4V0BVhKy7qdnbTvcOYSv1eNj5FOdptog39im4oh9a1tTlMT
gXKdED2VZL3Rn5w+b4JsAIOQnC741q7moWAu+yr7TTDvoRjs0fvaT5sobMR8rbFN1MS9Dv3Mq9K4
p+f5V82nTd7QwWda2aoaWCxuED71UgA/N581V99fcwzrMeYL7PnYTuakR55TLMMcwaQpz7XJXtv6
rzAKyzDKRfDyf/dtWkLPoYHZyzZ7suzR5BleMR2KAJfSu6+PrjRgG610uPzUJ/CGFsXavWg4bRRP
nj2MJY8V1fb4Z3MPd0xCrdMlo6B3EqL47YYaDZ4+iRf3HEG7ev3jliOEum4Cu+FLKMNK6SiVIh96
QtDdiY1pjuTSCRpdVduyLTqgA6etyophzFDFmp9q7Nk2o1fQN92kftyrTpLi4PHVW/+T90fpYyY9
fYWlXnN9cWl8tj0NkJRF3Ari+lMV0WBrOF5ls89WdgPF/+bTFe+YK0w0DepIvd5ZHmpVSLVVH7lB
0fahRtIEV/6IsHJ6GQLTdDrlsUcjKGxwnMZAjPdlWUNuBmBcf5FdjlUYs0YC+018CmAThfqOXWrN
7JMfEj0r/ORjULbz5cRtu3n+F4tX1b6IPEdRvk8QQzwQxvV2n8/5avffs1nlRCtgDyIftTTQkgjm
IincNaibOdjwMoJ0i91HaOPwoWcNNFIgNd/aHsBvf3sxPNCNRrcXDFAwSMgLZaCU3oa7UwPfwKPL
nMtVk7/UmxHYWqEW4yHgEmfdCh3HTUm1oPaou+5rfrClkc5pq0isc3TKjnHP4m8F8SURjZJkiu2a
jGaeJVCYhz3sf2S4o5NIZESBPrw9NB6W3pODmU0m3d40fqWTxOaO8a/xK6ikmtCmp0YsnDb3JOlp
MBcFV89SBvE2/O5QqxD3oxqzfiJUNwQ2NOkUZ41t8VlDe2EBrkiY6ap++sarAyAGT0vD41j1EbHb
iTxjwCci912ithakRuHwU3BIfbqrzdmFlp2CTeV7EzSS4zjfWFMjXMZL7YLtt2NKAqGm3XZomjnb
dCSZfcChPA7gKbM1XciD0HCIM3puoMQxQ4D366psZ6vi0uDkh1mJegQ1TpS7tLluAV+PpdvffJlQ
uPzeyQmn8dQMpyqUgVKVC+/dqM//UOTEdPF7UCyAZVSC
`protect end_protected

