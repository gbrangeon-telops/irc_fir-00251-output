

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
BwHHaRYHij9TGTVh7NqyF6fPKvSJbz6zXpDQ9T0CSRjM0Tr3I2/EoB+qBgzPRFij4R1VpNLIhF/W
jnZk7ILw5g==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
EoffIvgX5Yh3KSkMHr6Fb+Y16CSwhqKyrZiel9vaFNUa3EtfX9ml680qKyH6k7Lt+GT7JeOZ8tsv
GeWg3Is5mnBMAsR5XkmKmU1Mf0hiU70CtdaVxbMu+l0K5NkyBzps5GWZFbpBi81xyWc3mZBrsdOP
SKFV3jiPDhzIXFusLNI=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
pC+fmAQpqkr0vqse1A8SFfJnAErWB2cTBoy5W2fu+Qfel2Cgg+f01SLqdiCqUwM3sdVOYKq280lw
0KlccFWeISj6EGy+UhrlckR4KPE0XJ2GFpTDwr6dIxS9OpYPDM1MXlxttLYJRqT3qA2yEzsidST6
0i31grVO6qNsjmpW2d7uByo9M65VEOheITjyvjEpcaFShH/Xo714T1rUj9u+HOahJ+Y/IZt5BXf5
ifgOOsFSC4Urhn+vw7WBdTykWaXAuPqSgZ+BAzkf1tn2a5qwxdC/nJyffVluJZjwqKsS2qOqxdcW
lV8I6VmHkVrsFF7Im+SIdtLtq6ajfsK+Fu41Qg==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
sjA1wOpImDpYBBRjnwY37zkJTSoQvS3OSqKSHwre5fBAKnkrgUJxozoTE8i2Z5d9g73A+Dh1Khan
8gYd3xbR7Bt78jJM+PFuUbVx7c2wSRcHOAp2KIXVLTpuc4ycdBn19YJhb2UIFhm80kkNGNgavUsF
mOqFyOQQiDU6WY7JVI8=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Yt106ecWVBUI4xOZZkRHweGkZD2nlI1jRN4H6Fzc3EkfIh+DLe1c/sY05LO26DhXbTC0r7f3V5kn
SKvkly14VHuR+p2mt2PXxY2kZUcL6SEF75Sdud7O3qeyYyxwzbLXhAk8rv8ESHYXdpJzGlAIPVhc
CV3MBlzutogOhAPHHcbRbukDx/ONHomfzueq+JuKHmbmSP3Sji52yPtcq4iLW/WcLghIBdR8EZ6j
UoWFDA94p9C7hEbP1WkZCFdBxukr8LSVfTsZyILoNCYLGaM4SAN+KSvY/r6FcDftOrSTK0VkVrNX
POMgLw4WpJ2xpIx+qCPH347wGbfYnUgOpgfHdQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 39232)
`protect data_block
ynUpLydV+00Z/oPi4ZxDPJcTWqUu8PCflaRCU7Ta9w0C+PT8ndflpdiJb9CFJ/Z+8qQKaGOKWxmA
3yiODs2MobCtPCKvopFx8eRmrgptXbeZ0uQg7RFtutZAseWRYR+WfXu6/4UzW31c9kYohoJT8j8f
OHYtTY3d1Gxoe+TkdwHg2ygX4KTKEZExt3+ePl96fFVuGNks0mAShx2BEWxqBrT4PkykIpN/BtcA
vJZ4JS2BJ7rFAZJKr3IQFMoCr4SfcjnlyRIRoPPhf0XJj7STapsTQQ5QQu3AITqsnZUQrdGItwpJ
ZiOaPqO5aXGYuhqLO199Fn+ugYXDR5iF3eBfRBQgkwd2xlG3DkraApkuW0akW3MywKnzDQ7g4MGM
p71TlTuMzgs+yTqKL514WltYM7wO2ZsBFGLV0Pg+1KABa5koVzZUgpE/B8uIoTgHqvrkqXURhW8u
tWn7oNhSydd0L6LWmwN92WNlC2uLuqPQZCY6U97qTzcM8ofqarPJV9spleRuwJ6LnTTB4M9Oi1l3
56LB7W5cjxETVRRsknG5/TQ81DJ/OKyCqFxWtNU89nhbIrRNiVrfJERLju+reeOV5TYYsDLLhuBK
FEwgEEUFmzzpMPv4KhXX2ok6/xGlqOAxBHKbC0YKHY5QBoUfb4q4pwwReyfZvtjo/EnD6AGc0D+N
zBtqUx4H9WcBztsNf4ubwzyDgwduhctYBV+mXbBFVjGyHnTuBvKfq0aS03U9vm7pL6oKIEwns0Rd
67knH+U+I5Wnb4ewDi2viZeus3kZpBTbMCR4OthYzuqUTK52h00eK+W74sikaNnpEvsTkYyKFS9s
YrMHcDkHmZ2mXMsa+FRvkZhhp9s9Wu5xzmR85BXPD7g4m858X5s5aHW+pYDin+Ojj01pv1LAZ3Qh
jpl+TZZuK07SWDCwTaLlEfPLtK4PqJcDobmm5O2z/sPxeGdQ2NR9MQWQwgJh0T4NVjj5ozy00ZTF
MYvxpWZtrkFy6t2x3nZIsyVYgyPdNm+UksXrMhglfNw2r62DU0jQDN5siPUNvlm9diup3hyBYbgo
exZoRAfjJaJbUacqTiYqhbFqud85NOovTVVPI69tge6UkBhQITNU0qNONqB0MMgOdYBc1aB+vODQ
9xZ8mpv1oO2QdexPoDjL9pyddTImXHjPrK3yBEqzaPneEcWvl+hJ0WTv1OKhjIiAX8pAVsL64nYb
dsKhWipOG5apc4W3PIKIEQ/RjzWeAq3JPwZbtztJ0Xm67QYTDicrpVWI6D3r/KOjSkzfnOluebhQ
JCPER6vWkQZQqs18cSHjyN1qg72Hu7e/LE49NwDLYoLPx2kpCOrOmWLu4uBQvVQw4022V9DVeSzl
hbB19+Nxqtx8d4sIq47blmZ/oHU1BTHyMpCD0VYa4PLzQZ10xlY4G6Wu0mNFijl5GV52l+qLxOQG
fHRpnJx31yp0tgnVckcUO8vXoMSOFR/TukyUJDx1hnllZtZNrG+TMxJpvMKpU668vcah4l36Ey1h
hSAtEG0hzpc+qZGcaE4o06OHRut6oIL2angR/uEkDzGloxwwjQK/in2zfWUXHQsvy4fWh2jRNXTb
DipU/FoC+GpUiD6gwmicslJ4jN5NcpH3mweDv3WPc6kabWX/peUrE8a9V5f9PxipT3T5pboebfJx
Vpcm6hk/4MZIeTHM8td/Hjt5a30s1lIhbetgejDFOj7TXyPVNuskKZWZoWrorC3H4sxO+KhaclQO
GvhyQuU+ZzwAlXHCnf/dRBzjBVuMHcmiQn9ezqtRMTZr0DDjhwhdII1I8pVEQyt8T97q6I7nn8VJ
8pBEZIRd0sU0LV9D4TKMR4lRmSeqQ6hq3TkJ6XNtyICYOprlH9repohmeWJB3HtmXaVH+m1Gq57a
pccPbRncACMVoq0akGb9WbsUNM41pdjTvLJ4Ce/FG69d6crtYerO83b/GOhK56cAZgdoBJFxpMr4
vk4464/3eVAnHlo21S11VmQVj2uwulRQEn/b0sC/o/xrlK1KpLlrVH6RzeREDzU4gRbxnBtZ0ieZ
e9Cj9EG6sMUVvdUl/MAsm9h2VLZeWebMAVNsR1Y0i21n8VgDA16W615xY8B5hPwubx0R6s9qjhng
ga1BtEeSRJ+1Zl9VFbaWhY90zKmFHp/U7eL7hAswWg7QyMK5qlpqbTSOp99Am6pc/qcfRFbTzLqZ
M6Krmn4okMYZCcCTIX61VAg3jMeIw3UuaIkarSh13NFLxI4/lSl6P9xkQ1qYug72Z/jjmImD3d/0
PuyMgEt88AVF0ziE1rPB+QnPH/aiSiQbptP+iP6C8lM1f3NnCH1/6hMdsCmptI+uWxEOZe46KElA
GT1oLRG1ji7IVoGglhCv0HNWVHgkOiOSR6M0ZXsNvAEryWmryQYHDB8gkHJBMJRFZFgjQjcIzh8V
wFfiwVK01bzOVhOVeKpxnyTEHvv6MACqoA9wXAmAl03SlYWtOYb6ULt1GeYljuYuDJK08akfmDgb
gInY/uAzaxb47luRxc+5umBYTaHATS+NKcXmD1OknCktpROI+sUrk2HbrVhd+NHaFPH3R8hkC5Bk
HExMDDhz4npdDZFH980sxZ/iTroM40Li8uFKjH0ArbkxcaajeYhddVUY2wB7o139+MIU3h3UFOFa
pOeofzwscQTYKC1RMe59xzF6EkTGft0kDoiQA8sN2hc1im+gvZfCcC9+cikbyaMGnpXpwsBMssKq
nj5PTNKmScJJJVZAa2vr3Lqh6XcUJQIQ3X1PFA7+VmxnLuY3E5G+C+GrYjOtibFR8kHjzXOy0sjD
L8/lk8+qk95TYcgufMCGTMqMkaw5+vLtylsAx8JvriGNca+vK4IRX0U9V7s+1edEQGbyek8JJOdJ
wuWr28jZKRQxI+uj8UlzDnddJ7d61MdYDx+mZd1tkzw0dBkvj/lBxgVqFJkPJzCFpRyv1q4ecBZG
RHybPGBs//gRTo9Vx0CKCJjpy02TboNfUeigFH7CW3OfvsyvAlwv3n3/5L/dLiiyAPsyce8jf6rR
0HUxQlRVD9l4hv30PQdaACLf+chs5KbgczrGkIlKCpdwT9aEiz3LMkGk85mlbwhUz16BYOUNLtwL
HhmKHasNOQmKRhAs1a7QmIVlZkQmGI0oPlhpm7wJe0Bt0KGRGOWmYydDajEar/TqzbX6S6O+d9n0
8Vg+ihTm7lXU0EJaSwwA9A3u39EH2djqNY+iyqxlJA3KipB0iFa5CqDRz/Og1HYDDf5TaMDEFg0n
IEE1bQas4RVPUJIXQYLv7dl7OoouoZ1Fxj64VlhjnddeLt5pcAPicMS4G9C7gGH+5WgEbyS0IDlb
Oe9D/51YksJ4JfW+hoWr2MU2Kg9FFe7x2n1slt8vRTB2455V/+bVJPJ+/FSzGGw15+o9o1JpXvLT
vkbdqzT4MzhuWnBNwIamXlRRX3/hOVWelXfNGrSaHaZV3FnkleIZyWLNevUPM0Kn6V4kKdN4otRt
WfL1WKIRc8yTz9LbQyU1lGTdSYNn9Kko7Tfsb1VodVlb9+m+ZDck9JoXoiHh0QgkPdOo6+9XFTFt
JHzMVq7zpWd3NdvFMwY5Xn48zxjS3WIMihZ7YIvQDEpoqYx6AUGra3pld9EfFjrbZQp04YbD2Xn8
N1ATJU7mqscooevjauEIBttE/I4K8qH3YZPbdSgwxS1ZPFaHpIl999hLQCHYhVlfmoI5qT7oQTjn
G8W5o4PlBCSzPoJ03KGkBWsfm5Nz5Ow33mCzSi0w9HxFSnLxfeFXAz/9GAlw0MBgo1L9RYuW/psh
vgPfpTjIGshZGnJoVM0b+vffGdgjiMHkSUd3q3Lxi5W4C5R9qkayFl22HqTym+v/QOcnVOV4tEMU
QW39NzD2ru+whFtlIx327qkHWbewX/ETZFP2+lNhLJTARXhPlBPCxrZlFqsWxZomDcH//17YkkEY
jFYFRfDE3K/WO7Tfw5mD54ombM4ypzozAQwb5N8ZjT5utkKADdWaFDYLnLnspIlyqzywAbu8oeqh
xh9in3eB82j4m66qi5MzN74L5eYHQB0zkWXxn8XZMoXDuI4dGa2DWTCJElPqn99E2jhp2jJ2JG2b
1RKnyqpT0+T/EbS0JHfGIKahok/d/Kr2YMsol3SljFArJwPxHFfBloZp64kk9UPafLDQ4s+biGTh
lmeqo0hYSCKm7meYwTX9o10jwaodLC4mtexpXYk2pUeS+qdc6lvCUIoxs8zbfMBOYrRlXn637Bj7
FjjVt1QQ2vdntBYde8DWPeJAZxqZD0Rud8fYTCQDBaoh9xidCeMnWziAHY4ZhUYKr4NEWWdbbn6O
qgmk1dwZb/0raA7qLuIvargA19ILBJm4xfXjTsIsMZjIoG9Y8fK8OoBTplWbgjVB8G88E0hKH/kx
Mk6AYIx1OOebkai6NsTE3BR4K2RNSTeb1++VECJAsc2AJoezSxcFehEt65w/7EgTX3+q9LM1gtJJ
sR8oSXXuiSum0qQglYsi0I+Li2Jfitan7DxPNaR9NgsZZJaJzLX3uEr9mOUPUm3s1pFCgByR/1eZ
8CDppzZIjrJOp/zXo46wbjVhapSuYflB9fL16/Z9N6tL60r/1weyqnsliZE0t25xXu7khRziMexZ
cVl/OIPXDSPG1uQf94vd6HfLoeVd3uVXEyjZ3LT8skaK1MA9l2w1XZ3KSUiCjelzaoENmSauuRtz
Rf7wC4RNuSXa7s2q1duc2h+JXplzwRBelFxNP1zAR0e2Xx8oGdZvwbGok8gwyyfH+f43DIfoVw0T
8oK22eZRiosOE0qWMfjA2nKqz0FkJplofdTZKmw3axeSAGIwanIFJwSql5iVzb+M5MxI80++M7Al
6rnWFOHaECNZETfg1hcBHQWrK3hsQ/M+fHSxOqnfJRcw/tbKp0CsNaePFtupwHjr1qh1aKXrqYAi
E2j19gNqaNInHGR/uol6UtV1Arb9d9X5+/wfhCFnWs4mlmczY6JqDvPAuoC29dt3wQAZWz8u0L23
pIvnE7mHj99V5UXAfqMd700iEWNGyCcSY0xzwYiJmD6jRh1pVwDoWsu9E2c65X63TeI1rcCs7t/U
ng9eMbfEUSHRDfbUnYFOjwC3DFa+EHLX+ZsAk6GsSQJEyGqrdJ+KWWKZVMI767lmmWuwvj5tAiHL
2HzMgE8tA1mpmOBLFcnsUj+EJZJjVY8Ez4xGStwm4yMqa7ukONtGqIWTtSTjKGSigfGmgN3Uy0KN
yHJK7cqd2Lpv9mewGLDn5LbhPWMdbbl94wmr5euoroEzdoDorfg9TdluJBXd6YihlYqIXdrtmvcI
Lyb6d7VAdhJpesZ7Qr7EmKEuPP545ALrh9yPU0+iiYdGsxrCcAvgf8Gnu6/gWkG8KLYj1zg+zQog
ZEcldQHoIndJ3X4jPUF4bxrMvFJpXLTZGmjmg0QkZjKW8LIwZMByJ1h/WhemKET0wwZYoDrblgZI
o1cfZMmQlHRPgGRqPmK+5ti/Cqd40uC1cKY0Q+K1mMUtXzEt0bW4zoSZikruFBBa9s/V7lBpHyA6
5Db7E5/RZMHqLPxdEgurH5lFkFNB5IpBjkI8QCERB+ioQOTMAxm1dycyl1E7J0CYoWtL7EuUt96H
1IH0meSX+k5gloxN/Xxj4VgKkqmmQv0RskRqq8hG67vrSXlANFbzzK5BzEHqVln+VjCacanOz0ir
3ugvswbPmXExoz2ByiDh+uE3XwxtKVaDklyHDob2+p4dLYi8YtaPgnybubrlfc3lEJsPTu7IUD7g
9Tp17IFYONilyYkGpdO9Rz6C/xSI3tG6dzrKMQ4X94Q4xV0JicybagmOCRV6Ji8+KuYirVzYmGz5
VQjaE06ITm2NPs0mmaeTWD5W67rngP/cFrnQu2uam5Xf3ol1fJ2HOlVjkVOEorzIv5gDu2Lo3yOU
G9EHlxCV8aC0hmEZJ1QgxrCGIEDfMFsERweWMzL2MrSFsVt+sjsy/fOVDrzI24JFywJ6Mx3eLFOK
JUU9CREAzx9Ev9nIBjNsQIrJGe3WM+HrGJMxtlQFeVmDpb7U9Rez+vKtQxDJnwwxW69EsDDn0asV
18yUXbQEK1uRO3f0Hs4f/o9LtOZHEG8b5O3FLdpqPkLjJVC2BGHvh136sZ7Uaq25z5zEGEt8LEbK
2qQ7iZ+bT1KK7THBsiPsiH7kairdOKTYJ3rf0qjTSPGtuQN32VNK3M/vB1ii7PMp//g9TpqUaSBr
nU4pN/3/wJTvEJZExMpZ8Y+2qKWNyNNrGr64Huj2CDx9MMeHYSwaNsS7jDA5Iw6DM/LdWU2MzoqQ
RWBsYefjVcHA7KWep4/xepMy6Cmt3CicHxaWYBWKlBl1QZBi2pME4/9GnRv4YAPyU7TnoerXdYg7
V8eu5Ry9+7OFs+2lk+cnJb1oKrTqHOZKUlQMjqZEO2Q0mDc7hKvP5keg6yOY967Xf658idjIHod+
i/nJIs4fXya0Nog74kBHdNTBmPAAv1kZNHhfrhkQXCFGCV4p0ToP+BSKSR0Ybimba0BPOVakMKi+
Erpf3xu6DHnrCDxDpu5mtzRhHz59strgWBcFfUjJVjn2vzSEdmFRiat3BJoCmqZOCgOy1m07UXKg
Bmm4FX5h7mGfWTGApnzYy+BdbU44bCd1binDQTXJHPIAnMY+EruzZdMwuN+rmmcXOgNK61U9kmK6
MIjpFAinXAEmtnVyG/x16xQmLa0GbpqkGHEC5HH88eMG4LMxieA0mCJOhzyWg8PZIqMMYNGm4ibF
CtLokl+lmyzx/jnR9aDA1pibZesgeNCmxE0V/VgSMVYMm8iLPQub3eoBpPhTwzob6GPf50VsWIjX
xgKsk0L1x/4cwytL6TM90AIHP/0daE9COqm7Fhqatp7LJ+cuyyNA8UJYWE69+J0snLMrARDP1Y9B
vIPba2S3sFUzYoZtpZ0aHPj3/Y4vTdwHgqwt5oWT3HamtLiSYINGT8qEJIqcGdLL8MfWoNE2n+AU
8OtO5mrlUfjOVOcweYuMh+2Wy1x951Uria5H3DKUfiI4DLQwL77vIS0sS5YALSk2NX+q5g402aUB
uyJgemvo7jYHGPqliKU2L4w+QqhtUiciVwU9n6YyMqkSqZXE4RvuBdV670+vtK91z6MQqyPVgHkr
QjndjAueKcAmZXziS4GQI0J5dG+j5hmrK7rUedIAhRB8HYBU2rNQT5kN+uBGV48Nv88m6ahKK0bE
l9/9xZ+AUDQz5hCYbQg+ZKiAYI9C+VVnSj4xJdU72vPlBIvh8Zg0yr7KEK4NwEX0NlZDg1+TYCFd
6c97/ZzeVv6vpzckWADM1kgLNNoDp1/bjDe1YVvHrFk7I3mpScVuXT/jnm7jX8ks16/MOpAloLT1
bwqNwqpq9yKrcJ4gst/AGAddAu7wShR+bFPjHRs4yHTjNdF1nlnbP+YcGNVkHpEzUfP8aMj1p+2p
5OQN2lwiN7FXKgX+mZ5gUjWXjpBzyKvjosh7jpbyKN46l6Rqp0Wg7WaPUXavAtke+6xbH1VXuXNn
W1kz7lHoiizJ0YWPGVkBZQ4u39Lt9cI0d8L4Uzmkj/UVoIM2kEbXDpt7XZ4a1WWB4+Y53vgJzZO5
CiqC0VjF9BHg/j5BUFwyTBDT9ExN6d46svAu8QBAbP0xTYYnvgYogo38Z3kPo3jLP5OwF792Q3vG
5Bnp5CPPF6F6MSF75oOuF5XdYhG/TceEjWvDKjQ8pQQ2+3BboJnR5NCMFdTJu9Hy6mhNd45fhq5x
hlaDugCytfSsDgz1sADicYXbrxAsWAT73ACT2qeR8mTv+IBQMBQq0JW6CLU7mjtptZs+OJxogmN4
OFfeETnXVPGiSPLMkVqN8g2lNmoSEyQOTH3i9nLPGecHXF2g1kp8TymCulbnzqgkjqOt+g1ZL0gc
9IGjLb+Nv5+omfQ0/Y1+3jwQyIvyIkjiv8hVfix0Mk/yDwC9sljGKt27NqpPQsgUARsAuRyuCX/9
n8RK22bWQZ2YBMX6IukH69vijYErlECyQvUDYFsWJzMsIqstkCW16/1ejqb+L4I9e7B2rjcmhrZc
ggMmdwxauQ385lt6HEQrR/+9k3Ph0smrXh4Wj8Mnh/MXUfCOcBbhOC8DlxJ/zopPC2wcD19h7XnR
ow953zH0motO69+Aw7RZpTEXG7rWe8wpv3FIYl38sBzvSMcwtytU/NCnFFmieUIOVC7I/mdFxRVI
5PvnsVD3aP0WSntOAKNAPywUj/rwD/6+HRn5fSNNxchPexmx3gi2rhphKcLI5HzmeB5elR2+dOqP
29bFkBWZ90vTyI9SvwP54yPec2ufm4mk5OTsKAlAt/gnV4kdb/62j1x8KjQ7g6PXjNA+4SowXgN7
MOLv9hXQLKwqJXLC4dvV5VuNazhklO6Je2pdp6VzGdHVxX+OJ9r0+SdbzhRbh4038wFRL8ttC6kx
3CbYRSZmub+um/9sWfkppyjn70jMvNoyDootoVjR4nPCS2m/yd8reaJkThyKOZ0X4y+pHkcUdrJD
hU46TrzNXYkQJM6gYnAETcVSy1bQpuO2LUhdudKh2rHl4kDtBQXemD2smosta7p3HORjDisyhoe+
QcyDDG7nu5zOokpcw2HfevAR0Lpa6qKQcElS1ueE2ICl/NlUK6NZaxqVhu0EsVKEoj8BS8D/XBST
3GWOp7TxUqD9W++jnDSxRVDeyMfVuP1dEjS8IBteCRHXegrpxmMWV3YoSA3lWHCiT5P7Tj91bWBe
eshA+6+5fTKbuKzO2lPXueGUO4977FsucF2dXqf8pKmGJHisDjjikcSwocYFIACHQO63iryztC0v
sQejyHrvtq6cmZRMVU8WbmbanKf1/Cg+0mUf235vY/gsyfNYOh00iDWg6KsT3dybxHZ4F0hrEhiV
49VOR+JUVYrVo9GOqsnRqjgTR/iq3A4U70xYUgc7ehUfG0+h2bQEIZLDhp9WJ6YTGOghCMm7VLNF
qyYxvLXtP0dY11R1Nzo1UQa3UP/rQqSjZf2Ed4Oya4DxchIT6ikkMR0FEVNzAWmzCYqlVMv0irjk
6DsvhNXrkYDKBCM5029cVAdfQR5lfvCu7jAmTLx6SyNOyZb2oef9YDZ6IJ8KW88SFi9GRtpCUV+/
wEHpU8jvOxWCSKMsBL6J5JRwV7GFRYH0cibHM2Oach9/yRbyjCkR7EaSQ4Ro5qW7XzDH/4Jx/55O
an1q8X/+jIZckSFJehXCiK/mAfpeH4a/qDAeTp6NwpXZ64sVt9tkGQOFARi6QFaOTkZCV5U7EQyY
Qc1kp5v8MhjpVYnnVln8evm3nzGckSNRy059pJ9d+4qErpzea3W2JQg5Lb/vpPjxH6oSPeTLPLZE
wmB1bYwg3+hZOGW/Y0nHX2jxunidJnqZ5IArdGnCTCm9GvwN/We1cmOGmwB046iT6XO2ozo5+Gg7
Dx5Oe5QtBHyZG1cFRYm25GAVKJo3IBQR3iyCk8U3Lb3BR6fiXq36lLmioCJsMFVQOei6uxUu0G6X
PkV1o9M2haHQTG4lGyNDPP7WU9O1Ee9yjK945kKnu7JmpiHkIlzzvGgziW9XvK+SEGOwLdDno6Mm
pl8Wl7HSPeTLHhmAOrq74YSvOnEb1IY60i+ujKjfkKjV6HWfO8KQQOSRrbLIrXXlbe5LeVYzARQd
1b3QyPtd48MVrTpkkyZPwEaCZeOIDr/zGvYwVr3JmnnjHv9K/1NIxF9Fte/bGxgIGdsKWe2chCXq
YnpC9lIKKSFTAEKlsgvWmly2sF6sKCTuyl3vUhE5xHyQ/iqgN5sdStwHy+ErUmC+85Tc9DW7eZN5
TLlgG2hBd1T+D3WpplUB1wSkJZsF9QPt1alWvy7XZ/x+4iLy0uRtbg9JtOnXqeDaB3vKpKf8USeQ
H147cLewUqlxPrLU1Mcc9p267OWAFL/OiVIdym7eF09xlt0ENYS2cjtTpNUaCNdQO5xNI7A3aWx9
Zljzj8qdbYHyGE9WRSBwo8L1oP42Cs+nHqOD5aRJsc0GRStKkjkT0sgSTnydVC4QnJpsCaOk2tPa
9x891Gyww1tEfpIpCBIw59fJu1xKVUDsI3diC3wDR3Iqk8rGEJTy9H2vYNS8mgDchxmE7+1kKRbZ
JtEXFxtzqvAg0owLhG/kKFcLUQk8lMZB3f0X1Z36B7mH79YHf7J/g1SJEpUalg+1AYbsldogbmvx
bTh+W9WgOkYH87FNBwqrWbl+GVTXLM6X8MOxdG/eUiDLgxt/d4pFFyha4nRuJBa306MGwRc+p9rP
yPXJth92Xrqyoue7o2HA0iCTppEffIk2WJJy4PfZ4fadO3J7ztXN+3U9JF9P6ftajbm/g6Mh+Tg2
3dV0brc/WQZqBV50L3CskDXCcCR1CW8YWYWaIUj8Mk/r/rh+k624pOcMA7yNIpVbBxP6BNTsohe7
z6I1HiUbxe09HJP7hK5FnENq6GGZ72Fv2i3gy3coIbFajUA+xMYZ44xFF5/eQ6qhSstLpfMTOG9n
ZJA9lyoQzYPpiVZ2gZoBmvoLPVbGCIxTuI5K1Yg97s/LbsDr+l45494dfKm6iPtt1n2byviF6c9J
lxFUT5RbuYhfA6m5i087asKuc5CbO5KW1g6SbR6tUPMKLeAT0S+2HKqbe8gB4yH6nrAds2J390Ta
B17uK12CJQ4mpnQUxqVNQsKRTetlH8sM84caDcAA0btQUsZhZ814HmiCa92xvmqaBIlHlDLTi12k
RaQvg/kqnukeoJNhFSVZ+3d9Ypj3roCwbeRAvfCCQzrf6Gt+FfaOJCF5YCKBKcPHGpkbcikphnTe
5UAcKUoFwbOONkWzVBMjIfNeHK/g21CxnM57CqJzVzt2PlBbucu58dHFGyghUa/ZARJ68znRr6Xy
0X/u3axPO5XFPv0jrzIPWUH6Oz9gDUVcieSMEhm0TWNXm/fSEOT9K8fyk5fo+6PhVNuA9XkLLpAG
Wsf7Ktp8cFOyvntQB1Nu6yCbrEKk0vWC4QVKfuRmmYEjq/jf8SjFUlPqJCqnEanWnOIjgFICdTP2
0z4+3yEv1m67MzpDFtoDobMEZMQQrPFZyEQQoCe7tAm0n5zIXjlD/msIkRjtY1WSyHYOs1Dl3JZJ
UKWXhJnuoWDRJDCJmc6FJ263xlp0ADhQytPxwUpADB576d0TrRsMqAxQGEqryCKgmNBO/wpNHb/4
DPwh51mF4aPdhdJBSuoD6Kc8Hbwo6f1UX1aJKaVnAnzFJJ/YQcXlKtkICZLEaJ0y3+l3fKb9oJS5
gvt/TXmgWZVt9Gysg+M3QAKY7+yEkJzQe8/TBgPJKyWUQYd4NQIJOWnOSR/mpAysoh1b9EEFTmVL
jN0ci/c6a7yh872v/lsrQxZa4FfxtWtdnFPFrSBek4WaK4qaJYxnd9I8HsMTemnJ+WYVaczhnxLK
MDQyBJS8Y73Cq3QIGqTlpiJmmezsf4kiNtSK2IwB6j+cC/Tlk3phBB2iaoWVqjD367rJ+5WwmGQf
r8Ci33RQWWRkAW0TK5uIGFwobMAExuCs/XSXXZnKZWqtBuGLc6Y+wX/mXdgdBVo1wJ1gBeIt6sjN
ALUBzGg5DfiwZW1f3e0B4Eg46xvv3jvp2zGlkVS9AtEVgx4SDnfGVQOMWoBTYZ4KfDqsnCDMdwpp
8LUOWXkMvhWMh3iY94EyRJDKsIhnUO966HJTBa6uP2ZtDhXeXJFVhu5eusi1SUV0mwuhksL86V9J
AxdDr80NYweuqsRdnAv9UVtpo/TtlUCVA5TzAp2Y3x8tf6fslRxqXV9T4pjHCz0r1Ces9C/uNq69
6UBovxZfBVGAmJdzD8ubBsc5R/v28Og5GxLOtluI+/bKVawHBUh62ubLu/sJvG/ZKi3eJTOyjXJ0
fzAb+JaUxLgCrSlcXduiJBpwodWkQN3slS77Flmchufsp6+3/YtR7iG7Y9hDOpCOcB+wFgsWQeLV
9EUJVY8oRRirvcnW7W2NbxBKXOzoUCgcF1KNGhGe4KNE9cyOkeuqtKqHM0901PHSsW+d+sqDwKLL
fI3KVuuUhkqbYHP66PFU/2vFux+V78+w6TawTqgPnB2jlJ/F7dPb/SN1NGJ2cNZnWRutMzEG0Blw
fx//JQfu7Nhk8vpo+DMjIXCT5/W0Z97XxPanr2d6GD9LWPDRC5iOSEHETfNdTVc7WN3+sSgYXmni
ddJjEtMRRsVXb6rms71RPeMVeOZ+Rd0x0/jT55/Ccg01egTmben08QeopcFL+P2kKHgbiOymW+J2
Rzq6Na6w2xDvswGrlR4uY4P0RL4+XdpRcXpDoNGekKoNd7S1Z8JFu6dfVLXhwgmBj3Ys2m+/Irw3
g+pDAQgjdTkOJhMTJBe2jU9hI4XNBcoUzfpIdn6gA73XwMWmq4qFYJok+9ch7U1ZO31Ud4GoXGoj
lvlhcu2GLhXdPpPpuBV6DAd8LQu9hwYDRDdBl8ioTz5ZwpoUyh/TKuPBfa+LRFO6TdGh7YSYz9Z1
qIGbMtt3NjDNmA0YA7GpjiQaFegklF8zhH2p2B6xkCFSdUZnzf+ARJyAkmwa7KmcMKMSb3B9m2k9
0V1wzI6TRXTDC3TpN5PjF4J3bXG5RwBHyGKYCbdp7FB0PJ139yD1+drHGtxzYJIG+BH2A7Lo5VBX
6tFpNU/IsRrOPzwzMhVvANfNJGGTa+h1EgvE2C0RlDkVR9VYPqoRF90AWiEUqFjojs/pfwp7Wc4+
mjLcWY7mZ+7X6lFxKSz2goZXiVVL5YOjBB3tWteoUbg92AK7QzxWKY37W7D8FBUwQGJ8EjKeNJFZ
VrMZB7DeHvTkEJd79mITWEkl1dKtKlcQswXlUQf3lA7AYtkoC1FZWarXhm2dRNSETiL4SBmXqflV
N5hRAiXJxiF5R3FC5tA4oc3zYbUUSs0wt59j7q8G93xeMfMpCA4H69H46pXgUSVuQc28JjSOExdc
vI2tZJ76EkWaTKATmJ1XOoMtWLBnNZV5wGLMJ4/6yaz7TUYiYoR+k1TT2R6Z1CpKRBBGBuXt6uaC
oWEbvJLTHOvAPkephrTgfQe/FKz0oFeF8Xyt6pqrWrUbj/sEmr7dAo2HircTnbxK4C/YapyeYfyH
TSKfaU51I1cHBhJFLiBmBfTvkeXR+kfaYuhP0oifrW3kBdE/t31RgYm+VsT5G41retFoVmmk4UvI
cHBVWpoFBFcdo66e30NlmUGPaDHae1gtaT89Bk1iOTnyquNzOCOQE9K0dhc3S5NaIYwaXlQQH2Ff
hE2gamVB9a6dYFQer0M+pg6ikTqHIRv/Z7rtI8nJeVvVMFevnkr3s53t3Tt0BrW+mTKuCgVTPBef
2Oq1QfKKHE/5NAAHPL1GLu4bJTJ/vg2XwiT3t2yID6jpwM7TRalCH2FVuxGt+nwuoxmNc0pV84Zh
MprzqXND9pXH30XHmnQfQ16+oHpJb20UaPUqwORJMH86Svae5R5CM3skb+2DeRI5rSkAWS85XFu6
3Q1xwrtNFADF60h7E/ZeIyxgqCsYwUTW/sKb2nDotPlXqaeTTGr5ouvKPjgNui0fU04oe+0qDz4v
NmaZV8iaPW33wgKjhcOr1OFGKflgyPu5rdf3uJLBpQjrK1D7sjrY1K7vrOGnYshMYWoRsUL2zub8
wu/bLIjxlRTmZWd8oifAbhqnSx5fL7YVnZ04OnrASN3KyyR2UFoM0BHngoJHZfBPwwZ3wVSbxtg5
w/v5eHBUNSTyaHMOpdi/bFkul4XGdffc9Y4TTIS59YEAccD3h3gUz4Barr/hMua3DpD/pe1OYX2q
JHI0jiDgPQncQzXc0fmTUJMr+uflHgRSFKvoRAC6vwUZeh+QfUQ9JV9afUqTgUG7oznrpWpvVIan
ILIJ9lbBuIBKb63/5vqyvtFkalqR8veAIE6WOpC5yGOGqq5UfpwHvq3y9187cEbcCbYJ2rsbBfoI
uzECnMSNmi5sx6WmUM4D2nSy7nI3MTo57W0o5//lCaVp3aOlPTH2OIHsRsiUAcL+KzBq945/Gmyx
uLBXcZXmVH/k1ncbYAQGkBQZdgFo4m3h2HMl+gvVn+1zrsQVqqz0Al8lVhzmB6XSBkJl9gscLET8
aGsZqPhI5LKXcbLIIxFPfRsDwh8RrOghQ7UBzn18upG9yWJgUFcCAislWGyVjISXc2SCcsxVuO1m
fmDp8EzgaXSPglP8ZkDOlBE02hY+Pw9BijjKiQEDFUeox3iuQNCZJy4PnAFh9gJAAglApRNFaa7i
Kzs38Wor7Z+Tid0O6KGvk0vWLifDdFV4O1Xy8lSQfnZWtzrN6ue2Q/vwlkw7ZC4qv1wtbj4FGQ+e
n/wGr4AxoI3kni0oDaXq+woBKMfB65Q52n3m0RU1A9R6mLlJYom9+igmpEC9XgfOygWtIQlSBJhl
Rojtoi3TOA8V6C9nxYRjYXg/t2NaOUnm/Z3FlaMeH7Vu82Q4RyTS9o1P0xwDTcPwyoVjBVgySAaR
j27CWwZDcuvto6mQVtQQG94NdEx4fbGV1Lh1iU9hMnaU8qK5ONCHdB2aIccgVJaHzODStxFsHTCu
pcyZXFA/lPylrW1V5qs4sXuJqTL9pWhRN/HM3hMst0XEFCz078KpHYgRpjsO8bzDY/aDSqoNE57n
aJO4xBEIY4rDvNl1UPF7Nse1ICT6jsYk35LN00PVF7/yQp3g8Kz4SkK2vZOB6Mrdr3yFMHjlwH5w
EBJMfuSGCiVVKdh/7gwh649AYc9NNPWWAoq52fE5nsoqki6kx/ywcNq591aZuZT/V9rYSfnEQ/pm
Fcd3Hw+60JGQXsI0I+FB393f+qPKc6oCRyN0AIXKNW/ggg6U/+rql3eHvtfNClvaOB5zlgYmNSJq
yZB+W4RoIw8oECiSzdtEw+EYgntKKOZeutSUski9dPArARpAZps8SKRJAMqvSCJvDENyeH1ckjsp
JkLgHH3MuCuTTQPgTh7CMbRCn9fYPL+Mbs0ckVWBXIP6g26SmP9XuR9mTkv44SbNojGXJeDK8XX4
0cEVN0ACs2GlF/CIjZrMHvAmYsL4gZPwV3fstH0CKpIG8npzZP70w9pqNuCMDsE3tkMezvK0J6/r
ezwmBdPy7gQmS5HnX9idERrp2MAhcPqkMUiSf7Eup41xPWKzoH9Ag/Ip86IJu7+YIEZP7qR3ZXx+
XEMn0oYr1dnbendbb6dQSpJAERC37nuCQ5rf2zh+hGjZXEVyNE4KhsZ0DEfGy/k4FuAAuQfv8d0o
LGjOvLfmW/90wRB+wsf0mkny8JJj2b60rb5wd3iI8vB7MYP1N/v5rlMmReB8MqUluQAUk18pQptK
YKLLXRVqHBUoi7lW6ar5xbjVrysUnBuMh4UyrMQcpBhNCkVw5/irG5A7/y97sbrUv4gYzh/RM+sh
EbOG8X54tRLtlGRd74/VNFQv4Gimkf3dHw/zziXhDXRenUCx9OoNZT42Eo4e4pW6QCht+t2/l8Ge
ygBMze7af6lfh9j/tLFAoWcIW7PJk9CpKue+cCZJV3CaXRzyNJU+THq8z3ot5a9qIoFPzXC5+uwY
Y4L0SJAbgOw/wQC8ENqErjurfwVo6JKG32So3P84NMSn9cqNH7JOzsGr9sYls8GGYqXXaosGEfGC
oNYEe6KKIxBJmSf0MkonlgIw9ddOwN2O+YK3MXhI3Qqo56gssoOE/XyySPrTlfPYhks/0TNzrCno
sz6n8SlzOhuUj+dw6mIBHcDIwRznkKhKXE/NmvXLcQOKuNoeU+Eq8H+7nFdC8yF503Rq6SV9Knyg
UDgSJIWONy53h737SsGSdvcH5Jj+qFJrHtlOwFDNrvT3XMQFV0YFMPwXC/NXhHCpz8624iGTXqVm
NWbIEvdKBX+KRaVtjjBFeiHD+iFgv4yOJTUaRkbDhSYzyXiAqxcPf2hv+I0d6U8g/E25pLqT2lJI
55sy5Qs8iq9VjlSAE/xVMGxCqcGNhsiZxPpwfxLx8Adj3HSuCM74YLUdjmyb1POiRjZUnzvSlTM1
cezEFSS23S4TTRKIRC1j1aY5kaENiCFgTqcsF+R9nvoiJbP164JgJu59zoR9mzoaEtfLoK1CTbIk
aVX5rDzGjIGL8PH+OLF1afJtky7qAUSv6IVE9D3OjcOkZ5KerrzavjnBhd93EWuFotQoiK3XDI82
yZHTBzI+lX5vOtZxu/nr4P73wEpBhLCT4OiFGtFa6SVHjkOl7dBx5D3vfEEAEbBVWVsamg85iCsY
jX8H3YdmrB9YUnBuviKkLLy5KMt7R/YYcMMHaVe2Kcw8QKpKL5gpNXTEJXCybVASK2hMmX3+cdG0
1hAzmZDRUUNpe3TvbDQvCA4ivqTTk7EFiWdIUyNXA8gtMcCydWoZ5z8n/bNRTfWPmWficX/hS8Uc
DMNlTyj0fpeJhKYACYmISl4+4ZztxCUGOCuXjhouGaKlipSemI8xcw/DyFxS9tsjeUMlvsxrsYUX
CZMHOAPZcSoEg2Ql28Bs92jJgHq2X34gLcfnJ3gDXUFY1mipsIU4QsXlg3WZQMzRZxSyaiRXFdxR
YeKY2LSKWIMml1EhzIz/KNjOk934JtheNdeWYTPH8Y7lMrL73QR0jpgQlBeiQtGUA1i3fK6/1nHW
zodr7E4k8sMGhY6p2o6JVyCjsNVIRGNNCBJJw/T32b6LxPXPxS/nLA3D7cQFv/pWUlb6s8AKNk9R
M1c1HaD22cs6u0tSkOioaYRuY36B447ZBkiqqdFKY7w0Ts3WR5ca3PsgQ+qRe0opbTTJMvTbPvae
9YDEMJALwqI5WAd2xQOvxh0fbeE2OsSDsqfAd6zLIg/PUUX0eoAD2uVsK0es19mi/NqpvA2kx6sI
5t75e+P3zvvPY4sNjMjgz/0m8emS0w5ZOe6iDHDeQGRRXEQM5ZumeFoRBzCUWIkclixNs2Nxdgv0
q+7in1pWjuumI4pRemfbHXy9ERLeHxSw37crvOE/ARneLXT6PWNhxnOXppvHxaJJWByQAG7+Cz+5
2wGaTLKj9o6c6tadhogZnv6uxnqg3qeZAXiT2LShfkxfmtME6Ogz6RNixJTJm02lLpRpYDhj7Pms
ynX6bN6oLJZhSuiVLDyf8Y3jVfAB1GignjXvRRyx7pYCMGj6OO+BaA4qtFoFrmSezP1ls5mxn4Wm
2jFc2dxpkNQKmSkMkzyxYPmtd6Y9YLY/t146gG0k19ELQf4ItVXnjPPQTwLNZmj9KIqLt10ys0v/
yGtlTvMHKb1PIEGIYrOzl0EjBGtkzacdCjuAcaM/i2jX+6OLrv2Kn5qhtJzPGOM+dwtqdylbRjAs
SAQI+7oq4rquY6nmUEJG2lShAM2X4EhUatMyqBA4v4EDZ4ISbMJzk+TXkFRE9kpkOyyVD66sJa0d
x8ugARM69w9KtrKpfHzHN2lrS508SDbUqgYjQqz/UQXqMVmM38SJ6hijZy8hskBICSBSkDnPE/BE
4fGK2xK8X/Hp2R+ZjIvBLtMGcTZJRIHJTg4dmxNaqvMgNIfRDPnsV/e+4jxchx2GnzZtKZHqfg8e
2xdncoiaXHNZClz0fw0HvoNBJzWXK4LYawpSL7XIN3jHOXuCPaA9fQ6rfWG/DVeOR7qpQ0H6TS6R
cjzu6NrcR50AYpZG15KSeKqST48G8nI9yO/aWhwvHaa7obLY+35LgFKcbmpVii8bwRrjoJlsxOPr
tMV76AKvsuFIfp8dkUz8t3JibdHqPAb9qujdK+gTz21e1ZTD/5wb3znnX4TkET+RGU44MR8BegP2
H5JmYOfXUHi+ldvYPXLT3P3d0e2sZjpjhlXJc7bBsH7ib1LuHLZA/lHyp5hDycQCweOZXYaOKUO4
lD1JDU/9isiODJKSfInBcKKp3/HOm6h0nQY52cW4tf/Hn07rmgA3fo/idumnqoN1FIr8ysSDEt47
TjheEYWILZD8j8EpkF9sLNXM315aCg/ILpyYGtBodmyxkYUIfgONqkBjF684KrQyfQ0YGpZJWgCj
HVYUHCBF1mLzKSVZdqINukLQOxr5woCSTHDPvu3LSG+fS7ZIpq1X88Krl8J/uXN1ulJczJD7Bf3g
gF3V/pYXCFhfmtBNG/6WrjJZ0yULDNT7WXCcPH0SXVoh2hVReb9OsHclDyxbenrKmZcNkVOwwuN+
VNn3SqBfHRZeAwuCTSOQ5WP+QlIrIf4Io+NVz6YrzCeOfoibKQMNg34Yn8xWjVPGzUCX5nas7JAD
OpppvXGtysDsPNXIfePgf2hi6nczOmZbTzhWeN6qVOzCDWeTY9go34Kj0bNlgxENpsA7Phn2yaLy
DD6dTYLywPHSnND93ujgn9ZnNyxAhOXUC7pKmYDgxE84UiOFeUX0e86g9SkPgzQvo9F44krzxxvc
jx/8oFaL5YBFhyZ/dCDr23j2l7gm7Ltd9+DaF2VvUDdRUcUdgEZPGT+gV6S4MeJwjbfk3XanwQoi
aW7sKMr5OsgTwCIsGbz0rB+PN+/+L0bbnDt+kMAZ64hXRbUp7Ce/XGPCNu1omCk9sByfsiIp5PCf
3ZIIrLAzGEmP5g0q1QT46uKLA8fZZV2Oi+JMu5cQvua+8VbAHyJABrAZwcamoZ8eSNNz1/PpypW6
WF93nx8Q2xQmdXDYHY+ZmlG18y+du6JYp/KF/QHkW/6tRQc2qAvxMvIOB+fzTkTEYpqdlYK54izf
lB+WVyf9KOVWgTgluTympUP1DpkTDvNnWB0XWgSSlA49xxtQOt4xdj0XKJRCQ5Er8Z/0DaCl/X95
cBW0SWymRsO0EQMuPNK0gybsrBy16HYHHAJFLhlRTv5wQ/D6xeJBTz4riPx4IewpskzVtsz4K9mj
WYej0IMgUtFvUKlitoxF3iN6nS+x7V7VKMJug+gb5125TEEP75p/4h6TiiJClBMxROfcOSyxRe62
Rtcu12zhRnzTFHVGjytdPUFr5rkJ5kGFNfaHrtidrs0c8P87lUWTgW78F+k8yNgu/OAWeZFoI/qT
9Z7qj51hLiQPYhHcBXDg7UUhJF5n1XV6cw5Ktw/zi+msDl8+UT3piFwYNAOiuVbB/EkfnIklSNON
sTqwG/tqJzDkIE7keomK9B4qxAePR4w4seB+MgA48lM/BM82j1DMFQ3dpLgVpAL6Kdruoa5FQwIH
HRlkujGodlR+G9hr2nYFrW4RDQSm3LhNV8D1ArrlsbqZUSVPzhJEFf3lt+llp7HM8KO8eIGcNAY5
UTUAkxf60h+MWQ2vbE3GGr18NyCVwzBqz0H2rUHOKSp3a4C+CujyEvblIyjLULOGYGUTbYcZazXa
b+E4prawpT+2CvKSsQNHnFBBrYHDnHuj8ij2okbXOcoGzhtsmwhdtk6MFAEeprpu6PBbsBXDjDUN
wepCd0Yzj0KOH2kkrdXRMCmAfPsSzWRHI2Im3xbSzjJE6Eiru51e1z6XzdDFPvLb9YyoRxkf+7xQ
/R8ACMXDCXSAnM9cpRuyo/Uah7jY27pK63wDCj2ZKazNG1QnN7owB9CjveD72vw/upeUa6CIQlhN
eY+8xXqWO+FUtUKFOmhdshsy8pqfoepHMKExd8CVSoYQygwTXTIEQVLAuUmafgr7oum5+/+R6z9d
ULK8eaLbKtPhdXkcrzJkiQoLWTz5FWZxK0NUVuJGEMyjCP81AYxPrU/3edqBRJgPSwL37pQbgD3V
PV7QPG+QWPRWzO4sgZDynm7W/S8lSo3FCX0uUWY01XPg1Sl25rhSNuQeLh8OOP8vPguvKG+q6zG4
/CzrTFset6jZvXkVslXf3uaF0dIiQsG7Od+zldi9DEWU4hGeITgYC4ogHuqc2/0amZa2huaN5MZQ
M5H5oL4tgzOa/z/ezZgTWmTruWrEpmqXYZ3TcuQskPj/Rzy7W4bgfjKuSAkEDtbFAbTrV5PtLmeo
M/XMiPHlmP1NrUn9mZ9bhoPNZ1xi8bb50sxa+jTzA92131XEdcyA0+rDmBSXq2r0KDU7pSeU/Xfg
UIA/TptUvTzz3iOXiCkYJNKkFQiHjVID8Q9p8loFTytnBUqEoIOVJOoVAfvPyg2DlOGAlRq8WY7Z
22pRx0mTzyf3E87KwVmJoVTn3eGHIXeQhMfkviLyBNsk3Etq+x1KPA1KCmV0Z8wPHtGGlbw3fRty
e8kL1iCofmfxu0uap6Q4EVuaPorAnu4zPnGRuPubcWUIfejmUBYX8TaM82EGhfsb6xwYjUVWEyKm
MbqG6NqVenr2xoA2KwJyoNSJedcfJNuUXn4dflAjXOzYid2O5OaxWcnpwCTrEU+Xuv+Zx3VpxOob
1x486tGBMY/vmVC50QzRTP1zTzGHETOX02gL+aXywYY5/hDSi3PdtbxhXzmdSUGW4MH0qpL3tIGx
oraML7AYJnFLLXozls4gzqgOvcykYS2MeIGTFQqQdXXO5qf7woVsx1hswTrgbHeCu/LUKXqD4p1o
OVz7noPuw6HkvbqQuGtmNYVKuVgq3OF5Ife3t2qH6bmKwhIA+c/CDjGjTptCCg8y4IW3kX7FhnKE
oSA85DxkmcUDwEA4FW/VKLzi8wq72CUwVmTFqnMw2A2XJJ9xcdDqulV73vwBhj8kNygAxlsHPKX8
iF9VCa6ZaErFw7hNaePAWVjWted6IURk3lYHwdepE785BePYDiF0pAVQFfgjFSSKmeNRAa+KIPMc
OLTAFdfJCroqo+GL81sdLaqIMa0D375tzkldypTRPFv9bOZ44rkVabTJrsP6CN9L+g859NHvB34W
yTvgYbjzQdwMcTBm4liVuONJ/D9j+2ymyRspVHfLj2jK/CCPmxyQHTIVlJaCTkAAylhnDowWVd35
Lr6KEMrnhTnyCwRo20jYaQARvK4fN9UDjPJXfAcaziLQJeb9mCpyB4ijFmI6TwTwE3+ooMOQw2SA
rhHE0A8pG/NXn3p7t9rs+GTRBvjodYZI+CJSGGieAzxmy7FaA0VYfIP4dRgUjWEBIGYjHAORfPm+
/SB1p0OgqF/nG/biphV9w2M97EmnkR57RIuKeoyDMpP6suU6PSq/RkJvawHSfDSsnykpO3Lelsws
2FrZhPeZiDEbmwUtl5SLPPzwFjBWf8roNiqLg1l1mbI215FVhudSOBXXBUwzrOWgRIRFLeIj1h8U
ZS/0CrWI5RTAa5demDJVo/s1DF8hnpCLZ0bWkVQZYmfpA2F+0bnZoL+M/wQUacV419K/bgQsfIrN
X2IvPEFz6hyygA8bH39l57BqK3ZqVy9rc6gegbilfBsfY4RxFdyLDV9gBjI2HM9ee4Rbftjeb8JE
kqoIp3sHKOWlsifnPzVCHqOyaJsQTKMqsIvn1kekLBSfAh1Jg/hCKX8xJvKeafeaHADcFkX2K8fq
Rt8nklgQ59SPnBUNMRJB2saOTre+FPXRmdnsnCU7am+aM7B6FmjyVl1M8l9016eziwiz67t7HkJn
IpTRYfDb2I/sYRPE8OeQ5whgdDDaB3IOa5r4w/6TmLsz8lYEAoVN27pIbYOYYQsC5G+F1JcmCeN9
Mjc1V9mzQkLIXS5FYqizfmdx8AlSVYrfP6BXh/9DrKxF0KJ05p4JsVMC1wRK9Dqz7GzG4Kp58MC6
i1g1bGGS/Xnrm90rv1v6Q+ks7eWT58F8e8J4Aiaf7KwjiLXCKh/9/TpRHP+OmN5LLkbFSgjpNIC4
+bfg2ypVQmdUek1SsPuevi1dyhxzxelSkohT9jSnTYcDI2A5p+h5ex8wKDaSvDIL0UqQrsgplhP3
v1PRI6IE3Agul5XgmztgEwc9yh6CPe7DKs0702PrGH03tId7FHZky5fTBn1AEzN12x3qEXcIfGeo
/ODjY1Da90vL4DI1AScx761+yyEKZwngsNiZnBN2LFqIWwD+efFq75DxYC6O3ClEi4TIzHu+Amps
uBDd6Pnf/hT2fc17E1ufQ7UQ2RrlPkaBJCSLfBfgfiUMzRjuxd4COj9z1fI/t6G2iu2vZp4VgrsA
HWlsG1BVYpo/NVqHGa603RKAK4d5BdRn/WHks/Sne4qjYja8n8iP2euki+Q1N62de1VltLBDwgVZ
86IsBgmrtCVyH28grmFAmJNYCN0HaaxJXmxNTosb19cXnXygeYQd6jyolGErW4TqVEI8H8e7JwVN
lYItWvKIJP3PrRlK3A6hd/kYBEq14NXAsg7G/vhAoNRS5MLJNwVf62oqvJ0nmqYcf2Fjkye7YMkC
j4KZ8XJ/FqWI7P0WVXpPDRJFo5FifaoygnxclIWUd3Ygr2JZg5+ku8ORhLkpx0SvS5q8IUBGIKl6
fQSxAzwzoVW0jNtwlRTczDpT6mOldEp8YtUoXg6f2h0BP9HraewqGzzZbhmVRPA2ld7bCRqRgH7K
ZOzjZFphRqSgCtE0igxVB50Tvc0CrjUEBQxRvTWAO0mJsv/5oUqdNXDhndKtA+9f8iLNho6nMeDT
zd7lYKBZfKKYPww/cHBN39Z6hKrlQoeFRoVWwgAe7z8dFFlF+061yXuJQfyUGT5NjnP9EUYB7Itf
4n4mLOritzwmA9wV62GUZhCGk6EhXadzbMs2L7uosQvgGE6QVLku9j5ULBQpPQzU9fQyGwVPeubD
M1s7kRvyGAZctqK02FYUhutJXEzY44vu7k2MJuZ+QlrTnwN/GPR9bPPARwyQpGk1Qk70WIomzQFF
adTW6LiPdp5I8SJdJn2Js4pcmtfIMComTG2czycDAFPVzfVIrqGkxchqm5XxQ9GKtBSpDx+O5ugQ
h1PKPulawn3tQrqZ4UUNtyRJoyuOlLK5cC0t41A2uW66wdC+2RFfArEJm5slKgw0WfJ9KO+NcLzY
KYGx3I530eN5f21jAipmM+11WVcs/l3OmDD1VkG1ogLzNCc2YseSKIdA0gj0phZEpQL4MT0vL2l5
pX4+8pjXTBLJ3NbknBVhv5+LJnV4taplj4MPWFShBOEx3Fpz6TRhcgym4lKqXowdGirV1ACwsbmi
PAgwDLqwzEOWK+h39z7ryqoyN3nL1PQ8N7Zm6GwWhB5y8sefBMwaqujrItGyjnW4y0j36EZE3vMS
g8zcVRhM9ZAmBWtON+lBWsu9cgtv+a8GLr0Z6jLM9TMoLoNw973I8iwCfuBfoFjltzFYJRAfmhPC
tVWe3kLQKQ+4elmjrP/GsJ5ncsqOl5/AsTocClfBUHylga1+sEZBdnVcvb/vFAMlmLuuHBHIlsGQ
ivj23/vRTQfCU/X7IPJaixxn9rjzR/2qahE+T4TK3Gr1qaQj5nrLs+x16RfpzI5xtf7nA8VXFzPV
bC4MaUnEE++juBni6MBNNcLaiKzLyQFoNVCUiYK8Bj2siNLTakugeCazkIzqKPd4/BaOyUG/QJOQ
i3gBV2jmeTPTpIOscpzbV2ZYoGAjphPEkXl8mKFGsWWOLd7BAHgee8Uk1jWBCMgpwQ/XFU7JBf04
Bs/kLX81JclLPXqknDo+uj8POP0qAnfRbWu2Nz9I0lM/VgxhTebmT7iN4BzNKxcOz74JUhzGY0/X
VMXnR6hQEZNKW/RNa16xytsRBQXn6wJ5MDVbY/8JdV3SoErf1g2i3gVKc8jijYurTdYVKHoaWzTA
TOzLU86BKz35w60n0jX8rvmIITaiX/T7gPc2Pz+2g/74KWDKe8v+tpHHVicgMJv+irmIbx935P/b
3XnpKO+JkXwylnhOC8io67EZdn4LKPrNUGXoARzthDMoNcamhSSLFFd5xWRz/11xUQujbvOg06yA
iqt4CymjKacOlsNzxdHwpTnTOZ5wizf63vWmVr9RACZW7eEbkc8ygC4sT8iNlMz5gCz0SUd8Rksy
sWrZa9JWcbt0/O2JHRnpl8GyLzRpGCIvxwnbYjnHPszPEsJ4DVsXjY5thnflIVfZbqbrk5yPUUiD
Nh6LbZyGg83weE2+OlKeQcmnUf8e+6CM4g1rGYlQtUhXvQAGEg+9f6sCH4ktB/jladaPeVGPcjLJ
8ARMlet2PYukYHz1NaKRK97CHKcPAwkvAus6+2pDTarLDtIyLfqYFveLCUZ99fdq7QcK/kpu5/Zt
5YhhlXWptNJTdl22zOjljZmKp+dioDMBWfuvk7woJuaekqBYMX2+s3jwzSzTfuCBheGW0NvO/qeT
rV2KIBRs7Lk9CPwIRbY/YuchKyTOv94WKSrkwOkMWHUkDJy/vLXzmAlYrWQCoA7i9wjk5mXcg6rv
+vQt2LARwajE/jTOH0I9HwoQRI0ZesDiE2ZD6Aw+JpMHb31HMX8MWxEk9qGBLCzqzSDj4xhL5VCR
nUrAmmHCa7rxytLPiunyFPZOXHlt60QGqtmKXmq2ZVnVeNv3rN0zFHNusFuXada+iW29424JryOT
KXXsqDl3wiU6PEUDrxxu16Syunl3VN7BKDrySs0gbGyBKpGBNzo3foZntsT2DTpNDJD/HXr47J59
66DJWIA8aBtqhOmVSveHKZQ1Coo9Mmc9krVNiGOvBq9Idz5rSPGjvYI3LxTIw71TKeBYemI/gu7F
UvnwD67g+6u3uD4+GUmWUANsNqoGRPW4rMsrTy/GQLmg7MXETaHi9AEtjc5A6WhTUhpftBEADoMJ
u/dpd+xXJFeXWhV7o20XIfuuNEnU5hmErQ5uOQJh0aFxw0l+tjyWJMItKVv5IYqkV8F1IlPeMrxj
DROfWuIsyoNqnyna8OmPKUaVo40AVI9hNdj11bUmwjcTTkCBdVyr3VPpb2kLfjEMfenUbRYSy1Rn
mcXx8yo2lyMdse7rjDmI1HjhyKwZCIoFpBhfaDkDBAHSOsvnmRYTbgrgFAMbQUgFYhyplCmzDzpQ
Yb4p1okJRmamfoTP3xhq7k/TF3VpIRmVGZTuO0J+t+GXIlfaXA2QY9AR//9vZ5dyoVnOGaKYmIhg
1VgjHgosp3OU12aqMgmhSIkW1Q0BeZHwQTHxnqdeJjvBqmFqRbzLncq36McNkfbtK7BihhR7NC1o
E7s+9b88XX5Hsg6MU3S6J3AGAiZv0D1Q9OnpJ2nYjILfy3ovp9E9TCA+uKS0jpQeq8IU3N+ne+MW
VLTS7PltLRsEDqhRTqzZnj0W4IccXuyJneg5fGOg+lv70WquK+JYzshXLPuv6OX4RxKI2F9qbDIz
4eER7DYF6+mFghU5XUHH2Sew04Ii3SCc3veztwPpDkjfrMOd4p+JUDI447jm86SZD4ug0rjo7rwW
pB+lNeehJowabiY1pX+wCceCLgct/F3LnjhkP0NIfJ4BFACVHx3QnQfqxy8P/i7iDGLj3w4B1yoH
3na0sL8U8HziGrAz414Cncv9AYdoqMhjm0lRfCHDyFQhzTC8pWW+FePS6v31odaGCwj8gsUQQp2o
TQJSgoD3faBCyFuQhfXGifdPCzjtpm/zE6EANuCXbOc3jyr80OOZCmFTj3SKkJKKRbEFKyJtcfHp
qt8gWeilUAAyyK3xM6WePeAGqNO+eFMZPc3Ika70MybqUk2pMX6UYV1fv+fipA1M9jHyvN8/Jm2g
HftMdHvz/QKkFXkw1VDgCrd90weLGaOcGe2xWSMrviIbhV4YC0I/Wt+KdNTF2D1pnSBiIwmwdMtv
0YiXhhp3w+tGCWvV3yZ12XQoOkDhhZy+ZZiUi5my5M0qkmVps1MXO4iJpROOOu50YdlmUTCZwouk
HwnfDkaLGXCpBd13+bsbkLnANtr2Xi3pekv9U+nvcmCGI4WaaOLbgbXuySEaQldaZfXNX+SfxkbT
WDF21lls18d+OT8OyXiTekoo4yS1HUQ9r4JcKVxsQTuxoIExeyeskXfDxOWv3vwvd6lHJ47iIGsU
b9qS1z5TeC0hFB/8Uj8cVb1R612GJQzbeDQy1tCogfGVOtmY0N5QkxWVCyD0VC7N+Fl1mCMoHVhj
1zfDsBjEQwcR7gJf6gDk3SdAb8SN8pAUzpHNPF6l/MpIWIxMc821Pa7I0ey1AQtvzD7gz7X69l81
zSHhzH5DjkGDWTv3J2WD3utS/wbg923HQaGH+qGfiyCcSXrMX/D9JLrxuktffaCyVwwmBjSwg4I2
2iPD9zneZ2VN7cg1cdtT+//Gec2nyAT2BU/MbzTFj3bonABH0hHbJ5cW9tXMT6BcGePz/tPchYyP
3bXKBjnnqlINMx8O7xW2Or8OKoY+0fB3siWHySasOwJGU/sleCMCagG0jvqxwC7gFTdlO8aGouNG
kESlh85+9RzQAnPAHuVpLjP/dsQipg1iYpnRtTx7csBqRlmHsYvaZmn0Df99RJ4id2dLdzG0cYU8
9+O+k/rj9BQA1LWVP+1EzewOrx74XDeNSyfVfCBIWEstCY5BZtST97Yq9F/thCDq4802vnvCnLrh
xMW8zxGazJ/CYB1a+sYjKUMFNABkFS70pjuMyXvmKc82kuldZDUIdVmkhVgaauid+vfjiiQvPWXk
EqoJ6BWBzYSKnqRRz0TBQJWYi52cF8v7MQcdYDrXdNIX5EFwspQxfJW1YOxfO/FW9KincOyqGdr7
ucIe99xRMzw1bl9NZlXOHRLOePhLFK31CXkELrwgXRgN9CGJcAccIaWQbiIeUiglElcdF9izI7YP
aCesevFp/aN6bBdO2kdPIbJ9r+W9alRKHnauy2yAfOWk6ZBNhVMy/M9MClWwaIAfC9nHitBg4q3d
xoDA3hkGYryPFsFmPNPkVU9FNEutE9EeufCo7BsqQmc9twfHHzRZ4kvAebEu3Fs4mIoKeLRyxvAQ
9cB9neb8s4jjjhlqQDkESVQpRDlm/5azMJV6vuDf+ExKzAxLNUrC9n2HqDX6hTwIiyPIKuGGwBTr
GKyzYVTpiPiWBRK7be2Ka/CXC/AlmUzNHpO2fTxDb3y2F+vUvf4Ode0QJaoL6VBLbJ0D22jBrW3f
ukoilx01r6+1FtBxpP7R28+fzq1aWyrDqOYDLf69sj0871bLkGmOuLjqrQClwAxCks83u2lFlvn3
5dbxDOY4oTLYq/qQ+BdY9B1QFBG+/9DjjydOSRxaCSb/HMB6BiiUuaet+zCtyEfF7t5oZSuzGSnr
Z4zGLPBIpGwYgasdZumJFwKL/IjOYJ3hkVqmPdKQYRGgWPoGaTTSpJM6+kHmump/trd2DLYN2Awj
aVLuXXGWWaDfZOVsh7f4MjDL0NLffkExh9EwZzDm2r5D24pcp+9QDDVjDQ7q4f7525NHTC77Yi0E
FtEG62j+Ht1FNJqPe4ELEAbm65Z6b83RIDDd7wX3LnwDp9Zm0rlaS2HCW+Fd3Mb2+pdWxXKIIRkw
THjUtXxIx+sLU2Sfmcl5QOhKA9pHBgEcAUlMd922/atzY7gsKCtvHzHQbiBIeUeEdOnA9rB6bbHF
OFkBe0Gq1/ZT8n9+ERFfsXFa8QXh9SpxJ3MiWOQ/upFWTrs+VFmsXu5A/1TaVkZ4wUiBeAX66enT
qEZgBkWwZjDyEkQqzdP1u99nfVSIUm/Ml1pNx2a7lWnqhd50TKArAzjnzJG3PrCqtP9s/uW6CZIS
1J1MSCOOUSG+fWH2v9xYNtUbdl0IqMA0h8h1EP+73n8W/aiEvtYWGk+GFjOO72ADzdJgSFjvRt9l
892qPkHid16b2lrHe3R/75o6xqBghr+mrN7Dkx1Gn1BYJjGwHxASXhkR4O3JbCI3QfmVQtZsuBa3
0vCAd8ntfAAWPSoeOhZnsVDluSXawO4nFZqzQjRWDDRDELhRZzXPGEMyCEddxlXHtZ4Yd7LuTCVJ
rYGRDpgRrXoxQgsEFHbDOI4hNrl+5DsH/+iEmTfNtDfUN3PzaOUvLnMaZD+QuGiXHMGgRInyGm/a
ho7v+lYdrGCGKwUYmaWgghr0m3GhPNF36ebsNFDdTO/tBc7gCE7egaWo3DZkL0mbpuaUXbm0MQ9c
IsvdZ/S7kVyr1+ZledRLjhADBarcoq/WpYn45aUav3az6Z0AeAa1gq89cGcGC4bwNQF0BJedqrAJ
o8kn2/MBDk8OIFwh/W9ksSITKaFEeJCxGZ93FPcRvk/1Sj8Gh/hFb28wW/uYnYU36CW0l3Xni9z2
hyo/XLPEaHR3dLsyTh9fxOOa2QThzG0hPKK6fjP+3vgJhSdApUxvI3Q1HnM7FpldXMvUbdhlXZ3M
fH8vmGspxjRU1zBpahw5xRdtlddkxfqudZbkrVSw8418OqH15B+LgAhTQ8N2/JBWV/Lbv+M11/m6
mxwL6CRF3PgG/22juaAvjpqPlLyPO5huZS7QLws0qAHNruzWak15lmlmftwU00S+TZvLnJLVDy8a
1UDfVqAKLnTCsd3XMndYKUisI3NzT/mZGNi10/JIDq/O1bpJHmI4iRpKWn0PZQViIyBD5SQV1CMt
ruweBf64rKKsv1XKHOphFHKjVqAvYHcTgOZ4sWARC51QqiPHrQ0axi2pUUSOJaLWYsKHOh6ayT6+
vai7KP9hqSOyzwERaYeAgYVREDi6wzy6kH27sGFIBW6x39+awfFkWwJKnuCq/m6oBCXgLT1FPJW/
5MLHG4Zh17aR5Y0j0+ThyQNA6ySveokI2GjCa6Ej8WF6WtWAFUHGlGGELNoNLgzQlulhkZrQ6xDx
rUa2hIpLK6dDiAzEkn5s5quYEA3htKJccupy8LiuXqir55tzlqLI/yYV8bItWK0XcQlH4hVJbngT
bzwpR85UCWsEme5e3N658MItvAs25hJsL1nKTqm2n+WzfMpMKSqMYxRdy4U0SRsndhnSKsAJGD0d
hGOGJkZqNsGzFehjxL4gLahL9+o1LMbP5KoVXs8o6dPbUFhQZyx3wnvG+eRtc6slqTXkEsLVdU+t
WBROvox1Q7Kcv3H+7eNKv9zn+cWmw+qpx3v6UCLQl4HeLbcS/RO1QVcHtgzV1vdws+0aQ4D+iHRL
cpyqtQDsjE6ERk9pmWql6azqsv1QeJ0rTGtWgBPfwEX8LCY1iJ1WGUb1a127FY5wIenLrekDDN7Z
duZZrDx9BZNbj38RMB7nAgHGQdtpJ/iF1A0XD9Dp2OorFKxumJZr3TrJkcfeQjnH4/nCoNJekJ2n
aDEI9aPOy4IAko56PghiTTCrdHWA3GOlDwbWhtGG/nDb/X2x8xFDJBLtiFWX0o59BqhiMJa+f5Eu
un7h5YthH5a3ClccW60QKoQ+iCIfmXNn0E3c+fTbaRDAgsEaqvaW1LHSV/3Zi+ehBZ0jkb1SxxdN
NVEqs3zgBFCtx5HeCuh7QoQQownvgSYdDAPD1j4Q57tQO0m7YBafoC7HnmQPUv1A5zXBBwQGNWL2
/PBLl8UROCB/xynqmEQtQLAo45C9SLudv1Ft7+dfC/NSoRfXNX18Iqub9eu5hW5z4H1NnnteEl5G
R6NunmudNrLrnYsA4HRNmUCMlPOP0ECJBEa9XJMOIB8cXx2NGOUvUHsHadxBl6zUHzibWbF1hRPR
SuHlopza0fGkG3FkBihZaselNO02f1SzY+DX1cWINA8UELw2nj6I7lh4MzTedKarqhW37br+gHXk
uE6GcIzJlHLHMZLGryZpp6tgcrZjwIoBhR8AFuQ93V6+aSHSg/Phm3qS0uwg2LcmAjTAeQxC9spL
PMNnisiR5A1bmflc9xIvfXwBuIc8aCWjlXXd1I9jCpaQcS+mWYIbg+oVtSG+mPt85w6dx5mQTrdT
9b/cSGRzKbWuJ+XnBFOgOpxOYNoIxGwiLPJ/S+UVFMU4F9cruHaqQPNX8Fmlq068IlZRuJdLTJR3
V46oRRoOlotEJp0u19IOfyIwiCeN2k5xuOkNAYPNkfl4w6G8Q+T1SMfJKOFnYMcma5h/DDH85RlY
/Ih3/37LHQf9yhyPTW5YTYyYWNYIqu8hqEvaIQV3Xf0To7CHsj6e75DJwQvREGjHGIIphBnvHlnE
4trwIXKxr7f5BOB4+/dWSur+yqpe5UP9Eom2x09pHg/KXEg2qPvn96FpRJudarGFOqcQDQm9IHYJ
OCwi/O6GijwZJkOKN09GD0O45maONu8ydxUY+NLzHXKGgvYCA6isXIyk02WuQhJtdBAh/hcckTmI
s8xSs1VH2bKbeXko8tNwcSonkn5Vi5cBwUq9eOZ9ckNvn2ovPWQs05kVcUidBDtChBwF0TtY4aaO
JuCM/Cyk7LRKyq7EgTU1LscQv+CZ+1vehEXAvESlIxC4mWIZtejs1HqpXxoP23Vvn6Af98kj1+ne
kiizPZtr83gjWNh+eDSm1ivPDrlcexzABts0OnqTJq3FJqsDiqLheevQGNxep6oIKEUdTVUbR40Q
QRsGx8PeZ2abLM9ZG+oWcec3Hk+KF6UygvOeKLDS1vnmWPsu0rHIDHKKZ/G0PxXdbVr+8WLKgHlY
lsaZrGOCqVQkAAJMHkxz9eyNrYPvfsZEt91xUnNiAshgKZVxbY5kG/lytLQ/ywH1h/GwKElAiuQQ
EmB3mQ1acZYfY1WTW89EB9VmVAJSh40F3WzA7JWuUrN9Bq7Ad8+T93Ca6PV9Uf0fdLJhmdSbMRRu
SmSAu5tW+C4hBTn4Ap21PESpZcI4V/BBmnR92t9MkIH17aMm1+ImUz/pyNFR4p52wL0xjRjKe48K
BtT3qertFCGziU5zU/sTtl7FDKz46DfTn0rqc1cOMX/+dIQnrRI3T21XloUj6V/dZZNxv2BBROgY
4Do31pUos5ACBa0wWSR5UXuyBVYxX0twxYy//zXMp8h1IN7OOQT+KSdadnaxiXRS7w7tSlRrjaF2
7FiTlsI0nKcg3vg2YLXlde5FCdmcIPF13SSWve/oW3BIABqFOGUx54cxx1N4o57KN11RInL61UtC
ZhXVXdM938QKJNGA3IHvmPHZddP8U4cNePyekqJmBIpmgH6ZwZOSSFfjZ2fyfgJqX73d/uHZ9OsQ
YNMORAFDl2EQ+q2kHhTJdlNlIN4yeDAvJUqsqvzmUETyeDcoFVlCjNNXB3JeKqyyR1APVeTSNFJD
KQcywh9ePvlWmMEjADAa4tWKo8eikHUEaAKGtfnwBD3yV86V7qIKpWDmbhRenF+f6qUkQKPZboTZ
lO3wBqertVMw/A8AEDE1O1j94DGXcHvdiRNAsBHCP+PK2CPT+fiHD57/vTuNpEh66zIBwE0OJvGX
Z8m17vYxiZj0L/O2nIXxCA1Crkpb0rzC9JS1N5bh9nlpV6dS8MjNkToSv5gqixJTjWI1PJxVskTl
ASd5DPSLBNW10L6jpgZ2fFDO95C973E1SZ3zsHfyADIS0UeF2NnAlct/uUSftUmcw4X/9GWTgCLV
FrRm/wBtAg0V9MxWTVflte4OVJXRuTiAAGFxPqkBEHS+ba8pvK6eOES/8MzvNHlVXr1AJx0+rQIo
WmCjv/r0oN8bU9qK2m02kqcpCYvX2HUSew57Vr+ySfmpTtytpomI8gtqC2GNgkN3sYw152CS7xVm
Q3K3omIW7sguXrTE+TIvSyja2nIvGhGF+Mva5VtO6tfmgA1mHY0l0vdOtgRjAcfvEaawDx/lagEy
wWpDlKytf/6Bg5Qcr+CIvGM7IcKBVYh4h6lyp6r38WQPRndDNO2ytP98P9Ew77tu0CebfZHRBPbh
lLDtOOqFEafljSvGjFmuMijN14hPONkS+i7Bd9wetn/vVPUcFwB3zMOEFqwKsnLN9XKKyNWnJByf
AyFAJFu8a7YW0YjUc2XazDGLZWfj10jyVeIfJWYLm8FGTgnwAogwFOAWZXDMVG1/jT03/+zYrpbE
XrcVZY+gjURFfpoNEWSaIwJsrFKA/GAKxaik1/QIkAwXNOT1JdIa9zyGmt3/iQhQuFWZ0u5ROdHs
fpeewhvSf3vf+W815j1THKDWBVBUgbPJUZ6CFhCGUX5YeL+ekK0Bb9wrBTDo5gWUelzy3sYbtfLH
10RkyjWMH5CaJ2gJZGKy/b/ICWq/n3tl2t/E62kyZUtjUPMkK70mjpgk1OsVwwsG5bFOIDaNN9in
BM0hQBwROGkk05mwvX++ubXztz6CfZNbQlZvq31V4ZN1ha661yus8wixDWN8t2N9iDz5DnWwVbH5
jlEivcuHkiaFFwiOXsbdaI9HQxijt4bJ9q5pw+R5K1xDWbko1pepfL49dUOtsLNvK327x6wq5Pza
4zU5k7ukLlDd8bd2NuDlIpUsaRK5buEjIkVbWJincSYLoD45Ibvtzw/C3VgWK8mjg4bwARnTW43h
13y6ZEvXUf4SKlcS1xnj47gb3qpODHbONZht0JGuMje1kJeOnbXEfjVWhc7vFpWAXkJtu/kkNIdH
uM+99mhs9UMZnokUw0J6C/2jcbf2UxFIU4TeomS4VDgvmGBnvtruhX28vP184dRKUlI/vJSo0ywh
H+AaoLkt0dmKi2b8iWguko8gYFivR2wH4i4WXqWQ6TVZj8vxgTKzcEeH3uX5wBy/2TGAiIRgdDQq
SvKIx8vV/L3UN/PhOv651TUgrFLHp7ir0Yqfn3Hqb5Jg13vL9jaVaPcwgoIaJpRvOMDLsCYnI1Jm
JVV1xo/cBmTGI/tNluova5uoX38Ny4a2VC78lDAFo0ToMUPUOZj6+EpM8Fy+vMJBGwKO8WFKqln6
7MJciWkFqg3p4nkaZhceUEDYoqZB5KurLpfZCZeNPDvw097UXUEvE2josGDS432O2moRp55OeHEP
IAg2kSjulVz+ZWfJlG25nofAV5FUr/VZoGIBAiCQ+ZNxqcNAx7yKPNcf0BMF2A7MqGq+jO41VslP
ZoZ5JeZxmUrndLHZ/g1291fDB9BqIsDgbhISajRBJZsN/WIxDmZRaL/rytCYXh1OfimfGEJYFWpz
5kmgv8aid06s42IYby/Ny3c6TOP6dX48qWGXfDcrFOLZUs1G/aJ1i23UaBLrD/0kwLBWTwJTTv+U
qDbFXPaM++fA6B81OXJyYtvL6vkaJHjY/RDowUZJDN1KAV4Gfa3WfKVewP3PleDOZ+jsxjtOwTjR
Bjk8oAiSxZagXppUQG1UIdodlJn34JxZrWILzgVbIO7hsDxFA+n9L8Ir97fA9741wyH/h9HhEomz
Hb9HJjp4ZIJCQ/4onGX/URhez4YCAtgSj+GHlNEWI0Q+lq/thJ7oxnHKQcatd2pe0dw9qzA6giNC
cf+P3ylSwbkniTgTjLpHYgOfzayd8EUFpQgipZkFy1PmmSFVSfBBUj5oLs4Rv+I77idnEHdO5Qjo
no7m0cSiOwtN8eMx7V5lipClLMNIwWnJF/kuRmeeBiib9Da62jWr8jz0+Elo5UaHv7B+qrKtJQ49
dJAzdoVZ6W03TW1FJ6ydcCu9fupMtE80jwps2KAwGT8m0/qfQklnxYK1NebWVGuW4hYEqMWF408n
56qw3piHguAJGxSilpyvyVr4nzw06W8Ue+XBTKuHieGTfm19RP2geXxAhzxVkm8YtjVRhRzbqwtn
eUpQC3FVSscUoaWfx44JejA6t0UUUQKYO5yyA4ufFV0yW+9JA5FsjioxTn+P9zUPaSy6EfJIn39H
U9WqS9AdLmHbJRn7fDwmyFw7LDbwxr/H4C8teSTilthZwuxZKuTBP8G5Sbklh9kbqQU6RaBYS2W0
YA+WIBdCYHG3bgr1rX5H/dcbjQnpBBbuwdI6+05FlfpfNKsohjNEdoyk3TCzwulPZvcR7DERTqT0
dYfmL1LXc8qOW1Fu5GvZBIqKOQ3APj5WM0/0Cx2ogzsg6AMU4X14kWMkx9x3AWRU8oHkjzYi8Z1u
dWo0S8Chr0TRunFPRG6SlW2PEPNVBCtQuN1PeTCeof+diPncmq8m5qwUw1UXxGZDffSiJBRyHQYq
+jB5+kar2BiWODf1iVzq+L8EGQy7/zlQC0068pt1EAupHn2QJRFqlvA7i0lltLMJD0EcPMP7ALhi
Sp6KOELpaHygqbh9bwJsoiAQqOogZxK69i+aMNs2s/KHSx4tUuyEGAAxey5iIcnEok0KTd2j14D/
dGmfFzY2pokHX8i0/C6W1Pf1V4RodQJ9VfKbYipggrB396s+h0yg3yTBJElHLRFy/YuMvIpyQeYi
D23F/X8NU7sr6I2yWT/fGZUq09NPY3/BeereHmIQLhKpJRNfhw6NKBaYrqZvxi3NWHA5ifJd+AlU
+hfEDRZZdY6MIeJ5s762w4bcYZE3EkwUzOxrzAJtiMrjqkHvuxhy4m/hUJjSprr2aI6EJVMTLjlO
jXE43I26hhAx5/W9wiDFk5nMNp8UpDClSsC2hwwccbuL1JHo6S8C7+inCf7ClAgQ/JxUdn6t/VX4
Ykp2jnBO4j/0OiakR4SPrQ9P/wKcqOQqAgF+p00bS1Iq9+6x294NQCSlMuZeVtFF2oKeZQ9HRcjt
liDh+b9Z73ZZDu4WDNj36aFfw8o6bvTVeXn5sCSdqVQWnJRrllCtbRQSY06NvgWmdyn+npt4OUpG
zYm/LD+EVDjhbfDHQHj3w8/BQHwN8tJzdSx0AMAKGVacSEQ+uX4BTNNKhZ2/VoXAZN/496mTpDyJ
XwolD8zJ1KRIKFa9PQ0lF77/GeW1MaLHbHJjhxTnpaW6MHwB+oOctGiYZkPo4VVDW6OLfEDwCj23
QBV5P4JqPqhecrdlsiFl7QAYm6IquAoTpNnzYAvekCAfWgzWE86bXzSCOfybr/zRd0+WwkbMzaPq
AbvyqCoU4GCUNjFxU3xxE8wgmpRhUmdmioEEwfHS/9IUBwjc4sZEppJJ2s2iRAdgumUcjeB8/i4G
hmO5AlO2hBGXo1RIl5oBI/JJWHSCf2HTFZb14YAnhABHnpbuLt7vDNarRGiUdF0yESFpUFusutX+
GZvzeIwxgBu7O9kp0mPhWpqQWWqfSWWvyz/bNi9+NX+LGYxPqaTQMnGMWOA4diy9FxcwdvIeyQ3P
IkcdjW5dzxHcPTePKtneccByDvd/Q7AOet2jGv7aq5mzkAVR9TuPtm7TwE//PPXSLTvX5+9gp/6K
aoFN9/Ta5vJnP/FqfGPfZP25vq3l1ethVXxXWUJGSd52NcC7YyMbG4zWtyPQieN4+o2zkjzZfPNU
uMZyEAIyfwi6wFK44yK4Uzijy4E/JB2IFNG0friz91R1FegPcO1SgEs+rM+5NZHUzLM9GdD2/3+x
PEnh9qkvS7NL0m/YpCEwLXX+iKeR1Nz1WobYo3CIxjqYPyMWxn1mab9fwDKYN+hKH2kknEcgthv1
oZ80dR7JOITaPwsjO1UoTItJYhiIQSXjkLYu3adcr693StOCfdo+9ldEiT24Omvw68lb+IPxltFO
i9hKFFkInbYod14y4B+jQtlhLRLyBwnjTdkuTBo3wOOncvZeTcqqZJ2XKiTv5v4NNz1n60W1mGAw
crOWAQ29w073rY9JupU98rLa5SIdGdbwHjbQmTohZfmF3uKVsndIJeYjbyIVXEDBtCmkOxEl8vI+
KmwCEF763zNKIC43b0WDbrMI3Qv6ZAL/LautuY+0Lqr/P6mMJMKTDpPqhcpyUabfzhKRH+FoeD5I
08IgKA624E0B/dOW71rB6FUD9Ale3JPcQ5dWNJqkWhNNoDpsx1berMz4ENG6UiuFd+xwmrV+3mKW
UFotDob9SM1N1rldOSxZRZnD+FSlBrKtkHzs5ckSHJHNsVhCLIQoi4VZHduAgw+bTgXUhZtc7edn
5YVxK1zCIHEMwBHqfsIhtsfD7PsMlGfm238MdMYlnf9bq2e1T+LlxyAyoEC+coAMna/BOa3AmUBA
uEz97YbOuxr0SrK6Hw23eXE7nJe1Q2zF6YD3ys8x6hpNp67Fgocacg1bgeHazn/tzvQAfYNRPOxh
QKQGAHo2TyvEU10yorsum+r5IclKGODzFsYPUX8n6e17b04/m59ywbFgKqJJVtFHMUZbuZy4kecI
o0zWQMOQUe5H+LhAya3cPEZu7HszkPruVmmZ57Aende+b4EwFQWPLL5GKR5zYBdgttzi9HLuyGZs
kdsHr8D1rwaEMwBE8If0/FxtR+EqbLGG5EhnoVjzhpYWKbtIE9evscXJuUHDdNBzKMjcEcSkycEN
fL1KMIF2BYulfP1+pLjizU43+LpdqO3KQk7FplAk0ymTcBHUCu4v9+PGaBQXApyZuEA6A6R67Tks
SGxfuZ0vDQDlhjMnsaS2XX0VEP3/s9Uak5R56kNPK1y+xGJe6VWZU/srD3O8hz+rmQCxoff4eP9K
EGkSP9aUL1huTQT8SThYjleEhdV6ndSJHM+lqNBekkd2e+S8r/t/Xx+g9BM2+JB1Hu2IzTfynfWq
jnC5a10g3HVC3ScUDYevmDL+acS6ettdCsxJmtm39IBNvqiT3qKLfmgt42XwYkJmVw0OSD8ECYhj
ofx6pUT7rnKLz0u4Aav5rLjRaMeyw98IKoOHCK6pBGtf1kaioLjbUGOYgA2/1fLeL4kLWo4C3cOK
ojxgndEk/KvFx6m10aeAuZDSw/1jsY3UIXedHi70LDD1fLXQLxDaF0zKS2c5XCy1+LgGGx9rg0wW
G7AJBEvfVBtRXZwntNC7hnBAmUKw+3HX/mTgRV3qdPWouoTqqqdIBJ+jM8LsFLUAPFSrQh8PEiEc
r/XMY7LTbkqWboo6Dr5KSifUvxEqGOU+KQj5j93fLyU+dQeseqYAnnjVL6XUhzWI0uGGFP6C1iwk
kHrDRWKUeHDKPEB2U/EFti1GOF0pBJHghgCrxAErGDQ2CiBfWwJPFMaGz7Tbi5XeGtuE6bz+0WWo
q07P+yDuz12R8zjnAekD6CJN+QohxwrKk4018gibR1BHcvYM5aSvlasswVjQFybrVWtgEBp8YlMN
1KqYruQIvp3tijG3zo3fHSH+EE5+5brRM8rmJ8Ug3oorMhzJMmFkGBJTaZEpd/ZXxc8IJHGWtMC/
F/RBy8+WjQFp7BAP+07wVeQXJVDicttkkxWHis03yg3AysVaz4ILHV+r4x0manBgGcO35XR9gBR3
53DQzmUOZpjeK94z4Uvv7MxqmoFBShKm7J0uKA+INQVG9Vj558S+TqxL+Y45VUeIWQk2LKS1l9ml
y6BnZgSzvC7wnYp7wYxhxnbtGuT6qRNKd5wetmyDYjWd9C/gEp7LlmcB90/kK2r8M26HD7G0nCVu
FRT1iWEpehOGNVPW13Xqh41KFR69grxHRvHTcibX5at4i2lW1iPYYKs0xmibZr2glaJWA/teaKhe
cid5rspn6VO79GLhjYqmaUElEbAGIvqBFpELUVbv9PN5wODd+uXPGVUuVTMPHUNxQBYK1xxOl9M8
3cyJSglerXlh1UKPemSCZYppjiCZ714FdGIM30wp5y9wmgzaEd7FHqgNvB7gJ2jvn2HGiHDqDirJ
S6X5O42W1m8NSm6YHiDZSWd/jUQjWio7EbczWfnrLGy+BMdNGkb30xDEN9yY1sA1rNIwqkxiQ8Ut
lQy83q1zdQF3tWV8k6oB/EycggGoPP1XcmS2XPVd1YpDF0BJnwDECTX0yLM8ia5WDCXF9jswkL/V
RY2buKE7DtLzOtHvDs42A0VMxoPGLv8F0iRKXbsmvFel877FxNz1/wygfU9BnZXgvCtZA53+wJv9
n5BPOWmKxWDHEqqGDQWpiwtpKHCSt+gJiWCBgQXAPN0Kt8r5Wipg5FuUwm6eg4NaTQlqj1d7Z3Ga
mNyWMH+MKcbCm/SoqEjOnygCiP3RxGT+OLGlt02bhhK3VHH8L69wLEdwWQxzA0t5KBt3rwY6Du0d
FTUfv7aoC3TgQjr+ZL6IE1+ausM9tkeBRIsEf5g9/XK1o3X7EIdTu3LXWH9+/CtUyyl+TCAL4Klf
1R1hS8yOw1PIqX4cJ9VYC2HgrSOxpXGj2ICP6RkFvGXoD0TB4Ee/2rtlOFj2IwLdhzfLUJVoZXkk
MDUIWaFWGH/+zMS7FGp+QJc94q5jJ6B0F395mcKf7J47ibOP1GUq9otfk/9E03MHLWQuRBkFmn3F
IC+orVHukEYRgrurvOKe6eCkFlhCo7V9ozQ3HWGWbmsdlbXPJ5yqu5bc+Th05Mf7m/fa0RZyvtNQ
SlXdEbaYBV5ZjTpjs0NJSGQTdKFdtnMu+FWrFGQ1+VmJihEnEJw7NoegPFFCGWwlnn9YQlFVjjII
ulDDBlljbw0umRmOOGpoEG4zxk4AV+T0NnhX3sZReGkll6XQBXKCmKATFlHjR6yqTRr8Au9aTTIx
jID/vNv+4M7AQe+xq9xV9FqTEYHM0Y57bGCW6nS+rjGLKAP2Nz80htCTWz+AS4Dzt6Uauvmfd2HB
RDBIabzwuCFp/M4Hw3y1XKe/N7bwBseZwWdXv30+kEcptKwGFVI5k4H+6SoYsdQw3gKLVnUJ035s
UuBPWJYyS9xve3COjbUTwZer3TR7rIQbrXtg30/g04LjUrLSS8i1c4nrEEK5pzeUX6XVWZRiGTWc
nQe0FE/y3mAn4isxyURHWtaVoOFAqu6ZO+npKixv52gryajfh6imGloTWn7M7PBw2MvirUZ0qR+d
Vh/SepJajHFpWsRd7kSaL36w93QUYNBcqbEN0Bhg+qClKMWJ8sYOR34z29eaKpAafJaziMrFcdMZ
vsG4iEf1RX4XVNlJEX68fYRMXEIsYXMg8cnFd/kqL02H9e6TlFHhz7GtvdNFqE9BGKLdrn0OFD8L
ZYoxhFRxxkNwLQf3CX1mxNHhz3q/XPaMHsQstO1H6YQg1H+P50ia59NiZbR6eTDf2Z2QAXIzu3nk
jVLBqccG7HymPn2XqidimtH/dLO0jhR5574Dkow/tna7GVCtAQNeLCl04dToEE4Ea+5cdgQVI7Mh
0wHkfZo0kwCtLMVRUOkObaKA24IBK3f9WNUm5CPKiswR4vE8XKxQh89sjpYbaZyaSMxKgPoFRPKL
iu/trOfHAT0JmxiwPfbCLIo4Br8lQcL+p8nNYRE+NAAw5vpJGk91lLIu4qqd13dC43wPLlZ3UjeU
GhYK525hsUT60o+Kw+eJtCZXSEPJZapevAvehMTGTaC2KpZw1BhwetsOIItelFBbJQFmEAn0+Sxl
Q8jboFErolU/FS6gsZOJSVrQpdzVUCsMRVws5BdTOoYU6SyoYnA2+5JTTnQ6RUCzYG2XT35tv39e
R9i6WO5C5tJty68s70Tz8rc5mdtQeJnqi2DGa2eDQSbNQo110kXRIUe2+1I/Zd86nMbvxHwdz0Pf
buoHZOfEa+Cqfy2ngL/f/hjrrBWECFC9ZjOoI8y1H6ODZdCpFNB4UkVvcgvIBmRGQ8PpVW8zgTvY
cf4h57fAsrgbv8+lN24Sqnf4IbRbHhASje6jP2BrKvF6cTvEDJTh0dzo901bSuYIiOBxNlavoWQA
maypr8JYdnZN3wWSfypNEHKdKra+JJ75QZ/3rIOfLXjgq+/hFsKK3d9aDmSphQl1ats/HmFzUpwe
II7xkEYhMpCnvCKbl5NnOLHkfdFd5ndjNrQuJsgg/bBoxgRWOgjAuL4WIyWkUe0JpfUbYs/ZY0m5
RoVxMEyDop52zO0i4mkxQ5k1Rs0CA4uzc/SiZKAxseql5ymSgETnLluHt4iQccTMTShHmiiCeZcO
QJcPahkWaj/eQkRnMN9AgcRgPM9/oBHF6lJVc2uncVYTKV8UngUdMJ1wtpJOOL68IL9gFw2O95X6
iXUuKT2EL4FaQv6O1uTa3NqFPzBnv0V1OOgNWV6jfpc0+DOU7bau2VpGHol78abLdwsYRkiglhma
y/PhBUyFRUk3qgkaJvJ8/fesSnjubaqYjjDSdVzCpgZuyWAfSwobyuDH31MgHyrwnb9ZkIbsTOwp
qNvpOkkIoeDxqrrZYLK3jYvAu9XVu5ualqBgzNigDaxRBwMLR4V0OOPnHt85vJYruz5tTix3CErq
h672X+UvSnWA9IzeYXVCNivnZvz7qPsgjv171wP0CWmMKENl+lM/LlkvmjCDgcvNqMrgKTMlMcGA
qUAwE6PDt/ru8e3lsG6M8eWGNVqKHBzCFPgXmmMRRJKEUSNudDWG0VcBx7VqvFB/Hx+sgXf0cMG2
cRYFP+uOruTwMja1uqj+Z/2iKmnhgjfjiSUPv4IS/6OFX6EYmq30Ts09Cd7NbEYANPBdbcy+58c7
QFNTmsWoLr18U2c6x0+HTYEC6LvVZSkcR3yNY6mj3J3t616vjlpGWEetmFid4WJ68InEBYkO28Ob
d0qzQswQvgJZ5JBt4MFJeSm0nbSMb5yCxTUbDxunwdG0zS9n/HPQzuQn1qu5hlVi6BUQTlcBeHhB
QtxwPjhNWxS/q9Clix5ffb1iA6FcpbYHfcJ6qu45Hy2C5v+/lbAoPxLUQTKWCIcrM0UThFalEEOT
VAQf1i23mmcwt3BR6ZKJUGCveYHRHxOlhd9G2PJxUSjJ1aZuG+g5vKq0KJgzNjMeIACLv7lY0FMj
p2ZzB4N1CS264KncMd174FqWkvP4Lw2G0leWaPyygdSxAOSWuI95v6rfxeMqIwNFnJE2oafTJe9b
6nSzotVjpudWAqx3oUj7z5ljQL5unh0+6I5QH0ay1ehkx2IE1tbQUuKWfnjDagje59YEkLA8FitB
6Fsh0Jccog+LB1VcBm3SdabdFzNHQex1+Y4wDrMtkhW2XKTjYrcX43iZRENbeB4oz0tdRPFzYKso
Nde702taL1O116/Coj4yWr5zDOI+DKNiXKpm/jaJTdiBKrBVSlS6yJjKLYZprG8fZxV/7rB0ATsX
GudD03EwLnwjYLO806tBGaIXGGaCQ+9Aw6y1KzImMxjUaOjODlwpzPks1Y5xScPnTmfiQm7g+w9E
WTbrFf0GFUs8yMNQPxL3vPNoqUAglqZbFiPWmalzcTvC76+3Ks9gckZ8nXWwzMHxXCmPqgzHt3NZ
szazscm3KZEkGgnrrBECj1bT3s7GBbDi+b0eTohgvKDe1oudPPLuC4j5sPvehaIUl3HtXrFVI7Zo
DIHxG657Aopn5p8khu2QF5aa1j/b2cOujBd5GJilNdAYTn/RZXjHYRTOdEVAh3Uw9G5EUFH63b2s
MNhSB80GY5CSWqu4LWJqvzeZ+4B/vl8FJgmZ+5EpqL3w4L2dGOkdKcjIMteOndO6xIhbLqFWU5dd
mZ/2qjivUmQAldbzLYwcXe7iRSweU75P79BChdSsuISc3RXldIFn2JAPc7Bckd5Z87V6e4ymhkBe
9z/L0+R0lY3va9DCK43W1UJI+FWOD9TUN+SyZ1DjKjprDJk+N2DqPiPBQUuJLPrGLQ4xqljWDtBq
w//dJRgfEaLsl7BtSUmiFYmoLDkk4VybuwqB1oAeJp8BZ2uYsadns8999ZMVpoCdcjvygi0Brckx
fAF49GoBEuBMxEvx8pTW7wPcgeM1GGVSQ/uYSU5FoMjtVXToh/DzsArAletDsdlNcl47iOnbSEHh
qaJva+rT2MfB6hz7ZjAQ967M3pEN3FqfhlbAXIsycZPQM5ovO74LFbHa/Q2QN/LK6ic6CY9+Y3oA
cdZZfjnow3iKeBrfe8KdBwZtF5Neebwgthl5thkpxmJQpFtEDuZtQcZpVbqb7C08rr9VWEgfRlNU
dvGsPFNbg22iZONzG4s1X8NLKld/mdZQ1eRLB0VWSVcTBsMb8xWL8KlOnGdi19N2qusSiVNCgnxm
10QjM8l+ErvVmt5u8C/ChMzQIANU7GCJN/GDb5i3aiDPLn7piSVWEoDcdl5+jI1XNotUej2m7yKH
JC1P1Bj9PqaosTD0jpBK+uo1HmLnoKYaTI0tBlP1WjthYLc2iEuAzztITr6dPsgq3Rs9/hC8/0Tn
gD+oYUEPZW/U1+6FOmphXDt6aLvibOsBMuUszrUZohv3iHyxo2fR05kuSWE+6vUQrIdWzJPYRG3Z
/LOSSjLHXt7MyJDBMu2Gm3tsfzpdTD5Lm/82oTm7YbbFNfvaHwgGABlb34BBjjGCm4FsGDTF0P0M
L6Lxiqg5zbCH25h3sTwJImI2QjCJwIz7ztj0OeQ/NJztEnmgi2ytZW8Yg/6fY7a1eIRzIb4u2fXu
xHzi10tBuczje+bWAgjF+XZzx/X1uCXfaTiRCZArHyJZXr6sb3KjbtVlUXu/orzT5/EozG13YisS
Ug+QSRdJkahbKKYaA6IUJYXe/D1BoMitrnjfW2B/BKyVJhiK+oMBCqoqLXmJW5AtZNYUYzpLoqJ3
R57Ux6aXROzPgm5/qxf3UjLrUBRUk7zKgWbTClJyLSfs+aG/a/W9kiZqEZznrDvnwnHixJBeilZe
UWBhrab5dbVdMZrTFrC5K48k02MXFtjYw5mymSOivv1WYyf3Qx/nNoEUYARbvhZQPb9TWx2gcyM0
SzZdAzo7NRLLi9r+ziHzol8mriIPIS71fUkyKZ+NU9uNINGJkVrlubGwoWpc6YWOOOnFNzUxc6nF
yriC4rBjcBKoQtcLlxENByRdg90T/Zi78JSGU4dsTwzdT8iKf1fdXOxGvqnWNrnFQrcXw/EWzQP/
YgY6sxP1fDPeJG/50Irph/L+ckrw6PsE23iZFlQeUBaoin5xbkCI3Wxke8DZq6IR3wFEcnnvgQw9
GmooWQWrfOST9RARvrTyKbx/yZCykUKBIKH4vZGlqB2BdCC8GtB9D5yEbIkui5DcWNJ3DpuaQL+d
UyMrbKT/fh6zn0a3qiCQhmT7ZxlKsmRrsXPdNKiJJ6t+tzG6ZnOHMS+6omTsFWr0rYCSQ7s7L7+L
lyp8mralbpHrJSfHilOWlHls9qL0hA8SZZ/T4gw0dfudD084nRArmmbZmnG+4+sLCd8iACOYYnKx
LnNMN01K84ZwEsQ4Qy6Sym68XGSe5fXFp1NmRXRo5kqbjBVp2tMomHXV8rSBWyMJBNISokriX4Uj
ixdSfTedKr08YiW23WnbmaIqXwqQOEb/gFCwpyoE/+Z4XtdP75nM9YbLrHS2hfGH3Y6LhpxEwF/q
g9GM7w38uydVqYr5i3kre+YJEvZmwoDGBgKuAA50FGYSk1bUxpHLHkNBaablbaAcjQOacz1+GUgJ
2ioxdx/Q76ufBidqUfD6VSHriIs3p6/QvMcNSr95FpyWJfRDUoE1Q/hUl2OR7visebAawbvoopnp
raE3OnLcpcqTM2So+Hl/FqzoalnFWN6u7PUdwdYrtpmsQhh34YZ0o7Q7LoF3vJyEaSMIdx5T1RM/
UktyOqmPfQX5EPqziXi/KgmVTpajZ8/Vg5ZTpvYpB2YK2raBDLq32Ea6JbpjhwuDpXJ04MlhL1OX
idrZiJdm+88i1Xa6yWfomVeFV5nJ42Krp7OVXHIXVcP5y0jrWDnf4w0Ahk1KVJO08KXNrrs6PAI2
SAvQPFXCnzFnAypaEXA3jiAykly5xnf+HK7XbKbn+25nxSznCREFXZFl1QDT2v0Jtl+18w5YUvTq
sv1HCtG6TO5YljtmfUUyknowdE7wfRXhFHAOmtlR4Et5n/kibuuk7NFRS2iI/pnnQTfXbDBBP7FK
nHwG4iF+PnwOb9FXdGAk9gu+bEY3bSNu8E217XOzzGB1qaCMw8N66HSPp+Nb5PRZGd8fM8uK351y
8ZPrA0S78SJO9nIw+S7QED8u7yBHu8aSslHD9SXDjBwLeLaPia7oFyZX/HbcqrTOrryvAIbkiJCw
Y/nwi1pXzdstdwAq1sIXZ/fIP0vbLZHWGsgek/UnmZEe5I0qB9dom5YwGirRfDCun2DPzOKTOwaz
C/NuP/swwH5DDnUz1NuXFu4+1elJ7ccGes6m3CRg6w4j+lYUHmq4wWa04Oh9OuCppsi9SflqnDP+
I6qaIHHWA+AxTVhBx2kk8RryDgJg+zZJ7oNESt4EoOpcZcpwT682sr2/MVPzTv4KcSoU7whHRLOT
Fpunkp6kiLERIlRZBSbGtcD7N0ej/urmBNTa96rIKYDYq125S/DGdrZi+eUrIslZiQUHnOMpaUMO
Uxzi2OVM5FagSajrVlJ7PALdsgkRift+Wiq87/8xkq7tiuSYFI2dU4ztrk92E+N1HqvTc6RBC+2i
/YQObRVBjGxWuM/LSiePUC1okZgAn0oauiV/6Xsivkb+1qyHcB5gylHNWquefs2rG9EZUzPGIfHe
Ji1YMd77vTFj/BMbWietQTGpihnwKgHNHQnejqrUKIA92A/Zew6zcQZOOxaR/YoNFYGyE+kTrvQC
PY9VovocyagBTLUJs7zM5AV097wQ5N0rV+1pRbVMtqdW3fR1XYas9lVOed6rRmjd7iuwlQpVVblf
OGxlgubFnIdLvQmyS/uidzuV4Ox65qp1B2s+3JKOVznSAaHPmYII5SOxz1gjWnls11D9NrljTnpC
mgSLMnPJc+h4H/FbbhnWjFU+m9y0E6be7WwsxnszE2/UzAod4d8Jb1MT5m/g34xraABH4LijAdgL
46h9aYW6bSacrIE+OhMT+cqYIuLW3fwj48mv4/tLB8RraERNZxCPvVV4GjX048ItquI9e80fJLh+
h5AR6rhl3I3DLVC4AQWGSrGKzQWFMstukgi7pv/FVPiELw9jrkugtqpxRoSfFFfAJrNhB+WTf7Rv
r70FaizXWmXSBIBoJv3wP5dqR8ODWdTvZPWwubJ0WtnwW4pI9lErNTb4P5dIqb2xwJC1+BidV+Vt
JxGdUuWNvfZjQKqfgUPmjWv82ZE84fpe68dLaEj6WyrskLUFzK5Bce5Jjn/R51xP8PCyR/RcKhX2
XRqRol9keh/8KurVEerTCI2pv/O+jcGG174d5U9kXLas78CQ9HUNma9cEZfq7Rq39n/hDFIvqflB
WX6hj0ZbJiUmIRVRKkqyUPJX/4lNcSKPQoLjDp4HU4CWU+UKhyxHDBi1nhuB4ArmfmeJ0w0vLT87
bpJ37AObBeNjXz6lcawLynzH2BvpEBPDklQNMKYXKhvLn3uzZb8CXzxdD7RCyvscn7JwmzcDOGl5
//QNkj4x+rvcp1np6Aij31oqqRdVyW5fdFWKV70trS4J7l+yNO2RIYVm+IRY0Pc6GFFsg65iWLkR
m5cbAjoWL1e/DATKW7N/2z4kkgaG1Tc8Wy1onu85P25gI4XiqcpbGDGN5GIeZtozR3r7hiq9FI1+
JcxHIJnug7OUCn/I/VRXAbiS8LioIQDnb6vnRqNvKrq/SverYZe7+FA6JoMO9dNihkabC6HH+uD0
FwcR5wXr71IIaFLFY/KcloMvLYCidkPlGYsrIING0SwcCm0wvGm4GZJ39q7LB/HDyPggHd3TsRYz
nln6yE8XIG0x/PdDzguI0yvrpQVY2+WKIHh3ALnJ8i+oBa5LEuubyWhjyGBOzohrI75L2ZlBmfaM
I+qbnwwniorWR9Dc1Ji02st8uvTvnoYUygCspEmJP+5VAtBTq7x3K18Zb/0TmIasAoGD53dp1UCP
2Hnt6do8Hgedf02mIZgnfG2eS0orxfnESPC2jefg81HYyrzTUfub55tXlGyi5ld5OQz5AzAPK26m
ztjcetbQ+uQ0dOnPo0gB7LrjR3LCUKLfAK0ixTUltG36AdvFiz4MSsmgUBS1gKGzE+mKvLdLkvkk
ifedt4nbyJc6Cm66m9RBjOlArtc9m7o6GPc+PAxrWL+p+bEh3O1sRVN89M40RjwwoDlwMt9ECgaJ
yr0tu1kiPpl1FqTfsUrRMHGXR4xgx1WRoRM02IcgolU0cNG6rWtsiPWJrlf7wdVFt4dEsQ5OzfT4
jVNdF0LVW+KPRI4VoDTtAXfum3Yz5GxnJIu9viCywtaplDzcg5NSOdDu6cW/Po3Jw00oPlZ7aDDb
QodbZ5127nDtoffxskGUnCt0pqhnMdlB/wwxV2L0L504DJw2Was302GDwIjKt3xHdAaZJ4XUoSRQ
QvY9C7li3Exh0gI+z7imsDWFb0Jcsv7fjSQFuB7sRfWBUOaJFOltMHx7q45bSEVoAQ6F4CEYM9t2
mYFMSdl02+MDgD9jAHR9U9ysk6IVL3usAq8kPf0zmZIY3YEZsVaDOM/OLaPPntwqQ/5qa0nRF3zN
ndNEpXAFBjpqbjJgWHbtH90/cbj0ASG74aN0eu7OVZQx34wFioeykEywRRkFFc8ovXxDvhdNh0V9
PUcrDfEwE2MypLg2FK2MZt02a/g0rXziKvaBtQeKtRrpjpsrm2wb62m2JywwCv85qBjHO9akvh5R
JWWS6IDej6MITckj/mXoUgMeC3rznP6XxHi+hxeclLOstHT4h6GjTV4LehikGQ2UD/R3V2adaEHy
YP+/4skcOtfXXGO2+aHIYafdUbP6Ngk9OQO5gVXrUqDeVV49tQ0IDracj/kF6GIvDNyQ2LN5hM/n
xCvhPhBYx9EOzl1KvGauMj7pXP02dN5l8NQRQ59kkhN6S0XnIhXa2zC7AF9cPDRZ9t8UtLmOEIhG
XtkPlDh0jFJk9/FGthQ3HIOA4uw0IkEPVea2kZPk5QyjUKLJ6SszEIGF4k+McLxHC/LZnNK2LtI3
A+iDg2+kKE/fcTOGlxuqf1YVgior5BjURNTLnThz2aUNid3XUcPt9O1a73A0+bkzRH4bNqSN7x54
d/jE9Z8iJZL/bdreScgKcxNh4bfH6F6Qt9bpq2itvoPKQVbGdep7wl/fYvLw7Dhs42m4JeoPrxh3
AesQYdsWVObT0gG3tSXLdQF4/wXY/hN3IjPG5EBUkgoxptTdC0rCTLkvp9lFaa/EfcYqMpST8590
FRMEIWkQwmobLf5o9WMw3ZML/0ZmrtEZi7x36uefDqyDR61D99T6Inv+ACBjTaDQT4VzENbvcl3N
011HvbDGiRT9uFtyYrfJVmFJOVo2o/sPhDk9c3ej0nLzTkJBM9nyqwYYgipugylGo7VVm+3mWOc+
XS9rWrmK/pk8JCL9Zp2mn5B7wHtnNGi0VjBS7qXQQRwQdl9MIdBWFchmTUI0lWE95K/pPMm9GgXe
I/FjsDNwTQx+/pOBat4JYkJywqaP5DxvBKqc0UUJigytxohunKqH18pppENE6eaDFXSrVlJYJENF
BqYTehVKe/PYSOXc3YgeqXHY2SbeEfGYKLhhJgKRk6IXaF2PkuB/o4qfF7lcE25oWsOWsDmYm9Dt
Ta7nhSP47MHAHqOp2yupQhh5x/ru9DlsyvPb+gDD0jTGSkeH1iclSZOTwcvnkQagl+5k3VhqT5MF
3hxDBkZStLko+4aqaPRIrIvQtAQbHUugosGgQVHWG7cjtd2fGbiojN8u7GujVryePW2VxbDZx4PX
0z9HykgGJZ5PEb+izBngfhyy2cmg26Smym4He9AIWfpaHx6EdKSDh05qLxFgUoU4QGTZ5DdXQKwa
dNX7OCxZUp2P4udNewkPXlJWOaq2hdmcm9dhRGZetMJfy1C/eLPFEyCGrE8zr2OARAxbhCBvfWbb
XmFg1nwe/n9cXHU2nVQ1XDFNubOaXHmUHg2KE404x4q0SXdv9JRV+BfnwjWhuZgcVfhAUbwgJhSc
FN7PSiAwMGjB2q4wl4y9aBwP9GjAPfer7CyBDwyOugwXqdqT/GJ162l4ZV265EkUKKjzq6GIPKO7
ONv0afMHg7w/NQLRwzCAx1Lkibyn1usJfoPtNUPqfv+2QK5UlKy64BHW4sdiLg8epy1//OpAfi+r
KS85skILNHzhVBdllNYsFeWvG7d7KUCBUAga1yCDMYax4Vuqh4mLfds6VyjxNhQaNKEi74V+wWIC
qufosYD3G6SQ/imwTVX8iTEtADO5aEU4DNYmHCPYOJ8aTaVKQxtH7erPO/9hno4TPnRoEM8bbPN/
K2eOmpnp4OaWkon6MyoggDZrR1YRaWuonpiTfYLJDEJdXGQ7tt5GWvhIFr0Td6PmW4vUkwCEUPuW
rdBLKQ9/9SpBEqOnIVvea0GB3ql1nBGnE0FgA/+CDhYyIeP5Jov/EsQp6DcNorX0j9te0ZhrKHJ/
nEmQ3zIbjTUks8RerzIJBZSkZhAOJxBkTRSdH2+BDjFfoVuRi+ovVLgBaWYyGh1eKiPbVJdMW3r4
ecLQ9ICQq7ilGl8HGiwzYad/eRFRjsg16zp5+WdIAAZVaR4Hoa2QFFv7Rdjhp+7QklpkFtawI0Qt
9yNE6D0HEkWGpLrgisyVVbsoNXvgxozhZ4QcV6uZAm7/k8jSXJgbx8No2KoUUHIF7X8tGJiY+Kl1
diIzdpYIbSluSxHtAVLsiG1KeFRk8vUTl3TwcqwOJbZfPMmru+LM6BnlVnlFLSbQebsA2ylblTyq
3kOwhN601MF6pcLPHthXBzfxmpYYM1AR6Up9T4CEEJi5lf4LqbBfW2/nARVqIhHEmW/qlBJtDtwO
UGyUYPA73rgT1EIPHOijjSs4BLiG4Ip+iBJCHrcfNuc+YHzJ9goaRnFBP3G4Q3oDpaHWJ89KVS9k
p7Dt+6lhB8XoV8LoDVJurFi7zbo1SQEkcZj2bdVtCgL/vIcM/fE0a+ZQeVL1KCEoJ/6N+lmqIOFi
MkE5LMZArKFSu9oNBurq3qSpVhbU2xby0tlhbqYHBBZ4F0051U9St1aun9ZW2uSuO+JQQfry7JPk
YGBR/m9FL3H/8Jh3Bu9wEjPgcy2WwLCnY8bAwbe0fkgs73ezZXiZMSz+aWUu46xySotPluWT5pBE
klreNADOQpqv8X4wyHlbSI6EjmUwLDuAjOOno9DCNk14m8JyrRMu1XwGcZnc/yyDoozuau3Zm6aI
0Gb8BfQyGodWGSS4EYsqO2ghe4vuho9wYx0YWf1QVzOwhOZcAD/aKq+0JmCuqCbffwCWoR/cMnQi
tEJeCvai4W/fS7IsIjNXbDUtkYi+zEjXZyQIcjvES0lDAfgvGaRfRS2moCTyngBI9Jg/GbLEZFOY
4uKxbgg84Nm1pL3AFdnb1cgH2VRt0z6RDGk0WquVjSt6gcYWOuv3NHsHMwQzfJSAYmpEh/xWk5Jt
XqSZyUqSxz6XmsOxFS7z8dI6z2agNJo7IaUz5KmZlKRcrrn9scnFShWIlqSkd6q3AYhfhPjnLSfJ
oF/uUfC3NEc8YHkUVN0+Gg+VN903qnv92PG1oKyVrKfm3s3gowc0PiOH/++2nPWtKaQ5DIpk2FqH
ag1gzyhjDJctrjBq3i3LeXzFjR8hNn7JMaNNWalt3BrTzO/NMHivqQDXt4asllYkOI6GOiqgRHyx
hGSCl3r0fJf027Pqi7CjfrY74zNy2XAR0a1t4g3MrmsUcHQ0SzrANFqGdjlPZv6NMd5zDmc4kfI6
R/gqqPKkMYXa2ifXYCe1XXSjE29ZDOSIYFiLgBM8NqVtXpDUt7Qk9RSVMXEva3V7wFK6E0JkVa2H
NJ9bPgmmg0GzdZOfB0qQX4ypIGjTWmtg4z1uikbw0w+IZpfEO+vKWrJkZcLBtp1ZcX4Lh36e9DeS
LuUVZR0q7wlxnmabdUuA5GGZnbSHZ7XIJwxFJjzFmtWAlvR2Rdu/Olh/UC4ELRqcOPWwnN35SMuu
JCG3am3rf8m4Fe7S+u85pexmiF4J8zbqEX3yY1/mZiwmHvIv2zwmXvyTM8juS5Mos9zY3B8bumCL
k7nDkyoHOJ+lWYyIZUgXzVRjmvvrq7OmdqHWH4+HPh2JKn4ZD0knH8Yk/TkiX1O3/uyyR0wd2gMn
H4vH2DI3YEx+rD5KjTxETRan0bO8jaUbpTusw5FjA6svgY1/8px941UyWE21RFmLw6dRMYIRDBBm
QbMMSl6C9xhIfIoeUqP5bXYUJ4JtveUH3ZMIMABH10PTGukt1p4YIU3cgvj0LjzTibUUbh/LxuZn
5oDLMmRJMnNzPByL4UqBDj7GOYRDO23pTR7no/5qwjCoKxybHNwbBb+CJqnMweqs4H7knIuXVwL2
HU1efyw/yMc0VqdQedKv3TTn/x6szuypkoUtp7+Sc/suEmYOfSDNPQGyKVEgFtj9kaZPcofj4us0
aC43atXjlxEzbBs3bnPXWlEsGMGecpqfFEs0u5Ss7zGP59a+00rmJhIgwxh46V9wED4FwGnJp8lE
cWyuEljvluuE6rS766yINd+YZRKThyzqVrfEDwAO1vfUOcR/mbMMcmBI3Tn3go7bggeyxzYNLFqB
vPE9y5p7NDYubqpsoQ4gCM6zd0bZojM9x8cV+a17vM4y6byUvBX45fkrtAbAgucfn6eacMkbipp0
7YbAbu7Uo/KNdRpuVcJWW1bDDNsUO3WnnYABm66VOkwIUhr5sD+aT1eqxUQrCo78/pzdj+iAc5MU
lwjXRozROddr8yZOAMCobX/CiAT55tlXoEJRHKvLrY4hGoVREpuSyo6XBWZ2QQWeV5y9FcyCaJsu
nxjru/Rw4JoB9f2NpKcpE5E6sznuXQhGuQEBqv0+7K/HnO/bblyqo4gnI5JX3h4UAzO6ieXEp0Zj
+tbNCsZG968I1XbQKNlnmcP18aw+Wo+AHwMQXQ0dpHEdhfATcn1AcEGIp0TYNWIxkgNXGQOkHA9Y
Eiyr78YYEdGMXfbYD+otA4vJHzfm7bCVsyhE9LgLb/6Wlxstx0sC+0HKpKNOtrTETUeqbb2uz/c2
OppVKk99/YwAZD4tFTdpPvrstuJiJwpJa+ddBeVUn/1LY1bi7vwYSHBTOzQderixFmOQSyp88k33
1Fv4bhW8qWCyT03wxHD3jMiZ/j+dDirsN9jMPycY0ntw6lz7MgaESDgjMmAdIRdZpCyoGNDK7DWD
wEZaFBUe+Q3zMlkvmTjzux4hYXgB7bguZld/wdSDr5DYt5dsyGyCANxGdR0zfM5olSdGebZzmRd3
cCIklFHU1PO+Bc8x3F8hehXxXjFNiTbdCyTdt04XStto2j73qzmExI/ep12M5uAiU/Vi57dYRsCV
x+kt55WLMgFktNjVpPrGL9yjdusHdCeoEv5YnEmrEyfc0ez190hyTEQo4b4E83kh22+Ab7rPOvAn
saXp1A+EWTrZ84ECYNNylj/BICrYpfxe7vQgIvtqA8/2I6Wzi8lEupvd7FvOSJsx0dZKwtP3qsmB
laUhGuA+vov2fnUtzGxOJAq7e3Yr5OYkKN9xKAu4W72grjl8QGghua2gRC1zObPpMVOGTw7LJ9gg
AMD4f7xAGCiH66oxKRyy7ZMzVpwXffvm1Eyk0x0f7AXwKwwoSMt/lnyHM1gZv1rKB5Nm2e4yVsQQ
1tcBJYcjubLVUd/VsPq+v0ykJeZvVByCcb/aNsSlaZlwRITnmWYGz6fPqrH2HL6hQkpLECtscmZs
fkmqvGbw7qVDk3VE314sHJdKV7CNWPskVNu+2sffO+MtPWJHdbADsHkAGR2jO6HqD8i7Fw+XHG/P
WN2D0a1sHoFp7WnnuPaDmb7Rd8rwO4AVHaDFU4OsJqAKkj41kQO9bvrH0qhYawCdXvhVlq/rjalh
6mC92p7UKssBe09Nvv9pgO4lOZu010R9/Y38ZPCd80xGND9IoOvTV1uV1ALXeYcF4vB9u61ZVTxh
eEUCHyRylxh7qOQaC0WlYDXsriewtsHSpoFnMyPeJLLvyFK9tGck9jpk+gT0vI1/FBpmLAO5F2AU
6KS/DE8b8FE5+MnZLeGKe05nAS2X4wRxMjwQL2w7BQAsdULaRpo5ng0vlC3t4I3hHw5ljE8A6vP5
2Zjy9XTO3S2I5zna3BIGWWZSMxeNftg05o6wOzMQ0mw7G4IbymfV3yPTtMQ32kO8ZinE0MDwdOLM
qUCWNo0rzhH0IHWUMHmtCFgCBllqVygtArb4lUWkBLg7rukJlhy/YLVYYGgz34xolfqpxZpmss/D
8F1slxmqnpBvCodAdyJpvOYQQs5S5OWFnnS8Sdflwg+KP+llOw3+tZpCKhCDJkahWL6CkMbyWbSE
gE+4BwwznBg5G7pg6R4EqMZ6G22aML8QR2zXxJn13zJP81WItaftaoBH7IZml/ddOGObEHrf/4kp
+2WmNH4V+LDYPACAYb8sdFeG9p3HqctLs3CJiYL2VoXYmGC0b+t1Fb9CbesaFvqt19yJ3gS47dBP
mQ+p0QfXu3TIG4cIHI6wXu4Qj97A4Ifs7gayIREH8Z3ti16/Sl0iSe4SXrtRZLn7AjtJOq9d9EoI
iGbumTIi5OarCt1IPcNcKTx2hIzWM6G28VXnMjuGN/KDOVMgHVa1VX6oLzKqRkyvpn0/x64Tyw75
IBxn2/oSgv2tMtixpWp97H0Daf8hRGvx4VJ5BczebXhSwP1nqODrd5k2BYf6uJmOx2abwnYG9H3E
U7lfCijXWr0+cYirLecuyO3P5blrSSJ8P/X3BMdIUiUBoZD+qqxcdVD+QEPCplcZKz/nda7xRuz9
oHqYLVTgIPoZo39deQfLgq5CSMDk+LjdgD2z19Au0BuCv3FGZEmrr0xkHfRa0r8b4ONHky36v1VR
EzKvveBL7XRwu3CCqpovX2TWKft/uzWIeEs/OGLdFY/A0idRSHBdOFHAt4aZRmzORxyecHGuxCoM
6gtjYjzPsXYBu2NxEdzHzrfsZLYhVIO4fyMrMaSzn6uP/zfEyj2yPy579t8GtQdxzpNHWiH8jiza
E0te0Ccn1Jn5cHS4ZtjZmOpTL6i/dXk6cQWHy+CRMWbdRxQx9ue1eUrSEXVHUpumS4c2Lvde2vhc
MwK01jFV+l6UQDOuhYuNHZ9UZYwxzLsvGNf/rjq+vibg1z1NX0vHZ4VcP0yT+DhrDEKTOiC4og9A
gh3cMAmrT8onrAjYz9Vq4Q==
`protect end_protected

