

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
kNSODHF2BA8phv8L5aZNyOOK56HCcQ5lgKBxF8hcTzwkWRF6WnOKZaH0cAk+oZsvi02J9SlLLySq
oKFSyBG2Dw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
df+BuhfNWqGLyuHwX48C4kdWet0FAm6osy35ZO6nvLm9LeYvgiC7d+QWQpEp/leK8jaqvimQleVB
qNUNsNTBZzVm+VZnT/+N9fzr+Kn5brl7DACKZQsJ/J0EK++GrIymGQB1+7LWFg6RjvqxHctXSERU
pIxXjKUtzcqAwrR0kd8=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
j4klfuw/RrSoDKuTiN/Si4GPF3r+1zWV61wAeT879HAyso4ajbQGVJETjBzL4XBayVtdsViewbVc
n3EWjppKn7DU95ziVUsafFQrG5PCVJ8TPZUJisZwRf1u8N8ojLSjd7Gi7vpDvGySyTXx9aoOQ69U
XzJmTqPAeaivz/FLFyjHWzMuc078i+06EYa3j0uxrNsDH6/IL5syM3QcJV3812LlPGSBhRN9Wynk
J5AcITSvkzy/dqcKICGyxp5ubBr16BEoG7l6F/VEXvTJm/kJnHW75YZ8OAQ3I6icKjHkLZysnDlK
KEU2K5X/pkwYnpID2ogdwsEuEQr/xxo42oEmKw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
AG9C2Ti5ZMi5neBsWpJ1qwXbrUaWpaRO8Qn1fL70JVZk4SiqmPlFkL5Hz8GrFfE4eBlngUFZoung
TTZ2IeyMWjxhdHHDVda6+BqJtPiX+FBQnaCzRd4VBLDnB8KUn52eheU5F9XtqqkHq+oJV3U19TRZ
Rq+NhUtknFhYrHlVXfM=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
TuUXpu2xk+duDJnZONHfYiEzeCuzIA9y6Ut5Y0LAE72Cfiq+aIEHs4lmSaypPxj5+E8SKfd42Iqd
iKQPBy7GWczcAr4hdHMLEortigKfhxQvyiAB00CsQyuj949i0l26Eh+7iirhYh907kSXNLc4JeDy
uXkHZzsX9mKBsIZLMO2TtO0R4ECsHQbqo/hSpi0B8kY4ucdqtZfLpEsAJ7G3XH1L+CD4o7on7UAz
BPPpoVV+VIZR6heT9EgSZTHhg3uYl38G0Ezv8g8s1cbXnSuowx0B9mx89vkctBzRxFOLnzsFdBr8
DIKQCrHZfdOhrNHz4ZkgOrKjCDpwEkMA4ATVfA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 26464)
`protect data_block
/o1hnqtYZzVSqeA3QeOL4UYig3DsxqdL0c052Q26qnV84M5MTmdNAx8j2/yBZHq2fhqYesgZM6An
rj/hvd5oDDAAI+fPak+0aJ44ErzIcmqvegkdKPj5xuusQ+P19nb5gFEXFBox7KmHKpBLcMIzhnfU
KechdOEeCSIRxSDmPv895qy4n7Nla/Ls68BsDA504Mz6tWKX/VAJOxx4NisSElRsQqXw967GfniB
rETpIamI4pjKnV1sFr6PEy3vjJjD/XuvVvEmMG/lDMnpqG0db4OAYsV7EbeV/3qO/TM7RXlWcJVd
cGp788H05ExciqmzCWNZtYmaKpHt1voQm8QKuouBXbc/QtSJwThlPmZO4sJ4TP9I25ftcwHBCQzP
zreZGRKVk25yEA4mnkLjLLb5TAAHAiGh8/M3Lhu5XKsaUzWLeSsxmM2OB2lgAkgpY6YNz/nARLpD
YXtcdVALcPNy1lsI7OL0BRhIsjxFtWMxDrtKAjJLLgCA+C5k1T0/qFXvNzhbEm9/FE09p3oSX29r
/kjVb/ClLxuMgx8drb+gIWjoyBIQ4v0mvz72XnpJPfj9Usv/22SmICTxYBpJ7epJiCPYZZx2zFIj
ivdZtmZYk3g1WFRTA9Z+tgqKeOORHYKDNXj9aJXUVjFSuQE4OdaoHUwv6FZ4xSx8pbYyTV5HscWf
hR3xHlYo1O1mLlMysaBqvUfmV8YRyK6NInahRdhD5JJ414jraQZy0kmYtrB0WK7bsIBzlezWXtol
pejHJjt7eeKdMI/tLIoDzDG0wDx/kdbuA8s2Z/RrJyOduaR6mwKGK1fdBCn6TxUvFqOcQbqu0fxN
IeFZBmd8ACT+IQnTx0BnazXz2iuG1meAdrJY9QI8nBzNY7D15mhh7UZMJLjSuLsvhTCPKCprA8gK
EGjuCmoGADpAJCGH85AJbtizt91yOZmirfdDkyPN8i8E0oOYq8RYV+Ho6fFJQ+PhUVlAPlVc+srO
rUh1/L6tPhz0ICRO1pm/0iwUPoAellq8ylag6eaF1WDHNp9qlibjNx5SfjEIAa8mVx52zTxZ6VBC
9AnukkDqC/I6ukdI0J8e1DORo4CtGkXiNnDIJMHl/xmhK26uW10/M6onzCphQ6lg26Ut8f4Zh/ht
veXGhE23Juki47OGyAqVK3Vyb7yZ8QdfG//UCU1P+hJUiGum81izF1+mOf8IbPBFSxwu5K96sOSA
lFp14GasklhY13dow7xb3IA+rRu4nyt3m8nGGDfwhkMzIKQ0+zCiDYE6zIK3C1w6aKYazop+3s3S
0npVgd/oTUOZWbd2LVnR5KgEpz78dDBOooHR2Wla//Oxma8M9wgqSsSr+/6O0aYNVvfI2tnpG3iD
yRuA8DEq7rp4i3iYCWfO0f+UNky8unzcSWqBte/bA7fdM/RcEjgIPCL+H5vdvIZGq11khNMTJftr
vTIo/mVqVM3jl3yHZ2xcUk8IFHBiLn82wohAyxdRuM7luhOyXbqvMcl4Qhh41B0dza80hHx7+Mi+
Dpdwc2z4LDrcL2/6Rdbz1d2fegWo+aXYUJ+DoNBKphRG0ldUkMAArTc6++RAEddGRA6KyHDRI2+N
p5NDLWdV4i8DxaesIVG5ElG5z9rbkCNEHgDO1/2+J7xqsN2c0KSq46cWYGEpRLMK8fUJAtDks/LW
fPURUTeX2lMM+N5Z0+JmoSSJJlk/MB+bXBMr+PSc+80icYk4YvfoBZynuLsuKpVbEQPIsww0rxFA
9gaDX63lvLafEPU+TytTanjZscYywXCXbeYE6Ve7kIooRtKH6d/rD8R6ZZgZZHDMe5RwfqEm70YE
WtCMqE8g5+IaeAoVy4LnvT2DKmlmaMw+2RnaBL5+L8Q7YQmsElYVWH6GNVTtPgtvtumv/eXWMqiq
deHLfqkXe/ZV827QoK1BUaAFk4KHypRsXLXFEBxZ+ipHNaNAXrtxERM3eOB7tAivIEvGoWYheVaF
4ek3YAw2E2mZj+jc68ybgY7EyDbz4os8HUE3Vclq3cNGJ7il/NH5jSk+A/r37MtPWbz0s9JsGTi/
0ldjwHc82gAeB4PHfctNE4nEgKkoQKqBf/CXiK1PcVvINsQL5JX/KlJgYV12FOffty61BCQQWgAc
1c9LbiCeaE13hODXKp7P3WkfliJAlWctxfABium3rcUhv7xaYQn/fEzPDa4HPP0rcCN1P7DqlnE8
MbO58RmGteN4mhc++3pdflEEAa5LfW5TuBV7GzqF0Vm+x7FDpblhY6oF5CJt6tUWId1JGX0KIjF+
gE5HDuAo4cb9SpzYdJcj0xuieGTn6aPe5P9Z8vHDX59kgKZc0VbPxvnhib5GUNj64A2DH8nHeivF
/XzYiFtst3FOMrfd4OrSzFTyHsZqYw6svGFyWGi8ZD8tlpwKlFNDgD7HZ/6CeTpnlpggC1wG2ykz
imhbV206VXbHdB/75LtOi9G+tUvDUcYPfJQI5SerGuOg5Ud/IRQGcL3QNFjNsFCgYY8agUomJtND
tfUnawW3KImF2oHMSBvXg2eA8YjdM2XJ5D6IKr0SJ0wkAdT9ZzYA7eOCpEv0B6tLaZItcp1+lvIP
pwawwrMUU08a8b65YuzSprv/S+c3TuKuq4VF2qVjWS1Jbz4hZDQyezHGTkVHviEDVLr2IRTHOO8V
5dpygERL0wdtBxfhYECAnuVSxJaPCCV79ai3ZGZjRa2pKJ4d4MiNAnu5dDT9C+CiauPpTFWfuupj
+4FTIEfOAUnhY6kscM7f0CHKr89S46guV4nf/9rgWGgEV4dhG/vamOGPn6zwOMzHaJWNpKTPFAu1
4HpYz2wLgFPqooeLC1Hn9Sn6Y7KOzjZ7KxbQ9+4ek1p3Kxf/yutASCSJho9/C58aiVkf6fd57dKK
BI+bdx1ioNPovgwlLd2T3jg5DQ2sfAXdQgj0e5zCjmr+a6KJfdlfpYWkErlwd3Zh9+Suth+uhEiU
oe63Qf+oiPphQj284t4nslL+VIBea8FFhm60J3WjVE/eYLNi9eEURdAOua0P++bgPtYZmKp60L5n
OoYAq6WDpCG9mT/xti4qJlqDfm/f99ZCScPIW3e1JozrdIfWgiS29QATEAU9qlvVBNtQhGczwfMJ
TIGb1x6tlCmu0sfyqGxOxAA4a5U+vsjvsoilpQp8JSb/WwGqcfeIENJ6Xuk2QPIe5E1W1bGkQ8J2
BUZK+CHI9LAACbyqrGM1UYbC3BxdpnXQaEsfvEOFqFtauUN9xk7DAN/1v152fgGzCpxgcEaKwrtD
a0WEhmgEC8jFxcGKWxf84wEC4PfEyNZeOWvYNWSXsLmhOVMjLmxDhq1jFflC8ZJ6fjs9NDAxQr3f
LVdD+xGbZa2z87bYgwISwBFyH41Wz+ETwuqbzi0jGecTimjvn0gpAGhwvnqjjPShEC3K7HTfPZX0
UGJmYCim6VsQ7xvm+doFXO6u3Bsa5p9+vzWKOWKKyyAfXjy9tNUucYIUT1X6cF1Acxe/gM6H/zsV
eRiWaNMI+BkAlFOqzVAIszU4vi/j4cp8jDNnDZMChkJHsl0FZeR/qiTMtOEsneiEWxehOcuJ4beP
So0xRPlg6pSnxMF5i9OS64nwN0HCV+Ff+1/v13dmSWOf6ylRF6RDUkXPxbKTpjlIViOwKnBXMsvw
WIED1CrZ29iy63g39MrBQ4jspr5Mlatfh6OIQ8cn24tkg1SvPDpNPO4C9vbqMIXfLrZ/6L4vNHPQ
CVGYbo4bPUYE/ADoGgit8b+x1e9YiuRfa0S0+MGjSHDQPbw1btUxwubs4XAD2FrIX9RzWQ77sLOu
Bd/dju6uIHIxAAkHbiUzepvV5WYibzFITcVOHT2ks9zwnk7z0UFrR9caeqPMlpBlX2iPgl9/pecB
KryzBQqW5JFSWYkToxc5Ibqo575Yiyvk+ZDU7YiwXAJaR16ZpnCikcwPalcVaXhwChdoUypsazUg
5V2+rGhHnZYRTuUA79Fp9Uyt1GCBAkydauwKOljV4kPmlgV12V8MYaAqo0ATh6agEj7VulYZMv7Y
+u3SB+SLo+/gG0Bp4MoSd5veOPZL0w35++0xMexw6CtBMCUGr1bO7AxSSqMA3bpJjUV+jMAkXRVz
lULbftF0YHtPzZfeIfzTILug9bnu9mARYP/MWDqMqux9dfDwe4GqCyDZoHuLbxmL5Q7YTplD7Zqv
VbRCdm+qL6wA+HeKcod9QVTogulaMZ04vmQ6iUYF6v4kujUO8Gbm2Gz64V83cvfdxU6v5+ZRrY7+
Vh+Byoqhk1UAyw1OOdrmVk2WSlLZL9c4WrSyslEVKatpTiKu0T7jBrusM+jmx3HA6AxXyBFvZUSC
pBInzuPHg7eB4Q0QYFM57aTfr6OBa0fKmLLVGLL+Hik4RTBatd+teFBqZ97ZoYYYX+y9ivQ2NPgf
OdnQ/k4GyVNLF5osPtkLikdb1JGUEO/DSzgSOR7KOjpGTqo3qIDjJ8VckAJuyquUy5JLe/aRocnK
jC+Qjb6flhnYmrE/0j2Y1GtKrMp0dg6JwG0UNZA8Tq/1L+KPiJyFu6zuGf0X/roVFYer0dGQPOCZ
SqBpAOM9sqzpiUni8bldmeqakRJ+/Q0sVV8TqyMSlz4S4Sn/LeHRUKcEU7aWShSYTNyV+/AwgUDS
Yf4xSromEALpMNLg7VicmUXG9GaZYr36b7IHfartFrlvN4pIdrIe6dvZUeaBtceMA13muN3yCjER
Q2S00r8S6jDmxsSqUflC+N6v7tegheL+MPCvfkRf3xUJTMkOePxsrUXycAib37Ugjxe26SvmZPbM
vz1+k4q9GzkA74ei7z0fXu4Kwa+9rDihQbGcGUHN5OceGSikHYrOEA5koIyi0GLXww//qNHqVVmA
NRQSHMiPSp5cfexddLEI1BTmpkCj+/iuuzBtUAvici9SF4xhcLgqQKSwzAvXGP7E3jInE5u0AyJp
SWInLNMZ4bYb/hgASuNwLk/jPjA4UregeB3gV1ZCPnT1WJUTJ+F/Yi6AKFP10EVptV3/8zq4Vyy/
MooiM7eoq2LbYbChO0Zwmcmrzm7gQZ8k6PbzzhgZXWpu+17EmuWf13bzTFtnODLK4tLOZcV58loZ
dOvGB93JG7B3CyYLPps0fosnIke3WAH2s3JHG1yi2GhHIGmDcr/tyiH86GTmiqx/eJ0VqbE0ySHM
wuGbcMDlAF34oOQ+hIbIbi1/Czekt5m7r9PUqrNJPvjDAEenPgXnkA4rZlOZQJCtDsY72VCiRpVP
7/amxe6lSKbA+2uEbsENf/nfSPP6/3XWBWu2LDAvMfbynKk8n1v1GACyJ6uxMQqfV12Inj5nwrde
ELcdlcI//C9wKfkNxkFEaDFYAOuU8THEMVP6C1/nf3wGk5+nNxkKzbhnHDpHWOk+B+swvKWamySi
laGy/QLq1KSJG522jGjdYY/MWybwMqqFRyr3RMFvqX4La9FyWHHWVxo0GvMDQdr2Gf6UTPKqVoW3
k5xJ/V5FjGmomLy5Jyes1UkNnxxSjrBQNqmJRM6BHakLKYpLwFtFG14x7nVWPv3Ny3RLTg8rjGE9
xs92HbFFp99dBCUgGa8UJFflX7/oVBIaZZv2tskKJ7i7xZrkVRNNDHDmRXez4oy8LHUFMzUp/Qno
iVEBnPSXWYSRMlK2RBZLPlJ7yhmCox0WXHL7Fr7idv7zDkFdkEHEuN5QunOgPeWsHT4w87lxMjB7
BTbJGkd+ticODMEpxQxbWIFs2BtreEwyGu3jQ530R0GA41eIfoBMZ+lKU55kIJ4+G32G9meJrm3U
ziFcMeeFmKe61TlFMawC3i88v3i/mpDHOwhvljIwQfP31EQKMpj5J8BjewqPqeePgrYgEFSWymav
g8TzEv0uldMzcgwsZoIovv5d3DQ//5tvJoIiL3zvEBWJUMlwFzkmXGOhbT+zH+YJwxRThJhRU2j+
MM7eN/diSviTGMlA0Rb3Ji+0fC0j3NcU8Ol3XwIvLL4Ij27wWqqbjgElh/5qmVyy3aaKAmPmHvU8
TFHX4y6xX5daG+DiZplWMQRvG3XhgL4aGtKd7B9konL0qElh9yZ/6xuosXTkj3nclyz5ie3WPrQ9
0WnfLUS9y19kJ+PJAGptb18wdwHHQdZwe4KuJwB6Z773FxNlNOBzt91nIPG/nQEy9R3ceXMZaJCt
FtbkfMmEHkOkOAjd5cIddI8R/Si/vf58KaIiZi9eD1zkmjSZt2UL7zk22zw4b0uAh05ztsWbxhB+
iwusu/Xkjz/4N6kFA7PwCQbD7VRIIj9k40kNTcmRyyh/wgAYszRsTb0eJWT0IiVqycMd4Zuco3K0
lXwZKK13DhacP7unSsgJQBkTupYqEiqCvEbxQPZEjl45/apmvY17HmQaiZitcJ2l7qI4CfUi0ulg
kdj7K2ptqZIsTjKybj0/zPpXQqDVq066CW6UdO9q6iuSK+RL8LC2gDAfTommjk7Mu3sfdM5mWQ1k
7+9Q0ydJ42zKnWBxEdDjbkq7qIZr2ksQMQjb7ROKtP0nbSeb72RqfSWqdUcn3+5fWzFHX8Ur6BxJ
DInI0s69UM0VFDl1kFqlosjVqf5xdpIvI1W/2byh76/Am4OS5w6ytzNflCPHer+gtbyY7dvNrIVg
vSvqDleHd3VoaxNhlGo7SOCsLqa4xPRHHD0Sok57Tvf9cbCOVTBRnsnSkM1hYIRccanSnzW+6v3u
W0Vn1/Bougtv+CD50Sn0Kd76vtf1Fcdt4YAW2/VqAzx+sI8FP1/Es3/DkwgY2PFhjIR5XNIA/42G
3O/SeLs3ut9KK5ylxSSiQGVPO8qBt049zDXHtNli32xDaLv5rA6o2u/0esIQ2MQ8li4akmThMro6
nd82ysuCf3IU4Mq5pjctrBRNsjlkAwaCGfojb9CPIMA99AJU67XeRWb93K6AI74RZbh7JbhhqoBv
enauizyzG9Fn1vlhhun1EhXXFQ/DF5On+EOjfM/xW0ENVqQIDoBpP9uR/vaypgZ7L2U3LUGN11DE
dn6QPKV09KAxeT4WaW5RUT1x1UeIK2aXV6Gmrzru7OGOvRVHbf7ztBZR58Tun+wfjWXxEPT31SdC
MIFwXfvaJhy820RVewkSstTB3AHYTelrH3mVqW5BrBNxdLGBOiKuScho4Cd81WvV+wZnsv9t2p6j
ZdhOJEfZaXARW25CUXG8u8XdhswsNT6W1ZT8crWBw2KayTrVbZpN7C9XTMuU4d2De/7dgQHrHrKI
3dF8Gn9upZUxoJ4QH1KQgATnvQC5hZDfxMC/3fMKqX13o/C+h775olsx932Ja483woGIMUJrKzHY
fMFedYGLGQY42cXREhnABvqLZf1pBK20RYZzSAR9mrb8YJi7b2aV+8ROclY6amSAFLImMsO6ksnt
bDCBjaFFlhe/hE+NZoSPJOS5+cetRvpIUMdyb8yJbd3ccNLzm+n2n/NfpyS0NY7rYFCxdVCRPP99
1/AVLncX4z1fZU+Naj6sir2KUGBLXSxsPDI57V+fHoBtXwQIX/IOqOvOZTZ4VU9pVburNZTiOJiz
/orf61ETkYPT5UZaf6DjHTUcoSiPh2ezc6R8saSjtHStJ3fcqFBFC2Sc37QPNvnWFQvyxjDoXcAZ
nMGwWbvacXAORCzoW79ya5K4C3fSZ5p2q9ab6f2NFKb1gs5n0TsLvXZib7EQ/KwJpw2W7AtbjmjX
Z8w3+f2A1l4OirLPsnvz0mcd6dj7qm3keaUchb/oE4RfPFhXkX6EJunyS3zwy8axkM2U7H6rtj+T
cfRYx4+T2ZhI1vbbNtfZf6E2Zaf9TgHc9m0GbqANdHuIQ30buRPDpznkrn3zh6GXYWvm3tyRBluF
H0eBm7uSKzCGCaGDBDQRMk54pg0SztlEJLJ2NcOmJuwHtf0TBR7s16Z0Q2IE/08sQ9Id5P2E6HZh
l44fP/tDxn6vtczbCpuuJARcHyK3roJsJXuGeJTPIR5v9cLuvWFEWOrpPo7ov/qYTWEfuW+xVV7k
zt4j74+h05nllDFGPxKjxPGbAdGNJE74YLjUwh0xLI4RtXrQ3EUc+Ygd57tc05VHijD93e3bQl4A
Ag52bPYexk9k7mqEpjzu2FcJCmFt6RmpO0idKe22VVvQLAzLVBT/jmrhjauARumOKOiSDTxZPvqO
fcgXd+3BegInJynRrLqliWBQDSzMlLMLC9jfmCs7F9OuNLQjWM3IADs+F5/MHxr+uZcOTjPaffc+
tMfrI3123asgjG08Ls8qxZD7bVMss+lXPUAKVmbB37fFgvxSm/BhrQxnUyk5Uzf0Ol11C5F1YYKb
Kwc1iu2NUwlQ2xUt5BWtf6lRZfB+v5k3eCk+8d5tjYXep+jMuY+q4ztQcGm5rWd77nhGJNXWX80i
CIZq+KKW6zkHdIjz6CosTF8AjUNhODHtADMiwzeFqay4iVvy/BtiomXKuudbs3EgcnyvQ4X7XmTL
uHB3u8BQMuq/ymd2XtUR70bBadk0HKQMMjqgjbZx0RurwhcDTlsxOcJ0YgESRSSZD5NA6sKI+VAE
ap08EpjxNW97eRWezZyvhDSJBgN+4Gnp60TMkOMIygtpknlOaJXvDll/QEyU3lI9oe9gfPrpiB2O
51BVLsJTDlKPBv1pEc4/rKWRH2x923owju7LHDbMdb0+xk5zue+FGeyh+bznm3IgB9xw8DNY6wvy
KK4lhwUO/97RPYxXW3sQ1MyGsPT009kVkhMPe3+UPmYAVWv0lhAcsXJhdPKi8cZl0rWAqrMOhpd3
FZAGNSgUw2j9+pJ6Liwxv76lfoy4AMIDKue5fs0sdPB/99Kf1pzID8uopAmnBkIuiorvLHsn6NA4
CxK67qdRYiVr86r7Ljy50d2WdlP65TIfeb29PsX8twD09fM7ef20+Ic/B9kEAn6wDZXJNubTcx9U
mcCyj+tMIwBRbLRx8n1+aJmnx+pLIZrS2qjfAI7zQACW5kxpP8DYJr97t1O3TsxQenWDzprrOeS3
VwFUjQvhicHLnEbKUnrS/+6Ea+V5WAWiGscJkFvAaJwna/tfKbjYY4vArGEBXbcPrUtrMMqliZzZ
LNSkDlVFEIaC28+WN80HPM0LIPqA7JPYnWW9+CkA+KqCAsf1M/0uFddOu3OlQOl5GaLj1ngwfykg
DP9PoKpTwumBgoods+hOBj7onMy4MBcsBSoLLHkpUkTTsXSyeAtcYCj2oIj5UnVSFUVOduYxbqpW
aM7O6tplSa+cSQ3MnPh5BYcEjoW0lH6gTDkV5e7AFp5BrjYojzMnf1s9WkI0SkpCrlATcNc8NUgw
4mxLWrlzoiVeaHntbFPrtCZJIGykqpVW6l57ZZ75ErnFoK8dVfLuCwuEAnzpHm21ejaJToGQtPeW
8+Ufh7c2AmPFm31bR71CzG9t0T6+TksoogErHqlw1yBjzQrA0tZbLL2eXMl0L7TPOFBV5tvqj8FH
am51rfH3m2Fj8A+FHM3Bzcampr87ockwnWvOVp3AHEO1ROYYpreJZtoCefTaPwIgfz9zFskSxjg5
N4w+IrQs/VG/DpAUsvHsh6tiFkiNsHDecsbfnqcrqsNOE3ODKd2TE8MeRrLUeT9TTYRc6usNCi4M
U5d42tljug1J5V3emA9ylzRYiMgifHtBBReijWXR5f2r50xi0d1lnLw//bti0imqgo1cngwqEyaX
Mr6PIZfbl1WYyBCretscx1Uao7ClSx5NLFCskdddQ1okk0zEKF2n0qK6AMqKAcso7F8tGGW0NIPt
i90GDOL03Ii+9Y58z+WKxPRuE+lSm7Ul+ricrQacFMv7sKF5eIROjnX3e+Ajm+tiByCGLXKzfp5C
ig+oJwg16nPuR3knO7iaYALpQcEAqZ6VYbZne0gatp46qIqohopUOTbT+cZ06KVHvUHL8Rc8fZmQ
HuCtE/uOGOxWawAl8ubbDvOmLllWIdJxoLjyh5Png9webGrBdmPyDP4NPO6w6gss/ZmScA4Rv/20
Ao0bx6mEZtr40PLors4AmfHtHCops5opwnCtoj9ByTF3trs8svDyyX3maUz4xRnR5QfeLhYNxW0X
agswgHxIa5iEpmD9qj1ean/u5/LWTzaOhi4bqfM9m32HAJFrb6U5cYSmxZHj5r/hVVrgex8yxBEp
VftftGyKxEjjxxjZg4IIRFgJEypdI+LRmiSqbMf5Y0kSrecL2fXaQf1jN73Zt482S+1Vh0pSDyUe
nFBtIYF8ydTclRLROA28jJbyaJbemtI2VshdGEwGHz7rKojlccB33Nx9LCaaIo3cffReODpoDBrY
sprbsWIHqy1AiIAM1asv9GSNneosqHW7hG3GwmCdnR8UUDaANIXNvY2JSydlLb01j9XgdCiPfqjj
HClErfSq1e/sxp2gD4GYH1IthIP3+SIa/6TsI9xIxP+W/nesd3esCzYkFJxh+j+JXcvDqaNv4UEa
tJUj6eepMcjAxE5RhRZH/P9TmXhesQhFu6vCZSUna041c7rJfkk+zZAAJzaMWo4dau/Fxyrp8GoP
mTDOEEpw8Ff1V7p0YtiyT0Qttum7YDdu1S3A5ssCv5bfLdZd5VXuAUI5NuADgDh1AOtNfkz1ODdt
l0FMvoWuUnIPd5exzurT0iZD7ZXM73oHDu648euB7drjBIl4DtvhSV5JOJ+oUsiwdOBTRN5RvPIM
wTbuGFz618WSMWZdnCjAwsEN7od7frXzUbEkCuo8tsfejd7TLtAd6cgFHdfQn7F8cKoN410nmvcO
IdgvuYxmEnN40QDUSrFPnH7w5+cole853h4NeBuyJgWXhfszDo58kCS79/UAsG+wsPlHEIb7o29A
EpotQ4WxLepXYI1LAjT7QU7v3SVSGKYjDFULzQZDB6+cq3Lr7Ca2aLDpLrg9bJjpfJ39s8aT3rsa
H/P2z8UEQGK/2IoKu4pb7as5oC89XeKiWs96PoMtzjl6rMTjvLvthT7gZhG81S6FsByYwW4yqe/c
tYI2Q4PSTYGEk/YHIeA9jnLjPY/sh6kbYE+B36DJbwzcmoM4wpUKpvK3Lv8kDjq0iaw2sMSHYl3b
PQP86Lwzkt8/XN1hcmaK+KV0ecNlRYb1ptCELSymHtl/djOmZsY4qQ5XEfJgbyz0rSTbxyUeNJPK
lX6+MetuWH50NwqzomAWkMGsclKsg2U0tUzKRd+2DxWThC3Lns0jHRnzpf1liHgy4FGGhzdQhlTo
e9BaS3MTxmOhdRzR+ThpEUDdfI6BIi6orqI8cjIwy0TuAAXgzTfXor6A64uJUzOcrU4O2rd3wDA7
O4R+Oz27gEVwW10b8YEI3U2QFLQD9R3CTmahzJHTZmSNpa9SOJ5T1sTkToeYA6k3uXYkGtaBIXhV
HU5IY+HIs8rNjTAXd8/wonj3hHGnbwmsvqWXJtY70JJNc9V2mZx/lanDjLWy4vmS6HpuYBgpamHY
pOJDwczRdFuKU7DZIKtY997A7OIyZwaU8mTuvBu66o35gpQlbg4P0Qu+AsqJDhQXC1avIlvC6eO6
Xan5+salEGYJ6kZsF7clJp4oOiZmAX/X1Zh9dllfokx/ol1ZmgfCGdUiYXRC15XGctAr9l/ljCi5
e9hARpA2sy/gZfFbXX4Hu3mN7jfGM61GpG3l/nhMq8lI6MJ+N57herVatChETLMC91XTV3d19iD9
IQ6hgPP2OYJwQcLi96Wk45lsbiu7rnt2H/UyHchRtXRiOHJgPKsY6kdPjoDmqWXncswizQwXN725
TBEKtdhcq7uFgZIoV5cJMqUP3RnOZy4VYf6n9p+V//g71KO9xGMRRoV7o2TfcMi8CGhmcze9g1uy
nA2cnrPE08o6Lhg44faMxNh1Ly6i/WbapeaeuxaxCgFVBfZgdWJ8nz5qCgJFEXIXXHh38W6V85Jg
dSqtqRxdl4OrV4A35aIkWJOn47LtyzeNVFtoTD5HzX5k5SC10TUdKtcISoWskG7IEOWMjbhQbNvH
+vxrClo/1ywkxHzXFUDhFWIpm+pirBSpAx+Q3/noBNJB8FIdvBYU/02/7YSSoMT7Le6GYWq+JECl
wJEn1Qvd+h/sffKNBie1gfpoEl2bMAkBn88R6J/3HOoimtgaYiFQqQ4BWVZT2UxqHClIhpitz2H0
GteCgueilOmzNduv/1Xf4n/lQeevFYL7dNRdBYfN0aistmQkg2Vw3e6q7vykN/YYBLFZc7Uqr4ld
WjW+ailxERhcCVTlZGncuHofrq3310S+pXjAnzVskeROyCwP9e4GukRlqxn7dWDJLxsEkB8UKkDP
HPRHPj5NXTFhRgGy1WSWeQikDSKGwJRElP59tnniNAgJHHkO+17li/cW1zi4UnE8LMYPnbj1q6YE
9vagiiJ9bgKgdAVFDO7D8lPW7rjqr3sLXKK4HgYaSBtr9pssDIZ39p+yJN5qznEaYmwz9JES5XL6
OOD7qTIfPQ6oRMaLVGccQOu4EKbFSLTHEmyhTBJmbU55e5TQS7FnmKLsRA7t7X3aW6biVEPxKcUH
BvF7aziayNH5WdJDgA7hpb8HI8O6TK+/5x8FXdZ1xQKAh/FeinV/PGYklQiIlxML241SA04pb77X
pZ5sf6Xis4wKcXa61GTUnTQmkff6Wf9egSCguN9kCBkyuF0PSnlQfoY0Z8EFkfSWES6damx3gDYG
Yfznqver2/Z6tg2OTjhJR3LwY+oOOiM9fEvo9/pwwaEjJQnFjvTONwQGuc94Eargj7Gtf0HmJxOG
cXSkrLG/X21CFJ5L5SBdGKiMKJ8+MZjLE+lLywYz2G0aHI+1n4s50TjxKCn/jUPe/lXqelrx62bG
eILa8qxpQ+y5EicMUxZf1qWzsLwIRfD4WSxAmRKdCoxX0JKrWrAUO1Xgdmrimbd/bAF8TUKWd75Z
YcvsTcKAhXyMUobQgtJRQmaHFiq+LUjHnABqxok0AeJFh5djGmo6kGGN8WhfXOTFYdkbg7t4G1Ds
xR1O3al9ys2E8+JOe3jXEn+QRsZOmgyvhkjAjmTViBDBToclN+eLeBp29oeRRQlj0hNWPoqixsKr
+ebTdqFdZXzEJPw0DpZ0EsiO3X/Zwu3XMT3aamy4XpjWGflSww5K0HZYamsxTDvieg1o0NikIoZP
SNEw3X4JjVkWH4nYlSQconVf274Oo0YqPJkk12G6e9vFw29VXT8/6B4b1XyQkc8QjYoCY2CM1a+Q
/Co7djxUfEQmz9mwm8aeIjQ+VyTaNfQ2WwPYIKE8Q4lwu2PSlCiRbqy86T86L4lbpBqY73Kd1alL
vt6z1wwa35w51sL4Ronf0hUIFGS/YUrki891CVVKYxx6imX3vpFVjzHjQCJdUfW+ilrRJhX81SoI
aeeiSoiHqC6iM/51NaOSIdpqlPrsS1BnlBoEIZgSyuVkn5v8anmZnvup/RyxQiVgPZ14/RU720Jx
7iJ1kyYobMAn02SFSMMK1SyB2lZ5VuYuWeoK/9nIV3qhbABXiZMRvbq7b+wKFhI0lwOsi9nR91VO
uQKTtwSx5Q1SsTMbXvpV+cuaDcCr4umu6h0QoQyIjkdd0hiGRu1/p9SaGerOH/TBF2dtUAWrGTRX
zoQ9xgyGAgS/2w51VcOzW2xzkuQLfp1O7loAio/guTcAbAipR4Ntio1AaQeH2Fl63UvJex1/9bvT
pgZIbkHQ1UcOiHZnvt0yTXM+KtRKygQRCtfOG7TUMMX328Jm3m3XSxotTFb+iJkBwVoKCnA0GUHm
Kt2CRFmcx8AgJfAtxTEhaBGO5Q7IaGy8eFupJ1Mavo7IKmLIGhUt8V/GBIWTmd4Qj8LHvSF7VjWa
F8UkPZRc5TgNPYbygJeksDHRwShfETr/ram8akiQ9FaAXgMSkE+RBCcCAyd1hrhrInmrcVw2mL5U
o3hAkvnd6kTewmO8Ii3cKuL56ZOSRchb0GWMX+d+9XKvunoTOR1ws7xB2SZsAqeij+fRiMQarPwA
aviQJpaeBcQKXrnBvtHhiSpTGawXSTKIu7+mU8ro7CNqG/a1T9+op0aKwQaVrxxlgb7qlswlJWEy
LIOHOAV4Qw+USCDGFPosjws/2b4gAB5QYUZ1I7PUP1e6NHu74A6moT+MN/r6nl5Ay2QPw3s801r1
MHUp91mnEYftfkSrh3vJCyNri0Sx+ZrjyvTk3rurRbJAvhe9zb/h77miTf7qlydkVUV+TG7ACSA6
O6wC58r1iT1PnWyiQS3St8qDEoNhBKKKuzOfyhazyMDsBBp/2zi4rd2fKtwhEPsxI3b0N7/lkvjb
qxCty1t4AQXxtLp8RNWg7nwToFn/AtUDkx2fZVRkF/VZ5mD6E9denm5VODn6X7sTLUHoL8wSgwok
fKHs78Iwrwp4GUjR1rt9wlPEFuLRW+ahdnC8ZRZneYTE2eM8ae+B4FXLul0r72sM1zZFTZiDSr1q
HCYKExRulF38JPrnyEdvveZoREKY1NgEcDk+NqfL+fnF3FfYzCOadQZ25qKjkhIaHsDTEQuCSnKu
nsBrNrZnicMxKTDyRIIjDN/WUUsUZlJE2vlufFXYrMiQgxrrIMWapjbbdUJOSLy9Pir5eJWrc2Oq
joeKuez1Iun4Xo/t9s/TVu3aO2m1yHvF4h0KNLuZpSyZLQDhdnTG6ZVcoc0Cv7k3jyHeVatf5ZR7
mcEUnL9Qta5mRM3VqzwNxyo71x64e2IfsftZD76h6dJS/mMWcNPgIVGqu6wBLvCi7ZDcxlJ6e5rk
QiN5zgJhfTg+iT2e00s2XJMZVWcYkG1YKv4Ouxt6TWnwCetkF/uV3jl67tzYMBuUy/zcawVkF2J3
nFVErqjX4snVir3DEZW+iWiqIgeOgTQ0yeousawdKfwRuoouWHyBW57+MWPqdfiam9WIfDAoxjq/
XQo0WRhI/kIy/bXc9pOTDTRfA4W5xb/v6vsmdxOyYduqf+7hShWy0mpgBVZAD0uwqn7WD16F371u
preWVUtY3fNHlXx28v10qnfQ/3PlLCpLSaipXf3ZQDMpAgOk85R8lJpiW6RnocYiHGBQJUPkAprI
Uy9FoqGmSwICGdHvG4ngbfttVMz89DicOUdaFOpWa7QbSzHUmKXB84FVhgHw5uZtLT6fVYcco2w9
8jY3ffLMw2rViOtdrEpzFDTXkLtQpG7cEzml6PWsBYy7h12aA7a0A5z6IXPoBGh8ztfWPloDSJj5
WgkJjUVH/F8lJ6hUIrhhO5DneQZgXEqdfEPGYt9bgb5CKQmMzN8hRNUbwfRKdjYiTEooI5XvIfzi
Po3YPHshf/tHZA1zy811O3O4VYCNFiTp+WLn233CLGOkKC/fvWiW7KwAMBE8m5Mlt6kqqVej07wX
gkXl4Miilvd2JMw+QUXa/ok3BONvHbiL5yrZo4gMI/jKftSVi8GgWzavLOJ4zho6hmlfpZZxIS78
34Wh3ttrf1vYF6S8OacegsMEZoQqY8YIE0DucXzKFenBbgRVTGrZ9MDdLfIFtI3DQrlO3EwmyNF1
fEZRhq3HIFGETAJgXAtCRiGTJceIJ/JJMMDnoGYuAG+DKeV3Ze4SoQqPzm0QPNCzG/REuuSksx/x
xhUwgFW/5nNyhzzCL/uNMrlrAy7JPhzTJcLW21OT7DL6LHNKGfMx8LpfCd8+O92YlKat74tLXY9j
CcRZ0ocDgB2IGGdRoEbtNEuiH1qdAX9CHbiuoTnwC423VdiM5yyF/FkeWB5mc2q4psYg5AVqo7hz
/GaU9u7AaIaoejgmS7Q4p1HQOGxoZpCxTOQb6zU9fZ1aRB6FHChzajzZM20AJIiXvcskxi15Bx+T
vImoJuKdITeEU3xQ/ZOrTQNjK0Eyg1+jElgVc+MovKVyYftTrNZ2AwgWvnNf8TRTPMI+69M6O0kq
zi4tIHpGrn5bPetoZMBXr53+Ylgyw7kHXz6Vg0SIOQIL1kI/iQVCGBNO/5ZAvfzbENwIL+9l0m4N
NVIjNuULSQZXG2VwHsL8RVzLIALuvkZ+/YXh6OzeO1YH6L6bmu0icctqjEHMoYvAcC4efzNMGueV
/2AxbgDlalEqtgupDvVTGaUWbAf+fB2PL06VHAm76aFzTcrXj1nSAqN4UtiY0U4Nymq0LZ0VKpAC
7mXR1c+vtqqSxqnv6UlE7T5CBSU+7mkMRkTDhgz0Z9RcOo1P7JDO4VhuxeTV+pTA63X3shRWUYK8
kfy/acAbru4+0AdGlaMeT1xb47u3zhZGuwvsB74aFBdup/YAI5vpmDOuFQGtxesSVGqu05onrfAY
FIoKJmJXyahUFJffCzuzEeg1n3jecA0kYmwcZbYu4r7gPMQn9n9m95xsvFZOg9kfHhG/JZfZGs1a
Cvudcx1eRvaAv9j+jWc154TfPMyCq3YMCHM03d6RHofAOaPryIqotuYFpfNb3yX4kHeHAdVnf/hg
eFD5XBtqLgftruHNXtP7VUL7I3sAFjBWEGS3pca4jbnQR8e5W5P3WbduMKzZ5uRyk5WmsEcllTtu
ugh1ipUriuDV6ot9cYSiiwAvWngky0uX6U2qQFE2evi/okTlQyyXGR1j6HFcQPGbwusyTOZHRBh/
PNDq/OmY8V+CgMrlj/bxgjAnvfBHvLRA6bQ1aS1Pkgru3liDM29w0agUOYuWRWPirUNrQLPDXt9E
ysUsy8yfaVrezw4rvVRJ3IZ62Bbt+R8gXKUEAdj0xKkevSHcoFwcPHZc6jW5o4Q1NMYpNkRq0YO/
vYt/0HCOn+VRXRhrpmg+Ud+cCQDOmI2tlgOYe3BdsCaOtxLdqT9YjYgeuBXfk47ShdYEWUgRywBj
LsP+CS+PngJwPOx1OnepY9jdge+H8PYpUluiVUd9fNb5cuNSaBn6D651FBH+yJLBmyeNCc1KBRgr
xZcMuIJ118ILFXSNhCpzL+oK0+jbvPSB+GyZTva5Nsi6aCq4KXUYEFUP72xhXt6Sn4eKPKYSUuN7
/MbDw5qi/vW8HR2PohLma0oS3R8pJmoaz9YoSjEzcQ1wx0rwPHTf1CkP+iY7GnMbOQ69Y0nZykFf
uX5MbTbCZPOX+7jc5xV9fxkNaucckEwCN9kWN4Lb3iThmN8EQLoU4xF80vgK0OVWGrlU1rX9wl7Q
g0HC1DYPrggvlOq73JUZR6aTMtWIXarNhexopGsFE90LQZIwKRxBnZbukYrD/po/+S7nyTYhTfZV
DDUt/vudU5FlEg1DZ7DpPhd8eG1gkbTL/1yB32ABIptlPR3IAbf5FInMehCEQw021oKKBXMiE7FS
3GnkLk5erCrR+k3AMYXXcMyEh2m3V6LNNi7eSVDwhgzm2zSl57VE5mwcIJNOTACwNh/IHAzkzi1x
vwLvwWbcMk6TlFE8F+Z1l3l9CUqyTnT9bkWXigVzlztmGk8ARyC/eGfTb/fpjh/9h7bceFU/eQgY
sQd1B7fABgvttjn6WJS6dRRwf35b2xm9+dRUd5qQLGxUI+gr77xnIzgpu6ITZkACrGkSr04vGQaI
w/dFpEyvcvf+5M/g6JCr4KoMkiT/1umQzOvS430WlMeK3R1Hrxw6IJhoqDUGh6aIAfpWSwi3wQql
BKR351+JDbSgRjGhKXWNd8ALtEnRRz6iN8r1h91J8ZVFNwhUAR1WRG42Zpcs/vo+IgR4Jn7zQ9jU
OPihLpk+4KrTeSTJBtKuujfqtOIo6OPX/XkY/dtrdcw+gCGsviMSXzYziTykV4EQbmwnTxeJRY/S
gv/5YGRiKql7wXfcQ8HyuW/NcIARmyfeJdmF6IUPvuM/hyMvseDdNphfzLJb1IAekrCKOZPu478f
5CSQT5xXEpZUsgy9uRUHu9LSQ6BdW2n5gzMEY8dJ9AWiFjwxwqNLLXwfU63RcuxDWJUN40Fgdt4U
XdRG4Okq2iu5D49R1/BKo9ZJkLY+Yiissup4M4WExwIi0zfQHlqIp4SrOn/x+f3dKTp3/M3S7dWg
o/tosl6zJKmnIjC3R+BnkMPL62T/lCXtCjMqFPLjJ9r7sAK7tss9HHVxJZ0YfRJFH19JKPnjJeJb
lwRQrm4xDDzVt4KZUP/oz0025TajLK9Fzx3DOu5CMM6aSEzUsPIz2f4/AOLlv3UmQhjFon5yshaS
qmSCuBhw/VjWgGFGim536AlZ52uxtqiVIan9FlVq4JUIs0U5dc/lxIrHerET9Z2lP5cwyHGqP4FE
nw2TE5dDoc4SSmGrMRVDiqVB41UZOGPxSmj7WlobsW0qFzSNaP5smj4JRZ9Grn/M8tQUEdgBQYri
vKoKNr1DmMyRtGQLsMe9joMAN9sAsk6/N9XiCWBFtXT1eFrsCttUVndT0deojUaHcJ8ECIAkcxqm
ZlSBa6QgO3MhK2oNZMHKlYKOa0vZUHATEHOOTdndp+pzjmIbJwtHZ9F/r/BgheRwMdtK/gmzTXot
SMx86bzNlYCprDsDoxwfDIx4U+tFgm/L6iI60nRl/IC+RIkOJcRY3o8axfWRlrN2hnr0Emn6+UOo
vJfm6KFZ0uFq1xLsM3v6X5oSZlmwk8p4+EBO/Bo/w0WiwGhsURALh2OljVcQzV0CKmox2Gwd3Plx
CPUEsFrsj1RqTAl1zsLgBhiXOQoSvFYGzsUZy/1Fms8IFXFOvKoLTrOPfnp3a6bT/AXSD0KnZ6Ja
/kG6OeKpWQhM++zHneJ9NpHHjSM2kcxOookG7RPTUP4QlcUvbEtkktlhSby3Wure9ZwSRDjTLJUI
NlQCjKdqnRvDVsdCsTOE6yV418pVNfhSMAiDI02WWEi2jCOvxJpaidi/C/Cs+NDs8fczb1Rhskl2
gDJ+av/PlJVGpzUAirsrD1+tVOJR+AXXhG/OCn1QAuXwUX39SXNUpHM7XAV0WjYtNKMhExjovxxF
ZVZyh/IDSCsLxSAyAVhPVMGHDKb9og1/alvleRg6HLGKhaZBe9wZ6zvXlICNYnkRkECaIr0mGw4I
Dnbf3gXxz873QIiEmoltEHVf5a/XODU5R8B2ZPZju51R0STl5MPVi4zXyRJUk/X1kIyLYtFVCr8K
b0JL+UE68Mats2Sn38Uf1OImkWxNtf0FD6BXLdPso/Lkmff8wWoW5KTjBTJ4XO45MuxcGoigwjz3
6eVQerh9GgXWNmmzgscdfxOwX7hA+U4ClPcOC760yvzIf6QGnreGOAVmwDPJ3oHWP0TkloOBWIWo
0tuQq3LuOHNR5NAjRKOq2ncFkcEzCclZkkfFCuuRNNPfKbJDAzvTWJYM6frMNaDMUbiP7virTFL5
+43CDSKqzwDCO/U5N2jXT/KhxQPN+ArgpGSIlVK8Z54xc0C2qA2OYknyKZx2ej/8nVHvFRoCKSbN
jg4Dtrg1NQ7IrmFQFYCcbvfm6TBWCcxH8KpTOokEdnmFH7vVBcex3uttWetmUe5eMQTePfmnzLHE
q8Lx/gPH9chje7O10gVrxKNsG8JS6GPiTof3MLknAYuX8MvoBod6+g4LsITwvZEWjprBj665Soc3
hN5XjxFCzQkv/eI37v1oXvALxckMBCijIzLZfS5Fz/VxIq5dy5brGnjhcFDhNJFYTivbtb1cvP0F
MvYZpNpFtngIb2hcaXbXCIxLsBiFMFAgV9DB5aSuv+Gi28p6z5AqB7bvqQmcQGpg87L2GkLWfx/m
a2Iooy9InszQFWRmVod92qjY4wwAXhxND3WgqVso4ilsm+9SAl1U1OYxH/lJoa5/njlE2cIvgqBg
PsqxgpZyIi2uCGuKNDD/UjvQF6RC/QBjt+9SrEji9bvRaOTelWxkIo2X8F15N6uSLO5IYxjLqa90
h6O6q+hBsLVFwye0r7mVHwv7NKxPPgS0b31HYvnrj5pp/flZxsW5x1j8s1RBTy/1TQ4Yk+6jBodu
WChJgSmnp2UQuSRkfB91myPkuyD9mKWbv9h9uWaE8D+8Vbm6nJ36A8D8u7zWJC/2hq30qh36NpdG
i7G9MkDS5TIdVtEVTlV3Onto6Jx4mf59i3VjlvD+LCsrGSMoqi8xoPosTBffATmkWzzKYoAaZdoZ
WbcuVrdHABQ8m0UMZN7iI9cHjib12sy9v+0TpG67Q/shAbRPSoIT5OmWhOgaXIyxC8kViKV1UR6/
kR5h+UqYEtthX+wh71uWd8udyqAy/ZEkG0b7LmIBzecTYHjNNs895aO3e/XLIyaEhBBL6lT2CJrh
l0c3lMa3NMz0j0cp+wmnC0iXJ7/xYUdCP+czI1+iWW2ICZvDqB+J/5d4EOWVzAvolEP1Zw5aOTcM
y2BXSwYxOHuHAYpOyp/KWKJbBeNBFspq9FMVxrxXr8RYapUGN+5o1PmxzLYqL/P+0x1vbx1TjpN9
ClK6Nr+curCfI0pE/4k/9N0CcEoQuJZQQ97nawzKZTg8JpcYAxTJ9QQb66j/vik4GJw2j4p24Cko
+a3vg+bP24F1Vt9o+11+799kpqV39XEUzY7TUaspJyeMqUqQ854vW8bcOwZf1ACcUl5N2YrPgP5J
xH8rEVE+pJ3QZtpzdKJCvSjQShfF9b4mtaL+1hFxRFbFeGGZ0D+yHeiXtRF9liZ2Sp0qD4mEIzC+
BqUW5Ld2GDai5VIgnriJmHsy2ML06DUChoJqCDjGRMuv+UKVkyxm3QOtqyqYBsCCd8MCN/qvQspk
k8dggH++wvSgKz0RRwv1PtjuEKQwkVI+OKK2YLpoMQf2zUvlNB/V8/gkcIF1XQ0Yl3hXHz5WNxmn
XGAF0Lu2TCFqslnLRPbWOzDqS+axsyghNkKlB9EfMDUyJRk4P5GgggwEWnj2Qm9I9PNHe8XWOjBy
cblG/2fQM5v4u0e1S1G4/HZyLLKJISSMT3YRRCD4YSXD7nYt3FDat9zFe3uq1MqKXOMsq1YX7Cqo
UvtUbL/eQ8+vPVPHvLTlbWM/BWpZQWiiv3EYZolhTBTZdCVOLx4XI8UwFyrq+5kCc8yvuE5+mcCW
Pi/2ZOFtSHwb3Hb3dIOoR58MUroKS9g6FAZxXIiA1zeQnkI7SFvmt+q+6KGthXAdNVFF67XP/xnR
18N+fngIq1x9LwwVzY+WSAizyI8P8AEruaGQyT9B+ej41bwF9h7j7bfYuZ9CKYe0wUbzJbQZC7+A
E+XgfGfWlffV6bwlDD9Y0YPXnAQ0r+/y9R9VBNcJbA6YYAalBPGpgQ6h/f1/Unzy1RBZ/QwSd2/n
WhND9tQQa0aReYQpnNB8K9zRo7nGwX8V75ACC1LMhbHYgbAehZJE5AsyL388pf+Ij/fWGqAXSb1K
7XY3/dpjkOMX+rJo+QzY+sGhHADFYXbUMlPTeyfezYENVpkJCol+1cPwx8DKippIBZLRfZMmRl0g
zYCl4TxZy7chAh95l/DoykhZhAFkenU8AEnqeL/45r7xzj0BQghqEO7BNRDNvSz7R9OmLG+eGNie
K3Hf5obPepw/ugikdrf7+vbD5j6o+vOh95LMJ4msqNHsKWpkjlxdqezjvOTotSOOl4gb/epxhLV9
7meM1NPir8bYMJeJN/wtbdzPSxTAj2gU+CeomaQqDwIWtwU/RTtHwii1x0cm/Iuvzmk8jbXGEY3X
fEaA6BbZ2HUZsB5Uma3OoD0om6iPlq/kO+hfUeVnciCRvIAe8Ee5K5t2F8cbVlJo/gfycTH7kckb
nVmJ9z1EFHkbIuK6JHd5fR1ac4Qr1I8wCTqcMl/GpFX37pECxmff3khZsZzC5CZQmeIUcG/kvrc/
sN6hqdcEG3Ri3Z2JotbOo7spgwleLjef5YlkO+eVsfKEcrMvtKBu/LYfhF8N6uid4FfGQu5WJ+Le
q7F/WF7ChsXcD78kz6oaF2X+42poC5xfcgT39LHcaR+/4D77pmqNz0Kwbz90+UMSzVb0wgZQ+jFi
JrMFTpPN/6BtqXATlS1Okgsgl1CS12I7k3j2DKZcEsQq4PdKNNWva+/6B0joA6wDSOZJ4RQqC+Qj
GmqsTPbARmXEhgmfU6+D6gGjylhuBpiMwqJqjnP/rgiBVJ54cJ9zcVTk4hFlusd1rT00XV9Dhkrk
ZMFOGvZyr8IjN9G7dcaDAVTqu7Sc0GJH8/ctlbqbFdNns9s3eT0RBBbhHQzf8dEON35x8FmPX+qO
mxZIDDkY61d/C3HdCGlSWaHzJSC4DWRtT9YufgqbHcyKetm1Kh9ToiZ6/99JneDa5udq6yZhQWuX
zereeeYSekjvg03Vb0UPIu98Gp/8itrT07eW8WY0cKDVJ2hjKQp553vEqsE3jH/iJ57iulvB8nGK
M/zsKAxbp+puTJ6YUW/xn7NHPpPUC18RAd7ZEOhvE3Cfi10Xo3f/vFU3CU5tDaxqTGfSjgBSmPMH
ral8ACEWQk3wQqDCopux1F7udK2LYEIoO9CaA2uhp92WYW8dh6cp2hJIOoDxe1/CM5jqbocgOTok
er2iJc5ShB+HotrSR5lJi8qSL8wW1tTZyyLxQ+JlUD4JcJ5XcccAZ0qIIbZBHKf//2PSMUVG/1yI
40YtBYgscEayxSVGv9be9JZZIFeOT5G7MbT5aLmS9dQBc4b4zB4fq31aef9caSx/0HNGPxFSKohF
Yn+hTpL3GmgNDet9tJNHBO3/RlLd5TYphOMa9oc1wsdDD65VCjqDiDrTfFZ3JltLcwRYlE3/NgxI
mEPHTQ/BW/qD8T2cdFZWUuKVk3D/4Zzyq35BRaitfG8ki+Y4k/nIuYflRmq7SwIOumaSV16Y7H+t
EEp/CUeOI1sXJNasgClKwbEwPmiYY3Nyg2L9/635Cqbu9mtJR6G/7P8gEeNFfOUkhC+7W/xiu+xr
HRnIzysRFSsW7f+ZI7FbOvpRjBoe/O3ciL8ful2xFmfB61IPkPOIeQcGwbv17CbJ2WKHiUHRu1yp
jBP1Y+YF1b2/Ch3rg+FBW+QJ9E6M0RJzv8OGlht0Amrrx5iA3v0d+lY7Y0FEDx/Wgem9w4JzAz1w
qyLq0QqUgDGzMduOwadQlEbMLNveU4+vHYzuO8k9QDevFCgQNZpdlpoOydQk6gHOO+vWhFTdcp23
H7biOi0bGiwYwxPbP8NNPHiMbV+2IUivJv5nLZ9Yh5u/uflgZziDdL5SxxeeCI93vSJeNgVRCg1v
Zjw8yJGGm3rWuFQRwMjUHZ/uBQHFCOXXX/d4/HUz8avTR31Wnx7wKXajszmIpirUFuWM2fLUGVOX
y1tl3YlxqR8qqZU1nawe90LORLB84gQocdJTVUqwNk4rhpaUZGpyE4H/fjr1GTLxMx2KY7SYp0zJ
xhdTLPBb4s/FSgUOvL4NUvAAuN45DBQDHHAO1Ggv8lByg3hAhnk423XY4A11KFInXYzeFM4+UfNo
VdFEwMaof1nFz7vfvzH3KB/33yKY34fNfGYQRJzSuaR99G1gzvJ9wO3EVucp+jyoxTn4uNPF7Iz1
UYEifPaz/xVH1AifK+6O+KMB9/7M3sndRr9lF/UxdQbt2Irn/Uz3i/6V+KA19FAyLKswp/49HV5a
dc28VS0TmBDw8UWNqcxlQshcZB4mDsPd4n3eRRZHpmccnNdSMj5M2FaThiPB57FqbT/AO+yc7uJo
UeXbrH5O/nQOw4uuVorG9QVAOhFhdpKFnjlgBolUFmV8wh3fDkL6FfV7eL4JIBWB+NFON2q9FNGb
plPVO/lparD+TK7Py9VDmUanfMoIRCDP0PqOvO2HXyjmP93Aoi06qte6pFI7zz/FW6hhc3XZbBVH
q1ZLaSHtVp8BiZg2TXY0VZq5tV5MjImq7RaamvTr3FnSWcqjuBGOjGf4nG+CZfwKK1nu5fcX1+mj
LZDRPnHHM/K/KO88b8T0D1Rnu+iEnq65V8NP8jckt43BhJxr0v9uV+r+uJGiwDIJHVj7kvzgjZde
z7wrURs1vERplBn9dguVK2n1aY1nef/xEzQc6WiXrFTaZQ402gCKOKBu2BK/WKTrqxVVm7En1+Ph
I3bt8ril8WnKJ1I0MeHx/Bkn4CcnGBe5o6Ob6XyS1lz9GJ5bfO4WdmdlUdA9YPnFHQ8wdGmIf/nw
5HuGFdQn1ISSrf008At6mxJkAFlNjJYfJ6pai3x3EBO4+sm+5fdFa14x4WrO/OqEiQ3Tug37VNl2
0W8FKoC92F8wDS9IH8ziiBCl04BmS9i4vmGXiavbo8x5H98A7nhFZqgyK0cA5EQX6Dh2M/nTrfsy
NVVcpdUtfc8eJnwau6J614L/0ZT4c9su8iy3w769DlHaiWhrRSQcrXrMxBqm5kBJJUitiJuwtAsx
m87KaYTRdLRdKrSWTU0cH5mkrZvBDHtvHKqww5rrQE0oLcmK8ZI1BlYwFlRKh/+YFCUQlHUvISdq
tgF11RId6eYL7CZLObIajOkXf3VbaGwJSs0FY3aRXad8droWG9xYnyL9EeRZdC1+/HJroXXYb487
DeRxkHlZfXyuON0xcR/M5w2vippHLVdJnX7jpFpYPf4G2pPBBF9VkIR4orhCDFPKEQZlFuE52upf
oVR4JMZSx673U05B3qtX14YaQyNk51zS/BOGhV7QNtsa4Q/8uca9rNfr6EmQjuwNKhMcE53do5WL
mfKKStl8OrI6+RWeIEgaPpEOsjpKvqwWlqi/w4GNMllRFv1z4aWwyBRzbOl1LnocnWnyQwrBhH3Y
FVFSS1qu4uHeqm4s91YTSoLM9d/Yw9hJAb8BnNuMiJiL/A+pTPcMhnB206dEWHKLywq0xHAr04yt
O5zI1sKgXa9+GXuxVQPfO/aeFPLGyryjEdrOgsCpyq5UttxbyYijYAOsWKe5SuKYIGv4KHMl3+ec
DcDxbl0dcKSqxZfdT4WfNTQxBQ0Dl3EtZ+RFi8zz32OhWaSQRny16ubb8rb0kA224Fzu+Pd+QgEJ
h5dXmU3zqH1NkE2LjZ9kYXU2LEhAdlBC4cmXcavEjtfz2YjD/2mYzNEEEU0hoBRvf21tPHu0Q+Ha
FNmB6KLN1Ecqgi0Aja86Ha4MV9Nuhrnj1J5TwTWb4E4M0oQhV8f1tzfu7r6GqHlBIrUzTGL23HPH
FD4Zz0NrrhyH1wTFDU/MjqJtW0PKFtxEoViyJBe/Lr4zSrA5Akfi5D6WLW1EAEwIYxAYuWJYiFUG
f0mxwJzj6L0mxKw2aam/2+m0dg8LYKPG4UZeoZKq8/4qVufdNvEV/Hs6XeXRzYE6Dim3M7WaSTAO
NMhhId39OxVk8DM8u5S8OKQcVTczfHlMligAB4p0usTG0vZ9kYPwYcsQ34griAMsj/p9ro6co8Zd
qcwneWByLxdl+mFEPgQMwHw9SBLMqZ7rN2tfjIvNOQ/qb1114M9T7eNdL52TWDlqiFKoQM3fYzyI
TO66PrKeTz/rUurDXl+Uu0WmwH35pMyYV7Ro0qRRp2FngjSjt3Pl3Qx/qSVWp9iOHw4Clw1gZpm3
2pc+3NnxzAX9vqO9tEEFIBhErp31+RWqA1IlkdqERyz5QLWMfahAq558HwrgGwthsQ7uwLKfg2Jf
/NlvhAsKDvs6WsNTJMLgyJig/A6PlaffXdCmJBITlfaS54BGxGYTvTRimpVy/YFHFggPKGF/ub+w
mY3YVccSqT3boARcYTdmawBWmdm9/Wzwroqzzug1kKZNRf3iehnU8/j4YaIaPYzsYZdj18cYgmXL
VOP9BvUJk9dNskqT7uqT2oHYAJdI+GPo/gDbUbXmzpJd0hw3I220JzSUd5B2lXTZD6SyGz4xawLZ
ohqilpNvAf807KYAq3NMBqAo+dW4UaAkHzGyqJZ3f2C6b6oTk5800WbHVIPL8qZQOMshsA+GLT6n
L6bdDrbfSVqe1DuZIp7WvxtVHdAhPxSKu4Z/Zg5QLM1ClkGicq0/SLhMZNdV24WYOvkyeUEp5LL5
fKNNwC5ObJQ8Yz06X9/CNjZshrkBjzBkVadwsDt1g1RxgAnzEMFjFzeHOTwwtRJUAre4EuI3jd1t
7QSmvNK/wrvGrDE7au8U8qn1J/k7fD/B4eHwg7HFFuRRuTa9HBMQMlg6UNOvX9yJY63FuDLdt9ZM
5WRQTvR04SrMtTVlKdaF0md2wBgpAHuJ1LDDPSq/jMDidjp7m4bwRIMCv4udLSLTmyV9lEXaiSFA
0PmfLrW4FlHWCyOEKkb433zgbxUJrF/CPShE6u5r52zfy+KtoJ+R0VhJVVGqrYfFfPrdPd4PK8S2
rtT34WXotxRjNFmvmLWjjoBwC/IEtMZRCVvUW38pcKjaTviZtG4QJd4UxUv+9GRI91lRMNJ8aokm
MgiAtm7V19FzDHrduIcdN+GncrGgUQDRSlsYnpeCUuBJuSGdGMf8Htcrszkkp5ksuVCZK3mG2RNF
gGMyD9wQpwdrRmjWOZVHUvsfvc4k5BttpX/TTXDP3ljykCUCLyZIQKP+lWSviJuYacvmQte0MzWQ
hVNzuNnNTzYKBzdnRr7kJPIeO+wUZNiF4XS3GdJnYunaa+ZE5xOBa7gg+bXnoDtM4iDNCoQE2lZM
bBudu8Z6ZafR2Mrf5KnDMtTpHIv54u+V5cksQ2BBb1Fvnn+pG4Wm5xPZLIBvYN93xWXTNlmXdcXk
j7jgEDK4AJOli/S9yNwqPLtNzew/tkgJ/1vcnTAp+8hM6EFpIlBdKoCOO22ujjRmVrD9ZEsFGF9B
h6EMyJB63eL4Ojuw7wQntmbzqDOiojQfK0Uav2zTTu98b1usIRxVawblXlzyp8fda2vEf63WVmWI
xXY0WfWwGJvZG0Y7QZWapEV6DYDSt0Y1an3saWzcRjV/ZBOw/yuK2WCt6SCBQo8AElhjEg8n/ok7
XYdCYeIe5YYQhoEgcqV0c5fw5nOEyLHorMP5H9Z5x0ct836P9FXf/EZipXnEojC6JLle8WKq63Ik
h9W+tHoZhkEAv+/g7u4SPXmNFwh8GGkTY9n+uPCTXu2O1fFx/vXjF730MRdyXAS5c6rbEuHqiVJU
tiRrjw990DlXrFPkzcyrFv4MALYX2WDqjgQy2Hp+NfrCtWOTPEMxwY4B4ZlDonz4ThqzFlreIbnI
HjzqlyCszE6aAhazeJlFGrUQOlkWtS8fvoWp1XDnzJZ+7BrgOnq9lV6IMkYPcl2xfC0VwYNn01Ef
9/H8AC4BCt/GnsQZ0rxzmYyrO6K/gNf6vGuUpSP1SVNs4TkDf0ScpBaZupQ5ChBMKIviTa7DtWnw
DWtvcYGyBhXZu5SFP077keSsM8UAypyVwgQX5qJMFTtANknev+wtNisM5tedEDXydiNSnwZ6VClb
cDtbrORP9dZvz2+B+NaAjzsYws0NU72gwEuSicpP2QM+Y+JAPkAy9z42p6nKycJNzWIFFb7DocI2
46LEZ0yipiBB9T4T+QW8maclq7i0/QWAGIzJRogGeyD4I2rwYZuwft1bqPfGnS+2zB/sNmlrDTNi
J0pc/ePRwSfgoMwx5mByfaqeefPqs3yoZvtCaVP4VZ6X5bkQ+IYku2+4lDc0WtfdGx4oq+AMX1ZK
T0LOV0QvhUnUxu5gRunZHDp+DEhixEfZEA1cUbIAPwOpLlNDA8o5Sz/r3pE41vAKUtNIRQLLsr5t
+hV3edJDv+9lEd3GcJkNc+60JlpQaTPu9OWaHQZpMlcD6PBflV2/m3T7IlYs97oU3cbX7s246NcK
KUlIBe1JMNTR50HlZLw16jGRtFJhmvfCi+WFjbBtk21v8fmUpgVeBZgXupDPgiG8Am/vS4Yj3SVZ
Ose5JJbrhYGRdYpjEPW7mPNk1P6ludXypNBgjmFnal6dr5dvW8yGhWDqct4dLALDlhHgWNkCeuJ4
ZItqjM8odvPdLdndEJmgXDWhyF+/Y+8dAlK54SbG4eWZFN9HCNUFyxII5x8MIx2yR68FyOg+2CWa
xPX2RRmMMBPLWuDdwl+c+B2yCARB5m7el5SGLyYFrbZFvn9HJyf4sad4LlE+E5I1tNnM4i0c8oce
2uLLK9cmJtKKRgGe/Q53Z/PyT9+7s5gG71GwqG6SOrypynwILYW1h+puq4BPOn6QkzmnmmEfn5G/
SJ6tWqfvcvvs4aCykYAexQGIUdrF9UoJ/d6mitI62mh6LwOz5/QMXcnpzRY7F1+a7UjopwT0PN3X
1nwXzknPf3e7xPkNm0kwmK7j588Ei2rt9jPBO391zo2u4iLtf1c+4C7YIeqEnzZrotCM4fy7cSAF
j2EbyQqUQEcYjmrVgR23ASpqPieMJWfwV1cWc+MMGD4+qn66ci3JpG+wOe7SdBXw/Kjn/H5f0M4T
lDBcLB3mPB07WH+UMb2OEGqShXsL2oe6pF5WhN+WkR1MdXgAAx0Cms9yK9bbMjqpNo3PO7d86mH4
aGLrQTLDXQwZdQsfn6X19cefRh5nbUq2IzudhbSqBohD99VoHjv0011QmDe8VPds/IoD7iuGlubi
q5qMaMtbUSNT9mYPFiOAn33jzpfMt/WKhWOhJrJoqP3zWBPF5OpQUxzk2vn6UrRvsjux9ksFmVad
ByUMavWiL95nHWr/fnzMqSdnw8xp38BrD5O92yIiyisjghvedl89DtWNsZ4qcKWodle8Nkkv3hPv
Zv2tPnxbFZ2JhWEXbednPKx1oNz1Jb/mFAaDsEeIjmsULKngi/ZnTfdlh1Z9rD1DJMqnCvO3zPcs
Q8bnn8QlM1Vcy7Ybwukr/RZigk470ZrMBkqUuqem96D2VxFwFagUy7bxqdSRBbU2nnCC6s28obh0
s998eJwHpNZZ+EQa/fVeapRdwCUIdg9mzMhmjjCPSOo09id8LVL5curMiQnf/flUR/wS+wbW4PkX
9g7F5MdH7sVRBKYIdRgCsVF0cguH4Um+ovvGd7juyuytXf97nmv5AA8My8PzEwsU2b4D249IytbZ
uz2pSppA7nEIxyVDGo3RYRMLcrff5NM9EqPLLmC2Ub8oce9RnRqrmlHYafFq6OgeS8bByT8VnAFq
j9bvnCIulVfWZGbF6a+utOJxdcYFTpmL9L8LMdqGD5Ag0Ge3OOYC8hdBXm8DgL62p/eQ/sE1CgXy
C3+CGxXkfrc4kCpOBv6JDMS3onfzC+3oQrR9jBaxC5lsbcmCe/JVm3PsZUDrHV291R//ITlo+UgB
10XBu1+az1qa7HXpXWyW6SMtx1lzmd/56+7+pjhTnA2BwCA37z8jsz0NAvA88iJI/Ki2Scd8nYJz
jd3/nP1S7x/rUDfQywjwNutAhNpx20GUDEHzveKevly5fYH5SdxfhsyT8xJL8dkHviTBmEWA5LCR
ijX9z5ak8RCGzDpV9EFymQ9w5b8pXz8jkshcBox4O1djs5DXmIoJl06HE/GWTfaSYmHpXA0qIcdE
zj5xyq7lCAX+y6ad8WorMtRvaB6diahSxqsBr9s0wzGxe1mbCEi0FOscXShD6Q/nHcdFCBaMvIVx
hcMKMyWI3g4ieV8VkLfruPcsehDBxH9iKNFH1PN0wvqKfPqNQvHcub91KbIOCwTsaEv1Jsk2f26J
iu4cR/teA1JSyvbXMeLDu0UEnwtWCxg+jP+cer1m7gb2YYJmO0Rl8H5nMu6J36NlF3t8SCmObOq5
Gr3OH8ndW6rVzCvnq3/kl9IILb7CM93gg23KEX4Rl1F16oy7pRA9wx10YP/KKnxLDLjq0gqacEJa
294jjFco29rK1AbRdp3kOxJbft2wCvhpQJNRLj+3NTIyfoYCq/Ok2EENeG9puVlsfcV+qXtAExLc
EpjHb5Bu0jWYo4hodKJnH0cPRg/05Tvvk4kVCQu7TaykZ8VUW/MkKB7rUMGCd4dujYdFZPlEphzx
FSSKnYqhOIbfT5TpGAGbd1pjZgRZi2xQTHVWi0qwwgLSc0lJYVC3x/OuMzze8SPbYjCN2/X4XtKM
s6uBSbqimKG5XOdBqSMizoFO/ECsywAqBDK9Hvf/oyo/lV+ewqgaolgHbmprm7X976VY0au+ZW2t
cZokRq000foONDhAv7MlhGPY97ILz0A3FxYAfPCOXju1XNGYsU5X0zPaqv7TEe3Lcqm7wowOYNcq
9rsQIIv/c2iq+mR1TdKyut4uR74qA3CcKX7tQEgw2juGyyDkII7DeWk9Pv8rQToK9Y7DtNytIslO
KI5cjXkOtv6KlPxMZsnFH0M+U/dImahWZ9zT6rlCgclZwKY0BKZDSzH3agS3ic/7TgLqrcqIaxT9
Eu/D2t4zAmbWK6ztTS/5wzllq1pxwX4CZTKyXMqFBlIcFDwkzWoSOnfKHNk6YWrtSY9tYJyNJnRd
/SbY+2s6ED/YxVzV7lUJIwvS4iyaVpK+bqg5vDOWUyARnlQEmoLogacx9EvpbsQ5wCmetvBxuAoo
MTbOq2KCoX/OJT8Djugw0E79dfeJnFYSffRA0TkBJc+kHspeL7FMo1nHPdcXthB3QdTvjOrUQTKj
1kXfqvywiu7k76X/3zkjaPXyBrmcoJktq1W7JfQKKFCLeg80pKclqe4mr4v0jKjjIkHaLv5imuZp
abYdHWhiyvUOF6cDsBYTNS9laca/r5byJTnm/n67oJFQdpBTLIJYUzb2ozxamGN2tHtcnptQAHnb
JHh7uFTpjGBt/fN01Y0DwuOkJ3azpHQhUpf4r3tiKVc4RTfXbXLUp3ay/7cFbiguOjF8VNnj8aPo
OMbbEGFuJDMP3mzI0mqzOL0g3IYLON02M1KRKEoU0vY/q1McHtv0t1O3SUpshEDD0bU/9onEQFPL
m9OyGq5+WsKzXVN40U8K9OJiksBu5cO0UM775rv2dEc+c1lY10+EaWrteAY6sCtBqCzMXBMJLIiQ
kbSgrXzAp6OdW2pZz3p6dAkzUerK5lgDB5fMsNOlr4hJknZzW3xwzQ0yXQtdEVtvYsIL16qM9g4U
cTI6k7cGk5ORdo54o2Nrv3i30+1gyh1Iss9xUlbYFBO0aa0dz6go64XuKFSir87BC2I1fQTun5qD
uywgBBB/z7WHVnbm18RKgWFsWAEmecBmkh8CoZCWPljQTcVcB3mssh68nWsWwwHPIlDpf/KKbcBL
BkKmcCl5l8ClzCxqR5Gry0vMYOh/6YvzXUheuX8UC9cNZBbebCkB31wwBXS4n6suVgVEfgwcp7DU
1EWnhZFopbyh3+x7GXgp2wzDkVyinVSkjIy37LBMnRUb8/EFys3eLwQwLQgT5FBMadkl4IOqVOs/
1eTgOUtDnltqjZfZyKwAwmX3pm+ODkAP+JlJYzvjPdQLztGdGnJ1BU6/XSzU51eS9cvZRvvBop8/
li7EfycX3S/lk9WphgET0rkQXBcGW6FtoBMsFd3CK3i69kvHWvsLhbqqm0I6zDyzxrJuUkO4xL/+
1ghdfibAgCWgd70iOh7Ch4Uko4oPYe5UhgHRCNcxJ/inmnUYlJLJM+sv3FZwRKo4PwhDWrAXCE6Z
P+V7ejX5fERX6qcwUA/9z3BrFeQ7Q4wGQJM8S7MqWKgljsvyn/9UlVNkioSZYgSmIi0nFJnegkqh
HZsmyGsIzTHvyYec0limZwEiI7U6Q0nrtSCfOeSNXjdGO9R0qarTmjVkMbnt+DjzVIxNXYex9V9m
k6xVx7wpwdsz18rXbexGRtPr5rkS+3ZFnECi6fcwku3h8Z72HOQNiTBA3/XGkQv/2yYGCdpdNgib
Ar7KHefLU6EoViT8h7U1/F/XqWWmKNPJhomKjXzZbexKNFajVgpHyAEeSyaX2psOuSQUpvRmJvBJ
UTtDcFZdkfhamTorIbR3fL/vpDCivJO4P3tc69/HnYDnI7xarThwdo+BRhuRcS6Dyy0goIm+rxX+
CsUElzIMhmIXB7p3/yrODu6NNiuJEunxSEW1A99h8dPoel+Y2FXOJpk5k3OnnAN+6Jf4DBlYyHzO
zT/T9goOemNPXxfwpKZX5FvNEKIH/J6yAv80O7tkT2yTDYttVM7lIIORcQaF4H0gLlRHBwbvOGsH
lMRY2RQdXaOj4e/JQreDzxaXWYHo8HnXVuQOFP2IUJNUmaitg11ERCR34nxMAA4L8VG95xk9xX9y
9kqVGN6V1oBTVa0+HSI7ZTRTCVwXv8VWQU65AoPAKdZjCW2vBYbnet0ZzV3qgPxGeonZPgbnnMMI
dnKUM5ckZ2EY/n1e7MhdVCb9qUaA1imDxlXAIYM8mr47WX14f4FzhUJAdoq8rnTqyx3XZEgQbz+N
KK4YnPz/lGVDmHE6hK07JpAPkPanqPdXDvmm3HM5UwblrNHn1sXRT/XUlqt2IGz243LNJR8ROlmK
pw8rQyiOLnWmvY1pmPJ3qoP23+erK/Hl7RqeegkiBLfyscduHKiZ98Hw6sHScbDA2fTe2ligEmWM
ATz9o3hO0yBUMtOxIMCxOteJKYijk+BtuikKTJnlmcd2FujE8wMOq6netR8AxdWMuWhPzMyaeO0M
B7y3Zh2vb4HI/JckvsLe9Wlsy8ESvI5hvAzNZSuKuIadvhZPyLYVU1edC3si5JphwdeJy5KkxsO1
V6yPq1bjUALKLYTwSkxUwQ+8n3kDsN/RNHHBNVdpICfzv+/j33n18+ZjAWGK9yZAphEZtc1Iy0ku
63BtjwB1AGRHVURLLImN5ceA1jiJsud7VgzuSXOQs/k4uRI0ZkNN9evBPlYooiylzaY/S52UJJJB
VuhguE9oRXcYGZUiysVKH2a/VYF4gB22BGG/FCIcasz4l4LtnVbQP65radjxqw1dmSTIAMJdk2GG
FI9oXeTjWoJpPMSiRP0p+dKQCQX3nX8Wt/J38KO8W/5ObysaEsNSGy6S35d21KKDImq8emG31qD+
uAoL1uu2V7c25A+e6DNSRy+CXZdLXqfpjLZyeoodGNFikCPvRH7JJS29j4Fj6FQuS9zZY61WZvy4
49Lb1AJ1Wt+KS8pWvZoyIrEoWg/4n5iu6G+uo3vkBiAdzVcRbfsPThx87fdkBN3qoTfp/oLSR0lG
QYkYMoeG2qfiDn8NEUHEW31HrDSyAZFR+9raSLoTbJL6ds7GcDQDYeRkiv7NaM2UtFsWY/WYbND5
g7GDKH3bOb6sVHyQwph3sOSzXyM/tlawhRdE3L7lliToo+lTyasZUprWB62SnVHWYzQLwhJj6GYW
C4JP/XbBHKqRzhmb3aiNy7lZFpeCBtlZrLyASgZ2VonMFNOG2Zs7/BELSfgC5Ccjag27JjNeGXW0
9FB2bczbnOQ+4LQdM2flg+UthtFrhG5H30ibNymBDQ78sLLDBeiRGHyaej6iNXnKQoESM9/2sitn
qAw5H7WaW2lIakJw4rbz0rzDCSZVGMIcmE3CRY49LYdQWdEqHrig9pMibP4BtrhVWnova8sKVT5q
NdW/HarAKR1uasMHVWZFZpSuyyA4ZKDfWJgb3R4ChSFIBXWUwaHef/Pr+KMLL2HDyYos9EdhqTyy
UUuYXjRHobFhR52otlWo5IZienv9/LiqNZMkyK0gKLWPGcvPzmae2iCB/7gJ4j+LNg6Fb7Ab7Ixw
jiCeJ/dU+BIgEAvwTCm3W1F2S+OIWFaQTKM9wn5oevOXtotJ4C8SM90dNoArVbYWxzydAP8O5v3y
HcpRYuORg4IHCIYKos6V7B7yHuGkzRw4pjz/ZkT1nUNib9SieO3ocmPF/vCx8NVBkB2m19vvxeIW
BYRw95Un19iMwuWM+yfhXfgNzbwHkjYCq3Czax1iyUJXTG2VLuHuPrpR1hXcCUWg58dle2LJ7Sjp
k193GUKLxIenBSH1UrMqOdAea/FtgJcwFsiQzqtDcBqtuKjzoJ3JoI8fd82ArlyQQSjfEcyqnmBQ
F7FjFPHeOZt6GBAiC5dqSyKlyhpFAxpsD0vKDW1DLw1AmXpOHnR9KiqtTgjpSZcigWitPe4o3mDe
vdn5f4Xk3bda0L/9blM5pn7/Sy3Wp4LmuXabx9JhbbxIEmfHHvT9wtEPhQIXOBxiCZGaohk+W1qU
AaSAQ1RfC8xJvojWk+u9PolaaBHrxGrQh6TTJZmssgU2xi+0vTRfVxf6JE7bkHhS75RcEA9+a4Qc
q23uNeOTrNd4lU3QQeNScE51e9i70igM9Zs7YhKOWKigg5+YJoL7/46G5rmEroAJ1DaP1Oe5AT/n
gu1DLnTs0Fzuk9Iu1OQ/jldF9n6vt9BDwFt7ZCmXyN7rn0Wh/3025iLBp+yS0njcPCaMF35c3yfc
PLZc1XXGz2uc+Oi6hNHQm5yo49j0Q4EMB35T99j2w/Ps+y+l1aspYhOyJVJ/ceVPnDzz825Iugi5
+Go3uxjb8LFiCERKAe6fwHo+At1Y7+w7WfCB/2Uf32agTGlf6iQuRKJkfda2/bMP8UMCgXC0tR9L
5No3J9XKSNxSaAz5KK5owCsvUey52N53YUSIum+Yl+lfQGjS85VCBHJ6vh2+UHxGLH7xylQVN7yu
tnZNek8Z0MAkoyZh/G4HSZtsftFV1XHBoC0DB+mLj4/7k1OI40gmeiCPrmHDCxr7NjCigsvZN12h
lXwWoZUUEoLGoqcwX143T1oXZ2Iv2ktxxqr+LKWS+TdUgJPsljCq162yIx7yDnUnzz8Z8JIOJrar
j7k8o2Wt9xo179BK2rIkhCgS8KghxwTtPtmvR7z+pMkypZnvWpOmKvBGcxMq91RQSGWLww9ceZSD
XK/ipBP/eRig7svIGGNW8d8PZpautPdkcAE+BUgSIMyposzv708ilOA38AWRfzpLomrlaBPRQqiW
/0S2xhyCHFwFyaYs/6fFSznBONKQXm87NwKTUquiTmG9YrOkftqhpMO6DK+5Jf1KXNMdcv7Ec5WH
lvVC27rc62OKd9QqJ6mq4ItuWhkbg63N1apqOsRd49FACsHAJrkQL7TfCXUMc2xrvaD51DI59a2O
B7O30ZUFTD5RnLE/mEBor7q4EqMUvy6RiSMVh68xu2oAnVO+6JbHxTFLcOh9DBUOClm9ho2N9n9R
IGtczNtOAzQ1d95BDEDuSSVEgqaSZPAZe4idFeY9REIfJFKQrpDEpr5EkvEPO/LfKMVYpa6I4cjM
POizDAJfw3oeo43HjWcHl0Yp5H+8Nkk7PKizcIoXxTXkOwEOFgsj+zForQl/YifFxKjt55uapkFq
rXm/8dV83Z1wxbBz7eEXlJl1UTody8fgVBggXjAh6MlC4Gvo+AapyTCzUBCvSH9XQQHDiVhvB+Ei
PKQ4Lclyn/E/TshPCMVVkPJlleuBdeh5XkTuh5NCMP1YomxiflCW37L7wUHutanC1Sxad+ZQZX8x
ptkDkARfyoOSJwZIMAsggcNDTuW9FSrFl5FgaRe8HV9o7eDUIywyiY84+kDNr2O1dHZ/PjAvknWJ
oR11RMw9eFrAZo2EWAC3Frngcxdoy5iR0h3QLOrWTzAMOy5YxhDAO5Jgem0Df+VmcDxKPuNuMvoA
xbUCu5ytiAbOYp0VODvH7nGrn/XmCij9b9V6HJS1Yuhy00ZLg4VUis5puVG4dCoEsFBsT242NsJB
dLdywvM1oS6/sW0L8MHM5GPqj3MewMKSvFAMVnZOuFogIP/+h36Ym9mxhSTYjawnPwCRssRnpdkN
N4vKGrq3wbUEmxrD83sBHQ==
`protect end_protected

