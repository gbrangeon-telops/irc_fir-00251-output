

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
nnA1LvIFtXuhnEgnrDveU5DQhO4oCdS4/TzHWVjuSWRiJTWamPLe1zKRcIJ3OgsD949QJsbaygaN
jpuk7BYNZQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Cfy8I58fHjYLB4BFaw/VxzidETwabyuF6c2nxAde+hbLnyzOfkymKdOr4Pk5oDTY4htTgTDRWzMe
dytGdfmZXjp6SJIGysindi/Logxabu2rWzFmbsNC3Q0gro5se9+3qoriCL3M82gnhvX/joJNLiXg
rsFmmSylhS6v32W24xg=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Gu3bZVKL/oo3WMbeK5OSi9dLiGmyQy2yONRw6Nst9yei3DenlP6wnhfHYdkStFXi/uvWUBEeZ7hN
0Bmqlib8vQ0eJP09mki40prhGAwrKuqYt+2JunlvLYMjlmKGJOXPgQJfoYTNzbZDTWMAPlUaZkK1
oZkHNa3Wtk5m49sk7N6rE0lY6V2L8UfgTL/MmCwu7DKHNfTBd2W2KricGJ6ICGb/eh21T7mo+KTw
su5JPh2xN6VOnDqK2JFdz2Fe2UsNNdpq35qIZsc5dRna+xfhp64zhbzGUq3oNeTCYYFL7/rkWyjk
xMfq+Y7aGpW1qrNdKLCLUa3C0oRubzA+yEUHPg==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
CjIoJO7bPG0vgefcLg3HndCtGBfDCnGBCSVZItM/kv6K6ZpvJnvEpEF/v7GEKszxgiutC8bTrPRk
/jMI//klbN/ln/AMlW7lDqpJ5wXp83c77tloVq04bnPwc3DaApr08oK3Bf1H6JgBuFfaRFUfxoRB
6anIIq6YC6xrV65+910=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
D/ZhWxzQ+2vaiYn3/fV/u9o/WEb/ogG/V9KccsPCOCWeaD6JXzbX1wTvk2mHL3gwIIjopxpeK8ct
Dd/kho1WYC462ZEZ1ijvlrdcQ6jRucbVeVK20vWFMC1CO9YW54zFCdUIFDYoBjMQnJ6IU90guAMg
K2P3LVnqKNh7XA5585Xm34QBVEtkbFVGa/nBjX2k27AaOcjv8CeFc7ihUp4B6D6YzM34GhHkOxNj
NyMvVJlZ5HBA7JHakPw8PSgdpMIr12xEOrEcLpR4AR6H6hPW9blh2XXVPneGey+XXrhV6WAB7P2G
TGbniILS+ojY57htkmkMwgWfAakIRm5HfiYkdw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4720)
`protect data_block
H5MNJmP/TWas7XN3GhF0KN5LGypA5CWmLReKpZZ+aLxaIGpUOk3ZFpsnkWotzbaxBCXx1o2aUFE1
WVKw+NIOueXFsCnTumA1gtPoxMEaWb9vwgPhMc/Oe6E2WNjSV+5/kVnl1BhiGAeoqOw3hZGJMrxi
TNnPc0cV7xI7JPaGP5OhG8NXWIDGdjIEJxvnR8VQJaAKD6z/9nDdz4GeYDeH98ZsO+OCyrleYCF7
GFAIvmziHGUfj4aGqRS4y3d4xse2ftmOa97y/p2E1rAjqpGZeli/6cOjJb8y4efXvrls6UK6Qftb
P1ebtptfGKb41rbHEmikXVMcar/nE+jLVaGNo0JDleX3IfeyLifW8qQf1oBV48npxaimAU5ZLAAX
ICHA0QbPOGj/NyBnCmxasZRsS/JVAsrzaFQk0PT+ITh2kJ/xGDp3tqKcyQM9n/WHmFTEzIWCxrpk
NuI21FysjVLrHOJNCv3GnDASnNCuIaIQsmWn3Xjr2HVjP2wvZlqn+jpWI36qRlrWaGXyET8o6Jv1
dfzBWChxrWgNjPpHE0+sEtflzf+Qhcyy16P6oYVeS8s3mqsfZoJROSfUWXM/AQE76xGctOM3+hQI
NohbrU6FIRaEUDhyGU6LoKVCPnvwuVY0eivmjPnHRap3mL7z7jjcEBk46l8cddQ9GuyoJe56Oot8
+c2L9mtO5XsPUR2+22SpRPfr/ZS66Vmja4XQNl69WQ2r7bkPE3EcuQwta9oPZEuK+tQCtvFQc/QI
h551+WR45y7ZtNFs1ofuTYqSg77qp3comfIj4teE9DH4jAePiHTs5cudbQgsR57dj2jlJWO2Dunx
WTwuP7utCztDZVGdLZekVRfAkj7bAIWez7CjqSlfSoGDUCNobgnBmdVvFJSBTzw/kBd/aBFANdQM
xIzY3ABaPnd1MvWMeOK+kzKUsldpEMXZmA06rNjt0wQXDY6l53TJqdUKwJG2ijBAm0VD7cHSysyj
CONo72tn3M4TJcJ8FnGqRx40iRyB2lxJ2VoP1rUBjokpVvOfW4V9CzCCaKb7Rommz0sQRr5P/xlN
rIx68NBoJby4NVZQI7Q28AjIGXC5LgtGolJa/FAThhzgb2GOLv7/ZeugUjdPy7KVA7DNEzo7lTZg
3QUP2QUC0KbwhgzU0LJR2Rggh4KXqm/KK2LrK4FqMa/VmFqx5XcgDP1/gA7M5Q2HAmUp4yyPmiAr
dkqRNyu6tS7KgVpcXKtSVjrVvyPM09zbDAQJKvWeUNUKRUdMJbQcnFNeGC55lH/I02ipyzulDR6D
uQVv8qgszkQSCzpKTneLb/YBGidYFZft0xvg0KIcnA80CBmM1gyQ3VCXXrWRFso7+lhR5NS0d0TV
oVosl9cT2MNImNDbtb82S8EI+o8/a09JS5cs/dp4u/cdDcWZ0iFoa7ESV4UU3yi2jnrDTdBrzbhR
BV0cwSje+IeXOtnmQv1sYkRgR3K1VW/K9vyuDftc+kP1yPb4ayCSV9lW5xMsEB28doRiOtrXASjf
qSYYvUj0+REZ1bXqkhrgpNGSd0Nk+qvBboZEpdjPE6nH7XvlRS9vRuI/fxTfKGlixlxZYqm+GXhK
dewB0jvoPB4bk6RCwMKDmtJs0rDUgGFQFM909fjUNZtfFJVnUyT6gn+MkSfFpOUgCazuSv9zxtmD
UJ+B0iFWtLWQxV8uLtJeFcX6p+N8z1P3LweJijnkxZSSZzuLbz0PpVc+kU/dwe4G/vLvsNSmTlG9
OnnXf0KjY0Vd/7G5vEKhe4Zg7MGaFUVtSJjGQVhGpMH6DKdcUgoSo4BvW9365r023xA162PwWeks
jc4fH0xcY6OQqG9OxGdFssPTnNC1MYix04uO4rBdJfcs5bwy4mBgY7ZN43aitxVFTplFT861V4bu
SkCqHacZMpdZP50t70ngydlDI9MPp0swrkLHzSIxHzNEmfYnpXd3FYJ2As9Soh+9zdxubUcikijD
ZznaReV8Fmxpnc3ia4m8wJ63ScaKTMnF1V6n0WDiAfekTWjyEuNo22O/nT82rk6xXsAvd4pNRD8O
BomVUt4cytGIURIIfCsYLJ0DMaFuVBo1wT8qw//Sd7KFllrOptjJBNU2hYOZ5c8ibGrF520dkb7C
Lex7ZaCJHfvqeu1wYzoivUeEmCAVawFR0kGrXgpiCV9vgnshDMSJEyHaYCKmPsPHJLqjy6D5pgcc
/Z9z6mcS37cGW71IOUb3hQueSZdgOOiZAKO3I5KKX+755LyBcjTTnnmwUHJjtOPDYRJ1l8NVZXzb
vgLU56yMtCz2YfzR3CpFacuU7pp58XdubMtnkJH0hudw/AJF8vEV+8IKMXCWVUylkC2QRrYbM7il
w12wRrxbCZ1lUVcB6hVSoy8cEWGu0+D/6s7WLs+mJAbHvr1EiQzCiEZeqEulx+/Bvf31Xjj5kAa1
zneBw2IVaqBw+6SinLs3fFaFa9WxwdloMKLSKBi63DEgdaAkE0+E/XLnxcc1W5vDCFdY/3PBbng0
jDu4jo6U5PomzHAAHwyYVss82QiqoWXVDLP4p1Y+sEBjczj6EzRCQUi+HxI+6Q5Ide+N1X/Hlzis
FnLza0weDItzKDj1klBD+Gh34ZKv4NYHHctUDrx8XAHozmy1Qn8HXYrBkxpnnonwoSka2hOPcKJS
OADMVRXHLnducYmqCV517BE5UxIU1JNSYUidbwIAn7fpYplhT8eDwBb4VJ1LBdds4Yqd21IOmJRD
kFsANH4iXr0Hlh4lxEZXUw8oYP0LHfUCs75mhOs2ODwoMaeSpp/e8HxYOC3UctrTXnMrt12Yv9Kn
NPwK4lZagKT1hlyEpNPwz8yRgRNgLKeH7GGcLrtJ5WeBuRrOvsx3W+VAVAhfytkAP9WeyZFP9FSK
Xs3QP250XyJY55m5Ci4DPjB3x+ORxv8AFLdYXiDpxN0bWLJfO9utU0KvNILaDJ9mHVoifeDat8j3
ys7BUQnoOBFaayEHIYGtqxzxYn14lL1QHIvwVhRedEed6DKaVczU6pel+79GAUUuf++xsovHWnXp
tzTO1e1VU1TLsf84raw147gjPBMjlZaV6Mi5zPlbcZK3CoDsY0aNBTzYHTmyhX/ktq4kU2FlaXjk
2HNZuDqBO3eET6z4a9FILQzXMiwyLBecFKrb7LA70/7yNebfl9msSXsT7Uue0ZC1v7nZPcKykrR5
tLpup+lgO2JoO6mPxaEXvDrg2uCnHspBWmJlbLamN1OO4Hab+KexcuOFgpnj5XR6/0hlngwraq/k
cfbzaip4ZtV/FF3iU5cnahi8HOWNDr6AjCfCVdYnXBnfxyvCWkVQzto7hHVIrTqJ74Pz7E1uL2Q+
5Mo8rsSafYl1ZgfUtVk3mzrpwCXukUxbH16ERGoG+/BVd2BqpG5TWklT04g3JhiSeIOl4qYKXK7K
ZCcktdfxE8pG5xT88WjnGnMe6aSZiOcbgndsPkj33wJ2K3x53W9tTTCuvIYqqc2pFP8SmFUfcYkB
B4gu7Zyg/hmhllPipnfmIpN/wvgM+o1CehvzaZUK8tMFPZ9guSPK25ar7T698FmfNh6Ov08qGZ43
FEgL9531Bz+szRzA5mP3iLer6mwyVAy7kGdGAR1eP3WQdDTfkQbk1r6yE0O0DosnPBRDNJhFMH2S
bnGgib8D45Ik9iWt9aXkch5b8DPjcRS9XJmpXt6HqAx+cCohdc0L8LoAI0u48DAsEr2QqYH0bMR+
bELj83xr5FAxHqAMdO6L35S28FG6A6yKipqwYv6m633g0hsknmRgE/BZ5vOZqQu2EEezpCa5uDfp
jwattyTtrrUNtAb/FJDuAvS9P01dEeM4cgV76N09bMitM//4FQuQf99sXG6nuiQ9xxsVghNMLMw0
h/evXssuLrxrBXOP7LjrTGjZYKzowPxP/tkaIJg0uKdEJPauhJ6lAHWdRmrdh8Cuhxos/wcLJsIl
d2vWVeriw8vze+OjsmjPJJMROx0psgu60N5cq2VdDPT7qQtimd/Mza84KvNZZ8RVhbFjZ56ybHu0
DqpgH+SlJITgUdk5PNna82WAOxIThS5tHz1siY8Z1e3qNCnahfuSneIdqoUhcZqe4AtqTUSVgOUz
Xy6vDqCev0OqbhafjYdB9Qwh1wL1CBmYWZ8qLj6jxmewVgETncaQ+CD3WEK+ADAGj0bDW9t/GCDI
AzAZXIEynLX+skNkG/EUhu4o9c6nKWF54reE6ZiqQ/zc9CrTiHYBXx04LbfWeN9+ELun1ItwmSf9
vCdfn2Y5HM3WDosyULO/HiylOIumwtKD9cPQHFcYiJ+l1qcL9mxFEkVWCJ5NDlIDVC5caaK8A03G
qeGIwC30aaSA17uai793yPESNozSOdkApD+JQ6qjeuY1FEYUcRbMjbV45ydwga3W28VDylvgWjL4
edorrz7+UCN0bWg+qgEcxAt8WBIgAiXGtJUgouCcbOkNIq1L35phWLt4jUWH/9XnMR1m0GC6adiX
Jho8PCYtwD1z42ogv32VIwt6eNJQUgXZb60Yqj22EMM64Z4SbtqGZ5LdGqJ+dwyvK2MIiRifAQAL
8tgST7I+SwJ45/9nm5sc28X8hlVubngP7sTJr0qnnrKiyW5QjFEahWoqS89/rpejJ4i5cb2OL7Vb
jgVApIMtRcJuwtbcBQd6lKP4R0hv6TaDaNxe7/emF8ztRi/mApbggDK1pCGEXYtdzxFSvuUbjaN3
eDBY6+3Tw/ohGxicCRicOC3IId+UP6M+eSHv9fya06RYzYH3CT+p3pGkg9hmtbGdeENecjvOaF6y
hqFbV18K9X2NHpEyMkScySYfrSjLFX+Rq80W6D7f1Fq9pcl+2Em/rTY9A4gSqUsTufNrI4nDF9EJ
c9Vtp1uTwUwR+pNdlVk4iV3WTM6PwRqQ3PwXi8W9otrtAJ/d1lln3BK9onhjsosw2CjAw8U5v7cI
lCrjbxbja9GEZV2tuR4tgfIhV9dBHcd2pok89rsly4ddA4AHqmQYilT6rANNVl9M7JzTDzJpK/5J
2UIerp9zDFF0fX1ggsCuqCcq6/lyEVt65Fr5r6s7p+7zhlEUHLa+WLSvhrV/h4o6HfNENL2w6UAZ
KIvHFEN9YdX8EmK0w2n753J00fCxKav2ZVM7kdOlXJOlRCqFGofTg3WoSbW61IRv7jHut9tX5Q3h
bydl4xwgBYObyLhf1KG+SYggKfYdsY1Pq9v41eoN9JgCCqYpph+ohZ56vDQZH9Bx0rvZIEb73ceY
OxgyDPofO0GFGTJ5nnpfl7bEkoHn0gDZkst90cyFxH61fKDGOhBZLNsUntZ19cIe4L5F5e0n/J45
UsIIVO7Fti81aLp05MuQTWepULxHUhLMyTdM8n/v7MTK9nz80PLybsCtuiEnS68Qocjht6iuzRT3
5ubf68Qhfrvbf0IPANPMWcD63uwEut7k20ofoaHWeKet6mYPZAxCC6LHfOqYVc+Zcjd3zBq4n+f0
vN1igGtYlPGNkMSt08cU1GNX3/ricqVZ+Tiq7LfU9VaOJJ2/jbTJBd5s5C032/P3XnbZ/HXPz1XC
66D3v3MksiKhF7lF2NGhY1BQXHCDi7oOGaEneMZv3V5ZcvIuXUS3HXCozVbO2GhwJL5QTSER/R+y
/Osf1oMQDM9eE9TrjFyo1a9dQeuLEAMXPWDRTa7vb0Bh02+zU8ONGryFatMjy8JPF9YPXhe/RVy6
JbHMUS2rOpqIQBuVsMX3KNKWjmF137wiR3zoKkq/4TaaD3dYO6v0MlwTcZI6aURhFoHd3a8wgLxY
y4DfolBGbmRNdG5LkyrORPMMrkKdLEhtIXUJYfMIgmDWncnOQ8TayJVb9pzasQeUUdoEeYeTGMuj
XvCy6dSqsotFp93Hgw8b0OOVCohFJ2UyIeeis9ZTMv7ttgfRp2IXJqliKwI+ozA/KRN2/ePsaiTH
hcU1qlSXcQpMfVZHmrFEEE8SACGalQJ9SE5qd7s+PXePPwItyW69MfpSVPsYpwV3ghIpp/zi8I+T
si+R7seXipnSxIae6e3YXgSZjIkz2CvkbPh7jlPRDuq/Rmb3Uk2qVTqov4/8aWgvx0ZHloD3b8Pn
yiN8nmNenBzNzFYO8Qtg26izJcPyqH8J1YKY4j5k9Z1ovK6ljqKHSp8BGhh7YjQms4mt6P9KxioN
gCTIdOvFer4PfDrreQPL2/IkrdCNIRT25EKFJVXTUUlh+HdxNxEltcXt5zscbKfuLWYah1Luoxlg
Sj8+FbLe3Kh54wOjj1UjHlv5KNjn5aTFVIXkgBeqpRNNlEfF6a8EGEC1UYsSfw==
`protect end_protected

