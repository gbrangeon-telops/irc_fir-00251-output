

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
CZom0vHERP+sM9B2H0IfoDUsJRy9riNTVWFr3BZpkrcd8N+2GrPBLGYjWv5bwWNFs2qiaRKQWIBH
5SL3Ros2Jw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
RCliXKg9Iz0QVLqI8b9GfxxBU1GhNUODWipyNqGvNd7T9Syer0VoYCIXvffp6DiDgM+PWpXEJgNC
ZPrITDndrkqwjZ0UurJqd8Mlj+O4jokuol/hbGtnMKDg7LMTP/mcm9YRpJxuqv5WE2ZWUtD1WAlU
7OzpzsPnbliZhM0CcXY=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Kq4rQuO4iRu44woH6WSrRyNcsAgSUJbnevjDngvc9cypuoYRq4je1NTd7KtIptAfdlUTFMhOQTcF
fyvMO0ctzr5YXTPO+6ZCPBMymjnbHRykXwGANIGORUKHiAy8zVrLHGA2Tn1n2komEaNoM+u8Q25L
d17PGNi2LYc1A9ZX79yuNo063Qy3QX5dSU2poXOWXHho+u/vL1PlOKA9tvs+dS7HzKYxYNEywyjD
k9FyesJcGgO1rBPy+iEmTMF3cKMWOg5VxnjbUI6qOTjL5ZYgIsb5KR7Wy+RP+kUhXE6TZP6qsxFC
3QU0aGkYLyynNyIHyyLl9cVQHtYz+x8w0KmAqA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
3w3EGD6E+efCt4Fs6HRylWTDMnbDGksrBmK2LrIuuDQNpphsT/R3PC062rFGmzFuJg/bLf5Iafea
N+aHJBb97H7ueY9YF/kPUqJvkNizbPUPQpBP/2fJ5zOg61lddHncYUooATB8NAF2hcSBgU35x68X
0+ZIEJC/w3FOSQwJ1Hc=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
sL/FJO3bDIPRCCsg2DyY6eC+YEqAvN4pdWi2+bTJiJBIOsoCbIwvgrvycADXfLHet65F7sNM/rTn
YIBRQ62HHXK4AhEPCYJ16a+GWujel0mLrgVipEjZe/PIBzOTjqR8RXDwI8IW2xOJhTKtdJhHoHnZ
fRLpK84QgF3/ft41vG+L+M5INzunmmeduLlvL3yJO7PaDzNzZxm4Yb6qxrxT22OrC7GODv7eJYeF
/B+o0KrZLuu0VxgdWTSijA2jO6/yo3BIW6TSbvbn1C7fQYmUfGWF6ssH9kJPORZ7fLwb67UH+6Wy
MDlUpxP5xevODOWeiaWV5Hs+S3v9MGrU5a5myA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 18352)
`protect data_block
7tg1IRgJproBcGu6MQ9jJEvsoA69Dy1Aj2b0X4A7ow/xImR2NfGhlWV3VZ4e2F/+iBQ/5WG1UsXX
9bb7mj3qeZQOc/jhQ9N/ptyLw8WY9H5SVqwgh3Ikh1ovARSu40acpBFffhr5MUViSfTlRFovacc6
LAuiopZjIT1u6/2DPdBcRryUEtR7INYoj+RTHT9uhOagE+DJihpXedE+Go6XPADCsTGqLtgz4wU5
P2IUpwkJp+M9DhAkFYIbFwZLcu9U6vq/4PK0cIfAmsUyeoLD8J+ixDF6lEAflL0J4THMlLFQHFS1
XLuOrL0cU7JtdFZsZCzJ+gMOd9jYre2/eHvCw85ewuhZQwy0VNi7EMu93iu217+FPE4TGYulvgGW
TK1jpD4/c98xDvFPep1uSyxSGYc273VS9DHoRcwn/2Gk9FSxOZWls5SdNH6E2FOJDxoi9/6I+Pio
Q9Jhmw4KABSn33/JaKHviuM4rM84NRudapF9PAqyKHKuHf858RSrPjwm6MFFS8dcTrElwgZHc1Y6
Fl92R+HvIDW3WSkOB7ogm6OkGzPHTPKXr6Xw2kuvtHijUPuVxvNBTFIhE1CHZyKo3uD8RCFP83ia
x1MKybLIaph58jHLr34f1D4nUyLONOonRH9oE1jKGjGTU4Kmpp1eqo0msG5GSUeiPivcaKmveCD6
sKxQ0/CtKnFDu/QJtdDsJ+4MpNw0CLWWsJocQeopzlN9L58uqcLBdKW0nPE1l4eGyHUhXp7BpfQ7
n4axLDbFL3g1hbhvXcH7M6hTFg9AMgIQg0Ic2/2xUyOCT1qENcRgHwOZHWLVR+4hXisoXWCr0Qhh
D/u76jIQgbOqkUg95dV3yxzjxzMSUfbfKDCiFLU4aw126ytRY1v6ouBh2pmA0WCkt5Wc1hXFLpdQ
A0FwLJfd7PLWTweiZC0EXkrV70LNKKTihMAstxwKZZ8utewjfYhRDwgXAGWX7AsDm8uJYcyDIFkE
8rCmYCRWZNDxCnPdBE6OxSK2OjSVrNO29mG/aeSMM92LWUWFjqK4u4d7y6vTj3QZKu9/eUhLc3a7
rYCjyZ0WPcOE36Ala2y8shEJR0QqGvuyV/TU2JIRifxDAdoqXngahy/IBlrFtlsvaqUf7aI64Q8V
8R6qoa0O6EQaP0Z8Hq+JJ7//k0wlBEXN6YdQq8lRtABy5OQEXLYn33cDidLNsd5MeXCEYRsBIHbN
4D1fw5LfGKTaxIU24dfmJWY2Mx8IQjXLGBPnPFoTWb4GJ67Tt78zgAJPLuxxXePI3C3R1Gr1dFwq
20mC08NuQ2aZDe3ZiUp/5YQO7EiJRGy2nKhoCzUB1WBx8Bw2iuGjo3Z1LTnjGR0M5NdF2N2XV16Q
PBPVZDTnW0sPYgjxSrjjOHZLel6LG1gTgP1ALHz5JRD5TZO+Y2Flq0rzuSUv588rPleUse+qcj3m
sHmD6m3zIpMZo9Ny2RFKDiNez71TyTD0Y1EBtHsBk7z62dvsCQbP03hWi+6DlwDxdz2navu4r3aW
u5fbz1rPfhUK77ceID3euySrIhfUVTYmCv0bby4I6YdpHfHTwIrz7wfNw7kqNTkjSgYRRr4xMsZQ
X2knheFRFDzUvgKhTtThCZItqonxSThI/CgFRJWZql6uCyqFmAN9tOa5JsvLar31Na21FSwL7+Hv
1r3EirssL3GScEPqyFk7vlBcMde3Ep1WJwZh8Iur2zCx5Wkq5jmGi308khqyB5EG2j2OveymBw9Z
8RIChrbBI6Ggxm1Mj2h9D/cfj4+I4N5J7S1I3oZQ5hqTGt3vfNRQmWubzRAXKmxbkY8B7K9ulMHU
bZ4sUbufHdjv3AAhqBjbrdApXW74jt+3/KIYH8PXa4C/Ctth+iXfC0ylTEkSXmFwiv2plMBE3NW5
jIRR6yOwQ37DrQd8S51S3n1kB/6aojR7ImD+UAtK4I0VWCTQAWiYyJDZyQvbyqCW4GdKJQP1ueY4
ekbl47e2Nk9T6TRQYsOeTo6KsAQ1PhiXh3svVpqM/3p1LAy61KeRUcXWoq8MGx+1WyVSbHTtTWDQ
IKi/7ohmhK+uu/I2QsAdTcPel0Np9Q/L4EQZz3n37YoY9gtRXJXn0dicjsE57XnOSNNuOwmS4y3j
oZNrQD+hMXJKAn24YVoHlunaqK1Yw4s/zHfGHNRowIw5v/0nYCyUiy/lUJZerGMAyWC6/p9b8k5n
wyEylIWoCCm/CohgzAotZgB2ooUYF4F4DLnFT7rmtsiNGn4q/8pvbMPktEN3NKOzoF0oen3wyOng
NV2oHspvxZJKOrcVNmuchXtZHAOPj4Q6HekR0/Yo9ue2QkKdQfAf99nuaD4imb4M0OBGCZUW43Qz
/max1ADTsZu9+jD6/gu3gtpNH8qmwaRS7kLY4lifV+XOH2sQmeEkf8NxiOTcxMZR2aRsQWIjJpOj
WY2D2fdm05LmbMg3lk3skUTHRM3einzZsqxWK4TlXTAnVR1C5RW/JqVdOcYXAO4Cfis6gckN8iqY
Oov+s6KsityWJimWAIBAYwYJDylf/r5Y4V86LFDlaXgcls+BW703MWUmfn6n7NS2BCxpCR0TGkTX
N9KmpKJE059WvXnBmPJZXmw6bau65awyuwpbmK55GUkQEMi7v0VkWyT8ymU0hx6uAC8bs9PiMZhT
FWeq0CKMLYoDnk/lhREN1ulAfvfza5FUoNXX4HzOWIrS8QH3dgS+ETbsLAbz7ve5N4tEHN3jindL
3LbY/EgVoFiYzGIeGJzjcfTjatiE5wbChx5sgEAEYPflfhoPLwxRs+ESuAkYSIsrfRvZxZMWh+sd
jGC7d4Xg+CdfZjcJXm2AT6pRPdDo4wd+CRSP1T6Vtqub89d+ARNoOQPb9RMdve2sENk/bTYKa+Wc
sch/6xSLDlZ2xRP9/JWhuPvxXxcvscbLLDzyVtu9Fs3HcjLvNOkhNO+YzzCS69xi44xo/mjSqXU2
oK7tw4+tkFGjuAAwxzf8K+IdiN6yh6UrujnCgUXCsieHsAALUR3vC7bHYzWkgruWXPC3UvxwU+QH
elImI0n4Mi2HcffB9oIyw6v5JahqLWBm7Wz2XLSwcAx/JUVp0EjGc22uedJtjD6IP3HLiEuVpBBS
qzRm88F0gU3f+rKbhBDeqy4wmt3Rnc85T3EAmUG7H4HleFbiAG/Z4gaaRA1bN4bBZmzsrR4JgdKW
15ZiaSHKc5ut7h+SFpj7b3RB9tmogAU0BUudXfVkxrc3/JcBcW6AjWjmciCT7Z+GkA0rKB8PBg88
lnMeW+bmRSo4S8KB5W5lQvmXzUnuL0lPBH3wbbbCkzE/Z66RlwBqqUPiqgYQoL8rGcswMAEcvYvT
RQqbKgf2RblZvwZpnVNQbp/nlXIdRWiYq++S0uzPvjPgDNIA9EyB5IklIDeDtdbFtkYMqOGOOQaO
ADFPB5bh6sNgQvI8OZAh0M+HzsnU31Wk1g3+PtwFuQDSw7UHuj/zNgwFl+M8oVo+fMO+L8MT2vkH
hujKXnCXqZBITTkNInKdAQ0KUMCuaIfH1qPZDQgMczeEb2CaYZwszaC3A9iXWkxXovJPs1Sa/9sy
U5rLpNtA5vgbGOpbRjopU0MG0X4HKgPagTzRAMbpRSVtcgdpv8BlC64vuTNC9lMNZM2XuHc5rwky
U9m3iOyKTAOsRdUIG76m8sUpnLIxjb10Gi3c991+m7EHEddwmUE8bj8iQQydxEPGjnN3u/ob/z88
+p0HsMWW+xXKzdhoZPLmvsZNsucvoAsYPls3JYuUvfTBsR80zNSpqt2pK3/xziCYows4aMDck35Q
Rv1v4Ix6SzI2JhQTqhxyFZcyMQpTpszX+E9ZueauxHDW1doCIloB1kxhJdweuApGy8Y5v7Jntij/
qWPRl/8h3SFzniksIYJWHkxKIeiP7H5ZFPVQjjvFE3l23nfsTGcx8VJPFWZYItFwwQ/xIw1dv6Vp
Ksp+zVdoFadRjq++kd7Y0qhx30RNMNtD4iR+sW02mxUWvUoUzg5wi3WMPft6ILAcKoyUmUqfpbW9
s7pEVr8gPBqfDOm2IIw0q3oo6ZFcmClKbWY3JHW6jxbGzy3/hp6Zyf9o8IkL1HaGjcBRqmRaQ1TC
iJTB7w4prwvKss9+ogQjW7h4o+ZHpKSoinfFhwQQRXll260RUsY2+VNB+pycffhgI1ZSoc/UDxa4
icQyj56Ve1vgeshmPdN8VqimgeFBq/7TKVjomxN0YjQXlcslZH9rdwnRtoTX3iPHIZxYihS64gzN
1tKgoersH0t2m3uS11cHdJPeUPHm7kzqC+kltzFN8StELc7qA8f++bT86LcdoXNceIqFaUtdrsJ0
CxHHMpd2x51sLKYkyD998BCxklngVsMM2znqT1klNpoPSkbJDNY9XFE6E8dIO3L1I10AIc30wEO6
uRc5duKT9g+SckKpclDbnx/qDt6P8dfn85tPMNKE7OLBLVhTwyK8Fow1nWzCZCJh+S47A6rg7Sq6
oY590Ea4HzzC9iolt+iIvIbCa7rXdJGrEksHDCMkJkwS2DYiz8Vhs1404fSUHaEpF151pssHIVQT
/5I3fy3eM3hZ8mIWGrXENi3E7OQOX6CDy8kuLQaY6TBkOPvkEHKFekHNLURv6XBfITOX0Yu8++3W
Ea/bZt8NrF32LT1w9ShtWIP83nzg59K8z4IlCzgsSOAkDlxu+wEKTAkKq4yyhUSZG7dj+eKnfpeK
cBaOojxrpjs1P8Se990xI6uKcMNXx9PXaR4MLUywMg2gTpT+EEoBELtNDY5uimXucU8XxRud1HbO
JyjF6XS4XHunDcdDiAnsQr2RDH7zrVC4LyAQIzt9JUOSUIwo4WL8/S7Q4GS36+fcAuBxdwEYuBgz
7u0SWjpAQAlMJtUEnAWzQFG5C68U1D43CRr1hCZw06dP+HsqGXjX8BF4BWe2IoE6CibVE1+fr3Fe
bHc1OPnB6YMwHEfdZkqU6dON0Fxp0ZBPKcPYpEun16fVPL96moMNBhyFYYAMAm+peOUltbATNxna
Wg41uavepjIw+aJFbb5a8V1pEdSuVq/ZWq5NPtrfBR2EAiRwFFAKLihGruZY8okmo5OoGFCyJiFC
wHmaOHa4e3JJcJ4LDa0IdyoYhjLrzpPFksWdawZ/JwmwNMwlnGpJt0ENC0wOKHPZnRaCerPdkJEL
0FMb2norIRXxAOxGsq5hnMcEdf8+W5u4Aio9A9fNA+fkVOZHxzjiOhDvrHxBZb29FASFi3WXEup+
/gBslYkgnKYodagCdVAqYOLomjBnS9AIdzvbXNibJCMUffugYgdFvPSdswe1+5SIkpMwFR454Llm
ahlJMRXYL582WtUNDKXBHozou96mXwJeo2duUalxBGwPpLzNIgIYKpYsR1J1q3DH0TxcUdd0VtFi
2GQBymk/4VWPAslsllm1KtKJCWM4334lviHp8KXOLg7nSfxmt5ktDRVx2QyNllYl9tzuzZCWeHjs
nkB+48/8odmgcWn4gHMPuGRZO6MNeOloRW7rHzfXGn6nOcsZI2tItmOicmmmGFtJ/ZRPBaEqn8vb
KAcAgbtiFKpb8/cEK0Ok3OAR/3NnLlajygIfLKOWM693YIIwKnyqobSOF23oQhoHpdr88cd10G/N
KKFJqj3eLZ2T/jsWRE4x18gWSriY6dHFe2aQJQc1h17O8LJ2YAxbFrJni2zKEs6qgDfNT/buRp1A
PlscBUmGe9+SFK0JXNiT0jLZjRTpyvpN9e9BW5IKMj8AU+2vsXG4G+Md0nza9tHCodhdVsA5IE1I
kgcI0i1l03Cl0AD4sTJes3h3vuICl2TI3lql9EHz2DV6NxSqBCl6okhmZi1A0gpp3tCyJSbnm/99
iXuKHT6AaFxTm80YDLD51+Zkp4r7GxyGXf58nOEipbSL4Gdi9Zk/PgUl8NZv96dXbWqPL0dAyOHk
sIGuLP29Hk8wkqa0g97gqzsximtZI9/RrDJRp5P2Ik1HiubZU87FxyK/KZd16q4PD6LG2qb5ZgNz
6pRpocKQJpNb7ad4rWdN6NLJY3nBs83gFaaPJOtkgACuWytqrkMOmBhnlX0khe0qWJXsPh0kkJqZ
x0D6AnWAy8vrtvYpabKLIwOpZ/mGoFfd6yk+iBPXyisXOABWZTERLxBHxMtdGC9CwZcfaY+04Df7
t0Xevt5fzdrtZWSNV5GTgV9nSPT5uz+Ef3MWVZPy90xEPc6UpA3TQovhOsmJqh/gwg+13fNmnL57
pYBv+TNIAF4RfiY8F+qqEPo7K9mgE8VC9GoZen4/lqLXco4kERPfoKjED5hGG1D8pcS/XEqqrC7t
l05/68N702ISyBaU7qh0+FKo/SwxEXwG+5GtNq9PYr7vq3PnH40nQ1msfDBeGuD6NhWjohUBGCx6
oy6qJj5UyU+QI/WGhMwHsmgGgA67fXyBf4Ibw7/8FH0jhcwlNfreNP7oIIg2bqbWdsSXFV81Bk9t
7rqACF2IIBMOgn7VwTH6zfegiHSDmeF98SolK4V1vtlfuv3hjq+8Rd7kiV0geRMWKkujgug02nsn
wa1ClusXghnNdT2Qqqs9wJPD9BvQ0QjASgzzBccasorG0s+LbwpZoh+irwWqQ5o46ETeT/P8BDC/
iTBgsWV20LcMDMFDVsOv5qe7PHZmeENcLr22XnEWmAlpQrZwicEwRugr0PvcVA7pQTD6fRNSG6m3
T8kNVP37rnLlOcwM1TF9+8Jz8dR3JcU+/0s8XKtOVBb6AVfncI/eXVh+6lOFqeyBeZ24d1u1wvlG
9MhRGQBZ82lrlBkRRM3JWbk8XzVbyUU3QuRNpBXMCIWMmxQo1W9IIrtoPoPruc6PHO3hBuirN4a0
g7WsOJjU6CTIEr4pIEazW5wNR65ZNjmfzAKmJdk2P54PRyFnaXMhCfA1zHoGYWbBwTfBN9S1Nm9b
0+QT+cK6GV95wQSVq89iMcq/OLWKkNNjYzRKzUX0L0N4goWcPtC2kXFJ9cBMRBlErGPi7DoCzNjV
d6YrV+liJSpy6pWFrzedEb6/h+0ES3cSKzbb3JNygJHvMmNrTCkVWoGb+0IMvUo/aa8ql7mcR01T
9mCWvKHbPSiFuEtMNCQ085K2NVSZ2KssTSKvOJ3DLIuQuRfL+m1cnCHwpJh/q18PkA4ehnd/Qf1u
aQNfBKb2F0zpnItvB6g7e/02Q8CVtqN/idVIdKmUP1/PJZ+uExtdwh3JAlOMEZbFqkFMokx64clU
Jg2WskmA5FZx9VjFekgopnKjgUshSceYU19IWvhFZh475NK9Rf4Mpn25ijzsw873dPiHMa7XdgDQ
FXNvK3qFSmxqbs3cwGKcAmZxivgYs1tYWMTAqpaQ6BMkwU1MQxh2ukTc392urP1GhgssQk2FgF9E
IJ3FMFKmMjPA3dWhoW/YMieKnmt2ywsm3P3vb0cK9ADeFvIx3HQ9u3E+31DzvXbSaPKbFAmcNjp0
gm6TS/3oBfrFurUf/YQCvvoVEJmerhysZpUplWfG/P8dRMWtZWV+NBVqAYnpDcwC83yXHAEyGJqv
sSuU/IkNdb06Q73/dw/f/T7mCRaXp+Mf8R1AC3CZ6IUWtsn4yFzJYoo+LRmIvGVXJuby2obhExwt
g3n3lHC4PZ6lpRLQAQMbQnD2KRqRyO1ytfM7de3dspjfj2hMj5EyuLJ+gHLAgdMeJxURx6a+T8qX
4Fu8aK0oIHL/qIogVnM1AbxJHtbZshqKZf2klb6ZNcjCQkhjVDrbHPpdOVglwNBqt8QGT7NlGt+l
Ng+2ajCRf0xRLO9M2SzE8jPS5yByZUQbuZ0t7W++w675qzh85fma8CpvQmDR2VaihJ2evB9AeYSI
42mbx7KkLqP4HIkAle6MLIpbdDF71QMkTthDsDnBjVu2N5hgL5jKrcql398l4R0aT0IqPgEeqKB7
ugrgNfftP5nzgaYyONA3tiIAtiNn+JdsL1TZbfQzuLAF1Cd9v+mGc88mPG+Sb6CpFXpOW1iLcLub
m5GXtaZE6S70Qc6RkFOweoEveUAjciYpSbkkK42XokCUkjHaehwwmyAkg9rHzUyX4iiRVMrXzgIJ
7rwUMaQvgeJHYSFWbJO7BHEzJV71tkcB1H7M6QfboO379vUN2GYl3npx4P8axmPd1FiwRXsKqCVB
BMrCpJEbYrW0AX3Z1LuGgGbqvEXHMSiC98MloSiMPGp2l/IYevy5HAh6iy9JDKYpxFVEBf/mCvLk
eYFQPMYZ/4FWUOga0GTO7U2rfTfpJq7K0wgsBW8/KvH++uqbMicOznIFeEpIO327zrI2KyGdC9tg
YN9y9ZbjRV30jFlWvuglLRIDQSNhaZUEPqj0xV4Gh4NAABUKRptzH9O/3s5VsDE2baPYMwd7K3nC
JrjFgqoAhSJdbBGQ/fK2ulp/WnUQE49xz34yx8VVwU2UvrAfSyJAiH+dZXAslr55VEle968rnIgl
xCZdguHffEDCssncdxKSem+iZdtFCDD7+5kYKFL/t0jyOEqijt//1lD8dJLz4UZnlv4SLlckP2A7
f9ElBc3Y/GnrqRxnriNzLSHnbvGV63rrotBjCZjouiOAkS7qWJcNA7LPVxS10JUwg73IQu4cw3OX
W+KZXJx0KCPBSwFcz72Ux4oqCWd6r4N0m3uzDZMZU2iWfrlewIlnfPdwx6dOxrcXfRd+uTtJpyjF
OYSC3gxRxWkKMM3OuXyS/OLDqpeUnKUNXNn5sK/Lgt6Xla/XDJKamzFmwNVQc1KmilMkD4M4xIjA
cbt9nEv6teH/vXrhAYVs+ziKoA9sGnecXWm1TUm2V+Nz2l/X1ZSV99EXLcPL4JN5xAM+ws9g+2hG
ZjH1UITWZb5BElaoJS4O1Up4yu8HsNI2cOkrdm6nObdpR1qlVFK+Z8oG5+P5328L0HbaM0BY8s6U
82msC0dEJH3isnWvWwKQm+2k3PPemjJ0Cp7UgXy/RjRO8D3GVoWI7gAIq9Y3GRsxf9OaY6auYtLX
HCx/9FCq4oA47FUTp9tjUbo06FHFa9uWxh0+22qdob/OVBCOgnNyIGT22yW/BS1grokXFm0K5DVZ
4AQcapAWZAZElDJXlhp3FfZ4TzzgT4EejkGiXJx5BbOlIk4mjbiRyLnHO9Bn4nLjCdxJ1Udzq/Us
0BPuXw9iUYDwvupDokN1xOZmH3ITVJZIOudV8REIns65nt6DDF1zc5G5w08oxx+cx518uZKlX0+u
/atcWGE3UHU89TiQdIK90LdAIL7dnhPCun6Iq0fEh5JpN8WXzpCXZ6RxqDzS4pfBB3cgLvoITOpU
ZHocqkzET+7rK+3zoGD3pmPAu2sLmzJfcHBq7Ns1Bb8W5F0//sY0roBS7PeF5vDDMfAlgZ6Udk+S
VN9fLXprOdkLiDguZBCNdi+mxMxca740b2UOTR8q7JRWYJP4iWbLO2+LPbKLxA1zidDFJ+hMHmtX
Y+DoaGISDjA4D4CqIhWJI/x9uZZs18Te9Gm7u6mDUmgttqM5eAKev3m7uDZjbJ1qEq7FBMnZLcZu
SzjxHNkIz56p3TOW3ZBubLzBNIeTbeoBYWqtzPyr+er30pjfqfzKpXZ9ipmv3T6XexFZOBFPx3AQ
YLIsm9BtNosn5FQajcv2r4fKQS3ZjWWqQIGvVhfeCC27KclYuhfU776PsX6+Ey+3mS1ifJYmTmNn
hBTT+qKGpxMLOmLYmVvTvNnQfMk6j7e8zFshcpXtSz5VipSORdrIdz4Rs8w/5adSrsZYpxk5GkW6
71X012/oXHVymAsLBehi4jDAwVUKpD8rGh+ENrSesmUbXHFJGQz/EBTcxC2zkQ+COkPrrbgf5En+
/DoG2jqkG9IEka5A9NmAsoYj9hKPHOvJZxv2aJO775uAdViJWdm7qpNla5m5o/aYL3P0dF55Mq/J
uwdrdqdHHdXZJSeSbKLSRDnlykdaoSF2+XtHJ2iypJpXJzu5jO6gy0UEC6bw/4Tum2TryOUlRzXY
zmMLN3dnE/qHnmIll17++6hZRLp8LefytLo/IzL/o6dB/+oELC1dZYleCY0I58R7KMiRpzRqjKRB
dX/MF3Vf/l2Fb1ZHYl/2r7oH4j57Pqrvj0nHu+s+Xw4EFYB8axAn1vBlvKSnE59Fn14JUz0zvksB
tAUthm833dIoWJ1BDjY/atDQAYF0Q4/Rhdo5ghqyPHCbSl+fZWKpUhoqC4p/YyzpPWLC6H42NlQW
BQIBz5gG6/Ya5f9iiPl2NGDbgc/Oj7bVQiaRR4JAaJ4V+eZN67llN1QIaxO+djWIBMHRmmxo/iRx
yt6rRl4hz13Ixaarq4ryQUKJVKsKEC2cR9ZDku9k7jlHPhf6uqZB2vY7j+XA7wEM5A/2ZDENIRbl
spdcpTwtJnJNMY1dXVxxuMg3nixARIQXWU1ELp36ABo6L9xugV1Kufc6Cavvg8ALrxfmv1s2Al/t
YHnmzDhY7qseTNvccZEh4puYbcqOmLjU3Lub64LulZUjR53AkvqZ4ZP+h91MLbZIzxzvJRiicE9X
yu3I87gSLQh1dgcedtLrXDIOcp37Qt1OqypPcM08uLImiYsreXkEFD5qOVtE9dV2kwEZvjHvtnRd
2X28H+hHECuczTVOXgs1OwgPmuo8pAikFqjHfOK6/cqIcKEe0ZvrmTY5pjenK2rt4U4YfHBWv6mS
9+oMvbg1jv74xHl28EJdvl/f5IOOwoS+zGUrthLctbK0zMe/CUxjPmX9ljOclqllXDQIyeAoQJnX
ZMcBUer/3Kx6mMvWBOMjPSx6Pc8xoLLEtU3oRCt1bij6YvC3GmK4ooMyxq79kri5zwBpkHJGufoF
OZe+5jOch866o9d7xggCeEwkOHyh9M0YdP9mFeXlQG1nCB7/0FV+6iMi9yTVZ/Yamkngwo83u8tC
RHpXQxu9qtK998OT7gj5m1cUhvt6LdCSusJZ7fVgIrYQmIAaoxEwB1562HeHv5GlX9Yo+CYuoO6v
SiBZjYE2jM7yjuFRZtxKL3T4dmiX0h6P/HKqsxccej3VleOnJ0rGDrgcQ861hFEVwfLItARwa5FP
avPqcDJrEKBhTC6PK8eJVZIgt8YU0LhZQ8bGSIEhQfj92DAdYKTlO5/F95Q1kkofIJPe02aQi7rU
EfAHnuwijdHiPX+IuzkhNOqFSqTPKvRJIh6J2F518MDxh0HL8YWoyN2y9pTpDm3qwkW0+zS1I3dn
XH+AcqiXecqYpINCve7TAmuUpXaIsKQS/LqdlnsiaPxacNb/r2rkusOQIccsdcM1LAY6udAGnOJX
O6OrfVTSYoylsx2zdlzevKvb1PBt4MEEoN4UB3hseHWSYUr34/dOcq90D3tCycGmvTx7PSg64rTL
D9uJ1mW0kttgzGGVm7HgMwaSg0oPEyMI9+61xDSsSRLx3K0HKz+3tYi3IC565ToOOMP5TifKUNfe
ZDuyh/jhIA8zdd6BIfgMrAZT5E5vR8on2Lvafc2jTl+f3MTV5G9gFn1hVkJjmiQuWqmjbYZDVdFn
jB94phq8654KjdYc1bQoVBN00So7o3hA3/EVgxaxU0pm2Fp3JVJmgYQElj/h7pqc2DJhQJ/blY+7
AenFc9R+cj8n9VcxawVy24//rGmEAaFy3QglTlAfcPC/2vBcJybelJCJ6ka/x7fCJMotQ9wfMW06
Osc0Xn0peMpHmO9OW2odoHjqukvf9d/1pCfnET6NufVXlyjmUXk60owG6rRRmVgPoSO7bAdGbEl/
RbFW1Av1wVuhYIQSV9uiW5wFX2GMgbNTA6y3TSRIwtcPz7uHkvRSXGqq7yzTE8tGWoYefBeKFbwR
7z/+BDQcuq7iCcopc2PmcJPfDpgyFo0XggZMCgTNFKFHfPkPHiaoS8b8F7D+2+tFh69FV+SY5HNi
4vlkSo7dTcL5NYCFlxZThYSov1TM3Sc1H0uGeCOER1X4SUAAWsSc3k+zpQTeWi5Qe4Wx0QIneggx
rkMn5bEpS4lMskRmJkKX1LRl+ZPLHi7DdQDZsf5QB2MpYDV69uCCwarzE/+28IF3BVucACcAsE/r
bcNSCaVEJZmaQyQxbzyxRPb8bmFm9xS52Ehxr4FgjVu/3LwckimCIw0Lr+R8X/lYjlwz9Y5zNV1h
0YpsK/lUFKWX8Agfy1efmBNncL/F3busKvzFURn4qhCN4bVqIhsq+vqJNvXMGn1eClz9cJjqebvG
sCb31RC0Fzaw/2PflZrtu1aNuiSzNse1BTj2kjbulautuzkH5Zt4Zf66Zu3l8toYKzkD2dyF5fRz
w/SMP7p5Yw76DBS0Mcc+1GzzSfTaD6KyrLyQuQ/O8+ncgUzUufw2bPy5w73ObIZs/5BjTN72v3vN
0MfanwadgBYlHHp0b+uiZbLpbiO2ElyxP2FfSvUPHXcHQ+Iu3ddsOgS+0rEHd6zspRmV3hbXdkgT
frwiqLafRP8QaBlVZidjqEgP5d7sHQuKI44PmZlkKNoCNxlgGWHWyklqpB1sKExLh59FDu8SBZ+A
tRxbeBycZ79ivabaBuPpEcL5JMlT63Huw3ecQG4GOd6LcSB8PxdcVIjiw7eg0Kcei6kRrZZQivfH
mJy59jGM2LvpssUlTQFaFbj16rWsexGBczmxIYnG9eUMQp2YXBJRFiL1YCnsvLgf+4oJ9oy3k+ng
gb2MFhqbaGqHuAMg6pYkFJnlA4A9gqXmGwbHB4JHxAQitgRZmtvCqZXUSXftRq8YdYeT0pYxz1n9
jGnZJk6t61inSJjWx/yNkwsNpscj2cWxpwkTEneDpOw2256NEnZGSTBAu+u7UUxUWVbaq3XuSzzL
UFkeIr2DfigxODhrAWYfSakgxaByfaaG9Fl2UZ2pwut6Hz9IM6FHKc7UhUU5bMHWJ02liFg6eRYm
uUyUF78dqGstnAvI5hqvUTCmu4JBAMwd47t/dw2PCCKhSVQn1K+sfmbV2aPgcfZ1bxcVXwamYRu8
LjoqgxtctBEON5nQVJP7EJdCbt+qUUWBVY0kX8dwOcOYZs7BohT/EmbXz/kfC5vxPbAj4BYJe1H+
1tlnNFboniO1fogq7JpFLNpFxSVnTP/Ras2CuhQZyfRkHa36TRnvyqMs/VUHThSlvMc0UaqKhkxe
xYn0rs3MwG+zt7ZwiFfwz3MggKHpwWqUgecXGGd1+m2g1U4HpcGIZeh+LZQZsJj0M3yMCTVIToZZ
6L77SZM0htTpElU3TPLSV0lyzGsBKa39oY2uokpowHkjQHBvdT/d6bpoCURU9+lxhz8MyvLWp6WN
GHyDGga2h0vZlCXaB3M6OAfxaTBP6b5qeWxd/Y+wzVaPq1YchPoOo9K8lmLipCSxCA98vVA0ZT7+
Hu7QsrMlPfe+OOyp/i+oUStQnmaeZ0bvlfTlVuuyTLSbdION02UipZh7QOzrLCaNHegDt6BXynR4
BwulEzlu525sSz8HHVfc3DutPwL8T4Cxo4LSGU3iAfpX+EEjrGmQ7nvEzE1854GpAJDA3UiIKfWw
g06M6CQ87pfxVlfeVu+jxWgZKbjtS7pQQdhGOjyye3H6AEnBI7BVjExCaMvTmKpPgDjF6IG9O6Jp
eP+MarrZx7h15IL5f9qOQ979IJdUs3mFCu79JNeS0y/dt+po6TovbxM+GG4nDFmffLgtf/gILxso
znEGH+3t/xZD9nNxyEYP5kyR0C4cgBEgQn25xA0vIbQBQj3b4taa/KuhAjEf9KNVg9wI01SZNXAh
Xh7/lt9TcIw36jmjHTJRKalmFCswCO3SDRnj8c7dridt+zGdnaujPDoqDvOZa2Yk4F2l7lsSH/D5
lOGTP80UJmQA/Sy91kBVIPNtXeNjaf9InqM8uO3qo0bVxOd1dpgX78YV9ANXdkLl+rkyyxpBlQcB
q/glIeRrEZkFJbON3kBG+qWgMtNW2/cSzU3L0HdV7Louwc990nhXfe9Osiy06R69gaJeuZ3DdGSX
4h5fyn8oqTgkJSpZpxDrPxQ/p3sbAO0ZZ86pAtHW0ZavSca61vT1MZ4jyeRYuoQlFkju47FXyKlJ
vKnaTJj4BlH2ZfPoFrUiyP72F2W2S26q9cfQdsN7AQiJQeR1fd8ZB4NcbRqvE19a84mj8xFe9Ypl
wcExifIVJzP/beEdjLWY888MpgicB0qwJTCFkqGvAI0eR4lTPqduBo3gtODV4jO8MRnEoMbDJLjB
6cRDMyy4iPuy/vA+F2n0aPKjzAXm6VWIpdxumIw7GAXf8H0Vxy7qCFmcPFU6G/pafFPnxFm+y8+1
cw4pN9LM5uOoMpo1X3Q2MnVSBpag1Tzbl6q17QSvCUuu/J9jtmLrXz6FDQniLQdOZTzx0wRvN50L
JJOko4YioT3ISFTdFnGXmQzCHhfm1hu4NwEXjDED8yHUi0UlezyD6SgywubsYo2jisWMr1GtwGB9
jGcpHhdFvSwivXhSiYLeJbL6YP4ygyT2tkhS+89fx7lGc2yr8MKBNH7gF8cgh4QQugGI/pxhwzjG
wCICzDGDOb3xPD2Xcd3mLZLUIY0p/OHj+Dc0ZL/SQtaQWCvxJl1mDn9vCIMVDr/jzkwvjUv4C1Yp
q9nRIdvStX3z4D/yzkMA3JBM2LOwDCqb6z48GB/NIlxK20d4VJ/1UaXRrHg9sgQAbL7D9Fh2L9hC
oN68fHWJ9O4SX2HqY86AOqKCSDQ0FM/3lInFY++r/tdwbRbnDrJyUTJ81VFwMISsXxXio9hMTgch
C/CwtYn7oe16xuCk3egilRCLkCA4C3/YzHnlwIVE/xm6VFlwzepeK7s89QwVHaZjtVomDNDimguG
ZhSSPWqlNetv6Dii1plPPqqRHrXg210aMWG7FzugTUFnmNFJu3Y7zMs4tOl/Fps8rkNR/OGW2XBs
/BFtTvwWfzf6t+Tfo/rVviT2zZO5o7epSnwwO0QnckT4d0sQQP7xacPZBkutQdpGjgBPmVUu7AlG
sW62KPrCwv+7b9cmQYlMuaz90LefLlGQksiBbioP/SkK7phlfqjcDNXqgY5olbYU+m9rIwzY2cNi
UXfeVKmiyjHsBLUZely8bobpBNZXy/goi3CVrB0RYtgcYGmXnUkaFp+qeHZriZLuYkmW4LQ0gvSU
VtHgdhJoBP1IkWI/5LPT/gBUugQECcpyn7cywu3kN/QOazox3DzmwhGrYAJ7Uawi/hQxXHPcK8Am
2dHfUA2d4rFQl1iDM+EX6rV++qxn2GBZSpqDK94ubQSp4hP5BDoCfl4v2CDZ7va2FESRHViSg1ZO
rs1215WY41TqcSUoh+MpLgAkNUCgrDYsqDjwN8ydfIvFG2N3Gy0tlxGp3Nnd/Biel4dkmBhCyGoU
oPu3a6nnKTDUk0zVyDTNhonDQ7QDnFPUliOt8YyRoyxH1YGQQtzQ6BinpPY3OyaWjeIulKNi57uX
wlNcuQUxXnNfa2JYWyyXvdSNi6c7iFHECetDLtytI0ttOtJE4vQH6F6KoYob80DN6r7Sc51EDYm6
5qNn/eY0V7hmE/Z8OJTueJkO6wr/R6v8ichQEct7z2w0O3bkO35/1ltzkFgEgiLQa1C/VZOraVub
Shdv0ltroAP55sHxIsnC3TjFC2grRoMkyd6qAvsDXtdXfBjQSYcZ4YqsyAYyQnOxGG+pzYyRmVLr
BOAfL8O1TNuTsRf0sGTJdhgfK4+3aD/rHN35UIiDPAlTBvowjiEDu6qhJgKpDYRE1LUcxzD4gQ9M
ydGTeCo+CCQdbibVji8k69aQBWDH13kOSEYN6K1Es8rDEB1VPvNyfsOFLl4DxOnsBu8iTqX2hw5d
t6xzMD+ZlK/wxg6xR4Hgj+vqy4VP8nNO5BbG3Gyrwwfu8S2UEeKhaKS8nX8y49TubhaDpDObfpRe
0TKEZlIX9Zhe5KXoHSAXpqbZ/P6phVNoKfHfOxVdP2LKvv8rsom3UKoHDhCubMg+fJn4LogEMGL3
WTn4yoUkVsZNAIATv8BDKPbWPiwhRTxFpg0y7M26hGKXMlCNrqbvFMK5NHY54YNFJHb+vn49HIgW
1K6YdqDJby4WHBvQQY6FWxEKO1xWrlJJeiUpaMPMALEgWzAQvC0QEykDTqjQ4+5t7LxOTh7wI/wc
kn5aOabzkA4NX06NMrapxHRWA18IFx4JGN4RoqzBJtnBONBja0qpud3gjnndNfjDl+MavYxgoKM+
QNPMGHKZCvGT1AJV/CKle5qVEglG/pAnMbrXFyTvEn+sRrePqwJ7db3OQ3bN49HcgVXf6BvFftfs
2HwHUL0lB6YiBUaz60lIJM6G4As3wbNQ57N/AmUVY3Erg3XFWbXdQ+AQl5CTUJxD/feoWB0tSasq
vEYL2+pEV8DxaV9SI7x3Y4SoKHQ2LESo423z60cs7ktlHcHkLqi9xSNN6Nl1f4JnPvIUvb7IeEzL
2bZztdUVc8RTbtwOUIaHtkaNKrmvgz3lYBjpDw+u0r4ccAlesPhaQ6+rnt+KpzUp0S/4VbVVNdj0
0rHXgSxOEL9edqCMh2axyCS1VYbL3IzTRFYCuHMdCPOKUMfqtOc4x9rOeiJ4eUIGt3k5fwjD0TQQ
CpYEnpCpuqXNMxeUhH3PHLSYQkSuB+tfdwmfuk68blYahxFFypogiTFKxrPHw0QbfmB/J7p4ktb4
QV/TT0hv+Xd6SIcr68n92AHMaBad/233Nii5gka3IfZPRktH6MYSjKqOd8oEP7L9Y58yQDI5BpbC
LZT1mSWwYshznQBJk3HYyxmtmunbktaFBilOOCsnIJoNsNOk6MA/l8Dc9n+APm9nTOm6o3p6xgg7
uyDfLPA1xkFvNvti271qIX/8otqubZFg7vwX9H3oworVjW66Fb2A8i33bZyiBf4FXknk8Ikn852d
RQf9HB3if/oOkha8bGwuY0X6o6cf3jwt/WQoOBqj6uAfJRduPoPEC58Ya6uXiR/RoaNfIySIlTKm
WJfbq4z6QM9wd3QnPLn+cfBj81qjzlh8/6rDrwC/Fr6wby+dHmHpaM8c7xJWdyR0r2/ZzkejFPeU
Yfs5fOqpPzbpARBlVKzsIpgsxeiuQEFi0x/D93qPV+x8l54XxV0dml4Nlps5kUtlADU7blYikpyk
/nFLJA/HpZl+QSZNgT+xzRYb1gp0rzYhcYyDBRd5EmW8RPopH0GyldkaZR8MSDGL7zVc39wpc9Uv
xl5F1VrtnPHxBh7z4fbY09kzEcaqZna3tYey4iwQo6GgrT3iR0Gxi+9AKgAerUzWHK5SOKkVZmzX
3xm9ccxfNvz6mmOl/ykR0TZkMTCPK/NVoXZMmC2ZtEZe6UJdCS+KOFMYBH1rRjRGQusQFO8N5IkE
wSb+VYTTCkY0KUnsZwzTClrUSZt5tP7eSzDMaAYZo73YfwIA+BWC9eT9lKlgY6VSaVg8Taw5zYbw
gLpjq362FNkCT/gtUsfqh70l/ZnTLTuZcLuAusaplUmNTSp14OnG58uT5+gM9EXxWPsNNXQLCwC3
GBdFKs13s3IItxm1aiVj1XTwkxCe9Zwy52o3dHPg889uHhQN1pDecnvS+KtfWf6r0A+JPGUmTLU/
Rp5XBJCuLp3x17kCyklF8Ae++9ewyfrN1tXLev++Bb8goUTFufuIdJfpuBtIgarjn3y3PEGkCGXb
Lhzhw2IUTkYkb6yT2vaSfy3HqV6SiKnQ1ZAR1+n/5J1Qau4OFgx0ZQY26eex/GG6xhRZeVZu/WF8
EGDlyORhE/C3IaAWaTXap/dqNtYmiwxNviaCuuBh4pWxCZqJpxBaQT85pbsDnz/gVieqHVCNz0WI
qF3g12sWZ/5qRHpF/3NyOBxDwz3AfUL0vkI/a4daLtGPRv0klJuPVYBLs9t92yDsAG6uSmzzkD9L
2GS7Tq086suYWAMQkeHu2gxociiE5Na87p7U9NZboonEKJt9rrWAVRfLWDy3KeMVYgDOUJPi4Viz
0fFL2lwfNsiLTGuzJqBBREF3NHZjq7oXD9pNE89QX9zEIsbl4kyoCiGTWRlrHT/RYq4NcF3NCZiE
WLDquHWd4+NR4tvxaSdwfl3C49KfxSxkWwavoD36lqRHaAFF9jWezeicOWHJspHAyOaDKC/W28FE
El0mbxj5rJf9ym2r6KO7K+3syT/O0LeDVllO7RvG//n9rMhQUw0lRoG/LY2scIOWg39Keyy9VroS
n1j4MAotKwYQCj0995bfNQH4DL9y8Ozgb3ZWqJN+vurGEycRto0nr86kVSh1NMUMa9vnrhPuqqhE
OqZbLP3FbTginY+Gc1tBZDWuLH0KRBAcgbgxIJ2C7sCrdnHLsAkrT/e3sOXrcPHIaYMo+1wzROpv
3UMSl2yxwVcWLLF41U/vX3MqztByAMbornBm1njpUBKd0srOxnmCfd83JoSJ+dvJ4S8nhTX1JZeS
5NAtJswLVbFtm6pSLLPhXGYBVBcSBT4wet9621LfYmQ6LMitR9tZKIwUeUxDvp8b0Y69N9hSnk4L
gxCcvxdXFpiBfKmrEE2vKPG1qLv7zsAfmS6SRutELHGt8fh6KbEct1W5nS1Pvx3XKrkcxLtJLS/2
tdl30syqg5NkjdCxeSQcBbFUGLLo3Qp5N7P70KybtXlmzT+ooUExsY/d+54gvNdF/b+DI69YDALJ
ZsULB9kwh+xaRMTR0rpkLRBG5ytWYBNLyxVcJ3o8nraAJBHTSmLmrisgD7DwYqsT+4jJ12lJnZWz
A4RvRqO9qSZ635aAR+e/PpbF9UWYPLjnaElV/raRelYqnh2gsCVK/Kn53135m+gaReBHTxWlQNST
ODZsNH60MMIl6DQvspaaZ+ZHE1iAGY+PYvIy2im0TOKToHyl5ukYnVf9o6xzwzmnT3LBof9DKfUP
yIhuIjIyk5aOHCXW1ZmMscABJS/rWZ4LHyVZ6zcXMaTkdFESp83zYjwIYIIz09/qWxAIUPjHPMCf
hKkbnJidMQwMTISMyAUWm8IPYYMfgXxoVey3BYmUgIG6AnEToqni7zJtTGpW/keK3jPPYUcsxaW1
ffkJdzX3Di9pdvjq9ughnmG2UC678t7avflPCMVQeJB8Ok+m69fFfw/E62zH7jVmp7BK06BZuwFy
Y3cGLx6LRH0x23AxmP5CF5plLXiFHNSD13iPXF+A1v8Djc1xaBWH4ZOUKbVaTmZ5mA6urRrQwZ7y
+y1S2oOZyG8udXcZbHixKeoGuSLZlAu+6RAdcmxNRJ+RbkzaIw8FepxtoV3vGCYLNC5FvmSa5nST
pG9EYrc6THwD8V7bM25mD2Bs/wvQkaQI3fWCls5/xDPBXJIt4gD9COuqm2+e5aqAgQdESHg83I0x
yDVTOQIrcLnbKbrPAQAgUCD2SUNM77CtDOTUBFooyRSco2p4EL2/AAr3AG9a2mUMbv83ZL57/7qp
/BYUlbLW6424mLeZmr/Az343Erxud0k8H7KKVok4HCkOahDG9xaiYg9iRcOwIPScusQsCOIfswNa
tv7xelOqsF31c2IJH8zVI52xSYDnUkGz7VDOgG11NsGaDLEqql+wLihNXP4+uUQ7Xcz8uOWifQhF
MysvwSk4JVOcG0wrNBbPawHpyADTg5g6HQMH9ecP0JoqnrUpOlIawzU3/5ar864hqV+6vri5Xl4p
tA1RFanmM1vkgEbCEsG569lRBAz/JaPxNiP4yPNH3sj7Mh7T0Fi0vPbFfzHyAm/lyCFT3ukas2hU
SiwxC9h9MTNEV4x941P9sCxTTenOLbEwZI/ImemSY5dJ9CmkHzHrZ8diKDMmkER5mD53Cz90Wvsn
LP8wzzKETGEbSQiQRp5PWV5JdJSPZQwCv+Je+9STU5OR5CPuQeFeIYVslk3Ex2pY9RVq3hawckbD
BJJ20xsmEN7wcckQGjYBpt156/F5YgbsqO6T8Du3ZnVFGZKu4+5zQiyglmOoicjyPmVX6Y7P82Ya
jVrfPjVavB7ZQDNqQXBlzA3WZNvXkqjsskNPuiclXl5nNWNf0JpLtrn0MwBYYTTESfqxxg0iLxdD
h0f02SagtS10/Qmc9ERks0zEpmma4hvIMACyYqzAC0U6TiOZNxtV/jBGJSh1+DqyUQUCCagbJwYS
UdlaoLtbfeF4MIO2HOOxkLxdR0fIhwC8yL+P7USDxdwvHnlqJTiNneB2xhDzlNHK/PtCrtoFVAxC
0nTcsOJn8ltbFhqV+XylTG1y/Zh60nxb7j99knZb6c59jHmKYclWICjeTkqNdDLfzi9cMK/KtKN8
Y7n3sr4qrr99CngoDPd7+dN6hmzqak4GToSHMUFBj1mwNPFBggEtZ1k16/cmv8wXcmUSzannf1tl
K4Y0xPtfpwPgZZx6SKfWY/zcJIQuBV6hpWwfn1Og4wPnbd8U7I62cTDPiL43zn+5t8Zfxz+XG/1d
2Ze+eRv0uUJK6Dv7MHUmMztR9nuWzk344Ck2SLm/f3L8xm5ZyHo2PpCfC2uJZXbKZgsOPMnNl0lw
ve3zq7Jwe2WQRUd0xzO8SyIBqPvHPjJK/FFN1LVGMc9hhGLj0VSorugfC7Qz8TWRExPbTC27VlQx
WhWJEUTIkGKqgVo2rhvbkwSGDu4cK3kau1zP1hCmKG9sIpFRFRhcTOAzhCI9IO/D4QwDUgHlAnKH
LOmcsgCu9vmAMY7o4VyH4z6EB42n4UA8a5ValP6mcGGsyKjQjNpjsUQGCDJQ8ocqJJT17Uuzj4VV
CHPWlTfuEPnc3uGhUtFhMR3zE3MxyzRgzuAyNKtvNG9tMmBbtZqWLk9dPFrxyF9zt0hO0TjMA1wQ
JSXT1m2/E1o8pGO0DjxOiPD5CO6Co7p8ZNYS8On9ZYPQvoWgVUhnQKVzhMc+sDA86XW6ssI4IXYf
N7T+BVAa+KLqIJi5lkW2SpogE1Y1LBHloaN0vhfGBwbUP/jKg+YeMWMLrOuC7mKMj7fs0bHWkKGg
Ea10D320Laku/RRUctPBh+XTx6aqdDkKj84Mnd78EqCGl4PQ73U+8eDX+eXyhhLVmOhMsLw+UhH4
AElwedoYlLzbrmIL74KhSO5GKk3No0CubWcXh7HJGpy5hbNxmDJrVxhoVWA8rbgqyQDOsPUxH7Hr
X36qeHPWb8Yk3jKohvpCzE4oI1lKi0UgjgaMywtmD30VPQojaqBcLgqXaY3yvmFs0DsgJyehhCEB
5TeFVZmKm49jq8ysBc2FFoQl3FzfM4yXu1jF2C9ygo7N9ZCYzP+jnot0chftSjEB13fWT2AGRrWw
7e6EEVgGA0QSARgMu2hvny7wcdbw3Ruy4KOLNsT8FOhfpBMsXpVaZMDmN2zCI2BzbtFMLXWxUZx9
FciVTM3PUPYALI7ribojgGIFIiAmWrmT3dp2OdRVnBB9V1q5FQr3XtxQRtvHrmOvIFLyvU7izqmt
MTYBjpRe4c/qAYw45cWAhxEYmw830SmCfzj3W5cTEBCuSm1JAghGtL6GtR/46QqWyMOFzaHx4R0n
kjFkhQEUoQ1xl+4SYZWknOCbO/iVC5JT0z21RJjFnEONUFF1zU39w19efVPuOE7+Akq8bYVFV8Hg
S3l6HEZ8KjD6i8FOkBQHUNQfqirhzeXH+YHTlP8NQZnCV03x6Pdho9SxNrj+cadLnq10J4pQOR+C
w4ifC86kJPGDDrXFzL9j7cys0PNDqNGPWRRbqaRc9E8URLF2Vs6tmSVrDnCmP4neq6Q8FTZKb5PT
RD9I+ghxK6MA5yk7xQilBfwIOiuMtZ9kjHPxvldnHKSUKdW4G7dxwhsWQmFg2IV+960+QWSZ9MB5
C6SCqSLm0G9g78YQHfvIRQy/BsaUZk7cS4rkxj6RAL2hAE77oCZNcZUrnemlzhoGG+MHRKJ0X08a
wCVecq4oZG2BSwA9eFf6kbKLxFQ6F0eOWnG0EKiISjgRkCII5/cemx5++2M91jqAgAJSso5bXp/f
NarivsuSHMz/nxOQGoSsZNnXFu+kOL3ERjaJHnwWKA4e+yTu/r2137mRIxIq5uP8sHIw9HLQBoPH
mEjBAbTZvvXyr+1+xFHM+MeKkBXHnqHFNnwFpF2XFG7Wd9P3JMZAe2vZcwBN7lMEfXP6QTcZl9YP
Z5Q0H/JB5zLaYVCfBWLGC2k9aKAfBp/nuKTIcL1v33gzXUpHFV4MIyJKMAtV6nevA4k8tMNDhLwo
MXCTFQxLWAbqmIH1eddGqoUGQX6ozjMxOZFVZexbYvjLN7EBPombmcy4VR4erXTtg45Mr3JN7Nrv
8erEuH33JHOfMW2vSEp1IQQbheMfJT30dmd6bc/BbP9SCFQUk6XiF3EJ8c41vxA5YpYyBL15tDTh
Z3g8TXNR704NeDpUseZrkFA5a7E9KD8qUvObRJViDH5OgCTROfey4wP3EGhdaj1My7j1llEcZR3X
/h58FcTtofnuAK/gyIyRzBwdrmFjY7TVMYjVfuPZjteC4Th8kHlzBimIQkotFTswXcHZgo7nXGyj
0Jt3Xi/74tnGsgSVWiT8qs8aA2/b26esJNDc6iNJOxAmuTurkVQHSlX+PFhw34CBHJE8tHx6tR7Y
bK48X4YXpv7RlNKqyRj0ef8nn633SVFubSGc0rAG5eZQGAJvK5U8Z4n05IpbwAZVsdxyFX7SMadC
IFMaSX9/Iq8FXzj7nci5UdOesYJDu6NDUV9nK5V8Q6g3hmXy7U7y7Dzp3I+zPUbck9lQECK5i9Lf
IFVmIX4cEI4YTM+cSp95mc05ZPrFe0zFaegqyRfXLiycMMiOUVZq7c1cZzxgoyJl1XrCxfaCFE9Z
35/YNNmaCHC/Ui+mNYPiSnpJM7YVSGmbSt79tMioJDobK1+KqY4Ls/8OETxqrkNV3aW/wsqMXeRe
Y2NzLNXiBNfAwHuAAC4ZZKgRk3GDKY0sCLPnQrK87GLjqZZRhqG2faQa5QAtMZxtMLR37sPkoAtm
W4drBo354HA621bgIhjHGopxJytQ/0VKiTGJC8xs4Pc4DpofpwoFAKSOPZgFvPPuUdKajBYBy51c
MEorlBvK/AgGYW11tndBpV1Wmr3qFtdqptsOp57WbYhhvGla5emD4VOuB6WQCvwzfVccSJDa5BVp
96Jir2fo9Mq7e/TG+90r6uoZNQG+BmWPWFSr11ncF6sKPIk4aDrsB7lHbIR3nTFZGbk4/5AZ3CGc
d9f0SArj4TvXGIKOklrJml7EZQaFDVbQz+gL1enDO6ds34YtRwPLtRRByMzV8Ws0QQn4rMuQC+Mg
Risi6lQOL3bKqeIhdPWTt82osJCRHGhHlrLpMTwvgIYDsDTba3PrAXHbOrX81Ik+B5iT1jYff53F
eoFCj9aAu4+YD0bfIdGJ/MtYbfBsE+A+PyHonIyJBWbsVjoaGJN/ijolziH8FcC56tpl6WY2qvQH
/HfQixUxN2Z2qKLTFYy99h73liQnYZ3X5F9hSDMedzoXdTwquFJzTOy3JQuRs/siSqwzVZ0wx4ta
rCqv8ENtZizadE7/DlQlsSm+ErHdtaGnwSGCZcTj8aN7JfQuYUI1s5xu1OpYh1ovdfwMEDi9Aysg
icDuLn9t1hrZvrttsr2mCVM/yth0CSWcAgbC3v37jbiNAgEXO9bUqR/0I9c8DX2wlO7UpnSYX9dg
5Cdr0ILCWEr776g6/gk4N7H+AhAntdA+W+W+/s+nggRU+HITjEqhr3n83rSTpjqPWjdCy3dzSCCU
OfNycF6Vj8BhjHSVfoiFq2SlOqMjwqHuLRUwteiLH/mq/kFLUHl2FSB71jRdcyCadZ8O+4+IN2pS
Diuyt1AqpwjfO0UYKEyR2BZ4pUM8fZ+MO5NIoTpnFNNXCi+2wVOJ7oNi8s0NpjvhywtpqRmW4iIv
q+1stUHoGVOEitu7K8FX68oGOtmL0NWRMG11LDIYr8gJkar4gOXknofJoIqRQiWqWzE02LIwkv/t
63vZAwWTfhIirUWsFau0zH8RGSKtXEkxT7cYSelsAhcAQB9d+YNUeIwrr9aoLHCjrqBarO3W7ao7
N9+5E53GUMACqno1kyJlS28VH/t4lZC9Qf5lMdDvqP6wgEg1XtKVYbrD0H1NoakdvH0+qoYiYEbl
Mr/JAlXvz11s8WWNl9BLbe3B6Yi8TQy3w9gDmn0xn3wqoX9ok4VahCZZpdBME8WIahm+Z5/nxQnu
fkZnBAx8E10PsGnNt00R3yJ3sNiX99VOzm1xOMG7w2ZsNfuMtVLK9ycmYlJKzsKD3G2/wyQ2lFIW
vfSaFRstZ4eengeQtZsNvW0Gp71nCLvhSoDtKeQMk3i8ysjf5NXVQ6RNwdiDc5nS/4hbJnCma5pc
wm699OG8Qm1iZLzdhSxCWMtOoMYhxWmMQ0KzhWIWIEevnLKVAwRDwUKwwZRf1NtG83ggzJl/ZMoq
5ZdgW9sg5CyJkw6bAZM1u2fMA1QaUC5EQHxTuKa2xuUx7mz/nphewrn7oZNoDcUvPRyVvRE3N93h
vqZpTd510vjhXEXspFQnQMhdcu36RUDxg4M4T9Gud0+etRQm8h1z1iAu9FZ76ybInJ7Eck6DCe0J
pJP0+pcOGotK17SYG1ilHICRZSRFaJZSibfYi9XoO9L/4zHRIxGmA0Mg4VgIykx2l7OpXduyEQ==
`protect end_protected

