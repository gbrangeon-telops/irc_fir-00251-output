

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
HUpwfbtoJu5ljZH1PD1nirfZUiqEH4rdOJmHG3byOsiHMKK3LegkCLnxPuPlk+MO+z4ctY9AQVS+
qDXnVNabAA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
J5amwDwAOhmwY1AI7aPhS8ck8cUzk3ZbW/PSkoxcoFtS5AuFiIpCT9Eh2Lt0JzHUUKx72jQhC4xP
E8DYUPCIo40JuI++9z5fK4HwpQiCOB47OP9CCbDUXkdRdGgF4e6aIOfD40xCprloxnLZWVs0yawE
2eWpDksVPZ7exWV5yp8=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
kHeSBUaR4Gb9xyNR7/PmBoZ6gckk9p1h7+VOSSxhgJTOkeDKrcZOdIV1GDgFDrDQ7kzRgTiYYdNg
fXk4UhiKwBVyrTjV2sMzg3+WqoUQIK6Jy3j+rnKZ0FHbaJ/B0H/GfbBoAdHe7Ll2JvXvA2JrUnjB
cZCpVeHDgAOSHC+pzlRSIpPSacSQtQcR7XQ/3XaxnZYRC7uHkv276AbG3wIpLBG2zxIX3ZP+ackQ
pH7/JslwJLo+2yMp03WDL60KY4dKN4/3Cbuq0p9ZXqs2Y5D7OEUZNxyvOtt0dnCx89ZP9OSkU6+U
STforoN1MyOGgJ2YZ3QN/z5I0fk2RYpfEM9JsA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Lu2s7AKqknRcUE5f3UmM0sxhb8YGklEChkrpjNpqeFmWrHZVTV653SjxOWSucZRxKRWERgvAD5Ge
f+lfXprxLknFOXVThhIZcoGHsP1dAaIYcRFINHuR+NXvmYc17FBsIljnkMKM4grLGNoBCK5BU3oj
+OpUaEAqYZcR3Ny7rME=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ZNNygMQdh+aYmFNm+RRdz6IwBodkqsu7V9fE3BGXF5I2MBgRK6iGinaX8yLwnKR/gy2F4SnWUzqm
SM6Hy+mVD8IIS+xm7ukIVwLbM9+0zez0kJn+qWOW6DSjxPXqHRWy3fQI42FtwyVBs6pb7/W8Q9NM
y83XMjmhW9gbYNHIHq5e9D7ao/9WQ1Ytg4YhUY4H4cSzY2tHj3tbIsVO5Swzs3K1mz8KunAK9qzN
WNyQE7ctUOauX1bPhyKN8vZcKzkl7x8jPe9GO6BDBcCZS9DeY3P2LTqajNPbMa7b+rdlszJkVZWF
aXg8+G+Fp5cfd6qUK77FET8A+G+lv6qs6bNgOw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 26160)
`protect data_block
k2qjANX22zXvKLAnaU6T+bEMT81roYUMpmvcIOOl/eqAmOuPp6q7hJiev+60T+dTO2AY77+ZRieb
ap8X7asOAdfejkdaPWH/R3oiWch3pAanLXz+RHg5f+x+ADJGh67H5LPRK5Zx6oHyyBJSDRcVL32H
ei9D2I+xIeJa88PCNxmS5QMBW+c4kujEM1kv6D0NqLDQPAdmXJe9W1vv8NetVyOZAyiKaptUALiU
m5JixY9GpY5WGJ4obALpbOEYCM9xK9T+BLjaYvl7rro9UikJi5w2BB5+1yDxzk6Mm6MypkW6xHXr
u5/IHYN3yjwBeMzu1GlFplgRxOfJjDN2LwotKNxRs88BFpUfmjz2R40MTRYVYSITgdLMgWTZNL3V
bUHl99Dv3p9sAs3DR5EUPL5GrKzY4so2StZJZ8muJKf1iwsCiOEm4W1EBMj3L8ZmrzTqQxTrCPsj
6RpMGHKjer9EPj11gnhZMPyWHIr15sbAbza2gr/BcLqnoPbez3oYbP0QnK+ZiE/n9SMeUklFD4xc
P0rN77t7DK3edM1u4LZxyByvXp+Ipian4A+UwWdejmcs/YvHwehP9uRQWltJAgKwHMuKnZjTF9xG
x5dIJYtQJqSDD3xrHhweJu437ai79Qo3ZZXbzOJjK4skNl20PtXAQQb4Xsud9qLBNBkuOAisrJxz
IXiB9EzHrR1TaYsZm73RZmnWGU3SqGmYPqYCeLh5brw5ddwXrsMKx005r9o3uDU7kRAdPm/AlYqk
CDtbdnSyW/3CfPJ4I//+p/V8ImwZ5awH7LHwTTzOo0UVYy8+WtT57AbNgpnkLzd0zDcpBZN4Fz/p
D8jPrEmOtQX053unIANqJR2R/QNArIKNE8VL3Fo9Q4lWsYvlLM0agDnOBO32jd3SaDfaYzFf3Ae9
xUk/awj7s8Z2rThvH8VC2X/7hnpz8Pbf6stVdvBzfxUIJUR4QCSsggdNCYnJkGELR69fY2nTRf3J
2/kxFDGRFqfw9IJ85yzqS2SkZjSo8oYKScs7SkcsrIXnaMrz1/V8bbw+wXWB682SGCNrq8r0FjXP
qGEgLUDLTvvVJkTeLLvFMs7MS0FpHWzyhipCP7Rrtl1VTBlGWkjHwN3U76cmxRNERzEF2akuQZlQ
UNl5OJVIHCMkWYNDKZ0HmNN8Y1y1rQTXUivaDD1gg1B9UR8Sr/VSGZaD44vmWdiAaxAO1l3kekCA
NO0rlZFTcYxavsO0sIahxxx46yQ4hqSfSH7TpHd0LRs1vNZ1moXJd7K8GAQl/lib+1LCGQmxgJ5o
NYdmw5DFTznAo9eCGlXZn9pDm3QraONz9Aye9rPYYbWwEyPqsMjsNUdIuQ9Zaqt216ONPIqHpzkB
sOKskLoquae3Ppl+uW4T6czwnhs6F6b9gftxqXnpC25VCJ+gukoAlHvSOlwcf8p4HsRo0PvZklHz
ZFGflx2TzdL5MYmrjnWr0cnswHG0++ZMVGP1TvFsZNPC93XI2gEAJBUdTc92gHfdxA55xedQmeCB
h3BxRcfC9yYeYG7w5lDKNsZKC/faX0vKzOs4mpBGBreIvDUxQNspnnZ+2+++2mPJjkiLcgmX/Iwg
JLmpvk0Q92EafmB8YRuHnRya1/Ic0fuKm/+EHeKGVye3qwgsOCyOntgTwyIBXyihBylzvOwcEh1t
86/Ld/rwscwpNtq+8whb/7CIXfHsV3P86Zz9EUiLVyTDVmu5HWHu1+Dc+pIT4dGExqkryYCMkayc
PCGG6tM36Stu8qe0cVhYnYPCEzo8trAqn/nm9Kk0hL5qhHF7j5TNc+Mm5dGUy2GdpnXfbvyZfbQU
n6zP/qj96gDwQvDus7xIxVrvrmbJbD9+RrES3toK7dS/DK6KV5xqAEcxUkUdre6zaFK6X02D+eoR
w7Q81C9npNTbqQ+njiPTqPGs0KsJ5IiA/GLF4zX+pWhU+ld3+EUCjkMBZFRuTS9XqzEHPe9hICn4
r3sFqe98kHBSfJkp5BAp8I3/SM0GrQhWM86TrcBGCmAkqmOSMVSRigtCFSkkx3SdrYYustRHgujM
ch1HIpa/A4Zy2KcqZDpdCGeEh1bFqyW3A190lTXIYDfzvnsJeYFTMLGgIhBp1u5+P+USfwaQ8GnK
gGFNTYIb2e2gLiph8gnWRxJPmaGe28/dPclwcK/w1o4sgl4CZyj08UQ2NJQNx1xcH6/wI49kBFum
bMB3TtEK+k27GDUdgUvt5IT8uH7rMxruIqBtHYjjNbyI86DxvhqFM9PgYqx79rPtGJ7dn0nBNwR0
AVVf9Cimd5bDpn+ew8wkZAuolHPeTXLdfxOEbWkfCYCShLoSYsqYF7x9VMMAWyLE3mMrwRLJmfBP
YPotDHKhv2+KVwMTrejZTZW1pdTnkQYS+XXYZdgyvdCNyq9iQXyUvODdy1QPk1tvI+OffeJBrCya
xmr8Zy+blBb+burDoSxzxHey0rZ114pGyXdBTzXgpvMO9GZQaRtYXbNDenEiS6TEtMG8eiik67a9
A6U/VsODDp0hoZ5necjkMEEztwfE9FUebKjTPBmt+u9BgOatkbsCAf/QcdzDNO03zARgyUZIjL5+
0So5sJvRkaWiREvif2D1u06bh1QHB5Ghw8bYeSLr6Kg0J5ppDUZSndvjviwujr9gWiVV/DMfGhDo
RFnG6cw4ufl1nd4MKPCNVntjwz2q/LXauGXyzUUgxoThglJ0Nxj6NuEYdCr8YiLDA692QNni0nSF
5aTDMJ0BFCDtVxGgvWclnyZXXTesR3kpb+wAG6qVnHCKdxXlvu+tzk6pMrlHcFmXJF/qkKb1O/rB
r78DJ0ajUEo3E6kjRdIAGY8XcZ8vqFLdkhLMakECS5yU61n4krV/K5db5QIaPHaeJh8t3QhVONPQ
7vcsDTw3Hqs67vgwAo9oTV42mq1pPy+Wnf3oolO6fG2Px0rppsc59veUHTm3POeySRk+XHSh05K5
tykPNhI4upYe90rAYa6Lvq5e8sJuD37nG5I3Io74ZFrgdB3ybxzf1cFnu9UIHW6/sX4UHIUO0lpn
sq1Ug2c1HH1EsdoDoP5jr8noXOSCpoLzXGDAKveAy4bGjXsybsmU+rEsT6mgbB66cCxeUuwyFzZp
RSBK6YbsLAuxdP73uEn0PjdWiOiN4EWYsJc7mjC6ZQxeRGj6kTckeUj8t3NS5ZCWhBE2Ob1YRi+b
GVxIL+KOFU1ZY8uaZWHZ+WYbAi9+ZRdUTUJPtCDsjJXJZ81orAjVsZ1Li7gIoXRk2+aKfGlcnLvd
Qqbqg5TSLTOv4pwUF/EQtRWNT5U5MyZpytpqmR5ENpkcxo0db03fuDBP6DfHBA+Iw5D4JdNgtJCY
NXv7uWPdz84QXZXPVLlryq6mOkFDRPSLyDdk1hczVbcDKOEAp3Jo4XJbO9ZwSreWFRybwrxXs3GF
z5iTVdvneD/8NuHKWMQKsPrwuF1G8zCLH6fgBZRn4YuI9YGRzmD9ozqgv1NFnynQ6756+EyMiErb
FULq9LAP7ndwRisSfKXUUYGzUfjWYoOQAX6KEreQfWi1Su2hFFQWkhQXkFxsXaS7pu+rERFeJQJ9
p/SwtPdujVdygGCt9kiwZwbtR1lhqROoIngiz48jv/rK3xI5ezD01SO45vwmjCynQAcPehe6yk0H
HUL3fvoS3e961VsmIdfKS/7ARkoEDr4o4WuEuGW/bv3h7Ipa/U8ThBTNnXFtj9gjKw0hVNvpNWF9
8a8jQxbbs6JecvyaYDU22y+/bGnuGn5g+0rGiXuS9pOR5IdbeaB96ZdeQpkn2HWv68nJWYlhsyRE
ctIgJHBvPs/tFCaUY8Tkg3sr8evGYif3eG8lD6JSHFQy6era3GUqKS+hvSofcu2Qbypyv3wfsbNK
JBQvBXy2ckd96nMBxf5ICwpJ6SzDjKX+HRK7hWkDlnG8G8GI1iZhyPTnHrejO9cee6bTNufxs1Xe
RvIOX1ifo90vW7WYaYeV4uQpmuakEnoYSkAt9DOTLblx3V3mb6KE02w1Zag1As4VJ46b6p/nMyL6
KLVQl3fWMKDLvFwLN1fILuM1qkNJyTlOEfAEPKaksQ/05Dcx5LS6pq6sdwDLXOWod/I3+Yo5EQTm
tnatMyo5uMIkR0V1LUCRkCvtB5AMfSyrQlol7dMxp00uXQsVej8hFn/WHbaLIBLb0tCpHadXMRJI
dIMonOZtT3C9c+uSvWYvoR7j2rEPU1+mgKfSYRzWxPQNWwprhIHWhQXdYBQPJ7ICh9lZl8eiIJ/0
Yfxxtru2UIEFxiSIR8SV9foh4cCwjROkmmf3LAvWMXNGq/fWkv6bPkNtHSz3YVRQJF3QRfpprYk/
ZYhccc5hZO3wcsJt2LhMeaioq/vl4M/U0MRQ/i70dx5WkPIXI+6AFa6Wn8/U78szEU2p+m/GLRS5
TXccdmppC7i382/0Uj9poCKn5ZCeU2t6k0kWo5BTIL2yUiPW1WDVEeGnvbEYD4KA0zuOqStoDuOY
qkRd239ZDveEJthPhA0gc610uJ41N+im3Qkxx7+JR078TB/P9ve2vNeBABffO/i3S4hD1z7eeuMh
Qi96yNeIQOaFMfnSMKRcZaW75ACfAaW8WvcoSflAkZG2wWWZKATXxzc06rwpY/Rpthalhx8y1TRH
Apyue9T7STg4Vv2Xsl80cc9AlS4ErCCsrqn4CRkthbAYaYk8rYx4STUigFWcmHSLDVJK0sFpK0+U
DnOt8IU9uYk7SvCGV7xE7smAjAFh6x19/254ya0W3VyXOa2oGWjTGA39wjRm5H3h8ULd4ZesHjGS
xWZO75kefyQ/qv0mPze4gkpbidhGw3V6cY0Wx3jDTDgbFTwbERyFZ5M25EuMsu8rPSJR0WjWXQtA
ZvlNi7qMqkTEKyPFM7+wMg5/kt8QGs0IAyVMEH3+sY/jE8avk+Nm7Ai0Gd4qe+wUO9PZWrtMj4Np
n3Xy7Jot8RVvfX00DOoI+LXoLCvUUMxfXufrZiyPG743sW2RxgtehItn/Vs3yVMVkrOTyzasP4im
jHNfN35Lgqx7kZzAV4VG2eT7svlRAPOaY3cmir3oLJTPeXbiB+o6BlCdyVHmWqOBtFw2j8CANeaj
4insuCPlFDZ2II46J1al6RN/RnlWQuaE2T5AnFH8EKIoPSaaOBC0MRdVleKz0L7zcoM7EqkH5hWx
oNtAmXMmI3zZbEbbDMqO7fkTXnk2X//C/mXpOxvfFLti4mTMHt1Dx6tF4dK/1NEuEvNSkDDEXJaT
Ns9Jx+jaZ0aMWX8QWavFSvlZ+cS7WTqH2dZySoiAJXEsPqa5i/lIycKbW4epGssj6PAHGILaLqsC
R65uirHUYxqmhmR7Pj45j1JV1otYPbZ4l/KI7nYcwf+97MuL/8cPTpw+AaLwWA1ue0eGbUWa0+9/
RBVNkGHx1goM/NA+MZf/hucnyJLFkt6PIZV6KuJ/U+jNtaU2PzAwjTa/1HO+RHfJ64dm+q0/wWMC
FbF3WNWmEJWjslXLF1gBPhpmWVxQ8VXVE2jJ4U9mAiCAhuBsVxa+Fm0QZgc3qVHsDR3DV2RHofv+
wPJrvrMTxwtBrM9rOV50CewAWs7Fuk+LJx2edAllJoiZmTY5BVRhxCa5jv5TgawRZTCK2qEGVNRm
dr3e6Y9qyo2a8yNU2VKUnSd+1bzB1BaMs03SqMyk9CvTYP8uySE+cpkpDR/V/30i9bcT6y81KMr3
4FWMuvhgFdyBY4v+sCQjBNLbRiDJB9M2ix+fe03bHeFYUECENpAZ9qayCgnr6K16/8hNEJpiZqlg
qb8s8MHm1rRylv6PBRlDGJahisA4tT61yfyL4huoyqZRQttX+6X0XDqW3P2SqLWsX2XM3fq7Cl4T
bc9S+TaWqoK1hIfS2anEGM0PXydq1twxtoF3ZFulCupbWcN/nT/UJ4mx5otWEimMXk+qUdHUDxE4
6B4XU7cpB7rI3aU9jJrFgA4JNfbiU0p/Hx52Ad/rXtCoqAGInIkVDFTA7qn1JTUzQnfS6NSsw/Bp
62xYmiFQYX/HL4+NBtxGiamfm4E05us/e+Fkwvzh1p399IlmGYsZJWsk2o2FMAZzEK9kTcbwvupQ
g1WiYoY3rQCA0oW7RRFhVhFzaVLXMHVncO4Oo0E9m6dby42Fap1wvtlEfq5KiokXuV+FObmbnqEA
aIaFLZZZt3xVDuZ8ql2a+anwT5m5qgsCnviDrBQ5g3+CeaAgxsVm29HgrX3mScgy9aQSRv29c5ag
+d585kx2VOWuumoGnPZ+i/8WhBPbC3rQpgdYJDBilNmqka7KfdJI/mleebHJBY8ULbn4J7WY2CUA
ThBeu5o9OcVoqacDgYXDKOarq1CACjFmvg+PkYJf+n3LAdobDAXqVuJhs4rjyIei2lr9RDLj/AzV
ZdXna+7rEIEC6PqbVUjMJi1X8Zb7WeVu7kr6CBkyA7bTu1vQtyACZPAO7pTm417eywJkrZWTszCS
NYN0sqH447FpwNvh+pt4busXA5ye9q+FLTuCKzP9Kq4hYz/UO3Kt7c8IrIWxJQ42miA6W6ddEHyQ
pRs/w/JscooQiDESGKzchKMbZuf5ksJ67bsAlyHy9mQYslCGTxNM73V1w4MwVNhSBTEgO/P1KH26
dKF9xZCyOCWgAw41cB/SjMi+yY5+VYJjnN8FyJULnqAUnU024hMdtsnZ3xwCj0cCIdN2XUzfMvb7
Up1d3PVvhnBgDBpxomFQ1xDKljr4xw3Pb5gHMl0mLJGgIgSdpcrKWwdIiQcv1pKp4Y5vlhGSNeP8
i1Yc5I7AFc0dfpJM6zNiazPzcglzvui4SyG91SNAs1/eYOfRiNHxgoa+I7klHk4dQ01cKPCCPiaW
ue0BQfZzJCMm0JvsjTUNtW3aM62f65fJXghcTwPG95s8ZyR0DTZa8SgxBstGRHN1RXCgzrms5BiU
LhX28i8hD96vaPxQfJdIY5zoNNlxp4I5VjVLjhiM9Jf/87OrDZofYXMMLGpcUutYQAJvcKfl0y2M
QToDNwWqJyJxl8+epTMucbboPlWHiEUgiYiK5Mk2dv1fN6h53N2fnX4YkLp4/UAxogk781P8eeHg
RhxrCIVEPr+VJE8o6us1MZUVbIdgWffTKIroYrGakVddKAaXFFYKVB8C8sf6QN7Pa20G7iBllqgd
sUrCts0lk0CXV1iV8+Fe5crM1tZfCtY1SXLHHDaLdJlOdjkew6UtQMQXcNrGIN1+VtAFypC+ADPf
3KzVKxDrM9IuPU8fytcSlhwFnZORSdL69fieVbsEPQ5QkJZ+DrPiYAZT4Ltc3MapsHmpkUAeGfN6
otIsFGbXurIOeASVJXDQ/JbWZo+8+btEKJSmhfNqRQagulWz0G7MZAJe2fM4swgr3bFkT8r41mYW
hqa6+Cnlu+QtbQyWCddPQo2i5kA+H343p8BmiBDj5MoCZRr7DWvkz5LzuqknTLI6HIfoKEBxaM5j
NKH8auTin92cvexrIP/nNIVIcMCplXIQrwU2qKpQC/YP5PNW6rI0j4A13UPXFSWmeCmmiFoPBAAU
hS1nh9YMeXb5HkZP43aG5btTZWrXOeAlYCK+vxVUnYiKlYleIdigJW1oQBcVes7dD/P1iqncdLPi
1OTD4rVfo7CnhtJZD5zeiotTrmedqaoLUF0dUmoM1R2QmZ/mJJMXQjPJbhKUOF1O8EyMu5QBs6kU
qxiVXetv3Dar5hO2RBSktAhMGLrTqA+LZ6d+RBdsRhWJdscGT20IjEbtrTPlr5Kj18FuWSyiw2XH
6ZH1hDNFx8QmE80vQXMVMRWieafxiU0o0peA0BgBFMtmTrCfuoQ9TfQTHQh9XL5Ag7+XPhnGoIG1
f9fxeDSFDZxnqGgy9WHYwLwe/aDB7o90ROERtc0wDmLmijBKFw190oSnY3JEzna+j4MuXg47UQNc
J5Bo+96XPngcaR0JTVyTV2daeO2SpoFX7JLTFssF5wlE7HRjYPqzWaZSpEuEmonpT2wdHMxdCaat
BO6q1DC0bO8i3CXqE2WFzXpSs/gOrGio+IIH8UxygGZrdbPMTN4i3oMP9CCekSjv3ZnjHxtZttOk
8wGn1Sq/I8jqX8XwlEnyK1HUogUQJxVpP3teBY4NvMCIcEJXVaNnX+Bf62MUqXpC2/BbM9+K1Amj
unNip9b68GrRcgZ/Q/3uhisaM5re6/ti5D7jFJmSRh+mffQeZMK9AMFFNQl+nBdKHw8WXwHMez/2
bb3EtRNzemMgT4eGmjZyBkLWWFSM0jCXSEj4zuSr6GCyt5lyGaH10met+ykJMRT7WtDeJOI5LkKf
C46uOmf7quM+Y4qHDGNwuonmUoJ74fMc+2wxXM2SlU5g9jKCzAy6PIBTzGOcli+qDsGGSnLjRvX8
1DoeXjBbQ3OtADc2aXsyToEAHOwXgs9JJ5j62HtoU3M80gwVT8T714Cc/XbjHaJ+Zz0scf0c/+Gb
PU5655VwwqaQlKJtu00ZZggPo98RRQli9WdAyY+cRZ8WfJcj0pEEC8VWvQ7SV2waDIpTD4HbkE4s
zxca01Qpiba9jzg30CPnyak20geLzpGmEFBVeqp5iTtF74/ZgjHA57tImRYLmcU66FoaYWlviNjd
llMw1DI0vZo/rR6ud0rZ8owcjvY4tWwTkK/5k0Vj7yZtPdI/Bx9BB3QGJVudDsuxi7Uy0L997BV2
tXTQHpT1KYKM3SoJIAGIFCIqep4sexz5aZms9nfMNugC321QbYCOl+n9i27dmRjh4KUfRqLgCIad
FlNv1Ujk/WBHxaqI5IIDopx6DTC3pg7Bqx8Rgp5Mzg27sYR1752AL/FG/Tl7IaKa/dBtBOrVi+oo
c0CF2NnTust03UmaNv2rC9LNGDVQ1v2vZQ5u802mV/7qHOh0xkGpQ5Qmc5V4FatbHoqFulQGD7MD
goMBQ0W9A85k8wLC9IQiuyzYU9EKoz6TfA71bInIrLe/qe9KKaZPl8HaRGLF4bblvCr2jKT26piE
oaC439qLeUrkp4Cxyj5KuWPEfJvwNjmbwE7ETjX/OMG0tPWbrcYlivUpA8XpNfdbdfC4LT5NS/I6
GS0cUoXcuwX7rd+ZiIczT6bl/AQz7WREmuKY9YJwzy/OOkBBb19bcfiMdPfZEL126FVmX0TroTUg
VavaUDvInvrnSGNVg9qcMUJagCPlFAKVWixbl9G8Y3tmLFxrix3vBj7SOanYE5L/33nk/PR9UQdE
blG6Q5R0lUCpae+RY1aHG6Wi67BpbXynqcQtctPtKdlfwOW/ZpI/EwBf67ZhEnX+IW1EchOdjxN/
5dN4dJHlS6rQIUHe+EdafV8pzIPdmI1UILFJ4CUwo6/D2myPZeLZwi8Iea7GYDT4uXsW6Ywgm5ub
sOQ8FX0qhMUiVvCMoemaGgBIzV2L7vDq+OalvA8YPMOL2/I45QXxkS0RGRGbxwPsz/NtN3Iy9kpu
DAwncsv28bfmTeMFwKOXY6gTz0LR2yd5IMU6NrnsDwULjLHkFMAryO1wmQLZ014Gzy90bYZ4Gzu/
hpyugeom3LAVx2QArUq9TYxuKtVcRU/1wdrWgQussetbOdoFLixQ4g77NBbUgjwS/bnUKfAyA8g1
AuhXfxrXSPjQN+6ej9apgDVNvG9T8O5bchsxJkHDOvsXK+BBNAVZK79YVNSXfy2NXEZLEDFYMs5r
tXIYkGkPr/e2DoWP/4QF3B+4qC/Z9QSTLZCZr9mYjCh1JiUoadrOA+ywXBnA2dx8m70gZI9I6eU5
FawGsObbaOhtgi0ZFjTQvEB1eVs53Bt1RicTAD7Q8ch92ZsRzDU/rQfmVFR9m9bpzeJUaTUt0xXp
KfzCymIP5R85WV0yQCIT660T5qTLneLa9i6r2H6KJPHrIFxTuoaIrqfYEgpC6yaop8gopXOE0ARh
QxlNjoUXHhwd8afRunBGSnhU+uwES0OUIK7r+m9f4D6bFsY+VB00ojFeLxEfd2IuVAX4J5mAr0dY
yKYFeYujA7f3bdmyGWoCdi3AWcyh57naP2ywLEQQZyL83VNUF6jcZpiN+66KH3JED26btpLp8PX6
rLMiG7ecQpDCRegBBYbWVu9KEzOVIspYwRkED25fTd5TwpG9lieNx2qLkMBEZw3SXCKFQUgcPvfG
thYR/MSTzCeyvTJmN64KaogtPD06Y/QQLiVrNlWViS8qUxdY5MMbRMx8Y8g2xfSMz18vmp6YPDjX
wEIAl7JD4vUBP/83VzIcJu2ox+pcq1j84ExW7JSnJAhtwE48NVzu34THta0pdrekUSGGqEI9QNhg
DmXMKrclem85KRuIJ7t8Wp0E2Hy4LPLI7MjJiCkWFA4AuE906Uwo/5F7XI6chMPZkFdsriBJvTKD
J7FctKl++jzsNrvzDHA9rMa78w0xBDztZtgR/YVWWPcTJ6VOXLh5ofvDytwo+sqT+TaIU0LVO8SL
79d/7s1TJBuXpK1ZEzL9dhl9C0DGn3TGYle7oP0eepPArhZyNEjY8lxHv7BeVBZcaSWYYEFaPgeI
Dm9hYjPol1tGP2b17rwZsLpCCW2SLqTC2Uf2Q3U204oapuLO5qaSrUJCvLu9CbTX3vlIfox1AZN4
0lTyV2p8vrPIrZWDn/LixDsHlKzkGr4Cqzfolzc3TnnXvfZ3JUgizNYwZphh6jhkQIh1z6I95UZJ
FYU1b1QJESnboZTf4wJXCsBzMxLDi92aMVnpzHPQOAgEojzVXX9z7pWoGVjQLuxev2lfAIq3cjI8
vfC0yrbB1RewmqBN0gl1knoiypurm6LdCCI7ozEZcHAo6QTWi+6UwCA7XvBECpsEYqCQJEXU1QPG
V1tmCqBPJYsarzyqB/ScIE+c3l5ckZ79aIOMz4LfT83d9TxVgjOXOGJ4gtq4aL1YoW9X0UhIPFIr
0bADu8/oSaHBjnfXc7CWJFoIY1jowKCOgsewNjHcs4TV5bs8gfwzGRlyNUOHMXWgD9jUvbwGV11b
3YbNUgK4V3yqHSjNLjzc+g4bLRegM56BHCgbpWVXNyj5xIBz29JlwE7M0IZFwQZBeP9zNbzjE+9p
ocd+nUXiIrifWoEs8ASQKjL+jFla1dEn7vI41/GowPaTw2aLPALBNpIFCVkU7pXLcSkYzseOgBv/
fIusA63FhJ+GpFwzpUj4MhhaeJUJ7MQq0cV36t0Enm3CVOd9oVlWu9M753m/Cd4yRifG3FGWBh/h
4JwuHtzrF/SLpHKuFHmczVqcx3/V0fkGBkqFTtN6iAZj4L/rAd0DPsWq6GkIOr/zPVTCCEiFT9Y9
JmfZ8qclpLbV/WziKPVsVMVe8CSSkfDfYUeBCpcWlA3tDpQAB6glhwpnp7ICTGktsN4lvKGp4j5O
g6pz6ioU2pYvrOebXQpym6/ObfGGzB+rvfNfSZy7EcLMVcGL5Uy8FSk9NAcI6SJO1dzk8pKvufdy
nCB2uKnxaTqgRq8sRq2/Efo1oe1HZUCsudWix5LpdcX4rAkJTGwwgF7/IHuWB/IF6oHKqYoGb5K0
LqoajoaUIKFiwarab4EPqAB+P/UH94qABJgfoP6t3i5SMZF89lCgPRHMDykyCyM7mSXh9KaybVYj
aNnzB+a7RHppQN8qO0uayG6VXxLttVBaMNAjX2XN7Eir77+R1FCeSGq36IkNZV7gbQz+hXHaAL4K
SA58PyEex0umgPK/T89LokEl7NbeahtjxN7wqWIoDxpQINivvHpjqbUBeskdv7lJiW1x1Hu6/oqr
7O1BRYkZo8/R+6xnXaX3Ae2sZ7FIcWIZYYzSq3PxJ/WMVlUuysgGhuQBAoH4uoXL+bFhjX1duEzL
Iip0W6B6aqkbxhGUcZ7PDhA+0u/t4HC6q27cJHhVsr9qBiH+ozgxNLcG2EDKlfDavjmP4l6U/Nj6
PlG7K9xiyGDM+VqAlQZkuirWqOh/iLBf+Z8Pbcf/GVSxRvgxKNuv5+04P9GBqWZbDj5azdgQ7f1o
keSmWAe9UWNV5QuVMjH/eJL+dNA11DvPrWh6m9wN0wQZfX0Tq+aPLAcUOgBO3x50XgDhWk908DRn
cG431pycRF2UOw09551vss4XqWew3T4De6DlUP1qWgszQixMjSPPWv524aWzcs/ORXnUhuzfeljL
xJZ9sLvqa5Y/OA+JLu5D6UccJB350tPiUGeQxfOzPd4GMcunOcvtS5gYbjU0zf7nycl+S5jQu1kY
oFo8uTeBnxDYck6ErQgQsy0R4g0BOgQvyFxMZKVl2tkKVhCs2D1VgJkWHCvdLy8eT8Ao6aDb9+/B
66aKS2bQhXItRAuiBKzAmcXswYj2+2PzR48CMTWRqcF82rG4JZNzeZrCfPU97Pc/duUVOERBPvsF
i84v0+6CFxgOu8538ur3S0PmoE+hyuGWLU+VbaaCev2O+mahe7fql0mr8nWquBRLkZWVWQs8zaoy
rUZdKvTfFVixBXFxZ40PWqvBgpvDm83XDA3Kr2qz5zmt7Iu0zCSecseCREUjpYWM1b/R9SjvfacT
42pPM3IRjVZbZBzFzTi3sihgQsrWF2SwCVGMPRGpYiCDFb5R82A5l5N96BOXvNtseTU9nk0sjvz1
rOXUvsVPcws8lcSmoHA3cm45Wv6GO7aSAcZX6CIrTAkAP3sgzUUEhiaLLZgJHPEV61OgX+QavaGP
vzapJC/oWfTSYqV4rntAANUKncL1ZaFC5c3pUOkt99rBZaIEjzJDh7uuXghuZkR+6j+kQPF3YCbf
ctYvQGEQ2MlTOlkkKdyDBnWr8NQpf5ncW6ipsRHsU7INRF8pXEJZ+zXx0txxoOt4/7TSkmEusmhD
oVHzXOyz3PBdqcfZqyjcKAzyBr9CixrZk6c6ZuBDjA+rnOa2WB1YhrwctqeyGzfhIFn+GRxDFdHR
sbhdkrmjypNHWDh+PWJ9DOxtIKBTtzEHItYM/OHR1BAs/HP1jgkSKRtDU2qf6yeQxhdCE/aGZ7yi
y1xLrViyZsgF8CZeJYKkEi+c87SlvGkuWEbeWMBHfyuR/9SUINxQWt7u/dZd8CU79OZ0oC2WGhsR
Hw2DKjFzdLmsN5Vq8rc1VAASUxweDqjT+lzD4Je6h9l22Gy903t+RZBr72xKDhTb1gffoPitCfM1
psr1YMkx4xaV8FflFyUwVV4/uXFrHmRLRK02hdQfLZFpNLtAtxVBstStwf+NWHWByn386m2ZHknX
7At52YZqe9Gx0OSBPGnJE8FT0HX2CkLfHYhvbfghkv5/DaiYCRhgfrY9Sqdudt5qvyrAvJaFpLeG
P6tXn8P2Bn8ZP7zY5nBFzQ8ABQy91HTM9HOe/p6bj2BoFJb1JDdudjwWkjVa4oWxPmOFgOvDkT8E
Uh8ofN4LFq3S4/BVE1WeQwd6f0craMolfZW1Z0I0U13OTubdxNOGri0dW5Y5oY3rhnwpzboAjhNA
3ffZCkh60qB+XkjYcTFioHE/AFCp2wL7XUZZZKyHSvwv4JMKkHTNGEaZEDWd2a10f3E5l7dF3oo/
3yN5BZDb62wu+JDIDO+oL9LepvLMuBBxFZBqH19Y/n0HGyKsnHNeICapy+ugMVxupPmuEB9VKq1D
yF7xrkcd3+B/nIzwnr36Uy0JrUFeWGsT7YNjUyF/Ln+IokO/i7ox/JaSeM+2CpNSkSAnox1AcxtX
4rsXNLmUI1X77EYiuJc72KG9HtOc/wB9TBms/GEGDrNv9x7PUBdAUfAbLvyTzGxTsDci6dJLozPg
FQw9yFBAZqSwgs5uL9T9Fzf7wgkwnAc6JuTKt0RYSv8cXUAfoU+NmKhi9dssUd89CwbvFQxN9mc3
FeQ/mG6YeMEKS3q7zDcnWE4mvSSRTGO5qXUX3zI05lPPZMC5jfqVv6ZfSC6ay18z9V3NUKpc+lix
lP2BSN6ZUfYPLL0Oj0H5KloMkH2gPLb0QY8ps0WFS8FD57g8ORKNFaX1OVdvygjOFbPDlF1RqgK3
v84NyZLTvZCS+Sn1Az9ZaebLHpnq6fvlTBAJByoaH0PnMcWBeVaJLKqzGMYtLHO0ffJPhfdS+k7x
MaxTyXotl9HS8v0kZp66lJRNTaYxueH7Z+U0s3pzcS/+Psv05eWj4Nvi99WuXchLSemVEJbbKJX3
CXY9oyLltSlla8Qx8bPdqB8ucCFblowLGmNYXhndWDv6J0UagICsDtVgx+sh7r99Y43/LQuhYSO8
oGjKwXifVcyhr6LUYehfWnTry7vGOihBGSNSd1TAwdzeN7wZzMZ0LTZ5M8EFpZYDHOt+ErN4yxMl
neGZzdocQb6fDXBWzySD5fyG1c1s44E+wzra5C6Ff06h5rWe+M/7AYO9F9MY6KNK1sSQqaQIVykz
jWuIcxpZyVuKKGe+0j3aZvhj4zPtgsy/bEPpVwO4X9SjTuzPil2gV8n0BwRa4n+s4MoKaHLIFTdD
gEU7rOU13BrTRHrmzQywidWT02p3n71aXo+xkfpUSfFDXEUc+ecVKD2Y6vwZE0AlJngE6cXeerya
tjpihwHAfGAZqFNQntkKqvMVM8qvwaRVYi01SBYLeeS70QrEBG1/ZVRQPunDCLqOnkAoLZ0k0Bfr
FioBFeJMjsvWWVvlxwk/Fr3wLHuFMQeZjoK5ciWdtTnGzfepB2o1QhkB5OY6PQ4gYRpjE+7X0vbJ
FooiENHDNBH5WMPvKm6wrS0bAG6uC/Wb1OLbzLxU1tXQegkV30Y3PmdxhiAlMnY2E1qxWVcw9JVg
R+Az7y3UtXd+WFjF0tGYRYenlXaJSYWPuNqqjLqPe86S+U91F6kEFy5H9nsPpZCv4vURefNs93y1
r4L6kcAiOeltDzeCwqC08xwTnCbeN/vBaGpSiwaoiRVgsp1e2NzSXEpLi/NKrrRX3loKutiAU7yY
zkz0ufqe2ZPBNmKhHL83evgfffuVf6kAU/7aM8f/w/egUdVz2yU/puv6zvvgfheQPDQDYIeL+srb
T7YP6OtbnisXfRdaKdnepCKrzb6KSz6VXY8PWSRC53s7o5iAxYQyNM7Ai9NN//bTkKW3O7RTDS7b
5UJiuJFZhdewdBcr31Yq5rZ5gOLLnZJslUgNT+vCRsuat7VD3GQS9IJcggjPixOXQkpn0ANtuGkj
+3aeUIRQf3+7BNtTf6MRPefNJLMaHb1C3Q7ip3gLukekCkUsxJrxIs0rhLpTu9FsKo1wmhE2aitJ
kkzHZNBEvRG+PEvmpKbZY0iJXk9hpqWuQXpDlaJOPDYHhQa+WPUHGHTlBDUKBFjg5+gbkr/M4mto
EhSrbN1ZE9orp/KMhjzTbR8HPu4Fdrk/S7rMsf8pYvfCcmh4wqOVEF+vLIAmAi39dfEiEhxMkH5B
rnzDaSlJKb8weOwMTygxMqYLC5lBY3ERFGiEpY7/eWhEb2sxiF9rAUXEqaiFpkcLbg26NHEwkzIG
wqXV6Iw3a8CjGWFCPLTwgd1dO+N6JOK0B4wDKzCQ7KPw3t0j3iXfJbPMvgxa1b1ZVTRUr/dLJwgm
v6bNWjEhMDIRUriaCeRxrDz6+6040VdtFvNn9dTNINvqwNcOFHTcmT5SugbDJ3NYMAkrryajuZHN
8zAXMBIfR82uiL6Ota3bhg8HEHafTeJnjtzdB+Rsg1kUJeE6VFaTrpqS3OHGceg5fbu0G9QEevNJ
56hCOiT8QlNgCuvFLW7O+4TKTUlCEAaoXi7WoAsfNzV9MgneuzsIRLTmALUHvuZ2Yp8vSK5OgGCN
PsHt9PGOf3+aU0GbEVUAmLljeCjsj633UntRu7FsQ1oNzBpDDqCiYMqW/VKjKoonXbjlWymyZrnV
4CRGVrWn7WeQrAbq2GNzm3CeOq10GeRvc36YEF94ysthCdrGukrcbG8oc7q+hEjgiQvUak1tatLu
RiNymFrkhMk6ijKx4xVVSIASnLb4Jblc0p8I7W/Ea2TJwTgiyf0VFaC1OQdR4zcauqizUJtcQIAB
C76rfGUfeT54dxS9FP1tNhDlc8Qz0WiRzsOj0ZqLR7H1b6GWn9T3EGD+WL/TTdoo1zqeg+tQ1Fuz
V/Px4Kzi30x9tgWcd2xyAqUvu2hBLuzB7INj2CQSJPACMX6aQgZezpMvIj7rcWVW8OdEzZvNs7Ma
6KETRHv+X5qBdjTHQFAevpERrUDjogB+LCX0e/3hUJMiZq5ZOv17U5P2gGYBObDeemfMu1fQn8/G
dRJtPvwpwt6swoT8P1YFjItL3JhujA6yEWdYr2KrHpTLBGx3Y4O8PcoY/3Y2w2qqgpbgFJbEbAns
wDKMmX1seW+6XCPWktXDJAS0wEm7i+D1kcwqSh3h8epigDTadHEyEXixgjrhsx7tRx0PEpJq9e0x
PELU42jIQOOeoI7Q7jQHPDuDLVAmkYGIKLmpVhsg2ZcKh/65CLPpKzjjlPWb6EsQP0oZC/rQEZox
3/q81kY0brAuLyZXo0VbWjTnn+Y/CET5O0fRxRA64J5c/T14PMLEHwO/esNzfjGnZlGY82Vn1leA
RT+uQzFoDzwb2giEJPNAMmU2Bm4K702DtkGWCYYfS2KCsshHUE3Ut7M1Zd80uMtUOUkJgerM5WcG
KMfR7fp5a/ipxn1ygdAZdgHFw48Op4nNuem0S7s6zVa/J16OLz8VcMCVtBMReoUXpfLgnXBndjJz
Lvr9VK17bBrc5rLPWtKic3dt9dPcNU7qfET8quzHoHR4WaSHgcbGwUEQXNKjp1+MTE6os7r6jGNb
9V3DUj1DMNgSegTxHWCBzqmKMAyyFAml4AoBuYfDQRexMinFUoaN6s0KyU8ypoNRfSX64HSTNrbq
tpLPtn8sZvmSszWZM/Ljeg5dS/E5vLYqLxezHIBpCQFcs8JoeDRSTeJ0EWcO9BzQTtPicUzl/mlk
bYOcaclL0bG4n545G13h0UzIygqiDQMPO6fRQNl8e1TmU+899pwB/La3kV1kgFAzi/fLo7mMsfSY
xms4K4O+O2pcnlOO0jyMt4dN6OS8Mxaa13H4nPWGesIl7JbSM97BOQMyXa9SR53zBToIMLcbmRoN
IMGG3z6YlL8hiqczrl3jHsiU2L0+qIdOr7LeWXoFOEgWFdvAu4eilu3D6dDt969VQAJdowocJWw/
R0gzpJJ6yQi2JIX6cB2MriBzoDUJRg5OCnKYP/KbdVW1A8S1+FOT/1892YKaqgZni2ZNH2cRjsCy
JXN7Lrf8NIRcnyQnmCWh3s0jtyrVYNM0EczHxcc4yvqOU8A4rOHr5uSds5KsGPbk17AVKdIqQZCS
Af9/w4IIAmbAImGKRwQ5ERdeGdQdB2JwtQDn4NMGfczn2sQ3ut/s8Y2DFgfA5Jb6tXmb5bPcsPpm
EHET0Q58uxaYB9HT/3TB53ufIchLqcUII7wAZKH4r0A5iCDCGLp0twq3J3EDm7bMwHvzrdvowsV7
T1/nlruSxHx0+q4M0ImuqsLHcThKsDO9QpYRgw69FWOQxwYs7zX+L+Z+Tjl6uXjcAjF0C6d3mj+3
jMHfVoSugNXNejT6KFkWY8L/1cUNrlYY8f8XG2FD5Fi5f/6p7q3HWx1VyDyCIuR/StRM8iL6co2n
II2b1edurbtsUAK6Z/KlcCdwRPbGGndQ7IZRycnXYiRWsFh6PCLUg5MNk9wKyN798Kpx0akD6Y5y
w6B7ewz0HibnhEoqA0ZYe0PQifdAId3/R/zCO2JVGOqIRoYCck4VPKv4NGORwd3XlajdoQUCDape
JJNKJA72QwhWZOGbfCRdfIjnLa7B7I5hqjAkQcGliTGMVcawHIg0wwHlpG53VJuXXUsHzyG9pZnI
Uva3XoCMf8cOSIoSXnRBydDYcNYob6uO9WGskSTxEdR/AZ0Zte4xCnyj8KocriClWPkysxqLQ7/U
Zmp1ZBWMrkr9mhNyJ30MpjkgLszpJ2n1btNArtyZaAde5X0Jny4sGnP4yGZXlVqe8Ny82VaXQMu2
6IRTtJvDnFTxu9os8jD++p3rUMRTyO2eMG6qdvkIHYFT+sI+gvESz1IQt+ZV7tikuTinSaJbK9/j
j7wqHyurLs7tA5rqspe5USq/tSKlFlJyBqH7qdSm973BlrOlaM0AHmTHz0SJfV5+OhY1s+1KOyxR
OO1bwdTyQQG7EP+v6jJAG0hMol6Jq4h+8ST/ASB1X5ro9JaemA3ZLcjJXpGd85OIF6CRJqlDivqY
EWM88juae7GCWfMPYepuWcDGOpobv3yXFeSp8TStlxIZMUeWlBova6ETEkRyE079Bfx6noDjpOPg
mS6Gtp8ea9dUwHpdsXiqmNm8kW5nNSY0q3zTj+KYpwE+l6FgejyxdXZrfJwJWX3lCUfSAXVllXKQ
jxitxPmphNtXeogUV7fVFAKqxpyfECgvOLgZm7Gr1cwVcK331U11FoWvczJSNJJjczIkWIcduDux
mqLHqgfyRfMY8O2JDU7f+8DEd6Jk2pKrZMNY2F5nNf77P7Z+MQ1qSankpIcbS874NGwYCTQPNbyy
i8C9AMUWibctCxr/i2w7C81Y18SDT/Q2LblEZj5X6MjDzqllrLrb/QlugclQCq5ZZm8HERbSZyni
RU3S6tbxkgFqWDhXMbg9GWndk7tEJSYaKrUxFhEslnv2mtIwqJMuV7eD1lSsQJ1/ztxcl9/VonQ7
yOC6cGwWXK7hDK3xRDu+Idahj7VmvXHKTYrLBP6h03VcqLDTevgvvoYSoScOFrysk42AFvbeVzKH
HlVkCJtX4mXFtuCPfKg76wRptnyzDhcVmndnYvrvX8V9UvEHW/iF5kTyi0cK1AzWcsH6hCrSuc/+
nKOed4cR/Eq89BK2UKj6s7d7aowt+dr8knde42qj3wQEY3U8UCgDmZxKFo/s90s4mSpCdgmYQY5l
t6X2cZWvIQ8r8vz717PlEo/pset81Iop9/xR947LMZ3telhyrjB9oAihHFkkGane+osq3HeJ0klc
2ljgeJU48Xpf2hnWr4CpRnUvkWQmFcnhCyj3+cna3HdQhgZNiaZV2tUQasx6BdO4OsSY6V7SOKSK
Y8qhQYoqs61WkEi+c4t/JbFjkVF26Ul2QN1D/4wdF4+6VolUl5/Q/MgXjaH9F7VCuBYpqe3E+sQK
Y+9vSsgHC5ZVVaKMFXKI1q4MgNuYosshGK+j/vXuu0Gdr4rL3138DSHkj3t/p7nO7pEAvx/PSKRC
8Ans6eDsOyb3J1EtTeLzY9s4J4xxr9mHGRmhxAGSAWw9evtq98xEWXtxe+QaKvwCEigDQqHGspFH
vk5qogHBK2zMr3nZARkYrfz/76boNTD6biQSg7xpzTS+vUIhRkqjhuovnNMirPVpn0fxA1ON+kBb
igqKMqnoYAPgOCrq7fMjIaFnDlIyxHCOy46G0X8vVGtUgihrC80XOnXdgSWRfs9O/H7wK23OSvq3
thUfvL+5oRJ25fzIpQ5vcsxjMRsp2m16GhrOIxK4R0joe3kqF0Quv9SWwILLNUAtl+YgbxcLTRw/
A2VtmUGMM2MWiLBg9PcAHtB3qo/MlwWRn2cagez1y8lmxXH9vg2D15ISVDB65lk2INNdZe5PjJNY
HUZFw0PvH4K8Wg8hXaCpz19L28yf8n6eTk0PL8XpbUmKRuAREqcGQkzOXiYbTmObijb+VJiht84E
/jhAW11VogYyKlUgmYfPLOTML0i0jYYz8VUHrXzKvuT4Qug0JjQ0DwM5KpnFFfTUqlY68vzh43ge
IO6LJ3fNHzwPf9kKm+tJunByVQYOUa1n+cgrpemFh8qw9+TumkJmoUg2ggSaS2pojnksrHT4Ok0w
Z5HJib9LPiQO3mLXzvzbLYfbQbP5Z1du2QVxk7kYS8pKqi8X2jg2lapwp+aLf79xxYpX/o/SRgRC
nMij9J4RpETtyx1hBEFSjcCuO2ExcVud0coK1m7pma6GNoQhCa4aJ2hRhLuYqqDpScCsSrpVCbpD
MiGkKqVmHyg2Ss30/5MJxMGOYCROCNQW3V4Hz5LywSuGFerTeRGhwhsSrZ0D4cUPdMy5WTzXR40b
a3NYxA3vKVjqAPPiKYtHKWxsXd+MWMozk+s84EkL27F3/z2mxKSEk+6P8n6iQ57e+S+4mUYWxV3A
lr800cB8LWUx6PkzpWQInxz3hP9Of9GMOQCUmXU0WmF4yG1WoURQC7DspkazNe8awpKumsLWbSyC
a4ZRusWtP24VO0J3/waI/FBXSGJ8bT9qO/6QQrx8kYbieO7y+5BtSllYioDSuy3roUGYi/QjUAgD
IGItxUuUwLbw0JQuSuVyj0hG+mTvMP8TiGXg0Fv6NOmj7qwL/IkgaRZCOKGagECG2E/3Yhl+TOIe
u6SF3pTEjsh7ZDsLOoylrH9Vs5GS+ZvNfxTEbBhtL2D7oi5UcZDxkXXT/b+wO6doIZWb2Kr/i66H
8iTvY2y94JavLOnFPlB+AFvw+PiagF1XxOPpefieDUCs4clnoE7OuFxKhf5dyxv+84bN1rGu1Qoq
BGq0O6bd1c6N3CQJyzK96T2MGqFndt6NqhqfOtQbbLb1Ho0SqEbJQ5+x/dLGxiQFkhSjIDoCRu4b
VqhMDEJN7NfHCUfp69DqkaqYOdz1+0pA5Fy9++3BeA9vFj02pLpIpeFfim431i5B08Hb4IUY0vwT
pYjet31zlydCE2zvWzaDPJxdJyR6X+2ohVipCBJtJ2G2rDyT3m8WzJqBWqBO4ouuaGMIWfT+72XV
PgSyauqmENRFqvQVcXIxpP6lwMw5G9w7rSrRrFLjSkeTCL4zEffApbkoA+Nix84WCO7IQ2aZ+k+t
SjC7ChL3S70wYzApZHn4YCnKy9XLQoxjJL3XrIoMKAW+uqqJZP5uf57uhqIOLcDm27dqwL8sSNX2
y6WwJiXE41V6MrpBRw9OTmgAhKZfIokkJZ1OELV67m/3HrabMdCmsJ+P9fdv8d3sHMiSF89J5o/x
R7JBcj+GcBuRMVoMYmgzEoo+9K4QY9gDMAWoaIlwIXqIx/DMBOS8kR7INflxpy9asinzI/MJLBaU
CWbiXYdt6YosDsDMd5y6rDSHrpDIinYjkScGCql5FWzi8g88uaJtPhMxBJg2yhk6kjHPIU8+GM5E
mSwgoWDgb9SAVIF7X5ezOSwiOY9MvntvnTHAIKLqbyQ2CddkifDdY4Uspv+0qINAzaZionB/0rVc
4uGBOX0OQ5x5mdW5aYvDniUxyMbfN4nbamsAjANBp/QAubTkvrwEAtNFDTAft61N2vJIwnjFErP1
NPvgpCkIrr1VmL51zgWt5d2H0KzqP+yg+lO9GmrlgazzkJWxft+FWbqxZOmIbO/TTSC8dolRC8jo
9Mz/5mQmNIbl5lFBU6MQOSwDIDKVpz5M5A/H5oa3It1x5rqQfSG6VVJjZqkqMuyX8pBt1MESHbta
zeJvhT1BSPUfL3D2xgW/YjR4uKmq1s9VWyIfGlhw6CEDuLtpGG5yYeqo8FnRW1MgnMKFllobCI8U
Tt4m4Eel31eKh/Y4XjXXx0zzlSmuxvUpvvl2JS9rfi/G9oCnCaSAbdwMOnHtSkrcArZ57JKhaaif
6nO+ELEKJW4W0ap7+MtAsqNFdPSO789Ek6txXUiG23BHf8O2KQMsaQoqJfM1VjV35u15SRFmyu/5
3R8CeyJHvXfMYoPRe2ggnv6PXeM0H8PQuD/Jt5qG4GoVsTI4K24jFuQgjNi4Hfyl+pkY2Kl5HCMR
A+g5jeH+4VFPkKc+EnyyScrOGmDhxJbrUB/t4CW212wA3gaHrLRhCJH/ZRZsF0y+blbKc7XNAQyj
qF2B5JcQec2GBWQ1K3PbdlIVymSsKFEMk0/eDGQOmc2nO6lZeMtGHl42NWJyKCWt0+0xXd85AUdB
Y0a29hGIrEa42nKaTMypGQ+H2UJTPTj+r5UA1iLIG4kCmGOZWK18cd0cCaGENNPfT9qCjFpSLClZ
RpMp/FHOt1LKqUuo6BkL1VUUQOaJfztiBrePAGpN805ZjQxx8/cl2FPeNJ4Xn47n0zhSmVj7rTJw
pzxVONvmSmV8cCFXxzTJFjvjd5SomkX/bj2Kv1QtR0fLS2XgCoKirWa9KrehPuWbT5/7lGNKZ3/k
gtuXVfjZVDDQMXk1Ey0Cx/MG3RgBqKZswA8QqwUV/dxdAp2gSaVKPlLpfSXoX7vpsXO47i0xCpxZ
BXOSs1Dj4lCfvATbH7v1w6OGMKSl4ephu53Z6bsE6XMldL0nj/uDueeVQQopgAVtmmPxS8dKH0fl
qsDRwZCSIT9o+g1cDQbUL6kiDgffDpErkdd3a2kRtlqUKsUqnQwoGmKbQM5SBiI+tPwlD1OsAh14
ULbIqxtbZVMdD3C9LFwyyKrpf+eUWjZwZKif5Dg18XkbBLq/ugBAe9CEAPIVhflNy80eH1BzjjgU
NF9dqSuUCjsQpKkByNTWKfxUnOvSF3bm8Wd8g5PfV5rhhSNvqY+5nqtUKK52+q4Bg83ITJj/q7st
vKJzW5QqCK8wcFjYBZTqC6iZjTeVdIWmZE92A+tw7BavQo7y9aeyU1Y6aSZF8PscDhRpJnNYv+px
SSZtEk+4Qt4CfJwIuy5N/dIpvXLpimzm7+JlGxPbq8gUguGG6CftJJPhusZ1GJImfGC8hX4/d7gh
6GfzW0sre9TqUUIFC/jgZ6FgFmMSx7dpqbsYI3wOEdZtCIcXwc8eHvcwnQ7X7azpNncuJrgHWKP0
4WNE/sqaL6xhEs1OF4RKjuOPtsnftWBwV3PHzMGKvkMg2ImN8RET7IGzIQZoPetDIQ09gIkYrEwd
3M55NHMMdPtVTZRaIfDhULhMogq2fQvQDp6hhCYeXQIsjUVOLRX+m3THym++dxeIlVWDIRNDbU2X
HRS/fiR4Z0kHZ/GrwjnaNRxwm/rZlrcsVtp9avSdB1pS+iDQcUdhBt4242mC86VrZj/aknjDqWnH
qfUflpEKQ/qAieo1Mlt/7kNpsrPNUcJdgwODQVK26zZuQQYE2oEMuAJJ4T2RZasn+FUjRkmNS0rx
t7ReWs3l0xQiz4rntPC99k2WMfncBxY721ruqleCH4Mm9E4acFGvVggoFL8jqGtmjykxX8/hQkCW
w/oFbHWwUmXbRTf0GS1Wgz1fijtkYZhEBoSK4vqiGzYfl4LragDDcj065m1Gc4icKRdshii/EuG6
6P2nId8WReh552caP4QPVLaJmkoe7oqwZada1/p++LcrhVGFRXFuL5lxCBy6jGAGj6axnrztSvr5
/DyRsKxI/7PmIl0KfqI3YC1F5w7SRMSlRgvjBEWhkE2evenAPAKA1B8Mn0iewQWY2kv+5vkurT6j
Rb+f9gHyx8rXDT2jvddyduA5ZZ0PijucjhfwlN3eIn8+/XCGxxW/fIM2LX9SOuQQZI64uTzEer2+
81ngvqvs30b5B1O2nyzTaGKWc2jJ0Gik2gnMkooCP9HclMREwXCOZRjQY+jsvFSIZMuWqfmbK/dx
U07Q8BXaIMRELUqj35/nhJ0B70KwewpjQ9rMJmEpuTb4ycVlde/bzwNCZ/G7DfsWiCpGsplnVML7
Te5B6YGecrW8kxO26Bx/cZajL+MuVEkwa/wRGnHVL773EoE0AOa5qJJhkfF71rhL6v/HQxCa0mQG
1zjir5JseE3DT18Ok0GI3pzF/0qtZNQ6YN+EonNwY5VEkthXNPrjIBo2tzBU5a1L0wdTN9qhCqmj
9FBS/r/FPZwf6VltbCNjZReVGbBQyXaRaDuLcZeCEwAlC/2wr4yQuRowRLLHrV8cVvtfimOig1JC
5O7HdyWcsC/jigRuATLh5D5roXgDtLfA/IZrnrJ3jN3DxjpamVUKiFe/dV8gzMlel4NmYiuMEG1T
hAgJUJi+Yde/ysmfHK05Pmgp7Dfw2AzMtxrK3ObrPTrl0pwKNtVPfpvsKHZfmTdS/PBlYdkQGEkP
Y0Z+6Zr+WgsVjDbNn9DB8w0sXg5l9FBcKVVIEh4sz+vbH4dKPdizXbbd5ITG4OJW0g6DDYGpzt1/
AaBLt+/ZA+svELd4XcQbvH4/iLVf59gIBZumiMFq2E3kQp2mY4hXakNcK5oDmw3zy9TEkRKeOxAV
T2OV90zJCHMklENs/IdAIM7zd6btsWXMd8g611CfYznDTh5yx1XYrColU+/WePCL9kePtd2cstHp
N0JwSiBxtR7Zt+n46KLiHyz/QjjV6YXIiNBZzX3UIZZNDjE6IUwzqr0bKEq7vs64sw0REQhaZNVp
yxqqp6pgwU6B66MXGnK9N7Ywkthr0yD4xODHzkMAgzcvnr1eqQGOV0/9hvpcGGqBK7wBdPW9P0+a
7XBg7TxyHmTo+n79adIS9B28g1/JAUuY9+6knmXcfJXAeEHQ/mMcDEEQOwOb7ncnO1mF7QbSHVPX
a4MiBtqhVRaZUaXijaijyAXeH12F7VbejZDjjvLaiJMySzfCjJKkUgVUHBbCQ5JZFtuTZdlLaI8d
xWfocwe//xmjgCsYvB9QcOQ2XfBbnlX1bdlEW1nJJ+pnnh+koOznH+PwqzdtTwZ5NoJjuVi8MPjo
Rgl9uzjVzEeGLUhlEB/zoMWUa2rrHpy5SymQDR9C1OG/mumz5R0FboeG8d6osYL/Fed5/pf2TtYs
gm8AT7jwCe+gcbO+P3QwC221Q49xFog0FR1OoRRpIDLwVBOaNJjmWx2D+ho0IYlwSWpnPljFLX6M
oFdMX1RPK9TzQSSrvmlbEZNYlSu2+Vxb3xmGFSwbWAHUvtOYkCXmT4cBxpiPCwodNYhXdgCOrtVj
lV08bzHkcZbFaQDbdrYP3xvFEjknwb2wLJcPOFqu9YE0uE0R4v+ofYi4mQ34+3VV7kX3VtX+OS8a
BztmFKqLNUbDB2vke4teUxEWY+wMQuXXG0/cTGOPszEviUREgd6c/2ALHuGmjZbeqgIUWWSVlXIM
Hn9jgeTNXQtGHlid0K1ZUjDLP4mzk076etmYnJSc+Po+ARdd/XEhKQ35hUe75UkORtI+/VC+Rx1N
9T9ppWOyUWTKIbhj/kPldfxczn8QgZVjUQ3/rEFpIgDqkyfpWIygx0fcPRbWwTcFSqYkMKwOxPGe
CQGytLYdaFyW/zwa2rr75mpAfnDn8oAQ8+v6wKzXvZR/0NA6/vxXkN+Ze9msfhjBRxbZZWVzCtP+
nDh+KvYqHXzwhHGQ0eV0MpkvbsH903XEQYQmFbrvLq91/CzR/sJUMkIfPLZJrmbU/ia1C5Ux6IRF
1KMPq0Yp1pfkIQS52Vphi6qXtjOPc1M/0Hlwf1okNMBJSZxye+/7z3H6CGERjkTIlZuzrEK1eiCG
0b5e8lYkJ+R4ALt7MLseMDsaEIU8u51Jb2F1KCt2kpeyLnlzqzP6gxW/J9WgylsfhPi3ILjkHYlT
W6uawLGKZUTStiGRo5WA9vjOtHgKF8TpF7UcO749GWa+iNwud0b6dErvO9mshfSEOEMKNJQWYcii
jK9h7t+J+1PCVAhmFPZRObi/lZjVcZRKwOagIHITE0MIc+N+Rnf3SU9MmqkpP1J7bvDqOuPRI6nW
Uz8q9Y16RJW9WGEF6UYjAFyhU3ERccGJGsTa9uyC7RDb3tUPj7b1jWtjbP6PWDwbCWZIfMRZK1Kd
9wu1+3YFuL9r6tANn20YaukO0XE0oJjblLnxrhX8Rbj9blLSI4m9LZ+IB8GanuwR+B+cKg+C3SnF
NO3y1NcRNQBdcBY67Yv0GizAqFIFtw9aSQBOgNlJ5XFqVZbgMSWIkzYJ1HOOHNuahaLKbolXIw0h
hNwMf9EfzfDcaEB1/nWbjWjzHBxbvkEmvb25Xm9alMFv50/Nd7Yo5CrDSjRcfI9Apfedtn6qVrNM
/JtTngB+cbEgNxkA6TkEDWvgFQiNZgDeVO658Lobl3sQk32bTWYCW96LrFm4kpC0sR4pkQBQw+H9
WvA7sHGMF4RxHOi3TanoTF5DVXyBZUok2gyQDuJ5iZEYx1KcQNYRfV/hORgHSuPVGiOAp5dZfh0P
glZMKMgu++bGcJMUUsQ84siAnKfEHuHh2ERO51Ib9sXSMtUa5mMYbxsh+MiWmQi3NwcO5aXVMrM9
tpRWZbA8gksvxqc0ra6e53EKHi3q1JtelMPlmmYlA0pDn+36qVjsjg8tYT10hfqmp+qOMfKUYzMf
sF2+Ldd/e4xUbo9cN9tEqU09h2w43tUJM7TBvDiwQG6x39WxxabtyRyXgOqgksnAFgvuQw1dyzq7
wCgIMJuHbbuyvJHEhikd4FD7BQVeUZdGAZv+raHGAd8s5lzp27TfVxTcwfzKZNOES72mhFkDhceA
U9TZpURgX1kt0jNoMtgroMamFw92IqZI6XPeIEWhbHXH7kdab8IeKtbullgnXLyycoW/3sx1VpZ/
lFZm7Vfrg3ur2oGUumZnPKLiFAPqOY9yDOTw6wTiXw6GlIDuAbbCbP2NAd7hn8WEYR00CZMxh884
aqUHN5wLKmuCqXzOi9rJ855A3eKTTPR5Le1jeMq8yOFr0jvxObo+B7YWQVeuPZScxBfWr7UPeAbY
Cv9+EpbZQyPZYjiJe/a27cKTKbcQqa3AsLh42lL5mZ1LsV9poVCaMkGjI7achoU3V+QReMsn5uaM
DEmHZ0UHyqzn+d5/YDJ2Vk3+8s4nanWiKFPbhMCVWDppkGmAHhfGw/Ok53qI2HaGqyPEUyK5FbXY
J3pt/CurL4hiEqDJIqRAdC/xZced41M7hDaoZh+FApBr0ele3xToh7V4/VcnW6uQxJqnJ8wilw1d
JiR1sepErIp8ZAHD04LHV0L2UodzIEHRWlh63S7Dj6HmngJlkn01legUAYSsZkCESl6o1GPGLqBP
5rCDYwvmSmG98/vkK3p5bsJY4YK0rgMbUwFn5wW6gTgEzX4xhw+clwp3IlBPpBrh5KhGH0BGmS7x
bZWAZZWvz1zJLBPkQVFPhMuuL50JuoZ078+JmDDmxaKghGeKaB9u7kg+ZHSGIhpy3ldXCdBewcV2
GrHgC67IM75X3IY3Yf8q7r+COtN/n+qALJRTfEhVTh81KWMY/hZvybUvxSTcQdDJGxIp2hpTp+Sf
WyXj08qhuRki1XgNG3doNnFB7LlFYE7I1S231qs+CdcUUObVXzQ63R8WNIXIak18nMujsSAsZ38c
or/4QCimZMDIs+yoO0903Kazx4YOQ86vExXLKfM0mt3mx2hDQrPHbHulmdD/FCetgGmXbhsTddP1
hVxRa0NRDXoxsbcDwktifowVMzpp5yKXkbn4LBDa6JbRrRxJCINBQu0AM6zVVWvRomI7jO4mTpm7
PxXWqFdtkdMPFMglA/ZHwUV6JT6mH6alDYqeUzybuUsj+P0E3zN8NiKwXh0sLof+VNQGR4Dbm1RQ
7z2uADVIlcWRraQ8hZDiEOmuiumm/T+GarwP5FCvyt1/4OUfD0ReR2IzirWCZOer9Ps36hyYcWqJ
Lg9kF3zPvXk+RIUxMgmCqw5TF4I6nw1szkX0lOs5IzUa3ZHvvFXyDgDuhJuU3d/35PZ2CMZxcUzw
qpqJo39+vVfNKX85TueoQnzMNRJBWAQvdQVZon5+GLb39qBgIpIl9ekQZJZ83JTF26Gc9U4EEaWU
HT9DJTow+pX5qIRA8nBRRLO6oPs0frJMupJahbsLcz6ghBeIj/yGJFsYvMiLO0LGIsjLHT0PYuRH
BcPZaT08UXNM4TBCL88nnExyYV1VVmuB5opiyFt1Imsgi1R1ZD1PGvotpWzx4Mg4YgOhpqp48BX9
FMWexHlUdEsaG9SiEU1x/nQ0j75GRzal7lWKiY7CMh3hY1AIz+lK/rQw2FBK7jplelWmVk85Wu8y
K1ziBMjhRfbtxZFIt7qU8XOmdXJJJTSHebgv7Joxb3o65z//TQQAdTL+/F3F98shrlfPaCMOFEJE
i5+uTJMWRz/fyUqTJ4IihOiMnVQxOUPus0jn6z1g6dXMZcMIGMMCf2yHcWQvazMYoA0IPRlMxS6E
qnKQdsniyPf0FgKyuF1cNHdpf0K5EwcGxPg1HgjrMGBGhj4/fxxS/Amd/onFBl+pYX6180pBKBBT
nXwEMrsU6wg8q35fPQmfmnntsrzWL44SX+AyCSezEUNwnon8kHLWf6WcHLhxehILChomddajxRjX
dPsFducASHeOPHaFdysc1Y8HzB8kGeuyhWaHoPJmyFksxtB2wPTM+DRx8y5sN9UFfx+S/YyeDl7G
/EnfNjZW1ajcWZsbFteu+m8AIgMO/cJoEQfPdGjeijqhvpZasLBpO1fqUS4aFnOsmEl6R5uM7tAt
viPJOaDH9hrxhWUBQpSYLy6vgz9JWTp0CjQq3h71ZwWlweW1ayp5UOWgynmb11uiIZ9+UEr90pgW
xktTbkwsYFtZ23eCLv2DxAhp3oVTxRpECKSKF475oQ25FI8j9cUB6JP16ukL+7YE4cHogLY+zUDN
FE1Yt7jEvWw1m8NSxCzYcp1LEgxVOAHaKEqOFr9imuFku2UQJ+WxkXRxb8p53l2KWSJDXEPr78Rm
2p8swP4c6t2j7IIewJ4H6l7vrisH5by02A2Lo3ib+CNwLlTyLef4xPii/85zU3ALffq5DIOhMcW0
AvsiEUkWOgAyyuP4D+QYKi2sCa3vAJYG7wP3EsgRIRqOmKNEoWWNIgSnQO1oQFG+MwzRDQM7S4VH
pRq7J8KKnSWui9/kqx7lWdu38ajwSa7QwVGxcidPFukwJRz+pSqz2lqpGkthiMXadQzML6grSIEr
/47iLtDzh9Z/3vPJOHwsvmG+tpQRbYlsBQUFfx/xpobrlm+gaNKTHbvu2OKnepYU5dnU65tagMbG
rHPDInkTbS426gX1i0Qswi+RG6qXJDArTRPQDZsPsHmpQmjVQdm3WHnyis+D3vwtAsgQ3kfjxC7v
3Jw8itTKOxm5OHmPwr3urlINSLpNhwK9fqxztDNvIlzCbegFuNVnl7km3FD0eOWwzm8B5cfEYP0r
n/weukjc4i5Bj2UMEQIq/0NNGjgPnmUsiz9Zw4yOaCex8cImTKkTtHqQ/WYiH9+Megwj4pqSg36A
iQ7w6d4IWWM+a7Nt8L8mxawkMdKqN8ui3+OUlgLXu4BjVFh0yZHbfLPSY5Ur9zBlD1AKSpEn0InN
kFFlVA7lN89ZzRwrLiPHTPvcA1OqrVprT0raOJM928G9+C7VUuw5Serj+qMrkGdb+brsbZQjIwoM
1NGMLuv8JwQ+hLogFjbVjYujFOu4hGJqJu4cn8jbP/VoTSwRumOj/rWgdl9zy1CGvinhyz7/gNum
kCbLFE9jzEIQGjHOcFd0nY943oEjnj1XPOOXIYzjpZsln7ISlftaTK6XeXc1c9Pks0DGX94SlDa1
3+NRu1zXxEWkE5ECywGxV2RgQr1R82nVwMK7G47q6tHwEccGV6nS8CWPXdKTwt9nFLBhJ0dhEGTD
59/qzfwXIGIzo1PSJiBEAy0iCiOJdH8dLcpmV9+MuI+GqNVJGr0qeR2ZoOnKA+wUEy9XtHEPIlu5
fgn83zUPhqsj5GU1DjobyGKGzbbmaNVjF1xiid9NQk0jqLP+1lr092nARnqLneZNRfV8nEmE1O7l
0F0hoeh+rOyawgemo3aJCQ2i9FwQDT1QO2IcsLVtyq0MTags/hZrMoJmwZTKDUsuCn7ZsQL7Lb4e
NwYR936WxmXn2d8gw5zaerSblREsW7AOu+HLqmELtx/AO1t9PSeWOUQKdMqtPUMAfWX/UH3F07C+
/6CZvD5gx+QBDSI4lQGPoTwBnSOvKNwfM62D1sZh3fx43XJxkHulR4Ca46/5Q5J1b93JCE7Xs5CR
lkoj7IPi9Wvl+Zz5MCzNGxKD40a8rSyPNXER71t4miLtrhZ31Dohq1TVF1HN5f6yQZYb5vFrQKZK
pINQGdj+WzUqBfBLhV8ElRyIHPgaTu19DrVf6NtrWIDBzTBtvwLuaG8pbTDugGbP1xyFbjuKLsF3
GbO3ZSvhIGBbNTfFWgOPzTNB0hVxPjOH6xeBz7M6xROXPF+1iQQIF1hnj7CfS8HDnKndlXIhfMyW
PM/KI7L81q9Nq3K8aJtPHmtPa+9eQWb89XsR3gnoc53YJ9dD7NIB7B8GI+3y10wUjW5GJ0T6j6/X
ycVvqQj1C5V4rgwkixKCjJx9615PI/dD6Juq+TVsGZ7rw38kjbIdR2X2knIvlSOpKVPbV1/7lsSw
EZFmGpS3Q6MJyg3k8y4I2K8cTjBgftNKPsyBJ/x05nMfK30OR8pLfade7N/FGxYvkgx3HrEYLtxV
LvnOd5oBzD8TI8om8KUzrpsOex6T0Auv+5K3rAwZsqZPfUqgHJJ1XQJ37qtOa3q4+pcq4XfUoVkB
e6Sm9b9l+Rv2tb5XWuYlboELB2vtaYFupcMgybm4nCHoUqDziZWv1/HFs4QR+rKrpqCxAV6+cf9l
m6iQvJIFwd+p5EE+O8wFSDLnL0Z9QMgxpVGHVXmWHg8KPNp84WefNb2suwMgwU29VXZbd860wgtQ
20PGutHz1lgzXgoHMmRHdBJb9BYA4tSkw3Fa7GBJX7onSp3SQCZeFY4bnr4i4XWkflwxOLmeH/gd
MNrapPGBIubS33aW1M6nK0j2HiEmO29Ds+tpCOGoBqhcpcXtN20AfL3SLiNS5u9vSaLFnYKawDCz
3YF1nNICfpHP1825ibixkRMazJWbw1+hiuDqW+AXDR0g0LK1gMARc796REZTxTcZzBZnJYnJoFjW
TL1aL6Wmq1mmdbpTYvEn2TGjlcALUzSHo2CO7joBUyiy7czyDdPWD981z8DdHQnjCvKOmsiIKFTx
/MGYxfnXAYfch0CcTBVMAxh7yvySnFg+BmjeMXxtIXkySwJMqw8z2Q3wcpoyUP5f0bEauWmgBlDD
vwrT8HZYgwb0t0zsdV2AV1GlrWr7ih1mXpHREIQ6a9eceVdVUjI/T69yWTTxrTTu9GPJqro/Wvqu
1PHfBctiw9RMpJxzFB5HzWe1M8h3qjgZOf9VjDRH3NC3oiD8mdBZVPyqC/KAb98+8Wm9vOC2lwV6
+x41FcTUzUS6D7jNXDu0D4SiUdQW62cg8HjrDWSInNCtotQ/7FxxPB1Rj+LkBnQwQpVUsW5R4Oh3
2t1jf2KyHnwackbn3dwHdJqKSdppCLkaOodTRN+aoz8TnF+4tqAoWsvD879Dk7WxuPreKQWMiBRf
7i8DjopMZLlOY+SL3j7CWHb8EaiUemertGWAxw196LzfrjGU0KMDoqXwwOoPb8+isDjGFdoWsLQ9
q5wacEQKzHiupd7HwJvtBx+ezZnxwBfg1je4RXMgNZ4Ob3I9czLm9oBHpaIfYMBHTsiP2oM0Yzl0
P1WAgNFFjiJbJT6bx1R1MI+vfG6xFSn85DWA2UUeOqgw89oDvZ33xHrSXlfrullCKLYEQLghxHtk
b9phx5xU67KZOGJAIR2Os9tds9pHTjtpEHWYnElXFKd28ppH1Y+s5mSjUQzhTjrUA6gSjJHJLG5Y
PWJvLtBcinwfBXeHeAfhgKQzVskOAK9DdKImWqCPK9w+7u3SfPBV3yiN6FMR4xBQKIq/vqEKM9TM
k+gE6HzSIP6obXzEce2gvCHNYkuRTQrWx66Zn/pa1XQLbdhVToQYvKZVznceKBVuOradoMfLi/Ax
no8VenPQ2P0NRWiqDJ9n06u4WBE/LWM13/Ptd6WRefdBVSWEaminHoXUoiMruZPR2asBd5WNQMnx
c4/Hhd9hUnjK3duPnLOCfq0gXH/cCaQJOIQHA34u4G8a20mGISwBYVi5a3rhSMjPhlqUhQYmkY2t
3uRT0rDrR7ihauIMwspd/2j/Z5b/d6YIzMhuKb7LZtseDtBgLfuokjxcWV3/p93Iw1mBqqkxukur
AGzLPs34/VtlqH9p28xD3XxHm3xpqqXpUFJpM8ZSFWw/aLI6wRruxVTZgTu7REuWoFAPrxwh7aR9
P5ecZCVXPIK+V7/8JRhTGHerpbExmaYvmEh8YICHG4FGHpMrTQQaHGLSSMgDkSWqK/XvASbZRScQ
TiCXYbKkXH5NVMcbGmSdMxY849ftDebbaDuZ8PevD3e4fry+DebSOWaM+tsydNPV27nYRm+dIeng
dSVDo8AzLN2gIjLRqlimtDbehfsZwoUvlKL0DmIaRaQrWg9n7rGEwUO+tEDxOGafB+lUBpAof8CE
cwDVNL8vAnrDrwvAHxkXZoIs8xu0TL3s528aLNRN0RpSm1u2ddv3NbdqeNfFIP7lYFpQww6RYa7I
sai0BdTEhC1GMrNXYr2y0EGk4WiJl2l9bbaMjsnXm2Us3is1aDvf8U6L+GU92v4L05RmUiFJIQ5T
O5nNQURz4bjIEjm1Z9f/0vQkrgWWdf0T52thF/okUleIRU2uTkH6MBsx/qg8jo4FUJzts8p4UPSc
IMd/h/FZQKoaHpLnESrRObCy3aOibj/9Gwp6QKAgrlk9tg1y2z0qboJQ+m3dymnROzIGobC4iUvz
8OfNWYxI8z+2H6UBk7XxgOP5QFWaWHt8QEp2PVl9r5ZjHu0+jXUraANrtaSqvybb8+cYsTSLkM3g
H7L01pO2IXT0ycgoag/zg0jw4BqYA+5H6hF364p2S4G76WtbP0P2VxHMEmpDHMCtY/Sj7YNPzKQ2
d0ndHrpZt8SuIGlH2Oy3ddE9OSNyYdpRpQLRf+VutviWzcFPXr3sdvUO1wEk9+K+VCsFCqCH++1D
/pSfFE9HMDFbPm+f3XaIohFLNEBSe/SRNTOBo8a66Y+0Oyv0KsANcDStktzyPeV8azOVF3JPdk13
gDSZ9gSlkLWHqVjm6J4eVybznxtIWB8UuN7q932O3PuNQexHkOEZm/dzenyCAcQEbZZXWXqEQGlG
pVZPxY4A6G4C6c/NdCavDoqVHqA/L/j/ATDEl6s0l38qNuP8uRSQ+yhGLef+PxYKwBBDsj1Iz4ia
ldtnCdP2MZDLSOefs1gpHDT6g1NzrBhEd1kOd+0yHBKZ/qmpESJkjBDp/0RyNCCH33btZy33LOAi
EeaBW8A67AfFrDiC5EeFJkMkzuuCMKfTl8YrNf+ruhBqp/DeRAV6EZkQLsbD4n5wk6JF1j7KRddP
3h8JoJJvKk8tFpDQuyfe0DRydjJZHOqPiSHdM+GiZQA0nqodigW6btII1VRdWEtMSeBB/gG97z1A
yi2EK9/HOFA6Vt4R3DB1GXwcyvQdkBzOiMoK9aW/Ze86STXUk3MOgMfpnI5R/uhQC2N3lRfFUw8S
UW6dNH0BH+wZMxPNz6sbjrmUGFUVm4229ADsIFG+N9OYBMW3Gt4zBaKk1YP9LpdsUQpuJhODDKvs
9pjlx8CqTRTM97Xe2xoxiCBZwm6zig8CwF9n5tfgOcmbcVmRVwgtaujXtio0GEp07jfF2M8Dayxb
Ov1Gr8bBJRfQ1e1YQj2gvp4XgXaMy9qK1EVwRphu6uEiwaMwIqF2my3WNzJubLBxwoC2kU7YVjiE
nOtQXJ6bvkryZXbISEB/kFnLtz2Xykf1qslsDQzJynOlhbTzriUFPkm+tP3QupKZfxyCT3SJpBmr
Fw47o+iiEypXbiQv+weoo2k7R700zvbuOWmC7SkDaNWg+ou1JaZ+Q0bJ3mONhwkeAU5Bmd8geMTe
yayTCZ6GaQsOgMJ5GJmJgMr16HONBDijntbp7EBsU47NsWWtupt1J2YERD0ulDpJhJYs0yKNZXEg
tHd+3/fKbi6FYpO3NyKAPk9hBPliTUxoVNu3dOCeiKIsbbq+cnDUERpJyXL6xTqQbf2cANUqvqti
2y5KzBU5JMyB+/s8g03Wzd91p6tLVsguDNVmZAGzUa1A/DLlyXXH1zwSrpIrL+j2n8yrnI9HVO0H
drkDfxy/40zNJNmDi90CyHiFNHdeHwFKdVvrYJQw/MlqrDAdcOTInogNyr8u6EZ8B4V2DR3SMftM
M9d+AuiuznEKxymfWd7/9gggo+rTBskBtClAcSU4JiOWzelYh1g+OZh6p8toxqhK9QVDIFc1rOj/
pJqw/xsJSDB62onjf1Vb/98YIah0sc/OJo3yZUYnAGX5iV5qVvEVCRKhKObb5K4DZPg67kmCE1Ri
BClwTZmgvdlIJukBLBmj5qT72ccGhWMHiHFEE+4PFyrLuTjYpx42NkMyOHut9Jd3BBBmnhwbWg2i
73l35y1oS5CCKoSwFWsYlqtZYDBqJ2N/qYNwJxnVVrX8AWH5t7ONLrWLeD/puDug+g6SweK3vC1H
U/oBwawY32/q6uS8dvMJ+5LodUQqYMEsRESlvXJYYz9kyxVgee/Z35qoDk4/gZZ6JYx10rsOCih8
TBYW3CuSmaQuwmA2p26LUWRC+mkwMtK8fYuviBgQfpFQIDJdGeMmFtxER0zQLnL/KsEoShodnNDN
267rois5/iVhO5X97QPUZcPfpb7+rrIhqZ9vJjbi6yNEsc6N5mnTYXx2O8Lv/edkwzHBzHDI/4R8
2Ar5VfN/aCQ8fI2q+fNuJqY5GXUE0BCOHgRCDLqK5ocwlcdBu8LL7Yf5OlzxPUewvskBx9Bxz6cy
ZhNUQ8QkCVjRTxf3CX4WClaYWos910n2CYMbchj6WSOQjxMVvUF/akwK5g8cuFz6K5ktDAeES3dK
AutTPve0LgDSEISrhV3qVVdMHjNMVdh91cMnN6l28IzR6kCrnMvQa7kZDqBFOno4sPkAjW+jNl+E
vBVnIm0EiKZ+1duLHxMg7VNy+1K3zlFKtRKNtrDA0sJjvjfsxHG0uVmpFnA9tJhoeCsOkAeNYfOC
C7ea3csjxus6b9zhjlMtrrMsJ+Fh9U5kH+Qiv620Ej4J8rwUmYoHPnaLypR6pq/un9KWoMxz1HRk
12TjY+4PzYfSiYW0TcQ1+Aqif/GCWF//4L9Z1+g0R/0bH5KXKT1zxo+/22fzww4Q6ER+HfUpNPEo
kWXXsuuYpJoXbZV0HiWC6Dntex/mPvq71IyAmRRCYbOCV8A4duz+TnpXHRDAhmuaqxgKOarxMV0G
twQ97YYpa8CPMMw/q1nuUaI7uTdK+gxsjFcAcQ2P/JsgEXXMK/A/qXqdGpLZbULv4dsg6X3c
`protect end_protected

