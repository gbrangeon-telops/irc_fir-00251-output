

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
hezhI5arYh5Ll2LsYr9SKRVb8M09iAN2m4JSbciXeqmprOA6kAYKyNVYZrZl+7uJ9rCbSy2t8SS7
C18wuehlMQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
iG3qoWxeKUs22C9+IygRgNw/Ob9GNJdHtLxrQAtYdMzP86eceFi53EP4Epvud6QFqZ+YCcJAJz6X
BiP6+zFZ6SCjFFuXw9pefFKNSIH8+q7UF5dPb1d06lbHzIZD+3mRDkhnSZjrqT/zLAUZb/IQ1Lbm
Z5oVMb2d2CoW5etMngE=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
lCcH3M3hshWBn3vT8V7Ds2ckpLb00IXg/NREvwDTgQ0x1n/TYrAfJvH7lJwH3QNYGbvde2S4oTtp
dxVz5eb3NKybz4CG1wYBC2N8cyfQblBGlezgCm3PFTB/fb7+0CJP6o+JNkedc2s49uA9zPZB2axM
QOZ+WiL1UDOqHRt1CYUPiwYxRC9z2R+kY3HwbNnbrtScHXOfjyqwc/ifFZR8DvMU1CEJYRjuFvoW
cH+V2gM6YyOHMcuZuaYjA16MxseT+50plqCZJKvjkYTDhSYcuZeDAun28dPbdfRu3AO52/Kq9gTu
MLy1G+7O2B+746vqe0NC8W62Tyb+rHxVnOWRgw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
NvvNy4fG+VCfM9NYumsm2clZ8IZDrJQ3Wi+cnwU6WbSkr/joDlB0ZRXsdo0mhVbkhlHdY0OhRpkR
3RYDWBuljULA6BTyF1sag+KB46HFjV7grhZmVLUbBkCWRKYz0xq7bDcNxf7s4evpI4rWpbAGWyJ9
TlfOT5npzM2PM090g2k=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
KN7EzciqITw/PNwj48fL1Z5o1AjZa3hMKXx25N37JjIMxkR/++b3PX0LoYvLH1v4MmFRO2F2HE6o
+A9StU1NJwej2oLxLD63NMJa+VjJBFCfkNayO25s8BHSFsZkhjc8mIC5S+PHU5t+p8zDOXzJvXOx
j/qM+zNzxFnZOpagckJWraMSJbbFjRIGq2RuUI6DTykdz7949XyxajpE+pE2TrgIaNudJhMJkV8s
PmKxeai9osJTVlAQyTdS+HOwcKIcXexlGTP+JSkiagntbBuHEhDR83LTtvkaJx0GY9b8oHB0RXsI
Jp2E0CkC4MgVpkaduxkwBZ7NjlyO6dFeIGiehA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 35376)
`protect data_block
3BdnH5/pzO9bLLKq+2I/OpayvkhO9Gq2PNj+FhzM0UU9r7F4SMtjqBZv33KhElDm9hfKu+EXNHJK
eFg+fm3vkOL/UJc0fekDxlWaq9LlomTYoU+QHfuVGPqCGcTknWgKrcxgu8uQCUnhTPeZbOAekxKE
FGy9FyRJXdU1BD0V4Fp+hd+n90jOgjqNGuWfeXx9+yEfl1k/DWKdSlpiSh6q5P+xoBSIJ3YCmKuI
DsRmJIKH1XROdKEkXdSKOX2ivIi/L0NKSeApytGWfTxb0yDw6ynt0MmaMYJlF7/iarzDPAuj+Fnf
JSMgvPh/ZPxA3FA+UDDrU7P/t6fy3Utm1kJAJUFZjQ3fPScgpCQsyBNWCXjWupgqiKNX9pQ9+4f8
ybV1Yau/uIvUMBRprJX0SJuP6dbqT+0h5wnXY6I8VK8nNX8gLqJrAlL3HHGSAdYWjn2T558buZ7X
Pu7cN8f0xXTKTJPveC8b/9EcEMJocdJy2/6J54eSLGmrRxUbsQ38hoAf44ha5hfPTjZux4mnINZf
CEhYrD22ta1PkHlg1mNEWCElsYQ9NvBFEtP6LEO3FJo46/BS69YdeE5d7a8P/j9HODWHJ9q/8545
ivHWYXB86rivYopl13CISsvllMSsUGMSU2rt6sRZTEg+bKTSHqwqIpbS5ex1jjHpWnTdKx730CVf
Fi6FCfkCCYokDxdWIGs5aW7Fph6fFth9jKdPbYRKBW91DDrg8Ohh4rkiPoLS5CmZi3umpgQjDbPk
CLyjIk66lyTzgFz2MIIz0/YOgMr0rcLt8dqOnmYghiHCCu1o2PvSEq0yUm0YHGuvCvsgKK3dU/0J
FZSwacRlYC9xpK6YDx9jiDc/FfeFgtR/Yt5O2R+vNWKPBvpIKS4rmjixaQQ2UYvcypw+0//RJuuD
AtHG0tXeahu9hLpYCPOlP5SMuEuloBkn8BoNwzH0l8Rva0I1rw5roh26l4zUrbFgRWE2DCKI4aH2
zR5J9rHVr5gykx8Hr0hUkQhg5MfWEFzKjSur+/Y6Qo823T+q9Joyq+QZ05U78LPWyJ9DbKoVYqR6
3wQWRAlqZBjFRP8l9pqrxpzy8A+74ZmqwlRg/GDXZ8n79rEhzt+ybaOkS1zsa6986siCNluBQxBC
iy3VCW2rmRLzVOdLMgzraT0fPboYRXIH/kgtpgxz/pS9OdJhhVOALzzqUFeGOrlpq1DCeC+XfBjH
SlrTs3dczCGj1/lIURy+2nWnBhpeNBMN6c5UuRdxlbKgJc/fQhoUEAPE5CsQ5y8kw+hwbbNnGorE
UCMIojwcQdrswfQJgQwAJlMOr6GL0+93X5ZOressvTzTvxBIKUYZ5n+xbictwZOrSNZlPoXwlUsm
UJOsfmgTl+5MyV4TD7CaHruzlLaUdX8E8acKyrFIA+AHVln13VGFSQjae6gELhgHuzKSe6M03dbQ
MrWQV3C2UkGOXTmJjWvVA82BUJLsqex5VatossrQHdckLt20lzOvuje54o3eaHHya4pdbtI42hC0
B3+8afefT8nQkB6OjaWy4M5o27dcHUh6Z7qlDPzKZKofZVg7Zrk+LwrxepLgxZAtHqBsmmwgsEIB
zQtcfY7jAegYrPRELT4eLI2zYzmQat5f79wLQdmLiwAzzwzlZIFzlszM6CRR41/oTrqW6bE2WiN5
3evwdFMSkTGlyHHr7FLKkh8HZ1qDFtKQKQpiarsnhS6SDXtbFsOD4YJv7uewxksQPWiBQWGngbPJ
UW+eEAkrMzZ6KtZT/QZLGUU68vt6jEuLLzfJek9zMlvmncSRXcJggisF5zsd0X+pJVv7KY+1wwsK
hl5EpYJ/hCGwG98/1NEgvB5vgmtSAzlyTE4txcgMFC4R47bS2jBTcZ6pAc00GDf9ET6TZt5iReQz
EgZB5aijBoJajOm2EOMqon0V03O65VVIMWX8eY1Hy2NyCsSWPVvDSNzQAADJvVcpUy5BngWy+gXP
nn886B64ff24ZoTOwgGG3kmclU9QVE616B6QQxAEb3Iy+Nt1t139oP+n8Nfe8lBH38upmafqaNiV
JhoXVoPFMq5MZXjRcKOGYFaTJQNKUQ/AeIkEgXIw5hkHPmxH5PlX7ncNgWPxZ9g4CKVaJTGWFma9
6WuxdZmEegVWGzW+dv8RVD0bIud2fWpSA6D4935kkJ6urYjs1NB0UHBD+T/uhO5fChLTktfW1Efg
OSE5oQmZV8wjCPUIJ2y8gALBTdukeK7NpqvZr82Nk/R0eDqJa5IUbWQiQY3ZCoFZNHHf38vwMfYt
gVwvwPPESduevty4Fo7vpdg9QPredWW3SL3J2v6pH5XUVEmOs3TKdZ5PZh3xzO8es5QG5Sklhwri
WT8nTmrERdiaSXQkIOMUn/ibZTVmg/xtcLdduu4rCvZf3cHnMHE0zQgMNsvoK/tW6Sr9ljrhjTf4
vHGlzGD1h9eiiyCMsJ12itpadGNxNt5mLSg86P8nxYYPuU2BQnGWtA54MJSkDVVj/3FzD9tKyudb
W5P4NLPchBXbVZY5khJSO9l6NJyWh24uJYVWw0w6gi3Z7QPYpcXKeyHmT2YQW3+YeOSVPvf6jLZP
kVNunt3C5W4Qr59JTdEDtjMYzdpFjEcgOOCZYgVp9LHwKXfeg8X/fe7PLkf+p1dRqvpbqaqr9aeR
8k4GJ4vF4+Y4I+yGtHJ/G95iFW2qtpVS4M7tVXeClPgF2QFWB2bQotCV70rnZwc5lnip4iQ4VypK
joaerywgcT1EBUEoK2Z8asq3OT57ZpEZylB8o/gty1l1RVdz2LaoRP5yZsVJN/mLTqT0LZitZShc
R5y47xdq9LwOACQe2opRsWzlvHyE48BHbCzuh2QEZmjE9T0L7XdUdjcnm1NxwIa/qYVoUojBrkKX
Fa7n6Rl5IW9NfCnBFOFjSxYWzHmudjZGGFeliIF8NKtdTGGbB3/o7u2p6ibmTHAFSSV1Wu0RLMgv
4d7rMPX5KLiynFPE/K0nlUbodwwqWX4UpwW5gdvj/URmIHSn6VNIxJjs/1ULOAGnGRCPLJOse6tT
jhDqi6A/8TKzwZp4roBuNgwHbDR2T/7Nb0TXx67iZ2iLVDBYefExTnvWCKxy/e91QAYBKuAd2Akj
M3mpTjIbsuVL2MzdtTmxmdUoJXUlt8sfOYXiQMaDOcW0p1On8nREb8i+ecakxCxvagRcC31SjFcC
GeyoRki3+Y0ECgsHde8cEvcL4YMnthjcctaYBj+N+vu6WUe++qpZZMhTmNzDBw8THTn2Cejw8WOr
8ZDAWtSymfPkKtU+e/sXAC1r9R0lm0LdVfrIL0Qr63bMZPrNxM9IzcQvqGE7SwtAB0FhhHJrfkC4
qwLj3j8yGNDxkJBpzER5NihMTwg9SCCrS+YU9n5EV+uMKBzFC6Wyj54D+9QyGzdRo+9fQ/hS2R4e
y+ZwDAPURyjAex76rA/04+44fumFAdO5EW/5Z2SfaN7+M0GmKOz4O9up4Xkpuv8VrIUeNKfnv80u
o24yGA0BTjDQ7LBm9aJW3wX9BywH0h0IKACJ4IkQDI9+C0epsmFDdqd07afsN+8UAzsKQxLY7jxU
JegC3YKHhKtrJugYAmnlbgS6hWQByJR2v9kor2qZOvhqc03ia84p5ZtzRbeJLXo8itCOD69idiwz
okJGH0I4vxW8JEmbGlToNG3ftlWK+VoZH+GmEeuXotj7h14YE4lc/a4nm5f9SmrAE/gMlY8i8ODo
D4DLcC5Ha0CLQOrxs9Ehl5AM8rdmXcWlvy2dI/A96jEVMbPnsODuHsXIYcaAT/Fpia/loSpGhWfy
1VuTt4DkPeGh49TvFhbEkcYTmN7bVARD4kLxp+AMvNKzlTpD2crHMYjSQw5j6I/ms4bDh1Epabk5
pPFvwkEJuHMz3jCRF6C0FYjVp9Yl/mrFJmdqQMgFuctGT8bt/4NIbCL/Xv5vngr411TdZbR24uGy
KSOowj+VT84qEQJpIYqXcrjdrBK8NkCvjrz/ler+euUzFmSMA1A80pBg8LfMxgbFaPq0wy3syG9Z
zwOjutN3YCmIK+WIyarRTwYIMj/wI0ujGHEovPOVA+NG+3SIRmDjf4GY1WeIDo4nKJrxEdUBcoxJ
+OBkynb0boNrGAsWxgyBHONAyCvauiAmc+P4v2+76HK2Xal6xLTwdiclVD+qhP9CfF05CFA2C4QN
nAda7nGyYUnwlIFHlci9hcclu7VxjCnI3wy5vqsPaU4odrBQ8lAR7ZrDt+31uCJK9813r1Y93rQd
G2jutkWj3xY/wCmpMGo6rAU2jWwLj1L/iVXYg2Nm5wNlqG/mIhnX4k4cy96N4HAJpVR5vyD9jVHE
qYkh7zjzT10cnetJeyvjWb6Q9E94wRN/E8vvdZGgsycOcbSX6Kb0ZUZHR1pPD3MenOWrff8J0EbA
PUviDLiAhFZHF+yBWgXCA1RiG8g4YzREv+u1r7XAPs6s1m7mNZx9UW+gTCwYDPuMZN/OLG/X2O4V
pAKEJiJxAQrv8maEivTesZet2SjqX7mHspSzhQaevddIOF3cHnxjVLJWPUZgFPCpm9l5Zhell9NG
+Ky64ZKSQuqqgkY+RwZGIv+zZGmEiVNqgdjpsOVR77TX7Z4XIs+6gQpDGLgr2M9MN9iDCkf/aEAK
TNNhm9ZnIVm9laCXlOhrPiyNSH510dOsemB1NpI5aeRjbrJa8NmnJrrvDvb5poi8ZyHL8tKRJ5T9
GupnRQ+pr3N3918Au4wEZdCugIlIF6jrJ54INvbbIF8Obe2C+gnY7da995lGY6I+y1O9wAPDX2Py
uxCa2UTMRUU8fuCKH6dwT7WXY7Ly+LkrmRMG6xvluFXdiKd/vC3ZI9QInXx4Is4WTcM/3img/dvm
SO2s8iwBNu0HzlSxxSQNq+/+5raONfec5RN+gYpmG7Z6PRVSIzRrwuDireFQcKNggxG0sJSh9OdK
7fJMetx9vGMaaiP5xz1l2cliO6rNypQ4z2lkKZbCL5R/f+zVIAQ/gq7AYXktHZ5QgNNT1pKqeBx4
kjv7u3ljhUUpPQg8rn7MfN4kPPZLH8edv+3y+rq9YRZFd0ZY+K+t+7cKkDuFfab0iq7m7l+M3VQ4
uc6LWctDgyDCLI05gCCYU/8Esl2y2S6piAPo8jKHIu2piszFaPzWG3N6ot3QOSNoqfQ4eepColYx
21zCqfmZhrWnWDx6VHfTM0mJim9s+9/OgmpTVude6wIZRRotn6/aB7pWGfPqKCpWdY9w5uz++B0p
ufWah1TPLkGFYY9KI8oSh9v/PF0nFLbwbCdmRQy9SmItVTG3W0QHcucPM379/BOcX/FYW1zYf9a8
5/uDe+rhAPEdoobRkl5EksF4f3BsqcE1OtS+Lh+pottCnptX2DhlG1w3IaMNMFdva2+8AcYpJTbg
JORMUzybF1XGNBPUN0L8aG0G4QYLh7yRJDl22cX7KUliurJGvlMlL8vUDHc6jNcGDw4tSqXMYq2k
ri61HgIZ3fKUjjZI1gXiDjiZ+eUl03mm1QL6uSiZqh5vjHO0oKbFfiu9lXlVXhsyxTtvFPAJU/QF
wgYc7j7frlsYU8RMKhHNnyStbMuEE/uwJVqQ/b3otI3vVgQyJB0e8D1KXxKAy5cWeWJ6jZGjD0AS
3epylIDRj4UMetM5J43HlnYXhM+97nGF0DTTxbSlBINqthXbPkdPYe1QnUSnpXQiBWas/gMEQ7CK
D2KcG5oz2b4V0hXGTStjliOncaHN4m+Q68tFD5r51crYSKz2bvUldOXJmmhvE6Bh0/2CCarHwtnQ
lEP8dY2jF5nIi+3fvpZjJeYZU4mJMGxnfUd0znhOGY7WFQjXMJAyrmKH3tt7ggY6oJ4EvyR0Ie0y
hKSW+wAlAn4xgz1pzT7aDStM+V3g2b/d/I59NcLE+3MOQt4JDZOELhyXuCqzZep7NAYrGE2xF2Kp
9qkoNPyqRGNgzg1lgnOKBbK463EQB4uyXTjPaeKZi4tupeu3/Ap1+EozJZZBfGCnyKWmOjOjYDAf
QodtbB98396QemHvenl42c9BYY8qyg0LJojI2DxL1LXaoDe3vCuiOXvHhIFm0XYtkJIud3z92+3m
8kE7HOC1hwGxbLEKMIR4v4SNdfcljxu4SMhWglmpcDgnEWaHDz+oic2WEk9RYEVeMi/6vBgNXqpj
fcSXn09t9akR8crgH9rd9qU/YhwC4ulRG+2v8Qy3gn2xUSPNd5hP5M6GIw/Rdst0NWDXctCMtyeN
wUT6BV54UyjBT+7fJV3yJT8UTgGsrZv1F36le0GGkopvfPmeYGsUeDSG0eXNoXtvKNGs1b2iZptz
k7N9h43v3Ntcbq3eOu3fXefkURQL0xE+DNiJlrPjUhTNPlPE9gUyhDhj6Drn0KPL4h/5lnhtXGao
0sXcmWEGJwqcHlBVogQAXCXGmSLZXuqJ5PZ2ciKkxU9i6ybPG4/e39EkfO4jgdrxD//nioH1qX2B
ETytop1HVexqb+K770x2B7GkDg7iBFeIQK5eFSu2SBAlCGflD/tR9qlSR4q3Xv0cBLCP6iB+gX9e
sB3/bvnlf7hsimpyxDs6AiZlNuByfjpBpP4RBJ1KMD0Ff+D07j9VZZDNZs17SGTLiHsJcaxgzQOM
aXNN+8Mlgqmv05h1eEZ7qIsCs8iNXqRTUGfcyKMfax5F/BRQoB42E0bD0eFu7zIeetLuWw0o4T63
DvSCeTTTMMrvbntfATzOlZLMX1Zw+3l8TPODW6n/bzLspMbc0j2RxlZRzEtwBPAjsf47PyT/by9h
NtISA8e0y34BQdpLgvdpInphImUeGSBnfls/U23mpdM4SpbgmdnFGCxGjl9W/JztdqbM1xiWc6eC
ULfUqhbAElTDNRK3MDvY/6omnE3cE+WmZQgLa/z+BlGIKHI2TyDtaYQJIeuicilAty3MiD+QXs1h
C/xfwIvgE5oYYw0R4Scos4hXKx2NyI5yeUxx8cESVcmOT1cOkbAL0wQmonwwhrz/VXw7wZFMEeD2
FoEEBuMaa4VcK8vu+CKHC/QaBfomu10MoGPfTIokYESUefqiQIB2WG5JUnxmhUs9keGpne1R03tz
o+TkBJIl3fv5hJtgDKga8jqhm9djKMklzWvxpi0raV0psc8IOWjmPV6bvhTNEElxbiGS9ruLp0rT
8/UbyFGddMDb0AuZmVHyYz5pi6FSrW/KF15c+NJOxVrwFeFfMNjVUCtjTqEcwxm8bEgyY/cWiLDX
VnN5lzc/lObLb3BwKANMiIaMrsWMIIt9E7UJsXSxEmZfwiDm7tr/HPejApCzTVSryPi4JDlxiF+/
d7zipB2YWRR1vnE5mH4ti+D7bOMMHrxIkqAfwlCVng3NVK4syaMpELu3uDQ5/1luPh84E7Wyt7dV
WARGeU1/59cJXWIJI+gmxDJHzLx0joNbNWsnU0QA2o0JW04DOKlX0c39w/4RyFBLMF7Yy+80MNz3
y0D29RF9UkM1gzoN+ma2avoIO//VHaCfuz1pHqKY6cMlR+MiYfn/J90jV33NWFfLEnlQsZrkHEeB
G7If1DvJzwxqi08aviI1WK8uKzjv6aOfZgqjxJ1Uy/S6jLYQXKqUXc8gdmv8EWtLjuLZC/07q+H3
xVd81GxVvAHQWyO+ApSkJqd4I0e15wL+aGsUHU0PnuOXMwdIgztVrbp1+oO33BXSum0zOI3vbicx
BYO9GpxqIcZbPM5sKqaKYBjO2XvMxfO/fjzkZZT6QB/TpojlWk0sm8b8TZgwizTAeIyRV8ketZx8
h1z5F7Y/pd75I4ff+sBnRRPhKQhAlG4mKMHor+EXwJY5BFdtnWjqKwEahkMPzHa6uFo5EE1j1+f3
FubKSYBME3J1IMNzCeYfgHCL8hhDCPax/BdN73PZokT+aMoLm9rjLRmUw/QtOefrMEfC+7XjczDp
4/ZUHNEXWKLo8dNDIeAzUfjCK0ehNP1bFKNfMgWlA5pBkt83bDwoG5IGG0B9FOndOJDO9iFoVhKw
d5nCgKYLA4K+/qdGEkLpp1hA9LHDnVSqy/3P3Gi7nCzCFBsf83YxY7nu/oUgKlqeGZJ8d/2yNoWM
01nRmmsR4ehLRvrjBg2NFDzGHZmyl9EUy0ozziZ8U5cIITJMKpST1DSgKyf2iF6CLEaYPTtuG+KK
I8kt86fihsEm/hpatXFfodn27NaN6NM08f6zNI6dO/gbYdcrf+Z4kREk41V2MYrNQKE12XB1k2YL
z5LpCr/D4yqE8wHa/OJd98D9xsjiQ4IiRnliCZM32zSqwCRYL4sP4c/C5b/aHdz8wUPc9w7NAqh5
OaRoqIofJKQZM0ikbMd2056m+MZSt4leFi+SGz398mNBapbWENnAp8sV7EIjzEhq/UMnIqw4WI4P
YDzOPY35YqyBogZ2tzao0nnH7erTauQsrSlDpVpw7NtYjUTjnxsj0Ta7A4uLYRXQcKWxF68s7peP
CNQr7HmDIrY25TufCaW5uohUC0NqgEqsdK610yda2TmpZPS+cFVBRcPy4DVD8UMXIkrZUioH1fOe
vApZHkNYNXx/+pcto2jHQwZ/p1y+TlBfMW6/8r6y+lnTKSC05xcxCIr9E9G7+Vfr0UbbzCywKn/S
PWeVtnD/px0gUpPigNasnU6OmjerJf56LQ0v/KMxg98IN6r2Mxhu2nxcSq6YeExmUELrp/I8jra4
HyZXizDoWX7piz3ggBGKJXFOPG+78Mq07l79etmTCFph5SPbArNm+8XNJpUc4E7gJ1qGdNJYL2hw
mizpklCDKpc9q+6njXDWoVclpNruFRXhzWPZBK4+nsiQUVm7GzZ40+bmsHy5tg3mfwhwUgiN7xB+
udxJGD3a6+Xs4MdQzeyk5sd0vJKPB0LWsaqzDUdUhl1f/QP31dMwlciM6zf5rKoykF3stkj7LSVR
zp8cnLw50xk3vieT4nRUkpNAnweGzsGUzXPTvklLyMPTtduScdGsdG0lIfe1/7Bmlvrr9lViBYap
jEfxvJ2uVaBg39dLmzJZyjLnRW2Wl4+xgZSpbSYTZM7ig1aA8P41R5H32E/cOO8E1y4MjHvdij8d
hGLCMhPWdmAdEafJyqeDFAsE0KdN8Y/rnJ4ABTfiT4ULEWK56lEkjVLYk6ID2Xh3lbPpxPGNAgRC
FzuQXMQnLRTuT/96582BG37RAUxEQSWOK9Fi36KjBh1WdaSu+0V/K2y7EDOUgTnezLP+pINoX0FR
W+0uTuRUtYhiv03okfoKQTwdHISHPL4nm0B7LR+mdso+l0aB4ix/m/kbjQFM16vrExAmPwO9QRzQ
7UyIr/Ql1phBA248dY9TUV2/CoWRM0sQ44VedKFuwO9BCBheAmm5RtWAZD3Zsblhf+4L0vNjP2gG
GF6IcTAGj9eLSSXgJg2kNwfc6CW3ZESVV0CpILYBJAYUTyFZQWC9r/wW41F6PSMKUoy1zxhufYf6
QCzSSaoftyxENFFGdmKaYhtIVGx9I6B53Vr6zj4triOgVDZ40pb0u40xarVQFKwgeU79HZbtwsab
tXsDeg2jddw3uJ0F99f8GsWN93EYIHtm9mJ1EZcHESdJURqq6Lu1IvldOQFH7QjZ5umG+lmPIa4z
hqEzpiYt+QL5eXuZbvutnC4E3j3eZLgCNzpREVndv/vBMC9kfbojulWF7vvSojFr9YkFT3b/v7vX
+o37opa+wiLiiKCijrJ5XYpVcvyLMA+LNod0XjUTf+s0aTb0WuU0O89+cMs95Pl16W+QPKIJWZ1Q
r7BYETVRJuEjwLv4TozjKsdbb9He5mD0oCUoXO61lWarwunPELOcUzxXCZXnF/puQ8scBxJ7FkJI
ubDfM7VZrcvzdL615m7nnxuo+bwviqgNvgwXT2WpiI2GsTBg1QfPcLV826FeApLYvanIsjnYkwn8
srUT1K02mVN9fbtkk3rJVgW9y6nKeEQ/QOqdUCobEOcVHkAKgSHHQVGwKLEINrd/CsPDykVk198k
YP/GWQWmVcxIFz3GsE/vZm455qdt0FEJLq+31sCJRJqNvRGmEpD4nRQltp1/Sj/CCKSCh+NRk3qS
YmCnI0pKgNxgwS/4olTVtquycxSRvqDt8kgKWha5xxJJPtsrWy8M0KIGqZg1cveVbftQg7fy1qk2
XcxJ8LF1laiShVp0dcbXQ65Q1rjWcYwJaEHHyk7fGX5GZO09CzVK5Zl6WG7VVbhiTq6QomYwCcx5
FGLzDK/4dS63MisjsRInBa+E2kCNxLKYksNh8PAz7a6Vz3FliDIPAFhLiWXPlYl4k6NZm3GNIeND
OLlEh7ucZGXgRDnzrekdxCDv1k/BdrfTpnj5UvlGmdZihWSrKwkTt6RXKRZzmp2u7FlQUohfLVMb
VeBdXzyOjWB2mJH8BY/GXY5FHKk3BzZdhAw4Js+U6fcM0zPwd/On4XvAfkkWJNuh4UnudocFBEsA
RClkD3wXZxDp69yWJG0AUJmugjqNQoxCMkzmmaoiyL9i4b3Bg1gkW61WCHiRGD8O5L6ZViML4qwS
qIRduGk7SjUw6QTkZslb46vgjlWjjuQ90rd5DFRLbvH0Bn4ZJFw/+9wC/6pIQCojOQCHFTDD7I/7
kLb3CWHtTTjdUQ4/R6YtBRsFfuvKXQXIvhQM6qKy5X8fucgCKrxfa6KA2eG6RZfiKKRgofSpnO50
CtbbDCs6isc2dr54IbzhRMHRgWK5eX9mUzMoXRI5QaOdFabOvWqdrjQId3oRwg0AyQPxqbSalPcj
zeKDBbUnBiMCSM2+7pumhfyf4oy//8TfH6ldzkTaxo/rAt74OiiB/OreT+cdbxLbdY7+UZMgZfUk
d6l9XW2pYlY1X24cEQNbOaOvSzfHXzQIgq3tmYIiGVGQVFJyBBwrkqX46k3u24ZpKIY1+q95lnUR
qetDobBl4CxrduZV8rF4A3bFy7AjUnrOgCpILAnHs3LUQxCQI9mAQkNxCNmoE4ixBmS/sh3LyNi7
PDV+ZClrC+kvhhdSbdQRR0oG9qgZgjmyRDgsljhDdukXhDwrs75cdmk+U8gAwbJ+g30uCnjy4L+t
uMZkU6NOSFvLF/STUkoXJX/ZU/T2FXapUWbNwb3uCrfTAFDFzKn3GsZcv2QuGERSL3WtooOYaXvp
jrvoLu7AHQ/mrrPKUJaruH8ZWlPtYqHdI4I6mKio9w1pZcqWkr8bBEZQhTI4OZtCZ4QcR5gs54+H
tK3WbfqqYMdo5o+ubAFq41HlT8y41JNIpXOtMs1iU4NYs/9nOreDEHyKENLM3BNavkdMIiV8gZQ+
yvyrN4ttNo8TRqu3l4b6TgUTGKK9Q11gXmmmfTyrgUq5N8p/Fb62wxi41psCcfXsC4rjyBLgZEFi
qqUisdA+Ij0kWFnmb5XMS7Qje/73EzoQvMda3dRj4ueq/syswJXDdlUJQGH4FovVnL67E3NlWdwN
hy53dXASqJXzrEOSM0ZnhIin3od2TgH9ZGQ7ogCgeJ8pmc2Atr/9lay/kCCiVPB8z3RTDHiZXTsY
wKiGfaHDrCTYADd/+8zFJAH3sHnilkQ6qmcHliHhVWvhISRFz+2A0z/2CEV2TxXEak0z4IU1qiXL
1EYK0+FVFGccbutpOlia+KSMOYyBLVb16R+WdIKX0tvcqik0Kw8ZrawA6J2BPvLzN/VK24YB8SAC
yV8pdCS1wYuKn+ACyHyGzdQhoDIsEdAiB1HES2xeyrAjIcVVAb/Ip/9fTO9A7BmeKnR4g6oupe8p
atkiFpGUPBnYt4jxlVHIZAFVfNuXCdWghHXF14mVtpb421mILREU4X4tDtk4DgNQvT5UE/y2j54d
oiqIBAo1nI3+ZSdV63crMPj5TiFc9XBN5sx7nAITyORDoJTMXDOBOAM/VyWEFOJherDM8wEqtg/F
Um/LRpmil212I113VHSh1rqllEpTa7HhCx4nvj/NQ+B6cQP1x6N9uddJ/OT5LAYEBCfJvNn+c/aL
hIX2JKcvrQ1OPLV/yhhhTutWD1afHoy1+TDWWg3pRp9gjkLpDmWBabrcqY8W6XodXlwWVmcwIngt
rKI/qvnqT54ZBW4JWlSXJ0IxdsY4qvi5M1rFbihzXK82ld298DDIG4KT0OL2DByPmFgpNKRw8H3G
vUqMkw1t5/5+kXXGmX0eeI1JOXRyGVV0TFdp2vJVbUK/+rOhgycFKyCBZrRB74IXFcCJ4bR1SVMb
dwvqGB6yaei2M7Xv+OcqliHJOeBbPc7+t/Tl3ula50VJD20FS4xq5ykhKztHoy/M3OztRsXDQFf6
68xMsGYwDGKIRwMWVwSGLfaHLLP5ftxRuVEiQid/h/uqNtPG4Nt8MWctuZrQEHuI4b8u0BjbPWeb
iVALU89UDbbhWfzhjktHRrVyfjL0bMGnjShkh5YKG4qWqI6dJJ5PgBPwlsgUNdMn36id0ijMKnF2
0Y0nfr6EmUmRiA6PZFZMSB7kgBmTvmNT+vghZAXbztDcqpLqLsdoOycdBTloakeJ1ZCBfJagfX5f
R7kSDPuWj05bEBoX83d8VTAQydnd7OicFAV2l3DMcOX9Z63P0Qi5eEHGP0tGJ9bEoiIR+Z4kF7QT
2DyiBQThImCrSTsBIVyDByvHFz9n+KILZqQsqNXrZ6JyllhDVlwKI7jtvzujG8I1Too+HT0kIx6+
uW+gHvItzTt6S6HkQUDQuNBKurSHZivLIv+qfyxIyUBLSzkkoobzrgkuRRkfOa1m28GH/e6ZhCle
to9vM3ETciZb/gz8dbAlciUAh/0QSu2+UY1LWTqrHeYVBdk9F3dVxepdcdWAqyL3M5+1XAyiqtHg
9mrqDjtUjm3+bFba/f+PKHcmiupV88rCg6mJXTKohwEYYUaVcuAVNJh3SLNX5HginsW5hnMO3Jip
g74Qcgb4k67s5cvzeJB8npZ/NXQNAnpRSiCU4hW2FcdppUSrt3JOsLOU4NtRJmJDW/mTl1KuqR/e
PrX5JAsynj3yq8dKzyrY6QSVxrakAO/u5mAUu4cWAv/47Lv6FTH8IpzkjgTdfy2goDMUCdGpup54
zRoRuQnXVU0c1ZLBO1pzrt5E3/PRobPk2vZPLOOSP92ZJj1tayzqpf15NVErDsPqggsEf6v99PHq
THWSADGaMQZSJ31V3U+h6FpydN6p6Md7hoTKo2bPC6pLC1L1wON/zTHJMmGsgBochzX1y/fspeZU
lxUz02Ty3ChtqXTukC8/kU4/Uhc6ruqpN4bPGrQPs94ZhpufHiQc0x2AQP+XLFK70mXxGe+DAhkS
b5ONBmnQLb42FZysHsBPt3I/LRVVg16bylq8ZjE8aPTW+4oj5UH7JF9n0MfIbGli6LWNn5cM/5OU
4XX0Ai9F2IK8RhhusbtCXUEjFFRK78qnPDZuknbesyRdH0dbE9cxiwmatHAT265dTrHsk0JixV9P
iC8uwn8adRhvPumLxU9vZ5sjawm+MmNA4Eh+1Qe5kXzIX42Tu2iQ19amV4t5f//Sub3fJxGclWgM
tiQEs1xCokA5XqvGx76w4scSRVB/98f7SMw0omLit5K6WW4hsZ2BwdWHo2wg225tXUr3MNNxrI69
EO1ZyfOgNvButhSsw7KQYIIhIQ2anCh9c3YbwOMabpw/RSSc3UK3VG8NhQ/WvZrwfJ1S0T+qMWPg
BthQws+P4wCYJ0Bw4L+/rqffsuRUH+4GtbVJ0moMaHxAc/4i1RGgJSDmPL1nfqLYhf+UF90stS4j
mdbXMtdDwhSZqP+HvuHtj0JsiCTuVGMlhc67ZQNO96UfaspltQlK7LrXOz6jhOhIxosKuPUOwwHb
K5ER7KOTQrCvJROe9Ny3avF5xFL5G8exO5y2Bd8WPyd/eA6EzAJNNDGvR5Y4VStmaad816d5vstO
76UWCmr717xscvrMJOwUfQppHrEFLYvaDdAcppYBMuE4s8BApvBBev9BXCzHtGG5OXDL2WgDx7u9
V2HdYoWuLl7Aa1XJA/kPJYbTyyS0a/peper7MsTs1RqXWQeQ22ZXyuffNJqQNTXnCNFYUtLTp9p1
WjJYw+Z1/gPrvQH6yti8GkBKn+8ijPaM0cwwWa1tMQ9RWn1D+34pw2KmLBeoOeVV4jMaTPAkCkLq
DDR5NWcXAYkbM8fTc2hHIe3J84aOeB5MsGUyvTunKSgYMn1GEonpKHg8c8uH5bYr7V+xpcxSO4DL
mBnhJXfte5hT292Pa/iHLeM933KJqeKqf5EFjuS56aEN5m1CbuYqxKDW4MHkLgiHMAjbTDx+UrCt
wIXWzJ3iOvoAQPLiAVx7p6nuQDTdC29sHrgv/8Q9VhvLlE24wneEFXm2+poH6K/PDr1N25xnC5W7
zrsTHWv94KruWqm9qyL5Dlzk56i47ZoLq4FHa51iJiXjjFGMHpLCm1zg0WLDFcU5KQkyP4wizsN/
y9D+BKKh/wRthAs4CBKxF2YpN02ximrh5L/1snMMFN190TSpvE6QJ8Xm4k/1Ag7qcOOZza3KAYP8
zoDNPUseebMrv/2QnvYY6E2KNIIkqr6kWXz77BCujzJQf1RX9AxvEQfw1UvvksqU+y+C7AO6pp5k
ZnVkJx8lD3w+V1mmyWcQ2YoF4eD8HmoussiQ/PWDAaOBXQCDaKbeuwflBrgFrCQb96+H4HaE8dqH
4pFJxPqwYKsLZIkrgzbKb5VJgtzbAKOpipiBFdWTI15xDqYd0dz88P0lIYoGHEPl7MXz2HBO7Oa2
b7UzJ1za38p24RcqpNRnDiIO1pTfclq7WwT1GR8hryfzZmMzxhlSIs9VcVr1IPqLj4ktoG1teA3F
Ox5DxptT5clyG4jbtsPD+zdjKjrrOac3pFxDQnj+M28iAjt/QW8HrcAoPpIXpB6PXOHI8Nn+pudB
OLFh5OhXSJYTNEGHJWl46skVg0qzD8KPS22pWwJp7lYikLbOvHB8PaedLzLjUV9G8kZDS0wuRIeu
c9Y/3qK/RD718OXxQbq0NOOJ6pzseYPXrU+Z6xSFUiolcfzpmyCmHe12VZzc6/A9K1FPRm794Me8
32zvX6aDjuCt+IoETboqe6h9MkLSCpIJ5KxaI7q/5+8ZsYS1QeADiA45dKfHsH+vnZaBQORhIJjj
62LqIzGp39DMH6JmztUlW84eBNM+QsrGkcCTyqZY1KFi/mRLgoNheYsM8Cp5gGNExWITjiTGl3Ii
Nq/gQLOYXvkAG+FuuctXcA7zNHLR4g99xaszqQs6CxjSiihSfve53ET7jv/4yXoibX22f47jd9j8
U8ZYnqoAVDDBX8pB2fV4AGH1uuqzuqzg661jl5luUdrtJ+iARWUsOghj4r8mJ2wsd5nSiEjM30xu
RJfnAONS9tfG+kbultVLVcCJ1cLBpTRdnhEFBhY3woU1G1sDM0nqHtHImieIOzuhq9HzxsC0W4le
JwmQoS6/PHwC+zYGhm1ZI/N16KRg5a9HN3QRBOgTxLhrceoj8nf0dhCXEpeliMRD6BfVb/QfReEC
caGOns9KYbRdkq01ThCxO807yU3Cwo1rAfBXerXm4XLkkJI6q99F2zRwwQXNallwLUJd4EEhlARP
vUHOqBBwGr8F5k32NRHiZWG+EaxSsVEfzP3K5/POo8VHHg8XqRKrdSfEKqCS2SI/oTFDhReibgj6
AuZArLmSP4IX1XOYU6B73+p6TaTIj6xYBuE8AtWArUExRQOZCMf6Dez2jfdH+N5gXDWa4hOVX177
UlDDLh3Ggu247oRQ7lE/TG8O09UguLJRtJwVS6jEt9hmAdn0+F3mYPL94JbiX3+2MoqVm3UwQRxe
bTwVudhvF8+7J+yxHn7iRSi/PZ8GtfMG1KkxOHBbJXyMIjG7TUyClRhPIXyyvAF+upzrYItWrXdy
7DjtxQMBIsmIj265sstc62yoFbJWNM3OgRteEvt/WCnHbmVU5nGzGJxRyxJhdi5pS3TMyu2zYJzm
k4+bLnEZveoPunVMEmMfM/I9cuRWEn84nv6d7kcOlNEUj371PpoykAdHesU7AYh8HNSrgE5FD14e
fJJF/+JQ8FQoD0xt+qtDTPBpr/l2jlzoH91EfKl8OqkH8NgmqMT+A77IIzU7cHQB2w8Efmh1PC9Y
MBN5JRmPsJz0FCp324iReX0whg15j9sor71dTEqp+wMHDvCpX66PBaNU+eoKWiTDKG2ZermYb+G7
ePAxELXGcM2r/4mR5BY4M8GIjM0R/S/V8uYf3SpkRA3DttYyV70sN1eTVJRjfhY6sQQ2bpaGiKeN
xxkAk+tZJcrOBHMlqdzD/j9o5C6U5XljBlbPU4IVXI27O+sqDUKuMskmXKSCpJ/NYGjUvSmhUN7k
Mr7/+meCP6jb5LOfN43o7FLj2/qxgws4X3AdgBglOQo/8GkBQekorvNyUhi20do2PQuLB8zpophv
k1LfZPPw1CArRJl+6DJIO44AFsv5ekUPwX65dlKm2wI6ssRViESeokViIcbXEHKb+a7Ev3swVnWw
/mfKqqKFmE2E55MLaT9G2YdOP30LlSjSP43EdWdykfIKvdddO6CSul1sWYokpNrDp74dnxsZqo3p
iRrNQTBDxLosBrLTvho+tzLeRNJV5aXcuUjcLQrwCxTTE2Oci9/mG9DlUlqG9jPVPOG5NmHnevHg
pbEU4i4Fp2M2lmlXBTI3wQFifq4s5DzDNKRqEEuo0TBSch9mzUgrprLRMfDSePbDiMlavDGGs+Gt
m2Uy3jjwmJO2Ku+VdtYdIspo45RVP+sQdePl37XqgrREJ8fk77A5HNxJ8l3zR3xxY9Hed7gvXZFF
5PpX1CEePxzijkMiC2zANbm+7eq8IyrtN6MCQDSGqAeW+xCh+71PUn4XRNLrC0XeSAX5tc10BcWf
l4J4TGtSjtKuMaoNQFVVQML83YXKL7cC9caN2LFxpQ3Jsmby0i7FZhLqE878Rx35xIdje/262dFO
wyNWd8bWZmB/N+fM82kHgWsQltrxwGj+bVaTUC/CadGjXqLIv0wnLsdZsInX8mHXbdwXsIUQPBRG
M8gsdPq/ZA3jDqKKEGL82YivGcNAmUbBks2RVxl1KYpO3xATLcnc1caKeq/cuCCNMBhhRaVNfBJX
1y6tee+jd86wBe11XPnJKEfDIuQaxjS/T8C6ENik0/z6EHrlrPGSB0PhbIj8WkDWh5j7t1j52jDt
Uhg0Qiuj3tGnwqVhMl7OdpFtBqEaVEZmxTV/okm53GYw0rb5q9HCegO3/X2P3fWWl4pAqS/oEoDC
OpVf6XcDhfLgyecGygsfxv9RIY9VRFLhu4bMpvDb5fvn/n2urWrxq7tHO+ao2TrAvCFKUsuQoHgi
LfXy7khk2gvZT7NL+vY10PcGaBagdIUjr1geB5l7S7U8byQlhjDFtvEbF7OswRsTBitnPqH7EoS8
yc7/uv37hGyVlybFs8RJB96ppHz+ZWUngz4nSkDgCy6JtQWhH+w+vauRyf+jzDvMqfz1dtGFNHMa
qwK0XMWEahtvepBFSJrQsjNzQsu2n5DfG7N/ODC/qoe/2olznXgxRatTJwxGHQgGX57ts/rU8EO3
T8RLH/v5piWZ6asz/Y6rbsuX9Fex9jgb6sPBf/fNDQHzZuxcedKTE8kzhk+kGjIHNvV28ZWBeZUn
lmObJN/yW0jRru6FQUxr5llASuLpsuLZyf5cRDGZn1uPjEQwPZvDNttH2QauvAj2TCApHpr/Xr7V
YfkNsbU2rPBy7mAH9jVtgFk/kNk6RUnjDtveWDSg35IWUNVGwhgxXCKivTgnp3PhRiJujJYB1qy6
1vrWb6fcZWIRLFp+d1lWygzb6egDNJKADVR8MeSM6OpumoxSfUWY3p3kTroO+6lirU7c+K5UPsNt
XH8AMzHQ8BeZiXs1408ikpKo+DUY+R16desWi9tiq1wafEjk6yc2zdHL0TSnLG/L/nckSqLrfg5k
mkr29au11ga+C9H66GCFW8GWuxqpyQ2xysNDgIFZ7iWQAQAHWpObEOm9jH3d8qeT7BlJWWsmYkra
Lszu1fXgOtkJNK/IxlEhyHs4wp/W0Dk8l0zpEN13A2IiQWb4FxTjV9/WFbrD6Gkzv8UbDL+Ibrms
4utJdkf1KsafigEAKnzCh9YsPmCvDIiHWNLDzfAcDR78stz+v4beT62O2ZHbqJ0XHPs6jA4Sj0dR
OLtHNTPgzx2cFDLIRddnhRqG/oUwlkImxgs+yVZdeCKIMkoA7MUcn3uyhFZ0bb/a7vjAdhiaP8GQ
bavhYIIIw/aCiUqZsOya+TKmeNnkBLnH17MZjMfNsUpCFJwHjlu70KhPl4GWLhSoCunLw+rYlUR9
7dQl927yf8lzxgsxhqGlQbpaFxjOq/rppN8dTkcJw+uO+aTN6As+FDYB+d8A5+GqJ9JJDKk1pKtE
iKQiOUS8TaGlgyXU1JpqIoqHnV29TA6Ssh+LQ8uQBON1XylVKN1dAgOi+sabEFFUWVAWWLo1zU3D
XxdmkU2pZcFK/GPNaY/YqiWyxy5gTX3FmxHTN+VgNUq/l19daweAcLGos/Yvd4W8Vjb5I5ZnecaC
VHj/uP+YIjZe5qhfvgqUXyUzNUxNnbKuUi6xkIjJ7P+gFYAnsfp83c1EWFMuMkPIdOR0770V33nL
+N1prCTDaqBvGCm4ZdRh6SpZodPHobF99O14e50+jchYa7xPwZYfaPqNkmE+kp0Ef3byPwP03KCb
9xYUhIeZr08jxM60FvMt7MqEMqkD1fYU6jylqvT7ue8yiJ2NCQY18cHs89hMruZpM6BDa7MQHGFY
xnSA2FCntK0KF1VYBm4cg4YxW4jnqa5ensT7gEqvj6cC4qLOA9DkEHyMmMzPItqaLsbo60PbLjRT
8Zi4ZywweTcliAGqb+ezYbHsdntep5XW81w72IcihAdyFMJD3K8RVRv03wV+uVn6T+ulCOsxGq4O
5yoyS/V0+H7BXVmCRC8sQjPY9hg8Wi7yXGyXDJyA0UexDpqGyUacT6GtC7us3funMoqw2b28vInT
7hfdwIlPddcYvUHs2MF2GnNDvbWaGLXcxSpmuyo4fRfqhCXe/Qp5xvilgm4ZELoqU8JqVZmBAQO5
9gQZvNP3tucK4ouumLN2fFKcCinqo62I/DJNQJdVeE8TGj20hrVJ9IswqIPxNxdB8IiMj+Tpcat3
pzapy1Za0StKHXmCzqINbCSf5VlEDg9ShJsymcsoYEe2Tdvb7ikj8P7m+flMTdWFOGqwTgesWLk9
bSz1SKkyYFm7WubzK/ZzMByLeABu7RSnRKg9mDtqfZQ9HUqE5cvz6d2XR5mDpqoz1yj3nZ/bPiY3
7qYESfNdgWwaS70zF39Fn8ahcRK3zzc0Q6L4EmL/iaTJyF7giWYzbsg9YjCa2VY6Bp9hfj/5Vysa
ltdlt6qZ0gzAcFUqKoutBWbOGGknr4R3b02ZzmhUxUiEHZRV2peWg2YJoJ9I89VPafQ6cr4Dzijz
7a+X/ThMsG6xsL6jNvUb3UxiESe1K+XM8LIjg8CUnVSd6O/GFa3McWYDnZXkFQmDWSfH0KHOSPyb
kcyV8FF53d3G6szz1B7ihn3e8IBk9pEDtoL5QQ5QoJARXMUlCpkpEvN786zHZLOgEGyDpyAC7KMC
kDBgXzeKjqF9sTE41ZNQR+g4YULmaeK1jRGOXKy53BlMF7hQb6Xooe7IN9ETqA5oOhd8sbqeduDr
H0QcBb5r+SqoIdW13HOcAJRZHMoSa+Ehgrv9q4MZ9Z44t+KoIlrVkY25kyMeeBionJbg++r3Q4Pr
bhLzRbnIYBDLSRKsqdUNQsPPSeCyqIrIdYUqGmWgADxsBqyNU62zUll29z9xxYNVAY0AAu5ZDB6H
kdzAiWAzLkeRAjih1QyLL2C3GSR6PGLlxZqpgJjdqeNEdeIyKLZKcMFFlC/lNSfYNJZjbvz+MkqE
vy0YPAB8/SP1Y5l3cwoa5HA5MbOVSizadu7lVgSYATtrxxMRJ0+sR3/9541eam5I982q5d7pQZ/A
lEXwFUarqLMHNTQjd/To9gE8ewvcA4EfSQaDgvJXR0+juqOqgy2Vrmf+EHUwHzWHPwoxqfXAFdXP
ocGkz/T+MKvgC8dKPw7puJf/55S6tbZohvfK+UWcSSDI14LNi6AD0sFUdCaiO58MzJqd/qj/ZpmB
ZMCk+az868ATGJhuSxtoFPuxvbVQgA1RHPBUCXhzxZfivylEUzeda+lZGHhsD2vK/kAbu6T+koY1
5BDmidJg0hxyVZg6qYVsIZIDzfEVqUaoTtUbA8TFO2pSZpnzYBsBlFxrjqUgxSS9w5VGyT0kOEBz
K7fPq39iF0w0UgPaa331hO0ZFgw0Xg7UqCurHFtX2kIP6qkgH9pR7O6+59iWlPKb0fCOWGxE943G
sqYryyyQoETo5AEv1GxAy8ws7Xx8af5afACfIFFussRq/NyMipXasFJkYivlqQGQgA8SxI+AW9Zv
/POFaYz584vIdyYo+VRcyV8Y3BJF7AX1KIpCmSVgtYzr2an7fuMjkpWcR/twoZYG8HDOA4C3G7RE
s4S8GlLTgiUQS7IzOhEo60LJLeVECbjBT0uDn9J71cgSUEK//PhmQFovufRcO8LZx+fqOs3V7n0f
kddeuEsK82eNKhexQVeFCC7PW90qIYVHZQDUKVkblH6yjXf4ISq6SeNOQKeWQvYB2Qs5rV1PUlFo
wi3BbnHF2OBBa/zdE7dy+mJQteKk1x8unX3SkaJmIV5XHDLoyRF3LK2ZD5CkvhljCvAxyAfeC3Iy
L6/KJABH/WqbfFslMFlx80/12eLYTbNUKvIlutzjUIXEf0glKe/zcSy67Pap9hnjaLvxCmat0loa
LJf3t4RDnVoI9r+pvguQY1WTavBBhfV/9Hw3H9QijzlcNT0hLhkaXYBY8cutBTEUGXYbj8y9QDGB
5DBMD6ge2R0tzIiKQmhk9/PzXJS6NelgGURIrSckxXMdHiGkRv3/7ZIqu7jP+Ih6ctyxy6otghDP
rl8j1myb81I3zC6UbaN4VQFZFrPrKNd+rcdh+OQyjkUSxfvcASco943zxCiRfe0GsdJP5JwS+3L3
Pxsu+3R+Hm2eIqhL1sx+15sTG4EK7o4iNWkBTmQsbxkj7j+uUM7cnH+WVqYCollisl2/6FUi4ei8
4ZO81bw7FS74xNrH9BS2iOzUM9xj2KCWSLkDGrM/qGl0WfkD/0PQoFSrfM40XqiDr9L6Gqem0hwr
DXPsuW37lpZ+75fgdw7mFjgxOiHVHXQ5gSZ6q/GeJ+cUrH9Wy1IrREcSa1NXiEusTApmEA1g0NMw
v3Ib1TllGEUETbEsfXODHUcPE1WSfqe0HEqoIpN0aj+GA/o4JsDbcOlpqQEeHXr5Cir4GaBLsD5q
5KGf2PO7iCZPYhJe0H/yR6773HdhJQOpKMkdVrb4Gq87JsZN4jXnugqtMgyQ/d9F6YghFFPBt8QR
ko6rIXOBzCNLkg+A3iRjV4V/trCN9L+mg1YPtzXVIuhEnhURKdGJbdMOEdPE6E0F02wTVcbWpJE3
iP3jVBGelVbOVc11QMWI1L2p7kf9J04b8dbowhHG1XTwp+nY0Ex3qFtfF8lfe82tfFd/bjyroKKt
CggXwp+nYt3e3KUWcB8nkCXJUoYbsLfJRVm/E46DFXCkkDYwXEdkAqvg4jqEcFtqEDJS//W1rxWS
K322M4UD3d/3DPqZVXlTELlRQ/OnIJ2hgTwwIYUEUefii6qLOerhMubdhAZNQHmLu53Hj+5DTBjY
XAa4mf/3vxvcgKLhhDjONbZx7vF4gXEsWGLSI2bjiR2SQb+O5U3mTWwyjM6szDiOO+EZ8ZVYslL2
9niUvzxe6RtAMsNpCPQU60vKyQjdcInOGWTq3Jw87CPoRZA4saW4LdhYAyeowmaRrWQMxJNnXV6A
zR9HgiItGpJqndiceJERatrfsr4n3eZRY7AkcjUO4M/mJYXxNrDRxw3apeXwSiSQHbCpRZma1lHz
JjlKG+GwBUBD+4EVzFcO+jTr5aEK6bNGjoT5V+tHYEQoOSluqANIvWEatYEYD7/K+0AqJNzPn33N
d2FkhR/DsBKkEftuPX6hyynoifKfev/Bj7s2O3lcLuGlEMYO/K+6t1+SX+OlEm1aV70rWjqLDD3y
ArHbtrKSlSng8iiVvCxfXnAXGcJe7IuPjdutiltNe9/IGhBLPCY4pkvKkH/1z60lHleFiL6KsGiZ
xsTvCudD8pTMWZxzTudUs/DOd4dHWOohDoB1Rumw/qj4efe2cEFHTfXGbm7FvFTPLgxYqWx5Zlvf
f8Xh1EW/ys5gY0AZ9g4CMabq9yndTTnZ9kBrD2/ReyjIQbanpJbB/vtrlpxElRQxg7tW3Es8Cogi
si9XCWclNEMy4/YmbILBZS/knmA4BwZfBblavJuZ000S1qipofNeCHX54+FtBdsBHtR0/xVVj/dv
VBH7yPLF+1tnIBIyraJFF/0N8/SpahAgN5zUPye2JibtvHoPUlXbg3F0fTx5rXjhQtwC+wekYdAn
KCUFLzM2Qwsldbe9vXHSb/LJpd/IRy5BgwKtoS+PrRnz3GTUEmbT3cBL4mwzs5uU94S8mXrFdqVa
zsub+h5DilpWBEyMmrSnuqDReXehEFYjB1f6TWvKlcW14Xtdr9XUOOwnCoq2dyxWHIwkJNDGMEh2
kzRmNdDeMW6O8B6/LemH2lPwHXfhZwI8DR0iQf6neQU3HuKMvFtm799rnDH/I6u+4jn1zXl5PNOp
exY0y9HmyALBk6dmPCA0urjVBxtuj0nIUoqfIsjl70t9zNuhrxL7OnpJUAksr6NuNCfLZAL7riAh
3MdNHvdTVsG66xgR1wFSQI7EmHw37B92P/2EinKy176HxU7jAt3EXuWS+xDhrAi1eJM1fGlMJE8L
BXnb8cpjyg/TLbRti1pLElDdSgjSvsK2nELJmZL431nSn1+VqJYagEnr8JjV+5qhj9Nvrpm/py8C
rwykd+6IenD3LJtw+f1myEKhztr2MaOvU3LlEjojDLgx4UAYbZlPsJNM3/kVoB2SW82cOpbjlvUs
BbuYCHT6XpQkK8b3ioYu+z2s2q7za9WctbxBhZ30ZL4AbtYIgT7J1DDhtG5JKQYrOmt43H8IsDgc
eQqgEppqeH4E7MR8XnrtA2M2GrRuBvdwsbhbcYKorc6PTXJ6lA5l4hnTnDDiGJwkUGtgkQ6Iyh+t
GspiftKDFj854n0hL/xU6Q56qpXM0brLHEOIDxCj0g2qRfUsX2GPq/edu5Rjm/2hbHvtyJmK5zos
kroYNYKTmy+XmtVEVMexo551RySwey+ieQhGL9QG5wxSuw9mt0JY/I+mmKRsaQSL2cS8qXTC1Hg9
fKX395uenai/zVWzFfNFoitnhW9kDonBhqNBc0MTgYcRpSrpj+xbJq+TEzDby0j+GGeZF/pNTgDl
OOvmmuVwgEY6RVZ97XmGIc3/XV7/2a+f4i9l04lc2SCI4uFYXadNWsEEoIj6YoTYcj/GPJvhTtRg
D9MsrR9S/48ygWdhscHvAdEow4aV2Ok1c0g7CDzf+hl2OINHT27IS2eP/GrVJvsnV8Ok960VXaTh
LZVRBeOdZl+2I3Yjvs/QQNQfSLABgS5DsGXpr377D2MMR+B3WJiiaovLwgIojBUpgABlCTIN3+P0
KNGOFGWefZQDStc98i+6pPep6qKavxbJqJsnAgG1EORfPQrDsc1ln3rJktZcChK45h9+baNqsCt4
e6P0Y8gHJHszYI+dYNR6ysfhE5nixBLs1MM9O4ZrIrmxaSvsmXCLnfkRGXkV1Suooxu2jalVyOvz
cSky71WWx6++7UGVYdEKGO1cZ8YeW+mZ8kOEzRI0OjDWmnB4YN7piBqKoSBHILIdwStKEraobvwI
7kv2hDcdv9X2YEhjSX+vZig203U8CaUHE6nlTTIU0xWDwOvshoGrzsamBE6VB53ccScdzfVBIYfa
bYe1+jckcFuavH92fr8DC/KYKx9CkdeFTADxgqDjvOK8Ze/aVoXn1K9XoJ2Y3BO6S7vJiqkYL2k4
6UV6WY4THXMEPSDqlqQy9gZGVfoVWKlqpaUw3S+yyXc01XA2HeG3rLuGMVJ9vnzh/aDl96IcJ3XZ
FEZ+riIaPojzY/eHGgc2joP0IEiftL6jByX3tYqQy+ihcoCj6H+3oOOcQz7IOl3RSuXHJ5YRjZ5v
El5h7XvJfcK8YNnBpggxOSg9JKI99l4L84lrQ3eru+OAeDwSti+f6LLNpEGB/1q4mw+Pzmhq8aDO
/6M5bwukggO+viryQjcXaJfGyauyfmoJxKtfGU0UFYOyr4pROy/d7/W35vsDHTl9f3J+GTzM8DD0
apaUyUoY+4e/C/6K+An0NpJmt9hhlyEWIqvPjkcVpGL4Dgr5UTZijmxJIbSa7NEWZe/JSuiduS/p
SLFmeDM6eZDsvb6NR1JveqRNfwFkHfPW7yRdYQ1m8DJbqOWNtmKbUgw2BgGQyr3vHfnKty2TCgoN
mjrppoG+BS9TYFAKm3Krqj4dcigykFCOjGp3bxg76MySGjLP0Wh4HYbM3Kv1Ye+oqQQZaYBjwAeL
TLFCduWI9muqhWuZNop+3cXolrqNzu2/oDRK31ovE+Nytm176E34q2itvs3r+PJ0aF7+D7tprlKN
t+1CvpLROSJMb9nc5VDjC1ueYVCvxDIh0u7DasgSX394+wO/W2M+D63WXhL1Gpn8muSQgruagrew
o4197/DfskZWeXxjS87iaityrV7RuDYPZGVF3A7YQLSle9AiJ5igMwaDTYphRy3cvBPlnaxKVgim
A1RI3zG4k/dfQNa9tbEMn48jZAfLeNDC0xSjZXmRI0JvSS6CBPyJsjd4lsT1upN/4O3ECGKUSDwx
bnVFNs2XsaH3eA6BTS9kP/OEcTxFVfxYcfHb/OblfByQToKkrjyWKXt/aKpROrMS7zA8ths7RN2d
NF7PwZDUkUtejxIBjyBVTAr+ZtqqJbox6ich5Thly12Wwl/TVFJ/EXEWlh/5YYxvmlfEehJwb8uX
QPdgrZa0creU6r0Cb3cOZ5sYpFXwzEHfAGHbA7B2NtnbgK6D/8o19zDarCphXBphjmu89Ehbnuuk
Z96jIoHDCAJinXLTerGiBkZprDzRuvEwGsYJLAauTZR7WAL6sdRFPkUz83Hn8J+cMp/Le3Re8T++
s9m1nNPuv7n00NC3k2tpMyVFHz/aPZ7qxYOHodFi9rp0jo7HcGLvqkH5Dbz1F2DdxuX/eD8k5Hpt
PSvY/gz8Gptg8X/dTPqhmqfdT9+NtQS3nWJ81f8p/5X2RftOIg5F+ACF3CZRFb1aSN2tvVtqzQSn
ZqYu+qYKlGYWX5fGwN2wY8MFpw0JkOaaWoebdPdPajaJkmWcoZy05K7kXfN+Zxo2oJg2mQNxRo5d
kZcU1ylff+M5a3I6NqDBj6AgkndkmCE5qjEMQBQQUJauxwg4KNAf64UcNNWe6oVUNIMTO+0toRe7
fFaHNANMpsj/AMMrVQUjIOR989D0uD58XaJVR8xggNuxJiELbJ5eQ7kO2256UH+8uK8SFGfWk3y1
xEeqodHeiif9MNvFPEXMD5nWlYfhKywex4z1K7vlmqXNkH6fhMDlJNX5QROuY7QiMbg6zKZwoPIp
JbKHHfrbk/ZATzrGn6iChNYJv/eAAN00dpYRRu3BMCQz07QKfB/+bPJrKiziykIvBrpLG6nimtK3
rIlE3Iax7twRoU9pYozPeYMhPq3aqkpLVLez4d8UcNM5pWRpkzQqOnMsMSVdguWq0trrzfl3irxZ
mBDc9ZT7wf9kr+wepHuUeFJu+FQZukrWycvfLAhoukUp92N90WpW4ZcE83rr4W7e1wWeRh4/7FFf
S4QVKkTjKfHyYXFE4Slfrxef0iL8fO5AZ74nBSFhUJ8WPpcqO5dhu7AUqbNLKrJK+BQSUN6xjs0m
mnsBfxBC0MvOAykk+EyDX/tdaFe/8ybYss/kNFBiuh8BeZbfwBank16BzRkocS52n3QSbOyrXDau
VKLT82A0lge1vnvivVCVCl+JL1CuoNC0227m23RyrV7t1NtHh0RDUXLvaAceO83Vo0i1+GDvOECf
+ZHTQOSYCPOOSsSACsqTV0n6Aj/9+Y6Sr1eEugKzwyLYSPJGINcROW7f1FYlUWVGAI5TPf9bhRyw
gYc5cXUBNtWpK6jH7OSG3aMAzlmh8Z5g38XO3j9QcQGWq+qCt+lKO3N+LkpBV37gBcJwqfJE83eO
vf4DuIAEAT1V324ffARsBFuCVPG2EdB0dAU0n/ipxEJOoJ7jyo+y19MkCIk8AIXowDIY1mLNw5bk
gifHMo1me0GlXSUlobOafmqS0Q3jQgWUi7KgCeiuZKB2TGAkwU2Rlfj+YXC/R6gT+cnE2Ii7ZpGn
wJtBta4d2yJUF28aSoFTuIC5OhRndooLTO7W8b5Uqz8QtQ2yjfaEuggSAwN79c1U/Pllo7ICUe4b
KNJIojkehIRTaCvNhVhTDrZhSvd2g2OoYVwczlONJE9Uhr12c4n+8yavMBUoDRQfPZZpWOpGoEaE
uaBFrui+b6k8fNBxjdCGpiix3iU6D366gqVWmUC8VUElmkCzQo0ctQ5qR5RySOm5RCoQMs4BTcgj
omNmNWWFBxgNxD9cOAkJc9/ijwaKS6vKMt63z+eeFXOU0/HjDK+XjihfDfbzcquQlNC0G7jua8UO
AIvO9+kVKssLLH/T614m7HhYaPpPvZ4HUPxyPdAb/J7Wd4ZaMX7CWu7cGc436Tuo4eeUVLx20t4d
/0U+DDkezlCMXfURwWmCm4nGk/dlMh0pczYF13MM7Bf4ZE7V5/eSsq9jjas0ArDYzvtpzJsgGkzg
pwKl5jkGLQfHnCGGLcP+txg+eiwoCo5cq9e5XaW/ccwsbtkSmaxYN3ZlhhYZIOb0qN061Yv361fP
qlN1/GRPUBnKo0Fg4qA8EO41TgILkePJEqEyeVkVuI9igtOfGlAzSJ5IJwAn/mbF1LBjugGYD+pO
jPTSl2KPs0AUZ9Jn0Qs54JtjLx3f8WMhxY+mx/MT/FdSgYECNT9/xTiad1UWBJupHiImsFbEFlcf
hTTY9f5+92jPX0CUMigMkM8Q6vejamVMLp4bipZGxu/nh5w/mQOfWi/tCXU/B1oMzWI9zW1jIq3c
sLs3yM343xCbz+gWXJvwP8SFnPyOP1oYlwVoXuBXCiNM/bsvHEkMwKn/P8Ye5JNp4af7rn/nukRY
cag5j8IIpS7jcLVYKemw6EPxuJkFQy2Hr8Xcq423wM3vkuCKblJ0ECVtZdusM75AeCLg8FFpGaqF
Uy89+ao7hWbDlWDnBUz4uq9r3228JMtTv6m1nS0XD36ajpj4ZMed7IrS9jArfvAPB0mgVv4roJ3+
jpkKdt/D1rVNqaiekHXbSOLt7CZY7pVZfkNoY5TvlZjMcrJXC3W2NX09NAgmZYEa8s3x2Q/KlaL0
BaCrvTqciHNYuTmwasdHvre7t5/LIkJ0znyKqWOq+QzgYOmcQLcVleSu53MVFmk42+CxxZb+Riq7
wnKS0OKt+OwNEViKWZRVTQx0r82/j7pwNXIQc8SxkbH4Y+m6KFlAm1TWLsIl+yMQTKy5lmbcKFrF
ZpIyg3iA16xYkPqMiwvISEXJP+Mr7H/U9V93p2B0nlF5lXNQiHoDdDOl54CBnxPiJy8PJY3Vw9Z0
VPd86WbBSPSM9iBJirYZklA70IWxt+zcKklJ+wqHpc30WWkrC/R8Ew8UTGGWtB5h5GaIMdGg7abv
UqaTHGESS2gIbeXHXzKw1Wob6Wa45tnGRGw0ax96SHySo8VYUMQjfwHoMQFL4Oeo4GHoW+xgyxtR
CsmKBUXbpzKsil713ZsfcoT0am0i8eFwOKFeLK+UtiUPDth681I4BOaeLuzPPLrp1EYJhbId5Yz/
JbKBiL7eeNUBU5ExfUEWxsLo4dz+xQ1O+wDEA0Q4UYBCUXvL7SLyKdaGVYjOUtDJq6c543zmIO9k
6Aj8R9mNNKdd3JSq+kM0L9wwgiZRDT8ryI12TB28+5sqNBPcznCWWOlstDn+vsv/koAnJVuPch8y
cSzGO+dmxyGY/+r6dNrmLGqcYqhVY1igNCzLSG3uOIYW7HIjzgpnUq5pjT+JcsvlVty9nOdZFRWE
AMovEdvuMnGlKinqrtC9QWnPSgKFuW7fM+jbavWYplaQztNxO2mKMjy56Dbzt55FSr/59bOhtfzr
IYhi7ZRSrOEDA7mgljxXrX2MOwFA6Lnxl9B8o5Dy3k1kP8L9Cu7OSqhENNc75zrAkj5g3VsiR1oa
CUKsIGVaxYdZELex8zVfKJAejhY3YYsYyczZYPnSgp0qc6j+aGxpc09I/qzNlsRJu6X8MsYFPuzg
AFLyLXrS4cJ9CEK1Ga2q9L9GSE8w8C7cV1/0ws87dVqCzOmPmDYaNrKM1Bdd1Ddkqr8Dvew7rlsJ
rQi6GLHCCE527VAVX44NZCJ4lyLDjPYHZOIuaqw9VCbZS2maH6rNZ2nDewWUHsy5eVUcEyMlbRjf
J38Ce0Pp1A1abzXxxqnQVCqM9AC4GXnjz/IzNdST8eUiyaaOGQgCwk1i3iN1KJoRzavxEtiN529H
JvUoOMU0mbdnKD3shwFIU3jTYLSpap4E/g/6aC9Hky85yKP9FfSrrAT0mojwfvdEpH1v6S33cmqe
1P32Drek9Q1whgZsl8jAly99U4P0QE5ag4wISSLkQgl3FzHyMdAcZ/gf3HSw60mOvbJ/i6oH1rlF
LcoADV/kVzTz0SYV9Ge9K4JX42Q8r0L8mcopTFeX39qaHu6HJ9ScGs4UbvQUr255OqkMP7J9tDUZ
bHiesxzEsOULMKS0Hp5kQlMeo0jVN/Xd/1ANKohH+yCDrEUKIshLTktN+Vc5GzcgtHlGcvy3eYuw
OdZlco4nYNfLt+Yr8sfE0mErib6XdATLjDLZfUWjru2FFEBDOGPvApGN6n3UoxgOLvifDraDi5q0
4IAuRTALQoCtsDSM8iJBN8MzfPEtwjTzTgmmX6a0hGvACB76xxS0ddRElD/9J5ZNlfQPKYOrnUy9
sMQBDg+Pxl/JTdRHfF2srJChvwOJocENUz7J5cUOXe0zBodD2Q9b5pvrmmxrzh0oAFRozuFJ6500
5E1wfqVCWHEOmOw6MyKWwBaHyb+PsuSZ/WIraF6EOui4IuZZG3E6b6DN75WY1A+h8QKxW7FEGmSe
ICLbOkPEvCW4/HnmHkTnpI2VoWmME4W93u6TC1EzxR/3rwVgwSQsXvg93RQWRoKKMWGXCfVOkEGF
jJpPHzRDupb0NwgKwFxcKMl2/QwRCyio/Myn83dOqV4yZffIE6UJZ3k2SgGMSKUn9uRxFD+L4iq6
PkkzYz55vpzNypmyXh9jlmPB4w0Lo9byi/kdhh6HQvXJriuPFS5bUxJlMU+PkRsRMjzWLDOSAdq/
qnSIigNn4udE1Bc009PAd1vnP1VNeKFSzlSn9WQCQUeDIRDfwmR0mkfUgfFtpzANB3vMSpl2m9DZ
acrcV1Ym93PUaOvUZxNYmTSThFd291StXvn5dHsZI5zhe/Q4L7bXP6zyu5lxsisUc85Szh3nxI/N
FlwtxGyk+7Jl+gGT4rfAt0fxID3WVjzE02O6thf9o7tOwH+QjRuwXMhPf333kLai+3Q+FAtNsmTM
zwIkR0KKikPeDhyTTEWKMWPVuQ9ISHuRIaCZzQT47Nym6MYuYnekLcjvkp4qZEHWBybv6Re9yjt+
ip3AOaWYmGtzjMZKhh4ifbzPpurVJGoNxmTKX+7OUlWE8PO9MpuX3gWCbcCLpU0FA1DZz4Ov6Gdy
1rF+/TUONE7MSOOH5J4dCfd57gK9/Lg8iBe+R6ryqPMihawsQcliCkmAnnOdLk/fnuSK7bUJurKh
CMKsm6xPsoWi4MAHXLy3zQPLy3rRssFMcUNI01xvk+YLI3Nj7X7D1Bp6NfiNSIywg6Xb/6bdLSWp
jK6N7ONJVs7Vzw4suK0gaiShQYLGoqjTBwrZQ1rpLSs9aYbHpDYs4F9QAeurrRRvAzTYjYlV0NI9
HXdCW8WuI60/wrXMoSKW+50nqmsRYnleMyiJ6olfkQg9sZlT1Pxk3My9GUX+O1PtvgxC/JoCjb95
0iabDTLayEVQN5cfvBW5mS1KuP8DTwok9CyKQetlFvU6gFHE2HPxRmbZXdNK5ixjaB5nmG2vHL8y
nqLmty/uZF+cFwfwXZb7b5R7xmdgpqNhNvlbXuWjqVo8DVJMj7VlHyV8W/YVHqp15g652b43y7ex
XJFU3lC8svWvv/Ix6QuyorJuu/C7UEuYLtT7laa2t5x+VM+9EkxdosqNUntY3R1prATAmlqmRLTO
deICXfbtmxzkvwy7jEPQzlJhKeqauX/GtYhhj5DCM6z0f9anVqMQGtfpXnTVW8vOJrid3JqDGQzW
Ofi2Ih4efoCgaW4IJGNNJslNeYvX7eQOZKGPs2ei/2Pk3AgoOqIOaVLooQQgemJ+rAFDB7UVT/VN
bfJ3ltCcF3RdqHiITUYV1JTFH5AHisb/VOhsmgtkwROdPdBJilPgjMVEjMUdelbG/h/86Tl+EGR+
X+ZzGak/rsdzMlnUtIku0XwMqOZFFABCQ2X7xNQN4C6d1WI/BHai0rnrxIaRpxLU+1d0cM5SHLNx
v/fevaLLbcC3/kMmjQqedAyLYUxVCrG8eTnjUkfsgiX1D3AgHBAVHZdrSbbP8HyoxCA9pndZj7GO
xjHrmx6GoZx+P9TBe164AynmclI8c8A/nSE14qiMMqiTSYZKynEqC8zA216iDcjzIKYAbgPck0S5
3PpupBssjBhMfaLqPp2c2KPGg4OpynPiIIF/eGmkCk9lBA32qQOUTQUOAk5YBH37d7cNdw4OF5AA
xqwWUh63llKtPwmCXHG95gpQ0IL+lmQyjEORZa+sbTCwpxh266fBkR836uBjXvg4r5L2ic+ESSJX
4amGn/RPjm2LDILyR4xBC5zFA//xW691duTGKygNSjiBUA5hL5IsqbxdmGD//sBeNfuaHTIXGQei
uoKI4hK81O9K9nRrxak6E1uCsVQ9bTj44443Z3nEy5kewcH6S6bxUf5nxa07nFrP/igkGk/Igm+M
lW+bAaVONFGDTsU5m93JIusGHX50t0nXXVaZJgl4IPD+GKMzBGNBv0PdaHMAI2Me5r9PdhYczLGl
IY7NOC+Ia4bIbP2Px/jplDVGxRq8UWCwzSF2V35lIEvyRs9eDW3DvEkA6q4UJMLyu4nIKpzOCcKZ
dCKRypBsF9LizEiqEulbL3iae5v3ZEUu5Qui7AnIxwpe7aF6ybVxFndFOejFHTVUBcd1Bor7AoWU
hXU/q12huAW06B0AMSxzSCYROUIXPyYAstdtugiujfxedoqXWBwUrBk5988r5lTTkSUtyc7Agial
/u4opxy2CTj6k6jmtSEosyO0l+Vlh6978gqcAhc+p3bc7EMkZ0TuuzZgA8L1Vfr1/LPuM/Fp9n3z
c26ggEnuJGEz6xmkmTO8RXD9UhRLANbpNWsKbe6nQbJnZOZTGMo1dfsVRw2LSD+Xe9X8Kp3XpiLN
dHIAwnCugshlfRIbXXp6W7Vs8ci1bBdFaPfhX9UBaCFq1mox9NBQuY3FeQGJoqs8b5DyU2FghK2r
PewmCk9XZHQcTO/dlhToR2i3CpRNGdmDYnIFRk6lAT8PblJjF95npwh24o0/81SlZqfN06rKNEOK
8Uj/CR30EcJrRSzeFP9DXbBV26fJ3uZ2Fit6E45aeK57P8SOtff+pWTy8TlQHYrv1C5vL5l2KCxm
z9SA1kzcSY97iYdju7PKQxALSTKjNmU8gGNSemQ7+vJcKPYTSFM21/cmwrHOe6O1LqjSRajiHmf7
aVEBmhq58yGtCS/sUF6adcuS2xT2JqHQ9bgvQ+T0oELEMLlqmHf/jM6RYzVxBaczVOcgTuyRfUMI
gxsgtpCntQ/fUG88cIzwa0NKpezE4ilFSM6l3xkIVU8RnP0aF70G5JVrWUxbmzXpShAshDnQrHBn
/A+UGCZIqPdtwpJShch4HqKtcu6jK5bCwEk6TNMYsWnhYTLZxN/2vfJMu8GrVhEeXueNK4CBZGB6
leRurVQjn4N4lnb7Q0M5jc2eKbZvqqpeTJrL+jz8jNOgJdZ2wgjmLtPn9Ic+hGI/Yw7SlSBbThEu
1rkeFhFrIQIC8sQQYzWq+8vJuvn0/rfPG68pMH6lZINwDKtx9htXIadMl5TEJBnDqwj2O5w8NKcg
j6Q07o0+ioJZ9yFjzp6wCWM52lCTEGd9sf9PUNiwB/6Jrr+6T9XkGu7RGGsyNn5lVAOtWZNjhlAz
1E6/SY6DMob48dZSMHXwdPztVsSo30pmmIy8tJxaTyErpGi7EglkWbWl9A8zij5tVzFbdJMEqKe6
14X8ZrviZd4QGZBU1awN51ChhCDP+9Y9j48BdlQUZKmIF0zdyIuXyStApnD71+up49EeW4R0QyOb
tsFgqYQAtIkhy7WHKSwgMYNolQ2nos+EaCYwy/496ngV57QU20yVIktEv3e3d/N8GPN4GZ51pqHN
oT2jWM72sU6Lbyjd6Z8Wonwq00XmcU/h5XbBoujI3TgM2FROu+aSyd4ph+fIoOOI/ee1fzR8zkck
urL/qnKNL5V9T9rqKb0utco8WJSa4HaFPBcstjBs6jYSG2arvT3VCLZYmUTdY3tRQ67mMbqOXt1S
NDQbdwaz1KSYPR1PWF3SxY+9LatJUA13a+Y9z2W/NnaYXm1vNCSyv5+6Uag3n/fpmn5mkRUw+WI/
P/VU0xbHhBGGdv+wAXP3iGF82lus6odvt9hTpzGpIyGX/OOy+XlFOwn+Xdxr27OFP5DwB8N2/xRa
LKUryo7ICV3u0CXd5vcL8QMTE7Q3guJYgtVPBKcHRto9SjOSx5G68rix+jT7a0xs2/cap9RMvXfV
Zopztwh4rHPO1GvvT1b/kmqIYLqpZtPjmmQe52kBMj9bj2m0lazmOvVgdFFNOwgprKpP1DBuY3c9
S5cOpz38hU/N8XIQpc0GrwwXiefA1XdJrOpfI1dcTJOV8wOTFv0+fk4/rRUmrdEzMBMMLchT9fN6
SIn/WC6T9eeG+tC5jHYB3CosFHA+M+FyqMNNdKOusJr+EL+KPkbbDKjZk8xv7GOP5GLmfxu4CnBv
qecyT2IxbmKBm5DWx06M7AXkxI8fu1WaGKcOQVZXQR1ihReU94go2GX1woZW3FM5/t4iGApx2cae
LdWUoJXfCARmKsI2yW4D5Qrw1LPPvwZitzWLuqcorsnrPPdRVK6tD4feekuWYjncoX8qRHbHzuKd
vp/SJm7psBvnu549SwJ3IZUUHjw0LAMLjkXRGw9biuDh4bYx2qHYDLI0bcSBwaC1CB3dNMHe5HiC
wCrKdSqWbWxCLarPZAZTQO9V5g/+HCHQYfHGARM5jS1+J6139art0nINwIF/9xhvMaiRJ1zqZ0sQ
KZGvCVe9gXrIlpkn6ULLj8O9vBxca0nk4C4h8djepNaB3rchlC33eGaMUsFAmySu17tn1MMtqDD8
DZ2zZIwK4TGiSRYi1SppEreaTiAdN1e5Hcb0IZkcfFb/Hxflk64d2YPEYhbLFNjawg5mXp4INX/O
UKDdsL5VW48uu5YMtQr7vBbRnqcgFtqGMDoYnEKoCx+I+ZdD4h2FO5N/No3KNeW9h5/25T7+DUoh
+iDkcb0HTcC160VoZ272RM+hdPqPE7c6J7ZWrjRlqbm2mbL7iMGhBf7UKEHQbmI/xW5qBC4t2g8F
flewVohWtJFf4JC6uCRFgIx0GuNJOhFwgHfSYPGx0KfDTqw01qZhcprud/P/GVM4/bNm6yvWCxnl
9EdSBPdNNJQNMpOSEQYsDOxF7MOPwOdI/BuJSfAXB2jxYLr8bChHEzxAEpaKnh+BbwPj+ePshFbk
MNCIMePY/zyiiOeNdOOsiebiZnYyV7c/xRUy3afBbKk2utiWORdsCPRC6cBJB8P+El03reCSZJRf
e2S/sCLu561OGHzG5zMUYINvKQz03bZHRjzoNbdFVaxP2tbxJeNY83M6A1NOSCnhJq3tjyG3cKDY
pU5ZBIJazouzg2hS9g0Gm8sIBP6wRcJ3Tv9MAnranaUhiXxGWohPpGMuL/HohObyqPYAwBsC5TY2
3zOq6sKL7qAZBhK+4HZ+ghVedRSbkJbyI1hJ8JkLhZJPdxI297mjCabr5B6d/uldUAFjkmj37Z3b
EOZGL1e8mn4uxT0FxrXyFyP94TlnUBZgasWip4b3VPtP+jHAIx1kqiiEBzbv6nn/1SfdSYq/937H
JEP+F6W88u2Eiv7Ox64Vp+pZ7DDRm+A31HhyZcvoYSgzrpZUfkx59fzT7OA3HsUTwzaj7M0KIh4J
gi6GVg1kakIh/L4yKRZXCB8WA42wdz4M5r+kpUpGVbCa0Mvl+41JIDAxDvVTIl6kjoYTbZhDxjAf
0sALTGX5eYWGJtGqWPAk4nAptUblLHj99mpNcgHA5HX2/oT4ZU6VoMB3OayYpA/UjxSlRKTttpZm
WREcbmprn2ieRs1/gLOryq4qrs42gjvGSa+Gpdi9aYgPSUYGV+JO+fhD5RohilNXHj2MhIfx+zYW
qpXSuEKi8J0GiCpxWXOzbSHkO38mO2P2udTyceXZcUwa3YdBegs8hdlC+hMTfr65jM/UVqomuNbV
GlWlnKnA1vaXd1N+o6aZTNg1MrMwAiDa6k+wzfgAYkCX5Q9UXTm7MERX58q51H9K4kUhGVYQu4JP
wn1GFzNKIceeKAYV9TemXFkxBnnaxRqW0Cr8vxoAz0ug3X4SkZA20L6HHBs2eqIU3uqfTciPnxf9
E27+JuvXb6NmWC108u2pna0MhnxBdsAk79wQHCX+8sJl8s4bZX3Dgd3zDYy7te/tcgLAfAgDnYJ4
I9Srbmz426mM3gYZd7zhWq9CSzkXTNsO9K3NkZHZIYNLLqCSvUf7kJ2y38GhRvFpEnkZZXWPG5H9
GI8O9KYL+vXlcdpYqNPNSnTpU+bSst/wtkuxPFHwU0A2YIb1QQ86c/idvkI5WP3129kI//U5y0Dn
+SwA+s/iy1dY5myJKV4PMS1AwyM6ThH64n5TGRmsoNbciXQx1uc1zj3DnrJH+V6M827UM1Myy3fZ
c6+P1IZooKECE4NU34RmADYqh7nQPwY2v3Ju332JaKHrcmTzxfKZHxMTnDhkC8us7m8O9j+25KKU
2c0yErwt9xdMYkPfw0JAstKR2QsMR+sg3MD1TMni55Br3HsluyRMjtqid6WT5HprCHfMcMIYMFv4
OOHtIA+H4J9Q25ad9ZqlBBxek9djUFb6V7s5ddallrt+TvssUNilI5h94Xu/LN5FX8jFgHRDds3B
lIE6VWQP8cLkU01lxm/RobjCelhu2lXjBptqdxIeBMx7QnlME+9vNjbVHFRRP8HdruhPlgDAMT5T
HFp9aZYG8Cb86DvgQXTgqXRvKR5hw+MADa1JXCTsriYBNqu/aXPb990UXCHA55MQ0FULUipYxNVi
VZ7PQaMsaOXxeEQU9qn+0zgGWNjsogSByrH7lTdIJKCl54eXTsuqz7z72vomzkCwLDdjh/rdYvJs
KKybRtSU+UARCTnDfZ7O4TNr617R9N2xZiMYPQsmzd04A9DeuSF7YEvoaX2JAreqVbFgNiWffWvP
v3tqkXbUrUnuQ3/cpsp7ncSPlW1nvM8ERSCrRvGw8GvbvVXSIADQLRzP5mPF+hc/Uk3A8XcOtF55
SgXBlyNzNlFs0a19vzPBYG9eS/XY5NS7/Zqg+Di4HaVk+wRUe6AW3gEB0+3tOHhkBS9X3AyDyHLP
95uX1HPMQCNNquRdzTRm5zXGGp+vvXDSNuVpGnSSvb2E3eyhdGsVci96k37imub3yMGCKV4kHF9l
5hYMSbGbAh9UJzK8UOofVm0tQDH7YLf3WgoRByYrILUkHxVKE9tklquKsJaBOCTIera6DqUZkQsQ
oIGLXVgu3+D6shpPG79hBvUyWKR9/oWVI0ygwmsvgeP3AWC5rA9bV7ly0zQpZhnKbLu4Rda9odcW
vQlh+OBH5+1Oyz1amD0yMObP+Dp3zPHBVIUrOyP16GuvV03rXSjr+lwtkRC8AkUGUY6+yhFvwil0
wSqYcdvIVC73jJMA4nrMwqRRAzQSAZJB9VQ53bncwW2TzdgZEBf1G5SbT06HE4EgTlpukgku6vsf
yaJ0QyGds9zY3uhAwdajWu7af20qarorvjKpXGW6c9anO1gwBtBvd0QgisT3MT+xDpw08cdSatzU
cdqxb3HJjrkl3zaaeLc8ddZS31QISItAuT5C0xa7rtQ8vrEdv4t54Or63xqMOxSK9CjFSGl1R8g0
846NLCcBn/9yMFjMl/VE/pTETXi7mCs+PDu4lra9BNAy3WC9tDI8tDfCdCr/bM9STeFVkTdFRzk0
y5Bh3ewxbl2YpcVhb2h/m0sVhypZoIp2l3k87j0wtDs/ESP9v7WPxYpK25iUcvbBKoIfCva9zSSo
SkU0Rt/ZOw9QBUQ/N3qNV2j5KlObnqqzOAfBUquy+/Ls69wBqZ3JBZ4QWd8ot3tZFTekKlSkLEMA
vvU4dZW75JHOqvsNfj+Cy9fbtg9qm2coldjCglhadTEpvkdkeYdvUEgWN87RZsLPbBMtnc/qeF6z
uPcXUfr3rFUJI4uQMQR98EzFUGydMn0cWC7GiUni4w7VRDa3shAt1a6P90Uk8H42DANA+Rm4DB15
OxVyu2ZhsEnWLTZPJ38dhR9yMzsp8feH5x1leFGgy/IYff8Zval7A5UzpszKtObQG4tf2NDkPdC6
1m9xVyc4GtXPvgqsfvppq71+uwvr9Yh0GLqdh0O9M1nOyqU6+XS4m0ap/Ok1Uu4dGjWMrCo+7KAe
6QJ5yeGxniIlQDIWwpyFkdxuHIJTEAgQWwf8ZZq1+BHMy83p41Q4Bp0GtWi7kvxI9BSPp6DeGi3X
duj3xC60qTlRPjD+kEc7fReYpRyz3VGRcTHBTRf0ti+EbBZe7xU747n0qLD5ZuQ7PRRxBtpAXXmE
0pTdvd3QHSgTfBKUx6rI0Vsf7tZTMotGhF3yZOBel40tMsCASnXSXAZWbBz1a69jQXLm1v+oJjDa
rpdN2lIu1GlhbzpDF71323VuN8KLJRjWLNS5yhabhnvchA2CC3MbvEpxhve4lwekn0KAgGT503ga
5te/yV5yxcx7BQnJyQU7Q049UL3yat9AAVnJ38GiRJ8jROJ21yS018i1HptCkagTX99ggvgAZV5e
bma3tmV92qZ9lhmWUSxuaMIx/knVZ0+8B9wrQ4KKMuiOb55awrkOipZ+tLKknQP1Csbi8lCvtE9R
1zpE/OmPJYU/vKDoFaE3xYPUwM9ssr8xNoamxMmH1fJbCeCIt7IKluDtmWewvF2/VO02+UQaQK/J
fVUeB9b+VTqtPeXEGZBD9xykyC1uBEwXFbPvO3Am+vXkqwQl/qU0dUQmgN+n73lzZH4HlYjgkgNg
k+Vf+oRkkcfBDWaS+SjXrurOR+Y0YHzOJay2XlTWvr3+RcKzRch4D9cOK5iAQ34rLpMP5ilr0nM9
72CxMIT+sRtX5C/fVcHUFr2b2b/BCM0QWkDeliPAr7QcIwTjdJxPsBKuiUG58BJB1+KCmc7BhO3R
2ncGgzCTieOX/PTiQTjiYKF51ikO3Xn//bDcIWi+E7CWL+wIAPRwm1rWoI04k8kKBbvBr0yML6MV
FGsN8aOT42x5Uq/v8ViUOw8m4pThCh8yM9X7iTOY1bDPVmULJ5s6lriOXU+byoXH7WCQ3y+qM4uR
0rrrP5T8cQLB8h0GadG6mRQZavFA83/H/EWY/dqpZmE49XAS3mUe4WPmyiNIhLKJqpkJcXprTTDi
3ikYgIKnVm7hHPs4rLnqw9/fwkFwhHzNnao6ZADgHI96xuAdvD8GQhfWa23LgdXCoGdvMqXfxtox
8pXUQC57nSyNbmlWmmvlJKvAj8EbDxwj2r/FQFXzm+iZEvqz/1GV8OSNzgDEvPAFXwf53vzrdQap
sOqjA+tyII46u4lNtKIB2tJOqasvsxcUifOVxc6ki6KdE9xk4TNIZv6BgXVwYbXF7YSCPSe9VrIi
UE+UMEh3KNJ6mU6crEEjnm4CnmOJ9IA269pxdTqxw7qw7+5DuAlYPJMOYc6y2IChVd3amru3XU7d
tA+YI5CVx+3K7TjXL3zIxk/LkmE3lcBMP+5dcIkWptOrcwlpZw2rZXDwWc1zzKkb2K7BinRdHxrz
tiT9BHUMU8EhdN49/LXt6j2ztcekH9dyKmfaPYc8tGHABfTRyNQO4s+I444GD4u31isDZOZ8Hutn
ajBEi0ahn5khA/TjGo0ah3iLqFYc1+yF7WHrdgdTdo1h1dhfawICooRGJP0xbbnxcEWJNzbNAMnT
rb6+jKiE3qFiTKiPSXP7cXr8SHFNUhKLo+PCPrXiOycF18cvSCzPUAVXB7KaOtbEN5OdfGTpxnZa
KGpONZ6ZXnfs+pTDMO3AGT5B8hTAi376mx4HX3Y/H2OUKWFBtzQmjrahLvwkoW1kADvPAEjsUVV0
G6XKeRrYCwVzA6nH9jbRC/TLs+8GQwomsCwEhNRXkRAaTGfuFjo2KNaIekfAbyF4j9z6R8Nvre3u
qLMliLZyzkBTAu2XQxqsT915Kbzp7RIpR+/JBj7VsTUfD7pyWhwK/1bFCOkbHJJE1/DZC4mXW2KK
9lP6jEGrKcIgPwxhaiyhWa/WPJSLBhpxXmP0UjdtA4SqhDZnAhPjaeOdGQgHCKXfU2YSH1s2qOKD
CWz/Dh4QkmSqzZHKkwic+MZN2Nnd7J4mej9uk6g5+6jbIdgxiR5gVGKHsoORdCDZBr2cntuyY/Yz
d1/reIiD3gGSA05VZqxlhR9L9SfaL91Zwe7eB7/DPsNrzgfEBL6W4oQQ/ynlffoh3MIvRwl/O/cy
p2sDMSYefAbDPavxYoqSMpbA7WLaLc0yuASVG/rbUMKGLjAmcvl3CoXmVavX8nCbGo1TXinuplLZ
cvdbuFpSrZ7Vwngg90jLcQ7evtGde+g2buJ/uaBagAgl9AaM2EffmgH5e0dR04JjRD1yA0eXwVYA
6OvWOnlA97o8A+y0NN2etThmDxbVc02PB/Kf6Vlu+9l/hpoRN1Zu/BSYv6sGacEwsRT2g8RcKtdq
CfvZd8VkBW/flZCB+zPdUqRaQSd6k6/bXxy+uKyMNX/5vR/GE5qvlKE2JlfbK3/RscwAM2v8Jzk7
yMETEX11KJgCH9VVwi2+Z0pCPSo1mvm5P/atM5qBIAF1vpu7+3vVne7FR+R27GcBLIbgZ9fjEkzA
E3YzPwkWJqYClzOVaau4Qr2X6afZhNqYz0IP007BfZGuyD4AL4ran7Ynvf1ivyRORZUjCc/0NU/9
hDk2eZUj3mXfzNivdsIL0PQ1D248MYDFSl6DVJnbzXMiAlUewKGEpKQs20COVNMuV/UyATzFq4fG
fQlLfJeurwD9d8ezfi7UiYOKEn4Jo1c5sD6nIuSrw59ZVPTUBnCo6mfbE/mYZ58gZqF1hUo7h0Qk
i8HENJRr6kq6vMeDFJN4xG2DGPbLrZFVm+hbVpB2n5eXyIhjSXNcqhBM0VwMKqlUEIUtqHAoXcw3
aSDd297IbFSslY5Gq4RbolsRcMRcfByT5BrrCwENq6IKLQQiSt/jRQZzjUkZ+K0CAMd7WIJ5ix1f
dP+vYKqRYkg8fKQBJsI2xx2U1ZsWks/Cs0Ny5T4FoyBS5kYeEp1GxgfJCw40zyUhVHzqIZ9gMyDF
IPGySIuGKdmHHa9Bk8GrUnneVK8q9pDWKmHAAkIDi/fttNi4cQp5q2weiJrw93nqaXfrJ2PJKMEX
2gyB8d6p/A+3K4jeksvQ0eqPoJabiVe9uz7PcxbsW1jMNE3WYALJfQjr7V9W57q3y63xUpPaNrhP
e9BGFdickH2cczNA9Q4A41sRJpj4ubZCBUc4jF9cPGMG36B15JgWsg2q9e2myfRrUGadMA+oz1OO
67PUptPkq9vX52sPsMA6oAwNfwE9XyJrvgT4qiISQaDA+yzLVg0dqD00KNA4/003itptPzuXO57U
J3u1ioUITnFk+0YRRQASCfV1qffrA6XxGnGyRvF4CHogUGTFncqkAQ4iFq0bWv/4jC/5crLSielc
71BWpOiEC9gJQNoqA2jgEQrXkXTSqASgFFDZBjySL6xN97JSzzFbDNt2w3jNNSyMhyxnjrhnsXtU
Psdc1GVGycMflkUO6UWkfxL+UDBILZySvLfqFIGWhsrXSPzxurC9V9ae7O8jEtU5ju1FCHQxkLFv
igCbxFWFxt1eq1bnBpvKevlIUUzSib4+LWeSmTvezRn26GhvMYxKeiN3iJTv30ElethPqDUcOspt
zPlQ2jd2BYaFTB1jZ1Sd+fgla0isUR3sBWjoxNwmfHvjD/XIi5Zfc5zTWQDj9o3ARJ0G6KY1CDNU
/pXxIPi8ME+5g8EUy8+VB/Iy2CpHHoNZaSO1ptS9xG/88a9MyjBda16BSufNBp/84mNINGiC73r9
winWQdQ366zkTBvHQO+bvOA5Lq5RnauBDK4AscptcMwaJOe4q/LbOmukxiiTuo59gidK5TRkyD7n
92AJv6qkvHRX96e07w83SzN7MWE2zcr/wp6ZM8ruCKnTGGM+aPvz22MOfYfSMxbuIkS0G3+1BC1W
DOsm4ibqnZ6IiJrZpm4nW2QzpfZppFaWKTEB+o1dzkSk27JSgyMV+K12KnZe7XrAenXUQfzkIVHL
K3z02Of+jRH7CZtZjSTIULR4RnE8WoLqkoMwx6IKz57eA7amdOQnErMjq2vAZCIH6BZBu4snwvZm
sqKW/y+YweSuSPF6Ao2/28dMwU9l0+LMuYpj0IZGcWmUXtXoUH8bG8YD1yOitd5b0DJ2PJ8pPJg8
GBIaWt4dnPGAqlLjSrtLaQMID3T2tzfwUbtOFR0/fGXETYqxHauJMiuj/4pDov/qikNdHGsiVt9o
mPXhxe3wSnNlwSLAgFFfqx5tCFc5BF/ey5WBAsNZUdmoFXa3/L7MDgtE3DZwDR02BzarRdOAw7/G
rp13gv+959NGfxbkJtJqsXLLxSgIb24GtFUiY5qXJnqU3PXlWOchAsG6VAkkNfvH2yvmZrKaYuum
bh57UwYS1H9Uxt+70iBkhlVjkg04q+sjJlGFWiTqakG8YErRFiG1bn5ovvO9o4E2VObi8d0xrI5R
H4WreOcN98peYEqzPsYHDr63CnkTX1G9tUzkcsnn4a4SoxxfVGChg4ZxkxS15nNed1/T1DdfM/oi
5eQ9CumJfly8wRyq6EYDTCv9JdtSAhXALB0y1uqdkhUAd9O55jQWJwHKY8j+78j4HUFW7r4gk/KK
Srz8jJ4HFw9NIIDE7CW6nSp8J+IwaBkIMMB+AOAtnoWqLmRLWN1g3IOMR1GS7pGLBDm0dD41dCzN
4DRflEiUKNwGXX25nS7c0d7wJS+pUkqhqzSqJeaGXqwzIQx/GxaMa5yifejywxxztm9qyTMzSp5+
FOR35H+vF/uft6eThU9MFJpJIzRdw5vahK5RYI5h7E4/LVvjymeIZPWyayud5QpZsOuxvC0f/RVQ
bTb/yFM6lFfHYb6ZuCR8tI78S9NWdA18Oq/s1M5m81a2aUqZt3bDkl783vMNL7PrRkmeA8/4omra
47n492fnMoEzEoM5jfcBno9Jn8OB2Zz88K2aiSF+Bkp5ptkMITpVFqKziRt3KWfzKhoM8M1nvsss
Mf0ThvU9D9FUwxVMXxzWUSeOGW6/dRulabmNWkXHtQ6151bnMQZskg+prkveAgNUP0wTe0y6OoZ+
XxSQSdBMSVA6a8mstPsjeJ6NyF7H7stdp3P/luY6wT5E9svBmW6HsW7HVRoNdJbcuSK8EzTWwzEJ
OAUDlQf6nsEK1/BKoEUdaTJJP0K6k++dJ17xXO79Lnb9c+zZt236PU3RYDihnSEbSBZ9i2usuZJg
HThTD0CLGrk2z2GhUUB3qJZBQ94WyEImXfdWAAR/Nevbh801/FQtZVj+sccQEywIksENWh3J0zi+
eZWtSvpE020Jel8lbQuHf4zZ0EU/DM3t+PvHHOfpJ3Kp2QcAWIUZtlLpa2mzJ58SeYPs5fLgcuse
17h2xAESYp3vmVFJ2QyrHz8ZgLLrZCEzTBx9Be4aDdsbrM9cjUkThAk1YXNPFkkYLBN/Pn+AnxrF
T83sUW49rT+3D4gTMcZTW+3PCdScw/Phz6IAcObwK8eNRph0kEWIiNhvCdXhQCaCubLBuv9bbIJB
QXb73mXojd63vAqWMt2CG1tZsAnF0VijjOFk9L4Z5wCkdKrDXe3TeNte7phggVUgPBKp9Q99MtEc
aTntFTg/IMwDjgtshUOIr2i0B61qjTtJuO87mikzmL/1mtUDOdaxsuZ+E5rYRdaas+ldBlDgTFHJ
C74noakaqCXkvVSo5gkPBlNL0WVYQiClYblfNzb8WUjFIgVnxcmYIMiOHe2X9lmkFVq5cBBc9Xrq
wruipkArHLCTCJu8vRgA8UbyMbczxq8NHb6+WvdXs11FoimRbAFdfZ4N2Ug3V9mGY8l/K2JgcS1b
f/y4/HZQ9rgL4cVM7Gf32Hj2L36m8WQoUYozdsaM6TS7iKfDPcCQZfNYxh9DLgmMxGjkfPR12TQu
lI3UTOg079pQfkqaqlvfZE7c0xBsU5S/yTKIjj3artkgabtssIV+cy6+Ui++3yfLWITOw2Q0vtKT
W0ZflKZyYm6nke977KDEbHrRewFl0zdrecQav6Buisfq7BsSuPraEB0TERWltsKCIjfqczqmyhXD
dIUKDC0cF4+7l/fj2SpliaIrue4BnVy01/L6ZRhr1euSR1n4o6rssCmNc4FzF8VSvQB9nQC0cqUF
aQjCXl3vqy4qWKaDNBto/LWONnubVsVvSpdCg0i99tpEVm51zPa9mmswCboC4BSV+QzfC29WWXd2
Tf0grIpwXW8VxRwRxs6+kESimhOCYc1oHNR5c99kt41b+ypZPY/kgakb9wZ8I/WAbg0Jgi2PDOEU
xAjEP5wR9Cko33FxYbxhsi/WLhcQmUpaP2D0z7gPw3kFhoasYZ3fBWzpJWKlWiIUxGW3Zx7V3vw2
5tCflt9w43daYvRVWpX7/E+7WTd3dK0iDXCG4f3c835Tk1JP/iVyFJMOYBu8pPXL1+caDW8PYeRu
Q78VEWqQsfjEZ0q5i1mYt6eXsQbhxwm8qt3jDwRqpsriziTgiQ4fR1F0q5y/ZuGu6SdRwMYT1QPx
sx7ouri8uZPrvF4e+8wAMi1Anok1aN+Ks3Z8UYp0vZq1wLbnKiCxzyaV+FBmm+DxkrPU6Rr6T8Br
IDdbhdSILLuK5vO9PGbs3GOz3mqSOyCmLF+5y4QX8GbvmOjlIuJFiOjYQJEgLXSkuvgR0Y4RF1IO
puWzr4Pel+6X5qZRSIXzqTk4ggEKxq2HVa2ZbxrDf71+ecLU7u3OW2IMrUqCp1C5jpiLzhp/HKx3
zT5VZu96qTLU49jS34YKk0l/aS9r6ZZqhGCNCJqa45+7Xonm11NVwOaWEv1G/pn/yyD5XnKqGwqa
9lof6sri8vkWgP6c/MFVdZfjnPJy53ZT+/9tVVnYU4Pks5oX4dSEfmoafPqjU36KkmNhJIlnWeCb
Ip56LRHvv/+hPGn/cMgI/8pwYc6L67uHkmG9TcBd6PWCCsYfHrXWr9YxyrxyNu/hPrv8+uekTPAT
CaOC+VdsBXymrjwQHYPQNhtEDtC6z7zOE2HNSDgkfUuHsNAWegKvO6UyFtHW2CvJZiV9esfYJlL4
IXx++Lf19pFUvzCnmDUmChuPSEiSX9wSbF5KENJBiU7BpRBIDrIR1f00BFwTX9qKStZfzxKuDYuk
iQwg94/ewT0Nu3g+BE36nXXpgJvV4GfObkYzFN+lK4sXJ2FjhoLZnpo49ptgwIZ8Cv/IykGu4e36
k3IYxF6na/bOfEjE/9+P4GQfC77KJf3JLAIAhR9Bif4vcORbzhE7zIRpz1Eco7oWlZE1MEecOgSy
TkSP77AvZ848B+YIZw1D6HJRWoW33atOg0VlG5CE98RqpkTcae5KnxIo2QHqwr9sO+VIZs+xINA2
DJlUDnEYj6KqpETQdCIj4IrE2+pn/KZZU9nh4B5boP7+K+l/Fqi+2rV2Fe4XFymgG0scwlEgb8Yp
jab02pVnIYdtJWawTUJLPRfDLNCwv1+aSka86FzUhW6XcPVlc/xi0itUtiZrAg6h0U7xTKDkcS+X
oAauFL4dXZY5TJ06T0zjKXg35LtrL/Lm7HE0t4JdOCQ3BZC/TGeMf6T2x51ZUhMO/pPd7086Dw28
4u+4oHVlJntb/ogzi9Uj3or3AkUwLDyikCTsm7soaWPAlxtfeLefMwUBqC1donptL+S96bMI1y9i
UTqO1raq6I+8sqxax7GCaSAfr+fOM7ZtAUm2y21khfXZlanc9hrdD8lWT8OAD4HJiEmf07fLMW0K
1/vgzgLGfeEcuQ2km+Q94FcTNU5YUnIza3Ecf4zel2L5yHdxAxQbmwsYRJrGrTPg7g91tNq+JTl0
EbBJ0sP11mQO5BEydkmvZ6zIRbL7+KiAL9OlBomIZY5Lb2r5ed96zq7qO0fyS+zoijtSIYVntL+8
M/RqLb6jttjrs9R1mvxi3GF4spzObiUekYAfD6TZ6yOGyGW8vdmOq4pxzx4bhw2YuWq7qMg/mEk6
ba2O7pjxlNv+bHBk9xFhNO4R1UFAtfndGGMUz7DVOc+Qa8r9A3MR5HiHKYXfjacvowk6Q1jvvPWC
4hEOKQ4tFsnb5P/wOdh19TSIsia62eUfiOXsHj1rYpeZFTMvdgOsdRJ+w3tWAZktIPM13qtPMYTw
PtZJ4Ht2EdS53J4iiuCmvj+0iUUQPiv4JLYGELbZJeTBMuV9eX5HPYkRHUj4S7vEM0UFEa6c4jy8
l+x9HILogG6jjV6fRl3chuVUzwYaMhfgcTZRBIZab9IipmdqTLIW/pDV+3s9C0uxGxiJBFH4DJT/
hkFHcAzJ4bHx8K+MfVi6nc5QG9+wnAMSQeU475LzzbOdNT2M8r48CczNJHX/G2uOSykjQFUzw5Jt
5D9z5Y87LnVcHZ7GDgNj4+6+dDBMCx0HeJ5KS3/32eUEtiGwKB6tJvWbvgCfprbQv5T9fB5oItgf
bJLVYJzT6QVxZj5hjtzxmD7a6HWEzjHQ7xbzDJdEAB9g2mCDRK+r7rgt7iBEztp45NvaKpGoIwR9
fWV7Sy5qO1mre3hSQz6+LwloAyeVdRxnsc0hm13Hf2YxUBh5rkCQZyCJsmd3iL1OKmPP/CUlLccH
ut1gPva0cxlWXKRLWhfxLThBMVwHhwP/L9tLsttbtzBcpDwLqGr4vHnvdtf19dYjuzFhxez4r9oU
9a9f2r26OpLqMd3mSmeOsgI75ncYZ548jAvYPtZb64fCMd6U8ncxU63NWNm5BKfdRVJB2laiI/Fr
vEftB146cBj+zkUzi4xzA902w9qwLFddG67QJQMcpCLGxiwLx6V6uYwsexcldlQLJ+ScE0w72KG3
5uANBpf9KPcVOxiT1A8kNZ8XJbpwQce0PR7kmEgR7Eoo5H3AxD7KI71WN64Zy2gHy5XxAkwIp2wd
x9cxXXZsTjoEJNkteLTxts/q6D5pr7aEzCCUAS7JMH3Q+weVEW0coJUNMqxYal0WWvxLS1PbbsoT
e2b/9LO81MrD1XXxmFLlWbPVpsqznWpMzkh6M+Bn9W7uVqrnmvvf2P0CoYKBNNPGT34gCC8l4tf2
+EUEYD9Zk99WMV1WL5pHz0eQ+tgY/wMWtYp3Wre9Ja2CX1Odvxwfq/Y9VfgpBGHpibDwdjzDtrKf
6RVuBTSMWWLd2oInjUSYHtHcvfekHjkDacTu81R3EoBH4UnSgNFodbyz+VlJmSeZASoQS4Fufqrc
PzdtdPccQiZ+oswajG11K4Oodp9eRdzGvtHMv78JgDCOu0zDV56ABCjFQSFdy2iPgF9Lc2Oeq/ZZ
iTBGDZS5s9X8Xwk7Aa/VWZdYf11KXf+pes23ZjoLgIeu0yZXliWSOZ6SeNMjkZONROuWCz9lyzD4
/K9zrd7LNoKowq2uQQC8+zGZTKlpmr+hQDDyvXHRfQAxoDxJ0tTWpqvcOKa6X5gB/x0hHWc4oktV
N3RXTTzS5OOZvNzm0uczzMcejk2+hPG8I3BuwtvKHYxCGE8wPLLg8nTIm0mp7XvWCziG9uGYrsIt
AL9Z9NREQ3vkD7IQ4uM64VxgdLNU5SBoomjJxGa4kkk/hck6PYt5GTC99ygqTa82LdeQlugQM2Q3
dgyu2XQF098zQGPXZiU3G9KiRKl/X+RF5K5Nv4DMhb5tngjdPftZwCy3ObN+ZJ5g5MIqhoV3tw27
pA7SoZyWbQKb3RBp4eYvW99gcHMV/1KH0clREhJyGu1VfqrenkQYRMcqdlZTw/sOm6Zq7I1EvZVJ
gj3U98wRAsHC0pwW9/+rkYrnpEqF1ARjUx5kustpF2GXF/uSjV9phgO5MXK2cB3EoLoWLv+sMKkD
ZcxEYzivMZbi4Ao62xdXCXfjCKTdG/hx0NCiy2zsk4RiDQoGsylNfyMYyWHZIiudKl/NCos00gMM
aiIKE+Mt3EHENIWtA0f4s64g7R/bq+xkBrqNVECZk/K8dBzfqYOucjXvoVcDTAc8jXoB6597GUfB
r2EH0akaDaU/NLtzrbRlvf44RhVqh3PDZpYxM9edOlJfbusjJoshUrvXRx7DH2+N/PM0D6nXjo3p
g4u1nI/foRm5I0dGRE24MGq9ivGigi80fjXXklb7HN/+U6tPBcbhVU+lS474Gnmd1xmDYQVYbBwz
+ccxoJV/V/3IxUDW9J4TjN5LgtNxU+RWhjRJeFm4udtmYCJHE9AB3rWPaIbVmInvg0qynS4kU9na
lf+49UYln1Rv+fDWhsbO9GXYTnuCMa1wkSW/ztAPKD1aSj96fWsuSVtD4Ip9igs0hMICZBd9/n0/
BPXXS36aWvr+vGHFfTxaH914e6RD/nwA5xmsuAAmCheh8iqGICFvOFxCdPJx6SlIr2kXbi4ICKOn
ko1RU+uCrWb2qdeoaIXcvWhiWb+ibl0hgoqAPXHJ5gDM+bTyA4gcEFKiX+Vx14ZSxTI3j8CufbR+
jCygS5Q4RCil/EyLLS5Dy2hlPpvKwREBav1G9YL/XgiP1m5krA98PTULHlTBX6DujJGhIKmdkeMN
LZ7/4kdccGPfJ6YqIMn0zlVLpNko5slE09/PQGi1QB9wOcsw
`protect end_protected

