

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
gQ4CxdvWgnieRLRQ2AMwpJaA+X4QUP23A7mcpTzLH1nina2JWDwyro/SbR0koY81VxQ8tVNBYSg8
3s+EjSEjvg==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
gPnHmBrjBHDleV2Jfu7AAgNyinLiMa4GswbueiHBD8y67DvELbF4ryETXsYzyyRC60JDgiQTY9xS
mNBL0n+tguqX8nripcl2WvUcK2rEIU4vEmrY5Xa0k52V9uCE29ruqODz0JXngqZvaosAn7R3hB73
7cI2IgLWPL6sayUHq1M=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
bim7wErRMWV5FSeSCuJLdGVUUYEH+U9HzwEGlgElmMU1LE1rxBL3MWBw6E1Qg5kGmxPZcrNQKg7b
PLZUD5Dv3VyvXW/HR3jI7P5DnwdmPcuCjrrkZwCh4jjzor7rIj0AM8ubprUHwkpicj6rKGNYRGRi
+lmT6hjwlretXlYwE1YClKFDSDei0UBfS9a5tRfCcNpmoCaImXf0uTOJ8unbujREQZSIp1snYBqM
Q6qvNMpDqcLoVSU7OrgHQdnonXWYqY/ILDCjdL1o02B+xcnkuGf+oGCDs8KSCPuzYvirbLqI8N91
feufkvRKEcc9+CQ7U9kVuEQ2Z+MB8XwJtiWwVA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
HhRynIQ+TRImN/1ISEgCruTQGOfZ7yQ0AeSPRr1UgeSXeBV4/j+sqUVwy6KpjxjyOB8/Up1pUaXk
C62p4kvtT61bX2llnNuuYjikfaIxGUWJ2S1a+GpileS7Ui7iwtZy8qreshTy7qb9L+4SycH2S0Vs
ofqZzZCA27OgdUdAA0M=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
RhnO7aE6HcfX9+ngWNOvpaRDGHOLotkXich9kwwYcDEBAwcff538vS/s9YC3iM7OnnDBzfIjK9PG
hZTnV6Wbh+heW3iD6MhhmPxC3a+3h3Xr7G6V/gV+8tP3qbjwLdyiI3Y3Tl9GXzeddtSNdvaD6764
1AS1CtRtG1cyGvfnXyGxmyDzJ91rqIOqSJbBOVjL0a+NolFyEU0BYVthKlZ39r7JI1kVtcM5XAND
LnFrRp5p6iEzVZDFdricPTs3V2FwNDnZSvZ0QADHlENUl1ofRaFRtXOEIahTDRwJJzBMRTba/K/s
3AtKBuzpWzTyvSqo+1PWwgrrClt60fAvHko0Yg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 12608)
`protect data_block
dgz1L3uk9b3RupngcR9NQCEe/fz65+G59UL/KkecdLRfwtvJWQvKa6QoM+AR+6Eka3vsmae6UaMK
Bp4SxCEtzajPrjvf1ZvbkWOqmuAgcJwBDeGAxjIlLubJ7bGIGk8cUxmrZA76WtNVRH+iIHOV6Gdp
8lCEKTOBWxB7MWLVqgdNF5APG+bCLBvyFQexNH6UMC7c44xJpCGrngGdtFmODdN3ITm4w5e/ojNI
Q1DblPDkRAanA6LHQY3NpctgKUxXIf6lTzjPgElqBsZK/tWE7PFbAp8egYEREi2ef5V3N6mBxTKC
feiWd/5c9eaUOPDolIFFjnR80LxlYZLikp2M5IO0O/hWSrzP3klmVoaOPuCtu4ZmRQhO4aDP43bn
FZABBcoGH3qpDHa9UAUuU4YXIIX177nj4sf3dgYmaHIUAUjfma/P2d9ZjfR0SlyH00Si1YovL0cK
OAp71qVCtclebJDczVuQgzHs/1TgxICTUNugwtd29PLy1/pCGrjjk/uL6oed9qJ8wqrTXY2hkvXq
/q0YmxKJdXYza70hRf+zB7iLXNPh3gkwOixWnwkir6bBGhvJlOwf4RI0BrtH3fmh6aFjhMzRflJ7
fSm2rcUZDeeznHPrdrKdyVBUei87EdpD7+n2+AypiHTRwHJBLYpObvkzvLybx5t7c5wZXxb/+0Iu
xKQ4CT/+HEyMH40t5lkvEmrR/NhvFZ7VNYISDeyLMP+7nEdzbNtvwVsyFmGY7G0N0gbO/Q4hyZJJ
1YsY7/PhRiw4R0YwwlnKvJ2toQcu3FA7zTnQY/9dbsCokhQf0hRQU1ZeS/fKECNFGDWod4Fl6FhJ
HqaakiDE7Ua+NVqAorO+Ix7qxbmIHUO0qLdqyq6OIdrQGEMFphd9EZZ0ipIAPmSzBz2QEyitqN+I
Ct29icc0lY4tWiFj1k0xvAyQSDyMNYyxhgUOvzOPMKbSMtyXyI8Oarcxpqns61+9/s/rRfX0mnAq
1t3lbMFxg+BoNBf3ZuKKCaYNNJSaE5Bl+8UhnCTxkaP/ys9EOL4bKQyz/7EwK+MJAGpKdnsomysY
/e3Z7FP2C0dRu7NypzE0q6doa7xoDp+lIiGC6/m7xkgLcezCppt1LfGvmeClFLqwb9rVNTWdGxdv
6jjLm9ptRYhLL3TJUQaPionSPyZfkG32SmBcEglYheUKLNuNXnm11c9YKFzE/o+KF13lVxo0ihrA
2nKHSA4YjXFOqA5h28QRkvDhp+7kvlausspeikdhLdUnFqlIiPCHmt4+G6lZP803jnXx0cHlFwDh
+SPxd/ilXBTkeLtyumVmqu9bepOgzhdaSq36UBTaD2vtgZpuPw6HZ2jZxWRJRWHdFst5sCufURHO
L6pzaL5gxzU4/CG/v9z0UX68BjLEkpPKrXfxZ/YYlaiGYM6l+R0of49GWBaGVtxjx4B/Sl/laBo4
S0ruOyMlEWLP6EbiIpeAr4Whw+qN3a9VPNqlmLXfSAKQ8VZG/ZTiswMshH+d3VVaYUt4GvgpfdSu
FEA6pe8ulRHhEoDcXZ5VV381DFrtxnGsfXvegjeZwVL7OSE9hs0WbapMv6EjVQ0j8btF+acZ0p9b
LkMCI4fV3867aDiiilcG66EhsfC7WzOmOTHxOpYa+PEO4EBa5p0AWQAJTsO2iYoaStUQW0EOM1D1
AEczdBk6hsoG9eDTy+kbgFVUEw1K3Isj9qQfMZWVBr2Zq0X9jLxqFyi+OyIuBhDRLNeOxCFyQb3S
4r2k8Nsn4eWAnces5iMWlUWdNi1elq0Bt5c1gyCUxGXoQbj0QEu8dNFT2DKW1RSXZjK6kSNsIO9/
eBwsjtCOlEVaqbrR5Lf730N356w4/nSXObY17Ai+syoKryh2JG9EcpXgLaLuuzuCmpGnh9eQWS5A
1NIRm35WEAgsf7nc46znsyMoq5EwDyjkRTazQOPEY+cjKYI8vtArlsppdcA0gJwfunqOrfWC1X1d
wKaqX2GUJEYVXj3MdKiB23VeFSQIoGlL2Sr3jjpv5OghAOJ5xiOOov3cmYvONziJ8cnWLBW70/CA
cN4vYzqHmj5EF+/e44QYcdlH7364kUvDjbCtVsJV9OV8pootXu/X3lGwWAQxtOuL3sQOVe8oKsMX
JW7Kq1WeCCxs8YV3LNYB37yqLi9s2VJFTqlp9+0wKa/Za1qY/y049UWq8ZujYgQD+7o5K8+6RQgg
3jMmMrAaJtqnqreoBc6G/H8IpMzCOz1BvElMojB/s9kUfN8C2o7CD6qhrspFN2xp6npNnsXMNOGz
uz+K7PdIS+n0hjBIEMaxtTisVgzpfgtiO+Gl3R2yanQgWHLly2L5ZzflJLq1wavPISsSocAZRIdY
7GVco6ozDHqKBVW7A88D6/z+UN0eKcTT3g+9kEnslJcSqMQmicKfzFdcnk54drn4W+bl6ykd4toN
svwyZIkflh+GaTnBgITSWN5DuIwB9AoLaN/PW+wDdhUPjFG2CJ8eDLkavKxJatENBPtsCJw/2NZc
+tUEXZOji0HejHvWdt3C4aFw7w+ed5XRppRYm8Q7EaN2r0EeLz+8VlH84W8lDdWEvoViKTMJcX91
HpyCEdk/b1OM6VqXyHfXi5oPvGe8uASbgestBBJPxdALLtmCO9XKAywT/ZLq4RXNztjpx9c8UVWa
zTwopDkR2I7u2bJrrr0Xn22d8fP4yBwoLlRvcxKP06LFqym02QtiTjHGbxb4UgiV6zGcBSXLtR16
ZFvBvEAJwiRGq3FBlA3J8dkr4FXI/aGzBOswqdMcJ6gYVtQM8Sr6JJTUWBvExnAS8g9cCKTvUYrT
LBs5FhkpTn4qU+5LFhynBOdtQicfDiCB1L5nkLMoLRhdEAAoVs3IWP3JpFQkvFjOq0Ra7BdrlLCO
QSx1JuaaMc85Mk9jVObFvyRMJFq8nTHlDxyYHWl+/hpXDsYNJJbQ5/C/tYv1bCe0/uXp+FPf2yLi
aGrFtUImBrVmK04E+kmidgYLnAkyAaLg/tBwKZWPqf88nz1ubxvQJPhTws9rbEPg1npJECPO3Ydz
Ur5EInM0VtKMIHKTp8DG+mVLHPfbmtPO1uBdFa8rQ2c57sbHw39uCilnxR5MmmkksVi6PwRs/Ta3
+Jw/7HE7jT1rJHD7SRFt6HqgLo7O38mu1tQHbPv3FREL7kWCtSTulSSU2j9yLf3BCvTXCf2bS8HW
6pVwaPmX+yVU2sFiFLhBUV9iPltntCrDRpf6s3GZXrum1DF5xiBJ3dLRRW2CAVtCGuZZLXZq6sPi
Djnqbgxqpslj/JRAeXuWotu0T/dp85WenQnWhEVf/hJlJIXPdCPWiXrxnQdUrDEQzLd3BSNMDQFd
sgfs7EIdph7+84RC1/SCw2pdsWis9KuzDMdTQH0RUJnDgsSACVvephN5pK3n6su4zsR7JhuyhLPe
zhXTN9HfcpwtOXzH9n6Uoo1CGwxrsBluT3F9PlxTVFh1Y4J9MYKTQ8ilW7MfnE2w6vZyJ3jKdRDO
oVu1h5Pl2NW5X4PWQ9pfe0xAZyEimo4pf805Ft1hfXmXZTEZTmyhe9qNmwwPhrv/vjW5MHDaQqoN
hnLB7RT0ycWMYCd42fEcLhLBLIQFuzTYQ2wn41eCw7l3bo1pEHsnAqNeifr8CWnAV3HP9CNs8Kh9
rZJ4U+mKisq8lMtbaHr17ZZaAk0YqUPcUA/56DM2h614jIf6O2OOj+nDN1WQQDCrvj5U4u8AXBJx
RzO7FZ0oZoD9it2FGM80nYU1mOf65Qu/9U/DnUc7+6IdtD0+vaurP0n2kE3GDT4Oqq0wwm2gIoo6
Lfi2Rtp/wX1bw/1h2aRyxV1kw5lTOnvMXS7UCoVOeBmHBPS+U1vuMiKMgOLlFB7fCxioqaYAJ04G
5MCa1syEGB+XR0dklM+VSdaTQP1yk78osSYWG6NP3wKiukCR+VfCXTMldUjLRcHGA/AgSnTPZyC/
5LVQnOU27UItNHq8UO/7wVV6Os2PkQmdtBkXiLQwouQiCtvj6q0EM5L2urzbkBFx598MBxE2t2O0
38Qam0GIcvNVNX67gk3kSVYmoQ6GDubr+XGVY/AL1Prvtb1XIfMXGwgIodClSE4BdN2nQhcn92ID
2G3T8xwfyMINMtvcUKLgyYHdsGq9HNTiusumnmVRk1PM/dYvPrcfUyotfxpJE/mu9VqYRufRNl3a
r/McJA9UxF8tveHg/kZo/EToF8I/JXWXMIK1UqAxTxhFd2k4uv791iZwes9jJiIexh/narpN6ZkK
16GaX/lF++JVAfTDVzRGEZgoYNOzBLSoPtEEM3Qt6zI4RrEAqWfS0CUgkZZ3VfGUo93y5ZQ6MDPk
aE9HNFGGTygToxd+2peR13sUmb1YlRhHJK/g7W242FMYzfThIlIFG/8Y2slnV5d8QLT5TK6IPcGS
nthX+8I/dEWmExvjWgLOqmOjopQTrPXb6dSfrWx/eJEiTG/Swai9L0UKADz8+7gtkT/IMYMWDJDw
4+MxFMmyUy8jJQLMs62fekjtUgHZhB3MfAH5HAYTJLzn+JWKIUxRqaPcPy+AHkCzciCEAqh54arX
XrjwxWs8vMqUhmBzK5rjJUz6m92DStlb5UtQOnThaMArnMP+9OsB+JCGj9MirahUeGubHzr9Prow
p+Buq/xxtPk2WS+BNZEcHlb8nZX/yCYKqPoLy9ebHteC7/rYi0YHs1YPShOYF+RNNtQ2IqvWZrdY
Lfjy9HOJgTkEmLTHV/yUe0TDucdJsMw24Ed/uItSHyAYLe/E/a9d0o/aHOamNR7c5zuPGczBZ3MS
cxzTB0v1T9PZB5DhZSYGzsU5oFuPjri1ayhjRYdA+scw3+qq0njADQMCbB1pwUC/VoHFN97tEuj0
i9CJVrzc1sasJJZzc5gWT9Dq6zNoTHH6ml9Lp7evDzlUj4u28oM3KA9ANIT86NxoW//mtRmO6aQs
pex0p5ig5BN+LTT0Jzp0nSOvOLs9Pz6uFHou/lXd7Y1OgjJKR9uqOSkhCahYVa/BgyOgqb6PM48w
Zg9Osedaa7cZur2m3hdQCAcUuXR+75gH27Y/FM1wPRck3KGObn2tk899bkLi+KYbnvqBtWLFziS/
oXx/nnyIArIWSxbjeuU93j96UfJbkBwZqP8MZ2sIpuHanbNx8dmlqRylmz/FP2mRXzAdHdgdEHyG
5+hlNce1vDP+5W3XN1ynG6B0p6YHY6zE8OwCU6yS0SqWKiEHwpEX9hG+Q6z9fifz7KYIMw8a1Kt7
VBbNHpXLmmCIUbwNcFWpjaAydw0IKopTbiHOHM4fSZarJoJkRJZM8A+WD60o4BRBoV4BbYoPfCn7
JQ5wD1/fRbbklZLNvd+X4BjwnpzSi/u5XLQGgPkCt1jaE/U53T6Xlmk/OkL/L2nEJXDfnZRsHn+Z
/8A9rAofLJGWXH2H7hWIyz8fQB+2vrQ22yORNMpnJkplXg3nF4tDC93Q4a/vnR64w7xI8L8bExaf
7BV8GLH+jlywOSmqmmGfQ6VibJGJrwz5WfBQIesD3zopw1LD241tbAfSbfKtvzSIevBIn1bqpCVD
wRoX9nQjjyetWS5M6gQtTxbnqQMbMBfe13FOgZKddGV+QkGFuyLiH8aLOegFW9+xd2iBKeZygrJq
ym+oAErj83+neNfecNZCNY7Mf37yD0dYXleSz9hIGusM7VIoays4ypMkUcGufZZUUvXs7Hyq1yoG
4vc9/FbdDTu/YouIu/dRs6ymT3JiNpYTO9C83AZnxfWTISPW+q4gVrixPmKNyfLYBM49PtyD0No5
yaROJO8/Td9XBO0l+QRA8uqf8foENVWGE49IOkhZuz6dR4rXtYtf4Kd1UwP8qGxkojPIBuvjtA1+
zq7eQzkAPtKd4APIAuLfBy6OelL8LVNZvfOj7N6PNAy2Hy6M8CIyZ0PF9f7b7cuiuJcJ7lg03De5
MNjJeJjObGIFQ7q7xXDBKEi7uxB66b3Ho64ixe4Thwbjn+NhupKYqipHPVeNFHs0f2rZtcz5Lf5p
j77tfwjDQESWHFf1nhaVHCc8Wi2rxd/yuiQjMiSMrKDfOSKTB7pkhSyc8cZnqLtbUnMiOivZ0NvC
j2jMCzrV2sfPKRWKgJCInVMYe1eLuL/MnOgrI6XUsc9bF6iUSBsyuQjRusg2BQbNMzvs9BjPm8h2
4McMXx/NfW/nTBwWQamIwwKHgNDXrvpgm5gFwDyDkd8jnNzDGptXAvBjIYQ5yII0NDUwOIUWsggU
/qewskGicR2X7682/JnvXRsan3h+55dyzMin1rnOoNe3GRZtQnlhR5Xnpj9mAv7zP0F5n1bTteN8
Xnz/o3qiqt5fMQ3jE/l4d5MRGE4pHwetOQ6iZS4pFCoL08s82j2V1JI17hD0+u/ZE2HIAV/Fm+0d
6Whk6kK7sK2GeODU5x5QDMG4U6Ah9cGByf6iCV5db+MDWX3sU00MxVuIsL+ZgBcNxOheOx8RECVR
83oYgzTmqk8AMstssaLimkB5rRyIAWJL8Wlw2i6tXepenfAwx5Si+WOKEQezXsoZVhJTdK3ztn3D
7PB6xaerq3MvU5NvT2+p9sqX7DuSBgg89WDQoeZU99gcvOGNJAuEx8kymTtToM8jzeFmyDB4PBjr
ENNcqBOR9ZjSLke3cmlbdlttYFfVa6Tra5ca3u0QSRp7bhEEugipBspZLnuSa26z2VGFgG4uYwQ+
VlX7KMstXPKAOjL70yfpi8kem0H+NaGCzpg0HfHbgUH0Ik/RwgN+8BYBRxp/ioJB74MgY39XpgSa
uXsTCT2ssAus745K302yHH+dCPlna1eJ4xMeVqWvCG/zgmrJjXYpf3JF8KbFapFoHRbQcDkJHUOW
CiaumN7VuAH/KhY1Ip4nKdi9PZWPT1ALLktTjEjdkdcAr6snrOEHZtPGmNrabTeeeJ/QpcSLO+Fk
PoBvviZvWFSJ1nADz7xKN0tqiy9WuDHZkhfNJ0clZI5J7gx++sf8S3+fsYop+ZujYpAbfoxYkCL+
SN2wH7pnl4El0Ff0GrstBZEtF1LFbpRxZYYv7PuFWOi+gVF/RRIHSipfyVtq+rMEtS49/dat1wx+
rRaCc+J7z0NJpteH2mtNJ4lPMjwpcx+8J+BNJpt+nFXiarn5HY9VLrFCsr2LqA/okJ8xAEqZt9I2
cVRb+Vvxuv+fXsRcWbm2srzDuMTgQXxN7xQmnybd2IrbjU8z4pYBRp9Uc8z+6VJIxmxeUmaRtA45
zfPnVG5z6qiuRHpV7Sjby40A7cSkD+oS9wSkyZqUd/+UEETR1LRwWa1WGXDf117ty/msoyW5pyub
3uIX60WhddWTrrGtGfGTa+HHdCJ+oAA4zlG9MUlKqL6mIN4qoMnN0s7qsvblEUE9A305DAH7XyJu
EcEE01woDzC4FiXMKf9R+xwqcqGnub1AXBN+GXYOX0NW2DykkpvOWzKHNgHq63Mb7sI9wqcy3YcQ
dL4AZRQEWGhGn7x9gTp6r/c80FErXT/33pCgpN7c1NEu+vQi9Igee/8MU5hwKHExtoYo6KHOaxGv
JB7NdyanmGBHEd6Mg4P4IKqqWlatrr4x40mNLcVpO7tmrKCkLVTNgdw2mBoet1QKAZDIJniQVrIF
tq0rX1JoMJKmHLNedl12t2v2jHkwL+CBcH5Q4EODAlmlBcY7iVPmaHxocdI7VEbzzpPRaSVYBXdj
1OMz/oLZe4vA60S9deiNfYQws5TZWtjLzfJ7JKvvfvRdSaVedn31ayyxTDSBkuSDoPJNTHGae/Ku
+HqCSYEfdekdiUNfNv0ZyZJrPAyDOgDndZG/tNKW8uXC9rBZxeb7PSymmh1xlki7dlhRcMIYZK8k
NFVPV0xZGSub7mJqGI1nhDD1de1WNBGHnU1xA7VUAZOsv4IePJrabc5UMUhQhzgzDjTVlsJsDXzb
7znkUQ/OCuH0hFhKGsPjmj983KBTnFhnv1tda1dfg0TB+Hp9jkZ9+zA3v7+A9UT4WJ7CK+KOsIk5
njjA8tVf/NuzPMiuCFXqYTS16lSCx9GYmEk/uJihlznQYffeboo5PShBMwEeH5VMFswxksQlbXZL
zSf+M9zew+SfDvw/+yFen3PI9zDzingkCyXVJHsJ+9p/GQxOMnrP6jjIHrk+ldHo6HVRetkJrA4P
8l9x7ko2BJKOMSYwyxCaqtRzFTUMXuoSNBuIzk00G/kXS2XcUSZAskT/ECejtKjVmRCRfG7pc+z9
DbLgbyJbUo3APdUuJb/GrckB9EZORVnFYwhCKDpfG8Irl1/Ge9GAzFOTAkGhcpNHZQQe2IvIGr92
XBhL6SEtARePw1l7Ab85B4UJv7UtN9mB1FIsjfBD4Ky7iAERUPz+fUTTCqdlU9V/PHBStSUZiubc
3hKJyzTPaO7Bqx4J0yW8oXOCBYBfdzPnVw3KkiSyz/L4fYNMpComdBjC8AlBNxS/+RhAlD+LrEQY
iLibbr6aE/wJXFiRANWtp428V9w4Extfn5sdR7pBVbyhjc5LfNbmd0owoJiInrE5qaG4gYkPiEmJ
VDSDCml4wX/ue8a7hgjMgB3aVInXFKqnVGM5tINiee0uyFzMsXoUHcrb2JHNF0STp5EpLLIw8ZdW
ZXoGX1vOWwOgRi9czCoL94QSM65/35pKZlWWq1mZYu6mAn6Z7mpRSx8IE9xYjzj9cc3fi0hMPFqO
kLnxcIWmIg/m598c7T8tQw1T+o8iQ1n25n+FQfS3zl1nj5FJG0jCrkyZEV+O1zspMmnAi2Yur9Sa
aNOgP2nyAxe52BUyklMfYp2810PqklwDyY+DF09+ks+upauhkLwqai6Ep2P6HHBKLmBg9jSj1qBs
ht1iHXWnbJjjZCRuJiJhbSzUjkYUzJZpsutolsEpiIAyNpnurq+MemwbUCw9DhmTiqnYUc4dyfEt
f2tqc00TZM5E1WilQ0mrk+4G+PVV6s9DHofUP0+/SzbkelDiyMxd3vtPsCFzCciznMYYqIhzyW4l
1fxlXCcHNIkcEfC1lx65ccUVgn3G55fcdiHxwN+wmJLEoIIbJtDFoDiuWXJVGzh0sPfQgcncKtzs
koRTFbaql31677fPs9ssYGgExs6MXh0QJGEuwHJnNNhfZMgwu31H2cgX0N1yQhYS6lE0PdbrUiaL
nGs2HWglNsaV77YspHnR05M+6RxG4uAWnigWPMKgBfoJIoYNaiq4pH7cIuYzD5G0jFcbdlung3y1
VpR9jgkFH+b9oCk5m4Ce7e+Z8r5VbS6sNDaKCC3gv81E/7LUS5LwN8K3gkFViYaeaNoYdaBhFTLb
9ApiRY8b9wdMBNUcdaOIBwrvw19m2r7iFO56a0SHVuCfumJawJ36ezZdJLAGKOcbQ8mXttTS0SQY
jmfNOQnJFojRv0Ba/IDEnKS4NKAcBRKuku7hvImMXk9khbfWXFQyKn968EY9THvmUfd6sfeLMQZd
xOf8ZJRbwBo0qysjczm0R13FYtB9lJsyuFmWtbCcHkQlh6V4/9H7CBBnzne9dJlt/9GFOVom1PM+
vB4EgBZ4yeh9xu9ak3nKKauyPS46vlFZS5SnCFbIrDNMF4CL1BrlOlmrh0SLaW+JkgZYAMOVCFLF
Fu1qZZfq/t9Yrqua4YR6M/DmTszzBSX4c71dowuEpBhv2OvvHhQCcK4M5F+weTqPLEtW6zmLLcVQ
hJE8NgSo/B8r0cT97zRxKLmLaOulGnEIgY/n0i3vpzLwKYws+1FbWpdM52/qP9oGwiKB6Fa4uIYI
7u400pZ3Jr/i7lALCVGB8z8JaIb+OhSrLgM49Fx6jyUV2AhYOAuOEjyBgB1/FsMCo0UBcG8kbb4L
Q8rvtfBnzRWGnPWQ0qZygZizbKd/SBj79u/GoKICtLQRF7zF4uujs4NQ4PHH1mYaJYqbpPtTFQ2+
gLZiEPDow+zK+09JLW/Xcg3/wabHWVSJb9Hnng2tFwRoO0UsEANDT40fIS6R/qAbk4mz0YduL5JI
WPJz1jpmbCz3ItEUCwAK0F5+KwYYdPBl0rG1sy4L8/qosRYdloK0kZvcR5sdbdEWXnn7HXSTB0LR
NAw8jLpFPueJkwfTqj5wcOQzh7lPJPLj6EVJ08cCxUvDyNjoLdm0L58+pidIkpSMH5k9vhALdvE8
Ly3sFgoTApTEOVuZFiBBlWQI+bEA5hj81OsdV7oguiXzJIpPGjyPm4qvUSkHHqMkMTJEF8yoksVx
mFOLOwwOtHRiMNxmF4F3wt7St6OUDtN6i/6RO9c2+5QplbSPFtQxdFiFuzYxYe+mdE6iaAWOEMsI
tAAbTcAZo9XczV50WYeQG0JF6PEsIXvNH7nbhWEYeTZhLBv08XT2/M1zRHNHVAJ1QvNG+5mRbghq
kIacxNhXLfSFef4trqdA+esH6h5XrNaHUeb0AFa0A7GGZI2VWzjOxD+TNmA0wvcZFityeKyhc2ey
hT20WeL6v+zIfa9RRJevbZQZxjiiHTEY1j8remNVIHgEBHxRDrdXcTEyZe6mm7wCzGV9x6pmrtnS
af+5QmfVhXIwr9OWEoJHl1blrCXMTypUVI4MN3lUeeFwVuS06iEcOeVgHen7qiz2KWw2tcok4LQu
Lp3muKbPWsazMjPb4m6QdwISxhW5mxnIVWB62wUowROGth9zNd5PTQQVFPHADtTk1tdxUvi+sV2W
3u8GpWqoLDcfyK7EZ8QBByBMeVGfPVWgYTUwBK6bKkhFoECR0HyoZe6GKZUBzt8ctaABV+Id9vv1
KFUIKIs0SbBM/3oz3AllII9ev5YUsLm2CnEkIzWwAa8KmbBnwThUBBLH4naneHZFiDUrXnMOelbj
WrrWiN0Ev/85i4vqKxoGfoocxV+69zhN0rYLBSvxovY+7jcaGAI2C5u8GjES8a38bjG69iJMbztg
ndJzjSpNR//qQEaWNOvMEGTJYfWZPAu5pqgeAybq3iWnrMYtpcpBeHcfC9rIzV2gZQ9iYBvTrtou
Nb4h7FDLFHvOTNBeIpi2mMD1/0ktVYfhPOuvkH7c/Si7CqdBLfdNbvR4OUDFhAUgxeInd1e/aCNi
2EHVfDrQZw/moYM3hf5u8o2GRdY17G+L/gYfw4zFbDh0lVpY11IqRHp1kL0xaQ9hajlDmFb2SNeI
PbCdiV9gLkUsM9H+qUvUSdDRJ6aIBXZmjyv6P9el44zL6N/6n6Dd4ZUq453TL51WcMtasxmIhZQl
KN1ZJUmsQl9rWxyyuChR7KULlHPsIcctviWK2zdfeyaottrxGwGncxvzZoXvI2N7K9s0jEgh33Ry
cGK2woCp6RDKz7kw8damjvzZJ8cV+i9t/m1P3FdeRSk1BE4I8zCoVM7tdJexHMGHW5vFEx+Oc/FV
N1skyQHBTQTQa6M12sMpZjLX8J5ih915EamhxlIC05fbm2nGYE3deWZgqdTmbljPBtA97n/o8Yg9
BJAA6FIEF656pKTL6YPFanAvr0aMghHdgMOaB1cVvGJPSFLgpSLoUmkYCJVpEbsE7esyWvbx2rVc
dOBzmMcQyPbt+uMqJSXQoFYOHNDwBU4a/9ZgSlvzqodDKSKDjvIpYOJ6+P4bcldMogTc7w5AfvAD
1j4hO0L7S3fsZLZYxh70HNSUsZMWyGDyb4A41w/f+/7WJYua3Gf2xLN7LC/9z4p07oSV8n8PQ2C9
hIvBLvX/9X26iTJJq1AS9shfJuVoC3P8h4WUkJ3ZYSWi8+qvDW7r4L/d4D2qM191gI/aLNX75Vuq
rFi1dVI85U6hKHd7AiBiwgh7R1EfZ9f6nyePcTo1NY1z6XB6dy3YELhVuwW06sUa64U+gqgm1exq
SwbYH2MNTQQIUbJ/re9iRXLkCb43dSfL8XzSJSsnuXkfSk/5dcetLjQsMCl1BScv3SQsZUbpq+bg
NWoaA5xxpERTE2V2TF5ApP0eVPf3BAJM1eOrrsLLSKNefZeZxXqiWF+buWWKSWRuZJX+PBsSGLfr
cFg4Ep6LY7wmATvpREpjSOiSh2FQJLvWR5e+6zN5Tr7h4f/V8kKC8Sxzqxrc64Evz0IJ+XLU/NcY
1e0k4sBiYqq7vv/jC0HZJ1Oiy+BvcHHp2T+hoL7QdF1jmzifUbLtkjWt6czO6O75mJ8ihsSv5CNO
3P+ISL+X6ABvADVSmMeMOgbeRrTVZwiNcyWqvzwdwI5gsCeBNYujJalAZ5WgON/vOIwQgX/VWdCG
+WMfhJrOLFoy9u8f0gcxysvPVpJiV2ng6e3PjqpLMuAJTyZH0l0mtxCKCbvbrwtZpEV2bInCBk17
1MIqDIZYsCT+skGc0oWxg2p203FrbsMx8wXIdDgIm+siY+Rq89N+K/9mRonz9+3kNWAkfaqWEldP
U4GNWqW3cmYzXbePS0zjsV8mtl0GdxeO4x2jG7Zg54zt1mnzBtqOVW/EsBy3Jb+fcs6p4Yf/O84U
sTWcWG+4Wb8KVhI5jZs2zVKFv+m/CpLGRYVivqKj4k1QrbM/Aw9wLWSjKU1rPH4BspS3OBZioU6z
IFQ7eLCiOUwTAv41yJebNyhqsSj8X9tkd9YJ5qXTZ6kQFnwl0qytaWBndgU6t0aO8TRiTxyhzbbc
8cjlr+QGyEgS4E/vBkBG1Q4DfW04+1qLNqqXqXxFggDliGnjsCGAKiMou3GCwUh0+FaDkFFK0/nO
0evJX3moaIa8AsyYejHOliyBb6XA4Sj7cLKw0qiYq7KY1uB2Uv0NrB9MexDBJwPnwY0F4ZhLoY5q
PiJc2Qwgm7ik9MikyPpE2DRBO5PDOSsUtkGJI6YOY4wfu5lTVJbw/5VMEkb1Dzg95YqZEQStl7Lx
TNH7z+03okQsmp/wusmSsRbPi+PcRhqeDG3pJMNK/F31xrVg35lVuPbZiJrPFkP9IQdGdduplyRa
djJIU/A617PvVzGoaoHXZ5F7mNLxBFMnlR1hLP0/4560SueBJWMeDr5DXTCtplra/V6MMpKGcVi2
yXCynK5cRKwVpi4Uple8c4l67ijGKwZtbEOA/2/Z3okjmu7NjMu5O1uo8E/keA8vhGQPFHfnhhMp
g7J5DFbXqGTI8gXKkI1y4Hpge6fh/xMEoclJtnjdho16qe05h7Lzhrk1OAND78/DW1r7l8RbI/RO
OM2E2XjrZgUGDjhdXkZ6lWf3M2LH2fyqX0aywgHZrsfq4SiSC1SE3B3PW5NXV+Bcebs9g32LWImo
5d5F7mRpoRtxM7DCiHrSVK2wUFoPBKAHC2SfxF8qr/9WDKGcP1GsslsyLnLY04wlaE+RFjDg31yL
Tdr5wM9PgJLzb3OQK+lReg81+xlNVr71cGgcaEz6aDGnfvtCN6W/dLNqmnltHXG0Yz8k7LbmH/Ge
BMEL4ORS3H/hHTDmZzVOf36Q94Xekm+l+1J1gs9fV0ht9LRqsL0f4nu0W9r3+XbUPjTMxnWGXEPL
BFAMQw4UQUwIJ1nRfFYYk2eL0N+mhmQwNSocE67Ile8fcbD7UlQZ3p02MJiiTVqg4rFFzINJ9Wvk
5kFukN7TWkpcIqyUI5tfwxw8JOGM+S/I41HgvTNwg2pAFR8HviDxn9B0rN79QzJUu6+S81nNsC0i
tXlJETlKRPmU6Cg39YqyxKBwpD/M9AE7N79wQ7aFU82egjKdur/+9YM9hXsnvchX1AODyD1iCV0A
FdASczR9Xq1f5rLa0pwtCU5c8Y5eog66pWUVk10xUDglUSEf1bgvO9fvZbYN5zTsdJEliuf4TpWW
IKGpB75Xbfb5v6AKLheRrcYSGcYLaG4k4xHsr0aqmk0uynysGIFXJBMa7QAZgO5lvIY3l9BdJ2A6
Rx9Z3dBQCejpoa+EKyA2B1LdoNU59T1Nejvs0HAjJlbhJGf9FaXQ+/bzKk7tuD5PeJ6z6kjYeqVo
Ag/q4KB7MORVmtG5fbaxU5sTUa4SL8z7lmL9Oc4A9ba14TyihHHcBWj1SHbDHGbfxk2WhYgm/SUB
WuW+1ZclmzmK9V5xCeSe7GapXjEqY2H+AYYEsjLblrGi4FNuOHB0U+ejeYKmWO+BK3XRkO52x6IV
sEikjoice2u1QdzqBmvq2Hb6x88oxegkQ1v0hAMDsvasizzgK8/7n3UBGaEe4nLBlCuXO9ShlJb8
Q5NGDEp8IMgwh8NLjzGvR8BsLSF1j5KglpD5i35iq+xGRxrs9ws90ieov9i7cpTWPgJcPGBqIaml
JOftgmX3Rj5BjrhrziBXxblR62n8VVoVf5dVtNrrWfrWtAdjdMDYKXgUK76Huryc4jjFzYYKrqhU
7iJ8IzzLtWwZY8cqYkGifV8ECfIz/o89ljNtRYTULcVkLKMjVGlMshxRSioWQEDPAFqTrGoQqwJS
vmLr7dUckWqUuW9cSOFG+5uH2faOYgBKTkEvdniwps2ReetGE5FHVhrExnoAugPFJrVxevYUdVy1
NcyYKBTDIN1UcQL7xyi+RhOLHGVA8+anm1vkZpQ7QgQ6qZwFTwcTEEMsD95/UixIz289tOIfmKv6
qjJv3zLQvcoYa1kxJMXovh9NRMuETSDiBRxfQsty/qFmYR9LIy+mcOrJtjzALgwnmjYNOMoFxK16
ypgvSgYU9HF6g+VCEM1keZ7f/G+C7pqHyrTgs2zXNRAqq4G1Vr8EtuP02XFuwIKOStvwIo56bQ+Y
FOuf6+kLNbbdt4SiVhYxv8XmkwLJvcCLwGSCEK2IVC3RVmP6dElyk2nocUTRkxZDqCrz+iYA/8hD
FytuTOARDbH71Abk6xuUJpcWaCW7pDltVLSkLi/pINhsajJBf1F6YBy+S23h4tBZrbBpNo4UIEak
++UGMxLuPWGoirP0tKkeESMRxU6yhCAVqWM9LsTfGbaToE/jkCCZjsWIkX9Gbj8dKsnQBaBO4mTH
kyISHHwnke2P2zuWCrY8AwurYDl3KUKG5sh217zJiz59TQn71zI1ye1PSHLX3Ts0n7voz5jFaKXh
Zn3zCUF8/Bvm81ryqOlRviRwenPc0t1oWUFnywKeYsVbnnHlKKMV36HzsFKozqRocbB4UPsxqSe5
UvqfsJ3QKAyHHNdFV288h47LcntlrNlw4KXDDyC4+Ogdg+Em86R6i2+wpzQSRJlgLEKk7yOUIW+0
J2D8dyyNW/Sh7COHdgHSyYc3SUGjYvRtGXw14329qjGdU2j/yszZAj2DjWzbzoHJhjk3dkLj5Mu2
n+LOHbKj0d6S4c35+CQudZR28Oaex+Mhro8aJjyN9IIKOMpr4rVLTfzo1ix33s0LUUMkKQoj6tPZ
507tXMiwGAqT1meS9edbgDJ2FBkQBorg4/kkhNWZY+TjXfyBoaOyak9qMPXYYtAS0PdHtTnu7VI2
db+fdHgrajTvwIvRiKnjqdKs6dG5TWNnlfOjlDf66MJzdGcybdWaIOpBt0IQg0V1Oju59mxbrhJk
O5pEYbJmnqwNqm/LzFka5UmNjq7JVbDTjtISCiwIQtCZUhIexG0A2BOBynOGhaj9Zhq8LNADNa3T
4Ut8MO6/D/y/v/lgVTGMYhmXgIocoXxTUyoH5W+pi8Xa8oN+GblIZtr6P2ykzH82qm48r0kDA43t
xOCPcznotvTN+Anez4eMkcT5GNEkL88TTFSL7lCZlVR53hAazAQE5EQ335DSv87/SeMBk4IXqrRr
1LTx4RzThDfFKFBOBmMyl+Gwnq6udOc5mgWtUHDjpcvbm1d3k9ey+LiwzBPCD3P3tf1UH/3R1UuQ
3yQ4uG4IAHp1KF2PbASLmYVrNiEW6sDPpDmf5k0Vm5sRUhJ5h67CBntpB/u+WZJ8sDdybcFynS40
srQge6+854M6/ZoOigGAL16Hc3lCB2Z61myReqbcK77ztf1yHjF+uSGHO/i9NFQbhbgMW3E5dygT
S9QpRI2oSfbT9P3dF+LxwwSb/dZey74ytyuRcYnSZOhPJZyuyH9qdpKgIRH3McwOV/8AFrlV7rgJ
qlFEoVuw703Vs1EHweGnYjoa7piCtGVLxB64nyGe3QeQUnZqV0yjO71mjcdgvRKxYeNm0n72Bx47
1A6nJq6r8AuQVRgEXPXfPLfGX7b2I7Nd8xAnoMgz7FYUY51qPxL0hLGEEuTLLBNv9ZMJrReMvNOB
mqAQht9Dv3fi8Lo5qH+31q5GE/rEjQV3B9T6npBL7QFAmlTUfqoiaHKxpTxaYBoKeHlj8BtEZLlM
PUBNRvkYATBmcjSD1Cnv5DIREV+21lLhDgNme4eyQi2XjmR4VyStidsUU9E6cdd1HgAAL/3QYLui
O61Yg7uNB0wNigb0TcNajWo9j+HfFMl+MRxmK8WPuZa/nYYvSnObBAw89EaWqdOqSrWi88TCIMKP
ev8nYONUQcKyVpbdeU7b8+P33JABy52jHP0z0Td9OxRkO5Hm5bJbyi6sGPyaxHeGwClJG1b5JC1h
DKixmPnqLIQoPm9bWt0doTqTWBUHDjT9kdyUSBxUSgeEJDa3FWjphpJTIb5XTJ/rCjoM8eeIhV8S
jKFaY4QLp4d6jFM4AR9wGTfjYxTfgzolXWqyEYtBmYoZnjcvKnjZvmWyRDuadt6n9BxpyFVJHhNT
OK1gV4GtlYhHKwhOcCQJeFWHkUp/LGkOYJEZj34GsDRTLCK5trELn7t7V9VBpr96fEHT87wJniim
8DirUEsu1D3FgJKrGoyUX+ficuGO4SqlxrSfXWIbdmPxfUSU8WehwwOMVHuriMMAFPHgv3ltzQNj
iVEZPgesiW5/nvLravFxYUT/TRr66oZg/NZYBjh+Po4xtnpfw4O6otVnw8GiBt6DL0fFQp2dFywS
QDRuIHrB8sF++ERI7XN+SPxBcxGLc3LXcE9bfULUSwmbUynpkG/XwAbtDgoUojXnHMdNt0FFXEWL
+mmkiG7lmubyjUw=
`protect end_protected

