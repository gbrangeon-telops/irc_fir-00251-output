

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
dwCKj5yWv0+IePBqJHT08eVU+DwkTeU5oOrKTCm5D5dLE5fjKonyT8s7ehOuYqmaU7hbrj8cK+dG
v6Hkf9vaEw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ofPimz6qWDPfdZmLTvO15AJD3qAYPdAcnxW7u3A5HKCVeJi1plo2JwW0CBkFgjSMPqG4mB4Hkwjh
aser6hfQcfNXvJ3JUWr5ZS6ezr5tSrAVnAOcpabYJ2vlFEce3rPTiHxnx3vwSLvA9frZJO+K8rqA
zTaVjBo7aLNhP54LcX8=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
xVx1mMvfUwlXTa88EF8IX42tnG0cXSGFt8ROQqT5GxjYzkciIVjF2lg5N/iujDWrU+m+Hq1jVN/S
7L9ZrnRgKz1GFQOxHGVlrNSRcf8Ej88lKuK02N1SzF4b1/VUH6ht92N2p/ROW4dBYnWVBpIxhF08
xg1QHd1cs9lodA6VBrB5Eo1G6aluz2m9EBGHigHdWN9RnmtH4Lso1/y7QElbZq3E4/diAxIYh9aF
1JcFvli+iX9S3ENdEluRyVweVryo5jTYqJabkRWFuo9iOs/Ic616lgSVONZ4NUl4ItIqkTq/gP0J
z13d7iJ5zyP7sku49PKKDfaHMGhWx7ug9eg68A==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
mm3ysnbGmWPGigjf3cW3nqCJ7td02DMWAwGM3y8Ir0JjWwms2hUSloczYrXXwus0KFJrOvbcp8EI
afa1rxF5AlIKiPd5moyH7qLa6s40f+FTseHQnAhUIfuaGWVSTafXnP1rMlydXotX0OgXaf8ss8Rn
aesy7+qw+4loCzosrzM=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
quGvQtw6SKSqCyA6Sp/eeM9Ow8TS12WLAPu5jebLdqM/ryW0A17A8N0thkaJZco15r7Owh4nFU5l
KZcrcDhvn1UKmGv+3eWd84UW4QDpY80dJTTq1XGSt54iFPTL0Mo21C1hbrKXm36H71Xi6xWsaAlk
nLsOCKMEHsujeF1naPb1xFZWSlnfCp9K2SB7wEzz8xUdktOS4rqm8CvHN3HMePG4N3SsN68l6nRq
sed/9GKEvYzA04tbQb5NASiphn6udoZq4W1cZDMS1xzdJ8v00rtDdh9Iinn05spY0CrdzbMqalEN
NkRAqp28PSG9/FiSfEP/QtuVq+XzCkevSe/NZA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 83872)
`protect data_block
An4KFWB3oFHRrCHvjfEBwgTXHw3e23vbg6Tzo8HzsdVTjdV+Qm+A7A+1EZzw+/MbKhLkGDUe2m9m
XefmofeoPFIfBWEpy2pnDRJqCGjIbNBvSt76YqhPAJ1eY550vD5Yy257imTknizTjtLCHjKiVW3E
Cgz6IcWHAVnAKmmd7z+WZX301wkB7TgWsxkPC8XniBRVK+zRvuncJYrDGSD4Snfh7XUwH3g+x3SW
u9BMeghZHmsYlTOwfanAlTV+kLyZqKZFublEiQEurLEnCuRgU7h+0RPrKtybsbz6CePhnSJ6NLyR
wmCo0XIRgSxMlgG5WbLyA7X2Y9W+ofsl3nAqwfA89tK7fzM9Y3u6AeAnH0/ZHLEVmyQ1LR9fzdZc
Z19CuHKPhfYAaYkbSybK6MgoCsRT+4GY75zeJWggtCiNKQy11/6s8KCi6vxiUqkDfQsyPCpMPRrf
kTyC/0yUPTPEJzKTGRG/m+EVRvO979Ti1K3V4Mh5lK0CDJQqwtK0v38hak+/VxXiLiZ13z0WYcDf
MutKx3wmMbRcAf4+2cOCa/cSE/m/S3b2LBLDogjoGV9opXQI/TdjETYHvRenukWOX4ROeJnYFAP+
hQUpKLBNtgt5e2eYXqOkKnqdmJsNNnk0Z73tGj9K/6cYz8TlUPGhzWWmYokZComct5ugdFw9Plv4
EQe83zAJ4EcIrcXT0Efi9Zak+B53BkDFddf9YeNwKzalVMYGpeO+vbVHrHksIB5Sany0D0i8APKw
THpiJ9z9KDgwTpYdtZQMrvoyRyfWYkIk6+riDtJjOHUuogJDuMb7CH6SqqRnfzoJYqHqz2oYGeVB
O3PVp2l2NaRrRulyKdZ0dPp3I/WT3OOxenpzEdUIs44bWchrP3Sz0feAGJhUavuhQHlx3+9vMNQI
uuXg5OQq/gAhYhfUfzKSDI5WOUFu7N4d+N7Z10TLr1Dh0xxF43ORAr7FjaGgsXCCECuBh4knf4Gx
EFLGhzYuKFx90DrinrEnbCYF27dSY9ga5dE164SV+2yoIdYu7z2WiFtvBQl9jdmuX1kAy6eFrpMC
hADymEN6RufvsX1d4CLC/m6JN3MjlKN0aZ61l+XMpILBGw2u+nGKCCoWNagftdOni2VHngqJUkNI
1VSrMcGI2fofwl5/YigF3LHjp3bTUgyJAPq8jYYks8N6+tPA/XYCt4MF820xjbkXGSDtOjojSXcB
9zDi27JcMjjHCGJ2T58jSLx2ZJd0ZSwPdzCEfhrEBUV211iDhXXMZGXJc3ny6ptnpyIQGa7VIU6b
pZndeMG2mBamdW4H3XTgb0Y3Yj/+1W7lz3s3/rnqYolROg7MifSE0V8D8aoKOSL3RUD4clXp1L5b
QxSZGtY6AthggARYu/jM/LwrNJQ/rCGjtvjtG67Yky2WM9fVrU+1oJ1IYAYkthvHrOq+zWPHHqbL
pvyK64vv+F5EYxcqE2DfzJoUWlEj5EHaer/MrZfOxOu8RPWt0uLvLaG5f7Q0Z9joEnTNRdiLtbuc
FpBqX+Q1xxGRpOBFUjl8wt6qRc5NqiVJKuvS1zy3DRKbqP2aSFqR6kkvx4AmP9M03lkKpLEPqgSE
wymdd9/VM68xFd2llPiUk2qSi9Ec4zsii7wFv0Ec4OYeiyVfS1SGxteQTmdzXxEZsJlDpy7taqFU
p6tVz53Mdd8xSS/9oA66pw8XDVa6Szsqc8VNdKK4Dc6ggLNZAviJRAnHMzVs3kZBofddxK1YExrY
wwm1bLmGDF2Le7KexY0J8l35XqI3cSCC1Kfh295xqfDjPERcIV/6LUm0iFFzOZc3/zY6VgfdUFMq
ahpAqRwqxLh/Uat3umZzJR7o2TKQ96rHv7yX3RdfenADeSMGnT3MGS45y+ZXpxNBZZ83Yfu8Np8K
yBKS5ul7UOK4xvJC1B8mDRMQaHXUEK/bNByCkDzb5tLPmpSRBdMXP1Vh0IRq0voekgjnr7O8QYod
CLDXH0JALWk5TVhHiMMreIvpsEqSM91Gf82Zj6Jh7rXOvn7brBNjV0y9DoilqDY4yuGyVoMeK0Ds
FH0MxLltK1sbF7Th8wgDEzWiNnAFGSI+BtwUo2KDaCHyzanX56rRQJ9ku7iiaqB7D+KBb6Wp5xNy
qqm51hoyo/W0UKN6uL4jUuadP1+GNthTlDa5DURQMdU8qspL0/TBwX7qCAYTE3NuF9nfozkkxDP4
R6mm5pXqdiMZCcHmKTgELwVvyAEjHoz5zAVzVKQVSVrBd+E54Bfa6xt1Z2ixCN9nQ2oXDSSjX3Z0
68ZZHiPm71K8EzSbZNlRjRwx9i3G3IIb5Vc5MyCqh++dmIXIKvKVhLghgciYO6iul7e24fkRlfoB
Q2FibTkRzbFpq4ijTpD7zClWZ+GU/z7sCXVol1mVLLsqJSD3ixfrp9GmQuGVoUU4t+nblgiNwixK
BAAZ5OTnlC6IEpTMBXQDFOMyNi0A0dzfqPWtTIHQ3G+Q700FX6qA+xD8ACsX5Or/EIMLMMu3U9bG
cDUL1haJc8eDRwG3Jd7wSJAV2wHFUSSxPlEzBc3o7+fsL7VfTPeRq9hu2Up9DsB0FcuYQB2pjJ7Y
lik/iBm9kprsQT6kZvvoGnsuQRuVU5QCYg9LG4K65NL3YJ13Ptzm0Y28/rNYdieGwp6+FYuLrY1t
F6r+NFHUyDItsiINBByGCb61uKOwWYztuodby/G7EArIy6oM6KePhyb2rjJ0vAD/fxcOUCyLbQby
mUHPgfUB/mwZuFiKDPlhxRE7z0sHmBiXUqZj+vCO1ky5yI4+DT7MKeqXTOt6jmxsyQV+6/58jIuH
OfxBjEaiXhngABYn4nbPxxGoKSJyh8v2FVHEt4LG0FYTE0a959LIPea0LEIIOsTNzzMY+EpmmIRU
YfKQPdhAFZQ07f/hrJQtLU7shJ98gcojMTq6eCoeH8b3HF/NBueJ97joFwNwpyq2LnJ9d5O0u1w/
2dTK37zFylrmC82WxGgxTklk111mi7Jn/e4ufLbW+sRkkF7x50P7smph9AhEMgF1wSqBDmBAu8Ox
4+smPZydWS5tNX23iXdz6j+a93sUXYoPOTscrQmbG0olJbZrknBIH5hz1qDN4SalwOt87if6g9eu
rPYPrXKldvucB65xMmWt4ZfJtAFYuDz/d0VJxUHCO2kooTUsPFLI83iJTpzAXbORd7lI0jeU0r5/
Qj2uHdWV2eBtL2kZ8rqC7CZYBkuG/1i0CCdpJSNp6Plu7wh9LpOwDUyvqnLaPo8s1xuE4CtYLpcB
V8kQKwWed+KsKoMRXT7XW946HFTVd4t1e+55lNd0Yi8fEH/oe9BzWV2psloLTWGPiQUkUgkhtpcu
q8cVuqeXhLQHjj7yGhLfBJcRmyU8Lx55sYo5CU8WwL136/aZsJO8PxyVloiIwkDNSKqqrpusbD6o
jetztQ25c+GJK9uDil/op4imQp0Yi93s6ph2k9anaj3n/qCf3Y3uYr3u/rSNFFgq8njphakrrFqk
g5ux2nsV7ZRM4m/2GergFgLKEUc+qpVwX8nZTRZS4no7hi8ZQ5ijj9haDw8orr2PZkRoqMkLFf2K
Gz1tbBGCOKQZ8ETBw9MjU9WoqB31WJGL58RKAsyo/GL9SN6RJxiLWa6Lxr5D2XbSYQRHrZ39I7VL
MGFuya/m2ErUhikrQCGIoM0dillIju69E/WA5M23ykLBp3ThrmZ3+zjQz7VyN1XpXz2vnnthqfid
MTnRCCy6mZBQW70Qt/mqmkdb0+QiXMU7Kh5847pvY3fbNyDaEFKJc/QJ+9AXsDfjxNy98L6HaOo1
UCPtDDcwvo1CPyQIjmcFsMNqE5skJ+VQlaQnopN2XU9/kcZSsr4/4s7x4stYJlajo5ujDGZGhSeX
L3fArAC3yUbT6IXRVMfT2CuTs84WN2E/ycr9bvk5MZyC15ubup75my6TU7zG/+Rzb/2DnPFvzHfq
l8ZXJs9b/VOYHnOXfqSs/wlT8vmCq/KKdoFu5TjGVkr687zXcbP8vfJM2+aNm0A1pzB6oH64jE7Q
KUxh9MODK8TkTm1rrMPcQIaZEW6hYPmf/QW7E+VqK/3FNh/ODpgbf2I/u6fvz/pITojMpfXC2FQ/
qo6OmRkd7xKDVUHySQ+ii3n4W6qGScPEjQk3jf1FE3d3xv1cU/6wMPa4U5uDWUA/W0EVqMqeNLwv
3YaVNm3oIrEd7oSVRgPEkGiCXGpxOMfyMq1pz/4sQuEG/PFx+HsIMQOI4BjTmwSywObJyPg+9w7x
vlBtgfPv18nqYLiYfv2n0EVybgUPfGGjDsMwKmkRgD9m3AidRk5ntlLparE9heDcEyFWHds1Q9cS
PBQUvKQG1yT9yluu2K1CIT2gteG+1LaLyLTnrjO1M2RXA1zFFnPyqlB/K6ECPm2vDXFBisOoNxRJ
Roeb/vYh10Ddid2Bv0GQBMFZRal59YVHyfm8fJR3yPSDsUkCu5hL1cOCDVow5CN6Ru9XYH0DdHiS
/T92LUVuWO6yCyZ66jn4L35no8wHVLPV4mRKA6KUHVY/oH/m43ZgD8WSajlw0cdUUmoQtgPaxZb+
2ijxzwP3R+bdUogkxLmrT93BSGFQEiLKZFQmZPqpBGCO/GU8kcOi43PN8F3O8GukRrDYs1Xm6AJG
VtRp7wbybTbE52LpUDU+wusPqOvUgMF6YeH19GD896xjfMHjxVegZ34WjhZsn35hTYDjvcyOYfbh
L7jT+1S2E5PsmlDPqtRAHHcNu5O97VzSpx/6piCC1Dpbzq17mmyl/gf1eEt3+/ewk+y/16f8yW64
0daSusi/PD19j8QjRVg47SyfJemtJOlrZYXjyqD3nk92ETqnd1Xy5aOMETmVWQ8pCoVzWi2chIGJ
qerULY0amBGTRfi8mw7CRbLuKWGrcWUu/Vsdv+3yJ9saGydH1XSnQR8EtrH3921xHKRUhtx0hZd2
HjHkdXp8kzMF5ahl0d7lu8bJLQAobQV8XPINAeOS6b/50qOFj2Ouq2RpC9Ig1bvR5Nm4AcSvhCGY
eMIvSyU5dVlr35jCtTFdaeMk4YhsgUvkUmHRU0KHnkolkOWWuCcGMifHdzmn1Il4jQRTnFXIAxqq
ZhdV1wD2IcMUC5zzUzrF/D4/kzGgD/RJkRMXRWXawnAYkj+Wf5a0dB56ruONd/1+EMayBoysJ8Ue
ydXGurtZkt9WwaQZzSbt4l/SYC3URBc5KpzNkiNuo6fxEvpPImcMrUmj2EtC2hLdMcqgrVK8KQCG
wNVewMpXAyjOvDdPOiIXikpe3KXAY3yaXf1wKi4kq22JP4zVF9YEUWfDebOgV4VAhok9akZrGnRY
VaIHs1ClG0rGRZHelBpeT1RsKCeB8CzEscNNKPUd0NZrw4PUgsIncIdnftsDf5GsPZtlWR0ztag6
Hm1KBgFewFUCFovusx6DtUuoLyjS1uz8KQnsu2yCjYh4yLnlR9y+td5bEqW/5zoOscnJKp+ycnut
odSDpcxukFa843gxKVScTF5Z5Til0Slzz6wLgwOb3uVFS3GtGP7z6XSKl78n4NYdlMZpStbOQz8Y
BPWiIGTRetTacaR49bBuqo7zDkAqCW4PcL1JvhJ7DRbZNUWsE0e6H5MF6racBslSseFGpp5vHmHz
JxqYcx8wwyqeLS5gEBjs0vSM5bYPtc+bn368A1ehwGCTJ+3XJQ5/HE1LbOgS09qWiyalpWCsSLKc
089tLJ4gMXQTWiGVYdjB00U7C5c7oE4TF458MFiy7usBALKmGfDjXqTdg0ZXFlOFl3isbdCqoZdi
vKDrpZtJXaooVDJblaPxxH0z+6XAiDsdUZN+RkTaezLm/KGdeUVYK0oEQld9ttXGsBziEwRGdnB8
4rYJTmdRWeeqLP99lg1b1v1W7zS8JlFvoGhPF04E+6ctFU3u3v1ipK5tcYnet70BF7Vp7jqHyxxx
pbkiPChjcnrmzMDjQOnHpHxDD2bt5zffYy9CyrgYkSVQ3QO1FQdVcsL2goCB2UcK2yBFF3AWk49H
YmfL43iXpP+HlFY9looVKBnZwaaSBAxebBIvu2F7YlcRjvJleb1ii1R7+Z+XtCtZTItqEIAV9CO2
K/iaHldOQFNKt1cOEC53osrHLb9p5gq+enBgL84pp7hCmTLbhNLGz22SRey0yqGlGkwIKuK5LM4p
YyEySwyuAjE1wnyV4dzUR9dxLFjHFeqsd8huFUgsLAvXDRFiwHg4ofdP9j3WZBkeR6QIsioKpvxw
EJQyJYRJlekY28dCJTyD6iLcI+VI0IBKe6A4oLWmQkdeXTQlzAAA7siBUXHXFGfTj713LEydoA71
Eg7IUbO3GMXOxABlEZCVfLqdacHnYp+FGFHI45pK5bIrg39Y4cZ2S/ZYOdARjXY99BKcNSqSzt6H
1oFThlmU2RBQgg1lwM9//0np8lapxojX5Zaj/w5JT/Vyi73o/gaD6F9qGth6vWrOqSRPz8B32tpL
i+KCakAiVN9A0q8bjjZgVEg5jlgiEsuequMBOpv1DG7FnxuH065nQZmZQvVIo1DnEbFDpyzOT+V2
BpcrrEo1Ij6wASBdXJQCXsW5LJMV99RjKbolMvY3qP7JodUvhIQHWhJAf+MLqpap5SNYHUg8RjQC
MmLKiP7R12lxLaOtyRfNcqZgxcnnsOFCbR1yFt+oN/vyKFlJGOKflhCO4pA/QUlmw5f9Z0Dng75m
0iu9gpKSHX0dyQLrDZX67c9SMYsf3qkf7oLFLAts5uw8UAlUMW4Ywqp8nHNTSQ87R02fHZU3CYyp
XH/ZhsIZQrRvLu4bMuXfdqsXc0fN6QxVeb2WDFj8IMs6lF/48FD2lZRIu0nm9wjVcgkPVAyeO1LE
a2dDcqT77wxiw9Mr8ij+xuT2ABJJjbSGKg3X2y4tCueo/yMAoPmarEKmYatRja+r4wrIUctr8xkx
rCjwmcCjLk5A+vLG/lcrSTbaWkFiFPa3rtBl9EQaDVMd6W6c2+9lH8SImJSP/6tQZUoFA9c+EAQZ
cCKNNSpVTAC7TMUol+RqNRwyJzT+nQFGAtxtuUm19U+YigqcWm+UWlEA65vKz0qpK4AOFTFlHXv3
xOhh9xEeASR7MbfP2KZARMypwCiDaHh79b50XCrPzU26EHfAUh+5IeyXY+izEQUbKsgWDqitmYCi
5SKxIlUdZiIfit7iTlXflGKz8mhzA51Gee4ADnyWjQQIP9IaO+aspVg7Qo3B0vY+UEMdMfyX5ICU
uNOal0PeJw0tXVkSyZbXb+J2/SzMcEz9gqBIgtnZKAWPNtZ9KWxO3G7BHdvIn0KrFW/gbX6LLQ3t
fGWy7/KExhAE9hiTPx3Jei1FZAeC6wa33Bsun3eD1sGTeqLJnzWKi+tkYi1xZ0Zr2DRQTslUQ9Y0
+Dl1lvNKIV/wQWJjSeZ6Ua4bM0PeHrNHF0B/rDc5edEv+97a52ZwhvMJOSkxWXoOYjEcp+8MkDSl
OCK/DTp2sQFP1evcaBxSfyuGHUwyCKFmTzAi1BYRrc5rMPlBqzdVkD+L7lUxNL2x9gw9f9L48QfP
muiVXDeg3Mjgclm/QYt8yXbB9diloMKO+D9RCXLmRzrxEAb3eAauUSfPte/+csvVzLqQPUonybSZ
vulWTRCySfxjJ+qOcEbFZZ+o3oDs5ixnAGSoO0zl3UAbWsmlmOtLQYixO0sFNy3BAu8v1OuEA2YG
xXq/fF1W93bdgXtU/mJyQvr3oi7YY4ytKv/6SbV0+K1GNIQBVt63QRG/OxLkNIQFznVeO5Tfd8Zt
kW+xP43vtOTf7QkXzQtlhBVQnBZxf69QTcQVKvH2L5oCLeycm+gmg3xb0hOuVPiJm5k7JWYgduPV
/jqEuB1lQok9OMYZSVbSW+omJmZtzh7NVP6G9uWWWQgECMfzefm3zBgjb+wOWmD8TWYGAmbdNdk+
PlrL7uXyUwoXhwwkfss/etO33+45KectdP2IJDLiqtx1WlbcpV9yCOSafCx6wt9MrzUN4Pc1BB3b
0RXYup9m8Z7pVa3UzqiTFbAYY7iQxAc0ktag2aHlpAhge2Sw7y+YKDyEVXMHpJChs3T8VP0Gh51g
ffx1fhg2Q6oLVL1EQrz3gZxelbhzI99qxUS3kg59CFOjOaYWIYb3olj/XHKpMjrURDZuOMfroLkf
DjG0niZMmKvElCTINsJQPnd9ajsMAdjn7ZCMyof5ryDRWfbrfoa1aCeFAf/alVycQxHW+vg41XEJ
KbgU+xvyqmEQQ4i3rjU9bni3lt2Ksqu+cZZlLQCZ8HcvvsRBvk7jKhK7C5YfjvSsitI0J+8GULzW
ldA31jZ62YSDLy9+4ZZn9D1unaqsWgmWiw2dmxy78/vXTY6hOxWX4I1jJ4WDc0yo0sV/MLsv/v24
OJtN9oYB4dVYyix9S/GwjFfCvcSzV/KhYHCIJa+pKDQH9v/uMKfovsDKWc22cbKcdxnuElOnpPVE
KOc4o5cO9vPwaJzu/ZKqF34nHlJpQhLx2PGDL0qhX6ivUlYOTYjmEVumAKbiOjjCW6hmErynDf1m
0rXvnPYvCPvsMfr0L0DEut3lKLeGO33orKC3JjH1+qkcjBghaz/4IJ91ikv7VLBMF1GcQjHzYykQ
D8uxGuZlr8DDICDnk+l2ozwPk+NpWo8x7k6L5R61nIRli5GKNlpIhJe81WvlsPw11E/2/5Ux0+Ns
pG9ztrRAXvDzfX2ixYa3S8Hx6jye2/QWgFLD+qM06AeCibYr0+bDpXI4sYozlTbZKjaOBymuIvIf
JWWrZmoWJ16aXso1dZ00C6rEzCpEKK7qjTnPHG7nuL06dNyyX1oeO1oILQolH/gJul95sSD1fQ+A
Fj1d72vDR2R6y0YrxhkWcT7shEHoPpHcjwE3kGsAuCA+PWKMHrN/nSpEzCYxvH94CjZmjRhlN328
os2xlw37whuFaw2vDHL+o2D/H53xyQDbLcHJV58Jc9FuBObHHofQhuMqmjnYCNNzVakf6CdfWPKC
w0P65BxljaBMAe0CyNGtCHFyFVJRey2hItw3M2XLlo5jJINMkBIZRVfj1JTp1fio5AIvmFFPjHbA
JChTDI0tVPzojx1Xkn6VdLXt6LtzhDu15foSUCv6Yyr/0HvLvg9TEqeclPERWgErz0mjqOaAbwtJ
jbeG+9RQyS1QeKg9iOsIax+oHcGJ/pLZrtoPjl/+T6gVujPxoApuWUYUuFDyDBgmzz+6WPUiaHlt
oY/x446deCoc1+9QHLtcyteXCmT9/d2GRlPNKbg8KAG+dqzLTUBrSceGAPSCCcMQvTzBNdkuwTY1
BaJOPWxHEiiYIwAxWkNDthk1yDW8d5DT9y7ZPw0WCXodjYigxqp6NRguXiKnnPlZrBpXmFi7QehT
tFeY2aSeblJfDPS6oNrCleNlRh8ddMTzT4d4UQ9BNLZ3v95WeQl/GK4RG7GSi9nSVpzOfgBOWgTO
D35v1Ks5eKK/BrZBUZHuAKfSMCWdvPdAof5qOaWPKmguceiJEd5tUcB/jHxWEPCL/ZSdNRlJfyMM
b7QUIALCs+MI93UgZ6UmjXJtdr9Lqj2CpbWhPy3Wb5RB1XECgbOYbS62n4BSguxQYTYvrs6T3riq
tdSGSRZjIJo/pXsr3DYcOXhjadJOJBLWik0SL7NuFLeeSw/XKVzCWPJ9RrIPC+5ZAttdBRTM3Khb
DsXxnKUaPu0LLMd0FTRK9kns2xzHCH6IPAjXVc7GI+0DRU0Q88GYLsbmSt5Tmk3/fwHVSfnytCaK
V4UwOPpa79gMTNizqwbls94zsIkNE7mDDobaLFg57lQtDjpjziZDygsKxyhWv1Kj2OTv/D/zvCuX
ToXp8DL4yIqPq1exEM8uwQm7TOhORmFbj6y9ooETANMk7joHFn3ynCBOxG9mPwfhegclmhPvGKws
VAEQfvhvoqvUcus5vov7+hqT8MxOzDk1UX7W9zYo2HDONPkXAchpA5zScb66IeDAoOSYCkfjgL7N
Xv8q8JZuAb0IFgJpyZIfC5dnX4CnXTQLaOd/iYvOUn56tF6lGbVQMbFNSITSjna8D+foonnFpPF+
FekJvdqn+saXSme5DqRMVl+ksKNrzDc1XdBtxPVI5OhKuSlk5rDQKydfTBPoKSrJNzHhXACtup25
b4eONTIUhDT+6XV4WfkyhN5Yf99u6RtsqwHgf29n+/gzk0HP94CUUOExksYNXJhn1MtfEZlsrrCV
p//Y4Quvqo4yr/WLEaRimfKysFFc5Np2UNgJvPm1jCzx5JcTw90OLXL2brxKJXZX6d40jAtRuiPn
8Nyy7EczHy65XAf7ZdZrOD4jvKXuBNwchmaRdcuaMN2uoHz/mGzedHqz6Oa1+AF6gbPTb2cvxWk/
g6rDS3/KBENFuuZxD1W8YDybd4OtXjyT4+euit8CvyZ8wH30tZvTt2bvyrL9gAqhoWWLBaWtvn1r
6ynfO5EnaKqhUBK25wTcoC08rykbJwK/+ReQHGPaSkXDZW/grWrJBrzkzgycVmDdrZhAx6kAeBPY
zf5P8JlZLAgT2Wkgw+AaROBEm4XkgYB1bFXfo3TOJTVABna/Ic1GwvHRbXRUJV+PMWU7nBzGNjeU
nxpCOfWjFnyXvKlACiWMVBBlNv5bWe3b23iz4qZJWd4JHjHYEazd2d3ke99Z+qRGYfqnv3fWAjzL
RcGBM6jG/Uw/Oo91Z5TN0XKEjavF5WgXBj18tplP5S9tujSWYIj4HLGJRhkTqG2NrbIIGrAu9NzR
kEEZYy9juygLbew/Bi1cYGQOeEvBoYOSXUP20X3k8TujkHzkhWC/44SSY16Jer87vAZ0ocS9zK5h
nH7sOQ3iCXpjkISsr8ftHoh56cwCT/B/ytmQBDuYaGTS/lsflMZqPgBr4NOOyTXOjzK6lllU4g0S
NKySf1tGCrgZVqSE74H9R6NIsTy+ega45UUtRCRHT3qjIsmWhE4kZf+te8a8rlpzvHTHM//c5FJa
lKVKbnXZ9y/T7FysTQ8wCCp+oIcHIGhOdgirmKpckLPUIQKJ1ZjAFrFhapEw8o7VzJm21pXajHE4
v9h1beqzwNUkumbt3cXdizKJ9xMP6V2Hu7r6QyVqea6hZ2xfTW2fLpTQ+G1IP62zplbMVmj9Oikr
1j+oBaOoeD7wJiifZX2vHKrAPxF8CzDwec1t/ObcoHga/p/5wkcXE+Nf8UzZpmDwwYC0//zFfLSg
O6PS760pICONvcvE/XwwUSJu5TLWuVZMa8i5z9kYkfNDWckJPqsWrJubz1j63J/DrOrHdX0crZGj
uDXT2WWD6vmiji9XUyeLYWtNgeWP4eFz7nPdThNtfwJBSmLW1M5U3lxgO509AQ1Qu1BhuPcypI0w
xvxiVTjdYl5b3CLNXuiy5+sH5P2kb1uLO/pX/notzCpo7Y2IWgHbkNXzPnkmHGKp9DnZ9/BGv89V
pAybOtGiCjEGasjPyktKeYaTTk4tUMdejO5Ta9iVzTwlO7bALogGWYdyO1YUXPOdEJNCALAOd9h+
69o/dtzQJ/kCUjbNHsCzJrofXSjeJSxS2Np6j01MzWhL0voMTbljPZyYcm3eMyzgwl6LXQfM8Qur
GUk+6mFUcLR+1LgZUMDtJeEDF22VWJxpApSObbtg8GrMyljfxzSmS+ovxeYOsA8LPKc9acBh6R5Q
xc347i3XluXmlL2jbofjBSAQEXQ26YLNsuC6+TwH6Ytr52TgvkbsN11dY5fhhAe1YIP9TbQE5ivj
1iuwRGaedemm+z6yDpKklRJ+lzZGenBfYkzL01OhCIirfhbV0M9tRtIXZBN9HgcsiI1odpHvNBFl
/JhFDJr9jKKJkazPyRBAQu1SnNgyrhqDg7GPa2kpamjnHukDwhXE+d2nw1pIFVCW1jXZYUxq+Zpa
QmUQND0uEXUo8EJ9BSlJfFHLiBFzgWceN7yy0+tDOhi40mkWxfy9hxzQHUooWxkfAVvEp2UmIzWq
gv/14v3x2hhvLQFKxAjcLFZeKbuKc8U1/UR/EhKLEJEbVgsxDPT44Odf9+NhrfeOLuvFSkdFAqFM
0nylLzCw/ebJtWas4bKoRO0/DeI7c3nMevLGDhNV4PyI1bAid0YvKhoLC4z5chrVYCqgIpF24534
0XVddUTN2ZlTG9+YIaUt/AiZJTAvTJZK0ScDWCSNPmnohACj4Yv7vW8089gzdTrLmlLKDaiUMaE4
Lvh7qE7xHg6iFe1Jzh9/0dWr46Fsqawfm9BLv8n5q6k4wZqhOecn/BL73TmnmaB6yS362N/t8sM6
aNc2wNFDRxFGmnv+4iLhaPFWnBJzmuPwC8iEwXyP0+ud03Gw0UOBB4qRvHb9S1KEDGId0ryq9foW
IPqYpeP6jL4GKCjnlC1iqSYVAzb3U/pX87LDuc97aAfbOse7sT0aTRycSEdPu1luZMFBLyHf9fOy
AkC8QfkfzdZ9cvLMAkVBtJQ/Z0NYmSJKPjaFCzrBAdN9M0jHj68KPplHcVJoDRf03cYEPA7X497o
+gLvIb5ghkHJYsvCvYWVPW7SMZNDVVQL6hgdfG5RCcDc0HCjDceaELpWulxgG5gVEIxXMGJbcu8s
M/wi5X+SplGvyVijBcRQiDX78IsqX0ahf9wjbQrND3s4Gc6N8PQpCaAa6Nq/A9iVphH804mFGMpp
GvIHnvlG2Qi2e6d2ikE4SBCUcqr/MUzV8SdAlqLwvogpgRYae1InLw/V482naQ8yRVmKCl3pZztB
454tsWeTDhK8do4Z4DWRzlZWmA1+Xz4lFhZ9zXndtdk1akBv5tnvcwXrqidGwMFI8C2hFQP2f4Ve
D70dQvqhn4XuKc3G2r/w/6jc1yyx2LiANUcypYQEawitmx5EJ1J3nElHAuFx9NdHO3mKkWTwA9+6
TkwktQJgzqWXI4xaQOoS653i+e5Yo42FmQIuBJ/Y2psv0rqew7Noc2DS5EbgnEYcLyqGjpt5NpBd
nQVUPp4m8BzqFpPTNMN4sKfYxyXShoYYGtJrlOCmKfgpJ5rGhlO7mByq2dobyRl8fKmGNKZn1168
uFMa3vhaidPlpJ9ccTeINVwm/t8o184wG43YNBROyTs3ltQv7P3T+u48mbNWA/8hudGJi2xx+AOH
lfv9+dDkJFuqPRyCQBk6oj7LQGmb7lXtrnlHGBrCyJL7cyN1CTqxa+bPg1NpJBrEOBe5+rvf6nEE
A+E+cfuVfb9E7NKRlD6KrbCqrAE67hSJwnnEOxB//zjs2xB4SqMfyw1wwFHJ8mZlI9tRBNDN0tZ7
DwDcbf3cuEzwQ092X55JXhwEK/Sa44Co5Zo4iL3SVMtA5DTXpN/oy3L9a6N2OXhF+jhN+1jA/rE6
1ClZ4GIjjDAtFCnan+QzxlywkTg8hUsuf8LAJSJemp8igxatcwW/0zHsiDfhEDh6TC4ZsrcSx+Sj
hwJ3CAimuV1MzPlKuJ5e536H/jeghlLsCIH3iOnMZeQ3jTYbgOv3VOG0pJh56d/NyBExLYaHpKXj
m0STcw5mz+HiBcw8khxd7rSvNeWlU/2t2FJMXpNkHkT/UiPvOEmZkBJI6Z8dTXKcVflWz+JIKUQB
+/BnbMKMw0If84iKDaJagwbkmL54Ow+RAVQDgFUm/4VyM0nQauqSF7XXMiIt0weRAwNdxElQTzMM
hKEuwfwrV1HuXpdr3iXGf6UQf4CBVrTO1jd41LQJeDf0xZ2GnmONNF+bw6dlSMuofrApJ5Slb1EM
/8TZ9wg8lOp/7Tm8CCvNdLf8IVEMpDkEuT18sBXcagI813HV5djxyxzz9QOldQLOJEg3uGeLePwQ
bnHrlh6Z5bUMgmKW+vx5PsVQCu9XvoSNGYwUUTpsevMkZZoiOvnQQWxTpYnqcfw2ZJIoN/0M28m3
gxN+Hdq6FBqh1YDfpiuR4NMgkh6DkMuWURa9rDANej2T/QmiJtOabD4N7Ds2lLjOPtdtQ3Z/NKg7
Z3hfAXhImJS3gCAdxjsNfHRGSVAjwJri6psB3tkBQ4oXkEI1fmbb/hZf1eaI3LY8qAo7b3Mb+Lur
cgVvI1cEWW6pYQMcMvkvCbhIPvCDlsETQJ8LXzOWlWyrzAhR9kImFE4581sC2DzmIto+vqZnj/4O
LQq+/6vXBKojwBmsTc4sqbrbQO9e7zRH2OCHZ1KzL+9ZyFTCoLRqCsAUxgmo25ITlubUkxFgfZkM
xHVxslbrPimUihKDn9nTzgn6EdAPqpnNxuGKiNZnp0luJhDRmRfEjo8+wp6EvrTXvLSUj7yHXhiq
HmUC155Gg4ZWn7abtSBKbq6UYO3VbfGqjP/74+6ADehKjFB5rzdyFVZuff8E526KtwE2z8eHyyBW
QeskwrU7ks/YVjnDRmat0k7rei2j8ncPt6NlmeUtLybhemTpHklsdxlSVgKvQAdgYK6U7YaB/jxs
Xgei25Ddaxp2avlgR2oHGzlEcrKV1nAZqp3X/6p8GHkvqQpg/qAtxdH5+gcWyo+KrYK6YbXmdPyu
BiRFVwx7/1nGYjU0w1QDhlhJGLIr1eccdX4+yjjKq1JDSvyswO62LKhZhD05IKa5xzQNkHA3F+mY
XDGsxAeA1u3jqpAuxZF8JfkZUUQy35OYLPUNehhpc3aY5XNi7f7Wp8wrZdQwp55iD4BdS3UKmbj3
ouD3frZPfrycit6Ob5A91IkZRkswuUYo9CzR81q1b6hOPLHvBl/qjYbRlJyMc2Wup73JY9CMfN96
BwmcmOxTL3QoBQLUPfa65BNj/6tst6vSAJy3ae+UudYAqWepYkQQ16S45pElmdlgdpkQZmMOqIcg
aL8Zwmpzl+ynWn99bO7Ie/zAzYT3ooOxSyXwFJyN3e9wBTPt87RuZNI/cU8Z+KlAiLjOEfcCX1Ac
TIF5lIvS4NY4M6na4JVVSh+z0S2NgfYPrSQoE2ad6FNkSkN8+9wgdGvOIHwiRPTH1GwRP3hFOs5d
75/Qb7qLx9ddjT7yvKEm7VQWsAC5fFjgAxhUy9EEwsxQAi/mWFtcr5qTK//80TEX/SHd40ijwqyx
vxGsR7L68AJixf6gLEVBh4jTmR+/g6ap6X7aAF1yZ+h8jWIuw5voxERncqGhjNaukshdZaP7L6B+
aR76dXV9kEEd6fueNMSTjqCFyCxcoFJBFiY5IddfDtQWUTQPLxlm7IG9cgnunyZUTcl6Iw2Il8oJ
eL9iyB2erI1XDqOxmTlV4y1DXbBwiKkSrB2W76okllXh6EFh6mJXooE4r+IHmmlF02/XqEEI2g6a
/H3F4T42jvNLJpAkYeD3+7N7CZTLAk0ZgyVrbk54FPPkaqSsSQMubQCWeGRLlMbOAjdDenTkLiaV
UF8g94WKJyzQgH2oRJdgnfSo8qmbSgm5Cige06OYgrMC3AwWiJySM2jjiuqbyaHBZmZJ6kPNste8
3stTLe1IwePCuEYCZvQD6h6plzVWj/IxWEVBGjBY98ujdxVYvCe3jhUpJYpVwxtb924m+Y3F29la
0EmFgAjgrcHtK/GxEvEwCU2yNSyCemCQZwIeD5HgSh0vH4JXI/SHQHElZUsTF8ZdHv6SMFcdDFMP
kuqqFRbsWq0ReuTaEhDY3mdkJs826IFoy39eTbd846wEt78R6GByIePIPaHfB03ElcfncuFOaJl0
ixNOjYL6+a5Zu1bg52w2tkMtu3xODqhRRLO40vhDNCCb+sFiZSglV7+6neELZuvvPyee82270AYa
cUj3PkE44AefKAQx63mVn/uQpO3ocy/ckxsOA7JlLKqLYQI6yf9PbA5fz7Q+pAdH9aS8kBOjT/LE
7VivtMK/2EkYwttelLv4gAwU7qN8/mNRnXBYrzv40dngLsoVuuQ6DRkswJbTbOi72BmpR3Jsfe9W
uKpdV6aKNgKCEOvArRWGDK/5+HrvqJurA4njtCCeoKzysgRglVMgVBP79g8xnHI3KIVjthBzVKwF
yyIj8wIoaAvAs3Kg1g2ykZtYaVNmXlWD2zulNRr68al+GU9XRz+LWr/+yk9Z8ETezMzEA6tEnnmC
MqLwF+RglY8sSW4/Yp40wlsMPuNjQCIUK9Nn/koLLRPubPKxzwymJ9jSLe+gZedSU6kr36VNe4gn
jHWkbmqumJwUSZU8rIKGPKEMIgbn1xoYzvcZ1I31PRnDeTvcWjmpDWjcKkcwu4sTQAeegSsl3YUl
pzUPqArtzi7IKrsH18yUqr3nph8VJJjsiMesXPwonMGj3N5hZYPFccoCg66ZdOS3QEzhCkiQgzIQ
Wdxl9ATuWcGxhs3BT7gyyl8FtB2dWAeEqypXK2h4JXfmnPCR8gJurt9caXYPLNeIgJd48cJJE3P2
pJutmHz7ent9FeWh137fAmfv8Pc0MYeI11D8lx9S3CvTT3/Y40DsNBiyVCoLqvsuBWuXHt2taWsq
wi1ERuBlu0FXQbjlxc1JZCyxl6b33Nf7uB1CF5o7LSbNYmGEALb5pWSKzrJowSATL2C+561L34id
sMOKCW/WQiGGFkFFoP83Q1yvV4skix9DyXpawEVpOB/MogrN1NbVuPgFqYE/6boaOpJuYbG8B5jH
L0mY57rqaNYRvAxDYZAsXigvXqZ0fD6TYRRF/utIeZ8twBP624G4pvxq32G8Z6FUHgDF/tW30o7Z
1rN5ODJOrz+k+CRRhBOWZO3uU0AT9l9OgijM9/CVLwRW9YMkttQAL6nzkflYpjftP23A3LTdQrI2
GhpDJ7mQ95JmROkv5nMS/m3qSlVQE5IwSdvYMzRiM0sXWdtPgEArVvIewilugTgm1vZ1Um1ovypG
DrQOsX0DxTjnM7vXT/LSAqHNjSkQBarkTjDj5OKbJ7p28Rt1v8n6H0ZnzIYSTYI4A8q88fnj5pqY
INFUeAKW3U2DS6xvIbHAIu/JBljDtBGPAhKuHCWKdd4ypdrtRlgpE9P5T1Se2Ry/AfAKBZ/OJ5wN
FIACkbTChTCjNHY9R5KQs9iKMgT3vI/A42airHuJQgB4HLSYXVA5l9H+2VBb1pIt/V8kDGpgpnS1
xltMwIDWbHaVvfxvUWHxT6VHPGFIszoFqP2w6GtXzQ7BIDtgdQgawHEaCmNf5Siis/vQ/PcYzOdU
VU+ITKXBLYUBP/vMIVZiJyS21tTK0cx6a0COK2Rj5u0ptIUg/3TQh3ieqW8lTD9j4w0mMeQpnsJ0
+i4cakwuoGXtmvps2F7Pu9bAmRUgk8RROLnt+dR2K0dqxBtwjZW5akSmnIDTf9l5lq2YzYXYXvCq
nUgtEMaPxsMdLPr8WhQWqWR7jbJfasPuHDMMmvOhCcD+5iwg6hlTzATNorKLldskgLqdBq+ZQO6G
lCnFUsf8fnzAeNffcxHgTZWy1glFyp3SDFFNVrMWnz6AQE6uEMcmWyCkGEDeeBXaNsRq8A4via8s
ylgRxAXUaffbUx9E1l0GkNDfddDoDOnyFyydVqPZp4/tMXwabYD7LJuETZWquPJc+gLEYqy+0pS8
kWY3DGijDXUo5Kz5I7AYuAPX7+boshGhC/8ax2mji0eVvP+qtEYTBTPv0u9znVcpTEEojC9olIxX
JA77Csx3lq7qbVcYkT1gBCfYPCnQM2mVXxdXSWP9KWvdj9q/f/uYkwqGbOLLbC6r4iftgumpNCXp
Wo26zK5QyN7zk58BR2dRFPO7kOHTRN+HiDSqwXZc4SbvJ0zktgOU/7KsvLA3OZbodM4obam5umfF
5E2riDnxju8tgMX+xvk25H/mTui89uJpt7iDtvibn/SW5jnJpY1ykXHm10DQI6YWjgHcnoiI2J1y
iUoJckvsSkkAM2AbjhxibPnBYSbjjIIvIgx4fHQCR1mCfRVJI/fciMCwwqbd0Oc6H6aAM22lzNEK
zgS7d/vI5nDTUOuKzJ87pU7w2KcOJ5is9rjp3610PsKXI6CYEsSMfflPTjZC2/sMHJp/DT4knC9l
O+MAWBakG5GcFwkfAtKvFs9ERjMnhEntkc+uhnZHy2ReNYYSN0pvPCWwEjsJmKgYQVNHd6sIO2+k
XwK6FQ8qCRDzK6/L41FDgF3FGcPZXjb4VEwFtHJQddYF52YStA8YrmhLB6m+5Dl4nFONVrgxoahk
5jtTnIlwvUUtXRAQL3mCl/XILG34HpyoedzhLQCX7R3vczJUItLdNDNNNju2ZH5eXPi0JMqbdC5b
Pon9pT88hvQqqJSC9FsrjUmOOnDNSeESI09p9CJ0/T/I1uTk5DK9GF3TcU6j6nIcbUExslmaCJbc
HDhH8ior+b1JkHzQvyJywv3w5p0JTdtRKgdFJAYpGUHIA1PNr/rNg+eWgih9J8JCADKuQ1b9PSj5
jIkCZDC7kJCcE2KNQcRvOXHxAscjJTvsb90xHH7rywpjX8wpPExLIaQtsY5DJodYa+ZVaapYs6Sw
xVn/bvvFhKbch03QD4qrJ2Ub1Kssm6BEUHkj695WQ37C60LGiQen8bTqsXiBfMbi21I+zTkeq01t
YquhcEPH86BkvpFztSo6bpgHNxCwMIlLNoyzNYgFtv6usnde/jrcL8xCK3dTg5/2UuWV796o04te
XFXJe7U1NlC1hWRUTNystt7DWItXIZv4EWzZLwC9XDGB1pBSLUoCDU2V4z/k8FXXjA95DdtZJzNE
5QRww0fFEubP/yr5ocYP/JfQX7BfxMHc8URWxVYcEPtpcYtiGYMD0ovtlP/U244x9tgNr9AGnbEK
yawip+ulOy6Jw9xLvK4N+6RLpp5RuzCHgEWa93dGVpVo4bJ+YagaD3kUjkeEmxI4d9n4Y9kVwe7K
lYBrWua7nkM4BMWZKQB0qCKhmuaAfA6+T/LHnNio03uDZ0+8POSoS6Zl67sn2S1Vm9vKlv1pVVX2
L+K1q/IV92YaybhucXZf06HrMpaofb6vkvqwhp8HRJ1M6ZDCscR0qGcRe2VtfYRy31zfQAze93rS
LgwOAkg5pVtKR/pDMD5Ue2fbIlLDNTm3wDv3Xb/4+8dmXeet2xn/WCkKl43l498PUybsLFwPYvxn
bwC/iPx/eWTCT3fjXGUPYQQqIv8cX2b3mV4fQe1ikVvsCUoiVtZ6JLh7pjfrd6/9mHpQT5vd089M
9X1jCjI/3PFGxhKz0Ng9wCBJDibm5H6knMczckXYCzQdh0npUdElS5BPkO23B6rmGHQXNJ3pjTpo
vIOTciP4e32JleccJKpnLZwjfgC6mGIj95W67E52+rza77dAFmdNVw+ECe396RXmKQtLdXNUnpWr
6m3B+7njmaq2bb+C6h4sgWgigiy145fEv/UibX+tjBIDeqwOhiwAj9RsDLJ4LyNYX6/V8E1d2B89
8kSqiXDCRAhC26un2XFqqBNRXXC7lz7cxONp2+5Ajt+1lPdkbCosICVjE4Q6RmHU/PtXZpMP3kqr
IDd9iIRyAcQyqv+QMqiqvfTN4N1hBvJdUd5/yJOHMlSyhNa7/SlpWJToh6GrPWCVnED6MBsB1XYS
6TjdVabZXWG6Vne70ZVDj2dsgqFaDojrdYCJnDLFa5MLcMfsjkglbNxpHchbi/BBNXGYhmlDdPKW
DOSRbUaiAIHqk7GxdMDN1Shmatx6tvB8YhLUmaFDNEZZ/KDmpKcR1TdKlAl8HE7aivFv4vL8tRkt
jWqEicDJCGT9Fp/TPd9iX4agNiLLkNHGBPlIFMC/u5Q6KFZPIz4I6D6Y2xnQ9E/XM/YES8xM2qFv
NU9raYw4MWC3u20z2NzuCNQe3QbH3rnfBeVCHsryVmqzdS8y6dvxCoknjDM0msBAcEfLfJpO2C1D
hC++BfYmq/y75q/a3YnHSB/0DKtk1IjeIHv7gZqW7a9iPtemBhjvrTZBcAN9+ypDTmCl18LO6oWF
l413+Ih8Ef9AdL0ILYuQl7yFqbe8TUIilUTgc6xkjLl01rNiXSL6i6dT1yftWmiiURyqtuehYjO+
xxkjwfLGoVhbZOGjrCZ9/GXxhY7J24q1Rgq+e9EMwfhckqV339YRgeM+fCOODr0vur58hY4lOj3I
vlHYF4t2VRIqgcndjehtQURz0GPGYRWRJ8wXmw3z5XdyVAFtIF9Ay2bZEh9mC+30CIo9xMr2t+WE
0lv8G3sKBUSyVBb6HOOy0n9Yz9oPQDNveEQICFDxV9m/8VB8pCqHbebb1bwikRkuCKgXBfITPOnF
/8Hk/NRHixFlgTeR5odvhSCkxtuuav76V15ntmIPqo++38k9Uyfn6N6y+bEac4YqU2HeV9tkJ2Cq
BQtwbS38HF0HEIqOyrQVtcEyqDd//walfLwt11Pz4jGRyDxKuzI5/P4iDoiDRbi7ijWtNusboDAf
V0C9e6AoMlDiv4yeLstmeScmEiFpx+uQlbzxYetco9In2jQg4f/WQ/vNe7QxJnOeSXVAJZlCwl8l
5XOdo7uBpPc9sa0UXpw5G6/Frs75tp/+OhNm/8wlS65jH09cOUlwFoe4csJ/pXS/Oa6s+z0zkJTV
PRlndOFPFczp674GBwPJkfq2L7tyKI6lb02JRt44HrWBORiDF6nICOE9zIjapUTshdxQdviTZdHx
hT4JgPN5JtPqB2rVdlZakTpiz9zXQ+e1+numrk5A3KstXU9de7hRFw+tGNwDdDatX1tWC9gjVs/7
KuSOvSM1ZlJMLJTjcJQEdIP2Ksy/o0PPJ9BL5Jj4/5fGBroVuzEsjRqvFDkBcjfMszI9lB90xEP6
6S5y/UoOoYkzzVHySOICT6knT0xrPYn52FCa7qs9jUqqK1PgU3ZMqcMOpUl9n/kDtff0PZIeB9IA
w0vjv82QJMLJIDaw9wLfMaZ8Fg5fQQBHg8PMygcLZh1DTl89zqp+MU9iVXe/oyw6iYfjedN09yDo
TTGYveZXB+WwloS+cs9Ut2Bcns3zKS40LWkhCz7HmF3qa2UOynN7u5MNryn+P4slLyWWs6Lihb4y
TENJRe+rnH96xfxihGUElStmKUVeNw609ujfNSrl56LSTp8XjepcsE9SV6KZMgmK68nhKGfJpttd
Sn6S9Gc3YbqzSYn3MuVe3lT0YEVNEaJCydhb3Gf8HSEamTwGtJN227/2TAzDK1fEWG3AK3XmB3Qz
9eMpQkfh1na/yDc68ugpN9hz6G3qeeggYBBQiZwH7iD4QFCQ/PAhSLGHuayIvz3BP+tOSngCWv2w
+VHBhgJEayVDj8NWDYLqY10fNaZNlT5TIs5jy7I7Mag+8AC3pib+FMdTjzkF+iC30ncH+4vAEqrL
lu4b4belzUqZRMQYPQE+NR+Q+heg0ODXlPbUpEFa+dtAyVKhwy5cL4C7Az5asD92nn0dE2OLSQYM
hKkGB8waKuvutXpqBE15cfNaelJXQCHIO7yKk4lXlakUYbBpmJXjl9DrwCNsjBJ8q3+lJecQ1VYv
iHzictuRvv3mTgLW2S6l8rxNV2ea1FqEp7ddgA8QLNLyYrWQawW/rFgwetlMSr2FfR+r8GacDI1x
c5Vf/UZkh3YoAxoixYT3A0KT/hcjNUmHSZXcfcERC30NCrxW3ybOFa9eYjCxQy2FabzdHjMWpTUr
QTXmCxPjAxu4CF7beEuwd4a0SnmlBl0SaJmW0pujr3gguaMMcRg5dYE7QVslkIb/eZPWcHZdu0uV
xsPWBFTht8BLIl1MUxciuCdgqcMLIom5BoQ7KXR/06WOGJE6wZd3BOYg+7jioT1KGrIyv3sRWAYg
LsuLmVtzlHT+JNfzEW26Owab1ThEAdjYMrB0kdE1UwR3gsOQzKJLNby65jVcG+8hSwfy0jLmCLBJ
IjK1UpXMXGbKR2748BD33jbRK4hSyDsoo2fKaoxf8yCFN131uA8UOfFWUD0MSx33NGMXKpEqRw5F
C6zg1SgYGjk0trlN5QmT0kIDeTf1kzUbqDtPPzcYGzeZTtUuH8naNVF6Hxfjm/TgEqhPBfj9s4R3
JmbcKM5uVrq9MiqTfe8dL1pvNK8Gt3WzVPMnMVww1Hg4/lhkmiB2GhAXoZPqz+VZPxWAUBGVhWcZ
BEy7oRVx8yPBQDvp8wq509MVWvUIgyR6EP168RzaXHLqE9C/l1NVJh29x6RGWWPhqVBlrUGr+zI2
wLph+A20LSr4g6AcBQ43FkSB5l8FyDZ/JWY4aFixKII4FvBRW2EhEfYDOB6hZ2I6yTIuCvUnqUVL
ZQOaPD29p2jHI6IiTmj2h06kp909fORW6zLaJ+u7x6HnY02nBQgYAjeLtRosgMgQnEJrDPxL6EZG
PaxDTAMOFykDZ2YSJqgsEUyhLyo3Uu6t/SjsJYoZriFew3oNKwJLBJySdULfs2yEPrli9zYxk2wl
qW1/rjF7iOF/4OREZj7d3DTtvUenogYZH9gGMcDFHzIw2GSkRf+Jwe14GCGLWWnUo/9fOjD0nS4+
bYQRgKHqc1RTQE0O10/TkF2XmxCDcURON7KDzzy3iRVNfSAj1qRRtkn3TOJ+dvEthqqHZCoHNNeu
PxgOXzWDKhX++fepSq5IbIPhR6xGImTRRYfCALTxMVVv2xxD7SYV6orFc8s1ns6mqLkjqfA/dABa
LR0ewZCqeuzya+hQT+LHTrZnirVLN47MM47CRIv1MljxUOolCED//VyODyFtpMRFPUcYHyImT9IL
KMHw3a8zhq9qFTM2aFnoMIzhExCHZ6Nx6vm2Ej3PZ0No6KCvJC7gvuZWyBXhneLU2ocjVRqmFYDS
8qQ92P3bi91qLII1GYK72Fl9vFI22XDDo+/mr7ldggbk4Ou06s8iLe6r80HTO2w3gs9h2DotCHLB
52IysVRJnZJ0FyMe6TKcKz61FZCLCRMJ2kERUIhDFhJfVC0rnzfXQc9yZ+hVyC8I21WvyL5Z7M8M
/g+2t0sQwy4i/USUsiZGL4OcK5eiWTNsBAZDRw7KFbRfPhvbU/2ZgZodNUDmceWC13vXzNgG3xUN
oWMr4jEet+xbsthNoqtn9naWkoFl2yyOZ+mSWVCtBbGNhIYmbtCalWfsh6wEPR0mgCU/yYwmLu8y
WanGIXZuuve+SeVW7JiwWr8kO9QLr5UtDGqEWNqwUN5pAVuyiaGkmJNceil/oJVQTmrX/2DwpcR1
9TVic1F+DzzCLjzxFqq1yN5k4zN1FNUpStiOJFpvWpMVgXVd+s70QYncG7uqVSyzbDgakUs5csBt
ccfAZoVVZmNQhhois/S9vgEdNSLbEKKcBZKieMxx5zB5Nj3i4v6qPUz4bFjoBa8xwbR3jJH9YqvX
Z+0/e9K13kYg6xfModB/vH6zXia7OYvjexnN4xFFVCMAajkXCWOy7s6w6HZ3RzPtSjhuTD+CuvH6
mTUjWQZarQNaAInosI7/EozUOOqqUjuh8eNwrNVzMOL6I+f+aJckwLs6penSgmrM67v5PnkesnWc
eZCtS9BnT5ZGXVmzo2boBIyqZfcyCkzNJhX/WpGolM+jyC0F5r78I2lOVVh6Fp8mvjvItKIcN3G8
0adJvw/grqmthB0+j7acmLDBehJUoxjRbp00vSZNU5Wr4kxCtg/WEdy25pnyZYoAWgAeVmulsxKN
aTnsi3GG9taBK0lQK2Pxth7slv5q7321ndjj1JfzyN3T5hMeMfsYhVAQ+NtZQcHOvA5JkJ98jV7S
eJgO6YUMM7c/KuH03qzc79g9lxMIFpym+0MJyQawWMeHMl8Oqt+8Py1ivLGwiiTtPkbGDQYirX6R
RL2VdrRDyv+SrUMumxucDoSHBGu7/Hyb6Al9/Ns8suSajP8er2KwjOP9dTt8nrS2WaPRKkKHFw8l
l1w1jys4jPj7LUFZ3Q1Tom49IfypJQtSopszkslNBN1Vdaq2l4SuD5DlxkkszWDX+YA6vVIXUn6u
rTZbf+DxY0DdhQF/FyKrQ+g6CqLzMZjQrXiiHX4HPHR4DhDVxO26UEs4WnlXHKyVtDIjjzrimP4+
wu0Uwcp09BE4+jSi8RbR32g7giE93bx61iZMtRN6y8dFuFTnyZnYW0qYt12ajmFyqd6rkm7A7QXV
9SgAlJS8/8r0DDzszRcbxkiczRcy4+Mh+8brQzmbrNf2gn9Uhc99MBWq1DKy03CI5JB1F5J7LubE
ddbEB61ck2m6Wh3oiQ3LOp6D/NM9t/ZICwUF098jQkfz4I+O5lEoBSrGhxS5XjNHPxVYoZEeFBeh
KfNCrBzWuWrU4iCjK/Bhy5cqfBkPp3mCSRa7IDz9WFgj3j2Fx8w0/mOXnuSi08xHWNJaSi5Etuqe
qg/PaEw0wZ9VnwqECW12zQoRfGLEKXwZsbWge2OsDQvnIWj7c6DSd4sG70x60kYEA0bu1t0E+k71
0sA/1eeQnDIO8nmeCZbdmKysIhIzTJTFrVo8kAr42ipmfUhe5LG7T0IfEH/EEBsX92tt1D6JT7gd
4IzXVHGiGy4I5TWLOpcA2w9luCjnV0W1Wzgugw7nK0d+fFReVMfOAiLdgl4m//KBcdb/l7w0PVIe
0nZ/fTOe4pTXzwcrPT0604D4c6RJdhtfERWBQ5HlpHUeK8hvHkl1PNZEIdfUBezubYUQQwBMBui6
KfTJp+x3U0X+nW82Gfv3OzBgkfyHzhz6uk6WdPAcWHqB6E6ho8DhxQtueiXnGanePUsLV9t1JwWX
87cdHuQDl+70Lfa/K5GOznKtYMZMp3M+oGhoYZ9tXcxM98r5OufW2JkiLsTMF5fbb+59iPb9I5qr
2W0aNHduvEC3F43BZjPIy5fPbKzhi4jnZnmcWpkCtzI6Ikza8V9CZi75+s22+imzhlroE8txiw45
UOum3b+D8XdhLb7K1FogHuvKoniGfxaSrzPcwe8MpI7Rag5GKOJMlIsZ6VyTOSaWUnGUn8CKl1Ii
U2bjoZs9ZhgvfClKZCDclSuBhoHdwRnQAaVHYP9F+6IqKcx2lw10zdWAwIx05sMxAUaY46lSIzIZ
RK7E9M1U798HlSq3UL7HPWwgK0lFO/gSoV3KjElRtJ/YhZcEUtWQXIH+BswIJWijuixIP0UkaEtJ
I1m3fJ6oHSmiC0TSUH4XIfMZCVhdpmUT6LUv+LtiSRlgNpFuGVr6rQc+175KQY4dyNYsE4SPJRhv
hFrGCBWgQJ22WbBI6ssqAcy40rVij4R0shSNc6Auv4yyT3cn78FZWNj4ANGQkC+VyABa8zxJR7lZ
AIF4ulkTmDvwgHJ7esTuAYdoZ9evydi7mpLAwfhN1+xddaNH1y3irVGIi1cZE1Ddzy83YcvX4aCk
W8R7arbxi4893AvQjqtcpd71Zul2Ok/ZQTGkHC3eP2hzTNY3cCUiGKFzEYIiY/YdrjSSBb0pvheF
n/uGvMuNFWyRKhUDS78PLrrISwJhlx27X0N+cXmm19hYzOeBwlNH41jG/c8l+N5jC13aJ9+ibDa2
skgIAjUXq9Eb5bH8kZi5YGlQFlsp+ScJPaADZ+8E9f8k0iG1NIikJTHvKyZLfM3n8Y8V4pT9ML+0
ptC75Khn9MFtQtsf9owTnoC0qboi5PxLcryXRVJs/FlubIFUrOONI58hwivL2umuld1n6EjnCAyL
rukukb4Euh/keZrLrcrv0xFLfmofwWaP4Omf/xL+czguVpCrvvCFdtJNwQ7T8hVQOYHNbgVnnTeb
VFiBAj7TnAQcxj2mTs0RBmaVlUr/pmr6ZbzEBii5nSYaTX+nhWkTlWcsjKK/NYxWgvwSiwek4MZQ
IZFx+JKIoItvBDhFaLzbLSrB8TU8AyO997amQoWf/aPuv2lMSLFrlVQPuEs+4ZZDgRdFkHBlkfxf
rSbFhATyqQHH0RIJxKrAbZU5EFgztlJnMwcDN28NnuvE2z57MDSK3AIHSQB5b6WQ9GjhIhy8ZbRR
vm1kXFk4ZyXhxsXodzSe3yLl7icozKB6xxrqSwT+NZvjpE0x4ofVQXlve6pjH12NDhXnNW5W1yky
fV6q1pGIUF3Jbcd5qkOXoxDzDFTQO78xnCUuZjbO85MipmEBym7RDIGLxBhcqcQgQ7UAasDG4i1g
3p/xOH9rzwdDjiLeZGf8543rONr6NbUY9iu/KnPmMhYMZI88pnsVwxjIL1Kx0/4RyQQp91bgiSaj
WPuwf1j8afL+dTK51qAW6DvWo1anfd+xlsusZMbZdDwXJitC0En60CBQhe/BV6/F0ssGV9VSMXuQ
uFvsnjUYSxzks0NKfqzZXJAykSBCUrUOK9fYhPcW1xlNJhjCAzdGbDL0JfsJM54EfTRGIWTPGT4s
fbUtWnKZtWvr+yZBbGeKuooNVoUigRLxiIO3ZCOE4wq8ItLo85balzXLKUhMzRgIozXxKippzchZ
9GgMtO+S+uqI6nbHDxUava4AQ4s3cenNEtL2XzVhwKHo+qN6sH96GH5QmiW628mKi4g0pPBa0sD3
ZXmCOtE7696F9b6CNWiSpBcmQo1SzCZoJwsohhtKuOemOLk1NVUvAy6mdLfbBJlyr8Ve0ecU7aJV
Ufjr+q0CaB8gwxP4k6Z6WsHj+qf4kYbQBrAsq6VDeL7uFJd5QPdQUu3B59/m5CPmvW73qc7PgF1A
2ZWlTWPZEpsRB+joc3qeb0NOjshF7ZSYDebWIRB+em4Dw/FZHb41AJcSqICc0a+WWSL1u7i3/xm3
C01lDrNmQYwy7VlsjEWHZBn0xMfnsRL36M+sqaLvloxoUDM+nUpH9tZiSt1CJQpnnuuFuORaQoJQ
VN6DRqudhM7YD0Jagpb7PBLSn8fmV2RrTFlWDMJAH8S+qlN27nlUUqDm1L1fJiJ5japoN7MDNYad
D3+S9Qp3kcu+kCEW8N+7iBWKCQdJceiQsVK44o5Yab8yLDPkCowXRZaZR2sYLl7aKpc1Lss1bGeg
GckoG+JqwRJTNzfzFH+I3kRwFuXmdKq7fKWSajFdb6UhYfwQ1bBaDxQkfZHge8R49p2tmwbYydGn
41alLsR971eSIuXh0X9ED5dNEJOydTL8hSdznsW+WYbnL7q42gEVa4ASGl5rvNidtlnBpu/nJoTO
pae0TC/yxqgmOWCH/h1mPAkJkyB1idd2DrZEgG7IT38NQNn/6U7uXKIS15Y4JTnQ2Gc5+AkGAadq
z70P+HG1MetXqoHjoxGUb/VVjSMhCnRA3KUkP9V3V99MCX7uZaxO4kuPL/2/NmhU16vM+AZKk+CW
P3/LcBRrwn+yASb5tiV8/sKpLEQ9NKaWW/7xU7LEMi5koaMiHwP8VGPQ1Gen2cf4Xkl32KpNpdge
PAM+pc3LXES7nHOYume1H1aEHjbr1FHJixFxmUYqSymkUO2D1t+Otva51PCzkwXuVAL1Mh/iTG+/
HQAYW6ybPAWGvSQ4zklTTPYSp3qmdimBQ+wY+ctZpTPakFMMU4rAdXqNU/KaW3/8gutWNegvGhut
kaeZHLNBeGH6y39Pl0irFWXtvgOsAlplobhT+NrNEBCjUU4fQ8DFEgwSVelynL4tX1hkTO9Lk8EA
SpydYVSTi/DDhBL49cAv5SJqQl91ihCJ7P9mw4D0xc+pcgB9+j4SZhEiI0OK+eSWkCJ9apeV+trX
WcegSkz1GTTmxQFBTYhNQbBzFyxxWrkG9FZmb4l030E3zqM4gjL2Dr5SvjMhWjpXnw6jch/nwj+2
wfKNve1jM2LSlomEzd4Q/6932ToaVDbmBv2LcA7N4r0E0KHDhV3j68cvfZlwQ5UDtirotnpinegq
6fSJauSI3YId8vxgl8OJW6FvULFeRm77kYNp+ZsoShFWuYAn/BdlpyipGtI1x/5iRevE4fNg+N2o
n3qqKV5OQbUteVFEcbDjQ402Nh6WmqWXKE6QTCZWWcIkfyUoLQCgyfKdY2/XZ8up4gYVk/2sQfud
4zQoKYJT69VMBqvKr50WuUcXwBrhKU0PrV93ffWQBv1d28p2u3nv+vLv1B+ucHE19NkdYczOh7gM
EVYts/LSC3CkFMOBkj44NZIWLFIi1hO3C3OI83uRt2GjtsoyKjocEHulT7dQZFVk/rYKL/1qV1AK
2O8DRN/um+0AKJXUQhvIaLHneF7w31m3bwNRAF+PrS0eCzdDlukIToA4BaLIgqtBacFlC/0tUZXX
x1g58U/dMraijwxSs78X/9zlBuu/rx+9fTDwt1q1LENft3U1kPamrAoDk2qllJxIcq/DX/9BIX2R
9Lu5Gsb3SVm2CICSYlNloFQg1PVknR4tfsnrfs/y+0tR1czF81tLYEewvVnKUA/lbllU8/od0wOT
VEeMPLgRQ+3oIOzw9YoAtgWuddc0MiYswf0L9eSg4w7x3xwW+fcmrIGAQt9AXm4IxTRHOr5F+ezc
NjPDU8snh+mAi36KGfMeykVYQgf/zhJLk9GYTao7lW2r0/l9uA9NgYBmAIOmEqZAr1oLCivDKMb/
dkZStJEw64pvQFx35maH/ZErGc2rsmo+fpVqsAUZTziz9ZsrwqQT6HnhgsZ68kqRwAuPThmQ7nVb
OfZ/uHPKhaKW7Mm4yMeIe7rirveLVNNu+M8o8L0oOPgrPYhncbMOTOFCuNy3MytJ6R0F4Fp1KNoo
TJ9pGDP3OMGY/KK2fGCLkTuyFSeqaBIPo8jf/g7TPn6bh8fF9xecmSvqhbBduQaw8WmKExhAJ8Sk
9XagOq8AC1QgXJrA47WWW6PYhaTDUhQRd0F9nhfScH3NO+dVa5ER1YCdc10zDM4+6jI+OTct1N8Y
C79eZHCiIaK2cwkPmwQlSZo/YmRVW+Pu+TfirbGZxAlhpyM6CVaLIh6glRT86XgjIIc0aaPGvcAD
hbcHZ00HvrEn2eu/+DotVNsvplKvPuHBPR7/8/KKCGJiM1T8nPo014Z1bDJDMer7hziOTKHKGxPT
o7imC6qOt8wCm/TLPqNIkE0O/4devgwCvhxBklWD0yp9E/6muhKY6k2zvg0VBLOGKDyTx8hKVdAv
VpQb1CkpfYR59MZFG5eZh4PPcmamT/eW1/9IHJMuxqX3/iRhTT/GSZAzAMYQwDtPVKZgJN1rTX1k
y/pg2FGA9MRqdpTbdT6pnSJF5NYXR0Ww9fVHOIzwJ8bwnazJXNZCAVg6KzPY3FOpdx0NLX39LBIk
6k1704aqHQriq6DYBKy8N1RIJb3mUx5djgM2X03y38z6EWg157VnaxXSKzDPhbOOm0041wjN1Src
7QxjCs4OUPsj6URYSwMx/8/RFskXDarfjiY9/MAXeRERYEr++lSAfQrAsVrAGon48tfEgqdnB59u
AeCIiAf9qrnJxC8LW+Whsa2f+j79EBQgoQFVGVn6wEeBPXLTPkoShLela6x66C0w9VP2oDrxli+c
nqsTlElQA9Ht2SucUevA8w4voDGYTdXFvA9MKNTRBDzFHKSruqNBQhf8T88C/Y4SVwbY8EMV3Dkw
llIev/haV9f3ZK8udSk+/SdDqeJ8fOzQNGhFf52LjRTGzfcrR4Ak9IXxGfyFNvsOV5N10yq0vAnV
HvEWwkXwtzk2QU4jtBpUHzleEoWJUYmU1olcBQ8DA2COxyQd2CSc0hP+uTaPUfsDXu1JQ52YZU6y
lhuVRxIaU0WUr3Fg9OjJ4qerqQlFST4C8jKpQQaN/CyADphqthhUUlOPv7E5MR//71MO9ySh+iOG
JIvtoY2mJifnCvxxIzx2egQXTrs+UUk/cIFdHw2EjOUkjQmRiKu4ORUpiVzx1sVh58YjE4cfcmYf
/agt+I1/x/h6eHLouCOJBqyR1ilQvilQPEiqUsRv44NWBe4iImVVK8P3UHr+rTIKkfCShVdDq2/P
PDdFvN51FtKPlO7hQx07ElLuvrEvtChsqGeytezyCGmcvOt23NEyeHCJJxpDZqRp/a+cuFylyyS9
5a3lqjsQmgnHAW6+cwpOO8LLllueyqpcOcTzIFRIYQS03Y/EiNeqvfEr3W9OP4Ws85QfM19W5Rry
ptUQNMhLfQGPfGT8yexuLW4tVG7MeFhKu+mmwRK5rusZchpCIIdQFP5NH+JPmiPIP9avxqDG2RDs
TU5cHUfxiwC7MQRD9QQh5CijgeZEGQzPG4qluwdiXMG+od2d9OvtvYwk6Z4dK6o9tXym56YnnuZb
878/OwWoV4djOBciYunqNW5c5LmBMW/zn3Y/sf3HSfRC6gS2BnYWO30aNN6343D5YcMhJ3StyWcO
yhngd2G5EbeKeO9jgAZaA1p0fws6qTgwipdxcRYzPgY+HjTxBh0U/yxvvU1BKdVpFP1VP9UvIn5X
GmyPxvlxhutD/UZhIdfEIavFssLpKqceV6izwshv765aQ6SyHPEfLO8j+5Q2HKVMhQ9MQCznwlYE
ueamprfy+5dQVqQ4IpO9neC0BtcsgNI266vN6Lqj6Y5ijHK3e9vo4EwZBMhBqrQBQzelOQXpymFj
fn1krTqanYxNlwt0RzkcKDxr33P6mBAsZX26r7fxG8OG+7jNayAsfhCEZ9RwGpjZLZlaETDj/ynN
FHiM8g6yV39C8lrbXNFKDjCuqrzUmOMSbXGhmH9O2Hgj+/3jMJIUyyslKSZrLrNODr7Dzb7DXEVS
P9gOv3q8tmy+/j9eo6pt/esKUm2YfeuCDWFH/3/EQU/nOyqGGVmimveIJU+MHlqSVAt0+4DlRtJP
iI4UvvZdAepuA/vX48BXhTdQvfSgSQ1HtQUjGZ1Pxy3ATQTfVsQShGzPhfRShW+8PF4HVYf2TF4k
vcxXAaDGKuCwgEp57MTlMsjcKLGavTPOgCCi/uJZm/vnA17ZdOrxGMwrAO9w6lfIrn1HYHflm8C6
PjKVvGRhVteCqQdFzggphAa6jxuivSRUf/chjb5y3GSbYm1Lq7sH0RoqyxWxjMHqdEr7qj0wLs39
masAS1HMIcPtIvuRv8FxWYwmSw6sn1U6J3UBNMxeA54LXd9Hz85XwyU+YEQOGCCttsfI5bje0ZaV
PbcKqBEhD0XW2/GNIWYZpCx7QAZirp6zGDCD0t1qChQMRMARgz/BdWMt9LWrm2uz2/REOPRs2RFh
5Dw+RNlAYDQZJ9DRcHYnUZg+y8BqC6lFSsglvGQpuVUk2I8eihzSViVc/t51v7WUuI1OOe63GoWq
xIcsbt0enMHym+2Phbem0D3qLzAhNO/6rJRH4ce5uMz9H11iywwUOxzhDnIeuk4GE3KfW/4He7KS
0FbJYGo8/fATIYmYvxw9BCZoeaNyZfXgasPGXiiB5lTBjKQk1odf3d964sj48lNWnO6FRhdt8HdZ
RiUC3xCRtsC/8g5XNCpyLa4ZEH6iOJ1u0t78QhLvGEaifxkSMaQ4AjR+7hBOS4zssO0+HdwbA+mW
iFS1omQ9UCRK8WiSniBtorw9cGkhVMSpEHse38Z6mR05fVai5lf2o0ThCmwdicwofb8OOvsR1chI
ZKUgbqvY8SHd7cEScr5W6h7vvHHzd6EeRkJdY0JFCh4TzDRQvllBsi3LYQVm42l4Uub9E7UeodtG
w4DE+JdK9QO3IxRFwr7TmfICsALS17oiFmG5d7teEXJtjSE1gZV+aNeTgS0jX30FxqDSC4wGOx2A
CN05e5I2Lcy7Ydl0PWnJMItCF9ZOuQRtsCP8ifLZsq4NTwiYGJl8hf6/zQnMwXfc/uvvXf2Tixl/
gzdy6BYryaSeqRs0SPH+NoW780geWr2bNNWBON3V0aSGls/PPmRb94d9Qd1e+4jNt8D8nzfLjixB
Nmx2jMArAecdTEc8kzx3xcS9Q5BTMs2X9p7aOAUQG+2Vy7PVjtVIb+04uraaYMTUQXu3Zz6PYcO9
/U0uRx/rjizJw3FcRQJiZSaDyl1tZGT67LSs0oePz9SGBiQCJzReYucuX5Lh8OCgSmekVU/MFBNv
BB+b1vIAsmlu6guW65ZVhzeKgIKYK8e0frUr/aRj+poSD4RNRYJfl7t++LsrVXgU+UzHi7lD7KIS
UCYIKqSXgxmIHfFi6Mf2WQVQ2IRTJVyTyJTKHafuSEQ9fW6k668UPiD+HZnRvAdueXgJRgkBQjej
l6aLXASwdtrBU/U0OliCpjzuwB2ejQz5zULOMmt4aHMQB8GpVJHj2l2m2XyUZfAtyjlEN0oStA/B
YWXXVS7Ps+R+LUSl3kHY+YexflUxwKxkry9dwJpeRHcfMsgyVxqQMCgmzHC0LuQLvP7DLsj/N+Ja
L1UC6av7DHMTcX9EVPdbJVmHl9cctBLxY2LcU2KTv9eMn1MumW7Wv6H55+uGk7Ml4fEgNjdmetzP
vyS5zgvJhhq63SOOWeKstBlE1ndO+MXbb9ib/5DFdj4cX+6w5jSRj4r6Z2Ug1x2rmJxNdPAAniFg
c/g86g0ksa+NVQbGOzvphxLTn2kWocYHbWjzgoC9zLfiJpUxBwovdmIFsOBxb80s/J8d7ydQkrwA
J8y/yaUNL4//yhT2wRgeYXmLQsjndeSmQQg540qeyuk8IVhUtvTPzhhrw1MerGenUDV6zHTrLXKb
tKPWsXP0KMprUIKRG0K2Utw1IMCbKv+PJhqa89CNGqb9kjDCjnEo/QgLO200x8jAjUlfDdQojUx2
Up4+GW98wPVL+z71/nIC7UXLVuLywk+ahhrxx0FCfJVph/Y94kPHKgv9FcYhH8JW/kkm8Jl47csz
C7WfUpIyUua0wJG+KOvySH8yVyFa/32UMplVK4/rZL2Fe9UBTXuYXoXU0oadsPi7HNnI8i1tFOct
r6RsDGHDTy8yb/jkYC27n3RNIy9hYZ/XMUXYmhpPcaKc6XpstNORKVYNKgYLe4R8TJBFvCv+VBzI
BxenWeTXQgeFPjGTM9SVzim7lLbzncuJf0DoJfpBqlHl94ahV0vsiXd2EQy+/4vzHyl83VF4X6Xw
6pzXl8YPeN20UlJWxh0nErd8YH3ua4TKbKMba3vKmlAnOetKCAXEFEg9HmdyD9VClxRVAn69dMHX
gZjgIeJpNV9RalqGLMnGtqkuW5T02my0nhjYGnlNUQVuLGrDLKMKXMk1DvPj7niYRFPdtbUj83dB
e41Rqbx6J7Z1+u2mN+pwYw154ysPSsv/v0oe47FDk98QE6GviO3asvUghaNfwBeImBKWmu3uxVHO
Yc4aq//fbG8yTZ6wWAYoz79SKzbCfb14OaI6SDwI72sP3ltTyrynF1uusrGWpJCo3T/vfMGGGB33
29YB8cQIMxsP5qlp5t9sH7x/N7yO6MyGH8OKrFjSurmjC2QMaU2d2sLVHX3fsH+VKGtYlMQyXaeR
T1BZKgazRXXTIaryyU+58tuFecBZmobpX6yWf9r3wHheWlWjNdL+SvkqHBWeldpYp9CiLaQxLz7c
wLv5q5jhSk8bAXf/lZBVjTD4ZdJchXE+p/XKk77OLLgR1xHFwbS2VmPZEESrEg612mhxoPNb7//b
Irv5KUNlY+g6E30px2R/Lk79nZOnq2t4NM+7Q57EPveRUiwSTgz04Jr3g4lOdSJ9CC1/NYDz6AHM
4AKnBp6PLScnqkB/xSN3cxTyA4WYfvsDPzp19knJ4G3LFFC8imPO73Jttej48dUMZCLD60hpA3je
nYvsrPGiuyCl6KVczgWuaVmAgTuw8LAAdwk9iA/VCrhAdHCODyrvEBF8k4hW2q7ncw95hq897icz
WmAkljd88sW34YJSlOwB5dFX4gsBBQ4LMmpOZoBASIGXvwuZajcaYi9+vvGsxCMjaskUKmChpPxk
Q+dD05IiIJ/j76+NmijNqmUkau6e/ei+eoyitdmVTPgUU4ZEW2dBHDF+IEwV1fkpz8XS4ol9Fgbx
/ElzgUP8R7kcSZM15bLRZX452HzyORdwVd+mSQNJLOvQKOGbKQT/g3zWPvT349BaomUrxWdyWeij
QAjjOyBHDmKJJ7j96GehXXQbEMff59Td8YAu2Vu9khiDKei2xJOYeCWC43XupNtk2vU082NMGLsH
RddFt8bO7ioo/LdN59RZzc22E+FUmxyPMBrGkIwxBhKzVMWzPKfsD3HzmN75OuQd+QzYsBvrKMKW
nKJ2PSaTEmGf6ocn3PspThP7+2+2kfPLttwjY9wLM3iLCDEes0iMqLZJIbHNq6w0+0iNDDeEo/jn
FzbhnxW/0kRM1Zvdic0pZU4MoeKwjtNME/vcFAw+aXISZaKPmLozSPnPsfV+FHnuWRhPbGhl94y+
Ov2ZMJu/qthWNo0y67UcGNHyrpZUlCNlm+OnQdLU1LUQfBjUBVFWWSOnnN8rb+HLy7HGYDlZe+jM
UKUkI093EbgZmNIyYgOxnP7IDaekOFAoXZXwYViLCsfGmxVAAMYT2rvNcJdVt7O/Gta9OfuZkf1z
ZMxRm3gtSAwuAOvxjlQlALVdgcfim8F5h7ScDXEprLdZzUAgsnSv3DvUOiAxwft5/BaYyWFk0X1P
wgI5szA+gXj+mOK2XeG67AERdJ95+dure2uKbNdf5l30iM8bisq8k58hUUF4zwfh63vEKqnt4TKk
ITeTUTrGPLubSicn2uMjAtx8/GhK4zf2Z7BHHFdkjSXe4FP3tDf0HcLuCXmS750fTkNWsMoncAUt
i1SePGeXgvpRdc326rYYscVyYAFRLfXsuonp+eHqgce2P8bwF+1Gl/ih+PeJMEoq+sp8VxeCCqc3
8fDYsWA3kQdjRwPUscpd7Av4U/bsnOyBtI+XCHBtrzWy/g0j3qPtPKfvEuyR+4AN9y2gCsHVNqDy
wesQ5W5Z1v0iToGzBk/d82C3oClEyaFS27e9iSN9BWP+U4/okiM7HaCDLezR/VVYdT920OBu0YPn
IcQzY1YhtmolVdGXQ7TJ5X67VNAk7N6S5SMdsD+FiUWHnRHmvtbVN4RSSiLgky2cbLBblAymBWqS
mf6AOyjaGbEzbHhlltTd4zxtWGUwM6fCaXyIqBAX1D7tBOAkXfAp5dAP6JL+rS2SlDv+RAIdtX/0
XNxvuRGa3TORFZxOmrSEBMZTjRs48dtz7wlPJcoGRSuY87cJdBoZVY2RRCFD2KDVLuNiVd04TH5J
LEESASnuOzBZJ7ssFRoWs2rY9ohXbLAmfJtcyO4ctg+tiGngVA3vOhh60VCtgmVO7Tv0X0zsiekB
ekHmbyd8YFFOFyy4y6FoXuuNw/xqAodlpYCCJbkXAe48EBzZvOoPVNk0kyqIZI/AXYIFhTanwKLb
h0wqxG4ElEeoabWRLRfwRXDO7Kdd4LwgMAUrlWUGguiRmElR2XaEWb/FaQPnEnFidfeCyC9Vt3i8
VwTkelhes25pB3hE9lwjuWhf5PUUtRgqcV5ViYNMwxSpqTFKQ+ETB3zUMJ3IZ956GVqdy9k1GfrU
z2b1ru90JTVSfRksuA+uvkS4IFggIL9c+anBkWbMB1OwKXArun5wOSfv929puWtt0KyYwmLgq6LC
I+qrEfBwi84tAiELEaqvL5UPwNTIbkr4u80omH+h0CkCTn8TFfNOiThN/4n6t8leKtE98UGFEBjp
l1eZ5Zyx5MTMGyrqYDG8lzx90loGNVHCk8LKhfUlFTa4TVxDyOFp6fKrWZ3myGrrm7A0gzrXyLqH
g8iTcOVyx8ls9QSclWdFzsGyDxmSVn/pRmm3PQov/Q7ehGAd2YRNv5TdamcDWhPN0STaizdWkFKw
caNYn83II3SMoi+MZNJ3Mpb0Ec3c/fGfRhTZLra5bxk1HY/wXQTl/3dcYKX44cxozVEUdP7aoNWj
uE+LG2rkzEOV6+YkgbiJp45ScHVUQcfgDROWgBGLhHYSKBAi6ebiuvS0PYkw1sk6uQoDgFJ9HZy0
zTI0K9ty089cU36DCKbejPzfpEo0hwRVpNSZt5RWsjfAuAmr+aPsg9UkcOflpMeTAc3iXqieS/eT
IbhgQ5yA/H4mB2fCnTcOSeu2hH4cjXgG2D0KdBUliqV2NgDx+ighXIBNl+k6pbzDPgCWfV5Q83X4
A9eE5BEDh0o7FMfIwEwYgih68fVeIYE1ZbH4e0yS+t96zfFbYFa7AneOq5q0aDKDC4nrVxDH3S1h
7auA5ojGnQbxFb6DG6r4oNSfe/h6mGdK5mIOAYmUjpMzgmfO19YeA5AfDHiJ/h/2bRTgZoHhWN+v
dRNENSq8f68YnMnVDV8X/8V1big6QevXaVaBaYnkH+3yD+WyXi/5dsnSRAU4PtZZENLg9vAA1oni
+ZHrpnNuYOZc6bbBB0JCrJSgvwnIbUsH7YOHMgF6nYwfZnivBwCrNM7NCpyRpT58mpbSs4glDIZb
OSmcIiPSRdE9XKeqZqaRtHPnXqJt0SXBhkwx9bWU17OitqU2d0u/G3TJ6p8Je/NTh5EBxIcpxhDR
+h7WqAf8UDtLE+MYOFHma212+2hv5bhvSSXCa5Yijz/+VEI+DDkQ0peSGfMtTc4Lk3LlICTlxf3n
yyVjo4dFLvKnSTGxNGTCssldmCBIrLuP0lnqQpHnMhYsGQ9Ke4vf1pOFFzjNK6t7Vj2N3Hup0jYQ
1vuaFUVhePXkvhfMb+vbf607pTdyerd270gT6G2nVq+TvOpRjH5pEdmZME7vTjFdOi/ZMdjau8NU
caw59cthJJXdkWFRsVwCYihuAFLksZrEb2GWnOLgs8qRLMhiIIq7sSqNGwx6I06SH4okcMAQxxlC
E6+fkWtXpru2/79ly4HDzMbS0yZhd1DUWfizC9PIKjD+/t4MXW0N9rIqTd/ywEg/i1fbX7AonfqM
wjVNd2BFI8632BcqVVtUUeHBcLeW1g7Y1oDdoaH3nY+B1+/5MC0enwsdUj5SWUIJoJOHKeXvLo0J
4bmrgU/7ksWjlR7HUsjx/1I+JmRrQZps3AtjHGhNXjQ54TDlE9Wtxw6NJ3R/xW9UGSKEmnqHQaos
hvcuCcamML52WXt7SO7yqwkFWrCrVEhw/uaz6SHkznUvevBb1VaugBh+qtcpRlHDKO9NaU6cnem2
/LQRx2cu/feIh0FUyoZcf5cP3LXIWg2fPlQT4CDrtxoVqOdOAMq4tUGwoEKFP59jpnIY/idJjs24
Irx2gwNa/lsMzcvQjmWTL+wlQEAHFcp/oBe75uxPV2RS55rM8pVEsRCXSqqbzVnyRbkUEugWPskZ
iU2dvbByw9r6owrmBtmggqA5ej9w4EcndwKuSIMDbbCtsByLDaMYgnsNYLEqMjGSd8UvbqdpOBmk
s8ocij4LI066t2aFaSMu+pG1piDp/c+MBfOqVu51wgZXii/9QDgLjNQf1MDnUm2wYMsUvfIbPNQ6
1OXkiU7XTSkb4MyAA5I2BgholiuIIwcidqFCmU+JlMMZq1nIfADY3Ho3SNu175EeFscH2VNB4+Gk
qoC5Z5OcCjX48K8ZHm2RDLHgGcNDYDUEIXzPh//Fd6PeTg4DwMgIU56TLk8A5Zm/QABq1aU1SM//
JNcRItq7TDfDUP9M1V8K2qa6D0HaALBeXKPl3DjiqEu6c4ilEmRgjdzjuIJAP50Hz+qL1v5BcAy1
cNX4GlB4Y1F1KvG/Px4VjjXpjz0QMf70k+RbUeYQC+4I0/U/yfZg1vgLDx47wopnz5fEvQeW8tTv
8FJnGA4xr2jDjRnTuPxVFNxs9mbq+olWfgb6d0zzeDojkeaedDrlL/+DO/S8jr6v2eXoPDjcmYS5
xyyT/XcjZlAfGctx4DMRIE2GAkda36U4aCM8AtwF184LPj653J77ENjeFKPXJ/alnjh0niKDovKS
j0CKak5/g+4Uq2+e35EcSHKF7kiccJhCGOMWodT8ZZnaEPcg57yDI1yeuuo4shqFbfFbp758cfcf
e8xQgIYFd9o8Z7rLH4x5gVhe65dafaaH2iua9rsRnV1+xMkGg0/Jv1j2SHkPimnIsIoW+U92SlrJ
oPfbdciT7ACfz7iqXl5/zM3sp0cOgs2142UHOn+POU0n5N/BvFTw62B8Ck7PWQxU4D61pMG07AsV
On5GENgnP0Hsl3DRoC4Xt6paQe8wkxPrLsRBd7kCpkZ/JmjfyVcmRS4mEBQI6Nd0G1FIhFqdE1oN
1DS4KVbVxiiTt7gMLTh1IhBkawjuXWfDd4PfJvnRtHHHtkxnlqQbygVHg++zVgSRSwn7Z+Cxe16H
rJ9d0A78GgzcBK7juxPu1A5w4cuYGfeLlL3sdxkpg0hiTpCvGzHr+oFqQUI3roh4f2LFMxq7/3ky
8/a8U6z2XrU6FToKLo/vJZ/DsEym+nHoWG6QcaZeZ4IdH1oTmUNk2Y+uq9VRWB4B0g4Hs/jOEskd
hbCiaLvC/IgOcde6PWBy3reBzNbpU3XGtxu5rnCrJpFO7lEd4d4j4JkppNvMouci8CNNw7OUkA5n
AZKC/mAg2fxKJSDxKOsQJqhxGXHTrMay1+Wn8SKGvVGnhNfCMRb0aHBwas9aNb/jfuGa9T0rDKpa
IoK6tQVEih64QGLoP2QtEo+Z+GqH+MGqC/0GybWrSAQbNI74C+JskKEmThXO3HlqEYnQAIYNzgJL
OxvydvsjiA/1pm6gjj/df59CS9Zp4DKvrrEXeP4ag686HQHcnG/EReFj0ZFGffsN33QFqUkqDxEI
7AQoqucv5hKpklbLNo1zj2mYkkebnkGAwLoOvvtt/dmxOP7XYb6VNamcUAqTWe34VTTMFaK6cpIO
zN/TwuQx4CH/ZFaopkWxjNL97pi5Djn4VF2X+XQSToyqAFeI4BAqo1YiRTpHDMCcrQk8L8I817Ih
4un6NHWyHRio4OVkMfx7b61qNSGm6q/jK+Y3ysYar2tMQpn10rpjXLE4+NgDlYEcwhH35qEZJEBp
mbuK+FHJ5VfIkwkxn1JAEunI7kcGaaHXCfgXfwcNKQQ0SotfqCV1c4G4y6nAtHunCdKZpFqtqmFZ
lf50txeA9PxMXdvV4VrsgFCT1uVonKMezIh5+7JWk2BU6M0i7jkN36WzX6AhE3EDpm/CrPMgaNpK
jtlEFjfqRIgPNYI20sSwovvr/QFyLuuWfgbHyPMJLMm8bhYlcqfH+d3QLI+b6w+RySAQwJ08RPcT
xv4GAlux2jLzY6MEdHAYx9cOlLa0zmhy85/dsy/nlLYMl/jaxNKOQPdBGs2SlITcqNOI93UTZHZb
1rg7Lmw5NZFHuWMO+ILTMJoyTMLYxNX/SgEsciqu3QbI4PIBz1liEAUjLLDz/JJcJCiN6959xVGW
MikBpRrT3rB9Wb8aqihWzbkZPMC72bbuVDrzs/+ZAxGA+vKKbCICbwuNUTfqTVbN7GYIGe21qDGO
cFuvvTgIlK1VMZbnkQTq9bsDR99bvWSvE38QqupeubNDZ0vdaP5HLU2Zyx/OTeJrwHHtueSkJ0xW
sk4SdNyfMbNnZcg3eUwdTYTLs6bcqS2iHjquab+OFB9pyf0sDKmUmIMl71Wl5ieU4p0LhUi0gOVD
nQBgZ514vJIUNWGOJHzhK/bfTHqg8fm5pIBiudrzoP2mzFjz5ZQnkgAnXE8Cl2V0SvjZ4YFMgd4Z
RBlK/3ON6+45pB+Zpih8+kpLrHhMOCqRSQtP+bt2/s230E8AOeoFvSwbwWmWGybPmFfhT3HzMEwc
9oN0mgipD0vZjrFumiq9ez/9J3eq19EEDoQx7orBvHnmCkp9uk+F8nBEvN/YcGseGB+p0Pyg1Ae4
hWLC/ntdkK5+GBm4RLLEjnczByhXpS5g4t/J6Pr0Di6UnleTT2hZG9azkev+IP+SX3FlGpdfjBRh
SPfX+gsOnxamU7YRJhACgW9QOT6ARzxc8q7zOFtLG0Hc1XLUo6BKyrFd49EUweoLwTYzXEZ0Gnd7
DDV0MHpCDNaZ7iZcHJ7VPiBpk8B0JNgop/IEB+0HlFkTWU6548Qtp3H0992bNFFfiAqqn6uO7UhT
mLNedYlKvbHrWM7VTtyo+S6R7E83yOToVNeQYxotAJGO8aaeX5uItdXpFXSTsk4VPblxt7wJmc/C
BnVv01dbzSObfBCaOjc3E1xti7rkgf3bXHU4bRIbc/6gV//kDqezBQvXFRe7iX4yR3eJcOTitXk0
miHqQ9bWLci+xJ4Rlx15I0CDXRPb1RWCxpiCQjk/9yVVvjBZHdSf3Y+XN161vKY6B2KnjwCCP0Mc
ZXCgAlW6FdjHHrFzsdk9pZOUpjHmqmiPdL0tL5tYA8i6AlI6NZ7BYDLyD9Vz8BXKGGDu+or6iFwF
sp5hJivhUDLxMc8cwm0zdOXtTNPhMvk/8BxxlkcR9VHBpKH/K6nQQS0P59saBu2TgjHn27ryre6+
0OiaNSQcmNZrVGwgHZP4mji39OWz/gjc63A9YarpL4unkU7dA2kQQEe45sY6e82sNSrncqk97Oju
sZaueiJ2J0Igk48f7gCBetl7OHZAtPtlqXiZwOj2yZdM0Lnwoizw9yq3Pv0ot1mz80LUZL+yUcW3
fm5vCyDgO7LB1LYmfTraHFXLIQnQRa/8MVJCXENC4qJG+vNlRhN70E5adWwfwhXXN6fgCJU1ofga
Jt6gUhEWujra8g/E5qtBasjLr4u93qUrkpmPUFA7JRCbS7eqlQMsI2cGfcVWYBOOmnaFwdvfHt2I
qEPaTiwkAgYbFXypDt/sp3Zz59+1wHEVPl/1cLx4WgJueYIzhkCLqGRUyVsi6QHb1AVlhUMl8i+m
svStRLptItcC23cRvAt+vi9MJxu3jAqvRXffm9IHhxtMDEBOtWkZVmRQhRoP1CHH3tjcnpXlFtI7
M+rQ0Y7SVTHaRyUdiiawXJ3m3DveP1JDXuiUda5NKpVbCcd8e8fW3IeYaZggtUWVfQrZRK6flU3g
HiS34mODTeAQmGhypNtZ0ywHyHjbbCT6oywxfcs8cIoH57QgewnWRzkHbKH4emJTK5HkjPC0csSo
oKcmvpV7mwlyazcMH2eVQTOA/Oo5O1D9dskY9SSJCGJGRWC1tO/UniDRCT0QLaVSP57yXO9nu2nz
W9MogEFZjx6IoKtQBtGcaklYzasjSf5KVqKgaATtqx4jq12EOvDHCLeOrimNACYo+1xfByoNG79g
I3tNSgvSdiLViAyq/B5SduMCG/VfzcT3gi4GNHQYbX/+L6wOxnyRWjw1uPDiD6q6JycTindNzdpg
I53bayQ2I7oT3OKIICjdnwVCsymQVgGYC1xEuF/O564Bq/j7JOX/r7ydjCvu5FV6wNU9163uC8Vj
mOZDN9HGLewp3ynwrl9btdKlffO5Mz52Oek6+vb25mpR8aVNa1ws6Fy3Ij8YtAQADLX2ccpkJqff
SWFwsZp8vioeiA3BnDEtgjSOYA8pQ0N6ZSRFYBmuGddCilmMJSyqLMbSUCUh1emtg5KD84r/WfSG
zpv+KhFzsXp1Pg1Wkb+B/m76ZzRuXX7rPyiSpaQlyEXAZ86atSY5mQjMM7XNlgwHsQbvEFjAvmO/
VTvMh8PRDgMCjGguunPBET3z5UfNpgNWE60smQyilZnpidyod5le9fDpf1UtqnNsZn4DH1ebeO4W
nNk7BN3Sixo2kCVp9QIqgE3ytBm02IvOCcXIGntIEdLTzcFnY7n7WnsveGUgM/1hv8EkbrbX3TEP
ayE+YbEz09Pr/99NZMHOLAUxvXYfSnCbFH0xTaofvhenx5ibduwn6+s+PPPJWA+m42deluRBlI9W
WA/HDcCKOoAaMFQXeE1goPd6sihXRAb7sVZlZ0hkBsZ8fzNPv1Ysc2dtY0G4VTeR0QEeIMd6M0Fb
2dww0synivC3mt6erqZUFd4hP116dQRq5nB9VsF507Fwj37/D51aZXSyMMgtoOdhcwuwqbpuV9VL
Z3d0wE9Wml70gVKBCUqzMcc1WGGZO/e+wM4olpIwWdczP9eG9dgO92ENizO/NNkbOwAKs9OaAu/g
fQJyLGDy3iA6CQqyo3mZLZk2Fi0Dh7Isuiay4RAMauuUb8tuksYsbLkLcztQcdE5vKiUz8vh4fxV
U6C5cvKDb6FTwtLED0EZSq0rATZ2Q0L9vZImljlfb+vRumekDPhk9jq2OVP3VyXWiGNepvHIZJr+
sjgETcC/AocWY+XP4faeBG4jJBaxl+u1sSvkJb60bzhpr40D7IAkwuWfThaLyg0OildzdyXwcLtf
b70xssDfi3EY4N1cROJeYw8fjxj0wH9dwWfRQdA8zzrI9HxgNAAuZ9ClWpBvPk7x1ZgZ1/WGJdsR
72ktaSuf9Hw9cQKLv1Flx+ahNMmHL1F41nQrN+SPklG4Iexpy/vUP5zjSxJTv5LgvnSR/gTxGun7
pdGGebvSU+xWV0l9zKL2oMczyaFLKb3V64r+8sTSO6k3Hz3ROLvcl+0VWFtWdKl5R6GeKxJSoMQh
JXor887N1UKYhNlDI6aA6kdU7s4fc9hvC3wNyzk6UDuFr2elYrWeJjDHCPrisficdct2vPMqSGiS
UmDCCg8iNlyQZ469wS5v7dbDbunPJ9i+08ElI2Oy9QIIocBfIwalBX10I48oabRx9vvxn2hUaC0+
E/KFQXHyNhVRszp3lleGLWlrrQMG2GUyYDkPEkIuTAw8fB0YG1nOCZ73YIlJEFggOZJxnni9GKEP
NslfTH1XLwrmp2Fg9EK2DFuWzOXZjiVU32q2kuuxGCnyjoExUEz7NRDtey/4uk9QYvbJPCOIBOAo
K+WcqFZsHaKOKdErPX3Ga/FmOYkm1J4ZKEPnVFHECMHg/vvBQTV4jBJFsDNvQlBIF312MM40mn1V
tLy+vtBDugIQyWzBnWDP9NFhAm5XTla7eVhqm9P4oX/fG1y6ldVj9oG7TDNAgClw6ho0eABKv3V/
xEGwgckYLGzk52qxU+jYoK8lKK5pGuAvfSFsQukac4OPkLvMvO3gziLfo3DIS1e4wpwlKB99PsnM
GoMjiYS+hUpf/bV7XEYuLQNabl1OO3ZahF7hquxA7EYYWSecOAoOXh/rFq8S5cou5FQnLKSzNoyL
NsKQHo5+9VswtU3TGmHYF1D4ubQ8yU09CH49kNugLFIhZu4ULd6qI+TThvCGZX260iKW7gkZc6Nl
3jY+wsVkvoLj4ey7d+U69foSaTWNPqhpopxmlKGCr2K5n2gWNVoasrf1Fj3LI/U5HjE1mOxIZm6Z
4Y2ul9IwVOgLi+BvV4PA2HIephNgHMcfW7kYzErT9+xceiclbd07S+Gwbs+xhrLMZUcNtuSI3fbn
wdjLp5V2NGKALN/kGw6OoPHI7AmSAWpcDehM+GDJWLmL3Iq3SZgnyY6ESwwaiGZ+KBNP23zeECLk
WvLhpINeHC21qmfAciQ9f9W7dDw6z6mH8nt0Bw5neW7f0cjlZyCQ7YKM6121fmrx8T6tBtWhWDjQ
SFeKGuPD4b5WMDVR4sFiApT+QEUO/t6uxPFzu4/d75w6ubdbNjk20q5sxiiuJa2pg7qfSM5g3ISt
usz6oceHM/2Pin8PEvjXWJY/u0KfG5gDLFAV7gvdZDf1oT7I29W7aOJgftLNMdFeiAYxYRbYJTsf
WY9wN0FD+zBqdgz8+TC0xpNWPYTlP6KFyEXdGm9fuIpuHUjIJswbY3FdAmdz1aqA+XOJJau38TG6
5XXifLYuBFzVpIBqFpEisWKczcY/GSKUSC54pqq2CVFqxmGCNTS0/8lInmKPBProl5DR5K48j4FF
9nKV1ZRjntSNSbO5ix78nBqfSxpH/2EmaBWfXt4LPkzUmfMjqC9Msgy9Sxv2HY/rqspsfzGF/YiO
axLEvz+Zl1wfpdkhIipgqRyMRUbBfbHH3U8C1FFWTJ7Rn2Vv3RwvObsc46uXygFAvy/6+Cm2L6bU
3kCDo0DikWR4JfstK9jxITs6GZs1kJSb+DGSVmFhS3/Fz6wtynkiHt1sHyDwSrY+/u6Vsk03VvPE
aliN0bFo2y9+gsXGKbqSohuVRVBJh866GnJDJQtgIRONLTHbG3Spt5wauQxlJCkGepZ8+tEaJjEO
pGRGCafnFOKfKC6SK2dwohiZUlBVN5GuVLUq+rI0NTATepTZ3iGeBk1ELMS4eHNqmWOXcHpwJrMO
/xWa6re/1TCmkFyTpQ4DsuCfKVTmDKXBED1ZL4StCCa1yKg/lx6DIKPQe/NhAxMVPTY7xvEW8EJT
Gwqk1JITHOzVdQIilASgQRZ1pJApFZ4eVidHzyaO0FVRijYkp8CUGptc0WF0j6Z4YKIJujoEuPHr
hRLUpIOfq+KcVzY0CS1lLYpoPqEXzUBS2RdRUwyQYE38OpMJbUlyCAYyaf9nb971h1HNBDXmQ4uQ
ifp3eViXTor7kegGWEGt1/RINCMUCf4Fhe8v67XWiyWYtj7c6QMqd6qkpGH4l3y8rr0vCGvqh6Oa
+kQ1Fy2trb8ShFQRW1i6qR8KZKClzaq/nQXVogCVCEmWGuGI5pGNfjyRwlaxujgBS36Yv/pKbOpJ
j64AXXZH3YWnefPjR6VPbEh30mh0Ou47n/aaeDM8FiVaE+eiS5cMDys8lyx1VSNobtM0AWFseF80
O8pw6U5TzD/Qfdl4JakcGKW0TWlZDr+N33c7bFgwpESrz8MTDj64DI4d2t3TyPGBgthqVhtedaVS
CuQ3MADC1PYtfgsaDUkYonkF+3eZIs4AeenzlkxOblESln1jJiyciMc87wQyPlxU7kcA14hzNZtC
9T57AEZemNq+zvkinMbW0AhsorxYPCNC695FxtyiZlW28RejpcJdy/4M3DOUGULHEG+s0TV6eMeT
yD0gDMJE8kwtu1iMEmj0+anYE7Thv8qF5Fuf35xT0G7cqB4h8p1UJienn96QQVzzzI+5/Smrq2TI
JQdDDEa94kaSDDsg/S/sZ5BtFvfP5WpxLMms0lk4fBj+nS3A/ktDvU0jdUugssd6zo4KOLZMTRB1
Pomrhhex0/FAw2fOoLFin2y8EnAZ4mqW57YSI7CjGx6yn0WcQDKqzjoVF2FWrHeoKoSgIJviDjbV
EFXdrBrpUW9LY2/Ns+42cKovnYAo1WsNYDjxzJ+Q3j3KmszaRbYY1zMiide46POr7o5oJ2Bo3DEx
1FfO0DB0gHiNqQ9K9JQ2nC6Xtl1BbVfXnymoxsNgarCKERm/geVab6q1KGkJkFK95SAN1ZMzCwU2
N8iCQ1cmuORHbuYaiDWt3vvUVgrRpF8ovKkubtl4FcwI3haNijmXQ5R68VcSzpyFkSCWVQhFdZ/a
w0kxebgmoOP8mSxXfscfey+GSRrDFkadqYYgJcQtmeiZu9Q+KsQc+QiV7UuT+HT3FSPy+Z+2LPgk
ttPFkGNzsBgGn7ZN/s65/y/etzAfzwWAQvVjhE9egGuTofqM8D1wNOAqw3qNddXVIM1/6nUCdEWQ
jXp+jKMYgRrXIUtakgDvYGr8LrWuHq/HBgdBlluaotCimnkvIq8Y0DN4OcJGTgiU9rwDV4sR5Dp9
i/hpMzvxKtX4NUSr2dUlIlJPAbYdgkqymRVY70xjKhaM73bw/lXtiP7FKM109lSyRpVKRmRrVzzU
hmP7n0ylC2MK5sxqf7Ln2P/f55zt3UjEKEVvzZimn229NTWuBnVtQdnU7JCtQkpNr0Cl7EjW2cke
Q40WSGjfNZ6knukCm+QHqKTxh3WKEhlYwzMMHhLZSVCA4JLyIdQr3mGVRmLXtaHsWJ4cqtZe4V+Q
wydxu+pvyv24xvxicIFzraKyqHigAq9SADOc5xCqGznxh8LGmJhA/gkHtKoEC6m0gd6nYlZpJfAM
2o3btS2nECld94LDU3yAmbg5CpXIIrMfPPZRUW4NDzxEVSquVYvJHDH1VqAo9d73zoDFslbPPaGQ
8VhmLTYAWe/hD1UlzRZlqt52DkU0McAjTEFgPu1dNjsNLD2xOFq5B6v+oaz7bj52TqMmtr6bLtWg
xSJow2lxZJzq0lQK56BZr1mYu5blLaFKv6fTAjH/3tn+p4gDvXJ8asuvLfLjaJ2276YH5mfTpuIm
Mp2Q4sbXiQymiEXnH5fSHjGWM4sfYruVm8BAx28p4Ypz/YMyKoBlvGu6ceMmldnwXPCPkWjVJ2OF
rTu8yGIduKFT5dYpUOxo2nIZdLhaDOYgwZvRTDYj71gDIq2FkdoMx7kL6RUXjRVWYJDTPymJJtZe
TM1BNq9HhUzA1fyF7tAmAEF9UPZpmNqJHXeXLHJ5UX5ZDaXZw89byzmz/aRyBB0mH4wtNIIGldp5
QCEb1ouYTTHWaJRnVLsdjoZwIcLih4W1+bsImUd4lN+ymPKJOcU6mov7MAsDygGBnI1D/lq+Oqxi
ItbL1HVRSJsbceLQg8tQs6zj2sdojqv06pKMDWK+GvDLh6xCt8pNpfuXm4wspqzY2WMsg/oFrceZ
Duapqeqh/GE2GcS/5Zz5Tvq6kJcWMT2eJDSy2tQuDV3Cf5OWB8a1jC4O61JZjPgA07RRmlgGwu93
DqtcTHyFwGDvysArPnmfPPYVsJ5J1tZ4Esls7HzYGmdOb7GloNMgwVOOIzha0Xx2ex7wFLpnQ+Td
vCkVxA9i3idYIVHnB83qLsKPMs6rjGDfKqlMxOZzkFiXcHBd3n1z8Beik0yEQ70nk0F1zwc8TkR5
gxMp3Cl3bNuB3uncS0Ds3ScY33ZC/7jBwJvPNAP4ADv8+Zp6JsI56QswidCaNDrXc4hoVsEan7xT
GAn6rifkbejz0Ls4SCzYF/MTuT807EAsOAjw7+QyDLCMJNVRg1SIlZ6LcDit/sflYXc/0pjBQqi4
8zT0jNunSaCrkTym1aQZXUxdyF5RiOYbN9+dYfwf8vnrU3/cLHFpxUOJ/OLJLOwiMjbWzXnS+/Ki
m3RAzlZUop8TdR7uz2nJ0peVjv9QwcDIUChzZTY95huEcymAekNzdEzm4N9hevWfUDWZxGaDkBXj
jrRNCaqGEoDFugE1KUnJ2Yv+wl0aAxWExOKBtTbk5fFEl/c0f1DZIZAnUBmAg9PWE/wGDHWDP3FL
6/o8LynN/s+b1BJGmZELI99ocv8XPibz9VR/0tcozx4Wfl53Hy6iBGQhszuFDa97otG/8NuTH1eY
SWRwRci+IBJLB1z+9MXBZhOtqvnDxo3CVGZVzCWLlYY5GXrnYW1A8ZW0VtOAVKoMMVdPctpE57GH
Nq+PM+FEq1TnLLz3qSpRvYFygrj7WpF8XRR52j6TkMAsAVBp7qEQyuxsSUYORnp+w6NBzXhdrYAa
ETbSwVZHtBr5H99KRcoRjrdCLvXPEJBM+rQzt6RFMK1t1x88mJ17iYSXWwDa+oJAEVvvyiOq74XO
9IOTTd+DSOnY7C6VqehrKAfuBFt2B18XRHZl3+oncovPcymzwIyAdWxbdvGSlE3dIvX5sLTuKfRb
d9muC8jNOgywhVXiqz7/2oD8uw/0nQkzzmfvvaLg5kzoNrLh6rrIvL++ljdykkuHgg1uGQfOsSwK
ush9D7BjNI8tTYEm4FgoXwlrgS6fWHkfWUefv/9+NhnEds66TO8bny+nOYxSnOoboOeNApozfbDp
91NISjkzwfCeHJbYAAcwhDBKQlFbYZ6ESlriQoLE604BHM5gNGxrjuz/Y4uEFCPTI6XDs9IJranl
SOx3y4vGgcE85dnSlBqOhHYpgsUL1euVQdKVBCdeqWeNGDWNHWhReASixQT1r1ijy71ExvAUemB9
ukLdtlxk/n6w41NVFgk+ObsNsDo9E+xH8SQ4IaYqQgwqUh2fPQ4nnipfGEQU9iu9CXaXENYNNSv2
2VlfhimKkobJRvooiwxq0SV5TxE9EpVfbCc/8SrK2NwWzEcZFCkgoWrbKrh4N+pu7mMy+Qih/0Vf
/67j3+dU4/SA4GqGYdmnFYh4N1Ci08SDUrp8VKxVUo5AOCqyWy3xtIWE5vpjZq+cdRSKxepN3v43
ZlW4a5quAelFQwSz8lF7W3new6TwPBA7aIApLrkwlZ+g2xaPZr/sh78bcsUW1nOvRAIII0/sKMSI
Pgz8/CDzavRQbC1SUXDzETCRK/YmjuvtWh7TYrQ+EVhTN3PNbs5NlTTIgLA9XDZG488yZalRgomn
3L1Fk4Z/XIaNgyYzNkXNUf3rniLVJ6sx0Lbx+t8w6f61IPziV2++7pBXZ91yGZ4z1Dt+jiGTzc7V
BfW5bAB+oyJHeb0ZAoWm2ozonlXSHvMMGyFxY1DdcwcDI6RP3CsewkyoWbCUEAeY2okPZI4FzHSe
cSqNl1M3Wnaq0Vg2iQ64q5satZyAsmAjkfk+SZYeGJLaFBBel+NIwIT8IOSvSJKecHgRRWQtr8Fm
22VBBQqcGl5PKle4jEKNGUY1YwURhuUkX2qSLRZjcMRXnF8EVW1UosJssonbJitFEUA36YjLDgHN
4sHFOz52IRu2wg9ncFBq+vwj5bKNXCPyrvjnwsmmEmbxiKDdwCnY+6OUN93FD0fy/wBS2IDZdA0+
GtIvAJNK9k8kXBYD/8Z/gCCwds0Lk+aQqvw2b2jSQEJkZWyCkNXSGov35zopbDTExxj7r5DoxhpP
GNgPwag6TnLdAQH4L0blLWsimnDtBtlIGIc23HZa1kl2XOz0yneQIeauhydW76VgXQJJoOwqZkzy
Bi2/p3AUruunaXtuubIl9iwIRoubcCsEHKvk2V4G3wGdF5jNgYJfZmjwVBchvookdQx5e2fxn11B
hCOdZrOxC20w6yuocHskn2FUJVpAH36HUsJoshzevMg3/hXi75YcV6QyHSNrlpVVPWtzqRjI36uf
5xFrGSQKSOmuIwap7TiEDWGBaymYVIa6KTF53Ywt+0Vg6V55yR79vdkOVXZNqnrWSdO/0ESuhuUZ
6PYAt9SCLm8LDIn8Dbn5BQvYYAeoqYEj3vv8zz0OgscXiHD7timUCygAmc5k9hyfvuMZjouCzxFL
7kE/rT1T1lUk6lzokPobb2K07hCjrLv07PxwLKSUpeYvAOoNo4YTre57RSs/Z7bnYwdc0/Ttau8R
30jQko9MpkH+WACjnhdpDRu0caP7z7nK6JHmfx3NxgBqLpSfqRB6rE/mKZYY5FB18j/lFn7RIpqD
ScdV4QYwJQadSKd3lIRWc1MPgohsvpy+Ct7S7XoOhDlRnzBlXuoQoP7KlgEt/aurYmIkWx4rlFcV
CehA1Fj9w31eic4SdWuE4TnEgTRrSaAzpLn5na5Ol/XUPaLZL8Kca33p99JnrTTtmfo0NwND2pWk
rrZGVITnej0qhu8YqULiEKWyLROnj6DjKTqitrpOMvW4MU2ZlG5H8zCaJpEH+dbNEph3M4F/7RPT
TzjR4xIvPGJlYyogAuL2X2DxGiFkHKxRivkDMBuKW+8C/u3fvVs7Za4sNDfF9RXMnXtQhpY1Z5PM
zHDlHSR8cNaCcASOazoG//uBk1rRgEjA+5q25fn4apvnDp95E/Al1AtZm0Lo+MSdyl7Ru+fkYNZo
hYp5ySgozDhCMraGfFzoF3vESfU0BBNQn7aKMrj6HHDc+5LI0C+NkAAIDfKlU/urfc5mR4d9TE8M
Botup2dBp9APA7u9yoivdErUCGe4+iEb9M3g+nIIetn8S92ReqMwzOPw/3xLISLKPwx/Oi/dRkQk
yJZ4pFUs8ET0UBXcJc0qqYsXQq/lRvVr2vd1WgkM5qJice0oytkZfa6D7N75B3age2GyYbuSmxc3
mnbwttrMb3RfLUime5KuUw0kYMBnrsvRKsl4uxhv0ox12Gj1bb625qBWONsz9iIMUW7Ry1em+400
+sZ4LSO20BZYj6vR98ClITkNaOGADWBJyenG1M9fpNqM7NKFouzD7+7vfYqn80XFXkyLDrFlKwbt
TKbIGVUcAm39wrdZ+rgSJ+fHY1uZgwtB60U9wOnACadlGlOVZQeuCEMcZWzDJWi1KX62Wc/Aclbe
d/vqNGZbfUrYR3f8bdXcxVGVBih6XfwCeb7vz5f8X72ZKce/q4jOqWhW/eifywvJlSTD+Yjr0miS
UeiJZXpdKQLTmQadzope4Ea4tTrtzxQqLlo/l/ybNNwZA0Et+Bd66tluC492bHRzC+NVFa8SpiPE
7klQS3nkbFUUeOHMQM6SMjG59T7PbXwFywn8AKvj5vVCpP4Rp9xtRzoC+qaEeRqGYr5sHrSFq5EH
opRhg78GrYkkgDfM5M4yaN+Uppx5+TsU8oXWWED2dFrk2Nvfos5WGbQjNIWP1enYELwxd4JCzV/x
kmlVshYKebgNKtI46YJoLgvMoz4e2dztGCyzGeRPa1smtVGWg1BY/o/49z0D3GKMo3nnWM9bmIy9
WlNnorfA2fqPB7vSLC1txAyZUSJ1IRnegVVSUbOVS/BCQwg49WEsAazK7j4usdnnIa4YtwGmYpvL
qpXrdBjtyys7siWJucyY4BTShz8eEHPdiHTh5i1DiJEudQEikfWrtR+QMr4LYKUyA0771zUWBLuv
gd/Ykjqlpm45eD4NAS1g3f0a8YIuW+3RtuMG5kb0Aur2KS7OjdKh4TvFKfLNedIXIMfGyFKP3pIh
lUWsD0UiaQIJM5YkC4S/YKEmI4FkX3dgl2IONmtgjLAO2iNp4p8YRN7loiiSfezQ0oIzGxf4XwZn
s5RMZBsk2hjIBJtd12qjQUzV+4KSyKeXsKZybVUj4py2YIT9DPu5JdMxrzi2iaTnzwgvp8Fj7tk8
siZa0B7sbhq/gpvGSFFu3lewJv2vOzSlLDN9JpdHUQQkXnlPuGkuBh4ag7Eh01s0rqBD91Qj8KyC
qsEZJBmuNMRe2Kk92SoSaWV6+DbXZpA00CBs6J1mIpEIbZZ1bOiG9EDmBgLGQPYQJvmO2DPFxKJw
u5vNwc35UfQSfdV85+rxSc7uEOkuIm6ixtaDk/33icgUqpZHIcjljjgH09G0F0T3I+GkHJTyEK3B
LtwuG2r0LQvTYR+IWug9jSrPd1huWvyHhV55MM9t8ER1aj1bVXToaU9nLwEthqGdLAG7/m+zKZOI
haJeZ5oGA4jfWuo1zbVlxu3OJgdI89vNm58pGh4joDsIIciIUoEvTHaDBrJRAWOCfA/NPwRhSvOf
64nPaT62kliyL5rjPGfzRi80PRGARfXfoIIN1xFBkMSuKXqF1e97fwJb2RchKNev3xjKs0+Sh/Ce
8/B3EIf5A3GoDBWkO0mZ/sypx7t9REXI88tbDSFe98nW/1OHhTLxiAbHTp0rxMMUWVSmhcTrPZSZ
RSZYJ7WD01FqAE4OpMrSeLaj7LbaBDuYephJEDlq/Urtv3m+LDo2NCHNZNS4cayWkknsCytUoox+
jYSDkoRVaqexOSNVqYq22cWlr/7Ef3D7sVuju20vIPAq0af+6z8dL24iGIfWiI/B5hl3GiQ4L/WT
YzbzyOMMupjIC60NC/zMjlJP2qxT3k8QvhUpO+4Jd49rCH2q5AXolaST/p6eeoKV3oVSdcvduRqW
tMG+tAxjnrVmdgyCxN61dliyIzVHy9D5Z7W16MdhTI7NospCPaYzMrlFnyIs7Sh61ByELfvfQjLD
bwCvUXZDRc17pFtsYMQoZi3qPjYKyhx4oL/7O4vuL3LsHIIl+oLaCHUMwMncd9Xyf+/WKzUgszTW
AQ5O5TT8Q4VwWBEcHhhoNK7jKpXC3MDQrXn8Cfy+TZCT6ewxHZ09Gv9DWc8PwCoRPL0nUCud9USQ
Xmf0+sAc5dKGerYdDjGb3De8+3vY91NmSCks4398vHETZOvKIYos0VDxKG6DF2mKtMwpI8nBvUYj
HZF5bUdoK4rBP2IfL9/ruzxu8oAeCZT+FmOOiiczg6vm0dxJ2BVn5vasVWe3n/FTcORYPssM69d8
b/n4lw3BYVVSOkrc6mMxizvWSe/JDYb2XC54U9qtJea7CyeD5lDsy0DwxQug1q2fX4urDYY9o6PZ
3l67wzG/M58Hb4CQvv+cNVZbw899wVy8n9v2fBA9onGbINWCY3X/0rKtTyePxbfcwMZ4AzRjev7E
3LMAS90Wxkq36NzBEbS/a2MzxxAAQWXq/XV9Dj41wL39VGq8qMO3xLjckHX89YfgFQlTKb1detO8
9uGgbTgj8AgBRjyJdmqrp5/ssJpd8u/MenOYIN9rvmoOseOYKKgGdxcmYwLtOjKZ/9Glf9bPcaVn
6Y5KKq4iZNIX4LPSIp9zyhOPeW2/snTNm7cP/k9Tp5yAfnAVamDO5PczDXOo9eOJzwIlXWDLHZ4R
58yP+hk2pDeihEb4TrxNn1E+2riVjX8T5BnikCLypbD9RSpv4EI1A/TPfTeOU6HkFo8lZChmVN8o
6/iIyNRvvDIyv6xGD8CM4LGLUP4Xh1DUzMHDpScrFl9+YLdauoYGWW2X3q9a5C2Gt7SHJaUgHdnu
fnr3jgds+oTOY3jaSPSGSf+c78li2XXibQc2aKvTpS8yu3xA+4tDSrKFxtmc3dhuRFv7djrx6pgW
mPm58O2tb/6wjRt+DAoZtOhCVOcfgwqOzBGHStizMtXfB2dTDACF04ucfhdX9BClySAsZ/O42oN8
5Z0JdG07GPjjJrfnEcl+1CRH8d6Z296c75QdJalmPHHFy+xeGR3GBTrYQvd1KcKSno5JX1l8Ir6m
CouFh6ZwdodqwQIMHjONLgXSLGzqJ3f3T9izFqOgpprNakorAD2u02Ugw1qySN2DMuX+7h1KONLj
C+Z12TMehWZUBgxmpxFuiNej5knJanKF97A6gTCIXcQOwD9J66U5RHcWVnGh3RcTYAbCsVBzFw+v
E/w+maLjPV8HxXJQ20tHMRTSjtL1FtpusTgqjukT7ZOxv1MK/uOBg/c8xVwar/ClLDO4xhwp6qzO
8kZVntFWuo6U4scELC1HcTYqp7NT095+dtsb1smrJ1i3bhxvuP/njZXpdNf/CnnE9QJ+DbSQ1ViZ
OWLDvG/exh6WENirykQwnFqFPe6GSHMV4Y8fpd6AeZQsb5BwGEwwZ2fmGzaOWFW2id9k3ne4+yOv
tqhiOGIzKTL8OJO3t7tD7cHhl1lvd+dGZdyHmjHnJXQtaXRJZjpyWve2T6HvvNqlNnbEKgYRnrOh
WY14Bl33boXHUrtj1aHp7VUTx+t8rk6exsbxN/q+jxtNwBesDa8puWZeIpuK+a1WoMEd8UTPWkTC
6ADLkXRNsxlJFfiuoG4T/U3RPgv7K8R9HNTaJfPh7b6zOlJtO+uyUh1hvL/Th/YtVuWG9ES+l9PF
8a5KavKF8IcaZ2xlt6TlwKpqcmlmn8ApwXt0ZrutY1vpBK3UxYcITlu62Vj8r5iZJ2Vpz2PuCm5P
UQljsULc21VV7dhX4OhFigKbYBw9saLxosrX9sul3asPOk3A/x7/Hk8hYD4Z8m0kPk+JSPbb+lUN
qC1oW64Lo4nRXi7orNK6mmcfiOJ00ekekXlRS41bbbMC2OwLDVVYpwBe+ReKL9/ZIbYhVhaqHB3s
hvy9MW6ygHm49aFFIxJ7fts9H26Pfdns4IlSK75MtJgUWUtvpx65sggfmNS4g3BPNZ7elS8K+QTT
JJQ8VUe41hqQmQl/CubN1mwUQ/f2Wi8GL/EVgscAn3ArntS1rfKT2BZ1L36CLJrKkeYJAIL6VrsZ
ysaS9nvZwBkjuHAnxAudUaSuhqw/GzbK9AaJeVynS4Na8nsmv5eiMErE6IrQFkuPPDBXu5npku05
nDmVgmWT+RQ4bpIc97XmAmxI+8UU0FWRGM7VRxy82Yu+8NJANuGrIyeu37O/0mErifBpGAl/V0KZ
WekJspXZBpI/IIFwlpDHaNzHfKplvwDMoJJoJIPmWD+7fRMHe891fXP4YKPAqpLoYMx0G1iiyd7j
N5OelnGaMQ1ZMXcp1ah3qfd0QAZhCI42Wr/y6/Q9vR/MHBNJSZDxs7xRggZVFILinM8ztJOEVRaf
X6TkGkeHs5OKiULK5/Uy1Pfe4wYnNajMun5Kcu2JgsuQE7+UA7TNWiwwNn/cBsly6j4kqBP7fCEd
puOrcH1fxR779qiWq8ygzqs/I7eLu4Mq2BC2luBOeEAFKubGIcOKNTYgZCfKZfP9CIVtN4I2mn06
PH/eNdwo3oA7Vl3/sk0fhNmLOHKRkZaLxm72uJrOoeXIZoeoK9B1g6zfwckRfq2VLmhDMcNnjWX6
PCYR6L03f8a9zY7iVV9qFbeZl1jW/WDw4z5QAgxw59wi8dnSh2oC+nAodJYqknC49f7BukXwiDaP
sOs53ZbFa8aAjALgd8OQjZyCJ0TEVxpUEMEo13Y8XhnDnZLcHklxicEPcYD2ANqEAkrujW/l8CX7
g87j84SdSN1H/xDEof6k75d7mGidNmlSvffOLb12+GBjxOyfGY9oLMh8Eq1QSHBJcKzBcCSZbezH
JRWyxJX1Mr7TJt2mjft09Jl554lvgXgMYP01mI6zuYUzv2zwkOLrqhlpjoDt8twxLK2h0xStL/sn
Y03OknePOERbRmTM94OTtpeWXyY7u/R5hScZXAR7fNJ9ztXxqeYtCMl5ObAnoYyqBPGqoItJbxpt
q0ND4dScoj5QY7D2KdgyYY1pR7zWGxpzs4KBBSBs8feZK7qRGKT1C80N06nqpmteH46jxrv0iq5j
g2UUHrz2Q9Nmkvi0/+nXRuUir73hLUoIAPzAqF0Schv1wf4oL7Chs5hBR9TUM0lSGadww8lj3Kzk
t2Rg5Rar67tcpVZOnJoQzRhJNapiaqy58cySMREeQU7IIyPur1ey1Kz0bWBZj0vD4amZEM7PgNG/
1Y6l6CS1rnfP9UMt9Wqdsubebgj6A87R9KhWjWuBbTbSXYUbD4EtTnTkxP2Iq0YdBnvzkXGN1/l2
XxJQr9zvEQhkxcosCRy2e7Buc7sNtNNjD8SXqs20Jrw3hE4dRmVQ6eKLDI8JG7Xfc8CUgwX9Bpig
d4AXMSEvbAuHVw6iLn2F1dzwwfpC216213YZOC2UBWO2JishV93bXMCWmcBMARtCIJEZurxe2u7X
vjd3oLUXOZznmcWQivXnec2prBhcACCgzCuiypjJ6TPtpGSdjnMfIL/bWjTftF+1W+Jlvnd9q8g9
5IhEefwaDGoNrasIaiYr5M1LKlgSPcC91zGR9TBw6vPlN0PC6jc++NY8eXsQBsIVm5mDbQh14tqT
0MMMjW/iKSVByWOcJTGddyTXKDTt6nbd637R8hwev6vraI22+MfDYLWj8M44cPWzd6coNQdgj+fH
y+BiZT5oHEQRhIn9zi71ukztf3iNdEAHKDbdZO2TSVA0LcQLHs6yCenxTwSeEOhGCiUBkcmEU+ps
FfTn5gnmCCcqmmaBvy8zLiJ/wqaIKSgIzo2dQFVxQ3IUOCiacT+3/r0Jm/G9m21H9OSdUWC02zRA
0P7ZOIc0kEn42YlKvp0HzqU0HriMqBSx4ApjgWmYYJYonHH8WFfjbM+WaBzbDMIOMSmR2P38h75Y
oqsFJj1gAY5AVazSTCPwk+XwoAYiKSf6xHjQrVr4ZG65JQta6MEJMB96VVQccOOuxElM9qi2eWlo
B7L0ChwY6epax+Vy5TnYd9T6FNJVOar19lIlsRIghtijHmk09+H6mH5gIAfw0qtU1xQ9jwB7iSH0
ygUvoxJl3+V4TuXUIvCQ5iPQHo05iHH+yZBEyt4KsMx7XHV68oSdhUjd3D0ezK0CIKJIfsttExiJ
t8sxg/MW/fd+lZxYlbvOenayTAFuyLJD5anTPL6BZJJyYP+XK3U4F3yLhGg/FRopTKhgkCrwgctH
EEAeaWRr8lUQOod+lbEE/rU4TB16FdJe0SpRmS3J2xweTL2s/7jTs/rT1RCwrtiURT73cBYfeqZ2
Ml+oHajQjNut0qntlBZWno8OuwGsHzqlGVEVux/ZN0ZxWioY+zPzS8wyCMJJ7BWo1wcdaqEkWd3u
b/wmKgA1gq1fMwlzjc5Az4NOinUDjyheY++SMB+/fJ7yd/uwgITxEecXg7PR0S6QGwDILZnmsc6K
S1j+TPVwbg8Wfz+Ivm1vA9gMeA0MP/630P1faKLVKkU2Km5WJapac0kNtHm+H12rfI097iGERVEg
bernwcDTKJZKvfvqbykQColCjwmoj2lUN26vTpY16eWC8yQAksmxPJ0i8CEjU9YhiTn/vX7Skeb4
z3jr/GCheiMvB7brgVa7xC9GQU8nVuIy/A12ex3X6qLagf8eu9s63xPG97Hx1XmFQUPAuepNQ+Ux
MOvTRfDqpFuOJbNpUMKCLgpxFexoeoivY+55zx/mxhXyitQgI4ul7FHFrTMwkgW+2HvWYT+4QlBg
lJReraGWDsldPXpPItKa1BIeUPcpdzwbSNksquEW+T9zwru2OfiTIrJl7X7PzsE+mQZcW9EafcIr
5eK7yTVbi4NBAxKFHzpglUlihEu1WAbJPbu82A5MrJhbfKT3iCoT7Mu7k7Z9c97C9zEAiCRTqbKd
9QgwqmncWjMwYzpaZnbEI9htzcOK85vjFVzBXVcqghVRpbO11Hw3VzczB3xPI7yM6OtaEYhiZNSs
PjMfkrZh2JaihSyEByVALwNwb1NSLsydBghSRGPjAbBdtAAxDlAQMBt/otS97KQaG+Ne7D8HVxoy
kYgHiKJ2vqiR38Y8E4JHzCt5pS7vbUOrLWsCmcYZCTf6AgUSq+Nc9o299maohiSWaEbdQ52a0zXr
A9bgTdL/oQRLQnw3+fUOZqvVrC3SNiB1boEOYcsLtrfV9sjA02+7EwNyOLJHY7juKkK7PP9n79N8
l2lAM3PX0wXDun1HIk2TLOtPP6Sq9/701q0NmQVrXcPaOdkBoVVmn/zep0KOwMNC93CHpEURWyrN
h8tAbTMWO6LP7JN167tRfKhgUX3ynZ4vAczjsAExYdYqC1NVKuuP3K2kC+K+lI/65lLpXnzhZMZE
q1JZBw+/zdUc0t6bLMheyHZ4KqoW57Sxmxif1Tv/79pHpl79MmwT8WWjihnmT7gaPVAiBX4ICxzx
OITHDRmJMqUSUXEUBZIUYmk6v5B88ceQnxO/XklOYCe5DfG7Lo+YRGzigwdLk5hTB03mPRXrZR/n
WV5EV8vITzIeEC+CkUndZPrRqTEpl4Pj7DI7a2DzXO4ZNNmKKr7FVs4SDc0gWcqcDCZ8kgucdZC+
BChgZolTEvHyh3a4EeT0PyqjcdenpeJiMoHu/iG4Dc1oOo9tKuNXusLZrnKItZvIemKJaP9MZpJn
Wu0f2XNjxWi0pWa/Qtd79l5y2R66QYLe89/xkf9+4Sv2G1pkEMh6xtUS+TzaVdGiTicPpC0PogN/
icvc/P4QUcOOdjpd5/se2S4p/cm0JxFK6RHtwNx9FUszTpSLLWH2YCNGyKOwzM+x1qqXtZsqtoh/
I1fWvSThs7NfKIEEOdzojcpRdYrx2pi7qwRmILBm2HdK0T+DyMHAE0j1m1cJjJwZa8jxmmS+lBlO
e/Y82rtnKoZ9C9hF9DkRPzLoBj1nsNB1pq+2VOa2AT9Ow/VRGuIi+q0m9KjgUi4w5uprNws5s6bv
YcMppI6DKU/CNVkpIJkG8EewGEM38Vhw9AKJXNq6xLtiaVRTFmajUmRI8LuKomMaPA4ulVZhW3WG
/wnArQyvS7JNiZESYgdgAWt4VW0CdSKtAHCjwMNC+K6p1H9Mbdz/7EwspW4hdQNhfYHAE9jRneEN
ez0FNcipdXOL1ipE2bkkIAney77fOcp/N70ve0U+Hk29MY5GZXDyRLj9d/bPlgJknhmVMvxbOuvo
8Ok4lvhPKwGAGJ0Iff+7lNfU5w74wYupBoqcSBjRXGFMmwZMoVxGKeUyIvCCvqAadcxtsjUp21ug
RUihObteQfTAL13Cf9YAVf80yhAyzh8D1ibVe4cM8UjAm6XEwoQ5SHa5AMAkLmnGusWBEHfZSDOA
iMwBc2kIjeiLUrKjzsFcbkSrjYBu5CaMxccaGltdEH31RT/R7pLiDZv+TQEMqYUbxTzKW6WeMCoB
RZY0ZkAKAlPfGBwruywV04Vn0qhdX8fPF+5gRyG5HjplCPj8idqVbZ6x75WlzR/U7h4N/aYkd0tC
miQk8r2tAqyUhWI0q/5ugAX+46OLUdmP0dIcBq9ZuWo0uoCmJLphbmnL1dgykoyGo6yfCGBasmq3
+6Q/kaLmy0QXhgo571leJD621c7YmJUSem7Zb9NycIfNzVLI8K4Tyag1qOwVlNxScgcPU0Qanj6X
2TsI3XRCTHcI5DDU4LPlF6d2oFuMqAc1OCGx64O6F3vgIh6DbwZaY9fyRnP38Xb/60a9uKxpZ3Rn
Q2JbmUWnN3ZbKiRxucPhFf6qL+7grtX8he1xA7WTkFEbXGw38iZZy6VjhrtWIeeElnW17+rrClSs
yrElNwnYFguJpSaO06XjhrWf8DEBx+4oIKk4KEOSRdMlzl8Prq4hPSvu8hE3npCJvDBbNpxD1Ziy
I7I/Vh4Oc/KSfgNWuVsKQo5BPRxQ8aE5wn+iJnt8syftE/5/qLNjfB/CkkfoIqLuTEUtkqaHxCVX
gxZGeg5Ha7Yu/D7XdBPqgjSsfUZ2vwdfIn+5ssd8uIC/XvOJfgZXCbxZ9K3ZCQqohNe71yKSqX6U
BpetgYQoDR27qenm3O+TnS+b1IPOrWXPfU2DqnfFlwrMCrhsi7512WKEZqFhwnBkz5/zHEy8NXHi
Q5rysbhqyMHGwqjYBut6DE8PbT+hlRAeC+/n5JGfcBM7YJFPt2fXl0/3LpuvEIjOc5PAs8V7p7pF
IRCcVxV0cJu7fBJyFRKhPsMywDhwQPIkhZLEKhQjK0BI3Z2YvepSbxGbt8fDZRBenIuNtK6t/Uix
eGxGoSHJ0JEQR46LqJRTfFot1yBgtNcAP8aTe1tlSemRYbxNXirFPC8oIIGKr2NCoUy+ReUlKlj0
tQ89B04Qv3o+PB48kdofaaEEG1NZSdfklnHHjyy0d/1JB5n961Y3DVxoWZ2EPmIksM+/wDfFQ6w6
VuNaPmy6CpeQ+FweUrFg0dyelJmrpEBwEmA9LVKOH3kbyCBOBFxK6rzFM6JkmDIVwGTd2E8adM3u
QeQoYh5vPLKCOXTGjfDJY0YYoL+xpuN7rFuCFFRoTmlPjhkZRBqZfi7jPelGYjjPdP+oKzxpbZqP
uOmideOIcJckExgYoTsKCJkYVNQL1zK89SIPWXJNRpi90zfrig7VPZ/oZk7yYHU3OEPYBx2ZL7+4
FeR3Xe/JMaN/hk1khwyi56Xg1HfaIalVIOqMsmWDZPusnztGbwnDvYyuyWFvcO6m+YYge4l1vwTw
emyEr766fbVYeYu6QpQi4nZ4UkO0wOo9ujdtmhReFERCGxuUKzrqPeBo2F8qRcQaZm7E1y/VnyHf
xxaioKqp3IrcuNEakXDnLAXqKfzwTKNNT2tr3H5HEonbWoNA8lg7bOzh0xTHzyKNDgohlDASwktN
1AIYjd31wIWH+rjmBPZhtiqbTU/AwUxUfYD+jh4LOoXvq6ykENJmsT9964iRQBWpID/5xm2C7xgM
js6YW/mDh+spI9VfsCPTeP1iqzlSOKNtUPbUBvMINW+XnRs6shmnN0uyJjYB9OkUsGVeK7CgAsiT
fHlOXiCunEK8T9zUQliVTHiSJdRSL07+7ycAAM46J40fRBeLEzx54wN08xHMidC1PhHTeUwuEHna
GLwj4tbxRsx2HzWpknaEreJgM4fEce0FR8gh9twfHl7yDOPArWrVs6hJRCtpQpj+Zk0z9GgbXd3l
3wahrHxEZDKRvDXeuk3LvgenjwEhqka+KuZIz9huHIpnQxgHuHI6pVhFTdG6iWHSO475RGIwo3+5
+h2Sk7RoxrK/9YWgKspQ0c+Q7eLGYYESu14fOTFgXelIYtXkMN36B62F6UH+vj1qD+8LfR0GKXMZ
kEtdiumgyzB/Ids+iAiQrxYuAzAb3Q3MzOHSPirb/o5pOJ0jrwD421CFi8gNvcXpzM6LqdlNTwBb
mrHGSHmOL8c/apOVTy9LpBOblbtqyRA6jbqNFT9XL6D8ROUxl8+xaSJcZjssdi4ptCl1OvPL0u/F
umpeBNCfaLzY2kuw1gptvIvQoLyTfM1x7yRpm4BLesGtgFiNCTG1CdfEifoai8k/2Lvx7JGdP0iu
nWsyX9ZU0tnsee7luG/nz7lClTJD89V9x7WrqKSljByvj9C9eZqoulH5KNbbqsRMdasaDOwil2WD
Vh+vINRH2rEdJyVinHTSnQO91ut32auRcHWt/N+EW+rK4/Z2MsuJI+8Gxnxs6zi5BDg1dG0958Ja
mjNc0mD4TEDknrTAgLynA2KoMEYO/M8vfxKAmO5lVIVXhwLzSNPwe7BQQwUEOVdwau0XUt5JOPI/
BFlIIcK6XGBigdX51rXCnrewQQJQBP/c5Nc96rAtsSeaKTSoMxzKL5p0gHEbw6KOT6Sq1WICrJHJ
5X1h3Wv2vNWrIDoe9s4Jefa3fJFUcoJmrByDspQOIaXdWULZZfRjbmOqnCf4ZvGZ1wR4kartaewc
bW5O5ptCMh7QZO+lYa18w5lYfqyJgtovCGdCR0TdR0ZlRgHn5eUIfDhlGZNh31D8Gz9PaAFEiiFE
RjdvQUsqXlcgg7OExnnlW5vO9flnPe9jIpet5JBy/paVUEWGsSh/8WcayponqUM8rtELsqu1wy9a
paqimCQX0Ni5K28X3uUFhRDIVlGz+UtRjU7O46TPBfDuhB0yhwxALkvVV0wcfcgYkesxtCgSrUKq
ZCOH2ouA4gD1xnfsGIe0bgZQM6Ink4ttUexCVtfYI+SSkFSIARce2803sUmqobdoyxZNT8HSDY7n
vC/lepLK2ALi+OszuTa3kwV6Ov+ZXRWEabwaj75G5JPmAJZrW5DeHdpv4aAC+vaqlNVbgMHcFXrn
fyP6XSkJU4rxZ+qsBsa54mweyvm0QftNCk85FDFBQ5yBUWIFNhMKKjkCmo3ccam2EEz28QE8n0kq
/4trMxK6mpqId+h37VDE/ea9UkrnVZO+Afu9k+KtvzkzEgvZEMVonClgI+vm6PJtbX/Pb1teroOc
r8DR8az+Fitoo91QxKdqLAfWHZncjOpdCiVuhvdaD0//8X65SoaPskYym3tAZbNrCCgh9oFu44Kr
N6teRnP/AFdqZa60kfaRZs5vfSPXdiHyh4DhR7Jqtv37UK792btQRDmRWp4rsXVF1SerD/abVBqU
ZuxVlteBS397mqx7hB3z+4mFGriyEjmU6NgrkZ28dFlGppTvpHL7UiltjE1RD/ahAHlSICmaMTV8
ni1bT6EHTDHOE+YO1syipXoT5mRScr1RaAuYARkPruoUjeCb4CYx+17/aYqPI0g7fAMJiccrY9HA
T9nueR1GKeWPnfKvkHuhRzoSx+hPmXivbo3EcfoCWEiFUPvmafO5SM8mLjpRGl23ETfutjhYFIPh
kQahUR3BCnvJXdIBD+0SXW684pyLhhvyhnANDWYyBL2UkY24Oc0BzVVPAr7G7+MX6KEFIWE6imDL
tA0Ns8VOfaB3xy9e5oyd4HxpUI2h3HzIfUsyUXi21NLHSykeTDTjqditPD/8P4OiWylPBzaCH4dh
OZeek/ETeRkWqJJ0424HznOB2LOtXCb73M8db8zPfIIokifAel6K4uOFef2cnfUxvxtcbEW99Fna
5f/v57IAZeZgltRuSJvJlpU3qXpiTU5q6wlynis3ysBHkADjb9EgW+8sr2YVi/2wFjToxPzGXYWX
qbXdwlWBrPHMekTO0V4DwbwmGm+2n960jkD+h9HUIM9mdikitWnBe/VdAgnt0+uSpUlufRwoFiCy
TJcSKLnGXJi9EPGo1TK65TbwO3DccrghevsqWM51RIR7Df7uSKjfMEBQeNerZ8My3Bx9CS9TcZEF
o2ARbcQQ3l4o5TAVfLig2mX1YwSPEfUpNTjUvZldGhJ3MBnNVmQy1iU7649cDtwm/G6Wli5WDLN+
PhvPhaXibt5dqSo5OMa5H2b4qzNwv9hVux5vmHdAJD1HO7BcnF85t0O/16zeOcA+ulbV4I9Lzak/
c2vT7Dyz5FSw0TGprcOgEU0FvHmnwyFeDk0Ri0kbA3zvn8rwktM3xuRTEyo586XH9jEoZr4J0Wxp
FvVCAxth/RB5B9dNLS9gbTNx34dUb1rhUkZi+QBshGBu24VZHDhrIwtdsX20Ih7UBRQ50l3Cxmo8
FB4Mr6WpJJKpg5OkYowksBObusCXbye+Ek9YwZiXXCcBwGH/Nb3Y+lUlPS+kfHtwHsmjQ/GtA3bE
6d9BNkUNl5kq3sWx9C5uA9MSmDBLwTTVZBOdJNlu+3bUl2h2ussvaeliut6uZ2PEbG+DgFIi7+5o
6KFSe597kMKzW9oQi9zBKJ0rutV87+Txm7HrRln1GyX4oTNEGf4rE7e+UTCUuZCVuDXNVmmzeYje
GYw7PbemjMZ20b555rpKCJE/EO461Ro8NVdZK0K6Yxe/aau1Otx98RvMDyVdvDJGrJU2/97w3K2L
y8PiQCQcnuXT74mAZdvvYXIG9VPSNCerfC59EiqcHQI1xeNU1givO/ME3TeYkwixZhXulotXZDu+
RoozUi8Bd2qaalSKL9Zi8URAb2AG/gH6kMeltxM3m0+laEdKl9oRUObvwRaJlqA83UlxgOHPjtrf
UYziE3lqVOxDrTSPrJOxdqLkKCgVNBVFNk6TIQVaJFsZRAV6WWbz+bRZmEWX0rOsCpT0Tn6VZKvm
6c+/f9tv+wxEK8bP5LiUt934jjkRZ50AMOcRTdPfMH8Of1utD6/OAToOGxySp6OYg9V5AVaTODt+
6NlQQOpCpALxG6JybSJEmEMmBFYXvXHMriJ1SK7fAKeWggRDYfJCklhXlFkRtgq7lJnm3Kz3YUQS
53jnxQHIB6pE9FqIiGrOu2l4mPmY9QdxicNVBRvUqCEGlbVAVJzitCJEejQ5fmOzrzCts5E+hyBn
fQV5NsFRlIvuj0zu7d9osok3/xojkt6SO0AZFQVyQ8fmEokvWWiqPRrlFcamAThYVxRo9bCThytt
DCrTDXAAU84BsZGS2LAamXUXfNiEhNXHbwmWtG0soJFJPcsbI0EYBHGkB70GHFjAix/7XYEwcqNa
vJ5/DzCdVw3iJgQHTYVmWDAIay8buDhXGXjHClReh6L2CUZ8jS56Zkm1p5QVmVLmgQjBCRfwNbK+
o5gOjhiVW6iTIMmH74L+1e+u1dLPm87sMJD/dZeXFtVbArZ4FGYNzApNi8jK5AvuUokmQjwrPIxd
9eDpj+tQ248zr30iYeP7SDOBwgALEiyR9nwp59ltrh/LjIPR3gmztSSiJF+De+lKmMPpwdGCOnL8
6J5l8NY9MA68dSbQMyFSooHo/t89hhOPDslPoQgDqDP/xt3nCyiwIJHqUf+CBHQB95lA04d4/Aqb
lX6KyNnepa02erddwjQTI4pc3l7PkWUg23CtY6c3+thxUJZIMqEqsbNEMzKE8KuQR+yOn5Ahm/E5
3w4OmukhcvoInyqggPw9a2N5DylCV/wAGMeLV7nNJgOGXL2KCY+qgk4VGoA6vhiCNbs0Y+QU7sgS
CmLU6lfXTMJGkalccVr6aHFovLbWZjlEYvcyLoSo+JVzYaeCun1VUEV4uhJ3W+geonXAxZRiGuZc
Cx5z7gx+iOAadAPLdUTlT6SKg5v17bLtPav49PD9qlvmI9ODzwfnDRipcHCbTEJYT+KLOFUpKc1M
V4ZjWhCNJwwy7NLfvmAzoC/2KwM39HIx4k0OfOPEsrQscrgY3fgbu/3m1UO8yP5IV6d61498YudH
RWWzVrrCghwptu8WU+Fb7sf4p+YMdpYdvCIIqM/tspHt1AFV/EHD4ZwP73fMhexXDWD3Qfwzq8W4
3zrDkLU/VhPlBjOv2sxPbdDvSD8ksYYniSU0NRV3VWiK8JkGvEPm2rzHN0+KuieDpamJ4ULttPkl
6jNlXndkTz+G2tZIHgYFYrdVFZVcvQztyH1qV6WtBiscIAdMXd8MncZzQN7mLx7b2NgW/+nrhjey
Gfo/Gei5KCoeX1aIfj7VzF3hMZONFF5Mo9GQRZleZSBsSOtt5zb+daocdidRZaGMntTHw9WNnDZ5
8OAM9vzMAQCXAXDjuNpdcj0cir+jMrYJD8JX4uN/HfyrVJcEAkJFWn4YOCKMDo4mJNgG4YnhZYQH
7qNJcNYt6cRtRBdMJdcDDfBTsFWdeoYIMBSMVkEZLMCDQ6EIK0f2dZTijpQCWePzUnhQGclEVz0S
zJbCLmNLLGX6ow5htfDcGiE68ONuJK+TRuh1mc0jvyl8KWrqvDwa7jPaqywjKJjR7LGb2+08Bb3d
TI4rMHdU14/AD667Iz7pZl822oFOGumprbQrwQ9Fzi9fkW27ZE51zW/VM8veJMkFnBOmnErOiM3K
EQ9S/lFIwOw4qUmKCGAoZofo+izy3eeeJI4VvixVeWsru47IaeVUJVqR3PHkTNUVOQj4VY4Neu0K
CtKD+zVCx6h97pL7yqNH+a4hGygtGGB9/WKel4bUjaCZHZnpqRVxn5FbasZyWCQt8t574ApYKScc
tm5n78ARY1Pdnvf5KmlK5v8XH9gGKsgCRxnYqKKmzsi6lPsp0qcJLyYZUIMlKZngBsHDSo7Q8W6W
Ietc9CWKc+UYwhj4z6F+Yt1Z115GkAAV70oosrcAxMVUlbhLA7B1rs0c0W/uRdkEFV8KNAZnkFgp
7E5yNpkq7enHvQGB1zOk5ZWuDBnaSgEgXUhRTGLu21OFp80wOjOdpGob6nuHtzymwaTLPd2/lD7m
Ft+yDdxZ76x9Osw0XdQZq7iDzKKpezfqXp9dA1tyAtGoOFYDL2mM8BGMGwykil5TLvAURIJT0qYU
RBjY7/nLX5OHYdTGQS3iUMl4maJDLkMyfabfhIMEYs3Oaj1Pln7k6Sz+6HmIlC3fnYgCDff0kbt4
nVO1cKBTKzdobE+OWpixIU93qQE0vcDKynSLtDMCarVsjr1E8BxEoLhKBEbnlnvuNeAVO1Kpkzoq
9ImpTcAQxqjZolAko/83Ki7ZnlmpB6qFvpvTuonXulKW8NutpUJfA4kF1OtqNQ7EqD6BVg5pReOy
tZZfLjbv21XYKV6mfhSV4hXjqRnCKHyU37SB/TFppcVMoZBB3nU6XovZxHCZdgMHrkkmKq0P8jUU
ViQPg/2z3Ne1Fj4vTUD+19Uk/gF8ydiVZKczzUln2MF29KTtXBlD3aw8EuAg1A1XyQbgQ2e4HmFj
vqU/oz1Y0NEQ4LnOp9sGv4eBR21zpDhp9+GTEaqlj9izOZe7ndIv7ovyn3B0RDTcz351FORT9OJK
FrjhQMYKQkz7k5BaoZuS0PYGvpNe2Y8eFoSf/x5mlHkmY3Skgyz3capkAjwqSMtd8V6z026PC23/
yFo8S98SQvUkCgOKtli+jucbqCzOtQasQIO8jnggztxrbIMdrR56dojzZ/d+HI0YznUmC9S9/5NM
iaLjBLKIcWkdvEuqx5tIYLXbUSXUJSxsm8iYWLpBjFyFFQPiggDgKgOefsNookb5VXhlaFLWZTxH
EsSEoo/jTartfYNuQ8g9DJHkTFyDV9kHaa+SGKOI+1KfFCfXnFoYpW/C1TILX5uu3BdMAxmD2O0/
dooCVa1znq141TtlRZY0iaedjBBsZw63qsiCh34ETku6Dow8hs4aZL4SBrHqQnr3DTZ2AaqNYmlI
EVsa/dqyShfT2K3cJzicIVMC6Qkm4yy58zBeWsDJDkwumv33fs5J6ukrP4+wyi8Mbf+sLQ8As6oJ
04tXTuhQAP9PU8ePWkpor1OG2KJQ/d5sHjhFH1sW4O++8O2JZNvSsVZu5nklUlaMWOKZdsx2bMrz
76GH07lWnCz8gNPPTGBxcrbKVJkWM2qHDJKhwi8mfPlZavAwsur9FGOq7L+T0k+ZGCc+CTBbSr0L
fDwiK3bZxExmyZ7cpC8pN5zNQoWSeWaKIRXg5rt1/yG7XGTkdW8cDassoqEH/yO9RH+hjWc8Vv7a
NghRAxE8MJEKBaKhVKF6AXjadBUnsjXKW/1R1Xc+sBya4/BA6a8flHkKwHud0F42Z/94vKeE2s2y
I1184BVp8Xh1WIEdAvrjitZ6Wmh03mD+q9vEPjnp1ybjC/TcF47UKILb5kSEEAhXsG0Oyx2rARZJ
f0tEWVuzLVuwX3f5hcW3fdglnsUXKMMY5mn7PjpvdBltATkqp70z2rrMjx3Ae2hE3sys3WwMs1Uh
D2K1YgRiwbaodIaG6unGXV5fz4eKMlhyUPAGK+tqbyFXbIwJu7fpXI0QK+0/hAjTIC6Y5fq1AQvU
DX6ft9uC9WRUUzB7CP3hsB58AIRsW8fmnALgB0hnnAY1ce5+dUhAGe8jdmgY1C9kcPk2cC3kYlG8
MdRez4R0cIDNt9ICqiKGBkJAF9fOqUdcEjNtYVbyrvSyKIFwbChkhO28vX6x5xtQN/G1DFfyR1Ga
2dE58qcWIpIJxw5RdhmBTs5QR/8zETOl8NGZ8NFwOKbBrcnBlwyDFBZjxRdRJ5K3I5Fu+VBLegvE
nhHZQgxf2O+WIK0ya1qZ6F9rMfnwVC0wHtZ9yWfLKBBki4ICDWc1fkRXlVTiWRlMq3/lcCMrIbvb
gVP82BAiRCJsUdVnQSBUIdQwUFCXBeM7PzBo7BcfNaDmUwcndzs20QBOMaqdkCYT6Ww2HIfnBz41
rSmisJzgNvpLWZsZ30BxEwzb8BmdyXV25nwveuTUGHkg5G/zsUbtcavzVobfIekeFibJhXMSsn+a
9hGcilkqg/oPBI3L/n4szRvO4TK6JU+Q+MDMXcJW+pdWPZ7EAvtlrBZfFPItr2eOuMCPRvw+9r0a
RF3+41tNQ024fYpfQbOlKbVCGwC25HHMBCZ5cTioczsHe3ACQSQqenLhekuCMys/pEbpr5kqj8RT
tS84URAQxDmk/Qk2mI3E5JvrizjtZrAwXHeCsA2b7pOQitFMlRK3GOb9jvsju2/5peRV4Ph0xw+g
ITRyH9kAHERbAMIwlv7BZ1Shbe7AZYxDAtnzYM2tiT5JfTmFXtJXR4w8qvp6oeAmSe+AK9M1IKO4
GL2OznlBMyJqED7VjpJJkG7LSLvEP0MD2d5GmWa6kiB0ItIs8PCMYHf5bDBdDpEdFVuF3TW8K7jw
axKmfhUp67cL3/p/QxApEtUIL73S9hRN/Yb2kJBKyTOMB9Tv3lTKFbwD7PXbb8ZKBbBW0zsO2lid
a7Pei8zkMUxDfVQrIHNxHf3beShdyzi27VF7HjbL9C4F6Su+9ziuT74ns3Q3ZXlIykWov5P+rZvn
jfNRzYWD0JOFGB1IilIKQJfx9OVchrejvEN7OV8nVit6MKG+UEdy++KB93HNFrfRYLmAm7wXyFLe
AWyWsYdKdqwWh7OQw2fJeR06bGGxwKjBKs2ePmHI3diqNViXK3l2rd5oBOVvOU0HXXhiPoVPLJR9
14QMHIIDpZwcKWV72JjFA2S2CvauUIftm4b7akynutk5+KW1V/o+g1u6Ff5gUlFa9+FfcAWKvfmK
S8UG8BfnKKlr6XEvlczxZM+B2KMNbd0t+2NBNNYyUMwiDGTpOioolaTP9KFLxgRY8J1Ukq9x2u9k
28dZBBJVa1Qx1m2FNax2n/PTYz3u2rGJfxVk0zpdl7Dz2vevo+8N4vr/1qALMiaD8/FT1NQPgNvK
iMwER1Rnnw1jGNztHhgtBxUsOJTyAV7rlENg/2qNgox1pAMZJUjl7xCQjtInZ+9cuXYHB7VeAd94
VCaXwOrt/Hz/MXOODN2sjS9nw27STunS2uUq/0EOC5tPsqVc/K4o5FvA0KtTx/fnD+9jYiXbUPxi
xzHqw8XnbNLc7zJcEKYY+aZgCWDq3bH65PAz2BfVj/q6/3zv8Cw/bSsVpERfzDCxHMTMvA5ihXiU
zXlKwaGR5g34dydZF3Bdp4/fVhFe68t/1t6NPEchogiTi0qhvDwHLZBn4/JtVOa/GKeXbGYsJpmH
aggfi09bdB2z/qm6Vh3Jp9wH2wk7kKvwYpT4XB3NOMcnmeIt4e5ZgYqt1bDMXqqA1tDkKZDKxEUG
55GJGcMHsDL31C9tpXmbdfYUR7AS+89MdP4oul7fKIoL8f+Dqc0hR317V7/4QdtdGIhQGrGldbfl
ATdm8/mHZWBvlGfxkGzOky+o4aDMzDv+MHoiGRIp5vQRw/0j4JZMOjdpCqvau2ajN90iTatpQ8g0
b6juoMUEcEUejqc2+ilWyUW4S0AHOkWu8sITV7tBWYHPrauwYPG4nEJVs8Rm/ib733jvzTIgH/Vc
QqLOvrbuJywd/vT3ZEkOBrSbnYvXrg0qcz7HkFxPB7CF4sSx0sN7yk0x7aJOU7iPApXKG87mxnzx
zwNJKCwaxWQ8pttdQXr7hzMJTjCy5lk8+uS267bZM5SVy4vi2SDT+D1tHq9Q9jfDXlPa8mTjlnIN
ywH+7qr1FB4JOKwUkYh70TuyqaedLAAnX2+TZhkOKO8QCQP1THPhW8V3j7RHvozK7I+NzqkekCw+
91jFt42zSdmCiky8LXVRjFXYaTxj++4nIQ45WFadyh3tzvwakMgKBdQynaEpKizczxsQ1VzoIy2q
Pt34fHa4qvZUycrBLApYrZkZGH/xm+CLF+rIwn0T7WFJVv8Tb0KE5PDIfuRh+k2n8elo5lQD5Hot
JtV/RY1k9L7szmq0/OUjFIqqizL5qc7ZaVaiYXV9YTZ+dM3B9s4AKsUT15+xkcSH7jKGiujPjDtn
pDNF+KUrI7k8vHXNjc/MLLvbD5HrgP0Wd6z/PmIqsNgjbLuW2WZ0GW6NTxluTahHqFutA+859UBV
EZ6exPNr8NoyZ6HOXYyo38dKNb8MyWebzIQBcg44RYuEFOUSsFqcC2onSazET243LfJG6/io8C9k
iUNQJhX9WanXNlN1nQ4Zij6MWwUgvMPkOn8Q170hvKpheCjwYvJfAAodmiLH8tFNHg03n/jn7ajV
WJuUcC+wmx/fML+tIszHZ9W7rPfLh2fUghArxI1r/cW4wWDRI+XqZqS0HqNY8C4/04c+xNK2HAqF
eeLq1UQR5M07duieVD6fBMP/0SHaJXxlFBcIf6KbFQsgyHxGYXBJKURy4LpjzUZF91BPsjNcW7RW
wWhoEhj4PJEddZ9nPIxNNbXRfrEMMZ3gYZIJcW79ZBKnJz17OdtAvnzXaoobxsu29SJtHHX+IvGI
f7zM6w3xT0SUI6svihY6cjXM3i9cL9uW5aT36oeRoaC4bBCZG9kavSSltKHsxtHEs8hGLtpAtUus
z2WDfe9TFmmD7sCFgWcunrpEHoTTvKaGozZMXhx4JYhHmTWGPPYtcJFUdz/An+29YsZbsG6nGnhx
64jmzu8FlDtIb/hPDWp2ciKylvCp2bnlWoLjmFkP1qnrdchEREHkqEfsgukZRAihWg1MjABx5ooe
HzyRe8HhONzNpmQoRdJs3ivp+4abaFxY8cx6OzBaW7zsWHCGaeL8BarKDgwyiaHm1mzgJOdunPjl
XFtwhv++lB3/3pyZIAikflLX7cKfaim+Aijz/kdLKf6UMwJrhZK+X0yLPgUx2emzLYLx8xkXq4gK
aJGEJz5YdSrhpyoVmqr1fQhii2H7OA31drAmfI0qgxhRockfNHiDN0XFWUuXA9xlsEb+5HXFByOX
TuRMYqzO+DYDGC5pQVIcFfDH8DrN5CUfajuYJYwUiNP9EbkD5foFU6/yaVv/yBB/xujGdytO/ufc
RKZImMEbrDv6N7vCL6Ud9hu9X61fzqRRGF1SLQQbr1/DnkNY4ygYOyMvr3hPy77e4FLoVkirudyF
LlJcfY4rYe1OT8qUX2vxCCI/EHAcf6L1QL1OzNXL/vfNZpZQSs9uFpAViB64nxf+NACgaaoKVzDw
cDBrakOSnsth5H2tMrXqsXXevbcoLq7GXMX+YS6YiFZS2yxU9MQjlDXIt8xni0c0h7eIcAN5yLb1
G+W3o1EEtXlS4Vj+rYotOqJGx3FpG1La0osKY4MdnSqwxagE9SS6r0RAw4qLzRUEP8bSKQOrBejW
FLq64aFeyluacaXtiWSnWTlyCJomFmWtqfmafxGeavIPWQQGkoJfNCofU5WPRcFy5XpRO7v/YgCb
g4Ar5FmUZ1dAU/3xpwCu5Mza5ybwldCWXo7g1XMY4umW86C2r0gX+7NUo/xYUidEvBr/LfMdBGad
sxk42EzQXcwXn+GzY8tvEvX4sB9UbJnocPTYqbuVW1TkpBZs4cuiW11+w+HiEt5p/YRqw/OKYdte
fZoMnVrwkH93ukvB2/Hlown25i+hnrk9lSUWrfUwqkGNyNaGXMLA0La3yMvplLtkG/nlFO7cezB9
jFe86emQhUVhWUTio2qHGw6MyjqGrO5eyjS+YucUhsDzoEtappKMhR5YFB6cN+muX6RWJOYlimeW
ou3MeTQyY5w/DlooMYqIE/RLaAvtOWWHXh4HMgUhLICrQxXckgY1FWpWDa0cG2xsZFjdEAdtA491
Cz/VzyXPnsw0y2nUTzutZHXdysk81+fIaZY08X/6DaG6cXvu37mwmfX/qcRQv2qaeuL/54k1yA3P
EJrfIwFaYkZzynwEVzSm52gpRANsnoANPJ+kvCN6+R0RD+veLNhCh3Rn1izmkq9JPXY+qKzHP+CS
sw7xJ8giIhvdYNkjqU5CKLeqF5jaDoXbFRdyT1itbsasb1nvX6GZAHKJRgfbDilZVO5IrM7UGGdY
bLs0EqLzuU4W71wllCG6+AaWYIhMvikBqjyusSpbYdPDu2d1qXwxUsS7yxMSyRdoH15ZxeF/jXe/
C72tfAJm0t4bsoPpWEctPN3FAbUgzcnuQ7e4KFT2843Pt8mbanN/lkFXbSS7g0+T0Z3YLovCcdGO
+q845b38AuMs1Sw4wRqO60xHXcG4iO7pb3jh9fdjdaZ5620GG1gCDPvPwf9T67q1G3dJZGSwUzgs
/9RwYl/rBB7CWwaP8olO/8Rl4u6IU2MaLZv9/sdHuAX8Ny/1OLoWbfRrzQBJKcM4kwxZTau9fbP0
myA+0KaDM3PdjY0xNvZFicIQ3bd8BIniJGJ9+ntUp4rOTf85Rp1HMYtvOZ6mF1hhy5496MTdjgS8
G1RTTofLM2XXsD1QlzJI6cnRIvP3fHNABBd5QGLhOVj1/gEuump+Uf3DI8QBv1Z4qMZdD4kthKHm
h86QzUBV9L3cqTZBH+4mCNg9bWF9d3D4iogezbJUTdcW3juxlZCsk6vf7aa1M0YPMl60gOs5boPL
Uy77rr3EpG8hsvrh6awAnTfqvCqGTVGHxsTAdRlO5QzxDtaSHKJoYGR5xQlsDocbkhOJhkFOReU4
Y63g9iLfiuY0FLfBNYZLGseBh0pa8Z2sODW90yGD96QiHL/CzfjKKMxOkueNKztvrlkY2a+2sRHS
CgV3dL1z3G5KeMW9QjeUyDSswp1M1gAYnlADvLfsoMkHYzJl2VKvfGSXD2uumi73QXvXzG2dmDXi
v0xWqcClkyHPCcwySY0xl+K5mwDwWNpqPuOhlusuS/BC72thzC7lvPCr1i8/oozBTmGFdo5zKiBH
vxGjZlssx8G+h5u4b0A4+9VPMDygJ3qy+r+MoRASNQ5eYwQr0QMqrFw4+1xLYs8TX3bn3cFAFjaJ
N8WpLJn1uiFBL+Qt4VYEG3mH17RwkVl9/+sL82OrfpRe8AJnDMT1Nk7SaDxXVgV8SmjV2DnC6ndk
3QoOA2AkcQBNbf+hXVYjXpSW3u0cYTJamQnHtSbzNjruQrm8HJNqT/MNRiDTTsN47US2Bg3yvOK1
eCrrS4EK/RtrNp+ItGmEyf55m1t9P4Hn6ztCjl/kVKUV8LWG2zervD53/i6FUDtJO7abjmYSwJrq
zC+SVUzAxH8GJMOshYKEZ8hM6SmnP/faJvJqhsZXK0G+XKYmBOM1Yl4iIXEfRc+U2vsF+NDaq2Fu
bBD9g1mKN0k8cVq+9SaVvQ3EvUGIGTjYJSOpzWOhuu7A5kdSvEyfJ5/QGmJP3D247C8pHV2WoaPA
D9sQJAg6To6rAyxBvOiAKmdA9Rczo0hFQyVnJYUjogPQ8j3JMJFyal4/9QKEUa2M19sz6e+VLt7b
t57jWn+WibT+rCwfiiKP99c8knuySuJ9c+wcXQMlpP6wxoe+dSRlVb0LOZznYpeenjMo0ETKce29
oI0zKYW7wf/fC6SAdNvIQbIl9vZvGAOwG8X6GTGpn/HqBrYiil4Ra8qNGRGgVhfiJgKcW0KcgLlo
dPXejW68h5ZNd/BihVzXRjqWzTcVUg7bXB+2swhLqlx5Lg/UtLBiCmh/wHNM6yvXmb3Il/lF4t/D
9/giGYy0c2rNL9vXCrU+zvBxwsJ4A8dC80BVBZRbjrACsel6XlkktQ2aP7mBvPWq+BrwJQnvVEcf
EIR87Ae+0GKVyZoLnGaFh8m3mDUCxM/lxekTmbarDmxsmnMAgVrm0fXn0zrywTXWuQgCtTMiZ5Qf
zwNNxJS+jLLsPhEKI2jN4Vca+rRgvXbBl7LaaQnD2ggg7hN9kREMJO6C08ylS5HP9lAAqc+SfQa5
1qnG7+PkkQHyh8j1dDDxnjNDl8UYu7OdJWwEQ5Vl5StS1DtPPlHzzerOll3rxByumQUc0r2GZ1Yq
/Oa8cZVhN5hjXkf66prG8bSPRtxT4xRilKusdqbNbKoRN9mvdwIfQ/0tbfblaU0pJeddIpUqHcRa
nEG+8YX6dKUj+zQrEzC9G9ZKXFHsxXGWaMd5L8fR9lN6jYmUnINv8z7LtaC5WK3v2Xs2GdZHhJ2f
unKBkO1pAFM3LmmrqW1EqAPE42Sfy9/NAvfuQ7gqht/NkYTHatnHH4Gp3kVoptL3U4GaDeo9OFmE
hXDs8Tu1LeWw9yFbvowtJ1LXwWMNAcAuUEwXJ+4KF1KBb2jovlRaQUKI0fViKsv97Vk3WeJD5eYR
zvOvujdSqACzU0PXTXkepETolhu90x22i+Z33Xn5jMmn4iz01BdGkwZtpWcqTnn72qAIzeK28LNC
LOJEgboZNvpFxjXOXwPNwjSHCQ1OGC3cXLVj+J+/vqrkiw2o+PNGbRnc4gvCC5MxWMUBQEiW6P1o
WXj82pL/lkZX6KBqVr+ZQ7HUz/TFocYCokSrCecNcaT9kzIUMJrcjwLUrAkThtKyfu1GQfzvUQHH
Mvhn2HctFmAQp+VfH+h+1k2CQV2yhdTi4DNQK/ec8b2d8BDz2R9mZn5s6fxLzfLSCnKI76yERGfJ
MokeLsKQQH1axA3bCYBsGz1qt4sLcsvznntvGfC5mH9cNA82mRM27lk3Akb8RVm82JQuUjhtdI2j
VUWVxXVsFq8nOrCoUR7ImBSZSzyO2dboi49SurWee3zM9S9GylMYUZZcv9HiUa5Zg47J1qIkpiAA
aszZWHu2PXMcnHmmhTDVz84hAafBUPGcwV21YmjXF8ElI9IPXGQgta87zvzv2+QZY3jxNEMQozFY
wD9SZys+5wq4/09h8aMr62PpGDhgWfRP/Ya0LfYjkSqSYEhSDqct939Q36sS4ir10ZXMfpUqhhMm
9Zm2DgQ8/sF59QY3unGKj2nwmpWLQAACrBEUMpEVQdBVrej9rP0CpeHJQIzgiwxkG1nqGRxWRm6y
SvUCQ+ijAhsO8KXHLrYcWcWOWLYxR89ix+Vec1P94TwTGk3V2VfzOCZvrLY+Ry0Mk5kQ0MlVC4zX
8kWW0PpTVuImQC7bpxVO3vHyjJgVVhaIZQLaU7RR9+ZTX+KqKeuZO+6ekGwOodJWy35ISgUUQLzU
UkJnPr5np2a9LTQwW/VUvP47NrXdHulKfev7XLEQDzAAvHns67OkJUCNF+B802H/l/2NCXEeu+3v
/YsHFFvl6YoA3EfmAjEmflyHELbhwZsWpLz74qlJynDt2DvrNYEvkUGO6lFogaiik8QaR/xhPytJ
ykf8oxxjzr0wTqGeE6TyCvuoV23UhLI4XPH2OrilJiCkh6pgloAUa1vHQK63AqDgi7LQcGXklLUt
ZlduhL4zsBtl4ll1Ramg8kLwR9NP6rRzdIk0SAOzvpuNPJBa862mMUq75LuXhkYsJ5Qx5ZK7nkW9
vgCyPFJOv27leEJobWa5EDMkri+K8xLnmJ/r+feLECKrnXYlPDyPtSpkmoy+hrToM0eCjJhp+mQn
+fdg2+i5TWD190oqSfa0f59K5p8patnE5DDoQJZmWBQiv60ZK+3/gE1IC87ji3T3E+EZ2j/G+DjM
Hvq38Wvr1AO1Hf1hVVvbm2NmSKn3R15EzRpCvH9rgx1yRDa9BB82Nc3kKT5uIfNA8qJrRP2aHMxl
ZX+Op5rxLFjrWrvVURQQLe2Si7ZxCIlM2KCdr+dSGFo0gOKzotn3RPGc9pnN+qVwstbm0mhgY/am
9y/HGYnc0wuI3frmoXTeqHqTm0Ur0ublPGYZ5yusaS+eEbBO+lpQtoHfjK9pP2VikGf/uj7pL4vh
flQ7wPJ0lAcZH1W+l6fVj0377vJvSW9gTdY2gID9Yt9+AOkFLJZZZr6z9hvTO6+DMCsUDbmL0aVk
b5XIo45AyDpboXiJKNQxg8Au54QQ2SMXkBKzi0gNEHz1sKy9OJO9LCy1u1fg0DFWKPRipklXCvou
cqsZuWWCnIbacFvjN39eTbt7xKTj1IMsRByaJmHGLVlnpWrHS8rSn2ri450lHKwyBOIAI33VqO/I
3R4k75He3SRb6TDZCHzhDr43hW1cweVXftBBbQgFa8DJJi6cjUG8UqXMxLDmziXEc4ABgGnF0fqV
FMZ8rppw2p8fzTmD3vkK9ZsTf2KdBEgRcE8lpC7HduqfMuPvcO/O0lMZEPPM+eietCOPclh7NIK3
nUAfLiyRsTxn0vQW/9lcNLmQQBfAPcbkR2P9pDrYno8mpLx4dfuZU0rVMg0Fes8W5ABFO9nZvlC/
PRikNM/yjsEsoHVHOsMusT0rbcNvVr+UCGRY5GswI4Yxdh4T878IvlM7wdfv2f84SWN9gcpepRuE
ARCp1H0YVroh0WfyB6sZNmlmb8wU5NBbxHOQzPek2t2no1lzjHmaLKr6XZ5IRjdo7wEYxxbAfLXM
vT50BW/2P4InUys7mHgHgPntEsKQjKnzSWBL8IbO+OqlHvLsVGIBxhQI5TDy7MoARkF42Skrv0MQ
3MMOsRVVKdF2P36IEHqDnT4Zx994c6+OEpjoAUIQIfSSdSQsic97wJPVe1FLVM3v+f9cg8ONE7vt
HJ8MUNHOVJebmIZzXsrYzdwZpLFswFzK7n19glHzTid4K8LaVO0FRB7LSo140hoNSMuAzhewCL/T
NMCCnvfMXaeX7FAgHTY1zqInm5NsoY15Umi/fy3jL3qzVlij5WtB3wto2a6FwH0UBfnaPtDnaE75
o9m/jFWV63lVnxCChe7cEaaFTf6RFIiAOUxwBK0jnmEryHimn2JNr4ge3gPfHDWvkqD8iml94rNZ
Xvbxqs1VCwlhR2s0tpuxYGgmXbQGz4qxxIWju/PW2sH3cNpDEFVb3zPFvKu22g/bCxjBf862J5/s
hyQG4g2F4RJ0LYBSo5ioMGJqyaw49keN5HNMUvTjzD6NYB8o0NcEkdwcCRf1tTEy7tCAPCGMc1n9
KgKjZbbYnsYsxuq+PmtH4B0oAuRC2VvM6zNAsuR4zbrwsV5GN13FXNAwCLXQkvJE0QahKeop1sB9
F8NuufS1CK00XwqZzFWLVr5kxRsX8fGTLgMoGwWiEVyu5t3FS5FW8HaAXNfmL8VHM0T3wMetNlub
JLKqn9YQ7khfMvf6oTV76VgBAnYHCBcyxmaUBeDmnixG+hz4hovKNluySZ9mJTJTk736Gg+42y1K
YZ0ZJg6XHnbHVqp+eLtarPHBXlmhFqFAHUpPo+YsFXS6rRCwMn4xPuNf5XsFy3O7B7L7s0bTIVDF
lrsHxB+aEDuV8zNyNvyrSaYqnVxBcKIE9eZRmzAJJxjDNWpFU3W13Zx/JmkOz+CFsEBajKHAVi3f
7h1WDmxn+0VJIhiNOIwtmr9Xw45bjd7R93IrL17kWaWsPB5OZl8qamUlJhAnV2AHD28y+jGyhNOu
sgfWU2TqZrpS+COi0FtvqUrjbRt0UrIpGI2H3zKDkceFGX/D5fSm1usDq91xrrE4eirGZAfI0G4s
0z2AMI4VbQgk34yBGnwXAAd/iKXjbFdVMbSD9nN93cPjmNqG8nhG1HEP9lReJhlbGLt9ggGAyZJx
3s9/o8hzsM/UgHy3nfKd0Zmz/BBQcH8hOve6UmV4uCD97e49P2chRSZipe9jefkGnq3nbM2nCqnO
wXMDGCrZy1bZRRYewtDW6bEcYhTffKdwyY7nfqqxYw+7JV49Jt+6hElzFjxVhNsYmRM3BW2FT2SP
rW3Y3BOHKKjlUgB1WVVAS/VeOQUfD6YaIrH67hc5FwaKnV0WP2CO+4H7wE5qb3i1qXu3ApZ6I6an
4F0rxGok58FKYSF9E7oSZ6h6dJiLKbzgQ8ZZzkqTJPve0+GlkYd94lYwnoWV34i4M6ronFrNLJ/A
2zDalBCAMpJ16rU+03d4IU3NQ1JUBxvVJV1vhSR+ibd/+bYshkxEI/CMVAiYBzQUlpKhy7y8RbBh
kI5RvBqoXU3Hn5ukaP9W/+3Br/gxAE8dhcGrE45Qr+ZtXC01kq4bjaKBBwRtilyUu4MXVJmfJhzj
G6tq/psDe1cw4U5/uVC8lME2gSAEil6HBGwCHvMY9uPpE7BNREbKXVlRaMMagxMe9HKwbGy+RJJJ
qQ1IPWB6vjzUdFLjldlwTtIrxJNrQ7lcmmQ9xv3euyFrtY/pdZyn3FyOcd7js6S4QCAu0HBLOjmD
s+xgP3dspwSsiEQ/SWjT49YoEXNhuwjLbCI40HrRuI2A0b5y+vJEzJHez8CcskqJXYJimBxxt0/d
9wCZkTdGK1nLTpydI+PB8DktG5+RKNZYJXLhUrCMQo0F518b96vEepe+wduOjJWsUq189LtuouMg
Guajvvo+kTmXLoBGvu9KOcy7vIOflXyPCejkVSSqc1OwSxuthp3sgg4wXUuQsLSTpe8xaljBOTFO
8k+bxWOrf8U0acYIgCqhLudreMW2mttFvnw/sMj2BZdLGCTsjFm7+lHzatrQ5eGuxyrXLOfLp+aq
JmPsS5seRD6gsWX98mmvjx/7c+b4uRfGI1RvoWCdarMjfHJ/lyI9mQvQd+Jmjf5FoYK1LZ7VeDhV
O5bcLacn/B6W9zWJqbYRifleQHozHsIMp5oCxXhWF+jDCQ/dp2m0jEdOs85GxQpVjfuXY59eLXw/
OWwSen/vg9PbydFNuOSTwCIJ63mK6XpBe0YO3Ca7TV29LAEhlw+99tv7ZTZAjFivRi6OxN8eaRyR
wRxuZwvQl/IxGhigZljLxWPQRPEcCdiSrYIUMdvT5MVXdkRMtJiaEOYmDnw0Q+OSJ5BZKpo5WzT4
ff++fc9cXSpbhKqJNS7TUDrIEguHhuo6enRYMYXcRvHz9fvboWTxlyx84Q6y2tb7YaExVuUPnKN5
HcyyktPL41yMNJij3Wq/z40A1tgoulW2DchUddO1m3KBwk5c2Pyds9AG6pB6/jsXlfX3TWjw44JC
gX0OSJGeykBrJxhUeKayCmew12UDVvIJcUWkOH1KZTqrD3FPWA50A5cMgcdWMTkvCuw8mSG6Y2nV
ucnuur3Ly6fI8jkZdMKwrIlgRLqkv9YueC9fSYiqiSbIupDS9pEucmfuVdveSrG0FRw6wXRnRbiC
7I0siMZUzARLXNUE3U1ZA0QOYhqxkrAP1RwHX41m2c4aGwB/OHzjxVxoLUBWLDmF93LRJZa4W6ry
9nfsLagWLEPx+aLAHlRxhyD7pswddUq6OgXGW/VpIn+We+P8H2QcKselLX11QE/Rl30QtYNxV/k2
dCCcPsWYjP9B67dBU2u3b3UMf5nahGRu/4bZXKZqN5ReKZ54tZTJyCCN9AakuzZKelHrVbLhZpNT
L0Bl3PBYnlDh+sS1RDjo0nSbigQhGKfUHK5PFu0e5jTSFa27YNyA0pMuI0u3C/kyKOUYBjLY4Dmn
Bvff0MBH7rZWcd99eKnwJuvXIxDuZPJNZ1YyElyG65NCocurX3Gw4Ee4DKmOEgEPGjPYIEBBn9j7
YyQt4P0VG8NkzWpnJwgLy0HnQRKp8w2f243PD/+pdi36BiVX2STVfYZ5S9uVfdFCNeUjA+O/PuE2
dP+5s5XbEFBrozCXCoUJZkpn+Ifba9E9kl3xiYQAdq2vOBmHxrRKV7KfiwlalQmtaNxrUdW77HFx
oToAUb9pyRBopLgh3lnOYzhopUxt5WGpqKFQQeVTuo6YGBkh2hmEVeOytCC5IgnFUu99EcC2WGut
RBsae+MrkZQF9WAb6Z6BD/ERYz0+rGqjb3xkiBNidWm0F9EQg0Hd5q1OQgH+fvjKoLxo6MRmpb59
1boGkoM0xbixDtIw87phX4RboFUQJ7Fuw2zSCiFe9OenNSSI+0ITVZzkP506st8yXHASS3kHBMAD
dc+hScEFc4CQI0/aJ07KGbfxXkeFxNS5vVB34akCUxYTkneNgbUu+AueHRpOzGl+DsUqIUQMja2K
jzQz/zt4+G6wr5+CP8Jsij8ReV4VEzl1adUIMkgxRXNJGGbjw9QXiN8aMIDhrDfQFVuDaIzuFxut
suG+ndF82wKwBuSPI5rmjPgLetgvM1/j+xCPzlBe9oxtUpG0wfFs/hVpoISOUgGYQ3tjYNKHHk0u
4uYOmF5VcvK2+D+E0dOERKu9l9JhSbBY+Y0kjzAiGjhjO+78BWnZmW0r8KGvNP6MRJcGKkFKEvpx
/ZtxujQh/C9GodV7XgcFyVsfBJrU2DnVxubQDc144ttw2HL8u1+yeKiFqQQB6LU9PmnFJ3w+SUib
D0PQ8tiUZMQZ5y4zVU7CVzRMaF9LqFT6pPxFA0El43x5IYYEUyhh0B0bmE0BB+TSulf2LwphIEno
omCHagMnNYZxq2ITta0QDQpfsVVa6T1GoS/UHIG4AVA7VUxpyfGyAj5ETVQXN3LaGlmSGVymDa2h
3Qd4m6NtXeK1a7C3vElsfvJnPpy3UsyCFMxaDfiKawazu9pdhYUI9EKHWVDHDrX26utCkxbdTHyN
opC+tk0RFDhd/32DnnWASFEfnCxwQLXebsd6F+DhdKdXMTbnMBY42TPGcRkT8KoH7K7I531v2OKu
d000NCPIKun4UUFmS9sTKjTupCYVAtzdV/t8IP90Z1nQT//ma1JzOrPLOAF7DoVwsqBDdWJp/pMW
0KsVFmNpM9ZdAXUt0/UimK66OQrYS5zdq+U9cluJ8P9PLqvCzsWqalih8zK3QXnrN5cz3zWE5ElM
Svu2ON/QD2WQfwQrU9wW0CtgpdQn2B3Mjzm79rOK6vlFE1tseWZJQObcByX84+tct4fRvPMTZXG5
L5BAuDusIOplUC/UZZ0OnI3MKg161nGuQWO6CNGTH78wL/dqyltZjCrhoXnhbz9RG4We+RQgjcsI
7kxC2B/HQ+tm4DpqJIQCtgTI+Rwml3K16JttyKa5TNhZHJ8Rf3ri9l3setM6uYYrPpKZ0dJZKlAT
Nz9zh9AcETHPi0M6SiXPI3+gvsoYQgljI36S0QpljGYICL+uvXPfuiDIdMb04UemsQbzOKFAK/hR
2gWQw259A0ZwKsGcr2ew8aPGQVc6RAVnT/0oC+M1YQCpNBKRNnMFuJLGZOZRsquSFqHCGpuMxWTd
HdKwD9rlcTPr3bHcVETStpMHQGaY5MITDY31qlWXHH87iRSIHu/IQThzMB9NNde3Zi/3sRDq5F8V
1Jhx2f5Sce1aPRcjTmK2NsdDqQzldN6T4kIxZN7IcHbmMBuKUOlnfdPsqYz4YHa1/ndvVxiw6dsS
JU0N6934r3iLG1qrZG5m/XWJDzWC9bdr8Kjo1R5wwzy7GtnZV9R/0Zzqke6y73NWhbqx/tQxA0vF
FqRKTNSc3zHZHN+DEnWSWu5CakupJQPNl7baQ5l/sEU+h9N2lv3JRIjhU8aN+jN1/3GQtdo8v2TS
C2FyGRIn01XKpHbuLzJzvx+HDpZGftqlr6zgBbrqy07K+Xu8VuboAvBr/IUZmCc8O8KFKtdLUokZ
5PP5mOT7GM22oFa+5Zn8q/iQcnUCSZ3p3a4PiTW718eVleOHq4U4u2gC5/znUiITsh2bT9UQHK/s
MP4z3DDpzQB82G4iV+W07ovlGW9fuRl9OaUO2qJr1CRTwssWcO9ryNvhg1/pS/X0+T1nEUS4LZFj
Z7iViG/aaeWib6aneZBYOT7HfFwkt8UNKk9esMkB/HHHUB/yeMOAZ4H8ch/rDkYC1SBadSkEJ/yP
rbu9PZLYL9niZKxA/2pBJPSyzRx4je1vA0dY/0Q+ktkavf2XRyZwHYzJTy8yNlNj3/qh+oc7ClHt
RO+q6Vcq2WuYb8UbiCpr6KSTod3Nu7uk5Z0haX7hjoCsCd6TisMzqeTOh7d5TsIpTKTgX0kbbzKE
1nCoWra3NJXQKwk+9/XUefRSm/K+CV3IuTOHntrw3mao4wioe9i8Spsg7ll/P69E9nlEPcjMAdph
oGKrYcT0H0H/lzjLdyTgPmesfw30p36hW3s/cbLciNp0bBk5LF2jAlM801XJRbROu2Q99xhqt4jO
kQZs9SDxgRfEKXSQsl7U4TGudTjVA6Xl4hFKA8MFM6zUCX1dxax0SeRcQzYWZwU6cnvhU6EW+blt
ox1tWfmHzdFjhF0eA0j3oVgkfQsYnE4IuLE4ZxqLRnacOGsmwxBtLKEb3vMrpfDEfw14ilQzQC5G
OyeqjuREwpyT5T1RpM3hqrFBoyXuECjaV/X6CgPdv8AGGc2BKUgivhRBHmWeoaPh30gFXRTD3lsA
SkzNUTJq1L2oCGDglHDtGntT/2zwuyA4yVI3MD4KJxFqvPKlsKMHmV8p/KLSBnGq6D0Vev8x60IS
dIvjOH3VuVLY+lbKUbQcjOKDUq/whWiOmynioq+qJJbeuNLoo1TMjuxcrCid1cqwBq9hx3fbqHC+
ef23Cj/+Ot1FmZ8BO3B7yZEnfGo/lijHFdqYiUk5td58rvo3YHzFPA36s5Er6P84z2Q6Ih90mPy2
mANZ6kd05F7MJdN9zgPhUnQOeUVE+GYxim1mOEiFxdabmbNL8SKFVggUe4laAv89Ez4+yicxUeFE
aHjQ0DhiAcCC2uLe5w9Z1DOjMGy3vWlHxX2oSelFT3CERMix6qcjjrq10450+usv9XxzWem6tWAT
hSAxE8Bxc7FXfSSLNiWBpxmV3hZVh9WIlldPcNHeO/e5iaDffuz0FGKDMNTWzw7CCq7LRcRLjuen
Z8ne7fK1NvvMfY/oP8A8V16PMuT94HpvleCFoZZAsuSMV2BJ94iyOAem+ZwJXhxKMZ2laJ11EZwq
ezU8rR+LP3d4xnjFj0wxm3HwwSUmbzIym4v5TmcvIgkg7MvjtBQDqQF7tU316fGcZ9bTK9RKn+Nk
eqZsrnsFFfHSUgxZXYFEm77ovkx2SC9f2x/M2YQls09favTC+AVSGXR8E0fhjAMtCcPq0WUQlKpq
z+BZr8oyS1bkvs0k8QGwS0ulcVsR96UWEb/pscuEN4DguHdItEWjrlY7ibF9O21ZS0IBpUgV+9gN
eY9vszWgjhF/BEIwIAukyDmJiM2MrgZ31xHUwvOSaxdbS1n77OzbEe3u8/SnNlLKQmKMpjVvdyNI
wW67YKjhYeCbMSZ7Zw/uGUYji+kLUq+uvKL/PL4Y1CtFI45DKRiJZzHReEkWUc+7r6bFA+H1TX7l
bRj6oNuL4B7HobKT0yi9Se/lxt2K2GnKpuJaQIFdp9Ji/AyLx4L77LyyKk9Q3acxU0Cp74trur+/
R6qEzstIRbXMWvodbpaLqwN8lOj0xesEUFe1c0Nh5hjpA+JaLz/LQDn9EoP8EnYynRYMb3PT2VoD
QLxIf0btvcQV9gVv1TeLsxMfh2a+HrpvLXY/geXPA2GYSh4kfyw7BzwJypV98S52JQWNFPL3htBW
W7w1osJ/TubSPVWbT9AiUmcevbpya+Zqss4jRTvj2F8ruxty7FBx65SC67vwOUL+6Q9x2BvHN9KI
hMPK3jAzvM7tRkOWyn+Rz6qbMbOztW2YvIe03PHtzpJWOp/aUGmf89EVOZ70IvR1tddd4Eqf6dPe
pwY1B8uSo4THHkt7ACAUyunLBLkEXn/O7n5AJ2KcmYOANgT974ovhmJY3mlMZdXzTqjkKRg4ooiz
bdq9XP9tYzSDyY8hobkQArk9/i+DcITCYvkHKAa3g8umEKgQfsJIUkDzwy7Csh0vAzdk0JeWZGys
6BszdlL0HGyZtPayCS1auStbwXfyjF9zfBgiR0F/JICcZTKy++v7h9l6i1a2HZ5kHDTCKQ2xs9i3
6S7BFlipkgygVGMu2rA+jx419AxwzzscQrAOiLFV4Y1pYvPsHQcCCWTa7qyMK5Tk64KvH2nBN1om
zSouByATePbxvKcvmVJ5YikHvez8e/rjh1o3Yjyk0oXkA/GSSp2nSzsralmWI1NVjiR7IQUFDV+5
E+Mw4nVNkT8aON6xUipTW+0w6Alt1ZozmLWEAAPfJKk18ltKGjxC/NTpeX/4G2DYZPOSXhwQc2/l
+4r4LiGkzu8sIHkwSaE4CBKQQfiOJSXP7UDAx/74gz+EJJ+URqffEYNh4O2O5y165h/tCFNZWC5H
Oa7QX8VlR41moeA/lWxWb7ePpC25mWN3BwuZARb2JViPRIdL+1TbAKinwLGKbkVI78e0v/ipjuT+
ZOpQZr1fkZ2xu3ZCLFa3Ur8Dhy/sFw7VvGyqMIysYdedzx23auCU15hJDaCCcviNH96guncXUX/D
gnvBGtddH83p+IdcMMx3ulORBNqjO3OKZckPfrNkdtatLD74QWKdxDrjZVjtdPIng+rdQsoUpLIa
x29BwJSTHLqsiNUCwKR4aNkxp5ky0KdzPUtly1AbqZGEC0LKxdln2a6U75wwRm78eWtjJSditkcG
qcwzVtKx/JbtcAIqblMbm4W0wx5egI1nzBQiSDjF23bbMS5H1VYaaLi68qZ50vL4ggL+irhh4OJO
Iz7YcF3xU1WQ9WvVbGS6ohI5jXQ+GSv4j7BjfQDfuAfYmgBy5TvQQSsrThN3oIph5Il5jiPRgzsm
EJeFG+NwQOU0MnepWvsiAG/42FAJZlcnBOrKwJdYKDvfxcOJaIyfjayFs7XUdjUZtjvA7A+r6gp6
rQn7hUhiLT+6rwYYvLmnjirhyGFVfpLQvIEeJ9NflceNtdi7ZhPWx3+bhh1pccvP4vJ5Q/in6j+5
jJV9tBlAYjzqk4a2l7TzYx0tET6z/doma4jq5ZnkF3Y2eLvAvt2j8Z/HKGQmWAT+oHOFZaFVp8qo
eXa3yc+dsgKrLkw+FevvwFBgRFcFfrLuk8GTS/CRdHkRcxv4L6J7IOC1lbPMSdSEyvRYAxA1LpUO
linGzbLZ7u5QNTbYN8RYaebyJWmoz8o3l3U3EeuHIq+bQvEECSi1zWv070RHAlNAPRA15++q6Ve9
p7GdL5Ps/ncM2fCud4AXv6obO+RgVTV/7ZZk1o684NpAXDgAuWb8TIa+OSBq9aY79XOcEHs3UjBQ
xv7tY0pdhqZwMhKoAkZMBDG2EUg2XH81M6NRl14ZZpp76yK2SPHfEzfbK4kFZz7wgcYAGGKReojA
iEjH2oWo3fZ+rO2zQjO1pgmDtpQJtRI15HvZ3MCPnW0Y6Keuq1IlYEFfFNAHmypvB7gGCuHesjmM
LNtq10erNcszYBXEPTY6pxlB6Dv68lnh6Mhc6L/TqaIMbxS7ZpVfKb8cqP4+twM78uJsZ9QKkCnT
EfJ27H8KkEAz0PbfaNFLyzuJdGbV67g9vMrukgsHI+qgdqTscsbWQQgVgwx2MX/B+vGWxME71F+f
4V51ievYgHvAsnyHGeDh+XkaDdJvNIGa6M1YWXeIsuqH//7px2Po65vOSIE5HP8ePZYYpgJCcsAZ
+3lubH1yH1L6yxW1sfSK2F6jAxcRV1f0K4Q7l1PVhw4OqdekIg31vA6e7uPV0K/KnExXhtteRsoE
6EiPJAGg6TWIJ/MZgYnI3aBS6YzCyzRI6bPpggXB/PXv7l0rdBMqUJ4sQ3DRLSqVzvn//YysqRgY
PawrDZoz2UYciBlml7FNCw3VdpEfPxmiT/e3LyjJXpsh9kz7+MMeKpIR10vQ2Abu1IMI094Fpnhi
8SuubrLyRmhldyKr76usdSb2a5Nh0oKLtk6bCWTPmVCmt5M9x5h+F1NntVPxTvwnMuFKFo0J1Rm6
yhA6xHkUHPPXZ6FxOh5UgOhpXcmHlYx/l/l3QKSfTa3e0HzYj9L26By4QaEZf5sjRUcYYZa3cHnr
L0F2duC3RG4V9GjGQ8dHkpH3Uma7B+7ZQmA9v8k+ZoTGc68ajeSuREl4y8Egee6TK2LsD5QXkjCH
xEHmMGay97iZIsmY9jJdLfAW7RlpYZTHKosZPcSYJtJCKitgjO9GDufgydS349X8zxt9Hrd3nm+P
BdsRo0CqoUmLlVRiD7DeJFNKhhc32celOEO/Q84g2h9LbGCoqNb+gaZKxKzpCBohYwr6kU+ZoUrf
gso5juZkyaKyLJvgOMHr10OpftPzXvKsXSbPGSLYhGj3MNWey0zKFe+5hTTqBycKl19CebzS8WG8
iYSNm7AeNR6ytVgHntfEWsmo7YBD+/wJCDBsVzd+ijSzc2GUI/D1HzKqq8qz4kXSVN/gKCzPRTvE
sMcIWDHXOIKicpT2wu44roymok51rx8+FzJygzof70ZqH4300826gsB+cHHZSigaqb7eWxgicVrU
vbUZweLY8qvNjGwxvWlbHQzg4SLHii31baAvqZ8nT+GpJ91QdVqwnxMW5XgFHMJLX1QoCcLzCsye
nc2ZpoOfZ1bwzp3kKvMSIijTN+cFjzqUiW41A4Ds/Iq89ERtLL/iPZrIzWNhee4BeOJczN0II5mr
qfOQTvhj5mgZDI4IdTRgWWouCQw39soxek9IKMeN2XpMFOcD1BXh9Zohnhi2I+Vg3NGTITRB6rgy
ioheq8wksFx8leRi5LiMDIzXJ1qAOf55p7ggrNXLkiIDvqQ5EsTNAo46ejI0D+H6wYLiY9WQye0A
WHbNHEpc9qH60uyRLMJQS9VENe74Uem/5JrELiHTdZNUYTNFnc5ce+o4YJzB6XK9d60E8F9SM/I5
G7IPFfiHwMzheKps7Dd9tmyVGqeWa4V8uAuIv3w3JfO5yb00uutLo83Rt9/UqYoJ5asz0KhFcXsH
LdCIsCFqMzEcIEe2wHXa2A+ZpI6i5A1u5dcfHHS/RvUKXqihQ5xeKQGwo8EhDrbM0XJIwr/NmU3X
XImkuqNvJ1UZZsDczGgZJqyVZYrJ4QQWLbURMfcV3nvqeAxZwFLoPmsihS0Nve4Et4RUGurAmYpi
qiNqompo6LMV8x8ZMj2GUnfUnjk3O3eFY9Oppug7qcDhEd8RPFDxUAW1IcvG4EsecnhzffWzCv7M
ktTXhZu05nfX100H4I0ZD3NQqdl9h3aJABg2ftJEMNU7jqA3hbLLg1EKqtaKYG7GlwU+xk/RFbiO
cB5XZmI6hm8Yzg/difFMdmI755RKcrZXhw5/1GiNalGkxD8vROjI3OaSHt4ZqxIlfK4riT4dDbZs
sbVoJs+m66gR6RpKvsJHxqaOhPH/YK5O6ZAX0hpxXIj+uSkFvQKPXFnxDI50p8SD1jQl0HcRzqVi
UxnaDhATiOTKYchZFThlrGI6EezkZmSMBkt/redW84m+HB2afnUOLaJmiKGU8JL+Mvf+UJy4EseZ
yMEOhyeJqN+HXif/dO3z5uF4ScJTK4Se2DUSpBDrJVv3HxVhdXnQ8pMOJ4+r+CDIrJkQY/d9G2Vj
yW5rIJpjhtlZ4DJc/uy9z0xGQJ2YzLEQHGK/phko5Mr9+dEXPAHG174vaqj3PgkkfgLOovJJDNVL
SVdfCD4d6DZS/kTnAzuxd9/m1VmOSECxj9Wp3Q6aPgZs9p302uOh71tVRG2p28dEecD1+EzoJW+W
kh05A3cwu7edtjs2ISVAvARLkwBNFdaKNN9o1Tp5bcRaBE2mxyY6YqhadmgM5qDWBlQMBJRV1+/E
lZGf0MRc0xdHLW5dK6niDFeFgpatdwvOiDp6YGR4PNtHCntGAeSfi2+Y1reX7MkHFUJ/2aqkPnke
YrLJOVFk8qctwgmJihGfrM8d658lZfAMbXKTjnj8454DGSbJCVwKbZUvOgczav3celcFt6sB1psH
GHudHZ/rHjgxOUlHf/n9WP1QhDMUGu4ozO4G6qoEMVJmCqyTu8wCRgCW7l7ExUJlvTQLlbMgUFnI
lXKQIzpxEdIDXAi6q7AMLRaVD5140qRN0y4gcvhlLCsfB3+1w6fGePAkrIDYGM+vUPkfpJy8Wo1w
JVZm3d1XYAkh1m+kVXrGEZbWSPg/mf1VKodZgK+6A5JCL7E1QEqzEzpe+W0OnEtX8kmNzTeGI+Ik
CEwf9u/+oTrJbYWcWKqo25x42KNDcBPcPYrDI1lAIHVGQGZqCqp8tLrRpCIDSGesB5uA5Gu3BepL
iOnfAF7IUFQqqWb4eHZpWBvQM0UHpHhm0SfIewlCBtgLEG14iBpApLlLWxzh4NdUGxVg7EN9OSB1
kZ7q2lUB6gTd39atPk8fiaXbpO9+RHyvS8+VvFqclRdFI/WJwq1DF+108engwVcuoRRCuxwKPh/z
wWx0/1+d0hLWhjySkAXa/rsuMJmZU05P/qwXJtNwxvH+9jbm1fF4P4YjSU0JnppoHTzxnrgpJ4xf
v96Z2cKdC2u9POAHvnSInBK+RtqknX+DL6eBUjDSWDX4D180UHWU3qBrxkgKwJrolAMBqzyU9pai
23EdTCk+vFPhqaB4RAbJQ0oQo3IAVtX7ubnd9yioTn8H7ipel2/xLOWUvIWj5y6SbQF+hpMjivTQ
7BgLfkn70rwoREQkYa1Q1FfUK4Px9zhQbmlrFIMDpDosevpjC6Eh+nzRJ91BELUxO4Wo9GTw8EiL
DfolzIZY+j9ONabLOaIEaNyaH5mIlzi2KGGkFJVTNXruVPRMLc0gOkQcpxkRf+MiKsyEQ3jOw54t
P1GkNZHUxFIvTEoEn1LlCQwgJ6LeS7n8wR/dkptZzhrOz6a0VPa9vGicFaD8OOXozqFGgFBAxIE2
cNI3VKahPNI/a4l+dMPDvB/cdMhyKXP1+Y/xryTRSKwxF5mr9ZvaJAOdW7C807gRgjHKh4BtXoCP
gi3MWBhAmGtVogB+aVM8uaETIV/DzVSrSGHZdKjvHGvLeHtH/sG2+LJMYDD875T4TYuiPdOKEGRN
f3BZca/NZ2437dIVGmv5q4rjmHKFa2bZu4nHrPEvq/yFge1vUXDmWg860k0dnkxN/gIXe1pH9Jk0
ScWs+BdVw25d5q51DhYj2NiGjQIUsm6EBSIFGNMnavgERnkmELVYxlBGACzxt6BWrJfSXL21L3yy
gOXIQck45pi6ggov1kqWNN7CcrTpvqV+Ulg6xhLfW5tAzsFkyE7SlmsWSEiWAMi4sUL3UzY/K4L/
HhYYv1i1F+CItn1HrX76+V1ZTA2Fo0c8QDpRhkSk84rmA0fIN8uU6Gwbq1vALGFO1YgBwCA/K59P
TmpJ7J+YgWG21KJtLUbO5B4aDwhz6TkxwT+a3vk3FjZuP6xPBq+HNt2cHDwIfpQKf45gRC8jn68X
3YT8O78CnGsN77OQGvxYjx1gKlkzTu26aPI6zE9TXGuonL9NvF3c/OZPGrBynciW1b7zod2BuZGf
C4LSw/eTRmo97BQxz0muiPRzLDQhc2nHbkFp1p9S56wUr8r9fiPsBc6SZuO0EE500pNLxhuR+Hbn
670rk4qmbVlx8AYoi2sjSPhnPrYapvyCN2MVsU6nxuTVVAwJX+PV2L1ztS9Af++4GUVea+BEMqrV
Xh4l7TRye1e58M2N2k/63xsookkaB4FbdW0yu04JOqdcHqgqPxvZ2TLAb7tMmvf/MqFyImVkdYUk
nSVTh37eZhO9OqSHuVXpGg2ZlcMoVxxLVtDCcIzA42O2bYJgL86f+rVt+mrEQ/aesHJHA7rDxASS
kRqdPdiHm6mmTjuu26kv6hrh1KleFQewdY+Mc3h0WZJNKbinrGvicQbFTJWZrEn9CGzNpljoJE12
+qt7Nv0SlKanccqAVOf5ow8bqEKqmsQJ7O8Dcgcg4xUplO0KqqhX1ktqhajFxU4Lq0VHb6TZRRCD
ZLJmAhEQP7jknpuDEya5GEieExoPJMuFRkPdGtwp5VqQsNAvZGW0l56kHbm8KeEYAglCWjaRK5Jd
5tYlQsTVkQbOKuT2TXsBWEWmrPVNgCSa81imcAMYHtDc56t2zUBf2mTIShaVQiMzL5E3YOFTDi9m
MarXqmgJOViMpQFKhQGeq1p2xWX6AKkdAelqSS8llJpx1G+Sk/yiVdHA3PSvc4q/GmxVnAbJAyxl
aqUM4HE2NrbgVhWNDlDBXIlJIdwvU1/Ut60rC6L9H2rdEEnqSuFscuwAhBiNXEgmqtgNibxlIdv8
1sm9yrRv45CIlxV4vIRIOjB1YZInOk2Zbcw8GOq7xedeXYB+GGY0t0IbldhE4kqfTHhazsIQvgTp
eqfc2O53zThmVyk8pUbgVofLpDBBrPvyBMvYgucmCAq4AHuvqa66aHa/SmgnkPQOb+23uiqf5c+f
EXRS300/4L3oq+AP2vQe06wiJb1h5/OkVMw00qGAH2Ozz5XesvBU02IlbzQ9+gcJhTxkqxIbtCJv
25BYJnHlSXMiBdIn4AiCYG9lglMX/xqD9hjbn3xmOsdLcF0REGRE/Vgqe7A85++DjU5i5Yp3pUwR
219HD3ONG0ykdxf/3y+OC/2jBIq9UQC5sl/+9eNYUmEztkjIDVIoY6cMdecXfx3iieQZ83qYdXVO
+w4yPPwm6Cq5t021B41EHW6o3IM5U0xc5y6dg8GWtk/PgAXQx/g1II5KFDzLK/YjEsoJzSV1RBGh
bNFcN7Hro6e31sQ/u0I3sm8XAwFys1mHEHkmlLwzo1jo68ybklbkRqebbZ6JuPibbPZomQIdPdiK
qIIU6ld2LUc5JuMa+QsMJFunKAGHp6kdCkU5xTnZp0x8LTddnRu1jhgtKpXu93tgtZLlcrH13ab6
2VVx3ShWN+zw0FgyPx/AsgsKjAr1eomtJCoLSuDMQnXKXOiEirD07ER7qcLkGqRcG08saS/1Y61x
xbHaJvtnHmXOXiKanLBvSp4ZJznLWe8FVehHujA9rhNlJDWQAoENDK8Tt2S2WAliVNnBdtqvHCRL
IzKvQ+aXhMwI/5hRZBua6vufuabXkOaXh5NtBNxs8ortUkWlLyDCG1qtYWeyiWReeHeBwJG5E5EO
y2DgXmfe4JWx1E47P0qtrF+FtduJjRGcu6yRUUbbQ8mrBSq0PSKLra5bx92ufhAGaMsHRxxIpQvN
dscEmV3AVP+h4qHIZwysybedlkkU/HNa0WvsVcNiYiW/xWSg7TxUPMY/2B5suwBSqsSKvyfPcrMI
B9HRpq19Xomp3X/Qjce9S/SYFzHVjR2npF/YyXXfIFZ9TqGbR6BKharBZQ2+XT49hK3YhtEsMyqE
ZyWWAupYLwOJkGCvFqZ/soCtEkPKw+nDL8/TK3EBknEkqOg9YURXcDxFTpS26ni+GgH143b5A5pO
vTQBbMOtMV8wNJ/4U+hYXiCA1quApz3hMr0GtFYgau4Db/2a32ATn7+fORgJbxvutGOkS4/uxrFv
DUoV/XnkkHBwvrJd55IaCNmKRLRjFezAKMN5BSiIyuOnT+mbddoesBSszhB8OK2TWPZrqIYFFQxu
XeWlBfzV8NeubN6A+f13h7B4Im5gY9OnwblwKlM4M/E4JCGG2vyAAo4qBzMwOBGgUG9EAcnI+dbr
/lqvB8WfhqxleAXDu3nHh3xyJZuTzlHYtsXPEpBvuJfVoxZyOdqj7EX+0tQuO90g/ApBrPYvlyLh
G9+m2fkyuT1cqVQcrwD3iEgV9yo4HjN13DK5JjIWLvmtOh6/Fylt35pl/3UoxKP71JTVW9KVFgwF
93bNtgCXl8Bgr2IiW0q8tbJ55v2jL4LhyxeNSER97p52wNwAp2oxNBGM3bSwQpeypkHfbOKyOH97
/PuN0NV6owQBacG8cEHSyVbP0Ez9HdZbs0+Y6ZO3kMeIHNgGJ/1siefg+LFuBTTWGp6rrnFfgSSA
ZKCxF3t+b0i8B9lI4IDV1W75g9tuA/hWPCXfINmXh74hfCpyKXLd8NBCU9HAWLw99cH4GPTp7Ods
m3zUSQJPL4Xmfq3RM7BRUCz8lvnqvSSH2nUJy1Lp2sClJPp3qGsMRKQ4B5oLwSOM5b7HBrhKo0Ll
WndpJIBdKo35ICVWnbyP1Ew2yxOYFjSCvC/6ZZkR5G1jTmw5IpX5fCCldqyoij+uf0HOZdQAl/6d
VTMXa12OCSDb3cVA90FAr/H79FWVtJ/ZHDy1ic+nWKzeMgH9m2z71xDUnCHwDpDYDe6hyuB2/aje
gza0BkIoqMzacsUT2I95sFQoi7Ph+dZRaSRYi23e183bO3Juyivs3m6LIrEShBfUH9z0pNAJaC4S
D57lDW2jpCXP5uDm8Df1DIr1//LmdwYhUst7C83CvkZJIU3V/RDlerbQCuLPN/qBMxlQ3EScDfKl
0kLd+hq4X611togb3BRkpjb1q7o7Lr6j6qzvehieZFUEgt22XFTsknk78BRa6jcCtoMygfU76gLO
uLyf0OveWV0fmPIeCQ8Hy41/8BRJtBSFdt4bbCfoE88PA6UD1lcDFm0lC8tCFb5ZqiYzPDmkCLyf
uvLiFPn8lTWVx+Ur5+7PDznVSpXHvST8oFwG3PSRrMbf1FahKCzVmOr8YRogwU8J7EihvNAGr8eO
T+OfWwBz31+zvkN1PjcJuiF4LJ4zIROQJ19mTnmO+a7tOLpYQu+cgKRZX4IWfbPWoalhc+ur3L3G
YKQ2slTCYpB0ywH/eJ8OEVGk2F2gd1X/aplhLlu9bP8yn8Wto+vcQ0X+CJXDeW+gAvlRG0V2CL/b
A6ex+Kc5pcCXrZwjXYhi/XWHpD6qgV7jiolgvmRsYQedYt7+c8iPGf7Ox+q4+4jcgpCv/Kowe+Rr
3I8vQ4XUv9PkPHrbMfZIYJmNnrHVF1xP+1uuF1FQPNWYhhiJdjrZAdzBoUd7MnqaL4jYLDOXyP9x
6bVSG9od1vUK6XGd17GGZy0MdQGmJ0XTS2+2sZRGeWo+7ApdaA+bXln/njmCcdYaaVoSSovo8S79
78rvAIrj7pQjUezqqngd3BlSVU2RRC3KI9UOX/EytT6+s5z7IpI59QVjpVI14hmWebi+jXM412Gt
4MQaNcX0pp6qt1HvDpE60PLi2AkhjtEE1hSKPGYWq6HOMUgRbRlrlGkO5yh4uPXlAxOj9SJkUfyz
/uSY9gmUcP3djHXq/UMQv4tVTI4Hv9IHJzhs6chRoMMSdihtmzEr6IidGqN/xehJBtZ/wW1JteMq
8ExbFnn14Hme4COAvhdEbTDunAtykTGcJICwQYjacp32NZPfV/6i6chxbMxzTeHsBC3WmWNYkzdC
B6++YwdvRLDrxRShpt7dirks/ttBeKHkvvmJF/Ijxs8VRITLhopWMTMVwioesD4/zHcmqrZHzWs3
pJ0Puubqyjv8n7zrAWdPk7HRTQriG9qfIfkDgH/50YW3Fp7OcxtSg8bPLGp+Keu80leJ6YArgWga
0mjY/LzGLB/WzOEx73lkNF7Kb4WkMyEjBSl84T2Os733eANttzsUhAY66y1JD0HyjFnEG4xy2JQm
oFGx1GBB5r1EFILmzgMmZzM3l1q4yzkHalgKXQ6OfWqo43yajYTsqwARzE9MSow4QiYnRO/MwlwI
CHmSczzPuYZVNPZDNIBeHJH3gZHyCbG7DcbU4250MQv3U5s0HKLMd6R1Yd69ooM16O0I9CjVqRuh
sqIKtGqnAF74sNgm4PVMe/kPwr+7YJQiAJGPhXHXVMA0hb7Vyk1a9M2ANzFfcJi3E8u4VUDe3rLr
MXfvfG3lc7uSFPCgD+x5BlKiof7sDV1d6MHOFksfsCvUwtqfE9oJpZ0EJpul2bhl91uII76RCdDN
ylNsui3RcDE0Ri3bPxv2j7U7vkD9fbCSuP4tfTG4L5C/lsjRQMeCMUa4B5SngPOyFDBhEfORzYNI
JfBp/hw8d1wHdZhG+gLT/kzoiQVjHGMWs56up7WYucBrcuxPoj/mHWtPKmZ8ddI8LAFVmqEpbGLL
PsHe2CFv84yL4tYh9Ms5+fF+Yoa28q8nOkoMWQgLbJGY1EcNgV6JnA5KOhCPLDf8qvnl0h1yLXcA
59eOl7T/j1SoKxhocOR3pKY+wczeTE8kSFgyoFqFV0MN4lJvjYkv5JLK5kmRMQysBZbwtlOIBvsQ
dy5CcvLn7cySDuxDIGoZ54vS1Gmmx6gOQ/PQyW6jwQiWfriB4MXWBPOZQKmg9z79HDHp6aDMgpkT
0DJanJ2l2nUH5kYRoCVZEt6n7fK8l1dQFnZH9mfS1WaVlHl+LEL9uEgBduCNnrO/7T9TciX8yvZh
V7eqa/y5RQ/pWt4bnWlwev+AJ9qpYLQJilD7Ye9vaoM1iNYkoI5NZ1XsqaDDKk7RHAGCrk6gr8vH
TYUmGFanxUxWPZErBvODBwwTXn3/gxJDDeZuWkS8dGcAqVlRN7Qe5ysEwKC5LVgRPOZjQ6yPBCji
7d+Y5IRITJQ+7ZVUDMtL+OKw4wEPQnhpfFHKQ+Z3TMXIrmDURBEad77o7kSlKxMiRJMi4pqtwPES
TEJsa1zF8MI6i8AFtTTQgMLAjHi3AsdSRZ2s8eFDzjncy5/kqbPnehqtu2JzZfHkTzYxTaRIe3C+
xbMnlAjeYBiKbOg4gx6RQCvKwasPJhIxZ5XfdkiRLtnoIFYQU591wMNJzT0wPBK6W67cNap9F2li
l/N3v+b+KJyoBdbk1CyLBwZaQAmtfjj30Ho1s3drrGRbGtm9fxVAV9KPBQ8fcbIqppRDI9RCCjWQ
S8go52F63AtesA4yVPIj2ElW5hXK9MchB814OiiEw/Uu+IodNMRcYDw6hHEX51vpWazfaYKCGY1O
JXeF0PyWXFuW3jrCuvL3yxXhEbPuRbHTj2x4oTHLr98Yb1JgHiqZtI3VRHoNXfT8HMmYHBuHoW+I
GI+ysXRov+Vsu2NzRU9YMBA/ycWARuzHS0jUfwuivyCDsv5vu0VHxrcJ641kJ4pxe9pb7Hu5Jj4F
CRjRAvcyyh45vCgpbADUQCJ/rPzpfFje3l2DJ6ompvFYEFbue8vl6ShdzR9nPneQb2J26TSuSufy
PAdCxXR7QAEp9JcDUEUu1k+bWjpg+5RGe4OSd1ZV/nK2plcnxCelG/9emiqx6nugvAh9q6+rZWB2
YzWc0rhgegh56HWzsAMiFcxYe6wLa7C4TOMYPxS66Ipimrocn4F2ABuqEvmK60b2sqSRAICiw1uC
MB1+3aJ9QUxgDYg9d4b8hHlQ4TJXBVYnM9SPb5nqdRVXuxsL/uzQCnKpB6AddwqReQU/t8Ru7uHe
N0zlCeriCZY/RFlykNi5HOSq8yKwbAo+1DPMOWfaw9YpLaPws1CWyxz17KzH2M3ZDA7mh2MMJJK0
6+ivgvA7O8IT3b1mcdpDvFEKoK4VLF3SKN6GwO30KpRyph3eEZAhlQn7uBBToaKa0yQ1TBFB/dSf
yCIdcAy2R8A6YgqZPB1O8y9Te+Upy0grCjgRYxy6764PcLXKtWp8Gp+EnIhfau1tyr77uHYHUHvc
85b+nI+kXj07+4mRT2oHwgCVxu5kB/ZwfQJ6hoJKvDCQtZYr/RO/y1Bd61G4en5ODmT09TEBaQRh
5FplnUqSf1zHcOo6enGQT4fyMRhmA+ANHuHwoYCDd3XIQxLh+AuLmMNTrSTAlAkQXCzf0S7h+hs0
gHSXKOg/dJJtJRAfJBarSPPAtp8u13f9XWZrh+pX7o7FAhpME6oKwmUVvYGr1hYodv/3XJzm8Rjq
DtWSBclWLJggA8LHTq0EqwNYLvRI1lFzwAdZBcqmPXvXNyiFrPXomSqRCmt5I6qGUNmbW5OgU7CS
iXHFHg0+qQHvoY0uyAh0whGaiPZ79k6/pYDE+k3zJPLuICQYcZnt9M4wchAD6fIl3ZlltGmAC+7g
yZ6hojiOqjWvJRqgI1A4NcHhKY78VqIJCSQOyDp126+lBK+KQL0mBMryLgwNr4+XelmqdcckdwVp
Q7QgTU/Y0ZE8iXtfXKSwBGXN8UJPB0uN2OlQzMlxTuEUrvGovEwQ3RHimpJXkuD8GrmRkxSnitOR
zTwk10WacJ8ePWuxUFg+AzKZaxfG+/eaItINnPpy3fbHvWATjp0nH1cdHTGjxJl/nStDKedV7eAQ
N22tg72mzL3JIzEJQ7PKh01PG8CqpQYqxmwLQtI6D3ws9J1gNTUrsuYbgZB97PmYIaUiBJBREZOP
9xfpzhj9WETcej582OnRCYhsa56gqN6k1b5j65nnsMJFE5FU7YwvE8ZuxO8klqO48FYC+2/kSfqq
GAGqJ1sdLibwiS7MXENglwxe7ZQDTHtT4oOQTTAo7xbDeow+AxXZP6dNuURfCROdx7Ji2EF/7Hun
RjfJKDPChV1Hnc/tEhay74TgU0sFrAQuVZGsTKfN0ykjqFGw/u89uIMdwVz6vi0a7OUvD5dcjBM/
QBsTxtcNpf7J3LV49OxyyQhjfQoEt+GP3r0yVW1wK4xQlh2og7WRsFS+Ln5txFlvnv8bffBTq+PI
Rk5ia/xtPEgxr8Jzorf5MRKk6byZrjzh+2h8zS1CTFxn1yh40IeNYtyF/C0tXZ2Xtlq776JUIufe
Z339WIQQxmkyP88SR9pvQXdX2uPF0V6X0uc7+TfcmWGPhj8WZ5vNi7mCfaRltElACWzwcVMHNUU6
xn3s69Ut05dFBRyzpx3ZPjJ/xCBMYtHKGvoJC3tJvKNrbIppWGk9JDZoUW3xyny4zeBHV8pcvk43
ivaCEjUDhxuXfks1N4iRvxMIoa+bHQBGRbBz0S9WRk0cBKoz0mY0q2EYuLHeJB+rIRgRO0dpCxLu
u8HYMBQNg1ecYuw9zarOGg0v4fToPB/H19yufb9+GUTLVYR1L0mMyTVvSS12Se6Ku4q19A4SBdBt
NTBsLms8EVtQWHIWOKYtsvsfkg+HImsGly8KwWzDw0I9pXkq4B98u1CF6kx/zr9A3w3YMS4gwnkA
IplIY8PR1raPKTrXxiwLIU1MbYlHBUdZKgrNwqI3iRGtONdDMPFfqPbHFgeKg3nPnStFP61+Wgiq
1tUC++fd8exlvaPscnopc2b1PutZP0UqlYZKCoWNIa4d6b+mbHC8jwXdfOVw7ACtnT5CdLhubYmB
5v8QS6XlJU20LswBmDosRm4mnlOkod2bV/eWf2Qodq+FzJKv6w66J4CdOpSCZuGAqSQclx3g0nMa
ybfHs64B6j2W+Ctnb5S+92LVC/DJtKfNfZ0APYACn+F69NuRpoxwNnwj3BtDS5F70t50VeVwxZHR
FhA1/X1I9jYWSpKm2fzDkuP0V0jhgyuP6IlDUTMeqj+JeoK+UB5B8ecRMnDmY6f1ObP9yvg1fGcs
nGPdHjtlxSwGN08ckyXIY1VeE0dSWPXwxdwfSuu+nN3iTiYadd1AORIASjIJd5lvth3v5RrzSRNL
mfjKDR3pmZpzYdMuQwGTcDB9q5y7tOexwjzGbVkaBSicKIQOkFdl5vc553XYbEDqgW5x6NEyQY5N
sObqAXPmUn36870+t736yqseTGsbNf37lW/KpgLH07HPsjxF+NbJyN4oYtxRpVNa+q41aKUDC5fn
nzV3m/yyuN1TWksbJhRa0jA+ReenWEg66cy7uBKv8WYI08uFTU0mQvlFKAmDeQknaOdo82UmaffM
p6wVpVZWtS4dYe6SsfRJX8yeeYSG3pje8KKH5hGQZONclmzVGbcpnBfcIMNAUjMMIS0x4lW+UQYI
TjYddh6bnMDhsatOI2cgVjqbASaJqdgdpV1xVciSRwgNbzXvE/OGHfFEWnZx5WcrxEakjSB2W4WR
mHniSHmYfeKI9+sbHSt05DG9YilZg9Ga6pZ4Xq+bwKBvnh3XIOBffQRDPKcSUq0NiB0Y9S/31bWO
u6exAL61ZTwsBeFparSe9yW6nn38LVwpY2EvfU5BebxaLUc9TCarPXBdcyMpxt9uCeR4Sbxm7T41
WJc3Jsu6b6GRb1MkurV0/W5AvAST1gRfvehigF7xLgQzASImH/XjnKchhuTSdhOZePqYkUU9VX65
2l0CIGEtehh7kk9kOBNUJWO3X6qljCmbKK8oqCiC4VdO/9oc1tmC/dzUhr0o/V26gco6X4SHH3V4
lfFDbEsxCVxj4ZWUcBGwk43GXboFh9AB6axhN06hx7XjjKY4WyLO0eb4LZs1qUJ6cMHUXUSgEtXo
8xa1Yd4neUFVG2L6sbeHdU/ItAlbx5oUoEFLeo5yLWlsQy712KVIy+A0tQXT0Fea0ySdnkEIpC/3
X+BBz3wBEg3lTLyi9JLeXkCuvYSRfIOJA5TtSpYJCafHX+I6tNp0ezRj+A7TW/vehPrD14cCl2An
gPM7ohjtMAyGUO7FTSRTXug4I2rhut0skqI7hSraLJWQMRwiy4Gf24YVfDszg3wMjGjUWCwP7Ys2
Y1IUlZpNdDFADNQnlO7EsdprJyB1N63jCQzGLpUQPM0nosEj5FGcbgJAwncNnbTMtTGzuIIMAkOc
Oqk81nepoIoSONbwMonWaaHZ4bb2eEYjjnLM+y3rUZj+I4FRZ8yE3Bs4qt54qnPqa1KIBZf6dpBY
rz5w3Kma4xIRgxXHbYwbjlRQjTm90jgrcHVNeZofsmqRTFqXO06/aLuUrJ1BkFz0V5kh1123Za9p
JU4Ph30IvVRqkcx9BjbmHGFGM/EjpUIFL6gfshsYwXDOjhOQoHj2/mbcJuWfOR7iZadqRUOqlEkR
eIfExPPXnmrN7K7cflLEmGiRnkat2RLt4aakfSQNlesLgXlPwrj0rwYJ0MM6Z0uNYnFC0GwuiCuk
kyOjZrjDTHK0x/Srbnd5zFSSAcOAVuf0icrRzFPFFmedeKcUoRpIWRHAPLM9kTaPsNkd0oYEOAPU
hOKEkeFDtK0ixsDrebjPxaUjAyubCoSWxQ1agn21UB6nHsYkaPkWCoie8mdN/20xidMmLek+CVou
KIJNHlxrhqYP86IWm8ZjBhypw3QRvWgxBs39/dk5uyp6vfgYMH1Jr20bhFidkFzNP7sLEUFdrZtC
tHsjuicmcmysCpx3tkkSlV56Uz+EGWOHAgNPa2c86fAh78ukdCU5kpgUR5I19oyQ+uj+VUyH55JU
vrAPVlqLfKyRpxVQNFqpmeb6kTr00HJScc6gO4lVxhr3RZPuxru3v8YobJ5jsr7m+lvIBr9o8HDq
vNJzN/jlbP4YWqz40sMD6rDlQQ22+EO4SmpAYN4dsb4EJz732Xi5W9ZdpKhnWNf7IM6SRH+EZD+T
t5sOZkf6SB4wSCR7WbTtPyyUU15G0yWUB+VFZ+gfWWOkYCiSYAanjBxk0urK9q8oXSynxiWQi6YI
YGsz63Aew/oQB/tG66sDoJr6jhhEKKRNaFEbubOYA7Hp0I9aOJdSF5WbII22W/zI17n98yXumk92
B2ce+NqaASXGwfN+V0Y/IuyDqtgEZR3WwirSqpPh5hgqHCP93nYWFSZn7Z9v11IvAOdHN0XUI70I
AmP9V5DGw9A8Eyym3VSMt7L1dDfFq9Lnr7tah3tqOpRQEPvUaRGI7tom42zF9jhsgyslD5wMDrdm
q4eblVzu5MTb1AQ95p8xybgpkhO7AXl4U+xO6KZu37JAPxS5DAO0gfaqrhF9eKgjQcwQg1SgOLtC
tOmY4Za3wteLGdRn0AWQDXUN2IN6ZE6POeH137dr8yU4Y8eqhSki5PiOzM4sDXfUuJ396XaGiYsl
CibdVlMpIK7hht7JRIE/sFWVLuf8HcOsOlcQRKM1GpS7jY8vLWYTjytdNtSLtNtv7Te3Osw4LHAY
dR2hO5O53bXjD6m8Q5wUOJ/ClZZojPeSrcwFnKLFIFPUpcktIAXva1gQ284yN6beJX34GD+Qr4i1
9Kl5j4l6Ql4+GarxARAuAQcOUjW0SrIsKOiJW0+n9c0OV1aN0/41BW0eOyIg5XDVLBEC/VRMfnFb
Lb1aqDETC8hgcCJSgyJKLfKpt4wlP44Dlh6p//G90cxswh4r4UoyvsatMdQoui51bPN5pFWF+nwB
YzDoS2VvS7/bWZgHzZdz7Ws0R9613IACGcIahsrGvwzSaNvnBLFNc6UzkIUKrKgDxqwL0mYn2dkp
Z6bMMGDjIXC8ZO53ioQeaOOGFeIbSTWQiC8+tdQI52jOkoZfPm0TXZWjuDL9Q2hCiKV/iTBvn72F
F9W7F177S500jDJykLGuCUsCOuD66Xw5rpcJiudmFigZuLlbtjo2gZdpe37CVn7AR5uxZUTvKf5+
t3OXm3tTUWFbjLgs5ydRXhPgJFZa7puNYoEgJdRHYSuHKvMmSbp2jbQxLm1qJlLznEl4TEeP8GVq
YdojDvG3PEVqEXLBBhgtXPwjHKhX0CZ0LLD5euv269cBjo2XHSQnL15grhRgrAnyKCDlszxcPSgb
f0QzPmy/iMPWj8tNqvsgWsPSvXXGewHrQz1q8gIQM0BGLFKTDHgWosTDxvdtcjLSPcmCVX2LoF8N
fkfUwhhZJ4+5gaEM8MKRwQiOcHh8KhScq+LpviRMjAAGX6fPeXLMAosmiICPYflP+MURPFd/A+lC
CYFC0b42mWokZns6QBzL8cJS0qm71iRTHiCdPleSBXROnEw2N4MTNmYlmpB8QNb+IjWZ8zeJCU7E
dRVX5NNavbkR3hX0HLRT1O/fMX82VxVEt9uRXL9H5i0ccEleA6jA+JUmSo/avQBYQ2K/9BPpJpsa
5BvLXecwlHaLWa8XUFDNPmQEfDyynnul+H1eGpEDZNqGbFU0OutDZEQwi9xhxXEBPisHry8hV2H3
QI/twtqzxWT4OPAoidihdR2KjVq6dG3gPlSC9GQ2Kw5/+LshOUxzSi92tW7WvK26+vJvHUtIcZct
ij+gLAf1RVi9np0AaiUNrSNxOHzgJ3FUpESpAwpsWdZMfCsNJGLZV1/10ZRtp0OEGzHbSngP9Si0
mGYmkZifoGFy3U3s/MDzYOhAlANXV1xZB4UHhnhjqLjA4rry0EkMZkmv/UlFKNSZbDXtlcO2xuC2
wWPg+64ktdEpeQeOaPZDKS1C7Ye7PqIa03YCoNchd/Q8afK9SrG6aKVoyjwgRNEDSOG/StmTRiiZ
tVYMoV02du1kovBIJX92L6oMNvJCesyiwMIBVQEWS+zip05XGYqGozhF4Jf4XKo8xDzkqhvbNjYs
DPDu/ZIwO+qf1q1dZYLt8gBVzpIH8FgeTPWMnKQsAnDkYFGb6MacU4nTn8JJJMfGYrWh4aqXBaXb
H54miEyCWP7vryX61kLpegXfzbFZS1lD/qGzoXEqbJ9OsEEfv+RQni7JicsTvtVpRCf6BDCfwwrB
gGRavpu7sKyMJZ+CDH9NY8MVLJWJXoNyLyRiW9mAcqfRxjBbUcdQogIFzFNwEwme4ylWukclHbnM
/3HG/0v4XodKDMA1uXH6JKrsjW+kzmHd6Uk8V8pQa2exJqFR0WqdKYiU1gK4gvBIbG+fiHOtjeAD
HPo5290XC0VNeyEi8JHydjcTtYMsVZP5Zvz0A4HRVdPgl/SFJi6ptyvYKA51trXroTMXQbnSUohR
kO7Q9/XmyP/pe7k9Uz/n/UeR6yJds1q3bNXZ0T5ENPXreFn7uBdv6HofQRdWWuE3YdoI4H+R8mEq
ezXAeZX17uXyBnniumX2L3/39glIxT5EBMbE5xXprP82BocOIEigSG2BlGLLR6kxrTADhn30Egsc
5JWwmvZF4BhcJG2y4FjU0DM+1xiL2q6KgJAyT5oZ+uA27QxxVEaqGVq31dBecM8tSJhd765yA86I
u9MUpQMjonhRSWQzj83nwtPMe8QYN8fWP1suI1Lz+D5EZB2olmhAVVvqamWFgxYvE5e/NSy5G4dX
tPw7IJqpZMLJqb7SAGyJ1XE5lxMyCWjoULvzcSQKAexFL+By6Hvu6Kv28pWOlN0mNuPyjVHw/D3k
7U6fX5PoqnPrle+i65mW3nAOkRclA1pU/FFDclv5H2E1iPr30GpkcJ1tsba2xaKBLGWYx+wrQ7Go
uCu/3Ncx2AXMgsw5PXpwgCz4XFZ1YOTjutQF6dlgWDe32eGWwLxn2qw/PcBWekTuaf27Cr8+ZEal
g/bsG9iMN9y7wdjpOtSjGFuDnrRj67NFrv21pdj6VED1LiXdJtm817jaDe0jAOiGGLKbKZSKTvGM
65StTALov1L6/IU+KcPJKpXP4CMB/6P7XT7uRM+Zo9a9K8ub65JvvEYoDyG7iDb3Ldzz1JjHwnOS
lc+wT5lqGYKR14At5sk2ucf/9hNK154Dao/BK5a7vB/6BYBDnz8wYmYw5sjZtlD3Y648ATz5tppB
adk7KLnbKayYKXNyPNCQC4I6sNr/QXyc4wOhqMzMMw/APB0cnPG4HIXeeJgbjFrRirLuGlwLtLkn
7wmGQ1/pVBotJoHQ9RoAaSeJCN5n8a1I2RnCYCTfQV22/WlRUTKe7BfdbY5BpOj6PLH5CfbnXRYy
HE8wRSKQL8bmcnnzyouij85GzH5zkr1fjyWlc9eRLL/6zL8nSgH4rfEMto7Wws3XLEQ5D6ysulXY
l8mUa7A3kU8hsKQtdWg7rZ/1BQLcfZFOQe2PW/eEI0JyXVxmDIdouaq1W//26rnvYHRuI7Sh2fY6
uDIaSNYAK9Op4c4vZk5gbe+iMMMMBB43tWID5eJJ4Kzx8HrSRLklML9a3H6gHYX85LELfUEqd7E7
g4QoazKHgOlfr+9/KtNe6khjFuUHXBirkCAHjSdcQpu8gwMakgTbjyOBwOzwp46U4D4/h43wYhi8
/MZ3eSUhWtBR3vd+Yj9dTT1wv59sAYMVUqPM1vEf7hhot3bb1Y3tqA2Eo+fxOieR2PCyCf4C38ra
n/bgtLwaMNP80WYzdm1zjMCkyG3HWPOwcIaZwnUSYzUoiBRSRadOsPBj68o9SUU1hCmGmvKEZ5sv
H5wW+DjOr6gfkMDXVrfZEqelhF79dUBL6XUbjhePrMNGOrGVomiNNOh+PlSOFmI1aYfd5BlCJSwB
fZrV44m+ydiDZtf/Y73UV3ZJ7T6N5i/PGRemiwbablH1pCLtq4+9SuA07iEZUqDCROeGdwRKvpxs
zTe1oDEOwvZB2jjuy7W2Ouyu7fY6ZysZ2FRwzN1L2rPB2R+GuVOkbhfHXrZsSq7dQ3flY3giU+rT
Yqiq+wKhgbEtCdLUR28UC0+bCLi30YN3oQheOk+zN/55DzgcH2REXSJHU5bXJXyV4LJL2T0Xr+JH
TTwkwOkU103K5L4ZFtgepGv921kEdbht0mxHjWwHAQ+oa6YkQSaxzgrOWchwXQo29QPuXazVjecj
QHQBqw+CcihNNv4IpZzPAOzZCcwg9SkGJXE5jjmpAOINPEH5MqvKlk9dVw5gqpC9K2bmt4tr15vo
cHvoP/lkDuqKyqValxUN1dXtaUZM4bhgyfAleEJamKdJhVJOUNH6Wnenjx6QnAZqT/2H1esHzkYa
k1NZikBebVlSfsVBDH3hwphb4ti8LDt+Y9Fr0Acee+tlGdI+VhHXoOzOTpceAs2RFGiP+eAk3YRt
sxBU8c5BrauSR5I8KgNvX8pqiTXt8fMuOKL0ZD0fLOzl+SqOeyGHanXaN1d2br1eQQD3NAjwvsmR
J3UjJTmeYo81g43LvaA/cDwmLtPCaj+55l+o0+p2Yt9XjVYxcHfcEbQl4VaaSjmVE0wIg/BS/s7u
nmVTwqBIa/OR4ZQEB6GqxiGIJmpAQ2pmRLK+Gc8RnrXsPHnl77xksimaVsGwx42zGv4SqrrGh+PP
0dwJKGnLU11knDIHNJdnW0oCnwVvEAbrJ2tUbMEqiSAnx5BXSZtbexolzi7WxkrIpNFRwvIjbef8
bepKK1pV5UI/ZiDZBKAPhECljj7M0KC7aJFoze87aC3K05IhRJDQZZK0PTBTPnM3EjPV2yR7O7mr
vnKzm2yXVpGK7/MdyvEmsbQPQF7S87NAW4lxhahIJP9syz+UdAPX30lciUf2QxJRc3uLMX2rVrfY
v7cDb/FiXQXBV/2NpdOGDB3y7T6v9Q4U3ATNYuWIqmNb12qzVWAztne1ijASBC2l59Cfb2ZKbmao
K5DA7MlXXZZoc8of1k173miXAaPKZyefprAxhi+It0kE+qdErFBTwg2OIhMxMWp8HW0cAo/FxA0s
3T5C+XqLMVAFb+GQsjuR+nPAU8+3sitk+crReyUZBc4wONQlzBzDDwW4c6M6EUf9lopVqXDBdYJk
5u8oMYAvuR6BZ4EJUWBfV1haGUkaudqM45vh4mWV+XosUxxOJnKUe5YV8HzOPEp6m2AihXft5eqf
KgSxGSZ+GsIsYLI7xr1+qHdCryXBoOJET/IG/vwwMeuo0bNiSn29dhV0l5zW6Qa04wyBI1N/g9BI
f19VyAfLX9AWEdwlKgGTUZ55b/U7H0k8/n+L3QIaqfkr65qLNGz7z33e2E0hL1qSMfwfISa40E+p
HS6m+lS6mP3esJWRK/RITJpiuh4elonneQIpamXZ9AJ1THf2+rSU9UFfMrJHmAtT/NaKB7xgqwEz
I4dJBiJvdMysPu2m9Ko/CNKIzthPKT9g/LA36xwWb9kSUm+Mns/TmdPWiXIXB1LA2ZyLEtXm6W3R
kr/meTvSk7D3gqiS/fOAQ02pKf86nN3dsVjWSkvAF53ZA8HNCRBp67iSkSWatcWdceR15YJRCjcc
06o+2OY1xtZ0GVc73PIshru1PYu1UWTkqPZwynFUVM8t56kwB+H/+rnx/Cx9kr91TghywsRrV5Mm
+aQWFq1OVo4HaLd6ZlA+KUDdYphDh9rEHOMdpuNjAek5ClyCLFlvCzbIJhRhgL1O/zQZHetuRRIf
vE4XvIiReipaHEg5dimjlF3VD/cDI1DzzwuZEI1Lt+M/mHSIfzH5L45z09Mj1x98gpbGoNr4aa4r
L2Lx2V3/rsIL0FnfmwaGrUrDHjIWTY3ETJgN15EGcO7oiwYLUsJeDsoo5HY5q7aZG4Dqg87ahM1u
3qUO/WpX2WKo+KrDhSO4yNugWBrajeMh/9J7aNeMocD2c7NLTb59sNy1E5J+SUikyHswT1GM0Rtd
X8g+kTzisiTxfExORReNowwLZoZXpZBc+Z0pTssn11mEFNgBfmOh9RCbVZr6VWlIK6dKGE9w8CSF
Pp/2vISZ/CBz9P12Mdsm510u/2WkOP/8vJPoML235KoMW901mSGr4EnCOa2pSQx7mTtoqMiog3mK
s5YGgz3VOgbBLXz6k0J3mjUn3/azUi+nSL3XHChOfdlFo7rZRMpJr1KioHi0sQPG4xjh2oazplRb
d/0GZqBsQg5T9XofbsLBfkfbF/lLyGaVrZT8s0c6CfD7IpB0NrXg0jHYhZLOJ7U5xfRUPLl8SzYS
v8CYJPN99dK1B1BUbxD7o8TtMHpqDaEgOLTfVunF5P0hSmyAY1qyWNpdyoa+wPNa5EWrBHyF9cl9
T2Mm1oclqE1y9e7Hi9F05xlS5MUkWMzlv7cjCmMy1hnuRe66yP2e4cxYEAa9gHH4daACxt8KEhqn
rc3h96152/OYVwE6iF3Cu8/bz0lhA9UrhZj0Ftweg0Sg1ZgcJlHXB6Xe2EhFOy+k8BV2o1STztTM
bRg1lCJ668ySpMkb3dpUOjcziVGm8Mm7G/z2hxMXsIGkF+XDqFwTvfHGvLtuzt9xd83og0ehXj1I
XrEReGKXdMx21vw2QSUTNdWGp1vqfi0tKD1WxoOLurp9sAuwPRCLbvgTRSHj0ejgh+iHN4tnPHH1
AuZBdrot2NqFjmi1XoE456TbaEnm7EYOH3ue7ALTyi61KW2xoHjqIIyyH9Z1t7TMkPyiXtXa3/W9
snchtplS+khYogPZWm6KNPh8AynHZjHbVwwdZs73xY86aA0xbor4zAAh/rjzYeDSWVcES1hdOmAY
A9xQ4tmCHumwaxpI9s3M5ccZkdrGW9giwSGK5AB81Z7K/mYmPjXWIFS86mnN0jYtryzRQeuX/H0f
ZX9Z09qjHUQE6H7akK8gq3YCeQCQfY+bpEKKtmV7z28pW6FqHbQWa9JxxwRFiJw0esxr43p0nKsg
2bEOhs0FX5F3ZBswq7FK20zNt2H2+D1jjnOF6hipeoI4jRmAykmBjWOarVta+W8FDF36buteXYvD
GlkOXGVRToNP5pQwPpgPvm+wdeVxG04sUT9V6Sn8PRZmYBIHVEs3u/Sboz8u35OL0TQYMCOXWCqx
GUVbqg6y5cDIRuLSvL8gyCm5mryctwyVIeA5OqsLjtS+dDAVWy0czfttO5A3hk/JO9/GG00GiFMj
M0sVVyAH7MtKY0rE8wNMSZ6gk4p7EXTb31ALHMjGi5rRs5Q4EjaG8RViYK8HZxd2Kdnxi7n9KVR9
Wn4HWDGFaWitKPxZexvNlOrmn7os9pvfLXw2ZfrAwRFPlqbf849FJ7KM7pS4C1Uk8m0ZjgYy+DYy
POmaTZ0Gf39Cm6wsEDbL6ynMF3OwCRoNa+VWwmxNesXqBg1LCpP/eTw/rFpXKJ7HYJ2qwLz1B4kr
TElGcZLcPw2OnDhLCSKcJAtv3ye8iY6g+hdbQjT0OCGFSIfGpYJIgw5NWqSr2LaLiPS1MYry1Ht8
kcXTT6rf1iI/pZ0NuE0EewjD/Fy8NtPIvLyEMXf2iNOqotXNkZcZqh9CnY3Zrjq3YTc4AJqbnH61
bTHrdCXFnL6niDLJjVP05e5/SzgLVenWgBwxis0ke8QxPYsxS0rVk3MNaPnYa2cD4rWfjFxgfg5s
Z4nQQDsAIzhsPu7ecv6ztuhf7E09phDbozW46ty5aQPl6KgcQZkcjOsJGsrtgrdAKpxZ3eZjXsGq
fV2afCZrbwZKMB1kvEaDPZ3kynJUKfAwEtDCkaMvh5UduukJPewIEdzDmkUlDD4LmbOAYJ1tTjC+
+o1oXzIE8h+rb/oboBAYXEBzgEkv0Uevd0JsLymqAu/pM9F3dBsLISITduWoIGSm85REMdofNPO7
BesDiAL/os0DDWn/XNAjrJTI1NRd/ECrYZ6zMlNBBta9rheOpW5ikSSfoEkMdWFN39AUazTbTorF
TY9jHoVU9dWyA2ceB0quQQAObOEMTvSItHkduPD64Wqh2nqiuI00enxrxIImofQL7A7FZTo/2MHa
CUoGqUp87eyXiPfU76u0znWjxm423z0SGCWZ5FRbk3Z/N4PeUHv14/bpOXIfIgQXgUAaiWsLev/9
20xJrF6IhKkDaGgE5pPcuMqBoVPW3g6jnwVA15h5NZON6wVBVuwCCGS9GQUo8OOnc5vpUxr/cCLE
APQrz7pxzEH1P63/iU6Qv3CmKEf/n710XpfbTtqJK6pVrn3jDDbXJjMWi8AAJv1p9NYCBFEvfWmT
K5Ujixo7a+FjhZ9kY8Fl7Wv6DJCjPM9oPmTF/dA5TR1aL/XsuaCZkodKTHb7VMn63r/6gAHC2hQ7
xM+6WaRQzCPDPdIcpC04Aked/HY2951r1vxZeUfNk5pTTPj8zN+pPfwSPsQ3+NpK1Lq6IRwOtkBr
m+1GQ6Y+u+IsSq0lyipbqF08GSDl16i1A40j6vQgMmc748DorbKfTDO3Sx7kUrWUEbD+pXrpOtWf
54umlVojE7luP2dS2sWUiPk/ilLiLDWgdLMF8F6Mk2Sof1ptdpiXoHgsVfgvxawy7ijQT256leAV
eJMkJ3Clw90fp7OpNjgK3yM9wf5A/WTaWM5cZ3aYPE6nwxlUIiPRR5GwnpnpuS+0/bIYSF0qUc1R
TqZ8TUZwAafjLOUWdJti/Ph1RYqjI4jBNX995HtuJmVRSGQFZhHCYF0HZJVwIZsEAk42WTcLGFO3
T3enjGCJGnGOiJ/FSL3Ycn8bI0sxkqwYW0A2tWp80lPTUE85TWFrWdeFFrhwkUFJlB2Y/W/my9SA
rnyPMbH/gcU8uIl/gN/Jb+bVRNCoY8744npUrmgo1V5kBm0NYX9me9fiBEwk6SDa1+lropmYvGp1
Wt7ekbQp6+B2GKL/6srxP6AX2fgDBmA0ayEmd5yaBQVLzY9Bwv7+SUPUI0LJHxm6/59gysAMXYcA
VJUR5wnILaL7wf7K+dJRsigcMEWFg+M57HlVmTLvw/ojnOpSKm7+2Ew78mSKNfQyicMypuaYuTeh
XgJ4/2jQ/58zUWJCTH/IfJb4iaTm6dLpLnCQSWQC8UYyVQ8SpEN3c97ndxNPQe4C5S12o2LsTVsH
KACfZwhMy4SwgG59rdVqyVKSR6VrascYqtDZQDP9bXHSlaGuKcL3SmKACX7w5t8JfCi2KYjTvcqP
GDvXDkt/qaqLvT2PqcIJwYoXiw4sgsqyEwceE+M/hUi5HHM3KepJ1KyVWI6p0IT4Id5t0mL2aIdz
X2jUDL4/3cmTt1oHURA4+ISuqiErupM6cepmz6Zc1EIj+sC77cxVc+bFVIxjyDxBrWyM3RpEKOTz
oYef1R9lHXv7Scem4PG7ovpTwfJzPGmO7CAfd4k+bUyMkcjyKjuOSHBtuYS/CiCRCLokBuKl6MDu
Prd5dPIjXGTZEAzaesr1BVpalsPJ+SEg5qchnwlXu2SJe+8itGUGZbZ42GTYRewSRYZkQ34YWPCw
itrSY0TdjShOukqVbVaTHr1qMnCUACMmhPZLKsmQZsmnST12W3QuAJI73dj++9ah7NgWjD1TjZHR
CTgVJIggd4/MfwZVg4fGMiF8a3u93mBrAn2o6wgT4HMqLGeT4Wod8fnyGj/ZobUsrKUC25CCxtS1
Lgg0wpL9JleGTjdYecyNzexq/rZ+6ZRZtwnVEW0486goA07wsaGiHfERsCJDGMPktbQhXqqrTY8e
J7bY7uZPc8KwQLrFhw7niUUmJ43R8zBvJWL1uWnxLQ1ZvU/iLTHBKjayTVgnmVFFgl5t8QCKTERy
XKiyLsTUIIxVmosybAHL4pu0Xq9f/DUW5J+adr7t+uyLtTeDOAGaeQfSBFWJUDVhWxT2B5JK14vF
mWZOdl5m4bfcc+Zr+AOBKaZJOpkRctRbwRzgys8k/zHguUYMhetC7N25KrCcbiifW/UL1dCUA5mj
DEWlxUg+93gQQ5tpN0DHawjvRTrfEChtPhRhqUiN7i9k5YOlaEqWNGQuZVoNm4c6wl16lqbmpYMT
Bz0qOMPJ/TGfBgIBGSznuPS3+62O5AUDgSFGPRp6x9mLBR3gsosVPM7QAeO3dqXfMtwOwOVz0Uij
4VkZyZDPpK4x1XdjzK+msF+jo79BoEyTu2+ViIVt13VahXqvVGBUpFYaJWOtL7OKeko/xwCMdgB7
LQJP9Mu0hXLxghd6lfh22myNTokNoMQZpGnoexseEcjJKSXp2A0P4Y1APpyvM0/CrJb7aRaFfNJ+
SVQwbSF+mD45ftG0Vk2U+SynqBYmLbdXeJJzJWJb0RfGY8hlXMOUTfk6Y28gC03PX7+JZv9RzzIq
nLY0fGYN1r3UGMFpp8KKr0Bp21pEzQ1nBJvA9meSeiwJlTOJ8ZWusi9EKpgWE8eJmLsEA2j2CNbz
yf+pI1q1sCwEkAdkXj3FLpp15786D7VhrGh098QSTvPz3+o+o+R9L1HO7keWK6Bm7F8DoeDDG4Bq
yA+HQONj1jVYk5auMGW2vjGXrpkr/ap1KV7GEWumBevul3AAhmG+Mwgl14xIO+EJMR2YWGlXkBWd
PEL7fKS7a+qyucrUxHiNZ3BZ+VES8w+butO122vL10BWZmUji2x4iVno6csQyjjLgTWusstrGwNF
F5RcUsuFIOEH3OyTlXMAUdRDVmW3jvz7DOkid1H8WGt/4H+gqeIoOdokA5AwGDEyypZuaJE5mrqw
fUt/HXgOPaHG8ceTBqFyOTNKD3mWQ+mXSw40+Q7VxUmUKuOg5gDzVGgRwvKMopi3TNJfWRwqPjvp
1+3Re0buwKQgNz3jh+GhXj969ruOb/H8VH0ykhJwEW0I08SNFR8wxWee7yiJhk/C/u+eHe0Zg9SY
0ic1AnHzPK1MO5nhzSWA+WRlmBJ3P/Zrh46yB563B2gF8Y515C3LMSCpyK8zW2q/CzoA7aTGxwdf
71l6Yz0MWNm5f4/euVMGXfIV8bbetdlzOHwTsNNoUKmo6d50PRGuwWX0yVhEQiOgU7eLmXHYe5yb
/4R3jnKNSl3k/w+QUrIYc592Vz1YtEAWsEAboDYVimeSRrqmt5ZYFjG7oAxF135Doh1i8C2fiuC0
RKeAGsLW1sqsygi8xuyhcJ4N5GNUaQTLa3wxdLqO31mMXxLHKfKFttwRqSx7asoXNCeryONErU3N
pdGhvRo3FAcmULxWImc+fR+l2Lm8362+WsyiR7j7HpxXu2N8OK6P/YYfyLz9lV8ADADm3UnASTZ0
3A/aCsITNqdNjqXRwYaOll7LeWctYIUQZIcGw8svWaWkSdq/yytRVRVQdFrPrl/60qj3mXY8sm5e
CWPRwBDUWYop0kR5o/JA2aSsl0MsL/pe0mHDypbUuBcrg3GkFB9Y24BT4nRriZKdzU6njmfmx0Lp
OudfoLqzlIdeKLvm2+YwQ8dQj4KXwDqfxfBPK7PJJ/CPa5VleubaYuFaYPDFdzwi03lJWEnQ+U7l
Sr8MUhfQKp73D/jdnID/O+kZr+U6Ojpu1Ou6MiiTMryi+9C/ijGMMFQSaB6dUFF3YN0TDr/umLUr
+l/yXdQAwxizmShyMKwBzv2BR/1HmmBgjxHxk4ZTfsFytNAlQO0NcJ5OCcv2W+0P3FHdWxbhlpzq
5VVW7G20m3aFZkF48Oo69lo52M+9z0H6XzWUKqVz80+faNxUnXY+gpOS0A/j6cS4x0uDAZpC2M5l
UNQ159P7X5XhcgGGxV4Ahb5d5fx986byY1K5feMxA7ScTqxxJ+4Wol+rCc6Q/52TDvFsx2ZYKqnr
Xz2tBeY3cNQ/mcZOWfIR2poLL7zg8HySrPaUhYXJL2x3jfRxukq7m1SkrDtsL+uO0ysn1rINsKqO
6RviGq+9p173gI4QN8oIAO8C0AXBG34nx8ywyZAKs838v942X4cY5TalSyB0bitkZ+Zg+Nm8fgI+
fXfTxiaQVrxwm+BQGWPazROJZXr/C2XVQpSNfC74+8SsOoJFzAMG7j5qTpoZPV0TfO6D7ltZICSO
j8AaYCmJ8ipzPCzItdx/QjiIInzlU8E4U4s2D7QhKriQi8rRIGB2AhkjMbxc0MFfp9LRFcVGIA2u
Hr8jEdsKfnuewh2oNwwnFmpcGyoVmbXX/lcdDG9aWHbcJfF0beIneiy8MzY7i6b0XlGJiyJlstXV
ynNIr2Isfzw2n+AyfqkksIK223p3W/+2b8OBOtQw2sb++Mujpp0SewsAcXt+m9MP4GRIbhHOSMdI
a0l0dT6+tWQ1V2DAOySqkSNaryLxR9+zKIIjPOGPcumjVxBi8paO/wKs/duWNC+o6KcXbtjiDK8u
jmV3VOn/PGxps57/gRZkBj76YoYsggkw1BpCq/OVNnVfoQ7c7OZq9mm0003WiUDRAlNVCP8tarUQ
zmaoOap03TaurmXa8cm+YbG2mKm/PB0OXJP79+hE4sQ+hDKtVuLX/MWBBIcnAPYrxqXRjAA9CX4t
5+Jdo22NXZSfjIIj72sPC2AgJVGwSv7V5szFxwB8AH7AST2kARlXiAx/egcUk5D29BXXu4FFsUon
G1vDEiTe/sJqBe2QgmgifsBLNVKwr5VmCQuTHWnPEjSm4OJj/YRmdS9Zj/WQeCbhpjphxFAdptYX
ppc4Y0pP1uNZhCIZ+P93IODT3rXPp4wYHLKN4gn/vOyp8vtADZTYKwASDRVFv4t5PfZ30cqHtiCS
uJIOqmFkFqkS/OnBHfPWMFeWsi69Zh0+kIMwQF/I1g7sQWVP9GgeblpR4wGh6gNNLkSBhXDRVWPK
02+ih1YD4aMjrFCD28Q4WzeoItwIeYlrjsmq8apRQO9lxezCQEe3AJM68wDR+ywAVVmnqs6eEeQl
8FmvTVrUBwkmdiwnxP8ioHBfTAI2GaEAXvmwD+7zscqAwtxMTPzgVzQeMjnzoWjcw0Hexq9eaKc/
E0Nrhl7/EkiSuWYtZOp4S2Wp8M3HkLzrn/dpBLbhwX2okmDniTrq9fx96lJp3R9BAAe3fe0WzLv4
zhVVvwnCE6dbBKyWC/fgQhJ29IopLY46ZHy4e8me+Pc+EfEyLOvV4bXxZ1Dy2dJOWrHYx1PUBD0z
eihbTCxvtA8ZtlbK207MrpoIXh8wWQjQeBt4tjhBUGrmZG9tDMcKHO2SjnjEVxmUCEz1CY2hbkNS
/F2ZCnnBHFRRYWtJ3uP47auJTTl/jMNTbg2X2cKYbqxWi3tqgxjXC8L2r4bMfdlCHKz3jmc2CKad
cZwtxiDpg+eFABaX7JATtUZa6Uef5962upbw5KL8DtA6lrRTiLIgQZzmvI+Oo/u/L9XgXONeRaHd
0pKFHuNH+isWK4t67KjlXTCqoIWCfCIbIvO1NbFEVhyt/3fovzJ7vkR2kkfvUaHRSxc9oUHwdkQ4
x+pmWrAv7L2XpoAbZmvILxcjcnxU2kBpViARznJg1PPJRnmzhcNPxvyyuhu5/NES5zHc1GuxrKiD
qV9r76h1NK4BcAnQ03EE/VDz0kHmAOlbI22jqRB3gZfwH35Vgn5pJCFejlKhmqEm2HtT5yD7mbFj
ykHeMJjNsjx4KuCMryfGxz5VDAbVozxcwzp/K1GMraBI0LOad0ZZIvN5+YeuCiuQKScbUOhqJrf8
Zx5axxAUYC/1rwAJyMYOkvujDNn32scodnIvW9RG9Nw5Zr5HyUYWmg3giCpQEaEFPV2f/tWK+adC
VgS0Ak3dOeOExATaFfug0Cp1iz84utVNL/ZKVKPwA5obtVh1A3B4/2Dkn3b7z+wHIkeS9M4OErI1
LBgodT4RU7j+KklGhwaVJ19n5451l1PCaB7WkkXlsP54wTBtHjpB2TogNzV4R9Kgxraie77hbFrg
O4tX1kH/CDn3lVLY/HTp3NrYhB/uj9Nptm/lcz9e/oJk0B4KFXhvh6ndR6P5rX3fR3h0M9ueo8up
FxSH456+d8Ykazl2/VNyA5DFqbWvR33NBHXJDoBAiTjh2giDymoE1q4+0M/CMPaLl5P1rD0r0q/B
WSIU3idloxYvu0/RcdxIJnLNi2qyL1bvynLbUEDocoTlvndfNoUUaym5079kI/12IcwmYx+r71qe
y4rPNi2UgBdgV26xN9ba2d4WILB5AoXC9KkwV7CdMPfrQUxpLRsy1GlR78yk2QNi560HmxfsrC6E
kXG3gRhNkPxEwvedhF5X9LXQnoToAxToce0rGxKMhDj4Qlg1OyfkgeK/qnoWC40hIV8pMa70DjbL
vGgesmixWHmZRZgn/YZz8bO7rbu6WhZLzMCK9bPzrGmNrG0rnaCfBeW95rLwSH3+GYDozfaGsGPV
rbpUBC7cobMzncFqneeY4fxIheo7Dpq3twAon45uGdhOuEG9qfrzi0MUiu2Ps6trxEFVazGXBP4V
AsPyTmqy9imAUxDE14pXrJJPCEg74HG38viVGoh4ZoTK6DHSIXF7Yqm1T+wukG6R0xzdAvgQXHAP
dCIJKXRyS3KI3ZH3kJXGW3gj5UMobpAA+FekDU9OcNCejoBXRNmlMB1PogiJE+yMvppcyIyKJm6f
1oNS2c7fp5oTFDdV7YrTryPc8VjoIJSutUe4x/jTYxlPSuh6N1raF987glDkrgp4gEqfcLw2tVpg
aaxzsZai5ZVUiEKSIWXgnhAdsC19TmJ1/d7PEiDhvIWxL3ct9a6YqS0Y4uzlrFtSxtbn9zcxKhb/
sAFbeQcDSjSOMCS+q/rXb8H/ZkBjiJvot+1Nh3IQVy3XjKXmydRUWbdDD9L3EKm0K2xDpFGPSxuI
cZNWAN++63QH4NS1VbcxXi6jNKH0beg6Az7hdu+EkZ/AVr6QbiSN1CiNBBohjcc9YkkjRMVMrdNE
KV13eYQYvqK4iNlG8407FodhYZPCV2yyUSqnT1ab+qoVC+MGHKBod2wlTxE1MgGvBXbCoV2UGOys
8bzGJRdHZNNiVGWfGSjedAUQMX0wx21rHssacB9/JqvsH7ZkPcwP+4qLCSp5plsCz8ury8wEaf1f
77FMBb0Rcrlum8BfUtZXEQogRB01ivJZ2PsRPafqh7I+/RIv6nmMc9KRtGOoJ2bMdzKCF69nKj1D
KXMOP3Ugryk7L48YWV6w1nTNDVs+rbOGHtcNhZidmST5u/kNGhN8aL8pi/GZHoJCusxU35ORulhL
R2h+dYF9TEWw+s7Ogy7tm7Dbyr7e/EQeJDKiDbkdKvjOb8VTUOfJByHoDC8j+qOaCVeilMNzSPNK
q/3uecZ0+5U6Ji9wfPNRngk9DMqSjDK+CA==
`protect end_protected

