

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
AEDf93kkZknTAYDLPy4q67UmP9O18ta3jK/RtCkxR3ZqpY2KlRt7rza1H96MUf+qsK6643W9A0n0
TP4few4v7A==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
erRjv8zI0elbdGyufePGLqKRctW7EMRy4ag4V3lsqysjcz2IbkoY32VNXZB9TkYq6LxuID3xgPR/
/dbN8HKNlVJr4fTV1LqzlQYnx177n3iaEwIdtrjwP76G8DtyrbDzV/JISwzd650MMmyKJtHnC2yw
alWuAIIBdbSW+HbA0I4=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
gdHY5LRWuJLwhBPcRYPMx1NPD/GuGCtHF8ywmbYLyoAM0rjTxb8zBoSHfJbS/2vKpgG8RCdZOknj
FMJ+fOkJbpOMFaFsosZ9XfIryZEhroI0pt0zugw4Ha2XsmQGqxGDd3IyGRBNvDMKRw2cnjSZz2Oy
H3SrajtWuLhpP/vuSzlhtnqryvgbp0USaL81fja6LLlPm2jXTcuqgEPsJwwUUhxjUSQyRtABTEvs
3Vjc63pIVZUYkpkoaKpA4243dOoRhazlhTF1c2Dp3uyCrdGZU4fWhJHW7m3Cq9Aw1murzYGrPLS4
eQrf4MTXbiMtIPpNK49OUBbEpUuLfnDwfATFaA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
fCQs5S/zt//IgxsFc+FuMl79LHVh3Px9B+S0yADLC6MfIDCRddIdSKbTMZ5DlFrngWDJwpd1JzqP
cRXcul8iGoVMrVmrEStKWXi/mhtK5UkWTAd7hoyj5zcI+N7wWWxU1eBAeKZQ7uML2SLN8mYzQYLY
98ufqGLyMQeFAWp64iY=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
rLzkYB2xv7C/3jKaA9rJ0Hz1NLTW5YORm+QksBhLo7WkyUXUd0Olk6yTtcSIC82lRfBo8f3njqY3
dhmWfikGbTNV7gixnGfPYVUvZg+xsJ7adfqwnApC/cK5eBJGeWXZ3Z5gEbLOhuRw/04o37fRIoCo
Rt8ZH/C+LE5As0rIpYw6uzjL55RYR91wP1R/rUwMQTNJ8XwXPkAbkuyw7FWG3uW7vEvZ/CGu+T1f
VDCUznG/Mry2818W/OOR+t5yQ5fYiXNh34gzkO30FRWgtIR7ZfOn/fgLqv2Iaq5XPzTdULGOHjv5
Pl+0fdEaYyo+sJ1yt8Il53T+ZdgLTjEgv9cjPg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 30320)
`protect data_block
CgQlefeY02q4f9sEBl015Xr1i9WNkJ6A7wBookLiXTcg6mmllu3VmBdVIUSBcupUp4ueF9OHac34
VAbu6esAo5qQSzH0HcS1nDNfATfQDhWcghUeYjNWDZJ2nzXQhZ1/ShvTkgwYUct8Ct+oLDOzsRl8
MZgZyj1kziPvcp1YwGhVhkwLGQ0O5QD/hD8knnRwGL7gUX7W0vVH44Oja2hcDge6L9029lvhIacJ
lD7taclXmQ8u7CVBWx8XP0gjN3VdMV4ngFJ4j95WcApz5d4Zc7YNMvNbaTgfE64N+jDtbNr8sWTz
YaeYbbQOZ4MdDTyAkvE35IH+MyTweSuB+3yUg2bBNb2gal5RyJ43w4dHc9ajAfYsoWG6wQNKgqTW
qS9udTmv753LWlykJLMCeJ8P3TSDsLGroxAJsB4N0ErSV4M7vKTzth6UTdOpusC+VinWKXstWE9j
xegCnoeGMFWaFs93umvN2+zYpW4ofiocv4Ot7V2AcRzIP+IxpD7q4RF1NLJglkBmcC+hbj1UN7Yo
HJ6fFkqaB0Sd/GsmhBDNFpsbEC7lQY80+BpER9ZkzpNMiqtLTC8PGzIgSdwbUeyZI3FZXXOWpSRu
kNRbc6n2j8QEb6FswMqhXqdcoaVFHohT6JnQngWE8p716givCzfBdKYzlgi0WQfJk0pybyUwRuik
f6Nq8MtG5mIA5ZTpYmb5GTdC2x2+ly9msWPeFY1zwGh87uA1tOhE6lfDbcGE/vsQWELPo2f0KHsy
NOBzNg5BgS3t37rsdR6O443rSNark/XA+9qal+u3VLk6+Du/OVxN/zfBCVrHoPHwgrEr7IEt3bsF
aNtHbCuFkyk9jWDDr2p+AO50s8i6e2QZCXWQ19+GDf7JAQBtkdf2Gt13d+Kkk0lA0P963Y3SKX8F
HlW7cca9CuBe/YzJCfOOqOQLSCzjuZBhQE80RX+W9lHPLA6PEy5yS/mCNKHOvC2PLEQvvLr6dOwx
vMvjPI2cx51CkDaFH20p9gPUHhRyXLl6p2YDRHvk1FsqbJJR6bQiFBrPVHNgKgtMR4FyBdXQUbLJ
y5F+jdrd6rROpiW8UA/O1lBX7Szoxnec7mOMP2wvurH0L6fRzSx7qVoiqtQhq8YUQJz+ZnaZy/QC
0LqrYviWqJSyLSP+yivYhJzvGVlKwEpXEFp4zOca9j9AM/8S67G/kGXFAtvtF5cz8j/A0UD9Fcrs
KCJm2DbCrml9/wEW0Z51Luw7XTbsk0dhz6VMwZaPqt6i9gljXA78izbU6pWGeW3XNAG5RtZbVHE5
iT630u2wC6cipjgakuPunlXtPvWS1Vtla8QzBEe0wMHQ0tlpUa9hqv1v0a1Jv3YUjuxMphFf7nb1
A1WP1aiApYocqRKOqAVBajKRIuU1f2Z0NsPUC4qPF1U48JS2wO3x0KVxPDltfC/DVhmuVIGcjBQy
8fyby1AnO8qqBRXOsdJasv1Jv6skSjeppTWx1lAPRAW5UHXNAIIXIvpFy7BAqXDgN3jIg0060NOR
v1OPqsF6fhtRSpHN0Q1n7ByNC0ah4cTHXLkjZ00PsN9aS+5wJ/wKc+ziL05fwjXC51CTg0K1qRKP
PCzR8BuQU4VrUJtWRYL0izynJlVEPkE9Jw1na+SQ0tSqksarXHSrzrS3czFwLOIqM+m3RNhyGTz6
/3hv575kIvVL1JFg7Axr6ws1IWSdn4DWM3R5F9SwPAM2444pu16/mzMn2QO6YpPeBTBiL/SVnSkN
IXdt/Cx2CiZCbrBtDPutzbDTIU3NZpKeH4zq9Upd7sB5A+C4vXhtisTSbUFlyw9oQfbHUoop5fdj
LAlej3RBojnl5FE2Wpi+rh7gDV63sTmWrRWNtdKG6pR2aEooMrGK2vzbSP4L1BoCouifyjWV1Tdr
4yESoRaBTVWe/XSkA/TQjxPzj9u+zG1a5rgkEAqF9Np6L04EPNzGpryqkfjp1dA4m9SY3txiTOXh
foRZKhxLoyZMzDpB2s6gl/ugCLAO63Gpd0INhgWbOgnAq7Iw3ECjV8QXTpjY4hUAnty5amS7s49M
qDGAP3UbXwKL+rdNoOfRtu9jJvRjvcwZGMqGai0+oFuFGII6bzPrVL6r0bbgvxCE/K3yAWn0Q/jz
v7hsXwWL/T+CpcDFY1rHvhVDg3Heg/o3rusPxHYM/QeFbtMCRTWM7icj3GD4VImCXi0thTUVOe+m
SaN0CiTti8+bX/JqpD+P8qNKJxK9kfl8vg2u4cdI/6Phdq/eQvtNVnUSyea0UKheKhT+4jcDIyaD
fzlqlafX2UC0T7RVUv4NzlRLFue/86bfGX3wnIYUokth0n8/OUpQq7xB+847hRlNgBprsQXXKGxJ
Ac++Hc/esXCb/vh0o2j1Tu5xJpJ5macRdnv5wXQW/Cf7LmgQMN8BrSKMHklUDMIzNmCdO0Kt0zbt
AquBH7CBQwJwDxAVCF2AE4xfotXln4FCbol+JU/9VOH/PYUfd5glglYzk85H9eVID4lp1rctUFZv
oadmJ79wMQ65XIaZF6M5NQDzijUGjFvch2DJtDzTZ9FPNA3dVccheKpohTASA+6Kxq2BZZNUSlQv
tW4dF28BbHsmIEtMcIzr5WB2b0C7Ehjfh68i7QdJLlcCh/DxHSl5enqcomeIZcApnzLS7XsW3Lza
a48qBEGrONGRlbijP8hlz04zDkFiMAA1LN68EXqs2HyWljBQrMuLn7VmhmJh5mQ7XOfA198e0kuU
nd8g36H/AycC4g9B1lS/AlgqHSPSqYAebSTcXeUjfAT8FRyzsf3O+SfNgo1DDapAX/mLBmw2siAw
soZIdW3furzQK4AZlIT0SE72hsLUIXhK313F5PzEUpjES4Qflxr8cmvi+3UMu1y77RDe1uW29/Dx
ksN+WSdmTkVr3dtZkD+uBwGCd6mHcjvmUrsO7ta/0esWA54NW7a0yvKZ2NGrANKTmhW8BuOqw3QM
eBpMGzmRmJNBD4u2q0wGmRii97uxfODoMJ/1adCQCdHsXSypIhTGFrleXszhVwRpPq+kFu6E+V94
qiS3nJnDr3/cpBMhwnTqj+TVdT6YoCWixoofMonX1N70uCDs0IyWtwftGmYIsJ3NEGi/HGcZfAsg
ZILFGTthhF7b9mcV3g72BJMaEOdHaqvLxDXZW+wBZ9hfd+5E4m2vqVLexnl+/swBhFGOtDqk7yDs
583/5etXshX+BZoglVM1OfdENNuTqOemNSUolSx5gJeB5/nEYvryFe4XOL2H1gthUffGyiFdSIol
Q4z8mh6JX7XMdzrsjfWuZA1xMfjSX2DfSpMYAr4xNH4FtSpn7QdOBdQMci9ThAqAn93keTx7t+nH
9R6bqzcgsFTgCV/ZcuYZzEyR2LI2js8VZUJ8QoC1aGZuXlwrGJst+CptzDRLQwcU+6QBMMT/FZkw
qMOmRodaz5/xdNyx1IQJQlWeouZhIhBX8ajGjPaVQJTAt7t2XL6I7M/JjL49Asv4AEvVe6u8hbn7
3oRvaHjmFvMHtvEWwlWWpU2Lw1fT2W1m7iHUTnLbQZkijMDbwpfLfYZtkOjHPIWNyrOdr2jHJAHS
HGPAmXYIu52TtRW2iMz1VI5Z3oOU3fvO6phWTrU4WXV5hAfgunAE+vA3w2gSnvZrnyTIk1NJKJVD
djs7vw2+OHGY7wzp2Xfdmz+FKHEpYMi9u4gWj72riW3cHEcfCQm/opzy8m43tdlRlXxYhpVidJrp
OIDdQEYQEz4oEVQLDAZFeudMHorORFrsmZ5RphMrWCC/485v67Gw/Pz2LnqG/raohNn/Bz2+Hqq3
QePSuALSonVwy+LiUM3SVzjYHMETUD50sqHU3IjdpoTdsgUwawMo3XJMDnw09s+/jX2JN2Bi6O95
jtdc2k95lPqaHjBuvkfHgZOnVqGNUTya4symbemmMtddf+N3j/KsERhRgh2QUgNu/beGZtpY9DaE
0NLzrnGhD86x3fSKquZv+N4jNYjJGqPnLQ1EK8KfYNLzkX1R6WqT6eqzONfLEGX33BCjN66xn09b
tsFYvPEA8qKNM8zHUmGzcwxOhNJE1N/I4aIAfP0r4njOdBL/BM2QASyqs6svIciC4+8Vnbs5OB3h
q7GqWKo+778zQllp+8SYt+TC+7S9agndm7e/eYdsq+rU1vfroAR5dMQCMUzyhnTqBoK06qlMnCdS
bxXadXpByyzoFVBD1yOtI/DNy5Wwa9ZVi3y2JalaNsRLDaxzWIjzvh6cpwg4p7tmFTTwYXkBISoT
gHhF/bwOq9uG3Ff80luyJC6diHB7Nsv5jnligb+vHtWYNbz+AEIDxhddmCVu1r6AebcBiNsbACYU
XcbCaTXXUpWyW6sSMhQQGqswM9ya5tq2pdKQcKybc05KdGfxf/LM/6K05zpIj3o8vQRaNX2taWi1
WNtVHejp5WE2pHEZPMSFVPb/5uqr/UUwc/jgd6np8Yvj4r+fU8MLwAJ9h7HVcWuI31peWAbXRCXw
8svYZ+jYqlLQb8L6IRzZjYev7zptOfMUFtMd5J3ZLXeoAD/6nS8TXVwKIAvTSaGM2P1zsHJ3+Qih
FGliHeg70PfNp25GJNBZhg1xDJsLEGWE8dH3Kzasleyz1TKnonD0Dk3gmfN72s9vJ0bbhcwzYkji
H51xkASHk/yigb1zBRNSs8CKeRzn4hHQGMXmSazRc8WJN5R36htXURaiqqmdvpBX28iV8RpYgPb5
RwdRwiY/JZ3S0yBrmBwOfHx3CwdtlQdKqHKaPwad87G6gzvQcCGXQ46BbD1lew8z/XxQF+WHjoAZ
TQ1JhW17k1YfdxWXne2ACdgoCQtiwlX1rZHnLGpHcT9YpFFz35gqzHDeImWhzXU03R9cyWqdGhp5
EHDk9d3nOmPN77bBRnDF/UP7xb8mg7n/aV3TMD99rtD1Ri1iP4uvzEbrpPwgKxzEeZcRVby97wRS
07SijSMh5kHjyXtz5K6/7xGmATwohgQZJyQRMfHWp7CLWoJpnV5oWMVDgPRx7i5jud2i7owXfI0h
CunIEzsJmTmc9G0nN/byh+GuysZzv3uWRQlT9XWWJ8mC+zv2XTMSkHqeL6SkowD4um8SX8giS6yu
bi18Bc1mFBFxLUW3jj+SbGveIROouzO8kPyVU/Gc/fVFwO3PrZaxwrdftjXVSU98rn47ngPhEv+P
H1Su408BjwY8XmXIejkfXgjcdg95oSeBqfykVul0nIv2tY0qk8SzJb+wI6DbF5lASRkVUVJi81zm
WmakSozjLwGWggpR2076lYKC4zj93JQ2DiAk6XsCX1U+Xsqcan8imrvK44vRGkdeQayuM2+kQFUZ
ZsLS/B90J+ec5U+JUHTjXXV0+fONRrg7uIc9YdAy7PguLXYG+0lE2BwE0Nl1nqeK/lpSsEMfddfZ
WmnB+dO2+I2u1WJvTRE0VDsL5GEhDxv9vyiXyfi4TsMp7X4GLQqhPDvzLxjl+Xg9T02O2y+uEdS1
kzi9MNIIb2P/XfRBOu1Hivl4lO9XwQQpbAduIsTtxQ794QEao01uM2zVKsR1Z7HCdAitvsQyDly2
t7yCBf/ATYwjq85Svx0OVC7bEt1ddaSMI3C4GQK6VLp3F9As5eVGeuiXMfAIQYq/OSQP+ZHq1JEP
x/h2sfz5CsE3lMTUj5WjeA4GhqWu0EC5JPHDKDHny6UwVrAV2KtneuG7W+T0an76IKIwa2YrYNO8
0YkK8ONNiZG2SaiKjJL7f2GQNzPQ/sOgT4TrXTu5Y7YnE5s87axOROrDZyIPdf2e9j+8j0E9uT0R
kqfnsaPsP7vSE79Lsj3rqzxehqkT6e4JTp6iARi00DgosNv1Im8pL1oZy/JoEk6B/1yupJx8ie7q
VHNwwcsP8aR5E4QXLn+hFSWzWxcKD7pd8Gr1ig0IYm/lBH4lmdD7eZ66reVToVPbOfB2NmEtGtjJ
c+V9fN63HmOkKpCZfNXKzhgEI70E9oyIzYmfRH+IFHkqzZO30dgSW0IWJdRtiSMnwENHbBbdrqUp
P5lb6DFDlUqO3dL2pORWkuF9UcUeSQpdmkvimfBzKbXdcij344ofcTUyBls3XMaN+Sns0S6oEkYP
aIQobyWRN8ZMoNq5VjKw4OzgWud+VJMR0JPFaQ1bM6MTXgKrmiKIs3mmX5DTzNgHVy97Qimy9mJs
ZwOK+n1/tZiJXmuMyrmm5H522wm1VGT/YWrF7Sn/aOJWowx9Hadun9iBaa4M5s7i5o1ChV45whSx
UHZU0gElqzesw1jMJvVvPzmQSeUeuqKps39gAs3howZvaYcmHuS/ohqi1goMUEzY+se0yGBPnE77
eGo3P1tsiJEbBNnhcjWmqVIZfjh/3KiW8KN9vH8ymgjTyB92ScMFV2fFuJ3gDb+oo96gb4Wv5mdL
WySp8f0K4/BRLFBOoavtb2rDqIQMdnZnP/2QDwN1SXkHGVi6WJx+4gUj5UdLWy0X9J9tOU2cBXkD
6RSYY5lywrWkDFsFL8EseqbNOkbh1D/NLPaosThXKNlBhNVv4EYaiX1Aph2qbHyGwxsw0nUIlEXx
ajwdZyzBfLZyCBx5y/OJgEsE4OLR/7iTmEAoXJV30/HoAS8pwZBci1ldigzk0LopJRh4+9fPqjZm
cxzFOFcZUTn3FaGMy81TAaowww4zwJu5Fe6T+Kke21Fpg7nhHrKPqw7d/b5HkO0kXMWGfULAQd3C
5jgt1X8SWEKjBOiaVTfH3OQoKvM2ukx/nERl0MCWGTsQUfIEHO3BfJY4y6oZrPuqG0EZU1XMGrTB
We1Rm3+xZ9iYRItrw74y80zEpea5d+tZ5wmC+evB8mdgr7mz5YA/FUAIfBYx2P3uiuxgQN6UYTFH
J7J6CvXWSyxvszYdpknlxC8vR7cPv4WCqpVEP6Vqz5mb7yMo4mXeWpd4xLP/bVkmykRj3feAvVnv
X3yTmdoOwtO+F8heZjEkGu5wl7xN2S/2Xlu5pMLkcuo9eD1vyu3D65bgejGRtYgvq1xfE7JGlXPw
KBSAdLz5D5csvAkNqiLGHctCitSMbweh/J6ibNndq666D+w7rKs4cbpULUNDDxPM8IHN5Wj0d+xM
MSiUim9hcOupNdAyqYKpYqIGR0fOSLu+T33/ycGQnTXrV/CHlO8vJZhI01Vvw7FKvC4moyATqKSB
VTpN6gix8yXN6CKD/9aJZCQekvyXifeG1VkrfDshD3jdnzsqlvKlINBEbR/412Z3K9UV6Lh20NwA
5oHkLdAn5CT1JwwckxLmbyAYUkYIGXXdAOXf838zz8Y1CmsYSEpotTpzwSgLn1bot5/SSQbbvF7d
CV76nCW8/a4XH6ysNfJ720YSinxDFCtyinEZhf+UzfApuPRluTOCIYE9WS1zieKezbID+zKnWZKu
x+3P4bmvfoZQy9kBCk56v6VQsQHdcMQXmg8//n7HfnXEMznCMJhhB518XDoXxXZpf1Oo0jGNZr/e
hoSR3sNgk7hOGl8zE8BIDnV+bPOWFvX1kk7CdI1KQQWzSJd8VlXN6GZ4m/JxQTU6/numr2TcAYUU
ZdLYgKFQ0XOkHqgWWHmDVPbJDak1/h4+IWf4kPHe8C9ly7fBA++ROLSj1TZ0XRyjDnA821IIbCZB
UUFADHnm4xiGB6fWeNjraSER30xA4cpx0f+z8hiPDjL0D7/EmaHZxtMA9dykQpkI1jr2CQIq91/n
Dkv2Bm0n2leotXZ+nXrXPaGdqSndrjbrDaIDWMcuva4KVcPVtZ0dPwPRLHLLGkmOLc6s+c0MRmlC
dPb2TUBjl5FkVT5+E0A/ZSvfZxXmYrPqLR1Q6PPH/44ds7oCVRu21BwUx+xDTRlXowtHh20TAbFO
ua8QDEY599vz4STvD9hunoKXOFPNGKPeeN3VhJ/uA/lFWO/ZySpt7NcY2Lno67Dbi9n1Ia0EA+Pl
TcGxnLZU03wAGPQ2mJTavcrTAqDrTSJe4yDwvoxZc2P4oqaGnXBjuqBbf7oNqBY/NzZW/BHWi75H
KYlTsU+RJxdy7Y+/ffoVqbwbu+hRHyfvrpg1rGdsmaXGeeo1sA9s8iG6nknYfaqrNcjjS0NY7gID
Rqez49v43EdjRvV45fLs9ORAIhK/9XhbQcWGKEu7oncb66VKJQ94VUcNID8vTp6ch8ftTwrYBMoU
iUmF/fvnte33i05BlO+osJDuyNWNze784DURqCJk1s4fvomFvuZYHUjooE7COHKyr/sZDUWGNLhr
uJpP6aIuiI6tlONO54uEjk6VRkCNu+1tjnNg3O3kXFz1JLnq0h8/SC3HO8yYTiumRdzGdSNmtvCC
9JT7IKuMZ1jqbs+nFgwAjaa8f2Yeb9IyPpw7WWQKhmBkePlA82kxguEKcxlhLp9/mJFDHmjZZVDQ
TH7tOKIS0dlkGEhD6+Ef1CmTM4Yb2Xgw0uYl12OgFknntm9DFs0dYS9Xcpq/10PgA2EsAQufRryz
qlq12vI8ZeNr2guFfpEc37+MYs6U1y5vRzVm4iqXdL7LzesZLLBIhwtTlJcU+asV3yY7NkUanXhV
dfQiulJ/N6QLh72HoWPLOVZ57RS42PnNZptbOzuz7ZvfRAR1rO+Rm1UfhA/ZpzwYw6L355HOrRd5
3Ci0BqDaDw7Y/3r9AZZz4lvypSOG8cuWpQceou2gmwpXSR110gopCMdGtBPQdhyyHsrimFJtr3Xc
gwdNc1QnjM1E/l9t9SvQb95TGQ7NP5FDv5c0E1g5ld0+dEBtbMWAUS8NIbRLEGEx0bWHx3wiupe7
UsRjmUfWk6RrD2qDBQJgciWjSDa+9m40ksUmNQfUD7PK0ynPwOO+x9Qwn6aSylySsvog6MKCRIH0
eAmeQmavIKFtlFwckvdOkjgSiIzQsEZSKBRBuHqEdAyu+g5wFKvTd2pS/X7PCDwvsal4FLgYBzBd
ywvxkMiI8PqUH+Dg+dvAXcURZ+aCDAS9Jq2R1J6Ov5GdGBNVXpS7wMOoX1MA032oHS1ugSPeJGDq
3mVpXpgEczg/AWpeEXF2SJYtZoYy7E8lXrDLdL3Els9QueVJ5MnLUHdo8O1o/eOwUIJoTuPdIRsj
lAeDLIdCDFelLnqTpWA5BaOL3c8gwmtFkWZ93Z4crmPMCB1BjOZZ9tDaeKb6Uo5jvvFfVkP919zp
nDpl6KVLoYCLibF5aIJn7yqkeA1rBn0CuqL8hPU/Lr5bUdT4AgMWQwzLtLvQ8L7YqVFr3hOOCZpE
UYKL6iBmwDozMXWg4/LtUzX7gNu23vbk9aCdLvhynmRyOhPXSiv5Y+33XWAXkRe0nnC3e7jkRplK
i9Tg0dcWypkfPiM4GFy+3qltT39YHm+kQekgnMZNM1d/157a2QuWyM5NX5EVwR4KlpYuQ1yFn/Ft
NN0xNIWfq0RYKPB0GhdUZSuh4ca9PiAEL16eb+apwVjj3fpOaNnGczEObTEVD4NUPEsSiEenFafV
nwurlhAaZ8AioIFoMiejAfFzlo/HfgAb1GCBlcmo/0cRY46FErB722OYWhiXM7SUhasZbo1BF29J
qAhNr+Ab7VYIIY3aobq9Wu7nSsZVLxqYv/oWoyZSCIO2RXAb7eTigvbWjdbp3T0aNq8jzIwIzGfQ
hVSfaMhcxfGPUU4EzdomTQMUBzkQmfoW0zLxoQncPWYicNYFDLKugoQ0YA/geF9e4Dkczdqo2Oqi
hLP5msJ01BwiVMO1apB/4IPO9tUf+dp+jCNMCqWO87R5UeevdskRSdfCF7Brm0PgDvSZD8iK4Ebe
x6ECi34QY44IignhK0fotnxMuRXgslLEk4Y4YMvGSRiUpIijkY7rCsKjNzGbKWchrlidITgsnDwT
QqwHG3pGlMkzCIO1Iua7VdpVr4uvvRhf7Rrj1HW9ONHf02nI9XZzPIL64mI6BbFVHvvSLhMCwyHp
U5mfgEBIU7AGWeRSGmQ1hylRpvmKKdC7xLRgcvLfcP0MLitAeDmoPKcOr70SPdWKiXSiEvNTwlKD
x85sed8aBhvSgGt9H1Kdal3ksbs7ve2Q1OvYnUCk8v5l7HtqiuVkv+zun9zJlsQWYUh6bVJJuWjC
jxaMk5MI5OjLAFVjNK6mfcJa6O8qGK2DuBD6GuNYIQkI5rz3cCQg544bsDg+qpjj3GV/W268D0PT
xRUe4StQuOstuQ5Y1iuyKAycbsOLsAQlcqp/l05ai4nY397DzLeDcD43we5om89RRsMz2XmwweKT
O0O8RZOdyu4pkUaqPurmjmWatEr12i9pskwP9kwRw3UJBOolBAaD8CDuuK8hJxEjaya1s0kYd2xQ
bJfsyzGlr689IVSfOfS+sIs3fMKkq67HHxzt9vFbJ2YMMffVPjnCthc7tEZpiH5fv5XfW89dMFmM
ZXYfnfxcu1oNHQ/pnaWK8dboAdqlzbX4STT4cb455NY8i8qEbXVGXa13QPB9bhcuAyKIcP7kr3+G
SIw8F6qt4eaZL3mJIAi2KsMf7BkJGLI7W0gBi5ZiKk5u5Ho2obohwd0gi6du/lqNL7ihse3odtkM
I9FuBvrf01WhrfV91WlIKGn/TJuzY0y0NHiBCEpnfTpebztle3FukWMz8S9gJ9YYlBRyxKum642/
OGSxSr3f86oZjXfdUfJBQpZOeNpSZTEvdU08mSHaUyeQdmMHhC/ozUw2RVq1ai+QCamxbBLJVB9q
zK2Sq5Q1RsE2cL6xZSCbR1S/hm5SlXdkI06JIcdnDo2e/Y1kXS1HZHN5vLJwXDyl2MB0J48X6hI5
+I2GT7eJ35lnJoJBQPQrMa54d8b7uwyWEoEzi4ox5veztF6xfIqlR4ewUS+g9RsjVPKEvKh+oRBJ
5iTswS21dnS4+DxOdIYwYHFrM0t58lj0bRk7vzJWb1Dk5CtBc85BiSrZWNCGnxvNevF46QjbC2H8
sPXDPfFlG67yE+t3aak0ebWumz6zyU+t8A4m8I6bm2ziLyx+BqABgzeb88Zk3jQo8sEeXIBftHUO
U0Jy4EHvEihEwFstOphotDnn8dxL5OrsAw3O6PviZ5K8666EiDaIYf7dMX4svRz2h8f8nGZy5qN7
fVjd8pVavf4ioRzwWGCC3AkL27sv/E2E0R+mF2lG5YuvApc0FqGeqbkcwM1obGJOkLlrlSUCk2OV
rjwkCn7qxS2Ooqis5rt+D+lo5AhFBgaZFh08qV1shrZMPWsxTMku0iDGPUvCKWyLlceCj+9LsGkn
quQcG8dEQr2pUr/AZk4D+bRAvB4LZAK1P4DgG0Mo0+qYpHbP1JjihjHrEGZSUbCfWmAx2eeiQTii
h4w7uTimW+v/gUQk7bfLb2GSfLiKO7SVlBPpkv2YAyVxCsGhfOQmEKuKOiYBne7aHUw/BTJINRmc
vMCEgorNhZJoYitYjJj3Q8x3mkDFieWNoluJQToKfL4GuVWUY+L18wJV4yw6FQXW9ilx9qIpwzqV
Z7zPHwXBow534s6voxlDhEpBSP9EKOoAET4a34SZ/3Ar7H/+tHaSssFLgB85A6o4Ej1dMYac9y/o
g4G32Jk3PShQroCLGMEI1oZfjAHO/2WpdSZFIGzPbf0/GymwzDKm7MV4eyJGei6fsZVgzd+Xtg7H
onXAdPNHf+PfFZDF87jHSmPCsIa5UQnxJJuXTwWEbnGbXKLr1rgSIcpDOPBaDp1e0w5pmWNBqUIv
l4YHiQSPQRXnr8tAH1vqblTuChye+p8KmSJaxBEG6IE7PVzJmFQxV0h8SxmFxrUFKHXOXLnOoOcb
+BroT58npq3+BcaIXlkbYLW+fqvqQDcNGKJWUNd3nVuP/HtvARbe+IGFZ/feY0ybbgjY5ynp8feP
JedAgI5aeY2bHFC5cZbqkxQCaOGIRtQYz7YjB3s1zF6farBX7KPfpPQNzXeEsSaMGllvVZfGGAOQ
RnYpZQk4lRKwqsiMRZhEpKsoe/ZAbjuTXS2smxBdD3MPj2pS4eAwMBj2A/bAFZLlxUitNrWRzlVN
imzGZ07QHtjgL252V/CBFob3c1Zd3LzgnQXTJEcyT7wHxiYNytOrVv61jKvEcj52m6avRIORt7kK
49wHD1nBF5fW9Hnz21za78FKXK5tQISJHJjEUlde9mk/Rn2MrthTD1Zrige6IOXnnUjUMMXuAud5
fV9N4gKNXJacuqFjJJbPC8gLX0LpGiivUYejcJXyHB/hl6Gp9XyemIhhdNKOxMAB+LL51gLk/OkZ
VHkn8uGFKbeyUACU8mpOD2rhGYDyYILlwdYNNQEWwyGK2Yg27GyCBAS3sV5PRT+57uwTjop1oOwX
6nsbABNsEeYZENGmAImVTRkzudz92Vjl1CqzgfioAqZgqXq/WUb7SFrTYnaSVUJiXkGwKmHNqsmd
2epFzVc3OjWW44JfscW4nNavM9P/O2INovJDqPIJ3e5JW7nK67r9imfC6U6ZXemtsGZRkShxqT2l
2+JEqmCUuJGUOSBCBAahfj3im0431oZLPawt4ay2a9NHq/ONVcWb5BOGsI79PteV5oojerSjiCzj
Y83Jp90AJPZCPjMeqvWZiD8kbSpnCaAjCxhYWOQ0acWbzvnPDZRixnP4LEUgFn+4vw6pPIbbmARO
C2WxafItApkM1xw4hXxAx9siqXx8xmfJhG6QGmH9lgrDYX3nLBB7NX8s/i/GxYYkEmIKzHLyjXJ7
3M7ky4GQT+tqlxGVujMm6+M1EzkcviKZOPiAHmdrjEeO+RfFg6Je/gviQkR5YoqREYzqBOt/KCku
1+xyT9xVK/RhY0goRGKP0YFZUP4i5w70SXITqe/Cz5itlRMs0pfmUGfBnmQ1RyLwfGGjLTXcJ6pK
m1CYwQSqjFLRg4Sy6zh9d8/D5MO69GBING4AF+fBpff8QRpUDIViUB5nAZp2mG8PTJwABYbkeUO5
CRG8kjaTNpiacnoUc6T8/rrPolF177W6XrfIUyBcSJZcVpBbfkGt6fuo1EpKzCyDbZYPuChZCnXs
56dZ6nfH9T2wegfP7nMjQYmqc/a/gWoCpnfkyOHd5yqUwR0DJL9vBdSfm/vWi3J97zT8/A8E3H48
TKrUm5H6d0WxcvzI1JKwKBr0zGC5OOE4SUv8BkXuRq7zIzTntoIveX+MfgcgLZRRGVA2NPce5bQN
VumwBQ69o4ETzLcItD+rMQhPwawtqf1LaoxL1sIWLKlUAflFMCSkuRSK0bg51FfljmhrNLEozdIH
UcQP8RNKUcQ4oUsIp7pS0oXccto3hOmvD9iG3G934Nal8tkcd+rJmIwokEc+t5CV35cIgpgyopje
qCZpmypZ5uz/U4gFC+EscSYRrNIv7nPOVS+yPobar4v12jeCyhh6q5S6BeBHQ1uugZnNmsPhKYvV
PbosU77eQJ7GDt8DDvfQSN7VeEBfuFqGGdvIV5noLfyKj3rLGkN092lrSNUuYn7VeZFtWEwYX5/C
4VaLsNRTFrknsRHLxF8mDtTqQdTUriImCM1bCMyZOt7dvMI1qSnUctxdmxloTSxVwYzmx8Bz0xd4
CXCw8rnrFzPFIORrNZ+9Un4PEI684z3CmZ4i6H4R5qyoQh517Ja5kiQpFfBJtHAmiQjXbGHJMNOJ
+3mHOo4StAWtARzZTSKgg4YifVl6SLTqpraTl7B1tl1yvWufZ86oYxiVPHkM0iS6yi6UrdSI94vP
KqR59KRqEbpzQQDykOx5cPzzmTQPKnQS7GeeQhckxbtXEVMmAx1VzGNTVPcBraAmSzCia7OHNVj2
P8CKqczco6MTgOAtgb0TZ+PQjiT+6mwTv6QAfdqewMS3la+1RRPTcr0IDnqdHMBmBG0botcWgP5v
23Dqg//ihXraKwb7jW+rFVfzoTEyboLX24e2NmZRfVFyex5MlXZwxfxK2RgBRaf6vPTC1bv0ZbEn
tLBo8C/T5eXhwXW67r61yNr+NwmUKLC4MaGgWruanIk0PzfHwfOA+onfFVXzFYiOWeWAOLAWqIEe
f6x/pt2SKw2E6ptAexOkvSME53VoW3rZKJYZQ/7HIH6ZIg4IgoNRb9ikLttSuX0zbySVoIVtX35A
HWQU5JfENRDQYVckujhO8/D0zVlJN+tJLwm7KCUNyAXIAm7KG3IY8whQmunXrHQrEb5mvQex0Utl
sYRFF5efgkhN6JX4BaKhTM/lnhpn+iNr8W9TNIV5EhZNOhujmDrQ/sDeSmUiogwcdL+/fNt28rKz
RFUqoj1wX6l72TNi15L0yScFG67bA6JCBS7lGEMBEoa0XtoO3mglHKha+elCNVT1JVwwJ2z07hyx
xy6aTV61qZSLNIJhFJ9UpOm/aUGntdzIZb1VRquVbdvWXZjUAu+G2FIQ2tBV5Sj6ZF9cenMnfM33
dHaREI1ONzCqjFscI+kK37TZMbgexkX3H8NCZKMtQoTRfLf4s+EX7g8HEh/5E6//8KnkYcf8W3va
dYr8dldUnmYGjqbvVWrOyStBFuixLM4lcT+DnCjUoK9n8U4ENRq6UvZMIbfb0MczjUxtMoy0AotF
Y2HuD6y5pb8PQ84um2+rX0XwGU47tw8pK6Wgur2Bwpo2OgpK4F0NDAtWIB7X1m2gL+VpqdBmkHyV
DPodNjG0soAwPGblQrHtoMacDQEyO/ye95chg3Yk+dpzvNQTkcWcbDmBzDCU/9dGJXlmroc9kmjc
sYvwuQEz2HCwPKUoVm/Zq7/MsdU2GMBjJ+nqCoQfXp1IGXnRIRlOztDiOsq2XgUlNauT4o6BqCr6
A/TLcrbyDqKIhBuXjS2rWqhL2uU7nBKdHTvY61Hhn1UT80qT+QQykN7hdA9bKJsj3RMI/5yHd+nj
3ZTVOFSD3Wohu8CNaCwgeyJhoS/tFHYzho/TT4KqIvg04scXxJtHh7gOIa+so+hjqrkQyDzRAFsP
QQTxAcBLInXOcLte3iRuK/uXZzhk1knz42T1z/nvduRZmADMumbHeFEMDmOgctTi4tQReZSKKawb
sdS+Aao49rIA9Qbly1tkIZLffiw/8qnJYPTuwxJkZKjGd0YtWxr4OfF/YMVq6b90yuIlUKxQfxTo
2vo6DqZEKTPJEiyEQRUupW2c415XIEJ/2qhD4rZur85oFwPks+Z+Eb6RomiFeWyxqbewNFgsXwnE
qtBjM+tixmx8N3jNPNZF1A7yrK43XKUfaG6QzJSSUCDuhZLZl/iee7iRFb8gT8qpAzAL9fHbeIxp
7DeMHX/LpKrt3bKxcjTvdq7xFJtuISgoyU6nu8Rcv3PRGaOWYM5YJ9Ysrl4VGpnamDj+GKpzHs99
XT/7IPQtybCIxPp4VWRI84JdxflS1loR5UpthZKbe746U6RvZtqZxWR8p9eEg5vxSxQsHiQahwZq
sZzQLHIJHcI4Fiq/ixAtDnZWslvQ6srG4PifAtrU/J7CkAdzTfGv77EEQrj8Usynp9RRCIcbS4vi
2WiY+HW7V6TMWcB4zkCz2deYFQ3kLXgX0lffSBSraSj5vnhssroMj0Sm7jeR+YQccVsDWx7b5eH6
Rej7qmdk6nxAraMewSBP/zMeMuFiUxkTgv1vbdmtf+pT+zziGYsc6049yTa//gDUWvPQnEhcSTfR
57fghe0+qg8mQFWcyxMjI7ox28v6bEngoASg5f7Rq5S/6C8OaKICTJ6wz9yDlc1rM9/4iCOC/Phi
8KPX2WseNQPwG/VVj7iO5uykCA8TQb13phGPWdihOqIwMV6nk5+NullMQDw+eTNH/el5FkN5SPA5
ZODS6+ppyKrDiPrhxvqfX9GRcybPBeV9nTiBRHjluXyP/lA2GoMf1VvsN9vjQGStk3Rw+TZwj+VV
avjHZPNMk5LPYLEeH+E+u/aFYwtCtZClMcIddAEJHGlBuSKanx4M7/ftieaWByuGDvU0CrDnIWXJ
umYzvoN6ZSQTlxtACwltJpnkT7xpcvG8jpry2Dk9aFfrRm+JfTWWs89R13jPZcdyYWJPC8ff2d14
B2QnDXAXXYNbFsPAmtNiHnT7PvqfpN7H6gLFbQRzGkOAT/pu2TFNavDpgvhjxgFSLrnrLdSZ/bWR
fOEqQcBX3WPLSb2dM5rsYLVKst/u19dyfuE6/lkcBSYn0PGHeng7FZ8ERLPYfH9S43qLVb7Duvu1
lu+cqCzuzrCN0dEEtgV7GrdZTjaTbrFdbBq45bfpUnjkggtlArB/EvYsjvGMFNLLcbQWea6i5nHN
w20XOhSJayqaB8FOP8+KQKVLSgv43J8/bIG821x5r6yVm3UNz3Tlsa7hfUBSy/Zp1HSORlDEgcI4
oHe8n/ZVbE6xfpTVNnymC6OXai/Gn7ORKtk29g1NQhwd0dttrWUoRfZzQj5yQ53oYlWuE68ClQD2
3E4/ROowW0v/m+opJ4GvmemcniRCjsMg7wQK4hjlM5bZW3XjNAtJKeuH65vbEb6EAbHLdMkMG/cN
kTWnyZdvyyJnRlf+MHoCsbBkHLl5m3BGJ0RxiahCo2oLZxsYYTwcUbYdLr14wFGMjvyTuoTNHGq0
UmLP08ivcRx+SdvmipkPqGgX8Op8Yff9dQ3Ryi04iFFxS5mjRz43r2kcM8+CtI6m9SmrL9L3ebF9
binILW/2FrCdpnU20sMdRZC3Rnb/X4U6ebUFVfvcXbR1Q5x6xPfeMkuNAFe0RcRqHrUtkZKRNiG2
Ek3CCCLGCvSW01OXunfG3lV7qD73CdXNEtgQvL2bMRHKgnHLDNTkK4ke0xwuTibdsznslTpKnnTx
jFRzZotPkJnUfydjqA9g80ZxbU33DV0mJoeydV17X85FaXhm0O0we8DMfhXCI4RQR4ldwpfEsebt
qh4/hT5CpqxDGY+1daHrHfRjFbx5qK0jO2hHDjzZwQHUvYF7HrefPKZayNIEWNs6bK+Zn7/3O1Lf
7ZbqITYyFxgnJB7Q7z5ztsms8EbuAEkLAkp5bsK1ibcJsaG+5bbfM5V5CW0NsaWWmqZTA8oChcp/
V4/Q8yMIhNOftgxfuEd8acRoqIV3oyyiryvJUToxARzTBaaN9rGn37g86BjKNIAjMcQpnc0psDGG
cTr4Uu0BszFDrosyyBWPYOlcqzvMffB1HRIbaOiQ/JTREZUi5rAODPVJe8TO/dIAM+FE1W239GHK
afTCdxkj0iwMPr9+jwmq5jxcz5FFQ+EzXsGYMATVpE2Gir8Mgw3DmgGLeb0a/pdKzFVRnn37xRPy
Df1PVqNz1xYwIh0GOtGXLJ3lj+Y5lJDWcIHAMILlxi/nxsIQ2YZ5j5PGJMsYqIkpVQciG94XPajj
5FRT4G+S/EM09ZEPvE2Mte/L+PPwqPVtcCS5gzVCZul9tZswoTsbKIpLIxaR0e3vaJaq3psIReng
0oueFuR2hT2Xq1ITskR+o8puKR3BPlZc2woqG9+dr8/sKpTzj+dlYvleohwoDBZNiqJzLqj86F6y
SuimCB8lh8bC8fXx+38dMz2ePRqdAX+qbzlxPF/QKQljJmQ/1yS7lGO0GPb58FNFWQSbhuNXxhE2
DhYnWOLz/TpXOo0YDTUv3nIdGaoFHEGeQQ0ETt7CQj0WZySAnz9fN1SJyxDGypVw8odMZT0Oy4H7
zrTSZVb9DHGfcMGanS6IykUO2KOHhCqi0VD0kyyEA0mA+R+Myw/Aw6R9NR5vS1B5JdzDFrJi7RQ2
dYLpAhHN5SrdDp+Nlzi35485eBF9Mpzws4rnyl24cs7pHxSDxhcR1du6WwAxEFf6f63UO+4hZxEE
VfN7QOvR5Ik6J1xYlUJxEHoLKMu7EdLMvWCi8ZFM4q+Ix+rW8UuiXcvsTNEeMsdVdZ4f4VnKP8i4
8ookmWCYVb5wdYZ6+z3cz8RrIX/2AoHTLgFbZGzigEYf74m1JvRQbq986YzJ4e62uDU1ZgB+mdgO
ymQswWT3eV7S1BnkQZ55ApcyW/2lIMkIc4ivjJv+uRyb5YcKFYaUSPMAvibqokJyGErhwJvejiKL
W6NYM05ojeWvG5aP/U0yUX1Z0VhoysPqyIq0mLDWEJhbT5PumNuL1HFZuB9534dJb/sKeL8P+dws
OCfWJytkT4ogVOKXZiSTimbGK2p6Gei7e5SKT+LgjvLpuwrlOTlTHF/0HElwN4fbJ+oZ44qFm+tM
WZEKYdPOqBkS+CGeERKCC/P9PY2LG1UbrCWXTeZbXPNuYkJBthoqobSl6jSszoPLodPuhAWEWgTI
OMgmgTVsD9jpUt9ZsBKrXrRHpKWUId4gSpwTP2gMp7VVwvLjWOv1ZRMXlbXoy+aO1E46Jd+CLwaJ
x+Zn8vNu8K3JZItmOO4A/AgO2CbWwV5lJcwb1e2kd1SgzjWa67UioTDatf2q8AX9K3tN/yNT8rbs
pOHhGvTqxafzlMBCgEPw2MXUCyHcd8bovJb+On9EWFKpy4psljhsCTKKH+8MDuQAG/UHm0QNucfv
aRnkHnQsfnBGGx67EX6ATEozermcQq9hxqzjp9fbUipacqv71U5XiDZEaLX+DEji07vz6bGTAivZ
Bm77mqUCYIahXEWcc1PuKSklgWKOlsokq1B2Hp1QeHUCwiSnwc2pnDhlbl4fcPrmAuBoLif1VeDn
TEXQOp6UdQ1a/izsY86spWzWA9n+z5xN5zGrPgx4okrk3JqOFmJ7X0OYl0Ns4FMdj3hMdKof624L
bQY0u2XTYRzOa/FHKyJ46N0uMEi6TegpR7D2AQdDxOiOJ4unnRQHM2bSo1xYYsVp6av3hIp0QbH3
g/DAK+2bIprGmXFC/I4lAY+q/VD2nFL8WbgsOjCoHlJGcIp38L1IP+Cse/B65Eh4Sz0fl4N2eKyE
TJcjgiuxKjohbiO2Ft6EGgp49pyIAtbSk4KdGZxLoASU8+Lwja3sCHLRziXoeekhajyMQF47+mKp
61LEV6omAaecQd0z5Iaz9/gJot3I3IbxsfVF3H21o12FWnaurEb6WlVJ89AlORLR2pCNMEQR0HgA
cMEoqKRQ3MXRWYSSgzRUEriPrOFVOQp/Fu7WCmlutJDIsybVb5UmbD1OeRzMOUVwynwaw29PZBBP
jv2lUeU8AstJwAYZ9+/y4jyHeFtIw8vP7r7Rvfpk/LH3HiFZXUHfwh6Cf1O/2uxuFHEDUwtHefEm
dH1w/EYMZr8Y1TSnMdQi4R9mdGOWuP7z7w+ol2SMv70hNoLZzbBVzzhmGoPvDtyni27pn7rZd20a
fq0RJI/hqd9qypKttFvTK5XLM5SJrbIdyoPR2r4A88kE91i2XC0eBsLf1oTqQL0QsMobnONwLmE7
54PVwTfjD4SSNgsmXw/maP3yvLJ2vemQguJg+hAjZqY4W1CPmeHYXDwDKcRsitpY0baMbw9hTa0p
wb/Rvyl/5gseQFHCLWGIzSgubl0fMxUBmAdjhJqW7ma0JntCup3DjVcYMYN/dLm7wzodj0PYLPtE
3CrIgQSXWEXed+VdV23jBbk/H9RfgiuivdB3Z6cG2+r2Ia5CjImJ32UT29dnLR5cgWvmolt80NXf
1miUrLWMwYdtVzGYjdD1aOnylo+qczcT7sJaCXI9pbWGDaxyoMlcupDpCtgEtJ7Mzg1m6oCYWjw2
NbdMK16FZkvVoEBe0GONavzpkt9iPrpQA0PeCr3OtTgvNGsrcdAnyd8I6z2kKc2Yker2B4z52mdg
0vHZ3sTT7IdiH5tA+5FZzALh7NY/mgf3NbtH9b2SC73ThKqvCl9ntI3vQdlTHBjr+h8vxtkmE5pl
hKWYkzEjiikZBzXvSw9PXuyrT5hxmQ7zKSvtBRNfNYeWlnKL7fdLtWpt0xN2EUJenXg6WVk+Q2XT
ze6R+RnkEWWp1KeKt+rAQOid27y+8Ir4wIq5k2z49zvIshLqspaOROyYWNlQeKaqB3ZSSq6BERJh
UQ17R2fkIsuhrdlw4JDywbehF3c3zzp7xIu1r+I1bor5AcvrRkjAk6X4UmROGVWDVGGs9SP7j5Ff
fpsYqoSV+9yfyQSF7G0aITlcpbfOQqJ8BkdkOe0P3ejRbcoBQqnW4LISSjc/mM4INSRCXCyxtfyR
uOcwUiGZBMb3rLtoiTFNwcTSrO/9FKDToY0VCt9jHZqpi73kfZoTiMTwRpRIAujcw2WtGIRx7yQ8
A7jOFXD/s/1GiJwfNZspHfTOP5IGpUa8k9goUm7OppAqEQbO9JjSIP7Rfk4YfyfwqDp+IMVOmIeP
F4lzaFU9hEMh/0Xb+jnnH8De9UWe11sqSipVghmV9zFjSembfJwFA1Fg7Lwd6qopqJ4zh8QFWKkj
7rx16MfFim6DMUekMmavoSOSBFbBf04Ow11OndQzh90hJJrqgoicYC26Ci5a7irqjw7/f1Mb9215
F7Tuc1pGmTvVPFkxwy0I/JXUJj6e4Jw8kCSWFjZn+mj9kGG8jNrENKcWTt523wo6rZChTtOm/ohU
Zn8o5MY4sc70unCBdAwXjdU+i/N3YkkcmoO8qfKyT6DL4rJ3wCJZ2rBjcXe4sEbLXqwnSFoQUpmG
aAf1GOUkAPUGXutDXZ+/f0ksUyYOMezU42Jo6tJ9sh/1cRrxL811ieUXELsOeJT/bac1is5X6ugE
TM7LaLbCUUoZud3v53xND3AKZ+llgMDm+1RmH8S1IopZEcTy4s7c9KFcbtGgpdTfj26lKl1aPerh
DDg1SpeunICoLOLfF2/P6Bs/pIKGkGuSlm76fUZIDPOq+Q6ADuEdCunoNtpWCz79TnIcD1FAr/3D
FZZgYKMgutz0Qkom9bPkNo/6/A2jsd5YzmMn/YORtSniHqPxqEZW5xkUPIIsWS2IX/mzmA6L6cT1
oHpfkIV2/LCKxyNdMJzieU3dYUn+SMR63ZmM9qUtgS4h+Qtzxdo3uMQf55N1Sqbj3UBsKHh/TVgY
72fMVwwenHFqCdKLsWtmXe+cdCApmgyscC9yVru82hQ+y/u9xbgSa6RrhigBqOgWYam9bi9KwZx1
GxnDBcecr6T1fV5Ai2xF1To+pUzN89B0BbRvgioNLQ+8ZEtAkgO/J8fQVabReIkDgQGJOB+meYhX
5BTWMy9MPmGTKRJ1UQvwMzHZcqrAZZROEaLXGVpLSoGs5E13Ki3OJetbETWHj9zXo0UqAmA5DDPR
9q2h6CCIJr7XsE3iIdGL5MV9Lvq2nykRSdo7t68IqsfL+/pRYaEv01FOfgaA4FfXVUJ2fYWHw3ZS
5OuTlx+70XYI/kmlJTgRslZ4+ldnvicyWolmHe893uhbvjzix27CTacMUL6RYrCARb0xZxGvW+BE
SN8szEKOzKJ0BIPtHGCq5ufrYepE6E/ZOqO3MThvYpGeurqi0M+CwPEw55NCMeoJJmS76s2ejorC
yriX2EN83lAINtZtjzNGqOJt/8GdDmFbEaneadrr7yUWF+3cnA/zByL6rPXE37wsSIUZ+UuqBbNz
9j3aUnBTOYajBLV528hvCJb3pWYi6sb5LWMJUowf475Rmpbgg+UxFIePoJs4vC/ZgWcHBp9bz7JL
Oe7/cfmoND1tWWgxoLjzKC8GhkWrBRfXKxnY0mN79ydj4+I3q8t1XTXwKEkgJ1GQmNnfeLkxOQfo
tQWMXs6T77MdT2EpNqQNj7ylqNXbitgI+p3fA8q3u4JvtqRnQkcgVHmr3EvLV95z2OwwQS26pV51
SUz6ej/cCi1xihZuy1DZshyKsLYuq05A4VfVf0o98Csraprqi7feJUwhZ14XoZCry9ZCuSQz1Tk+
5b0Prm+FQB1DVS+BFg5VnAcF4Z3tx8eNYpPxCKs4a4BNWSYqS/VhmUllCwXu8SX/+dfWK85zhXqy
u679uLxTt5/fn5Ii1Anu+9SLFcy5TNoSfAtuSJY2j0ZBq70eVrNpTKSV5hD82Y37uWvphkoDQnew
B2Edp8hdOYJMnvRTg+4rDd9w82w+AS+9qPsxdjeZqUQzhIB/CXV9D+xGqyn93ITJoL/24qKA3U9u
y0LJVlL5RwNcGgDmtk6O1v3t7KBTmn4U8Bho2BonaJENzOg8ktMATCGMehXitCnuwmQad40B5Vrh
77gLPY//40zwLBgo5q4xSbSaYkh2AxsQpmhahVTz1lnATFbkOjepp/1q6M3uO5mXdA3oogzfEicG
wcAC6TOfHZZhtsXt1smrA1ipLXaVB1/B91CmUBl9ZxX7yqgOmMv0nWzW2caDT0d9Xy0SM42DsMiF
eHaWHels+TX8L7o+v/KvTLeSYQ1542qXTiEqlT9qI5xzEqpdJORt4U5Y4VNW8QNIY8n9cpSrwC35
PvsL+VNRNbB+sqTixXSkMBRzTWM0aLlyFNrbgikVuILthPNklRhHsNtAGJmRVcrjLTGs7quSG7X4
oDc+cPh3bOuDsZ5h2mKf5lasK8P6Nmx97aoyHA6C54ExV4tfTIXAM7kLcOfmlMId7CBy2XThnqRJ
pcItlIRSJyMmaj+qr+3wj4iuC5KFlbffowcvku1KjgDSSrinB6xjQ6mPGozaeVL9TdhQ12jJ2WEd
Q8406Ix0wtdRW+HNTge8xPvp/N1OTljb9ci+Dk5cr5In7a1tQg2tWHKccYOGo0wVoyVa+9vKCcZq
PpDRMQp3+Xu+FkSI8sde/WugD96MfXFEn8oa9fDK/Gt8OrXBOrV6KlsmSd5ULykTelPSlVEmqld5
/qc6sSRHCSO1x3BJEsG83xXn22eUJwnlZzp86a6b81VfSm0AYTEfsDRw5uW7ZvMYzhGsJ3xLDHX3
ygCXWdH5B+GYaVwhFSWO50AqD34BUpfeS0zdmSP33q2JXXjl2Syoa7J8LD3yyAmGE2zcHvqlJpQf
g1iSix724+03kX+XAVHcNRo3EUkC6AeZBPNS9SL/opecUWbTo6XwrS69JG2iwRyRK8MGHMTwb68r
utQLygK0ga2czh1K983gzcttMm9EtuyhqMG8xWkifEyfItv0iwfB1gW60U2VtOZEWJQ6GGNPNFXR
C+D/lVkZFyGGLmtdb7ydGndaAEYh/jG/KW5ECV7R5Vt7+8zgDnLFqHx5fnnVVTtMVhtvPQXxQ2yN
P62yL5/34BGk+VQB2YpIDXIcrbFe6iYXMerJb8i5GmlpILFVT1WyEIzaN/h2JauzqXlx68OE14IM
YVNIShP0K+jYjD1Kbuxq8/L5IvpKhgUC78AyIYECbNekZTMMpbo9HGCTPlMO15L7w+Uo+/b7Itlc
0Sj2EesiYAbeTgGPQOyc6nLU3MEt7Z6HurHMYEME3xgO5ggA1uVMwdXW91I6D9Cr0YaIPDKfrSCY
PM+Pg9BqdIoppsqRhTbbY6n0wktOtHjakNqlmBndZqw+57Wq+5kYqJ9Uxo071ivc92HfHu4XT8vl
D6n2jncXDumvbZEZITzItJZ9v+njZMLv28aWXEMaZZ5b0b3AaH8AA2TghQkzuKPVZ8eFT0urQJVO
kMnEbKITAlQluLamAR7hTb7etySsUEncdPDB2DDzOtW3Ew73975FCiAOsvxf8l4Q/pzttvyK7678
/8qRgkiIMytmTaXAsvlpgig8xy7+7N+hby1W2YNfOAH0/bz/2nglgSfu6m6G/H7UjXlIBKVAdSnW
HxrIi8biwdWmObsfS9/wO9vqnyMEpwGnSKSY96MuW2WRWtf3dcYqyKL2vlhbE2H9KhtGk6u0BpCe
WOcDm88Lo4xRE0N+FhPeQiIO050kmooa/eOzd+0cxpVIObokzhhjAQVZ/LHaEYWdMM2dWeTwXmN2
tuajM8gIszRolo4+ND6423/UcL7nQsGPRaNF/V9My8LlF8U/sMhdUcAIk9Vuirm1RjOSG8058j01
H4yipJIL8EY2XFsGHZtB5COc0EfVPy7Ut/aDD/fKB4r9BccA0vLNhPYPJb9aHIcy8emlcEgGVi+w
kTy1DqqZ5EEBJVfuflTSjdKZr4Yph4nLbbvfSRsU9uJiDEmSwk5Nw1WJ9A0+8vhXQs7GVfes6t/w
pn/Mlhepg8LK2zCoCQEnuQuO+DwJjyRZIpVHPuZKj5nJngHTyl9+W4Qd0fTtiZAYzUIsDe4WCMzX
c1j32HKrE3aUPDsahJoGUSHIH5+206pwYJc0IC7cTu4NnCXCXScuhGReYkXrc3vhuyRqcg7uImrN
8w/aA4tQWJUAp8hLdOeIMb5Aom34JW1Czy1BliNRmuEGJhb6yp1AfT7Xkv4ZH1XX6ERjbkOSy+ik
/MaGNVt5Mx6RQyS4Cp6X7wffZLjY8BjAaU/TQCB3E6YJdF8a6T6XCxajvt274N6cgvi5ypsAamJG
0Lzkn26CzZIJ/D0oCx8MwE640TkCG3CxOJkycet0uCx1rUiogk3iFKf8sRGgZ24sugDYsMbLsbbA
3CEMvSLuU0+/WpsBWOQzBkNkwma+i5JEXi63YPx+fIhta8V/VL6UtffpQGVbyx6qLyhRcL9CW+UY
x04rHea4+lq1oNueLr31hweypIKHpu5FS0F3fEJTqpb2LUB57ZDAIxBJZZSL6QPDN/8RIq1lzVpn
qFm/ic68UUq7mcRwLbEuKkZQiuY8Q2dHuz6U9XyHI2BxTOtBw0NQqfyW2tD6CxqbCPwWUrja7a1k
ulUOsPD9/+kGaqtQtXMLN71bCEIdFsVehocFNMufPj4VwuAbw/SVTfkHgDkEslsiPL6ZD20NDVr8
o0gpLS/FVlMXp8IvRjvXkWF/yGxv85CcI2FhPzDWkVhH8H8mQmaKeM8zqPJEmUBNW/psFFg9xoIU
cejIh9SmWdvcH2Z/RiXmUt/5creLbLbU0KmD5ZDs7/pAKepYCr9as1wspu1zrP5k4qHTGsdFzZRu
hnhhnUD0z+h9bpTRD67lcexY/l46nMmg/JP3WTSHfNONICkp/ufWVcBVFchIJqNy2Byv6+nUJoju
f8EuiCaQkDWNkyH8vvD8ZDTj51I/U39OYfwyd6E6Sy6oFNMupbkkaq8ICY1l5RlNCTqm4RJbiF7/
jk5VPxcHf/nTHB3BEIxdy6JRz+W895/SvbIwYUx15S4HX2EPlxtBt8g7EDVoZVl7Mk4WAuBSuUGD
7WE73SUDIk2qxp2NHuGRa2Y9X92jWtpjaF5pxUgr6oGmBpl5ww5rp65dV/TAF9Yw7soG1tHA3mh+
rUuyzpGa+3IZeRWf7DusWGB6nKyezyEwUQJ0cUrrIO0e3Q85lW0jAttjGX+niQCKF/5XeSMX+Dcy
SdphIZZrxX9qC0Tm6PiTHIoVrHqN0YBT614+FyK5sw6heP7XKiA8fC7DE9zLz/qpsBgUwH1qBRQ8
h8FZ9fmuCqFtT9i5jJqcS6K8a20bm2MBXemNH1/ASARSt1y0XluitdgXelQ11YIet26uVAVMPyWV
vC1hss+bGuWOh/4nfY0BDBe85pW/9JT3Rn6UAyjzxyuONeEnncjZqVUIOtzcZoLLbvqhYWjIS1SW
7l92QtioTP+71HLBVKF1yJcbWPZmlUZ+ZHa+HIZm9rbhxoqotIH3JsAArxk54OYquksQJHK0IteY
MOe/ANwhHzYijau/MuuU4ydrskmQn2/h8QDG6FixABqAJZzrTVWhpvPAOFQDrSv98MbzWuiBbfCj
JuciI4jJa7QwBKtk7DoAjIK5WEk0404LZQT66VJwK6EcA58WR6v25pDYHN+Y4FunWxdrNTCoAEC1
mN9GZPIeePEwqYD9PVlprC3z+vs7O1THfkVbjxQMTLbclZ8u8Duh/Q85OZM8rTBEOnx4qYDsJYnY
FxphkTdqsuCq1hLEvyXkksjX7CWntQgHClyuZrcBdW+Euy7GeuZN0h471l9aFiJBYLNkbDsRaC+j
5U3SEwD22bee8pugTLqKUtp3ShXWonbjSuOgZjrafkQy0PfHGfU+ZX1OfatWc1El/ksGJUd5myfY
J4QNa/cnlfmGVi50UpoQRvGBxmhlJ2Ns2Sq9LSWzFI59Vzgu8syQcI3Kf7lwGAkd+fQykncb3ZJM
S/7qEiSK3gw5+OfplgEIJ3whLaohwgS/3NamrYNh2X9oKficYcNVTRwSBuGWoAYLmjbHxbTaITAc
MUsJ6vZg/Y851kUhr68xRKZMqkYVb37G4NaTeSOIPYCNV4AtWCHCt/7YH+zjnxqMCz5hJe5qR8Re
7o1mw3W/ELtpa/sa7H2oQmNrI2RLOHwHhTaJYiddQMqq5efAqjtmp6hCyKgsfuzE+Gr9p4Giv5Lu
UPksusD3nIiKHpvJ+Z0Wsz1PojWzh2u+2+0DkGZgPJ7BSCeDLgOieEy+TZETlwxyk6bSKOsYKBLS
/aj30J+C+HZyn6WjMMpOs7XOzREXybS5sv9tfnPk/9de4LuQM6IbB5gdjCIjTbC2YFh4HFAX2n2t
MHIODrkAgX93ubXurkTE+Pyue+Xh2a4lkOmvUcm+Xl3RzNYSK0FLT/AODmwE6DhCF2UBM464TEZs
24/gcmgOg/C5HBNYtg4dXP2SHwfOtZaUjYY5fv1vMQ+TcC/iyJ9jVcQY0KjC2u0yat58Hw1xAAY9
/MP1k8rhc3/y0VZi6OsJ0sqWHQ8EUD2W6aMn+0F1mjP0v7s3Edad+IJHeYueEnUDAHyatb1yFiiB
KlnmDxHnhDFtt92M7k3ozu2eacCyjG22PjokO2pa6bB3pKgfBW4WgZFVxL4tKlTbOYUVU7lPH9Tj
BDkVmFsmxlUkAb0PzYh/wS/0Ul4QjDAm2DRoRl1agEjQvSKmtaQFH94r7o3+ILASaJTW5i3npHWH
Q2R/UtRXPSunFSuatNDQ9AVaVMWEVlkw59ArMQK9xTt2g8qk6hpx+WFhr9p6v0KUBWtWH3oowZR9
tVyLBzaLcQ9d8q6rLvYcij4CSE1J8Cc3Ztx9ytbTY9pVEBATsPkjHWmdiu5JTCOn0+fdzbA10M3s
VOJEyWvWyJvMg+7/Jle/V0cJrZ9Go8pNSfRYRye93Tv+cnY/5T5e3euQ6OwlcfvX2Zr8abZ725YR
ya+KenZaYofim1xI0RL1AEp9TybzPd1W1FkDUums4mbYSypSHAFdYOUHCP5+/YvT+gctZuSJXuG/
AbgcuzW67TrBh369psfZzOwb9Y1sEU0Z94EU5lMHDVsPrJxGaW8MTPZECXLg+VM5UL3gVf3LxgtA
+C+edxGHS+gmHUf0BUaL1DFWoz/qZdQwfJWGDY1XOzVK9d4Ew8xT25ABFV2Rvo0jbwN+sVlhpAp1
4BOgivixItaqXcqLuY5FsGK1nNRmrx07HzCqJunab6Z4eI0mECTJgimBbjIY07m1BSmxolprPfTY
TQ2q41xw8cYsaOv2y8dYWwYfpce+Oi6HZBJIjGE12DQKggzrCpp8vRkeDWfcwWc5ahp6cWpIZNGq
krB90DEaRiiXcSBsSJSB5ERxJNtyL44QZG5k72WBaTxdiY/qc220pQBjlAtNNq+39ZRFR7grz2h/
Id4EQhWXBX8RB9zemJ5zNwcK/j8F5G7WqitKmjTKS9OQ2O1ehEeFgBranKW3ZEJogKztOpgiPA5R
cFqNmNVFOSU6M8y5sFqgDc3rDHbJU2rZgTAImdbK5utDmAlod75znaUR621LmQltyCHlLOeG7WQr
HFM2V6oo82RjY/Yu/PQxlnInguJPPCfJIa5f7mfSgbNzBiBO303+t8S1rYucXH1O38Hl6dJQxwEk
DqUzOceHKgiswHC50n3VCt16lKxtXPnPZnkGCRp2Ul1UOXJm2WW3Pg97TLfFjXbKjHEtuKJsd829
bY5v8kIbYA8jbmPrA2TIXQGvFkDf92J9G8/MSQwA4Xo7ddKEL+oKhQmRJulObpZJn+a38rhs0kU3
RXE6sBHOJpOQplHipg+YGofrU6rU+6ovTyKLdcfXSs8hemZqZw0ItmTrb1xW7caCsfLNBU71R5Qh
wjsUnQCPur9KrNyaJOsy+BYo+CfBjgZoRSK0nTwXtz2l4Da9zr4sUaNxZpwRh8MtZcIWSGtu7Qk2
Z7ZggUyosicJCciOf/ZvfeELwEEsSDhvz1TFKLOBiSR0D4hV9kpX1XzE8hg0zbUF3usSR+ywpzlG
53zo94/zaoK0ni99YT17p/8bmQZeQObBtF8whrYPbh6NRf+r9VbYhDFD4ry1VVUdS/ZUKVnMTsng
X30lAYT8+Bvd868a0RfK0amcKdYuGjxKmvQU9oMP683XjcvnEZ3MhgiOzjTk0y/yGBRAN8ATTnE/
oK17q3XkGaIjYLXWTjBjwYLE38krQiTGxD2fvaarRY20gEvbZpfcVOOpGE71u8xnmUA9KW0FkL8x
SKsTMq06BQv//0Yq6mP/dfJeNNdLCl5RmIFhFyK6Qn483B6fpVzsjD/h5i1JQKS1fuE6sT0EC5W2
kMe3cvoRnFq+rUONDcN9mixOqgH3MIYL4TIYtfqOu+DI+pX75wkVt+MCAPgSR/spEdC1rKZ/1lhh
RGPZElZx1X96a/pz/p00h2zaAq6niU1Cy+YNVkTRHINNQPyhGE1028pw9rYrdCs+0XOm/F7uUIsl
NSR1FZ3uLaMBfIwkpGp4WWF0vVuQ027v/J+GTK36fdA6AVlyZTZr43Jc5+9luXXR9M4cm+3nvzYm
X39ryFzzy/goyUDQ4bVfqsHAIR6/Ql1GzyrdaTUVxeRXnaZzO6nUEfmFfDCAXVnD1shlXL76ko46
O1UyZjFpmCo62p3qQp0ZqMXbj1yv5vQI3mTHmWofWeLE9VQoo8au41D/brkCLwHlT1PJyq6zaPDd
njQELkYvfGh7POjWZ3vpGJtmLHcd/4aYJjXEwZdUm328X0sXQrYnPb0ZowRV8UQEH8efzZDiPeZ8
mo/O+RbxnSfTe8G/KKytbgAbMTBR61vkY4MT+XFmaOCt0AK+/1EPIRMde7LOgmbfpluuLHjK9uWj
iU9W6zWpSOVBe4YMeL8ZCUx5+74AIC/YOALpeGglvR6by+DU+LM0PkOfyVFc5BH2kCdLdbYb+DP4
1apvx3XF9rn2cd0MSO+2iWsZuU7Dxqh6gec5Mc3ByeuBe+O0oV9Z8omU3UiXufB7NO/FMN2uobGx
yj3nuj+vqo6XPiR0gsw3FUd5dAISkvKmWnNtygEXQW1Tmno5bGQcpJ65IsfSopG0gGtsMeL+zT1s
o9InYFzYPj1C5FqCH9P5rs6cxtp+6GKnfJiFhk/Nw8WeCT9yePNLR+UFH058p6Qcg7APrhRpyBBQ
la/vnEuFBQWxsIPzGf4xQCg3kUjfnMXw5X7amTA/i6oIKGYN8Rp00hI6YZwPoNCoMI4LHO2WI8ME
i+dTCLRG40S9tiqxqwCkD/Nra1B4ZaN9zZvH4U+uoEm/n4xUApT2vUdZUbnV3zUX6NeC5uYoQNBr
usy2jS8IqXdEl1I4xpwL8Sj1GSdSx2GOtTgRNySE04+sRC9BCH7c0qT6uOV3kP2Cuf8lCLvdHK+S
69PV1w4lQv7cga3OGRblk5abQC+eQtyVFw/1dI5sQaqsnonpRkgtCqUz1c3ZTUemeSQxkks+4KEo
rwoDk1njxDg/NZ7Ik47LS0/y+4/sKcXqP4EnS9YIB8TVjeR/vX1lHJsMH6z+GIb8RCYdR3mMgxL2
x3UMW8SUq0D16hLS1LKjo+Mgf5Jt5V2mOD4jl9LJkPygjhL50U50rBZET1+SHnP2rURWnUPkwSxb
WEpEroYVcJ88ZQAqgH7D8B8pvxo+/BsJxUlBu4EiEvxCpCHVPiCz6eKLsf/Wns0K5NU0uFF/AR4F
4TLFi5rY/wIghMerSRJCaIRugaZdXGn/GGeB2rz7IE1yIEQU+vGMN27pQFx2XNJ0blW8wh629yg0
1jBodPt6h2yCSUN9cKDjTMYY1ULFni4j1r5rmbN/osxkVBKaQ1ZDVwW8rTUQI+4QMRfGbYZvu0OI
wQz0/dxwzSijEFP2dHY/dh7iTP8KQ7PtFR3DzFH/Q8r/aV+4AYpOvSuXJxtDZhBCRsRYYeAIB+S4
6LL1mGc8u/SEpB7wYqbuwpGnLc0IjSmS9x40gtSiiUsEIBNOZvh+/NCkLIV/l1YZnz2+8Ffiq4gU
GZ+SLUd/d1EZBdQzaMI1TQLVHyNu83NPA5kb/FB71A8eNKWF7/KxYFtZF2e0OuE2xNl7AdqU63JE
dzJVHlnAQkThSJtUq2f6ZChqQ7Sk9rhbAeIGLgakcufPg7AFwOsoI/J4ZGIqOJvxgOJMdKAqZKIn
4MllxCkUo+nGXMiJM4vUXGFT37fvgpSSkwDh00BuspQ6+uySql+jANgG6kKZK5HIiKvncdQN30HT
xeUFY0JXisbCruFUIALJ0RJw3UhKoF5Ks2fZAjTTpZopraxniRxPvJ3F29un7GVoc/ZP16m36ifo
3o8BN321KbKCLyE2y/t2yE+k+T5URaxiV79HBNke4Od64JNoh9jDPVr48fdfEAbPINd5Ep9jXrGb
8ehK++ZPRovvOSqyua+y23KDpKJ4lp99plPb5Dxq0lKxcqkOZiriyYkEhuM2PLg8dsNoF+sK6dwr
NpVcUixFikkjSqwCLtSQiOBx/G3RYBVXxmGexDbu3wCmdN43kpc9rRikTldDQLVoo9aXgg6HemPR
68EQrkagiH9M+fS/jXXyCq6LGFIyk8KeR6sKlkCzLXOc7Rd1hRM5vJCitFW52SIQ6QP37UHy3xPq
SmP48sP8u2ipRyEmVbdILhkAhv+c4vEomTQohIMlziWSOKLRe2TgSod9qWFRhRx611GHLlfx7gvh
w8RYZL6C3caCFC4aF7hjZnNlX8rvYsYDZOMVkyZhhOE+nDwKSmNOdv0RtX3AQIZXrNbMBnH2y45X
bL/f4Jg3gecBaN6mg43Za1DYe6Edm8Z/BcZeki+tjtTh1lOVAGkETMMQO/HEoS4N3lGRw87hr3lR
3zeFlmYyWnHRdG69SduIKu3EouWziOJ2xDNfsiT9OY4dijhSGO1nTEwOEqgi5de072dBCPzo0Ouk
3Y8IrW4IkUP8I/8fNuIRwsQhMtqlphkOmLlMrhIuBCNbRvEcv8fl0LD7iu+nSMd4x5BVlE9ZppIv
z6481d2fCUaWTQUqY5HXVRo2u90oqRDHJgmQhiLj4QhwIO1Qe8XUPHLtp6prCnlWGKw+9O+ThZ64
kw1hW4h43+JMS8jakAqX0Tdd0tnXDWY2Pl03dC8Ku9XlxRcwDj/STN4XAfECiu5kunYaFZ/1Wx7K
XoXbJjBP+vJaitIyB82SI9fxSmaufvx4GX/wCm/GTI8/OMEEvQhQMaTdGVyLbHpR4n7hicfhAGUy
sm0sVw6Thky6MpjNNnCSOlvC7QUukEhCAAwikNSzItqF1w70annptWjEZIaTRxt1P6AbtFd9Tcor
4/OY1ZQZYRjlFTncopKj4SA4TEig+dH1AzVhR6dfsfTwHybt1ZvxzW36KmrPyrR9dzfMsPyN4MRC
4K4MgZHMjNFDUxKBt0KX55oMbquPFN6pn/p2ZMShJSjKt2z+lJo3NhXxewhmYQhes9xwJWrYq4Ft
YNFtjF0o69ixvKz4WyR6MjnOKc9JIucnP551WH8Jj+Nn69Sh2lv2UVv/ojWj/3oIyGgHQ1yjl+vR
fbVMzqzQQCtdJyfv8CcuRphspD9KtgyzrUPmxYkaE40k4YXl9HSBffr5fUzHTpQNSRpM2BvX/vWm
s+r1qaz0Pt1H2l7VZWh6C///sgEfqcwA4b0uhBE6btufXhmxYsXHCwjBni30apxPgbhDrWGGE1cx
5gCJ0u0gMjvoeM1psNCHrwdzcEYW1IOYoeJyh49wqZW8AbRq1/bo5Jya5J3f0lGI3Ri7lpnRvkgE
RDOcThSfFdF3p35eGIBla0Tg52ZcQXRLNm4NG0aUaiaf6d0sZZf8fp5MZGwtNmFeh4x6TGxQCxyW
KKT/5JHwmVxVGmnlphk4YnG96CQvhnz+LTSUD+7/lz3JMZBYc6wyKaY19yZBdcqBIVa98Qux7GHj
ZsbpYNn3leHZ6kidH15EK0TVG6S8Ujg7eI1aKEpUj+aDosasMm48RRzevjjKwjuegzzZS05N9E+/
kRBICkZ1isyd8u5v6S6J2Ei0GSOGtHjTpou8yreixCso9QLf4zIk/k0ou78Ud9sC0/+/gL7gRPyD
Fb0v6cWSIMNOEOTB5vw8LGrqtqioViC9hWIjY20uHgpvxb8RWeUurpZIWOFcKZbsd9GUjc7d43dU
BON8aI1KrwH2dz+rS6HkRCYVNj5IdtYhtdlytc2L9lmNvMNtyV9uPFAQB6KpyDUSMZN1FEk5wffk
2FK9UnBhU7QH05FJxVnP0RAeSzJC+/7s02nzV3KCjo4fz8CiSyuYpMLkSJ/ZFv339WBPwL1atdVD
9sdsiOotNIPQYsnTbGJDjIhjIIz4+PFhq8UtxZVx0adqKunTRObnlFG9533UDK28OkFYYTwzYcrW
00WUDs6ktyqme6DeZEFE0rmtNbZ02EAWI/l3n//ecvzK4XKTZ9GcTpu/TSfqY9MlN2SfH66twGVg
Y8wtvUbtIV81fd8bNqEWxF1QFtQcSJb25fxPG+G2oe661Ocg0sLu/17/Bsh8+RZmQJ7t3fKnkdQ4
XR22QUucob+cHlVJoeKBGV4aohYnvnBYebcsX9T0c3tBKbHOqCyxOl/pv9Ok9V7z9eiiEJHH4c/W
w5HpPeMvj14FQcI/LxKdR/X755fn2+KxzKmxMLcARpBsoEvhox/ddBfL88QPyuzZsPTmOky2c3Ho
C7iW5yAqvkBVwotnW1aPvZuypxVCnl8K9IsS6qxyVy43Lt0JoZToi1cQbhiAbDa4ushaLwnAOpmd
DRgwocKkwk5kjdfrZtlEGwbj8AmIpAwQ1etewNd4U4TXTWn6kpuSt+pJfEb4kOBhJmjKsnrs/1Ok
VKLxK6rVq1l3BhKwDhYvUkLPycEWUUaB/ZI3DQGseC4AsC5NNRgVYTjCzwW+ib6EPsiqVNnTMv7o
XlTJoxMG4OeQx2S9gOYevu9/GPGGK6OOXbj6CQjdoQXU6UIPvvS5Zb7OVk4ASdz1X9+D0Oe1sCpB
o8pzCJjse0shfCDBjMkFvgEMWPzbXV52IpIfNUllGjryztFmhEgOZmv07p1U4mS4Hq2kcyCo5hT/
FNSXz8fxS0iMHah/vmb+w61nRACDhgq3HYJPkj/PiHFrZsIsQhnZ8Y/sbO47nA46+YPxEIqnRbqZ
cHg1Di7K0dDbqaGwBrWMC3bWQ4NwfTWLXFG3BoJxmh64du1yU7MQbup6vXrknj+eqMX8IsKdcO7x
KrV2SzeOweg3aRFIOcSgns50ofwPLH50vsPV1I22rMRBYk99TzTUZnZ5Mi7IV7P5hilRDAvt9/tX
saTN0fFLTKHHPiSYuTJDhMzZJqV1usnVk0KLmvJTNYtLNMerv68opOpm10KRVbKNT4bVsOYVUqkb
iIXrNVJGnI+JenvGFA5FEeUBTC3Jh4ambIWOIuG/ii7o54pTcIZKvQGerZWWzSktt9h0yk3gnMZb
9RLHFrbqHulbbvaLQ/GKImFSXinPDZRDiQs6Aht153p0d7AAUi3I3rEaT0SighfvPEgm/JkPpJpa
6xm+pXgZATcP6iHXe8afkA4w2lpkDczOnhhiMUb7miV5By68cjkZmtQ8zRIxMzSMRpgALzMnSBbt
kwgToONoLT2nSwzrVFkAW1KWgqiJ2dlOfTXS9rOoxQIb8TxqxV00K8C6ugXarYD4rsCx6IT7juy5
ePtEhIs/wbOdwqqFP8sNSfa/5do9/dLJASSTKqbx0X2jmzmUMGyKGNY2SDzkh+ZSZAXPJs6e8DpK
dBjQ2ZQ1BTwVyAFHUOIETBHB318zvHOD8A84GBKMDc73tf1dsjBQP23p86BVEPH305dtAmJag1Zo
aCqiJ8ZvVvXSW/IK/xxGo7HdMrWG19QX9q4iFylvwvEOW1ChLJUj8y9GRCvFSVWzAMUKRmWjAtUG
NtZM90vXWO11ATtquZXGjvSrzjtMZsgcv5K8q5TWTyyVxlcz+RyVOQe0VhnLtdkaBxpxhg6XqVf8
BmI2pwlgl4DmCugwZv1xPC+8UQ4hsjRClEgDyirLCrGGhCtN5b+7R8/771b5+4oAtKfSZB98jHw2
wvdO2vVfEW64XHnLYZl7qnsdOpJCThUkCCHFCRYR6gJVbaJWqMVMzT6DsWpotF8ExDUe37P4INoN
LD4uN03TXyMNvPXf5isuF/Uj81mkI51dSPjLduOIVk7em4ty5OrfAsByaFlULgLAvXXNvNdagJal
M9anD3UUQsKWOxWoSKopHZhISQ+FpI5U1bo0IFvTMxFXCV9mSDi5IWGlKe8eDSxa0IcswxZfMLV2
2ZF5J81e2eAOU3M41EabAwCfVTPufaBhA9qP//yRxz6URsXEgpzWhQErUY/IoqRDzJBvQfK3h2OX
d0uMfOCGkMb9sW/x3UjT+TDOY83Sx6xNNKo40ZgUv9TmgKr+m86X6YKrMmDHPdLoGv9XXfeaWJcU
BCUe9Qe9f/ZaoYkGicV0yaoiAIEoRJZ/mQTOMc+D5gT9fkRlFpmbfyZ9nlB3VnSu59Es2u9VD7Q8
GtOB7EOej5Voe8DwpOWo+QnCgoBs7XloudU2ejWZ24wmYVt2/Phz3h2wbIHZb03ZKWEy2urW8vTn
LNbFtRYLBBg2ecJ6cQcjEX4txOwgzPztu/d/fQynabtRjjMphBPPM9dU+8Mvyq2AqyX+S6uRNICf
IHNQgoX0OPmyHAzEvpq3fqIc1xI2VUmXLI0rgazJ0zgPH89aVBWHKR58ObJ1rizFMXgnjqOIv5xZ
jfRuUnfTJr1zRrCI2GfDrdKOLEQUZ7aP0Oj6Fp1lpqtPHINyLrwhC0bxIwvKxNsGRNBEuZTbzer3
MqTEXIo9cFpt328Zu0DNWjqtNxTnhOd+5uAubS5xxY++CUzEmc+2vu07fbU5lZDwCOpWsr+a86fF
OPw97dDB+e++v2LQ9sBYOkD5RZTbbOM/3ZRQyHhvYmNOGN00SSw+c1nRO7NLd4F8/dTDls19QQgW
hVCvuGuyBxjYtoaDiA2cjLO0yketHf53fTrIDx/rgDonS2qYuwm16ydomw2Zai5OaeXUAyikC0m4
9pvpEhzS5F183wpBRCk/0BkFPAREMANsl+F6VLgDmhKJKGHZcX8IXnF/uAY3Q585f4c8UUNq1Fu7
YpOb79y5+mlRBnZA38qAJ9yTcjRwuCtet7Eqzsw6NYRcVFP9zr7f6QAp/bFcVEsrFmaE+szIt8Dn
q7n/zedi9vt+XYv5E6LF69VdeO/jr7tw+KisL31IsjCs3qEz7My5HbaTx7dzkHTs7cXImRZlJjqB
MOwTE0hSjoQUBEqhWC+pdfyXdvPU5/G1sUKw5SMvpPiqBpChM5Jo8cCSABGpyQw8Y/zQNfPvPA/1
UxLT8qZW6ie2DnfWPcGUu5B0WgSam/xABN3qOMh891V5gFAHoFgAtakyT70nKgxcjgkwIPjNdGrd
FYe/GCJasDGgI2HTP+QM6ByXheEGYxTsEZbWJVMuT/AES88LX973gHpZER9EeNTJ/CyWPGFEYIAl
N6TNg9WPQ7WdCYkFtEQ8O8PikgM/JfDbkADKoXAyqNbPALW3K9MQOIPXzMA5Z2dqzBZ+P3SZ/JdS
6aG+1Mo1omlWvGsfe4dQul6Mi7UiYg7lEYyne+cZCA0u2Xtt3H2ZyEIOYWPkd4DBr8nt4WSXhEEf
ebVb6+t+6k1zErNG+wgyemxI0zMg4uF1M+2Mod+2rB29sDIaN2zZi0VokG8t6nr0LuYAWf/eYG6P
07+NOs4f0sHE7jBV4jZ+GJqzOJUhuhppy6Hgp7Eab/UHFxvhTku61qMy+SfwdpM8SEsAejuMz3ZF
CZ96OTrhxBrbfUowqrupOC1VBZaNqPsOOG6muZ+L6RnoBGpozIaCfKlYXxnUpdXqfHfTSm5yuR+B
Db5GhfecZ/5d2Ybc1esfdtfsoL1asRl7zk6S/vFGTjooTN19/SWCUiTwHKyqlPBcOqrzSus4Fxv1
aIxKbR6HFG68HuaUPcRcUNmZOzuLDyuYQ1sIJufDhl/ZnaKNxp2N9xFCdoKALcmODokS8jO3kpl4
pA4S5c/2dsk3lAScN2Po0qpCtA5Of6/R7nZDdo8AG0pY9v+ozYAMGrnhF+4dcM8HhDRiDJKG4b1I
l3EKruqeTI3hxYF4DZt3dxcT/u9PNA5rAmts6HVrMeO6KVVwIR0yltOTcYg2w0UyLru4KnWHcY1n
88au+IjPYF1wEHIlBHuYXNE2KWPgQ7zcGnsMis3oZpMdfVAcb0030aGZALVo5qkODD839pnQpaFh
YNZNpI0HsM/xv73MoBYLaQA4c5D+8KoXVqnk8YkIYCIgM4L7Af49XSgtGkIgEPZTv047OvR6O4w8
qaBu5JCNfDomedDS+WLmtW8vCUmgH+v6KYLNDo1Iemc+lRiT1FHDqeXW7pSnoqi9Ms69fhhWiD21
MJvMwSu1fLtKdzZadL42M/Z/vtSwfBofE/a752sos2kyYIz2TRvVbb8kizzhcV428LDaotBC0run
7iDkFg4Q6UfFsPZScIIlhF8xiexF+EzQFvKWfHNqZgyB+uEbWGi8ItnItMpvmEyv0ppiAZ7jj0XD
U2hDBbR4ugW5yq8hdGP7HJwJhF/G2ZL4W+f34pbDXTOpvw0apTVmGExW/rwGstPRjY8+Rb8zdpp4
atK6QoX1O/KtwxYqfVeJKASZMbX0IyGBBaoo2EFSVTTJutiw4/WE+tSZA6EiFFMIwg89j5O28wqD
qMcsXpv9sVxdnftZHVCkG5Lyfmd365/PQs2Hl31D6+Q0Yym5IZU3kkoULg6UfJBalM4sr9XpfJCQ
6rKop1v93JUCuN5f7VNdsMQIpqD3QdjW0DCcsOYkpyGjpg0vP8TQrPOPzm4dgA8lnKmpR5FH1LHD
UDMIoeqgsYvybrePOPpeGmq5ffWNAI/i9V3OfN9c0jwlxLg56o/mHMdljbz/T+9BhUJtKCATScGL
Ho4mXVDeb4vGz5fsoRY4nN+ooWaffSQrtzxKI2meuv+KXjfEkY7nYu6rabUE/QWsyOGOZG6C+tFY
E8f/OVsOWfsNXgT94Y2BqdS/mceDpAf9vHgXBEatuVI6E5Dcq+LAR3CkILJfjOsZGJo3IkmL86lS
dVcYVo0cIuJJpkdalrN4VoTsI/OtrYNnvm8BbVvvL4uTvCb09e3P60P7kyYKFMwahrgolkx8aYEP
3HlW83mb5IVaJJtRjlrXoz60SGAW3c+/JUKp4ZkSKE152ozaiV6KRG1a+5shlBQYprmAmrHOCpfL
1dTzJYre5bc1udG4FR9o4Q69M/7imG+lRHCAh3BQhNWW/NXijfnrXJVxGYucl7CmRJ8thcHCD9CT
6awytF4qr+8TzTxr62tYIlWLiSJfGXleNs82FdMkDVdE4o1WIz8HfRgOWYlYIwt13tpDdRk0B9DN
LdCoWPvuAh8L35FlcjXFHOfLq9MTl6OcmtNr2fyblwhipDdzmuluDc5TLBLwxqz6w5Qbw+bNFlof
euVn3bdLkiTHO1CeSWE0oDWlGbyAmIGVGMv+2JvbsZk8qiNeqOqn9kA1vati7U5m3+viJtVca63X
vOTmOAF+7SJF1v36wbNq17xThsfyziOQ9PZBCq8PBZ6deFYDWpKQuyDm6qLPSIWLTInURVakWbIg
mRV/gw1J7deJRl1oG+H9FVqcSeUOt6v6T3ikshllJ8aVkV2JotLgXXYG1BWM4CDbxc/fzTOtJ3Sl
a1op5/RV6q35mGNbzFl6xWu7i1z9AWJlOJ1yosDsBJPbscPfTyxPkOfVmL97AX3pl+hVxlbZRSIn
6MEo3oouHZSOKKjoOq9nkhQ3Ua7Qfy7wsmbvXIAPB6cZzEs6ZEB4gOxhSM0yNcdJwBkzV91g9ydJ
b+0Wps6akHIsaqi4bRa7ja5/juY8rO/MQu2S7Sib3CuuuV5VMqx1T1WOlPmf6zogcnPK6iOZcrQg
ZdeaqKaitQ8LVev6J1s75FN/kXCr8r5OaBa3EgBLuIYS/unW3hWpgP8SHHbSWWTNM/ImvjwH97DA
7/AnoPltP0M96TTWybjbg/jTrF2/1zx3Xv2iMlDwTExsj9YAVn5SqFSOUL9gq52puY9TOXVpyktv
ZlnwqR0bk2exyHZ2MN4Y3mxyCK/1+5weYoYZVZ0wcyyEUCCnxOT+BD5RriKssN4CdT2BYjL17hFW
FE18l6xlVStsawSZgcNhzURijaccwnSmSsuCJ3cdwOg256VI+ResC6b3YJ6okjRwD/PkKVCwdacY
nyDuNl61iHLi2kS/gLZ0+AxPGo8W8pc94cvefYe17qd971OvpfpMicqagSW6iiVm+4Q+SfyqQNet
oL/TWyG1riQYSfv/Xv5LfRIYeKt8v1pvEuqlnct5Kw5+nPW12ODKcYkqtyPpNWcyjplcVrRobpzy
tbtO9uPzNuOKT+c8i6RiZTYZrSHw7yxFGRsqUTERGQf/UwMApcyaOVng3ZRDb9VNyFbvVct4bJKQ
xz7cCDKe+d5zvHww7a/ZboC1bzRSafhoudo1fJrqbKqcl62KxgRe9bPfszxRKu0dZw6VftM0lVrK
f6UrrEWrtggEa7jtAJ3kC2J8Wy+8Wr4w8yXN+WNgorFDKywv4jxyFb5Rs7yOvsT98ekLt0GTEW0L
TG+kSUqP2WDHR9SJJinntckFCLiXYJsEKmR40Z1nKJnxR0owgaf249hz2PvrudVm1bn3RkFnimHC
HrtIyuZWMZjacYWYhUf2CGkSuZaS7Yem2glZeXiqXD4X7/Dboz0sSTIWmjT6v/h1gLV7YCyGz7VP
1cy/C5dlCjZcJRkLeyTqLMNARVKYOASvdMGwbo+IeCTU7b19HkRPIlgmhWLEKLgdVEzBOXFY663M
yQhj+4QkWPexbXSggba16iNFDK40r20NoE2fuyBJHobUByHgGGDY7ec/mk8p/N0XxekQ2XAj8RdD
hQFEtjkSfhXZMgM/Po6fRfa2Zhv6TCH5v6a61vNXdaTnGSn+2tvzKyD0hadzlNM5/O7Tr0V+j40h
iQlDG0Iei0mzwQz2QmaQrzoRi3uTIdtffvUw4hUWE9dpNc4x9m6An48P+VqRGXPySuYAIpsOZgH5
9tdfLJv95StQvAUUl4Z8qg5uOjwihZS747CTN7bOyy1I201/xvIjEAPEl1di5/pySPUxEYot2lWl
E3ussp0ldZqUJH+gm298rdgesRVdj8g05cghuchRwutZJGs9g3erIIIsjtTf+3kmiufCvWmQNQyL
uVXYJJ32zy79Mm0peMteht1HCdgSnrlUskclMUwtQeDWUYoAGkSG4/20uuZuoacsO1tCoVuuZ7tQ
mh8Y52KluCDCwvKAIgyTo7Y2hlczCsfp3MSUtwJNJJ7YTwjJsM5wPOGIbsatUegdAeqgOrTnodZL
0E/Hkc9qOcA1BvWRG+Y8tuH5+2tAWQBSvNyhyHqHpyo4mcx0a9VSkTRyVDNk3FvWSKw0bdEafCTw
RbGqnjibxNsLdc1rqe65fowXDNMdyQnjUN3S8HHMctnym80x66UUgtMeW0qlRmKTuWuakJWqBS6j
ZN8VdOaDRXtvYaq3DgDIOjs+52ok9/WKFtMUeTH5YrWiahlm/BWHlBrOo62l+16IVBU/84ADS7lM
77xZTGK4/MyP++JHWFUEnRGO3uCITlL0+aJitK4a7vYBIbBO7amkfjH/cJlNOfLJ5AWbvXMy9MnK
vnfnHk8bl23AnASCUaAwO5TJ2jMy56lvZveQNWlUFdLuEkwZnXwn/Zsf7QYtwxV0JUmwXuT1wsn0
NVyXMeFWFuZsQ/2u30DwqGDo1FLbB5UE8NliyUoQAimq9/MsViUmVh8qOIOQ+fK4j0JhDKwzyHo2
vfmYfeA3/NpDBI6iLGLMvEsrXC9AUU2Eea6KGMViG8xAjaO871Nlo0jFNN/1Uz6R42V2TtcqspDL
wlMpCoZC4+RJi01RdmPPclxaakpUpuKn9rWNIsspUUZ9/rZLAVpIyP0bFA79neYJ3fZ9FuMHxWrr
WLiORBX8Yicwe+yoQcVUxuAVC2femLVkf+6iQ1Pq/XtNuchnpB+YM9vum1Lna+pJ5JgZguhBv8dr
INL0N5/DptCvXJxPCl403Kfo4fG3BMbyv50b3P5g8MyJUn2Mu1RRljhpqdzMGaXRWlpRzvN3kC4v
sk8DSCXQgLTp86y2QJ3Aoz7yI3IsO1wm0ni+htvkYRcoCfrCqIwWHafASPe5KkbRVe0Kvk+yamAS
D6ehJOAOabg3XYQah6o5VHGEcpcsPT3jTXC1WiXoKwvwUv3G1bjlNiuTMwMu1FeO1BzSJD0HwSEy
H+4t1gBsR1u/ZkXyujJz8032JAUo7IntI6ea0brjnjnhaO++z8tc8sOFRIJTRlikiWlBzozZudv+
O2e7J+/xH/mFqicIsIMGNLXcxgLRYZbOITVW6ini6ud3CBQwcviwh0U5Os3TwZds7LfNCHEmgFFo
WaQ32p9ODo6TawE9c2rHR2c9Ntm4FbUbL3qeSefGG5lDQmamtheGcmdC277WqNl4ru8Zl59iPHBi
QlfcgVoTAuyf7QeFMZXdVPp6v1m+4JCpDZwe4ZpEIRrB2cXRX4b7hj4RXkhoIUZ+aK411c6kfY1A
jhHH27Sdd5L+dugqhaXymTsZU5+htkj0vVFmln6NMY8Ox0POcirmVHfOd9cdcxd9Nh+X/Is=
`protect end_protected

