

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
WOJX5Fv2S0CzprysR8KMEndET58Nnshq5G41sUF8nyr23cEOOYS3xFWHzDNrh0BglAkKcA2/EcsL
0Mi0zP+UFQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Gc0ueCwDN9OX/N8ZykP2NxXOhHr0aqi823TAFhXP2T3sZajOBosaRN5Om/T8R3LfwK7+baNKGGz+
UJk1ogy8JwdYWmJV85/JpyrrDFtvClJsQxdfCiEg0IVlJhvJlhs6FCZi5Rj8qwlvbn+/sc8hT0BX
IEC/9Hv+yH9f2HZIeiw=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
gOAtaUsYvJmoKivS2pd7kBeODY1Q4VX+agLZ2/SaxV/BkQgGuuCLHYg9eGdXBmjxTqXO35IrXGnw
8lzEMm8YS53SBgfLbyNKtLJ5Qej5jTli3Hhz2BXRqoQonahfpMOh6WT/32Mi5HxamPl3+Ad8Dyj3
AbqGosJ8LBJRb65Babsp/E0dGGngj0nJjmmY8NHpqNTG489434uBxC5ykK4ltOheXkVJtXSHoR2s
c+RXEPDO94CZYlHnY9b3pUqLafSVqXTeYuw//0PIJQNmrXYuvkdozgm129vQnlKXVGzYsK5DUlRz
Q+VO09C3aal1Ga70326sWIG6XdhCFEnAfQoucQ==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
3INKfUgfMTydNk3PjPUP24H0r2p1C85cOfDxce4LgEKtine/HDrFDahWRWORtm3mNUVaknW/GXSC
5KErdi7NyQ5+CFdf2MMmaC9h7nGYKW8O4nbf09hLlm3blRBSd2i3h46PihYy7iaS3Q+Z7JKvWuiD
J79EKDKw4Kqn3mmg3iQ=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
YHV/PdEXZA1kC+N7hsk5uDSJPgfJRc2Sgeu6l1dsNtZhWFmXeBe9vCszID1P11I6wOICxCc/uQgT
A2JL79m9I3kuY9Ji47hSGH6+xG4kfTKsYaTVdl+16SjuG/YaIhBwQfN13p/8IGQ6FysnYNYR5siA
+0Lm6CwAYBXVRwsuIA3R9dSPKgq+Sbk3MQCuaqKXbxHiA5oAAI2R3Gz78f9hrvy4Cj5P6dJ+TbkJ
j9bOdpZE4W6tXHasCVI4EqJlfqQQ48uWK076fFPDGpd19w+K6NBgkvxxlXDC1t90ZvbdFgDD30L/
SOFjS0BafCCf2aKaRk8VIdeBs9pr4wj9gMwZYw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 12496)
`protect data_block
onN33vRFPA86MLUw2plHjWCTmJBlmIL96UxJA26erwtNzFaxPDq4wwmX5D7N4okzBDmmG36qF6xU
NRbSRIkfLXO4oVQG/Us/3e/c4p2XCtNuXJzbyvCD1VNTGprsweTFgkqvJJxZp4Qol9/SHgYd/o6Y
dujL0a9i2vmDAsKxO2V8zCBxNqIDnS3EwIvsZpMsnUllh1Br+mrpprxaCbO6kbyb/iOMmhHNRv7j
rQdt5n/IVicFiKXpRR+nOeHyH0J8LfZfIQa9wkJY1Zvv9+B0Ns+bYj35pU0GdnNchwkx5qWXFe5D
Tv67Xh9cEbXVV5W/f5XdXSXELedWDWrZJKxPqwswbsj2R2pIJEkOgokfgepqPW30VdYnuuztgrea
Botpgd3cCmxuiFjLWiBghRteznpa72xGzUfpuNnXhjYudhcZVD363jT7lExGQO9VZDJwoC0jLCI1
nCBWHKIDwFkYywWptr4hzyEqo+Ip1x/H7gH5yjBbQlsWv1WE+Pcn27i3VoyG6p/5RAnzngTouNmN
3ibqfX2ruMQ5nmKE0GTKUCAR5+zQlkxxyebot1jkQXmSQxa1+mK7dUyDHUCo0Qeg5uu3yjgyiP6Y
AUBTocGOc0HFeXbxj9dntSRcMgg/RCRk5gKWZXdzwvKuY8Bpb09IT3USxhNC3tJLsdSLvYF8vHRf
Xz+qx16zZNf9YuEef9/nsykzvf33D2h0hEUUp6B4RJu/iFAFPVEb/0DJSRJRGSkPVgNh6kava9hB
21rdGxUO8H/x5ftZJ/0znL8XinvtZhGkji8VGNA6+GTAyvFcYCQ5wF4SP1PmbM0rMIkc6+JoSZnI
b2BHhWVd9qKyNQ/z+TKthc2PN/uiSSfZ2mxIb5eiIApbIjBAfEtZrG4lJ/JhgIOOnoUPh06iciW5
JX2eR9EjLN8WaB9/mMSgzmoUhS3MiKbzcVug2Pk/Qaf0NntF0Uxo6Ycr7t3ASpf/RaIED3WMVIEm
5dBfGdXTj6KdhQT/Bk1HkH2M7Rhjf4KRcYR/e6NpIiLSpfMgT5K3YKhb0g1si4Doopul4KemkRoU
bIoVo/bmcQJAEMMgQeORfpyXHDO24qc45xc3byIb3gzZIRNDw/Be5dfq/pje5++4EGBW8nzkxqR0
hW9zaJ7KN7cpGTVSGrYUDwgDJ+46W7ltUZ5hVEcQQGKZ+Fv7LiGu7QbytIcfXgx2PvVPOumI9yz5
FcVkcxiaSNhtaLUlui0ftx3FvvByIf0gCrxKnLWQ/LdZX8iLfx8RgpTCecaHTcZWC7aSRsF4Att5
OHyvqagifbDBUuvWj1GP3jVuYOv33acvtJLpF44LI3fVusrIm2Z2bzQHNmRCahZz9iTWUKID7+w9
P0UnHJwIy/GczunOK0PbKE1fWx3uekeJ50GUWCfgfNFHkjM6xJY0j+1TH7MLCTuRqYYGGHGbaJiQ
mrteC2/qozqu4X3qj4ZFsBdZ8ZhwzWgj+KY+35Ky788ZvRC7O/Zvd5lDcM3yTNYl+6uOIWUTJGY6
HWaL522RCL3un4paOq2pKvHxair2a+aB1QqCo7ZGOeB9WK+AmflmFYRDWU4Ahqe/miHqoIKAG6eX
FIL//XY3lZXHn3gCmiJ1Z4NtUmi6kNX5PZxYkArZSnOSPuDnkuM3BQSK4fhcit86eujzEEQyAjR9
3yLPGse4CbSJNbokf5emEOa6wc0++BfBVT57IJ+e1vmx5Eu0dquV0ANIy9HwmFwbXrF+bC95JAMc
DJ3OHhHXgSosVWHrBpVhadPLalaVZhrSNzFOq9GnwqiHt5STuY0NaLsp82ukiGNJplcavHzrwWtv
Qc9q270MrsjAYgcU5ot2Unoz2Uo6lKsZNgBKgUDPsv9+Re6SnD+jGzuNCszMeXFm8yQlAcfVBmxT
wVfej8UF5p0RQdDz6u8KAvavUXAWGmcv9zGP9k/kHE/My6uovvtXPe3AYoN0bbVjC89EWM+DTvmJ
9k5MIP72LrsSjrge7+jGAws1TJRTKMbtn2foIXLkmPW53gxaOjKJnQw0PyOhfLVKqOEVwDmbtTOF
3RHQM/HTD6W4AW7CvtANzYQA37Y0K6pcNdk9hTon2u/P1hBiTsM/YS0kw+il6P7NB4nxqMwl8pDx
X4VcDU8jSUzRXOLfuhv2Ym30WYNuSx5Co4OSfImlDAiFZm9mLHhqHq+8znNv3b77cw8fWZgSkdTN
gx+KLt84DQnaf51AXtn3zJyjghco5JeSpFhkd9lmJOvlLLPdTFPMHaG5l/sR/jaNfxSmMSRNhWFZ
GHB40h7oy3Rs0ah0IjxXTq2vKH2G21cpp1XptFZuGxETfcKxgWT4lCNEcNvlRYECsVBxUYQkkpUN
HtDbqJsXYt43VPdg1U9fg9Es+QZ1v0LjlKDSgStI3+fGj0jyJf9x3eKxUTcJUnIc0PVoa1qFEATi
vnV1euQ+OhurHfUxj4iPliQ/giwX6MpL4rkCkhCDThw1Z/L3p9hUMxL5gXAkRVep8R8LCpd7gtXg
DEuvY1hS6ja7O3sPb/kkfziPAMb5ijmyAuhwdbzYoPTPRjDp3W74z9ddl5EpmaKy+ZTqigArzskd
gV+OGZysshdAjpGRb5LWaSyshciOD2hwXei0FElGPfeiYGN1qMw0TI9tPcodGJFydtAL+MYUSQid
0y5ndkoVarsFGn7wZU38rTr0lcpa62otxRoJ15XyOgZzcGencERm5YYHrJludTXM60V26IsTrX5L
OCov84ZrN11wCwP+hhs82yzCkfd0iSIUefy4Wi1s8mdWuDzAUuvrveNKM33qGCT/a5mCeq7uHR7O
RKujINkrmejxvZs+7Jv4Bxe8Jh5E6SgYClX6IDch+uLOfrUAwpk4FenIC/ENqSaG7JLT0/HY+kWh
7k+AhWvSyd/uA7EXpk25FU4P1rocsXbC6WzK6360Sdq3gSWfd3q81j4OGuQpuedn4x/9MC/XzHcd
WyLMy4vQ2iTqhhTbyHnx3RmT4yQ4t9gl8+TfRbq3lLdYF4rwGKN3rAjCIIzc8f2OFy+WmYGL/M/B
2CFIuPn5uHpRdK6vybQuoIJdKnLXI2t4QYnZ4s1iy2hhrO74nGjnrRQX7XzhuYoKaRVqXhFbsRt2
XIN7eUSHapUeYjliLwKzCRGgZkKpBFSWjoNrUjkHtTHmbHHonCnKaRepsxTq0vV6O1nove6Q4w3e
OtU0vhSV9ZY8u1vBfZql4ZfCipu0afozoNceISQC8tBPKr9d6l88vpR7gJ5SX2bTT0vyO9ef984Z
welbtFhdELWeN+M0qQEp5pJsU7hcKULDdCn3Yg3YIlmyB8Wu1MH6mGHGByYZtRfVw7xO5+IQI+xX
5UgMoBYZIu/MWEoHzCUHfNqImu8kau1a+ZByzP0zubxofb/RgDUSHrKkV6XcNbfuhFoQMTa25iBu
72ScErZ4+lCzSpoy53251usXjCtt5+PaCjmqBNQQ7wMSd9Ijh3J9hUMNmP5vGYOj4QvlXaKPuHLR
h+dhyhy5Utcpje16/kdlQ0bbOtqtRs5UtzXY44fRo0qkUoj5l93UQXGp53qjMGMs2SaVK0y+0L/5
GTXDf0pq4NRmyC4i3GKgYvKXo2XUo2LLYgB5nvGk2hKUuLkosvCRpz8DK5WSFpP6PYcrTY2licw2
dpkWzWwKcfwKkDP+I94HNdRZTAAQLfXXrfNMbOQj8fzdbGR9XmhrAjhHdQjo5HjN+3Qfidv/eeZZ
ZV4ZOA6aNUOMAMIdLLreu6pwDqXvUea3cRmLbeKMUgW+yztojhL59nE6AKtHQ37bNNnjlLUgGEzr
DLZzL0eYCz4XNwWNzj5N3sutBw4CwbBOMBSzciMP6HTGOeaxl0ywV6u2vc6KNgdIu48vf3Z5qpmc
bAn9uWSmqasIMgJz0Vr4Trg6ofKZ5qXwxnliyIKNX4poKWWhE41lJgTotqNIDPeNS3j1/pbYuIMv
IYnzAhQS+94KjPMLz8NtbJ92sSkCjqY4sMCxYGdurHinRrIXIBjIX5bpnQ/j8fSGkVPGzx6JjRji
1d/x021IygB8G4q3FaBEtplW6EOVuv9Q/uBFVXuUkYEnCm9t259fWjPFRIe02ATr3P/FODLTbxlQ
zk6+fO3tg+/p148KGvPCXFW0eRu2eVotqEWTaMJiMxZWZGhCQtMWHBibyiBmYMjHoF+uQFTOouZd
DTTi+1++z+EhvKRJGo67nwVFrf9YP9vRg4hnBn18ad5n5fq0kEAW0jEV2sbbJIMzS1BthliCRp+W
QkEPZhg8uSf7bUYS1d07JSyOJ1tCxJbCVSrKzBIHhZ8z0HU466wrJbgx43orrUzN51AVan+0QXP0
t+R+KGeOtCIfmApRjV7MQO4mg0lJUxf3KmnwNd+QfPncjbmrAVZ75iIUPuqsEll6vKryUCnjrbyG
0bhZBCWI1Zie3LIxThzvYPAU3Bp/FhM/rEDHO54Zi5Gw2IGw+siRkPy53dqvhL5Oj5iuIndQRmhb
ZL4iV5dYDWHW09rOeZQFdMrn7ITuZdXefx+8yY/lv4UNWy5rhOSErw1myavWHiMhYTqRzkUygoDz
H+oMyXJoTrFsLjWxXb19RTHNF70PtL6k5a+It4prm39FoE4javP7LqNqaAT2JJdnnpHD9s4BWoxc
GQJS4V90Ro8zULsrBG1695SKyl8szP3iuKKY/lLNQvGC2BF1r+mWO3HKxqgNrmo1IOTW2bx0qjTM
7X3RXjz5Edsq4ByQuFvYNoAqFZHGGhGaTN5IEkEF90fpPMwRRaaq3gNIFIG8k6tKKEMIleMDuyGf
6DW+pWrYuG7Q+tajQftEoBF3eVvrYOsEAVxlLPFWWBsgORAxnNh+a7UwTr5gO4Js38sPtTcpnyM9
YvEyoZPqcAAPwNou1C6a8nCH6LQDP4lMzDdZdp5UGlfjcZu9bmSli+hXwqR5PYCsCLre7h6aTW+h
RIQSPllsQz69v7ReQKGIGjI538UfMPiszHATdZQsRv5VtvPMN8ULCR/w5PKW4ZrLituw9zbcP586
Djv9xtbBQ3jt/VkMfaYWVcayATkfimCppuqf1qfGLOVaCOqaiMDhyFVPWjfs5n3CySMVnN3iY5k8
xeUVa23s1rN4jW2aYNtrZUUt8t9hsmAKB/WpPrjS5HQjxoy1O+oGvHxJCjH10uhRCirzk8lA2Lg5
RYFmIVrBh9vJiB/xxKCjeKb79kNzKo+nIQaXlcEzbVLJQ8F5uAG8rlhRvNL5mr92zIdZIgqsp+fj
ah9Jf6mLCEHtjoKxm3QSimLL3K2hsgMbirFFhLAOabkQFX+s4ph3qcJa2UtXmbpsTVQnJDZF8c3U
Ch6tPfeED5nShgijTlcJ+Q8XMgqA0SleYqlmRAFTFykJlrDdSkIFBXqgSGMZpSauQG8mvL8nUV0t
ffJIeUYBnzivgGiG2FmR0W2i95vCY4fH4SLLhHGawa2gf0xXBINtKekjFY8JNdEJlWhXmPrDROIw
81n506GU/9rmZNutR0QEWn6bhfmDnxxv1Xn0qt62Fj8iIa4919ERvEd77UTUJ6ZeDIya9Cgl6azA
WnHCdHTsTA6AKK3sIrUTd0m26yAXa/doEuKhw6eYfhpu1zMkG6ee+WaWIxLszYBN2+rPjwpGuWZj
x7YVNMEG6HIRcUz4biG27PLCqVQUwjK7lTLw1z6P2SD0jT7wR/ZiAoD+7ALu+G+YTIkP+oB5VZX1
znW9AnhiGLBH0zVdUuaHIZFAfKOviBk4Uy3CFTPmCOBuKbBemRE8liiU+InEBS5stTEpOV3PM0HQ
COCOv8c8XMQP6lljD1JPMKirPTdHV+udOAIzEegPmjNFgzfAG8sQikEErpkeujC8VED/NCDdJI0g
6FuuhZCUIDb1WNp1kFQvEXYX6fcDoHPI1xlQSP3IMbMe6d8oqTgOTv1Ldhv9Vl3KakTDgimSX5sa
W1lMf3LAhK7PvanYyKul8JUlmOOns6XxCX4hbfKNydGTVVcdVqF+Mj6CEKwWjJ4EUd25tpakTgaS
2c7HIONZLrhg1cRY8f83Lt6ME4B/f50GFntJLicXCw5N+0MkOk9deG6Xmt2WmVSxDT3ZzO/lVbdY
uE+qU1kl9DVE67QGMCzIrpTwUnPQy36UFzNm1khM5ypYYD5RrxDJnKrQeM1f3D04Zssvs7iVSyEB
vBZ+9XhKccFyPs4bYLTTbvwKDF68kykJvFmqXIZxTmDKGU9rvdbAG4E50pbJMd5eXbuPt6kYx+Uf
4AiqXLXq9nNVCDVo8Uu0+PT0+1Sm4B7wcOW1QGCpppkDa9RAyUUccmfxAyaVg/QR0e68dwJBQ7RX
3cccKDxxwjyRftmmwHSAu59iiVE8tef6Lf2/Uuilspgt6JCjZQTKkr8p8hcombgrc6K5rbYMeyrE
FoqNzHZkhjdF8nDIU+lZAbZ+EiH1r6bU7uj0TP468xVLJpiXjyNJGHB+WpVbaPoa1cmHwigW8F9Y
LUuZo6GpYnmPDgeN1i54jQt/Jk4YXjicGmne2JCVMbudUrAaEIzk65NYShWxFkY5VSy8/+PGvetR
zYtCUNl9L8z2TUZtibEN3Sq2FrRV69AWY2v3Ssdy3x19CZHUK6eYTBoDHA8Y+JruQ5GAoASLihjf
PCa3LkjCRXAMr2h7xgSLEb1DPh8/L52ZOrlgoM1yMnY0vHj63/Zt8WrVn2Rxv0xc/A5VMrnZg1Qj
hDZuFkEXfBCylBoOLPDS3tjEyFdKymPE8DB7kACzQbcs9aiRhZn+wf5hHL+az9Y4UUBLJfZ5Ltce
zp/YFXIDFzLXpOQOD7BWqapNw/YMOAAeAgR+K89kGELv/4LVyTRatTNGIyNvL/B5J4UjocSH32SK
30PlXj77znHfWQf0jrEIUVvA3h/WR2q4ZOXh7RMn92ALXz13bW8nBchcLMo/WKRDu6r4tG8mu/Cb
ae8gCd0obzVOrXNd3mbYXto9I97nnz4o94wmQYy5+eKRkKD5JQZJunCaSkMoI8RJ5vNp44nYjU+5
Jk3FzrQQ6y6rJlSNLI87uUw0puqTm/HZPmppNmYnYJ25OaxPNHKxRNdTbI9rpKBzviGfU2XHVaXR
l2ZzhQ9YuizBaTt8WwzViBzSMAa2cGHLPvn7vifsxFG5hMwzanA5eJ8PT3mrVMk8sHmF0QlX5aGG
LXQkK8N3KHTChTDNdGZFDdrdYIGqjEPHSIRYDmc64Iu1bJRINguZGe/k5iVVCTf3q3ua3uXg+D3Y
a4l7iR3SoeK8YWFbWHqkvQov3HcZp9SRIDatJ5dXQTlhbtJngB7wgQQVGrBOzNXHNpXEyfsko8hY
TIV0YfwFhUBnZJymzpIqN+1HeNWJWCffGvLnMhXeSOD1tNvwDuq1rAGJ2D/5G8e+d8R62VuGwbZT
xXU8MvCUlx07faZevnh/pM+dSTP/UPyI185IHN7a2xca9/0QPMOH1zxA0NDf7sbKWGM5vUbkOdWk
TAzMJnAkSyersyCy6UH1cg5liHdzcVCC/eFSxb61vgKP+k9pTh7U/omQ5IFriYCLcfkO2cb/bRXR
eiSPXQVx+STsFUz9icv82kgFS7y/Ymj0OaSN/wDXaxtHLWPmb63hdc/TPuJRrcNyRPHSZSres2zr
X6Ece5VjGx18HuhtAuCXQaXzCH1PfYflxuzSm/Xd8sqTnqeZY753ScOJpAmphJLYiquvVKCytPx+
nMBTk4GjQdBvSmjQDSD3R9GmtGeIumit7/zR+QhSq65wC6MMSYMz/56IIgZJZO0gajphgnsxWLmA
Lz3BzDt4uuqPC2XaFRp+LTduC+r57N04P1U3eOMPL2hVqdX7t+S9He4vj2ZBKl0SWHjrEog7gUMA
gf3CPLSzx7eA7oL4Jbg7ivuS+WQxFYyIX0aJaFrMLHMKv+gVx7v4wkY7fIxwhFfZzMIfwA+ko+01
vaJekEx4R3ok1QdTBR4P4QmqO2dMxPCQI4GyV+K0fwcaJ2wL4lHR3vBvvoTeg2yXeI04+A6W5kyF
lDgCROFQGDRcU5WHZpNkrBvWSXw1Pz8TEIGsuoHk5KKN3lpx8Xjyb8IzSbqwuD4fxx39+Fer0Txh
C1cSforrU3DU7ZbuR5tMZ3rSXwWw7YvhPAcL3TPbVv5wUqNLFEA6KWTEBZLrlAMLi2Dx5hS0aapv
K21ucAa8mkGp9uMamYidn4aHhE98Hcapbw7a9z7AEIWdGYKUnKzqwhij0gVkn8m8/aN7lqnVnQOC
mpD6NVTMUxmLWDhMvP0Yak3qZkI9dCD8RQszqp7zwg6a2uOmeFzoCxmR+J/u7OxiOJpNSi3OsGFi
oRsvYc0xDn3b0SKIon+lnYaD2DVFrL2oXXiJ3/VXHRtENj0QRmuq1K1syXvvXWbQzIAxyKfDLJFc
6Mkt/HVbykgUXqb7E2GGYin6rKrH9qSv44pcde3UIqiztzWIuEvVjr3QFppy/lZl8DV3U91s+KbL
GZuCG8WgadaIUady9IyKKZtD2avntaM7xPK8LYtv70kzth0loFMNJpMSQJhslNQjxn3QplQUkSey
x4z+oaaSi9gfu9KJlrwnUq/wUej4oXr+vT8LRDj+6JQi/HRXNWT0qRNt9SG7WvZ1RqiW6XZYu8WJ
wteTyg95j1iD5JixDN1p6INhTy1OiQjFYKw2zCKOpFv7laSphS2fYkNEeIA37JrTSV1hn5RAnodV
utTxvlU0xbrG5LeNiebvTqCjsN7GM031mR2HQJCTsDEEj6Zkg/aQz6GvpFSdeUgPcMsSi/2qneD9
GKeYj7GY0PZJq0yU0ls124FDqWhWON+40evgXJy3Z8agWL7kagtynKdNW0DnohYRzlOPb/UmUmYZ
CgcWZXiIlhtH04OurZ8/2QDEvjNAOMnuKr9bCmw+0n6brH9naHcVaWmLHoINZxHlWIRjiwgy18hQ
kg7BP6ChkOPhR6X/klZCJauBx8x8hCu/Cmp0tbIUBfIRd85miLIH0kV4MUnhWdtC/8qrHK6y/kSX
2kCs7hn8tR3q1YXJXzOU4/X8xdQHqdnARh0epdqYa3J2zU+OoQ+TQKi04LT61/uRa7ia3K93nqHW
Fm4TV8NC5/r4lminyNWSegT2XJAfQKCtnz1SAKEdI3gq8Kg/lu5VvMK/xI8klA546DY+zqc13wgG
L4Wre7cxl7zrGbkQJyXLjmVLiG/RqPdqHLuijhWbK9YV+TtgPtjvKfmAlqv2ApFoq6DbqbITpNpr
d5IALlPNvjCvQZWlXj0XfUZirIIR4vWja93bYNIpjn8kcxHW8xpfQIvb8Uo8eeSpi47eNJ+6kfqA
YLJQfndUO/XhY+dOtavz5f3nXZ6eor27hpEL8mhj832PqcHhRfYYd1VqTDkv9mhCY8GTExVnGNhx
zkMaP4bdE/N5Xk2REPZfnysx4w4pcYuTC1p5Mj2LCtSHiw1ZFchWp0L4qDfaPe0zG3jVYaIeT0qa
Yj436oAZp/ZzaX7QvH4+dlj6TvZsQBuciXjlygQtusl8+45g/2JM0O1mdLWH+OswmeehpNj3XLym
l6VqvYL5QiXcEFp6nr47QlaZ0VjrvGYxdzXRUzFK3hf5kuJKzDfrIFW7Z3yFhEM/yw8FLBva+MFg
53Sua8JLz4SO69DLG6fS2FpOvW5pfQoxzYCDYKz9sxnJbX2jRlDdLdAwV164/gnGo8yEl7aJfmY7
k7Dw09ivq7scMPrBg1OfGkrZqh02E3YAD769ZUJMq5QQDG5ivvxD1Ga+pDTYDErmUIIMuRePWQzM
kmcYICyyNlXrGPlHHgs1CiSMv5B3xY+8vBTuIjCm0NMC05BwYl9pmzy43QCbCuxCRnmZDOfaeX7T
UGUM623xwD3lND71MtXF6+vzZCKo0fv0YJKvD0LJ8Hf9GwqQV6ALR57STes/IRWS4hWDHVoSmKD5
qnIjHX8bLgPCTG2iHYSVGPg0rOQTaaJdpzrkRP4wXK3bbuadhKYLP8reko5MTRBUeDD6baI5ymjz
gCu2INXNR4mAssoeQXX3c7ZxM09SkTZ2ScbeK8B6I5mP32tuWsteAwgN8MOWPoK09HLv33jFa6ee
OMqPzKvVBU9AXKp8gEAq5ZhFcsSd3FKVpFytlZcrTYS0sOKjYMfGJHyiKXUYq4N35qORgqSZrbGs
vhiDNAoZJTp8zs12uQNZS3OG1u6+TkILyxwp06f04Ypao9qWJ43cR3XhIk150vXKAVI5WN6pbs6j
pdfYhI1aWl1kHZut1EGBErZdKNVUk2+6Ds3jkMGiLSrKPXyE2AHNBhViC7XOXI8zjrZWDyRKlf6A
I84/fL7wfxfL1rIju9VOxI1zcpd2psnJsaU2i2lJoMEq/DRG/Mhn1EeDrjhFXCvbfLdakkzs0rfi
GabPBSfisjLzbCgGRYmGtszl4iyj+lmmnlvjV9KUTXazXAMs5a14oUumuDJS6U4tYQ+tqbqOBVVD
jfAIawVmksWCRoDIpOt4pUXQ0weTdnoHo0G4UHSokd7sRUVVDIkQyeJ1fa7Kusd/xxZnMogVHH8K
gHC9+Wq+wT/bNddrUsYCeJDl+F4rQANr5MQQyTeo1uCxmTMeKFG5C4K5zdSov8fLSDpJ96bwQe/R
ol0XFrzGyG3TaRTlJLhbv1+rWetscfCTCuKW/XmPkWiTke/tv1FFeKMuSl1fBbw7SfJEpf/Lrri0
NhUlMtXbuDlLB8sRkO+PJmlkgosJupbOr3zQqAXXOgMOscNSeeYUFh2NFql5RVCuVGobNhuXgEDU
LMEj4biW/0zRZcSUaDyPRLvdoK0nycSKdD5y+Yh7+gIkX+bs7pKJxd95aY5VN9dmqNmJtGW/AUB7
Jl1ZfVrpuaaoGsJf1Fcj5gRf9uWAdqqRxCRYxafRh7/0/BbwX6B7kOL3FOxArTKbKrJcdqQR0lKK
wUrqTnmyafYk2eAJlmSad30pY8D9Fqry+v1CSS1tjIhe5pPsNxVOVaG1XFpd45OAMydFiwgu9jmC
NEv50DKBWbCG3UpmDteSLGPFtuvVm58b7PMr/7QKOak5PTHaoi5Gfwl1dbMMf3+cbVanBIdpD5LK
epc38w+vg8HvOFA0WWWH2Rc4DYL5gx3Ge0hGkZ4IQe4q0I4/Q0lpLdpu1adN1+uy7BNYv/coG/JS
HMvEU9q4c/FrTuD3BXI1OgBlYcYxyffKN3+Ju8j3RKr3tSU0ImMDhKM07gpnTzcjmP5spI1vTBJs
D7Ak5M/Rjni1p+2ORPsdHN3kcUAS5kIckLZZXy0PIhFQNZJ+wdmqBOGf8f2ldwboklncO+dFmpng
jpl6abQU+d/v6NV4rHDrZFsYQdNY7P5YQXdDwVh4vIKlsCw3zYgQkf5dfehbHZca/Dk2Ij84PPvS
XdTzVIveib45/WQgJqAGYFDa+04XzgIFMGq9MYjMUvbmqg85GvHmbPnLqrMQBCFy3LMvm40Yi34i
5qA/Niqlu4y0Ad+tWTlxaUu1Z8jlBE47MrmCcsTYFaAJcPncXnUjpPJL7RNHpuDMHP319V6x2iKk
+v4rxvua1EXZIFaT9uIpO+Fymc1H8FLBiOp95uhXLvNdU315IB6GHv/DhPoeSDdCoSKjnnuQp2//
wDdca0qZr3bx5vXfvEOxxQsl7hDytWeaz6+D4j5ZGeZkiQa6wy8BHYX0pukKsvIdWKrZz/i/Kz5P
tmo8IZ875v1upDf5JCKlR/8Pp1pqy0Qg7euBWjQuTNafj20wAf+rZp15yyGQuW5KoRt5WMryN8Xu
Rp3EKRvIqLYdtBpJ03oiLHK7o/TsdpdiaMZGIvnSHqyjugkJZJzq2KOILsmn01uh2lGUfTCcyqva
YS2ojy4rL18t9cUgCh/oXhxq0bL30y8aPXw4P3CvK8kpqpsqgdJhVJNU46P+8sUIi9WlkWRZrCmV
rjC4JrjsAKHK2zk9B2Nb1UUwjnY+wMGpjdJ6Z44/m2gZ9qoFjJBvQ099eP3C+0TEio21noKfBFnB
vDi4YAr6lnocJmK8UqNDuCpkN/suCNCXnFxzPpQTQ6Yz7tG20I5YOy9JCobNU/V4UFpqxhKIJiM/
sciPR3BRICr5C1arAkdxQzahGGN2v+ZLgzsfX4ew/vpBq+fccaBxbS9bm1087dtpB+Tq1SnKAo6x
Kit4F+tg794wZsD98BVu6SWo5yNfhn+Q9zvul7lZikuW18OEi/HFHswZMO+rnvjWPbp5XOT7xMUL
sa1lwkr5L+GwvrIWhzN2ECrEF4aiuG4/JbHfYVr5wq9URoGqz8AtLkClWjgBGYs0lOvWOu5E02CI
SzTORiZytclj7yNuGS2K3FIro211AnLY9jDtBUvKeZaRtfNo7dmZqaOty2b8q116dgDubLJmXWeP
EpFhD2TH4p0kTvMgf30eD3EfaxQKeRqg2exKvSpKx+2du+ZUdxs1ohQl2Mk4eVWrlNsw1ORxBTRA
R4YMpjRQUxbw7Rrqr1simuO3AfsUexgmL6aABLZoRkWDfDj8t4/p9BuIZavY53/TFwRh2Bhe4i9A
ouQpgKU1DRHRARHpKDSeUtt0dxYuu6ev+ktLEan0jjhCCgYuUG3LPkIf5NttanYPrqnAZ0bXhDsS
0x/c2qXReSY9JLrqnhVDxRojd3WwkbQ78s4ITxj6iMgCekJss56DCmwn1mm6CnF7hfRcamLhQP/S
ONgVnPzSQoPLbJutKy1Ub3QP2z3Ge1QUeHEc9VIElyXckIatInyy0wlcDA6WsM9CV8axkEVDHhWD
RD2s1l4XdRKPNEdKO2aaex189BgJWCl41xgP+e1Yz3NmxIIDe4TuV0JAEG/f3aVjT8uz4g4sQjpW
KiGxbK/46LskAPY+VKu390o9vRibwnvgDPbfj7pgRzVqclvNNywoe9tcofv7gCoWvu67pH/V74d8
AJ58QWI8htQtGSE2AiZ71t6Nckf7Wjc8JZCYtAqxKnr6jvKNn8o17zX0d4xmaDspwpiQKjUlKAsk
vFU//XU+V4lL1Ip1xiRZL+152MPw5y8JpstMhhs94ukejMHXiIQKgxXDaC2RIv8nXU697kkebcBe
Xk/KL7Kn8Piopsmtxc8P/LOHB9wWQssuAt7v964hM/NOn9/bC0v3Cm4UN0N56aazM+sdpDcYZibq
RHIRnC9Nr8EAxjbaM/IvlKpHq7O9dUhulwwFia8YxMHC1NwP9Ywew0Uq/udWHF82iTGAs+4ezo97
AA7pf7/E1Q/vksHrs6TDMAFEnVHAQFK4PXrIprJ8PYk+p4enJqod+k6oraBbJO+BPguKb5ZUopq2
P6ukulWVjRrbVOcz+QiloI3K/j14xTjZxBOLHgjKF+i7eTYmB1zmiI0wabEs1IlpsqTWmoZKF4qu
aPMRp7EXra+uWNNBQRqeGkhMDJEXE9RJKI6KjRi/AzHji/iE4g0tLqkS7iSKQ2AoUQVXuKmA1h6d
8tdDFtP0lOJlq8BhorfaDWBoyO1wUJsh0ykFPREcCYLg6wnER2G7fct4p0qL09DeAxjW1JncAacY
2/+jE2eQzh1UlPEoWnB4Whv541SEJtlwwBN2zwkc+dLt23Hmhk8duYsPAQJqUV4xjTQNPWHtHCLH
iNdzedu1GhBPzlVXHnWCTr5iNIQ0UDhaUl1RyPgWsJJtw+yxszTvxlQOGs4F1Zm4QlhRnn8e3yur
JrPAUbnDCF6q7islOIcKecDgXWJBUjKAN4RkNHGJspUMPUo7lLjaHKhsoShHIlq0mz0yFvDIOtfW
DWh6p8sSCWjXkflnKZ2e7Iys6fEYmxDwMl1HVqqKpqEJHPrY3nPAE6nl5lHDa41XG9AWHPk2+oW9
wTgiRlUEvoGJ0NoeYw53AJX8OA97m4Qkdz0j3Qbo5XK9WC+BUxCpGiBorNatogfmYL6UfNvpoHPb
Ir9LwAeZoX58KhQect+luws9MnhAiKS4aBOWxnnDNy6MU9LOvlFNfBcKWOBsRCHfuMykFm7LvVHl
mUGnt7MVVtrabdBmUu5BeJ+UdcqeZvkIGUN4V2q+UT/4dW8kyXEwfM0nijk/ctdBor62MJjdOqy7
t7NgPKLJGm2hidoxXMJ73YiyyIsnlrdFsod/RnOQtrOXMkBsIPokBA7/gpl4+TrXsbl85VwMEh6H
fvtQJGCbQtlpVTix1y4krBDI+8a2NvQZMmsqd3tzywKK9FJx93yCTtwoU6pw8/PWNbPYpgsxAHGm
dhCeX4XZnUauo8k7/GAI6Zr2A2ngoVOax43EoPGPyN5d6+0nDxnXnYXf7biDECelHV8S/5k1wVIH
FBr1xU4DHV2t30NlSI5tl6hZjV2kLlXFm6VIeclrL4J9tDuJNY42tj+GpaEDAVgM2UTWOGzCdXuM
kEVSyINHWgSsumIUbvvF7uJDy7CjM5NEzprJyXNnn/WKm+d+FOqCVXJ0GPzV5vtvBLHTpQBpQf0M
E0EQnyBf0r5wBTAHV4s2rw4El76pkjIBJxQCiH8b+Wl1RvzRaBPkB7ZPbP+QLL75lanukmD+IWIS
mZfJTFIYTx6vyUiFENGgY9oMxkkrohyPEQakbdsF13rSR3le/s2ncotutPp2CKeDwiRlGWEEGaP8
NcBLBuIcDX5F7MuLx80OEZbkmy2fzkIW0QhIwJ+9r7yp4AV28RDwutcw58BU7GESXBVAoBhC6wTv
PzuZNdTAbfXpkD4YkkYClO45v6Bl4aarCetWOU27LXbI/q8+O0ZOlrDmNHzZNwLgr9ozj5k/2BTe
V3i9hBnqUkfbqlbpOQCMfSBu/QvVWRy4eu1+Z0lKsyiNlQ19nvAcAUdM8a7t767KkdVpDhY7NhrN
ykZ4J6hdDzZVkWaCm5GdteOEaU8Qd7j7mNigXHxlvfhCTYru13lodRAZ+mevPfmv0Znr9FVYEttT
ntw79zsbTNfosa151gmN0L/JquIMHI0mkvOtYyy5Ow0HMcJx4BJOM74/bA2YF6Ol1MCur7zMMZ5R
U1v8FVC66kHI77bbOu9D7Y03tLR6PHejRMopSMflO9DO8kvcGvvv+v1pGvfmc/6rcrpCkHaSTRAy
md+mzll3cjhYEnGh80zpq0IWf3I3xQn8Q/QLHWXNDUm4PZqdP2E1BeYCHlwIht4Qum9XFbKh3AnA
qsbAONSWgBDtfhCCsZKv0/L1Ova4PmEKXI2vNzJznQp+GGowZhREA55r9yJZgmFdntRzOXeXze4u
T5zSfZ3uCWuRkirzzwRaK9wrBMpEO0tAZWPT4Ti5+oudkJDnv8GIfE0RjwJdZL02vDKJZ8NyQIdF
PEegU6Y+G/CUfb2WZSnO7Lxhnwq0qKhHfB8z52YczsRSfrm7FMo4AwRV9Rq/Ali4J5p7UhEOkPP9
EfOo0F65L/iF9tKYnkP9tlOShWrr4xrEL/sSVy1Pq3siUZ0y9ccB8WGOwIgl0COHANj/xHmIQAQP
8WzpCUMgIo+3YUqCh2Adla2wyZmQL0/R3ZRDx5RDiiI3WaDG3zkEhO/e3PKHjT6GS4s9vFqNTuCR
HYCKoXy7YumAcr6immEuPY0pDH6upLkHYTa35jOnScgLw0TZMgowjrfwx8kxVj8aNwB1Dm1hP1Qt
c5NCGxNci3XofOXOyG7BfEqD3LDDrG1+Uq+3+4gEHbcbads+IwLCyna5Cx301ahyHm5IhyEcDiAe
i4IP7QlilpFk0Bb6XYjiovDeKp3WnVCyKJbdbgqhKLVlK5QEJ/69Nfto5tJe/eRps62BBmMezVuZ
JM5rfClssuaSP3ErO5qZZNa2T0/hvYdKhCaNVCvP0JW0Z5PLulEylqCzOzzXLt5pRGDXs8Jn93gB
qIsfaJm5h+kIdB4Cl7gy/9miZIZsdj1q46T6gQKd8aVQc4u8en3tjycaiZ96bKVaGu336H5fziIQ
rVz3ciE7R/f69hXyws+5+A9ZepOfJfVbmLB+MxE+67NKdZqx8/I2r1/kmqX+fgm0lK4aO4ErDWgs
olyFP7tlkoSUHfBqywGbbb4DVkbBoRsRjpxt7RXlFSKOPEwFokbAeXP451Ok4T9VbPzdXTTlWlhk
Gqhau7ooqZ6tbvF532OyUlRr/KBD7fW1/bnljYDwqv/VxLyChERPM3bd0r9itW6c9wpESoR0VEIc
HEchWCLWpSZSdksGQ5gzSYKoF/0wG2moEWF6LhN4IVHwH97IsBByicVu0Y2BKplnLNHLW0DbRaRH
CVkWkmItoqgdcwJuaB8XiISOllQzbRIaWxdWnU0anUoES8aTkGI3pWuaBrF1pQLPmviTzpkmQrA/
3Qnx9+YqiWRiUxL3HWcH2Ofut0XwajLCkrlk5B2/2XGg5xToviSxVEQXI6XfALmbvjYrxHAdU/4+
yy2eNuLz8TJTCUhS7bDeu8be+Wu6QltD5zHOnjI5dbg+Aq2sqFBSDel34ccd39qgBTsXV3ggx/Ok
8fFJkmx3t1vX8ltCSoZQFvBB671umt0piAhFAdJbnn1ov+8ttIUV2EW09Mns2q8icgah/GEex93Z
i5EQNCuwArSummhIEF3ZTR0YQsY7Ke01lV9RGplmNghCg8WYQJidwTHXc6o++G+0to1Q1b4xeSQ/
5ltOZ4r+e/5TeZSdEzg/fB1IqmJZ/UGQoWTDATbwmbxHeQ/eADNPHTVAowAXI16SmOIGD87EJNKl
LWH+ImwzWOYWR/2krQrPh4dcSOpMYs22ikhDID9jeoXMQydqeu/Tv25tn9J4hxEFDoVPtLGvrJ0h
zr21KgrwRCjNRQokKQ==
`protect end_protected

