

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
MpZqUX7RHqqBov6r9sp19cCgAmwWMQKz/kilwg6KfQHVNd7thNhiMjNr9jWB5lhCnXS2Dmq96KWe
V2+V1FG8hw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
eHZEt9aF2k9bUkzJgCuA+q4yfEhMdqCEDNKyWFDaQseZ/ofqbFQAQc2uVVXTRkEXQs+GrviVm+j7
2wxr0JrS1Xw60RqMKKhLpfqRVe2BmFAKgU2BRL0PnA5WtTOSGCOmSJGfPa08juK1otVgwc2Gzis9
06D0/bVknfjjRpJI8Po=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
s0TU3tsqHiK9WgquIx4poaAXQ17I+2l5Vqn12DnbEwMyPpn0YeINJkDaKFxRf41aPK1Wkun6v9Z/
YYZDqYBgVO9Z0NMkbD4LC5C9cZSBdk4ezqdUWACnMS4IR+6qI0nvPM6pNZernzgmYtMGFsG0h7AO
2CLMNIzANr+bYhHkAqpdx/KPtV7Deh8xOAkQeNSD+8rjhU0z6Gg+2FjdPjkTgWwsP8xrTSENuxiw
xPh+QM3dvd2tDQbC1sSMu3CzeLQh9mMzJ/R1uFQDv4VC1TFFFPI7VMPMlrl3y0ondyZNERO3SeHy
Mn6aVbKjlR68QJuFwdsz80LSh3ZTJ+foTk16ug==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
uIfIqnJL93Nk48nDUNvQ46MGSw+0jZe8QEp6D5vC3ytHCm6yvGspxOPTR0O/6R1kGtbYGX5AVD6b
KvoAJRDP7Wr2E6PTOWfFxWtEHCKiApDz7UksHM1gqF0d7SCMfsYR0KKn9LnLJiQxmEJD5y64ve5y
9s0qEeMi9k4HxMVPc9k=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
XH+fS8ngHwfDFxF50DT7MdOHeXbY/uKmg7Eva1j7eQ+2X+a34Rn17d34wKLf1Z56AIT4ksXzo17E
WT5KT9rKAQNao71yUm+YQAunOwqKEPRyxOz3bb+3Zvx3y9p+F7xTeZFLan3KtqwByX5rGkNJtGjN
oI8H+T5FEpTIirQ9oxghooMSVVhKX8RsayssyrgajR3SSX0Q0ggoCOy3XtjsFKfrcDNlt7iEsMAt
+8vV+volJUxGGSYbt9ATDx7fk+pYKVnFR1jV5fEpxyqiZQoGjkjsnbN29jqgiZBfhyEe2uAb7sF2
RnfrEGY96pFoR0k3gse3XEc9radVftI75N7ROg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5808)
`protect data_block
o48Vmq6HiOrthGArL5tu8rbTkF/elcQtYf8vVaVeRYQdjygQS6vmQAsheLRAM4cZEj0NNRyacV1B
+HmS3pfpIRnExoRlsdDk+w3E/nkJeQEd/EqfWXU98XC86zTBKZE7hbqavXiRITaIrmZp3N/WeQzH
zOiO/SdhvVp/d/IPm40T/Q3Lygfth8iL50r+51IS3LsLCYKiAl76EPpgctZ/yURPd9DcuyhgAmio
3sp11mZuw3cvKykhUi3EwNaG9ob4xaFg2kbk795fxEX0ix5oUHyraokUuOoPL7dr4AzpbGPqziaQ
CNmgfbylGFOD55y9dmrhnat7UWaGLDOPgRLp17Clu0dYRfZkiJMLY7FS6lP9/NFDMC/EeyNnIL4r
KV7fzL2OhFQU0pG8CqcF6CS9dE2Ep7txNKa5/U9c0gZtQkTdlXjdob0aa3PqPwImFkvoIYDDGkxD
LWt7PNu8EG5wQlr+MQ/OM3EaCMjL8pdtc5rLHlYcxl+OqPt7x8YBioIesE5YHuz0XaDlG/z4rFF6
ZOySU5/LnaAsXCsmgdNygb+K7kUpBrUdGkhO0lMvPJd2dUIV/DpnD+qUd2Yvt4Ofz2WeemeMfZ/R
IQe4+ruI5YhD2OhRacYovzNoi3bZEwRWLoYW48KI/OOQt/VTOIl+4ze7aoZ5TWBPF8PX6NIlAVq1
twWhA7MJHPIMc2wcStaUu8KkHL81NsbWRRi+0gsysWAeTJJsYABxXmXR5qzFNk/BbNwQS0qRL9ir
twORZyjJ1f951cmx8ly8IfRhYqagdCuEHrp592ABBkvmHyFwsf9O7dHefyK+XGFJqrgdQOeHRl1/
PywMFmH97P/5jRo3Ip2sJYJ8x4hCW/PIp46Ttzdxjl19igAZ5nmJVi2J4rUW5FD3fw4tntOmlz0A
QyXG63jKqLqmuHakY0tMjhlX0E8BJlRO7pqxyfSXHqxf0yRjvy1gBP/vH5o+V5OtIgnwTSXPnS25
HR9eOu2nARwOEQU/CJpqBY398FWhYYTnn4wlAyKypmNhfiJkq6PeFvi64jKtECrbwHKagNlJQlhX
QkZkHRT9qdKJWEwksBg5JmVi+uH5Kto471WSnN94w9WNNU8vjRZssDJE4AYNXyJ8cvezDZJ1ah/t
sNcoc1QEXDeq+oT7zRuWPTcmffnCPvuiB2YxHc3Daw5OUkt8/eEi/GBCXyVp4tlRe/YSvz/4huhm
z6Nu29wHFd0/ir2jeO4J37rVizdUwyEdSDxtgWklR20/GIqU/jf6Vc3oGStvyQpT08aWDqKnLylW
3LsC8EjT2MR1wZ6Dzwln3co2YZ0mGTM1Uulblfc2a107qabNgvHJXbgv3i3mfpluMN9Qpr2zOyBD
XHl6gC85643D5Uu4z+N7xNgFzdFglY7AC0Kd6CutCxA7n4l9PNA9GdauQv2s0yHMraMF6dZi30ZA
nwTRPnbQTv8tm2b0GZb3PzVsgNw4ojiv+ukSY0BIrBYh5mt3B0SWC+UpkaeoDeRNdB4QG+4lhr0v
JG6J9AIACNfUCiL5iFSUdBvguIddyVsIMSrRZlxnjgYuMr6WxoljR0VWZv3mGYmrjsOYf6roGnl9
nk0jA6ptH0M09SNqt6DNtUr2y6U2tPXR+uD0/CBybg62J0LfSL/WZZoT+OT0DlBdsstl+gFXRghP
HFcs169TqpAQ5lAwErWUKLA/QwMtDXGz/44vAjk5SbPvGfIAPRbssUGLTIxLJotNlhj17xq0d83y
QN0dsXM8doPZL/aRjgGMj4fJ2tc8cKQeQOIrypj1RK0madko9uEhyc8KeS5ZHjNTwQADxv1esbqS
vX6qeRo/bVCxJ5JCSedwPQsfJNjTVBSusxa6QW3kwybaQU9cCuu0pdcqGliN8P2F+RvevvC+UG+C
YmxCSg1A2PJsfcjs8b3uAVFf24MRfRLlD6TOWLs6VDcmyvfIVyi7a55Nivjnmd+ocUn0D/hLKV/w
rphQtwS5YskkvzbM5spkFd3JU9Nc+9qEkxEaablfT2MWN3H1LeEcWSuvy9JNFBrdkLfptAn4g8d7
59YBpkGnomLeoP+11ZfMRnzYJ8+T+vL7/Sp+LMKXYPtLylcy49tRlskc29E78CS4g2/rX5qExiqS
35ernt2Duvzy5q2da/Sa9MhVeZx8uiMWMrJ1QhjqSJYzXzGzJ5myCpprwCmmV9z3jTxbxxgB7yv9
HiNeYgnvzQDYbNJPGVhKd6ielK3axZUEXaCqmQLC70hB5RabPWxqRvmCnSmtUHmqXPeYnQLC8nG9
iE1HTkms7nErBme8Trn73nP8BCMXRRPSgrXpqhM5pvCMnuidTAVoyx879Q3h4EKXVmqAvWrRcfPy
IOsowqzw7PC4chSTowqQSnaMssJR89xeZkOk4jcZCdEZNC10T3Sr1EV2mMW0hWddOwuzCkCiKedM
Z6ZiYKrcknLvMT+XKVdVul89a8wvqrUSPT4zSO/1vFI4lGuSujXdi4S6ORV1zG+o6q3Iw9BSfNe/
/vo3w9wez9Q1ShREhcMvkyVD1gGZZp9VDAXoIZpcn4BESdEZXBpV07J5Rk0rd/JlCX97N5454nUT
JGUBMApVZJtJpNihtAbqjvjwpj7OHoNeRE9xqRx0nV0PqsosSdHFFzHZ7Z6VbO9cMlhFvR7sCbVa
vxvojn0UQNihkQLcCblYNmsYpkzJU4M5DAWtntKmDJeaYvCxfOBbHtpUUfkZ+MrmujfwFFXAJ8j0
TjTlSnXFvBkPTF0ltop5mFdrNy+cO/m7w0phN16lGDX0tRlXAsfTgVY44bAKbbUaREzPe5890jY9
j8qHFOf8hFgBNKxjxAVU4LW0exoM9vJhU0lqVaeqAxxwD7pUKjVPQHNS43+57aOTIsn3dTkdsy9/
3LrbSWocQazCarFlb0M3CNzEmi0DMTPzljNz0uwz1IZbuWevD/3KDz1zTM8tSC0XsGmq/R/XMN+t
RTfZiCq2C8hH0P4SvEzixLapgN8tTuQpD9pFj6ZLuQzzyBwT4vZF4ty/Rp27QephMcsHkophxJ94
lMk/7X23FTCouPJTCZN5oRnHtnKD9Vyg6WK2y5lSLOwfcr9dxBlGNdj08l6ae70UDNUEM4OKpHN0
sq1yAA6E9OFxSqPGi9VYIYGzr18jqlCGGPwXoJjNvDl9NGb/9RnRraGi3dgP9iJUukwjUuDc6aWY
bu4mHzFIasNx6D0OEmNKUCYjSnYuoIsx8zkxxoQb3DW1Xrx73bkbAKYSwiR8SjSn/m+Uo2VUTXMV
NGYB/lJXm9od/8hng40AC+0oL5vDMvJtbC/APFIzlJpniDf26vq2MsgZucFCnODjlh+rAJwM6uAb
8M5JOMJEomfjWKxiU2KHfNyRJ4NPQNMVfK630Guc4N7jIc1pU0X5EWAodrpiAQ7qEKo2b3e+k/fo
ASeY9yBSL0b3fW1tHAeXPUn6vQozLTLMRp04gQpD8hqKQ3oZBW21v0LqSDQ2ROBigS6lQZ3x598f
h5WOqGu2Gg72Y5NkbP+jRI0BwSDNROMF7TDMI3jYyf4efltzQ5LIgKuvLcj28Tg1YHArkE/7P3Qi
DAl4z+GBvX4HIcVRY+f6BPcrxyQMBEbU5XwbfgpEfU1xLAJkiQwPj5sJ0MsPZdg9q/20mUEJcpzu
8q9+FYLuQ0xoOAlafAekzT0lSnJecqPebQOuwoU4L37WUnFT6RFcWYCd+V71f9jFoc0KSZ5uzSHj
zUeQu0BAeQ5g5C9Tcm4wclO6jIVXk1l84PKVBqWatTuk9g20fGqjPLLpXoGWlbPRde0yRlAguJtm
ev4OcTAf9yDOX4hvPkf6ZhATfiaP1qEQansuvRc/UJZjzmH5xy0+o2bj6XlcFL7wewGSrZ3+grk1
R/bDNOC/9ZNhp57GMzJjK69X/BWAl04zqld2cY0oSSFGYbzmHDa9k4mFAD3UrwKqj7o4hY3VfnQ7
CL+ISyM15HuFojieNvbk6vCYj554sffDzwLndMtyYnGl/jZxxIunn8rBmZatwejxob8TlqLKvVOL
1no0VtXD20KZDApDOCxFQ/9G9e9Q8V5TbuhU/Mt+46gSxqkcqUYGMOPZTPKtIAlr9bSemAfnmEdS
JcVDelPt0OWkAkA+DFadSe34EJKGZW/6QatRmUD8pCJNtyuO7UYuEJ552J2pPMdSaO/0cZXrid2C
SEwFsiCTHXIeAhwSzDuEANC5x2I47QT68pyJe3QtTnj/plaZ/Aq/1URDid42GFoaSOTFb2+otuRl
kN20YTBaz4WFfmlGWjrHK6fwz2WfBLpT1GXt5e+fsSFOKaxeAmiYXMR6jG+7LLceNw4PzFBV2uF+
bBCNYnUK9K1MFq5/cbRIlJjfHYOEGsb82nS363Wag/mY3jiGvIqc8hO3tLtXNfw1unqCKW9Q9QGW
42k2NWA2fT73LH3whhQsu2On+Byhbtevl46lYqdDsaaIfvMFFzLvgXQpU/ShtAnTVfpW35cKlgUY
8SeD6T+dXwFguwaZiQplsRbq2ZZlboBD95PAtgBJgCd4qKusq3ONRzhoAzN16vhgRQh92Q8d4zbd
ZE1usTmMrqLvcf7TqJQ4cypNWf3PmvE4j/yYxjCOO5OsA4RQsISkcTw0Gkb1xcyqzpT9KN8M3d9n
sF+K0owfEWQYrfBqn7V/k5yZrz61xuhsW4+4wN7r4QIpTAuz3Rt5r4YYw2nHf/pkO6IHzumRSQn6
x4ljqHSDk5XfLPb0gIt4b0ATAAu1wgEoQmy+4g/9aO8DyHNq6GI7adHvtDOjbAdlD5ci0iGTRx7G
Nmobe1CNUlRMLgdYiq/RfBYla6ZJ3Y6xq1dtpTuoR+LL6/IpTvQE5I3Qexz2PBOF8v4s3QymozT7
6l+tAJ20U1+eU30cr0F75jiFx2873qDgYJPDjdULtBBQfzuofL8HBNAySFDY+edjmX2fvwtKNyjL
tkcqgsY+ielIk0o+GgXXtU/D61NYvDbRNiPqqrFwthoN4YjkT76nZQt+gszE8HUBbThDLDu7eqwQ
sQvQRqrSd/RzZWURKuuH4/Wph9rGDUQQG2+A+KFb+DpvV9wmeojRmw06k1+95tNEMhZWkAynxLvR
g04DMPgSfMIJYcJdzNwtcBN5HsiVxzyySeuCe83pppipHhX64Zm+u2HEIX6KTAkeOZdG7YlmMiMx
hMR/PIrJqBXbMNT7ErJWGB3XwTgV2DmruqD0JVp1OotnqdS7ghL2Q7Wo20YZrWE2XccUMRt9RQC5
YXX/js2+Yo6wPRmDZjbYyp6aA+4ucItjUgxYVHo9LXEeSOZj1r8IkgJbkJt2PaQ8800W1wVKQXTh
ixOyteLEtDc83ZRYV8DKe5Z/y2ZnXIxeMjFNHuemaeI1TNgH9ejGNm0vNzweeir+S6yrnYofWNK0
uoi9b1kmfB8dQkROleGI5DMUzNEcTrtPIeYjDpRvvBm/G87hQlcUSd6zRT23pHuydh0J+/hf9qD6
7fWDv/kkJsBKWoQHQL/dm/v6M677QviIL5mK/2dWQf0cvrcqgNPjtHbj5diIz82jhwgxtSqYnXYz
X2WOO0ubdd2Yp4yHEB5sqaLWH7/p2sR00nrvDAboCPXsEJAhJqRUrfoMh1ALr0KeCepGCqTeQEtf
f/lMU0bUyouStHfvmXzygyTYB1HyY5UnyCnlBdqGzypB5hX5Da69FjATY/64vXboiC/GOEbGFDun
H6cTooCLUk7Na9CP3nZSnL4MgYnK0VGdioxzcjnyK5bJmaoc7fcKrO8fGBO5/XlLUhxG/Ies/HYh
VV341wyt1NSreU/bR33+rzvIFCAUk+3RODHPngADal5g5gJ3Lc1L6J5nI0LFJcFUk0QXWZ2zSMVO
+muB7nbb1cyddiH5C+fT0Rdhj4zQVudxSpXEHyCQ7FDA1AMO2SsTefuI0KyMnbXhvoA2+PxHaRJh
Y7KHisem0HBNLiZFyQfNEMewo+wQK2LYixnQnuWlsrb8jf/EAQVGoGNdTzlJBuxB+oNBAYyruLJt
tuJS0Kb6XnSpArv9xM3CJ1Ft/4t4x48PqcaFiPkO4+t86/w9XzDtgUI6aU4zdp0gHAN4OkfkeuQn
YeaL+9Q1FeM9JyiyKygDE/U+sUZ2dJRHnYI8SQnzxWDjm0Zus/tFjSHXj+UU8/TXPjx8yitnQpKX
PFSNukCrglh4cp8v/2hgpuEhEqeK13lMq63JIAJPsy7NH7WcOfSm9Od0RyvFzXcH0oKfBdZOzjQt
T+iR7juOfUzkTdW6qcKdqSlWSAvx0+0HxaVhaqxEJx1FDKlSSR4BnH2n9SE5N3OiQTo5pZSX2/yo
J5biViZig972MU1gVHUJlQmjBHozqBQSX2sj/XGFy6qSclKOOr9/c3zW6efaBBfVvH07O40GZY7/
9jTEBDI4fcbBUerpXulWSAugDQpjw2IqLHVIg6n0zbM4fz9T6u6pV+I4KtjyE2gwV6uZzMWby43C
b05Khgy0ryS2rXfwb4f3sXyvIqukLHsU/H6iyIUh5WXjDqmmBXQS5ZqpxDsmlSrtXeWr/QSXF2UC
vw3mAMVTO9MZdCgpDtgrgALt8xmpN/TUkMPvUCj/70xyMDjzSqaEmasMmwNrJ32UtV4pHR/AwXSb
sml1OJTbYc35Yh3mIFDQnQUq5h2oS+VN6rthW9Qd2Wj9hKUX92T88EGO8iDfMGfSlSNL1IsiZtwc
OxMJRiZz9S4WLwLbSLrPwxDjy6oZMyyZpw2ZsmufcADopZhRadaeXv3v0oxpOJ0Dfk5427TlJtMR
vfSdCTKceYrdPw9FTmh/lt1QQU7xqxHfmxaSduZSC4bXRvflCERFRuyWkzJBXSHcmmPZprWVvnX2
cHFjSGtJG1xMwUcGb9cCIy7cr84T9RJ4FUXjHYDDVgNZOgxncXJUrNH6ZCe1wX/SGzqGrGOZNs9A
I03s4iQ8B1S3s3LypMaRTnlWlb/YmcJqBlds0sKdKwX8euMO+Bi7rwtj86W9L4Lh3MnxYEeUiuCT
zL3RbIeGCmu5ETLWKB452C/+vn323u8XoFhh0FslWQ79Ku8jFw9ZUpz/TsFCjyIt5DT4L3VM73KS
Cd4jH28mhB6Zv0X63nvBVTyHa8SKmkvckPkPIQu0j+WczGhEM+sAskJPrHIBnxsSt8Yk8VHneKtK
y6Vq0/4z2Va/jKpGTPkx1kX6MkZJO4SfBuzuD43O7BiXxjdHaeXp0m0Gk+P61IBAiBB1DD7BKf2V
vlY0K2C8KAlq1Y0yvW96q58V0M//0nFFu4peGXUfm+zRzB04aejTFA4B7f8SoANxmZct0Iv+4gOM
+swxzNI2cjlw/pha/J1C4inmlcssQwxHaE1mtTY/lr0rIv/EEcZb3xLgetDelJpp2FPeWPfps6KU
BXzAJslxahTUiq1Mb0XAx+ivj5Q6Eec/cmXFVWhAwfcpIHsxwpMlX8hyB4TMWULdHjN1sXSf55Pr
s++KZ5jRp30LEV+KG5E0lba22s5BR0zdMZXpyce+06zg1BDPuROIZJ8JWqQpV0TPPZeUFar31lmh
vWeIRNL38rcNbrDim6vCtY/F3dft8R58MsfhsmTXSvwEEM1BkdnrjWqs51bRt2ZobZOQOu92MHQE
gdvld9CBhJpeHUKy/vRBNHNRbrwkgwYvVgwihWAXXI87LH6gilJMUM2TkjCV2+kGkN2hNav3aYNF
h2vyw1JYKpWoTOfXQJvUp+VPRcvtUWWZa8YafObCOjrvySR/S9GJplobdIGXF5aNln9M
`protect end_protected

