

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
CWO2bSovBvQ2ByFi3vbGk64Kz9+OlU+ol4ZycfRhtc5mzW4spj2ZUNH57Z6TD/HWbssYOjRT+UqT
ip6xHZc7sA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
nB5KuhofnITTIpXOtfG8vxQ8BtQATMQkEP+DmIE09Znrcw3yJd8Ym9iSaEwPi49QFbQ4UCNnUF1p
Ci6v7CITkdmn7C29rKsxyl5fQwQ4Yg2Y9J8sH3IMncLyMWd/eC2FXu2c+nIyMZ2PxTUPVrUjVKNp
s7scT7Me3sAj5vk8vEk=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
MNNArzGZfZxohM+fQiY689sNLR2SVnrB6IH+/5sMb7hSfawQFJxphTI8Kro2JGGDqNxumEJLUYrG
7mZGSE03rCaVpdhD6Rm70zB4CVRXmxwbIpEK83cCm08nMbZ8k4fK0avkhJQjAW3CnUztsuq7IA0K
kdwznIXZSyXH6lPiqjIN2Skr4/LMpA0PrKFOFlQVuPkT5ZvNvxenTGhCq9p/EpzKYQA/Q64z1Pcv
8PTscPeWEIpmqBcuycpxO0kwVqiQNRqP/TotOuVFkjYLePFpvLupJo2vDdC4y5SiD3RT9wZvaSz2
Bb8UYdK03OxRsiXtjWytUX0MRrf53QlD+4mRvw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
JO39BJFIHsw8fi/kSg8TBE7CDuzx+VxY3tt2e34SSpwe1+CidGWrS2YpQSFw2o2o0JVA8lhp2pEl
VW+YDwewZ52gevHf/k4qIWqrG228k15Q2kpUAiHbcd1YG0RCacsRIqlWdSiw7wc/2b5Il9la2dZd
yyMNm5GMzs0PBGaInn8=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
DxfcLsCbVgOrlbX9FvTGJxwVAV0OB3tR+6ByNYT/Wivn1M9TCrq2dM/5FWlDqpdxHIYJfhQjjzlJ
F9cbuhfluBOxtIUuGdHg2uX5LqlRjgmnPZ6fbuzAGkBvSUoSqWJpXOKWx36bmV4iGY/0e23H2hgI
ZyfwOhBcKKufNk+Nq7xnSV7GWSBSiZWYhL47CEdCY+E8EYmyeXyXT8RcA9zqsfKsEZqdz1rU0vql
DdxwHxaE1OVS6MuW2h6qgK3l9I9LyDohZgyoP4VpBk/e9sTSLxcSmGiXwe6zlvuSw8MrBIn34Ezs
uAteiO0K8WEa+5P+7J56z0wy1dst9IfRzCpYUA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 45648)
`protect data_block
+0tZ36JmWJEIkmUZpYX/a0Afr0vSi+bOiL7MKNCv5+waO2CrmJ4Iuj0zHVqeyan51b2HqdmdsinX
FlGEU6wOOHKgjR/rID5cW2MvAZiesdp0Pit7/fMaNiLcQxNT5tnms0iP8xKeGhB3sN0XuDRKFS7Z
gex4Zuqv0kLnBU0GuhqaiFOvgYDv4J+o2U5niQDscKXvTGX5QApOvwPnInH7pkndm0Gi/Peel6i+
grkpZxYmpU/fWSxkskeEtlCEIlKjFPNeKCsogS1Sl7vcVZZET107A2kwh16kaQIZAw+64fJjJKAT
+3IGKiQsDlFClBsjl1Gm+bDCYxuiKn8zTV0dqsZs2C0/pZ7EgBjtclNe19z8ZBTCG3dPabjhIEFN
ntlZu9e5l8x13tsl2i0Jnh+UCnzWF2sp5+54eKy6w2fpkhs1+pZaMSX0D+8INQdzDSXh0kDCz8GJ
Z/YQiA0KhgntSKY8LUd6li1EbS9f9I7zc5pG6hurBGjD6EfqTg4bLYvDRlPze8faPJpnTYXSF8xu
/L3GhI3d16kIOWhAK3qVsWz/lDV7Jqtg9/qT7DEwpaSun7DdzJhssw28tFZ2xsNrFEw4dNdU7PP3
Ut1SUDSpH9r9KBNiKt+LGB3p0AU8x0CeWmcAAXaiF9OqW5wbHnAS3T/dz5L4pi2voadZ0OpYdjec
mnGoYqBIJSPRjeyIN32N8gGKOgOy8WUU+BaFHRAH3pkjemaJVrvh50wMAcG9AMO4Z9DobA7WBXwQ
gTWv5BXgiVmika4v6MPJyFgKeOa30BwPvbIs3jS3xZGAhiGRfgXFJuTF3e+0CoPCQ+F1WniuRG36
rMhQ9tRakOHqq10OMagHfhqMELmH1RlmktOuWgqnZRIqWsEkv1KMayEIjHRWx5jZaQpS6xt17OWW
c/mPw0j3pJLuTmxT5GBmdE/jaSXX+mZQzjc5fn1JLRYlkPV8WKwyKBfiWi1F/nwlSYsB+Kun0Mip
xd32BxRh95qikYMRt+Q+H6ubq4usOhIbSE769zAfWPck4W7RB2M4mg2ytRSRW+SwLJ6AwPYy5rVG
SLs6baRHljdh0n/bfU62QlATKZ5DcEigq3UXFLeUkwye2XJU5AaOavON2emg9uhQ7m9Xf3GDJOl9
y1M63SiCA+klWW53+yN1izgLw1+HKfiatvZDdDtOF3co6UvCEctHdHscy86584oUNnFEKXSncxd7
HqgDmFu48lgCg8XG8FGm4S1sZSGbV3lEK5lxMIQ9yUiP7MAlqXaAul1YpvQYSQc0/8V+Vl0pG8pt
FAHxMQfbhQKkjY3WkCzv59f1PxmZFuc/c/ArQw3eCsn+4lYJ5QdwURmgQrygZa32OPrVoZDs0i2H
ovP/ZEOzItF+javnjUUOpJNv9g/cyAm1m0LZ6hD67I00LqqR4u2rdyvqqOpw2xHLxfmeSl5VTFk5
l3yd5qQKTkTMdK2p6clprpk29rKNsQdZygLNOkWNGq/2Op31Ug0Fuf57unqhGFf7wU0/9zg3H0Rf
GHX9wU9IjOdRyToSTmDa1W7jXuvELA9X14wbaUDG2UedwrInt1iaPv89hert1GWx1NaATAngtSnA
Dn0fGkFlSBxvEP5Bqx/geQx5/wFu5e0ernH6R8cEpbktRnLsIEhR1oivL87b5BNVb33gxR1FRMJg
3i7XRh8Y7Zhx1NHzgkLIsyRmc/3QpS2z7sLmn67owFtEKT5eYWC6ypH+6t8E80sfX+8OBJWcWodN
Oa7d4HbVLVQpdS3WieacIpLwmg3kf/StGE7jFJA+QMbyZB4apMIjqzLp3ZpRqR1owOgIYHw5Kdt5
wiw/JrCNfbJ4+QmxSUi8B8rTTna1ONu9ZItwUNv9SBXKhHu5ifQEe/Gp3yIdLwmxsdQnJsB2Xj7y
VftwyrOWNpdHUKUh0rVMqyYNrXrFU5l5szxLQBDlvhjSzNkrP046bwdtcWKQJVWY2pYhXbXRCehA
9E2Tu88k0zNNllN29sVj4PcQXQx5LZPpYoDZMEFivVX7Fn19/4D2Cq5yOUztmcKey9FEGVdIrnEf
EbfHolN5VlPT2kvBJkVvDJEjZ6d4N8hE6ub/yoXXLbpdzTCaY9xxc9Rc+Zs2RxeVSig3PBQ82AmP
FAw3I5fjyLQTWU1ICLAn6o4oJzscKfYpkBHaNdiGwslKt+njUo7JeWS5wzRdfUIXNmWqY9nwNGl6
KBBnjJd9MimBfdmCZVyQXJTvi3zJebZ9zryZLIHRSd4IdrHd2/D2OTKDMMREkFkPvvxjvO8/YzX/
YPCHwa/dTkxTSLl6nCi9ymSTFJslS04crN23jwZiMAj1uX6VAKwaa92zNmrpCVTlyKiJzrM1d0vF
LNJjiDgciSvROnk2zCFw+X9fZSw2ibn31d2OBgVI2FNbJp+emvmDuC6mkRtNyKde0fwR3I0Tf5u6
jqN3elSY2PV8dKMsoRAXAp9S0DhvFsPR4Da1BrMbqKhwPkzpVOxUQqh8gUA7HgrmCMv7aHgZv09j
KOWwgmQISPmcnMd1wTSimo44caNHLioK3Br6bNcfGx/IVsHFV+DF/Sx0kjvJQ9bRiCn5kEcG/sd9
TCF6xlkfc3DiIosMjp3WwLKL7WW8e0AfztiJh3x2PyQg/zM36ymgaYdAjzenNmehlG57VHcOFanF
YvAnFQcOER4IEvWiqCuC1MICHP2SJDOdwu8NPCEyrh4FVwRRQfgJ0plNNJQwsq6WMUtYVAS7T2yj
kHxjMhNoFHQDmVnS6LUocUBXW/+U6I/Y6ziCdWSgK7haPMkFvqmsHC7UW+LJlfeiWSHJlmj8+Lrf
P8AqfrxOfyJEl0O8mbexU1KHh5tRco6fMRKriCGAbkOhjGkjxJsHL8PBRcVwwMRpMcDX2EnAQtvK
mQb3M10gbdyUUvILDyiGz/3OHAaeGRcFJr5MNexfwYR2e52hoM00Jo33DHvVNSb5Jr2R3I9ds2KE
cXGMXPBgK037PXHF2tHYuNXkSkbTLRi0cucbs5QsZb8h3XT7K2NbA9woifmtijZP1fcBYWq6JQ6L
bDeEMOHcbPbCpK+iszeOKVzIp4CcrIKh7wRH0nGXz/FWHufsQt6G7wzS4AkUQ1gDqm5MFd0OZO5f
S7VKID37/oC7Wrf/CMgOfvwJ4AymbB0+iREts16MfFmDu1fqO4tEzTv864elYTF+RJuZmS5HDO74
h94jG0ych7i1ScSSM15sPetq2pTJcM6O5r4aGcYwWdSXVf8MJWVT3OA6dANupfOvjkuZ99kRW9gm
dmXdZxUo+CRJnyT+joNWeamN0yEw0fFz2PmKrVmu6njQWdYftXxz6xAXGmWELUQOtZXpKNss+nq+
edfFtam0zg/tq6QtTFCds3tpJZo1J6cmmDOgvFfw+oxAPBbP9V6lzG7i5/JH5pd1waVK32IrXylP
tKRHeH8UNj70wKDeGX+OMIuj8v9cKiRyF8kEbZgRpKMA7z4SwLzsgcQZJv+kfVgtR5gxiTA5zPHO
BDBQ3vHP3mAEBA6ZJmXDWAcqpXeI5YU5LpxA9zkDmTJ8YCNGSog5/9d2nhWOJUJGK7R4uC2zRKjr
10VZteL1wDNMM0931XXpKSYG8aqY84+OU4I7V4irlNg66XJKgjxfy9bpWJ1ocQsUeWXayKqcu5Yx
mH7/ZaSPNee94TaneuSVL6PQw82CVfkGZnGVbFhQmIOHmlnLydo9XXXH5zvFU4t5e3Rzp/n8HxF8
i4fyU65ka5aM9pQoHMP2ih6+zX1QjD3IXU+Yepowpp5UTUsig+RcisovdSg1Cg/T81Bcb0n8Oq8C
5P2isBrzpwv1ByqFzHOFEuVQEIZJZjT85t9U6KHbWr3NjOwiw+k1bDIUDDvH+3H7+dFIcWfuVsA5
g5yRgV3o949XqjV2FXSnOHaeMYOSV6mpls3E3s1uxHrt0updnbDQF5Zs9Zk/N46d4OIb228jpuHj
TouPwYTUVysQlkYTsWJ75O+TJCsH+8Zg0ed//i9xcO3SSr93Eqrr2NjeSUQTvSiwLD92H2f/tRW9
gVPo25OBsVSGAYVvenB2ec89w9mpTkEL41MU3vzMR4+3NR6Xts49JM4JGFkoH6ry9YpPRxUZLtv+
fFtKrqrYD9FhYsVDhveb2REPHQDst6tVeCaxdYhpae41IfbmyTHUmg8M5E9ZICFwKQ3jURgUFJ7G
cfUzVa7hXsjeybs4ZfUjrPHWxqoK2p0Xj5LsvAE74FcPB4G59tm0T8sqaB81hbaWCISk+Og/CQ/S
rlXaQ8xEzlV4PfyW5pZvF5Q+s4rgg0u9OhTH91JegT15fVQ8w3kDadS1aRA14CjzY/Zrh8jkVGHN
+2QAsygaaZS4Pgfe/KmwjuDu/pt8SfdiHjd+qUzGbPjhO0v5a5ipAnDk6xV/0nrsncm8OjxYZSce
0D9rkIT7Ximu5bajz0/YCuFivx5syDnTTAzgJn0GlhQNHsgcgDzoJuJCTS5VgbtxnBieE1UvPu3R
IXUcbnu8K1YBRlu6JA5WdQMdVKha/xZHvk11Om8Wd+eqYcj6M3QEeLXE8wHMHc4RceFazu2P17uQ
qrwIREgb+vg/YVBbCL4g84QpkQDVnY8Z+VbLul9TQDZA1I2HFmI/mAkkSOPKMhFGprKye2VF+rYy
w0r4MUV8IiPQpEm0UvYYAhhy3J0pqEEnuRyHRuqk3OMo7GPmf7uAYRhHHbMty685U9NZNnTQfBWx
Uvky5nJcM+GQBLCJksjYuJlS+Q8Uh0QMP8CcopG7/x/gLLxg8cZmMFmVO+J70Bq7l4BAKJCxSgXp
7lIN1ZU5xKS0qPK+3zh+jBWy+I/a8D+vPOdCnTk5rb9AojdYmV6g9TbGKmUxFlf9GrKKwRcaKWHi
b7lCPZvaYQa3tmG7r1Ttxz9n3xR60O1yzkIm8Z4teevAi21EAEbtBKhMOv7iwq+rTdTIRsua+oKm
Wpr2+mDpGRycbpDXn0E57j6Ig7X2wg9hIxd5tuzoOBFSudSAxxxepk7GcyFXec0tQseBhtMoiQAJ
TWlOBoDShDaiCgp4j1bbTeazsK8ABzKM4mCAt1KbjdvH+kqG8TI1VFe0SrCL/hUNYrSgo1W8Nz5J
IYgxUxoam35YxEnqLG1xe7gUKHqZFl42u37TaAIkRcm3dl0EsGB+m/VsTUTP5gYw+7L8vNonBDdF
3eXsZq26LHKDsc2lNcnz/1oVc0fTXmSvtVlZaQgts1HTH9XF2Mf//Cu+jhDUL17FkHSPQUbVdoO0
herMHiPBKx2Ek64/N1mc+9jgCi4dx5ACBS/RdTpaKyuxiKJYLiDr+R3+OUv94B9W0VsZzy37fwe3
pta/gCf00R+5uE2MEy2t8zW2G1oNR8OFg2Y9+HPbkyN5w/kktRsumsvu2kZVmPA++26QLWEP25Yf
2t4I0lS0bx6+X003p2FL2vFcte6tgg9KAKSZ1K5tUJgCkx1estpagn+GdlErFp4i141tFoPVFxsn
PYiLTnOAOxUSv37iiTojsG1TQdDss9UtX6Tn0+2O27W7vC46OzLVTGSGfaCIZWre/RkYFwgesIoU
2e7D4RNtxrtA58UhCk4ygY3NpVvaJl1xyXuKQk7Ea4CbmaLbnYryhVaK/6BQ9FJIzQWhVWB+ZUn7
LkZ5oEFh8ro/Ic+gRLYbD1jGRReLyRMqYFxHZGJNeuakDPCZb4IVHExcOQ/LBJDyECC8nnrWP/2G
k/P7+bBEWIi4O3VbWSMxp2JcqfnLn7IaHSmfsnxbhK/gRjLwmwSsBso4PkHZdrzheI9Omu93j6f4
Zr9IlSRAfziBnYffDw3b/jiJiVu20O9JUFG59V8E/Rw/LEpwZ9ryIgo3oy+xTy/Bwhp5WVlZ+jA/
pYnOK91La4De92iHzsULPWGQHOAYVGkxf2Hg2dOildipwA2G9gvHRKyNCrmdktMuFp0iskWHoivy
2hRDobuCwgGsTmJpZicSdy0uQ17sdnJCnyNXBT62TFuiF8TNj2BV/3UGeww9yVpNnVKk16l2cQgP
iWLyqbfgHcoL9rxZeCm6/XzYCgZOUYF0YLlvJhtYan9o9GnIOHoq0PHQxmuJYLKl3vbhVcf0IF0s
AWw2wEt9KXC8q+q2t5mbGFczsNTJSsDFa0GTlrSUzShaG77A2FM6oNmBweZ8W7pnKfKZvzofda8t
xsvPht1TWchhsxSDFYWXbxfpeyDo0TjFI2aWihFnFwKGcwvxZU8g0VSb2qRBVRwATSbUbg7MziTt
ucUiYPcIDbtGfsQE4NcRZONVswLNSRf3O2r6ykLNXKybLMD/0jbdfFsSsZCNAkfd/CZyGKevxsjx
dIA1jCYW+IYqCWkKFSc4WDd+TB+48jLLjNRT9mnKyF8jS9LYzLO6XUTfrmX+y+uS8SeL8pR2V5ky
lu27Afce83RlX8zHoawvEwYnj+H1n3HcvYI5Ad+kZ2+QSl4u3aaK70uW/yVFhLcBkLQdW+8oxt7Y
tOyeW9EEJBMBscZzkj6K4INrHo9Jm/+lEtvPeVO6CpklULdTGfON2IRegUMklfNzQJyMpWhY+cls
3VOmaqTkiJrxbgYJ61f2E4Gwf59zZHCgN6LvmO6KYEeFyCxDhJD7KLRFE0lRNl/mI+yf38Z3BOxx
8okIbHvF3Kk77amAWZKhKuCyTdQ9abvy//BSkMwbfbIhiIw1O7ZqSwShPvz6k27LY8XRpM2rZ1Nn
H0QcW0XWbUbrZJwrM1JzFp5HtRt3p99NQ0GGcRDdKcMpNzhI3wm6/3R2SUvkwz1CXkMPGgT6L5iV
zU6/TOYUBX1FQZfPlEpW8FPFxcRKSB7ozxNu6j5dCUXxdsDHkA6veKuy9LdCzz/Zyid8rop51bwM
ZIsg3NNos1HQ9v9/4JaYw0T4915/t6qAcDz6uh7Cs7zli2t8Xi7qi1B04wOSWkxL4FENp4SGPN1T
K3rZu8v+2hVU8zJ2Dz3IGcpyYY3a1aF2/LmYzFnKD9tjdNuQi8jnTZ5ct2RloXkK0plowHI9OpCl
cqiX9xNeCMlPb5KibcE7CxxejX9nVCghiPXwIdM+rjdwLnW5ahHD2a1PyDDbriBHNmt8eZTTigoT
a3yyytTkGc94gpjTwO+qwVwsm2+NOJnBDOEy1bWNUnfo9oRbGhVQDpknLWYUB1B5F2l4SXjO4pM3
RITc4HB6tWtGidHeT6+IWUSsa2oYDizRjijAi1GezOZog5ZNN9qWNxHheFWzMB77rLlMKxj+Xhfk
A0vjJRUHyww4S7M/ztW5ms+1HtotEciU1cJeXWmfnIOb7gLvokBiqzeAoMjuptZqjwMQNo89i9o2
3Ln9tg9cjL4zg62W3s+Zsgz3iVL7rkJDFnyLGkGnNMyCqbgMG//XrUNwyYcyvrRQa787DKyMenyN
qQzU2K+m+ya1j1YSawAkqORZ0AjKOT1wsBpuHheaa7PgvwtKeHS3syrOt64T721pYMy7AGgpbNXL
xAbjN0jsDonZ4qcK2R6KXcOyR4nR7jd2tgaWkiL6+BmKQVpW4X9WCU6ARZwig4FHenjrr75j726w
O4FFyRzVyfc/62J3LFyYwp2AfpN/QHj33EuGB81LDpu7ZNnDY3rpn6J7C6VEHEv7YYjRC1+4zw5H
qq3lZXaxnzzCIzrHqqA0U/uuJN4cKnGLcwxodA56dXfH6KsT8XI5hnZxo7yntrqfErHeIPpRWW2r
urIKME4KKaEY8YS0ravm9KpWNtAARtdEz8EpD9hWosy0onkOKpf4gn8qm7ZZY0hJjiDaG4pxvwBf
bC8mexQsvnUWVoVnGEz/ICgFNgKA8mEcWaj6fuRwpVFWFW1ogZRtl2ordICQl9eK9wA8L4b9WQ6U
i9OLoP47jxI7uH08MpffiCBjFH/LFe2X8gPe7ubMP6UI/DMmiKAW/shA5lJzR10+ZhOpOtH6apCA
oSorjzrNsM+RtLIvBio9UysMOQZwh9QqJom53yz0PpEyIFKO2TbPKIcUMkb8WojpEO24LMoe0EQS
HIwoqjskvH6edRup6jC0ob6kqD0B/u1rQXLdYaEJb79LhUZUgSJZ8SPqndRRLiC02xadWPwQ3vq1
mBcAt/kiTcyL4eg3f6kKo4RoQtZTYH0mSiHql0LaRQp04Zi+hO2v16uzo/0qaW8YgCnOxqBZXQax
Mb3pon9ik8zpCxhMWQ8wOtessxK9+IpI6pBtS8HYcy6hX83Eamjr/PQH+EPy8ZwA8m/YET2KnhOF
KqLEJpIWWn9L8bPLdoCriW6oyQqPbz1L8Evny5RmtQNyNKuE9Yw9W4UXGANrtpNflQ883AEK3mKF
md8MBpvsTzcvOMsnieyt4XEfMIcGoxYALQJLy7RwsGFqj2ubO3aP39YYhRIMtj4NTmW56ScMX7Hk
5++QTRPmQxVlNWgH+Ysd359RYKsesijU6wTC1YYweUPHyxa/xfmBD0zkFqjGJ2uc7AtvCxWMQo9u
sEr2laB/ZStugZghI7Q9G/igvffoEsKE0zdJjYZtUW5TqyT9sj5Ee1V1VOKjo1O/YzEADYQzFU9M
fEzzTjSBX9mPqiZwqInWLE03LTkNeFhJgB4DhMLLQKZV4sXpUvgkHd7jIl5A7y3tZNA9IokTEAvX
84gIgxzQMoPmLhQsZXMFavfILbP8w6b0y6iTtgjJ0kONq4cDYCy4xWb7Ad0A95UYGEoKLWfgbRKc
hSv24nox6PTOe/28PsidoQBoZA5Qysw91CJ0tdwWR+/O0QvqvvB2nUqQip1TCsJiCzXA4NUE/qxt
BDmx/zIqQ17TfghWZIIO0z4F9Fx2nNK7Qb28jZiAURMFyDQ7MUmo/7szqpgYnoFWtTn98PKftiLF
S0qiGrhwRxbBxPWzh0j4tmNuA1mCs1IQB8GPZv5r6ChvGZGNTZ++6nCAoiAsX1+qSq/2t96sE+gi
fNosDSaEKRxsCdi8SLqFnjKA6wFPMniUuwi6vKFOTLycmCKf3hcuxqFiQBupo1u7RKKSE0STWX6+
MyMhOw4LGHvHv2y7hzwm0yzlTFT5uEyQIDORedrEhw9k7OywUH9eA9EtP4+GeTCR0Q09Q6Oh/CIw
GQZxilhS6ZPngszyHl+MOTRCRA0KJKBuHIMbMpUcXec07z6abw+p2JgKcEH07IHbpDTVhjj826qP
EkSKpJ59kx5ivbpFp6QSyJWhwIAkWzSGntpWOV/VHxl9osE5Ny1dO/7pNgXB6y5y9jK/AD9LQPPX
hqXTT0gxf1UKG73lge1cqMxr1zzvNWUFqOnuZW39bbD4Zren81Ol0V8kYEpaQCBIBMcEZgcxG9ug
5myjattTuSiNLrmFMe2UWQIWzSc3uv0+h2h8XAtrF6DA2HlPosRBXmAzc2q0WpZl3+D4Cqsuk4Qu
SufsRmFS253D4Lzsr1pQ0PQkozqDYfVLQHeoZQxy7hjwEL4OO5ukn2rxXhMRrje1C/RX1TEZrKTA
KdKb/VNGS45nZsjfnX2Trw57/XXaPddaxumTDdR/VlSn+oLcgneePW1Ntd/TqHOAOM0klTk3+6eb
7XOaXKBp2CBtPLzCYIAunR3mm1mRD9eS3bJ9YEpzu2UqIY5yOjPzq0B0/kwoUXdyfz1FmK/+QaDt
Is0U1tlhzBwANIuuXhBEx5/jJBKxdIn+tHkBlBfdCJ3lcXNiNR7eps7LtNIFiOy/3DzplQwycnn9
WjvPEvkwd1KEibsjbFXpHvPY8JCQh6ZmTU/dusikFABvzvQz3vFcWgUKzvZA928A9JrMauSDjsDo
38vcKA7te4vvrTJGgtBumptRxNvWbHMCRInHlpeWxsVZK6T8BviDaAWCT3O07XdSpNxzluoBJTew
LS67GvsE9TPFYJ3G/gTaJvIaH8KfcrpELhPBCMTyOxsKQjDetvnb3dk0i3w8oqfOu9j58SJA4DKB
nm+cnWj4w1nqerU1bhUPy3mFDnnLU3e8aOEfxoQMbVBxRBBCqqqfFju0IywWQePG4rpYYSk/HqgH
yKw/92r9T3WahAM+tt1I5/30rgH7QfCXFIj15Ch007056YSf4aZwCQD4jrI4Kok4kChr5IvIJRMn
RVKHDO8okK4NzPjnUWNjz1LZhvoeVP40kHneotYyjYqIv8eY/4GfDpMZARSz6zwFiGql41y5JLpg
yVkKm82WuxtQPWPCN1ZfOgLMnNR4z0+5Ha9eSPYrsuwzEOc8SrPmAE5nBta+Lz6DWQO9ZumIbKWA
k10KlLUoIvw/wOjDPpCtnLbSCqIk4mE9t6diHBqpEtXkjuq7owYtp5SDC8JwGxnhfNFGIflVYzXH
29aSwDfo+T26644PFTjWAQ48nwvWMjF30xv8B0TlkV6y3RBQtvRZbND6eQgQNJuZ8yyk1G8HdQGZ
Uf/2fJphNC9/dXYNO1N0nyy+W6uPhMS/Qx+5637J6mCmxeJ77dYnNOEYovixYvuJASKKvL1Ca3Ta
+wd+5f7LFh5+EuNfXgU8TneV763kY6bRKqyLxSa0eWs6mpDw2M5MNw/w+2tdHxzHTU8pbmVaf3NY
nz2ZOuqAQ5kU4WGwQVY5O2AMdNKJ038DkgJ8xcVn/O6ikHWHu0gRFhgr98hpO6s1xl2pI6FAjSgp
bwZUcX5e2vgcRwjjM/ESNWM2KlOfpynFWAIuA1oPOds0wMdMz08wwVTJGmkH2d5UiNNA51czrBxL
e2FwLov3sfw2Lei72iIQaIi8oH51Y2/KuG1GnffBdNKOQz1cNHAHbtDCTb4NIwf04Q4TK5gujP6N
c5RuXbTYFkj+S7Ghz9tekblQfCxDsxNaBMlIrvmgMl2uEePH/jqggaQTLm73O5O+QHhXICB3jD/1
UfKQ9LLZjvpXbh56+yxfvdRI0mI6Ep+mL0ZdkKIoRaxWWLvXDUUoydn/tTmYLJgNhtnHWYd6Uvf/
yYsYfmmw8IkjyqZ5YSU5qCHGATdW+4jcXwlt4k1zj1dU3YF7fgqH1zXgjrSeygbMkduYHiEd4ObG
O1ZeP5xkm5bVnJOvX9YVvjk8X/yayIDKJ6Zzyfggp2P0piqhrrQVjWuK/0wB2cYFjMZymrecKejX
V+xwalcOCyJ5IPb0WmecRERhnZmhNpySZknzzD/QP9w+cviJJEOD0bdLib3WBIa2fkyQbPa27Bl/
nl6bLhe3ModhLmndgOn4M3BLyUDiYVqkmftwrcdrV8Anq238RUeZppjQF0LmlT2dBlVA2A2KDLzd
FJzvVS+yAXy6q6AKE/oJSps/15+jlJ2Ek7yBkzzq3jECXQUFIoyhUPQ6m34jTYcbpZrpExO/2NJG
DKhJbJxhhjSMPqDrxiDKjSVyqfmOTypKutc1MaD6aeQ6DE34pRyejHxweR2AUIewg/ZJd+v7GOpY
fKnC/gIiDwgiqIDRQMyXzA63UbbP6K9VMWci0CU4r1oIJHRakWEyHVDGZmmmaddYDLFoTZlJZyAi
+6mO169WYlpzUSD25CqcN7lBIJnCBSsdMDTTDkyiJbFN1MexUMFSvODI9hJiFi/TCBL0L2PD09I3
Iw524+WH+aOosgxp1OG86VXCCKhhaqcJVGYzcAoAxB9ooOvmTfJTPgXl14eK3iiJ5gKU+srg34Gs
Rq7QzO4NZpza3+pdyjGg4VOxVdQSBRTDOBxRaEtb9XxqOg/CJobX2f1Qalw8HflTGfo29GuhMacd
YdaVvJSu4Qcedqn+e2Hj3BzWMymaJqEWIXQ8ODUlahnFpBQSqFV/jvI+K5k29QwujXWUg5E2ourQ
4jVaXuNxmeLPH4n3i6y/fE+I5WmqyyFWhUVcYiFZKoJMrpLpspMUBfcaBL8eiXp1s67E8fzBvfgC
K4w4mnpZoBicosu52esQqftTHue4ftCgzJO30ib+jHXyPcka+OjiEe6Y5EhYQLg9Q8y6aNClVNL0
92LI0IccpqUe4ZfEPTmos9SwCxYXAHRF9zNREYEg2mBGl9+/ZaDnqFPQNGUUUy4a80JAONaP0j0c
UoKICrYDKdLvBgZznh+SsvBjhjfYQ6kH6Q/FvWLswzfhztPWTvBzOdCqaQCk1TVF5nN7l+r1cOsf
LCUwAfciKL0vhzwngXmWsV+hVifAD3RnpzONOTaHyhNTi4TWbQi7+bDImLswrvoybUGuAUjliazm
CwKW+9J6eY2UqBcu0V+c1QNZOoNU2+VYAvlunZcFUVBxqDGAWuqZ0jed+OdYq07WyM8yhoPdxFOL
Lg5kywraTTAClUEqWYkvA8lNDX8MQiz7n81ti4uYFWp+fUy8bL5kn2SMCHHO2M78a2bXNUGRRUiP
Pc1fqTEOZhwUXJDd/GVQZlcL4vlcle41ec/khTWlw+VFzjm1fX+E+kZvMxZrD++JKNMPUhnSmur4
fXJeVCORrPJWgsRPI+MfSdFIk/G6i2X1omYhFhmgkWvMoqvWRZa8FmfJaDeX85/9PdcL+N94JXNr
wV5TCQcdq9LPvz+RUu7xlu4CHd7nrcb2Kr1fQmV4Jax7NglPmcN1x/z/ytdQ3ObHVRiiANn+ujoJ
SWyGylUrkTXBmqDzYCq8HdeJfloW6pUURFOty+TR61toJ2cP8pyGsJMTCgNtLQrYoocrlWH1tHlE
MOJ13Ei0pzYEchaMRcpT6czLXVtJdHWGYfbmQ0Emib5Sl1gjDU7ZX7S2CyGSKh2PSnxQ5G/S/9u/
8GgCaT5TF1J9gR2W9lIii6lL5qzlB3OKg7QvBmnsiTdJpPaXWrReX304JZrNA0CfsKiWGI7JkyJK
/NYlleHPpyTZJN+mdFofM9pFpVRseNnxvizdBz1nHgEOPCSpJn3hN80ir5M8lL7lbXsw8uuRhzNa
lt4BPqOnlqtdE1UANpMPcJnafkvi8DU43Get3UIkS+zda1zOIsw0ho5CwkZGBGRBsBta8bu8tsoF
tJYtODYCajnB6cXw67UA5Z+eLIqOPjSreovIrwEfAYPGStvwH0wAx6IHn7wJplyHkNCMyxAm/PTq
B+v/yiPgsvCl0lGmYvLMtc5ktCYwzhn0yoA/Vqa8odlqw6thM+i71sCtVecku9N7U7hD5K3e8jyU
TgbY0JVrWhnMJFN4XYZzZL4WRzd3uVRyT9n88RFnbiEkx3CE/WsCNo/ebuIuSRi/7gLMc+jQn2/L
KCRwyILg0ATdeE+MxCIM497gNM75ci3JKg5ufhiu1s0TnclQyGC9MzaiJ/s+gmGSAHEreoPvjZLQ
wfJTPjNIHQiqTiPNsfLRkUGHnT69bw8HvqOtY0IJoEUTDWfRWGb+xoyUTELyHQFv12mQH9EUaRT2
MPBFZcO7hGsSkLEi1yP6er+C44RUnorghgcdtDhRrgOV1Z2fZUnEbS+2hhWnUZaMaFA+JKLobhYC
JAkaWOG8oSOlH2yn9tH3YE9h3xJ2qShON1SfnMvWcmMF471s+lzck4pH94DDlOqXrd8AWYAChGVA
EdGqULbhToMBcvNS2x3O4DEM9VEWi35guizKwG7eTjVL9Li2YqtZYDkrZ24fFmTeArvBBSFSi5aN
KtVy6kFYV7Wy1Gh48OUZVWXFGpa+xvGUWpZMv46XTtine4LDEwK1KygMbq+6R3puVQmCaJ8+0Zho
VVpv+PLaImOIodqkAsRbBqJApG57+qOg/eose5dBCMeR7ywS6wYIWHL+dInY+oFseebG6HfmyxAu
1pAWP8yzP6I3AYi/NtEeOPx9P0w4E7Iq0MrqvmdKMjM+0tUKNOSlYwrfpindplAhMXgiEo/i6msb
fRTnXHvaKRmCEanX/rzfye0A6JhgF3fdjXjTXE8ciPpwdpARMBfz0/pQAs+XZfaKVY7as8ewSlEO
mJAeOFe+G71soGR1wT4l2TsGchi4MTpskKiM97CuMxtnjXO82HSQ9C6HDKcAnWDBdjRdYegJ1ENa
1Fqg3oP8RnOJ74bWvyBNvvES9nzNm2hWjYq5B2KgOPcjEOQ1o/77dInw3K+XJa18p97bm+Fe+anS
gPILM09axCtO7/4kGzDSnucA44v8n5yFKxOQTxkOnJEFcl0P98Ffs0iMZIiXdJMC4jfUTSh/3h7V
oImlKrJo3CItGJJcc1CWFqcJc8g9QTgTioJOTp8mKmC4pSEhecmDvcvB+IPydRpA93Nyh471bfF+
M//C9gOKwrIwKfLI9yyppIQB3dC2vANUKwkOPf8anUpT6+1mwToIYzPflJ++hE4HS7ndpV/1rXOD
2b0sBTDx+9SYpgZs6/GX8D6uadNU9GrWqNcvESJ/z4LggduxgcNNTR7ws4U2fZFQfgxWRVBZR5Lr
jAPQ//ydRUN1lmJzw80WRfnYCV7mTBPC6r+6ZsptzKjBSBKyfrpjj5MOaiSW5jLgmzpQvHjf+CQ/
Z3+sgDhF3t+nifyd1WenLoZ/zu7wteUDkERS0V4GQgj0TvlcQt5FybWiyc7gmNcC2dF0KKGNhVjB
q+OE2rfnYm9T4pzN1bLsAzZ7musk+ZMyhBTojfbtuW0OJoXcQJtf132rz4694zTyW4SERdZS/8uf
Is3Pfv7cLYC5Q6sQQl02il2UbVCKU2vgTDVkLbSu7Ve9TGRWM/BFaKWt+lsyi6xa+ymdiLzFo028
Sv5U1CXC2/eK8qDDalQfefRedsy3QxWe4Lcd5vDdIfmru5Akjxow9x6epI7mhxz9ZI9LymZ2eGM4
Rh2goZEv/LPGYDv1f+BOmbztT4Rb1DGYMercHKJ3on9REF9AxyuL+XDn0mxPd7EZEgIzZhEFKbZc
iyTe7sA/ep+XdxLkjvaMck/Oyy/2Pw+/miQDddRR9ssvluJRiR0rHyo7x2m7BF1dC/N8TjZ0XjbF
cWFqw1V47ynFMvSk2vK3EJwIbYRQEPLHnO0czwK5LuvbG9GboR4ncZ8KjenYAskm9uueX8311oXE
JM/JIckXTtp3rWpfcPyVe47PcoJ6H5nUMHHsz5fsKeLla8/OTSSoJieYonS0SHF0cyekM/fQvchH
5OnkgvgQEHmtMYQma09UGC/GkHu+7RcDwPLxhRg4uOdeAAmnHLjd6vkAGDIpU78otCu0rXgUwsNZ
Flu0pu6NrxKCsfbPLrxwzYd9wtLF3Qct6RQJH0mMMEWRoowR3rqaqrRp5P4dZHfUlhrb5ExdkE3x
0oKfm9dgskwjL9rOJmQvjITJVvSDzC9jDJzHZ4mxl29RPzETTkjAe7qe6WNJlqla+Nd7DnkxmPKs
8DN69t2XNj8pzX8t9uB1sLSDYrEe6ivaG5dlytZf5ovwmLYoYEyKmFyg4THau1SietVpSiQdLdzJ
jDhM/kV3OQ0cwO7Qx8nz1ycbjNNyaFGOEO58Qup4MuNPxBNM2L4j7CGQPEaQWO7xRvDPIRe+28Y7
y9rH/vZFNWbQ4Sv8SW/3xI4yIela3jnE32P+YuKDeku7qOdR+ryJ+Dleke5+EgUlqltKItTm1Gpv
XXNWPVwmw+e+EatNu774/OLPBScVhHzDq++mo1FFZDQRZFhCoHjd1OpT/FKsUcTykxWsbfrD+leG
jy034jkW2Zzt/6LNVf0AMSARPBMVHizzfArZ57cyrByptvJtyNPYfayhfLV4+kj/bF1veFPBWnFf
Fioybbqdt8wgrpg1n/9Z1CO86dSpdwNLsv/ks5xWrBVZpVLjxLTYUq/aYYmODFL9QQq0Zwp+WWYi
BK33p1mI95EQioe3xKdjPHvgLEibzJDG43zdWC7rFTme6k47qYJjHt9tEhjyqmGeKADLPnk1fozu
ghzFL9W7RdugGKZgPOw/ksRGGB0P5Wo0gwd0JE9ZsOPWw9WrhrTtnD3LCj1xSPMyNqQOyDZzv2w/
aXaj+4ytmWBPdu0Y7LN0V7jJhKnIlvf9/9Vrki1ksaM0Tek88VwU7gHrr3JqX5VXBylTLVLBLJLm
unDOglcJDM+YeQKkn+EpEpy3WFg25dEvJaQbgHS418H6PdqxEC7sZpkTBzYC3MvOnAoLbZyNy+UO
UZ5WyCVQg8XijuR41VwvZC6TH5Bh9MLRas0HCzMBECEttPspjDstUN09cKGROLN9826IIM1EgjJS
qp++tVDUSQhq5cLRInmMHYMWQVdEEE4SEhdxPQoeegVXDuCkA0j96QRwo5EFkZxDZWHMvr+T6aXF
aPInPAVrAWoMV47S0pLvOuRsdceFbuUapx8arcIz9JAPG1DAxJ4ZpVDfLZ9kec90Ozm8cqe1oo/l
4MoSRb+1G48TuiZRqGylY482t70T35PNpidh1fHS4iPk31Rtqmm2PiZhHX3jESvRLjSisY4yCuol
VzktJRryL3oNysinWQFO1j+LKL6v1dZwiTQLasZd04JqFrJ8Igxz1uS0rr1fj3r5zq2Wpvb9uBss
pnOOxUy0BKlIvzhNM6RUrd8gB09G1j2EJfY2sKY62fBIgXnJxPT4K530TNFB3xMb4wzZhPrV8h6L
WQSKGVd0Er1u84FRbtywEH3fHFx+06oHdqhhCAhV1RidlmqVx1/Hm2BJEP9HiNd7pqqRoNj2DcUT
EgQ+L3U9aurk4lKsCj950xAp6+XhnfVgXomNwoLwgh6c6fNXAM0PuiB0XHiD6A7Q7pOwuD1opQlC
U4kTgBwldzzk+WEri/tM2+llrsFbg9jxz9LVjDoJEjuFSJdukAz7/BKDBPIGov3zAd5bdQo22Wwq
4ohhv4cCG1YG6pMYwlLGUEU1Zc6V7VpfTchLjyAtnGiGBi9wdI3jXwqJnLpd4VxbmbSOTd1e6vG4
5JMKBKYplsGf6p62x+78JYvMiSA1nbkwJp/NRyrRk17BMRmOWxQYODJ/PDaezuQe23NyAVZukCUh
2u5NeluIhsKMi4Ea37YdbyChVo3+jdMKbW8YM5XgdRlUBtVUKMvLMa5taDyiN5CxbeCxLB4LQMGe
7UvPWEzcAz7g15YKnJE0mwG4553TzwFAW/7itk2C35qh/xWm3BwmXUy7FPaEZGfibg8TZLYf6EJb
NocxpXxeipP4KTwtOGwwW6MDsay2PhxtKGIguSTFopw23mp+3X1JHHO0axv7CbtxgxM3n2ODSV7u
f/q3TotcW1i2Y61Ynlpw9ZE5pyUW/iu78y9NcHBNRQStwNdm0ql6DiDnlVR576lmX+nrquuRdXxN
rDwkpESHQfzbf62ltHQNMWaWMTKHaFodfB2DbnpDwxfjhPcJN+h9QEb25USIZ5XHJ5dh4cy3C2ZO
S52xJ7KVUG1ohjf5PSwj0jYUXstN8wVX5yIGS12Zg0ksnE8gHRwLH2PmiUzkp2Bt5iswITknUZUT
yOkV+dblHflZUG0q+FPyDMUF3uDnwr3r/8lUBQ3TCfv82Wua6KceDx8qB9DHtm90UJHEZXmglYpc
DWRqWmEcTBbiICS2h0Pc01reKyfDO2XvJhfoaf4zDFUlruDpUiAKsFe8hd17ganIArRheY2QEf9k
8Frre75xgU5SuNGqV9QxAMTQ/JaFLHA2VA0ZgFDKmbjLYxAC9kkBcvbWQDJ+rhyWaAq4F/6Movov
ww2YKulqvv98cCGSb5RKmFK5E5XqvyZxdhiMaBtO6CcgfqmgluUHu9sAMG2Iphub9O/MsphVlsvn
/A/PoiqjEsnuFJnY1SoAU6K0oNdmA9APqcgo3t41LvZjKk/Xfegh/qmnQr8szS+v6dZHKQp/HSoY
ip1D0f29F/T89qQ8FnA9oYtgJq7hNi5NGuMvTTdZTB8CkkNE81xJrijR6yKgI9WLxjjniggeozta
ws72Ig6QmqKNhehqC96g7hc1/Ymmx8p2m6/a/R4kZKC92csptwi/VbEqr1ZDDNiSaccM3TbeN6Ez
w0OrofigFVvjVLh657kN9S6Jt6kWnzhKQsu6fx1/0FbuRm9uC9XyacvgfajvRXYz9HgwMq0AYOO3
guo0R+tWGiNXICw0kqLbK7sT9JxV4nbzmURjJkrufRbxuGEdYdYLfQgXyAUHcfhw0zugA4odtMxM
Wgfr664fU5IRkKW4g66OoZoHcJhgprnpRADa0dnyrnB0dJubdTqAfrk2q8TO0tsMNY8sePEW+Url
XloNBXepkikrY0ByQ1u8IuqztoBnrzCuwuw9ktxrH8/4N81HwYrWCaKzCsI5OjVJVUSVaolBHsbH
gXTcyvxW+3tso6l1LHXG1NWLILLDbjXF3CRC6DNd5cKbZ9Mvgc55HCC1CVeBdzmXX6eGvPPXusYV
Gqt7Jk5bVu0UTWOFupa6GiQgk1yZllaKqS8/8OR7quTYBj5uyeX2LhbCAGhz8lZKF+mLgb2iU+ZV
3Qb7QSQymvDqXIXZWlRm3oPCf+N+hj1KTfcGPkeGZsMcWyMiTMrv66wz4pZqbbm5UZrIz5Xkt6OY
Mtzcl+jLz5Ge/3UbxQ7+kNMefb2PVyEudIqBHuJ6YVyp4CRIoXKhC6CD1XF9qhxRCj0d8sRMnPkx
UFNoNO1HBw5Y+lSCrU2nuT3LKfHE9s3WfzJrAh/hlwiTayaCwJ3ycygsRYR0P1QqK9X5WmTvGms2
WZvBIltWBrDua+5FjjC1czYLvek7EHXLCsyXy/A9WEz1uVNBEaNP9EueoypghuvDw7RGVfuEa4n9
PxjkNy8RFQviGDmxv7h8Onr4kLKyyaGbaPYnlmozcF15L7VOa0D4nyEd0ehrywY1thWqVUxgo0hP
NQ2hlfee8E1WQHDhBX/uwGJu/KnSFCMnuWT86GXYry2hYDH2orLAUxvtixy5zEokwqZ/hzywZA1+
wYdCW9eS1ZhvrV+xesDYPI4lGdV9ZF3mAX8cJfR7gdZ/IfpG/IJaoVzypio5SLrB7e0tcLmCZiJv
/vsm60G/xugewvNWIlAgzhcKafOUVg47kTEQdDL+HuQnwP/SDkhY/RUl6sssMuKqlUl9p5+oNrxo
SdNTv6unUuhBdcVodNDxXUiPUJ8s1SS1t/hMGmbxWQFLViRlGE9w5Wf1NZ2VmYOquoWkjZopjcHj
quIWml2TEStOobLFjPy2HQ7i8Z3PavN5ggEkWibfYZJg9+bmuXdxV08D53UPNd9YYGeA3P6C6j3+
ypu6Miy3PJfgBhk2mT6ShWPUd9uYi2kqOfxNz+g2rTnqkEboGPImTRR/1Qqc5llrVm/6g6ZH1gYC
85KXBDIn8aOmj+0q87cEBPzRvlB6sK6QDODfEDJpOL+1kZoY3DaqfOs9XO+WnZpbvGfmQxZlgI33
uXrRg/6dJKwmTUcJSmO9dK+hUSAAA+l9v+sa0qxzRwycXeo4wptW3pbU9uRB+4pPOlth6ual4bbj
KI9pyFLKBmiJCGnuAO5vGD55CBYSimEBHHF7IzwyLzKv9W9iTdhcOwO7sUU+haAa1S8fnRqgjlft
Ihj2YMJAeoPRi1KEyf3LOYZ3cVuGhQbjxse+7quikvFPftNFubVbrNk+/9W+pOtmeBcbrsZvzizg
OuY0wTbKmP3voHo+4ln5uy/bjlojMPY3BM3Q26AdczPymmwjzrzQeFhokWOalyAhaNGFAn4o+J7k
4wlY+37wM4PfcCnttDjj8k9/eENTCUORZrDDeMco2yrwO7i64N4vD0VE/Ri1Ict1odBEsYJ04g9R
g+N/6EIx2FkCaOj8KxSpoTbhH9aJy9mHNqrIzGy1yd24FpI3sNhRQFjC3fxjP4Nx7t7iG4vTR7Zm
m5hzDIUDPsMAJMYeuMQ7YxK5QCP5o/PZXg1b2X7cWXxW8hI5sZK3DDRSfBPaj3poaabNdaxd7bbc
1MsPCHuvyB9OtbvAI2GuAoOiPmoP/czOlgWAmsZ+wYoaPnfZ+lU6DsgptHR8Unb/gXz4t9y1rPE9
2sShg4OxixBWdYCz4qYc7USBoHs/RLR6Xau8pzomNbiXEQmC83OHVfjchSyOdmdGTc1dxTHWXRzl
vhWq5ATmG/Xths+gEI1+bNDFjox7L9iGrO2S7zPbNi7FL4U8K74XiE5BOEpINOLS+wTqoNEGOPm8
TNISJtF7J/mChMCeh9XSlBjQ2F5pE07nblyY2Zqr9Du/sMp5hMp6buA927G475BI9xZu4OVgMqhH
LvVc0/ziM7yd6hVcv97Wg80+VHPmSjjkoJazlxKb3nZFrrpZHHM/wcHMFAO8Yo/X+KQfRO1S7gF7
tMErc419i0qVJhdozw+F7COxpesfklJI4lT7TOezLevNqtQ9bTFhc6bEN3dTgXXtB7eBYvQ8CsPl
+SgHBWUW0rGT8adHUFmGP6UQC7JcnbgfbB1M8HBMihjlWqbDvbMn/aYowVyx0Ky1i+oUaTijACrv
oqsgvJ5VE+WN8fetv35e+c3FdnT+5x+gF6H5UPup8/rMMBsQMCSZlp8PtrHJv/RTNvaHwAyIqeoj
QYGaxZ6lu8GjrbIxH8pSkV3N54D26972KYzwbMzY0+qG9Co7t6qN5qTlgDQ8SyuOhAvyE1eLlno5
uMdG+1fCyuYGxbdGbHZ1jxvUqUQ1cmdI5+vU9ClwlpgMXsasscVdVW/HXe88TDuVkG35SMyskfwT
akFPRJHVstgBMI4911LiFNMOe1aSuMPW8M1SQZ6KPYRlyIwH7A9Br3RDzvyYFLnZiJyd1OkC6ppG
svpSjNWgRWcq5wbu+Wf0ykKunzANroDJzQ6L38bz4P09Foscu70I8umd2UxYw4GT9b2z6XVQ6LaR
RoERwNSZ/AVvUcBOtTFGATTkgYk4B7NddB638qnzQFAcAhmxPjkSJQOmqIag8law95SjOKn7IhdZ
M1dcZShJ3GIokciVHIiHLdrE/Le4uIfwW/ivr7t51ouQ/+u08y1teqOyJtd8Qh7UXPmQCGjVYrk3
aPkqTP9ORHc8eGSZmIweM5Snn3MpZY+Kpxf88jzQtea9x5W7+peSO3/CFHUZ/vuHlvuNWzymB/Ph
Zzub2GAa+psUIqQ+Dmk+6tvgosyqim3+XExC3iwnA3ccpuz/h7VvkCW1UI4Ej0FMS1ygDB+Da7gt
V5EjaZXcDLNtaIKXpZ7yn5dWX18I5IpMfTOAP4hen8kFumzhGlQtJ+7ooTGSffusqNM6fqqafxqZ
bioQucSXuK7b20hVLBcRNnJzMzVin2qL5Zh6rkdNsl+n301YnM+Hc+kkXRijE9n3lSpFvpZ+AnYc
irzzhjQspFLQjjgwbIwajcuZO6g1aPpE7h0YjgI3bBKTFtmzoWDf+qn4VzCrbzlyzUuypR/1GS07
cYMCvYrPSZ5LuexhFArQphk8z63H/nsMqJ4bTzM7yxZCC1aHPZ3sDRDFC+Dme8hMLfXV4FYmwfYF
gvdtttfEKHqiX0EGukpq9qwO+/IThi36aBFRCTWywAKJmr8AHLApkEX5+16Bl6bD35lC45ZcHfq0
XnXxIk5gUdfAWXP8WGFw1Cpukdd6KWOT8R7Sb5+hQEN6OZhL4agaC5rPrgxeGkxGfKTGQ0yNWj1u
ij63e59NTzbwSDBaXusjgcyHVsUTi2HLW65Nfj6J2FD0VlcJYk42Mbh54OZs69kHHw9btwAKYH4f
unZwgtTosvUks1EOFjSdVf8K3Qz8dr99d4boqrQ8naLtHS1sxcgLPo4+dzpm+o+tZUS/qVa31v6a
opwJz0kbNz9j+3Sx+1+M3tm8YejNrfOObGUMcHJ16gYrcN71wbW3NBaUsEwWoeeC+ASALh9ZiIAu
XWbq4hR358/cfS1LGjZwOFq6Fcw9vEguyBcCv1nJRRtMtatoGvDzzwrNQrCH1U/3mvr3riPfhePC
duEmCDbPFL8/Lin22GO5QS8ek9tpV7G3nruoyBz48koLCgQHapr07gEeChDCFwKbSvXeNET3rK/j
ILCf8dzI+8E7qjzbc+7bpWm3vZC81qBMU5qE0sBQVx0fhzJCWYlt4hKBCXHH5azKTSmjhwFAqUDZ
73Fbf7nn5IantkYDcC8Jvw5snSp+qN5IXpNR/n2qFypqTSNfCCU69iRSW2k1JDYZp78Gkouy0211
k9OOSpumylF5RT4x5ktrUgSEWktFZgk+aB2j2mjLYnWxDfv8jRiTNCCW41F9MhilCrAcIie5BM9b
2OJLES3bDGOQnODer4m8SwX/6bKP8hXvrJ0ohcczvR1E78JH0mjYLNZGuscVqvzxm7TuBJ9l3ClK
1CkVixiFkW0wYoOOP6nX9nE2UiUx0kPbhjl0mHYu0CcBEPGO0E08e16uWl9/rAKjcfFqkbIRYMIB
fSLDFcVUciQQsXvEwpXY1Sy4yhS5TeTIVMgepNoogKJOIa4MTk4HPIqUPkqAi+O+/Xv+7SQRHduu
xRtGV30W3XDo0CXykBa28SVWhoADOncyZMfOKPBWtCSwGja/EdoWbIN0JfQN1NQMCrcO61OFhErL
N0M6ULAkqF6XMPbwNw7j9WWHTviWhb+OEJ8pLoJWoYfPVXN9RnYJ2UxoHk8AZV3MG1Hgvclo7dJv
U1cqbzy1gM7N4oiCxCLvgkri7M0x7+WedLxr+IhRDWi3fZgGuEbwFyCC848Irkhnpf+lAdwowplw
eKx+S42r/LjxY2CWQdt4o02/dHBtYxtTluUV+tDK+15TM9aHP4P+W9ObM640+Kl3p9tQW92jayiA
en0oK+aXUEdma049c33YDGAX9okfrEDg+SuLG2GeBlnvClR1ckrnhgi3e2xqCh4ZobK4vaKcf1if
UkcEe1iAZ2zWPCWVBbZ7vGc9p87IoVXelg3VrRQCgh10da7b71qJgm9K+VI+2wR+vNirOENl/oXh
xBQInRwDoElmWyPFe0pDKd0VTYAW2nieSmxDClxzAdG20eQMZzveEGFpIYCkcamB0bci02KCO1BT
2Jn9Pf5m2SH+7EwkgaK3QdjMueOejGiGKpHrIAkbaSaD6or0Iri/WY1hWqaJupwThOC8RoL0RWMv
jXCRU9ebvpj8qz336E5jYJR3uVPCwg2nG0GifGMmRefIJLDL+49qxzYrDQ2ZF74IlmHVkVOOuHIl
XId5x8Q+YarSI3alQr83ZvKNmDNvzqzWyV5pY8U6DeqoAorIl65SwNNtRs0r9nt4LUCCkBGsWTjL
a8/1JTro9HMcSXzjp1Q8xmWGdy6Y/8uvbK/rwRDBhoqWXgie7bcV67/lCbAey4xrjhbzCnd/t2h0
QYiC+DSR7dgzPYQoQ/pvP/HXa0E1+Pyd69pctuw+HjnsgUvjKBRhc/Eld8A1IFHt2yZakSyG2OvM
Whmn2TOow628/ubxYGgXw24AHKSZC3GSU15e11p5JXo3GuzMcqqrwRIj5afzxQxZMMIIfDUnMCzn
aj928LL2VBc1sJA9GrY+EbNwWvRXh/R00ULi5d5+5DvuhK2UQxqgxPfj4CkKGQ3YaG1q6D8iliDU
Kx/6StMAhtMFtJyEruVJfvs93L6eFF4QSzvDvP7oneXTWDOpi30QrxP61qXNJzqS0Fk01ZooRXUu
XO9GDNaE8VxNpyGDurjZCIomZIi2xwqYMSBcb6tIsxLErgqm54SXT7+sEMLrqsqysUbjoroYDrRa
QbkILoc2cL66mw74KwADr+ectAo+xr0TsPqDuWE9v8NuNQdXn/bJgkyvlFd1DIQfV9lNFqTFcumX
/yhH1+kO4m5jw5PQRQO4dwGjKAeYZA4Jgn61pWubIsTTXJD2qhi4leq1OwQ/gItjEk+L5N/OLChO
WfaIbDU0lJOzVpnDK8MkMi+/eK6bJPUs6IEpYC/QBdTHESUvkZY29eJDYTiYplt4E/CU/kOJueem
Jrk07ZFqMVenOexpZOoxEiwj7Uc+QxHHATodod4VCIlWMDssxgC4UAJW2QY22E5+loSISWEdnB8j
8K9wXWaCVJm2Hew+AF7B//2EnWK6NN35W3pRaNWgqoPZlqVV8ydcZUO5NtxmdDHbQUOyd+0/Cgex
MzhrT2PAzYjEpEVwGNy4Z+/OIi+yMSgK8Zy5jaNU7mTMQ/J19FjrmqY4s01p5EAzouCgvAIYz8xD
IPt7gu2HwftukSa93/bGrwE0472f/o731z8tphtZCc+FmpXkRPI6rPB5jXcyth6YtnNpTA+dW8vY
X9fF0JKInhgQV2J1cVneOZOtEn12cXf+y59yk6HbJv6llrvY6rszkLm+byRI7aQQtLW/FTJhEtQf
yWpEMeFPaDrmojejNElEzh1Wvyc7zGRMMZ1yJPi2sFP4Uk9rV04OPTdj1rLgk64eedX2vJQLVeF4
31hod85qwtoRl3kFDN5d6O2RaOL917xJFtrQh+HAADWZc0amdWkYVfNcdIp6HnzBFPqBm2i03XwF
//5w99r7syMuK0oCi28N64ET74bT5S0YVjmzp5bJ8s2h31V8kzOfQ9yVmf1mL6OMB7qQDSuuxqTS
Vhny94+DVx1d1hoFbpDc15KPa9DyyHyfViHr78W6MY90oxbnXASFIQtgumv9NQExS+rbBYFtbTqY
QM/ZTnnMqlOTpMo6FiGxt2NHUJP5lpUvKqQsiw8oapdOYkkKFGsK/Uv7p7rrplN0ac4OPXyaxcKd
OvVubTrj3J5aA7eWivM4he5ZFYyZ9fHoG46K7Y5pRIA4+sNrDmo5+pRtNUAgpnfZU+7fsj//as18
w5pNvHgdAJ6jHAMYb5cN/3knnyQdHamoVcbStqJqJk5PG6LB/wQgeC8gqFt5oKl2qEzFdEgcud1G
TMRe8ZTZzr0hFFxw/EbSk708/7lozum7YGhwWwF0TpBqrVq2wH0bjbVMcAAPmO4Iwh9+MPqXzyB5
WmL0baOI7h6alPndaavkRFIglCkDVFrHF181tc170jWSt6xU7LiqI7A/kRlhdqn4PL53lwefczwm
cMXfdyN9/JXijvwv7WpbLryKNqHxhNiFxL7LKXa+Jnpx/g3E89qUdW/SwwJqrSblBhFNQai1UrYb
x3JH/YWd+1dEtWk2bK7gbwF0fui6Kthy8VDPOgFfwfSmPVhF1H1Iqy9bACkyp0INPgFWiETcm1/k
tTcxTmnxOjZmKpe7Te78+j7u9u99XHE65Tc8S0yi1OTT5/ikTvKtkAoJjUCA4Am9T8CC7L7R+OOD
jdyhRZ8tkne1IEFHlIpp2W5xXh+iggcfjzi7uUADB/Azj7zC1tz/cEsMs0xSra88wue4s4TE9g/S
jDW71DpiETi2vwR0Vtmsq2UjxwYUCkcn7ZnadVSqV1w8ekAplLZUUZsdyw1ObqPy+L4z5MC4ScQu
Fm6AAuAI8LzBxmjfSBdzMDCBSbwYHYBmSQg10x5XYlAL2RO3dhtBAjgv1RRBSKQq2KkozM8xMg/L
/F63I3TjbO8ApJbNPxRlkmppOhBRLEy3i8KGV22el6c+cJbBOdI31NNy4sICflHkIcS9+OT3mSnb
7jkhx718oDK/r9lb1qAYSpwcRKMhfkLHBrOJHjthb1tcrjcCVYmlaI3D/FeLRaiHbKXg+Zxlsf7T
FBVYrMbDX11z6OjwoX+i4ZIxWyl94Nxskoic1X32SGEO5Q1LQn8G3FymXpYEIxEB0mb7AUBfXGxc
RrG8BII3DQo2kd2y9/esWkAFc7wXklLxLyX5wIlkkl/jq63yBCUQppNaZKiybSANeHEhr/Hlrdb9
0Yuf6WuuZvvuDe3tozRMv2VKmAR8Lh5MEVXS996G6533kSXoOqLk8ph7GYuaiGrcHDSeaVY2T7mg
IWvRpuY8pQ3fNjuuKcIvTUCdexwNAKVuEIJMflwcsDjMcWqXabo31hZhmbPAY4k5ZvGjiCuZgB/R
s+cGR2HsLRk5eIdYFA5LVubCJMsegZtHQ3sTMnE3j3lIL7xxOGTD6bwCG+MoaIjvGo+wwCByTldt
tdSx9EdB7//WxsyA8BjSRvO1PlxBRslZySSdSP9VybxGhORKryFb3p8lPRcTR9+keRECsS0OHNVr
cRSmO+VJ3NiXsBYLPL16j/rvu+1b1Pz0tMU7aYPuC/CZwTw3FRsjiX+Vj7enznk2ntjJdcosLuU2
fIkLdKD5s+0+Hy7BR1yvAbgrkwcBUaSVqzSe2IGX8w4Umz0Hq951Cak+C0zRllWu/ZJcduwOt+ip
Q9j9mXaZwJisU4IKFEOLdF5dKiqR1GYdjkCV1YRy6zYIcJrcC7wOGABkCwKa1BXFV9OdHdSm0QW7
0PttJLwk9FFHCYMMs5WuFxmMXntHx3Z6popZatTZMswazhok8B9kgpG5aPeDtNcjza6aMqI5xAwh
PDoHCN5vmMzWgM2RDZ76TPsCWtzbnmubQuIffRlWSjpInYQVaFmkHNA19sj2rwKwhP0PZvfKXICO
+RGWkUl2XYkhWKpA7sCOj7ukqI4M68kAaYjWVYnJ/GMJaBWH3Sl93+ZHFr7IB5whCkhZ7IcV5MRj
Dkz1NFQNy+6mhSIFplSWh2kgMSi+X3x1IEkxcGJNGU1UKIiXAUpfYAf6a2jD57lJU23VVUP4qACY
7DJYrDeAYUORutSJAjq6RDE+m57K26dyX4h2YmLWlBmDEHKT/VryH935vbBsaHOABeV2D+L/0w/N
Z2AadWbNF4e4OC+1dlDaaAgR8RXNqDoaG8eG319vh5HjHPva+0epVnw4AzikEvhFrWpBEUoEBweO
YqUlePCZ7V+rjhLrgeRJFBk632Mf8U9ht0kekXLmr5/3KrD9t7xRZAKYTBuauAirVXin0AUAHZVo
YBZmXdBjjRzN7lH+B5+CHMQD103HOOrGGGv7S2q7YBXBN9AGRTBj2oWeWESujl7YVNlvfhzQR+Hy
bjiCBuwaXw3BDyIB6XG1k7wZTpUMbjpePEIOpl5qDpHqT/Xyi+NA47R4uwjeGTr+GOGWOd0aNHPN
JqUBVSntgXroGWFB5IAfo8lUKM4oAfow0XW6ic1UVR3KzpBMoGNHQO0ZY8qvlWwx/ylGey2cwD24
/e6UChOcLvh3zw50ORhQmC64Fp1GjvZjLeoIdSLqMRNmsB90GDUeaQ+Cgc3yhjQbFLtWp4ssZsg6
AGp38D+XgPfum/C2yLbIqrN79I+SWRUo6qn/CVu4ev+TiEQyOTpwBu84qbzq8G58d7sdebLEFTWL
jkoMKmsrG5c81CjdC+LYppbFDzAKxvmJhLHlDeDMJTW2C/+HubSOVMmHtkdvhTWKBkZhxCMpQufE
Qdw2ofdwz8knTgw09bebeRk1vs8Kww4rZbPKSUO0yLmudhqTceMTQ80ksJ+OQVoKydktyrsLi03R
dD2WmfHy9cJEm0svhnyaRVKfLDEA/Mp70Xvcv0908JuZMUv5ypWXWw4Uy1l0uTRJjmZyjLdh8X76
51MZTHqft7HuIe2ORePYPmJQyfx69IoPKBuX3yiammU3EwKBfbq3IJ+zq68LXR3nLBx7u/Xb8GNK
7BdZtmM9Yviv+0lq9Jp5V4rfTAIwQwVf2urRcdPtrybhifO389zQV3ltHcG+g5CaSOH/bEYjGrc+
JQ5v1owGAVPN1pKQed4SYzD8vCX33ZPepH3dQG8/nAussu2X54+AC/uMoubJ0/HeFS0oO9j7bt6c
AdIyPxFvmaQ6RC7XYN8PqiAfyQz7nPuGz3kuCnN+P8M4WeYGQxHDm7kPeLXPP0d/lH/LKSqBB0h3
8XGkYBFkd5gjDF4aE9asdYmP4z7b4s9KX3fyGKxLQkZJpKtSjnGfZ/Fo6VVX+58r5yDNwgIreu5w
CS1aHmIALNp4a9hie/+r1vEVAKCuVQx+uXIJlq6+ss2WYqE4Dwf2/4n5aocXHQcqgN0p/hjQXQxQ
12Ay3wLOWr6V+Au0Dj1CM8yZO3cf3Vec/Elc3O5UBmhaQvaSRSn0xhjUn23xr8B7HWJ6eWfSK0IX
9UYJiIpo6CUk5URX8o4OWvgpEU7YNEh09In9AbCnuhoWRjxa+Lu6a3sRVJXcUX0AuXbiyJukMotc
1Vwvh0ey9if0h11mJX89A2WINRpq04mzFD3zOJxDSYRe0SxF9+2xk82LqQcOxNQBIFIoX+91/RwX
V1A6h9ZOMWotNz6nR10KLCX3+Pq2r8Nvlw/mEazN5S5u+L1zNWIFpOQnPwDbXIEB6VhEb2RvSIMp
sf7oIeCphxn3tWJUnx1BXtob5LElVyv49wmvWO+YxFedRLTD70Llk69y9BBCS09nT6M6eWg04Q2y
jhqj0aREQvQbf7sDUKLjhQwcuZSggEhKx41UDHwhNP47x9DpbDsoSH0nZfaajlTB1Uy4iVMVcCEV
YcMzSq5GJOshLisTaSbt4dnc59TEEqkf+xoykD0DXIL/EBMIXx828EARQNftg5+aQMw0jDEs5LwF
fks6XjJBDupLUMEeXviXYBIV3/qPa2ioiSODf3N4mwARHN5963XILuiYo8YqjZamq9DJt1KPJ+ZX
5oWnOg8KRc7nSbel9AQPUsu5lBHZPmjQDliM3GEQBxAS8H3yZayzAEdJuKsv638f9tNelxSpoFCD
K8dwjjmR90jXuAGZoL61Fwy1NP8glk/AoZTJz7vhOhK+yyVJDDJZnVzJZrEnSMZU4Rly+JyzmXtY
IzVLUoVvOB9iB6btcE9lD5QXaouh3USylxu4ZVDAk5OJrOT62sAPblOHxkxG6WJL6MWOobVoiSs8
pUH3fVBT42igcndWUwbTuBRW3b2dj6jcRT57hORtH/lc6fYConh4LSXOtDgU0fr8eW6/NxqKR2+S
J4+1CIcyiWXuP44tB6bdkPqAmRfI8rDPmuepVuqlNElghae6Vs02KNUwqEogz9yMqZCqWovtW5IH
nl29UTNvlSOr4YCZnSozasBAARDF7rB8+3zZc1J7/kfWXN0goM+OJM1xYwkziSO+qN2g1/7iPG4y
hq3iAIB5Icxbll1xdyjKHzsSN9GkaQYm6J3darwt+uLPaiCHHtAzXZc92B9tW4gAuPRPInkX1qrg
Qbe2++g6frP+OzMht9qTSo6UEi7gMfQwNeItU8mnh6lKY/tUjlQgCWGzTNPpmoBGYz/MTUvxFhTl
cKfFeEPNOMXAOGtlxaxxHj4kDljW9jytOqIQM3KWsMDhC+QJH23jUTEjmFDY0XyqddUb4tlaFW0D
QtRo4hZ2cGy4JSnOLLy9iMXRthp4Mgri/4YaPWFOU0gMjbilHYmQuvecDUFsqOhA99QqppxmKjrQ
u6SzNV2pxeEiL2aPSXCdDSTLLy4XefTp5I5zCtEGUUlvw7KeZlR/wK6EhZ/AYfqR/4IHfC/fYpGL
TG31uq3bglBEtF+aqKg2Vj9siuZ7IiRS8Ynqv2sZ48hzd5XMTBeSRYfeGx9bKSMiRBE8NA+Iy/MK
pVb2mquG2Hm8XLoqCLAdgzCRsIICY8LR3M4M0bgPDuaoEMY0KcXhKVguGH7COswQlgxhkax52Yc3
ttJ+k9KfsvVuku1kJZYeMBcsbt8OOxZazx+ovwvRgsQOVecSvpJm/VL7aTM0MGLkLSL2C80lPtDT
wLLSD+kCD5+j0MnZhgxyFl6vApAImhZ3KpAZhCEjfJFHlHFAE9GRZB+pxILq/TKIO1de/LdekqLV
7ez2g0opdLwpFAwzadNudSF/PdpQ9/yjmmaL9xgqQlyNG+FxtX88/rFqxkrPsSbJ2/FJvYHAhxSC
7WTwY63kHoIn/2JIhNi49Z3ic+hYKG25WU/Qq0RaABg6y/Li9jY0JvS2L/qY/y1gubTD0YT0Drbp
mi2nqTUB78sHn24yywvMwAyA+Cm7V+T/Z7EJnPQLev8katw+UzddBbk0W6ZneLuydS8RyVmHYv0e
9RadPo0VopizlX/Xp9yf/RQ+r9md3TxQ1UlKnQG5O6MoZRi0QkLzoEPiHWOcLLUZl3eGJC1boSB8
MyxPSrh1rjLVawv5/oFOD2asG+FO2e2aBzR1p/kDPbbBUbLTxw/H2W74n/SYPSzKjD5/xyxgzcve
2PD9ZjS6+wSylfsxcDxTr9CFAx1ECVr4mut70rCCqsWq8dXM7l+SPJIR/x5MVdEvcR9i15Kjdemu
HAUP4EuoWg7CHS4/jPiNErNsjp3i1tV+vP2LKFuOhcGT/84vuCu5zSK4EnAhv7VlMlUUCgDc6mVm
JRzkUmp3vf7BMyBP/uCXHRiQ8bBpkLsVwH1l3PsZwGqP7dgLuE6xiMxM6nAXkSK0vdgPZBiaKWi0
ul8P2tJgMrx6DYIvotpQ7x07C60pkZOgo2lwF8QcSPAn9XDWSqAj599uFMYDFZ6W+AL4BLu5KYh7
/B+IPP52WGsdM0fEj5Qah0Vt5tTxJqBWFM7OnZ/UCzW8fqRwWabi6z6bjzyzFhn5GK86q7xY7BVt
F9bkzGYDuEyD/T2jxfTTSOdRdTTKy8WycAxaEXZ+qhK4avqBmkAGJLmz4pLK1Xr67uvoqi0Liipe
dSrmskUiMzJxzwqqxji3L90srfGFJmBtER/pAACU67NOn/yEHTtr//YaWsmW3mVi2u8niFDuPuIF
1bX2YFm/hl48Gkw/SORuk42Rk3E67ZsHohwXuCW7GMlSTdQUNcX8FL2ZjCktharO/tdg4/JvyvqD
S9tsEgNYFVJwLR4gIDs69u3YdALr3/RJjvHH6V56lTjI90DaMvml9ANx+aM3yNPNFWABMvbGjOsY
VL8nJOPG8iSYqt4YlKOqGXy7RacadDUDKXMnhCqntVWF0Xs5EwjkIqUFgHv6cBZNlNJ+izG1Pmdi
YJwS/uvaaAALYfzWy7z0f8eWFEAsfNEd71Nr/Lxc6z6CaGjeksThojpd8I131yThiJeTQH4W+4im
WpefJU7oiwWy6Ahxj5KdMjQ3fsf3hl/DsSwv+yuKSVSMCuQxWPHQpJbSy7QsmuGkguCktOBqhw9T
jRkrESXvw/ZJf1+eqeqDdediMb8zwSs3RLvff0XZ+iw2gNRxp0Bgg/JuYDkIFWoBh0Y3rHdrFu0l
iBzOJA/5+ZWvGy0rW4JqujJ3WeDj77XiFoOLglAXxfKxpry5pVySZYvOqg1WIUzPUh+JnGAURMuC
dIOj2yLj/2MisuBCWUJAW+mv1IfBfIFOTHbFSOPLzjLMc2c2e//u9ZHm/oOwQ/DnOkI39rqN5cRN
U1Z7YbPVR5C+KGw282KIbIMO/3+hgOUHvF9ap/dbfJx6S3RUWpnr3jXWQFqETWPBuNX3Ng+jXc5X
K6RfKJjmvkf50/ZLu9CCAQrD5v2CgxgyKOcECYvOd51zKdaJm9nEE00/TxF9XIoIWzI8MoRvVNTO
uDBr0v4neuXv9MsXoSuVAbBzN85b8zRe8n80yURbjP0iKNBwnW1CfIQzzcf2DAvnLBboMQ+T1j6a
S87bzdjODOF0LEOUOLmuHCGDC+QKFFp+eyxs/g4z2jgWqD4KlPTG/uskDi5WnMjR/7c1SSYum7pH
m8G4wga55QLk+rQoLIHo1M8/mpLlDGNfDytyi79t5lXyPAU9w71v5Uk9MRIzv0KBGFYmNKNsZuZB
H1vZGp/2YwcZhLFz4xmVCy11pUVfVdcVcsAiwS3EF1FMERLOLYGsY3sZCBbwzB6JnbOYT/OM/mQ6
zv0zHpqQIVsHdxlAZL/MD+WRNUXsOhJXvLb9EnfxTPEJSYM7QOdyT9igPSx0mQhVACyacDljWJma
VSuCuRzkCHMWUhLyt6l5h2ZA7+75yCH/Zdysq6wdvKpJiL05AMDEF6rqo/A/TqpWtjDTPFMa7i3k
u+rDVcVoyVINxIXvTmhSYqvyWoHn4MCoWXvOFBZ31Zs/nAFGm/1+gEt4ivIE1tct3oJDmBhHqahi
1euqFkCQcw/1LC/14sLADJknswboSBOlopZqhWKNarDly8474ihQWiWPSGkejY8CEd3pbnULCWdU
ron6qoYRokhaBnKXMOIS1CNs1a1hGozeb+V6S54+2MrzOJ436b3WLIWBdqQdRyqUXYh/8q9OgmCj
iyivQkpXLy7xmN+HGqI/kK86EKvsHAFVe88YQz4GpWzM9A2f5Jz95zT2xgFYb9jsX4ovxW+jXSma
/Bn7dccbwvUtrU6+A96bhgdZvZBjq521TIU2vAqMLhstAXvP/ide/ug3m9zx+/GpJX+D5wjY2ZRD
Ujyhp4wc/B8/qAOpATWPPoNNwqZmzGWkoN09IiWCBndXH82aTmt0Snm8UHWIhH7IyfvWmjDUtnMr
+okZo5aU41TFe8EBuPogM32WuK1BTZW8DAr/YmHhiFxOQbnFUFokLe3BSw2cI2SJKkdpmBDtXjIv
egX5gkizVGpn8dh/WnaYgwYd3pjwHndpRkln3XymR2JnW/qNrvGGAqXomjb206jJXmIa6ZrEh7g3
DIacdCH0PJrbAFbkcE+gKpdr1KkBroEe8SHA8Fb1REAd/hE1MRDg7RViGoBEm5V5WamAoqEjfisI
Dt7hTMKOrwVzD3y+qPgBkXY8w2EVvk4dDXHOCOWWQEy110tQAEy3ZmlYHVkx4hI5FpuyDSPhrEp2
Y4YQgWozsvoplgD2kx5s8rGFxakSH9pkAkjGlngu1Dt37awREraJMGFISuhE4s3uclXddZFsNrKb
fSxVFOH+gXSoTkD6GikwAeA2KHGoflnalGdI9LVJgwyCTasGPXgEgm+KB2HzXD9hAdfm9U2pYXgD
LGJuID1ha+EP3074NHXgoq+eHc4ldX9y+IZS6aJ2bnkixzJJ5u9ggNcU9dqXNZPry9jPAHebklbU
nriUg5IPQCu5ROcFpkgdnAom6tAbM3S2jOkKuOkMwF79Sg/0Md/Zy523QIvxaVpcMyGFJEIK7jhk
ALm7NAEcwa/l+WWsP4eJz9FS7YvHth+CFvxnapBNfjskxKuK/coTmpf9IrumBwVn250/Ru9xkzf2
hGBBD5L8gT8zvVP1DGENhEdqzni7tpl6bkQSTHNjoHP5T9lES438pX3Ixdfab6fygZeQKgjzn8s8
tv3DMkkdmc3h7lyBFBwkaxE0Mkpd55zZpLSO2L4hNTEgptwfJoH9l8l1E1E1WFOkf6weXCrL1hXA
BHrghDPtTLy79+3CkDzTcRigjHXEKo6MxI5KG+mgqAwQi371VBhn/f2FkyLRo8LhXOEKqXdX2h9y
CVFCiLjcqtjdoD2EC6D5JEp1G34po32Zna03fnn3ExeSk83cAOoLbV4wJLyUPS+K78YisB/TdOIz
SrkCgbkwp/lyeFRqdAXdupMnj1gP6whFk9PbEqECoV3jV47GeT+HGzY4w3ipTf3yCY53FpY2CInU
T4uuo362KjxwFWtyuAyT8VG1L36DGBKsPyeBNUwRSnu+2tzRm5G6CtX4hAUywz4R9WY/2RXBK6x8
3iG8ZEHgMRYRK1L0WaSt/C2Vm4+0Le4oU8BoXMTJGZ0UaZ38H6OrPHZe8WnKctdEWw4TJPEZbE6U
J/zSNQn1MCKkuMJGXqBwALR4CzEOle6AuVdyrzI66G3tDZ+oCOxiEE0xrJ2e1CMd/mk0sJ2FtS7F
rM05K636QO42pO8MtZFoxGiUAzeGFEJB/OXlupQFrrRvGhQzcVF5t+f+0RXLRgvJwNRttoCIqRwq
sTj5GGTY5i4kWLE/9xNwbKEbsu39tI9Ax19F6CNNOF5qo5p9yge97cIFEJnHM2Ag+VqOvVXXXg89
AujKUHSn5or5wSznp4I8H07uat/xnj1zyBeTOK7DU1HHGJqAacBriM4YR+xZ0QT6nEBAundvjqs/
PtAkCLrO4sh4F8N5OmtU4+2Q+bxDgo6nh2VZTOhGIG0ZX6tD8KPijCLCE5KEuOU0lIFTPdrz/Xk4
anYXOOwD1DsZSJSjiiH9DlOY/RFqMwZWI5F9cDgwA4dU4vJZ+Q39lJ5QXNJy9ZyduDq4CBzKtyiu
gB2bfQ1OKZh1Z90v8qmhYHXkBAxQZ9M2L++/3JG5hXahfBFIYnijK6VS/uwq/TksJ70XTO2zm+JW
vJom+yes3TE+dwux4O3WbGRUis7mitb/zmzuGoaYXblwW3xFcJxLhJnMdumSSkaazRIfDsU4Sa/4
5UORcPEnXoKN75TgaLY25nSarThzqLKZjS2S/Du9a6AtQ/PmCvoZRwzi7IAXTnldnlIfjzwBCR+s
pEjI58xUqP9HYZm4LJ+c0LMvdr0nZzsMZgEUwaexisF6KIX5PRWV/Bazc5+h2aT5XTpEZvr4piX4
WvKTW2Gckd1uIj3vWHdCD5eLRY0HUueYFZ7Qs+GxNkr7e/7xly98eREtl97bTyTaVkodZKHAXJxx
1W74N0WYpJSNK0amctKIsUbnRR7XTq5b1V66T5SSe0ITKf8+lLW9XHlnnO4fIq+QW6hBwPsN31RR
cslFzq9zuecEglNw5Sohq8xRk4nY++zKUO7l49wO1szlX1oPUsrN3/OIwZUfeHUQtR+rLIdkBm6N
pV14YEBZ+68jEnnd5wNhyHRIXpqGMzpXd4Oocouhg2gjSE8DsqAMhzpoP0xwhQBTHXClrqoFU8Cg
e6IODjZGedid975681ZvAw0ZM3GXIf4QfnPvLk9LGwObgWU/QkAAEqBE2j7BLnRGhADCT/9cXh1u
h4cjRZLSZdWCRsV0F2PgB7u26Iq0OmChpicYDhZ2fIguHocQ1f5HNlocGIXQlk8AcWHv+rmBgWuq
UHpuJ7ueIk72/KnHhd3fxdzFhAb+0IdS0JBSxr+YkdPfcvsTJmLDQHG4fzhsP2LK8Mmvn6BY3gKS
uxJHbp14YofRHi2jBODLGVg2b3+hU4PGOpiK2yjXhzR+a5gtmc3B9heq/mGl+oqpvComtB6J00RW
9dwxkw7uXnxaepBDuzawD6fBkTj019B740uKzBW0bKGUZxPUhAfeGEGuEwjkmNh8HD4277FV22rM
2fK+bzB41a7+HZAiJTNxAWRRjqnC7/WOX3OxwnbTqYThw64wLVC7UIYmvcOKdeWOL0BjTFk1qLUl
GF3LEHWFXye4L3s+iDGHDDNv8qSy+eF7D78vGdCsPuPR7BA1iPYkw/FxrSe1RqqUQsslOXJE7GOV
6I+4+ZyzBijRf2j2w4NWXpBdEvAmWMC2drZE3Z4NrdUTv3T+A62LFUMQh2GMpW7UiR+852hjodta
B/cr0PxuIx4XyUSbKbhrja1bS9LLMqmKLneEpanFfgUmvA2yuFWdBYjmnx9DjGAW6zIegkhwJvRK
plTMwvTqDmqKnr6F1NO8Y2r6rySShEHVhBhPrHK4AUyptJIghofI8XkHLTdbeI9cI/ehW8kTd9mc
1AAAsHXZwGWNuYH//EgEcoeDXLbzKprKVBcI4h59w7NChYcUSKLQ2c60Iorn5CLTnYkG7dgG+u/S
xjsVGLVdWawbsQXSomNjyIzj2NBEo1VtXPrhCjBBn9rqV7eIGNkIdZFtMtpITf6SYz/zgry10SQG
orW1W3QDUA4kSvTDqAXFvuN5DQNOIVk/yrgl3CdLqdbVkmzLpurG6opGkbvOMW/vbyFEwWpDB1sM
PD82h6sWNPyBQqkgGn5CR39PHjcdBvRjhSDwAe4zKz29dYmRppL/efaTMY67hPwwIbpdkTpwWALC
rB3hDec4UIvFdRH84DDlgoVDWyc3+VT80Glcxihyu9jMfVpY7DA2/KHtV/6TfGam7g2eJfwhejz2
4yNwOzMPtHjOtDCBIWKb1IesPQKf8LLHOT8ZZKojgqsaS1QVph0Wel+obUWYhIWCh4Jn5nRI8IBg
hYIjgipVZchthXb0fEYMEwKmZP6f2yCzIm2QDj5IGHye/BZ9z4OVnj1Y7ZKNUwVsOTqN2HRu8A3Z
EkBPftke4otK1ejz860yYko19nUx+GnzCGvE7xA6v4dELjDtYHevQpW6OpMa4b83wVNz7lUGmF9+
O44NqirBMV/pyupY00MCuu7r2F8mImomPdWsFwGgMtN+0CjvAF0xSiPGjCpeEA8MW32EvgTVUoG+
NGu86PIcfE1Gs7i2LJoW9ubh4lxHslHwOM7il2WONTIS1oTjXsVkVJ96osafcQiKrLmJTdGzVl3P
Xo80N6Tx69Jys8vpyxL+cC7f8GDYcJlZi0KFZWnTwWGK8P05sPjuMPxOVu/KJpgTSrFa/DOKf2mv
x6q8SV44S46ZTqq8m2qA9AuKxV7mKJ3PVm0uqs+2oRUI7gfH8NaL0NMi2oe5PFh/bMbnC1Q0YmX4
Kvgsr4uno9hmlOX8qoAa38p0bQgjXktcTOQ9g0A9PV5qMP4KCpWIgvHcBEut7EbxYuR6vEa2Q434
kbwP2pXfbsPnDZfPDcMGjVJevGwdMnfRR/YeOIHMmk10eAfrsZTn2Iy01h3vMd1jhBdyYGS3YfEI
VaRjSGhCwCoEgJ7hBt6xtcHsLliSyk1prQM1DLa+/cgCFQe1iUF2NS2gm200SZpjaH++E8/Ri3pm
ulUo4PhExlJrGmGvspi21Ld+1GEFY2i1QVtRUJKKH8qaOJdXCgyR8ll+dkynU+8+8URiFlXa2Rsl
IyvW5BdsUXQK14jDV9gMX0Mhh3WPx2jj9Bcih4w7g7gE0jXokRQbemmpyN8gmoJUF9yEEbw+b29G
AHqGEdEO/ZB/35wpmEovjakU4la8jFxqMRAD2bWIyPGycCtgHxnJj+9aVG9EKtLmN3xBkSD/FkKr
cv4klntbAV0vXnQExhkqv/qUKMK592M1dCGXd4DSWP1K7ywJVP6ubHwt2t1P92R1c787J6Jqka7O
7gCqK93x5G5oZI3Gwxrs0y+JxJJBMu++hv9AlXZPFV6eXYPgMVOvkNUMGpA0y7TwUmsHBySTWZet
3VunDEvkjKNUg5qAT0wWd8tlMc/rgXgooDQ21J9nYmv+s7zWjyUUEdleibvVcHUjWORkP//X1UCk
c0gjuRcUesiNe28NTdPKWMGWGuBQsVFVnKB8O+/42E4y5UGObG48G9QADalJNs+Le6A+cH2pIyg6
vUfHBTOe6m0oB9XCSvMitVOJ5xyaS22n9b4QOLWNvAYAYkSDaNHRWAYVVZjrajNF7TeiH7LRjUu2
stSKX01qjXHz2TZuP0gN8SXctw2bZwwmqTaStCkG4vnvwiKSr0LFmU1zDyZIfjrr1wDrMbcwnVLY
oulmwJeKNZunt6ccgHafDofEccGMN9yuNHd1DskrT05nGvBUNW30rCaUaLIss7IM/nZU7cxHP9oH
ZpxEldsWFXyHctWwtpsdQkGQtXt+AkUVTdqx7PAliWJ7EmjWTYbRExmBNe782/1w3sPGqfPaW0uw
Waf1WLxQPTQWff8hbt2gs1y0OgpK3OVJiJQoZWUOzE/T7cT7oL37PQSXjvvgfEp+OSbvUQFvrSJs
6DJy7XghWlbh2xYJh9k28WZIeUy+jyvjIlK5f3Yk46pSWectwtm50J/+QbkfSwk2y+nz2BheaCEk
7hv9WwJ2MU39QA51azNTahZLAno86399d61QCkjgauk0EgHctsSOBc8Y16OBB906js0Oy2B1RNvf
eXoZVrj4vy5vPaPEWybL5vj4VmHHRoJe0vykYiaVmHaIiz74QjaXN0yTd/Ki0H2VC2TCnarBlJ54
6kPH7i/kqmTbWf6VNoDq+N5o4wvOYu2PV+tgOYd0fZFxNOZaB1CGfahrNp+UIA+mtBdKYPGa8dM2
/IxZPd+ag5F9T0II64Y0DrsH5peOTJl09tmkpLuR26OICRoS1uMo45ETybxY3VNUIf1gs7F1hooc
/+GFEAxEwUaljMCh7TvZdH3MxyVlVnDv2+t1Nemx/6eEOq3yt6LxisQ3x5mZHp0c9/gXnx1dbMoQ
tcdk6ob8sMD2vcknzGOu5SC7oFBuN6aAKZKbxIRTXohvKEk+jYB21NXt0qgGQTIIu/Pzz5H6AzH8
otjWdErTJ1ZRuasQm6VcG1P/FapyfIlT/u8NoY7Y61wTYZucQoGfC/xTEP8TL5vOBY8V0MlMLgTv
B+w8ObI7cUcX1jw7VWClfjxMYtCiCeTW+eQM6+FxBsZgzG07v6SX4DcHNPyj8GLNPtIQlt1j2sYY
OXjVVvYdqtduOztL41BdDedl9VCs01Futm5I3MMyRwoUv7QCiKTJhCV1oIfIRB8gOu88/X+af7mR
rLmi0z6X3mc/r3YhmcFMJzD0aiAMB6dufE0/UbrxoBAqO9ts2GTQYIbqTtaS5wMIlGmrZLSIBR9M
qPqj3N0bFHciYUTuj3YzuiWBA7o5ddr0/Pkaryiy/moGFk+tiAPmdMzs9t3izdymnxW6AZzAdj5y
g/CHL58qkaf+/Zb2+TO8ll42jjSKP1+QqmZ8+5OB0/0tEcuLT4U/5zQxiQlRYpctn5R5ISvitsWM
1pk9anDpCTzcmP2vijzEL86YG51I0B0AYYbD6c+aWMP+zBCYnk7r3GWA+hrWYicuIy62Y9IFyP1F
OEA6Nsb0vIgZ2/gxXL0PZR/GOh4LZdtO3xWTEhNJRwAV1KosPwi2HZDfqU0i+kaER4dAg2d8hIa+
uv7DtWG2m/ocOWJyh8qbGBjQP86goRDbmvM5EgP0Xw8yUOO6dsbwBe/f/dC/ogFSGfgUp8DNA4Ul
Yowz+fomtRTqIurC+5MZ3llSyfqdjbnXUdueQKcMHCNHmKw+GgsEBeC+plWmxdjZNKvhAkQN0O6q
TVzpvc5+cCZAYwt8K2pLLxGUz1WZBIYSzM6DamslEnWwzQexmy4BHV9Npr2CYa6MZX9lIl8joGFA
iJd4vCdetxiMyFxPld8HevOe+q8ZR5hp7MblTi5M0bHvW9b+IpvMJS7zZmRe/1VpJjGX0zdd9gon
y1lT38JF/Oj5mqs9K5vbCX95bUeVZpzkeZ/PFApWiJEzeMlGSlwdJ2tLZj5Eq47vBKT+3/j6AiQP
OPP4JIAlz6OekCt6W7PVC36zPC43YMDgb7Lk8TBOyCBE8+5LZiS/GQhqJCfyFIoQa//xLC8g2qVi
9GuRl90jD5UueeU0cjAPNCYdcA8l/+oqXKi/xyyx0Dys9e/TRVRcGWu8sugldYjfWtqLg6Z6Xok4
O82j5syeUpbZ8jmayk3SX2Ur8ZDUN4m87yt5xXa02iUSYOZjI3djzj31Gtv3Tp7md4wME2O3aSaj
sUv+5vG/tf0rH5dXRkPeJSg0LfmZnhK7b+uiTFtk3fMQrmpMfuBabLtCDxtoKmTmB9cdq9ZRN0a3
W+rOPM6BCXVYytV0Tf8efrN4HXqE4wAIaKexqPpRcaFyAvRs44JTgjZ9Y9hxrNIEtKYZPGJbjwuF
iWnsdhu6M3mtL+ndTOY0IuUHo7yH1whPaHm6wJ9191DzRsw1fJfUBf+rHzKuFt2xhGQMWao3qfEm
gYIkNSOPLdx5/4ngSu9LQs8Ls7mydb6WmUWTSG1JhxwKn1ndeUhewTJYqVR3lAqgqGr+yFixFqd6
z4DtsHMExsc2apc/20uap6TiHmr7VrWP/p8Hfdt6q2whqcvSCTiHyYX5IOY1brzGWCNoDxMbJS59
+C7P7GsIlsIZSwhNjBuH3Ics2/VVyf1E2EziGdTUMpEWL7eXwFjeW/c0rabjCmW801wZbgga0vd7
UYOmQ6n090rol61ZPeGTNo1Kv3HXkuKkjwpkQw9RrwLvgzQv0DhvYik02MhRrucLGm6w+ynLD0EF
2+06QAftmS54kOdZw6KECm/zkwNDoX89M08BWcPPnjDSmJD6eKsS4iPgzT2SUCzWRnxTrPkeawmh
Cuz/UGxIRBVXdFmGv79R5EEBWdLLHsSjoOz2Z7cND7mHrIwmdL6Di9MRz2mZWT2ihVxhiVAh4L/c
UEMsDxBNYirY8yCJXshtooz77QxIZbSuSnD2d24UwNYDiafM5BT1cASseV5Iq6f5zlHR5Wtmr3tb
/fRVABkCa9e03A6Y98Gp9SqVpyj/0wdIipFBiwBGnhpYi6yxNPOdp5I3v1lIATQpLRUMMzYbuYuF
jO2k1KlL6k+xSrHN74jOwkrsDCVawbi9bx+XfHgC6NE+QFib4ysPNZYuNGgN1SUVshDZi4RgwlGe
Jib3Kx/0GlC5qlDg0TnfCfa5SCnNFHU1So3giRBdJD9Qpy1fc/MbOcAw/fPbIV4kQmgjD9KbZ7Un
FApVQD8LJUNQv5W4xehAg159Fy22GRZKPlU2vBp2xFxVc6sHGafXRSwiFcufkmdWeZfBN31VPSUr
cJWbHvB1TCZAj+U524LS4p4V2QxaUfx8mZTO0EgUyCBVM3+98iw0deTSg8dNyf/c2ipYm98Jzd+j
Dqoqp5rFetGq5q5G/smzP7x0rxblp1O/1r1cGGD2E75+QlLIgYhu//z0BWK52kIWU9tLjceRfVFc
1TlSVcLFd3uEKzbgkUQ8X26Wz8ueJ1F9j2U4YT7BC01fl0bl3t5XuuUAXRaLMStApr1hvPVlrtnR
MU0goxifzkSVwUhJHNJYvQkgfadMfHnOhyijFzV5KvpAumcEnnFiGUVjPC+dz8uIRczVOAkhU4TE
7PwM3/420HxurdUik0OqgN8qXFJnZPINZd91BhYmZQQSgZ6mHopwCRF6B+Q6U/eoKDQcsqBJkO19
BaRrid/cNvEVCkuwycq5KIBgqrIuBVxEsGcpXGICEbbrQesKIF+PXN931FOn32YfGh1zJW1qLhzQ
ArQDpasJw1OEKOX9looomNnRtbYQiW5fTetym/NHn0H949jugaX2GTEUYllyueFBEYudOB5BxNmS
Q6BUhYFr2yqE0Cp4IWmG+5u7p47j+BgW2KKnZWlkABHivxLyye/AYzKCI9iV2kmm0Y8fqgb65/5m
hHAPvl1xJOqKQTYXks5JmRhmYOYG51lTAUA/Y03jPHSDAv8Ic9CnIX26j5JoTv/C9jIBkl7do9Ox
OPm24dRP18DoHOdxlMNsMFRxTGYzZ0/uuvHt0UdrxuIYDgEqXYyttFdxm4tzuUGn5r23fBmwpbdO
kFOdKotQYpZ8XIutk/89aK/bFits/M2WkVoB+fsGGDcHlbHsFvz3FB7VDjpJUIKiT9sXm91FbaDz
le3x8D+Pa9J+T46DM5DnjyULOt4u64Mv0uhWy48979BvjXistXUS+UJkGwfa/eQu4w1U0arEwnPL
S3igCYbDqt1B64DiWQ3bD1+8QiDIohqzPRSbiYOXAcbSmQT1hcHN4bfmbdlI95g4PCXFpVZu2K5A
tpsudmniMpn++aS0Cci4fRxpkm/ZpIyMM0WejnVFQeuH/J2IcsARpENVWCy+ffXy1JyAdOLTPkli
7LoE5ykjpxbazulG3jH4lYO8W9+JBE3YoszukJPk28e7Ltih//S2RxEvNce1mZWrmmcNsvzSlHI/
zXncFDcfvUo//GA3zBbg3kmkBc7a03tjBxDlcp25nyGaOl7sMoyqSSLyFQL7673dqRLF1Lj7d8Tm
aqhyFjZcwBRWXw9Vg4szlioHcIRTP1p22i1c21GrYoGzs2+A5NsSx7ZD2agFjyFirnTZX2xRx2Jh
Jm329XUTELGHSdUQjsV2wySLt+BbB2NNfspH3Wchfhq4irN2g5NuB9jRfPAtLyLPw2d1pODekY3a
++PHDYfk15FRgATjUPl3NS71UAjy6zblRy9vH5qf3JaVryEdMWVlOsBMuBFEld0wbQ4zA0IgJlwD
zbNbCii5PkVAJ9m1A5MMn0vkC3eLGxR0MB26u9WTBGdYNHzXXWsinsXti/svJXkQVY5z3daTgSZh
rlgLKIdFbOJV1Bt4PlkybfZoKD8Xx++vnVVKp7u2Jp1NRp2eq0r3A7h7z/l6sXgNnAPPUW9F9pRx
MkNtl+6aiuS8TNHh6dKrslWm1oV2y8WTfcYzVImy6mHOVRYEpa7skCZ5ajpSWh3ZFve+FNH14RPt
OkP6hnyUnnCXhEdKpTxzwodFbsFHdvOb2EL7sYK6vEI7GZ8iw8oyVi5bnmav7mB2bJ+QOAbU0LI8
t7zUwofNhndDqt69K8IqfywGWC+Zd75o5LsX44pWGegZSibjwZktZRCfQzAFcrvOX61kZW9WnKI2
tM0ZcfI4KWuSU4mtTP7CwvjunpWgf6B2Nmr7Xswe2vyieQyAuC+rnK+NHlhzynVv7khYIlhcU8X4
4sIMNpgbFdCzlPRcenLCyRPCxSwLpjkf8jyjYU9Cz6E6wTExed0o8b9miwNtuMGtI35URKfXfFVt
/J170kXRj/0PyTVkR2NAmcDJNuQPk74cPL3N10NjI9Oc2PfG8w2x+hdX+rWWUVyy9vWs5nyyUY42
wOxPDPboG+piX91w5kqIMPXIA8H3qYPgDhibesYZ4f6rz7WcPMAuW/MRtP6hMKXUgJ3ClF+O98Dj
Efo/MsIQtQvIKKqlDAy5mNK/rqMl/niobaIwEr6dUXaGhtQ8P5PM3INtGjKIhtn21b4ZdLKw8Gf5
UdOUyHqt8IeFS96iEpp+SZRnOWlGOVnlNthjGecgjo6HWS6idEbwDAeNDNkdswlcdvXg987XXWnO
Q8H4GylAUr+vXyP1mCGMR2vOAo7kBAjcCQsdYmKOo3Tyeg+hEngt/16kvhuKhvpziESihvVEWZGu
ptNh3+wtFVD84Pwjb7LfFxy556ZBaN9yvALUXT+8il1O0RNDEKVfjncb/zC5Uk7REYJBB5ChYDd0
lmQbYRMqScxlYQJhXN+PuiM6qSIuR3Bye2iEDAYf+izezs37/5D0hJZuOhKBdSrob64dAUQF0Krr
uzesO8OH4K6xZIhldvhXKe3Q9hlkwaCUTQEnZrqf3miRHnQreluvkqVtTn60flNkFm6n5KaH6Ku6
2oinQI9PhBkM8zBpGKf7di7GDO14VDZR7ROUaeSebzkJIqWBfVt4SpRFHimq892i5hbADo8Cej3m
C2CMYnyxZ2Ngd2bMkAPiekJBLFM1q3hm0fxU/rVSjyARHA3BKO/ZntxisT8760O7VmqZZ8kSOSxF
aNT27tbW4HAZcV4F5/vdrDwTW1VLTb20r/D2vGRMDHXI6M383GLZ8EYhOBMB3+F55MMvGB9Ly/Lj
+3OJfx0L3G6R2FBmRmAoOqyrPdwjjkfpe72T36nniFr8nn0xKvNV6at9Ne7R3rzSDAMJV22aH52d
U2fGgBFIOkDrOQ5Wk9V7bL08uen6qbA6cMVLW2rNoqd/B8witrpzWdqgqob5PEQtOO8D0v2+XZfz
f34Wjkxd2PF/FZ8AC0J6SyPT/1OZuSEK2fOlGKZEarBhKdnKYLRhlreL0mI0lhG7lpNrj3KjB2Hl
WaUs3OGWRJyWjJDAUeh6scWE0LL6o0pj5BVVOqMU12HxpwgMM4swPvQxTUoFxq4/WZfQrrGyHyyc
I8DgE70hFBshmMbj18q0A3OwiYGXR8gK8zE7JxU66kmz36ZtHE15e0HyYcDJDXrcb1HOVJTo0km2
dIc4wjRURafxc0Q1MZN1EkWs8hivBgKcze9Cz0QXgyy8qCcKVHTq/cYNvEHM0hdCSKyx1gwHh4ef
VdINF/pM67jUQpyIBvRSSBT3rbEugR4ad/6h3Agm48b7rrBhg+g0ex73NOpby00mfKc8lKopM5xn
rVcTZ/JgO0gag30vQq7Txlvy18sQ8cD/6jZsQgqLOvyp07xRqDJ+KIxpRoPAaJOeGmXT7Q95/8LM
Y169my46P0ndvrT/YQiANamE4yOrTGdAe0uQUdM9P3XYh7AjrkvHU2AvHv+zZiQk4ZJBmUxikd5W
scslb2SHRQLIfk642pUMNB8bXN9hkuz1xFL+haBKGGCulg+M7xxPvq0Vm85NuCW3G6CpM8z+IGHk
awZAV2fKK8BDrsRUgYPxj7OlP7s20B84YPB229N2Te5BPqB21j2I0o7gkw7XCnx4uLZ5hRaYpBkw
9D9bnEylwDqEZxD8PCd9LscPbwErKCi2FiyjTy2fiI3CXjXFnlivE97a/m2rCnn7M2UWocS89KZE
AbhZBhEcUa17W6/YgBu+aR/D8L5PP9q7xoENHiCdH9XR38JsDpUp1a44eaezPK74QS1xVYW4Q+X8
PKEP0Y0HAVPBmBHbsKs1lqUSAsPavwfIRdEAgdsVmidxzePoWvta93iVcIzYmdLjEjTqoGIvMQHJ
uA490TP19yk31uMarzPDOpsVMr8/lmV7XQoLiy2b2ORhIRQUmf1r9zfxcAeyUheSv1M9AXqK6Fj0
lazD2NchQKI3guDIToYzzZXJB91yssbAZbC5mX6oxAwLZKkjyulLHL8dIkCGnRmqHFPlnBmWtKLC
cAXNX5Crc0sdGbqsGqzRytZPZjRbu8wOvPxTvaFjK0XkH7TdJ9tw7F+R3gCMl3BgMYwo1GTajcXh
LBygppi046fShtPoZZrrdF9fAR3W5u9HyuzVw1iRCskkuuJfrdEvj55saLJkoJZ58xssBRrZ0uxo
YcGhVec7XUmSfnuhbjVyffCug1fpiCd0YcO7Su/s0/THTVk+Rovp0zCzMI7FktMGqes489KQZajC
/4Ue2XYGWHPfBUeXKApAX2MjqZ8Wu6TcNP9JFuSgHzaOAiGPBPyNXO85RIACDvldCLN7ScWQOSxs
nD1sZAKs5z10PWDI1uqMtK9vs+Pcdgzzj1WI+amZlulbYgsuBqk2ac5oQqDdMcvkyN1JsXpsHXth
0uTLuKifZuLIkYgtd+dKhAniBZVvN+icF0Ej6IWIIQdffEGDlmM9Y68tO5l+sTy4pLwmE2h8r/aZ
rygRVCHG4TuP+51ItiTeAkU3xbMOTr7F3P2ZhN1DfKW6r+7PXfR7i4rUm+mgLT7RrhsJffLIWtpw
Je+wnlADXWVdG4QrxXrLYJWkrD59Che8/giZB3zZuqvZSNUN0I6moM79GsQZ3hpYhATHiUJ7xDmr
c8E1SnZUdqaXjqABAO0DLf2Hx+JSkz+eO6K+Az8VfL9XPu0qWwI1hAI4knDgmucG8L1A5pCu+Z3l
0eZ7Zk6snXYSn6W2JkHJwOLTimmUNglDPedyBcaNBLUwd3Rxsv9swdmeteVOM2z6n3UVE5iM+7dR
ut3wXHdo5S9O91hHkYELzI5mqgaE8Kcsl80aCjkeaDJTQtR3V+0xTTyh/tFH43FKPixDLPJju/lJ
o3vYvOWVbPIboyQvu9NnKsRzYj54ZyGQcjjvT1TnZalzCYI8pOpzjsQ9OofBAqDs2En9Vu7/ZpJg
ZVdK6MFQG/FA9ON/q3PzfGNbmw6gYNxuGssKohw8/7FVFjSOWT+aBAto7XFQTDur5XKlMuFmrOd1
YM/s3iFVDjc2iY4BgDeHTUSnVd+3/qgmVHIhY5UL+pIWM995k9oX/Xgtd8/zQCNh452rSMtlMT9b
uOySQYkBcBDt1V8SmFDiQpizqfVVcU25HafAOK0zMQNLCkzS/zQEHG3cMsaePe6ovsBepFmudKCn
25lYCiUyP7H2ajKevuU3NPPhS0ekqkDAgbMtsep82OGLskzgpsvtDUHr6Kfi6xagt89/q/bkXTmo
EgOeakYiozCB4QRmkdAWkL5ZbYOZL8MGpbucrfRfUlMbCPv/Lt/3CqbBlaX2dnVYVx8cQNALl634
bWaZ2ZHx4Cinocj9tETnxyypswfXvBUs3yfiJidxYq/SJai7351WoZIe5GugvDpBwxuNTWfrd6b2
KEbTBGfJiMAgH67zKmiEbxKFHsHFJ7LhT33X8Y8J7/ode0xU6HcyrpdyGg1QziL/8irew0V4Gbnf
/tqp20HN5tmbrGk8Xa3pTa9ZPkKGp4KnekJssgeNphXZPmaQnm2WrtAK8xNsh9fBDLfBBk8stJnD
H+uLXSuJX0fSQGDZouZuu6nBS+w9IEZJJv9vL0tcU2laOulFTLr9SEvq9zwileHEuX61f+3IKpFG
svqgk+rPEANbo4pOQJTSfGYMtJvJTnFmqzXEn50NqFkuhrks665ce1HoSNeItJsJrpmS6lnlKBYj
GG3diOjc/ZpNMBJ+XFYpvACmSXmapgj80pXd3VXA9tidsuvFpnHT0Zb7woxwz+QiJ7x5Wx8i+Imf
GJ/NiDCth6CzXH9whhHhqgyLN4tn3gGOH/0re3z6IyQvJJjMV/WWf+aLzU0t5ctNeIfd9O/1rLZR
xA5nlsoIdtUwDlL0l/TWMGwIkbPDoSURyLQc6Qi6bVOXm6Ixo9eA273FswDtC6qZPxyxuYysjwE+
Xsv3i8mk7bg0WvJMozaORSy63IWk8dR0HYJREm5LnDWK/7YGMhrAmVKzZ6sULluFcNdBPJnlD8Q6
69p2veDyYP+ci98HYkTm81rAvg70q0Rx9Vis9rB/ZBrRrpVlFKpFiQk3iOb8Sr5euJmFsasuSMit
K3FP8ZQTihVvu8t06StBtM1/pUyIsYcxss4AGRSCo8qld6sm41A1HZzF/Vm1dxnGdQosN2Pn1ufz
90fwtn4osHbRI7aKj1YAHKmAtkFapk9zcDQSBALTwtSOhWyAwuMF5KF0MmSxzX8XkoVy8gI5f3W2
duCZBIqagyQrPxzrGp0LywE5HUsJn4T/8ZZcWuGCbxMPD+Chg/JTzM9ykU8kh7FY21xpE14dvysx
1jJ3wrjkfvdP7O3iB8Xg3oXWIQF7MtI0J1GLNmCIcSM8oOEIvvhOGVCrzDGGapXOGFfieGLAblf8
tJkn3omnjzqdTwzV869nhyn5K1xVX0K6qJwOVogn0HiXLfGUFSitchU5QE269HfbWoRW3KH8wIes
7tQ+cnXTtAvSy7vkWEB65IvdXf43gv7paxpIt5jFSQq6lwqCOX08ToOVowcC9EwscXKRoiXpqtak
C94imHgpy49uzgeyDVnQ85Z528CNogXtnVDq2+TR4+TCfEfIeq8mci6yxBAX4wk4UwiJXbxpiQyH
5AjwZey7VBLQ1NaEE3qKFUPJv5OTpyu8bD2iAzlyulfjK7tI3CONDc9Eynu7EY/tZAz8WeyvdvIq
GtNbQeLMjmntOkd46JvuY5xT30wilr0RteMH+d57GNJ0d1W4j9bmhjOwhWNCPlZC8Cm5+5hw6njh
2vt/zCU6AY77ZfQBxYC5TXtz20xHJwF3dvpwctStNjNtxNml4Y+fDSmuc+6/upllJ65G58ozq+DM
dZ38lAoqxzBm7cYc2zuF8apF6tx24LVaaiGwaCUEjMDzufuEzvSmE1o4VBQqSzxnrZ+O3iLBf0vb
mVINgF067QNpAiWJZrZrEs5smigzqFNFlSG2UBxYEuzrrp6RhZKWOgkvxGzvBtXrnRmkuILY4nHQ
4Ok0BrQQDy7l81mOURfbscpLrurPPXVn0HB7GiFKWLHzM29r4R8X68HR2RiUzoJw7aROUk/wqKFt
BVt0URbHqdcrE9Xn1pf+TIPEQnX/u4aVdY0R96C5pQSJ8APj6TMzTZXQb+yn5pJDkbjtMzV/s/jY
VbuoVEvpg0W5PV1vzLiCbVvJE+GRJGXgkOAQOYRbze6dB+fKFbPc3KWso4OqhVA4zyvgNY6C98pN
dSyR459UMKV0q6f1RImjZdMH0vLWw/B1BavOmw/qhOslHPKDU/BLgd8UlzUxKLzmxB1dmNvr0Et7
ySRK0gcJJBgnvG1rnvKjF0uEyUzuC3TrNHTAnTbwVeY9iI5+AjjFP5QDOjUepJTUyhTO5FyMPSSO
fVZgQRmA0l0AVNcep1v61UotoqUFucNvd8NzVTumKwZt13s0wVqR4S3oxjxjyy7QgBbcg6FL9w8q
QCA+RoAIq3i2jLITjGs3iFQHZutPT1WKduH5VSjP7019BpELmtTZBc5BZDUevzOf0w/C8Ls4248x
D0EHrVdO2rF7XiVCpYaLWhcarUrHW4x8d8aKImq5bh93UR+Cs2guAmqVqDHS03mM2vxRFbJvy8nJ
NHEqP1eSOTsBJb094MJq7+wqLACJzao8g+DLpQGX3t2ewT68aTQAHBuEV+g93am0Lg9dbuoS8MBX
IoRZdjDApdXEcxWWtQ55RxXoD5jkNBCIb5XT3t26Pf+ZwwLexwHysgSFHTM+1RvFuimLehihktPI
+v5aT+TggL8wyvUWT+BMmkkl15K6hAslWvG6TPvPO0r9elAC1gzs+4vsoTscDMqEtwUmnHx1u9Vd
78KvhH1P/73uOkaVv+p3SyTiK6eCyxiyyFdgqulJElZiTDc0pbYZzDFBMLpmeCWyR3Z9DQvn8njp
fyxJCIkVzuG5HKsbSI3c53hEXt8280QAdLvlG4+4Wnft3CWMOSpB9JrfiPMFEi4uCL/ebqX4IjBu
F8R0h2fFQ+G0Zw14b4os+WR/Km6F/XQ+TemLz522u6E/SZJnY6QNLH/XJMfw1U/LfaGdrf2P93DG
zpQf8cZMHjOBzQkp+fctEUP092NcZZe7o/7qKYyfJGzBoSW4jEUw28V2m+9SR0YcQH0IQjtN3JDT
hpw/6kL+n2rsQyCTOCojdomkGfuhxMdmeG8F4gb9kxBhgXPAOq4dOjK4/lbzhIDPoOxbEokmIfZp
SUg4hkJsAUgFihQ4RUmAPgQYUDumQ3GqiUnliP1F8NB2x81Ghh1KpGpTfcTR5cCcXgL+qv2Kk/cK
kfpDFIDun9O++wWL1rauAxpbgiFqlwbLdFs+ys9Kuyt4yBLgaWm6celD59W+4z6ViLd5RCRVY7YQ
iczDXjEhJfV0lEt6KfTpvY4i6uBZj2ff/vJ1HQofDcB7slPZMvdCr1gs48gaOaetpRx4jzTPn1Er
2mq1ebtbv3Kh568WJuY6LRXUo/5Iz3Fpt+1Clbje64VpyNEkxc21JV8GhKCIyKtjGa+EIcPE/EHZ
qEpTiCTtpCzGDWcZ6BzJknPE5LUsQAb7Qlwq7feU4u1mbtBl2s0nQ0saM4IxAMgVDehDV0GFi0o8
5nH+XxX9Ud8Gto7bCyok1cozq0IpyiyD9DqZARWu4VmqX8k10CramwN0MIRX2D2+9PGXySmxFz2e
iCDCdJrLgcZmEX7IuPthztgls6g7YTd57z0nIEm7SEH5EbIBUUBka0SIBxR9+Lqj1YXsYnCBqNrt
RSY0XyUAMgdDK2q3nlf/eCtVDABqa6hG31nV6BYx20tOzx6g1FKo7CHFj7Ag4Mgdaep/kdDInpxV
NT/QBIfRkxPKqi8twWBs5I9hqrMWS5A5dsTFnCJnqUETmPXFmqU3Trj7y4ok6sDXc7ZPpSZH7qSh
hte4jk1aKX6uGeMrUxvzmsseSPIlxVZIfVRferscrTuVLSAuCUiiDBiQ0pUXFVOZ2s+BIcdU2DMI
/7kUf+Fg1kCzjg1AdNZ+yitTTml+KsYWynAyHLJo4Wc0Lb6fazTEKszpcUcu+TNwzrb/RcTUAfYj
Fn25JygP6PKv7y/Us2nhRRG+9hByUVCnwWSHuR1UFvNwbHvVy3mxZi3IE54RCSXE4G+VpZGk1X8p
JWIGhn0QDkW2bVDrpCCQ2ceoSavohPu1GQQnow3GdCIHmfU91BeWHtf5KnZXUYSpeRyp+dQ3e7Lz
aWzbbHtFlGGqIH70CQvzFzUMrEJHmVBImeHOSzwbNp0Aeyr8aKTiaY6pjuiEH0A+T6P3XvrvGs1j
yzkRdzqzrF05//aQOFOjwrjIe1vebDGjbz4V79zSEvcxnzcKBi2A3iqdG5UlVlGureSwnPiXbJH3
0YNmtCB7OwDIEX4nzcZdUeQUxMvYPc2itbx7vlzSoXpsRpj+8xxK6MKvEzrOnIGySB5NV54BnHBb
2/2CVvXsljdAfd4ddQqb5ViJid3iHLPQFVOTd+ggjz10uCvPLiKmSy6jrf8QLt1NxJYD4okgWWqF
KlyLoauYgkLN03hiTXnR92OVbWJJa0d9yImDnujPr/ureeqPHib0v3y9yMDsUq2IOxG7sR/Chzme
WubggsD+1vD245OfUUsH/ekwfiv5yjUus77Aph2hQq7SVE9xNt+YN+aMBt3J/1C4LKvCu9EkqvyP
Z8OZXo8C5QSM+RNKh1Wnn314oRIkzFTfH0YOs/F88jK9BpYKYn0leX7BmaU1+Iqro3l/DsJuprEE
HMYw3UpsnJEuOC8GM/YCEfV1z5kn2VbwuwLx3221TfSy+FZ4GE+TA8nviQbq7KxgLXSdbedrRnhb
Wh715ubRQG5znN6zK3UBcf5VUFnorUjaSLyMf4URqhMcWQnasUcxR+HaygF8xG8vKDb8uXTScjrE
8NipSyFagxEI3IA8/dC6868a5mUNMeEq3QhH/nPn2JJ6VTm/lap2miqtOrmsk4TcMkx3UyQ36G6Q
X61vZf4PBD7CJqlAfxfAoNonOSWi04uo+2odxDQfBxxTpNCt38ICk5HFNhNY76lf948fhlff+FhL
QRa/L9/bvkU4VRg/ZOJjJ1Te7iJiIQ1eSQiWEz9prHzusWG6IcltnLG8TnX1aQ5+6DCrRyi0PV7P
g0jrZ/tBVsE+KkmV+PaKhFTFuNz4CvIJov0ZXrg8KfsQu6FZ10UlCoAjjE3yksvtoYZeqjdFu6Iv
OtfXEUOgVjV1/0EDBWnKpZEW+RS/UyS67iDq+9CSyj1jluQC1fIPYQHQXw+r22L4hdtjZv6sjMw7
KiozIel8muFK1Y7iHMYQSvQPw+ICqutaNlVFU59IJGH1WDh6WmhpRz0nfPg+TIycVICkwBJi7Gsa
D1Z8uNjtb4PQqHEqAOFpVczE+oxDD1K0gkLjqn5PNHQudKu0YFAP2whTxaAyJKYlvkcGBBfXjhd2
lemFj5UIVc1NVr8A/j1TPoVcLi1++I/SoWoLnSpkW5OFoknW0/Z4myo3yvvIh+w8IFHvDhFicmI1
HmUigkN0EEhNaFVt1GKDm/wSYDWwxQi/2VWcMxkoOPn7ugvZ6Uqus4fQ7Z0NUeJUQ5q3OHoOFTm1
qBkarMXTxxLCFO3x+eEcmLbkESuj572jjxHsjI3hO2lqvI+enpuAnYcCAvyKCen0scE4W5S2Ndlu
QbN+Z2ypsrX3AQG5VKlRE+mYze1P3SkK/uvc1QcKIcu9l9cL+wEhmGP2N6xO3c+aXfFEtPCcO43k
hNqu/+06dzuvAtwjuCTK0EiQTYRZetZdyig3AALYxoWoybHmHti4nIG4mb3qpNGEwDIy815f9C7C
COKuF6gnBdacoLP4AQ0wf6/7cDFO2oQUKMwigDQZSNxHOwOC+wPNYZyyFtxmuSLEszh8mQygVBFS
7TnzBQ97FZPmqUYepQSXFfnyqbAI2jmuqmfmTobGndGesE2/css2F9IV4aMR3pvBtcIX/s18PfaY
qW7VDBtPEDMuSdPRX6nPK3ZUWMRaM8BbAsPj+hvrejmTHXNwswHijT9rF5hgiq9aqyjCASgCuUrG
bHAQbdXJ6OkxHzQOOCuKyQXYe/oizBDJZ69lrA82A+XFDhzMvjr6lSA7MldPTcR1UNl1KoRVi5t0
l1ezLEQiNn/6Puk9pRHGRJNH6YddwWC3FmISyZMqWuyxWsDVod92+HBtocqYsk69mNkhbURpWjcC
BPWjm8u6Tiyq3pNv63t1kFXx4D9k2HSYAK5GakYZ+CQ+aOGlPaQMxxH+8st/UWpjiIA6R325liTS
jo6PK20xh+bu3rKE1rvaE/HNKFAd/7ARUX1v8AWHnIlzXBDFyjBCvasQr/enLZ8vZL3s6SbsKFPK
pTXrjIq9yeyvfNmKi8qP+fmV//1vxriJ8yPC5d2ObvuJPkfDt08/jUIrVgGt54/0ams3XzQo1ZV2
k6VdSR8b+fRGRN5GjoID5p96L429Cw/+jEuh9SrwxUINcr9KfjMp+/RvvP8B45sEQpXLqkaHpztC
VGhPUys9yvzpOEsfoMkUvvjzZ0O9sJOhWqic9JrpnUKCmtqxJd59uWLWuJN6QRKirKVtN29knR0S
fJktAhbBlk5FXNe40epunrC7h5B6k1xmw9PaCCYnhlOHAVeQbAKeMkvUyhUjC2G7QM1Zht3unM7I
tq4ZfdJJ9mP1GrODMeLfeHObMDLTGao2Rqk8YOpwvLu2fZZAZE704tkh2IURcCwRysPAmKxylR5n
jx0QW9OdX8mL8M+gI6sJ4rK2x7H36SSz5ZpkHeGKxcaeLA+aog7PIWCJPu+qSQOdAde+it5ZBLFJ
EqYNHWQfxChfePNuatMbgYCSk4k3bKM929IlVH3b9CyuJuXsHwuLSV/2hrZyG+vsSv7ch1UKybtT
vWmnZKLZYWbGeDmiao8xOlqfNVNBWnPvVLiU2Q1bDtxcNDD1apBt1quIEek2t+VIP5uPx1FrHqP7
S/nEu2Cx7unl2kmW2yqxlW+/JcshIN6tCitHI6kug7kWPCRxwgJ4ooXGIbAs88q8kCKTuLXro3qA
wfVFP32plwCh4dZiaVj+9itHgebxAnmUw4Ol8btB2EjtadWeB3PawjcmHfSYvZlpzqYUkOkS7mY2
VZITvHUokDx7Za7wvodTtcac9JNEUfeWO33iAlo5nWiBySMft0LPIY7HpRvLp14U6lhi5Inh+F+C
c23FX9M9Hg8Z8gzbtggvKxv338Vdjsbx7rSkEU6C05cEiTt4tso+CiUegB27g257peiVzxBmnLA+
a/+1r8ijWD2Xnl5mlZmjRvkvMjEK6FItI763GIHPWNEGOLYAL3s3afyt/PSbdwHqfH97ps1tddCp
zpSVvMxfhGnISLTpFGzHDPKYh7isGnJHl0XZttVGN1ALlggEBfVjBvEqPocj9mYcGqhUcZOBv+oq
pzeSw4PAO3Q4aGMxjdfBI6N26/la7fdMT0JkKCqYlzBRGNKiyKU0IqzqUlmf8rCvTypQVy+Hxm3E
YG+I1QAWpwvL8M1nN+dvO2k0KwtPC8npjJ+9ta0fYabb4j/kgLkVnInHJrUGrLe66jWmLWqkWq0E
R09IUxgKb+DgQt8SUF1kBBNsAfDzl30LeTsQYjXuNDjvolXqTSiXZsy2GzQfRi+Jrwq0AkeKz6hZ
ydOYGxgLwzkT5Net5G1WHVS6XnkpHx9zzMlE58ujSFNUbAS90awVFllh1/vQq/uI7j5Ad13TpqrV
sED5lB+X4ZeXTRrFy8qs20nCIDVpeN1Sas5ulmocop/4lNAFZRDtDHkusPMPspIeob+Vqcw3oS+V
YEAmOp2MWwSTtLzg9tfo/N9S9ODGqRyK1NAgi2i/hwo6SqaLvgVEg5AYCSAt76r235hLiDdKxc7r
DXydHS/QD5+hqK7fAQ49pM7PE1a7LEGnVJSgSj5EXxq0tGHvQ04GBv9b/V1HZqsL68GQO7xMpFKB
+sJSwVf8XEeedkfAkotRVftfZwEJIbdataH+SOYZgXR9XnPtdRT0EYYKvN6AhmVnUdtVLalt21rA
zFh0FsssVrE+CJg2enyIDEoxMfKS3ovtxSmk/IhNECkRRg3VRFpINKgP0CygvX2DwEqWLUPlm5yn
8qiRxjErF04fxWrp17u2v8vM0EO7RClFe0dRL45Yv17MEMyhe4XvEScPedLBihO6ZyTMiKpRO/ki
6vYcYdSWoiPQWTTqjsSqCzel/wAxEYcb0F6/gwuhMmp8ueIxqyG/pR5G3bM8gi91yBE3pfCCj/VE
e8ajM7aKCoGrXtF4Tbw26XNUkqOvkpK8nGvEjexafhqdlqvll0C5kQso1XNc60NB4poc8AobSw26
cBzZYHPuhZyKdvKmbDU4MRaSzNp+BYAchBRXDlWm1Is7TrIB2hmmfDnunDdC/r+M/lDwlYLnB65P
ib9TLDBMQzcjPebJoB/mh0Qk13aldqgJgtC8H68z2M/BglvjUL7a8fFS3SqqVg62SR35aZ+LCWtf
oJrG6aOb+vETDYDq9lG29IsnXlXgaJKumTt0rl6MCu4SoMF27+dfACIcB4xywR0l2vQL1eICfXvt
H12lPUkT6LxdP+Fk8pmwf6CsnuTyUT+3iOPa7As2x1BF5V473zWMDMYSYJc9VnZk8PBs3XI0bKP3
NIt4r2Y9a+NS+Gd3YM/y9m5Ywk5up+Em+j/3PFbDTvqUFUPhz5D7aY8+Fr4GJlB9/PKfmss3JiBu
5nxnRnIkHOJmK68OvKw5bm0LBxtNijur74q8Qb5ZmHF26sA/x9DGZrB9v0wY7LVojhV1lAcsGnU/
i+h2nVn/5SJyWGNuLGdeVlbBMD53vyuIQPvQqacUy/77Zn/UwKPvh8+QYfdHMoI2X2TtrWSJuW83
hf/LIblCGjkPTKzUuIUhsHPfpxk/wpjGK0DwHbYiQ2+syNeRqpABMS88ZXFpoFGOxHLXMZ3ycOFo
ygCS2tnH+9cpF0JVIbo0atITMYCx0d1wKsbsIwQXyJdv8RMwBCRUWm+Hh1CNEUZzV+3hZ2rGYQ9r
U+OQi4O4P+WWfNPHu+yPKtbmJdupi7Scouz/egu/wCjGK5Ae1KdXGljpjC89jmMAgRXSRnGgp3fE
dDZNHWllLzV5nMvMvVibdtXsEQzST3PpSLPYojfXrT5HB55MtjbiNyrGMrlBaBpbiLHB6oGMKSxO
zBRp5Fw1XNPSybxS7R44VcghZOHY0JM2nDhQt9C4OsAJvHPYrXVSXfik5s7Is9Hy8lu5HP0G/F+/
znFLb2oQxlgYiVpZT7VhS6CqDEoWOIzaqM+HvRCUvxF7JDV3rEv1Y7GeIBh6wIzDCF5pV1lAeiHA
QvT9OCfmf0poNDfM5C5VZsA9yAW0hX6fLWBFqH5R6bJpZoh87CVfw+kThLXi5uBgf1Jdo7YjtFaO
AO6sV/ZTuo+Bx9K9M9ijMUi1JAfJOmReRCoTPlXYUlhDSgSonWIaam0Kj+Xb4LmTQnnlrVE7KVJ4
0kIzzo9u903THDK9qfA/wggTGkXWpwVJLrLucseRYohxoIPTbxvZXQE2x4Lnc/V5xq02AYQ0YhZI
Zeep7OoX0CbEcMGYUIz3/rffat5kG7YvxqSXUvtpCRDjT5rKgwfyTfvi0zHSFA0v3wkW/g5zXxsD
OmCqKs5dSncIyEPmse4jLtdfUGdJMoz5Ve0X5k6TuTNjoaQ5RzgsgCr3sv3vo4ilFSaSILQqbKP5
w4vjI+7SursAFyCkEZWCumPvPTu3xgbUvpfjvY8YSIYFDNmMuvf+lvf1gFaJKtYbLAXKwh2kudXN
UBmTz/BWx4DRYajTKCmHOrYCpS/e7CAzpx63dm2quSX3pn5xpiLBJV3wTgBsoNWuNoTxqAeSAYFg
eQ3e0wsjfAmCW8trva+y1TDLCyQR2jTXdrg+xpzZn5lq9vRkn2g9kuMJzjQu5ItXZMQrb9Ezr2P7
GmTom1QggixcMMQ+2HxkkBlkNNe+/CCVoANvDBeUxiHE/dMc9deXYFKkmP45pwS4P6s2XCH7X9wY
WhC58FLxJiCrjEkX/o+mcdJntLaw5uT1K4obgpGrABEDAngZX6Zx+Fhol+duQNBTkPcYszD2KCvl
qlrGzlQ6piHB3Ft4//R2rFjQcADjpOGjP1+qGp4tBO0z/vaX5O8//oXATfYuqCDBTBrQ2JftJB/t
THOKWwpnxubJoX4SravFvQrVEdDwj76tkXgEGu51hZZFD0kB20Vx0g0VbvBhBcqavVQVK2VTFvq2
zI2Ko/saf79q57lSdRzcjW4KitQaskfYlDoZOrGXlhf0jl0n5HaUz2K1tTDIlvAORxpaQi6gbULv
x8FLag790fhuqUytp8inZQTJd+A8RdkLRTLiEFUEjc96TkAW72Ub+MGq5N6kq+ViipirfrDdMY8B
tw63eStzzdSfMyIeWj/rrDZiZYLgyfZuUdn8pTOyTh7TYOwTPPP0DOjquugIflmdoumeHJXoLG4V
LsdMVrYFpImNRtkMxv4HPuKkkIezg4GxtWD4azGdALpwbGm4DxyNOfQhqnrUbER90Feh/sWHgUC9
oV71P5dfoDCdIxe6RXmU1JAXLJR32w0DlN2iXhsHvXZJGiY08a5qd1IRg5E4f5LuzNgKJajzvNz2
JtCkVJ66sWa6M8Bhz71ofGtIvg3qtSMQTJZElw/4T+6kB+8A3N607ek1/AqZvwnarlhqvmwIjBky
QOmwWNzNW+CNVmeyfCjuYS4hTwZgTU67p/NMCbYnwWh/sW6FssXVe7KhV1Yk9zPHMPIEoK7H+wv6
hz/oTcqM3ntwINk3Xe0iZCPLDkaH9MSlYhI5UQ5b6GdWIobE8UJMiWhbYl8eN5JUV+VEevDiJvgo
ZMf4DDnJshUfLFbaY7gtcYzS90pH2+G0EqHddJ8xS/j3N2jrwWwiOFwxPTCIGqcMdbTxNMLHY1WL
MsX3I3tyGOne3lY7I8Tu9vKmpJLArDhCqg/EZiK92dCWOC7bZD3iDAwEkbf2cuwhJHxSTUgW48Pw
lD6mPRGe3V3KvvJBXgRv9ta8li8l9afFMkK4vNAJ5yU40cf9I31uFcgZKYilOpd9Yfh99uk+gI3u
A0/g36rgocSmSyH1wWZ6n/FbvHKl8PJGXa4p5fN8bb024ck+A3dO10D0dsEQXgEus4rR2EOuBWnM
37b3Ck+wGAJIdUj1aqOv490slgX25wRNDdw89fnyFwdVc7lPrSwoaj9J09TrEmliN5ht5y2Fhu/L
iQR9DxA7EFdT8JDfsM55PRuC6J+xDAUQ8GFe5PSLPph511uAE0T1+JeR/Zb8CffcY7C9kPCKSzN6
+onVv1wjqgyd/v6FAU/gZkwvdHpYlfLbveM3b5HwMhLd8H32euq2VKA9vZmDT4K33ElG4SvV3x5f
bMbkWckEgHOWj0s12XMssD6joB2w2UdfdMg+wH7GSAxfSJeetmRXoJVOLJI+3T4d0+n4lIfmDB+x
HaUGlX4UwCTb8sEYUW6zWGD7S6fUhe8ucJy2ORJxNZnNBAWgDxJD/i98smmkkuKyP+GrSsnxQwCC
ZoNdHEybqxMxEVmsIcpjA02Njx2MF+7xMPNPUhqC4Tvtr8s6ktQ+pxipWIY3KkahP9azVYiKWkMN
JMoib09XHuwBHfbcbEIc+EIt18poFuYbnw6tRLllFPuVdztYJ5+77I2/8QBBzR5NwG48DF++XSTh
nZMg+8j/sJDtzqxfc/pXGP4K0JGsasQlj3uyH53qkgNm7jY86CGcbYoYClF/p3QCuBbwZGV7ckWB
K0w7Pd3o2XEFtoF7rQlmTQoqjMLDeEYosKGXv3ywULhWUkhQ0qAZ80o3KVF7J5oW5RsL1SJ+IUlT
25ClmOLiAgA70rK+1nEvD/jYcED82+ym92nETmSRfbaaeZNgt6tl/a4Fd2WOCCd4WRpXUnF0nmDa
oByTAsix+NFqqLlXFTWIwjOgrRImMSMSKnOGhwBv9sommNk49RZUG0MS+Hga0T/7doMF8kEJ3O8B
WgbCBc4fgG4IIPa4W6gRvCfv0S7/qeOafCOijSZejgN0pT+NJFyLD2/UHjnsS622XB4la1pryNXB
3I+nwAiRwdsmnloUoDusUQ9Dxloi+LQ1xKRYVoynartFBxshxLuYuDM2g2D77PEmlLQRkzuuyKsv
TNliY+2aD6ye1DuFulZkrIoiQd1HPUofqlBRcM/34tkkGOB7YYYSLkP5/nM2B3spk4zGftu8/Suw
o+ozrP/jLGWiEyYoRtdv3nh3lf/IvJiPLlr2fgdUrxGsRglPXkwK4T4h4ysacRYo3KLSMrcQ23HU
QQbMWcBYuSvQsYvOiCVgNjUAfwShF7ckfK0OMYZAw0yefxFKRWf7cGvMqh4kWf1z53BPObBEOQw9
cNg5Qd60Y1ukxs3ZuT0vMQdd5ONw1+XbeGRm6eyrlsXhv2Tj+UUruhOe/lGsvdEX0hwxdtmHG///
1qpHuJtROnOZdn1XoAkGdjk4K97wsriItW6junp75xzs+QHNiht2Ab5PB5Z5SNCs2DT5yNh1Xyw2
YEdUKlGxMR8GjW9SXSKs/XN/CUmZhp5yd/sPEG1xaA0G20bdeV2/sEqK9ud/cyKUJPiPmJxz2fZo
W+WmS13DN1eHwQn1mZiIgqwg+rlEF3NhisGh/FBCpUWVlUZSLzB7r+LFAKxKN/D8hawewz66D2VS
l2fyodgA8d3HsQ3VB+xWD3ldB+EreMtqFc7rvfIUmruLIJE/LOAmCU+4JoIU9cJpKnAjL81HMCzL
mgcEM3w1b+zxK2K8nOnOb5KGqJAXQqNc/k/AdisjLAmqAEKFQsD/GSZhod1WXzwdJpo8GPNWuQPW
8jxyaKiOydKDWPnxfYlk8VmXu4jxA82wcYfvzTZ9dqBUJ6903A+EiQOdFc/pcbijEsdZGdSSO+Pk
4COWztgD5hTTYgpYhgyddsj6zJbXhdIGNoR/RsON+tBvna8m5jtICLtfR50rJwoPAgh7fvMaIbMK
eq4w7RHF6bzNkR2ceSibv17kOkBjDbOxd6iEl1siSmGPpYGRvjjQC7Ntu0cvrHRpefDHKNpBsG3w
X9j/FZmP7i8kB3l8ZLhngX1llmdO/tc4TkzrfcpoR+yWtMCXv2XBHTCHkUcz6vo0KoY/XrJXQ98x
HxJawJinODCsDKZi+v2e1N0ggYY2klvqoc2YSXNuZ6iWaLdiO+5Tjn+1uva7OMW586GYHn6VsbEG
6Zpb64LQ62FgK/qiNsWZMhNfoZPlD1GJMaojpoggLP4qC3PCimvYOHeCebZOc75QPcFNIov8q2d1
YkK0Gak/Avd1vbTs0ueyzINKqq+RiFGNp0/Knl0siaop6i48wvpAjsC9afenMRklCRLeAFDT7UFh
i3LS/o7/IbmH1fhy7G9SIu9OJ7LYSN5svfBULEY6soXfFf/tYy6TiNXqNmwzRmMkLT0w64zXTIER
yTBZYDQKnlmUKxMkW3ynPAdHaOLANf9oaxQfw51Y0M6pb9vO5x8EDvcvpzvEw4hfJ9ua7UeeJOKT
UcIzzV+OZOJlq0DOfOUb8kNEMWjPIR8NhzPCxrkkwpGHaDhn5ois2xcZIG1eRg+30w3V9Nxpc3ZT
NAYezaYoAtWAjTOJZ/qDv2SLyINNsK39OUNj/dgUm3FIN3hUoIJncou8IEV9woRTtk9YHcaPJJLV
RZOpexNCcjnP/6qLGneSRd/oRXvDIiT88mkJEJNjwSKvs1WH/62P8LYpOA6DW5AhT2L0chhGKQ8c
nSyW+g9I/zKiSOo/v1pZyiwFsg+Mv9i363rE96jXiRyOBdo+1UdIXgSo3jJYZv4GbEdsYAlngSre
QKzd/S/ooZwxjO34o0B1yM9QGnw/skgCWVq4gF6umFKJ7XeFKv3OHUkbsYpzZor8N+RaMZDotpD7
Jn22RJ3P5KnwUfeBKxUKdRLCYwlzJAiMzejw/1DHdagUjBWofiYeWUY2seFmOyfKGioLQN4rOpbP
80b4leDTpuGavWK8RPN5z1JuLMmvbeLw/PIdq/uVeQ3JTT2znHh/tGO35Wv0UcHXcM05JhfEFgum
6fnRfQpH7qMtocVZth/QTEiKENZgt8XJKCTZxq9k700clNCWAY9bKHRGh2CdCZ/Pm9uz+FiGclrs
xIhXZDbKJx8xKpTIiUc1NlHhW7kWMlzDtRpcyUpNlEG6ud3DK0eOqImGdePvW7pevS/JLAuaeijc
nfftbIC0eA/AOTEjxqskSWbLA+4rZWkDF8DZU2ib53vU8HFaiaNpLac+G3gAfkulm7hFMiRbQHpj
WFFJu7jYGQXx5if26nTSyIhLRxNPoevcZDLnk+L6p1D2Vr6owuHm0b9kLrI93QBMt47feWBHieT0
ePo/DtGe0s6ONLHshbcO/kB274mrRbiXwjfLcikbZ1AX/FJYQxsFTNkBJvX5gbeqnwsw+3R2XqrD
y8EKkKY39Ol4aeyzanvbAIvXP+n30w1bNfHMnyrL9OTAyiNAwLusu8qG+UMVUxIQ6AMWd8+F6CRN
i5APP6358EWsMwN1Qj857FtFGNgzOVUbCaEzNk+25X9gESdlhS7jF980OTLtvha80jNJFE72bZZr
1IS/7D6L50kpfkAmiHbpQLQVumXUWcaTRzQENMm9F+XpH57Llnds5Jp8iiEooq8yWKkdaK+dw6bn
0tdOyoefh5kMqTGNdR4QFfsRvJQaTpgNbRUdPvYA05QikixUJ2s+cZrceWpbPNUYHnHysaDRMoip
Dk8/1C9eJ5ZsxHjJnmMZWzgO0PyqTZ1Kn2akuyDTs53PDL6PWkUonVbytDzx3hPqIwibbcSDGjbL
V+KFKYlVqdlK1GOn5Y0Xhb0Lgcrw2s3d/LPcslPxc9Lnj8yMBI3oRVWQ7jTZv02+baVA8R1spJ7t
P1I9BzAdn9szlFKQwkQv1OSdkcIIGE9grT9S+NXSSinTTouIcj1/Uvbi0Ew0fqA46sNq5HZ4Tiuj
Wphs2ggZt7RrOlN9HkpZTraeQmhQlakco3+JWJ/sYAVjnBTAnNnWSvbFhFYTBFuJ66HZQ4WoK6P5
vKP7QYPDa7nwgppTphEDXpMlcgnzCe7GC0xcr7PzfQs5b3yjIv6/+LU02j0mYekAk6D5e8LlNcOt
rNFGdCFVZr+D83pJAYpCkJLz0AOAWNNoIzaXH8ux1Z/LKUPchW2/jiEqCY6HzMR9nIpfJSYy84xk
FrXmgVTg2DZaRkQnZgUqfNXFYIEjSQrzQO2UcQBixVWJI2o0A56BSiVioacVoH8vAKf1XZsvm7Lj
/PJEwZkiQ4uFryRH1DXVc+qzXE/ZNjP+qYoYoGspQv3Ig9WO+ySO+0ka7qde/m7aZrxfUK6JuUgF
lKAxEAxcFUPYz/3yiXC9JTwQ09D6lpM5SpAre91RGdFAGJ38Ry0vKbbfGmZvkWs7oGXm/kzEBGdu
PLtBFk9evnFw5S3OlL8tZktVkhw6C8Z/2nNu8GunKcdwF8OtVEZqoArgP8gIobAZiulMBouKmLOY
fu8rexHsONbPnYao4H8tD+kW8rTcRjfErQzs9r6JPf8Z84kB64oJrNw1CvCMs8T3To+XA+6JpLpp
IdzO6D9apanSw/h6AiPV1T6rp883Xk6nEat+wSxEWU190Ygq+ib2g6K+eeqf9q+EH7iQ7qqG+utt
addrcUc0hKZZQc+ZOWEUuS9hKMQ5MG+JJQ7ch/xAEnofYqH3JOV55jB81+KKHKoSUKfAdZfMkia7
s81L1O4EyAKvpMKW9gGtPAKW7R12ZPTa9axuGsITEoGuSBkLJCXZgW4/iJ+bWTouBkUfiEv0HwJz
s+XFE9nTRQDgLFSybUIjkBm+qNWMKnn6ZxSBT6jI8hxBvwuoQhTjv8FcywUgddFeKZxcfNs4JrYB
u+8G84VtY1ZOm16iOj5Dfy4CPLY9KBr6SHy8AumoicAL8rAhrJ5bAsuTNBKI4vYrmTHNEaw0vyvv
m7ciH5f7v13wN1H40mIMfGpT59SGM159O7olkoyBq7SX+2y0vCCO9AOGNhFzsVfTlbRLP0Xxj+td
Q9Tnjf2j7c/3VOEifZc8gJQXJzSz/caw95JZyhX8kc55UruOqcOS3XTbrXchUIooHyRK1GADEoRW
qd8fUeOfDOS0THOuu4U5SSHxNk5sfiSXx58/ieEohIoeSg24tUYA7CXYq+irSHaj
`protect end_protected

