

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
ISK+8BrzqbDVc2hIh4k9UuGvqsq6yFic71tfszsK7KRf52jFUoK33AosGVUYsGH1pmrUc2NUQcDQ
LseNrcojiQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
CxxZHetyKRTjg1ePIJzq+w/Yg+inN7g9nkhYUjpPSXav+SKIAQvdh174FZUi0SnoR2INo+rdZ3gz
yq46XymO3b/3npnRNCCU259giTvnOJxmkrtnjRyUpOg8jB2jnHg/f/BlL3OJUGGiFonBs+6rnNvW
4aiU6ycFpLQsNzqRlAw=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
HZ1Kttz7DNn3t428AVZ/hrbCqljpJfsdfcEo7T7pfqxl88ELioDFFp9rVcvvZiZMU++45qS8CpOD
SfwcEjOj8ndwnIsrDamIUHs+Qm4vUDDq8EtyiGhux+pwMtpg8rH6kCwLDCkdk848fWRbBOGctdAr
AiQz4Fie2ectzKGEhjERjquMNqkQkhNIuEu/CSTnyD7KnG+FK+llVBavN8lxjWeDvk+quMyk8Dbo
gA/SdzYI7TCZkNEFS/PvF3Z8fPBK4pBWz7TyfdHacMjMkaPd5zGsPBmQy77xwc4m/sfhM7ZX+YW6
VBTILiYtg7u194UVgu4fHE7f45jr0jTur9wbVw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
2VX2NPBJC/FYSjnVp8ueqtxuxLgenRIKbrff8tdhuTb77js7o9S4OVH2n84fEyvr3hl3lrO9ekVq
VvQQOlQBg7Zv5/tFAeI5YFisgygYrqeX9dQcI485CaCpeN9nanYXhtHWROH+ZOYckBZHUhhjC82p
LnYwoausKSjsi+rXE64=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
HdQIwrCqCFDZv9OQZsva3DMtF+8TwiePvWLQndNAXK/1V46C6C4sVLdH6SK4FvPis45PZ52T91rx
x7mjaMnTgTVkK+VoFF3Ej7xzh/2PoR+YkiToyHCbvwHQXXvv3GAu3HyqWx9b4oOndnrx5Z1mco/s
lNgEY825qOfDqrTkPvvNBXThybVoOKs2SBHAdaQhQemuYVAjS7mEC/lA7vom+55/0dhIN44Q0vMz
6utkLeK9axPmrUz/LHNLm3BFQsfvacsQoIQe/Y7g5V8ehxANfnzft/Jgo74fJAU3odGS++0PsHF5
2T1joNptoFFljB/U6DScrAB2FxigoQal7I/OSA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4112)
`protect data_block
gBh83+TF5Spu2PmybZ5pLytJYDe1Kpb8j0jbQnr9IA3M0Z3zl4k9N9Rh9dB388h7DkxgPGbiFDuO
jJUxnyTiAsBHX1/z73ZyY9dnEAewvcqMLmio/0/YvcpziKqnX8T/KgjBVjYyyx3hVqFbSHHBdPFz
veatGEo2rQSaHyLnaEKhC4RsdYcLIzoWv6xCWr3gX7lbPEJJ49miG8rbouiLuWkfaG+oB6g1gzPC
1FeEa3ywnuW/iRjqKVuoygmqSMOpHKcsq2tOvYezCz/dvFlx8FrlrOzMja0/d8ttAgap8UTqUseI
XgDGVM49eEGk+oUcut5z7aDEDksiMsT64n6NM8npB74s4p/xFAzb8eNU+BrTGdqj8GlGYVJ2kaNh
xgeJBY/eSW1+K2YBlRnnlkXG/CIoNsC/LKvlOo+3kow0GVXfHBFhSBuw1PJi/qN6cGQg4mCITwOS
sez9XhskluYj7UvRwVjtJnxIcuh7BCHMK+A3hi03LfQiuBvMgTPCc+usfNwZGzQqnEW51lCW20fk
55vffl27AcCaXc4cxtie6avfYyjNhE+kLdcp/P9Tmj5qVAxpOyW/q5Tds6HCKc8kPRup+j53wVUi
v3F82RRwWKv+5941ELP8mta1zatTomoXo6UCqCKF+llElqnpVi+F61+0ptZ0PHd3Zh2zZ6n9AAb3
V/18M5+OSZzm+0RuC4t0H9bpb0CZVLXOGzznGP7o98YgIzZcHEBh1+LiLECWk9NrJ248I6pIphgU
pVQWcJTvdq8srEAyjuhdp5oxFQSFdtDei7SLyieF06A39Efs3M0+T/X6Y/hqZ4lOHd1uLBKLqdTA
sZYpiB5Z8JpcxXYUlYO0TQN+/39e1bjzqzrB+5JsftJIw1NhkOVpo7ZiARvgQUniND0zujvZHFdU
z1KhJ9/EVi1JLr/0iYZ4BlfN5KrUYeXKXunTJfQzJEx/usNzINz6Va65uC9WVPMadOoj0JfO8IQC
B4aP/t6mQsxDD+/ThC2773tBMHgVm0UscB5+kZ1N/VECn2ck6f/DC/YnMhtS8X9eIbG5JArPZrdB
VqDI3RbvXwGzJHnEHopJ8UiybqLupvTSF/zoqZb5RtDnMLLLoQkHmYfUfHZknc+bDksgrzPdBCiF
Q+DNt7WxbzSFMZ83dO9YNxWS5tNTJRJ9DAg6k56VE5LtLt3VuT2aoEax/xCpLNQyT8uZ5T6GIErZ
XmP92/DUKUsdZFAWh1or5vZ/gjlX0SQl7jGPGfaGuX2kd0TjzI7UgLEBGRHccRIzcasWCmeYH47N
GfnVzJcjgR/wWrL6euln04nwD6VQ0xjYEus+O/NHShtU/0G/iLd7QIaIrn2sqsTmjxUg1msd9I5C
9R059Hnpf1SXZ/CT/tO2T81j2OHLJgT+FFz+UXMsCEdxDqTsORKnJUHiE+Nv+lvbgU0kgIanD6kW
wlXJzOB5Co4SQ2TowHvdSNvvBfdwuyJTgkjWsB6gW5fY7afLun19WDfTkRqqiOkDf3vg10DVZI4r
Kj+XOEIlFeDm+TqaKJxWVt3DCnKigUF3TNmqxDuCRxYIpK/Npn3/YVpvjaf1SPfGWFYDJZZf131T
bCFTry66Zx4NUl5QWUET94gCjK6iWRpVW6n8YStdE81ttHq4+KCUktDWE39uXFWehWjmmz4+Iihw
AfaaX6wiLuvnBSxon8YLM+IVo22twHO4afHWitjAJRidhcrovEL1y0Nc9CDe/PZO5tQmQd5KR5Fg
g7tvOYsmGYfx7B6FHwI0PDIU74uIAmAFAdzDSAYdQmFlp2mYd+fAyLqsWiSH0ZzZM24or2bl9TNp
tWar8CwxQu1I9wbOg1voCg2DELoWRn1ZvqaLpghTWEiFBVWZ52Vi/MRch3Xldgtj4uRsJ0NQuP/f
sqA7vN02ZYgyt7ykgrnYUhVXeWfd5GekLJGY82c5KuJCWPJzLGZnguF7FxeJa2bDn41yH/sQMJqj
CgYD4FzE5zQ+1URKwOkiu2FnmyIE8RhFlXp//Ov0pvwgBMzroZld4A6QYm4tF0cAebj/VAxAQPOM
3HUHa3UeDh+3oKt3n9iwQ9ETIu7pebZ7LqUhtsEdAK1kre9X0vug7isTgd4rzwpBb9Eq7YpvuyEz
mkCabgWw5hs/z4NXUMJ7v9ecNcJJhAe0d45OWrBlw0Y5NwvTcg9WJ6j8FvEnZWs3GDjpMqKraz5H
x19TB9vQ3UGUkbLAt92JGh0FOe6sQsx3drIlVzeT2HtASVCWehFD8pB2bp3Tg0OdVY/8gFYjl8By
Ebq8U+Fi7Dg9Ls59TfFyUw4DU3auVNd22JvWqi0tfR7zv4DIyYyGKa/Ho0eHurFTu7xa5UpfxVPL
gHrETHlWBw5Mq7w/FIeVqQPlIEyTeBd5WXsRm02aHDMp3UjeeOR9hE8GjJoqpcOPE0S1wwAbzsjk
WKkKG5y6CfP/tsnlrSAjc/ezqxGsHtBBqaS1hbXepdbwo4+PpbjPQGneNIRiBq374t/DWN8NBAIS
HVbm7JCcD1jf/Emenj50rVg+eYs8nTUS7TSfJ/selIHArK/u9uwR/q/SoMaxgOI6PrBZ2d4lhZ8o
txhLIt9ZgRv03hp0htq5f4vPOps4Kms/qkSEiQG0MlJdE41j1i6KawO50AWE0PUtSq0kbpx2RKQH
wq68Nce6hNxrXy67RlBb8WK1HkZLk6zqxD0R4zFKxA4BnGtUtzSxBeG854XdsNIhNf8jrjB/nb9B
EybVWIG2Sfxwc5fDyDsEaL1ScEmMVFbDSHWbIyeObOnl2AaK2z+IHBy5jfH0+MBab8szc1cYhOD1
IcyIFeAxvvJhV1+LY4l7cWbxYf5TfzH/8p3hl+FbXfAnevFwsvbOVRkjaWbb+/+qCuVYk272bzQu
eD1hCd4qq38ngeJVCaibEFVKV1AMyMp2UTIQYjIvqGsKV653wjT4czf4lwq1TurK3CbfYUn60oBf
OrLpRgobimJ1mh/ExwkqBcZXl3z4kbWdFmc7IbJzbqyCBt3rYZLOSUlYPBhCLR0BOUVOYlgOYYaf
FHL9v+mbbiE2QEGlImNFwefwPnEncaJHIbyLR5thtAYwP6lvAnMeN5Ot66qeG8BQ6QuxeNGPBPFq
mkaWGXfTfq4sms8NPqV0jqYmKYhc4A1fBPO88n2n3xJlCUkL2wp6hlNPKUR2ba6Dn9MF3F3CPCD0
CS1IievP/k4rFzfxacojy120pLXt7Gl2ydJqQ6AUuoP07+6j81vWOO32ynrITkbbb4366SpfztPF
cHw4+vmhELr+OZKImUwHb8BjEKhl0vY3o6jKnHZdJwm3253Ddc1dhHpJZL8BhilPfWwGg5WVxiFK
YWr8BQXVGGCMcr7WbUaCUzPeqClFn2EoXpK3fYxmLkzbJtELXasdq5ausMgfjxSv8A0WUIqStH6Q
/3K3TwcrK8koV5bLHTz7Z7SnHbpwcVCgkx//dr/kU/7q8hDjlh8gYVTM5/HF3tiC154WZjQX8ltf
mzFCB3y7Uono+zvukN+TsWHIz7PMBX+SZObwpyLV1vhvg6zV5BtkkykKGr47kMQjIc4D3prmbkJ9
rNN4X3d/y76GnnAqCJdsMU/8w0Orc4D8BMhc3xqUsJDlw5WBWw1R4sgCerGYneGWZmY7z2R7cna1
scdgbTaHSkmWB8AVlzLME3AU1Qybv/rASYkIX6slv07JGOWTSGTf1/Z/kNtAn5PAuKqbY/kTJWFM
7lV4m6zEnoNmrlJcziFMSMlKncmXX2K9rpSI/RWYFoGAWJlTY09g+3kipWg6YglyzgwEpIm/JeA+
/FQEa6OwbEROktf05/DWR2LxR2QF1OjfYmLnQs2GPRnAeP2iCxo3OrrOc+sp3htVYxBFn+Y7SRFU
dYkm+ExoN/4+6blX7+www7thTZqXAD8ldmmu+2c22lkfDaruVMG8M85oGwwWXN6eY8AJmRKfds/7
VaBl5wk7jJk04DwI08Ua7Zd4bJn8uXgJpQIaRwcFMeDiQQZTAsLdeGnXVdCGJ1xts5wGYi//IcGn
Pq12upbJPt+3BWIrXB8hC4hgSexxJll0SJ43pQeEcV45/5hvqVDjBV5xLJfq1+q6+uBTE6iHSOPs
OCwMBiChjgNwACX4H2Btgh8z7xYLjgwJRePtT5N04b5JjAnzLLOsug5nwcS4JLe48fz269UUAvKg
itrT/OnuzRopj+qE1tvpbaoFN9/NS0lE3yaV7Vn+uolosJRl5A5UZQef6KuClOqwofQVtcSlZLIL
Kpc47P6J1a2hfC71MhD7WJwTZfuNSd/kQN9pf6c79cR7yrPUPZMWFoOEojaKImirXvQ4yd+5B+WI
DQMp8B+AYkbioHBkIiJxKeWbnc8KsHtwCQlq72ombCjD1fncNVaVfZSqxcW5uQOKj1muqG7Gugjq
qQCHV9B1damwk9UoAlKqw0HRcHg1laonrHzTxWUk05BInqvcR5Ajiek4Ne4BVxfq+EZIkHVx6UVx
gkr3BDd0GdMXcHnZ3kN+UEnhDqWDjUgGJlBV3hFf/G0oP90h2DFimPaHMGaLfJAG4IaFf7kTHz1c
/OuZyCZjxkO2v+Dld7R5hpKChm7cFFQLJEloa5ulrllapwJJOCQ/Iq2B25LmzZYD5tSvfetMmf3X
H6cF+zjBYjkHHU8m/JRUIB4mfvosd8NkJYIi7EZPR7BLyktgAdDQFy9oxvro98RmBoUqkva8Ais+
mvSuV3f0fStzgX1WoBleFxihHF0vQYCiESlHtd2Ak0ZSKJcoKVIPgvHEBw8f0P2G3sT/TTUm+aVt
9ZSbwsTGw6O1xnevK8OdVT7zl8MQM2QA7dKdtTYam2ptfq531wQ20j+fqO1hxiKRQFUKA81XulGi
rHYdhBOianv8RmeVqyck+TorHjEBE/V/ta0AZSCnxQhbnMzU7Tyt20sCXEAhg7b9IHy2MnaFx9aD
VZlMERFHtmlJAF9qdhYVYRDoKCjB1b2Cz9Fr7faashXdaijpl4CWV+iVtMf4u4bbwntJI+oT5A0s
0qQnl1p+jaid2GXEDYl3HNMTO8HxU/YkxDvD23qTPOt+0Ea7I/LNTxCvZfVvzTteu1bCrNOp3E/E
nIgK73jN5xzma1PMspOS32vwHW19mkLHpgffqXv/0pTn4hKncxkpe3gaM0PTPU17wT5h4MrvIlT7
0mwCJS4f5GxSWvkdC4CjUxsbHFVwVby41VLRvEntMWN8vLoqZ/qhZzVUiUj5tBiYr/hA1y97JAEU
MX+9X/9fO5/79d5yDJajX8KSQhoCzmUnVqhxPc1kGA+ISVCvWuVBm3N93Q6pFnt7qo9xcCQ+jS+m
PohZ+qxnJA+Uqilxj1cmkLv7ZTyw0x0U2ke5bGMoSWQFU21jv+3bZnApoevYdTrCYWgmFi+tDjNB
L0rao27TLBftWdaoWHOPIkQ3lyjpeSHu3/IttdG/k/lD+zwj2qD9Fj0lruPp4OzBtTAQqynd06vQ
XQlWGTOYYFA=
`protect end_protected

