

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
QA13xX+R/ACi8km79qumYiCoL95/JTNXmw/Mv/Sollu1nSewLnwk6qQvytLuy2zqP8g5ZHUfDkXy
dYJVTyRzKA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
nii8tC6PWRY1wcl+Yj+dJQmorGaa82N6txtyUcQdtmyxn18ohe6n/SpcWdMXBCN1HiV+XVlZhDEw
KvXEmx5H6nBr5/f6eVRIc3k7vZjXpluRFM7lDsLgIpfE0fW00UnX/0rMYgmxn+5+4dG7smGpX72S
zm4Z5q7tYiBa+z76ex0=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
yppU6wpcO6vEUEaOZTTT6jS7XbaY+e5Jeh6nknICBRlkmT5DzQmd7eWK0ShMWSlNt0Fv0kuxSdt3
PRQVKoJayZoHlh1UH0U//6ySDV8PrR8ZKYbnb5G7lC3+6hAsVS0WEHoXFsxe3QTXWezPX8OXISSE
YYTVzXqeBUtBDqueK1cvQyMM7IWnXgyQ/0dRh7UmnEpiOonlQALl1eEnWSxVZ0L5cd+jDbcSlWqj
VgoBh9A+IbjGjOjE8FOaFLUMzvKXmpjNiGzhwyN1qXczrRlE54AWkRUECVVEGR4zuEA7VTQH6H/B
e1HQhNsFNtK03nDJRyhoiacaeHGOBo4yneyZRQ==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
xoEHrB3Q0Yfcf3MYYTBHkrbmS0WN00JVFDeAhGuvxPP5kv5812Q+oIM0e+z8RwGLEwQ4F0j3UPw9
LR04YDkbyd4XfjRJQED6GhUyhlVHkeZ0vYn6D/hB6y5zA45LPFz5aqbLudigfR6lDZgyof50XSaT
wkqaJ1dNbsbYXDGYiiI=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
SZoZou8zrLQYkyuoYxGz7q7TKCLXDf41gJHR/eNOYbjhVAUcJLojwHpmGq29Knnj056DtiEpAnUR
HkNwqIIUQ/PzBp2ZRgLcYUhgAGFauW9u5fA3Qe79SJmVAKU55R6eP+5h6YaMx1oo7Myp8ZHgv9LK
0atkww+rNUFhc/kS4ivaypKADJgY/Slv1X55We59ldg5OMI3+jFcKD4Ow4Gbs5tHnIUzKQ507yjR
1wg0oIoTMEm7GhN3wZnee1A7XeomsW7IrTE+3/M1cRWhdrj0rq5nqrI9yilbmzqQyqntfJK6N8Y0
QQNZFJ8oCjr3X+2kFBb+Pd3/scpZe1PtOU8TgQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 20896)
`protect data_block
PtM3xv4vSWkzUcsCB9exhp7HS8LX2LkaQFx9Z4DYzOZa30wQ8hlurUPHPTdz0lrOLD3JZNip/fWC
iZQo4hfAHcg+2ICBWVbS8fu0Qhtwa78NfFJfTEGEUAlqtrLmLjwr2jCt8wYf/1w6N0kQSPkwLfbO
fgLFaQn+/DngNCNLAbYkBAhh9Rw0tIrboPxvkeVaTTD3unfvwhve2EsFejpL65BgNFZ/87bJAyMA
AwQ7l+M+CCjaiLxeWVeLZHhnbpq2HIoT/xZB6pUFSM0krEqtpa8G/sS/YLY3Q3U/TLBHYad+8HwR
cLyeAMvQfVKdP6i4OR2mIc66T7ejCV7W5gy9UAcbmGCMC2WFKvWBswdPtJpRBH52FFnV1mDGARzR
cS0ey3uECF9Le7zYdm2w+OO/GSTftcRtGlQFieqpc9xVOY8/E8P9rKp21xKEyfBxepm8O+LDMXco
d1SUlPqGa77L5r07Fjq0wT8bebQnunBOars6E2fQ4sSiTr/U12iEgcKBMFOaahH+DYGYXhN69WF9
o1oq7BJGEd0fMVjiEqkx0EsiYr4kLdYE8RU4l7RTK/s9Y/Zz3OZlUSE2waUxhSmCCqHGuhvjwSPf
YYE/pPmAvc28aUdJcEwLdjqwNr3ekO4Jz8aGK1IZIfQtj96QNWo/mK6Delxib3lYIZNLKh2YVe23
DLNKlpeiMVAOIo6unX4dF4axdR+r3dN+k+Be1pCcD2De3B4hL4TR8aLccHQLuW//AmnAwvfTzlrw
XwpfXr98sKyoSLFsA6NaCI0FNahpF8gAT++kJs3HEWECv7s+kWjNWd4mUBUXaucXufd5qFkqPkCJ
EWRYoLCjXrki9Ka5WhwfmQmIYhOsEl/kGkk4RQaUdA8AZ0b1cep9OItwqxI8zHaKqxx9wQ3PY4Hi
urv2aS+s6EyWpB/ExX9Zy4nayQJj7bSLx3p3O0MfOp4SLEpOaq2qPZH1y1FpNYUn5R8Q8DDdhFWq
+mgX8T4NcDkS5mbsII9Z9bcWRZ26Pd7OcCuRwSlLwMPQV7U/+DsKXo3tcNY84sbZO9m49HczsBe1
wHxYbaHhTyalEJiRxiL1SdZqTHC2A+5NZpT/Vq6UkrCOZCYtr7AMd0c3eetjiumJzjRdsIkiz1na
Ax6wT8w9ThGXgl+xploKHH+AZxzMlRNkWyMthHTTlU9UdEnE/AOKqygiBQZAoh89wA3xEZYiOs+L
DT/EAqzhqhRtAp0SRy+qTwfvPZmWnaZU1DzAqukEAz3TMr89olB5I4520bblARfoxiuR/4T2wQ8b
mnXLGJTJdhuOtvg+GZu39djwuXSeSIJfSee7A4pGxpa73e2DsCKR+3sHBtd948KblNCM8wYkTlCG
dgKX2U66irLlYWNVZZRyWxiYFLiU5/IFMqdRMFtRZcN0WTwxPcjevwFKsZQj8QrIdjVCORmIP5yV
mhiGUl+ReESHiv63tSVYY4z8KekK0EAB4/Tj7TDVnSw6HseSnLR/Sc/nOzvekV4S0EGh/gK1WKqa
URA+AbIRLXbgqacf0r0UBfmdd+8LE4AeJoLOl/EVZJoWq+e/Yg6ti+Z1RosIfFQL6SAeutn5FGBg
JAhHqYnnHLlUNzQWFx8OYPIBQEYnHvRhWnyeZenLa0NOsN/202rG8TIrm/rZMJrjdKsNQw4GNoGg
NnRfg1OvYzfHLFmYc2cwS7GDWSaWU2pcwHXiOhBWXIfQwJw8mYXPErA9Z2c9ZJYFUQW/DPxpAifD
gNR9lhmVgiAXL7kx2Qth9lK1mwHDzKBccCKgKAF2+HP6tWwUT2dW2btUm8mdGJSH50gIHtmB7NOv
+4z4NwFXGYWQXBtyvG2HioAtHky+kHQGDDwDL1/+TZ0Q9lH3veJy+IPe5smWN/PDEA5VV0oWDcq5
bYZQQokWxtdNIkA1j1uFob6ahApyATxzPkkVxXBCfDUXxIM1paFzn8KzZ1tuExw+Nh9UC89pFQOD
OBfWAgmR1hI/j6oYmzF/H7FECVo9zoq8w2kyoRh6v7sys4IbAfEj4mS66h98x5D+aJERgLKLZUkV
cdGVMF1qEmoBqL1VDv4/etxJNqqLGRBevV7PeypK1/cTmKH0039Ga4jSGq2yCGuQ0+nU+GSpRcXg
D9VwE3/CCJCYGlFo9Dm0CZDPN3PHMaVeWVozfyyTIRebw8P3c3tylc80J9E9t0xybMNm/7lbvtPm
uXgFsb5IvgX3trqyicM+QDln4+I6FR1KkPu7fFC+AzF2dqSeDyady/3cwqDINsy9VCwPaKWJ8TGN
cnNbwRTQPp4hH1/ySSE3dK2ZXQIuif5V0rPc5+ik5NB1EclryvAXHbxiirqBNE5Vklm55HyyvVq6
AVH4zDxjGhq2OzfZ5mnhewkbnZjASR/OiJJF9gErQojimpvRZcA8JKLzQfh6koFCi3QjxnPwkT+Q
uSOemyrsDZRnt2UL9ftIbah0bpwhMZ+8ihAKvKBvKqFAgwI72i5Y6m9kzxNtoID5StbAzUv13tz+
ziwQGyHNTUgNOQxfrGuCCwTmHkTwcRMRwfMFgQ1uPSi1mphGx4bjzgsw8/N06TVNTwbYu/rrYcQE
wjR99dPqqqs88BjjaN5by5tcoCw40HLccWngI9JRUVjN0fQC/7va1q656Ls93iM1Cu35xUnM3oo8
yIOv+YOQojmGyBoKnMl8sGt6O+jqqtz8tnsjyUpkZFhrE8L4MI1YQnTtYLOh8HBxctfRzAoX4Drx
Ms2rKfuiG8TxlWVln/5H2enkm1PDStzuGZSv6Z5Fw4RtMwjrcgCNL3KOIumK3ZuGngNddR6/eP/L
3Zr/Sgt7/gwoR4Q2+YOH7KUcuzDfDtEa/aQB54NL/osbl0mZC5TU7I85d2Fa8scBRLhba5DkQ+//
EQ9BGwyt/FrGETg4aZz1i6sb/kwR4msjhhTA+qdLB8yLpHR4vrW5IUZZplIllwMcS/sZreg52icx
aM6SGWEYVZqoOHoj8sJb9ugt25wcsCmiveanTAFemxU9zL48ZqE7SNLvTECFvNwtvd0ZVbb62rER
6PkkS/czz1WWPBs+rDEYodMReMIOFJo6GN/h706L88bAIjKWMn/CU/teXozmQgYrzQSSAlTdJi9M
zZL0dZtz+c7td6dCcTl2XHzy3rTiinn4+N43K7dRFY4Qbq2j4izo50b0wfsSh9qDEmKw/KGHSxz4
RjkGL/2rOsth0dx88cx8e2/48RRujjbAJ2DUQe5rtmlyMocX0b1t+4UnMjxjJLqEcmAEpDiy+WlG
kk5aDrKsQ6HtgF1WA7jpB4wjoWKLpDM4EFgejCbAOtQjVZhwaDGqPmZr9Ah4J1H47lKHOgraU6AY
7OubkKb1SGY10gTCLTvHXyyD+tsr/I8eNQLXDMg1S0JCRzyue1egVay1VeAlWovd2pcDb1dyqq+o
OnUkw60ry+WLwmdjtT7XXlXJQUSupK5/rdjI2Ddi/QGfwf4DBvk3qAVmAZm+rQp6lxL3hPAgBDk9
nCG2zPvc/5+i/RNvbFdS7bV82sI61GrlD/3k2a9W4BbMmgINgx9UshvB52VXpFkhWgcYWRfnb8IW
XF+DoeN3vwy+0lkmU2PkcQ+FU/jybjSqu1LqosvX5SGeXSeASbkRUlaOcV+cpYg2cOcC38I/4rtk
0Rg1iswNbj8eVoScMz2fVHgalxWeC1PKJSu9dcvBRYGpxmHYWh3C2q7ihmlTRqrvildkOK5ifkw3
PYs4AnOKtci5H6URP7b4IWbFXP7uIV67l2CQ0XJcGybAvgRoLlGAKgAfok4ffk43dLqfZKXi61ne
92LkHukn5Gs0LNv4qr3QWwqOVwoVMXZD48QVWJtTAqCSAK3lT/Tbd5qE2VlxlLDXlG1US/Cvtgeo
8tGyBnF+FjZBckxHpQvfiwZ3X6gDsUiSq0Avp6PQWowg1jUu760caDKwVy3zsWP2aQOwLLgeyOni
NU3PE4Rq7POUI910g1s8dUQqJx2N4nnYd2eOTqghNgc7VYBSF9y0AHAgIap7TcNEeETcAldDlWRG
rUjVfOzYAD2iqZYxlSrRbhT7HUmQzLiIHplm9ClM0lazv+C4a5dq+FLnxFXQSMlPTf7A7PDfZK3q
5i9ZpjF3cxm2qoo61Z8QDRypb2yzCj8bJHzhu7pUVr5bEHg1CTxFs0/wU4pLJRdLMgA2SG9Qcsl6
E0vAqgA2b7sjllt8PBTbDXd04KqrZ+TMlKqEtfOgzJT+Ka7kM+7WW/EnDNipz0W92m0JfZIdkbC3
HOlng7Lck8rHRwx6HFzbNcs33wS8qi8PFef8HTnqc20DoOPeAZFJWHI3X4+m1uPikuwSrRBdfmu0
IFxxNhNVLv8/eHV1W0vUkSmWWPCP0+ATe01FnMjhJA1kEw1/JZ0kanyxSif3r/pS/LZ1ZkrSd3BU
GJLFAEWSSvt5neyD1UK0ev3xtrG65q5Uk92AtQDkg/OjqbiiO5UUYZBDcdYu4NHdYUxG3xCa7hQO
GrnT7gLbQlVjoKrKDja/dFWwB92nv/YP9RhiwRxBd+mpyPuIGM4J/PTRFLrr0JDhCroC2S3BdSSG
qujSEoJk6p/gP8cEOJqAqr+5AWDGpKLAfj2H3FJHTGE7OCX1ZOgyutm4ZPh//uzmvm1p3nkfSHjC
yOeX5ve29VFI47wLZTitp8dgkKQfk2SJoQfVspNu5SLh+uO9Zgu+WQnEZBcHV0fiRn3Ihqp/MC5r
wLelu6cLGfbVkl6pSSGA7y9ZUdPl3tjlefEkY/t+UPGaroCtSD4AQdBD9Df/rg+2xIv+Z8udBdW4
p4EXJdMRSkOgpuvoxtUs1quyAlDn2BXDSMV3ypHPAcpoVc6CicldVGTIVA5RPgVOts5FMoSHg6Te
yYnwPy3PSOW/R9HQzLp8r/a3kGslQo5gEqjP57V1zJp3CRfLuBD1iigw1AgiluxdxAgnHHroq/E3
DYcmHD2INSBx9RuCx1y3IKyTMC3wVLqTmjyvJGvzIm23+Vv3jUQPzc1se+dKB9n2wsHuS95T6DqS
asc0QSzqNOKDhD5mxKbY2QWzMldXTb9zr7b9OzBrjh4gmN/bOP6F3OA8Tayuh0ybHdYLZUGp70uB
F4RTccnFXRwxWrDtSTiKUcL+++1mhbcsnB7GxfebWy/AHljIZQp7CkW0BlC/JWTC1qAeBarACfI9
pnLCrS+h75wiCDaYq8fDYymOPKVPtnRIrSc6q+AKKrwMV/FWUICOmJdqILEgj0kPsmrg5edznkTR
pVtGIxDSGT/dMIdc5p3MhGjLwNCXolGF6eB34YJBm0ZQUJ5u0HhDV6dQehplt6Sv0OvQm87DFlUd
PyD7+aC82VSDsSzjQmUFp24u2aU1+gi4jXKRndxOODXO7r6PANgcZVKStw8/r/YEQXhfDnY6/3Wt
2RCls0PKcltaTvgwSGIRDqkKqZnWcSNgeS5qEwPTggkFhHawauB+lXREvLSUmTH+y6o2eoFe2wF5
1cWR3GEsK1m1R+RGe0kch1xrNXqwXhsDCV6wPPqaRGTkWrUjHvMeyZzUSiHggXJK5GfXt+PrjWq5
WnAEpBh+3JBbeMJ7PuYI9qsLzVZ2z1KvjSWN9j2gVlPMoFkc5mPYr83n1Q0fNK+hyELclBQrhTvr
+UWAhrI3luCOuIVS9PDgHDuK+B6kE6UZIBwdfvJGE0AzS0CwfPqRj1vGkrr8pDk6XpBNYiMsMSrs
zuXzC3ijX7l7amtf4DqHLcs9lHuwvlOQAlNOjto+DnZiwcBxa5e7WqFJleQEskJh3bgbmjGnM4Xf
Bbxz01tdsaxIvlSb3KvCfoVOmIeAPQpZzzC8jTXHK0SGO6yTsWSz2NbfpFMLpA8EZENpC0BoW4YN
e3FoPc12lb/+X3CssEh2Qo+pw9EYoOq/J4uN5vGgixIqpuWptb8UksvFyTQ/svNI84Hj/wYVdOVN
tGSMTavonMunbcBwjTVtTbBRZHmX65B8sx47CS5RgNrYhUMkRZm9FvgS8AEkIXo4QFiTK2xyiq0m
IO24kHSNUk2GtVqoa06so/dsPGks3/Wb6qYMSb76ZlnPIwByhslcXMq6IZq4RYF8cpzt4q2jqjjH
HLF/rqVSAiEU5znWQHnJYPRIiLCVEbpix7r5kycl4EqQmd7zqBfPmfIRpQwlgJVFyeRIOnPGvLz7
lhBfKkSL4YMNycYxz4BhhfKTikjq76fHdjkUFFZV+PcEbGSlH79N8gK6ssgN0UKGIk31bxdbdUhb
L4c+NZR566TrWUvCHlA2MhkdUIohzPt5o1x/76UVsucLR+5ac6QqL5Fvg5vwfTbJVchgOaLglxAc
Bt4IgXYdPGEE+QqEmO4FfKJl/VahuZj+0z0ZURd6XD3ICwqmnpG/W3Szec6ijY4r7L1BZqsAc1Kh
rS0KvwAwUp3OUNao5WWZDJSsCf1Zn5vpfrmmdzVccJkNnIxwrVBenB+okPWdxq8pi8Kunz4vPj3T
638xfkXdAaihRpGTfuVfoBSZDUX/WkWqM0t8Zp3JihU+PV+ZXgt01R06GTXUcJlA6JvtYv1eMXCj
q76QhIUfOAIUDNAb8Y1ZuO1fSaebLi2UYzrTx8ik7WlmOYia8eMYQ5+BH/B9fedGq3leOgoI6AAY
LbxA2nltTLo/qhpp2hje2GRpB01+jJKsE33oLTrCtBFVhZY7cmT/xbuB/1kyCcZjYEFCBOje6+x7
8S2np1aMbApmDH2lPVDsIPJ5IMvetoeArDnalkfDPZ/9xCgRBJt63jXjkRUXKbYzgJCwR/PD7kY4
h36xMq8rgQClpVc0020plAf1eEsNDkUYlo4vu5b1u7q8Q6ScYWNxYHpQyw+XvJqzITbvo02m7jyI
ffW3TBiGKi7gebxjoru5D80uQa1e/hmClYrCxQ6vVZ9Jdp80oDMrEWmiSOrz/DDqlURwTAVYKgEg
iANvuyFRojNnR68FlGKozUJJ4Tj15ipq/zo1ZfRcQ8iFwC4bxKBM5cqg0EaXYH0FLEOxvxg/+nM1
9ZyRsS6+sEA1BOyoYkRWRUuZ17/+seq0JejTZX54fG+1pQKhF6zdcFngJP6APTNFwp0Nwvct5kis
Sg6Ukcdp4dMyWQ+W+9TsGXEJSrKaPikx6i0LhgwjxYB98XD4uhnJDvSiaF9Qj+2Uvb/zQ7D8gz98
AQkCGD+Q+jpIZDvV189P5igM1C/rQnAKXGxupfL0qLEUZjwCxTCSt2OFMolfJFrpuEzAwDk3RfIt
TsWpI9XX6aItR6NKtWP87Icl9vSP8cMUMv71TOO1wUK3M7oWopJNPJ275AzsxlhChNw2ZH+7FCzC
4Xl4EaIdS0XzKMNnehep/zlWoEoPaUn/csslBV6N1MiQa3YvidmbPJgarXedrxlJXc9LtSlwEqQN
8Xjc1GgpI1l21pxI9x9HtkKGuWcsVEZA3LihCr1r4OW4NcXm7cYFWzeHTMOymyA0d0WUhea+oVKo
ocqgSix3L/HWMjN4xjvdUo2XdeSLg6p2QI+rq09qBjBMaIUekYi8LNFTESCYNsczSJBNmCCvcJhv
OB7eEe2xAJei+LJntsZSBg++44AVUZx2G5Jibzx1jGRT/foxbse9tvEIiL/Brcvug6kt7aj+KyM8
6ANbQwtha8r//chNyUb9u8tmAPCOZ/FC6epIuvv6V3cQkhFqYFhTAws8TKGyfRuDC7iMk4NYObvb
7FlXyzyZGBjAGqHhSJTHUQbFXoGDQ+n9+2kKYtNj51MUvO4TwOT5uKlAAOmLBffEik+Vvm+WZDFl
sJvk32wc/XsIE1UYHfrMXv4exp+bW/nqnWcyGKaCY3XrYD3UgFqa1Ms2kkS1QGCOfSINdr09+Q5T
w3EHq54C90BZhf8zkeuE4DIMwQMuUnhYzN1K0z4zkjmePJguN1bD3J+pFskGXwsjubNWez232YZQ
qpPgKUSMP2T3mRhQa06Rj3lBBsHxb6lEKJYxSW9Aw8jZ06RiIPGwP+/IE8Qi5HUSnp0yqi5NqXyn
20mxsFdBjYlvnqwpD3TOZTTrFSWCtF7i20c9Hzq2V4sEbIWFC9VGzOJvqIF6Qu1zNPHyIWLIZPlG
a61amM2eNe9MMvxfMU4DCQBrtyhhYzP+7R+9rJcnnls7RqgHsyvd6Dq82ePFnVNM9Tk7bZUSXVf7
M2tVxeAw23EQHNq6EvX+pjVu2IZWDlML3NqTqJXjqYJLAgCkKd/R85Yip87IHxs/8WjTDu/ZhxNV
z1gWgYg6hnZEIH+DPA99UKmOJZ37anSWHl/YH57YF6DVhoJn7/sWb8suVg4gHDdyOvA9pCROro0C
S/PNYQIxpLxjLuDj6wInQrSDNA/iuOW4ivVCunE93cwva8jJaiRqytEUrghx0QCJVG8ozmsZUjpF
+cWayquNfIQKBCHE94ccZ7yNh3HCs9CHEwULrOZfJTe6TbVt3xC52NRHEPt1f62BHdn3KXX+2JKK
h732OE9+kXa7jIbPBvABn/CEzKMkgv+GovYTJJcir/cIfwE48a7Y5m2QsJBcKTI6/1Qhw9bAmV4v
fntr1AkSU1/SKu6jrks3qcFnVaEEckOcu8gmGApsLe5kxwOoXQ6lIgCAhmiza1gM9U3mmhwI48IO
QMWWW8PRMXQSx6JDWY0qvMxBTnpSBTGbN/B8/OdaoJ7iAIXFadotS65JrtDhBCsFQaUtY9ds9O0u
0S/ex70vunurrR8GPDYfIr4qObSzZb38DseBvx5SXFI/9DVLB4Y4yBAuwMEuiiYWKIou6IQ88ifT
Sba5rl76KV3lDFMEEjvRD95OGDUd7YCq87fpqRLAcEWN8ESPAhLO3re2kFjSZLyQ+EgmhpgtTVh1
JgY2MIDHqV4I2AZ4TDKzQe9yI/dC+ObMWjSNplQQC7pZy/HQjz0yjk4dMtL1Y3IzFyzr1qTWxbf6
atEIYR1Eq2E3ybA7gxmLYxuZBpqpFKPsW9oSiVYSBlCuGTk+YjYaecAnTMtrMRW57QsSxi/f5b3/
HWdv7RnqhlNpuhlAHwYfo28rKvH97CAVV2oSzglpm0zI1MBFs1kQdw1ilbMqP8qwQgW4H7CTkClV
a7hBvqWy7WxYn/66wh4bCPOpHSjBNwrIzOuIc4i/oykQzMccYcKSDDUxhl0FjluMlBnyVDbpyNph
jYMCnG7IuY2I0BkxS4UpojVOBIlSYnRM2fPJC3ecRazACzAU6Z/pMDy2irVk4MLsBhA250KRv1xS
X5IOaCGzcUQ0UC4coCIAdJ1FuttbtgSvq93Zda/mSSGYnug/MzwLfVo5dJP+6C3LxJ7pCaYk1Diw
ESTszTjj413tVzEUyHSq8gyUyXNavEEoqGo30D8pxxKVEru8B+jrPPGmoq4fdMNWDd5WRVmGJJmG
t0T46PUo0ldwSaw6fWcYzOG7uYkvjO2+2FXTHB4vp1shlhP5flYarbFG6PW9FUs9VvyoQvVv7tso
t28fBSMIOZkf5PZQCPzpecArgZk99j4yCj4pqf/abt/O9wCWNEhNYaE8WjZtr2eTDEKZ7ggeEMw5
Uiwd2zdmhxUUG9uH0O0sN/k3fvUanJOj5fCo+1W5xaDpSSBfMKrB7NUL0NpEzRGLwc4BUkX/Bryj
ewZ+Oma7VAUo9KX5ERwAdsVX7zGqr5Jv1HvDC3BctHKjMeKys5FJXxX4qYhPfM2dEsXIwp0wppz2
MNdJUKSH6LUVGyMhXGbw21GidsXnvjn+DxyC5tk57AWGtd6+AAfrpRsJhDRzwgAA3gVgWWdPUEyL
VZ7iKo0hE3EqQMoKWlR6JGhdaw6VDytyau6ZFRMkUvLXFVIA8jY+qPRJ6RSPgxAl5NTKlE1f652O
VLhdI+kPmIYmDOhaoj+SqzcfpRHU/fiZix2AhNd/d8NfdUZjQ4yZpmSiD18rqKSCkfNrMx4lZ4lQ
eiRGWVwoef59NQ7ytk8pvKVd5FEGfTh6oxpZYbo+KBJ6saeJPtNgq4tNMOwwpkIvSB6ODyHS3qF5
YAkaW3oMV1CE22o98FF/pqB0kWavWtx+LMZJUO7lhbpBZrZ31fsXaLSdelwpigSaU5hoJuO1BSSm
6dqeumJDd0tNM9nduOaUkgGVPqCT7sPq9K3/LDl4KYdVayNNu8iwsR3di5/j+4vyZ+b3jPszTk4b
0fLKr79eHlcvgXOdATwzMpA5eiHs2ibYPS35RQVkOqsV6so6xhARuJ9Zc7ORoDD/i6+kWy9QozA5
xuhMLSbzgeVTOxhj/XLtplz2zfqeUUtNf+7fWHivYFMSTOKxoJ/tdEwLoYzpu6sq3ZE85Crk/HnE
O+FmQUjXqz7ibBClECp2jZh5tMzk7lcDf+4jB82hYmDhO5MYopdfg/g9FEbIhjZYq4kpR4X53vMg
3jl1f9tN8Y9wF3tNIfmEdC90Fpj99BFuENdBJPC5dZ5tEn5zBxpz2samZPixPKidLp8DIzTNrCgi
yehFYENWkiB5jMad/mPngzxoFSvz0FrzLzDAU3DggIxPPsKOhM7m3EbnDuzZXhhtECde4lAz/ZAs
4Kc+1dnaA6SVAvwmBUMNnQD5O0IJEn0T3M2V2pTDo85bTbRiAgTaAJp/5ovoDu0e5XZLhY+SGmPr
ZhIySkfbZHM7PpkDyxlcdTYVItrpWab76vd0lMfqDkvfdqa8yL9oH84+2lxTNRxvGfKLcaHWZwG2
xycZFEdFSpGOoUD/Ancct8I8U2fYjX9Ywu92yOKqmorFaEenhnCXjUpJ2rLOT2n2G/Od4Vjui4j3
Uhm9aRs0CTU58yJ+I542zRA/w1Uj5tU8psoTltP5qPnY1t2OyO+S2km+WcXyFfx6aXVaP0OBqQQZ
z0BII48CMHXWnGYjCrOTHBV2W6Eb/tUfl96B48UiRbgb6aqxSM+fLGEjOiudTm2qbJUdrGgRZ0BQ
wtCULXqOmiiVycc3Dl3fJG7Qj69fHd7cDecgPUpcslsdLTrdkg+0eReBUBqdqw1GymBeBkrok8ol
P9wFmY5FhiapIxNgRabPOYPhNeZ9hQp+7FR4ghNwWxkYGHQghuVRbeecIqsyoHiiIrXg5+OeIPZ+
FgllTccdu85OLUQA0zWZIpuKckN2bK31kIW6laWFcVCfikVeDYY75+e38iSdWM7jk9uAixTF9r97
lH4dnNswQx8nRwFh227pQXKcIo5UvTjaKhN+29CKrheYKG6lad+HFmSkD8NeN6rIcjgevQP1k2O6
e05zfnLmrDzMxz8XORGZp143PUNbh3MvILIGmf4JQQlGtel/eGgWFOUygKEpOx13Jtiu1VkGDYjK
Eq6n50gSfg6h9SXz7Sy9cF5MG3+fgOCAbAON2RJ3bsXjqV2+BLvIJbKEMlbrGRHOu8EkrlsQEPm0
AmeeIXX8Qq1rXO29HC2ETsu0+XFEOwwx2K8Ds5NmZjcduaRnOFwyKAD4dMMsWDf/fRpUTaTcRU0C
BTf8yj0B9cyBvYpS8ZsaDyNXWaTde2rOdrYuYgwie7XO1CkwfBFNQ4xSH6z6naTcbx83/b56/Dxt
5Y9brcxi2AnWJgSxGMO4TuZa7IWXNNlkALVg9bFkQxf59jtFlM3AH7c37zEzBmalNc2QjXK3NefW
5mPaNr2YvlJwoMzo994kpqqfUZvA2wxYY9mL4sTJ+/CrP5lh2QtzvlURYAOChfd2iuBqq62WwdGP
mCf1PfagDhK1a1CGn3JFKQome55ZCuLmuErEXHTewN469upBAMIgh4tS0gAUztVvPru/Faov9Irt
Z7NXOBl5lQ2Q+2lZG8FCWZe9huLF3cxTB6He2jno+DKNy8aLzzMklYGRdT0Y5cZOk5VxewFsRJjm
2ypSIEUgXHU5R1c3scThBCMMiUBWQnqVFdvkykRg9WZeukRXrLXp922gYGP2O1PV6R7G2bE7Fa/D
jLqokc+DziqjFaNs7cUu9/NPi2ie3eycQjNolsePoH+MJ/rPBrPd3b4Z0F0rY8Kd+G+ksNkiNZBe
TrN6wp0HjLesha6xYTALGWJkicJGugqKRnEcyv3GzoYTscGpLJthDoW//WO7hLQ6/c9nnCG+AWbS
hNLfUBVt81SuU9MAVWgH5HBYUaG/7QV9t+7EhRqYb+4Le6Mf6JFbjgsTqgobuaMDUh5l/ki/Wlbs
BAUzP8TcdnTDPbacQiJek9Jr7TJ1ayyz0PFBDBRkMFlm/z92wBpwob09ArrT9ehQ+40owI2YVm5S
4g5IbBF5w5UwswaFGTiWRFlob/I2fANeb84ZcsxIj30m9d4cLMplFBg33MEBVC31RC6U8O+2qr9M
cJb4FROFVhp8BDzc9ytJ+kY7Gv6W70JzwSlzu90Q2f713GDSCdIpLiE94riAfXzn5EVkxfcUUitp
9+mYALvkMk5lzoBmdIYhFZpIKkuimz1IM1hPYs5PEGeCDgtyt93QHJuK2rW02VFzOdeQ3q4fzNXs
ZobIMOE/cEjuio9MBR7FeIICzLTR4mflug/RMvvhCoyXu+ciOtCDguNvYdZAVu4YMpnQdPcV29wr
de7Q0NvecePq3gjtGk45ROXpGiQGjGsXNT7NEvq8bbzVwsPIupLXCm5xRXh//q168HmP4D5p8nOv
HdwyW8HYypbUEEHEHVVkVQH3MsacR7awFWpCbCDlwRgF1PdxHvrMy4O10mku2odiup3cLCuTY0Qq
alAArjgEYEeNWYbCXRkcWHHz4nudcAmDg728hUlXZ9AyDG6IpytygI8ErQt7gvp1VowX/1NsQl2V
xZJ7rDYTWMR2fqiqUcDTdYBfCzsqy/WO9d8wj/PATAv3iBtraWd1eQiy2tpjue2RpueyfkZeEg6b
ySs0Crkh3S5CrYxJbGu8p2Ky1woim6Vgn1kl/czoER9ifCOZNkRaGSOU98SsXpQU0I3ICkNYtQyQ
B4PRrF5z8fY0ODX0Roce6yteY4+iGmsX3xYwvPpVnOpd2w3U56jwOm2adqYf7ed9/ljbsw6BoFBe
gI0cKQahUJmQxiwlX9x/QVdTBxJ1DLfE/X/PqFgZF6JmTSomD1YtLJVQRs7nQxYPdjkShV3vy/H3
BuEB0iTOBiH6Mo5PH6REUCwhQv75+OdnKDqSXl9GY5McDbJEvDisWqVymVlEfr+03FhYfVM9ZI8C
gvy9MB9Iov2uwstiZXyjj2rv5M5K+3+nCYMZUZbzuo/KRUqYUeBugntLOi3QX8sPkMMxgAi6zaeU
K8e1OznEadYh62LIiTmCZxsT9KcyHljsESsexWjNO7Kz5C2IAcUwqH8Q2O8WlCBnZ3cnwew1Pqpi
hRxdHCBjeVstExQs1m8Is6NzwCOFhdYoF37J8+iuKUNhgsDlBrHqij/Q4TRomLlZ12zDM+rvEWbe
bCCHsd8AjfziVVi8RnYFYG1gsiChnqvPipxTozzcz1MQHDprA8cVtWCt9U9tuk99Dcp0CWi4ilsg
8Wye4FRuHJkfC8IojX4VVRSFDBsbL+lxaF29NCwa8ViaJjiMAUczyvuhmCO8SwnDiszYSd5ZEH+e
YsoJdFvqfiQkVJ6SyesHuHNJ5pvffF48K4ZEqYtCvx/lHbIgvXU0+2Q1nA1x56hl3bOrDqtmYlnE
8mOqK7Ml71K+HoLt7KkrxE90rjW7NBSjG8LuAPCeApsQ8W++L0B5mzGGuMEOve5f2Ey6pZDMx6At
z2t9fTIsn46BmQNU8OFeA+qwOwZ1bgAmlj1zSbmC8QMGzIfuf6Am7cXhIJ9uZqGtDg0KZeR8Zkdq
Pg4ZgOdVtPe7g6DYTncQaVlGXWfVU7vBgcApMHq311nbI5Zt8BZXL4mEID6tcorX0OpE3hQKxmrg
txrYqqqdH3rClltvIs3gcltURs2VjiwfHwePpewPJBCckY8+YlAOh6fVsukur6WfuPUs2CNQzrMq
5VYLNmT9oWvCoGDNrAIxCgdliCeIq+yZZrImtJtPOw73tLjBvs5KZZ5OjLWraoVIoKsejJSfrXIO
XejqiigQPEG026PCmbHOFWPhxHyUrAbokqnltd7WyLKtRWfrtNxTUi69Vt7AA+3oR3zd/SEUijO8
Di0uAlwlYqGoOabp3/3ReKV5lb7Fdtpl1M1cwZZLrlALnMYEuCPxCe4JDyG2cSXZtF3X3eJTUY2Z
eCNEKquuSBBhUED+258WHSvCm6qst86Kdhu030i3WJ9y8h8JzbYuc2dGTYvpwxkMZO28gy9CLJtJ
bjcL8QGjAUp6fs8879II7a926fVW+l4tM3OWDOVznUug59Rgld0U/6aXWveN60v6E9W26WZ5Wry9
I7LZ7bcTH5SlPsylZ1DGg7M4gBJcW5kE0axl8+i7sV+aHO0LgJvCMKlfn9vs+5MNygL8fRCvh984
BrteVUIJEHYpO9t7e5QqYyAGSI2h/D6BhLnv5SDgRIOKZCwx1ZrTxD4YtFMkc1E61nqsc0ZGDPHO
JUdbXgHVqLMDpvKmJBcXkkStngLG5u2ggi/QZnBRpsNErR5yW0FsgPmXFZzuiuvlUVGhehX+H5+L
W0RqrIQbwikeTPiWtMoKjcXDp0jKxvCMDFCNfBHfvGbuxn2kwhyHDqmURrmPPeF4on9zYqGTc8pU
nTlZnKKqSM+9BePMCHBGldcA0dYw9u/zPYKfDQ/L98YGnBA6BsufunBq+GHA5C0gmnMx3WflvClU
XxKZZvHzoIOxMyzZnsrQJbgB60SHJ+tUWB8rIsFjIHnN0eYEkj9aYy48HsR2FPBHrwRqqSCMF1pG
jk6OXlKfjT/gBioMZ5XlF7jCC2YMsoK5d5z3ROExhxbMGZ+zdz2Hw7vExPpuO05WBloFXJEX6MDz
W9+QjVRpLNO+5Efsh0YpKof+DO1ttHbd4mEBsIQ57YF8qE2jFwvhMnHCVKPSHJeM8k1vfedF+Oqm
70dNmPjjhKlITXMyIvi1PwnifclN7SgKuE6pIAteETLEtRjhGh+ALQiln3nPCvYIUfAvslML1hoT
5+3Jwoukd5+ui0pOqnyOS79p/Mn6pfa+6UiLLRSCQVEDIS3OgK1mShFOTnRcWbz4MwWt4q7Cfl+q
Y0yWDUl3+F+ECgqEI35X4p3djkiOhWteVbw28LFvfPyMy8kjCKzap7AevsfQJCbtmDuNyB5ZKNIz
xek++1qATdsuQZ1veVJierwGiclQh5bzp1WJKU5fWtIj9AYLcFO3ReHdfpr1GTNUk0xJ9ddedhJp
k7Qg7aROIUkb4AAIfxyGyrSbT8vvQGHMpQHAYi8n0Dx7+n7yRsFnnrwDUz2el0cQCuMZJDFz1MRF
FadhWiyXv4DKNnsdZO/zaHTe6QdTxJpPM7TQ0A60h6+fVtbpajhnmjqP2WnNeD5MFkualjqez9cN
K9YBw8W1CH5TnEMAqp/w4OWIvB68o4WQpDweHqTNSAg57pSFvW15m1FXidXDaf6YhstywLIQUQvc
MusZbJ6sHXySf49X+7Pze5kyQFKtVXkV3Be1Zx8cfVetcRAWqA4Lx0BKy5Z8CNumwW5PVMMwUqmW
m6i/3/1bjfcof1zZ2/MfqgnlfHnYzFXO1EMo9W6L03qVI7hV5adcefCWs/75EOO1tRfo0j4RGEAO
vxiqOoEFWN5pa/+7eQ5XqDkg/vcX0TbiEhKC+48urcnYIVxIegSO5Kc2QOkAlfQdzgxC6TSqHHyb
JdMmTx8GE095jE8FpWEwvoEouK9PKVUwdx8j0OWKyj7PfRm0WcLNgrvQq55ZETz/+ZrHwcFb1Hk7
0hiePPifmjC2pFQHPGmbVcUh6xyKNpxXy67kQaTGSCu3ZDhaPFlFRfgsTjSPWrtX1IM3f+ksuZSe
33pLb5fvdkX8ibjVFRQNaNkAl7kfoiYnikRE/421x2osQFR4muSLxVh00SWKilj6EKNn6R+zrgiv
NC/oitxMWCwe5AvEkHi3goZWRLingPJpgKhwDkg/aQ6a66LYr9AWeBqy3edjObvk9e8n8iD1eA/g
DkOZgFNKVbpXdQ1zFipIDQdjYID+yAibsDa25jREutpGqVAH5FvVEbkOQZNEuiPFX4epMc24Wduk
OtIjdgpGyB2W9/oaWpAbVRbCbQFO0pQMnC6BQ/NGTqanAByi7mNRnHum0yiwSauBrdInWVY/d44I
jAdRUEhh34PkNrF5nf/pbqt1mpZfLMls0p551hc9OynOpSY4XXoFZv9y5q0dti5WLMX1LbyswgBp
0EWvjI3KmZI5+Z+42DOrBK5htYkvHR97UrDXyo4qKqwB7AjxJ5IA8ui1hmuHzOM8fIFkHWDJLaom
gWvAMggBh24WgcsrgHVWzQ3jABNxaZVA5tql5MzJ73Ik4Qfm1we8rOxsjsqZPv889jjumTTwzMBr
6yBZa5BhOk1in7Cok8abocGETCjfNyw2Vi27PhXVdXWBK6xWP8Xm1Y38FAHmXeTXhmb2OZjBDNxE
Hs+38Nv3t0Z/B9OqzQ+4aqx1Z/rlZkeHFBS1SCKJHUvpTzCn43rPXOxuEnV2FA5PW0lWlKkoXnWO
NpGd58n0DSVITPWJx+E/BZSs0B+OhOh04hzBO5rd2hGLBWMtm60SU4SWq0l7BfOyYFSngQ+DAzgm
cOk1sJUJXTVtUr9YC8TJME2nFemCNLUmQxlhofg0cy5S5gvbLSycpUhAnYMuIncCni7PK57ZKjoZ
9cTIWYmMeoW+dQwSQDrcpA3bUQKRrQjKq70beC/0ZrGDOSf3MtisSaqtJ+TY9Vq6xcz3VUeAgcjP
3FSyqyn62bvk6KYFg8KPYF7gOeljl8Vv8nS5FpHfzLCoekdab0TNZePa2RX9CCk5+D/kBh82cmX9
gpK9ilAs0NxJfhyi0n0tRrIf3zwb1BWG18xcCzWHtrXkdmJkPwhJ5Tpei4lYVA62v59Zuox9lyjy
GcimBHYoBwFCoRL4d8rGKtYcCBG2PS9eH8+2aSuOmb+JSyZ8jxeT5zTBu4CpuolEoVAHTxnVWInh
BQbnv49RqsLVq9AChiZinipBYKwDsvMU+a9EGaRTDZ4QSfXvqrvUV1ybZAyUB3yoAfSYar2+gtdc
H/68RsshLsyEJNZaCkmkMehcZZyezUomK1owla8mnqRW4E6D5w78XhA/48iruAXY3v5Ub9/Hpwgg
0RcT7jF4TInBMF1pU4GbWTjCYu/VlvknYFuiZs2ii796RVo3PagTwoJ3znHpmHLSjsveBTc00Zzm
M1xgo/tBpUxAcEDsZKEFgglxK1hL11fcUC14nUnD0gkVFibvNhP/3ty5nSY+wAhbT4YC5JLM0N4c
3ZQx61aNe80EftvFuZzYIzNXdVATmhOEIsVVDUoIMZuDyMS1iDxtuPCEih7JbtK3idQk01eBlrtr
4bVRRdpJGWrzQ0s7z7zs5XxhYqM8tw+m8PhK8bL9kG0etJaoTJYr63/E+rminhxlNgK1fesleu+7
oYyW4ivVVdEcLIA9TwyxcgO9i4rOKwBtjE/xiBkAoaMcYam5N3mtRKW3UQm6nxr6CVDx3TiYaIIA
HlWaxSAYRCxVPKBysUTlBifDT7vs9+MD6wTMSiXbKC2HQA/metIDDf323edG8M8eH1F6Ld9LAFN+
2nvjr2lzHy529aiuK7TvPEAxQZi0wBOu3F3HEKOkaoU+IydDv+iiKT6kKN9mTVTe3JPQb8TBs66m
f5TYxxTRmvbEg0ihoZcxugfSIDYkxWJ7PuH2ykOzzT+JVXNqP8FAEx6oCqutIM595epHEH6vWdGB
VuCxI/GD6CsBY5Jg4uYhnjRse3jakP01XiyHnucGHr+EMzYw5YUpQaS73lVAhSv04C/33EWS2F0b
S66nEZkAmGAItZl0xORStQ9t2yDHYFWgUYif3sBXAZy11Y00Z4qNPM0uz5X82UdLrMHLORAxGOQ8
OfE6MZUzd/9BWZInIAkuALOnqBAEldOBd4GbFLIFDWTgLBableHhfcZMWscnWNMMpI9XS54iFe5W
e9wfHmOW/eN7R4J3xquVVECEDB3R5+Pw+nmVL4d/3QIZAfjuw374y4qPj1gKA9YDfDWDpxGBgUWi
yg819gW3GK2Jlgn9QCEHgSSii9+LDYXchq+2f+hDkhF+pY63OHZok3twkomQhxAZU6q6I64iaSFV
xs8yAmRNbi0zEEsTDPtxSjOdwhfEyRMTSg75jxbQW/PDuODjhXpsIlAdSk+rYZBCS2vGSdr4BQGQ
BOv2Xx4xC6VK/lDlxlwDYMQjrGPnlq1xnaxSEvRUtKO8dmFTMyYEk4vfaQxcu85U/FNwTHWZtJlG
c5ZbN3U3QbXhz/2di+ka2bPs0YLN/ML6a24c0s/nYc2aIi8VQIiaEOodHK3taMCMuW+UCcIzRNig
6Mpu23dJ9Okmul6qllitvPCaArheVJsIakbod2hvjT8U8NCn30YGpd8m4gCaW+7vllExlqVXM9lm
1/aW+EOfABJ19gJSd8TQ5ld8SaiJT5nEne5CLn5uxi+5ycMNm9yP7JNZ4mVHVvStF68tI0wtniYh
IKAwbSkWdkZ/KzN8995wp3mWhK/Lam2vfj8H/XpSy4dmzkJOsCXD1WDsB9yLB7VRtT5DdggFp/pr
pcrqS31E/N7QY0WVGnH0ym83q8y1UXmk/vVsWJbhvsj0BQIpGyPNxwXwg1pAqBfmC4/YzAcwr7Xf
LCySDdGtvS7rKLNFomQyAxijHq+XEzGLziYSralsf4iMdUbejg22fh/qf1Owqo5S7um0giJ+daFV
7J/0I6Qcc/XUssMz3qeGKepzetg1SvbuOJteV1svpT29cmIudaPTBEDrqJbHRWlMes1exidMQUWa
yino40uGFzfmUB88j36YBQJWEzCybhqvXB86myTQJ0zQgMxLpsPZFTz5RGQvIsgacxk8cJ66CMMt
O/3AXv6fCeEyHj9RiXmhv7z3F22RBTlUuP8KJBoMAnSW211Jzvcl6S876dawN7b5vxK9S5nHj+GG
ILgMj02cN9F9fLApqW23RD4Ou9D5wgW7YMPoMJG/sRTyLJ+PFGpU5V8/kXNfa+lkByZYs6zio4jx
Dg4R6WsdlWs6ZQvjlLSqdm5sgh3mji4DxV5z5LW2Qj3NXLjbah8rDicQ1kVCWF9uLhH/eHYlhsP5
06QrCXvr6U1DpULXYRJa8LLuVpA6uJ8VxudkwDL8s4lLy1LvjztadbGvye3nZ02AWmiRVdmz6YSw
IGwWdHXHNmyVepHIkmySFoLkxIeuSbwfqrx8gbm9HlfvWaHDHxlQMVsOJcOcEaxjZjfg9UoBnyci
UFGIRXxBHDmqLn/OQfCigJP61eQtgdLkoZD53iyKOkj/S0avL3j+ivK2hhWROVDC1ylczKuSnDtU
9dh0j8jkuzjx3kKLtS8FLE6S5RidY+dcKRyUqRXzIh55YtxmmBjWnVFfegczHgw500K2EYQvYOAu
/4QJVD+K+u7TlGC41qZUZh4sM//Tx8HdpEJ4HGBg2BVgoieLSjqcic8caunAqUAtA9Os3by9F3eF
SMcCyhRAVcJ+I4BHyU9I2YXXKF408sz+0VlLrPV/PhTQHQLFBjnx+PRcKh58ITUi3BtGA1ESHAGA
gAOe17V8vcvxwpFymsMquAi4XKFaZOtw5JpW1SIGo77de6c0n/ElHHlOAHLkZYCtWJ17L0AV1ytc
lWyTFDHSo2RS/PLnPeLTPXTJi+X8ilUDn0GRsULzTn9o+fNw4LGhVRSTastTvmhJb/BwWjn7pIVs
sYa3daqQbU8aHNoF3RRGXF+170NDoKdWxTzSSOc/HyQapOlQEh2fTJxaunNoipqosg9i0L88R6Rg
lrQ3jpN6aS32pB5kfhttxkc1iRZ0TxE62Hzgq/ghS1S5P17GhPzUD4qoAvZAViK0fAVBRRDJOuea
2sAk+eT+5KD1X2jsHpDnW2C1gplxskQR4aT3DrOwVagGy1AMhvWTi6xan6ObfNcF9sRgwuULpsQ5
70xxcFOHe5Rdb7cTEayfMQV3xNlzkXVnnXpPoSSbhvmdwRy2rJ5Bn8dsqjFym1HMBCzX2crfBhKj
Vb5sfLXJCRRd0HsZ1aWKHqGJ0pz+ZBWNTBtrrpH265j2DvUlnhrs3NbmbMPNESKseZBw6aHATW0t
zlhunv4zZ8T9N4DvKEl66sq7Pw2PmUhrozBXjyjeslFIMxIBqWFN0x6ED6hEfjkKfqQ0bZJ1CR+C
IGUVBThtjp8I0KkG2bZ5R9wG5UcTLFK8hKVS4wt7dBfx/H+U8TusZtZdgzRW7uj/GvQ2jI48LGBU
gbVBB+jyg5rBpFiY5LFv6Mos1O28va3TLxS4yzAt76eRVPWsllvI//GfxGSzmniqjwAi+TOweXZg
jPL8ma2H3kKDIXAqYltcpEIKf55Yk/sJpVS0rfOpTuvcvIrzaQwev8QQQrwxVGKA6hbn6CTIMZ5r
7UvcbKi9kJ9x0SxDsauLUWmLLm3Llo4RzDedqddGJTzTlVoB7FHtrwuxYYkrfTtudiv8oiwMZ0uF
PbrJj33m8M3Dy2z2IW1VnNLBn3oUkD/38JlpWdxXlfjtZ4X6MZK+8luo8g0oPsh491x8Y+njUGml
IBtymkZVYXYxr0Ca+L7GOAjfI81B4rdvG9gJwogKRySa5KfGkwvlm/1xjD0WXTgk2Kq8GhUMqlvx
3gGNUt/qDaorud+dQWMp3R55UkZXGqYw2hLMtGw740giolKzafK73d/WT1X+LvilMCBYFmm+q9D+
FRUPkMfSL5/d17zV8klV0keO4ngMac0eR4oHKAu6zUpbxyRmMq4j2RcYTTM9cowkxADHaHPVtQKr
DBzfeP1u/zYCL1+gnT80TBiFHtzzDY26ehnUK2AMF6neKda2VlYQu3G+UnrkQcIGeXN5Qiu2/wHy
UtjcXbc2M4S860pXapKddEx4XIftSYAVmoLnRcPVaU1Av5hXjF1Q6sZulnwK+eSUurs9pUIndUm8
JMan4fm64f7ioqH37CGPMZjUtmkKB9J9sQn3FPANdoyv5x2kalN6SXS78yr8xEXd7maKbdRGMs6T
nhXvxPMN5lZTkAOfhyTu64nXOSbxtJh+nawsp9T3PfcZ7Lur0i7hZEFHCG/J/6rPZHWGChtacboc
RZGdb5qiqN4kaykWyxfoHS39myFuadT65WTU965v1YC3P/h9yFykFlxwChkzWsv3dqRPri3ujHpi
FZnBZGIWFLNVh6xfQML3cFl97MN8wblUPGNhJ4KdHheUcG1osj18hGf2qcz6fZj7HpbwJqyNBuiP
OdX0M6DHgZUlP15cC3JjNlON4+ZudYk9N7Fsxhn1kdOr7d9UPEa7UtZ6N0mPO0rxAzkm3Uq8IIs+
c6+Qgz4XlUvXS9t5ZtShVgFLae31B59RKhG6e2WksBWP8HRkeHqC1I34LCY8tRb7sZs3ltS4YGQy
9Fx4LZwly6QpmotaGSHD6LwljBSEKVkn88N/689khrF/F+cxnViStiVh+xLrrDx46e2yYz8Vz/ER
hN6oZVPDYHRAFMnlMRvIHhxYZs6z/XNaQRAEiWvudUATEnkt5phu11KJojFFC7qn5kMp63lYDMEa
CBr/HK2zSx6RVKMGMJcRwDQiT+dnfDRj6hDHTmz10u494JljiRjC3axk2lT5lZ08JYN7j7XS8/D2
3jZskKB17PMlwCHQrdAPDT9HOCFGbnImBDqT/osioSyk55eu/tCVV3cdq5Hg1pscONEg3u9gjHs9
/9FaPGOaue7AFh3oUWyr6KfpJJeUkZtkrpIaoy2MqaxSso/GJUvZ8E0TPpROMu3rIZ6Lm8+bbCkv
bt+9NH6fHxhBjAsH4U1+nCxr2f82hr24p8nXufJncxD1rrQrd9uwEYlR+Q2Vn+LbOMTCLxG0/8uu
PBQ7umxYkrJZs+OUM8fSyA0hl/vJpcxsxmFk+oQu4fPgPiy65XkJrFoJlp3rza0Hsy8eQHyqzEXc
n0/zmhm9QRopBNVfd09ni+rizNPwUuSPvnDlNCeJ1eOooPiLnqFEOx3BCEJV0QLkBGxZ2S1VLTtJ
eCVRKmwMZhHu7p8nCkCDA8qF374bbBvMlfoioWzJkmWzxRA0Xh7HIrOZeccEJEw6gvpi34J7nk7m
e+kNmkboIoCMlr14YFosAuUsdKOFc0uPn1NZKPGKS7KWWgpzWvH8hOm2Jr8dREHy7RJFDggK3mix
liIQAMHw80zQTDFrxH8f3oCna5u0gFWzZsGQUOfd6/zGiaMkcLogS9ia+He9pnVla2R3TLPcss23
mwk6HW+ntq5Bq2CyY3yuBTvoK4kOGvKJCZJjKs2QjInX//U8ZrvtyOpINqzHtHc9hYVP+InmqPZR
AYNZTo358mzP8sm6c+EYHPG4tqwdD3vKElQiy6HzoyDxGtkj2FExFjyc8uebTTtbzB0fCFp+9W6h
z1qefbUVMW0Ajuq9qHgqzJ6HYQ+/9nMFCe2nkRHDcQqpNY09UjTAS/Ce/Y16YpoNm92nzYIDws9N
krav+I55/YYxdeAn6sK8BYCWmc9YPlWgFxlLrZAsD8Ml8tR02RM5EB6u8i/2tbxN5RaffWoHyKZ+
vHcLPFxBUiGGbWHrxoLzV05pZxEGMyi5Jb6H7n7ZlqJA6IP3mAr0JJTa0bMd/ViT6d0PiHG7OvXd
69CuhKTwMlkmix6Q8wB2MJHaD+c1THhLvSuNqRUg+eg6pHgTOMmqbXpQSsr6vXD9IeUX9HOo3ieY
AnBVMQV9Yh9JrZ0GLHYhnGFi8eiiW8a3dNKUXJIKyWLmWEgeNjmItYThrMZFGix1qyHhc03HwMkX
Fzfy177PE/rFBqdzxGNey5cTxXXA8M8SyJPw0VWJvGa1hqsvf8uUa0QB1r4pKsmHSl9Sk/qwFALM
0HuJEsxXRfQPGsyZgmguUyhBX7M2918mPOZDyWDhcOsSvF/+ih/rDoWnW18941nejs1FN3Ov3chX
kXJ/1lJnzbHiqYDAit6aItWo1UdPvR0cSBVEa7ILxisz3M+VTVU3k+ua2KLJuOJkV8ZLq124+GnT
uA80YuKM7pqS9Qghe0hralS81cEksiC62NmCYmeLxdX0O28OpTGgiZqqLSIFMj6D0edxLse2oRiK
MyALEZlDHGTeGZU/MfQO+7YkkFyCMr2qUsOCySngjy8xB4T3Ow8lB/RQQcamgyqG8+DUmEk9p6yo
NIfhkpbkA5SXPwMGQQFeqYBODHNOpvEWAbMcgBnse3Vo0BZXrqIFlSBxiznFsZmS9YSDb9kyI0B6
HSr50EOjib8RQmwUOiMUK5boDcTDSh9dVxCBOc8eGg586q2TV9f5Qf0iFRAjk0KqPTTNZ09s0XsU
oNCob++bR84WN4C5tqhO6BQkrF8UbspvknPpuXNFc3yY6qUhniBStbQBN7ZiFD6Hqd8tkcKg5s8F
d6KOTPeBfCQpHas1s8z9sSxQy7XqvXiUgOZr3JWUGWO+zIQMWLCWqQVtAXy92PVlZX3q9kBahBwD
SwR3CHR7A2R+5xftx/hVMs9/5zXxfcl9f2ft7EU6MTUIvyXaE0GBrrVR8YvyWqrCu3TzDyxe50tA
zxlyjqKHrkVKiu0L9+jP9SYSAenUS1zOekn1CsH9pRv63u8bhHE9MbTBl0P5UPdZIeHmm38kcsU7
j2wFGkJLbj/Vo61zKcAKShEw77zEGLTZ1gHldRYfm7YZFZQPfJSr/P4OT7awyrPV6i4od2yaP4TY
qKRG7NKV0cU8txRVg+uK9MFyBZgtkajfEWIGCKyX8yAHf1keFsHGIogwyMQpWdDrpLADkEq+pLD5
/6u2XzI7GIAkd3toDWzOq3Kopi7l7qcnChw9cNXeDoIrE8hub9k2i9/3poPfRzXKyyt8p3Y1xutO
2AGApUy9Apz4hoLR/zOUXe8/5f00TnJ6YcW33XDHkJmrmvTC+clFEvfj0M+PFRWiL8TJs2UERSLN
mOuh4xkqKy4lLSo/szFCj7TtQaswbi5jo9SRgsMTa0KOHd6LCZh5YOEwRclmH+MBqhThqke0jZ3w
EUB7AhNiLnnwBqVsxz4baahjQZUeRQljaG9YQt8/J8EjjJTE1ODWvg0/QlP3OLnWCAeDUROj3nQ2
LcvQty2+BabrqnODxKIYjcIV5aMm6PYih6eeuwkga8gARGvBmMZIYRmQZDgYOeI6lWVwKS+bFjD1
TQuicqTK6Brw2l9WME+uN6/IfEWFVy7zx/lQfpmtezxM2oKPvfJ+paH6xJaCjhh0z/Fi2OBjJK9m
lnTIYw/PUemHmx9/PEEdu7PzzePiD2C0RDL/dw7aIUDfrKBfRf+a0LrNGEodTNB8dql8hOUBQ+KS
pSaIuAAiVj74twwAL4BW809zs35LSRbxb3hvGV5nawt1KG1pTnhyxXZOAUXrP7akVvlU1W1aSLIN
crnX4ydaLdRIx4X04k7eeZ5XKMaf2jDQQt3T/SXAFKLpqyQ+ubpTOtQ+shaFAkuSBrx3UHpesu/9
Ia5dtLdvRsiufoUyx3po/gpoor8UiGe2h4S/XDLSv16bMiYopADYWrYxxSTZl+IMWUmYiKIt/APX
YjnGUv1bDZHj9FsmSz9H2M6ZM0w4R/6Qs2a3hrb3BQSvoTWlBdLJ4nrw4HdLMeGo+28ftQtAE1YK
0dUayoxGTatf2sDyHhyvj6cYsCXEurE2cGa8lIyRc7Yq1xz3c9TGmyond/If5nH30gTCiGzioA7K
j8IjcN67vPvyZZ/AO8cn4g8Q2nHW9MXb4FGwjB0Gczqw9CJBJvZkuhpIBNwlgZLUYJZmnENlFRGb
i3t471cG+2cYwm9nzUsG+BRZH2BpZ7v09v0anx1VyqvSNY5TecDV+08DNx3KJaA3PQ5Lt5q3hond
gl3E5MGrINmGajKjBqe5qz0N0Ul6JKGh6+1i3WUhtxD3TNnGY/JPrPdfEOcDTCBZHm7+PDkMMC8b
z4XMoLK9oo8rvZY4AY1nGxMymQRxI+MI52M8zjCRrsrUNUJzhv5gQL0Esl4Agyvg60D55MVyneyn
wfiPrNxHRWva68hiz5ZzQ9KpTL2IyBqA80mlv1t9IL69oS+HTzk1058ywEChz0TxCnTLsIsj7L/G
+RmLE3ckenV6RyYP3/MLHHHPT8uUlWc4t20gLyph0evSkzcC0OjEgebHqWbg2qDwfr77EcxA7UX2
KRhMZAP0nmXlkO9sG96pKCdyj+SEakEszmAVROBXgMQZOUSszI/ky6B0HNwkk2J8J3FxtvyceZAc
w853Mc5VlumZyx0DyQuipkOiYD6ZJhJqEr4RhPO3ufxaB1QeNO58RVfFkSoQXNQMvB+cPpbnNTaW
8sqwmeuvUqM1kRoTlsvRs4aP+7GUoglOLrQw1TrVYGzHJ58lscv0YCyLEQl1mmn7sxAhVLhL12ce
lmrtW2mEd5/DazybSFBORLyAAklub4cpf4ccrM7PTp2X5pJbC1sROa8y4aC9zBqiLufS+UX5MlrR
+tphvsC/v8PqhIpNPfP+hsBYEnPmn1eU6fjPSbxvNU8yNUhXK/Dx7LurWzrrn/wnd2pszGbcgBwW
FyJ1+49F648LkhGq3lnSfEMuEHqiSaFTtLC8RiKu3QMFzdk+cKP/oZISDYvz/eMKnvH+7jsL8WqU
Ji77UsP8zU1nEmFHA7AZ0g08kLf8la8DgfiZepbSuaEdw0gEpvOnwoU8mAtl+KvhR5GRUuvq5Gr0
L1mxQEN/N0qMOfTawGhLu4IIPZUB7OTYoldjC0y24/iJPD77jE2G+Cvr/3Mwb8+n5uZCdmcrTfPA
t5aHG3LueMOEwMYix2aRsBFNbW/ykIQsXduVtmokiOa/owaBmagBY2E6jOgdOUWD7keBMbCSzFx0
JecH8ZlLEipWhBmhS0kP29IR+S8q+Kx34kvAg/s/DL8jaMlaSx2gnOClHTu/daBl3v3EF1lJzUc8
krkRT8tgq8BCMHVuGswT0Z3c8E5gvoBHMLSV6t52wKPJzQ2fI6ZAm1CPOuGdErg7P9nbMDBmmcwd
UcYaQ2HmpsUGRwGdby4F5PAYJn5PQvhVFcOsHPVJbl7IospkzZBECmVQ8RJPtWmc+Y6if4YSocTp
VbcpLri99OrcZ2DH/3nBfQWb7XDrtK6zJiClBA5hLJJ2g/0kMZ5s8unwDlidSyTPLgNoWdKiQwmB
Vp511mqPXOqvzDJAIQCQALDePjuAx/ZiavdExX+aU5rQqKV71DiAp6mHPYE7s17hr3acCFeobz0e
GmIkz6RxbLXmCWLaYfYhvTYk/B9LqbMVwdcGxMPJfuN7AVJkmBCfbJBfIEg1kdVxzVHY1jS+SS53
ic8iP01B1vVu4tgQwqXvQlkUqYZMxmIniB7QtYSBJkb+H3Nv5r2Pb43BFObWKcRUoReinY3qMW+i
n2usOY/ZPTXaRPWBaPAz48Jmzrd0ffb5+NCz4+ekVNevNFdqPoUgKHBUsxRd8wZf4LN8B0AaTKeU
XfG9X0M3xQ3b+FSrZJrR0Z5ebTIxfEQgIWlIO8SZhBOKVBu31889sRxV1LOnRAQbc8tJzcQEPyRp
UEMOInOnd6x3erpG7gze62wpS29niP5SoVZJUFBtox4uqh/8N1vhbD7pZQGfRnLlciFVwmE4ZJBS
qKgXDNqaogJpnZrfN8JbyxHeQHMe22zbPk+qQNk4Gn+5prinfEmkNB91MQo2l4dRM3p7UrpTjvet
JL6o7LWTRXsK/bq+7Yx44XDAKXIjHG22b2rGm7bNqtDrI1sJt0fqHwVyxeTExr5PGyLP4DzY2CNa
yuQW7Lh/KZd8Jq56UE0yF0APbTdATz0kx0rQ/uUKqMs1F/e35kWlnVL8gZP01VAMVf+hCOzO09cI
ewSTLfIM4kkufXmvr6BdnVgVf3Y332dtpltxvzFrdNzPNtFzDtWfxssmf5/7t4vVqYZw/BmCWOfQ
kussevhcROCrAiZjuhlnPWjWi9a7KIVNXetTk89ODHzRS9rpuPdYT6uFbJWJQxWrBDh3PTSln5hb
1Ca5/hJPD8fOeEi1jOYRA/4ZQfrDmVIC2hd+tk94uM4XU6iKpjzvdrwPib5YINiPMl+YSbC5Y/4b
V8FlAo3Hi9bRh83672agK+F7lZLMIZwwIwcOSZ6wxC/oxth4f/j4ORM6ifFkNCpADt4XmrhvthL/
Az3yWMq1mH14cEfmSWsB9dMJ4fQOSUwILKNI9zmeahtd1Nug6B3b3ylP2gL1GkUcLq850IVXB4V2
3tFcxpAdcXMX3RRKgZgmzBhkxiGMWMnOo+talvlWjtHf+uQ+OLL19oE2jRwXK/egLO3YblW1rZAS
dnn2Aa4szQFXaSm69jIM9CWLOZJ5avt7xWTs/Ygy9pLa+m4FbQvq3lB5dyqJFKweyOagoRFS3D9b
BUbRkdGwUEjABaur+CvU9/bkCBKZy3K3E6SiROPfN1OrC6UDqnrE/i9EJb8lFQT2Uk20B/jUpt+E
Mo1cStdiFsjlDTQhBpq2zV30szxojAf3S/aVcun6jWUOozfTLZ3w5E3z5KOlu3wrHIvc0JRe7/lt
XcB2TZNXGMyNRRH2t/ofu5LSG0OhqXfoiTwciRSW1kQqWvjaDKVoQHeijFe5Y5r15kzdADRRVCTv
yow/l66FW5TN16N+s8xWA6ZKlFwuUERwkGbQBm/x0oMfkBenM91MH8m3k9XK88zdtld2DfbBzCDv
RcXsl0ZJqEewZ40zTrClt5Vb4B+mGX7sGXVc/3X20vbR1zmqADWiibKAH/+y//mcumti+x9bpPWM
eltSwGcazDLTCBybX2NGiHkX83Q19Yq9HM7KLEa0Sa9PYFcDN/IcyAi03PxyImXbgVUcb9dnsxt1
mfrb825A065nvFA0dbjU1gDxsfC1DYUGS9AKmIITNUtdhkcOZs6CX5NOus64kvxryWT+g+1yERHY
xjmtFsLr6Rb+4DgDC9xS++KmbIFj2FaDJSYMUxk6EoZ4fYvl7ed9UfpeJBe/THMmxh2epVczQxfH
jiNp8Ei5SouBck86O4vlCstsfG1x9CctOL4MmAsfsLjymQ==
`protect end_protected

