

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
E82wkdGPZb/+6GZoDi5HpckkoDtuL8TGRb/JCIEDYKunG0ehlHY7rWSAl7AxBVkDytYXn4VY0NY3
tD816aZ/Tg==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
aN+8nTYiRF19Ga2xgugxmmkjykOIKDSAJe8CuGlE1RsIGMA/TeZJn/LIOmkC0L4RXBBy5zkZr6mC
39gWvg+KhH324/pLiKCLqvJkIObctxdk1QghQFlwGyR5AgwumO5V8XR0wkFrGx5lcmF5I1Ic7QCL
4FCmeVtU3m0TggWFC7E=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
aDXP5DZMSmAZ37R6bG0c2an3UXXBQ9f2UcCbZO9jybJiEbg3jaEsz9OP8BILMEuM2Gg6zqGospJo
IL0GjwnUkhmqiXNrUyuU2ZA9j5Qfpqi0cT39WDwUPJ8gireHKMW3Lk2XSOOhzAT2gL6kjlBz97a9
e5WZk5XJ4JpzHsyykVOoT9yBzVvTvBYrbMxRFsaT4GZ3NCp2/bL7FcAdHRGbG5cNEc+P//C3rwO8
4GNkm0wKVMVQq/2HclGOKJAykNBN7fGuG7zIF27nKqnI3IBVFzw28uEsxwVFMpLMQ1Amv9lQcw/X
S+F0+1sbjSvaH4de4WOv3cOUzYKQ/wzN6fSahQ==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
c+SPO+b2cpVqItr9nAdAKH8LRjqZZjyv88QHjXDKD8kCd5SL0IXE6XqQ/EIjme3B6XJax0d6vBvr
92G/L1QzXOo8P82zgbpcUFM1hqtYFVROwwLTcIHV5QmMcqgWTv/CxjwYFY9l1w/ADUzzHakm7vO5
G+sQHpPE4aud4403sjY=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
T8GeY0or01NdwqMo6UKJMUTsmtP7APuN0oCIY7KzFu+PsK+FyNTk9rSPzJS4j6dAZuNV0qTymCiX
Xbb3asOZtqkbmx9Ts0TBudlU37PFSlhj9aboLv0+uBJsltC8lWgypATvI3dldUNiHT8HwKeBDDaM
ge1f8g9YSSRm9Jao06pgbL/b6i2WQcOEh+n+/rJDy+mhlYh4b7sJni6U+KkkIH+Nz+FTmo2KpEia
kiQmZaPY0KLlWtwgAmS9D9WXDnBy7lDRle2NygR7a23rjPwxBp5MqpWylPuquQQaCFWvB6BJrqSH
TxLzvd+PYmz3XQMRs1MJrzzaNEb2P8EXhMkKPA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 12384)
`protect data_block
NuQjmFayU23HaOtjx9hLvxJ4STaQk8kR4ugKXYBETj6Jhe8hOIuJftVUVik8lYAC+TpjyEQK7psZ
I/vbL4F3O+NEknGNP0UvLjcOMCivHpbioOGGqXYlpYre4G58TSzQzyU70MloUnx/fkW8o+yQQyyH
G0Z8LOKq1gSUr04X8kQQckyM4Xk4j9gEDTxZzr/nGO6xTe1/pQ3pXxxsQyoCrHOFmS6ezGsbasLF
KXMyALt+rvvNYoza7PzBwgjsJmSIHd0y+CsrEYAsE8Y2Mi1B9dI7cI0GHKRcfgqoCXhfZOX0q3mV
BZyyUktZyamW1rOleduaV8GSljwLNklM1FpgIzUk8SATdAuHQBuqrIpon+AhI6L57ngRCtIytxVV
R1kqwGQiYwySn7MSn65Y7fkPzP8TDzrreJ176gYbiLuSGtllPowVIfN+uhT/CAwGt7xQqUIlb0z+
Xa4aaGvTOb+8d2eZvH7ejnD5YCXmsfXptbTfWCao3pLpMbi5q8f4UK3wM5FzAFBBier3Q6xT/5F8
vp3yePDgRVV9OZxcmdCJtlxhZe+S7hVPhP1vq4iFFqHOaG6hjyuJ7ViZtiTMXxnYCLVhSLBBzWnI
hiN3F+l21FCU13+vR3h1PbolzNaZ+BLnFNKqFe59wqZbvZZT1tfjpEEIp6H0gC0ny5tUuyJLLNOL
NgGq4Mdmae/ZHgxSl8fRkbxyApTmCg2nRQFOyXB1em1hc2zjxQWHpHHkv/FJHl2PFQ/ZrOoDfmGG
5A+10FDo924VYqvw29guAle9GLxtEd/r4+SRnxTbBpQDY482q8ZDN3J8OdHSwKTJvDmPnE64hGAk
wgcch8HpDuYPrHoLZVlzYRk3T3II4pZQT0m5l98+GMgCQFJ6JuhlIJDfkbVp9mFTR7HVe2A4oEv7
FCgqb3bJt0CWTung63wMHLJrx7+deu0x1F/KKqgwawtYW62c2+eeCaGoBOy6J7Z2F9pKF854eQYF
Rd6XAw95ddUpZNFa1UPLw1M8r7lD5tskGnS/7zRj+rdzKtqPFjic8ImI+buBoJp5qyy1qj/aJMtA
zQ/moXQJNXjBPriCjRGW1yhYnzoR+qdLtJH0zRppD2gY6KM661WFw2Kh+7A7iK0oPvehTHm+9BWW
DngkJdTpdxslkhyrVX5soyslVyI83AGCD7D5L5i8Kc9pNP9Ic5RfVOysZ0YiLQhWntZ/NI9w0bgr
9+K3bT8iqhZYqJmPJWHNGtASpL8n7TI43ujOeFjAalKHiOtsjmVXHElbX/3uM3Xpfdf9Hj87urh9
nWMBdgQ6LYXJxhGD8dAZag17wmYfpqyoefi/NkcKyPrdpNccZhhzgynjHwLKdsxGxlGTcWtuDb01
753MRnSsxJZxBS0Pug2spgXPnlm+WHwGNT6TFCrGycmEEz+rFveDDG0xubfm+A2nACEU2oV27cBw
zpGqNh/cAWY1SU3A9R2KIt9WnxTf/6RZCsJ2cKYpYEi9zFeoJMmrWi1nRiI+KOMZqTkLhhweHtg/
VLtRDaH4hDd2whJLD/JNP62J1k2GCUr3fxhU8pAsGnSaNXsPWU2NocJYKqy79Lv3GqjZhrbyh0c3
JJQl99Xqtg6xQqO05uQYLwFyW8PHb4bFiy3VApNb6cDnsTxmjQ04bPrTk1JgdTwGgZXHxoZm8n6t
IgFKrmKW+g3E09hVb57JoqH7h2aFcYVqdFEF/JN9TMGuOyu7MowZSzEMd11Pp3hrufg1GNspjm1/
uN/GqJdcvwraxQXLDnTstBFSgIsBJPrIuh9qJwgQu3j89F/VzOtBLnI21X1wJmUGYWuMCFtaHRYZ
NuAf58UxnexH9tHgRpGexb56QnCYGU/4BzHfLcwaUsFfsP7EU/S2Q5GeAfhca2e82NjMjBVx+KtD
z66dKLa4yOFl1poSWOMlFNWEdLpxtoBBr4nA/i+6b66XOWESg++gnEF83JoFTQzoU05g281weRDU
SChzG4A5rDGrQ3ZkzwuTKp2+uFHFBu2nT5H00kwzo0CYPToumI0MiPNtBGJ2+RqVNxx/LxIaWylD
mZm6vY0BUCvvKbG1JtFK/7beVy8Qb1+1PHzdd9d/5JCPf02SynIXXxk/XdLuXjj00IlYlxEcKVOy
detNaCcQAqvBxaLskxq6roblLc+1h5xy5lEqpfeyIisy7aexMtx92jDcp+g4/H9mZR4fHpK9nKmX
aumipOb9BDDCizWuudrSj6R0CqA722brYiHJvZm3JFU+prUXQqMrRwFfYfdwz4nusUu1/bcYsmKq
rUmMAf5ztZVdSUmIhIOelf3d06OzpMXSAF8k/7h9pecQ4rZJs+7m6+qsRpKCtHoaT951uCWU4Kfe
gc2mvkcT8nohe+CW5hu9n7RI5JtCLjatXIfW6VK1OE+4+Uc2olzlxXEMahfEzWUYKvSkZBcIJQ78
4iezaAv4U2S2C1ajLd45aeZx9f1GLUzgaFvn9LpFrf37RHijE3plXhhxII0Hj2FiZ8COV78tSqX8
0+nEtO38VRXBw6HNBdESDNrrK//V1FQbk9peR5GDCuSkbNyFIGDoY/duRvPBTMv51jKyN90pTMT/
bvno+kqz6jyXgH763Bx+KQgSJ4C0EmdIt/dSSoyZNH6nvxX/pt51mqEkWBRbD2dUrdOtc5OW1ap4
RMD1wvuuB8+pF491pibbwIQH+OZO/8iDDEqiRDuMUWnK2QE2he55iONfBKH9SqYqSO2HQH8TQFg+
r22l/R8l1oVYXEx/NIvSr1PRfZlsPZi+nUHM4K3UgmcsGyIf9Ao7dj4o7ARK4WRCFBOhRoCpYifh
irjp7nbW6LBze/CfjfbtF0pW3GA9tH3D97w+U2LwUZOd9YP345MOd7yCRwJk45o1hIvY40ocAUf/
KAZzmQL/2fljtwwZsXl5vv0NlJj+t68vPhVX6GQBozuGFWhWp9HAcksQYZ6EGock0FoVH+HjfkCj
LxTn98o5/4MzHTjadOWA+6h055omdUaIssYbGtc6IcZVUvS0vTyhjWNuS8g6eMU4k/Q2/hSCjGkD
e835bp8+mnmP6ykb3z70DIHbCQ+NcnSlCqk2RRG3szEdVPGUfqYyc7ta5bngWgSnjIgIFU3n5hxl
bNm6iCOVDhypsLulGAZ3KOSowLPwrey08ggFa3IF0wr3MvKwyI3jCAPzEMKvxdCEnHyNyUZcusZX
HAogoiByKxBZHe33mL4hmfdP7pxqwYNTR+1jIagiABMk5THCxvfTbEK2hh2J0Dh+IyXzz2+YWDHf
dbMavz9HewS9IzIf+JEPpi+CfLh5kFcdvrHqNR6hVS+HDL6boCip1ax53kDAGDGxsABqM96Vt9Yj
dXJ7vMnqOP0BHTKe4iocJcXxaY9bgYO6rbvRU9qYoEo1+5817ExYCJ5bPbpCJbpAb3y0cYDyoHGQ
bhp/+2jbq7RFCTxFi2qPGBuXLqPd8wwq+wqQfe/Ub77r7STpm7IrypEpr2RFLD0261qY0e+F+wol
+xwIktpH1b43K1lWlwDYg57fcvCTR7pjxERoT60Zm7lmN8U6XHmrGK8oIz1XHRPMNUfck25RgoFP
KeXgkw9Z68tgGkBMQ2ALAUIuRz9eYTBl4VeOk+tf0NDUz1dLGCXPwYP09kFZL+uCmS62UOhvjSU5
/3aYPOJhfeJr+9L72Jhfk2jC2VxJ83AeF3syptYm7aC4Hy5j/p75+G34ks9eZnd+QQisCdlWSJB6
+S8zV8NhT8DtDjblgRfYLxhSSogFR4tUVBRaBEe3njiG7M6whCmg9EJHzshVmc4oNZFvgIfu5lJY
V+qqb3mhpKhKTezePqy09zD9EclLhxZ3SdoufYeEQ94kPg8CzQ/2Jh9tHukaLVmHP/cSWnYXnp8D
W89qCmqYcIQ1cpfE8WdRZNjyVDp8YLzu6QuaYjJHLbTELbielo91kXxYNFtfmwVWho/sE1An0h/k
EKRf0O0YKbPApIkVGIXl3DC8AW9pdBvvgYXwkWkpRpFSv/KVAtBbxaMvz1IiuMGKFoeUsbIcu578
jjaI/+LtBiW5Olg42U6MuyJRfcAlCJ4wzU959ECHo11ssE77y0yQSs/FEhIQ38Ay9daXQIIPhOFr
hjlBkxIiS84Njed4hBzw/XyrkSiP/SM31VJmvZ0T8/JZHFluQDtqp9QtKlEpJHsBYxkp9OjTZvkT
iPctWMoOHaTT9SVeXxSvmJULKZnm+e7CCRkqPzvZvgyzr+DnRLRGhm3TL/+RfzfXncLR4jnhp0JU
PIciSf2M3IArj6WtvdRnGal8nx+/U0QgYJNRTaGJaBP9RGGJoZa98Cciq06qabaumgRS93cA9ux9
n1ZPH8dTYXx4pMcGit+/2Rz9b0oBKJyH1kCwqTlvQjuYAaw9lbV4bmonJqY2fNdfD02qLqbZlE0L
t10c2Ml82hXm/+h5y7o6kqSTYn20kUsTv3K3s8l4ivZbnLXoP4dkuh6x9E+LuhUuPAu63c0kTXXx
fA3OAI8+qD+B4s+wBLTW3XcnWSAQQ0/IYgfRdrN07/NCFSjTSk3NlOj0EoNdRgetySh3SzzC/AZJ
6yKt06Fwwbp117FvgRaU/u2aDBVpFRS0ngw+q5AWqgKrwNR/oR+U5R3QiMU+d/p1xKBTBP/Qujnn
9vRAl0JkUstvkuowkNwT68boo+FNSW3xxMl2kXqnE+qSt9rhgx0ZclkAePPwOJscqegpUDkBYNwe
wuEU4V1ncphlzPZLvuXqiyrLQmMiP7wdcZj/qzbI0WJFzU/k4/MwapYmjfG1mxucdrc2uvCfw0NP
iPpBOXoGs8uwchHniX5TYZkIkUYTvWZtTe96MGWAzwC4quIRUF6WJG8BSjLw+1TEowCN+URn/gc+
SuWcPPSi9YA2JQmea7zeWhCrslwVfkSZtT6MXqfuYjJGEu3AxRtu0GGyZkev3whM/d1hj3grs8Ce
5t4K0cIyby++K2EjWkJHb80GomZfu2OAYI8GEaIcfryffRxbqqWndQvm9K6998jo0vhxlWraMwqh
X/hok+QeDzIgZFQofNgL7amNIRpeVPevhnqZV91Q6CmEXjrwQlnT6bxWxMqh3AlnFO+fwS+2CsgL
aog2RNjPTUxmnJ89uFvOBcRgCUC5U/MXJDMpbhDA32CfOOeSHOe/aO7JXT7QYN9hWLtm1SES55e5
bOqnfatOdOMcBU3s4WrilTQhK3EcH1KtwwPs918N4ryreKcG95CfA9aEw19PrSdsXZRIZ5iymFkr
Pvyo4PTNTcwo20Be/Z0ocbmiHDdFiEWLmHtL9b2GwpFb9gHEVjG9hPsVzallgmyCvsJpApQIqeVT
zHhClsl1p+mpwJ8UuqUPlRa9zJdSGzTPmORu1HNshcLsD9edWnVDBHloZHUIGE3/6CqTY4YCgEts
c0/lEh98JM/o4UEDlINw0ZIdeAdRn5fTs3rpCP4ruzRAKh5BsgvqMmqkrAJBqrZ7PQyoKQih4Wky
f6+0AOGFvW9s0E9POyaJ6jXS10gyygh6P9/aC8aO1kTVy/hVSeRrSaGIWkcuX31V7jp8rGQkm7mC
F9hqGnfaSw3GIUtJVeEPq6J3qx1ETD75L6Lnzl6zfansJGSzzomT9mUcV937wGLJRAgxMTnHuV1Q
7+qpj9yXoVW/mdzVx2l6QqiQpqSEWf7Od6jPCIsKY5ccIhwnl7BVHzBB/3jKwlHpunNK7zyqUXx9
hNVS2kLklF3JYZrzkGYbHnwVlupscGkEBP6fLeELoHdrOBcMlOL6QmMzp9+rrzS5cVOrgoZa2J+d
jqQSdrBL3jQqTmO0UHBIORPQrWyj3eoXpD2Phn8gVGvoNjUuFJKhHGldUHr0DngD73WWYJJhstVM
HRWrBawKHNZuv3kzq1sRywjijIdfscAkxlsTi6RBCKUgPutNY9f+2MIjgF9neq/Hc60pBrgQE+yU
lQzZnv0QG8s9H7ieG/2pR+vVFcPA4KYtsZPa8NY6al5ZE2AUJL6Zf06sgys2HyVEOYslKQzQW11s
4Z8/gmUC5wRDSAAZMQg4qRaN3IKtkCkD2HMXqjkEqkYqGu3bc2NnfcH/hUF1+Cv8d3fpD4E7vdMe
dMnE6XQRYTxfH8l9n1vdQcS4+PR6/vDYoaSm0r25prGmM9U6ru3klHmbHoCIgz20qU+wGimk65Bi
plz8BtEH4iti+swmhnLSJaagz1c0nTbuKaKu3uzrB+SEgznnDDJp4rNrFcG7YyzAOaaM46aHOt9m
9enJbRC7zXylZVJcHkKiCfRQ0xMMOnEts5e+RBjJlM4kf+XhFzmhXRlTyyCwy6hEXsT/rlIEofOf
CU6wP2eT0WHyQCPDAemDj0ROsVsBfNK+g2BFAtH15tCHJJLalHYBm9qtstxUweCiGO2gEzz3AYpR
ggOfAW4p7Jy2XU3jji4U3FWjFGKRouHkAkRfnAE+23pL0gLRay1ESzTXE53f7XwTP5xrPDH9yE/g
lEBQoynVxDMcbjZ5xsoL84a/2mjbEXRTm9PWs2sqkOSdi/2fDuyjKL+FO3mlyxUly0xyLDya42Xj
4wBoP8QQyRSsQpr2cHcGngSlat1EjBCicw8EKCw8BHI5rfZRmNtZ7RSd488mReD8Wms3ZdGukQK5
LE0brij/aXRc7yKZgnV/Od06z3IfgPOZ6MCxEiFf7iezUBg/9Qnlw7c2ChX/jUI0DTP+nG6vzkTT
XxdciM7XX8CAYCuPZaQI0S5IO/i8mj3/cz6wWWAlV2U4NbmAgmT/LsEuBZMTN2kf7hGx09Zay7F5
dXjzaPoo+VUynapaehtG8n05sJuV2YZfH+4c5ok7I8acEc44s/ejrPclSVvT6sE3EeLqnjOnHHBg
+JwMdy5fS3TN8hVXwRu1iggarnb63ZODR9GxTiBRTQ7HdnI8sQY8Dkr/5oc6VYi8L5c7ItM/fdoS
v8yBS5gq15/Pcl9jy3mn6MHhmK0wvlf0gwiUyR3wHI0tJdV3PX+OHb3KNONvvezEmB0Oqq6TVotv
htCzdcaj9N9dYXCC18vd0KErMwh4UXr3AApUDq3XBZ1rtI7S2TiyuLepPKSDleztI3Eo83IS1UXe
6V4mJcjy8mu1gRh0o7a0SRjANGw/+zCLAkvsOczRlYoHDjgbkrJvluAZCzEiqYvkZ17CxIpKrIlb
75n2sAB96mGUzQFy70oUWB66GQGoowCuvLgyia710le+lNoHd+bWPGnjNfKIXj/Dzua20kPyNMAI
l+etvBmE3UWGeAfHqOC+YkQaoF/zhU+yG6qtHXK+tKTGgUMKyY210f9/TnRxH0dmKR4R4hluoYM1
x8ONGjIA/uKXqE15sFccDCCXCWVcHQVukGTWFZhUDbtYEOzJF3YL2i1w0MCaUeTuqeHtorqzPbxJ
U+4W5zyHvv9JTgNwHedSicfg7rzowhI+7h1mOn+sXiK3S7+gO4p11F8EMtvsymT1qQJl0RpWN78Z
T2HnfijITPGueJ21GyIAIKD+Px+3cnyi/+MOkjh3+LZx6hnOlazGOEtfEkrnmjl+AbCJvYoFgmhF
mzCerLuBmRqfxyJ1N3Du5jlJKnZ912v5y4+Wn7LVodrrNnkVcxxL11YKRaf/KTNMtmbvjikabGav
GJyQ0F0WLFpRMECMxGoQXgaRbrYC5E/IOkCMnEt3SdVWA13njZsGEXuXRDwm0pSTRn4kcqzM7X9P
FL7n6hC8PsDvvfkHKcJwD9qZnTY0vGKpBbn0el1aYcNrgi6wOprIHixkrZLriHe854zeeXMzwcyg
NIeBG7MKHU8Ss1DFrzah9exV+iDI9+WWNGC2D7SSQj706j2InpMTU1AhZ5Fifls6vZ2wjJi5Rd5f
8syem86fhPGLGgz+8mATr9OxqiTpNQ8sHJpb1eCMGNSUU1dFVg0dfLyVcUy/ChadKYBP0GVWx5iG
puqSZu6RojqoAd0d35eirYgUA7ZRQQqDudEgvyfqlD1heIU9gk+qF7s9/ZXUMuF+cSnfP3Gb0YR+
5VnQgFX13rfx3nA0iJ4mGN5FBlek2XnT6HCcPIDyuOfU46eVz6QjjuQlWF1UdkG6nLvsP0TiQ5+x
FFdHCBEZynBPQe6iwcbaWOARyN9VKxK7ueuBep+BsJg7jS5TcaPShieEKsSjGCEgxWGlnEQYaUDI
NchVvxwYgyAInDKpMrhCvok19mlxuxQyEvRU1Gi46IdCsGQq6QOxcsmAW1eGsCe+r0+VD89uWknQ
JFs1qU6i+DMXAss5xPx5CNbatCeux9+eENkNe6tOu7Iu+SkvDmvkdhQIqlKz6w2uknJj5NEHtGiQ
5lS3esxDrtz7HpxSgDzombP62OBTOW52pvg5dxXqMZYTYUrkYE1Y/+ip0fZZBu3FmJaqzvLR8dRb
7ryb1CuTXelawE6IVEwyOZBOLtcTKiAwLfi1O1Hm0TPpkMpo2ydyjRUBysKykGLAfdMdS15i+40/
OJx1oUFIh1W75uz8yj/Ro6S/5UEla6MQ6b4Ji46kZHxk9DRbb6VQkNoWZwX20DpDplf59YnSbviA
QlBGjxlCwB1pdobjwGSaeLvSJCjejEA7BKCfJdLFlqUzSxh+mDGgfwaEH18p+jL/zuGMwcv6V2GQ
z4MePaZH5mkMdQ7PzI0aKAII/sS2J9hu0WEbLSnTQ5+/ggvFTNhmha7hUPSjdfzu0YQg9Ow+jzcw
fnQgGLk5e7ULi9Ot/24AV9ZGljgHKvzH2MY4cobUL13Jb850dj8FSy0npXToQDJxkIHmogYUBp8B
ArMfAsBjfI/iPLX39kwqy1Ly0yb72jOWmwkgOO3jsrUqRVWgvQx5KYePoiZdiR/MKf1A+IBMpQWj
8HC9MqPqn/iqiOsqsCLs8r/MMUYUwYRJrm7qMDj6ztKGuwDx26o1fQAGXwe7ArxSKZgnEAdQFxIg
Fta/fYEQ/og7MybopCQhvNQuHa89PQQiGkoZLn3hrRrilThB8JvR8o6syK5vEEYpdoZzRYYwWiFK
gG2TSEAvR1Q6DV+YSuFmFlx9HQj1isc1y2sKMHly+wBH50U3WnTg1U/RBHzuAHiPcr45wH4l6BAd
/XfCdhsuIifMTowQ7140A3QEDB+YOr7nuE1OivYNoVAcQXSGse/gQJlZ6wBbLu4ZWT3KEEYlrTjm
L8qn2490ISgcivwKXBoAbn8F7LtFVBm7poqPIGpvf/xuIlUzfz3B20C0ncgaZxV3eQmpDbuGHPuH
Vmu4YnjCdaGNCWeTxQEc1dQJfW8dH79xbY06SKbMGxUsabYiobQMc7FSEj6PdhUTgnWdF5vAscwl
9EZ/pYRCgmL8zIoXt+D6PhIQAe+n8xVS0XPPJIaCPedcw/PtNrQVvcjskDACJ2e9PwLwWerd5Fwv
C6tjRMTqaqL3G9GIuq8iVz7gui8WqCE30Txbp8bjGh5WrrpOLIbZGjQ5rS9SdANleYwAgNT8AeJt
Zuszm0l/5nKqbDrHtLqSDcBfUXSYC4dkXqxnKflbORipHRXgGDiaLFWOGQqsnZlSvSN2tzaGfkuc
JggGJwJYU/+sCBNfPJc9Ivr7u/57VB32lb3p9rKZbpIDaIRKl74KzVVPidmxhAfgFmQNCQ5pKmBa
c68raPfbHIhg2GiXsrur0x/VBh0r92zN4EVIEcQQJ24kidyPxi2YMmrS/kaKPph22DCVliLrvnG8
FlIFodRi8Rm2yPBgnK6JmpXFrBe2DBkoeAZ5SZ7HBurNaAVTeR5TlFVMDufTU5lzLw/bsrYGwLxq
BQEemBMd8lRzOfA9VfN3+X09WvA7kW1dzf0BZ4JWNNicGqn4RLUsdZZns9r3WEmseY6HWkpr4cEm
lsUtEMagOR7NQ9z3Nq44GQtGwq2Ou6TwJA7RFW4dYQ2DzfG3MA+8Eoa1RSg/K3E6umybUiYa0f8s
zTcbA/VDLdXjzIdzE4IjexQZsOsfiCuBs3sCCHj2oNesW1vN1LSCGzj+SN/PdBtf3Lg8fx0MUpFk
OHhzxk1CdQUVqUsxN1zkwykCfubq6mAKpDtNRXs+YsQniaGHGt1WdhWECRd+s0+TEPPpD6yCNSZ6
FPP31liNUfsXb5xEVFOazXgLmqlxpOpOct75UPjCDTOiTw0Xzq3Lod9VxUq5fdunDbxjIfQ/op4S
yRvmuXGb/jhz4qe+2xe8PegdVISLQpTDQHsIkRV6lXlAb6m7Rptzh+c+y4ohNmRWgxGhcUIeOW8z
HdaMHTexy+nJbblMU9yKwQGBGaOOQXC+7ZTjWC2WeWr7khuEDWfycfghmIy8mafiETNWg5u7s7zb
ofB/36wAICLjqWp61UUXP0B6LjHEu4QUNqjGvSGRMjOWVO9WYLCTVpTnmZEjtiYq8WhC58G2NlCX
IjpX5Llg8US2T5wkmNbCxcIAgiWo3MGOzJZ1FP8gsVyiqs3LF2BjVSo+aregL9xvRhMTW2LbOxiH
AVjBjhXwopMm17BnyUplINCX9cccAzt4SxfL9K++ERmT3j2/Zy1qABnOCEC9KDcM+XZ2jfllV1yJ
5HwJMcO8yqAC73BFTprWCFyBQ7wu9guQ6EpK8KcVq2B4F1BIEe+rkweiLmXYLwoNzNOyZY5m3mLl
aOxBF7zqnp+Q1QSgufnL2b4R+L9opdhRQLRknETPRzy3fLuUb4cYtUUbC783LkNzUtbSNt//5aBk
ELAEvKadf6LibbrI8IPOjUEzOfDYeov1WhSpovHhKwqRRbUtGF5s63RiRpwf7aNW5+3sVMnkfGvy
SM/3MgZn30UhOwZDq3XhiEa7Zrhzq4ONC/1JwTjxQWBo/6U/GMrlNKJtmc7XfQX3o0niH4FzoXnW
zkT424rVU2lHDkaiSKv+cGxh5FX9wi+NfyHGUNbSehFMZQqY6uoUDhvl/ygbgdgF8lPQhxLr+4WQ
HX3NOT6Wj2tRfIyOiz342YLpaxAN4PQT5iawdrJuKDFsKheQ264l1cQ/XIHF85BWlijkNs0V8GNc
co1KMUQG3SPKMa2rIMN4iWTWP0EgweUFg38v7LwaFiFl+wnzZqLOx74PdKHrrBHsBvP8zUpjIRah
I1evIqDyyCBX/6nO7I5cQHUf8wlPlYe7rCS5zASA/GLesj7/Gwu9g5/sjOwIrg3DbMs+YMUBW0/X
xsahrZ3uPmjx3IrlLng0Se+zG0EhXIw9WvrTtRoQ/eEBs9n6gjM7hphIvMMZWgMSHBqjG0Gcsfw2
rnM97Y+3MiZh8LEHjiKT+BJbfvW72ml5a30P3q1PvevZoGIIuxE9OfqPSpnuZs1i3PQiuGbSY9Gp
NUUP/8+V3wla6BucbmQN0/pUlILYasAj4q8tA+324IHa9BNOhdkY5h3thiI6OQKibR5u1ia3TdIv
X42Kj3MIB8RIkKBwoON5u2pB+b7mdPvzqTkBN1dH90uOpFI0sweQ1c3pBLocTNIVtO1IvTXd9n1k
XeIwwN/edm6lTgZbye7NHKzX5AGg9LJfCe4MVaD7OXA2F5ysPDC/r3l/EXPNGR/YhaYnUwKkmj9i
oeFN9d6qYPHE7n3KCipV9AydPInSCyAx7NuRF4DAkLKtJd+h7R9jY9WLmOyLu8Y380yeVTdwDAfp
yap9EpO3igmSqzn2ugkGHYOGqBsZTb3F8gfE3QN4UMT2OF+cm+TzuKQYvt2n79K9NNxCtK+W5KIE
WYuKZ3F9isvssge7lu0TwHtzNKSvvTdMpYC3Bd2mrGAtg9CKcQwi2I7Kxb2w3boRauTTXvNPLcnC
0qHGirs4iqmg5jLM30S/JEVVaRm4FRQi7XxJrrp6hVQ9+L6/JKx+EsJp/wdfHOsL8ZTx6ChqCdGW
efCkMyYC4Orka3eJZbgdGPstCZO7Aon18FBJk5cHAuGrCDFsX7nm3lOvMDcpe6pAn3OxFG+M7EvJ
Pl0lLfFHujbdVYtytE2WzNzhS9d+zG/gC9jSYJMaXIev4Usq3PcmOxapntq/q5kaXu080HWLNlbZ
02R6HryW4XGXQsZehPMMZjubNCrfGhlwjzYYOc5pC1+2HMXX0rkCBoVr7SpaJLM9R4ESjtwEf4cG
g3X9iaw66jQSMlV8WBltNMza47LQmIQt5fSqFSIkfQQZEDqIUmVzbPbM9nU5CgyBR+ylVyO0sKBg
cb00FAo+yhIhpnypDQLm9OtDKJnTUSmoN7EEAhQl2WqVuoMqtZiNWRxLMspSMHbnyGXoFdj225me
vrgtS6kWeaponN1sli+qw0tdRhml90OIMd26wwFgh4KCLUzBnLzs3UxM2+CF6TmNU2mjqSDzfCeS
Adeq+4pc1h+LkFAqZnnwTRJk0GisaCh2EiU2cEFm/Zf6fE8WsfRmTI0kREaIrYXTc8MWw+TmlSU6
p1zJ1Mj5JM8VgTtXSTn6mAmslzYFdttdG/E5COpe6CDfqHcsd4lYuGcmxWQrZS07HTiQt9loEKQ2
XYBMbpJvc8RaM2+jXGQWmRPTMCrYVTNavClmGx5V+jpGUHDzkV+2giNdRufd36G+aiKKwZFTWRxd
Pi3FxqBqQpKMsjbN5P6iOo08+hOOICphXEXlu+BbdM3z0csYCvCy+HvIUW9SUMHNjfc+J+b8iZXO
T54GK5IFkek+L/SoXSTESP86lP7qsNfQEOubDUVM2/emYU/JhwMrrqpwi1g/noD+CvEC69QDaCV7
zAvkdJ5c9qW2yiME0Btlnw+dZ5tJMmdnkbFg/eThROCjsXIqYy528rYLr8IRavQVCsnXtWG9a5nY
pmy1BnAUeS54sTrB2724NMLNOLNgNuHU0N9GqWfpfNoG8DNSUL31UmlSv1H520w5ViTFGEWQ9CDL
SEWsEfvoMy2t7hmjTcFR2Y88UwI0cBDiUkcqtFZGEPeiR0KhMfRjzA4Qkf+c8yDK3cxrla4iQAfo
o1yto7nu7FHJmsemLTjdx2mjMYzNJ2b5f1xke28E239+Sqs2B9VOdVK0ep2D3lPup4a43s01XJGN
gMyfmBTorjqtf7n+QMAJAy0PeZTb7tx9xFC5TGqjPf2nszpehYVPO10wv8ygSj5P627h6MP2KFHs
Tl36vRkl83teJr3jXUnbcPp5+CyZOLgiPZdVej9KTH0cxMQFxbpOyklSr7VcEoqSfziAS6j/bEgk
vOKWL4B2hdwOySMn4yk/hUdm8zzwj5fvgeAf/zkM72pkf+8ljCDq9oDaRvSUceAxO8Ew6TO0D8Mp
CdqEb2ARDgsX2cQKfTEnFkAKi+j3W33+xtbs0GhDXFFIyvExE51wWGo+bQTZZ8PRPljKHCmRFfaZ
eqhZ8lLJ1+1RoAt1itoNkvyA1d8UWaKGb84LZnn/pPxdLRipFYc+p3PoBGaJOdOCULmz/MP9NgDK
RU9TU1cT24gpbKB/uSKwhKT9SVmhTs6PUK11wbDkJpvfbX26OVsb789aVoHw+7Bn81IvAojGfcDt
GxOU5JC5i3Ug2kQiqtWGExjoDIoM++xUP0pAufEz/qkJft15Z0e73CkYv6Zox1SLXBuVI6XfuXJD
z+GiZuvManZ5kTtJev+pXqlMgl9iHoW0Klth07O6cromJCtfIfsGe3BUTcWYMBAq+Fi7CHlIzMip
qdc5Z5PjMonIsccGbpGBBj6K+xTF/97+ZMF3a0KWobx9OqMKRbyXJu08cKVJkmuAk+8jxC/arUpw
hhP/gQiXnlrStmp9aIZ4i7XHwq4Murw8/Ing8TcZuTE/BAGq8dOw4iHdEFqZ+2+NKgZCm+jByDci
9ikH48AmSJhWkA3y8GdDXv/w+MvJXhQdLnC8FZDmtP1dBAUnrYIcstUYJkG19EHjn6/DDu1AVeT/
nAoffvCwFzhh7n+VV86MeZZBP+Brldj+iM7ullu3MGbtIQDcv91HQ0HyeGs8nAIVDxmEWqu830Oe
kn2C7M8yfs5bQqp3cGGudQSVHgmQeUBhlwQxZvs9elN/evdNyYf5gdLO3oF/ZnC9KMlHGar/Qvxa
Sm7rV8T+z8jOaxepSDe/mGTntjJyofvoIljQVjE8MrBJYBDuw7Zx4YW6XkMW4bAoMs8EorDiBAHF
7oVR6NRipKQ7RC/9Gt41fsXbdYMBlme22WMafDhLY2vKCVADqztG5JdD2ZbxZYK+hlNKa9I9jMlr
bU5H9/VaJcsXyHU9jJgpYyifBPKEQyP/ShA1TJltwu/quc7+JawhQIFzbarDWPKUy3vN2GKtVxnU
OPRcYEYeQ5ewecKSQVRdk9orW+iPn+o8xSUY9wCXGaB9RMwJGgc3ERRiAHdsvd8klPc30H/ZeyRL
Jy0JFYsl0tt5gG4vVBzajucU3hTUxYwEf8rJ1EChWpodCMppf6eAHQWi8TDEtRXt1ifBHrAGhpHH
O2cfCXVs8ZQLgSzDX55j/c+P1tEM4z0Mr8UXOf28HK2GcODSb4CokvQW1K0uCp5JNb/U7bMQRUqy
M5EknLXb8OSYcd/TP3VCyC6d6i2S5sJ4ZVFyDg0hM8RsA6ZfgltUfEYhyw6gf+2/N2Bh93WHEqIr
/Fn441ZnAF/QmRPWURxoe512pQ7koPUg8qS7lDDovf4dfb2GjYmQm0ADhjiHwrHBDqM85nJiEfR7
dlHkbn6oLT/Dl4vfgdBSVPC4tQtm+8aviEibZiXo69IiIX8/f4GFgg4osO3ROSXk3NxTCMj0E9bA
8ALHiLjPTicAPKH5ZWuJND85+S5gyn7nEo0k5ykQwCJBfeXjKuA9XhVwUccaKiOE1n7exgeWYXOT
PRaSrDC8JV0ojyW53FQSLfZeV2ZficgGeMhP0Ban1dHjEZEHmLKZXolH1Iubeba1ozqlBBfaiSAj
qFP5EJ8P2I2QIA1ppxf+f53C/kJgfqNIa9gpLdC+6IOu8mc2N+dKIQ9UnQujDX9rQ6Ki0cTwsKEh
tAQeSZ5gzbo98brdUNu0xaBCfgIlm0VYlnkkbkHqEB4LqiRDNYO0YSCS/vyHFkA73tAE/BVWn/Hq
z17Tu6fdKzE/F8OR10+4408ck6fYmdnjy3FZ3L5yAuUUkk7awUWpPz+PfM+ho9iGBp24jpQhBQJl
oTQXp4rNtolJcambQpQOJde9j3MWHHJBiV378rPnka78DvBkPLCiEStU3OCnGYDA1XNoyOP41NC5
1nj+JxpX8uy/8DSu1FCXUdwuKuUjArYusaFnf8inTQdH9b6/l3mraPO26Uh4z6IvWFRNhqDszdi9
8bnNC3R4CXg0xzrVosNGiweOWKE5HjY8M329fCawRsiUPYom13l3IHh38dKYBaRrq816wY0wRA1/
R4E1Z7g4dyIGJ0+UG6go3ev8TufG8Co79JiFf+K4a3cvWF1m3QiZcsXaHdmjHa6x98eHNg0EsRh+
ILA7c94B2qvp8xuQChocxCq6gvA7aFP+PgGLVEsq7yArTcqT+K6VgOYOUNO9eAiFfDpNXJSbOwXl
CnvQyitqO98P7oSl2fWDBfxekXGabfYkq6hRhcpudwQpaDTPS5a9IIgNJ8RWq4fQDHbFabWf+nM+
W97dLUlLTlWRGJFG5glWy8H7ErvtSdL6E0uIq0pUv+o1EzPjG6gnurwkAWpS6K9x/7TCjK18ftod
+beIIJkaleF0ZkGaW5wujllFjpxVVsUV695rwlyicbXKODRY8RqCXtLxx3CEI9Q1taCZpTN82ebe
XLWKpT3+b6PCSrZxUsl4QiXvztdDHXCkfrjB2pS908leanubHbAhD2Q9yoKOFA/UXeoC3fhphvlL
VGnlozEmTyz0cw2wU4Hqq/iZMlTLcOwGh/2vFvDo8Y9IXRo4IB9GNQSyBMz3rPkOMzpHvJDx7FH+
9yZ9TNu8AAlWCkt6FxqpSPa2Y66kCT8WlYuXOyVawmhPyg7coRQJQ/5ihTxEud2fzYvkqWVBQyv6
c3VDHaRXYnwo/XtM9/GRQiHNb8a3lRMG+D4hVGoe4ukkIkyzyfFVMR/B9KaOSQ22rYAgywel9lhu
bZxXbH6q4HA65R+PN5JkHzoDq/DnKHZGahjPHdcEqI08MtlIBeJdpaI/j3R1CC3jtDoDdIF5cMIb
KD8N139eMpQBvjm7OHUXUHWi7GHp+YsfRIEqm/GWl/FoMmURI2vRtv0n6DkiNI1hod/DDuHP1Vm1
1IAA7wo+zjyVKROR0gZ0xIequUfll3QaaFwfET9nhqXIzv/m2OfWOp91vs95sDGAW4a/bsIEYEtB
Wqcr9SVPJz+Vf8ZGHRxu7hwjq6RogemIvZBQFM5VAYsIda4sCXGYCur+Uwk0SnKOl93o5fCVi2b2
rjl5E0EbcLkTldcOc7VHeqoFTcWjAYoMk1eKelgSIjVOVVj4AG+/NWnLY0GJRvLccHoLdtTK/U1W
OX+DbmBLP+nS9c0p+do7R7EwUOLVZJbOx/0JQ5RWoNMl6rZJskCx6E6L3jcvds8vwXw+KPiWQnhe
DKOz2J+Lv4s0y0lV6alYrMAL4fzmXtHuJBJwDwJT68/CrTMf3Td4gF5SGPv2RsM4jYqUDQlVZlT+
yqZYPsFre5GoQNTJphrhQirZbLsfimBNVvbZ3Sofbm9r88YofW/sK/fSjpueFL8VW73heNBFc4iJ
KbXsNUR9sfUoBfSoMbjs
`protect end_protected

