

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
iaGK4Vux1Zzm9gBS3KKNmBXNdPq+lSqE3Nnx40zW9JpQDS5U0+JlSB5O0czPvIZs1e6N9M3JonU6
/VRFISTQHQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
hnTIGD4PF052NtQspkoD0qYNWsnDfk/EZli95x6g3PoDiWDo2i9hfthnklZPOTwcwwB/on/PGVLy
LOGgor+yT4ZX8UGtoSmScYDFDjshoGWHhtXrHczoGSF01e42zFHCzF3p+Kqif4EYEFLVI0b3qWfo
JoBwVA5mSGa7z6eKZ08=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
jM4x3jcOa6ByCa1VWDPoU4L7JC2eupLAavYhTE4GTMYrnvE7xP73g8zjlwq1G8Zy1ODZ+0DDopVA
JY2gdvefh3SJisXvlbuH55643svFB8C9ZXe+EMovXErk8XGGsVfWZZ9248m2dlrUXREntbWGdORb
Fvho+MXYXuv0DV2DKImT+u2TQDacpvX5e8ltSYsMmjYxEdkZrVMF9C544bgDvuCE9PfD8XjA3SZW
m5oOMSMtDQabvtrFCxaEG4NyuxA648giN43WXdidnKPUkuB/HxDMEcw9NxHOVNuLeVs7mrwTNW8a
Y8nkGhyssdB7pA+UlWrXAfs2U9Wpi6SjK7D2dg==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
l1zDcM4+iGcttYyoR8HHgtSyP4Fiyy45WEsaODDzemrDXcJaURYpyLa2UgO2HmqSNgBK4XdlSO3S
QC2s2wdlVLq0nr6twxtavd0Mc90p3l2akMlkawzSfWC3lR7JsZexWZNEb6frZfXhesr8/8i8wphW
9oH5nUnhDJDdlXi2xk0=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
pHbCg0c3yWoABGhh+X5xmKdWu54K0QNaj8yiI7dbYcl0s74Nnt3O7DJj12bDcjZRfdRoiT43bXo4
30QPK3Jr7E41USUv0QfI981OyCHaIYD9DzkFx/42CQBEOSHNBrRTW/rge+4hugPE8z0ogrEZGdei
kB3oPw27BqROJcBQEhzDTOz6PP5L7SaiUGBsXkKo2TeQ1sLfd6VNm52eUhSewTFcPcdSylZU9gjA
/KlsPUnl2PskRWTiOzVvvy7q14ROz/8yTOqbBslSCNrDfBQA/bwCsE4HN784FAGU2BIu6GH0W9gV
ySlMw5kMiPDazI4NmLxMcJvTd4Vi8xnRt0T8Dg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5728)
`protect data_block
RYy68068/Wg0pdhvFTPIpzG+Q6wbpqdlkLF69oWOfrL67yuTfY8tiexkiMNLyxdxgkT2HOnK3l06
d+Esb4pQ+cPSOM3Inbwfq31SHl8YCsmt6aYiykx3hZh92a5eW6ZoX9zMPNd9Kf011oB/4PENVLYJ
/HR8ojcvDaCWZTD729xUGJx8kTJfnt85PAn5yaMJxPQAmqR2vH34IATMSnr1vZOt2bUyAA0jdUUg
d4d96blVU3ySuRjqYOfVW/VzjooMGc1y0uZ2MvR1T2sXVabMFqaMLz590P2dvYC2q9774A0at23y
xmNPGiUdNKr1S4yZmbbsRAJTRy716M6ITeQG7voN3rFxV79BuZZ2zfDZRUv2J2NGPmVkcgbxME5U
tcPA1a42yDDocuvKzxpcIxMyEb4bS9hIYC8m1WA2L8VfDKa4dq/0eayYQkOSBZhUq5ge9AmuaBY8
yaIXlKTNs3+qioDQILLKvrOdknGW+1K6e5rm55FfgfBjlkWi++SUq/p8x4Vw3CZ7CqOe69t19VZz
LPg3F1FzFhFAWakkdVj8IFAhuleUf3932G9bom/NlE2p3qojprx3YQbYwehANc1nCTuVaJP1Q+uZ
SVdPnYT+fA8mmZU3VCsS/E1GtzmCnkthaOzSop1n99Uw9tF6krM1hVytrupTTkdUeaXGLOh/H6Jh
RfZgsPIuPcakNrV7Mj1YVCdZB2ofafQ8lOPmY28jgvHsME7Xs7Hwh9wCkpZQXIlqaMOom9f7A8uq
fSAQBaaqf/FriSZIw7iJGGj/qNTS9Rsf4q9GvoiO1OHg5rvivHq/Ul152tcQ3Ig9HICMRiUXRXcr
xLtRzmSSoLq7SOTQvmneobt9sPu/j9MKBrtrSxwFhJZJc6skon6YIQQBmtB80Jh5bMaYf4CWPzGB
YBW0NtIcYLfnzZJq7JvXA59MORTv1MQkq6XVnDNzK+/xm0VvGrPNFDe1yQsfplzDXDszcGwxkXeD
BcgV8iUvnoTAPaWIle9qQ5laLkf80Y7aelYX1QMvOkPcl/zH+/ZEoamUhe1vS0Kx6pwaP/sPfdGG
TqSxSdn2fPEiCaRJ27OtgBxkn4wIdbTNOYaxxR8v16ScEvngj+hMzcxv6zZGgLXDkO2TAjY4pzom
5Skfefk4VHMYxHhG7tP1JCRK2ZVs1PExh99bNV3aGbGzI24e1xGPE7xo7JBPMOByNSGJd2DlBOEu
L09UcogTiI9VISthwnUBVPdCo9JHxHBEfOPMH50XshxXwZvpZKNVGjqVI6c5fowc5BbOdxGBed1F
+TYMjl9VjVyCkV7hUhPLgmg5q7SnJQSw0f98WOudZvZYPNJSGmcSPzneMHWpipj+7Na8lvcnZyjs
2NqAYad7WFYOMS0t9B6Y89Ii0KCwnGO3uBkLO+2AYZEcvgpfaHHs1z3o1pnrUV9Mu8SHsrDXThHW
7O6LIreYxTkVHQBKs6AFiSpqrApfVx7HXa+MfBwoKtfdtufrvJA0zl+JOK06oX1e5lpnaMiAvsY3
CRiXDDl/TBoCEyhxdLiqFsxyg73Xy1XHc0E4Mp3lE5h4cA8xAkIjmGCabx/AOnoKQvHiYDpn+nsO
SWXrYfZbIQzuaobzd6pdNqY8Ho+hUO65uOHA5gtZ85vhnXL3aatK33xQjCJKtyWNK7lhPmgP1ebh
hosNXuDgNuaLRt/Au1bkkv4n7iDUyaQ9A0IZV+fQU0tBHp/UQ4uJxhy9WmCGW14zaIGtf0m2Rknh
HU20RulkPbgVQ/Szr8/mTHYm/0v3R1qqQAXCfJgCyQVy9ihBQQUyYLCMzLwgTLI0vowN8kBOdOoG
atkgRr62Q7s048i6tAhXSMzdKz63bLP/En9Qjj9SvxGbWiZX1eRPqutJ17UhzX+oULtCG4f3vGuy
gORZHNZ7QdIslSYgYk7oSZLyXkNYNjzsBJreIkawJ0AtyVmAGa077z+/RfVHrTEghlgvtCgfUxIc
rVjrr5K97xUrEdPRfCov/l4QH3Pq6NWSE1anoknrjJFR99JYHfTkDDj8eKxobQuL1XxSaApvJJxn
UxEMlC5Au1/o13olW8U4ixsCNlbDdfPYJ+to5KE30o2IJ/ItE/6eL6Rd87SG6oaV7k3lWLSQ1fwk
08j8Jcf0TvNBgxf5PheHqFGegpjJs9UVsVueiMtRNJZFdl+3wCOrKy169Ur8zFMiRgoHY907Yg4R
n8yUVV+0qF2xicoGymD9/zzll9i2UmGcMuImYde+EdDOHQXtWjCSLXF/mhN9AI96cnkbeYIEnwLd
JrFLCbzgg0PdZ4f13OK9tRM0rtFmk3h3n5DTXDWfdXlH3GB5dbdKOW0+4lYTfcVUeohM8vzyWDyV
qS5jTuqL/qXvxqZBcOe9T79lPH2Quq8MiS2WNxrNmHu/+XcbVCHhCk7cVG1+k7/zy9hFu9QkA9Az
5NuRnaqZJHR7giQBQ7h1T3z6xMAzptc0+OJ/7H/EPz1iOvB88WnTuWc0izilnsZAdqZZAtxTf9ip
stgqm3yPNEHrBbBn6lCrf7bdQEs3S/QRWgbv7hF2Ck9roqP3o7k3sK2gaMw3fbnEjFdoAhlSr26U
pAl7Q/DAfrh+nCmibRymmRiIANUINLT51wNI1ThrC+ZQxKIjHfznfDK0Jp5S0skpZKhtDxgBt+p7
xdxpgGyQ27mJdCoi+42TZcDCHk3bpEq+Se08O+RY4BSD+0E/y9kfZXs1jTZa4Zp9OaQAjX9O9yJx
xwdGrne0yTB2WrRoO0W7Td6z6Oxb878qEgfSJ13ZlYkaB1WPV0cNQ9xCTI/nFN1Rp1S/TrJaShSI
XPX83gK6Nlv+vm/AaHMDzBoy7nLVQsSU5IagOp05DHOe4l6ocDtPenVsqeDpZWR+8ftCSA8ZJf7/
r7/i9Db10qBv9f9GiB14D5zHbV0/62HdYD4xT7zhP792NL4eAxx7+zIvMIb527IrDdZHXjNg/yTg
VK3gZPlq1nNW84z6iQfcgDS3vKzrAMCLGBD67ilF49PokZSUe1oHNxtWuRENUcoIVYgPLBsBk9l7
1fc2BGSgkWu8WaggJGvQW1rtogPX9KIPMwc5qKbRmyKT3GT5Q8suHcRFjvhilD/soQupWELJrO2g
fydhlr8WGQq+3AMBc3yORjGhODJsX5fwdoNigRukRFSzAhJr0vLZ+qrrWVHKYK5LFfOXPlA/navc
jR5Lx4HTzr9DKdzDhonTn1VnbNeY5ECH283nCHzMYZldrS/FIXnGV3uRq5FOr9AbydV/eJEFgFuA
4HbM2vO+aqCWPzuEUm+CH0KZKMhGcCGed/hisI6HDdYf9c1f9tH0jRBL87mTxljY192lKOqiCk40
sXavkXGCdCQwajwwKgI9Dx6HLcwwcPDSnDqh8WI+/vZjyQ9wHm8bRuYdVXwaVSLucabkgOgayVtD
OPxzQoKUjYFG7ZArv0bU9bLO12YST1EYMynFIW75sJNZfR8+5Zi1xKNQCTbwESacZbk7PBiJdH5z
E/jFuoGV3DkMwKDlf9btvkRRq4V15rAvT2OLWwVCFnFgZ0TJhNtuHrw3dvrG64MkBkSPGTW070Hd
P46imD4lNLp7CoLW+EofHTO1dd6ITuzXChrZTLrdku2xdBeDRRUPh357PGr7w5xLhSlZG7H/JA5z
gcVGB6NO9Ajv0Hd0XrjV8vrmnus9Xe+kRf81L2xabnQcrLVntjhCi6j72ir5DBDRF7PIQ3CmHEuc
afke2BBpaC20EnBb/fCn3OaOmzo8WW91u8S6EM0EG8Pfrc25JvCv/jbr/hjyhzAe3rgRvcjT0kG0
M/ceXI3SvdnBFfTRgmuf9dEGh0PwjqnfseUXAZ81fFrc5k5BaQVBBvCHQHdRGXx84G1k5Jq0Jolm
WcokNYJGbSBk9KnWYVbQc77adVioNzBLCZdzdnH+/OPHW/1ca5H+KTkUMDpSJ76Nx9FCAs42gT2r
DYG6CufuPUjl3gHK97vCUfLXVf8KNO1pp1ilzAVuKycbqOw86JX9neKXwavidc+pMy9EKMWw0mwf
U3xFPpZaALu6EBpNMeQCoBDYQBc1aTp8/mXVwl/CsXXYYvnQUvoDrIGMI+BwBKpMl7XrXhJwaTyT
2PMYC3MydavySvihoJJ1My8Y8kUiNvCT23WJdRP5FZaV9SZw4PeobOnXZur0M5bIPZFCdtQ1QiHs
LWQB7ydUr3Uf0Ud6vDzEtnur9H8hhesGtzjFGJCOcetXMc/0jsz+capFCOXHis0IhEdYB8ijdZ6w
FJgto32ocxBwgqSbkppW5JtCds5t3FCtXFtKarpsCzJGKJr5YRQ6YKml5UwiF3/p8z+RWk38tpPF
lbxSwZv2kTnTggcbEosJXw4IKS+UYJ6+ZXRa2JHLXm1STJ8KcuKqWX49lsoZSo5ngEd+6TxHu3gi
kjYtUnrQwaMpfBBIABLMcGDseE9wY3QY/mJR3VIG9SrPZynIy+1WQsK6fvMJ+5Q1/82+5U23MApD
S1NFdwxfYPDI1OC21GWFDvTKERQX5OaO/nhWnAOAQVJXDLgfr04lEZYy/dJAGBLaOw8ub+gN6WOq
BHWtejRZ3pno0pUPPMeRRsKzHn2RrjNXcDvZDjlCDW/Qm7OQsHHLCidHMqogjkTRTpn9sfDewAln
H1JZ7TE/A0J1dGpkmmR3rzohcblprfa/dHZuJah8sA0IzxevWasBW68dhbJ2Aw+o7ahAVyODReFB
NcE2AZyc+nJqstFc47fyRWL23HIV+ksAiS3t+99tzkD4iyTtpH3+Yt2SANbR4C7ezumZkNRuF+cE
uMnIE10MJgtXHye1RFrJJCSl6vttMXJM2Cus7Bp//TR3DED3/W0yuwjriJDBvCEbBBaWz/4Ciizx
tP7v5TcLDfOVs5UqeQfpKsSLX7+V6UNDJR6gcJ5q438LZBVfSc47bgOpFd+5LKOuEmQ1+F5L21Ev
EM7bKllM0CGy9eNlrbI5S48L1gmcXpm/qS4DShwoB6gPe5c5uCyqj9qYZIokvNzoIgEXWRnXCx0J
+dKVQWO8pLiHT9uSxAr7QNpbiWZFMnzTvbyIIiaQSqMc3ENgtERaAn5duHtZTQUcf+4gG1P9NneZ
Tw+n+sYT9RfO3qhzbQt6e0DhwVWb0xN3tJGbj0b7vK+m1PcmQDq052jcbCZ3vk0jc7qw6Jl/wFhS
1sNWbAqn/KqH7FX/wJDcjd0Rm6zt7wL5VSYpeIt+NK1m22fh6IifcK3U/pSq9onkw/csDGEPdkWt
U/D8+ZrLpxGsCmczzm/AJAoFSdq/6LqknHyGWfkAf+wj7OwNdHLVUN0chw0o3aa7E48EsVN03jJ3
lsCuEAkgkSirhfDxIl8sewuQXLweujpmt7uEasUhRHKZiNi3jDhVgtBLXgSRp8ty1c91DeAguaPF
ldjq4YaP7kGidqIx/dUVHIj4Rdi2NBZi1jFnkoeIfmWnDPKtHfWedHs9COvPkt8gb4d4evKojp7Q
YZcXMVewqZDAkJnGSm3JwQwUuHWhliesyX67tIJglaCAAz8b4Mfo13XJcvTCY/eTMbdyscOHhd9g
9IJTmL/I7TJbuT/WmdjLvzGHnnHIJ+5rDPZ1KsUySn2yf8SpdiaZqTCXkp8dpfqyELWa8EICtg10
GTlqKLhyiCkUogCF1cZ2FX25HMiJi3tdO3tDK8wA+3Zdga79NvtiCfwaPvk24YkEn9d7V2Z2ViGO
h2x7EjS4W85tGfhmEMmOdojbDREx/7bQJ8zAkhdPwGIZ9zkfP01YXW+KsM3bN1WdipBRHNxKmlPG
vO4dpTjFPi36TSPuWHybBmK6hTJD8yKdElsdPrGCaejfbMjtHDuMGWosqdt1YbBwssku3zpTymUi
Da+Znk1ZcTFyUPm6I5M+T2fP9BxcWuNIcYDZWRHDzpkWAfNKTcC6l3Z2qodZ+n9pebva8euBJup/
ddVnyaDkCqeMex4V4n39fI7VK/CXejRh5ahwbAMiCTyfUOr/nhZpL9gwhv6xwNX/afoliYhEU7hV
JG6w4UupF7XcAJhOWHvkSAp/+QRYAVG1a6OugF6nMyzJc2GY09yxhxgYFex6HuJE5+NDwmJ/hYiB
/sTzFgslSzXODgLjtAJmgMxk/5uYXVTLRyQJXvTyVQmYOVEwHGdaXwFKMfCo64V0ApK5rmSFzA2K
Bxvp9swpBF8d3CDH1yuKg3eEsWqVWD6cZYeS/xW8ZG9fx19mV0ZMPDf9zG2vkj3EtfAT/ttyYetb
iDHkmY/M620bZAfLfD7dQWJOaRGzC9KvzPx6YQCNUhaItyiydey4hIe1FSOyG+YvsnjU9Z49mV3m
kKrKGqqn8qgGk5sMSL6LYcW21ZZzaj1GcMPw2R4P/ch6IoQ/gaMWjzpnhKZhfHA/NRAaYcJLeuvR
sS+xKbvNuK/QyI/jpBM92i7GE4SsLcEzQqt950mJEYZ3jzDjVkrG618kITQot9bs+FTxJrigE/DT
Mmz1VeZ2J1EHDwJMO9Lf0lNxVQMLkG480KBsh/GH7b1L2YpwgKli7NI6uI6NtGKWTSPvy62QQjpf
fDeQnBu91+cpDwz7Vs5LhjkDKsxy4A98xlA4QFaxGCW95CBEnOPnTzgyJUrLbCinQ7uH4J69dcEZ
AF1OSsy65rsYZwHEzSxh1sNCSEDsT0MTEoa+OflZ+oDhwlPK+LwwQWT+q4nzqt3YGE+cw5Il1xTr
0fQ0Wu6HuNEtNgym9ykklA45+XuFytZP/8ZxlveCQy8YKH79tGSccqlCoWTat+M+IEQB4QgKlkIF
jFob+xPds/XfPvJxBsT1NFfsUkVIyUJL6vIGUS3x+TF3ChKFZLP3c+CbBluaPnSbq8Eb7d1stAR8
WYd59NyVrHAycZjyEbfM0oJkmk9m4837+yxPaN9ePZhye/QsOuKGJiVLoxJh6UZ/lSSiKgY8oRRD
HWa4RwmkO72flDfSjoTrZwHc/B6CINUIo8K0tHQ9R5/j4fWjWrJhlmzJUrVs4dWUxjSPcm8+ypmf
TdHpIuBcTPNr0/dbpTPaEjUwWXRAPs1ibkxHvKtRYv3ceWBiSkG7FX8vM4WmfZ2N6lIlByeLrHlw
Mc8oc11sb5o714Pu4haJIdoj3hAGfJliq71ijG7qZnRan3X4KDnngCBLUu6HI21ik3bKb/TB17fK
o7pUazIA5yoy8gcFWjp2Ov3k8trMAVgcpew1OoAjwqa4nv5nJTZ6nUREOqf1k91TqFq0IqsfG94g
amFomMbjFUlL6lGTYcR5j0gF/GbBFVgIvtJwRlqNvTZw2OJ8TrqnHeTVb59e7LfoAvdw4OK44frg
p3MT2CaCWzs/H/8GycJPjmHCgc9DfMCsXKFcyq6EXw1Jduw/jgAYRBAxhNKsZGQUbcnWZ77IoMsf
JbPOApRTzn1EXL0/h4Um1EjR4KmbBBxWOHtebIOika6YuHORLypA7u610n8Zrd4eHtm8STX/iDLp
toAnM3vv+DDtiztj6x8CdYrgpELZq2APNCFnD0v7bkn1G/NGUwC8iFCG1cMW0O7mqiUYo/MRg8Vq
LJm+yNfiGnNlShLh6PRUdExuWGbqYLZim7wfNYOpdQwWRX6XjiYOdNqHm4Y317PVmIDleoV0WHKX
Pbf1CSQ8m3gNAZ1JQxYttsQWopphLjBmVi+jPQ==
`protect end_protected

